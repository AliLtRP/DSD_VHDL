// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
HfzhNFS31lryHL0r/A0j1UIryzGhUyjFDk7rjpptIlulp/F1+3YNHKgHaHPRRt8Aro1F3XPtyAzz
KObM2hNtYoBh0fO9peJJH+kNmhk00byQe9Q1cxIT9P8sc1CVd/tbMctU6xeyZdRjaolqXttbGLqD
XlyNHhwvwDtufroJCR6expJ7WgcfIKzgSBJPzi/edNI1RTAVKcJNEM4XC2DP19NA73DUOeYwU1Eq
zsoQvcmUuOENbTZD/J6MSVHHjq6xZBt8AVFkeAfO4Rl6QJy8LBUmNw2OzqvxZgqmB8oqJWIiL5pt
PLE/jcdHVBFwUG6I1B47RL1/s+akjdtUUH97bQ==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
CxAf+ZkajMDKig+955Yf5Gk/tPY3IiGfE8NMthntK0v8AtWPzkoA1p2xU9O8qP8sM/L9t/m9Rv9Q
76RvktXCM8mnt8kgZvyqiWZGHrXeBos5Bb0QrdjsOScf2kgwUVdS9KLfin2WIrUr4OBUU91RYHsR
m8S4IfwRxNecYPXj1//oe6TVm6/ooulRYXti5awXTuc/rCnb9ygBGs3+rhJ/WTdqAeix6iNLRKcJ
d68u8IKaD8zUgb1rSbE9RIoDHudDyH7aZf2KZ91Zvs52c3EiQCppTdBCdphMsFY9zoOv91qAx2tl
O6f5HQWkdmVfvj1IBPTdNJbPPpyynr3xHV4/Myh7dirsi5Zo+1Z4lnHIwT2LVhq5w1XALWU69Ksp
V9KQI4Zq6V9pn439YxZ7XnPBe3zjTp0Qk4c2SJaVlreQvJNmwD6ybO7W2/8QA2ZZXqrCHbKj7VqI
OGSzZ8/IM7PfhbifuYrsx/EplnB5VcnweyDyoKX1L53NNLj7/YJ3Yk3/gN3jiH74TR+ls+uMHafp
QPtgy+PP9FYYz6EQRupVrPu3g1y14Qd/HqY2icaewRi3dJzi/wyHXXlibMALS7tkYrtL1DssR4WQ
tz48jBVfIJGHtMpj7LjrIW19LK1YAm+owctg/GV454tRkWFf/ZuI8Il1sWXGkzaA71ZpcG6Vl2MS
WcG/1osTv/CFatnXKgRARPr+qfzETb8xPrV0kh+eOGd3W/guhI0lebUEIEwXvxuo6QbQXTaaLjOp
tXhkDeqOwVH0xRgVYkccmOah9qDO97+Q9GEYt+ZooxeVCdfqoa6StGz7qEWIDD8G6UuJBOu+O/Dv
XpxKb91zk/h63IGA+cd1t9WqpMxgwpQfftui3D0V3I43QEkA9qOZEKVis1FMOz9hZMV/DdlfksdU
au7DNdzVyUEc3DnqyCqrg0LY4LECFAd0U9sS0Vpc0Es5/CUPA0m2E+l+7DPLE/A/aCJVXLaSujRd
zQ58nvo+sDT4GMq+AUZ8JMDt5aRJQbYLalNyRxHE2BhcGSQH8WhIrGBiljTzokrqtj8UDIUBNa0O
cjvPYKwkPY1pZrjTq3QOCB56BWoBzDGg1N60YidcfQp7NfFB49OOIy+yg6Y5Oy6bVaIRF9uudmEn
+mOJakQX0epLNVGiL7mU4BDjowaEorcTcwiHsWPfN8XvL9nT5vwcq3EN9pU9o7ynYx/7xqqPaCzZ
JwB0jaDM1bHNTXwlC2yhbXtboF6zc9vKeeohvZfZKDs/h5apWuLbeqC+VMoZDHiYZEFCP+dlScz7
KLfdAquElnvijsFEPqas4u6jfmBKIxW9oiSWbC2TNGtwOM+EKWDl899YuSpDFpN3tP1lAaeiyJLQ
+oy50PQdq0xvrCFBSinXme/HAMZJ1mM9gnR6WFJqZqMTkbfEtf/wZYFVQEQ7Donw0CnDKJOF0BK+
2wkIyNYTazj7O6NqeF9WvbDuoddfdcx32EWCiRWDYrM1PYNV/XugWtTZqrpjidfBYfsLIWP660dJ
baim9IE3Q9OYij+OgIIJEfz97QhqD4/fY1XI8orMhsX64UkfsKw5E/tJWQ2VbO+2SyIMgj4uP0lO
XNQy4uZDxsI+Ghexu6yUe83DPtaCGoIpM6C/FQLzlkLlzj1J3enXyQJ26bwthR7QxL/EVLOT2zEK
A3XfWhsVpJAlS75cGGQYyikF4GqtnQrJIbVGQ3tZsLyztlA+tM2lgyBXf8eXSbeMxpsd3FsYp6eW
nDkUr4F1E9GnyoKn4M0eVCHkeSbt0tXAcYGDugrU4m1YwtRzXujtFIoxLfWLaf56yXAEbBSKsUDp
NHEb2dunYw4J7Mo+gx+3V6ZQjXMaf5qsYjhi+9Gc8EPopHimmoXNCdzI6P4HXyqUPx3fBbtwmPbo
nQoZtNmI0E4nhUsoAhu4KtJvuZD3J5iXJmaE1Z8gSJ6dFeyAV77k/ynmQUZ01eblKx1kva++pvfj
Sf/W+sDQiDN67edlh6ASnomtAY/WtuTNM7PqiTfzAueH0NWldX+KFWKbtgPf9MtNdcx5HetAeC2c
ciZTjYwiSvEJ03vrp+uv4verVoynIXoVWL9XFl3RRUA4U/0/lKsCS1mwLB1XYsWgvbzLwkvs89Ly
5J82h32dZlEahIObaOoZhmAqE4dzUaibge/bHWZH4AOQJOQn0GcGD6afEawxIxuXkuhGeQPAgmeU
EKohe05H+irbj9EQ7rR8TGQPQp5DhU4iaNiD5D26jnBq4pagjACKgqK7DsUGUaUkVu/HCeSLQOX9
P0KMUe5Beir2hh4guBxtaXxyPAtHUgtgJUpqH6UHoOyy1yadRxhsb37mILWQ1bHR7cfrdkiDp/uM
twgGwjuAOx/fcxePQAu4Na32hHIGJA42ZEzA/sfI0mRzB1iKKGjhdCZo3SXH+xrSVKvEnmGhho67
tHYEwTGOtDWgyTiRVWtH/gj1B4GkfZclYz88Z4hucdKESHJ5CT2/ODgKZkD17M/qZM0OKYmVxwp+
AYsJe0FJevOsiEMb1S1qhN6nLMFxNlnFsLvCDSCrbPj5BecG7NpNbi2F1eRaIfShFKTbB8TJVV92
Knue7gGyljTDFLL8a3dOiFUVw/uPp8mIts5R7BeT+58E3TQ0/se927ziAsQfggnLq/E2PKaWfd/o
XmRX/ItwUqboiRlK5T6pCFgKZ2LEXj8M1xTzXziIpwJxr2cyaejBs+MdZSNCmjsXPAuRd7PHwAna
3Y8l35Gr2ow4Gz9HsrIsTHhApY/o4I5UV0HnvABcxM0IMzYHDQzlGAuQ4RvGVGF9OarVQAe71JWY
DSHgLVJyH47kJbywsmv7oNhxKkREHeUAnqyyQBenvugYTbN2cfDPkJDlNPDn8gfd9zyDPaIh0Ose
HreAc8A+5rdc+X3lUN9xV+JMK4Loe/STo4gBf6qS5nCINjZwlt+gAgBnllJz+rfyR3wAhZYKiyga
76rPdJfVspBCpcihU/NiL6HfnuNxRMFXruVRZvAAQ/e5hkIbmyARVvnq1UHQa6rU++vd1FN2xnEf
HTK6IjQItbjGDPR46IUSDUv0vG4yvRbtU6yfL/4hlA/3W043CezBOJseserBZMf9WcZwpPIDmlBg
PIqmmoReLc4G/O/xZmzXJbPrJwzAcDkG9JGBTVKED4giTXcphnyec2x418xo1QbzNKYW5tWBQ6iv
pGlhWRYrm0fFQKyJszLh7tAF8KzoxdPF8hzekhHGwTTrQMRLNCd8cNx0jBk9BtcfrUjhf/FCBN/8
EpvUJ5WdzVtQ1iGBZwvMusgmA92bhfufRbdSAXesBfb/cZzcJwBaMRUlxDEN/re1p933tKxL+FVE
5/U5bdUHNJS7GzSpQ4AOAWHxrEUpbozBDQuUZT6DtgQ7wV336uZQE3JaX/T/VOn/SuaeSjNR4wAM
64UgY80w8w0qwaVBDwVzc3MAG8jJE1HsGRGZyHCjS/IEu2ijaYqwHqVD/32+UYhzglKe2g/jmYTQ
n6oM5ATUJJIH+nd0qnd3lIfGf7a6XgVYtk3Si6v6weBpykFncOgKIwQhjAmHzedYQHgKyZsDBAZy
caGxrhztm3pON90fwSuOK7cyOXjrlqUSXeVDemWXEbFHrVVMf05TMQUnBVy3+8sj7pWeNhwjAaXC
c3rUOXaTs1I/RD3gcOJeIgeTnqvNJgkVGLLGhhnc85CLY3zfvrrG126sSh84yjWFlhK5o+0KK/va
Chp3cBL5DGDUn81QMaO/lvbU6pGbljefLJuYCyeCBRa1iMx9Zr4gncHRwnXwLdBPONqXnCK8Qq0y
ciEjct56tUpG6OADn7wiW6DJ02mM2K5HVnI3cAhFJKekUcIQbUJlKwovEHcg6v5myKxfE+iPNQFM
eXW2jeRipw3oIbtISXfNwCR/ALvkbcDpvNhiEqsyF/IFsLk96vtVb3X/ES2fDLTV9d+vvBJLL1cd
zlKhgQWXvuH4eHPbeKzuNC1T7dGeSGK0/8NbvX112FmsbJppEYaZbf8aBj9k5C74cxChxtTx1Fdi
G9/Z8XlgqaGWwQrK1yhXiBsK+NcA4CrsJjSEWx1257elRJoEV+x5q25kpMyyTHIjGTLM+zF774NM
VwZmwj6SlXpz6ZJPsFKsp9Pb1yqnJh0hVWth2w6fd9x5jbDD5hXz+CWEVLQV1TRaIj3/XXLh+kn0
gKjDxmDBE58xXBJHzfnw6OOGoh5jD1hLM4cSgrKACr3ZdDriATh6ItrroZvGqDA/Ux5G3vPRN/UU
3Jpy/s8NhPwI+olTCojxcbe3vU2MivbOyhhV7EI86jvsufxYyIx1puT7arMArv0c4YixaE8xHmqS
8YtwGpoFNquAITPuOufm604fL/ctv7CF8eL6JvAgxqrUyWjUyV9z9ad0XpCqBqMdbVn9209rOLNw
G7NQB8LWmCJ0+rfvXvA2kocqLVJbN4zJ80V7qqowXADNA15/yol3Dr1ccZVds4e0fdbiXWl669oF
WVghHyf92suCzOu03qYBas7E/05czinDuYPde5of+N+MCbEZpJ5GJeSx1vq4X+eZPEzy3M//NfKh
1HfLcdqjPEQEBUYGkE8XklEN17BlKUTwiXf5LKytthd/X8CLSZYzGwYELfax7N4JYuLhWYR9kklc
2p7ltUZQorJv7uIRS6dS6SU71aHoCFK/YAQ7QC/j5e32Ahd3YtXRsE1aqJ+NqXg8Ug7gmXEGuLPN
egLAd9WltZ0xeWCwmcLnsLKfoqcvz9IwgxcT487XEBCJ94QXq/B9XoxE0/YoFOaXpXmY2ez4mQnK
dLeg3xrCKmJxjoBu2fjWB8aVzCTBzxXn25QA9pXtlTPpfiRTqCsLMwUoZEsqR0iV0fjfpECEqwsJ
js8FrMcVQcamJo65/ZkNyInfjwCfKiHc7DhfeQPKcmknKOU6DTdIO8ges5wjqPUkvMKtEkYAtGXG
NgbjfLyEr3xh8f8Wo/2xEmDKi+AhMxvyZMZVrasvxSiWZdh94qAsyLCIf6AR9wR5qpoNRmUyEdwJ
WdaIcFkirAfdAqzW8KoXac3Y7vs67+k+X9DaqQDg4mn/uYdCojVojOnDatl9IlZ4XW0L3nSH+g8a
HjpxQkW+W6jjvvHEIa8AdtUxRR9c63GSXbIltSyL5ZoSvgk6MkfOe8rWldyKYKJ4VCEC8yA+C487
e3YGBrpG04ZDs6P3igB13goEU06RlTWk/Ix3i/XX/wQG3wVQLIsr6XZPlB+qG/UvIOcNBdujhJA4
KHScB0toV+OFM07TiXrXK7DiBi1tiIq+O6TneyZnDexRue2cBGygx0CRfiZLluyXVeQoQL6RBiYZ
0spR5k3QLhyyuWLz7rTpo1ZVaJxwS+KpUkVgmOTBF808g8/pghkdR8kREKWP+Au3HwBJscpK2fq0
4MFZsn0BAszl1e7Znb53HPt3/xMPOyVY9h9QwzoJ+Omo26NsU5kHOgMGnc701HRwswG9nyGLXDwH
xb1+cKj5jqh9SRWcGBvyGo1gfA0Ll4VdTDYmWLy1aoS0V6nmQaV09EgBtp0GsMGpFGy9Dhy1BWuo
oRrIm9T4iwiX2gSWvOBQfTJv1mp43w+VaGjfk2LtWiW8zzioZiauvvk0kDLkwsi+PNNMxWz4A+z0
+z0bdCAF/0W0tw3dJZ+DLswJ6z3I15ayeHNngC+cTPVMfNsXIMM2L5hIAUVG62hVDy2uONHyJ2aG
EPMHGWiQyErkegww+1mX/QqydnT5TzMf6FjndE9FrHOWlJpepKK7JBWFsl1taOy9dYPacTZMNg14
qV/TKuD2VSt7oiEC2j2I9VAvzAKh/VRagGvKS6hYD4lssXUE+UItOK4MDj0CTe/xUk7h9p9Gu8pd
UWqR5n6o9yBelBhXhzBRBWoy6EezudtoD7hBin/DYmajc6cXHHSklXZ1wDwguUPqdqxcsoH7l1vc
r4PzdBUPghVAIs5ZE8hfl5nuVQtZncH84wWvAU4eNyefoXH7dsl4clduqX/oJKzmzB9w5ewJDKXj
2XdOgNTaPbnFKavy66ROIkANerlzqQbLRa7/RdYM8k1uUrV2QfrJCONOydtjrdwYxSELSA/wsggr
BAHSBjkLKzSIdh1YEbCmSZBCZu5MilnM4u36D/usQ3bEFS6Ab0pDFgDrYwC1NnDXcE518rxKOUA5
PVSxtCWbPExbVTHKh1Aia7iVij9Ao2ZHrHqG3Jg0PBIaBRt/O5XP3G9BhTAGn6l4w9qMXwqfpaP4
NbgLhR4y9kyuEM3fCo47Z2+tS3TKWrwwyrz61XcgNshjXEZnT1CPKLy5F6mi8VlgbguY375gOBwp
Bch5erikL0fDa+GPs5Y82V55TblmGpQErqD5qFVLZBwVfXC4m7KJpSEaHJqtmxHTKsHtKg5+v/Un
9u2FOzJm2gusUfdhGDS3d8uxh+B8hMVnA0mcpltBwavjzJJTLNdWk2dADvNkaAfs4iAdc+dLKZWS
qHCErpAio5vVmVo736kGsede2ooRO6OrF3bdZCToiCItwnZyK54DpoBXoa4xBXqkL3J+IEW0EMxl
lka5vzrmUxKbEYPGNpE2xiYptTxbj6DRZejzwszj0F59GEhyceErz+1nKnKrCUP4NZqlS7kr1eRc
+UcVfD61lluEAvzuXL5P2QO8lC0OK17bvbijQJvXNk7Ul3BzbqodaQ6yYapCzXyuaODOu657Q1Li
/ZHrPrV0cfky7xZHSuNze1HJ+DGLxQXbIlxdDgNfcQ0DnH/wbiQr8MJcyjyq6wOB2/hEJUWHK3e5
uKeCXDifO4uED0VqKX9Ycga8B/Kh/HXr2vgg2/cT1OrDLgISX9eqSzJkta28SBtIInmccIQWKaoB
67ujw1u+pgzaPCY4l0C/FpEkxwjEAZnQVnu1R08DjAcTrdEJNeqkfdsMY/Dg7oIyyopZULyNra7k
XidRRG6M8PDHbYS91uXwX2RMsZbCSItLpBNbgWOAvkpPFynMu41JUifDVL0IMaDxfe5MXt/uhNuD
81RnQkni3XtL9Mu8ih+LSK+b0KDQyfY2+/USEBExBWfzXhJqebXVI5pRCFtu8bn8YlYzU34D/94g
n5hdogbwrYFwgIa6U13TQMuVOvsfWfWehz5ke8Ekf+UeHJa2Nogpk0xXIp7UEAp2j/twpM+tJoDw
PH1aDfIhkWFGNXNvzBpNVoYTLk8fF62DV6BphCrimczh2pCiO93gKnPaZiZbBXEWsd7OU9mmsG7+
nLTugK13OIfMtjNYWKrYlJOtT0jQlEBWBGPWRja2fvWBMLkJASvEM2WmYerroqTaMCCnP36g5+o3
6nWwxbnNN5btjd5D54CtKR+LOStYUxg9aOftN7x6YbkBpJSbmRldvDnAeyiLG1XP+3/H0aW07vZD
0bbpt/np8Y8DPTnQf3Lp1cl1wyOdHE9/1xjWMpv6uz92jXwgxu9auzdCCxJ1d7uXTSR6sJBYAFDQ
jQtMtsy/GbMMCR50AOWWIHRcLEKAFrRKgQWFV8Oix9HXTrRCGheb9xyavpAOt7ohy8R5xr6J28Yf
bB3sq7Kkaq9dNmjQm+CRUmdia4fc3sjrsvPUwihSOHtAgh8URTiatHcQTg49wwuec8p9Bh16SRXr
oJjTJ3tLOtq45U4AZ36IJfaliMFVV1py0jFYGc78/VsQzwjfwPboOYMKS3gO3zKzuzvzHVnivFAz
9D0TKEB7D4Cecl5W767uKFNo1ypw+lEiOW/zixdRE8JKs2pb6IfsgJWfn4XnpHxyEUIW36K/pB5n
Xbu1CZD8OgAdsQwRJQO978vQP0c+lkxIRhXdJKoFg3zQ//3pEhOVTopcBEf8rCAWO6cyp4EFKl6E
XS92ll2rl7iDeQMFqJwDh95KlZ8Rn1sX9NHZ+xFOhzc8T6MeKVrot8KzUTbWPs6yfqLXlLUihxsy
YCjo83O3uxnD+TNWAU7q5Cth9Eyv+t4D2M0RNJoDpVNV0HSpaKOyAl4Ehb3fbg9qWuygPk2xoUpe
bxkxLc+xRwiff78vObXDAlBo4o5aMtcRi2yc6Nf87ji5OCTSM5rXCg+csNXR9UjDx2XQd+EkTAV/
56vW+EKeh2RJFiXokjCZmlyEZae5p73+tRsa5+8/frawdOO3AfotfPp6q5GPQemYYDtphLDX/sEt
C84ZHE70HkAE3SMitOQ85qnbw14SRzboQoXJa+K1/q8By3JbQ4ZJ6nIBVntP+Z+Hb4QhcK+MSK4w
wH3rIbUrYiyfxQrv467xyKAuE2jxQ/PKs21631gmGrnqjV8nrOTBAs7Q1+zs1lj+BV1Tx92KJgCM
FE4w/Ld8p+EeURtrPatEAwW/oKBGellnkbgtOAP2THBG9lha2US3sp0/EjSeoJ+z5E0C7c+9H18p
Qw/ZdgaX3+Ngab/n+ja6q3o6fJPtLvy1Jkq5S8fScsbYQgh8sGJzGmO93EljIJXwj/DlB2jLA8o8
dNi0VawhEOe7g96y7hNOqUWy2mfX44F5XhXoJJDreEN0m5QAYXnw65TH9zhMqd7pGIiPJ1VCKe2n
3AF2R67xGufUT/W6U2aXzSovBAzgbtGcpjNhCa1aXr3nCgQcrjTqCwUi8z/zS1dNSMm60F73uFnp
s7PjGRoo6tcu5R0xvQaoGkMNHUm5JX6JTFPUL8esuU6pzpF7e2PgZ5Up/d9ZhAK/pv/8/MK6Txws
JMxu6ZArRXFbwGcIIbYdteTXMZFkC0u3+vSntQvVuczdEFG9vMk/PqxX8u7q7fojuR9a1OTPgdYv
fPqSR04Rkul4l5ge+xQYSp8HOrWl0qSk+PPZ5M1yc23MgDgfJIwEfpa3CsUEXKCLh4sn6qAQcWc/
B72pfv3touTqo3W6/V8Yh08AmtSbOG0weVYUICE4pweTy1XOi+otqlNuucu+BpZSsEvrug9NlTYV
k/Kdzv4YoLWDZgwLWXiZiy1ZYCzU24XHC/akRI3IpRhPFLs2AAII9LB9otzzsXYfohJtjRK3YTJW
qkm2BHtekZOuimC5G37XNn1YCBK3LVZF04itwq7e43MmFLSBHbinaiqBm76F0GCDCE+nlslKX+8Z
uwUFid/0CHdnOWpe0vdQu5m42RdMsuQJDtq+Gq/Z2zCg+8QC4PCFYwEVnREcdEGPJNXRC9dVmCPa
ustQJPKOgdz5tGlEUhAU4xk0wv6NRBey2xMrDJxbNEm5hgEKfMEim04xpLNbszze40SA4t0ySJ89
b2bLgvMjGCkxZbpD/u9EcPIYL24ZJ2d0msq4BtDX9OlJl6EDUl2ocy4Fl8vZZertVGcGTw9bHkQK
VkBrTYI17NFSVI2CsgSreash4OK3cI0sr8ZUcJRFN8lzGxTVc0H6DzyNU+S+qogeDNk4aHsJTj8e
mHTfiu7U6EmnBamjWZrOWZiUZh1lSYQ9Xc298SHQvCqGFjqMJVa+Z2m0J5uTHq0wXRfrPIQ6YOVp
sGFmBi/DQOoeAVOImopdWmYolawxl+Mlg+88jAEyN49zIgoJp57eUFn7gxWuPaFOjsoItq24KwJz
c7zDwbi/UUTVS1muD65PePUnsM2iuqLBFg1UXjg0UsddHRJSez5SUZQS4Up1+jKQMuv3DrD0YZKQ
XPVHL9aQTgIKwTrHSf2sDvlM9yG2/O8ToudBzIzR3Q3cpryYcHw1oTLYNk2CRPYWbLqgwVqIm6m7
CJnkPIgbyRFVncGB24ohbUmglJFZwvrO6j0+2cENVNZ80+Rb+um9CnIDsMnF/kDRO4myhCatpWbN
X04kza3nn/NEvbZjLNBSXynurRQKjTmF1IcXH6lJjhsugsBw2jqskZYk1yi7l5ceiZiqie76n8FO
XOQ5tlbZLGy/58Nottw4vmJaLZ+u/P4KeL1yncFHqSQ61PT+omnjQvyOfbzjc3pOoeeFzpkkp2xR
DyZVxuQSnzQVJJRjUE6jVfsB4ETWaiv+7jlKUfD9AnhloSqDTK+q97d0FJ2fKMxCdBvwZ/ruyXNs
Khq2lfZv43jNi3Oq03E4GYKCexO3ky5JGEhYdE1jFqLtmT4x2l6pmR0guaNJPH/+tLLvBECQdvk1
mbRt/P+iRGmk8F/8bQj1t3KCSvH9JI50z7MhpSaQDjI5+xBpiGaSZi4Gk48CnP5lkgz3QZWtUAR9
KVtNC6+XVhqN+ArCtcQt0sEDJCFXv4nOwQZ0WCjHqI3ul0JNjw7QAH1Y7BsbQkqXrlcHWNAb99Mw
/NoNjkMKycUFdh1G9ByBMkVAndu04/zMNCTnm0e4bjKthfKkyZwQ7JMTet6cU262LS33p8j9Srmt
86l6sDbJVLl55ESzsk2utWvhRD67D7m/Zlt9mNfmia+YF78zl58PzcRHX6pjbd2oB28BAdv61OBW
uHnmB1WSS5l+CUoQFsM87mxdFKXkwuKSRNNpmMA772qwC3NPU5RpHw==
`pragma protect end_protected
