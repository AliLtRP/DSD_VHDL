// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:57 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
QGHaK4Odeb7eMo0uWiKCkQ5I4Ue3TBl7WF2n19KfpT7muSjBsSWWSvu8PwO+oTQi
cO76DqycsNdtybf3Uvr8aRehUQofc6sQe2Hdr4ZT/qmYKVGBcp2tBqVLLRcctO8r
RvGS9GMouziMq+fiAM3Zuc67kTF84ZfMF1CbvaTx0fU=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 7504)
nhR64ff74HpBM0LGykJKG0Yt8DE1ocjb9OvccxPK+SJeISDCNSreqYPFH0bF+zRG
hzbdgZFka1Y6SBYj1MT9EtiZoWaMI5D3Sa/g89VtYtBvsOZa7s17eoYYeFP28L42
vEqlm7O0A66cCMQ13SrzngRmj9FI6VB/LCfEmiBOhcINpesxSEzs0IbL1p4JDMXq
sHO5y/3L+G9sNd6/5t+YlhajxwKdIHyDTpZnouCOdyTQ5idt3Gi/sGsYL+7wXm6l
xqYqyrCwOBvmL/awODv3V7a+As7+bmcbafW8+XVQcZX2oPcdZBd/bc9tAVfnhwfs
iMIkYu0/eJ4WiydHAeEclvTcch0y6q4+ivQx2HPi8JkyO543wfL5iTwaU2Ig9la6
703LwtTdFNg/3NilPut3NmhiWEA6SCUtkQLgcDMkP2U/RSMNFyv+tVfEqOYcQv9V
l+28XJvobnbegru43ll0KEPbgWgD41Up7eWP8wYWcirsQzlAaX+omvnjgztztaUY
55ZrgKzeRjrNvhbwVFB4dJKUhhxsgdT7mOZqs2nduYlRLgXrr55f7QRCPpX3D7uE
1qpKCuMCohWNj1GKzVFwmgXJ1UgjKlM1m8+knHlTxN6ba7O9kNPESRJWlb53Z1X9
6wybC7wKnevk9gjeVyDLJnUCowo/zxqueLi6CT4lrLKgR1ddNKlzttrnS7wvfHJg
2FR3Q2cREWGFtSGx8Qp0oQVvhAATwjJT6R81wTW1CxNHMYmCoMHBHANfw9za5u4U
gO2+o6GqjAnsnrDyJVYRFTnw5YABWWoq9KDvqC0f+bpxQuyVXe2Aosw1scWCSgKT
QV07ELiHAEcBait1VH5lvNcvihPmu9CHuMgUHS+WyO0AGYfYN334MWb36jQhl8J9
UKcDBZES0A/rWwDvBslNoEbiOu6ebrNJPZoQyB7MCGfoJelzy5dHmcbB++MXKQk8
wa7qjLQE+oAScnTkhhH7smKXQQujCqLaGqJWCVPWp7/CFjO/9VcaRHCC0zTDjCCQ
6HmSykDgo+aN8kzGGWPLc7dMYiK5jHV5MtWLbg4aerb5Sa0N7+cF34zszf7Ni9W5
TrzUoIxi5LLR8yrc+yl971EGAnzYpGKMaBrGNpaUa8P2hb7CjI4vsxeAeW5klEyk
2sfW17XZU3dIusYFiYOOQOq7U9uYvqJbE+Bdzou74slvvWl+fh3K9yek4iicvU37
+ZPTc42kma2EmhfMdjO1qalfVFQ9vqixls33Ta/M9m4ngUqhJb/Wt1D/WFS8uauW
WLQOoBMPfiawKo0kfBSb/PRkXM16n4BJ7T21pADXbVBIkQEdGN51tqsR+igr4vUG
Tsuw/vJAEk2JI3pOK7M2TB/EUmuI89IajzhTVLzpE9LjBOZiPMAZXKGvjnC3ciT3
+97XOiAX0a5cFywUgyvYDO44NE41Iie6LwiDu4st/4h91YNDEUjxYcICDw1SzP6y
ogsymb67jz8836Y2DOi4jy3i34seXSpNkhxCT7JZYSKXhrhOhXcxnoH14G0RprDl
LcoPUWJ9I2tMM05LKvNw4yGuhKL+JhEc9gwR2mIGx2ZThrFPZy2KooJy5rOxhbiy
WRVOEElTSpoxCwgrUwp7eM8DGFrMezUnbj10dbywXQmu14ZYy+dfB4dpsF747CdU
6DTZHw1OF6NIsoWnxzdeG9y0EX+iefsdqj14qtYsgOKlWjiUxCdxcDK+9HRw39dz
Otb36o7cbkAeunFE1uz4k46VMVMYQVS/aCuChHZkYZKbIt1r5S1xfrAcTXqX558A
mrJiBOW0tcx3fOzsSeSXxM1K6hHT9ylzCMBNE3Qj4BH2TcZZ2h7qRHysqDPqUscK
VR0M0dZ6/CJt5jam8Cy0VDlRZ7+OtaqjeKpJCm4l6LLcoGk44ZGRGCAqgQqqW5pY
nS7BGArtO4NcnRlVbAl1RDPEj0T7q8r/LueyNUBRfOKoo8zIwvl/yv5KdsOHqFrR
WUWvw5R9bMci8nq3+Xba6IeNk9UI/fvsnH37tyVXyy1PdcLbIFMo7tzMW0zYm9Jz
lcza37cOb6XT2I09Nfc/Ld4IQcxDUXzQGidXjblI1dMuG3WCruIOdl0OrgBVtwpc
08e6dB2qu/NGTfJYqBYB2UhAuCpLv9wW+uvBHmrxHP+nsIe+z2YhUb++q6Wa8KeO
2n91gV31lEwddpMupKWlwwZAJADUJ6ASGwwHlskPoxw98X+V/BPQBpaURhTo4fwG
u7e0/zRIytuGG+61/Un7tUry0j6NbiIbj9Hm1pdgTIRcqhsfhe12w3PIvNmkRLLz
pkvNKtLZ2tcK5DjpumCop8Wv1w4eQ9BcMSmdLPcZLS8HoKD4lOY6viL3vdG11TeF
8R5K85CyIAw78uksVY6tNzKUhNdFaEfcUzxDamV3roPL7v2yVq3RW1AdcOXrc6wO
ACpJRVnLL/cPQGLwLwGk1V6yZXHJn4wNLLA7qXPuze484U7UkKFd48dKnwjnRlHq
UgAeYiRVn6wk2UNqNHjt7wa3qY+M3Xqu5E26gRMdjzLK0EZAxCcGlOyD6NJdCRwu
PbZ6Gx/oZrwAlLFdXn2A/XbswduGPsuo27BvpiSbgLLd5g8Ytebg/dO8KBXAXrE6
TGC8nC2UmvH09h119oudRXhbrcAEG4gTlheGGiw2B9bs03XWUD/aXzzQIHKkDDUq
oSuCxZ/ZGFOelnjQvhD2qgNqISLndpSKy0jPnmPFIu00LDg9ph7vsj01Z/tnZh2Q
9Kl1ddv4N6IO0nXx2lZz6OStlOzqRac6ExNQi0PvoR4lIQfHO53HB8TPEJGbBzjI
gwl5r6jqJHlkafYf13ygrAdisAcy+3F2UNxwjGyEt4Z0olz6gu6MKZwczUWuPSoG
smWJNzagcTNxyD67WQNreL59gZ13tEWmPN79V7EX6ywv09Or+FICBTlXN4v9LBFL
xNo76W6oUv0q0F62VKeBZ6LUKPPZXAFsVnj7N+6LMXNNSKDYx6UiG7mnLm0vTz0y
fsCH94YKHimKNoq52cf/AtqQmks5pzGaTLBNBI2NpVQ07rR7UmH+jZpvqdhjBHt4
S0E7fXQlnr6DgMEPNfIRYwVk5e6ADtDzy9pzEX+/7nQmSk6vn7BSGn1Bm5S0nbQM
mJNzdt42UIroJ8xtXcs0kpBEMwjyuuBDj0Lq7PD2W3yallW5WGikKKpm0+GVX6mr
TQgmCf2jQJB/uKBmGxSWhbT2ojYsPogCiypdJmACR1x/6lw/W69iBBc12YuPkd8r
a/qRMSz5SzXanFP1vuqqBQYum2T/2Vyg6fgAwvT9BHWVdM3NA7tH0e8gsSGh7KHF
c6MEsN1w+qqjD/GS4x7VSOumIRZ0RVE0Ym1ZLP/5rrSIYfAkCCDt40j/xpVV4byF
xukH0H+nYvV6SD2QY+0lPgFv67K1Euk6xnBHAzJ3h6sAxF3M2yPpuqbDFfWvOow7
uy9MX0LlSEXNC5kZW+zRjXRBLN5Y30ggB4/u7VOB+E5ZX0PUsdStna3ZkJK2IW0n
F4Dq8nCmWApDEFbRRrmQwNFUzJ7j1vSBKdk+EVGrJ4zTnVv5Ll9c19IlybxgVVS7
6wufm8VPxX2ikwcngvm1GMzyfGIvczZvXtdqIj7924880IvLzZ4AHasZJCUyvTcD
knwljMBFhdp2gqQfwBIc7a6fbG6oCmXujlmiuX6bqOHS+SxF3ZUeUcItVKU/7g6O
MY66P4gARFV95RNdOVpxuybejMn5Bpa+WEQAy17kgJpodccaBJXECKHq5rm8fU+P
0O3Ed0NZ7j/Jls+o02+XdayVOw9Zmr9nid6if+/pEqI9VVp/W24WtfULhVzg/aLw
51i2UWDxPe8hkuA2JnBC2Yxg8UoeN/cCjGGOBvR80hxhQoHLsqqlE1pVSiOoA1ik
sTeWN6nGCNU8wvkwbeLjzscRUZ/jv5dSK3uilY/lErx1t1rh9XW5/TyPJs5MMV4k
59EwXwp2Ikd/pTvz98hGgUy3uqktczC3Vseh0aBEBb7WPSDLm3xKfZaHvAdf4iWF
33Yr0z6BEYZ3UedyQ0blTJdBbYmV20WymtQHqKr6KOrfGfLyqPbce3xWHUb2u69P
aO2sWMq/5Snl8ip72cDI8U42d4z5B0eytg4B4XkAJvf+Kyxy5/XQvFhJDRK+y6GQ
fB7EgYLnntcM64pY7Dzgryx4ghZ7/Rf3c/fqvVxHQQd9zTymYeczVaSKYmOp7sBP
+Bmf6zdajGppHGpRMm9cTHOS9b2eo+QTtH4pnhbLp60xu88o+u1d6H+pbIh/UZUi
Pq36m7qOW5amTfkjl+Zjgnk/380wdxD7Seu/c9FBNffl59vmVnxldBQJXNuVaBLN
xDvh25Y41sJolcgckpV4bDoFxvKQNxiFtrG+KnzJQBZb5r80HFQKXUn3uNxzjGUX
hSKO5fGytfgz2T2NjZzzqtifrMaHc3zWz0ZNRRf9OSZek5K/vJxmy4RjmaLZchd5
LAYdfvYM+t6/rfCpU+E1cccWUzfO3ZuidmpBJOX7dLsReT7VIRg98msEtTxt2c7k
DIZJg3HGqDmUCPnIxM/onQyYl2iqcHX0j29MvbdvP31U7OPKEQ9TASpi/iVCiled
69TXUKtksyXCJcjEpwZhmD9xW8d0dtAvmOAk3kNafV3fGD372DcSYm3SL17LMykR
rzVd0Rys+TW8f2cjCHORRABvGyCeFHd8323ypCKM9/UwgVqGel6vCmrYPUPcAD15
BbM6nK7/577Vt2j8ZhzS9sbdf8J3vBAV1uBu4NHE17IIWC4TEPJvQj5786KGebUN
TrBFVpI3HUw8Y/7ZBLwEjxcHBw8+uJxRJUsmVyRsSgD1FQ32iwAcL5vnSH1AIoXY
18rXWrP2ODZp7uvQRv/qsyBFx4kaoUUI1Ho1jHk9tMT0WLZ0I7+AiUXontHq1bEp
4JYOoZb1x5M5TMfifSCqJTvX9UlifFlOenXMNKv2GEao/LSV/KIspRzVIeRC2bxf
czAHrSOkN121T6ggmdWQEyPrygEYzFzSL2hHEqK8pZv+24LXA7nY4tGUu5WQd9BE
B8cYiEUvUnYOAdXJ9Y6Kn1Q8XNi69gf9g0QMEguCdQGJOnoWOoVxY1XTUH9Dg4qp
MTwPn2ZolRrkDp6UetQtx6rXuztl/4K/NTrBDQkEYHcQbZK03/OZ7S6OIu4CqfTp
mjV4phZ3vaCXuAvF2WwmLN0smRFkAHoP06FVyCbm3bWtckMUbLh96InKsnNd78VG
MOdFMQ58/jG3OiZpCNMd1cZ9hqg6kY+sbNozfitBXeACanbSio0P9455NI06AkDo
222eaTfhS15LEE9oUX+SIQorld0WbuTj0cm4S5c6d9gCkkw9JCTFepG9oQvRlaLc
SdypdLe3JIRvGRZmldPLHF2r+kWm/uEjGRB5KjcCe9+HVbwxnQvxxR/BGLXkfR9d
r6q1ZyBLwri8oLIKk8a+oYaVCxn+mlUE2eGtrvsyO7p0m2fyf8DspniKNuMxo/nD
Erkpl66mvfvKik3HmqgfuXxkUNIuR7o5r/Z8N/9ormzolcPenbCJ6rz/Mlos0Y3Q
yNhik4bd2vkE5Qpjnks6Uym8ypTaDOpr2l9ZbC+pVOcmVtPt7wWCZKVgRmNURtnN
Sv1sL888AxdDmYF8RTPwlldsHVxXjG2tpW/5ro4Jw5yuYYIchCQu0Z0B+Kh68a7L
OliaY4iWSCvZOsi9ROAbK/oh2iFQWFusISDP8lZmTTuKVrxqylERqodAPrw8SE4n
9SMn0q8BHeoFUwp2GtC0FEt15o73BgaqxgwEF/ITN/y60DSMIF2ZZGpSoag9KbVm
Nvi9iX2DqbNvt99lLAGL2c0ysnLLCvawiyXngSVzTnVzGfRzuvSL8Uf6zKzT/D6v
I/x5UBJbANdnubxjHmdD8AdKuAr9eF7za2e48h+PlxlkYPYs8Badx1UKXuuQpOHJ
c80ja0Gx3VWNhe8JXLz9PyFN/G5ZUXjdbd8pv6bHbEP8zVlyyUk+Kfp/B6qnHFal
NjROjauSu4iRUh85moOzu6oN1nSWs0t122ozLiTL7TXf0nzFFE+ClPKgPJVa1GEJ
7REJablhOLfL5nMW/vMH5gCOrzk03L1+IxbpuRz4IQJhpoaIjjkFDP0WTEMPiXzQ
is+TRG1JkM0t88mQncxwmtRH2wQYYtZR3kyaUwLXSx9uquZ84Da5G3Hc6jcSBaGb
TPJ0s0ZoQNt3r9QvsfaKNE1Ldud0WI0YfOIhLTbUCBnKdL33ti6703E7weyS+WES
8p55eJfdFAzRlCsyxE88xG2HZtzxrXhBCrv3g6I95jiyh4yy4fVhWwC3dH38T2JK
0wC0K5n/hSq1zjDVAMrgkhFBZipvs0BqOFJJJYV6/p3vi+PZXqkLYDJJTPW69HYI
T/JlsKz7VC88ITuZQWl3XALNDUU0KSGaJtsBIMOJyOw9NCgzhpiPW9S0aXWbWWIY
Ez8XkLqqVH8xGhn7/F6ahZQcDusThKPBc49iX5MgZzbaKwNfMxiogXnkIWRIT1w+
3vdo80QFJoCIHDL067GPm6/EnJ5PX6NlJAvm9DJV5YGigG47IrM/hpLYmtbFL8sj
tyRCrhIrmEEXcYXzkeRfVTVRGLYTw4QuHq6JMIav1XTeL91ts8btzxQFJ/BCnUEI
AWRp1dzCLE0t06MzTFjM+JwuIUK1xDgs/814PnhtU2n1Pj3Ifl+8s3M7YRiaS0Kc
ZeMTpBcBJTBQRT+PiR6f5lHwrEdK7MsW7uhJ419gWtHMtkJE/Mq2++Sb0wEVRkiy
/mJcG4ZgYnOqKO3VgYUg4E/ll5yu6AD5V+dc5wSvvcIglPqRTDBSIsmvy/6+SoLi
nbQAO6GJRRCrbxGcHyIXLpi6SU2EH3zyPgaYdKpGrHU+SKhLkq3QtzX9pqWGs07F
jXcr4swuVpBX23k3Dnm6E4q4RjUIk+kuzn0lKLN2xQPSLbnoG1kR8x03vHsiZg6r
6ZS8c2WO82+GvDDpF8G4RhhLz2Tx4VnFNGGIHYqbEeB2TgRo1xeHKZJlRbp5tpAi
BIAFaWIrI4eQhZ/3sB2S+D6Y64WIjS5WKF2/84/7uPy4G6vzWWdwGGlp+eqfdUsk
d6v5U5E8LQ31Xs3qQdPqZAAHr2zDN02IUukfEVuRh5+15mGMMcyoGJv401QIwB4+
pR5uXCYwAw38QpvuhPNC6ETapTAvcCI3UdXNOuaJUs2D8MuaAoPLilio062jdrVa
GCLSxjbnABeez9hIXMPGOTvLNbm0ofLiggwLZOEZh9CmJ8487QVdeN0+1/iuSi3u
1fhYoSnHY7cj3U93zA7HLty2cJhvWNsLC7geUW7RwnL23+Ri+wOb33G975xvBSaB
8YqwLGY9wwG60xwwt6QNdsZ04WP5/oOJH3pOfqBp0yjKs9V2qCY5/RFwvAgFbE1U
hUWbeF48yo6NiXxGquXvVfis8laLQ5NRSQVsODsjLEVKxABvjQqzeaJ92zK3kV9s
OhQvGjIfE05bZl0iif2BZj85jRIVwsBJYoMrlg1TnBfhcJjYM+901xMeGG6zE1Wf
kuHGMQyPxbp9xbJcb2yOxF2vJEVvht4HTCbHu0aj6beMqEXWSPbT04rh023BaN2x
0KHrDUDd3rDtOeloDEaxq+ublEEvT8AuQ18bxtDRIQ4P/gjF8VmIDA1MpGVZp7B7
dbVaNP8TvN1ot+H06OcnkQMIP2bPuyNApAj7MlkahiYrynxknVKFqi4ZqY1B/Bfs
DQzK/TxuG/eCNgceIr+6XR7nY0u1P/chJlEy5zYom8agE2378xHNNg0L4n53DzAl
+9UZ1PnMSjaAEXzhASMQIitSpEuygPd0bo041KQfrnKDBR81mBePW9VKd6pT1jE1
19jV+XzoLwEzFddeKVB5NwCv0seZ+nWyKe309f4dhPsTlQrl8CZC7IwsqS0N/Tff
n8fZBLE8j/+GIlc/F2qIkPrQOwiwNBgtOkqe+FxN96g2dJBOmsILKCycYrse5Wip
hHpBfejIIta1yNZ8LLFglfNxA9y8Tkepk+RyhO6E1KLMirwVLaOHH5Lcvdw8ONjk
e853z0/7xPl2nGnmtIPfcThJW1ulAjQJz13m5CpUyoCdfJ8/PiUe6L2a7cl38kJF
HVKfIx5/9eDSzA5DfX4Jk03iC+4903/FihVhI9ONknDizstaXlaWPSko54UOQr0b
xQsWCMPHgLciEvJFT67N6nrI02vNb+i/s74aGeCqfaO/JenHzN3dUxIeg6EikaZK
WybW+Wtifd5e3Eq/d0EvYW60Hup9xsxAX/8IppuwL7qDK0zAMiVspV2/ElSVH2u+
fBdQwNXRhH6tMBQelAVQAvZc4puc8x/Q5yX7bOkmZBRN/UMHvwm56HJgCNFpbikK
tT5fVRzhPaNOftY3Kei5D2NILLJXLYUeD9WMc0dtZ0QGLVmHXHYjQ4ejCv9dkkIJ
vvZHWPFvNWdmJ2/4PR3+XPtnkvMVzs6Vg5e6lf5HTNuQvQwbTBnaAwUhcLU6vdMV
4Sg9QwzlCkSoMwJ14AUIOX89r0zofYvjLfwepmLwv3N5gSAlzzL7kUCw+mulBfWo
AmRX7ZYbXED8jinfmGr5oCGGQ0bbaDj22lELwIT51LWon8bkJWhE5ErQgowA329g
ELaTF2Va2WxMbyggVRPw5S87n1PZeVccpXbEOf/qYmrC+lQjrfZ3wXgK4SJbb/Xv
wgnK1p7ml3HCU12SQvPC0AQV5G9o94AAldOjIxebNf9zj9or9nIV/zthsMiRqaBC
cBhW7RKUM4TSTbtqjRUJvJ1/xsipwDhjrmXhhtkEPmuPTCPsViXNJsGzlLZMSi4m
bBwsBcU1/L7gk5iIkbe/WMbP9aK8lYb6ZpQF/wF4r6wNpLwnb/Vfa3KVOZ44hSs1
qHA+hP37oAtULZR55xvtaxPOW+PmQsP3MZQqkKjz6Aga6jI1rPLPZBuP3vduRnDa
FDqbPH2PU68OboWctzz4rsf+clJ3vvAfBt6m7TPMcAvKi8iah6SrLqITka6cgIcE
HpvePpJTZswSeM4g/FwUVnkLvg/nUET8/YLYADZ+0kEDhQd5xsWSJzXYuX92VfuU
zZMk8GTSocuBlDuAlywRzbvosJrrY/jih6ASiU4g3RpSX6oVVU4V+UoAO+0OwEFb
tYCiSLJ2STdc48VxF88m1CkUJXwHpi/LOj5X32AvUOQ4eQlkTxSlc0WWoZ7RDDnu
XyXEqQVCPxAkQW6B6ZpFKlubFWP0w+LSbxulf8B8/M1qaFCzaHatFgj2aDexlWgO
Rhvs0gkUK1QcDrc/fOiO7Y6KRLRaVC3WrSOdLo4VMRVXzf1LT879YpMZFJffMXOZ
ITkg2cJ7iPi4e1DII8pufiNwMIqgjZ0VBau0a8LQpzFucNNHWyqI3aJV18Uu68p/
oD4YK/HPcpOjJkNNeJw6F9pOGxoNekDDOZr/gjLD+yNWbDuQOvt9JS7kyyav/N8P
/pjeSnJO6u55V6mQijiw+aGNY6B1F8aES9q3jJC7NRaG4e9/uDSXBbZ5m7xSBqb8
/vwrjndXiLEMr9VMx59IlFmtetU9jgN52u867hVCEwW3TyqMYttycnZvklnyDJEP
j8Y92hljAbfurMtAAc3lE/q+zcYfdWuAwszt+T8HxPA1GcQO1VowRQe6XTYiYMGw
260xTRmG/unAEWppiRl2nDu9DZSVJ7Xk7gKjwjk/pcgHqoY6NtD+myuPmSvcbB5X
afDQF3ILHDoE1CRjtHuEsCDAAtTpJjQvJ2PcaC5VJnSTuyDY4/Qgt1jdL+YjKZll
66O+POfm6qhPqMezg7o8GV+Y35iWeHqBh/ZamblPA1nTKc8/lNCCiZxTm4Rl7MHA
Ku82hqGiFvPy3cJTsew2dUX7PwaYUzqPwxyOjRtuzLoq/+USkdKZYRTyHqW4cf5Q
ATqq3uhathM2CKEjOpNZvz4vCq/3KqJpxhTiJ9V3EFzgvypOmB6WVpj37ZdGwhGy
7Q0FyIpp5C3guJhcZi4AUg==
`pragma protect end_protected
