// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
gPhM42NVhEVTQ4NcpFef3MouRVKM0lfHn+1//9UY0xKl7rLDJGbkHF6uwSR1+JjPXkJjyCckSyPM
oTLoMOCZeWoynt0xDmtBBSbETWECmyn8yHtLyx4EDx0REog8KthHHftYqeC9ouQiILBCHyGI/0EO
7Orve0h2j1dHujnVHyeHkOcz4muKQsz7xhFThufNwH81DcWjtrHJyNxFJ2kq+WGEWzY1qQIxkJnR
NOiJ9UOC223S3gDTf6xp3G6dzbN2SNkt7D4D8NmkUnxJBf7ur488U4hrdlUbzqP7bufukQ/WvBZr
O/LDYtR3eKoTwmd/cNefdEfXtYECd3jwif/Glg==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
yg4Ck/N0KCATaYyManzECm/cg6bLDtkSNrqaBT8cBCQKDvBKQ+57gRGW2Ht86b9dPpM3HpgPanZH
/G9zIUW2iYlrYaYE5jBoZ+YMhhdSMRHJQOl8OKwnceS18keELa1hEzSkrOa90D+G/uw2rTYHyxpD
0XCzD5vjltkeE/okIm+OsPrtcg0RJyomyQZMffJMGM8gHkjRFCUAgivAtvhQZE9k870puJUOyvqC
tlDh4r86jEPTtb1EpAkAF+cT6n1zE6+0zCTStC6lW7FVMJYlZUIUDJC+E5k9D9stYTW/J6Sl9vn0
NXMuNL4U38KTAuRAgz0JTmlChv6nHu2zfxi1boVVCiD87VyGhtlBzqjo+cbsqpssjBPP5/4voPWK
OHD2gOaONnrJ+C+VcIZItw/NXamRdhL2D5IAAGz1pqBECJuVuQ0KMvEHPlB5PyRiPV/cmUb/aNmK
QQqvA9Lv7IgqQh50Uqjkb1Dginvtm8OXXrIXuP7d16yh//apNc4Ub8WwSE0fKMne/9gSm1M9JxVN
Ruim99fVK1RcP6q0UmxG0662fbc372BG45aKjPDMUP+e63Rnf/uUT7SEi14+uxOJI1fLipwqdiZg
HBGbhjjs2ebYOQvoeIpKaiqxBMShAkYA5jZAA92BSFpgkdyV6i0aANhUHl8BUVJOF1eXhm8f6SNV
5kighTnC9zKGPhFsTwMfrFPlrAiDZhwa1/NMhYkAhWiBmlPEyPd1QKW5sWS4uzkmjobpHxzy1+0z
BaCg1rDwsZ3fc2rBfcns/gdotqpg8QuWqfOKxvkH9IDlm5MWtbUnAGOpZtLDz2M8dIbeWIqKO8s0
GlvAkMyttbsMH55iMq46Qw7tP5DNfFBKGk6dY/uQFxwiED5k17ybtmuUQDeH9I1fMbcfqlt8OBbQ
WQHMICdOHJLb9Mg3e30oCNK1rw8YjuUv/pPRfGHRjMq3NRDt0vQGB13lzqUUO7znlLrXDvybLuu7
VGA3xzBdqW05t1k7mvLI4DudOOOR55Jv4m7xwVq8HeAj+qo5VHjJIPGcOqoDnlvkXP6ln/SL03XZ
UFDUiM/PUgsKxnI1GHihhQ9lYTbDPmMx071CpMX4R8d7ohaRvZpTEDsu1NzI6ODH43Lh8/WeVi7P
XZummt/EMhe/quhRdrlf/qMVqwUlSfkU0xlSWFcKTzQDp8n6VwDcD4e8xh/I94xZNmFTYO24oTrh
lvtRadGuREaALrfyrglFxlNIbpsvveFjR1dyF9USes7KQbWY+PSALh5TrkXLbkQF6BrXcK6IWTp9
+sLSSwPd24ioyjLaIP0Hj9KWXCH46qmS5uomtagW8n/bbYFbNNjQPFq793HLz44ajTVDRM70I+dW
F6pRBUJfzINpMGvCGBnD+yjsqWXaTK72aQqIiKytRyW5lpicrExFjRRn01BACk32I5eyZoeMk39k
KU3wTECQnzJqOMaLAb4w3dV/XKMdxTuouJC7d2W+1a/vemz9zdCzXscj3b2EL+pbrPCD1rcnveR2
0XMiJUV7QMOpWBBfckUC6c4QCby/BKk50+ZkNk8JpKFkuOODCWUzei8bUA/fP4DYiuM8x+Kq9yRf
qHxLft8unM4vmmtSvrHkEBnDveI8gTYdmChj+fgSB30miF62cJ5/8jchJwg55cmzkoKXhesQ6DhT
Wj7pGxbtMo1HwlnfaREV9U9YtefLJBRDwRR2Pozkx0J1fQ2TQh18dblp0AiFQJ4i/fs/zs2LbiIQ
P69tUbn7qRTRP8dsFgBeZWaUbpFQ+4/ilTYG+bfz6uDHt+AhhBB4n4d/laebEegz3b4ZPEnoOArW
kbkcpT+R4Oi+j6n9QriPOfqwOccJAIRmsG0O8puLos2pQhiWBAEwOR84keGVZkIwK4QkMhrr+geG
Aru0GzTG547lpm3pk3V176C4Urw32qpABI3bOzPiDjqSW0ASA2qSQkR9HZpTmZVxojAUcxMwTfGG
3vAR5jCRDYLPZi8xGQxdmyuEZG7++rpPSa1m3Estx5nZw6iSxCGzJ1VUTfZSpF6CxyWN6rwLKdeb
w9jdl+Qz0ougBi7wnWzULuVEIRtiGqEkCio/VUyvqM/sQBQnTsU7/Q0l/P+tNI6cv5JzCIKzehku
hb4hmRVVgTbMoBoJRS8jMqWslDOyWmOpxyGQ7NzcvHqUrt+9vTE/YsLizbDZYXUUjwD8heneO+g/
zC/eIbC0loNs+rxkfQZfipu1VbNwXbcLCRXl4ala0mZi9Riye7zR6xe+mK+w902G1yrZzIw6viAA
qZFhavcEGHYJ0SaZCH/VyxI1FggGiNrHQ1IC4DGVQMvhkKr7EC4NfN9yOZZn4DcgbnFqibcuE579
qzM6BEo4edmMxZ6IXApOO3HkYP3BnmGMsPUV7qbfLcpRhdF1a+X6BGP3ONeUmuG0sTSy37YfQSnI
1RvtwG4M4pJ4pbkBcOL4+5Ukc/u54PEPmtRmo1+sWgfmqRWUOudRaU+52eC0yapxOJHnAxW7CUVJ
0IFuMAVzEfEv3lllVbK/p6nCRFQ7zpO0iEwAmzgAQVkKEuMSTSPa8zF6iCuS47jR93fdQwiXIeLv
Ss5Lt4sAtiuz6ZTQK6XfMoj0bNZB6fdghCdpVJSbJJvddPktcSng/ekJCnIMg2VInwKNGnwh3O3D
bNu9IdjvcJBJRNWYD3o6bpFyxUFqLB3ncbAQNaNsKr969GH25P2/k9xMcsMYrjBfDncD6xG73S8M
229BavbJz8AQqIBSnf/DkBRgSu4oI35m2B5IjmEPM097hVepk8PEDI9adnsTOW9j/lIoRVHl81cO
n/b7hJ52SMGsLcZ7AQ0x1sUlGAyuhR56y8Vho9zdabolmRntkgqFWC2blmFB0DnlzGpckL92CO0F
y0TxAkAPVP641q9sdsTmN+MkASRPgT3bVnm9IW/DoetNH91mx4NUDbVl5Br6ZrvQdp2KpZD/o2Jo
kkAVLGZgmc+HzI2yy8F4/O61TaCdEojUEhbQk4fyJLdw3mz2XVBTke2wGVeUyq5DxD4ISuTsyWUR
6tkcSeR6acY4EqnoU+4HmIG3zCkkW+tYDdES27DuAHx0v5wJxHRnq0KcHhEVT0Zr4BaCc6nDgrGh
zbhfjfdvlrFxhC4RFEq22J5pEbo49oRkCLzFv7YmCSlEiPu8V4gh8dFYob04E6jMb7f1hcZocQRp
kYjC2QPkaWld5W3YuX/f4uD0+C9GgHfEvYWrU9tnUn4slsOjMlww8U7IUiWsPnahnzGoomlcFTd/
2Prn9lEGvkVFCH8eIMpfBjo08COo/trsEbbakOqT6CnSF8EtV3bQyNZ/8niv7/qpxavl1AgBHMbY
GWTnMhnvDFoPiM7gwCley4jQ/2uPqm2wNR3gPPc5doVKhC6GFjQLV1RbS2av9pAc2uGnMfi3v0Qq
adnzpxDPVrvvgxFnhc0rWmBV+lXRGtjsK0BViXhiSqa+aA1zTs5lz+KKPybfFXduUV1OJHzc97sI
foxE+dBEbYmjgI4lao6r9Y0k26fRSt5ekb2vEPb0shbcc08hoA43qlu2nKNn9jAcljTEaIEIy/s5
NqtrRU64g2HZT7BV4R8CKFiQH8dHk7CDAOuZvVsO1yJNEAFYu8VFSHJ8t4Tq83q/ka0J28JuYGg5
3ZqE6ebSE8jCKZYUxYMXWFIiEOFoOLoHbBKaduV7MprJ3Wh6EOs7WTCbZJwb6mBs0WJ9acVJzg8l
j4Ar/Qs9LvQP13HuMlx1USNEgTwGdxAqc4CY5v6AOMaNMz92/UzQhEtAhkYEZyf6sbL90VkL9Bvp
SgtSw0Sl0Qtk9mss7fo3KSBbsCj10ZpQx4Daw3lrkzpwd0M3ZRToQ5RxUF1dMz+wceOFTnw62feK
BwYk4ncXN/GoBnTkExSHBQSysKqK7z6EQ580KN4zeKivh+dkT3UAonmjV2z8ABW6EdzlT43yYaSH
CoZP0jLrIH/TH4EHRFbPJ3whz989yPCdEayiItC2XDoQUqzDR2tIdFjTAOpKQ97kOrQuqIU/LJF1
Q/tBeNEZOpWNgXLUXGBxmolLL0IYADzlsuN4A6aqfwCyj0X9WbB+oZAAVjcSyjNsqCcQvdw99erq
uyEahzeK5Xbp9IzvKiAAVXFGAlxyQ+yNd8Wc/xcfx1gKYBsFkY3WrTCR0VXE8UupgKyzshxs7eRY
DkZIF+BDnY7Xi/VAg9uZz6X6ZfHH62t3IhNoQ2hRw3kyGIWC5o7K2oH3kFVtgR/wm1oFG3xaO3wE
zC1thc4Va4uG7NITS3I2ym600On07f7wTETdj4uACOLaQwEnt26aalQhAYfG1uts/nZKlBmxTX6D
kSdjm0VOXYfxRSyDZ0tlX1UR3+vOhARhJgmhdvgPqYCrzEuIFri/py8JkTEnInYPNQRj4c02gGh0
n9M2PJcygtG1S14NA5uERzgQrK+IEuh4ujuh4Mw363DKlAunPjpGxmlQFs4tA0iw5OJuqufIlK10
UsAxZAke3+pvbf4hG/OuFGL3zgoT+IzXBcgabk0bdsDYCMbEuCuAS7fx3+WOP3wgrd0AleKAwf7m
DB2XHx30uCreCVmY8K70+1r9aLEW0u7k/2amEQ15ZtaJKjInWRa3NhbRu+aYasFq7k88+kJklzd6
MKPqPg5JrC/AeHwNfokykAu2E9L/wp1tWV/0A9LKvjJoINX/6XA3uI2d575OXEmj/E+87RpJ/pVq
bFhqzTo1/mboClxm6kCx2h9P4etSAjuU6QkTC0qGwk9uN9+Nl8R2F5JxBT0ARCWPp9/vprR66Lqf
b/Uub9Q6HUZ1yvC+MF+dPKBqa+Z5utE8geP8lVaXOqz4zNwy8qTYRjo4PnKHdDCNZOAKGvXPuFjb
I9WZEPxEK+Yz5JmBn77oOyKNWB/YRiV05ZKfqEZy2YqVkNkoAAcovWm65BPyjPhdc9KsI3PJL8ZM
e0HDeP0w/tmnO3rWNetO98m8LngCCinOryOGhrQC4e79bSAMwmHRk/0wfFd7oGdTL4ekRFmDeKFQ
76TrV4f9Yby680e4K66hbJ3j7/haPFUCKtfVFqzhUwIrWTaxASiIgRG2MQ3Jvz94iFfi0KUAw3nw
KUkAzcNJfGUahlKD/98RxBma4WruKFwHrHLaopggio8VZbXR+e0GvPpxQ5scMG/pX8OJ3e46G08N
wBobATxIwgwJzZ5bw+HrF7BuRuBxITnXJqcDyK4cInrxCaR6aIsYUKI2NijbKxxOnJMoiOfDLyd+
pkviU1qGULWF5u+6d5anQy46uLsisnVtNH6wGo0nDqjt+8KflJ6bVF6TcMXIKe8aidGzmPp+UKSe
8T0RBtM36DpTjT5WV/TrHi33UhuAmJvYOq8Yb6TJ6V3YaXXcmFLWoymFjsUCAl7MHF/X0iZo8JFB
3W3sIzI35q7U4Xq3F/lH5zFuIzBbnRPxM8X81I/6KmF8sOScgtFIhmDYvsZbBUgeYBqvbBxFQgbO
YEW2hPEXDaEc8R9QPMVMqTM91JOqAVeaDQh5cL/TUrZhi7dcjHTHp97VZ9PU/ups8zNkIRDvqiyt
t8mRva6mY5HWrEGc0Mw1IgLaT6fb3nhf0+qU6hmo9soLThjFiNmArad0X/RO9ZPTjmtcWXK5N4Ce
WLnUB9iqmUcoRo22U5KaH01EXZ4Slc3ygMBWkYfd2YUaQHi1c0A+CYIqN0cJlFjZ+3pwnQif5ze+
xJ8+U/i60cOHdj6MbwKzRfjRrhgl4xuSA1WRaE0DN6cXxojXabIejyEC7CpoLrWeTMAeZkaXw5rn
5nID4re4xrWUP2i2xL89kvp3S64MI7AvcM0uMJMT1BTxZQbt171ChQcrlz/wU6RftxolhZM3qUJA
TAVsJoh2vrutZMFGR31suSvp/DTKCPLtp/wiG+sFHTKkIifJe7z2WUu7UK/YODI9ykB9NvTpiKbB
vJWPhP0v4nMhCc0NMUv6ewWguSkoCYXvmQbn/FJTae9T22g7sK67Zn/sW2meWyBOa26GX+A7cqCo
JIgWnXAYfEe1fn7k5goIZ9ywq5CUcH50Z8b5ntcPhZM5Rhrr4Sv6y6X+gtoXEJ0UtrQuFgtEQAPv
LimNaRz4Bl0QFykUipfznRx7TGeh1pAJRR8sHEq0+gXJJgsIybZAfQIGeTQnTvcQbKnl5wWKi8I5
9pNKN0Lh+dzzMoOarZihShjslzmGK95BVpB2V8PQldqp9U699EdR0yT0OvoJXfkttWvZknZ1oa1H
PJg+VokP2LlCGD30vfOhB26mOkeNoriWze+7FQU4bGIQwAyYCwNdpgLIa1+7m2OPq3VI46eHr6Lm
iqpECuZyysoV2k0jG+3TwBqyJMIJu3EofniwHkQ4Xdnfg2Fp2ystOV0PhPjd+AN7rDDIJoEwBQ5z
TCOUbOScQua70GJevtkIcCo5CNGshd5qacZ7st9B3LdQcGchl2ES0MIlR1XexCh4YkXaX2l1pwfD
yMm3CkNYxh6OWdib569uM3eXpKyA4a4zUS70k6Bd12yHpdGez4Hx4o1qxc+LZ8ffSQ2d7hs/3gNv
0MEXGQWi/rqpcSe9ndWGBJK832HuECrlO0Rz7itZ840+p/+xbKqeOGPkcGmIlo/O09tQRMyd2YnD
3U5Y9eyFFSQiE4uoIx99fwcsd+eSO1ihcDPAcghUXZFT+oOO+SN62+xq3OOke0rTyeLkbINBH8rX
gsjnTS0yy/frCNrK5/eGPKkuBev64F0kgRdmWv+JFEKzpHcw3so56q69lsc36q9IZd3AzLDjd0aA
+vC3rgIZmq3Z5h32+lKY3zGyBAD2ratzF4HUmnBrtSs993l2TdVSHYgq9/qmWc3O3pJJd06N/ud8
4WdK/XcEATxd3JylZigeXgZPawsrvv4c265uicP2VYU1CmPDpPKXY/SNYUNMy3BeG8tSyyftvLDS
+jpAV0BqnBBYOJm2YhyTMpQONNiiKA341cm698+JMTXUucPdi7XoSykQmbre2mB0hhufbfvn2KJW
1MIr5vW4eJNlvBFESmhB2UFUzel/niNnbuOwUXTikDsIcAEWMZh6MX0rjaUYns+xZ9kkQuM8Hjvq
E1q9vBqX8OKBJvAwttFDJ0lkFNrxwEqOj3Ka2fBIliUYLMD8ZhLTrKYCPXiVNR692dY85rd0e61K
Vhjv6wUCAIyZfJO63CmYzvFaCGe6GUz5mWVmOM0Ks0KIIjCl4ffcMiUogK/KPv68DgXuw1rCgUzQ
ZMFTVjERltNwml4sSJ6NBZKkcgDxNVcI/zlHeqVaN7T7ruPNUQeFJlETAz4S+tcYda1mAHKRkieS
Yy9cE0U26PGbDq05/6sdDvLZ9wC9VOy/0sdNKfaEIuxw2qIuA8aABwXTcDVQFXdwlRw/NlFBIg8+
oi4S7YyngZsbmAw8N3FAGuRKOiEGBCjgwaBhA/oHYQPlZeUWZEH9+4RbOHaaBNf8+7jabGP7pIpP
8nvJy54k3gxJmXjNtkTz5JRqmk8PXlmJn+4UPW9PiRox8rPBPvONLe8y4Zge8MZGNY107YpVv3Hr
2cJtsMLlDVJG0Ko27oG7tKaw4UdCfPFZslb/fDJqKhsRmYzihl99EgzfvVGB7gXx4aAcwLEFFrAD
BP3Aj59zNdxCmIsMmKUYEDYwp/6vFwHqwl6SwkfmzrqBNFY5tNb941Qvvp9AkvfrB3Zba5R1dD2J
XrbCqd+95fLIlKoi2S5mzZlqyjesRRVnCe1k874KmwWC9/eRvgg2Yt3wDFPYWC9OpQowRLg5/Qsh
hs3tU9VZU0tZN7Q+n/6anrBqyfg/ZJZHtnpgxatYMSzOk3+I771hBmz4G/ETXEgJIDVwWdx4uvrm
0dz6PwRZeI/0pBKO1uOGWeVw275qb02VJqnNtZ8u+qggzXtdTMIvweSWKSkkGBGiBTSKhFd38sOv
vTn07Owfw+bF/lCK2HRBtBu2N13iBSwMMOlVJ31q6FFtjBroyKs9pOTDps7fEe9bWd8ppqWoHF23
0Zkjbdk5Z8TyxfE03T/hlBWEB6cvApdE32BOfR+r29EyR81nMq3bKF2ykyD00iY+gOXGJUmuc4by
RDoTCp3+3KX3AlfEOQAvEFb6UswXTdPI1tjGpU6TfPGhFBeWvEsLDHo35ovozyoFojrlUyHIMM4K
7xmWCvWIaliMTb47PWvjSsBRsp865aJN9EnBN0fIHWmLXPRc/NtZErJNz0aiWQ42bdyHhJn2X/3R
meArCn5MnD/btnO8SKGIx+UDCF0ITt5ORJe2vR1ibuUnqN48Uz1Qau1x995ccBgDavrH2j/HbxOH
IC3Yo3PY2Byqoer6rIW0iGQf6OTfgBJtTiVpRSPCDB8F+YmwumwbICD41NGAi9ML7Vi2qbPOY+C5
BJkHikTphaBlrednfmcZAHuduGtJ3/CpXTYACo5KSa5tcJlQEFN7upGyJ/vu01Vuz9pl17NELwSs
rUQfz6yOPPwVjf+ShytwMRNC41IPIK3BCShGCFJo/u+90MAWzhilzuOq7EUsZ2Dge00rUFb/0NRM
dfEMY1uI2XUryMoKQWnmZXtvO55qqzB/KdrVihzBLoM04u0mErCOqvlt27Dalvy7YWH2fuUiFNGp
qDUPDbcZOmKdRlTeCCmXqjv1Z7efMrfhPlgLzdcT4j3LYoBu/LgDFiKAUcENDHDrtNdjS+Xq6oNd
z4z73MVczQNemMdtnyYTh9Xz8OAlLwZEk9LtxtGc2U2PpHd63PJSAeMO1Ic2a5l/wK59+Frz4poV
F176SmTPeQ0lJgME8vb7uPOMxSvwrp9u30yLGGXiLLUKw53fXUSeD7YIshYjvxnXGUweX2j0xo/t
p44jSN6VBp/EVpJUcKKgW5fYoD+eLbhncoW2XS34taV8x6EiM/AxPQHM9s0mrLU6ig/ChqachmU9
NzNUkFkufMhuikmkBn0DqXbGFXnHHd7j5idY8gwb2qVkvG2UMUzHsd1JQR4vie9hcaCkjIId205q
g2ORdXrA9lykJox9diu29LfZrtvvwXZP+GugIQ4zPm4w1gMySj6I8HK+Q+rTwnEab7eWNEQ2VlW9
LuDx9zl4OLbreO6clO9SSLR3d66Gb/57r9KZaWpXA3G38aZWDB/JvF/45owOQ/fzKuJVK+rW0cVI
3eCRFTGnwcHtvTE4VBrvaVoTviM8UceQUeW3gC02jiF+e70/2Kk0qcsNAcYmTKJ86LjH9pIuNAny
s6Lb4gp1GUtKvtsgLqdDtE0cRQiJYF1ctZBYzWBmuXeuGOOWa8ioeNsliQTSvTECH81xPt4IApgm
y5glNlVMtcBgebsae+koxczGTXtSoZLG5drFWsvJmVIytvfL/hvdsmHLUg8wQZzygtz238rz8zrG
X75GkBdf3DIac0LjKY0OsR4LmjWICR1loS3p1Ppravb8gNDMbLHXmDKYluCDto6AtX+/KFUWJ5hI
rnurhpAvDQV1lNTfslIEDhEZUP3bGSMStVlcQOdOfbixW7qxgpofpGBsbveFkbu7f8pAD04rRaIs
vnEBDhiaBm5G12YsK+latdX+jSJPdLjiRxXzigxsWc+J/r74IlWjtU/nCHtRyasj/6v/zay5+FxG
N5Nlqx29SX5jbCSF+Pp70Ia53zOZMtfZdZwmde3+22kWXVHZZJ+D1olqtXre7BfRhIFLOQ0XDARh
cL8kfClnh4dFRiczwgBcIhgrehmJgHvXOAejPErOdev0pEbbpi8g0fyWfxvw6Ka+V9dn41zDtvBe
sKabidRgEUKfQ6ZrW8aKdKsYf/RuROF5ony8icLReVrHhlBBARQt8NnvOStuXsoQLUHOYymSyl3/
BnN7E/CA60rvTNiPfKxBR8iDPN7rqeB6mxi4MnAwPxW10MM6uHdsfLEbyTpilBxBtBAmW2ekGcRy
NVSAENjQJmF+n4VwC6vVkZysC9DSyvBnW9/WALLJA5W5yikufnok8hmbCf53aQWSLyTWr0qlQ19p
POTFDSIsR4QPW4UyNwYJu0eZIdYyFk7e/+BHPVLdG4kq0h+9JO6uzFYFSuUolwERqgW5tg0h6VBu
chOPkUMXNYgqzEU6Lm45X+KzlskDau17QJP/Whiofxx7f14ZilHRyPMRhDRcAjT4iRLaDQjykvfu
eObF/GEha0U3N7ixLR3L/l1BKAwf2WeuB0K37JVnAtUPfJI7ArEGYPT1z8LeMojyzKoV6h4oPXcF
PhnN58SkUGS82DWe8hcbmDFvbvU3Vok2iZ2KUH7PQG6O65IR/b/278+txBuaysEwqKsQNULJeJdA
dg933Vdt4b3VNTZ6mHAceBaNdA8QdrM8tsklqByFcpZetct0bunqm/eNUypOIRIOQdfyeLjOhqK/
TWFlPQ4xuTFFn0I6MqP1w4vTG2Wd93DW63F7HlFDPXpOFKX4nAOecgSm/d8607JAKqX41RXfq9gV
UU4vkjag2x+LO3mOcAqvMH1j7IdnOMoYPA9xqw10cWhln2mFppiE5kYGWOFXPsTq62Lw0U713ujf
iSgFiSHtzN7SkqPlxtHj2zKDJU7iVbvog8re9zD/VifMi4ij2S9vX19fugeav24HAI4hj2WA5aFV
gLSiSQmtYGhe3TvxX/FIF9x0CLDxcTTxepEL6T2lpQjyQGpBxOUghVf37tM3QiBh6F70RQiL908e
AU22JutUmqSTnPnTSzzZokMf07xQavPVtY1Hs7zAO4N6eYnxGCNe5PHHIFehLCbIytWF5CxAs9zi
xpv8w81rpdcWDYWkeRo1av0MFXGXinSWDY9Y/HqY/4DAwOgXurUVCdsjlseNNQYq5Xj9pZBURS50
m9ZiCVgbsW/6Aj3Ho+Z5qCfayC/7n2m9YP+nZgT6AwI5oq6o0NYVKAUvG0EBnb/IStU82w1E8AP1
j/tAnI1yCJg/Et2M6O4DvLOM+THSPfDMjV/zu9SfW6Hr0oBmbgwmiBfshnyDYevQB19n/q5+eLse
orIHBLTXBrkfy/fm4PPPDTBgKcix0JOPgzx7lHxr4WMARYMQkJ/S3cB0Oo+JY8ucRKuomExoxX81
Bddas6TDwviZyozTmzzlgwdW0FZ05XHpDXAnsST7y5bs9GGQy/CO8q1FImfG5HHclHjfRv59mVdX
deoiJIamXTDNJTE6sJ0pcPxLKKMR6o1Y2lNdg/kQrJVT8U7bP6ehd5qbj+6ZaOpYWPkdjwSSx6WC
R8Uro10uKIBHi+h2+GYhvgmlwdu9yyE/nbUtNbmdojyBhrkBrYc78mHYAsle+XpEHwqNED0s2ude
x4ZTwoDDiM4kaBahnVrundD7z1ppQeaCRW8LxNgwb86fHtzRV10wnt1yjzmAe9/Oj0xqbi1sHcpk
Rer2ZkpvtPuOQ6aRTXM75UQQLbNRWSzip3DAXbv74xT8L/vndqyYwxq5wb1webo4A6wPIUVguRhA
8aN6jV+9mFgzrmqYCqY60VyXUctyiyG01iTrCD0iRi5Fo0j2z9UchFextNghm03s4tkge2Qzwhh0
vopbve5kgyw5z0cErLUGyCNz77XAz1WP12Ml/08PTlykJFgz12KeOKLVZF51D3NYo84JBRh5m+mL
PvzRFCBm/+lMLxf9ckqy3FIVVXbWsw7uirLrfQ7oy4ReYHhjxppyTCyUZE3+oxdq+XxgO4lXGYxl
qNuuoViwrVmWx1PeIZNzZOu2ngrsXj9zUHMpSEJ/Y+c3yrUzry3dUjg983wgHCpEXkFpui1go1Ue
mh4IIMAs4M6OtqFjTM1xEGYiPkkMAVclZ1ItV8g3zqVZH2jVw5yD3AwnAez4oHD8FtxuZ1wakeHt
3anT1xi+xobZw1nQ0NLAxHDATNWqFqBdzSzZkXkjO3eY+fUZE6+/XWmkikYzrHJEmOVL/NxzlVuh
xKqcBdWH5Ie5WVEMc3/yp9fzHsOf23bKv4fn805EKlbiibF1VI4yQAJsahdKcLfA1OSMl8ZTyEWW
qtvM97jY0s9nt3wmG6l41BXfAVh6DyvnzbHpSDPFHHr+HrLBingLn+wnW4QISmaR5Q1bOxxfYDsn
LS8984MEwL9X8hdCyvJZ0ej7HJwhD2HVxpmxS83sNttxmabOKeEXJuwWidBvEdGV2Gw23rsIUxEW
IxrGHBRX/3j3cRfcvAZjyRcSHvDSAAU+JBKSuObr7P7yLE1pkq17yH85lJSRSjkGQ3l508vBULYq
5+AoL7AJSoS/E3ppNmJJ5xahsMg0k6QTwg4J2Gnm5NZRQEuZTDXF0MpX9DZ4h/J3FBXyrUyLU6Xh
Pn6e3pXB1U/q5RUg5Tq5mGzd/ISy55jL9mjzm/jmFTzSL3/ogrLbO9BulEvO1nsHGe3mwAbecAOq
z8DGGYIishCIXsDpkr5lBhm6IOPbfAcIDr8Ks8XofBgB4VS9MDIqKLTrdgRFmOaZNwljcFzpwrII
BTgo/+nD195omQsEiDF0h2FnTG711ICg0alQvQRHVgPBQVfeyEodvs28wOeRSOg+s+cpxiTGtkvq
YPyhv02xL+jaGNUr9+qFP0GMn1aLfezYWIFBrhQxg1wt6Bc6ZvZ/1rgo0ve9xmNLtMyQzvrUYgr9
ztYIUByhUS3r3x1tXgpVZ5j4XWetEhOrzG8q6m37XfnXbb32FaDCfYN3PGZzzpddGi62zhPO/NX9
aqkjHeCkZgEINt9g8mvLx3HYlpcmrnEB025U4+Q/0XqWxQ4XyHfNkb7C1jkayAEalNMGa4zJ80Xh
0Uyio/yiHg8oljGJuw64/UEWov201BtNE52KF6NoAxFxDmNmpSXDa0Eny1VqDP94P8CCyL2+vjjU
n1sqN2LfMemU/lgeIRhtgplzJOHADudSUUKdBqccqpQV3JW+BJc/ms0zClJ9cLoiG8BXNrHspbh2
gkr8VCB2PEOV5fir53bS2zwEa2bIRbsbR3d5TJ4E/e800rveVNuRmDpIx+/02J0OfuHszn5EfMUX
lx1HGOqqHtvYtXfAgLDdH0ELJTqMjM73RLVwfyvF6agWKSzZwyBf804uKDyYQJPyMZrDfjdexpfS
+dXgwAU9CVKQrHt0mQuzkLp9k58gAn5edAm79dHPu1UpgcjpUt1+hVeNORUWqz1Jwq0Olox88nre
omh6u2rjwjVVQ/mhWDymCzbwAUu8Y6juPIPczeh5GZhBzc7juxyG9Ps3ByNFcFVc6IBFl6iLyP23
ZrkPzrMYoOPWWTCN+En8HSd7dvZwsbjKme9J81udYU7/E4ijODEEaITfDu8JbrXnqsdPJm5AwnA5
aYQT+LYBEnMcjGUOJDoZrnOzpd8EYQb60vl48SLr6/7izbNP+JtTNgBm2QDMwzUbTdrOEbswsWPR
5WevM5JyKp8MOFvNZzVPHVUS0rCC/L9T3Qo5QuZlsSh/4cZE6GYQTj3NkN4v8r6ugPq7PCO5iET7
TYeIhPczRGwOiZUU/gUWqdP2tQFUtlTcRC2X1MWGXH+u2mkEkxmOexw/pAINDEE5LmWMO7xRRqym
MpcE56LoAEx1GSr0s9cMKghNmvXVVkrebuE+KOY8JMihifUDTV15oAjfpjpLUy6uIFgFCYbLH+tT
eNd7ovL5fiyLMBlnWnBtvJRsTKSqD6dKlUC7WLWo4YMSrGfeoNsvGq+cyDAGARwGwZTQuFhyxxDh
8nhjqCnoavG0BoZe3oPkbMC7CKMbw0ZwIxltsBulOk6pFpaGs6x418SUer2UHteNZkICK6pCaiFI
8XB4cA7B+999WD8Z2EmFldyotLTLKH5x69J4d6JzhOHH2coAQIneX5wR8ZloT2rC4V5Gcje+vggN
B8gsdw9yccdOTt0/+eJvLQL64Ymlz2lWl3X0CHECQFLnY3jhWfqI96fgUXmryl+bC4AaeJQvUJx8
0bojq4pjFeJz1tIDRDZ41kc4hQuo2d2GUKLD1KaPq1ZGkpLycx2DxxyLHWGYUE/nU1zWGvDPP3Q4
Q/EJWYb3rJeFMjf8/vgJxjRSAaH4/SyFgi23CpoorkcyIOIjLJuG7gho9/6WgV5ys7ySFndkI2oZ
KKPrlZcMDNNYqDwStSKAIsNcGgG8z1+HcJ+dMDCiYarK9Bb/xQ+x/g1I/5jjnNnyKgYgPpdr/REH
g6tIG4/ioLEd5tOccY+eCpJC4k/HfkQAOWlZX4rEJYNiFVV3BpxsmRTBP4pPfArUmJ+lJ4TdR7G6
+p+QM0zgV5x3kjFEPk6Tb+DaDEpBW4r2Ov9a/f7cTW8UJ08zNKzCg2OXlvMEVgoVL+SMuAzS6XdT
rKIoUyAFW9zgyLLEKHe6tjuTBejGxDnCMDeZNHutguytev66eHCT8i9nnxp8erMLEhg2JQxYidRq
wxnIm8My+uqab7YYe4d67V3sCKetWApbE4KsoVUZScKe6s1BRej9jhEWWn7ZQ2VWuYWcoav5QdCF
Pa0MawmL1py92Rclg3rkCK55y2IX8eZaJsLoK9eL5ZSphrvwlGd6yXkcGPLjp3cee3Kg2LOPD6bc
UcC2unlbgcHJvfSljpClpU0bQsv6i0HlN0QN9SPXfey3q6pOId53I513ABcUOQPMcUkPbuiA4mh9
z1t5K7y0rL/gDUIkUzD4N2YXSeVTUsRzN0+hASpMt5L37Cbmm3bOCAhcThZuM/59cvB45OWrLM5g
Pd0nOYJxfhtdZr3ilOCqlW2tZxH28ITH0CxPDLUkReMOEBNoukX05PpMJWZAr3P4Iw5TgO0OLaro
wzVT6hMlr+O9aKcwWpEjZ1KjU/NFktz/j1Q18ximFlTZP6JdN1FZ9Jj2h4ZtgxTuR7j/FS0IqNOH
dernP4g479MZ3lCqvEt7ZlD3PMM+YXwDyHgDlmPWrBJYqkKCEe8yRkJQYU05HczisvBQAFxpyKUt
7GZQBoe3ovlRYpOiE+PQQkmKLPXaAQmstRt7ooFAul7/r5prUhc6eguytGXlK0YKwQwdoT3a9NcE
z4g4yOzmgZ33ZA66mWMO2VP4KaIynyfv1LLYy7JfRSLijqTpGkMhtj766XovTXwi2S7Y/FtN7b5m
bPkwk/EhrB0PWQJoiaaBzdZdkkoaaypuha9jcKB+bPbu4J7tWfCfjR+qolTp099AAv3rfdyCruUl
swth7SdFzaFDbd6/smg2DBPt2pgaD+uFO363rFvjwdBL/RaxWYiBKwoCybv4DzdYJ3M8oSn4S+KU
uyVaI8CE5haF/jxIMeGLtA+ACrpQ3v7IP4S0xL4goEQCviHlqA7Zneay2xjKKMnznGM2kHSXwthp
FAvOLbDywyfb4xgbujMkh1mMQ/nwyRHO34E1j/ZVf+Om1Gnk9/1fepSONkH/4GxnA9n33abGyhQy
2E2vVHAo2hS7v9on7HQy3EwehOo5PCvWeJvM2PrkBcdwgb2KSL/YJSeJT0J/DaJX75pNRbxzzc83
jGV4I9DI5TzUtncWRYxh66D1LxmryrwGOahNpRmHCBWZ/THEsUJ5prwd6YZAjVd5kJqrFdji1W3W
JaztobIB4Sl9XnQTAx0jR8BX3VNt9HvjQWTwVhdHA3LI33TP0ljH4BaTw2KDBwhnn59trczqFeq2
I1k6fdXHA+MK1ydjWpbvb4MSfAyz9bsQ21z0Ofu5C6yavXKrDUDJEB1xi1dLEWAqorVM31PFCvaU
4GqwcEqsnETrkxJPkCsPokg3cFS/9Dd/A9O021yll8NLPbgRfEy6Ckmd6ENV4chhYVL7z2kZTjgR
4FjPRH9MddUM6W+jDxc/3nwHsC79q9qCrvO6AdxyFJw/xXXOvApM7AZiaEUQQaNpdcJ8zUsnP0r0
5mK6c5QGRSAiXUhOqwzHQz0fCF3xPrPola6Fm05qDj718Ww+UB5NJW3L5C9CtfJwj8dV32Ae/Dy6
Dqm2tqQPxvvZ7LjzYpLokFUxlqWaW6ysvVKR/s9wb2keIwT3ezU+chmGXYIksHSuOMbynU45HymD
7Zj+xYQ8tRvhvdco+Zjo6T/Zfa8gSymu5iv3pCqhD8XseK+oc9++IxoWpFKQemNjCHXuRcYnc1QP
53t27FlxaRQvdNtoYvTYgPEkG3rbGjid3aEKbwruMPnfSDeuBWKKEjb4/os3tBm9apaCuajxm1nx
RyYic2pQfwl6n3v1VV0GBxjajBFRC65okH8UmPf9aWLCAS2dL9oZxqUoEA1dcrL9cgxb+fWe3y5q
637VskA3aYEKD8+1ByrmTbWieCdQ+5UG8mdzlaOfiXnnMOs9maCIggadAMhTIAtQVf+fRnJxzc15
/ku8FwsYEe7RJRSE4PepkNnWk73rdY8reXCtGQB57cJ2P/Tgit2Dsf9tOcNWYGj6J0Jm/KpZ6ADh
qTfq7kvmZc6zuUlf8+DrFafncdeS/ZE7DMTQkbxb7GJwQ+7Pye4kggg5k+W7caLlehCG6MySUKrO
/WAEuz0hIPDzmSkP+fBSn72juJ+VwUK7mhuXHxIb3ssZkieqUZngvSyLOrt8QBXZUdUjfa+uRA2x
xpG2wPYARdCOtIYuPQrdRluqdGgwL8aASIYlbmewmDNYCreUWzlwtjLAEEfndWVEAUCtKKAnsI/D
dLgyujhtG8HWNnlqyQK/kihjzBjDvLNXG0zu0UPmSbW8ONBzoockKZQhb8x66Q22a5P7d+LQu/fd
DFK786c1ohP4iGC6a2UoJ/nin4K3+e0ik/rQVcapB4VbHGqxxCy3lC9NN3/ZS/H/g5avIMyDl6x/
l+qcWpL7kFAzebrJYs5vD3uD67zvXpXpQb90JfDC+6EafykvFXWbmDlyyhHvSwR1LY6VcnMEzp2P
YnV3CR8OKp+uZev2YzmGJLNAVh0oeBVcD1bD9oxbK9b5w4GCp8D/2qBwsBoDcosSJA/7vatKYj7X
Bdsg0MpHrXa/kjy6mPh0ofeBeADx661DZ7QNcBSgnaEcwd/0bTDFoAnvwnxf9qd1B9wjIW+mTsz2
4DXrsLmxu0HKrtaD7nOm8VG4ANnhtWjVFgUTbI12PU3023IcEWllVWin5e5vAQM8xVW34gIEsB2w
0H+7aIkzXtm5MltUZb3thpvG+/QGh4VAemWVsGZqbjm6z6xpvwy6ohkOrWKXzr/m0cIXr42BtHCJ
TcHTcRKGDJnXwYiSu5z3Qy7PIISHkUZW1DnrhvkQOdw54lFwsuwKCg6cLFCiQvsIRogMPlCCu1Y5
qW3Y4E79gx0ejepe39xm2Me5XWa7njZQ3jLumTDAOw1CiAkOX2ol5vYo5tkZMylgyoIWYzlsql9o
3pkX+BeH2ayY5ZQuouv3MZrWN27fcyU92rUcN5mKyrbjp46NKF6h5aI3VX51SaeEQ10bTv+cZovL
uL4ozPSpfzj4LBARIDyDydCtBHzad48UToPQBZACejLlV6TYlYm7PmqW+PrNzX5uiJTrleOs79Sz
1pt6TVmJ85k1N5d1KIGWVFslK1YBJsSfIf0JBrIra0Eu7eFaB+QHWnJqqWvoSvbqUcjt6++m54Gj
9WuDC2MOUw+LIqVY6yvcTuLh/rzbnwIrzrv5Lkttl0JcKaYF6F51oYTav+F+BlFd0/9Hz8AEDs5Z
lJwTYyywPq1Q1XS1a3qGpXlTRn/Q3J2uZEfQNFHdTULX5d2PXQQz0YwogfQ9sIOnkAYLkoKOigBR
+A6+FAxC/qaV6dKAkWUMx8ZyAZDRDOXNdws8CrAT2G/6oGquWC3XffJHJWcjL0sbxpmZ5iqbB8u7
cgerWvySPhjnE774XlrP8/bcTdnOQ4pIaVpL1G3P6o0Riqn/bl7ChRyre9jeMmNAd+lmXct4ZpEe
2sSfnfzDdc7itnkJF1ikuYQkTupj5nwJBqQzUslB/QUYQsdHZttUbwhw53NIL7VXRwlKnb8KyT1Q
kelEyxQbsTpj3WwT4/gU/v5r2sEd57t5lX6rkBP8RjwrQ+7fs9h3K7R/Qw/jegnNu1TI+YtklZ6I
mL9E6nmdcT2TjxUS81pxBxZ7Eej4wKPS2Tvvf2UqSLuu2Kuq5e4j7u7YeJx1pevE+dX5p/8Z+Cxo
QOAjPaugRuGwmAd/8AJioePSZ/80L7dpwBU+YSGcV3ISYku9m9CWESTv3UeHImfyZBGGiSkJErPM
cxZc9tqPXx56I4vjgyABdyuhpkzut0omC6nVuseve9AQBzBMyDPW7hAUQNv2eoCazLWMRvpY9q+D
KCxtODsx6gq9urBS3YXCq30LqUEPp6CzKCCEMlGgxxTSIADwnSJQ0B4gIjI4X/ZmiLKQCoSLynZU
EbJUuegrmWjB+Pztf9atcbbw5uRWE3U76cpKtc/NRZg2YY4Tr5w8bYKMghsDV2NxiDqAjRDAKy5Z
f8PepZn8xZ06LpTdVHrmEM11MBm23uROQN0UwyNK1udHQ39HOks7g0J1RXQZeQYByWGt7x+jLxdS
E4dWRqBrGFPNk00enDCDG0wqnVNAAaJwAmJM0a2bUnUXBgRZeHU5481NJWRfgPflkPMJMiGP7EOj
PxlhF1aOwQFfvwsfsnnt41b7uHRZRLN2Q5MdwFOlYXF3O5h9hIB4R83rgUycFn8EfV8eWZYlsLeF
Mx0bzUiWuhhGU36/I2wF0aj+FO++XcZ9OfyXYuzNzwZO6y1CH/rFbnypjYEu+4Occ1yJthCle6gM
hwLS3k2yRMhkZlpPLihNXUCHnPtvuGoRFjw9ucPhoYpIIpcrRoXkih0AuQ4vMab6XHjwBMPW5Jcg
QD5ngRdijqDx/kYpxQjTdYG51hpl22SbDa7O4GwFqoFGzoZ+ERc1yVYHox3IXNOIh3dh0tj9fEJz
da3Sc4CG4Ye55Tn0pisVYADhjVYuaDY8xtEeDIznXKWWMGDeyxxlVeCCGHN9YkrbA7dfCVyfcF8g
x/Vmo7w9pOvvCxilZOyfl3J7410RNH2Kxn/2tvyqKp8glJSHt3ixRWnxCBcuWYurtKa+PMCRyCVt
NkeZG8aUdTWJBV/9R3ynlmQZ2KUl4CCqKSLg1yumuWn6AQ6YODUf42hfwaVFoAeQ3yyJhpPxy1Be
xZyjAj4IWv+beaw9smlQZ0hCSLZg8dksxD15aP+Fjtnvz3YjDAH5vhgmVMeA2ARJbZ5UymEOE6rR
LFVqHUVCL3a57mTY4o7gvOdJOM8SjI2tmrF2NOFIHkv1/kDZ4lAbUJvt0JlqaUMgDoehjbvg9b4p
phmZ7eTnj699wFffXEe1TcLEZvK/uocDm3EShgR9tnvLYBpHzelY2VK9lRlyqLPI0CROvkmTAotO
I8qUml0/BCoW8zSi1uskyM5cas8Efgpx2j3djXbuHoJ0IIzdNQSD+fCgC+23J770c5OSdhXpS63v
5+wU3oDvdSmml5UJFKM5RKXd65VQifVnhFZIjiPg7ov5QKoRWNONV6hJUpsu4IKR8IXBON+/Wo8a
xrl32K/aScT/AXfDdp04Y/5KZtE0hFq6u8mHW1RnNfhlneTmPG9dX68Uly/wDwJTkzrpec+KLAcC
kzZvHb+BZgoib/MK5MNuWQ6CtInkzoWjDy2DVuSi+uAsqOpDNfMnXSh0BE4xO82f2W4fTf+jnR51
F6Gu875YC2FIZfmskFZhzauP3658QerFawhPeAeElSPBIzpaZZjGysin1bLFAhq/bmBj278XAiQ0
ERxkFHDZNWFMo94VSo9A+yk04l3rYu14Pw1hqnheK7AffnBE0ortI4nJL1KGbHTnyMuzQ5P02kgT
Hp7jdwm6S8BMDXjnD1f3ZeetD8aybmXKzTH8mJkrSzJIms/9/FVl2ZFGx7X+jXMsJxAlBwg8Pj2Q
xwFY86Exf8pcmF7NIu8dqE7V15YhWSxvxrE8axvgk8h+bij8q2TRxBGupbWSkvUAhu2xcOcN/QhK
huezzbOKAR1yg5s+HzKOKSRQyQFVk8zJ4/+xOpyMWQn3s5yeEmsa7CJImdVoOheGvy+ncDEW2+1P
2UoTqLStshNkxdw38HeTZpY8ka0HSAY0ptqUofeZ8mkyefXNgKTeS4a0/tl5aeMs6wufAVBqPBS3
m7d7eBGaofRBMBV+EEbZ1OfQlTNaq7ygjBZ0Gu9xJ9+2SB+v/IU+xTn54fX269IQuqVUhiDPZhxP
k/3U1bHqh09gHQnisZN8O+zrMEhbbiWp2jEN1GmXSYSVCn9Dto9/osUXtatNYR/JG79rf8HPruft
iMKFYmuh91tlqnNldg4GsK/WklaCGJyh3XO+fqbShilyz6o3GZPSSKF/g6jVPimReYQY0mB8Q8WY
6Iww2sOt2ZuAutCvw02HbGeA8xNNIsJdqP2Mm4QjceHi9GE457i5qgSflsmYzs9WqPozoRPStRKh
M0ddC40Ck38y/xU3KlDm/LLZPNCApVXtrspvmL7+1ozSDc7y6KrTfczotBAU/nfzVlllOd2qL8M7
7ioe9gazE3iDNHHSLa/I5Oygwt4593JTsRaA/khRyaGAZWtn60CHAMSn/AXum4GjjrY2R2AAiMaI
wKPutljWdP+QOSKCZmy08QP5qB+sg+ekjFkyeD9QoPw9WOHPwx/PP6z/l2h1/tM0eI+RcfwcPxvu
ekrFSotzAa+GwW1shdO/5CAccm/yDvJXAKMDc3I3+wV59aRRTC/zTMsGh78SOh0VcJv6/7wwG4kx
7kRlldM/NR9hCZ+ZqfVyq7Uy4TKo1F1sUUa+/mO1iO/0Mk2GJZdotD8ziAVhm0QGsU6Bp8BZC6zk
YTsLZPd25nHR3aSRrKJ9GKJ/lrGfkiSteU7R5n3eaSiVi2OWIrYyg1boHkbGo5Q0N1TduMPJkqzD
atr85/pVHc27AaGE7OahiB1ZEpElYTrkJwQYE4DOLK6/FRtKHEP6ote2oSXUK7vuT2BVWvEm6On1
fzpVP7INBWP+259t8zqcg3a9LYVpFC+7Pp9/QdmnXSC3smDLuSELsO0bezAybOu027mAWItBPbvu
QMsChLJ+tgLVXidGgkoHFzQz8op0ABp4hwNj6j6Jw3v92wnw9VkS3psz63E3NZ/NtXzE8n3ldKDC
SjGDR9LREsicrInWLJ+jzeWNU+rMmfTzPUzQpf+cNOW4yqNy9icXDqp1f/rfgQHoB3D1gYLzWvFf
osaHkA2sXae2luUUJczriFXw4BEN/HdGfVDtd2lZeFp9OyWdV0GqNkF91ilIJIap3l+8yIfE479l
Y3wfiR4tGD2I+A8aZdDdVSjBoLTp+7xsDB7yr88NJO0lLC1p1ReJANxBRCyoADqdDnYNajdNq9mo
yq/28GBGc44ZPxi89QPJ2huaPiWyI2nIx/azqy3bf7DaH5KclAAY+PRfr82xBc3+o8+WRa3Kf2Vy
++oTmm0FSORKrYKo3U2oW/SJzcOBYzMR6zLM1UjMYI5NcRa4doBbUNomut9A9jSr+0tryFqYnBzn
WzZAubtFUCi+s+rRIpvJ1BrzOi6Pve2/VGQl+mf9qAPxbI2PcC6EnPq7yqycxx/kZUGZzeVqVrmI
zKrVUtXK2vwSPfTxSN8OXBFA5XQ72Y4HNcLVfBW9nMxvHHWeZ8laGHYHDGO76DucigSf6nxfn8Ta
zHNAvW5EiEXDy6i4+TC5pX4HmphuobFaPt2GJWYbGBOS4T05hqpsbR/M1D27vc92kw7SOxlEybgU
IrrN1+o77m/xn+50JM8QVw7WnAy6BnYg1EpEVvYiCRuihFR4AjQo1Gmu2iAm5/idiFyLGppVHTvP
ySMykUBOXytl87/IjUDYmpJkw1tjDdaPfDuQFc2+wUi6md8mfJ/FaDS1qsGfxVLJriRT+N10Im3c
lUg+paqYa6Y8wGCLWfAO7jLgWU3Xa9XwCIURWtmc8rN/bS5Kur0sxfmzzGVksHOPCrrhxsJlDYaO
PPmLKVqRdoPEMhyFhW1QGa2ihyithgBYjC5v0kkb5F0TPHWvMbQltoUSmnh3mN5Lp+igbqilJAy9
ykgQCr8cf+HI0diyiG9tDuqNSEUuv2YlF7Se2yoOoDP/N5xe6KCwhH7/9go77G+AipdVmEvAm94+
l/eAtQU7NsEd0D/McBvC+o7Psg34cF32BypuGpYxFuefMhc21nfef3G4KOobCYpqPqAefj3VZBpg
pYDPGiYQI+cgV5/DWjHKDkE2fzEJ9PCMJI9R3lCwlxeegAa//ORvAczeRSdKuxpt6mm4l9hw0AS/
tJA9D5Mpop+ywf7Pfk2vIHZnVKZa6mESdfBnXkg+FbV1/Pv534oOcCHb669/jmkItYtDifuf3exs
f74cXAeMjkW0UbzEoCYIPmB6xZG3qTESQSFc0JyRLykJc3ULhkW2kPA99gcLDy21rUD5r7corlbY
R5+jO8r7X+MxjU/u7BHvhYUIzlpC98eSrpA4pCRaBBTOb27V5JvlQIBryjQy4YNnwWIf3IRvd50L
kElsZ9SmjGikDyJwQdoqGUBRR2YAA672Zpc03wu1a4xuUK1nzDsi1WkMj8GX4Zh6QMY9Z8xvyYDW
xX4iyDNB67PNjDRbJJjQ8OEcos4wSYJ/f3n7zaVw8zNbiaV5dFF/rlEqL5kJu8/yND/5fE1R8r++
bEVNu0UWn/D7cLO9JFKls1sGUVKKtyqRejPSzKisr84i7UUa7nwrBWtYJZ9D9WhTDXDK8vkcqUxL
bO6NP9+yqof7VT6mRhJyIeDZD/URuATHiyQ1Gbt4TlAbM6Cu5L+Ljy1vkoPYl6VHkBy0ZxP9e9r9
JXe4avFwft+IM+CFspARrC0dZCvTK0qECPsS/+94s3nwjLWNFyNQgNZABELqyWs=
`pragma protect end_protected
