// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:30 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
nNlXVYBHR0SLQU6TOUCB8H1NDinzREoqqhfNNnYwMLU4tgcHR3Cs3i3XxVxqckPM
dIxU0l3SVGhPLicc7GwpmsI2cLacIcp2CNa1jbN4CcQbaBTGUAVIykWoJXGDpRF2
pP3slH8XyG+DBFq+zU3g1AtD83S9Vf0ilOjite7rs0g=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 19088)
kkn50fqWOdkt5BmkB1BCVyVHGHT1GFjYuFBBj8SipIKvdSK1Mo87ALpO5Aw1PGEH
P1oa2k6PbKWuI7yDzdNkDwSGyra/HA86Gow0/7vi9nJBSgksafouKEusIr7l3fR7
WObCbXb1T2uxeC13xhMrbq9BmVm5bV6KIHpBt+TFctTqghfGxnTEnW/fAh4CFy9k
wazG9dYNDlCiipxscDXweB2uweBBrDSgn86K3mQwiHGLpmv7pKuHsdPYYJNJWtlm
9hIsSQ5NxTF4eyog0iF3TLWxo4krL0C3rgJANeiY9TU+QA/LLsZT9XWQGIvKOHg6
qb53PB6bZWHXawGuC+2+14VQT2CGEAj5njxVyfx3eekQszwejeTFFDKo9oHs3yr9
5kVHDYIA/0kNTUIOmwyBeTH2Bn1h+W2QzGgFpqdJ3k/HHuKhgsPNejvzsJXW37/z
4UzNonzKkhKdw4E41fKqbYNJ+KeyQAFF2CQqQ/Hq/YNZjWj/Z4x4laeoFQgrrZWE
siJFm0vK+4v0SzeyYwo6/5VXqQbKUglq5eoRfygAo95/vmxSZgFmQmj176AtpvY+
bYNpytuJFoQ5mEsKA/JDxR9/uHkTD78PlOzuBikBADmvrPihiDfY5A7zSTpfyT1M
e4ZM4COLEvRZ9JGKk9FhO63LT6fhckOQtbhvs7SK/2imz9sWxr716OjGn3Qfldxg
oMmb2GWTWUGNuK9mHkwZZfbORDUYelx4XJWDbC0jqID/ZGbI8rQEENID7EPE5AHE
DFkawneAW1SFk1s+u/jFo07UaQDCES2gW4+Tq+khiGW81lmtdV2POuQBP8G7s80H
xq6vza4sr8UoVmJdA4Qq8LZDMXxBTlZPgGI43zdw/KSBGB+aESYJmAbutZY19Dvx
dpnYcqc2oIpym8/s2VIxstjOx+HSFSLPGKLZd7Ba6ziXDDQafJ38OvjkbJbpR+tA
a23hJ31G+idZyMoFrogzh7J+0Mf3RtIOkooalgFSNJJOZjVPP+y2uq+pmz+3OMJQ
GvHwovEu9XV7p14J270vN4+sTQFpZHEMuJCO0WplTP6xGvD4/llseHloUr/EPl3A
eR8SzGLLjsNt3IMbRcf4BmRebTV9K1w3B78U+bQA1jGEuyKwvP9CY1/ahnqD4auT
ra6lA1COicPZHs3fFOk5p0XnzRkFcAfORHJSiwVQcXCj+OexP2+A0UAUC/bPecpa
IhTEj9tpNfHVrWKMqReLCzm4hAt+jBmYk9ClFAWlY0NoIjLi68rAp3wYunKK/57p
f88W8Cza3V1hBasJgW2OhO7W+QjYMLmqto+9c526nXGaQndXo/666+a0QtMDEw7C
CSTb4/5dbEK8fj5bGlV0sH65z4MUxEq49dRnlHvB44a+oNcmiuwxPASSrp0iFXPW
xSXHW6JAoJtQsxnhuBjjBgjAlXnvMTxj3LrkMOYD3NuCfc3RnunPfh/78wujUEZC
ekoVygJ0iLq64daXwwoOVLIctpjTBMRjoY2pAPCAJkb6xQxnMf1WOVegqWB9SOCT
91qtRGzxuGISMnM4mlCvd/aYu1vCf3itKOVns718SGVXc+mTMP04U9rfixuTlk5D
o5mflxjDNgDE0UAfkTBe3iVnxGc92tQTOmQ4PM5KTUOUDw1v1xvMiTlBBzE4T0zp
hklIIm2pGEkz4IlYFU18JmkgHnVkqavrMo8dOpAo5A0l4FeA0JzBL8vudBu/kmxY
2a2FDSOeCdEKBSEDyTa4gHA8QShbT+e6JxwtBXPQk0oerZOCgPMlfdrq35FxQkC5
/B2rPZOZt/ipUgwlgya6xfvoUd/sbPRM8DXmMeb1V0H2jOoj9yjwIvC9vPbSjJJ8
oQ9AQK4SqYqXwegqQCyLRDmBypqTxxhxFv1qNMmc70oyUcBUHZZtAnJ9n6B0Yfnh
7e9DltACmowns8TS6dm2+grE8/NK0l429EMMSY0NJWhchge9gvokyTdio8viKSrw
IOA8h684MdM7fvlHOmwVzCgkO9UamocetG12JR3tUSWjRPKip+uubgAHA4zSo5sg
rWjhY/t9Jb15zeNJtfkNwN2Ccflr/QMSLpt4CoXrh7xfH+LSMWsym91IZNei2vA2
NtGTd29F5Fz7xxs9qMDjnsVBuMpa9Dkasb86OZGee6gDTGOv/ocoMo8CvLODwXgU
9noWcqII0LKQFmGmJOqS8wVO97QJiRgANk+JZgpQ95A7D012fsZ0Js9ITo1IPrR6
CIYwg89f0jhnKWZJs5v0uDFHx0O/gSU4IJjM+WHJ8UnduOX3gVNRTrH9lSX7vwKD
b+PI18LMPejXYjOFVyWqNOcqC6AW5jBljVulz/ysEe54DG73ClCM+aj2fiQDb4sq
WqVCUl4USry3IajSVQru6wXWAgW4cCJkpUB4yQtNsRaIN0hTR9hceoK+vO7x7/Zq
ONNZQPBquS9P2dqWpVTiLJ/do5qS7/0AS5EcZKcALUehCM46FUxqkO3kWSWmGUVG
AKkPOQcKuuCoE/9EnyxZ3T7PSkTJHMue4r1wNAvyZ3EA8mGs1ub1/AH2ZXaggznf
u2V74NfmCX/k0gs5YbeycQ7qOgu06AUr1ToG914xc9N2Uz62h14oKJkZVj4xnR3E
LCuD66wTKmkgdY6e6MUt1v1Qe5PNyOVCdt2GYAf0Ae95RbSmUvRMjlGbJ4ddeOeA
9AsVywV4bKuDWWwS8TqyiVQwo5PchzLlrI0p5shawhD4A06GZVJRlpxVgauBq4S8
ly/xZBgwz74z3y5ynaZfUxiC1vhMhcYkiGcsfiK2D7tjcQ/ZHK+TpQOsnoKMCR/d
UXAX/U71KxvJmd3tOtk39XaC7TEx4VumOXWVg2Xi8er5a1YY1ZLPv2C+KoxsBJvh
HrDoiM0yBZLYlzxObMFBf4XKvhIrgq9jbzIz5HUrWqEfFPb/WjOURT1X+DYank8+
q9EepLjFFHdo/gFwjIKI1BZTAqZOPRml1oFNKqGvr3b/2ywMqCTk3FbPsUYrNa5N
iKFE1ysTTMugGZ1VyVGAdvgU1N3+eie1bB/LSVGDgD2xpTVgSAdFgcLFe4NmXXKj
ra874yL+L2WKC7axKQ6Jkim9VDBZwvO+nDHTgN2bECdoHY2OLAzC8wvIfqxY32RH
gRCQpziaPurHDWzxtFBZ0/efE7jdLnPR8bZE6NBTy1YQvwLBEIpO8vdWvXvvYCiI
aS6SXHCQpmxRg7y+0KBpBe93LuZHbO4OVERFOnW7ITzi2dqud0De2jiuS7CX+94j
+YkVxVsWszlR+lQ/JwhxpfkXuZjM+RM4OsKeh7RIf0LMsRhe40Jw1oIPXWZKxFPP
/L3P9D1PmfRFWQBkZm2X9s5nWQCnU3/4gC4H0IpmdErGOLxXzf3y7qlDxSfxt6Mg
uF3b6/y/DuyABYuBqeHfvUB08uzIKno/lRT6RapBLTvYbgKVQXZisOTtBGsPj4f8
OLNu7xeTdzm1I9IGnRQ8aQaQ6LsyCw5U4rWZmyCX7Qe5ow3kXNroii81HtRY+N/q
3BOfyUYfcd6DtKFuhn2sPEUZ4cDU/kdhdZzc1P1ItZI7F4h9J1qF+VmlkIY0qV5z
++6/+ExcfDL71dBMB9Mg5NTePekSCYKMPH+qiY9TVKaJMV226lPBH0DWEFQes+kg
fWlpZ9MCREMjM/7yxEyWgxDKVHDzPDvHNDHE2vtYIKxhOJux+dA+DEUBwyIVcYWR
EkekHedZhissXppGFbf3JbgWH9faqbHItWHpKEmE7ofVCfmuFECybPRwAIcAErXP
Epa6k9SM6dZ3+m1vwIKzIoxhJMpw0Kcnd3wFQGfaKZyCD6QcvYTDESqOy2dNP8oP
4+WHU7/MD88UH3XprrzCq/f/HinQClylXv7JE+Vb9sX6Q+6qijik1aklLqVd3EHe
Tbuhm3rPzjlLG5302NxF6OPbMWsYRxvRN9sulQtcrHxft5p4gV84KLURQQIONApu
vCdH4QyXipKO3JScPfRIkJFkfgWGckp8Yihw4b+vL7A+Qxg/Wn4VZd8D6OYDmuGR
EJ4MNyd4Ga+V5WqAJn3bGobWJtqkQQWhya9kZDxIEBSMEHYuklOiTGbZ7v7qKm87
iC1MoJwwz+H/SdOlJfnPxgLOD/C91topHZJvdHTUEYoZ6Ks2z8t0inMGr9jZfNGZ
yJp1/MVVQH869eVd5RufkEtX6eOYHjEs9gdH5bKbfSbcd89KhaeeP+1CWZstc0BS
jdL6Nk7gre/osF6v4ON2rhNx1F1UCESfkr5YW55gDpUQFkFrIZ4jdPXeUsHGMvSy
eZZkUfeI4eiOARjv8oLUyCUo4RcDBcgnV0Obif56k1ozVjkoAHR8DZJ8A4AorKaH
yufeULDf9X2v46as9d9YkXbnd7foFWj8D6RS/F+KejAkeXeunLCYGoUwbpBuTqFL
5mwLPbomycwraacdWaLzbOlRlO8saevxUrXVASSN9AAIWUHscrdtjXcNIqfWN3Lb
UnrdgnMUxSIohB/dDEZrnbPvBWmdGAyDWrqirc6DR1GrlpcjfTvyx1uaVZqk/Lan
To38eeFzwXRj17s52ZNjrkDDK3nV0o1A9Jb+p2r4saz2UR7oVJt907AGlVfBC06p
vjeU/4IeZ5P2Y4Mdz4IicN2IWTwk8qilXOcnvEaoRD2njWl/8NFb6yTXXGZ+sa3n
kKwGyoQont1YgdKLbNkqAjpv/UQlXaeiLcit5Ukt2fC4EINLd/4ur+E9Y+aJ3hb5
Ifjzt4AaOW531XK3kvekphc272a2vkqoa4jq6gA8BvHRjBiLCeJFUWGgQpkflWrt
S+lapIYfF6Q+BzmplNWN3aOe3R1Tz8nvWi22rVQ6KNZ3QRI3AtmG0gQ8jqrbrxD6
GvHy4w34o/8wLUiDX7Rfcaj/Mrwh21X9huIWDghp2w7TBMSeBJur7CLtZH++g8ki
8Twwm7WAEJGdFWfcPRPcFi7WADYOgvZ16WeBvGBAF4iRQHsTS9NyIMepdVZBlS4I
oIC18N9Z0EGHlh2bv9evuk7/EzlcSkBfsltxKwaARBjLAFlebWLu/Bybmt6eGqJm
NVfF9KrCpVVlFLgJ49myJfJfYyOgft9NaNHdKIJQ41ljbpKDt/XoImfsqnHXvq68
30umtGL7hvwm047TP5DkRzP2HYTU2n7LutN2hC4nMplSj6S+CPSVwig21ZMxF0kW
MdUK9gFiIC0EBm+oWLhSYGIlUdQ42lvAtZzGhQZ2ZSTI/rFiPf548+oYe9Q+m0EQ
SO238XXX4E1MB0pyu/vai2ZwP2Y0jo8qZLD4jM87Xp7wPS63MXqpcBW1JlSXNGzh
tChqeW6oK0nuvzsuTd+JtvQTLFwdiUCoeRZ6kDyg2OlRt9bRPjmmV9ycUuS6fH6t
wh+MSVQtjMFPBeY6zK47b/vKhSzxkBuIrcnjUlqk44LKCR0AZgZQkLBoajGY5dw+
xzxGHPf+QOAGwqnjiYu0+7k/2bjlLAuQHs9aKcXXWu1nXag2r7LiaLNeP3pQNsHm
Rx+PAzMuHsxFDq7lPRGF/16B1Ou2wyQAhqDUF8goFPH3SdSxyWKOoAuquYEXzcQY
VNQlIgad1IyaBbGtWWO5jBSwioJ9YPy4LeumByomHSkArWNEEIl6MAn9g/+yS7li
lQ3tD/ZaXBqRKCWg6StorNRbE2QrTlSeVu5r8mbKFsKc5nz9juK7zdGJJVooTXn/
RI8QMqlMLE2tpSdnx1wMEPYVo6cwxQf13YUwxupcDXKAoFOFpiZrI/YKRtJnFhKZ
wmP9WRq3VQsuvUIw//KtkB/rlsmj0g+bH8iGMslchwyhIygjbdXIxZa6f75VJ3Qp
PdsqD6u7dsHUfuLJlJbFCYEChelHDXg98IgZMblrmOjRl2m1ktHE8klguFUsxzMX
7q7JknzvOxL2x4rLj2hs4gD3DGFbEXiiTpUzaun4RTHNeK+d+67yFa48jtkI566B
feFhyzHx+O1Ja8CsCQ6i3dh7DCOohsP5/kt2kMVeeBmPOomxWtIvw4MO3oEEKLfA
BtNAF3EzDIH10Buf54WJodUkxURhutsp4F/HYt6RiCv2Rl0HDz+5GmF+J6L6g9rf
5zruY+HqSvm3K9bXg5edCK0KgeHodd2PB29sE/tpO+4sgu14F9jYtcD3kVK0kkz2
INtiq/EGt8+mU0BsoOrl3PA4Vf6f7XwgxAGh+scOi6ZuYEUXTD6z7+LYQjWMGENB
g9AJ2+S7C0qkOsIM5IsrPZ0+5YSugAGf9r1ahd9d7vKS2nvaleFlQiPA28uj/xDW
EhF5UkVUnyXXcGmcuVWWqbSaO16LNUkPt9FxY7dRUtIkVyWMC1NCkmIOnxKeZ1N4
9tiORRQfFXcPVq0U+K9JwhtoKcys5CKimFz6FEYpdd13RPwhmHMa9Nyfvgi3BQPA
UHXGpehXavtW1qGnca1YLFTioVlXZwBxM82f9NvYi2yLMU48+nt2ylpV/3eNSq2X
aBvUxisGQkpoR+tnKOO0ArotA2/Y8kwu66EZRoAZl3dkQU04lPrlZITOiIHZCYjx
iMjHCKBFwI3CHy8eQ9Kx0o6m/SmBevgK/LjtwfANhlgJS6jWFRLpLnCB0gc5MoGD
HDSZsRHIMAjoopn2wQzWiP9zykT+0MZnb1Uq5UwmTZi1QN0VLudaLnzphjNrG3aZ
vtC8wetNW0p88znz1bkwWuN8TRegRa8+fKphKbmbsyxUG8RoDVOt0xVS0AYEVKlr
RZYLc3n3Inlh7/MDS5g9TG9+L7es1FnNWVy4AtLmDuKcx+3Nz8fxMspaSVq2mM8T
3SeUGOflVq8aZWSkG9PHZLZJjYB0LNnVFxl+JKtVPpUCpkIIaNCJfNH00PvHqGzL
CeJctGtDWEWjRWmXPmdlDTr4zKNWelrz95WioRulomlohMZzsIIFk3YhsLg368h6
clwtwqx5oXBjI0iBIdttt65TpWJpItuzFOAPXVhbn86Xk13P7mP7lUPHjC9tHDAJ
kQDsByYiKX9NefnGRObrOU414TJQYqDYmHKm+ssZyTHOKDDMK/KW/TpPL26lAPqJ
1SPD5bBMWxRdMfDLObGuIuQs6vP1Po7EZELEDexjcWcnDMam9dIsCyvfu+eLWvTV
f7oThVXYUjPK28oaekLBZWROYOOch0dO34cm42xEny5iEu5CxvfQT43OxIIQTNMT
ejvtQNkn/sEVxHJMRwodjQ+XINaKnG9ZLjLlp5juff8gweVb+VEaXadpgZOjaSkD
3t3iKaNhB2KVvF0VhOLQnoVVe5NYZXhjG6JsohU5czsGhPm1H+TzAdjWpg+cg950
MKRH/MB0rIMb8y/5jD0kfK27azHsdYvRcrtly06IYUBT3vMbPctLCMtLuQLEsoE1
9eRYcn8jlHj9EdJCtHPOhcBiby9FuN2gOXGjFM8OEgkaCqDk8p+YbbjI5tBViTry
/foR+FmEMpGeIDFb+b/g+PBCckq80gl1OzRrJ6iV5LnU/UJFBhQivoOrL5j2+rse
BTsjwtTDDP23znmPDMsS6VroHebZv6oaMaYQyvix+4raYC1GzAnr5i2wWbdlT+Gd
Zt+fmvEBthOhMlt6gsdNwhoHaEzSXG7+mSvU2GcWaOIeAmopZ720zMUKLCMkEmYP
T7fsjFT1+E5/OKACkxnp5Bh9XvKaWlseWHuC39wQ5hOLqAhR4kQTG17yCYVnrEKf
uvCkUrVeaRmrkcxVuPWBZUEtwhFTyr0kePDTTaQHkcZDD4DMJDoKybPu3zg9DeQO
IndABg3Ac3QdgQvh47L5z4Q0qzX/Ibz4Cs8a+Ysb/A5dkkmKA9ck1VFrkXln/jiI
2/lLBosDX9X8laQZr7KvS/+tacVu/H5wVSgdmSI2/5Kq8o7nm20gcM/oaujhUuZX
mxjUDLel27GprSD31bNAcENXq3JR2YngyN63gNLVD391j3aRwwkYExfuphFozGr6
SaymD+hEuMW4EPsKTCE20MdX//yt3R+Af4EPF2Sp3MsUUMC3KGgYsfBbAG4+apcj
H6jBnZwmGT8LuyinNsdxOYCqxD7VDyV7nxs8pdEvxdqx4iZPBIfaSq6lR/IsIIz6
opS5/yvNNLqfBUv2HemC7fioyFmchxdL/9bmJY/fhlzbQUdHL58CR0B9y8F/an1e
Y0Yrpo4PXrMQ0+woj/vLJlk4sxwYB2P4Heb/nxJzlHa/KDVY4ElFK7nIvR/1N8lj
GTxsZCRy17yeIa6UmBEa+EtfSTym+CYFmHzdghMQ70o1BjzXhPwblRGwLCmOqSTH
faJzNbxMG+3vTCp/2CHQ9YUF9+25YbuoARPOvmBlBZQUBeZ27ZxZNjgI2sM6vGC1
aW/qjaPX+yC7iMU+BJwLaIZZBPJ0+0WAHClnqsznG/cLNSTjpjcPs4siDXirdKhO
vHn/qQMhhhsoM0Sq7oT6f3fjKwta/iOiuBjseMXAqxiiQ7NM1FiSQ6tI10icIIT1
Sa88mArGJkpjInYvxpRNrSXfAnnQ+//p417cwWK1WSNflQZMZSIlZOnatyOspl91
mpjpslYuxY9tyMbwS58TA4/9g8ub8j0jYHFODx/YSl7/41bqXmPXRD6Oa42LkWuS
7dfH4NgoBhWnAHWBMSuDDaGFvQGMXuNaYENrqpS4K3IJTHHdO/URbwO4YEw2Wx0E
+cLEm+Lf7Bz0HRBUnyfFjYZP2OpLBauc+1FGe81fx4ooXESmG7Q9EtvzeE/6RsZd
rkEjVnx3xbMqaAFe6Kyn0upV88qA37J1pHdNVrlCeq5ZRlwstt0CHpllav6m+1vL
73SKOZTp0uzDv7xBM+u4gK+R7oJYjgl0T9cbZTQlAUyGpUjnKn9OI9BIQgxjX+jk
0fF/fqPsM2GxKfV+2Tv7IixVWrjKTmY7B5M257rtmcYaGdiH7paBneSmqR8WlJqi
kBxepdFeZo9tRkBt5b5+4FoH9rVdlyPYsw0uvvF8o+aLzqxIq+hJNeo9N7cDzfOa
oT747qG3xZTO3ICfp6rE4AGWDSyx/Mv3JquZiPwTWEH9w8XDCHQUhmy6othGORBb
ioUjV2E2Fu8Mnc+dtoUqaSyVSivLL3yEYbLXnKZWq8mu9hqFflOkiuCsh72uIxhj
oCqndsaaKyNRKjWuFKOMB/XqTHupMaNlPERavODKUGr3gxel0d40mvBo+aUV7sJf
oXWdqRfQGoMt9WpGApsxsmMFqulu1SXayoBIY4n/gJl3gAYo1sHW/r0GDGb+B/J1
CnkzPTluPARY6p21oIJn9Mw4WGC6C13SNAEmoyFlHS+NXXke+MtDYX3s+VW08qxW
g5t6EQsIjQBO8Zq3KHsj3mFROoemzrGePiZQM5DhdGIzfpG1IePfEaKDKk5fXppR
zUHes7WPkB7BzLFR1TBIkFruNZbPljFJMW4cR4IcRHUGow1xC//pl6wEUob2tzVH
InHoX/oEbLqPhNx9HGnw5q71W3FQh+7Gl30vVwi+nPJNrw2vb9k8MZqJJL96YwAy
NwEf4LaWJf32yr3dY3YbGfJJ/eyVixkoeQfb7Sygx2tQZI/xPWl7r+OsGSw8cT5M
cj8nYcoByOB34UKaZ0+BZAeIKgvRE455OAifBWMvn8etwiF9A6VNDZJ0NrDzC8ZL
ycmoOzPHmpiWWQoCnuoAbmsMQ3KYcMIejIAsHJfd7pzR27W/Jcg2JKFV7NHVVqCC
DJyo8sxWu9U29eOky/qh1/9OWwsh409YqLvFyOrLQAWqiF8UKwMBzRSROEABDUl/
brUOQ7Lnf0wcKeYr5lrPj5pUNPmuMSsAbAOVC2Iup3e/ok/w3UObyTVN0FcoZQG/
3qJwcxTamy+j2oarll+e2Hi1IH02VVBpCZgDzG3foee12rgoiB9SeV2SL+0Wfugv
EwoMwGYSgSHxLmfe/+qyW5w0N9zXCDza1bXxxQJvNdmMBPAc5beEJq0QqavLLq6x
QlMqAWPMwCrpQskcmiDofd3tfnB7JIqun/LyKNTRYrM8TFudpwcPkEnfs5tkBcZW
/zR8gZCtnLJIgY6zZnSEoZUoY7UU2vOtAg4cFsLuOhHQDWtOQnbKphartLv/0hea
uwO57tlv6mysWAx6rXQuOZ6noo/O/qeXSBfxQj2CA8wlo83jGYyU9QPWP6JhmZuj
985TuH92+eKzBWvupOR75pF5a385g74EWax/VE8BW9Zg7beE2FtpdxfS4IA/XDLH
xzupBoucC49h+mBR4oIDyJQM2M8HYXa8TYUypj08BTDkDzdlK+vYv5Kl3WHfQ0km
h5FvD3GBdoJcpT7vxvkqZDiSskhmlEoG/p7ziaWUYhGiEk7Vd8RzBplM8+Rdvh8N
nNlD0dPBVjqwfVQ3KMMzIs4344IGWJls0o4wRJzSOpex9zMyJUNHIV34Xkr585d3
VxXKKrd3SV9LqHYvTgSjZx93Gz7LHi83wnI38nX3HOogR2MvuLxDyQYCpXzctYql
HxNUcRaEySXmzOrhEd58X+HxFM/NdPYXWGyG8irGV7tDIyBmX0zlWmpprItClhGu
e1Et1G+7WznzMJRniIk3jIFfDwIUdy85TzYKPFm42nUTxsQvU//tdE1OrF9E+fB0
lbYtBls0zAX4IcN8GTtlnwFoy6EGnhI6b7uclR68EXChKGWobdLWJ9PuolhYgGHe
gq48Ah+PH+g2q9cFM/yb+aqKFhBuFRhjGzhNmiJch/KHTcI0tmOxrpCUVRwmQaqo
Dzd+BDFO9CFrXWxAs6Hii+aFrBQo4UZZ+GzFJRtUcgPeMl2/nLh74PtgOZE6IiJH
bE76b/kOvoSJCRJYkkjfj4l4nhxPn2wrq/8+uvJj8JtkJtAfclCaV1mR+R2DHWIw
AGuzblrXi6EbETSyx2aeA680hdyhDj6xHg3RtoDZ7990zMXkvRcz/pzB3d/cpCkF
75DsYj6rlPjirvJ+hCoggtnjEY4/oWA1FzNB+ZNfAzxu7IAyIQ38T7OtJuo51C+W
vgTpkXTh54OPVSywtvpahZ05Owbnpg5rtcGH3vlMACXHx7QveuDTARucAkl3rN1b
2tr/axoHWB8PdYLlyM76uDGSGad5qiJjiDAdDMBxvuvw4uXzkCuhe+6R0vodhipA
7v2sXDaiI7tngb31vshTAPpF9DxnkC+vlOk71u8FNSE8Amprrik0hQm7NHVvlU3L
xN0A/bzMlRRlR0CoBhIljPNF7u0OK56mvj71s98wLI5Vo8TTFOO3L5Ga1VcsJWUj
qu9Yozhph4KQ1wadPKKi3m3b8X4sm1fFe0fDCFk9wDMo/xQvG8df46oE9agzLZkF
7EyIDh8zN+6EEOu7VyE3/7/aUPboo9CyWOvrad4N9NAVN+/McJvf8ktl+YsYnR7W
KJztd1UHmZmZogWoNFTETbgFsMkSAKWogX67oRK/GxIlywWAJvBzT5UsOaR1uN6b
2DKjCmi9buaO99Z33BoULHxjoV9+fu30Fk+vTUFLxothMr639XiGCLQzmL5pMSoD
Bn29esL3Nm2LMSfnuVPBk+MipwtFCb5LPuoplaJHDQA6B+CPkT99YrZBrAlknF1x
1QZ2F5DNytfBhi0v70XkkPpyyA9+hsEC6hN2YOWrXMKGRYhAo+WEhe3KnxtZNopv
o34mMU5s3uMbGPXqJAVlZZzRHveMZyiJoq1Qgbs7sfkP8eiqwsLDIlZOpdNkR6fV
GgaSH9i076n/yWlj/1zfmn8nG4f9OzMAM9VIsWMsvLEp7ji+a4WzOL2UwWvUnxiW
8F9AcxOTODW9GnOqOcd5qR/vFjfD1xeG9Xv+Z+A4aPO8x/2x5brTMCAqcDjXsj+K
TwkvOtqbd0nTIX9vj/XBgWe37co8zAQxf2IVBPls/5yMHFfh8a1YSan1ZJRWhALQ
1eGXXxBxppWNkYrm/qsZ85i5zrPx6XUJUgFrVQwOIBNskCR2U0P2SQfDs45R6nxZ
bDMVYT4BXtoDpdwfpjnNlz1E8i2sRGJGg1cwSNYXIfFTlEQX6oipv3bqA5++bDPE
u5naP+1Ioar96U76AgoM9uYG/lwd5Iqps5jrYHNvuub2bvnUpbNslaYo367+SxvI
lYlbJnInirYR8Q95sLHZ5Dp+7sfiFNAiI01cImLl+x5lRPKcK6HHh6xR0y2WYfJv
LNKP1E7+g9nRSgMgznVvYyAX58md3pkq3Ihc+Z0Ku0DP8TGCdZAgzuPgTuzcGt96
PF1ZXnHNBHpcltyjbpVAvCekxDW0ERQ7kXf1kpi8PuT4n9P8UlkDUANicUQh0+zs
yNKvTFde3PlXUKz/goMRtnnCn5Ys5APXdPyD81D8Sf51JzlEwDEuUqUyaj+LkumJ
JLa4xV392LOpFA82FulS1JQPNAhSOlRG1leeBSl6s4R6oAZ6UpxxfCOUI9W5F2fk
A709GxUvMlmPAbmJOCBiEzjrVkUrOCDVNrJZtotzD2yr9000gh9SC/hYAJvQg/1T
KiazX7hWoWIRNXQZZzmibL6WxrqQUJvmZbSAKu4WSggBbNmnQC9nOS3tGgarpkSU
Je899bLH1gCQ3LsOHxYs4zU+NsZgLYD1zk26P07nqi/c9RL7DgpFIiw+rmt32VmA
JfdQzXUQsLdykxq2KKDgd3k05iytiFyXbwHtM+wVTy0VBbNujEfCIHzdiV4vdwv9
0QloXcUTNYWL7qjNZ6VoHsT/Sy2JZaEdi1tVaxKKcIVoXKVfOcuW3WAQL7NyO4EB
m3gOuNfJ+iYTF8HaEarRkEEZpyC4sGGPVMviWianqd2lHJsogfvlJfg1F5HGgAcL
0p4w96N2xdmlL3BKtPoAUVPv0B3edwcoGu/jbazDAK0K6Y9H1BH+hoD8uQxyeKs9
Z3ljem+VlGCeMevcHyihsZGzHH1PNW0Cx4LOsdSZJ5iT/6UzUTWtpKTxkE7op/oV
PwnbpRIY5H6w230IEaU7c8iq93L1MOgcWQsc1za5hZsABkoNyLAWYlpsVHvkbHHG
QENY8hb1BA+X2N7kqdjB3eBZmJhWt58bkXdprz56B+2uZBQKH3tRsG5mxgGjAdEJ
5mqziz2BOFt5nUk8lM9oYMI0vRfAxJQzSjhDbFBJeRhkrkHMQquLyPNnb0iOVOAa
jGgOfNBWWZa62u5FgM3k+qbg1Ze68luBENdnB+iMG/opgTE7ES/fIoPRzNJalnbO
XsFtEWGLZHXbR1UnxylVo68Y3ePEgc7Q70x08h+e1aUkjxgYLfWqz/bGkZFUg6dB
wrliIV4JGn4ejcIxpv87EZvOD9fmtAdOdICf4sYnkocIg7xgQzc1CCu6aHrN/xM7
k/Q0T8f1j0CnyHSrXMw1aAL9PfWSFWL/QVsOMsz/UIyAmaky6wr2v0rsbmOlBk40
1UH8YAxmrfnok9mxgMZK641th0PaUiG30mCPhlhUymx1qhi3Q+pG8t+xLXlQbA+M
qC//om5Jbd/GzLZPSU2MaWYfcQqVb31aTllGEbMf8w6TRinSe1F6pzIHwbFX3WMX
vnzN0E8YVHXPEeiUMyryCfmwT770vzH6Ti7/Vckm+qRXS3cwHiky2A3dwiHXYqBB
dA4aPFrh/OR5oUBMpOzg2oTxDquLJekv+gbgLoSQJHxHdM/imcc09iZvHcFhLnav
2UGTDXSD7rcmaLzYfsPri8gc4edVGyTGh0r3aRoFFLaOTmjsNyZFxDD5hgkHub3H
ivTQWWCI+Dai5Y3W8FZQdC3gZIxep9X9YtOXaFCBRotCjqTijMqXQFyMV3wSs/+K
iev241bybt1lvE6esYZFslo0nypHknlu5Y027t1K9hSff+BgbTOBK6GX5SxTvohw
eAFmBinp5hUpdExu86FzFkAB3bxJYF/5f538O/6WShTFqx+GP5FvhsFe6NUQNXgu
W7MXtdnYKzNDzrOvZFSHfER0PzIhbcR+kTTzt9PrVLtOQxMjWMGBd7Lya0qkKwBQ
XaFs7g9xwrrwhBP21EVbNz1gEQAIlBiRZe2QCue3yJKUIzultFXA/2fTG2Yj8IHy
4S+CYR4JpG8CQFEqsEVPcFNiixjJq9jddgB4ozQ+ZrW6iOn73ti1Yr2w+cj0O85d
WJlZjKxce9cESmtouWicgpUtHLRBFEmTACV5zaX8aNFYiYlQH8E/KZ7A1yM/1Rgx
G1l3KM1zQBQ+ZAJdT6/DSaqtUOFaX91pHDHpBUVDr9DPt4mrRSTnvxiqxqlj9O6i
7RgiiBfsUv9js4nEzwuxkzKnePQf7XBFg/8fcADq2R3ISNpkrcTday729JojBUzg
DrZSRUKIaRmWTouqD2rPCDfwAhDIqzkahziTkaGEBo9ujEmXW4YxKEqu31OvCbyh
0vaejnpvCIwiDyC72tR9U0O8RfORiqwwqvRSg2u2Yu3+EGVzmkjHzNJ0JuOEH2DA
GBLysPtUdH3X6l4GhHU1wi8f/MIxcrhTRkmumvKrD93tlby3x901orCxVcCRTlWM
zgsF9ptTSM/vAU3LqN/BnCWlwjDoHsVPJrWbe20b+9XoB9OU8dWLQbe7pjK8PPK5
oicuhDhMdSM34ByI9x6DZFCZS84ie1/YnqlynYoBhbWBhCrnJdRWRdP2XNpy7TRW
nX1135u4baQM8EBGTh5WoKSwYiOjCEJ1VFB1R4hKLYyX85nT3rr2kC6zrKOjWmn+
0ist8AWGKxC1P66cS+n04iJyMagim3TW7MPAe8ihbw7OGJ0AUIsGUbF/fNKGJJqV
s6oGO9F7baUFjVvzLmCnTT707KSjiC2X1qXXCPNP6VnojZlbFi7mDN8RTtuy/33P
5Kc6c6dCCWkaOim9lwssHn4frRbAUqVnbqoOwJA9B2NHMYOje1uAsr5FPAJ1Jne2
ld9uwQRvgIDm/2dWqgfR3jH9QZAVS2mCUh4zq1Ck1eXxwOr6xXx+F7cnT/8IUixl
bcUS4PLKunDjSbFTMZh/KDthk7QcBU6P7Vs70kWUinRUBg3OOifLlhax3JmQEIU2
mNVW46O345czoGk/CZwy7oNjda8+HoWrRs56gkFc8ux8Yi9si3QUEwLL76tR596Z
n/TU8rKHrGYY5cBgjyEC6yTIjiPppqlYUzP44yux5B1e6+8XQsx70b1W7CZU2Mdg
0+O23WAXa1P3X/wdZWz01bAuDX6gMakdcGqZrcQE+RKIL9DxytUozYwD9y0Fv2E8
nOeVuky6JJdrPinPzTfilVP+7o5E78vvklL3pcAFNhP/gl1uyloAsrVkVsHpqWvO
wBqXeAenXsbQdFDwV9G33H6S5dpHd7Gydesv0Wo5EcQMwELtx9A9I7VuWq5WZnyz
R+R6xcz7ObfSTvorGJDmzW+xk3b3DUGjCLmipsycbg4ITAZ0LtfmpAbl5A6Lf7xj
6+hUoM2+XGLqBPCT0yLjumtJueSAi4a5hj3xYiOEOVMY3w97TgC9Cpey99JL1x5G
5wnYE/iXNgdy+mhj8IFSnQXO4Z8togq6cdmpM4t1b34ca46eG2Fc9Gm63MTc3FIZ
a/0wPjUE178vBSCHFoo+KHUhYJHrH4mr+5mZDPRgp5p+CMJgyPRF2rO4/xJNwdu/
K8na4hdOOZpIZDsD/kdMTg8TwbtTQAQq1LfbptNyHQPSIE3fA9PQ2CdBFftjN8wj
RxtkDgPUKrtm4Ik192QB91wJv+KsrkvPQwvRVa9Qli1kYacqRqcUXdweUeSxwr8U
LSSrOJ8P5wXXi9t8PA7r0MiJDUl0IEs5HVAhPzf0lcQKkcxeAnerIC9Age6DnrjH
KNe4ZgWgnJvS0PiX/Obm6ZItYqZDWb671a331Vc9A2ViUoHfmkUP5EhphSoFVpbJ
RePflrv/uyjNw7H9IXk0soUaa826fxMuz7DxPev+DvnueuFX5+nivaZH6uPA85f/
7UCU1QaJ2JykxVC8BVDljHrlNpQAY6P1jvpFrCSkrp4pL30DAa45NSx/rISYVSrA
CJr8yI/rdYq9SnbqNnr7Jxlg+gW1AI/HkQI8pQREy31PAJzSp/BDMguHfpKkJHWE
TTwcVNn0zbYdHsKpnwkVKb2MC7Ckit8m9E72Wow5d4az6wkBAI/klSw1jTeCUUz+
CcT2JB+j8A2kOZSgrAIjZ8Wuo3Cymr+nsGLigBaLHHFSddbT0J2swLlNY38F4mFK
WSOghofVpYum5rPTXqWzSvAL7EvLyrRWczn/ifJ6qbmUKcVQove+SUqrzMveQpCt
bsWHs2KGGfKmDqAjXjM35hO1y31xQKcsxagXfjRCwbeHTnIVJF2Lmy4bhx7FbAWA
7T3dYpsYxwSV5RnSxs0i90pcjl28Cihjf+tdBHjJ7Zbrj1FoK72dLpX8hXX+9ytq
+bYq9M5SKfsta05M6Ox43s2DY9b5pVyA+RPo/Ma+5o+54NUb4PUHIBnu7bGEajWO
C40qxWqfHf8m26DX3fDQV/Br+hlsMsZ2Dk15szeUqdzdEa02qp7kBIDqaqJG8CF9
98leIVYtyeW4YYEs6mur4Vbka1fUArng3+g7AmKGCsesHLYtcCUZOlEFmNHLzeUq
lzaM1yfJf55r64PDYPoCH1SYvCFWsDwCOS/RdML5Sc0A5VjMdFwb8hwREobMMwoG
MC7Qonw0leH+Bx2deUWIB39qLR8zfRrKMwdR0Ep/LzmMEojOsEao5iAjNYHvW271
Z7Y/J4SfHKOQMVPJ78Wsnop1SCs9lcpauwvREBFW9DW8ksIVpncCZ8VQ3OnWCAAC
d9aEqHK8Cs+WvB2fQZGWT74tLYCYmmJ6T4VxetIC8EPdlNJCl11Ey8+L1XvCgKGA
RkrFibxpdi4dLf1WwV2HASdhhpvpvPBmhDhz3W3lCIMJUOG4qB3tHgcDJATsY6uh
nO9nNNA6ifPhVj0Fa6/I2+VNrPhQAY2pGStzI0yd5WBAGKYrlMfO1siL99R6nnGy
F4r3Fxm/Exp/pQZXFmI5Mmki09D3MyHeUhMFBYcJY/9mbhYm084gcgA3lBUesvmn
VKAM+8CXkQaAOA2u3CCC37m5hbzQ6cvxEGMc8NynnkAdaAok3FTk/ISgFuIcU2zu
cDvYW0RghyvYMFVLKrTehibC54KopybHAcUR4qhILgBIzBEgbMuGeJc3I00nujE6
yWSJId8jMW7iNW8q09B8MN8REde6jQDvkgEAJEEXYPfGQ70xVjbxTbMdH7BWX4Mv
gKeJ0CBhmXE76HQlHSfqt10kAIrwLv6p/KEPbKB367AcrRv5gC4RYV2+xvGk11M8
sCuZLXGdk7ly/X4Wra94vnRmZEd1JzWSSj1wsHE/MoTULK0ecKA3PyJZIyNXanJG
8EjkgvaNBdAGycUCIdA5r2nU2gaypmcDpOgi6oee+t55xuupoTrP2OrxjuLnjg+e
SlLAr/GiInGvbQf+VOW4U+ZExdwgVysjYzKZnPV5/As0KNZVCdaS15XF4hPyda+0
Yq3Zk9jyv4k/74VDlSfNCj51c+RLGo0uCCpfs6wm+DRgXWGwWjuSq/Gx5L3AruiR
LtsMgjSvY0mZozCdgYeT5PxusVLCvFtzTaccWa5WRUm/1KmUaPLSPCMJ14ohoSrs
/cWXUUSuPCYuse1NRfBgvA9G0M8uUL0FLaep+og5cw0oCxtGUSCu9cWMAwipGEBK
/Xj72ZtYQsyOqg1PyeHj/v7t1ETHYcz/Q5ZGo0koUDvKwr3uPfWcgq3V84Avy5PO
obRySKNEi7P4THDuiU6+t96jsBXF5PLY6bQEp4ZbH4ajh7azLF0If7hDyAjRQ0SY
o4QBreP5Tf0BEQRsC07WS7MnxOyY3KortNcnbG5JojKvbZuMkS049oQrENi0IWvU
qN0FkVpc61xz/d18+tq2Hj9WUFSb8B80pRRH7g1PseOX6hCqzFyqEFuWsHCh09CY
TLhYZo1USK69DTAAVOSB02RiLai7EKHeDLDkduLUuiRQzwSNHz93Uv87HGIoLIt+
z6Y9//E8G+7B3V4J3bpBJBNFWU79RNejvAv2AP/wYDyh+kB5gz45myaGEVHiIJZd
pKn45AaRdfONHTzrDNzXmj4zuMdQ49LodP5BzWNKNjgd24P4pBJxgc6JrvsqGObN
iSAYbD0qs11+s0LpsXTcjIZuh9afm+lF4CI6SP+/ms+e5mL9j73RCN2gA95nNG3H
W+FoU0jL3uigRlMc/no+KWdNksFXkTQ3V3DgUiDMw3tUI2llAKENa/8RB3G2qsMt
kQWVpGEnDarUBhYK+e8VLPOV8rB7L1hLlHSeaDwpzfdvmEP3zRd7Ww59HpdFdpv7
Zrkxcr1MZl9ZLxw0ufYxVlG+z3Mb8eVWM8fWxTO1jo7MTiv9cAYtjBSa9hk3mNL3
VFibCsvHqqRRPjH3z0NZYpFbVE4EA61QBPDtrdc7+xt6mV+H6ce3wZOKtPBDYeTA
H9IsaUUDO60Ix6RYFTIXtQwy+6ByDdaH5If8U7dsvgu90PP79lA4TysyVhQocBRv
ENdZHYSyuKGk0aEqEtsNazjFdLNIBfYPzoI1NUBOXojiRbzOyPXXhMN/t2UDb+so
gjLqRBtmoTQyrldsPPUKD+ABEXuWKeWX4HQE24AkasNaqLGiZdHfpDqbya+GwJqd
iGBsjRozF0cQIl9lyNBgT3yOErjQrYGOwCjPUxFu3EOTcf8TQ5l5Xt/bYCk8RjmO
nMOdXvICaR397wvQ7+z2CykZq6CL9+qUsErsGKjKdmirpVd3z1Le6jOSydX5XJBm
2qDUw2XuuG1L+2RztEADdJNNMAA9MXa08QRjDOOi0MPz8Uah1U+qgCHOgRE0PcWF
KbVKOAp3JA4Xl9Wephlm8ZABcjTgH3OTuqbTSjbjqh++6xsMgmAptJOSAEjBXAXu
AXApwBDQkA+F7+KXua8uqzIaNkCfYCuTvjL4Yr/cl/2KYH0D7e9TS729uTOJ6yeH
r7ckYvuf84jZW27DoSMTdwO2SNvCzi9FvrJt9C6tWF0u0oRvGhK0KfxgvpYLTF4Y
qLdLJZobQCo5A8UkDzPM+TebJE69oCa9PKYSEAzPccneTc781O1EDSpMkoms4LQ+
xmAc/Bh2emKEcpp4rS7Op2QWafInKoPxxU1v+EcSkyu9mv+GC5pnX8EbSypl8ms7
O07S/RNqXRGM/U/NoNGVi2juW0NqVEXmIWuL03tzTbHH47Ig+5hdanAGEY/jqpwO
l9wpShNjPeiKY2JDcmQpppt7r9vrIXpHuXoMz9xSG7FUiQlS9+hHr49kxknrv899
O+BCR4Sviz1Pfgtw2iQAIDg6PE1j/vjwk0+dvtoHRp29VA+X6Trq5UO3QuH+Cdes
A0L4TYiqKPkZAU5Sqq0iMM4uN56VpBKt59hT2I5HZ/0gUSu1GKMdDUM1jHjLxf4y
Y0xe0yDH6giM0gtFVAmfHI42+zolAdGCj0+etvzIop1C2AQVPY7MZ4VtmOAubH8R
SjrVaBLci10gMzx1FJmmAyUAtmXcZ+s5tKA0bIDwRNpu/X4JSCLoUwR5J4//oUzO
ANQqruHxb38JRSjXB/KN1DWeIZpVFG9Of6Cx5YdET6r5y3CcFOsHBRwOS1OKDzK3
IPmEGkZ9WQO/jgoGGFnCAm9JsI11eQWWnU4qovXtZsZXD0MKQ9xl2xZL5UG+TNC7
177d5Hw9usPTFOUqpEBNCaqMEm893XOKgxLkWx9jYR2hu6FCJ0FvrIuFWssJpgEs
9qUzWtRD/XZpzifqHSQhuq+Y79L407PYzdofJTEnc8CuwJ0ihR2S8di6Qno3OUlC
+TSSIEXbfbUD+AcbRxaFclqU7J82wskjg0SQzxal9hMme1fyL/puBvp0yI3yOzUM
FJpKcvt+hGTGfolxsl0b8OOXVYrGKrG6bILt+fMNXHsQ9CAEFln+XJophphholg/
2ZL1vVklRa+519Lw7D/lyVdseWBL6+e37hH42RiF3V8pg6lHK4qkZsL41f/eETI2
Xdt9D5/QVVIVe9F9KT+LLF8iMtHyVTZHtajnkmI2LFMLSC/8OdBPp69TONaAVuRR
GMX/mjOZplIAp55rgA8CPs7SaXwJpf3D74Bi3jVbp0Z2NzSy/3uRxnPvb4O9BDlW
eRqrvuQk9d2ANwUJzqVkRbqZ20zZWXZ6ifaCzwNDn/+hrwon6QrWSruwKvhfXvBj
Y53VKgAjdjhCto77STKKmfKnfWrQHrcJVh5xiQQGFxGGh/MSKW7bV47srSN2UcCs
hhhcDi3yzyqyK2oCWlYiWVYj5AknfyphV5RnhqUboQfNc7s9mE0pH6SVX8MQzBEJ
JYmgkpp6mu6/gaqzwStFPB3sJFptbWHT3aeVdlm+Sbs3r64Put/GAPox9SiTg0r9
vPHorn/IvV4LLzyFv4u/Pnf4EW3p+HPuAzGatXlmLjoZc3pRdpf4iJRazLBg7lGm
TZLdq1WHrR0I/p4dvwqtpVUlAY27ZiRaSbo+Fe8rQsRD2EEdAUWHltlEpWIThr2m
wlhmU4/3SeNOF7RF6D7QRfPyqu3Wuv9Rq+JphZ3BspsrUGNksbBmfGVu3xbJnoFP
ybWOvDbrOk996Xaj+MoUa0s6qYLuggAZsnE6NY98tfYdr3+skh6SkdW7M3IQrKsE
bsur0ULtwjapo/iXYxfOAeYSow84B3yNbq4bzN6ThH2rmQi/sPwHSo4VmPJ3kIFJ
eeuxGfbNmNuAUDS24IISlfQLalUbXhhVTO5emf9zlHoAjtzGXcgshF+fdzKyKm/K
l+wp+QgwS/n0J0FTO8YfKN8iJ+A5nokGGyQNlNekTlZ0XNzGCV0xN8GKFFQat04a
Pkt7/5JVbEqhxjD7fLu4YzkbrIzHn6ksFS3hZLsdLiRxRtrg299zfp4XR5BuOtve
lpJhfAhtYXV4iyXDpNxvachm9vfr3XIIeF5St88he+1Xao/K0Uxzph9rBElfBib8
FWgvEttvHcGopkNYyAk1gzhGm968xUxT/rvycQ2fseAUwFvMJTOAdIbbyoXHYOjW
0yAxpZiEvjYuJ4uotrUHDeHVL7XcheLBkPV2sgGrGWn3xvWMr9Y5WACkPHXZ8nQT
it3urayDPJFChvo34Z9KvbxhxHVQgrcxi6MWrXhIJktu0YvR0uLDhV4OL8YBcyn9
Wn4eJqSf9oF+EBOMHU6xbA5CJk0FweVhLXicoBzVQSMwaMwMwt3uXwAAIMef0vxv
pfGx30geQF/QVtSb5C0eflkr9vsYgbkHmVMreQbqkAnb2PNiCjZkFXfiVPjN59+m
5XLnFi5fwBKDWwY+w7bFR7QT7iPKb1N0IcGkXZmh/RsMJHbANItWo4lZl49PHgUv
4UzHlZGLJu7KHr8KbxDt28m8YjbELmGhS8XV4vElBRnqvA97oAN/U3SzuNtjdW00
O1h+H4ffBRoail2kjimMl+3H/XTNt8rvtghEemmXARo7QNoB6r38ciRdq2dMPLhD
0C87wn3+KCK0IKO4OF+WP1dLssEVQSA4lfDBa093H8BiyoWzZb0I+Aho658MmSC1
7x7W/m3yQzzCfqLs4wBzjVVg7D5Azl0MCv0ncCxEtbfe5ekA7yIPfd8WHVWXPumb
oZDu3l0ZbCG5xc6uxF+9ty8aku2HzH9mXibGeJwgn7NkQ2cOqGBQqolWCtz/pPLa
QF2ORvMqtCwWgA1Em0Cyrv8Pe61hhCgksiSnU4goA2thADO0ASbEC0+BSqObdrSM
R872wMUgNBRMmHlXCWYDbVXtlVYL4HfdQgyCItt2Fgg6Y/euEQiFkWrYoCm7TUBw
9i+pFO7S/6XWsfE5/pW7VUD2Ak871ISPau+lRdrEp5up1aRSZofdg1G8qqWHNasu
UTR9QDe/n9xNpFCIL8yNN1LXo6Agf52lBDdO0MEQhBVOQ1pY3KMQTSqieezo+Oip
m1/cu0/FARtVZYLdyyuA/1zF49ddeRroutkIqVC6egOVwUGaNvAQP0OJH7mNBnng
0AG06t3zsnersSm4v5Hr769T40xOHw5dYhxaahPwbId7ik/hHqD3W5O7YnM/sKO8
SRVW8nn2j1P0zAOs7/GbuVeS1QwW3wvx9df3HumniTosr7O7Qnd4dR2g0QuZH8vp
px8Xara9eKjwiUV1Sk5wAZMMucs92jUAa1G5tqH+Qst+KAf30sdWWiStXeVo3kSS
aIdrf3bhvYSIiM5t8VR3X8EjKRLIfwMl2/oMRsD2FUDE6lV/Hr/rofcHsZuWyP76
D2kYMfWWkZw/Hk+LJvR2bbBKELLb54UPT4pUoa5+eBidditqtzmKpq2rrdKvlw3e
dX+csXhyVby77UD/jf3lpKq0ZXriopO6mmUTU/bNxMsb8amcVHoj0BDldN5ZS++u
Yq8hHv6UaUozACXivdwBnGsrb37SGd2E8Q1S1CW6480Fbp/5ur2VMOAPF5BaktGm
JRRQWo3K8JB1nxEWiCKi007HOzYvwgjXjXHtAXeKTJyrColMHuFU5Hpa6H5gfxCo
Dth6szGOGlB0cQaEoLKb3fW6jDdVlW0qCqq+m3j0xdHheVhhLb/NNFOSZT9WE3x/
8sMBQzEwQKfyGni06uzaw66/M0cscHkzspI2V20v2GHJxTAtXbUYNnyJxrE+y/vY
+qH5OdqsxQM1TVF3/VfURs2HN0xuY6clOtLvESdxZ5QowybBe2fdaqEvK9Ec/y5m
vXiyu7fxZ04J3bFPVnmD4YZMRkXOCDok/OgxopiKIQCvdO+6VS9dshQFdBWQr/u0
b7ypPA/PI/MbPv4FOoIzmhqvXTtuQA+O3W4m8CQtmE/iV4n6MAXKmJgTk/WLExjW
2r89ZcI29vM407JcELcYysi1oI7jr5wzjfIIxoqAEhHg7lcCpD3kgtIKKDQKrwDo
vW8cibuN+YZL1zVJueimBIbiMkTft4VcgVaat3hHQ6uOtg1ZbiPCuMYlhPmTbioY
awoTOKgK/wW9L2FdJRLpCk1aH8OgYTDBLM/JSech+qKzlBsTWVqNIgfyuEh5Cguf
nHqUylyU4XCqDomrNvdn08IrcmvljTEOO90PMakBzRFPvia026yA0bqL7xk9HxPB
p9GKWa0PguPgAdDR2O6ziruGLiUHcsWnzCLIWWmqzNOITy1kM7JHlauiqk3lu/Dr
hVcg6E9d9yN3tchT7M+8DqQTMdJ7PdImjpO66RGFMNTLvawZdbCiSuZf4Pwxdper
hyVYPJl1RbiG7MKVEx6J/9LvXr3gBbmyQs7UdjZHsDms0/d9rGIzxyb55u9jEXbj
w0/UW9JfewFs18CgygAHSEWlqpZEPTg7L3iF/tj033pSy15Wy4ahQTUePj18z7Lb
1CQGkFQqTAqcNP63l8Q9qDviBkHF9FHThQjJsFjKZFPFSn0PL8rRVsq5jTEumRf/
AFwNgpbTuvl6g+oOGg6+P2z06c3AEanpA6hsewuTBfVDk5HIJchXw9p4FYZ+mo+2
nMm+TKbAwC9TVZkpVlXHllqff1FkOhzG9xN+ho69ozbZj/12g8RyWZ//rifPJ++7
ISkWU+ibspTAy21xdU2z98HDPccY03Ro0LFQS0vLleuzwmEJTLLVkEked4RJnQ14
JHjxLaU7ACmQjahoqnC8avWocNeLT4MH3T35944qC0A+3Ii39Kc1MSSfUWjWr+T8
7AokBXnASzLYEmwsfVOL4xB20TQ4kuycCFHOuVg+rt0SQLmTYp6HxZ3DegxHc25b
KRgLLMukPrp0Wt5vGNvlcDlBp64Gl6NT7VKFfOnAgSaS4CVxO4jFtAWvIoEBSAN3
ZDjvNUljmK7VD/zBUZQwT7F4uFcFuK4ZGwn3ai6aZUwNm7b7sfQme+DSko+/GznY
KifJcRUj+IZ1MmE4/qSmnJNeQ8BfhV8u5JV6AmDG/89mOo5Bi7NrZzQdzBQFBnGT
oRVmZN0d0Pqq8MYxrCfhtuHgTD1W/fDA4Oq/0ToK36I4rBRbeD5rW8/OdDMCSKBB
l5w68oQrRixdi84WpOna3Xq8VTOM7uHk6IXCqj4Mw6YHje6e/LEkFNOcVcqHPamn
RhnF6aURbhFa3dLeuHyZL0HGHJyuGRC6VNuJb23qlTbsRdAAwa2pW1ITWDgSeSFt
JpJSrwcUPuONroiW8v2Tn4e1XE6k1L+WMESReBf/FowaMPpDPUr20lOs7rKXeHiJ
X2/MapZvoIx2Y9PnZ42Sqkkn3LKa7aqeXbCWcBsvK8Lc1/xCrEoYEeR3SWvt3Cbd
oXvIqNJjup5fcM6JaHIWEll5WgyAougIh0C434vI6vza1ibjvL9yPZJyLZ8GBAPJ
dcRbxBFkMZCBAUUuKH2Ro1E6mtWpfTvHUNZ4yzm6HS3t8Ux9IX5XesNnHJokoCZb
TuqVQ1YwEbjmFMo4FBwo9K/AsS6tcPeleEsT5pOUdePUo2MU11QGrVx0ikJmMwjh
T/haUyKynXq6U/KK8fzCj56mFRFAHZbeSQrn3LB0EC4MoKM+d0LOHJ/hEd4svsbC
3VLGTORXYObPVA/Yyc0TQg+kL5wrLb6JyrX94g6yTA6LcjWJcUkzdK0xC4Z9zaZn
ELetq4WtOYTXdnppgI44MRjMTVNW+5n4zIfn+pSqLVpaRlXiNyGf9hBl5CeKgITC
Kp5pOONctdCSWNvEKOgKwyckhisK6tC05ZbjkiOZVvX93pJx6KpqtK4zj3bl6dAZ
ma7AXmljJIJBiBEdbgHvbOUt9B0HSQGnYlY7gUga8NyjBFtgtZu8n4Ra5nFdAYn0
nkDMvo/d3BNa1er+JNsfntsFNau6Aiej2u8qKRaT3Gxw0NUwSvSJxt74ax92g64V
X2dhDe3Uqzy+ZrmdNPy70R1ZToLIYj1uNJAvIxTlY5A8gcR2LfFgpdjXX7mZ9T5f
p+h9sFvBnpRIZ5LM8S9M8/IaaCaue/iZuV4BU/Mms+cJLYSrWE28XmTj2qp8Eis3
eBjYavn5nGKWDtBquRL8Xb4aBTwOGygpI7xYTfI3/faHPc7/hAuCMlIg1kjoll8G
f98MiPQ4+zBaDmb2maHNzbVor0ceb8W+0ZjSWPcgmpKNURxgj53yTh4uNNCoOj4D
WYNL7YaooHZL1twnKcZyKs1UqQ3ZsWRBriYayTuPkwyHXOucPIxfKz5YTQxLYlsc
3fybujrKYUu8dRlRc91FURgbXNGp0PSKy1ccY32H3BNVkzfDYmBNmAt4lIgW/vYO
RInSyMKCrwvfZbYu58ZTjVkQYXenH0M0Q5TJcF5anWPj2fu8A7u4hM8yWSU7Dd3y
zShYvQuStaoM05a6CH1uXzsOMTCGr+rDhiM+PyEV35/u1eGb91gqigw5AP5ACeFq
ZIO6Gnj1T6eLSFOP2cIO3DYCtdLknvIyA5mw0/WPohnDVYddXwwlfgqOwGygTDU5
jwU8oLlqqjIQMh7H3G3YRZKcvETDGbTcAhuFKl/Ji7PNAPpdqgLsNGmrY0JAK4Hq
U86rnh2uDLZzZiIuiH1OmZlXj+kNMm6spHKbQe0+rhqvAub1TKOMidiqEh3gPQtT
uJ2dwaPaIg0bnaBQOKfjz8Xnzpoud/i4pORXoejgOCH082AGjQv3Ruisa+wreMkl
2Mmi8zfEKaTGDzemHDDE4kbvVKWdinJP1GLha+OlEFM=
`pragma protect end_protected
