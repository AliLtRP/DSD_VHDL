// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:43 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
F6wY/vjuliG5SEnk395DLA2nZvyfHA3WOrZFc1nMQCdw2xU8d1m4+EvRDlAEPhx5
PO0EeXacdEkAM8zbl7hG/TrPS5pKDibHXJSgyOEb27xDRcTlqPEzbfJ35O6VI+md
InIhRStvJCavNJ/QfNKR9YIXZeLxfO/ZhDeZDzMVxGo=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 4720)
qMzF8jNarATtissjx73n1553vVY/np31W5Tklbv0HmvNtErnI6Ck0fUJLCy3Mb0p
ziyveRJgcdBbJvG36oa4uat+zJLYK7bGxU6grljinWNr6J0Kqypg2lSJPpZ9VENs
6U2PiVgpcbHBXONovCk59SnSIvPFKyBVsMxbPXfOEovC4TQ54Z4VYsvHPDz9Zb8w
z6Jk6gc3mQJpx0Ra1b2gn1cIVviOKFIB34bheGJ2y5sywnwkav29km7/QHoBMA6Q
ZcOqQ5jpw/GSc7uFcinP5EFaufsLR3LWUe/nlfjQLDwksOdEfyeCKZOshfII3Osn
Db9oPayRVZKgCbzcsfGYLIvSpY4hMFQm58hAJj7YYdAafhJHTfg/ceMGG1uQzJXj
lLLBtiKE7VhZVyUzjHf7bdLnXppOg5hbOD+NinLHxeJTHPVwzSvK0PDabXhj2Q3w
ZZqc46BRMqpIZ9qi4lIG1BnzsZcU9wv3R4YHE4HNTCaKXqAK2xsTVndVGXwQt7O9
y8V7oFirflyPi2c2nF0zY5CvULcurac8uk8FmAGF2azKYTsxXR7fMtpUefxc7GWl
TCDxTlpiN8tj0H4So+3dV+S018JpGeAJOtayLQVQ1Mc/p3s5KrFepV0gmUZooNxr
qKKY1hNuXPnTXFJzshHdLW1R97NH87vdsivgdQ5yIa3Oc0VLy09JHNO9vAxMF+op
o8TwSJKQlx6FppZM6PMP4wYXW3WMSZuV+P/14ETglYAvtqINWmI6/GDYzQrkS9oc
1qRu7KTswcxrfxJ6V2W9aB1qGQhRR4ji9hfumIPDir45iirAnBoZBixWRmyubTEi
ONUTK2gIZd9ksxHUcidkKq6EExNbI49EkHq65V+NvRJxtT4inTTXkfyJ1O5DretZ
zfz1m2p92irNyNuuUXQ+sB66U7utnGlT+XXo3nkQhrE+jgWNa1yA7Mp4rfGeuiGQ
dlDUntQbsaQSiv6kKveHQ4F1ZSoKmYjdycpkvIoYdHhcZBjT0Z9bx70UpnTjdGAG
22Ev4oCJxBr4Y1W4G9u8Qwstozbd/ieqZLOUiRDwXp4xLwm5qi5INFbotlpf+vIA
0fe448zyK+O7rsDTx+ZyehqU/CW4aKbK9HlUF29M0SmSbBzF2saXH70V1hKdp40Y
flAds2dA6XOik1mj85YFL9yph8yrMNi8X7hSKoEarHrHU1oW9rGs0WqAP2+HlSU6
CoMOK+Kb4oBgC3IN25qzzVge2jf2wYpH+FfRNc733U3rJ4kgjEyn9eIM0jgS2/D7
rVF1yWyMDjMT0lIjC5N1NAgCjJBtHI8N4GFsulzWp1AG2wVxBgf2zm//sEDoaUPX
cF3xhi0lO5U6EOhVF+palXWH5fs8rRFIssBN9ScE5j3/6xnR6CfEVEfuIQv+eJ5P
hcyCf05TqMjLYkL5k6SXHUmoXqSh+iM5gvoqPBksoPrsm31zgSGNrtIlmF5Vqf+V
oaggDa+eH8sI8RycrpbTbPz3dnqpjraTjG8XlAw8MPxT91RIxePNknuiG9W+3KgK
fGKlYaZZtI7Wi0dkYGN7gB0nMtFt5pPRVvJ1HFa8m60ucu1WEv9rjaQyPQBhE3ZK
ocL5nWRGmrL7LwfbhZb93fZs0UtQewJSj1wkI569eCcX9EBxv7OYl2hFs4YoU/lY
uRvunqcP/HKgjXEfhEcOiSUhoo4dT7KA3Dfm2xq6ViJGmRlA76yISz9ZomoRgbWf
WAIqpPuDgPq972gLS/AoSWO6v+TnIT6tBSTszB2O0wr14vDMp/HHzObjaZt1fZYu
ecGaVaTK6cX2Fp1OyuA7THJ0c0p3OoPQ4zpUe7m1l/+G/OX65r/y1I2tGk8CMMiG
kmBuJy0VTP/TbYfA9P452LRHHDgPFae+TTS1aTg4W6vjKyHtVkr7pAVeoAwS1K4q
n6WgCVn8iVmai0TZInjMpRDvxcrjRDsEFd1jADAvQ2tkg258Uh2NoVcF4ZAYTARU
GrKgrfYTdtbdMp3GdZzrm60fd18gE4YpkVuH7OCNk+c6GgkTQCs+G7LFUmBHrP2W
qTeuHPfByfIvhU+t5619VponChR8SrtX9WkUvul0oyRDoBfbeXuEqnaAgQpYlyqb
+F6s0fQpOeABUnZsIrwieNZNPfT4AFtt7pv9D2Z1SeiroydSf5BoGqqXAbpwjY2w
VXCM4AdFzodL2M5qHX07q3QW2jPGK8jl3EixkW5YEh+pjhR1k1FYDQu/iSayvLqG
QlNC5u9ONRDnwCZ8nORYK5bLEyCXHKOf77cHreZH4xUcvijL/0h9HD/CEn4UkmwU
ghUtF5Y2I1tNtsugwrx/T5PMgqfNDfdDm/qdc4pbcjBEbF/UkW0Fs7nANmyvVDSP
SRb07accdeY0y9eMK9hIg3yxkcG3a50kCxoVB14oL8M/NMj+TavSe/RztRcPj6C5
zvlAp+34h1jWeEs23DUZuw5wwxil6d8hAaOFtE7gKbAf+y76nUrzjyDqxKYs39eM
liK0WtFD0D6FK+BUfYeNvREjbijuIPyo5xvN0XLLoDvxyKO4smVmn2vElotcUpB8
esS8obRv7zFKemDIxVcoRVOdXCUsjTGz7p315mxmRkYuQtuFnx8F8N8hRiCR+oBS
W5qRm+Egp1wF2GqVyCWyksiFNuJn+RpdT5M0RJ7LkOxxc9actdfLRBiMfBWD94Kv
2apbSKLYerbCywGEO6iwyHI91O7DrOQNTwmmaCyBJGCMyHKh5qqThCC5s6/rdsEf
crZECr5XCDeqNJjr9T+S2hbpY/AtAnuXx3ZKq3g7DlxIG/S9WKM6F4Tb4CC91wIi
TFMMU7CEkm1yOyBwyMBJ5DpptDOv6mGiIinR7TdjB6yKwcbM2TlR41HCHEPb3oZJ
QAs7CHuAE2dMciTgYAE5Ch/LJkfWYgoy7XOTUEBDgO87VUxNUWcZQfLrgerP/nbj
h4vc2EPEe6EholgdcgwPAclJV8zOMMCMlApI+dCCLai6hf4ftiWRyaFSxwrBdrNh
AVsOzotZKs+y8uFrvUYCJmR7IGoofcszI7vXkb0kjYjeGo86ImEnqbibUetB2lCq
eaK3lP3uvmLSkbyKBC4Xzt56RD/DJN/cKWlkG+vRJG3D5Kesckn4IQbaBl3SN68E
Q1t2wCJUezZKD4jlrbW/cAIBIC14qgKwIXxU7F9ta6uQzPGihkp7I+CID5RPgKO5
oBQOjxRSObTG4TzyBSlt0WEr44QrnpcIwEsNqMHLSLh5KimLOFMX2WbbphX5rtAq
9gyRTp8oBIovDKX+bemqmsaz2Uvwsnch414BgDJEo0UxdAKEN/Fusm4pvfKDDbpN
ER391EhnHsGoNrwLIVMoTWKd6Ido3z3WWRYpd14ZpLOwItI94Z8pjowjWo0u7RtU
pcoxnUcdaOwOga6y1FKoJghBCMmCILaiGE38Q/VriYoIx8+h4mDNLsm71puD3wS2
Zz8t6Gfov2n+d+MDDeO8tILuoDlP7dVCb1FK+1019ASqZ4r4vD7NHyCAOdB5ZPJ6
gZ/Aio8s4xmTsMJQFRoxbx74E0FpQBz7t7goj4Ie3HB8N8BRQMEQ0ZmZjYZOl0Uy
tDK30rUB3FgDu3p5pJUDvjLjDFrTcBTme6kaVw6raayA8pdLyb0U2yPeiBewoXMG
Eey1jnVoU4VLlgxEVsXk1HCn24Bal9tQUSWCdlA18bcqqKW+9go+oPyah81mUBgF
ko6WzRLMmE4KXVgW8l0QTLj29WPGDK2Fsi1qiAVvB6B0H9+3gdLyJ5K6Aq32Wsoa
rN2zzbkV/7zZsPvvd15rDlmUBq/nOqoA+xqnCws6FKeew0P4mpLTFol38WyFC2zw
iwAQWQXTFc+vkUN8zegRRPrRZMXoRbisblBDXzNBaRQtlFRypsSrsSryCB0GLhDB
3HlIX+NeMneyhQaNTX8SVA4FiRquPfy8Il63kQNl7YM438YkcWtS9DsbWvT2iQEx
cnlb17Ctng7FVhNSBamPaMyNLbkI3sbDaoFZUPGgqbgax8V4LCXz6YxL4mHD8qj4
rdMrJN4TCE7Vj3bsKfUH4EbU+fAzSkPGIwTtyc5Wguo2MHcNEKpsDrMdUdG9bEtO
b+FZlpGsdizcwuFjL1G2iC5IN47cXDLFywMDpKR9tKBOXexkOwCPXmq3zvraceVl
KnFDblQPrc6p097a+uVnEgF8GeZzVxhADFx2X+G+Fr8iku8sJGTip/gSEehqN2gf
vTmJ4eEGQNeAWs20ck9e4QhNf/nVZq6nCA2fD7Mmq76fzrbPAY8hIy0b754xBoWZ
H3dNvEYLvDCG4j3idX1LCNLrkjCM9ziEVf8qnonWZSu4UahArTRiSuJekaEL4xZI
peGGaj6g3jApIH+oJf1BokhCyt1eG7jOKoPGuctbxJ0UnL7Kpz89ZmLVUMek1z20
8iJSpA9EQbvghDwPQX3er/aMpdViBUQHy6GS21XUp8oKVT6d+ZvVXBHrVhEetbvg
fp1U3oOXPbdFtwF7Gjges5DZw2ykYl/BdgWvQ/dRlmAMi8C+eLYjJ+PkWgjKEuxE
tDy9p3ARHEwzO8Y9M/X78pqKI1bYRl0SSiCmVjR1aKpd/lEoBxouOfYOh8/g1RoK
iH9TIt/KBOnm2Bm52YTrJ8f1jWqfAzbSeueZj0weoGtrCpGHBhQ9QSPBG+gwZYnS
mRu3lei4zXpvWAvSSmg8KtuCIO3SNBo6HZXpDT1ZW2PfUgFxQa3ezbJpdAmSJm5l
DoxevSffxRzSlXw9XwjNcdRgtVIoeYBgH2P0rZ7OIDTiWqUZdJxjH8oVfSqJIuIn
e+7pE1lgBLQF/HeYo1MO8O+DoOFA4aW+U3dsNt4m9B0Rf7CBWBbjRS8DzrMJzaIx
kfsEP3kM61Fuy1Epl7Jh3oRnlneFSERdEJlGAWwYiukxFdyBj2xYtk9FqK0O7prV
C+JcMq02Ktt8hA3pL3nP2fbtX5+HNWkL+8R3RdJjglwnCHCZgfifr5UuPfg7ns1i
wR0jaeeYbJvfXgKTzKrB9PWdRFyWlxgtvn1ZfC+kdmlr9q6d0et3bx2qB7d+rwrE
ajtP+MFu05PofRNgQFNz+HEDtVeVAq4EHY5W9gjskoP4pyMpiXZXUgBgN1KqJ7Mz
WoQx9o2CO5lrUurlSJeWt+lVOJ9/7/KdOSNlH7cmbpHgLQGO2lzofx8V+CV5OB8V
c42RQ7fW3D7j21BaDQNk1mDsar98I5CyQHeYVn1zyiKw8ojlww1rCzg8sEufa3cF
/BBnOtF4B1+roXif6MqKc/yqFqAtbcu8oBp9MW6ZiDstSUf6xV453In7Qas+XKW0
UP0gV1R3aQSYLJP6AeHjH+O0yZDdtTbxXQrlUDf+iMsjF/m7ZDPwMb/MjyA61Bqv
ZAwSFM94B+mFgCBV3KNpplGJ6IyJ64WLbEOQrAp2yZ52hdFY8CpqNFOfZWV5BBYR
gtKAH3qiMp6HF0nfWz7L0r2Jvct4S8wOfRkbi7sSRX7yGRzo0q5pJdVWTH7MiLPK
dmuYbys910Rz7zTUd7Q2IwoUXPxteY0fJ+UrAUYsrva7GTFpJsaiNkD+77VPnD9s
4Cun/ZoMGBKB6rlaHe3ohXI2vLGIbjYe1q+6W6gEf0CHlWv2CT4prOnVekOX0GJb
LrHbj+Qmdh+EZc1RsnjO95FBGuzhivPr29XOrUixEfhjHd7O+BOWZkCkgiIBq6qx
scgj3yqPt1nltMfEqZXQ9gG1OVS5J4MbKsIS8AZYKR24DuZrfmpPZSLVnbmnd48R
fBCOyfo4o1/BiEu4D2Fwaja64l69FRhfVWCIe1tczg7USF5RGa/5s7/EF1fkeCol
wc/e1Eb23YYJ2VSvJRCi4Qu0i6PQ8XUdh8Um7WY2OhP7WMbR0JQ156ZSwTJm3XIr
4aAUio++dKWA532nBtVssZB2Mvs6Mz19PaBhR/eBaHVxMF8ESEJncBiyX7MguZEV
R1tCJcYOM5tittSBGKq6TeJqRNMNBxZNvpzSykU2PD5mG5vRz1ohMyIoFfCjFqPe
k6Nm6tPfli8Z9tfwBM5+MOzmm4R7tOiUhHrqrID/Y96OAqbd5H9Wp9FhDFGLK7GF
cty6bHcHNgw5wrUpmhBEc53Cu3YSEp3Bm0eFWV1h3eSOp8rcj63tkgPD3Pg5WtWm
fF30VqlkCGW1UZ3hrlG1qWD0q+x8aa6VcQWzVIONRtbWSgrT3u/b/PL1M+TKQPru
TYWvgMoso0k8BUWSnwJJdjZMz+iESjCx17O/tpN0YU/EVXwiZPvRVo80OOPka3K2
f9XeY5F3Tm85+8XK9GKCRA==
`pragma protect end_protected
