// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
h+x24geRF7jGLY0X1ucM5Zsbo8qc0CFSY/wm3sNo5tGdZGpHYfvv/FG8OKoAghKm3c6pldT/V/Ia
h1XWeFb4HjNrttunGxzyQcBOiYHpZ0u3L3b6MEQXURP7QkZUcbdFzuUTG/CbAcjCwp9g9FGfuJpL
tu5xTmWTzSf0KECxFaR/9JQT7hlnQwU/KJmWmuaDS17UyHCCaRdjgKME6zKH2PnctxrS5k+pIQgU
S0yRFW64c9ScqybFGcf/TWAKG9PlfcBuFvUTlUypiHnzIzenv+fbgQVnbcchQ3iZ/3g85/cRxjAJ
TtWbVlIA7rvfBbX4Mjwdcc36KdfAQd5GsVbmgQ==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
xvuY8V8mTGUgP+bZuZvPTvyt3B8T5iCTHMo+sWm3DHqRqX8Zd7GmXL50QYg9XGPhEpGjHcS0jRsS
PMlWrQhz2LVjMWQ1ijC76gehzDNjDRj5f/UjXg16/AMXTNedmFRlhekzRf7denHqeGBOyLCDieO8
qa4wxRi9j1hiX9MMSFGQf17TwYltQc8sp8dde/+enkH7W2stEIGVfJxsLBo7HdHYVgXpc1TsG7PX
CFXpsYhMDmqz33+372T7vzR/nhheNSzUW581Pk7Jd+UJQ5hj1RodvTiQH4GqZasxDmOwL3uV0Cld
0lo/ewdyQPeCFdOSglq51t6RTx1GqwaaOujtcIDCm/msXHkkCvWM9LnRz8YD8oT4vr9x5o7Pq9/q
U3M8kcPdIY6NiDzu3geLVDH/zbFF9sqdGJbw7HgHq8cgKbwSTz+/S5j9cgZOsXCmBy3OTtiJzEKU
UkZO5EVot7NP+QI4iaajrOEkKGp7oHfbn0+6+lf8UiwtYq8aFu3t8dBJAN+WRpKQwva/aqt5zPOZ
SRXb2Va2ZpjhUhpdC6wri1DZ7knbu8DwC/t9FfljVvr2v9kuChH/hoNxzVt9EBm4WF8Whtef06Y6
T2mX/JPdv3mpoDnq21qcIS2cTaLhVuP0ZFR+L8du4FpVDWB4OvyL4v8411AsAMcxzw4zu3WylHpo
9QnFi51LHN+s2qlQ/BABopuWQGTlwNZSQ9lMS2mKn2g0Vh/zhUDla8ZCd45fAT6lJh0gyT2Poecj
A2TAXa5vmf5VZZRIjPh8yFld0sRml/MONwpo6EctoLmXPB0rZQ2QmQA7b3V1VIYfYMwYSz92jBnU
qzMNKzgyUeemuwvP8MXs1olbLwGOUSBNO0m5pWPD1Feio0wYhWptp6J9bakAm9iq/hp6hn7x1vLS
1j1X16gJiFNdvTZW6JyQmwtBSKtvNjoJhrvCFk8fIwieoZrk7cGwR81XEyhU9P2cmmhg5jr+yhWG
Ji8nnCGOPyxczG0Dzoc9FUvqxOhx1nalX+nw3FmrvHo+hNhtbdC2XTEenczOVgBYtQnxqz/6/MLk
39gWLZXaWmNLjSA5bAgWNC8gFIHuHduvv6zEp6Lud+PCUoHjgjBKnD2RJXEvlvDx+6mBXnxv6Z+k
ISzjZTwdXhWaO+a8V6Ke85g1eT6obEQ7H0x2UqgFvCYlbxHMoDOrh4nX0JUtx7mH7lJO4T5kMNNk
WshdryjmR3BIa0K+NPaHVY4ygXQl8BH2iAgkz8VUllgbGGruz0jwmbfaUd7hbnr/4of9GdgW7pAy
zjk0AjHEM1yCMA3/B+9TkkmHHYdbt+53heZoQcZfGwADppCAdRODd/2E0I458JYybdtGkho/8sGU
iQTiEcOglrLflbEoUlzfHcvn/+yAluXnzDqL9DZeE4t5doJRFpNiO4YJxjticyt9560XhuhAw8po
85nMcIlrqLWzN7WB1IDP8SOogd7lm/2gUkiFpytJ7/uO4ahxV+7g0vsdDNhAmJ/d+bvUv/kdMjf3
CWgc83/Sa1dgLXmqdUTLLLMlpXj4EeJeFA08aWEwJfQtdFkG9FbXOfxkT4I3YQNjuFogfr06fQ9K
vvAr2CoPKtSUZT6S9/j9jRd6lpWYJkDMP4pILEQ6XxvjIcyb6N4RGIbv4BJyBtJf91yU+TIWU9Pg
Tzq2OvfSuSGTokg5rd4JWeiSgA1HmV9q7MYhg4ymddPY2bw6ZlxlhBJ1JQrJrmYc01n+WN3Adgho
jzkYHA5BCXYKD+5BPZYLTQzis/T80lOPbN3dhl0oTUPYaacwGVu3DItYz9QXp4KQ2/npAScPekON
bd8Ot0EPFoj47h9Ok+Lb/2g0KGdrPNuz4aFGcS85zKZqE8LqHWDXbe9OX5JIY/zC04qdtShGItpi
dHeFZ0tIbYov2mdy0SC8yTOpziHo0ZRyipPI20zdfHjFACa2Ic/R39z9ae7yEhBJnShXZAtdpfOI
RX0n73wcc6y96pKeWt8YdfNrmZUX2FgAx4oyH/bU5BWjLioCamlTyDpLWL2pLfID/VQq5gQ+a+v9
qDhwoUIVJ1LKIb09hLqUsY6PBr+2MxKsKxvNCk0Sg46G1W7Nu9+TwkkHnGUUcvJeKbYaDls37lsF
Qu+JL3X7/Zx6LnGm5cchYrrR8kPXa4uOHuzbq7l0dMg7wI/fvevETYaDPQ6dCDld2V8KF7UVeklT
nclnt/DkmolboGyVeOdIrw/T4XkHRqZLVOFr9KxwwSnV0S7o9QE4uJIn9bVKoSKyBu1sPUdfidZZ
/AeDecaOlGO2Y5uqBumfhPb4UHKg22FmGEPLBbv1vubNASiWbfJW+7eKjRdDa0XNl98795KhUm6g
YVtfqaGzBs/7E3jzrh0wChPGZ4yU7O0hB7mRVHwZVPdA6iBwf1Ao3LT3ve/mfE+sKRDnZAHK271u
Ya+j/mqWAWGcN8WNCt80LilSPeW0sh64bNTrqqUS+JFK92gWBHCloBB423FJwVg2mRNKBCpK4vU+
sUDbYF1RNLZI7F79vc+QJe5dDbokSA/mMoDy4iUNIYQg30I3OGJxlsHY9wgo603lgV5tgpFdlwil
m9NZgXJRy4diYC4IIlL0nNUqPid7ZoKRYTLuSCLURVtRagKwzzSi6L1gqyvednsczfYufunVErNV
Dy+sAMNbgC6QVlLbwKdYkZXFqeLUFdWM+5b79GrUi78LSLGHOs/s+COneynGsOJ0zHRL9b9kTVvn
a9pd8+reAwuGdcVVHt/5NNiXseEsEAtDII+BsP9nZ6Kvhab1BiUaJR1zY4zm0JIz7R4OtU26HGGW
CsxC/dtBzCbi5G43vbKMnN5Ax95G82NoJNuqod/y/xPkSVfausD9y6MudyRbxO1Qz8YNYT8WMR3W
eEI8CM6TzwXE2tcOyqcfiC+n1/ni1i78qQUnTW6xtcr/wgPRXNb4ztOklO24PA319JwRuMy4xLWC
4jNxihUU8eFyEsY/OOc22prKNaTnCyJcUzFGos/HWRNGea5vjPFMHWeHiRCK2ESWT7YlTF97BkIB
fJUeBNr2QtsogWfqkjFy1tLWstHPXdmKvk8Hv4Ax9chKesIgHBhlSdrlEMHh2LWuC8XZKDb9GIES
txKICpAg4bL6f4Vlzi22/ROIX02ry4IV09jCFW04Z5JyU5RWrH4B5iuHj2SNw6BenTuqj5sMvdS0
HS1J6erYKXnNbWUJo8z6dm7wOatsWrMlkO/WuBznnXZVConUuxVidUvWyKcLf2Xj4iuXkgAYsiGT
rvvTUTlK9lJXpgrwGjpK0WWX4X8qxz4iNoaTFieqeBV6mHBLWx4LV8RdRZIQifKUx2jT8yjfIfvj
sGqi7tgWwDnHSmcpWjUFBml+Oic/wHy2s7EjhOjJHoJQ2a/fabNvbBVHmD/ANv1TxPtHEcmMjPZ5
MXup0n9/DeBMeIZFoC8z66/dq0nYoyegQA98ayYxXTfuYAzabEtq/SzbyvSKO1VNbzBysSr2A/wm
VQlYfURh6sy9tKAbLDlhB44o4mwh683vJOwgJ+Q8vrVGZUzr6tYEP49YVEN0vkEzGTSBEDV7HqD9
3u14lThOPHusU/+X7PwMYuoAb2GEzEfifBveif0waIiys3N4uFHy8FfF7Sg+Li7tjlEVh22xGTbB
qxE9wdsvgC/eO9NL8TShpKaMEzQ/Nz/8JGNwL9Cd99UU/xv8rBmT6ldSZVpcAMOPIHbwBf2PiijQ
kuj4iGmW/1EdHKTKZT7Sn9n6BZQmFrM+ihUFCQ6t5/ZNAnOcI5i6V5fZ+hOlzrqUA6Vx6xB7/H2J
94+HfEx//SQaar8ZWAj3pF0OXxPlVFZsdJX385YrKK0J1qCOjewrexR7hY6QHWOLJSeSztwA2wR9
fCUUbIdgM9TG5IvpxANs9+7TY2uBZ19++QODOnBY587nN5md/CHJuXzG5ehKLYGhyKFQvA4lmdIt
CPbw3D6+MhLcDrs2Ebop4j3DUm82ssmyG/SiK1FT6dpFIaVqApeAkJzSKcT9z4Z/8U0NDwPEuIwQ
/iLezDKwT3GbjgOmAH21sv0uDRlEKfcscfbYwDszCb4Z1zuLcvqnTQJA8FaKgUUlGDw7hx7pRfLl
jj5p9OI4P2soPwDgzzV2NE4a18GvkRpEkMIdHoyuBCSxg36nlZWuK4L9oqIXZKy6JcXESMFuDXXI
0F/eIFL/fcjlYaIuZYeIroyDveryvpzUk6CZzgULQlaob5+afgUaeWtP/OpO3gy1CCDim31ZIrjW
v1ctJe8NYEBd6+Gs+LJ/m+DAbQzn/HnBoEocIwoLb8luuHpZWc3Dz6ICm6fU9rIl6HvsTB1ixT09
QDrGlEf1M70rmjtva4IwBF/EG8Puas/58xUF+I1NI6ghUs6UNUxEWOT5tL90/bXtZS9G93bS5/gS
qnGtyBPRp3u1IYZg8/EHig7Kr10iazT5vA0eAknd8JFIgskRb7FQhyWGV4N3wCa+Kkm2ZBI4owtP
hM7pANYuB1wlnTljoq4chwyXmAOYSyiMkAGRQMnFzlXBNMTrcK2vu2xG5+DMAwLs1Jv0IccPXhGN
6frG7YnNW+aMY9v4XdJFs48LBG9qVQ4cIPUUZrq2bg8/aNTCov6MzygrwUnBKT2UvPLGsn+VKtPh
zxCyHYCrA1VD3SXHhWRT+D3lBUlpI68fIADZxq2sDlhoRpDQA++C5D49AyQcmt8KCoyF245kQmio
1jBL0d1Pl39puH96BF5nT+lqm6t6PbZi9RD5MElWy+pR81IUeiOhylsOeQ5PMATnRfZysFzLHxkM
3Du3LCZ3BI2cx3G7ScvkW6QuPie3cl26jz1QM2u129gTFMerkH32gwxDBY0Cu6Y+7nhEB28A36jo
IZe/LIomjYR7qdlbgJ/7yzL8PCArKS4Wx+3pAvZBCzQWSFcbZ5wy7zASMnl7rj29eLoxP0xVGAom
gQOXzjpW0JMCxVjHvuUMf/Cc3KT9i5Gfftqdk+6Zfaf1gsYu6iFD9qQd0xKSjqDOCNw/kRRtywe0
a4EYz/635EkuhtR+kEu3SoxujVZ/07dH3BWvk0b1JNZYKKCNi6iwkiwbnu+rMDjKaCynGGNt28cq
vGLG3ltRvkhKZMWQQ75ssaqoO6mM39Ej+Pk8Pi9QmE5pGnxvvXwpsXDXIbDlmE4FcGH6B7FBPyuB
9hd8C5KlEy4rlj1riWMAhlIX321DdTAYIK6FNDybB927gbnhIAQUFWMQVbnuVZNiKXASdeeT8+2E
IwIQXzc2jdXDVj2GX9Jk+Ffw29nPMKU6fsdkKDClGD/pPNuhSx2pvOdPh0l2kfch85pNsQuVNYu4
SjGaBIcthK4t2AJxtp+2qSjG4CBkT94X7j4SqVR/9gU31OgsO8BJqVahEr/li96SwHPw0LZ3ZYUS
eGx7eCvbzme9ngAGWQqPul4zK0YQLtz5r+7mDyGCwvmgC7W2iO+hqMXfGNuhZt9h+mLtMuBfq2Si
ds7ktLZFKoIU1gu+owOYKO8PvCKsbo0n/mfeHrICxe0gEs0DIm5kaH9dbUdJ8soCOBQPLoM/xvHN
LQyfI6aNYNHjOm09eyR3xtZZ+8rDeHhmGtquFV9lUqNS2iHRkiao2/YEq6d/OSqZDFp2XQQXKZjM
5rdgLBPb4XSnB0zKmIrgj6oftvwhjgid92PlNLVWwDN3PjbgABV+v6sNZyqaIg7/JBCeyqsjZPP5
iDZmLIEmWruI308tmOQWRL08WfOVfEqncZTGIxgl3LKot45YH83l16UQvxIhizSNAQVzb6zBQH/u
3wkIjdzlAT3pEGhsUqUg7Sx2FXb9I4Yparc6+aw3KWNh6v5ZsHGalyWmPgPTPg5ZjAHVHMwt1MtI
qFR+H/cwPGOcQsQ+M5cpNetfyz6G6dhs6jApA8A+OA0kbBwL84kzZpa+KVK2CjyYMjOfxUXVmBt3
DneRW/g3dxFDD0JL+gKVZyxJUA5a5ZT2u3FpQXb90jHVQxEpYZX4iMMwWXJE+rYY2Lz9g4698xcf
I5eGkyKESx1EsZc74AtRDHFc4UZxlTZZPzT8ZtuNj9OypRUapMvjP31fkloVQaNBrWJAVXiwggKt
IhUOfuYS0lgtnS1E6Acg7MMtA7swAGsRmnXf8jn9idjjBO/jkazy5ki7fMH/PFF6p67MzEg64bSf
2kMzBGLFhblOyH5ciX6tvGoj7Fhdc5jndNAEoQugT1PQ2PJg4iEZVqMv/CNcBIxvsjW8YdamStut
VB/ty/UoCzz6rr+D/QlSOPsEUm33WElO8TXgh4NN21KrSKyfm60PpaHSBu+K0GiMnE4ufKaajRyK
HqTXAJUBL7VZ4tz7oTFWHNOKRx4s/dsnVWVxJsdBlbxB42E5pp21PJC9/inZ7G0FqEQjhouyEyo6
nWqQCFi6N7eNnpGKJSdoKgivYwtsPwYbATOaxF+fxOOkeZJi/CVbE4ptfcVUV9FkO5wEaM4O3CDV
Aoj46mPW7CpW1yARr1ultR0HhLIlbPH/hE67J4Rxj9GRhck426KD0I7RT/u3B+MZZ9L/nMUfOzHw
lb0rAMwIE3O4KiDbAVAA4MNAlUAwfQXtTH0MNeeNXchxHeqJHq1Gc3wU0lMTmndwUDpc+4pL5nkF
qknNmW8JOtJdncN4tyIfDtr5q/oLbPG92RoOSoDZGkVFf0NfQGHg7/mTAFak507NlYj4JJh45Vwg
z3ggrP4zr6Q9vfwr2ILbn5RRisADjlipLhXz8HwHKs01Sxivs2rwZBNdaDWfzHOClN/csFqy2kx3
QUKyeA97ZcEUMAEzorcUPNQP10pYQo0U3E/O3pm4uix4zfnBA3AIp7Wo1I1dHSBWIQVvoIra/Kk9
E6kqx8M5cl3qiY7VjfFpU8OFEldh2WWcJsTr/eWjndO364tb6ONbG3jXfGgs//rkluM3afcF1TWP
RbQSH5oWDoKxwUTgT8r/J/VQMCq83UbeMeS1sWIrsBNIVsMlt4bZaDBssRwHyCSYymiXcy3Bwsi3
quOoExGI+a0tBdVR+CbzGKFFc5OxKOcYDwvlUUfovXGXYujZBMG7ucirZSOlAgsf3S2PEXoZfFTY
1NJMc2zO3rLRf3nMZ/rAn8qKTGV2PtjwWBfY99RUD4aGhVm7TnExO6j6NnAvEaq4Be9mD2rn7wAx
i/LrE2pu74zvbHONzwVQusATxMjiHYpaZbLc7xBKhVJkQLWuBlTNhOqf8GHMOlrqU1jo9O+76Rxt
Z7F8ELc0K4Xl2ixiFodUy0SOzENCYWOh7TEbn+SgGA5Rx2ryNb1erQJpXVPPDiZI3kc84ke+pF0U
BOpu5lSMzJ779qInQ6wFlNeiuZXSYDQ67L0v4jPV1PFKpxxSPEvPO2f/wOkYFdnNvoANG524UCP+
MebeFCkEHotm14QXAyrhpm8Qd5RfwRLbxhkm5XUCFOF+WkYlSjpfrvl8gaYCXAlApPeu4qaqjNV4
WkvZCd8K3q+6FWNtI8uefgs/RP8NM9XteZegQ4fufTRVPdWcrSwthFSvUL0oXb3fBHijz7vbdryc
7j+RXklHcXJhv7yQVIVnY5jl/cyDlgsXpkgUp8AiCFbQK82hnb8MGCsiRXzb6RYxZLJi7C9fQpY8
8v56ZCVCs9Sny05VYz5qOgkfQOMr/L3esaTYTVkT/o1QJ2klRzlTinLgM0i10VyF40wr6/2V99QC
MHnEzFCP3kTuz3hmKe8HV4LKguQblhqCYDPiFZoliktCsScQ3/edm7dWozZ+Noad+Qs6+SmA8d3/
tKGcSDbHmgwmQ1wmcui+0973L7FDJkOxstvIUKSDLRWHmYz/7sa1DGV6rmFUkhpRH0/QMUMrYB1Q
tTApEUSnU94253gQ42mv3MjGRsl4I07++cmaXhUppBoJvSaIyAFF4ndS/SsBP9nwjpfzwHwmnw3o
FE+xYKggdR2mycGYJpQv9WtxlfIFxKij3eWaca+5d6iLw/zNARGl1lfnZ0c2LeOmWgvsjSH+BFdL
xazs9mDVlNRzLZdASwJUx6rBKrKuhYNHUIP1HTtHLpSJchheoQ0ceB8YULa2tM5xxuXsZCabwGfg
O3JOK8Yr5dyOKmW6HDisK5Ofl48vDy3c3G9fV+4/MC8qi1UeYzDv9qJrhCRxfPvAFi76DYfxaBM9
53MXVD8lCf1E3S9PDvNm+1hz5MsA0SRjc3ppynnaOAXQLJ7WmiaU0IElzKhQwuFtLj9ma8lxf0+x
pXJuebupe/QmvyW2CR0WSpv1v/ddJg14ratC0E1R6d4crG8xCSOiky+ygwyZ8cGWc3KGpfcWwWHq
1mInWKVicd3hPlaLUfKM7oPfZ+hl6XEOcS4M8iM+UmVyx6WgTxb/7T2kUDSeREAEQ8KgJw/pcjvi
OC8ZYiPiteIJSEXlYUtwFn3vOBavT8kTcN+fO7IkarNWv1lSqG6QU9rDnLBPKM5Pk/MJFFK18gIn
Mh0BVOVM6UzeVkrybtrYPG9OieR1CIkNTbqBe0EgogxplJd1EK4G9KJSplJGDBLmW+cfl4PLUpOS
KpkbJOuuQEeSmpQaYdHRdHw/ye6Bstsf8DhgikabLp4Sj3fsn5NpMS/GUUq5NVDlsUB7DDGP+NZ0
QnPeX2VUuyxICpDR6yGqavd0Jx5uGi6vPB/F9FATgkwh6LdRxWKOchTVC+1EgJ5qO0DL+lyHRK60
J4FH/7FYYWHuenGxT37Oe9e4JGAuDXKidr674GXOaxL/MrxnfnAS7tOJafXL03dm6NQdut9CiwBJ
U/AySWWdG2/VeBzksKwOEsJl676jGGbWMv7KxBlb3D4Ary4741BQV+GM8RkYAL/1LYv+5jg5+ame
L5jfdNCx04eHnkKVQwPQy29b8ONb2akcCRwpJMR5ZWMS2qSAEKI6ag8B3xMRCPQZmU2iq5bCIMvH
aC2kZh1gVq0Ay9r1nlAGCFsmd+aY9j3XNhEYd0H67oXFzk76niClQD1pZCGa6NX882yeRpYfIXRv
2hquKfi6wqINxIBvWKeKds0t3Anl0FxnxxqpsXiJtEvpTZwScT1QxJZVTUXa6ytMcC4kTGupyzVO
RmuRt2EYv9B6vgFwGN+5aUSHlBj4KXM0be9XOJY2iW/L+oO0o5G//QN+co9VKZKOc8oWwy3iwYgS
PnnTTrgPCMBkBmd9azWZMKLBqsV30dBLovlvfkq3W3pLDfoLFhcEixddcs4ctkdOmlnJ0yP0umHY
llN0lRWFax5aUaw8EMEeB3dfWMOi6mrlX7tRBvYaCzQ1vqb6XjeE3VtmfOFi1LFAxuKdfRp02/70
ZKzyq2ts5K+o5YnuPE1+xiNG1szWfCG6uczK3LAi2m1i9VfTYN4TLPoP5Muz38NCAN4QCKadQVHs
4V8O0wfgS6VoPrBuu+FWGn6LMezA4T8gf27LEcaeEINsOe5YkwJDFBsAB85nIMCYHrvQ2JEVE8F9
mwvOlAuvkSSksLUVRhdKxnmzqrusrP1DaqKagCGEn3poaRp3Y9LyY79bUwRNnOGxN8K+ZSnYQ0Ao
AMkigidQdDfQlVizb8eYr/tejVUffatFsHBQJj2OUZCw5nI4C/bB+Dtub9aeXHbwFwa5PsXksRNK
YqB1m/7dl/VIlmIXOvYifEgx1012CB+7OveZ+22aD2oJ9zFQ9LwFbcD9jU7vOESi0GsQtTKkQEjd
c024CZ/2ibeWDMd2SRbmlUraxpTUHQDltm1aw//FCZpCQ+ggV4v8V0Up5D7nUI10YI8uo3FWU7Iw
sWJHWBKevY9HVKOewVNfJo8c+yBvCuMxEbHI91lkoTU5nDCwzch5Gaja6gjaqDHl4LY5wDQdwoVt
rj5GaUlfkldB2701KjiQCLXHktlUnH3G2Lzw0KR5cupBSrmxo71WFRRSndoPOX+m7HeaYQfb7AqF
tOmsAASyDXoYS4kypobPSYD08bdCpb9rZSQvVE0FluvyDv1D7yvTpEqyAR62FbUxSr9ULSqJ3e3x
DBPkNsMjqTVnibuHEDqz5/v7ESz+aD5ErHNPP2HZTQt1iEvtTy/m7LF+ECaTSr11ywsmUDlPn/iu
hHxoDMQzCoI3sRy1FgnO4sXQQ7/mwZf+pABo4X9oAbDLt0nTord9SEo4+94YmDAsPRvvVX/f/HlD
j1U4vWV7ImeOa10ZcGMtlziO0u6P7WFPY80acWqU/mqQ0dIjXRGo/SdeiPt2ZmjBWzO1nVs8Tu82
Nc+WpbLNEjFc6hSFje+7brDut4xusHkWc0uJyPgQffCtQh9dfj0geA+qQlJTfcsfF1ZqF/uFUSbB
oOw8ZmpywgBIk6QyoAQV42atyscki/xSSFiqUU2r1yIUm9JtcY2Yxbpyr7cBusCtisLT298cyP7u
+lZJg0AH84iNzK9wdc4qDaBcBNjKm9VEXbt3qyi41n+xlCjl3RqC2QFL8btMK4o1kG50jEyfy8oy
NOb/fHDY5mq2rTGJFVYL78Vos+O9Sv5z6hf1o3o8AVgV3R22X00vKLWZkQPW79jtERzNXsiYjbsd
uuXX/0xXHdNlf2jJFtDrxj3SiZVpAoE5ubgng+OQqSD/wHLdI+wvEKAusI0kDBOgPhulr75ypC0g
QSOC9t/3QGexiaN+dxrkaKj5JHle6eXC92A0A9FKuAClUKAJ+aT+xK86mCc9CklijNbvWJmamtEc
U4azJuR7OAqsDKNtGSsloKPosjGYRg3a6Q4oFWuUxoxLTIY4huaiL++OGGg4ZhgOPxXkC6LLjnW1
DZXIDnalqiiuWP2QUhFsbSpeg4lwUoQn1GOHPRJVYmWwHy5R4iUyQwWgKjCeuOOW3pwd+OXGX+pN
7kbfbJ7m8hmcpJf2oMX7l3exwR9gJ8zamUoV066STvl8MGGnML77quU3q7V++VbMYD3ySET3F46H
cax/O6SIEqbWm4wkxXftB5FMhWu6LzUyd7Nz/EDbXppHxDcGZL4g/jcmB4XMw4eXemUBxhgitspK
5VVT2XA+gimarcrJ6cQrgKMqQx76qr9MizBTOsZJYlKP2xEobqJgZSrdPcaCVp+V3gZ/LKtLeQNJ
IOlFQLBidTMriboeFh5bCmuwT65wbNvLJXbdoW5lQ481bm43cFDztnUY9ndnxreu8JQmEGqZhnSe
aeK6eDR1U5MxeovcswDvWwXAq1poHE7CTC/pMqXAurm9nVy7nhcfFjwA0Vkq0yGLnRz8giNiF4c7
UUx88mMa8SrDivp7DIWKMnYxTT/P0rXBsWWuUyj6ylpxpMnkh0G/I8zdJD5R8dcG0zmSeoehn9BO
iD+F7wr7OmhhNzYsrvGals5XT+Jfg7mFIaWvgI8idrpRF/M+y+n0uNdsgGlElVK1LKn/Uj5zOIDF
A/z9FQKEvnEC15XmYNpmu/lHAG8lbTWAE8IQhFmawNb9EeBmdR7ZTaQc0P1d/u0BJxz6TE8/ShsJ
b/+3eAKokLndHIc57pCGXjIhiqtXpb2SVDwk4L/DYLRUsRydhv0yDD1rbx7BFCBewQgtxsu1zotw
b2AhwvVcc6dnOmAsJcMME3rEKn9QndxGrgOoiGtFL478KcYONJpyIEjs/ZavykD5fmqMJQUV1VSZ
+bGjeJgPjzsHqgxWW8DWBmxlbs2JKTWQ2kpcu6x3H5EuxJXTU/epGRg4lV7Xum0yrICetu5uywiz
jaHaBeWBoIgDYwUWsZ8vTxgn0Odh9jK1zMQyJQhTdMOdlJncUdybHc6uW0USJ5YkabKzzCCJDVzy
1pyOU8Ii2UZ0WJ8py05puOiI5plZDiS11mze37TVrSn5jiktcLvunHmyehy0JCwbxHQmdP3ImGLb
ATJiGWh5yfGuCeY9vqjOhSXSQFZGMnzY5tHlZd4UmqIMUpz6qIKc823cl/QU45Cip5Sf8H++h3C5
Iv4dBc+/ueSWlBnGm8wqnv4K9IAWbQ4lfCTXNrNNu2bVPDPbLe+r58APTq0op8pGW1Om2IrWStD+
zY4IW0z+1OI/xvTxvCkTaK0+ok7SyVlvXZSOQNzF7g2Z6Md4HclgLl8znjSjKo5Z43KhIiQaUg3h
gN5G6QK0PVAJvWDBKS9sgUhCsH83vGcQfYeQBNQ89tTeOyBuFwukJSIH+4y+kCqSXNiwKap4y5dA
2JWoJk+iG1Bplhb9x36Vz4DjI8YF3CnrSzvwQ9ftDWYmqdQXWd2+yxLgo1XdiX/UpIUTkqfjG6EI
V4MeqN30R9qOmlNOSmEH85yL2KZ8eC/0r1Vws1WyI/bnPOJR1m8IhEj0c5AfQRniuj51wFSy4sLU
bmjXocGeAGrFGU8Cucu8Ej13BQoVVmf8f1ZXKrdtAvJpfyL1VJyBiCtXoe55DgTZp3TB7wkoUYEd
NpYNIqXUxi8CxvOclL1G29Jz/rzeUdBj4Et5UkfInoxM2q+47HkrZJOm902r2/DRbI5grJZkdmpj
weDeMcBZoUxkzR0J/ZUVrfQKuJswlERWhNkXRtMHOtS/seB1+0NH5jXvDG1pzylLnQCB8/GAjX5k
jGg7SvzbiucNeRUtW+dXPlEiG4xifAbWywPLAcMIOtpIzgOuE83rwWrHODg7P6+ZUUsH0faU6Y31
ZZ6PaZ6iNGb9H4Hga4xQuCqkrkc1+vMaZ3QEM5TdwIxe86VNvuN+nfPS8tIpVC6klGh9t5n885i9
s7l1i4oa5s0EzEy4PQoRlsjNf8kj5trC0xtXligGgHOR6uqrec6J0tQ42HQQVGpWB+4XANjV9Uet
hk8wARRH0NkSYxZx3F+XUcrkMaHoj9+rALrvmhZNg93VrqZH1KiZsp9pri15pMImGQGFA+99sAot
a548cBYXYQnV68jmKHYD+r4CGlsvAznLTjCXN6w3dIraFdUJjJ8L33CWAb3qjM8v1iMVvFs3KCgn
SvIawE8MWTcaQuzav08yXjY+lX6rvQUouWyLb8NsKGU7pyLs4+JgB+0hqZzZx2ulmyfmZxkURqR/
uPLUPHayRekMykHz7W+bjyfa0XxhFws7LZVK7ApoUYKBHKZtyThXUDG7Fzn4Et/W6wB50GQFOMCw
gxJAPql5fsJdnBjwH6Gm7m1jSi/DFdKXarLXPvy+0hdJl9k3lNbXbieFRW+Q3NQZzwgp5WWaELID
AUsG0k3PLUIIfCTBi55BvVWUGvcGN0bI0n/5luALYoMPNeKWTuwNuvUgC5n7rBbrpsfeDYF7kqLM
n4EuH+JhtGB16Oc3fEOxioA0knQw6uKNRs2o03ghCHbHMUf2V4I5cirvK7Y13HjAKnruiiJyIsYj
8OjfJk6eg0d9wZkN8mZNX5tXIj86pJns7dPzkOhb9DILsZHirO5cFrovjC+jEfCnCCnAourqlPVR
TmQ4hqa/CkBTBRPQULFfQmsDtpiNy0bqoZqaAaA5a//HjtXDR0wXzwhrbHge9nlL2o4PI7abRcf1
84pLx+vG5ijwxaqJCbobwYkRJpadkr6lvYb5Le8neKxkqBl2zXKFQQjXt6vtE55MAna8iP9v6Rxr
Mrr+vmCoH73Hef9p53T86ZMBNN39K2ig0RssBcbjolhvjCPvEVgomgkYUuImk/MEg9V/jFB+aJ2H
dnNKkYCeX6FhIm828NUjWvq14we3kwIjQoCaqHa1cHKb4mGG1m8VbXba4DWSxJZuI3PqJkVBflrx
sASDq+WjchkfYEhiVAsKbyuxbDtG7oAdbAdb/CoPh4uGs1++wBtjYRis1/XBgi+kV8P5qSd/TdTH
Ppp6oYUc8KPxPWBCpbUSFApW6+OWuYT0SVfiicECDUuZTgF1s/jxJFUzQmP45qNgbxOssqzwd5gG
VTUIdQuiroE2XwdBTaNhW3kUmQIFVbtk/90ds6FUVG9hseQbV5/kppm7Mn/CBscx8hVahyiu6wFK
+BNmgvRHSLzYuKWLQd/sSKsLx71f2MWOU6btIFboJcuP1Hf+oLoMYIuCLw+bd3YTOiqEV/QheChE
61XDiG2AF6FCIfRRh+fwHpwjAiogD64bfQpRnT8L/Q9KsbdGE4JwfTSmUwpyamFn/NaBZfHOO7Qv
vqfD1AjW0PQQv/kbl/zAPbI+zXAJrC8cBr1NwccqySZ5i93uGYYI/X0mduCl7DDoKxLjXXtpINi2
/9kZ+LaG7TC1X7DvD10eRGIsmTYifrJdUqLQzxoWmMoawDTk49Kf3nOXDwHcyuRVtrwoIhTtn234
Lg8SvmetRn/YuqlFe674+1YHDjsFKg==
`pragma protect end_protected
