// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:35:26 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
btZ9qlZGYfVRY7OFQ+3q6rH1c57S0R1sDizP5inAaTQ9nrPu4ZdXpOMQjL2asfVe
IejZUyL9IAkNT4jTvGcjfaRUjH5BMwFYXCowtwe4KarmiUJBwYtI3q09nSRLutWB
OrQw1IvDSOVI7u385ZJg0qiy9U7fX6uTvSXvDjLmuEw=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 6768)
l85Xx7Gp+SAZN/MWHylEwgvAN53c2jQV8NC4r2gfXVGrYV16kMpWU+wSkwmd0kAd
+8jghxBxqEw8iH7zhvQRz3j+CqXtevTctRol/tNjm35fHVAwoSs9SlClDaNT20D5
BQQK29xXg5DVPBKqRPfyKni3sJWWa85Jeo+lacyXxCwNQUEInK+RFeSipLnNbb9x
HLd43HPzxBe+LXOqyAHTUfEdur898p5Oy6/hBGkEfzLMyPBzJKodY+eYuAmYUNrp
olpEEAuvbLfgtHyGMHfJXscl/gtD1aTussKgNDYXvXhFzhOZXhkMMhmnaw1MtO2P
Eehc5roMy/+zIv+OsCPEV3nkkOfUX+4bKUctWXVyPsaNyY0uHPNFztpBgpgSlwrb
nGKZywoHr816/28LpG6VB4IUeO03LMEWVX+g3aiK9rAeQdxZXQ8sDKpQ0dXTE1YJ
fVUKR9hkrQp1q2/6mzltcFs5ZkILur6YiLWstGxfQ/eYCLasCcUidLwGGRWlu+ru
A1dKHcpw/GQtwafArcJQeSfJ4s7cF3hhWsbKrDjpxtNZscLpHcpIynfcXdPHDyL/
ic6osT2y9JsJZMdFB7CqhBp4IaHAtVZhaxe12QPPPQbu6yKsnhzcMyUWIdxdarRI
bckm8rsU3sMDcGu6cTMk37vUp0GEsH2ONVzAcalSnGREO8YTo+uMOmO3vn5Yfg/3
L02ckbvifIoWsI06vCEaEINOqCFNrCT6rCb4qYyiXQsh5QIILf/xMN9D20OYIdva
HtMGsFWc5XirMbv1R9FQGjTnLZAmU2TTbkZjgkx0vGO2MtTyEfewrTYmCFVncSip
KmIgdKPmqICuVTzvLPwPsBe1CfqLae5Y7+L2so10LyFraZbqVSMLu9gSX02gfiKo
v4JmsAGhiZo2F6nCr2x4UOLaAGegvrPHC1Ddid1c0WwQ77e8aX5DBXUwHlswfyGs
k2hXi+GoesIKhrnTeyNkP7pYpIhVhIYiemy5iGaTqLllBnlKQgmPBDqcHDMJYDZJ
yLBOBE2IF/buFNlbi7z5I896yjV7+3r2B/ljctH8tnMZUq/Z8Sdh31JnhR0e6tU/
U63caAgKbeljkZRyYapanIDabKaRTTuP7POzNYEFkle5k7HaBn8/KXswYKVABsZd
6HfZs3aeVBHp609qOya6Et2PkgRVvB99W6246SEtr4M61Sk2kEWzzql+qZj7XEub
fu6pnhHQeJU5fA1ZHR04bLvvqKcLuZNBebhVhbFzo+9ur+QspleVKLHra8yj47SE
pZ7ashUGogw/Y9kOWiy3AULrA2KmJFzbXGggRvcGqYAKMbq74yWdxGIxM/Be/OVX
XW4qbvtDnUNhKlOHvTfu9WdEBJ+NY7cEIfylvf6cEsJAYyDr1GOaVcVwsR/Jkq/v
JzDmb/EILzAeF27xEFIboNNb2QCuCxtuH7tk8Y3oUcMcD+YTWHTncF4r+WOl6eCU
BV0J24bzs7v9wjxmrgt7U0yYX5e/GvLlSRSuMf5FU+C8k7e5EwGgZLebmyfiTI35
vyfDvXkaoBO1niC1azgHCvbUdhKj9mllh7wpAO46furtTp4zqJsAUedDtF0hsO/c
jKHMEwezEiE49DARkgyOtvERyh3PaH90PFfVtFiXju4DjJNg+FjodPXWYw3Fu1/R
HXptgw7tsn/idumUpgUwgAxepaQl6MJb5nId2preRfyL1/7Jj1BQaCnavoEwOOx8
M0zLZYKOzOcsKU9xObU1ADRCsxleSd+DWPX6KpvCJJFYu1gkQp523h0JJ2wwCume
yZit/GpWkV75gRUZf9pK/KF5kmT8lwl0rL+LyMsq8Xlp2N86SMKbkk/jQ1xGt5kB
/RNq3JBx51V00mMcvxks09viSZ3FrJvDUKdMp6c76gonZ8KKyY3g6nJLhJdpPelE
7YZqcwsAkxQ2OzEWuwy6xaKWor5O3NJxWEwIu54iYX/D9vXVXuieQjDwjAdiBzl9
9fhGcvR6zuZe7vwV/EELkrahtSPQTe7Mr6RLQDF05vuKA2sxW1/Wxt3AQSGZohZE
60BVMHg2J+gbaOZ8PWakVK9d0oR/+cJzGpPm7a72N5upKoWJwmwU16gjvzuFjfBd
yHYn+v/mEFnaKlOxa37eqnjC9vrHCDQgaMoHDzPgCL3JvDMgr0UtZqwRxkSbNUy4
SBYrVC4LqSgKk59DMjTVpuWVpzt2UhS91RHQBabpES3L4IIA4ToAb8thczlPuJxP
UzqVXMnwi5WnPXmGBAu+CpGwrliawv6u+m0+moMwm0I0fAvJuFacGZUWEwinbNY5
rd9ulsbHlu+SUC876blG7WagObRJDjQKd/rVPDYb+HfQUKjQztpEvh1gs3u0VJOd
Ypki7u07cp16clFrzZUA9pGl9pGzgAJCOaHvv+8E1KFHuRYk2Hp5HD6CeTwDTo7J
zxC5qOiQTS2gJBWOrDPT+fD5McKyRGZ7opbnm8MgSUkjv0RkuYCnWLTFLn3lJ7Sv
Y3tXRTrIabRd0Y030z93C8TjcdtFiYr+7Zgg/vFVKrXU3klg9hRuHioquMIKjGFp
YSvEkyqLf8QugVJjLPcfWVxqNO6RJ8+jy/zRx1oj3j22aWYx5NXgcUKArR3UUTSJ
5XV9C9nTbH1P62kL3p1Rjv5Z52OF4nM4e0yQ2XpiZdeHAkfNGQrph6bsQx0YrJw5
IHgGTiRmikUVIrmm9f46jsrzZMRVnCzKgnXdta0FSpcuy51NaxvRaSJrpsJXqX2h
OGSE6DwNabG8UvNGcgzJ8hPyHhKa5a3UoXbUJifkTsh3s2wgUAgAV6y9L2/CmlJ9
YJ33Fx0K2pH5kRYG1EcC9RWfqTuz5FZpEMf9zcKqSGuyfImOZ1ps/LInCvSEB5UJ
Sz4kkcfQD34D6izrlQICeK83q2zcvvnIJFGPbL0PkzeUzpY4dhCMnG2j2kyiSUET
UCGw7zxrCP4N+pnWNabEKZBJvnyvm8Pq3ngby+yyiIXfu1hZNmT3G7UFUw/wvdVF
qSrZxDfgzEomVnAbMAddnoLoTWg7cqatdRCdzpg4IlcPSjY+9l1IIBjgEJfPlf/8
ZmCQ5cDs4QO4m3lt+SkssYHJkg3kD7dBPTbYRqUx8ryfWVOW30yWV22C67jzACYF
xBGVx7MYGuLq4T946DgxgBX+q36Ld7t6N8GRV/TO84eMcdFN4TZw4MC2d/xw1fkg
lNj0kAyQOGSUVet8pDnjyE2R/YJJzAQvEwEIunvjNknUVg32M1f1dFl6daCL6obj
LTpneTs9BdzC/NPto6hP3h7ExgVDgx8sIZKxxpXFdBOBp3YjqgItjkuKtCMxRs4e
OZa7SfpHylAwPlmwCv4xNoA6Krln4lEdfq861adlgzvA5F2sdV1RRCndjmzLZ1ia
z1fdMaH7HRRzLd3KF9igaobaFL7W7t73cj5ny5IuGdY0EQ821Pig7r1EC5hxmk2w
vAd2yfd/7piSO2XqZuH98VY2vd4S8SHvUXZ53UKTgkklYrgawVJhV3Z06SHMMC7e
QGLJF6N8TgkTubmuLs0cz3bPOVSfcWJwgYW3HrE1jKTyyddx9bBAvkyJhAUlADCA
X0u/Y8rfyn9gpZTarNW3b6tsrAUXtObU/7/xksYIGF8fZapBZvv4bbYJNvzVPH/w
7iyH8vT1fuxjJfZCHeTh7copwfs0Rtb4Bv3U0c9INNFcITIELLXN4RjIDSK+Vwa1
TtVmUgNnEH+VQzfSlNaXz9aZ6nXqibSViXZ7zeGqxCnhxIfvp6WbrVATTUFPJ0Cc
/e3Y3VL+ieSMRjHFP/r5k98UA8Eid3C1d9oEK5tJvqWZilydpUlDezs480avEMoA
BhiitRb2npfdPN7OOuy8BsD+VM/4Jh1WFuNTb9ppqgqWefM0ARk3H0Inc1kYfH69
EQnjPHC/1fB6MbGKtsbBSjKvMiQIa+ncZ9TIsDpB86+QWD2z5F5I68jQ6aQml56f
tyaPsyY7f70XfoyDUzAadxqF65mIvd2eozyPdNJlsT5lEaa+FCNl1HKoWzL1p+M7
Sakw46sTvNDopgd7/z+snrp5ULkOvDeJYjSOvA3gwXFbeBUg3k5ZNfZ5J7/c3ogS
E3Uk4728/QVRoIWG5jEuZO5R/MZGgJBRMReQ16BuB2IfECykoqcJlUymbLz7ZLIZ
nXmU5enx/SCawbVWT2ZwuL5fYNC7ZX9Md6BW8fNzPA9gtL3NxbEeVlnBGWZMwAJa
pyWsyHOwAT+nt23Hi/VbNU5g55TB60QlaNaAw3KUwLoBzbasBX18zj4k+2ZzUe7C
i4bvOAW9GD/xp2ARAUh0IOEqWgvhqfpWI7X74uWrAYI0rsXyvTSLk6AKkAPTldW9
i8O1gd2W/EeeHiL0yyd421n5C8UInsMrlY3/vfNxnJLMmUwOS8hSIzd6qsYe1jhb
XCyyNcA6dCceys8pKNAYB/N0Uw8xKxqK/i/deWDaB7yaPXZDlgWlgBe6nL1+VTQP
1pvMosCptQwG26GIIW1XYdAeGnH/3bM76GiU/IWFDXzDSI857yr+yVNaS0Kn41rS
Djt0WwJrYZcux6XUD+5ERpSp2Bio8BBB5jcFXWk93SJf2+ezN6zNetdSePB6sTp3
dwaCGc/2SO3YaKcpRSgXoWVgbkRddGdWqCEF/9kxMK+dm3M0DVgM1cjFkMPO/vXB
ylKalL6t+weKrNIIGanKq+aB2JrjaaBig/Cc3V7qs32q7WQq6KN+T3RX3EKFEAwR
LTiJqjZWHXYqIhR35rsIXGauPoHu/rlVB1f8L9t3jrJXwsPygC8njCqNJ2OWn74d
YJtvLBmVJ0tkvL2QzMS4UYvVV2qmLm9Yzwq9mmgOj/CRa5OFTsRwarwMRxGYyJMc
Ye57+jkY/ocSgjrid7HiiD6H8rz79jSRkUhq8dft9+01SMe005M2//l5kWLGMe0L
7GxeR4aQPcW0abaKRzCGyd6B5gpzyDLgIgIdwMhincWK1jbfHVoxfquRkYCvLCt4
dx3rJAX3hyFMV2iFvWwxTBLy1jemx/PfEMRf2GHVQ/dKbImEw4F4dUCd1oPnu2WY
D2tqaDeWRhppD4xBX79XWp9ctI7s2kNr5WdGjOLm2dh7yf84mMIEPxKOs5y9ydWu
U//U5EbJdD3ulHKgqvxsSE0arOx8Mogoyu3yE6bFnOTt1HZ8mE1jMsUB6kXzmYeR
eEraOyEdF6wH9x//ntXzgcsQ+Qq0mypXKcyLm5j+jBUyODNhI8Ad0+ae6BDe6gmS
+rzNlmSPB7VpBR4YoTcVOJHE1GDLRm2a/390H+5S/JEbzv27vAQoco9uZ0A848qR
hmoCFmBOfN1YvNqldZZhtpMt4eJqHhim40gzFfcf25VJ7Uj/VtFpFzn9ejuJN+Lj
/rurq8Mj/a+lpn7/p5G5fFLT7qs8K+bXCVJ5gzMYWUNNztLL2nTVloezyIhHNYat
dePV/f4J92wTiKADBG+ctNE88ebvKsZ6dPhC6arvjXzOI/NjY4vYizXQ9GQN3c3z
yxcCPqhsPJw9dTYKzfXioTx+tVlr0y3j9VLKTAbUKcqDv2J2iTay21IPuSq02+ks
dwDdF8RixXnDbLYwEomN9aWFfMnxUZeCzZamkdJbprP9YlnaX5Q79ND0Pk3sPaD1
oUpzRISM+Nrb01BA3BulTCAurq5xxL3Kn3+UJTqth0rxb7MDAwx4mwXVmgZKsxot
ddL4IhhCkQXKAyp+WH1nnElsOTtWgTW/V2IMJ6VYe2jWbFSMkzQ6rqToX+xqVN+z
26ypBEm48vt814TzqbLcC/gq7yMbb/odY6CZnShPjyJ03qLQCEn3va2aTtcc+D/j
sFox6jFtO8pP9Yp6ndlj75ETtzx4q2ePMRnHMEOPH2PRm4zdpN79B29WT0FR/VEd
TqPavzJWyJqzWm8ltd5Jg5HnOHfMYzD7neGEbp3qJQBxdMvMvwMiusSoK/fBY6U/
Cbk9LRGuiUUpauerBGoINqa+q+AUGw+/w1zrXQtUXcindwjcuGYMaj9p1KXqHb4J
vYqeWPCRsYGnFzpp5klWif4miT359CmevElFXBChnOn6MMDQV2+Z8Ydgm063COyC
pcLpHGBNisiV+0CUV6rwJ2xJs0dWOO8BKnbVcrLlxsvTsKMnDbdvWXvwwstXYDV7
MHm5mD7qrFTRTwh7cPG/9vn7CDL0YgRrQKSvigp8xMP/vWEnna4ybQIMjB0g5ZuL
HTpl2I4GownlicdppymZT3+LihJUEtlcjI0u/uC5O3Llm4LAyuFNgJzpXrUSxBMF
iyoZrU44j9aU/ssZh8qtpMk1CFj1QoscXObpIB5I4tyGqpOYnRnEkX9NwxZiWLQb
dGusQ43mdBm0jb5Yi66dHqEwr7wbqsr+ePVX8DBRY1GMssh0DPyiRiKBLs9f3fVB
Hvsz6GHkVbDuspcwHura58OMTBVQ81qol44BJsGLq31jNBbE0wpibkuF3zq9wX9o
vQd0WhN4iClhLbxta7CqKSdOdl9LUyE3JXaqAcdheT8lUj44aZFIy5SpG6/fRcRb
NeM2Xm1j7aQEvHieMlE+NjmSLTVxqHIa0dpzmvq/IFmmVDSomIhnrO2FeTryzLPz
8tTHN184Sg8+ZkQCE3PV3MfiL54jo2w8i+Qz3KomflIALDWcYExAdrAmhposFO5K
tZ5baglle7T1xnokBSbOH0jYs7BopPSTZPMPYBrw8YKQFt067sxEIj9jXPqce3S6
oXAK7oouzye+T6qn+fqaeI4X9IlLUsqaPD53B650K+8zLVL7SxiNPpYvId/isrNg
AmBRSb9KukLqAaRp8ENtm7o1NJz4yVzMMaW+8YPdTHd1mJOIYHmnA1HOjW+rQh4j
Zy1Ke/6OjOzsDYInByIfYfuOMok34Qzy9YgygC3Eddcu832H7q5n06+RLO1+VBy1
SftKlBJ8yE1DJoWucqAQZS0e+OHfD9el+Bxyom2tGYspcByYHyO92W4qUt9ytnms
E7JgUl9lYmcVMxy6mlkJ5e6WyybWmegb1hAgOgqfrEXGjFGrniNL2+hlvLbsOjp3
hQDkG6Aa2GdIkPtxjKTdkatPpdmRWpcK3lFKD8br3ow3NdO/9HyV6u3bmQwOoumh
kFOWBMSAVKMxRNDpmOXnr32YCbDy0GZzQX07DmPhfSglHxJBvCb62FIRSsxZTeCM
VFJeds8WTRT+LzVuitvnC1IqmWzWyMP0NVzWIem0C3R4BCZb6RLX0GuI/PvkKJjT
8cQmEheiG1/BjIbrECzQFncyt6feemC74+s5yJT7LVTWMPL+rdctLG3c7K2ipuPO
txRxLpzuWmg9VdkiZhC1dUeEDwnkAPPYtHktsvbXmItIcdtZvFQrVlOkZiTsa7Jl
vZ+XN6qnM1u5/wynzV9hSLYZRoDCPSZpU81ytbqJ2zneA6+f2NZB1QXYpigsfGlc
by3JvKPz3BpA8MYBDJt0z/tQceg5rv7gdyecnPEXpVPp5RePsEkjUsdYYokkh3Jp
LvTDpds0IJ8RRHAV9pNbAHGoGdHgdQciFYLGrFtF/5kzWTIb2DS22sN2YVamLw+5
xiJwx3/XH5eVL2l7x17Fcmk7KUpt6mN3xi4rm9UGkrtJCSBaRyq/ELaWsi+N8JlM
8dZmblrCHneILk9r43PGPjwFkhD4SVsMiNSNuqH9dD8Uly9QqZKyBdO1x6HdiXA4
gt7g83BfFv009D0BOgH6c9IFK4ye67iXbi6eRQSRvNOgIbVEnR+KK7B5M/xqRNpE
/i5gX4vzSCejIoBzYxIJ8y72DxR8Y+yoz1T6gYDi74I6PEbh7LKleSJ7AP2zpIEY
zfbiwq+hnwhFlIamyN2tQoj9qotLJMA2o4vASEioQjYomYRz+1aDyJ8h+kQ23cs1
z2l4oqoG1hVuU74aMRQt8skHocMOg307yxpWIGuXOif2vgWae2yp5KL0n9R6i+uT
715PdCm9p9Eomv2teFpyNPEfLUtFW9y/ujseMx6qRERpekdN7UKoDioAEZGNzQCF
aTINutTrv6vwqkCBzA+l3a2pYO3f/dlae1hRnIv7Lm6oVxk1X4qgFqSCCsR7ZVua
2Dq/r21FUZEZbp1oV1iIxMhg7H43Bl8CeSZwpyxahAAv4+QpQxSqCCibOTTn+Ned
gHRElIjADtVhCkLCL2Jru2WGiJxIkeqAxZ9En2skSvCIAzY/0uekbz1g6nBUc081
2NVuwzVYgVQ5v6DAjI7gsw/UpeYYOShgNzDv5KC8TK/bg6IW3r0ui0dmB+snM2rh
SSYAeIr06x7tHEkAd0Q/Csq3zQIp38A4cXo8zEaYDpnvPQHLCnNEdmV0/r6uKx6D
mh54pTnmOL5cUtt8WfyzayE1nmYZWtrul9QohfLIjIiDiUkQ1vljO5c9NCFzdBlD
z6vk8E/q1YZc9Cdvgsqh+hk9qKln7p2AQhu9rbtcRKcJSwHXVFt34czWMqZ45mNU
DrTWVjfyDQ//W/m/XQjRT6i9Zq4mn29fOS2PztCJMGFiVhGwRRDhyegMRnEL3i3a
eMuK15UU1WfXJrFFAxC0v6wu/0F2PpSohFBhAtrc96yX2jVZ567bKpTksDpngz/8
8d93uAiaTq2/IIAjMlzR1nyl8F9ATNnBHxoLOIio/RYFFot9mdivYgvO/Fku2qvp
a5J0+16Qfc3S7QOc+0gAM4alyscQE32FCVUd/WyLNohSY5k5c8/AdAPrvjTjWXs+
4aH47adyq3CHzLjSoA6oWO4qVdRRRpjy+hPb3dy1ko6Xl+CRqgNGiMdqsXWcylzG
4qz3pPTaevjy16jE0fthRsCK5w0eArLjKXpPE/eRvNnEIbhCSO2aKWur+zHnHuQO
mpTvOkeit3vnRSccvfSH6YJlk/fzfJ58aVy/335kwAWtv3ig/XHGlIzM/PjHHxxY
Heu72/3V6/1hvE500T7XeZ90k8BffdudOWO6jErM9kLuTlUDOQT+bp/yqMp8vw61
FnW5OmHWv46nSoM3T5rROCUpV2BkvhHusi70tT5Cjd6oIoam/lyoezbClnWbUgTI
`pragma protect end_protected
