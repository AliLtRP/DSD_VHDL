// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:39 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
UPa+CKtex7Axluc2+5CBn3NS3MZkLQ7wBxDKwOPxfv2sOvdLOOIaX006p/xY4pnL
PSm+xMHvwlrp+eIjV08CNp3+3AvsGUkymAaTglK/wlD6ljhZGgaI6rlx6ibK6tHp
dCAJS5QLwVRNs11gnNnGH+NTpkQwVu7Fh0OUqjdDwic=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 3184)
dS6EQCGwoyr7AFEcIjEg4E/89HlsK4R4/oP9CO78DlgcvQQSCQL62VvKsEpupWxx
m2ymjiMaSC9Reof+HenK3pco7yvUktxW/ipz23FTDAWZkrmV68dQgbGiytHoo5JB
3y2raJOJ0mvj/9Ow2+RkXpEKj7G/ME4g3QiX93qFBJtkkR7+SlZHZFhR/dFJMPSq
qW1NlB3FQa+s6s+Pjv/1r95F61S+h3fPfpyZplzvfTM8fxefMubtbHDpwiqcQkbR
BpF/y1sMPbKLBrWX28vyYXlICK6Qdkw2jDGd+EScWIkII1IjZF/yKk9lPUndr1j8
zk/PNTYM3s5z5dSDAQL3UY+qcuKXwS1jYpIP1eQYMW7PcCfDcST5aFCY3B9OnhO/
bXWIGv8ed7yqqX9CBpPqJBj+kh0d1Qbhv3MmAH5TKd2myySfoc5VfeacnVtUavuO
iJeXkLGBJ2h11saerPUMyMDz/eKhBn7ojDBMRQ01Zpbde0HD8lbJY0Wc+ROVrq6y
BohZWxxNWSl899OMdz4NEI1nJ4TL5puConEIFFmT47L/iDt7TnOV/lZZdztfHV4A
kdYdk003vGkYmNhAro3S/Sxm49KaatHyrJ5FDmOzuXuISMWOB2fhsrZNiOkh8YLb
Udtki6mJclMzm8R7XHO6eC11t7e6YCbkooJSf5gqwXTvedwT9VTqG14bkjpgRUXj
sPgboznS9hW1LMccx4jYAg9nFfOOP+p2VkAP00BSWvWb5S41lu0B8O27Yvor0WOw
LBejqs9GO4tisl/89xkvinu95Kb5XFW4MQpWlX2T/3bnZkNgWBboTS4kIVurBzbd
5AEnqPPdJqOBeLBBqD4OTz0mVqmQB2Ef7gcr0VwVswQJbAaYw+BKqWbZ7Y3X5WFE
YfoZDY62AFJ93w/eEQhzYcOdJFLgbClkjSvl5rctzyGJA5EIYs1clnBBp6cirv9A
dFwgAKIobcXWmENPSFRQZRZV/+eRZzVleNYnBTsz2RoYOmb2qvDsR4D21lxW0e7P
8UGGntN3J6VgXH9H8AOUzXthRhQImvPvbbObu1wEBctkwHGLALSkWgkx5H/rzs4U
V4f8vVcME7FAU7YQIHfYdGM35KAJqeHA5gilHCwjl+q8WIkwRKFDjxRo68UehhvH
LMtqMj+AhTOGgtn7hHcO9r0iWRvgmGnzsw9QkmugZtcvfEqndRiI/bW1fakr0QHK
D/rzPmspWuXOEZ12y79TJLpz2G4sMAAAX4preCMUmatdQXjqkqol2c2IN/ZbwPo1
r5sd2p1gUIq7+xYVqDZHx4r3c0BoJmNaNzn4eX5FH0yNgVfd+XkISpbOu1LG4CMB
GCPucaTCyA+bozktEqfg4+hwjgYZoL8C7JE1d8I6P1hFANzkc/D/AUHOCiZmSnmW
omg7fw9VjsTGrHdkeKcy2oVjl/48nVnEwc11Fwvr4bojE2pM8Af5UAvAhI8t6HQE
cJ+nOwFgEmF0qqM7LZMG/25H2RYhFtbJjKtYZpSGI05c5Q332pEQ2y+h2/4Mjhoy
XBNs20ly39nNNrgmlKK0kW1zKdNH+oMh6osF8DMJzivUqofXLB9Sv7OSIjqiM6WE
BbXURl8Mmn/g4a3fWhgT08NrgHc7pFVVD6ayd+L7UxjU4D+6kgXSbje5dKbqk2ZG
kqa0yXwxfTw8EL8fCeMoMc42Mxawu5JiRhBTy7vj4DeTyaUkiRy+G+SgcCBel+Kx
oi85eyoMd95NDbLJCmjQwg/nTLEmiQqTRXCbtfmNeBTEYuQcQY4dxAyX3SIUOyzL
KwfxPdENBUmMVhVv2K+rtw8hYczSh2rfwMkfTDHdajPT82t1adHnz907x9XHPcSg
6EzkbPj1P4pZM7Uptrbi2xWwds0KgvEZUInETI5yyE//2VKIuQdV3S73vjrmWdrS
KpiLKjj3LiSBpptj78dJl9mhtfIlO4WJNBAq6Uy3D6lDSF9xPrPSrnnh4E5i0BJH
Ohw3hMVZvht21NlAYlHcQLuGOwbFO63zHJ+KdoZHEXtRG1knAqOHySeeKo9AoGrp
GNVACDO8F+GWqHrIvmgVl3CGG/GUGXJjsWwFNcs2xe56loSCLH6QMCKuOXy15YeM
8wilExYipqDjahBq3HubYAQiZ2s5SszG+7+y0f7e4g+9/62gc0kd4clSihoNWgcO
DZ2b/6HK2mOLmM+7kBrY6INqsQaCHJ+JRKa+W8pujyEN+M5Cqy5zd91Gqqdltnjq
tvoFIqdbfSl/Pmh/20ki4SOqCI9MLM58v5DMbasdzINfVtaGZ7UQouynWF7eA89D
E76qcnTClBfcSRWYzJ8fZO0hgcfKi1Zoy3g0EvFXF0cd/iTtz/u34/o7sSFkZ1/n
i+1iiTPMm5RxIhMo08ickRp7KHllnVuzII5FHY4eTD3XEs37jS+Mh7WnHwJXbx6P
Hgo2brND/r0md+sdHVQ6bfKtBcSEtV9lyHP2Cl78B3iCq4dm+U4Kzgk3Avbb0G/+
zU+6E8mZQbr7yH+keQw9EjW5hKdkOhmFxcruYUjMC+TUa+DAK8utSnbwFDC5p3Ud
QFRFQwBwV0bCUibF627m+rirTZPotOOHOde0T3vOoK3vRs5WJunviO/UC7p7b2Cz
u9a7Hr1TbCLBQnmMn4eVg9nvf8iGVRtLu4+8HoVpqZPORT6FBHxUWxIXB4SOGXjf
BQLV+UrmK/j+Jhu3meQV8E8NS/erch5hp5D+tvUAngiigb/ziO3Qrhx5SR2XBw9M
wHvTLyGBWB08AYjR7QGfDMez24nnXoCaWYbKLZCQBl/ltCp/CTo5DiWO2lc412YZ
+gKBuByJTcgTdRLtUUBWvvXQjmHOwOtiSz4Xc84Sccjb4qiyHW4fqlbOuFvCjxwJ
sFUuXHraFUIlaCfZ0JNk1ySp/5pjp2ERf24fljRDdof7d+3I9c6vp88faF3muQSo
f4dGzm08qDgTGtFlpQOKnRFoPNXxpQaui8xhHDb3uI6o57gbM6yAK7iT+pi3EXlO
Z66BW/U/bfs16fHutx+QB6lNoeXaacXsHVmWnl6m8knMe8T7dJ3/S2UQCOCCH5Ap
DyTEb/j1mbxufnpZyRg976ZLApbJKHLjAOCL/QMAVH60vNUTNAWe6x0rlarbQ/6i
o8kmPQZGqNOwZT/i867WwBgB6bhWPwInwrV+IIjcTgKnSyU7ywmL158+hDqQEoWS
ZcxH3wvXsBs4Ql3EYgyTC5t0cPQlli2J+OoNCW2o7OA2IksH6zI46FneXC9gQLOX
dEz96cQDTxfTrTQTtR+/wFxN+cuGOWQaX2ZGDfo1M9jUCFL3ojkBVaetArgb3BSa
e78QyWenJEFcknMauPq/2/rWoRQ7y3OQPY/+ZOXpCtGgUZGSb5oQJRxC423rcSB5
T/u0Q6qkzl2kxBeMsGj2EfijRqWGQ6sHltPKgFYhPer78FgSC7TRQQdTemd6Veez
82iNIrRfFmFqaCKeM5k+7lXlA+FzGXfS9IT84AdSuSDdhjcxkmx6wYsmao7LUyaP
GXRGLifjcfFrVgbzSW6Jp0ptdcbkNlHVD5FGlkoo/4+mgj5jys6VQfL7EPTu50gY
Dwk70j3mS0hciZT2Q5LlMvcCuEp6gSlnfviMuBmcJkXFT4NFup9I/4gsPgHZZdNR
DmK8eDBBTEZxeqPPFLKbGmFXKMurt7wcFR7annPbXXozY/ExJwoyeaUG5Aop4awx
mQ3Sn/B7S50Hx99lz7DG4qejCf4ldbAPDVOOLP3nyonZkWangznZomMtqya91c6z
cBblUBGoP2bA888xXfWekU0e4M0/ZVxX+v2R5o8jqTkrRi5C+CYd5fU7CE32fvlU
cZsa6IRJbB8v/YpRVWkQPjEwDJJQONQ51D8+xRyGREfV0hmKC4c4bx9FEJQh1iKj
hY5wgUJdAmhsJ5CBTnEcO76WiG1HzaV12PxplSeTGNin1+ql3xs5lZYwa1bDtlSn
fg3t97kZXvow6MsrFCeqF5ePE1CUgLzTD1/a0241HLRcXzLNqoeTMdn7eN+sTcAd
JhHINEXJwe2uv4snA10/Ymh0hFpFTZgOJE45eTgBWvgY8MthLZETZwOFExa8usyn
hPd2U6TVCKgxnVx3ef2OBE3c6z9whTQcTCRyo5PUTmmAMT1e99r0Gk8UJMMWET8a
KzNFH7jKNIo0YIa3NDmnl2ldGFIWeTimW4hd68hKnS+7A973691k/hNC8gksWSur
K9wfkWLNy6p0HxjITM5A9A==
`pragma protect end_protected
