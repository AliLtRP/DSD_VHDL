// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:47 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
HDyzvUT27eHP/g9ijGhvWPwNdbGlQkN05QdwN+jyEZUUuXAWeCB4+SCbC52PqtUs
SFaibsK7T2MQv2UUXhoWHnDtxZerRGFIJkqUWeX1VwLSs2YbdLo0PlK5KriHk7UP
eehcvs7R0pSPS51weleDOX5cl0PPMl0dm4G6tGyRiuA=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 41424)
2SWfuNetlum2yjk97r+Iz7tsKpCS6iq48QNspHn+jafBAGUzmihgygaQVM6ySKo6
qVE2iglTcxKjlmJlZJjn3ivb74wGLuaW0L71z0N+xKxvE8AkhhXBEk3YCV7gBb+H
MP9QDULE6yLMKDCOM6f6x+Fykr6jm7F0p29G0CJj+Z0eaExn6bMv9ZTUX/vjlUnn
HO90mkaDEVhEKgFKflaRB+PO6arJINcDfTiIees7TrEWukaNOcRcYVI8f479ILpn
VXYwpgoXBYwMiKcI7HM9NjJWncxxc+1HCe/RuToBotbRwa8MfN/FGgDF84pwiraf
uucYM7sCmbO6ek5DMt5jssbFzrg4TFiJ08zZycVfTW07Jt+cE+90fnlrU9EZYxBX
+7lOwQSGyw17IUoBixMsPAqn86VL3SuX7ThLe78qX8Aduix2nQV2R0LtjXbk2q+P
5YPFEjVVg9u06ESZCYQIYn5FKMqdBAxTqUtpdT/W6RJ3x6Lt3EEE06ii+EqOe/gv
FMFOjqZ//hNO6b8I40PsiKfJd5dwZbH2IFnFJro/aKrdYUa968kEDqSrfxKLxURm
CmqJrNl9AtOFo3QblT2K62h7+h70pGkOjOi3YsDUz3v9G8P6e+aOUMsI4ot/Bccx
3tp/ibEci8Zeb1s0LuB0MEp27mPGlSGRFeCSFfCHJLmk8/ddap+m11TwH66lwr7y
dOKcM3lmylgHbqb62149yXREJIXf478aSPF5pInmybxyIbqcLsVedYxiCCBSX1yt
Jff77a1uBZNU2P9IJi8pzJOpzzqDW39OBBO4ZkNR8eOUWpeLxJ79WUbQlIoXWDHJ
2ST5NeUvexiIZYidmakCJZSpF58VYX9c5gcVik80zFznMOodFJspgKObR1OXTvi8
qWT7MofPrYc4pln65LlaEtXo+1lOSsUZoMuQp+JCp7kyJu+tkLAtTpS94mbEh7Mz
QQp2evnEcFm47X50s74gwJugeFTJRLUp7HsshFl6C5Lt628FWbFtUgAqX0nILb3J
79E5PY4AOtm5yHJypsGIUZOPDLwcYoqRzww0ms+VXDROqmP9xivwtyPtsw8MSrvi
wC/fzcLwtWAz+ZYZMMay3fLt/v4S5YYIrFq4VHgZC2JAM6l/L6QPpe8nw8BwXNL7
zo7k5GvD/VjLIeMURMFFYI0dw9AGPLXHmW7t8VP3Nfzspinr4Z72F3pwajnl5qd3
IzYglK1eW3g23HfNsXcDSMkv4oSubaSn5sBOPsF0gYsM5jFoPm3bPNOQ+HTs4AB4
RUajZo4dWUphjUpTqCGo7+x5RI4lxIuUV7WrxhaBS1eG44P/Z+bVu4B094mR0En6
FIhTsdCWrZ/4M9at+pA7QWJD7b84hO7zoFQhVnx7oBSNt7azQ/KEbbQxFAp0n8Vh
Z6Zna1S4dN1tKg5MkuqvSrVqQJY2rKcpYoyMsRqpt9Ed+4RPS+kwS4QRSe30i3SW
ObS9wAcJcCr/gvvT3bRY9/jFXxDU8yayA2Zw0HZowJCaYkXwbL/cQu4WEZLCZtXC
d7jiopFuMPrFJ1ZYmf2Dya0+4wpOyrkErB2bWaQgRXuk9WLjpApaUc8qTB760im1
7fwUPIz0CdTXAd7zDFeCLX7Ce0I+aL7qs/DJ/oqC6H6UyLNHPUma13ixbnqk9o74
7EJ00ac6YWnlKtZc34ggsn5BVNUfElDnw8wubgUzKEivolHZBI+k5C9FXjwGZWqu
5pSUvN3x03Rd68vxTgoJHjNV5rBIy/dZ24Sl25NYQU3cGKeV57odwB8PXSZ59sAp
OptciDbyEvTxQM4vPp7TKtpZKe8XTE9ZEyTIy7ZPtmd1YmHJFzFIirt47AyV7P1x
XtL9JFpoKqjJiN1ABy+cOHL8g6QVkoEpenk5QgoWzklTs2bT6T8t4polt939vhdN
M2n7LzouX+vJHe73sxS6R4smrLtJPvfTqzAOv1gVUryxcSBIsBmSKhyE0SDUmyqy
WKAUNsSRxw7cpTn7KyPvz8Gxl5qmWetTI6ePQSlJAXVAlKuNEtDvPhpM5stqWAr9
qmcyhxGLbtzDUdXxvLctkWh7M/37+dCpskcsvO+QwkuEsfGsJtH3kkWqgdmQCGOv
12HDlJGKHuNlSCErSxzWVNCADMEj1EPe7Hs3cZmCyiWofolPAw9nDzIhkc8BL+ME
5kjDp4c4cFgZHogFmC7E2IqgAxiwr7ktl2xgNZDHUp4DteTwozAj1E/+quG3NdDW
5tZ+1gkmTsh3xGwCN8Z9OI8GHQesmbpPnjJagXsoE/Zhg9WYoldqRky+pR/fvR2a
QykQ6euskv/AIs7ke6q0lWKMNzXuwGWkMtx3xYhu0KIwntZhHDsb0u/OpT6jZYnv
UxSUstI/XVdvYLhHOCN00t7jE9J7LIXXDLyIKf8hvazZ5JicSLCtVhR8LZzg+xmL
oPxZdZ4ghqyFkmxL75ocj7Xy58aAFmF4PgQjjTXfT9SzJRVnioQvscb2CulRtIwn
ng3bLhZsn+avg+Lc7vJICk6GGZcm3pvoMGkWPtARl8ITcIJuYW/hhz6dDhYtHmgO
QW+ejuWDCynr8rud+Zh4hs3EqVD4jhBMcN4oLLXzzR6kdL3f5uF4ev6jPiAF/ebt
qjGmHKVP65LUao1wANa8LeQN3R1akwwYZRfVVZjCcSiqd1aD1sNszDNQPddnXqlh
nHiSoyS11vUOYDCDVdN/umWqGnPo7rRxZica2TGX5qOOp2Iobr5l8ZvNqi8PpmQI
zKnx+zSAXYBMzOW6hyhEZfJLGTX+iOQ8SP9f9tlsnyfwRtf4Ymw6LJuwjkbvOqeG
d/fgMk8nPqW63ud4Eth3eTgCcwv0BhNYDdifDRqTg3btkgN5hcX8Vqt/AXA0BDhM
BC/KkKp5AuKrlFFkVwgr+ibMPDQh79sOddhGbfWhJ6hjpgraqAoA+9Gx4ZZGaCYr
+8fdfghfYFdZWgkP4HD7corVEN5NiSE3pITJAU1qIxerHd5vVoXP5RrlISn9EvqV
eV4T4wBPDjAMMGmCQx3ai5ZS5FibrQeSE179BkNpBKB4xP7JQK62H/WONtPsc1ru
AEUPpiy7YCkLOSdy9OX5V9fxfsSLgcjpjioCUPxaCmJGvPa43IyB/6GQ/lZ8Q0Wn
pj7yYokOYPdqtJi4Zlaga6rlr6HfyMO+obc5Xy8GJnvgS5W7KcOYPkyA4igoDfW2
CimJOhMB1yGGgXhVVNZhig1MfhN6fI17aEQ/9gdsv1tl0ef/R+6WtIB7cttY0T95
ftU8rrRcNWZCpKbuyE9BhDU8yLCL3iVeEsJJ284+H7p0oMNDatWJxF1Khc8vJ4jD
HEIOECo1huKeMEV0NBzIk27fx4ujvFBP32EVIB23sZ7WWzqMAYZ8ZAozhspTdfFs
PfBOaIpnjaUtjthnVo+E7BKYOhCEb2GMhmTgYvd+vCwyhu6yS32EU4gUggme5kpK
hod9xz7lx5VRzgEYnHqePxyKntfQwRsLqujAh4Z6enPqpYoorFwHYGOLiNvCdrcg
XkKD2UG+TdzMTZQcm/rSRp4esuBKCwmYuPS2ToTv0U2uI97erw+qwQ27qHV4SEdX
71mU5Z7OOVO6cbbuTYj/h0qcvb2KZrNS9thEi/StfyRxNxx2/2BCQK3x1z/fcQEF
XzL30GQHFoGBNFCdZHSIFW0nubE+ghNqA8HyfxoxgCUj5BKPXrFlTNtI5YcLb2+F
Vt8mFEunejB3inuQMnowr4B6d0Wn1t143x1PyKbAdLHWsQE6BUGAONVEAKls19x2
cjxz1UkLYOq3JOdD6oDsdq/ozCFq1H2Vi6qo3aa8HW8YSKyDkkCcgTlTJ7pQyCuC
iMdgiWoyEedeWC+9YPscvbdNT/glXCyQAGDY13jF63IdtALf5IEKUWQAKuZHRs9E
0A5R6dBZB9TK26t3C10yoH9RJI9KS55RDx6gQw7R1WHBBz2OtxDlt/J/IG+sTAOb
WcAYAXB6hb9RtkTDILkbOcKT3Zj6tpKSKJXmTZrScfFHjSqv4Qmev2dSJnmjVubc
rxFzIeBaqlbRzJv/xhIevt6TCsnWm/CbI8tiH0cD7eVguC3UVVrMmHJ6LtQSwWpn
QHD7ivFBiLPk/fsBVzcbB4UvbdsCunxEjsrsKjFOCrnXZX+TKgSLo4yhVmaElteN
lkmGDDTsSwFv6C+ifmWLDn2vXqt8X95R1nlmxFcwejZoCuos/XLIYq9VAhInUgwg
VW953qg5BZm5t7dfRmpFGmN27TVw8FK71AJq3YEluXVquby/lVW1fA4earJoWpLL
aPIh9xSXvmyt6SnusjKT4YfcKB4uUCZ73+MQLOgShStj7qwhsVfIrpcf+ch9iUvk
Ml2qS+TOsH2YhGtvz1BwMX7CLMwAl9sXxTE2PoyoqMGVANagk/XuDwldC3snELEF
TsWC+qxIR94iRdQqLTVSsBD3B0yeOFsMIbUmKXtNR+fOsGGiaqsRGdfDsGNcJYVA
C7shi/P+UC60awN7pVSmYWMyii+oh2xXPBs/EGeh+RXsnrmFZPoLzgwWuKa+ETWb
xraNBqHQ1OORuM4b8U5EDYaWfOVuO7rsMs0NzU8zfF4cbkkzNqwMzLpFNbLtDwGP
BOq9FqvKLJYi1yegtnk0ZQ3QE7xwUDS7qUZHcqGBLwg71D6xZcM3qQMLlGHGdy47
4MNMHVrXOBDTx9G+aIq7oJMyizO9NFHIh8Qjvyj7XfMd4et6zrLAuvwzUfRitIag
qGTnxoy8trn/O228V4fVy/xKHvgruOs3pp1S5MrGDhFVrPMvRpCg9rGTuLoeK0EB
SpFZbc4SmdfHllQlpkOt6I1BAXPjmKSe4aQK9nZNAd/RsqaDoPyJMCid48RvrE7X
5fCfKAMjL7eXOvv93fU19lDm5UifPbwGvRrIf/xqdw/17MrKHIuzLVVyewNyDNe+
Gor2CmS4dhsI07pC4jBbXeP9t+S18Smdoh/SOVXW8WcNiPwR2wSiRGOCeSS3e5Ib
xSv+hBhbuUkWDUFEHpO8gvQjKFjyqUUuCTGAbF1b8OqbipJpCVrKWcZ4b6vBPB/s
4OK1LXfiEDi3TIEilDdf6lyHYhyDIxXVB5beQEJ5ZxqV/IbwX5xxiGftzZybkHx7
QnxA05/ZyB4Mdk4UXx45BWo+2RJdPBx+wQzbbXe6J9blp740dl6hmhfoWz7NVWXP
unOpPRPRuUKBfappT45rRcwKJpOosrUDgn1519p2JKF1MkPbd0BIElGU3l/77xW8
oPvHZ/R/3ojRHSAqBm6w5xbraZ3AZ1WEL74k/Q2GUk/1/+W+EkmZUaLjHl3HUCIu
Obcq8lcpOlUc0DsRkgbfV7QeptjyP1cT/Can2m142Mgr13funxJMHbRG46CWYQ9H
rm7JVNk64nLfCuVXgjr+F0KaPQEZBtIpS0OfNdf8eQ7ygWwyYXbObKoPMa9qfGOQ
bIdzNBISS0Pa2WD0hUEuTrl3PQAGSr7HTWTPHtBirKJwIeati+89CWnTgTDkgmxD
LvEzcJ77l9TsEiGyWdJTDfhyMndXK2BUXHnmjJJHHUlG0+Zvqn9Ap6M9SM2XMvar
W2YtQO0+54AFKPzwEWuR6Q6mJcFwgNkm0n5jonlx6PzNjWy9c5GxpceJ1u3NIYWB
l20TYdHJ7K2xBm6OP6SNBd7ZWkZdtbvedab//QVh1IAjc5AK37kD1Tb8xxh+e4Xa
FzoLF79OTSfoX1Q1OhjhDixSYnv6lv6HGfTFzjYZZ2xzt8ofTsEIQCZ57ePuFC66
NbePhhE4dzqhUnEHrd7XWDwyrzdeyEQdxQlWtD3jhriLta5vQHxOcJa7DC4DuX2D
gEWL8NQ5Czv7zzAcEjlqIxBvZIr1+RElOL6VzTeuV00t7cV6NWqy4mCcW6weD71r
X+djzBXveq/BptpRJAT4kX6sDwChXMjPaHtHoB4qqF9UBp4LJqsZpdefeVkIWEf1
Chj1F5US38WMyMRYp3AQOV8I6R9GA8BnRQseKuxUivfVHR2d1GYhc/PRDlaNuxYu
/y4yO6ABZ8hvg9Y+hv9tXfR9+8LUysvr/V9EG3/KwAXpVUgoxitb4NzFwuMbCqFr
15bW6fhEwrr20QlVKbmv7E+JYEwm7i4N5oSstuJux87MVSwMWwsGG2USpt/w3/3h
aRzesbGuccx+iVJ0uz/QmsdBUJTF78qzgGnPKFGtbZSrWy91rkSfbGLgg6CQqIdI
E6rBhbkonLNukXCF5EJFxYVDjOZB/pFzE9+jsmgzyFa+o5sfqU8WA7ah8mls8LEU
O0h8cWS0tgfWBluatlXioPQfEq6xAdJtqXZgrWSA2dO+tHdb6sBfTaxIm8OxV5pE
L7Lv1uLYPVywucm4idNoEzXfu5OWK1yHL0Dj4R8Im1TmcMamKh6WDQ3LmMGLu8M4
ky9+EORI7J8T7eT1DHV+bgeHMJzBCFJYmgnNBxjbyhPX/6lGgzOltHFVbnlCdq1W
iNOMewc3XKORc/yzcazJTRzIivImnxi/Ts2O6ABwPfHWJ03UxQq8QHWSoOii7dXj
JXnSRvTQlRv5y3OaGYtThFff+2VAt2vzG1S6y2R8j1tRQFINW9pFKGjCuYFqNV9S
88iLLcvpR+YjxUERK52jPkp3XVUcT0ldnjq3kcIWYSIbhzWulUEBuxvk6ilMDtdy
MiBZLrdr3lG/ZRHxsS6PH0UqzYNkpxrIzsXqbkv7yj3qi/nYr2IT0RVrpJZ/jOpo
oV4S9xLp8wYiggZYq78Vq3jDZ9S1gYB672NCLy8PtdwaGLHis6usuPVYOhJDa32S
A1eSssOgsXkNHJ2X6A3QtxSP/S7Am8XR0/c18UTc963t7ohz4AbXqt2dWXFDgcqS
tCNsllHndwXNPtk/NfLxMVT3xclz5wp9mn5/OLNuMQVDlWnNjbP5tv66K+JhyZUf
25rGLhfWtbxl3GhDxa9iA/nwH1rfZxspDN6w3FN59QEkODaiONPw1mVqaMrV2i3d
1RbCjjXtSihSdoH4xnlNqcS6K3gRUApul4JaGDIGbkRbTAMfrS0M2cq+IrMQF7lC
ie9aoHlXfz1KK7OLwiRANWv4z5V4g/9RCNiJt8lSf01L2gtWoievpk7mZsYGnd3x
/UiwCQ9OfIif310ZSo0zFoaOLvkPrLmNWmibpzjvrTzn0zhDEHtKdNWsrhblOPjV
gmaFH26Zmk5gXGbqp7uRr/znwnnUub0sfw907BqOxT98o0AEpRYuy7ecg1Kwvhah
lJuytb1lZ88lU+01SYasVaRvrp6tZ1Q/Lev/wfxuudM5lNgvAq5+bewd3KZG2JRf
p+pfhsd4H4pfQOwWF0/A7HVjFveFCxQRMCAVe/OrauEO2Cr5+4PM7d8RCZIFutRC
f89puAdR+SgsMMaUwpJgtgaE9PBnAjBiJMSkrrYykxlJXOgGQAh/Z94nXyAZoRfJ
UY94gW1AgtfkejSr4RTVFV6+tBkJXzU5rMVpApzc4KuqpGJe5GhLqSmQ0tA6ta6r
mpLbEC4OmwV7OgebEQTbRORFIpUTyHqg4WdSQquLf2NoxnEEKorwUB8hmJlzpbEP
4Br3VbaajwfVlH0OCNKwMoTPlgAYupv7+kHH3Sokxjbgji3tsOJ4ayLP9HhdQ5pD
l+qm0AscYrZWdjim8j0dhSZn5CMYs6iCAfUptucjjVmlyz2C7JbmFj1HdnsF9IwT
8HbzW8kBobwVWfA/Mrtjlue+zn384T2p+hAajec2PDgWrL0k5bfdnyBqqjNtb4Hs
+oAwCBClzdzn6ldISBZ/asB6Zi+dXK5+QgyoTw9lwRf/0PYJIqWNr2UATf1c9J4I
Lh5SmLU2Y7wIPDGan97ARuV5qW9cAraN1QEKfSXFLnLVU8BDSy8F2d6XnbczndFM
GaBSf6L/i2CCnMMabKF358QJn56Mh/4twlC9ClDygDu++ilqn+tEDrMKAOxyZ+mg
+TVxdwlXBXIiEcykoA/zwGbxgiDMlIIbCCyY0zQEcOp8Fwft+NMcFS+m5tBg/gGn
Zw5QA4BrYsUyrLlW1s2gjfuDAgzW7fGdmp/DjJP+5OR1qIf7D9wz2DrIx34/PTW0
c+mMs3XVcY7T10LNptn4jh9SaxlESwzr6Q082T8U0u19NZC7Ki2kyQXRxaabk+p4
9Y3kClq10VK+lOQOuTucPkASEXwzH8FiX5R8GrKloeQzaC8FdGE6U2XSeKHVBVtx
tqgPaPIal7vfklQhLlqxmsyUGLPX2U+cGx/MNCpeJR5f4NuaRG0RDSqJ5NSIUrI0
nZOTPqhwkOVBCu3fa5IBSw0C4AxCZ+Chx3cdudZrwGFHD2iWzHmL2kwSV7MnkLY+
2D45yDkX1YA+Z5PPh3hKyunxSh4O/Su5dJg6CW/g2quUw2YwR63Gmer+PRkBOAMX
AKHy3VsJhIPLomUkZuksxjvYhYDZ77CjXjiTkNSkaeWu9cs7sk80mKSq0Bh0mnU9
NZzWNmPQynYrrKDi2hGDQlaU5EPp9oE/oULWUslK+Q+4xR+d5t3n+mtYylwH3GJL
ps/aTM2fjT8fw8aJn7bkZyoqAbry+hQfiwxuaanHnZAzO4I+p3k2zgma8jV/ugoo
unBIE6HsZk1QMIVOWYxdHkkbptqcM5rIUvAZsMCegmqa9+hbAOOidS2/+FXvCSBQ
Hvg+yDmlXW6LcwgT2Wed2SEgXYw5GyU5VkN09/RmMv24qnLZYyAOx+KmPJNNMIa7
2EtQLMkbEKWRiEpJEJD+P7s1gcNT/ad84aiG8gy5C8x+J1RCsLb/6r+4EI9Czbbw
SNsl4sEwFqEaqF9cjdjEu1wB2zPd9XwvoCnALIHe+m3X4ZbikkIVuhnIwXrCNcb0
kwRHykIdre2jCpovm+KUDZfDZ2w/almbHiYVAVIlsmE791McBfFF72yOoPgGEwII
JO6BTVbUL6ZGnqJAl9oLSIb0twqaUEmL7WNLEcW6j3RmcalFXPLndz0flpzD5Wj8
1Fz3MiqlOG/3h9IMHyFdooqzaBLpHzrEIqJ8lMlT7UnzTpOsqFjOrgYWwxrQozD9
OWKvI8xRZzQ8yskjO8nQIWIDod36pOfCpWe+snI5SS4vhcxU/kkacLngMscMPyUZ
K+Z1HwFpcu/hG7+gLbBCwVUMdTPFPG5W8fLeyxNtrKzsvKmZoP+X87b8uTGEvW0w
2Mtm5nkegckBWi8ulxadYjrQq/PlogSUPu/YBsYaNst2Wcfeiu2uXpjLj0GWay9X
x7bbEiuTQqL3Yo8B11Oa8e71Vq1cT0A2E5754lb980IWICxSZx+4OZ7eOQXZo8Rp
D98CFctaByeaH2oTJQqBjQKt7Mn1rYh6+i7wF1c53y1cEsBZGMO4aY7sZKTuajgp
mz7AebL5HoV9ZrlAI4JCAkVFg422aQYCesNzb4F1xh/BxQEjMOkVU6IMIlwYdj6I
aiqeMnraU4WRRnIhH6pYjcwlLlp/1F6lybvAcG7fJnCkgyUGS6i2n1zi7elc1TKk
pfnayxn5n81nFF5k6WYdGQJ7nmlrvXzmrKZYoLYHMcU/69/2fB7yM5n1AkW28dL7
samtJgO9ts2aGVZ+nWTpbj55me4MV0c+JhKbNTEsd5VH++wkN1leUSnK9smg7O5s
S71dm/1uGjJ0rBje5GDSJMLD5zX3iaHmBN9FM05UNGPOQ0ooRIAf4pRD0KLoO5rq
Z/IPr+IEkoT6zY6SindStyKzg8AeRl2t0e+1tVul4WvLQbme6auzW3DOL3RXPJ5b
o8KaMB9wvUyKf7s9smNLW1pJCSDpPDG5HNp2t2oLwz5CleMRfgRotxH+zi6WVYxW
8LhRHlMVRdqx2jJ2yS2znE4GXxYK66wK5ubpNG8Ww6RKo6SzGA1oQ8390P2YNSA7
UCxyTWsWH/JIROxqITQfjvO/f8UftxiSk9Uy/pp+rgC8EiOLh066Q8+o78v8rXs0
p0wIg5xgosrJb3U9/fL0q8P6upQIWMxujz2hnSTJPReK9B2bzowjm9r5MDIj0hro
A8b4gBvn7q/BOMthUZXXCPnclDDqTNIhyA+9QUxKMkxbXYYFaDcxfnzUt6ZwPxNy
l4k4O6SlbSs8enoMkhiRO/iuHR37cu6mlMgfaW6/1jk0/jyXU7qpxu+4uWvdWP92
Nao47uOmutTUkmKSe8oIbvoGsZ2QCcy16knmyYquCazH6QT+M3tDJ2ha/2jBgwix
znwhsFJOCpSFsFBrhH0ompElD8S/P0+Je8QopBZeGQHP8Mtm2anYDPQszBuFxJ0E
pdblaJL5dV3/wWnDmYdtJtAf+lU7pOL6Gly1J8OYyaUC0ybjatJlOmqNLL4kdtWU
WJMpyO0kxhUDkQBFPJs2NZBgAoye+iX4tk5tdg7F1tyxxqKGCpfK1CCNN6VLmfsb
i26ERuaONHYYcIQsYP3W+iYVq7L1WFW1VRcg1eK3fj0d5cq0wjyqKpPq/D+nKmQN
ge02rtceNq4mCMLyDRSrqp3x0IjQL7mEYRH1sCiGVf6UG95Ps9jDszFCDcqpDFdL
dRt2z09AHhi5ZsUpdoUqmILeLJOqbA8oFgP6bVgDBynUDZRSu11JTeuYiqtxBR99
AbbZv23at9Lv5cQFlw+9RryQGzrxmQ1J0odpJdOH3g89pkeXnLzwDYm+55v/umZ8
8W93mD/IUoCJbX7rQAoinahySbIW/6mA9oUBiI2iMSaq283SympGj/Qy1/V+5ZXf
Pn5576BGUN3e9P0owtpSEs/7E9sX/vTHFDgOdmPTM85lJhnbkuDqUKHodX0UofRr
c/qqUL6vzdrAjgxXZc8P6tXFlxuQKUpVk28Z+oYa6utOHuy73AUQuAAZ/EyktkFD
6IdDvIQbuRe8feyauIAetXHrzOsmRYp0GnVoqh4Ykur7ALa4U/N6jQ18FelByN1s
GzTXuX4Vwn2kFDaXjT40Z/BNIKUKwrQWNK2D5rBixplv/IdyMhOgW6RFFF7T3ueO
3f/Ma9NIZZWiOosAASnRnWKNXc2SaUuZVyneNfRNInp4Y7Ft/ThErs537SNjMX6v
VG2DB5T6fAcKv5FWtqj2Gn7ApEj2FL0hxXF5cILuu/O/MifuhNsDDTBdiHv6GeEy
cpuJQFFNJVCH6vIeQNuoEUDCmYZ+DaoFbXxkybprgXtMi8K2bES4n7y7dRvKOLDA
x+APY8vyhuFgDwrTM9KTdwANBHi21n2gvLWQe+sCVUtgzomAINLcaxmbnYLS/cEC
zIgIfI2J9+y8Xry5kpmbsgOHQ5DN6H6ACDDDRckwraZy1oHAL8GyaPq/Hjq8P5wy
dO2fii+H7AJb0QJEufcgHE9sTYbXpYMlZqMRj9doNd+2Y4eN9n2uwzTN+oPNOJ6N
O7ej9U2EfR6XmZFIS+MnkPFy3FmKOQBmnqXy9CV5RLR1jDHdafl2PwKfV4ue0ywy
jPT9Kij9U2H/Rtp3Klr/s7iqLpzICNjfXtUBxkgwaO5qBLdK24s9mKUWF/kwf9Xy
YtyGFH/DU0rxGKVscyz8Ts+zXXQtHyMGtT5ZmQpslpfyXBcK1blwJbr8LvCgJRlA
hStwyWmi5Mpsit3Lfpc247YNXqlHaHamkrzwERZj8lYMEl6FzUf+eBFoCYeKBiTk
Uw29kEjWm2lslB83JXUZxnImsc0MHkf4b5SiHRZ4KPb8OcKo0UQijNPYF5Mulqlb
+MmGE+p7jvOjf0oq3YyIy1X3KgFwayMrx3mcPusRvX8jV3vf8bw2Cz+5HQw012Im
AbNxQoU9JpOSUKyCPiBMblM/tq1C2m7JQZ+t8oUJDiWTVZc+RRlHtoxkH4JsFzgP
QzhYDXOfftz5RnmUgxNrDARU+6p+U3FfzLeNXptAcTNOnrkBrU/tjuV8TvWWh7AL
t2kzSws/TZ2z2fY5wZoIj1+eHJi3dCprGyOs0+3oeCb4haZydvovw6cNCGYnKbxH
pzZbvoxe7TbscqTub+3wwzTPTt7j+pwdWACg740TNj2npqy+MBAwU/6019PWrcqr
X8xGakzbBUZgiscGjQALaj8PywRMAiyyz9tj+ZbbEfHEN/vO9gLySWNSz0Gh2uYk
Fxs/XZb4UZ4Un3PxFDMn9X6Cwi4JFHVVNx3C4N6AUMYrJ2nRHT7pnSDKa4ovBv05
KrfpzCTiON3cDPLcldZ+i75obCsRSjmy1FfzVmM3KAZ9L/aQuCBrJqAIN1Vh0LR1
qMD4bc05CH5H23/4CRtAhq4pl2msXnUNC6UFsF+tzlkbEpFIm9CN5hgvrNPXo3Dg
97u7dpawYICL6le48ru7V0rnCRE13lDZIZd2NzU/2/grUs4V+mFVm3tJ2xum3x7f
aveKGq7KNb7g44WMJhW3cl0pn5SrshTBho8eE2oWx3l0TnsrJFCb6I3zpdg/2/1r
IS99TwWgECORe1feW2pMAh7vZp+8ygY3+h2yVaU/wtt1tvNLzFvrYRnbQ5Ab4JiR
JqyZPhvQ18PNfWDhBFKieml4O5Y160kaWnDasB2RumloqGfLgyXbIFmO0U0kIgYb
Y3byUZHjpdKQrHVllhZ42Vez8M1f/MDrrKc6Gj2RY5iVUowpZ0R4yYtIWTbiAK8e
IAw8+Fq1AgbHw0nsa75HOSioZWAJEBizvCb3BCNnWkldDEMqTZUg4lIiR2/Orbpp
Ykhd0sjlxAc4snpHKd1iouCnkW0QDF/RgkbYyc6PSf6PDz6kRa2CBzaC4mlxCTgH
EgWYKc4aTF+d7jGCEqE6P5CBdhTt4Zogstu/nFiUP9NjD3NAz77y2dZZoR6hH48q
ds74Yuol4ov5X9kyRIdoEdn6Dj5UtGWNE0fIXi28JbhZhejqOn1liyc0nnEGMIds
qptgvC+rtynxXBSu1zjvpiNNbddF2b5ax0VSL9aCcK/xmfPoXdIuchNLGTtpibW0
aIlIIUdd0iqgmPqMHR8X4X07JoLuaWiVBnXlzcnjIKDLR1UYQwvQpwBSIjYm0j0U
J09FaB1Oxwhax7yJyXIS30casCpVWuoHgsCuV5TCWfVTsezrk7i2fkEjjAR3hCF6
UD9E4NZ/vtUvtyq/c9YDxW3S4FC4c/WUQ8ELN759V2OVozaSigDMwkXrbREVmS0J
Og8OGl+VJG5BY/5ezmKBlOX4E4CWxWwTYYdMY1SOSc/n9szkFg4wEmvxNClmfazP
m8FkYtPdPvY36YvJPRrsTXkZMV8k74+pRCiX4+ta7teN8RYQ3qIIwpXfp+g+/BbO
iPOgjy3drTHysolt59pHTGADNx+LEMyvXBsQKgx6fJrzOJaAlw4aybPBbPucM14x
tD9/ubt71kN7pFgFqwpL4BKeqRBa5IuPxvkIDsgO2Nc5TswC+gjazHE+Qd7IsKua
CPU5y1T8elMEWmX40L9ByffW8D9D/YSGozq5ME6v1so9Tk1dxxRInhXjPbAs1Fnk
rt/uP82OF7flfkLQZNwEVXPx3oM5RNnqNcXJaj1S4j+5mQ03sdvg687YWzenBWw2
F/OXLfcWQY8vmgCKDHTIgsVgM/PMYAAVEKyXmH90v78VBC5yZ4ZHXd5HRck0GBzj
1f1j8YEIdsfbu4ZBqd2tk2jAU3L5klZuzB62zNWx86ZSRYafIo7rJldtcHimkrdk
Lz4xIkGV0xpM+lmbZr8PjTtus9Va+GcKreTqEU4zlHViZllUprHeC9e5wsuwR2EC
1a1BbKKmshsGy4CF5p9MjCCDHqpk7mwJPqol5vyxa5evibxCMZ8to+qbmPGiQ+Ki
INlb9OhTD/zJmAQv7ynXRACs8c8Cw984FeiqQKyyljEHe9T4pDAmncPbj/F/j+1q
u9xepu3mUgF7jJ7qGWGcykROKdUcwh0LQSRAXMnJMudZtV8MzC/yiNv+c6kF9n2Y
5HDOQJ0MQ0swTG+BOqBhoen0S5EE7mLqLCJpVKmteah6MRCwKD9RwDqb6M2CyiIG
Jyf/pZIOdv+G987h1kyxYRHcFtIH45fqpLUk76PslXZf6KiHBETU3hg+zUiFBR2D
/sR5rc4cCYyrFpefLL+/pzaNCdOK4lUyBdEHXJuohj30sRUn1sCHR3fSc5ocRm2d
1NsQjgLZ+X2jzMjn4WCTyuMwqo9r78x0mvf5jNSaj5wYXCJ4iAjxn9zKgsB8TGOr
8tLqKPMsG0X4cr0iXJUOOxqsordaLugaIHhry/diS6yP878uZzfgZl4rI9w73Nu3
2by6GU7h2JkpLD1saRuVb3XXNAnh26Yx0+/3CQVNikF+CQHU+0T8AmqmwovEz2pD
4Kqg6LfGodD8xDF8h/Hqi01+eqJlCS8VPN9uXbp3zQ6e/7ZKd71XJgazgg5Xnq8h
mAwOhD9+mFNaQGKa2mlzi/LKgAwZm7P3o61eUG+Vw/dZUBRsBIdgzcu1MUBDDCGR
YxnNzKRG789ulDeUMdTjTrvHSQb7AXrZ6BFEkRL9ufb06/iOdHSbzkMdlAs/NziZ
d3Luznt+yDtGJscp9piuZTrf4kKghe3zD/UsziOxdPZ2vS9coGZh5LvOX4I91YMd
v7RSGwGeg8Bh9dKFmOohSU6EqKcVUn+HY1pPlrvBt7ciWEVFQvPLdWrFOa136gif
IBbrhhcyKWV6Vmub0tf5/kJDA5WzCAC2RTFx1RLiC6f50rChgBqb+pw9uasq6adI
HhBwU03kxXle83wn3SGUlMrP8ZC1TigDkq2ZnBzwlXVaRSM47o2aGA1SLwtc9qNe
E+U/VsIYgaVHKhpAHbmkFJSwQXNXzxW7mFiSzDpWDPZYDVDfU/ituyWrR12DSTfX
Z715wASyINP2E9V8uOz5MQ0dSvWI/h3gz/cFsRHQ0LHiQ8i0urQU+3yjdBxannqQ
KlZay4SLthpxAWT9mIv2CNsof9bOzKRGQxDqsEWEGIL0obJk2DQq6qLhjSPI+bcr
7Q+Fui4iGTZDy6G5cxLyjFnHjtAPz4y7AGkspGZuyRcuWjJETRJ9uf54X8kt0Dbc
eiYvnzzP6TQWxc5H5bKTYQJ62k98s96vY290PvBd19ScGRnVhzkjAzn5XGu/1pWN
WD3vZQwbqPRvbIAvnU521W+dpNIw15HbRgpXoKJT1oOQz9AfKGpMvYyb6e5i0IxN
2BLgdbsZ0qyh5DgJ9eFotRrgclXjpevU85VovWyoXKQtkqJDqnIzWdte2XBbEmg0
Wr8sYh0jZtaNXAXLmGshiVwXKvoTBrx+/dIG2HG0YDIriJzcOFhw4YDzwzUPXQn8
Nk52mijE6zdJaJN/GOGDX3vzLhM/+11C4h7yagCiiRhmRdCbkgniZU1x//cxuxLZ
Sh9tAT9QKblLKxIhis/uNOhqu04pCSENkfITM5QMGIc0UqITLH55lqFFTStRLCgw
1gHZxpR78Ec/S53VDxzxKwchqb7ZxaoJAv4BF+xGrT198l0kh2/DKRpMDb8+y7Dl
IvucKvVJq0tL+kl6kIU7YhkL567B0qbrRjWGS0B4WVVfoNRuFFCbMTKxpBRDGRRT
Nk3xb9UE6ERI/+50v/m5l4t4MQL+k5IisqsQwYVx8K2cknnqJeOwigoQsn+f5Tzc
EUEqIpRETWvxRmJYwiNQLPN3i9vY+LpB0yRgv2LD7b13ZMrLzPUkPIWHzuayQHqB
u4IOUuEP/fqmpVRdygAGBknY9yRCaOQlQ9AnNTntVkGomAEJD7ocEA9xS66VTQLi
7DYyCG88oCDJhSyBQSnX37NQz9A4v0fmsrtZr6j3+ZawZFa0uiNNx6h1vruK61cw
LIBYGhtxeoIcMRBWeqI6UWrBwwWKCSG6T6dBKla+aHKavIdL0kFChJZ3nPhQaU9c
lSY/5qu5Q+OjTpPY6Ck5/yCNgw5asERgpBZp5T0DdFykErsb3Rgsgr1W/HveejAO
oIbEcFacd5aVbpJNeF5bBEx30tCtwB8FpoJP6GJgqw2earFIQC/KUb60NgqJE7dq
FUdAZATk3oe1ADmFYRii67tcqfu+u/EUzRV8lxOG+Xko76W60IXf+mGVqFA6h6lY
lDolzP+IgsQ0vV0wp2JG54x299nZTYoZfIvigjRfD7QEn5ReOvADv3pzGikjhsz6
ZmXEpsu5pJsQX+lyag/wJ4TzoY90Nm0aGWaevtT/rSRKgZTMAM1NLW7LvlwR2kPL
D3gYPKsTZ/pcCcXGM6aqfcUZFjU3hGYrIcbR55PdPDTKXLSTHeAn32dq8yoBq1Gg
dAfihRRkshvJaZ0q2gFiX7uLCHp/2oJwRB5ryqF83drHA7VJJnsmQN+pToccmRlH
gwlrYLZimsQt8G+zm6ufxrC3z3XagzUgmnzKzMwNFZJxoz6clXE3f4ABThADRaod
HWRYX8QKkCnHJ/NZG/ip6Dq9neLjjZGe5TdoZsgkXJZ9wGzeQ2OOVUeBK0I3vbTB
PgHROMSfxVyVoukW7m7+OHhW/cX9hTMC1G0zu9gvnFZ6nhQyzFfX3f58AGvhkRBN
NN6mydTP0VP/wWskAZqqnzy0Ylq/mwgb77rflAkib5hsWsWrV8+ONM1RFkB2WKIt
6p8cvWisURE8EmgbCTpRfuQvbCYj3H61p5MSuAXxGB7FagqF3LMW22cP2Ie1Lsaz
W4YJZUHjpwlgikrMY9zfVFtn0uvBX6RhyxQp6T6m5qrfsTVPWjSJiVVO6dBc27Qo
YbNmESGGs1+Gq89p18EPNZBo5wlfufBC7JlGh78HYvpIqYz+PSlw8YehZslbPMrc
26EDzZSmiFAwUiXwTzYjSYG7iPEEanH9v2KwAW1j3yT33StBtkWwrKYHJw0BMEct
KldyDF/g3ydH8Gk31iGwWCSxgVWNLdDPVUvyCRxRVPlbkuW2YD1Cvh1k0PMrrIra
Soa11J1uquUfb2lK2SD5L/j9oHMXoFSAVDZ61ToPKKeCvCAcTyFX+lYY4OqRf5Yb
pxCiRCDvMg+IkrwyzHVBCHbNYDwoplhY8SENFviBlfdLtkneOxcFKbdzYLjKjA91
Vm9BOXsmQOB184KOFEpE2fmJDj3GlBe9H2au7zvh1SyukCiUIUChoV6l+iOiNUE3
twCTbfIinX+LtS0MgOuv+1GA154LJ5BsHyv5gcADm+CTu7gdD2ZcTyewpfttVosz
SZyhdZeJf9KmWJfxsJlbVzhDEVQ91kkv2k/1/vXF8lnnGZ5SLBvlZPuHjHR11JFH
5otvMTdbDt2YkcDxsnxp5yPgx0r6Koq2NLzI98koglRCfmiIcg9oQi/3hW0ZEP2E
aeLixmb1uTpyeqxroKK9I5mETX6HzJkXcv2NntnW/FG2yf+MvDmQrqY7UYOq22fY
Pbe3gfuvo+Fg1Jgk6xeDhimAHKk+TcosBXAzO4FjYFHOSVx5UP0cKKc3Z7ru4Iy5
FivIEaB3+bdATw6y5jIxvdtKlV72bf+9P7UPh112m6noEbpvOSmhStG7JcyianPs
kUYtutRoiiPZz+nyaFJ4+S4+Xd5xE8s9znBA5BoqvOhcwoxZD9d+WwlUnUJ1bPcU
BiBzP1ARIj4owTWsDWujiRXdi/SpMYnwqhZ9CAiHSvxJh1iZ9Xf949ZbDDonDBGl
ovrOchBiMHIY6qLppB8Vy3QP4ijOrK0e3t2XLMs+Vfnct+DSdedTn5Dpig9QN4pW
rZHGmw/hLUStZTK0V6r08kUAh4LEqgyj9PK5it8ukCeVkhs+WoO5s8VYaG3e993y
CDYKNeO96rDye/JWGCg0FYl3AY7hpd3sxVQ/9PZukUyx1RAU1bQX8DB1Pnh2nrNq
BbS44aI1i/D/09lJYcgqYFhjgZdJ7eJuriUx3hnhibQ0BbuLwqSfPQFcHdTchPNk
+ExgeqEKxN3o0DQb2LbIo/3DPZ1Atk8UHobg5m9SB1O/B9H8HD+MkG8KP4iI8fTf
NMU40mXloglGMwY8QGYgufHIb9MPKi6i+IVjOZiVJeN/HnEdmrFoiLTCWia/Ufq9
Hi1Y6hqNGCFFdJFrOZv2mZ2BW7vVproV4Tj9X2CqGVQkxe/DtRbYcb8AVCd36jPo
eJmZf45utWtqd5h6FGUG4MjWDH5sBaBthSlpnS0t32GJtVpdspAAcJLmFsPuQdb1
C8rFAzYGKd4SF0DUuBiC3MsqSayE6SgMEyxeMlJhAfJ5gqlOSFRD/Pd0CYsTmKGR
MXGLS3oZlqYYFt/lkH1jqexa2JIMDAgTnsnOHk60riyvyDT0dbCGE5Ie0BrpTFel
L2pe7d6o/gaGzeF63nUIrpA4oohvwSv0q3zZKIExj5Zb2xXBqamxrCBEUTTFeNAt
EOxXrVF4j+FrK0sZ6QASrvivnjHWZoTcz45ZI3uYGho/B1D1jHdB05yLubbRHZfR
JsITDsIqawpW/Ig3mUvMPaMt5RuoW4e2v+MAsw/pIoW5rE2YrUdUEJujn9vtgMd/
XnMAwj9lRbfJsKgar85Mgl/WTJ3wKeqXn9IGM3jvGVeo6gpRqEoBDDHRb5wW/1+e
32/qxgL3t6b3LRNPjQa4P1h/G5f9Hs00cfJPx9F2ImEv0S7b1YAs4usJIO2UYp5y
O77nqxfrzR9mNk0D+NbJw+LT/bLIG7q2ROu8sMfjPEzTJ7jKBDrxw4Ob2t/Q7lfd
GTsSKltncPt5Vp8/E/JuqOL1lxv+ye9AFTpYjVZKZVxbqmllDSFCYkf6eVcnZaqL
LGRI8BGvF/2fPJx7UtwgAnNPuN75HMIDNoh3ODe+TjjQY9g4g75YDslzk7NBi3EP
dXarnOs4YF3556B31WiUwknwq5tAdjiTQIPncqT3HIZroXIhBtBiop8r19M8zHGf
c9XXiagyh0XUINnJebEEY7ge+G2+jsKFKnTn8JpLh9qd4SagbJFrHJx/ks4N6HMp
3nkt4jX6Wx6pKCZpqCySXlnYtK5rtqPUTIYNiEXMZmhQ+kFu3dtv/SBFEQuerHRU
N6K0MzP+ljT11T2CBCkEyQ0QKDvMNmwUJBq4loWg66bHJO1a31BPDNRKQvDNTpy7
pC9s737r5UpUUFM9T6/DCWO09PBD+KnUq4wicsTCDTph+arKrgsS7qAWQ9ArriRh
KTbuguJNN84PVITiWr5ACU0hh5ys4j+XLAdSkwcaP49VKTaYAG9Qm3o5y4/O5OeI
IlPv0PSK18eXiA+gt3yRWD9DxA//QaQQ+WNCcho/x8RI4/Iwu/nd6b2J0LDE78E+
Di/TiEUg5xx6T/WLoR+KyBZMvsu6XSaIPNhNgvV5nnkd0izp5hphLCUJ7c3wOCVy
mfEqZ4dheoLBG2g6ODMUyaOH8KCcVXIUF7zkuLFTrCu48kS6I216IbbrjC07R7wg
FVs2c6A+ynG0YgKVYlPmsG6mvGTNAGQAts7UrRQrbLMI8h64FCe8lxTk1DTquY39
pOkERPd1EZxfn5a5ReEp3SI8JhhWXPZ7MctyohaEJK8ekp+y507eC7mPKdA645If
dIZEiZy7Fi2C3u667W1yeBfweNLNo7C57jDnBy5Q+dcLwRoHiOMRRg013iFMrDjx
Xu5HwEaU3zCjst6+UY8ETFlOu2SMV6vUmcGG8wQQuY9J0PrTfgKOT0DryqY7rPY+
nvZBxCyn3ofg5kYDE9uMQvhkF3VmVnCs8DaIgX5y29QJwTzMHkkbbkrnoevf2Kma
OUdWnbJ/MzAcupBoC2AJw5KtARAMSHi0FoOSoRVH/TpPP7Xy3nX9ke3RbEahzJvx
kNfCiwR/65Lwm764cZrABirguPbPTji+QFLd+oyMYF9stoE+ZWGq/og4KKRmPhvD
MxGC8Dsl3xMp25qJYGYJHIS4CBEvgqvGMimaAdCDTpyPlGPLLi48copxzp/uXXRw
tSay38JgdhCpGp8gNUz0jR6tSgUoawgIKhoPfw+cKCj24jw1dmHBMKICuz3ev+RV
dOM5hhZ1gKQJqYrZRsHnpKGnyyWQWKVpqRN8nvRfZsZ6sFME+6mkOiVAjstVJUuu
Mm6nuFJK3xKDlDVC5fob7hNomDnHMGeXs+tWpy25Rb0J3Oe+XEXgXy6vc4vAOpZU
BPKfVoTW2SqGjClpOkKNW4tGsNkRRgjJluQZmZhvi/lYOR244Nk8ui/4YORYr4HA
+LZdb2+Etu4Wzy/fuOCA0STLhzDH0DDCLEanJ3/etPObeafq9kadte40jycyJfcX
yfr/Wl2eOH8Q7VbgNEOPdkGUesdqNLywJpU7ucB/inCnXYm63W8UnAARE33ZdlWJ
OPbQtOMynFjhXATAUMBvhuBVerOsk3aOc/dT7ui80KfJNBWGjfuCm1T0GAqCvUIl
CgqvYDLfe4S7DO2MHtrd7XzwJufEh36leB1QIQBlFVipDK17voGYrh2WuSH193pH
C8nZVkNauVEho1gJd9KqcWg46WVaJ8k90lSFhl4c8Adgu+S5Ka8G9LJ5HSY766Lg
ZwgYieITPMnIW/8jH15kSZ0NmwQ5ygLxUuRaw7kGFpXHnJNTtWxFn5r2TwQZW1ms
8WPxfhUkZy1dr+LoAdM+BgO0MWy+IhHXbeQrOB2bYqy4FJ3w0yW3/MI4CP5buvl4
3XMfEFcB0zaiBJSBP7E83rfyKdB7w10IKDLuHW8fQjubCw1FOvxmuVBVx/2w8Cla
XeXKUG8MLWCCHmYjBRhHy+Co0iojs86Q8mEv970IvlSixTZGlAJolj1fZBK6+UKD
uXXpIolcl+ytsuGpNXvmJTSRSYXNSGp3cIoQhFJRSAk9AvTK3XX8IBWAz6eYnVTH
URtVqkFXtXJ/dHB12W7xrPE6TmW+YZShesEQl2RSnfReiw+hXxoKhzUO1s55jHt6
DG+MsIiV51PGsjBdrhuYBA/oQoniDgZpwtCysKsZ5hWLW9b5C29qLB5+gJFNE9Pn
t1MTQjNkAq8pju1HuG5HX8SkajgJ8Mz5O1NdAaucILkyo1ue8k5wAtCp1VOz6BmT
md6FoDfqzFXUo2gFnvHO8mCccs+6wzgIIpJiv8DWerlt+Z7yHdct9HoJjSLDbWba
5TIm2iC8Fhs45+El9DVPwdF6xA0aww1kMSzsOdMaJ+T+1x1hdOx65HZeXsWvwTmz
lWt9oOeUkt8+Az3jgJieXwGit1Mrtk+TVqP8dHd6kh3ZyXojjU+9WXJjFoWgoecA
om0FFEh88vqnsmRm3lajpRTO7xKpMVSYK3zMCXYdqTzYjbID2otrfX1oZti+X4ez
D9alXFSqBqV4mGnPOtV4wkGUSULh+K36YvIGymmoTqbNKQakxXjvbISPGOR0tCTI
R+iWP+l/2M9raLW8mTYOIopNd0uLfetFUtI0p7Ndxoedp99eFVPsRL1EO9Uvr3Rg
Sg62s1PBBUv1qEJscNqzavY50LZ0EFDrkqTPKHURe9TM+zwkVaP3//aHqVPcgZQJ
9PgH19nLsko3Sl4W0U6oPw0MF4XAQpMsa5mL/ToG1nMlgoAx4+WnS4EWPf2rgO/0
0OnnPK2QcDgoJyrPZyX2fkEzaXYyZumHoe3pB92rz2Uuz0x/cHuinF7cG1ybZWnl
RYDkmUx5h23LsNCzjFJuze06QTdKfhXkinPPmu3OkOjChhZHvvPgOkycjdVkGJ1u
/ksO3CBp9EYVRtw96P04sgdRlxpULsG/Z0uKcP1RrV5aUiRM+6YjLGZdvwSW7SAi
m4+aY78y7c4jjJvQzrCLYedfyIyizWWEWvCxEiBmWtepbROCcNNefKWxmV9xE6Kh
aDGOaipGnCBsIDG8yMsywFc45b2nDNQXwgF+A2opUsHG8CPtgcMEoxUTwtFRzIvR
4C27MwG8HpVbzX1w9nu7iVqNGkB95zfL3MPf07vW059BoCE1HglQFkHh73Xi3zmR
/l4JyCGvxH+qMOe1nvsPxdH3NYlsvSm9XxNNsMhrKkOP2VmDh6VNJ/1ekNAbdGOI
adCHYNOPlWzo8ha8/p2le+hSLcGkyi1/zFbNIB86DMl/lYg7Rwr2syQOMSxQ2/wh
tAq6/a69AGYJDlIvag4jB2MWpg4XswpCvZwIBYPoxTRSLxaBqYKODavKiQwCIGVB
BWJrXyvoG37M+Mo3z1caRiqJL7l9QGUiQCT9IbYCze6nImCzcvy9rxZ6FsU11JRh
YLS3/Hz5DGLeKAX8jCCzCcJT7l0ClYVRgaRb1OVXScyXDr5RDyrzi3/RXWEI3TYw
wzM2EX1DPq6ALruZBR6UYxmMhzHMmwExOd5Wvqsr4yq+m83Wh5tY6MUwort95xWz
6uf+PDWkZ+oWTZxbLJXMr5B7o1NbSBU0ECKhtQmb0A07HU94dfkBP9slJr8ycO/5
VuMZypVnr6UHCrSXRvzJADDfIrwVprIm0Hf4KuRfN2zulVe6QwIDKoxtTB857Z4X
S+M2eL6yVlQ3denbD+Ra/hRMwNFhlXlON0K/FCjDwTcx8Wb1OeqW+eR3Ozfyohqj
DimH/MWYylKEwdiA3WqUmCK7wLbqLCzA/gfr2zWDUhrxdheYtsAy4zWB+X/v7W6n
43jISnSPoL/pnTPXvU2pz1KVqUB6ly3zxUlqNRz9nyKzO689Lxq3Lfz5lO137UZY
sZmjTXpl5WYZZiTQGqSVcINQpK2Fq1Utbc5ZsNfUsUlD5j2ZF1INXV/JpUjURR5w
Mc7MtS1M7BdxF27nALdj4zDoGwQ//hcNTKgL8uoyvxeT8JUaIiZEi6wfX1xZ/dlJ
kWeaCF3UwR3ALEcziN8LtdyAJ++ZFPbfmfHjDjkTHTpuCHaV8zZwfHH/tPSidgtl
MdywgIZiXs56qyeIepIYBlYDyIohCDaUoltSNLimBmUeo3chu0mbaf4G3hm5QZqA
Ac4zDubGtU8IaOyvm1Z69gP9B35oCEko/Wz/NbJILpctZeBe4Ya1xCNsikIRu4sj
c+Ccz4u/SkpKP4oRnKSP8ssZa3ecnvJihLcjdwfsEPndjNMoQxbwduA2UBBE4Nbu
+0aHq5l8JcmIApzgpA6A0xT9Qtqa/+ZOAQ8hXzLK+yFmqQphV6hq58qGMEnIovwB
xY706x41oIa95HO5jHekVexlKlbv3TkIjZ1O+zI2hXKr4Sh5iFnmjA9GA8UuRKUa
bQZIRnSREITnFO91ID+kPdN2svBb73khKCdfunTycBUqHKQutmZ36kuCcrU7cXHo
hBA2vmRbOZoYVWrdYfOfrwppJgbc/ZtOJJd6DgXkCdvY3yNToN/QHR5CI0PRAQkX
rOb25YhB0I45sKwybs6KSwNM0gQbvvXIpveE/pFNVDd57zpOvZ2NRWDqFEhodozK
qp9ba+Kmd1aISug7dkQsWFBZcH6WQaJEB4YDNp1ZGGJU+d+LJSWSXUNsvKowb2a+
UImKGmtYc7dSuM5QVPBhE2wTP8/PDyH88yeM1F+aN0O4rgyu+33wat7NUGDrqJcF
Wp5VePyfJ3Ara+xGs25pYAHlZGXpIyvgGPYwhBhKTvlissFMBEs5cs0xoiLnReO0
DgveZe4mpZEOWmq7bVXexrsEVOyKUTPtiOKZutJ8KU6RWxf7S3HpQYCdkVT0JAEE
GT8l7QHLozlTVPU4qcIe4wh6mjkAfh5HdxCM5a0EhQiDDgIRt8NQej+w1Q/pznBs
POuk6UBzM0hJs5OESuTpfB+nc/VexfooxLuGW/m5t9X+K8jFYU8W7c+Fnm2uYHXc
1Y6r6bRsaBGdn+Bt4/EOL3J0fNjdkAX9hLe7dn4I8+ONmd36MmC1ypU09LGIUuUa
jFT8j0WRXboFhvKPFFJYDYWeppTssnKRDbiFa4/J86g3RFlTJWzDULoeSAbg00i9
xMvUduqAZrcYVUoC/0IhQ4KQyzcGLr4b0palPhSU0b4ZBfXBghDxnT9o0BNewPSU
1GWbzvhbfVB8KbuydAWzWIZSnpootkau6xu94+c9ZMeLGuL5SQ1myGbqNM0tvoAR
3n2QKvxhIc1MzJ9SDMf49wPfvJL4Wgh/AdtGFuzbljgqnNfD21Kc5B1BghZue6Ft
z9/uGhVglpvqL6aFWcYX4SZEhKUvozGxvWS3ic0QO/V4avqZproJA9qRrgg+efK4
tFRXCRLiKuYJSLaWURwXr7Avjq6vs7nkW7jTAXvaYp3rPE/eBe3j1g+ALPLtEbow
U+3oA/L7Zm4GyoG/6217Sg9nf7cuvDEnxpQRPBWHa8waCS/AbOIsYceaA3xTbMVF
2fFMB5uxRl02rezBZ0y98cqEM6Z3R7X6XFx/oNPVo5TKVUSmBfXe3zoy7FvapLXu
4lqWmTcXWQpN0HI5HBhUGNxhwok0mUAfqRBCKIOfs9fG0a+hbvkA7kCzVTpz6e81
Vsu/xCllvlMonXqNmj5fQUwy7P4FUPcZz0n37TN7Qv54QbwJEbHwtUZsnpAjUGMD
2DJHDxlY//Qd5x+hq8IRdKSVWdNE2H8btu7h1kvF1HgcDcbEml1gYSNmhZZtoFQx
NWVrrwGQG8hkSPfVgnLICuHekqJZ4CHXQghob8zu6vDE45HIj4IcyCsZpwORl75r
d178bCfzCG8CUTBGWWWWS3Tolxcl8vNpBRJwG535qkDYYHK3YWp+4H2zoc4J5TtP
DwHpNpk0J3TnNNNKNmXYV3meFdG/PrGSikYr620JRpVLxFPBGtDHI/trs/+A3i66
VVEL282IkYC0/7xIWce4hSMvZ2Ief1kasbXikzAcry+/n4oL1+n4dezUkahxGZOn
58CRAckLLj/RRM4AYiDMETbWjRuoIMhgi4nRp741D5dcTdabo+TsSooF44HxqXI8
npDo/gNUHzKVGUw0Qvx2yZABqrQztkkL4wudYD5vaciLaRszhf4xY+ml5Sxg46ha
gN9I5xl9cH065Vw+e/wiBBhpXA0sSI3UyVhoheiO5+xZ7WoxTU2UngE167vOL9Z8
Xn/gME8pk0bfX+3la637mdyQ28jBd2EVTaaftNU5S1tPqz2h/q4LbBMHtByfDOoQ
x9c2XBFltXIxyC4H6oNzz1vM8USSUtDNg4YdB8o6Z7DkQWRvSbHYLlJugS4aeaHJ
SphsEzpJQQOsg0/HS+5an0oJK4kE+NFuS109j4LVDTEOr8NF4NHkLsiuNSPtAkV7
e3WIK/i0oSW6Z+4937xzUHAqDXwwVy+gIPhl6bsrEHgfijKeSHTXzHJwWTdsFKQC
YX1ZQkzug/zo00Z1ue+iesOW0OnLfdOpJX8qeYYVMRYKyaj3hpqXK5hXvFZE0lHt
n9e5UL8xsQ5wOWySJjs0GxUlTb89VyxOqo7SDo5JaLw3gnpXMo20JCkU8qi3dbbH
u9xmf3Qeo9ia2IQ4U3qbolhtnXo1XJLi+Te9DIJc7tI6mO0MK3nhwAMo0T/ackHO
KAONrwledM9z7NiXffgfO3LnsIGv/bquYCoQHiN5SuVZyxw4YkW78NaQXXMnR6jW
Tl2TkB8utsNEkBLPBno/vGy6uvgQQH/1UM90BVZ3xyAfGhMIxUTaaclGtFUsYmtj
aCUYiO2AK5bAQ/Deq7rdGrMNDTjUXLVqUsnyc3ckhms5mi+MyWRgGNPkrkVvfdyd
PY6Y4Jz1s2THOlUiyiskJYe4tIVPql5C8NBaAvttwWNvJdSF2YrcGKLFBCKwb1Qh
J3EAFAOxuKUljPbqqyW19rcWAF0M4CG1e6EyfDuaGGBTLf8O7bG4EiTuHhe39GjQ
CTQYjuhT1DxCMnqMj+w0RKSE2qtw5ln942uPqwFTyD51kpYfg3J21dgDrFa2fCiP
zm5cScTvwCH87n6IvoCgFKAWzi59Aq4Ie1Tg6y2nXSDOhkQKPCTXJmp+SwzcUP0N
WxkjX5JTtb02kllHfKqhj+clEXdtl/HNAoTbmzbUmF6BH9oYsQCX0jdEEbU15Jt8
SnTJXmOIP0yMyuZSqxlb8eO4E5LvYJXW+vtMJ/lvOeDTJxomK+GKd0N5IvMX4Jue
pENusOnR4+xdB26atcXo/5M9GhoEa/NbFCuPHARr4LtpE453uQqesMwLZC8OAsDU
0ltH3THI0Gkobe0ON9VH63egUqEu3TzaLFE0UTX9vAyljdRXzqkdq9Ghrr9czea9
lrJSL29QJueeyDSWnKi53sE7QxRmPHc1mR8I3TKuO/rLCGysMpNvBNmam8DTvJ5B
cf8XHLO25VBYagAHotidp1tqLjnviKrS4bBLCoWctfj9y5Vmtfg98XxzrWGRHKZT
lW6CkI+XoSlfdbXm5IBR+p5iQ8E2w8QugGqQC6SQvKnLBFmxvBAg5AB7t7w/+P2q
EIBZORPBGw+op+JdGpVC+pWCRIqlnKxGXZGv4NqDuYc9fekAoeruoJ300lL3jIw8
dOFv8Y2I7mUDgkG96OPhgVDOyfkyhRVmKnk2+0GTt6cBdeQbOp2UBtdrXAafJqWb
UYtIAU4YpcRGG/drE+1J2O+8MJx16d5hpNpjtt65rvUK8js6AgMpd5i9aWasKYcR
DKRqxuWGBoiW2sgno+MY+q/9YFPs7A5l6B+kKmAQe3wtoRViV84aHRvQt8XgZyse
wuKnA/k7UqZ33ZXqYrOlceToDQNnCTb1w9SoqccaBmkLCZPu0xaq6moGtxev/50i
tpE21FTR7Wj4Xsz1c+CXGsDQcUQCGqL6yk+CVN5ITEVa4tayyZQc3E6UtraMwma9
kna4hw1qgYzdGJ9d+PFhKQqZoyyHpwsefcjgj5digwL46TaPVbo2e8NrgTc9Kvw9
epaxV+/vzYPINvCbca8UQTh8Z9hX7B+MKl7oZAPb/s2Cep9VFOKMRDxSTThPmP5P
LZgCf5NMK2/OswgnqHriuDK1ZRqEmOSF4lu+qqfqrIgv5jaPZFKNfodK6BzTFb2G
z/RLJDg4MT2uKGyfaGL1twpC5tTE60WDJufgLDOUzUW2X6rQqSKfUOUP50M+/vPd
hL8um2UlHP6wRcQ2BFjE+lh5qEusF8Ar/VPFs3pLEgiSuejh7nobdAn1RiGvhcVe
vD1ShtT4Sfqig9DFB5VZfrTZYZNXI0pROiQR96H2jPrRwv6r9Fl2bvlgW2PJynRr
x5aM6ovJAver0zCxZnwzpc51Ve6rlMQk1km6wW9q83Z0jMnEiGD9FvZahRbF5et+
XJAjVvIQ79kheAIRnOWLwSWNnFayhFquel/M5AxUv1LBTgPsLebk/MR5b1JVCEhp
FXVtOQVJsSthGIyJKEvJlnkrYkujEdAxemHI0NHX0n2tQYyYUMYocoDe7kEMDpex
ViYCjMecHfNZZoRUCEnb/MEiXgLkPvY2RFaKxiRtBKuY+3g3WgpW3/wwH64dNr9H
ySb5ri1NASVPIfxNkz4bczt2P6Eu7y73XE8CkjMEVwc5Hj6Cq4EtSnp9TuuWalYu
UcD2+DQS8akOPzX/RcMfwq4iUf5ayKChvHrv866wDB3x6ocvRWLeps1oADnMa42C
Odi6cdzyazo964S3eSgrunCZqvKg0qZoMg3wzkx3AUvznvoHfpOflVjhwiC0PnZH
zbtM9/9cX7JPx7ioa7d02vqdIeQkxiXdkuLlXA2G++l3Er8GwpbOpGmELYTDeXsq
07t4ef1Y2WEn1Wx+sL/f1AePrrmw/2dLs6/CUUT2WS0SZM1NJMn46IflHhzPwDo2
5oymK4R3/tQqUPjImqzuYLGRgpgS8woZZQ1Yb+GQngzGHcNASnYWF/VQa+QPXHiN
k7J8ZIpbr0N/OnY6umR2+WSRHY7FzVXxv83gEYEhQJ+8GSqTzFVGHI+Yc8OyAywR
hm4bpvu5zjXSROp3UYQoE1TfIQbTceN7OOxjs7A3zijW77qpCiM+NJ4tB/h95oxf
qZtNsz+fFs0q5BPXN6A8PevJSDJjJXJCU6A3L9cBmhoUlkjdCpQS6xnf2F1MWSli
ZG6amqVyGpXZJ9Nyd2EBBNaf7HPTeLta6zhErOmsPq2hf3XSge7cHuN6f/sonaA/
NgEvkMxZ4wfCijzLj2MITXdeYdCM2Wk4YTCN+QTwZc6Jtia94OKRrOz5HYthO2yf
RwqoZx6/c7lg/CAjeqI2cnYq8PkRieFj3+xpYlImWqVjQp6F3P3lY0uZXWq9GyWf
II8eXupbr23YZqIMwiQQo7x1na7VkuLmT7/szgPG//hqn9WWo5NuHpKT2la6yaJc
H0Sg4HYa9jq/C5TdaJVOUiwxxydDBjRdU0Tnp2uSw3F6qGxkFU0pvUzYL2dbZ+FC
Jwbm4YENGn8fmahtOE8/Wrwhwaxg3lyKt4riS46TN7Eb/SLcZVnMti7fUP1ox7bT
nzM+yy8FuENFigr/zuqZxcNYKUr9kA1Lh84V9eDQQ8aQqaX5KUpoe/LGMrvaX2Ih
lOT8Nx1mla+5BPBW+OrpzxNwaweKDyKAuOhc6a/CoBBoUb3WySSyXVdrXO/S1NKS
xHhsuPficdQSzPPeIDY0eIsPxB+dRJ03wmmtxN90e91ThvigCKUY3IU9tifwCz76
6ZIflKIc47qfsoWy+6fXX5sh3y5NEM6j8KRCq4vhEr7PgxfuUAjOPBMRk9wsfbp7
fEB/Ds3YGb4oKCb6EmPwybN+M0il5X1M+mH03oDwXd0hArFjGTqtIj4i/7I5Yx+J
fWU+hchJDSrDc4H/HBOQLS1b3pTk5x9ACVs5eYsseqoLHEv/y0OnK5ecnsAKFUJx
VYciSM/XK+OH6a5Kr4Tpk+DgFwM6gUQykEd4GG7bAcPfJIvPG7rSwGiT6zJCQvuz
5l0SFR11Ul0co0mcOOMztAaW9ad/VUpLRjXZug43jsjRe/pq/+StY2ZGxPX1JuZa
EequlPyVm+dymnVzC7W00hJHrjgFFBmRZvNLFWavUgUwpfAGxLV42blHb+X3Ns3t
sWE896T9AjBQaRHhvkVwgo/+Q/3izPQgo2Dju4hXy/NJUgS37XG7Tm1j4PJfvoPt
Ctw7hz3gQbgs9hnIqb9ivdMhf1VD+AiRKHUtABMo/x97Js2lRnEeeN1mHYuaL4oe
3m5ivzP27rATzyls7eUGfSb/i0sX5hBGZOjrRJwUqMcNFpQjFT/FlM/j+xQq6KVU
2amtz6gvVGHXERcrygRKous7ozNYVgZfY9HeKOle38hXWzZiscEam0Bwjb7OE/no
FeXW44MnGehTIuSmV3ffZNzJ0RMLTeWU6TLGizON+KE+BZU6p0dlHrFT+/NkC2+Z
B60rFBBTHCV6J6kRu75+jR1JgEsbrS2dHqgaBERgbM1BCF2yGaSQbWpchq72Bjhq
pk9V76/yagE8HWlbwzZEKErq6LX4OOKV9MTeYjzwkkKEV7tJLzoVXwLrP9mdMkIb
JaSyV+IHfVzFvCd67bvprBCw3eN4Uc00uSltf8iWkabOhWYwheGoXZkXLKqLltIQ
1OGXZwcjFImmEK2M7vtxbWhMejQrf9wLaXZJ3BMnmv5O43WPcBj2TAs2gjaR87Vo
4ng64jGfaWTIin//30pe52h8Q9XSMR6AVi3QZbePrLt2EjOUgHfaNFWiq3zXeLI1
qDYlgS0oA+p2Acoxp5coAsK2BVltN2gPtL+55Q0VXTF/H3YaSkOrYgdGkjCUkc7m
0Qj8VFK6iF0vUR017wL3jAPxf9QOj2AbzmVaJuEYuKZ32mcnV99YadDLHc8+IZpc
7iBEdedq/KaKWmRbKQf0Z762Zy3AwlsuLU5roj0wSxPLHfNP3x4oQTtjFWlEu99P
m8ahD1DNO10F689b2LkKk5l0pQpYgPX3uxnZiiiTFzeCmk+R4IT+434EkG+Zmbae
4wWSMlYXeePPSSBRJzJXTYtiqXtPwpsq+no/NV1qWwvKH6POALk1gzpwIlbZcu1h
W2qTcqHKPv+H5dYmsielTInpZ/tXPLlBfKc8VeurreIc/gVnmjtMjSFcpkwqU5Wo
0YBzcZ8jSAzqC6XXxYU5Jx+4M9d4ZBKFOtHL8OfSzhavM+ZzL56hUJdkMG6t9Drs
TnEGvF1c/C15sEVCTwHl3wqY0xpfYpgm1iIJKwM1r1dyEmbUG4xxMXtLMQNrB5ec
Q+JPZpb7K8YOCu9d7NmurOmY5CwVNTO1fHVwCMKRb7a0MQB6SpC2WXz4IiO2nOwU
FIgFsSUYSH521EaFGANzZ1lorOeNnyQtS+5ejpNoPcNd3aMBzU8d7cVBbv78B+/H
yZ4RSWi7IkYPcU25/SGE7mYxvPpRQA7GHLqdTvtrysmlw3hs189C59J50TPiT6gC
chymiN/Xf85EKysCWkwg6QRWuD4l8sLomw3FNmJkMP7dyFoOvfiqG1IoFu+89L+X
y6YJvgd1o+6PoSuhRVcov6gYNxrDTiXLJ22sNW/VX328tADzUeNTrMzgS5G/zFDH
hnmXoStrQZEVpDk8egT47WnV+BOi9LVY2rlZn3V7nTnpuW+VuRtWPzd+JLp1sjB/
/nCVX8yF6Vup+L1jOMmxULgjXonAzbiC/kNb0zEKtG2LTka7fQ/nesSpDaOD4POn
XmCJIsjDY14VZagktzfbK0CcOPxSwxo11m6rnfkim6YZsegjZH23ZCVuBA42sRks
etuw3iaHPEIxevPvyWb/Voh2jFwPWxgJF9jDgiUDLqVABFMkoHp1XM3ZgaAa3HUM
Y1lp/Yu1l/YmrUGeOTl6gP48/HtTOdVbx9xgQVII/IrXxMWN/lcrTn+9mZdgDDvJ
uMdjtp0Q/CHYJStWfVNhOHN5eTWMoRy8T9nGJhkUn+21A3l7q9jZ2AJc6O+4DOA9
R/Bt4RUaaaxUu5GClDbSXLC+/H/wCITeRUC7qCitjzUze3N8A1TWHQpQNBPumBjN
PLw96LEDfDrFotSl8AEhu65fk7ur9XSySOPezH6NoewKVWeFs7tz2vtwC5PD2wYy
RT2rx/ylmXwUZFfH4wc0KHclQn2mjn5wrLTyUvz+eKJuIH7YvC/zFMoE8ilVyO9G
7u9Om5kUnt1+z1WyAGbAGHwDFLklt50Qx2ealUxa4lMbD+A0k6Fzfh67HbUug9IM
z0JXK8y46yJbbqeuDPSuyFF9+TGQfBZr/3MOdvZvHB5hLXKBy7zWUjHkcnUhCgGh
gJo2gj6USS79u4njV3UykObPrX9IBPz/1GAV+6FvBTK5NtJbtjnJ+Mg7w+YFsxsm
eGvvCSITrvXbyzxmvdmHK2Evvd0ouxnfN9SqbnuE/vbzBJYFJyhAHyo58c0CkxAW
+jnvy84u//5ODISa3pOL9huSMD1XuGzse0bLCQWGqnkp2r/s8/cRBGSHeWvVKFH2
LpmyoNCqX/2c2QIG86Q6q60VV3WVrLe9pvGzqRIO0YlrJsBqLay+r1qxTRyRFVRX
waUCwPxgOOQqOG3laowwFGDptEWHZXXCKf+t5bIMLj2ZOKw1E0UsH/fSm9Y7KpxJ
nm8j1eM8BgoGsSb51sU9UnVi88ua3uafSSS1M07klBXiZi+iKILxeR3UBFsS/NOW
UynvxvlYDyFpNWP9PsIE1jZCEkYNFSS9+17CD6LDX12iF0TtcvkIGId3t08b8v9m
JPoBPy00d2j0XRdNmlAlfiW0Cc5s/BPTtQHWlrBg68X8DApbOC4fL1VtRLD4LaAl
lELRpOD+4tz4DxF7csaKf+BRPkrr7GIteZIDVjRO7W6RKRDAcy+PH5b84OciUDr0
yx0d9G8m5z6jeBlVqi/ob5KY0xGpNOPjFcWBLgMRw1dUSxbtBTDaCtcOYVKqRlFb
HiiiS69oz380s0PozsUNEsm4DA/FLXx8FiOXfMV6v7PshJg0mORZA4Ifn3KogNhj
JqLx/ClJb4RLs+l/tMK90NRdhHhhRwWaAV3zkw3Mpyeupk84Uj53dDKMtdu3F7h+
d3PHOxxHUzwDwwapPFaOiuO6JEPW4lyMiViQoSVM5ETscbpNqL+m1Ml+Hk3AdmfP
7Xii8rg6CvTk6gNshNBkpH2fd3CRVLamGWq7aHTQjkgCIlEXIL5zsKFumjZiicv6
dmvx1o3EMkQmDMRZztzulBrPtJrRjTm+wZ7C16Ha1tnlaC8PZiDgh+EObiLRce28
mdpRhbNbSZ9/BYtmCj8mXzPMD0461tomjaK0MmhjwwX7ESL3rBoLc2w76ydqaVUM
XheOzqTqGOGMmA7GMJrTdLCKlOYTge2vXXzCEqRjeSYmcSxp+3wUEOgaOBcHfj2P
B4XhIkKFLDr6H128aOP/Lf2M8fzVNPwpODc0CIA2mUonSOcpcKs2S9N9+JA9qcHY
SNLpDfcwibXgVAEQ2WARN2gPat8K8S4WgE3B3AblKwh2+UUMXwLZTaQQIHNtKghn
h30EIGolQpoVBAM/kQtjnULB4/ctPR2Olwpw2/HjZs9dRZuwhNd8ob1d3FeQH1am
Bt55ms4ZuttlGbkYocPSLD6jOl/GkIRGb2++CPTMwIJGzsiMspsj55yM0qxyu03Y
fZWIys4jnWkjcfZCUh2+UP3clfbLWBU17AuydU8ljkivpEbWa+LPq+BjJ53n+DEl
mUIyrTbxwUR8BkNFvT24Z9d5zNWjcIZtBFOiZYbjkhir6sJcMI+t9Y1LQ1RbUh0Q
+GF9bfVlEGKhy6X4cYxRKvqxr8YF4wXbnqyYm+jiREW4+V5Vh8amCHRgGUyJVCdW
Zv7vX7hq6sjaX/3I/EXAf/P73k7V0t+rBNBJshvx5P2+2mBYijcDtjoe2BiblmBa
k6awNiV554vbzAJ34N+I1OvJw1DmOp7JRnsgoweIxHveSNRRxuD8fhKcQtFc0B7a
8jEjHje8LfA2DUcEZ5GYfTM7qdxcDbikkC8A1SupvTd4wR/LpA77ZEqra8pfVtSf
a/2/1QsbWN5RRuhwTSgP75aG/Qx+6ysqB/3Ga2wYVzw681p7Kr6Pnb7yeOFdKfXH
nTeuOdv7OQ/8FyjFVqsWGdjIX7pzAVsNQJNuX1R3ijb3gdlizd1/MWGnm8Ec+oHY
lPtfOL4JGwSsCYomg2ZT1GaNWrDK7Nkigf90Im8Un4jmcevZ0ikRfFdJu281G/0h
ErkmODWh57xQPp3O744UE/mMtWwcHZ7D4iFcOizkHyzo5AEcMjR37PX53Hj0jE9G
NFK9vf8to5YIrcI01+6dswyrC3C+MFf4vK25CzvXm5NaO+xtQ++WO6Z/IkeLJBTi
MqeWyR3A/4KUn3HpJW76kmGQezNbVd3fBoNBSvv1NwhkWB653zhNQJIk4PHOHtvn
zzJonx5RLVUEUHBXdB9rgem+xzUWKg2DZgFOGd3KmDK/IUA7j9NNoTrYSY0Ex7aq
WZPtgSfdSEFn7yLWCXaSLQ+HVExVeeFCv0W61xzgxR8g/PyVvmVY6zSGqTnPVBt5
YmQWI+WVyPMQac66M1LOiLqHha7rf9/4htomCuRHpAdQmcKd7dg64YHgIM18WMs5
98IIFZP5ZqfVicTsqulJO/gzoYBa8/u+Bz/IMxysUBi4j6BdQoc2GgyiWoPAIeFT
vtO8c3xwmqTnCIQxT/hmqrHEqtywy4lphNkR2VAnuaNUY2u9b+mdWxRbwXOg7bwq
CRsMJxqwxmRFLlBxEuhmPHHqV6+0Sy0kPv8FqXBSsqLjejlpM3TRZwx1p1j/CNJ1
AY5b96eRzesgZoqV2O12bcvaMFuQpb8pTXW0PjxWXYKLlTWBViRkqQgY/Dbje+az
fU/286HD0QkpXaAgH+Tks0EszXukf/xEj7ANI6RSe1lT5H/ijsY4cK25aBEwsez9
/58iE4RzfpThe/NNgxMCpsH2HsMLOKzKXFBbbyT9uZM3LsE651ZJN66TSmAj7wPR
5nw5RoLXMCe/4e4MwkLXzwgnRLKS/+vMWN4wfvElGY370iKS0oBtAXxQhoBsmteK
b1rEvSSmoXHc0XDuN1jp35g9GkaxbojuGNGANZYp897re9K4qarsRdMDR/SzcCT0
mhmmW+T/yy6kZxwCbRgMynq92xXkT8XMaWIA55llC9/iN2TMaHv1lNhxXBj6q5Zr
pFMktAppvm7XRwYGZQCn/9ww2tGh5yG6g6Bz0R2PnaosMR7xtZooyEMy3fX4VbHP
p4XT+d5uz3RZ4nev6bGxOu6QVynuC/enTRgx/rQ/teDHrdlJKOhCWzuXNYDz6lew
g4t1o+8eTaGuqhaY75IBjqcl+Myj9TrmlhiwEFkwUq0J7sEpggO6IWj+FylPEcAQ
Wfos5OwWQQcgR5OSOvurWTS7nJSjZd1ohZhlh62mEKGFy95q3+oRggbCx2NPgP8Q
A2FkzryJ0AR+IcGvkSBl5MffvSwOzBWtAmVA3zqEzPpAGRXuMNsQZutmFWVWhzuK
2+zx2jKMtOf1NIC4Ok/n+rB7Hgz/MivcvajK8RWT+ThsTzgCDjEcWXpO9dU6wqP7
CxgmoX47PBKO6aVyeHk5qi+iK6QIudIFaQrzm5CGcpU7CRFcTskGhMLXnQvQib0T
/gPFcFIkQzjeW0ToNipp9HRqOw8swxiexhSKF8QQME76BLHFJmqJiz3xlt38evqR
aOvNwDX7OLy52HtiLzX750lDKaeVxCLZmhegvo9KUZ2bAzTRjXlp5jMzUMUZQ+ae
C0v0NWLQxe9P+jjH+F1URg52CCtzHXlAQnOxHitzMlCruSr5OZrg5FcqDPWBEPEK
Xpi+WtIf3Kq7wFZCFukhIF8Fogx8fAfTDrloGxUzuMbfRjhb0AWXNVEQ6FPHagyL
o0YpwP70FhHEA8AaMj6P0zgcLdFAOTD7WBckZh3xljSJIP3NWaWlo7wrK1g8N7O8
v5ub7SHIaIoAO6NO9oGQvPggjYg/4DYer7CY/NEWm+1oc1WgSmTOEmzc+pcKC18e
jpzDNhxT8ah0mc/SgbS7dyJfK35WQvMszCYJ+4iSxtiMtf9F06Ugp1gej8i89tHK
RuWwxErxXJzjYD3nvKdpyZQv/6BVydbqq6s+jocBwoXV+Ju0IRQvea9crZDSZiWL
q6WJC/s8EAeCMbPzbZIrheISBDIn4M3gaT6I+VjT5pFLhpMFwkHr7M+eYbaJkVf3
IhJ0tGII1FHtdNTfFg+i9q632jOLbWfzCgpaL2+HeslRvQijRzTPw3698FNxDyp4
k0rUtOA0yC95aParL7XCKWH6xc7U/2Lzgd8zNLFVw23Y3fyB/NTR5GQSD5Kbrs3w
J8E4+vbd2b8MLL40lNM2isl9R1Z34Zz+TX5y8TYR1Dn5aNuZQsV4Bha7GAzYU6wM
qlxpjx8jryO5QaU7jEcg8KhXc7hvpTzUxe0o9ds69LohCcLCf3aaLa4bbd8sqynR
9qTh4USZhkWI9Q8b5Ap+COwPL031zrMjM+IFypzEbmwt209OrNlRqjMzf1m5OZvz
sf1o40v2P4qsAGQiEV7EJW+s9Pn/Omh+bQs2eUOWfvXn5wWiNlYTcC8luK+t+688
Zdid0eMhSGHJinsMNsP0Yxx8S3cC5aLiHy20JX0TcRgb+7tOT1YZkhno1Txn3VUE
MyiPRaZFoqVm5+k6FZuu66lUoRFhymCLb4U/DoP4ijB6HYYet51YWYI9PWj/PC0H
j+syhzXMLUEaD74Df2L433WX1RK3ga7UTVzKV1qTdmkDRkSS9yBiK/UcfbqnrCny
io7fKzfcjCUahmD1b8yB/hJ1gQSeIuFmg/7nKaY9dkTTJvhWgv4OJAifPfE3may4
9LXgtdSL+upZOz/QBIeaMglkKvPSbBdo3esuZRkMUq7W94GIJ2fWCW+Ysqbfl6LM
0HdKNDXhOM37lE5xOpxqxgrHt7c/ftnXz7o/01oQMUgF55M78CXjx61m5omg7eqS
nRDqtiU0tGws2SXxBN+kwVY4j/J+hEtS+CFeNc8aH+rG4hpptDvb5bbBbKvPbvWr
3UgjBMNIviqCJZImatBDIbwvNb6bMGCVUUnSIOF6dGAGxJnKhfTj4WI5q3JoGlrZ
yWgrECSZzt0StXTHxpTX9Rp/737miqrrB2SpG5GB/9P160nb9yBTr77yctCwsUl4
sfECvobU3F13BG3OfaqXcVICITb8etXBNz+0q22lLOKLvzRY3Xu/8su43uomlati
NTbrYuzYmGBEkT3rulhYJ4voJkqaTkDJ3WgYSwcxn0jJ4Ky5lmNFQhqzDunxbBwC
wkLvAw35+2d4V7GAIdmtzfETEgfR5BhaJuoL31ma2ZFRygPa6LZBx3gVAzvET/EI
8Zgs6HrjDFxcKjojyu5m7MKBqX/W/mhXD5jsYUOprilJqDZJG+We6YVersQj9F+c
DjT67hztktKfjo+KGz+kQOQCXjAfsIAflOLKGPtP91XDVLf00fvIxJHNh9LLEpIH
YK/JPtIwb1DHWp38MZI8oq4X3OO3KveMEbrrupfe3qbsEzF6jgpuMgi3DPnFEdYw
4PndHR5m74hEQUPQQJDH34+T6iUu+4wMNiyGQnaHSuzzeXuN1PXTJXXuUTHEztju
s6+syrxRY+M/Zo+uzhguF0+N1aG8+XCOcc8URZK+P4ELHVMZfuZ278wp+sLGuvev
SHu6WM6RcMSTnj/ldzAhmydy7N6UBzJ0OKbAFRYQhlxZMkizZbw4hJmD8usuAZoi
jULnsp4en1FAeXBatZF5qywY5BN6nCCGKyJd+Ob6OKdFPBkuXiothS6vrehkRO3s
8nnPmB1swBLIWGmazeYxjmjrSpwcMJs8ZUSWU0OYuE2hjx9tDoVCKKmEu65GN9ul
ero7CZfWaapbdO+zzLRsRxwySOsWkWkkgyuNaF78z6tpc8gwSXiUbUFKw3N2/pvR
QRPNqItmoO/DNVoV4QRNyjTZDNgOno6XoKemAgknZWXkD/0DGEYiAIrDA2u24f1z
f99S8AgnNXfypyjX2Q069avl4ELcQAVnvRgcTjcR+ClFfBKQaM0NFyLQNEMMGwCc
i4UVA5o1BPUIOWthB9VQuOJ1gPBH6SDsdYCvwJw5X0gV4mY+5bOvH1dpFCQ+ERI6
KPaadu7NBL22XAxCOiuh+smduhwQeZkVRrXPDfOBnHNUl9qBiUarHxtEWdy5FOJL
/m8n8tJ0u7GzYyus4hgeQVvdVArCzsILFgtbH0tfZwLqmAtnDxgYfqrTLMpAel6P
GLKZPU6egzIPZvtnTpddszIhNoYSIBCfXgJzzGz0rlvx7rvkjybwGyLMlgGl0k72
lGpWQCPPMDLhLX35/guEQlZSqb9c6N+NFn8Upa+R0dNjlaLAqJYfiQVOwrTZvHpR
o5ULX9te70FF/JoNMJhWF5g40VZ3hDgRwPJPdxxIC+PDPkuAmPUAUhX+YkZFW0Rr
NjvlNs5TgaJuKudDL/9mYF8HQunqBTT7lDxjRuewf+jXuO8mP/tBaQGNUPj4u+xa
ZcPpJRGVauS6xXFSFJ3VVe8SqJm8ntV5SwPHzRHoE74J5BIjCURUD65mWfR1TESL
7opSeBh8aRlGXuThaO8j6sSJNDSx+t0OCHmgF1evbYfUbHWLc/PAj3nAYfXg/ilP
y2eX9SS9hpBAuEgzyDIhxCwT75dr+ViUc72w9Rw09Skh0sXnc1m8+zt0sqwlUjPN
qKVWdF1myl9jTrYe9t/bVXtnoFSyLhUMXUU/z3ALoINStOUn5EsKW6iOAN9aYSfu
/Zva+SxY0j1KjBZ1LUgfPgjkwwbSxoxQTdMzLi0i/hK4Y21t9XzNxgNRzKjHFvHB
13fuwljgx4lihh9p/gC3MUcgUOKYsFgTuG2NM5q3RSbBOuPitZCcV5lAatoZo/0o
iznHPqYh7Ne47gIfxZfsi5LoGoNPAnklnAo8p2N10jv4iJH+8tACbuT9pVI3cuk6
VsCfBelc2o7iiaKdf3p27ANjbptaTMOfONg73hr6fHZ1EKAx3pA3jN6r898DaHEV
/OlnVjDxBTUrAFpW6MBiUjrGMSR6etCgW8HeFIPpfoxU3Kla+3MLROM2WL0LkpBg
L42J3YD7CscH3QYNyr1J3MMmksXohfblqsaEKbzBXCLvecONKhe+vS1EHUyIyKRr
6zbkQiRCuexV1n0NPRXo9xPAiD+iJHMfMawXEXPvDCnJZXdWnm/k36Aby3SJPKXC
LaZqsnpCX10Z/aPriVdpCSLCOiWNdyAt3xhrFKtZZ7Rjn0SNjrPPGC2djbQ9HP3g
x6QVn9F2Ivb3i4j2wGdJR5EuYgv3fiNY7STH8Xf1Ijxq72RiPoj29xCVheduiQQz
3i7Z3OFpZ+hGETTtrhyOBBsoo61DzE029UQ3mIUyM9OCp97KdpRQ3+HCUmO7Z8Ux
oFJU+rN7PZnFv5fyQ4cqeon3zuKLi9klOW+hKVzGdJICU4ecgjZgALRrqFrP6e2X
eGTChnS9THgpatevIbyICfHMmyGYkK27npsmWYBOC4QrewHD/ZONcLiKt7IfWbDB
JMsAx0hYpACJjcJ/1RjmdKPYmA3ODaOFcNCCtUcPq9nSmaTy6ctM3Z6LKHDxLtZQ
RLImW+XujUcTSu4AiK+Y4d8woa+Fu/5Up7IHPfaNBCxeJiFqi+g8hvq1QtC1gO+K
9zv7licEOpw8xv/9+pzCCeexGnhZs7bt1wJk+Nop+kBI4j7EmGlFiXvMfWTYQTYz
iQPy3AhhY8EI5DkCeK2Nhf7RcvdIfgAkghU2BW4kyC0duETBBI95bQff0RDRmtAZ
2FR2QohESUwfhUDoBcWHGVyGVha9zL4VaVpDnVMR7NDy9Vr5EEhIZJLqAuR5OpLx
6CiaD3YWk+BIUVjbD56MbWbHsW6vlDGpTT1UFThIIOGdbXcb8cZ9nIwvrpZnCes0
OvVV54RCrjWQId546Im1bLWihX0Fiyd0FtJKYR9y6QQIso8w6hqwp7qs3l0DTWAV
Q8VZ9UP+HKdxhltRcxRq2AQnrXuVEy2zyUpKt2MV/i2pj9KpD5XZuo6GPudZ9LO9
nCQskov2Swx5DVnhLpTagiF2R400ZT3stlm7kDPxKTKPjBFg5oJJpg/PvX7ZYZRK
1SrxBC/4UE3aaY/iy1YgE4INVDcLPz/q4k7bIRgbidY9ywgG6vI4CE7iz2b26V7A
jaHVLNJjZxf+mKZ2o8M0xDI0gtlq1xaBfHkp2qGkoXxhiPqGW12zaHb9PqriHJDS
gsYVYnEcoiH06VGGU8Dhivlqj5QkgnmoRuC7cgl9o5WZX1fwZ1UdcjYurmLepYJ9
2qqo3WwoZyRLxPftmJXAICM2R4dxeEOHrmc9S77lU0boYR5eYdJx2l/7xskW6Waq
Npu1kEIW2IfAvNdHO1TwcmLRo+HM8/Oip0WFGl6YvJIF5AWFPuGpHCJ13MU32Dd3
UNryYUD8OR4ZWmXv354Ldo9x18zwwiBIgE3n3UFxU9jN0efQRD1XvK0ueCPsy7zq
iIFq7/arPoEdi7WEw6CNr/oHHCANP/n6yLssfJ/8YV+PZKQLko+8Wxgh3+wIkgji
vNWeJlxxt1DEmw3qNvahbgZS+IhQmJec0O1Hj9d6UKJCilFZ9OFeJpRa77oJGbqI
5oGdTbtAv6HZHcJJoOxhMJORN+BnO5KkDfpIfwZgsNlLLt0kjM9GVz/alstWKA7J
CUpefaIDbtxIUlX+ZK7fnewRxeESr91E/rZ9fVGKtr0X1bKeoJk9h4jvsM4P0enb
KzZShxdzOmvMx2OTHwo66wJxUBRp2GWv9ROkGk1VS1GBED202c5S0reS1dg5quKX
hxC6o921PQsfosUT459uXR0xdjGoqHd0HCoEMNJPitvJY11mf1PdHIshsX8O4R6T
o0sGipU38+UKFs6KvzVARzho+U53mYLuq2bzhfFDxohc5Enh9aDCZvlkm/rG9epu
z9qQZzK5W+nvBisY3bKcUR4GTst2YyKT78O1NRM9BdEifs81X/zZRlmPNn1lbezo
KCTN3lmV9+emto+AZE3o3sFZT2WUWv159FWpyxNQC0d+wdXtmo6e5cEGrZuYCicu
y58R5hj1XuXdfrADoi9b40ejNAdhANL/xFOmvTof6bKwLqlznMZ1wpfQPjgHppg8
KVtM8giZT1AQdNoZb3SHdWnqF5EXlwwLNyR70jlA/936ZtUa6TWrUQQ5+whuzqu+
lmWbytdgR+WJtFlwMEb4NTpSJYuqUw2r0E95GtfBKeUnf0+uAmjILRwnsU9JQRJX
d2eKT8lU9B2Kop6YqepdlPBJjhOAm3wUYOln0g+4rmkh/OUMEDTB5iflwx/CkoAm
oAz1QsXTE4hJ2RHqdTXowt1+xX63xUnbP/gK+83M3DpBmtezxcuA7IjSlF2WJwCt
vH0w0tp2AEkLa7Ki8qnUn+jwhNUUUtE45bvY2HBMMqX25sgX34o3YvnbP+v/nyF4
6lmmIhRhJEAbDZejJFf3EpffxkFHePqPV6+J3mZ3WXQyteMqv2xT8zjKNQhv2plL
tYjVkwwLrog1ExGzy9w//e2IfjGgjuTtxgn456CJstEo8RbP1j6rXIfOcCg4C/WN
hLVtblp1+4Pvxc7ftaaCLPjXeiHf4WY2aDKqCTinWXF3zcv/fRP1G+5SWHS6Frxg
Eq/L5u3zUNATW7+GNqsQ0ec2zpkR4od3k8+iSC8N1xsiDB2KVO1u/pGi8IbzWuOD
XRdvPvxaqvJaJadXu6NtPFgsabEJVQbDUu3fvCWXR+L/pXuxw6jcyOPZ0HXnfANN
NY2g8yFtS3tyZk8wuFN9+NDL8ttvC/kSVmV6et0pFnZv+dvkPw8irSWxydYkhK2h
d4TkdiOWeVSRHQXt/8dBneWPRO2OJdJF4bxXZdKgOKsHbwDSUpLr7OD/lid8c765
lS84zIrwgWCpdqr0HDDQgRtnXfLxXyhSrf26jm1UMuZxI/YoXTPhUT6ap0Fkc+iu
ECSZkQQT777XBhAGV27Nnu06XiNJ/uRN2h5jUJuOgHwC3oNen9n8gNmbsoZPphiJ
RfG4eADs0v8/m9ZWgQZvxAuJsYR/+D9TYlygX5srvf6Y4Gep3zQg0jr+5Im4W6Mp
8PuUGolukTtdmotKGbB9sXHwsje6kOqRyc2bg+XgN6z34PNQBkeM0w36yQLaiKGe
TdvFBiFZiPYXV3mn0wlM+ZxOqKQgrLVXhwitIEI4T8b1z5dfOwXVS65FBQ/ASTnz
g/Vx2hKvqMODpHY7Q8aNRxa2emFqCuLKk13XHhGI4kXYIE4JYrbcM+wTS/8icElN
DvFAk2HO1i7MiSECI3ZAAWW7GbCUZF6LCfj6KzlIKjcfhTE8sFW811hg67VAL3OD
S8ml7/KrLFW9mFevRrPQuuz1wfPJiqQ4CkmYh2DQZgShEOyK4iDfk+MNqe160vNA
qa2aXtbywaHbQrHfFC3i7eACDNnBhImQo92Pqxg5OQvbwVXC//0N1D/GvQo0LOfW
+d5dMm1EleQvwkNY6f+zPE7rkhrHnZ8fB4OmrWXpiiD1/qvCQ0Oh23glcZrgGEdm
JTB54Ac3x/wKIWGHk75gMX0om7YMiEGJ/XIsmG/weM5H1yJooFVO3JXi2gR+4qAB
P3H76pNxEZRIwETNgjmO0IBj5VeqQy7tC5bBSKnTI+SoqfjZCcJxF0uHMLzUUhPa
vrg3h+rzKywde3x1PVYdj39fsSmXOJyQ34e3AY15RJStb4uzPaoYzGAU83Kv5qbu
48xpe1ngZxy3x2A9bMsFwytYMCISlLN0YdLAhHpI7d3cGLL7ut3vY83Fq54v94oP
iRahXyqZYVoc2znSAuumFGAp0lIvnlu2EadMaZaqlSyjxGfzjpnmfAIWsT02tgAd
354AwqbxJ0sDqZn5GRQlWQVO4RWLIAAdPKwdIO9E44JTka3bJovJVYbNt66BkLRs
P7A9PllUSOW2LYAvo70gX2YISjIdnB8X+MGjz4pO8EPIN+lu4j4XvSNAjCiuUNcy
3dDbajfMyzTA6pdkQebtdvt84H40K1edx3/hpDcwXH5fMwEFTIradxDmuSyQVR4F
EuKbhnVlg2e25ORRGTf3fuu+dAN/gMpFnQgY9xmAdNFJgqmewGJ7fvBUZANwqw4+
D8L2SPU+Iy6hmgo5DVIUIJUkh1iIQn4wcBKZhSeLaDIbg/R0jroUE+kthdIPd/PJ
5Bs2KwipYqaeq807JNEUtN9c2joAZb5ynR1qL8VrhkmRScUlngBZR54i0rdnF2HJ
CYk6EdRbs6qdAsq6719uRmmgvg1Rh5VqsjFZD6PN4BIoRF2B+D+23SN/oPXUkkxs
DP1tfptuIpGU8RSPlAG3sXSjEoSlqiAo/Op1oXThH66GT2WEHihk65dh5Qe4IMW8
WSS8B+8ReZLVifuL5pgHGMJnQdccARCbLBmwCtALPbNkoSpyUvDarJd7vM4MaPcZ
yL1gD1znF+nptb8RoitLcST39EycCZ8AjilTSUrWmR9OMoLX5NHa1Klw13OQuLbh
QYpTiqQLUt4+Z9726Owt7o2vx9RPpUVN7mA7RgBUnZ+iZ5Ixo5cp+yuJEpWpeZV3
vwgUpEqPQAa1jBLWlYWEDH6hv96Txxf+dAlY22DmIni5RMdNI1olEudcj2Wp00Tu
QHpdlMpZjCfNjsI3SVIyUNIXzIEhSs+n0CPyf7qQlisHUFiM8cYJn/71l1cDYBrb
tkOakClePOcK2CufvwKHR9HxNa+K9TxnOFpy74hTz/w6JTgpaTi2fwgWNWfeXaeo
M9cl2kTVWqu1VF5No3EO7ofrEVPforYWv1q9IVVdTQUXbZuUIhfiGTQor5s8QbzV
bzJKVQ8G0GS6AsGUClwg3daPiFrbka6KSFMIyQHvk+ztENXI3hvgX6/nfLoNcjRl
6/e4eW4i/pD8cVyukg6fJ9U50d2AZ0PdDHO9uTKbEkH9aAn4xe1XmAJUyXnQgpkN
lux5haesWtH/x3HI/GtOFfJH0eL8BGaR5TrV2rnIGaB2n0CW+2nYkwpEeJjf/+Zx
UnEd5+WExGEEzKeBnqm6hMp388wEgiLbxCKyXCMR3f39/QSX79782pcLXlbNVRLR
sKAdSuYq1Ntd6Ipa8Pkngsp3xe63qPvIMh4MxR+3dcaULOTpENFD0kAxXeAZr9o6
3NgZ69067MEG9IB3zTCsK8ZN0SOLvPwlEhRCVQdKLfE6fMd2nUH2v+j83jubjKTK
HnEbp/rYvntAZp6sVlg175djUItjM3bLFUU9NVyhPGVKNdM8o9WHPDTDE3bopmG1
mLwESNyVZmYNnVG0Lfl2ZsRL9hfxmfvFdJ76uM/F4l4aUwJyyu/bjlAi3fPc5pYL
49wPCpPXGw3pcocjT37KDoct/Lo1RuJ+8exd+NVTTeB6iGo3bH0zMJiNAfPz52TP
rjZlEgjaXYqSkle9LIqweES4G41BuAiDMfZoZRZnxG8QNt/7xq/HDQuvfzYBkbto
ugLlMRCO14sR8Tk2ePn8GUsl7NEI/gxrGq345+R+TeZ5wYy/KHorqtFdAo5aaaKM
YHC4hB7zowlNKRifobCfEnlTwl4Rxzc3F9Xx845YyJ3777HIv4Btdel/SLRZW5CY
WSkmy+R4fTbYccsTZHEGIgEC55QgxJx6TuXMxwn1az7eHs/dx7LS/UMzTLGL846n
LAq+E9nKiLff8f548V0X3QS6LL9s8AL+eT8HQx4IVx8Q9NIiTXI/Ie7MTkt9DDA4
UTczOf6LPJm2esAY9kc71Glj5bCU55QL8GfPDEK9iYQQRFQ24NPsYEGFdmACBmYz
uplLs02Zwr3nmaEL7jU/RcL43b6nHJduFBZ6lOyiQhIs6h5Sz3bg/IGkUmrzZIyQ
V7McAZq1hutbC3G1U5EfP/Y1c5ceC1UiX6WIZ7eJRwdmHFaSBV2eQdooZQ+ayGLD
pqGzU6DwNO4bg7UkC3zk+cl9Nfp9XQKA4GVC91mjab/IelkQ/BVrBy+ayZWkOjsU
CRvSDasN0ecgEKh+Hx9EBDWT+bX3CoRUNZ8mDMVuwhK6zTEH62/vuUoMVeH4rXaI
mMvS7cowGCubh3vAcJHn77VWKlxGbbJj8vICogf/QTK7TaVk9KBXLlWJlFDZVPoC
bwPojjhePpFJEFd4fiN+JIhkZvg0KisU99o4YJ43ZsFW84K5dF4srTTxqVmtD65Y
6wTGcaQBoh12pGVZWVyhFcYmSjvkgEX0TwdaeLJjfDNF3cH1yyNDvZkvmUTRKXEi
/IAHBuObtSDyoHg5iZ1isr7sUP6PjbBiCDzxGK8aUV2aU3eNLCG7o9qPxFdAHYbT
ZRfr7R4zEVdViDcA6XcACU6oTHErM4fcvfcv47NvAt7p1sT7ZQU6bTsvTRCKejb4
vewLjVPM+YWGClZjTPKHUGZ0ZpH0eK+5WjrXMc1aoc1UL89OqEP6YYgko9XAZLGi
OELYTTTagwdyCTglfjz8WbFiMnJz9CPJfgkbYfqaKHyd1pD5M0Na+Fq9mrPaW5W+
BhLx3PF05glwFP6yz3qwruavyXmLsekyf6CfrWj4bK5G95JUIX4JcPb7EQXS3C0d
w7rRlDj14XEwzLVxwJad03caHv+x6QJPTtc4m2gTe/anWDn6eQVPRsQmlLkVFT6B
jVMNdtYiXrapKDq7Hu9YwTR51mWwVbkLW162AA5y7KNzwshglWHYkavtti9+gBo3
qKuyx2aImbv/isyi+Ngv1oVvIUSl6Ntn9hUwnKFmgyot78zSXTUWWFtj6cwE/LhL
RhSb/CDmvZHqNFBvKEaP/lYFqbclZ0dAHn/spqSzRtDeGRXK/5wNI4OQQ73ygP8O
ymV7ZSKvBUPJ6e+LrT6wO3sZHngzLTzP9fj5CsBJhXm4NQIpTexog9ZL4T0CLUyX
QaRpnwpQhFXD5prQDGs2rxKc1iLK8Lb7Rhk9QrxLI9v8b+E74mSEcOMbuHhvu+ov
MrId34YJ5Dqtk9VKcGgepIlcB0oyv+cfr4+dEJr5ZhX+zY1m20ry8jAlz8gS1VxW
3dGJYhlBSso3gzETDqgPWlLJ62C1f2+6ziKTQ4dD0iLWcvr2wiu+tx+/htF8WJBU
KEqKFyu3OVE58hTctDHMFMUe0EyybDZIKXeYgQJxvx+b/EKHJY2CpFPl3N1ahedY
+z3wBgy1uDNp+tm/hPXf3hVARA8EAUX/m//d6KOyMUDxBK3vkEvq6ljKZ+JVjz+u
eLIEAHWC+x3U6P9JXVGMP6Hrimj46Pb/gVgB5mnMpQv0kp9KZPSXINmyeqm4JqH2
RgQcKI3gzuzy0SQ/s2ZWcRKdDsekyp1KZVy5c7Ez7Jymsj9kTXwfJUY8l8tdFoId
8bQ63+UeMz7HBtsWEuDSxQ1n7hBRnWEJbSOYMShjtboRXXoJHYWHfCydvTOk5KAW
oO6CJwrL8MYQR7tJKqY8fnmBYrxczY0TadjaXW4TaiYhmTTO81HQ4zzZfB4OdCLJ
93QKsf+Sq1A3E1Rg8RX7pujV5+Won7aW0qDM2XHQVnOhcZcp+YqKyMGWGTAh6rnC
U5lqU060Zox2Y11wPOHKLae0fhZ2v8zTs0PH9XYQ7FpZd0z58nBrc0rYtpwjnA+4
MPq0EYL/0r8J/VXIyVAuXFExMsik1gTEKtuNJc2IgJDZzxzckMuA2qaIXyDLmzBM
vEgFstuKFy0hKrtiLuEa8j1iy3xs7qg/BqeOALnsDalR9PZeNRSAhcbqImHF7rxV
IQ3Wf1G3YVDw5R2oN3jcoiDehiTpsjaBw5RHgai7D5JZTuNWgd5Z83wD34RPlBuT
8SEs/sxDAHPOdFzmuZwi3/ECZL/+j+9FPGduYxdPvu9Vvp+TmI0Kug12iv+OxlaE
qZbuQ/drxSDwUC5PJNSlMqsdSrvNnAUrApO4QO3HIT6KRMVR/ZQohjzOTEzELFEr
LPMnmzczYiIoCbOoxNZjSBtfCbQOKMfZhC65MgdoLyakpgM1aHr9uq052O/Ypkbj
7xmrKl/8Gu98elcXtAWm1fnwlRtAhzYTRb8khkWzImk0bwAN45MmQLSYMVeWjiHg
mnDHOk6glB5BUS/+vhi52XDzN//PIoWslRNvQXcMyQWYcFfe95MO+NuNpDSfp9Ae
wg3/bazy5y0yaes37eh9c5hOngN/cUh8y6yjzhBHMCcKaZ4FsJGYVRFMjX3vj2a5
5cpPzNXGTlBscjhc4hRk3AmzuadhcEbTHg6vP4Ktib9jRy1eZiYpm5fPEnNOFzSh
quYrmFA9GyEra7UcAdaCHrkPbTts0bH1YZSLo66dmvM+lD1cWdEOtJCKrLXAhMnL
IXexCOiZ+DvczosyVPBm8Vofwpz7+ZfxG1i5311DW3wfPQ+r+xZNKj7OxJ/OYP+/
q+RrhR3pLk7H3f3JYuVhtv/fcOnjT4+Tmnlxy+aKz+TKGmXojqggIZ+qnVkgJXnQ
kQdg940Br5ooka59h82DrQKfuzDWgjqkjBBvj9M92xId4Zvf1fhpG8OU66gh0CYf
dOCDmcMRxcJkXXDnLuefikK49x0SS3tp7KNB3dcFbt4Kd9Qu4jVY6RO/je1cKATJ
nafkoOpruTAtzx8eRezdtn9Tv0bAUF9aSIoymsOfKm9AZ1PJCEBhDIWoB65qVUqk
Nb8yt0ieUe3isQdVqnjP7JKlSdZO7DBfi3UD9PlB3NRF9lafX6Dbyw2Zl/iuwdp9
3rcOaFYfnrjLFu/xW7W9ct9wFx4AWQTkTpNBGF7T70KvW3BPtO+s6Nl1/6fSbCYo
RRBRczK1laJ9/ZuYhm4/RjYFVSkQCzNNr/+7FaQvtxv7O0TVnsz34/dAW8iDtPBv
gQz42PCfDvRLiPgDP93DrRZuw6EoHl0n2YdkMM1tbnTZhOQK0ovfmLt2XRjUq9Au
lviNSvB5G4vIMxP6lm71H80HVDuJSYtKJWPGnWpGqHKFJO9Q6ySGh78EPqas/Zlo
GFw0ZEvyMwaGHFMKgarAES0Bxr53hdpB5T3jIubQNH4TPBOXnLvvBJ0VGhNoj928
4wrKiZwXb+LW/B9HZkgdyIRVhxyvBFh8sjQsPKCL20TugeN8CXj8XaHAbhwEVCA9
T7jEChWhnxLSsdcdmV29MIffNWov/6W/NToMfHaa8pEp/nu40rzUfzoTJUv/xf5P
SvnQMiNNHIW9IISuPxyhE89slICIifp5HgiFnehhZ1jGAyR83DWud9ugWASxVVWw
VQBQDddgkn03t8Af1Vjpt18tIzqULT3P5Tst6IBoZDnx7HK6UMYeaUf3yurBRza8
tncZqKlh65+hOH7IB5raQuZomO3sg/WpI6X1DjhXy6oMItpIdwCiyr0CX9DV5BUW
U2RhfIVoqB0dMrsAmkkTYuqbqQxA+N7oJ2RInK4OMW+a3cwvorDUz3FUt+FBlti2
jCsHi/XW971i0UW3rDBDvCzgoGI2iEZUNp0TfgEn1NZ8M0osTICmRJcGm0ZrUHgT
67yHPwn2R1jsokVwcF9wChG/T58KPHwSnuNexFvbL74LcochJPE3SHK7NH9P4vTC
N4Fod9XpaykGYOzmdn8OkUrk6HT2IX5EhJWPxKTVw6Phbl05O3ADnA5Wk8m842/6
fShLxKV+3DnsDYh/CUy9Gbux/bOvoq/zc0MXBEFjF5qBG2E8wmRODddsMThsaVLv
wWBNZXIBMbCI760TbeatwaWsuiEF54TdQKaPSxMr4ap8ACmjbC+WoZYhx5DksRFF
APJr3RPbh+Jpsrx70BE8V8kUf+ZuCctW+Vn23hE0eMT8FMQ/pcse94SX5xkBjWM3
sI6ae7+DgiAksQ18k3O+jkYqkzMtIqUfeaWF3kkNzdLGOPUeHSHa4dTbSpcblRak
jkREYwhu7n/7xOFzKt0IFlKKr8fyUefiJ2dk/rQMc442HJz6UJTGdEZ5dJrq+Byd
CKP1KYHyULzYmXzPqsD0cPv9PC5NW+oFNUDKTOn1+m5Lmryg1DFkvBzM8Vqb1riw
wba5llmbHhSi8SJYPIyvEFkMHlNO7glWVNS5NJJxj9Sy6XG7gSRRZ+LAZP4iK00c
XSoVTqKZYf2ORNa2CIJ39knlAIeokYc4FN1Njl+2bO7lTTSzia6KqfbpDbwSG2i0
o3CGUc/AEygV5gp+nfL7tLW+sqkUOHQfivo1pU1P1Fde1jXjBnEDTmg+5ktmCZFa
rvB6agDqhkRA5gcQh4RhCIcJve9kyeduDt43HROzAvMVymTIfleCBXEYSVINmToZ
tA1ooa9mksw2B8yFrVVWiFouuagycu301GzjWkZ7WxO5amGYdtwqHDlEL/Jtw9Sh
Vyz/ZW2BuzF1VBGJUDeJhKeB0InyvXLdchX+OIrAah+ZoKU70aADw8Wy8BqaqUll
Rpj5/iRi7asZI7PNEOXrYDGndyDN4Qfwww4Pprxjw6zcmJensKyWn9oldjDXwArH
LdjpHs5xDtgV6BXNBhclmYOugLqS2XQXR1FpF4cXRq1u6JWz5t68m5var+MSiu37
2X20RbdvnxpTx4YY4aUcqTgPOTiaULDuSw/71FyLpxCgvnrCxGpwb0bBmG4RlDKQ
8P8AvdewHmydkXVeh8y9OI3i70kbU3KC10VGLy/3T5K/1ZRYegj6e9U6AlxEphXN
TbAxF+RKeI/MNHO46xfz9FMeLCL0YJPgco2P9M3VEsHYFAqNjy0YCGRY63BbAQ3X
0I/wvACy+0nSJs2SLIjCsmA3faxnTu0Qgsd4C1p/S1CIio+v4gGX7HVXZCE2oBFP
C1mID7R3IR4tEx0lS3rJR5pFPNVUAaZYBxyBAEc1qDenJgPTGigeLLblNQi7UG2R
+H7GnZLLUwkDH6gq70iMRgHGrx42MtKrtJ5BHYGa3dNpsSrJ/pWtZsvXRdlKwEn1
UjS4Veydx8vh1PcNMMB7xFNRgDbNDUFePdc3iob2eKfkwzVTwoIk9ZZmXefmNVZC
DJMjS/qnt63KchBe6TQOljledxsaRurI60B4AaVABf4pBwPaNz+bwruqMKzkSnMg
GRDzS19bd4uojlE/cJ4yndgNLw+z/HjoAvxpfIUM1eTMkZjTrhT0+jqkbkPyPy3C
nSHcH0eYJdRZqJOpP7FGgHkQYN6UPHG21P0WP1V+qCnGmUqkaTte6YIEG/2Dxm7l
rVAgvbYdYkek690GxTpeEcNCHWgfhaO38zZSkuL8SXX59Q21VPpaEPRlZrVvG8Jh
GbpPLNb8WQxLs6IZAhY1jQAHTiwR7R8ZfoE/PrLgKcHpeMErS7h88//SqfV/QQCP
b8GWEl9wBbDU7NHX+pOEw1/xxtu2skqmdYlNipVyxFI0H6NpXdZZofnKB0g+djYr
fH0jZCTkhOE3WcTYlPU9FBosT2RkJBUnjg5vzs0mXCKA7jfqAmlHMzs3YVaxQwv9
jqCPfo2RP2quRpHQJipJq3xZAD5OUu0PeyZqCkK0dLS1CkpkstZ7GDMu9AYCZig+
fkbMPKRf5O55vceYghq51X9rP2y03fnHw2yh98UtqgsCupyz1ne/xD8Zzi84xreE
a37ExW37LiDvU8RCTg6FVwPCUdWIzou0NJs8AY0ZjtRYNp32dfVPKaMMwBH0ZgI+
thKaaIed215FjdFeopJj3cu3QTrsC0H71h5auD1gwVhYV0z0ykMXCebR+MKRoBu2
eS6jDsm+EN/yLd3JfprRf/ctNfNsV00EeGjDo09M2HTEHQix0nqQ6yTLW9fAq9cO
N2bIwFEigsVGatHxGu8By9O8lmo6VRN6t8ovp3KswmZY+yAnlWtiWOyXmizugZ9d
PxrH1BslfWYvrLzdgEkX6nwlQ3EJ/i7qRnOwgEuuh7FBI7sz2EZso6dGH2TqBwJG
nqrXdA4vkHt5fu0CrNG2d4pbdCQJ1MHf4UuJSEkT/FWOfy5Q8JYlK5+uzaVOIqtK
LMxzpoNz/3kfilC8KgmyPQdCjp9MTqbm0774zYdQaRtFw3Lr0Ts70zP5zZFQuzgY
Gtj/qbTQwwvHKXfSrK3kEeesC+dg397AcMjLSle27MNXpZ/F9vPXXQEHjgEd3Xqp
nqwvAfaxV1hDceF/HjtnIdulw767yMJctm89QGUOes51FAs/IogoKQSBJTRen0sx
6yam6KYtnd+xa74o2oTkEiAzAjMfGnrJ6ackZVSRPIHYIuOxa4lHQROruNp8p0MA
lhrYZ8ELRlurcfwtouQAmCRw2gUwEX6B3lbNQjbVgYsgbfFcfRecshztMbF2l4EL
nZRnV9AtYtW60KvAUM297MARmFHmzz71c/FlPdfq6HBuvrzj6528y5DvlXIkYMaq
UyUxR/cE1Jlb/3cKS4mvsxepy3tDb+xgjYYx8L/KUKculEz5GsCMuM37Nqtv3zT/
gZYbv/bY3hfSLih60ZfW3qLoWjhfTenwR5hiL5+eU/MPq+SofNu8UGHQoRjdEOnh
MXvMMm/iKzn3JVtUDqerlTmb2ARj9TX4CQR/jwMEsZWfth7cUEGl00DB8ujwqHCm
fq9klmrBmHHVcpNXXEK0D46smOjPAq7a6gKNzXo+Ra2xQCYNqCdMFGpQnAXHBNLe
9RKVV52mkA55R/3BW3ya0l3KWxLmoW/y0cmddC/6ZYRMKQUKIalvc4Xee8yRZyJn
p89ovdgkGMGcyHT58Uq5ztQ6g4PkWCbyf8JPGR22hSBytSwaC004upgre9RGx3xI
k0+N8opZWJCgRp81TuKuRBUxsGbhJmyjGUIh7GpaHV2nyalAretfRTStm73xyLZl
AsFjMv6SZ5y6Rulb/rnNziVX4fsVgGXm576i2jLwVeFt5qNAb3cVF46ngo+5X2kE
GHLuFwsuGtZ30RGZzEcJq+P6MmMBslJ1QvIS74vFGXSBclbuNggiIz4GN+DKEd7R
XUjvl89ptggghuuMZ7qcxaF6f9Mx25rOpBdTbF/d6e1DEfBUYbyNpNUR1yAo373O
6ecZKaW4YtpgMpRy5nr1YdGjLzueyOFzE1k6ydDXi63YSd3bn5WcAVreJZkQlAGt
asvezobo250cZ5lWA7OgOiEfCHxNeykrqGgLnMwfov5zIMqQJBMUdyyjcjF0q9Cg
C2apXBHrf5OAlHlGrcbiwP5SxKJDAyq8uZCWoISNOK12FkzzXxcQinNh17x12iws
ARoc9hKb863iktWHOTUTKX/3B+odp/8pB//WAt0xtuRnfvS7og0zmeBag15Z3fsl
7w4acXi4+Fijq79yhaPlazJuWF9/c7rjMTScgn09vSmDQTCNw15+J1QYa3YsoyPr
15/GITCKxnP6R+KUw5eQV6M2kSWzx9fivmqQ7czAWMTwnHVIhLzaoNLhDwpS4M6i
XvVkam3EG8GaWaS/y9ciN2YRM+rO1L9Sbz40Osl6XRN6NHYOwMjDAIAddFK5KOdX
wUneUJv+6huRottwhyUZ6gN1vUAXypdtDs+Db9svhkBemxzXmOxS6VRtcOwlRwpS
WkbDiNWlT9E2LOZnhzt2Xd5Ulvjy1ofnmE5+VMI2+kvvSVVTJR2PAi9o+2Abth9o
WNTGgbina3tJUjvQBpkfHW6KocKdbibLngPbx8G5G5rXvbgxPNKC9B5CeSZp9jxq
YyxRsu9GzxQz4rM+/agUJAhvuG7hJc2KRuaiX0eNoP0cMtTz4GR9UHcPJkkdIg96
Okni5wLTV10g/QvMnCQe48tjQlMOtuhIToibxJ1QfTuuvfEC57vWFH9zUiTy4IBP
wsn05ESWnp361UaoEoBEbuECrzVLLz1E7aJt8jXE6SGkfOX8gjM0hyB2vYHcnp5x
lQJC8j0wQpvL9w8wDiwUiL+R/YVXmRsCjul4+/petBBBlD8yJE2dM1mYSAh6NyT5
QeYCoE17/xb3pCroT9WY7yW+x4wXzFPxLiOJA7vRrXlFz9Ogac3CS2O9/kV+ON1N
4jm7sgIFl5Np0cTw1A9/LvJLVpf/BhHnKwR8k5mrpQIZrH53mRy6liODnfMZltUh
rn5jmQKskVMLmlnMNmylYGNnSHUe9y02TdqWvbdUg5/UbiUnTNbesBxn/Bx4hkqh
edQpe3O3iBeU1pKUuEW9FCmWRqq/LknHek8F6yrfHeeETLsceP/C8Iz1wap3rmUQ
xnNRTGhZRlweKYmVZIeHECp4RNdr5Rtm3vPeVC7BkmdOCl6fYQer4PGjUJYxOhvJ
/4ltkzHcGBnq8bfu7Q1dKdCVusBiNBg7jV9cmrfTImzg3OOlieqVMGza5M0Rk4zC
WjD04Ws9yFrHY9LuYbLwnMwIB1hSr6SY1M5u2sC+q2Jd8gr0eS8uUZ/auPSubFos
8giI/p8cmkVQBgwhVQP8/RZzoiFtp9xVUdzx1WOkHNI/qfAYcQgHiTrTAJ++a5j2
uhmZ1vV9LlXKzcahCftCpl2Xca0agdHol6BHOe43C9JX06lc6qMrHpFTkqdrGNUV
Wz4FwBAJjd5z5AFmoMaAxsiVt5IpbrkwisyDmgknpSYcdobTaw5ncPEFMcMH6wGr
vK4hKykY6IFe2eqFqlebJXPFXruTs13k0+H/uhUGJoHGeL5l/bGTSptVKB4tcVq2
3B3L73KVx2EHPJjLWboFRhndRwTU6Y/dmqZ708rE00MNp2LrJtsVMFYR0O9BzeJb
FXPh1rzQqMkXyCgl6aZfdnNnrY8wcPChJU2px3Lj0itumE5UqKqR7Rt7xUCTsMnt
EOSapNJ03TAgLg+pTtGnM0h80qtvndddJHHH+uj2obsvm7vRqvGsrd2snuFyuI4k
Yk29ljBfrMxgPewjk+EMixdBu8HV9vQzotjKp3b6DR92k67Lz3dJlZc7qrTvGwD3
qEc/kkRfgi3EhS5ICGqjQ/G+NNZKVbPJBzeXPju10e8QP3ACr51gSqi0xG/9b/fG
sVI/7rljd/7SFE+eDh0h/4Tq4HiYDX7bdZfwBJ9HrFv/J9+MbO6jeCQ3IcYNfPyU
VSzWdH/K65GspfABbBq2bLz8fSWFAyTL0msIT6bZu+egjjpKI64KktGjx6J/5riB
Qq0RxB+V4uZpcbj80L4iVtnLgO272hUet/tdGmRaqqjMuHhwF0qXz1ixDgw1kOvH
zppHw11Z4GRzGX4dyv/KpMKT7IzY2nBWcmzUY3ZIHXjEc90hU058abSDKVcyY1HG
mzVNI8sgOjdtiPxI/0RBoPzdDvh746cE7ZTdMQIk15B/DAPOrjMOqdH3aU6zEHzT
q9kE7X82EzUDYdS54U9jXB/eOv5vXQIjWxYH/G+M+uDPH1PoQKThG5Q69dF0PF3F
WfsRqdNPZlhesjEWUXrtRCBqlDvodYRHPfjLf0KEs65o/Xk58FRC5MF/BbKxYEbR
LgUnYApLgfrWxvEtXE1HcYdAgowUQHeIYko96n2jwyTT+KjU/auAsniG0AXNR1hl
aaV9kIDdf4thzmlx/i3rNyJDpjuLX/42RBQSU/6WJj+rn9E5n2deLF9kVTm+uGFZ
EHU2QH/ySadNxAQD8OKsylLliwAHxzFwrh/FUmmnYHuaW74ZK5LVcDTQDRHK4pIV
7U9hjAbHgnZ6jNHU6B4fymgZwXxI0zUz8CB/sxBIunrLVDUlSwZ6eLc8Z+ED4eRl
n+xMsAIpAJbZqdsIRyBeX2xLCyDOMniR10+uH253coaJWGZXjTj3BRbDO4+0k03h
mXtzJTj1pI4lJzj00AGk1NP3gmD+WbjoCCii/N1rbo3lWIvvbHpM0NGXZoDHP4kf
C52tMcFDrj/5+Y8YB51MrMdRa2FsnWKsZ2VyBndrKfbgqBspojxDIpp0ZrO3YLQw
4RcCGA2pHRKzb/mWfLPWU3WzDKYBVTG5scAgNPoMA2Rul5QZU9oRecYPji+PiDO1
5uAVBMksSFrw5W188BQxyjPpZ+i6+Lt/Uc2LLZsGsJWfgAgI4dzrJRJ33jYiwEQS
tkDMAq4TzZxzy7/kzu4o1Pl151tXyYXzUUi5kfy1Thlwt9HTVrRq6CFUE1qVqZ3t
+ypVUoF5GshEOmRdnZXtnbP2TxXmv/c+UXqG19ScuxxHfZcTUOZqoPMhHQkG+SUz
+veGMGbnkB8yq7YAIwqFRQYEnt3p4BLkbg7lCQJFsoo6rRa0jsn63MHucYphm13N
c91aF/qhuynYeV5t/KcG9srs1IOrYe1Nz8GwbcCX2dQJ0E+8XKLQER1Zjj+cMXgr
/VLI1t7FerCuHbToNAZ7kJqn3fJ+vFwrIloWbBBRybETjd4XJMpO0YmhkQ/m94No
CVOOF5UaLviHWnYQsLvCpNNYGLHwNVAzeZbqtWzf5/8fTii+Cdp+cD+5RuNgFokE
G5/mdqZ5rbiVkygDwcvita9gpTN9LnzKUIhYS5AhoQLUsHOHp9feJFgwGoacRFBx
b0tvOqlu0HHM91I+aKNBkHspFvIL7RF/tENSbrY9THdnt7SKvEq3Z+3NbWxgBe/8
6fr39t4+Zv05Mkl0jjYIH/WwjQydo6SvR1jhRrChYF9vTfgHwMGhTzJfPnzcJ1ug
xY5RBJOfB7EhijZ7OhwCxW2ubouWDHOd86rFogYiTawhyFZS1VbpKg4m7YlHA+LR
zYn9Q2uG/DbhE3ssXO+zULYc5RZuDT2LO7QCUxhb+a/voU3t0RM34x2ofgd90c69
pxQq+LqIGOD3jZROZyfXYYqC3BwIMXZLF/6N3Tk5ivjbd+cwe8kuvkEcQL4AujXq
YFzzInnPDP0+hwHBVjkBuvos53uNgsL4Bl+Kp2pPgOtmCobpKmY3SOmgsCxLUDGX
zp1eIk1ztOLvA5Mh8XUdTI9hWiSocAn5XKr605vK3ahQO+Lm5DUDOxFq9bX4YCZF
o/kWAPv+u2pgJ8GeYAWLL/r7wJb235vrem60W14AvIZUbdsLqQ33Vtr5FTAMDN8h
0gkX9cw8+40RQTunklSJxQH+VxtSWIQNC7lPZ/6owu4wD67I6wk9sfpKNetiEXHw
eFh6qZx/6ogRxtKne9U1jvpbyaT2nAD9HQ7f3/yroVpjXrbSseuOI0oCUsI/ODEz
Pi5Q1IH0wNAHV7drb2CRlygoJSvakV39w6FMmUkvdsIHM2sq2p3FgZAhBeBV/e9a
sEK3nNxU5sbkyuULAH/DpxIYo5zLl7XZT20qUA+2wSogxCzPt8GQXLHy+2IaAOZe
YV2rVTKYdJVpmKWTq7Y9EVmRjqUIQMaxywVRby+EO8mL32O2mP1webf9G4lLbm4Q
diw4WGAtaOCmRk8ZQXtpcj5q4V3cRgKfp6yo1Le8/n9CWLRSjo6TFaXDamh8L1Mg
KCslZHjcgdRCo2WLaBIFFvax4LP+3fj9m9i1TGwyeVzcsAZLb1UpzHKXKVYsGWLr
dXdi6XT5VH5BnIj1ugci8kfMYeK7JcWuyQYPIN8oxDKO8XEdyHYrp5FDQKDrHWtR
npcw2hqsRvaKR2ugUm/fSkkjEfhuB+EL1+QVb33ZLZP7EIao8jRg9vcBIJKcRKnV
agPtu1YYJOIfFp/ag87vOSDQGQ5ApX4K/CZx+ANhSUYgGjPCpB0CLkJr5KP8+PQq
uOcRooOpGIpAarToLLj2R3xhYInBo7Vwl04EcaEgGx1LsNwvVWd6mb9ySaIm7/ur
xrt+AGtma4xlPpwkFKpZv2YEz1lh3+7BPDjHyuWEN4WYQ9w/+Q5LxIWdQZwCwRRl
P+YLZclV2yiPl/f8TbyQ2rsnNsC1GdwFqXalDn9Vld6t7gKif2osU+M0Q3a5lRZE
VPtCvh1d1J9AqRqD28WvpLwOc56wCACZ5XiGqi9k+CuUSc3g5cHWwrjzZZFPG7oj
ab1h5usv5OzJdDEdILm1we+OmSpjEsSKLLVFdY/aSnTW8TjA3Hol208pGFzbxVKR
`pragma protect end_protected
