// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
mdggavBAwTuv05Z/c7C4QWMKCrnvgV4Ft3ILyy60r5FqgIokLpZgYxy/RG0u/a1wrZaMKmok1Hq2
SoCh/G5H/9wwFqNDo9UjkveEiNrAWj3KBSdqCwiWZ3zf8N4iExY0HRQvREn41YS8rVJMrcm4YEoA
mG68PYJWikrhaIvRT2J8wQ2A3Zwo6EB/BCUICA4F890aiz/ijxGJGsT6H8Vom/NqWv84YDV3TmZ1
8oBfv4uxiOtOMGktn2sFqW+pTQsVgCSRwOR3dpgnospb5ObUirdSYN1WdZ0Pko6x/+KVEuQCKep0
wzr+uFVDpHUms2kPtjjiPq5eFtNS+fIdLQjABw==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
6ERpcQJzuP4+ptbyJRhEwRm4tzeoyT4tZ2Nvoy4qVlk8b97b3uWqXzLz6fSR8o8cAhmb/qiU7aw4
+4KBtiOg4q928KN9+6Nyq2HByoIrM3rCJL8apwtS/CddNdwGmO7FnTBYXu5srhfd+cqgm2ezawPP
wWyVwKSw6PB+iRsrMbCh3svHAVOPJbgsHVdIt/opFlU54jkYk2cgy0YzYeFyfV+xwEN0YDr5jJ+8
jyVSEULjCJwP7QD+GhfoCypYDe1YQUaybQ42GTAzLDkvNUofUg/MTQFc7Gl+mgFQKCLhJHNkbPk5
nJCI33SnKugDzcQpR8Iwz62v221Nv2hWzfat3wiMGU+GhkV3iYA9t3EqKEakDU7to0kihHVuRgZr
r7Tw2nwoQ9XuU1NfBzrvSo/AJ7R8IhHXgdITFpn3bnft6Wr6eubhnd8aDIzvBIhLbuQIWOWCBuFN
s4liBOqqD0PRWKA3yMFE1m051xNzPx1xTuM1gKUoTjop476b6UEMtRUIwe8Rp7hL9JQwYnHYmN68
mEq3cb4b09MQk+zisVE/No0tSakGXCgJdWjH5TzzZR3MsBziM2UzXHGwea/H5RgZ5ftROAECao9V
sIUgg9u4UKU4MzlH3A5t3H5QaoO2EbPxZ6KiNfEuUJprWRPMjiIyCPCOclNiEAj+W5rtiLHl0sxM
3tXf6RyxXnrJ/dF9jCgcguhbl3NGnF0jkMMQ1B+cPTd3m2EaiadGX9g/3vxC6IF0HNphcveCOWJ6
n4HZOawqsI0nwpvP00S4GSKKrjQJH2HcGzgt4bcQizSoZdeeIv92xgikQPXU7QZrazN/q7edQd9y
zwcrvOwUIzexeLXyCzcunjbPs7QBEd1mNQRr+hWbLek2A+sVkOtyAf8uw9GoIHaZWRqlSQ1mnuJu
v/sCQ5b2mQ5DbYgxZ1Eqw9ij0MHD8dPfboqQ2kQ2TMzFaM3ZNqh/+42pwbPfVY85Jk4TVY0EUSiH
aMwvlLpqPwPckZWoJ7NfCfKd2r3Vb3+dd/pfWNep+v32Gg1my3O1SGB1MdfWoN57/cIzmFl4S9O2
GuCFuiiWGuD2QX5Z0ZFgQFzHRMNEj2OZw5k2Iph4xjk/p/HjBpdS/iFgarxor/pG+PoozikPqdve
9IvW7jY5iK22p6P8hTUPCqfvoFzGxhp2rH+Ux3LMkdF31JdIU2uNHwp5q6fi7Eihw3qifbthseET
IFKS/Bg/Fl2Xe6tIQy945PiKE9Wpr0iTySYeiz3OW5iLYGXBeQh2ZJG90OuOU4s8jOmQYNHJmafX
U9I7P7QvTiCy5R3yv2O3nnAZhPZZ3c83F9JixRFe+HRly6NxIU82nqQ1jLuebr+rMoe/7B76+4Aw
bmWSQxZKFkSkGrSRNwJnqa/QAs1DQLmu/3OCAH+wqDX9p+EL2QD7nZ/+JqdoXSjUOGyOVklTv40U
zBhG288o1PLKGvcHfoCOuw/HZMP3hTXepzNXyVIXuHohAxXs3kyrw08ZhPVbxiZiKqcOMWU6nBTV
96Ft38FNc8Wp7rG3gJZD9ucbQflgwUEmRs3qEc8BIGZVJWwzG5KJSorbHuHIiFaTBzP8s0S2Rykg
AugYaU4BArJ6aJRqmMU1yJRWjBFuY7RMV2++Y5NNvb1/TCtORqkDO8JRCSY4BdcqPFx9e7nPw3I0
rEqu1l9vfH0ftVdsvU4PF5zbnMlNfJNlVmcbCy5iaGBUBnPep0he1D6ZXxZ0IMpdMBpBMW5HraA3
xh8+uDrzxOk62wQp/T7tKy3RIhfsQK5EY1rbQTiT8Qk9T38+Ssg8M6Z/+Kb0l9dOu8CJwUENBwfo
alAPqfV3caq+DVl6o6j6i0C7ijHttBvuFEdHzl8IUL7Fd59pd6F0jN8ZrizY3vWFRHRRKXY9EZqr
v1cXFVnNNJ2XauuMO90RCo+2tac9gs4OK8UmlgYGJDrTFZ9j5smcmkI1qPnEQtNS8a4IZ68Ee8B+
09dPEuvYvE53SK6kuGilt5951XL7XgqcAe8ZXIqEZspnl9H+ommOPIBTJV3Nk4E36Nvko5eG3M1g
jUO//8ONwC0lcOwPJBQuakQRwccM40YWnamvkMyXr3hvHYqH9unjutn0awZku6cqLH7U6CD5thdp
vWge7I2d0rRUmIpFchr7d14wmI8rdzyvl1xm6Z+Ft3gs+F2s9/RmUYvrQQ8N5ueWW+ygMOvtlfpF
1zNd+q8++RtElxM42DjJzi+7FRV847FXU5O9B54Sd/HyWbacnE+cBtU67fPiXYeWcP0qGdMaVpkH
/66u+sL/OfR9eM1HiNMNK9s9NVQxQ3Jdvk3a6nH2wqfSpkQ+yX/SycvXvMtKxqh3uM+PZnD5GrY9
8BeiXIVjpcRhfOsdpXEXviQ/xNGSAgTBxj73Yg4ZrYWO8UUqw2jiiQ2czQ3HEub1ZCyECWzRQNmz
0/+9FWJpbc35Rb/Ab6xi6pdBabN3VGEn4iXtvVfvhTdGCwGbyWR5VjNH+EqXIsPIh3VmKLHWYnJZ
mdP9fdldQ8eRej9zu3QsEEtwasT060ImVXLqe4A8OsZ0g0B1wy5qFJNFwuV6Musioi9/+Cg3pEsP
VF+GWzhW2FnpCZRJiH0EY1BUAiaPsVDUWRlp9UUBKXOcrFj8vd36az4jmI/TTGa5ce9PYYyCFxfo
kxdRyWHmz6GF3QdUF7RwWQ+8CDZlANG8YGu2+iLVxaCODOYXkDrzk2LZGWki81nIuUXr2GBumG7u
2bHfVRtv+SZHmdivhDE7HEjEUy2XYucjjxU8Vj89pMP50111QyM90SXtIDz2e9i2QNQIAS0ZcM1d
bel2qCJUym3ZA5yGNwyvyMy6Z93Z0kMeln5biPiC6x3WnUjQH4yxR/B+l1FEFl4NKF4SAfYzR8HY
OWVME3dCF8tcZgeR28l/mn7KJadIDSHj8pNZMqputIKym0cNYvJBQfNyJImg+VoXfFfUsJ0pOVx2
rLy21VWs7Zm2yHjV4cM19ZY2OX52RueDBRf1GHwghLpxkzsj6yQyan2cnt97dgcqsQc9lmCGdtfr
10pcp6OlxHmwCnb4S6jHer8Qk0VGWWV2Tq+1ENG4vhharDBRw26yKgyqhx7Nco+JN5nPpaHiSr/i
t57k64B/D1C4EWNHE8qVKjyUklYd1H+BRE24nG6yKoIOhVFa3tL6lQdI4QntCmp235Fzs8MfsYkJ
/K2x748koODrh0t3JWaIlmsyGRodKwmt1IwLZQOCjBLc748MuFWJSMcL5tWJwCispnIEkZhpbS7f
Pa+UIIvEnzFYK2JGa6r4uM2z/j8txizcGxp/p7uYqnlTGDnw42LkVEg2yccun3LTZw9r2aRjZPuP
TD9USRinD4n3nPCK6lC8G5hNsoFELe70wSBW79G2Ch4RvfbPt/vGGFF4dcX6ydVOSwEpycN0qbgN
odQQihy4xZir2CSqFQEG8SAWR6xN46H0/D3FQ0JcTynkOO7ZmJLa3WDVq91y/3Y3TQZqoGN+Dh7f
K1FfsUpdNeNbMNb/4DHqWFtN2UZiE0B+A2OsyP+DqujD/rgmZ4E6/XyU3c2uNOyqW7afkqAvip7X
k3bf2EAVV/0CWJ1THgykb4P1zewi0OHxuOwcHcsfR7SVoymJqRq1BlImuU2T3PLEWbGCUM6TzOJ2
r2XuK3OB8C4PQyRsqrkIVSQE6WKGqx/DKQVWP0zGHLIOGpfcdtf6SGA5V8hYm2nMrBdrCilhPwJF
5LKgDJ0DGayDSYqWlrXQMi+eiU5GI0YiEKh0XxWCarXgH+Bujp+ZlpccLnheo2AZLWtODgbHXENH
UejFToGTbzh/Lf/e8BQGkIb0s+3D/svHVEmV632GmVVNTSM69NPHIHUi7JDFWxPfxK8xdO/a8PxT
RZDpzuDB6FNin6ri4a4Rzccd4zYzvmbwbhOsWwrYjCxZJ13Av6V8qqjT6Uvj2TkQMndxoxa4dBzX
CMKtXrr20NZgBIlO08rW5qPTOE5n470+Gis77A2C2bpTgKqlJvHoFacYSuacx1nWeROg5XyOB6CT
BtXFEWtnW/u3ifG+RD9Qc+wkEoT+nbKCH41sjJqgSIWRC95t8dR870PO5pD9B4G1LBZLQN7I26Im
YgXoCP2lFS965RtqLaT72YYjYnIxi4uv5XNJ3k1rv7Dd+0vgd9pmqblp3KEQiVek3cyX4kFpo/Di
m1Q12UXBnJ5/Zfp7YXArAXAoQpXcs6Ct8atnT7MBGFU3O+o1tEQDOB+GVdL5MV25IQE/qpSsUpaB
dntBX6xuF2BZEtWYh3QUjuJftYqolb29r4tpCe+Y91zNt0qTUZP66aDybkotcOkBvr/jFFZkhd5P
I5N/oQSU4GIU4zYMS16k9n71IpzitSxrzRUPiofFvVQ+0E6/AuxwbVEMxfqVT7fYGXxXvY3U7xaI
IhVFbeEMBjMavlIKbePcWxy5bcKsSxm7w0YX8aDD/XZl4t0gKvVH4BWEQp9VvdXa3ck7GCFvFWd1
QoRQEplc9CExGWxFjkmjqFU0MvTdy51WPsfAaMWxxEfSwdJpESpXlwBQ+pJUFvMltc8tV8UiH/D2
tB2Huc/LYRZwuq2oWfYfdhf7ITCiZJtKnRtETpZN0KcXLhLc+x+fiym8/bnzY/mUCFZSJnwxxnOh
5fhsUCjWQVn7+XGYMyhJlc5MHi30dtyvPvG5SzaFVpiXpBpP6tURp5UwsLzGgH3dg3kJsfbyDbI3
mbAP8meauKU6o0PTMqhPJ6W8EOrjiiNG5bJUqYMO+8KltH19Jl/XYLQMZXduAdOWSBDHLMKMcoeG
tJBlaotc3Ryj/7djex7j/w8CpDCNv/IQay8Q1d3RRg4dDo7nERY4RmT9K4Q58jiweOQyVtjTLlxQ
ZxRRrAnDAahsMpoAS63tfpjm0b4DynxBttS2XjXthOGORFRZVh0SAIEW4vvl/iB5L+obQlQFp2aX
RLrZmAaynBUT+LUDwehcKA3fWHT9LZ4z3DnG0cQfFkGx8r67l20SeFX3Q2WEiJceG2olXxsesvk6
Tc0n2T4tque9K49WnczHlRD1fkupvkirOf+CS7NnwrJsER78G4zMjZUxKaJfyaskMyMNhW9TdAjf
T3PjzmTR3aTZR5zXkDv2ebKvgSAROe9CI6mAdtFMI4ITvTlEzJVSeRZgp1FymAl7mVdWQ2/hOGEF
VQH4HBv3b9T8NS5A1UzVUC2+inmFgQpXSrMqjt3jWaQsIBaO3MLG1stTb51m3HoIrKnjOq31+Syf
u7SELegpvqbE3x9a3BYWtHRQQkGnfSM3zXcf5KSlxkeXNZbraBlsmy3P1RoTLve1yT/7ZiWcGxfi
Q5V3WKczuknUxli7v7gLYOzU8Z4aaInLYqvYiguZ0xm1wGoN33RZ4+AEcOIJ1eOsaWzf3tL2fEEr
tKin0emiQRB33bZs16f2IifdJXICKIc+lUe8NBTHbTso+ayUDbYxzoRn/0WWeifCrnQcGQtsgRBS
vS1bsPmhZ5KQKP5dUt5JIxSHRLJDQDabVBb7QM6f2m+gf53LcuRzDSi/3nv3fg7HK7GAt1xmDtUC
hFEb3gtitrOa3jGYSF8OOluTdZny76nOHgay4lTHBwDNKHcUZXmIooU8LpAPx5RgFDlJ5omSfb/F
1HleE7yHOAVkRasChhnKajEDq1v/8uHmvPAr4qJ3Uuu6LGh5k1Fx25mpKxpl5QYAfDgoniZkujA+
9iTBOLZAA3jRWq2b6y/uoEB+AxN3KuA3D9VYcMXXPQLVUSe+lnTUI64lgqb6XBLSHyUyt+NmYvK4
/qgHfxgY6J/JzPu/lmebtqhV5oL828yd1rlnEw6aZHcqV/GSR2Rr8DTHFB12vjKq6JpWKeTPRLuC
Ymt7JZJfGULVznfbIYgHG92uBtyssu1vC2Aoyj6F4mGcYdfEhQdJu1fc9NTczbSN2Vefd7BQ80pi
TjiF2K1rmMH85BD6xEPw7kM9YIbYBdjricUBFygQzUh9SJEQCvyGaS2QzvYz2llv/Y/FLL4bO2Ks
2ALONVFUOvTzVBOoezeVOyq828pdJ5QMQOrQl86la0ON5aBQf/yOhN/Z44055TYp9Or2Sfyi+SZl
E/q6BZWTQvubtAOAXTxH1SJvypi71r3BmrHQg63ovZgNX36IWBPiYlJijNO7hSmadO0mi85T5Ysj
AmQDW5GGZCNDkZ0XKqguqZXF0IqWe4nMV9/tNjdx8kg2DZYVaUKyjczQu6x2GhRx3Eb+GMwT1YgS
UzogxHVr0zbhQeNpZ86rV5HCXtKWOsD7iGXLYW8okWYTkbqA6Ml5WwJbG2dI59EeGrLqzsYQRBjD
IzZ4xgBC5oUiXVywgoLzLG5+kq2hxVMmaqPXOy8hxAdXvliov6qvWaQ44lFjtlh7toe9isc2ZI22
cbmUwVGj3rtZ3O4eON+ooyu/ZPQTCsrL4wcvYBfCoJSFJix979kFUeazdfKOHl8jifhzp1yEGr0c
mgQ4yfiKm7S4J16wIFwmJ4nHeXM7uY/DYBf6QKLheweKNtErx6uvUSr06V9Rl5Tqa7fVbsABp8ap
EKNasGsYkUrcPI4qzhKZajVLqlfgjScc3ek4xcM0M0fYfb7IlYYhmXQWx7sX32WgsKmNtZWMaYJ6
qEz5gEhFyweY849eoelYj2XEca7YxEZk9qtMJcjRYDcyfM5tCgcOoBPolhOnC5W+kmJOvM1SXKBJ
WGkHt7dHBadj/E7EJAD/gRtumTPfVi3IppV55kuRATCLOPccGPjbrmt7O7zDkMw6G9JEkaKjtobQ
PNve0psQuV9Z7fulvYdFAShqMwj4/I7acSaxM3YFkfMrzUEJv91t+6O9HirEcda7Lx/tIp4hXG7B
3/kOYyiOzVGP3+/t66Hj3lMlSaGqZmJto5E07sjuHGlbqRTVoGaOS9Lk30ZMqQywtDikrqi38SxH
L7PLHt/eyFjwa56IlWA2+VEGCux/NM/M2JCSWY4yHf2t5xJT2WM3HLqWTthTKS/HcdM8YL12wyxU
l4pSIbK//g+xNeHqinf1HhBQl7yDyaGV7IYoHFQwwlNk9QPQ0xUPyr86ovJUBrDL3KuD7X3su6vo
LoGlUKTVCPKCgD3HZDE86eF1UEGoNo4VodDBmszK7C2q6x/f9Q1MPFN4MLH/YXOXZcQ32EC0Mgpl
85KrMhXMxoSdJYKi1kpP9vxLQ9qqbyN/W1+EmHhlQbma1O5JiN57TxxkrziuaXSuj0qWx0JqTTXM
rhqbiBRE00Lbsm2zeaNHtFJKg7xyFE+cskr7jTTbzwy2YWH9dcvQ4WLnQ3JTLQinXLNqE9yp3Q8k
EhntpF3X1ODZqNXz6LrtU0HMhe2xzlC0BPmlSVNOJar6S2m3LIMS8++U9p/p9CDD5n3Nwfv2SWSA
2dZ5ogBkmyDdxGYvQOYiTD07KJofsGIAQezYZtxfAQWpU/D6ERiKJ3AqQf/AQfQkSekRKizXMsbh
hredKjv6/uwdpp5DCOVIYSXI3mJ4rSAZPdZWBlX3UOwh6bPcn0WVR5t0IKfPR5iYzsYQsuwJcVfF
tKv4k3KR2ztBRD1eTdoKSzZS5PWaq1lJV+xujWUhPujexmgkqxhO5rVV8jPNsIzasHYy0utxKjxD
SzHRN/TQZ2uaFYntMpmwppJ3708NXnarMV4AQmaasnMnQQlw91KjrVk3eXzFzfHAdMSAtduGNCpb
TD/KGxKVsQD5Y122/Oh/fNx1P+CVHRHZNCxmiGdOsTDSmb0CaXmN8K6cTuPnoRIKFJMf4Slcf6Se
dD+x2eVYwEqVLR/FMCTkMS7zamn28FwZ5wF8hp2TkVnzurF2hH8OqJJRqXy+b5nj0bIRnCru/dyn
BoC5VwZf2hTLUiygUSrxW/tMTRtMMgTfKhOgzZ0n5KrEbOVHsjHzss6YyRuYPLVzLK8IGL+iBt21
Yo+uFpExykF1jX/8ifMqEwVuWvV68zDJHL7L5Pm2RzxOiTl8rjKFd9E4uV0HYsSly7F6k3NMPYub
BOMnkIab968ZW3PvNe7n1dybrN6NjXIY6k7daqoTm4foJ7a/XT+3L8U2IQruMheXz4lFo9Rgugju
51N15d0w25A3BVD+Y1bL6yfJoc6T3t0z16Fno9GEYGsS+bGDscwV2ceIDBrKjw3ZnVnqH6Q34YL3
OqdQI0V6VoWU0LL0afcgwBp/RlUHLXrkFzYv2x8PJS5ebr2UHGdoi8rfUNSKiS/PIfHDoXd/U3V1
Ncea/fsEW93Z6zux0dk+SPhM8BwTmTOHxGnkHMjiQq9f5jDtIrMkskgRnyfK09ceQVNFCK/c39N/
CkNB2J1PC0Z0pDxdVsKCWh/bqeZ95KYkuU4MMNZWPeC2rXiG3f6Fy01j3XcATcavcMu68YVQsfQ+
eyZqLi34s5cKYh0tMAY0968+/ezG1hK+RGpqMGVNT2g57nx7yuFCnmP7FPTYfvU6jbq/d/EqsAo7
IfQNahXymaT4/e0+wZsewiHpFDaC4+xKVoKS2M6SaOfD1NdASj/OErGOJyjNb5UYmmn8d5/1WDab
vtAuMrLHlb9oQioKbeGUqneDylrYhO6u5j8GT/mF+CDnoU+Q/x3Ym/w2/9+Yg4xSC2zy8CsiAk5j
Iomu3QaTIPZCSpGpUrbV87jTBrrPTN5QU27AoL+LJ98HWsTh665qWvjMe4XESRZY4ZWFywKE1dTt
boTHc6/LDux5biOnd0q2AmhMwK+5FtKaAyx+PMBffyXR0fbKrk71poa48CSuVqIWSacBfBAw+XpN
+sN1rqkgAT8lg1/poayPIh6Pav2Z6YllZdb04OeIZxiWkbl3XUvtSBbZp4QCeASC58x7aGddtCwR
4q6WX/0KoUvkAfoWHNXiO0hsjq3/RK8+cj9ElSthivVt859GPlgc/RS51zPCxAkw/eNA1rGC5vAa
RdmPIpwPbrg0N246+yu0tgYDXUrblozXDd13p/zMa0L+gLLFaRQBDw1LGN/axfgDLIKJLZLK1yLp
STkdOG91w665FPSCWit20jzvCnOXROsELnKVEdwP80FenQ+DTvlF99w2g5MpzbImTPQziiTRj2xH
0pYyt3YnRA5YOp7nKMo6wzmbB6cYzW5wHAkqyH31i1RRpV0UUkRFBTdCo7sp5VJpOuLJ5Yx4quMZ
pm6X2ww7EL4Ra+LB5i6d5CKlonXIHuy2gtmF8WWrzmGjS6ePzXLC0PxKuEv0p4HOUR9IKtdnFeUc
TG9WU8LyQn0i0zFSsJ1MKAfmsQZe7ZbFkhgrF9HbhnsRaw0HRvDiDqCIclzxAOSpykfnOGMQ+gyX
R5MEBkmMFgv8a7ApJj2EW2cM7kFqvLZOlu3mkbl7aoInLykbSCfZbHih7KmCUk9Ws9XnjLIX6ppB
DGF2f5/tNsIqfCmaD0eF+nNpsU/yUiVxQSxKt9n9Gj/4Pbb7+PkYhPfRg6HJqvI/abGV1agz/X9m
otBylIAh1J7vh/94DndH7BLqy+MMrQMGUimePPemc+iehVKGwqQMXnoR/C0atQ7XG1jpVOrPgy4V
9Zh1iu5/1BOhox6rYWAkQmaPJfnZ2+Sog85OEg3Kf6gR9xWNWFW14fRURTiy+/4tf13KnotQK0xo
Efgv1bsW/bFg1R12jANunDac05WJFeXc7f7FryzQWwmcsHGbnaBQa/6Uve3VLjDFRLWRAEUjCmGw
6WwIZs0/n8rthEV1RZ0+VBgGxJ5p/nzo6RVf8MHHQkNV8XbgcscTXT5/c76bV5aQmp0qhGsnc2Zu
OLyWg/6jgxG1kuNlsEawYB3kEqWJXcqrsF7+adBpcoP+me/jaURCJRqj4yaDsdPhS7ajTuVJ7PcS
TxnEjSN6quXuqpqceXZaeJAuM7yNkRBHoLAtw2zACOt5RHwCHR+nvyYaQeLZbx1h4tbF1foou9BL
thdQ7+7Iar4mix3+i8wF5c/G5Dpqvy4FnBrVQYqlOZxis3qkm5tiMjhVE8KqvsZyY/UY6N7ZdqQe
ixnByxZvFYopHULq5cfMjefIU/BwuTCbkKFxIoRV8iSHV1y1YjVbfLZf1kfuXN5UMtyXB9Yf9KIp
kmMqdorURzgTSJuHLzlW3MGi/IkD/LSKw6Z9KWQudIkd5KA7gV/yN2GpfDDyssfsPtrRJcxW2S1Y
Ex3Ygm6c7szhbCsaGOlG8H+Ag2rrm7BAACtSfS0vTs/1SG18+iKeYS2HcwRKyyVZzNWr1UjGze+t
2Ashwuq/EI7Llj7prssWTW7MTtCywPPYurlJzGvIL36Ub93W3zAnnhUJd77bU7TUlP3iljVGlKNe
STddll64ATtTmPS7SXLjkZMq88QKB9xVucEfqDioV9jFtM50fM33O8SsQyA3U6ED/qp9euwReBvt
Ss0jSSyJsS0nfRnJqvb8dv3CpuDUg8tuuSsoeF9UnahQWizmyJd7m13aELXJcaIyl1puXcx0qtDU
FwOga/gCWUQ+TC2QUNvghHLBzlaeUcodabZrTtg2qKqnDlHEAjH6LHcXoo63izZA4KGUNTFSq/PJ
p/dZhqeVGtPixqxMjoTnuq78qfjc0byxbrmhmIXg24pza0knq5oOlgTjCLFSl0fcH71htu0jEqi/
BpbxiXQqjuHjrgtel6O+JxBfXkt8icqcQrDvhAljXiHgbHwBea61q5H1sRwW4n1Kw3RJ3pIK+HGa
Dh4k++2Oz5yWEi24VxM6faySPJMkAobiJABXCkIHQis4tnRN/mn0MzihXCjpgJ9k6JMuki9upD1v
9CSKJdcOs+Riz6XcVQ4BTdshpD0tgTvF8L5jL4NqHlPSsdGcc/jPQ7DG7BNZhpRwt0ixZ6uxRhdk
6/2UM6qnt4aH7Qh9Zv/kHNw+93PsXnh2dSkr55RcLLrhXWVsq28ugU/IgyUjzICQIVrnmaFuhUdb
Qlvv5hJk1paGOTKplamTg1BXoUqIREHxyeFXtqtVFsC1ZiYjTyAOe4FEoGEnlLh/ZtCQZKj0CN/h
VIoJfEvwbkDXM60oRT61qCPsx04u9ORxGwlodVasUldKC8gnrkQcBTTu1SDJXXw/wfN/9anm1w3q
NsAakjKhvJ1StTZHiQ2kqZrYfMC2aedrgZgXtNsUkEhuLS+EyEzd6vqRkxit7XQ7VnjtdxGjgql+
qaV/7Ugj9MRvLH0XFJk2oWJ39kSzmtpm+EUTnYyDW/3IVKtQmZOV8Mbg5CtHtakP5LwM/Fm6fhaY
HYPT1bDC2VLa4vRwOodEVcBLP70ffy4RH+dSvv6MX09fZcSS+lli76KfSpSFe7H1TkNfeB5kfOIx
lp3SGN3DdQ02HZ7lak8DqIFRg0kMzFi/2ACVi9+G3HW6TWJfToCqE38HjMTmBe7G/j1B50sMKRF7
6mZrZVUY/yqSyOE5v1Mey+QRp2s9/4RW0HYi2/Cp5yxRto0tWhdmlnJ9GW28MLOgo/5o9PkJAuq/
BSVu0zeoVag1UWq7SVdmxPa2WiAiWP6WfvStJIWq+S88PagWPz+bS61AmsEDCwquvQ634ijXxOx6
KnL+9Gqb98fdmjQxU2QMT0CTX0u7ExwI+wMix0xpuflrhLjUAbI1GgIbT3LjNWuFEBQcD4Q0nZ7W
rl6rrAKnOLgv3AFUV3ou+dxcGrgM2cvZXVQQI3XbewzT5h598SadlHHy2d+ZUnyRpNJ4PSBHUtUN
k+3F61sdxtd4FxnjfzUHTZRxSrpVV3mnAtUuTV8TQnlvE01k8FgdwkaGwfAp68XNZLUj89ScYzrI
XloeDj71G92+lXWHYKU+QiUa1tOfieQr/0e5EPiBxzLxQXqRK5j0hBIYm7MI9787WWIXW51xOGqM
AspOzufaeuoCR4j7KVfnghoZzM07dh7O2+ABne5ffRNqe0deMLaM1e7NFqu2JdzZd2XzH2g84tRq
TZRw/bHfdyXI5EL9Q6E6A1P3sMpWPiBbxl6WZaNuE5RmacJMorw1YpmY106f8WAYqNUFmtkTsK0O
Wh7/ggxepPtLNQho/U1bsdYIy/sGE9/694Yg7eoLWodIhDv+qWJoG1NOx2XWZ3vi6yTXb/eV55CR
KBgaq0g+UlFkBWeNDrjNX8kr8mZRrbimm3MKoIODrHGvRlbFW1/RMtZTjf/C9GMHVvjdcaynvhTD
3xSlndHcu/g/+Eg1HbHg4fQ3aX3H2FBjq4YIcGVSk/M4J6kMCCVL0hBUyaM7OHAxIy1WersV95Ev
A+i7SbxLi6cbeeTontiOhf14DrPZ9Ce8bhvzO8Qb/wiHnQ5erMpt729OjxhgwWesDe40Y3DDF0v/
4GY6TY4m+eCjjpJ2knkFjFrizhQWUuHnrh0RWmYiZMnJ4tWPPUtXxcmi45+c0gp0ncZvLypEjyu8
VpZm36fP5xnfUSjyQ+OW+nUtlIxhFUBlWQy48WPaxGPTg2Rwpcd42R97XeGTvAZwf0XnKlTiGx5z
hjS/wwpC9r37ILpx9Gp4TAYp3Zt8KTENenboXGFj1L6Y4cz9tTrd4skLOB1m2AyllqGgkpsL+AEr
SmOUl2ZnsJ/ewFkUcigLr3++UvZ0lB8/sItcIzeJtjPfwrlasNaIE9RAV7pm1pZf85cQr2/D4t+n
JwdAYjo9bIGyncCcgCgnrNdfrwmcv0vypIjyMuGHquoKddvffdiZ1FpIcGmztpvaM7BMIJlZPAyN
ZPqJBZ/3DXAKFh3SxBC/c1WV1QkzvVB4qeH1P2/hb25NGO2Z8BDozHfCrD0Hmdb88ZfqvFwYKuEI
/KhTa9tFHjiDYf3FvmmxU9Pkp11ZPi/ahie5d18EKokF2yqtuTRxhCmshClK7kIur7A1sPx8Dt2a
L3CR1Bd/8gkoEwtS3iDutDjNw93+D//bjCy6qg8nzaXIfmUWN6Uz5fvf4YhZf8Y6xuYjMZMe5dgu
9+SouNsdyGWcIcSlWulR9adaQoyxlKEtiEzVSL+D2Vhe/bGH0mWdf8LXdJIdcldFZSJXH7d3E0TM
vfgQf05dgCeO8wKF6+hmuXH+9zfa+w4rnrTvJKWNBPhZUcBbOVYp6BbY40jeXw6seAK8RqCHQASk
JkjjJBTPYikbGDOROxqvSE6Medz6D/+Ec3NbccQyLiDDeLOIJ+zTUuFetstRXPVthVORSxqSUBoc
P0JJJ6Qt6rSZaI2MFybgKzmY+wVlZfNISQMT5mIAicieePFagGJ4LJza/4b25ze+90m7he1hXxzp
j8mu0S4h57wjxNSw6azk5WOc6XkiPm63liqHcbwFXry7qLCsyaxNP7Ik5kegEHnU7SRtQD5zircB
wpRToyczPBLBJUv1BFthPBoU4m59sZi1yCqS3P3Lh+rfd95Zio3luQZocm6NKIL/bU6pYXodfni1
YzZkEkMqmEV1dFzh3dGxj0LbCWagHtvUNNtKxZ3AoqDrrapoSBA5LXWNWRsnprtPBuHSQKVBoObx
r/56DnXzjl6oGOzUDD47BYb/bE4JfCLexyOk+3D3GM9X2FhQXrLNR6LQ2Dbf3ZiP7Y4+a/UazCBf
uk+Jvi41hC78Ntr7rki6dYNvcP8eqP1X7JRuq8CNoPKICYwU47XERVVKlO9izxhfQct5OLIx85BH
0T8I4xKNMSsLA1T9zHysoQmPdYthcsyurH8xiraC6vQ+T0XViYYuVlwx9zUbw5fqYDuCcV4Klh17
7/rmgLKYilh0Lgl2RDQopM3EZCldKCpohZDz7AjJy0KV7OV7PQbGbvmoaoGzWB/fCKECZB576Ybx
4MqdQ3k9sna75M0HAtWoUfogiIszq0bWYtNrGObPmwWA44t4+L8RgfIkNsMWcaK137FnfXFoFOTo
JPjggtmxwV48aWjK2Nvc5wz4lU6IvlHLCs6KOo+E0B/WgcQig5wbSeuF9NOm3s6efwZvbF0T6y0S
XEO9Xpk9tJhNGthEGaCkDtLRyTkJmVB0jC1hHuSvasU8EsNrckbvgoPT6wCh9MJ82GWlup0mVq5M
iDt7OFp5Zf7rwbBA0XYFsstS/1bD+Zp789Az/Q++JcgrNugQQBhhWpmQc4rFINRCmDjUfrw3SGXq
Ka6VHrLRdnwKLc3wMNqDqtHnlyZ5uUEmLqEdJ5Y9yXVM7c2r0vpAFjZnACY0/g/C6woX7rXN96Ya
8xD/IGojoJf94LT8+GUcRsq8Gb4PyjEfbonShJnRhFUyYcWRz8rCtE1kNO54hm8iljfAMq9RoEhz
Fp+P2CHp3Q0tpFeG1bR6hrytcDFBeHIIniV3jTj9i+xSennBMe0c1xOlYX0pDBz8gGDkDnhpFevQ
4ELTCe33DWzhxAzhfPPoBGkDoMTs2TKjGUKOzNgckSVYf3Q3az4UFwO+pfUDAXI/oNDuOq81ejhA
X8/srO0sWaovFxHfv20XiRKcwBwSMVAlX0CjgWwTthgFT+jVb/jsTgJUyzQbFiRqVcrssOYcxRJs
UbLjcKb9GE5tQI61ROKhEy6BEIpFggqRcy79ulw8Ym6DrcmUQl8cvI7Id+pePDtATaztqcyYL4at
kFA9eKLWG6lHXV0WziI1pw9eEK4RzBC6KNLRwmkxKgtZpgnPnIs8TwDqB7buVYOf9StlIbCOPV52
T50+vbXLVooYBMYCO1aC5iSD8sx5y4Z0lwS1mUd9Nbvy6jactqiOeIkMDK/XgdVoPuup8VuuGJQC
uSqWdBy5LYnbjILRLNV4B+skOW8NeADuCW07UwibPmr1VYc15J5heRUUSiMzBvyzu4ILYK7eKt3K
HWS5+hluYPEhOSG3mRSNe8uQBwUQCSSvcklK3P9vAYLsX06MVEaMxPil+FdRO15YEcqPjRpKBOLA
11z/VcfLZU8AXZT7zbnfvuZRiftf30v7SKHoj+ZrHishe9zuEaNzYcVW8XIVpTGa6Ni49VOCruPP
2yZ8WHlufel0TsbVE/Nkrap6Sv400zYJpmrTp3Jj4qo1+ccFoczwy9HWsdBOmHNmhFY6qyWNWQGU
6XLQZBShH30OzxFi4iK07gaVtyMhtNfgkqKL2tIuv6YINCXtAFyegUFB7X5DZSWZp/Xdc23VJ2qG
PzKjbkriWbE3p/n3E9cmGchFEv4i2jD0R4VDKemm8wvNdxBDxGGIxB42GsDDc8DmUOFzjf9su8Es
R92aDpq22mLju4rR7rO3iru4DZvDsx5nrkUAZK2zwVuhJ08gxgnj5cZf3QYjS8vS9GpwIqGLD+Xz
omZBszOURCFjN5ePHnCtkEBOeLbsb/sGXpmu8ywO3FvB2YJY3QGIQws3ELGV2Mvy4KppvO8Z3IFV
vnPe+sY26eM2QCKZG2N7kYmzGPXPywaX9FkxpzEN1+doGke/wt71l0mdGxp5n8md2ak6dIe20M4Y
ugyKO5Z2Kf/ZKcL/D/+t9y3RTSsH6g2MZHPx5E683WkdT2jrnIlS2rfU/ANgHz3HGXnhHFvzic7D
tGOwS9XbWMwPyEdqrCuQJP22qB+zQxIp/N65QyXtHC18QUZ6LDh3mTXNcT/lHEYQ0ilMMUrZ5Ntg
m+P3WmRNiqPSIPTR6cJ8z0LbYNvDkY441nLrPGH7Y24nOx2gzFMfWDd6ANRf/mbxT1JY4yTHtq4r
9z7/Vim/vNbE8rH4HlIx1dgQin30sWUhzI/rstlZNKZubrmtakUPOXF4Rjc8vaHBWGo4sl9SA37Z
xur7C4asH/d5jzxBPjaWOO69uQUk4zvwdyvo57E3dfa5NAB/5in7hqdzWUlEx21Gf6KF5RvqTuPT
ynrekhfo+2zkoP4+bMErjmeTCDwyBoaZ4s0VjG+9RtVqTBHDYeidO8g+MePffJ2prhKX81jKggvV
vrtB1qcwnDeeYn/n4aQ0cjqUEX1uBixXDGH0wEnAw/lmfXAozfFhIqtCOjp5Q/Fm9fNDT0lR0C/k
ozUG2Gdg1U2g3KwFXyTGWEV3Pii0eGIlPZGwPGKZeATvNW/JhfV5lQdDpAE8mVOkXWnmCJyoC+oY
NtS99zcejAlsYpBAMstV4u3CtbuhexcD8cp/zS190yi67pC7J+TvOCLNGGkXSPPv1B4YLt0+AXbk
ZC3ZQwPmLsCOsBPw6Az+V0NI/EhBEsEAq4SgsQkOV7wIqtaRdadlZNKma2e1Zge2PjNhNJh+KsYO
YHswC9UfcN2yBqW7l7ubTl4Iu3aOBhVYzmkeCHl1qqqFRbGxtIb3m2bmFjCZ0Tc0JrRmt/lMg0DH
/ufe7FqByU/VrPeV4ZKcHau5LIl5q00qwINYRx5hMtb32NZ0ZGWIiLKEu/wPHADZkbRVBFPDgEV+
d9XUKjK7VkfDE2jav2SytlfbjlCs/y7xEBEDfRKQ9aiHTUQlv3MXb1TL9qV22Mjkm1m9PM4SwAwR
Xfia59o28zHo2BlZ+vtk+Ju9IKmg6T20oN1gIVHGC4UU+EAiqn0dY9UkpuwDfri9I2jav8Ph/rLg
daMyarwf49rL9ju/OSMGlr8fSRnwrlOy+t26R224ldlim4ncxdMK5/0pqsCDk2Bj4q1OPY3E+bUP
bNdxeTKD6uSwPZqp08FNLBxU6lvpEP6IKY+ErLELsCTlVBfjDiHFe99KGMrRfE1+MozRHRu42kW+
soOvzkRt8dSPlGeZ0dYzpaIBjM0SaZbIq3ixOv6HoaMdBXjmguPq0Wk5DUD5hIQmGxc520hXrYzq
4WothQ1fwbvMPwHyKoZ+GyUOQ5pbV1sBHxnHd37NDKFL/k6syHREZfWKOHb6w0rxe8Uhe2zt+TBZ
xn78mg0AawkOJoV+57qFcVlu0/bwsO9vRPu5QzdCouF3jhXF4lZyZDGlBbZNieqY223DEP+89KZ8
zIoL07UR+24saPCZGSuThzaDaMot4K0ixf6gyW6FhSIXLR7am08OYeSo7B9BmCVhS9LLkt4+HDnQ
6NuHZ0AY3HpB24oOJ81CLYwjI3UJl1Dbuv2SJyF/CkZIZKDbTQXy9FFM9w7IeMJVgLxytrSZ20um
Ij2pKK3LLRqLIDR5nmQpbxPC7UXvvl9RzXeDJh3Ftz3oRqpvRw74DPfTUJ0mrg6qF8siwirQlhZI
lHStBC7/WM2bEzbVG70DiYBGRhEXfNi0P4jhTYukK1/7ORhHCJ7kWYaAY6XOYGk914cWGSTYgRM6
dHyCieVB7GvYm+iDLjZM/ZFIkUv/gc2zR6F7qFk/HU/VtP7HNHNxnDqvziZQAr4IYZqPmlIljevK
aaR8rx41+zY67MQPzmyARI42ac/rlX4mFWpoMx+ATrTv0s7xmAHdisKEskJ1+FW5Otvbc2+gSqoO
tSQwsNrcJ4DQQyaU9J9IUOYwtDcoGQ8MzUaxfDuNDEq0/MaUf5U5KgTZ+p/RkhXhxAFVuTfgCnsz
KNsVzNHwxdlD4aqVasxgSfpSNIUU7h3SF0+1YfDtGRskMEff1tOsQF7Ube8dzgnXUrJSgYotf+x5
qnXLbuUBuO+02+vjiYBtPjX5CZlPhnJcBzPG5wON6KI0oP+xVwGzPOaFzQn+Y/k1guQJfH69kRmR
qI5qOX8IWtYCmwlFlWfXCiTZU0WIJCeWoGqcyCg+iYFj2QnsSuDtqmPPKgRLaJfbk69qzVbwBbyk
RHwnpP5PpiY5reH3mTltypm5eyN0hNyLfvCFiLW8C3alFDWVeGvyCzfTzc10UfLzb9zDniwqvG8N
U2bgf6FQujDe/YSY7yZqI/sYohXhL961WvLUhLbjtCyP4EKofgTgyjKDjuKRRjhbtyAMB/If8Osw
D7fJhnzIFlMvCIcoaTBo0JtN/X1Ze4zNWibm5NTdd7TuVCIHMYggsvxuPd+YKw17Scp6oNZJ9TXJ
V0gmhwws/d0b6OEDI98nYMmrwNF/XIFbPglDYcvAXEXYozoAvZF66ICMjYkIm3RWR8oCaz8tb9F8
ppV66+qFcFaLCtAlWEMWWc5NGpW3/jJ1b68TZCMF9vmRvf/MPrJih4IkZHFudphX4qAetru7wpAK
YSHZb8iiFVD512mLRYXvhgmmj0qFAcjJ4VBw37pLNQdHF2mdgMiTHvxVviZAxySt0rCspQzffcJn
xDQQmP8124KpK28jcJdhZF10O2aEMVVLGfmEgV13LmHR5t2I/U5zJssZu7ahd3XFtn0X63Kvtwvi
QUuqFCRswk6ePqk8qhua+KI+PNlPP6vkm0JHnAQIjMBWFd2Q5MSpSdfdhFtBrjn3fOnoFUjwbTMV
JRQzuJF75neSqlDAapp+tdFUjAUbsSmrUZGTTnbulnuHCYtZGiAFgk+soX0tJotfadxbv6AQe5K8
JRevcVvW6vdl81ilqvwzNYqI99p1eAOKtWeo5L44oQ/jh6ZDvtWmz3ErXKMKrO8zWDhYlKDqElpE
pCCWJd85MaGukrGCqMnw7mpT11zoYk5O+Pn002h9BxEQMkDqdcdM83IlmqMMlZkqYt6kYWgFuMgx
hZiIBniTykGkga9Vdb3VrnI/cdN2mpSM/bIWgsdOUOXZJD/C6YGqCEJwlpNTiARUy4EOGXRp3HvY
AQRxk3UnEVOLLEGK3T2BAwR3KGukdRGvsu4DscJm9oqQGHuKqqwFr/uIbFZPpNHWP2zVSPta2ESp
j8yPkxumDHP//WK5XUW8oA9a/vF4BXfICkKXx/fJIJ79PHnIRCbTCHrffYZ84owHCFX9HGTyfhwa
6Ssz7ZAciUk0gJA0HW5t7cB+sTUlya4Nm9ulkvjBq3vpvZ1FRWWAWm+r/azb8aJTjlciFKgY55Nl
kYHNKndBXH1pJ4pCyobO1uFcJ8BhtxqiN7NkU3OYEScpn+EPo7mz11/ErzmYvMozM699wnqSZaBB
FKzVR18xHxgopm72wK0EPxjVGHWEu5jUuTg5BU6nRMwyMK8W/5jjbJplm18l6vTQP9McnzYNBAos
SV90SZJQSB/K2yIMcnUmSdNiNkVcdrWruvPX6qAs9an6LHSRExfdL3yCylz0v5a0KCxbyo3shuSV
Qwa1+JQ2DuCyHJzQo1uimMJEKWkDhgK88ySh5QFSiaGMV5OrtgcheoK/3ipjudDvw8SsxezdVw7j
pVAC7I2Nic6zwFkGAOnPcnXJvr55xKWB33lZjHoLc3dDPL9yWbfY6+JBY9mYgodhzUNTf9Is2Nll
n4SWOIqoFJBnSnXoUBGFGpayKeazIs+X8yQJdQUplN8rxBnHQBBB6LBucxNKuoBXJfQxEfafDI6/
IFKdtqxQTPbMeNk1TSo410wtBaF/bm+ZrfvgN/Wqhe4jbbw5doceneiGZqJNn2QIid6bNslBXof8
Qag/LB6G46JGNMMs2uZGqy7+29z3biP0RFcjSou+ocQ8rhOGPEdWsbmQxdjW8gmRBHBjgY9LCBvf
nqxT04yNlJpWBlmQG9wA06ihlXHrV5BNwvp36fPZ8UNS3/CU56ku01Pq4+HLaOnSyRrCCub/Hqsb
VsuTapPBy+rA7537mjsNq+IcrloPU73dLFFi3FkBr6rEtztvPwpzHt5SnYaGqZDoZHRLpyNbciC2
qObLzvUYMm1yB0HpS/YsCADacuLK5sRIZwTIu/aVstlqCTzvNxwfscIctxnbBslcXbiLcxQ7drrL
YEsj/8kPwbrfArPPaJKJWPxhByMynqpgagh4jsstvOURXGPUW8d5/dJSh9NH7JOQTVSeFeQnKDUO
MPOvjmjhoPYagi7LE0TwRQTlLe5p97Rwozkj4LSk+jIs2YMoxueBYPWTbQXMJJrUcKQ725GG3lir
fyUQ62yHNbIdoQYM4mtaIEXJmgy65XdkPI8gfDrpkw/pym0ybQaXiI9chJUo6QgNCg0QMesAz7Te
S77L/ui8JT9FiG8kp3rcXMuahfFUX/17Tq7rKQ7eXbNjO1njb4spo8GqS3VGZDenuGcfqqBbgYs9
CDi5CIPs2PHkYH0n/yXzMm/nvOjzNn8YNmdfJBaMrvVY8zK/ga1pkOVM+igDnRd5hlhYMSvJ1Ez+
YlaCUB6jGm7x/3bngXneon1L8GCQ8lsrK64EGtFHB2UPctyoWa9FESdYTSA3VLjbv4VUqVNse1iA
RvHZyoNfioEbk6P1g5YTcFzEI4F/I14cUG09iiXVapgKiqC05+vj+gE42pPzlYwE0Ra9wvhVHgQT
iBZ96hnqvQGduRrfxJUF4MkbsYcfkSmi+OC77w2tGj4Ycb9PurGGw5+57WzHo7oQjzYLBFSf4jCT
k07XYt/TMV8p5ZdRwHyxfJTUaJmzgQLP86rAjtUEEfax+vmk7lMWRYwgLMbztvo73DT38cucLv8/
hzJueS+xFmi/5aYW0VBlTsreeHeAR+em3jBYlTGuYzh5G2ruky+zL54bC7GMKUsKp/0xnOQYmvFh
ITQSgmSUaQy4NURF+gKWJt6Z0axeOKTm/fwRYIjpOp4pTnxbv4xfSVQFrtebyZ6qqRdx2gtEtmEH
0nSmqPFmb0XY64FDdlxjvnM/32wYgm4yvM7F1m4xOPGcesCdxkkKVbKJM2XgW4+HMLDE6w/BZg9D
RpxbDFDZfDB25rymXmkpMNYImuawUzE9kz4/nbyoK6XqrHdzrKjsIACeuGEMbZS2GUXQmhCugk4q
h0CNXxvbMqT9Vb780Nk4W0OWrcE346VcwYi9tuXta0P9GihxW9u+WPwMevZme+C45btswlrpbijh
vMyc5+Kpm1ViQjFcdObIVIMHMNjF28oYH8L9l9KZBIj0tJTsuWflDf+mpi6iqCTdANJXfQFCbmKF
3ZZWZ8qEfECxtaQtAH0EvKuYqJD0lsRC5ALfB2Bw/flEoh6gO/2ZTFyF4Sh1D+L3/KUGQJP2fw37
7c9FIOqMr4wexeyJ1UTTHHkAFpI/G0ul1LEtONiOaOCwgNIajAW+4DapNujiwgVcj2injEeG8l7c
F76ASqu8NMl/01LgTh3GqotB3zj9jZjC35Vdg0S2JijVl+XtK0I2Wmdr2pfaFB5fdzFQkT3gB5NH
R1lwWE4RUjTTAG90b0KmdRjxFmSS5LNS/V/V5b+SVF2zOSXtH3v6Mm6bc9kc1ihZ+LIv7EohdoaI
lRxvE0KjwKgVt/7cQTa7GTE9wBe7RuM4d37p1x331AcE5tINVNF/e9ZjOdyvBEQJdxJgQRTTrBf2
LXwBXr+tdzBglyfKIsj1QncXQf3FvsB4TimDEbJ9ZJ9jqHyh0xsSL/UPIKEd3DY+uushYG/dh6HL
48yZG/+1+xT86J6ZK6gOv9O/e81RjZ54x28loLSXKx8FKMClvN/ULcWwBhsg0JRgWrSmwUM6LD2q
CyqdN15RUyY7hwQvzZ/KDhpFGWi0DVVAIQWyM1QhYRB7IgakBmKTJmt9GVDOezHKf7sNdJYRY3H5
I3S+AlOX/5G8G1sn5o5a2I2Nsichr3k8a8cgUrmlXGXDE1DB9Ub8tf2Q7WeFUMJ6jIi46xw2mNZe
CZaANH/X+XsCiOZZEgtECkarVeqEwKyix9r7m0cwlHgA2n/i85ZzHfci8vUP2KbfR6cN7LOuk145
fPLFB1AN1Dn/XFrLOITGQ6Q8q+4uQYPuWEjD//luqRsB3WBA1dWVIeqBLm0sRW1YvB9YvkgbGUGD
HxksUXYudTa3D0cxzoh7u/mlw3obfRA9wkXDZQqNBIwM691rIri+xfyuS6NI5J6oUEObGWXJNHxq
+w3sveBDbRQGhQJZ94JyPGXN0QY6tLWBIpyhxWVivtCM+skK9AaarAbDCaTWdCce+dKLpeyIRFe0
tIMM+Kx3NQtDqwLgIQLXKYmP14Kr47P6WUzOC092Y8qxR3S5wfdlZt5hTkduxujsOYlsBmhKoCm5
u9bxENms0mMPXXwZrFvffL1fHwPnV/eajPVbdCwPGIvclmR61h4i5+GF81FerIer+8jltzoGwJYe
jK+1Aj8DktJMp/+uNjSjDXE6RWEMgCasMX7qmLuUvvKnJIOxbPa8jvIKI6F5lzkD6cW1oql59wdr
xRl7wleNPYSYxCiizHjmHYnsF+WjuVpiTIaqpsm/CMR5Sv8Ycy2IMB+mtR+SuQyF+kgEw8mBIAx9
evGL9hEy37J+OvZDyy1dlOOQk32dBObft7qaixlRlp2HgsIenv+U04mUT4srbAydxfRADS5k0x1y
IwReGHVgrAe+LrdvAis5z3QqJT75ilwdohQRHJi6f/U6KCmM8lMfpZ1eeBHFVfOoVzAvbU6WgSYY
ebSG4KvMalYsyOZKKVx1q8y4MwPaMNR7OOjIXvzr15y04mClRR4hcO6ah0ahq+/yAjsMpqH3n2AG
F11sDv9rvLuznYJk1SdpMybsgkeZrIyYJSInvmYp+NtNv8NMHcDcn78Iw39E036vwdV//v0G50Dx
11KDukuoi8Bc+lr88R6Gs4C5rqM8MA4tynmyfWOgKcVXsO6xh+11k9M6xJFnaD/1aUES9FJIGNTF
KgY+OPR2bLxa55Uh2yP7ZEM0u299kUDj6GCRuv0bK3c8+tRILh/ZOL4wTv+Ehc0oQGnSVZmzyVEz
v45OG6Be61PXlsZkvCAKzVcI0dibm9utcGgpAr4iZtoUhFRfAXPyGOZy58x2pIaRTGbt0QtwTz/7
I0Gty2oQ1gj0i5knl8G9V2wBElE7VlRHbQ4BHlf27sXJdUp3LVY3tcWDcrsWP1GTIsFeci308Uye
pG2Sq+1Ff3sYphwy2DDw4r37klg64XqGXynOl0iujZ5gdJbqtOWPOJ0nHru5ot34ug5eI4UIgW7K
YXdFTcSUpNZstXD5hZ7Ec8G3rFL6whMxWQ5aUXZ/SGZQIlMnLeRWrPeR3d4C7AhatwIzi2nTMFc9
HZiFUAHo3oakTfHiSW4rKZfPx10Sz6ic3LW6+aw6QtxNC1gmj0FPuG52G2jx28/zY2+KuGCdIccb
p00ig1OY+fgyit8N5wUVMu1P3a98PIrIDUj67uXpx1aCUPCfKM4Hu3a1NplCbjZj3Lv4yWyNGVcw
YQaqPU7lwTF1XaGJRSxJA4NLy59T2Ju2ZMWQavTy8wAJYk9J3yuU2fndz4s4nl4HvIwVw9Mw38Mb
Yc/mdV/YB8WAsQUa6anRqTh68rGPuTCtXxQhcppHM/U+3aZ8rtCudPbcMDSSpgg0pghHF7hXyWkh
wQ2VtrLBaDQfIZKquSg0GpfgXqZOaW4gNVSPoMKjsgduJ2LKKfvMryRwRau13Q91S6n5gp26ZHHr
XnvDpon9sU8Iy7js92DFoH4WGnFSp3js0s2Y/r/hRWJOgGzDhBJAkYisBOC5m65wdtgS2AFEJuR/
iS0Vk7C4/bbKvE2Q/nd6E/fKWYadagutVxImXMRTDZT3NRMSwjDcEsJH4GUCP3Zvrs3qGS0DrgHo
9x3YpgtyztPIbmTMNuoGDnEPYgrvL66NmGjw6zL1m0uqvA468kBFpT6Ffu8nT5W0ApAFKowIaV4G
rT2/DF4xyVXktjFFcqDpxcfp5C7XE5vhy0NosaN3hs5qsRcavk6GrRPMr7zrCqoh3ReVYZzH+AkG
oAhOwJuudcjTghfWUNhId9Ue3Q7T0koSWnMXCIvvJnfDiY9kazqhwELLr/P4XBb9kiN+2AMIqMRp
f8UEJNL5I+ZIhgdvs8qIgL9Gqy6J65FM6ziCYgR6p4XZmeSmAWSXRqTNVh/w2NyMSZ8G7I0F6uje
qoBaEHzRHrfezFeNg02vCG70fCkZWNu3H5pg35e+znYHDvrJF8xHVYvsuCHzcynQfSg1U6LHnTyZ
GPi3i+3iqjpYiQAmlXFygsMeA2O3yrSErRyu/Hx5XyMe/K85hwD586Q3XG03juLAX3XDq7xKySTx
20ToVOJ7pL/VJumKAknkG3I9whnMGzLkAc8aARgUsf2IxdKKZ6TVByRGpJm4fbElBedSwL4oA6VG
H5ueou8zauvsyYMPdUUD0o39UcoLc4GAB1xjFXF2hpdvt+s4Jvdun7GU0yz2IvIhFRp6nwwmx4YV
g5/017qwVr/mmkwOw2sUHl4MQubcE/nKoWgDHcvPgPNMAELlkwnckR5/uV3f3EZ5QvG4Dgg+6gCH
LhtvK6P7RocISldw/YmUn1twkgpawd6msnbORpJXfE1pcoiWieYMKyoBL8pFcjz7YnVu+UU2s8oD
y4WVqbBPRaXPo0ex1tzug1uqEMH7kt+GQqB01pqQ2O81uz3rTuSXQJ9wlN3WzpeMcP+3k/VUJ2gR
8pXCJWv+ybRgPvW7rqlLRMyDhr3cLLr88DQ9XO2R+BKKScqpqdzCG2jUgAbxBJeyVp1gv0G9PsE9
RDGISC6q4Yt6/Dp47TDiLST6nGcH7Dbl5Y/hKGLhjHVniweaJnKjNzfilK3jdTd/IPU+SaOgC9so
zj/ukWX68kKWSE5x4CK3TTcoFmVocylvZM7+H+v6zgPqPP2MSC1kPxveQGRZUgu8EbXtUIgIQFXa
bk3KuGxisezOgdk3IRTRmzMHh1KHnlTV9GHuKrYzx/yImenlG3t0XOzHcQk551I4Hy02N3fcYDie
oCmYb0o1t7AiZzijxTpCNudzzk8pBlPk8r4IxzOVKqDTgEcnKCR15+j80EoOHqNUTVVrHqx0VPUN
3VzzsAqtUz6CUYYZ1g3XUi+gGsVlH/C3Bik/yAwFPaM0cyN1IAHNwqD4z+VgIDzXBboODW+gjEc3
B00vevwjLvrYxluVkCeHfEKNQbMy6AJ/2hbA7kpvABHkyQwcNGuDbnt7KHKHSQWTLTS9M8k3rxFt
PpL/ge/Ys1uyRXKi2lUyCO8ov/wjBRjC3KvBWUn7cZnXFM1433Lb2MCSkYfBRvoYXJSW6jKPbo6u
HW/MvF+Bt91H5DBwCjodqbHt/IqN/vf7PETysd/AxgccvcxF/h/xiFAb7TDRd/RS6O76VGL4bWVU
3g1GNBYBzoysjh8lgqZFsfjpMpUdbCtiF+gk0OLjByEWPLAtSAkFesy4IMUh3EWsUwJ0FEo+upLV
YcCW8z4kMJeUh7zBae9Q06XtxfLEcO32IAE0ybQNniWBaOSBEDsbFtnkJsaDkQ8tsN6e9+uvGHOT
2H0vTUOmpyt27IO1jitqv/VFyf9rWcSBcbf4StwZlvF48shLsAYn5Czt4ZR9s/wWlp5cHspFAlt1
W8q2DSZl/8rp3YArTXIGTlDWsCHmHONZtnG1pbOUamqowwxnrjQEZXM4e30a3L6qykTrEgW1XZbg
q5PcFAIRne7PerWKjJ7KyA9ISWyuoln8TNK570pX6uqNormZ3rg0lENSn6jDeBLxlXlYZfbADhkg
BWRovvxluSQbE9Vcn87pcj+82a5kGT3OdY8M7JvVQD2X/D3IUReLDGFFWLMxfngp0bRcYHyZDaot
L5LVNFSdBgWq1DC3blyq3zlKzfKhaU91qYolqq8pWNJd1asSovBegabdanXz+Efv4YynykzDgsm6
E3+htZPfyoS4fghaGeDgm344anVfY1aSpNjynlzfMbBxzgxUF88dUxJB2WWqmNSPqW1eXxzT2UMB
+uSy+rxibQKL9TdpzlcVshZNPO8JmXQqepi5n8DN6Qff1jNvE8rkg3SZilgbr0OO/5+LJFGkrgaP
LmiG9Vi0VTk/OfBXXp7ZV9Xdgrm/WJ5YtOVQZlLlR8GeFJiDMI248wNiinrH0CegEsMkkajCmbLk
qeWWk9Mfg+ImXLzWHdP2VUimiZBsdLAhuAJDQbC2QJR6VtD40sZ+u+AKC5vYE4G5s4ejBahr3a1L
UAhM0xWdcxc/PIPiEVP0uNqhYiNcR5bvXwPFjnAJs5Xp1I4vP1B9ypBKewft06FVkHKrgcv5apDg
JOLDt10/7+PGE/gMVRGRIsg0qza/j2RYhlMOcn/SVFOlNuEX0/BMhuA4ZcblCcGRHOTqfl22I6HB
rb1I+4oYGTYIthSdsxq4FiLC+jNx1pCs8foGGQOWcrQ2BTh5xGdCPhYQweIHNRIuzvfgsWA5Vmj1
PhxXGm8fCz337+3pcNlJCZYPHDoOXCybQp+uHx/eioFFgamo/kRJRlDNLVp9s2q2cNcRwQGLPuXN
DWe3YUhg8QDlDNUHHLGe9Mn+xbKIRqQ8/B6iqud04gVbG7WAQBRjFgUk5fH4MdDLb+4xHabI++1s
CigW8oa+YwQGlcr5wZnzEJwBY14E+zL1tp/Qa6cL8UbBwYPgArEfeO4ACrwNCGHeGiwr4fAUChVz
6wW9CpHVMjlGzRT8ftqzDfvZFw3EcjKLY/+T2fD5QAtA2ylp7UiKlPOhbyYnNDTpb1W2CUuojXv2
LEWMsAtmxd8TheImOedLbmHTPCHWdRaHV04c99nUcacbF59D1IO6Z7F/uONxpQZI5hd+h3qnjNZ0
iuZylcCIkHDxTH8gmOwD3J9pJt85a6Sax1CTfQ7Ix+e9nPIamBpPRWJoQ5HixHK4QS2FSbA2bs1w
p4rNbIEuvV9vBaxB2hS/anlbtnIAVCh3J/VwcqWG8tYG1XEzV6K8kv47/acY5Wx24JDfLgr1QfhE
ug0gOrIUxVAp8+0Qe8YPpUzadto10wxm56b1qdrpR6jmSF7JCR4w8/ZgaiZuyN94qcmdRFoI4lrO
TbOREymiplqU8UMjcYxvpZgDtxpH7ibJeHoufAxNHy89BQp7m5034oLN/6ZzqgkTU1E/AW5FDN5s
1Ngo++w0zVyMLM6ArVG8sQSJBq873ucsYE+D8NofKJqA+te6aNIwYfzQIOOZhTU2JLnJcHujk0f/
Gyzgyj1LAL5g3kF2cmjqc8btz22QkypS/C1SiT/7OA46ban6OyM1+L3GymIiEeeKGsLfn7kIMC7p
JdOP/QVBHUaprN+b39S1+V3ZB8+00YLIRtfobzBjQOS1XvQCFmzILZ9JVNWIg6bMdvKanTrl4tfu
SgG9/OswpPt3HVC4BXk2gDCw6q/5SVz3Bl9exzhkb9R2jN/4YQvHnY2CZDUIPbLJet86vVbGsN2b
8yPJRZyNcP3C3XJP2iAEurJP56s7jWKoLRGRs6X/zUsh9X+CzrLYgaZXAiQ57wjdAjlTqRvOzK1p
dic7tsdqh4tapZ5FEGh44ljZLISLWtwicNZVhTN/Knt3CAkWrP1fxFfkSXRad7z88TLWk7Q86YvP
0D9WJBGAeBrYeAjcYH7Ayz39Q8YfhypE1y+6E7oz6h3mnhTS1/m/h2ARPHk8PBbGcvK6T7/AB8eP
zPJFqdPtbw0kHuS7AL/Q1vKdb/K5h9dwoczXb/XXpOLtkkX5lRTIlBPESzsxdIGP1v2Fft/QuSj3
HOmrH20WKvjXJaNcxFpwjrz4JaaLMAIOgKJLtvzw0J9F8dA+VjN+nelKFFjMb7GgM9ZFxVjX341w
F8dw2CsNm7U2sY1vjamwCEDfDggsMreqh5ZpvZgJF+OFqep0cODzN0WJfpdZwhiEmXEMbPewkd6U
/ejO7rF1fgNie0zHcNRabDm02s0PBpZyAsevrRpVQI7GSkBETW1Q6yKKx3ODDBKhnQaKrJ0Cy+dB
hBPD0vBIGrUp8eLNvGCAlpFl3iUcZ9I6g8gDyhgHIGXJ35IPUWMPs6xLIXKCbhy8Sd4rkFJqEbDe
3aWaMGbylqFl7u4V2n5BDWKmAuxfAiDFpK2X6wN+eFVUYS7ylviInF2IOMnxeDn5dwVm3CnF/9kp
pue047J4qMS3XLOL89fbyYtKPnMuUa2fJF9IoJSOfk3KflOLbwc059x8SsnOkK6jCTtbBPANCdct
Al9S2Gn+0GY/iYPUXIRz0z7fzRJgQsxZml800im7Zbl9ogMHShRkkEL/J5peTm62Z3RGCDfuEK7Y
+nxo0cEtItX8ey7tm0GqOFsDnJHdIEA0ZIqwa64EF/Q+QlJOFlajVDE3/NSzduGc95q7387svFmG
wcWqvCjwdf1GVauFq3ywQNvmXGbLIKFUNWAADTg/wZqeJsM67LtiLPkAHyoDdhnwZooVR4Sbz8Vf
69Ovk6Et1w/R2CWswtJ9CsxMSQSgQy+Jt1wmucEBB7v3PuSRhk82f7sGLuZ8F0RJ9twHuTN4WCO2
k9HyEte2OpLgO9neR6/+S+3/PH2rCKOC1QLDMDEgluGHA0y1gusqjIcCk0/NOF3rB4OwxYPtI8QO
03GejdZsPCqKRmKmQzeBPDAadRxcjGGUeOOpE6mlIYPBFNIxEoYsG2FoA0e7LedlMrnZxQ/XUosm
NhOlaZABMqB7+a9W1GLpQQUuA1GjOuWY0yNxofT15SxROthPybyNtNAlKw7fL7PN4ccFwmKFl2yf
P8xVL2xm4TGjBpOlDZZOMJgVFQnK50ojARekqslitJehk8lCvAb82m8xE6Oi3StZbTYNxlBROCgk
kPgmX1xTiL3OibOql8UHGETrkfqrZL1KVYazdv6Nad0n+/51z39a3N0tIOO/dlfmizjafPUS9Clr
QN2KciJbA3Z/gQ6CuEfx+S38htu33phSJPsjwRvMTpNgRGjxlRqyx0EAyX+mc78f68KtcG80P6DF
ChscvwYDXH5Ue9/2PbeewzFZdCkLIXi1yiIe46reBv8wI1W3QfjjqFVg67ZMnzb3HKCDdCVwOVC0
nPoGQTXL9dwSXah0BqlieGuhCXHKlWRlXq8Hq3kHg+1N4U6YFlDg63nntCKWfpkoj0YWbPZJbPOl
Et/4B29UJAAHdnO8Eo6czLpVZ6QA49NaW7sHRJuyvbhncTBhnCI8sb1FuZuNmrj0Yw5r77x9pSRp
8oyyXABkDRV50OIjU0E7B9XYfnT0BaVrclPRrxIdfTZNdMlua9OORhGPpf5tehI0ZKxYlX2pNyFt
N+Z15L1B6sH7izD99PP1trQCRvRKKV1QSE2MYEKRs/DTd4qrmgS4QxcB2+B94zwgjzlhEW4XK3+A
opf6lJ8DDugqSqyclfOb8CnRTpksxHalhKO9z0G6gJ0b2vZa8zkqclP6TQUCEgS7nwaLy/4lAvZ0
DFaBPIh/qNF6/ZPkVmydf9V1PeqJdQT4Z5DoDMtduJZYauCK56ilW9/E3IXngaKMGC5p0nQJ4iqV
Kdke1Nab00AklnqkJXToWn9uoapB5Ig9DyV7BBttpzArfbNdle9tF5Zx6K7lD6H2veIJVZ0Ndjjh
PLSp18YjP2yrI4tKvpMAVlEuckSfVKZejT5YInyQYYGxRx3w7FxhEYdXOB4nr3awYIsrUb3wn3PQ
t5ZYc+1GciUTIZ76TNbG/Dg7kNIGe3APvjC5LrAmY3DJ37ywMfNBR0iNdY+nuta+fcHixKNmCvZe
iiTyN7kJ7ctDL2EZjJXjob0Ro8YFJh3rGz6LRWM19dmaW7KJXjhJ0zGPpr9IdbL6c5AWRz8sSSt0
wyElZSkYasmqguFXMgSRjnedqviqKdEjZt6W/HHTv8ni+iaAtfZtkFDWHko9zpQutw3271AiiKjn
CqpHGxNwWzhtHbxqvMWA6fhWI9BGR7mrZerIlqOF4QEvlNc9dmgTikKmu6twH2Uau/Rnc29Yxrxr
QPzVF3+aw4jD8rce9TuydXiOyyFwbgOcwceNO77homUkH1B89o2EAZJAlnhqawaAUOcSY2o2dGbV
54pafQYxvBGVfNMV+EXA+7Dv2a/OBBUdzc/6ZZfFBXSgXwXO6K9GleDKtxG+E1tEDo8dZkmHLM/K
omvBfeuUadpiZZCoZgB//LxukgUPMTdrfYOlOLMaRu2UKHBs1q9mRnqt92JmRQJnh7YyZ0xL6fHe
PEaI8S5MneljSJ7hTs+94UDezlLWSwkwpb7KMoUd+CT3cAqNAfQDj8F0do+oYyHWQSfjwKeAtYxF
bcxW5APWz37ujKT7P7G5BTC3RUH5IFtPnZx96VEv+0TPCUTatAdOvro1eAr5YlXjqfwyLhafNH3I
5LkOlZ9+xFoNH9AbsBJr7FJLHp3G3wLJ60B7hKQWym8Ir6NzmzD32gObMVhpTQY/U2ImFppsxdFh
r3Hj8dUtOniwibF4mh8N6ZC8bljWu+Vzi5P8eu+RpAMeL+wqPyMRBYU8glEqOXJ9eLqvH4BFu63n
5dqDHRW8+ABV4OvwCwnH/FAnLiw/SIsaqGTx+NfF9ReK8TU9y3wyXMDPmkPnziDH61sP2tiHUckk
si5gqvzXX7pzmcuKAl1zxyrnH9cuOnbNIzTi0pDwf7gpd9gTXLMJZ09ul79aQAo4va0iymn4qKJg
7AR9dHp24CYc14aocVWKu8DrkNJF1IHSyBoYyR1y6vYh7MWBARKy/+vwZ59SnW33dJCwg5wszlqj
vug/po3P4qhkwRuhEkDFX0nZrKg1ClErkUND3U9O4wVV8QGcjYpPh23pjPz5/lPeAisqHUqTJ0zM
mrYN/kkh4tn0uc6oTvvPmflrkTZY8bUFhA2Lk0aFu8RV5tlroHmeFCrUb92rl3RdpLdGKY8uBGI8
+LTfdyd9E2WPCPmU4sKI2R4txK/WQn19HVdbrLYPgEDS2PJsz7egKdjgCZEQdL7Ej4KoNoxP9Rqk
HtvSdi/lo7RDrShNeCtGKmVjDKSYbN6+Cdj00x5D1mFam6tl0P/SOzehgFdbwPXGd0EaMHoUeu3s
XGzUgi3WEtqDLio8WRzZ5E9BFgKQCTsv+th4PFtjbWAPlgINZc2jYKMog54PMSKRUyPV6iMNQHhO
gIth8AGiQnoENjKe/YsqRR33m3yXBlsQf5LeCwWwCEBTWvmzXqtTqDmhBYL90b0Sjp1CvFVjSmSi
r+bau0ikhHNJtaEIpG00u2EqpTKQX1K09yBYhDPmC7o3IdyKoSP6T9nwpXIA/pgQumAUtZAyOE+1
BTyXSBnJ1fj+ShfIebX8OH/9BFeMzKgNOHO7LDC7mDwD83QBvJTdd5QsiiLEEjo/9RU+F8iTQADe
MdskUoy+ELuKPM2r40J/HieQROYjcMJ8AZz0/EKY7qlFnSpzMfBWPBESQ4Cq2y0p7vNkeTj7ATnf
O9KcTjNB7f1OjHIfsRnjZ/cHpKcUavrqIcWeMFcAfxos7ko2L89mj87vo1gAcSeaPWxzlakOi7Qq
ikzRiXgTElzS6IDWtZ3N9rZo1DoCUJG3u/rbe79NsudbzZFSoJlE0lAjHmwCTDjL1JhuQRdwuH5X
XmrivUewgF3L9i3m2jv28x6v50/BF2zT6/5IrZGuRmEGb1jy2c8W6N7NXKC6EHOZhNowp0rJEPT3
hNDN/YjxEG6bYgQtk58+xOUkLfj3jKJgfMpg+HA5HZY38JHDKvN3+MLSRxmGw+qgS/k7+1gbdzgP
NHkKX/ezaJ/0qcPZ6Sf0CC1piRU5NPXRDp1PFPnVHSCrePkNwxd8eUPpBL9JVAttdLQLP01vxyTX
2ENkw9QS3UbQB2qVE1Wy5PbYqb59GvBwdPg9tb3bJp/QMO9ZlY9V1t9YGWS0TXCA1THVLMkWgbLQ
3+jxyWdIu6RT2GrekEgXXdxopwoGNxAE6nmUErUAxMW0kExW6PMzaYIYRII2wyBNrc5TwfswC963
mn7i0H0R42KYa+FHU9f2wimbXG43rn9h7ae45DVu/ow7WQ2rDyFFLJqPzXnGJMJE1Ao8f6a6AKyR
9+CwIBoVCMUx74xfjpzK8n3/bNAaUglMt8l3IKMHhlKDN5KP/+tqFaUykFF6GopgBbqJeOWxmpAc
FEpLClqGgIUj0BYbQtnYWgHgFqlPRF0Nu3tZyY9l60krk8lOlpltCYt4MFVAQAlOurymZnUKaJ3L
PVJukJUNvwfezDQ//YHRTEVRaipLsAxyMS5/ai10ZGkFoYz1riRwLATbKrw6EcxVf80oixDAxhzU
eoyjuBUVjTSCFkrLOPYbgrDL5iEgmwyxawgB5ERLABd8d9fu5oLvKTNo9qtm47k73uOilEiMdrs8
TVz/351pLqJNJXApBan3CpUEDDB0nSSE4FMTJL7+wu8MzjTwSiGyTZQcOaA3zHtBxtG7n5H3w0xd
QGJtjZElqhoAuUzG2BruKw1sD+x4l0j4sRz6/0SXP+KRuNxRmM2QJpj0+sdpZU7FS9mRVx8NB0SO
EhrC0Qb0f1UaKE9zenHOFjuwf77qaG9Iyj9mgao8Pp9VZh1gUTXfGRWtj0Jb+cfn2gojnNIc1hhz
5wnm1DpN7rW+ToGgc/9QlgVKbAM9EUsixoeb7EqyJfwcVjrSndLQjpigsIHsU+MfhzSkPjsTTxXk
Zbqw2k5io/SLhW6BxGBUrMa1/ty3+3eP8U55j2gqkIKjoO5CAXD8bLdv0lubJxE7ArbvNRvultk8
98BVrO4GdoYXtD3Q6UQjZq/tL/LSE4D9SSofN+DoUwqbD6ONnDANJcdjcedPpYGjLSQy9kaqgOBs
aqvaBzAoVtQvzaJvVn0TfS8/1eXpzN9kAMovt87AodgSuKpDg+5FcPaMDTnVbISuKJzrqERd6H/B
6qrxDFHn6+529uX42NwjydKbaUM62kSwvgHuz8xnj/8+SvNO4bMrbzpwPJIuL/EAVTrOVRslDrVB
Jx5cPNMm0tTK/vUb5m7pgWpBJ1J2/7TqcI7G4KZzw+XiQRbQpZydy/B8n06LvPgBCcVwI9UN5YTe
+Zj9ip5SffTF3o20X00uVi7Jj4ry9myETzM6ByMNtrfEDX4UqxVdP0EkDZ8fUo/9UdOl1LnOTBER
TERLnUjOKm4Sdbmb0slByW+CLYwKhqcFozWWoUnJO9aQXLHruqAXnSGJbsJ25x3joGMC0w02eA0f
F9Fye4LX/dDEKva3MDGpKnOGoyLiyn7jGQ2nMzZRnrvHMP6Vb4oFLl7KYoyZN0tGywe5xsAdI+7K
ScIlnsOycv2Gl9I91cWssEOLbl5FcfxG6mCiVk+BRjjVVoT8hLzT8F676Mpw9Fziq0oGstO2IfDG
hok1W8Ljx032Nw2Ls04FkCCrZFfjEG1ONIfu2hPFGuJ8OX9J8sRW4Po2R/qFy7EbylENeuklXvLZ
hz7ouiqfle9mIAyTZ62dBTqkrhAfrGIBmRQJeBZ3HryRd0hAVaJUzq8xpKCvLYQ2LYci4qQUk8zK
mLUItKVzlkLbuzJrpp7kBV0uOCHk90ogH/8RaWLQrhFdZlb31/6MZKCfD4e6T1ftkXRwEdxnTMP4
jWTx4KBuUG9GDtLfz0ORToRMMjF8EO6EDbptllaRyWbV1PXakDA1UIPWGdBlL0tGbySpR/MNCmU1
y9HGuQfDP4NEc1P3PV4F4S3LgYeJPAEiuOZwgrp35Ks5TBXb2nJubbmYRzDvLA+gAugLL19suF71
hGp1xRBLTa7S7VA8ZRhL8UeFziXcpYKbuNgwbnM/51GhJHTLE857+RDw6DlhOtTVxAP5AMkWpPWc
CPb0Muk1HZfpRxYhDiL853a1VEfbMYGiV4d2YrmecFIruPj5toR8EnQXy5hjcXPIY8miZwfNBznx
47V2vc/FUf9NDs5pQeDsedYEca/m/3kpIUqqZpxT9YF0PHNa3FR70JI/FhbYZTNLSKSeQdcjxL+7
9iGT6SKVtQAP12sRwP97BeqEWoIiYmL1H9Yd/KgyqDDSuBl2T36U05AsI3HE2VEuPvToOkAs/cGG
5SdmT9vr6LS0TprEydOy+V8lw8/hNdQg7TETpR/xjtWOybBqsJg2dFzQIwlKtBVqZ8PFV6diV8wf
PxRiKLfNP5l3GDc28gvRNII3AadYg1+dXy3eTwAI+MnmOO7Gk0OeZsI9gp6qR5bsGpusLtnqAlZH
5hWPVbx0zK6s/2rn7vye/1xeglF+gneDog3eLRaHsOVXKLGT4WWeEEFhYxRVPt/eexlps4UEX48b
xryN/MMohPjYPVcNBq6JtFNETuzolw06CtY+okfjoY7LMQWYH40gVkj2vJzHX6PFM0CpFTIxI1Kv
uKQjoJIkQ/I+JBwda6uU8HT4LG5e/4bVp+++mYq6P8ZSY2PdIYwptPcgGKT1bzJVTaP6waoBQIQS
nHuZndSlSWYd8X0y3ellww4tvt89WvpEbY8KZFtkU+EGRDFvQuBueSDB5oXHi1x/zMggZNQ1heW/
suHEwZDJ6MTkvMx/94ON9Eox79beCzkW++Pup0Hl2kk7D4D6qcBeFrTOYzT2CHgdkJ8z/QrkheSM
T8Zs0foAj8MWR2ZCWilDtp+KAbsWKLUL4mEga+Zcq6C0DdZM/68RWeuuAxcnJa7quEJ7eVHvn6Jl
RmA3VqE2gcH0bhP0HPHHXPD8S1iHxJhXevh6cBbGcqxBr6qrhiEaAtAku1UtaocpXnV8cDM9Wwwv
SmAAEVqoSL3jJ6urL5K10pznFZ3SgUyoMFRB1mRJ2AcXnxHVknmWq3LiM/UHoQFFcOve9oq8qRxQ
8yc0XODvf1v7z0HdK17toCsTYOc/xNntdUrPQ6cmzh0rpBnUooi7Wf5dIQ8lwCpnElaG8u+jnpeR
ROSXld1tWVNxfOi+CSHK/xWCi/azKpjAnqBjdMeIeHlq9jPTv2C/q5IrCkHL1bbmugMKgod9xzj4
xoEY4WU3xLVKMtRqN1S/nl28/4n23vkQZ6vNy/kcDtlYQPssSLnaLsGUMQpWv1cvzH5cxY8svqcd
Ei/UxpGFoJRc9gzioHdHD2c8GuS1xgIsoSuubVL9FKE5CM5LlpeHW5e+qF5P4w64TssbZAkEiITv
8YI11kTobxUFd3SgNMoBwl2tsedNu1lvu+1jkvHwKQVimYs0PWV8fD+wONK6fGywfkwAtSEUTZFm
a4FkwEG77SodgEhk9xGIgSTYfKncq2wCswMgxyYCvqRHHONU26oIaqw9IgVdsEu5wCqfrDiQnV0t
bFwyVtloei/LgibXT1TJq51O2I7yBcRJiZlsmqGyOBUz5D4InlgBg5c/tohR48FzDXKqPuc09Zmm
KfN8yGmBYtxuAGzhaTnRND7qZcPY54akkKZ6LZgQqU4KiPjISIs+UFjQ9hnD2laA0b+Uvox4wJTx
AdSOrZM+gZGzhM7Jj6mo94zcLPXoE4d0TiigGbbQo2Wbi5sZc6SDM5F3cHT372BJ6bHgvTjGhM6b
EW4PYBwMFauPKtUOT9F9o9N2elSsF+GigBvq2sjA+3bSxbb9nT+wForZfDYu7gPgpRc3rztJT4Ne
J5tO67rda4O3nmduWYmoFokfrDRG1u3k2fRq4NWTwgWyLgYzAEZV+W2C8H/S67q8b841N/aU+cJD
LCRdeC/T11c+rylxjuDRuKdiIMkd4cB47nlIEusz319cIu1qmcxbaNPj/XB67z17E4OVBa6gA2KK
vb5o7vw4Tn6Sr4qhlNpBqcJxW8/TkPqH6w+/IpG6cyf+qLYMzInmUkS8PiYQNZgULn2+c3L/bHCb
It3Tz+/Tc6pAqYhPEPQhuN01rt+Q7KR5o8AMa0Ts3xPGZLVVdToutYXr0HWQ/CRf/H3GJkHH4du8
ABenRYWfHpgCexhozJH7rOc88eL27ZJU2mYjUze3PVhi5PHXYNIIbaWwCkQcxCYwvmhZpOLGM38p
I2xqahCDKpPiSmUlC9LwrI54aZCYUGATGaHHu2Rl3uVBR9HiX5BmBAJT0xVp7u4FPowgF6LPdQ0a
i6cNO0CujjYY0X3tpKqujzYfeShkWiV6qZlvlhSWCuxlcFCxVmaS0PXi1OaYh3+TI+JbMCQUetj4
+mws+L7rsURn1NVM8I2QbnvkD/0FYJ7hlizfWGozyKwYMqh/n5fceBKiT80QcVUGnSrACKDTw1S4
2Cc/iZfgZoC92ldtLBZ/WBmzROSyZYSzW6jpIk9e64GnPR4CZTY4ZMl2MMDSFZttzRbcPZwpRGcQ
MN1dGPZ6AQmW0oEN8KwhmwQ9FaKttPaI8UvBTnB6LOLGe5zFw5rxZQl9PD68lBJGO6gglHRIrqnH
xmYN9kerEZ2IkCUOLPydT40iJaZSt2jBJl291tVWignoKG0wFUO511u41HEnA8AV3vwNWpnoQe6B
+m5wCYAU2r7iD4dPDt1oAePlK1fyUyU2UpsMWv5DpQ1eNsFREPPlajXsh5AhJFGyT0j+iIKdg0E7
9D8ediY7/Bt2G833M+2JTbtk40Uz/KRBG1EetkJq3naW93lweKzZ1NQCyQdkc6Pxez4v+RIBDBeX
IjAYB6Y5jgcx7EgAz/JrB8FG9K4e1sQnbY+bWQZu6oSj17BKDp1jXO2FsvcBdwDxxrWJJDTnq5RJ
VMrvC1XkQFFm7IaTDRWfhHKuo19NEeO4GQ2cVRA+MBStGbYmOgirRJIdRP66O0ZlU9YpqsRSmEqY
M/toJy3H0l67fZC613PkSpPw23p2XWNLr22duJuIkO94OwIKbfpurg08TdvHFISGYvqDJ1xQu4WU
tVg4GQoRcQXY7rH1kxkn+XZfrHVlyd9zO8uxCWEvw0x9yu0Z0pSuTLU3UfTpHjcvv/hgG8ywS22S
OHDzR9ReiLVqBo27aAZYk8YlMwAM6EY3dcEH92gylJ8qC5cTirjTc+rWtPbPxeE6+kMbXEGBMVCj
4GVmHNgjZW2oV8Vm4t+y3pfDydELaW2Xmx71CpLu4PLxyF3nFyg4/qxhmEwOOYlOginVEaeyVOXV
bdzK991Sq+Rn34uvXPdMOhtZDFP0pbF/OvEhvDpRhr6hAd9PcnmcCARfnZfGCUEmYCDRDwDBifDB
zsIN43YbDDu7ReVwzaLosrIxt0MeXfBSuPCEzMvxEMLThqiSRt/IsD3ZHAXDiJOjjIpsWG90/N9C
rd4xCMy5XyOy4GlgIayaYBpYKu/mnC8XWIx5vPl/mBDNf4rrntOVyps9LL7OsQ41j3yb4wSh9WSA
M3gIOPjwYDXQOUYYal5qAzQUfpNdAAzdaiKm4jK7isJDX+AETpkSGU/rx5LqQfl9gLaEZwNcRpVH
IsHdqBJl4bCw2++EfwLKuzMJyW6D5xKbDnlA4uGXQoOeeVbA0dNKqdToN8EA48VlKc4syuO9rz+g
JmbI/lH9+BrQrrqk9KMmlxxykcRX5c6SbIbDb7rLdJA9tOVOqMOV0dof/HaI5I43jba29mmEzjKq
JguR4+C3nNXbh6WktynlvJuMZcoNVb+SBUKGRQVmKYrICOhU7VU2pN0hWstkfPbyZmuwmT4C0nJ9
17jp8QK3ClTnNZ0laAeWbt+dvlx2mAlt1+knI7Du3+vgHRPpz4qCvxUFBnurlIypmQrCDDK35xOk
24tCBnXYoZkHW1J1eNXLqlekQvuKUM3O7SdHwQeY4HnSrQnTpTSaQRcjghLt7RfUaSP+be3iogbF
hL7++UJvYdvtNu3ehb80+PsYSNCXvz8VF8TTh92qaOtKG874xrvWRRHS0R064wsfSyMfsGFpdSl1
Mx/SuLFUrE4dLtS6tsLg+g8KNjqkLDvce/XzCpuI/8dO3lBqw7PVbSBGhTBTJJA83XxniEl8T/HJ
GYwMFrdGMfLEsqtZjebW0r6xcIwYeWAI1pPHc/Sih2FMvG04XtbuUZ7aD3OJudvDq4iJp/ja9GU2
0xUUoIUSlic8xeVv/nd/IIWdNVP2dyxe65en6DeNA8k+vNg3c0sXjc1AHXucrKeaNK1F5cXiOG5X
jcvrrTvXTUJ2V3TQnZ0eDG6T0N0nw1++MHisaeKVWpQStkRRvNoqMIRfPkyxUehpowfrQnvaM2wv
hWt/Z0CXvnhQTe8V1iRHj4uKCs/awfWU6EFnSCwDR4qC3h8J8Ev2MJuK6vmSZRtZdpVU82S7iLyt
6gduqQvFsRe0AfV8trrF3D7AYZmeDK4VgdI6J89ZdYifbXrW2NsoQOJDByJN0PUN0V6RJj+qXcic
Ik8OrxnefpPNUmvpCChOlKCf7/ZdovcXd2CKh4FG0NpIG1SYRfY/QgnMWA3p7PIcJBbcSkzs4Fp4
iePOnkVdDv6b28GiNJ+/q7Z2nEzGp6KYsWpKHfHwP70e33iArKQhCErvvGmHT9aR4pBW9/b56MRg
8VegekFCO8EGoj4EHkNp+KSZNSGC2Ew2uHTCtVbaiKD7u3kBAwHXdAxSb88A5AMBAYEdEuNc+2Q4
5i+r9gv0hG21pA42u8lQaVMR4rwzf0/WOsoyiSZbOT1DZh0+iDk7znF6ry1eJcRCgRiLCwXf3YGW
dIu9bfXVMp/4zeh3Yp3JIu4KrfQnEEzSyrWltam7zm6ME8h8ZTt90Pb4mm4YD2HOcujsSa63iJQ5
Kf2VSEQIZMMjZPEFnPizdQsA5mU2qpLjNoj98g/NYYWJfjpBWPqXBhRCj9R5gqxMkyOcxvtN2bhk
EBZslMVnqLOuxajeky+6EHpSbIiI4xUdORPHMyJuS3J5SQ30KAEzeAKsFoLXJdDcqDtuVIuB/oaA
EDKRTokGIBbLEq4udPhWtqSYC6sRr6QlP9QagKzyDXLSY4mhWVy3w9ki0sqMGQ3l9PlcjM1cIoZd
uKolzIq+8f/Quu9GHVfEVXcLnCw44PjqAzOMSOGF37zfInv/ZhRcLoZJsKCk/dT7vf8FGXK3bsju
fi2TEwgF0uLkNScU/wlxf98V1AQEQSqQJ/hK9VgnW/jcnu/eklo5AmA3FZo65B2l9znyN/+/3WWR
5fu/EwLdy6eoAxbhx/54X4sFvcYXkFmX1SWD8AUeOxfi4AnBtcfoOOYb54uK74uHbCdSUaUoolhk
NluwWBPTK5fRdLZbSItXQYR/H+OElWWUkzbHRiODY7b7aw/nG6W8j7Fy926oje5/080LHEqwSp1K
sy3TLLevgaVrXH9hzf5ezvOFJkjZSoaZulGeI6PceI8DRUvHS3niehE/iemgK2wAXBuFZG+QMOgv
Ve/YaGpfsRfebr4k8plioN3sKAXxZZTC4XyYQYveWJ+rWzvH449XSFJQJ0w3l1YKjW8x5gpV9aV3
xbR9jSTO7gtEgp+eckxGema2Z+Yn2RtG01XymKPzrF2S4HZedRyWxhzKguKd6ptiGZ2uVx3wDESF
WFTBElLGplmNjg3otNkKKcTnQZqWoKDkS3rQanFMNVPV5ywTeaF8d0etmvq5TP/v0xZWmQZOj6wr
EEuVQVLN/RECcl3/jzcUOyR43JGTPhNTSm6XKwL1+wxIZfEplu9OJygEOevebqQszjNrmdOwfYwQ
FkWz8F44veC8c94XG07PnhPcWQMj2RWPnGmrjif/n5K+AQfsDGyKfpGjQ6o0cki+JuUQ4vQmdPex
utAnrFJiqQSA3nklTdxCZnyrMqYAug5BE6lOD5ReP1JiaB7gvngRK0hT+7CZYhyxYVExCOan4QTl
lyeogGnNmTlsheIiXznhLr/AI6hn4UJVFPbqjXmKHqvJ5nPwckPTYUQL9AhUG4y8LQtknP4FzTrf
c/MUDTa8HK9LIAO29sRr53EYPRgOSC3axSNjDcAYa6a22wjrVmxpAqO03NbKbZgpDmcwI9aWnQPg
BExKLiXm7dh0eBBp07vc1gAekvAzfmZUdwVNlHDbltX6Nwv0/kn+SnxZINZLt56JrlT5zQR9/joe
vn0w3uzU9hnKYBX/LXMEbnpLuIru8VRzbynVJJrD82i4lH6K5c1GPeeYK8ppd29dH8csX2Zn0vPn
fGykHGWN6mn4JCRHWwO4unlRzZNaLoBKcwDYrlBUeKxJvX/sulrts/wdo/InOVsEqKDxOlgTMrto
H22d9Zy/CB9zCOwwRYKMT+IMzujDptf0i3mIDOnlgAL5PB3m5oDZFFQdFVoQ+CAyq6ooTgWbCEvS
f83i1IZafocakzKjolukdbmWB9k+seFszQAyyMK/AatFLMd04UNrMFe6CI/pDGt4ElZsrCNlAvRK
4tf40YyS6v9KHIFi78PrBwJU1O8gqrI5vV7QsJ9CVBXQ47wINsFYhUkPABvn/RD+ElUeCboTjsiO
yZ0D1iCO5RIyYQuLtbHWZmgbsgmajk7tK6oaqSILp/iTU55JpxkJbv61EZh5V+zFc8GvllJ2R+92
g5gEe4C8UJZX5uX7Yc4g7/JH7PrCyRBMrlV3pzfVzKtWwVapGtpiUA8DMjr+Ks6uKQw5iRj0LN6C
E1a0ySLRs6QmWrhTZSm4JLWfuINdDNSoDx0oxr94DD/+AK05d8Uc9tvJEbthmSczeqoJxuWDxjEn
kvyEKlgrRSQl0ni+EqtRnKjwHwg0ZFjhMGSIdEFYhGrgpe+Cpds9D7yZSDjQ+8p3m1EgUz6WIj40
zIp3EQ6EZ2y4AJfq3QoFfOxc0gIEJxHlLdcaYk02AnvJcGbUB9x+TGxVcNaRf98tlE2cSsVpLXsR
rlkjTLCNHcbwN2QJ0kcUhWE++MchZqWTrUJStxOPrG1GHaYUrPF/bZLWrufG9JMoaHLDgm3WRybW
KgETIfKg427pGhK6duwN1bAD09gXxOEP+BizMMpSu5K7hZ27t/4vAKAiwmHQ/SrzqY8C3gKcudlJ
uYxAv0Zq26/mRBZGqyIpz8E0kShfemjQtnF/ONZ6NrXGArH8RPfwIx1+6Y6T1LVypwBLpEqFeTO8
EtmzM85mICuKxZLTankdcE6PZyD0kOTtvxSIKk2yu7cpcvkE8ka4Lzb3/XYNfs0gdJOQ+s7J7XPl
fnCCifpqotW+1gQqCa4lL3wpkUZZKwwhoDpXIBJDtDIyBIXO+2jb5cKW5NpaJtWXf410xIXhWIyB
uiAHEIEGg4rs/cJmQsM7/QFFLuzn3x/Ds5ZeKSAL8Wx8+MIfWC4vh3MKWuWi0LnEpmivwTm/hmru
HDqaAQuZc3EGFzs34qZ+fGmTFlkrrIII+bjq+g3bHoZAYUUXJgfh7d2cbMW8oKAsVKNrTdZ1h2Kq
MGDliMOu9YrQ9bxTmPz/iRRZ60wiqd00cjWULlcWxj738HaMxx5fojZLXgOM9O5gmWM7p0KjAmqS
d6lDvIgKBvbza+3JKdn2JwlaPo7rJoRmqiaZ37vJShATZTeH3yIMfaJzlenehEY+x/88SSdrbh6C
YajD/KkpOoGWhKOZLIXCD5NEC0OH7AAEggawAiSnXoCQRADj3kvlrWBIWLmIYsC2GaLyqM7iJTtD
Wh7++9lSqQ+ZpHl38BzDz97lWmg/WP+RMxznkF36qZX9fgeR/ibjkAUdU9GJVfDttO/GC9iXY/xU
aEE1xQO54RAZMO/M88EuD49d8AqN/hTEKGrj00qmhaY3Ztl1nVd6F/UTloN1klOubPMT32GuWe8T
BgaYjh/BZkftgjwoeSluGv1MQD9lYoso83QI/LGbNzDbxby7MJTtmD0ZeAE0VOjJfIAN0f+w8xAf
eYO9b0qGa9BPxeediyPjmCZx9R2ueI407gi8iB1hH9Z0RIJfYnzrDBfvgNO74X9hC4gulnGQgQOb
G2f24aaRiMVcBoPWQFERR5v/1DLspm992IjlItV14GuA2TSOZujNEJpLirHD07jp/FqTA7/Jo1gm
FPspwY4bbbQEljYFyMbt5fe+/2DgLSquJ/Dj7W10YC6CTRuSkcop0WVvtzQnWyUuFA2V6CYQ7lXV
ZaM9l5szH0vkxENQ5G+q5hcMj519/jOWZFZFK123pedbywyMgXUzVy0SmEG5Xj3bqgscrMFvEz37
1+1W0zCExlX20vjJTnVyf3RYWPGiY6uWQcFtirN4ed6ZnMJuIhiIIkWtPaalf03vXEhQy3W3Kn8R
/lfZhMBeIWyLPvSylAxhU/mOnVt0U8fox2Rs/EG7orcjc3+nipSbHBdAeqYNrLGitPp7KohIjJf4
qCEl5RDzNHaxLye/JWEqtXM4xm0koS6/ELNah81WI+o2bg4zby/su+y9yAKfLE2bxmXnMBFS33ER
i4Mk+myUQ6mFHiA+P8052mRBnxztFzYdHhcgyVFLkiISsbsKY4HTRfHCCYZrV5OJ6VfSOb14hg9u
gf1wr2w4Eievgy/nJQ1bGyci8iuA9Sab4QaQDcGOfygAJK+vute4IgSQSW+rvF4YNNwXKMBiGccB
LDz5LcVh0hj0M4Z4pd+sYncyksuQ7dkviPTgRY8mI4OMspEjYJuxgYSCoQgdGeNX/fTBFcHiR8Jd
j05RGasSdtzgXrNgwfW+dgBsbc2jGIDAWBmmXr8+wPg8XH1IyiPsdtFb28mDayei4MS3nCCIB10n
P9odBOVvW6JgnDUoH1PUeCH9f68/Z02lEZb++R5QDIX/ytrs1mJulACauaf15OMP8xCNNV17yYAd
KtwBhurro0oAImytih1Of1dRSaQwNyaYirfafrPJaYT0b6rh6hhtVbNn/A3nQGhWjoQpVOEJEDOG
OCjYRf2jXfbNuxNbNhztdt30+lhu2hXQpN9b0fgxqqIePiftljAXYWu11yye1hDd7qFggYMNY9C6
2Lp6rw23mhtnCd9IQZZx6rojMxx6GYzUZwh8ui9u/uRP4CrybeTOkyTPCwWXiqiJndT2Np0L6d+V
Bwic0tmQwGOitgtvETPrOFhulty6jPoKmKvFJ93sSy97QEdbEm0ZMlDWY5ff0zSHzYYXbMG0k7Cn
js4JeszwsIUQHYF8xSwJPJr5V7jsx2iETSY10pbTxPcwjgjlz7X0Rawfxlwxm2dRGj7V6qlbBIc0
SyW4zHCdodjN26N180W+c1T/vNYJocnAX6D/KV0dq3FTmWSVRhnmHd1TEtOY2/XT4YMalIj5tupi
y093sxvsy9Tdzz0QugqOZ6P9HchiLNSdcVRL+H9qc5lcu7e04URlUGv7LtWeHjrokVaFVytVP9+V
BirWc62LJBPw24iW5PE0ErN3eMjp/fQFmlPsJupNcmWkQLeT5TAT/SYEM0HvKA5u+VdoEbF3wo8D
CzkuOUhGwho6N+rA9W70PcOmhwCTX80gjXxOOyLvITti3+mtaDh8PbwQD7LaEeA8SROrBX9/705E
Kj5/svzG5QejjSGmNnaQGIixbnkKiLFBazDT/CGUhrDc467YJ41bW/WBk6J0XX/rCTv6PFERvoZR
VJzFLq5AngpTy9IiyXFU6yTFgGi1V/a0CycreoOeKLix0Ho9or4kuPjzeSXX1Go7Z0dAe2LQ/Bu+
XyXBoqDEl2ypbIJ2LNMzQMwGiW1Jyq87RQKFOZc+yTnQQ723kCngNV5qWiVVxdFIpy8HeAstXw7T
n8sW4JvpGLtehdCMlayCsl1goZ19h+joCH6koxn5IASq99x3NETzsLJcG1eVVqHxGzRWp3L8SgNI
J5zrQRc2yohtkRFsQyyYv9LF5OmXQd77cWycgCUrbbDQbD4datHCS86cvFOPsw98AR9PEQgpoNEM
R5xYK5ggdFNURM3cm+EYYgLsSWuKl6KfGaJoOiEYEvC1RCypF+wDSo6rbFyfE7m017bnQV4xgjq3
1enUHdD3owIJ9zrFSEArQkIgqieppQhyB0R8zZWIa2QZgBYYJQF6+sE2jee8cDolNpT6DIpFWhmy
QmX6Iy0mB5DuCAaBO1k+3kTUULFXSGVRbSe3idGMcXO2m+L1hXFC4W4hbCAfrnaHsAmiCojKPcqS
yLSoO+zWgKmqTZTXphUaOp/c5nALydu6JBKoAqMgneJpwMPnnI7AvDAK4v3P9tlnZES3OX1cymt3
vmMBNuRtMEQypaUsihYk/DxkG/rNJlFvfPCcI3m2E9HUKjPAyKghQb9XrrmeHyNn+/Z+hYzbIUmf
aqwsOSIhB/chquAJWUNSLvuAU6vJpDAIiV3CHJI8Hx0zveXFUluXZeZZ4YnUzbiD/Re9xECpv+34
BkM7bX6ggRjeG+JocwrMP12pmA4QZoOTlenv4cNI5wP5FZvj9MwkwoHNdSnvaJG55OxskS4h1/hH
aJAw+6sZon8wtU4xjvTMRSPeS8fEmlgsXWTJoYTnQAr5Ck0dIsEMRzBqnFd1wjeR7gO7enMAMmzt
e57TNPWL3TPscCX0bD0hQUW77HmcsYJMB7synwmBh2D/ZQl6mGRSNqJfDgoRUGHD29whvAbtFqNb
veOoIj3twU3hHl5oknJFkI062nk63v/ydNAHq41I+eHxGMv5/uZS+JQnchtM+u1/8N4sp1P9uXIC
70fse8HwEL0eUUppqWvXbX27VYOmpQ5gss3cO1lAaCi+QkcKAvJatmsinC34Z4lMfVGC56RtpcTL
7piV6BCu0AKPSaacx6wb+HXdOwWk5T1I6EwQrQaAF1yhW88GbTUP0RrlPTjdCrprS8YbrrpEVyxd
1nQWWbt83gla6HJu5sgrlbi7klEfNwrPMRgqj10+VOB/taCbtKBV8z7uZkQvz1iYr1fPkXXf+0w9
/uFk65thAbw3gC6BufjzdFsiHmlz51BVVtaNaVj2tdecp3XyCaGjtDXv/Lkn6oCjBwLNyxn/Mde7
1CBB4Sh8fRomsCAhVNR/anltDjGAA/xi2ke8Wr6c2tGVMfaGs+x0vmkb2dGkQVvunz0UQ0njXXWg
oThkQ0htig8L5zBWGW3RPidm5qnHzBZOpzf5jH0GIXi3OJfu6EXapBRPSk6ZRiKb7qd2FVSnluYI
5F5t1hkXfQjpLFcA0LuJxPWtPHIFe1Tg8zVcGaieST9vuuMVgJpVIyP7hTvZjpQFqy1/aZMk66iP
cHKq7es3FlFy8XPj3CJt8j/fmB9WJjJSuZjmlYYcSFVFVbPhvQ67PP8b2DRQ6hrTk4IbgwDRLzi2
Y2fmozG55ag0HrYcb9mTUoROFzC9aC6XjjKIEgomxy1UrS7bmeJ8qR1KujYOeme5qg6z8MIJwT1f
pYrVmUdkchIlvMDx5MhkebuyhuPyvg5AW4sZJ27EBg2iJ9Uv6EvzhImLZtauvmhUmXkhmIbeMiBf
MwIpqI7iUhY0fSuZknCBi2uvnGVu7qKS4HdGN6cz3Yy9b4bAa0AuvTIN9sbduEqIr6/6WJ8vRvvX
/EQQ2kK6fVeSjOWTAgdEP3y0cp9RRblqAbvEpFL6lhwD1mG+vSzi84XztC/jRrCT/paUWfIiHX11
RFBpHTYpVs4k0H8FCgzj1O2W7Yb3jsIF5JIhaJkBBHyxCSvPMeBMWTyJjFF4qKr9yU1favOCB6aH
k+nJejVQS9N4ZdB48qtp1/X8Y50ldDTWVb6SGF+gMl1swsBb7NV6wz4p5cFl2iROxi6sAyiieF6e
b+WlemBgEZHlwzKLDEw9svjSTTGNtj3+m3yijOiv1xw+IstHb4835ttae73uWT6MzF1+6xCLqMnX
FYQbUel2NbBHuVAlihKyGCBEvjIEvEN/DvEABzBftWiZwakLPWmiwC/XnPU2FWJVa7v6SIec8RMb
Q788gwpQ+gfx3hR+3vW8Qde5GAhPaIs8G6rqQ7Zt3z7E+3+16rjPevkUs267VhYYg6SYUllmR0oP
iZYggaNJ1y/0LwncQR4hhLRnhc0NoJ82Ux+1TZ7qIkBBuZcXYoCN33+jd0Q8tu7oMAnFzNImfb+i
4PqVpcguYNebB31r/qhHs7YalwvzZum0szpFHPV2EdY9t1dKDgT5uOB1esuq42tcrk7AMJv91XOX
u88l8bkcKncfYJgLGYR3nYy0yZO+a2WRbheRoPxvZIsIh86QyidJTbBaXIFlXOQVv7LgAUxfYfNq
SXggX0F6ADVxZHpdBkTmpC/vDhHVuIuDNzzcKCaDJ+od+xVEDihHxnvy5DxP+ataxslgfhkph4wU
hchGbMOhjl4ulIKku8WKoeKGnPKLGwkVVabrYCvhc4pmWlBEoibdh5ytGoar8hWc9uVqjSazNxtc
p34DkhPJ6O1a+bGdfX5+4vpR9ncZdY+/Jl6WywN5kkZd8oPRJrfIdf5sLSV7XzVU7GtasJ7wjCSx
1kX1ENKWd8SzfO4AB4Jvfz2RKDYyNgLJIGYdUljG4PqgLcrjBtj0JRFNENcfIVmB/6mJj1YAM9AT
yUjutV9y2tNkMWun35yBlsTlLpFDf3Nb2GhDxvtMC1PjVhM6yckc/i4shwl46TONM0PnSannD7LZ
SU7dzDzFfMGnr7HcPkU+5d2bc47gNOZ5eZS71uwduTyMRg71IR5v9zc6K3zKCWaRmvkHT/B/HGAh
36KbkgY+N34BRfjBuz31d3icjmZiXySY9iSEKJh0f9/NK600Zcr2HvCoQmacAICTxzF1Elozf+62
fJ+6X/Hrdv6cFL0INOo9vUFUFrjLPDgVrAmwRG+KLYx8uKNm1886ha8rfO+In2QN4tHfYJwuT0xc
wbyogoJ+9VHIjTJ4LAadTVttfRpm+0geXNMXUSaU9AuPxjEY1g+a2chBNLy2T6e19yleq0sBvyGu
2gWxPbpiKpszwYo+Z8CH2FL7dwHI0107ZTCn22H0PGZpivTd4LMoEQFHPMUERS5J7CkJwLAaE59c
7FDMVUv5moWQ/5Js7ljwMDMJdgWwkq4KHDLIItHqafMeEM1Gjk88/hrMUkbs3bV/RApdguP9pFLj
KnS/2Ngt01VBMkEDN69QEihcqwH80w8q9sS/at3ZDLglh/nS/eq++3RDIWMl0B5W1aLGo0uzi6Vt
D42/oBQ5dlS+R8kceR/5+HOqqzDDemIy6h4+xBlBUV/1m/m3o3ClCEAp3hjF0BnomHsO7H0ho32o
SuUdP2CIXr6o6HTT1tbwVN8DdrN8BpymE6vWm7EuZnKye+sbd87IECGxDANWLldEymY4I1lv+rFX
v3srsZPP7ZEAWN4hc8XOtX4i5BzeSt5shPB87n9ozK62u9YVXCge2Reu7kQaz2xPI5wHx9w4Drvp
jSMTXjv70RNrA135IjT7CxmfjiDyVVWF3ARVSV03cxMyxHgx42o3sl2auK1VB64uMUkQS9Q3O8Y/
qUf+41Y0ZQufvSell1mAoZ0NBq3kaeorvafPPdEArXE26TGTR5Tn6MYNL7HGmyGNb7x7GFKTseFs
Iq9MWeK5w2/QU/8aPA3kfkuQVM/3hMd4w6zQVh8aC1SqljPWxCpqcbTGu3nyYcVxKGXB2Yhrcawq
fTYcc0hxyFgg+waSbI2Exh9iFSw96fhnFMWPHND5LqBJyNEmGcKacBAJT2Yf97GRK4AXJ6wKgryy
SbS0q2B4btNMbMrYQ5PGGNRG1PbvFY5olXNNcRjtKDZaBroRIHTjd3Zx02bfL4OW06m3xRG5utTo
5/l+tF2bCZNJoAxEsydFw1B9WhXq6DgGJpsf2eZ4L0Lop8rKWATE31L71S67G6DtdiuOgTvIy90w
N41ZAYFLz6ogCx/LqBzPzCWnLOPUMNmuTitScnlRqQc5z+fT1uApGm2EfNLkVwkkdI7RpyojDAf3
RpOa5o0/kSUoeQd39ofwoNGQff5sUHbXtxSwLlwGjIkORfr31W+lt/SgsPJfDuDXrtUb+h6XNd3j
33eVd6QMWpA24gjOYO3mK0W2QLWP5ldDfuXwP77Vzv+1ZIU1fPbBicIsNVLY2HqLWP8ucbA/1Obg
EoIHYPN8PRjFWvFcsMfMX9Wp41HHReRcfqVkCillzeAUSOS4PD3F/rbHZgEfWvocK5xXi7xx19Uj
uNPg7U5XwLvy7XwC5TSu6+J0zU+2n796T8bjGptomDHnlAC12jhFn/KtYnaW3/a/pOpHSrF6eI5/
8sCXMiPmxq98PM+Qs26nv3xYjbbOSH/yIo5GgvQDTHr1RteaQwtR/nki9eLNQWELcT6DDTnBfe4G
zcFFLgHjCOicRRLCvc55R+0iQYXd1vjQlcRpOMp0pjOYPV1W1ATE9crHJ9A+PF4//uH4vX2KyEIF
X3Wf9mDltEfPPxbHrZCBYHje4i9CQutKWqjzxPjlW4pNmcuWy0s845LspFtij8g8hLJ0M3aR0lhK
mkNVRKAluyQTz1xnUiY6NZ0WTP6IqO88tADYvXaLZi2T8Un7/XNKvi9D7h+JbQMq9Y/ZQt5JAhSK
VARNjQJEYMJNypiR+MiC6yhn2UzkeKEXR7lcu4SiSvXb+eqyXBwWnP7U9Cytf6OVMTnXjqX4fwMf
3AgUIZqnb+wMxH3Csk1HiYLVlZpmhxD5zCfsQ+wPcSnLSG/Yo+90DebGOYN8EVinQrK41AFD4Geq
enoKA8YnrVAc4YDX8rTUhdrwuiYG+DNeRnpctkhS2LlrikM2IRp2MP66zJqXxrw2ii7g93IH1NL8
+cF1H8RdyqaJUlh4EQQGrujMh9Z37oCPruysxdSyhX5ZWmgDHMgl1DomHyYtH1+iBU9Pv8LW+1uS
Rta4IC8KrsNPIh09lWw4fMJ6vFv4kob1KBowA6uoIm0F5cYWRumQhb29fSp5H9BRWJXlgxg7dxb8
LovUTpF2WWAe1+sqIXCyMVpSsBWjds5HuDnzI0OykxJlVEUVxRaY7raK8YyQHEfOf8bz5DYsrp0V
kwYizefY6Df4Bp9vIOGX2T0LTRErIBrfzpeJbHhOW4wOYgMx7ZK6FZPYYD5Lhgfy6QznouP2J+Nt
k7YtI94cbM6dlkko0gHn/BU3j11wi6vueuthmrkOK5f3zZeAowh68SPzFAIhaJbhInWJOfG9OAsA
3NJWZaS75ZJ2HWwUwQzOQqjuqtq4n2eCGwzcv3PD8DbK4ObjCIeoqY6BJK9guH+vaggCDyWyVjSl
8/d1PDNGbhm/xpmtvUg9hMMoSGb36THN19FXUVY9WH/mG6zxPsY4DGJ6eZDzSNwEcoa9aLdBFU+9
tTdMq8nHXsz2vwNNksvg4aRX1OLLi3UTeXQxAUbspbXnfhJCqutxVgbclxh3U5VnLDyPObxdyArh
Zy19GfPxP9Wc9Ap6O7WjoMRYwpcZPXbSjqnSM2H42zrVBZtDcbSpbbfKTM/T35O1G/yT16WV0Wly
U2GxJ3tBLAhlpQGdDXkQ+U+sgOzlDksZn8yEO5tQryIH8uS/u2LvLUSnPHDgEGNKw6j600uyQpGf
37TMq5QhixnJWzbt5xCwfK2QkjOSuwTZeByfe1TWc7K6ipTuF8ZtPg5O8uQrTzt9PNtEbhlCvBKL
mroWIydJ6BemKL4ryl/gBqYX7JaeEOgnpLTJ+9291ngGUmjF1qg5njRJniF20tP8esU9KiUto00w
YGSuYYKuNV0l6niaWqURe6sB4e4/2vEIsJU27/J01g/B/Frop3Mf6BNITd9oXAIGVv27Bn437d1l
b/01pGc8dBVexojeOj3Q5Yh6voEITNiie3S8l7sizOrM81iQNXbEZSt+McTvIgXK8J/ACZr5wCmT
ztULQeqgoZXUzcLvD7abuMOg6tiMCm5TODl5IQxJU/ySCOxemqPykv35W3KWBPimXDw7yDJMZB3S
D24FCPAIWtibJ0T54kygv+mpCq26XhjzK6jbuXzpMJVJnmomMjmRmSDrfam1TnM7B8gqd0uQqRUt
tNpvifTVaqUa74p2To1FL2dXPn8GsZw3R12/NjL7w9R7i2YgVZUm5HisHQXv2w3U4HT1RGcDWWMQ
uHH74JVg0pwF1mxWQrnbrkMhgcF9v9Ltw0nHweRX5DHbOgvYOMSGSPWTo4OlkjnEfCtFrctuZMWZ
HNT2fS26gMTFZWF1JEk9kAkRwH426eDyHc3FeY+RdJru1MxDNTTzfYOdE0LLh3P7CTFPRLj/RWIk
v88TUspcppc6AlMW7bOjs77pFeVVQPTG6Kin8WwkCJjNNdJOtOSdPTo0oHh7FNdGTGf/wc8GtiSW
OsnuKQfYU+PpcczFMG+cuSxPcnoxecAPS+WA0gMaFLybM47NQZiwf6HOe9qmKURWGXoGgb5xIkgX
FCDaGrLaKFQnYvCpyYteDpL4eIaAgPdhQST7Ij2ktjyk8hixz89N5xoePvfo442FW5XML8Lzshtj
WpjJ84SpX0a6Ogp+RT/f79fqvSOhBEbiRvILLmXQ4xY42+nwgyhTL05D+9CteRZvxcr41EtuFwg/
6WNvgk4lukcDlwHNkUSzvGRFsKzVzQthsmZWR00u983bcfiQAS+7qDayJVPrd2LvrvW8yBNGKNKn
kY5f+tklBTjLV4CK0BIBn6q0emWgtPf09voboE/lh2/uhwCpELYqRbOOhZEeOri1MfSO0fqC/ii0
9EZBgM19GhYwtCXc83qVGej1X6iPjFvGdf8o5uzMeVCJyeqENaCRfrEzszHKgHRM89Vm83YN4hzt
ZVfCCQmr6+1UEKwAID4O0tkCYjSkhqF8H8ojU2tjPzGkdH9ySpYBp91mkIMqglCoP/uDZrXNyKiu
9Q9VMMZBSU22JUKLi3mNOeWBu8DKN7y30t5gbKg3e7eqJuV4xYmGHESZI58nABt7aDQpZ/7yTamq
3ycjqsbrWo+zPYq0BgCHl0RvTohfjB47Sp55heRbbAu0PgYKcsnkajLi8Kx62ooOiCfQP8+eRKqC
PVas5tJIP/Ow0xqlwfk9Za8nTzxgMJd18cert5WiMxHr0zFEtOxBwZxEQkrFAaD34J16kC1U8vpv
kbdBMG032e1kPyWjEduEzEO25+ksPIvbTXkcyzdWEJ22tzWDcClKzHHWkfecC6shTbAL47Bptlld
tCEOqj78/TGTKz7OSt8qzPqbD9DnYZDvJePsyhm5VmZo9MaoRHD3hhZYRC8jwx8uHEmZqi7g9FrU
4ssE7pffx1QnNjPq6+ZFU0k3IUoZpgLFfgiHuUoKGUs+nWRI8sdT+AJl0K2wKEtezU7oq2F9SbBu
a+wxR6jbGnXlWjCgGDvBCvU1mLUWYltQH9Yp0ZxUO/Uppc4HXBmvMNhdATM06dzHHYQyxtIT9hbY
3nkDT5F7gmCekx1FhZZbxrOpIPv2SLaAPe0e2uLsrkVJya8wyYslAtitjd2hnk3quY/EakBtHIHc
2XXoaKj+7F1c54SAJg/Pk3W7SDE9arrX76xoG5C1bQWMVf7IC3jisDooUevqGLqp+RvMUExnHbhS
GRDbRCfEsTxRPrjU54fjWQYKG1eHrSTD7Irt1AzZpRH7g4KIPE0mEEcQVTfxh2/wwCu0XHDGZkun
Z3xXNtkr6aIOS/WDrZz7B9smUJIbOoEJThwvo6NWPtPcOxqeC+rxb/Vvti/VG6o00i15VARtNsr8
hiIxSh1BJ2yVoxXcVdzoa2CwKBPuBTVU2ChI/r6Ki/R007CWgiouFKv3aGb6YnxG2Edd5/kQOeX/
YRrkFfS3
`pragma protect end_protected
