// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:31 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
hl5bp63oiNAxAxRVUroigL/EkTuq4zm+yqoIymbRv/PHBAZ0RD5kEXV7IFA2R1Pa
COBYaAdUwrgARFdcbiQDUeHIrEcF/RAxu+IOLy6HnAxTw2Q7Bhp/C1ZJhVKsNZGR
FDZ1thMPyGk9NaBDdLVollNhtCXLMDoBGW3aSgy8o0U=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 19200)
+jip9UwtfZgGkjBY9p/cb00/WDXCQKsweXBTRaaQzuReAMwKeFQha0UPVCd04BXM
Auyq8SiGd/Yntp7vODtu9ObUWkVYGDmJM4v6+f9iSAYePSotVoxRYgEkQNrPFMK2
P4oWGKwxVvP6a4Hus4SboBdUyPevvuLOfjiOuEkrrFy5zYIbVfT3LHPoEs70P48a
xjPQYdmIo1zI22LhVPV2l2tZ9cRS3QLHR72RZ0HF9G+IO83FG7/SA/RZAFTYro72
s5ybY/SGvL8TZnDUqKXCIPKIZSoA7fMVMLjg5JYbU7eVj7h3/SYa2nK4S8QSc+a+
+t+8Jad8+8VxRQN65G+Xqvj4rp86byyTOUaH5fVPz6zLczF2t+4xzxRSGJ1cUKFw
0QKCmCOf8FQ2wWFWxH03hWbSfW2w53qajvmGshouVjbSg3tMybaatrrIEiZ8wpiT
SHMdH+frSWJKaOIKbxYcW3+Az/f5HQkHX7nqJl4EOz0ggRp10L5vExlm1jcRJ99D
hGm2IprMQQAn6x2hVhEZckoKCtSyGHIe0OLBlgUAva9oS2MK1PvdD5qammt46qOZ
7d16hxW9dSwpOqCo+En9H/1eiuE7ESfj1Nb4uhJrZFnT/QlDZfqieKy/FYuec092
gjKfnnspl5fXuIxBhs4Dlw1CFtFNu9FKRMoLgZrkIkIjp2aDKWgvapuvylCvPe+i
vl2sZdOL/v/ysiQKGnKzVI3DtB/d0ugnNgxrqm9a/Isi4CYDh4L3jqwQ4NIj0VVz
PZc8JzEOur9VNUIrTGCRwi2QWyR+5pLjEO7hoI4q10nLAxVgLhFxf2O6S2s6rdRB
8E80olj5p53hRypC9ukLKwwzBKg0LKjzkPFlEKJl5fbmkQkhR3Or9LOw/33fICkF
31iFMKY/y38Rw02lBIYIPlHPYUWNZ2vb6FlJ7YXsrJBpcD84jCQ8qonTT2MeJmQz
/qQIy/vKJCEPHNUHLRQ9yBWxiilcToafnlcD+UNlUhD3N5s6dPsVV5kvdHCPiADX
/GjqewhuECxNa9Na5NseFqjvOrzhTmVPFuPTf1ax1gP1lCCNPAVY63r+LPbgX87Z
i6tu/KpwhewihkA3D7Gk7mAze2bGqTxzRACMllDmLZnecxUtEi9rxirPWl3vXcid
NQBLefKSDF1aWmuKEjUODFIr0XbMHyLTMTnuTFE82vD77kN4CH9W9fwrwdyaeeys
dOEhIelLr3GDj3DE62dHQgw7Yv+wJ1aFSG507Oeyow3hxgis8uUXrDxBT3oHauSp
rXU6ANJ9UBSVepn9M+EJGa2PVuEiIoAHwajN2JtVIA/gqzML2I4oAaQK29kCkYOI
piC5doPjhsh/MfCsun21KfOxn5LHIfqGdGUnl3G/xev5/RZXHsHdlIIevVm7zgoC
EtzE2/CzV/8NKJgD8VczRQv8vj9pjfSPhQOaoGsdueRI7ymyDfg68kJb0lvB+Z3+
xMvSvAjvAE4RDvSgGf/h0H7ls5GIT/Y3Jfj1B8TQHC0D198G/k4XO945vscyF326
gdWczEVVI683hGJpT73kXBsB3Wf32DfdD451Z9tYn6m8Bf2U2QU+Gd/uVYCw76OV
+NweZd4AXPD55E/ZYQV3THf7XLBrVtcUgJl8XEQ2nZnES71iM5k4MvP7XbBNnCjX
dDNssqBULKb+6/n6hm/zV13dfcfSNw6hFo9Hsa7pfzjBZH5RLXP5aAeXJFB5/IWy
/HE0MUf+h2XNi/Z9R0Mrl+fpwy0Xfb6XXA9j7tXynr04u1doddeysVo3eH82+lik
aOavFfKohKg1hl5Irj6+PEQ8cbtcLz04uib5bEzqnID4YMo7urxwC67M1dnBcRsp
r+mzsGWn6DXjzXKJayz6xexsJDOhabiqn8WZaRpikpXdhDR/PP7/ksr2cRrEu72a
hta3L0UDURF45BwAo9T2ykav9oscC+f2bWcNAmWGQj6sSQWbGHtzI2JjbbOro/Dx
wdXgAEXYodTlY8PyyhpiFVuZsu5oO4ZJrqtbOMF/y+ZqlXR5kozbMc6nCNFk83vn
Vw+KxcDMajSNLeltTmU50Fz56OlD42WoG8H9dHRpdM3ecXs7KsoSBbBzUI7VCLh6
C5oEmWrS1ypE94DzRsaFzqmxK1jxf8Pu2mzAiBvgHrEastMUaYqPQ98HJDqeGH5C
Hk65rRTD0XejEpdkJ0g69vyNTksDQwHb8eddl4Sa2ok3hQoJiseLLIN4mHe0nt5P
0zrkqDNERwAR6Ir5ziaNdKZ7b1Qz62m0Ur9OWG0XHyTKDx8rnb0BWvp8fNeajtNH
5X1pCWGcp4ontv4CVugW7LCcsZpvw17A7MBS16zjzQZEQsZmqKLY8DP0s2kR1vDl
EFENAwo3KcXNvjr0E2govU1mS+spg1VR2tWHFP8pXPtPFhVMwAbho/lwe09z9HDC
1/k9NcIzvTFT0leieF0YB5ttM4hpaiMBBr+siVpE8uaeDK5WN/RL2mmZEflxl7g9
ZClStGNTR+0TIxcYke/IYTOh8dLnznNk3iRrm86U6riEg1zE11X83vLIS84uU8M2
x6zeGtL6L3BmW6f3fT7ZeQ6PyPCM4nF0vkAVCwLwHToIZX17KD+ia2pGpsxpS4QJ
EKxyLRaUNu7QDUqSrJRuqw7mlqAN6+G++dDM4h42UFC8G3UiR2Jn1F8oZmSHcmdW
9GHEejHC/kkN67RppV9YyyI90ZACGScul3vblSMplEt5go/vCtX1cM0MOmf92uU3
0ktHMQtjOD0vOksUAyzcl/AJnlduIJvwCzvL4cfORg1JY4kRUHYix1+N/2i2tEFp
GSkB3lB6OXl+xD5G7RyQmAdt4LaJZgDuxCfbR0PEZ7dCTqcvMOnVp/NBPYECUmM7
nutGiuq9ZtQ+lQ0XsQYGS9LdoTNYx1v7jqP2YT6XB+zlTj09Xm/Eex66b7zHwICf
5eDzwreck+ew/QnSzMCLyp+yjiIX8AppGiv7E8xSUwvKG/fKYGfJy0j+9Ga9HFJ4
jnpWfyFrBc4XTt9Xx5SLVXO9MfYh8RAfmpQPDlLZuYD7xDv1xbtH00rJnFaYGC6h
KIqNnYdcFZzS7HBmi4DcoMvAEnX+/cXU27Qfgb6AK+byRBSocwpnD5OasGg8cvY3
QzPzKLi96dVhBtcmvvktxM8tt/nvryly9frvWwkF8C4nB0BAdXCgl6MNN52417YL
oqbX7hyB2OHn5ULCnT8d+pFq9nebaPRTxqCd3o0UcwlWAmFbmp1NqYzG8+MXzQlE
yGDQFjB6AmTsrAc/FoOap7dsYtq3oHP9M9DOd9TRx4cFLE3Y1y2Zh2eouyBXw26D
gyg0a6rLCV+CxvUfD4wFldDT6DGBWnYPOYQ5MIE+Hh7ka3TI1Z9Tl2HTpa2WDiSR
qrtjmZHkhELZJcdxz7tdPqGW/FOT8hwCefxu4jLp16Arp2CncD6tEKuX2V4ZcTZR
UeiuSXNgak3xKEL73GmNsC8UE1AsxkU2PJeTIHYCvd0CqRsRq8xKWojznwc6rG7C
nGo6SS43HuqCUMx7A6+UrAhf3yfDLIkCoRYh/hYZlQ+/Jg47hP7UlVfSD6VSoEhT
CimoSEMyvwnesS2lJC5S3W7FaAvrWs7shLIDwTwysNq84+KhoQmVwgJlPDbtMxlU
k8wXq5jtu+xD9S+qU0e0u1lem0UQogQOCIuDgItuDMdsTkNcB1yfGAy0fWXDPk7/
nJkOf+sSNnfQaplSBYHWnGsl+EgAQaMJ7NOFfeRaamaYZt4l744GaaY265aD7In4
jGASoWTlnNLEZ3pX+Q01LuMEBWmmu274sMN9Fh8fQbIruhy+CWdFKWL1W+n85N4g
Jm0xb8r0JMbBJKzFAIHoehJl0KMnO4+9/8SSJwy1mCtS+P41RbhWYV3OOsAsl9rA
sR4zjPiS91zh4ncIHusms1jRj0vhoUkcbKP6St/PF00nr1YnImThDACFXpdRvOdn
xPL1dh4P0u5QDL25yvH+pE0pAod+yB1rBsxZm4pFJ+yA0fq8gIDeo5BNlLfwy19N
XbnlUocVEDBUfqFEtJbgHrFZR9+S6gg+DVVTmpDAH4DfadFWOeprqub5n8Uwm1Vm
ygjraA6z+qS6J41cRMSM+YF0UwxsQ9LlyIEuUbu+QPXhc/z9a4LspKc5EzTFa0J+
sA9hNJl5s+vYhfWXGzfgaFAah6CkyPGqHm6wA8wRxnojl/RDO+ilc0ujoegGDgAB
mrrtjkAcEuT3mLYfTpVl8RFsD1aJc+1PetDJyA0CJt5WJwugDufV82ZcOTi9l9Mk
IBGey8r1kUgVdZicOBTZs+jNwNH7zq80B9KKFFXOEpFQODVPBwi1yMXYfv38uFrb
B5uZ7xq9dKBtTKWvQJiijr6s3q9a9V6F5nugW/Qdxk16VEMctszFqjjRaUwjQrxJ
eaj0GbGb2ZpXByJLlUWuLK+Z5Wq/ept1PEd272aUkNCBYrURcKxMC34zCwr/uGJX
HrAKPNIuBZUmzSPSiaxI+8Ard3TWHZO8EmzfTMxnOGZmNOPBdwFw4D5wNVWwqFeD
ahi5HjaTf0MIDr+ASBqcFz9MH+kqSeNaeRB5c5J6YYkOHcKoCg2e7IHDUrXGmc0P
I3hTB2b8S6ZnE2YHeFQJ9Sz9dI3EpBkaaBDJ0WuZELFHekoNaJlaLBAeITHwBRW1
lcrIWi2Zrgpq4miig9BSqt+OIE3r3hx4IQU2tSZBpZORHOwI1CUJyaClBEa3bBAm
k1QY3k2NmxbU17L974y8hURclER3xSMZ2p8LZIZCvpr/7Uln++xRYAaphssWjQcJ
mFpe3auBrmbKmGuikyM4HBqt9Keo43eE21jETrCyumAzh8jitgprB6S6ZF1jNO2+
//KCOsUnK02TUW4CoFtMMgPjEqz5t/ipOUSzLjF85PRIK/ZxFKyYg4zybpcmwcWU
2Nqmtk6haxBrUchf/zexreCJw94S4QROYO+DU1nnmf/oiAMAmvvS8aKLu/lj1Ta+
z1iFsYeikQPitftYVoHZB30kVl7FvrA2s+uNnVnd5O/jguCunJ78BYHaLSU6+xfc
AWC7YMS2UkwlYZksQwMEw9fZls8lU05npyP9qLIvOE17wNdHeI5zLvfg4uoERjZ2
Hrg6pgszjVPPaMAnITp+UMZIQ8wjbNaWGApxygVFaFGziA67ffkI3yB2HTzBZJ5m
f/b6XsCQQW0btg6FLz+DyIAKdVfHO2gLvG7FDH+5vTYwR69Yz9LLbS/fi6VpH4Pe
jwjqpmNhFSC5YgKPOzOdIT0bS3/9Sa15XPyYj37JXdvda3s9q7VheSGyew0BqQqO
3o1L3iKMcri5D/ZBeRRcbLYsgV7hXXhTiXA/i+U8QVkdTQljaU3EVjZh+Mi76DAW
peFVXH2eBwdiy/hAxVT2hHe9KsxZ5pBvl/ggtgKgMHKW3bFouSc+5CiELEeZ+a6f
gtHOeYQIH0Q6fD7uvocSDl5bz59ohcDsAcewPox+l77G9xOakfDGrC4LNiJuPp6Q
H9+h7xr3ahSxrM1EySbpznEjjarhhMIRhGS21IA4k0TCondjqoaZW0WRrVI63v3y
VqcMs1OOtNhq6Qj8nHu8MJHn1xixRwY5VaYTvBvDy/oigR05yu7t/dZXuXMBZmGw
ruahctNOo9zIfMVpixTntu9d9nro+aFxcUdtQOpBQFMn8g9JENMVJm/zSbo/inUw
laA7OktF5X+Y87TlcQQAJqvz7ACxcF3M+WBojyvIcymHnED6SUa2WoLVdXGjw53d
6+6ssDQmUzzvcX+l2OyOFF/7FyTfnwbj8R374Gd2YxC8SgK8F+Pkzbmc5yuUmLDI
TtK4+HPNwDysATqf/j8/yum43P+GzaCXRCOg6XTLhfripyRVFTFPk8OBGGzywTkw
7v4/G7tWUtBw3Mljrzg53jkJSHk5n2gydX8/ypkWBigMBofGCD1oP6d9HWsgZMj6
L7hY1eDqy/qJbIZD6Vl9sNTuxGpwhLVZOCGwfxIUZMX9l8L07kCTdqWFj+5dUX5P
18OgwMWd/E7odh3FFhMZZmoBGoJtN9qItqnPKqNt4fI+k7lNdhDYRpxQUs/O84zh
WM4jD6ODfl1lULhftiEktTG72rq2wWEAadDmAw3dwAk4YmKxXEDST6FH5BM2b6U0
TSTFVD7TE5YgQ9jtaXgtZ6bK/7yDPX+Q2tY36aEdk2X1hIzN0+KA+gfC+H9mfIWj
dNrwxC0xGuDCMbVCOltowA9cspz8E8ZrQT3Ll15i6ucaJD320e9XeTa+VE1eFMfW
y04Te0g3kvjZezJmikeRQZCum1ykStFd+Z5pnE6ucj28T6lW5755GwHA4MeDouen
SIR1vItgRWs7JgWevMpFm9dQ12rIXzdLaExbJLi3yPQoVqIjQhmQDHREzsKKioMZ
yPv6Raoe9pzYhmcfoBa4jojkm0tbKY6ij2TrvZGIoKEuJ9TWURrBqRunenqwYRG9
i/GF5t+KJamBNUin3MZiBLYIZfEF/mguL1SESYvqtOuR/VXby77Z7aP0e7B/AqWB
83x7owNdgU1uPiTbiH0Crzaphm4gl+zhl+WkS4sPOOKBa2CfaULSEnN74FjriYQI
gUXsS4kbY8AEhCNlkxKFNpjoX8bUf7sA9DYGCkAW4M4Ma59oiPR0UHRfM53x5swn
j0mgwEsJdQ93eHkleeomGO03IvgeNbyXocId0O57/rVQv4XdY9an5fWza4YKSscj
fY0ySUYGUshTpXQqxSpWpC9UpFWr5L/iuIi6+JIqRdKEZkptFGDINBXwRGZdPqw4
9khcpsGWs5H+v3TqDXA/lla2IuJkx4fWi52Cwip4wT9btz+fVTxWZzsUvXHtIfHN
Aa5ZZVrqVZESaO6aDI9PfdHx4dmEwzvNiUR8NuPUcJB4ZMgDnUybRkWoaHSAjbAk
HCzC8JQxjmsdpX5ePAOGyLOPpj/h+8AXrJd5f8kTxVuK4Lxz4nat/kYJqbYrXLgn
yrwSAasT1LTFCu9uRFOjPI+UnW50PCd39cUlAOcBwpeNfuG0CGLCMsuhEUE3cksP
QJl9eGvot80f0UxNK1iIdUceSF4GAJh/r6I6znjk8K4vN0gaHuj8YqUL+Eu00mDu
yOx7IS9YT34XC3C16W6BcwKDscpxje/bpfVK5jnq+iMl0aKV6M+J2dy6huGdUVQ1
O9G2+nPKMBaFK57Cyok9oFLVtFmAnc7VIv5sQvITggeV0NNa6fxA1ub/WLs7RW52
14jvve154kXrnyJqOwP6KHBoVwnsy8C/0ijz107DDbDeUmbAwLTzhVgPwhOIJsQZ
JgK38UBIQk2xuP1g5M+7Wmv1A4lQbSkK46esG1qCLdSV3JwA8d6oQ+CZgOYWMQW/
EdKxzdbEXEMv80DId603GycNjf0kNaA6/6c/yas9kyavM3Z8j2ZZ4vpY5hdSMWAo
FqikvJLjeMZNQSoFvmwX21EED1y/7Ne97wtvT88PyTWaAoNg/FXT8aouh8GQUJs8
IwsLjJQZVH2nzroCuH/nZtuMo+ot9EeOTNcEUzZtWWsl3aeYOuvivi13wj/eNUx9
Vwt8j3Y3Rd+nD170NfFIwZJGoyjeqWpurRaxRRV0m7F9yrFv2pTny+zQX1B5Etj5
GgmVxI+M7OFGBXJ0a1P+AuYDcjwE0yRSVmWirHbqO8LmfYyym1S+o5Lds0PUJPCe
Ipjyfgpdm7Q1fvJtqZz1wTgAd2FhKIfsSA09Dr9f0YSITAY5Sbqc4ZkLUGyQuP2E
8AeDjypeXyoUVUu0lxYbY73TOXgc0EJ2DNGB76+vRNJ3Als2wBEhjHjOlL+1IXQA
wplTm8hDUMIDSY8ci3GuvfepHWd4cYzCjQljRru2FqjBk7E6VeI5zFsjlUnLO7Gt
g6OcO0vQ4TsBUGvS9SsO0D6LPDWCFJTAaDFacwLANG615yMG3CN2fjtjuTmOQiQo
NkzeyrFCIsoDo272AQML5hlVWm9xexqvLzXplm/7rQR9PdOIIgCKlYI/OxdsundN
zZCe1ZPpFKpN90oqYVCYHBKBZkCccp3h+NPf46BLlULzvhhYlqcyrnQoNgBRsls5
gM2/izT73HF/Zw1ma6of2HkYZ8jN6YvYnXEQWqy9+dxvO7s6sTXxhLp7VuG2Tni0
UX9/UuXYe5qqnMzK32ZCmk1XARUos/cb4m5Nqxe75IHD9+xhI+g74AZKVbJ24vc+
lpno+NCRaLP4F6I3Z2zxCgNxOllo8Mxq0XHHKz3IaOhPNU+9smIcQ5yVc61iCZya
/oP0LI66PNBS5TxhnqtPtxppQOvWGe8ewVufUfik2ZMLygcOS7BaNCny4shYxCg9
cpIgfUMdDfuG1ika4iFDM0HDgYTfNuy2geLpKE3ixyfLwHaPlAFPl26B+NQ8w3Iu
HP1u12EhfCur52RztqGbWuPGWD44IilmZ2wl2FjLBLbxBbsQaUUdp2CbUJk72Zgm
8EkC0WInpRvbaJ3ftsHu6VQWIqCDwwnhkpmB8o7LIhGtOaUj05EYnZtyZyKb1fHE
iLoXhb908F6zSdqdAj+rAC141REG36TaD1BQNndSc3IT6dGk/VyH6BhucV/+TOgX
hLb5t5QLNtc3i3lFUEtyK2xQVVpU5Iz3djszpXfMBoopKKK6chUNwWt6mg7rQgnT
f96GNHk4jewluNuklb+fYfb6HbA0nR6Fez4xMr8NhzIe2VkWJgTuQXJBI8uXQY7L
RlJfg+6ehGJSw5E507jSumW/Xo62y9Dh+Pp5cEUV2KcNbn7VuSVyxDQ+XBHoORUC
a6LNabyLzSYfPU6ymxARHFfE9u3fra9VjPH8ZYURW6li6B+9u1mXLLgTdYlNF4Mw
eVK/1FEvx6l3j+EDRY5fDfSJsfn6pfs9DwRz/kCBmAoslwPQIQ//JG0RbUT98r+s
4/EQtYT2xofnyuHIEAI0banNCMqAy7O5GfP9CzfcazuH6Hg6OG7ChCfc8smBmABA
QTAIs/nHpaRndoU7LKvdf5vffb+dYJ4kfH2ujfwCZ00PPFnqR0kAHnBszGruy1hL
7nbQSFMayPEL0PvIveCUwiTmIUfil90kIbcEekvVq5/+W9DLoNLlR48q87N9VPDR
JE58aO1JuLURbSVF0GfRJIo4sWq1qZy71t2DTE963ftBA4kUq43koAHjJzSeza++
XFA3LpRCcLmNtIPhYfZ70NMGJp0RFuqoBs4ZB/ECOgW3FfGGpCYir5SUlxpfaMVT
xNYEm+AscoXxg2He0cF9HkCG3xQwazUmNpAcjYPWSeO27SGvrGNpdDoomrW2C3Ne
cGSYWIwZ7+L4O1jKjsVODjA/E36ik239MFCsA9pqg9JGVVjGyWTbxwJcYSEDXOoI
jI9JXZNozZfGn0O9NtWUeFO3/L5aBduyo0Q2bTinkFfUHORurM6g6sU/Kdh/Znhz
sN34Q2XJ/w7Ex9vrdzZRvwTyGzTLQ2amNbjkpTZTUOsd8WOlelUmLR7ZFrC/2DJK
jn1XK9vYs0KMOXlDkaf6oLTtzHwyhZ+9JAUZvwEAnltQ2N9jVoZskNepUfAS2wLI
vPP/hsQBzslWT1fP1PkRN75Tm+Vhe1lqRP75d37sxF8RXg0KZLyTtr6yVl7hWHO3
eRj7zy/rTUCsQSPBlXzhiFfbnRhiWzEucOxqzqiW/ESbaYKqStKRQzqfkrtjUiqP
sWNGxQK+UYtvvPMCo0jD/DbkFYz8L4YhPPGMAgHV9lGIRsqKvBe+eoTSCu5UfbM4
lsWm3FhXixJQV6qqgLJ28R45WqTJUYgQxXzIFtN2A51+ZbfXAxd5U9deqTxN8LAn
eyk076Ba/4lWGs3arUXQHkxQ9stRF+gwcUvISHiGxuidvQJisVz+WZIhLAceHdXm
hbtdepBel+zDUjxE7GcbQuYkjkef4/b02z3kmYI5t7JRHSmgq7FH5Yb1Oxei3nAN
mxf2/AdMfegic2RWMpcyjWdocviI6+TSEa6O6nL6mF9BO07pPGt19BMPyegFJUh8
3nN5ppmvGQCcVLmt/zTwk8BM/7Ptoii72U8YeYj2ABoXt1H48RsPWptfxmw7+mCM
5o4i18fUuKnxcgNn7Ac5Vexb4L0LdbSAQNjLGOZC4sJncxjlL46LmuHrLfFJG3w+
koVog2LJqxR45mq9u/I8kfkNX8WWgNLOVlbNpgbuHyxFNV7pjI9m2U5bt0QNQKSd
uu5Opntt+0TGMqXSfRNDpcS0ARssXDNSw6dZl7/TI0cBEBhhyu3gUpZfVWzGP6E/
wEVj5/VCIwRkkf3+WrYl7DyBK7dWSBO7sOuFWRjA+sci27n/Riaw8Aizr5ViSQME
xjqXUoJVhZCCiEr0U+UyvzSl8RfFFFL34JImJ8spVHHzOdJdVjAa0Qxum2M5aXsw
i1g9NzSRJHzJGkyBDLjwEF4zqJYPx/M6zLzXovzDZOKzea4eLPbk913g8kNRTMzy
56awz33k74bn0DRiFBk819vYVZ2vseIst/Ffrn/Kqo+2xD1Qdk2xtzxMO7avpwAL
ZL4jYq4ULN2FP7qwkXik3idUFeYwS5z2Z6HGEU4drchahRReMWgKVgoUQ64E4eH/
VXXwfHFSwI2M2nuYQLojFyeNq49zghX9YMmGweASk2xV1CNaKUgMZqAIKSGUAh7d
efCDrFWhCWLUD2JcCkQNxOoNOemqYGsLPybyd4YsN519D6TahGXr8pVS6bOg1A4r
duecDRsRbBAUHwYDUEC9RGbLgAeK4aTd2t1byVI/rJyfKNDHFdv3l9VVslrkSrJR
9GfSkFRK4gkc+PXrS5hy20mi4EA9dYtJvbckReqIr2ocjynv1YvAnZQBQvnruWqR
SxiH7oGDIGDwwS4xx79xTSkf2Ks4a+hEqi93tMtLUAytNQmY4LYmXc56N3vJYAda
WYG6dP+RjCXDI9o7hOWAfPVKw5V4e4YChSWcQheoU4qMKQ1TZoMCAkmm4dde1rtr
Wpk7dy73bm1uf0KWdwn58OsgU6kEaTGLFgX1WrxYBs9T6ibPBD4nQMZuJrxnj3Po
6Ng4HegnHOhSvefZzqEnEQMFCz/lg6/yL1toPN81zjt9txnQnGfXhkzcGVThM+DO
4hXj2i619fSKKW7WePgVGgHpGtE1d1WlcYpbNKRmcGOpHpuovDFmr/FrNq305d66
WkWe3g6Y1UAL/8V33RyHAL8hDiDe0tXu5EXGBXNgEWLLjMdLwZOFCD9Fbk9zLvbN
YG5K6Yv2vqYOyTKoDvOPKnDGrYjWFsBAAhD6hwcOCtZiC4Jc5YNuxqD8RjXBcTB3
PSw2n+9tC4EF7MsQxrKIQJVt6ucuKpIPFf4skJc6OqiXuDKr6RmBCj3/ZV0Ay5Mc
fHhUem47c0FZFTOPbLX4rW2SCf43cPGsZZNktcmAb6RGL3uJ/JQhzU1xUQPCg/C/
ahTsKU5dtxG1Oub5sSC5/eEWn/Zzct56OsAH/p3R1kBRV1lAQHFngjCQwMXDJmxW
8aKG1ggbuILE7emDuk9EE6OQAUUZcbcA2CbgMDwXv6bPtHbcEZps40dKAtE71K6x
gfXYYUBqEnLhVBFH9tTuqXi1pEi6Z2DGUU2RJug2hYjcEIo0UDmtoc0eIRkbxUDy
ebP7L63YmjHWbz9fi7fjJP+Ia9Wv/jrurUAqFRu9IQkVCPBDA+yiAm03whH4806X
a7F6k9briOyPT5rtysL6vgSaLJCLZLMxG6SM7YuyCgcFHvjcysdQgkdREvPYGDOc
19oh0AZma3wOb4GNT5MnJVVSw6TYNKvn8/1ikRpZNQJb47ZqKXuu6Xh7M1L1CpLr
95lgDoQIDMBaVR2wqFRAGR6D3oaeL9V2mSwQ5GR9VqJ6/zwIFsGttS9mNmTa0uB3
uXPEDJVJKYozGPv2z99ttkPZAx69rQ5UxMms+Ggy/UoFHv6oVCk8QCrzOYgwPKDp
yMSYCvZ6JMFtw8fGfgDU4I/DZi2ntaJP9EmnEX8lZL0AbkNZaiurY9QU6G3tJRMq
arSF156IYUDNvouPZntx6ikI6eKMnXSlfFWBwncmNuSbl/C17q00d3n8J49wR5QO
BH1jU+a4lfX7o4GaMOB5ckbXf3RXl9WDfhpSRQ8AKgspl0TxuFU154jf2KomKqHN
5RRS/5Li0WHKIGtkzNRP1G0hhLmOAFM3psJPKWBqthTFxFCsUdHBukwQwcllnPFw
RX8XNod1fdRi+wZhasaNg7ZJKz12GbKOzclMo++uTBldRMDcMxjwGXYzK0jXb/Vv
r22tPljA6kQTMff7xG9aM7kMeR1jvGghbp28lZOAAX5XCnvJYi7XvNl9b+qplwmg
7n8ZzaC6MKTgkrmVNa4SSju1UJ5gWnlIvN9juwmdPEH8c9qN9Bp1+Ww79kKr7FeC
0awkAXii+1w1cZc/MAbLfSJ4oU6UBx1mwtU2JM92lPjV+gcI36m4wQeX7FJJaFP4
HoUDuBOHu3/CGAgdB2bmW4q/4Mi4ZfP5tvYEpp9jcdhdEtW9cx60Zye2mS1Odd2m
3FbSMr7xn/rcCuVA4HQYBt3Ay8xp/zJyLGBN4DptsfUSiuaTNdWiaQIMDRvWLWnl
e9yiuju3qP6HsgOK6O7uqAqf93M8rCLNY4gfkwqFOBekiUoDFxcm3scKZU4GVX8b
caNdAC5mzdRufvF7YSY7oe62qzZ8OhGC/gPDl0UoLR3NqF//P99toPqhy92T1W/a
4mRIA2LSSCIZH7t38eWnCgNDSlEXlqd46FWJzzRw5zPtw3eMbJ++jZIzSiAWb4m9
bUhdK09oRkN+66XBKrQmjeM4ScFIN2xTXC2pObQ11E11/sm8AfIzD6VCxmGuFsTk
O5lAI6gYxApJ1AAANVsEJGuuCdqik5zr+BU0jDjdZwkLa3V+X0i9Dy4OfmXjCZhD
9OF5tNwwcG68Ut4bUnzxUrWJxjXkwUxxqZvg9aX3xAtmQ235Aq6PjXBfMhMhkMZr
JWXz6UInB++ONG7Q+8JQpdxsY/uXcwc27mlGs0mqrE3yH5Se7QRyDjOcQrLpuzCf
P/nwIxTfv9d2cYpAkvF0O93sZSan3mZmCTQ9yM1uHvFNtUrQdUpCJBhurxKyhYK/
r8dJoSRHgZ9KYM+LnHWCxZLoyapucQD+u+qcuNFz/VPcGaeM8pJa5EZqUyT2W5Jj
zoC/Zbs129f9xsXm57rbZ1iOepPL70RSgqHDH0iiWwK1/oyxESsEneskiRPBjcFr
gZXPDoPyRxc3myW9aXWbVyMh/PJsXpnbkhJGKbDwcgdoUlt4hHuRsbETzIk+v02U
K38ypNsrKQt+ybw1kSQX9WtuMUmGJVLRJlnSyJeFRcf/8y5uEPo8DPPoFVjlmLyx
J1ufsEd0NXpQLJUgzMDAsG6xpkcc2lNi99BWCSZgCRus2LdrJTkgSoUES1bIs8Yu
ecxjeQ7A61EtHkZO4QbGFhTi2OdBJZRg0FgSNaCuMwKXtsucuVGj0brzchBxVwTV
43WBauULAa+QMzYMRvKvGtpgYTCjM1kYJ0BMaQ9KvL0AaAZh4niPNgPcB4AMMeph
EPWRW8cREefBdpmqrEDOMZNJQuKE4ZX+awr6cGHioZv19arM0/D0DMKtiTfvDg7S
rSrDN0eYwabC6YAtAQESDTkFBWV9JE9YW2lqqFFAeJHzC8kqXGLRlbBoeTyyBahA
L6sT5pP2ITmUXg1EouNCT67e2CYFiJ47thBmNd6IWoDoc952dPojo8Fl14ijJBQ7
d48YjKYGAGj+pC36hMELhBoTeGIEJOQvTv3gh0crLoQEMUhx6zx8n5BwhQKsYUwR
L3j22q9aBcboWBugxarjJ9nLYYFnllEgBFilCTuqkDdi4zUnBLXoeLHtjRwfgLNx
fmNQMAf+AqXjpFo0/aXQeTE3c3eTNNfte9s2kMf57PCZsgVpeufvrd29DU3Pdor0
5S2F7SRrZMBT9YuvxjLcPaJkNQbCTrkzO4G4UbRK7yPns+fZNRKWlH90kQLE+F1i
0yV2lfpdWoZ5BFiVJq+IYRw2+ShdFHld8UVMNGxzv8v3MCMwThucjU7SS5ByMMdH
lgUFaMxFQfx+QQtCkSv2r/GpDWpfaOIBzwhnnR7dN+IvFCtxImOf6FX+vBXsxk2Q
i3V4zEc1CWcxu7ciEocwviJovBldo16+g7ZDp5+Viqw+1cN9KyZOktZVZ0XOZYTP
FyM+uG8i2dJUrrPEsU1H3PJkYUFDPSAd1pl+TDnXeNkPmi1vUnfD7FLcnMoGNWGP
BUKbRMbctAvxIPpPhWWpe1LufrktQoRgoghxma+QUV4QsmfeXdnUm0zbU7ACFpb8
fBgn3AY0onPZ4tPWqHLvEnkodkCO+KNYRALiKskyEDrsUpfqtR9E12ifuQPFOEtg
mCDciFam1MlZcZwtmSLJXsqWj2Yx4ZUwJLUOdWD7n26rgqm4aTuSK4M2aw9iAU+R
aolQKE1yewLQx1eCOFsRCVQjlh9bh5A06TlRC0/69PAXTtq3TpWuKy0UVBJLBaA3
0GarvSfdsUXBeVaJ6hJ/+BfXMO7nqtNe0Dqo6Th3Su81L9p7GN3ZILoEYlE7XB67
GIVuZB0zfVuJb+EzEmgaJ6PmHXxbyAjTt22uokNTeT08/y9d8+R5NUsksPvDw9tL
Mcaz6bpU+D+kELjiBNBSbWirjSd6pAtmbw7kOIwTBx219DxEymRmZVAhLMshzl1h
LEqHMYEnA29ltnuTTV0dilFFHTS0KbJQgiS2YfJ0q03Hb+LDCr3hkiVMUHGyP8cl
iLGPTShSsl6BAlhk2tskYAzcmDlW16hwR1U47BbuyQgitR6ZLV5YhW+KGYDuVNmG
O+hKXKoVkKn5THIhQLtgXuUbLGn08eKcj7u3lUkG/+zLkrvrNLMXYjVdu6LQon6b
WZpzMn1gZuahE676Yzhl15/QAimj6ZsqreylKWtGg5B/CyrMmcge48ifUBv1byPV
aAYDG7hjtOtIk3GuXpcHnteYht9eyTsp+aidGhUo3hXaiQ4PCA6BQG0lJ67cPp9r
5ctbCjC3FgisMlHI7iDKfFHK3xXK54t5n1QPktYj8FO9FUwq+gSmnb7kUc4IKlwI
3T+cGrCbYoE30nFdIddwSItwP2opCZktsJovrakgo/8RBxLER7KCN626gsnFeXyq
vHadOvIZLrDGvfyGQFEiVN8eTlsEPc3GgNebd9G99ZoR4EoTAXA/c3iVWi51FCWR
nQT55wIyRv4AfEOnsVadBn7yzhFJ3qh74aiB7lIH3bVFOPDKFlOyHTIf/rdxTiGg
tNLkgXk8ljTiA9M4J8szHS83A3ak6Yg6ZE7BvXLuM30r3lW8PP3f65SWIS+hZs0A
dgQCP5GO8eDybvsBXh+dRAFGxI4BbBpOYdPZWySdt/sBPcIPdwNK8bcdeUbVk4gu
SBnmbk/llg0hjgFr3qzqsRgi0At07Uw9uaAse5TkXSGEhTZVNLVWl//Ee7Zd2YeE
qDV2o4x57s8k+XPx+iJNk2LoBFo0RW3Ub64oAwEMJ4wloR7x6ZvZZA3RhQJ4Qk8d
TDo6w4bvTcDtrLO986RdTlzf0paScSFO8qh6wpjUtqjI9eczvItTrkMk1V4PeCPy
UFAR6TQPpgXuSvYfKaeumsyOHFCzxSqQPMPbxTOD6hIJToW7HDrPN7DrP2ORQyvV
24hWYfM5J//Zha0+nMgbNHlhzzUFM5MQXYlK74RRLwXV6vFp+Yxy4x1DfIRyaTXT
znebJS0/b6o5nj1Fl8VVF3i0LtqlaOYPKMODEb7ulp+3ulZCudUWVuUe8vJGzsvr
390AHaqVvfTujMoD3q3KB1jdWuHw0PWxGy0xMeHZ0kUBzC2LKpO1bKs9NBgJRVH9
uVyufLGMio8eAdegTUqFy9bltnHIlIpks2E4adtv1eOeyTFQjoeUeMHYxIGUjj1J
qx/Q2US+trO9n7+O3MNsgBDbRGnFOJFXTJU5C36O9ksunXXihqc2RitW62TDKzxV
4IwvOp/0koPrbGUFSrlv6FaDCu2z+TPqQMKGUN2FSCmfQze2g4XuB3+CUE8pOP4F
5uqRsdprDvj57xvy0tzIJuwleE22N7Xaa5PauCE+Tk+hOosmB/l7bedFu4n6EqVh
46b+bE5Jmr1FMNsy1sF/LIxK4GAnOgPVxY1tlEvVG2AQsmdclfzAGmFYGHu5tgPB
zVwnjQS5ioGLXIqLBT5lZQuIjVYlQRsSEnLj8qplBwJ7GsOMJaciPeD9CdMOEO2W
yoWV1FCAD9ua7L6EfodTVlo8px3TkHXNnkuyPZ9mYTwEGvOJ2ggCbZUZcj6RPgx5
aJWjBlKMxVlFtub87plfzcQQY+pytjtdm+GTz2vIDYNerpDLCV/drhc8fGTSW3ni
l/AZvQc+FhSnEhpH6qaKyzS+KZvMCcu5ToFyKlAticK+iVnla59c0rlYrPvYTozE
giny4WZwim4GpksXm/s8Zb44SIvgWQZdfQkh8njqZx6p4I++iqN4CJTeVEsy7Nh+
VGAOzDXdiEATY4EC8jAB6OPByUqNFrCS6h0CveYxP+XNq1gdUHh3VkSbS3BbYdj8
eAgATcaWnkm3LaxdK4SMgE/P9JVMeRrgOxB8MCMN+ghG0ayvj5h0jAIeTkxiCFgb
Yd7U+rM8qdWcYCVeWSNDmAC3a2F1lkS4fvZ42DIMBs/mttkB+37z/YGJG6FSkXDT
jHuw3hENUQGok18UqbWjaPk6W3KktVCDXMitlmbIaJSh1UUImIJPGx95dHnTzQSd
EiotHl2Cf6OcC/kfFa8qYbaX+Yu6XJHmUaZXAQqa/6mzSNznOqsrgiQJuFtuTjdO
hzfDgc/b0/aogtuqwtW8e2sj8N5bKDjYdC6bg7RZOxXthh8qvShQeRtqVOrb9sTw
4P3IWx33DBj8J4xJw9jrzhb7rz9ODoDa4mlyyKHZYCQ700hCGtHjGyXrHjBRqAf4
El2jXDnZeuqzUTlQv3Ne5exRC0BkHXUmFK8jVspNXKs/z5AVk3p4w1hUhUkq2JUb
DOZg7vL068rDlcnl6Ojabk3HWAn6e8rjM6Yx9zmOBYbW6uqBnMvx6r7gBM9N+u8Y
/CICPtPNvSYkckQRGN57K7yA4df0hvBgm/Yc3YgU+zWpVBYn/iMV/EPVjB/AB5eP
795fJugevkx3bx3EFCJ5rhuR9QJmlOEZcJGU0/mfXWhqDnbqOS0V8P1IMtO3rrpm
+lENKStyUtVLRJx3D9R88ZPFFJ3f4bv6eIsNdYhLZadNVoY5PdPdIvTBuC85wC1W
EMyIY6koaas8pqtLF+fAnmMM9EHyobJNQ7U6oCwlIT4hnSl8coJLK5rW3zEy7VIQ
5WCZE478sWQdfR16n3Frw1LvfznJZI6eAmfsGmIlaaVb1DEU6RDC7CBpXogCOKVd
fQusWAPYtP6p6HpY7x8UlLumrZ/NH7EME5fUGE1Y9Qw0W15vDtf0dxNIX9Oh8YBz
MmRghJQ2KDKaa76HmieVrQp65VLa0IQupyst2UHInofCUbffjJaegL58Uiza5aMt
FXA+A/U02Jycx0xo+1+Oo07ziUDr41tGvGVMnv+GvgwnTcVQ4HiB8V0X+DzO5+Vm
EVVqw/G1j1gspYvxK9etv82gCoxKjis7urbf/Lo+bWDxDtWb09/jX+gWX1d3svVl
TMI0EFSu2wVkHFVb3CevvkxmGb3jnQJf/HSVuxm/GuEOVvFzgGmi53LDGvFNlzyq
TPjyiLtF9SLf9NMOcc28ZvxHST/rK1c+ZR+P/1YNNLgYkFSzFgtpsgmlhPAV4UTB
DzQ+uVmWYTMhMNkBWFtXXBNSotjehDGothksJHa+Jgr9j8aKjrZcWCE91wpKVt9E
L2yQeEBwZjLv9+bvqYUmjSImtrOo1no/r9ZxwL0Ya+pdUkGpjGtK6XivoofdTrUm
QB2wetovcGbrGjMejo8Gh5l2ACqih93nREfUo/daFMuGyDuYtJivZv1r5rPXQPHc
p8GIDFmGleufKGFQ6mz8F3koyxjgZ771v6XZ/yrbF8RIfys7JIS4h6/enBZAFir7
Jv6NvK8DdNf/5rtP/xRRh6mRrIWSG5INdf+AnszfsLQGsKwoFHztANJWWUO1giBR
vrAaWi+If2/p+91CBe6IzecNTUfJ8lrke4Igu3wWNN6SeA0a9u33xE5y9t3f3yvK
k+46sJEWLYT0KsDxGUH+zIn1YwIduIiOX4zase55d8DzlMLA/PcTepprHAke8Rg5
mRRZXeJIkLVXXXrXlrPCn9atAKNsPZnKLVg7/POEjRJM3661TK+yMB/bBsH5Yior
MSE1bKeFWH/tUdVuYgQzVC+kyYAa19CPr7IULdGFg0uxVaEyi8f//BTCFx4s9c5y
+79Z13iZAppuyZ0EDraIGHuk1TIdNN6NNvrJIbtuQST4EhxzHYGMFPd0XYu/fTeI
LRbLNrAtdB17BffsawhaxUyMkZt/njTpcrc3XlVkJDQZB/V4qR7z9S8NXAlJ+cYl
Km0HsPNrHbEQ7tzTVkdcqnwALiTZq3dpFnqFq+2FHGmp0RYJAsyEt1mtqQvhxKwB
pa2siaGKwJexTsxNBLXj+YT+p11gdBDDIzC+MRJFZ53CQUtcyYPVaXBSLtIxWKxY
IrrUTbIrLkqlRPoaIyPYc+JmkL4MixNAhYjosUlKTN9GMtmY+4yKayzmAescZLjN
Yy0h/ae678MrFDys7e0nW6UF1MH4wjDFKggbdPPNI2DOka18IkHsEXOJ3tQ/xGZY
tRmKBU/KSVkGMbAyizbfEt0YXlQ+8vEB3SaeVKPmZ2arXNzoLmfJDs+cc2yIo2fY
RCPdfvZuSpDgiDybIQlngZ/ZYGMXxCqIge3kdxZ8UXk3HH7wUqgMzxzZF/8u0YzF
AszdohcFAwijKf4B2txey0UyQoNEujFu519IvzZ0prH9E9evs9b2wUsfCEUQkX0w
fbmBdSXZYbw1ZleLfFtlYVWhaXlzPDabBUH64b0CxmOySBK35O2BtwF9nwJm3Q3f
X7N95PLX4Y/8bvzFHQ4adFhm7gZTtNfRt76RUAv7wdVOS3fQNLg6SrwhVRWV6VQr
9fFEph7COcEG3NG6tSltJXaKQBhkC8xp9fGFaGebjtlzKkJx6yvA88qo/xvB3oiH
Roz/w5Dr+yIandq9WOrK4/dIr1YyAYExC7F+ba4n/YaKWdodWHJd31cB2L/zDbAr
/60xCosaNilmNounLSpiBZZtoHnPLtqubBvfDMqRvyLS47tPtEO+hkfHj30BZp/F
nAOCng+Szc+S3JMaw7eyvF3i3F7UXFHh9evyERiOkryu57QWP+7Wx42Wgwnx19vh
lPR+XG3fu2XV2Y9tUBQ6Zti9Rky+1ehbj2pRXk2UGi/jh5w5ztrlhzR+oa1fqHh8
8WRnZzZZ8akjvioAXQza0yD0I1huWVbA4PQQbjUAfBWGQ8yzG0CJPAo2JFgfeMsR
BYxLtIobWbaOxSIMT9Ilbwsxet8taLh7UmDPJ+/Ns50X4+a98wRD1r6VMfXmPNj1
/gHExP/QQGp7cs5KwNB3Tj7PAf9LwBAXXFjK1PNg6ve2Czw0WkJfKVxVGeK96Nhj
H6IitrtA2tCRc7pWM07+YlyX2RoCa9bbKsN6VQI5BRT+yRvzsO4G4o+n26VWJCBq
7NZLVhoRqFNSqRz/gk55N5It2HYHKO8drjcNfABImZC2P394z3gE8tIzmjtRGkXy
a9nxSzCkVwc3TezpIDVBB7fxBcEuKRr8Rdi3WLg4uXY4bqGxDQnJbeLKQTwG7UCQ
0Dij24zcmGzEUdKbcqic1NoiaCt9Ucd8srjUOs5Gf/vbGvHTA2vElI6+VAlF2WNl
Qn23lM19YvejV/dMX3HjqdEcYSxjp+LXYtiV7KvukYUzmP10zyIr45bcK8t5oRPt
/jhh3xqvb4PMooFdV7azmkIVVjuFctsdRkEAnk4ad023xTO970pfNJ2A5h5CXpB9
IRFrpiSMBq1nSn31Jjz4HAb4WgNBRUJZs5to75OXtqpLi4EXTNsBoxZg9Nwh7qIm
izu9tfgAij6ePs2bDNzlCrIf5nVu9whJ/MB4G26xsKuez+SEswAL5C2TuH2ppMEx
3k/kEAtNuJoY3tLGlWFCeEzxLI9ClMuwncB5yuTZa5cwa1box3aDMoXGJg4NRiaw
EmegERcoD5JWrMT+KQEU6/3p3qeMYCJUcpVRXOmfYgdYl5BbSAdcBVjgs7HjJ/Zo
q9dgE5lZrKUnKLnlgDWuPKwsIV2S3IWjEa0KS0jjFPdVWJ+Es3hHnHffBjfdc/Kt
EVulp8+1prqzGUv1x5SLJ9uqJq8UCT1SF67/nWuf6jDyTfl17fH86Kv20gzlqt3p
JZKJd0hFGMqU5LyBW0EXmduD+84LaiupmGtIiSEwDJuHYi79njEGlAcGgterYwlc
ymneWqq4JvmeDTRwvbd+wEFWuBrZp+WeId0TU/CvDNrjyD7MhBXuyrRVf9Pk6hFQ
dCedgTDGUeOfDuMHtxssS70nEME4UO/qDszpNI1akI+moIJrErWxjYJJb5hxixak
ZyXBm8Fv17ziFuseDdaAAse+Yxv0Yv6tEZYTasDWiqC20Lm9++mVWeO7JCIK+DZ4
enXuNov8f69Qm5DHE5L0QcrRa7iL6U2HDgyFs3GUV7VfHKvdmtDH+go7w5IJT43D
wLLhlQoBMbjvVSdvH7wY8ZNkRxLpv7AZNm5EexYwOrh6VqJOVy2++NCnNaoeEkqt
Zzk0kDEIlYo2oZhuguylm8/Aw9qRkXvYdfbhRg+S6ttZQoAQSBIlUbSmMhgTYUo5
I7tb+di1GqKRpliR0UJeA1Vf9AVC3QFuWEEjnuZ7QR2tNCPH6sambFqC+mMSZ4oR
ROBxhT1IeIEKda/vOhCTlyp0yBVnaE6WpgBzvSc3mItu2lPJDZ4XqHGxvKQNpDYi
ZYmbUEgciqGt2m0VHYE2W1w9QBrB44Zjau+qMVi0MUKs/2fnXubZlqLU3mvG96OO
KpFvUtsMBrPCBMnuxx2reZojEvhqQijJvFOrt/YNsBZsdwoXIbdIeNAx8PHQsV+h
Y8+SoSAhE9s4wBya3EqNgX6PGd2Gw5+l7hwZLoobAmF9Ra1mBCDQ7ZabWIw8QeIQ
HkZcdEu1WN/EO0lM1MVdAtH47heioR6UClQIduT3trmuUdFWAxHBaodV+jThHYxs
EsbbAZPwSUcTBe+Zp01xE5FVsWRsiFD++9ShmPqy7jIr4kkquqLIWPlCvWCztGIG
S8ElaGgByYtr2bCGA4Tu7NWnHjORTozEiksZClUgxlceemW6sy6hwGWiVbUfBKEJ
8nL6v+gVo6Zdwa40PvXFz81ZMI+N+yBn3nM5Tn8fS9aAsga+9efi6zSAdRSMrTJc
8TLEding2heOYFbNDpwTIqi8FN4wnkJ2yMn5q9SuFK+AAu+po9L7sYTTgft9s4j5
cedm/fuhpcJQfmdXSbPmjsG8/EwDUhI0lzG4faO10+6yuuMPkvXS9jGKG+DLLrzd
dBcLHJ6lqMPSW92CZLIGn6MzlE66ABMay4beMycPNQrt5hhjYXJPr8v4rQu+qz40
SFNJtN3URe/6BbpoNmwN8rgJWr6DzAAaRASzG73WZr7XuCDI+c+yhSlMWcbjdOrh
aoz52+fgErl2hBMr9EdSsVS+LC4d67OnGLfZRll+IcxyX1kjmLJmbW90WZX3w4Gb
+4y4DYJ7owwk4a+E/3477szYFmMNw2j3AADQSZM9EVnxu1pe7W32ObYg9r8yuIYc
dmOv9PuQ12SQUXiW4KTJWjS7pXgZhui6AxI7x5QZK1Dw0m2gxgUd2tR0udkAtUlR
lxTSU7Dk48j5jCZiFgyT0BVEkZLzE4h6pfNHJfEHU67BkdCpWqKHOXFm03VYTe6i
K9HpO5V30ZYCaXa2PysMLaI0Q8aIeMmUT9/bDms5oH7FP1GbJiLyDtsqCjR+4LHC
YNdaCwyU16dFXCPQCoMfQCjt8tzYGZXO9jysD5N1QEapSLN0jvzpXXZnIXtAxBY9
i7mBvzg2tSdmwiythXTy8wN6nLuoyRWwns9U4wIbhDAd3MNOa8MEvk0a8lwvKXXN
BNiYGdXo8WKWqMGnL0SYDAyE7g99J09fMgPfpYAgVsdd6I3x4T+eh2gSXNwpOIe9
B3o9GWaa/6dD8Q17QaxGUpZFPCvcvrrGmCZJszzeN5Ep3IKMvFIAyG6VoJQoL3Xw
4xwFDKtuQyytDAsEyxRv4QwpaWzyJ/1uX01u5U7O9ZdP9i+/n+NNsyh442VNgH2B
iWxG1QwHHs1NdfwuinEa9xbDLOsfVparr9kTptTnQwH9iGNhdwZsYn0V2hppA7zG
tjJemiusZzhjOpCEPADpCmAqhqFwnrZJQ1y+IQ1iDBVTYNT79VbwQSodYcMhsHD4
cFQbBaPVuTX3FtpMcogRMGthfs42wNsvpL8QtGe/Vja4oOoXjYXF9zSdt9aG7oLl
weBagc1jKICSsq1MjQSAbymvzSNudbNedRjd6NKLF2qbQRNVM8XWgpId10Y8Y/vb
LaoqQFOgPe+ZBGNxrz9NkcCCjDUz4rYExjF93bLpfDlxUrPs7UPAKI9Q+6zLrgsR
dIqG9nGzU5KIZY7NDZx2t5SBc3xBwAw14RBAdHjOEYAX6JZlcp4FyEpjjTYw2hq7
I0x+xoz1kqxHBLna2xIEs/gLeGh1hrr0vw6/OjqYUjZZjAmXJPrK15TIQ9kCGsEq
R9dnYaRR3A3ljtA8Dj7WAo2KTen7hSbQgvZB74ELcM7hFTXfjxC429/V7ICdvNSN
Lwv2+xWiVzzlzE19VfMvYNqmDHbIiyOtwXNv89H0eX3aQiuz3cAXwogQ/M1q1Kar
f4gMYqeis02SxRBYxXkmVCEA8wmUlnQ1RuimTw9jEX9/ExNjRT/p7Ym/oWmrGN7F
u08plvnwk/fIxgwLBXdPecqMYO5q2h5d1x3+phdkpoeHVV6htWo1Q5vj9svRZ/nd
iU/zpTWOdmxBzURVl/58ERtf0xXiw+9foC3xnJWgcUQ1Hmhvh1x8h0v/eJ5kSkl0
+d36WxjSTS2bjypn2lXAWWIR8+5YB6fC+hwEZJ/1t1Qz25Wax9WwVCp00a7bZkDX
H4yrUMQkjjshI1om7XpOztuiFxSgQCWaAd0NwnG26nzM0zsjEy+ZATW9t1HLA/dY
HuTqjcImWBsE43g4pVGjJXK1pFm1zZWJ/Q3lnzOWdXdlxJEksODwKr94ktXEpIkX
t6XvdgFMlllTkxKorlXxzsJLEmsTbxREht9/Q9ksXPim11biEyV0ZhHWW7mVzXqW
7xMsFeL7g9fJ3RaxXl0suvR0Wi2cUyh3N+FM9sJM2EMYBfABmfxMqLU7UFNj0pWQ
12PTv4OpiFNfMvzGo6x6lb+rc5u+43rC2RIV2DfbvFA9bGZJL2NtB3npXIc2Cnxf
K3Z4ZecTC9LZUTOqeb9U0TOZZc5sTvC41G7UqQA/HmEU43puWajc+T5g0Avpwu2T
7Giii6//G3rm1EU+miQlhXcIulekOy5SjKsWWmzVh8ZbbSQT8JcNEmzmfHgwf8hN
5ncxE57IkTeo4ZTVudjKMyog1D37s7hJtxx8dQ8utrzm5WpieaGodhITD077bwNk
DKLI/zNeWqa9jYRKmANbuGPcfFSDSgA4GGP4Y5PO1g4ipFI8JqVOCFEA3x95CwVc
TTlYss0CKwNsqsesjs8gn9OJhbeyF20/89sifQjmo/w6YJAbMXgjeoCGVMsUReA9
5gV+8svCvHMsdAz+rEaWjB6Lf0LFPTEgGIugrQ105MG+B9LfxIdd29yHQnnh34zt
WwSA3xBoUuCHFNswL1eei8RuIG8pdLCEetpiB9TEOybDY7tusjnt+nzAjqvzqRiV
ui+geONwt+93/RL8iXqfsKWREQtE6Ny7cCzP2Sw2BZvV3hHCj1Tngg4KlWZ6pxPe
Or/Ytpu8NevrqyxiJgQfa0rFV/ruzl5FPbRy93zl7i4hSCp9Wjd0TZNiFn1iiSLA
cRbx5IW5W4EKTtzuZIxdRJSeK0HVt3C4qM+aQDCOEkbPzQ4Ozbg1wHF+pesU76u7
7oaOScyBYYWa+hhB64FPp0DOPyYqKuf4gzg7dIW7y5ENDnxnINazylaaBEtjNbqC
04IxtHiNtdG5HQDJzaRBQBip+OdqP1LPt44IPQVuk7j9euZrMBliGdvauQWCEu4k
fidgDcRRRBGlDJrHfopiots9LDmQG3D1dQohjLwTynfxh1wxHzIBd/PLwAnAtix8
zSY5XbUboIFJH/dAcFa/O4oxidZnw6Oi6VnFahpYJW7kpohH05sd47tomV8G951f
rW/noC9bcHNqiMioGYLFwFKPxsiIMHy7tBRyHmTM/kXctBa0rn445vAlm6pI/WGr
VhLWK9f/CZVkGN2/8F2HM1HsdhoBFdDGI70nzfyaGuuiZ3D1pVf74A9C39WC70wK
+2O77Bpx0hTIL45BV/tTCTG/nxPzUIKAt2mgod3/VG3MBf+Nrr37rWKYJPUebR9E
rReq8MAlytSd6KeMuFFjCV4qaGxEpmBEAxmVXLEYeKc5D/e3hR/NF2ZWn9C0iFUM
mS4HhpqLKnw0zNj2nxpKpiD9Jk/JQJg97vAsUjldoF8Iiq/l2xmjTuQoXkyjpoI1
zmwGwH7Wb+toWm/rueQ0u0yfEDbrV8W6LP6BpQyHWLdwfJMQnYfIXTolnjqe7D/v
ZljdpFST4J1Z8T980Hac6gvVF6hclRHZWp7a1LwAa89Agvlq9fGlqQKY59tK9sii
joRAORNixTOjzNHAb2MwAQ1lh9DZR9xy7aIxB47ppFfThhH9fT39LDGtFXKkQEza
EPi+x5J8DDJcfYqX8lURh9u3T29Nskof54vrUXhA2a/oUoPXOPbx8QnLRs8FZ2ZY
eN8O0HOog3tUPFeIMp3P1BFIOTjoGrvE3aHRYMxQ3Yns/RLQsN+oUhJqsOhYh3DJ
Ikb9Wxu2mO1jWKLBUzG5t1uNGGbfrio3zndH1ag+dZdIlyguKYzFsr4xbhzLOl3/
GPyR7VtgkG7h5MJ58i4s+qC8ASxyFmL+kIU97LJa4eQi8GqYTZ07cubuIq03jP77
QehBfVazQJsNv1jlfHiy0GMSZPvtbsu+6n1wJdXyAHDF3s0TNpvJM2ivO+oBBQx3
Sa1SJRIAfka7QLkOzwMDxvq18vBh4S5FG0Ztg0KnmLt+ctyeQHLxBH3d4NYRuIBL
p0Z3iK/rVrJBxpgdnlfRm3Yii8obKY8pdemjYhZCW/0jGiDNAvKgXjx3GYhiqKhk
x41d2UPocRlx839iC9MkFztN5etLi5IwySPoWvBMNbDEgSB+qYmX6huHor7Vjeqq
DrI3449HiOEkwAh5bLk5L2mn/3PBWI77I0/OgYmq/YjVi/LI2tc77OfVxI4lVO37
phbsSfsPuPsglEJ29rQLzQc2GVgykcbINI7vbY/ZR0yw21b+zcDe60vT17LDIShI
zQQS0iCogRKPpJWGn5E/Pdj+Pq8IXaR4zhhAG7ZbqnVhCS8jB3pyx8zYqK6rmcFg
OPtnOnQyStBn7OCCTcbXxPP6LfomHR7lUOhNWkJy2XjJbCiJPeCtzaI90qsJ8CnK
RzBFmpX6nvyTq4D8MCpJKxed9R0Jk23J2A7TF8BBCeI5M7BFKXfaIv7kreRA8/kj
`pragma protect end_protected
