// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:39:11 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
NTl13OS9pdrDbGq7pvfYZ5qRlfWiP84nzOikkLS/iYDcwegrn5646gKi2nw0zssB
loN1YwjOw1wh0ImIPv2ZmMZS++7aquCmX8yfGF+V1NNvyciAY78HQkrfhKI0QywD
KPBAEYYsGCgld7YKF9L8lHWjFJfO7+c6Y0X2vioD5TA=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 4464)
zLr+3TFK2fw+qo2DTPtZurXQVZepKgzYYxh8DdEO/LfnS0LkWVIU3u0IaGIdzPHo
TBLjjeMB35FXhIOlnD2pJqoCee7n1I6n0XQg6+MFUm55IxOzGCB/TW9TnARoMox1
R8eDl/vrWBbuu1eozWf2doKTmuP5n5uNjo8rZX4wZKeLfErxR5J+M/91twxHc8P2
NaJLNFgGBGnAv4LuNpghjFlBhH4RL5SnZtUWooGa2RNxcTb+nMMdiiHclOg+oioo
J65oDwEMYTQbE76t33WbCydWJPR36QipLlYYzBUQxxW9h7H0tos6IuNwdUrdtLdb
hiXb7Z831hvY0D6g65ma9+wzkFRZz0XE9KCSougAB0Tc0dKmbCAYWgrPoCqw7/KP
1bAh0oLM3BwVaU+IsA9G/uLVaUJ9XQ8cVbSJi0/CGoucSCn1h2xaqJwFb31LJ1gL
FhmTg14Z0kkvk9TRQHgEqoUtPnLElHEsrW/7Hgj9hS33mKKIviktYXw/v/+XpCnY
MAp/pyElcR1pl8zbOMvrmmBGepsVQmcjppZY6ctSR5IH/F4NjZry1xH+dBe2js52
89MoAbzf18bvp8dDhv3D65UalGGRBzbZY6bsvmob/GtJIQSTbLNMrxIDvE5GiT1x
McB4amRUxVkB9SfGkPnkrvbIUZ+es9ZJOkYUL0tzJdbZ0Eq+joj7xmqZwez/l4Yq
1SbJEZJaWkKOJU+tpkza1GwfRisMLppYutG7VSZQuUN9D5lzJll1tL8G96rFB9HY
VlSPuvUc92QhMXeKbdma74evM8S3fVCv+c/lQQx/ByWJBd2ctDEYsUM8nHLSiYSy
LUjSVfnReZnK5cXyz5CQ9o4koKppqTK7PahmuK9R9jW1Oz93IIhStmNFcEtuTlyu
ctmE+fWu2JaPFsuJv3wj7iQRdTqC5tCqk8CQ2e6C3im88L6M7QhJ7A+Uqi1u8eQv
uniUWHsGSUwdtSx7iCtNybfLot/2KoBbpiDvACCs4od/O8xX9mNkiabwSBu02NIP
VpUP/e095h6E7cpQsrnutPKh1h4Wlw0VDundfrz+TcZ8w3xLiunUBjKs1ygcvqTD
kXyhWoukxfjg4DHOH+uspWcsQpGurqVKkh9kEOibFhICs3XQTrkkMbGhxoXUbSMK
h94z434EPuLK8DWPs/sD/DeXHvG+1oPoAnsTvFM3lhI905iR8T4/cFHJYASZ01aQ
WEWkWAkkX2W4SO/8d8EPFcjYJJIlTDU7s4yAqoGpr5mLu+8iaUVMsCdxidrmCopN
388OMDKzf2dM6glfzpR/QGBcbn+a0hdUb+JMHGxRPg9gdacdjekXp9oW8iqQIFx3
Xgb7MdVCQ1jOh+uiesF5LInu0m8PnA7tYUvnghPvq+o+5F8nreg/fbad7Yt6XBxt
G+zM2qiObJMQusfce2Lv20EXmh0WMtsm3B7Bpx90QSkM/u1um6sz0nSFqA55KkKn
6uUnxEOBA86fDVhouh4R3I10K7/Gh4gyxYmQjKaniM4RSs3ckGehkl2CGMPBf12c
E8NEczG4RMJBIqmCduacxN19Tb+9jnyP5+qMLYwOgW5+rxwgDS7Z+Gzh7OqLlUJG
KRw7KQGOo87CBpXo/eHSW5lXuus0+9gG0eONP+dF053PFEgD7W+R6h9qSy09nDQH
vdnkj93UPozfaaK/IzRyMlg/Z8jI/QJ0GhG3sc9wlLsgMKeaCXMydomSlJze0i+W
BUD+jh9L+PSgy/nT+tBe2r7tgDjFhO+93Iro7RyJNryKSp3Ldr2JqmSf8pTG1bP3
Rrt3NU7zgBBL8+FHN/P+Bh7bZiltB1X5eopwzHpFcgI/wfsbxUZhg01DJ08rCwa2
sujYJeEavQQdklFUr2ANirbdMmZSr8ePe4AAsX/VK98kXdMdJJ+0uLEVdwjlHcxD
imVJZKROx8zffcsYcMWVPSEGTs38mnjnVxaRjukjT1ff7JiHVhHXxFxtW/z/7mA+
GFnijFZdWuMNv1yyDDCYXNq1D4g9ryZeR2cm3vqDZklDL0cWfwYnzriSWcINvbSw
owrC0pgsqieI0JggvRgKlVnghaF+UCdFHTlaGXUJUDNuPZ8DJH5+u1FCzI+bo7sS
vsb2WkdCjGBskqlkHX/ZKfu2lpx2Uqp5fdudN7DOuugbyI4C8gCpSFWFxkqRcGuA
Rr9BvwhTWj630wbLcbVci7pRdiGYS6xZ3plUmyVdIa5YzISCQP/RxkxV5OjtLU7S
/olOE2AE7kVnkCMTbqGE7xAPQNOf+rOBMS/tbaeZp1RSWP8vvCHtzbQjXzBx7s/0
o94gH5y85G7+cRpRcWlDXxolua1ZIZFfg5r8IcnF120R92rM5aqQxeAmakYwPveM
17D/ZbPjY8FkRx8mGTKxR3iQn5pDhsfKv9gff6l7jVw0bIPnQ9Z9jILJRY9iKLsO
8hy7PF/woj7ukHyMeT7wRLbB5ya7McD6XfuGdw9KcR04mB51e7jOuVvbJh1JW23x
HgdgvSF5xCuu9bKnVMhgM9oslU2naFEUEs6/0du62o1XotY0aPxH52bRmB9yuF/p
ZAB4YkozNqFZzQqd//Zchv5o+Zq7puog8uqVoHunsxa4WO6M8rSlgTKIUqSLE7m3
ap2QTMya6PaRltevNP5ff28PuuuZ3i3aUcakTBaX0mIJg3teguG056Sa6uJJfV40
nAzjC+wttrkpnI6fI+GnIUmRSsGDXUF6tKDQqB4G5oinraZSSvC+RfLwXMt/PjzM
VkHuaa42NDscKDl5EXK1nHWKLYHB89Xdi9zA1AC0msu8pwgVlapJ1DKFDBPjpZzm
IGW6Viu6gN12IOD1d6wmDy8BReqMKE/3ewFkRe81QciOqTRRY9b9gCB95qrcHBAb
BfKA3VZWcg2qoHEmdiNzdsgwqF4F3dVER2/lZu6j8xO1AJTD58SoHG0on9bAhPlG
1WZIDLpeSAlElN0AFBO1Wp31PaGD53oMtMwmD+vyeIrUFe8dKdbQWw/JRvf27HU5
BqzyqSS+ofI1p/YIGg+r8eoczVT3NF4/RXcWNzEfB3mMjnfv4p7FQHcIzevcFp+I
uwrpAiDPzM89R3L0b9jmFrsy3b63pmGo/28AgKzjFcsr6BvopHrRm0/gdnfvslzq
zlvvPRrrkmlJQlw8jMhDdZqK4Jc89pRJUlZHjtCk3B+Kc0omGHWwsRazEQBtvunr
7jqbAcVbXDG+7ioNx9exZl8Hoqzh/rN467Xjhc+Gks5O0gWsK121/IgX6QXzUiPF
zBhf3KPM39R9gaHHMfIIQhVb+8YhAJ+Yj/HonKwIAaXyYQC/PgNecrMDkGjm9Pzp
VX7lmMO0YCyH1RfgitnFLwM3lHlQVADhptcWC5FaXh5pZfZtx9Lg+OZpFdVL+0YC
zDyB0pqQGaswRlP+iPcb2tiM7B7E811cpzl7qYJTW/UhprFuBH2Jtgg+0d3YSZ74
rYsLJWeLfnpqLVBcR7rIDvVntObrjNrq9aa5kch4heEewgwjQhF0d259rLo8g55q
JBvLA7lFAJtLGllZptUswEno9HU75xlwMT8rTUJbxbagPsocIpZYbHEBYqX/W1xt
5v/OaUx8EjNzmzpujHPsavnEffoZkMT5oFB9xTHMllYdAAyvD9RcRJIOOMSszQMv
Ix60cD1t6pStMyLbpV8V0QBF/uBAfJ49fs8x88Udg2jz/OsS4Q95yhsDBTzMxBxB
9f/AB/k0qBOragQ/54EYD6ngTJHoJ/s+lGEam1Cus7jOa7W5VFr2zOnJ8+Ko5Af0
D7z14t6q+iGJNpuN6lQmOjceq9VPcWOFByTGm6WaDQES03GUxUx61IT65CVKChU3
xv6HxnWvuFeFXkZpJRL9BK5OygSZM2kRPlw7YcREcbMN553u9C97P1qHf1T33wPa
p/dfKYWf3q4XurTVVLQS9Mh4SJd5RSoMAPrjSzhM73/kuEwZTG9Q8c27kIYVzfav
T87a/I7/zzxOLFICQzPM8hC0s90gfhD/KM3kjTT8GFATzAl9H3RO8/4gh1KZnLyI
8GgFrqr6EkvH1htfN5nn6wgr/Po1IXwkiK1Jwt3ZmAXUSjqlvYHFLENpYO5JS3ZJ
iQKed7RGqBU7IiIJ8b3q2bry5i3BeTNJNAV1qjxbbiMn2MFs5NNKFKCkfYL1MBYk
yeiSwNFT8vcMRY3njw4OaxYq39rrIo97QjPS26EQmkr0psWPaYMRWkePhCylBom3
Kzv3YGDJTj3LKV4TDduEhq2rd8iy/9Jq6zlKYaoPZsAFUlaUiN2sZhLh8ujrOYXn
hs3ApFL4TzUsUJJ4YBfk/pF424gt70UIaNGCEZNF2zPUGcVKmfzyqtLfgj5WhPCf
MtB+YHpnUys2BXEOACgrhgwxKummHBdTEdov4sW9S0js7rojZXz9YwuT5llpZC2J
02AFzxQrgyxAv1QGx40qFv962KxAd2klbGSfPTAHPT7Fm/fwtztn4S+ZTXn7j2Lf
C4NnJN63adKVZXDSgwak62K4FHr1OVy4q0GIp9bgzh+2AjTybBhngpNCANLrX7vg
pzq8a0VtMfZ5GELNkkfQ5hzQ6U3deIG6VUoUy2oGLH+4KJvh4iUbI7iOQ5SDeSjm
Krizz7v8G6TZOi3HQ/iZSgF+KOAUTrQipiHfzJkeSFGpkeKTUHSJrqCVRKYze5eJ
WkH7r6LLgROy6SdMeio6aos/7gMrw504wUinbug1kaA1uhLTH+E2ehSwUPF//ahe
ECJxHdQVXC//TnbK7rxDmMlIF/LHX2//pj+1jpwCys1CFxFT/tQckCAj48on5kmM
NLPSI/9oTUMwL/G3/2iXpKYtmczXG6QRLLbFWvXqvJIsgB50CQyaBAnu8c66XKJI
Kzr+JCFoHIlySeaZ4H0RJahBN8JO25wx9fO8NhdNFv0ZIBRXbKpnzMeAIQJJTt0p
Gkhdt4XqDiVlXXtGUWyF0mMdrKMdYEpsfuJwKAx+6uRZ7I16qnnX2KHST1e0mDqg
zVl2bINPRV3CD8HjKhMsFZDzaHydODxL4opjapxOoAUjKimwVpvKEMX8f7p1mg85
tnZuejH7XpVoYa6ZluO9AjHUc8tZay1QDtPFgIYnsSoW8QtQ7QB0Pn1ZoMuRvl/r
Q5Flb/Hrh4fJ0knm1CwMDxcmbMK6SyWKSjNNMYwOKIr0GalOZcQrfUtyZeR+d1vL
envlxAxZ22Xjo6A159qhvdujq5G3QfdCQR6NoyXt6nf9UqSZDRE2SOpjjtwC2dCt
a3dXqHvX5/SVblK19fexe+86Kqa2XGawfmBnFtqtwCtp+QwDbrylEBKYs5OP7OTQ
wgsC6LIQctFtUa3QhFjffe7gTEu5jlPJ2/h03zpjyjyHjpXzC1YjPik8k5k4engn
8E6N/2Q5l4EsHMTCvTgNjGvVGOOnCP2wz9q/H2Ervs3pLvUFW07wMeLVd0PRpeYd
g786GfwzS86/w6eOlOej0mU03482fLD9kYEAGF0e8HPcv9iKo6tTZVc0DkDg2T5S
w45fotKejS4Ltq+hK8iqBpVekNEhX+IqWmH++RIWDdAz6p6CGwFpXv/DB+2Dd8jq
m/HjPgmLzoXr7vnWXABxzWjso6Yi4Z7rbizMm86P7qdqJ276itNo6qmJUlI7K/99
nN9E/4QiiTcqtXxtlksY++2yFLhoVGJY+J5kRDVg+RPqvnowi7P/qOcEjlYdXKIb
Fl0BDJLmmW9xuNogscfULXOyoWE4ww4vR0ZN6Oz3Umbd2Qq1UBB5HKNsJQ/f8m74
0fYFst1WLtoBHU4BhzqX6m9Ej5KQ2ZU3rolkCp2K7T/9u4ugoXFXbwTkJ+rvfKnV
nNaE+upqZn8/rRNy+8RQDSXDjJ8CqoaVgxIBv7n7UX6B+PpcbIAazzmjOjyId4uK
oKxew8iEuLnFYWDdqCy9loW/YbJ5f5steUTVsOXHmm/M1djfiro0eIi+xiuSf5Qb
`pragma protect end_protected
