// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:19 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
T3f1UYGafsy3zqDcpnFkbI7u2NMfcUARmliNFz8rpQZ5m3IMvr5FXR3m3A8WZXFk
T7QTQCKocaYpbawJZwbY9Zx0RGs0Tph9lLRDj4jefbnod6Qk7UiIWYOXsR2xw5gP
bLHbfjg4ahK1sks/6b4ECvwVtzdIovdY2tkvF+u8V4o=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 72784)
XsS9Jc0LXsCJvhwm2aTN3unbauhvZ2vOUS3z7E7CPjD36QS1eYEX7P7FMrWd5XOe
ZO8a8sB0gWih45kXb7j5FR8JaZ8XW2N4Bb2/C7vtZwPu6+nhYYbFDO9LqtwxebDG
Zwg7SzkKIltjbjs1cecBUOzjcmVD2hoj/7OWMx5A/rOmBe4257Lrhg8a6ctjVV3O
JPQIozrJ3412FXpVyoHzmDNUV9Y+6+FLD+XZBbwkgHd+P7yVLmHolh0xj7H9mWR+
M1Yhg86Ilxzbev5ITHOek4E/dQzeJGxkBis9X/E3kiPS/ZzvFvQFhUebbsa9w6Ec
DbldX8y+4pjWfNWmUpOkbc2sfawOOGBwVHtvZcPMigY0nIE5yQp19thM9nQEEO+o
zA7ANH+dP6Nhe/H3RUWfgxI8kD23JjcPQA9HbKTao0pdzh37YObdEUQgo/QrgZ+n
xWH5Ik15jviDzBrt6oxSS6h1nweCis6jtEB5xCeE33sjl/BUOjq+dXrSGGb5hhm6
7UBH2jfqE9W8Ea+uMTh8xU8iIOb7j7IoxvmeQ6AgX1u29LPsjAgnmW1Ft45BFP9w
z27v/RZ1tioPpjoJ4GcjhI9o/xJd0AcLd7m2fv6Pf3CwVPUMouKjFxDAITeWaBXr
6Nb+rPY0DgR5/RUc3NL66mhP4IFR9lSMPtSPOMg2bOWzks4+qbAVvUWyYv71kEmV
FG0dGIZYFGhIsWzz4lH7DfwDKKQcq/zHpjh1g1rQaO0H6/4XNaYHOj835cb6LBXO
iIdERhTvHFhFIfcQ0r/l0Bmno6Mt16DoeBLqyiBW62DU6DWB2zHrKedHpvISUdb4
QYRfv8yJujpgakya+idPGs8HY23DZaWzKPFoOocp5/cv9XZNWzwmkhnlqzY9Fbbz
tuNyEI4bNrjYYFlLFGKrs8+iUXMxjLp7kOO8/kYAxMF44SdC5yJt6QZcJ6hW3HUu
2yd3cYQSRckI/CLm0WTkgimf7QF2Vp0v9NNwTc5IE43NV470rlqQrE71RFIoiKI/
74kulgLT59Ij7LrkdU+sN2r50Jzrl6iV3JZCSt9dB6QfJmDe1IXpwhruYVjlBrCX
fDPO5OJPSnJZSoJzgqB/Ah5gTYOXLC+zWGViuCEavA4wsyitTfHNxE9JgFfWRGjm
w3N12i3u6shueXvDuBcZ2PgQfm9ZFBPQOoAti9ZrxOt7/Ai0Cl/6EMKj/1FWW2Q5
UE7obOLQ8qyIV3kmkJjkMWSPwo7T5ih0ltFnuA7EpfXHa/K6ilxztr3Crph5Kn8j
tXJLKw6hazGhKYJhup4DtF+maBTf0DUJd7tgZ/8nOpkWVbAdD5hKHQcPsfOjRsma
/C/jhRvqOFkahIvqYLZF52zbXME0znYCAPTn+JpoWTUF8fti1JbwOL32KzN/OyqV
Vm9m3MCdh+l8ZZoyHc3eT/5LXpeTJy/hjuuXgm1NUPU/QXg7MtRoo+y3QI9CXIvs
QUEFamPOsh29YCX6Qkg8I+JF/T2i17X7XXehexnBqvPI4qhLcwcf3XAq7cIqH58I
Aj0f2yc/rnprjpt+HqW/uiCRdp/J2FbaYOgeVN0ZE7dUVyRQkfPJXXRj/LKFrtyG
jeDa+rhGOUBEheB+TQZmoHZAABR0prmEioI5V3b2WMJRjboVjWw4Tb1JQk0BsJ6h
QYuaBMtwZziG/zYZPTTk30gAGfFSYb5zxDQ9G9tYkQwD5ac6q4CUkbgqaULwcbms
YK5Ay83dyHLP2OxKDVCQ8OeNjo2TXXY2867E/iCXlXLR3Dm4K6D9vl3a+1T6+eIV
1HNsfQvbRr/gSJZ869PM7b6gjGZrGv1bwArXVVOpg73H+WnWgvWIQwlnEJkeW5B8
EdEoqC/VqFPf20WyBzavZ00wrts0WXwKS527z5ZFZcNmYa8m7cO5vJ8hZcqYgaWB
T4Kv9ok/+PVQCH9TXAtZIhUmKKOhj5EJkBIU2BdsgT43uxZ0S4ul+GV9jFGAfUBN
XT4ullDllVIeOEAha61PFMBk9oN4nSVp57FLbmru/HLzqLGJ2110skBffIudoIEF
WeGifRavsfNYC93GlaQAY+9qN4vb1rwP4rgJi/prQyExYZtTTcJWec5tyVcHHgxZ
cVW6pgQtfhUPVRHi7HTeBt4Q5ZYPbSeHxL6kztMUW4Ni6C2nZmJbXQlKVCLEcuyQ
dFTyk+GGPgMmf0khMBS0IYzjrC89L6kdryXL4649nc8bkoT9dCQbnXFsGUSNQ9LC
LiepLu8p1Rzu9qA5UIJIYrLLCXW9MCgOzjfNWPu8HiBFJzv/7dOW7kD5HB0zQcfD
RVJEhNAT6LL9Al/c91nTunNm4R30/I/XtaLFaRyHvBd047CBJ5PK5cO6MF+U+BkN
pClbolCEfwMUWa/qTduLXvZxvMPioR+ngUPLCPpjfcrmXCKs+PXyEyszNtc9wAya
7wZqjsF/ZbpEJr4zTdzOX2T4NWrjABCAgTDoTpWZQGeogEubYirqHrI8lZlPINeq
vyzh0G6rloWBtrv4lQSUjRMjB5q/71pPr3GRYzyUNmSbYtA3PTJfMoq4z8n+sIXd
HJjHj5ffV6vYlaBlwx6qxD33bxZ7rHAXYqz4Yj6TGTDp82Hi//riC8b23WQVuJjG
dYghz13tGjAUWpddc0cgqQm6PLK0LRLGKjwrolSb2wIHyLYbPGvmqTId6JyUDeAy
S7DKYcU4Qc1IRgCWyFOMLstWIOrG9KtyRi3u+CykF4nZvxxvLmTSG3yMUZEmUxoJ
NOkDfa9VhEZiXK4++aF6dF3lxYofDS1fM63Gk/wGH3YArORzbAP4AtLu85IMze7m
QqEJlhjTI+BGr2HEZaRySmhpyMcUm1hND0pKRhr+Uq/zP8wrDsv1MNxYxNXB6mgu
1qJ5RiVzB7iT6nT3GO+OYHpAUlB8KRUIjI6qGUoZkhXduK0tkyJXWUmh8jdTt2VJ
EVlZ0sI15h9fvtZIeO+DjGGZUDTNVteH8p4Ww6+rM2rF5nceLpyidNPNHFBDM7Oc
szaUYeUJfyH7yQsf9OkHMj3UvRJIkU2aJprUbfZW06eruq+QruRUYOyL1/aiNC0R
5UjMmQIldSUG5zUnSw5RqNkydZXC5cSENS0w0OOEBMBYX+nTFNtRUtmf0IQ5xpDb
kze48SFUvWfG0IIwu19qshgkmHgd9rJYihcCEvwhYtS3vP8kNp1kDnf49tfi7DiM
BvK5I6LPHNJyhjHZShtdDreNvQANiiz6Fh5evpy2iXFDEEWeYfw8FRN2ZiewYgcG
W4FYCfsKLVFvT73ZKAKkvdSuYgGoP6CSJZMZ3HASko3Nf7kmGplD3/KhyCSh9FKt
rFu/PLV04cJ5ilYTDbVWRTMh7pR3ffRGV0ujDFvhrtQY5AASyp8iQFpiA9o9aW67
xCsH+QXb+4U2MW8BV1PZuh4hsU5waXEIifUCnhSzJvpFO1fGiEVCCCWK8ThOdpmg
TiZwqroZ1qY73FkMGMTP8JKfNXsCPej1vztfqayzALasyWPCN6fxyOAmgmD8PY6/
Eb+6pijADSBK6HLEd6qb+LWDC5X8jkVcn3GIf86mkKO3vQGiOlL3m4Dtg3v2l8Jf
1Rj4bOfVyRuuYP+S0n8OFV/0AQEtaA6kxTwBM2Z+PyOYPSnZBDmIdIKto2IXzWGn
wmVM9sQV1IouoobEBZ0NmGnjT1omgeiUJ6QVTbaXd+k7rSZKrTaeOgkCF/owTsg5
a7W7xx7Y/q2u0lusk1kJ+uSV0ys0bEudYUlWwBuV7WAox7C1kL7T3kN+VA3JAOgF
w9iRdT7+zlVXfkrFJoUlXr2sO0Qq6bNulWlXQPE5AgoH0oEcg9F/u+TXVDssCkEo
DDyQsf8K+fGhtY3BjG+4i1YnKKrcYwRh5ackJg0ILSan/wkNEfFJtirESrCgrmlG
WfsGQvrIois/eiIJI5MxxUm9qAToTLwoj1ZDmvvxyS6Sm/bcRdsGnUiNDB8X3o3R
9P9/gXltXc/BdZza675zEw4xaHi2NRgBJLF9ov8MLhw/+JWgf53qDrCOnsDVNRJd
Pglg+j9NVXMUdSkQB3JVaIMrs+YBZafPQf+QsJyfI9fVbEI8NsRGt0x0RFI1V/JD
5RKVrBePWDYPBBplU+4hzP68SBJ4KU2KKuFcGS5tjiv3/8RnjiqP4OBOlk9STV9B
erLmCZB/v8sIWnEbhaZ937wgiapM6bK0J5hGXdEl1KHGY9eYiQ/0y7OkOmC6t8Hr
GOpYpEGtzCkTnNgmwBqbK+TYoSd/4VsjZHCiqb0i7GxCP2OUeP/MyB2OQNAtW1wc
kBgN1hMEVbxPeSMguIanjijAZIt6+XqJazNQlg30bXC0f64OSC3M5S36BmZ+f5ZA
Ft84usAdukM2K+hjvptQlFU8AviJAGDf1Vb4oaOFFDp8ma4ghUKsB2g9CLypW6L/
12oPKMBI5pFciUlPN0sNKsdJulSDwkBBiaFAsP4LcDZ8214DhWmaGa9/xwxyC9Uh
JqLYMYGwFCkNNzcf1mf6qNBzI8Oo8QokrB8AQMD4BtbRvsztBPxtbKi1i0EcCnfg
41G9Cx+X5HOzabt1UkjKZ4a2KLbL8JrDaod36q3MyKhgmhsdWBechwMgRfK8Gqew
agibzly4G3UUNLH+5UfgOiBHg1CyKajMAyvGjYnsV25o1yqrbw4utxoiV0/3lI4C
9pcXixNZm8oj4WrE3IWYrSf1wotcSFd87oHNrltzV2JR8ZpxnUdF6N6jWmdDGlAw
CVa2FvD4ho3Tesv3tz/uXV8NOqC0hyI153soMHcMWZf/q5n9HZAhPNPbmXXO4E29
2RY/B3CwR/c9bfGF/PkrrbvJ4dQ/w0vsUFc3cLTocIu+lDdUs3cdVOS973HXNC/1
Bqd5MbCQ2u0yERAM927KawhcrXp1q2CTfD3l8ZE6KKlrFlaK2cUHIcIEU85pMxo+
8ufAUC7EOqOcQcgFXoukz7i2Yolv9pBPodjeb1iuFLVzUjwhrOruVL8+6tcZ+FHI
+ODgKv0TKV6AX2JdensR5HMuzTuM0aybZgC+OZo8EqhVuH+p44gurLT2AsP1ao3s
aLj1fDAUJjkrUl1oQL2VTabUJFbmayccHEjO5qLhUjAyI0gKO1Jsr3sIPxptL2iS
yzWor6wLLpEseSay8mVJqefHeP7n+kd0KCtDoWLdvfEfzF96/yVyMZVXKCCQwrSa
10bcKlDciJRGSvxOxq0SyJp3/f1PEUDvLu9zcOLjawzhTgeoERjdAJS50GNmCzej
ZIyArx9CquaecfPNxY+qjQ+hELAtLJyfJOXi5ZFi6qTcEglmv+aw08yhNuo/QbX9
DuIhtlHebOla0hAnrx/iFxyYTC9BT4EORHMjsFEflK/Bc2nVOqDoCULgx9EXGeCW
/VczM0UPWEBizwphAHNwOvR991hkGKSZt+6h9CVJTsTpDGIFc+6Bo3S3PwXWCEWN
Tg7JE6JqSk5Fw5wBzWcZfLep4H28c1E40Hs948Gw/yyy1uqfkbgaWBDb+ZabkWWb
lqBFtio+0JB9k+qctr15hRajwOF1i7blDP8gPxi16B1Ia3LYoGPPAQq54BtNEUF+
rTFJliqLaA+lX/FfH2xrCPXZj0pLDK3+j+lMgifyvVcFTkFjzlWizxqp7ng8Dw0g
iWXD8mINjumLCr2Jut3I6nzc8Un0pCTsozTmobGho/bnIop/5hgGktUbBaLyPvHB
Ltwsvqwy7gg2UEBfROZXtQLsX1P6oOY3ulLW5GLvbSxE+e9+nOR5WBytSrYvHyVW
uCKxrgKapo7TzDiknGBxGQ/NWU5pPVm1sAXLFAWoGuYIgTH7Ta56MYNIzhQDi5P3
yuipvZv+x/D8hHln3b0Dt6CU9vjiNfFmXp/j5R5raFNyeYMJ9xEh5bxggg+x8KE3
8iFAMP/56KLoJ/nKm1/rCcKVGK1F9QYq8J070d79goBSSBXTzFrhEeK7kAogYiuQ
1K6ZwpGFOiE1aHpm6cithF7Xy0/5edYyXQdoKIFtQMRLZWVo0qketJ7dxKGkVR7S
2R6LLbr0dOaKMo+kYF8q/NryKQUSyjiq35Q+Bd+vIpxAcCgI70jlO/7jMnXC7GmT
XjqawYxV3QchVNR+wQdreCkiqIjH/it4+LZ/Zs6xIN0sKnLZr4rFPuEiHqWmeH8G
KDkrtJXNRM3ncvov1nRToX2IXMCWeP81/Fw9Lg1EkCvuFhHVrgmMaY9kN9A/v+1v
7EVyFNUvyh4iKHCaJiCfXTKemqAE3WA2/VFHDMAB9BJTU841AoCegn1ilUo/hwRP
PcKE1ZOo6ehM5h5JHzp7PJtOphqFvx/gjMQroZ6vAicukSzACMlS4XIL74KuOtv0
rRKs4En4wDkrVT6nuc9prOJAF/toJ2pxm6htf4ihVqNxSf/PY8b0jW1wrJ6Yvurf
1UA5q9RbTgTjdjGEn3c+Jukq+eRRkMGjrtoxQesSbDDIzfw5vxXxkB9McZ/I7qg4
y7xCsWC8CH2fkpYQy14+HEJEmd1tTa2nLYlRtxoS3RABxGPCEjQUWh7pQG1GqWOd
6koyBD7vIVpWAySagwyh7DdV3/ppJ+8oEjmNGiQ/CohlUK4LKOHPKwpxMpkUVWQ/
q7wfZRi42qaN5dafy+NAUkftSSoQDqXqGViavzMDg5MGDqk5mbqU7jRkslVOU8CE
oDQwSnGvviZC0IIwuY1E9TKzh10SmqWjPKttTfcW6d6ozsIdOjra7VsKhtTuPkvt
ReiYqMxwRAFqxCCSpt0KEGITz0MbzyV9K9W7Ou67t0FkwzG5R0XQiFfXZ1AAq9J7
EA6FERXYipn5/vldYAmmC+RCKGcsDLJDzkkKguc9ZaOxPanUuyARMObhisiwhX0j
ni++X4J4G28UqL4O2iJ+hochpxzgvx3oIzhVcGEW55HLnW9E7vhXRpiToTWys2KO
EXAXbwJcoSZggQaqDT45XF5G6cY+oPYPzmuDM5tngR9jnNa/fMLDTG9GjNMJ6Re9
FJjxtlAF9bLGbm498zXdMCSMa0Nd9emnUrpFID37oV8Ut0uZSFaot0WWTJPLd8Ci
CAjPaYaVW0nUHirdBEalPppP2dbYBkkodlknk61HSiwSn34u4NNhbnUJUDe+3Zjh
cs/WAFxyEhY47reiUGaeAdE0A+w/Fg9U/p47wlCc/uZJW99y+xkuT4mvWRknm0Fq
gTk3lIOCec2JSlS2+Ld3jdS9ltG108656bqn0qKmZslD4RBEm4keMTTUqSemNsz1
KnJd0sj9O+0x6yb0LY/ZkQpHs52Jp3eJ7Ho/gr25zY+ek9wo24fTj+/bcThVYrxm
nwH6qZqVlVAkJrOBEj0jrbzlySUtf/Y7h6wSX3P9mEdyXWGfcZRhaVHFf/XiifZ3
Gnxi1tkBSNnPowHxGn1vYX6sKMLWIk0XEViqZx3kl4Vs/9xbhRb4iQ+ubN1ZycIz
YRLLbHXvMMhd7dhyfIDdcB2P55dx+zYPEBruridSZmkrdomOvXfGS4lRsHWfvxjL
lNbgQwyyrVHf7wPeblNR9ElPbd13GorjZNZjHnQqDkRou3OJU8Ky6cqllouLD1yV
93W70lntzq40i1tI2569xsORJ8eC60ijUhjP3B+XumpvbvP4AW1vDEcIH6JIhBFs
tbBgGLxEe1wXNhb5vvuxZYUBuW3p4h3hyXz2f4npIMI+MswACQdy5tpQ3Da1YuDv
ayWqpcgDroUGir14gzM0wnsTuwMw52L3zaZmmBgEdRa7vUryxw6BTz1SlbrUzB2c
V3Ju+ZD/H1YvS2EdWGKjfwxvj/7+0tcnhJ5SpByK5OqdRFROXqBxPo/kHK9QbsVb
MXVU7XhfWoNksXhrtytWPNVCWTb0A38EITaTC/IjYwt7Rmwhl7Rg3IJekHsPlkXK
PY3ARTrWiZ6Id3W+MaMQYav5RKT4jvFEj7MRuCZeURCP5aILit91ieY8Fs08HtTo
FGDuKwJOkcydrS0dHpDYFit/ugqGbV4MqoBGP9v5zuGv4NP2FnErtDyRF9NrCIvR
BWncEdyrRkvWRhaKR5nHTZWmNvZGm++wlPZrjwgtMd91+tGjtOjaXpY8sFhjhX4i
c5t4ULyyUpUrHbuHOVRrtB4dC9iSkxQu0Q7/AcZ7mehG+ecdal0AAuV9zpppH2cD
2cEJR/irx0Vj/hgoTVBvoIjq/6t6mk5GgMGYaVqJQqkmtGm9SaA+MhbrMRk2HVkW
tleeNAqAxjSPYJBCZG3grW8UtZdvLhjqNEDWAsqvJJs1KrO1QsRAyMNCOv1wHJ56
mFLoVjyFGapvvxex632yA6kWiHTzQ50V4JdDg/8zOKSSCjiKlVGRjHA/7cLgjp50
Ua0vPJqYzxdm5u/QxQ2OGzbVPYCsU30J/akYREYsHhue5alwGQioWinhE5VNT1eW
s5Q+AG91P/SCXfMNwdanExGu7HjDlBN9rxZw+uU1XQvajmMnVa3pDkgactOWeo95
5le3xxIILReSfgXbLyFgEtPCk836DI9N+5laYv0MLr/zk54UvR/v8iU/woPt6Cxi
jlvSWaOm+8wbSZkuHdyKETST0II4FUF7SfM8BHOjqvRIC0BTWQNrUVFxIdfq7IaQ
2lUgekG0h87oIkxPdaZtfBJNhDlVA0bvJDbAk4AhyPL2yH2PUwEK6hvOEon4Yzij
JeVPdzxECmXVDdwDoZRoc04Y7q4TpObvs019ZzVjnSZDbes6k5KgFDHhpPghcCus
uuPr6Q/JIU1rdazk49VhINz23RQsRRp04oZEeRijyA1tjERRri3cY/TwqengkKkI
fnQrnq+iHjOB8CCF4Muk+h6N1Qp6JxDaythhed3Ivdp8yxX9FsPG32cOYQ4e9tiu
2iqL630ShLLrZbyG6m6A4XosVlGAXycHJ4J8Cvo5jrjZne7d+kn1/5bjWrfTvy3h
+1PPRHrmQcw9w2Zse7c6XXS+otWAqiduazo2qBrqoxEQWk+go3P1700RiSsjR27S
PP570dO/qRfZuqLtrvST33MefzJ4OimBD3b0ZNdwxdIIcoJqYabIysAAfk5kcXQo
LLPeizGJsfHkm/XXqWi7YZgKS7iDNjLpwzEQafm2SMdjW4KX5YWAshQtUmBGk2Cx
jzsj2tU6bvn6rbCFvIrbISncwJfW3MUOkEl3Ot9iPHd/MLu+4dH9yIHlV3RIkR0a
ZMphMfsGsEkYjGxkbnHnl9x0R3Dvq8UQN4xoskLdnqqloNWkXkcocxVyI0SMPmLf
FtkCXeG0HjMXRYChAAfvnmQQeokyZcpYJ0zHIyiNddDQ2L5BEiyd5KW/Hs4AM0bA
4bJWcRBL9msYSLFeDKkocDgmahpRIBImwBXemq3sHFLKbhnxkpc0SrTYElxL6qLx
vXo6+kZJsjbzi2Lg+UdJUvyGasrUwNGckaiSfDXwEGTv+BAGUk1GgcEyeVPJv+U0
M6+E63fxatARMhVlS1OBd6HvOxbdnsUV6ANP525K4H9/sRPR33lW+Z4BdngStMzE
h6s7FoN5v5zRwlaYMU4OaKW660UHtraH8lBy+B5xSLl/9NtBHoaiQOwFEcRWc0wo
OqY7SW9jXzZsEKt2PKBwQRd3QviKIKvTEcmzwI/P9OO6JunWFPdlnn8lJ0WnKxkH
kIP+YtFJhLM8mRRF+TmGfPiFoSlFqr3GI67TZ/rJTcE5BmgHm3g5MMZfp+FVPOsK
t31yPjHu3JgxWfGUYAqJcMyv2T8MvM49AuxvbWQojAOQBnwyqHrfe2qd91+gW2JQ
MI3ZgVwlHZFhKCuiM9UwFvrY8ttYgVoV0vllpuvgQM/NwJ/ufYJl4QmPYZ+Cq5+x
PbCVL43kXiPrVgPquBESOFLJRWf3OxQJRTFyKWhqlQ6Xq30yDBpSZ66sUzURM+ww
EPMbmFQ8yHZPOndb97vkoOjBUwVc0Vbxzsyj1vuktIHX9zkOCZOmTUt/Ojrpa0+8
CKWPhjX886F3C2+mYOx5mcbJdtfyHUmFf/PnoalWo/82RbXYWwpRTJwcN8T7n7Od
w3JD2RtL2gLfVEZJiV0bj43NE+dTHS+gJCvKZSpn7R4kF+48/lZ7EIBcZ4FWZx/7
QBfX8Kyn7GHsS9xExYawcpMhJMOy7hFy57S5qXynofdBkcEJh7LtOHL8rY62mq5S
FuZXrmiYxkxBMRMK8VBkDHL13Th5BKDwJsXLa3WZWR0SmSwZ9JtrrN4bzrDbCSH8
A8mdnG8vilmUf7EZuQa5sTQufsT/3UmiE7iKiX9EEB+EhceAjp0OUl4PtCPcqK0B
/axjNrLuZZa2NT/rLKAKhxWKGnTorEa5o0vGdOYwgKt7r0Fv3EBNuzLrsjOlekir
2Hu1aH7YgM47Smiogttfgj1NJIbXrhd4KMIAF+/1ZAfKEqP6CRSnr60Oe+ky4Vsb
3PXoH1M2BLungdTDmydfNzEVQ6FAUZvysqlKgpYMB5dxr0kkQksqGq3YZUlLSJNO
MtrlEmiV0iwqYTzRI/ibt0YfkofeQw0Tll0+QAn9txleCJNImgq1+2gPiTHMbcSv
q3L2Hx1YtWmE3sDX2dPL6VtaST+qpCZn9HCal7wIcnvoJgefwGD3dwXCdsyuKsys
8yIgvuJcdNLzwFlXhGVCWJV/5iPu7MT5bwr9gtButyH1LYNAvvRp0ITsRiwNWd4b
zC8MRjcqDlyCCPJB2t5fdiJxcXzX9V9WO/OH0Gg9QiQ15sbemoXUyVL6bAjXyixB
8bCrTsTIK/W/dYRf036ZML7QxVjUqQW3N6wRfd1fPgHOxUgspN/iO9ow7V47PImX
lciefzCrVRf/2wWOSSrPl4V1nkR3irOyQfwHszs81cvIOVzCC/51ocaj5kcx7L2a
R6ccuNFw/7j9sYyMTNzmDQ4fFOGt1/1wA9n491cfhv/pmPHUKE4G+z1XlN9fbt/4
a5lzr4/ACOkTFG/U0A6VOgU0etiOrWSATwgG848BHrfOdiEOzhOYQYQGIdWqpUVI
YmymLpaYoJGCnv5s8M/s10NvHynohOvbRLPFa10YsuqxBYs3vGDONRJcPkt2c/F8
qF/nyxrfS9hqvgVD59xNqBihg3/6qrYOGbS4snrY2Ma9xtHvXdAkWli/DuMMlBov
UEaZymohwOeDy2Cswks1k0XVCq0JeNWGY7kb57qk03RN9a3byw7Ptoda3u7Bt2gY
C0obzB9eqdFjUy43zjEkmJpElQ9lC9Y2QG5bvxLaPPSKuHtAse1IysZbVJnOYSYv
3sS5fSnqEmHLioVWlMkiUdqZJZ7XZfZQg/gAXZKrb6UC6MxLTChynSytpbRFvjTJ
uJONfhEyWJQANRL1QUGHck9QLEtzsjxz9+5e6h+/C4Y+sAlyjtWo8N5v45GBnDFn
8ryMYHpzFN6l/bY9Zv/xXejFdSGM9xm3ZuYh6eWWx533iBsLsv7okijWh88DEVkm
it+o38WKdBsCs683idIbddAkxndWDYoirM3UrxBkbanMbkBSY2h1m+N87b7a45f4
2DJq4ecwc+nyBc4wjF0Nj6FKibpT0mU83DBewNoFkVCYxECZ9zBmQtvvUHH8ahCf
bI7CscbTTYbID2PNRmYau9EHfwnU9f83twf7N2k2XIUJ2NrSJaw/VQ5MKQzWhkj2
H948r+sFZzA231elPYoBgP/FcQy74maXTeMJZupmFyks5XyJpu+LEn3DcsIdhpIH
nKs4V/k6gh/Oa28sKzRO8wqFC69KecDYvYBx2TzPcUOgBU+1F2zCJDJ7s4/KzuL/
7I0tyayngKJnpOJRKPMtToo/kte/Cqe/j34vz16wKH1m1111qRXopaH/7cs53emf
GGuFpjS0+Gt4vLpQmBXoN5JD+0Hwo0fgLSfN4+yO/kQyIzjcHpGswC/bu6CQa+DQ
oNZMyTZW0JjyZ5LnxKXF/1o8MScXKLW5ohHKNNxBITGK6l7B8vmN/li8hN37Mi7T
O6el8aE70+A4D3LFg6SOByqZcvGbK0Qt2diB0Pj/bqU0AIFNZp43mNlWuAuhsROS
AWEG2l3aIBgPIo455q3Tk1ydkODZrqPYfftK8T9pA7SF4o9+ym2rFnzT+rm1JOaC
atq5gvDpzEIOkC0l1Pph4id+fuImbxrle7vyAvdhm2eZr1De6r2eWiQm/GBHbaV0
nSiS7kQCwMXt89EZwHwJwKdgO3c0PyQGU3g25b5apDN/QfxOSTkQQZWbWeE5c9xM
2Z7z0JJj5y0URAzhWYVVRiYZJxea5Td2fbmETTKZwjpQ7Z/gGXkq5edlE4tjlo3N
NE0lmWheL5RgHdhVAioUQ+72HxM5bMrVjaLLSipj7sUj0ucZSWR/Vg7hKwbW2XYT
BjvxZ1O+EYoC8e63lHi5+HG1lN4UU+8eWxSdgfxI8i4Qe3ddtTNJOI9t19ebbNCn
eGh/80DZVYTT6i6ebZatFa2W0LkIKynVyQ155/21FVsD5RZ4vpxixZrBMXxLzdLg
rSDN7QrZUKSiGPrKybiadzTYIOrWhasOlEsB+KnFIjV4vyBILylrLdbnbsf0Rj5l
yjUOp+0cXgElP1zSGCDobZSmwH36PZ+n5YNyeBjAxURroETwez1owKK/gMjCZp2p
w764lK1Q6wNAurGsTa5LrOArji9QgzUIjqbwborLT0yjjJiTQ2d0OP712gRUlq9K
hAwe6obFMyRTvbk9ntwbGHCgedYQ534x7vHgItwLLrf5vcKX4xTYDYqF7wYZr8qE
Fb5wEjAGJX5XWD56+6mcYyY/DkEmqS8G4So//Nk557ZG6u/d5NRfR+ysRZoYlh/F
ylj4iOCZenXEo1+lSz9gi2EpKEZInMnHPj7zl3/bQBH0MfH4imF808HH0Hi/39jZ
exd6M/dJACPsFgTCAblsdVeG0+vxcC/UGUGhWJCDHoo+fgdB7iWr570aCltjcoZ2
tbc5Rhj0G9m1hsStl9ZUxlOe1hCA9PsT0v74rfDBSPO7fH+tR6IkgIJ6lSlYihH0
LMd9jGuB8FhaerzAUY3DvaP2sVX5FnVsEC2PAjPMGgCEcTAcXTCDlhV0zrbPRhiP
QU7LMypNIjy2AEqmx0UbxZtXM0L+6+ytl6jdAbdaLPtFvRALfMh6Z3g9PTm4hhpC
B9FSVA7ERA/WsvB6Ov7IyHgFknWpPrVuWW+a7dNevA4SKy1p6Q+PQasXwl6wg7Hi
riiKY4oj7aMkfUPSxkPjm0RJZ+3a0EhbYoXAQiFOyewfwve6EHusbPyXlWh59tRy
tZGpltDP3OCCToYXLpgN7sZLQ4SlLt/OmIEqudDFGhLrpA5fjzYGz6OoVumm7why
VXTf7xrYsjRrDWDtUGRMPPql0iHpvx0HIT8nTB3x+QcmQ62Zmjav8VVsQmuuSJvg
pxMahD5xg4AUEN+11SqM+OCsga1QjhRXlgPn6VBNkFKVjSX2dMg0cRKSvY8Q279K
viY3wtxPMSTnjm3DER/Jj5wPI44/m1xI2LivZ1nihmaXuQmt4Ooq/NpU8AWktdat
L/86o9TcME6u/uKhf+DHYJ69zmHSW8R+hUG5J2Y2c6mD/1t0tM+ckr4WysJV1xDT
ujovejREtwOyGzowgowbAfSkdreOx8IyzGHAa+uUHsX09V2o5Yz1w8Px6S84niFl
A6DNcoujBIlby4TdZBGnuHgMNU1SWOFhb7ulF7l+yu15s4j7GYRLve2SWcHFlHlN
XKctxPqkaqkf0LJIC+G8u59bUGAFQYWKIdPD23BEOvqN8r+1Wi6vma9/Fj+YzXVV
XlsvNvF0QpRuKxsaS6SCLeuqBQBjsobgV+uvUML5lw+aMLGADhXBVgKq43FOuwBH
do5p57YvB//mj0n1Y7il+uYYuqwELId+A/98G2HPwo0Zcg69HRRlN1ikYkACc2MZ
4N+fDspSc2Tb/iJ8nV1pPJCah4Vw9lertUSeTJutw1x4cmZaWxt4RwdM5cwTbozA
v8eB3N0S47UslBq7tcFD928dZh76RPQ8SKBZJC0d4UyVXW5fb9XvIhz4Shvp1Lgl
kPUBCkjeDXOlTV13o7uDL1bg1rUAkd7uBZw1Tjp4km1eMZY8CI7qOUbKfeon1pb/
4r40i1YUpaMAoqvTse3df5q9SmAU9aHsuvvkSHr2ej6y0NK71tFctin3SCauFGJP
DkO5Zun29ecR6LRxjAFZJIapqSQ2S3gwa0M6xbnWTcsk/0zZHJg7JUm7a1LH1+Ls
nwLoj7a6K84QmZ0mDQiNJXaCJgRxyVndxCQr0dvHwaUeW8n+Fd4pcRZC+44LCCK/
CxLJnQj/rXhRVeeaMjZDx0V3noDynSd5mAneTTDXWLPIHmIdUaEbsT78Nw0I1B/7
xZB9Bo1NVYrpz0Uzlx9vKsGU1L7xxIYB8bUwxHlibv54s9UrZfkdgtB1/0wkJWOl
6ena9h7uqwsJ2R8Fxe/cxsksv8H1ZdhLSyfMryVF2lGiB6d0AGxmlWJ93R6rFCew
Yo9kAvPhHYVn3vx+/ZlARFgKA8Fy/tti2r3nOdLSlDq7yzeTgLpnNdVanluYGiJt
pZarru7mdlNfmGt7g5lzdECkbdBAcU0JgiksyEhn25bAa4P8LWtVQofiDIsiQA4j
2DYRjoKlAW8KseA9ric5DjjBCdB42WNU6ZQWRrGWZlhXQtICS4JN1oaq/VTK/0ww
UQ8GixINDhB/WoTF2umVfeiTcHruFH3gQwUPs9zRne8tHtNU2Mguqwl8tZU1DwFA
1Wih6zve7gBtj/amJ01NCDimLPws1LplK9BWmq8ejyH7dJHIG94Eq1oeWqPNplXS
9MM4WM11KyD4Bcn1eiRebjKPAohEglbWQ+RL1LHzuNPRFA0ZpnL12bfgb7f6lRy9
QwGyqrYBxSQo+pz0G5+EzSxIERUMS89thjsfH5W3elTrMnsnt3x1xIHu9mmkyoV6
GX7jYf2OtRB9brGo/JmqgTTehCyJQF/P5BtqVUpUoEAOSpoIrYHPCoxGXOvmK4wa
n1pUcGhLIl4qIWPTgWswDA+xdHArc23oPMBEDNj6KK8ens6beYoco9qDGluE+lhx
WXk5LMQITEw0sbalTG6qamk/hFzBc3rWqOrngUAu39dTnbS+YcNbGe1CPzWG4Sxu
sW2TtNU+x+EObMywYrljEVaJFYusn/dpHhgR3qcMYx7N0Ar6d6NK2AYXWdHTb2zQ
MNEr5BbpXLEamVJNnh7Pqild/keH3bMucZgmnR07TP/LEiFt/w/c+gm5P/mgp0bU
2XS7Gb78eKlnePTY0xCvYU6xGBxHIGZbvVeT0nYDfLjlwnscjhhlbu2IiLAHDVtB
rzjnCj597Ox5kqH5i7vs/7vRe65t7HchiuC8oUN+ICQ634CLtr4l5MjEMcSkQhoD
USA3s70SuTfhCAeE5rlL4Cm0l/ZHLnazMtZbYQf2Ie7uAZ//keGGNgQF8w7taLLg
Cr+6vOZ4LarVy0+SBu+hFir0G6Vuy3dJeTRbf7GEwZnpx6yn2gMmwPA7UkXsJBvx
POJppY02g7bzp2T1nmbIi9/AD1hrieltLPnY28JeDeNFTXC9IKjV+SVLPD/UGjV5
0slVKtqA3ZeX3jMscU0YxTQ4pV4xJyNBWHlGcp2yMEH+OnbW0eQJLMUIFen23ia2
/up2RklV9FTisrIElbsUqJZ8s3Yfa2Doilo6zyNF2NgAK4JF4rFyYPs+pboA6jsB
gGsFqqG3nG/5DpBZo1MtPSn6Rx9G49BRLru4RM+taPYQA/J3bYjajcak2n6Bt4b+
4PB+rwfk+JcLnRi3z0o/gOnhhZtIC1OoU6Y3yPzxZZLKIWB51PTIhcCnXxFCGMZV
xpuYGzc5QgKeeaCTxxvZXp9AXqxtde2CGEMtS/QvWZYrWMU+BoAySWerdvsccGLG
Dm7zWMWg0AtRLq6i+qiWw1+g8I2nluD60hvPhj+zjLX0KSNrujFYoq4xHm6YOysJ
BJzI/l7nxTAgqnBidiJwFj3IvK+aejBDDN/plb4Eh7eX8yHJrzel+/sLwJsr3u9S
kkuE2djbmnPlquWRHpdVj6s8RpjgSuZWIeWbo93U0dVAXkbqZqGwh66aJbDmkRhR
7nHF1pwK8zI5OCYMdys8jpYPZuFm0gK7Ix+iFbh5ipbsR6Y3qssFoH5mKwcFV4rp
bJPd5kCZjdJlOI2fnLHina4Y7AGj9P4qWgTT9VQHtSUSqlS+kGt1WKTS6thFK+wQ
qfbwbTBVnCkQe1Dm1cN/TJdU7RoN05tnA2pk8t80/jKyKgOWwpC3OxiimrnXs5KD
iSj4LeCoXDikC5QAJ+PufvtkHNqiKngUAUBYzEqmlU1xXChKyyW/Hcg3LPKC+Qh6
PhKDTSOJ7mfFbigtjrfIyQNrHGfSvEtbaWfZfTTfFcjiCwO+R6LARamypWEK8JJ6
CyYLHSgIY2v0O7KtbqIzZ4K4YanvxZSVPGkTMkSrOZBHI3C4kGY2t8kKWpTtDAvw
cFkNZfZVGWSKoLgVf98J3Z7ekcxch41FDQm0sxEl9HJCJpPU/KCkqKbJA8Pt58MP
WXK84jCaZ9W4UUUBmTvJbkORHxjy8CXSkniWa/NyqqSYGPJ4zdhtlj8zU4DWHJgW
yg579wa3KLsLsXsL6unlHquZpS/mxVv6lGbqsMjB0SYueD+XLawvb7UnKQ3+qoOO
gtN3PfFzUPP3KOLJkYXmDZCbltbAGQMCYJd//IqD0JJFzvxRRdMzGrj2eCcRSmBL
jJrIXN9yw9Tn4nm/09ghVDXgMaKoZFGv6W4NU8l/KITIKaOVemBu0Nw2HsQcgpNj
DWsnwctLYSwZmnXzMkV4rfsK2Hc75GCMegHvwoY4f5ForOS+AlvpiJXc0IRW7Az7
yZVHRtJvwmyvxbkHNtw92RvC2bZQ9itwhKXT1LLsFP4yVGlf6Db8yIzdzWjsker6
XTFpS4BJMyBCudH2jiqBBuqbcuiZ6DaQtt7BuktyQrWeY2fJw5c1CI9+BjLyFE0A
lpYUFOGAXLPeShXJDAoWsAKqrY+ehKZ0ZdaGoeV4w9RhMhfjLqlDO1yDWGKHyM0p
CXIFt37Ti45Wdli+QhVYIvgOuMfV35ykbEZHG8txVeLQdYm/gxAL8Ucgp/jxOOKa
OAMQF3f9BetbjbZIGpDAEjKwlRafl3L3R2FzCINt+MO6NnUgG3RWwWtp261V3M3a
al7WneBXt/0S0MCoE75NhNzfDxZRYvgaU74Nh7/yrMWRY1Fdi+qgkOELp65YtiXQ
M3M5R9ctXm0nDmoQUBy02UWH0SkJQS3tNAPS2hXY4hSlUHm/7R6ShcRR+h7lI2dH
e+h80e/JXBrKzdIxkPAwi9PdNA+yrtbK30ucpWtHGa2RiUUR3e+oSoBiUrnZlL7a
cRzwFON+mWdI7rDk0dMqeQazJfHEcc4fZJA6a4zM49CRlZ1t7P0DOMjCmVnJxzmQ
/VUC94T1+/6uE9QmF02ByyHWJOVo+aS4vIyFSAomCWWE2++lUgbbpUgauEd+fD4e
w/eiqEbL3JfzTaQPfLhOEV/5INvkDbStI4A92a3mPE0tLCJFsRZaYlcS6Ac7xnUl
1bs9zEilavkRUgE0rHaLliEBTLynQMHMwxtMYb+GgeUCE+dLhRsXTAK3iBDakdx6
4rJeRwaHf3O8F32GzIyAf5i4IvlkEkGkvmBNVaTF6B/2eziGmr7auPQqasj+cLo2
yxY1lcudIGoCWZo54L1GhwoiTTPtAYhQ7mkoSLyF7714vBrfdgddFhF+YBwXnfhn
cy5Jay7c4ZuXpPN4QSACp0DszYBmhMc3hwpyEtwqpIatcAVGc2of6Vj+miPJZON0
vh7qWGsuiMC5Xmts+o9YVHKhtTKpkr4ApKHn1Qf3/8I8pfgw4nI5412caD0M6boy
d4zJKFUVE5zYGZXKUJf9glwfpEqEcYq9FmETo0+SwxUaDUFZohJrG59+LjWdtz9o
1RoS7saKvUlNbiLJnCxjO5Yu+mEkn7QcIi70MY48yR8Gl1N1Y4Wkc5peerIZLTQZ
wQe5AUn16sqMpZeBpovlZQK0m1rIM517htNoxEf5NYO+8WeJLEu/dyYw23C3B5Kv
J8+7GBz0xuCM5pRreD7INsPdMZ4e9hLDznGJIJUiNC+r7ZZPCTG77oeRLYkGzpiS
38GdRl3gu9KEYrdPuSmSiI/oZvACWR6t+eYH7ulMTyNZQFMAH/KsarOIFloP96LP
Hju7ZKnkF2RpU2g6Wzb8P/eaKUR+nHtYPkMl7qNHh5835NKprmeF15qByRZeaWMZ
xCn22qZ64TV92e0d8r9mbv2DKjryyLTGOWEjkbmGgj8517B+jBmtpL/43IaHa9KD
CGofb/a4MdMIMoVrNgj6XYkZAmxiLXvvhgmRyyduawV3iAgNQ3eHdlOxSFhsT4LF
/a5NZEtR+Ir+uTgpCTo2o/eMxC5ywxlM8Vw90eo5W+XY6pF1+jV12N/TW2I38S72
sO/bROyM3h1Qg/JnrQ5feYyu2pZgMxRhM+rKJ9XUhBL2njNgkbX0ZmXh1TINDVQ1
XTBx36pIuphi/AG0UlDyI8rqHe0xVktONcwOT/Ag23iP6lBfrHNR7cFs8Qs1/tEV
YeccSd2jKffRYATdkeJR5XGlvhKPpCN01P0bhhkzJOTq/BT9u+HB2NAeC/qlauKm
3RlbAoxCwQwegGI35b2Hx1ppY9EX/O+8iJ2iZVlumJHbrpYAZPMqRXcrUeEt2fE6
Fst1rFabjlXS/5cc7yWYDm1FgdTBcpguEP71N4Vd2UU6dB2PkADPsJGE9eB9CqAr
jKu2YO8RlMoD9MpAGgucYG9HwspXWYRKvHmcvYWU/Xwyc8qUx/XwvOGd7m1eJV0i
F5ivqrqgfbLvEl9JNYh6RhVmN/eXwqg9WkQIWcGVtbRimp+3Ky3rXgafEH5F2vBu
R9iNPZBy/dZUl9X0OJE5LpEtsfni4H6ICLIkp6PDOVIY97G1ONqd9ZsC5LcjH6K+
otvPOL9G0M4s8/IYnTMJXsWeBMzf81oRJG3MrINeVcW/817VqhWrN0C2t51KGGWS
oM6vH1nlQCzuBUHASeIydwAzAr+SHVH9FSqVcwb52czweQTSN9SCxiXCMiLVb/rn
aOS7F2Ryv1QxklWvc2pUQdPbNocfkAx6bWP8lIAWqcLe8FpaMrv+GH2O5UssGcxA
Lqhsfe0TOjoJniEl9PfMyyXwAOd7OnSaVupv6IJomXzfdlFoxNfx87xuVQCqa9+B
+nkx4LrXnhPzjkh4sH2ogHr9hVlA9oKd6/84kQhYPy/K6FMxcIYCrZbqF7+XA7XL
5cEeuchew2UpGHeJUmS1jSeDVV55rtX1M73MVbrt88HIkbOzqhIm9rkTI55xOPGe
tTws0JD83+xf/y+/Jtzk1Ix2on6rfF7uMA4DS4Fio8hhIeqD1slWJ0xKDt3Wh9gq
BFMGNXgpb92sX+w+mP0fBIFSbS+KMX081if9GfpWGlAVL3sfKS806b6IR5Ki8c8L
byj2+L0BjC9Y4urehbYkL41nqi6dtgdf82LL1a/MSpi6MHgT6oSGS9uldfKZQqTV
dfORQmqvEMPEHNq6j6OKloiyJzifJ3B5Emjl5JT2453CUaqkXtxXr1MyjmBAHBnf
iAAZ+o7nCeUtv+ZfnRG0hb49AFo6gX9p8PL0WC+OQBBxaZf3HVaesUm2pM5EzBkW
1pxfGQoegDnEgJC+HEZszYWCeJrqahWsx64c1XLQzY0hAimE63LLKqb23RJ+HcY9
4bGDfuSd/v6d2QbY4SPG1Mj0uEUJTO7/MCnldr9jxfXzNImcFuvkl25bmeCt94xv
7hNiygFrSAKCEo5a1Wc57SF0mYqTFapWTG9h19ygduD+0ke/1HQBk14L9aY/35je
of5FT7WVzMlojfeHUkGnhwFT880MySwCCMCMN8/xd8d+T8w1nitI3kSLf612yiNO
n2cZAuZ2Hkp6CIzx0i7T3dINfqjE2bj3YWEtEi6bS3maZ6K4XZo3YQVeU4RX5dYp
qMZNaA2RWLa+FabZXism2M0PSqZrTr1RyMITpq8tigAr/x2mnST5tKXTX2pjkKfh
w7kFz9Hzqvq2OIN1orYG0sBW7aYWPNTbQQwWbTyMhln+345F+5pOLV/ynUKgbtVk
PrG7rlZzPE5PMWOilfEL9abielA0jKJF5cX/3Q0kiAu0ZS2q5OksZWxJo5rpu870
S6Tmqq+8iuny0klHiF/14Dvd8s3Q5VuWtnC3pAq8iwgEXrfVkyxu87EWohpnM+Sf
hQmVTrWFznD0iMQtN2djaLckRupokAidUulMCjjyBWzMZF+KMplAYNnao44dFn45
WfXZngFGz5m6qo2Rdl7/+kE44JJOXZcPNTbC+QCRKAEAcV2dLQyFP3NtmddcTW8V
BU+HViW4cecTBvU3br01tEniobnYXe0Ga6YD6JxfVqLeZUJx7ppaLO2DXShe7w8J
aWded767Z0U0oiJzXVn1yiHF5e6DN6dlrY7CUQY9du5WXlmrfV5K2bBpUrpbSiBI
VDSs+TyirXBei+p8/Jmh18RGhAPZ2VbvKATJdbG9ig0YAosaPT/QjKoHSp8i+zaf
NJaoPyGE+3/F1fECkyBlIZ8HGDbA8jFGKubGs2NQQ5WPb9QNNNqplXpDTYAiX9+y
NHmljqzR2PGhwSm+FCAWP1PfEQOR3pG2nzgJXS7hUZLKws5S1fl8gpkvSFGibg3K
VVDEhkEI3DJ57zZm69wEFVKAfhVbOyu9Q5DpmnogrbuKjGuU8gR4TxXudm6sxMj7
UZpQIm8e2DYv4XIqlrzNVhLj8xq6xZGImTyiTtpxk+hbHHoQF7nijLfYwb1tz+in
MYx3fRXzD3UTzaLVEsV5MhZF4vrcsE7gsYrb5grfWiDAvduVrgeQ19ME6Ifqpe7V
nq3YnBJS2e3vedlGbcKv54lAgrVgNvbRYA7Z2ZUXLduv5b9LgZvWz+s64LB7MjKK
hXZHqSTf5/xdULORiRyuTg0y+R9vP2e8xBsia3mD84clYb1tQsXckHofZt/6Ksmd
h8Mbc5Yk0VL2NjsUD03rdOWSJstwwH9qtzdSoPQesNLbLWSV0b3Ks3a7Cz7pM28J
Y9TbLfOpXXThb2+mIJnSwma2JTxGgbVbgbVbMUNCrLD3YzjXlVXr/v0FNEKRi5V+
CD4JNXgkCHt7H0qrJ5S20SgKn9R1QyBKtAjayWNyWUxG/eW9VPFvG3aWfUQHUIsE
hqdRkuBkG4ct0YzK2hg1lZ1PNY5mHrkHrP48EISRlizQW/1p7DKonQSiTY/UeiNW
F89ibHdRYOEzBscfmVYYQ+2jXsw6Tb+DGHnbzZkuKuqzYwufKvQX5ZOS9eRW8Ujs
bSt9Jic9asudOoZbLo7bX1nhibj+abJXh4JxlLJ79n12uxLfnMyaO4OopS6zcjns
OVwudT+Yy9Sw80pNefqb/UExAR/EAADdfxQ+yEAcN8eJA83Ce7ytFN8w2KfUe1Qa
9JsdjpHg68E4FvYXhoTYOcPP08y2g4trY5WObBenx4lXlqyqTaTBb1H2sLgTHrZ6
/eLZQWffyw6qjYODcgzypnMcKD6Od7m74CxmKBtY/1zSPwoM+UasN2o5F99vWmao
6zwYon4OALmPuPAnGhqIsMU6MjG74tjcSfYX1Eb9kfIbRj94E6tQlDVBgyX7JSdJ
a87Cyhm8HfT6G71ndhIYhvPuBHYhqFe+lmdyNFQXGMpQq6F9htrlGcLp+s8SBPgm
+uXPP4SpzQ6dmFAHt2NCkiP1E9C/7/hG0QA9qh22Hh/GBQq+l225EifJnipBO5SZ
aZiQPSFCsAix+e3vB3I9Lfirescy8q/rQZRQdAvZ0U1J7S+CqVKaz/Sueb+nVLm5
XXFkBKByN4SyTJyJU+61qj5ya+Tv6eSbQhyrbTAMjD5tKf5Uu9SCq1tQW0wLzOmO
tgaXy+HvFP4O5V3REFB1g65C7TxZAOVsom9yLzG7oReVEJ1xtncHzZWOeaIj5jL1
C4cmQsZPNSHOtk4IxNZE3KyP0KvOxtJV0RQWe4Z4tUNltabmDFRN7OkhKJ0L58Qm
vhGy5o2O1BjOSi7MgPjt7nFxromo1qzy7lk17kcKMx53FWtPiiLx5NIYqHBnuKII
u+wgJf1FKDWlG6gurgTFOT7CSWfoy2FMxZ2br9L2toioTtvpAD+/oj3/I/ZEBD86
ew97pIVpjTZsSP9gWwPcQvEUGANH1gVk2aWQDlpq7Vs2K6waGskzgyZAlFhIVGmD
/1azLzTddEvZvpa8zgbKGtlYUWfJ+uxRaRSpziYpID0gVRvIAkkousF3Ui84xsou
TwlQvRZ/OW17UoMR/aYTYnpOZt5F5qE8DVSBRqcCsWbyNYDnZ+xAiQrn02KM8WhU
oQCXd1PXRXp2/ZoTCC+UIQCKZ0osa2Rl13u/U4TeqgQxPfEnZIiKfv5nrlM4L9sk
nAGTg4VsH1XhmfLfiK7kVNm/1zb5CajFpL9aN00S4AU6vPZ42q16EMDcLxBGRFrw
PEAxVJBStJFViNu2pxpKEPEhzEwUEF4Bd9l9/ZdJeDsiv5oK13KiU39KjVu5p2VV
pHifJN3Jige3y3JRrgKRnX9JIuQaNj+Cq/euQNBYYyXjH7qnEVSRP40eHfeV0Fg7
QnIUT73LfKGT7KWJY9j0epGrzOIzKUtHGv+9672CgXv6jECiU/6MbIX4aaaugD/+
4MAQMURPBLM0uJ5t28wiFjto0gTi4u+x1JZjLELusi12IquR5NG6EF7mw+/e+ltz
1xwbIaORDhlI9m1oSHKTXao3mNCCGF45zbq9OlA7INUQ7/OIOWZ5dIHSV5FX6NSt
eiIbUfyOlnVEdCdg+zlykTFCvcNpRHi5rLODC8X8gUMJxzpNJ8RGxpCckcwFxBAj
jpZmj6DBxdM9++pfAUqeOg2eGEpujhWSsn6Tohuzqz9/Gd2G2Xkla0KQ1Xq0EL4J
KKliNgIctGU0ZVW+vQeK72+7W71UGiuc0D8sW4oxkLnuhsMe6/GM48CXjHAaaf57
AWfGdTOXHMbdidXb3CVhevmxFzjbTD7vAI7GGCwfOCHDg3igLjhDrENIgQBdrK+H
GOpOqfFzhXV1RvilZxHI00y6S5/ashXR7xthi5h2b9MpnpSuXsqVbQXcu5ykH5Sf
ulEIAFVAaidX96AexJ7+Mw0bd8hd0UlOeHQqf/cL48v855ARkKzJgmBPuRsH6VZP
QVKa5l2slqh7AfAhpSA4qXcSGLxq/jJuF4AP5ZeDZL5zlE3s0AzZ/ipuTf4L03lM
+sSNxLZna/vhcKVh19iVY9OP/34Mky4JzDCDlG3YYu7vVN7wWu3OLE+1VGppnYhm
njoA+YgP7UfZhP0/tPzgfMdIME3CulE1MTFyN50mRj8hTnQR9gJhtEemFaYkI+Is
5YfkamOg8kY1ZQTob/QyfYgq2IC7K0Flvn7T5f1P61y015Ksk0YRcm4V1KVG+lr/
sZfx8aubC684CRwuzJgkO84JIfCmlvD6dt1Pblr6+u83VF3A7K6NyKi96mOTBIPE
7ZsvNIKYm/RZzlyZNLQB6opfpuzrMkxEuUbXzZUDRJypoXYqXqam+OqAEWxXcoTF
KSI8gtN0Y7mWzhLNR82sTi0EyfBg5o0ZPfmzd/Dbm3Sj4lh9Lc8oiP+DX49yDnLA
lSXUaNC5353OJ5hbpKy5D+8E86wxiA7NGxs5iMHIoDdbtLUKwZc33Ci60NrS0Ad/
bGBXKU3AP8K23FU1OKU72oxaSzdcisdCu28RduNI4rib/tv18CAUlQHSBVFIOlD5
J6NMqfknKUeKrmQ93qtZkpEsOKTaDUZqF3MGLp7fdJz3kVQsl7JHUuJG5O0qXH2Q
yTtt6DvUPDOBaIZU3j4HdamjoUK0WCFuThJVt8ohBG190PCFryDa0l6BraxYibxj
npXpyCeOOwrouvk8wBx1Zr5Qjr9R0uollpQHt2omhCd9srYYFp9PY9h4sNUTG6KS
XdFDShphmjnqIwYZ9qWr3lRvARemnXYRxTMVMxF/S3P+ya7CvnYUYA52DoQxyEoL
Mnj9PiGJCMNRKvQVIMK8v8sok8LKQdCwYoSynbmgJYfXOGU6b6k0ZWZMIHfThExN
q9hiv/IzxpqbEi7UiPJmv1s0PjIuBnOMzNUiqg9Z8jv4UtXhlqXxmGOn5ILqBdRa
kfoNmMvIoVh7qe3DdJzO9jaSDp+0HFZknwaotH5IK3NEqz9esPA933/QGzv1BKmZ
rfVZB6P0DKR9zCz2YJmJT1xJvq9oa0eEHk/PrIvwfY6+p5TZo8kzaWI10WA3XO5k
sBccH59jOVVZhN8UwH3mUctt16TdG5/2x3Dp1d2dWLpQz32tO2XfJ/TGcWqINlCz
ZwGePqjeMduYJFRZWsc16Y9h3h/99kQmVrbddGg+yAvP/IwCAzJV+VqFz9s/CuO0
J3hkRsFODs35hD1ceIKi+be+4Lz42o+vPEzbH91YPefd/VGtFSm9Ajs2MEyNL0gD
/Q3JG/i/ZSIfUiF5M9ufiPF1WwRIGwiYdirBSxCvhKwlkW1PIpgOB9l/rzw6YKlQ
3jQJDwnXBPiN1nxma+ywcOvdBGA1gvSNB+8/nm7z6hxdWztapmI+IWMCbI8EUg6C
XBh1N64QHGs5fMN9iFXTCJd5tcaGU7BGZMFcFTo/McqB2Mr1N91ujSN8cQ/89iLp
GQbNd/SUIP05QxpFMniasOT1u9avVk6ReQYVETeQW7JmoOmi8pyFuPqhQ3xN8yZD
U85TX9x4RwsDR16t1z/RgOis1CctqP1jRjw+UL4G8ARitqZIp4hKFRDKYZpEaMG1
RhUMB1HNp32NS947VwKvfo+Q4mHMZBEfBW6cyIRSdxxi7OzcrULMUh7L1NV26fNu
YQW2J0zoaqGZQh8GrUt8J/eAXcqE5a6RcJWQ0TjSbOzv2Zz3K0R8wqD3gt+7DKTO
qB9XFcaZvG6+j7JP5OpOdoqvRQPlK8k1y7LOtcIXH+VWyE0s6Juhx51rzHoaYH0x
3cfeA7L3VMfO6HPJ87sguqlkRjMX4Ts6s2uqubEfbzIHxkb9yDNIFvprxJvtTLOw
sP+CU9g/dY0NKHtSaOBsUXAEUJLmnDZTQJKZ3SSzreD1e16N2eLIxJ15Kqtqdjng
44/FRy8GGN2kcX99LCNvKjQx91qBbYmiBidat7nomvw90Saegs4+kCWpSvbsxVxy
qtgZZFRPS8aN7NEmK2LfoGlCpHNzCTK48aNYY/Z9TfCW8jFa672tEsXJfLCT4Kk7
CDoYcrakkH9hCFJKoJR6SX/Sv8ptNDEKsto+7GBR4E33U7hEv4fgys6BuzKFy7mb
K4x/JqyvYDH1D2HnhR75H7XFg7+U/cAMsjwyZuoNdVw4miXlKpKgbDtUYZ9uKEBI
1B3aAgHdv8aSKRY4xN9m7bnsBLkUqoKrLG19z9LQVLT3sIZanxdBfOq5qYQK5ij9
lGa1wCZBcN5hHg6/870+rZp42k7Vb/ZLOZOiD+7bbtVWLL6xrPz41ldvqnNl2IA4
eR5G7kO2IsETPsu/iEG0ihQl6cWEuq2z6l4cBi8mOkvHkhWrkJrrLzJM4zP6+HNg
8/yDHJz554DqujQUn8ZpM94T9RPRkkLTvnNhOsnrQEmjmHFcPxUFdS0rneQ/qJW3
k3rhNJDQQZD+tU51ldhMWhoKM0XCpMIaftYWbKUK431e692mHJXjuiXJp3O2hr3C
I2svHO6oD8xDF6vKWVEUyPzW0/X2Xec0PxCy0LaypbASdivvk0VN/vpfzjXvl7OZ
+SPSt9xeKCcz/6EVGYsAhAndUYbBCNpVSXJLx1kGg2tqK5DMSnl1u1Sb2LXdnX4j
UYYm+jm5r4YgctBhOni8qZkMc7nJ2iJ28KqhNQg+lrBk9v68ICKhreM8CwYDgV7J
uYLLcaUFvQ07syul0kO0/sGbd2nN/Zpl8O8c3dlPrhl1Tshj4bct4H/pOtFCTS6+
5n9r5HTwdFNuHk64uyWcEpRHQFhk/Ub2Tp9iCqL0zQtq8Ffv3yQsndA9WgoOmyQ8
UnT5OlR/7XbiTDtQaTsUzf63IEtRViTo/7/eb9fqYDauS7O0qhPicThAYB1AjJuH
OYGvc6hN3qvLTZZ0YH81XpXojMswqMrm1f59l0fzHn7Y/EQiCaEi3aHKjkgXkban
rPXrrd6u6Fr2Jq/lrYpqERGCLsHkWO9QcZv5s/fVs3HUNnykSYvsh+gMHykNDhjj
d6aAwusdZ4g5TDjOWpzIkSdVhk3wEtKKaFZrPAbVq1A17KjDGQ86fmN/U5dlWQR0
BcUNCrW5IYk+0DY8KI4PwGjSpxcFMcqhlzpY6Sm93/qOXMcixhE8YXebkx5VIsKy
iHImSKNhMfWUthv2SuNAE1vu0VBEbyAaiwWZjZecS09wWqzSyMSbnnqGztcAgZtA
5yhHrZdfJyx+LGqaVyQsp82VOPTUACK04ogLNga6dqaR3eN2QXaqNlXwzSU2r+QD
jLQZ1QfbRDApyq1goV2ioLZUFMcZxtGqujueogLBXtBGvUwKWuwXBrT3yR4Mk1D0
P+/WkZ7ftKewxldVxpknwUIwBHAczVYdwMDFmSRA/fOlDnmDjTrJPF6LImB+1SmL
F9CoXurmLIskr0QRMT3vDf8uA0Ezgnh/H/t3J8elrxwDT8YUeNjhPBSN70SH/aLX
dEF1gkLsZtjT0T79tWXHzrm+5vQu+0vanNFAlir/PRLXiXajoR1r8Dj260l3iFHF
ufb+ONCWKIz6YyRXO7paibVv1aFVXT6+wmN4orbVRbS/BsvQwYNj1z9bPs7rRC9y
DG8J0K43s+0r8Bc3BFnbwmf2GJQWUq8G24vnzg3Vz4lZPEHf6QzqZQKEeSLXMuLz
UcLve8AZlOD1rr2NzyV5c5s6cccvVcRyLq8GLAoy2sBmGjZ6JIgbayGbUZS4cafv
TjeEvzlLaNvLD09PGw3M8DTkiP61jNLNqDn+C6lqI0a4zCN1yCTOTwPUnQngAOUU
oowwTh4SVcBCVwN3XbAdn9xYI/ukNr722Sygi/iwRHZltl0uF7yY8idnm4zEN2dI
t1HB1qE7sVHnERJDK/t0zMA8cOptm1wCzCP87APCA6WCTqnqr8ZU6K95Sd84qo3e
U9+M+Mwc+p8Wl6gFKxa0sjkV9scL9hUZX3C/SdkzknrWj0tpRkyFyB9sL2jTpFlL
x3m03dgogkqc93OM5RVpzs+vj2oec5ouCZF1DKs3CkgW6ZbV9cyUSTJCc3P2hur/
4hfSuD1W4+nvPfxtd9y98Rhj3EbjHQoN5JtRgDHDjJS261BvuB3mlgRaAT4pLfBZ
XYfmiDZlRNA71H+NsIgA7M2kNC/WpAKvHVfB4lfJoOmi42wIOE1+8ZTa0h8qLa3T
UdeJ6OqrC4jWjYr/YotsbSbtt7FZc4wgI2L9qsWm2oyLLg9rbQ91n+kkyGusqcS8
4OrIF9Wsn62xfn/Vp0qxdKAoqQ95mhIMjm75tDGMQgOMNuraZhU4KCKQLkHMcxU8
KpT9UsL/FPB32qRoKtDDLiVCro6btqCx2XAZd0v9glnLQHWpgOyXSzVBHsm2flS1
haKjWeE+xMUu2jEebhCzKIkTO9x5X7d/StufbHbSwsdMTZgjZUWK2Mpm27+pNCo1
Wlh0pHdNBO4C3JvgytFjjDtwoT+CSYTsY92Tz8VvfXwXLNRyDh8nDNTVkOHxGoIN
TDzShCHpYCiBfaL5Y7VjVTQ6JeSct9y8qWzkWOaMug80HfnOFlx2thW6AIb1Px1j
xwf34cJutS5gyOgXXglOZCISKbUiMAzKFWgpQQ1ka7z/1b1JuxutRe846uudJV0k
18Blepq4VzZf2aXyw3nSS/86ldgzlZe04DFMUKYuXvb4XlNTkxxVbFRX94CtDFQZ
XH8tqeMjj+oqYT8Z4NKjynkU194pCsrGJ5IX1GwWnP8fGF1vUFVNE+VfUn/altlz
A5mCgakxViq0K3pLq3oHykABNl9wcKF2VOPho4MxmvGovEzocFZzfxhfS2BCyBLm
/4iEC1NK2LT44NS549SOu2LUWDmKZLwR70ptBbaRYXOoOXetyytnO+r1Cd1eEKZF
oonw4431aGuELvPRJivft2q9F7BEjrwJikV2BIunKOozRQTEqgb3BpEDrCDy1xTO
IXeaLxx+H51ASccnjMKamc5ejLiLn2RyS77lvgHy3to7hQxm8FuMt6rDtsLMgotb
EV6Gr7bGN5kPUd/ww6A4G2iEDuQKU/G85IJRH3vtGlX1Tel/8DpM7dNrgfgXP2dL
EbP7DRstnZQjTKwVZIXVJ/F391iFsgZKsaXs3SWsR8x7iZdi0//s6XJuVediYi4u
ZiKA9Q+EQLmh4tQyg+UVgVssZ+6H5LVrw30TUMtK8AHwnkmxloTAXErTxzc2VnYr
GcQNsWZ6P/W+LsgWHYUmAo4uTQgtvOrYHCBewo9pnt4oBr8HMbbc1j8xKKmQiQek
0hJDSzqOkCCeiCnTyPtHef5WVz541r7+Y8Du4Sua4GMcq8xSIeo5FpgFW99sJTm2
pD0353OqEaiAbc3G4M6Dd7SqfNPuDqAryCfnm0X1WxexaVYMmWLE+CgAHvgEz585
9zYDJib/o8yKYUe0rBG2zzg5nZCdoZ3GVKjWq4bLb5CWsGjrBvL/v6uYrjj4+RYm
D4lvReDDnZGKsllgfRhkfD8KRHhS6qIywQ7u/laNrr5cMB/nlVNMKuqkcDui61ty
aS6yDSbOjosBaAjOh9LZWPpXh/d8IfV4ze3nRXv/DEsxHMQKJwXLnwyxIx7J5j5b
/R7Cmmot7RIP56y10+2LQ6hVfohvjpqvxJnJsFds+9m01qy1TWb59kwDftZQg84/
qkmYmomLfDD/E4Zx8cpwfsX4fgojfbp0vrNqQDlOd0swKRLl2zeAnA+zhDVemeNX
+5aguQlCJM9HCz2/CnerSO7QXrKLSMB4nOygne3Ew9HrlXNLOcz5rTj5ZTNeFjzj
kChvC1cRgHk6YDqEmpKEC91ZtDC5rPAzqmRRbTJdZ8UIYTKUnqrRtRasCD1pi1oB
cMy3ldG4Gqs/ZJkh6Epd5bobJnwaS0UvU6W3KQkOqQLR1Yhu4sXO4rxhveMBqCFU
dUfQolZZV65yBrwc6oskp9tVfOHNJicq+oXwHsO45Xv2rLzro1d2TrFtDnYdDD8W
NxboTOKncxDaj3uPQ9wHiQcXOGJhH+uYReAeVwXtHSzH248ptfXYDArmhcbLe9Oo
HXmkaCZ8VTpXZeZOAfNKx+koqBiysTMfkMxTaKhGDKjT2vfEMwdPlY2rMaQTLox3
QSkejZOchGn74Hkcz1YhntjBZ9Pu1IHywa0LNzoaRerI1pF31ouvQD3+4rYzq1Fz
/UosgZrIh86VGOLvJFYZK5oyNYCDRi/OoPVrxaGez3fVdMZFpdSYBy5xfBtSnp7e
27EmzgARCKMQWMHqmTDjP+Eci/l2amGntNde0//7ZP8MDeP+ql6c5KI4KojbrXXb
h6N9nmvHFwOr+feuH/bNfeTycD9DwSlBDH1KEFcpNhLyo060uW2NF5XUpxVvgztw
4vhSsadcTyXJ3ItBdJF2E6pxokwPakCEDBxn4OvmxlqRATOBYygjN7WRgE+Hfgco
Ch4wYn+fajZ8rqEe6ABwYLf2M1dsNHBR2VFaCuutmEkYxCiM9TvqC9WvHrq3Lctv
huwrChMC0oxrsDdyZeSc9awMN6jrukOX6Jc9d09Yoql2UnCQsetjp2AYCfaMxnvz
Z3Rv15Z+u/iz1YendADQxT+JfxG0AvI2LmAOk5koVZH99et6c15s7I69WbMV22Y4
y8zNhUa2E5tHM29JFTPzk5IMSQtZglFHPiN5LqMjFxQ0Mtr5yoPIlj1p2o1nXK4x
GAtQ7Pw/GnC7UGvNjSGDw8PXOtMllAJmlNYqZFmFTYP4DCBIatyV7+Pw46TtZRTs
mtKJsLxtYIx5CFu5uSWdr9iTsyYm7dIT5cYALZF8t8zUqc4fIDYGz3TMK0lTv6ZI
gs6OvKbgoqugcH7x3JjMMW3JGvasg4ylolWWMWDQ5zUbS2pI1P4UJGmkkIWw/VDe
UWRXTMnj9JLnTs64/H6BaNlgck4qkRGzJ8+rMjoBe7U87yDnspdy7tPj5e8MXrHi
LjlqsPOT48VkAnGL7/ArSVQp0+2BRZj4vp5Y1B4262brj+q0H3YvfPM7ThTESG2s
JJmxNZhe/PrpGJ8Gyo55t73OnHyiqmQmnGdaV5YNbJd6hqQVwCHPjv6JQGXHjrpp
OSsQh0cWeaL1hSQLcdnfCws1t86nLk4r4FLww34rnIFns4jt8yjZR5pMGuF3zEGJ
v4XKo/ZIQY+ONvK1x0JIIhCNlA5Kd6z9k2uFWkuBiFghx0cfwFLocHaGyuUMto2n
03JgMgj5CRDyxY2bkZdNGtR54Ux6lqUo3/db89MJ9RA3/zVHuecXfWgzhFXsPhgp
bU/+yJ7MJgKjXWxOvSU63+MI9a0JZX4DIFa1POdY5NAzbkE9tEssxxSRHFGp5noS
0VOMOFgxd3IqY6LApZBbJb663Ef6RCmomqwPM2DTLyBe1nXHkw4gYQqzM8O7HMQc
+hyotn3iSlxD+1SSfiqVEj1diWemX+f9z3xlzUsnF1DE3zCEsV5fnB/pFuAPxIjZ
FGSGWWRqKVEKhnhsG11Q5gPPMU+qJgMON8LupHqiT+08qIchK4jY56tL3AMIAZM2
6U5B1rzj5fmTKVopCuctwunJZhJB+aiqaJOd1oFRTBIiLrQm/KrBlNBDVp7ut6r1
d1ckOMNcx9Tt2s1iOloQzPvx7giKmCIjfxSeVM5Z+KBIgQgm6k3PqmdHslIz74aj
BDbQjuviJdj5DbrqpPj5M5nWrGN/CzyjB1S3zq5E+D0k68DI8dhJyURsS25THBWL
y4yfpu31iWH7XlMcpgUgBaje+e3FmOIE+Zdmkjs9Pqv2GnbJLqk2HXVK7t+Sm36J
0SGjqh795beXet6JPxjBTcllzVaR/6+LCETr/em+HqYgMRnS1cg9M/kYVo+7s0O8
XhFcEQ7cwrn/U5ALycljOSwJn9gWGf6GRDE4GYCl0+yxEkuXuWlq127ocvBhtma3
LtelkaLXFAiPhiZxSzE+d3ofxLY8cdekuw7dG18YXKQbRETMmeNsBqnWaFJ1vjjB
JR+VWdt2AUT7xh74omydhUWQJNbv9GEBvYrEaHIsx745vVdRvtF8JMF8t5fZ3fjf
gU8xtRsHBu9ldKxXBI1zsu0enzZhb35996K1A1fV9xNARhB30cLJFHCy6QmRaGvh
offSlwHF5zdXW7W2NWfwqO67wiKHp8VfAsz6+dA1P+HkyX0OnP5Pytw8WMMkIV6l
QdBJdXHVubvGQdN+Z55TLbgQhy1QjhEtsUxcY2FzGZSwnn+W4k+bGjYztBgimauW
jFZ/jv+z21do91mPC5Z7dRjndjidQWqVWPTJCsCUDvuye+dbdKN7Nj3FaXfiNJZL
OxcHar1C0xkfKfGLOz2ASEgEdMV6CTzPs2Q82f1xueFDnxh946DTEZSAPBwz8mxO
YXAsB4vvjqMT97hBjArcVa88L2lU6usm/yIKNUdcDSfI3kfAVlTGlOIqJ+3UR92g
s+y2xnonwjt2XLDRjf6myYGNCzcivHcltny/z39+z5rX8pM6jIX5uvlITdDQUTqr
V3HyHfgml5prTnM/uehWLju/INEE5vh9q3nRGzXIpzWVnOm9rzVQiV9H+43vnyq8
zc2Fv6EE7nh/B1twW6T/HQKLeNkPFwnoXS2MbPq3VMhrvpaUMDU9GxU/08QssdO7
vxhmIYD2Sl9iH8ce5YL0A+97v024PM2VmeHXDqzp40Lh2zi3YBkQv92hOCdXFLnv
0PXkxxBkcvbW5Ta4zhAiB5hRzsWNak3lfuVtiyiitqSEbnKoHC+cRw+e47Z7Rx3X
ik1AdidwZRovHM55DPf8f77P9w8TYzguG6gfoubKm+LpIt15AzsGrUpy8+AufLQq
APpaL8T9LyLEIfpbFljQ39nfzo3Thb7qsDox4Wwrbokj2Owgp+OyJrkCFQ8IAdTK
bQAkJpVqnx0D16EpoaV+EVh18ul7xkFKbex2rZhs7TSmFZ29ZbMMNLMmacrlLVuM
iDij912UOrWY6LEuI59k3jjpya/lYjTqJowYyrQrWPRXnpugQSIGoX077RFaCghR
+awgpUAd2G6G3YAjgJhzh6Ihk7Y0oiLVrwGUkLJYoDtnTBYqei1Pfks9UaLmfSx3
dTJhH2Y/sNNWFg3cFtFDnyTP0QPQisNIOx4mayCvEdTn0fysolR0vnVSRAHulE2C
qmJohIrYr/Oi3KJyDrE/d2SuCviujjvY3fCFXTrO/AIXfCTNQ6lJQt/xrOulzGiT
SvzVKNvahatyQTE21FqHerTOM7Qu0URBRyMgYYBHNmvMibCdrvy8WuUYSv5+dyl5
yCFcrl15fxZCMn7q7z1gPQxYW36cr84BMFfjCQG8aEGddepGrCiCCl1jmaIr/a/f
kvSZGxysJE4ygXNL2ZrfCyV/nXIDKhB8ZGJFJr/HS2T/se1tHBOZ5x2384gAk1+M
e2RyC9548FIzN9wpqTkEwzEXM4ttvkCYk2sgwUePntHGAyK2e/CbM/TIMmhAxXJV
jXF2y1QlbVDun2wBGC8OOJaEDtPl5iG7aOpwM+mQWU/E/GJla30mCZ9lsBABg6zG
fflCctfVtTn61AQ3qZoYh+7+lQPO3gQTnSC93IOoGET6iQbC3KIZzaRM9tumV/dB
8xyLbY3xZ004mCHiOVQI6MGJjAqdtysGXFWNJ6Tb9UAGBUo9j9iQxjFTYd2Pn/9S
ZFl60rlM82DJ5VVhiA88GU5u1pNe7Z1ZzKsB4ygqWxZSkjlEoPslBkO5K8WNyyRi
RAAQFZ7gCYzauKvtp+MDU6cQWX7lldLj6IoNFM6WJn/2/yw5jHFlyG2+6XOoQrN6
rK+Bv8WtJ2VsuJym2vVrOFJRpIurP+zWH70+IQ+Zoc5VIO3KAWObJ7oOrLPi7NRZ
1dUFyV9nUoQj0gJ1mP+D4PGFE207ucv+rTY9E4TlWh/rAWfA94D5tZjWJnkGLnYa
PFOfsYb8UnLl8umvXXpLQ3m1+74coFC7xmCLqWzaMGpZQ+7sYOOSWFPpR9JdagMJ
JXv28YN0N1GHtusAcJ9d5GAueNDir73C+ifEmp9WVYtuPOht4aI04PAMWKV/AMax
qr5ho0CyHzVCRDAyw20uCVAUWMyOxsSA7Z2BiNKLUPOXzB/l9TxhPSHVTeuwfRx0
blYiNqU9qcdbAyLgLJQDUEYGyQvggDzYfxoCrugAp5Gq2XMCnvBKGetqTeXc6+So
bhGY3d/ob4ij6HsDIihXubz+oC4ciEgrh5i46+yHYsp6epEn3EfviLCBIR/DLNW5
w5PJLcqTfy0ZsNmGffbOKdrRDtmzmxg7szZ7O/c6XuWts4Z4kA10uffNmHWDymdR
vu9GWkt0+dGjeS1lyUETAnuPqdRrCuUo32pdCHFBFhmTwlS4qvZKBAWneb8vP9XH
WctmL5e6gOaDJXX1bjB2GlyZyTVoJLQ7WVINJC28ahIq6lgIJtQatI710/EpQeFk
Vn5KXthviO1uJRtSPL+zanNF1lO3Grk4WUfGd6s5GfBnzQx82h1mtec5BDv32rwK
YZZaZjcCqoxI7MRnvO7EdpseZdsp8hcLqkzfvnstqa/5b9PH6Yee1ZSs47NvjHP5
fOQ4Y6y1EkRIsYPq0th7JS0hoG9ti4ORlXmxpaT0hwTpedicpdBMF10K+SMqyDkS
KW3C4GBtFhmMQJTSn00T6bXjRSQcVF+0AmrLmgM277baFIRcsmYGwpqZS0ppZnyJ
o4Ja90k7rAr9LO03NjO1CR4tEreu+0ElReSaA+x3EEXKcGZ1h6v2M1k4geMepXh9
gvuOYdzfDfycJxtJCAC4KS96bljcZwn2XLTzPPpSHePPnLl3DYYEQzoLA93uYOEg
5JNq07JRbn5ZrGsO5poyz8UuWBMzKlp0dthbnmgQ1ZH1XQ3np15yzCiC6EWEP855
8CBakc40k4FHLE6s4qDtpXtu5O9kHl6JA2YhzLc8iPG7NwfWvMLHthGfcLLcHjva
XxftOStBWDyVVSf8NHQdRVnYp9ZRzZwJvzHcCMGgnnuDOnKQeZI4T/ZayKn8ro7B
qxL1roTzMuBPySWcEF5hOzfxtSzpBiOuOHkM/FK5+pYLTRad/iBJjADJLufWCyMl
rCBcC06U5e9ugebK+lP01IuKLu5Ud++LSb5nTUCm9XggiUGMkOXztmJyrmyLVKfe
/GzHD5ipBYWR3eXAsdQaTzdMD9ubtU1R/bM6uG2k4Y1Le21RsUa1H+wtbncLHTCA
GhEyl3rrmtGFKEUaxaU5GhiNU2mo0/pOb28jkcR6rTWGhj+h3Ktp2lvVWmMzcOB7
LlBLUpl3TqsqcZapsm/TW05DT10mNlFPHbcuUe9ac9DYHIjrpFkE7+gjBopKoVGh
U9OUbnhzMmWuT2Dla95TtO7Jqsw/nHIbneR13+4huqPMtMA0fsYvJpEE7w4sDIVL
HakFmHD0xK0vuW56iVxN3aQfV+d7EfA4txV8h0xsxcfe8MTzTVMGxbKRxAAQGqw/
SUoLB+kPtrETkgnM1cAQwEuFGU//e7PwKPknlVzhoTBv6LGQQqk6+aRuOasqZ3dX
sBQqqmxu2utUxVMXAVVhx/uvaGHkuU/ixGNwgmWw8UiHzwNZM5D9BVwOsxlV2LRk
CzpLPStO0BABBX+xoNxmUZpLMqa+Cm9oBGFfTDtQO3IcAJ8fvWosPQSTF34tCQjo
9LluF46PJLbB3QafbirGtQI7np4HKG2CAHPj2LC1wXT1bM0qxzfHf71oAv1ZqMdf
eueMQNrQNMqay9Tr1F8hQ8Zy7GtDaPc42ytAsMmKNWXCzldHm8wcv1ke5ueUc+NT
cVGAdgpG94Q7RpWs2hfiThSDNolj9oJyyteQeZU92U3Een7EeHowDbEgE/sKaWYx
yCpa5X0QUQIYXKUXL1QFpcXhdB4Vo6IMRXF8zwUh7fvp9JX1/XBO2BJ24J5plVOR
wSGp5D3er0nAYnM2oaEJfSYxbD6wF2SSA5GycOd4FPKwgUXgzNEMwbPXATH7puwf
F+5iGpOZit8cqh7PUFwThsLyzzZ9UwPSenoCe6bDKsLZtsP1mKGnhjXsGJG6r/5f
FlkOwfMUEvCf4Cxibl1qaF163S2r32LpDUPrMNQkpdITIXd/PlSiKq1HhB3XQyHx
itduwKRTknqB0ZAtKpH4BadRZPBjkGqyMWYA+9x8oStdTLcB5rnqgjP+OW1YqUs9
Zs1r1bgTu6Zz0NmYb1eV8zqPZY5xmjI3i/dpT5OJKy9F9Omuh3hfev3CBTZXuA5c
sJ5aNLJZzLlBf2dajl4GnBClQnEoKijG4f8fqB+TE2p2oIst1+bO4vYI6w0PqmC2
3KdmRCHB9YUKPQsXrH+j3YrjhiWeabqDaoh//i3ej3LTcoHgXtj6+dS4ZkIfImsN
Tjt2sG6G795GPCaZPi1JXQVwJvgQwWIDNHhIWNdXuYbbS3EdafiXxBaCWyI0dZ4H
kCvqM2CmGWuYCuQ50/pug546PZ6pI24P8AJRhq1cIdcjUqcoV5E0hJN6t/6viq/E
5SS/gZLBVFpJxM73x97aXUgUHjX/22IdECNsPF0CMKpyiyWqO5LFB0ldz64uYEKb
mXlxWZCCtDYkxtZsJg0dArqPH+FpjNdc+CA0Csq0SUlV7KK7bJx+C7Prn60XW4/e
aQqNC+1IscElbupQYH8uTHKIbDfvW6weaD0mz7mDlTjPzPb0oCMl5Ro9uN4ey+yP
1GwckN8/zOV0MXY4sVxxzTSk3AYj0O3Z1OGI9drVVf3B1urCLJMg9oU28QOXahWr
jD6mgHWcWa0k5OnTS+CrO+dzxUeOafzP86cKbauv+L0PMPNPEOTnVRLhNnQFZbEx
Sntqxz4leVEc8fkRFJ+kANopU+bkDzbXx3X/5rSQI7ePPvlC1hA4TkmpZ/7acPFB
AsaI269mqiSVTp5qmqd0vFhE+cwXknmRf5GpFBgmzaYNIp4QD8UGgvYD78wjByaZ
S2BJNUku56as40MHYXPsjSu5BLYVbhkPjueEs+eePDGSI3+3qwbvaBr5BMnIcAPO
VzCjF7ORszsyXlc65fyt2WTjgKqAMLA90ORGKRiagDSk9EgYSqOsgCshOlbPFJrZ
OeBTr7qXDls6JzGUXQnZE/joPNwYGzccvSMjvguoqlzoka757FxRqisVNSqovo4Z
/QOsowtUZzXRSYB3RquSbwDZS8YPvDUYO1gTdvHsPjnNbN3lCbOffl7cyYaqtJE/
+5ND3xuseOwyXg4vc3pBAEErYyWeDSWOUmBCMuhPPdTu7tBgVRb5m4u7TcIzejqD
Apr2o7UfZEuHj5/QbBGI6Td620Y17RxH2AiwYK92uMzFAMCC1KZJ6xa4lfkW7C0K
6IesuE+Sm5qEeZ6Ligd2+FceljHiuiEelijJzmpl/CZHNVtAkJOvMotcQb13SUVr
2s80yQN9n8z98zdxoqHbxvvdHboqzF+uAwUQMcouiX3z6ikx8dHDS2HAN2diqd6z
NtiFLmVmLSMKeJjhf0FCwuoKPAlADjGhAlqsKgbBXsF3hUoHTvihNYrCzuPybPai
awzFpvxgama6jdflfHxo33kvFX5RuS9XrRrKSx65uBdQHYMXo86tVErDqDVol45Q
121hG0HCISIrSdt0PZNgHsLnOac/0tq21WoPdCS/xFSz14c8ZGxGcwz3kAbS2yi7
r/HbyuDJ9+32OfoP41Tq2P+me23ohPxjSgJvpjP+Mi5hTRmuP0dAmGHA7TVpVJyT
hOZ/Z7hvNA9J/zporCGduj+uhqV91Yl6XjMcTFDvQwXUMTcDA2ECQRe8IqWvzjbf
4iPWtbR7yYqoCv5kPtsTVX81kLYmhjf+vNUub5KlFB5vE1IR1kqMMhimv7SEbSBh
SOBAtXMHYHcSD6Y4i69j0gDzg6gh++tyGQROaCQfa9qXoTHOntBabi1zyU1ijUEM
CM6nP+YjHILRVCjyHS94mNqsZkUMj6/2mM4G5rNdpZef2M+Uhgpt2oSM5G20QkNp
aqiO2hXqqG/vEduSGv6iq6+Hy5Wu7K+cIMwyD4tdWb+RLad4d47VKiUQKPCTQPQ8
1kONl+tqsI4PRP2cpjjAhK+/uPgakwBNkqjeqsH85xo2alTektAjCAgPmcfYqm8V
UNXrY/4OANcqQNCWdqofFGYDkiTqCTdXIFIWckOgM8fZM1lIHm9cBe1xMr2ioBSi
Y4pbjsO6mMOVwj5G+i7FyDY/GNCfz9vtvTCIsi/QDXKzAdhIBUHKau+ZfFiDX0P0
VatRpqL2K2K47K/l51NkOzldbk/jSWaCvCBLdP0prAFH7K760W5ax2P29kjGxOo1
Jyw/km6mYx/fu1rNl5U7ZMG1mPUXiPR9Betifb8nC3+qQD3Y58qzFE8v6iwP42u3
xFpIpgtTSpWVen9BA0flmVGBP2WkgkT2up7unpuyNneLK8Dsmybkdxb8Mhyaanih
pXXBldElJlC9NYLZTojb2wzKRozXPMSvKvvIsCwd+DIZjW98b1otd4tDaWTAF68t
AtRrFCzcfATAvIsrLHgGyAIaVU/yyVgJ5qMIC73E+8fBbWhMtptrN8OVpTIMCGMn
e9fbpN3ZQSWbSTwfRWYRLLahFT85aSEVWrZXTh8kPYg/ewVB6KKnbJ+I3FLyid92
ByeebwRqzRZ29HVLEiqvY+ABZSaxvkkBV+P8j4rpfT7joALAAMS9AxlZnWLWL9xD
hREGyUfbUyawNIiM9oP8MUCSbd8EeZkccFHRsHb52Iv103ivMfYCA1mqzl0fa1vD
620roBUjg92gfRdfs2W2kvFZw9iBeO+DJLh+g5hXLuKJSM2vtYdHHnRSHREeu6DB
BYE8HY4IZyf/YKOk/twTb2TQgyiukXr4O+XZWmriowyBApgni4l4u4swQ4Wb/avF
/BUFp1K1BpvuzL7/K6FmFeZvJgNW/1bEvJnSz+Kuqi592zi0ovh6rPH7SUGXJ84d
La47d54C0Hil+6hRmK3j4PSsreTHGleX1Ud3xsJdwQ3CefJdVc5QT2LXT+UzYEuc
X17/FAZ5nO9dcOUbFhoQQlGs+1HO0wbRUBrPVTVyviDocdkHmx6jed13yECu7l/0
JV2zh3eSZEsWzygRUaa0l5/XCEKhcJvapU8X4gqOaSwi1HqdyGhWLMvIgSVH1vdw
nY9Fyq7beIh7pCiRvhGL3OBtMwtiOLAVazfh+TTJvneXHyNWN+5u7TgOPCdAYAsp
/ggtI/ap+IQUdEcHrmsTP8RR3fbNY3kT5n7yMLrp0adc6B8sxrGkB26IOpiIsDmX
xE3+qihW+kZxxb/wLu3bV0XTv2heBpGHAnPu38geI7H25yuKuSmTyya4rrS5NNTA
n/WeY1bGn9EpFlu4GdQ6oHSqRt7BvcP3RfEhziOXiAb+IfN/VybBp17rY5KxDLFB
F5XZFI0SDspSUJPOJfwTFsLBGZ8E20prnB8XJiM0PgbBccu/u+IM0sS93Gt3qBfi
hkcaLSAOMJPVAaSRsqeKSZ+d1rXFFGIytQfMC7g27RN2sKOberbxVVGws76z7Jxo
c/MkZkD5402UvlldTsunDncPeBLDBg/ccpruVNVQMGm+trlmG/rAz0jbvLmR6VGg
xwDttLEwgRH3gRfAnDnm3dY5dEuqkX3fzPwG8zOY03c1GCzPKR+VY4wLqBpYSIjM
Mr7FhwCgeEh4f+WCTLEcJWwTFdOzEGzaLeF7Z6H4xvgvVEL+eIIc4KL73GDP2tIG
3qJG7a8jlgk6jkXTOoTCqsGtlcJusWV+bjT/Vovla7Qo64BrmIbiDsVx8Uf4MW62
G6fikBov8uzpteDTVN3zwMCee+q0dTAhWbeo7bpiyt1Nor1eeB05PmMyHRHYBtpc
V9PlkEAsUApqSBQVANqoNRmcKfMdpq6xYTYhjBKA3SNBzp0UPXWsUOZoA283secL
KmEgE/KJhlh/djDkwmydqJ+CTig767k/3kYX65nSwlfI3+DFRUMzCH1n44SvRrrj
r87Il3ATVxk3qDtOtDXWE3uZq9P8c6z6fDcjXAWOOgVSzptfQ459ROnnHLyDThjv
/WEx31z7AY2hYTCaYmDUXYk+qbaBz+HpzFi2THdVsL49ZJj+DM6uFXtF8fapvYNb
r1yS3wtVCvHksAYX9R3YOLjGpbKZ/py1jLKuRuPzxyE0bP5I5dio2G0D2D7wTdf7
BCLffuLxmV+501+qXKzOg0j7ublaKwGJOqMGd5WReJ3dYS/hRy9430hAauunAlc0
Hso+55TPT0FnpImqIbnppgVzACi450LTfi1HQW7TamMLhnOnUxGBZBHT24vM68qH
RFOVSInFQk5nAZvjrtMzlZ1bJnbGY2Y8jsTvw1KQTUxtv2CHOXpdbjKIzntB1Wai
K9IUivXCtyYfsXfC39kJXGwkLlEmn0HlPj18m9Sb7P9VBaZpkIwfATXdSNjJCSCR
rIRU3g5XD+dEfDqcJlRXW91S2wQVy+OuMVBaBAunr/WzE6o8RNqHnxL5I95EyPgr
5K2VMCih7OVBpe04tyjQuWO+WiotUMzhIXrF7olkcEfa/51Hol/6ilG2l/lxqz4i
T9MgFxqQ0A0SsOX8fqLqYFQ/44VzAskQ8J4APN4tnXKdo6F0ryV+x2JASJQT8oq4
if9/kcMrznbH4FkWJs1CDsWa6rdSYjwhgzA01SjKF6odJ+xFRqCWcdbYMxIrPhw9
utoFGR7vOsJwEiVXSHR57H/V8jOos+MfZTh/Snen3d+UJ6Cv1uGA0NDh1ZZkW00A
XbRyKe+CPn0Ga5uUnbRxIKv7bEaBUQ1RbvN+Dvd9P1C3jdsRr1xfj3wlW6UCCaAO
sHqFBjdQqdXWRfhWLa8bsIKbIjx4G1l0N1IioKwhbDney6C7w9XbxD5BdzwiUNu6
B4hIhkPB30s8uZOW9a0yRkJY0d0ekHrVB2ctcUVMlq86gyq0laApDUITOEvKO1iT
imOlToTHJvqRnX5KAPAntxsx6LYQofoevMPEe/oYmetKzAadMwt1H1LctZEPggTk
5ZiE83vVRrrHQPqXvzJGKK2niflDDIhL2246SP1x+W/Ey7qWrjZl5ah1hQGhdNXI
6VJRxrr8xYcYXpMEwqzk6Xd5utMP8LO3K9zAfPotWxcm3EO1KR+aGOM+09jY6Rif
pyNRZ0TOAyfKxaomSnHEs5LX6qqc+FbFgzNFiaapB61VsN/drXP3fOYvIkIgWAed
BcLv+qWqXl8dLHV1KY0R9Z1OZb2rdvCwCo4woFhb83Rxxnw8uZQploa0MZjHWRG8
MpLJIfG5NmoC+R+kIbvFmfzPvUNrSzmY9BD1Vmgc+YGoAKLmRAEYIjIgtx1zbExr
QnwF546He/GBivzS1F/c+CaN1QostNWyCvQqA0Tz/d/En4jx3x8ds/V0NhhOAXly
FI3yQZuupnRoYRjmGSeQtGqSUxCvi989PODulK2osj9bjTXBcTpfvKrgai/4kaMD
iTidOCT/KorSb8N0+V6RvCIkwTSGK1T0I79GWKP9aWXI5CfsiWNVtDnouPqht+Fd
qg822pPBVEDXY/qfkx+AYY1rQUCUz2ezaIT0rpGHz1E17RqyLkg3M41FB6AxjtqL
M7naU4f45xAc1Xr4QD4Gle5jFbtUAuLLDbgXShJzqTKjezu8p4zfIOsuqH+ECmrz
68ouNpn62nurcK6G02zNdjDiZNS6I1C80fdZWXX7iIeMmhfmQDc2IYwnukST4bNE
qHfEIu4h8IcSCofUS81oYgLhBqIiC4NVQowyK+K1mf5gm9Jw2usSnZ/EMDX7cOaq
wfLE7b3QI6whnxuDA5LQ5XLYkCVhu+8w/larkG/iMCq6QLZKbGxsgSL755JkhZCi
8QkUGzLk+zQVa1kTGDWbli1ggNQ5R8R2k/74VSor9BKXCsuZOdAIsd/vYmrJ6/pr
ox/FMVV7xYgkXJpfKeNgGhc3+NGPN7fU+uer17YC5k/Mjwe0vneJIcEZcrqzHH1W
x6x/0ggMGeeQegwvuw76KPmfqw/RRIjQcR/XzlSkIx98ErsbOKRjCY3b2dUB69Ag
gKRLl/Zz7Diz/6RwK8AdhIWlc6eT4aVfdvQG305D96+tXxAJbr3Huo2cE0X9zPJk
eLdp6dtCqkwaCXf/N3XBzb+/rPOV85+wM9mkBaCecc1pPHhwa+imsoJBQquBFhsM
UBbDOiLi9yPKSsr17WPushybvgC9fki32QK/F0E6FOTJULdycPIqYzdtMfq3KAYf
6NXMj0KZ86bzcCTVGdHUdgq0lX0ZBD7RbenpsmruBpyTazvhtWh5PBhsZU6xb6Fz
qsXGJcTl0yBhVaX6/JTTVrCU9Jvs0k4Ylg3dCk3+ecu9r5nEgByVdR8Rb2sk/laZ
fm14YT7no48mQRrAARgmgHykBu+Bdjvd+TN5ARQzHNNXh73BqnlaNkHQ+qGe07eG
UjpWgBpspcDtsx5O/8NJUw0KdlYZozmp2cfizd92BxVtDyL+VOOdePTP1/nsT7hO
DPKmWEO8e/xeamz30ZHplhVllU8wcs+IDNXhqzLZeA6kmWJPS/gN16lmJzDFcYJB
QKr0S6no7eddL4TK5uqWgmBZbgpp+35+TkGEaQmizb5TbtncdEtQeZMfbHUgDYm0
1cCgVWpVyvHye+h+TWtq0mIVw0VcOY0mJsVW0G1q2GtcGbfy0uKZNSFVosDkZOw9
MlrKA9YG6M/BOky5q8IRMWv9GruuznXc87DEJiSgPOPndlekt02yw1Q0UtfMYnzp
LbpQ9ZtkrLCH6d2CH/NG4ZF12nb6BrFioFXJkLbtJWM9ZVhlHj4WmCShplMAq1lr
1H7Izp2PW85iWNR5zvJtt5k8rqhg3wTPZiS+iHVzf2kfiXPvt5xkc/V62+X2rNk2
lxxG0xXIpxif5bTGxImsz0d1I7XKZA36R6OTvmkFzy0YcS1rxKMSNs7fPbd8h8R9
5YdOALfw6BCtUG3J+YYZcqZfB/b5Y5oChW3JBM/tBvrEIu33nDvxaAKeiUOImK2a
qsu4889RmpD1eD4TzlOJnUQf7vHpSiZjiIVC0sisuhaOOm7ElxFHGnh9VgMRO2Qt
ybe/DOH9K8PzBbFooLHwxcBTYWcrk6j9cPecBSSKJqleTbMBlbaYISd5ihUZC4ZS
iOgY3+5L2u7NaQEU1IYQZkCIAIeYQumdPgVDWCtJBR3sAABF41vO1NZnX+Li57pR
/OZ1VGbp8OxadMho8oLeqlKihUt3zvRFDtec05/PCWtC30z3pBjIq7X10eqL368A
4uz8SyoKN3QmcHCHrLfRZD8A4OtrFy6vXwKnxwutNEwKUOo68DZc9EoM9jCBHglU
cngwm9AHVzslIcQEhKQPhPbKRRwOsKvhXgRmNLRnLxDeSEROZVe6scsXmZoTy9MD
UkfCcWyDNToxM6bEQ0nppH8WgxIoNR8fPFOSeXjsYkWuoKuYYGA8gFmPK4htW52W
zXi8WUKSu+AQNTuPlCtZ2CibyCAeBLtIpkOGdUEPVSJlQYMMmVNnYJ7Ntlnh9zPV
6UmYsJZqLofTQPOZHuS+Aq8tRNyJ2rIdl0b/Nx5FWl8/YE/rFTbqiO8jedx0h1lN
wKXdJ9WMvxQGBplGah15ywYteQWClGntw/9tRPSF6GZt6eu+RSm/N0vEsf0ym5Es
c2MWUIZ68lqa2XdoXaIe8CGsDpNqc4CpGvOmjZ+A3DG9T7krRTpaCM1/JwYCBJzw
gyfWfZfJxcihELh8xRx9X6nteCm0CJbXyUs6Pot0DU+Wt2l+4wXU9Tz75gZbycer
GAlv9YCQypMM8ed4EScpPsdNGr1+JVgQIzaeVsDdFCqWob2zWZz80bOSrlOQVaxc
X0VeH2b9v7H17LFiipSSQhp55ZP+OcF9uZO94VM3jzz8duzUYIPHSiXg88+sE5Sy
Z6JfgEd61suw7xefrZ2ATPFOLzddJgFXplvBOFwGvF4sO91hQbcZ1Jqc8r+o9DqN
4aeS/beUO9+9j4/qx9VpFWBJ04RfSrAv4rrvX0zxcGwLPgJ9CIKWRlAaxvHjLWvH
4CNpmEO77oiomaghLxFaChwPWcksKru0/SQ2vcKknbBq/h7Ry4LgREPFBV4SeE7N
2rysIsyF8Qm9aMuZQrEt3ZxF7FYs1PXqZQlz5qMgqvgBSEwdQ4sn+MjgFf0q2Qvi
kGAILftnbuiz1z4pGEKj/s6s3TgA2oVAsXdKc++W74I0pEUBzlZfAlEZWHicosK9
MhtB+dIn0Vo9DxXpqugvqdVsEMiC6qXm4U+/nlDNX2OImsT+53QBvViM5P2qeCqH
UiHN8CSOZnEA3eRmjrw1a4p6AH2SL8/Cn/wCKvDhmLrQoM6eW2vvMemTXLa+Sl1i
Nq2yiWOP/Z6N2JiLd1YvIEXyOFOyidRz5Nns6jh8jOzIufFLsHfilynVZxemWbPE
agXFoy9K/i2vr0yUVxMg//TzUKjMy0giJk7o1nb8aIkhG4z+T1hZPll2mW/akA1z
J/F16lN3G2DmIyCgD6m946JAO3uA4n94E/cAPRmkoC4la0bjEBZgx7odiuvcKAoQ
0MqQOXeuisiEfxKuyZtcsCyv/IzLdQZuDJZNBMdPCldTPDvF4U6YNs1ldBVas6Fr
JHac/ZEdwzUrVc+b73KNNaaKyGIbBdOW6DN9Wdck2wTJSad6PMpP6yyDwGbN6Tac
U4a3VDhGt7+Mzc4GCWmt1FLlbpTZp2f4/s5W4BwYndl5W1/jDVF0Pcu+eYcmSbnW
eZCrDTwT+QPBXRZ7JGCWfyfDPQ5cNaate/fFB6YvSw8Qty5LSNE+g+Vo0lw7HmpI
qCuARD9OXvmf1JVy6fF5mA/9mu+qXu96U8VZqdnN7cC6mxT5Dm7DVwG0xdyJs5lL
XNGrseZxxmBWI9bWCRMO8P3ipCstQJZRPv103Z/qfGD2R5X13jeFwEGzDEf6XVls
XgXRCYIkkNv8p7z6FAOroKZG2mPXULD8CepXMkRnjd6U1ISw6S7wNF4IPQYgQkOl
J26gWGAm0haa5+BJJWH3Sv4jCiDMntOEMbytm3a97ay6OHX3BnncU49xQwqzhuDa
MPX7QbyJ7bmAQM9KJrLj3YewWCfaTC2sw4sNQ+WAF91D4/JEhTMs62jsYJ4m3+N3
BsnSn2/nmQDtB+QyY5GVe6eCds7i8lcyFvEupny8OT4SLyYVDSv3TE3Q1a4Ykr93
TnYDb9jca6Ax/ZsWe7q6Zqic7rg4nijfH6mOgP75jvIheFFq2vLEvZjo4oIyJgpw
1hOLQCeg9zTT8hfvXijv4azbj3azs/hT6MVv27+TL7iP1luNh1fvO1bP9xsHhBaV
Iupypf6ZTojLh84N+Z0swnik+baTPRg4UqWSHhXB/k1t//VPDh4ErOdrcTiLa3Pp
+c9Z1T93GzaO84JzqYST2jplbUQeqjXPNRiFSgSKIlH3WMsQTQZWGmsuVdsYyT5C
lji+/ZtrMm1D/7MgFWcKNs9PxsPq6pEq0J6UUpMzQbwr2Dh0bx6KM/7xetAMrGmO
zb0I6tPDdlKv6H8/mJ6FTRYYTPlmB+XBhqCghN/cUbflP0cQC+4TByWxBrzEStzO
Uy5HKtnutWImd39F3fezelj0tAv3L4Th2cvnj9D8bLmEglefmq2S+FIOnufGhGg7
ynlMUKpcC4+zgIj+smN4tkLmQLbH+/hybyV7eXBqAMIeszqooI+Y2NoSz0XXEJnk
u+0n/+woBvEO0IybugQMFDJOZN2fJ18zd3l+zla6EkfDYzcnMln0Li0voEGwzS4L
ghcI1h84r3llTAwOfq2dbUnaF87hfxni9FQ/rvyZZwxsdIkG85e8WFH2U095PP1k
PGJkhKlFSpdbfud6VbQCwfhDFv1vbJwB/5/gyJiFMjiXInqDdKtQuJ56XTDB4ede
9To+KC8BKK5rzkQ81JxsQZKaFDCqRzkNg2HOaRWNRlHcCqgHvlvC3lul3eGZ5E2d
QDJ7tuHIsodMWF3M+yhnbzGg+v8abcYNbgGoek0PDvnXWvY7mkFVcC4Nxpfj0Jrr
uQCcR8nA6PAFpuA8G504K8b/gq1C3zixmFeoc9GFGjYM/qMgS6Kl0MhUkiKowDvg
P23AIE5u+x8NzjzPAA4Cp9zAKYZjLpmDXheb61KVxVKqXxWYIzF1SX0jlJapvDG3
ZBq/qBio8MNE7u8wMV5Vt6tF/CZ1Ifzgq01dPNXkbvTD4OA+I5mW2mtK74fuKgOx
OGq18Trw6MLLNGmOEjUAWHz5HRF+wYstFoNeW14vrMa5wO7gXZwQf3a54jImmPHY
9FqgVIhqIipyX4/p1CQgczL5u8oE0tYxVfXV2ctfVXhNLyXuq29X6AxW5Yw+ltOv
vvQzl7JvjRCYyoAO66MogL9EEYyjPCfAY82FfYJV2Jr5jrvhezuyVld4IiC94kX+
Eu1wjQ4Z4gQHcLGxyNTEkS1H4Mpkmwn8GZS9hPYKoa2vOWRrKgMtkf+4RwJx5tU3
AJ+Jt972qZX/0KwWYNRAvtnWiLiOrF8eITUSgHudoh/kXX/UcJvUSFPwW3rhffjY
4qbshyvPzRe4qIXul+Wlz5/luqxuiYtFB+Xd2W9ZasCbemV5gSBzLqm2oMGXvySK
rRPvxNj1PRpr7ArFnB6aOTOwGsDdurcgptCWWuCWmbqxPe0VMkU2qTyBE4RoA+xl
FXqy5hy4ralP43JLDWQkZ0fUhSFwlSgZYcU+anTO3Ydqjz9tnKgcmpoUCXRn++4z
dnxck/1WW8W4z4uzaxg65kDepW59/QL/DFslFl8fz/Aj3a9J0YUBgHLSlA522u4U
t3asGf1VAaxmYQIh3HQJk4tTI67mZy/vSBxKFEFmaObPMSx2dXzjDcW92IGas/RH
qQtWG0duXOAZtn06dWFiDpVL9yLa3w81nhEvMTAVkoDOYRff/zssca1c/qK1d6ZG
vRp9dfn2G4GguDKKz5FjImMXdjWI/UUosZveX+5gelxq1to2g699Xwj/GnbihIiz
6PRjndwpgmyqQfl4cbFf7YVyL1H8/Ofao4uKFgytTewvbyMHmhs8ZvxpEDlgEAdm
rueztX3h0o6pCvluHRXhzMtIndrf7azBbljREXpTX3+y+N98QYns1iLBRU+I16+6
zk6objmg0P9ygfa60X4Lw2CCH3jYlteHn3+X0/dMcwzH9tI4ndVPB7MJZ9oaTmLL
8bTXV6MVu7hYn85cPaOIU/PvjfXegkrGYlTi8W9vDZ1vRz3whkUmjlIiexAyf/Or
i7NKedCzb7QGTzM1fD3DvoxL6fJNGTMKSQuEUzvJvUluxOgVhv/Nm8c3edr0qYoS
f42CBwSGUcC/Kmi9Ga6X4qTu1JXjOKBLbF/OfOtsFuvmFojVSrBskXYbAzKKoXCT
aWT866G6P07W4mo5ttu3WfdVT+ZPRsdxQPR0x7h9zOP4rjucmCZ/x+D1vbTWnUn5
17wIRNzHKrCJoT/df2oP9+RsofiE5sJLMxSHmg0owss/sEFiZNNpplq4g8LtSwXa
0/deeYUTT3OOv4RW9Zhk89BNUWkS9uiS+xnNWQqFJa3fbm1KIe+iWY2xoS1x5lFm
PHCpD/Ials2e8k9yNsYVIJdIXLKoDaEdj67UvVmROYK087EhL+yfvh/gZvWuGd+u
FI1akwi+BQ9kvocEKbkH/TSCOISNeU9D52vOnKY9IESs4hK/JaFdE22VCEpWlJ3E
K0E7nZ+TFV7B5oyrX1+w6Xx8P5SyEoVLpBoYwwQlbU4GXtcOaA5ztziVbTkqJ5vz
+bwbOXW1zzlfyLL1H2twuLMnSB0pVvscO9gtE6h8JGofEFP+dpKuvxi908s/9+Cg
KPTu4XSsIci5OGomvd0gNg6oHD9OVSJ7/kCqklfGTMbP1K1O1dHsfaRg3hGgn1Dr
fondrdHjdH1yZrOSjO4mApJeP8rpxHpB9GsmTD2Ob0F8FP1jm95wwXds+jAte5Z6
HkaMi8y/5gvDldExHHol6/HbsLvn7Y/V2e6qroknX9N+oDsOiK0uCnxtzxR+Y8U1
C+75kLwALOCRF48rAPzHuo6uU+HqiTsbpwmalzhP8OGZ4rKkBndsqvVHLo2BkdnZ
ZsoDD4rDmPJm8uMtTvAfOfXBc3+6aQPb34kl6bG8NyYzqFnoj5NLSm0N+KBW5cXt
C75Yr7F+n97WRdTN9KIr68jv9RjGQKGugL/bjza+lo2nzVV7XlKuciKwsHd0KY9u
xymLZ+tms8LzodJsuGsTiJHkBkhcGr4gSSS9izRTDK9Tdj1Oj2vJ7ZQH1bbR8NO9
NdJN7vccHc+WttgE59z90KtMtsfP0H0LUuemNTG6hGQGuF/0wJqCZ8H+H8DUdKNR
BdiwgGpMMvvW0/Yzci1XdbR6VQ9j1Zlq30QTES3IH7BOn7H6jGARreN/L2m76XTt
lpssF9RKohSK1p5egz1O/m34zjX4JDg5tOeTi8TbCbjCrP/V9NnXtEZZ3KEb8WWd
PClcdoEgnSJ80DVgvixXEYRK9oD68QI1IY1X2dl/vh1TyjwoohsDgMHvJRjoRJGO
eBJU05rLzUmzDCLBBLzZbCylyMhW/XA9cLd65cCV5LzCqVH12JcfTJw+qr1hb1NA
DajwQyYe/YYqdY1kzkFf29a9eDVcEgYJ0ADT+NRURe+ftQJhmsWkHFboFLZFpCfO
ek6JSsiXir3XgMhvD32ZAib7+UNLEIHG3cKpmw/JHZWielwQKMmdyKihIL5XknJD
Fru8ufJGVk9JvT9m8nXxLw1zSq/XeTqRLbApieCBJU0z3u9NuPBh23V8CcgzPUBZ
sGZNADbDB2v0PuD5vCwhV2j4Yf2DdLQZemMyBdQZmWxybzLnRn/aHAtd1zRSULE9
klk3jjVocUkqJAYJp23HDGyjTFRes3/pz2raPK4LLL29mQnwCA1wr14sd3cU2AkG
jogpP2nyAQxosjyWOKOYMC9bBj3wqHhI8tbX1g3pFaLSyPp649H+EovmI0Z2mq/6
YibjmeihRPdTYcGT3/hFECKqG6vWmyRfDYmHt85bMIGrtCvvf1CV+jMXOHLp/aL0
CXkOKwi8N1rv1bt1dHQU/bKHZWaauda9jGoS80Fq/bUwMKnam6J74Qve0XxzukMA
Z3KpQqASvaqa7L22H27Okj6J3Vh9u5nkHQQ83jdlhBEzlEn4Q2alUTHwjfDs0liV
yoMyhsutd2WTLUn1kATrrtUJYoZq/4X/j6n36x1S4D6JASmz40EYy1YgQziri6kD
lnG36gyRqpfkEL3fFR4h1cTi3H3jLx1XorlhZOO0DdLfRh9l2BW9C4YV/PfNZprD
5lds+i49HydWpAuD6A3EB7k14OT8lIxB15CLl69tWVLh8A+XmOYp1N0w4FYNgSuX
ofYOtr7sFBeFyBS+TBs0/Fh1bpkOOGeCdzWzeEnyUQYqUOZZWKzi2njX9+SzGqfD
EYHy4LPoZXK3wku3rkv4XBAFbFZtZByqt/h5MZr85o14UzhSRFXRaxM0boQtK0J8
y+318ZSx0az7m6iap9v95SIAJeUb5h65T3fqSqF78KTZlUxlAvYSnhazi5fDI20k
z0E0CXI/sPYq9EOqKc1o5A/sZtXiRMgUHGkwwEzP9Z5RSP/KD4wII7wUPS5BFGJP
7fYaA+6fCwOKOos4HWsweqf1PX3o3c/YNB8BYyabhH9m/LES8Ifm4BAtVaE49mB4
YWiQ37B+mngQjUKLMPW/QdJLKEHKjTPja4yZTl93E0xveAvVqOEIi5q1fTDPZSId
u/ph7FAvJLYvqqiXiMWzS9sXcTnDFihayKSMeN9f/n4Zs0VjTQBgnZMwiGGVRaDj
zefbG1yBnN6iTz9g9J+lDdE9yBT+Yo6DWNWKFTXmcBogB3sorb+lPCarqaV1Pofs
cxY9yY6zGl+5zJ+GCrrKRb1IL0f1yMQGdOavvF0icE72UOs2WkPzL8IU4urK8chm
pMjSVRg545w7PNgko+i6UsChZf0HLdRwSrm1YKZYRJ35yZMBpNU8TdoHqbF7xYeU
mzEQvZhGDFUNyQ8cIhBs//2kjO3SueVMOwCrM1XaAeuYQW1qvqS1xMQIvVs/5BYr
6HthBwymNerDcyCoYM2LlxuZzm/nw9yMjEe+7XPgGhCUsABGaQ3RJCWswGu+p8U5
bDmiW0+XBmWh5yzLlOc3+QjuwKxmEo1FpK3HrHVBPj2jZdqMPNP77XVWXfUIZH2j
y1BcqoFzUUhl5VXNGdf233maXKRD5q3Dfat5iv+uFP95GY6E3Bd+fVwKbmfmpIMN
ZQKikO7wDJ2z2UoxTFY6sNLBsiQH5jx7H9nb+FKY+NlzB87bjbRKBc03R9wOqLsU
J3EXqnixMMMsY3QC1bVDMMICfMpeVWyTXsNwvjIQF24vVr+e68WwSkrSBMl1zI8G
688R7FZC80yfzDSoyjzTGUYnbnrPNbYPlnBB+YucyIA6q2CNHFYmvhyq2wCW2KFZ
+AiqZSw1vAXSkleZ5swf5XMzYD6fSnGSq0IGpbF/N17h+7HwCU+/9z6mxyQ8b/BQ
VXp6mAQgxeZJaB/4R5bPAG+7foQ2U0iwSElNFaKAdO6E6smysghspnubcySnPj7k
qYHT3g5xIo9ZjRtSal4GieKjCgGj7NmaW2aXy4nlGvmCmcNcQVcJ2rt6Qyu7vWU1
RizgXpLmweMiR7ViylM19witsiNwGRMDQ6abvxTD/CvAoicVx1JAUPScN704WL9T
vUxXXbmD3jnFIQ+cpm/bg98MVqWe3sXyOPL/ik9p1kSSmaScwiCFw5z4aGQaK0B6
DhiEIV86DUsQCEW0A55YoCcE1ROvBPgk6leR9EOhJlTgJ7D13N7zmpifaxJHNLcP
pj9cur4sjm1cOcbQPMOi6MnjiOxY3cIgDhDKUwW6A0jJQGURjRwjaPwTLEHm2xAa
guXj5+YK4hWMMnn8lT8+1uXM1g6qsftFDJTyxVrSRBJUDXiruMv6O8p90e6KAVLM
7j+fiS40jYyrK1HTKt35dXjsAbYRQ50BSG6O2xUmBj7ZWawgCFeVLLZ9ECuzflAM
OHxNpF689e1lG4MjLskLxzX9RqlDNDIpjZBIQs3MtlAmZ1O1ayq29ygS4OMJ/LLB
kIfWkIeWBe9y5BgeoN1HxgCHklj3HVOTOA5TmqK7nwzD7JcgR5oUJs56J5oqinXL
E10AzOGAr7N/Nc31/WmiupXrlcBIkiscPwBM15b0pbOzpsXGmgGzXwhzVaGHUqta
SqbrmyFR/2OQPVQ4s4MGf4JS/HwFtS+XNIRhXNyZJxm4aZ1WWKWtwva74YsFGZ+d
wXwO24T7zTsL/0Exj4VFmpuzYieEx8egUYq1nD/7yaJ0n4ErJ+hqDpTZM5QXtO64
RNQwUupB3RmQYaPWTGNMZe4kZ9L2VWJ72nSgNqsIu6fUOwCJORi8sLz6LFUnwJ/n
CJ6fNvFKJtL2eZxwDb/TDtxvKqeW28luD8DS9AmsHZumMr7Xp1yDaD+S4/73Y02v
Fxcol8g11+ZAFArgUG37ZfOOz8fV8ORYyZ/B+hDOWsMbPWajJKSToi7H8/uqwX/L
ziKJpNc7yxhxLs7OX4WAS3beGwwDljdn0AoQrTDRUf1Szc9fZxMWOugtnpZYZ/ih
dR7p3hpF64NaV7RY6cAKRkXrNwExMDcYJEceK0O0L5f6xDrSIbvmbGqDgJqOEWAh
4va0Rq+tnSgKj3qCAvyVCYXCcbUoNXZYictu1fg+J5M5+YCs/H0jP9DzM86Ks968
LmOdQ8NwQzlmMUOz6jTbYelvBN3nWlK6mhpz/tqSn5uPBN7J51E3jPD85KRcfxz0
bQmJw0Vhs3uF9+Nz/tMz8ccul/M/iKlhkOTjrVsNnSHBhY/yi9p9jx5oM6Gnn6Lt
bSyxuNHedGIEZ+ivTDrI5zpsPU4cpx831jhnbnf9DKQVb+g5MPwfjrfyvxFAZfLr
cC0JKK1mTQxNyja9tMda1+Ypq1hOHDLZUl5KByjeYBNtKu1uystxJGX5GFnr/cXa
CjB7feKYkMfP+HAZawB+qsYcbel/91mzB29+VjPe+vMpEYpsM4BX+oiuvCBUXz+w
s+nlxyiKZ7Gl1WUP8sbDIUBaQ416zmaH+nLu+hhlGPRoaOtEwhj+oTBZmXZvZ5AO
vC0Oo2YgpjYWD1fM84StvMkjKQLxOC3rg79p3WWQM51XLLBgpYEscyuakGsqhZ/6
t8Xg/JC8+O/kFyzfJt2yphW+UThR+AhNTUVzr5nbhT2PcSrt9bBc/KBX3IpCV+F8
cI45Yt9vVDUOsQ55WHvfTJgk8Tq9ES4NQ/fW8ep51LUs5GGU3RKfUQVVX5JC7WfR
W204pxEmx/YNXhIq7FsdwGO55gtUGTULN7DUhZaDIJxkf1DWEwrTksaA9H0B7+HZ
tikn7XgDTgSAb3c6rl1PoX4m1eEAkLyFV7eocHwZV58LmyQSLXxSbq8/X+NjLLom
ZTxqmYFc6TkCned3tH44ng2RWZj/bcC2Ns9+HjRpKiLw8imHU6AyZJlEO/fY+88e
DlakoYhtaOMVPD0r4kIh6fGPELV59sRaT0jwfiFPWViRIZTzrmSnmM+CToBxhRS0
cHHYopzGB7GwVtYdml3Qc7ELNSQDJjnQ76Ivmm067poEF3wcHey13J9YrzHqyRF/
EJHh5bMnDsyjPnGCpOP1pEDJbhxTndtYJ2Wt1FRScbeLDb1pBiTKGSt3xq5Vg6a3
wN8KqtWrFsGUNNhvp6cScL1QdhcvWpbf0d4zjjZiTwKK++hDI4lgt4JdwPDZ3qKZ
h0m1rGHFOaetWQmON4kKfBjN6BDQxOtnr43Sgp/BWjb1ThOD+ZdNqMnmOAJsXAaa
gX5spY1Ih7OFGfnSIb53a30yI1jNlw2xCbdOB8qlXG3Y+h5Jd4I/30RP7raODzZE
KQqD+XDuxmv65vGhf49+Bus3UAIHUTuTEROvzaMub8Uk+CICaML8AkU0i/lcgBsY
LjAtaympQdAifLtwAbeP0aU2BwEqcKWIZ3YRZ9cSmsyjwAvoyiitUiexPGTuRzqe
3LPL+7Cw6BtshRhy9HlEiv3zxmxmdcm9xvEmajsi2qyXBD2zJIHyJh4hdu0LFlj5
1n8wiznP+NFwy3AklAXCLhNvj+XYqqI4ew8FXxf30MiAvqJPjSoHatPcdaw78Pe0
aL+94jusf4GFwVK05K+upiLkdQpLROvz6QgEgUW+VkQuSgJjw6bp+VUAYHpGALDG
V1KNbeaixhqn3byd7yPWGfLqGvSFYmDD385BsywNrxJgqFNgvu54SZN7SyenASV3
gBuuM2m+QLYjmkJ4qolJeqc+rRpYs6paW7a9xdl3APSjZGOIGE5VYKUxP4VhbSaI
OJY6nCBwPWffg2JMa5deoi+z2FNq6QVgLqmTl/QB51oRF3N4uQ+Y5xKPRplIe0b0
/EgKJ1zX14WnDjPiAl3+uBZjNeDO61/r1hbx3ec4Ic3cnC0+ab8+WgJONWWL18UQ
Z/HCXUhxZT5DUv2F+ZQTKgJ9t3EANDjFHBoGktuskT5sjUX2GxscnJqeLrSEl+Eo
M8HRgUW8xmQAhK15qJXt2I2GL9gFlEhWghOyUp9NMwMCoRzCwvBPZfCHWG13hPEk
AJzI0WBGBjh/eDrTuMdQP/pOSPdYUkS90PbzyTk3Kdc1gycsqhhc5g6/D9X34HRL
+FUXYryfZbIkTx/aA9fXlJMldvoM3ZHUzzS2ZdlC7du5h4YdiWHseWdZofwkSe9m
H1eG2u4ul1+cwI+2/EaQVz8A2i5hEHh9hROjeamxuzXr7cjC/yqAgqWNLRReKwEw
kKyo4JduxG58tfO64c3VGtg3JmV+4sV+brDY0TcONKUCr11UoZie7TzIjCEU7WmY
VMw/AlugkHkrmUpSKNbOy1xp21CUnboVoeGMqYQdTCpPfWS8vmBvKN0dd6rb90+G
RsYqa0rtxtqNMc5Ld17t7rdbfB8YEJtVUeZAjV2k8455xBxfwhY7KNMN4+FgKtkL
Vl3p7A+WZ9Xw0yyQV46HqUzRINr6wtVZ1ySk/FrIVRaN6hJnr1/ev87VNHh5QqBP
3l5U2m24c/DLdiI0qRCNtYOTmCbFbutWvCFAzIu8UkLPPr/iwu9PvGEUCnpc9R37
PkS8mON3xPUqSqYrOgxJsRVnPaWISXj7uZ5JrMKLf7sIicTw+S4VE8ATxxJ0EXZ6
MBcHurE7xPsneXabKSrhBUt3saONhewOLrw6J+y/+IzuensU6rOaZ/uQqdLMoEuh
ImR3zPJctgzmJ28LeNDRWP/gSpKjB5NyPNdvAD5ngbCSkhGgfu7/SvuYIwsqH80F
3mEbB/aOJmmBd5nUVMoB/AhZqTqPuMYFkK6EDgGPCt/785g5WKuD2iGlbQ2NOBaw
c07qdD0thmig85mHFAKlgWAhssIZ5fvwwxbhpQ5N0O6dkHG8tP/qtaUqCSpdhH6h
uk1MSML9YjOYwYvLPChWn2OuhnbH9xVNcQ8RxgQuYx+wDtPgKCuMpBA4cxMm5XGd
HJ6qQV85FCkaMqBrfBgr+4gjBxbZRmCU6jvJp5W7dnfUTjW+qLTGadflzAqrOg0K
Uh7Jlzd/sp+FLOVlo72abg4nGSqJOS1gGK7h6CDJ1JT/2Gn9zyLHsAp6VsOlhMG7
mX8Twm9YyBGFCFU3s0MkuLlZKDXXPQZC+OZnZJ/VUr/uS9Xy0ps7ok4dvSuzIIkC
oRkX6b97UKoyK44+BBX436umZzXLaa0vz+mqXqUuEHss/mRSNW433IHfNrn9x53b
vGQiz99kaC0+5M85mLju9WldTWsUI9+mugID8kM7OsTWjxQ/rdihA2mnPLHHpZ2t
nvS9soQ+67fPYitu2bYEO0YB9KND8w1em8qd9YBPtV873i3lPHzJxOhF70yDxIp5
kChlaygNJFKfdl9xouDK1bpKXvLCTE8jdSA+v7y0SuiSWY/dAcwJH6FcHJ7B8Uwt
qCMwX53I9tPP5FNoPlK5yu4jbPdXPav9kshcLJZ689448NqIAKEwT1DNDiwU9ZAw
r4i38fdVqwKESPGmEyru4/1JxnFwHlX5TTouj5nJmgzP9KzVc9PY7UCPGwnP7Nsg
+GHr8lezn6aY7FYfIWn2wH/oZ+typOpFZHeu5AqABJ0I0QjiiqZDEJFT3VeSlsS2
D6zPzWq+8U0GSTxd4MqrRTegN4KZvS6uOq0iOFEOs983WonWgoP6buNTfCdtxAlJ
Q7GJV9eeOorVK4ubefvEAt8Qj5zvyNqY71y80Zoq9HAgvftjzOXdKnYQRM4UZ22G
GX+mEP5BqUM3zThkfq/IDINblKSYRaAKkjEXz6VUwXoqKtL8y+4Q61ToypZDNDbe
0jm8n4vPlcM6X3iMrgkEjOoHoEc+UjkljuQwP2klsQTzse4bcs0g2+9Ao2PSfw7k
z4wtDytYmMz/Zx2X12Dm7d9iNYYcRyExchI6CMPm1Vj7HG3hXD5jTk9fXrBNahJd
vwN/2qhxJBKURrSc1x8xZkUMAR2vcHWvuFqcxHMvNNqgv39jJrq9UUrgUYvufs/9
+16F/F4N0joXmNXc+to0FCPtCsixRKS94JBV2XW1k9e9Ou0jAeNI4r4dSuDqBHF9
xOb6wj/6yCtyCZYLkPErpbb+aVZxWx19MXm2VGU1CZVOzBSb1MhBeVsEBHEiukZx
jmzW3uJ9223zX31DRThg2s6Dt6AtnAOl98WORixaAub0RseE8E7+oN5wXmcqjyWs
VNt7KY2k1xioCgxPV/4pRrhM6AFVxah04miqiHbF4yWsp6OrxEr0CXkji32CXpmp
cao2c9SNDfEyBm12LDv8rH8jRbMBMuL+1L0aUFJCp8T8ri4cRt1iGLUrGh6LdXK2
ETpknra6xMvkiGA3eoykZTHd9fc44sFCRxKpkUO5Hb2gWD+1wtzUjFvdOST7KGtz
jXt5mmR1yFls+VIPdUcvTU58+SGJGj17KfNZ7f1Rw3vHJBfUbguRXjX6t8DsMI3Z
mvmb1KE/bKRlxt3zJkFRgHTZNlBckEnx3PvJdHZpgHS2TGsxtwBvcCjoHzFHrDJY
sRIaTnQvg1hfhwp5xBwUfWRFV7odyYvsysrW3g0+Sl6C6/8oxVV47kSXSvlAD8SM
NU07HeLpI1ggJE0IpkgRwssiN7bYFKQIjeq0ewfUbZLy5at+LzXVOZDnhO3iUx5u
bnHE8J9u5CDE6520fwWAm4ho+6/4SiEihsjHl7A5ZP+jVx/Vsn+bDUQirTuFDjwF
/R+mOi6fVJ2uuJYRJv1r6vOVYCtfT1EXn1XRlywDoPk4rXAm9pohgE8BUF8G43jv
bvA+qASjJHzvURuk8aRn9gjKWx+gvzSTR1T2tchaoo9lYkb/dmCCbt6/liwl05bf
kIv1xLzIIlVMgblB4j9+EnTCpu653VWsvVqj2AgyYk51zhy/2fUBPFnSJJGwOxhE
VNIvbU08lefYtvZN7AcWINLJBj/ftKRjksoyhOji/9FxVV8vxp2FRPRNCp3wxzm8
2/BxdmmjJfj3QLvNc5oCDO/CDRLbPPU/6OaJCqZXDT4CaxgUk2k7kUaZKyGNVjSe
wDRQw/nHGFelbo4CBPh78U0lEBWPGmUZWms78jJjvJJg8DkX3KH7yqMcA/vqfPur
vgcxx8yZkOUkHMokdqyceSh52BxhRl/oT73Je4q9wuDZAHb1Qv7EUyR/LV6yUsK5
eF9Y+7SHRGpldntuFE23iK1Bj0gFdCLgM5ncx7/NfVqntmBrGXEfsj+81p+sfih8
18kCejh0v5J86iWkpvdz4QThIFNQnsgulpCWtlz3TJTkjTLqNb7gIqR9E2aOa3BY
EaBbaXNKWSW+1paOHr8z7yWHDkA0aDpXRlPxJfHOpsKq8oizVJ2P/O7PV+ueT23J
iyt5d54hSqn0zLrAw+gPSc1q0qm1nlVYBVZuwmCJMyVTz8MDs5Df39V5SFRNfLey
uhTAAaPTHTsqblHoCA7NSloS+0iDI5dE2BNfEAhQUft1I5d80antM248+wFgPv/I
H4izmvaFrtSVmoXw2JChE0bvBhPU8od1FJhv0i5rOv9NRFhLNvWs5KvCM+/XSPO6
jzNby4HsW0A/pUZmGNMNiA+5NN25sfQoAeIlZz8qVYQ6C6uBX9ZLq4z6g/wPNwP1
HBiLwVNtzT4a7qJfuUYz+Bh4eteoddUyIrwEx7fssFDBnR+15ak893mA2TKs/bzm
nlm1++fnUVYNayKD8QgU0lgSvnYqYlnLOokrmALiD35uFgWZMcWQNr3ltTDsQwyo
Hb8BBRDwSVZ7NI60jct5K5UIXmNI9MMVADJH9sDamKwIGOa/cpB/3pCX/mMYEq4o
PFYUhoGR90yPVkmnsKxxUdGxRa5NbDgn0O8hiBV6pr+zx9xt8ocmLhgh5sAbMtYb
cKdl/A4ePRX0RCGR4yhI0Pi+gAJq2qvmuB4C9TWzo2Rz2TUaQe0gxwHxXEksrXe3
E9foz9rHP0wcgcm9PtH9GU5ChqUEOY//ABrMAjKqLsLPciUP8amVsfHiSFBYBKSb
PrbYHD/I4x4D2ob8bZ0ZgVGcfiasXrD7yW/R3X4oGk68nJIBQ19/WZo9xiB9ujJN
wAzYyPjQvENCwuWjuZhWTvOieIu9U7mFBK74dZ+TFc/YOPVkmiR7lRHontyxIlMJ
PlrDbyn7qF86RKz2xJOthMC0+QooD2KhPtsJr8m2QPoBCcS09Suqd8jRx8y4RkTW
LyKcfQT0EWGYCSf6M/8uouzyPGdowk6O74XCatasMi4OoGAje6SrncJdX2X8AQV1
BYUghPH056o/e45CV6S7x/tys1WSs2mwfw0gluEgchcItCtnBoHtpDVKnvEmhu2T
qAjrdUubEIp7ScDSA9/61qFncOJCQRci3Nz9QK7xqk2XcJBWTsW1HaTm4nKeDrlX
gPNnybHMEcHNHv15fm9nWomav6O+6m9Et916ZPBUrR7yBneSs9Ob8Xb9kU3t+TU6
g2EWSx4MHJMB6W+uJqPkToqazgMhSA64nEurr7lq44VKJTwlOwXwbZjvCBsJ2/ji
kZMfVQfFWD0CqWszq0vnNVRybUbTOThvx0CfSIrnJCbl1cXuJZ4ME7J+FgchhW6H
cCjPlk+sTtcH+CdQPLk6I4WlAvHWZs/FM7ARTWJoCCA/n22JxOcyxsb3G7BRQEcT
FQnrWFWd/6MV38vOH098OFinZMLghr2nXnfMRPuwVDAnEOZLqXSY0MsJXtKztjlL
4vzvpnq+ZfEqqqiGNpw8evKU3zAimXASTy2X59ilixUMbOg6nQWZs0jAg0GgRxCx
OJVYzZDzuXm+BoiksUSWGdX+G1rZpk5nQA91l9aOOrBpiehESiglZMKjr9Xe3FK7
/TuOs21nRwBjnsYu+mM9vqq0Y/11+dXpUrVTdraQ+5cGMMGpUlwKkeKqH5uQmIg8
4iv8TzJPl4p2kAJgvxzhmV2wlHSOmNSb26ajPc7L2INs8XR+cafQWuS4icpBlv05
X7NDC8VMQTZnmgxt7NkuuTZQlVu+hcGd4Gys4M4qulXLHB1qFQ7xmOSV2UGDcRMx
CwVPRJsiI23TOVwYt/BcwadKZydoo0uAFysHx8wIoZ6P2+bjpJhofrq1R2yoyAog
9DXXWq+15dnpHfIhARcqDOy2417bOMm2+v1rgp8uK/owaCR31Vw/ghlDuAjLfXCb
9HQWmlsftdq9CZhijTliw31bmFlvLLpDdwkW8Un0LDnBEAWKbQcFyweX98EitRrV
Wl/Wm1IfKRVzcJfMmTtXLzSKR02uzXkezdq+bGGLzv20jrqaVPFkz0p9xnQ7R0Z5
5euNegTi0i4rGPdozuhSDZURNIpH2Xnc/vLO8TXw3JXZ9i3i0c/N+2LsXhUOLSJU
yJ1xv5nC5S3gYa0RjWJ7cEefP7tWM1cGUrJpqtwLU3VPQEm52hU5me6ON8FBynW3
lv64fJG+Kqp41QeyRauPinkzzWni9ZkK5jPpL2BTj6qGFYGnNZI512oItzklDgz+
yokIJgFwhhubkwf2LcUsRjDD/TzaA7Dsm70UWOCxCAAh2Gb+N45b/nv4mnbSfj4I
vAGCqf0OQ12Kbrk9TNZP90TejRfZHlsaMzpl3pS5Z/X42xJwPpi67mIMMJmm9Bzm
7Kzbi2FvKnUYdgV8nX8R/X3GZE+AjEaGOPJM6J3+MyliKB9eGF0q830L8C5Jo5lR
V2BHsilrhhvtTCkSYzQ4FxrQju6cfQ+jdjQHYE2A1gMpRAXK2nMJTTAoLyA15d0t
wicyuU4IbfxueCpszPAvpraDp54ssfJrwW7Y3m5fxjmONuoEM2j/vOQyn2x+Jun0
eUbK6Dm4kWagjNARPSKDwGNoWZUAovjmGkWLv0Qs53lMBZDVX8UpPtMK0DNAeDOB
Dk7/14wNc1andCR5EUCMCZ2VAnxZfwgDIcGqZ75n/n6NSQE1Og3oMI1X0JVvrMvJ
gNRoDnFw/C9AapuNoRxvKrGZf+MYxqw0upDEFK1cbiKZZk8bZ265clRzP0GbLRr3
vMpxBzqhx2t7RI6Yqux6V+Bz50lcI9waTshkEZ4LAeDsglSTH4xI8BrsJRSN+U7Q
qsglZaaRiJwgIak4Xx4J9mx+DinzcVxuJTWUgDBQzFM6h9uISSZY7LbU8TFzIe2D
UDQuMAHk9NFSnuLnro/S0zLATXcN2YJ0TAUUMD4gW9n8c44sRBH24thpRlhAFa6N
LCnCYuBokaLafTFIwcrLZjn9izYr5up5oxkgLhR0+cxC7I5vVZjDAI8QONSUkQcX
R4tPkGdjmkPbPzTdVo7xxI5ycqmetlJFXUVMMUgxrOeVh25sUc4GHrCWPy06jZ1C
vR0mczPHyJDeyvPl0gnQ6DHoytN82pNfoWaZxQGCa/HjE7tEo0DLhinjlIgX+Piq
dPHh7WO1j/AcHHrNes8vlIOPyWocSu6/36KUuB2An1zsnbHABecEaqNfRISLsRb2
QwB21LIjsC0K8CFKb4Dxm3yo5/+Zmg3EyApSwLdbzqevsM4SbdEnHcCOnittHuPp
oOEzsqcVTF73WkIT/N9j6FburXp7IDPvM+iw3FiiX1zlZK6t/tUvAvrCl3KJdvhf
puJVx0Q+3EFcGeINlobN9KMitmbOPX6U+9qa7PzrOL57JQ5GQJNXsAkdK84vHld7
l//AqgYGzf076Da8s6woKIfZTSQlSEmK3AZacJklry5WdHNp+R8bvokf6Z6E6amd
PN8AseUJoE27q42dcLXSWFHyCpetJF0iJUwhGfUQ2vQAXjSJ0KlWZPADsktf2nHM
vfrtbVuGO9eBbO6/N+VIhL/EOjPw2gWs3OpTFbvVw9HQjwVKXRPW3BBTnZWkNbJJ
LmxD8B5hnqIgUdvkAYeItgK4rjT6cslaCagT4FwJ1U5XU4JuJKcYUXPFzZcWBIzJ
hqAKGUskYFdiV6zs0DIj+pKwMuwN8MfTtxkYHAr3cvNXjQZlMUwwSISuTjjfjQEq
x2YYN1xW0spjvHJof0Z3w/dsaawKMd0a7ZsUIcGQk8Vm6o/7kdaSKf/Ibcbz5AzI
f/5uJrfIkuCmo2x7caX0oTGyO8w62fdXXdDJeOZJ4nW+50olIpUKk+xo0s9dN9bH
Q2eIQAcy3yz2S0d4BA0cjwEkJF8nQwztWJjw8iNAejK/P3ZAR/23mxTuaM9CI3v9
ayLBxiG5zwe1weflUIvK4ZhAWB79YrgkrZ9owH2ufSD+tSc3Rg6UcZCC5JYh3DBx
Agm9dYv3su6+qdRug0Zr2rUiYqsrAuG0ddfuW801cS/kBW5BSuI9yG367vEQK8me
PueERqVaGl8FLsX626v1q8mSXvDsQtuU6GQHQVvJsEGJECLDE67Bfl4GLUpBtxr9
T2+rB8P+42iaQu5BcFyhCTSmDwqldfsFtzltAGf2i7DmwFyk7XrcUAGehH8tfYKu
FYIQ2MDtM+rpfYd1d2PSt1X/CI1o290fUsa/+H34Gs6D/V0H4Fv6QrVzjnU4wMXb
fcxui8duS7QW5tC7ndh0CWrpd/VgSQprk835EojVhLc2LlbeerZHDx+7OdHr8VNC
cg5I+8cy/mN4T1GbSU1NUNaOE838vIJrs7ymcrbnwswfx1byJSkiWf4D4OU6axwA
72uP+1ueooQ9SsogST0VB6t+Qv3zbfsO9oZTL1oS6Z80r7mpCWqoPWx6K7+p2x+u
RBY5QaBvjkFwrn07BE8X+Ad6gB6xRInMqy873x+Rz8MmweBSCO0vlaIK28Gnb0q2
+DNfBLo3fKlsY65U37d6YAmQ/VNfyqPh1rnLRY74bD/6AAgPEbsK6Jb4hAmxBX5A
UTGD03uZbJ6Ymg5bHSog58qfRw9YmZFVqJ8lxyct5Vg024CEHrdJV9uog56uVRTY
rnJYcA30kcfkTJGNE+fHhLwWjorhyEP1XMaK22rF03DkXrbk2ODYmXSsf97BfL7u
sy+tVqC8gWGWsvnWe+rWRijJ/bLAJdVamCvtRTb2DgAFGCzhv3YQz4CgYHCFumSf
llV4TUyMPjWBNVo5UrtyLRFdPkylWK8QLKYKy2ljkQkSIdO+yi9OHhxcZYDslwWx
f6IjydTv1WbQuuKOfE1bUKEHeVEMNBSUe5HD6tpmz/PEBPQa18ch5AwO7sRt90qq
Xg89xgO0Amxp30vKrAQM+n+HNNZffjgbNG39s9CE9wpYn/a/1MpS9sYUmqlxYsL4
FQNxzHc6fSqp9NGEk1Dgj2FI8HoUTTBelt/BqGG9ZQRTCsFDAeLlgjNmrKS4FLzY
F7WFtGsogquMmnI4YsJ2iMeA4de928mR7SJKg6mXvOmDc+9esiEdDd3QGqHfS6LD
ADC6eQtguW7CNpgBAYfOKt1OK58FBg+BMG8LNOzhc7FqbnonopihedYIDCDxyq3H
vSJVOV5O+I+An1B+5JaWoLUfJR6rJLKrxvwrbx54+BC6VDzYRqqtQVsYl0JkDIvE
Oam4IkxAT55H4xH6x7/0psF4BqLQGRHhApr7hycJ73+/kGRgVlwdU+0K5Fe2egXr
3AFP67LkKMRc1ZUzGK4PX1InabDboyTQjftQ/7Xqs/jCwpfIl9rnixOW1Fwg1fDJ
OHGNDO6OSuWLVnlXOCAzoR0smr6SqRlqbg65LJPU1qTMy9MBt1RdbAU6SddGX+Kf
1BouHQeASjWO+uKdEys0wSGpuz+yROgd7awkOZXsPaxhQM6zWIUs4aQA4wH0WCA4
y5rgIdTtZnlaM+oNmZLaUQ1Wf54CPFMKpMcshg1Tz07B5XEH3tqbUc2MoYXdHIsy
Mfif8DDosBbj6vcUQoFyKWsTw0uw7yJvjzchnY8tnaITp0+CPXHjZTiu1QqJ4GJ7
DDrAqIY5eBMubDcsK/faT5eCSuU3wQZ79WwjhQhlkmPOhcGpUFHXVPLvajWlsBJn
0UFpUVONz5EAI2HmtzAi1IlgKzfAD8nDtEnG8rJ6+Nl/aAoRsaarCtGtJBytB/wJ
gCBaJ3K9wob4znUhPPsaHHYAnhxoDE7UC3DdcHh7cIDBMAKSHXnpbGxQuxNT/U8G
liqAzxVIwx3zbxRgWDm9AxcqbiyIZGI21EJwzgToNF6OLewI0XpZpkpAIW0CLn6z
1traUWnuuHWhvcOVkndz7la0Dk/qTxqBYueP90+nD3BdSwJGzgxFq/DJNxhzZSP8
PeM4bbU3AxOpJyl0wO2ctQWTXvSioZdf+yzL9IEIUDmctAvQraI1n5n/joREQU65
CvG+4aHRjJZSiP6+8VQfuRdDJyfYeGjWBSb2CRTtZOCpwCnQNvYRvLMwrlIHTCTB
YIoAr4CsKylARRGLiwwJgRnvb4otkBV7ohTI61h1XJgHIw+Jz0rV4sAkl18aZ/b1
Wo6Ue4RB4J81lBzjhkILCB1OYKFZG/hS12oasi7IM9UOEc2jI3c0qutvtrqd0v17
/neYFEoaQDkG0dDclCYi9lpw1SPwmgWeYjolJ7fpQGqvwuZy/Vb9rKm3Dz19phfh
tBC5HYusrxGFrCEfcRWCKEKw8ZMQ7iusmxGgXkT7KafbY+fsm17A9SzSmjkFt/+G
3kqdPQdo6KMkj4nQ7e/DwI2G7vZA1G6S/+tfg2sVkSwPX2/OCoeaaLYRnCWIlnrV
XLMPPxvIVIQni+BqhiVpz7XO7cBnOEUnmf0MpC8jn67ErGArzGQUvCM4s2fbLKiB
GsCqMVVcRg2Ppvvj9EaHPlyH1KD+/uW5wdM+l5JtAklErZfh35pHshUmwFrB4t9a
mlvpYlrVKyASdBe9OaI2oXJnYUAX1NqAcEKQpMvZG1YzXwmSAsbZdHxh+iOwIDez
2IH4Mt9enHHRNTYMrg0gLVUo6gy2MUtx+/tpBosHuwugc7bHb1AJO1zAgQCD6BYO
UX/oWj+X36KzVwzpEnTQohKz6slTbT5stWHk0e5pLQjb/R+YpJuQTmkdx1mYSoRi
3aOt/Fz7Lf98AE2Lab1Tf6alwtqZVrPmo7Oh1EEArvzvhrj+xJCXBpQxAjqBc1jf
ywVH9+d8fNITBSaJU5pd8ks63fcsz1cg+rHotUgf4g1CEFQyz2SUaMspdxFE8UH0
jeh6wtmCj5FFWlbzLx2C/t/iv8iozjsZOhbJuP42DuKwPoF8oxZA3ouUoMc7aRcm
Gy7jV3s4xjrdzabyblKiVeSY17a2+dCSHzCVjOiyVWgY8rdHRdBNwA5bg2R/it9e
hxh6pfmHMqIPFqjFUBnGFtvkM6CN/Nx7j5u74CHaKbME4g3uKe358ZItza/KK8k8
3c9/9oX5aVzKjodOXXxte/gegzqSVDnq41OkqH0r5/VVvX4ScEqlpDzhwPqP2pwi
4UksnURN90UPFeeJhRgLFf8ihgIZjDMEQawgoDmSmdDyzxmDX6Vsk4T9+UxWL6Lb
vZQIRN5dRHC1NDs+v4dg7nljF4nCHMy7axsmiULwMbf1wHxmb7/zzKMZSLOl1gNq
1z2llb12dgsJYZbA605vDrghPgVLmhqidXAbhYfqv3ZIuuBkOXBM6mn/S8hXGREI
f4MGkMrwZjTf9cMmGxjjiSzoo3V+7PY49sz5gj506SIO/F6dMuqGaP5EFepTDU5B
uH7f0ADDtobPSPFAznY452zQjtkdyD3foL3Pfksvipu8Rl+K9SpB2h7gabGfW5bZ
2fIhhmCYpV/KwLOW5Sk1wOCpoke4EnLr6jEKN05cyXFkbRXj86JriyUFrRjjrluO
gYR/9iRjR/ecc1XXGfQZEIpyGpyKwsK1G1VYBua8zAgqv79gBTXFX9iELXsv+rRn
dqT1ThAGVf5Njs2J5qo1rHc2FqvIo1r4t+NGdzVuWAcGNtiXZVu6xc6180+/byQi
n/t4xESnU9p9MIalV1wc9S9cdV7A5CIQVb30DoZlJyH4usiCoT5Mj32PgSmqzKp1
W9RaRG33iRqrcl1mzEsTBZmNtiqJXfwOteXFtocd+IWwmcPKVMO1nKLpFzFywVh1
+F35YLzdlzQG2tq71RldjaIyX7fZ2kjllsptqrIZ4JZJRWhi5C7CprfBEiN3ksQj
y8fmj+wGI2PpJBc8oWYqbc7v+QnXaEow57XGcw8x1XAU6PSkiLsY8hxir7QZmbtj
0RSTDDGSARM3wT+n+aJVaxXY7KduQT0/J5BYXFnleavEK7URq3gr69dPuPOze5nM
61ACaf9oPBJsaMJra153xbqKA2H3vHbhS+S7FBhoVyTPFrxJUoFITHRz3E8AX4/d
wmxfrvZzCYj0zTmdeiEfshc9S0bOGXl0NjJ3hxzUXdCEKy5F/32JDX3kB2OsYzWg
C5DmZiQAO9wYerQfpd7ieUAW8YrH7UbpDtkkPq9smwy0NU4tj6rwrUb4t/2oijom
yxEo2lOyiul6E8tZ0kByRe2JiC9SIKESYtcBJgIcm7UOrF2LaOaWfUz/Xefw0GQ+
bPEODFHW7on74NAk9XHZFkuy5IQp3ssGGZxzqaRoNilNxfP6C+ElXSLMEL0xadQ8
5OsbVTbk8wno221sYVG7It2EQnBnz1F7eR4ucPbTKhIBP+20uy+yl6MarXrKe79T
nF0mvU0ej0kal6kJ/NyFHbAp1V/x6tEewr/8WV2avShP7v7z40I6lTmW4oJ8aSxC
FeDPI8mklo5PliHYamEIk/pcM0pXW4xiLzEsK3vBNCM0gzzaxBERzYH7ytJqErWE
sO6nc98cdpfPpAzv8zra9VvN/o9vGaoxiBCCIrjqsppXI0JzsJYW2y9t7fRvsssJ
sGErM29kG5yVYJ7Pnz9OUAkJsxf9XRk0dQj/5oVKYrAFDnSOG0uo+IslCkKVN+yL
VFm30KVQL/Q7DWoNMgAjzch05EWyzDN6w6xgKk59HwQBr61tA4oETBK7EJ1SK1bx
dqQWi0jYqMvJ/zQx4+D8AL8DIvCKwM9hT/D7YSWx2b5X9NB2SUfnLnIkUcTrFdgn
ikBcr00Z8NKfO3+FQU0oPX0aSpTlXXxmzz0zR7nCfXuuO71z+D1x42GFmk30PbyW
GQcgZuwyVkU8DWOjzUEugenxQ5A6lNwLAoHry/GqZJ3aDHu2bGmeTLzoBlj0DclG
iKCrY4jRovauEq5aJES7amXuK+A2teweV1FKX1Z1IVfZYv8ylan78dmFy+hFNhW3
gbHZfoBJwH10vdKfPTap+xwvwigPd0pXwrlEvquYMX+KoqycxEKUOVXOJ466BsIz
NbI3ZkLFmjAHPUdvRdWWMHH5k7UCJV/vylKIootu6kFBo97JE5Itc1pwnQ1B1YiT
iFaAh5x2jRA9YNQthq6mJXnTveNN/8xG7fiaLaTKr/r9r4obLyu5C1j3Ubu9Jwmi
ezV7U4Ta/iIn6Yf1bGDNNMvINaP6nmBpTNEIqbmawLheVUQJoh6mP6sPgJvcO6Xu
CMDpFCFnI5Uq5xXHzKK5PS+V6Ge5gi4InbR3ilL13b/wxrGThD3hpSdNSjXeSm/O
W2YIEvXl4smFNXsUhl85d/TsD2iAmQ4mwkAI4WXjuebAgiIDISlf2QG9Bbcg4Y07
i21kiuqgdgbEcRhGm+KxZSehSaF6WLk+iD4P8kxRjv6z2hegCRc2KdUvZGsN9HQF
9uspy6wwPZqsLltW1OXCmaMgeS6xkFJAcQFg8CEHlFX0fZ/XqJAArhAw8iQnL4fa
QHpMkXM1Rq0SQmwwJIGQrg9fzbMmQpx6Y0sUAeriScbCokmcuR1I/vjM7QtMK1Op
CK+UJpUwzwSOoCc+aAqmdXEhFzFeCyqm5wHx3M0dNyylIxzDV2X4DwnJpMyfPfS5
2WotvM9qZP4SrDWzcsd+YaUrx1y2wSWGMhK8En7TakIXxsnjAZKT1zPITDCkBTQ/
2PZN3MvHMdMuCiSV6HTJhZ+9Nl6ytZmn9DPc8yIvzF7Fuw/zsjD3m1MsO7AVsCbS
4BBgyPsZZ8n9l38eQH/o8f+6oybqby+jVZEiFoolqng+hv7T7T52Ic3mVy8jHJ8a
Ak08HfiKhMXTI0V/723I85U6dFnNRpdNH5D1RR1j9jEfb9QxW+bdSA0FBXC4+cJM
ARzTXdSKsQ87ran6cwafXrk3CVanFxC1J7C4QOdxcI9UX66wbSrPn9FK2Cg8jcLw
6YtgPNNneYHdTk7QK1RvJYrcmXcqe3WeU/y45Jvk0U2YvxohfkO6bMK5P0LlvZqj
EuMlsIaAnLZ/+PRy5tfrlKLlYB6AHmSEUDzK/OoLu3H9uNjUVz/wySuWm9bdmnzG
dr1OGycXauxUIXA/n6kqm+y0bt1YD+NlShrdHMnYp/xKlrmOAnmko0ThI/WPvCv1
jaEawerB+oKZXgfyAK/cQXceBRN5SyUyiog16HWqY1AhGMvJTigWZ4TTLbRuF9Pg
CA5rI22732ib4YL6c8UXsAhVvpznA2bG4MZ1Aik64CuS+7ciCQnoK34OQTSmlla6
f78Iy7pRj9wut4sODbGb0QwJUmW3Q2oDV2S3FY4D3Zm3vAz3/kln6/lobiF/6DXl
AWG7cNgyc9//oK29bNMHRFWBK51r8jbo/bMbnzApLiouXjSPGbDFporEgoHCUlWt
kr3p1wqM8xwAzxrMU8Yb2K3wYTUgGm1ylLNjz+kMSAEitXbVSW+eop5OKxN4fnrg
o4QVIIOIpZ1ZUQ5ZSG8gZX8rSnA4g4mZ2jodDCojIXLS4PA5mIlEGy/JvLh//BeK
O8e85MY0lpxf6L459eZuRDufBvE9kJMr499Ht5LB4DgPN5yEv60TcE+aLrqLZmt6
zue9tP/Lyt1ixZn3Ae5zivvK6BTPgLPdX8k9JChqkS7ibPAi+ZIeSD+Tgx8Tt3KH
SAjRJ4/8beqxLtCKq8DiLJTambOmLz6TB+CTCsmC/fOU+QR30t8VC9G3k2Sx3HHu
MtiINQrVAqPpKcthbka0H9z+y/u9HV1TiEHTv3kCyN1wy3uwnFoQTLxHa4zxafvM
7m/fO7WUhpTlqvWZKBZATbgq/5Rfkog9Dk942gYu4mrlZKcenqhtkzmUFuIH+I6Q
kIv9c/2fBtozabrIb24jYlvG4DSUdLI1AayoNIRFkAqWiFMZb4QlHR9con8z+SsB
M5C0g9SHUxUNDPEiqeB8crjouaaCYXgujyrYh/F4fO0ITWaWPTw52eLIZl+lYJCY
d9jltA6yxaYYJDav7xSDbq4wSmJCYBhbWFaBmftKXer2HirAU2UEb08Wwnoo8Gxq
WIUIWTeCYwcrNIIX/Gsw0YxcCkwxvH2XlvXOjifqbbFSn3KufX4kytvH+X7dnqpc
sGl+d9PZ5U05Uh7bIhnVVL4n57CwHQwQzEBcps6pQWdVY0VKMjiRVgZAPbVIox1s
gFKuNo+WxAeRfKBeUi8rcd2N1i5g0tNqMM/l/J/GSflL4BQ4NtE4FiS8l1sJYYdE
NQyCsifUHpphX4U498WluWcr2Ny6GcH/ukugpYP3tqzLH+W9TD0m6g0zRuMmDktp
LVDdVShT0b5lcxdRhswkGcuUGsfYjle7bE+e++4MZVZzowLp6QdjxY3EpIM3QD5i
5irkygb/ZTyKPGZKNpiyqz8P8hKpGoACnTTWGDcoCs8Wzyp8v2sxQtpNINtENZpG
qT0/NVZFCvF6zBGZLJoqhyF3W3pWfdsnqJEIg4468ILRroylGajI9rPEDaAFTd41
msXN5jbHF3hm2wyu597kKrqzNAd2geQEvQzqjW9N3df7zlLDwXO9MbOEv6E6dazb
TernfWscYthpAP8nGzXEWDHuGxiJgPo2/K5DFgciqIXH3G8vJliHkF+jToW2FSFC
HXC1bBk4n/7h0HshFrdu3JFgfdZ+9VCnPWyJLj3tzvV0+8nulvWGv+0c7gpC9iRg
OqdbtK4fsArSW9MDFHlpEnfMcYEeGNlJrMB+T+1Mg1SEJtPWj89jIgA7Xf7Po2Km
AR4a4Wn9OB/xYXsxeO+L4pt0Mdg1Y1PsqknKsM/iU9wLqWnAgEZVEjRwoGDwpF7o
zSpffVsl4/b7oE65Ty7PoQ3t4SkAzojk3k1ui123pGbJRLlmhJud37sJaY2MD/an
F2Srs3cFzKtT/vfoyRrgQZRTCl4noPsY4Ms8/d0GEwSadtXQqoLYiVSI37FbJZeO
Lsh+NmLngBgPlpO6yx6bta8HlbCUCY0hxD570KWg3s9ghqIlXJJVsVvh1S4ivXWj
49+3Zg3F4sjz5q+Sw1M1xp4FH0nS5Gm6lj1NjDQwrlPGpxKxHI9Wi86SQSPAqza4
/I5WR1Y8t++pinv8tuXWDBl1vQCb6wkGjwhSETEK/IA0pvrVzouR03PXYu1qZfKa
RCcoMZVLHSD9Ab6H1oA3GIaNxShHLWqGkDEHDFfV/dOtEBm/FOjGA5bfzIBvxGwX
I+wpoWnT7AW7nZQaJSBG9yPc9RLYIi0wrX+beq5wFo2uydslqViAfLCHQTNhKH1X
nrwh9e0t4JgqC2tV2qEUTAHVSJF6iAhmOtQ0idTIgOqX/id6g5S0kkX3Px4CyDJr
7fqPtGoguFQIHPE11QhryqVgDYTyOUS8hMUT8ZiD4qKv2WE/Mu+dkKUYx1fPXWBz
OXcUdO1EQftNCEN8JHSsC0Np7YIZFM7BaJ0Biqs45Edn/5NY/0BcMm2dbwA49VTx
JtpE1ion1cOY4knCLpCrJ30eKD+pPN+SrdertviSY2NGKeVG0qTpT7stPBTe9IqL
ntPx2cumZpRMe8tt0CaTcfL/qgeesrBFeist81L06KGe2UJRmhBiOOlUVxomr48K
94ZrzfbQ8OVtBMCYJxby7x5GYDFvCXbyQPKP73Tfn5HaJ+duv+9iHH5t5mbRv2lD
R4F8GfR3vD5BJz6vLiZuNbutjWLrJV3+qF6FgwXSBIx4a3xqjlZRtl883s1oK9Ii
xfukpnVGvYJKG0kLK3z5IV28O3fFq7Goyu3xb2MCJv9qD2sl0nhzTuBctVdy8elb
asOnT7w2lYHIOEzZg4M2LmU7aVzLhFTAJWKrB4BXQpb1uPYTY+CgXaf260bDR/b6
AB5tziZFkYJk85kIXOsf11AdORt3LREZjUv8cFvLRc7Rv4fpS67UCCF+/uIXt7YN
8rK8CRQZszAjmCHNjC/6iZC7lFI7aiQKH//JVHRb3xgDZYyG2XX6X0vu/vJ56kU2
rpqn+dA8iGNbN/+F2AA5a7NVjT08v31Yh96CELfzbes6DrczxK6+vWSQceaWerkL
cWtKW0rMyAm7m1WESIpPlDTetAOVSyKWjNHAn/e9xAVoxai3h0eoRminwzxZj8uO
IQl+xELmwU+LjO16rVzGqO8o2BAFuZbXQLvUK19n4b+kFdC0A7AOPUg9E8A69aTO
+BCHrH4bRoL+snF9JaWPxJEtXQ6d2FjZ+zvxeT3udw2m5Wvz1qUD2EMwzb0chKM+
6oGjYsw9Qwzsy9WCBqYG8kdfmY5iMo94eBSd86X7OYsuGWUOz8MI18/IXxSDarrr
Tlmfe6jJ5eMNlqZdVl/ZaL848iKUZMG4dfXDtQHvUv9MbyRlmorIAx1/Eu+qiYVI
t9gxx/yXXFBoSUskvT6gpYhdLWrl3UbmnGz3QCCzHmGyhTpjKXx9GbBtYrkk0A+p
QObq5hYBqxFVy8CkOB6I1f6cM7YmDb8EfhrV4LZCH5NLJOKnbl/bTja+RuArCkIV
Ks9kBu2B2CekQCVxRuS5Yz7nGOZlFlFiq4xOxxcVweSKhV2Xt5g/3uB8PRtrt/uS
LHFdeJM3lzliSQqm1EkO+gnFKUP89nOl4I59l8/w5z2+AAiB/bm7nc4Ecstf/W5i
KJWTHr0VjOgSga5azoOGC8YRBkBQJpA8eyXgSN7qHXrVKB2HL/Lz6W0yAcvcJI4P
LWC2gZrU28otNpiLmUtFnhUiEtuxq7PTlxUnp1fZ0113bYLzyIL1SLhedRIbpqOe
oRiKlLhBqrvSZJVHUZ980pjmCRETkCNv71d3ZOArMxa+3nNtAKewSyTNvZapxPcf
GE4VfptlcaWSoBI+AEI4CeriT3z4OLQOYiFbZ/MkUdPtsSIA+ip391Uum4GAosUf
KWWQJMFX6WO/GqiJxYjnQPD/PEWkA0Pc3rBTKiisaDwGR3KA2hXnzGhpfiC8E+pN
FyngWn9roB//VuxYIt1EkxGrcuLLDOXcNgTX5qWDfKeoT6OU/qzwWTNkIIc6c/CZ
FGW/WD8+FW+K4sk/Y8RUt12eVnPK47X/UZCFrg+HBGjbnHTSvqc0/q9nwv7D0AMU
2ItAZNXIuRQk0dZBpDGGJ5PPu8tzPAmJSRs+gDKlzL2bcVwX0kW6cZKKJE3A/j5p
wxOprYTZn+D+q57v7a+Dv+1MUiO8hAlNk8H94TkZu3dvhCS6wcNTUZ0B2XoVBka6
lTL0laG8wpBtfBcNRmq+9t9pQ8bvMcUsBvCYMSfdQCNbS1YcG2ib7tbpR9NtBqg5
lYj+LIW9dp/SIqNuLQbAu3NROW+ErQ4n11lb1wonXkr2XIv0wAqe8apPxLUzKfCY
LolcUAu9icVMUF1f7wBwWEuCXnT5yDI9C7qe1DcpA7DYUMlforAQWpzqN/4GbU+Y
7CC5D1Nad1iF0Sa3BJVpoXEDInb0zq5OvTPFutQvMObjhY5tFMXXoV28ChIyk0Z/
+tT+QwrzTlLarK677TqVr71cFVblfAd1RQE3Oc2fTAoZPB93QcYsIiW7z8HEl5wy
sEw8HsyAFfK7L7a69Lp+T199RdQvijEVKRMlwelxP+VJ+1JZP0cJh8Cc/yZXyphv
GYnhkF3TnF10dwBfWoGq3lG/cCKJFAum4wzna4uScENlwJPqiKoeRpfEk3wJ6m7P
bXWDAAaM2C/tKNied608pNH53j/S8GsBg1S/G1rqcJM0fRQoKd69ItueZ/ieUsuj
kdb7AUWpnXv/6g+XZqsnf7y1SOACqxUXBWvDFzWJtD7fA53zrjLzGUAq0fEFRmX+
uLbCzwlMKHbI04rvrftz0wMZh3FkFwKExCH/f/kICRsCN05FdIMoLf/1BWmZhOhT
B8fPbIr31z8m+YP9OYYVpuvTnF1PK/1k0L6r9uzc2U3UumcbRkxUcCC6V20/VjfB
87BcVHePgno67CUWCAP8Uq61N3UM2Orpq75HzpYyWom+VyA7OUziIHV8AzLe47KK
BHd1VQ87T49HPjYIqFYgrd5loDjFcxT6t7haf3kUXBIKOWKhzz9YKhsfcYTvhQSP
yvnQOdot9SOpmxeyQHkCoy89AESM4xwtvI8ja5MKcu6Ezki1uvhZqJqqPHUe6hZ1
mVz+ug4aXMDixsMko1gKAomZN+75bgxlCBlm9lZeoERuneOOXwfVX0lhJ2+h+6iz
od4q8e8f0DKJrmQXLRtoGHmESc0sHL6Pny6ChM9jquxLfPkcPIkDL3GLakTiipH9
lH0zDnfqqUzDwf4U7qKeq3oPicTrboCZCQ+HHaACYlLglAUGpfz2I21utVAMx+gL
NMrimpBMCxrL1NLxKtWbPZlTQ6oqK/N/qYlnknUM5g7YFxIk1jEiyMZlRnYN4gOV
A7CBsuBzFhU94qKBNiBRvKhzX7pFxfCk8pJ06KcDsmn0YwcShRAIXAAZ18JIshf3
BSVCY0RtQ7HbfBt4XR7uBwpTdADXjWcHIlkziBbRi9Bs3Bjf4u+3TgEOfCHMabQa
DceudkIE6bAzN5UTM8Zqm1ziQAxCFhvCsaXp3tFIjQpj5r78RgVkNm8BBB/7Y8jB
sZvbdocu25coWS9gByBFgaW+bsRS7TpB3Umzld6kZwosKTv+BqysJfyhkS16qbTi
Dyc5HFqcatQhHzNHO0mfyUfIYkhIxI5OdijxT4cglX0kKfEYigygveqkyDwpUhi7
5oNPZjAdocOIJ823Eem5sz71eRgjE6Xg58k87fTvOamCFVUvr8xFnW/brCQbMJU8
9c+71dYHawb+RhaFj9bXzGA1dihC2TncYQ2Fw/7Q9u2VQveIiD9GWegiPqJnnsLg
RNtlQdYqfICJ9ywNoWBIYTY1GFgyR+eT7ospZVGAAlzLJih24geOLzxpuHU6DOpK
GF1lJlxoPzjrmVdyfT9LtzVv4TgDP5yb1c7cTXVL5OND3LgUdNelo7R2D6lHHpMU
xvzJ9v7vmFCJQBGLLt+Vpq+C3yIeTFCRtCtKIo5NfCMbNhy/zjkCL1W/RfWwDKK6
N/7haLJqVsI8VG3h66WLqDaNFM+l0P2rOXeLpM9hBwMu4JFGhcsQHaoaAqRPULtk
I/sfH/uuPd+vXBwXCwtnC80kk5jKKsDsmv+x1oLKYEdK46onLtSUrdfwtEzIGcVQ
PgaN20lvAicUWa3Xljh424sNxEsEia7twjhsd3TRnLO6RcFz17kDK8BZDlVEQSfe
nXLRiwNSoGKD70NGzJK2YrvJFgwxunmTqWRkcj5svk9OwHz0vOCYKRWmcdPg3jcG
ZEJE+JL245QbxUn3V7FPEPCM8DatcYsKGo8EbS9zfe97wbS/d4QONwCROzEHNreK
WBInUPatePsGJowrX6W/wisYPV8ElemErzLmqfhxOBzwHhswCJiVJIMr4/UrLrIC
tZxS1RGfHTmg8aOtekkK01FnRHX5zFpNgqyrxw5Y7mrOv/YjXer072opz7wHMIu7
fy7JfT/yd1wQC52h0FwL3R9yyhaEau3k/7Rnw+tzBc4LEvLKvg6gTTswbxVuTkWI
KjzgHkLoMq484CULr49oBvzti9ckg0KyzwdZ0ZHIyGcvCCSxhHVowQtVtf5DdZmQ
5Eu3jFHKWjYr7W3NQQJX04Wf85PBPaj8+ex7jsPtWSJpBCidbH4vP8ud1hM2UTQs
VihJphFlOc5TOUP4Yx+z8rRcfXmFDN8xMMDKoIpz7ogZT9YysS5aFcfKTUMmAts/
30c7ia9pHWpAOAsfsji2XfDVLnH71Vlh6yi0xXMSyLHSKwsFyFo87IawqLJYQ/Z2
JNWNT9FIBGrteqyCU9vldv0XHVF5CG/fSH0Izhq/sMaF15p5yTnn423o7LzhHARy
uHEC0tw1+90XTPt6dtfkraQYP+tZkCiVRb1b1E0jijuRp6rpmSHTm6VEJ5Gt43lU
Zm3hkYZq1gnj8MNpnFbxu6FgNrH3yJKiSwmrQRrpRQx2tupCVnsOgY+OnyxgMZ3W
dBgVslvCoobq4p56+rgU/P+FqDCWW/HUOHNzvXg9QJjGLfTc9p0h1GFUls3vuqHa
PoOzmrvL2gJqw91HkKCp6k97IZBTbxoYtWlaVX3T7hVZPnYK5vKd3NUAUlwx6GoH
LYeTLCiCBzGy+F50cEWPQntYKJoSM+IFqDeRF2OE6YZKZLMbEptqOtJGcKx08sPe
zdMCdB6zp5WoSouVeO9DjquxyC4+7KdM8kMYNkI5LhvXhCwrmy+sH1WBG601YFSk
2jyP5x61STAgDLHMrniqiT/SOrRnGVOdkbnrGH2wNwLDC8oYt8dLWRTiWsTj9LmZ
L75KHoIY6xG2gKp5SbR0ZMElhsOcDftdVTwj6zdSB5A4vnlz3OxWpmqa/WQOtVL8
zDQ1Z7ELtsD1ZeY39B5kn/XS8vis7I4UgJocVz7Pfi4P5hO3thJ46YwV6vw9ZhxM
dzEArDa8/Xb0tT7XPCR3rZfX6RJWwjyqRQK3pda6Mkzf+FSuaN2Mp4krHlfYdYKm
g5Ywt4+4Vj/t4I+Q5vR3nahVirASlzEwmTUtctOILTnPQPJImCvnDQUfjM/a0Mbg
PuWjA2ehz3CvoYXF9Af49q54+piUOxZ8XdQCTIkkoCd9cJIb8M+IXHnsGVz5lwzk
mgbHLQnq4X3VDpUUoTc6A4tKocUcdZ6Bjvcg49wxp5UUAZ2ZHNYNtrZjs9IUYRAj
njEh9FEm6P3uj0As4Ov40UBK7GfC8/3XfHGkvohrmav8Z9r+3wrRu7hYxjgpYfVt
+kIXif2jMAzVc2gvnpr0iKkEy/vUP6lhYpsAd9cTlQqujDdtzm8ppq9A34CJ6Q0z
4G87NF9kVCezjByqc2N4IPSuYVnH3wYu/mpZtNi6pPNQxlnqaZeG0khRU5CbJsMB
4yYMGnbDv3g1mpvvrFsWmPEK3CI/o4/j4aviWdLXaLuIvAhIK5QrPnN3E7PlOCPI
3o/JQAVDL0SgwH1qq0f6d4g89d/r8gGcTiHUKMMtfxmcOlc8j0kVr7wM34rg22f4
NRKrvbbi8e/Y978hLANhyweJivxwdSUu0ywoVNTJc/2OA5T3FlVNGzc5DXVmWX9E
uFq1IBgjHg0J+UXBSsDbKx+A222sx2S5GHtkGLkFJ7LSgLEW+dnUNj5wud64eO4Z
5Z/QdQe8v6wEuFzmazA/NF76wE1A7RTGlhzVZitFnBukWaEJUNevpnrmIie+ESrq
YyesXFDNV7UmS3zrZFyPEojpIqj54v2lg/XmyXn58QcGGAYw/Iq0YYhkIcGkoJv5
x5dBRxB2c+LXRwKLNv+qxqBZaVAZPxbMJH4JF65/dU9QaKJ/kDBhXkE+7Fb8gdAy
RonZxcrdJ25RsCLfhxFb8UP6kbaTblvUO5bl4vWTyVZSgNkkDf86BUxJSa67nlEf
edgbElkuWaZq1AHkVFIVX8jBJ3oYHdnXZghsHi37YaQzij4fIHXyU40aIw2Ibxfa
zPKbmbxHR41TWH/e9OQDlRr4PlIC06yZd4X8uKJoS/+GIqatgBRKqwmUBSsR9A59
Xx5H4UzpGJBIlLvgQ9O8yrtFnQoy9OaIoVLMmc4V56ijGjs9jbtyRvZJK2yGzK8w
1Lt7yJKBRUzoq5Dl9BSQqsvymRtgi5KuoTaH2tA1JyUTRdjnXzZqq1Y9OPzXK3Ge
FRmCtVps3jO09IeN49r38GivzmmV2ep8HRGBbUD7jI7OBdR2GgQibqqzmMAeGqwL
5TP243gmjJ1T8a2jojxPwyGWTqrcrxLQvfVbVAsiUETmkf9dKEHPlN8cXmvCjBdB
q0oHvSjM7BBWBwNXjd7U95ZTyLZV8WLfbhXKP3WsjIOLEt2LlUG/QuZPszcwMd6Z
U36RJOnD4gokhkgcpBaMUZWJqkMTW5RF6AdtpVm+I3NwRD1SAugeDYxGISTI2fkh
mqupC98apXY6O1I7sMSvbqYTLEI8r1sc7NtWpd+F3NQ1Ww9SsnhdL4/GVL5r+GdI
S0p7dUlhLMJ/hcgI1L7KuJQiZlGecwJeqH6eFSsWPNmmV6XprKuYg50E+mwz5pv5
nEeNyVJFHbS/UoFRCctAgMk4L6EL6drnJ4c9T+yqjcr1L4QMImf4tlYyCP3+m5eh
1qp8D3LxsGC647MfRyI+rhkRJFJSSQWbp7jKShgYigNNE5Kf42i7VmtGziHlaqNh
+a356bazjd4kW2KmYApCNIZ2FIGIw2Q6QITlaDmaDRBaJkTXbU4b+DIEziOgLz55
sdLaGzCap8iO3jnwTZQkWLTzLzV+heTdgZikDRFW5eyvwNk8Sk9uNync8Voa5YLM
LYYx4wHH1pciKrC06PI4mc7g8900alpyZ21IOk0t3q3ooMHaUG/wBmlR6m052C5O
0iYBDboMzCzenuQTzIFlonXgKBZmQGWLesOED7DnzzRJc0y8etiMv3f4LcOWosR5
jwUJ6V0I1eaLIOmnXnDpd+ZE2lW3veRWUneGSYtwVCPIFVZG8PmAKhDuikUoyPon
/aKAucQCnTiwZUlhzxuq+UvR33UffyjwKSyUJaA50BrkBMI733gdvNE2qdgF+SYf
2SuIFdJp7em25seHSG9ZcjT6PuqBRorHJv3+9TZVnVLMPVNfbbbu6QawtX+pkZgo
YD7BTWzHNbcuYRKg0iDa2LM7pAKTLOM3N3RPb/EafsM79+2qFUZOJrrun4ktDsGh
HRka23uSFElkV5D2Wbip07kV5tgI32rV1oCg+1IQdkyCJO4Z/XSCIF9IwvGoBFnV
ydaMbVvSRrzqXl/Aborao/DsOJB7IU/P06P5IOlKTZ1FvMK4z1uNNLs9B/1ziLO9
80BsPFMfnxVVUgKZWLReM7e+kesX1r6JKhcWptLIgUbMAFpnka7iRsGi8hjy52WT
L3dgi7wojHmtesMt+oo4kb8CxOW89FqsoweMefgQsAfRj9uiTPlk8WLUNXQq/qtx
5e8+WYWuD4h/6QxJA/ueCeKeV4JKA79jadVznfpBG+AcSbhHbWOl6qY+Zz3pBtYX
QzqfoDJilwrxktPN5aJGfEefv1nr+4dGw0RhUiJAJisOrWM26Py5SDY3BJLhIs8w
VT0go2Cg17SawQgLOWN6sjQeHm2NJ+/kq89YPXnqC85YyCmJjwaLBr4bmnGEEDPW
PnRhlmGhoP36ektSOFT0yI3gk3+6DA6m5jwpdtKc4l9CUvgm7eRRpdV4fK75ebuQ
NzUoojARSnqJMdA1IGLrmquaZt7wQBHjw8RzYJEYoVD4FN6JyuFToVfvMu3o1on3
lgRy9zgufY2bfzDhjDPxaD+fytExvUYLuoEF/JUq0VBW6zLkB1PkQxeWM7eERjhB
j6t4YbTD8heXSfqGjk8SpAVEapZnUKzSG7yIQF7HyPVP7gwDYZzNdXOGu/MavCYn
yfD7pBzQvdHk+nPcB7iD1v7SEmF9qAu7R8XYiCg/ovtYgmu4RulvX1J1Lo6m9OpH
YKGWXDy+C96FM/kKEHd0tIE2aW4bduAqnm9FB+ruymfuj1+YXA3OrL1YcFYiZY55
dt8zzPvrWf4PyxorbYx9iPeTwFi9zrOS2FZQWbdCZti7OowM0EfkPLBQnjpUKtvk
WHXHDvn8wztlwE8j2hlmjZ0Z0Qb7MkgbmQyRWLuXO8S9N7MPftSVpHXuYCXwxL7b
WtDbWRMjLshzC1ArAP8/3SGTjmXYinH+AIL1z5H+zk6gR0cZwoh8dBmHq+AKBHh3
1KFdRUvPwBWpbfdHhMnNIaY6cFcx5gXSj3UnzPKmpLeKDieQ7+vHru9T21nrLPYA
PL+EqD1Qi7QZskeSiCdx91VxN04vjO0ydQNCSVxYF8XGUe70o2R2yGd0x6i7NUgG
h6dvhgjf5aXkO1Yx43LccIYdQXmrk1+to9DDbHwi6fK5lTzyUfA+c5Hk+hWVwZqF
2vYEu4aMjjqV1Z2PCFUcMfQmVdbNjRvkDUIJnp7WbIRUDcCV7ZUkku75DmisBBUQ
f0aLBJrICRMdfW0p2wxAe2qgXJHwqp/6Fz+qr/xHQ2lbgqfHy3BVLIIahWt6Qm2W
+0VHTueM3XRYamoULIiJQjRtSrgYA3MSW8NFucnGz7qaMX+dhPkON2cuYt8bbWaw
H+CiHggsDcFYOTe+6sPjUY6g0w+wlXN6ZQLymmCOTn2jtV1raM+fU1HVIjm312BE
8oUHILS/UxvvOLHxcfyfjZg+O/19vE1i06LPwxZSGCApaeksLq5oPoMinlOsoxaR
lz8qfsjwqXh2QMWvmPPQzruFI5BMF7us+gW5tpKMqVxxUNK8dVRQrAx4wPrJIe67
MbUScwquBLxNgGy5WS4JUoTZTLkN/Y5pVb79VromQ0sWCjSVGMXZtenItZVg5p2X
6ftkMVvF08Jj7JbeM4iZ8oxo0XqIi0ztbrrjfyFE41f8ZY1CDiVszyfNYuH23Sci
8SY8EBinZtGZYZTQDzntDNI58LCmSkf2DfSfXavoa3UE2rL2PVfjlq5V/fx9I1PN
9giFDFFoGTiD0r0F9WN18SVxWJHqKi9R22wvi8COiQCNl3y6Usbvv5Vgqc4+dPzQ
ZA8buN6aCOHrq/D6RSdhRPY1Zy+dQayCT2cLoUzANerUUCp5eX1P3L7bslG8vTbm
8ivEYxS3jMM9lNkMTgqeqA9e+6QyNJtVeePQMCWwcwq2fwV8m2xgu4DeAIgHKMvV
Uxhl6wFIlwkLSyVP5doN000Y81mlx4vJ2ImH2MDEQSKeUqqcUgjEojANfqibheW0
Ieua0C5ZicRlL7vHVHlXA/or4xr/T420tMrL+v683QT527F8cSG6A6ttnrfmNI7G
KdKAPyfAQ2PcCPolcW6/WhfMVPZOY902RbJJvfdy7JoTthKSrcC5QqV7TUB5Iz7q
4NlCl6CFhGTHUgV9TP7IGAmBQKUFLj/p04+yaj5ARi8ZDZrAmSc1vB/w/5XAlmPM
J2gautbQ5kpvBieoKcl9puGjJ9iGflpLl4iYJ24e/piMIAtcU72C6LdSfDLyagZz
ktekWlmdjmjao2IS1UnlDAtdKrJTgXFfRHMKC/wQoJh7k29ooyp2iG774Jf8sL+D
tzAzOcENORwQPgcrsBl6IWdemT+ovtIxJsnBhpxDZ7wfjTNTuo3dGGoGIeoxgpDS
/z3XqQFoI53EOhXr9gz6E+nHcQVL7nVXnVcMmt98VNXAHWep5hpTUouWVIUcckQ3
OR+bGp2m/MZ63DihgQQWxb9KVZ/J0Uvxj8HXmXDcL4OF7NSocfRocx61SGpAF/wV
oo4THakvANSPvTR9SpPDBbNZwCk2QbAcKVV/ETmjTG/6Tyb1pdt7hZFd8ZxuVR3x
5KprFh/tyXrC+/rH88jU6w9HjJaPEbrOs6L4awIaOqnl0SmT0kD8We0DXitNUJCl
UGyLgT9xQ+ptmX42qbWfyg7sE0rZX1U0NA/SfaP3slcI34csHriWXp/kpo/UvZBU
NajTtGPSwkjSfgJupweLJAfFKuCZbLzPedxcwYFhiQbvRdqn5Xqlg/xgXbGVysU1
t+2gNGF5qlelg9J/XXAb5e+wZ095oXNt/ilmuCuaAuCjiHVawRhjGemPU/2td+AM
hNAUk0fbm6lsbtRuqxvF5PgqA72MYUJ3yMd/OZVP8gTXDijpuKUbtgStuDNpbe/I
JSXCbRC2pfj3psbYBOjxiAofHZDvNTICCmeeUsaGygT0M5xnm+LSBT+ZjKev4Szl
Ud8kY7EyS3qZTPhfWVDUpc+tEMZyKEJGVOTjzuIGWi2NTsyur+qaI9dU9/H968lK
h7rtZbRgp/qgUoj5zGv8SkgVqa0zPcjHr0YsUy/ryjpnrkJScR5UxT2FDVU5jW4Z
ugazjkZRtFZEPD7yuG7cumLGudYa0/4V3p1YAbuc+/JqsymixQUgwAqSxdTFHc4/
I8fa+/ie7zC3hPN7R8NhcrIppK7olFCwYJQlcmVaHRYfoTbJaQvQVyGyAKpJVqHP
F/r4C3sIABBExXGusFpid/0tOuW/9wvZduQqhz9EHf/O9oKHtPbQ4m27Do725f5i
FXNLEMvjHljqVWu1exQQAptN5EtW9gvUwYZ5pZrTORuYke3VknVHTutbRGXoldKL
HRTdSpVyrJx+Sc4WmSjtaRApSh9iai3D/Jg6SU/tJeLOe86zpsTCdtGwSmefpKgM
HfAExZfE/8DP622b7ezQgJyhp6eJtWH9Ctaqik2FFdGltrfPgggDHTB8+yX6SPni
MJHJkdSvE2L/SJsnXW9UdgGp/8bI5IBbys3f3qzhCZ27hmWXGXWSHDypfI2wvSKg
sBvmSSMnapM9DR0FWjGV/Clanrd+wjI/T5vIJy47LzJO+NEgr0IH+9FhEo7w5IwR
rVltOimr6PTsj8hJC1Fofsnp4WWTFu7zGz5kl2Th8tHS3mqAzFN8hIQkkZoqy3+6
xFbgDvRwmKRb5fFj+0J7mKNIGit3U3eQQplzgcFeB0tYtdfrfGYOH8YZZOJc9UqG
S7HpW65AZylYlpPgpou176A/4LwDYyEgrakpuQJo9OuM3V7EuUq0uFo2kQQbuY6n
o00bqoOuDed9Gr/K2OKvxcqbQ54N7SOnJ9iQND870+TLDnGsJd+DbEY7qbZRM5Rl
8RZyLJZqW5UhNQweTndnB0DOXNj4X+VdCTqcaVcf5x3E+h77GdIXmqlrQD81AXNG
HA7PQ9M7gGwLAhKH+sX1SK6MaO7z6FqS/I3Xx35VT3bfJE9rckQZAT3NtfEO4mNJ
0nnb7wnXi/thyu9URz0PttWN/iaqxKsrezV8MwkEd3SPOC+L4HSwv87HBI9+GUoN
l5ekd/RwpQgYl4Vpj9znDcOye4V3QoKyG8IiYLPHwTwsGSbzkk2MQGrhExtuurSc
Bqt9pNVQP0WyVtI4Q1YzQiJN99fWD0b8aPPdcHUFgmMDCB6CmmmXt5FFI4KnVQI6
bekfw0wVq2torpKkGNPwZk8xNaHPmAc7YJtVcvFG2pasJGEnxKu0ck4zIoBROjdI
IxbywV/opjaqYmWn6a5Wv4pvTjkQILTAnncVMOPzwOrASQZ3y5voTKb3HklVAA3e
zUgC2RR5qNfzRBUYMi3K0IG7OU0fnT3yYLrVQ8z7cvLIXLyWk93ewXkpGUkynwE1
Y8VcJ1HCIGJTowuTxbZbDDLSwVv67U0/j+mFLrhLj7C/mKUX/LMHZz857caCeqLM
jr4Vd+X4b28qw8XbsgjvHpXnCeU9jksYH+CZJMHvvbwBpAzgVbZamcvwuuGxbDW4
PvaXNBC1jnrfCkHsBlYSWjIcnV62wdqxDyOKm2aeFWXH+lTsDl9zZAh8C1c2/fvG
+oPuEDu/cSh+Y/HiCpL3Pw45twI7sOhz5Y8psD2Dqxga9wnJCUXkn7ztZYMBjKU4
G1juJmhJa0NFGtYn79UX5pT+Ta+8Wh39aveUNPY7ceA/j8f9kvKe7DkIwekizdDb
g9eD0trgscDiTezn/V9TbCS5wq7Vqc9SjYitKjarHw9aeO+cmK1In7zRu0gX7l0S
XYOYhDOQS5J1Mp/cxK0CZBbhvPFrCxlf6ZOyH91EyMPEfO3NiBc0PYgO18m0YAk9
YdSUc3ZeH5U4L6Jn/2mabcRG1etweVxmM0PIFMXdDc9ZpVatUX9bniaw8/qBTki1
gHVVa3YZ/vmiwJKQ3vSK8/gwHFcJxDQNu28Fgp4redWFi6pQzPXRCbSn0FKBCXWe
J08HfGekUjPfCa+wJucdq2+XOFWZuAjLjPyeRo2+7RES8viJotvdtI3mH+gaAx5H
7ia1Gr98/OrfgDNeoRhM9BS81BcLnZDVrPGyU6xazJzPa4hnQKywMTent/EK7/Kv
C+VlEBXx59if68ewHz2L6UM3QJylMcbBuPJNpfveVCKaYIgqBNYfDqKenJmMTF5e
97jv9nzJQAdni16PZ1oa3xNHRFa+wzn9ierKM9iAvH6BEl4kSD3heNqPickxKJni
vam0LejTNojoeHNqClxfAmmiYfH4eCWKN7/70z8YdkMzzGYYvyJNupIiEB4dGt9v
vcR3RWRyvVBgC8X6ubjyci8Sapo+chW6EeQ/rV23T2L/vilkNk9Ob0udqtymfHQr
yctqXcEaysV4qfzCM7B3ohiWMU9mmAPm/7gwdfRcwQ7tqR/+HggUjMmJ0d+GLgYE
LpW4SNhj8mAuOz5yA+A8Fre0GDuuwObc7rsolbWu/WCuKP8eqZHo+LPGR7lQ1foI
XY/enV92NA5mWfOZFFXhH1NABIgvAEqEKaQ2S916TtbQX46HZaB1iGuU7nl3AWkA
qTD+bm0MkG/r7++monTfCJDzw0kPGdNANFliEDLeGIVRwl2pwkhromHO9l4rBXjU
o5rPTHRb2oos7N4AnerNFAMFZK9QLOx5ljlkQqHTUKUhVeE9gXfPhFyRahLBVpRP
14VWVbR4RvFy7Pi4oZS/ehFBBAjmIy4Frfhy8I0NBQjN5MTpEX4giSAlE5fgsE+k
BOgeJhv8wbil7NlMLkHfyguba9BufXmNry9cOa7hRLjFz48qf3g+B1saZIBo3x1/
satLCDk2LYAjU+KwnVuIu1SrzZnsBzb2UAVGkbVJnmGh76IC2ReYcIE+8ckVnIKK
KS3TlNGprNnc36MqPFv2vEPhPWxz7rmq/6rKrrF6N0A8O+ScRRPqYsXuoi1v1Jb6
7k6GKiCgweYNGzkMK9ZoAmXcj7tNxeTGcz9B9kF+u5Yq8JjDKPILQ/jsSVaBa1VH
qVInzlgbPX+3fq8bVrE7/goEIPFuJmn+bJiNDKVddBG11bDSemhIm10F2ee/vWXu
wc9rvuNLCm4lLTMUQK/mCHN69r8tRGuJ4plzhOrCW8m4jwhUhD0pKMeA5kqCNsyl
qFyqqWkTjimb9kc2qLk5IgYhEDZWBktMhSWp/UD9ClcNg8khYEQkYZm+n3hI8AXs
Il7Ek6TImkGskoUNIaI5vA7ysBrVCZrwlVQ/RkvFu0alcyspjhaQPnEhb2D74r3x
iomHmO97bhSAmRzQ2sLZ9nq1158p3+4LyaxWAbN2i1IEbc+Ni5hzuS/1T2HOgm7Z
QSTUDPikxVAGTISQtPGcNjZRs4l19NdO/jngr8vasQ138rQfFfGZqMQbDpPjkmKT
vvv8Fg1vGPXfRM5ALpxf0d5br/McVWltHeJ4n+N4mSKWD3kJX/0PLOmHVac6zpsc
3dyNAma8Gy3RuefMoTNu3FpGbmhmjXYKBG1SCl2d94AUmvqgMNdXJg6dBwxZNp+u
wraVRkkzhIZKftD4eotG4GW60lIoQT72O3B9CpjryxfyQAbVRL8VA5aHjQ1An+mX
8U9GQDBevRNcSszUPPeD++U4te1Aza9xgtM50CYCk147a6klrZGEq5ei2yILjT39
8wxd6CX8nwkpjiKurg8ceIkbb4j27TyqpH2WSu2C3opVuLDWP5uoVSe9Of3E4ycI
oJpYxKalLc4Q2eQ3SULECXXw2o7dnEo3XZ+zCnl40mPVB/KXOzIb3MVZ4MU/1WMF
pnkc0xgu0HV8U6spoTyi6quNP68oKnmBgUgiNYWWxIBdgJ9pVfYeQXuy+jm6e0YP
5y+Iy+m9ttcynzaWmLKCWjEOrFCqz1uG5DljwRfQ5EmDxbW/ejoiYW04kI2lnVj1
pGt19Vi7IyCCM2E6KBmAX/HNJnUIUESi1Xe5KasLFqhxnWKCqYRYPnqtc9i6nCih
aaj/pvJ3w2yiB6LL9eutwnYuxQvRxMOODYAPRflHmRYVNbzK13A+CWmlYPcuViRZ
BmDddhaBu2wJVGH9JvpLyVSEDVIdmNblrjqxir2miF8jl8YxUJcQbV61VPiQmG3U
v0tyo5wrcJQYEb1S1MoI+BTxHQk6FS1eEyKpmxWEyv7T3U0xeJvV1mcuukrR0aJy
IQ2PT88pEU0IDgKeu83rKjK1OvaxSAzP8eawC9mPVN2yQPlbK1vTWHMQySuaHDRo
UjjazQAPGhfKt3LE1PVAssYDvF8zENV/Zt6lkNtm4yjvyrtt5uyytvF8styi5zeB
NoCLNlDeGXnZDQm9zkjET9PF8mj/jjeyn4CklL9XjG1pu8MyODu7Om3nRegE++wX
IM6IPNxlfk+rVflOtCD9FlK0/VNSJ1eZCmHUHxrtWhUmFyjGP0lRuUzg2CDkgU0b
bI45WvTxVclXGR2xkZ0y13YKAlqF3dRSUy/MH1dVsPinbCK8VAAPbleyTe/OVnLz
oQwB/04RoM7WfFS8XFyIp5ixeLKhYeKn/Q9KCZhmHBJMv7jL008UBssoHGKu1soc
w6AZI/e++oSCevl1IKvH8sEPWvPH9tUZEIUqXeOTMOCNfdNOTW3KGugI9/jrZSCL
z+sqwekGtq5QBFvP6S2+UdvOYXXVnp6cT4SHX4VnyEC5gcYqnagvW4otGNxg8wcd
C4qXKj16iT2cXo5gP3R211VZJQBDFMPVK0gQcZmNXH2Co5AxdOEH1Lc+D2SL+eNJ
ht9fP7aFhZItiugPwFy87vDRXmL4Cbs1zUrbyhKhl8smymj7gV+sfq4XyB/t8Dm9
pUxIQlgHXiAoFewTOedd8EB1tZcpDRnkpEokKp/M2M20HEeUibqNIoE0GhXguGTk
bWR7VuPDM7MKWiZAcCu+gKRFkv8pW0h7eij0Fpxp6gQOiOAe8OqFEjlDbIw5ljAJ
SAFcX2UXnYid6txWIEumcxtg90gJOf4YuWePB7eddShZ02XNNHFtQ4x+sYWo9T3f
NLpIzB5oEDn4K3Zfwm5Nu00jF01E7BVOgcfVDZ4TqW+d/kXb1IlvSEXq5GUh+WVW
GVYLWGLgNWg04SYjtUDPkOOTUo3UqgfW7mkUPLO0ZuwWJPnmqOknvAz7ITArE2vJ
m6eLzWLpHXwLjVUHNprQSVNEETRh1bk/ujpBt9FziNSBhGldNMUlfv0XcmevhPNJ
0bC88mNQn04NL7+cHGztRGgAOQ3fe2MWdVS5RSF8PqzHHdsY4oGjAsie2ySfSvZ4
ySh8gOQCmBVvDWyFa2Z2aCmIS//83ql2wJZEEbLn7sRLh0rjTZ8OJzXaKV/oKKyu
fFwS1/47j+uTIR6VJ6CyyoTwpLgeyLjruZ6KbRDB16jMT1UjSbZ+/D0FWMYHW6gA
aWzMmx1cj97fudinnGw7TnC5us57gkEb9h95AaPUrPRIPwq0Wn91JrA6bCcbKVuu
GCE4J3gExjSsqRSJ+xx4mxtpvu3ecFNtHFaTNzODyUa111jK5ktG5naZ/EjYoYPc
bfd04iOfafPUVUqyUWTD2ZgzLwoMOXZigfsOyuwD+i1sSJKGXuj1N0+2/4T5QENY
CpxG4un+aw6NwnYCzO83Gp06pHhQ1jgK/oqD/QvBNBvo7MWl6Dxfz3xs/zebnX/u
VJG2BMuGWhZWqKsJZksaFsL+H3Ngec3FpA96rH9FYJvFaHGNnTnpWK96X0/eCQmk
W73aAUE5lo/SUXE+Ez4hy9FWWK4fyVNDYs+eDEJIMCw1fluZ5OJoEQl46gIAkIsM
KG1Qplb5GOKpX7ANbAhlsiZ9WTNT6KEjnzjyzv2qKrTn1Zbf4opv8Kpj+PLQHDnw
/K3qOelXXN4WfOwMnTpKZKKZCsLuBTL3BgHM5+rbNLt/NELq8tZSz/ZgNm4ZE3RO
gcCpaTKwoqOV/XzuKYtcKof6px5fZTJLstBGFOIZ858npz+9kWrVyVA9QNsOBEsp
r8UK5jFhFqeXXuWkuu2ento2xWzvF9rh+35RgfSRxDdnsBomQsTd0oqX7spbmXsg
bvtUt3iOOdtbVy4bhjdpOluahJZfrHHqZi+It2qFbqQ+u/Z1hydCrMLoKBlbR1w2
kr99PfNPa4CRep7SDD808n9gfwJNekfAn0eBEKot1j9lNHX8wwOGsag7+h6WgZvi
J0N6yUEcfubFgK47zIyUlzz6/SnkmwnvzUiZEsftvpDrnJYeK4K2Fzkv84/9L0f6
XtYwv+wxCV9IXCPAKsgBpARVaw/CgzMD/s0/6cbFjRfSEf9xWeHTfLIsNLONI9ey
qvQNbGNqqHQrOhNPbNZUvgJTC4D7OGixvCLeioG/91Er7H1CuEzesKKn0sKTnnXW
Oqjd5svXWdf43itFOjB24uepWuXNlpl1eAvKSdtDELr3oD1rLhrHelYnPUrzlhSd
UQATVbkKAB4PoeHVhaB1ar0AZAMZTJ8p10Ex4p3XHhcfkBRoBCHtNzbV7FrRyL9y
q3xNqtmwyauoFyzWd9sbY8pzHguiG1zgDahlXvuT+xlBB5BCeUUe5O6NGDUIYgWZ
VbNX9KPJLIAt/M1/hfZQc8FRAV/5X06xHNxfVW6PbUU25HokVSAoyNN7v3TRtYFI
qVNg2V8gZn7rp1cb8ZSnjTd4Xd6ibxJp5VjN86BWCSdyeRuXYE6A5cGH8In8Pwlo
jzPrN5NdDOcV1Lk7TS7xwcruAJdvBXLKoQo4wV7kSdzjsQ8Rw4D75jz13yKE+FdS
fD7iVIRk6w/8qa9/Xo+1sw+g3bLkipLWTmt6rVExb77lB12pNXQ5UifMmteN4aeT
3GiaMmKE0FPJbVAdFVIAblac+eyHzF6CUpfBQl+Xc1vAK5CmnM73oipEQ+7/AJJi
uEhxT7e59iKvZfx22BDbVbbKpLCPwjBAApyvS0Cj1/ig/bZiLvEvYTWrLBOIZ22t
M3j+h88CBdnqfQtAvpJBfTxKEcC47gVfq+UPmetT8f6nESTe788cJkjC2fm+nnc9
qGXY4ILHCBRhTQBd2bnuTDETg68N0OrW5qaMhQeLbowYypNNKcySrPUWVBtS/crF
ZQ83F2SpnvbYyphMausnC3FvnS+dNBuphHK6N+DxKzcZXEMSqWYeCTpddTJuvd0u
ay7TVxzBuMzLzc14YJdVmvQnhBDOqENmFvLiP22FupRftejoPEt0XVfUwLYogMqN
VrEPUoDvHVXf1ynuWcI/jgi0rx/q0LYtOwV8bvxOKypsXOXpFT7TeMnhCVkuIoGE
61ZM2Sxtc2K/oSMr4xdM6ZC7EXAP+9/2NW2I5MvRt4Ajd6Gdmf6AZJTkENg8rWL4
mm5gtPJ1TFYvzi3ndO9ar5xO0qS7PxN3rGFGlI5ZxAE2zqGdVfWAFO88CTSH6y4e
6vLUFAK5iyiM2hxKB91rKoPi+q9PWMnXROYUar5tigGxADV2EwO/lU9O7+6oSvXu
EkJ5Fh3Vph9dGMka2DWZW+UUdFHN8DRpdC+YuNuWVT43VbzpGqrjm/k8dMr/GXRg
b9H1fSy0hOyh8zJyEDT8Ota6CSiRhSaqnCNzWm2PBAbExCrhxWPwxc+p9PwuwfP7
U0NYVm6CGv3yiiXY2o8Z3Cy/s6PNF6DUDVQBSs+nT6LYFi0RTo4UTKepYBGcg0Jm
cjPyPWFbRDQOvzV/PJZzgTCWMJWy21/XDPOmGnoQL4peHQyl/vs+4mYSUdGA7vo9
8MGU4NFUQTphE4Z4VpubZMDTc3Xqd0T/7m7DbA6n2ACDst6B9dm9bC5SE9bCwy3U
qaMz5Mfgny9mZthZ2ughCWGIZhhyGTySxnoyEIWVrefrciVYO9ZMX8eZpRC+uAqv
cePFhL8CbFgrgjqslcqzpLYPFUnJSHALlenmEGN0qCPLk4yOJr5B2MeDYcgwpNdf
gMfY+Nsj2HT7xDyZ+QZ3lLsQENg3/DZGqtzEsYm7ILWZB5tqCSeUqknACVPToguz
83/4p8EkBCfjNSyIjSDMtiTQTLPr6L/82ulzZ9seeTj77oFUVl165OqOusVbyiaP
8OFn075JvJN81UMWZO2hCWVjIdvlFBpNhn+d08Y6xGgfHU8995XQTdP7uqbVyEzL
CGYT71ZQJQpyHXEB9Ykxbg9mmxOKw8jVa2Evq4y0AEGRWb7El23/8SGo3iBfYGx/
FC61Hf9XEgoYWMTZp6p5tYg8l5wuqaUtXIjluWc9DIXvPZnx6Me+aXKjmPF7lecV
Y3fMhXm2qHYCUgAdqoE0TulPN5m3nhoMYmcZsWFqPEjVMYPmTxp4jtC/jIzRynNb
zokW/oVPmjKUyQYykxgNWCRylfM0LdT8mUwkVjLMBVQGVBAkLHIi3fcgwo8x0c3d
1gWhkjuvXOLv8NH9S7Mzl3tBNdPlT7DGoAaGB8oiaZ0TNlE1nO5qs3tITXA7j0+a
yDpu8OCxIOs6EjFTTOqG93wll/L8JDowpMNciOentmeMq/S8X5T9goAZejobmLTb
R/E9CE4ZFkniIXfYPAbY1hYJtrzeG/CONd4lB0Nebomj4q1oPLY2YJIUs+5rkJzQ
KbrJZIL3gUoL82oaB1D2/nWj0D9PnZF2gLTdRkD1rB8kJJGuivheBo9Qcd8JOllb
5MJ6lB8dkFUBKYaLZOCq3wl3Z4cuaMm0vgwRfvQC8DrmkvOHYx3rHuFn3dPximD1
lGa9piNoh2GyEXzwOJpAT0eX7iKmRWiaZOk8Dcx3se22getn5JUMd8P2n4tulBeS
XeuifA9vm/ef5H03zGF9BZHtsgCwr4Res42FzPZf2WC3x9j67eTWOYEp9zh6Rt9Y
ZcdKeIlTfmfJo4o+uxXJAlhN5/D0eYzjv0YeF3GpMQS+wHK21Vpk3M/ivfGXP46J
zdx4DSi3UWLfAIc6n4SEYR3wrSNGVQks+HrNH4pYE2KrU9r8Yrud3mS9JqF16qH+
QnXLaOBEfC/pAiXve7O8lqV1i38/TaMFGxslbFQ11LnnHE3e5nXDyOqxo++dZd42
+g9SWVncueWb+3k7r7WnMX2whE+BL7RkxVZh5FeTOr+LGzB6vSxxlcY+Djjf0WJB
Lz0hj94A3faC7A803x3t5FGNyJQAapSCTzSAG6EnxAhsNwgIvmEmlElLtewWfoAa
hU3ZiCsihXcDSOUkWCgL4lQ3wz22d5ec66gmfBv79ZD1oqQQ9CaELdaVS8rlmac6
c++ly0av8rym1XQvdSrU/xF4S31D9t6yJMXzuv54AfmEBk3C+SnG0cGq5SqKObUc
Q19cccr83XdIbwz8DuHxRv/2iKN/9rFURYYbSjpB6VPHqKrIv5/D6Gi+WsKoLOv7
/L8bjDQLziDyDHF9bOfwk8P8mjuZLuBuctLn0rYP0d4zZcm5Ufr7EcdDV0ZYcivD
CIzn047pKZ1CifJ4j+W04LnumHjI0nJRUztF9rMCXHQMbVt9k5b2mWvvo37gw5WV
5/aDBPfdWw5A3RQOBz+qJQ7I5gHIvON/y6+41n2VCYbtmyWSCPks3w0jYmYscpr3
GkkR0Pevo7DsBLWqKzm36xBsbvFv71lax4BCiQ1vcunF2MJz/XPuoKReDgdAejH6
0Wp7JdyEARrL4gehjEZfb0iwP6ijbRZnQhrKk7IbyEmacvPGitu2kuH1k+/HRD3i
Z4bFwc379Ud6fRv/9mjx+9xOjQCW5oDsiCL2H9tnP9N00GtCb76GtBMII5cfQ7rA
9ktegWZPXMixhKcj79kaMWUIctcl+3YeL7k1nR3xKBh9hQVLU3WDx3wJp6h7EI1r
sFeXcOlB+2fEqrB2WAKPNbLtWwJkZyVm3okvRL4j5BPN9NQDozH3rvV7Cn8ZIQRd
pgeQXBxnJocFO64wEDfeX0f9AO4ro1uAx4sSvCAHOncgrwGOxnDW3tmj7ylvQAUd
Ua46TEuo36f08Fh4nJjNMjqa2+PLICsaUDc2+bBIJH4rrT5Axz7I7hntltkcFC1c
muvZBp/kxnnb63OSs2m48RgX2c9+oeIsKesg2nqHUkZhB5744YmRkj+OT9o1Qn+z
8CasYEv55fgT7Pl3+jaHy6bcy4yBltVmc7LSXQm6naaslUv8U34tr5dxqYOpz9lS
NqTNUtBLut1NOD6Y5YODO3fxNVGLoYQXWy2zV5ldr0cIb60tTq6Z8LXX9PSGXOs1
BCc9DmfrA3LNRB/Pw5Qg9nKv1N3fE0EUqO0F0NuUlFanuFs/GDQSfGQtbCW1utIH
voKRbgZP1btlbx0hVF1euqu97Wqzjzhci3sC2dY5qcWvqsWqxf5ZrgtWyosHPCBM
eSIoTywH5qwHfec7h4n0JcqwNajqlLOGo8WSsLBgXdEW91QrCYK2CiDlE6PHdK2m
laXqRfWWoRXoxRu6W9EpAZlX6Kfeoai8bqK1PTwM/gewTvr8gnkrs1V5+S1Xu63G
+J6+ZhhNq6BeACmXBsKtyAIEr5M4N4yJk/OZPkzP9coGJjeN9kYYvlMBhayy6OWA
JPs7Ttm5fgiex/jxJ+8n09AWM7sWV9aM5wfMNS81deDpxw+9airTPpBaUyKiqrom
jxtRvrTKwUT4maqjZZLAsCM/0zH7rwDXXhy/saW4jXefhE0ht49p5rL2WY+pxje0
UN6N1KWOVNAbbxvXfzWd7Imz60xhxeuPlWqqjs3asP3XPuujOzL0d3Ey/UwzLi3w
S1gCQMo7zJAYDe2uzG1h+xwwBh+e1kyrbqj/QAf3Ixfc70zc1ENC8uq7bqhv+Abl
ufFME8ZrWW6PsHedlKjZIPK1hoS67NPDL9prOhw3IV3J0yUruqCEUf7EdbxFCb6N
5r0gTq61+yK+Koi6YT5L+lipgoIdFOVALGpa2y+wJ0LIUp2H755K/O1ir4bH9hpN
YkstL+VS64MXpklu4yUYveq/LlS88wYCn9TMjJx4aUk3wnDAv1NMYZdefKi/Mk0O
+a0MvrywR6aVDQfBbEt+FGbaa/gOxIhE1ojO/SCX5U6Op8kCDTTGGZc/w/OAtzi9
Qj2GiBzC9X2MSpzuj9u/ONxE2l7st18yhPJ4vR7H8zcJkYru+2VbiL6ckdxDUvQO
TJbvMHa+/VYjSsDft95TKFYSpwNI9KJwune4fTP3xTVxHLRu3ZQN00TmdtvgtPcI
NYNsRLPxH7Q1PPgC8I0rP2hJqISpMR0L8c8T8RsCJi3YeBrQ/P5VUxRKtdBpr36g
rJLbCN7gJiedB7trdK0GkjIAO6UF4yOkAO7YjkNkQQ2MvCNADRrlG2oQBLlExgQl
IISimsDkfevWdHHzWiX3v692LmgBDwdj4MNWVo/hS6f7ZqXsgtwCmP3K02V2X+Tk
rkMkQVvwOUP8qLjwekuWKdo34t2uR7sLLWcVXaZjNTMcR4+uLJ8z1GNJv0YieJtB
IF04bjo9v7YfPhcCH6ef3E6gUOT/OBpi/Sh/xWfiPLa6T++Epon4zDl6GDHLA2Cq
V8nKpdsOYMIrbPtxHZfZuiV5uEP3DTwRHuYexTIXdhRCirMrYCA0poW5/yfE3tdM
qKwE1b+/FFUdL3J83lpBhWhrG1PKGXUYSq+DVgIodLiB8pH6luzPIRMvshk+teAz
8/Q/TgsXUCUaJpu106SZCFYuLHVU4vmdqprmXzQB2qOagen3tnhW1g6GyhdbOY/d
dZ8B0x2ZAKyWb8HJGAFkiEwxcOJpdIW1pFjr0A8T6QIC5xQYIK2bNXyH8ahCXv2d
AxoOvW/DhJrfimNVFncOCvQ7TIYTkLJV4bo/7+kjhkzbxFlinlDbQ49DZkKd4aVA
1JFsyuFAzUbotSjlCFGXnEndiyTumslyxtOSqESBsGOIncPiZ7mlGyYSvsps4pP3
bfQmwY8ra+CjCn/3gkdquUZcvIvfntnKd4juStiywKvZcUIjfJvKzeqM5iZf1GNo
5YzZygcjKtb3TfjY+IBWTxxyV5bCIJ3qOi0sz04kmVR8ttfcf58RBeHc8G0qgsh3
vlddpXYTJFVt1W8tKbfdwgKBYiuakbyTFCfak+eBPFIKEPM5HvjWBxFEPu7ZoFFr
wLr7ekXEoi9CMCegQzox0+ASOu7+DbXFrKXGIJs6mTnGR9Y7Eg1Kh+G+5mEm3x8r
5983rfu/1/cl3LrDhaIjNs3S0uTvgXJugxm6LkER5UZwTr8V43QdO18P+XRQus/H
zR+91vM/t9J6JKCgQPry43lUQjGStOrzdJ7CdMJcTE+eLuexEf+j+fp1/iMLW5c5
5aQfv2CBjYCvUfVNWHtSFLIsnum7sdwDejlLvgxpajVP3tQPPL3s4S7SLEDACi8n
XquQyzNSUGuxZTK9XKgvKbnamGKFUTvjkP4MvXjTze07BWnvdqucOstNVcGrTSq+
BsDtG0DLj0LU7PF0c28U3TgBHWdwxab5Kls9NlOWvjwzlK0hF5Z8BSBf5B7YLRjL
VzoNqAtzSF9qXbanalF3Dgl4BFkNpgtCbrk6tgyxlaHBwC6iNh4EP86QFN3J1WjL
Q28oR0L56tP/EDxyDKJcQf9iLVeHKBJqQlLNNbmL/mRyeOVvC44imu9e0Bne4f38
y+Jd6i9lwp1V1hdYvreKswpDIlpk/Nzlnz7Y6uicOSdTkqf5SxIpUA/pEN0qGqGT
dXJo9mJGe3f/Tybvnaa9wvm1ckBxoymj2KvorwSFJA94SkLLykxFTORADGKxs146
m3CLbqeBb1Tj/egCjDcCqrAdyN2sQ7ACp4QsMhjrzlVVEsbUmR0B2dx2tnj5iFg6
AzIElCODSa3WBrsVo2wcsmQ8oHtZUQHgNof/8k3ONwkwMachRKfSWaDo7+KIjOYO
+Thx5Zp2havzzBhIK2reXrfEAvdPOiVsKD2QiEP0BcAYDn8ZB9dJN1xlcT9rZAzs
Ly33opSbx93Hiz4Ueobb1QwShpGigldG8owtdrBgfCzQjNDhVLqmobpYJ2HsIbig
QNbiHAJjS91ppQviw2hEBW3wIZileHa0dj627sOQZYODf8Fqo0HfvL6xfB7URzb9
pKaK/MwgU59wM4W+BxAobSasRWh0vyC3cVmw2BOKRjXV5rL2pfPaguGH+XyQCPAf
rYw8D6Lynl0sck/MmZm37dK1BaqVvJbUfH7/2CHlIN8063vPf1vWXvELvw8uwtJb
uTLJ8xj/hJW80bWxhMZJGfHC1oNfR8vm8eC9D+XyINxw/XfUcFFpTk29b6jMF73T
1TjVwSzAMydqS1LIIHNuLL6p+XWhuuoa2huc+xkEFIbBn4btU3YbXAswc6subKKs
n80qTT3NgQw/7Vav9L48CKOhNdYuvK+TYYbXNUgCM1bCe9GhJUAsHhZDfh+wWeCd
qcQQ34yQuQ0eQWrQHA9jVT0ZYEJLUif8lvi2/8aNWzBYeCsMuIDIBebtNmnlPjks
7SefrN4SMwp5TdBGBH4Xpcgo8heRuYaW/oVg4u45DoUJLkxE0fjVplsNlD1pDzuD
lspdnK3/WVgVtFnCrRcIyrYv6EXACACI8SxGaUTNXDWDtlbLAXqvptcP4AUwlF5g
/TwWqY3IzOlF/toGLX7kIgyDtM02mPJAOVck9zvnFwOCub+1hcvNZjql7zYqq6Rw
QIylEYG/YLGCAvZbxScQpA24cwWGu5HT9to7+T51ENYYaN4B6AjGBQrYih2JbBbK
qvAbZ4TC6hIY7Hm3d3GSuhERdjkW3i8QMQhx62yG09LQDnPWhkz2kRmt3oVBcp/R
O/XW/6dr86G2fTNqbjk0khxCkJzJirmnru/8aZrPgEepkR+XkrJOeiO4Gz0hDDIm
xvHZKpXG8dtGOD2GLwbotzOObo1mSCXQrRGJ6n2jmI4P4c8eNSaH+phDkwI/y684
RObaz8tgcNB7t2854nQR5z4GDlsKna2a7IqAlJ7sqWGap7HidGzfXPxkPCW9xbAj
rgm7N4S84VgJU5BO4/XTZKB9nnAoejwuAqcuqrFzEPSleErFEZ/m7YNw8VaS6vLW
c9vGfX7uO4z9evMYEyV4Y1vvg6g/bWZmbVJWjp2A2WA6tpegtyXOfsp3WzX/+m7T
+5c29CehYlKZnM4Art6t/7DQf+eGziYB76JVfErNTLq+qoJpto8ruTPs+ZfJM2iB
hiNWlXfTzpjDinJBJiSL4603OjWjZiiP/IklyHRmybcUzjLo6Yxvb/RXsr0fII3j
taQuspozlWWyZr4eOGVSQMAPxp6aHRLIErDt4nub1w91kdjulyiITqWPoVjlb5RF
7oZE6gTOyn4tnV5mviSlu1dDEUC2oQ8TLHF5P5zJrvyvjrpr8H+S8eWiYoD0jaes
AFDFBiIxrU0TlLws2H1kZ0PZ+ZlDy3lJDSk5q8n6t28bE3pIGtzAUMZRf8rxVgvb
DhCsaIOCv3cJ5tCQx/awFcZTHekYQ7pL8ptyVDRDPto24lZnIm2aPiytB2tjIVT/
h5dL8Pl1LfbphLVdMoDhCUIP0dHeZG6nUYVTbZuVRcwg5BGSdXgNObWz1SVzQXWh
l12EWg5SolPotqYhJVYZ7zyBoWxxLFGhXXv13i2cbw5Sa9N03BGWua7PVDLtmi3T
9eTmYR5JLRwsscbWkCBGDJAD0sinBEGGV/HSWFjI3ZuTtU7IQiaep32toOafjO+M
DYdT3WiB4VlO4RePwgG9URFMoX+gpVk967ja0NWnb1Y/T7u7CTUSqne1Oa0V3Rq8
5HpuK+OhsErTY17ucuJAc7i4ER7qWat197s2/dlCZzilNI/hdWRh82AQASZaLzkR
MiRm1fDkndYjNsuknB8EIj79FUOD/Lz3tfZD4Tq45SpS8ybZmkT/5Gd1/ukDg5U1
z0Bv5xyGrMJnTy6Cnu6pLOiGJ/3VVVTQfT+4PpVFbbcYPkXLuk3GCUOmyOZqdPof
QfQ/RFz96cUt1/7GyDIxKFNdK1naX5F0tHnBWGyQ88si59a0HFExewNY2MldFr5m
QVycCX5GnFsXY3KiboUvPHxQ1zZ7C/XRHluYRJoPKIlB3l26g648R6BO+RjPCxHz
2aCfL1/8emt6mVFnJpmUGKg7e/Wn+Y1z2hsRZOrfzEI39fpC7PnoJNV4xtT0WClP
9uNrJLNV6hCu68a9dPrONnEWbFF8w3tgnHDCkb4y5PsgoLl8u2No5cHObY1elbB9
GT0DeXHIRq7qmF97Wz7SJV76p9y55oU8SG5qJeYxqhQOpV6R6dvFkKDrjnnFarB5
eZDfHmnrLZs7vJMEx/iwylXxunshe7Sh15FnIPeyLW3m6063GXWu+w7VXJr4kWv/
bdVOKAEoe1x6F2OIsdAWg+JVaBc0lTxKeqnVGjUU3wNuctARp+wi7WJsr8CSqu24
jn4LM702zU4rRCCwxs6CSTLvceUKMMKC4XtFpN+kQQBVJ4TL3+lD8NYqMKAEk9WR
flsuz7OnI6zqS9d69Mvudz583RagZcFTra1D4Efw6CnlYGRDhsQAqXhm+OGZaEtV
I2vzGzL+byzwt0GxP/i1+Gtun8A+iqG6WlTDIk7AKCUj8oGOQap1xNd5KxJ17S7z
Q31Wys5DW+cl9mXuLLdM4nNpcT4H2lwf5S1m2rv8NFJTFm3lLCMrtAqStYc3UFTG
uyLL0AG4A0eq/fupmwWIbtzss+hZiAWs6h+tQlwSObNHnysSGr2tV9fyZuoRnhSd
MQ2wMZQqv7iC43bNSRcg7HzR6LLJiQUwyx/6YeBMZvnYOJ/Cdvxf+XIN2KF3iG1P
Uvbl3RUVh8OjCb+c/xW22UYgwo4Gf060x35ytsbgBUqe2T9H+j1NXEyf6CNvOY7D
9JAWYP3wkQQ79mkTrbvSNvYQCqmXQfSC1iufEzTNf95Hbd5N79+D01AuGJQg365r
nFOmNBCn2R8QcNmI7cz34NAMsQAG3EuVbCIBCESfvF0lBc9TRdRhCqD2eN8osNJJ
QzISxe8w+E64xLnQA0Q+cSNmnnpBD/w2Z0cMVWYNwQ5+ZPmh7iDSpzDi7WCneiO1
m8e2eQvDp3CZnW9QZCenWUVSz1T3+5zZ3PpBd1mMR3cO5uAWAhQAtk3POqh1YK1K
2+rWNskSvux1WdSBAt6l869rlngnOUgxHWmOS5mGVG+rrtZvC8CEujN44BaU+lDG
/zPGsO3fm1dGWCOwo4A563d6vxGFBQ4ScnM5g/7NQ4K19FlbMA2H2XOId3Ry1phS
9XsjGH8tiBo5sYGINWy/fQvlhtU1kcJr3rFx9mjnNrjzp0xlNMXfVl519IjRS8i6
mHBMUYohqdPEKM9w3fzUO9FmaZxMf4+BBYI3vOk/35RsTYxJmNgfwQL5/hnusNDn
MWlt1W4S+ysvAesfeCtAw199JrZB4mO9sMAamsH9Xf5PZQks7gfR/Q5q8xdDfY9e
DnhMrs52KVrdRnV/nGIbryrp7odLD57yUGgei9omR2DgzJO+9oHsPfSBpFYy6/Mh
yN9yBkjgqgzZJ1UtkOGTlO8AlT3sTJEyMNZNyZCK2WF4EyYlu9t7mvwEdjJ52VDU
sfUJ6NpM0PpUsHixet115Fu8JGKnKQyFQcalPp1bIuJr+e2J89X8cRSlMX3ro7Rl
KODKs3tVNbqZGLeeearc7fMPsCtynK8lpcv+8IbarNNID0m62i8ElXRGT4L+xx6r
TrNwe49nKBpRWKxWP7AO39mkwkeUU/nVavcGChv3YvN3OdRZC21we6QbSKIgrCLy
xR6AxlF4Gv+7V1wHY4DHrOlCw2Y+CAHJpOJLg+Mkn8USvPkYbRkFnAZjzNnqyQn8
hCk0CRcJy8yaYBohnndlcPlSe9ih29i7FEFpTxW4unbSRRY3yxf7FleVKANMa1qg
4T2PyIT/ksDLrXYn/qAILW4Rjoz7jdEIaPE6igcsDQ3o3TlQRQSOriMVlDnZPrRR
ByB0WdTaoCK9nbcallwpivV7AdEyVKbVvtMueurLnqGDg4zqQhn69t98KA5I4PJy
l4Wwv3K4PjElKset4AEYC8I7+BriBIlgRayybdCPTQTE5sAiSNWUd3A1oI7xKg33
9ygI3GsGA7UafaPi55tKGTq7BSmwUARwPfNu5gEppAd5wNCvYN4498hVf1WW9Xus
OVO81Tg8V+Y4PxSjSY/ef5yzqVW2gaOcTRSOmqb40oNBScRheR6q/1tMEyMhlSDN
rWvoASDMU8kXp/6DCXoysR30+kpmjaT/5tZ5JjDMbt/RiYeN+3gt6lSEKUgCWEdh
fVmwv80hjELulICAy+Aybe3aARo6ySH3CB/pHJ6bqsvYclb42VvWwWtPQ0GPsDAv
bQ05jch6cIa6PIxBuPrylHE52ZcDWJ7wLez1s9U+PtzOYLjzK1Zc9hC1Risn5K+J
G8S4d8kZqR/py7CDZ8BX/RUuHKkP0sb7m3YUJYLlLh2oYkMdzqGVZ1HAl9+ATeV1
EdkjTV3YihvCK5RpL5Ws0WqFBN1vJBhxrmdWwHC6TYOKrZXXKLN2wQ7j9ZUJclxb
iwndR/+VTPKxxG0XY2qKKyqPFtLs32ahmI/Df6wJ0L7x1FIe2jTFuTGM5uPVDduY
69w7v4x/yeTnA42sdVpnhqn30zZH00WLfi3TIQYRvB/pYS53WXbt+eTeF5+eXpr3
EiCioS1UD7X1tC+dh7EDaMUr/FY7FH64PXceBhcGXaFlE2Zkow5YbFyYyXNsgHQe
HiiLCgMbP4tQz2QKV2jyi+zQbO/bZqkLsUHMrUg1vuA/D5+z1IN4MADUcx7sATW1
MFPi2Vvt8H07nORTP7iTdjT6rmdH9oDnJi9JYNC0Ck3TaqX9Ov87AUVp/GkfgAkC
kqdS+oYka1ITk6sD4juR8LYu7DPyeeje63TpoK1Vzm9IefnEoouqskKDnLGrKm88
HIGYnYpkRkjoCiUvZiPKzI+rrxRAQnLHOtwuym/sX84vPU+mYf0Jq+c/ScNGppTq
N6Phym5/OcfVlPkk4zpUU20lxP6h/avchxBFSQoHlA4XcyDlf/Q6iqLa4ed3yxOB
Fnoi4I1JuZiAAmMG1wwKLh1XeM4H77q2Y9dxM9F+RdMK4hyqOIW9TBTZFlOMSLk9
Bf/+WM5DInwrdANYvW4RGFjmR2BvIcqLhWL3ImRLP0MNG8dzlpavSl6QZBEsQm86
i/0Cr1LDgoY5drW5X1vX5ZDHvnxsQfhablr9fLHxcZTkb5NNJUJJgBtbNSQmfDZg
GtL8juqfICRTm3+Fuvcd8HCbdWpD2gpiHMhDOWP2GpudpjMP94rwmr8WcDSZ7SzH
9Z/HCY4+im4bZulDRYxDdU5BhYG6bUlEbIY2Iz7ihgmVmHWghXxNbK/Ah6q4hpij
0vBXjnWu+XdrvsITsyTefSTWnIgdveniYo2XIEdm08gVdVP74ePXNkcCCZb9cJQb
/oWuTFOVRXZaqbCvf3BDKnqJkO9qUG9b4tdsf0u/o1qscTMeZV8fro4XyJ6DvuGj
2GtQLTeVSgz/o7UHBb3+b9aTtmXomN9oALcMzigq28I785qWRK5SUHm+D2CxtgAl
/NlXGakjezBlouYGlSqdXQkNfBFwNCzk+ksgnHq25on5++bgF5qosgkFY/KoLc7h
1LTVMaJgGMn0ufa91busGfR/88aspJdR4mS4c6kiQBqzhsHwDiBzWrS3a48MNdr9
E9NTCvMNCNI30gVt82kMXXuvPLWWbu5wp8+cBHA0tmS1aGg92lxg/7SbLV72aBAS
mBCU98GS4t1MRi7WTiem0CeibDBMkynvcz/vKG3MH0w5LyukeQuVkteWz4XdQbf7
Hc+pbk4R1FAbvVZBdg+8+sR/lEP10hCKaYnxcyjgDzCNlTOqpMYRH+CBSS/mChLv
JYDfi27XWhQBdmmMVtcX0vIJdwDu72iFoeQEWfFAZ2QdIbyFqe7I2K8pEO3BHf8W
bGDzs+4TWuU7jzUolcWeoOydpKzCvr4LGas8LqgE5IwvsKx/9vrLfBX2KylpZtxv
qPtkqUfel5yWh4jy18KJ/nbE4ZvzDu9ifI6jEutNtbFNLzI2IAlArNnK/b57grVI
TToZcHo07xZuR7FTTN5Maw==
`pragma protect end_protected
