// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:37:06 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
aFuDekOdfK+DUXA7BlgZo2JOTviADEmSAx0clF4l9OT37LfANWlLEZs85E+/Tq6Q
Eg/NDkTYPI9zQBaJTZhwuZ43F0RnP6VQGVKZNGxk3wEMPi+bUxgLaYY11xbozz6E
DtbYOpaxH29SjOUazcAexSKqsulA5DJ6VXI4PpURldw=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 9824)
mhHZmdyXSgdGKjNjgJagbxXSM06JTNpaXe7CpPPSnRrMfRJObPeKnIvlV/9D73/x
uL5LBNR14NP8YW12XTuMehGsHe6YRkWk7v9Sr52hnQP/perx0hlOJKmtAnLErjJV
1kSMJC1IC/fQ7hmk3MZqHoSyRklMT9fRsZjoojL45Al4+nleft7jVSFfec+SynNu
libN5Ph0P8IIrNIxvfNj/nDZyb6q1+Fv7qqQ/boV9QPYfccjc5I6FWHVf/hf2m3p
T9CPg1BOACQYA6QgxvhzYUrpRGx00Hg0/M2aT9nCLPbcyPrdZGfGLS/XRquruw+W
/SMXShuXwQvBdPZiMeRNtZ0MX+LHjlq7kjD8/CVmHP0A30O0Zxr2BKq4nElwlguN
hLF6KvkVxlbZdMw0yhbguSZKkBYkF+Yu5WCirewhkssqY/VzlpWopeGBiyhUIO3P
wIolMvijmsVhGK5Zm8s5hjWfbTtfB76lFGnKC7lJqVx74QfyGlHtk6RJmBQA/Uzh
h4kz0gkux2kUTKo8xir0HOjS4JvYMLFwrrism/GST/lhAVuNAdRopHgYtnBMEJ2b
lZ6Mp7OMPhBh3mu0k1FmDx438HBpeUaYCOqnFnP3mkANMATDmYUtcF8FUCUHKD4p
+w19uoGGee1wIgVnbnLqvIltPZNeEMGo0pXNMys19bUtqAd7wFxd4+/47bo68GIO
dHBheGMf0Icb9FQ3VBOhYq7f6K8Vky+Rwya5E29Qaiyqgl0h9LbkJ1LQeUOJ/alX
TA6UggXTbmo9PDRWJPuXL7mFKbu0erM8GWXiASBVzDN753tIG6eD2+SOxs92L8RT
zt2m+1xxO0YaZIUqXUh8koYLr37u+/A61jP5sKmOHBHkHdyjS10fhsBDHOn5PFyR
1TuitxkeN2dWL6fAjVbC/V6llD6R+mhvuOtrde9ctCb7EFxovWYueeC6tFxV2TjJ
QsL3ADwfmswedHZFzixduYxHnMcadW9O9ute4QUV8mjaagPjKk2kMBMCTEThBLwA
1+5u5ER2GcX5nagcXTrItc6fwrlPoUxWavKVvOhMXCutmfPy3VUj1sAUrdtFp3Kz
7I8ISEgB8CtBvnHnbvXqmX5I5xS1IyEjr2jbC8meliT6KjCajRD+loK3Esdgxdjn
HK5m6jc/H+DDAOPq23QrjqNYf0hR7284Y5eUJNaliXNg+IO1sVzi9egEUTXVr7pt
5VZte8CbwZEjGzuOPHH7z/fS+/+e/FOI5K/CY/txu5JGpB/KaSa5h3p00kJJiP7j
NMrVCmIae1pnveM9AmJZ1HzAZc2K4/+woq/zaRgDqSAKj7HC+nMe8ahumSBBDhOa
/6mQSwqyQqaUNz0rtNyv2xkeaIJTljWbwbusf4Wt6J2KmYnp4wTgX251e+2GhfkB
I1vUM35Au33LDkGja6WURyoCbP1SUASPmN4a4ZZEMMqO/NJFMJLhHZw1CyvYCWWP
Mjmkm/JzjX4g4w5TmOfiJsKAdjsYFSPecmj7F47NJOAigP5pRJN5xlgr93KdDtXI
Rl8+6lzNePBGNeiA/wJgo2FQLdwMB3gS3CxEdJN7nuVnWmCJAM8UlYqJyFWh5QMD
zPJnN7j1VBiyIKesy7MiCsiHO1+4euUGGwE+pgpJKO9xDu0Ky6xVg3ioyVmdDPMa
yvNqDMK2hS3U4NNdLmeS7fBaxLUcZGMMDbCn4Pwfsex3lCelwunYGQ8Xr0i4uVtY
x6kAF6eCO95Cn+c2eS8Dtt2Y9723tpiNnzEO9VUlI5DWMRoBJbgBhbCAnfS7En+1
cmphoVVh0g4kRoenYC5js58I8yMBWMbclS3ZZOyIK2mqGKWtT5mBpp8RJIPv4Zcq
5Nkvtn2GoNiVTlMd9bbvVc3MBmwTwxpCgzVaKZanaly2+wuVyNvqiCg8l8pCcgTz
tISDfbsErgUBc+MOwi1PpCPMVvTY85JguUK1LdaYZKrw69pJCT44ZRiQ12QVQLZb
jCnZFINPi5qvm2fcWUpNO2bb7a24xBFXURZBVwJznrHEyTMWSnPLexX8clmXQ0Yp
bKKDUmI/N7TTQ83JRII+Et9KyIHNXKY8vgJrPja7HIIdtJVOm4hHFqlGed8E721K
bYheWNLA7npjYnQg+JPy4eoNYISugxfLAd5fQXbpHopnzm9dydDT7zBqibSLOzp2
NGzvgbgy8X/HgZ9rnn3myiwxMrDn1Rs9pXk0T6rrM5cA3BTYSTfQo34N5c6K4v7X
tpNwITfoMfBhRNuIQ+QPEQTdPwKIbogsoditqQYjfpflpJJXfS7ybpzGfkAY8H9a
yUFqoOe4GDEWIroWAVtaZfbRpnFnXjgGmHT6dAQEa1g0Y3+loCj0dcmS3FtCOYWl
5sQF8YX4VcNYM4eiD3Mk2So7G30K1V0t5O+poib3LVBIomeR+ZOgyNEXGVxlKK6O
ydh04u7LT4MxRLqq96YcTYe0dXCLVwFGSJmNpPxaf8z5XvalQF/79im0M+VxrrpC
UsqYQ4vrLtQBYiAof66my7b/NPR3EZFwNBjJqleJr8xd7b77hmsZbqZcOUJtn4G0
2Z3C8g6dBi4T9Vgic8ewaPCKrfefJcaD6iHcYyr/mdPkF0hPWsIh319ZEdEQzRK/
b480HMlYBzbtCnloFBoD6tZHzC0+1JgZ42fny4yFQ7HwDuDWEABJPzkCK3NbjVJC
6oqncnlfD1Dkz6kDjuKSv7yo2p59jK5DjdTCIAZM8Ce9/OxqjELjYKVe1cXD8MoI
WwMKSpX/OMjYMX1OYaIFCv8oy8G72brln1p+Y2hNc3E8LUu3ISqJaJd0ZDc+djW5
cu5iu/6qCryJBqEkfl3yQQkjhXhV1DMx3VMS9l3G31w7JHiS46br2nE2l2PUzYuo
NIn2hBwOn0CzWfueDO1EwrMu9COc6Oe8snM6SE0jA/bs9b7oX1BAf3hr2NspRbKV
QZO5RBCNgLq+49ybLoDTtPuE9TV1UzjjxE7ZzolAV/DYlqN6n3+IQjxMBASd3UjF
mU170PSt13xXgjLNT50FpNdWbQa/EOHhvjRb0OtnkYwte6cQdyF6svS2K26XVCnB
7sS0pqJ/LB4hpxXYK8APPcW+hhip+MJbWLyxujKBEoLBgHqjZIsEssGzpu2LISNn
Xj9irjulA9zqrU3NIymppSVi7e+iVpPxx9yLzx3pFH3p5F1v1Md8ICPr8jQK1AEB
nDlLlVALXEXneW1P7sMzUfO/NZ1oCTmEHyc1oIL49PL1NziXmmbvbnSzAEvJaV85
L4E/g9DGuJslxMY9vSZZfjJlLwAR+BXla3z8FOeB4qi6qOgRyiqjaerfC4yhy6vx
ydeJmnALAJS/05k+/hmqbUfkPq3cmpVM4N9a7qM27xP9rpl9XnNFXNAWWDVar2yv
Vj5K3xKhLDkPjz2CzvOZLCJTcoUR2ERtElJqCDN/gV95k5Tm97dcLVlYnOXKHsE1
hvDuC+3pC6rX+VigwGcw7iM0/vKyxSZDQ2gJYuUDt3oyMnUodzyIDqCF/DBVcSn8
yXFL+k3bzsUMhiP8L3l1GB7Iuth3ErgYOgCBb4MYtcq5UiEBGMEvf7291AjA+of1
3i1JOx5wz+pnYKNNoqfupapHKShf/Uf5fCWEaRZ/Mu38hhIt2M5FXYcwms+na+7x
hfYfm8q5Y9pnebshoQxZOxFRBuL8hUNQY2LIhDOEMrBNIxCnRTMbvWto2sziUOJF
BZfu3W+vWVsqIkDGiZMmAZ/ieHyOp2BMOv3twqFKaUO//yahxZbISoZhrg1Vvmaq
1hLOFOLGNVMt84nX8wh18uvyqArLAEMpKwK4vc6AG82Ym4MRt2htCQ81umxKDrKe
kfJaJ2/Sjpy/nVcp7trECaQxk0KBO+3pm7uBR64sT3wXaQihEVo5TMqHC4strt9Q
THyLRuiZKtolexfV3Ga/hd6xDStzzfWnpnaXEFFxGj2g6ofLh3af6GO6EPZoXgJO
0xbuVESKutH5e6bkt1MnsgKoHCqZ4TfDbLyuYjFfkB1faRMABuLkWislYI1R0Osi
PXIzwfvSlzq8V4c5umr1eQE2UIdX/PvjvMV2VNwOZEjWK/IAbfulMZWugcNGNVV7
yyCIS071Dt3vB30zsUy9instwQVEslRoat9rdgatZMBI09RqO25zVodxc4ReUVIy
wi4AbXSRDsYlRpoq4kv6mTWy/A/OR66H80uI0rNIwWlEvDdGStGTSGhFrQTK4ej6
GwIctZZoiH4iZ5qVE18rA9ov3Wr0B8SUNwGWJT+RenBQjAVeuIP1AMQScNn83x1U
1Vl8W7p+TU1rVAe8ym0nguDbaf4LJL+Dj6On3GvfvzxsQjGyRaJtXHxhXdSq6vIk
M0doqZ+leVyLrUdx9T3FkzKnJlcvg0MX9wHYREIL09zerzSH/5WrMDubJ2Ih6vVj
7VSyYdt4XmLhdsMO3xIZv6yucqMf3kCCfsRyqwvaB4quUIcywc6BQnVpyZ19BTTX
PgyDmp8Hk2mlKQ8EakbkN0iOOX0SOyeYSdDiTjJkEqfjHj4nrzHmXJh8IO2rIKB4
hVc6U5N+BY/MLBrp1pQs5XEe9gvJLpuWWQBUbqrOBg9LLrd1L04SpX8z/9DZHgfk
3bpitvKFqxjinNl21ioD28H+9IVOByJDXC3u/gl/8uOlpk1TfX3yvbUW6umbACT/
A2LYfO8+wNhlgcxKomvG2/1U/vkA32JHgGgQV2K8ZyAZ9oYUSITWHlYVzKsdfEbx
miM8mUVXmXv0/kpEQ1hvYIvoznr1nu7s55WhWFg3iUvKTXxMwTw2is3VZHEJCDmh
52AAAV9jXaLFG4/Z/c1LCWL+S425WFjpMIevrYPc6Hg9vmGoPRmBvwvXeviRu8js
twL5La1HaC5jp5S9cuStmtx196rlfIxYBaHsnaj9RMW2MZjT7syrDE04lBpULbYh
V4mPIU89Ipc+orWNTanAaA0qM5rB6fLdhtp180zzx2o2wHu/s+LYATJcZcYY/vFI
48A3Oa5Kc1UTJbUbLf/haALaQiN1AqtyMUK0lnKPAFYS6RNdk8TxnG/zPCEXcUMX
TBsWxUFAMW5o2yMO5bv7CCKHArz1zeP3rvbIew879qg17PeBOCdsu4LBPkg1j2Oz
TB3ScGUOQVLvO3aJmeY6ltHwnuWECBGaT67AcpbxDAFcVWO682vnFAr33Zn8Ng7o
dAtpal75xrlbAv6K/AiZO1e9ZL90ZzVSx2XQQ003SOBmLPMeo0oqb1DTZHrlVZ4U
HOYxqHuIf/DKwmQvczVnnk/js1V3yjtnmdcgRAj11pKIhqaAq6EHV/eem058Rzt6
aTHqUytI38J7v2lOo1gGth1Jvd7eYsfczV1FZEv1Z3YMwdwkj0ap92IDy1ipRGlL
R/1PGRkW3f+i/a3gmS9lCxrqkSEBvQOCG8TuanJkC9lEUc4WUV5mJFD5m9t4UqTX
2m1uZHg0ud/Ycjw5/4akjDJW4RNmOG1EIMnA3r2YAHZOZmFh/h+4zGuFDxL/lPd1
XQ6jvhUZcHfdO768NQI4+3rzPj++S7pxBKLi/vWdQ3mSD/v7Pw9QVtg5t0MsuJXV
B7kNAZv8ZM60OCJy2kuUr3k7nJPL/bwxcLlH6/2VidrdN9pwDV5GIRs67k8N6QAJ
puaeI8hkB0FGsvDQKJlPE4Rx9C+SziwT4vpGynt2aSw60Zs4+gStCj90Cr1m3LhG
yhREiXDuX72l02GolBNgzlJv0KUkMmP3f/LiFbZEOSC4FEaMIg+y6JgQmdVqT7NL
ThqEOp15XjjOsYl4/NBVWJiX15yz6ZZ8c28MoJm+NJ9PkLR4txcF8nsoSeigKRLL
aZMwRL7OrGjupihgTG/JFMt3scK/Lhfpl015feHefkJeid5I8KPgWZuBOvK2kH6I
wMfkavCqLV/NtDq0Goqc33eBCJHIkcHIsvqycXeDZvhddMjSNa5PE4W0nc8qvudv
71dU18ygVQ0UJouaXCooPqOU7scppf4nkue+1ySpXsTjFMICJs+xjEFORJpEQb66
vsmFve9a3aA/ZKi2yRgJOzj+eAsE+7mdhYF9ngQfQUYxt6VDEHcfz3b7RqGABQxS
2gKLE6j22NUTZ1Z7cG2Ulib8Aog/azOwsQ0S4Gi97AKhb4keqHt98HHyewrXbPSJ
EtnUOYC1Kl8A/oB1hSF/7h2w5okuaAGY6j2I+RwMaihI6M8QwR+nfHrcfFxhe0yD
tMSo2V9aB2XIRVvJVRp5I+H4hBH5YOntZNHedo5BqBqqrPrZdPqRVA9tvUUXdHcH
4l9FM1/kAeReDa23oAvVtMQEEg8igXLCGNqh89l2Vr544mhKyZLQIXvZHqL7vT4y
BUOP65gbW7xJbNXNB4Vts7+ozwvR4v+5O7Bvq31/iC8/d7oFJVR1RptCXhX47KOG
rs5ur2TrX9DviRqLgVgkuIsTXwVgiQKIPGxdq2GjCu+vwdZVGr3CVKkBoqZYEFIv
qj/91kID45KG4B8ZAgwkYEGRxwsM8w76Ci4AjaABBZxkFeqsXb8diygDFJ+5juCR
YkSGwLe1cHpL85iEvBSOEX408ZL3/r5ZJ9DR6276u+1wLLIr0HAxvq3N6nBmMYZU
YY4oOdumP3ZhgTxDfImZ+VfR/AskYyMIxxk+z5G42RF1W9P//PMfUBfRE0nKq5J0
JP2ipPJFyHct1RsC0vthDSO6SYxhJ/D8IoO8YsaJH9AZsh/eIu2wCkcJ+AvCkdjs
sg3h1IbKwxPIA9tY3UIjFkRNvguH5oJUisYTUJNKmHmhhKVS6Xyic3Nw49dt5y4b
N3+e4XT6i7iup5AE3tDyBUlDXtX+7CibKDoFKRnlFqYUIu+TYUqj2bFFuznS2Fbp
Lk+FE7Ct7vjz96Z4rxLMq5EIoW/rRwnLWv3B0kIZNqDE0i4xsj/KP5YBtOAcN/Ts
/rhwiY+30dg8ejE5N0EgMQAk0KbfXqRSpek6x1TTDo2nrAJVriKARXvk2lwYGnAZ
OCX1jHxWGj5Sjk9PUISeJ/mrYuJAyeJTkY3XSsjwRspFF0VlhycHcTkzx1i1Tpaa
Z2Qe/VMYnJUxZaxSN3fK9/a1/lFZBpqomZum4lPgrC83UmgkdMoNtF4zQ5F8xUJA
JzEsoDkcapz6vh2tkZnLWQ+tftfkLY1XgYui12THZyu3QMqos9ULVvWZIhjs+r3B
Hmw2p0Xk4WeBfpUWDVzGyYPWGNTBqouRy+5bYDvD+tGcGyiQ36/+OX5iQatyp1Tc
6Mg/kIh5N3cxs4PS4bAvGP3ReZev4NFpXsbgMfNFypNB5CfYYfw1TgYCm9agh3ql
mLMgp3P29/48px4S/mFAWVb41E4xhzHPdxu915YKKmSNzTUTFipPAfApO856UxQ7
R8ZLwL1IGUfJqVh/Ga97yhMzQnOp6pO/hDb2GgpbElHDAc/1QGzztBX51Uhdx9BB
c8Ybp6/CaEuVe3iM3f022URuhICfDP7O96je0V5WKJUZuF2LFXbBET2CvTXeoCoR
M7OdoAb9+eI3+1eCd46ZMyOkJ30/P7lECDflo8O5JRvFMENpD+BUiV3Fsc0kAqNb
M/K1XbNyPI5fSJseS0F7qhhi6C3Doi3fiulYWrH9RkYjXSw3W7/ZfTtG19JTCQs4
rkzLy7V23QhLYTK+W5gw/aRaSmByHqs9k1IJlzWF7s7QbRkA4yLQ0FWqZYk1kkgC
3RPHYRUe3u5FWmZvoAgb1Rqo/4rgUWrgcqizvcmREe872jR48hLmcrMArCn0vCYU
pouXPlfEc38PMD7lBzUgG7KSuZ1+oFdXz3fdv4X+OKdjusFhNZCYRpZua6oYI01b
1Y+z9ZCRFCUYQQelKHt7pSKcErz2I+TNKHF6HtVY3j/k08eRPp9rJkhtxAfw8eji
x8Hz1k7O7DZ65wInOBC+wcmWhR6JDyau6ptdaen0X+iNcFv7EpJOfii4FmLrfpcP
Su7ZWSgzOWMk+Xg/eQIYvEN25s/kSCkDYP9QbVxDfmSvfx6x2it3eNehJa0+lAqk
Ft+JjlIyLz2l+StkmrXeU7aKVdYq3eWTuZ1SLabgP3GD4Kn7FUpLfYpo2td0SbnY
gwi7d24ioJNquy3pTOT0YPd888oaC2EmZ1VBL9r5mTRhtMd4GBQcPCf0GRILzY8P
vaIFhSKeaFtt7yYwVVgbJaDC1CIVDULdjKLaGPbxiI4FVGiXEulgKpkU+6zWGBbu
ZA0Sr2F6sf8SKUJYW4oKPowahuLW223nwn7UrKF4DLcplhptRZ6b2bgeym/PGcUP
AB3Ey0hiVJ2Uv2n77BtCDRy5tz+FR1EFjNP09r9qR06ax0w6vF2+rtQ6tku06sX3
InhVx2jW6sn2vi5AL3XLwPLwlSw+GgPSOTQczP0aCCVBg8QacMSGlnKYHnwu+SG5
zgB4hjoTPBsZRS7etvzIRCiBJ1Q/HdY4d3kcQEWctns3Gxknls7Oln7c/7VUcTjT
w47RNZEdIxmMga7+ynq5zzPOYR2gOwXiFgE7pfNJIVROVSdGpQnVo4ANkh9U701E
p0Hdpo98Ws9zTwJYxBjLPZnsLOY1tSf7l8gCAAN3m6EQvq6bXMcDQ/XOdocVjuTQ
SX8lM1jis8Jb9aqRGGSVBRt1K/WpOpRbCeDeZIryZWPEnNdmlAZsSl1UWrxCNhkm
tyPE6tPFG36O2mkRIMrUvhZk1GYW28LGXhMjZfE2e7lAhXPFeHfmR+7nAsb/cTh9
D87F2qpQnBgJfN+nQKRTn9ukUILCQwN5jxEKAQa8cvpXGd7uMKvigl2wg/Z8KDkD
zToBEmuJq8tLaYsxdOGYYOd+s4LxjO8Jm2oV24wcf+jnXuB3RZfDbFzgPwwCyNou
c0fxv9XeMC4P+D9EVv7nBC5UYYwFReKmE9BNp7vE6bRRybrfHk6Y+Q9b2ujUSY1X
h21nslEKJe5/XaF8xSv94EBFXkfWXNr33ecyi/4vFJyEJxnaUM7gQiOcL6R9rP91
M9pMyEcGGFNgpF4XDuc0Luq7C2ZrYFdixowJosis3RaN5cLjwM70ntpsDEEl2shr
mL7kxBPksfIyynyM9+diEKpNuYl+YILQ7w3oCMzlFBQzK4DlBduQLwMYaSzWrVP4
Vg81i77SxgKg6c9EycBSseq/ah1kudptCkpE1UiizRpFP/E4kqbcMkN62993md34
EuVkHMYQUsWsBkaARbIdG4Hn6KgK+01r2Avy1RtaKQDLVFl790WArGGO3t5bTKbL
wqle8Mv+dH2u/WLHUnH9RqXq4++2zHqvmFKQ14nOxDKf7+seZ58AK0PXGs1HXRF8
Bk1X/pTe3FiQHDEYb0RKwQBwxtezM55PSZ0WOTQf/lhqOUrE1x2QVYKnLpEt5ryd
XYXfE0HLnHX0KZhg0HEwaq+QtNvUKKHfYe+n1pVbliTV52nT7G55LGNe+dywFg4I
oMWKJhrtoSZHV2A8tcoJXa1xkPSQ0E6nVqw8FUMAJ8rYKaP1BZYILgU3aQCYRpPc
HOWrcMLyk6+Miuet3dAXJqxSvBf+px7Ojx8WIs1KQSkDyQW1m65G5H+dT8Pmjynf
aIbl1ttz3POGM05KLtkbu3XpRpxAtrhsh24q+7NrNbtz93gXqCEUnX7QXcz4N0VR
MDaD7fvfkmKxBdEfN+S6u4fGpwseQ43dM77DpOKyCpLmRwLu3zX/5sUu7RxyBth8
NXvFI0aj9yOvJkI3Ev190fE1gzhsNPUi69SztDJqu3vPERnTD7QwgvTqbewx9GK3
NwZrr1EYJp/J13Rl5a68CBpAKOKc/IdzmYzRMPpl/EiyLgEi0ZEe+IoW137GFwav
JJ6TcYgUlAk3f/Vl7qgQmQPqFovZyPAEZQBPuRkyIrRK9TZWJNv9+eSe2VvKUpIn
E3tjg5+yuZY3bcPOSayGCBAMHhQckQks7Uy/VojjmeMRiUVhan87pYutfWEFDk5M
xrIZ0bF8nzTT/hYfaRo6niUqQzvH6ydAIsBxCkBMUM+ZxswfYfZ+shDZU8JHqbAG
+NTix0vDdx936Wt0wcgdFdrmGcG4O3aOl6JZ5f0s2JSvJhYhRnvPOF8itYq2mN9C
jXlr82sY6O2uQ21cmm4QosVyPspkTLjeLPTETjJbmFW2WRUam/9jTZiG1ArNku0B
c5afdBzIq1onyyzybuc1Ko6ODZSKScE7Idegpssa4FSIK5um64hDjGNGNGSTA3DX
brr9Qbkd2a2yf/8/afoCEJWvAgi9dtRPrhfv75TjV6mub9rSEw8LN4m64zM/wn5v
dxfF7zUIm3QiLv2e7yeQvS4GecM5WqJHiVNMVLs2U40PpbbJBC6bhsQAwjJC/slo
Psmc69OekxWuEy8S5G457OP5yhU4FLA4E58PXwnyeaV444H0f6yLfQz1RVh3g7Tc
BUa23ub+T8vP1C4HbnMCRvIGMYwaCiNiyOJq5Up12IL9rPF8JboPTsffZBsyf5oE
MQZRJvtM25SwrM6u7NlNYlSsXeVywayc8BafMF7lEf1JF3kHi9YkUB9a8uXJqs9l
YbK/hc/eDYtqrN2ezlbfmy0sFlXdvFnMFpfwibyk9MAFh1O0XmqjAytXDgkxxks2
IrauydteQSJGar0BIucYcZj2FLwd1Wwd82OU3CTy4HavKVbMXgi4NDCR/6coAgJH
SLG64hLuVBqvZWrB+N0WwNKyxHVAYxGKRqtFVmegPyC6s/JTtO8K7QQfnT59SlWG
IxZ+eMfwk/CZuo+x8X9Mtbu+EvRFq3ToeYXXuvd7xzZUFiPHNM4HQTRRXB3613XZ
JNqoalrrTs6/r/B25zVVr4ZwIscA78xBWH5FFm8P44A/wuyWVhkebQuJlkMw4AkC
3POpqXWTQKWV7OdE1ZvETGwo/8QBWgw+THvtxLiBtZYs/y+IPjAlPCPlKJBHBTBw
S0DH0hI62c7yvY81cXt9qXhbg/OzRf6TGL4JpBVeVeqxdSdMGK7VIeKh2p0LTYbr
sHm7uoCZCUPPd8JQlBr0wNyofokctammeBQTVc5Y3P2I0utA7qveEl9fqfvZa0Y7
efirrKY4QDRp7lVZP+c3tAEw2LKtvrQAcxU/MLEcwYMumyF2WQkz7XaN1DiLTrQ6
vTTHO2FHLqCoX7xZ/O0tunI1ecK8iCHQ4kSROJAGYzrTu+NYO6+oJQpu+riS3Cpz
u4etMBI/waSHJwQxtPUM8a7xBDuiI0mfq87zaBHay8+/OSDp+yGmt7oexIydCh5L
hvwi5nGEvvOB3PbOMZM18VuUUvSaaPCFtfPVU8YCAZQPp7LpnnpAOZhqm4VyyBPq
7JuJ5sD5jGKeWuLW5k7Qi6XmYz7ep6MT4MoQKWd0L4eAJ+cFN+VENPgb3SkKA6Sn
joI/sELrpi6aXnNH71GsJg/tTZhDDRLccWQ9KI0i6L41o6C4kUF0R8T/G9k1ZIav
g23P4ZBhYOcwUDpfG/tJ1mjBYV1AHNMSpS2HvMEncD0/KodeyUmjKrvw6MtlDgZi
GXbdsA8jMZjWHov/gxKcYjTgS4VwS92B6fQaiCalYW4nhL4SgO9n0nmV+WB/O76r
Tx4D14zCH+C4iWmHTEMD0DflwoWBsuy4JedSmuNJQRMblGHLdq8yDExy45x/TPyp
rrhe7HjdFRVQzgWu5mrwS36AwKcoKBLB73oy4NjS8KyjI9tzc+AjgLyebwvayD94
uCD9109xh0dmO8GY9fgTfHeV6zvUngSSwjaENVgPWaOD2iPvN7xuuDI2Bm174VBi
fh7OeR8ycep5bq06+EsCbYS9VrGKiFQ8hrx8JP3p0ySQanVCInvOUltscpxFYGO+
yTABOIA+aDTOdiAgzCC6fJRfQgFJzIzzDZfsqC2kp0lCp3AxDTUBcokZhaNlyD1w
xzl7QdKulbJitudVzIsw6bhMurpQLrKQ2HjJkDKxD7YNVztE96bLhbwJP+iI9I9d
pKVZ1q42DWLC34M9wKzDUv/vNzTy1OF1ikCM+feL1R4gbgzl/vtcije3IvgVh7RZ
TCfumLKuEg0qj6e+fXlGkqnQ06yLNzDlqAzHjk4MYMbmVH7GRHUzDsLUdUbaPtJc
A1tJ0w2JprY3zq21cYZFGhpKG48OTB1/PhO9BxJas3Mtrj1MwHMpQSFyJAEcGQBj
2CGXSF10x6402RzO+6QOKWIMGoOGVPI9N/soUwPZ7TZi7Vc5jYcP4SXEdMJ5FQ9Z
QBYuIePe28XLLYSmZx6IL7yE4E7t+qR12leszVWxnoFGOCQjddYzJHmbbaWdeW+i
0Y9di2LYTy87gW5wRdcXboPuyFQfvhgqyENxDn4qDYpQwe1scSXhZjAk42dIesCQ
DQVvXRnGxYw4rBPZmc8ryna8GCojyoW/2YrM+MQ/1D+H+++2czCrXDVTtgd+eNbl
4uzO8Gn6C0/yit7NGNsZhzQuqIl0YGYNit1qZPGieGv5DKQZGlzTxSDeYy4IQ841
8P0L6JqULnq5/oXCYzx8Bdw6/pJ/r2xAyu91ZfUQJUE4iiIu/dIyrGhybBqAGq62
y6MnSahwEYAlgvRN6SO8zacB/3R2ySwW9KqeEhVHlysO4H8nhIIqUcM/lLJKkHd8
25B7xk+0fblJ12reLm9/jD9yVfUZahrmHNJhaNyOKoATJ79/r52PgpRu3mg9uJEK
fSvmzvryWwK9AQQcv6SSywELFpC7cazuf4W7zF4oYd5kkyhYEkkzosdQ7eG391mf
5frx9J6NSTamuFzjMs0ksyckbL04vAfJbC0bxS6QQe2gqqkl5ILjnxeVP+4IiUkm
1/A4Z07EkhKat96SdNr6sGgHgTZogos4RVuxAmI6Cj39CRZP+Z6HYbHo+SrfNHYV
4Bfhhjko4ZltAHAIP3l2ZM2EN6GT/N5L4/U+v2b7fYtTkh40zhUrVwQozBGLO5Te
I/yrTEVyCj3rIvzxjbo5Kh7iLJmABpF0N3ECa6hIjrm8UFZRnvYCA15474KDqpTC
jC7oFqy5tDtzoFFXC9v63B/Pxi8fRryAIBXcM1wHIokdsachUKk98d/bas6kk7dv
AyyhZRaSO4mhUbZXujzvqAooKZA5wJFxI8NOxPZ1nnZ03UgrZqkEOWWcC0khjSu+
ryl5u2tdlllN+7JQoqszGZ/IB/DirVmXy+gB8sxD6R0=
`pragma protect end_protected
