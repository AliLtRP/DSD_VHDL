// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:56 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
AUVQBiTngXHKPD4SG3ZOiAjk95/0f3tNAIk+i4fQErNIRSnKehHvjeaZVFmyZfEx
cbdsO/wyQnibvulUVzoma/vi7Iki2o2IuDkB8dPuN2e6sbO3cxUgxlnNF9DpjJFc
EzrbEWox1qOI9MB/NOLts8YA/oKJe+SSgfRHcC/GO6w=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 11488)
w6EJynAps23+RPZCzGp7Yc6jNTBr9yS/+4vNOVvINek1U5XtTOvGnkJkiuZsTg7S
2ZBHC7XHa6HrJRa3xJfkuTMXMJV/q6I/6Kg/mMN9vD++xKluowTARqzd2ok7/QeB
yC9++wyE9m9NnLXDv3k4J0ZXQCFTUSsSK20o/nzV04TdmAUwytbktcEtGBBx7n4m
P9iZ6Cbm1YtlebiUU4DT8zQS6sphz0ljUxbfP+HUAtKFKBU//5XLNz6UD0mVzb7M
jEnkZ67E8s1tOtGtO4pEO2iLx2dhxWd03Y9Wb+gvPHwIBp/yImNQPIRmwp5TnLlU
yZR8p6dYcyvP6hfPLSVCewEokTbseDHLHAM/vejNzVLp1zVkCTI4bEdNUqvpJDcT
HPldltu8cHXp2fDYcXF9MWq5Cr6koFV2WWuIKCFikgcOlwpOsPgK+1cDIDbNH72Q
UvxHt5N1BX2wyYRifunuXRJuuOiN2MgnPKeqYnd8tr9RdpnbtNy85lX/xuLMPwnt
NXaJoXVom3oecN+CUmx8EYLXvRS3Z+JHz+rYgapDsPXeGKVCLidJvZ5LrW4Q1DcT
+L7e4SKMmWw7cVjYVd/amWsl6WR2E+opBE2Qo0AZdn3sfvPxIHmQY1d2f4PJujaa
eKUS5nDbIgUk+nJROvndUtrchdweYk+9rN7BPcA/k3CMpwo0qrhoTcW0vP0pOGpq
tJXBhTtLsyca8UmdUHgy4GlCquM+l80g7Nr0NbYgzdqo54gksmOuiLXb1ECwCJ0r
m5dLZVRwGlIzQZTZg2/7rccbfwkjzSyB2Jz6fkv3f8nY49i/ElKOROBJ42lX19Qi
YoLhTY+y8v+vxTkm9m91KygItjNWm9I+8h+0BYRFUUBsOA5VoGw9xhaWbHFn9QaE
8NHY1a9k6VYiN86oClgPO0uMqa05GLgVshdTEndev7dSDbiyMztKmaMIQbFtzSxm
Kxqo3/vopFazma67b1uHWIDK1aJxfcGBnVjWOxQYzenVTlTGvF/iume2lTXM66pV
rQB6BxaD4ERI4s459rV6WY5v4ywhQ/aehK8X5yJPacP4Ize1gBZwacJs/Dq4Yyv6
i8lG0Sjp6x0MnD5zN5BhTYMBCPbeSwD3vqboQrmGSutHRP9HJ86P2nDnI2x5WRGJ
1jeGr8ACHsgctXUdhdJNATWIZQDnXpMVgN7Lu7EEYZDB1a6lF64xSM2lYDTRzbMf
AUhNfR4is4Becn9Wm/jsXwthOfTZJPZ/vF8Fs1/Z/XFozU0AUWmejDnHthHKy+74
cKtIvFWKPPuqPq1WL8y5NraZR57nys40oWtuwGo3PMrIo1PpRZtgpimHHzhByRvg
9cgk1y1N53r9aaxT24Z3Umr5cliDaWHMd2Kc/ioeK5/nAe7IPJE5e6McO8rvel6A
kRMp38j8phB5/JXlDnOI7GB7OybvtVw5I6sVW0vT8wrsyslmOgrf212NqihSKPfM
XJ664rSxK4+zAP7Lboaa+rIFynx1yY/An6MJRW5a4RoSHNt2FBFwpCokeh5vpefG
qXcZ04NbI6cB8WgWpJaDyN2yW4ICPM/nJdZzQuTpKey7622F6MbakBV31eyO1fui
tE0WtSzw1vcLfJzCboItNXwjJnnCHHIqBl4IVTuYLOOM7KwYM2ukEKhQtK0bw7TM
N5tVd0qKH3BwoIPlWWxmPVWKCnVdwU/gWzzbYxi3sZLhauu3Wxfilsw/XEgjjz/V
5CrP5q0bdZuGuBo4LERq36vO81LLQy0BZDqQM4M4UkwhSIihRixQj0PJJCFPr7xt
CJqJWcKbYUosENaBb0RPhXbQAUSmn5yBq500GwH+JarliIdSVU1bnVu9g2ceWKtd
N0t8F+j7+zKWL3Nq8jqxc715LYwgxSUJ7wFYouIbnUMfHZNO2rafeG+Ny1q3Ow38
VdkH82UjIvMSqaO2I3ZFEEEDPGlTGjVUD54yqOY3nyTSbdDVrnyz8/ogDbiwqCOd
S8UzfVw2SDXLobfTItCMYuL7lTNYE40X0IQvY5/A8bTItr7MaHrBSWgQMZ0oF1qg
Vxb89Cn2tt5/JkXKBpzxNmCk1WSf27kTpG1f4V6NMOITlOuqby3sIw+nLZSrPXhV
hId6fU4rUGU+W8YXQ0qMAFy8sBnLQYEDSaixjxymr1Rx5CEf7LDt6AobRcMthH7R
lSGviFMwLAqAP/Y9lXPOHEF/tRD602ex07KkZFvQoahcdWawSRXB2BQh6m3ofDo4
hlB7r243AhOOKtnUp4qJ75pyzpyxr8XBvayWT+ximhEosMb2hbHYpq9j+A7d5G6b
Q7svO165n1YvoOQ5QLaPeR8jUxkLKrXmEDQ1Bkp0FQxCHXwemXDJfaofGU55FwVM
WK1KXQzoyq+W6GaDpAEw4AXf4frhsyOLlALdEGj9CQp4hJbAim3ewdBkmMpgHeCl
OIL+SJU/eAFR2ugzmyZAXxgIyCxqhJAA+lRw9WqYd5tZibrgNjRYfDRPTOsAovep
pjPncDnjZ7fqoBiIf98q9dR1EFUdl07EdjJf5Augoi/BqzjZ75XOrRVlrTSQ4npS
PS3JpB9LCtHi1mBF7BCUCsfn+UDRHnyOkaJXDScqP9JmTgrA1lmas3WisdkDeCZ4
4ObOal2tBioEInGaXqgvAKTzgOE/3mjm6/aMdiSkvQD+grVeAf122hjW0MwCgB89
URI/SXkLIswlUDh6Qr0qORYS798XvkP0MAsPff1FFrPRzmDTUkQl9BVg+0ikMSw8
GeEssejOez0q+yw6LMF3iXd5vGkubphEfZUVo98V9cSPhL6874nIEqEdcIYtY7Qd
g6b7GQ02fVBzEOyBc2B0XmwFZzG+cy5wPDt4h2PBVFkDQybX2GOFS1jt9GqlYqxZ
7xtMKP3Oqp2JTxAiyyTs1TciwWlCw2iPysdEV1h/Oc4Lz9LfmuBeNEFiIidjIFnt
G/d7mfE3Q4mGxKfUCDpwBNpG67SqvDX/C7mx2ZW/C+U70yQ38rJRstLk6o4s1s1g
o83aJo+HpsnQDLMOHEGZNGJBBu4fZneQs3m7VdBZOczL9gbPQsG1nQdHLoSCaSqF
u+phMQQcjX5IIsbEdxKS8eMZsNPa+Jm7HDam8vPzE3yqN5bJtK2srrn//kSZOQ16
1jh3baE1DBRTMGwoU7M5mUfGBO1/tYG+hxnaxnBy1quS8FCLpxHtU44X8pJ5IXyC
GDzBhge6YlTW+Ta9b38xtH+JeYC6XJsPNAftw1a1zl8SVerfD3lNn8GKEptxSZNn
LCBexZGe559qO7nhcxRwAbPyHiLhrcaox/A88kICrZ842KgpkHh9ztZFPffjSsvi
zefsNHEDlcXekm5uCk9Fz4w1P78VEI0sMtDI0uq/jU6Rl+BLQNPdfElGqrK2Dnnu
Q8Z8PcazChk4WTAXQ+1U9jdwJIhEj7vg9Oweep/WPzcSHvYMxa9OKaPx+onKH2+E
W6AHLjm1KKcy3WE1rK1vBdARQy+Kg+jfRoNcKn/2koSqXP/xhNv7a0/eviZkS8KC
SCVYr3Y3iZkPkqVSHwEv8RXUMP2UB2su7PzfKwVMNiVvDQi5+NkYezmlPLi+6cmt
wB+W7ztZLwl8yM7CQ9tql4nLAYWCphOQeYr+l0nIguaDIHY0CBFbpREaRUwrcmTt
CrhNg51tn6aqEecnrjjjBfh7o5ILjZIsoh8jXgobvaGcCkXXaHg1CUlBrysa4Ecz
Ao6RYxOouRBVBs6OOCdiOfS8c0v9+kI3/63rDkonEMRkUYDG9xAfkrVhCMD1T3hZ
CUlDlXMq7TQYod8YxYY9xaXzx6aBaRN/ZSYEiCwzEz3Nw2dxYmRpY9n8Gc28jw6D
xGHlOTXZyLLU0fTjfSwACOYbefWFtVlOvUIQRl2t7Yl21CCwFQZrqGqPrACV0PRe
M703rrQGMNzZHwUgutkC79aW8G5q5zx2aRXyNl0G7b4cYkyS53JgcsjtchQeF9dj
XZEQ/RLnRzie8RCBVxmwm2ucais2iF4zI2RaTlxr0cEdf8ig9SlrtR0Z05CWmT2A
gFAERrQcSywsglKmw5AfaK7lNov5d5GFFaWsHaPVHoZdh9aQ/kVSHA4CFkJem7kP
gGWUVV+nxPVl+CjGcjX5C+xpv40uwKhSz9QIeFgtHHuvDLaWp2LCUjRQWpMGxFRc
ZlkHzP4bHt9nYWTROgDU7XYD7kjRAExp9aWU+jSpoORMMKb1NwVDl8MR9eX3GUSk
5kCRA3BkOSDXXYL7PlhqVV0tcgfdjufwdquZmrSpYT2+kWCjWxU/RAty5zTZXx9Q
mi0LFXqvG7flmzsc6U/kbcJU3ZxxVdrIi2Z56RUDiNdXjqCz4IXcZoqj7Af2v5k4
BqLXFlc/RiwCzBTgMXZdddlvNdUi7yfLXEEfl8/ir8PCVj3Jo0yYV134tQzAaVg5
Q/Z5JTh2R9Wn+xan6GvARVY3sjtjXpo3YmCpKgx6fyVwMktMJasXYzjN9D3FhivR
FRn7NU8vXWpD8iEaFIaqs1DlvyMDf5j22ejef+JGublvOhRKZKdC8EYnznHOCBpf
ah2XkEWGUvVtdoO9x/divzWh/pH1x4sH/8h7sqx0uqWv2gBhKkCM6HPo3V+7frdV
8Ioolg3d9hTpc2d0VXxQFr8XI2uvZlpnv0jOE3JG5qqqCO6npVxDbITuMVo/hMv1
ivUYSG8Wst/MiA56aglXmptbZpwZuDtISfZ4fiJcG4f9Ltqy5+Kkmn3OLHOrzNm4
JkZgOWMS6LQQzR80WxldyN03rrw8bW5jBJ+RIJ+zmCzpD6BbvEmZ73ZzMEjqY5FB
2ZfTvaDsjZhRdsODj2/oSB7MuDfOmc3ExXKhtFDKE8CcuyX+KgtYWwX0w6ctoQuS
PaC+Ytj53LQJkTVJ/lWnw1dn/RB90OsglPAL1FgyLWNN4+uOu5v0cV5xvGQd+m2A
8qKiznidlNz84NdVJLYEX0LVSoYp6jx5YzZSZesMFsMlCdJtvHeAlySwb9ena/CC
Bpg6G+ApDAo0QPIKu75NTB+EmvrJ5e2y8fotnmc/vkEvAv0QsYP3yz++fwnEqJbn
hY/6il7/GYPuN+vF0pWLScRT4GjVr+S4289QJaZ46B2JOHl5/9xzmphCXQcbXopM
pVJm5qhH7v2tfi49UeVZ9cIX97KDD8MjRoJllarsdqCqMYmP6Odd1rqcCTe2xS04
KyBPsPHXiq9q9GKTDwCxUG2CWy8+gJFSH88gSHL6ICeyO/aFnvO8P4ARr2rOl4z+
C+DooIkr+7I150oKb5lRRflO/mSuhtHo3eFnTRmGtR9xepy7IoOR3TafGECiCoM+
dtOvBU4zYyY3XoBZcoUgBWjHtMTsjPIrVwCnl50Kyj1KlQkp39zmavbMHQ4qH4rw
gq+HVZgzZxS+a72/zcw1tJBYWoRTATYvViLNIMnzG2iAMVsGsXTF8bXk3pfPmsx7
m7kkiSa51xP6icJtwYRV/zjEOxe8c5jek6aJWDDAv978Bbex7iOA/yCYqroUqKHS
SXyXzuars3wh1/WvCikLaVGk1alob7PrbVfQ6RcGboaH+JjGJz0ys3xw6xR7Sdic
zIkq0BbtxzZv6J5ndpJXjjMZ6XBXT3vvaePq1S+o8sw65mz6q/T5CA9wa0XN27bW
oyQW3GHtDvvFXRixkXhEmxeFRNtSLjH1evcQet13Nh/XgAUt4SXLqOKrIL74YnsI
T7sI9cr70hJbbAhynEBfqHVmYEvvNsQu2ME+cQD1KX95UbuYpRcY+O5Kwlx4IsHt
VHPoxq7gCuVYsZh3hQU7VxjHLFC91apDHwikOK4u33+nB3eQDomSZl01rUb5c81b
8RxMMkJ/KARSJbtKN1ZW21bQRGF7sSPngcCZm6VQ0IX8Kh3/cZdp5JZbiS+mflGk
inyxjwqXpUl026PbmVx7Uya/vluH6+kXQ2yh413Cc0V6q0hL8ferNVV2mc+n0D+Y
38OIo8si4ur+bptSbgw/LPhhqKazD3BfAz5o3xNvE9sz+r+bhOnCJ05lnTPy3ooC
mjSXfY3+Q8ybs446xYhUzzl4VcpiVIiXsIFuCsTj1doPsmJemVLe9tmA6v9kKRgy
nTsK5yEiRbB3rmH38wvfwF72WAUQaxNhwIWj86C5rHAW56AWxJpDjpF/vNQDKYYa
BcuiuKYUwcSUk8S0ZeiX55tVUJ6LnI2UfJtAH7C+Pa2RC3uS54qlmqGGZMCRtMQE
odm2uHsRtVD9GMrQHPnU/y87sLfSGQJr2sHkp6upqFRiID+L58Tw0Yu15vhvXjF+
7w5xVsD7nwFIR4+F9XWd/6h+Ezpy+WB6DwZcFptGIr52WkbzopU44j6L5ZW2pRB6
8UrUtezcJqaReo3SqlxV0SuMx4VclP+TH/sGBnFzl5Uxim6ufTy3MW9T8+FIBVSG
iod7N57RMQpEeiRPlzQwAa/GZu5UtcDLHfXxdm1ZC/emrbKm7KH7TCs0PVJ3V4Od
PMEJRkClbizCeM0Fo01qWMaShxNXtXLUvFaHEhjpIhQSgOmSd0GrTiLreuVhX3Yd
7TQF31/mLd/RX+VeS86kKW4bXrBNMttNUDcyhaQECoiORSciettjFr0GPYHCemOz
R+xQmNzomhZgaHQCWeS/Ll1A32B0mBJxFF9/DSVYGrIC5ImEYjLEXm4VAonkTGvr
01l/UpEw00N2HZr/fqi66SCVkVHhWsTOP9L4bULp6wDX1NALKSYDsTxibJ/bT1n6
aEOGtmuV+AyqAFA1rfcTaqY4PKcvToUaNNkKGDzQoafvLq01r12WcaOeK9xYgiPt
NBWDkGtnU8a4C5BPP7GUbupxYTIll4PO7Kdk1fsLg6Oj7KIsTq7ig3K8EQTPQUqZ
eMJAr0zNB0KDh/pmfvDvZk+zD192vKwHSYtCZiPrET1yu6y1MtU+bKbfvjT56mwj
mBXeux4xje3m3OqfrWL9D0ytPdzg2pSqsXPHqAvGS5RA+TYfzDEax77ECNCo6OHT
WSaOtpixaRFBEf10ume8/Hg+1FUaI+XgEPMdeenE0vsm+BxsLfmqt6bMxhlpj0mO
pEO687yqMNRofLi+BxHZjV1ul/49+ZtjnA2RjtBrx+mRs+rwTm0cQ/lF6aKvvDoU
/xvgUqSsb+jfHCTy1Ghk+XymTdB44qvVhZK6yDpcdRYiCfjSLPmpMfqd3IjzjlF4
GV6smabn18qcLxS8TRclIWmPmhGXioCiMfMClpNgvZgGNmT9fHkXr0FxCTMHkX3L
cgfzxbYF/w8oypXAE1t236z3NF1P/Bl2Uc7IQPbhQoGZPMJOzR0ULZau/822+VHq
XPxrufsnMpwxofPf7HZoEz5tkK8wOTwjoLlHkFpkOn82ZURGv8YYQz9psSSpFMLR
O9MqlmJJm7yvD+exgDHNV2F9bL/rjPBcKMQToUPWCzBGbxKg5owsxMoYqQsq4k4y
VKAzygXMvPBdWRkIi+NUIJSci6eRkqT32xC8SeVG2jtG2Dt3SUI70kczhQ0WCP1U
pV9qsRgYHc7N93OWrCez/XOHsDaumhRoEccgZU8peClHPk4trKFE0TAQ7tD/ddGA
X3BahVNZBxHWX74xzUt1UyYXy8ZnuS00vb5YICpOWXz6GKKMp1Lhfye2d1l+jc+X
pgh0DO2iVbQA/Z97s6ghLlL46SElbP1isSzbYghapdWCnpC74Xa2l7sEK4FmiLaY
P522VU6oC1cF+baV5AcXAJqr8xUSyRH73xHez3YNgJp1ixwFghuXCfOngbf13Ujk
citOJHZSwniD9dc1+fzAjFD/Be/86pK7hVF/X0cstkuVgd56MHhTGTQ92DiJNPPm
hCIZo2SMy+QniqsVN4Y8gWkiz9SmSD2/CwUblj+LXsk3nibPHs6JHFv0l3JBytfv
3NJ0sXCl5NgMr8MMyz8/nQeOtJhYWjKMhpOV9M8TMAF4Kf8FAQPKpSi8ov4orknF
J6sQkr91nGR9uZWSnEEk7UuJSTNl8z87QhxrO0HuqOrxBA2McMFD0BxI/821v8oH
GI9T1yoH6UAGyVJGK6CxaBdxOAdXMO14znIN6ie+Pl2j1+t+SLdwblYfde8KoT1Z
AMp0/sG6cx3USRXDcHNCvNQaMoBQN3KBHgFKbuUuAiRzX8b8roPVd+c3kXt/iw8C
tKICoxUAWFujR/k77w2v5PC1d9F8jS7mcaliBQTtu29IIf0mh1jmU1vtK7kw3Ci2
RALkymjtswjItaokI7PIwoU96iw9rKUfJ7c5LNAryVPJos7wdHdzyk52iUVNpPM+
voZ0Bi8u8tC21oXr8KulskL1oWBGduCQKIRXlnXRkYFUN4qSn8CP4bbFrULHvKrr
/KTbiMHNowAG0VraC72iUn7rjyb7+qWzx9jDImiteOrTTHei1HRfBFYvuVDMAyJE
hWKSg5DjWOLw1Fj6++AmlQr3i0verrrnVNXTODe5GroaORrllH3WGRxkz2HxCcxG
xoDO9Ydu9ItomoYMfTNPqIVmG7d+WebOt91pjCSLEfIIt1wTUeIbhCxQ0cGB3iqT
13C/cWsmqNpdkNxu9dddPsRDWJpUxjdgQy1WI8bHEO8oA07uP1Jo7QbwQFfo1tk4
7ecfi8020viytc0Pl/2rQBjFFYpC9guiqS2F66xPZnasXTI2us3WLvmLruEAgYAZ
5LJLIByQHeFIghUkF0uVO1EpeQbd8FrvmaErAXhqvKk7+6Q5rMxRdpXs1EwoQOVz
QZBcKHBgroDSmqY2F69wZF4olcOxHp4xOL7kHme7WTp+8hnJpAzxIqCFGVWMk0jk
RQZFiHi4SmAzsyLG41yYALwsxstSiqVC4RA4xwjEjGzXaGHCtVT54y64ggJgq8wM
zAmMnBnTYZRPSIGOj8AdnIz1ru+yM+0uL/hjC7O9mXVgR/uZX69ojvbeYtQCrMmK
sZsE4LLc1AVk09nC8VF6MDlPzqkdASVa+ah/HydqbQjeUmrDjqrsjdepIPL/anay
7XUVoAjzHd/mm7UO5qo1O713D3TDS6CACM/hh+SpTZuUFR6HL2EhP9qOWR+AcjVC
9n6XsT0XGixVVfTf5/gOzfpIL8TzbxlAjwLkNXGb/4KirJaLSHKq0jLmJeGTjAKl
oxbCSGkJAqs1DoHTVj+RfL2VByNUlGGZHbBNWK3xFdLfVTP7g7SYe9MM1glF4ND1
g/UOpn3xy8swJPv9kEGNpxO3uBnOWxom3+Nb/KESKvW1yscJpVXzMBZ25P/bcfch
N1OE3csp25HgbsZasMJSu4b4fLRRZctkQYujOr6ormPTtcNUj5Wk90ppM+QtUENH
VPpTeuPPro3uIVD0JF9QgK6mtgc0KjG+Xgo9AEavNacOKPNjOp43HaxVCN+4ozhq
K1xseX4CY/TpSIEcdexrltZqWb/tS9WJfHQwr5ZiPPROSEfgCZ9AaGqOrp2cL+BM
46bdVeiXxvFg9qVGz8BNojCbgVYr8i2CCOp340Xab9c2kdodlXB7FnrDqb5q5Muy
zmmpySpMzd/wxWN+uktovuqs2glR4v1WN+RfpSOyKTTQVrNRRB3WNYeWGg5k3nCE
SJLIVV7+rXnFQVOvS57y+Sei/GdWiUW6/7lSsajfEK4NPArR9MtqVUDHu+XvfL0L
fG2mU+Cf0bMTI0igu+gUpv4tZtBRF8XcMfGkHinGJ+OQRy/6DXAyocvO7JlFeou1
zRhkj2BWacuV+Ur7Gi+zff3cz5Lp06c+nqIA5dOKo8KfsuoFFdNdib2pFPhl4BY/
ATxwbJhmu5p3Nz7f0t2MJwdo9sckyJDnT2YD9n1tedPAdUoQN+sZgW2I08SKyjdS
7w4KCprFuUMWj3PYKZD7Gl0Tp9SlSkMSmymsM+CPPkJFGGMoIyOUQA6ZxDy4YYJD
3mQSWH451s75LdUO2s8ntensQEFbjPIhEsmjJyAhqTsc0gnMp+iof1+RGmrOOTXj
HPoEBtndO36+ex9/0uyef0uACzXZo+AwIF4nw9q1gUyy20hyOKAXA2jJsjszSEEn
e9UGbJSk34iOqlJTxbv9jagEx2uQpKUvvOThpEfUA28TTsSjLHr+krEFAjY9nCWC
0ayEjZ8ela+fSgFgR1LjP5hieU9yDt5WV2wGhMPwwSDiJjn1B2mVGKGIenlZ5fqw
7WPS1QfEIgPSs0+Xppu7ownEZJV/OSDWoKTKTp+XrLSFPaUTUB9Hzz+9VXztfAcY
NzWzZ8P6Uco5nyDEbk7ef+yx3ZfZ0cME+nvYBkCnouosm5Kmqw8dETz0fDQIRBnj
mimJSJverumbMOBYnpbjN4ENvgedxuZz6ReEZiD67ZfPRLeO4Zm3/0dW0Z5gvna3
BzzGgFLDmcvZ2Z8PRSWCNILjvbvZ5Ro6gYcJp8Mmf15vusPOn2XyxY4DB/NLUumV
/qyTpCByA9vmmwY6iHbnrJIy3pCSxyCm/mPXALBxMpWZgCfVfUl+RH38ZtimnQSm
mJBabS2++bgHBhPBXCNNjJY1vyAFoyghPtuykjkMvCPDNjr29D8LZfqF12pDGNZ5
YC5e0uNG4v/TkMr1jajwUd820mYGpj40lr9zZ7t61wa9aQMXbMYjqUJ4mzoYKPRG
WQKjWMzWVuBo7E2+/DGld/SsvZagcjbv/5Ls43zo/kdqml6x2+9vZ8X5T/K7oduA
er01ZykpcIdXIAXZNxtJFOSaU341qm8qn7L9CuAISBOjDznwR28Na3yPr4CLZCAf
NSqKpTWDlYssSJqlurTv4LWH3xTm5SFT8v4nSBjxOp2C1lViNQxBeuuqNtjKTR1Q
0cje1UsDZyDEHZzeloRs9Jp2YcK6KL2H57HHd+azWfmJLm5jIf3Y/UYw/iixmmoc
+OSbSknFn0Xko7o9Z3IBkXlYkESDs9d7JM7sWcNEI5YDKxFV961CENzJJzddjz70
k6YgY0hhLxuXLdqYsOvn1D11ZZ9vP1Fhu4aJgXf1sUbUQBin9i15sKyy40bWGLoc
BaU8+uCdjUJMyg/d1qme0tbPfXvROVhAgx/wZoomFWdfs1k3ab203TpyFbLiXg7N
AESwKkjbVfFrnB55sHxsWNK4jTGlUZcZC3wix5cJsFlgWMx6bp+qqrW4OukcVOQa
UqCCF05phjMnBFi3YOUo3cIauoNKqb5Th21X4j6NbeamY5WHXFrSICCTPIzmxzrv
NDWwYhQwKSUozjN3YpxqS9cDRpTMDC8W0+El00HdLYJt3pZvSbJSQosu4Iw2i31T
Wpm68Xya5bbJxGqST2tm2xG5R30ziTwDcGYZds8tSDLmnOZbxDv279kmaQqlxBQn
gplDZGpa0d+FQ6sgJec95J9+xsiQV4T6aON+3VSLOqrsXOL3uShUJWDzM/yrgVY6
r1YZ11dKF1/jXJ41uDu6Zvw/WhwDPc6uHbrD+ZSpoeShKgxgR6fEtMPj9DSGygur
vkXPl5ZDvHxnBxK4pwnuJwg4tlh2C/0wjuwV3fPvLuLizOPEFUlGfSNc/6yDAoZF
jZwWlh22vbZ2rMQYDPCUi6yjIe8mp/KvuxtT6iTxhjOJRxzhcU96W7tY/2cecZlv
QowRzJ6Dc96a3u27lnAeVUtKaprhjRAe+dVOTCQ5gEiPHytpYbpaH+k/6qjpNlbl
IsS+nhAnmQrxh5awPRE6JM74NtKAb1e/peIrdo8yChzfB1lewIBM1F7EMu+e9Pf1
2JpjKq7q4YELQiqRRq4JysVwRWoEzvxvyQays0Ss/tG9DL0s45wRFXHoA5h8/hbv
6/qPTgvIg6ftqyQy5B0n6JHO+bl01Dz7Zxl5/7IEzfO4uA7KT3hhhkfPTDMotUWr
j/pyClOUV3ktC9PSu6JcaLzzN64dcolfvGJd/pJh5IGNJ+OOpvItD/Ogq0LVrkoN
m+OPNZKl4Fdpnf0Ln/Sm48KyLI0WrSjcyGSOZCBvLFrpkctKJSeHNx9Pg1HlPJtI
e/qfO77XnjBJhMRnQXzCFkp63Q3362IEYQu2jFBY9KhZ8uoRWr77+TWDxb3jvGmd
LW8J5zjXoEMd3jKxx6IdKPXByrM8zcfgP0SxjFlv3KwfeS0VIvQvaAzze6RzQNCk
p0pfbG+jxWiARHRY1So8vBTtWq6xfPBIJHxP1ooaSYa8pqPF4FWv0u0Xt73gv9ds
vKTGnw2mGY9qKXo3jJErOj0JUgsDSuDWdsM5quHetzt7E2a3l8rWsvJ9kTbgQkGZ
fmIgm/oB79qrrYLiEfVf1U4blMkYtdE1QwSfviHFcF0BZDDujB5hkgvhLOcRWQYp
n1JOI+ABCn1pcDgxatch3XKsyYOzMxT13YjN/o4de3ocaQhTte+X42r35hNOv52Z
VcDVnvB7ft2Fz4NwKPyiMaQ5ZOylYoVHI6p9czCVQXy6nWhAbkUwqDY8GqgeUuVU
mU2Qs5u16BD1fuKh/KT2sUmce5DFW8jBoENuq1guto2geHJOWwvgdyglMgkM0QUZ
F2Bvd+w7Xfe2UATdiodCzntBMogLReB4vxTHxxWrLGot3Nuju1MU+ieHce2hPyxq
AHFSDtjIZOXd+bsBc9MBjTJ40PRj7lNSoHQGozXbmKjQsbks+t9Z5ksGmVKueFfr
rdHWslRCY0Yr9JOnsIDlDrYKyLz65SNfUsBtG+BDrgpLnK4kpe8WtaM2cTocjm0F
9SUzxlJ6+/H1wRVBhfELNqtw/GDLpfwVLtwZttuzZEtUbcVox07URn4viPQo+TRo
0sn+9xVi3L/UtrfX+HItxMnu2QMWwldw3ODkilz5Go7qG/TshbaU9BRqzMHvXjZp
toYwjvGShOBOKUdIMY0h66iqTd7LjSCtvrXlm8LMmLCR49LFLSh/EF+gGrM1gXXU
laXpPMeQMAXRDws6d64xAF8HXctfu0ryURhUCF3YPT2yqmYrqTQWJ7NBhnq/XJ72
OX8BQroioM9kC/yXb52l9vheon8kEOPvPYTXXtrqy+mw1bHnP+egC2aVHnT8j87u
Tu+Tb+jkT8NgyonXaW+qKywNkIBKcbJN/IwAM5uffvoB1COOhRU+nXfG17X1IuHp
Q7OFZWlFYR2IezgwB7gI/sLPDT72RP4Rlxs3CVuNoV90WNJu24w8cvuvC+JdPtdJ
uNeLU9E7jSAk2ozJ6bxs0pXWrOAq98A4Han/o8lHYDjArtpC7DuxLHwnbYHEz0Bx
VNCAOgGOjljzJlwgAGP/6IVy1J5rmABAhlDo6IymzaZO6hqTVZHQ+y4B3pDl9iqh
6MHRRTdD8/AEtr1YF3ugPV+UjW+cCe2Sm+59Rzf0cIFqR75Z0qSIcjSA7VUcAJwB
tpN/UKneQHys+yRjJk4JLYsX9wwNDRVwwQAqCNoxZp7JNKd3NoLnxXV6b5+lyKmz
aH0SaGrlsbTgWMVhDNzXDWUMN6rWWZO44bVNbKFqQ8iDD7uULulO6CPnWNbbeUec
fR3q2vgOHHR/SOQMe4zDRtr2hrAJe2CNoH32ZEGKqhO+yCzQonv4ZsjlBAZap3Sq
yOpfoeqmtZIIDdpSemZIq3rfP0feCdnBh1yeAitp50mn1/AzGl9JUVplyKUXGnm4
nI6Dn83IsEr0xa4DOy1bICf1BhSWq3GtsiI7Mj2fdiNeEZ13RvzquCQepaTa4Dxm
FIXxdKPoDzc/PDK16GIeS8KDWcbgI3DiV1ge06YUVbyECGkkoMQh24uqFNsgi6ZT
As1D0nQ+M2ep6irkOMkbYH9wmP8sGGHYNsHg1S8HlEyeufVFxQHNmPoN4L5Hq/BW
zXyNMIl+2lg1VcWogZUqb1styWvvK2X6pgXmMkvZkgqGVmLyaWLYAnkbhtMC/PLI
Vrj/Ga7RwXZsix5hRiCXxLOpSM/2D27p6QlqnuzO8RI+c9vUBQJwY4Jlu6iFBKpV
uoW+C61mDjRzq1wMMvS+Y7Ob4DJwxVCZQ2xKiUxBQ7BV7gxn3rMQCBE0mZiYtth4
8TIb8pe6/NfTcyukUGzHSH4YXF8nppD3FaifCufSMNIlyvO8YhF4Rc1slRepFrfO
F0dopYGx23zM+wJHf5zLiM7VBI4EAcaaywYrfxwFpmxBU0Cb10sbK39Aaol5LLyW
T+67Cjsj2nSVMrAUmpv8tAyCeCLEAWrG+PzpCATg37pc4QqTRfxDQRaS3gTIlkIR
bq3BMCsFqyHq91lyKQPwo7fAHfb78x+x/ZJ+c1A4/pdtcexu+5Is7ufo48h58Dw3
BqPAIQTD5iEI81jgSNA7gsAd0M/fGzmoyRdYiC1siqQQJEKcJZmwuLMfu+MZ25LH
U18YtDoGiOta6GASSBru98pMDQQkOTQD8/YABoWys1FyBGnZFcrDNTe1YfkQ6Gs4
VrGjM3tHg8567SBAZrSjFZESHVZbammSo8SUOtmfW9dDW2yTIgRVIGlgsmyaOhvF
efou/j5TqNcSK0bgqkzU5AsDhmI5ft7OJd/ZZ9Y712g3mC1NHASAV4lmkZGwjIWm
tA90/P7MJoaCTdUscvrm+3Y+SZJQjQFbLq1Ugrvw8wsd4SO8MoczFVrDM6FnR/lP
ECkfoMRhsZVO8EUET9yHrsxQZHwo1kGP1iIWnhAaWJjptEgJ2aojvXYQeKfMFZbd
4LclTLoxcxG4LSgP/WutfPzm+e91OD6N5kGvQ2+JzGqz/QAZuqCqQ3PcnhxWES8A
LPD6BDrVfg+0NpT1jZ+qmeewSXOcjA33mhTXVBwVbHwMnTdQXx+gXMCYgEJptLRT
NzGGxFsZmUvpU1C4JD1UUjGvJXD4JfGKxVASXWqw83lQydX7ZyRqYPjFDHtsCeoS
2kRDrYSqnEmSdKk3veDvpKasVrFjDtAzRgIzGWDpEda4ZilyBuKY4VPosgmnOjgv
D9NnvultrRvfSBdnmkrtoOGQVZa4ieoFi2AHZW7X/yNTq8/tbZYIBOQrivjFiuls
0+TDzzYlSh/KuX+kiijA8HcG17dxV3qXJTq4gJ4kTACtJbG0Xq7wS2hlymery0lw
C8rjnno2xTAt5wVi+N+Fg0Oda7v6Y/P5pTggvIDLQlf+Pf2Rh/Tv+BQA6Nz78co9
AoclU5KQGaNTwxS9jsrTlSFyKomNcg8pDz90PdHK/tySWSyV20FA1+S4gBXsawW9
VFYMbIQFHolbzYz5RgA+8V9/dQRb7OXMDZkZuVKNNZBtseWEv0lWZkF8GdBbl8bB
xRKU399ktc8WciQW0Id7XYJXEexPtawXKGncm0kZOYGg1Z+aVMmsHK/4MauMpdYw
BG6lgsy40K4NQPTWFkm6nmUTEnywzMB5OZF+Ltqw46VwVHU/2L+XHKpXDpsn7upg
HwgV//1j+fevt/ObS++XK8pqQInpQfut9HGral1dRgq07TaHX923+X+qAeAuJV2Y
DAAmZIfUGO6LYudKvKbkpA==
`pragma protect end_protected
