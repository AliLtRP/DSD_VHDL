// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:11 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Ax3gkhsboV2oPbeRkNTfV8+eDv6GvSKxM8Et29JbGypJ7gikJg5e3+/VM0DwVJgY
zlEOM2tSGLCYKd7VAtThXdgiCpDYcs2uBvdp0kAgP3yLYdkM/RGApLUbsnHwksLn
8PT4YYU6RrtIy/OKXf0nAdE3iZ5Ch8O1Ub+i1bAfNNU=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 21424)
z5YDXVe7KiLI7Xn9SCZf4RGZ7pISlBc3J37YnzO9cnVGHGjgeVcA+ea9PHPp6wIT
6x9NXNFA5QI4umJWyP8efKxUg/fFFcEYsD6Pg56G9Sv9Gq3/TjiCiUjOGOdP6RT5
LYo0Ul6+mBvFUtkuED6JbJnEXzv2kvM5J2SjQEb/ogMde0ZYRhsnCTTJ1VF5p57x
vDQ0Np8mSuKW6FrsNJ1JFZD4VMTzK42aag44wWKpkXYPjPr8/aVU9odSSbXRB/c8
UVSQbU68LrqPcI30XKCioc1FBgw05cEKSk/RnokN8eWqE4xT1vg9G6vIgJf30dEP
ofOZb+55TtpbDrhi2VMRwnFR9qD5FDSyhalht/RF3TPRX64DcFa82yCZCYufgxhV
B0EFvY3nkOEO9GVyMCm5eKm8/B+LceazBt9t1W42AtDjDEAPX8UzYckBC5519fCR
6OIauxhdKizpz7/gTs0+eDFesjksS2T4YL/z5YpEMSxFjZM7Hfa5Cm8PtLMt1FbF
WEYLru5wkjcD/58v4tb5dqdsmQLaFzdFfC41PeKMhLd06m5NtRIftyHJ+ojv3903
UFframDHBbcJx1Nip9FWXjsuGJEVX2pFooWPnkEg0jfdn3y8XxGMPWgo1uESg2gr
S453AQ09ZaNIeY+fEX2jj2huL9jfeoNKs2MOfGAShFcGBf22dNL3AZ3tYMyVP/VQ
cLkFEzEBR/nlXNvTkzloKYeQZMi07n6TQCpEcDfghnQdH4tkDeqVLSj6W8Tv347I
FcEks7FBlIZrxNOBce4uIez++zE21Yir82OFWEtB6EHEpeJ61qFLYYsGmaUaRs+P
t6SnwthMyZ2+fIK4JkN8qLNsKr39hul710dAE69tsPhfEzJF46RtzQi6DWS56U1h
5URdAuxB55TEQZo5XyX76vsSpARnBqW1xO6p+4FnY7B8zVMYZ2f9SDn4SA5x25RB
yojFLQZCldLNBKP+uLc0Rh/qljbtPfRMkrSFxxBWrJaGPXLSo/L5kZGWT/diXTeZ
/w0sbmM+5GwX1Iveym1HXq81NGS9tuzfLfSh//Hhni2T+bKBxQ9PwH4mPCXfE1lR
0tb4c4sJvZ4lTQHnJE0UhkMGUWQ6Sk5uYpthQGdqe+hKYGPEYbN39fd35zVeNL9F
+WUOYp9/bojQyDYg//LVIha8GsXVbTnAkxiy5pHFIHdpk1wJY/UOnHfK6D/Mby5S
79tfKb7qLrSGD9K0O5I3r4pWZ/h/xWNtJZL2LPSAgj7UWr8QAKGSRUHmMzg5axuS
WXllzKRkaSimgH0AiFWaCOm9uhv6FDY8LYQhqF/FeIwRSUsN3Qeu9a0fM4fncx8D
MvnSSK3mmoASLW9mRM7esfYrN66txRG5skGrzR6cTB4H0CnRBnkiyiUIK8yvcosW
M9BhoKc6Y2M6VNFxOpeniYy4s7m1xH/AESG5itC7BC794tjH2168NkxAMqSkNl3g
2H/hpbk9RexWUru2EzbUhJUnbuVm/jX7NHHWvb4c+lOis8AUCCPJzaZ/TXTJ+Nry
YE0+vsPE3JDMfVr/0/UjTQHj7FLpRDpWxCToRuH4IeVKCn4+qLXP9sMyIgsmS4Wv
/8mJK+CLXb8uLHOnNttVo5fwl4rqKVt4ZQSitzN9UzV53PTxH1+nTarcRTCGgyWV
EW0e1gN3fvfcEWtEjkMH/3qacEynmwv2bYxo+4CQzKzPY2drBt5FZwBQak+KQ2jP
nYetCDQHAFB8ULoi5vZULu7ar9mAXBwyWZ3HNdYOXTUWegTjt+PDKiP8Ccmc0XgP
jbQfHHx7+oIdyjEQdoHv4PsZqM3hgnv8Xj7/JspQ9vTqXMxL/Y0ySwyFpD2Wt8k5
7+9e9FaprWeSd/jKDdVJtt8mDUt/IMWOXb2U/Bwbyyleaw7ZfEJCCLeadceMLDFm
NmqjIZdyTbVoOOWSm23SfxHcnFHhJ95SCPeHoqWEGp7XrSVaH5uBvuxS9asatWgZ
1sgaMq5+bMmFqjcJWCj9E8BloRH2loHGwd1Ql9ApRLtjEIhxcF7O3VjliRyTHCSc
k5D38mrlw7N7Vuvl9eW8M7/68mj99L6ddXiiIAQzrT3WYcQQFhWPXugd0hGUgYJV
r0q3Dnjx4dKA+0ww1/0BCU1GNx58lNb5JtuLjb1/yaXPdXtEGtQiVOEU5HjCE4SG
wnHxSzlZjsXsq69eQS5OpsDFbYgRZaDL9cMvx6iZ2de/+3umCsVE4jDifxYhDZnU
SFCta6lAiR8ZutYrDh5psyOk0TlKcZytxHObqhoIeVZNNuztfZNGdzklVmwpnjms
Mz/OvzsxnyVf937mian0iZj7W+ZAGHeml+ynDYGGht/tFsuyauUACQwgO+NLq3lr
Ip+1oCyyDN8BdFlF7xIq0JBvTr6u0M2dvGJonAf7NpuDjaTbYLkBKKClacW5gkne
BW4HqdfG4+AXK4A7+72ittygQCnxWRQrHYLheKiDrKP1vLAMmDe8OQgzg+jvQW5z
fBSf9hc/TbtPyET5e5jtFlxUKM6tpopPjkyIFh2iOYdZZYTyWt9CmdAQFCG8Iz28
1axW+83/8O2K2c1C6+ay25tcIgSfQ0G1GXRpAReqT20eEtoaLgzM0RV4JyPgsFQN
McdsgJlJL5i/SS16zks1EPjkclMluJSgX+wWDhXw6mSJ/vXdb4UDXf0Aeg2HtnVb
6IAVYB2xfovG4CySi+p+gELrTt0Sn+dmge21eC9ArlQQTRfrKDkVQMUJNQQgy97U
tuYbHAMPVpXK+aUPsLL1O8xtQd8Pb9h5TRpGzub8+0d8ffGMcWwr+vZ+O/8/K9tF
MH+42xgkLSDxrUPBMSQzy9GN9/EUZ2Lfp7BEHxWroEjgPGqbTOF32UoHK8R35Wbh
YqbH7RE5XNWGl2BfDgKAN0av0lnqTJG1l+6JaeaadujH6G0YqI3otZYIfb9nQ174
EiTx3ryVmduN8GWcmUGCyHOSN+2nwoFXKxp55l0VruyGip4O74L8qjBvXZVOmzA/
iJeRbfgizRreTDB/UJnJysFjebN7iDZy1z8qwv65KP9tNMMPpuVzUddPNjZJW5Qt
GSMlnXYyjCstH3AD5Av68FsaZGvguxOibXY5dHhfCx82zuiKFZsaB0NUQKLSxlgs
lqp15ImTBWLliF+FIc9QZ0RArMNZO1RiIT8Li7lgnEwL1WVwlVZxQRr7W4CGIwcB
Azj59Eyxm8xwmc7di/s+fd+lZ90aUnsyDk99vNXgh0ykjYZV+29YGvLZ3+AoDOG0
1Z2MxIdFI6b++3fQIdDu5tcS3qhKKkKtkHFOhYEKApSAJFHhtK7HPS8lmoQN5MqN
e9jTCbnW0cYDNx8MR3G0BVgPWO75f1yHZBgYrClh5LrPB2DqHf92nI98G4H5cSBH
7Q66nR3A5pexrgmfntJ1LbtQdDbK50nuOZ8Zdg4DL/gzgPPs0m1W5F/ZxTmYNU8P
wuarqsxbga8p/R7EALvpfTyRbsml/SNtyWY7cKSJJsbdznjnwfetsiin6o3eMJU9
8PTwp+5BTwescG+zX9HYwEeEsJh8v0CF9wABbktez8KX+9DiZHPr4opNOgl2Stzu
88k6O4zalMq/mluvEu9AWHtjZzXU5V1Qhx65AxhmilKukcVoFgjNZqMSluCJb571
CxZ7lmutaBHFRa6e3ZamBJtoOCN1hC86X94LYEZE4i+puMpz9KmoiITmEM/BM0cx
R6TKttejcaalg15jAYGZ72oMpO8clqR/TeJInikiXlF8ifHYBU2yrk4ev1Jmi/o7
DQpuIkP4LlvIKPYc6PgMw8kai4JDVIGGih1VM95TL87t2fnW7AZ2My29q6aWmirU
pgSQ0n6uX3PqFNinQOSJQIsbjmyQ5so8qBRp2gYKc+WnCrB6rC6/cqPSqXcZxT0j
2C/x4hIr+FsKSMty65vEY7c2I3TzB6jX1mU+FJ+Av/e+TKqfgOxde2RSf+17MtdJ
M7qtWWGN8u210tmdj3ajhpErCbsNA+RQbiBBpNSGcTKIFAR7ZfMOMCyjmELJAr9x
vRxYgR/0nF6C/bp6sgBMzQzCZBC9pY0L+Mf5B/HnLQb13N5d7rARdKqcv8wLnWwJ
dMMfr7jbK9AP3mHW6vBXreBuTtPpr0rklawS0m1yCkZdwqMvfVkL9FoomR9JNG6U
Sj0dadqgBHMD7Q5Uv3hZM64s+iM4EZuaXaU8EMPTuBNUNCxKP8Y5uybkk+t1yt68
SpZ7PvOp+9UkSue1O7sLqnMukRHuGHnS2Q182nkZMVZjVRgC3oB0zdKMZj6eKL4Q
5Qg7ijbvUtBvWyMA82MJnF6ZacyDZRoV55aRn1PptBaAH8ZdKNRgFuopbraHgWe7
/6KRPDLSxRd2+pYtr0LtAOUhv20A8yzCT58lt9P9Df2UK2U/POI091hB/aNB1DOg
Nr9lVYnwSjh8PKy1ZboLlXrjpIwNvlFytshvc2Fak+2ZA6C/8XBQkQErQ25vkGfw
n1YC+07S7AUSMTOaK13F/d9defSWXW8geBcDDrQfWJ7n5nmPRJoWeUp9acFjEBO7
RRZpQiRZBwVZQZWpU4V/HqrhT8ej22E5uls6lFRVNxZ9xfpL2oytNwjReWK4RmQx
67oPxcQGpgt9eUbfNcHvfAfL03SNOK93IrVfc8DR82hXWt1UfQOcvoZZxNn3fy2v
Z2VPwL/okyIkdAStvmRRS5Nd1NSVOb0rxfDUNbBrdaU63MvlTc1S0pR1fIDs1y/9
fBMZQP8Eb+lKThp34G9TveTPlHcLf74iumn2OV+EQrWrVghLqUotL4lmewftBrgT
vrf8a/SHKp5ByFqGf1dbO2fBIpSftHKDRFwRbHT6B2y/Kh7NxA1S6+OGYVMl6EOE
QIcHMpmLldBhVsgyHK98GTwdHa1K4qFjrAKS1WOfSugzrbXo2EMGnkCOz8PffRHu
x1GtZqvpHbQek98aApM32KNs5amleXCcSllk3v0q4M7nLD8DULpVwnAz7i0mM+VP
9bGYwpqtk3HTIo5VjKukXlglMpv7LCS0L+4LJudcMaL4kGYWCndpLVPvVkDjo6T7
/Zrpo5xxUH0lxF6rT0e3uBtQnvfwedqZ3hfLFxNQEJuJTtKFbjV0c9/BWj7bxTra
nwB+lpwCyidXGjEHHZhL1J4ZRNyg8OE1Pk1G1TSik0yafLjbCtxmrNa8amy79tpJ
Op9sjXkLteXWaGS/uk4LZbKA+Txny5+J0u+f4aUZ9XFMy4QaCS/GTKUMt2X8mpfb
M/iFKk+OkQ6kz9Wpsq+2MDXWGlyNsI0nDAyltCIXo1RS7+WTDfZXsOMCh9qZPX7U
1wgfzX+twrRyc/wDcZenMTdGC/HzuMnZOOGBp8knLAScfqB/5DWKszwCEwCeNwgv
UaSbbcjjX7JXQhRwvF8UgJR6irw8e2qtNq6Bm3aJIk172izyPlTXjv4C4qn4hkSe
mTjjDK+0dK/k2o8V99imo7i87HyYUrN85BySP/AmIk1mWpHEiSCVXCglMqwoN0ex
NSRoxBmr/eFzwjs+qYAFkY8OQhuYzvu3K5LlR52lgazDw2czCtVS6mlK2j9LRLkj
6Hyod1YI4+6uDhdEnEqQcbzNZp5+hsk53bc2NGWrX4+gg0soN3xI4CND5AlbbK0R
CcObntHYfZrA93JKM6ghRzqAziF5dCftV33PqCs2qYp8TltCEMNhZZ+vjybqxPzY
iWGtuCIaeuc/tc7RSwxIIrNei/QH8TXpevEVOE8JJYS/k6kiEx6tx3U5O/zzYyyb
whraAsiDvDciF+GfmaEuG8ChCDxBLZqt4R2k0BkV51bB9wc9KRnmjBi6e75WFiUa
M+FQ/6cDwuhWHa1rAr9jqPqH801jkO5oGp8it/Qbv5GvEsjSf8Ic7riw9iCUMCtd
38Ee7j+Y1tBIugbIOj5w/QiSxRl19RC2ChEk7NWdd8YvMT1G6w9TecQBogOEemGu
X++6x7lioJrDV2KPbq8wSKgAc+WLHw7dJ6GnMapzdJJg6OVpprmYX5YC6PVVyI5w
+uZAGcLpwCGP+IXUtX656DksuEg//RprSk7NXtYpBQ6rXZYM4Rt528/pn1fwl9GG
s5HUYKQ/h9am7Rh2hBKrgHNsx0hlBtAe31Bwzv3Xq1M0k/JQxhGrVCAHbf+uq+v+
sTt1TzmADGdgxWD4IFw43nycxa+GvWzZ+zR512SJZ6F9fqlQIrvw30KNsHpsVP0f
qjk7gMAZaE7WN1K46ooFw8I8A3XxjpGrTWF0FVfiM4zArswMnqQXP71JazZkrWtG
gGqyHwhWfyfQ8qczeX3PDvSs7kniDTNElqc5jiyvzHNu6hb7V8c30AnNW41lhERN
xIjqDmnQa2bim4cWZrSTLwke2Eij9ALzylRxXL6uERm1mUS+7RxxR9D8oaE5V+NZ
Rf03QCtqpm5mPfpzjF2nZ6lvcZh0EHmDdunQQ4G3sGRoUbcXpcs8LDxHPuVmjJPQ
gRb/fLRbcFPfl4OgtqSEB+E60lGKRvpHK1whz+uSu/YXagDbzu0xbLY3Tcbi+PHr
PrzHbJExSEwmRUciQ6ChNoL64HsBCUhPKKjQh7tjU00VflY+nQEftuQXVTn13RTH
jJjwlra+7oYqvv1Snil1abIj7B3aSOWJZz9Z0LNpCQrbSrJ4k2Heo1gZooHx6rEB
C/MViuxwJ2fiVPdpWNk/kQVPSQZrwSeHzwq28sHxgQm5/lDpV+N7YmGDrfiExCDT
DtASt3E2xS70WSRRXlPLV4YCURA4imYY0+Jh4hX3cw5sj63keR5BghEa/zb5qeih
p6FtgvZyQGgH8tC9fraLnLLA8t1RfIoBjQcEwx7397KqKw3yh5rncDsAoO5TpQ70
cC78WVBbFpC65TAk7znBhz1XBk/bZRc4XDP2/zR8y6s+lGREgMOgpiK7XQvJKhw9
eSDXxJd5VoZDIVhFMnoRpifX07fJztoieqNYQ4EoAByy0UM2rWNNZG5xvvQOXUyY
+FTk6DR/QR3He4AI3Uv4KqJ31pPTBxKnhG3pTv9vvp/yhz+L/u75O+gDJoRL5wpK
xNCb4L5gbjMi796MqPe8cS+xavWDLmtydJjEDXaq3KJ3a6mfMpik3pjjWDBrmWw0
zaPjAXlRiZPjPfmUDjM7ssd0Nl9kOE26hcG+r71NfYBnZyJ+UQ6o1MHoVTx1e9NI
6ZU6ajPxB3xG1YTK+G5cUoVAc5eOjs7dAPw5Kaz6/zgcOzXtKL+D274em/RVEyFM
5A/MVKxF8QV61vkbd1Q6HSdPIEtcoG68ZMlvq+5MFnEFFYmVPa4wmYx6yQBkn+g6
iIRNOACi2k+Subjfwan1nP2mqJxRQdI2UqJtFAHRupkTeFB3OIkSdWYinh+v3X3p
yT0JV4QPi4cD+T+3iQscDSCkLnt9OQJ2jOOn23jgL9zKjmLN3+IlycwPjX55FQVS
LK0DVGjWmnC3sjpTLw/Ah3dikrmStwuksPukCzyFcXN5OXCFa+vE11TEORY7dx6H
nPtyfSMEHUZwbPYoFgmAYXz0iVQ0y6JjyflWB6Ehr5GNHGWX6anrfw4m1mxqe0pM
k3MOVGoQyAVCc3k0wMxB2NxxBLrNCREDznFGtij+gsJXaQ14wJu/9SCgjryFtIK7
c+55EBZeOX7oqOyBltiWJ50l2MMjW8isPPxEnhQ2Jg/GDNU1+C9Gbtxx9o6Qusne
9ygoASHyE/LtUt90VsE0RbdjvsLCKhE0Fzr/2aHUgDe2z2Un9fD+VBbhk+u7ZIsl
LXDcE96142F2Oabi/ugEDTtRBFuwZdpf1C5MCyavqCuEuSY6Z0H7sVdErvQ7T0W/
WG4bQAzwMM+FWovz/GQkFZGwgG9tOfnI1v62hUFnajmk39SqSpHfngnHvQ0ZfP4h
wEah1VamtbHcWXbhwXj1Jrf//ccQULMK2poRqJKgalxvST9k0sIBt05iQH0TdIcQ
QKcftM9zmEx/VzI0rfTT40iGZTMhosd4IzwJezVhcgGKcoYvAZmHofdbL+K7Adzq
MNpLhUFL3FJpwgGe5JuF5PjY3RF3yEOfE7bagfVFnoA5Rz3RhfKC+rul9q6q+09D
N2cXblggJyaw/HaEqEi/VzYutU0wWwaAu0fdeHyzZU0mg/jk6d/z1SVRZeKWAIbr
X/CMzbzRP6Jvg+rOgufykj2zxeVjcOiHRA7PVizeynxg9bXQEtr3tHznw5tYOvBC
Lx9uGqKq7A6qDWijyxrdydOfiE2MXASIae7yw9pUdqUi1cnQtV+045gRiipMXvfJ
Bx45spLHO26Hjbdh+rgqnxTei/FdNC88tXfZTG31yD5bjc+FwoyK9Vc37BOGA5tr
cjqf4+SoOr8u/2WPpzxqErMHI14KekbsZJI2bgyczmY7llTTC4ezaMxmIDsimT3n
VJ2hP2SIdYmAG2meD6HrDYIe/EBfJfkjIxkKK2vbu80eLFj48x63Z8cFiFrN0l/g
N81/+GLuZXPoKAq5Vk+6GphIsRYM/Wi8LuX0p4Uevz+lt5DVfVoGJiAPSYWri04F
G7VR0zrtQHqWiDR0yuQJD6erzOLfTDY6YT1Wy4QQiWWq6Dai5Blvnu9NsjrsCoiz
8f/mlphTkZl9go5Aew/flLAOv2IfAtXyk8Am7FW0c/mUGnGzqkok/DERNBpWJHpr
lZ8+nCcuGKT9D9sYsmnpTX7iWgk8avnzp/FXhMlEjkWejYqY9SoD3M5CzFVhax7Z
sCRvDD2Vx9ccg0zfzSv2L0stKxxjPK9udjNTfGwjotSpTagmf3dfIHereSNX4Tji
hADeH0shhfxymBODSdVO2+usl2nLnMA/XjaB1jpxZZ+qYb8uTZJnCt1ON2NG2Ql3
CzDRdx+s6cIUdBRCLU+d7qoniJ+2L1JjMhsP/L+1kyeQoA6LuFRTQ/5IMWFPFZsv
EbRoWG0FNDCkMzUsWKly0QsY7o3cTXBIKlkyky6ilqN1URkrTHAog5WPRU51+uqS
R5u03wTw27AGOiZwMfePBIjDuTfin4G33rNGjMwT5gLsSvb/9DlJdxrFksKzWGPT
YV3ivZmqsS1cmWBQbM1bk9aG6Vx20kzBX/+4BPhY/mKInUCZLt23OpExp6ASN36p
wHoxeLyS1aP5pueAqcwgqt8x/SAfVQsbGaqHZaOkYnS2w8dpJeu2GJNwGhLvmaum
IfFdRwhjntxLfR73fysnRk854TnY3GCVFqMQ51JC/BU3ZkwaRA256ZkY7qQ6/W8h
YesUDLGdkGiq1TSePgsulQr/rlxsVeqjiBSR1sgvy0jE2YElIvIDQnqtaGocLiBp
t0WC+XF0rzDTVRpTVRHIkkH1RX/9LWrd3IxFgVoJjIvzEq8+kIGZmLNTRUDJR3Q9
c6zDu0srBDQpFnPeu6XOd1/eP/DeabjX/YHYxIcAjqMrEtbjkudCsK9EEyH8SHO1
WxTK5PUYkEShVRZmk+q7XiP98398CQv+T9GNjt+zUlmG4OgCK34xMDZqEhDIg39Z
L44kYWsy0BlfdK2WJw4+Xz7AicNr90ZViJNJFSA9eGtzUPNDAHg6cgSA3j2Uk+kf
kxfqzFuMhNwA8Y4vu8Rsd2bCiQB4WAA+xrEeOL4tJnlHL09kuZ5dRjudUSGRFU5M
GSkAstlip91iuSDyCF9pxN3+ws8PaUhI0glAc71zt4HGLPWNxzMDi8jfqbfWH4SR
gO3TOg59TePsrpZCt33Oyw2+BTaFygsdbEzDzoux2XOBU1xPPMcVtVaeAOjsMr5B
dStBStGAXCxj/VzAmzxap9M9eYPoecvunn+XQKF71HbISNN0ewhifEwpXMEBMOjD
4RHjiU8WngufrNn/iizX+brO7jAGkGkxOHiTXl00Xwb/16bFA8Fz59rfYUWTSBLI
+xwQVb+FaMSsSlrzJQ4Yr4Y8SYVZMjX52rpRaEC5E0kmjzJ/soihv68umbkxM04X
+hIOm7Zo7bYbZ7FpTjJ3BQsuu3J8Whztr+SrCAoahf2x5u4PyjYGQXHVuhuo6dwB
HXVwVHM6NP0bOcnBQF8SjFD4kAc2hUtURdSqswkqvAUTofL2LtIvWQYOdQh7k7qA
1LACM+KegLd9JHXlnBvbR9qgSyl6jLORrAJeI/T37u9q/rWsl66Dh5WTzN4zisSd
Vg9+eRzvANDiXrEgg0G1cKv/RI4dt/XScYZwWNtLzTnikQyTFvVN37rxId1fyzCu
b2TF822JPQy/NQ7cNTH+zJurClnymP4Oy8MBgIMmQdHnCE0cEGAtj5f6mMVxCfxp
uJanLhEP/phKaNHyWZnHoFQWCP24ZKYvDkfXs+CBm+uI2Vkhs7BZPXGxFzM7WXsd
4Diwm1XN4R8ibVTTUtJZJ9+KLjlWp/tOyoaQvjSvAf3nRGPOU5axjKdQH1+nf8X0
oTSm19/LXvC3PQOrgXpynRGjw1mx6bhxgOj+969wEuRuiV0GHlIr0lADJ3e7LOCb
8fTcVJ6jr9l595vL9qq+LUs04xj5TzlaR7bZ0AiOmB5xWGuECm18HAh2Dn74DYPs
UWAgbje0FQOCdSQr/gG7D9lH+pJ2nxC5Uu9RgNzszzNEs8ojEHMDVkYI0jKTuGcq
uLtTFFB2zhjSWZBHEfrARoKY/rnUuDc1MpwdAmzU//My64PMCCyusM5ocCavX2Dt
sIdqlk6PQ2O8dj9ofLDbkhfiq7dgfVyLMt4CrK0CcYUgDzV238oQt+X7LEdsc2ZO
7OpDATjy46O+r3eJEkuMhr+bhJgkLzhDenxLIgLe7IrkaaRY89B9z3OqCyP6mfcR
C7iBrlkRWqsJt9pBNGZOtRz74UZXzaVpSLrpgEhEktKT6NmZ2N6j0kI0D1pFLmqS
bwBV/0vNfdo+Qf5r3r+5UPL4exQCOxbfUQl5pzJVM0YXnJtYZu4IVqvtJSgL59SZ
VANQtKK5rHkOmxWgq3yJEx0oy2AwaDO6BZZB6TwNkIHbWSidBaZmmg3lWdKY0Wn3
6nafzqOsAoN6FCmuwmLx7Frm3p9i/UJb+MyDOcGwpik65+AkVafV9luOUaWb2NTC
TisMU0YK2418wFD6+LAtud7zfT3i4u0AVmVChEUFyujqwyVOn/J3qzO13fClgqr3
e3CeYK3C3ZccngmYpBfJ6ju1KZ6HASCOH3/eSgW0+7KU9X/BdJZjRZyybAJFu0Tu
UaLiRhGDw3RiYiLu3xIWJS2iai3RVPKSylQpmN3exG15nn4BpOAQNUDSN3vSWqAa
pDo2+cMFOwfr2KoEeaKL0ydymM3JSddaJiTXL+YmFIVL8BJbt//j3BI/3xlq924M
WgTJMc/m+qdgx8qstfzZWsNDa83uYcCUv6B9TfKpZj9u98p2yq6DssWcpeunbqTb
RpD6wY6WAmwn2RqUSygj967aQ5+OpK3rJ5JPSmqPrH6Dw7UKbRsJ+R3gcliYUmXd
E6hnkujZ/ebZ+KfFQwMIys9+vfdQqS0WEgqMGqVBSdc4ExzqCadJuA934nEg7IU+
ATdY6VAavz7OMt7w6Q4mjKK0Aw1WP7kBFamxziu0IuaNf2fYu8AS9QjIX/uD2cLZ
OJQcFf7Bk0xDAYsOFuK9Hp0Gc0yQgpnUioNSpEyvSKonLQ6NdGL6/xeGeZkmr0/7
/ullajElJjPggzue/Qu8ZCNfn56U3jatlVZX/tFfBF7WCCNzDX+Mfk+zF3+Jmnfn
Vv0O223xRzr6vQEm7QceqxpRp6FWFX+ufC6EM12dxAyiaFpRJ2Rl64MvPR+Ex03u
6YFGTI023DHDGMyqGTNiyrgQkP+1dFot14hfxDKoRCJC12U3uLS7F/m5/i40lHoW
fTq5TfiaXxYRllo4PVem1OfkW+3WPYHTcD/6Xy0hJINgOtAaeL5cZkcW9K3fClQe
1wOXopKLZIS02Mkj3QMi9v5VvVfJKIP9GtLJMmRGlVWQG1xq3HYizrCOeO2z8F9E
hxOK+eZDecDOGGpW5hRPx+qmxXu6BOgofWRVEaWsRTeiQSI6hoieEVWQ9eo8VFTd
ThEY0aHl22F5Z7tnY0axu1At7dFMX/bHD4l0q9pg7jHKWQcyKJrd7bTC8dbHXpTq
0CSrQMNLsnmlna9vkK/lNs0iycJwqq6k/rwEXEyUE6jbjn0UuM90KYSBYC18XEm/
7dP9ReSP+NbuG80SXhdNmL2QEFKneyQmOAD6kb6MePtMhK8gteoaW1djXaKIUPTI
nzans1IGUsrecCAht3UAKKAzHbnCNT1Xl4bpsdGA6o4fCgMxafZ0bSmfJ3OmVba5
cpqhVmrFBp3g1NpYHd335tvmeRqIgIlw4aWqzt6a/Zf/3rd79Ot19ClT/P/DPHBL
Wd416vuL/DtYTZvz78pDG8TBoBjYONhbyGEcKahyoW35a70sXze7LMk+zAwD6Zit
LxwSV2cLbLi3mTk3XpXsBSEciHUoYcg34jgMiX/VVHgB0k7eAjs0yfh7oiFmgTi+
ZEZQNLebIvJTpEDgFB+j9qyjJGLX0af4sTsbouej2Zc6djDCJzsslRTD0uAUCVBN
iBVa2YRP9bmsiRpsBL3IhOe9NL98sTV+IkG36YNMYw7B73anaw4C2qum6dZzCet5
p9hBQ/H/boRtsW+Bk+DnI7Fpr583R0nBltkU5Lr1tmLHh1IcdL48EQvkizN8v4tl
aa4noROIHtmFE2UvHY0quUeyZXV/BsblUryCZSmFQoE/H2DUr0TPNe/gP8xcpxnt
xF3kBl6RxsD+BanxrEb3may1EmxXLMoE0ctWTgt6mA6+oIjSF1YcLQ3vqbSybJna
R8JkhnuULQzf1fF2hyQUNySC+OT0E8q5zXIPZgb7GX4WupfGGLsvw987tMW0FImg
UzPNesrMRdG4eZqRolvPyWLjNNuWo6zXqilc+eLQ0bwywKajXw+bt+FrL1l20/tn
Jn+CEhvfvG1hHKOvR0afxUOuDEKL0YxEyLfZ9F0MmE1b0Uyq2odZfHWkVHPux4HX
LBWQM3s8jQESOeamaMhqvb5z2Ak5wUI8TrnUL4Kee1MjHHAFoX4pv4PdmLcDMWcp
EK/0bo/i0q3T15gKvDiW6YB059L9EYTNpZoPIpuuMCKeFNaqkrOetJYh6MXWapnB
E9x9YgrY+3BPpJPf8y3G3vKerb+jsWUpNK7TWhmOp6wjAmZCsqyGvxxW0UDpRIjj
+vxc4xfLnaCrmkto1w5GVfBELa0gKB9kP7vINh5gzuJXgSY8KEpDvwCUdyRIbfv5
6181NkEWNCqLFl0CTpTdo79R+69epKD8kJbElcbTKDUm6CW7BpUNC+0/FUWKemC8
ULmfX2iqWCzm4RSO7KeMQafyG2HLNLiu8vOh204TMqf7OYSSJ/Ght7h85Io/FMoP
ruYG9zyLSTlwgbQrnhSDnNcQc9C+7PYpjreBaV9qk9LZaoJlZKP16gjuNKZpTdGJ
0nAVXF08W/3NaFN2deQoP1Mijbr0X4E5FCHpVeOKCUEyhFLwq5IlqHPgnbV1An4G
AgO32clzj16CR/9oKRSIvL4nug4TtxmBG+PX297qRiMmT1VIPXX3SceFG/ff95Ml
3PYbfxq3m728QSGXCkHp3sE0A0NveGjW2pDC3de9H9PvxTf0fSUAAdxeFj7Llr0v
/rXqLy42Mwl6m2ulJykzLECuTAb4bI2TgK3EAYTnmUR47STEG2XgR+P98D7edrh5
sRxi0TyYjKtPfwKaJhdrz5JkxFo4Sdb0IQ29n2PAxWI8OZDh0NpkuX9zZhTG+zFo
PCa+xPjppBndz4DbrAYHLQlnR85g7re13vffL08HUzqbxH9+dYgGxOfxz6hTXcGc
i5jSJrW4XXZf/Rz2pDJ7g42yjZppq9MdHGApqjb5AmGFvT24ODWMAlVhw2vislKk
p/UC9znniq4jUg2zttIA4UD0TAO5Tf1O7L8nCm/OihoralubfqHXlVc7kob0Hobx
8kbebw7rp3/b9MQDUMVJgD4adq7mfPX/8SbRqBB/eMkQPJbWmFhXkEAYDlKGh483
XxoXzdO3baCHGLQoBuspnrgnyNu579wGhdaoVT6AJRdcY0fYsNEj9eZMQLZcHbih
KG4dmQtTfqZuGVzFRSO/Ip79IEtWd8rNUW4C/oMkzEDk+Y47xpe1ShGtbVs6t9nN
owV26FDlUnKOV3u7V+tZXh75lYkwLRzbj91hAFt0qzj+MzVqr4+regTGpMcE5gj2
12kes2V+qJ/qXRH2+RdsKkPALfIIFr7vJzZAQGNP4rV8ZJ5dtQmq/RCZWKO0wpGJ
Cq+T8AUdBhB5csCYSOytuOwkb2I83WJIm6DezuBFowE0PttgygvPIL2EBUUoeyEA
tKR5XiW6YTyOBm+xJ3kmw3YK9HAmusXsvURzR+2r1UmddFtB6k6A73jZrtSs0qsk
Gu+UTHj2n2hrthy3Ef9fn7fLJHlnX94QnJuAmYNYJnt6/QBDYy7lGkgOgckCcsCy
uxPm/U8WsRjf9lnWcFVQDwBqVtYll/MNP9yfZ/vOYu7wriAfbK9ECMR8Q7Q7uWnl
gs3KjYI44451MTHY6rEYBTpLI+cL8RTJYktdUaWvuSLKyekE8vUbXEDmXarQc11N
T0xu7NYdSXsHwNi6JhZaASHI79pN1+hAHq8Xt/r9Ofk+KnD44trP+Gyx7WYDKFKc
UQR7359nVX23smOXslGe3oAs6p+XQssFFWiUtthdrAEZ05ml1oJwQ2KcKxHnmu43
ejAekdfG9pLsaYweX+u5NRZWSxzBsDOTve5LN+F5jzX/mJKfFonEuU878Y4Lgh7R
DkeCqX7ueiUjmYZrD82Zq9oxW+khLho6FmLnzc9N42W5tWDgbYjB57ZzJSZ+jbYR
65g9VWDx3gA2ua8gq6pL3xlKyhSXZV39P5GkklO3FR6Bc6aKpfca/WhYB9QwEjA5
C1wbTxaGz62WWVUJhGreA8wXQ7uasq9CfMYc2zE8kB7r2IR+yCF/oFYXyaa9I8Ud
ylhvkpsi4MUjLpVap7+9wRYKFclho1wqz9id5c89ruxW1mTaRoVcYHtjy3JdH6ou
L8e3twkXB28HDiMDmQczLFuaTlAmvjWWGLM4c97XzJbVAjiR0uSXTc2IylBJt07v
dTeLYZcMkMKf0+fFdiLzZWLP6pYuUwJA7c/yy43EI880wegOk4JyogLgxmGtxG2c
QwCUkgdHjLyOsn3tZTJRpfMuBZHIwEuJq0t/0INEQ00EuCe89kAv3Y3gSxtKMEFv
E+aiWy9F6su7jb9UtTh1O1EhCI83Tq0Z50vHofUMHVwcfvvhtV1XbNf/MmBEmpc/
od/9X2VVyuox4a5F/eGkkPM4npWH2NOgjqobRKmgpHaLpermOrjs6buvQ5aQoCAu
HSiBEaORKku/ZlSGCa+I93vTGUVhX1A942Qh5Ac7oS+0BnBngiJS2ORe8bSLAbIO
N7qWt6f6m+KXki/VVTCBxLwkbZCf5Kn9DKo3073UHBtMCkBUYuiloifIS7PrGAyM
wAK1LgqQLPunmy2kVe8ZXryjugBYorMW2VmY9Ry6VTF5+NELn4XjQmWC8Dl9c2Kb
cY77kEZ7yC/TEzc+IMpVeozNKGchMKFMj5hyYexk3Fbh5INCiGjUWCvzB0v8m4uu
7anSja2+mPS1gEZT9+qdmHNbcI7SOr2d3yFcHt0Up09S1k5Rf42GCm2ruQOZl/kL
DkaJdKzrl+Pp3fmQ9xiYiK4vT4BH0xVDoWHh5LdIOt5FTeo+u3kMoK+2gfbORm6l
4oH+Wf1ExBf6yhCt1XZie5QmEZnbxLhCnvj4MxJJ+uga/4AdA39li3NGc2sKwKLP
s0ig9HaKAUOX2PGw+A9NyfP1YvLFCsctGRLJWltDoIdlRP+H/rpl0UFK28CPLhzA
F6eE/9MZGQaeqXSqoF+nO8JIHcRfxO7yk4L69EJ8H5W11Gb/mgY9jnp00q/ZW/HF
IDeUIxMaYPHQrQA4Wz9pVYld1aDc3S+QM4Ic29gGqi75FPY5lKSwIlq6dLYTL4VK
11X/agOBN37mb7qBBq6jXet90QtFeJr1yzVaX3G8eco6RxVaZOCC46pZzGu91x0j
+AXntLMl6jiyNrfHZZmXKigVSVknpCHZKvu1jFFp6zL54wDj1bb1kCu7Rune0Bj9
4t7Ii0sfzR/HKtntgNfbIVb49hkuOdpgYRsAYD5ul2kT/SKdkGYWVtiQqCz8582P
CS6k+twANzM1vCMFT/gQoz4JCa+uvXWPypOoA3aL5GXezwrCkrzmFfMZlsTDBzWl
HHavQg2gC7meMqRiMF6s1Flw8yD56szZ6jEt5QAimEmTq2jFKxE/F3El8MOP/iei
BulqrHmHOPES2u69fAgCpzyFjOtMGMGx204ypjguH8PyXQjGfIsHTSlOdd+ULKpe
WUGB3AvfiRiXio0pX1Qv+yejCoTpYuDzWQiYf9nECXBrkGkBmp2jysdI96JC3L9e
ziYslN6XzngLpdrX0bj7oXJ//k07UAVAw/GWJhaP7z6KyoWQeEyhF8Ov+RxjG37F
OqUPfqjrEq2n3ALG0x37vt/uTnTmlbnDB7RnpAHjGZkGGL3FrrArv5ELg1kPjflJ
Tsr12XXTjb9ZD2c9VEKOt6u7ROlzj58NPWcbPfW1+JK4zIJvdXtdnADUI1ljKtAq
Ek3zfJl9K2882KGqUhELgfUQBbCQLuzhU+sNK9LoZuuaxeWz+Yo0LIrUzi7NpUiu
kNpRf1Otnnsxvwj8n1HmP1RAV1pbijRiLej1QK84CcHkpEo13orJqTOKfwqkNY75
pc3+pJLDEs6GgflFpHghYB9Ntxy6fTZAr1DchH+TjeNCZ5aa0/HueQHEBEsireJi
DHj0P25MvmWmOkECOZ0tLgvWe3vSfLBcopXFZhC2sgppxRfAsM2JJELyJ7//zcRS
pf/RVjl9vwq0/QfVaH68svHHYrwBMmmPs0Y1QNwJ30zlg6SVpwv+CumrRDmRyxye
/9Hze8yROSi1dotyKmKQ6Zu0gCxndcRXQvwN6yKQNUJIyt1+bdNW0Vu05DAkOle7
FLnOU6QgbaSITrDTo0KSTmpwJml/zXniEsba4JXN0Wt0Iy9Lrb7szfMbXCkj0RhC
vLJGaAm+4EckIEraeWW5MLTlv6hhXOPWpSFAqIDxHTyNaM0PcNDlf6Sv8erUFyhf
ux6RxdDTuqZPc9X0qc7U3YTP3D337h7PcfnFVGe3UID7TMMg2HM42h9mI83KXnMl
ukb9QSfJgnQyGIh5mA63fERIwVnaJq4yTxWuBPbfGfrH0bHj5xcTWyC/4NyrNiQ0
9pPCJPXLfaw8IP0AIJvtIXMqOm8P75VXvtJ0pfZHnGy11+LElekYy8N0HAhtP6+x
i7SQw/xZFl9Ceuod92O1ai5onE98iifwFeOZwqcufdGwE0IodbHVFKVfjkymcBuo
CJF66oUO+8uk6tdi6cO0gpVehECrUfCcBcnytZNvrsXpuZpKTNP19WB0Q/qwQJkO
Lf0UgB2eSz/tSSI6q6d+ClfGUPc5Y2RAe/AImD8XyvRmSxaQY2+XAEfyRE4wf+iX
GJ7CBz4ie2ZKtPqgRjoEAk9Aa1wpxIBhiEOIczCpmquGj+9c+bN+lMA2seHn6KrV
qIjsbI04h1tLv6tALWflCWdsNq4ssB/tQbzAJWmuJiBTfZ4H1BzGkqm9gYYnipQD
gwNXeKLNLj4uQUHFHIJbFn680Q82YA/X0F7eWsMKYzYETYiOrGffjBE18XClmNqA
YM7+954axre06nRDHWOjSIo0kYomE3lXW4DZCIFv6mQYawJIrkQgE/pv6MwM2V4C
41socQ/x5//JxfwKxE9bOU3sdFuLaQzIcmLBROtxW2qkIeP2kZbW/tLGria8aRUn
NKKCXbDGkzee3U8OT557lWr94Iy2xEEJRQSJbMthdzSCfKLxqbuJ2vU1Eds2aNc4
SjG6gsWDXpbia6nJYRAunRJODLmuauw3k1Bv50f8pbl77ZeG5pgl1XC46iasqj/0
UFncZBH8mBhfCNmd68m5x50+YUqHSgCTTsXRHkH2Pxd//HCiOunPKycuTHRkDT+/
xZNfKCkBcBshvmms0A4oUit2MPuKEYtSSCryNzE+xRi4pikur74E6C46og2dfYvx
RFnGyjV85aoa1uSC3JJBPtGus2POWnqFcIHRk/dHC3DmrM0l7H6EfWtsN+zQXGXU
0r/PAsjraMEyrtCTo1quLiCFawgC3gibkmLvlKwc8Qx1PHccIdoaK9xCwPRvH3sp
yUNXu5Ls15Qs46KSZmXxo3hlmoAaW+UWsSVHIeA6OIs5SWvTMux7UYiiOJ/bIKw9
4f+mrXxXFmUu/EAz6huKZ4sw8H7V+cQ2JLtZ+CrCKO7Wi5EyVkM/sQlCwMvFoB7z
g1ctqgPC/6I28UizCbXMvDJlTIaHHeh+2ai8lfmvdFT+HzSRaxhFv6GVpY8UU9VP
V4jr060Sr2v5X7nJzDZKHNvAN5gUF8As3FfT7rTPl2V31iAOWKLQrwPyBUBgLx19
SaqvajhTgjLJpm4ZFny6SHzvjK3mjFheNXKwVj3ulk6hWPviK9OMSViSdAZWi5th
ghKjiVIMRhv2x/jR8Utc6rge0HJ1IrhIz2DcFbASXSu8kGLpCbziOrMyW1Z6gTlf
xzoUKl2+o3rGbGQAMO4LTdvz+U/XWM1tQgRXRhrs5eE0HspUOZimKFruydRdHmty
+ZSvVDlXqTNm2pQs2p6aSQ2mYwS2IukEPrFO/cyOnlTyPWqGZmSEgKjkA0cs0wyY
midxSRr92FpAWzSJlISE++aEAlnaaERmmP0UhlkqDsQUxxMYFgCd0wtuubimeXyn
DjTKQJ5KbKjPUaVuRjv1hgPct4owzh4FJz3lPKYH4c6HPhfKNZD22Vc/A9jqWpWw
rSRHrkTfsgZkVaXxbT0P/cTaZKrpVeistry6w+jWP9x9ntxaQfqqR7gw+JtM9VFB
1lJL9nGk8YO3nxncBta1ndH8eRKDz8HIqBV9AlSnDBcmlmBWMHyN1/YDz86kaxKn
P1B5S9JpJQBk1ezR65x5FD88Dsv8hOtOBG8sUyf24ALdWCCOkS0Xo3Ttm8/dXruh
G6xgW5q6zwYMpTHLMo/T4mzsF1BE0+31VjpCAMsyImy4Nd1VyDELmvA0eZY13Lkp
RZoUu7+bNHvCg7+/P58Yuz2NqE3fUqk+KNfPtrUz4FNqMk5g3zYTZIfelvnnPVyq
zrpcEHeRbCtvq3a1Gd4ZdWU9WDLH6ZrJGVrDAPB4oGopGS/Svhc927sPXaO4/XiE
73Z25b0li7XRrMGuxb0Vl/Dypj4RTNX6hgOdy/3RKAoeSOEEH+bFLgLcNGDTGvc8
388Rp8Y3W4chSgsAuGuilbDEoYQxSOA4H9gXE8aOj8uL94LLA5UPOFwUE748/0jg
0ufBlTdeJDC9LUCRw/teSCUrhnWtclSAmniM1Tcgog+di9si8At4VeUlHEhfUR7s
YP6RWhJY0nWNWVbVNy4xJ+OADlY0Ul5Fmp+3rN5r8K7ghRsf2vQ97QqnCR/2OBE1
oo4rRhTfF7gwAD6OGC+LZO4Wk18/oewIdzJhD/UJe8umXPdPJM5SaYLVFOOPRTfD
x0WKIRqOZryz8+/1ZXKQrDVP3nylG8h3QtW3+NoE5CXCib3ptCtHnklZkHoAydqo
eg20xjQ4u8F+1pr8fV63y4DxoFyV6r63mfesrvXkvDzOjU4ULPX+tukiMeZEx8C+
R0LHyfZ6wGCSi5PdfhDF/zj+TcOcFW4kAekntvfktzY4TOQh2S21IP8WfEldreso
NRsAnWHgiAV0NBsjASBFx6qkDfYeT2uRR9EMtstm8fdbEW+FfDY4pUiliuIvbo1j
mJYD64d9NrDW+r6CNVsFS8vmGxMKkC7K14V7E70Q3wSr8Rx03SoOQjfWmt84tw1k
qR6Mun4/DUmLpQBQMY9S6vZS1ELqsroMyZo5H2beh0jDJxLgTT/aOQzDvPQ4l2YA
Njc5BkcygXozUrGyEij8dBBOize5sEvOq8n5GkAY2nwRO1EFFe4JBhIsvhaZNn6f
jasIAdtun6TW8VXMBpcmijotvPGX0K6t0BZJd8izXKccAO7tOrbD2NuOpWHVcuNO
mp3bffuh4O99z0UG2gL3ZYruRx7Am2kLyTiZshcevaDKEJDC/EQFYqw9ENTV2QBj
nptc1mrqivRhlWIn4X/aolsi5Kvrjj+AMpuph2xQCUfjVjqhAaS3tFXf52Xpo2eR
lJPkIUOTYKVyPATDkjeNZYjY3NWH08rBJAM5YuijjWPLv8Wkh13641IWGXXeuMLa
wU7LpCu5GkWavXim33NCG03X6NpBh1LX9wPPPEKsqGQbSVccAuZMgs2kaJYGcqgW
xg/Xww52CI+rAl010f1elCH/DcU2mez776EQDa7g0N9qytfZpurwTHAzoL+fIojP
TOn56CFOT0gkE4DREtaEsdiysldPJhdYCF/zuozGfHh240K2XL68kks8+/n8Ox0g
en8B008Z6pQQ/qscD2u+VbtS7rPASmaZ/rI0ypTtBUjJ03mvhMTS4ltTO7wjWXgk
jfwAdKfvcVY15Kj9Woj/60mbU8e+vpG8xoNVa4GevlGiV1zEefM+0sDG2MA2zmPj
npAifPuOrY99Yz1TAmnWN72rH9pOWYHJm9qSUGrsHYzIq8J48V4uSO1XR501ASe7
5M4ejUvWdB4S7M+vx1rdysdyWD+twBcxHdJvJdQmjVxR+ZsSGpWWP4S6tyNO9a8S
AS190Ty9wxKMwxSbfldQXutzDSnJEFacAIUq9h9WQqJSBeLKWjR/guS/j3Z9Nl7a
Z28LnTPiWiTX73IfwZtRdj9F0m52f4Dqgr0jz8MG4zu6xkCIQKI8gmlfHKrUv99Z
CnOGffRZCcyPG+//rKwxyAALlJKc9HHtf9Jfpk8MqByPVdsP/C7m7fWhJUcCm07D
RkeqFahpHEggyzvVdHzqTlp4jlE4M230ozwQsw5qakB8KiIYOY8eHWHSkIrZZMIG
n3IHWFqhZJafioyjrMpBrCKH/btRb43Mjrv3lAb8WbznV3w8jBysRq3/lF6calUT
GeqhCex/1OEtkWAOV6VUOWh/g75XU3iaLSUQVCAXPt+BZjHhMCcij073zeaBRgK3
0QwZ/c1Xl36vnXyzCKR2Vov+Jj5aaqB8lGCjI+yUez7HR4fiKCd9eh6cYsE9vy/0
yZORA8TCfJOvVC7miDJG72MMCSyKeBBd8d67bnONxPgvVX8Jpk+iRX7w6nxDRWYt
BHGkPUZ1hEnC5d+HWIAvCFNcCcANtBmnjt/y0utGQfTrIgNVR26cTFk29/PMcBfN
NSGm5XaxGbTg9+xITMvBJ5DIT4BmccZUpBXPfayb0TLPnqHABYFqzM3WD6DCAq4j
FYLIl/D9SBsd7qf1fEJYQSjk8xzoE3aoi+JOxS35vHBtWSoTkTHZUfQzIN2F9W2R
aO/U9JfOSfU+WYGxZOs/ve5j6LQUqcokDzP0OAqYxLaBd/AvlZ2oxK/ev+5mllzo
0N2GSM9zYMgfCbF5URiVdWpj8BINxr1WUgNLHTP1ZbRAiG+VYFew2cUFbl+Gh6GB
nrrIPJ/OPVbkiAOooTHWVhaib5o8y0j5I1NYWWMpp/8fnrHfRqSjuh+q0Uq7Edlj
Sp4ttT+vPdXU07BX+1MMY5UOhJcMPKYEzEFttK1IYT2eCysjFDbv6NF5PLrR0AKv
dibUdldFkH1ihXgygzs/Z29nEwD3INtXOWqbdGwERRKcWeJM4XXVIE9HqsRdhPxn
POksvhyMziCe9dkBJt9MMHMZyXJIvERtCvKtS0xTww60muLHQz19Z1eZlerU2sdS
vJccSwZKyG2fjA5yzWw74ZRrPTboHFKzuYpH2zE3tpiGWCSgZHOj/EKt/4S7hHL1
DRaDdkhJA7XvDVltKBmm0Y5dZGyXC87g1Q3PCKX12zufdsGhmWMDhh3cnmstUgmN
Swh8n2GFVMQf8dimgI8KiZXtFOOghBtSmcts8qM4TKi/V5rruq8axrhXeAiB5J+a
myyNcGxiUvvShMy7wZIYmF7d84cgpAVPnlG5npMa/F05KHmKjzsOvHGZVlvJRaH9
adj+G+E0mkkHzXCgzSsoDleE7lnwAYjgyldCyNbDz8te/rQsqNPEcqBvryhJRYGq
ev3n6YoHyYiUhYXv6DcvBgMRQUNkHBOl3MDEzn2kz8dVl/55jjL1IrawaDIhMuNU
Q0L8di0Gmm2nRdeTqIJQ0oh0WKZ1bsbgLGLChbAud39Qr/U3nxLQaqFaXj81LscA
GQduWjputmpJN6R4MsFWc4JqJHUkhL9RszKaxGQAtBljTpvyo9fOny3UAfxd6j1I
X7/L9L9DLfKiVMBMe2JdqoXSMYwEXFSJMsg7+ssql6VkNOxau/7YiiZlkqSeWJC5
jdGdnINRlVjtzlf5zaPXwMZNqn75ZcVyyOzp95N3Fq0aLyWObXZSlbOGx4QCy5BM
6jbZr2OaXy910fGL9CFVdC8eeUDNHD9LY+HPYrkXLx0sd6MMueT7uo1wt+xBu9HI
xWcDXTzKvAJF+qEUlh/cHHZhWdQR0jCjXVsstfzYIhC2O3N5MDFFoUyVwYSlGPHg
E5CaVC/ulH+tw5vaDW1iUlASiN3Qy/+qMNkpBtY2HmOLysYpmpTe/6XjZKiUFYG/
GjGC1qpb+9/WSd58YrDoKXlKQVlTR+E4lDGggBuyeeREHE1s5kGPEEviCJ8b9U9E
++QIsHttILIudJjyBR1GNyi0DAxwgSjNdIjJ27/MXVOGbocGLHnhaWDUQJIUxoBf
43EwNrK8CKr+i37xjkRUS0HPCkVCowfcWSMQGyAc1R5+A97zFLHSpTRaBZ262mUU
CzCzenHiQuluAye5sx0Vrvok9XcryMaRX0FlRTZujnMumeoFS+lnCBTblrO1aP8U
hCnNsZR/oP4VexQ0EoIWd5HnBRBrvSqnpJ0fNp6n7LfV1xL6ku3qM67OGuiKnoVi
grAzLBjia/mcIUKk0eS33Tx/2PAO8X5VgcscYrxqxD036U3S8G7Dbo7U0jk7Mmi1
S7SGCrCxKAB7Ro9NGcAUUsmzxD5UpnaH7Vu0rS1rjKcPfiiW8ZbbAXG6oGUETRGf
3lhOS4aIT1B6pJ9Hkix1aZUOouGxLzGFJks19rFtqRabfblydo28nM09eRKTt9BS
OaMD6fbPgKH4pw+0Xb8Zusm2NOP4uJragkWTXv71mH2h/MPgAJLQkV8TE9CQ26CP
jiJiZbSralgpop+Jsmfqq5SfvKKNqx/5HQgA4Kq0c8BxUpug6kZyDiOdQgz69fqX
4fRU+YIlv0T6tnEcW/DGufwJEZSbHf1v6N/X55MXG3NYsWWWdHUl7n6vu+r9SWYr
ImM8w1WnsOLoDVSZVtDcyemMee5fumt3d1UCHgMK0njsXn7BKe165kxiOMY1edOz
yGbJA7wdTnUvejCEmyC84IFktO1keHeQvTywuGxW+Z0vNf6brzIcsFIGkVIH5WpI
z0hwMfA6Cq0XlENDM42esddYf1saJULRxFRtePzbTlFNqFMhJiy1Stc4MgsBLWom
73IRHh58wLfxhf7OjpgS3+mnLo/nr+/XcpgnLgAaYmgl3s13t+AHCPSHWVJITO/B
EZ4oVJsAes66eU7opFF6Zn2j6bmvXYxLRlpCbeMGgvrS3D2kYBzZnaUNaBHXikHN
Zy6aglfRgCr61ow7jrfyQv4fxvRmf2j9j5OpLfYeX0N5OW95NzyIIOexEmwq/nHN
N+ZgcgCN8SwX+ZpN6O6nRbbz2uqUMG1OljNV/jGfRXdjEPiiar1WnB+V4WwLzmzj
tKbvMhB1+dEI7hk43ZI8BE6sv/5sTs21LdPmDwOIQgA6fBAISbIaiFY/WsXGpQU0
NpGq87a+jVKHpxmnpE2MfTIO30745wmapY2fj70JWwfYiD7Fuz/5edHHcnFdz0xd
J268Yy67y30bToFAUAxjINU0cV/In7NziRlWc8f9vMhdmilZOzX8BKk9VXMl2DF7
Q7TUHIQrVRocCAuDTxueQ7LAMaXaFw2qAdoU7/EPAKDQtp943e/jlelnr9Ix4eDQ
Cuor46LSAvJzVXpgh2RQ6xiD/NhVTg8LH6s0PIl8aMfiqvc2F1WBH+Q373lq9TU1
M8/by61CVP1zn45BGP7zE/hX5IbLE8m28LTHjygeZYebGZp4+7oD2O45vB0PhdMT
3+EpE91Ce75Jl5PSQywU7Pq/Adw8lV3LiMDRPwS/6nv/rekuSBIbnsLlBU+yv/Zi
tLLr5XaabUVMuq2R5TnwE1r6P07sieXbncoASnStfn516xuG5/sJN0sB65kZ0QZK
a3u5nQ+rNagA5GPnWtFZWCrq1bRCTnZt7nyFaeJeYFWLgzWFb3AJOhyyumV02b33
o8XoDmEKyymWWvpXq1MaxFB+u6Qf9GZ5JgGy/O49VnIWmVPL0MlQzHZg5NEJGS/P
IWE4N/OR+ApljHwqJLxpnLopdkMFH27RQRl9Db1TEFkbTkGIKzk13e/HaXTJJpjk
Gzo3SXsZG0c4zq4l55h9mAI8fmoki111LurZ7tYyGITkkbKZuFSMKzcZO6x9aHV3
/9kyC2Z4TmH5PFnKREKF/NwCE2tiMS3SNfoCD4VikTgFrqeI5xUXFNuuNvNY6286
wALh5ljQ6upA5PboURCPzx3cSHZ4xE3vYPzcR8/ouz0ZZ3cL8BZqFAGGfg5mfjXO
AJNamd4wbxn5+Cr4SuLV1GvDj0Fc6t8pBUkQK/2eIpU+87aC9XVN6TwHift/WgUY
TEtkIWC9FdPX8WHEf/3+qUUNAyaICXktJmVvmY0jA8Z4QO43POKpLrWI3dUjlflp
zLx5YImkdVNk5n8ArZdW49JX/4iCEgLHTPfoYQjM5RHMDAkvM7olUtqZIxBxn6NA
z7JoPtE9IXvSnBR427/2QhfHU8gVq2dySEmp9T/MlYrxZRJcaDJ+rRFigrQp1cgr
ppQfG+POWCMKNRzafFQQsgpReT11x213F225FFTk2qFcawihSUdQSKrMBSjwD/3j
C1N9yOFnykitg+21BjXjwFyN16N4+CGR5rdCLdZnIXZ4LO41hTUWziTe+HC09DYL
4Bjmmn2cWtOPc/MidGYujtO8cwGuCA7yop2+qXNmTxobdw7YEprpQmqKmUvWzvjp
dooyWGEvyZUR56KiQyUKH7huLWHfvk38GvQej0fI0cVWfbvTgUymAWnpbC+CrTwF
iaigEI8kebo+LnH/CY3ZvyBM4lk8hGJeWsjm97NlGNR2aVBJt9pqMydeWMdcWFzv
QMePTn+xSwp90pPmWS0o1gpnyzDThbRqixEXoll3EUicovubJacj25mDpCcUn9fw
UlSWPn/tHMi8JmcXgnGWjV1/zv+WwtVJfwxVN6vrLbhTCPgr5oj07R5Mct1vCfi1
fvBijHht9kyp/oQJlwgwdVRfzX7Vj1tuhZu8DA7o9M0WxhDFhVpDknbcUBs0eKfF
BE4OfvNLkSGbgqz1uAkHJ2dCP6GsAIHuws15RlhgY+cPFu6161Qgx/TP35B13gt+
nvw5M5GcQpps/tmBHjIv7LpT2TNX0uzmb1hpYUb76l1YzVEthSA567yug1Yv8mRF
dk9VU8qxLIiC5pQCmpphpynjFbayAFZmNoHdvOZTvanb0wZZI0sBudHuQZKZJ3NZ
9dBTqLLONDhR4/3bfJLtnPZXTfv8njCBCRVyWe8i0jPmnCEf4rSfD8X7mrYD+Ble
4BIrJUo/P0SbCxHFiY1jvCf4Kg16C0r13bHhCac9jvk/UMkTLNjOGe2iv7zNLXSN
rNag3P4VTwAfuOk+HUZxsbH0IZXAUauVzXF4Y/P4QMtF8N6LhM3iL91vI4Kf7Vvy
gYYAAcx3f5+RKNP1X8Gs9XXtbBwt8BrB4OTVOI7Rg5fv1T0lzojsLgM1YED+a5B4
VEaKXEYhNbIlZ9wyd8rBCjG/ziOCTrX8SOe1yDWcCQsUwFJ+ti2UnfYqXA3dg1SC
2xYdaRNmgPlfLXHO+YlLzh2XusYxfZ9sLl+OHNNX2NSGfGMz0fd1gosNqaE+ofYu
dc52hle1WhJbxwM26tFZ60OenDShvU0ahqPzs8MoFii1JznPLxE5ZR44bcvRlA5s
AEBUujoxCjMhu90aDaCzVbcD9z394S4pIyCfLH7ezYLAmJM700UXtES3vwjY+cxq
5oSjF7kxgyBxhZVSMlArV8AECF0ZQ5PafD7CxhUH2ETDjFRZcnSIYCqiGRV35tkX
pOb1ehD8F/q+REhhyX8VFuS+blizF45w7a+VLY1Y/CvvSx7/a+T80QURx6q94yWe
YAhnhmKrABb/yvYfFv4DwnfDLDocp9M7QJQozWBNPl/6wud9xrts4B/zYGdIhzj8
iKA/G7Pj2jSV1P4m+a763zV/5CAudlG5dQhHkbQx8EWB9JhASfgKGQ9Ssq7dDcZN
y8T4SvMcTmDnAloaM9OjZx4LDZF0hh3Yx1vr3mbEY4g5aL/oM1FTd22Q/0yYcr7L
UTIy5ruh9g9UMUk1bKtz0VgJ4/75E2FDF70fWlDoFbN5179+QPEXmGSxg1OHREJG
MVgiyTzLZmkTFfW3bDHk0Vbdf8SrXCpJbaodKqtCmI7BC5/W1C6JdGGI+0teWOOy
tkKxhK+EHzmn5C+cLFjHwKOyndOE+iYwUb2xij+rKbYQhKn4gQawrl3Kd4UxXX7d
GAEfe85G0LquqplNGQWM6v55zB0boDGziQIioQPicuJtW6FNw+wH4+1sIBc93qKl
ajaZhfKaFmg+2l40hUX5PPrcON5mu5DpIxE+ua6paThsU5v4bXbvWv2/Ohg3SbkI
zFLPYhMNhfW7D1NEVSBtpgHtFDJU3xY8lrTJQ/tQpAbiGvkqoMt+ysxA7HxYuKV6
4LfQ912FbcllmWF/Y8DTnLcu3hBUjUc+y3lfvQ2L3SDHXXDAPITDMBjvNZhXr/xs
3JVPFCbcFlpOZGfcRT0Bx/5UswKCF9HCHuia0aN+BucPF8cNsPng5WB0XlRmKldE
XD5KE5uqioLImPII2bIMQGNLwFa+QOInBnq6AaHqd2EcXPkkykyT2mgJVKx9ILog
BSTxTYWkBsL9E1/6E5MwWyfRw4CNwUoxUGCT1358WMykTT12Coa5Bdw+f9nhNQOs
C//SL/gm1jsYcEf+ilRm+km5QNtaUa6BbFrXCpReIXVb2SD+9HaUK+zX6wkt95Pf
dzIMrfTu+/OyDDeVxXoR1qz5zm07Ae9zo0YrM8I/2fWJc4TMOZtc2o++oDHDJt0X
Aqoh7tjO16c7HiAKJMsUxOAcWipYyECXXavrsW/3CwGo6dsMbjqmDA5KKXv7OGLB
N53gU+TxILfTD8iOp15sJx5oPES2etwGeSabmWmhzmC4o08ueMtCtoS1bbGo3Co+
2kxEIG0D/3hZL6SFASoJ3ZY9ac8R9AVJSAtKyOlj66PC+s9xvfi3a2/fRslM5wDc
NqeKJCgqLFZhLgsla7LUDgloHmbdR5mPJzS17P8RW2tKttloV5QWoJoI1Kmx8aMh
6UUMymxkopyT0oIGo7mO7vC5frhPnY0tsIZjbA21h15fD//kmdVEXX4uXus8kUG8
rCK+Q6cHalgM7DAAW2EOvY5o3ZFicJWE6mUILGXZhbuLa4gpauSo8Bg8KuzKQ0cm
10CSwClCy27B3Lv15/EDaX752SeASFr+Zd529m+w/dZHRni4oJOhKRF0gZsmAoHr
q+ITpFeW17GBQyO7rX3dndBa1bboWYUPtnOGeyyPw55hANcrb3Fb9RFoSWWZ+QeZ
bgYJkA8Yf7SzZ1P+cPTiYCsyWCaJyhxQA8PmAx4R0Mx2eTNmD9tGJOr54n1rc3HT
S/wSSJCmwqfZQMbqrFL8AG/SXmxIpE1M3yYGSWirP7xuJ2BCcBg5g2kP7OU5L4Xb
OZPr8rUSzrtRKDgcg8m/0if1GtNyZqEHn6caBVQAaepmTBq17IHmQTzOk4UkHGsQ
MBlv4MNysqHZm5JUew5HXvVNG4PzXX9W46RO2UMGwsrkFeD6xG7cW5nF7DA3TIFq
rAnFh4EpS7bhny9OpgzywNzBCnVbt8VfwbxXsDoeJPh1TGDUxphTsLqgX4x6NqcM
B2y6urEh9WeQnTvqq3ZoafKfT0Bdfj0CSyHN/Rmn7s3vbcsfzwBk0yWypbrwx90R
6rQZUf24V7M0QN71ZfRo0PVLlXNh88MoCYqWYmkcp836dmTdX7Y5rBJFN1c2vmc2
65KjO7leSG7tKb8YOK9XQanviskJuIAQwyewBH+LL+jmuJXsK6R6zrFBXVwQXPs0
0xWek22oHmnFek1oyQ/2fH6CftxyoXRr4AXcKjnaIuLr5iGSxHXIA0NB1FqkguBX
/ILjsMbhfidi0iD4L0DdjKwryCDeXtNHmMbcwVI3Ugmf2uprT9T/sqraWVWXyMB7
mnFwqnzGUWD+2HU1Tijsp2iACNCgdteD0HOvY67qZNmPCSOsAUAYQyh1oksH1IJ6
qIzRpBI2ZnoWwM55I7psJbUlqFHXqKEqiEKLrM5CRhG4jpRmM0p+YErUNJsyflvN
EaIIkwth9dLAw77rz9Mmqct8yiKwGvC/Y2s4nCiekHQrCjzAK61IIBrAjVANlG4h
TBA5xHOTE+WkuqbtisGpwg==
`pragma protect end_protected
