// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:31:44 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
sHaobEtx8VF3JzzOdonr+gwYiO6zNtx5gH0LQhp5OLNHVuc1D8DU11kdvV+ztTrz
MEC5J1+o4u2Vm5JH82FmIuuk/kN+Grsgu5LbcJY7YJiwxaV1BlL97nfHjXQKgUWy
duJRre/j9ai30yIXUAaKbbkL4d45kwFVPZefqjfZTzE=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 4864)
kU2+vGrO38YieU47CdB53v6Qysrwk5J4NTzEdfuyYkOXdQvhXmBgWFEPAc7jZuFY
kJC4VNrxT+PEV2+GvBNDR7vmXj0lUGJxKw/uZs0pbVh237H9VJftJMtd08gZp3kD
TJry1aRiYy/VuD1sOQfF8vf03xxSqqhHnqdNsNgrU59dWD+KrU77OqUMGqL9M1+C
yYSErDARwEGBguM9gRB56bwCbfEFddCBbbxekWyj11NidPHyJZAhg5hC6njQybRd
spX75F7jMDUwAdOLsYoc4XN2mr0scuSKD+ZJut18ZRuFkTxuLkFl8APefVVfTa4E
59bnRhUMfWROpOO7R/r8nu9JIlu06w0+ugRqbjCZfALAM9MeL/tqnua3qZkgzNMc
jtiVYPO3pw+wDC8Yd4X5PZHFbu+9mqJzt87t7ecGk4gj51YHrLajwrNhRCb2dl73
T4rMb6Dsw8rsCFb01YLuOrJo//frLNi6eNjnP8UYKSu6wPU4kwaO+SBEIa5U+L9c
f4dcLq0pxctqJAOQ34W5KqXprKrqTfxd0m263vv3tz4Ht0Y56TCUniFjfHcdBBVQ
F2RAYtnTwaVDo2lmSRKlIhErjfe5MjHQRMWsU2Zj+IJvgbTTEot763YEE0B3eddl
DRhwxsI8FIAcCwtqmwBUj2HnQmbWwaJYCNr2xKKDw0AjtS3gWduIdi6LprTRD4AB
NtYuMJgrnLYJ6xMa5IeiA2MXEMNnYqw/qKdfBaV1+lWvgD470R4sGbQG/rtU09jw
soSQQU82fB2onANMib6mYyfNtBUjU6HIMe0VDQlvhAAMQwydK2sZGRyaktQKegd1
VTOXJ4MMaIqT2LZQ+q9UwWfQbybj1RxP8BLQ1GDmwVVvDekhdbrv+C0n/Kd3+ATf
JS9DnR+Ke0XnSBLU5QtV9SYdjEUjUZsneKRir0ycAvnPwO1p4lXDkNUk4C7QrgUZ
9Ot29eeWQIRG++F5MpS0WfVtu7VQVPYCxnJwPEtABz+skmjStESSX1w3Kqe0/eZI
fho+alGtbo5vuSD6yJ7xXYpQ3e8X1+FDScKKQlSfmgivxSKcX+NnZE6u7uLsm7b7
SKA/bomiRBot7rA9sPg6K9/2B8biEXjYqDrdcO4tn1sTljnKU120VYd3VGntpo7u
gVBHbu4CGi5KgrfFeQe01o+zXn8lNJMTZ2fkmTDuizr2i78H/xh42a8iGOLA8Ixk
j5hisZiAWv1BQDa8VUQ1O1nzrGEfoOP1xCLGgxN/jm+NGhA6w0ai6gxexd790S1x
vJkWtEqI3r4LWLbXUBYMhZyu47k0ujRxp9UoXTgWSOnF14ejNTRG1GVHamcg20Uz
DkPgn+CU12mGKrtA8W2z3taMGtxJZzhoJY3+dZczSvxzBhQ1XLqg75iwJGBdrbhb
Cjut8hO/+lDk8lAvbmW+QYUN0OZilbQ91OXjvSGYeB0uGwAwgsQ/Yl0+xSUE7Eub
OQAVQkM1RsQVK0OPCphXOgROvlnxeTB7Ah5yL56Rb3QY/ZZR200yQ0cOcGXN1J2V
0wJYfkgSzFKjh9jRxxBYjK44c6ToAROHu+2CJK6KCoT9eHM6NrjGadpxGj0vA91k
9OM3lWaxnUD502RbsxTgQ3btMZ/DQejNzcHAD4YqydzLSSXMIV58KIHUtVQltM06
rdobbaaowILHvjCYdW/ZVjkKVaD4SKKCjgcn0+9WbH+9q6yea0DwYoRwujaK48m/
8HRtg0ggMvA3CFED1MkVZ/uOBAH3vBLJMIyur0yUJxlL6eqYupK3+/twKCi77Stj
9cb4o8D2jF6yCG/qWD0+la23R98yJKYuKtMI/mbUYuYa0UdbH6N5HhCbCyrbHJjb
8s+GNFbiWRs0vyC04EFJ34p1YzakA+ByGZIJy5hfBiY8Dik6+WlaPeeVvHSLTV+3
J1yTHE2Masuz11DQaYejgX7eFew5dSgyTIdy7QQ5+vCAn64z30D7qe2CLaLRZK70
6yaM+D6fI3WZnjTVTMJw+h4susViqmenJ6cpjANZs62GiArNYk3ceK6B0t/Ih6CC
37sEDZhox9xV/YCTjLnD68U8sD0L7zk54QO7sKVTDvB5kXv2Px7CePu/ZFgE9xGd
q0KlMz7t1G/W7JYikrp/idxZtHBX2gExTWrHGuVKYee37cZ5rS5qMs8JmsoUE4p4
2bgX/MuHpB/+Z0X4uI7sWTCrvOIfh/rpSjKDAauz9Wlk/dhsbFMfwSI/nyPyLOJC
RlgN4RIdeDvk3AIC9/YqC/0zvfNtZvB93TPRHUFguQ9nEnMvN4bhXEWFlA8qTvLM
d3VU3eiO3Aj3b/c7nWurIuvF5BSdG0Qf2B9hlAEAbmYGhfZpHBe9MiOJaioYmbci
mEbkGqb1J1FlSCx84jxh4WIRG4Zt3VdIHIRSeNV4QVUL1wKQAAzvw6v1mrETZX6c
BKjNvcKgHsi16cd9cgU+5mB0b7n+2Y5hk8VNOx3QsvAn3zidaRtGwVz9MgiMpmHl
s7PLythH98nAP4Eexfz7xC7QWh+5LSydjedfchD4VEL3h61YPMSsDq1wYMPf4oXX
TVW4wfr+ieOF8eEijk7NcalW9gajOA9JHWdRKfvUQXmAfYbI0mxrUvDGQq5vLJ/d
Ynx7nLvzc64o8LhGQeEvaxxe/AvbiVIKumuGgUUziEhaQ9EEZUlQVbTgMeXNv0PH
H56Zf1Mf6HvN6K5B6JtQ8pIpjGdVrBS0ZjolJpMTHJRPD5maKfl22qcF/NIi3vPI
ADjqSCyC1X9PPFspy4fgorRVvUtcDNrEIBCkopNR/np5dXxiI02CaQAmV+IrctED
gJ4I7srwEJwwLmYj0lvEZvHHlkCHcoVMEZTnzqxutLdxZMqprdt7H4cftHhE4Th5
tLp4o+8IYHOG3iecQT3zpM1tylycAxCaCvLQQp/acKvOvthbzSeqzryxwqybFasB
59SCC6QZsT6odKLIMq0PKEvP48x4kM0hIBG9fJ5Y8EDS2YjMFqCY6zOlpHLAt6bX
sT+rPRUj9Jmh5AvvHQjwO1jA2Ut8XtDE7uY1G/pOiQbiFjedh7fB3ixmfbZFA2CJ
jLnyeglw+bZCE14e99isj3g8yR22GOdWRR+D+Do1CC7xRJX5fPql5lAYn2b3n9lU
xJLoq7mQ9V0YILBLu8w9KjgphJfhIBRmiedSJLdi5xmpKFIwl5mfFKqD21/VoIjk
JkbMqVPMMNunryiM5/dKJyuB/IxdndO8g0jE7skpkUa9j5ibXAfGZr7WBCLCj48H
+v8BQNne7kQP3O2FVROpVB3YFaz+DI3pbvHA/3CTUpLoUEXcADDruuGI/9l3bI7b
YS/zp3bdpmjGN7vw25GxL6CjGOBQAC4J0y7gacOmt6YEo3Mn2bjRBfc37Oi46H53
KLpke6y/TuPtwT9dvlLf/AwzOlKZIMIXLXji8dT4LOZnTRJb+7s3Lno7PUER7N5l
v7Hcjra4+jHHhZthHPTGhY0xQLpcLRZ3Tn5oBiDzMx9lzsg4wz797qXN7IqprjDD
YYQ0nSAOeZiCKgFGVSjYigfDUg7CekzICt9u6zq1UEI+A0FEoUeP5SfLwYMjaM1e
9pmoEfX7xwYwKXheEkZRPp8rV8fYslM4uUurSLT/cqDS8VYDSiSdEV7O1ARKK5bY
mpiTIZ8TjESkiFpvzV8ruY9d/5hza6XJzHzxBi70oLbuGRP/VQ12e1SwVrQoo15o
3IYQex0oLiQjn0WuwGNHWvytBY02TtbWzzOgfxIefqWzTMzg6T4ybJCkWfsWUPcF
Tg2SE6iprcduHzq0TC0+ltlKITbCQaAaACRhUYZetgXA0cZL0VWTuSrDYmCSSTwO
siuKfXrBrrgkvLXrDTB1AjUsZXg8DiZPrMUaQJ0zOCDulHu8BFD/4ytWBRqZSIhA
eTbKJ41WfbD4Buziapfd5bU05A/HRyWTgoRnXc2BCXhthGWR0l965qd11K/Citk9
8BAA0oXoCSE0QtVYTHA26zoyXw7JzR/Ra10n1spw/MbMVqOncnH/g1zYyMqcqAeB
44aoFaHOirpN15ra7R2NTArlldzGaByz0hpzAwFoKVbmHg7om/A34vvdx4fNUIk+
nvGXlTVRuKT3VejL7xsd9KpzmHJzmp91xfIJyC+eMljWRbzkb4/cSa3KPveyuwxp
xrdiCtjktIEJHJ/Nv9koXjCtWrA6noJ9YRv609J1/RAqEUAh5zjPQDdqesYal3sR
lbPKVj1oVIccJifHTw3NG+lB2ZFuAd3TK6UiHAbiuroUKaKDR2JTuDTISiHb5ooJ
7oK/aNg206752SfEJNagOoItFAIYFWWayQfi/p9gMuplJQrWfjB4txqYtxtzEwXy
7EtNXWb/cAIHuT5+aeMHBj5wfdu5XgwINQ3jDa1jIFLac+ysAZu/H1lYuN7Hqu/t
NCjfm34NtscEotoY79EOqkr2t0qL9r/whwoHtDVkZbaiqxTKZb1yNE+dvvupAUQ+
eHBrwVKG6jhfyep2uCZcy5AgOUXzjKNyyiCI02YQvdK/0kgeYIw/FZH+LCy1bQyC
FzBiMlZIp46jVLSpHyed/Swr3GrWoQZXbunU1VMAhsqsRAtClZ/Pxh6oiySoXaWK
BmsW1W70oqSByYtoHF7lqUI13xF3MECxPyjrOORvuWjPELVd4KshchGzG3pPnSPs
UygNfa5vzUb3hT76MhsGfbFtzoVv3e/7amfsXIaV9Qc9ohWGL1yPEUe6P8cVtBqy
29tXxTyHhRq0lKwKn5G2LdQZTCJXFpNWlzuC20w0zO2AuYLbPpRWx1R6NvclQYZG
6Rs+IAWobR614IDJEeXzCIR/0BJMsAumHvs2ogcAfqYM9m9yX28GPPJ6uGnargvv
ZdjArpTA9LcUU3xFrLBO0jpuwqmO/nb2W2UYvzBJXV9B6emFcDfLWcYSPH5lWH39
EpiE5CjdGvqYPsvSWLiVoAYP+3NFayJlBFPi3XrF+NIGvt8Hg9dQ4opBYl9B6p0z
z6zterDoGkzS+vckFwFQi7OEwDkbJ+Cm73K6oUFzdBMrgIMV1V3oh4xIVLpJAtqd
f8FpweugzpZz+29ACaOhGXSnNkpIsi5weATe+RSXPb/CVZ2L8s99HsLiK5bguFyt
T+G3hiWeTSn684K3BPe94ytJxsaCidlk1DsM5JqeyOUe2gmpj9tg2AIaDgiWod2q
xv3DOcCqzvtX3NlkKVklkikxFpnqMf9LIHkQ97vp0ksGq7vafth4vPA1Nq+gK2Ik
+k6QjvxLeyZrAq75bg2BkCtMVf/OtL5VY1LdBf/ZBbaNuP/aXOcgRBhNeCfTwciT
w9zceqJl1IOYnEWmK1JO8zLhBwD7GMnB1j41NLMCAzMeogQMZlEhc3WBOZAq093Q
i57Upw4mG6NOzQnHy9zbKAywM4DrYYbXcq5DzuDG0sAYVSfYHwGcMVvRmxYBaDG3
Ebp6PlhXRlMcD3KYfkVMVGqY9sezNTmjkwlIjeOkq7abGR7XvPsUsz6qDEwHKe8L
rT+CTL3VUYoK1qcJdRZvk9FWl7WkZofdlG9rAp9ypHgCXEyxN5vjmKWXh6/FbZ97
UPYaQ/dFQ/CDcIo4pZ5f+ynv9oRLIjCs8/k8iGnlax0K4RFyfNpQZCdYIEyjzFR6
qZVgeLvoDKSnkpQzeblgoNzmKtXP+49oLssZ/tvmCN1fJooGFEMjKDP5UwMiSYTq
2chUYCuSOeOWY1EkVwGZKcDixZHrDeR1Vynv2Tb2kwCieW9zgowSOhHdORnTVkiV
WkfK+VXJ8LSo4L6DM5Dcmf3BtVkOLrbD4NINkVZjnW0LaQW+hk7fUk2s94cLNrzx
82lVt4ZJTk0Cix6Hdy7ClC5OJsTjMGnfMbxj1D3uTDXe0n5vTl+FLY+i+w43iWSb
yT8uO9twVjCOzwF4SwWEZF8+4eZzv5v3i4mHFDeJZeaWCgNHDHKdemwy1eGrLmVE
c9UxM4GOv0pv9ZlVV2ajBT2RiA5PymZ7Y7pLRt1f1SJGa3nHqdxtKuCNVdOczlQG
C8W+JNDfGqMDXBxdL9HZ2yd0nmUqBqkSonNrk2CqX4V297YWsj7i1Mk1Jxatelft
jUXymbuPaR4C3UGu0czZMwtZ/fLm7SL2GB5/L+H/KzNGD8RmhDH/twFA9shoYOvX
B5jTgMT3jlzhLFnVU0X8OG28/hblNoIpuXyDe6vTsTT35KRasfi7QhEV128FMSMY
aDMG4oji94EuHiG2iv6mRKURdL5jl1WzKqVKtaQaUN6axhyfgq5pP1kmlKT7zeuQ
xpNuPcRRn/hOJH9ku4xsqLr2TnqmS7dyLytD+9Szbo1EZnDQFZtZB4rL1BhqKPXV
uMFCA13fijDHuEgWBSXxSsxN+l7Hbexf434hNABGo5n6sNDDJ6IMjf8Q6SapIWs8
ABUXCyiTU8BR+vdIipQYNv4ftI7UH9PtFI3Zu1UdbcZ300a8Dq5knQigx29yPio/
CwGVQqSQu3Swwo8nFqRtGw==
`pragma protect end_protected
