// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:24 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
HnInvxzgwBM4pWmGb96ykkg+tb2W/dfguMpmvYhLM7Aw66A/EyGt2h6lU3wgYl9p
9uZOxAz4fMT5YploW14il9hMxHXbB8/2vanHeWZ4O1noN9F51Np3S4T++bn2+Ghb
QiuHZlY0Uk104InLBn3p6QoQxoHGcQhAcP093/C4/UU=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5904)
v8xtvwGekpMLu4sLkpmjcq4/cKYyp6ik3Li+uOdm/B0D/dgHkGc20275KwxINCXP
oRW7epQDPfvyFXBtUquQAtWQJPcnDYqsRnYYCpIwD85tb3XggqThmHKKq6exnwg7
TycNrnfYn5sMGuTbpg8smEmUDgUJtAfgtAAn57VANtgN2ylJbpOnIxfUpisjj4gQ
qtjsRgd8Yd3TrAbTM58dlIZVBh+aSPW03a1xD5tTjV4G3l909/dyDWp8s4Uv3OhZ
+2v0w73SopqWMX3+roxNvOf3JXuqGETb++tjb8XCdOdAkCv6wzaE5/MyJq5t7OAS
jzfoRHcYeUHBVCsjcKpnJoKq+J6k813iwnq+PdAkQYRb8aLvxU6Ry40qwXoU6eKQ
3RyWe+rIF2yq6Jy5axHlQq6e1YOyCe1pvt83cgX6qmrWX97F4pabdB1G7gocz556
my5SkasDw6PN9erwmni9s4CGa1N92pQrv9FfFLBCY24JK1p06T8OAUr6/yZzHeXx
fZUjX+g4ctr19MLUXgCERVjQ37r4rVeB0Ax4fJH4Ih/szAGCbCvSA70wkwwu9dMq
uBm/HWc4LYuHP0qX0Z2zkpjZ0OT2WAUcQ4b46QhHzPa+SFQV4MswLdlDcr0+S9qp
rpKBnWjxCd1aEi6G74tvDb9KjENEOKcLt3COrpM/SWa0Rtg0zrMitC5uffRn2jKY
6NMhXKEdz00PP9/TJM3kq9Lh5vp+FRogtEuvjF1fNJJ7Wq994cgvOdbYfWW3bknV
76crvu5nnrjoa/4yrjUYik+4x1lsrYKlWqP83vtr8c8Ke+jVnORkndKzKFfTR9sE
6SBAF/63mM1VjNsoKoICNCwjr9I+fa/TXm8joBHh/4e2BQ1eHUHi4WpEeiYfDOcO
4+eOIQ4CBAKOZR4rTlVE1eFoXweFndFpZr+8EQwQRjqmCR8LE2pHPvMa5l1mFWWz
U83eCfK0Y1urRShhDKvdY/lhj0xa3cbjZpb2xaQ2d5KmuwIEVGT7Anskqe60aA98
8xbAThQVuag7Jdm4TDKJ3/ahq9biMHECdEWCY/7gBlbr+RtjG/j2YMJ7artsk3+p
12nBSOYt6Ruokr/ELH0yVYOaiCP0ZB/BvS1Q80gmvNKsIHPjVJXRLw0QaR+Wp+u6
+dg/6iot+j40ZLiOu3y5uYuncT8xcR4aYG188LTbURA7QTK1fdr9zxNgferoiKhN
ypXu0lYWqaax/Ha6BonV7JsPolTnNC5Ptolk/7uh7w1SlB37T8cPKfs7E6OJCWXD
YYvFSpVwIZMBSK+jqwznFu0gfOR97AcxZBSVwzgNYPo6dM+Ms1gCZLMxM8V9eDQ7
OWo/8J8n1tIQWtKe99uAIWe+WP/fq4/cCOI/uqRp/tnH2mtWN4bmYwjw9w+SzzsV
XJGSTHY5G0IHRhtuF/qYQ/V+qDGawoy0Ldya7uZgOV+IMnPPYhCBdcIB4utRe1AM
bOnmAVJgh2hHC9opTp232wPrCKmB+Ea23Guy0QjUG+NoPyUJ7+qnBVnRb0+UnDm2
NsDgxjzwv9vf5O+BacXHaPMnBbeyzEhbSGdOsbXBP3T4yprx/5dMu1JYONa2319/
nJftBxoD0DrUIkF1lal0ACbXB311m+kED3v1dJfMu4IGfCfmpZiHoGM/EDc+RBhh
K+zsnuGrEYstzpR7b3bxBKyswZ79OX7Xhvlx3OjmRggFCbXxbVkdN7/05fcJMuHM
Ur7Nk1k2vPXIPYJYBvpZWUt8dlGCmpSZHcRr5HRtKLlUl1B1lfRaEIrkH207ZZ7x
VBF4P5ZDX+lor3MeHGeKiuowpGWsti6o23res6qd9hA+r0m34LVE4FfI4TdC8rcp
88oiUwHvBdyzv4T7VQFnrb+txk5QeEFBLa4CQk6SiSKJY1nRQjw+euHAr7zUM5OG
DMb8lSMFF01gkHRNmNTtzi51QzsBja315RDm1BvCVUS9vQmTqXSx3U190y61kgiv
gZz5w5gnrIMvUhCVOOxP0RiTmp3dRgEDLckKNEeIoplBGAhrPyfKNKVWBd1w0b2j
9DPO2eVYCNwB0bae6J8WPWpJOk76VmmzvZRAiuPm/y0Jr9vncFOgu7Hia0HHina9
eXBTuyFeKMmZqGVpfkBhtjg1gWnU+7+VfogSZQCXS5r2rfLcnCJD6zAK0Tynj6nT
s5PnDZrV4uwk6uPMpcU66BOJV056L6Srxx/iWa7TUuvnLc4S9qSJ3bR/FSRS91dg
9/Q6saVzQzSg0AZrWCX9PdKg+gDS8MQ45p/3uZ4EIdiS7dFdwXOdMzLowhRdtpcq
dJJBEiKzfIGt3bzYQOPayXO5jAGpDQ3BTUjpg+f5c9cdVl54mP0DzikYdS7lNLKk
PEmZmESVfTuaV6nAWuUiM9e7RoIIoMeDjzIg16gvg6VITul9z5Dzn3ZSEFpNytm2
BdP2pHcP+2K05v/Sczw5yclzxLjzhEEnOcb/wkrnVYvCJwUTCzG7xJOQyNv5Ao7g
pUwqXqQV9hldOPiItrSJQFvTozPo/zbnbgRPUPkyHPjMhUzv4Ofhr6EDJVrFdtLn
gTp5PC5mZn7IQ1O+bNyJwdx3/mIjNz2/fbkXNg4qwdoDvEdOq4WIlbvmf5gy+caW
HdI/J63IjzMqjJLV2DB6EhjsED9lu0ouG7jCm/6QSf8tClx/HOlHkeuYDncdVXvp
wkVPzIw+r6eshgPN75nuuiR8fl8smPI/aSTQvslCP5KU+zasFhxhhVoKwK1qcrIa
5OfnDthMEtVO4rHHrl94Xcd3/gf7m4vBa1eWNcYMn9mVsAP+/oYD5OMnBRHyZtsz
d4I07FFu/2DjwD+jVYrkvqKyxQaoAXqlirkQicZcQU3/73tX+V4ZxW57yZnHEldM
SC1K0raIHtzwffOUJyaLp/xST5ULUHl9brxaWL2NKRC0R9GXylA92DO5UxWLuZ/Q
T/2eZ56VZgnC38sqn8NMWXQg5aP5s4eXj3c6mJZkyQKB874cpv+IgEbdrPS5wPPq
EAvkPFUX83FstzGgDaSXKfttB5sragq10OzhJeS8K8AFmszkdH6/IPNC6KHjHnrA
I2AhRy3ZBNhqsLhp0rWSl2CxnyngXc0kpkMZ5Z/ISbfjac/QihLUY+Ngf7IMFKH1
uhAN3QndyXSzss7b8KwUc6tV8AT1MVw6JqoSRTWvcwpGNG5jkSY33IFTOfOvx2Oa
DozNe47VEpm9vNGdoTycMpLXR1f0w85/krFVkkwLG6LosNTKrXKafdHWsbU6x0v1
gbIVldMAJCbLBn5bPxK7LGZFaU1vihAUFWWFFjVwWBZwuvHkeAtkrHeHv+fRgcxD
Db3c3sgzJb1vU9iKfyaT5FeLUKhiZbBvE+Be5sSBpwTWQAYezerf5a5/Y/LOEIp3
FoM0mXpyQ94RZ2h6rCPkIam48TleiflgBcr/RgpSCdRTBgfpW9XWtc8/vsuUS+Li
Bstg0Vn99pvoWsFYYMaNlKRx0OS7FYWEA3I8Lfiu3gTAqcJaFwzmqkfniTxDOQX0
UHi8p4WXzBPYg35yp9u0BMNJY0ywCTk+ol81QiQKilJ2dkh+NRkqDnmZQIPWChHI
hb2iO9GIdKh7xLs+zQSBEqkFjJJ0o1vGlIZRxLn264Bnz2YIFSokJ7hiGNWAi8gJ
l3Hl2HYOKagV00D5kVYSHIlkNs1FPm1ABKwJaOVfNls5tFp5YJmNBl7S2PUH+wns
zSSnLTi8qf3auQQ3dTnTaaFfJ0HvW4vd3tKYS/wp4rTj7VMkgiuirYVa6+gB4Im8
yvVl+b67mrdruWRd0g0xU4Y60SzbXxo8bEm50OLdSF2GqsORDZGeUO9yzoo+a2dg
3y1i/FF/mQoczy1Ui9SCtHZymepIb/IhJuoBWJRiGC/ucn7asCXJV+fZfIaHG/b9
qL7ilOhzPn935Uo3e9Ke2BmVosQv/KMTE9GCxdLIJ5G6PkWQPdXsMBENIYGVubxG
YSYrnv8z+JvwlKLEWa7Vd/JLEhhfZu7PDHhY4WVwmF0SpYr1klcNqDjT8EyICVG3
UUXJe3u9bkz4nB0gT/fNPeVCcuoYQkJZFRW09lbXVuq1puNi8U2Py15gDJr0hxMw
Nclgry3OyGgaeEb+8lU6zeSpqmNq6IBGbb5MdCZLZyOnOrxyuO+uFSKPN40G3ooG
XzrNfpY3x6VurjHpWTmTMhCcKwwEg9u7iMOp1B7uWKXaI86sJm7LURuafUkoWG11
pV9VhrGDA3pvjfrXlEOoNvfAH5nktF8y5ybyMXenPVj358kYK0dbwFjo4M4/ZtoJ
cB+EjZnDVNs2cXD0f4OXiAO4ZqVz814c4mwcI05OrDuOjGNXWBs7A/U6BEJTGUbu
jLAcY508DAZicrjDcM4Plw3fjC0jy9BAA2Zx2l8kLRfp0BoAQeEcRRCQnWbV6luP
wLpvSEFCBMyIF88HtBfI43eNBAFu0haeRTXE9aI+P0wO71aY87oQANwGKoeIaNyT
mBtZZoxmHfyX4/JQ+jmkilBPUhKldOVB59e1aGGCZoTnJ1jb3HVMu5AiGKy17Dec
PjTkT3ihKZZeLRZA1yXr+mOZz14XSToT7jUYgtE4fI661FsS4Let+N6oAGpj0Z3z
cH2SvqOik8UWWvLgMkSudBEIbc4L3LhJWIbYgZ4dCLWypt816PQOPo2Do7B5V644
NyTXjtj+/k8glUUakV+fD9xtivRNvMzXyrzXuGn6LK4EgArdEnDoMuW419QK06jf
IwAhzJdbMehU0wRpdryFxxwXcNuWtkod0BBuoYJ7GJSbwLASNbIl3xU4RBm61sO4
n0E4b06lSzX5U3NTqo98p/daDF81wbPokvLVQKNTqLSPlgSfwcg2KFGUMCORtxnj
s6JGh0sOW5Ovv7/e8mDNQUVE/D/kNvzw3EsqmrFcEoO9VDw9phqeYUDz/TpJvM91
yxrUq3+F2gpSRyNREWeXhoL3TZ8uTW3DiigR1VeyQv5RXD6exuwqqF4W1kZ/0TIj
18/RgooKw8xxHAR08Xq7LfpLnrfhXDYlwKho60IVi1M8SCeZ5e/Ceqga5ny6tTkR
hwIArPlQrec8kaMkL1HwZDPUDNqCVAgeHAD3f3/A68JHeTcbOzilYryM7+mgWrNI
uhKWRyCceAfFWsz+eH6k90lTkM6f7nTvejO0i8D8JhLOBylue6LjP0PzGJPkU3YH
jOzwMqj/FLlQ8bzTEqNAnyeN7WR4VlPaIz/u+vPSy9p3tv1+h82UxaEBahuFxes3
90sW0i8mSOkRGWL4lNaC21eXvqcDmiBrIQEAIhQvGtu9YQEtGtgd3QdTaMCjoFVM
/5y26OL86CxNxY9aJ4KXUq2auMz1hYWIZjs9fvHPPv0ss784LPiWsTzfGrxNklvP
ZQxZ6Y7tK0ETzTsRNl4RN5C7LLAvt1be7YcuG/faIMhnXNUhoOvp5FB82lvYJqjh
03SA51wb4ha+eyo+GSGPmfQYls9bDlUM7OAftU/RWitQDXpjLnDJwzjlvchur/4u
Xe7L9ohplOKIydYSdKR/LAyzEnUIW6vqxy/XxTSr/TD9gBURN1blGZXE7YvhHZG0
SSlVdQiAeVGQiq5kuC+loMyEOij9IwOYXOgULcJxdEo8E0wHAdrbuUEP00pEN7ol
6rJKlguO/OrYseRtxpAtdGpidBM72GKHEt7ebCNTkHPTU6riKm38RpdgkLYVOV6I
rH7+ChVOpe9+7rIX/PAL7QMG6VeSZzRoaKmxTbpJS4a32gq0d14+lbbhp8ksvwaQ
BNCZDt9BP64dnIAYKSTsPpYGhnr6zwwy54aXCECvKAstJVFTNyROGqoN1fFS4r5d
nTNgqpQkjpR3eqp+jq+5deKEwfxuTtWJkKvhkT/S4n9R5f9h7fYoxKwb1FYGHWCJ
VV5Xu/2dm4E4WF2CwUcFcVMSggnwmMqEovk6ff61h6dAebw+/QV8uq6GzPDZKRQG
q69S5o+9faQu2fTBQENh5mFxmTLPmj9jgw4hN8RUS3MDAto5qk+8YJEwSBGplw5Y
LOaQiWhIRVDavbFY3nw2G2684kIqGwlM+2HwPj11Pf3evs/D1QBy+1ZW3bLvCsoC
us6Ap5CD6nRTR28nrcvarxxeY/L67O1J8pWUeCDeNAvjGXR3sey1v+ayx5CQczos
ZhHquyC5N3JZEVcO2ip1w0rhQoNPiaIucSZDJtTsy/Dy2DOvFlS1cCRQWU7Vin70
kNwmCUQwMjqelRh73Ni3Snt/FXEyQC9hg+cr58sme2C6vwuZpWr10PuP7/lvrLwt
y3iWNNHRlcnC8xbginarvzyht+qLciPGhZ3y8r0fkDPG6yf3uWl9ksr9aRCzSBIw
V2UVminDUDsTSx7ht9OXUtaJ8yggmUG9A+9KS3c4pVqGHnQccZg6QKqB4CETZSnt
NIo4RWc9QOYaZnGdEemhwmiNzxZn48OKaB8ZrjPEme2zYM6vqMtMxKVyOwHRqfUx
+qk8gKxZYvUYe77JiMb6HcfOvDoq537fN67DSwYJAnavOMPtjfhMvzuMP9K2ZYL4
zHYBHfu2cbabxMZKaE2rmdCL9QiVic1Q/PDDrOdhkYYpdSqF3nMyR98MqHs4DcTt
enzgqtEADHb7vd3ZtnSHaSJRVzgmhxDfUdaCt3GB0tfqiXzcSLpNrD/LPFyM1Iap
0Aunv4yl6+6ZnYtd6WduRj+Bw5booxRM4FbBMHe+B4uvoVXZ4kDBo2EqCKk0SwSL
gv9+S+y2XfuJc1NZrL0blZhKO5FY+EOLxUIBzXaNmdhXhed67mIJXOia/LKvM+pT
K/2V7tTFUNaIwpuyb9TUMGYdMVaoJjmovyOLcnvmmxKtfqePiLkTw0jTj1+YH12G
MmY/+mMWPjxW+GfBy5assdoO1/lZjDDyhOF7D85lOoOg2oNhP7e6NyfKK/rof+SQ
aNCV2b2sDOkYAv7kB/x6cWAYgzAQiFGaB5YV3Bwd/XxTccskV8qQp3/kas6t/tQd
p8qMXXpWjL9k95pZvKJ83twh31wGztcS2npgVr6wgOotEs1OW8331vdyix4TZ5oG
VGZEElD1+USQ29DNovwBT2+5KwApZuVqTWz/svVdD+9uv4k7349Sh6Br5FnFkUgi
H9rVAdbj4ndwi11GfXGIkkuikq70V5UReMxLcpwO+Hg009Pf7vJryxsvt0+MOuQX
k8ZuXWw4tKXAV6UVVQ7ocSPraeqIWogvk5tWcLa1RHs8oL+T7cHC1ydrndQy+538
gpFR7jAi8d4LmXuyqIcKbS8YAtGnChRm8yhr45TPORXrRJj740fn9QLao1JApkE4
wk3+Xz2RqdXmKFuaxBSWx7cMrHinGPlkufGaZ1Ebo6h7ZnNSkApCzfMnOotUWbLL
wFNsijQSOjEAvHPdizZiqMPTRu2QIIZS2dg3RDen67ZVrv/ZJscwFSu19IVQR0Ca
cySr3PWQ2vJu2b3X2+mRA5t/Fv6/H5cbgEGSt4TWIxl2LlzOQEFA02EST1j85Tb8
0OvwwbZ0yn8jjXenL5uGqt1/+6mtSm1k1hP063m/mp1x5n6lupLHNyuhcXzzPMnw
iCrEy7uImb2WHkuA2vZekkGX1sER87U33L20X6RNhj/3ihFInicNRgOJapfuI2cW
hwS7pj+CC7us5XvLkdXl0fzclA0sNCdEP6f5JNQ1wNq/EhXDDMSZy8hNL/SoDmAU
lFOOEclQ9NvJRfxKFDpVW5tllMzZOcMtt9IAgX1hopmlKZLHKEJ5I5UbxPOvgUif
VRuWNNA6VyCuDCbKJPOz4XS/SvxO4rjq6fGR19FrthwnF+k4+jOP04zUsW79bLdU
/nooVnLaozuylJHjzIKQOkhrwVq72re8+XaK6eK5B5wBNtriNcabZXK10pW+ZD2n
`pragma protect end_protected
