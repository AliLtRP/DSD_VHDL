// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:35:51 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
IPP3xpHDfdkKZuYux4LxyS6USEf4C5Yf4QepXujL19fwcUGiCo5481Ey4NbiWg4I
Z5aA2Yp3Z0oX61JxMz7INxXc9P6WtXQxDKjA5DH77DRUGOqbJSWF7GtMLJdWANCM
uSRn6zsgrzvAi8iUCl8/KpTNYBiRJrNbyXpoAru/Jn8=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 3488)
xA6LXWgZnFsPDeMo7FNbSqOexkP0k8rMcXcPjjd/5gRPU/+ZA5uquJSSFmsRy09H
sMBHczK+D+pnXfVsexxG2DOUVyO5dqfEy6XZ8xHT2ecc7t+9+9ds7iQkkxzMTTd2
zdp589T/TUW0RioodjUXgRvcPNPd7QYQMCXzkxwHz6Y9EtE9Uj4ris4QRir98Tbi
DCejQM9gSF01mYqyRU27s7z8iH4ZkvE2R29j+d1SoLxJaQ869+y3XAaz99GV3h4I
ej2Ve6nM5hzvZmCWBVm3uIMtnCRLr1HD43nZgangeIUvA5Z/FZKVBJb15RZjLWT7
bUMv8Wpz53awe34vpE4yz8BunkNBhNZ6+dK3nNFZHTS8EyQgnBTF6hQkEi7Ujpfm
/7ZWj2c2I+eUtQyg84WKet1xr8VboshbXU70fdYArLD+Vi4ujD1Pq1RHxXhAa+Kv
77/ybVA2vvGM+bHWhs7AKfQG4srRNIpvte8kiCYI4LWOhf15OE906dMDKDxs6+ex
r5ZzXp8qD0F/Rvcvqf80YfdzXMhPxwRXYsY/aMLcsV1TvM4jTdmpaCBgGUcbp4og
/4EQd5rMroUMhGgukj3z6fMrGqOu5gWb84LzOt99S4d04x2GKRil5wJWOeTvTFIB
84fthQqLAyEPvs+MJ+hawtYKVNJLc/8vmW0lLCt3J7gpHs/AkQeENaR7V9UkuVk8
6pCd1/Oe+ZPMG+roUYj4wvI1vskQzkPsaYzw0qjgYqYyCsuEXFn0QvSGQvML4cKG
za4ONuuEJYPX3dL3Rzsmpk8cu9dWmc/ZJeRBzUjfyZgKIJK7ZGaFcl5Uh9sanmpM
S1BcHbKEMWPO7IKnofriqURO8CYqGaW7y6dOXmBJNEiM8WpeqM+jV/99S9Hec48H
bhvpCZy8Ta/qI0VzlTos3V0DGCHKbmKJCcbFkz5BiCsWqgBx5AjRHM8X9cD/9Wxg
I1gH9t86sNGtdThbZ4HcO3zuXGi52jtFMj0E5jx7Kd24xX32Y0Nz/8jqjJSrv9W9
sU6ZAoa2RuuiOBWlMMhjU8juEfVvX1CNn1pV5Vw6D9g1k5atn4pxJFmgmdaegRET
/IHldnfTW78CIDuEn/rHj/TOZMuGp5myMs57+M/hh7qg0Lj3ygqiCQhFaom0+jzA
BT80uYNSad2o6Zer0pOJrcPd1T3/oA0ZZNOYFTTvg0pPMDXMxuuWiO1y/whAjaKg
DZiJRsDPfHSjlqzptrQOUWXLXx/peZaW67HprYVVlSwsPJ5DzK4hE8E+WDW2b6Gg
yEOREZIezL/jv+JHfQ++Jz/FoL9owObhaIAlJZ3z8rcC8YaM8YfhnZTh1llaU2vK
gWNbngr5uQR02f8W18FEAzerxtHw7JwA+RqyaRUuX2AoTYyPyOzBKXstSyseWVGA
CXKfkggvPx4HCSxVgMvJmKR1k49/JWeWCiMHa4nzWsLUPHd6If9G13yU6hVs4kjJ
+GpB/m7allDEF9u8AFrzhG0bbwlVesgiATyC4qA3c9LfClgCHvO4lpaStKJmB1aq
G2wZ16oIr8IjIAbFCdIMUP5myyxXgxWpiRIgAB2+pa+soAvo4yPTCBkoTSwvruOk
lqzkpwSvwi+wYRhU4bLP9600Udpd4JvFoMVfbQ93pz7z4BSGwDddlFg+NdSBuc+f
i7atMEX2F+YUz7FxjUHGIwVwz59IO+qwcxrKBDeUW5GhZmUE2poL2wJ7htdZH1nt
H6PnVYcjhoxzC4GSnSxIR6iByfaJlVzLPJQ2x2Mnx6d+ZjOZJ8hVKQcgLrw2oJ+R
wXlbmpmlXWhka7iJle+XjLMlAsYc7PdBpx3OFE28UdilE0zhBxrB9GF6bfyCmDMj
/hpr8GzADFpEbE/qaIfYEC+ttO6XqbsVuS19rNw/cSLwH06fpQOU5wRVjPJa8EHK
ZOFWA3xRObQZQg7vSbkSX4WB7yl7TAVAQmvqmaOm4vwwG9A0GRjCcibAu0pq4UO1
2jK8TZ968iTY1pq8cU3GiJzGYMe7k0LDMols8/aMmu+nfOYYDEIVPGOYI7gaY9we
jV+lmItGU7DoJzfLEMMzO83CgrgOO+gdVD/TodbBTL0+pgzaRtbW2E8FlAidHLLp
VFyf9GlF7KxTT/JX7XaE9VD9w5m+TaQofP38ji0+omaH1cEsw9d+EZfefszSRAGG
mvvFky8l36m1YaUR5oJYoSGT21UL/KTVL20J+1c89e1H9AtnFU9XZXxCZuz5bEPF
Cy3iKJolyP/XzB19lyGmnZ4SZA+jz4S4gsprY0q5DB4G5Kh6Kb7KV81Vfm4favNA
HQBSzWEruKYKPrMzqGFx6nLZ1QQqXiy7TzOiS6zNlJ/HFdL9mauYamyz8YcigFaT
frAK3wKi72KhDpWdh/2RhSqvBRPfYrzjkcKL7Z15uo4VQ4qE2a/XsArez/bIB4jn
MFaogsVn+XfFvT2PJedgFWTGUS6l/MmjMr96/akrfZ2PEVBcQ6Qe0dmrxeLwjVLe
QkvsyjOg9znyJvNFUiY21MYn7hD6FO2evl4Gw/BeQBi3n95oZd/cCO/s1RglNVZv
Hzws85E5+me10hmXGCIsU0MI+T9X1W99ge5OZ2NnlTFq1ZBJ6Knk4xws0HPf2ysF
4sdcnICIOMdNl3z8PtTFNNvBhWJvHJznHI9gmxCqnRew+/qzwvTHsR84Eje1XCKy
p0c+lk722vc4XpFIt5pzM1jUCWu/4l3yWtruBgsDJkaZEwyKS99/it2hI4n7Xkcq
5ZwnONULjZTXTaaV7xAectghz7Lrfnqf8ULd2kL0UPJtp5zEPIqTpCmBu0hTH2FF
ylFosWcMzTj8hsXrzMZEKE3bU6l2z9w5p8j/qbwpzHPJordDXpBi7gAgQ0RA7vAI
eIN4EXVqaZdC0Pn8Z6gXCTxZHiKxW5oynTlMhZaT146EsjyhBEaWh14lTEhRXE+p
lx0xomMC9GYfV9KqQ+xtQraiSZV3FurK8sT7fb7ce+3WgmC6vzViZ9tvXpP3SKiC
1QRR+C8eV/C33mgA8mRhJfPufsOn7+RJUFQYvkqW/VE6ZiZubbMq58kEcPrcmnl6
OCh0G39GU5jOOr50Cd20cxw6uHuNgUaRQKjqcDgirBUrIRP1HFHTYxdHRwl37yPi
CT20FRWYRUkjssmle4rZXXJ/7PM8ooG8pui06pRV0uqvnwkvEnGsycS6KIQrSqZJ
B/lQwxxC8+1BM9MU8Lc+carDX8Yiae4S9b9aVlCUBsPo2JjA+SG61dHKD/V4ioi7
LgsV3j15+OwqEv3pZ52egHZse2+pfO/nwV5ljEtAoAjenlh9HGmqtoR0+CVCqe8d
lwjdY0FQeDcUYg8N+bRkefudLRr9m5bXytAy2gGhuYkBfvyviFUPixM6/iN5J6e4
TEIMIh8o9hO1wsTpbXKypFxppA+MTzbeWT1B+i4h8vVsevqq9DWahqU57doKpDsQ
QIgC8oZV65YZBOlHLKXj5fa7D8Zu8bkXX7SXfLiqlhEEZwBkj4xJ9LafrIaaHxzL
dcyswYQRyNBEYOM4/7PO/iztW2+Tbt+WZVyoENsBQIgoXkISq+HiCgpjjQvqFmLv
0BOxQmWPS3E6My03Ogwn9whg1cAVH4AKMgCUUEkkQr7yPeGO8SSaWqvg56+Dqith
28GwhThOXJNz/Q+hV3BFrW4IXeFncdHUD9lgeDcDvc/9MsXOmQVm5uWZCNKDxjqR
M8Q1PjH+KxRJmyaFYAlaCdgkJZCND5TyMoF993NVVNebwKi4xIFm9l/fN/jjPc9W
pDuEkokM5oNrfGML8Tfa+Ef0ETzuPyWhLWwSaKcZtk4205ZHpZ3fllpZugl7q8M8
QEYYMvtuCIBZjYXV9T3f9rMnKLyFMf4FyIvApbeIdbBCcndICUqATYSzpT8WN32z
yFuQrzif9AaBs/xpDTbY2QIzoyEhbpI/41GJPE5EFLvx8lrbOU0sQheXcyjvwnny
oRU/Yn7ExhuN6ogNF2fy28bdgtWdn2BeKJcin9GZ+KLX9madNn2hJIEcTbMedHWg
WtPJRDiDeGSKiJaqEotFqEQXbfMDjbe3cj7g2NldmSPw40g/RrO4gQtfGjMf9pTx
dT09rRQiDw5me8KMCvazV0hSf5p0yIrgxS8P9W4k0hIRWFbtzunklEZmJLq79I9m
fR2ynFtsZYA9vrMlks+LcCloqdwoVn5kmm7H6lMD9q9ESnsMiYQkKAtjdBFRXvye
WxMGp7HXF8GK7UPWcrfvNGpbpvIvHGcJXXcktOe6kf4u5i7n2ZIhfi7p2XZBGJwW
yqX/lvKIC63ahA/dPM1gsd73GGIP3kq32pWkdncfwttO6VNA2LDUwPE6d3vgpWvS
urz4XvHZSa/fljjlDmqk2XSwqyqOOGnjhTpcRMvKR8rtRnw3rB11OCpTM7TdJPT4
NmT1sAc/Fswg+98h7B4eV3hbMjUeeVhrq9bVvwtNAY1PNdtY4cqRQgF9n5Kh4V//
3UNPuX0ctW4V7aa8lKkSWbxGOd8dtboOPUFbL84tg/itNOjaUI6E5Sa00HAwOXQn
hZR9ipmhHrhlbwhdsYYKyvvgn0GrAo2+GecVsBQrmJ1oAMu/gFhZ8Y1APnOCdNOp
/QpfvjRPGuqh9QIGFwxiOQ55aSQ/gXETOF7oWPFZOVU=
`pragma protect end_protected
