// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:51 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
LfKPHR2pUCXbuI3bNFJAHn877b4cSI59dwZE/Ewc5grEE02pmApKDR5RTbZkUN3U
OA9YuS/gxyidgqFQMgAPJabaXfiGk7TP/DVjYHUTkog9jMJBihhiMmkwYozLDVlc
IxGh+a/wOvJlHbZe6qKpuCdJTem/yjFTfunp7Hw0F+Q=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5712)
xH9YLno6B9o4YxDhG1aaRDalAJMvPDc1Zg3Ju5/iK8eGxPI87l0PGaggrC4isBmf
9dsToXQ5m753svwf94/wK8FQzEVbYC6rL8cELzbBQJlx5amtJzULj2553kVBClbx
e36BswExAnecHzfANSmveFjGB55XwjK1TPoj27C50gCHR2l+4vNOs4nbHZU/sm0v
+yHAwyEjlhrJXdM718g6k0OPoRxilwYNPFkRPTtRplj7ZP5HKruJM/vax47czcFC
ePJEBwyWeaiih4NkO6JhKAG96g0dQgcfOuKPQpbOsmA6V3FxogzucB8NmLy7U31u
WvPsMpljWn83V4Y/zx+QxBMcifGw4QHRvUEB90QN3fJ8jGiL3xZgOK2PLE7/w3Kk
WgJ5GGJipwhWTIzXwci6YWcx9qgyOM/fezzKdHkmOIv4QEHRqqMWz32902A4Fy7f
7T61IQXX5dhehgufCxAvLdXOy8fKvrT7tZALmow8qu0cCwUO2n7d/SUiLWybFaYc
geMurBD28dQEVErFHWAuI5tcJVqmuwE78FPzmA+YQ1HK0VIOKYcl4kp+tZaExlrM
nwzhD9o++nr6Xv70eE1L+wzWTuFwJtvXadfbVSOHKt0v1VpiIbOA9FMkvFfZJDPW
JjMDvgvsNWdJCpUmNmVVIeGn3H5VrHb0odttyHYaZ2LEa5yghfLgw9npNt3EF9G0
Ht80y4xHVc6XMsdo0kWaEuywd+pelxtttzBVQZttAvC9y80RSASn4HL8SomfzC5m
ArqGHsS+JQ6EF19gyvKnSfhdvVwODuDdsVc1TTABPeONV8DeGcVWGzNvneHW+ods
TDPPhWhAV/Jpjw82X0yX3zTCXvsr1bnScQPierAQaRWkFNYNl6Dfh1MzaDTuIelT
o/C2W0siaCMlSVINsTDs/mNYvakkkpoUuWDdv7WU6Ncr9f4jK1smF4+GZIWz/nd5
RilubFktl0pP8gPPd/W1M+gxI8Vtqj9XirQc5LUUiFtLYCNc7XTC1BVzU7Scm+v8
VIR4JmX6sfKlgQlEL8xocoGfVLaMJtZ+fNAw+J9jSFY3G22NoM1G1Dy15N989jJn
5OAB8emJ2znpVy37jcKWGLxQO5P1BNBqP4FjfJ+AB98ufH54pIvV1Hapkh7AivNw
geHYpkJKr6j557nXf/svCbfYQWtTFGdfkQqT2243SUXHg9bMWlCykfGs0mbfoLPp
cS77hjiTjFEN+FoDS0Ej6L9/I340HfPc+VhgfgzDsZPrq3F8s4T0S9xOnSG9K3Ma
7/FofJ8M1Pz29fih/2qIdpjwWQljcxZ0cJHvIFcVfkKZZHq7U89xNenGujrwiRsN
BGPkC9aOyGOVcDILfgjSiQmB9lMzXnkK+Dpj9h2xKlQDomX9dfd18wp+WuBvB9id
WdEvSp/+hXUETlrG6HoRfMJozgZu2IT0ntHGIe0Ec4/bHwo/nVPNytxJDFOin7sX
hEJ4e7E41Gs8aJWw+Jlh7EqeJdDFf1+3DTqZeBGMG90IW/iEruV7IrQOxN7ZAp7a
VwYh5V1MF546KwIIKtBTQM/T2PKAWQfCq0tvlEV0/pR21aXYiuATvrmHMJtfe5Fm
JxuIddYQ0SFzjUAcQRapi1GkXjB7OnzBh9C3E/x6qqyZYALmrCl+K+nuU9pppQln
aQsAr3xa+w40BXQp6uNuy79iU1+U2m8wSrf8FyxHLs2AXXQD9o9Et9TiC+7Xjdso
gSRzazEoMKk/S52Namw23PmbWYHhukipjbyPkOjEKDuYzK6x22LxCex8zBmiSgvs
N81qGCeokbW90iv8hTmOBnktWCFVOIM5xDCeMFqnKnsgAusfe7kjxqNYyAZVrfCd
Q/RXZaYNY3R+J5RpyGE87T63WY+1iMgpvWlPXkCkJCDEVOWz5UDbIo3kX86iwUge
KRmQvzhjp2Rt7ymgwIS25+aScCwr94MHUauTUWUJZ03lfMK6IkZqg2cLn+Anmmz7
xutG9IOoPfuUlYx/VicBKWlM2LsQS4u1xPqb/8GPy2XxKXURz1viN2HPqooe7Ys2
3z3zT5eE4KXg/EFw0MPqJZL3yLA6qR4HOStfYP11v3SwlMvN+IHl8PM5cTtbjCtk
vXITeM4TRjUVqN8PP/+UlD0f+Et4jprcPUApGZBppmWSTDgO6r+8jCDpTvB6rU0t
gXfDQWgacMXK5MgaAaFFFToBnnG5z39Ytyntbr4ICh7HyOcrZsiHWQzlZebfAHKD
v7mbbE8uBU8na1YRZakBMtTvGCiVg6+QyZKf1qVu3+EUvpL6Jrz228TbahbJBwYV
jZUavl+cMkE13E8iqrq90PNson8kHY5poRl00yYEAaaZXxyP1S7FSggHqExAB+e7
pEm14o5+WX9VmCtAwlpQRm/kcdKHDUsyayiTy/H8/hFFfPZfWFQe2NR4SZ4WX227
BJ4tRGlj5yU609Jb37Pjn1JGqBwBYdsLm1P6Un0bnX10mqhzN+vGDnrvQyzpNlqg
Lkbk8tYViHkfmz0eHcnIVgTSlw43HK0H/Kqr5UqlArSGQm5rIvL1hHS7sUNY9bhr
w/HpOE1jm9Gw63i0AAeeUiMoCgdsMTRssPeGvJ1kQWt3OV4nBXvMA4mM3t4Utn3w
717NSh1/C4HobSEcfvq+3i29dHZLKi0VmeKWSs4c4ZR8EortUk5bYfKYF0OkLWkp
YRhbLwfozzV6OtBawQ7AZIkqUfdynQ2rxuKkUiHGAz6Yll9aZC3GMLuDhf4B8v/3
QLb1FaQb8AtxqxSUkZW76sUy0M9IXx7UswbzcQZ9lgB/Pb3Llhp9QFEzBeK7TmSt
bWnHK7AsSrgNuNFEofbcIdZviNiTHvyNaJEVKOQogAgLEScApDAYBkPInfQFV80i
/iKsFjs6zVhUK9gSXgv+wvbj1b7STzj1dqT00KFPMVF40Why7ut+99QygtsypyQk
E/CwbnUukqV0FSVi6yOkpn05YctmYFANXLgVWvR23kRJgse8M/y5WQxnSX1THBX3
CYewmy5e0fiuknovDSaZfKv1vXGCQ0D6/jzimtyZndoDnmH2kizETTBb73f9G0wa
V5xnKr7HNYv54pAzPUU/2wXtSrjqFP5UDSl4NAYEPYLSSqC1uuxrLrYHvCxqw+Sq
16+Mhptc9HJSU+nMpj1kM5j/9Rs8BsGTqpQm4G/ler1RURmxWhleBCa1We8jdcXs
P8yCXsk3CvefxM3wyukqn41D9qeE2PnDeDveLkhR9ofudzaawMIWBEz2tTI/xOyI
Zgv3maRAx5xySbjr0Bawxt9TNbgqvG4KiP5veUQXEPTrMK8S73QtJ3SCBl/qwM4y
n5yJHTOIVSfqb8sJsBU2vxRu/ZlQ8pBushWG8klUXmFUAsacbm9uSMI8AuhSk6JT
meundWGdXsh1sGc+egffUMWU2NbbhqMmGCNO37M1IK9X/uI3NrHHdXROfF/JSTWM
0zEg9eTgvq4caw2QnytLP28tRm92ifSPl/iA74iQj3dY8bAIw4uBQp8sjo3RaaTl
mIjYb8ozC3YIxYnTgGl4viP3GUoYBF528u2dsrStGfJjOCHs1/RwJdUMu6G22xOA
i7ucP0rbpbAbNf1RXuJvy9GTpyf0dMo083Unvb7HwH4t1JH9H/GBMrniyjTCnUBv
sTvroj/H/og8Vb+QCfFJsYXlilvm+IBK/LiEzhuLdaFi5GNEhlWnOlp7dgmqL9Sl
AHKIHfCtRUco1ttRpTq9pFjP0hF5lOg/BPae7B2gTPRbEuJolIRUQATzwtD32aps
OYV/g+hVLv3wtvSTfs4qt1yacSCGO6Ya1mKh3nNLg18kWEcs3+Whx2MH5J+h61ZW
KEVzEXAeVUO0Edf584idlY3Zgamo0cldwJDVXm81+Hlf/yztZIreO7cEr/tEdJ+W
BKeimOF+axQ41QcSLO7WdQwulO+dX+KUYxeXAF4g28FLYYcZKe42NQ5aoe2p8z8/
+1NXedaprmNXjuV/rn34NFaCPJmn3AZKizS5PF9yhAge4wGSg3nuMm7eNSUCPO5U
UsE2JbybXSYjHUk0IbpR/s8aakZ8uLAMOsGucDKtmN/VElBjbgT6hDlaCK/BEu/W
7ZS842kjZeihoMObzUxxlS6kMcVvwy6FfohSMLx2tB5Fzm+j1JA2RSnLi6MPS1Fj
AEFE+EjktbK4ksVFU5QZs0FI/akQBUW/p2cnAZNJD5KwSun9XtVanDG5DI5FqLo2
bN7P9MIJ03u0TQb/5+C0T23eIIg452a89OG0xhgu1mP06wlzbgA8iqYRTq46FdE3
pRCa4dRsznwjvmywzTh0jFqfFoq/L0WLfn1/A+xJsAUVlM3utgfjLEDx+maoYhOC
FI317iY1E4g03ggWFmuCarulochRglNDePb89fsmvoPbbB5DTdNCWfk1fn+I3m1K
T3YVAyooCXbiNhBC2EDs9uDIsQZEKJH9nr/6j/6cdl6s+ChJRibI6MHC5wi77Fvh
6GYsac4f90EENc/DJPirwQeSkwqpi4Fofna/1MFIAkZ3V24gOXZ+HuiBpB3clHDr
8n1knyWWMc5A5BJ7XkoeYEc/N332xXxTUikv/yLgrCjgsmP2SYG6cWlsAlH/wMYj
vt7E1RIlnvwgLAkmd52tjYIRlhitGlfKfnTveqEnUe3WKctzlc2j8XIa9UDJAZWA
THLT2KWptCMUDNwI9Hf30y/lKUdm9cLJBqPtoclxXgXVcpSXWYX8MebttkhLHOYC
uSL90ufLPhQbSwmcGqgboEsLTCV/prD5Goao7VqmDsxx4DgaH9LQABnuVkZIVpkm
4DKGg9PxQPD67oZK67U9+YT9z4AjI4WAop/bC2p+wWa5tvsWk3qm02UP1sNzGcK7
VgYACE0d09tMU4AZHNjRpvUU8oNop4+TCeFxJmzzFWW6Es97PiIvS/KuOb5JznyR
OB1ZSwJeuJlFoVJtUDdXFzrggkATVukRZJ+Bb6M8AVorcoWDDhuX0/KBZDRWyvxK
6OABApB3ElOmQS1N5iy7H8gSpYb9qW9T+9N6A66jannWyWvVbwz1Nn9vajgw683x
/1CVmSArHXY3/M8e/rEM64Sx2JbjJEpi8TYbVDSi3xKUS2IuaGO0136HAqSuRfhg
w1hnBLl1DR71W8fEO+VYm7plzrKyHWemmPeo+wzVzz/9ezxLoHZdrNMQG+gm/9Wp
0zNBIun933WQKtW+ibxMeVASZgQTUpTp39D/VMgB0jXjA5k2eV4QHTjFndc7jNeE
cGlweZ8qOvK7L1zezCiEg0u+qVC1QjD2OOgaXOt8u1Apb2ljW8UzhkI+KC5rfPhA
kfuIJTPMQtS3U1scUlbKHi3+KjjcoikL/PeVDjsTb8SkRHloH39j1updr9EBy4C5
6HFxAdFtB6iA4isghSKLLjhPfNy2xUFUs2JJDqkMDQmlrEVB/UqhsyLjQgalUvAW
I/5Afpw4iwub6uUKzliqdsdzbSlbk3IEjPZPMukf1AImQllWWBTQHVj2idJ9YAKG
cZWI4+ZEduzaQ0i6jR8koZlVBFg0Oearr73x+fqjqm83kqA6jWgmim5uMIBnF3VT
kvDGXFcQt7lrlu7iUgIAsgAMgAidgl2ISheRuSxi234wtnpjvLn9gwlgsHGGRk6/
gDAJWMx+vrDiPhVdix7uUONnwS705xDxtgVMWZa5QMIS0hoslKCPCyY41UBCLIY0
Y86pro2EWjUC2rh+IfSC01ABXK8RhtHBFVX8jjSC9uuuJWE/ACvdgbL3s5gKgWTs
yCOs1D1/9QrJnBiJnvzAT/8L25Wy4+oKDs2m79DLPLOv2CK5z4Jdm6sSJODmQjn5
jMs3CVaPJdIz+jIFXgp1IGGlCa5kK1o5FWuxKyosWyNQ2b6VdI7RsnvpR4jV5J/b
rsQZA24PPH2ogilwxVl3zxj/f2SVR4lKt0T1l5eSZHLp9Fa3tjTU9+pl2GL2J45K
znMBNn9tc9/kP/YxLm74wSd56L0qtqt7v40t8q1GI83rsxt5VyGkYqHq8mjSA80E
7CF/BMCGiBhSEjtP4/mWxiLzgOvz0ZxILPrSb1gStsG6hm5c1jtiItqj5AHAARcq
X4yK1xG+O/vc+7nTydbzuEq5ivdIR7HyjKhPF1C0Bf14PI/yUPcA+MIFoATb29mk
XX8ZDd59vQJDObyC40R1L56OVnOOFb1rqLmbyhwpHHsDaUIwwnMPI8s9qFvXr/Ee
JJe+4IsKvCXDZn54j6LHmKd7FcGAc8Md425J6lWKOjtgj8BIl2/vqzW4WbAX/ltU
fq8intKouz0d+MCqyi9N5+ZNvrPPXw5LjDTgcSqNu1J/Vb3SwKknRYIARvQG0OPV
UKMPCGRFKFXLLD8kRR4bazo74KpmoTKaXbZLMDXOJ3FnsTcs4ZMdkxQt+tnxi6aJ
vaF/do4PDHeuvc43kMSYMSCMGVKBwCDiakPRtmFWJos/ci1rcKwlTFz3H3E0kkhR
ROdrRYw308+iD+48ixC5f3TqivZ2JeqB1/tTWn/XlkZX62QaYWZOvVQCWd7k/Gkm
Sw2JS8ft7u++VcySPzCRer7BrIvo/rf9KfcnqNgplI2wWYiwQKcFnhC81YtmQEtb
+PRgEWGjSyidMxHNnAcOsVMXH7SBCNQzrMLeAlm3e87HauMfByLxEja89nR/hcRu
l0n2x0rji+JxGs+UG0afgEgmvp1emMr3U4xb99v+OOlko6IUkmu/h6NCThpz7jzV
Xc9YszRkqzZF1Q1oB82onfp7kauJB7IVk2d7IhomzkmZzZ/j2E9UMR/l/XZPeFx5
41HbAKgC7VcW6ZT21Q7spUQj8UfPZPDDYJ4QXOBGLwz5F4MKFkmgXJY3xRue/UdX
CJz6V85OzxVmD1J5yhB0P9MVulL1H0RVmNLLFiaYDPYNNMHqqEjY+vHNlRMc2Wws
OTeW8/uzizynBfCE/8RhanMOgBlp4XXBZISjJx9+IhF1sA87Q9b2+p1h5BWygB/y
9XiXlTLWxrxRDJQl7I7xtqHY0OHeqW/Pj5PpMz1xYLuexSZSKeqgLtBR2OoNjKEr
2Pe1Yr6DsTYlaJmQDuwpoMG4kgBJciWeIPFlaVoR0iLGrfcPuuIhSuy6h2GAEG/l
2aYcmPfVaZtoNs5OkgRJiAGgAVuKqecA0GpwK226Vn1j6Q9exCTQDhsBpuKzSZaX
SueRktWbyHJFkYnWH/bEdof6XObpt2Lejaz1XS4lq400A8XMVDBxdQYF+qsRf+Mh
DHTlSjmapv5pZsswEp+n+ibarW5iFjHiAKs4kRv9fQj2xIsgTxWRNdv5py4Nx1Em
WVXtZmj2rFST0DdoYeNmLR3HwK+Zv77ttsL0BkpJ1lu/NQi3FHAL/pkAfp3xKjrt
yVrLaMgfnb9Fk+pOf/5t6+4+zX7ji3IO8sUAD/oWLuebB94/QwD/OTYAM86gxINe
TwHY7M65CF9iZna7PPwV1UnsjCe8hGN7YBNxRRWmt0RswH6vQibWVdP9kuGf0l1r
730Blc/jvyrmqd1N2wVpb0yI+HSx3YdS8eO64wngA4vhC8Gyh1JIoLxO3NjQRYeN
t1zBpe/zHD7ZQEQ+pcEIbPBocXXOgE/oRp/k52Q3dysCbrBeUGInu4jOLsqmkIGQ
`pragma protect end_protected
