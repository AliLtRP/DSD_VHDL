// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:50 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
R2xost1peNx8G4h6fwEBjgE/3GFNx5GbuD+JPU2tTbAKJmA77GUVT8eFj8Xqn5RI
7H+vNVhEGcoO7XzwdNm4Hul1PnhWYk3FpYDuOGCWUjLQi/7fGzMEwa450vIV1spB
R2hVhU0NaID+7Ow1YnUwoKt0p4iqq22DRdjLs2PCBlQ=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 18368)
IlSvLTB2R+pOWMtXx2FefAGP5ulN3HxqIGX6N7/vD1RA28DGMmD93sXIPdDTotDI
ZGVr3DJlkqFnzxHdu4lnlHIbmFQTpId/nCcSELRMLoh6ZZdrgVpaX0sZccCzgsko
uTIR+Xag+6GiWfZDGzVSJe8iHnsSKPDFcePrtHQPCncyah9hi5/gVOBWYU5s3+Wu
Ti2cV3mOT6g/jnRZjLfrZRDSyHFbKumiuC3CUOLLkrurUEx3au772Wj2RbLD9YaQ
DL7KFS/knpXl2K+DJWgJndcs15YPeeM4/Hy7BvyM4R2c487VtTQD17KtADMUKUUD
wtaRAmd8yogiSodJb/rDXPlD/bDqe6+LFDaL17mYanHaMr/0+QwLIkDKznJGH4/E
jIZnz0uiSDgct7UFlSghojmJ4et5F19E475WNFK9Ug0SD2pUJRJMh9RB1mAYGZJx
l/DKx6hP2U4qibfKPqNlrrRQcTgQKS1WTInnOu0aN6QhCXeToMoRH29hK6GcQ3XP
b85nAFab12Fpv8+m32IGSRO2CMYQqGORcprE36Koj2c8F/rZi8BZ+4dfHq2zHtQX
n38tQ2a107KQD07CRJNkdo+2oaHeZsr/0LkK9k8qcEH9p3r1eX6MFyErgHakAst4
XAht4k6QF53Lbyh3LzHGNpsGjGcJCfFHn7YdyA6ROAuf4hfftTqHc5MY2y1skW5v
z7kk4iZgPXbHjdkenIQ05VUbOyz7Prf0nXvDuWkQkcDhqPpp/0xKwwNRHG8HKuXm
F2v+9igvv+u9fv1cKk90A5zRfteMBZhhFs83AsCGOZvcGXuhcFug7ZbJAWzpmyVC
sZn1GQfAdgOd8z/P2DX8X/liPy3srvqbpl5fS/JphZrpMVLicYltXsyTlBPf31P9
W0wpgAhINGwUYxDMjRDnp3rerIOGurpgtKQ/zyIwr0bzzceX2WGfNIWswyi63OLB
ocjQxHGmxHPh00qwMvrl8XeULJw6UnmjEh1Ss3ZzRny6LIWR5KwsYmot21Ed8nRP
+P5laUwQEp0+bE7N+/eRnzlFO+cZ7bOFFYt9lyK57E+zOQHohd/IhitqHrNHokux
sSr4mYYXypF1qTPxr/qRd9GrtuWvmja6Zc/sGk/WSt9wL1yKAs1JjWWNC7m8EgnR
KuTkrx6mrHstChI/gl05Du/RZdYveWiBmsR9MXM3dy6XsIRcCwSiD+7bk0eW6vtq
rqKdDfEE5aBDjuljcg/st7CbgJk42HJQ0lPvrHoqi/zZfPNv84lGVeAdSZ0rmmgQ
0amF/5+WkivKue2+boVpxtRTeWCPcbGuJX6ivxSPkACGekEzRM589qKq59clzjvQ
oeVophVoZI1NGG9ubanqGVy6jyfeYVC0VRt5NRR7pUwnIWPQblPZw3wmO1UVbRrE
SgDw8SC5hgeTGHhhIVZlwo3O+RjR6hAUJy+BYGpn8k55xl5M3bpg++H0bWYM9ypQ
uHzrHg7k8CzEtszLYkkGBL1mR6VXERXCLbZS3ks0lQFrtdVNSOzj0NRoMvMN9QDu
pIJ0ZLH6zRf6NSkc1OFXePLO+6GLIP4GGtbOWB5geGtnUgVp6FWCDW+lk6nWlXpu
pY15gsC4yfjQyyMzp/C7t3XzzSSV4yqK/5wwi83njY2VpHZRC7yUtQ3ja4JiHA81
Vl+DJ/+xoV08GamARy0ibJFOugN8R0zKPBH3bb6S7gzacmfMnE9cbg3xXqmFWYP7
qV6KUzoTqkPV51T75Lh0fqdjnP/IIfN6BmyCA7d5ldAL53htcnEFUYA1LukOxYXK
m+kbW7BaSfQ35RQ2wm45Rr6fdKg3YwaE3ez4GUmuYegmH8RgzsgoNbOJCIEMt12F
H57EIcpooqwHyIKVv6ZauTFOWpv3J3nkT3FPum8DsotUkoA+YI5ANUzFj8lfyASK
AEOOqm30ACGSdekC4kJpwAeJ39kjwjtgX0pohWN43nI0I0zdORMJF1vvs5yJASuq
gTB84QoP1eshXrD5RY9rNTgfbDlbIDazQj9FDzfwD2wSRY5kyaoSF+GTHYu1XavC
52hX2ox5Nasisjin9xkQROrnHsE7tIu3Z0xXbdG/UHqp6h3VGH+XedP7ugZf00k/
cO+3hllLxAxJNsKI7fKKXVjwba8E7zeXEzcVlIIMJx8jdekye1f7PMGKE+YQL8Rn
gKLiJtiUFW9lXDanBHLL0XctZDLrpd3O+FPcdJb/L2PGIbBDUNE6mJvD8NNd/Fln
lca+rSPQsZtgm7gH6OcdiMh6u8jQssNZanGvevuq41j29Mw84XU/bsrnnwU3gE1v
Odo1ZB3mJY2divPFtZBAwzwegt16XYqe2vhvdLtS5IiqkrubV4mAKcMjAhuL3MQ7
2xn9O4r5loEYnWzmiXHmzMAAQ9FitUX8C5OnXg6uEi+wOSH8t6HKEAiRsBpw1b7m
RZ5RHzG3WHI07A7qhcDFJKbGX+kAT8ipitkBWfFLUMxwPF/7xnoWOsMlHF6Qgzh0
nis7xfwv9eCzRFO+Zqn7NybygnYwWjLAcKWfj7HNMxxMDVfCUG+s9UIkXclZPnyd
XXk9aVii8WfxO8i4xNbenKqHqVbEL4j/tBMi4YgtbQmQ0AmaUKUztQaJCE0cB+Jh
C2A91Z7L4s7BaJZADi7qP56hE5POICPFCkAYUIjbX+2+NQdVBmTgiu0UugSstfD1
yFl2TK1E2tVZHMJ35OhOJr1p7M/R5L7dtWNUasw1CwTJHzv09wdZasAq0DVVpYRR
MiLV4Xk9KVdHSCaOTqo5UOO36wJmciuGQa31DNuUUDoxfVtlDRCYnc7Il8YOdhff
ENyiRfPqxu3ee+MReCsq2w4lUwZib9Y2y/qnMast0FoAUtk307K2cHp8wVs/YmiP
JLv59GJpMH+6p/hSD1zuTz6vxLWW0ZXz1QCbMFWs+24/cBoh981DW9RFQ/VKv36l
y7g8lG7EDDfLakB6Fwo1CvafJzvgdgTmbGhfJHlJl4oIiOsJzKi4q9KYGINagm2Y
BjOGRO4oa3/N4WdWy3bAdPUl+Xd1fVNyUOJ3BnLsYEYQLBWhjAUOxvuMZPobozY+
mzJVmDagdxZ9NSJlxwR/e5YGF7b6o4nRrACIKQMAM044FCk4JaL+w1Jtc1F2/bqL
3jYWKsQu3lmfcDG9mL32R95M9DE3s2GIONnGvQQ+4R1DA1JT2Oj/SdzVRYHuDL4g
Cf1N6Vitcs6XcwcQpf7dakHpkjGgnUbADOJQZ3OsRya4Op1lZayM720Un4tWpwd1
SRELv47EcrlJvOL0UC7ayvbwW6+c4h7vFMlceyxBKssGKglfisNB71NlSyPMoakM
xnEpz3NDUcT6iK18Wcgr6yOUg5OhClkmiq+hUYZJOiULkNL8nHwlbY4rd488iBUl
q7hWiXY77safdpe3p/Hrp0R3VZN75M9z9q+ZvFqYq21dDt5USOCEqDwIOQd3s7iR
8tPFfNYzvxIZcfK+hq+Ol6T99W5gRbHnihsZmMxG0gRmZ0bnmjmP3Tr0d8ndgtF8
fklR4Y9iYPiPx/Py5VYo75qIqub8OSJV+q9hunhADU7WX6k87BDfBkjCo4KWxnMJ
l7cJhrXiYy2WPCbbP2eETSJIUg57hdGuQlHVjKVWjtyd9CoSsQAxhKFU5wWDa7gN
43RKEVl/QOcRaUeYS56KF7yJQ+HeG4OYrBAUg3ZCB3EG1orrCB3gBkQnL2Szcs2q
fnODzpXeM7KztF7vORfN4ml3BviEed7XhtumpWXL/rUunLD1clOnIrOVxc8GBFrS
Fd6e/1RvhYLUZf0bHLerL/LiXTp/RbVzYLsNfAfnBsgzTJWJ+NMyBEGAUCpy2GHD
6Da6Vmzxj3JWAoMx0qYVdza77rbKAYQtvTNVfBZuaT5NMU4+a9pRZ3dA1M1zvQJl
W1RO0zv5sIE4jOSgB+XGFx4kFM+CeFsdZ7+tsFX2XKeKfbYVFEpghJVFBDcKfHP0
ShNV1itjGfMxthUIIA6CpRle5Q0qwAmQ4QZ6xKeJGzCNeV7Ml6qqzQWbpPu+If36
3MjX1kKX2Zjhld1Pis7mXtK4P/5Z32aDP4gt92uvUwy1S0UB/RYuq8L8zpN8ljuc
BEx3P0HtSFeeyJIKSiTkKcA9wzn+OR7joPVIy6n+ic0adKIXHBGhuS33m/brJ4QJ
QrABfy/0b2PMMKnTF0wqJrIcw57LqDCTOqWSwaHRDTZrb+e8aVKuWMlqFc8s8ZC0
cOh8Yx+IQoYfc0TdeKmh+KN+h/I6cB1P+tzThQooigO+p5HmoVBNWRahh5UMMWJu
UNU/PYmTnnJ0LR3rl4hM1WNr42+BQ2nlZXBuPmHW52Jqu3THN8lj6U4ogrgy9KEE
9gNFxa6oP9c5OU6jN7laktHAm5ne4es7D0fCJA7dHHJOTS4Dy9Sm4O/AfSuCqkQ4
X3lSf2qVGHCe6fImMSe/PTvEG88n59qKji1xe2qpQeZLAlBlQr4ZP4R3vfoLas4f
oJnqsPM6YfrFQuWGQQYt4hXmaIyyfS/A3r+Qxg0OxezRdY2HgFAI6QczZvvVo1Z5
KAoBTEYgmehn6c+0RlFPAqwDEyQ0mpulJd7BGwX7yyOxdiqntv3FfSPHXYGWhS6n
NsJoaJMiCZO3/ezlotYTapDNWLCMQyMp9RHFAFdFHIZKi3RgYkX8VIvdCaM+4M6t
jyQsvILusO+5l/8jWX+tz/TMwhPqlh5wMjjpfJx6S/JuRkp4x77yzwuNGczf84ia
rfMLSUd/gTjp3VIHzYD+lEa0Gbd53wmu/80o6+cOROdExZNJQph0BtXJZVZVPywt
hEJscsxpDENTBACayun0ZF45r9YJHEru2qlm66nEwtNduZ9ZxALZ71NtMz9sh/N6
tgxvww7T/oQLHTpoZl6NI0E8NJKVDXfVkpX1laOJvpyrowhSqsM0F9xBPdvkyXH+
1CrMMWwCVpImeKGs6Hdl7uqBYjWZvQCLbPRgkVG0k/TqXHcJP7pbjiKC2ALCyJgo
9A420DCUletksjx0BCLBrT/fYJNjCIpKYeUbPYT0D7zp04fA529X57LQzHiK2EL7
MMMAIgy1NTy/++hKuIpBSJClbG/by0oJN6wCghsCDq7YSOdkdShZHEsi6h5XyYk3
pH1tIOZuULluiLgamwRH26Tko7xCPuctmR2kTkiQrItOmEZHD+P1QpdsQ2RDAQlv
37/wntUcBdu2OSD3MlgtUmm/9fnXc1DNNTr33o3shay0CjHnpnOsgiVEMvVrVaOh
5TbXNpIXdXBCGMXKBo3S4/40qhjzg+1Hu0S+MK5LwCyC+8wXrCaoUlS1Mpo3SGMC
1FTXF093/kvY0ItSQMNsR5FuZm0WHUbIHxhdSVssen5pfUj+zKfsJcukQQNoorJz
HZKSnQs8Ah4Q0kO+I00HGCJs1tYcpGO94QcekheN04Yq1Qx9JFO5qxYm6bC/e/DF
qoc2cmQEd70jMppKEyJ2p366++/1RUk0oyiAW5YELjee9r3kdwABiiMm/f0qBwEa
cc30PKvge7oXtYfxydUUGaDTwRuUBQ8UAl9cAPdPD2VAGoLW2phObMA29Cew+YUN
ySHufdgAkmzHUkZaPPF6t6CZM37uDWGYcsw081wAHdywyqDqxtRs5YniFrsP8BWY
IEmZBpTwlnhFZJkK8/zyLW1Cz78e7jmKu9DE4MgIf4gZ0h/NCoDs+EsudamKkyun
5j1TrfdZgERQhFcVHdE7YNQn3AX+cMtyVBxkSTpXF9E5Wg18sDdsEpnEG8ueo5R6
thTqMdn+KW9DjCyhXj7mEEwyUcZrBVKtdrcEfixyUnIAaDshyFnDh4QKvE6xs9lJ
Rwz8qa2Az5mlmyDF8VyDMW884xByBsTwTmvekLn3/oIenBfZzGEmYk+p3cK3Tc25
uJ03h40e8ejOM9P2FRnpZ8QcVDd4dBO8Ojf/jbeoUtvNLRPnMVHUcZ2Z0PPxtyfr
0apH+crRF5Veb7z8iXQ+jeB7/Ck63TFia39gi7jOcSYus+KFWyXZYTwn/Nuw+jQu
x6YpTKsl7oio6eAeCrbhh5ocUctm2g0drSzsgYgGH84Zs/QkAuohgS3/hYuAIsKw
Ayl1tVEBXBD/yCHv9vt1RMHtKEFrI/JQjDyOsJotZUNA7/xnmdpx4ceoAPbf9xg3
J9YYCSb6CO4QCAFENZoSNqqdfNtK29E/wJQ6mDJd/YeXsqvg/0lQOQyynP53dTtl
lE9gVHyK6m/uvjn7ZYdVumT3d8y4bXvVhCbWW2bThiX/IAo6Ptc9KaZgCexoz6LH
ebsNISVK95KY0NMCMdONFegz1BZHnepz7s2PIST7ssq1lOEOPWgdWTSK8iJVR867
idtTZLUsXOrgmV7SLowo6rlq0uZO8Dap1XgXuyRNDVnZYm+V6e2OIejBdZMgOacK
Ebbh0Qf7j9YrVPELiHHEtKUeXkN9WkayzkZkgCbwsJPk79KjFeSr9EoHlVTcJiLU
rTU6+o1GK/sgxxaXVZTfEVA59RS1LwpAolf7KyoPYGSwiqeJHhxpKp+cAxDlG4V9
I62HqGC2tX0xfGe1xRATYG1OpfTou+7O7M+pmsWgTzaCawr3lzz7aIbKDLGHZt0n
aD3tX2uXiSdfHrLHOfghe0OFM/Xpd48ggpyrZQU7FuODcVHgu6yphriE+S/ytacf
QfdpnLSJnGU2Ge1i5v2kJkBpCxqHw2JAUS3kBOAbgb3Qf9RLo/9zzCFBwhJJ1Hdw
VVfUO50L0xm7qk9+CFRO16ga8J47OYjfolLdtmR97ZeFssOCVVlrwM64+lBjaGbL
8DdtqmxFYvF+tBQmvVuFlFdAynUzAd3r3vygP+Ijpok5r8jOzm3ecaXBlp3kAAPN
AKq27fIGdNtV8TLsEnkm+cFgVPa/puL7n8GIAR9U2U82DMLVb2R7N5txvOMDTZGk
Z1cPjjdKgxLtA8tgvJni1CvbpPAqnZOk3m19CUZsvwr/Hz+WRlNvYLbMd6WTm1pR
pa+bIptQTxFIMYmt93Wh/nXRE4ZkIn+ye24qLZ+lC3vgh2Ablf2xD2DRawt8zri6
xjZK172Np769rK6IMahrnPTv3vVomfGOoSyM984R0VFlsXg08EvZrwIvlGDUoyE2
FRivUDBsAtirHoCGI/NWk0FA9UihD4zldoK8a/pRKIPqCGTBrS6aEuj51JYqfF4N
z1iipbT4a0r4GfCulCKC9Lb90BdM7lmBdCqq8sFzPXyQQKjuhUEl4Q4oT4ZDLYaU
v10gZxzGJfw06M8wbFhanQiToh+ilZ0Y4uRUUrnXrpfWZNVMPlfkZSFIZUi0qQea
6bTEiIF2NtGDKyCsH7D8Hr4AqzUllrP4XLFVGnUQ4yJ/TnxJYwklI30Ve7uGTPt7
LdLu22/9wxkfwDDdT1z4mV0ovYzDHbbL+Ny2EFBMLELku/pBmvYhbP3Z709STpi3
J8pFm11t3w8zBWnck4HtUse/Y/BZj/tP/ZtxiWZDk1K4f+fgQzcelnp/nSxm/sE5
a194dG0ik5XyEYo4nRdaQHA6IbUZdy9YvvxY9o2sf8imSCfL9Asel/O9DcM5gOo8
FD2tK7fw0CgUS2hDSXGbsKwOBPrXXBMXeXcf9vANTjyjoCoD5zxTk/Wd3EqWNsub
dc+LQX8MwdfSpA5GqdxeZiXrR4Ea0rKiEcJlEkgmh84RU+Eh8TXvgowp96fe37bq
BrTMV7yzhhAcgn0/F+bfn5gSbmPMoYMfzGcdDsEmkVq1sO6JT1SNvCjYhXrfev8J
NDqwnbwAcnWXeYGrUkFTLhMA88O3gLNvbtTRBGoybZk0KzOGRP22b4f+c4vAjCY3
cmtPmo7XmqjhYdV2nGPbQzve7XgjdMFecBxNxqEPyH53PiM1C/xRhSYaVn7dxHOH
nCSg/5Bhp7CCKib30MKiZSFUppEUFOCIjzq3GF3S9lFXAJyMn+Oej0J/u8PXtPwa
eZOUhq7hOdIEFtkUUrHYcdzTjqBOVn6sgzCedVo9hE5Oada9/az65oijXaaYr9bM
ecE68/AhTiIF5aXQQORDBRvITsy+ZM850oUDDUPoIoUhjkAaGiKNE3HPB5QH097i
aYOIJjEuvbZVQRACZsJv6E6OxTVkHpX6z1DG2wkAkL3GF67N59SA4ncYSVY2Jbaf
/tter/Y0odrqvv2DFcWcMT7KRP8xsK/SU+yCBJbnhxO3lkDu/H+QzZzxPPv6N/dZ
VvCKjJVGpXGyuxUG8YKPv3oXlhfO+wW8X/LMGIrTHcQUlvnW/7AwGp0cZbny5twD
GPXhK0PTr8FEejxK7zgRHPrwKYOxmYZX2L+VMtZ7p90A0nlQkgai64LUUis7XsYo
SYsHrqPJePxCWR09S1E8xV0hWr5W7saOtOoTQRyqWob9kgkAg7wYSN2FKW1dGYol
F8duGbE+6GO00ifkBzi1WRfYDvpYulAE53dpmwykJRb8NMq3XHxjPkP+A9X2tc0g
e/HbsM13ZGaEE5cyvlKbX6hL00czJKKRZL+8b7D8/9h4ts9OgjZ+FUWaw7jNyvcd
k15k8FNVNY4o15QIiZ5k7zYohG/YbUDOdQslqN1A8XpCzKgOWdVjueGrSI/mv8db
iuuxgfG8IxC1pzZPdSTXxiaQVjMLA2chJYQs0dQYq7SnXAKvSQqOOYnsejkd9wJy
VODfNEA0uuWoGqP6uN8GCWYFBZdkijTEsys3hlJWazmujcaICN1DHOI+s2uNTDQq
R+j3kSd1agOO7mv60FB4dqOinq+DOf7Kl6c20cAohc7SJLBxrWv0a52bSbXO1Jfo
HFgYHzBL7S6y+JXjjhM1xEUdq8Rkg+5/02I3S4vdbdUi9BVvENaKPcvoS+KwzQMQ
JdW9oQ0GVzcklaOr0hwSk8Yyi5Ck82Q35C4vXAMeCwlFHBWkpwYpEV0YWFNnVgbI
80Ra0scjQKzc5071yPdTdf2010Xox9TsuylvHdo2OAEaytybnshQL5qy2N92v0UR
BTnWNNiJAIjRW/TEoSsalocLs38RxIxzn0o/Gov6b6meycUW+rZ1HKf/a8Jsa9+1
MndIhcCkFcIz51rXhgZvADpnWrk5hPE+XGRlIpkVmxJwlE3smlY5IOitx5aHGQb5
kVF2FXF4ATwodulhn4xSLptp0SqNnM1wWnv7VLqi4cK6zzrKsjanVfyjpsG+U063
El1FKKpNeDDo0rAisbp95cs6GBD2QHuwNG9fCtdyRnggcDZI8jYGf20wr9zMKOgd
bexdFxx3y58refou3pABftWMxDS9P9L0aFtqjiNoRy1lLDU+RV131Gtzpx0RAGsa
Autb35wlEujMYH92UVgcVRPAgt2gZ/SIHETAJEU9pXvCmBqeAtorf2u6bAld8CC1
103DOfGDBJfdZhKw9/EFnc64ZgZ+3fxLClzaW/unMDuzqdfzWhj76R7gdmzy7a/l
gqPhN3UG++DfT/rieygV7G3fLVIZqYSRl0NRYag7gwR49ichBdJ+nF6pgpFSiCT8
HDFs2pErZbJ2sJYVezfgCKRNpzx2/oLbq1Smw30VsecSCrLIZZs2xXtAjXuInvCa
2L7bQEYYqe1Gao5BqOOyAOQyNuyXpk0HvFGjmHZHwgfSSgoSPM5c5Ab+Zqsd5xaz
F0eXeyCMkyYMhi6JYmSKV0r8qL+X1KnPYmUmaoRaO6+RnyXNYo3d5i38Bt4OV6iv
EK9dGbnPbcg7s3w+qgy6yLo7d0t4gCPR/i/J7kiXMsbpURFoAd+Vyhfzj45Fcxz8
G0saYSay4/zg5Xk0CEuvwy/vPXQvsN9uHNajHpDmH9UfdXYsTNo36a7cthwHliBH
2Lw3vtkY/yOLIHEKa1OTQXqeGHOQZgpeyul+IfqCJMXbQj8oysvhp9DxuiJbj3NT
LWgEh0vej925dlCLRkvBarN02kP3mMI6c0Br5OdQvOXzI7z1Cenl9lbME/rnIlWR
hqPz0Jj7IF8/89P70rW8FRg2FBmVbkfh3lfC76ZiXJ2GMEVGB7fB745DnTphPiKb
3so7V3kwxAglBQWOXtj2Cas5HC6UE5wBusbfDkZROZilJUa8bNc4Sw8wZ+/AuQfv
3JicOVHES03ejYCDlw063eZOJ6tDhiHGvPe9rAkfePn8T6xBUk8XHdx67ZWurrOd
ftgTFgJ8mTnCuvKjJqJokBjQHXanyJZoZqQ542d3FGmp5rHCPM1L7aEonHaPQFhp
ixxzUMbpeyJUgd0grrD2qMavrlKQGsJgtkqmHG0GKxhiBrooWnpoRbgquvylASi0
RNu+dC0/uLC9201pexRFr/6Z46Ug6JlR7+POon8Z+rIkMzVi5vK0wUMXbYa9xyoe
D6q2ZN2R/+cXo7mS2+dGOPVvr4Kc7V5J33IbCTXevghNmAK/1dDgg5kbsFwhClGz
XxfaiVsGTX3Wbn+pH8bU0B0xp1eBqi2KtHCwEqutokt6bX2FuXEgiyP4K3WgYz3I
CybxGFHOlklsROiWAokIk6dkhajBiqHjnvhCQnEgokcmct1uNv/YBZZL4PV/zyjH
S5jMtFCC+fYz3MeI7ClqwPGnuoukbAe+rjGQJnn80NvEQDWXLvhwW44rQc75iWxI
elswNgtSjnbRYKK9tdMtLWUiUodMonaImsrfyUWNJqasWlgZsZN05nSbvSNg4p23
sSYUtQ31PU+DSIGP+6kX3bbZqRo9eeJcYZodNyt9AyAAgBcTkk1G84FwYFWgWo+I
cy3rk/fruL4grlyC2XvIgqNxwNG7WwQS+w1rz8Gi9hiK6ApDpBnlpOeDmpTGxN7W
3kW4SKM5yal3Wb+n85txuCZxen9CzhSg2PxwYeuyOxe0r9SqKz1Th5wdNuuKxX4M
5NUwoEs6p7ZNzUQUM1HHqqoDTIgvIKW2eyA+5X2ZhRwSNTtU3N+03iukUX1+A/8+
Apmd0jbYfJqElnfKVtD3gZChxpHsVF8Ley9b51fgZQoT3P1+RMEtpJosl/CLEpWd
nbg97hqIVSvhEJzEx4K+cFVcFN6jVHgP5FKib3MXvKTerOgPIrStsoxPoY8y+3xy
ftrHXCPK/pjslHLxO2L7JWTY1dvHsSPAcMIxE55gQmcTREtezZseTX8iOtiX/2pW
nxnV43Pm1jRXkfJ2xrc99U5zQZdxY046o8ke15LoyFmDIG8TfNqAtz8qT8Sp5xy4
+g5EKalv7725HhGVWrKrm3jG2udgPDrkFSxK5P/KKOfIwbqQVvfXsQaxWZRhXG9o
rI6sCdGRi6cPikUAk0hoZFgcVZusUKLHwsg106vUhzkJ0IHUF+5wSSuzjZbYFTa6
TZRV5yf2Nd/Ius32d/4EbUrx3rsewKkAOCXNHzqNFsSWAzovwIQJ20P6cwvDRNZZ
XTB8BW9KeZ+Gb2lEl6IN94qnYk/tVTELtc3btbu3ZlYJQM8aCfZbYrun0GRFGe5i
ZPm7ZUtOuPERnERHMC1cHfMInnqEJSVTR6gctRyknxPb9RyJ4vQouHGQCchMZUuQ
5QPutgUuXgVkEpr6GC9+nNFwgSyOOYVJmacqd7BGNUqRwhhroZUjdXSQx822hlkQ
UCGNGrL6fI+XZtPbiGWbpfzDFvnWf4cdwXzW1beGMDI7W5/+sWDIepxfpcZXKr4o
fDaimPwfoSta8C1gf52uEMUil997+3wwpfLmIMLhky7hJ7YTujwQZNkyoEj+UrR4
pySyQEE1jVsGTuEgutTuw61qXd5l3BP39gf94EeytnURIfJs+O9fuc+Cpb0shSQp
iGPxFS5OhFuX3qdOnCn/fOZDgTdlxzE7I4yHMIvU3kBMKYKbb/wLE9D771H4jGEC
anKYYOtg62QNGlbGDucmcaGSjeObvq2qUf/24wyhql5x5tHeGpE1HUbiBF2ZB2jo
Jy2sS2nKH0Hg+oaOJYyGDNqAIpTG70LvgKpbPZpGC6dR95oEnq32vziAGwWNnVoQ
mYtMw3lkA2Ra/updKMwTgGa9/OxjchAkYLUUxJPkYUVnxl+b/vzVZGRlHMuBQzCS
GHVxuKnWZG7Tvft7S9TbvO66Rr444gilHI6eBtzp1h5NJtZx81Evj+p9FHXEFE9u
27yii5Un6QB8Jeyfa6oY/kjLsWimSSqaJB2N3cbKOvGkU8JZTzstOlsEnrlAKgmk
wcuQGqjAuHrOILGmYshB3gzXcKng7spUogFs2R+eRKqweMTZSkrEUdyX/PPLaua7
7UqY2XlnC/ob4pnzvVxYya2HMOAm/bT1luybthBB2SGYKJM/PXjN3lXL7cPKHKGq
cboKDxYMQyqX4hLbbWC+hkjork6PHoBV6tg3kokRh2wraFjLZJpKMjQQOLDFbrIu
xLO3I/s+dkaIKkOzCTLgvEpOAdkmXMxcbf9ctjwD/btklAC2nFExZ21ANTovQ0Fy
N6J7gN3M4Fpqaj/mq8xZqONDx9cV3XkUwiXb85kfx/aFX+ZqyPT/pOWG7niQ4tfU
HAC2+R9sR1fNvxHI7JY3oprdtokqUPQeSbzvCJ4gSsUP3IUp8b1IHlFlPiql7Qb3
c9q59CHbCrmuIhME0DWZhW+VUoYFkUDriwrGaamuqoNXVGHS9v9v+5yYY4nh1jvc
NZNYmXr1Ont/CfqaF1Vwg36Whdv4aTQu5Qd3d5XI5K0UcenLSGfYeDfAKswBDtkw
TibG2IUMHnNaAbC0UmI/kftZ1f5AryArPIgLVoRWHdZSi3eYCTyigqztzxDzLURC
ecXidfRRRPV9zM3pmIZ45eGjRYfLlxWVSSGl2Bc+izecpq/Ixof0+e6zzmUlPgpl
O4xl5svG4WOC+eg5d7eu5ryJ0Pt/AgpXWLs8hU9ul675TI9DHvG132X4RzLyPV0+
r4HMUDVpFmw3MNutt49vwRn9xdSlSbh0cfH7Nbklawl/zkF2GzmfPm1CyHP/SEEc
MJChQmOYt7JZG5fojGgjjO1nOoBn9vAaXBrRn2mOPKxxkJqA58ASqfiv7YXP0Rkb
8o5968ZGExvgPwqbjZjssopcGvyPvsOVlo/SEMMK8olvQUJCgaqW/8OVfe2Hp+0D
CgrlMA5nItVGQNerepfD5AC7vr5Ypt4xShZ2YKBazNWrCYtflzeIdDMSkZuLn/AO
CNpQEuFBsUVMi5YoEBqNN42sbUSW5jgmbct87MOnxN4TkPHzObQFKLXLTZKhwcpW
4imKOWtzOkowL4QZ4lwNKyhgSrpETSlYhHwQRdad8496CoFp4dadpTv9VhdNpaSp
TybGebTQ0HGNFAMbyMdmAUSAqRFfnIRwdW06mG4NLe0dV3aWW0zFG5wTGNCp4NtJ
NJCK+7VlYQK97Q5rLT9OvOEBb5j3t+P2Lf6eY9FsGuX3Y7uDtmPL+ccaUevJAEEd
P32uyxAxo9qgNhaznvELDp07kUqXkSF85yl0SRxGA1eQXGpRo2HD+J+Or1ggzpY0
yIO0o/U3/1Hy+5WEm/OmX59RoO/MaRcV+UFmNBPU3ZzLRVQ7NZErBS8JEBTvJy+r
wq24FQ3TKnmcEKkOp+GlMIIHeDfRaziuCxdsFlZCoBqTUm7g1v0FWiAuNByJ62S9
3+taMe1xCX2BtuNvbglnbL8tjNYgP/rAZRRUck14KLtQpoG1pw0DcpJEIewnDXiA
u/FZk/j/PvL5NO2gZDZNJMkpmlXdmyF9R0WqUdoduhsdyXdaNm9fQkKPhaHHEQvC
ZozdfwMyy5cSCD6nxa4NKtRmR7IJb3RdE9Fk0VjGQyfiprYQg+svA8b/B3CNLyUG
2DyjtkjkRxhxT0hFXssJ/rzBI1DMXjNf9hCrjkyHq6VWSz1p5xmtFkZtFPKaxdWE
Bn+2r+IaW7tZtdB/kyPGlP8Q8NSpniygVNm2jMlpZCRMFlCI4pVeAwS9sbiVd2sB
KDkIv8UYnZZ509Itc0AM+h870Wxaqqb+KxdIu2ej2h9Uhr2bxfwx1im2OcTg1owA
9BLUHcZiOCLaQ7Q7+BHx/+++Lj1gAGG2u5RvG4kYcjHEIZ88eMdcLNsNqV8dqbtZ
o5ku4Cih1IiwRLhhEtQ1Nd53JvAU0yNdwAp5At80CsLkV5nCWkcu0rc8odh3WHtg
q5RSiA+RICT8xaJUQVmNHTSFymJj74PNMtS35yj0dMCswEhKN6sd64l22VPZC4IK
9bvM2Lxe5WWLPIzYMxeJ/nSa3/KK185RE0DUGx8l+OJQ6xTVFilPGUqKZtxba2zk
z8irrpUh9LcEhLKlywTFThk9hNEKmqLYcGL9AQQchwG9KeH6mNltk/Bx16fyNiCh
H/gjvSFPYBF0FapcEaMONace5BNiOjyXo8vz0ZtrujLvr285jaNWSiE0RTtMFdPM
ZOkosvBUFU/OvhDOh41R6oslydP4hkHGENKfGdOfTKZwTvc2O8rdyY8/tubt+eNR
eMzhDyMuXAUekAM5/GhUoU0OZhUeLhrEbAajDc9lrY1TIORMnSBL9A9tSPXtCuyf
lupPbO7Bdl1mK8BrfbNuTG+vnn/ffiY2gkYr4QuTJGK5Yt2MPgD2JuVw8cW9oHuN
HrezjKeQfTkI7qyUsrS+JpDTlMZCOdqY1FEdnPZFacV+RQU9+saEqSCEsK/89SJn
JA9wibDS6KiJNZCuIrDfo1+tGTiTsAjhxIpQwf/o8/coTolNl/2nBoNiT12FFlIB
cOhNm+r9pWuY+2zKRh7CfnAhE0iDwwpGIIPU8VkTTy5ES8AiCFU4SCFodeLv1w2D
3R+/agU+ceOrWykG9to15JwtKezwCufNByyn/CLSVE4lVb6eLSLfTwQqHDllSt5Y
TameTUQZTAZSmgd2PguhJvWG5j4mlZLqTjEhGTPai/+oEjSCbtjkMZ/Cift/HGCf
uJh1fg1IJJ3K2Xs2yYDapplLR+wQXjorXfZ3SUD2st0WcTxVAHBbyF4Xh9eNW0Zw
O6tSqdtBPUTASzLDUPoUwpPKpXBatfl5x4X7M1IDhzByq4OQzwqXXHNNv5iVto4T
yKKGDRIMscWxai7ynrbTlojDVU/EhXug8tdd6UzJvujqiGjoPucv94jKr4QB012u
9NPD6bCTPui8K5OMS+bBbnERrzlgy0vQZUrUA43wpM0Qx0vTnTf54h+XuifJ7I6G
SmjtXtDtz9syMcAXe+TJ+EbDHNlX5B/bGvb+NdmDqK0e8U65bC5QA/bSd1GGM2f4
bJ4EJASAQwQlt+RAmA9oIulE3OAktIzhCwn3ZBenwxSQ+PAetse9BakbnMpAO6+s
MTB102SBulLigWSSyPAQdJ0O3JK4wJqvNn0qO+7YaNRvJdVbohb8wm5Shd5lJAav
IUHg6JFmkUHfXCVlwd253BO+dMhUJvIn5wcXY0JrjBgRCDndMbsl3e2hnsr3RN6u
Bmrl7CigzHmvMiZk88rxoi8+JQiN08Ae+cCWsCzNhOKTFHMyjYKXZNKFUnpjrvzc
7xcy8zOx0IXse5bpaazSfVRq+ZnHLDEJz3mpFdY1l7T+EepB2svjVbHBDeGlsRWz
G3DW8np0pAqFOvLs2Ai6oOsz8x11k7wUVWAQlK6VEnUO6lWSkiBHTHVUHa1XsOQw
SjZGqRJdIM5CnYQC8oHUCdWD3ikdrAxQJ6647bRTuymHu/FJU1Kh38pCgl3HGQki
IuiJZLoNgQVm3AWs7IHEcqS901RCtqn3ZWsif+cPVuqLUhkydnnBrx7XTACKsjkZ
MjEPY8NCcSHnaXMEXGQwrXqONNXZvhc75IoTFBfA2y8kzjfFBUBsQSookGCxLr4O
BVlQqaKI8dpvVtPybGlpx1YzDOVl7li/kj7PqBA77klTWeIOur4gbMI7On3W0w73
WfeNY7fdW9jqz1YhZQFNDUPylDiiZP3qyrWdHdihpWVeYIlb/PR8OnYGxjoOB27K
gfaRsf7fuRvpU1PJWDjptZQhyIi4E6oa2HJz+8e5gA6qsj+K2rAG+YNiFvHNjjDl
4qcpPjuOyX438B/nT0jtiHPUbjAlOadV458lFwLdvrEYS/9D4mR9I3ypUgnQTe5l
hZMdkGAKwtXaf6FmPRAyRjegqluTbrOevW8G1LitC3ryRQcQ3nC2wpYRodK9to9O
yaHGGuEQ4tWawSh7re+unOR9VZz4tr8qH/0mCTVNCREABCFnX4xkGD2yYeEPRQM5
ElisRwxg2g/if/zQSmPbN4PSaLfJITnzB6NNRUcyRwxVrWWgbpBltKUooQU0Inh/
HvO1vG+7ctQZHSqI4o9OHL0kM4LHuTcqt5PghhQaDtoy2sf5D9lNsE7wLoCZrp4r
aAmpf/xTYtZgu7qjZzBsnXbftKDeJKBZJLfPm+TuKaD1eLLWht08zkl5dfz3CaRH
UCfDtozTof2SBbAOoOiSkXdXiHwixjl3Tx55e0AP5xiDS4WtllOj6KMl0rQpck89
tv2UEVj5rSr+g2R4prAB/Epv4vf5y+rI5JNwx+5nvJ61MG5rrgKGDRtHv4AoewMK
uK6Z4OFS5wJWv7NwAXCdsEVFP5QzOdmR4LiAbe1FOeFULZJTsgLTv4sT4XrItvHd
EK+DlAy7Z1xdtKGhjaSsv/s45DbeQIz6zIyW2ZQvHJpBoI5TSnP51lBBq7bi0u2j
6Mp5kF+m6ANmgwjjej63xHOjU/KsQLjq91pLK4zorbo0HJ6yZM8o65m6UlmSB5qf
nvvunf/drDGOhyYUO6UE55NrSE/6j+HfZIDjo50eh17T1+UVdGkKbYKw1icedW76
yNz28p5tMuOVPYk9sLjLjLMrTJqx8ltiGIV+2IyW0o1AbyvPGg15HcdaSQdizSFJ
874y5UYHtAv3X1ZQ7Ukf5Qep4Lviit8qe13oO3KHkefU0lo3Fku0uEcEwNXSzgEA
gCXB2KU8L37ceihOI8pqt6bPiDvkTjpGbmPDb5tFAyZNF8RayhL5I1r2ZJjYxCwG
+y3BVLUgH9+mcbeOPcpFwoxbmqCJmaSpw10d7tE7zArd6Xe749inIaPRYUTi8Yjo
v0wXDs38WJswzWdNBh9pPJRE977uE23RXOM2Lavby0TYwN1uMxaietCSupoYgWD5
2vALcYxsVMGioAnlaa/0IlquZIeGCHlHBkm1lmvbFtwSbMRnb7riOg7VoiADUGQu
UEQtL7I7x1FvuraEbxz3ayO0WLyjC5kz11a3RcMxO+rFyniqbICE37oJC7p/LoNU
7Momvx4gQ6g1sOyhFmyJ3SjdWBpdBxTtfwv0sF+ec1qgf5CW45FAiFRcXZjDUQUj
T3c1FvUWRk5+cp9vVU4f7lQFxIIEq/2FtmRu8c2Ui8I1APDfknxlJiFu3D0V8Ght
C+eNA6SmzWFqsgMEeBlM46NikVR8MJcho5jMBdDGlYEK6xNvPv5YgIZtxyRxMVWH
UkwGdwtU3Llhs6HrL3VJEhXJPLKTYOUthk4dW5qyEg1FV3jmIDnUemKt1hdax2Ez
P61Wrfl6hsJPOfEOoVQbPAm0qnLxff4aXfOA451ZgUlaEPy1ajLz0tzoSEN7GNG+
WOnO/kxrtU14S4DRUipGtY51XL3tqkTXp604zUbL0m7mD2JL1djnS7UwfJfOB3lK
x4cKMqR5r5nyeNLOUdYP5Sm70hB/+Ogy2cbgHikRAG25v1KYo9zdUgorXfYCvp4T
M5sNQSC4VhYdaQAaslSRk+TJXOiivmn/ZDlPrANHxDdscy+1M2ysa18e2WGsI8b7
ZIl7JPlnEGe2Uiw9EZwI0iO8nOdDNIw7Swen6H4P6Setv2Qu+NHB2CrQ7MQ26nbp
7MpkU4/yJCvue4L0cRq97WoVnSyG9axuM9MltiR2JZ+6eANzOFFQOEXk6b6MQgrS
FKR6Gv1Li5hHFKbVmYxeFajP61PoJi5i8PxJAOQl5GaUrQjgajatDObBUcVM3xnT
fv3y5zxCd1CFljvvOUj86mi3y2Te88tfXNzouIoihwqSBenMTBsuCtN70SrLEOfQ
oUUHTsSsU8fv8kV4o/WYgux8Xe+wtEXnebj1qyHv2+LiqElG+6vmLuVcpVdvRusU
rUq51j22RZY8coDnx4WvPkwkSyphUyTBBAdkQMcNs2rPdar15qoIPDX7jFPAOQqm
kJ7vsSL9ZFs7mr2TXxX+Hx4sm2qPezWNZx+NyucCH5UoYpjQnlpKgE8478uoO3k/
mS1vsP3ov6g7zBnvroPAehoeotkIRUVfbB/xm781oOYEYcbk053IffOpbvBtcORd
PAGI0H0i/FndokAxcN27z8uKpLxfjCwciIna/tUtm8UH92ZrYYfrxtirI/l6jK0c
rRHtGvWN4X8l1Bq5RpFMZoYkcBJY/QXjazezAn2gjtgIMF0/oAsSLhH4AAlJWMwA
T8RBB2BLH0gw1KcADaveqOnnuABSDQMOUmbstAHC4znMZSfjsBXtD+tgnuxdPO14
+2Uz1rNAepv5dUKi76AMT69QRVI5nH7OC2vB0iIxDQDDEWkAgKRUFleWtZx9UftT
v1LDrtYgakSA+FHwRk0zd/SIjUyYengQj84eMTRZ58rU47L5jWngt79GcYLwr1Zy
WrKvb2dV5WZEYYrfec3LURe5bNF8sywmtMjLG9LvMHF1SmnhZDwnuQs6orhPzaZa
rU2VsjVuXGIAkiakKZyIys7XtSGpDC5TktghOwUuh7QR/oGLx/21v3f13Oyco7po
MeeEemMmxJagMCYndYE+ORQV997T9+qhMEZElddumfLeAtZmk/sk+w52RGksBgqh
LjeA/b0wQZqCbEdHTKq7XQ2J8ytWDsS98C80xyci4/fQyZSDZ/xIg4SA5QdHSJAb
to51bALprhfOSHJlrG5R22F2J+owMikGNUac3EX6fgjGoxCkBPWsdYd5UbRUHKkd
W+MveqhBLOODXGM6lO72lHjgAySnGpWZOfqaBX0A2tkNuxLOW9cfd71cjSGtrXrp
BRumDgVix2hxj3QQ5XtbstsBFKm5IWCWUnyajdVrak+vDRohOQ3Y0VwmLHwsbQwR
4V5t3hAuH1KUbQzBbqdMJ9DV9r4hqvj+12+iXrIcHEYMJD89MRVk9OIPxBN7oCYn
jcxSxNoQE9ut4ljwyuQtNKfX1Mkwz4/8R4adf8fMOpnUbOS4luozgs1qoIslY/8O
uC0/IknfgT1Dn2JjtOq50hJvhnP3kZiO1otDnd9CwsXx4j4mcugTGBL6duCWduCl
u3SQknBMsZu5NyJco5J05DU/eeEFqw+w7MKLwzOCl8AEJ+NI9SRwtTWfCPpg8dT1
8UMoA9xJAmsMDhqHq38FCWS7o3+t7r4ckfjSSgyFNxqjSuzcB5pG3KO4xnvBQLZB
+/O6CbYSkCCKQ/6uMFZgqfIXZD08d2mO5PnthPyFYPP6BflJrsRE5go/MdzKC2JT
jEWs88jiy51ZMvjJTSbYrgjti8quwfh40wyfzOO0HpvVcqGQw8r/YBLI0XvKTk2k
fM2q8Zau+vixC9NKRfyyjeh3yHv1817fNjHAyDH8mWwjoUqjz54YZ6CbU+jYkyNg
a3nMVQK2JJNmo/LOGhSHxXh+pY2ddsXmPWJrjhsVZ2sHnQInzgYXh6FJXu2XpCrw
hUOwzv2KgU6Hg/fOJOqPOs58G+Qeqh9OV3pbVu+EGzUzEHZAze4QyFargxFr8zTc
E4RJzH3y+8R5/4Cw43DbNwwH7Vyic1kfTVZVLF/RxyzXoUMBZ6u1q5X8X046QS+0
7n9fpxFAO6QBxj0Rca5zLTpcJ6kEBzNXTZZVMEih7+n+6XGds88klJh885qOnoC8
QLCSmJAC8UIxy7JvuZd2A5LfcKc36S1lwLt+XHxnU2gKPD0dPaFbM0TS9kZIBx6p
SXsxxiYbtu5Vb9ajhVUE2g2LJ+ETElRnCXMWKrgon7OX0UO3xhBqEVwlOmOntqRr
vdCWMppsE7/WM8qvo/iQ8+8YRSyYhS8J5+wVysk6mAizlfpBYEs671pImmHeve3w
xqWN9qFYkfq58VPa1dxR1Y7JCrBNlm3sLFlP9gwbRkcDD2lVzlQPIEEhrxkI+VHL
GuVN0r++AH5juzFWU06iWX2oy4v1SySBwPa3MAyBK1Nqp+IKofx0TY3KlJuvd9DN
jZ4lU6Ls5kNBAwNjDxXkD1i/QNdkCoV8kiDs/0+kZvIGlc9nDNCZ96TAPlAkay+Q
NSifxojfIOukYnwKQohRzahPQgS/9MbgbpqolOc36ebrkxYIXYC8zZ2rN9qsU5hd
5ftH2k01cq6njpWvkYMzJEyPHS9s0qoWwN0e1ihNvUar6Ddinj1exbWrcdfcLTQ4
IGUqbWF/gH8TrUM/3lum2lKnlYt7ECGJE5nr8WVwMKNr07Ze5HfhSXi1rBE6ccad
DT/ij1BnaWVVtbS3OuF1S4CupxuyO+ScEE03ZL7wy/rpgIn1FKACYDWU/SC+ebFN
Ze1eEAqQmrn6X1SKBFbaZv1mUIbW+nwsd6eeJLPl6cuNRxSvilYgb+XUht1xRwsY
K8fQ079VQw6Ib6C3V7TyylBgAhkyTRc55phunlUkc1jiNrNtnrytrEZK1mrr+TFk
XkDkVeXIZmyEyhfimoBvSh4h0/lf1fZvKNrB92cyN9Pd7dYe4zSQUf0BnGqduqxc
UTeFwchvOL6rollPODdrd/hVPScnmmv7un1mPQZOKPEdEqAy7NIlow1AVMjHv9R+
wtlVVrA/vbP/W5jnoKYqVjTL18oH25KRBZ5xDUtWamItP7VR7Jqp9rnjucDs4ok8
Ye28NVy/AeG0H0VcxsHH7fAvjek4lglNddU58D6X6rptpTWVjhXQZAdr6DSTmF0k
4y9heAukA5Z9y5aEVCMkq9dKX7UxC89H55uEOSo4q7jnrkSQierQARX4nlybf44m
duGgeLqDSjykyXMdIgHwSaXcG9fyroQ+76RxFPWJR3G8Z9w9F33rsvMjUCwEr3xO
/dhkykWMSLe8Bo5O7fZShU70PxYpky+AwwNGd4Xkg5jdbIE/mndq4vrnGJWQ14EC
CmA3XrhmaxagH11+yDpj0nrrurJcFf84RsarDFPn+SgTklhqyRj+suKteAVVJovG
5wIPbZ8B5BMKun8ID1EpgkgkCxSjYM8rl9pogyJPKt2lbx3QyQtLFcJ3pVKT4fyn
uCyCRPxVzuWnyRyqom/Pjhs+g5aSddY9PvdDmRZStrZNS/YHB5v8kBZ02aPSjINh
xPYBZViu6NUP0YS6wfiHhm7G1ukLWXHX+OZ9khTq+YOUOD+3hrNOyc0CX7S8aq7F
2YyMrhbf4KQlMJeSZN8QMPHk8s4xlG+C/4x3ersFtJhKMOvLc2a4Jsx3by3TqNCb
RTEMIWsR4rwm8Qu7X4e3Y5nt9hs4nWMkdeZ587ufR42hNvaJqihXGCDqq2wiQDyn
53cJrHJvRcf5shkWz7W7HUXZBJz6IeCgKZFtXFt4rSINeQLLAOfl7qSFm8FWIzOs
wVEG3x9BOhaED4Ye8R9DLPiuy4DY4nkdaL9U24HtYvq2XMB6zMij7Rb47t9LMrb6
Xi8+oKmGBUwOUm5mHQiOUOM6t/3k6B1QJLK5zJmstHhHYUdOKNMVZgz36ONh91Nd
JteIAMpuiPF6061qjQ4bTGCbdAFSGxDLxJBvcALAFPBCEqjusliI+R6/TlR+PJho
+2cT3cBjH3VagB4L8KFLcy+1hf16fOhTM8PDJl+eJNFNt9FT5xgzmX/yL1C/yMXN
zHgWF4f4wRFTlaGMrgbznwHxxtbqFwnGXNAJsLL+MTmT0bGW912n9PMro4qqXUHP
tjot+xBw4TpRvJ3XuLeWppgb1DdpG1hUZ0viFhqcDB3IgXeuahq+GTPM/W2i6CCr
fdct8McGnH+lFU0I0JaKXlM2Bo8vT4G32vPSd0VYsUM1t2vHoDfVoIDqE9+cd88N
i9ur4vmcLmfb3j0WOTwsw/cJSvXaoc7ZSzhVLQ2d+fY/FZ4PTvLlZlVPOwgyddUn
74EojSUIi8b7TJXHyE0YbgwZRIv7Z522zZt6kyqKfUCYbyKJHWoUKp7x3VT6pels
IzFV60Eco46IU3pLm5IS6qOMN+I0KXPyuDrP4jmgc28w9sr84Tw8buE2aoXpjGcE
XSbfnASIJvV2Dklzh4PkH4Jn8cAyox9K17aYGhyKolJZ06m82YlnejDUjGnQ4pUT
iRF4ttSTV45bC1eiAqjD1n+NVn/V6QCz4XlEgJXf5bIb9LUsp/O+vm7pAhMU8TRN
FmpKsUsJJqJnumxaJr0BHB9MLtWEn7LoUet93NKiVLyrZYzEH7o+/j9SJg0pkHGr
vSX3BhuFl/ZurclystLzKeKI7Tlt4RzA4zVlLQTqMGsEx2M6qKwBiwVfrHnDRhou
vX7t5TD731MgPdQUGaLuWNISLuAqpcoqdtiYClSzK4FDkJcQWfRG41Bd/PonGMV4
lUvPRnq1OoEpRdsqFtShBqWqlbGh1ScojiFWsU2/y0XdeJtJd8pOaUMXPppWo1Ud
ywlSwFrJ9BKjni2ZWlxSKwlUBOwn4rMwYDTHrRGCY71uuT2EF+NnKtqLjyfpX9Am
64LQLu/1ypE048vpL16b101hRxTn1vlKfLGCLwHDEOSV2wKTFv3xiPhazFOg/6mQ
5B/0Tnzqh8uUcgIRnto1kQ7iqe3/utYS2ccXHtVGpbtyV18xFJvAFRorevuTfXEd
9fi8d0xz1tZZ0gIULm83AdY28m520dhpPiZhkyXidoqDujn2e5snTvhdMoNY/ZV1
Zd2L2U5+zK7xHCqODwHgR1F7mbgrBWWcdfccMSpDHbmtx2GmHoKgFTmy4bQELA6P
Srtj+D3+m4SDYSANe9W65VpIVdf58e1Oa4Kx1pxgmqY60i8WeoEXrAJOYHJQ6K5R
H9EeBDXbd/wgvDsYbEKuK8NRNEX5phKrhJgpPPRlA7f0MS8MqweZoUspC6HpbeyO
frXRJyBVkXKSLrcpT5YhX/vjq7NfikGW8ldocA7QhsiG5z1kx33W8gqQlv/xkQ8J
YbbZo8o2b2ComwYUfo1HgWVd2zHnyKsRtnNRbwxm9HT1ZDXl7UIFQZqGdsJCYQr5
ZsIkhO3CSLBiA3HcBV2PW7vD1kt5lZSGFTV/1yyKhuV4pPyKm+omEpCCvJCypq7c
Ip0Rt4csjTnJhmJhkuPhfXFLAZr43ZU7kD25vCxYrtpqzmdmQemKjPScrSRn/F+j
nPtEyhWSSrgCKcrM5wKaiSXW2DKHwaL3mRLgxR37DSkMN2nx8Nzabkc0mOfsSlU2
v5R7J4IMUSHkU0yGKzsMXUVUDKPAPuzW1qxxEj5HKIk/jcyJvA/mmQ3Jx7ixOUd5
YBv8UX+upZdwnBRP5RbjU/UpkbRF7m3vfobsagvbQIhPd6Uyh+PqtwUy/N6Zv8Zt
WJ3VYOcwChxS5b53EZdOnqt5SxSfo4DwIAIzgmFTcZxyBQovJQq/EfIm+cV2D4Xl
kHFECiDl4mLMj9DZ0VLyiwPT9XHvf4E586Tu+brUCEbakhs+0CzCcfK2iCviq1sa
hjHRJIfy2PTVzvNJdpvcyfqoNd+mkXYKw903ztpC9bzjC4Hk+TEpLEdYmR0p+j7B
4eKDM3/Xgcrog/NEyJZu8eDiTI4sIt/JZo/lzNH45otccaMtta+BdOtvJALc1Et1
s5Lr46aT7POXFXl1zPMdGdPAfvq1v53VchZ1Blxf5jrqJuoyqlGvDC5kyxTMy0ff
zKqRDjdCnYJ8OgOHwhX4lBx6MJOzTu7hdtfyskTOaSZsEhFI5gy4sIch0v1f34q8
ULgW8I1Zwc0oDzRZGljmXVt2WZB4DHwh930H2sBe8KFWxU1W7DHqnYqEkBBvlFOn
hU/XSlXpspDLj0GSTl/CqKS6OtsB7g9blL8ykCci9wM0UwKUYsFw/3Gs9F5aJY78
Ub2o/YsPIqc/NJ+YeKNAatA0KkncS1rBgFYMsTzYZu4pJHomlwkKpnW0Qx0cihgW
TVIAbdpzVrLycVN9beTuRkehurf946Wt6zJ1bo5cSFEOOPc1Di04qN8WjQXt0j/m
QUCed4TH+5qxeMfAxTOM09simZL6yBJRpsq1iTEfP9yK26hKUQtF5Cyw4EjwOy2i
FZD1YSjv1oPB/7IxTj/dANVcSYSlGlHojFrgf6At2y04TrcJmgMdH1YoFhZzyrCZ
QxDEvGf/iw9oCkRyPpRXsFMo/+LO2EWv+c4TK023VzL30J3y2JI+MQHl0etNbAFX
GG0R3De4QRa8gMm794XNaCduDeCpV7kcSV2F/IBmsk0xL/kt7meN23ahItXllaCt
gO+sZy7cWr6tEKyXUnT917Jm3Uy2o4n7rPlBwNPjwh09Ag1MoERai07NXaIt1gvk
r1kmONnH3s3UEMevzizY7SqAL84YMv/2sXunQk3hR4xi1+QBAQOVPAWKxYms1dMn
fvVu/oYedsR2iLLz2X3c2EepnMBOeYHk/6QTtWl4gHHPD5QUlBeiypCijiVH5HLI
w8qNxToUHzMe12Nymh2aIbmvE2w03kGDYlkRirHsWhVxo8t5sDMM9QACyZYbdQvw
p/IdQfVfthfhxdSbXAtInQOX1YQk4PGhyiN9ILy1ggPweWqYv7jzHNlOc+ix6pN5
FC8jSMuNYY5241oXShCkAtkKl1IW+8cDI3m0hvurXvY=
`pragma protect end_protected
