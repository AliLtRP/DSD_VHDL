// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:35:32 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
s0xqSmtFnVqAswQGSwTnHRasYV9dr3y5IrutCrNBdh1I3CUM0NgH6UzMfhnmHMZs
EiMrlUrSeCKkMSdcxbfAqHTd+Mf5+QAp2daab4hUuyuvDp3E139n65/rIic4vSFp
tS/OTeTvb4ASZvR7eAqqyOtA4MqNWp6NAZl/RG6CwPQ=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 3840)
VNDBwZUb61JOreXz/6X5XbO4Yg7K4efOP/DFbC1oSnx03JVgYJk1T0X5ztqFo1eG
Yj3qehohJZDCzpHQR3LuhKrSRNicvQopf3N1V7ckUSD+p5Qd9AeQc4nBBX0RjtSs
TdAzwZwkFif8PMefICsTt83KQFCZQ7nXka5IasiXsl2Ddi4VaFlEUB+Ld0NZABZL
JsJaOybwTkh5Xt17vr3ijwEYDCbqGZ/JwKTuLSc/DDW8w5eKAT04G2BYaAUmmzdU
LNUSDpCEtUjcUauR9Z3LIvsnCYPoQjfIwQi+yBz/AX6w5SbEpLckSiPCqF3B/H0r
kDSpZ4618d/srXUk9xU4EebrcMBGsskqy2Pc5IfrjadJLrEQa4EZ+O91WznqGpuI
RqeZpVUXo5kN/vI6mB4iMvlGLBORKyUZ+IYGGMk43M7vtiXDexGOuuyxS9pFww5M
+zj0CZp4px8stAUOwC8xFq2eBvcPJKIiNu43sn6FykesGzBNcQV8lLMurT1XJ2TQ
9CUXQ10ZQztmvi5yt1aXm4aNgOdwUGfg9niNq7NOxeRvgEyTqVg4Lk2Y/ShXRH7J
BoieZU28GsHaLeMx6MV5QtOLf7pYgS18WhMF9NrdooUsQBKqmvMELy+pC+4Q4ip8
nhKOMV62B7JrzlmQTZfUNofh7FRFuW9hPGkiyUI2Sawqga3U8KiqiRE7mUThcy58
u1OQ8Bzyn2hx3cdrsK/b8m0gr3kw8zOwwnecEOvroSzk6Qhu+t32Aw8+pwLLpu6Y
prbzXbCHTpLwlIIbO41+tOUjr+hTCvypSGnCiP31hm8wgZj6QSIME9Hq9aFwUFBG
RFNTwuOUJhy1JNCpt/1xSVObW85nuQ70CTLugK+udq5qPAN43m6LizhrdN04x0ni
V9+t6Dm/ktIHMV8VWAraSp5TZiqvBQpkc5R7o6e7iQgfEjBzRyiX+GVUPfGMMor4
HCzoMCSfYFCpovQpDxze7PL4KLQx18GEHCihbgVjBlhSjpZx4lRKZLq/Hsm+Ijgs
Dv1Ev+9LEXuEeAwAtOmX/Ue6nJ4bvqClpfXqiz/Z7vjHXi+srk/xD4/nqx+a2ZYG
EHOuDkjEN31Fksua+AcbSkDqIBgBlPs9GU2tmX+I2ULi/XQxXhiAUjxzaioqXE5p
yBQcS5sGMJ489WQsarV5TUPFI4H/hU5ii4wwtxqGhyBaPixuTzevnb0RlxPsPBA7
2oGjKjp3iloWYOZ9NzjL5L+HuSc3BAKzmXFGZpoRVEB190jxcMx9dke9yeoiE0Fb
iSKQxDR9a/AlJcigWFDHzllSzcJXA8f6c5Jl58ffbWK1/1ULUC0pXuTgPg6ViqaN
9BHJh+mUgEhf5lzefOrrHuIzWYlhzlv3f0CK/Z4cCvt+gLDg9OYqZ/Hrqt6vJp+f
wjKoh822TK5p2WzfhH+mz+BQWRJISYNJqLSaXcBCwgSGAIGbpvD5QClRMV+k5jJl
3/eZN7Z0AS7jwAhpSF0JeIY9Dh6Y5vakinR63gjCfAxCEleIllHkZuL4L57VO+LH
6YNO6xoSaj+lJJuuRo5e/oL1wcTUEklanBdVzSqgIexVXu5EPyxTAeSsjtFXuH9d
SQTThKJwRS6BF5l4saTaCtCamkgrPdW/5z+9ErbfdZGSUpe4mxUq7NsiSwwnb8eq
srQWi6Un6/dru+zVWcuVZJhwjtuktFxe70/nIETXgnekoVtYTE1RPKNXbDxYcgX1
0FN6lmc7507ktRoR7D6U5gcY1J9ELowcoNxX1fwQto4e+YNAeexP7bsmNfd4pSPU
4n/aWKNGbdSmG4qbX8eO/8fVhW8GDI4cNCtHP6nUCL1xd2zo1IjmuchA7aSDe3dL
FPgltAOJj6UeESe9/gxSgmLM6AsBEgSk1d3zg4oqit8b9j0YNmI4sw9ILKrDx6nA
JTMbeggrnQ0wQ2ec5M3YvUFbY9K392F4usz6LrC0DuOaTtlWMpAWe1gHc3Y/C1x5
y0ovoPL03mPJkk2zucaZo/BpdcamSR0Sgdy8L7cB174Cw+wgc0yTW1QZjOpEhBRR
LYRC5YEUnZMSFejkpGDE+7BOfl/YJc/EX/TtpsHYuS4HXB+0Mvu9knUlCfTiDgdp
70TFTVb0hJiVmD3B9tEiEVGdKutLS+SswJVW6/sQ1nTGHz4zMh+DxSaStYPzBlA4
OSy38ag+eGx/XNNYcoQumGOll1os+oft/xVYVdqfJBO0qs7HrUW1yuoOVabwIx54
4UoHTaFNxJ2U3/bYmEF6yJDLUpqticP+y4YY74Yd99X6IPSozBPJW+UM8tzEYZCm
oxdvW4OAYF1vH+WzYY8zSeN4uyCyptFbIBWlkeB40DgIrYHrxmcaUOnTzyUc0DpZ
UHlawglrIGyvcNpR/DPl451aAKF3IvuRfIJ3djLAZ7BvC28xfcphRDd8SivBfPNZ
kXgc58RIgQ9pPAm/UeNP6BDBo/WGmxyPXolYL5RyzRu8W4AxQcw6sJ8YV5njb1o1
YHGVLbDD8H0ajlJPoO7hsankq+wO99kG9xuVx7cGgNH/YZo2f18/y05SR4kqkark
IM0kxgU44OuBiJRbUSlzqkNIvLceFCm8tMAQnegQKhWFMaAsXkum6gPFShaO2OaI
fPRTtXehaiGLmQ7x7LHv38FsZRWejqi6SzHn6BU8env3Fu58b346TQBmwOL+x3t6
hlyFa5/dvcrUuzKGmgxvtRgsyKVzthp+PXn3+Bs2HDHdHbl4dvjX81wN48x0/LiO
3yYjqxJBXyOUa7jKDEXbfWAfc6UsoPF9TOauOapDmD3Zuy4iPwJMDcMMVrMkwmke
6X3YeppX7uuPgysX5r4V2Kz41dQsNQGWCHg8rttZsf7qIJkKzLaIeOn5sV1nu2uJ
IoQOL369jNgOPMNR/X8xW3X93LkM4Ofi2fcI7z8jO/3WrP0QjKAL+N8bikfCVfEb
Yv3VDFKBuumLeJ15H52174LBp5nNHI0S2C3QKwoKHJ9gbGs77lJvHicDPYSMUY6H
FM01M5hiE88AYY26ENty7bK2f4nUSa37EVmXE/GxxtiecdVc0b+oMAd5uzDrfiil
6J8op1JU3gVwnY9wwNmXf4Xpi0ETE3mVDnTDFWODYKCbPgL6D/6sqz1wh0kvcVFe
810E2OmNC1SzuO1E+ktaGnoI8yIyenNW38sx1gJgVA5/HUSPxwVzdOLQeW4N45Ra
pQvFIBXggUo+3D2E/YQSgJcCZbjj1Gl8hbwPuhy4f+Xjb4K3akCaHRCRY7TzmRJe
Q3MuyjpUY9l7GthFUQm9wO2uoTEtai9mc246nUds3rzeaphDyOcaVYRMBcRJ2ZlE
WqM82/Wpzeu7lnENR/strnqYbXL2CflsrWJtWU7sR7CqzuO+0Bj8Dss7MzEizypb
ARVF0LijBJAQKbry2LtZ5G3nbeO32HQpsoss2Qm+kTjakYGIByHLBnLLPtO35sZz
RA6aAjnQ4bqpjaTe/tXPly7kkAtcN8nlZHw9f+3jvkH9pdbmo1SMXwqvn6oprVSy
FwxkR2tlY9y3YohwnspX2C1BJqMQcUXiIxWwhG8u2QzARqavCz72l9MMrKtKobU3
IE3GRITj62PhQ0KdIHvFHqFnOi/l4Nx86IilxyRfx44zJV10hSEeVkuiUY+k8J9U
MEhUD5i17p67t8z2VnaTkT5ESTMFy6q9/VixhwJrIn9IKQ70j2l5UsPkruAnt4Bc
2H037dTOa6YWy99pOXIRs8ojhO3vnYj8qdc5CXfEH8ty7lkoZDu5unf30FYrjUiV
+N8S+vCRmiYd6VLvwfNpzd+qhjQU8hha2AZZ9eYnNunWw16X7NdWvd8QgCCFMsYC
twsVttJTY1lBb3k91YtUZHaBLAUSu+Eqg6bmvTCwadaMsRWI6bpGg3NdQgiX5u3x
m/fkNRRgF2P4ulHc2dm4SukUxBS9nhNs5/2e4k49N1y3yPvhULkpuaKmdD7FgLaa
9KZKIX9TOykNKe9NAUk1d2P/Pd5PvDBpqTumUzIFZawV3Gn1Sgm/RRsHdnyR/cXO
duXuNOlxoFXbEM0EqdXaT1iJMMmDa+luuD8c2LgXgEECmFeQ1MCdtz0D/2RqPDBj
KuNT3b4XbvL8lhldaqLspQ4WBGDtEV4lRzUzcR0AxDNmnJ5IAS1znxNhjWxdHBqr
zROXfR0kxoQ09fWhHDyCPyzLQ0JbnlLcHvcLBXlsFLPqk2Jl6BT7m1vpQv3ybP4r
Nlou62IU/l84l4Vt9F0RI/cOuO1R1IQOBa/eWUvVfY0h/voGv9hkz9OcfEpQgIdh
1VKSs+FcBhoCbgRiLXEdUNTvB3rjnZo8cwEWEBpfbx0v/J7gOkdL0tTlwTrdmW4N
FVny94cAYgciqFHAaBV0xjB0IvmNXO7vYGEAT8vNJCQ752JoOflxXhEt8GoQo8Zl
uoxAldQ7kKAt3pIy4TNcwNpFuUCco+1fCLysBefx3H9lxkbWT7jA0KAAHTErpFVn
tKAon3XJNZHTM4dRjRFHwRYobYG4ObMqWE++/Dm1U0QrTVIQJm+Vx7ztIO4564a8
3CjQZFHxslw+bLHCJlvG6hWw3e6O4UW1+KsqL34HJ+kuCEFypWpYUBU8V1vUAhz1
BoaflMouQZo234SqxpbgzvMY+N0nLu/9cgSN6Dg2pNc3usHNxlFcN6WGXGRG1b4U
vr9ABP0i5XMLPqgvF4JD21iWcMdb7yXhQyyyUACkHAlCknOPVsQJurFCj5H409al
8X8jsKVCiapoKRig2Vr7RNc575+fda1qR3XSbZH1DLFzeyPH+y2dLxDmAPyX5o2q
PLHVJHE7IwVdwoBJht0n4JylZqYZDzKlWh19NY83deAH+6p0S45RrTs1Guv+9Elw
NaI/zr21wC14CNMSzWZgnKqPdSdvh0TJoWoqzdPLOObduTm0JcW5DmkVnktMStrP
qKUuv5LwzMTzSSCW3Wd1/7sCWB32H84WKjS7+4YMAVDXD4qIgRnpVqZGWbw29sGl
FqQ9NZRnUVJN0tcaXuGAktT+McNccVPZC17Bg5Z25oR5owNM43y5fsqpDF6sCuJ7
Lu4BPqtXTc3/Fnl4iIedNMH8eR4j/EsQruxTNesYp3K6qWas+Yl+MkzbO0cP3wTR
`pragma protect end_protected
