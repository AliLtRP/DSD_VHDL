// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:37:17 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
WL3KidqaSHhGdC65V0+SYc3L7V20B032tvYqb0XaV0VaWTJEg0TBwqys4s9Q+F6V
G777JRmgqFsQ62CdjiUGc1LOD2iI1m4C1VEouQkTVpXKLvUzhLu8gV5DUkBtzQV1
DcGabdeLskDaJwoMazBeZY2jL7x+iv2Mt0B7Aqgq5RU=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 59904)
osrFNSoe0JO4weNt3n4mHJiXXLGIjnpf6mvj6753SCpwFrrr6VT7UzW6s2miO0UO
ZGI0vr+T1AylBTfHQP/+rhgTnVdNymPY5ZWGPphG6ELGDKJZZrIrRs4Q9XcOu13U
vMh7e+KYA03581wk5lvLoA/2NiWBRtle1/RfColyUUUvZfrpX4h/cDHTefknHnB7
PtaMMRCJlaR7CTfdr/NGQ5AoFc7MKt52/uT7hITS9en7UmV+p+xrnwyVWOkcXUPK
uG8360NNyCwoUtLWh2LHHKdFESdGzJX6rP5tJozWlKYuAFB5XzCezbjyCY6/Ygt1
RWEuOkiDuoVUVt4qj2jlOz0+SQCwkpMGX18JC8u+DzCasvTJq9R2zWwFNbm2Zvnt
Z4irOO9cixD8+p3qqtWavC5RmRsMd3brxYXEgLscKyS7B6AiGZGyQ2ANpk/7/fC2
vypTZeeie/BJFyoiI1mu0G2vJtCWVWk+J+hXunbAL9iCR23w6Ds6HZGboCQ1XXy+
AeqfB1vk7blQUFIF5y9BNwyWRoys6AGJ5d4WkYwc7zbsslWfvpKd7KPbvkzRBFxd
VMSHksKlZ3LmQSJTFofRnJ6H+8gdxjO3tf60ljf7Jf3kipUdYfpumw+6HAU5+0HY
wmP+xQgBwQ28MqyCwGlL/O2vzWDnh8dDSP/QsFx6BllfQ2SEAWmyRj7ONi3Aqzld
j4lBw3xVFGWB/cT756xzGmwYz6UpnITacxIKhf/Qhf9Ff0L6a0bqCYPEQkRNnfq/
QX3C7HAJbcPT7RCtqxNnae75ZT4i7X3yFACl4qsjxNBwSTfq9ndR+HrFTn4ypxrA
mJXEkozD+/6KeUAun0XQ+EQzp8uMidFpU3+cIjsx3YfCXrAEArc1UKZo84DZvyi8
r8VNDoQ102pjnfTW0qBcJR7FacSuSG8Q29AfmT2I7EhwLIlDiUkG1z5eVqg7EXJH
f0mOd6Las0yUQmkLBN2vK1iwWsmesqqNnvN2l2jcGjME3QUpnS7E2I9kwb2ti9VQ
MsagWSiYzinCa5A1oGBlAwgQ7cXzLcKFOfkUbhkJseJT/gxRD3BAZEANDfbP5+Gr
7pAk0edHo7ay1AdfVuwHakFnhtuEDkqLO4Qqdt2vZyntfENj22q1BR974g00TLpL
7QEpf4pAOv6/UqQExE2LwxYtz7Lr29XYZCp7Y5oNoh54aMPK4LS7KavkaAbYFlHd
5CAtSMhyDJsQIWicsbhIQ48PY3+nKSU+n2dihudCYQomwX1DdwYR1ARjs10bf/lt
521fwqYaA4JqHU7CyLlja31oOASkW9MCjYLndd6w9dmQCM2ywsAz0bI2N3ov58PN
Z0MitSxxJn/sob+iu/7IiWq1JkW1pNXktyQQDeRmU/e8PJudS/4qo2qZlfhQsdO/
y5wUj4MATC4oWNvZEemrDipdD/URL3U+dJrPJ7fOaGOVfcmFPQ7qlrC1Z2wBcN9G
7E7mEJQjMNgTEkjsKmwAg96FLcSpOlC+nagmyhMEx6fGmK7b9CQsTsoB27qL438w
mPTJKeOuhT/6Vv2OG3dh7VgnW4jzKy8N1hs37toovwu2RQzRoWw+Yevzh5EQdvK6
toyISqX9hqPuqysGn2jvSur0bseBlFEAZFG6Xwos+8uPtKAt1+JQP2yIphSYkDBV
cA3NKi52IH+aZLeao/x5v/a8YtNO/BjR25BYfUuodj/Zaln72LHTL1zNGg30PjkX
wFQH+srbiJ/P7kpTefhiBibd9W8LZJzzYPwn3JBa2qqklQeVvtjmT9Bg0DnXhBQC
f1aKcH/CqqDRdGHxsUGGTjMBBdyT9ECrAawqAtLBfcoIacbCAfKOV2DFpy0izTID
uyxgB+uq40/1t5y9Vbmak2De2G/lG5jRGloF04JVsML3zya8tDUSSsousW6M1ubW
ZHF4E2GttP7vFuWdX8c4LSqAIF0tEnvddPafGWySnoR//WzOhyYtcX+AhRBXd8Pb
acQFng1/IjAHJYUaUWqF0P7e4J70Faj79Xa4LBZdxBz3RKntbvcCxdvfyOWDVah1
psP81NXwb29G4trtStvwPHjfa/AihwGc9Brl6BO1hCelzc601n/7M6g+/o2ft8dY
JJyxohD/ibj8qz/zhsR0xkdGXncsrYfSpcXawyPFWvlKFjz/2wEBIBLGNPNYUbZw
MjEQcJzHBuHITi1V+IPiC7Zg0t1+lLeXnzFe9Oo1idwy2/jzcb3Tw7X0+A6CEFJo
E4YVtMnwYbmg0jfysRj4SkfHMjUdedKaOwF6z1yN+INft/LT3zRyo46wM1d6z1/5
EVBATJGb7yO1hNkVsbLz7xUNA9v7B5SH0zbUkTdGNboqQ86ng1bGPE14Lpo9Rzii
gNhZBhGz8gn1dxRkqk8p83Z3qZLVCUr9L2qVJdH1BUr27VRAKwE1KV+KHl4iyV32
nl/xg40iyy5GQlG055H50dBBiSUcBNewbgx5gy3Gr0WGqslAAolpyU13si7WeC+i
eTzR13nVvgfBaTR5k0iaOlL3PVk1zKYtHIXiel2niUwjBImjBelfwDXBUhyPFmHn
EMS4vJeUjKS+ro2CubgZa0Dpbpjs3wn7V1/CoohHJvE8wL35YPISNLtFSVbAqZ+K
f78NqtzbHAgOrctGuG/KuQEY1p2HPPCaYdIOpWzCaXfs/BIClly0PanBw3SNiEps
dA/mWzGLGgMRnOW5/pmVaEbVXm0QttLnykFuqXV5TKiS0/EYCy43q+xdm6IwKjpR
8FxSzde4Qk2YRrvCByLWS2eGhMUDlU/ytAZ8Pz78rZuTTyTlB22HJ+0Nc42OVKxS
sy4KktRuOCZvdkszGDxnlRK8YK6DokAgaXV4zsMRSpIKEYBgZie2XLS8Iof3FFCp
NKXDK8hIRrmIKIUaci+97Rffy/1VD8qKfYYlqJCki0xBHsiBu9WHIzutasz5KV4j
lAUSJ5mwn3eJIyAWWr4zZAdjH0RFOScj1ZI4EN3PXqGmRu+xk0OpHmUjeHyrarXS
D7HGDXQO/pTXEuEyoQykvDhhROzZCT1XB6uTtvvfprs+QIUkyBbxS+OgoFMkeSQ8
wh24LILVnd08VIea+qxHodiy7c55iEgSyeZHuFJSFPH/+GQJ0PUnsef209W1rzsm
pEFCK/eWPUoMe3+cnGGxIEaJ5XWkHRiesL6xqK7GUwj12v/hKucgzA1gBC6+sOsh
0fQCFuiShfsqkv0QxR72dUVAHbtWjwSaNkyfvgw5KUxASyUG5tUKi2I6WXhiudow
gcWObiK2RUVwPJYQEu6lCPfuduisC92G9W6dzAT8v3kaOkH6pNOtd/+aMASz3aJB
XElxi0R1bmhSB1y/vuHqsAWpOIQs2IJAhT9J2yt9IBMLRsIvoovOYe+Mk3Stei4e
8qkq7RpaE1QT56QRhfoVr41aZEBhxMb5+CUwSw6kNQiig4JjUp8+HJz4jvnEkXMB
Micxe8/j8d33bVBk5k9fMCHKDrs5heHjWiSXKsMGhTqmD1EVh47mESkmnc8Fw7Uo
hvf4vk/QW8ZRY1T9n6TdEJp2l9tgrPNbqxlJOt9qelsb9T7kdrpEMsAsziH08ZUH
eUg7wx5PgWPsSMr1qi/gLeL45CLaauCVqhPhNbe/VXEdXsaOYP47gEV1lmOYd/BV
czZbarKMiR+XA51P6rpAg7+cL/UnEF/+EicJZd58mnEmg5t76vUXX1xQ+8QPR7Ne
xC9myCGfk5Wmory2RMDqs3sAKMTy04D6PBdE9lFWKWuoxFsbKYGBUdhJoaNZPnyf
68/6dF9YCWPC0VbMhYL/KmSfjwEmWsMcxotKqBIV/O9LzyHEFy4wrJzRkoyAQDy/
MiZKXia2xCRF/6f0gNfPT3nW5gI7UD4pwy4Qsu29Po/5brrFWWKmHYiu6Goydu5L
LRLZrXrlnwLK5PurSksfg8oztJgzb6jnUEanpGJp3sWlqS1IPj3nts595hrlizmw
cQfrj/sNO2qIuLcX5DVUWXrNsWB1S1bP8zdd6BkV+hU9Nt1hoj8rzUVwmNampfCL
+2/eoxZueQfgd/eU/wNTiQdHqSPcg8PIItsojqFz+o9iyg89BRYW0oZ0XUkrSx7e
zzb3qgsOfE5Qr1wOC4gObKMFCL3B8/PnCDO9sLNwV9Zf6ynHgBsY5HDh/VZ7IXyq
QYsnh77GfB/tRqW+La9c7j6W0oMaP0WBNdIFAp2KVPE5/P2ramrFeFaUt9zlne7c
DS1U6x6Am/UFOxoekLKsXBfWyJLQGG7JB9LF9OFyga/4O836ycg6tFv6q/4ha+4j
1mAMzge+82sto9ydfA00mjRMaUpYtkVOyn3Yq4MX3mOD1LQ4JTPBx8zSNiE93Cee
qMs5VNJYIryIqUXurtFJLQSlHk3uV7KqqoV57yUIGzwQ3rtBD5YC3TuFx+H+d6gO
AO0mEQQoEiG/j1tFzwbQzQzcabqWCHCeBTMkk12HUzw0cZaOcIj0So/RBsBJM/ui
0IKLn8Tv+815OEqsaW7JRwSupLn05kwmJ6KiS3dU5CCGNasjRgrBuUoRUyGjGqxg
OgOq4C9FBwgjTu/ziEVtKaks0Lu08/5YRzFJYvwbzkoPscmmjoQrR+8kiqHWYOfX
nL4y4KYFGISEsjpwwcuodT+XhZp7sZdJ++2Xh+9kb8NYuyLRDtNeDTVe8t1ySjYt
dnzvbDgDshFeIJwV1SJrly4RyIzle6AViZXzrF3gOc4IyG/XUd6JH9pe/d3Ln3DI
jEggjCfBoyUmWkZFrUwUDEqnTPE4pTT/b6yPu9JDxmzw0kVeSXdQ/m4bp2DtPU75
sWK6fSmpWeoziAp6t6MdtkcZbzwTcYtMVQUVydpllImOkPzw3UJ5mana4EA4of7f
BzC1cu8EmAxyBKoBX2XHc/78fouBF5sbsuOfu+RRs+yiYRRfHnZxULNGXP/FfqpG
caWTG02PoLuPC5UVha8BB4MyXLuTseXeps0Qjbx1oKEZ/A//1+9fPS3SHAxihAia
HeRDGRDwhiltw17dQunqplMMF4b4KE3pkQnNT78NnHCdHtdGkJTyBmWOfA7UdzcP
RGMpEtrvjEIq0VMmrcLiii5YNbPUpVgLzxz3yKvkKqF1d8efDiQdeiGaFSmQP+Nv
OK0ypTyCJ918Bqmi5ANRkpB2A13xaFF5114FyMx0X9X1Mcu3huedyIztJR437Myx
wE/swr/0lA/Y/53xRaN6JmeWeeZ08eHsnLx2VFXdf7g9gwpgDYq28PJe7yB412WC
KHoDuxaHp3OWzRbQptUiYtPUGo8ApEATC8jFURMUqeseZzNJmuybUGtdSSd3Bnx8
4k6gR4gOkSc1GIIuzpoWF6wenGq44rsu5bInBZJJK2RmXE8b/sN32q+qM6jDqM9a
NHYm3/3BN7yxxjwGtAGTwtp69Ph5oexdoPaXGlC4ux6wI4h0V/iRfdK3QtsqdncV
/lYZf6degFhjBPaa+yuqZtBQf9jw16F0HjEanpnGce1ricaZ8Ju71FtU2DiMEOyt
3Sz7ySKbdAGAzB/i9iGIRaSfgSw8oyQ6gk8YgKlfIiymoBL32WqFN05WUUvYaaQU
vRvlacVDR6bHonFVknUkasyd+gFcJpaStfb2YDUEyA3LcTfn+iqASHsbeAKH8AWi
S0CxiGfNAoTj6ONoyTBCMdVBsrK6BlAhutoNVtPVdWvSUg48pvsX7n6idgFXS23i
eTEbCnO0YLVcG06JvScLtn8Fg3PhHRVqbHlMIbO5U6w5Ya9gf4DF9sIchA6k6mZ8
SvXv1yPaVKwIG72u/Vzt5BfVNXxTOyBbhOKt0v3RJMEpwxAYs+OnxdP1VTQVAto4
sxRSgfobPmHurcuzfjzb/dzx8Kcm3/cnpEGQTJZ1MR0fVS0+CKU7SnJMzh/L0dj7
3QGUn+Vkbp6rNSCJr4coSnKS7A58NQvA107Kb+MHKGyF0KZ7XUpNXzJ+hSREFAJ7
eELTHPhuIkvMYres3oxuZw+FKcwSAHX9p9fFyQZqCzScJCa9YTkysdh3D2+1Tmhm
P5/76zhLpiFHFVLjJqranwQMVwSjycHjuw8T1/uQyOQgN9cF1CmyBCagC0RStuTF
h1m/do1Vj146aWC0ol/dhL+x1V4sOzR1/S+zrIV6lb50MaO9TjoAUnDcq2leWaWy
eYR2tLZO/DpFGSNps++tn+/Scls0c27lpB3bx0pTm8ghnJHj9O0jqvDZoQX1Z4HN
fXhEVN9SQ1ygsqAd91HbqRDvBlTvuUozXNQ7nDB7uKUxOl9SFS+MBzVJ5CNyrrn+
q1LOn/umLHMFy/fyBNyyCM25yhUUZ09/n/lEWUh7WEDKz/fXcOW1mIc2xscyI6To
JrE5lsr18qLmVAzeGuVUYH36Wai48y88wyr7AdJFyzTeGH0skyXvVtJqYQmvq/nh
b33ot7W7hausBjTTI+jmHqWpkRvV8TzCKBuw//vG26YRzg4gHEQw+WWhcfvrmXSo
Cj4HO88siP2zXJOKVoKurNJdCfNltMluttBMMeipsOVnHzs7gevIeI8G+UVdUBjN
cTqO/0ChidyEtn0Nj4rNHmiqzRZHlT2gdJLVYifVkxoHuqcCU9p7i3olSpr5X1wV
3EMqm6cXV3XkPEjuEIRcTIqdm/iBOaZwhaIQA8NaMzxf71dOpRWum0+2hiszOse6
Nl9KON+0Gznp2m3FPy9HHizIKbN8jnMYrJG0xqz3c+g1meiExAIHW1TSAKk4rCyc
9Kdh1vwnc4vJaECMuSLxg0lOgS1WcV77u41WmXbvpkx0jnuv5VQ4tvfKyMq4peTU
ieJb/nwi52BlaJlCUiol3rirotPryyMzdmwtu2iKWL53ovMt9H54HXchmhS8kr78
KzuveiQnPfbHhn+WSx0axzjEWllAOo02RrHg5/ghNc6W4U8ijbodGcw7MJyDXXmv
IAkhUQe1PZAB7XY5Hv1Qprlc4Br4ZwodKPmNhrvRBylThVaaHJGNC7kmydOM5juW
HF9CIBJyS/TEpzHhl3NFzqgRF3QxoPBggZtk15hMS7+yf2J/5Lz5v2fLjOG/2bVr
9dfhJe4Tb498uEI7tF1u+q9dgiqj8wL+FgBjGRUbOzg0wQGB7XXoKQrcKrc88udb
MgcsZGuTeu46LmNYzw8qzM0OpQesjBCaf1HYgFieZg416GemUTtKNU8jBIrdb8YP
ZzAWgGWX6r0z17qRF+SrnWvYAi1RdVXwod9lpw4e9wydC5gW4+gaW3ITkq/6rBFz
+yCFlO930GNMba7CEMqJdwdomJGDJPDUFyj7qP6kDhOh5/OuUQrKCQdml2XFC7LX
BeHIOGJioiplFph6Qbb1tQqiSfuzei55DSLqgC7B0PAcPYHBwAzZ6QLqiW1khGjl
W/vrkdMECH58Pfu2egfxnjuo6MDs0oLkAKs66+rXufuFykUuWW7B5SMwTd3//3zl
5/E9ZKAXNNoI9S8+QJuoLbzABzsFnVJj8+H0Ysk0jk+q4YSMPh9ynPgZ3a8Oq7fc
KR8x23c4pMcZiWD+nCt85cAXKMkaY74FehX1Zymno45ug/r7f0wN0tcps2kVsbZ4
RZVXOsCT9fcI8tjcsROCrhDMWcoKR+cyaxkJ9mHopNJWII5Su5rhbOfHHrjRuWVY
ExEgcCXgCTPlIiOkInvCBo5GkSp6R3wZ8vsDlsB36rTCcfKHUAJ0vaghDJzDYAiu
Y266B+2WW2USuX7Jk2rW5xxb/H1Hl/22kBLN8BdfpxL7fhn4KL1ZEqTeNqOGOhyZ
Psr7Xfjd/lK9JOVT7jnyE/XSOccuzmAOpCFU88vnNOQtVqj1/wSBS2iHRemRrunF
Dg5Sa73WY83T7QxI8Gg4Wm8AJdtnuP3rYTLxhliED/g8R3i8GTvW/HO7EDojDsDv
Bn7vjaX/SSpYwonqgefVv7lhZ8wZ7A3MZoXHm/B97BSBlpXQdjIOmNNYFM8vYL3D
49TUGPrdOrXwR8d+78iB6BNDUxX3CdJO/TFmcYcl0opIyCM7WsoTq9kR9xjdJ5rc
SS1UZzSndBQFk72zZmXnVHxqfArdt0PPRRLjVG4YSW7RQo+w76B+5P188KR3D1zE
MZ18qMSHpjLjdn92I4zWqqRbmCiNp8htzjlwlfuohepfWDp7La0CBFCRyh55rGL2
mh2Bo9PKNLMrUUDKTADjxcnGxG5SZSosztCS4csUTMNpILP6kvUluXE47T4UF38g
n7chEHMD5hZalKTK7mMSmcZDSJlDNkC+CsBOFSiVF1PxzsAgV1zaHMo4I5iOdEch
5oHes7VRw/na0Sl/GHTaL4n6xYKJpk85kXmFH7KZUa38DyVuzgaEEMcq2I88LMi1
iNUSOdzovU0H+OzG8HwQlDZwyhWsy3UVP5Ik91aQ7zCTdTsNlp79jMpbmbEmlywL
mdPeFAW8x0qzY7Cne+nSodT6oe0TjlyMLq33etqpFNxzKWYIQ7c8GEVLw5nACATw
SNuTlB6qq266gFfRLYdoowSO5eOGaub1UHfNJf9xQOu0tQRFA7BFR3+8XNeL8zm1
FAZhI+ktnVGHlM7bOYcU+I5+gLtjXTw3ElbMlMPQQV6UVq09qVmFkdwpJeTGnb9c
LGFXDY7vvrPrnzCmagfTPAvm1TI/VTL5UvVZdcBbS17MURWHK3A6QpzwhtS7O+a9
COBPf1izJIGNFq6OBD7iIXDtSpqA4LzehbJl7a13UwwJGaBgMioy92CpmT/2EPof
Ea3xgcZJGP31Ox3EJyg0yx1O1fVp+LIkbEi8v2dUj0/IZMi2rD6ubrikFZspM+3O
dKMuSeqwXYTnOqWea2iFN31iP+2z2ipI2yH9IxAZJwTrXMh+cpDwcdhMu1gxAmFM
bwhsu0cg/Y9+GF2ix/7uS6ohUueCp+YYsY13XyI0b3CdtERYKwWmip1fASSP3TQB
UIi+uIPINLhVvDae7xTV9IutWRGu84cQECUt0ovlH87AxIFyC8tBHTTpMhqw9Csj
g5WdpOqjQMrMb9Z7NqUhpK8kh5c3wF9bX7N/s65m8E8THjQs9lqbcUBKbO1NXhnp
rrxa9xkRhhou85Emrmcm3GQyPgi3rMM25w2DIRNEBEMnQkvE1UWfAA+9WgQbnwJS
VWLspZnQaUavjzn+H7kpzSGCCQittlAhwz1jqBKY1ofA5T65tP8eqWa7l8phpdDU
CaSE8SCDoRYKZZd0flczGHpuSDa4IXZvjGJmyKT0BUwYdkI3rNPGeEjpI5iB5wnm
LNRJeWT0gQAwyuS8QWe5DeaQDK3J19GTfg68/+zyG4qpwCPRtJj4D8bfMzegD/7n
Wuspq6BTiQM6Bh8KnIRZMogrDzYzM1tAreoP/fTAkVdSJ5d6dUZ1ERlrtTqKgMdz
wqEWvFxXs4tanLt8cO34BMzlJ5+azWdRMRblQtAPaGDpsQfkz8ZrX369p34nViwK
gPJ820w4phnZ89a5IrMLL8uce++lTbx50yHTBHv1Vd3sCSYUjtutv+/SqVp3oXMm
qmE45Wk9g2pRRy2XSmdC1qi3FrSp3tsIijvxe7Wh6GGmI81U64uWuQ7zwQ5pTAdX
r0IwHgqTVoQfDoyxagJUye/2xpWWsllDgjq6IVu9g4Yx5rv7T8SV0PyIAYIVNVxx
9UjAX8EGjUvNcmp+ibDeNIXc+14YKZnBCDCsfb+oK/T5Uoac3NoQQwoNuCOsgJdW
S2wYpAMTkkUT2xw9JsQ9uyr9iKwrd4shV2QlXimDn3bHTg62eBcdrbu+6xHPl5Pf
wG9bCiJ5piiX9IFF63c6ckRZV9RTrutwPL5XdGejdw0QGo47wZQH4p6ZjN5UK309
UaiBQXIQtIYOiH7DujldxfV6Zk/fVwwtxwuV/t1JXqe+Mj/ZaxRbJJ0qmAGwXjk7
AGl4jJeCf2bMqDIolMHRP7Ze8wRGUqY9UMH3Pa+3co3WhjNZboSuL8hFce3TlbBm
jzxx/zixAX4jQ91Okcu4UJp2aqH7pEtjlYaRe4qNP/xlqh2QyG10riXpY7P/xMNC
sfjLNE8Grd6PzFmATYNYyXSnOOzQHOjQkQ05/nWx3k0VH9fWop5jY1r1GJFnBhkH
1fv5cu1KzhBJIYAoMtUZXGp8UX679eLtvD4RcNRNgIV0T+ZfEY8zQ+UIGT3JfXIq
+DRzRo6AfefPGJcWeUTvOVTM9foWy4ogFxVRRKmlp8Gw9wVq4xb2oJen/iVEx7pS
/j3fKdST6pUCMvVresqBNBa5V6sExhU9egT3IpRYdbyQN8Le9zrRMCgeemZsq4Dp
h3erNWAlAPaWaKqHEMzEJ4MBXhlJBGkY8PFdVT9pxmokD+0jycN8EArVwew1Q0qp
fZ2NGP8Kf7bzcJqv6Tef7cUkkUVouv4wwj7SIOxHwvNRu2Ol5NFVbNVQYxo+62Fg
4aAJpCFHWOzjCxxuFXsjrjalq9yPq78kRBETBMCMvglhtkIYOxUKsZbc+YPmPuE2
5BO6465tjLU2mN8dV+XiRAgbzOu7Vq0f5wvpFudmvbtYBawRd7s2Jhs/5TmeeLF0
orIiLNQ2l400rS2KYE3WnMec/okwi2JAkNyz9rZ4kJ7Y+OvMuHThfFfCg31fTBlt
UuFJyIZglYPVXf4jmw1heYpIywsvcBmE8frvN7hmncjTBVwZeISsG7x3K0dPni8Q
pO63kiX51y05VuaRCjkWzuViplJSTocfg8yTQJQv8TGNdfBdkiGpFD8c+eHbKwRE
7XMUBlIQeTet2ywLDfxQhlOz/aJkpBG4sXceMaldWFgnHLGjEQ2/HhTCK6cYKLNi
/+8DnDJP99PX2XJEVjs5G5Su4dBPLTg7cvY7Mrs4M3z6K4A9g8YsopgISRLgA6Tv
mio/J3KFXG5thQzBgrQ/FlosMy9TF47Y1zBth+8jtNTNvgYxqaNr+eqoO7MncQnc
aYlqoofJ4Px/kj3o5gPOf3sZl5Vx/PhB/KW7ZiDI9VK2tjv0ThQ6SeX6xrEBwAMR
7GXpHoOE1zSdQSE8PulajM1FXdHQR4b7p9QZBUjSIuxGJQcYUR7KdLDe8gbKqRYU
af7e2+6jQtQzyVl8OwI9UsssPKMeCpQBkd+8fWTvvS8p6Lz6OoYFnePGyUun7+3t
EC279uFzSw7RShNv7iyAG0vqJPhg3sldQfpMasTvU6Ua7aCt3EdhK/aRz6HryEWH
TddhXs7TQ2Ija4xh5mNb4fs10pNFR+1RAB9RvAgMGFpAmB41fUElHtvvKLsGnyZU
P1vhvza8FwSDgiZbgNClqbjGQdb9z9HercmW8IozFtZwu0FrgijqQ1JN+k0jspeF
+enhBXQzloXHY4K77Z88CULDR1Je6SV0m6vDAxi+aa07TNfaEtjykih+6ZOeuMF/
+8iTPzKo8p0Qim4FeRP1yWssSlf7vbLUXaBkIhg4+E8NzvEWnT2SpSn2YVNl8a+F
dNqAT6McM99irQ+EL/mom7KiNSfUqNlThUDDCy58R/VV/nHcrPyqPl3dc6tRaCB/
WQGv5FggkKX3guPSQhBEZSQqIUNbVPrpx/8lFO5H3zHDeLOwV1QcT7Vzgv3gEAyD
XlSNcKH5arCaqY7Jg1APl36F/uXkSKy+rOtAMXg9UBGdLIBuMX05I6VNqAdsmadQ
IxP6I3yiAt+26d1ndvdTQyalRz8e5HTKzMpFwPXxsA8mM+mlqEhUbVRY3VaGIbjA
fkJnnEO/wD1nPMJVXljtEiu2PCN7ysi6nvh/tubdRb0t//ndp7TIsegLk/7QQuMy
ehboldPTJ6TZGzze7qIwZkUPOxz3Un8NSAYRMd/s369HbvrpaZjBV23CFzqzAApr
Y4VD4/Whma43rTMx41ohcUTnUTWW9vhPS0YpR4Nt9qZKJy3DXy6lziLW+LJ1rIQe
kilCEW4fy2Jk5MsWKPuN5JFd2KlnQnOkcDpA4SKZS4WSGJ+JdIY5aaqgGOT4gkaE
7P5z/Dea/AJIQn8H87pU5EBT0wZqjIpebztZe9FiXx0iSZV/5z1vwGyChU0FYUHE
v9dTLh89/qn0IZWaxmo90lJNZMhLVZ2ohoCgwRVQ4GpTQcrGg+VcHxX2hdMlKvWa
Ka3/DnR0p9X+XgwIK9Ajr1B9MoAVRfCwQK0aCu64ECNaQGCptlEGdZB/4N789kjz
Bgn/O+cTwLb63hOrWpQ/blvZe3S9VDT3AqGICNt3V36YCcOoOBLUFJW+5AKcawJL
lyqn2DQs4R5yqDs3KuSODsTS+zzg/31U7mqUg3gFjsK9cT29r7E8expQUcZJoJlz
xshAPQ1xzkd8AdBvtLEst0/u69mvjmNmAs58To/dq2Tnnlg8CXeXmkM79CHHu8fl
aWwAqjZ9JQkEh3YxAv+wyBw+bjj/pCHC/La/wPrJjOecofsAVo8Lw1KQ6IpNPz1x
dK3tzixWnblwPZXPE2CSGtesg2FkxflzjHP2F99HQ2R7ah0bEPC1tZm9vS38rycf
soG/p4p7s6L+X+DipTNNvdc5Sg18Px7mvPL7NvMoI9sXQ3MzS/rmiUP7qXCatwqA
x6voDQJdWHE9olWoBcztz72FID4ljVG04QbuHObr0UYFw1C8DUKluUvW4yKtj0rf
R3jmiAV7hcviFe99yx26vmBg+NxQZUlcU19ksNUMdmQi/T0764fV62A/DFz4+d74
NVFlHooyGg6pfrKxl3SXK5F5OlNNdHOYN6qzNz0cfG6oIg2z4Ba5Hr9jjKtV6N2b
52YZpCPdOyASpMXT/o54dsbu0qE9lVvfkysxWldhSlErhoF6gRi8kfk3/p5IVhM9
YkwmA8uWCBgbyuPoAjAbWoWdimXDZRZ+nEF58cD+l9myjEDFeCJxRA6tod3CfT8N
lXptvH4SZjxioK0gvNZuenvSiUcISM+esPSfnZVa2QzIizm78ctEPmDrAg3MgkHh
4GBbrjI4ax8uiZs7tB3/QmjyDeD2ZLKZPH0Dp6oRZGtJ5KC7cy9ABhKYuPZl+MBN
djV9ZvAVTtmz84z64q5mBH39htgOQ8vOMZ04peBUwGY8l0TuTeMgRioU7ynzNoul
c/32mYXZR5P+LHth7KVueoMWbcfJcXk+S1rnwRCmbFmGrwUOvCJI4rGzm9voCBXP
/SP/CoeGXBApbLxLomIDKu2GAyEmQdlLHgCz64edipT1hZlkTcjckWDguxuV1cB+
t0Z2zImuK7IQX4TjHbWTVfw8fMzyUcZmKcW3dYnrO93/F1jiLl+VExo5wD5S5Xy2
4OBT+vB+XPdb//kkCkOVZv0Q3zKz+gzRaawMMNaN6qdnnabY9j8d0W0ccuaBrZ8j
sAhmQRXHenam4izc3EldBIh59zepOeCyYJMt8+FVdcHco4zhSY1SM8BwxXXeindG
kMak+H6172k3r5KLt61hzRQo65m8JEXLYghXOsQhHCHAF9kmnts0KRH8Km2IHmts
R8sG5IPsD3aec4l8qqIwn3KiZ40/sHw9uNIq5VJJjhHSGOMbGIpLDD5Ck1a55vzM
IZi5iJBNsyikpQDuNMHQOIKlwq7farun1XGZrUyeEKhWrjOdyYOaCelztfWf9qHo
Q/b7JHnP1HkidTTc+WsVyLRs+DZlaDohB/U3frzRc12WTjHv4vUxX+GUUxASjD15
ci1uS8OUlzFjvs2+lAsJ/8tv6N/x8qc9qm4sqc8VisS3ef82DBgZGI8LakqGH71O
Si+x1AihJmUFJZhJ1BYBc9SaVhLfWMOJsnC+hNmw841CytZOZ6j/jwrbtl5sGBK4
ofh6gxKwenIVfLjHte6EoAzJy6zk7aUuJgaVpgLiahw3NaoEy2bztJx91vH9VIC7
e9X2KVzGeMrb/G5SGxQA8ctp6d7CIVEbcLG+RaX9Wl/g8HMW2+eS2UicbnQROs0t
2zb+NlyqZC2hO0twYEjaebjIIjt/semS9I7YKFN/RYVlMtu2eCf6W0hF0mPk/mfG
l3B2fkizut0KVfEvKte0u4YD5XgFywpsIGvi/fLlnG3iehS6y18EOATLOwPzNr3J
PrX5D9AFrT4mI7o1PZIe65DlTUmmIZWN4+M9fuXykfiaXUd3F80HwABVZQ1XptfR
W/5GuAH0UwcWa0O7ZqDLC1P9uPSmCjN+KPZXiTUasoIQ5VrWCWcboA1baifLPx7U
aCCxHD40xS3BXeLt65Xixj+nAtKhHPMR+QRoXhTISCPJ9SahZKz2qxkr9ut/+X19
bAogNVEuIdavbXtl78zPwS+PqA/Rh91RMocpM89ttxk7yHRfK9XHqIetuMqm3rVm
bhhRNN/nNYnGjAgVRKdu+2FxjZw8jgYK+8LtpuEzOaGWzL2g54KvcuoNA0O3gJLT
UD7K1fyvajYqoikMtiQN9cqpRwXRxFWtupCwi/w2egFi8h8lag48Vhz7T0D00mVP
oIsxKrPpqVVFZfEEokIX9wwMre0d8DxMJqwj95LfW4EWVaKIZmlgVqd+Xc4gc6wO
Fiw2ap3IrnHIUo/wBzacOd4cfSRP4JHy7rUUfjjOSBnz8tN6LJNVha0s2YlHiDZa
sGnVhtzz4v+z0QNk/ZBYGmzoo9tpy59V6y2O5b1p0Dzu451TzxL3j4C8EGDtapWs
5bzNvJozkvlsgygdcAd+wO78ICJ4zJsHPXvbeapIVarCQqXiCl0bNGJHtlGFWTK6
cUEeZFyZHksVK9CkVVcQ+3i2/uvH0PLaOzGIbcmuv/oztXzunfDvSNFbyWQmQMlT
BegBSo979aIK3yiS3KJmd3AvaGhiyBv0/4ixLIdNvNqxlJQaNcS8VSU/+BtgmK+e
SQumFcmEBBAxYMxhaEyFrBep3rddtulOQiX3/ZzGhfxA56IB5aTo+Jml5u9SPa8C
3NLPiyPwtTO+tE6F6CRnir65ceksO+PXEXINVoM8MxP6DbGwkYl6Y7DmzWzRapWm
it3qbd324z5V4D94u7Nb57Fw4lSGkioIzkZ+o1okbt7U/R+3kxmONfJXEX4roNB+
m7byY5LBOjM23CLcUx4n6hMGFdosB4Z7Yh4qMI6UfO3rWIXOqB2P1i0LfZsfLW1s
xyGPjjFyYqnEyxBntV/I3ferQmugdF3Lhy6Q9a3lqBqN6lpPY+ZaIJ65jk3eQp9o
z7hLpjmhwpQ7oyWILvqVW7T4vDZGIXUzMbu0FWRpvvfUEkZnjG8os3ggs3WnqW0n
o60FLVwsvS/K1EJXiVKWtyWu/JF5dY5AjG90i5qfXPzoDMjxggPb9xFAGj4iH/66
xKgf4LGdjDG/jkLNgqDB4LKAsl9TQQ96Dbl1RqIGFFYumoYxuMCFdB1cpqekIPg8
58Lv0pppnbsRtdi5ZGXdhzJgxqL7Z8hl1v7VuT3+qBn8SMuzXgD5XYlkaj/AA/x/
zGvxp1gew/007DZEEBVPlOGFGP1lkZd8ROQNSQEDrEBhqy0saaNt1fLmjFh0TSiW
hYfW2BwquskudEpjOTk4TpAtlk1cqDAFrkffy/mN0wh15e0LxBdeYTemx2WCpjcn
0jJBpX1ZcevKu6x6vRVsIfVHuk2A9oIrHgkrtbauqePzA7hetoKLjuugaDumEpu5
pfKyj8RMge72waS3kVVVgB/h7agWHXOZxLfy4MUbmF0IbLYmQhiMk+YHZvUKMRCj
Ht9UqHOJucT786/esDNsWQQ/HoK+FNIzcqqA45oz1n4bKcme1BA7qEgfZEoPUHIn
6zyQW/GbJPuJfylvIzuqFXHUOrjMoAp3/cj8FPh26zGduxiFpBlCX2yoM5WsK1Mn
elzIiKgZUc5dudqFxWuAh/w3/58VQ/MRz5uZch+NSIYLMMV0A85AA+YRWZcRacTw
me264TQF9LBclHMqNCwvAOC0MohLaRlxNiEzZaX5jE9W6+eOtWiXkt2BL2WHYKfb
nJfiIWQOLGrQJZqhzSqS3HbC0AhD/3hnWndY4417Tg7Kd8YZEN9m4OyfC+AZ0EZ5
xFnm06xrFdJB9YI0hz0LFuCoYNnHGP4/kT8XpIgLglC6pdqPsAfqOdAeGXshh7i/
6XhTD2NuSxW/Wa0REpX+gemBDXZPF+OD/d9e+ARCiSuBHwcAs9UD2W3YuSGvlso8
XKY7b2DL4CdJHyKCSqIo+rpI6szVOUyc/jybXedpjh4+XDjWHqHG73eDndC8oRVC
gxp+Aud7lECF+mYyYTzJw3khxlI6gnC4gOif3J2CA4NabWqHvB9WlVmCZ6hfzjj6
HUztj4LIfCd6m/l8fWWy7SSD2Ao9Ya/p/pm5c+H1voMq3G3EVlSq19TNOl6fCt21
ZujrTjp/6OcvdUGMrDQfVebslrkZUHLpjhbI9EqWdB7TS/tcSIahOyI2vbaDB64L
gAfHfrBdQFD7nixQXO9UZPLE33I2c7+5jYmmTS5T9iLVJSMpHSGqit1914sH3Zes
fDjVwpQiyLlIWRvK/8k/RKBA0le7LJq60iSiC5HCQicekG+HzKgWprxImd0dR/Zo
FzWzQeryYAyBO5D+CtWIDY6rI6XSTN3LcamUrl4CUhkYUhKhtR1HW5QyJNTvta7o
+J40t8sdcjpbimlYE9aT5lQYlEEGn0h2N1D0cvmGWwsfFjYfjGADwOTAMsTFpsFa
vmU988z9WESWeZpwdPEMPBLCycBENNUArhZGuj8crr1G71hZyMZdXFn8M9jrIEzJ
3s5LCuJ3v5RE13PJ/16IKqPFYQRRz2SiVdfgu8q/Sp2yP5aYBp9elT6okDyJ/9Bk
k62FFQ/6rbP/ntGgnou99qjkrcEktoGwZi+sZY7/hTQkzgQUZ3zHRAGvrmrpSq0J
A6/KMWIQbr3S15raC9orYkJLTRudkoYJVtDxCU7y9mZC/CTJ43Il5pYS9Ho1DPam
LZdYPGagcQIwI797J2uGzRBWD6gHTyjuYvxRJxrffMxEbhMg8Ja7RnwTWk81qgYw
GBkxUdWmmr7MuB7X/M8td4aS88dgHwzwJoi2+JzLnJ6VNVK6XzqF7W2M/RDwQ2Pt
irQSGp+p37XSqqXl+lWnnOqZ9AqkhuqD3Kk+aDEpD9zk3p9VdUJ91hfLolk1QYMd
NC0vXIy1pJBzkVmRLrYqc9FcaQvb9k0TcknQ4sRTW7Dnq1k23S6BKbOgIP9rRNDu
6ucfNvgTvK+N5+7Zu6WvdDOdjnUQ81eyImDvtIgphTfajDqaF0qNiVkCToAmMhJf
MLR3eqWWihoQ89OlHPNI1cijlHkAd4nFY3WHTUe6pmfIsIbcbJVvumNE8ZhWQe2M
rw6CojThYvUbL1Wc9Rfz4UaVXakJst+/0TFlFcSr4M1+X0VasJ6Lpufw+BNW1gov
apO/BLrGZEkUEb+U5IA83gP0Qzj2uE+0t9/xB8+iAOXIczWCChJZ327er4e7OEeR
wzi70e0eMXXl0EwM7xsUGrorh2CgJIOi5rJxQM4d/Y1iqOkynch6fJn4AJhXXUZI
0tK2+DxA8JMDC2WdUNeDI3xRPaBAmRpfjaq2+QWhhY8NagjnkB2sjb98TXsvyJ70
5V2mcWKKK7aKsmpaYEy3Svr4EtGMisPppwczPzUyHcvff7RclV5HjYHqyLm2hX8z
Ug31xq45egGDbVNbBz0j0WcWWZeuFrsSIY4kp+El8sC+OVxmphAejTeP6D3Y8L8S
srj0QCuvH3xFP3H/97wL0LD0tlcVBpzoZMpGWVH3zy5puLKCEAgap8NLop87ZGzt
EWDpVABcQns+8RDsJqd4qFUuiJ7k4FT3qnveUzkrel3wFxF1MWmi6gGijrPcwVbc
kb8nEdjLXf2zmg7IVppwE/5vwkZUTZYyeWsrHibGyVi7Ai/LpMnCQDPWfyniZZGW
nEo7JthNYpwEYqLJHeSOAOOkXS3+Fn15T4Nz4sHsK0urBOoDFBvJksuvnnDbeLU0
fRz90Iq1RNWYeFpJrMIHiDi3wir5TyyYT11hkFSg6fQdb3lEBq4cH4/JOeADeJ48
kkN8EfCpK5ITv0w12RFpbPvNuG8CiYA12EQ44ldtdKUEw+1MZyp69FDUxCu+Z2g2
LE5mXye0P9nsPTFV3COk9RwnGzwnrkFaoR9G8G277o865XdYdJF1nxc4/uQzQl6Q
owEleUrteReSlK/JUISQxewQFCoNQoVIgn4kNWUdv+hKqBtS9vAdtPARHpghkMcU
BhKo7Wv3kefPJkz4QXOkbT4n4DDlPYWxz6HHJLDfk739uOCWTCp5kfH5VWZOqG3C
VNfCtLdMcBA7FTDY5mUr5cD72pRNhi5B936fW6OiKrFB0EsHqwX+4VZPcmQaI4cj
A+s9xczDA367/QXdqWIXX5GLN94NMT/zaqdw8WcdzT0G2Y5cNCHAbzEpWTB2mkLg
FEYICYUeUHT1e/e6elYky/j0wIYh6pSNC+mlSA8/F6Dc0JhTOXMimfg4EJwquAQ3
Inxs33aJGTb8xicu7Lk/UviYKMbNWb94A9ZmZOZSnEeEmiPwTK68xefqD4adU5NU
oCAqD16YU0b8v5Fus4JLqT8I2k92bIYh2QkZ46/xYPytCRFEZjHs14JPC3h2xNfJ
wQgfTE2ZNYGnACh7WKfFW0wcpFGbcQy81SM+1o03evpEctYBarw84/EDB7QC8tYv
kSownbL4hF5EmTGIppPNZSHYbDGSh++nrLFqR0B1/64I6Mv6vtLGO+VPl/R4pVaq
Zh2BzNSrzYb11NJIByOiJbP8G3+RKWXVdVD1MN4+qs/y2GgAJJh3mh1Mkq8Xj4/t
uCu/NrJ3KbkmOK1xMorYMgjh6JqazzeXmma8LZcQK72sUZ7Qvv6wcR+5kUQ16U1g
3xTkcN6wor9OMybxKsq+YffQC+2LjQHrdIQv81BEXoxw0v6PJKxEE0bSHCrp4x98
sVGAtX15PaV/1/e3uK/jjP0BFzBCDiNd0dpYOH+twqlE+gYc0egmzim4tnegshfo
gizpYINbruMqFmCd7+2rL6U9G/LqbUeYfyAI12P+GsxUk6SPeupo5fSMJv1gbN0Z
iStS5I3XbGZGFXRmrTCmWTWWgvFBZM+cUClh2D6jkN9lZ2EqZT3wGsnZ8AGYkVzJ
wgLl4/L4MTP4XV7x1uVv0v1ij2dCCVjAG9QvRpVONEV07lgmSmAr7KiFKm/eg8mM
jRjrD+knireS4s2YWoU/cET3CcjC8p4rs6VYzstBJQGTn7n8eOI0gOuRvatWiOFV
PofT1lKBSAgZH9QkINjMaHnPpXMgID43PbcUXNb3Y14YWKW0SGJMCaLxeWsKdGKV
zggzsnuRxVV5M15SISNrMqwStSDcdtRmX2Yt2u0k/QaBr24mNKEgZoiZhXO8Eu+Y
nUjmbA2HNd/7Zii8+Av3okcN7knMRleXgnJF40sbHz3a+0qR38r9vjFYWpj7P3iv
rbNpJvpFdZgTHe4mbdq5Xf6ooDdcXIUwcikwPGam3LorG1ny7POy0UcztwZ+3luP
1oOGeOH5ZxrHmpTDnC+0iV9ioD7z+WNhLsfkAD50NyqmXKeIm+O77jrIVZ6ZsB6Q
8eXp7wvMt3MXvxUAc04jfwJzsT2R0wRT6XtDL2n4wuqj1bcFqFFA7yCfys4SQrkQ
77sHdMlGRUS2fpISo3wXxmub9RUYmaCVfI+IhKElZTzoRHU3SPBPMhvhNif6PRYy
x/xXjPaCmAz4I8eFSnsuFPrOXAkyQ35Wxr8fKR0/Lalp6k17fNooWRTCsJuUvT29
jB2frmgrlHfAv1l76kxqMvMn3h+IodSQ6vHO9jMz5Sk9I0y40HX3fSkRiiRTWAch
odxPut3fsmBkVykfMI7xioYKtGDnGdReeMZCd8i35JF/u032iGgbFi5Op0ibZF0v
GfM8JJVB879H6OGSiT1EeDFpYIvV8xY7q89VnhmMc0ueLYtA0GVHTkjEu09wSp5p
LNGiwur06f2p42HZtkFR+qXWyYlNR3JtiV31/6DUEXRZYwnbAI2r6lkLZuR2N9hK
GWinPBlqx8L8d1C/WChCUbtJQR/TlNW7Zvrkl+xKyYLieRn+LxOdYgX/1uN636oq
YxuGwDmAyMbGWNKBVTZun1jghydFyf0HlbSex20SGhrJVfgg6sRncKbT7/f/qopl
FiBnT98uj3Wor5TeTJsi1Qh2JNc4PYmJ86MjNEC4FomsWpvqoPQOpGT+W6Z6Mvuv
e8pBvjuc6ENjV7g7hmk9spExqMcmFmoZu9456KK+C3dFXNQprfBOBVwoIjC/A2OU
SpFt2J+0aljKwqIYDExQqEGReox6AJNQ97yoMs/+PyGIWKmbKpUEwmHL17HKm1ni
+0RJjYx/ggDPmVW/CYElQrWV+xhhROh7ivzz1A1Hzz0uS/QlSENUUc6NsjBG5I9U
h435t23AzR1ZA87PEB7U1I2+0xaZ2JK647PD7npfGTBpCjh7K8xZOoDbIJIMSjEP
TOOmvzYHX711K1OmStU0QxwTE0N8DkLXM5H3jeuobe8ZqStZQYCdFnhIt9O4MaSh
b4kQknCP2ccHCGmAOBuLqXMJvGb3aJHs6lCa0xA6p5SiOGa2yOtZzAaF9kX+GrjA
yMe+6zi4goNsBKyxfD1i64jeV7lPo83U4E4bpH4AvQMqkYKeLJK6LrR9yrNgGikg
jP0fnFbrO8G5pZt5LYa0+dou9OZzsdGSbZNxLEeg0Rsm6gSrnRaL9xmrcTGzHhH4
G02qi+EqQsskb7JFqoYOxMJT8foJ/SHFq5lOTPK6ciT1DUs2MoXxT5AG+J8lludm
99y5H7jaUvJGif87RGusbAnMWuXe0i4gIZIQTIivCaZuhH88pxBY/UGPW29V5CXb
fjOxbLJnilU6R5FQFV5R12fIj59oBjXV3TbB6MndYsaVehxdOd8GKH+pmfH7FKiQ
JWiV5qlYYAo8E/rE05BfJsQAMlQF0zDK05+mBfVyuA7ahIvmoD/2/ivDJwPaOooL
qkTJw6ewbxTY5luQixk9IVgMBwWbED1WpV7+hy8FXQRDa4QQ6W9IOkSgG5tswisI
FwilQoD4+GnUsqPt6TacHaNm9nfyj203z4R8e9fDioXnIy2srWggtwBGngQg5Dgh
K+yKJMLYJ5lw6HzU0mCy3wb7qDKQVBqGw0WSJ6gFLQhLDAUvyBHT69riQdpefCYN
KV4cPyUYOdD7k/Z5v7DxGgW9YIUN2X3c1YXrh1Q8R3V9u5xtwvLBys/QCeV1oXz9
vQstMfMNpiYMNHvydZWj0vLwLuJQA5odz2f6+vFSC5k60Zw3bcHBNx1+YxOK7GgG
rObiYVOT+gxnUzBtb2Cbbkccu3JhaWdXNEf1fKg48+UOVV4WC7MwXBFS+6MEJd9O
W5O0O3WJtQ3+iW+aiAt/hthVL2Woe1/3OgWqsrowC0DuPeXQYzYdrM6vDzrtk7Mi
vwlWigzYtNECh6uqr/AXHKpYJn9FhoZcE9qMVRVkhod6EmJWefH/TjVICIk3Mao7
MW2mO5RypdHGTqc7zt1bwNsfLTk5xp1y35GLyTvzQA6+fJuhEh5+T4KzFAwZIuDV
hmx3/fUwUlvJQrZ/9dxWr9WrDsLJP/STsAAJZeO3WQKYLe8Xf1zY7GH7qF/LEwP9
rPohRJsE1VreQBPjhzGTdy6KobWsAvLzQe2Hx9r412oU7nJ/z8xTCmuzb/IDnytp
taG621YS52heKDF0hsZ0nI4zJIRkExNty9xksvUGfyeFSUzAEuCmlZGkYuqdaE1j
mCZ58XPrYsJwElp0qAAE0GrmDYhtANnlu/nbWaU+SFhWvsbVn+3pfTA9HlW+sCXw
VcnJtvWvcPAREGT3PagNtQkb0LbZPJ8fIQ4hkXjueHziKxEpwTkiPkUVs7J9/gI7
Ac//l1EIWrDlPCF9PVvk5mQR+F2Kj93BeVTYYy1FN/BcBMLV+wmNoFtYxdC2CU6G
EMgvH2Vvmhr1benJIdHG5RBWZMKnkFjsaFJ/9MtDTtrd+apQVHC3TMRXaFTmKuKG
a8LDhYqQ0SEy0r9Sr5ItmuVYS6hHTmJHOHzszRgY7hdKVTnS1+dh3Qm+m2q3spgA
ciKmobPX+LJekvpk4zTAuwgpgmzN/WZvpugqedvdowXGJ9+YlvnLkGoB10L25/DX
UjDTs+DlYoLGcVySnnJzRvJoAcd7Nt68cNnnhH0ZZua6fs7KsOS2HGHD9tWLC3ep
N5ubnZIGZdUd3YbWehZMLanZnarR5qXYFxZT0XMlsDkhiX4QlMfdmTDtGDYsWmB6
Mhc0jrp/tHJwKU7knlG/dgFCgwcRLKjQK3whnt+oL/RWvk1QjBRC/5xKX9YuZXVF
UTImMMqAjlewtt4q64j6xxBWMQJzCXOnQkL5fDGrBf4UgshX7o/WBzo7w2eoluvs
KnVw6v7hPD3ZKcURpTsGxTnH4PCEfQrRPhUvpMoJWOynOhsM4roXoEGAH0OzAxav
86yZIqeR8V4QixitkKI7LUhphR/j05i1NnwkQ4Y9sK/vQOtZRBRNeUAZwwLI75A4
4pZtiUqJgAFq6hNGtleHueBdQYDIEeYi8DDS4sJxxFDgRgo9PwOz8AAdhxCjMHUO
XkbDUaJQy4F+1/ExTtCSGPCW3xN2oxWo6/AtdYJXL9rPVbyQU2lxZJacB3d+uq9V
C9MYn/dBc8J5YdWzrF3xxL2EQB6nDqNSxRmwpFaRKDTfYeNm0coULPOyXm1eKKyH
D3eVswPP9dqfudXfQs1/sZEaBY0R1MPPMJMvWs2QQxLMmnG8gqz994/KBSwPH0Rc
+Cc6kE+gsVSSFm7QxJAHjhrZqGSTbYrBvAO9uqWe00iRG3uxaQo8efasNHVNSCyE
ktK1DO8vJshlxww7YkZ6phIycF1QQ27w/7ix4eLCFLhjmaRGlJEpCCWCQQcMms9I
1PLNsrFQwwr30yD4hQpKTxDZ/yEqbh3kANTfa6V4lVUnqsC9adyhFN00NA2SEcgl
M8kava7Dl3dsQysGG4HmjtTgqGg/xVhDjCc36f+vJMWf17aDHYgy668mUOcLSO5E
Mu2BBJ2jW7IMOTdCxdnmL6QTnNkMCuM74xZePiH53zRKFZJE4m6U/zR/nLabaxvM
YavT1tRECTz6dFZC4mB/1B/jf1rkP1kl1swZYxx4uMKmmDqF8gtorsnKzeZu4CyB
tTVsguJsx5fW2Qmug8aZBpP28cUIWeWu/w97UZ6ZbnwUO3xPJCCT1zSWpF6DLwt0
rFgKN8g+6/OiTUIMUcJXu7clVi5349FoKad2g4Zx89zSn2bAoGeMvFPauUFdj3e3
tCTKqDjCbbKC/nmNnpjfgWaqJNyDW3eXp3XZyMR/Q/t/N16PvvDepomMnmB34rkY
TfiUKqAyTKt/SJlTsCMZjyBu00b0ykmCskj3sbY3RJVWIGPdlGQqElBYGXvMaTjJ
hxOfdFLvq2mJB9KI/pBzv+D4453Kj1YwvfvHTA5rqij+WTMY+nfyevfM3+qN2v81
5KWluiWXH+WyHDIh6O44ce1lVz0vxPS+LcCXb2/vHhYrdv2ke1m8CGfws7iM//QO
I8rC3JfivOjSXu2A2vU76lyGVP5BtW74akOQALjIXEiT8AEsZ7+GLRnNkgaLkpmn
zuaPIg/e2lYxWkjs/58Ooe67HxJshFrhH9xexhJrcHcWShU1XmwqMSxH6icYtmMq
lpxvneoKHmm5KHIhZezqq0yo3NVPZXi2H54dGlKZURGckl4FAnJ1CBdhMYbB88SD
U9Mzf7vyJm2LX/WMYSpzQY5/RzLg8LO6Pb/d1XuYuYoSO3b78mVXn7B9G+8Tw8ho
r+NrpKnoznDGRmSuyvjZJafSlqsPM6/R71sl/IeZrOJGlfv7R+MBhm3xtt9WfXJ2
88PEsJ+NhLIdSdR3O8rl3zVhVlZkM7+RJgn1pBfbEyI7gPHulCitEvVxscHAFqmw
zhzslDQ1Qc+JeZOuJ6FgbHpI56IWHA+NKQlFDXh8TMNxgVZsZEkNf6Vw9fpeukcj
35A4cwsu6wSZ2aB/5OclMeOclUdRo53C3RX4GUynBh8MKDTWEZ34hJbh1amCuW6g
T6yc2E9eSSoldzRI102yDYbvGZ9hM9Zx0c8m8KbyLH0HWEidWJjCx931GmyRPb94
f9/FTd7mTejYOoJKeUFDWo/SRID/eOmgGkHs8tlUPV+oPi0ChYhtc2dtMf0SYs+T
V5vKdMEaIa1h+vvZHrKrrKYofEoWVF8E0/gtLBeBPv0cAtjrEs9itkqBHH5f08Kj
EZ+ShGgMq6AfJ10B+8O+U/kUbaeVTbBpnJ63S9xCbKFQ2pqbHLjqn5ZP8Y9/KQmZ
02Y5bCoQL451hpFuBzMWpMwbK0b7XeihLFnFI1Bv6K68TYZSE9KKejiKOWcusj0L
uFqI2wT+94M7dECPHN9RzDuYhj6UIEeT5t3b166XjpOAgET17wrWPjKgO4lzKERm
6BOs/SJPwTfuCC3fBZbGMoSRyilr68BxQZ3Wz3mg8tanMqyGGHtu8i5eXJwR6zWq
UkRRGGVociG03arpn1J3j/pEA/UzY+QneTQmAXSTHdaitzLPSh4jf1W8B2voy221
NVg7MDUkR10jp+pmNHU7QeAwASUSIUcsY4aNcF0AFMsEhe5R/80nLWom7j2mW4ze
bo+ZXSxweBYgkMx89bKfdJNWFFjhfMSFoqNMFM+dYGtC5V2yh+LEjQctJElRNH6i
zB0vX+FPibYPuywOyO8mTUH/zTvJ6aaJQjm/4G9OgASd+nG2MRFFb9iKRZuZBS1l
fb7aGS3tu1uW+i/jFTSV0/hIeaSUZr9VtpGwHUz8/qCXcGsJATZvbeSq2GGZZxcT
iopmGgtEeOiGO646/tE0D/e04JW/JIkLlvleKH0Rmux4aAemH+MzgpOTS+6wJ+Ka
/zM4VF+h/D9G1PeRvtNxsAS/TCQhoZKUHCTTK1+os7UCo3UiMLXik/trPlbV7adL
pRLLpOdiQUHXCiVdXhMv5kbGM5MSg4fDqrKgEwNFyfDgQbTlckPNA+YTiW8jNO93
QBZ1DkJsBj3oUqYbWnFotuHVjRynUhOXCMg48WfEDXf2aYc9aLhXTyul6I/wigMy
JwDciZguN4bzI0nUqzmbCoQRN7nrE2x10xcrRTQYuW09G0bd2K+Xg2gHC32DPqhV
m0gkNExvTDYf465hoYvL8WIjouflF+sN7D92T5/5qR1drSey9g0qONYX7P51Mkji
7jecb4wrd0rZdLrfyXjcqTYPpelKarFvzczkObLXsg8VtU/s43SBz+a31tVyqW7e
QMfYfXMsIdy2eVUdRRY/G1XpzdgeYMzdiL+t9g2ZhtitvDj/4zei3nJD21t96HlL
N/NCuO0Or+S6hSlCF6hQsbN+nb7jitu5F0juDMvcGJ1/PnHqVDkEC/ljt6b3+AlV
bHxoD6m6qaWng2567lbrqBnCZ5N7jt1h0OhDtBua2lKFuEclZycyVYn81kIT9+71
4muvBAMbSt9EcWVJOyZUTvGCQz5WRmeQlQFDn770Kfsr3XlBv3S071AEZ5Jgyxnb
ntAS8c7krD9+JzpquCHI0ORdwMYa3ipGtFym1GrdAymJTiQKNsiMOWdmNAq8tWq7
uLKYNV/yVEc2PKocvwaAUtuRwCYzQfuQ/lFy5mvTSFnIbyeUv1DOR7xKMrTzhOnw
GS+W3EVkCHPiCkMuOPjjC/kHT3M7Kkwj/nrjIV5/XEzc08CtV4vr4zWsTQE2Zddn
1DB14NI0EvvawJrcOKZUUBRHmj67kKBQVSUTCewOoPYxNL7HWzdQNKGEzl0cdkn6
MJWzH8JBnAO51Av37KNxwdeZuMw4GfLqtTGGJvPzaiy0II9DS/Wftc3zV4jBZLpR
hQPl1Iz1UMukmUsgraoB48cOtPO/e39P9j0GT0ICG0ApO93RGoU28HDMkWcpYDzC
v/4fhlgjEXlH1d/GTPofxLfDZOD4SNWUHbfbNTxUKE80Z4XiU4eZifnDos1yO6JT
saUoOb/87vGLtGkk0xx5TgHV/Jdmy7yeyD1Li0WSQfMYhvg7FrBM+h/JqIwIk/lp
obt++mQqPY7eXMTkfXvjwVhi4DDPnUxOsRNceF8OdM+Zak7aA2FrkAWmNbwV1tAF
D6zr9Zu5ch0aJEdDMeqbIxClv81hYyDvX6N3HzRSq7fmWPy/wSZboqRmp5M/7nFu
7MxpkRHD7AdgBqEguCLVI2M//r8ya0gtaxwW6vjh7CsgL8nd8kj6RlEhNYH0iVoV
kYhT44mPQEM8vcLW3dffxyQV9tZSP/YLM3wZ79OaWYlvGyxHLpYFM9etLOUs0fA5
CmnBNOAcCs7gFChk5vSNQKIZc/xhte+fN8ATvPHdymimaWi+DZqa1d/T+jc9bL8r
wGHcmzoKrhtBP4X+TIxVQmBSBuqy/enpSuQjf3hLd9Gnlc0vwWNvuZt8cOJ6VV9j
KnTHoHFsAvkLlYcnp9Op2wQ4i9qpliUnXpA+PYD+kAZ2IxwL7LqK8m5ru1ZV1kIp
5CkWgeerl4KmLD3gcFyqVE+yFc0x8MC0rdeG/Jsnvf6+qRecl6jdql8lUYmZ8MDV
W5DOks03Wq6nuRIFSratsNsGkCneMGyBQyB9F494pX+fJmzsRd8jqQnLfi58miS2
99k/akz8aecJYwHAJFTXLZsbAWG98IsrwzmZTnV5sQLVHPIkoPk8JtvlFMMVFucL
Wla1AFVoOvLV5oFyEuhdfJC+UCVdvCSVb5Hinns1SVcof3/8uYfEGzFNNTifn4C/
9M94lEZHZwr5vynUNyp3La2q/UKWWd88SKXpJ7IVekllUbft9YkYjMuQCV8XXPay
h4sC7N/zeAonm3XpCsS0CvtZCPyNQBWkrvy4GJkwfMDDC4IGsHPKrBGRvgfiURIM
U4uRQH39+9YmVHzmnTcUXecekaQtF1DR3i0vBEkau00lSbmbjSFpLiG+Gq+Wsawx
SmnepL6tseua0WQjv9pGrdPSKTb19bMbaThRUdX48QU/8bKU3MKgRKec3OiwxTdv
SHMJt7QIrHOs6p+pff2V51mYzJN1OvZp70QTVYzrTXdRp3HhfTqfQANKtj6Dkov/
IJpXXYE48wJ11F8lSkr30WYdtBnnwSIsm8rCwJOm8DGZxxTbu35hc29NRuCc+1mx
cbpb/KkGF6SRiCR5v4Ul79zwFhc7+Wi1BCy94Ga9gJFKLZIhiuyvDsmys8Hp+SEE
MrNUUWeOMA38nUmJSPfDOZiGmpQemDE/qs0oIGuewt+6ewQx3xMyU66T2V4qqH2p
dE8wVy/gt2CD9agy+giPysd1wd/80voN6uMb93PyAU97/FPZx9ldcMVDwtdaqmFN
1G5R1r7VxUQn3/rBNJe5E6STYLFus16q6AdggPPWtM3b8cbE2bLYeI4YkHH90GXd
cYImLEcehJWqad+WoQhH5POm+KYmsLIR/OVEIO3jPlPzLkfgaFmqjlJmoWrvKxEL
ENd+0SMFV+1d6kUpo3FXJlAka7vQDlNhEKf8r8TrVVCLSg7dwt3UHnt2c24GaRM7
p2UOq3kfb0Tz+HOaf6YCzf4MqZ0PXyBbHqUAb4wl2jDRv+VD+AfEEyARvTWMQu2I
T3V9nZPnpGSPSqGYts60t3FxDxKXc9Pu+RDVwotfOADHmRaZ4zsza36wlRvXXZwS
2IrzdAV3bjAXD7lTL27jqCSDu9GIofJybGz4IzgaCjmDDcbG2obM2s+R2yyPqKTS
JNCOOG/pWkx0OYXauGdT1/jnoRUNdCwUa49gFBlr9RxKCCv/+iIpNarwwLFYuqDl
yCyxVqGu2YntrJqIxIozyBDQxF/2oAs7OjXGSh8UFtMTV+gD6MZwDC1mZK8+lM4/
0Td30auWLhVaxiBoikACd0JDTMQGu7gmhNHiJkXEpL8DSLx352JPYTS7BusuR5Fs
h9Gw8I63LQ1w8UomQZuDqr8k7CGTaTiXuEIbcmp4Mwyb7pFQb7ch5o8uwkrMYwpS
FFX39xxY1Gp6gz2sVqPR+8fai7fyaJwwGC9/D3ry4HoHQsCs/0aWTrRuhupd+1S9
BTqylUVG7S/T7bsTwTuvjKQVzUI5tk/HlyX2crkI4CE+On6m97FDvp8+fVo95fxl
gQeZxQk4bavX51i76g1K0d0MPIFsAW9+viIrqAQcIQ0a6y11nzw1zvPUE/x6XvkP
0EkCnxDzzOoNDj3Lt6tTXMvhMnz6yBGJjQSTE/zjiRcwHq4qtskjS3r2q+3kueFE
IRqzNVMtuAqXckLra7Bi45pXvaxxaSv4Ngbohy5j3Ltz22bOFNezuncTEzstRMOP
0RuBcQp+kif3Pw/n/v0PUz9TJhF5pmgj3QdiJPLTkri82PKRTcn1eXRDZLkMgOUF
AmzUyJKaAwoZEW0hc2/yASdioZf3Vpx2vJThI4HerKp2Pi711LRfOpStQxHBXcni
mQLNfrdfjbassW5qkoN4URuhH51WLRogxsJev9L3o6AltQD+XKrAgkxDf18A6GeP
R5brs7VYhCwcTINaVhRuTKCbi6H/0c2Af9554ys3j8oENYNS6dpAITgbupenb7lc
e8EMz2LB4f89A+pzjZ7ax4/h3iVMoE8eI8d/VwiHK1zFlxIG7r7H0raMdUUM42QL
ZhFoTZe3Ms1XoP9B/Jwm3uKTD2KGZSltyny3CxA3EtlSigaaniCkHK2baQa46tBi
1HqK69sP8x4JLD3UCy9sCeZE+fJfdP1UaCT7P3f2YfP/aSRu0wJsi8zwNaRj+ogf
o2GbiyMbG8FM0Jau5G+ay3zrEzWbO1nTWvG7gUMxHyk/lCfYVzcMbWHyHKZNyH4U
CgmbxG5wHSAjuY4wqN+VGpAwCer3TN859UTlc7mMJXPT8ZyZRMcezEr7Yx4tjL3c
A5ObFISTNsN/5VCUDXqzB6HisltFYuPNnCZw02EqWA0myQzpeobVbWxZgiXLQyj9
bYksU3WLIuDzN5RyRy6GB9ex+1mXleEqjYXbxXnZc0iY7utiSbJQBqpNIvnCpBao
ZirFLP+f1C9owP1A6sPO0x4Jo+f+8ZpnsHtuqVGGFKNVjOCUcNscNxSNKGejLg2p
xGY5Dc1QZH4BJIIzotue7Sa4I4KYoDgkAQyDiNbFQdvMX32BDpJ5vIFCCQNB66e/
59r2E85t+0ZTQqFvlmHcmgPrAG0LpV5fSFPuC/3q9eBEXhnbd/JhbmahOW/zF3k/
zp7dtBPjBM06UfTaNLpkumL2EfYf37b0rYnEgvbst8Eoe9LwkzZ5MIQZW7clnh3e
a1FDTR26bfAN6IQbrBLy5j5dvg2eHP1APzzomURhabgiy380+XJUDsvhUhYnpEDC
N44lK3hX59HAVEeKkF7dmqMdljrhiBozYuwU5bmwZ+CnT5QtfHBfbbjTjW5YE2z4
ezntLM06AXEAbOtdPblNQ+QI0TXrFtofBUkJsFqt/XsbqDMq2UlgBtA7rs39KnKe
f8rXD3LLz9gLTDoosVcWzNQJofaogothGJnmTBRiUkr5ZR5U+uHq+emVYP8MGilH
guhcBdbUs61pTGmtX9e7fgHGsqWV4o9LnwFq4bUpksx5gzzZhV/uIhZIH30dqNOV
Kecw1AijLfaRMmnQUC8V+3P37Zc5aCzDNYX4m9ILYxXABnQHWBGXNzfpck+VnWoF
uEowkTXa+9GVPza0z0zRiR3bjvjxsVYHf02wU7onwU3CB+okGJNo92qT0x6Ux0df
rBr9gk9J2Zn9gqd6bahFanc7UU8AYoR8rw9soXCDRx2hjB5EKKKSr6h3LrwS+3pe
298lRg2VsmwKAGA4K8e3NUVrKEle+ookdrQZJIR0+B4lNUYZa9zxbI6zMb6Utazr
/JYd/aFbyPRNevZoA5y/AW0dULfE+wSXSrXXyenPyPCmBuE36mki7QwdG4z4BKnY
Jn84oFbAjYxRVoV+JRLvFLLXYrT/qS82RmISAl1Pcmv29bGCtvHXSB2UKTQue1nB
NYx+PAE55WWn/0TAMK9fDxWOW821LJpalohakRBY93zjvivVmpAPKp49GRP3wtLz
dqzlGqz5pHchmtBgR5iRHqi9ll/jFhThetJsc1wSrHwG3haKtsA2sgiY8WjAKy++
gHZnk/+hdqvCSHR9R9n4hisZb7QraOH5RPjF2KydEJNerZZqPYh8uFDYCKnf3p0X
Y61lmRnAEvG/6LyO6f5JGp7t8jN40Xz9fvnfS9cQNtyOJ35mN8Tbs7RKfsDzrTr8
IxG69CxzP06YTvoeUhn+MXWolJaaO46djqKENG1e8IBdkcek5jPFm3Se2neKSkXa
6ORZZiZD57aOcotLGw/KpqzPK/Bu6+DbW57N63ira7J5GrJ8JJOQNSOQdStKCAXi
rxKwGJkg25EGmJ+f8vXbDYqQe72zMafUNXe/jt77OkwBmYC6wf0mxNyWT9b28WSm
qzc7rLHOOsKDooHvajWgYGi5jXX74axB2K4pGYLY9KaUwqPbgdTwxUmYw9/WzxeJ
pxu+vPIPLKTlN7jlFlm7uPKnoMmtUScd971861p6qdUzvARXGOmK3FaoIdz1fkmr
TExDItLRldK+zGfAcQSyvuz5EQdrpWmFc6PZUmUTE0NgQJiz2IPQXepT9UMJhLGv
MX4GhD7Ca4NN22LOP/S+6k08zruIYTndKlZ0Vw+QqM5JQ7NQIWhNh5WdPjZj/+TU
Cj7lBTM+CbEv+lpvv7ERaTiIxiSwp/l6w2rwZIEtDebn6AUnF41M7PF9aVuF4ziD
yVbhI3ZMgb2xgns4/nLDAWbG9ypMh7e1VNyQC1wuEXX/n/X9SWOuVUDV7HSfDOJK
eaXdfzPO03Yk2H/aUOZud/BRJmzxlxaMJvrKSz0nuHpq9jS3+wB+Ytz+ovC4J0gn
j+RvaNHLUqfKeIsWLFjZRH1TPhhF9YiY+Zb9tCLP+DCQT4bSDpTN3sOJiWVdm7Ub
u0z+BSaI3/KZ0h3sWtqjtPSDfn2QBUecN3r3Flx6VziBzvZFVWt3zCBqxAu6N4YS
qAw9BesMr6+MaNlivNz7U3HoNw4Nv689a/LRTEG8XXnWLoOnvrz46OLyPRce5d3n
RBse55y5Ccd4C4OC7zALTuCMqkmvBtvLUKcKcqne2XSbAkDfiZmLeqdFWFwcgNih
JRoYxMhBJZen1bDoLZ902rUIufMBxT8qeydt5yLG0EijvbEdrWMXicIuVvVe60x0
nwiJURxMzwXLEKqW53gVpLW8btG/UWzN0DnBUk6wdkiEHKkNqRmQasz9ZlcnmcP+
dz76H9vQaCMkYcttaXnIG5FKDkUoIqwsavtUjOSEzkukrlL1+w2i4pEPT+eX4gMr
aMg/vXg2YEmTR9imN0yVafe+smGJ0M0ztv8qKEDgVgskilnUv9X8TSfF3YHCvzFw
au0su/2QeCBm9H0VyO9O/8dXqNGWXsJAZBosJ2A1YTTb0nTc4sHP3RPNceFXWieK
LKKTwfgSHciQoDBvi9BCh1DyJW1KQN+BEM8Z/i4O6MT53HzPhk+ZlpABJ836QmVU
GYmqfwGsSLDMIP4fSiOtQaEQzveCXYwtmmHNAYBlmMV2TKWq12NWxUlfRhHZfYZz
yqTp2d9MT9Hy/of0ZSDLPsMDOFsKxNyDgGjIkBFsT5IEYxZsKQISH6TX1XobwqDf
GNZXwkpuL5pFMaq/zEg+0+CzWv2mBLuburK+kuYUNzcTAHx7LHb+JeSkwji0nQMH
QNNnMOENTtfGdrUZvF6NhijGISMeQTk2eVApDiPwDiqo8FbdZj7lIX1sNOugJ+/0
2+VUD6UBjVwWLaaUcgNxGnx9WsX1HlQlg7JWQKhg0A5kvNMoU3uNdA/0N4c9Bl9R
ERpW/szbfcQufsyKScN4ayhkQJhktGWBEtF0kw8y+Q0l9st5GW2hkgs3FzO04pGY
VjbEABalgWXXqHgS2Oj2NQjgPkqtxJuVd50RKA13BSFcGxdv91HpT4xvymXcR4yl
vHWxBtXHkCLaQkmCrJh2XdqIpNTZBrDcsG6E+L5W1nxccmUAjNxBpyGJcr52OMvq
kowFDmXNCYMglsrlKmnPQrQcgdQekalTTzGH8Xm8ZiLZ9BZRH3NER8DqAdMlybRQ
jt5g5dqj6gkgbaF0mMav1+wg7FuUjdihW8YsdaGT/whyEgOIxGFxRa50H78C5pQj
zYorMnEtS/wmf8zVmnMDPNiSFpQZdD6TD1vX1LB3njTdM+vNdhmVSZCENOO7QMkU
ZrDUj4pfIwVR9MxxIpNjEIQFjlnHLK8OBHHBqvEDCaByclISXoHyXUZbFYJk+iaU
E0AEtfRF8xfEgwXGfnNAVe9XMsHm5kRHVf7NOm19wHhLsI/a6J1WNYGs6q4RRRev
zLpUjxOkeNYNf99ZjcYcnryU6rZvYxfA1OGwzTr3VMxtaajyPVKWw2GQxfGShJPv
20IEFVE/pzKLi3X7nOwB/dpMruiV8Du9ZJ14d5VcFnPOPmWKwF7Xdv+B3wjIEua9
C/DhbxOnd0xnbFNu/OtYhnsOOuiN3bgjwIPIPTw9k9Xmnlj9nBCAkydxQDGuJ4ov
3g0OzAgbOsv2vRK+FzvwaH1YrUMTHNCBfRzTixBWHOR1rifNHfqpbCJQOGFi/xr2
ppUXClBqAUpMwc44sjDaQcWXiACb2uc+vDBeAC39bfqZaq9P/s/C8zG3ylLj9hr/
tBrZNb1+10/kdY/SwIBLJH5P2+cZb6efGsPjPZRTq2ls+O+6gHoUpVv1R/5aEFgP
q/iF9/c2+5yPWxe2q7MQFy8+p/Nnn/Zflgb4ejRSDxbxDQgJNBi7mJeUJU/H29+g
Q9c/SCerjGDSAnLo0x4dqtWF8cxUMMfDo0LkS9/vytHXcJnHO7EBS5F/HozjlHD0
8JDXpSXKdenb8XcnTqg2X/ds6TbSsy4W5dfBRpnC6vjxa3ynIwdnzVvDGcjpoLge
5Bt7Vys68eqwFsutRVQy/5O9gWUARbXiXQlCw40IKgtq46zqh2Mlhu7sO/HKA1yX
FwmTCxAVUDDRzwzVnXpPvrGV2nTYrXa09hUXuPNakyBwAtuf/K+AROMlPjVKX+mT
EXR32ub+3vSz5cDM0TMrrwVyTb9F5H60Gr/4V1M3at1ynEr8GyHzaVrnsF2lHtmZ
svMfKr4/g0Wc5Or/Nh9nSDwSWaK2zv0WS0fgn+23DlPlZykjoFypM1g8ywK+cXk+
0R1O3sXwEixIKyclDvPPnO52S+03z+vUBOy+E1IqyrmmTawvr7W8pmdZx8GnrUHf
POiHVZY4ZgtKrO340n/L0Yxq5vpIloL3wcVNInEEiIrejueWjMZPgEKAZ9qUi15h
aiUWft/OJNZ5GzNWHHZmzPxJg6dZOdQ5Oj3OqiIsxBnNGZtwBbixTb8fi9iAeHHY
Rs7Xvd0gNPnvj2n4tJCOPz5AXidrlMzuGTcRu1Uyila1spkpXLpNnSwj6QbfDDNG
axDWN8ztKk5LudsuaNmwgteWX9usOK3iERXxVgdRe5CoJ2f82szUBJFWW+kXwJy5
FsoHClMS0BQKJnMuWl8xOhXjptRaVJNyj3jv2EVY7nVDtRoV+JWXlTBqS3LB8N5p
j2LsLh3r/vvc50dq3Ux41o5Gk6sM1iMKbFbPZfBQ392PYiBNU4RHY6lD3nAvs2P+
ssv1Y3AbHptEDKUpZH982OCbKiUaBdVFKt6uNsi6/gHB4JdlFVRvn9m/m18B14wJ
EBU1MDRWw5zPqyLO0SqGYIrNy8X7jGEjovGQjJJulRBR2SHmJeejZ/MsUwlyTo4r
eMzijRnvmsxny2C2vdNHIJguC46kDk+1ina9eReIbqESh3GB0v67Uwqd636nMNfk
59GuPv/XDtpbJkdNkh1sgNv+2AbTLcJkIui+khS8CVbsqqZfb/7ymfjddMBhDahZ
l+YUO2eeenN7lBEsO7xZS46jnQH9iwiHE5TuBiVNNoBiNtS3KsJoZ9C6KNuwGknG
VaMTpt/Q1W5QXTWGksOfg7UHOqjTBqRdXWBBbYdey1mRT90PjzwGduxUqTrZrLlR
4BX3jOlhStIRppZstlYcOhAk7mJ7lz8RqYEE07y6QEBXMe7tgcugiUW7Ljcsu41X
KW6jz4AbmNbTcHwVlePrCgHfD0mufNyS+PO6uPefrPTR1WFtixnQYUpTryj4Bobx
WythB0mxgLcuT++deSCL0Dff7gQSvxcvCqWW5ZV4zCcaxC0nZJxwJsuIRxEd4VrK
RAhBecrrDgMbFR0vRtp3v9Ndo6peJJroTGz6zwoG7gGgnUU7vFCCpTthEy286Iza
1CN+fN4DPtIhczAOAXJ8IfTLBAhtA8QO9df4b5eH5BehuMt20xf/47w7Hl4dPn9t
5yZpJNyEQO25k9Nei/VETZp1HiAHTvk181m+dfsJtYkI71Gndpl9Wu3FEmO6QNAh
3tuoksTTyNcEaFpkyb2e1e3zxDKAhnRVQIPIeAawbO5ALTmOho6q6rcLnRmfnZoo
sHBH77ETQ/DYnNX0gOxNOzYoMWtyvosGv41zcqocGCtbQEazJWR7FxFeytQ/aM8x
b1tpZwTcGFB7GiSQz8vA6b14Oxmp5AmPU3KBHFgUgqHyMGbXK1HcDjmKrF+psVY5
5yAwp1ZdE0PcrtAgS0QfJOrS8MZYk872dw+OlKd4GMUfvdldDNWUn20c0tydwzzy
GsAI8Dn1PG8FmoRMebrzNmdQAsvJTmP0iqGhYsgg8PJMejDRZjhpXFZPxHKR5vSg
2GgZcDhIkeTSXKFZnD5WxBjDnrtfkBq/WhrSDIM/eakZ7mpMl2dFJTgH2fE6W1bS
vQebg4+FAEHuVBubHlk6ne8TkHwmF02Sj2GHClxgEKGY2R7NGGhycMiNKQ2sac4G
mkfOTmbySXx6gW9ZWli6LxhSfU6/2A92Ph80QG7ovCxkM+vAu9QYboua0PL5vMen
pksvPcJkNkYB2zvLg3t/4jzgopJp7m23oT6EjOI86Z6VffNP6AS011Y11Js0GSGP
zcup1s3ksOtrVedEy9zZAsjgLVT7q/kPt0HtnLKtPc2+fI3aKuI3XVsh2vBUN4gr
q7GCNm3AZdXoq0eIzL0h/mgY7GSM1PYVSLpupl+5zc61o5cxmJOvcDf7gn8Kv7Gh
cQj0HsU/QZXbnYnwDFUPHeBIgNx89rEQo+idim0H+ZSoPdI4zlmD4PIVmu8VL8Cg
Q4bH1FqkMuba7DJO2iLL/7D3aRfpeoPquo7SqpMB7RgwPDCem3JUCLhKzPerXtSU
BlW3RCqOwJroEeb9sJcZHlfw5Bh/Z/uCJZuF52SNker+MJSw8o2UGo/5ZgLX235Y
UTBwUnsIw06uc/JAPGordNDJbrKDxlqF91z9C8gUIxPOXfR+4EZb2hiQ7T0o63bm
yccfA+Ps+NJauVIPNuStpn7GDAcVoRWxxbM1/PDsO5REA38+xx05NqbTx0GazSl4
oDhlUYVgVHvs+r4VRTswxvtO6akGEaHLywYjzPF5DzcQq2Nz1PbqfaIMn/+RcDk+
d/6bMMO6durzRjJ3JJ76eAaySPVN3ZiwMgcthrFXF63WxnPltPeDPpolav8F5cri
7rcFgTvhfIfTMJw9ZeqRc6hzxkOp1ITX9sZQp3E2lixsAXS8NLGIgcc9Q4pGaJGJ
GEQwOrf8+mdXGoei9OjqmX9jy3I3qpVckVKwZrwSPh2V68LtFBYQgLvQ/Ac4mxSJ
oyp1ZW6KMBSDF9A7+JGN4ealc0170uSU6JXFSX40GUDe6NF5hJzEdSQwnDWgoTq6
zWc6cNAP30/hIgyS2r+jMIuk9Ulr53UkKX6fAeA+NZ9JghWUt2agKyGWkYXE0RkG
ZySzMMUkb/ge4uq60INPC2tMPwgl6XU+fAWqh+6MmXpK7HyBXBJ82kIM4T0AlI6J
xnxjrwTRyr9rcUG4IY7aMsdDeyn3U2lcPRd8leYIojGeiO3jbJ3A0DV6txl/owC0
iPLnEKXpPVdcgeytGVUpaWx76O1bJ/5w7moX4/cjYVa6dQSuKDxlXqc4Y3tVZ/AF
0KJX3lVHedTV67LDurFRAhxUlCe1t48LyWMioPq7h7IKgptdvleVL1OAnOMMH+sd
hoKzCpSdLJB1fwaFL2HUJ9qBq+JdKbik14PUM1rmT59RhXOUAP/oEIVp6Y6Zrjfu
F/yiZrrusJw5wPv+oKelx/mDZWh726bTSiPF/mNWWugKdxA+YQi+fZkUsKQynbpc
YqSzQ+PWeOcZTW6ZFVYkZZ2/Yn0vFLvZb7aG1/+YfMZYD978ueVYVTIYSAfGITYG
2UYiKhhldkmrJOwxeEGWXRWGkmHIJjHXnz2RTQ3EHqnnhvVy4+uWI8xxqr/5aH2C
vIAPEN/c2xrpRCp8or/PwU7VYPsx+qjRxGdTIxrlvYU5Ep8fgeRf0QQAf2IpuMXq
ziu6QBLC40IP2EOFH5Z4JBaGXJjASdwTLKLM5bSBaptectvnIXhnJf8S1s5ICsMN
bxa/w2pLJIp/YXy/Cr5x1GQu2bh/oZ2ALp2VUO57sW/9UDnmw/D4DsJnLjUR8zto
930jwXiw/vs7TyQdMhngnoDH7Y6nkVcP7oPhUqJK4P3XwWbqrJpfp0J6SiPc+aWW
trFQlxac34CJP/1qK1GU5aRCHP6BGCirslJPq4lIsdFRhb/Qs5YQxUtRI/3sjfrW
8FEaCFtFUaKwdjbr29JfP6sObMORpIu75tXBP2x8OvIZVPTRmCZsjSfcaNnUfz5A
IidCbXbpvT81HArIKOR9JkevjEEwp6DF/HNXPjX/kNBiq7OWfDMK8CZrOojakZoN
ds/qU/Qr5ayAWZBJC0yrcznPofvmA6g4+Z+jDWRWhBUZBioqlC1fpEImODOYX6zO
2NCvYw0tcLnXZ8g0wGG53gxkJYhbQFk6HN5MZ4b3mX5i4mFflRMf6VwvMDoDKzja
d03c9bvL8YYheSqY8/q69TZaE58dXOpq5w/JMaTkMMmiDle6HiyPOhth1qMMmDoF
/hELQnYLgkxminUiSV0fMzmQT1CKHbuiuAhdgAErW1I71nJDZRgUIp43Msk/7OBi
TcCIPwkUFkm1BSH7P71R6M4pKTgCAqx8zajV71zCPSUYvjWNWX/v894VD21npYab
SEQ6VbGNLxObHVzINLZHmC3LN8qxpv03iri9RJ7PWH7++tRuFRinu/uNSndYiSkS
SqnOlfemsAcCzgGtXcHOkfc2/5TuAZ1ncJ5BRy97TrIb53bn6nB0k6pNahr2n2To
ChcHOgzRosm4+tnPtcBkDMGiCGI+ZGeiJeFVzZXwONPobgzPVr6yvmdPwPC6j/87
rO4+Fw8CWNcuSGavH4K6vsjfp+VI+kU2Laqm8TIT1FrGih6NhVFQVE8FnxNKtRxB
I/Ix7gBUy8UmNLg9Eqh5OUo63SwEa2k/bBAYUMLQUhUKqoWSrAoP5u7WtXb+XoNs
tr9HULjXzTi5w0gAJei2x1l0tSdSg9tLfySNownbMdFt/372cEp4BqbtoNsNM0+y
HC7NFxQ9yMn41iqRx/I2ADTQc41WiiSJ5O2WoGRFS5+pYebt6XGInvqNgVuisiyM
3ZC5/r7FOxBIPDm1gWKU9Yu3V6goVzCvn3rhhgtQFcepDUwwuFFY8Ne3Z+cgWnBo
ePlZsfQqfvE+TEvu+jJBdnSWCZ4nSKfBTzyu3dzIjeT0SgDpdUFc9VIPDX/ED2mm
yh9ubft5q2QkhJm27gD+Aao4oAkMlpCn9QvKX4Q6nP5dXfFGMpFdbmVAmZlOn6Un
UpsMLp/N75uowWmN1xqkBUgGX81JBg/mpDOEGNehjMJsSfNMnsCAowJ/rivaO+OB
F3AeAS8LyFX1yH27tawiuDssTSzafCsN8AodQ+YnRQ1V6l5Z2SbEkLpN3mj6sN3c
K9m837hb5m/pvTKR/XCTU0F3d/DdBCWcRQB98GUAzwLECDzTiAYsjnSU+QxgP1xG
22L0skPZ9TN2Nbf2dfC/26ljGymHB0QIfEgBPzpllOyRUnOg0ZLKiaxaqBXy8BEv
CQrZ0lLC8IR5xYGT80Q57eq3t6GBSJKCWPm392X13NX+lzXvZYygTQvoB6vMypE+
TvkDiaDFaEtKklpGqQ+9bp81jCnDTkstJksdX/LaLcBYI4NQ7J55ceO9PwN3+xyc
gWD0dzo9Ml5sZIDxKPuBeFfb9EQ4KDLjtzfM4dzUsmOHQ+hWF8KI+7OueeAQonbt
UHZjB2NmQxMkY5bpykLugSJbSdB8La3poWkIrwzdSfiRFsk+j8za7EA69fgV3uL3
9+vq537NMDs0K+P8LJLnvmkvhyXhg1IbC5dw9r8zPuB7XN5ff1jGLrCBmnZjtMRO
vHRbf2RpzzeP3JFO/vfUgpIbtp4B/0H4mDVCSd2ySr9iO5EpC+Gw89HvycHxPmmJ
tcSsXgYIqGJufp5K7/uaun/w3DAz0ufBLpBSlxvUkLTzlDjyJjyUQt3xCgzeTnyG
kIxPsryQbcktBeKdCbQk4ZW6JzBeqfiGuW4EcHXxamHwYKM5kKY2h6IUVrlKT9vD
Jv2O0yUG9tvpwuXKaarJlApV2i0sClWMCvFqHW7uvsNsWOghmOCZarVSGNrb4zph
Q29t24Tj0DjIdye2q3y8d3SyKT+i865eAdJ+91+9S4XNaa4WEgPDptW/uEBGY9Rc
UQIEpj++Znr5VfdJLkHss1oVqzKdJOaM3FhujZ+ccEDMu1/noELTjI0U06xnhTbB
CUREyOjqNhXnaL2xX08OlTwno+vRThpBt8dMS8cwN2n1s0EIxo5bQpvttuB7NNNS
YB3KEdYucOL65LkjRuag46s0QtWuavBGfGveFnFFh6yyhRTnzf/nZO8+zUlcnd6m
KqY50WN9gAuaVr1FNkv7apZejXBX/30X19HRayrM3G5wKbJ7InUQp29KCDwTw3PO
pv7o/my09yB7FMt4/F0kDXHqpI+42RBPGM1Te4K6aKwkcEkrurLCyWZaqkMaU2s3
xwuxu0I6n2xuPxvn6uCLvAEQ9xocdLyJ2u4uDAigrwtgwcQafvoVJHOqN62aa6ou
cZSSxLBg9U6fE9ZMMGxYShyLFN4AlKXX9YkYrMkUGmP24J/+k9M55x7xYMdaG4g4
UVelD6FzE07IraYVK5gQnWwTTxDUVZs6nLsjdmbOTiSieLZQT/9LTDvQ6ZyvAxuZ
CUWFUHYL1LnvkuOhk4SUHF/kisvwAJU9XJsk1GGSS3D9RlC5BKF2pfRS6P/dNvvi
kN5RVWOaXbYhft5mLWTTX//NlHAPbkQuhidTu5tS1aXe+pu12SVtE7NM6QECSdPs
jgNkybJtFrgF+Xw1mAGia38NAUZx1pvyYEE6e4sUVMGG0HkORwZ00k1aWep+5bgQ
MweEEA3/wgbMkKRGpEvogGTKxkRTwAJVdHsVLKUXtGSvkebbjcVf4FV89nHJIpV6
i7kGNEHyvVqn/MV9XEFRJ2Dp1It3XGFhNobLIbCvm4sUx0jHVGEMwmmSxyAhyyy8
GjrDdzzBPOR/0gv6K/Lz7yYvMEo7ObXVmuaZ6tmLcIlMi0c1ojiq46VTw0Zsd/3i
CG7mk7Ipy4lCOMmBK+e8VJDK6CvQ8d28uFrrhiNqfjTO70BaS6bE/q3PZ5Jr+rp2
ELh4aLW24XlmBq7E/CAalAOdHvTdH29c95jfr0y0JO/RJDaypi2W8IgbLq5nd5Kb
zegOu+ldm3gxh1icVnBYEMcMKdfDz52RsWhFlSinpmnEpQQaBfCcq+4rE2OPoPuO
QkOAxXe6zrVlxOviQAB0tgepwfko9GrP2H/hUO6hX4Fc+eeNn4Ke2SnjbHwLM8LY
iAsYAYCEFA56XNwtf+MUZ4A4RbEgLKgm+Vsm8r4IBiXp0MIfrW2fn5N6pbTDPwLr
qsRXXpMtJxUrei3eCIge1R+XUq/x+xPnE5AYPVWn5Errqi5j+eMuA81kzP4Az9AQ
9TKU5V2sTsp9lUnB26Ocju5TScYVazhI4e351BG6+xt3FZ2H5QEP6ElZvkurGM0v
GVk8IDgafKOrKdYPATeHKR9DiFqMsY9xM5Ju0k0KHmcSxi89SQ8WPSRG1Uq1Q3RF
DEVY8hA8PRXFrx6lDbvsW0RYLtqLKkv868y2RxGz4RTh7rFoxQ3XpScu8ihRgI9+
O3BhZ6pAoI0Uz4kPCenHWrW6SQHTMSTLXrIDmeL4ShKLMnh0Yw8s6O+aIsfpr0tB
k7zfjFMrJpjWjAKmypX59ObPCULdMu72ul/uVTBwBkk2ks+u07brmK/xXES8VFNm
3rrZAcXCAOnNJT6Q6+9enNjBjEsxCnVUDt7a8MmPapCSCDish9Wi8xwXPr8cQV92
AhiDJdNaRryNw3b5cN4zRO0EmQqcPaCfufSqhB9NnvU2cCHTz2xybGl/jmu+u2qc
WCr4QIguqPTYgAtb+LykBsCE6NMflroBZWBwGheBlk6Tqq+thMJarPYdlI52JWIk
su27hsEZfwL4P8z+7bNcYFyX5DUB+/0rISH5lSBwtLcaOwILnbt2J3Z/mXbHs8cR
8lL5YcApUXU0cyjlDo5aZNoAR3KSNsQiazPyQlSA6v4GHBCKVMW08fSX6lf27fA3
PxTYXA51exN9f8qOAhnu7keR0embyCpuTlVY3cZNM5Ku8Tm+KX8LvkmawK2/s+dB
oGdJUQawahNUwoBVONjNuCHzTUDjk1YUO5izkZKGU0QiPu32BtP2MuIXPHgpK8g1
QwKwwFm28NFx75oMkoKKVe7QyT0DHwGBvYV+CpfN5C6U3oTXZPJcv3agSALQnnuC
MjDOb/xVF57aBKjhkcXGfgcBw+zO1pGODU2k60Wv1VEgvZxghv7NpIXknUl+XvAT
H8Rm9N0QC+6ZTDu+aYJZ871qAK295VYTEOnd4U7+XcaTidlOmaX1CnO6RVCbL+3H
+aUua6s1sAnJCxqCOq1mqU8k9kvgwT2jlEausmMKb8VETXAGoHlWtMomcsrBdKoA
elOsRlwsSDM8EuY1wlAULFlGTavIi+0M/XmGbm8wKE7sk3vUPDyONWjmmWqIXKu8
XeaFiKWumvspqVq1i84pQ0RATupermGbIn83h7CEgY1dGyFyMTC+VyTfLWkFVc0s
v3eU0WlCdEvva4dGdbiZi7Ds0cHikvKUzSGp5OSrf5wLsVLD2wWQhMbTSGmVCwnL
NdVXwQOflc9wXzm2dHx6j3+dqUWlf8zZYlf75sKss0yM+xeYOeI5d++A7IGy4wMM
u1ErukRsZkWY3Q6h3XKW7dHDYehTFhVTrdapQNN3g8YfwAVFTuk0TPITevLBfXSq
JPulOCI1zzGkfNrsKosatyg3eS2uZoFLMdknuBUFZbZCcg/0YiF0FwbCq/DHICWq
OaC5GfuiTGWTLVpVRI6VkpsRPo41q73MVJBKSs6juUQ6+B8ZXTIB8UgCG0zC3zjv
L6PkJMGB6F1A6r0Bduv3JjWqjkpgN0YFlLmJNAUW7ID0ARW/jZczSq7uTQCLkyLZ
BOGh6LlEgr7fyodgY5h2B+vUn/tuiSzLG4OMdc2tWV4DJvePHVC6ddZSc8EkVdLx
SFnNh32Jtm2XUi+DOXmpMkMJfcs62tzcfUdk7b298fKtdfTxBTDbYZnDA0J85ABd
Uf522y9iSEsPdlgkcorOtgAGMVyWqkMYrGAm2e8476LqJTEzx/4WJhkNLAVU47ed
jek8BWL9D5PQYkyKiy/xx9Fi1uxQ5Qq7aqVUzyLlWic3EEwiZPxGP1LngJLiB/TN
YILmqb3deXMt2f4Uy+clbiA9IN6H4VM2LA2r1SsfwJ/Irw2T12nE+8t0eMOin50n
NZfq+6GKCq98hgmm+3H63Tzu3zSfRfRe7HOACoClUXeimy3EuewF5YxCdk2uYXwz
0LkctzHm1tUH9v4OrCqRq56DtegIdUjpF+gMNxJkbTfDHRrBA5/DkJB5paD4ZfEH
8C8CMnWiysZrDdb1XniRWGSW29EIeqml2hRu2Pq0B8Ot/PzXlKP2Y9Q1TZCoU4/Q
+37H3RkXR6yfwMbbBWQZQfV81wh00JXoQbdD+rzCSWL0jvUIFd4AMMGfGM8CY0cp
wFbu98zstWJxCRo8o46ZWznl+rUr2mkauW8fe8IRuWeDJ8lY4fksho+wQXudUaY5
zAEBZv29PJrBac8nbX8YCtfXMMM+vN8U6w+SWNnN/qv+inoF2UTduRB0a5CAEu9M
EOETQsVZKNuOVvowqmhKJ2inqG6AFh7NQ74ln0db/QLU7tdFV4itmzmwe5PFFucs
pL8Y3wf9EA1DJykJC2xlhR4tGBRilrQZcC1L1FB/vrOITHVFI27ONwq6NyO5aYps
OGXk0sUra6td8WUxLVeBqropQNjusgCISQ7oEs0vEQdYN8JNBiKtljE3A75as2fc
WJVlty3Xn3YRK947i76vYZaJJWMOOaKn8kcpsOnfokG+KljGbWQe+nDsQdm+9CXB
Cxmopv53t6YIlnUayrxdMEk5+s8t8vrZ7NDvpolakTT66XkfrAFejDKHFPHagSfT
2+F0kQ9ix14ajlHACSnEylsYFlcN/MWjfG+upJxf4+byUWbDRw9DdvMfjVqKO5z4
QUL0JpW92Pf4KVBOonfhqglQkJt14BlA4bk960gLPhBaePDHbRyJ7R1BI+ycM99F
CRMys2NbmN5zZNalnPhdZfvCCBr5yrZNzV/187U7S2QXdw+/g3avYhQgk1EZlplL
YsT4bf/cIxn2btJ6XHRQ9vSPu7VjttI7mFGSuTyPzodmnpc07aphsVCiT3CWj1KO
hHfDORvs8Mybg0ImwiGgf9akYa0Df40HoxX5WMzn7UgLgfysn18Z6cTK6yGp9Xw3
V7Tc1fEz0ejSWEEgY2Rx7X3803UaEMvdHXWI1GSQZGkolVa+LcyQ/FUDWaV65kJj
zLpwMNgf2cTwrv3Ctl9j69BtYp6emvfpfi9A/lJkJLz9hebHegqecN4IdOk5kwhK
Lhr39m6qPBe4jJaIqW6TOKZegTWU9YIHWOWXZmnEK10W8fAcw+lWA+IWvVcwTnAm
4Y6uOxpA01H+Z7uyl/I5V0D5jPAvMWfabfxX1AAh2F9qtHbYEo3fQLBWHFY61yE+
qzBBwEwUjzpaC70XQa0FOBzZxJY5V6mE5yzCNg4KTHvMg/2ZZNCnMafNPmXYlFKy
Ui0oBLJKgDpxyc+fPtdTghXzQCagdtCgGsxzzOSqPhjKKSqLlY8kzWMejvCGxaiA
ebANuKCrrfFsVyT1befdnTJ+XB0f8b/TQu9IhUvWUHIdcDtYDWoDmg2ZVJr781K2
bZ679K7kt8PM8bQZf+kY8f9udwIbUEWIFUBaA+SWZHcmdr7hWr5/vzh3V8M1fJnC
3x0eEDzj+zA6SKo58VPoSOTRm/H3BDLp3d0jls57aj6VoVtZUvD6Dk96qwlwNZqb
tiDYz5urZTM6mSCtsh50kTdwtHbb30YtnJZDWB78mLcmAt47M7GjgTpb8rfV7SUl
zymAn7L90U0TaMxqcO9nlu9amZuL5E7iD4gKlRpUvqRqu+s7Tyazta0aB/mpOtSf
FOO+bNL33Ybi9Aj1CuhdvRjRck109TIKEKDlTe/Yi3yWeQN54LtW0fjOED9hXiB9
6Aqu1WMWq9TW3Gdu9RGOF/ep3ZbkSS1q68EENwOJPLfiYP+v4begxA8Vtd50eDgv
D0v2U9MFQVboD7aE8QaBvO7Ei+0nkClRW9UjunRmvDI1KDxivv3spxcRAEK7d0FA
Yd1UOAsMP19fBT1b0MrJhFGO9GHxakgFMKiAbHDSeN8+kwN8m32yijJxMtPde0Hg
wgc1phT44fVr5rygfo7R6KkbrGWdNJNdu5RrgDKaG0pXsmhnKC78h7pSUKhKpETD
RfotYxBgeZKic5Vc9a7uiPcxuQhJ3OFxYMxKCNoyVhn1/q+/KqKIEuGjLncdb6jx
25wNvmJ47AkIl7Tjv4X/QSqS246TvbPyZWfdxTeE3csHGFrTHD//806rT3ioOF2Q
B8u+vyMUs9vGZkpmYkPV2m1DZC4Bv7scInRtajlqcCtZHing4SBSj69XJ7/CKr6h
b3zcv8q+QNlE4EM+HoWh1k0sg9Q5+8+z6qDk6w96Ch4Obb79sRiRnn6nfLI9tuDr
9InMGv04wCScaYGbQ7NI0FFZn8yVCtDjT3b6+j411xoN2pzE2E+HjcWWQFbLaLmQ
SE3JxrhkIj7QUArFg1cvUUt3rJugcQvmGtKkluh0p4kjyn5qxUYy3ekHPZw5bLrn
iHko9DtWp/T5D45YiAGTos/OF4BrbCJYECn02sHfsrup6sKrDxV3wyOcHOqyRftH
SlbYLwwkzqSk+dt+Bb9s5K+xVt9hEnkIuFNpFdxynRvBfdCg+jTMLDWHCBragFXj
7j0KExlYdi+54KyPr6Xbd6NqXpznItaWt6BjLLaHFwvPz1zH+vdgYdN0x4dGJdgV
fdAjRfU9yj3AK5FX0kuauWqxK7anITyz6NcZqy5MJcMTCpDI//MHe+cUjkDM6lGT
mQu/DCqabUylv7oHPRrbXY2ymKGyb8ehJ5kfEaqf94fQzMMnbDb8iOllH9o4Z7+V
kQtMF/vP38AWws5Ly7jOcPa0OF756J9ixC2hDUJu/2ND213B0kOi2NvGxvNLzcC1
lIzC2iIoE6g83dUQApiG/7/Tfhmtsjyz7ijqN5qUcoCncxy1hT/8d+iTnm25pJdP
N1KMKshN4BZ3x8Wv9NuErh37o0QHBScmQyj2OX0A2mwHeAmP5HqqgCMzNhOPpN6p
wpHuY2k/3323/F5C2oKprbB3vUiePLf7jb+sXwOrgBve4k0S/0Le7TLGoqcBRZ3b
roCTTdwZbL1pUZ70o79/qsU8A2AE00SNZ4A6BBA0749UZw18PTR5ERTBTOW1oZXT
ALwKRDX9i3osnOj2mi/wNrIgMoDzCE42M+HzeOvo7CoqeFfuAqNLCy/ZBFyOBfdO
4Tzh+7z6I1IND0wlHnNE9Yjgbcu+OBMOgnyV3awq5ANSLR6eGfMJCuITzOS9jPxO
lRlfPILNey6u3T2R6OVuejFjt8LadDH4vcra+PqZvSCnEDPkTzw2hMiCyr+ymheJ
sZyLpo2MgOtX9lrp4+MLuDFuqCqNt8iX0ZQUAEYqUm5wdd2VF9qhYGvJMt12mXnv
TtNn45+DQ9X5QhAXUtLfXgOVJm1AQRPvPw6Mos/j0nh5a25Z24b1TPTFX5LMKEyA
pRHK+pbunA3wsYj6ITklUVEMvgC/kcwCZvy5BGZ8WePYPl2naDXlCour/oqANWY2
dUJSaRLkJOvBWmqKfkBTL/O6goOxEv+7uzAWzMWQO4zyrPse6DyaIZwo53bg6F7E
+zUncNGp2b3Kt22DKh7jm8z/Nq1h6YBm/uvPEj1YLK84BJ08Cl3qNBXPNoNmIYym
KEmZeDFWPUgi9qQXknj1VcU0gg51Pa6NzIX4J6jQ1XIz9I4cJq7vc7RbdZL/0+pi
oBNBcPP6WVgHVMcaVWHqzZ7ZSfRqoLiOuxtTDH6ugXa8pT2IXElMoodx/v6N/xxW
zizK9rbm98eKpsyzRAYU/lTOzaGYn/mzZ713in+pgz8UCQxhWEOwyEgtfbzVYyFD
0I8G9E4I3K5b+W+bpDZLMEbNgkioEJP5DVHn+NIC6pjrVlXU5tdnEcPuA+eaDHI2
WoJaaI9Edm/lKtrkcE/P7dtUN7h+kQlI47vRPUcN17L0fCJgJxXpmfM21B4AuTqn
Q1wjptJq/mZRJzKW6r5dr9t+wEpW8IHZI1CT+0E2hVeCon/Bj/Vx0VbJp+D3EpLC
fi5EmlnjP3zQ4amBa5oBN6z/6RvRc00865RIkqwDFIGCGej04TdzSA/qP5gjZxqk
xdiGWPGmLrcQNIZB9mBRTDg/ygJg2QfX0ckyqeBl9N0qw+YD0qVasaGziEIDiYTq
R6gpnYxtVXMwRdAe/QzNHHUwNNLdq5KXF3t4XoHsQay1tmiJrBYlNrbLHz0HI+lq
9Ka/SdZ2JBDSJecnJsCJOTxYCfGcgdBTRFQlbejQ86/8JZTNWu1jmlSGAr2clvMx
qxOcZPS/TMRUriA8eCmsNtj1M7WGNpjzbDi42NiX0/BiViEr8yrNtWsHx5o5rkxi
PHLExJUKkymoJFIZfQ4MaXuXaumDNCTobaT/ubP0CEEbsUBR8BAbFwiA/rA2ACS5
eKGB5UDPBAorfdr0gOJBXyyc/nvXZEU6g0xsib42r+YRrdwqqK0mcG0crnN6FOf0
PY1H4ne2jNF87fXNuWG9ioS2MbdorkiIurjDIMDydY/KPwtAl2tnmv2Rr/c9eg7t
tGhkAYaTzl3W9RoJouu/UxmmCwS1STS8qm9SE9M7DszRMhe/CVl75Lh878PxAslC
1cOLB+AuXD/l0zZZx1rYnU9FE9p6NRaGgtWwiGWRPkEc5KfCkPO21APsib4GcMnY
Akjfzrnw+1r5BOmdIhxf15xU8oa2tHDG0Nktyobafm1q3Dcma5/PXCCNAFq7ILKM
QL/f7oAxxNUL/yN2tEbXn7x5QOmdJn9SO0vby42cnLAL+QnesqGXeOVmxiJm368o
ixn/zWv/5GqEPc5eB8NJO4kaxx11C6G+HtRIQuveA8g0cvF+x/6NJAfjZnAXwLMu
etU6NVMPTfU3uKrE7mb7G82Xba0TUxS4JmctLZ3SV13cyH7INmXS0IrHbkvqFk5b
7Ps94Bsh7/U+evmqbZy+t53m4e+WZ13hVpx64HEzyW26hj9HcFbsCQCwM4wtCMlv
X51OsRyL91aB+R8Azs1hcxnacFnTHUbfuZAtOQKHjMeLnOwhZE3iQcPdAgW3zQrP
JAvGh2Ko8yWdP/NI2/9JmmmN2nWuR1GJJvMT7fsHFKwYRvSChh2vBTwB2ALhL1UZ
IyIeu0zEsrAN41DmvHjKe98+FQh8WXERGg+Amhl/USBhewh/7agcKXqC3bzUR1YO
byQ2bUkd1MDluzB0pn28je0M+E5pUDd6E9MPnmqgdgEAGJaZvUF+X2xlU/Vn4dkH
9TZhoGPaLCp3N1RkccbOFFAr0PdtUs6TH12ct/7+BTXP0EJ+NfYxaSHePqdcnQPd
mRDSuraUQ8Zoc8kpqmo5McBeSCTkjxFW5uDOIGim1HFgH2hkkDjyQrMI0/JkP9Zg
Df10AlFEl4sNdkxWUH8QqLM12nH480tTs+Fwg72InvpwotGZeMCbvpGqUouocY+8
FJNDG07HYcEn7U+lxnk+r9wZMx6WVCuPRpmBLTAKDaPG7IbKQclVDoERtA+BYsQQ
vK3ky9k3TTZvOk2V2L5FYUOIDtwyUMVz+IcbZzlbeGRW1H7uy4Hyl182R94tkPBY
6J2HekOHQTCA1Z8Tli4M+UAo8iHT5HC3F5kiqJtInN7yj1bqYQ2jzUhEBY+pSpSx
QM3HlakEZcR8WHhARukR1py1kc5bcHlayYjHghvyGVLv1xthSeuh4NPVKyKN59q+
EAspufJnlV6bQ2+9k/Y5HjxgpJmwuH1f4z7SUaj91cA9qpxWq9k4bvXgHh38m3j+
PLc5y2oOd+P4zgzNhj6iRBbjga7rYsYDpOErT6+BShQohbtNhIRUJoAMt38h1QnE
gJVNa+JDcSeFvzcgkTh7PYCro8Rdb8I9Zl+7b6p1zfbxLJrFAIpLScnd3rF2Xc0A
HvU+6+aYNNpBQQfNlzpxXxmTFttFYKNs15Vg5Sovm5gjBn6BJIfq3yuMwPcmccpK
FPbsctfqNpfZtBqkzt+IIE6nre6h2HCXoiP7ZhNUCTI4NmUmeo6qNI2xDS+Nt8Pa
xE5S7JYyCQJD4xr37jl7dSrRRnXhF9SF1W4HlEVqAkz6SjJxvgEPDV5P6Pcw+GsP
BhXVWibK71sQxgyjwWE09buXvhoCnlYDTX6kYlu+N/ospdZVhQ58FXUywjqCetKB
k7dSrChOVQol2mXz0/H/oGzHP+hDICOlFtVac6196VNj1p3CwmAr/RStAr7ded6x
cXlAztANXYFaA64nd5WJQ3SwA1iHFBfUhwABJqpmhDey+37BqicoQvTxIVzx5rIE
nM8OluVTv/7e2T0NJrIF5yWybwDq/XPCWiNQa/kiRX0u4+hAEU2Z4M2qP8SHb7Y4
51I8i6Lrjomv9Obbt+clyN6S1BwRWVv7NhqXw5Fbm+qkuvS1fhXRGsRH4FInjont
PLyi7GUrvdoNDYoszqKYYkKCPKGNVhN6JD+26Ghs640z2fLCBGiRUZFq7u7fPU4V
tdEfhN3s3FRrWiL1eXLzR0rI4fK6WwktR9/mFz5DEKT1ZT0dx5hTgRP4ufqteq/D
viMY7DST504Cv4sKiq0npf5HXqF5oeyW5hsZQMPmqhOF11AC1mqcK8pPqbsMf3kR
K05KroQgNnjuibS0TGPFOaWoHbCQDI2zHmUhvAV2QPmxrCBtiNlKptJVdD3q4X8H
LsNNwlOl+5VEvtVkgV77frP04BZmtq80eTFKcit9d6PtzyVxw83QKySx6xrmt3J8
OdOmpP3TKk/BJELbHArNpKKQnqJ3xOovBR46sUPIUosy1ZO+QjF1e7qIttiMwTz8
lSg4nDeDP1GKqNjoesg3K7mg21nY5cO93MwkcQzd0/Ph0DTf2LKeClRmahjCFrCq
4GDzyyVhpafvGfaDBRDzPNZIDv0LaTxDCIjJKgzJairFHAfkLQ4J/zX/9jB5ecSv
nrY5TPKd+HANKKcAEOSaLtdLnPHC/udU4UZzUXht0Ea5M21Y2hCLTbUsJjCMQ9Mf
zvH8GddianfpwrxOOrtuQIFKM71L1XON3+9PLcsYxFmSsRaA4PPpGR0aFZ/326E9
Ddiq6xgZLROvL7AOn5I2hYZ540jrH7MLo4OTsbuptk8z/HNYYhPl+DBdmt7yxTFs
pqfFALOqS8csdvS4GcpU36ecs24A93aoDjegtXOAciD5gThEmCdKJrvw5Jx6OL2z
NF7UUa96hPccg3VNmTfu7EBne6AS4+zYorog8MragZEyo4/RR/HgTbwaX+sD31CZ
ln0si0xy1CF/6nXVRO1+Zq6mezciquAGhGeUv4nG4Z8RN4jc/ykSPhSBQdOsBZqR
nFd8LiZrP29W/sdaCcibo6SR/rPxC3cof2lwSs15p1caErqGWJ7674DqTApe0ejx
kL4ucT/GpYnezlVq1xL4Bit/03FzqFAv7nGm791zIqj8MoKmG9II8ctEktXDTzKy
sWZ9nRZwA5ZJvKkEU54SwQPhYn356myaREkhoydN96HV7HbJv7PJHTjmzI8lFGzn
iZl5GBLgW6rSsZWDObJj/uw8BSKGAPCHuMCs8qz7UqVwAvm48tMepDDBamqRbFRP
N22DbeIx1FZGMGC5vpzJ9E/133AeWDm9DG1NRV54tDGeX7B4e44G4GKQRRsdARBm
URvsow5KcVKOCydxsDrwY23GAhAIOt/rqk5eq7o5Fg2zwJuxt80MBe69y+Gc/zeH
Nf8jwZD7rhzLbCprw09RAkKOQnJ7utr5A0OYKjcu+oUct6WmdWMHHZYvqRy2qkQ+
PDQS3H49N0CwvxJUK5TCosFSGeK8j/R9snxm0yCXAtzVFdQoN0HBYD2JpT5zcWUo
k5JaAJ4HxKzvjULk89YwgB6Vi58RRmDqpOMRyEThxZmGXXkTlAqwMdOGjKfGNWwU
172FjpMBBtmOt89AMWrStQwOVl1gB1J5ICNNDTC6rm2JFKTp1ok2hj0+myucQzbe
wHR34sDWS5+lh4TymaECL+FFIZ+nFWztLlm/8CmxK0D5ycEio0OspXIXguFfv9xu
/YkP4hKx9biBey0FOttC15U4gO7Lh7l/dUldhjTUIjxy9QosXTbREqe0LFVoQcLY
1mKAFz6/slmHr5TXwK36HcuKdVXVhCU6U3BCZIO9oWdGzf8yoHX2bvqW3E+E9zFb
49f/2cnazBbnTwoj7NJZOiS8dtOGDyyy/QtNNAvDpBSOI/G66XbJxRctJvdgzuYE
NsBshhc1CWCAcvmzhuHOIi+FTZhRGjH1Ht0TGgJxQMMkZG7Qp8k+3UD7IAA+Q1Li
bIfNos/2wtkJyK2ByzVn31yqeHBhcBUyqQeduptYrSXCtceoqDyUOZ5LVrPOH3xG
DSXxoTBr+Lk03VSs00bVTKUUOrR5UzazZYuTu3TyFTZsMdv/RBrZYZNzwpesWYH2
4+3IW66OsmCCg6/MGdXjdAqhxDAmjhaR+9upxhMbuJp4UsS/dwMK9VONZSiX/5Ny
z+caOn5kYxktUJ9SlWyRYX07vcB4KAk97yqf6vDs4KF6Q6PTe5E2opQFw21tJyTD
PP5bhMDVtyQaqyyZildquiA8lTCYDTtCnRlCiWdpDIe3HAzyeUOcnT6yCHte4gWv
yPyL7pzZOMUnl5zcJl9NMmVxgtLVVkZ2/a/5FLKjxTkg33no3evMl0thnbZGYfM2
rGq8wgyDM+hZ/3AnRiQek0wc98xagFv+XMByRhwsW+Us29LrPJYU/017nSq+PxH7
cLbhNMPMcTlQP0CXnEEeA+Oem8c37zCLWj8k3ncwD3hCqt6YrkxSgESb8YlfgpdG
Il1LN5yFarPgUiP4IdKMHoPIvlDblDN0rHE10yt4X2glx7v9lHNd1bR+DNk7mO/s
cCLdEfCXR0z48OvL/h+WSyDJ21e/kl9ZHvsDL7mcnmB+tcIo7/2LqxJq4dmgaQFC
s+v/ZuUZbTW+hzPDGYXJf8y27UEBUGEzQ2YwHdgtPKeuk+q3eBrRTAC6oifTxTBv
tUy/9Mh5vtovp2Xc8zfMcRiM6FUezlcYF3D5v+Y3zsBJTt7bZ+6IE4uUpvJPwWzm
LeSQYLRgpKrltMxX/mvLfuZAxR080AP+fCX1jjDmnt3IPtou0ZKdxvCP92uSqEzj
i6T50KQZN2ma1nqQ+ef1NKhaA5YscMXI/TwA3atuzWyD0HAbfnW13mmbSw/gOE9P
9oNWK0f2/0z479YQDgSe4t2lUbHDqeq9n8yyvwOxF3EkvnRXzGznStuPOnoH56ID
6PNiHUfJ3GUz8MApFcnotN6M9HA4clsRg+IeQ1aHc5eCfezZOkiOPTAI9ZDwl1Qv
Qkk55RA3F7uPksdKi3261+HREzgETLjGy0bbhae8jtuNBZCMxgTY3ygDyTfPqz38
cz/iTmLNtxQh0DQ9jF2oV4j4Am4y1vicAvzZ3YRd5hKn2Y9cUGN8maF8J+I5uxeV
E0e1DfnhCNV0E6t1sW2gGy+wWG1uR5NslFi6byelTbNx5aSg9oUFyiiJshHDnZmL
WyB8DAwJrecUrzBEQdBzClVoOx5PTAEreb/P3WjbF9UdecxZDAK9Lt2GvyA8RTjv
t1E1w+vwaet+LVlwFDWlzz/4xNk2273hhGwSyuLecxcv//zT57juey4aehm0IV0P
dc2iOkaLEmqTXYQAcIvdfbqqRcw0dQsSfqp9vyCO6JBLXhI6sw1E3dPcAf4Ygk25
m0QqRUDZNS5VqOz1HZU/oL1uNlf4pXhNC+58/NY0JDPHv6ELxnLEDIEV/m81bUQr
aKX846YbTVpp62RcbQlhVzH9o2R8sbthmht2wEKTPT5tF3r1fOcj4qOODb2b47a2
aKRgkTPQahtVVnGTRJp7H2fcc3PZuPQSB822zK8saa52xxl0lH2ImMMZ0LvefoNP
RSbPdLKw1t7XiXW1KWtcuavaWhQVcs60rce1LkcMDerooitUuHfLS9+ZsMgm9Uou
VqYGNyh2O5acXSzxOlUIV3ewTLJTAw6gOPx61q1mkRo55BrTv1lP5AoGSyFUT4k8
iQOLH0abRYTAkij1SBadEwiPrAxTAJJWGKA94OLUF6Hs+mN1eCFGyk2G5SewkJLU
bOsFNHEGGK+Xf4xv35Tow7r/miNyYCZPhY4xgjEvhE18T1Bljg7eIX6sS2Hpe+0F
Yv6F3+yl1Av8igbfy7nOWAzJuN1F+Io6qw/7Oy1X08sm2uFkDuKFOWkpawIPN2Ox
FL7ISj7FWjTBJVV9MNFE1+3/xeSzGxHLlnXhk2cZwcPTg3maMRj7D2ZOlB/502Vb
gfC8VHnJKGbeJiTjRVLV+t26wkYqMp1uXQZnCKdCMwdCJvKCEjRkk+27PoUTmhjb
BRUk1xVyvISqQlOU2kHJF1heoGLxQ9+3LtBaXsDNPnSPxMBd/TrvhColOoDe4aXm
yc39wUyC+aWpVYk+yZhyPgLhM5Qrf7WGCYdACeNinZNRZFiVRcyEiwUyCalkdact
hp3MyGQLLZhGRSKdgSGPN8D+xOSWdyDJ43xSj+lJAlEUwNlT5mv0QG2+FcvYZjB1
GzvDYeCnA7dEbyI8PQ8gH2l5Q+UEzi+BoqEC5qtd1iwlCh92yux7aRczL3BNgDLQ
SG0e2aR7tt4E+57pkbZo+pI81jslyuTkdt0SjBwOe6RMS2mru5u2bbAhKnbUlnfJ
Mudw+SYcuHWrlFXAe71LyFPqzu5zK392ri3VwYW67XHnKSAihNpmwFgzxfcCJMJS
ASQZz83atievNNvZlmndMlNt3Hjy5e33WpH8Yi1i3wxdjpupE3dFr/MoFU4MlLMR
ZKoXX01Cj8m4L5Kh1yBnAjbUOFk+yhb5gDPIo+lYgg23myrSiFCAo8ahZIGhueV0
F2eZ6LM7rkg+eGfxLYGZRf3K9OA2ZZiPiCDL7ZLmhjOp0DzWm5OzGLt+F0/J0r35
VC7KBUsyM+mLag3rUPtk7WZTyfQwkQM5W4pyIIW0U+48+3xrabfr/8dP0Idi7CnT
dFu9VtsSRuZyRk1p+l9WjwIMNyBg2tsIJGhFSN3BsBpbmW6dS0ueutLMdwDdrBpe
y1sx5zp1CJnFBNYhrx89X2dsY86zeu4B1O2SXGoTTwVZfFyuesZk04QYV5+nWzax
UHVR5kT6uulGGLbqHqk5pHgLAIviyncrLaHNK72eavJz1skAd2yoCTVDX5elymqH
z9h1KwUqhGFCehP0Q2WCaRLppNNfFkxzgOJ7TO7O9vW8qdxgTomyLED02SQRxvER
BbdoLhH08kQKYW6pb0a6vwvUw2wf5hUBnPTaXTK6piBBPZl+jvmZqRG09APnhw2I
xUrnNiBeM/srlNb1nvfRPC9xMXoNGbZP4MS+oZxwtHxOcAz50n2OSqvHU7h+UKD9
KxaPpTypG2Vy39HrsODug46+V10xLFC1J2uBkM0nWe8YE362JyRPMQGT7kC5ypnR
N3TurGdPYAHPc/Q9+UjZSBHF+GJFuQynsTwz9Jd0Q58DxdRIgvdrqLDSqPiVOuVS
yZ75IsapXF4B8PDjxuaeA9Xk/q9D1sI2CFQch2Xijs3idO2APSFBLnpTPSQAtflM
9cfyb/QRPYpdrXfz+hxkdBnfdOYIU9amYLo0/KLUaXdHQ9QeK+w+7EBL6lBKbtwt
Ooz7Y7Pge/QKrv+BuP5YHJOsuIF9TWaCO1FAzlRkY9c0Ovd4tGVBekJFXuxNXgpR
Ym646OiHVsNdxePLCMFCaI2toPzkonkbsLDfvrzO77kIDCNXtfZjL29E1wsysKpR
WKo3q7KrKtMtmCWheHFquVIN/2VyYfOcor1kNjrdn9UZ3CQzDn7Y9xnZtRUvdIuf
YPkgJilfCEB/18E5+ADAtpx3e95HtO5KKHF0gZUpT1wXx+6jXWxj8GA2UOy20sYL
PLFLZ6Pepa4XFTi7p792uGUNgM5aTAVmrYecankwCFm0dRd6YjvJ7+moWEsb8zZA
zweTVwYx8HRWpVUmG6/aPqyZ3L4Jeap0yJR4FNklckgo9NfmCj7rTld1k4r8Qb7V
OVaGWcN0gGEUv01kUiH2pXdEyVUxRQGGx5PMqdXDSNG6q5TMZrEgRmcqJWBywD4m
6RUzH6CFYWhi9MhZMb+NUyJyxFwOoc2QyrLaJU24Iy5113mSHaUIeiyjNTSrYgui
/fzeCSnZphVuGphuLH4GPD2R4Aqz8aIXesyvmqXsw9b277v3Zbb5CUpJErl4Clvy
pCkH3Ht95woph+H8hwOjLTmASOIa7OATsSPGwPrFBp1IYSr7nzT/UwkqId/Wm/Ct
AFaDKm3aDKKW449IDQ64B/X49fPquDpEktJeev6WzF5wLpUDjW8SGoEjJ0u91qmI
dq0bn6linUao3r3nDxYtSNMr9P1XdG3taM9NCLomoHEArKzdr0ahkls4XjlBerAn
pz+4mpFrwCfSZbTEaDrdsJIqlQBT7nPdYqFbyL4XALdSxRBrozIZusAdU0pnihcy
cctkdLhAfzGl6sWT3ZqfKkqeM+q3Y3R7GB9JKuPSU2bcCNRcVvECFseeFBRTqGsn
/4ROV5pYRQr3NSUxuKGuDbyd92gGizaPUbAgIrW62eGZbylrLq2HHK1GibZdp1gU
WsE99LeFAnJ0I86+zhVvhw8RhaomPzzxrUoJ9xwBAT1LonzZL5mlgqipeE/qPLoQ
SahSSpItOhUFzCVgMREzKHBDt+/6whGedRaXwl7Xg/LRX9821m19XGLIm9pyh9qO
YWtAvYyfIzF47OOR1TAkeT4bHvBVhS8Ihq+ZwYnVqjBfuz1JsfNScUggYPRV6P3W
j1k7yD2WILNUYQH107NmIpNA/h4fZ2Qp/ggs05SC0FaI3rdTUEg8oRvkxIsVDVUI
Oew3ZKng3E9T4BwhiXWIsbHUIMjKgSggagNOOqRl2qIbWZmrbuOFF0X3fTwQivVj
zK3j8qeDpuTjbgUGMkpNdz28SJKZ7aUICLNtLGLP4vZZpI97GO7ZM/eg7DmPgKDc
LfOem9iN2MfAml7mWqRhWeliSyAZN6VdfuCW32Vu/DEqfSynB1Yc8eJzetxpnUXn
PWbGh12IQFqbz2u6xegc3ixfbBv54Ov5kQ4YdFuewLOCGki6XO2OzJbK3pc1cHg7
RPcf0CDdQ7ONVAH0kYCpozzoAtRRjBzYlZ1BpejTgNbkjsrCphKFdPQOOEiAyoOG
nqijj2AocpJ/KGLCr2SzkWQ1QEevJNCWtwgHpw7s/oaPDtq5M84zxY6VMu+NH6qa
e4tkeCfOlN9xyIAdiPTG9ceIPjkiKuwYQMIm8/pN/jpveHn63xT7qeKvKl6mTj4K
e3O4aREzJWaeAgckeEqwVVFaVWQyGT82ZRjhwTpUmvZ4GQX7q+0LKY/Fjb8kSKN9
9gizLVUk4A8D8yqLVx58nfHvem4A0JDg4SyhY8IwKe9JxBHfNhMZHRKB0VI1lIIc
5pKISfxbA12MN7BOVBiwC/HgDly0GT6L0f9ud2XGmsneZmIBqvQDfpM/oJTmO601
5J+tyjUhbhyJc7gadzRBxDzud2Bg/gUTA911XfhkRXAQsErkxHsflBBtBW053J6X
vfDmo1pDCTWcl4360aVc5nb5fs3QJOOcmyQYvaWX0YtbpUS40i9pN/0UOqop/Yqd
JvWPMXMyPY0dxca3sZjjGP2kKkQIYgHfocqvp3UmcohFUlLlVp0l1vGwhSSeFPXs
Ww1/6V05/qdDg4XcO6OOiT+zwK59hIXFWKfWrlfrn/xFgwYdlErIgKOpazAyWbhU
r0IyMBsaTKht5RYxFziQgBD0nDq5fHQq+KUIzOj1wu2+kJ+brKV5TfqARu5A5m/Q
OkTf+j2oxwklFDNcGNJ9wCo9Be5tcQ48dOVr54rLpuUMp1/iC3cIA8PqG/rl7vdv
Xqq4HAPvRAciwqb1kVLwak8Q6PIG1cMwFcErfHgxEpghH37feqU9D3fIp6lynFKT
Gwess3vq6FKHyajRfhlEpXNCGL5iznKQ4sB31vbhe154upOoZHYbySM2dn37R+5e
1MWXNiHdOp6s4goO857MFkRQP7VQsm/k5ApRwtsv0iU8V8ktYpQv0Bgqqf6RJ51S
Djwa64MpXpu4h0MD/6IYQO0PxKAy6hJN1I3RdK3BuwYvxtg/+1v9Gzkj8LenF+IA
1+wC03e4PgABRvwObUZbbKXb2oO5kxhpbB9xpdmJmK6A8mewZAJll6JEjpkh8Nsd
PlGoWfD8UO42HgqE/l5wu9whE89WQHpM9vJaDrpeE5Zwk8kznyWE2ej9wbsnd71e
Xn1Gua2R1x5b+vI9+9Rbm4dtNDnNPqbNHwUsMDxD1dR0fhM0F9i83Zc/UtAl4MCf
k79FacUO7sbmoNSgqQxlwrNYb+rRrXhUQmZyTIQa1ls3V/OesBcw72SLBHXS6FlM
0Mi5cb8TpD3T7/BUr7YaLDtDWqP+ScMyc7t4ZJsYVEXXzye8dgDkYoKZaytAAo1S
5LMxehRcxJQbhec66YBmFoQ5j2vuGxeRwqra30jP4aVpNY2PtqRrbuRynyQlQJJ5
g40LFZ3aJ8j3qNBpOBuOPpMpmJ8+VlNA5GbAit1uCUPHBqttGEEaArokvpESnOeq
rLaR/FwYAP4s/yrfcOqw7qN1Py0JKmDuIqS4FYrZ+QcKI3vDZtOoQu9Sg5KUNfns
79jQuDCCIOeadlxcifCUQrmLG+B4KNFjw65aKGKQPb8MXVUCpDegGrxaB27+0vfh
qNzst61LT4se4R6aTRfDmq+cHLhbv3tugPIq5aSM4JJIFgO27In3yyJhBi4Khz9j
5h0WXGq9PbVT9hVHRXL8TnNYMfowFkUL2Ae+K8xP0cd4oqriO+FgVpHMcRW9PCAY
/uxrP2bKJjSjnhojlEO7jpEA3s7iwxaD2/avDB0HMHeRgN4dzqhVo3YOs/yuhCaZ
5WtxeIbq3U9/PPD5FywjYxiRLq3UFUaa/B5NlssYiiqKyK/To37lUizZUo8wIJu4
dlu4uYBpveXoixBK2UqE95NpRaitAwhTEUh5g5xDY6H4Q4Fx5En8fSbbyOwpV5/H
ohhgId/qOuVmxAKokMB1DbuhWrXUk1QPGjEb/ahgVbpbhvdkAV59ZG5KjnLVkm2b
fLPu9v69i2wCYANYnhufc9geAbSMacxYOTIM9U8CP6WIgJKbHbJGYRqeI0R6A/C0
VBt8KfwZl7LXoNe+BJ3eNvG4rsoaVlhEGuS4qUpvysgfnZk+4G9asWE7hzYWg5+1
5lIe5dpVVlfZHNpgPsJ2Xcwkau9tzdrGpwoRk1V/1hbOQhf4tdF2sAf3Ql83/zOx
jkmbhNazFBwUqLXpLkyVQg5kdnIkeVckspU7BZwVWYPSTklInbcxbmlDRE3O3mY4
tLtNg8Jll7UVSL3e3iErDinFCExDwcY+PcoeBQD8e1KhL3fp+X6YGAtJTtcma4+f
8mgAlv0Sl6q3COGRebpJKIoTJPnSN1MqZCWbzkYg99P7FhtqiBw02zPIcZx9Whtf
8wvRFHMbxCEY9B2zt4sqD3k59SutufzvF/xpO01kcBoUQwYTVnFD6wxrm3PNzky8
A1YhMIWSTSBX5ZWHFkNYkfl/WY2xzOqoeuktU/CV+VLulkvY183tFeyiligDwWNK
SfaFjEQ8hcvyKBuwCuk4kyx0EyITIHJdvfYeEeWm881Aju8iSZ2bgns64kYtNAXQ
qhAQhcbb27xeXJPsKkIphIVx7Co3DuvieSF/UiZccBnGOiiInNbpI9cFcTSYf+xD
kCVJIQsIzjoGrFMdL/go/onmVvbktb5oUY+Qyq8+jot5k+68Nkd3rP6tsj47hHyF
crI3yc8GUotjW9INPOwmDvLb4zgOIva9uPvnagDblyyrS8ccWz/pdFN+y91+2xTS
Q/NeyL5SdfSafkzPiBxDpv8XEyGZH88T9fKpzY9efGGCM3vZHP8ViSMeBP59EWvm
dwQAFOse+3x4WQWT4FlmYr43CnJypz4LY/x8z1C1KVZ0kkfT4jT0DJ/dNxRHx+yw
aK0jueg1BrxUPCXTNzmj26C4w4vNhCMVIH8L0Udhr2tv3S6ufCy5hFPeI0aERZ+x
j+zjpS/p4KiVv3mQKgcY0ZTgknJzWQe9i+pAE0eYX7KWd6Sb9io6lp4BqfEEMpGE
XR8J39vKNthvI89N1KB/U9QI9CxosH4Vs2sc7eJwejM3q9tGjIbU03kIm1d2PlxH
Ju3w80XROuU2JPqMovZThL6DOYJ9tg5TQuMwR+oVphb60v3VNLS2c/HfWDpa+67r
CkTqSsLnai+CVoGp3aCt0LLblaVUkGdjManlnyhpYejHnT7AuopQb7Ge/V6Wi1uL
z5OCMxnhImJyPcV/2qc4iqHkPbFBUUtSA3sTgpnHKDn7SCBfhHhQ7l61q6/4acOc
AUy4tLb3w86Izup3nK64o95bn9aKe/kZ4rh57UgZGEizzW1OLTcbCZGRNkC3+fAo
jC5c2YldtgMbGVYP4yCc/bBWCZzt4SiTeZ0h7zy0ZHNvDLg2N8VN0U3K9RCLfjdL
COmedHGeNG/cDniJK4CgLmYKnolBnYJCJCreOvCPs4fA7J+Rnaid8eNZehFYOZ6g
vPlagvc3wXyxyTojaYlOoBqrFaKNaEOWzNSta+y8gFkyToqj+1PkpqZBl+OLNG5z
gKc9YHX9vizBSSRkIkJ1J3NhyAsJEtf6wD9BEkoPJdPVcmiLioDLSny2jMFpvTM7
0FpQRZJFAJDaXAujz5W3+UqfM80iidtb8lcxWXnRPkeGoCiP2DghOmL/Xs0I1ui0
2o3+123kpejszdAcvBpqGDDQyex9RxKI1C2SydpBjx9Pgw1+2sCswrE5gDsm4f30
sxVqRPGqB28R9cvVFAQFgoRHhfIC0SY6Ytp98nHHAvb4QknuaWMlxZxZNiXN3Tfn
PVhtHwjFlM/GdWiiD2+/kPxqUDPOqPMShCOXiTcmSli+iXqMVnrk2rmKuMYjGr3J
lRIZ4dlWaQp6/Tpmfent512wDWvX4IGp1fPRrwK2ilcycDNMmIfbvb4EvgcrSXoH
Z5gQ9EHPPPCHrw/fs9f8YRnuqk4oP0N3k1dVg1gbO2wjEHsX5JTN1WMn/epP5UNS
zYpX6+erlMLQ14KDsITh/vAqTmro1Lw34jtLr/uPFElk6LbTNiYxUiVOsgmdSsTA
25qBnl7S4Y8qe86H4EbFxyKH9g1Whsw+rLksIea2hjqbf5vLcUC8idgT4irrWWrF
db0I22KusroD4aPV+L6XjEhmHYWCnNSY4ExgbWrvB8CinDWdxs489Tp/Hp739IBh
ha0J3ESJXMQQndP0CjDGHQGP+QpM13V7u/pQ4wnDT0vPzCoFxdwN78V97iLbZXMs
CBUI0DiEtIp4wHFB+6JWgDcw1l1w98DeKJ6PHPcm3YAMgDcCZR/mpbAnBBFvkjBC
4g6ynrKyRu7C7nWgGUJywq6nOUdUqxBZ5o+bCDMx6HmvWtd4VTU9eZVfQLR5SMOz
wl/7M5OizytOeDOY9ewT3wGTUYg/P332AMaLaYNGMdNxsj3guL1yUuRcpw2CdgL9
Me3ShUcSl3lvlFDlM0hJvMjc+YtLGBLs+zle76YmoYA7m6f4/bnnwbQ+a253cVUl
/VhOYjR8wlFkL3fNF/9jn6bMa0LHTY9DQ7tLByza/iOMRirCkibzpuKx/1RzjfAY
IKwjfJCrSe0XhAavUNt3G+Z71s2UXN+nQTYqtPUwESXwWm6wRcR4Z1cnVKfgtApv
AuLSNwtXmsOg0gq61PtBIWCMd8yFiOis+I8q+zMruDdoxmR5PmyJ0+tfNZba+dCb
MlWofnGus2efril2RyntJnA0j83jWv6j8kgkg8SglIuORFFqTCbOctOBXawT+ejn
WBT1+3m5SCLoohxUnOtWEGYbZhP8hZxLIIqkPQYuOo+Gmx739ZW3NZ4ORkjXraL4
XqyfXWnIH+i3dcOAEQgFZ1+SU9vkwdimuz2wOlSWSNlqEXRMDaghV/bDV/GXr+/i
vW9crNXQIPjR0qjYpgsmUV2FRvzAWJHNIzzG3wpB4g8q8Z3rCg1IULxX/oGSCqie
zdBRA8mC5hOYwwop6xxghiQdovfaszt54C6Nn+bVoC0Cb+uNyNbY76UdWOYJJd+h
db+INhWr2289ggyumbsY2FFcpqXdT/oPXNuPZhomp/DsqcU16aWuifhnH29ePOk6
FHn2sIlMN0sxRuRGr56ypQlQjlBBXFMiBhhYwxIBmcI/jir20XLw8m1CQyl4f1j1
okHIM4QFFdmF3wknylR/ZAiLrIErSx5Q33ekDMLCo/Hliz7+DPUNPCD7p7PlZW1J
wdck914XuH/sixiFzwKPCaWL+gNALtfwz+bxH/Z2l2ULICzRjvgneIgFzVZdC2vn
IuumIn539LxqNe6RyHdu1wjbqG8m/d0k945TWHo8Gli115+hBx8Lqk/IBt/blp/U
0qdyj6d0VidsDfWG6ImrpqzKHycRJw+SapRfErstWkJXYPxk9cmfIHE69z1x4n7I
Cb7TGtmpgS5rGI7aUZq4meVHQesTegrL3Tez/RXq1sjZjFRl9/akpnxX5okfDv2C
xjbhgw9b1mi5H+bYLvbNfNDDG5xgtJ3p/s9YKtU0qyCLo6NxorMjST62cbU5VOBB
RV8yL1Z4NZotRwFmJZXRQva0wSljaQrhThGrvhAeq/zFPUaMW4r3ohtkdO2LKZH8
lZ0ipu9FoEb0FRbPPbYrUqTcoiXzItLNDJphEbuVR8dSbXy3uCblS2iG+vUt+3r9
HhfltA//7mh9c1tAn2MHqQxgNun2PbvDog7SbURvP2zHknD0B8QEUkE8uoR0MYqA
li2ZnXso0kAFaWr65tD7VLYqCob9A+EWB9FNBTvfGsauwfBtBcMSqMCBuYMtvOUK
qHBvAZkUssNlh7/l8zvn3RgiLoBUGK63MOF4PDWW4mVem2uOHT1s1pkw5hnB3Ha/
ZTuzmFjyUIq79O+CcCNcgrzwDFdROUgvl2EpEhWfVa/9wMaviCYvsLMLgKTbmE4z
2s9irjTu8TQ5aHSYQZhjg/QNQWpAYdAZ/GpL2EilR8mlwrEd9NgJ3CQhYq2eMBcZ
HrnKkpC+3gCZ/3yRnAJ4/kcocV+OY2e/XzY4ICvwpWZHI419+nZrNbWaF20CK1JW
IDTYwziRYoi+CykDne5LTsqfAZM2SKgYkSYQiq+oHN6U+Sf7JgGtJQ+OE5R4L8n4
1evauTn5ZXWqkglg8TJqWlA9X6sc33pS+l2RXbT1HRyVrskyjkXS2+PhCIlsdPqV
SdZs37YIzwpQSvorLUBM7sjg8mgN+Bz6p1SPppcOnPSsBzwdmhRY6CpB8Q2DRTUx
y/w2X3qoyqeISyImhR6T+keBFoqthCJDYoxVeAM4BN3XhI/loEuWMgQVJXMbmD8R
l27c6t0g6SVRAObw5WvCQ2mHkxMUnwFwE2I/xYs4M2KItsz6ONXpWC/LM4X68Dyf
HrsJ5BJ7+fAHRdI2qLnAF8MYiMIYk23YfxSGqRm7ZnelpiACgNn+7WfWA8ME1dcr
Nsdbls59w+kztCPCxJQ6vllI5psQS/Osx0ae+q7dEmYOKDP5YskdoLeuJCsOljuT
GxqudzAGcsEt2xLm7nELVK9pMERgo6QIsLEZCRAW/VSuqihVV/O6brS0wD+S02q7
ruLjq0LUqVXTKeiGvw6aBBjYOhyC/a73nW61VJzjzyX6KuXX/DzIoc/3yYf1vb+F
IEg5UezTqCywfMz49d0V91Saj27anSsqq6bG6bs7cDlhHAaXg0RuCPe7YT2qBF04
Ugtk7c0wvcy6tdktW6BULgw2Huzdl5Euq4JbTRvbsNkhPNjs0y0mgG6Bx/13Cfrs
iphyVPsW+aH7Bl0Xa8drBfyI5Vai45uFKZVTN8MaaiTBCvZ6VGhi34P6OXWr49OT
UctqivdYKSeEbE5xtfkac0NApTBfWSLke+3psqdZLO28jTdiNzgW3FEbPxjINbIM
xBTuvUOKUyyah6uLzyW4IjDx7v0ZhpL2pQ+Pp3+Xp8sgKexS7AgkaCwJQYPIjeAj
TrtqXGyfEfD8M817bdV9UIR3RlGNhwFMMBzmcdSD5efKiID8OAdQ2CvnhA9+a58+
2ZP5fEyziHTDo4qqpCR7BWbwfwapXKVJNpIkNc/4xFl7GlVD1MK/cWafaV4jZohM
Vob9XUxvKzipPC5cmgmjlTmGcIgANBN7jqVRbo+aGa6EW5JhKUwxu9TGOwWTbCRK
G4XGWxcocRexoiY6kLTN7T1lWrW5lReK1lHzuKcIyjvzimGdOkjqjdsB7NnuJRdK
ojEvZRqY0HInn8oven0H2RUty9s9KHvR/tMNiV+ht/bM4s/OLaBujFVrx6+WaFM9
+gJTidP/zYIvYmxB9kY1IG12jReB/ry7l4r+L7knVjQZ1qjN1iKTKmLalHI+rzg5
B0zARjZ57jc+XxNt+hcZKEolnsu+RuGLwmwXMRMUIEXKhnTmh1mukAfK8P7AHjFn
guOLu0ewGY0b9+n2glV0lGaN3FrLxq8/R7trC5zr9GbivJAKJewx8b8c2kwc0lRH
47XhW7WyJtmndDbDFzxnldqgp15hwyqTlKRn+TLwepBV1+X4/UXHQ6WkHiuUXhOI
Sp5Atdn/IOP/1io4lY32LMuiaWmsq1mHGyCeG6E9PnqsZ0+zzz+JONd3KvLM2ZWS
QUhSBg/5pMzxmxEuKx1t6yQ6ppnWC+XmKuQTT+3mUhl1mBSgESSEHrwMsV60vSVx
cWVxc7c4xqpi2cq/x3rbjJQduwDx4NLdqhCWjMqo4g2kKmoETauEsOSo25+QJ46E
KMyjpnO5yTnQdbcJlPo860Kn754QeeFimPyP4RFrtITjAw+Php8CZ4O3X7joPcoq
CQk+todlb3N5UFeWpDpvMMLp6i9YS4dJMbaMOUXqHWeXOTv7sJ3NjO57UgBM//dL
oJSQLyMmw89i+P8XayTw5xHENJchixvOR++WiUzRy3ZkesOAxW/Xlks/MZ7BIBiv
ToM3x3rNY5qIeTn7kBLNhmMcxx/5muLhb3GFH2tfQCVBukuM3icVz8e4AV7UPopS
i6r41ypVcmixmQ7wNIocn8HS1VEciAA8Jllr7AQ0uBq75THg2pNAJZLUv9q4W7Rb
DeqIJTtAxG0v6i0QiHI7DLC2CtO0w7gw23q/5sE4SgOENEwx0bkjo/UzaTeYem4Y
DkxCBTzDAFYhcZiz7bhM3x6LAA5xl8D0OkSOhyB6FuyK+26PYIofEtK2PnbfySIs
T0ZHHfK9X6J1Pwv0yN3wpIix1/K/werjidFfADyKTmZFs334n8FTCWYglZw5MXTi
C7teiZeQjPHB7PYDi42SfWN7jyd2hqGaugCOHrcaq4Bw1Gu0pqHnlpUYAIrJD31m
A1tGuMMqpAzaxWLmEV6g+oQumfgB5UZxIP8JDh4MaTUkm5wULU0zZqF/Ra7a+gON
36idUsVTbdgkdTpCzLvb2oKyE7g4TGW8sLKT8jmbgN+EnFcxNf+BAPqOiQY0J95B
Cs0OG7PY6ANUdrTwqfRCuXbUqH8CQVnkVBAxQg+4blVYYjmUyeZw5j1/nlvELkX8
zI4WYkwntzkXlc7YXBsrpaYX0BnCLWdEfTAmIY3p8mHM/7MZYaOUL9B9twIc5p9m
WpKk4aO1y2ZrawXM3vzWV40T7HW5Hk04EX15JbfQFOBVQ6n9vgoQnCvmK3nw3Kss
4R5+HIHvjQCg3SaEkIjytMzqcN7t5xrEiz+D3rQLxS+SmLEKaq9cgNhI3zud5iSL
155pIxsqfae5qMKldoiWwwH1VYKRtwjPcGY/JnEOW6VDC5W2hwUgthu85OYQgpFY
FCdMbfFMvubp4pKz4YYxm+GMZzk7IOn11Br3eDofPDR5ZNW2JnDud6Qfq43j8IeB
m66dtn1smYsewVXWpm7uzD1/dc4GgGkJCPpY8g7q0Zi/KMHX0hG0Ggr7TszEcT3V
U6LiGGGkbzkEtimEyt2zMvUAh4KrVRHci3ile+xfnQI0G556yH1A9970JBWD/bb6
nYqaUIGvKZ8+MaEJ59yA9ae53VCDAsqWrx3GV3wxk9fvcSAqEQPS7EKwKDSgFcaT
YMP+eZHht74upMadzVROJfGMcq0ZzY/O/EsDPzCtfBNpCclJw3zG/tFq7UR98h+a
jY9jXusQ5Qgz60dY5Pbztpufhgs1sEOAiS2/4SY1bV2nHvvqGTyAOtAD0l4pSdyj
mJtbpFeTL0AxmO4XQ5Q4Kud7X9Ys+oRTSCZwtn8fs7JMqCA7U5PhpPwVc03xCYL9
SB05I4Ig3rmbWxrGvznvoVq70jtgBqb3ZfIwg/xNwNRhIUbAFtq05wRfdaKk90Kp
bM/mRgGVv+ke+x4Z28ozferyIRwddSMsOvVTZg4PV84SbQ6Sz0S5ijaT0g55nRGb
KQSs7xDi00v4Z4/3k2eVeDxorowE+ySFj1rbpSajD8kpyeMbIMwtQTpUQx1b1J4R
HHAGsEAoNgTu4IbIOM9J9PUJrRbDYuVncTJbVGmpxAOpHbVG2teAyLxnEdS8gB9y
HEx68J7Y2ObVBvpe+WwzQYrePv8zmbKjG9w8xSJ15GeTeQB4IyE5jWkNYDe6IRQO
hjpQw5Efz7X/mQOE+anuxKQ46LQp1soB9mPeMqEZZytANKM9CMjVT6ATs1s0m4gF
WEamCXZZBmPW5JYVnpRCLBJhxvngyTpQfexXsaxCQGQmJZreJ0nZb4GzLUE/hcn9
6YRmF3L5Ym4GSkDKF7Zy5BK1pRdbmxMcvN0apcV+2+Fd2WmteDlGGnhsfjgJzYCA
DwJk063/3At5VIxmI1q2tpZ5Bcc3tmJJS6rS2ja+jpE8sF1Yd1Cpqyx5dkDqZoLb
Mz5cfuebZp2fmM71LXgi5QccmxF8RF15PwNUGl7yWG0gMiGWcIfrKE9wedEaipy+
wD5s4VkXCMbwMyC6Cqb71njeVzThi/rZPnSFlFBEZaFeynKVZjBImCWKzNHuPatV
Dvwgi3SW1k/CsfZO4JlfFR2hjaqw6odZBSIhGv1i3p+bBCbFu0Goa9wpVCmzybEs
tw5WRIJX2pfE9kge8syOXoJTZ1da+T1gIvzDI5PahUpFFSTA4wvLLK+iLh5Bf41I
dcMInd6Y9s34ZFDKUdTfjhmlIuwsDH8Nv4RiR+lwJRlkkLI2CLE7XCz3A4Oup4dJ
eePiWR/7Azzr1y7mmVzDORRssibfUeorylRW4lq/YopX2B4mTN4w2J+TLjsuVsBd
o2b5NvIpSJG1Zq3m0RzDQIs+kTLoKK9wAAIcmNxiPE5meG58Rp87B5FwoV1k+mcY
sNWO5hdjpvP9V56t6nRQbaKTJOH/HZvQGYb47kPGHgkLewKj7aGNbZzlfxfEBZ1i
Q+b2v4qrigZA3dT+GbLSwiEDnAb4+KHka/ANAimKrdiu8vw2UC9Q6tZsJ68aNwo8
INWQx8o38jZ61x2bfOaeWYtQeJuLOfNAUeuMPB6R+tRaMl2WM6UAtARs/lmkJ4/W
Uyhxo3EY2uflMF5XvIoyxDSwmTtJpV6IFU8o2WYzOM844KmUbTRK3Q8YUlhsPLcQ
8mEKF0MhIF3kOHtGwMqh6lcQfx8kBqynEqiVk+D2aGEwsACsbIthSIv7TOj339DE
TuHZ9DpNaSUKlpw0OTA1EZ44Z5odpCEn5i7PDHw6ntXdPZDNKwGdTyQI7XVF4iUI
aWrLuhGehmIwh27XRMlhmhISb+GMsS+JXpxYp3ypK6Ai4NQbzTh7HoqXzCIUb6bD
sraLbcdbXlt6+Q9h6kjdBarl5h+X/cevnHbl1a1lrpjVk11oVHPrXhu0F3JL2WCB
sNvQhpelPntiNj3tUq0vqnTKf6r+iXueXpL949rqK8VmFeA5ieUW6SVtmQc4p3zU
idnCG7XmyR66vXVVD1X7pt0BWNgX48aA4aCwQRVZ6TnhRBIKDVAemg4w71elePVr
CYtf4sZSocw6DdpADKGdlVZ9GoJzAikPFh84SGLZ6RakYkdvcWPtp8l9lHuwITnQ
wOhLB6H1V/saFVgXbVfiZBDWzKsYNpzTya7QJWpdtI5GwvhC6mpK6mxKkEy5uM2w
aAwcAHfR3CHc8r/4pTFrs+C2ZUMeBM2kJSZfuilFpjUg+eOmOeFT20nRvEihXydm
jj2csbmpTxmoAoZx8CE3aFMoe6+YZ7IaNXM6XqgX37flV+P+SI07RePwWDKTlvW2
dUYK2v57MWPyuzb+jzLD7yp8Zb7vQV25uSsgi6L5A/saD5GAVhjv5Jv3LAuZvAru
UHJbyM5jRS+41v3CqZk4UMeNch/7Ew1f0iHmy/q0PdIeM2r1H5tPAHg3pitD0iBn
fAZMhAFR9ZMJmQ80evrWKWVMoNRRX23mgSGTGJdIT3NJ7ens5rGF4UMzdOv7exuK
vyum6sLFwJx/2Zc/UXNmw3VSUFDOR4+9AG9Hc3eIbIAE+NqflRQIJoqF8MvpqUyV
njAxAyTXiDVSSNO5zjnvJ6pbT0siFiF4Onc1BGf7OvzuFeW/DTnERHhel3b3yY+7
Ik/XLkUVl/r5C0oFy7XKnGze4gBUsmbLQgSINRCsZHuqFb/FUsRkN6v54w6JZZyG
5FrUlZXj5EFOn9XAj4Ct5Hf2AMhll6GohEOIsHrJu73LK50SWwMfAAmIOyN+F5lB
bnGXgiSmwly0tHpbeVhFgZX3daarmiDSfEedvZ6xmn59NsGVSqnq4JMVq9eHNwZD
jH28SzyMY4m6UmIRLlkKscn9VLdYnX6hPrFoIJ77xRWuay+2Wl/JytDBGaYG8LFT
GlJksXbLvpVfPQw0NbHlGnPzkoyOeFxqCb5cM9kP5EpnSgwBPqcnTpr425u5eXrO
ppZTbWrHIEaZ3x6ulbJHLT179gdmohf5YLGkFpu09DPITVsaGrwNI61QXkpT1JbA
Vug73elOqS669E9q7n+09DQOdoMeSxGW2Zrk0U6T3Ie26kcIjJb969S1qURhraGl
QHHeSvS+Cwl97JNoNAM6wLMlp7xlya4deCGsTucAAUOEhVFPkIf2N98OhW4ahDel
73ArvdXTYsw8i5lJH4ZR7emM0kQFLoqjs7to3cay7qxZAmaE8umvKofKwatoB1Yr
B3lOBcwIyeM3+aAZkZLJRLbZQDkYEjfZ7K8BywUan7mT+3DNeFajT0JxLXoXZeLq
Cd3fwL1mzVlckaaAdQ8Dc9Dw7MsZI3XfQz2eu/HZIS0yGAkacaMgz9zxc1dDG2O1
eUO0j1inS3cacnG9B0z7iSkaMPhkYGIa1uIwgALGYDHhIxIGrQdW5AzvPO42S1qm
ohZkkmiUgc+1tWIlwXHfSIA2/3ZLprMC88SX6BptNdSt4lOkZf+MDJ4QQfjJkanc
wuTaXsVRqW84Imj2NewZvKGy6gFd5I+azLa3QlG44SYsurecUlXXtN6ul3fAyBLx
7wMDhV8qdb/NYT+oQivDNLJRcwk/wdQzuTv7xFRemv19dI8JbX4Dk+CtaSJAgEdR
Dhbg3zu1YOdyYWUiU/meRKDd4EIcQFNu/n4LSbTrPcCDujqI+ifmVk7grkk3pBGf
R+EbrwAqxMiduUK8dWT1p+OHieuc91VbV6RGB6pC9D4tpLiI4xoEcukwfhGpnHky
v5p6BbGimfeU05DLCG5jirRberyEB5SMip7kBRHGu0KPt92c87QpWgEF/hKJGhk9
64CN7P3VxCA2/74PA0EbgyOKEIyubCb/OL+fs4jKjsvuFc3nXD1A6qZ7HRidDq/8
mBD1Gn7bk3fZfvdkt+6UWvN60QNEkxj6yOT/Fh0kIJ03vrRslN4lK+TMrAn/Mp8k
gYFpL8kY2WA1kOLGxOrTKaPP9UWC4Lw7q26LNY0ZJB+ow4HILj+xyJtp5Zskjqzx
aXnB0Q8wmw4SkN3qFg5UMits6LXoKg1fsFzn7jmgHhH6gOwDHYORiaDIlgzxbZj/
6ayOPmznbmkE9I/pQCVI3nQz8RRQNFjgavMBVS7LK+FDu2vmJMlkvHRyxtZQx2Gq
wDe9xmSmxLviQjUbOEfhl8gpi5ZlSvb9/UvFwiFF3YNvheMaVx+PHFjeEF0Crh0p
RkxJrPesPQs65Vmxzs58yitNcx2JPx3zfRIJ17tWLLflOtdNRYNW+Q7uZfhVlmlq
lidi1lk6fud1cCnVf7eFFUicfFScuf0CES6vKRAUsCC+bi0fV3k2IJF92HtoaAXT
PQsejni32lTrsWPqb9C2m183d8+GrveAJSLi0Zn8QmW0GyYoB74nwdhPgvaO7+c0
PhISwKN5rKEdKjo03+aUuhe8g/TzSYgM0gCgz3CHC9G7KJEmqq4h7XzWNCJuyNu3
vOkjQJPnQ2+WSVgYiYpoLGLKcmnveOtm0bsimLMzzzOtwJJ68NqFiYjvhMHZWPbc
MJn4sL9POCfooVRB4Ev2shYKxmo838ZE9+3lla0rZTwIpBE7rCAfDh43hnwfvlyb
SeCSQcrcdzxcMbb4d7b01Ahxn+KS9xE8fT82hkt65bevaVLcsqDWLHorJr9eu7Qo
8YbK0jUis7rRiegCmdWHM84+hcAGmqETltrvuqcoYubUPnPno7nDonf+7XKVxjN5
jhbLqrIdS4LVL+9jql0JjXtjYm3IBUmkn4kGo4o7a3+BxgB1MqFMjqZTY/bJB2ea
A6hmyvHWYHrgW38aiAXyDIcUZBY2C/acELDe5zfr4ZqEydutuFQo6krWoz/U1Z2Y
HvnqG+iF/Se0ttz+td4xmbPCUu5/4KQntGZhfQO+JnREDGdgXFGMKYMSY5FluCkT
GDEnmOjhYgfZLSApHaTqBIfrQ6xJQYn6azgoSZoLs5g1g+oQGBxL2Q1+S+j+Hzn+
wUsgEnxfEHUSJrqFiNxwrRzUOuwyYJN6abN2ceHPzt8YssY7t9jI3ckCHWQp+P96
gFHOsstMdXyr+/WI/zsDrE4tgUseLVtpzhuxioH8dqSiMBaUWz2ieW5PeMxj3dPw
UWd7tvfGZRJvSk0eEY7kcEHzMV2rEcl0FfSjvK0LB6KbqbYeT9Qp6Or1j/O4LjkI
9xwpdGGXqQ3c7Pp4jRIEOGNA4Ezj/os/Ke+Pyj+KxThd9qQo0dBkD+jncRhKb5y9
mjzNYPB0ktbdCCwCRAmALPwrWKI/tPvkxUp7hubissmiAgIkTM2TQTBInVPzCAkz
Aul1gxP9kRoNcASZqft9xkaOV8Rn5VfbGfPE6sJ2NPZdXuJZaGRcvWVAQnGOOG2k
ygKfB3oEO10Uy4DTyrLNL0GeL6odTaD/FaTY4IdfFp5GvLGnKQ4yqnyCjWvOsfk5
QdZWKS3bHoYCs6C6ixZy3sEzhKljNvPb+qtgJo9p7PrRu3VzfskgwcV+bgBZ3Z3I
A7K0l6hWrGurBFYulmp3J02+/78gW4F7RUNGowmjntYEduVhU71DkLJmJbB6Zvrf
op4M/PEvVQQbtF2QbcVH/hy7a1p8nUk5zijC05RmAAaCXNGKedyR4Z2SaLyAs/Wt
kITvdmLupvPZtqQjdBcp4dl8aIS2SOvgWjUapcAGcijR2wJV6kShx+DpS1ftS5Xv
sOzINEFBrj9u8vkGgdrDQNfUdTqS/ECZahvWSmU9hRDi0qUn3LAkhLCMLC7BexOZ
TG8zlLqfdRYY3RRUkDJu8AObcPh7+Qe0iNEgnTvArcW3SX0uUwoxgBSvx3tXQiYP
2RCWklChZ1kzYwa4HDkPjcRAwwhPEylo12gTsVCj3QSIoYgFqZeFwNOZ0SzzYT5W
EJYVF2saa2EBQZ+VBtSYcEBjq4YNvHCkyiWuaAeiJ9YiFW0LMlC3Z8vDkJs5Xi6p
7doIhtl8wgEX4tQlbuaUdUnayuS+dSfmCb7OY+Wd05R5uupD2cOgVyqAlyd2qXAc
BqV/T1ww4LuGhMp91ujhK4g4Dq7Oh5URm4OG87PZxG0S/L02hSRVlc/qrtiV0w7O
VSsqaq5kpqWAbU1/gsMOqB7VwquKQf3QJm5u0kcy/u6Txrm5FE8c8rKqgz5Xv4hy
wzFWKq5ezu7y1LZiKMyikdmq+pwCoAbrNb93R4oJt0dTn7/8zpVfdtIdTocWtxXl
KmcT8wCb9T+YXxfFVCDP+DgQzrETmAEsDeCRbQpPpeWD0PwcVm0zVLZsaGRGh/p8
EY2afROTwZs01q0Yn03feopPtj8j9fUta44QYECKNrq3L5ssI47IHeozmaWAZ1jX
I6jxovVoGtfoyVwnjvNJ4noPMF4dEtoVHXLWm9RbvCUbOGXbagD4EvMlA3DMPa7p
rFXB9W5dpFhTpbNPqVfUCmJ8zFM0NDjapllER/rWsL0qvWpsBSh3BVspK+/RiEgo
sANZ41t3hg01I0S1qi1eyFoVnO6UUGKylrCgg0o4NIAIvE2biFKbXsBEKY5i9tSC
9XZtWHe/mX0dWh2ReQO8PPefXTdemnaDhtXLFxAhmQGXmMXuyAdpJTod5n0Smeqt
6awTsCVXXGNF9i3wA1S2sgDBwtSIMfn03XcPx6zjWc2Z6yiBNQauh6aj/CavfoLF
5xPxV4bd+qY9pVjItV/ltdBdml9gNMcT5hHvBMyc3JSRPICfEgeZNcXTDO8bZARq
xCqNQMgZ88JkVzqLta2Go5MO6g8t94oZzM+fGqJXHhODKTv4M9u9gjXuRnnT1KxC
O6903CeCyC6pOBBMn0jVbZDa5sQ9+x6Tub/qg2fwLV/NT/hFb1yg8oZlOhkwrcJi
YY8xrzoROXlFwFb50o7iO/nRGJebCp5B/wf3JCkekqUUeOtMZWOGzDTvL+dTqhuq
s8iSEjD+W6e5XfGvNemTGMyqzDMbQd6+r+TMie/Jx8VMtE1BCVi1siNxAh4Wmx+h
73nLhT0bB3teNOtDXRsojyY/Y4P2LvtpVARMVRAUOaS4Y4Q4B9Pedz6FbSTi8WWA
E9iqKAgzsDaY4r8sdInfrPSk+aNeyPveoiT7mFX1a7UapyqByNl83ZMaPli/JxHR
t1e+D+Kj2klqoD+45UKM7S+5ArhLZPy/kJuHqx5JgzPATeA1i9bujDPfjRgc2aEd
GSUAV3nvAmnEV665p0nwJRWiqQ3BM796GznyN/x/oqgSIa8XTpdCY1+IivYOGYK8
BHpT4sIt3FySXO1HpV17aQEgWTKAmPMDDluN5fM9LPnaUDgWGqiomOXuuMPS3o70
/pfa6HTrn44W2Qh0PD0mnXOueSNA1xVSBYoMMMYwSF3R0jQ5ZN4cgS1EFEZ0vTxJ
C50+03tb2NOqX9CAe3gc5n6KyJG2IbhtbfmWiSWiDiCrujri2Tu7eOoA+gg3hpC3
2EkJPvoGX7pEcdwNwNjiljW96HGaIzaO2T1lgsOtMeW3x+WbzeGabnl8/4BiQPYf
1dQZTGQhs4yl8L3RcQo6U3mZ89Izg8TNE+t5J58wAZtnAYH7uxzmUJ37bjRFWg12
KRQ87KjhrxPSr/oeBcMTNb6uRIwUvc3vXt2ciO6DrJ9nOVdpXeP0m0YSlNQrBCTS
xyqupWo/Op0jiSkP0w0SWicbA+8M5kboOmnetFSw6dTrXkpMrqm3BJqhWnYwJZKI
oGpviptErpR1duQlwhEU3nU2CBBBXwzdXFdY4qaiqE2I2v43L1P9ygJMkRK8KiLV
MweCWJK9DIXkaGs4oGbelnX89HiNgL1PdzCHtx+GEAfVviGov5w1PuxeBqaJ5i1t
znAStKZ49sjt9bw6kk4PUhTjm5jZfI48OWuYnwlOLKR5IS/PlX/S6bKorm7uZYc5
izklmePyrv4Rtjq2CSa1hPoir2LAbeb8S+4J+2/Qq2tY2b3G87XSv9HFwvHt/zM9
K3Vi752VHLjIgRe4IzJRmzNLxFfJp62vVQm7w2GIfS+s/S5vIdVcIqqnpshhVYHJ
bbQZDTbKkPCY9Q09fTSj4dhjJMs2wpfC/jrIAZepmLERKUIud8qmbA8dJi+v30+P
7nRJ1OeZO5klHzrCbZdhp2GJ+AHj4PJwkv8NXmlk101K0a2t2tt0PItR63nBGg7z
C7RHtVLUNAy0HTAiez09Hn65cW0wbwF0k0KPlOmOQWtpr/LPX72vkFkmP2pxW7BG
nChQqwVWE2QNtUom8NDxi2vaZgNtOs5P+Z4UwjzeN8b4UgaGvXipm12iJO4w5E3r
m83gFWuOuR3XYFfYr7mtULNIq3qKKmFoaa9wDZwGsGxDnu1SQsnzkTC1goO3/jb0
ND4ZSciI9JUKRt98SRL+0wekiEBC+MSb/ZpeNLmt8XJMWBAkyfcuOQHBFacGJAcW
TXmhvXfLARE5MqmglAw9zRp0yoiJ0oYk9QbuFyGOxX1T4UVgURZ58IcfrsLK9OwK
WQgImGS+KqTPM9oO1ZJPX4F3DPPD4jCILmZMzP7SL6Z+QdSQJp75Njc+i7HY1Me+
HuKGb97XnwEI3Md/8GUHL/p+q06EBwOaa56pGRisjZmRGih//5LarrHduyHOYwEo
JSBuRFB6tg/qSwipp1XQXljRk2s+kEDrpQ/QUVPRarEkH0FhVipwSddokbGL9tE4
GN1w4r9wGR7h8o/P1Sa0ZarzRbnoaWEFk7Cf9ekrZfL3cHtgmDIQNG5cJgSApZvq
BcNVA5/2R0DpfybISIjZ8DtVAXkFNJkrWwlqbb3h6BVB4BEPKAMad+KPHtsuY1pX
y3wr/13ZtCXsGPmshxQviRjmZvNgKB3bIHMCeZf1prOSMNUWu37PYJpiMRvWWua/
3xqVwtiPIi2yHZbZeCpeV4y6VIL/p4/h4F8/owDEblsQrHhhVPcfWZJ6qVCCp5ON
4xl7nIOIoVOY5ry4xQWB9HuqD8Q1RnQmlrgwAAg/p6O11WeTWVLgfcELW+ZuQwvg
5GX6CUtABNsOqYRKFOjaVYn/Cw1XvcrBDylZ0ayd82aBx8k1YD16Mq5L0eTuJYFn
O+VhUMFw8UPmpldXozVnPOwQhc+FOe9/cwQo6igkfpSzymu29vo5+x005a3cOnyX
3ijRH+SmhP7aa4qORtjh0LJcoWXsV8AzyB6tWoDBp1axMvYZ2DUhj48uJkBMd9Wb
yaj7RRwjLs+35ZfqDobRHiFhYSVA7Z2YP1UNXtUotudLiFky8+3Z5VPPT5oF+AnH
fwNMSdvvaGRj7GuVLWFk+7nipNjGjjee2DuwnEZNMIGDm1pW6D5fdlm0+zrkJ7nj
TWeQqlFxWE7sBYj27PZcVvqj5J1QVwFXnB0R6En1TvPOIL95yQMsyhMf6tpkJEmw
N3XmEZbWO0rs+40WzUk1PVMQlp5bxsbJWpoTZ83lnPsqOkBaUSMK/YD4vqQRYp3X
8T7V11KcvbB5pyZ0CV06Q1KwgOj5+/eYZPcMtR2P0Dlu1TOZ5Nb7viNiRIK7EH5q
Sb8QEeVIlTD4Hl3FE8P+QC+/eGtSflbC91SlK2NNYoF2ea03H6znURxEZ1Pv/e3M
9anhbcCVv3zQU3F91Vi73B9dUuADw5fH4kqMJtS/kkbATpRFbXDbaoIMHzxl4K6L
Ae4jBYPfHsWfyY95q0SMHRdert/rzlpb76/hs+J/OsyfxKsJFBW+6XIiZiAGlDNz
J/ZbSZDHs+6Ld7kOiA/QZT6XNjl3f780SO6+31koDA3dsNYjOdpV7b1f8RXAXTFf
OP4FZkoPz7FFnQHmNvE+f2b9HqOApo0cAgS0yqoun/BxYBLbf4C1htVQtnPPR1LV
8lIQN8yStHjlBTBzBgHV3KxY/f8waHHJvPtftRs7LsIkHWUOxsGZdlh9b9LjR6ov
LVCyKRLRw1h3CDTLXEZ5R4Ap0+CPt+jfOYB3VDXSA1OtGPquIxZKFy9ibI0IjvkR
ysvP4a0jFhyl1bXy0H64mJzHQl5L1O6EHwhpBJRUovMItaCW0HnjI9A+oDUAn+O8
sRLFXbQyettQ90D7stxsp3OkvTZS4SBhnWtG3dEq9/Ocfju8QJVzAQieDSHHyCwJ
xaXKbfb5kwjn2Q0kuILptHriut97DdpIy39vjK3IcANYnellR/NU6gXI80sUKYPq
svyc4KL5iG5BJxVhEy1YAxHx7J/XLsJOF6aK7q/xU6K13B9E0ddQw+YK1F6oZlzh
VT48xznLfz+R80buIhLzSZk+FStHRumMcmrtVuPSNyN0zF1fRmJusedkr2GRR84M
i94/zpjo7Uao7YiHLcKq2DMj11rCGWqLRBXQPGS182+0SUJkGaEytU185BSdfWGk
uYdgKOQi2rWieYOxUCsTWOxFkI+VQsrNeHoJPakUTxHj8SdiMqdlDY0nhLqV9yL0
Yt5HhxF0EL+03Uyx4NiIfVCmIsgeWQxbbfcVA3lGQbJJw/yW7Jh6309cGofolPDI
nUq8829iS0RrQ6nrBF4mkfFgAJDf3orvG6qqaugJ2qwJbyguNLOK6RxbiiHNy+ep
rys2dh+AC73gE/oj7bgC7VYHzYiU1heuMB/V6uycgtw9x6UCfdGIM1Ay/nz9xxN+
pNso6D+7xhyhlccOSlRscLi53AmeOP30Wri70PL7KXG4+HrJN5+qEgANSKSsJMX8
StKMpqv4L27rI5REfC3qBF73UDQxyP3mXJ3kpUS9iHQgDAQ2P7X5V65efkuW7tR3
aTa2O+xcDkYWhqs2YoyOg9gHpiMUjbqQEiybzKeIUDJ5c+ynZsr3/xv3hvlD4vVS
eqKR3nNs8THYhbFw2l6aQLmGi24L6YVpaM7QWX57U0MkxVhq+XS9wQ2bTQ5r5NWJ
2Mo2Aj58wdxbjANoRndxuQxVnls7485o6MYMbNVmWGGYv+1/TF0O70kdA7M1rCIG
GmrBjRuqK1G5tIPlgftcBZia78mGbfanYiF4JWwfLsN0x7kiADc+kjobMiVGfV7M
Ag0CXdOMifGcFxA6OE5ID6dIL7RCKDR8ruvKqAFe+VO7i83vbsUEpqX5pe7f4i4I
jsUi7uEUEIqPzc0FE7VXRbCLNQcy2Qzp5YzV8ed0EiVyeAkIZPmVOMTcoVTSh8+c
tU8Xw/0GI6KdSbf739AeOrK7VHGxL/GU1FCzWnPpfwLqBrbs8r9ylqlRA7fod4d8
Ll3SHF8FIFeHi3B5UF34tbz/glh5/2oKOlcwbJy+6iJBCrelF1MA6f1rto9v6iW5
W74nu8mfS9jyqhiGq+9ci+1IbwofoTDL8iFRAvgeNILwDpMcQ5s5NpH11xAltQw2
ggeAIkyLDrwTJCyiP+v1q0gNNLBoFA3PtbwCyNdrodnMzbjE4730HwSjXcnxNMHd
TyJZtl09eGVmJAVJh8K9HPncfg1KHG+DfNXS2QejhVrCUw0J59cdpPpMHVod45BO
ASn/Mmnbnh5/fRFKUH2LMkUPyP9D55XieXHBfznzBk2qzksqq/nDvlLpmTYI1e7u
IcqkHMVW24JW1u37U0k4z+/WYn/gB17c6syrMxGQRnV10dybaDg55DJW8y6wXTkp
K648HZ7p7AN5IH6UVGmFVWJsIZyRK6sP6P2zzHlZ/CpdvuEo3t5IDDeflmejo98t
LCCkYSS7Y7bDdVd/m6411TotL8p2S8nQRX+4HJBjOX0376RBod6aLB7pGWYI51Hz
UCM1WG5njm5W2TKto48E6YIZ4oUaDRzz2hLE0gYGUFA8DKYSjPYj78i3bKRgwCEY
TSaSD+DiNxEPUaYPQjrGP1yLHhWqD6Cqir9HwsZdbBNgTsh5tm6XCb2leL4gYI4d
kfzI5ycPctpc0ldcRmPDIMEc+yCobhJV8jGau4o1j9/sIoNTX+uzwlb1n0GcTf/3
hXFgfArOwEh1v0RSQGlDHJXxjFOumVB6LD1kCBcX8Q85ou23xUXTQNotczYybl7+
BW1yixOpaQMDb4dmLe9lZhSGU9agfyMD8VhDYpWomspBRI0aTgHXPDMBTyfTIsCg
G0N+J1S4fvKanHp/gpqS8EXAYJND7UYeucThiwuLewd9hIv9UwtT9ssmRmg+mwKO
XdSAeTiZl0ISecHW/ggoSY0L7DxXdW1FGUkw14uNYTbh1RtW4PAcworDeMxTe0DO
R88bXcEHS6Hg0Z8FyUwzN5nb0aAUSzu3oC0dLiZdS0bmIuznN5YjUIYT7O1lfE9D
6wVBbouE9BAtHQPtzWcWxGHg4jb6RhH0h1aRqBt8x6z+CgGJlT2BsJmoBuF+13aZ
j443PqIZ9pXz86TcqgObGk+X26+Mom25CyrV3oQqMdsOw9R0629HGnGsvV41OvJV
oUUL5dD4qiLFdtA+LMz5JqGB5eYv2GSuU9GU/ulgaBW5GwZjeAbYFaqQi9AGHG4o
lXcUhLeC9QKqxLvL5a8tksyImbQlUPCtweustUgf4Ep3m/X/uHmVDmidubsZWrSE
Jgc2kdfMSqwykZ+C/l0aD94ICzWgtZ7A7wyuY653Hh/3DJrc6qEM4s2/MJJu78Re
sMgWw4VkCupo4AZ02r82fEJPTuQP8UAUYHC7Y7+bjWQ8yGcwdvJOCu7OiRwDSPeK
xd0Cmwd9iAlBk04mFBBztLmQRI8r9V+29UrN8SvuAOUeXbfkdbteI5DZBSjSAV7q
OcHTcmnONZegG0eNxfkvjEuxDofmtr7oLtLkeOceiDoZTGieeR3hrDXPwWMTPsRo
Dk5t7GA6Jk51u6eqFvAh6wL+ngLU/NR7cbS+f/hBhXleRGVZYjrSbZYLIbDqagZh
ou68AFlh2/IqCC+8Jzbf5LpTpIywCXYPtY4RqURjZsyepUzastJ8ChiZncvHK9W3
QT4//J194YWMzPwG+nyMmUsEbEDVLE3Bv4h9SanjDxwW69bWJt6sTRdh/rmZ9CvW
o5466i1kbByqber79yQN/1Anz/d8JfBAiiEwjtpEoiglQS9RmArwh4TsYoHlsmdr
gQsKdMeFM8k7v/BJPiEuKI3Gx5Q/lPNhNzbHD/iPEfoAB22pGR7kQjxLmYmbPEFP
0VG5GjwnLz5L7esY/LHELyEJSLZ0a4YWdUAU3fb6C0MWcHijir827h9Ln5zKGD4c
7/2FzbviS0fPBwwP6WbE4/ZJAvP9JzikCRlYJE1AMO/1HeaSQqCRW3mhDofFmu9Y
h1B6tJKRcCIiDZ0d5x24Lee7lYV8rTAO82WOw4uFoZTStCeYdYTAHChwUYu+1Qs0
qeZbYTpRa1eMeP5fD9o1I7nHYzJDENcN5NoryUIq+oe0dSwTTAzdGKc9YopJl2CB
qs/Rtj+fORVDEvMLaNbtyOEKBBN9kxbbrCaP68rj0Vn0CwfBLg1RPrSDri2ebqL3
MsfU5fSvgZewX36bsewbtKcJiVAugacf40SLm+1y71n0Nfk4xbV5uxdwGaeepxT8
qlVP/uwCpCTazW1cYTaf3BJjN3Bj4iq+b7Hi+Ech12nwaP9N2pJsVivkXIO7YtgI
uVQzNKbku6+0Sw8NtJELxDWR2o1J87vAIbxY7We2rIyDTx1hRlw/Cy+ouSlqw9fM
Z06Qhv1B6EaivYdkbC7pVfuo1dP4FbnjxvB9rCjXuvRoAHI0nJVkpMoGcsjrH/c3
2u020aEo3XCI47MBHyBv7UUxuBfHX1nn86TBihu/6yI/OviM6I/8CeXNHfMA6sRC
lyzkp6gAginWHsjJu9mD9snMHCAvXH7H7xuA2sNeGXQCxuqpydOjMVB7HFz4zejs
DV13Mk8POlvH8gFbMbAtz5/D0iqNhwX7WkGkP4UGo3G4D70tJrkuIlNZekiaq4Tz
KdVfroWjtXHYc434YtnElH8tXMF4Nmn+K9WhQpKW/yL69+5PeeNgaLnD7hdpzgwJ
5GLJpmXxkAmT8eOfwprbVRbtuz39UK1cbUcBfpRtzKWtSeTyX1+nyZzQaCqU7KN5
bMZkOI34y5K4xquwhuSu1vGfNC1xvteelSOMl63uMx08FtFUXH8c7FewfTHtyuO5
znN8ViQufGZ+l8olxJX7wpBIRIn5tvvFcNr+GO7pDLg32ZU9n5YKUt4aFfgQxpnu
LZA8SreipfwFPljbudTNXgHorlT6KUM7PPEK/GR7iUK5b4/fRvSYlk0U8IWH60M7
jITbMbrgfonwEn3PaYD+FIwoj+k/LmhARlhfDioQo/Lsgs8dHP+PMQvc5Ic8rpdo
rzk/X9qq0snhCMK6Ydv1ZKSdRXn/qYapLPybXJOUAiv+ySSZVfq4FSBBF3LVv6vk
xeUDfBeTf3Udq21f+EhZkWOXpolxCLvJxx04ywp5RZivF/ZwqkGY9roDg9SlSC5S
NfDncoQ64f4BA/NRTUGFSwRW7sDh7sGL2GqXBqa0OOgeQp+zCmZbxBkSsMqfGBcq
I/Fj7zAvvnJTaQG33Hp7fAJ4XaF54SBPS4aPxSkQPQczAvr1vlSHKFmy7vWaj3a5
/75U0JSuA0UNk5QB08ZBo7PirMg3Hl+/qfYzONOJFX8UlQUPrVR/FgZ0UpyKOaQ8
Sol3Syir5AwL/tEtkqECBGR++1FLd+i4rCwlOxG397gS1kdlTi2cb3W1Nk6zOxeF
0Ez/qLMBwfY2DxU5CyRTl8Uev3IGKXsKsF05CdBLEjUgXIG4xUBMySNkg2Ft0lY6
8at5m/syhWuUHewqGm5slEMFicXH2Ka3tlMXA8t59lB4fue5B8Jx17YjeCRufJxC
0c+wRn/ACppqNYHU+sost9B8fqD25jXuwjvaqjkPmqs3snn9Otnz6FfObeUTiKWj
mXLcU9xmfAgtaZwjXyVg8FEEC5XxUFHovxnY6elErVEDG536yMEjDG7HUBMBIo9P
vc1fEEGaa/KRt3RD2H6OV+XlYRFOwe6RXeg+KxrvpZHkbrPs971LPwdBb0kNbbHk
qkTAEfO18qzlGt5/nYY5qM9lKngFrf88THKFaU4SYz6J+OgFU5ScMk6yFMnJEtCd
p+yrwRP/2iu++o7VwMS8x5IJnT/+UduSkYLasa6KAjc5rGfM1QGEipBycHp5THqF
bNwBl2JYns0KC2YqFHLi2Iiak9UO1zNYGVrHs0k/dzY3t5QVYjBsoi6PhuYgcPua
z4kZRGqQuy8ALlq7/vEysJxZcLUG+HUHZH9gO0E7Kaa/CGHhsn8a23MeOD/jcx0K
FRMaxDf3ksYZVM7INmP1TTNJMVLvYN4PQO5SCaSLgpvy34STUOKji7f4ytc97Tih
4rHEnIQekQbBNw/uaKxb+FktTENOnkAMTC1J0Q8ZUEBi93vk4bOaCodJJZUYfs5Q
RqNRvWa0qRHpGovGgspLA362/A5irop0+IZasncKg71At5Ey9oWpXhujt3nztVlU
p1VgN0PVQrBCfYeQJwwp5C7kms+UICBr3o+PUpWmB5e8jQ3JsnxfUjbMs3yJVlYs
ImC0aD0cRv1PWin5AuTxlTlROqZxMUXCWbxvvm0ALmVIKQIQqVD4LwMdxJa3MuCw
/VeXZgDaEha0SLmTctEI4NQGlJ4kNPECYaVnqDON9FhaBbcWHPK1UJpJ3PPH28Qt
eOgDagwwNgQgq0Yx9/Kd6+0V7cIYGmZRD9kKWBF2fZbSZvZoHNdy8RkX9hEuvPlO
/ri2Ubod+o8J3RUFqz/QdKyZZRZm++O3HDPQmJ375if8aBlBXkozJZQkctBjTD+Y
dMnUihcp8yjT33ftrB69E73zyQhB1aTRIQSUtRBruN80v2PcYwfxZbGY3Yj6Gpli
9L2n6IowtoGdwOj26yVTlqyDSTQuoQEjO7OHCoHyvi1Fw/ToX/P2StOt9PYFKKrQ
kkUC3l77VyWtuFYJ0MZo94tcxNDL/iFxFB6aSiUM1SwnkO4kiXq1GZu21OsINNh6
Q2DQJurmKGP+CirgZb2gYA/yhoEjvxhRYh5gssQuLyMZmF2Y3obcFL9eQdLDx6vg
xZcDic30LiqNneeexm0kx2IkDTz7PxEEAzA5Q+WfR06jWsVUBHz7FebQJNakuy39
0V+RzvkjfcQ2f4Z1X5ywSum525Wpc31kCD/hdhgoJ9Jhoqm84EHb0j8UNDoTMeyD
PRrFDRY9bAf8CntfenVnLbvoTvQyPeBNpOAec+s3koXb1oG5aFWBFm9LPZPCy+Qv
iPtxRpoL+9/oz+2cz5oYhdRY4zIIi528K3EcGNCHTf97tA5ABoU+OpnxY23RDaFp
9FMulDvDGYoramminsVO//MDMt/a/8iyj0E5+Kkqbv07PH7KXtH5bkzIBBGw5OEd
YJ8RIe9lWsZXQretVayLskKn28gehY7o7wb4CGhKgI312XDtSRAYUhe1xAGzqIN9
l1OiPwaUDewo8Tr6e6ncauEK5oTIZaOwLojJrwz02xTXPl6VdXMzrduJzj7Uwlg+
N7+mwf4tdnNdtTAVqcXmm2Kxd+k3n4aH8z77B7NKLyJwlXUt6BticViQmPOT4mgl
pE+F7wi8J2ujWfsaTCAYU/G+52H4Yr+UoSTWG8mwDy96ogN+N7DKkTT4uB8fp6Cs
vxrqDK94JNyBOb51D3fzcJIYhkM+D+DcwEFzRrGP6ggxI/HaiRdZn43Ore1MG4tm
wVQG4Nn1CeYVpvHtAB9QqsGshzCar6TUUR4m1qX5eAi33wKxbgG2Akwww5UHR5GW
m0w4KGWiMHwoxl4tikOXTegJ+YY4LuESR/Ezf8FtcjV32B1v8zhbGrs9fAsCciOt
`pragma protect end_protected
