// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:46 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
mlhYE0MXZGHbSbmoM8/Wp0McuTC3kgqX9atgtAUdclVsYuw+erZYtLU4RbwHRv9K
CLsARLfK+diH+ldzsObfcMnGOX4LPDN5XHphj91+ZIVEJ0UDf0//jBf6QQ/b9KEK
szmxPUsHSB+bV9zVcMzK2Gz6hTxaxFKdxuUGQYisFJg=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 48880)
a80D3sEwztwir7QtXiDOWXix4FzWrxzz0jTKzD4nHPzYsndEDnulMWL9hWAfWbuI
BcjPzlfq+LvnVmJ/9q91Fw+gaSqJxlgEJA8AyAiBRyOUPSTl1kKfMhCI+RR7v/Jy
Z3d3mYFebJ5C+HaUcrQ3F31zfeMKRBEx8ZyIYtQyJx1Hg6EILNCAfCDzrCU3xDh0
9q0ggOz4im3iZH8pEHDW06d20Et9pSsY0hb1EcpZiul6Bcba+cZ/p9uEaYb683gX
PY4jeNhfjy69ArU0vGJMptLtqWlOv3Lrlos/xxAnLJTYRrmjE2tPlwL/Ns39fUM5
PCA6KwzztpPuvdrlwqFwrgsOHqbRGPzh/3Yc5FJxV+yItcuHNlEDpDNZi+ptS9Oe
HNWCKDXAepFiV+aVJ5DqkoiChUx+UMUYKXRdpa4wrtFQUh81QvKn/B0nNS2/Z73q
0KbZ4Tj2AMN1DtQADtNts7/4ct/nHQaToJwqMkwctTDB7sftWNTWkN+U2QtsjcPi
11bg6JzpLzhesn1Gg4X9OqfxS2HERK0VkrRMxBSfdnqrWKMbNC62y3fzJTT1noAp
jyeQWV5+rHjRuaUv8xTR0jn7ZuwEMk0kyjAhqgGXwM7vYB/V0OvBpiej8I2uKT4V
IXRKBYnqroP9ljk9/red4loE53kxPn4gc+C5y6T0J1auP7cEXIlQxpQhQlX3V6ve
d92ZMD9TyqkaHjMecsWOZOepPOERsIgfCtTri99In93h0V3V2Jc3Bwciy1m1QCDj
B40zaEsFF971GLptiAXN2lLsXVzikhvoJXibIwMvSeG+gEiQJAXE1CPGPSuIxvxn
DqLvcPTby6G/ossgy0NsuRmskXRbxC0LKilzOPrTU3DZ+F+nAiF17dAYSiLl7nyZ
TlM0kN/OavhgnMBRkS/9aKFG07BFXe5O78RZzpk3YhM6yoKKdOXtI4Vn4JCdc0lN
1ywHs8Ik+DQ3xmUbyMGZVRjmRww/Zt3ju1XUE1WajvyUZpd4WfuKQnfVr+qwp3gq
FC9GDZdSb/7jJ34w0sMdQiwGZxk5h1EHlUxVtOQA2YMRAYHWuz74nvkcW4j6Nqqn
+q4ZR8lnRl5uTrgUuAU93eVnH0DVQaczyGl9wUElJx07l6b1p3aeD3Nrgnd0AA0c
jVGd4wvaAKDHVjJjfx5zfBy+SFa0TrxzZY2bo4bSKBx2/TkgCsuTXsJc6NdAlSMc
9Qmr+HeA+lcnel3jOJfXKgaNQ5HlLLvPm38jqXDI/iOypwrMjhvcmbGrVCf9npN1
TWCBDvrwYgjYMte4jJYzqVzvtPpyvZDkefhkfWZHRhfRddfxj7xy7CurseElab3E
i7ASjBpbE5hm5Asf5Eqaz1aP8apXjomcjZ+bAGmjNpHKC+g1/jtosLtmwBd1/QSi
InrzpPs2RxohqKl41A+295NkFSVZ0BAAl8hznWUuRrWV31PHi2d/HPyqYvG4X2ok
dkiFOoSDicYX7gE7c15sgRzAwrIltMfuoy+LcAbcfTGuc6uaQyrkrVFph5nspVgY
BDV8tWK1S/GekUvEk8H1wdovZfgkgFm3Cd/3dJgM1TBdVavXCmqQBnuINs6VleXO
CBVrNUCtmlr+yOkk5+Jkj+GxUjIzpVcGIpDLaSBEM3yL2MZ3xtvYgaVyESL08g0v
QmrMmdkQNsu+PBN7mB2pWcS3VZHtxUBvqGnaW5rOQoIkR9igPBEhrla69KBWAq3I
MA4O/7yLavW9SFXQ7CpHyztMbVWzsVdNUoHdhtBUj7Gz6qQ8BoRZVQDuA0D4uIEl
Cd+VMOAd6u85AcZk54o473mjNNMDvKkRrC1mNq++MeKh3kgIdKgkgNhbSPqU2b8M
LLfVw1Zptq01tOH2hKRw3W+PpnYdpGa92Sxmy11+5UAbjWavtycl8T8oWAtwMFmZ
UV200p6VHQg5UnSuJ9n7nn21gZ3FP69AwwYJs4pEQtac3ZJtt7p+/PW77qBMG6kd
W4TkPk2w4JNINkEUGJSd4V9RxQMjlSlX945ljur6T8tcvxkuUJ8dDwzrT4tjX9aP
PniAfTCMsQFuc7lmUA3LCKCpUYRC++Rp29xz2EoK0xolwct9BT1L1kXdp07UCZYx
F7tGq1GzdVU/RuCozg0R1L6TVXNqPuwYkkf0smNr+xwWdR3h21FqjVdu11K91DGr
lVN9XPPcbgGVSRQ6nhs8Z7zHdJcfz+s68vZinmUhkP9IHnAfBKROqFqs7tUl4Edi
P6hrdb/foJvci5ZKAeFkSJV9UzBrAGShw6veS/bz5Nzd+iP9kH8Nb5CjDIIWR/kj
/4FPwzXlYVncqCzVPYFt19LXxg0YxdYs/PWO/+kBf3eBMovjxp6zld8OtFHBcPwv
KTca+yqzxzHjj8wcJNijVFyf9vM63ZwAKlmsyMj+iefN8owYyi/aW7Lpvud9SDV7
NG3OuFyJyT5LDmtdNmfA7dyNiP+ecD8l+6Pcc3vsztyAnNDBxv2m8K8UdbnRGMYk
CFP1eGLlFRk+lo4iero3owKX2uAwSotp7VlJeb6iDyJAaReuFvvko0f0bU4NlZ7i
v8vA4u+wD1i7JNS9UdBWES4KL9mKAroMSSK36WvTn6bCkEyksHOMZrTNE7On3stb
fojk2TfK++s/GTXW7Yk7h0ED9/dwxPfOYf2LSq6XHgUyzepaDRC72oaur3vpWhO+
pcCVNxAIFWbvLX6Cm5vZERLuAu8PzqIlNfdyWheCRdO8i0QKfZav2GUnUCKWyKTB
dEs2LNaInTwhGB8MmlC6Q3FS+5YzLgxhqSv4JdyWGb7atahRbbJeDaFOWpGS1m+l
vyIiMCzUYrAzukMTVqO//AsuDZ47m/9jzxKN4x3Id5J9GhzinrLDRvm2K6jbGSU9
xGCYfjTlDOJCAxtOhiM/YRLD56wryUZngskwm33/aWVHAbjDJ0nOKw1iGBvKrmGX
7p8tU3QCWfg3+bZBV0FfD7yYsfIfm/PprmwEzMZW0yRpv5EqhnRvbB4xBuvjgS/J
zMquvP7eJBvL7mpsu36i4dx7Ppc2jqA4gMrrhW94YjfZHgHQWVI2zUQIXqTMX9sc
U1ypvWG7P1SBfdlZV8LqLR6kMZiuGeERDnVT+iIB9pUwm9z1uIcWJ+7ZcqrBvhfh
RGVgRDVd8gMgusBgyicyt6BBnbO5W9uj3cGaIRYpOnbdDUNQboBSJNe1EY5Z5aed
58FDM5KvQKSifmAJUrroUk1+vp5g9zrO7iIiLT+VGVAzD3nH85w/0YHoP3/IMGtX
383iVew+hI1Xb9m+GZdXl9zJUTv9hacNz6UUnIy9gDbMrO5ra1g1FgbqvOb2Z6RZ
zMcYXYDrafRmMYsYGjRckxPnkUyjrbTwrdEngKBIcfyi31yexuZY8AMpll1aMuy6
srctVMqN7YceMz6/45WG6kov/nzZlif/cvPEwqktZuczVYuEOJc0UB+fjdqqS3lD
EmjZGZAx9gL8So5W22Sk6mqYSB3gCVPWsQLqyKSkVwldN/IUCBJnX1OvF1McPVzr
3KecdH4hHJ1owXNGznfn/HDnTbGWg7NvT9wHeGzTBNUYVzMxN0gwbNMH6WMhdCCQ
bPSHCrD8DaDLCL8qeQBsgI7fzT52kG1cIc4eJeAmeCMBQgxAZdLl3I15uAPJUU3G
XGoWtaKonUY87oV9R7i75KMzvTDPqUrJ2Disr2WFay0h8oC6f9Uuxh7PbfPeaRp0
tSIdVfR+7rEiwSZRTs0PmXs3z8UGSDohaLEeIrSQQkXlOkVRVcL+OYm8MwAN2P1L
JsFS6TxkvKskSOMTuV8lhCE+5iTj6NloOBR2TyNk6hQgZHuyxQMTnsj2uBkfTKkz
3sJr4EuFWgOS7PF3gTG/MZMyIbZAEp8O2aWC1W58NGmnrv7UESzoRpN4gRxzTQc/
ZScOa0meptZANXa5sR1IawPZyMlLoeuDetiGw6Qyq7sOQHv80A6wWnJ63xeSdIYo
iwol1ILmZaJYpi0F4/rfRK6Tv+fXL0e9tw2ylretBqpYnK6UHT2DxN0qs3syML56
jD0Pi+ZPv3aT7xphXqRST0wcw5Z1c+MCXzpIL76auTUd+57RNzeMEaSStNw22JNF
iQNRqzqWBp9cQmu02e4vW+vnjhY10AjfHKF1/dbfQt1wli9Wnbd2VBlq5/pOatUA
vKHt59C9fe6EGEWVx18+Sc6O1kQlYxrFW+FNNqsBnMrS5eIb2bmp8xuHaXk81X8t
7+BssRaHcdtwGvsUXT5BE6b502U0/vTDyltJaDF8eabnjFeHaeTEQz9qPs6cYds6
LW8MGqmui4CxuAAkRKS+JVcatZFECK9kVhJ+oBPA4okwUFdP7Cww8lxh3bTl/Q86
rkok25Fo2v21ex6WHbnevFS3Divld/od2kjVnwo83LZihiCIzgF8hJ9CinSwbmdi
KgNWdj/gwk06w1XQmcHd6A5F4VUVfoc90RXA+mnOg6ZGxGoTcLBSax5a0MG5KTNC
9q6eFYsJDOMQ2ZpOXjZ+7kMWO84zP8HlrYJUe2X78dBO+iOxATBgzLj/psl54WMA
1Mnx6Wj5Rv/X9ZwZa1zd7dLozvOeLBEzBHmNXZTiYiHBZX3hWcUjNO6O5Nzqyr2C
E0pGTsapRtgpGlle0f1zXI1QLv4JaRJenZlDegHqTFg/7JwlrfH2TkgSLA6PWcib
qxhQ858ZQdflXkoXGzPVU8FH8Y8uR2g4M+kxgsN3qcTa2a4gWijiiiaQmlVQQgsY
VfoWK8iYK4W20NgO3vzg8Nq9VMooeNyB2jqOQdF0b9QYtVBYjMTTrJo4ERZQXdvV
9/a8HzMdXPy2MUXtmZtBth82L2puCqpgPBX65pAyazHNCqOFjkeg3COYbzDSUDm6
QniSBJHJjd3yCNWVXXKA30QH52Xy5YbplnRS2AsE0VE3Sv2yJHChdlnCJCCueRcn
q3bfuHITx5bHM+sqpb6L+wcFDDycH43WA9qzUMmwkNtdAa6XzTzjP9dHNhN7pXlv
8Zw14oi/ZuJuddZqCrJzZwWMoQY8xmIYPCpt9JAvBecNU17GP40td11/MPmqz0sE
/uS5dw+xiQlrX1FIqOzjotrNVMyAij+aUuH6Q0UV5j0lLo6M1r1HIA12ImA6u90r
QPyE76XJ5K0H44hol8YNTrfNlzXhdtg6IP8KNsdbt0bi3MvaKVfBRqkBps5VIcvD
iBWjLq2MbbDdliU7ji3rK7PEsA9oEbLnmKL7cO/Sx6lAymI3plkSvywdr2QUfgp3
0whL+P4b43YnODpzrz4mwGMbte/9LMFX+KpiyxBocLGKq2CZRwrVGFOF6qVVtueI
gUfdvCOjm5e+STPrLTig8dv4ZnOJLw1obLMoyyRtqYUkG+Q4iYuao8uUVHJG21Tc
aYEadsPAIyarc+NxJomrevPYDyX8wNxOWWYknzJAXcMt6QySyESrhm0b/gk0Chwk
bN/2hCMVn6uizq8+Jem7KfZCK9uXlqvBz75v431WTPHT6JvnQDimUmFg6o3pJ79o
zVIlkqC56fvN39fibk71D67NZCPAQBaRTIOxMtfUeKbSs0Pndvl4HayNe+jGwAh/
g+h90lWKwQngqQJOjmDkWQyWwYZyQ90H5baEPNGZQf8zjYVgMgWMeDnA3SYb6Bdv
jgtEMMdn7qx70qWycBzuHNUwzcoYBqdJCZBHOKt/3JeO7tqEHtCj0IzEQpLE9RpV
cZgzYIpD6xDTMZ14tIDwQmPSR4FXMXsramK/GUiLLvNPvhxP2JgRvHzVqkWe9rbh
unbNpWnjZNDMNKxHilcCvLhYw0VMSN2gjqc0nij+I1ZAZrG1OF2KWER7MbEKurvO
1oSYoEy+NH/AW8iJuAuLVTSJgPzISf7sCSAzyh7buX1LWuWz7rrsbJcLwTuGoRcN
es+QZBpIfTQZnXllaBcCxNBV0DiKvSxCLRD7nIduOjcZxV19qOmakfA24xJvdIjE
VgI46/VeSYQPeqMtnTixK1/k1i5frUFhNqi7a9Leovav9gdNW10BgLDyfHdvCQow
JOdcIMuWLnaRGKYkeYRj0KbtXoALeyMxgJAfGENGQci6uybVZOdmmIASkTklJZ47
byATVtYgrUVTab8xIBDr90q7eDCuC8zPUNNu3B5fK+6SQjsd95/BqLBpDkZi8+c+
v5SCxqanZ/iGoOp83U49gTxAcHFfN/0ZnGcxnsu3BPchAfMAhlqMjTZx7Zy6NTE1
Wfg3/uUntI6MmqfEeq+t/ean8jSj+r2+pxyS8/NwdWyA+xkC7qYiqHJe9NJ/3D/b
uPk8wqiir07aXpcRpKC7dxNX7LlmruWlsFNZZapQ7jmWWL8ILLZO7igVbkepfDr9
Img7e1O1AGOIeVbIirlwoEFMvY3YjM4Bvo1oz3UqeBPTd9cxi/kN/qmuociW4LNw
NSY6rfrn0L3eyY+CedOHbzpBXelrt5hbjQLZWl+DiPCnhxS4yYqaNKm8FBuZwEvx
PxjbQy4gZPUYVbwWIObdtErFfaPsfA4ujTAWFpCq8C0Omgv2255qL26SD8lpYn9L
gnwNluxkPqpSlANJdjPlAZZWwLEQxdy1TdTQ9MLfvcNj7ZDiySY57tc68O8jZWnl
If46t6g7GGj4aq5VSCZNtiHnqXGwjW2u6ZKLml43gqw1n0UYApml1GBRSRbdBhlU
z1HnKSTZyHiNL8i0++CQU9XucHup3kgnVBmoFqqtTL47fcEeowaKxj8S5RM38/ya
tYYXw6HndO0mDQ+VXxcQB9+7SAGyeNfv0+JvF+WmM4TEhUA3MfiG5e7WA9KaKqGr
IsdBJX50HhgcfDBnx8KnPDUunxR/zFxrs0+tHaDJPb27dNOzqLGhaqyH0PVlvgQn
fpvbZTlMfClA83D9hqMzd9M+Mf9iCY+LPr8y56SqieN4f7i4K/VRdvtkIQJlfzWu
5SWfYHTKHCDbkc77bYtW3BGbZg5mteZvj/+2+RWh52+AULzrinq4XJzAGRSrPDiO
mwHHxDdttTsmbVTz0Pk1nbU2Z25Dcb4INCK0/fcKB8NHA+Vtqlbw9mLX7Prm18Rh
8YlHukjQ5cgnbS2hMgTZkg/hPWiI6tmUxAhEqo8eSDpVT22bcKKDVMZxTtrw/oYD
bGRk4+JcROJqBu5LEjCGk/CSOLtJnQqJxv9qwkQsvD3Q8OnzF0oV7Dx7rV3AYliD
1sfHddLm481h804fyw/ORtdS6ZpgQYb4N6N7xBk9R+p7217j+GRFwhNW9zKdisoR
uaU9oDkW5PaTgRo4pgZQWDew06G8MdVkk0a/6PJa4h/OyLz1kevNrB0FJ5ky3A4w
0rNiWHjSw8N+yXbV9XAKtOUW0tBbNNZ8Ig1V3PVR/ise+V6kCAKy39eab2C0AGG5
Xyd7QJrkVhKHC90npmf6EvBtw5JV7nMkoyZY1kG8/CnEZpHmikqDw3hzUCuP6gVh
1zi8L7nXqvOoaOyKPXYCBkow2sNizFr1R1/5FKiN2KpvxCNHMSQZUpCfKx37Lgz7
AcFgNkD6iDwqr6188eDYm4OPJTxqaXkog/nzozaW4IdIjaIc5hSRLkupb/srPG+s
8MWBLeeAXKIgaGSDbyHMlDwJLUbgz//nvOGLzZwz8B4acMqqqzoiHPn3fehuGpC/
tohPrXGxu3/5tVEP7B7+/ahTnJXaa/tzvuq+2jGo6x/g6pKtmPxNyznLm8TrEnou
8gHwb6gpiSrvJ+eFeK1l/KHOEMlsoXSu8J/NYTte3na+GuKsep0WD4cmYz7Fo4Jj
u3UQbsjSn24er0GsOik7trifuWNhh6wuq2GDvqSrf5x5EIM3CL88isn2a3Fahd+r
+qxLFyFTC2n217CjhyLpYzsJh0eJMFBPxuSvcfcG+JGsOLYs9rq0f/SupoFPn3a2
wq9EtvXwSXeqbGtU1AEMiBtgtPz4dVQuXZyYyPlfpSjwn4fkvu9QG7pmPGVXknJX
JOaLGISdx0QaF2T9YgfnYd3l3G2twPfJGpXJy7rwNnk9YAqoHAkvt6xQu4htpRKl
Y8I0jie8PwvUeM3m2c9CHv5PmzH2FCSQU7GnUwx4YNhzZRmlJT7E1l4IoC7OUgm8
F1e0y+WqgFILKj8K3mf2L8Uk8FipbT7OTgN5bIyxs2Wk2VUYHWBx4XyCd+aBv2NU
KAnuwrllo2pVRkmrG72EeUWBmaQl/aabDEF+1hxsAfQ3lXHJeaDVHEeugrXqFh0r
R96vfxDDGnN5+1Erv1QgNKtmsuCi9jG5mkiaURqdecUVOEfEpASKRsmxaDRhh0oB
b0WM5srcsjRJaI7MxkSmo1OinDGQzP9Q8jM0htN1ZLfSmx+73zXC4IetgDxybh5r
UP6Z3Usiw+DRRpmoKBc8UuP34h0u0CEN4O2FNXACrKI/gnY6gXY1F4VpKkcysgri
O/Rw4AChJw7mH/IIa/XhrRR42kCrDgGj+/Ac77awhFVjDpWDRC8FRRxq0FvZp6Qb
NEFGSsmWgFIZ0PcUa6yKlSj98jNHpZKcL63ZNqygM4fVFHMrM/+WuIEWnAVVX1E6
5r4pqklDO5CuXuLGKMhPFbKBrpOb1AZZZv1w0B2IvaHooFPZLs+AHucgWUnZDaXi
aalagt4fWTOQSkjKhFWYrS19IxT6jcsRZl6C+LoRgd0eyrD+CkVyyNvZTDGuq/eP
ozSHLvTRJqbXkV9kn06qKCzhEuVZ2YjVZ7Jp9i7xlUUOONxuzHTxazH0tOxodGTj
GrOKOk1bwV9h0CZp6L2Z7L5n1AHppSXWYfzzA8660Zovo0295sOI0Q/LuvWoEL4S
Li88PGgzlEP/Yh8TMzR+qBPsRozSx+G6SQBfqHvVXgIGRczwYfSi5CuLrZFbUp0R
f6o3Ub9cyd0GKzP5N4Swx9mrPPHKU1zLekSqkl9J/e/3h9BuWAc3Z5yMyCjhpaXA
mLsikh56BceuLnQNH7kJzmycwWxfCO1pdsGvXjJWRLDOLr3pnPMBZpNVB1dS1Urg
x+gEAKFycJsn7dvXyXbiTlAZOlYDHDAYfrWiFfHsVPxGCeKNxNFpC3z4RWCK1ygM
YuzgXj0AniLVMfwYI4A5ZIu1bBg2DP8peTePCiIP/0AiK57CkME1ID9o0pmW0v4F
l+RBJ3rtwyv0MP86j1bGtwawFv/0FUn0VckjQ80Yxmyr11+P2Dx6do91jHuDzF/F
wPuyuWQ+vhzrvmEMGu3Nb0CDexU9779t81aw4+EpLcMkoMSoCMvLVQJ2sbLaV24R
IF3LYmA5eaeYvKT+Q1CAxsfupC649QDb9YdaJ3Rxy5lhho1Wqb2v/BOV/0zOvcW2
j7ppXw4RFMId734VHTbQVcpFtER36we9YrHnQmMF6cp1jYU6SU6UtvqSik/m2PhF
PKVGsIlBXeKvI7rsq8/t22Pg6bTUXxqMY+VFjo9xRe0rUGcG9kECpTxXAZp1/7ij
bALaJMgpYLdkBtTwyzQ1lRf5LNaSyJMniXaeS17xBGhVd3HmH+lnSYJtiipVlSsu
0QDyVjZWLkfN6Bv+6HKrQHM5w83twPVQrl4IJKh7gzBaDyRClftl9gmfWIjkpzPK
i3xpVJRjNsWBumqfpMcYxsTZ6mTWNAGKzJEJWyWunb58ijaxx/5Ym2t7K0hkhhkd
rZdM1CDKWf4j8QD91se5eFJMIcLTQLYEp3V2NX2Y2EPKzDSNI0ER+6t18T7YO8FA
m7StuTwZiI+sl0SkWni98nKt6bNTA0Z56ffPObc2+zVQnPOVxdFWkXYMSWfaiFsX
3BLBvdh3slGytVD3lEGVCXpkEfS+O9uVJW7l9+iXGFYGYvRvxmKhKxbO597rGw2j
QFqwI1VnK++IWv9gRj0s+pEG9ufURxfrr0bzia5EP2Kb3Zx1hxfj5D1iHdt8k8aI
alQ0tnkEhuesFELJ6x0EU7lLNyr0Bf9lSbMl/NZ6PkUV2AO9DtQ4GQOjU+4tj8Tk
mu6XpdgkQMWD293TvuzYY/Y+wBX1Exg48+dngi2+OwKqUT0jaOJD+lCqrioMFRtO
OkhbKFAaZ4fcBNEjOUaE8I1CR8K3Mzn6bq0irMq+FBXBjQ15z0QL5IqC0whpnPiW
EgZGs40ET+5xpAJwkReYGK2g6XR6+gZAxo6DNNzTpmzLXZnHorGpppAOoCWThd2T
hVetsEu93xxWSR6q0JfhQNOWoH643G715+7DeOm7onTW3tAyOVoP2UFxygkOKjMy
oZb7RpFZPSDBW+1hbIHs/PqqApFtQz7/wAuCFsT+ZZ2Jrm4eO4jCL9+Qwa088VTM
L0L5Y22h9Z8/sM4Atedlh1BVRZan6i1/WIGdQXeUSsmQS9o8FVUMYok7ha8bZHsG
Wi50BVlMeq4iT+U5/wH0qXH+XV7xlOedRUWgg0ESvBnIO5TPogz7qJmZoaijuNDQ
3LsjtkaOWXcFEk3oLDKiWTE42lUDGJYAPC1JYjy2mulFaNXQw/9Y2SsgWKO4j2Yk
jaXYkQgsrDPRqA9SoHKDjSTReV42BuEL+Fd9HhubQJ7+0PHF+ock5ebwrgUwu/kg
uvNmydW6DeW2w6Wf1T812KqgYSi2t81oX3vdU4DZpDG38JAQgcwZ8gCrJ2+U/dlD
tXwjB/tNKnJsyh+3P9Np+ePkwWDUyCcfbf+1ggN9o8xw4q95xG0s9eS8dSo8ZLcR
2YANI/bJs434TePVKME+PXRDPqPW/Xx077pksdiXZF0gAVQOVz8QfVRfcf+IqJTV
ImVq9PK7XlVbKfcIJ77LkR7TYfZHE5nWtDIfoOS0P4H7QUX8EhVhepHCThePGre1
LsMW7jtiz63cATKftKZqYUHtO7oITWhiZiLNgeoL732abBgcNm7ekrfzxSZXgAXf
PY/YvylNyyT31s4wRxv6LL2B6foL2oP44ownmXXAx08QqoAnYInCkPiW4ctIy6cE
U1ezP5WtNXE4vTDJTRCQuFnewDczLgDKUnEDdV/x3TSonTMg2FsO0qJmhlaWGj3l
va0z2QMAPxLpRLLGP5UB+BHNIzMngTU/u7Q211U0tB82Pn98s2ZkRjmhiZFGT6Wc
O5RbXmvmGso6mCU3BydRaPZqH+l6YV8m6Da95LmvTjpZA3FPGuPQZn8kaWnk+aOE
DY0NZBxv/KZF6UWJzEMSblkR223+YiFO3/LEulPD7UUlVZjpLhhEdUFI0cP0SnKi
ykl/UL/hMfUxb+YS3h4BHr/W/VzHnUlZWafe6qb9G583NaTV/3jbfX5CfpMXImr6
bvn0jw7qEo2om8nWkShnlERQhCbRIfxqJ34WXqCQ8i3U6z6ZP4vI4qRgVgSBKj+s
bBiVAL2iGoYtAHRkH3JXYPYk+Z8WmZzPt9g9LnPjeDg99RG69gLd709PWf+eR/Je
LewSQ6391zQkfBeiuRgI83VCOsiasMdTxXyM8a2RLjxfs18qvKrX/pv2BywfB38g
/KdT886nEY4AjullBpljMN56NcbX5I5NL+ZPLOK4Zm3fHEQSg/2+Q3Z0tjxxtRon
VFkmtEHiP+AVCZbhJBt0cyG8Ib+AtcmweaJh/cKeNZE67GCUev+BAeZdQumfDOq8
L8e8VvnPppBsWuKrF0dHkP2j/9Aq5cMUv4Zx5J2Vwn/iAW3qbA6FWraeo527WmGm
01ZYEhzUrbJcYhoBgTT0qY4ONTnE0C/LkFIlQBQTB6XepQCOWJtAeDpYhm97SDBl
vKQh6FNOIsbf92XadPyaWat8r/Bgmt3HsxjCu7V60XjU9fKKeEzX13Q4StoPn1Uk
Q2p/LQYNFttScum91DxicJbdT0jJ6sIhn+sLjLvJ1M8I9UHUs0aoQBjCeDz3HinG
i5NFj8MKYwWRSEy/3V7bQEBOd5S/+x9OWFeQe+SCnjvZcqP8gy3QNNlW8awE0Z09
K6uxIC0QBHkPx9wbz7iU/qPlFL5T71FAyN3ypITTKXDfHfkx3j0Y4AKRTEb+WeAV
G1XGg3hyHMN1OgLCSy3w+ExhSLjHFVYKut5yEPD7igjnRx3KGT2aSx+HZbDeHFBU
Vz18DmcUGa24uUNi+EixTIsua9oeLIfpIlGw8OL7L1m59IlEI9a+iSwr6w7XQKRC
h8mWxc8PNg3oTvwQNBQn1qwD6F2tprGJpUjEeXe67twfMhxqsE82osJZPW+HFa6a
DBXrI0G+wiKZ2VP+0UNWCzZ9Nt94qx3wo3LTt+wqxWdvLX0uMo5COvDpWZEuQuPk
9+2fCdEQMORzuy4YuKAkq7DdSk6o08feQOu2SliqGxFbG3mo2eqVaVxt8YAs6oR3
xhhDu1pe3ZSj4yJE/Tl0UlmB5IY3sadxuZeOXe9xP8EIyDFTYUH34UyJM/bcZZSN
nB18IA571AL4mhq8eCh2PWKeF1bKsqErRLlfDhIauK59zw6d+MTwNiKsh6wKFCyv
JJB6dCHK01axm3IaR9W2KaQFXctSCzR87svmbFzJNCOJTkgtrYNL+S4S0efbwjYQ
8YraTiiTaudEsm72eHUqWtrh6lNI8u3lQh6ldPWY0fVjbYnxYBKcFqYv/nHmlujU
btWPOAbwLp631H4ON+UtU47i2kplnkZ/7KNiUkODjE7PKEgynyQb0qP7X4i8fjpU
E/BGOWQ6bgHi8ChD9A/EEmXwX3QuR1awkvFoIgs7pVagTfscBsfzW74uF9qlwOXt
NOgHd047t5mwvJ17sDDwDbvL6+9PHX1j3Ou/3Jr0ZbClg7l9t1D9gIoKloGxfIDZ
jpkRmD1UdoZONPWY14pssaj1T1E6gOYUjoz6RJJ05mM9V7oRTbuf64kJS7t3/sqx
O59Bx7AjokQmmIrYDzqW/iRmhGAvZkc4mBLAOBuMqZo3JeEy13gyjOy/hFA1oByL
zu39c4pH0q4IhwTYOBXn/Ii8rSKV6BEdb0Div7Akn5fSaX/0tDJ+6J7CKvEEqT47
/xwqN93LbvuBPXQ0PfMENhQhpuKWXxpXCWUkfXTUaBMSdUJLaWuFSCl7FM8er27/
AXNxagiSYTo9s5gaMVXwewzppOoYbr5R6/sITeijSbIY94ZfD/G7CB342KkIiy1Z
WreiMT+f0FcivmVu6ykl/goOcKVFViMksA1Mi0sy/i1gpjmqQtxB4MUvoy9RIQjt
vyq5//GLYwmWoUK7kT3TbgSPdP+gbQxNKA5kdQliOEVisdkbycG+BRoK205CF0XA
Vybvdd87g9wRbTlfRHuk9Uu9YmsF3pzBaH16z3on6fEvic8q+1FAJvQsRmxhh7U7
1zJB7B/KjjKtfZRJDQiKFrcqpMWZ+wpgADjWjmp07vy0dTeh6VjlEHR19F8qk77B
AEwYGv2oY2KCaV1LcP68+dqJ09f5zljwSPTPyuRE/XpZHDWRr9mcnTjXXtkeVviU
M/Wli3FhBslD9hT4G0iLaakn+sZv9m8P5EI2lC6AKyy5aRWSsmGxZV/XxeQpk7dK
kGZrBUCuzHUYS5w5mVcarUhzOPpCwO5ANhvB9a6TYRuvKrP8N2FXjbW7bO1jNbAy
UGpsdqwqG6R14DhEWLoT/qI2q5fzt5w39GdHzKRqqyOk/z51WbO54bjn2OA91bz0
C23ZplvHXziuN33FLMygIMa/Kv1YsyMvzSw66aj1Vjl7QPnE4+l3F+6LUqQkzeYB
7rfkfwYaCyT29tbVe23quYpk4ypqo1oFpyKWsE9tj0YNwHk1B+e5L8JFZb9xUs9c
ZjcueqNEygWUMCmAiGQaRYzBzt3nT8/n+mCRXGgUBk0nZQJ03l2/BBqfOHHhglwF
x1YTs/8pmXC8v7jaJ3a3Lvk75zGua47SiLgZVssTlB0hjIMGUsuSAgDDf9Ds7o+i
dlHZQ1YWmgpCp66s2i7zvva5y12Eih0NFLIuii33A1MiBugRaLfLWhnZ2PjO1Pu/
nGxi/oGAQaBZGOnhpoCXIYD4I4cShNOSJEROuZCBZ6A8pNyvXuD9ILb0kN1pu/CX
aRNu+Cm8E1aj852MixolM6Qo7Cd/axRngza58d6V74/SebKRUazMd2BPh2+Ojq9s
dmnTjeXPPQ9R1J0Qd3ffv2bAyxgIJluiknxdz5oFG6JLPXYIPWtM93bvT/vQMWyk
xSXNzh8ocLFLN7SVTS1UzejQ/e/nkgBQ0UW3HHO+Xf7tpN0hKVBj/mO1c/ZaANy7
OSFL/a6yLebSys3YLhq4E7/+DwGpsyyoiYjdORTHkLOQxO0PKxwr91j8ckNJo28F
ztZ3FKgWcCUYwqrv/LKhduS0mL1nOkOqj69J5adL/cvxMsm9FMIdC8aLFE9FhSaI
oZ5fOsVQaAMAhWpFoIACBWEB18apFLfTCoy966G5Y/gNCfin2FSIIlTQYQaP94Fr
v7MZitAKee3zUbWPyyCgIf/1DtSsW/aBwDu9pFi0zfwPLgKYm125P/eb8IjFekfI
bFFk5d4J0bAtvejX9eoh2CHGFfThTKZE8QIclV3WgVBQ2uzbutfvvvjF+eohYdOe
BS4kV4KbA0SQ9A43RKONBsh6mwkXuWdYeuU48XxAAksuZVXN1DcCwx5o9+yUV9s2
zEVvpCFDfgphY65tF2dmCLKlNFZTx6rYvGeqRvnL1h9wUDbvoirM5X+nqv/wArhl
zoQjGKGrvVFhxtUTfRQ46UwhH3JvhA7e05XTzAdcP24RxhsgYm2DUps8C+g4NQsa
3jPyKuRP0Vmb9xVK5HWfUaG9fWWjX25IReMFHdwOKhHJx3ED9SKjcEWsb3X0mk5x
9F7S1+IizX8qmTCJehgq+u+F+VjsHnPj46m8/cwbwK+I5/RKpb2EixgLKQLisQSr
8LfDlCuLHsCrdcPfth3crb0sNdD57c18HECMlKewseX7vkW9J0/onCUZtZKeSQJ+
5oHH4ycvAGF7fnwOkAns+1v62+DzG9XYsEWKeYM3pFnttB0b/RKfJjErn3MSTnfA
hvXeqHRkDP4xvqkW7kdQtT32ryCWYb0Kazqon2hzI1iac7nySVUnu1RI52599jDI
hP0+NUFwtTwL2hA43sB9yx1LZzvtpG4UaWxImH6fGu+JB+jrRopc0equwtXZCP2d
h1fl3iL1KjUyNPN7/b+nXjTnEZG832hv5TUyy+eU4K4UpuUosiwglh2S1PKXcpgo
n61E32po4lJilquH1dvAYhHSNLFWJWDZm8Xy66uH4lroFZFKMuYacpi1mpt0gj8e
g/cYndAtR63du6tAXcBpDKrDFK5PFJk12llhjm1igb3sRYG+dNUFa1UGtyPuoXzN
rj5D3VvxKNdmsV4OoOKoJDiQUxrU5IaeE4Kem1VZRy4h1QuQokdJpH79xFDf8BkA
M2vL4Az3pjrJ70yYJ7DIYuYaNkhLrGGlY52XN/JA4lIbat2L1zEm9jiri/v1Eu11
35kKNXzivNNgsxouE4er3SpR6hPvuX302UmCCRhTWWXrKZeSQugTgnn3eJAo1zeo
NXF4FsocUcYITtIWFdoY5af9LEsi9JZxzGe9DEkzFDLsRrMfBxSzc9rWSY28HplX
N3jYCQrQ33S/Rx33w5L4QFOqcP/VQdmuSc6M/widkcHsLhUO/uuHNj89GnRcwr9b
N7+/kfbQLqEsqJGfVYtJ9zfxgLflUd7wFeE4zEet+g2qRRqmwRHU3xEiCSiI/hC/
Ywitt7vgOVVr2jJa4/xV2QVcDCX/KGgs4FZEvd719BVoxM7w1P6KcRh4GAUT4Hnu
6MDSLNwo1uVXeKKTkL6uFC+Z+6/9hDyRePqkDDcJT+GjCCyvykGZeiQyj2WdlDzZ
lZuQJyntsXTFF5Ehm9Vhkx83zsCU7u3qolFlKrr+097g4dBMDATz3oX4zY+hq6Vx
9wzRmT7LcI21vAJl/5OSGMCWFI5woU/JFNBTXZMaKlk9gSSztYOk2gJElRSDhOUq
kiULf8HM5cSUjoivRY8qvb5kvpYBcb1uNf2hsLiKE6A0B7eB7vWyhAiik80F210r
GOR3NcaJNMobCAV6xTuq3adWVzaDHKoWCmQTybp9eQDiMoi56lmd5seUy+g4B9mm
jascFi2aulPXHkphbNUGr9jSGaOICxSrdkKIJod9RunTxBtAjyAQH3MaerfnR6ZX
adVRTpst+lDhE53w+TwNZmCdBlQ/9HT9AoGr4Ro0TgBXuY0zupCtV8Ii9ytNU58A
le/YGITWjt4UBkT9981LQH2Osl9ucoOXgvRuW3lmvThE/BaOmG83g8HAWozz2JjB
vBSjEj57xxpa1KkOELsc6umrvHmoYd8ThETLWVj7QUgDyVPoybbsKHEfTerbFKpD
8RcxJ5ESVO+oKJUL7hM+TGjcWegihdR/vygGjhALl6itSKqcbwpWnJHmKa0GO7oM
hZmLdKOccGkDHMEPHyokRyPKeCCvYj3sPRvQr39+Mcr0v3yzlQT08rD7ocSKt7eD
kOB+15R/63J7jCW8LrGV1zUQlepk6UDyV4TUtkwEGi9229CsPEbESGFYOu7JNsAw
DbhVhQ9zTAUUFrZcvQTEHcr616kqgl+JEIIwLaOGY1LARAaZInpRh/vJQGutfx0F
WyAXEJvErf0aIYneYm9wVyXFuj+1/Tckvo1PE5aQJVDEtIaaNy5eDfcabovg4fe2
4haynhlE7NmoKiyhL1X2jAi+Za8lZbWD+MWHAFeBDQ2NagkzJoIQb7mGWGtYD0RG
Ac5Wg3DiN7Rj5IxT40u0uo6XXV4NNUa7X9kSby69oCu3G8Ba8tRIFNDG+LRCTGnr
2utrIK4UJyjidNlLURtmW568UAQxRvscAc/NzL2kLhvNGeVZTua6EzndRzq5THQD
tR6YKVQgf1Ifnbmw9g4m8O55VZx8hmEyspIy05ZlN9YKe+pXdISE4OX0TaD9Fi8B
5nDq0CR2jAzonJQ87dGroRPeic0r9Fiz7lezPrllnhMTX7bm+4h4gVQj4MxHIU6n
fRwZkqqvtTnSE2W4vtdn69+CK2nvCklVNeVdal9njNezzh5ApJM1378t1r7lfjDx
rk9p0POaoY01aDWLYdrow6NPe09n7ahX2WDhZya8MqjHABn6w7TES5bRjZwPTmJd
vD8iJ9jcCurYqAMHW+6+GXWQstwnd6D8gVccDRhOhHenArQT75kkiWydcQ+Xu1MX
QUSW0fndnKQPXWe2U9MgYYJD1xhgIwQ4kCiGgXLCxCzbx8AORng+2QMzn2CEplhu
v9bW+vN2nEeNmMuI9bKdlgEQykRVyhatvUT7MYBqtNF5qUKe+iO/fyw9vLPw+MY1
C6CcSf3rI+Z12I0eLfHw/fZJkHrw6St3p6GL/V25gyWECB5A/hjNOsO983PRRPij
csEjqv+lraJFfnVE+3gF2fX1HtB8cm/yJqylF3bxxElpF3Sd9oiBzrKT3KMyYbsZ
uy1bFVzwsNBluz28pBuZyB00V9WUD/joAAM1aS5NiMBoQ2Q6Xat5dMsGaMIDcz1f
j29Fw6wRfiQQ2JicXdI8elWiPvphrAGDSKZ++YbY8yP1CQ0Bvr8Z7tDC78oIx+7t
V+wmF1EaeASuYoTWB4nVp2aERshhqm7Wi4j8YvMaEVkC5FFHcIYJfTyOkIoHGzjp
GdOulBMGB95NFIXdAOMMyWrr6QMfaQxfP2rbrjQ68f0NdKX86E46FfQvzlsWz6I+
E3/Wd9Tuui6WGfawi+hVRFIANS2wuBuB4SoHJCWGV5IVoh37T29pzbdSVvWOnQw0
yvJ66ONNB0ETz3/YNEzTW88MxyfEJ2p0z0c1nrQsWT8AenGpuiYFIfaOTIRkIjVM
MJ5ZGPNMK7pL1rrixV8lDY2bVM5B5VkSSWXCGqbF8HsxQWTn/l56qcIVWXqon3ZW
/8IxWvIbIKBtkM8BrfU5rzkRr60Y/pzPyfw1w58OmiQCZxq5+SFCxFC+J/Xm87Kd
XHsPaqLZML9OY7zyQAUOBOkiT+85UGe15+shxb9sz2WaHTgjH76ARfc1oKJUXLw6
lPpp2OQqTeCesTlKlMNxfJuEEjW7hdofQOu9X83H4E8vgCXA9UyWA8p1mzUUqG6z
qqwPEdlixrdOnrIWljlVsojiRdNOSYar9tz/nAFhsIzggEIw6ekTizGbLuJb5Lok
MEL5SqKbosRiOMg2sQg13SGcGv/Cx4RHj469cDvwo1EbWCbfadlbBYyw9kuChThY
bx+zmZ+2cIRZUCvmPdrenHRnAnPoYNjZD0HedFhmgTb3SgFHbHPF0M0TQeUXmhA0
DvimLAyhnMHOY6ErBsyLeBX0tEZc/WJ/57lulUVXFxblXGiwcdH7MPrrsq/wGwfN
x1S4bMwn63b4O9gaWns06OYjrLmKgQ2Km1/oNefN55O7GEdvFWxiSQoa8SlM9zOH
Sx56mWX6zwioN2iBM8HM2smo8ihmosUhCobiY6EP7IXRIDxzRLrzZnDP4Rj0B+Zw
TZ3ZuMLCXi4mG9eQqYLnCCElM6j7wn6kPNzdP9gZ97n181G6yte5jWuandR9bvYp
jg5JIcLDA4UvDhKguFzgwsnvwV0LKhvOES1PwsEhyKAEm/KyQpjdolFC5vYg3rmo
vO2VAI7iX/Fz123GyY+SLNCm9eUlEcuk1PTw95Ww/VZUp96hFEYDRiCjG0nQk+QS
oXWDUDVz3T8cTlKStWKtyjT2zb6UtTfcCZAyIMibrPGDmw1CkrJf3Dx31mLDagYj
tpAWrB5MacW81KqY0ojEWXX6BVciPDZJCn+n1Q/xKiAVc9hglKHaQA+RUpu/MT0B
ZRzOrfduVG0yv+QEr6AzjH6fZ85FPbGKOVCb5ArF/Fd7ZdCst843M7Tb/gS/DfhJ
jjeT9MmwimD+xmbtxGZlLLZ37AuPXFadlbJ9Upvs2fCEm4Uiirfgt2fbkBE2RiWC
50BTNh7KqFYY8b4T5XCiCWIvHIOuIV0YG+m1ysy3PGY2brFp3QA/5BWV/6HJEMMj
HsJiLUyv+WIv3TLtXICzWmG1Er5Q+CiBBtwZ9Rkve1TE8icyP8YlVIEwXSX5t00J
EJGn0QF7UWr5W8c8U9PoLlCudZTcEPBV9Iur8s4tCsOFx5oRjnHPRIShuoCStN5S
Wn1kU0V5tQG9bnAWuLvHIGZFOlako3OfeGLzCb/riYwUNpkcsAom/Bm/ttAPeEgK
piiFsY6RssiRVMd5+mRG0cyuh62yg8xnEhOup8PBgel/myJ0w8xlgBImIpDZYCNC
MXTSyQ9rt9WuRjU0sbjUHlTvg8k1fjN+vB9NPnm98VIUXqVpT9H+SF0FsaQe0kbd
BOEtzg1zio0SyZ8X69qyr91iZdnKWI2FNJiDdQYSJyxRiy0zTYOT6EnVWFd/Jume
Cha2uVEjHZCya/3+oUKa5V48nXLw56k/rW6SuOc5upatJIv0kOX6B3czcWZZ557w
Rzc0nPi1ZtLoC0/vKM/Mfa3MT0urmia4/5Ua5U1fA/txQ7KOOOkmb4hZiadwLFr4
XHSdVdi6uxjsE63A7V69uyMXquGRPldxEkuytUCGcMlQco4AZT4SbAs8mBDHku64
hlYE8J3oxuJvsmoewBeWHz19E7fjpEiwOkniEV0pWJyw6H3m3kHx2c8B1vBkA9/E
hZEdpO/GVCvcpBptgvsdSLOVxcIOWekcOetvYQ8kx88Ka3aEYWcWMBJ7kfcTOuJA
/+xtzBbqH1zGMcAeVrPKPeJyJz93wt+y6thqys24eJiPOIofmFjgN67As4SY9ZUL
9syDmUfGJj47A0TslyG9Tsfpoc0WShsdl2zhAY9iPlSHJs5jkPQxPlu6IC84sOjZ
eBpXp6DBuGrtYNxxAw85/TW69rLAZnhZRFCtHFeuAmlresuWKExj3Z2FWWRpvKbx
78OHOtGwRa+C0NX5bQ5WVQXtQJqxdI4NIjPrF5R1jC+avFO0J73emuT8d841prCp
0D0jbUSsgzA2PTJDB3bChnrXbdwXxyJryb9ppCUyu2T4GtsBmChpGRf/QbqYFIhw
mw41vsCNLHk7cTMSI8wJSgqsUEXNgW+Ksrpp7YGcbC0/QycUipHFoOx8iEG8nhTn
OssgoCbbgBa2CjDxgsAU4zfReugUxP5PBX1X5EOPzc7k42MKVQ2H2Iex5mjNBvzH
S62daU2iK8XAdfidR7zpRzKK2YLhRSdH9sqI04G1CP+dedShe3fb6O7cX2pBj1ew
jzGW0pee/GxqpfnTiCc13HxfOxoqUp/UqTM9Q3EPNr2R41+57nF4Tuw/2cZYJQ81
E/JM2SjktNS5pArisetT3fOgR+5lJyPOndhSe4tokC2qDMrxvjJHM5shjLy+Xu6L
56x87k7iM3nOtaNLXAqVkGXiA1P+qwb3mxc9uQfXJGropO1UF5QnFP4og9EdJTg/
QBlTp71F+rzAUUmEpdUsA0XFB9RS9lSh5kjvM4l4FGMUT42WQ+gcZNtFdUSENX9N
GOmBqrekT2jK9x0UefvbAVBsmfxDNM5m+6BaYBADykO98EVro+2U3KWUH43m4bxI
c4f9YMFfERP0Nwj/tx7WQ4L5iwAhk3rHDKwrtiklP7D/ytbkVE/y7pUvEhrLu0+n
OkrTMDP+4a7W0LjRf0R1fs4Dp32rLHhGUpT/CWwRFTsyfO2sy872ozERPryRVvOy
B6zTIM4IefTj1Fehkf3m676qXNsOdD8qxZLJvoBJgKAPqxHU24FUAq4/sZyrkvUV
/HJZA+2qi+BP92vBhrS6fVJWppJVqmzqP0rg3lx2VZWE7wg5pqVE12rXzbiC6W9/
O6f9aNQmCU1y/xpaug6BXwUJ20vdW82wApQpROT0yXnPyCsBe4ssgUO2ubiqwzzy
p6gbPo/JgcsBl8JsNSQlBrisgh4kUrrcWY9nCeKDkgOf5rVIbKM88TUpyrUo7TmF
jun7hjmkHi/aE4EYcM45yI3EgbPdyX33OHqtJWsiIclZ7A5VZkMqmAbcCzfOWAa8
i5JUOp/QaCgT6GLZy8ru0tfZHluDNvYABVRRhu9bMp6gIjgWUJzr944/ZHk+zT/D
rkfFBo6ef48dI6Iz66LrY6frLVrgvIsW5B/s+2xTJaKsPw1AKZVDIVd27mwjL3MF
bpxtAN3suzB6KAPghB1do5K3Wk6Yslgj5LQkeovy1hMxyoWok9n5Ru1nz46paKN7
tg5VUc1r0Grg91J32Jm8UjRVmfeY8dBV9aZmlaDA7yLNPNACw+9aXhjvWDbOrtRq
7L2ziMgPVPzg6zwIV+0UeYWTrRun2hL+RrSpG5pq5j87DRpjiB/+fc9bx+LDUffH
A6tIAoet7xT5HEmaTKhp92DX3ENoCAm/5uOYQ0mR8aCDkVt8MiPIZY6kKQg1lNVm
A7/1akK/gcJMrd1IouTnqBL3ircK7g8LoC3Z7KnZww/OO9mjcWR2lAImsQX9X39z
XcyPeKwj5l2mIKm6zkKrGFZFdJ6hoJMPWjlx/Yn9hdgJA/kdbLXwDYVz5GuSuf2y
AFT9lR+cwGJ0hWR9nVIrFqyXebj/MDsOBRurwGEy7PXqoCUFBXc4n9/pwO06VkX6
mUlf0QfAylCqbpTFFcv3/l+VaAcCqBxsWc3P4k3W8PSgQ5oF0CL1xeCbTkWZLL1S
ftp8yPi3ulrjdMUbUCDRKuaSsTbSdLGDw1bgRl1Pq2ZfWUqUJlvghSuadL0hKEwz
B2JRI/wsdEsXwg/ECSdPVCZVBqQifbUIwyvS8EnMGW79RH8jHshD5/ogTF18g3ba
gbX2g4YzVjtQLb/o4PMfNaaQ/nq3nNXh4VW2G4GSBkYEt3nmxqSlyf71ySxsbcJo
NqgEIT/DbYzS28Gdt8OHGh6mLq17QLZEUrpaYRi4vRHUuSj1L8gztu0JC+NVSsga
FYlyuGi6t9oddsfgAPxOYJZW+PfJfpkUdUQKvw0cH03hiWIfCnd4IZFr6I1/VMe1
lhVupyyl7GuvoOzCduvFbx8bzubG1wTumSbqFYmOq7mPaIADOawtWKY5ePNrfT/j
6luEEg4ucVBX71E9VtURXdwg6Yhwawhcz/EWtIX+VW8XCmCSvB2JDld/F8WIm5wk
TRK1dpj9tLagiZD2TMVpy4swCUrBRmmQDQB5Cy0yFJ+UZYpoleWX/anHKYHIY21d
HNYrvTx+ngAYvyz682qOm4vS5V1XARSctuk5jOgnYUEeOowjiH2nXlVJG5Nolbi4
woqcFiEcLJX6bhuDLasW8OZS/mvAHE7oqyoqTlFDv0Elssp86W/4v5VRvFdwO1SB
wz5xZoVPHh4eS4HdAtPY+JhVry5M+KKsMPBeYAG88xqNYRTRUWVSJwWTyFvEWNEC
b0uybg5ThA20UwL6jhEePiFp1VR43BGKdfrLAXYaH+jqazBED7jxPtiCIFzFhQ9G
CTB23/DQbmerTlgOAqaHNGX3yeY1cXa5oZeFIe9p4uPt9Ru6p0qNPJz8EHkhE7dV
kypSFby0xKXhroO9/stX2gWRDTMKbhddFs+nPQnW8GUvzGk8HPdN0hrJ5D0qXtmc
2nTfBU3Zg1Na00v50Sf6R/QKU66kH6gLsI3xjw3A5J1XJzKZqkHPlUZqjzgUJwZb
v5FQSDBJnRHbXNu1MyU6m8DHZocxzwzs9clmGecNxoszes9eX9JeiNBayO9Q+RHG
Nxj08hHrFgbaXPKsG0v/xr5xmiCAT1t6gQCxQ55hsI3HKYxoI1HyVXx1Q2oUb/+w
MUhoaMBN3QFTXLPsV9ZMqVdLEo/IA1MX3lFwtglTDbLUqKtczoqi0MckkiNYHr/8
yLUQ+UeNKUeRSDgl03j75nkfZtpNaCxTsdoDYH5cdcGoS3y8G7rKVp0db0z+OpK4
pQQOBVYYrJ1rqr1IU9cfafQ/qT5rg9KlIWXOV7AJ7NqViDChNqgRJ5SiG2DEoMYw
o9rkBRyF8Zxy8wep3fhlEr8RAdGqRU7mp7xFHetUt+e25Mv6JukIYpRW+TARG4ZC
ieLo3HqbeNbsi8n/RkvU0mqh9eM1u1EQfBFzcSGPhLcFT0unULB5mzmmcOgwYJgT
XvTKx4ftxokMLnmzWBmw7ccDMR9ntx5vu0YAC/diGpxCmr6O7Gdyxffv1eZPQImF
SbVfKq15PTJh+joSaonKc6aCdv3RJTa+ZUGtMhyvsb2N/71Or++G+t/0KYS/WW3L
+UWOT2+iOxpHpQUPHS/AcsV1KaqsmVxk04NcXNXnoHJdETaG12LeCE6U28c7mXg3
FfwUeLrNkOM/GtjQicT+XUMFSOsdz45DEL8+nQpPX+aNZSxlonBTEV+d5sfYYF13
4ERE2zRIvN/jdHPT5ndbMcgn/0gpngip5p5hEKMHa8nOYxnWab3j0jgHVU+RsaZp
GFalTXftwyJXwPTwK5enitF98N5dx3JQay2tjzt6SNhAK8zKDhtNAyJfZJ6IkxxE
fX6moYZpBsvMqNR8WbwU7nAnuRNTz1YFsY4+Ci8iERYlQZTTw9S35pvBOFYVLZoe
dOqaKFRgm6t08mn/5THb5lhl0DJ/56kEkr8K0tMUlmEUgEoIv99NVx3Zqs5WaQZf
edZq8NEc9Fz6dEZjISPX4FeRSvJjVraq3ghnxKdHsdN1GbyFH1OazO1rkF7IhztV
vT7Bc+HvX1UOITFXQoDgV18ZFJ2FIfEGndApgwRgMC/eNXGjhV5y4vGRnFb7R5D2
6lZy9grpKBYXvLMpSMq7GJ7QxSI+U/8kDC2lyd7HNRJpaqrNs2AUcnWHNsMfHFr8
wiJb0C/5/0u8nMSG4mpfsXdIVNb6eCpWHn+lKOaJsmf9A8VpEr7/HyeifiZsnKWQ
D6lVZy1XrF3/OpdtWpr9i6NpRPFIPN5PfB8M/zyPGn1LY9UZ+Z9pvW+G3YR3h/p5
YgtRGbN9iI9IPK3ES8WxRMwB9u9Bjg1SVsdq2iYXojYM31TdfFp4w0p7hJZIwpBS
5RJwCb/vQ5MNEhM+f8KurM8ZoOjUtTljx5EC2zTdncsxE2Uy/0KMFjezOZLb2CR5
GIm0Fs11hI+fVOjLI60D/3WxDOK4ip3Bt7BUv4yKaRC+b5pArO1fwtlVQ+51eSMk
cL9Y/B4qbpVA8OW2ZV1uguRgfX5IQQ2T5TwRzaqbMlnxqyNz+5rrgbnz1BD/Bnvr
/wWEdxlVX02gB9Ur+tArvY0z5gH4j2Ij8SXieyQa/Pt0bQpTi0RshUuN5pvfyNBU
i90gxd7XVPImxTfFOPBOubj5N7xHBunMS9T8os5rr6qzAfyDIxrZ4JsSUsOlIYzE
qbqauD3MhfzdKfTfv6sSTPU+Brz5KB/Tv2RZeTf/ZWdQf7ev2wWu63Mm/lfCoVB2
qpnibbvSbFUqgQaJMiMYRVmzSJdAmoO5K5g2xjnjV8pfEQ/FUdsAHXnYvYorLPln
kLjODZwNzGQ3pS8FD//B4CtWE/aiTxkbYuM4ja/TgGmfaeOF35szlR/FNt8AqQ86
7cK0ddKSttkcw8XdNJKEDHQ31s5xo65F7ANRFVAuDmIkTunatCZnSDfpFKTHeXvi
gABXZf0rsW2FkCrBnzx/uxVDuxeoNjc6ztCLDLwDJ0BSQ6VRyY/wUjks2PNQCWKq
Dskrcwm3+28yDfur5aRkDoaCHzczKehQqHC5iE0Go413ubtjTfReXZH4rcHSrfWt
2Gg34bkB+fRcZYB2NyjE5SnnfqclqZpQaNGQOBiaYxnK1Cjw2kE3o9RwhrlqAcWd
OAJSdFgsBv2NahN+U0aSHhkegwmuw9HLwfA5Vhc81hjl98ci+PCWg2GCeT37jgGb
puA5D1nSxVjmJspjWg6Dn9x1BTOoRom8m3Yg8e/PRVRxjkreZag1UlELvsabWk7g
KpVcpGm0cwi2actx7K6D1Opi3dkUCOjhLb6R8zwNOXX6P9B3blNrp1IT4CQUgR6G
5hWi1vP5nAmHc1smxQfwhL6OCsMAL4xYROe/ulfzxb14TZd2I3X3sIaGu0+K2ea6
ndf8ESz779z5Dx+BEdSP7DhYee9D0QixARC05IenMRpag9EC5qZtW3t5eI3ug13g
XzNoMb1V3mY8pIfkQHM8kvqwhIWTa7jgUSqmo25ZabjzyTVF2jF5mTiyWzMQMnGI
7x3z0nNqHzFCK3RNk2bpRRudqMheW8+sysozHh8x51jkd6TnawHU83T3GSslC+0A
RBdREz8sybgji8khfIVea9aZbEu3Jyn93t3fvr3pHeNcjLdP/Bbk1JbTQnePJFsl
2K+wCzzqgrYaMpdK13jCYSpxLSvCVnJYPOklsp/GK1R4JLxJzmv2/C6k16tSrzYX
6XXCnuXvTUCpfo4VRSVtxtprWAiUP2BSKvVUOh1UQd7kRnCxxBEDXXcgUsOBCEg1
kEjP7zUKc1PzmfpkOx9ohFyjptzLiU8NtMNOrBnMq6iazoc8RaGj9KhrHeG+y30i
LLqMQLfMljNwQ+7gtuOj8UOD/NQ2n8U/VCD0GFLBEZy/Bcjj/8Rc54B3PEmKF6WG
JSJUvr/4oOAk9byLwvtV1EJMJxeWoi+8q9Txf7+jRET9IbiIfvHmwx+KdtOQI8OK
s4DYYqtx8mbXDAA8rwtX2Mqj5M9cxBb7xhkXNv4AJPe6LRe2fSRv1pWJ/N5zx4vW
g8OSUkEOwMfj5qsJ90+O1MAJlhdnJmLEvsDO/sZ93SC3idnI2TUXbtICyAbif1oX
nsnsKa7cFJm7RJ6JSSyCScws7RdFwXBifFYTGAmV6H4rAtptcnOfUp9CJtcIGPW+
/kC/95N0q9zo6MmxHPjtkIJsmqbjcUSC6RRYi1UCyPO89TWKN2Gh8XytIw3jfSSX
Eci7DXd/3tV7iWUN2FC+qahpzc8aeqCI/yV0nVrTDdEDq28Ah6Aa5Wje9RoLDgv9
cfZZrq7VhvEC6jh/c8RDw5GaJ7486qkkZj6WAxfJWPDv9gPHfDt+YLKbmq6fufGC
K3iloB5y1lU9HTOKrSqvRmTFOJJ2LUO+7hX9P2IUMZfOsoWhdJt87JUguzbHKWvN
fgDEQvosyD2ZHSpPaR5BVRgbwEbDTi4FG7He2tTUVKpNggRlP+GNMqrmvVpOUW1E
HU3N1HkJbyHK8wA45fexLcjEv5y8pPY3p2sppDghPKJXsEi0w86U8F9HebZ5AS7l
wFyUOTPRW/zTZn6gCP/8IBrEzu3dz07AqmgGt4HIzJGIqKp0ZOelQH1XDLS5OUed
rksNXS0oGgLReiPOkKcDAMQy2v3kF5CwvzpcAtZVPO4iBL+4lOyC/JaYuqplNq72
ay60d14Z67u+AFkpM7V7BGjEQYN7mDBUZqQplWCFzhnfwfbw4C/zQ3EklYZDMie3
XDcAa/FlNdBQfnb3zlVynKB7v22xJefkUmeaHz2QbfiQdfA/zY/nVFNirk5ULuSE
1ooBMr/7edD4jxzhFJXgrRAVS7uZ39IygG8o4JeBRFJU98ZdZUH4AasMbymeBkDN
C5rvxf2bdofnUau4fX9GJwU86PubeC5RtY+6BQOGnkKqPuo06moSYoxtMY7Iwvxn
xqUs+4Fo8KegO+3P1CnGy73EZRWrxKtt3nm+lk+qa7ncwR8U5DgpwewasUMv3DBs
s4+uZ+oFH+FVHJi6x6pTZzEwZMjfpvHRinlHWwVGtGrQ/S4U6m1/8pNvVRLLFneG
av1cHMxfwEDOsf9OyyKnR3pIYCxJgTbnUj7S+FiGqj4idk39fzayzFimQZ0PAApg
v5hOPSqGYsB5s/UJm2hcqZG3MzABPRvm/tUFTKYPg5j1AUzB4NpUw7iyWZ8yvj/s
vJWBw/A75VjOt6ZmuokKUwrQLV0vtSZygNBAnMvDKMDDhiX8XAskws4u0ha8NN3y
WY6vsfYyZ0XxuyxI6QZk/3vXSfGuixbGdlBlAojYkfv6K2La5PssN6yKzitBG+zI
hjsCwt6EId354XaCfmnl663heBEXznafEvB+ckh71ADburtdE1wCqo3a5pyJiZ5O
WZQUbVA5PkMjF3jr4gkLrtcHs8fFUJWSGU+iLLI/nT2PAEKenUMZkW9YEuVBrqK+
2JvyDSEK2YkJmD7a8pm/f1QWkEhWxf55Ajmo5WLJh5kMQqk+FsbmWlU4cXiVjQWI
PC/PPME4gR/aOYJYN4wtx76TDzWaP1VZXI6lGplrj9i4Y9yC8OkiYqSgJhfR4WXR
iUMeN36C6NJOsn5IC606qwtdlsYpBvYhIz/zyJenJmN/VqFGO1Xpc0aLGGuN3nsh
wuH86M+tU9VZI6ryjBoIJ7yDOZpVhk4Mmwo8OS/D2VaaMkbqAzVRrM9ayh1Y7tZA
jvM/AW5XrGeTzu9yba5R5HuCU6qIP1XAlO5oRO5MrwpGtx4mIPHihXsgMBdHtjES
YnoHJD+AiK0qkLkaNvmJj4wkCMnYzul7BW23Z8/c97YGVa8vHasUCBQC1HSmnRVn
LqUi9CagmlRQICfNs+ZmUTHCFO9eGVX/9u6ANLJ5X8pGeHqXmBgVF2UFqSmVwp84
yjWcw6sKvYmzxt8dED1fLSNrZzEgCsCo/JQ5G+FTVE6mLKlbRILj4KuqqkobEQrO
TIjiVNAi6zgEMNmzfBg7kFQt0P7/beo56/wQuCoRxtd89uT6x0bx9zjcltf1xDfJ
etXQSL+N8VFoVhTVfHMzEOmXpnc9uTx1Y9pyB2btFFglvlCpknI1ZGdeh+vliRC4
V0LkPi3nRk/IZQNYwERMWd5nsWNjlguG+4QYPOzW2ILFRb9pyf5fh78SBKIiuxuR
8fubEr08hL98MP6qGQoyTz+2frf/IR45CttqpUu46V39VYdPxZaG0D/opkI60NXr
+DSfEqdVFl7KAefovCF6ij1oaTqFZMlQYDCbp914wflR8dgvw5eIFmwwxfGTZLkz
T8oYR2Qfg7em6JUVMuUYwqWQqLp4lXvToLUJXnNpFnSVxUo8j8jyJal96ncYEfmf
Gjzydz49e3OWNiEGcR4vTduIIhjh5wWPNBS1G318OAbYdrn31MeKq3utgEnSqpBo
K3wldq4sBr7REksZcH9Y7lnQTYEDiXKJeqXW0+/FGNRGt3ThmjvxB+9eVYq6MZi0
GuIW5LvGxTk1jcJjN6G7w7zbgGgmhx6f1SZswMK8U1VGZQNn24RcX7gJDb9AQ/+y
xHLle5rpNoIo68UeVeJzfvTT6+I/1QkH5VNE/zwVcogkwcRTQMVxz1nJ36QkgwzW
1IZdeNMYLagr8X9TSLZkvTrGBLTdy4qRwtqM8iZ0vnqa4JAxxLs0/OiksKm5DtUw
x5HBNrBcil45VSeLDo1/v95NrhD511NuiX5ewIyXxad4sB61EBNfSaSuItrbBWCo
92qrc/w1LihawTNeISD0SWWRbPP2pcmLt/20WDI0Dbx+HaPEQMpZQc0lnnlaVoi4
MDWIYW4XLKbxhllLS6cMNuVcHj4Gaa13k4M+mCbEK2MGL242BTTqsxYopKpfSRtq
E/muDvESJZHifK0bJ5pxipts0sobU0zrMJCADI5ev34yiExKTzS7Ot5CMODpFru7
X+/p0rFBZTMxBr2i7YcCIuxI6F5RxHCCDZkv7WdvF+4ZXwOn0gb8z9UvKePtBLbE
l5XH+CG2rPRp2JdzCpNZUEdtft+3lsE5fVZJfKdb1cimBpYgDZxSUle3OQp9Avcm
7lpxblHmL2uzcvZUGn18czJKdBGKFy2AmTNk/A7cMP/oZY1JoDxXSFBk9KXybmMT
GwqpeswVUwJEH0KQP0JU83lJcUXd1SfGLRDQ8hHZiffepJCfASWow+n1Gn+0CEgn
x2fbxKJ+B4A4Qg8hDeVbCRH9lz6atde3s3POHojr2VUjPK72WoXhg8epV514D+gR
J363IesVyfPbEpR3M7W+siSBu6ogERLd6B+PiYRunR7jMpYA4y26LzM5Hm+tXgJQ
B+cMsfL3NFCdYkByrd6qtwtNLSdo2O/d9gFiJ9rJVIwIH7284oJs2m9d3KzXK7kw
ez3jdY9FKCn6ZkEC2nSqPz6tH8HzVRyPcX4VJk9MU/45ClGiEY9S8X4ISr/CwDPZ
NpzO8NMEM0clYyuVRJuHMBmg90+Zd2w2svOjQmp9IVuN92TA6ENzO4j60hthc8FH
YFQi64OF5KRC/GXKfs3hKYJ724Yb4kB/7KtZQn0L4OzWIL40QhiMY1ZOhkgf38NO
hRFml+ltBe29CrUor4XxVEwMLsVWLuABjHYdLzhsLkUd49MkgJQfDWyYj07yD2mm
eFMeIANk99LCGxmdzg/LgGxgg2WIDIkykGAzVm4ge/cc9qne5MMPjFXr7K0nlc6J
LCtlvUeek/r1Xp5KLhr8et4orowUVk9QyLVaPvWZVNB/U6mn/XGapqW5ZP9Ne4QR
x6HAVqqlX1itb/OUgVhbX2VG8W+3fpePyj4aBsZJbyYzc7mi6satWUTrI5juAunm
YHp/l5H0yBEl7zvTnMve+hs5RjJKfK7Hxd7Xq/2/Vh3EkdQridX2DzE3L4K70EP+
QKJyUuwZFOn0bdI9ZgUFhwhNS+S6mzmxFfnbmWLtr3+ddr2mpJMforh0EDv/BhTl
TJ0xm+OT64O3mBBGNNnFcv5eB5LyJT67tQpl2OKbCzXlyTK0MYlRad3lb0SUkATm
LK4sUD2MTajKjcfsaVCplZ6Y0qzJns7fxL9khkqpdZrxMghRTJniQ5e8Sr1uo28n
ud3fJiPclVf/WW9yb39eQoxazFYlH+FLHEBkMQIg+0EaOALWNiC/DkeNfmXHAhEE
KCghUVu5IuxWeHwJI8kZMucRS12mSDgeiJ4S1y6GvzSEsYcFBdvPzpkN+NBaoABs
tFrnuKqav1ls7h4nK8wI8X3cr97yXx+X0I2g10ylQ4Py5mvuyY47kKZqIFDPMMR2
csCSXCAkAMum/zHiVOQqM3U/OzkP5I5lpD+SnAStMMB+7zvvS9+jgoC6fPRIRTl7
e0/CMU8STqJnoZVkzLPXZqoIpeM8mB+bmijOGKqWoeHr7F2jI7fmTJaAaYpQ3DjL
Kxq1GZcpcrqsVVdfxnn0RKQ8Wes5vI/lBuoisdV9zRE6TkI0XWJEB1IXOrmZvATU
vzTchFXDA4R7W5lhxo//smdiPIJBnO20FgNOGtnj4vparwH6svsQVpGmGt4FW8Mq
s28YwquwOLcN6VgDadnMXXRxYbYP4FQz6gjGl9IwmF2ZefX6MwPabVLim9DgmRov
vBshiQoXrn1InCK2iWnPVSjSGUqE8+qKLLxKBL7rgPrDPm77EDs00oP79ip4/48u
8h/rji7VSiud/3Ip9rVUeNdYMWiCZhuuQ9r0arY0SiYCo+T52KtUdajxQLnQ1Fha
vhVWu8MhI9sHQfSGrkpB5SQX9meppTxDSWqEWzVwJK0ai71GRhoTWbaz7UjezTIm
iWh0bFi46hXO15fZrD3LekXgRCbTAfeTja4blYzzC0mASJKAYztB5LmP4B0aaKMT
zyolHbw/e7Mja+EmhiUqB4K4PnIdiyf5dQKzubnMhfed4t6bB0ycWqDzzdBzt2zv
OfCiQGwlo5hYCTMma96+RcSmwvxUvCj3YzAZT9ivGRc/pbM7ZHsNyL/L9vzQovN0
yvhcZaKn5htQSUzxBI7o/yZTQYPgcuaQaBGva6egN+fo7tN2R5jCG6MF1B9JlH+i
Q6qmN3fqTeUw1xtb0I8oXMup+AAUnotoJfWK2YysFVF3/knpqfwAJBW52CgNGvJ8
yJuDEFvsciPbd8rwFwECkNwcav1kCbeOmJhJfnPV4Bo5SQiCiN3szL+mcW61G/ee
Q+VxwESTrRl9QsM+fDnOHrAk7otE1+nA7cYXpeH9GY3hSGf/H7JEQpRcg3Cgzzrr
5NhjQsmFWiXRmtLxBLRntoNgy2FuztZN7T5Yp21GJ+ldUQEBUiQQZ4eRMAuNaL5o
fFC/b0mZSxADfEolxAAKrtknmHt1DvWGglLSrXREVV99DLA/kBzYHTYBCypD5Tqt
m72x63+bEIdIDLl/Ml/Bt5Sc7W481UpoIV7w8s/PA5+9s+FkvZ9Q4SoATwNDyvep
ynN8V+v3jSNWVT7micnZmxYDXK+md/9MrSvidC3JjbhQh2HzY75c0wfZMX8cz7UX
xY8NGcnTz2WrRJc9FMArNuOrDh6KgZOB7H1DE6gkTel1XW/ux+FZkAd47E/+DlBM
e3vEt5u6o310jtEST5/RblfGRCPNJSnPx3TQ1TIMHLjG9fAgpcuyLM1xSyLS4WA6
Ed8kFL9oiF2BKr43G6jhC+dei7FZzEHgRrh4aZW/48c1rQD7m0ipqhcN4yrdJfVi
1GvHCmm2FrjqVUYTiPXQSzuWD1uc/RaUPSKx1daCBuJbP5DhrvC/jNDedWj3Khli
F/g2ERzp07EYoiWe/z8SkJ7di+2Qxi9CuD4ev69Y1K/Ofo2YFOoO+HT0BBuwRsep
DIv0cGqvZvnAqCiEj0dczHoenlSQaGMx01eXknREunIifP7aJ/VP4IRM9pxYgWL+
3sjk/a5qQg9+xItALI0zu2vrxpzZyJhl9o4iJOrUqxukwwmmfM+SV2VJ24p61d4+
36EMMNm9AsgWit28OrfRIwCf17y9Fe2Eq+aP+5ApF5Zk28gNPprSGGtSWACG39z3
pfk9dsFcwIU8i+Gl7GnuMKfZBcbt071QV4pGgv+8OuPSR1NtqKJfyLWj4705ielU
hUOscqBnnJalOSmzdWrunR4LMMtD1HUOdN3EnCN6ZgIqIuiSyr7a7HT9s5P7UZDX
C2hcoky64kESeVCFRC+n3ThEs2nYJIQk6CBcWxsMCyGHO7CydE5lN2+SIyHrKVNo
1NKOLgsTS2cne91Zcp/ZYYyTjR7toWefsbk9PAFF/74xZ3fmgvnDjHS5eH9byCms
B+WzCyViRe3QdQjfmlzzmdMbZ3r/AzT45GopXDzpvjaRcqZYtt8eiTmqyt9lw82w
62MpTBppOdZrmzeeI81NmTr4ji+ZOcx+6JQN53qz2k9gzEg7EoMSneOJh4bTNRRF
A+a0EO5QMdbyjaMkTStHKqc0GheXfFO5OR2nc5QM9p/GcnWmowOc1YI0DbrMW/vf
jx65P6mq0GRxgns1yz6tAdaEbxUEa4sF/QfqVPMQs34KWelJw+2Qc3jmu30I/RJo
kxM2g8wlWoqH/bxlwsho3d4jNtshQ//xzL2+F5IlIlFv/UXwVLjzXa+nkRIi/3H2
/gC62jH6KydqrPVS+LZw0GOgn0uYg7bOlhlAGUiK+fp8/pebcKUvZ1qIm7gMxvz5
ow5SMEWBqG5wUQYamfUJNtOgeIwufZyPMi3ZI6DkBFe5W5vxqeBC8cO7kF5K2/9u
IpSlZkGwOv3JbgXJCxJat/h4BY7WlWpMjZp40te0d4N3H+fp/KQnV9fYwXOWLl66
o3dWXAu0KIL2HgD0wUYTGs2PRP4NSDMKR1cDYSR/P9z5UltkH22uXaB5orjxvESj
D65RLmi9lR20ORvqjXM5IDfesgwtr5JTT+1vmzkH1odNNJG2XSxhAGIzhsN+XA9Z
9ZYxF7P0U8xG2Hn6iKwnaff3C46zJ6GTAWAnu82sZ63OCm2RB+Tk39WO7Wl9gtoM
ikCScDbNZJM36RIehhm9HnTJRR9OhsLs1PIzaH+hrBijA5ArPpLZ7LHd7ne2j2/z
njdDAjQt0OBOyyonr3U+4RrIujXOR3mvwKyW3KeWMPiAGA8M0njIfce74thDXPnA
VRQsV1vaWgMVDuD33nwUxcGWJZ7DhnvF2dxLYfumh028mktRY/+MRTWLMZMoQ9Qq
8T6nESntjSCjEkFH0Eud8RrwONBtNDygaYoavLaTskE+Z681dNd5ZeqzysfTNFum
ljgmvtLeqi+b4lAMeg4wWEU/TgsJaDVENruqpHcZu2ULklhbT2YcLQ8SRrMYU+/j
hhndfvK9C2LfMnhz8Z05mSj1PAaCf6rNdxpr9x0AseecYC7Ek059Qbn7NvqtjJg7
C7ROnZ4Qw7GrFZ880Tm8t9m25csRZceJtJ6qkjWS21WOyXH7gJKMXohNu1g1T2oN
pixEUb93gt1/Oc8GZKSegH+70gkVCOEVO6T+I2Gy/axMUZ/MMVgpkqIHO8K2Mb8Y
tksgBivSPNnnPROOHCEmcMPEhPMRVzt+wZwEHyNahjGPYV0L++/RsfimMCRCIKYh
T5tn03POo8UjuDJA9A5alH0G+4Lt4FtH2xVHLgCB7VKwEDyifl4BhW30HztX8tzL
4xrkA7FfzaqpXJ96vvp9wxzDvkLO1/omqi5A4WYeY+zBNeAdt6oTFBJbAitDehre
wkuBasqD9c9/40jWfZ9C7xgout37+SWYVPTHldbbeMumxVfp2w+G0Rg9AZ3tEj4M
kNJUsXTPcL5z4WDmciEvGmAIJJfqiyjYLez5xfVLAGLzklQ164SE8bJ0BhVzXpqb
jlyNB2wMRQSltXiZludP2R4miQwG/qi7Xmilc9XjlNsYXevHucEfrmm9MPidXvA+
UPq0ILWAQOrMBHF1YlUc2W+Agr+Ilc1wQEd8IeABaUjV5+H18ToxCVokI3A8oMT4
QRNdq9R5wvJg06uPQ5bYkHkQjc1RzgdrjXgV0BB2ofGdwQuajuuNwMZijKE8AtB1
EB1zpCpVEY3vnYtxz1myLUhOMiu1SGanILZHO18IFGwhTirLDGmqPIoLPXNmHHq5
vFmS9HNZxC+2ZI15Ja9epX0SeQC3jn7JMYffFefoEQeqGFoJ6goIQc0QAeVTt5F0
GuFVEIM+IIFTMQboroxD2LaVpp+0/QKwvDa9eQpfxOA7V5shy3+Ct+smFJDYVgta
BpYWDDVWOeVLoU7CdsR1Of5PrJw+4PvBYogKbbT6jroTutP4V1nOncMKn6+QRbMG
eaIzSJsUjChLtVrO40W/7+R1VT8GKDnfyp/fHzgqssmbhYcNDhOSqEH8Ha7xvL7W
KMnOsbZP7fhQNV9i3jFGPIkPiY3vxJo/tHWnd0nvfCNAFp8Dxi9BMg0hf5whqY4J
zhJpdTCf8qTHgdCyoEhNeP8vdjsdnQCJq2nyRWmTz2j0zdGC1MKM+yM43JkyOR72
BdXVyteYXu9I1wqVBsZfabhmiBg+c9GzQrUUWndX68ilMmTIJ0u+YqptwprTCQUv
/vaKRCYe56EUmr45oq979GBvRWGzeb3iKkNOT7bgoO0sZCpgXQQx99RCVePUg0nw
2GXuO4g7btT7nHnGLdkCDsaAcG1+fHQshVN7l3YiaHcKtLhnMf8njm0l/zjtHC7O
OWMBoRMdGzy29BLOAr3KbPYZomI3h9aWD1NSmtJN8r+QmLzuojXvC6RlmExJrmZC
Xzu+5RESA9JU3UtwhWjXxNrCQQdlmxFgkNV4ouvll42fqqR9CjRikFE5w+/rBRtU
Bt91JQVmuAxo+H8sRsX/D+0+XC08koLpzn/ikFcfXuNvMT0+pwk4TfgGJwRxh6ON
pwNVEgHFJtgOQcO2OrL2WGnDQ2068B6Or3JAu4450IbR9lQM+jbJIPHpBZTYZa8z
rMPicFLsXYN1Rf0wv9baXht+jVL1d2pjjkBwcL/AunkK0oFNO9xkBL7QLmuNK/3A
DiRxvSO4hUQ1/FkvITfIW8/Cvqxlq4x+An8Teajuev26QwvKk1Y+yeUCWcB83SEe
V2Xg0YBTcht9t/jZvNfzmxtPNJd+iuDKa0QnMNEqTFvOhmFezdrkqjFme4jVp1dk
c5nr5bIUygTGeDck671rUkFzdnE1T62LElMwAJzNKVjisivVzossb4NqKuk3sgRX
xQPUYwf7cpi3YbUCDFhiIac+pP3EVKfD9ttFRV9mKt0k2xhG/MTe7mXYCamwDAKT
pv4a4ufC1l6ykgJv0Pdfq7wtiC2atLDCJfCVnSRM5QdmTb6XGrVvwXbE0YpkJ2tV
VUHt946pEmHETDum3t4jAFopI1StX1TK2XoDakKDcZ8GXd4K1caNbYX4s4074zV9
U9jFt0Bime76VoGrOtGF5WE7MQzr/D87RagmV5GE9DQk9013fofotTgWNqFqWeiT
oaYfOMuYYbmoEcLc7yZPT8jRS3MQKRGPaZEQDDWtpwDuvvqP/x1aSSYUVeVEBnRU
FP74ZoUAD7E52AGHGd1Kb6hDdw849jA4s47AOdZWwJ5nZfTETPOyx75K05w+yRCH
ThDGV4PiIECSGrw7zLTkw503ipsrKOTV5dS8Yn3ho4QVor7h7Us+SHaKNdIoz3hh
nC7ppf7Rpz3PQfhSKlSWyly5r7bllqLB9MIpDQYkU2Tb7rP37bMZgYM2rUesFRSv
u1mOmZxHeNni6AVOpEgARPRrCXDZTsSMkmkgGwBdncta45vWH8gTLb9rZbRqzhIc
5QsCpV9CzO/jOgpcTP/EAq8hKdER1nK09UkiOl+XlJA9hD4AO2LEeHAuZG+q3Iip
2tUpcJ2d2wNyXf+iYbpelDqfviDWih8kOC0yyjvmk8Di5dFE5ff1Fg9di1Lw0RHK
FuoBFB2qXEdO2B9pDwrX8pA73d9Kureh4vVzBbOPGYfM3YhEMPL8DdfwJxSuAtMq
8adbqc+56Lp7HmVli2DwgJNpm4XKOJj07N0juZyUif6Ght9Yww2q0i6dOio11r/o
nsC735qNOq5HXsgufiyXzHgxFiukKEXhMrBqDisYniAq7a8J8JpTf1onl1cejJC1
nI9zkqJAMg7y1eiMBYf0/MqEB11c8eNSZNsRuDu/V96kbInz38M71GmssdOpuaVD
Aev1adcPQRuRQQnEhpcVuhbasS0xPnV/ObkOQd6Y1XX3IM3lYHTp/MgYCBd3mqwz
+XAisIVtAJ9VAIu/qRm+n+xzf3QdCkgv0LxKd6j6Tc0ui8ZSY8oE7EKxNnMYowPx
C+SbrI0+biUxstX+vyRJsjhGf8/ogsVsKyf6r9BmaNxp01mii7YyEx5G12uX7JL/
sSC1v/Do3qNCzfC4/tYJ8O9p3YJXmy/vv8HZeWNk15xCKBsdDEAE38RXB/Q1woe+
pdIuoVrRWr2oAJ6P+Orhfa7RyLaHflNhQfav6yNr+64YWp63H2ux/paJq+J6jl3D
vwFlGaE6AlIh9LgV2DT3S3oeT5Pxju6iQpSGNMqWHum7KPsmG5ynAwIXuDjroQU3
EvQNNAtkpu1muFNjSOM3Shf7eprNEr2j/oa1ex1mdZN/3m/79YHJH8Kd9dESr6BF
z9QFnZTPvg59lNx9Fq2yQ3GUQBFCRc6qyIWe0rveZqb3Ca4DzrC45xpSYSigQPjj
Fmmqf9kEGovnC7V78VGrYc/QqgtJDmLAMoi7ub4NZg9VoMqe08oSOwxWM871q/1B
IhBl2dUeo5rLl8C5OYJXIk9BZBC3vWYn5an4Lfd2F4qBFGf3YdNSunhCN5vRBQ1F
dH5lrQkF7qUejwP7OosLKpy6BVtfOOewgq4koiL2gRlDkx7sT8jDhPzXQae0+Lmu
oAuKREAMGrxBGMN8R4/3BR+s0F81jNL7S76q5BaBooMxdPV0AZt8FMmwAcRsokj0
e4OBaD7E0ghNBVH5nygJT1AvyPSUa+J0g6NIk2PlBRusQrPBshhy4AsZDKceGZuz
VJKVKJ9XtRlyhWpfcJY40OucIivrmMD5Y3b28HyyYfVfvxo9Zm07GMc6WnF7uqo2
tQxee7vFiDfGYdGfFUOSb934neBTsHp1R+y6dajYcFSEaePbqxyq69QHredFohNX
IicRByLnOaIFYlNJd2FS86Mmi25t9rDyKHoRU4sijeLCgF6LuMAp9VkXl5ue3D1D
h38B2vydAg/B7ytRt38KZM1fdY5IZJwGi5IaKAu6wkPTjrJHbR9WhMzqZHzF/NJO
intTJuM/GxR9sxJzf43n9gZvTSaSugXdLMTwePgoAY0A6malAAyF3aaKlDuvGHUe
+C9k8kVTrWX44A53Ha/o9Vfobmet7wA9Sur8zVzJKVh/UJieIT1Y4HYR3U53DID3
MWNKGnBex65dILQHFBtiUbwIIxgYty5xTKioOcB0ftzD5NWNkMAcjrXgE5O7+pxF
9ARIWXUGdgWRq/dHK3OeuVOKEqVpwwlr9eSc9b2VrCcCwXK6C89xdU2sUZn42oRW
yGwAe10OHRNJJxhPVcCSvzPWwI2MJRpJQ8HQ5w9bK8x/A/woQkUp6ilI49DCzf/g
8sPOOb+cWLr77Zzn/qGlYRDv5mrOpKhtT8vO6FsLz3fYwn28fE1Ihwn1bh6bmFCS
pk9z2W9V0o+Yfv9Gzx8mcgHLcF8IyQvwoTpB6uf/FbR91FlMJK3ZCI8Igzs3gP69
DTvO1sKogelV7gWwCIjbNastL6WIU5G0MWaELEXC7YWZzLgI73L/aIQAcDL48RAy
w0XPkXuU+frrY6WL3m9V4bTbrwWDCxkX1ZnIoUEjACIbrMQW5Ji34QfR44m+1ZOd
T4UbUDadj0Rdk7zPmOQxg+o4syP/OSZ10NNTV5WgnOM1i/hk+ZDLa1Uh2oyMWrLa
NR0te7kPkSHFrzRXWnciNl6tlKzNx6RzFeqXzFPKh1DB6IwEtLnstWKw2KBa2d2y
e4LtUGWpWZdXY36HfUWwAkXWGhrvz+aEV11BWCqKoQdf5wwl5iVVIuK6VC8BYGYV
Z8eAQcs1vtblvEbbN17mKioZIaJ9U1BWebs6d8zBnQY30T1eicddu+zqBs185v3/
7PbolAoB3eqcxONXQv9cTNw2u5a+YhCL4Fienso8zTgWvGzabjkppdzbwM5RabC6
dJTbIO8QUxpEgd7MKgQVj4CBx1Y+jLx8niVnZaLM2UQuQTiw7bRpuUW4rjUP/ejJ
klR4Le9QeBAmDLrFK8Z+sCtBlH3bBleT87nbLgZEaru+c23YciFhEOJOBgCSlP6i
RQ6ip2f3pP6dn4OlX/hwe0p2ONqoCIkqe3nBWWC90nQxewJuB9NTLTLyC0PI/tQk
sLSZjPuJk/Yz3eEb+hQ5ss+gp0nwZqm8SNGtaS/yHIPAXqDVidxyivK7BDOPfLvB
xUp7zPepNclrpRIOF+DIzyO4WxdNPNpKgNnQvWSpW22Pw0JySpOidO+gJrJCPjfx
rozH2SN8Zqc1n+ItBg9lIHvihzmA/GNxHpn/4VsSjULD5IFQlk23xdOo3xSWitNz
iC+xJV+ZImBuQfarjcVygE6XN8ojzLpuLKqqTcX1nJQi0c1FEgrrUdu7JxFBgYMm
REBKZ7//e/zVxsIBZSbSp+Tk4EmfNL0Gua1rny7rMKJfyQ3es1fkfF/j4le/u2XV
KSd7TVBMgr7qX80YvV/9bngXyuMOzgk2pDmqr7FNuAPncRiBapGNW0Isfi+yG9uG
mLyAAUHB+YLcbJ86ZyDVJaGjFQRmBuAmKzL71kDQFb5tsxNeNLG9zqKG3ymzwmJR
YXGiIYxFgJtzll7K41p++cTlMz+4iRlicF7FbrSOuW5fCnDebzcU+AUMAz2wKvkl
rZwP3t/NYVzdVdgOAu34eLkhRlfXp8mz3PwRb3GN2Kgm6rOvLOOqREVIFfmsmh8z
sut7iB2rreU4ePiVSVFSThteCEjafRGVSbb6ZTaJ9dguD4jhEiYYOHvQzJ/yu5pE
wezi61vGM/Hv0kVZG1Syyxbl3X7wXCawWIpFlcPF9Le3hNAiB0koFWiCvuckxt7z
7rD6cfMC8uSKJor4O09rBWtbCpVSXWqKlsJtB0dwzeBpNvrBuXkbeq9S6FnIsd1N
QVuuhU+Z5Ze/n4Zi9Ulk9YqD1On9Y7kpEeqjWPFb6hiWg9OSuC9r5mKLqEV/cNh/
bIUAVyRuVJrFzu+qpBUxm7lLGbOM7NuWnncpksrb+nG3eNo2VeaA8yLZfDrLHI0e
kTmcRT26XQsssnQukmXbfpf4Q4ttT4QikncD1mbKBc3DI+ZphtxhUCAlvo3Bbagi
DQfLm9VUGqPsamB7sb0My9+VipHt0qlZ3i0xv5rD6OCleh98qEFK9u5S2GeBg4Zl
47qC5hivH46G0a8S93LCj9EAhuL0YRig3KsR/B9KzyauSx5Kd8zt2zsaLl+RzEAG
8PW0tIudvFBgHnlfsfr5Fpaw+3imEzmYKbenflQLsf1ha31Mf/0kNELneW9TYUDo
0ELic4f6ggPSJ9iECMp13bPqgZr7YnEVjNQHfcEgmqNF5aXh8REW6nJkGZAA1HXa
XGdwAfdWlVtb9syFSVepjVE0KI7exWa+rsxIrGgUKWIU6PlopnGkcybPGtcsjOb3
+UU5NTeNaM6JzLcMLIz4ieCSSB1GVPzBEcwPIUfaNay1RiaxNtSiHX6y89TIBFXh
0+wt/hBGJgsQSddSFpig+PBD+stvPfDwX+KMDI0SiA22bgjl4BovulY0NGeaXoS/
H6fbrkljj3HE9u6ux1tInL48fcfJzQ2ddHs0SyMCIX4o/miClzEbnrgoygkqC7g2
6klrICjBhiEFBn7aWyWb6R6gFFiqVb0GTaTQ3vMm+mjEbxZooB9hzI6d/Qfw1m0M
vkylif/jKqu208+KmuoygBnLQggNQtIROdRW8S7XZgfDyL9RI/Lrv6K7JRPWthKg
H+l/lh2nRezgbif/hM6wk9enOzj4gHVPNG8QVuLIkLAZ8LpWKlhXRWvQhmTzJ+Kz
pv7Jq1RRciJTDZXeUEoTxftKEUQgaKz57FlgeZKnLIfmd0f1epoHbJhv3hyLzrzB
tw5ENeGYdI2MVamM+WQU6bPlx1RJt0Dl0Y57b0qiBcA9rbZySwGJ0bAVa6C+sEPR
lgvItbF0MXuzGbBjVM1D9orh0rsPA49Zk/BJyg+iR6soi0xVYdEPC6DJX9laKvzJ
n+Pv7Ib9qtZ7gM0SYc7DIUaKfyCFUU1ljnPDyitHcvj4sxBgBj/w7faL/ToXxSRo
tGI7KzPbVoueihfv+HOdIWjGS2sidICzF8fV8WCAZkINtdDmmGpNS9gX25+PVTTv
Rro5jRkjfZHQ7l8ZyFPx+sWv3hPOGYny/aLPku64POUvIYkAhW985Ch0cPY8yXCv
vG3iTlw3XFdOgJ4vwwticvX95sMVv6VUz5HEt94lWWM9KvTOxvILWavvtk6LbDqa
3Gxk488kal9WKjtBcd9B20fbhMpmI96E4oEX2d7FHtl+LHjrqAdAjRlfbw/0sgkA
V4Sn0208oEhsd4dHMpFpcFjqFw3oRX1FlHazJ1ZcSk7I+B8TO+EeYhg92VaFyWs9
PvM5HmxZmWAraJ976DNJyegKIJBmyPwiLTPJ46Z43fbcjxUaADyI7G1EuMv45NBN
nBlWc4HIy9fGuIaFkOnTILKrHIG9AO3U7olW6NrwdxZZW5DCfvaOD8MFDaenl792
vanXJY7QvIw/RcBO3uXPEPAwUHvoI2Xz8FfS3ChPVDcMS2vTqqu/GlZDPwcPRjQb
DVMuLrX4ARRlHxavS4l42bMwmPRoW7i4i7VsANnyyTrg4k1JjzPBV137Dcj3BHC5
Hgx9txeyqZ94kM3OQICgocAoDEV0xM+DUt8MH0E0AYyhw3yvE0MdyUg7APC88DTe
phXKZuYDr8e/r8s9PwlODkz503jDsLoneRaxpOxE1kl/A+42RbiMuMxE3vrcxMzY
h9gshvtQshGwet4iJukM3awyu+rSqFcEHEdV8gERpth5L8llfNEKSP7TQEdr2M38
8HVc8IKHWliFKR/4eD756EcGoM+EaU6ljWZHE/q8vUl6gFVXOMQs2lXazIlMKRIl
D0aeVr7+pB2i6xiDTKJfRNkctCdoKf4tATNzFMjlMFmRnXMHOoaI4YnTsJWBrsSf
1OJuDEDdgZLShHMYOz5LfugdLhIba1xazk2Kz3kx6p/9Eu79CkhlhUk9zUyBkxX4
Kr8O9besi4YsHCzzwmf4hhfM8ZdDwtc56lgGjjB0dB33DNvxwKoW7mnfkQKgTDYp
mzVvru9FHGTI/9vTn35iMt2DW1DZ9gRca3OToVZskZxB0rsdCpJUwc5m7IJt8/b8
Pw60RfTAKi4jt+frhoMuGGM2Y5PTyYXosUIzDbQXEqnhxE5v3PQkR6KqWi2FOj34
JxbNyElnmuHFFQOVdXUkU3LqRbe6knN5Iwy4uDtOhl2S+FEXq4E02RsjSo6ePqfr
ax68DaJYnjw51linjsrDu7a0s/kR/3i2+pLh5bxdXiYPUa+6tFFmNeMi8GZbIi2J
smv0E29Mz7J/7uKSi42p2P8MEiv/uPvsG25eCtpKQx8J8aeDOC4tdgsvlezXJGpG
JETUBnkbKM1So3kqm+/JPcqsjW1hlXVLVGHsJhxW/kmNtKmwgrJ+y97OniEq7nRR
HVGgt9C5XomVnF+OJhrFtSCPBSro42R5C3k0xqOdGywSKixfrSu73oQQNfQeV5Tj
XS9RGIi+O5naFo++H6OQj+CDSHxhC3b/1KLEC4Pu3i/vrHQF0OHDTVrRTRoe5Xcb
gFK3COifpoLeclkg1eIMZ5WKfemehyidGFOPtfBZ+V0534XoQXfNw2MeyqmQwlB+
M3l7uxHr+Kfzzn//q5rt+m9ESurrOcG2XINP+c8haXXqQCI0uFo1DP1XJ4TKD1Id
JyJ2avRb4htTvZjdZNUCwXLLVQ20+Oqb+6BL3ADmi4b9q8aVzXOhIncXSiLeex9T
IcGxntgZ4YWZxnZmkliksLzN1DExFi1BipTTy0GI7M12D0oJwfvzcbzRaKM+yrsj
OlVD4anbldiiA7SSr0hRshW71rucvIFAgbtIDUp0J29Mtn0fGYgnX5ZzuouHW3I4
67S5t7rJIO6aekaYfcRwsFzJ+kIk9AVkwClGbC/JvpzmS06Yky71WdBL7dOJqpJk
lmL4tRkI/+3FUgmhGzoEQCC4arbPi8uTKaW/7KDjocQXV/AlTYn2kCscC5K8L3TP
x92gVSdvFxWCGqSSpNyoGRbuv6TULiEqBRndqjt+Q6E/zIReN2/Eb9ICoIsoR4Yp
TeQfFvxyflgd53I+1Uf6SY45gKC+6rT9ezK0DcIIPykZmQzpYqea2K4kq74MSQkw
2a6EoxQldejQSyiAHC7FEkVu4OJHSGtrgKBZmuJWCoeKRI1triIt1k+t8Z9COr+L
c+TTz55tpT5g4ke3hpMfC4H8CEb/dZ+86fNCdIf1Awqu6YS6ySKIiJ5FsgojZNqz
l6uFhWZJWfaFZSjI+VoROHAqDYvQHyWoiJLq3+ID2tYOY+d2FoIUFNGKq50kKh9t
FvPfq3ltmUfgeC68dL6WK2nnXkHtxmfPsVdZSch3IW9aevGiTluIJcFMWM5/CZ2K
ta47x90Ra2k+Zfc9YaJ2nS1HRQlbr3xyCDD2Q1jYx311hvTfhWd+CXymFNnFfpuJ
z7q/tiClPD7YSVYovmQR9q6mZWQ3QUe3fNReHYjdUmCsPNSHhvzN8Xv7iPloX3cV
ToGmgoDVk/E5o0XIJaeVqGGSicQNKGPfwC8zzUDfZnLYdhyjuniUuvazymG/P00s
N+KdRM0sKqUVtTyK0tSsObWfdRygtjNft47HGjPK/bVI7WNrz8IkAHNHybcB/iMC
DOkWSYuP1ejifRkigDFPQqjs1asGyJ9BnjPbu+PpG2qUTx+4qIQBqxuyV72Gm2ch
JedPWRqjVSktf5LSG2+asb6JSUo6NeUfIRJ6JN3bKnP8bM7/GCgoo9106Z7uLwAd
+4xQKJFxCMGI+y33Ug7uxKqZDgNUIsaM/ElsNgQxJDgDoPoMBRYt8GNaYg+vvcKr
1GxRTfTOlHYDwGkTk9ilBzYOcybFCxL3nceBnB5KyCfcX1CJCb/fEOLS11mnxVQv
VNQ1TnyD6j/f4rmVD3RBmYF4ZC9JJe22IMrY97MuuGLWJodgPNmnLQbl8wpAYIEk
TMuK3oEI2Td2NyHT+uYYsZ5w7jButt5aXyL/a4jgm/YWdy2qi7Nsg0uy9YfWltiM
MyvMFbSxbKHPQ3PmhXCZ+ZPd8+q9F73yNgsQ7XRiDDyVjTGoYshH6Wy/AUGLwcvQ
tDMY8Pqhjj0tdWcOFqsMYxZpBB4Xkk/jhWLY49bSk7aZw11FpC+6GhFALr4a7tbR
aIneV6f9vrix+WL1i9QHOrr7TY3oQdKpxvCvVyhCDfJFtuqxOjiDHcVyOLXJNf8Y
2/2YNWTyGBLP3NbH+wtThympej1xIbwa4qa5SX9RQil6s9IKXeBsjrP5NZWyCgOz
Ic/b7KgwZUtV+e0kTuSPZyNjRtaLGUnv9tHTik5A1SlzsuMOvL0+oxUFa+duz3oU
boPXdMl4AQ9+BogzGgklRF3S10nq++DjoCaToNc3ei/y0rUn3tMyB4o0hfhuQCvY
j0s3LdDYCegu73zeAY82/orA64z/qHZzLRMlbnulvd/UejVEW8gcAY/wfh4apbPM
D+qhlpPiwaR7EczZ7CFGHWjrA2i+M2bFLl1c/EXBlWvkwMbgFnQwnstnZFr3rbTN
mv+FtmMJf1vLDHboTV0Pkb8c8b9vL7HhVho/O5qcXpqUG3XfCShNwM5jsGiumKK+
lX43Zn2BIdQYL2GOxchlMuJwtChJiqLNVM6IOuqXaXuaYpPGscH52adE6fR39D2Y
5w0XKc4b2zNxKIuvs/vCoPU3HOAE+pFKJuL0zF+FOrc49W1iUV7BbNJr41Zt73HN
MQdxOr7UVm0+vyATNLaSvSZi0n/GsSwTN0h/QIMkO9dUXZ3vBRep3Y1tDgSnKMHk
A1LCdqZEDo05aClnG9v20kR7DQ+TPD07YdWAcKBD8AEu6iC+ve0dMwCluV9SM+Az
4fDDiO9USSpF4LUtNRFzGtH6v8W/SKJx5JhSo6Rcf7ydL3y/0oSAkVX3GD1xokWL
AUmjKmwzfGBic98h7iZW7lYNKPmgKQyTxEsSpbgki0oHt7nRjONF79aQ/xgmXWOe
XmrpOhDT/hlDQ8lJ2zJxVKKr0/0XtUVEIW9uHl1zUBqz8BTkGFqMAdk1MQT5zdNI
jHvAU0cWw2ZPtjAUL4jEwKkgY2W38PP5FHJ4X/MZV34Wt4IfxtsQfh2wmFadyTaQ
do52Z2Dfgnd9WgNCULk2f7RVSV9KBf3x4r76mK49aTd59i+32pxppX/ehUM9e/EC
ICYuOpXRnUUbycx24KKgmNfmnThauAqi60b/U3ulHefCXN+1mmys9hl0SqDehjn1
IkcYbBnzB79Q1Wf/uDK/l5mrI1TDZFIi1mBaVFssjRxFFG/hkXNLiJGzdb5Aqt+X
jSjz0TVglr+upuPd3QjlMieYfmBmglALIGLQt3FCvePaI9n/W569asizkQub9QQZ
ZtCex9PhPlCz9ccIcsbqGcwbILJw66Lv2Y0sOGzmPljl4JtS/aItUgX036CRG0HN
5dVrvpKOKxGtfMOb8OlY6NtZcSiFyid+FjLPwBnYJ/phS+8Ak7hyANWacBpEVcKs
QUlKMhbD8zsO72fKhrQhdflk10KayQSdATPk96rDi7nOM6OOUAxc+cyXv9qd8csf
UOTO68RdK5W8OQfPy3CW37LipHEXR5tHTKVsh0nsXe1TURTVgiK32iQoj3Iq9BqH
XKyiSiCnNkxDoPcMMOJVEFMKn8HuCbfUIK0eL1FJlu/J5/7lHdK49ZXYXB8ZzHSK
jvCGMMcNA5fbMy/g8TUbZ5tmtrGfgITtGf3MD0wmNIqpzmxupoBMNuD+XqIhOs0x
4HZ/UebYMDw7HAoskA5M7EhwaslxMga8vAQInjuDltRH0X470xtC6tauqVHERE8O
VKiLkBuOAcs+hEW/ZozokXQEV85U8zNoHHVUcDnkJtfMN4Nf4Tw9cAkIckPO+WqW
R7H7W8R0tgS+atIjTsmduKHTfN4RmSJ//fQ0fqI8XMHfkdZG+ahdGwkQ8xDVy8na
7JWTEePK/YMAT5KvKQH7Jvkwbe8vTEQi/4UFb7xb1mXo/92zGzwEBOwP8XCASJ5e
inq8KKGNAeRv8e6/MKjni0AvJ8L/BkuNJDXrKn4b4QD+T4wAqXiBujOtLwIiW0+t
Rc2OJPpjQ9b8EIqF4Rq/MfX+kRIGX/DxsT58rfjdgDeqrAKaf2IOmnfxbQrPufyW
R1rumTPRAyMbjcHdIC9l81h44qysOrsmvnHuram38Eyu+yZBrR358fF3XAcLFg67
75+jVA7JVend5NrIwCNg7lqAXZPz5vauAaVG1CjHeTeYLnbq4v8v54+SrsOU08TA
lo+/EFy0hXwFLahApuPZjI+P7BioHeXn3n+pVvbQTL9TvTDSuqVye26JP1lcWWQk
0L0783Z2C/fA9Esi6D0PM6iaBMyrS1+ZNdj5p3iw0qm8c8HhppDo48y2g9VOxiiU
q+6jqIyUBJFW9q0vkpU1zJb2CKAzBTXrbau1y8BzfL1QB6FtL8Auh+qbp1c7yFYQ
5wAUsUnwnyrBFl/Iy/G0rA0TdlIDSs/aqLqQDVgccoN7Igi7iaaOi55QkOkwX9RX
Xqv+yju7Q5C0ke5Qb73fA4cwnj4PCnB18FMbpR5m+5Pq/QjnHCc7O1enKgW6dJfx
5wF4waW7HtfVTdLvQd6gakdKBZ09TiKP3QVb9iKmTPNLJlfFUYa8bpNEL5bUasHp
Vjg8AKR8tDCXpZFJniqBJmbgePQwu74f6SVRFs2bRXv+3rBZdI4siSa16GU155ty
0q2DFEBP1Gn6+AzM2URKYTf0ueJJhRPEqKdDLNfm9DjVMKP/uRhHWlAzuecAlTe/
COY5PtDsmOrl3Xa5Fj7wuEItrC1Ysy9Nx9pLDEvxAwcFhkqhzKMJGHqTsyRY38Ne
B5fHaxlU/SYAooKr+oiv5HlQKZoIndHsTJ9pLqsxNQ+uK8/S1hqz1WT7RVsrGmlh
XPM6A/LapVCuYUSRacPOD5TXujNcxXxKmIIsEtDShEXJ7JG2xJIleYf5/2lmqZdv
A/xK0a06y2AZDVKonV7jua4XqONA7HhwoHczh/hOQTE+fi3GCu94rm/Zp+gsokz4
NQg47IhH+BqjKjsJjmw7FMAq6Rtag9z3rcACyMaiIJrQ9aaibRhhrXULAEi19p2a
XW/iV+tX/V4Y00xVBiCrpu1av9Wy03bk115m30yxIpj2CSHbpgAMb7Wn5lJWgKpn
PQXcuHcmURhRXPZEo+5VR7wUdBnfmBVMuvHPoB4DdTOrgiDAs6iWD8iyIcbScsWh
jCUNIv+AbY5IdC8+EAV1+KBnxnyX0LA9ifiAPAFMaZgk0nH4Q2NPHh4XzGzCbh1p
SLO8ODTJXjORI4f3keCXF2RUUSkCgWOEr1ZBsF//LJOzVj6OBoq8OssUJECbgc7g
CFhVGafuYrO/URPQlfpSEjZdXRpIDf7yI2xSWmHiBbm1pd1KpJZ2MaJg+Ey98P56
p6KFS0B9sZIT7bFCE5fpte6qzWCwlSdiWlzpqIOKAdGa8EfeWruGbt+GMO85aFwd
lkXPASPJMPCGp1W9Ev5g1E9Ix5cKJjzoP0ioPrgIoZ8EtL3m1d4sZUaMqSi6fqyG
u2Jvga/1WFtmTo+IOcjnPinEaMim0yFid6oA1R/8ZfiYOhvXr/Oqg8/sSozPfLay
imhPM+l4C2Grm7lS9QV6VYQJF4nsD4RXM/drAAF7w6nNJivngE7ZNtEIZqFnF5M9
E7zzb/hH/gdvjwvNLPdCH32fRX9wrwzGpoZcDRU912w+zB7Z3Inf5shLGIyojIOk
n89RIlAfGJ7kE7UdAOU+wrRw5R8nUeh4ylvNzDzLqr+PoW3/Kevi4I2WsscpFf9i
ih+psmr0bp260h++v4n7GI6lM/834R8F+sDuMjApxRL83W7tF6+Sv38t0P/4DBBs
ujGD4jJHY+r20eUWQz52C3XGPkZo3uzMCSL7DRdbQ1wlgJLMJtylWHyzJrrY+Jgd
fxjDfd7d50q5wCyu4JIi58yqFsFFj+Vmf3ePb2p8Hf1vzMDxrU3I+umIhqrAdATl
2w/CW7vG6P/I0W2cX9LHEj3LFfgfdMoXb4qrJV2+6N5sIepUl5NT46nvlaLWbMv5
p6GT42LPRM5lnaVVTfDUySEUSNUePmBkBYJzxo1NXJY9uUBJEaNJ1iTuA2fgAbD/
YnuINZfluiOoHYPBryXAprfozJzqbPiAn2Dkuz2zM/RMjISPBxLMp5MxUqY426yK
4WbRPI56cusWheZOtczZ1VucuYA4JCrQTY5suv5dt1u0E+Unw+klIv3i5RZTYQhU
mAdsfV95hTrRjq2oT/qfBWvqpsql6n/Yw66UMNGYskW7Ih1ay/VsoQvRoZgzgovv
HN5wdqdZS9hDRBR+d8fkHQWPZg3oFNuqRAJJVz43DbPgRllWFTjTpM/exCMyt0Yc
ZeZq4fR60Q+X58oFlfXtWArsashKCWqztIt7gioxNBry+E99QtO+xXWebRoHWHCd
xsaBue4b7h2fFAcDS4y0uwtjLVHcVyXHAp3k9gx8UNkI2gA5z6NSpJJceXya3cfP
/c1wY++e3j2OXsWsaW/dJjAE20q/d3iWDuGkmO/1CA4cGpaU5DUpZb0UH8M/Q8jo
uV5PAoKfHAnMVLUeahiLdjwoE+lLIUy6QLXJn6PrioSCh9qCrdW+AkpRUdQO7Iuy
+UxAqe5hhPYWfim+1HnHM8piZ+lpALbnuujnlgICrLBf1rYWPOqgWc4DZagepmXK
POVFdamdl6awl7WRiCtB86d2jtbPJaUCPoIqJ4iErAw5iBvjkZCgMMj+4AidPnBo
Rl0Z+Mgiyeh681vuUbjtr18mEXS4OZgFV21qdD8lCeWvZuCUukUnTK5EnTsEwVLn
KQEBaq2rBHKaxxZD74fSw0XKNVxId4T4Vjq7rj65jo9nGTONo4TkEdzJLyNK18O+
dXtuZdYzKpFBQ3UwS+BFq9w8h4E+QTtBVl00ngt79SIAsE2f6BqzxgciW1VGvvt7
4gbxW3YqtyTa/DPjsdSAwjxqP2uvMgwDV1KQPxeE2iQNXSylbgjc2oO2kARGZv84
UzkudbIGnsTo5VlqiJI2SWgo95NehUcQhV+500WG3+Wb5nVNkeS7ZGO2dgqCoi67
/SqgXxQzFw/O2mPVhLP7iwOcg1vWfSGbNPApaCawTR348cBfnuBeWRfY2NpHvwMc
0ohJOSRUwAn9yFZFKfXt6R5aMNuRYPy+18Dy6nCgCZ4wUj/wy9dw2R72ieIN3jiq
YHyVYG+COuGNdv9vsVwi+VLlioqLmGPpc2ZWicvbv7nh2dF11tKtT8Y0pdlt5MWw
zR7kDdOHeMx2Wyn5KqcIlUq1gQIySn+ErNxHAbPzWwqqoWkzywr0454p1Z1WOV/G
uvithU4PibYs4XljFk1H4BEDUTJgFc9Bxkqpn512kX2GVApqLvkfbZgnJcmZ891f
EqK8ZiwskHokRbZT2dOs+hNBMlVQkofjnbFmnh+7sdETCddlTtzF6aeNn7Aa5c+0
NrPOYb7BW6deBAroOYCowJ3wPKLOI6D3VaLtv48/R9ZP53/GQKuWNdVsn8gIWiA4
J0Q1ynBHfRN9eOV6SfcQLf2rAn1sOz83UWo9h3Jqxo31aKXl2AhGWChBjNt5SYWO
/5d4n2GdCQ1dF/4PiQATOVE5A9Z5ogVDl8h9uhdLSO6irgeC+58WmBo96Z4tuGWs
7tykI3Nt/T/wyYUNEdrDSsH1utxaC136BtNdzvbvdC8gB8sRzfZ5r9plp+txbI0X
wQMIAm32pkykyLwucX5NY2i2rfmtT9nDQj7tuj4Q/oO+F3u4k9hl6VmrPj0kGk8u
HymuttWSgpCsOkoRelp8uNRmy6HGK0p1dMmtvgff7BKbgG2iy7iMlkrPh67p27PM
WblLsP1nCG9NhAnouQi4loDiQ5LXA00IjS0al+xpvQO7c245ynSnuPN5vW0fjbL/
E065IT+c8YSNwzmQYNMoHkD0QJFJPqwNFRWjiua/zvvrde9/ZN7D3a6wL+YFHX/f
Xt7FVCWYlzEY7kYFhFE28f5zXHsN992RDVU+cyJKgv5DUVNAKrEgbsqg1BwI+F+j
z06IQTcIB86JcJ9m02lXvYPJA3z8R1Hu/FNJ0aCowNL8OREZzg3/tSbDgErqQWjU
KWNAIK3HpeXM1K7wTDdRy0AoUgXGxdhYQkszbkW7t71hh144l+lGQlBoq/Z7SBvx
z2exUkFGqilKBMUnruiQ5ETKRGNAArLUPHH2wpvAlxZ4gr51RQKLHAucSXQq87Bw
U/R7OnCP5RFmLcpI7A4lu6a3BH4QOBud8SQVAa2Lm8QAS0dPpyXdChzYUWJ1njaC
EzckQd4btWT94sEhskl3LVnWVBliW2MlITtfwklM3cyEp7zsfWo9+kGtC6MOYnbv
w9/7R8Rlhb9BmyZrJmmqC2bUruL0uYpoz83zapMw5CLtQUyGQdp8CBSASodvf/VQ
+vpdejsw7/DyZbAi60Swb4imd5nC6Cb23R38FH4DKHlQMEBBpu/KhSTuMs3hFlFR
szWs7xeMBEbLv+88luX24Zkxp0hplFo50PU4fVbvFT5bi0UV4mhEz68MaeUlyu36
26WwRXxm/4u2ONIpqOPKTXo6whA4sUHlWHHa+sQiw95JOVG4ljlg7pr4wvXNskfH
R0Br89ihva3po3MdOsVyaIhNcdMWwuznelWJXSMBxS3PBdu1YhzSQZd4to+xwpaC
1j2PePnFFRcVzT7iD5/Rf9aATCLkvNs/mBrK8Hjz3+br+JmG8K/lvXL/JlhnH5D6
b6DYsR0u664oJTyKMF77MRusT139BZEcuOAsNEcf9XLXA23k1YWauRv1Bljrlvxx
pNXmrB0dlR8nUw8xdRs4/jvX+TJOqKN2+X0VGvYsZNVS89l/CyoJ5FqJ/brANcQO
yVqNYbphBhnwCWF+aKKQ2dTQmNA50T165yTmh8OBimEWWNJWzD9GqSxgVe9TuyU9
wyKesChtPn90f1wB2I/mrA2cucU+Y9U2OB3Plwv7htGm5ssySaMLoPTdiJ+lVviZ
YURBPDLCGipuSmc7KpnMuN3v9aziresNWXoYvWy4f2igNEhE7OuyQFm69MPHtpg8
aBn1QJdCBc3w7GSdceH9h+21lT20e6zAMnY25HqLGEHy0fThZpX1roUnD5Ie8YzU
XwbE3JaWLOY65LmnwcJCvkWQ13AqaOlek/7Hx6S1CTydIAx0bCGIF0gpQx2MOMV8
Dcw8WxMvYE6YTD9nV9TPArA1DOY6vkIytWL7QbGWmfUqnl3TFCziLYTmMWFWENWc
sKgQwXeleCA6+q9ttaExw9Ap0mJRe28NUG4mocfmSn2pbJHBMWPbYNCcT7z320hx
CMa1WsSg//rpomnR9oRjBCBg8tO88jy8v7btgZ/EC8m3HYgCIYanUxS8xNOlKEAt
2mWvl1WwhH0deqRMrErbG+WxV9/1M9r7FA+KwIzkPxVsXZxKv9bl6cRusBq7jdB/
FX0qR4FNbgPlOwTEHGD2JWb9eGBOn4v9F6iswqtu9ABgaVHf8HtE3SqFGMDmb154
N/qUCgKyKhJiW2N2lYbH+bnvFRn8K3hin7GndWVRRzDayUaI33ucVMroXsxs9Ngy
Huut2JBIIBQ4LY3nDyoJ9QwR+XOhq50r08aCfm1vpcif3mhuAW94l8xMIiQaQD6b
n3ES1MpGptWI0GGjpd+e9seT4JC+BdN3ACGDbzNu9ymuS6/vKaS8/1Iimi/G471K
eis+uZf7Fcp1cGlMb3b5m0ybQMyvKYJlk7XI7t7UM2iaqpp+kwOdaVVGNRLHf1wU
FDDUGXqSMsd7XRc8MXr4eNaC74A7FFZjm40YG/mzsxoMqVmGoEPt//+dmcHOABds
GctfpgoNjYekh4MoEOwJH8+iOm2h6es3Vih/cVJLUZwDcd9hscu6LYZIgOpLJjzt
Htq90uYkgmzKxuzKzF6xlF5X6RpKR3SssJ3EzOV0cHkQ5LqPkqk/T9HnPAmimlyR
M5BtPbGATgl+gATgPlnwXfR3pOa6+81/wRh7W4F3oBcf27WseBK5ki1R4YKWwXIj
jaIY5Jyt9kgxuHqu8TwIs1yuzV5E50MYW9OikhljegELZMwczapqVnB37MVZjebq
EzKuUFccjf0yvyyMgSPxP3AFXEmrv26ikdfSSZ6xoUlZQva74af3Ov0/U+D6F8/b
UW28GU5VxU3YrIifoVGx6+2Mh7DZJ7wq0iDEvL4CCAgVkReQ1+L3XywOkCMHM5NQ
z716DC+pjMSmqiRr++AvyMUaP2/wJZw7pyE989mggaz/9J0QVHubnWFjVeGWh0LU
oJMum6ss9yWwxK9mANmdMxm/ubsA45DSWZcIVjbYNq8IbZUAyT06WDjZVomD72wD
4GTh8kC1/C5B9+PfZhtc5nmQpwYhc6PJl04I60a1VYd8fUUAiPsc6C4QuW1nz7Mt
Q8WYFcvKyN0anMLPiMqw0igpseTBCpY1Rm88xyST1dWDIDdRLbhirbC1EgkuNfDd
bBnx7SQx6n/RFSxd/JM6JcPZ71cUKgaJqxKcK1sxU+sh2pjjQGo7lQA4Vopo6Fb0
UQDQSIP8vGvtuc/q0b9tBy6Uu03vxRhtDIciR/cQMJ3tRBZ+kt/VRPOxg/sGhUvM
wDWyGppGl1tjMw7NImzPmp74crA4q/WJBKliXN3ZAqB3ntMI++87A07OxkSA+UeS
4nDNd+ipDJzvxn/7C/fpqP5Etj2Aeg2h1gOAa0xkTak6nelNUcrVyR+MFHCWslo/
aSWKP58ER9i46lsSQsB6S8iualGc7moIezZEZlM3LaTsWnuw24wYG6haS/3xKJPA
1B8mO9q83Hqww0D7Dam6XPg7P6Nu8ZcvV/XzKlBBzMvJy1DL7oH0Q3x7TtVdqRNC
3svc3Jg+v9dbRSqZk8kZ2meuBP3nU2I05R64s4iWStSdd6wScJokxEXqHZ5lfYuY
3u0D/ossBZ1sPxYvrSqaB160gz8lnnCpGOSEhr8DaKBSQkjyq8OAfVkgUSuDjFfD
hrLDvlrIatcjchcy6JzAcMXMlOoc7QS7frV5PSNW2u8Jxz3+BWxRBAXxd8qEvijj
27w15ZIFj2KOFtZ469yakMEy1Cr3WN2coWo+2mp7vAaGZ8grLNGjhJ5XxU6ekrRa
rFCgC9qL0LT9RvezSMBkgpLOKKq17dSJttzmBtNGh/fxRZGE48egwwuyv4H7D7IP
iSjSNtoRvY/3wTALVBQBYSC+eUrZi/9DQIEFLih1+dscPiYjXG00X/4pLUrhfYTk
TG16+BcYSu9CBEOUhBBbx9b9iQWH/ACKJ9sOWymaHdcTIEaZUo0xppP2yBkr+h5b
vvW/0Oturx4aAIA/pVCCXHBSxOwrhQf+6BBg96n+YYnIfQNscIbPhezCcG3pTFzK
xKj/ZUQ9wYne0ar2RceqLJPN5kZZYikVAAXdthaNaTgb9M+sqMXxTLum+iKLw+ui
G1gIBS2y4F7QAFAdtWZ/aFOkjAZasF+Z7ejzZic9GoRnUx3+eHB0ARUOtU8AfCJf
0g0aDct0Yvm5dxARbP58IBJBu8FK/0B2xfpgWXUM1Vxx5aDuFSq4pxepBx4nvwdk
8A4uy/Mz4SyWvecpl/EGn7wEgTyLNSnI8aVsgv8OYjJKHJ98k2b6Dh2LoCxGh3Bg
KOZsaQD9lkzfhJ58d8zJIksJ6tgNhG2Hj/95axjMMzLS3ftOJcJe6OJnNli0AxZG
cvttRDlUnAyEfzLvCILfyxhVPZ7XSTnLd9xbzPX+KoQyK9Lfw1m/WRmDXhcTxFfa
+Wl59OzlxAqzUSs+dcPSA824lfQqLiQpvCMqLDCfmGSaB1s7FVFFRHAorGWNgU3r
WIT4+PDUjE2M27gwdGUkyZZ1CkIT2rMFBy7sHoMoySP6I6nebEdLUYEa0Go9ERzL
MxdHGrhV1gksIuufUuoVwCOWdjdGg05PER+UeRjC/6ue5ixxQiTMiR2hI4nXZ5la
CSOfukYloQBAj95msVusQfTzLBf5OG/KX8b+tJc4a12Wa9zML3yCAEIL3k9ukcxH
R4IJGDN48DRn1Prl+0uXkQJsGYx33S5WlDJfFX3plYCcBMLug5KyYHfRtPoSIY9c
w8sAnyDOovPEK5fQ8prGKY4CEqt4ikHP5hqv6d/Da9+l4+W+7k6cmvGoWinR8ONV
l/s6VyPIOHBI2egZG1I7qxJJPQZUgRnwrUs82qOhhj9mXuZSWE7qDaaSoFIBMFrp
+AiipFogIzcg7aDzPt2Iy0jHaBBlj8xOYZQSCd2G9gBV/a6E9EPPNb7v8Y8PeKjz
RUL8JM8PNBLpfiw9a9xQWZntrxgxWRWO4O3VuKbV3ioIfOdUI3ILf/b8F3Qcx5Ww
aEE+5v5eYMFbHwYS9slCZngMSbkcGmBBzAf/7FHjCcjeOtyOTgs/rZltyzMm+x1S
vqojzn3YQUUx3tsFw0npM1/OmKSHhjb/FYTVaRg1RZFhDiag4XlL3pi7WIZz5RYc
uLcyvYRJQ8Q6dEjWu/KweF/V78RWhi8WSpNEOjbka/b83YcPV299qfl8C7k6lvoP
pwhdGtAP0ruIUJcVYeODMVD3ad7OOku/v6xfTamWP1YP0rN4wID9lxqrobFILOQY
FgXORcHjJx57WQE6RogO675DO8oD9I05ai95jlGAZ33u1xcjUsHrqzNyZ0P3p51g
FjTREZLIqoQOKLgFWZEPeJyLd5j4zi8cMxS/ZFifOIdZsF6udoPmjqZLYa/+p+YR
5IDzvb9jPe92n8qq4PYFMWF/ZPa3XVPP74G8ENzZhN8Eu/IXKbxp4g8qPO1wBauz
XIi0HAvkv3S0ZtHvHcOlz5hkK1to/E+MiBi4zpl1bSfqTOfa/TVzWOiTE02A3vZ1
vBEwxzQePWEhCiz2aUWx+F8q+pYbi2istKeSaQDTUTqMNu0QP3YAbdy+fQJeSjuD
qX1OYVTMHCVeK/UuNQN+4X6Yt9C6vucMfe/RH2rQSpQf80DKrEA2uEAts5lq8/MB
gmE8CWD6PxahaPiuxQDdAFEp7HHeyt2zBKTsQwNq0u5PgUcIXtD55mwxMueHgq5R
Cn8y59PBoqWxICsi4ybMGI1Ckcv9ZL7CojR0TYjTlVYkkW0NzxR3Yks8V8gP8EOW
aG3WTpUnXHY+hOVUmK3jD8hL+VMZyuVxwYoeZsJxHGR2sZgW7LtbUIvS6qhvsT8a
piExJSSP7zed5sfeSqosxOGDz15/KICiRn4pkwECLQZ6zhT8M2Hh9a6y78/+b4Mi
FwVHr7TdPNnVY4Mx+I1VO+R64VMrdcGtcD5ud/A+LupPsSI4gFn8L1yDBrqy9Th8
cvVV2l31QZ0vlVzKwxoOAFtQr3Of+RM6w9+0xpS1z0tSa8BUzvxCzr01R7cpeyJy
k5uzuQCJAr4TwzRprQ8zcZB9ymKiwretu7E8093cOkxRM+yqOm+FdXxqUmDN56ma
kZuwJjxER2lYcjsxbBkuHcufEMFJF+7WFwH1Z6N1OUZQOw8Pbr99qrvq8r8Aa91u
FvJXUbT5TQ5/vP9wyVQt2AGBR1eZsYYPxiL3aU0xrUntBomjNr/jdAiOiFIb6+fS
jw8C2J/IwM1PS0a5vOIhaSDy9XuRRoBwfbJEWueFeB011vaDqghkEoUZhjANpP99
sJA2wr5wJIQ9KC4xLxZCWua5rczgt6fHbLcgPVna75d7JjiSoeCKydVOjlEgBOtl
kxyxQU9itN7tuD9VO3p1v+UOHXPhROYNqZY2BwJtbZUCV7WJ4ANRl/y0opF+DZpA
oSEjQq7RzKqRWP2NdH+DpDCCA3fwY+1Q8D7Nz92FrawrSSnPkoq80Cd+WCjPR00c
F09C9Ej2fsvbIzQepITl5xL44WksZWCfR1FApFT9Hsn3HgkrG/1aHZhcEs22UrG6
LF1tI7VjNmsUDFW1Qsbya7OyzXRuqFI831mvERkBAfc3DZxXquEhG/WImXDDudGg
LeOLUIj5uFGzHmTcYWwye/EZsmpe+K/yexoR6suFbAEwnq3aF3kKoXyIhI5xdS2g
FjeNzagfoTisw1U/ExKWSXFruV9NEt+UQWMujRhxElvdvTv5RxDE9ptaHczutLHl
wf8wPdIfNVCtBH6h7y4yLztlpBRGYomRgrg3v8qm4DRT3MVP050SL5mKc6OslVqe
GWXiXoqMjZON1w/6R4VPiVnJCBZXQ2nRGou80j0HfdTU5tOFDUF+Lpz+lr80jJic
4XaLMemmhiOdSVj2gj1gZ+SJlrgioiiTxlcBOFgMi5zds1qDCVebHgL0GUXU66rG
zhoc+m1Ct1cym+dPSAD1XCnZ9+j2Fg3ik+7mAqGgUHcGtfufg8OZgnSMtvN2ACED
Ea6e91ZAjHAYKbMhyx9UdAMKZBO/1kx1Fr8LgH1dYpDOeHQQSTEIqiJdQ1ywWXru
TDbpM358HcO47e6l34g7F7e0cI6CWQ9L+YzNEJ0kBFqFxJ0cnD1a7hl5VVHarRUT
F3/CCrIzicqsQ3jK3OkLE7vOLJ5/MWbPNnvXwysStA8AIB6cG61SkNQfz14BUBdh
r8x/VCFSqNpya+pm5uM1KgAxRRIaEydXBjMdTq131EugP5k3XYEG/TqpTurIK46l
AelBQFFaysQbp+AQqJLbdu2VLh1JJfPc4GChwhEkB+MVoLHFvTkpG/ygXKbyuxdm
GbbDHGlHIM0mmSZsVr/I+EEkadGepmlR0FZ1Akita6GjDutTe1knxsI3Tm7TBZRx
QOmnpNWEX/Iy9eJlDImcxmyz8rT28G0y9C++FtTzSIgNaIuX4BvYhxX4CRKtYwHu
aen9PXlLByzbFHzV6S5lHuNyDsNWa6O2m5zfzPi26LCpnRiWU/H1mXP+Q/ePcazj
5JBcSKU4Xx79TU7NmEFjaUOHmLd6mR0e3NhkiN+ZnjY1upMMFz+A6JzfJLJXTuWz
cXFANfRxYXv1SHd12uccA7UK5CE0u4katdmF2J9n5M4jUSkAxGRkCGYvFx0Gztw7
yIVOUWQg0DUa6oVL5gFdZFrcObL1ppmHU06G9GRkwH0uouqrRSBzAHx8hnbpuKpF
cS15g2W2VOc11SFdC2ahgwX5MKp08hITQMn2U0ZH8vAVkuEllbCrRvzf2e2Ban2v
NSmCVBpSDwqD3PITiVlQojCgjP0ZVp68n7DLjSobvq+WfwxNnzetaiS4Pc7MOE9w
B0DnLX3gx+fnnwyOFvIFguloAh6yOOMgxqAv2SlygoWaBJxCGm6ZhBj3HAUy+a0e
v9nrv083Vd4eMxv8dmuCm1mwP5Ux28OJgKozqJRsDTmxSQCNPx5IvvYsPKoFKRJd
geBRGTlgL5WVYzq2/Pif6LIqV5xwN46W/fozGJAnlrEqP0CuBkD32dh0SR5sA3zQ
tC1PDOpbgutX3IxRLP+ayQZ6qYFRPZntn2r4PIgWqvWBZQ4ghUnjG509ZMSlPQpF
dZlk/oS0cYZLhmMHy/+/kc1r877rcjaU0R+4iNKU7Aub8bGj5YRSYlODjxK9aiIY
oORH/Fviq0l6lGQ/XoX4AbkMLGq59IqEt6z8cnFMEpyJAiYHm1Anj+pa1J/8v5M+
N8S82YvQmSO5mAubgW0Ue+w1CUxSoHP7D3dBqE7YdXktrOovbWMiv5ILqvevF0AD
NVcAnmGN1IpcnFVmmGVcrz7AfJrOdGCU+7knjYFhIOaFpIL7ggEeO6UCAuSkn8pG
jAVhfyk4KdeRy3BA1qH2qI5Y8EDuplxj0arNrENP4/AfqeaHJsc/d3si2w6HXV7F
SbAAg2uDdDEwxJ/jTDlEvZePmgQ5Za0nTDQdqGDkqRcQrSQG3Q8k2dDQ/+aP17bI
g6+49UYQtra0I4CU83CPi8Bnja+o4yNxC4Ov9KaZJ7e5rxPQcLjcriPl+q1zipVZ
lo1iP44eN9VmlzjPVmFj7EiPXph9EwmM7yeYBo2LSJjTrKRuOAu4IB5TRJwVmhRv
EkgoWfbSZBeyC7jKo7F13stF/jyumtVu3Tmb1WsZ4eExYYEd1QfYwt/b+0NazQpF
X7hOaghXaKcIDj4b63y927L1PA7m6HAuD0RymKZVyD1003kQWhLPOSnNGzZz7k9i
fL6hGo3//bYz6P7n8aP3BGwW/fY+EOS8T7y2p6Z4tPv5Pe6Q2KkzRwue1vQaM91o
HUgG5XRG64/AxD8IoUFDSqpqnjYI+KiIvagNGd2Xcvj6cSMKw1dL9KR/T6G1nFVE
2vXGhR+ABFHccle0tVvo6zmrqoItypPuKSorrOSHfYNwy6bLX6iyzm+N04EEdMYc
YcT0t8mqlNrUFjeyT5gZ1mTENjCuRDTPRkfrmqqhz0dfn+G280/B8Nnipg1HArFP
FZvGaUYmLiAT7R9mX+dK0wa14iJ+BxdvZc5HqrA2KvI9Xwv0MY/+ndfHE9zyO8mS
wwMa5C04gNf7Jg3L0pGeedXOwd7RJimLKZ6p8l9QfMJJVMBACyIXjjboeOlVKzJp
y2/F8yYIcBBW0wdQnjvxPEVQJwENAtXOcSY2SbMvZ5zpVnttXuAVccoHuDOUFwb+
Nix1GciOl/3ZhOoUil+WYHIpUC4ExJ4OoqP49vEHRec3h9J2cCnWhSmifRXH/u5U
3TanSj/G5cyc/TidTS1UoHAEAaL9PCROJO99SdJ++V/ztqte0S+GGlTdQOM8Rk4r
bR1NmBBemrrhx4FrE7B7KnA5HOd17ZUVcnwIJaVE6W08hIvgkrsRRpP2cBY/ztfQ
mouk5ekfOOLyrT6uMS6UCH8auJBQdXA+sDmaqfGFcukFmDiBDaz/W6J+DPRqSoMx
JYAvSeJjigN0u9ZZqNio1CAviqXtNG+Qno+FMVeGE3fK3mIPeXyuKcF/oI0mGpKq
yPahYtIIN2oMK+tlLZaY0kpzPDk+BxV6/TPiJQu+35T25TGzrvf9My5NZIkNRyot
dLRCpys9+07L6Z4qrsuzjFhWqdbXgj0XW9LOLuSGlI7anAY7L/30EHyhefthQDaU
/gpsn+pHVZXbwLjnn27r1++Cml8z94KOApRmJ7Oc89DoxlFs8jKrnu46VQ1776VI
QwmG8c4dSuKuiaF6QDDLu5Tje9gY1mvAgBjZgfCPDQNV2C1XUurISCoX0f5UYDbf
zdd7Py+h8ZoeUxgiYnjJwtjbFyBdquI97lDKRuXIZbj/nv9N3w6ChNzH8B1c68ko
QeFrxOXl015kDCsftv5juqmGxi0lgHaLHPDZ5d2QEZpRKfeYpCLEoR7vGlK2UXXd
Bw6O80w7p29b82eS2NoG5dKrdQ/ul7mb0P56RuO0+WMJcxPacNI1AmVRWvhP9R81
dvj1bXOY0A5PfL4Lxq7i0B14EiENLaJinHkmfbZLw0yQEpVipBtz2blVvh+iRdrL
0OeX4fLfJ78aosTX4H5yX7Fk+aO8iWP6CNY603VYvSgEoF8d5Ctl3Q3RBDLgC8gc
puTg9xVrztHcwn0DZK9HHXhjGMb3Qwj9dedXI5HvwojwTKc6Xyk6spujQx11642N
8hBS4TwMSsDI6iM36QDLrD03omR5OWeVHOC7lfaA+FWBlzFAEhCzlw4KpNpO8x2u
yZ7VhL8DxCzF3JwtdnrH5o+tu4Ja/XVb+JQB9D8fre1Wthy1l/NXoQ4vKCV7xEB8
E9bI0g5yl6M7KByh1QuLzpR8kn7e+OUAHGnDoSEXw9iG59CzxW6k/8v5UirbGH/i
N1wE9CPuKC1f4B2WlvGQEwbbaPo7crpLyd1T9bIvC4s4PiCSHqdJ9F0pHcf1xTXd
Gc2z/MD9wunxzyTGZWVFQkaVLzgYuwwipug1pDVq+QoiBPfd0aX+zrUv1/1dZdYD
HRojDBcNlsoWUMR2/gKe10AAh3glcTYsVWVyFa+f5Al7SeAX03ahR/+pYZ7GcXtz
2j3c8eGh+LK75d0z3IPd3jx4q5jABxxmulKuE5+f15519FQfvlbmG8vdfuI5fBWy
mpb6kYe+mwmqqZ5uMBVBsaEBZvG6A+0zjeFstz/5vP2vY1xCK8ONTvpW65RsPDRm
yI4DGFAT6/+zn+mWLBixkkXasF9agN/tIMkyk1AK7Q6E+djSpiPOd2DOwKEvfP7Y
KNEuGnuLagMV4CJK+5CKXBK1s9bC9skX3/cMr+zLN5+5gTNx1I/U2DW2NcgrRayV
MgwRC52hGZOIUP876U8D3Ptp1ndDP+YtEmccT3DWVB3fa0UqP7YCQoQ+8bZBIpy7
2jUT7twFNptaAk07/zl0gpKwNx5IVB/9EK9PwmD2aUT7qUjMazClJlJlO0ZgbITj
04YY5xiUta6cSbzi1UA5+7RbNukhhbCyZ238C0+MwLI4v2Sceq6JRuLvSIJRMKze
kyCorSVh4v84N9LPnsY2ZpUvE3qezrE5sx0Xm5DxDOyPlsLzTZsO0u/q1mfPyAj/
3d/Z93rvry2NQTO9sLt6BIeHKOcdfURWZVsysfgbirYXq43A9gfUmhqXQqp+dygO
kGXPpPYv/0W2+B89FzlqXG8DhTlEr/QMq3EBaoyXFRLfMGA8AdlxXlfR5IEaMVo7
mChPbd3BXm0JcQTRJJ4zwQ+tp+zAVK6EBxHTHXhxaeIS6lVc2QU86S2F9WBazJ0Q
nQGMA/aEPfaE7ob/8AGq5pG6VnqU/6VCiFhxaVfZDR2qg7gp+6BxvOCP20nq/3WS
sIMuk28k9qEyLKDeq8qhg0KK5HV2OP/Cvzs0O25CkglwXVp5PgavsgBwGWs05uwm
wi6tpiPAQG7ocHzfoADlh7d3Y8jX2kYe8I70JGI14/ZMGTqRUNl0o2g8x4v8ndaj
hx3/qHXqI4TgaYHGfS80SSxuTQkH8M49FWEPmZKBww/jrZf+oeOO3F6zvtolSQkN
iO4a8dEci/ueCgtnoVI/GtcpQYrtunelcIjVE89swDPLCVS+nyERg73yfUHnynAY
o61Rs6AnRiZlPSKEv7mPell9cDQ0NVF0HmftgrEsVTW5Us/uz4WmrRK8Bx6GdeL1
EfGDSgp78fUYQxqwmcnWsgn24pt/YXVyJvS9SV2RhKBSm0+476lcq/Cnzvimw+uy
1Tpo1AvoJZ9ar9I5xGLRZpam/tooGPGkW0BVVjsV+W2G4vIsvnmnqSq6EkMu+j5D
7afgxE5F9slWC+4H29ZuxaUXRnBHsqzD2W111O1IhRV7NiGi/86shQB5vxUYsfdi
F6PlC/GgjfGzlPyiOr+YDTgoBNtbs1EaMe8DRLMoWA62DrS37ACfE9Dm0LbT8h9l
uEzGPcdQxCCpqZjYyJsJb7o1sLa7tJu6WKRx4j7qbT/ak/9ATc4nmmuwhqcnxSZf
9g3mdvPjZER1RFzjjLWje1bLxw/7EVAaEdtWuzwitTQTX+4WbDgTTvCD/Ir3CYzq
cRlfGEQr+g8r8BcuYK3BohfSgMr1Nvkn9NCahH2AE6/RLlEL5T3EVD48/uOqSPi1
DSJkEd6PFAtrIikM4axbo0yU8ePFZw3HZxxmwLO/Jsyn1FTbR7TDE4t/4zOtYuUa
/pHRNaHBZs/eDrgRdmijpLBcTt2LNGGN7ESfCmt/eN5Xc1wMIazh/mGIT9uJ+qWk
UTaIs92a6qhNaSDjziV8B5EKaxwhu9oNDdOgVckrkqKr8on4jM1Fhg4/ILy5ZhY7
fiyirG3GfjYmiS/LFQw47UW3l8Q64jy8p3164jpE7jF8VhYCn2blLBZE4ubcH5Nc
BAUCDuaL7+ISHqL85WsPUySKF5GoHy7afZIp4hJCz3hLUPogWySzuIOqSMfNQ7MH
mcgAwieFlpYmqocGPqn3yrp9qHjrbsLN0bi6NHIN87WgusG7bVn+7SjC355LM5wx
NH5hmnze5AMRzCo/9obPjNGx+BiuED6d3s7yKXtef/8DN+hIK0GRN03DC6O36wO1
710yZgD6Hg7qn1zn3lj/m6AlD7ApnqhsxVlS/zTSJFIXeaUlb16hl+BCEOQKigvL
xvjmPW8VU2QjIEZqDV8sjMUY6JfQldCO3kmDZK1nNWxvzPjWdbYTHNWAZW9icCAs
xF2pZCgPZjmjsVL1ZyDAM/W/l9gNQP8y9hYHTbL0E9Iayc9Z5CsAUEbzp9IQczMN
lXRCOwaik7lxPk7jTy6wCLDBHwd+WlOmcN7Xw0BtMFa49xoxm+L3F3dHsgpd3d1L
QFqiF7MvA3crtfhemW+6UbYzNxF99BZIPeJAKMUxl4brPfDPMNWpqyls6pJztuRi
3n9s0JmDAhdmCXDC5qPggmbMjk2zFFt1hS0DJL71YNCBXGVb/8xe/9W0oJlhZ9We
dCGuyXYHloLgmLuzH8zazVN/YsU+AixSwN0ZK7+Wf95leHLS/MIgowTPArNhHrRC
w/v/qBZUf4EvGB1+fjJeJ8bvRJRBXJeikTrpuyk6fwLvY7HKUyzTMmA/jAkPX8Wt
7MCQ1lOjyqRulfEr+XlTgx9N0r5sfcEwsjXA1g3MkB1LtqM8kqY8j3kL5tHES8K6
z3P8CtHPZkm09g3SaMnc/qmifR7vnfWZDrJYP8eqxfKVDbXa5rF51zxMnKMm0KP7
jApdhfcuOuFEP3e1fnFjXE3ZEoR0R0eywqtRp23p1tmMPkyQQlfh6eIG799GzDse
7yv02txyn7POE+Az1ulhc2v1p9uB1O6H1FmiTlb6JyCFgipBdJPqOzNtZh4tRi9N
284N4TclJ/n6WnO8NBJNr5b3q3zkhG2mctsis/eOAkTpClxgumov3ojfKHFEMXoQ
1LUO5Yn7Q9GUmjvMZkr619caVvZY+IgprpHOsLJ8nWLcldQwS1HBriF7hDtQbwC1
Q531egd3y/0h4Fy1OxY1WUkSXm7ERZ49r85PZ4uW5W4Afq5Yttco2spzyKMnSehV
PRe3bMWylp/qikiqmKETNxoym288AIbTRyVGVhdWB6lRbNWibqmlKBPsBrYB945r
Qm1Ma0ITXnGVWq48EbsweXFPJcpOzszg8FuD8B+LFYUP6Os/SPwzYHm428NvSEyd
dqjwueWlcAx7aUXNvdl/sJx4nc3zlu9w51mS7B4H1eTUYoIuczcsg7c3Oml/sRoS
hHHSHODLpaIMN5+sq7Ssg26cVIRwXx/ZgWbLUz3X0f92sVUaF0pH7bM1aZN28tXf
+SjzvIlZmqBItzWHrEcD50BeTvmBvbgjPlPBFoubWz70dBRwgsm3a5K8TBIY5OIz
XprGRP6Y/tjygBnaO+TU47m4UN7YnDk9vBl7V2ouDmGNKcUtEGMOaRFgL734ErAU
a3xjF5Tg0AIPk0eiCQp5sa9/n8qoNEwkxUJnYxLguSnUlMY1xrQmcVidZSvXN6lA
DMi0UVG3hHnk6W9KBCg8GtuZvpcuZ3WUty8ITmBDJS9iw5XJZGpFc11o++iEgRF+
dHQ1xAIhONEVTmWg0BguzL0RvI7o85ULakOgzRo/l/FKyt1F7QNQTGrYZoMLoTFI
UfwtgVcz1eDi/mnLCsW6D1BGHZl399YsVricVcHldD4V8L8e88wce4wv6yESg8eG
kqwEcVaXmSH9iiLsK0kGlMwoa7e6VTen403m0h7KFV3Ae6+iQudQcNIDtfM19luN
QZEk3+i25+He4dKo/PAQPKFE+Z9hqG8EUiRLf2UEC7nq4r6ttuUBq39e7+o+ig/b
ZOvuWwzYk/G68MiCjLcG1oTCPtEfmuNwPUCt6u9yRjvvigDsaLAGCNYMKjeI+R39
+33uCi/VTzBnyNsK+pGX3EWYsfAyfHuFovc3ia91ERml01TqIqcyFCgCVNiOJ37V
C4HNsjg1kKIubV9wakHNMFi8EcgLOy91PDgRWHOoyElkvQkrFH/iImKmHxcmRO7S
P411MB0YPSPw2a8vO4HTV8e4hUIoQuwr40/Q/GMgvj2YWT+jQlKxfYYYsUKGUcXW
UBbYHRf8o6DYL+g6rviC0g++Q48kQvjSm4kohMf4XP10KvjP6Z18BxlD2lpQUVMQ
qG41TxU1JFbrbtYjjaGGnVE4HnawRyKCtPjL7Mn7KSWvHNGUvFW22UzOuYOCpuxT
RuoX1W2542K4fT3JkUPPOE/NC4w7SCceyN8gjckfAR9buYtB2on8DiE2yLizNMCY
9GFweaxArhx/ls5DedHOmzRB26uG7/n/LXtMx0WXl7v3nceye4gxDNTd0EQPFGm7
cxw2hXFwQOyU9+Uhlvx9OQF0w3YQQFXTsodftKKmBxoA6wye2yfGctDmIGPYtGBH
Socq5Ho9qpIPItFJDzFA/L8ouh+8yulXbCY2UX5/Er5fVvU1pWnO4wAGxWcp0kGq
H1V3VjrDOrrCcrT+HAcQW9hKoQ2l8IVRGEPKHnd/VvZOxdTakpKClKYHwuMUYmEt
ckbVJzsOsSfVQT8giswFKN6G01UTtc1w5ODPkK68NXrGAFRGlOxS1KBV2Z+kKjRy
vrxSBEROHWTROnUjIZGOekGsFXGpKzWNU4QtYn/aWaVku/4a3PgHJJ+V1WoHPLG6
Kl5e7divGybkahr7fwUGEIss+EKNVj562Js3GxXWo0ZGH0Eu1OyW969C/6In2+GH
Hoda5ekRt5XnzaQVIYR16TtH7eEGILPqV9Yz9htJ8hnYQFKEw1dEoFX6P3ycqmX9
m0lfS+DQDLXhDGcNSkWE80v1vbPTS6lKbaVZlwGGouEFQDAJZR9VwjP+YYKsWW1S
la2eGPMOhJ/Q+/Xk8nzIp7iJ2ST1ogDy5w4hR+6Rq/5KwvK7F+tkIE2kYMfVJsqc
yGPElwXOZmp3onsGKjf2EPWBN1qKZbPbfzX1lNAcIIVH8e/qe1o58V9OvjCw9Lu3
i+3Khxmh6jDi67uWfhuHG0v22mPwuMHUJaJTdR5CcI/sKRixelz8MLbbAVOZuTc4
xFeHLRhadKU+NnKjo0MSjXaMm7xRgSWAFiyY+tVAbPLvJ0hqfkK3M5q15Do5UQW+
ynXadtjXE+eVBC7DtSbcJsnrTNzwEcmEJVxjp9MbguTJRd8r91Gk8TFtznyJKOih
A4tAWHZPtLSKrQ/8YtYqD64R7ODVN7SbI5L+CNzogV+a1mfsTz0e3Z/v4aOLW/o6
t9DJRTPwJoha3pxXDrH9gkD/ChZF8nOS6Q24E3SQ11QLe6Sn6S5jEiHivhqt11Mg
XikRzpQBCKajb/pj371JzqtDxsaa8iUTUUzhCPJy0rTEdO/At647Iir6PD2O05oF
EW20unH3eL8TUQPwyg8FLOzsEWsxGtqfbAlWVi6IkrFgpWIAnag5Nl/iOtGMRhhU
WjR3Re7TZ4FysjMsQrvMVrJBDBCJtmYe42KRuhkj0J13zOssG1e2Tu7OyERozPLT
F6GMGmPjLzAGMqxvvDlXrVGUMwob7Cocc7sdG5e6JA4DRsSVNMU39MMJd/PQWcuF
tYcNlHxBCAa9VXCfuJfnLNnEaGwjnP5WAUPQ9PpzorGhcAkhb2p5Zm7tEZy+bzCG
qM2rnjK2NBxkE9/doMozvv8k01YbFAImb7qb1VwfqoqLBMzGPt6jpSQbiaeMifVo
4+Y0ennoVr4k0pYdaxc8ZOfXJEie8q7r7OqVZhsFmTNclMp47NyZKE3AHLnqjEC+
sq0PKwcdLaxtXsd6PU2//EXGoz4HAeKVHbjtywq8JDbE1WBmWlI08ViCw9ndrpTJ
kQtcijk+VEcCK0wdaQQI3iffyWv65azzaPau+FuikbD8IQ7c/mHED+4+pYIbSYFk
tIF56X+7E8AXMMoZRmcn/Fi7w2MWMuC4gyvqX7dYbeGE77uZFMIhyi2MqGO1h+bW
WI3GgVobZmF2tqNkbftINubkv6pQ/axlXuDNTRY2Q0jYYPOVH/AC4KkiOh14SDJ/
AQ6BIYx1J2nTUlf2EADGOcQsk9x/4CswAEOUT3uMATctbd0l8lPu4DT07vqZ0dEO
oSpejdylBnTDXOCQp6P42k2ROuNDMxSUxIcBDIYtkf0VjLmEKEAa6z0RYFlVJgba
aP7iwVWvyIcGKA9NSSg0C5DYHeYurYcS82NAl/1KC8TKTTq/kAsnip38R2FKhF3D
fx9l/xUnjoM2oGare+t3laHQTQVQdUIYBp0HOUZZMtuujU8kyzsP+rRDW6t6ZYPF
gDOIFuDXu5dmigzVuMN2x8Lrf9U/eKbRdTO86Vyq4nV9DGrxyh81MX+Dz/XmXpGR
T6wrkxwo8DyCAy2589I8J3+L3iLgJkF9186GzGk8ILYkIRIi4PIijgD/MzP9TIGe
Htvw+4hKBHRks3hXNDnNbU13r6qq2VTH8oiLafXhF0HPWXbuWiTCEcd0+HDhsLma
PJ/2wQprbfq6CsiNoAwYGgrWgkiitSd0tPNGNHklVattjGVA06F1MqtiGM/xt2In
Fixm9sdc1v3wwPgDli3ioFPmIs1FUiDVOc4gGVtqpBa4Ft/AzYRhG29NSaVTXu5C
JU/cuSFRhS1wEleURpxmKPrFPTC9tLUapM/tWxinXt0/FIypdOqbVU++W1gNfIw0
GfWgwHKTknp7W9qu982N4YQ6CtJkdD+AW/J7CgZJ7i3r/a96xh+A6Bves8kJBM8d
I3yOqxsXEGJelCRC8PpL47F9oVVZqP3boWoh18cDi4I7CXBXhabt4D74uVPJuLI6
hBFjLTaWKBrbB/nbGRlqVe7GEMPNdPJS54tEN29FOZPdPAGDcihIwvq4b2nq+Loc
DXFRxbAvWcZYc27spYdsG3nquYMBSlR6eVYCmvGT+gYvRNiuoVUut32ktVYombjS
Ad17Tvbm2brSkyaFsKUr3g==
`pragma protect end_protected
