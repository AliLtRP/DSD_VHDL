// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:37:10 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
rj0ojmBn5r0s4B0NbD/xQ9FuHFz0msJh++nwf+lKt/OKwVppmOgNyfHXGrbCLHfI
FJbAQAFdeWkMaDAGyD7Pm1af2yOyUmOWZ8xm2q0GC+aywiPjxY7qj3m+AONHvA2L
s6ctxBuxPq3DyWLBtRNEUkTOWi5xBJXgBNDg5sWZ3u4=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 112656)
CuCvZPNWvVk2iQ6KFlWdDKNgR7S652NxeTYyYDkOUIeEiZ4fhh3J9Cl9SDKdabET
qUrIw0u4X1I69CZdBo9h92EhxS+s/lU+fE4jrHlJSar+kBrlvyuRnPnop1Alh+wg
Pxl9oqIVRB2Vk0GUf3IDBvpOSgGSafYy9v4ZomUZk51gxnuuBm87eNAq+xCkPFNk
lUPKFC2H9YfyXVRhi+5tTyd/m1tKOtflj1x2kLcfB+acUGwI7SwRepSZBMAxn9S0
FptqCs7tTlKaMS7YMXMwN00Q2E+hpJbG6OXAbgbVVQlvWG1MlKsM0PovrAZK0nSQ
/ksIp8yDMZ5y1bPDTCESJCJDcHAAtyYF6ovwbcy/WkgzBj4thabBUPHk3ljFJmVk
U/J3hP++jLxbue611DdWhN17OFw9z3QiGxrm0vPpQMKWnw4QRsN+OQqNJuBsLFTC
bGxhX8TO7Tgjmxoz+Oy6/fsaoyRQWyNxkykKHqHZseqPuNooNPjXvZ2L2FgIfyUs
S0hDUVfk907tEzB1TsuaOPUUsVuLhUFwZo0MTkEwRfq4qgq+Hin093bXSEONCUDz
5Ns67whyB81OmWM8HBPIepOCoEcpV+wyMYPN+nSr93hmeYmjxsUspdzIqxtqL3mR
NVOC6yxB2/jRAGidkNk14d+obkQ4qnqf25WBiGZnFYdDVnxG2Th0ZvFSW3q/TYEM
aGW1zMmkBnh7sEHEEzN6OWHLqyBAGAtPMI/y3SzyptGGObF9jOQ/zNMkwGYJbBm9
jzU4aQBPJstNfMwZbiTbhkhpuFlvlvRh7On5EmjJwWJG/pVKGr4hDJEr6f8q/jeo
YaQaFkJtDI/AQCKI6y8TJRgxQu97gnnu9UkR+KDlovViJiptLiVgV2LqgJCLBsFp
z6sGSmpXEyBIoMG2ODJ8OAC21Xcxm6ATW/cbERlgZdR2CLb7ajDc0DqqPsZJ3X/p
gmNMyqyMA86symlI5VTQ4ZU5wqLToqQs+Hv8aD5IEaLHLvMcOzHJFmuQ4yLiXdq+
3SvVI4S2z5yY5j2oV/vC0dPvjNYMCSOKq03c7T+mNLHLvJJByU8B4YbHGCyrf73a
1y784HBB13n03AHy3jQjnQPWkxV1OeMmm8wfzsdb+5Ho6bnWs3dzBaVxuSKsfMVC
+mAg1avhmBGk+vpAfP1zyXOeJjj06MSTqeXK5bonNDa0VsBFIeNOxQO5E9/3U8pI
GF19jdTFQvyGJpg9BjcEZSCeLta3DCA3wZT+6Xpwsoj1XSi1NmkMQDd87Jzeh4/n
OrJIK7iVS5odL3mL06cAn9jYpRDu7TehwHjEPp/vIVIwXMSxDRisDLru6fo+44sG
VW6b7N/d25vdSg0EndhlcjBooofwp4gaF+8Ij+v6kCdJO6MVLg9Zqdd2+Kb+geYL
/tfZOZTpLxRQOcYlFR93GUrZS2m8u96N29s4c96emKUDJvPfTnEQfonxAzHx3Gpk
HbQjj+vG03rwuLkYt7Ynh73CXTg4bRfh8/PugAuRNfoQK3wJ1OolK1HcDlsxqahs
fbXC16BEGhQpnS2zEVc3WOdnbCm8K3Rv/mPg2m14Ad2BM2f4ubyk1XG5yoXyiRkp
fnjH1lL91GQfkrO/9khpxz0CC/RBbRyoSHSt8EohlhR5N+AuoNq3K3X3ndjrwJJv
OcoLD2Bqe/qJKPyCPDtW+aOdlfwzBJ2mz+ylwEZyhp4+vVyP2Vl43biXmCdQ5jWB
TivaQVImaK3gtoQO52rk2L4vxD64UHTFZc9kPMQvhoWshuM/CWLuIHfGYZZoupjo
WIDZlenBjWOsceexpZG7+JgJvVIkvNvHz6CMRHPqgSASfAEFWCFtWid8Ee6a5QLo
h2D0daoefNRKXUKKXAA/wiGsUsxbqyZoIjd8/ahhZZLes0NMijMyQR0r0SWURF2c
ysuQFcLHO6769HhL63vfm6rjMRzCPTX0JAOPMuYXmzSzf/puW/BCcmJmrhqMnbcz
tAY7+Mu4tCq16nrmyIgvA8Y0kHQfS97tLggYrvKzcNdITUIxvj2Qoz7kZbqkbdt/
tbfkk4UK1CH2MuZBDNxrNd4wuZeG3hWlVczDdbEChGgjEE0/wdXsq8UXY6eEv1X7
7QBZ043hN29h26D4kWlB9oQEF9i1u6R4FoMX7Ef9cbWeZQJ2Ggg44moscXuTYZVt
CL9fx3f8M3vIBfK5iJNTm6V+dtQbBL2Gkun1Vo2O/NHAv0n0sGOt3czxJPGryhhK
UpYfun6fxObc3mNBgMjiJJWKFoWoyxg3XuCz0yc/3aFZ8ValdhAOR7BUwmy4KGYe
N122KN3rtann4nWdWE7pSeMhSBmEPuzaLdr5b3nj5tNdETqxT4piLpduhVSg0CGw
FbX6uXWzhZqRnEavydPbLpGp+e1H8QEjvTCOvlsKU/37M/nOZk6i9C3SjqdL4D9Q
8cVxCXi0wPKvCk+Jz3S+pUIGPNqLHg1vATagxbAzEE1U+M5c2b4KeG7D6JagKWkL
hi9ApexWjx+DTfC02zeQoM+K2EDcyIG/0Ji29UzmYAQqJjM0vN0qK/1Cz1tepTcm
KG69OAB/pVxNMK/6Zu1fWkPYfiqOJwRo0OWlOAotHOWpzUQatYz4r1x69yNUJIII
cKsCje+mxmVdcLjLUtU98DsR6nGcupntzyxJEjjdTPDjt4NEDPbBaS+ygomz0oob
ccCeEi7Wzgtm4HxDvPLL7iXi+ext3DeH4h82w3+gzJhu/EFVsa74wV1chP6zKw3D
OCIeYXfCPfgr/8YAjpamhlt79QxaVqPH92Z1wU8tcnVOQ95Ny/JYEESyBabB3+nt
hAebd0745VafOdOny6CkDQdTERHUl3YpLw61sx/00zThWBiU0a03szSszBZxdlhi
QQXwcvDU6KghUf3fwV2I7+arHlJRflwkJ3MriPwbL7ZJ7b8ILXdWWrCp2I6rH1CJ
e2AWZ9dh6rLNflNqeTwfsZF/2IKG4UjOwQkmljRNHsmYMjrmSnaMNP1f7HtwFjV6
S+ioJkMaPzprzhWBaV2RDWhbNkH2u9/l+w/RnpiPMKQU/s+HgT2EmKfThR5NURtz
x+LSU2Gn88yCle8cMDRKHx/bqy1S2k5kO6wLJ1Te0uW2jVMSqeVsEdGHBMcHsIVT
FEvmfNki974WuXKcLMxgmco8Zafy3PRvJ1ms9D94gvJBJ+E4IGBWvZHyep6JxfDe
SwdeZNY/hroxAtextiMsQROv+Q4OnSqC4QUdMm37sASrrqGxfRAuRcNjtbJymB51
yBaMXxCjUlRhHt1J3yVbg8QpIfOwuNKRKTJu1GswcQ8HHEER1k8Ta5r/U0YMN0Dc
Ef17v3rChwXkXSnlTpkmXA2EsraXoeCeLAfwVhW4GRRxdjLCV2hNsRg/olXG75XW
Ep+PediMYzRvTg4+t+khqrgTT3/3lan//NOPREpTMF/C/0TdzD7Cr9C0+eRpdVUM
B24W9ZGz7G0qm3eqPO1L96S7k/GH3PKnS3k5CKJTR0EUDtXDTcTuvqqU1tsnFzGC
OP59SqKowLDDoFSqsc/AE2cPvBqP4lMm6nppzXD5UJf/EUwUPqDhD3njH6TFiApc
O06qCwtnVwOHMvd02Cz5draPcf8cwDvxoeLpxS2AktSMwA4K+1GU2mRJ658LyR42
B55sBYrP8p9vCw6pyoha5n8N6Jt9OTsS5osfMKz8JevR0w0YZP/m+bpYH+A47xy4
S7DlEyu6RlFCqJW4Nb1QfXN663pzGFdJfCD7rN+r8amm02KCB9YjehrjTw4Yy1tC
HPjL7OmtwTWadK8n4RvDxCjI4hcpeixyNle+VrgH7eWgHn6rwAu44EVJWAAZ2aFu
LrpPAEPF2XONUv9tkzUm4+Oi24LPI2idqh+hmns3By/KUfgi/OaSFlYlTILZ5qLb
YfWugCCOWSUSL9KTu9qUD3ZGUSFU+GZ2MFbKXJb6udD6IevQI4310SvtxIyazGC+
K9/gJYa52P/baVk52lmQPCgFMeAGcoVk+8tcAF3f6z0Hy36NrucDr4DhJm2kAtrA
UolzVjHecU4byuIVn2QSk/B4h9OG9lGorbOlr/foYQ3wFK5RvzONH5hDqhsPz/Ub
osDBiNAQ4VKFjKRsguO7k/mXw2T7eNJhi1mPk45tLJjyHf37YdwqlltFuR7sy7tD
kjsPzRkym911nWbnheg5yj0HOo98ELFmi8qyun7kdYwk4GcihXJay26ThC0m/9Ww
koOpBw0NgSJ46Z/tduLqcs3AaTr2TKQtEL7FcZp9IMGPcuXr3qyJw6xFnUXpRShk
/VjUrhd++bexwy+I0fwjWs2Kff57SVUjJllopRmpdFv+VyRO65q6XzkvPbplUo0S
mffRafKHq4pEInv2hbQDUpQJCj3m1hjNFnQKxG8DCYmZiqlfLMI/yKYiiDmL+lbQ
DE8YX4cvGhe5yts1Qs7aeEde0VZ9qXC1mflJgAhjVzrnJOHyVKKzyjPDvEaQOb+0
NmwkhbbJFk+D6yQNiiDrMrNTX1yAAyqbz3icNJUtOK6CxYqyazTYXiiOaTTk7uh2
Eo/d816p3CIxb/NrQ9UmCoMnBczgslI0Sb7TN1h73wxLnRJ6j5FHN5eeUiyYds8l
hMC6glYl5hUV9cZZGjVVUW+gEFypkuQd4SPDYQsE23f3LWRr04yiAvcLoQtT8J7h
IfdCdqJWfTwXg3T52iv/XtdMK5rtScIcmHJIi0Ta4+poW8KglR7DCBSy+IZbXv3P
Z11/IMfVMn3S6eKNtIYSCIbybXzo78SOScJK02TvNArdXOWuIQgnl1ixMpTqeEnp
S8jd7Q0y6Fq2c9xleUycWLIGvxie5v8p8x0PeaxxW64Gt2Ezfa+sjSlS0sM5DjBW
No7vIjNg9aoUelKB+0TvjXxmXMPRl3wzQZQY4kfNm04Nx9wtVNxhNm3ACvkbgNB6
UEY5QutihP99aHsoKNJzbDndwNv2HhEJqyj/0Upu0rQEUrRJNYwht/21a+ICeYf5
YkoCLJTYuNBtxAxlkzOhIhy7uea81bPj0L5umq9GNN4QLzx6M0scEs61KmfuChEM
dRCCCZ4li72vxxvgEMgQbFBe4b5mmSnTzD2y8o9aftLgS6GqiU3RKwaf5WxZbJFF
me8jIhT0YHPRS9ZKNW6T3h+pIGw5vAJ5nm7iqSjF7832kAu+T3m8zPJG7FZ8ycTf
KU/VfllEfhXWb2HSK2h+lZj2p8IqbMBlzlKA6VzpBy+qFKgBrJufObxf8spbXwDz
srH1zyJNyWHPgnavvCyhATJnPIpdYqB1eVi5J5YnDz+E05L26hpH3YGWVd5ZwSmk
Aayr3xmz52qc51nHiz9yMbCr2X6gBOGysgycXlly7LPoH+81EztxgP9SYKEyO1Kd
eVIc2nvvx4OBNVd21P71aIcI+4xZXEmC/CRIUsXBAYQw6dE9RsOHhVOCFhyxjV34
4PVLWQwrG7j77bpStknHkbrUas5HbMM2NO+xYMfeDHgKaKIbjfetkhhYo4Ki5dmD
G7W/3OqBj6W35nrqPxb9cle8pFlWm7zlg5I1944j9ejutCM8+CNdii6qi0En+tGG
f+dUm5dLwe6rwwoGVDxsD0vbkn5SibddxQWX5ipy5GVqp1CtF6v5wHfED2gz68KO
kdy3+cNCBSrIbdjwA9gzvzzzY/C/R2CChw9YjwgHHXbEhX8Eqlhba3G2cDcYHe1I
z/SJ29XpRiNlEfTx16HW2QVP3PgqZANB3bMlA+VBuIiQlLa/dpjw1IfPIytE8joa
5ar4Hbx0GIB9IiLGCUXEtGkKUjPuRxFNnKpICWNEssUOWFF8wfdoXXOxWVy1zVwK
qyuMfdCo1w6XcgAWVfJoRE9Nmq2rbvBbtEMlMT0q6/vhO5e5IlRHDaNVsK+0YUIv
4GPQ6LlSqNHAlgKenHgN7SsdpRnGLQNvOe455xdVZmb/bg3hMSUmz07XfC89XG4I
r0BUZJk4qoWFQXKXjE+9WMXWUgX9G7Qag4JAV6vmk50Y7YEG8hMLD10JD1FWQBNQ
7JcxfVLMvEqFoU3E1B5coEEo/X7Qtcs4POBQDIopoVRZV2OWlGTwLlF0AFbxRGEG
ZDq1rYhHK8mKUbMju5Cvw6XDHlJTC2uxh/KyB3GXBlZXACqHadPJqn0cZmmkpLwR
x0X1uYiTRoFeqnCwjHT4ETnqVh2cp+z2SqDGsaLGjfwBvs6wR4JDiSin2mUv8w9p
yED3G+PMdkwnCb+MD/cSq/OByF6qsmMk978Mf9LkumgM7aKa5TgOac4q9TrXhUA3
aK0kiku35OkU5jTnlr+3vzea+aZfXnxe+O5E+QY0IvkI48eN9TLYaRX0vGRDrsVS
sQgoO3r7EUpfxzCXalQAE4RBz/zzqEvKfmK1G42M8BfUwW6kUV3edLz+0hL+kFbn
ywRbSvo/dCBTYMMYwdV1uD7MtBm7/o5nsIb8qAqIOBQyG6qyfS/7RUZ38pukzcqA
o+XIKWrzMyYc5UwuxDwdOI9cZe5/7Eag1K9XDxBQBc1tIib9T2eUYhwU8yWzr6XU
4U4TEcYYqq/gkHlAJ/L/ybRj7CVm7fx7jYoinwtlga9SmDssW4eaxDlCc7YPwq3l
sl2v+FucatySiMZOYnIV0ysPT9O+RIwWiGG3b8ehpvfOGG3S62qoxFTVUXK1kD4o
Ga997ttRowHHlD7NM/xoGXOJBps7v9lMskTo+PCriYgOUgKDkShePUvg53GKXGzd
fvlO/MNDRvni00xqoB45dHkBRmtmVf/9R21+wYbrf6tEAPuIYfaiPx+jaMWMcEnt
9ww8Jk5xZHdsOUvAj8XJ3X5TjaVyKJzv/Z5GI2rYhejADnlYfDbsMSzKH7HbLIqA
MJfStENMsGv72rcPs8D6cMk7Y1J7syi6z4Up+l4fjW3o7h4gw7bXmu5/KDVRRTDQ
lzpxjlF1WTJYB4ZqbMyZZPshiaLv6nmrUwoHJhtv5kGeeNlssyEklxWPkEFhApns
Qq71wHB7fAcW8/dTOxESZvm+Z4DH9ntjOh5cJvTqfyCexwYT0oCLTOowoBZvJbgS
MNOb7+0xmv2lcZbihiJSOiaXlIMrBqNBZOngGekzxo3B6udAkCkwENRciOO5nRR+
IiW7ErKPs49edQ/Gp4KCGzXoTnIZ1c6HeFq38Bls3ELELtrSvJlKnMSHhjLKKKtz
jI1077hKcspwzHHUh0pbFo7gZW7I06wW90+LVeX+W+uqzFkOv7h16P98lWBIXuKc
R2/YGgrKHiyq4xnKhDODkwdUQCoPHDUy7FHgZiwssLqmNeFY8Wu0/R6HeiiNiTsk
EkWoS9tLOWbce5SvIZfAYugLSsldcGAnNwE7jFaGuQUqkeT+qUH2kth/U8GnYvrM
5c6nZQAPE/M4CtfelMEcrHwiIuC0v8NnNXen7TVZOUs9Ckkko9qHMCmmkwZYMbXC
3OwJquaXus3WcwI2cWvrv+DVNSGR/7iimnlPmbgUn859gVQJtsVl44bHfxd4gyIz
iykEjInuXnWMqM3F+tF4XyQwQmDacAtnfgmnDeIL+ux/ZzZEWFT5s+2oiK4rWYxU
EaO96NodlK6i5XL/+WL1UD9G3h4ylGzeQTT0MkjM8UBv8yxpn/X0xKlrQLEHLHRH
52Z31Mj2I2V3VoHNfU1LDQUZkynLPLkEV0+dBCCPfWqrMbsA8qUmBAsawFLn0acd
ELnGAYLric7XypT/+uI3v8Pgn3SQOBJ4yLQ7FM5stb17q2tHvq33fOcp6/s9aTrc
tv/sKaLAUPbsvHNpeZjDjae6lM2IuLINaBEXtSMXQgwXHsiRXOfeS79EHZop26zq
r+th/1QIH2K7moWiHiz/4ZJAgOzg9X8OOLriQeAmGEB/E+IuC/y8IcTEOsLDkh6w
O8W+gs1I6GM0ROR+0hZfTcomlCxmalWTlN/rtikFEPa1Lz+IxU6XjXde3CqP538q
iU0jD3QGkINqi1Vjs/UDKIlXa2yQLXuhuHDxxE//WnKiz44Fpmo7YeKL95ODnuXl
hoNVxi7kwNkbdzCmW4Fi7St7d4b+EicIBL9wn8gzpv4ScICSRUVIFOfK+XDHtbYr
lG1y9EzkvRP1RracmeqO2Jc8nHj3GT4R33XsjOI9Tuqe8ydEsUMRUYhDy+oroCJQ
5vKVzbWiHZmQrJfofomjuQb3XKBOGKxJ4vExu8XwEwup/zeo38zrmScxV5pafxj2
aFlDYeFHsdc2Xp5PQQc1InSbSksMydgHqXpKQrTITK+jqUJyqPtlriOd80bhdTrm
cpKWEb1Uob0i/0fk4RZ1GsLJqBFTRp0NFLufWKsX4PRFZPdz8Qr5XQCAEe0uqmR+
IgaOcN/a/qAWvag8Le3hdmIL+iKh9dFq6e5+YydMdpoCLsQIYkQYH38bTDU9Tgej
lRgCc68NNY5ivlSFgKiZm67YGjbkkPlQC1ULbe7DMUQtoBkJjLJ4VjKYNS2hOI2f
+FmOIRQf3apo33lTz3W+nVeo9g42LlgYg61TxigVvadVS4JKBr6TGNsB1vFCu3E6
hVlwmKifqV6owDDrfRZJXdl8muwY1LCNzSFDbJn1bYIhkOZz0eOoAdg3HcGev+58
p8688k9Iv1hgLBNueG1wThxpLC3ldDT6lIj6d+zBmb02dD93AxQsDXYdeQV3WskR
QWErgtQHf8JFhvLFjEaH9dL6NLRxfElnoPW9BkbrNfUAfyJbQf5izNiLHM3HBwJa
970mcDJ6v9FpCme5doVNSOymdvJQxnw6rMR2tGezl7O6OPWnwQZrKciMpe4YaUBT
k5MLtHD8vfvaIEZ3L2nYjE4zuRGS36XDABBUHBt14MzVAVjisg59rJ+LxkiRa5eI
Of6SUuC4sFRxyYGJ4ACev0efMtZle8i/E5W+i9OKr8s/1HRfD67xSnGujBj1H2R7
xWaAjpluNIA7MtzYnmDVhbkbHzy24hoZ3zz2NXKeg/juWSZV6xAFD/x2H0IAZymz
fhv5zkNVnT2tf4YmLw0UJeiUdpSJMzQHbdbdvg7coGN7bp+t4IUNSmhDfUIJVpt1
eDsVKGGGtE6dNMKRAZ6G+2jrlPepbbzi3A/UFK7nCSzkSgPRQWzgkXWBVuX1nPiS
+3y8dIOI63GGKemdYkccjNcI962jXxkKDigyi0mwTbAO+qvMHj2zuV3iJ0PlLg6J
XMf4MCGGcCz1rWnVqFG8YVWFxuyJPXcgZQNziEKeEaLQx0MBJzK6/olV9nrqCI0V
Rf2/vtrF6IaBpXtHRe6rZohl1F5bsT7xMfGR0w7LWwR3x+GS1fnMwP3HDw7d+MC+
dWv1sXILIrCGDpQX9eZjjDEUiH8sE+2rbNL+h/vTNNS3NDQuQPrCg7YQPBFL3uzi
mNqFsD/1yxctvxlKgdqE/9eC5QjCQeAH49EB+8jvbtenR1JLnZmeuhY1cA1rodpg
EUYuJEQuXnIDaW29MnIfcU+/jEyXhGTZojmv2wVvJ/pNylXD+2VdtmuglG3GvkFC
yZJV7mwytSX3HgEMGUsl2Ym6ewrw1ZWa0pKEwO2Km1fm/Z8dD2hbBCnJ4RDW++A1
p0GVyCRJ9gTSkknOCtTyDKSpaTCGM9UYgvjCXxxgmIC/m2abvBv85BvvhwctYeAH
Iciz7AD3d90A3N7kN3ifGBtWBdxxUdYbiywsofKDvJsdk/dEqJwtc8SU/vgPLWBE
J5GbBUUUmxj/D7lZ/CzFsHoWrhW0W5evhsm+/KUJ/QvyVmZ/FKHp/Ngc63Me5r+e
4MqAjSuLB4bTtezSIXLNZb0oAh6zCS69DwjnN+uP/a9Ckr6wZuPvAUhnelU6bJPR
gn7JG6d3qXGT6S1GZtgKCMXbXpB10UadWpm1aAasJGnsAwKdtm1EGWy762twe4EP
ySvlxUldQVMWJbNvznyWZ1GKuf/nEY6suzVbsnCVeL2b7fVm8PhBHRk0P8KozisT
Pi4pj70RpzrHPJY7J6iemNrw3xUgJNXT+G2jD+wb6fOU1T+Z16y3oiwVchzYItjQ
2DSNjBQ46nIIZU1qa54rLAWNMmQcWyllQ/xQ+igpV2peQSyzeXQMKcL+C0WlIlu5
BvgMwKLT5RajwqwO2lhy8XJaC1QaxUwcEsv8fTIA9zIbJDHjUB6oXRtvVMPBDQgW
SI1mneVeBGKRInqBQpZ1k84vGxwzMkjV+SuAtbbgw5LK42lRCkFhlj4YrarOcklD
F5fX9fdMeP6uwIRBD4LAeUoPlzfO8+XBrLKVbUJTLHQulcbAf2YYWppAzVzY2enk
q/vFeQdGE5sc063KtOWGQ5spWrxzPDdHVRqoO8C3qfZhohuxIb4LE3sOfNjDCKBL
KvhT9o7VxcdbaYQsI/s7NJCMPjsky5xwpAmEhskC49sjcFZyc57dGarVVKnGJURG
yQmEzauB4ZDuMjDA3STumhNpPHo25d9AODwtpHLt5EAZZ/GxtVc+C4DbHSstbMEd
FSy0qAii1icLZOJYw/ztSZa4wQRN7TzBd2cnyhekCwdChR88VYWHzAc4lzsGIg7M
+/kogg6U/zLiaj0ZZx/Ymnv9sgoE2bG6rcnE+3VU7vEMBcmzrYA2JMyx9+GcihDo
HVlU0VC9vCxhzXhUK2Jd7Tu/dPM+JyKQI0xa0eL8Qbw+9JKUdPI1x9PA+jQg6FYx
0Qcfy2osOVgnIuAtMi+fSYGW/zU8lUzi3Xxe/Qi82wASFHqKrgPlZWbTKwOsibNy
k7dITfX7RduR8jsPWneZGoZa4gAyHBS+PRFP+zU5pw4j0E76yMmwUkaPir87d0v2
JzFsx8kYDBLnjlx1HICl2W87LjENmk8Mtp7RzTcslmdeQOKAr4TcqZWfWmaWZNtK
eZ9pgri/L9KOjh75snUQBL98eRv+3B7NlSGl98NrVxYLad26fGRQtJewco/R7I+r
fGsZDaz1ohbiKqsu+OnveWX4vUmR08jt9k8FAKUaJvEqlXyafnWOXLW4JB5gkTGf
F2l3WaEpYsvVbaYHQMvlnOGcosnW/o2LJ1QPK7oC2nFMTtoO4QhSLzaq9MA8hiuc
7OOjBMHMjl0B9nRrqtJMf1S5WlWrlknxu5J4jviJ9/yPinA96jQoyWlHYEXeL5Ap
wz4eiVEMT3ppTcJIKG0stqK3PnC9258W4gjjR9pBzzvhLnIQy0IS8axNzdR37hRn
K+sOrlPqLqNMleJq/I9MTOGXN6Gl76nOT691oIRjH4TZW0H6XBzW2gnUjYTqdnj3
CUIR0k+Hr4K7SIJAikmlXYQ7Jp+EMehH6oeUiPJLGg/bFbmqnXpjYzrHocAw71wk
WYpfg8Jl8lWKk5yzo47gYmw3Rr6iwb++Jw2BXnR4Fd3AC+R7r6PglfkZlgbvyrsV
vOjeKBwHWAFGHncYujPAQLrwa0gQ9S/ikaDcd1JUzUItq7d96+g9k0gAJDqvEM/e
/+88E8/3Geckd7vw19l6oGa98r/wy5ICUORSR2aVCLuwv95qe0jGMnHZha+wdzbk
wXht60/x/nMzZV3iWFVXWHDAPU9dRyEvcDfRCDRQsWAv3fNMZ4F3Vsx6kAId94rH
TLL3x2D0veGJkZmG4moKV/YocMIJTR8tnz9BRpODsTXe2pBB4W7+PJAzxyrlFNZT
evRfe1yyEP4nGs2FOLf3055zaqHmhzVoau60RHQbM4jZ/YV8+SMc8p/VAMPgIYMU
jZXTFiEj99epA0XZ1iH0bDtM8skuxqUANwB1pxlQwucRbNWowyElIdLqSIl2/qzS
FxDu0w985I7T+36TLqCekODvu1KwrNOZa7uYbiD8Aw/9B4NDg/3k98/9XR/Betwk
thnyKDv8x2QMBoudkRpAgTt9rXnubAeFXKfaBVhD0D9eQ+ahKs62qwFmlqgCB56i
5PYdm7fIA0QAkVPXlnEF/G9pbSkh0gfDm6+0dG6LWdnVu3CTTlqfBWv6w1OitlaU
ZGq6lURbrCoyarLbPHtUqj1y5osQl5Lh0JpHshf7gGufXOEBwKp3G9opGnGDhF5H
qnfEmhQzBqUHguxyLPGw3xNt705OEjvAxXC84qw15mkMZS9BfvLjV4Wd9jMi6g/O
MKlis12lE2+0ZIsD+SuYbgxNBv5VaaxcO+dtCg6J8QieMbfyMHiNpgWKCHVEtOEo
qfRGmwRKtbASnLp+JszQ3D/zXYu2/uWQ9aSEeP34y0ImpY4TEd/4rYCupSOFPtgk
eNqcCjEjV1lVEEQrCEGSucICrGoXIIm13R626zDO+R4fDUEoadto4GJR+Y1VoBSv
UMwXft085Ri1c0UFulU3Tx3MCSA3Mr+6gBCKQm3Q5npr0038q22iM/hheBBvtjJv
dLAjLZAT6osO+n2LOiJJMMcQhUdUQAO+8Be1rSJzJVXP+b6nv/Mq3eg3s8FXh0Wd
jYCrbf7R9mMFw7vjFyA8rnUoWvbQJsWWJogFsSqFsDIAI/U0ebY46puDh5KzL0vC
0IKQuHR+fDXRCKdM3dKjBU+BvXOWhot8W4kkYVqhrCDZirA6A0HXiMuzfXpgF7te
UIlijWwijG7RI8g+H8mO0JIr8J1i+EISLNYNx55pOjaVbeYAc+eSbasBZm7viTZ4
RNhkr94RpTM0iAXn1tkj98pRoRZxANz5n9wwilgE8nymS0l2feXtH2C0ib64byMC
2NzdBbGCqhvzbc10ILZI1RPT/hLQvSrWfXx5i5hPmQ9ZQURBJ3AHhsvsPx9nvdSu
YbHeqCp3jFOzjH7qn/ZNXavPslymIqRxYZb/mquW/hyQly1ifOrfGXF9HKy6xuOY
kYvJIuJqHqsgjhMZOWaTbKH8aAKIKsTYxE9lT+kG8RdY/1Rrn0PATaQp/rPnxngn
t0UXUILKnkxgb8KV2FRNaWJmHKDBTX6EXH9A+7Ref8+DLPsljKOpDgrlONmYQH2i
K66+8pyLogEmEBmFo/pIVwHcELxgn24GKx4w8NsfvMpVipbaliTinwO73AKektgT
53RekhAlUI+Vj0GuvFaAXghi57D3/vYAjvRa6ek+yiHNBHoLGG71KzNDsAiZrTey
DfSG85t3Jd5fv5xbMhL8Lu09PHK+bq0KdDkQUSFkg5MetMP+YyMpSGi8rUdNaThF
qSC+Glc81hlggrd4AhzK1dGVVjmcGWGcscFBcl9cgXNYVCexg4VGkpsPjL6ytxHh
M+UHwYMz/1WHKMHFWEGLmXSb4pztdnI6FruinIEJ4ZiwYDrv8qUoA55BasN5x3SY
XAUUOKRRCQY1pX09v6BoQ86ZP1kC/o++SblpXGOm2DLoDVW0sKnWNGWxzT5UWH+M
ld1cBOtx5EiIHJyhTmlJmQK+Uo2tCpZErzK62uGEcbOtNtsdk2uxaaTO++hDBdBx
PTEFaASXOzLpE1Vle1t3Epg0P1WllvQQFpr5yKIcALorOxPgD2tS2vbV7tGLhUzT
euk4d6PCteybJNxwAJpnwv/KWnahOBr/BN0f/unOZdmtpQIqA7v+HJKHjWjHNSOD
F9q3OPXQ+s2Ta9oxamlCB5oUKIB+eozucpNLYVAip9+EiQcx8BNO1WUufrJJxBzN
42bL9tvtZgm5kqMJazTxY2T9fOoUQlKUoHL7+bwJd0JHhMeoOBr8qd5UeBQ6hGSi
Xjmdb+QatIOkWOtnvvKKo3Fp2Nn2BM6JP47TYkc8rrQheDs5MEZgHvRVu83CGxdD
+zRsDB2iCttHmPPagSHWdES5L5hNDYkw9vYfeArIFamrxJCn9TdLZj0GgAUTL7ab
Q5c8hl7HzxGcVuGKsrfH5f0U+XSIIGL4oyJVbpEe5jIsNdTMskIzX23znQd+ocbO
491FTcvaih0ndbaDp+glucebfBw00K27/PDxskdL22h9zFOWNl7yKx55WSqsBEbu
icwt5kk38gnwJUFpAuYidSIuBgrqAmqOKfm21n3eKa9lgF8ewYTMRcODgNQFNdYK
mUCMexaldQtb/UhomzTZ0SgIyBySwygzkrBvs/O6ymN1VGtqPNGsbCryQ/CJGXnv
C0or4tkhsikwAGjY6tFU9q5+wZlWNWIOBHWAPqgRXqHf1vNFuwn78b7NhIDB7hEJ
Pg5L9lexjmBqfQ/i+VdEPKi8oOH/z5qxBXhsBPNR9Xq/SabEJmq6zkkv/ZYaALOt
QSR8eTyIpc3EPblRscne/FGrK1gHqiBo3cjsAXp7yMaUkCaMDhH3DurNXZ8cWVXn
F+YPWRqIa0i94MlC1jtFT51N6xBv2yX3zuIb8545FfuVFfx4OLjzmsUBmSv0bWH7
X/FnQjJSYFBEk3K7imSY98Pp0PMM8nTH41e0P1CiUmeWlnXe0nwXumX9dX9ORRxc
kkn4iNGgv5D0oGw5CWTJ4PxbHBxnU8NCLBlIWtUKSDq5iCKoAM/hSK+EnNF5sq4i
gRLS0hvUygTEzTykdeAk0UFUcDnWEodQtmW15mkcVXx1oj7a0flbWNyi7ItgO+qC
mbFCa+ffpOaaaDBDu3BbZw6/kv/N1BDE/1KFPm1UmOAj7aiHHatQqdUaxnV6ASpN
mCDgVdb3KERjMJjG0l/ww17sMBTBLofUfBM7oPWqxUBdjVbY+3cgxmwe/01yDN/F
qMz+3rWaoOaCL8k8utYHixeO7+wzm0N7+HA2UDk+gdN78LdIUxDeQt53F6zkfXx4
cxvWC8jIamDIOg9SIg+51cEtEjdzvDW37xzjO9FBLuB9RexioSMNx/7HXbTxPd+Z
j1VAcG9aud9LN1N4q4ETcEu+OCmDS8Wskm+BsZ53ud3XXSK2TlHixnRTIg+kAOaJ
beh4uOkPR5QYUQI7/TaaNs9I9mk9t+IM1gWk0ZCrvr9hJ3BY5dJX27QBZLRkXza1
b7J7h9otEjO62Fm5lkLaw8fmuHnqmSFDGYz3GZcVeuHPxaidAhnbKd6YVr+VvvhE
+F0HZ1MPKQq3gFR328UblCVZ7MjTdoOAVfRHu9YnZvD16Ea6XUcRlejGNqVjNKRC
Qis+11XBhUnLZmqSvIFvhk6Q2Pt/BD/GolwYDzICI7tCex4Q01R9jSJfPrfthMW5
l0aiiS8X9x2sezFwz9AhebYCu5JfCqPY9xSWgkG2reiW7qurOe3Wm9DK4rgAWK8f
bgdTficQWCPp7xIiRMXL3Yj3XUAKOC5SqsITCgdbVEwnV2eAGqKtecg7lMEuZqAq
VoK8WgRFt6HrBTUhysAwLBJ8oW+hiiAWbnp7sgH89iu78pAH1OT4KfQclBqY8Dv4
lMAFWVu9nmtu4EL5JxWDJBUvqSzwgBTfg/pYq0dlrWqQduNtd3ZK7Mj9WjDiCekZ
iBYQjaw8/GITPm2x7pxoZ0vjhMPd0yJKg0FssdHoGBLvq38S/D+qD+tqVitMRfbO
JbzGq8Q7HPeaTmN8xhOXrF4xwm0ndJ/WDZ/EbZQSTUVZN8v4kkQktfgv51h2Tc5Z
X3x4jJ3p81UOGc6WvFa8WVRF316eyIJCpKjiTVS7rHfnGLJ6/cozkv0xIvcSiDNA
5ocIdiEni8BjffxP2B9UWgwQUYv8AUqJY3TwM7IepKWJtH8EM+WV/XKbdk5RDJr0
j31yhV3G09FkEh7Ur3zUdMlInhzlWqZFrTFWgp5gtq0Va0LvYVxdpzSQnP4dsGLJ
FvodsE+H7MwNoFAGltbSgA09g6V0bBTpIuaI2GTPY5/KV4Kx02/DMjwEgOFvtgf5
7IX635QmmGSk4o6F0tPZ8VWKCVjx9aEDR5Xy2KLMcsn+M5fhUtcFxuU35rTOJKoz
r7EbwT2NP3s13phaIcKAMTIRq7CyIarjS79Az8xg9t55LSS9+ZBgETMuRG9VWToV
4m9H/L9dhXPRfsgEXdhA5v6YV3JDFopNuym00v0+1ltPj0Y0cjf9odjvxbSxzuNV
GuruINrC+wY9zqlSPjbIp0dORmSaNgmKsmF7g9XUKZClqHy6+gt81KCEfwjgnvft
AtoHYq2t2ypTtFcfWA3Mooy9l4EIpK8GZbfoQQ8RdMYT+HCxHsHG9uAy/v3ndfEB
J1hyVpDqKM169dvNI8NLx6dKJDh1VC/9QnxJGQz6KR/mtUbZ0U8A1AjmHqGb5YEq
bkkm0P3SLRYGUheYdBWfTAMfm7A8A4WJ7YpWgGomXjodu7rodT6U2z6d1p9Rd7uZ
1DRcHFEEOrYrcOAJrq0wGoXyKiPleYS2O6cCEVSkMucej9/jCZAlmMNStlBbYKwI
rqQT8FsflGPgGIQyzwQiyVXaBieSM7a0rvsHUzFt0xnFkssKGsn4pnY3YwJdmgvk
3mwvzM6vjCoxYRAhn5Xo9gLM0w5WAwfve1/VXZWs1Gy/XhGd/U6JNfqviUP0R5qP
vdOIOFRDCTQzsvhCKgtQGjqrfeF05kyRIAHgrwNIcw6Ro08Sah3Hww26jywOLQa6
kOX0xoJ7iQIw2vFyDJghFteiwTeVi29hNJaK3gJjjGeuV0UzIK1JPLm5jDN0+sXw
KwXRBOaruNJ35rNnaLf4GVwWYQH2gwzo+c+Wfs1cDaNmasiYeSXXsGpex+k88m0G
kcUs+MtjUoQ29WQSqemDAJ7q52xu2nQAe+JvMVX/uNw0HHmjcvHgvv+MMJz8KVdm
yBs660cLFE6SEcp9nrcQdurwnbXqjCGBaxG2kfx5SPWU+lwbTLvOEwnoa1dMoD+M
XQRJiX1otVtlwXtGAcHwfcJY7FY8z+0tWKhZ867EtemDDsGqKm2hT+o+/YUwEAVf
xj8h6VLTiPzSjLaO59Lh8qDkgwFpa0Uu7LBLtLeKj2yfj6OgZHz/zjBo7IZHVr95
ASPTjrQUbedtIxoeSewg2fy6o+/c0+FiWaxOFPTm9A7Rs6r0hbfqRglINwcPVAbk
bC0444Z6TNClXGBJqA2lcpFf59l5ly3dEd1qEO+b6W3XgxTm/h+LVmswzjzEwZiy
chshtXFPC75ehcQdAiYwdpdkheBaZbqh1Hj24fChSj128UDVmdg8Ghc7/bnp3/lG
Dr03Ak3F1/0q4bBymknlzTVppJ3U35E2X0YxpPr+hPuENQosKn/j/2YtMoxST+1Y
OWmDJ6qsJvYamhn/69iTHG5zC3/0zVymdE46Zms+oCJwZTsrry/DzJpa4FO+MecS
MV4ofutYKc5j6aQ8PX/j8PGLsIPH54NW/NePgE5Ma6fdsMXU+cv7HufyeEZBZPq7
MCaMbwQ5gpixLx1szftyyVc7lwlaJBzLEeNQ6qeXStS8sHJdQx3Wagvzdr3pEHYI
UipuPT0jCua9VM0HxR2aO6riZyKDz0qUE5AZSsSP49tG/V6umh9bHBbOCQAlPH8t
y9ne4mzqRgx/zulb8BFbIc8N29/0Juf/QTsn2+GjMmKpcNdHM7HAkm/FNe/mjtiS
GtjCzHAEr1w0w4pzOpiiQu9ki6TdHY9LI2a3aIHrJbnfkGtto41lB98xze+Crg//
XndkGukFhEv17QAghjV5OZ5PtXFWOFqRl3HrKQP621qOXSHmGR2cUlcE9sxScjGj
Egj4lfhc3Xsv3tKKH1/bLj9+onkyvAavN0z14RHJosaCDf/AU9eXCuAYskG9JGx1
Vt1KnvCmRDcwku13kuQRlVnf56LJZ02567z9hUOKE1TkiOCygPiKVrr4idxOYLFd
1cRGyDaLGBf7F2jSl6AV4Gdw4XBGaRg98P97cqJ5lE39W12gY95wEWIIfSB05Itp
px002SzUxclZf6TVbLIv0ccZQTOGo/peRs9+T0Ly9hiBAA+Iwhx544kLJpDNtoBu
16iwOcPSxi0HAXkv/SY1sVg5QhDAsesH8jcMBLMyKVqcEtfFMULE+6b2YyXtBrGe
HIChtKYe3vdWkMLApwmIeGtZYAsxxBJfloZT6x3y2WEXFqq4y56mZ6hVSzhuHRb3
0vsVR4vC8gFjoJ2uLvatN/+v3B2rHtf1uTqhONQlODN89PfM6OnziyGG4FtFkVVr
52AScAEaQM/BN2r9k5y76i6wMhlRdh6aBbQjCr4s/x8sr9iQXmOXm8xU4VE+CbZM
xCcVrXchxNZ2lbwB9cqJzZQmot00yH1rwkr0alucL4PZPg0B9nICQ1yNGlv3xx4C
itZo3bwK9IOnzS6vZN3/LGgpuHoGI6pob39e+QWyUkmHJnV+6OccVTHu7yLM97vA
8a9KRcOHAHyosNYkmyYgJXe5l+5QaS3zlgWy4z4sqDZzKFQnWNpqcgSQaNrJemOF
qfhL1UiLYGYlwMS8PqFIoFrFkECra7/ifl18DcgRsbhNR9cMDifEf0+Q6MTt0gsI
ms4qz6xJ3Z6vmqbIwpW+rxIJ1vExKhuKyAo00OyOVtE+MvnEErQ8bnNJt/OYND1Q
D2XxaA577qVIgAsT9nOxKqlrI5e0dxroqoCqG+vpzKN84tthKOayWbAI7P6atOxS
iAvbULc9ThjrP78/hCpO3jDWq4/6yZNCDpY5A0v+zdii5XnP/HssxheOMcbrj6pF
bBaNxim0+BaI0cI1XQf55ctAHSwkClTPSl+lTzDO4Rs1ZkohifKQqZVJZQekrzcG
mQ8284ozLWOelWqncxy2DdfoMpPhBVe+HMtUgOGD5OtlrFdXf3aKdmtk7v17awRZ
+ofFyl3S4oHn2pfz5LIE4PP+iLCNq+o02aSXSlStylPFJ8oxniRsVj+ynSz/k4wC
oBLBHjPZWPs2fjfPvgxqMJFLON8qssDmxDKdyhXD3GXRJOBy0UIsdMgqx7rFa45M
cNmSeKdLWE2SBZRw1ZCS0ifQk1YNVFqUbtkrkmiC5cjFkaUuBzfXNgTNG+a+W53n
ZKBXuXAZQkGAShVvlFJRouY7C+AyoWCTd1KeBX0Llc80F0oG1bhslX+YpTrXdgo4
iezWoHSbsTdepHdEkctBTcO55FpUYjKq9PORtyYoMzz1DKrGdyVOrOK85Nbgxe0N
UqN6KUWH/msz8INulf80bGoHs5ubHr/P8YQ6jNluGeCgzKbiZXEd1fiHevv8cylH
78chqIzAoi3F+i7VCQas92EZRdET+3WJ1+wyZH98J1dgzFvkiqSTZerfp7Bn/hag
K71AdhZMBxGE0v0JVbo4P8wJwe/WTsmi+4TYWuUHLcL5XNtvRjaoVrhidCE7Fvyp
EEJ8hwTzVOeuG497R1wMjpsAVUBOXyyfMlrySg0q6WfIpHVNg9iTSRf+i/rKC4xP
X90oV0q8ICf9VIpm66oVc0L5zE0tU4w+VN71qvjEw5WYV1e3P7zsnZVTyi8bQ9jQ
sADr+HJMsxydnFX5YrSG/hqLHNsG8AdNCztT4XjHgcnGn3c5XbJUREQtjfyAEdqM
vrnMQHvV+TJc50c9Z0+jSBcLIX83jReJimyspCq6/hkN/Gmc4eecNC4Q0Fsih6Pf
O4Th3qcDWf1a/vJsAbFGQdWrTSqTv4lfOMn8L0qBewuWt0TQtxrxcr0rJolBn+mi
x139RaWEPcuSOkJxPI9TmKCg+W5QbQeqxIKLVsEI7oL11kz9y/Lq7+8DPmfgMp9C
1em2l9ENo6aTS75iti5y0aB5KV8mqQiJEiOjgL4cqV3r40pioOL7NlhNNVFmfQIS
jB1wMgyToqRMkFHJIZAeyoy9XDpQkmNmCZDQ6VFzl3voEs6WfnRqUsfZRrBrAaf6
y7WgVC5mn2fke1S8Uezv9O/leW5iDzdIvOp8itb/YFDTHxc0WO8xo1bkgX83kSeG
FEpliYmDBFJd9k3WwlXQklftZrRVAIwRE3GOVR5hDWJxHFEJnmy3uH1TqUCmpOfk
Q6X0fkyyE4xOzq35wmFNvuttnnT4CWYDHZb0G5PLlkOADMj2TvEtyUcHvcdhNHXO
VblO1PmSpkeUutW+alN4ze1ZiV2CmiQ2/2TX128GCsQbd5SeUA37rfudUKwQw0V/
OggpVrCaUf9hD/5szTAfxs77I0w+kmKnOHlDkBsrR9dO7ovCpNtbrsZAJmwWL1gW
SRMuFrKl3neBoNaQyYC9WjpwJDVEu3YiCDZv+gJJeL+JBptOpW+ojSodn6UkPwBX
BR2fVg9HeL5+gO7p9lzS+mSlvxAiRFfiyyIbpBvN9FGqrnsLL1DcO7+7OzeJpnbA
bsunqp1Iqe64ej+n+aCiRgcNJxXRvysTPTJ1H0vPsveiQKdXHzu/oRwRZ5vMKA9e
f3vul7iPwvx24af9BqpEh+dkVxODZA6828XL9AxqblbuS4XBbX8qM/nFoS0NWDH9
WC6HnNei3bwea9YVlZTEB+Cy9w3pMVqDut/TRpyKvcNHv+YypGBVfvwRig6z27o2
MEU4RQcqyfoYvkASF0YTi5N8pOuiV3oWuLKxmw0HEJNdjxRh3s7lbeAYgP4pXbOJ
h2ciNLs2IDplQM3EVRaxQE2X4FoqrhwZOOmAYCFDma7ArToBhR5stakbd8cmfMFr
c2u/Rc9z0YqbmFh769Oy9FWqB0PjfXJcjakG8gZs74U7/D6dEBTh73vVMzoM8Rjd
XViF0h52mMpYtKb1Wb1ArCRgPEKc9X/2eLcFs7Ut4JyIZDuXet3rOpIGKRqTQcZ+
Z8zxbZzmcmPxdEzYgK8ieUjEwLCgI04VrTddp0h8G5bQOo06msnPoe4LTiO6VUY1
tekUvuoq0NSDM44Z7hI4fH4262+cAtvtWA61RgFo3hy3baIlH0HMchwX8/p6dPz9
E5L8ljsPBLfUIkhQx6YfyBtU7TxdBDck+ec8W7+1VebWaA704Sf8kd7ZWMW+MEzq
JyyN6IdMKSfshyJ2NfzogwcB7V0HwRItQIxbqQGVRG2FEfQAfwNODetIqe40qCVa
O+YdZe9DKlISH82rRWKrhmpsFw8xo/zh2c/hg/UEER1mnVG4Y7hQ2miQEfO8D4QU
LURcIPNBJDm7g8BjIOVA5xivffft4sxkvKPAWoSwsy8zXDPbGkUoeQoaX48nS+xp
L8ip0F977eqhay1O54mOJYT6i75x/hK/B9YMLSXF4YpSkvKda5yg1G17bBn9VY74
hoT7FyODjVyJxqR8SArwTpdnveUWBlAv1MlrUB6vTQ0luw9/COlI8ff/m46gUEIg
TqARCtslp1hp5rPZGYHLK4RJEVK1xtNj/hfw+FAuciTxwdgTGVzlDr6GfV2jsZCo
8QwnvgsKkqBmIS1PxxD6yDWso+CGB7StywhxtjZEXiq8a/1HgfK03NpIREKqdz8x
13Hls1no+REYMGTk361aqqlSiayMm4xThmVNuVxblTg0tK3bxKgvrZeEn0n+5UEb
hOCXexJFbQnbh0WPwdUJ3fwJXcliWxVDyTF0Y8KqHRmOEuIGUnYRoks/SRxtqvQj
FGF/A/1mGcG6cApWp9GyrWAODxXljSnlod5yZ2xk/UrEzZv51rs0MzsGnxj+lvgV
R0RPCWwtLCoA1dT2PekmjD8nNT2rufl41WMal1opgMmZ13MU7VMe3KV/smOUUnWi
RZFrs26eKBUpW5WZyrbq2TnLZ0ADud542gI+OJLzDd4aSLoIdTjR2tRZyA+sVodv
fcL4uaQ3jJBdayEkj9HZILgfEjIbVNN21/+hxTRfV4NqIZZPpitVRo4apmbiqfoP
YighEj/2m6a70I9Ju1OTWpaynz51wbzO5IynYkylh8/l9SKKdhu2UKuZYWLVpLB0
o6K79jOKPiFeSR2rQfuymZgXydBWbowcFbf4xPMV+6/xglmW2/IDRGH6YqAvETuT
BeO8r4WAT0q5l9zxFeEyMyN0cRXqSek1Fd6nrOrdZYZZa+27wSHVjS1ahoURwBqh
jQlNVq/4DjVy+1G+m5ca+xhaJJjjUOgcfSLbRUtkzU/ccJfFOQPbd1Svx3FhdzSu
sPjbdIZWyAsg+DxsPIu4Mq/FnukE6cyngX8BdxDqu4drRD7Q6GJ+JWKik/FDGElg
zkUUAJRllWHN/aY6C7NcRoy8fI5OUZ6lKES4M2O7O68yJqM5YO3MFXpMVSNWDeTd
6ZO0haI/F2b2gU4LE6N+8YXeYkFW/K0lUvYroD/kKDiux68Qg2SM05gx6OViqY2m
ZA+5I/iJ7vvRR+/uP2tQksMP73CZf1FHFpyNnDlnsApGfltFAHl7fxzLSO+CuWEk
3bGfGhWEE2sTrj1Lpg+nRKDLWI7Yj6q9qJgngThVEXT6oNa/LNPjIy6xNwvZj2Ld
kfV8aBF/aSjpi093n9UsX2Q1899+X7gLGFRHpFCFX3gjgPYFyHKyihXN8J7ahurV
RNZSMmyhLR9sYxuN4xrn6eYl8Xha6VBweR+mHeNg5UOfdPHxfdfWJCafpG6tq+C7
wFXAJDYAIDNuxcOzVWAlx+xXUnAbShuFWAV8wlMw8qjx1yxSrrK93gqEktaSpugb
BYeWqis2zuKN0jsxsJRUHPROt+BeBUjDcQ7FiFTELLj6bstLVOC0ElQ0zStbYcef
vUZEJ3aef8ro0YQgBFy41EKRuVPcTDS5atOw3Um5Xsv+RfJe1HHHAAkdSpHquxO+
+XFC985iHkS0Z8zWwWQHXqAw1kLOaI9/mwgK3bUc05JTqE2VL7kHn2pgo3CalI7R
i+r4sqcJBl4akJ8Arc/qc5gyMRLKnQhx6yRPIqv7s1YrFOYuhD5GyqZnI011EB3A
/5//5TpFCPqM+qIoDUd9aYh+U+v6HQM1ltjZD4iSi7HkHKh0KDK7oO8jOi9Hz0mI
yemsTTT2Kf975J6f0cbjUsf6x7I9MJFZt0XVZaKG8GR+jjOU43YJhPlt4PR5x7C+
XGdKEeZExuiGx4sTSVL9c2QuhjtnbW5qn95Ce+9yFrUEkjTllaRnQ5f+GbH/rab4
azOoM0IX/pDev0XH5FhQG1qPmKgdPvIBWiS9FDTTVqVB82YBCwc2ah1ZsAkhL7nq
Or0q6aTaPAMMnQBKUwJDl9OzycPB0rx2M1pYEHc91U/FW5aEwrwdWrgncOSSrKOV
6l5eX++pCfqV+VWco8p+MaKUPXyR5xs01Dcdb3PBfRQa4XFQkQbmGEfkyX5ISlFi
CmiXPs20DKkjfMVSPrd2VPrP/JBovKW06dm0yJJuZc/MwutyN3cYyxS00A4XpFoh
BOubd1PIHdB7HCKjBa1CHUCrhzzQXMh8OELOq1GvLzLeMJ1GXv6sAsWEUicMIJnX
mRfn/LA+KctqoSi5u5MHgKnVnzrwqgsrSK2ANufHKhfLraz2sTNrEgRpzSd1qB18
xn60/p685Oi3car0Ctm5jSQKr888UMu+9327alhf2jDTxWrpW6Evs+lehgbn+6q9
DCS2RmJ84DijyqmOfsR2g71+IR+MbWASjPxTbAlp9E6BJ1iIB1v9fLfYPZZ+7Yur
rsCpyYwOLYRBhhBRhRnrlIAmMVQlitFSO6xPhjZ7IIflA6wfQMsNU/AuT8TUSs33
nPujWM9NTraWaCTxaVkmZuBtQCTrW5z7m3NEhDKmcmnsblI7xT8sC+bciG1ONYLs
i+bRYzP/1swzO5GoSigRjQ3G6p07M7FMREAd5DuQ2VL4+XeAiVED2UV0SMHVo/Ua
7LNo5gVAMlDxF/zW3CCT/JualaIJfQSiuu+MwsgIyOfIAGuEn+5wQg03Y5C19G9H
cphfwkwtDf1X1r1BVU1LYYdUbGXI67lfIFFv7gGyE8G57VkuA4oGEBHCS7axVhW/
wxVexUf+czn3raHKSyDq7ypsO99BFfDPwhrdfMyilyBoUpC/kCWN54mjzmhfSy4F
gg1FvxqD0klofQHD84Cv4YUG/NtzKZvEwAemnFcLczeBzUMNABquag/Kuq0Xzv6L
/s2d7z2z6a+UA80eZnxe4iCVdo94jB4BtV8zZVq50vQLINgp49GMPOYKOHobtwfl
q9KQxha7G7C16HhC355kqYni2TOQsj9PX0HOEmmVOvIA3usjA2AakBXsIW866TSp
Pr0U3qPIzk18r0/Vm7GzX42wjE/Vi4CD4QHgPBbTTPSk2a2NdoUKsHTkiFoF4RzZ
2BQFoPRgXEY0XclJb7RzHEmBczXiXIHUXBdn/4p/qLZ6kbQRSbEeHZ8r3i7tYiq/
Xge8pAf8PoiLKbgZDz/J89I2ol6R3qSXRygRHWwzHDljCueFkhq5hse+zoyAoMxi
LLEuIsaWKNh0J9ajEodNtJQ6pBkQzCFOqhbeHpjm9m6jTK2plM5V800QOllLG1Ne
iBC4bU91K4uNA1h5J+LHgdCDMH8iypk80YgOy1hGTXPtBxLqYilujAr8ASgWRD6a
CpVXLobfvNvVBvhFaIzRpI4PTCer2u1HP0sZFB8rgtxmbDYWAAqw1iAVHRMAVaQI
Z2yYcu+hi/ZzR5LXLGwSS8yTr3SxZS3zfuylKR1PEwIWWSjsuLGKulaR3/AAFUN/
467xI8n28+GmDgKL1HyowaxQagYj9vcYYniObyd2d21R2LTr+Mt0qsMkgdOMnnI9
SJTmsTDgi4p+JyLSBmP5bYcEYcdNmZVM89OKi9ZEiRgsWXnTeYxSNSvnjCNbnCNo
bC8/blfC+7Kh22O1KguFGWMUYqo/oyHJDo8dkU8T3oRH+XwZuNQmcT5WrCDc/PvS
4bCiD43wdLkU+qkG2YOm6JwrMTRvKD7mvCRD++jUaaWHpa7mUi2U3QnySugg6/4M
k61M1+NHbpIArTF5S6dVoHkcny62+GtUM9y1yKTfr5nMBsCIcLBCnefzwlrPMPuB
dkJEBh/c5L9YCaXYfXO9zGgL05O9FwC2k08XR7N6JaqlKsxRFFsqTu7QyPkw/FQC
QQ+x9dgrq+YtQEPUaMEC0zaVqWZmVCLrKNXV3K+1iui9i7xPBEYyaEwWRts6/Zci
tmSBPUy+8pkGq9VzTbzZ/1iSaWx/i9UK9f2V0LE0QUQ12HdJjEAHBkWViJS7JiKZ
IMYQktPCzCR8x2ZOEBIqazZwBgZePXeHf/38S079O7C+OWWvm+rQ5vfRzWWWnoGC
VOpr9wAYB8/UhpQFo/vzgnG2iT78Pw36BDuBdsEdvZIE4ifEImX/hXNqmWBYEmvS
jHLh4rCozzAD10gCtkzYlml3XUuwMh127T5P1EpiONOgM+nGarc/w+mm+MFqW8e1
i9A9lUB/oQjbKyiB8GDMISfIqx/q68sfXEy7v7PmvHC94ZTmbGNyQoZ4uNlEvNoA
hriZf49rAoGeu8PoHSsKlOXfetyz4MBzE9AJtN9tfDS4i9fTtnIyy551tucqrY8a
sqDtEypMkN3nWRgCWV8WE0l6/IisbHG3aNrWOZDSAEplT1bzfy+uH2/pZXGYGkLs
kLC9/9whEg6WmRqR22Sjwo7kyaaAOJQ8+F0H3mMuUs97TdxoyeGshsnOVuRczI3O
e61YhAPuhhsjfinMFaYanQLxqkIKSzH2gs6FkwKHKUdvGNn6pAn2YSx2ROKCdzA1
AEkKx4ioiTScggB0gJ4doSYBq0b2mJNbQ5IUqDQBaf/gI0tL4rSKEakjvIT1U4yY
NiCsLh+iAQbGnP5BsP9tg/Nf0DezVbi/AIigVyAey8n9ODI/DBZOLlitUsP2Oj9g
FbnL299SKK5oXKjIbv7AwmC8VH3+814U53wAQIEb+aUhG4KqZJG4kCjuRnv/9SxO
BtHI/2ezG3tshanL78g6vy6sLEAr8deUtlyrysd1XDF8w0i+6zaPgV3v+0YcQXU+
+YHaLpRjIToyizxFjfcfYbcHZKxQpFCHktUG3y7iPwyh05cXG2PTgYAB4V/mwGj/
L6tttjCjweNIcYVna/atiMRVcyc499X1DWVvbk8vJgIYMgkKD6kSkQHpijPjz/rp
DX67b0nyGkdiQb3rGVgKF5RVM+LLnu07MeTgTdfWS7yf/wbx6NkwF40a3pLpHkE8
A89S/DpwHTkKvgScibadxPzCKgLjFeylB3kxf9xciI51q3EyzPWXndhYrlq5m6sj
WK2lRuC91xvTRei5RTGfwl96741M2eyHxsghgqUSpVIoEZBtynpZ3CH9iSteEguR
rVGX2gxjiVueV25iV1saNGu2zx6qFdgtEIcgnEAcxrheQRctaIRSxkNM5zGdqWvx
+9bcJ8rsbCCIvvGMLrl1ZPrHKFpiW/Bnqwt+rnk6YjD8IQ+usSf0abAVs+QbHr38
Jepi7IvhdKNRoC70KR50BRQ0wp8O0S64vwpYPmE2oSNtYTyLJx7v0kDTCAjRlLVe
Ds2GrXXC+mDWRMa7PHJClqO2wWrvLKKXLEjUdbRlzatvaThgZ8fAuJvG/JyOnrdt
+6+tH3L+z9q7OQkT+AjNbDR1kXDmL+JiwJP1iyc3zSGUQFDybJ7cZFGrT4xJemlN
dPLZ+L3QzAxAj7WRi8oBDVET+TRi6ybYM709FD+XFMQkMPJqyld1dovfQvYnUNNm
27VKKFNx/nkUeU35bOsdtttetOhDV5zhKECN9eb7RduPPwkje65pZphjJ8Z1veKr
dB/OiS3m+fZB4Tok5CA4vmRHf4lSJixWf0pwFBcZD7YVsobu6U4I9MPmfx5IxsgU
TuUg85PUpaBg5filPgioMWEmlCvU2RrzWwBQmL2Mcm/i1kVQuwgkE3tzc7ST/gdn
NWSwMSsZOemXsLD25QyfB6AXBPAcdbd8y3deBO5oS003xWOE9vn33ZaH1bG1nFwn
gtydt8O1gHgmH1g/hct8pu3vFZHM7MJhh8NSFYTd3tunfJ25A6H98WhX9Lg4kwpt
aW2rOAMYW6mG2wPf3gUJaJ0/JzBg3xsaW2foF7XcPVn7I6NKFjVujl6MacwFzwwo
luMwHJPP8ZuQj2jI6Jc3CZzj6g6Ylq6fIXfFwQ1NoOzqL2QXRoqR3yVtvh1OzuEb
FIFytAgXhSFMLd+EZFR0DcR8ziK52Nis5fgA8oGIuAIgQOf2t6pazMIGW+xIY4oQ
xabnrLzzbJ2a2XSXmWGMx1/Bil5vMTfq2OI4jKbZ3rRrsgBvRDYgdGkKHufGb7vE
Zi4j+pY21Y8eJ8Dk8RwdLMjLHlpDh6trXlLOhjfg9bvALn8qjK04IQxY+HCFzkmn
b3XpgtoQia+IlGcTpjav5hHJCFjbC/QmYCVQqY4hOVEKt57SJNxj8lB4k+IfTuc6
YetMl66bQWuH74D6Tp2V9lpUAChVLCLtqEb2p70DwD+hkgebLptI6t7iGAD2BQDi
QNt/4wW4KpkRfBtH/nzbR7OsGT1oU4Po/SRIx3mNya1aDQjvsdbB4zjYXerrPo0F
ulgKinVl8Y7/zJBhBu0v9UP3fYuafcFtMszx42yuV+rpVpEN1H8V9RWokOHULNzz
GV40DxqKBz+j3BSZ6RWaglukaghh95NgrpcI3g5PzcWZiYw9RzCVNSdDssjz9fsE
wJvziwyHq+EFTNLMlb71uJtXgzhFCdrZSZ5JgWiUwfRN0OOHML50KEtPhEVR0PHh
3kcX64RkR36ovpYp5GVrnFk8hTdkbLYKvpiC31qO8UJB2LZFdlnFZzP5sdNPYujj
d5uJBothcjzLPCwsKvHxxAtK/ZVxreAPVRRQo0//nA6UU1z6saje0rrt589kuQg2
PrkYDIPMWnsz38YMH2vGnot9ZwughfxoRZ800FRvBNUQoiBxSvzWtk+JTeS5lSNU
gRElOEv7lPb0XrxB2kvd5aOYekhtctJmtqZPpTgFqNecV9PIS1ytWzsn/wbmZpaF
LyfodVDQ9g6c9+r+sC7QnaFD9xq5vNxziy/gcVbct0uuM7rqmO32vED2yMqlCQ1c
EYDumxBvynT7yH6+qp+ifEFojQRTj2SMsIPvcWv54GdxDv0l/l5u7Y0z26NE8HNc
AoU2bYSF33klvLZL/a1mN/RBxCPoUB8CApz6zhj76/BMKWuZItgBdQV0OSC0VBpf
btCdfX+BSfz+AUpGNkXaEFTcr1r8RyIVtx5sIVZE6Qr0LiaHs7+Q/bxXGISaKTs+
p+29aqMjw79pf5ID2GgcU33CAqBdV2L2vCRSiJ3WrJ1CvpnCxaEEIkRKMQGID8/L
pABtYFSQdPEpI7XR6Gov8ax1+BfpyyWFeUxEAHx6SnfWdmh38cLTYLfWTfPD83/e
2fxqyO8SYAeedSu+Cw/QGEZSmJx+YaGBbk/p8ohZWQdgIR9lLMEypHZ2i6YgwwuG
kQ4ULmPdCI5yXGUa0kmUykL9XdOIGPLyV711Fcrxk+dMSbSchtZr/f9A3aZ92hvr
8AASGjFlIiYsX6QUZCXUvMLXiJatlgnEQJPkTU3LTIrtFDkZcdeWojAzOap+rQ56
0pmTq3TjJ4Aix/S8x4jAUFR22fKOc3VSnl7DVnoH4yqP9xnYLOps1LHfQjVlFpbk
DvzBGrNm+671eTHj5c+tPdiXnAsFCxqC3t/ZhazYHHgVjuV0iI4J8dqunluINDai
3LO+Sq+da9GP/VTQzXpH7Gr2FGUL/+80jv0C92dugKptMsAIq6aXGnqviwgTuA7N
uc2Nszo1fWNYkWQ2tyx/UXXrnFWzyehqgCea1xO8syIBgWjslT4QwDVeb15hUlH5
2AGrgZLHsCl8VjdL/6G4rchQ3C6OMNVJ0ghPLnEb6Ok/ZSdZvdUMpy+tm9G0DZlW
jCGttzxOhx2SJTFNTOCD+JDns3FotaaXi7p6AHHAjL/ZBavcpA233n4hg0L5mCeK
aRUXXaggRqEgob0IigOTkYamcXfNMnj8+8vFUEnLoEsXaaphfSX7XW1/ITYaxBN+
Z3/4SsJYf60N2ckup1iNZsHdZdkR4mrIQwgRImRUmE3AH18eHdreFaA5sO7AYSmW
KL1Ev/f7V/LdoizFVF77q9QcdwPShPVYiUZ9C5crXyN8EMbf/TVCKj4Oen3yXY12
X+N4s0xYCo04SUKPeQKfnAPO3IP02WUhsHsijMbR/3VZx9K4SeN/EX6hprcQmSNP
vV+kwvZA+s/9I5XEGePbgEVxPG3W9mlw2PiyBGwVx2oDuDZzDjiK+dgTp1KS+mXO
4cmw0mf9ylvoFrMqduDK+hKba0VDFafbmD6UdPRBY3Gt4x68hA7ohSFLBKwpSkgc
kPm0Kjyf8PejCEIKSfEE1DYW4Meu2eeha4dJx1P6EDFav6ceG4Zo1KLjrUUWUhXm
ezKElGO7thfd4HlYqN7xO89Lb/2nHmQLN/qMPFZY6GlV+jouPEjDAGDVmWolVkJn
AF4aUcYTJ9SPDLS3M1SDd12oZi2zo0MWg4f7Sp6Tcno/7Z5dfLopDPsO3S/d7P7m
dmEgrTEtm8dUBSJn/LMxM2bHERmgqZvR967U6f0nMkiD0SKTg2bMmnGo+HijkYTh
51eVer3QLfeLuKOCs0rEscoMCox+EiPtHNUENwgW+TymgdNGjM8SQx5Oo32hIxYG
sqiRA+fm8Hk9/Ub4iPvNQVsf+ElJtyaKfChx2dch97Z95qybGTHwJ8PFw/CET3QN
ivkj/tx1Dw6cmA8/s7BWIYCgw421sTluSiF+I7NGypTj3knxZ75JSbgcYUcGazZO
U4zJe7qUIa8eHIPY8tkMXfmhe5SzdSKQ2e0zkg0Yiopa6Ir7KQs600rrIUDypcTk
vtQQzcnb52a3Bbe5RcBDzLHoH8M22V+zugmCwQalaY7bepUAtYGPbYQfF4SDs8Xy
Q+g56z+fUJWuMshmDWBZCGtDY7vFl6BJHjSufyEblUZvEz1qZFE3DS3tuHbThJPu
1etE7z+iFB/lFlmpocFoF/uTftllcAncc1IcyqX2AdHKeQAgQWMHmIwhvvONIsKs
o4iuC3rfSc6sdSlOXXaOtp1iY8iL+mILlxjIh7SvPxviSLJyL+N3wp/HZcquDDDd
8C0emF8d33zMAM1ok2fMLoKD2j9d36GjpbHYWiHBpoA5wZ05wybVvZoA3Cwcj3IW
kUxDx7yVvv7B9TfzupP+x4DQoJuoelay5UU+94d2x2LNftpAC4X9CwpUKKQWrpFq
g1dZ4kD3LZsSNcOz8HpO1XTQFzx/1CfwtA8kQ8CMfeCSipOF18QCXHsvbRs6VMLa
pvKG+n+Gns8AvCfC4YQy5aB65Za2/xr7yd8cQ+DqOISoRjLgsAa028A93+p1NkWF
SwxXXwkLHS4R/WH75TP2jPREQ565cdlS6y9OuiVyg9coB5ULDx1jrEnmNonO+ocn
qPRimeRcMSjU9D0REK5VC7Un3BsQvOsDTfbcwHRClpS1Qqvo6dZmoxzvwo0zsyj8
Rx3tFXuYW+xk2Gt26HeYpOxg7zgbm1I0opefXk1heXOwwWQtQNJE1mEXkBEpD8s4
8HzO9VnjkITX1iJEGQs+yzmlG4+qOrM9t2fZbp/gYY09gYtZkFetJQFXoyrSscqJ
dIlyScRCcXokdV7evNf2U1SBfSg3Q7a/4xIGYRA2imVK427sAofE9WUJZITktI7p
91U589H2ZeEoRvbSD8EpGqHeE8QppyMCT5OZxfwdcSHt0sYID8QF0PzBIcH3eY8q
MbGrr+af4tdgDKOfM516ShreN0WLLHr3IkbNXiUbrvQ6XJvM67pg4Lm8Ow2qH3Gc
j81f/qcksXfeZnlaOcpcqgCQ1fPpMj3mwLHhkZsvQK3FXWkgrjE3v35daysjVYie
Y6jqadu79t5QAL15hIMxM1r08dLnH7A8CiKD4b+POcqm7E571umVkdfV1NTPKI7p
O7+tD+93ZddnD7Hf3UmXYvjaQFsm3l16IxwJBKu1SpTGzk3WGgBlNd6AEwEBYVcA
aJylq+zU+JDn/Q+kyw3b7miffHdnumSKO/4rIFvGyPUPlUjs3xgpbkni6EvNF4+V
Mngwo+LVQiH1Xqs9Z1SFNYgyu478mgaXTrCJkrhbNHLt7GTfjhE7vuphNDNcbkzB
g0PEr5zbwSGvXSAsSZrXKpQpzQO8POTFuwVj2q/ksnRhzbY7L3iv1RRG7BSuQUx2
OWDQk7zDMY2cQ/kClH/cjSFGrTnuGRSxglydpatBUL8N+H9LLeUG66n7IRfOKlUA
wvMQhnsXPMKoJEHu9ml/XjFBj3qx/d62fuJTxZAGSvZS2nC/18J1of7JibEkL11Y
nDnnGb7s+v12V8zUpDn1XvGImOoxbSVEaHSEoN01HQ+I+gsyH9FOktLQeWUCk0Ko
y/rNHLZTwUCgvIt3wGJ5BwNdQohjUJFWT3WPSs5DINy+lhzLPOwhehVrul2YD21s
gZOya8Qw37ekc+vDajoZDL/IkMKXnO5DcPlCQ5ccflR9indDpaRKkAaOrcZv7xOJ
j/xdOjXicE1s0V4sxQGFhMENhzezsT3Soa0pPWe+1cEElIuWZJbDnNp6sMz6f4j0
/3y7EcbD4fioKAnjEiEejGuWhDFmi+E1Vne9/EHoYfyyk1U7u1YduTGoMyVuiwyU
9HwBecD3qNnG19JiQRl09TZQfLwcQVNrdKPS5ObqF25OKGRatt5jlqkyGs5PcGUE
0NhK7trBQ1jRyjYQsvsueUEI719c+4lvzeiUHpJwu2kyZaoFFFkR5RK0X1VK4T5O
ClwZhfxMgsbMAvCJf39jizhZkQigXgAR8dfdZStLsRBFfa7FEGGAdFYlZ5143e3Q
ndLK4xmDlm17Nk3yVcYutPpRpQqosXQ6EVnBJbmpq2Pgg3j80ZKvwSfDL3xJUq4x
7J9sYljTNizCX/AjzS2iPccMGrqNZ2U/u3OOdusEq9hfkAX72muAhwArKs8DDkSA
QPyjPGcXraGkKf9bCMAgObfuMkQs8ZB5JpPVozNT9n4Nszd7OFyCO+Rs1KcmH3Lx
vA9xZthlWp3eDnDufWETZVkIq057nKlu/5qKKOzrWTGdHiCa8WMFOuF1fYbjCQKq
IIdIm2QQ5oK3r7f4EJ4A52HCSl83Nrq5u8eADwQkH4F8i/WtVRR7jaAhH4xfDuCs
ejx7VK6zXIz/jUHstjBu/j4MqM11fFN1CTzMMugZ7UOD+3Thcif56Mjhk1bbmuiX
6I2CrMuL7QfXwNkW2cl64gxmZb/eiKqGA4uG8ufT9vsV9JnRnvk4aHkPF4yFgFu4
JPo5nYgEg5dPIOVhK9TdRKkncIKoFmOSbKcXF8TZqlumAhM2JGhFLRVLeKMwE5F/
wTQwWFK5F5R6vUWmegrAkBcFketTfcTCj6PiPa7h7J36yCDh0FKRRl9fVUuVx2SL
XUAuVO0O07duF6lS1///csiy66oU0AvdPW/iiEt3os80P8wc9K4cm3UvymZXvtWO
YA5zC9rFULqRkVqQwqG8QORplj3BIdB3Ehcb+VvPtsRBZ85hrj/bFJ9qTybkiUyg
XFekXpP1qCwpwZ/mMg0UXbUgXr4Z95a4GoVkx/M9CgRWrkNyB+9/w2+2QNn2S76J
HvvntkZMd/pho5zjLD19z70uxshuAlNBrzuSDlOwQ4bBMLw3bGwxe+XgamZBBz8U
hvKMxX2lIKapGL5ChGfsMZAP+UYHR+ugQSJ6CJ9Fu6WUpMziBh6xgVGdfy3GeZpQ
TOj+5blUupaLvZSIeOooriqOM1c2y8H3I0KIEtFD2veiIKFU18ByOuSATzC9viif
3oQ/L6XscMzssxIp6PIls3VJ8a5iZQIjXNjzZgCitiOISbpTKaXo7H4ePtNDZ+zU
H609N+Q8GzUQQ1OAZ/OLP07XhQe6mPsaLeKfwtB1H+OtW8IpSKlafgzSBCpLJ0Gw
qdmETXw0IkFJisvU40eqXG2k4cERn/+OcbKBE6S2DLd0MR8FFONQboQZp8Z0/UiI
/OCat7cHDg11HKpZV8DxeB4V3jSl7KT5mJSESkZEIbOtE7kyRYyiepj7C9dq7B5n
pi9153vogx8WCrALKgfexa/hFUZker3l7NON77Viiz5S/khT+9oSZf/2MxZD0GST
qiIzJQDf65ThXwBncFsGidrePlrJ0Am7zjtj4AEU19LaKndJdTwH7yuAWXPGN0M6
89CTKbSL4oSB3JJqrnjvzR4lTvnzhQWCJPdjXfayvkRi7kznTMotz0t/W7udeJjA
m6+L62cyB4cK6k10Wkl6ECc6qAhumDFB//HSmklrKq5JVQm3i/RLpVo8qW4E6v59
ZN6Atf0V+Frn3VnJRUSwVC1U29XHqSjz5pBfE6pEr1WUzd1INY47GQvHlU5uHkFh
kdhtg8oBbUj8jZkYSV81dHc9dI2l9JKxTLL5bFBlv0ljHMmiIoQJXTQOehfJB6ji
PAI8Yh6cximkQTEjgHdvX7gHu5u2e4efphgmqwWsnmJd9CHnrLCBg5TUmwsodzdw
GF5weRUM5xv7f0jhLQIVaN3wYg7P6ZrCSXMBhyWwDAdvz4kFVvy47k82CisLgGa4
zv+dWGtir+QtHM5poQxpOztUvCJn3mlTLfV+YUj3D9lzd9LW6/JsfcJG7xbDpjiu
6pGRmw1PsL0udZ7u+zSpxj2OTNqdt1S5FeA0DUjFpLAve2HqqrTrLtpV3kG9idC/
4J5boQHak8vrM7MlyGn0a+98/M9lAO3ki9IQ+vzFUTfTGuhNvEdEjO6xNreu++Jr
Hmi4OvjgureMXbDEpDeCHC+GagYNdc+r7Hl/p5OR9dSFCHQGiSMW3XmFF1P/kxaG
wI1mHQz9Mdq+5tvd5fZrz66S1VPRiQOPpCqoq6rr6LhlUsfEcHgrJMj+Fg/ir5bi
+KhsdJGfl7IwnALHBR14zntr6xJOMqrl/IMlhAkUsKUdDqJaoyRedYVh5MVAAxQR
SrZk9L178XvQMtpt0rR+LHISMcINXsc2InBF7r+yOAwrCJOC82HF65eG4FMq7SsN
7TbNCJP6gs5KGZP4fOwbL8GcmpChvN6LLmQnvxNCG4w5QVIstruLAfDcGu8+Ldnb
zhXvjdIlpsD0g0InjUBcnbLKI/S2gwGHFtCUz9wuFNNaChbK+DVh+f28CM7TzUv2
ZNppZFQuBCkX5QjyrvPPkXsVZYDeywu4F3+o8Sn30jhm3LXtWkk55kLFSOa3cB8w
4OypXcycAdjudsn/R8pgKijYrZBz/KhktlbkGwlRVAzsAMeSEQrXYcKl+d+Afsrn
hBUQcL5PdCrIIIDoYOgdg1xOtWxVJyrambQ68K6qitPyg+bbqXeRrhU+e4zrFTJj
Fb5dyXy7L2qHwfsbkTeUm3xm8bBnBdi6P60mYuNosiJDOxPBIkyrGQ8nFolYuu3I
KTF1AATDrOTmCTZJYobQQ7l4xiVEaLmmWzR9+rtOTxz4wkn1F326FnekhWWyPDn/
FsH6D/SgYM3Oo8JHiwkxOuyHMs0xf1dRGj7XRu6GeB1pUL9DhqPDKJvo/zjZi/Ub
2G4aa1B5sbUsjV/x2ZB/AlsNCv6b0evUKQ6rMf3bQSvjp9Zb7SIgHy6XKPJDk/XD
904CW0t420OvAj1qLPQ9+4XQvnSaw+t0yTVmcxbgTK3zfXvl9ARhtXMLYapPkWEW
meZ8q+29swRsoZAJ94JR6bic6s/JKhTSSrBvczVwtsdXFXnGfrrhxDB97vsW7DdY
Cf47P6q62q4CmlvTXpGpCnI28GLzPvGB1P0KOeSqrjJgHpBxPI/5xsQWKO3wFoLm
COj/ScULTvGoWBfdjc1bpzvSl6bPZXnPFzAlCX/gMchakq6CAaEYskB5D9BsLq9Q
IqDcLyHi0rNVwbFwtQGq4Y8fkzBOGp7ibmk9NJ6vC96M/v7NNQe98KK7BQSCkcY8
v2w9Wtg0JtDGetxSmqGC6aIDkBdbfITv63jAfNBkccMnnExDCgG+oNR+H938BZPY
P7/pI6Sfv+25Ezac+3DVaBm6y1AEt2YzhfTn95pUENDp2ob1R58dOQxDMauquFNY
KvDjxK/np9iAqqkpNB8qFM26NpGKTAfZS6/0Ajd28koju1f7SoS1N/zlByue8ZOC
Yh9Q6pjgtRjIwQr0SRIte9CBIE8seN+wIGjRkZ38XA56YCa1cPQptO+XhSADvStZ
w6loG5XouADmLiYRYyCepbYfxYexdqL4u9M3a/0ez3hv3J5puVqmy8gkoq8M+r0a
jPZI4OwqHAW5OY2lJZOKIV0HTUP/4Y2ut76uRA8AcOyeGhcod6guNqxFAhkJAT3R
yTlIMchBk9LmbQRaYLf4zS247NGio6m481Qd2jPJ5pNkIjU0bzPhzTmbOVrjWqwl
G1N9AmePBBRuAJWviNvA4dU0l1cWy3ccZmTteO88xBFSX4oG6Sraaf9OOxTL6X2q
8v/Wy5TZYud2AYY1i8MejxjI4XGiy/QpTCV/1a6orfZSB+fbp/OEU5A5FFzdQ/5H
WeKHpeeiSQGPN6Y/YiJnIMjtM2eiVPjJpIg5pJxBoEpWxHREXi5DUYX9ay1Iw6uZ
97CPQxjnHfLM5ui5e37r25Ko+qKtrPlzsC1sqY5eouqW3p0Oi/cgkZ7esb10qegW
yirWCtCgGvFQJ65V9hOFcqHvKKEOLYS5N/CfQJQJQ3OaQiZA0Cr8yui5Do24NyAz
Y6q+CjcANXVtpdTKxitbLboj5vltkzwRKx2PA/4USzYKTnfgPRwMGMMDfHwu02l4
6g67aBL5u91LpTxnYJxDMM1MN7NW5Ng6UVvw+HwqMsDxsu7khg8bXDmK1fD556NL
s1ZKacoXswU6ckoGvvV469JQfbtAIax39Q+MCroTg5YssvL3GLZay/RX66nV/uXi
Ne+DIR3CE+WIMEhuBlJhR9Ct8o/Nv7eCXonyvBGG/Ejm96X9JGARaMHAh4LaZWhW
vpqH4ofhGOFEDaIxXJlDy3scF88rBvsLXolpbQY3nRYOIKy94BmR6TbemCwTrj7V
vtcfIeB/7uk/Ow3Qw6uqr3pAoO3/TDchTSV1AHtOwcg9JReiSQk1FjoJLvMlnKDA
K17u8qxI//9OWcQaFXaXeycWTPQ7P/U5Aq5Gi3U2dST6UFJajvVFG7/IxbdcOhOy
059DfgjCce0Es9vzLOR4mzF+wsu6YtpxI+Dc7t4xV5QWkskNGl5LbgrUtVAZg++o
j4b1YMoAml3XTL+g0en17Y3c9zAKWbX92lFlZlcJzc3fiwymAVRawyp11Xlz5tPk
N6iFOmI+FKvdOS80EMhzk5OBhBEeokJMYO5ajyh+HQZ7vIBTRPB1fzgo6g3wbHOX
DzmjYmIWZGHWVxGusAbMs0gVAwWxDyoRSVgbVrMHuBnqczQs30Pe1VDJ3Xp93EFP
TWo0LVkRG/J8h8YDQsxTL5oFCmxFu4efDC2fZs+jRpkWQ5ajfZprYahr05KytGBP
Pn9cdPfEzUq/8UQBxaTPteiFhXz5qEumX+6zs0/jd0OVhTdsnR7YFFIaP2l+PgeP
W7/HDwDGaN4B5Xjz8lvq/Nw5IhdogmzfzwmhCQoGF8HPRQOatDlMaq6PPDfgIlPy
0xQNnrhJExgH92t+y1JlbZqE6o+h5aTGyMWCswIQtN+X/jX4bhr+eJ/IpQ62eIQw
+4Ey6ebEzebiFmGpUSlnGqqKxKGqTiFLV7mi3ilmdVJj7Dv8Ycb8In5p/4kmmXM+
uMRVBcWglXeU2FrQE3EPCopw9r/FeomdbQLqksaLf/t57ScRy2HDBNjLv+PVFxJD
6RU32F2xMhaET47jLtmzLcT27KepYf6djxsyjWJo909X1QsKrnR4Ze4lNh9+8xJC
lrKox5pPHVELz8fPnw+xKtqXvTur8bEr96gzqIdyhVKrJrqTQNh5B45CsyuKvs5b
zW+8LjTlf0lgGutF8sGC5HWvhL1rXzH5Nd7fz9yhFeehkWGxIqxLwUlRQ9K+XjQO
wqWoPwHQSutY/L7gOhGoRbZClHEdSzOWOlEMlgCwxRgic6b9NWdDfH+xsChZDmrJ
LzNd3h0/eRBOTUhRuz86H9OyjL8ZlpyaI9Wk33qbVqGfT8yO2C0knWNOVWy2zMAo
DqQFJ3fsoBvRdTmtLd/AEdTpP0zLG1aP1TxJ7ZlG6QQkecZaN9xroRbHT6sYtwPp
LZvuDmCQJt4IYb45ymxRyqF3QwcfHnJOB9YTAo+V1ZQj84ACeL4q4ER40QBBWxVU
IcDtiDMiNA0OTkr8GCQ75m2i2UrMNaFsMGXbtY20x9yZvTB/BxmQE4rJCbKiN1NV
U/dGjo5u+vBmSekB5JbJCF9hO1Qj8BC2cvVuoLa+W+lVLIgMVEqnbVpqfpkFkzAp
fUZhGxjRn8Jaw8wwvODgBiSLornxkUI0aJ9/cToNpmWCg0D3bRgDxBZHVGGX+30l
uXqrbDjVsXzWov7HZLqdUEJVcijQJyOca9GxZpWQxWQtl+eQVQf+DuQaUXfQIYVl
Nb5n2PGaU5GQKwVolbrmAIW6x00Tf6PIEM2AU+ZM7iD6y4jbJjRAe17IkZhBlBQ7
zoWpfOdHoS0vdJG2gBl4mlrrA8+dgAH12PwxlMxBsng5vvnYaGRtJVFCQjwpkDl9
SlEcRWA/uOuhbrDWLct97k2slpy3FBl7UjTVNNBA2bD0g5y8GdP0ahheHxrNAAct
8IkhA+Yrr5Emwt20uEnh7aU/m+6qb9SCM4D4O/5fs2oLMDfZPf5Y7LfL3OTfnxiS
5AdB96I1JtAOV2ERGeCNlHyxcPon+9zSqhFUWSpwnfAK/I1rESiOQjTR75di5aw/
Qrg9TqgUMrUpg8IiywnejR8wdc5LBCrTzNbJLMu3bOD8ecI4/6rGboXFPvNBpNmg
1/qAkKC00eL2sV9dwlvGnin8XbD0t/f2OYe+QmeNF4/kaZ4jlJpZhNvy2iZFgqud
Lnz2BPkAdSJe7LchUkCXE84JHqUy3UTz24fZtrWE9lijTpcZGlUgbS/lYqaxLOVG
YfYNVX2VKbwVkQ6IljU175xxg5DH7/E2knC8CPjX0mMAFpDjzk4R7fPGZctT6p7D
ErO+F1YhbEN8pWR/j20OrmJ23Wl1RXTaQ+aCZ7PLN8NjEQqjGVNd6HKOOJQEhlT9
M4/06f8yzld3evRdtE41g4wI5u7oBQlrN+p3H1i+zHRwD9W+nkqL22n5onQJCyTm
K7jZp4JLe6VuRA6GGkszblw8dQSPzeZBXy4+OSGkhgclXv8B2DollRizgSgouhFo
SExq9ItIUYkzPb41SLDy2h+pafKBgsNL6oKLDMfEVSQtVSgGrtQIB62Eu8q5ODjZ
fNHHijyjLjBwSTRIpl6Wd0W0tuX0RjYJicLw27o7jPufMu+4UZFLSCiVFLpVT4hY
8awClSGHar5gJUyX7rtnVEEAaYjLbafCxyb5dYhQKgGs4hsagCfWBzr4EIUpmokL
FVdLqBLZAjVQLY0RgGr1se/yJsOS6NtvTh8chewY18wSpKQKQ0jVjRNuhKjRSX79
1ex18VyXJi0/CAiz+hXBsCHuuM4qAvdAgyGMm84Kb+R457GXJBMFB0sqo8nf1ncl
p552ZrCeozdtPzFwc9ov+Uvu6SfpLbdBc+W7uXMtdSR357LLTAV75oJxFsJl13Za
rpga17EQu4BS0156nH3GDG6E9FG+bUXtYcqNAVgt7QRIMHj+m1OHQyU/JSHkkFXR
Ui5JdaN0wFr6zzKfXE7LSJ3befJDn6FXZuK6X4mzmr9B4ncTYF7KFepdLCTkOCox
zNpDI8IMK2ev29r6OFosltH1bIG9vNti8NU+3HYH+ki6itrSQPtCfd0X6TIq5KL2
phONq0Kil5RwrYRKVzy+ZMhaJjUZdDA65jjelPLkpPVzDPNonnk4yxM6FBNea3YA
13VPKKXge7GbrmwmJy/5Wc/2jG/ZeCrrz7iJrwp1/O/DNxuSGMDxYffQ83aRqPK3
RZSNwsYxZViFOx9E8jtOq3SvaVtpWA/7ntLvoTDG/k0W7o+VbPoY2tgbmqG1FOUS
iMfxf8BVzf6xG6lgTHVUWsAc5HRRjAahY9ao+0ZkQYjJwxV7n0ptdMlSEjjJoA03
+xoEF6hEkBdHI6IyUUoNi+NljVrDGCSN+fPgNTmRN0WyC9C7IT8rflpdQWWsKfjh
QWkkqwsPbkp5M64ZL7V0Ff5SEgC6eQyIsV+iOlrgCbHWq2BjEjD6MfZ7TzrsVi72
Qo5jmoiCuiimvtJWB7iy//v0pm15QRN2cF63QtT+AmibKulQAhEJeQlBlfrO0f0J
xK7EKaYzgOFsOGka+6gRwFxEJyryn4I7ykPhEufGfS+MOQKxGDRa+jb65C1NxBEM
+jSX1zIe1eevqtdshCq6obRhgDsgHgvC78vGxIudwch1V8Tw5FsqL6e4m5H9C/0i
NVrbE6FXi/VXZOZSnl7Dzlxbefmasa12hlaRbHK5oWCMEwJHO9tNpVprcx2DKhlD
OisCAtMhSKyrn8t9pVdIhsN74/vBqaBpAviUr/MFohCUOx6pV3bG3QSA5O3fQGRT
R9VHPbEmUiFl8/rM32bgShKpcYJl+apWG1zDb08X9VzVaJEfdKlParRCiy+4r9m2
IA8lxCbK/n1iy6Do41r7V0mEWpX4HZwbWsKX3n4kDZh91bFpTXgA/gBbq/sxm7d+
gXVSqsHTy0ijyhpjLlith7mpCk3KLAL7oacc+mQswuVkZjlmzvf7iQa3x8sMBHDW
jWCWWmTwkc0KlPc/N0r+ybRCFSqTLkUEiMKbndhsvCQ1mB5kLfxoniMtWauzv7oj
m4kZgCi8BmyCGNz+XEV+fBi0uphz+N0Z6cUnDc0aVsLcug72cd6MlVYLW+RR/xjq
JO38PDJ7OXMCgB+FVaEj3wT5yBzJ7oPdI5yNHl5NHCoo01ZZXM9XCKYpZzoonq6a
8h+WSqCLccl+5dudURTeiaFM8ygJ775IgZCoeyM885WkB6lOpwXRWy06HWO61YE4
tsNW7oP3UOpwfKf7+Zor2CuLk3kHRD8Ek9tSkM7qVbNctyvjGtqnSOZiSo+2hC3w
g/V+MmVP0X71//jHxRl50k6B1/NqufUrBUQKOyhdIU56Df5SpTN/SGN89YB7ixZ1
1fBnSszyY41HXnOfnsS3guS4wdS+2K26uo3v3IN1dVewgOKBqm3iVvA80ELdlktc
5F+WnSClc9xs27t4xAcfzaMjFU0tCdvO1Ln6d+SovpJlaSNxc3lrJcd42VolMy6b
hbEZ8p0aPBkefApez0STv/gqf6pXWmKcgUtmNb5ppPcX/8OhAFKywza/99TBEpiN
cfOTB3mbMfjPeQvWvriDs1C7VdlOxQx0wUMzmeFkC42yWwDqnt98vQNtgDaviXDS
5hylnirT/N2aBJi7UYqbAzeE6mq5L+sqPutKQmE6qKKLq7VFuwT3AzqDiu8USVj0
MCS8Q/6Yk+1fjq3IYMYk41vpmLyYxvI5VJmdg1LoOb23SQUOGcfuhnKKQNeis8Lv
yKVr5wSXcY/GLKTJjg8tURdoaZCzONWdXzfZwJJu2y1xGczY50eHlr2v//LFqguj
BySfXKnOtS1BwNYIsa50EZtapCejKTRyldOnSs1tMYl5DSjtQ/eSgUW833u7gOvH
T2h8wW1MSHL2jx6RFQrggzKrvqf/SOGb9cbrbgEZW1rr1kMg7IzEw6ST8d+YZi3p
oJDv7a5mpa451r/M9o8CLU2x0iPFkY5Lec9y48XcdNPzd0xk4ZuYvpx+Tvjyw1R4
7jTufWVnQAAxf5diff2VV+es1zgA0jCbW4e4ZfYxJFkE1+Sc6WSLRxP5kKX9ni5S
uJw4V5Mi8Vh0FibCa92Hdjb0yDCiL9Utjvhvh7uJgNbazt7yh+EpPsVUskba3xSL
fFtFyIOIMo3NlaBLyU+gUzNZmwjerSXG80vJ9xRqLfh6g2YjTwixB5Vyi/8adPrJ
AJT124nmzn5uUk9C0vJV7tLaM2HRdjYLmtG4LUo9Pw/FYQmaXVBeVmozczwNEVJ9
ohJ2G644xshk94c8z/9tcjvlacRG9N8xbTBZjAwLOMW3OgsUPNWjTF+7IRLwu/6K
U+uaIMVPH7sccNh50h+y3m+GXY+PTrZD7TMoFK4VyfHsTDmcu+H/k691AAeK1mSC
Yx+KozDju4IeJEUOiGfI1nq5Tnf4jSdMP96o97MLy2UfD/lfwjmPuSLE4ykJNRgw
DtaHIAEDYVenEDZD3YpXdRYVTS/TypdWgt4RYFWWMkclqyrbf3PhMex0ucIyvHPT
tEilD+3FsGi4mCLMtJ3a+/ElpHv3L2OtLr8WOw8MVbcV7XLmUrbGWnYL0e4abka3
Z6rOOfrgp0nLahjn0ybXxQnRWO1WJf5AotCT/4V92fBjmjUbVQplAW6ekvu73O09
QNH7JD1ko1/I/cL1Hn1Tt1JD+BuXPmkCZ5HSECMbVxQu+auJFLECymIIt4wQt5ZH
fbvhW/sm7z27wcZucr+qGWTwOjqYtBFZIZF806nQPPFRLix5BHyRV5E7opwXZtmk
R7pzT/JgYB/oDVw9CU4uQFOFRIyJ3DGJJ+XIfT+fjyPq64kqaaXMrqDN0L0bz1hQ
87UMZesyJEjkDslPLw0Zz6OslUCoieKGYIAdJCyikuZAR70oZ8UDFbUOyNeh8uBz
AuLL7w5QOYofmH14hOSVG6YU+elZ6eMjoUPHXaQbx/GK3m+26TuvZLX0v0m08WNB
78gKSoZBz9tNsDpptgr3W+7wyEcdhgFHz7zBlyjHSR56Bhp6KhXehViPD8YdP4Df
91fFiZr/qAyAoGEtd3+4zRd/fzWwNo4nhCNB/+8v1GAl5ULSjG5O8YeUKj7bh96h
ACUQ4w+UKLuKjciiLBWsNk0sNegrllPlTf+RA8HUQZDGiGHwI5yfGmgz6+Rc/fw0
5lBJ8QwIon7w/vdOBa+8KTbZnswG7MqvPVaFKkaCT1SHwCDI/IfFVsBUyTHGj9ot
Q0e8/OWUmH9/UzjDVki9dY/8xt8+BhWzUP4L+yQuAWMnyYQJGjUenoGALhxCTHvz
sWPVJeTL3tbNoZzKyoEMUOjYn4Dr3dgK00y35vtfzR3vQf5QmXxOmO4MAwm/zOgl
bMoeVA9CHD9qfSVY4fXCT6f8V6jrO8KdKsM0NBg6uLR4N1J7DvaqoTI6BwGMLyyo
0qnYtatJunBHMUcyP2TpaP2IzCejdCh4kPGHRX7tBqjrn5qlN2A9OdFAL1uTW78E
BhujaAvIw2bWK+d2W7F4J37HUOQ8ptgObzc6kA5c4SBEKtH/ksFJzKv37KyvF41W
LE5nwcC2bRWFta7SYzjJ4yyQ7VULgPmcLrJAzZffAiElJCNgQOcOmYr0JvZj4Ehq
IEj/Cd51Sk5lhA4tUuzw5MgnkvjJqZXIJUeu8DDctHLy1fuH5mXcMfyp8grIe87S
ObwrVMTP08UqV9e0RvtLIS+SjYTbngca4o8IGAJeKd+U67/c7tTTCBwXDQA05EFK
c1rLSysBKiGKarAJHbfG23L1U91kzSy+F0o93TNGxDXqW4R927mFX3KBRdx8PZBC
bXlEl9a69IkYySzKBCixPiK6wTOoBy68H89fBSD0xo7lL2YJ+4IfWNlEd5q+LFlo
fWG6VY/IWTmzWsLET4x4TMPq8lsgESZ1KOWi2r98eRnMBCm41O7QyBhSfkcamlt6
eTLx/q4tK6QHSEQCY3cJr4WmFmU6wtLuwQ7SavpNdl+sN3juZPH+wnYQoC2Cn1/L
juJ1wTwVOoAYWVjKmrcPrRcxUrdv8VsVOzE7cfr5jcUR5wo7pSGAFYX5FSsOpSpG
+vou7KkY/Q3RqDOVPg8A0bSReaTfGWc3FOXF11xbBkCJrtBSda/AK3N+pPZ50vXv
XAwAa1dje3LtgIYVO/SRwMtcG9FH0gCb7dErGB3JDw+oYavE9oErlSgGQ7lNDn7V
Uo7qRxuT6eB9lvJ6LSmRI3DSreDRrQ+gf4f7QmQu0tMshcWvm3fdCJssgbsoifA0
uxD8DlMOj/+ssB+Mb3hDAwLv0kJblySHIY+mtBJw5/bl0tqOWo+MKSM1RWIghgBY
Wli/mlb6Bf4EAeo2zBpFzF5yGtraovff5d+V5h6cbgDktUoQPsYq3d1zVOdWVWtB
YGOBDreBrct3B+uYzTKTOLu7OQGeoEfv/EQj25WLy98JbV+e/s5a6uWML4u0BeIf
Qma+YmnvaM0MTDp1AlbBkiFq3hwCGG6Nx9iRAABMpVj3DBuXlGz3epewmYVYiJr2
WOGOgkP8MBsSpwoRPDoUrR5OEwM6LkZEkUqWoPbPmZKcdLmHbgc08p7brdfrECq2
WIhjw/K2W8PpIzBAy9jKmeauD51SC24qnOp/bAnbtiLmjELGFGLLxuI48eMmnCuc
yr3hCt2dbERXyVO7zKc634IYAPfUekgHg1b71M9wNcS0qX/G7o01KRtSJsyioS2e
jtsIB9cNC57cFtSATGXf1pEzHr+NpJ6eaXLfKGiiezaTXdE5MDdgisRVh7idskBp
l+QNQlTFIBz5UXM96NwOYArVTSMd7ltwMeeIjR+4PfKZsvA1JVMqVr9wfrnW3ZpI
YG8ta2LCs1mdewsgY2hqzHonOugKX1IrzNpw4JP64HgRAYD5bCshwvT6n5MLsXkR
1OFnS/X2LcgqPgiB2trWydv558+k3cLF8twG/MuhCrk+LEkKZqt4p+kfYeHHecox
gcPQDZ+1r8QYF2DGZ2bPsiXcIbp8wVG3ZFp++dXQXSivbhDlKIpdVCa+DwfqADrw
eN5VN+Muxnh50K3D1vWmzc0E8OW2hWt3XJyh5rj60yB8oli7i+k8DCvOPg7P1lAo
n4x0pZygWrxQbMXdOVpKyIFAemwFnCaSEzIUpNOf0F2l7p6e16zfLg1H2k+YJ2W3
ESpLynDgvbi7sBKJ90ttlc9W+1Qn2UHej5nAPuOt5W0u+t4PHuFyYbVnlOSTsXl/
5wxHO7rCX4H847CETt1uSvB1z/8hs/8zJDtZcU1/p153eWS1Gat8n81ZpyukkFFu
CUZ54Yk2ffbd+Spx8j98fnfL1RacJwn4YTcz3Bpwkn+sR7e8hyRLQDyO3OZJ+/PT
gRQ4a9nVwJsPhR6H9YKuv2qhHbqWl5H35p3muPQjsrqpAFHHHKkx3kVAQD4Ad/Wp
oSwoY1klaPUmz8uYkoAGd6USff3GVAMBeOqhJ/icb6+1mxDMSN4bHBfMjAs85erE
DA2mXrjlQLWeehZV6R+GLDn8R226DZQl3xjTwuPJCrd/B8HXN0bSkTFhPBKCMm/B
C9T6RFVJ5FB5RTS44GoiFJ/R2yhqMYBYWnvS7ZxD8Pw4kLVeVy7npBB12lZ5G2zL
zQ6AYA1uCXbBeTMqBtmyIeAmXrW1SP/NM4eZ/ARzsNWo1SM3MpVo1zfmEHUjinaR
cn9iJVpHPC5GcPT2NS34dlP1bBIcwmr7Y19uMWVWnba2N/V34mjBd5+HX1wgBpoo
Uiesxet/e9XQTn+uMXeabizOjDU+4uf/m9sMr1EpUi6Fi35N/0HpP7uG7qpAWjYk
951+0w/jIaxpdXDBA/v3yDI3S0Oa/Y+q4tfxJcSSNl5x52X/j6jWlbW+QAc00sKn
QByaAdpdp3o8rMjMZgf18YVENmmC67sXOdDKZ1QjWciOI88s4dXpohP2BSE70MiQ
vZJwSo37e/AqmEqXvYpwh5lTI802DvSf8jOVG7kd+LvZRGA3mOyMhLE3kL690hTn
vxzaHT/8CiyyuUlBaMGUymWJ8OeYS8jsJQrkJSy9dELG8cfb2CrxoXN/5oU097VJ
jGEfyX3uQpm/cEyHANRUN8odE98xcelInKwx6mAYCx3cpu3eGCNXu8vKz/6rEhyz
fxGhvxmiNkGnhXnypJEIL+hre/P/pu7CvRY3C8VoMgG0k39BksRipidKbNdDpZtj
oUTPGI9PGa+INzqMx8wQMvlid2h8/6lEv16CKuFUn+000+E0s+fIkkCDYRrwHvgI
KtwVVHhg9XC4y+f/sVsyM3ah3tWQoCNj8of0UMqXzJyJCrkw2jfBS9r/xWfcZoyB
LjVXvJ1xvaEXq6UfrDp5/NrG+rSyD0uIeLm7fZxTafkO4bm0aW+jp5V86LWcryff
d0h+RopUddG3eFtNfIt2ICS8d+2DQaahzmRD3dPFY45FbcPkIRY3ececTenZsEfG
n7Jr9cgzq+JxHXddt7Ree1bEBkIB0HNKnewDb0CQbWJ8aviQJy4I7ONql11HSnti
Xm6EaVTS31CwvV5D7xTI6S23HXtT7/JFyEfCjFHU/vgxvBm+ip2RMGqtCYJw038g
+LKtJW8ZMN+uZMA+XcIT/s7z7mOL2sAuR52nFuM4vKp9zdPP5ZXbL2BQRI6UfRae
aYBs3IhWTbRizZpOw3GwBykT5z9ziEHGmfGPKLPo6rXI9P9CXjp97J5US6o6aF3I
IZ0kSF733Vd/aZNYefyVjPvyMv2Lr4ZjLiTa8c6r1U6cLx+nyJU7zdzdIFEow/Tm
y1HS2DUv/eZ3s2joMzgB7rd/fmz76BAh7q2jIj8XvMvuMQWdAyc0Y0gFbkYeF65t
rYA4/CHYrLtVouuQCqJvukjkye/CdHO8Wst68nbTqfT0ZUH/FLrEP5U6jt2Fp3cj
gpgOCgkrp8zKIPgUunHst9qSCRbpVMAYGEtOVG/U6ovhxtbydziIDJICFF/kOc9W
InLiplD7Ms1Sc5Wk9vUCqTY7nCzNr1ZC/6Qib6OfRteqvFLBMluNAwotOLgcyP7P
1hkGcZy9UuZEmMXtn6zOM2DN9ZmlmJQooABPBUN3m3IjiMEw1Cvf9eVzNhAeyRpw
RzNnFW2ErqImkvdqBwmGku/eKWT15jp3t8SQzN/FWTIZI1zLsJTY/SE+iyzuQ/be
6JV3XT/SbpbhU8NQXkQWfLUaOg6r5ESjtI4itl8rqNkA8Sbq8Z8de+ospGHUUJOk
xqAdFbBvAxde/WVvfKq4Jje+80zA6wnWIo/nS1TEpikrnt+ykWb317QV/EYrjZq6
cU+rSvnAFTLMZyp3ag7egmyV+qiDXJhYbTRgy2vmgE9HZ9QmCSMSqbGH9g21vNg1
aOtQYGkVJFCMSGB1Jr8+A6J0lZCH9s2TfmwYHlW4dkoQ6MPWPJbs89YViFesTcKm
XXbdNw2egCZV30rTPfvpQWhVuZpe8e/Eeej9Uw0lUo9XB67k7UAMEwwH29HV0sl5
4WCK8CCzGYIACZDAoomoOqED198FvuI6MJvhgu9ATNYlIYWexlwMbqTWG76yPnE1
cNfxJrE/Pj89xY5jgvU0V5PaNWsxtKRFf0nunFUpFKM2l9hc15SrQzw+MmnRsI6U
1/VWUHPebNdi2Yokwdzl8pF2/QNVZyx8dMC2PQSyCQMS9IycroMIX2HxcG9Xg6Rc
cJEdliapDhIQ9dRqZXVeAn66dJptKsrv1Cfi2n9yRYQXZuFuGTX66FJbEWPRS8wt
GMn7gIKZoW8iDqcQFhLFTqScS+Fp6HcZ6JSuAmoZtaOdv/82BEjzZfedwkSd9H5n
0Hx5yzcDss5LCHKVycvGdymNtjkQKhvL+xY7CoV3bgdLEw+SBUhqSPL6jKaTGWne
sTT67++jUfc/Iz7aqrfe84jLTHhKugVe82tGr43pTdXuHhq3nLkYz3TD+8rA+Drz
Luaregp4trge1fEcg8xErWvm2SPf5vwH++7T/gdYgoAyw5g7XIQ/kE4/9rp8Sg6D
83WIVf9/HbrkkzS3FgYP3sQJb6PCX3XI+WfQqR5uKW1Puo+ivpOxQBL2I6dxb2Jg
Vzkrg0UjwvOsyP8exar3//zrikChtH6sGnQyi+fYdnvQBIYHxymWDwsJqHiYkmlu
c6Nc+5++VaUaQDoG2COMxezVdX0p6N3TMscxIkfg8zqhYzLPKRfIU/KF3Jv/hoX3
I9pde4lB3DOHqijQ6dLOoHhdTUB19UnVJbezbcZKUVQ+gEYf7EFlogg0H7TzYPpR
+CQZJ5o5R+wc0cJVibwjAicSWvmIjngMqOhVDjaJk2bLWkWbqePb9latsR1bfB/3
fx7cnfc11a8iBb5SCmiPFzsHQ1JzBybVUwqQDRrdL76ReDM4MWAUczBr24mT/DUF
ZYGppWB6Wrl1NXv2wdJRjWjH2t4l1/2+ElQbiHFAhDfQ4aHrCgn9REnpGlcZJPGu
HY9+FHMkbEAdqx9daCBf7vSNrk2I5i0rIfCgcZhMQsXWFvo3WqFwApqDKTZM6THA
N2Z4H9NrX4iyi+102gztbkeNyNZidXhFN2P8G2nBhjT3Vo49ItHj7d+lE9dY9LLr
qIClrRRNlIfGmX0vL/gjNz9pc/qAEkvwEkeOJ/kmhVUk2SVD/dJGTbPQV+O8i0zL
byIN13b+5uJ5JuTnZYjsO48Zj870pJ5Jp65WxaT9q1dpeBx4HOHQWdfg4Q+TEFg7
IBMKV8BCV+WuY3xSI76hm+KMfrpipJaZGR9Kgd4AePsj/Pa5uhanU44sr2CJFTbR
MdPvtXeMjVvyLMJy/C8ocbhI0pHfEIL9XTD0S5rVAoLWAZNSX9rna4eyEWuF0gTv
+9SQYMMl1bFIyqe82tXX3iLSYZJEOzqIYnINh3VYFvWkhfSqeC08xxqL2kJEons7
e+5FmLe76jt+ntSQQCN1PkjaH+dTRAuF1zdRIzVnqZB+iPJoVh3QBvXBiJ1C3XCq
W0gqvnchmGbtiGJIf/78gtJFQ+81obMvbs4r3HhRsvztqjWwnYaAEk7Y5N7uJMLk
OpJsRC/4+YD7nQGk6EQPTHyrppTdwFFwR8XwKHxro0seS1Y3YfgCuc+s1hSrfOL2
Xb6eZVLn7ImvKAeksome1H/UNxy0XMJhjia8paBzj2D2u738UA+5+6DoHuLCfLjY
VajZc1ZUETLkljtDLNzthg4aJrIUUTuVOyeyfng7xopmylQ6QOz2pcacs55F3sb+
YwPkOTNiQYemwjw0pOk/4ApmIWEbMkYtQDK5IHZvU4Zwtz6jCyaAak88ZEKodyIF
bRptQBYS3Xf6c+JT+mGv6zZI3PYdd4EboCIuVOpHM5cfYtsg2NOQMEhOCKtwodUK
jWNCmrHxaQAh4c0W9bhuNGhfB2KX2xVth0hxOYTAviyCNnEVPylrM360xKhoFV9T
/14dFLBud378UIC9e+oO6+EAp3F5edvVMckxOwEBhlzalPdtPeqqqhw9jchRMFT+
8ycnpTHwdy96cJMqhLTbV+U0vezGI/Oppsfc8Npiaf+psJI4eVaB6LS41xnam9Uu
rcFDry7YWLMwnXdTyumVXSjI3ZvFt0V4q5oSasPq+m/MpywHhxAagsvas7tCZyFN
1KmerNsymYYUjFlX9cKchK99OdesbOdJJUVr4PXFPkoiEsfpN3s/PWNcw+WOXlXD
pA6pWXcxVIZzuPEbljkp96fmOzt5Rx6RhX8Z3IvsmWUuoD9k77sLuc3odTjr9g03
f1BqZvwJqb5uLShycqqlCLzioVwgog3DHGACjvs+g/IDfodNHCeORxjmZx+dJXOI
7nIyX+GOdXz9FTnjttaE9k3rKWRLulIW0qw/6bGoQhE5QP5L9EcdGR4IwZIL7mrv
NUtoA/adqEKeIoMMQahvJqqhIjLAv9zrMU2qiHubUMaGDKf2VEZU9i6qnaGAdU6B
SO18qLf7wQUH7rhq3xPHBa7po7lacoXBsdbhTD8UhA0M6zuF/HQPlRUfKCuw//Qg
KqgM3128ZFXp4zD2HytJ2Ug/CPHK3MQv+2kWeznUuiVSPhDbLgyWHdYq1li4PiAR
u4ncHKVaqnsliDGKEr5gqbP4rsdM5ydPRNIvuG4dPBP1dnlhJ+6CpNC/v0HR2Fmq
67aSz/5Yu/i2G1JyU2K+04DO9WV5KJda/lnsdPSNrQAjlWr1UyRlBb1CRh560dk5
KacM04k2WWPgyW4G5f6aU8nZyEE93UN83wd6d+fP45CHLsaNCqWNVV2QR32Iyzjo
vZv3ew8ez9sysV03aMoASW98gVGfqofWpqpawOAlRySE1kn6wIWInXgjPMq1v/9k
2UFguCBtmWip6nth33mUYta6Grfv3WAUCux5gE8Ei+4mfEEJlqEetFU3n+d4C7b3
J1KgmyHusZUy+2jcLNFHsvpMVZdLHaPwHgeHIqXtVmsyWgT/2SMAv4Vvi6/EmPeE
1hv/yd7hSHDWriSBM3ncRdOVEaEOnjRFekILFrDe8L6IIQm2tHhFMiPEX0Wui+R2
cnMct5TqikN+xWelv9Gkz+oYUC42Ke4Ha3ZIR+TXoAGKXm+jZYs1GYIyZL6oI0cb
idPHZ+j1/uCBWra1coOGDxHlYAiyl1DglTKAkJbza8lnl7QfNehayWr22PbIPO2X
4TRslxweMT3eMgUHoSymzw500ACKn/Vpkb3J4hbqPk9lo8yR6JcEpV5H0KAcdRl0
k+U2SJ95wXsRIP8F6bYkHj+vCGf/O7BkPZDhb3r5z0M6acIRTgKt+NatUX4E+vKx
0SllC+lhYKs8XZGFAY9afsmy4+QXCmRkTrN12akUM8auooa8TNihz4Ht70dB/6yL
06076ofiBBGqssh6i3LITxGlOXs9qV4htsPojmWsZpn7gW13i15p/71NIxORNDLL
k/+usazEsvW3lKnCqKIhsq+CORKpatIIgKi5xqWga5hb/Cdm+PwLJZdfOsJLijgI
GG7KvaRoaAiSVDmKq/Rho7fL+Olu6m6OYMI9tExGPjOfi8jNb5sXpIdkhB3tCaCQ
I+Ior8VeavztZyzkmBOPUPuwKNI0avyFOpDQMMU33sTdwdUK2O/5hEMpYia6iiQz
FZLDKs4lDXWlanUcYrsZLf7yAAj5z/nukboBRy3s9fmrtotGGltWbPoCqhtlx052
vUYyptedJv6eDngdc7bjQ4CFhlp6b+WGPdD2FTGAj2sfD4hiMMYRJBgBNa7z79Ww
q8sSqYpugFVnFIjZKiN5hujgU7NuQldyf8sloJ+Va5TX1jZBasM2xgCacIljn12X
lzoY3JululbBeL0kqulqD7XT8inwFUwyYT5J8YyK+r/3PwD8F6tArvVqv1vG7wuk
U88VRFfZPwrwvSyPSrnYIha/etmuyyhCRBCZdmkhqiZUrMmN7k6CMPXdhzBsreIb
ZqCPrZ0/RK6NS+7xbLVmrb9XZs9Nu4T7tfte//dt4IG09nGQ0muBmK5bMQo+MSAJ
geDbxTWph1uFmO3LqphBNCAL6EIqzfS5+wsJAHrpwTEiP/ntqy6dWRk0caM5BbO3
lVQ/3Smv2IxomN9wh/m1G3EEbJiRh5YM5F4pv7HvaDeBMYKfwGJJmjDTujy3GhpR
Au7138o23p3KFz+wGc7L/PgkXZcTCi8EgPocbSvWLYOfxRETFSwVYLwEWeyBj2c0
abkTjukCmIFOrarAewPqyKCIMV9AcAtBiC2H4ASv9v+s9qOCTeJo6I2hhMCK27hO
kYBb42VPIdmjlGb5E87IAjNui1nAXFrFwWo9mWxNmMILYTs76mwva/hCmoiLVn6O
0AwPtEIhulw2X57xKOT2ovjXSPkmuMq/PpXGmulMj2AoMQyrnAK1D+FVpzg2Ua/2
WqvoHZT6YluBJkbEHK7tVZ7oNNs4KIL9vU7zjkGGoaRmvqCCruS9sNqeUMintkS/
6bPUhbpD7gwFsWp+Uq5MCuw3G/a7WZdhAzMxcQkq8x7mPPXhZ0RjWpBeGJVrFE5A
K6dEnm9BL8QZ8B/fepfsfEZ0/meB7CL8t2XDOh8sm5tYL/rSG3dqgqd4KO5a4pe+
ep2R9y/xar5iXo3J3ocVfUTTYbeqd+3i3/hUHyfdGCyDia1hyYnxrSZOfLhYTsyQ
5S4pI7C4P8fxU1hHsXLSRd54ARNtu+WS+MLMbmQcrOi3shGASOl92fo+zF71PsHP
u1OrsIbDuiy0E4d8jEsc4av1vzJ0+rwOoPdKTJI5+BW+wlTKtP6FSGahBXLMAl0P
BCESaassuckGO9kyw+magDcDXAlElDlIyJgWCkoCVxi21LlY3z6uT3LCrxEhbkkH
GUAGecqB5E7+InhJvsRfYJ44MWdAuP2afHhTCBSgMT9H9SOuX8R++jt48uDWhGo/
A+Aq+zYbGqv+OkHro48egwkVwXOeayJ7n5Seh12nhNKanl+jYvvd8+rVgvjjn4k8
CaGANka9TFVmzE8eWl1k6shhgCXZ/QZe0F5BuSlP3+RyjLASah7C0fIj3ZIXPU2r
Ld7gtZ3ffk1u1bgb6w32AerLyGMG1tDW/IIuyR+r1EgshA3hzPfrJlQfxxfL5BG3
fF82H85nHBdbFGr2QvGThT5sNOm40/P5N5e+DPNN2daOsh6e0F3A6Z44ZUgZ/5VZ
dQxSjROxOr1pU1lCVV+cm9zIMQr/G8gHtVHZkyeB1WEk43wmDiuqKJPO8WoOX/Sz
LtAUMtcW3IZuITK9APSHxBfPPvZ5wnw+/xj1dUZVZ42uiMf5BFjx1FTeO3v1aNrX
lxjHsssl3uN0xwjaprwB31MccrxpTE1BdeqiIksqjgXxLK8YmHId8i4sAqzoGGhv
ZW8uQWzq9jnWMrGSgOW6zP35wz03CW/y7TX+09U/kzsp0ZTmfOVu1pp/Jv16YhdS
80v2Zob4toIST1e9zMCVykKJUoqsf2KhbAohSaNyY7UQNg1NH+UeqFweIgILBcR8
qEQ/rbyC7prOW9pbgGcFPnb3FjFvkAdyAQaQSs+FI6Wjo3ifsRD2xELOyh4s/Zti
/hl4aRhsGBbYxdzPHPkniA5p6AZviwGp17uDDZiq9TYtOgncPHVXNyY0Nn91gRNk
QO0X3v0BzmApOqHapIAnCC7Wp5T/iK/3ydM1fkm1nsyEMcZmCt34ZAdqKtT5llRn
8yfW/B2uVYpGCZDVizM3XL4UdNlvZnmWhbm5mB9Jo6T4n3Cj/Voie7WLKF+2u+X5
CCDqJcu8sI6LgHCiinJszbagRIJ48TziQlcTfWqed81tilxEZHc0SebCkC1s8ufF
Vreob3TqEp1vji/usOn4rlmf+Nj5wEUNni7TboD5RIYrZMa/pQ7hhgaw0LdzTlqy
VyBfWTdNXnacQ9A3T7tCiNc67YXbCgZdrFxHReqWpSI0UsfuvPPxaZ16IYo+benG
Hl8ZlmBS71fzPw+sK0GwS36a9f07o+DahY416WosP6oeNbzpnU+JW9nmO8/zt0md
5DxmapOkWeO5o42XWNWBO2PObzJ/DaUJeMpGDE1xjrPNlLlide/bPr4UbTHu0xqr
bqbuvzOtbNXwR16smCxQmO1+HMJuc4W8anu9x7yJGiOPrEvcACKRXpy5VXW5kvLl
ErorIychCCyrXEclzFmTx2SmtIYJX16Ao6H0dVFddztd9VUBEAy/CVnoljaTAGmt
KhAZFzNbgd51hgo8J/JgA4nTxFmZjR1DNcE6jp7qyagmXl84L00VLvI+EumJAWtA
zHUf3mA/ujNOTc+jCh4gOUpjmWFuvINanJX//slW7D6FVVCY9r59nekZSnztHraj
eu3XgELaF5m0V8FIaFql2jo/8hIUcAKoZsCSjrgTtcENtFFfl9cHihsizjI1rxL2
rPCbdN9nyJQ6IcuLjhN3LicpvmuCSazIGx5f0/y6fbrodBKnEGwTPus+j2b6jHfd
2lT4G0BQjbUh+bUT/HR1qbmjEm+PszflpNF+24A/hY+cl+bskEwD/r7D9xBTN1c+
8h89w/xZFi6HHnY4wz6r5g9W8mehm9XB5J3DaM/fSiJdTWepBsUuRKklU/m5fAUC
cdNjWmMQWhdMzA5HeE27AZwWSMWza5igwQGE2AYgYqlYJ3Z2+S3laPqtGwv3vaFG
86rln+QN5C4N2qene0QeUuJimKgLihtA/t6w+RmHygNK5cOLT2gaL7yCe1EDKaEQ
8ioZpf6bUUECrNTEbN6+to4Yg1IGjKnASl0GdDanpGBQJSLUeu1Bf3BPiHEymgmT
zyf8V+mM/ZfIPqhYNcEOmCducOpTJfOsuQEj76Lc5G6f22Vi7y0oYlCZFKDRp6N5
ErPqo7+tM+BPiBsk/dlyWymTrQxovkSmify3xoQhPT+zPoxDorogcUj33AiToysm
vK6oHgPzWykR9tLZmZM2jQWV/k6S/GfVhFqe2jVEaBme4P9Wdfwv5UC7em83oc9w
U5irarBWF5MVY14ei7Iw2fEgbxzJtCYPe7aSveT0wOo3uvvpoCGXaUVOL0hDxoeW
OPoXFyBpaBQlwjzTPP//JcuuffFJ5e0lLkWjKYuz8tRXsqgYqkUv3toyZ8fT/3aL
lRitvXWFh4r/bx7mf9EIEYOeujEGOcXd5rAkrvfpZpAM1WU3EP3YkTRUz9KG9RcD
kfU7jcCMn6P1K7e29R0mPeiSOL/RT975uiIS773PCdthQTl/71COIXScfkNBprha
kVjqcgs7qOzn1px4/BYRNzlXzUk8q5RlIc0QUWUqS4mS/h/NbvINe/6ia1SWQ35t
zfa78KQ9UjVnzxHpvrrhCPGRb+Nmns1DtLkYCa9Pw/Lvc7aVATD2JZ0GKkXiuesO
1IcVNMDN83BfizRUZWc6foPSIOKx1hgiSEXoZUlaPu7QKDpmB2M413cPgbfMd1YC
9GeFI1+mJUTm3RY1Lx7zsGFuJfYiQqdV3XWz65bOmG6/2KpFqhbJ3duVCR8uP79U
zrd2hzDqhOd3wHC1LINft32ZRFirs+OL8UoXq/JqJRS0zYoiHpTslSxSyYPlNAOL
rOW8VsNn73RZh9g8Ful0SMh7CCZ+ggNV8ssW31G+7zAmAqc52VS6XAMVMwfCH8S2
XZlDAiaxqd2JYFrPkrEylg2KYcmW1dUmzlhPmGuaLJS6QAFRqQ4aXYNeHni4OmBv
k+VZrDrB4Zxi4zOKCnUBMMEesAqzjA6YC/u6DpJ3fNkYf9VrR/zmzvtaxKGHSbK3
i9AfpS4yPjT/aCvSU2Nf3FeDIkEKPxcISC4GajZV4aZWCGOdTYf0QSxeFOo0s4c8
kT0MXvbMAYMqSPUYsqAg4bXSgeuFG4sf6MvXpU3fDNq1WUpLjFQ6OGcLYQ8nJIos
8h9JUf0tKiNMcsQqoLg3HeoksBPpOBZYrBbHb7BOsi8TSIsKGIHB7Cxocos/9PMe
WanSKKBukElx0Tss56zdvVuxOIP7l4YzwRfKzxC7kq5z5M77RJRDmK/M+4u3jzRc
sNUldeZnpRF8PWnaxFvZW48lc1J9Ty0wXCjvQnUO+iNyB3P+anjB3ovwBC7q7uf6
Yjf07x6ZEuudGnykN9vnNnn64LH3IIXcM8eRt34VU+np7aS8RN1XlsmGdR/r9rjF
W/ogk8VCUx9Ao9skIiqsT94w+GaBPt8ESHahjIvjRTa1XmCJl/Y0Ce82XS6J9uwk
P7v/MqQ9l4dG5oAOckw4F8GjRlsBcqrJl9mRALtw/U7hr8DC3WU3kW/gsFbGKn4m
F3gDgcOr+Z3mNRmkLYJ7DvgRvlBAanC032J+UlG7RKthSsJIWu/N7Y0yv4ip35qF
SdIN7VuMhCTDSWDsCgLepQbhE/4jES5sNCRZUNPp+qtK8XAzsj9mUPxCNr69FxPt
8lBi4RMaO4QJhUksBaDLhgZ8xMR7yg4pjdWJGxC2tuXfiyfZATsMQMZgZyMMVLEy
a76yfVbHtXF0/YZ7/UB9dkKPPTomS+VzmPEdjwZhtxrLw7Gh5F5fZyx2plQV0nBl
AcMdlOHFSHc/LOJ8s3Y5HEsbcFR0cKdUCxs9LdeZFCULATLvCu24zfiO7BezRiTz
A36ufdO7TbqhF9rqfGly7iK9x0FMg1rQzORLjQkvKyRkq4eGZhqLf4JGcifjkIdc
nETOX61QbkPT99+033rvpB4jcF9kSXFz7beQSbJzAi3ykakYD8hNEkyLsl+G09s1
1D73c4N5Qf/bO8+fT0v1mkd6XpNx6OeDCC1cxpBb146yRQh1XTJ3NC5HA6d4B+oI
miQ8E/My6KhIEZMVt2fK6Y9oKjiA553wXwkSrX/q2yces1z5r7KUbEG1tVyBHuJM
nk66XpDP2g5yauacAYb7iXRaaiHc2LvBOuRG5zgmZhrwTwHfKDz89aIlWwMNBM4f
5wBnOPGhNa8VCzwwhBruT2NHYDTY/GRcRrgA1jQetL9DQfxoR0wpQ2jvKDFuYFc7
7COG6UFN8HeJJvHEKv3m3o0zzIdUX3B/N06x9aCq/GG+LaQm9BeFOczr27bcV7Rw
K+06epaYYrXERja+j31BGhHTkCQqR5AodqcrhEhHVz61H+qsr3kkmUzIptnYMJZ7
61B2GJfWQYVUBH3AIg8tNW0iG3+5Z0LG6NLRTJEIzfYJYXpYpFlYNsFV1iXbYL42
fulg/BEjbmMX/JiLpmxs4wF9C6APhHwDPaBech9Sl1rXism2SWkz8APV/swne7dI
aiQMQtK+pZNhmK4OBjPVImJsRaIPaDrpuitrHAHL2RTV2sczkhG6L6oTbw//yEVe
+NllKj4+mI9MuW6rY31265pMAOD/M+Z7XQFre6FA84XhJdCA1R9RDV9fgN5CKzLq
dtB0GGalhJvr8txf9UrixCOyoP4Cx4uwZk4fhVGUPj8zBIR1ML8a+Bv9L7+OWScL
Oq81+7rayYmysMW5yCPIQAFV/7LUre1KKm5Q2XmLvhcKzQ9Nt/AWnqAIOWhtB98p
MtFxJABLucOLu6J2KvS1g2Eosnz6/ufTDOvA+FvBPc4+Dx5KgH0Aa8nAtg46a98p
R5JyP1kYGYXQMsVfL9dMUYS4uQJhgCNn27UM+NgfzwMSD6Ou/d4c5Jz1VcPoT85A
BMnrPJT//6PyLXJjsYO7zIZ7emG2m9l49N02T1lujqXXaC+9NEswvzLttdlglbXi
7vIl8a6oPgpoZPkk3216p/EoxvKAjPs53sro3sSt/KPR3/jRqfeZRl34pyjr+u6/
O8+yhFhLj00tcO1P9pABTAAdNaI03g1xFCfvsHLQscyBnynuaRsDmdUA3vcOQNQm
DgeFqshrF4UcgV5m5/LjfdjAHsMY8xRbqKiR3b9zWMiGkONw5azZHHSJeIFt+Ei1
f/kI/pYYt9YA4W5bFnHSx0Cs2cKaJ/41jyU2nZ9CgrDuUWzeAYeDb3Q8XsAV4WGm
YWawx56r/Q5hynevQSMkqOCgp599X0qehQ8XiKwcHFDAp8G0La+uVuEoC3pdY5yw
CXMPVr4wmsV3FnX51w3LWsz9nAn0BqWlvhSJQMbz+6Ae4z4ZzakJSff08tXJNTYh
sXowjzyZ0UjaRF0CoeJfcb7MS7J9AKkqHvK9GF705KZCIprGESsXX9T/SRxs6/QY
L8VfUMd3xt0ahKqiBDuCmv3/rRR0qHFHv0xkaR9lMzviHJB6KYY9uyF73IoVexL3
lyE7ji11+yAMrhB6j5ldsk9xK9CJgUq5y55Cl0WF7p2qaSkTeKW8oQwwCmVX/uvP
GMEtjgMnP9SWYpy/0yyNQq3f9P1s8ImGWfe9LDwUFhlN0J7EA5Dw8rXIIbOxOj+1
w3qFlZ7hZ99zumXwSOs8aKhMbwJxvQ4vc888P9ZYEJUByf365B90MfZbjLij+A4l
3MFc66YKGtwQF2IPSMiuG3w7yyjWOOi63o8aOwJNnAgIjcMfNZN6vrsX52HCWi5z
PmWZtcga4SGvPMzMl1gX3AL0G3ljPRnXGWGez0YkRyDcgroRUyCTod9Q9uDlloGf
p0CKS1eGUw3WuSbKb1In2gVs68e5jpZDgysNP5MWpKjkCabfBkZ7+sxyNVLqtLxM
UUWD0cExgnh+sLbed8s1t7pMrpaeWBtSa5VdqrEgWWAD7DVMUDD77Vweb1lcP0ax
krCkKySCOoDm/QOLd5h8fWlQebzQFnvcgAuF5D/vHa+CxIjmyWlpfKdQJ7ytRtbF
W886wxx+z0TzGIm/wlVOSU+yekc7JtOsg+e3734Q2GB32l80K9iO5Ktev6rvXoOl
xN3gb8FTmT2qMguwM1ROwmN8YzRDUcYWXILtjecx3OmTTAxW8tjUVckh6x+X5KOt
rqGVPZhQsC9ZcN2syd7BHL3t4gklSqL4SwkOOBK0zfufrOhqlMEhXlw6KuJiU7hS
I0a924Gy5jrkR9NkWdYGz+dkATMGXBzFLQVWgTxtzjdjpkWaTY/z+63/99L6HzUL
je07Ysf7Ynx2Hxp0aSR0GCjN/GUMgjnchsxbZzcHaz4Ywp+xfOIdR2FExMnMpQU1
jXjzuoAc6bB/QeAo3vuguuANt1sgpKLHKBz/RJzETXs+LLj8qLmmLtdyIrW1ZJZV
WKdSxaJCBxfNlvC4BK4rRAYQK3FFkxqWQD8y3v0vMkswl2H9pvvzDxtZiQm2EBwm
auVuzdCKrAV09hVyBLPSDb38p4eEJIIR5taziBvk5c3d0Q6ekXQF7MpQhDaCMy1s
WkepsXUAT1gqaWaU3COvQi7kHZj0rSbpglVjzYxlFGKMJ5PaJcWR0NjJcAOq9v6s
XSwnLPcyYwNHs+lSqUQjozzR8r4OKUZDnQ8yRBIyQXucbj6s0+8WCQgdFlZvDAn4
JQ2n4+RA8kkocSlQE985Ah1Dha1d4gt7Az/ffsoUKHhv55OuBbfHtijTYuPfdxLC
0AMojNquDdINqB0GVsfRPXOspz7d4RyvGu+djGIVGXyxtzomSl9U2SDkg3bU9Zrt
oWom0ihWaoMrarBDNFPs0pD5yHVkPhHjdkSAWPb5jyNEuRKtHNqSq91itcv8SIvn
mD0lksYkvwkXPl9qFLa+leqBRQle+I8vHoaDw2ArbEY9nqoRdsqluw6kggaR6KCl
P9oqJBAGCBExSS8vB6SeFO+Woi6ycZ+8FfoW9TaTpQSbJfwo4PO+URueyLL8Xtgs
7gvEe3qgQt4Vhcq8bd4rx1F+T3pdNvqzYjDDNc4e7Vv/2J/pPCPpAS4kmUfn+1Hv
HwD2sdWSEV/O+5jlkO2iQzKQDGCVxcKS1AeVDq2J3GbPQB3kf4jJ/vb1XqODckL3
TnPQnPSpzzz86ec/c991yNzIyqwutUX1ouAo6DFISPzDb0EsH2llbROLKHOgMSEh
eYPw1tdBRNCNLjUVOe2F8eIigFixbR/2oJ+S9dEOBJQVPiEsXFmkEWo+nIlVGOOn
l0VXMitU4817jFM8L+BAXIqEI7vd0HGZQoC+KZtgl8456myC0YgKcklcrwNnMK9+
afzljDhkb4o+SqSL2HLSISHLjsZJNhWfV1z5SPdiiPMqqAEkwqZKPa8tqw8MOsy3
TmNsbCCod8A+rxXzAv/OMQHSjQG+2poNcX/b9gobSI1IefxSrMuSPquFLqUBHWmI
o7pXjV2UpdnPDn/I0UYoVPtYb4IFGaC1CM9Up3U4yHGtN/MOLnBw8B09wHqS+ml2
nJurmnIOeMX1HTB1BkiAA9skoyvrCWsZFI9TLOEKysvydkKA6PydStd2Ncd/yivH
J6RywN/UKQ9aT//X6NSjkIDNe802bBH4nv9rS6IZhA7jCIlwjV1q3VMbE5B6lQ2Q
8CNl5x6R/cfofw8+jP9dutyXEWxUi4dbRIReIqtqNOd790lT1x3b6CgFnnHVT8CI
hTIwJr4KpORJn/RBjpA+soAUvNZ7ci6cwpfNrFDQyptNoaySeHYDFIkAVDxWmpFO
2Q/ZS9tjEP2NkHaAlAcuhi++DegR0WPNM5peguRWK4WyyrdTFQqP21sAb3sHGjAq
01NVVcgtrY2FO2zCbcoVz6MDMHsGQ/d+6mm3YT7SgOZ0fH0ub7YPkAPJpCmX05DX
CP+kdOf0LpRwEIYTLWXn8svhiXOVG4l9ED87IGql/sGdPCWjCRA0sfYNmS7DeZxw
Ln9K6jUHXaYvPqSwAjEYS61XIP369UTUxVxcSWoBXOlcvug6wItLkpz+OdewUVl9
aBPbq2EMz8+tCPUdHcIxIlzL+fROLTTRCUzWFDG+7ONgUzmzoJICtS5qZNz1zCQd
9OCTDITwjV4mKwjpBllbsTjEy1dtdQuIxWmWorbW0TTHEkhpdtC/KIfMSHpW14u4
IzxuBOiVbe5EyBvxGJsEGPUPmp0A7g8MkAmbRoSYoirOQrvBoy41iSSOn2nZEW7s
4udi5DE/SKrDSt4R8MG2sEujmcEgeZZMFATF4AyDdR3wfTbpdD4AwfDCQ74n0UP/
t9dIAJe8ljco6mSytrO93EO1bjIrWEURIIL4IcygVsRPR/xOW1M9Dn1KxP328AiU
PIaFmyfeoUwdZPXuSDIaYh+2KK0fD5ZG154+1WPxF2nVpTFnWqwQt82E1tj/87s9
wyB2iVGOo5Y9E3tYBbgs93rSW4aeNPjgFFeHI8Tm9L+uGVZplc5wjvGwpzszl9B4
6rLA4bZBXjjZ745WIT6uwYjbA1T3n518yztwkr15k8NkpZkCYmnrQhjVQIQ4L30J
6JffMj2F9TMyAsl8cw5PflR9iCWvEzF1kYwELixfdF/zOcwN4QDGxjA0V+6nRHV1
0QnmyVMU5ODmB+AYKR9g4zdw8g35vQ4zmtQui9gKYO/XcQVsfv5PgrxCfCWPccX5
CxVIJ1VCAcfusRa9oPDA5Lyv3xqIYJCAfUGBD1SV8kJl667WIkxrv2lsh5fBUsmn
IdXoBAFYWNFKP+RjVX2QeyquRqKz7uOr1t3DMMM6E+t4SvaqQSRp++LmNMSDcsX8
+WWXy0+hnNGx2nJ7rBrUuQ1Esy4XkVYOfhmLezRyDzsirXAIfbubjEDZp/OFOwwr
tBhXAhqlX9N3tFbcSUT9m7keOAK+UuMkjSB3107/gTBIOlcRWEll0o/puEQ6IKkl
Yr2KsbyALs8Y1HG2EPeSHPrJcj+QQhz4ESrUG8H06nKf7RAZq3Gr+oXJJTgxHVlh
gEZ4I4JHfoLYVu3LRZ/dzM4Gqy+KhtdwXckJDuQ412w8YG9KPJtixbtLO2chxFYX
tZGlybE2VFOCOWbDPr/o4xuE83jSzQcGfEOchMea9X57DYtSC7SCw5KeHRaxlLmh
43BuC/wSqYrVXYeGumsLvvnhigCpkvcw5hngMF+ao6goqpRyaVFiVAH2U4TO7oBy
58ncXQipJBtmjJ3VbWwnUOgjaC/QTzbnc/Q+HAkGe6ydYcXSo58++tBQnwIIr84/
zi1KwoFxLpAiR5i208Mnq8OS+08tj8AIJgEJ3N7by8ZCSfn6ahRoO39tB868Tuu/
NPCGODOxMK/mZUNbeHIJoLI93JvsdTJHx7XiDbgslsBW6pXav+MX4WIid5tdi+8u
8svun2NtQLB1+WrvyVWA8/69LGGam7X75phQ3SrAi7ugXtc4qb23nhFXyxzB/BnS
7JTTes3HgNJLwvp6MKpRfO5DZJco9XoF42efNPS91hQa1CAw6k859Sq+ZuokJcq6
mRWW3xjcAFCGLufurgotYK4srjOmxD+79MFOPHJHGDoKL5HK5yun7DxjNaeQxqwE
0sqEnDQRi80ReFU4Jr1MmhAw7KbizzB+xXD5Gk02RrLAGTvn1I3fkTyGz1u10S4I
DbNgPxlqesLRUpKtUVsJ9sK1alQ18RDMHKXICU09YjQ2Ewv/3079p1x4QteRZjOa
ZxLocUNTqjWby3UJ2oS6atbOgZnXz4M6IpLUmG4HueQh9d8RMFFHLypxnQBz6l7/
2qm64o3/LVgEwbI0+GyhR9e78eHh+vWFBBW2L69flco7Iwx+KaxHExjAjRA0MBkc
AsmBGzSLsbIzduKn+qsLPbk+SGz+ZgnWtWEIKjgm0TAiJTnDj5PbEiNGqyZOy39o
Zsn86esc7A7daqGgyuypGDHKnnttzw0ArH2kd8nH0WkIPDveGmscXMfmFCkRmyL0
RxI4jxplB7e2z+aZFQHa6bHUMHa/QwDTJIe5lUDjOuC/7DcHagZFgBYxC6vS7Wuk
oUWR6Lg1F+q2w5fq3e1yrhUe9ve5z284bBLM90r/ahWDxE6fjxngO0sOi0qFi/do
+wHW+tsgZdiCCMZ822jsYCXGldlhdGmfy4uRLKcC5HrgNDnsyr5gQ8uFhgBroCE3
B63myJ8n1lhJ9H3kRmVrGbiwnJT2Mty8XpH2RPlkQXGQaqMSllrqMX8wGYZtTzHo
fx9QnfUEY1P5CL6b3tCOmv4/OJfT0BmDo4WPNcU0umL/lghRl5PYUFGYCTHgjWP9
R2eCoi8MkiASAzQPRFaAdeNS8jK52B3E8Vp3JEJqk4FP3YBSMaqKSNKlwjW+a6dL
4HdF6tpgKfM2iH5LYU/gWdOgAqQUqfbPLaQAfD3u3W44cALRPpHTBw8hXfYAuN24
0fQqJm3Ib99aLSi2YPz/oO1y4n03oC2gCUUtt4Cqj/OJ9JZGtvkq0eZ/m3kHj9ob
thzAz6JwSeSd4xiHkmLNtGccilv/gv67NokUzwVfoCSy6lAihDwrsBGzgoPYRH7J
lh4kfkrIuGpX8VZBuGAH9d+tBNdk13M6CSDufLVRyppRm99w/IKD43LMAzXutKKD
i2fPnZYofkpYAYiaXalRUK42hv5wRLenZQlG1uhy4e8iXjI98/W8Ft1+tmrxwMiS
HwrN0cmj1ApufKD4QKENC0mwMEm4tLGAv1m4f4tW2ko/gnPLzI2JagJgXOpjIhPY
xdhuy8Wnjz1lo8sgtFyrW1eeYTwtOz1lm53WxzxV/5+czZv5V0/0YM/iVWt+iJWH
LArp54sJtfHcbStG7Vz1fGtLHue4vtlf+4/jnUWmr3sNaqI5VSwJOWDT4o5+wi25
TgysPp/HKXm7k2lHMR9GdSGBvAGvBQ79ZmYjzjQVDEZhQZbFzLCEX39BAY7VIlsk
YUP38COHFln/GBp1YJeL2RXO2Zp1u+g2njBNojxnY1mh4XywlU1t9LckCQWuH1sI
Kz9xNz+++d+0AsOHZOCecfwL8recld4rWBE1o+K5YaBGglfxV7TDvQrZauGs6WU+
Zv1nWquGOkw1413EarJ32/73GNv9VKA5spLKMHrRmdHRu7ZWRwthgAouXCkJMeFk
ns++qImumj+Q9M4H50EQwfSbjidTvWgjMPtVuv/r11CIE+IqD5m924IbYyuofS1x
FnRiCz/Ei5CGs8ycmF5kOtykeZ0FeFv+XScXzLZniYp+xdWnsewpReXZZTysv5n4
rLnIljkTTAIyCbErZprgxGZB7t4CPKuAeUtVrqeDCSnO2tqCzCY/AsfQVBSmaWes
0hYfSuOaGrvrHKuBPoCSY+ZBFpe1e2HVvFbRglPj2wC2XjnzrdQ+1mjgG2jRh7na
ff9oddCK8ApKmMMUSVy6BxZ4YCrnEPQgHE6H1B7pVG2OHvRK8GAmP8IKxkdAQocq
dSWNnftce/R2Kx//vQstMmJLEGLhCPkVRLGqvM6T/WjZRDVdBz5c04eYCA2zEn/f
fmVUFZE39uzAy6thkaszYuzFgGwh9fbsQ1Ne10QEMdbSYYSFykDzx5YMXgSfP9W5
ovYSpKSTkGcH6nS24nqlcr6erTWAYHguGe/y0dTw6RG1m06I9xO08s9tWNpcQahZ
o6JgnByMfWYkjjJvIF3Gu/mVtWVavH0lmeJsPvAXODkc0kTyZnoLTtCfBMcfbvVu
pguf/RmzWLdtoqWZG+4ayIL/0R/2rJC6g/s+9Y2ectHP+e4QjaTeEtMiEDWWtQUX
qlWpP4t+uN729ZiGLAprLnIHwIa0Yr/kdMIvow2yNbVz0vQmC9evdwjh7PFEdpeJ
o85D6fnSy+tRXS7wWC350kMCBUwdRAM3ScKxsAa3L0Lyd3hpg/9GgYIiZuEwB6c5
sg/7taFvnPft60deoh/T07jc2lMYAVTqrublyJ7tqUOByYlPsCmitIQ94I5pfD2d
ycofbIERvCn9paAui5ICeq8h1O6JktF2k4eih8u0FM9X0AqVyXIukeEZb4B5TxwG
maZXmotTvZ/cxepRcmZWC5/q6wpKgYdA2jN28sy+YU8KC1gEQ4u/kAzb5Koi3ebQ
RupFxa0nOltWqp8XFuhG1hviZjbFMXdb6N4BLLM9RGqFRy+bav5Qx3cvD8nEzaBN
FZcAibir4U0yVQMqGR3mVhrtClMK7et/Nk0+2vDExGMNCxUX5OiHHSlflK646XZJ
7YqlUdv6V2cJZnsurFP0Kpm9w4+tYKhy9rp+185bnyF818Cb82RnaJa+0fO7oNXY
WvEWIh5nvxUprPo6gL3qf8dI14tiySIVeESqjQshHTkVwQW56jNZYMkqmAHC5Prz
UGSvO/Wns71Kyn8FTwETDIhtjUH2w8GsRXqqGg/plZP1G45xpeH4KmTMIe2C0iKM
RS10hze+wxQsNraSktG1koMnZXtVj7ovCMJOcBxS8PizHbTYdJTBgpQxElybmEYH
EJ9V6h3aVmIcYnvvTOOZNbUPQ2WzhQCP6p5MALdwWwxkEd6aylPpZkHHS5SKv52R
a5H6GH5kkhgg2dO3WoIXck9AW2v9xKBkfVEslf/gC0C+LSaYHMEQhAqwBuS+xD41
cr9K6uJh0eDyRMLK1GX5XXpIjXfUI2vbypklPgNGo0gCnKWTh+G4GgM1Db44qUl5
rRcLq4CoP6qKBaM7M7RPp+Rl0Rn1mf1oIgwTIkAwuUU9qTvfviOsXpc8LiUPkpy4
xSjpL3vZ90c097X73mB28y0V/jgTqBP4P0cqGkgD5Cjz+LKQHY8tQYkrTOxSq5hO
TLcQJin/pqIApqA8zHH/th8droXoc7TqnWhO43ExXeItd/ghuxjQ9P6ERRNx9JHP
Ea6FJEREpPB71TEXQ3Yu+Wca+DvsxIk2Ed4hfOf52PSxLqTURaWxtgrDAVeESZlI
gN2Eip8xcCeIEEjCwcppRCMnAuXSMQ9otx02NU4k55rV4XZ6V8qCzUEwSCmaxqb3
dST5RGYV9Ng85kmgHIvdhQygN4VLed9eoTNf4PnWABw0jlia0qpBB2Cr+E3u1ZCM
VXU9V5CUDi3jnDZ04lvLdI29TqfZutxif9hg4TbXoSesgHXUSS/ZhGOGeNgvpGOZ
clx3RokjF0LLPdaMxm0vl0Ws/C/L0MkDS9+W3qOgNVuOarfeY4TM1Ay5+AX0g5/l
0+WpoOv6eg6pR9kIai+ihvQhkM0TVp3AMXZeRquPgpR4PrAd7i7U2IqI3vDFtAes
ZQmQIKOR6KfTvEWg/aVEo8XXfu7ygXHlcWii0aHbbBSq654BS0ct6CcapptjRe8i
us0zz4cIHaHdqIyKN5snDaUqsu9BBMyZzFsbXjgC783JNgTJUm9mj8AaZkaewdi4
VWK3BbFBSjPsaWQltIyGCqKiyYoguQ+4n8w+waRXhKGop5L2pq+rxx9dd9IApzOT
4pAZ3+ddFZPzczegUFlV+5/NKb9dY2XTU2Dtx3IiqqwfYjO6Zt1OlFj92C3InlLn
pGEIWwRD8POErVisIdWUjZnfTJAM33MsNiknjiukXMMvonW6ekUUCW/s1iwsm+Ly
M3RljMQglUCZeKLTxDF2x2svl2XX7/h08g5Pb9tMn0hFuu4dADpJths9OUi3GEkz
5J9n0vAoRGzD6HM+Vou0xov7QwkpXRPuWh+PafLXXPoHHarXOZRcFbt3kQbshsJR
0Sp/GqsRdXWleDIe1oPOKakPT5/o4WHLm6ZtAts9fA2MkIKKi5YD2VCp9/CR8X4I
hsk2fo10eqmc9ejhrIv22hZx18sN7wHoKPzvBmQuNkJnt2I8B1HsRK9UM6p1ZIkT
8zCb2CNMPchAtQ7PPndso/IS2HgZqnoPX5Yq0Ab8WWDegsnNbUfFpRIDc/T28Hv+
eDpI84xBVx+Z+6lode1V7WM70FUkpESJsDpbzrKTWf6Z450fH71JUUEb+hob4bA9
IbNExguPEEMTpqLH3LtaHXIYc2tkMaeXbQqvnrQUIbYTRUeobVLQjZgRA/jJMzqa
tMKrlHibKHKlBrjfluuTaWZyUlTZ2YMiHx1HoCKuNB+8EfHeOjUVZMkNC5ov7cyA
Ap8i7IdWF8xQumK6499bVQA9NggL++rB8PNoQY+dqP6Y0bJtRkLUSpQBCPjuBdid
n/7u0j/O19cpRC60fwl3Okc9nb3r9ol7jgsNlcrFZZxSQUgSh9D3dIP6dzzHFkD/
AKAIYyZdC+G89SfY7745r0rVO66HNXtNGCCFQLgfULVRO7MPASGx/aRb9WDdIpxo
cUlzvmEtlWh5YJbBCJtlsVaZeFnzpM7YkR+sgXvRB0UmbkbGM5Xis2XYTAUOGcUJ
tNgKYV8n3IKVjt7b8VeP93B7dZUS1/0EeW8607yawZDBgZIjpgzRnwLLmmghANKE
YGdw+TBqZHfKJbW//87bDquHqj1QxR7RJ5ZsnRsO4LVh+lIancJLOrj8wcCv/Nw5
IjrjWx9+I7oekVv4VEGpSyQp+LbzKZSZhwqa09UJ3BJzB/9Ap5Zzv3osHdez5Hx7
QsFcAnHLJc40/RdKBvmjpssIZjFTkgylkFOcqwPrJB+uPn30Ba2RP9EnZLmBU4Wa
jVrC1A+h6U1Nx8PDd7cP4j1epEGHiK9NpzMCQDRaJtLP0Ueuxu27StGMuqibIX2r
5xuBwXSpifiSzIAJontfPWJiDiv4pBEKxcTkFf6NpRIrDueTda3CMDqn9sVp5/nq
ITTQA/5T+1R9i16R2WQo/xFvS3QCEE113ytVqTWXhBlOPvADIotH2lFcQ4ZMOoeV
Wms04mSWK9hL9Aj4rL7hjxCzymTVvXIGvsUpO+EutkEwCApo6NafdjIyEHrxOSUS
bdmv/WZCdGhvwgHRuharLqOWxlPGzbmfBSZAC3L1k9U1gsz1RMDNqeva9GCLLmvS
eug6E9VWX6zJqCiHqES+BwbfN6N2Qh/z5VYtyUIwDeke+ysJy3LeDuVjVHvOrV8T
oRjaMmR5VZemjz4eCQgbrmC8Jq7Jlcs82v8oHp4RrF4shq8ofGLR1Cgz2C/ukl+x
lA9d3VzSKLy9S3XOoxD/pUBXcKAifgJ5tgtCZ0V+u46ntw8Nnts+03zH9nSD24w2
z7c4GuCg+JCOXOZZGAUMj7s3KM56rXtl4SZERaV9Bc/IK9v+8zXq8tbpkOVQpl3G
VPFObASTD6cdXXz/67rqggXDhkZxrqmU7ehAVGgWzazYqu+gk8vR2l5gIe2jXyIF
5wZG2Nf12c1hqnP1a5/K1Fd8r3si0LJHGPOKPv5oppJt9NE/OG43gF3hqEr2S+d9
jSZahuahsH4hwotrLDksLC1wwItJVX2Q73NSTUSN2NdpRTo70A8uF/58ZKGnnESw
OQ0vf9V2B17vYqRUzrisVlWuttrFetEjvm8qNMsFAEE3BK8pK977WVjtUvDgShl3
g5mPiMiuhQrqCRiszF/GAaf2t7tTGCHP7d+mBus1SAU81cvgj5V7U4zIWdR+9+4Q
dDs6HBApTzoaxQcfO7cwcV77rwHBXRsOXQTAm+93FFPwtjrNl2/FXnHeT+nfBXvf
RP3142GPa4MIjdS4C0mu7LBX/zI8PHYrBQXMhMY2AIGAkYp8g3wRGo+Cu5jICWhO
YJSmEb0J+xq0ztoneC51uVCht+9QWU/ZL8rNUMpYpOXp0FzHSaAKTkyCuEWGoKF5
HgQO7YuH+m070/D8KR5h+HihpfNsQ6QUS/NEtxXja3U1f8iVUnFgN++Lk8TkaX1p
7+jJmFvJ1jzup0Aup7W6PD0vVDxhrmnWp+elhCGu5e+WJiM7ud12quQb3VTBZivj
VJ48lN/3ukxMTTkTS3zmZBBmpdwbsbwLqmN0McCgLr5m9knAkNUbqwoqD2zuoWvz
HRAbuytsE/773Mn2GI1ADWV+TjR5SoPHiR9nNNI3bB6VUBIjRZbLu06Szl2vk5Ao
Fk19HvkBGcSrVTwcCnhi4VQt+fuCWRLvUjQrbu2gkuvhuaTqTnRzCXSjJ8Hr9JvE
P5SWqMtGozf0Sc1nsYRoIThordQEyy1HRbhsnkj/a5bhFV0j2L1zBubegB9vn05x
sU3nt8jDoIEF3NP+yRuaWb2FkFIUHut+dzYYDsUkGz4e24dhAjrflsEWuz5YJiiU
RlOt3R2XM17vEN7CdnoM5MF1oTCrrcDInz0o3zOuG9C2CmkT0gur9qcQzc1WUsZY
GvzLP6nl4SsGT1hH0Pm1n054MMipTRDW5oLSJkl9095vpII1jE+hpBMo6fXDGAbw
ysJIR58lQtnW82PRCraV6CZMhlJj1n244hsEqqwl/kWdD7fFBabjg1OFjUF9kScx
3AyHWGGplB3bj59Av4L08Smsm17NsUzQIAZpgWv5FCnj7h31UPoehVecSucCpd1f
Vp5KOrt7D1rhArkOa89acMAYFxdJoVP7cgoURUmoMcRJylZnCgFLIcx8mPeVhj8M
Fg1j7tmhTu5LPobK6CRBux3hUASPLPWrPtHBYmFoHLGwVb3Fs5LWknCwgJ0xL6xD
L5H+2Suktu3SKJmha5vJwenW+7EbioMh1QKSoHKKdB0z9s9DErc3p2voHqHd1QRs
pdzXQa5RsWmDeLDOwZELflrWBQQv/a0kbztMtpEsqUslikAOPKEsUGXvnD7ukQCJ
qNgbN98Cl45PIM6U+A/AH/B5BtKC2UVZDnAr8lBtiQauc9zr941gxHJOGa2gh0mU
hNfQr4FrqIiOSFT0c5rxo7IBkiyVYfOJa6NHEulIelExD7nCCj49WurgAgeyWN1k
ytAbPTbsp0vuiklXjFhpUVR8Pys9HRoE09lxy1N/MDwe6m7e2DTQLOj0x0bHax8W
ADfyKMLiP2k6/zgirVhXv8reR+JoLvjx2q49WyyVXzXVzZ91Jy8gCHoh5NkxOKjI
qg5wqnPng1cfPnSG7cZwy43D4j22IvDlHkSjzDCIr98/yvwwE2T9+mJ2/5wx6Rhc
c600UTfY7KpiWzTKdbesGqhm8Bmz8Cc1A7bX3hfCkKTh+qESSY2C9xdgDOd+ore+
3cP8H+6kRn8N+ROF8K6BZi3wxffTU1sQdONtxguaeAczwYLaC4EtWzLbMiss4HBt
htpYUOesbBdBN4CtFUu9MgXkrgLKUfoZaGmCaHHZ8tfX5lC2foV5QE523Bbez5A+
HqYkQVDR+gStsdA24lW1Ps4qHRzspY5pe9GCIVeVeWDrsNFv/hXAFBEIy/BmWaai
kDdhpshWcnZrjUnbD3ABphsiclWvNufTqkqjNG62i4tI8TlxmC5Miqgy+5qfwdBH
cjUtUVkQ0aq+QrmWFGmpH2mCfCqIdOtmzKbo7YQSIP6zy8SzVugQ2Pl3zm1IYaGr
sbQLMRiHyBmv/7lDr/Ulozdm+c2V1iHYzDjQZhHLXw7p+GCmkirdIN6/KV1VtRe8
LLzig4mrN8VJ+UX84x2QugwOdIfpqZ+LcGHGd4DzNI2itDAyKBqMPV/+gNhDPa1D
06JFxNlh6AX6Q5atdQL1JQUm1UD+Rr9SFKhZMtt77yqba81GFiG/6xd4kXJAsrDA
JgxiS9VRlAzDtxpkggoDWisI69oDvfvRGaa+jen7excv32rhuz8SXsnX5TxXb32+
dltefMND1q6h+lyTL77Lk1VBdkxzXM9OnTNbjYJ6GKKlPamM7PgrVmGLJ/4EYuqK
2bInxogO+lyExk+dWTWr4jEwbGBB4RBqqdVa6/fdfjl3fXEh+kt7y6tQQtR+LZXW
qivB0pGhPnUfrphRUVQhFItI28UoXlsOD5JGGpLdvU2I2IV8iIiaFQVvbYUJIyP0
zOkSKVAuJ0D56ehPGEaXlmZhEOPdeahpnsw8J/K7uQsuRRrH4rIutcp9Wk7EDIge
JJTyxxZaUzeDVsun7iboM3R11R9bxdcCmb6sqn+FA1AYLQeDMjf9ZQoM1SzE6QmS
AXOsUtgNX1oPmv+6lkrVsF8w8mfJfVJOPiC3d/s4Se6VNs5ZV+NsmV4QzqubW/Eq
UxuhlgoostSu5bCRZnL/V42mdiiUapEam9wLKTLEpUFWpYQbWBO2Y6WcmGpa90FX
3ym4UxJpwiIqUiiyB4VWW9APwD1Bx4+DvJjBorTgzmOG7+p1B0HAG72tTYKToRhj
LBeL+ZPaVIGbu4OCdtD6dhfRYiqmzUdJ/EKmnX7GsprXAvcwMd6vi2mJXzR5674X
4Q/XFX/GGpR2jZzA9UDzu0V174R/gn6EYxWkwSvs9ztEJj8ttMA79zcjaYOtY8NJ
BvIpu93rddcop76BANSoZ4T4r/U6oMcOJozREH0eUeFtUlJHnXaUo7uIKvKaAYNR
JM9wLQzq6MbmT4uOEeoDCVMuLesXDQwCrHQWscPO9kvej6DkeUh5bpaYcXUK8lm7
ungQ4sbd6WnCL5B7ldaX09xiAyOcHaNs4hW7lMco901E8vAfiKyFohuBzjhFXZLj
JJD7Vm1cYaaRDodMTf2I1b0dwLqpQknuNjsS7Fp9nIfxwQDW9NzaTPH9Encx2zbB
wEagERZr+k48ooy9RDMBkpw7c19WpteHbc6KIcKLfXsAIyp1KjszhjLm7u0Gov1p
heV1BhXP7n/5RXasbV5scHN/yfoh0Yg9acNFXIABsnaKGWBIbMb4ewZWKqN5rvqF
Xphv3iLW3W6pVo9nKzsWGTvnOS/rkQy1AVQ+2dh4wwZ9BOEgDRfiZL/jYawUoHp6
LFMfSsJZZW/uzZpek559bzST15UxInooUtg0+EHoYsmcg5+iNKp9XIwpe0svRuao
DlLQZyfUJbUSBo4R3dRjYm2XqLD0D6A8MR4Q/JHwFB3e8nyxLMFuQdM26jMKjqlx
tBjT4XhKJIq9bhPrpHQQ2tZOJxMRb9eoj9W8FOkh9rkFAe/6yszuL4JxEsf+hzUH
yOXP9hwfLdfGr7Ii7A51twX0TfSgMtb+S9jhJkvlA3RndleO0oviibHjL4gTCclW
40S2cOQtPga4QYU8saIfIGebR4Qnk1TBzUoRKD098aANd5hUFyIB95GRK3ZMHUvd
64CblPBmIY13ZNMNaOWBIoo0IrtvnN4snDWHjY/Iutq0caE0zJCXmJkrfM7qonWW
w4QE8r/fEPbtkNKrLaBtc1yZXm+uWHs2f6Ywl/GIVAIw5LNm3kGZ5ivMJ9VQCQcH
yLzNZEbKMCxjVlJWaL2mAsuHnqLcQ4twxYv5M3NR//x/qMt9lVGV6qzSb0TH/OP6
ayDMV7Rlvmc6G8NAhTtTLyERsDrqj1owjF4z14q1+QqkHunFgWLaasYKBdFK0xEj
5kTUWq9/4tn8Rjib9qPTq5Dvtv4ZWhse1E6kDZUurp1L+LyJFuRCLExxTgxOp3vb
YSyg1cEplMJ0uVuaDVpECOb34tKEeosoprlMyjnBQ01xAyY/rSLisbFdA13dHruX
g+KmislCYDuGifDwkWd3bO3iduZe7TTWKyiqVYSj3w2w0ygcA87B+08QFKOjnzsz
YmWjO21x7GvG/wWZJPcVgFPQqwPyyJ2aNuePy0kbScUpB9WuaYb+jsJ2wd6alqIN
MIb0tnL3Fuf2jNdsTHdrSHnN3gt/x/1YwVQYduQanP45LuIevml2azHUop0MgfbV
CxW2DCOuiuEKpV37r6eLQga4wOADFg1XMICqo4CEE1wPxX+AWoXjRSPY7rBnsuie
L1AwAUYpmuDpGG+p3jk7L84pHUaHhPxaNCDZq9w15emnJcnkDpE1jT4eicTX9c1o
ZSfpBoADdB9FYDZ1PoDHZZRTSYlQEguxaykxYTUI9T1/jweFXSDDq7boGg7Md2v7
WeqP82uiVu0MdI64unHIYmbsDt2r3Wf7KITU3FylQ7xdns7C7TZF/6BGTcobF3kL
4O/okv+KIs5fHxMMCwQsivLNT7kLU4ksMwXeckZLP1HPUxKiNc6f153C8PB1+pmu
hFUmhqhA5blPuqB+EW2qYBoDuETmjMVdPqi3Xwfg81oy5kyp25Z4UpFyIU8+ibwp
QxO8ZvY/ga+eZ2u3QONPbgj86FrKq2JoZkphMdUL6o9d/qrzRYfTnbLqbuYVM5yH
YX+CkYVaTNtTBRu8E19QROM8t8qmS1oNWt0zTgvsu1/2if6iMQkG0u6i6ZytOmmA
QER9VrrQ6XoR6yqMjq/K45b7tE0m+6Hv55spldjXqTTDjVLV8Qi5BtIlNb5rJbHo
FyXsn1+BZSL6QBSTH6X6gRCNTPutET7o9V9JXu6lQdJU5o09z0gvtgEiIxfeLIJe
Ni96zJ+DYfDot33KRAppBiQX5ukOSKoDw+lcpQpnaS4bvr1GHRujxHjb/Zc+LS9T
iOZVHGJfFZJBXqtgjmH+0Ro+VWZA5IlRkTv/rfAsTrb7ZXOLItCN/i9FnYNiKYGO
+15G1k0Tn19gD9IzXRhRNwpFkS0ut0lfz9wbLbzq77o+GzA4mamm2WkyIUFFSRbX
7SPWG/udvGr8SAIjJQwWGAWnSDyTMw6hUOctkC62vDpUOpFY8aYfvbBPTQy0nBCR
eVWRakwXWF4/zojNEc0SB31MnkHZ75SCoqexvt7aBhYWQ35DHk6ZvrlXhi5r1p9N
/iG9WvNYEO29q3yf/708p0czuLtLGfC1lM/nx1D/U2ZB1UNDKa/sScriVeKXn9qa
JnI4n7+mDcgnhHctO6h0oB/CfSAI+UDrJucO9cKhnGhlm+Rk3ACb1STpzsWyX4wF
Np02OxiRbx2JnCuraGFkNPV9M9ACBmnIQiHeErU6l6zIZTR44QdsYWCwFc11RhnC
qc++zEGSfNkFIFs0ghUQKKQZ21dPh0v6kf8cbvIg761fTRk+6w7AdvCBuiFc91Y9
ObMW+gbGjfFvwSF8/rLt8T5cpf9BkmznUZb1Ec1YdYq74ftgeALK48meJTyPf4tz
+z2giBF+4d0t8sC/FkS7Rm5H0jprlU5cwROiYsO5y8RaPdyYuke/s4mfxnsje9Kx
XyTdwaLQ7sib2DxPJZi44DMryen/WrvIS21iMmL3PGVptgdc2WOGQC2DAlVk65NY
IiYlusEGEM/3mGOvfFGF/1WSKNuo7vS/3oP40xKDRuewHRcw6GnK4wcAYgnNITml
WOfTFPHxeKTVEyEYtgfIXMSoUfAa3keJGlMTrwW4aXXPmZsrnqAa2XL8GoifS6E4
H+O/r3ffAtK3wUACNpTiz3IuHWElksZMZnpQtVu3qLoEEW+L38RpC2ySizB+vT20
yqGKZP4J5UBa+oMI3xS5C+zAPIVj6yGPLCf6uWF8Jvr43NXFNvGlN4qGN1sJU0LE
8rNYvO3eE1BTvjQ9lQBmkc2s8F/KVQDHbedC2tJP14F4SER5ZDJe/kEyuQVHEN/C
MHlpzoopoJtTotS1NaQtrRa04/6Brml8jnhxooXxSdOTfd+IsZNAJJVLCHouBqV5
kNskqKBpnD80YWTJEG7+6p7dA/av1uuQhXQi//AgItZNlOq/22NHBZU6HaFAlbf5
2j4/0uxlhJXaPNZk/CBxo5687ESOLnM2hHLCJn8r6sleZDvx5wyEH3W9DDYmmmVc
IgLXBn4NZqdFwHSr9se6n/HFZTEBNud+S8O2Gs5JbQroP0en4I1JekPpspnc0TDX
rNZYtHyrpIEu+kz2tljapx+bNeaS3DF7sKLr+Du46Pie/CJ1pQZ3N6DamlNHPQXi
6JUMa/zNBo61d7Ki3+oxo+pOc73KeF7O+wa3ZgKx9YCykqv9+QNcr0oYdAm7AUHD
Cs0JDIYqdVPCyRF2d6RXuzwAKP+TwdS/rBMLIczORYdDpmOVa5EBS0RewrLXKcDg
n4+5UJGPpmwA0yorFR8kWzX8DpzLRcEWiQr4W/coxhDqxow5nl9CtdnmSXq+MI2P
kJQoNm1x0QjtVZAZqFqRCiz3aNi0FWIqtvvUg1ysUapjNKc+JSKNsEi3PdxNEp2i
EvGwAFJtzSgRg+Ev+lIoDMUgeF5uXriMEbVl/ZcwSd0bJ4W29De0oTK2a4YbmSU2
WqvlLNpCdZCY6kKjCWXepc6T8F21X1iNfzyZl0YlacquBDATB8H0EzbRxL6nNMLn
RTKFFIjaGvQNu77Mzc5rm8lc2zr9QT6YqjponyUxKC1kzyNbaNC6uoNZ15x2fCXS
AZ6Xm158olCIqWrzuFJn/ErvPMlCPAGo1/ynvVyY3+PjcRwlyG9fuHreT8iV+o92
wdRuoKoDGGKS9ZZfUgGRwhy68J65XPUbFEV4/APKnU4sNAlaY52GaUn3MUTvFvVb
R4yF1GMx7bt5+zgdQ+QhsTVmkCqrpFukZ+9lZA2HVn33qZz/LoUTyILyWU4xmtrx
qZE6FSVRhfW5A9jFLEsKq0aqUdydXGlsdCWXoa7CGIWUYbQUz9cK/bWDWUouWY4o
XpgGROq6AeygpQ1HTWhyrQIgCikQnop71nrNmrVhwNvqoF5Ah+PontQS83rcxTJ0
+YGYpmHwuSYtChdLjBL38zt4qEPmRaEP9QMXeEBjM058B+zn91p1vEdksxn0MrzQ
iD0LBtNhR6lsoVxjvWegCtFKwAfy3M7x4ML5IwxkzQwp3Cz2RzXi+zsGoKhZjkSt
5WLLdxj14YxGXheYm9kylDMGuydeaO18TZozAQMrQihaxku8VoQIeThTqbM6tBPA
cjZgqo0C7KDoWEobloIZjOfp8KHbnJLJNPw0Y46JDdMlsvAeK9diY64CQPJw6l0P
/ItqESFuZwOFVtAT0VKs5wV3/FcwYDoR7fv+PIEW89qRHEwArKet0ZKa5wV+2P63
uL3dmCEICwVZSY1e1RIM20CcYEny1cKSWQLtS5w9uDQwO1Rfvaan55Nk18c+3NzC
7pJF5gBGvsdiEyBTJ+gm3TeE+91WcnMuQXTwY4d1cO5M6Vq8Wabc4WZNyuqC0gwD
lzl2n8vx/BvJma+3qPqaJVAmmiwzaC8l0zBXbWAMd5DLl7wJTUdyDodjOloXJmII
Deqm0/IkRr45eoZpxgRBmfsb00+FhJCd5kNg2Unz/Gt2vy8zXI5rjgbo6SWhtUOT
GL+iVKgHn05s++ytXR1moO+dIaEKWQrP5actJ1DUO3b6Cv7mGmVdCqXYjjbZPpFd
EgQSHGtJDMAU3y/alNCzrDMtdUiE7fBOd4QJMJ9VPhs7sY4Daji2Coo3LA5Shg//
YXh+WzqBkyUxD4KItEoOg0xHCwTPyjiJiFUXJ2tPOXw73c2hqyKzpD9LgxbKfb9N
3yH1901o2X1M4gPnW2VGKxkaQMXI9kEzFnl+/8YhyxEJqxfBIht3Oztpf42bqYrB
8BvJaQ187bErScU+3FQqzNs/Lw0uD+LjWdfabhL1RVYVm3tddObRqvvJMXFiTUrn
uNJMo+rhZZBaNxt3Gl4Dwg5B1FgjYV5LwhpH1gQwlXT4adufnOYsVzNkSeUlEyeP
hDRKl0MlDkJ3gwCi7NtI8e/23zKXBdRKoRg7LtEnxdYC0HjMh+KyZChuJUnnk3bc
Za7yqsWT7LUOSmOY9i7aHHFLv6iWtp6ItSTXGukyAVqT+f5qeGfQABuVho/6TsPD
LTOjlhnRHKEzlRXhz2KsRUThzd2FPjk1DFdZSwD8XkfPKz9rMQSKiVvpKupJ1PWR
V+34+B0NWeRNXWJmtKWn1oWDY3sfYdfz+o2JStw27eUYvsY6TIxyR1Y1gsvuk+47
Q3YIt6Z1EskTdNpDe7x/87+5dRNeWBSnn6vGWH0F1mRdGBq7Kf3uNd6RwS2VlaOE
rG2N7MAcq9Tmom+hu8OvysnXfd880m0tZqS9EQ8vmII7moEjr1OgyXcmXyDWckel
K7vvPS/3Cwepn7hefjMzrpH54XfdY6cPiz45cv3YkAQ7K/UC+lBpsVDnScVDnBrT
gUNol6ndHx3KDiH3MbRiXdTS9hFuVcj5dUT0RBMC5bCGvfa4r3Tdu13Mp6EzetpG
Pm7Tq9qzQaCpbkIi3EEil8lhg3l6j2wpW1BzDYu0pxEVjTI1GyX4hnBOBr53YUGD
l5sznvU0FCCXEsFW8LCH2dk8cTMurV8+aMVJSvIG9XuBK8r1vSqYuQrHz6+nrrbX
kQLtKDnQgpWDfh5JTLfONBT9gn/5e5PtsmmmLkOdhtnSNz6L2geVk0tr6unLOnmu
XzyyRbaKP0dLFMyNfZYFQ3ghscWXqXZmMnUbN1uitBhjdpIhDcy19Jw4XKiPa5t7
nZ48ovMDmJmajbHuQ652/6fFiQeijOvW/QcEi9Fg5PU0BMxLArto2QNo+9NS4l0l
sLRxzjorurPiFocH4xKKTJc/H1qMUjnM4yCHPvd5h2KFf42F3jX6qtUfDNScX1Pj
UCwIKJv+nIf/bkKkYma0xQ9eMCMsH9UvP3sDfzC6/KhmXx0zmAeYk1nCDIaBYcNK
NvnC4OEcLoKClRakiQUt0KMlMOctIRVUeCpdB67xxGxYQJzUmASyfOnIijntxQow
ytYt5cyKEYOz+jaxncEmO5j8Fy5AueMo+zqsk6qtEVwXdBpNE785Zvxw1JeEowOR
1cOsL0yUQQkZTJPzG3iNPWZQUw9xJ7aTnuyU0nTQQJ0P3qNFRcYAmgqaNFpXsupa
t4i7O7/hq8DB69THN3HfGDMIH5PolA9DBGQkfaDamLZGDlg11TcUZuyBkWpUwCoK
drT7R2biOhsOVHIcyX2Harz6djo+qN342JruqnuR4ZPrz6cz8wYT8usNtYQ0HSP6
yN77KkHLdOxNa0QiKtAeeocunnWMH4J49QPlEflZGID1MHeoeLaIojG1PXvsytsq
ZrxRiTxRyctakjPVD3eMllZXcKrCXbP2azqlWsAtDtviRmfu+JapdzMsT7X9c9GB
DDH66tu7ef1kZ+iCxl2e0lFa60uP9MCPPiEy6VEfRjHiCUq0nwj8XFnHSPXzwuWc
95t00302fb1MgTDGf+FQNZJhIWl06G9rTysOfkX89KM1SmPR+UNGOrXPay532LNT
qPxCsi/1swb4IsVDbqw1qoqrFYvyZ6alpLM9GfsTN+YxqeAxTN4AhR/9LAPx2IAc
BGIMmumovSHfO1Sdw3/8Tl723PJsI4Ws0gm3mapp65+xS7EGGqLzOy5TD/D/cOe8
G9ffzqW2V/r9rmWc/F6uIrf3fwUwbJGpl/Gqumj/bHCAc//e1aqXhGnjcJruOo/V
JScveE9PXltNtGk9NfshH3IZhlPSS31TbivU7gU2w+zoidIX8GioRmpH6MbhymQw
TfwQKo1urJNCUTxfnSzx9pPt2j3bk+vDsyBJ0giPPVyIJ/F8CiPA3E0csguqvX5C
pw79X3g8uJFlocyIzszn4nVwhogK9L1qHAUEtlLp0kYhdX/oioVN4XflB1GgIt36
B8+n9wv9yRho0JCXiiFeXc2iF5Fz8orixwSxakU8ZfcmEsJiWk4adHGIfCwhU30/
mAL22+dUVBMeZlDP2dTweaJjp3MuSwh9bwEoxCzy83RFbPNyIYqTIB7dCx7mbAh7
a5NBpbW/hhoEkLtanjjQEjMzgC1VIkXXaxUZYAbXvTXF+ImFXsSEj7aBHGtJJoH8
mnzoWXOKSIGWaWgdmy8IpmBHECznR+yJANyl+ltCUcR8MztJn1dyzbj+IK/8t9p3
A8TJOgpZUjHYtdjAJgEy0evnkSABvSb5HlZ5y+/OBbf21CrSNYxTJDTojcUmec8K
M9y/1LNl2pGaNuLsK5eheU2ewY4jxZhNyQzA9hQIKPKKd35BEvUBVmmUD2aWnld8
gm3ZkdFexCHvPS+LFVJ/BQ+8vx7SERFEsjVqCTxOzguLYEl+AkChPx5oko3fmsbD
RH23Kw0L754x6mHZZpiQugq5XwINelnXToIuh+noS29duAE/Zt8VIRDruqx61QrQ
yLOJowAsDAJ8Cpuo7lI2X7pW6/doRrG05jev2dbSZZ2gL1+dDKrC8uktGhfAG7Uf
upZ5pdj6+nWavO3gjPEPq6r7LLseQfShCLPR2nEVPxcKx/dRR4MSpQgE7Fscsb0K
fyr8Apy9cUfZ4hvPn4sQhLCAVdOwq3qsIPYIGAbP3Z7b0wgTgbat6yOSZ8bdYb7V
Z8KgpHPxYp1b9aWXCfrKevti6XF1GjJCQMCiDrbYDz0e0dVeQmCu4OSG6+xtb62M
OEAgoUn3oChCISdyExWJBbOr/1D36KaBb7P1kXRDjzYaFZLc6pUAzo9pto662gdL
e3MxW4zIf46xSncwyLv5/7ac/oq0WwKX3z8zMTSzsncc+0JZZmAbHV2LOVNnaRpM
hT7mJzjgbWXHekgitJ45JTIe8VhVTe6e9tNTCGU4xTtcHrwOnEHLh4Yt3cQ8TAK8
HFlxp4oJzzoHt/qSTUz/8mSKckFpdCAvWamrYuU1A7lB7UpciZrbeV1PDvRF+e49
er2r5XS0YIWyrp9eUVi3FakJjT+VZ1dEsyjHXV/eThNwmw5W18MR56eVlh31BzmK
czBJg4I0sEWG9sqO/dVTwkX3ZL4Trk3XkZFVSQRq0ZkWAHlhlYlsBCjtzSD7Ql/W
nFIDDJZ/Q7dgRIYlZ2BeI7kYa7hfDKYJdAQgScnZSyqvJ+j73OAVqgEOIKx5MpyK
MBDvv0Sq08UOQvls/aImHFoaA8LKksRCPwFwOGB3/cebKlyPeJe1cvFX5egnKhR3
KzjUepmq3N2AU3KKgDYMlso0UPNhB40JIXmMjnK73XYIx0IWVDoAWo7IjNg4TBEO
8K3FtU63Fq48DFZ4k3K65T8xWPM0Fy+sSRFTbL5LgwSEtlYEPlDBKdzRZkPLqRGK
3Uq0lOf5x7EkV7zuRKauaXdZ/cBgoUj9ojUx27ZsnOOYCyex6MGv0mKhTTPkDzuD
DWQqcdV0Bpqg/GeFvp9Obw6Wn7m4IsAPeoOrU3nkqNkj4MfacXNmQlPJEAdiX4Os
GRyfC1+7wBm+XlX/fg4fWkoT9AYwHg5aHoiKoW5ErFD5cj4sm+hRr20SKYNLtu/L
mvxd8h+AUwhU/TpUJrVCHfOsLe5WoZ7xP9T59h41RqfYrLJ1MvDIFc3bK960E2II
ljwpTMSX/iIjuFH4bmCmF1VGHSZ4vSJZojZuX2EK7vDm8EojcXOxh4As0I7pv4C0
mliXa9m+HuE/OLz7yk4whc/9paVb/jEA47NMQjU55OBMZbr/ME1/Q3+NHwhIM75f
vFOs1Q8NpjuBEpHdEuwt2FOyF5BsIMYELKF+plriMr45PX4PiCgvfN/IbqYOzTNy
3sHTvfZI56oKdl+6GyH4fJuO2ardRFeJblwcr2GSbNXT19Xn6vwQgmOG1xPyp/sM
gXt0+EcK5MX8I8oNp6YPxundaFnCBIRFukQWNTsZGz4lZ/0go310KjIxHhDszTBh
OnWIvSHMyclbb1o/JXxUHpBTkEBO1rDIvyEmRX2Yv/FdkwpiPsPourz2sy7L5CeI
2wt/lMee7iqU4PF9+DJDH4y46VCKBQyOcmk4XBPplhaLjX1W4G5FMg/dWM4m2zNN
qwkM3YWvTXCMOI9ZnTo2zdXSIXhXy3Kr1WyeXRbOm09iLj3HCBQ3SOxOfKwx1JkE
x/xrAQXbpAL9byqZvUDbX/o/QY2WNqIZZ8liu6QhuVFPdAUlwg872aRIqkqphzXX
+WJRr50AKuNkOE/xHvsW2vWgs+Sauj8MFMyuW9WsbJ277p9uVHPlxwvhdox3BrQ/
2CezeUk3CAuVgqeI5rCQaGc0yIzyNeMCoSvUsFC48deL38R1Bf9Qdzear+ymvCKS
ZD2PCK9A901BR3oVzprPmO143MJaLxEqQdVSFf0i2WHGFCxzLh4evMUo4dn0tAZe
zP/MEQKkRdRcmGuqHjjqEHQnzt1mKrSTFFc9eYihUM043uyqNeuZPpPGPSj1s3HS
82aB60NVt4HjBndnDYvDvM/Gedd/z+M96g4KHbghNGCHrDiptis9vT5Pq2rw4roA
3PkAJZ1WfeDzQTS3f3WB43TBXffrkpHkA1j2BRp+SLztBkIuqFRQt/EeQliBdCIG
GXhlt5WMSXRKsurVm1OW+R35mMYu2QHH/DeR90NKTzjyLGB1fEH5ZccDYdVvg/Xc
HR6mE2nP7BKQdQHEoQYIra3oCC13MVG3B8z5NcW5GJgk3msZOQ0CZdiE6wzqxKwQ
YEKmZQ4fO9FpnWG7KJtW5i9sHUlzNvdNO32nfHcVHy6H4HklKNoZkBGiuXKVbLW+
gpnuCn3FpiGO66unVxJeXm9h7HEWfw3muwKPfqf8HqF85nU7Nz/kISW6xVLm8nMD
Cea9WdAfNVxuKK4k2qmMLT+pa+bVDuAAMqoG4Mf5Z34IlZ2dr/IDnA5XC/CWQsUC
pr4IKUq3sXExlsSaz9tsZDjMGRdNiwrBYC45JnL/R8Cmc/19cvJn70e290VgcCaF
bigvttnxC91p90cH27ay7rhNnDnPOxECpDid+kpD9lZpRLEZP5f/18BV5BwUKwVk
/rL8olZufIGFxcXY5Q1SLmUHtiOGv6xVhrvZm5PsCLcVykIpdHp8DT5rZUvxq0zM
l6pSZrURM1msi7hP+tNucedRY+oAEAHUekn/lhzKuV1AswpTDvX8BYrVPpx3yqPj
nom6DpvnIpRcAuW28gBhEwAQJMwraQimarFHGs8MO9nCSDR/pINlUbufl3FNkHr7
AH3yZVNEiSJgtB7Y/oewNk4GI73K7lopmHXnnI079qQx2z3mZzOjQCcsdR+EZnJA
THbKY5al5BNXDzDoyh2CRzJFY7cVlj1usZ/gWQNXDYD6OKgeeQ73acA87mjy19sw
3jBbSB4XVY4uGpGKuOfYyiNN9OCab8QXochcvLBxaavhoruPwlIOMO0zSExGU6Gi
dw8EolUOUEdbBwKIbetP75VGiShTmp1Gu67DaOM1MEfkzdJeX4TU+/+vQ6h4Y+iF
r8SXTZvZq++/KUeJpidr9AcU6yZP7Fq+SgbNt3C8im4cK3zX2VmG7O5hJVNhDXM1
YxNo7tOzPyajqYl8e0NlS8i+wu+1Q7oKSHmyhHa4GdrPaPXPoG1PPKj37w9lY+7Q
mV+L4NOIyAU7f+FFRT/4iOLyoyPVn49Hf/M32rkbVd8L7E9segnfA4z+jRO+iewQ
bd9WkZbk8s0B6+0U6meXV0hm4XxMXcAa0rrw/J54/aHS6CUWNHcS7n50zHrFqPHr
ceXlCAFziGnFhkim0dnR1ZA20MTQ2oUL4MqR39iPBeQmux+00oqyLqJISv/3Gt6+
fAv6eNd/610D/w8GA/hIeDa6nhYLqMDVSfbcHuyEINcrhf2yIxn1d+EU1g1bnvjk
glbHZy8845/zaLfMK6A0zkLCwmqSI3PXxmXdSoHjb7BvhGhGHA5L6clAkr+DM0fr
tNogXpM4q33f9YPDDJ/VfThTPbSSScDe+Y1molpJc1WvVdrN9H/sQ4p7vHrEo7Pf
qXHi+AoV9NebjkctuM808QAxOz7KBR2UeoXe5lmfMqkon+UPwp4sUEqvRyS2ORTI
8N9+P4AXQAU80vaKF5CtDaLa6au44OPfJ/m2N03aeYGKreN8G64bY04lp/uin95Q
3arU19vh8KRdfsqftnqjBnd+YHfFRLcaEFoQAdughZLPreszjxOnjcmIb8ygqOi4
McddJZc3A9EoIKB58/j3svE2hj7dxvD3RwV+MBoQcTr3DYSTtvGqOsfn6oWKN/rx
IvzDg41BYYIrMCWq4TWh/TkFFkdZk0BATp+zjtw0o+ekSNo5aUjZmaRtRmh5kBDS
cKHUe13FTd6R0JlC04MPsqL/PYyy4Eb9reBb9n4vWoVkULt8ws83sJrbGB9TR1mE
SG4360Uq/2nflinWVmabvuljs1mWvhsOj4GMHMnfqFxs2eZTyozXV5OKT3eCPXRU
dEIQrOgvL69efdYs8V5yBnZUAMbhatoVKlvRvpvCW4smP8JDI9Qz8SlVZys/13Om
H5WZGF9PztX192izyPn84JdbPnJZ9LWBd3VsaAzroPeIJXOsYHYgSt1japQkD54I
ztFL/G8DsUFWhkIIDYqkrPrUdhlw+li0huXr0Z+bgvAxpdk5oqzjw0Nku7Mzw9Uz
Vw8tC0oKVv4VcHc01rI1jv3mJUII0ebxHtXLkUd08OrWFtMDBmapR9pWu8xJGxcz
y8xXeTpNxPWRiZcdVJ5OnlWBBPPIZ5cDiMKIC14HHnI/awjdAOLpYW7KUrZgm4lI
YFUUCO9+lGDAYEdV4XwP6MHsPrTNGwbaV0ooaWQU2tcC8Iad3jIoN85o8EtuafFv
GN1MToQLomIL2u00ijKPN6eoTx1fOJ/k15VyVmW8xoLYrptpi9WY8LFMUMTf1UNL
+krR22uL1EE7N8cpw3ss7PKtd05mJ5WHe15QAGp3cRdlY5JTgCPtgu0GWbr1QFgF
e1HgGfkXl65VVKE3aipckdlp70BekLorDx3DAtxiYZUEFuNs6NIFKZ2DOskv9QZh
NA8y0wC3aMBU5ZbLwiK+vkzK+G8u+L56cWHj6qF5yZmiOA3/0uyTel7W0rMfYMJH
v2C1Vz2fF9Wb3ADw5chJ5omQn+klorNpy4n24mrJuyebAXMl60iRA6saJxQ5qnDf
eIjN7V8imaCCWKG14+H4ybFms8YFYWaGLVjPBBevQn1eOY1LrxxDqU4zke54lPnQ
GSqPFNIpe4So+SZsqY2jLv6WeViQqYc9ZIg7jPyl18FHuahQx6j4uWYxv3McT0U9
ZHZtt5ZBK8dhk3qRL8WsiIIccR9A/yZDkaHZ8HeBt3hqup9R6IDRFVs2coepvK6j
OyGDaM196mjt+Qr+G58a0P3MHwPILSVeoVZq6jb5S2jbYtmrM241sjzrjWnpSSML
tJH85ilsB52jcrVP6Jrkxonvgyg4OIJFFCxCgPQ9xV1srPzrQGLy5ijm55qXTdVA
Lq1WEowpsNC2jEtay9bexJQkA3o9DeRAuuilSicwLhI5if55E1UrxSNFjlNcZLiF
7q1sjlUcErbLbollJNWqFQx6Pp51i7ef39lllJMS8rhB3iehIJ8KzYLu190uplKt
I23Mjc3bwnp838i0K8hck/RF2fCZgqLESW83DGAqP9nLefnm5m3uC6VsO0MOGTPI
kmRPlhnRwcPakgWMS9pKUDAznqUze+EBzIBPxevsatFKrEVMIn3dx/s0EEC0EpJs
zyrrBu4cAvM8TgPaZDmOU0EvLe8rsawdk7R9YkCeAQtrkd+wCDASZubWFYgnAeMz
gDaRLfWbMh60yu3qdXAkfPfDwWQCI1k+VWOm7KvI/QyZ3oJuX6CpQ9aS+DBR2IF0
q9elhLEYjCL+BPBIr+/SsDj+ZpRrWjLEpSAFF9R3TAFL4ps4Qli4OQ9Wnqc3qc8u
2t9uPy+lyY1jRwu1GZu7M/p5Im1/z9namW4h3otKbx9WI8xUO87aL5SSpNmKwV+P
OI2exCWCJIEe2s5+RF1kqXfhDIC5P244J5RWwhFVViMcpwG3tm5WCebW4c9hbb7t
1YawQlBVN7pAbyGVBAnnPOlvoiz9Z7OKPqIHXyKaqBpKhjdAY8M1CgRRYZZP3rDa
Fy1nPKzVEAKmwO9UQf88fkL3O6sQ5Ap0iYRXiENVoOuquqggqL4WC3Teq6g6E+Qu
XWREsW3fYN27K40p153x0DYZnGIh1nkMflh8gw/OBIG11ioVi4l7O5M9C+zIli98
4le/Ph4sFqhSz/N25APcI+4Qu10dDR4aDoYDnApLXS8vAY/5yIUaZ2Nx5e5S4k5w
Kyw9cT+F1PedD2tYhA4ONjHqO8MnOBFK2xZAn11U8xD5fGwKwug3mH3EFFt+4h5a
Fp6DdF9FaB0HTv5i6rcpx/eRu+q/FlzhOHRXI6f57c6ybY79lxpSKXDbeiVXft36
uguaecQtzFKnk2gHpyhcNmwvt+iSeQaL+84aQc/nOsqKNJt15klPu68G0RO02oNS
xewVmvAxZq5ieAei+6Tpm66tFHsVEC+SGy3DWTd9cYy/fgMFOou6yDws3IWZ2e0D
Clh1mgyWIVTZ7HV1XaUBr6cRXecta3Ktn9MkDlQvAwNioPzjm/XaJBCfXL/ZIDwi
KYuDzPfzex7rhz0oLAneHtCwhUNvGEZd7wi6PUsIqhyK40xL4cZowexpoFQwEn/R
RDe3gf2qSavytoBDOxddZKdEqEDPSpQvgcwUGZRlCL6cIZZeZVc1ghKj4ZGSkacq
Y200w17b1YQXGrZ8DkOnVyQTvy4rm1MLihQ1HC3/CCDebjK0CEnXaeGVPuJMup1m
+hFhyUy09pJvtzvZuPmkVaxTXNGXXycBWYeUArjKHgE0HYstuJc412FPTTN+rkGe
zSFEpD/Cw1U+5wEhsmxLoqF6ydzicCfPzDc4eoT9HHFYYNppEKXbWOXZ4Pwm3Tmi
AUh+60LwfKogKIH+LbYVUwjiWu58d9b7JVSnx8dPvauSSaKYHQZXGHdZIGEsvKJs
dlyjrXPnwgMb6OLIMaSFmEL5eLivl12EEl+Vfew8x0k4mqOrNTtqA9MN2Qzjo02i
nLvsi4fjOn4B8O0vEV0Zq0mRlrHJXs+ssqKbT2oORoLkfyqljaKoPqWSCyu/6kLp
NoFbVeCQZHeS1J9EmmYxf8qBtfVRieIULLJw90pwcqnKM6nPyT+H1a34WZMTSLNf
nsc/v25B6YFAxmsebPz7DRSBPoitrqokbDUAihOmO4HKoyaTw64yg4sxDScUNHvY
11gNX7UDc4NoFQV6Zcu2HdfYKpuXB3B+eVZQkgG+1v32/JoWbTSVcSUwT6L4nISw
Z2gS9v6EuCkXVMrkqWd1fQ4sdwMHZEUC0JQ+WFYJwVioTXcSekqo6Mw0UjK4n89E
skdyTC+wyEduQdlrUfwtHDsWQvaWOPRltzLz59qz7bBfGHI1psQvMWWPKrOGTMrZ
RyAPVkO5gFttlldVgEG4FUlWFwYhrXhjzl+c6u6OMrLqL+/pp5dxaXfakBg7bwQL
6y92nwMSwLDWcFQkI+CM8Sc7QZYNEsyxvWMZLQbx7vB1j7U+jTo4QMG6OHRlu3aw
4xIue5v+84RwpBe3TFZuvKZSUQExuNtxKyZoqr+iknmdo5SvRdo5aFCspod6g7lE
fF6z0ORcUSzlstwzvqc3gDrYT+FD/iNeFRSNSMtNq3Lm1z9lFTXTQ3rZasAD7BXS
Jxd8/Htn4N5HJZrHseOOvtL/dFGtxZCfpkdbThBWn/ZUvVs2eyaqx9OvgrQDf5br
w/TwgkBhzle1psRO/WAPAjgaUvkt3Ks08hTOtUGAzwmBwlgz8R7gF9frc81eP0sF
MkWKy6CLhraxlBb/1DDbjc/m2LkbK00YVcLcl7HLymjYNqD8zQxxN29SWTYdqNWo
f1yOV9IiaAgGIBzYUK7PMMe5iHduOVYtZgHEMY5G5wM3ijumBtN2H1+tcGGU3QvC
EGhhnzYTDaex5z9Ewv4BBiTEb2gstzs9VZ3uiTzK8Yb0NiMmM6mAr8sseX9lenF6
kFFbxbhRNkRDNocTqFvgASwJrVK1n41WZn83YF+2HXiozTtVHETHvml5wFHIfsBc
0oqbDfWApsmVYRe1QT/eEo9G8ZQPWkl87sQaQXswKSsa69lZzj1u7H46kukH7poS
y24KfYQCsQVAvodDy2Bi1/3uPvxeewXdKSWWIR+XXR4HCmrIWuG4XxkNy4u4l7kb
6hqi84MYR1DYmR8TTFT8gCyX3dx5NRztJ0COZMBH+LRiEW+mdAcSbxgrhlWTHg0X
/5sBUqBzZ7PnUwKb4foAf0CzKtuwmCOLDrb0+WolCrLjzSjMLk9J34a0/q8kpj1k
3iI/zSQNmrKC3Yqzkhu0o9iAxQFg6o/mMPXUfoORpvPjcTL1MocWTVt1dvN7Ev2d
MkU0I+0xMNAFjQ92UeoMCFXSQ9wFHa1eIzdR1tKk/6ZlBpUBLaN9dGOG86OnxXRy
INyz6TVfPvHup9w3C5MWjDwh1g3pQA+xIfZHixOjqUWBLf2bjqIyfxlP5n46kEc7
8Lv/HipZYTlBA3foihnPWx9g9pkejrtWxxj88OkfDQCQyULYWkwN0VNa8j2pD0zH
RR9/wdEZA3Jw8UBAiS3vbg6NJeDHGEWwJyp2zY5hq3UKi9/nyOGin1uXXQ3RkDsc
UolAOE7QU6xH3JfWBsZLGxoZDrILG4Pl5wU2OFjAD1WTlL9Lqdlf4tREcZu3lMoN
h53aIywRhXJxyc9T0wwHa3wNhX8Hfad08V6o3HMWNz6tLXH8Xx1BLK34IdN0viaK
LCgoF3oUAW1xd8mZRMuJrBSSOcJk+6/bJTRlfL0BmDNJ2gGG0jZEgjpIDxvJzfao
h6KoYXsi/NxjNQOarqD8lGpMGcknpGm1ZPl8t+sJSgGgeBssKypHE95x4bEe7b02
LbdslwQx4v6YQfKf6ALI54cYIYUCp5skRcf9q04uiwb8/HzAGc/1CPTlheWaWvHI
y9gI5YzEisuM48oqzGdH26ZPu3OXDhnIoZcjzBatRXInKa7m/Zx/uVps8wniIPoY
SJpca2qTJbFnLrJ/vYvmpstgVLna9gegCiw0AaZV+K1TIMIVLdj8sGLO2JXH7r9l
IHIXEg87Nhi68rz++LoqJ9OlyVHDLC4LwLA3sW+jlCAVdVex9lLswG/CqKkYc3xy
bNTJ0MQb/JRltnPTOpxkgktX5VFVeSYhEcHMBrcOKDLJqtEnN6+ftVWxnZPN2Od1
UPwiLEFofpPCExwF59h7fe+0tCKEX1cQMUSsSoHKQp01yC3a7cINq4CkUPzV+V0D
WLRPZN239ZqRhJLBTpNDrhOSZQgTXvellArVvz4XR6IWhcamdUpHIz3ySbREQapS
PTl5F84cz8uxgRvFj15IerB928iA6TxQrmXzwBguk92eCUdIQ9Xs7VzZAVKgCkVb
uLyfNBtOERFWfnZk5m2I4WEhueTYYIIFU0XcN7KZXMDJcC9k9ZMungHhNUwkYokz
gIPM80tbOhhLWbZXZbnXqAOwSM3lXfiAHbIwhVS92wbSCHdnjPm4rsLC9DgbbwZn
E17YjQyTViyFOcy89kJbjXCbUdD75MUAihhnn7tLw7P2KcydjRgpMXXJCtB5GKu2
pN/vs6MmbeCxhEDjlo+aNuZzQKOiG2M50bwCDIKRGsRl9rlSGghF1S3kO/BPmhQi
fPncHrwo+t9Shh2mmJFvi9/v8v5e8TFCYqa0s2B7l7Ouh2OgAKey9TFQEyQMZsDw
vZvhAmAHA10fz9yMI/XgUfN8ILvmqYvI6KmjoW28UWDqK+9bPiBTVnpD+2B7h48x
ON8rA2iAaSNmPHrdIDuxj5VCM2t6IHwn/KjLGSYaHIsU7CU3fWSokETfaBPAlRL9
/Rmtwc4d/XxXRuhWyGwAf/4bE0magH1M0lJxJh9+FX9PMnE2H4/W0oTsaCwOELM8
/wnA1zfRY8AorJuW9O/qi29pRW8JZWjSvJ1v7V+TK/aVKmKRkh/VG37DaH5Byog/
CVIK50+ofhn3jfXOuZcEUlu7/9Ab32OmHiIMTj5Lhj6+df+dscXXmKVXrmarX6to
wjnvDuB4QxeljPxKZS5VzduxQPWiJ1QXzpiLUyiEs+5sdRYpCq4/Qp3ZG0qZ8vXb
Qe+aFxhk6+G2jnzvC9x/vjqcUVrSnkKlPzOcDAH8zJAZ3/BpncCJCScWI+MDCIIA
5BCcsB6LdEuU2pX3HQz3jdWR4EXErELHr43fpQXPUDjCqk6xjSEh0MDv/lBoXQiA
2J3UT5ybquINaMEJvazUHY7PzMoY00hviTNxEJu+E1iB1e6EtvjI/Y5EyXxTEDzX
BImvRTvxbi643JMtvMM/3a9eOFgNgdouqDPV+wRlfBRJtYB8iB8jNoPuKKyGCfVB
l+/l6JVHnM8wQt7cUzoNHPerqHWfAkKrepMOTxjbcYFdZLHC0yYtreOgOmj3EqyW
+4bOLVo8urC92Bo5gjFNLH8F5Ch/Le3erSnfnWJoZ4l+ba+EGM6bC98M4VdhEMjp
kSz6NNmHCEIrOL7zyqkZF/oEAKkKuO8mvjYitwpVKoIdiC2pFpDx7+Km2xcJh2iJ
ErSU9gA8tTIQM0WmfVU8aFAUpkdIusuJy+RPF/MqgSCuGEcWJyZcAu+CnAcZ/224
t1NSh4RKSeJDkr/pckwOIYEM7yx0qt/m8uwSEEO1DTc4rlLlkpGUM7HU/5+8t7xW
nYl4rsiRrZscyPUlVa6NI6HY5FCUtg+qHczcwqMcm3hFWlbQbt3ItZEc7aRYd0e+
Sl+BA5mJ2QFlP5FrQUaH+AK2y1yaYRJC7UTm0fVqTgY0QhvMCNYQINuyVeATcfua
i3LN7BhDldyY7HelhOXWpu+uMXlME3rbM06RpZWk3GCc0oETz8aXLQjAETPLtQIP
cnDyMj/pGE7QdpjpRYz81IizWEnHDBWS9iuAJdJ36CeZdOyDaNTmx2wdLFwrxQk4
giLhbRriIpypTdOyDhU0CwFDz5kBdMqU3ju9qMdMrAVt2cKvnaJkf4S6JFivaFz9
ZSQdTnxUFiLFyzlFOByYyMZ5iX2o+pNGJ2T/Zzsb/xlQR5bGaIJS2YPgswSbVyXo
+tCEyUDlIkMYLcxI546BTvKD1/gRymCrupd4aU4JJaLfKxe6RLIdchMysKeLy4hY
nMTcrDWBY6crLUaRk0ZfLGQRyStb594JE32WlQMirinFuI8WrG8OZlw50AC9WNig
jw/wlL2DQUMomLbCdVtXW7uhsV2d8O/YqHj1nw70mZ8oGAwLOX2xKugAusAb6P+A
3KNc0Wne9lMC/H4CdaYLxUWPftmyoVJTBPNgNNpvnoXN+Ds8IDpjGmsvLrSwdH4Y
RN9HxnvSp4pbY3lqRVasfBdvOHFXcEwVozVNbqFS/azHIJtE/gjUvauvmx0n6cmy
MC7j5UYipYVwBJmLlrTRB9GJCmBj5r4Z6qzgRZT1iZtYDVBXj2BkrkeKPPkANjdS
M+UayzWskKlbkEGUFGeo0RjqI+jcIEW4AR/ObruVx0GieSLCz6otMXFnb+HznCD6
Tm2ZpP3tsCAbdGzTT9tAuiXQF/4xu3PwKDJL1PJFdUWixmk+ZOyz/J3dlZn3psFf
EWD4aQ7cjuL53ixpWHNGVNHRdcieT3HjWX/n0mD8aHNDPbYNfNh6jKzWpghEHQu6
3VjvO8YP9QBkERsfSzQtsJQJ/e2rwlCjIiNBMheS0VKlAmp2Bq9cwrPjkXrCBBzW
nBkaZj9r1fCBx4YQssD2Ofp8CHZ8orPNv2N8Zo391SdloOUAfy4lUUM+5iikMuxu
lFKrDVQ9fowE1KtvG974ndKR4wbTTyFNkeWVRoztof3SsLd5j3LOyOVWie1iC6N7
oHk+YF5kcBATRmI+TASTwEW5lFPmhwvlp6SGeNb5JDsCDYNdHGEJ3hHQn7BSeuEQ
kuhAy3Jf8qTJ4wLqrpY70j5lcUkYfbMcvvr28jB7xbLrLPgzwfeDmWeVenf5QT94
fo+F+rQWI/xXicnKsxiniEdlyihTW1iM/QD3+7sR700Cq8RPDS0Obtl4Hu2zxNCF
sif9dZMXbBGH4xyoBHVGc8jqVP+RiffiWgwCaj422O4ejT3loxx35HL9HFxpAB8p
DXgUATtcZPq5ql7CQbjkGff9JWyG1w2sCiRrmt4fu/nmRXsGfEWxxc4FVc1bcPBT
kuh1UmZCtCyrRej3KqKhydJHpV/xui0NgcgWA6iYbaor8yP3OG357W4m3BIAAMR6
n3e6DG1IhwZ9dSj86bN31gFTnudfS3nXQ9vSTWZgAYdSswdlbMusT5D/Nq2dh2HY
ikRnkRqWCb8Jzcjy/Bxww+JlldX9u3w03pCjtasQJBZhROe9pxOmhXSyhef0JolZ
VN7Mls0an/C0qEH881vhsXnd/4eSlx6J6p+foNLh1orbPH/jIsSTVarMayWWSxK/
T4IpOYvoC8PryiOJ5s+LaQaDAYccwy9qveypOgJN9yxBStrvydifl2LN+GOCOwyk
xuMccWTmawOM3vlYdFz8HqcfbbfAn2VNYVw83qx86FDrGZk0AD5su/LOAfMeGb+W
Gm3vVtY1TmcSibrkRGuckDT2g21jDki74sSLrGqRE6g3nha9c25QJbzqYHzHJ6h3
wWeWQpMdl0nQvf0TLkUk12cj38agb0RjQTMA2B/oJzKyvlGJY+1/CusmXbdcgtKg
LGcXX+J1HtAg99fQlb2EEpR+YcQ/U/FyYmNmgS/+saTvMAn4RxmsDAQpoV6b/5en
g1huyh3D3xH+wxejdX+QfDBaQxbb9MeEbF048+t+3aeA+QsFRc76zEfGXHeQi2zv
nwyE14jfbdFthkJ47rL44Y5Wui9wWSdRSu+HXSgHbShXBfzFoi30C7kh1RNe0k2l
PinA9qmsrNJMnyL0Rp5HpXxmnNFJprOrfJ8PxcLpItZ+F6X4Tj9Jdt0vYzfqAQ94
rjrGrAPbHbJtVnVjQcNQArK/idTRh7RcnpAKomdfOpf5tmEz3fzv5nbi/4NKh+zM
SmZ2/VY/adHgqbKccykajAKLwdulxMQAP8NoDMmeQoWO6RkYZecBkwUUsiQfQKMZ
gutAZ7jHcJh6dw0UrQziBywfKTiWLFYdqMuWwEGJI0IKQfhkhANUx3vNhcr8Hsi5
/9zetTRGXi8ue7C4cN2vJixEh+5rimpT5bj9U01LV+TMZCTwVGUoHK11i9Zg6p8r
dxmh5aWLwKWcKFGBxAPHjXoqzjoYOs/ffYRFh4/ZBRe2lmwUrU3bVSfdvE8ZLyoC
AFoEaKA/r+HEND3512BtUsKQUK28wgOYqEjSexjB2SfXsu7Ufnw7F+u3hg3Rmsv/
U0RO4Ojx4cEaqDfwoRzzF+KP+ophM0S5XDzuyKnMqyNRYwGV17jIBkjbCnHlKX4X
JpndTygx08AFTUaeKrJE+b3ZR2qBzyrnVAUJIjo1HxVgEOl2MAOeydf5XPy6wFS1
OEEcjPpxX99kjBdGnw8YxVRan8SXKmHuhBhPDEknH33rBnWnegowInNfHHxRzUqX
vhbT0Pg6H9/qN0FbM/dggKYu/pRGAOzYbh5BepLM0m16YMaZkKTgp7aglwLdB8iy
9zAeZCkWmZRFcfphk17gDhxLjKB7n5+t+3yicCZoxpgJI4DxgxJruSm+Gj3hWLeT
gRZ0IU4TX6/K9Ie0rnwIQaL8IhH9xyc7eHdS/9WUZX8o6NoW2c+LR3QzFycUqzXw
z02YINGxrnDIY/Kop72Ljg8PH9YynjpJxl3eOL27DLQ6U5n/ZO5oUsqPgK4UFmLt
HY1SzwdrOdRNyVMII3toS9rOep/ll0Zjf5VorMErWEVGWzK58rRZZXM0DoojPUJA
mVSL5Mauh7sQ3XEFor2Oxyw/uhP4gIGVM2fzOg8+t+3/2Z8f3vnoZdJAGn+pXxde
rGrcVrMBK9Ko8HHUNFEt2kRPlIHHoOT3p0K6HufREw1eGuvFkYQav7nVVnh4/LrL
ufWTbHPcz+QiA8Dmg4US60m3upASxWWZlfmpMHkUX5sCZ3+EqVV/4XLONG8QqVPw
ZZmC/Pg17JXgmbL9yWuLAp8mdj/dUkQJ+Qe04uD/bVJuQPWGNt28o65NSdR6aGRJ
4/I5Ub2QNbf1Xunz6kSS/y3LijkDMCh5cwew5GG/RYVjX559Q61uYQWvi3Mr17DM
Ig6llTT32ZJ78TRoVGC/MaI6OokXzDUPBO4SRFWmA07bLhsJuUSgFiUBwBiHNMv0
Xot/k4muuDCkwqxBlJCwEWWsSi7XEAIi0Qcvq5TPyoeiFa0wDjrXAyu0NWrtsZyI
3zlksoGBdi7v8N6mhwLHi/GB6sH/bhKuPhrg/hls+nDhZ2zn1xRmR2d2znE3eMRA
Dia2gDe1OrNe7W/t7KqzJH4hIua2DOCuyZ6OmMcpIW4fl4nxbFn/TIo8CzjUUgY+
dK4SznnfsIeJdFYSRhNTs13lCA7pWbMn42orZPCZLDN/4OTBJ/LSaLEAi/ZHU1P+
k/UyGtD10xSNa5G/sxyYyT9fY6c5Q7JuT8MDHc6rCDfcs1mGCXT7VlIJyoz9Enmh
FSwrzBpUsnpvvIsPmbJuuTFAMy6PdhxQqvxbi2bPnFPGJPpqgDa7pxz4JJtlfnzt
JGIyOtqSj2fEeQklQe6kKk/Sxx7lSllminYFSCM/LS9kanY4fYQczd9GiatW7lQY
TlCPbndeIzKkDRyThe6qaN3JF86uU9atCJI+PiWUEJmoXsFK9kWEFZ9m36c4qfL1
mrsVOWJrLSwu+ADtYKqb2X4mOg/vBaSMdCgcnuRBv1cBOcPnBun/gvnDPiCDbBir
qNxiEgbdXUdytsIj8/A/JBKAlZ15HbSPwfopDFJ9W3Asn4C9HfSAapx9KWdna4YI
Zwu5BenaEW3LsKQycrjawbuI7mfB/sVSa9kxd12KJA9cSxTkGui2q552fnoy3Rdx
N/GgqAhzS0g22BbZSY5cBIldskR9EGEzZ2AsOTsrMkVWYQ6DrBXKxSO22HJWZw7P
rshHHhlJPWZ7HWGHj4kyVLWwdM8c2CE6q5AUDqL5WDBf70VM851MzW6AvhPhZOWv
jCtVpLDsUc+7hRXpjOxQQeDf2qRfvf62LFFynVLOPC9nbTXbnGyc1J7tO8pIAmI6
N/gYkDnJAqlGlhuoMEaDtx1EHuw80XNDg6cqADzv+YXwblNE84g2XSx6VztSd+vq
+4FnGbXQRnLS/ALL+yWWR6OSQA865fdQ6lbW9QvYodmjb/EhGMSlbVyDyW6NvF2Q
a57vG/p+u7s0xlAJuEY2kvdtRekI4us3hH4ACIWnk1P9IsTIzFycangTkDCtkTwW
z/6d5NIlB3BQ9YYZPGUQ5IEcms3Fw3rDGR0cRe0RlApZKCTHfTn8onrbg4cSRvNA
CmyLQx231KKzEvZmIWL6Knbnxt6shkhqq194N+YnldURiNs4Jx6OpQ7uvXwgip1y
IpTuJcCHmTpyk+3ZPWUS9jkwEOwsszygmoQBHGHX4j7v2TEvmdW3tYC+liakZTI2
Sly/kDZm0FIIHHppkDqQhouQQXCLOIumZtez9wXL4BSWblivAIcJGU31k4ZZa+CV
F1P56976DdX9q//s0I1jL3rBx/EDw1PkLdlldqwGyVHLNui46OFjeUlujeQ4O9SL
m9/cYphg3F23mqUVKVv/mji+OitjWmKQH4rVYPtNRdw+uZU00smtNytqCKKvgxKL
1aeTdXcLIvLg95XrXCkpb+6r6o1JglpK8NVD61SW9qDb7mjo0RmrKRLK1eYddZAl
QbMPSuJr90DCbGacl5Oi8DVb2e+cyELjE+pYkM9j3rIf3SGNvKyMpnvasW701LCx
QNO6MF9gH2KgC4gwr+8RS0KCqB3SDforEQfbmMX6LLTNfTHi5ocUzA16P/PFgaTX
/k0eNBxNtIiwUL8JoDOYBUxHNcjvaZE3BRJ9/RmiLlpxZgLJt+gzJM2WsiU6tswg
MHa/NmM6QgwYYjPDhJVdxsZx0Jh+Bk1oOaCaCqH7aDv6v0+a9crUS47a7GH11WUU
Zho06Pcri825J74s0IiAHChgSjyUY4DZdMRN5m3f6FaGMjaGl5bhbeR/prjQ92UZ
zF00pBELtC6VY0J2M4vUeOngKcqROlMkn7394w/faIHdVhTDh42ZpJRBNr0tCRO7
0FhfZQ7PtHbRERSjPAvaegHaLbxBMlKpH1d59DJwPdJrVE2GVhoWqxwYfd9UZOoN
vyCfV1uRbdcU3FyQlimMCRMy1CqXNI/bIvRJBup2t82sEHqoX31e41lL2t4pK9FY
Ca4g3zX7NVHitwe3oBG+lJC68m20XDfJLrtVY5/Fz3MAe347RVTwdO8X0HCUOMRt
ZB9q9+jp1PO8ZtrBeffTcRC8AbTiB03JBGrdKGJc3FmZpNp1Hk+awCzuAN4/Vcqq
dD+UGnTR5aV6PUFmXpu89G7z5PRlgKZlKQwp1Rin0FIYsZVb9GVnq3pg7iaKF0r5
kNNDHeoOQwDxzCPETmVYopN2wNU0R4/lFAYb8sB5/TloTFybv/8SJFpR0shZC8NV
3VNW3OrN2y7W0sTemx40DXqaEXM6rJrcY7F6niskkQjp46kXKGZHO2OWXx5Pqvpw
3WNzb2spfH9oHSKrCD37qz5dBIGk3QKaBCnLgWCkJTxGA3m3gbMqTMbaXcIQ7DOf
dgBAZs1GbI36jVRLo5JWY5aVcDZVsElSAtLuljBi8SW8tmeavBF4EJEooUi8yUKh
Q1ylDTUtWK/B4fYSqfio77d5XoAGuTpukuLVyXvZQljxDm64dDkqghoOWpkxkAzm
L8CBxjS5uwR4iVv3e17EW38GppHEI0Ies5/rdKfdveOofXv3NJtLWfEx9GWMy76i
Hp2aZLu3eEaYkU/UB26jMiz56bEfXjTxe6iJCSgg22PthS35GMRDWeQQPhiUjTUr
AsCnsPIx3de96L8VPsem7vUJzaWXv6bB8fxHRX2LOBLKMngXRjuRuKOa2PWaaBGD
ZlILUsD+ob7NlTC0r18AZR3MRqri8NjHFQzAkt53b6/+a0j+oRlX0hom3kqi2IoS
bqmoC9N7EalP20fYD4GSBnYwIfvMT3ytRfU7NdrKYHOEevJqNvLpCdZOFLABmr63
lT1S50rffz0PHhKsRmwsCoqNQipDLHSSicA5Gh1QWqshwIJv9OgD3iz/7GNtxIsp
veUQ6MXpl8rqGbse2x7A7dVuJ8z0LhqOrYU6If3sRtXALRYzmqbQOK+ma9mXo72L
gFoKfSVS3h+/8TWi6UxBkXTYqOXGNJWwL5Y7QQS6bDGfdBzeQBUM3OceeEhhC5H7
eMBgXXF8TpriX76A8ycMeNWgRMKsEgxn1OFV/bN9ZNaKuqmKN1y0D8R348mWSovp
/rz73ldX7bryD/8vKVFnk3mskH+3jxAcqsmszyDYQKOg6p+SAx34yPWY7vyMzyog
jXULx0QzFXhQlZQDZZwgBjxWRCrcrzlCoLBvAj3cnxnUOWHa1SHlPPidsXWrziF3
2U7AkN0r7Lckv5dTBKtFMdaBC2Lp1vfHCao3iBMIruXjqLiVnqV5rKadn87b2SeV
ti60Kb/bmMs4XEVKy1y5E+sZcLTt1nb2ORkQ95glPXyRv6EYkKYjIUuvUL4Qojad
8PXTnuNYO7tc7ow59+TNamuLNlF1aZPF0ha8J2d1oYwxfcoufg1ZXAm75N3AonzW
YPKg/ZznTajCm9JyKVbd87bkc5H7h1uwPtxho4/9ildMmoPKMHWDUMRXVBEYghAU
XIo2upz9IH+xPp2kUFmg5eVSaV80RVMlxRtOwBvNmPxewZCZzWed7lcyKuwQppRu
I4T6eVScXtOLBSiAhOo0/WHIX47QTw8v1OWcP6XtPAaisn3CU9DpvHGnAKaLp469
VlTVyLW1sHPlvQIPPvMOFOXpoc+t2q9w6dNTRFTxou7FPFGQjXC57IqXLGapzFjA
bk0Dv4QbBCcFBE3pYknPt1obmxE9bGL5GrLY7JGnGRhSLeNY3q1cWCyay33jayTD
f1ojXuGaZIz2+b6Uyp+/6cgqVufRe7HEomhHTyEH4lpGN1ezIM1qpoGAvHD9mfrM
QNypPUr1/dYkzr0ucinlENrvS1ERac+NFaxwi4ItK6px6EDTigNOo+JDY6RvzpDJ
Y9BPZIcnsCZeLUuD0IieP1AeeOGGDOxtFamy/t0a6iMBBs1s2YzYTtyc4+8LKgOG
UIx45uWYi1bJGpcDxo1/JkI4p3Ovjvkk6fvui/oTsSWvYfuZIwKJxzJUqGmUB9qJ
mtdTNPFy+UBmQqnJwIdQJRQ8yrXDUtOLq2BsmFli6DcYlATnW2OenNxyrOGzkwGA
XHa0qkWNXn25QRCDY4KuPYWJqnDeZdMkMdyCxQyIfdSW1+zE5/qdr0GAeJq1CQgq
Y1jD86FkDiIDhoLgZF+pkemW7xIha3tnNIKSahK3nGam7d6vLfhIGWtdVajHknDW
S2pD32JqwM/vdqM/YHGIIlkeOQhWcCIbDjy+kCKuyayJoLSESDQl3VqWi2xJMrHd
oLR/yKVSJL6lZW5eTGaOlwjZu2Lo7jvPqdACkBTaIp4LhWwMD4u08iyaGglhwbwz
TCNCIs/xmsihWykXnOobJk4P+5OIyKU66LEGPWlAZnRfeIYT5jIZDEwO2w+9HXy+
ZyMw2/HyOBGLpeWDzofkdVUKQxpX25esAk+2TlKcUMQhb7rfZfxPhJFkV2HetD0+
X/dX4mua8v+PFbMSDra93He5UkCWr04PcjivqySMdtYSwC8pRejX0hELbG9j5g02
FcqXmIIL1zfkM4MNWWBvkzuV7zDCbwRnUUIqvDenXZTLVyV/R+ANavwQjgALHlt0
tu3f3UugIaaMwCUB4B5MoIDe8XctWyicHIS8Cr7TgGUyAMc9C50tdML3mfaRlvYZ
jjT7BmwPuq/e2yo4SaXzN/pls1rb4RowUYdLL1YVmPNxQnm+xQBzTj+lS2C2kbwF
hz/RXY9uKltqy1zX6/KNYwL7yh4oY8OqEdUKxyd9DDot+mFXXChpfqjAlY0JpyDX
odJ7w6VzX7HEOlBqjtsuDgTWVfz2zov1SPuMYleEh6dYDnEgJ+4wFIiWAeRlTsBP
xrS6iZicDhjEYnQUfYO5Mc7/jk4bNite9t4JakUsffaYodjqxu7jH0IWIFDgS7+V
XUALquBV1U5bTEc+40XxceqhqNOamtK/7w/WfE5pOkrT3arTl5Umy0LRPbi+Q+54
VQ+NAgPPwvHOYXdfI5ZBCQpVxMhrCXbZknulwBXE1V7+GmaEpX2LAhFHGgxjzzsb
sR/bFQx9b7SeAOjEnkQMqgdhOLZjXpC01rlIoPFG7zpC4/dIlLt5o3IO8g3wafJx
46+R42nq19GgCtlvz7HM/31KlxsRgilF9SUBs63Tkg6F/qgs4MKe6YIjOk7BjaLU
wic0+dSd/UEuYhVksnvjUNHgTO54AmmB1BZdMtVSFpwdGkrp+kg3oSS5bmMUhIBu
43Mll1B8sSppqjyDYieFl7Npy1fBQYYC4g3dPABvfvnDwS0D6EX14S+LT//QyDIb
CFFdHFqkRAUN7usPkrX6DNlC+Jk4VRfaZa8mQ0//X0A7QdkyIl9CZsBYGycUU+rl
brN/ufN+NDfKt6C0B1fLp2J0cnWmTdWhFJVan5f9Tse/HkkTH4FpbW/pNcHTVhdQ
U5Ah34pGAVsxrWgUwCcjrI1WvcI/q3JqD+3/UpeQ32b5hcTwLqlBgwv/7ufnoXQ7
khSkxsoAZSEudH0YENMiHLP2/iyilCOqt7Ch4BH8GEGVpJnWC6U+RpEIkuydeXy7
YZw1RGH5N8G25INTuLZ+wPOgPONAJz3lKfIUHwyCrs/sLe80NM3poEW6Ctn6wWE8
CoGcaI6VWbMYw0ncvDjPo68gqlq07bGpfu+GkPvpr7sPL26X0SXqp3Ds6nKPtCmJ
/7yM7JoCOxPMePK94p2ZWTfsCC4MuDPjQRR5ZV5MSlG3lOc3VZ/wsOPeJmRLz072
W0JNtIzqLgulptAP9sHy/wiCxtQC6673g3RoIQIArXA0t3jdwwmLAtQYUkRvKG6X
wRWpL+QKoi8d9kpvL+oTeQ7L9jL1As6Jbpl7aGLttN6moOB/V1yIzV4UBieUkgxI
G51YP0h46k4alxS+rgijmeNhJhcQAvI9CBQR1dB4PzFOSk/SYyyBUMH3c8p2xq0H
QXFRu3mB4FtJsaeNL7hlsFeLC7aHYs56vE0Pph+O3tSJP2YS+0c1gwBYlm7+F6ia
LIQAuVIQk8wOHc2cys3CvLgweMGas3bcR+UmLYWXjHfcOdmFBrWzFJgorqjBbeZn
sop3DB6ztvlDF143U7jZSKxBfj5IFs5x7jipQWsQgM9nPBwE8sDAvq4hDTFhwGB8
0jEn/H8rMlYK/iRYAs9AOkgJ23h5OPi3oZiiyXFtN5pjIc3bCxUR+tP4ul+g0Cgc
Yeb1wvKzx1k18f3iTffcCpQVm/5yZFwMdl89akNfcxPzt/bU7R46ejuFCWuN9emt
ktTqiuDR8lNV6AJzrKjH7BFBsQ1dsnTJUEBnijZPj2YS1UlcLeH46o0tk02KD5gm
lFqFUZszeAhpu0KulfD6iYSFHQpeyojS6NHaf26F6VpOUh8jyhiuJESvQttdPx0+
1CAyVLAPGEyZGc1jTtefyFQz0X3+0UPFtRHUuex2+IrDuYxzzgh+EIr/Iqm1cMjV
At5ekRoyYWjxpJuAaJ/YtJtBjSxIPOetdHScpEDpfeqlYVvNp95/WZSN1IE+x1zf
JlnBBfIr/yaQ+MUOPMe1qto1Zx71dCzg+cHC+G6H76Y0dbUSN55Dfup6Acvo2uvE
E41+EXWYWqW7dstSVFs8mbpvC2TVA6ldV4ieOsxIbniQMMsS8tRTJpz2DU8vs/tX
FmwxMBWTF/925KQ8dyzCWsZXWeZwM+xyVtBoDmaTBNdFyrsoz7itiTAtnz0lTOTI
KZqmbI0uzGqyis3u9xBfPxKZOWOzUaaI6ZjIQpGmqqmzhr4YCTtAOgPZs6I4TdYZ
vyP+77G8QgOWLiJplQR3YAjcaRMo4/dFgAKjM75I9K7UNoAYeCgNIIsemXaiUBMm
3pURqz1COcQUVE7F3IHsISajfzLMNP0gdY3tbwTvn27NWAiE5y/MggbKFA2ar2m5
bkCbS9UUJML1T8HmBs62pCMG6Apqiybp0r3LDmUTof1/kbzQrRZUzoBq0JZRKVFa
NtloFTLHWOxr8wOt96lLYvVLgbJyS8LS9duyV4vXYiT0Tm9W9Ki6Swv60k4Ezo5Z
ueP1HZn09tX1FdCmFVDeFgik6djOYVng3kWFUZdtJqRGXnvp9gLPRpdVpSb3t1lo
NiD2YV3APYpaGgdG3/ATR3zrpIiXMiLa3P0wt0K0KujR9tfr8AMVOcMGWr1kZS5P
gpL6uFEsNK6uejz2y4ABSH6eAztE7HsYMYj/RymY1vg0WZ8BHGeZvq/UJRv+Xerk
7IpYlm0Ai3PWjOEH+0QhvVoJJK5zHAx3FTQznPRJrnkE9WyqcvR7T/2tA+o2CWlk
WTOT4zZ+Hddo/9sP4tIqOb10h8u1ZnuqwAA6HCf/nSF49G9Tx5SaJCaoBUCSNJtA
51NBDIvrMptr0sHP0VEKB3pWLwz1IEAOHh0D2bz6xnan3qjCPJaP1SXvx5k7weQJ
3lGWDWD4EYqXItBcN547z+N6DDA+tbfRnQz3LuoeQmMPj0QTxX+tWj+kIpoaoqOz
vafakmxJ5KTqSLErOfNtMBrQnBRkTS4z0ZpaF3yK1ZPXyol3TTyUBuzrzPD+RNDi
47nR3mJH8vTURHH8midvLNZR4ASQraGUE65zIkpLeGEndxyd/xWEkssnNw85/FOQ
ZdCgIvQYwmSYnHr0jyXZt76Dyb7iwdtXF3u1TgtmL9wPqyP27DFbqgadWr0mbfLx
x2lXW0YqK2hgVA6jfmpWW/s7l5Lc+ec3zGk7oj5GtodjCNoS5pSPF+ww+D3FojC1
chh37Q+60iAxdOtEQXyVcGDlmB8fw2wl0/UX8vx/C2ZPyaOdpfSjBfd7UJwEVcHk
ZXQ9EkNKPnTt7CVKdAKVQSuDg9XvvoYOVZ5iuhgBAE4VUCHe+IFDfqr/mIfYbr+a
WdUyN3NRcthY985bdRXlxFQPc5PvRfGqV1UiGwAYmJWWx0FfBx8JS0jpkH6w4LMU
iiZBSjmnYN6abIBZtUCokPT1cIadjkSK6p88T/UNh6loAqx42d/EuFUdy8JNC0bT
SWuC7ksiQhKNRtjb7PlyNGQydWICbJSmsWRvSOifDNHoLNkp6A2WLRo9XXHceolR
9Itpqjct+X68XJmuVjMxm1cxuAiIAP7HMmkLrILcJAumZpFPiGVQaCktwM2+Kb5n
ioCYfFJGESlFnPcoT+J5in4tXcprLbg7YQLNSpk8Ug9lGJJKPbtjjBluvYv/5pYM
5GLDsm+4sA0AihpsgeV5vNraVVSGv3avhLuFTt5fbH7eHEo+DM5AudDyRUTPKNd8
oPG0MoilY5jadGT10180dKoLbGwTmWCMgXdUC0sbnZ7Q3YrV/U75iKiIfkH0CrIu
oeinVk0X/CrBT5yJzhaZ3NKNDOAQWwicI+idqhEKf2irtBjihMEjXurW4gZMumZP
406rPFhCv9SPm5jpJwULmqsBQZoiqjrV4XYuoPya1eEmc0S7KgsPvvocg8OGOU8r
p8Fwgf/4gNMuSd5ZQXzWTRebWv8pMAGxNnkoUYGiYVN6rAmqmV7xLdUrAqg5FIng
j1+gVF9P3+0e4J5+RuPw7XaWsnVRXyDTDlbAjfHsWoRjaFkOhuehf1Jb+88zkAFY
ntaqCg8p0E2gZ010na8YsMceKEqoML7wmJ+j29ZIDF5oyPBBo7dbn3Fs0K9s/icp
vlzlwCBEzg0A3jJeGlcvqF/vv35goZFArSL4dJt5bmrfT6CAMQYXWi+wmhBdvKvs
c2qySyID1bo1Cy/WpUOc39Zs5S0+WDfhjro6XK/1eVNtjeArRosbiBMG9F8fNMdu
kWS012TLS8+bcHhDvAJPBquEP55u4JS7ycoHmN8r6tiQbszQK7z21B7bWt8ItCQ4
UN9biPLyXWXlPL6GizjzpxGp/kE4arIlC3esScgPc8HqB5ngy2tjmlQYGejNgStW
PWbe2SXlWDthUUyjlskfid7NUB7hJ726a/8mS1fvFhHPCu9y0tqZwUPNvKQMwbMs
bQFQ/CcAw2+ZdG88bdUkCMBvBj/1po+MEL0hbi/KWdimFQ+E/iBrSbpejQoMQPtR
xyIUXaAhGxnlawAw5husv01hyJ7sU/TQgkGYMO8QelcksB3COOnEEe89zZ57ZDgI
vaSmnSoE2UUiD/EAg3TRXQXoWvKetn4eBwOpngLRLZLwfMmPzBS1Z2Wy9oIrG6lV
3V3KHRui114eWpco0kWZCc0Zh/pn0HM9UODkX1hFv36IPD9y79f1PzPInciZ25qr
syJ5h9W0iEOTSA7Dccv6hV6+y83tpNkqNboWkClF7o22BltgKpTjnfLLkaZq16B9
JnXc/B/uzhpIzaCxWh0nafNhVSWXPNSGYYT2MT9LW8lc0ciW6ooqC1oqYyXPd75V
Q6u116CZZl74O/XxeA/44QnA83nUauqnStVz52GC9qLiyIk4m63zfwgei5uPDF/T
9tIFI1Y1LaIi2avzZVNgAqTsnYNrF5qRcr/qe3EvK1udASQAN37mmwNC4rm5uyp4
QoPFgEM56lMBKgu1cLc6MdMsnRKWWNhBUC+LP/XPua11zvCPZuWeKJu9aq6xKuhv
T8AABeA25jhDOgUXxqEJxqVLHjjOsW76tI2FYqAr4vhfuuAHPTY+0GtyTfiaSgWO
ODZ+2wGYpWakS7wg1/8m+5lORys+AmqNmmOvb/qbi4lt4QOfDu9Cq0wWH1osNblW
jMvKYRjhZm5lMzSCmkde6lfAfBefsunAb6a2RbIouJ5GzIrl18hIwPXY6yTB47Ke
m/AnXJSr//Q2WQEWQ8PlRKz8gYq3dihyjYk+hylQ8ot98gOABMcPomWNxig8RUV8
XJdEOMYEmS5kq1c9L7tCta7zVZ2xGzS41XKrTLWHhhaVgZr2ZuBbu6HrLBBaTcJI
4UbE6ccj8Zy9k+K4ulU7ap2TQUNKXJLmftaTesi4C0tAAy7Tlh/W4hiKjqpRP3eY
CZLzvdXg8T/+g+ci72rXA7tgHh8oN1bLTKkcIOuHqhDIcG5QkIawFT5nJ/CEnARF
l5UO8Cpox407LAgP5SAdEkKR4x1fSQz4bv2AhuUfOF1lmGw+/hg2P2rZtuuNHVOP
A7kWXBxWXPUryn1i/OK3Vrma3gLQ1w8+FpUxIRk9+G3Zgqmk/qE1yK7FAw6UFvcx
QARD6G7y5PtfcgtZymAlP/f+j2xToHha+xRLOWBun1cVNpzKME6/26I+UneB/4oa
5nBRSuuAKDekq9HD+iCtOdo6tJfdcJTs6jidDI40B+ikfE3h/hGdQ2GiCA/37J32
YAtykMkFpzI8rF1RZFdbNwseAC4IgwWjIKrhSzIdTCeDXlkSAbKPaZpwphn6njpK
lJ7enUwj0TC0DBuJ0FCzFCDhsVYg+TmaGWAeyazM5gL8lz+mSXd+0l2N1kh2nQhl
bq0bk+9M1nPqFLR3wUBNoWnR0o78KDsFHf9+gE2fOM7g+IoF+rdZUiFeZkbqc4Iq
7wVp2TQfxtqdHXDcswXMYs9ejEgPIj8wBDLp4xuDD5lxL83VR/ZI/bxuCXkeD12B
TWuYlfrqtgyZsvcg5ZLTAxAor3epo0DNPEv0zrQFkVrGmCeUAjbBJOUsPnKfOvqk
11ZlJDIKo3ruqbrbFD6+Aff5HUbwPlFMOmlOpfUgHYwMbGVvHbeLCol+bycPCTha
xx/r0APtT9XTBppwBZtraRKNVuRp20+keFxCLvZzpxPeMOQ7WuwsZpjcKGkXM7ES
Ir9XLzQsZLcDRMV4jjB5RA2jJBoE9ODjibBkl1qoSdXnYH+/rJzOzAl29NMV0B6U
DgcJCpoUZH+y5/2bR9crwdnpMVXxuIfM8Zg14CFFaLriSbTBDPBqDzGtta1lJqgg
0NEgP7wl18/8ztdJtUcQHHY+T9SibOpe1/P83X6ucxIG0eRAo3FQ0/b1PYIg4JdQ
r+rTPaJDSadjDeKG/4BBMvklGI6ptdCnlC9SGZWX0sgOqkaFKen/KUNIxt9OVwub
4ueNFZR4plcJjqoNV15EiWmeQhOH3EMMJbKhslvXABv2tw1mMYI2wiiW6aIjSVib
ZFyDeXNq0s69k1BvTApB+RC2lWHgpPvnll/pAN5H1VDfylY83ALTb2hB1tmUZyHL
Sz7LjFoQiiiSv1sUMSJSOt8bu4fW66iXSYG3qeOGLhz1Zv+30u3kRqQTxZD2e6Dn
O8EbU919/HvRsoHCEeswsBEdqhBTFOzU6OOr7SzRJ/YTXG2uZj0tZ/xpvrBtBBc+
CnqCT7hv5J4tcO5b3QXMUbCpVW4YD0HGcdSRN9o6ENjJAcOITwxTzj5syb2R3+xD
JZASRLxq58hfbRs4BtA0MWerYXQ7xA9lg9Y2nXZKKng65G3QxUjRJL2itqmAqQF9
G0zpneYZUBAgWMcFuMDSc33cXMDpsWfDBzINIk9T+pPQZuGaq22iBYpZL3sopiO+
aTj5RLHgbgGGpLfnNQUi9PbpSkttXnmJOwL4LdqEKmHdNCBK2jEIwVg1zkKcLnX0
clQDh+oju+JkKVcDF4aIScWAOByC9/kIF9yMtied8oebXPB3PkoR/WF3wMgIR4xF
gTh+y854XvA93kEQ6Ur5wBNjgnypLTq50T91KoaUX7cfaBEFO2ndgRXDb9vy9yQS
YD52DX610Gjy6Mm6CUEFNb1BG6R94imlY0iD8EPgG+qdroKhqyJA2VpnLVqIZptd
qqoQ9Gc2gRODVOBed99xbqTWB61c4+puaqpr4i5y3DZFs1535jc8l9HlwD18/TXk
2iYZ3nXcikDtLBIX+smkNKmkJI0Wfn2DmkMKUvN1QrM16oX1cm7DUL71VSTmjLzM
Vr8AAIfHHBGIE7xAyYi5k/dP+4TWRLxpeQ6TKeIr3AuCvLiVHVZL+crmQMIGsIVW
SW3rNEVcxCX/oVHyZSUd/Szl2AOWyt50w3/0gy5zSjTziP43gajha6pfeipabU1+
osPV7oumwO9Ku8oZef4uM5sQiVoe0Yle+Jg7SlBlX7EWhmHYjgmqLUXA0/vOoQxo
rTeVqWEYkFeGA3vaS+wH62hKxxJzzNRrlARAjeFQG5dQhJHIa0ITM5mr7BnfwsCZ
exG4BcU49tN+4qTL1uyBLX9qn+kdKvMNNKYWOrhaxUCLaB16Ue+ycYskfCo4DG22
NwTpNf/sA5XIeTJ9byWDjzeQkCleC17rjj7EI/qx50nOaCO5Dd60Cb33nNXamw34
v25SMZRmndc9OqPnmmVQZ8QpuwrNjzq0T2fK+kPLaVjBn4ELKBiAriLzaibLXBv5
fuIq/yajA2AF3I9jsXoIf1qcK2A85hq5RbdbwksnxEm+gi5tt+kjkZETqr3MpghT
gRBbR/KtrP8+i3vXxfXU3Ui1+1AZmBuXhazHjFJZG7rmv/RZkEjfXKS85LwskrPI
t8elyUcAtGpY6MqUg71vV0YwwZM/O9JSv23nyPK7ft+ZoZqWnipfA98KaQi7UQ95
AVPB8DaG5NQwEtl0Zp6SqlO780P3/JPrcdBtJBbkDSK6k7UYamgLOUEgv3SfhNgz
AaXzqMOYg7Xo9ZvSyxPWU5RjqUJceDfqAf87z0U93yFdLmXHzbJZ4Uc26ZK/2ZbX
SJEsqVxhVB7MuphHZc3+giK0ybzxcagjdeQio6vFqhAEmfnsU+lkrrIoSP3mCfK0
sOJb3XlrrDew8L+mjksub9Yqwvp9NttDa14B8Wk4601pucGrfgjFqnY33F1e98Iu
mf3R3njLFTVZoWG/V9V/qegVaCFm8CJXTyx+/bHMtqsMBT3YV0QkVIjIy2odClRy
0xAxXlvmo5rPuYJm+lOt3V272w+XuTFl4JGMo1JPq6TibJgsjXeRuIw2U58BkTU6
KB4ArOH4k2m7BjqrdTj0sWKXAjCSja2hWzykToOkUtO2Fpgv7rzvMAEyyXs02TXo
w1JT8127MkGKs5PCY93P11mFTOjhAv1hZtW1/gS8vQ2lJZPi6pLy5PN/1RXYM/d+
SPqWGdK6ftXvUtNOP1cULjUbEgZi4XWpu1Tp1EpNuZE1892y6wVkxRbxSUP72zKG
6qrWDlHqSnlXmJ2gkVKU+gs6YGwXmAEM9Majcw393uk3P7Y2fqecNrS3tV+f1rTZ
ONoVQS9ZWHkdXXj3ylKqCYCpOzUoDq72nIZw/CrSPitgfeqH6xc/oDUROr5IzFCt
SB/f/RxB0WK8aexg0MZTravfA04KXhacCfHGNSz4jOPBPo8NwWWp2jXhtsPfv0Mx
1sviw0sizrkd7a0A3CQQs5M2qxDm/ABtreSpZHDNoYwFcDtHD8zgLdeGYnPyN4wz
96he3u//Zi7OjroAS4I+vDI4fZL62yPIeI986W3OfknMKs3+0C1PnF1DRUGEqVM0
vOTTP3qoC2um1BTClUQISKjG/xHzD20q23VJshfUAefbcxU3BQ7EinnfIUNujx7o
62wzleXq0kptK6AWG2cyJwBcWjqlzzmeQkW32ms3bGy/BoXUM4lzqicxigXhx4Qs
0Dt0PzFWBdKKSUWIPtlMBTTQ0LVdBDnWxLKuIwudOqaQs7vNWlBUEBGl7hmqS3Pf
Q3vVdWezRmyNbTXDob/wwJve0RTvlli5l4L1SfrFWKtWY0jyfvH6u2SGr840bttQ
l3Q666YT+5K8flQVcUhNa+75mj+YFv6ayP1A5/Ovz3MIxJlbD9Tm8TKL1G/072Wl
MqwfNcFbd63Kn7eNmwhHT00A4PUACpgwCj898QNGrthCDOVu9nQRrhfvM/BV/CDo
pHKMFsuAbYc7kmRWqr3ppuHsAWRVz9C+MQW425bAOKC+n4sHLqUqvkrWUt27W3Qc
mfPOzaEfdBshBIsULfvmHdcb3Sxglykw5kwDKtkY5hHvkdnytxFszNTmXshxWwcf
1a/uFXUnEBatNkpQTxCSGkxDHiMY/sJbHmyl+tC/3wzydHKsRQYbiYzlkNL1c1Yj
MyTxq8KMjBRO67mFaYxVV0Uf4LtucNBV6VoMhBVFIKmYFYuuVvrc9fCiWpD2mkBb
SnG6C/IoEVbpojcX2qZZUPjGzvO51e76GueraXkLGBO8tU8XuTufGfGAfFVXMgdY
JTAgcrvpKX76Ap+D0zzk87bPw6JZegWCJauYVBkKPRRhbPbWiGW99XJNMveutRQP
DAN6Wr0+yBbO+Y7bsrd9WlUoyojFl9DI/UIZXyMxBLBHCAJV7IxAg1gGpx4Wu6R6
5nL7vpQc0qyAE4e688wtrpA9HzzOaRl0aACXRh8v3CHRaOwRUqJjq22I+MEkyVUA
QM04LfMCDyaMc9sahTlboKrrvhfXB52+LPq3JfOfnUNAWVicajlxgGZVrOBywJhB
/lDinQB0rB0VPM9Nru8ikJcWxClEc9OoZJtfll8DaxSgedHDwjBkZSXdx/Ujq8hK
tLe4sxjizLMdynuU8xKlf/iqn2tDcCQyS46kLBzFsebE70cAoUS57kLcFkZTpqQO
pngKXaulCKPTipH1a6374Xx6f9yyZ77I5W/zFse0D8NPfVmKo2C40ljfMp45pUc3
jNYFeXkjoN3oFTVO2HeDm8PAhn8sGCTM+XJsayyZoemps4qriFyIfK5LOOsCQv5K
GnYZ0g7fv7ikTH7hNHu5cWK9GAw/R95ZHmFsvsaCncftLiop0VUFXZC/wtkxvhqa
pBdQ+1nYtjQpPJ3hFvbBSfy3u3e4Kc4vDGx9a01wFC0wI4+mHc4qf4c0xTrheYGQ
n11liRG0sbaFVBjf1l+x0JINkZzT+MjDI9+SGvNats8cbJ1rXwMXSpZkQUH4G2Ct
qX6g/RXbybWuwfZv+UkRK0MveELumVZu/pydiIK83QDyeK0nDE0ialOjWllSubFW
hrSjRvKpltFqgvcmkbf1nLOhz6GiOFSo7JTqIQVq1aKufgjm6bJEQ6Hz5UGW0nBx
dkWJQrpTsUuNGOpNXx8FElPalUmejRT/1UeLGOKULAvF4I6kd58+xVh+gqaK8AXZ
RhxQHU+DPJPTveHU4hUfzyWexvULhIjsblPaZ1slbvUQL8ZPre3PXkUqO2KxYjb6
vbzLO56mtdjRtEro+SYroBQG5cbHo/E/9bytW7RDvQZTFyK/chHvSmEJtz4tdSst
+vpjNTa3xbbGKcbaw9Bg6S2hH6hRsFy/3bqvsR2z1lMyHztJOf0XTa8cOtLJzm2u
SQ77DHp2bPMOBaUcHwNiT9LX3TTugYuVTEICSePwimN6EAthLJ2MAIb19BAB+hbD
P/10PIAYCdPJbCXMjF2fl3EeVn3tOSkqGbOcF586CUveGQo+qO7ogFkTFDMYtxYW
2nlxZEe1CiDItQYeHi0pw6lGyG20NRwUf8ggiQbajsJRSc3pyZyhHcwJEA1yuo9W
ZTE9M/DCtLbS/3hoGpQkw+s791S/BuXDUrjxTHhWqei+yq492JURgm4RF/1A+2i9
+bNd1NAr0cACMvGwxUeA+TecXVsbqlkQbTLVWlPS4Lk7YeXaFsejlMIGKPVlS007
JjSfwKDBT6+9JvP6pVvpCGxCyAhd5EaGKNwmzwD7498T1ZRD5qW/LuHtMG8AGz3F
pwPGYmuKVTbjqSJHtz450JQEVtaG7ivFKdXDPdhFqb78My3YCuPQxtZVWSSxlJ3U
eYIyr+Uo7UUpjCbaCxPf9+kf8p4d+9Gu3SOrqCRweuyNHx3/MQTOFka1CO9Iz5r5
lce6j+snQ7WiDyDAT97P67dghvupqmEfFX/2QYAOEcPaSYbWgbw4qqfcP0ov1MEK
FwllNcLk9lue+khXzHaWI995Q+x8LWB3N15PLjIhrH7o42oWG6/cJhTgX14B47Sg
gf182JprwGtrVMGzl1TDUL4m101TX8kNDVUaN2h5pSSLat9CFHRlW4v4et7NMcq0
wQU+7cR+pDvTk+8jb7JhnKUV2uCoTipPvi9OQsqwjcBp4GHRpKvpP6osLdU4LCj6
QjCHcyaGkSp9zc2AhTLsKaNFMRD2aclhfRHpZV4jeevhOQAj6XaS5nrW8HwvVfN3
sq6nJMLYqLoWxR8YAxONCezsLT+3qgZmQIFxVivVvPuAqDr7BjlbA84c1T+d/Ggt
XpwrrDmZ3bsFZX4mHTNKUWcXBAsWQfGrCXd+crQagHfitCJLuLyn1A4+v2G6mF+Y
Hvis6h1EnJoqnxFWOtNP6TUccoPQmvF58uREmU4VaI0nr4Cl1UE4JwNa7zyJWa8q
75LLEUu4wOxi360i/+wjVea2S8FjOTSLBvth4qmTG8V5VYVQ2Cxs26GdQH4pDqAe
RQFx2vaeYn+IcDB1e2KLoIk4mpOCYfUj43dS5azied3rnOHsn18/i1pJZBXBov9L
3oVkw7s01hJTcgXmIlx5PnBZ6g5PCy2swmxuzVu7EetRpAJtYFTbpdTo/RkCIU68
mPsHONdp7JtsfaaNCaIHKQSOkKTV402jlxa+XMifkoQsrbyAP+xUMKc2AE+v/8dG
m8MEuAlCV0IFSFb4r42XrnfofdjGrSM8Krmsg6uRHTtHJHuQexVbRgCLt+CWBY5N
k3UmbdfCDTExlD5wJmxtMfISCuBZhrxrEUPRnusk74a1fQpu6xf7SALfeMVUyrRu
uCuW6I9Njh/9Ljr3xUB54HZVslRojMtIS7KnfKWupWowwBhrvQzzAGBZOLK+dS9O
lxUKKa21pQ7wWb0YZf+jO4ZhK7Hu4LkQeGw+biYF4SafaPfHeFxMvDUfrEOCiUso
2M7blwAZ2XJCSfMwI/Ujp779sbyZepJEFrfIqh9ycKVytGV0m3UK86sYHeql4M5w
WnJBMU/IXam+e9dC6LSmu7FIIWNnkdZwyBDA4yE0+PFG7/iGqHb9OY+ZiItStxm0
0lf998X+q8j5P8Ovq4exL3QG8s6mwfuhlwgzYbuDSMgmH9dsu7qiCmQoPVan7GIK
r9YFY3Orc6UMXg6Jt9HrQHbuul8nFbEJRfB5Ysz5Wn92gDI6u7vtLqSLshourLVJ
y0YAKHsaIsSkec30ynQF//D3VlLmEbh46p9NpGSmCVinNvHdLnjwKg2z8VX8bmId
s1Fkf5eU9SIEO6RMKg+D0o4Jk7nPc2sLk2XX+tCxHZycxFBn4D1OvsSN1/vJvzI1
rXIbQX6ow3Uovmf05CgTmtWQ6hfKYMWbKiPXO3RYJQdyvB9kyB0yYt6PLqm7TTEf
uX6o5MFMD4gPFXR89XCznYOqRl4gziBm79I+ZctAkl+SUxXKSRCxxlfdNvmeD4fP
dlzGELHLqKK7mTPS933Xzavg2kD5kGrlzOG8OkQbg+0g42y61dWtTqsqGaHF6Hx5
TRIcFDp2mde4AAApzOff4YmNl0wQC8N/Dnwo4Nmz+59NzUs9R6dFQKJRkbAojqBY
QJ4tMaS4fRnrARBbCyJ0dy0OjKxjmY82feK+SgiFCgr0W8M2hvwqiyLWR9XrKs+i
uQf1ThkYnbzkqRtLlvnUFG/o1LfiAuxCzplPwRpAlMEI2dn6sfTKwgoyH1OSW9d0
0XTtlahz/EjBuKWedPWj4MOI++bOxEDa6ExlZ7RguGyGz5tpYVo/+wRsJSsDbUQT
Mo1ii1+6vKJXzERIjulu0dNDDbhJnnxEfWNzLB/z8iSo0gU5Hv6WZTodTPLsmNL4
x4vKC0LVHOb5+Z+Gtc6NFruLAcGhWNjr1hO+xfq9SVaSrgkIaviD06Qbv+DDWDvZ
NQ6+qsitLgVaAZiCRKCEbgnvbDEQDkIJmtNkURM7qvRJvP0O71k9M/qrvw9Ewd1b
TOUxPUprYvVztOOB/xVOyyapS2fPGG/IW71ckUbQwjvD2/vzoR1/xx4sQ4ujMGCd
n8zLlIOeTtZz1znnvO4Je/rknkPn8Rjrwd3W0Lkf76H3ka2ffdKtlUR1hZ0a/NvR
XjfYGDRFbj44dv5IdC7rCm+aDMeESeVqHwFTcVm3Pd83Af9g1GgGsWu6ilHQRWUc
Ewjk8o+BAD0A2t8v0gMFTxEf37r/zKMOpszXbHMkPe0Hx5Y4oHHujQ7OpQ3N1ugx
Dnl0FaB9zgWJlQifHZf0GUuUsQFxPjMlieKQfrXHNVrRwkUDo4+8ncQ2Ws+AlyDE
VBddP01MfrJb2FPZbFO1SHH2KG07lxlj3bq8UrR7PA66oISU5ZQG/MGc+um6/Nfm
McfIMa7+/8DkNBJL7ImR0w1MqGRICL+yYmbbqt6G2JTrdWmfOd3olEBYW6UrH1ir
LIFyeAkXPQ8HEH0fUqSOtpxkQ7mfldmU9xu2hhfN6EVAM2e1aXnpJbckI+EiVevE
gcTqG/jpwzwLEjlXh91kQE1zrsqfDzLyAvGcJd761aNWwJ1RrTBYHNL5lAPrHCi4
/4nDmdgSVTMJJH7PZWokM1rQwj+vXJ2r9utf2hZOUXejnaVBUWGsBssMOfHDJ1gw
vtOyio89kIEWR2+Y7NYXKlM43EmZ1dDAgSD5TNDlJIGeHiD/XafJduI/JKg0UV5Q
IckDtTRDYrZyEH+3MDAC/FqDXH5Vy9pjFTryNWdoxj5kCnsdsFHoXC6YwK+6yshV
6NGtIyruMaNmV2pYHSEMSHxOp11edGaqTz8RUSyTEwxxuQL1LZtu9uUhN1UCTKi2
4GofuJNOIkyuv3FGzhs5lAdVrnoHvDytmSKGlFouJIC38x1N/yTxfwOijrsk3JZs
+XlpQTrh/pB6ghm3AIdqNIueq65v3kMHslkJABXdTM476vdPuARlSy/foZeJWUFz
rZ0vNnaOXWQCMgLyKWAYvKvcaMXaucaeOu6bwSI9cdNWZ7L3+Jk4W2IWn2vUHZgh
rDOY4Kf021kaxPplR5jYZjw4InZ/lybKrcy1IcJzDZcs+Q8RijhJIfzla3bB5ifO
lMfF7ft4X7Er7T5Uv0v9G/dpcg8JeX7HhRwDtmsOj7wyNQhtzQAUVvOZQnUUVXlz
5WQZCbeZLSVPXnt6zmMdt2MXS46fKzhh6ZqBnNam8rg3NKFqB+xUdic0x6nj0yeT
fTLU/gzOo/YaKI09fW8HPYaz9XnIicb4tAUbzmoank9Mmgjfi+a7114SfD3Hdjdw
7vymD900JL+jZtZxMexkDy1llFdGTvUttisCrjVTnYJ8kDmbVF75aDTu/zrIz+1g
S265NlLKeV5PGmRcklnyq4CjMQt4ylFofsGbe4pMYLq9sZ82YGcyma1VUD6y4OY8
WEYQ97SXicYcMY7cG7mSnwYbLyCnx7m8a7X5+6o+oSCmiNkI+o/c4/7K9s5ZXUv0
F/AK27amA8dEFCEPzV0Y4JZ6neTEQI7pVBsLmg7ftdM9OmTPngsFDuzLGzZFo1kL
/YRIw/JtaZA8/OQnfSI18KrJuBHYEYFwcRqYPhoblb+soAehSJVINo0o85EseWzD
3DOI3dZwGEgRaAsJAW2GujYnWWr+Sp7/Lh2kihqURh1cc2frXJ8fAyQ8ajK/sCYm
5fCUlhYSttPEH0Cb/4oRdMQHDU/krgBJRrG6tVwL3O/LsfgbyJ6rGf3aSu++laMR
/WECe1GZfPci8clb+ZrHdMQQruhb9XFCqN+9uU5kMN99TtR7d2SUGlTK/xkqm8Lx
T4YB9pWwFxjJs0NFPBTiQlRUG5sZvYTDSGukZsupV2fMmsiEsDRGmxIJzBh6GhKP
azL6n8Ypz9rCiin91YBmkpzAbTU9L2FpOk8g/pQ0vpNpIehhTgWV8AZ/baBgisOg
Ye6Gw0Ue8ugf/76cZTn9XXMqL1VurJ6o8UcyrtuMgGpzlHGCe0ygrDLyUih528rK
CX5J5eUavyg5hlfTnSDfJRZ9fnnLyBNF9MPlysjuM5qFOBZ9C4Liobi29j9StYWo
sjI/+zqd2oge+4psf/5PJ3EDLDiweiIRw490QyewMRC1xYybw0Q5ovVmMoaWC75I
vwgmJlNkU0HL28r4xAzXy8PPHJ4oz/JbBvoByW71TFMg6CDmv4Bme721OTdiojnt
igaaAKHMtgL8dupmi2aFMMZ3vTOCQ1Q9tY11GzDw3ATKOqkAYL30T3T54qv7V97J
+OwLzZdMJLHfDPICH/KA4snDsxzhhjyGuyykRIoAPq/5sbovKeQi0ta2bMBTx5az
RCigMES4iDoMmQvecGvsxR90bHdHA0M/tPaiJpDy8AxTziAsUo7fBIskJ6Y57qXI
Sul4JflyXWOTgThjc+gQmXOlJCCYLCZSz3Fk/hoFVPPKRJhfYcPl3KqJt9qf0hh6
ziIjt8AfeVPM4DkwPMVibAirMHv0RgMytD5l3lJ9lCMPOcXeniZlpB9N8X/ty0aJ
NN0u8h3ZPr/EWh6YqDOSwP0ITcgpZ9y5jPXchgoOn9PLpLyVv6Fsbd8JoijXvy+j
T0ku7XVJKNiP7ghtZW4cBwcEVTimYxe1izrDCY/G8V/ILESLEBCC5Xeq23XzTMU4
hPTqY8iyFG9r1Hdr6Jv9UFYAIVdmnGXEny7piVdIMmshZI9XUThmWCcBLv9paxAo
K8pxBp/ExtRQ0CzD9BycgJ0rQbxh6sZmYmtdpwap6+QmgfQSlDzfa7mL0OhOorUG
/VWucu/ep+sKt5BsW0SHTAF1anev0DOi6zG2eywq8okbUxP06Nb9ziYCySsTIhAE
J1sX7Ae6aGlA5YW9SiMLXbOXdRzXu8bjUhlHQ5jtkVvluup1SVCGAukFi+EkiQTZ
but/+eIgDp9IQrzfFtJO/Vvei9XoNNXI3MpNRVYaMpyZY6MKNBKRsNph9KbZnrg0
6YFLwgXiC7qEKFWATz9MAXgMYbIHLs8S2S8y6AUqw3+vlgBcHKyD4eS2J4fFHNaD
AZwtEAruNMv/UAHdH2gSC5kk/QiSI+9kCFm1cEH1c6DZxuubrGiKbFvcfl5QSe/F
NHq4nZNjde725eIcsCu8x+9OSaMKrnOAeTqI2mThYUU6qQMV71fjESLsIO7isfjh
40otWsw1xZMYA6iOiHrmCPFeo7IO85u7jsM7K+l0vrBza3s4N/PGKYj9y/aqr3Vx
1albO+HLxfAFFZZfAID/zpr/44B6E2VXoKXi+SS3t2MxiKj6ao/wXbpEdlB9I5av
tkzR3RUZ1kzUxtSTkwMTVj3R87USV9ckx2ymyh5wwO7PODTyJyXevS1rkmAqG+Sc
H7W4VAtL6vrJVcNfQ8qlzxNUZ4nIVHYjmdRh7jOd+017nrDR+XXgIsX2ZF5UwnxM
msRMqYOGXOwf+WY+dNsVCk59v+xg5CYnIff/gRUqntWXx2R7pJPLachmvfLnGn3S
Vb72PpFPbnguWVoYT5l5vBbTihQLaViQ1k1UweYrTIFn3wqetmi1wPRC/tlI0J1/
Sg1eSUpsYO40UKajOTlcis7qjslDjjxDApW3x/6B/qe9KQeC02Sd12w2yNoOMIq4
ayRbvvoJd8l5mV/2xD4ipGdyAxekCRLTvrbwRdCviQrxC9SBjOgAEpL34ToFDtWQ
KqrYm3p4JHogSS2JIfFVI362DI1ASk4rh3Y6YcPPmHfWfKE0bH7RZxGI42+qywb7
kdg7nQhneASGDy7Munx4D/dLKl43VsmW6CI5hc4gJRaqKrju2PY9T+O5YcMKtvBY
M34LxNvaz2i4e94sNogzsUVKqegvsdPYkhB6duuz5OgzuuzJFaTxvLlTmLJtV5/f
ZlUVu2pli0wsJrHgfzhMZcz5iBRc2gRnTOeyVOvC0dxh6OEwtIuXeoDTSqpM7+BU
pSKuVGrnqTZAoQpn1zr60vlmGPtZ2KNj63Ker3m/mB5Vf3aOd6iIG86NCL8bfgJJ
AqpxL8nKdyS5X/4n7Mu0Ryg2MITMi9JNkQSRpDUWEL4OQtrWMJmkb+mpyo9Qw7L9
gDk0M2D13HmThvCoMJ7HEs2Gycxf18+pdaZUbKapkw0GP/4qH7FN/yw2fqSMebvU
9RKM0MAmRfjJjU4QeWd3+8gP0yioswB38fhDrwpOUs4wrrrvX62kipwDgR/k4NrM
w7dBAA/iDNzdKXfxo5KvRYI/2eYFMAtk4gMGKrDzSex45g9ZFE7SrkNWSBoUNsMX
UygIKHp1v0IPbrPD4S41mgTMMs6vY9HaOurlbqGVmEgWLAAYpL60ZgLnZ//MHoJM
QJT41YSklEgXFnX/UugI/9YcserohjA4KlkDv3z3bBq2Hfp7PgvzwLitOj3XpLBF
XOaIiOF6VtdlSxDgiwJSOke+JQPjoUJZSIyNpDzKnnLiQTGA5HOBxWb7KVSK6tWa
/oDUhem1KIdcQaTnhGxvGJzbd+lUuch30B71ayhdDyqTfEQyBfWfgm/xe5Elivsl
Tjne5WqVFauZVTj9pR7UB0TFMxex3RLgRfzCJ5smaF60UxOKIyNcUPPR606C9aeE
t/uQ3G1iO2/uiZfbmGGml0WpR3ETuq5OLBYKs3xM1JPkLZS7F4smUMJLrcWIIfBZ
OZkfM5AMVITSX8UPtUqoI7+Vz+Rdiijw/JedP8r2lSgulNjqRJSVDD+JFM14zdUF
SlAY+E67Vn1xAbu1LeDzrXNWqlhmwoKfeBdRftqVRQJHsJcChwJk+4lz2sLTgvLG
G8KuLapWIz4zqzacPcu+zHmp6zvZutKjRAbW31T/6Jg2b2KUY/TFJP+CmK1uJWhL
u+UEP3Whs6OcVUoem+y4S9kLxKhL/PXgBziJRVTQzIE8O23b4e9d/VR42s0ZJuD8
q0gMtQP/wMkYpIzBlSLFvV6s7nGds1MafyZJLXCgLdxhGtZ8qwVXjfGvgXi/jw1E
d2+1kZ/C+2iJDVBD0mD9MZFQOxLqpsHM4VNyvWdS6Jpzt/jB4IjnWlem5cT8O6Lv
gEHBJDgji6pw46JNln9UEPnF0C7CHvoFqru1+PXo0ZE91gWW8ML7h+jgh68tQgGF
03kZmLurKeUsLlPuIBQuh2QLeJ/nxlG2AtVxbcqVX13JJpXsB839pn0ZR5zP0Ctr
NAQ+TfG7vtfRTHxtYB2DOduKQq9qVFienbEMEt2WPbiw+9MuPvmqlexmyemEgzYF
LGXkyI44oV2L0OtShtZtqHR7pvuAHJmGyLQtrRetA5TZV575gZtYT7mXZCU1QF02
9Uyb6PwcXxwbAzGV4Ch4rwmjcML8/UEixPF44gbIG2ncadXoza2PbHSdJx831Kko
EQnwnrBNlUkxhg6KjrMq5j/Qh7U3om20cSoCVpnrZH3uKs4YtrTAIvak55AXzek6
Hvg1XdohY5uCXhsvA3WwDTCxDw9/C8/YuawUgQUqcoLVSFpEGos7PPYhzqDguZEP
dySNfWjuR/Mv8vOCH0St8iCv5kIUWdFFpU0KLc//yw8+gzzJhRq+7e49z9HuYKCh
vfrU660MZ2eIwh3d1Vx/XXBRBLa+/IhHnhMGjq2hGt9rW799MWtm4tVG89o95wxr
xY10Kc7GoflpRN1pxS97uWMAGj/+KmA9+7uS+/urL7Z6ditByTyKM+SLz8GxiPcT
ZTDcz4jr2BtUa6OsephyZpE+omEjTpkR5FoXr0arEQjeQnLOfnI5NlfnmVxo2kwj
9YggvnkHPRGdjgsj35oqQUnTysyIVyif5e2QXCwK+QxM1ieKeeIzwZD3ddiJIyXf
3OVQ8BIWkWV5mQdyOGPvWQdyqqhVwj91dBjBPXmijHJaL7HK4tBb+VGSu13MDb6a
PrMLUhBMMSXtBAFIPaON1dz9bCjROda/br1vffXJRzKKbvo0eN4vP2TZuoTRUUCI
RIVYfW7AvSIOYxlY82XG83TzBH9JbRXT3o37yUivkjrmk3AGmUI894wln0gEdOCj
3uoL0VUOUQ2KLRVBC87KUuUCwoH+lZeR8CVABEnoYwT7HRPCudG2jvItRu1t57KT
j3GgfxhnGuXtmYcQHlUZyX5+lXEsugYfoK6WYImAiRDGTYUm0SoWVQ1z5LrSMghU
ZhgV0DrAmd1vpZl/cd5wRT0TOieBx6mE8tWuzdVPPzv0pnYwnm5m4KrFa55i/F0d
ACnlj6mS78cBCjBGpJXHqJ/J4rQWuc4hHaS0McNCeURayA7N4PwyHI2+CeITeGOg
Ft0kWuRUfpGf1AIpDLc14pei8cZSjOjqNKXrN09Kqeg/yKT/T2hAd7L3GV7ZHcmG
QWRJi7DG8I6tz3vhmEGoLtolGwRnrL8TDCUdZNsHa0Lw1UmqbrdnRpWHk/JBAxwg
8bPmVajp45wzAU/ETD1QaODUMyhvhKcs7TGoh4TDErcMGy01Lv64tAP2dGDqcR7L
Lh/MMrQgAPY7nU0RtgF82WfMytMqMuXwfmTpZoOZWKyF84uLBsAI8EQg4zciAPcU
q4uLvwmx+i2jFNeX3t9rctM5fX1ZTkZPScKEks4VjOwf+FbDmlRJ6fyqyqZEd3ZD
nWJfULb4zV4yhvwes22P2RAMZCZr+e4CZem5O0TXE9kyacpwGW6JviyVNkRsIur7
uzK2bTkop3gUflvsn5gS1epL7LuHw/P4wqVzDCyeMSaNVc5fuh3snQriNAUp8QoZ
wBtGLWrMW1QFXCoCbl/oUHFtDKnquCrT6KFa95tfXMzYGoennU1ehf+WNPp/WCpr
uaF6yZmxnyyOSHT36o5DzNYkjPzjqLPL1NszesumRNs0Z8QmubP12t50PWABHWEW
3D62mc8CW0hw97BeAKr3pi0PyCNNU8NSdhB4cSVqa33Db76nlb1roWJZngcM960C
6WW/qPwAr+IOjuLKW6DxB8Bl72uYg2cfo1O/gJhjEcVZZq7zTp6R40iv7iuW94Bn
1VdvkTa+s4ExQ+nACi8b/q0nKLQ+rX1yyO9i1KDZLR1AI8W3wTI9gGQsyQW14a5T
8qZcbqxfTElP7Spm8/6SGf9mpS4+WD375DwlLYuON/lnZ+EcpRFQ+egGyVJL3dY6
wafck8tees/oOLnRH2tMMNaW9VjliW6JCWWVGsDe/KPQ2snA0AfWxB7HrDxWV1SW
tYEuOaxAeeAsnnnx8iQu2JVV+Cz5VzHr7P8QjuHb/rCilZUNWoSnDftpux938YbY
OlF8jBzHPF/3dKaJb3zbjg6wYuUE/Bigr4pZfmbmyb/BO395AiZqtxgJYvlffVNa
bTNb8qKsNjwGJQ0E7jLqU2P+rzM2kw8JirYGYfnvo4xlMHX+3zqGuAAWqUH3mZIc
lDft7QmuOsCk6lN10Ms4c/VFeh5xNiTQcp0dcpEaFS3BEhdRq37cy4M+uRf8N4sS
Zqo3iB6/LdZnkFPA9NyrY7pIh8at7pORFPnvArbLmkRnvhOvZZQoafG3FVPRnw2H
VDkTQeeGqImjdhcgsship3uvRRVy+CkMiZt1+rMrVAIzjTyYHF0oMHuNPDkK/IjV
KDWZTYQDQsEFciQvXrwHhluNLqY7AHAphw5ULG9F5pmZiVWVCDsVwxuiD9Bqerth
ds/00hlJmLSgPDDuv1m4/i9WYrBdZEMjJVAk9MzUY2oQajlYPRiyNxLHvHDSRO/t
El4V3IevU5QJoMZ7hvEfkE2ROjSDTVDkFRfMCYJkeHFb7owXLv+5oFkO1sIT8pja
lxNxuBCpfyRaxjpGIcn2ozalj9U7bfoL7V2siZ6wwt7mQN5Yt3xuLTGDaPq4w+JY
AyPQ+nO2WnniBKmN31AdiDJ8IxAiDYpBjDPTzB0dtTT3Ahtqn/5ZhXg21G/7v5vE
TTPYD4w6TNbwsn3HSUdm6+YFRCqjOK8PfvplWTM56k5tbBSx8UMT3D84oJ5gu7fi
SlLwW6PLbwUIRG6ihmwqr2lpPbM5Uk0HS/wd6IT/bOofEn7LzZgDno7BbovOUPbg
RitV2T/ByiTVc8B0ALYkuogdakpqoBCuyQsyfS/R2TFDhf+7qBlMKFrI2Aa2I2hw
rHMubNi1yWP9i4JZmAJ82RqhPKdpuSiCckxtawo71KEHVky99iXY4sdrI5wM9F3v
pBAky75aarMPTTUJdqi8All7rG4mwA+roc1eIup/YfuVmJVhrnP2WfoKxhiMwYJW
GEyUrw6jko64WyM67o5cFbCQknq66JaZthX/U9plJL4QOg1ee51WuF8S5SlcUNLP
CD4PHb3guV7kVRuAdZ7MEY2VZzUeVN47oHAlJ7mSvjl0e1z6e6659Tohsm9Vx76T
EmXiDbw/tuQDAK0+osWqCKt0B4crnSR3kDF1lqSp3SrX7OGMVXQAPeo+L1cgbeh2
IkzIR1hvCKL/VjYJt5js/wpX5mhJBVqmL0cLbqQXiO45Ziyyo9NlXwBV/gcQ4JOF
bBplx37yWDNjfeeaQl5WdOOswyqah3WfcwyRJ6smM1UL1MEZVAI8kgFof20q3uiG
PjruSK1BDKHip1WbCYsjGLpiDUptyOCSxYVPoVT+3gdJt3eSmxjMZgx7S6EDwWKi
9ZS23vZlB35AyMKaHDxzmWvNvO+Vq/GrMsek3DwYQeRcPXUWF4yj9zu+K5QJu1We
GoYDZlwuWh250gKMd4td8iG3f2TDYBGPy96s4VQ4Inm5HHBUmwG+fqwd5Qzok5eM
ClQvKlezWAMfYL/ZSxU6gYpYsvrqyDFAgDgd9NnpPRBBdu/ElQsKopyD94xWwZdT
v7V6lQJQtCAP5YvLfg1b7NDTQaH/D9UK1idtHd811DePW3MgeANj2C5jk3JRIDnx
2qg+mH6oPzMqDyUw5XJwaYJmyDVfVZpmzsCnY0BV5opQysKi9R5HfNNoYfeur7R4
DqNFsjEVvM9AmGf1//HZEyZ8dGlyMbnTiQkAwp7fyz1FcvnC2XbIk0oxyREH+/Zg
q5Qg/H8KV8l/llxKBdOOGZSJ4Vr0ue/B6EKpFCfPUrYky/YScc848bYpJpy+iKyn
J+OrxM51BN/MING/opSUOrybPTddtuDrElw1Bg4/M3n2CFqe0sF/a9eScBXJG0CJ
/xi8Owema+UGZnEzkueLeA7mK/U+wHavWldMeWQfcTYXvJzURQyoKmOAE4CkEJCl
/ix8L3iOeu32hHwnuuMpVPYNsoFQjAZ+B05rtphVIVGia3s/q0CLoMFe+9eEtUJV
RKR+YqpwsetupjVgMz/ouoBCIxgdnzkYibFSd3xpUnhAZExejIf2XtYUNisMF9Ll
cw1aJiMdJIEsoJYIPhuwyc+ZFOv1CtkhkJjiBlE09X5IRE3W9A4MSrALNFwW9Suh
eRPDDXk5EMtP5VR5maQSEoyGv+7FtieNy1Zi1V/VW3ig3MJTzKKq0jvDRJjbKfzh
ikGWJUG87M2WaMYK89y9JGWSj1ijLzUrBViJU4qrnMtC5LM+qbNxrfhRGnvYDBo4
oTjK0Lk74gZntts/nOpX7Cr3dmqgjkCCJeodMXAap0Z0cxXesVdL5orNoMjpXfNQ
l5+EGhvftsXwICd4wWTG468SIfj1LldrtxM714K2OcS4QVo09QLO1k0SZj87+ybB
Rtf491V9FUl904+hKgKx0ZWfaV0Y2KQ4H7iZaBN0Z4QSwZ30xScRwEx3/3YsITo4
tvUX6XA5NW+7zOjl2Z0Kgs1YX/MDNx1Q3p0TYmtt7kPYTAa5bEOfG7FSqSEdBBiM
9f77qJFyP++2UHrYlxiPJ2ksdwba4RMbYkr7AWCP57lhAu57d+SpayJjsh0LUAzm
GAsNoEC9bS1bxkgLcZc/Dn77EiqTwfvucFHFz6HwFEzX5mt0IClqcoMM9Xl61Iq5
iGLDnsO9NcpYc8EzcivV69v7vRwaXeejRGMpNlQIFFoOR2YOtTQNi9kkPABFBK/7
MecdanjNIIz5o0THTmlwbmltSHAiv5yAYo/V3GFusa4zOYcOx6cCcNf5rptQcHho
QAuPwU4kLfpekFrG0BnvAhYk5KoE2ZI/qgHh9OqC4wbOdO7/658MVRS+2Fhkxp6t
UeWAWIgFf9cuuJdQALY/NS7hQqGwG5f3PHalUqlU/KGEQYeBK3KTPq5+R519Uox9
JYx3tth+bTP5bd22U4MzCyT2AeNIqR/bAMe0QSKkAYn/DHaVWX09UarZIWC1FnfU
R3UMiG7kLebdgtf0zQLYan4p4bNWbZr43Mep3cZ7mdV9DEfRHRhi1KOzK4/cqw1r
pNzWtiGf4K2oTI9qUxwvMVKOmJFy5VfymZSa/QYU1VgIapndr30FZwhAPHQoPaNS
zx33hbqGZXETU8mvmLATJGlqAgOGzZzzpr/aCnXL3MAIXB6yeFrLhlunIU68bCq8
y+Bpuu+wgLxkeskXRa1J3uynxbc3y4UegickFeu7+2DaCw1vDapikDZYeWnoihWB
g57hDSq4DuRMBGx/4FYl9/tB1SUW5iMnZpx7ik87TGHAkN6WJNAMnGmmNEQe06i9
ZFvTeOlSdivK126IDnY7FKaLxUWGvG1zThZdYGLNZ2jiFBH0qB2FhUgG67RTeLRc
3e5/ALfnZlz2ZYccKiEq1ldr3RDCmwMyN3XWTT8AxdWtN1UqAfPoZwn1os8gqxcT
sk/sodHJsY2mwWAf4tj3uv+tbc1WqB3pJ7OWhKGwWRR4HeQhi8IN1d1E7p0DRBjv
hKlqBqEDzM2tD793UbOhAdSt4xePfwNDo/mx0LSPxCllT02lsckoJUtpOvl4GNhK
PswZp+iWBIJK0CRokKQQTWdncULAsZSYJZ0PHXJId1cFBU+2L4VFoZMGoxL8auFl
/Z49ZlWJ+57lNjTf99+bvyBRNfAMnFps4A5Bn7TP3i+OMteHK0rFjKdNlNiSYxxx
Le+0Dnp5Hmi5ulbECxjNYwRpkcv2Xkt4vP+1G4Mda+gSkfKaNC/rDeCyspbebhlU
x68UFhedKY+lupFCWFb8HC+fulZQBIvWD/JOdWP/O3a+OA7+FkxquprqRK30ldlN
ESYbLR5FrJIHF3mxmw9ofL01iur5v1K0biH7pnrP9t3DUe8cjI/OIZAsVJectdmr
+TpBo8v88dMP/4D3tDU2UZiStvEiuSyM8pqeIeE4HVpvnztCDdkRmz32xPbKvHNj
EWbDYi1E9mx3YRUi2qHpC2BQQznk+gZBCc/Qt2GXGPknpHWxFcvsiDIgg0ORKDIG
6NklVfBrMNzOJ9z/dsPn6b1zHzux6GTuoBLcMZiC+hsqhr4eUT9OMWfIrpbaYKBg
6JRL7m52BRy3BsVCeTsnBX3QS9Ya5UjzKbVS04zNQJN3B49lQjx02EZZ8YaJr4g/
w/5cpPAghQwUmzg3E9H2x60VgHhGSt6yft9oYttUnb8Tk7FUH/RimNB28OYvkKRc
GbQqXesHsg61hhxP0qm1DU05D49jJ0hQaDZKob/gBqcUj8uqy8ufpAuOv+dZ/VZ+
b+Sm7lB5bHQwzDkwee1AdHHw9rRGqxvcIufufVEc0+3qnCltpuOdvFm4Wzx1wCNG
+YlZLwUq1NFYeiM+uzMvyrCChoZVfZq/jLf/ZZiGZXZrDnoqpv56fbX17/BnHMUz
UMC0vGWIhezq23zIjuouruEfCqQdHOCBMuCriGk+8X7Nn8WSV2AKTY5yQm/3MQ5b
pre6DH6tXSaK5le36FVhxC+rXnnvkD8P9eaCDK2jtB9fVKZ1qzSJA9rX5abKpINl
6lKY0gR31+PAmbeFhYaZgNwQwPAY/CQMVWpB1usWvTxIZLEtBDczfIPKXb+WE+Ci
kpHjEMLwNB78G5Ax9fop2O4W1JRribUkwT+9qKZafZJ68bfMpc2QQnkHkKghZ64U
iXv/QabxdvK8nXjMu9ejpjcfqXf32PtgnoqimrwnhsU60KKbNZ4XiKZk2ML3pHEV
UF8BxOkZuHLf+kotJPoxM4cGfdZjN5Tak5yUb3HmKA2j73uHiUPSutd9FkdfT8Ev
ufh+6+0CoUE3KpMq8/3Wwx9xtdBJT4g449Tsne25OMgZLGl3Q618dO3LKFUylzpn
1+1iCmAK9l4uI5JaUg0/jegUZdJWSnkbip/ivAaLj7N3tYaldrfq6u9/7mBz49yl
R1l6xWbeAEDWqBIZFlsROZl/e7ylEcPoOaHMNE2M1h+VwP+6qqgpEQF1NKPAZlUe
gYkbTIDpSl3LzgyZd5CjetOZMJjRGB26mmgHK7uVCs8894XD+YSvKLRjQljIOW4Q
3fzcY5S2KX6xngYg34vgcQphJ1aoPmX9PqP5VKLIlI1XmJ7f7Le6wWqDblb4m9+t
G6IxclmZSh8+ulswZ2zaPNa8LiAznxJW1fYesi3z8Q6ozA5Qet+aOFGsD0qVsPoq
B6HseIdzqP6g3Bt2IgnMpZ6ze9jbfuL3fUqz7Dm5yIhVyakr2KExKq/HV2sZOune
sXZxnvFcDzmukCCsKIsJvAd9hWVd5f8YxUCwnUrIlG1Md4bh+h+l3h4zqIz2B6Zw
73oZhyTrMhGqFKDCGMSDY2IxPa9Ype6FfbWs43dAH8fmUr5ambmj0jBbyfPQFB+U
k9SVXFM0aDVFLMWbIiODjKaszYH+XcWvBX8RISq8SI2F4glChA5fP4MbomFHg3gY
ZpoBcsQJ67Q9cxJtsFDoCKZlIQJKOtgS4XJvSGgUp9A4Ji+IVQOxUnaN0HxZeBMV
wRKee5gch0PwM197Mu1DUcDHKyxoUombUwrBivWGYDzNzMkY5ovII6hoYAPw4Ce4
wBo4vRIZKzDABvMBFlrHcI5nOICb06H/3TDr+7rnVW9S1+1ppRXWAV8h1FhUwZQS
P11nKIVZd9P1DnsBZHPp8TNpY7qvOFGHeqStoeJWWzDMT4OYvfRc6AC+ktn+PcDI
KoSdltxG4UdAr83LnrLb4dymdR0CSVOCOVN6QOe4VUl8yRP6Zs2aVdALMHnIJTIH
phaN4shZdP4AHkxXHHVwkdOZV3vCbYgtBObsXVMHv19gL/gQKjFaWH4t+jX+O1SD
Fa/GWiBJUCJtGP8oGmBkoyF9kqHOvXbid1yKqlUGhZTAXd32ofe9OyOUlsCZKJvP
LmgGHJtWSl3ERw8VvLJ1/p+e0gfNJfzAr6azk4PpuRUFZ8EAiI+hRvJYePP71f+o
RssPyeY8UgU2ZLPi7LuWO7+oP3aneBEY1dRycm/y4WzJ7HZaDehVPLApqXNQ/sH2
Au7bnzvvB/eSbdK5Bl8kKELBg+mVbUKICKBY1Myah32+AthwHNj6aqXzzucNKySZ
bu7jb6oVj7WODEHlhXriEAND6F4lYyJ79QmGbH+gwuMgH6A/LG7PiSVwz1P4dlio
NOneLA5bPHiad9/GkXsnkmme1GlfTApk133fyFReE/RuS0v99oM4c/gMFzMg3iK5
59/8iPKVv4l/03r897rXeomMcBvg3bGXpi4p7lorlSEoFmAF7lq9tPRPcU8uC2Op
EjTzHlwXBuOTf4gLxOX3R8wSwl+meuYIKmHXYnRsqwOCQTOETx/NnyM0BYHyXmTG
MNd1XJZETz79Pirw0GIIlRuXpBcXdWQ/nXs3LKt+krkO7VqDAxXkOWKHENeyWAzc
tspfZvzFdWZcw8oorX04Zk8s+Ut0aDeesCajX36R5wzl53zcV9LwQnfrCArPVS0L
5X6fw6kVHfkwigrtGxSb7fDd5suDEG33fRe/nmWri0dOHXDiaA/wTV/onLKfnoNu
CGoEgfTVzFC7UPoCcLvVhTR4nUET3v5LsjyPVL27IpfnyZ3vBggmNyRrlItQdlSr
jz0UDWLFqqFyVW7ieGkS5QBuRcbNRL3C/5lmjz6Tq/QItoFujQB9FWeMUu9CzU3i
gzQ8GKI3nn0azcBdkAkRgxqF+hZMwNgiC/aatNBV/SCFgkL+/rUE/bxlT6uZkTFd
mhYlgIEMsE4thAy44JJGTxcQ3VSb3FxzUsuEalXUJ9TcwwQGgdHgpXUfnOkdPsaR
qcYIwQxeH30B+QLjIZSv3/LZqUtZZlAzkYbOhBewVmrNtoco1tYjtcscUCGNuq21
Im4/o96fLQYpOkHxVdzb0542Ex8YUiXv/x0QfqtyoLS8KCCKwdySs6ltv99MrJyq
WHKsvzvRNaohlAdVe1C+IjocdT0/iuecP+0LoTHngkRHHEItmD8V4sxPtes6E/X/
29+mbs89PKCGPc2Z6+T1TFbapcv+1kMJqxWCZEtdP8je1VlTTi7nGO0j+sIpJEvN
sZ0eZYMWQ0Qq2R3i0VgrxwS7IKIB4U7BahWN/bOe9UB0bE1oOf4Om+ymLgimjqij
65wjwK6QmnodmdJRguEmAhWLslZbQ+48mU65+/1AldzTv+QNt2FdZiKlLFGspqRs
VVVmngsqzPnVMvUWG1rNPN5OD+mPvz0lDP/KH0VsCmYRjJTnjCLMVi8itV97sBkv
US8OSvcOXkJQsY+KYXM5nvBrxaJn2UobzWla5fkvX2J5XLZlDnjGUsJ9PnKtPmtM
5HJu2KX/+sja0ZMUkDPcCGqjdrGNpo978bPt0koQK3d4qhd+sUZ38jC8V6XyzCKy
gKDrI3SnXZHXovuNHiugmwi/1mBKLIBqGFArfHlznkxdEgQ6/7WF3woMXrsxKVfJ
pH7eyUgguANYesjsw0or0nCU1dyCNsFVpJ/i9ziN2fVbbqOASfAcFe8YmVtQ49gp
e7MmfwjfoJheqVzXwpcoRenc1CPNmiIpubT86+HKVjxXmrWrzYTagHizTzAaEP08
La17XvRMRudBeCq/qeCx53jQ6kDs80Rv6tX22XF9v/PWDto6/1JA7p9OrWa2689p
M/o+x1BzWoXN6R8zuqEe2tqnoiCOONkhJW0xvzwGtKSEAijN6owCn+OTtw72WDcp
J6pqs1UYxcUMDSeKJSWUyCgXrJpc18i8IOeEK3Y8QlH5EnNMej9Z3bXveynUH8nN
Mez0JcxqFi66tMezUSppa5YGhJGFvA5TD9Y63ZfSe5lVOg9m8C4RObjuQF9pLAjZ
QEVyV3WEvH4sSTuFGSUMTn829dDC/VBPWoLrH0iT/X6RVcf9U3OVgQFqrALVjXn4
ieLaatuEYtLyEvs20O1wvG83AJrqqLwLJhQKbdoa3kLjDoZEqcIjYpqtod/BgHPX
l4mkVqkKQASJauNnJKo5DgPo8b/RPtDHAE0whUpwdFulMcsWzyL1U9QOCNpXLu6Z
MIR2ECfN+ZMZxHxpMfTuS1873gH+444QMM6Zec203N64IsUU2DacaEp570YmoJ75
+7u/DEkm8LZUm9cSxJaPAkTICkni7DVJkIIGk6Uf9mL7El9k6MvvjkbdIK+AQZLo
sQbyULs0WE4fqZeaytbBihkuAWKzsOHXjga3RdIrHO9YcX35jW+fhulzL7ALiPBU
Zbh30a9nyaKpihy7rtD7jiT5if2TW2nwYieJbAWg4SJxmCpETz3c1pSvqHa5D+gE
hHssyjFGDXFy5k7Fe8dP+jPqrpTdkWLts3E5ltiqTTMiC1nCtqPDHWNVYUYxo9Wq
tN0oIAQOBSSc6/X/xlUvRL9Wm4m+alecIfP6LtE2cPtHDOMYE3e/qifun0oDosjd
Y/Oc1SkjfB47qz63a+N5EaNaoqMxUcZb+4kcAXHeKKJYjfvjHt6fyq8Bke7Zr1Wx
ZDZrm4L53MJlPupQZ8TPRpAh9yOXkWv/o3yg1+Pw1ZI4wkvoBtCt+7ldNN9MbdwD
56T9BU3D+/7mMp9upAn6kyKKVyxP6Nk3JKdGhAbxe5mSr15C7mwMrHipEnnVysm2
u7qqTiAavFfqshMHCWm8cNqrkF6oohQS4RzAn67UzgiBr8NrQFft81HHOLpTcs0j
13rcmcQMDYyBmEBflC5OhMs82uTUb6jgSc6ZI+vY0lqln14r/cMd2aF4LXZ03s4o
AInbXcLtAsdefFhatoCpaAzrywSHGaVbwK23rxYcSSrg7KP+SG8MEm+R9EG8CGsb
Vl3eoOrHXScj/E73Zk7a0GtdhBYqtwv3PzLmFOafkbZKDF30aXpcP7NLZWoDxIgk
ZxERYYT1FPaFBxRfT/zc4HqnTa4ej4Wqv62v6vBSl++aYWEvMA8Ml3aoG4LHzFBm
KrNK4VmPN2H00QkAOvzuvPWAjVHwhB6HT1gae+CvRQjYTYpzmTJuOw9LzAp8Pzrj
OtimPJpUeR4oa7w9PCbT58+wFUR4akIw1uq67C3AQ/qf1szoXGRdurgkcl7Vfof4
QCsNuEVNbMBhJEaveptteVHNlwRq3kwRcw6Wk2zkihlHrJONECY/E1oDfs4U6YOD
TdmQ7MiNtbsasyKSZOrMhqGlV0+z2N7GUQJzgGYk1T4L5n4hDOtgHdMUYHNXx5NV
dTJI4HadXNzxYe3XLXeWnC0wtE4bdJAd7sEIMuggP6VLwdHrKMLqxi6j2Nq/XYxO
HkRPCvSRhb17d0RxbXJMgy31pytLwOcDfWF98Ip6J3K8IBikviY0wZLstcwgR6Iu
UopFoO2VpBbOWqjwWMjO5dDaL+5x7G5CpqNzKALefgT3d/oSLAqV8sIIgq9WqIt9
R0AP3isxRr/rN9KiK6FCuY3pRj03c90YlP0sO9D2K5ObR7ySJyPhztSwXfTaEikh
Kg3M6F3ehuJtNKhJCZ3m79F1Z6+ARCKj2apO2pV0y7tdcpVbUu0RztHGc2RUFREd
O+kcXfv3nIIRi9aeNuoYWBkhaA62EIMlNB5Dail9YrI6TIeRcwf9AhDZ+H3SIlFi
WY0ExER8eh7dvgaX7Z+km3AA5KBd5lAfJG6L1FDYjxSBuvFpR7fTX1C8pAoHRKL1
zEPgDh8D+BMsSvqzWaaTEm+FyuPVPhmHivfLPkwOVCEr9kgIZkc/W6FtWsUfJHfb
e1f9/d1Jyw7DdSdR3IELgfJS+xVarHEZKE9qS7f/unJdmNKlNygcWYwrkcLrMR0P
ZnxjBiRG/aQJWXWxW0NouCFhRmidjZlsDBtHvOpkiLMgM6YWfNpzaqK0HCZmwXSl
V5nX1Rjwubpm4LKoojkLaYH31eV3XzLQiwHEX4T24Fh/gZtyh2rDJKAb9/lDWSQ6
w4hQE3ONRpDYNVV36yaVeTA58GwxQr16HrL/rVh7oGstwTdwUmuLIMaOlD807pFp
azurWQmQsdkqHfu8jCQ5zDH4o83cha757gSXUlgTThHUpxd/twUvlx9iBikajzTR
9843GRQJhgMn54SP4R3CDAUa6bRMX0nq7eNRt02zURtNBqjikDYq/Vd0ecxXKJAo
Hz9ZEUy3mbkki4cWhaTwllst9qLg4Lbo+P/B4Rw2pYI6fo4hxsssmsoPjwwKCQyk
ecKbkJrZD1F4hXSKNOuZJ0dHwfL5rXN+ryUyF2qQkNHswDvlgLd2NKEHPrhVXnAw
CMIWC5nMfhH7k4Cl4kJCHVKY+YkUuS6CHGsiMAo3lGcDhWObYTx8tlkuUjdSyBOi
p64FX5rZIBFKfHdJNgGsIY59VT7BkPJFFcxRsXv5fb6c9HXuI3knI7hZUpp9esAP
QnxqxR14Yv7H+CcbbUBcGSv31Z5/434HFx0o63WQAJiKsiJ8omIDb9Sh1Ax29qVw
xwqngQzg8LOH4oJM1J5hW4i6tEx0vewXDXb1Dg+JkUcpj49TCg1nzaWWxz6YumZY
PxpOxHBQ9El0HNYSTItONIV64AXjojBYzx42/x7q609be30V5clu1QXvevkP78kF
GqnsMNwnUDISGaFkuD1qDDOjLhJi2W7UhDBzVDZZRjeK81/s951NFfXjVJcisKe8
hnx0ITf8iQUqSK63SqSCkrEEoSFlZ8fEpMEuI4f98DhJ/bXfp1/B8cSkm7WpSo9+
8cYawoQa0Ynjq8fJMH54/KFa9bKtlLKr+OhR2Z96CaKq/ID48mV7qkHXSc4jOLcV
70CVchDjZIvrNFkXpD9V4VxSKOf4utIB6krfS3Oo/EWlrn5WnVGucR8Eo8JrYX9y
XmWn4p2D7tWih+LCZoYM0KDIO272LXYUAHdzN9AbDmZGgWIskQidsxj/GnUoRCC7
VB2x86JepQJAJXKAgyzm3c8bp3+2zrLdNepSLj0aS8KOX709HCVGL2sMU/KzoBBs
Qw7lLTWHPv5AQC3+MZTr9q3laiy+iyF1r4tzrW+ISZg3rSbnLr27ESpFLjIzXggW
/BYf9QVbufou/sceboDSZD6f2QtElKu/QNbtsO/WKZeI/Hwk7foP50TKk39dBNiW
Df+/dug/BWB7ZnqaBJJKyp+gEAnw2396OWgCHJlfBuDEQkCt9HmfaKDGllKRYsBg
IUFAWd1sJA9PCnFIpY5UgwJYxw95csZrP2cVCXWs++w6HZlJy5lVRu23eEgmUQhd
Sf9Ry55uzaXR+vLmL8Ii7h31CYyRdGwoV/VtMkCnVjkj6KuLIF4QVf7/PS5JZW7s
NgAQQ58mkk5CU/WcgZmLE8G+4rh9nWjKqa2TKeOTwZnsffhQMzVhduFAdROV08r9
2eN0whBJzl7WZE/CwxLqXuNuI2AbaZHJxgp41CS/PjS9Q1P1l0h0XoVdFtsmXWW0
9eZk0+l3tOwQ3ZVskU55F3jFXK0nqGUTJgHkePWBDIQWBoYYXJU1aKk4kG3qJ9mr
kQ1SR1WyL7C6XvuLsT4ZJZhEZodiFH2/Z2UN5Pyp6YRCqzdmQ4v4BH63VTiXIzzd
bUx8YnAX4VGabcXgwikZuvfaBzL7vP+ZfTxAMWcX0HtFF5qkU374nH7uLyPUeXN5
GzsCfQbZ/LYmswaWS1driPtcUlUfKJYUECWO0hgIyFAlxbeWFk3yl8icP+Hqb399
bWowgCgi4ja1ekQrxnc5jBfW/Gie7zOLfYbUKtoqZyPc6v4q0BvIbJ4vJgCx5jEx
VoEO+Bj1K8UL4IlEgUh7ubqCuKBtxsLJQhfXJ9aAuzxDa0ySbbjCbHOL253guJyU
BRCoufwEhmtUH7HRRoJgiLo9RsfljiUybU4QLmx+m7sfEqUA/an/Q17Z37px+wdi
Ewg5hztJUowSP+HS0g6d+nsN5y50etkUg6StSoc4X/IbwTExLiCoMr7zE4Kwz3/m
ZEd3BU/ERJ1v8RPZ2OWb2Loog4yiuEifJziutShOJz08jBRru3KKwBRvWv14Jd+j
eszchHCvXXZp4cu4eDTSkwx5L14Qu34ifQ2NsxPxdtycMP8PSnxiF5ugf24OI0Q+
HnZsrYHIqtgDtnqaC2FyLYnD8xiopwhApjtSjtC2AUSGfI6INnJwBstGCgYfJO1Z
IHOvg8tXoSOT2MRa+D/CnHl479GBKzHSNr8FhQJoPaY4XM9AJoCMvSnAof+IFwgS
muDwjXOfN6B/O9MEpNc3PwRg1T0YNcprRWtPEouF4naqyfdQHEo9olx3tUBZmdM6
OiOMooyRCTa1tl5frge/TAKGZ21IynOMtBZX0kPEoIW97VIsSr9mWsv9wWM9K4cl
t2mbPrFPQ4LKOJ4oRBLbSVWcsoFZmkprf7+KuqoGFJDgo0uCddMlU1NDbzi72LxQ
ofcB/cWMygGvY3JAeaAA8kaNCTnr3sJTIZPr3KvJa4ZGOhyYY8QT6KrMRb+JSwPM
Y9x8S0pP7mTpL/lB76hacf4r/SGV2d/ry5KOedtfkR77euPxx8yfb4nxj3FzpUhM
gxo6pkTxM7Qfm5aKaARbXeJ/s8GBwznZYgVJHdPGazdukdCO8vbrVE5KeREXbP35
EF28u3Qm6c0+R2hSke+A6Fh9jtOCkQzDtbbvo4YTQbn3NWsU1NjMNVHSJmH6oDPt
EkuCZNeXmkE7WgpE3gNZHt2vx5m3GT4GhctfNCD0hautFVx372Bps3VjORkZdeuf
UaM+cBiYxMlnzXGmqZ4DODyRUOQUZey0hrAQ+yn9+vCVuStqyoNWmqdkOOTZl3sc
X2m2VS1He87Jjp+3T7cqRVx1kSNnfZ9p7GD4B2QmUFJQSqit+6FTC5YIyfCv12bs
ACNzfSlyJre8YmrAnjoWTF3WAbn15HvBl70ka1xDDXWaPcV2nXfod/zyYvrRRb57
8dgVKh8uYxH7Yhef/bpjpRfAwiI6pxjCuKgc35r6EFJrUhZNNCnJIR2as1V+ukHZ
MG9R6X/Wj1vOIYABjX3EAPxSgtczBwtmMJuCBJw8pWWM1v0/fDAcqjPGIR43f2vg
7oudRgVudqXDnTdDbKegPv5uzuL04ijSD9vR9/CN1JCOmRh62X5YvJRAxLdF/xG4
aR6CAHgZsycl07kHV75naEUmb5nJKjWCRTMqMKxC3h+vTLcC55rBP6S5ZGtIS9ot
rI6GFSgIuZlqLOgmHljcg1D8POy2mSqdakdK1pye3lxIj49SWauoeP6oYLFzZu3u
8Npjj7EFPXreYJdzoSm3EghZ+f/jt8kqk4Eeopi9pJ0I3/WupT7UE4Y579nLcEWO
kYuYpv02gEsBeUNUhv6UP6FZY36cnWYiWT/3nb9jILnCJhTyvIq9PUQJoubBGfT0
A9gq/THdSTryg73KwOoi6E+yux7TYo77hzfysJCvbtob4D/E/eKJ9yNGWDhjQ6XK
PO2k09qJK9baaPiSinZsaK3mMp+y2aycEqHUYsWXTkhpKv/H1qyFDZsnK/280Zfc
41GJ278XSp+vqrgXRAnGZh6FEPYz5UE7XfOQa4WNu2q9yHY7HuuX7cRFVv3G3fQ+
C1IsKAmPJYisYSW1W5z9yKeCPROc5x7xznQo011f4nTPOYx7xTkI66X21jD3dSty
t834E1qpooeIxg0Mjz8fyE0dnpx9vy9RwW42iu/iaum5mGQFNA5TDLNTZWM0cryF
2NZXEhE+6q4hYpZsiRW0oGfxa41UBKTgBjlKTl7Tis8RFYiBUtdxIX3cDsykqnjP
6hSib4xxJraRVVaahS7bTpCWQoMQpFvrJ580a8OsQ9zijxzU8oRb0hY1m5ljeQzP
wVaZgyyxUc0HJDXtVuc8mvuO++TtdzhGOABtX9Qil+i+xR0ykmiPeUrufCsucd2+
Z1De60b9zlFY79b+aLnd77NKxKVkF166r6nQl5wRB/8Rp6gpCcu1YTDc1zea2O4j
ihqD5vcAo+7yGCjsK9c1ivnX+WSesLPvjQswGo5JJv5zrwD5SsxyPnlMUWTChk4F
8bFYHyxMw8DHp/yjFurYVCwuxxea8TYmlCR4yztqrQ/gVC8/ZJMBBx064E0W8BuK
Y21ocxkd2RT1zu72gQ6HNDq02UbmdEzEHacyyTNDtw+T5AOlAUj1EVCXX6ZxhBlm
QhVrCeQRfCZIaa50DqjMYAYYupN0pFpS997L7CPjyJlGiMMEqBAGD8vDZOLAoP6j
JwoGLCmzxDLesZHX2CSlAoobpXK1anAN+p6rqx9qA4Gudt4Hj3XTNFFPMN31J8gB
7a9s8exGiWiBjhopdNAh3qH9oqIWDS4cNv7YNPpFxduKty2DdFhsPkeD2ijTUWX0
GWaoa1JAJi/cAipNTz6JzAmIhYccZjFWVSAgw+I7cQEuadfv7gF6m3wst4ixel42
5ImgkyuvzfPZX/x33rhKO9HHAzinelBkf0sNGeozSJZ+OsD3wrr6rgHCRP62tjFo
KGwvL2em5NQ6/2edQiHFUSDU7YhsYO8D1dqqcO6RxYlYNYzd4hf6QOESzzkErT3H
yr5t2qbe+rNduHQ4LHcyldbmuFDkUQgx9wIk/LWdBCE50pZFJb12V6REVuXkGBrH
nzYKlsiX1IwxWYmk+bTHCMFndZSOaYYM5AYZWXP4b6f3spzzO2cZh5Rjxq3lJUqP
v1cvBFlwyvkFiFG3cA9i5yxWThdcG/fAYL7kuzVetZ2L9sXLz8EwWwPXn/UbAAev
vz3YnqGzR5hZ5F33VB0cND538BL6iMsb17iV2/88F45RlzBc9HGZKh9Z2zxRoHpy
lS6Ghtrj09Lz8Mv1M4xLmWEt+xsdBYw/bxVL9vYN8bHl8aWf9XNWHIKqOh4I2tCP
xTHnyk/n5QMsE4hjC7/kfOkDXsuQzFmt83FN93VEXa1FFEvEnYTM5XGTYIDL7ubB
89sTmSqWbROBHNyu6R9FyVkFyDwPbhgMbGx0u2IeGR6Kk7bsScp/P0JAM8wuXRwN
EYDIrltZC+i8AM9YRc4+7UeEeB2xLHBwrH/xgUR/xmrJ/PsWyT+D3Jb/BeqhOnZI
oC5Qb7IbCYXddLXOEDF2IcQUFDgXuNx9IRSoJVfYzfzv4ug7CHwNMymnjKXoThaJ
4lQaDaX6W8pjD3lTDu9Y/lFRh6ezeJDdTZPyOyGAp1BP8RaAOO/f4oP87yLB0Nb/
vE2m2sAm5g+xPVUsRMFVmXKb/uzv6gumcG+7I5WRIrRADjLJ0CaEvVvC2lbXBRtD
jIIL6Xbk5F3gGob0GjEL/HAwxYHqUsioBtsuwUHb5X56kumNnwXGNef1tHWKMylc
qktnsfTcfHSXsHco+YZu4DjsZPBlzawhtJwnPz84fwhg5zh6fpq8S5ylbB//TSR5
sD09IpYOYhw4ge4PpSfAtZ9H0Snpxg4QYF6bwH2kCHSYOJRD93cRWK7gbJHvMvRV
PIi3bNjHGCHRepzwb6wN+gBJO2B+XmhnIDFoDcan9B3LSp+tmYuggbzYbiP2fvlJ
ledtUvOmioG2mvewCaAwCU2quLnTW1pWqEvAdco7Zsl0/KVoKtpBW68YsFC3D9pz
zASwG4wMw7BXQrRyQIrZqV/5NaotPrkDq+ezK1RzJ6jBNLzibpKA1E/8RL8XWjmX
X7CpGvewtl8RU7UoGolSJRyAyAQfhZLBFh43Bpp0PTIEeT6dGot0KZYOZs3npuac
E+uiZP17leY1EbW9HMaKwSr1w0Dz6xHsyjAZH0fiTGnvGOd5FgJcPTyY4BzGy0Ma
nqZEAZJzLNzFjhqDIhSy/IkaBGvJKUtq2/b+NesuWSsHlSZsdM51tzhKj61LeuIw
HwXn5hYj8Wtvp+Dn37TjTpm3xKhZ3buYj3CowrE5QpSPuF1jqO1vRnujORqelyRv
vXI31gq0l6DH6w2yg6s6f8ysDTjistL3JdT/BnoR3o2CQq37uPibnsqTA8u1D+ld
IbYeCAgZ4Q/T2A7ardc8mdkA7L0vRzvoyJ2qTUxbhSkM0R7E4/8pdk/mcJXxIjUq
71yEmTQUX+FP/VGq7NFDhNNCheG9SHkE4LWo40hDOgxhK0C66zZFz0/XORGJDR23
J8pddNKgpVf0UDtjuMMgxXtZiTN1dbf0KIuVjZdJQOQ2OWcHJpRs0xBxKL8SYIWw
GexxFVMTPQ/Ug0JWWDN7BrgzotOm6oOt0qMLIFHZKUBPUeNVcHSSEgIQ71x0oEAh
I7AWyNvCeGk2JpxTAm/196yvUHtH/qoD03vmcxGToNGlutnjcS/xLreLvTxBdMAi
es33/HX2pqVxmw1hQ1gTG1AfvAq3Do+gHWwyXiEbgPZX6PQrGp5cQ2XdJb2BNFEK
j0gWupcFnHP6E8fZ/x21SPYXseE45R5UX+CmGrWJOWpF41WNND71hzDoOtV4Tv6x
qls98k97g+rNOFtGhQg0NyUITsAxJaQIYehiOYNsg5O4Vva+nSJOUCv2GgNLvQd2
81ut5iiP2SGnViiFaru8dLDNHmphY//AMuf56z3O2jVuTzDcMtzPUll2z7J9FRmH
7RdO0c83lzF7MxKbcNaBiBm6cyAWqxdll82ENVOLfdyc0aw+4lKhVAueYX9XdIkM
6o4fLPWYspMtgidqCs0tSXH5kC9D9IHxeHAHOEk8N8C1QZisWlE/ZgK4tqENiyac
NcZiHS4qbvW/LvrbJWMy1mJHnI/6xq996/wgxvR5VsP5WAA3QI3A02raTky4wmL7
0znx9daS7WHQUcKsifBSa1iSuE4mxhgy7pCIDkyC2p3AOUPBx3fF8XEadaCVjdX1
mNVZpiGViy0vznXAV+4oeJ012UWVOlLZDVi3poQswNQkkMDCiIYd46JA7VykvmrD
ye/U47xHI78abhwtiDETNeb2hi0LqVq5ySfSnMRh8oZ9FthkTZyKisaaSgah8mrZ
0jNnzBWK4aAMXrFeT7smLZxbzAKCd5ayuNTXbxUKIWU92k4Wx/RNroDDVnTR5zt5
RRbodPrte2hVr2R9r7x+TiL/C8WU21Zq0jUfde1acncWjo0gQiTm1PYjSyAyaB97
hZZZgj0dPtEHe7YbciX/jFyKG0d5eYou+1a8QDuWVNoBD0cAYqb302/SxHT7mlgR
k50ViFY91szs1ci2Cy16u2hGAcI5Whizf3E3qnCJSkA9eGX2dh//DXPxiy6e1EBY
HTDh+tBGurTyGOZzXCA9z8RkhaOygAIhmusRwiFzAOLtrhu837YnjIGi2JjMDMYs
+v5BIvPb+KImuKg15kPt3+7YqvDVDhn9HjcQoMnaRLfeQaPFKyXLPQb/4a7cyIku
oWySRYU8Tj3Scgdio17Ki3m8I9D2hdHlcEx6H+yeF0CJNeOkStEyNRE06Atx0YW1
vGYwuP/Ir/Rs5H08VZ6UVC0hGXzDVfNXA/nuTbtE5zFHnA7TtqrNxcO1qDvMBdop
bKyWXIjoqnHKNDC1o5/s05DyecN8UpKkgRKgYDvpJHMO3SH+SJzIBQ4V1pzE+YJZ
DW0Y4cFvTaoMhuAG0Lf/rUZrMVURuOp0yg+z2oTFCBy8c23ldePXQmUN2K7+TKeu
f0207wG3+SnYeSTb6jhBJWUHfQ397NB0WBvDB5//9ha2Nf/hBhiZzY8wxmXJT87a
PInIHQx7uULF9z/DujJFVA9lPcQqtz2SCdUsQCBwDY7XoZQQMo5EVhsHPJTdMdty
p0e/u9T6QIzN/BuTuD0fPLF6b7XQ4/ZAxVp7zFaQHsYenairDE8yQtIRi3rMUFvd
o7NuMj/2PuRxJHatJrghLRH5wRS8gqI65moMi4bQS1QdIC95iVLk3LOt273Ns+wR
dIPmYViVgtgChBLr9CSBv7vxCHz1zMB7h14h1ElEySIte8oly8pJOxRQ3Gh55QKx
c/ADcRefaZJHhmOMtKh1QkQwW4/+ZFQ5qNHfh4Fnl+ciHCYUKA7jWozU4W9nHVdW
/YC9LbaQESZIdzjaPxHfP1cds+usKx/yYUsbWKa+k/TjvVGwX+UL27wpJP+QA3gN
f++feMLfsZYEshSIPrULZxeD+/HgamO0AFEdxF9QIFIufrYS5qFcjyX2RUUX3I1J
XZlOjwh0yBY36z3v7f8Nw1yvlivDWiEJC3gL1IIm4SmsvrKxpcqIYOi13vqpjDbw
crEzkN/Eik0yUiVdy4U9cIuq9SrmcZssV/cyUIGyZ+Ny6fdkFRTcbcbiVA0/Ux/x
CVzgcxISEjMplLfJIDDZk3oT02lNzHKXPPniWtmteVvba7URRHb7DozLpZnIF29d
yCl0OrjGIohQMoWgtUA4JIcPf2+MkH/mrD/+q/lz8Fo3JEa4kxs088op+UmNLYma
orlnE5D3DDjz/DRILhb2uWR2CqmQcLmlmRaJiLfMlRW9zoRGf0RPoe5DGTv1ZjE4
gTRXVZ/l47RtZrWlBDbyhB4VMdgH69M7X0qbdHByvzVmocZ9XKDmYJcYp0OzcZos
E86flp+BLeA8opCl0j+S4DpYFWxuRnw/ktbwlKI9pN15DGDCEMnyBiOMXTP/8sqi
K8DpajEqfjHjji0rZn8chOOLqMyNkyhVZmRAGyaegLuKRsAv0eldzL+zeX5vivjp
sgze5hMy0NnUc+w9yEdws5QRN+CVYmZ1QgJspIdvI29HjNNymzzblUqX3ZeiKzQK
FXzwCgr0ZBYNcLvsZSVIy7iUD2Q51VaD2PrbI/xStI28SElVmKafwJXB9tkFVxON
Xiu9ZGZE4HKIk0r8Qbk2IXURoXhpzhOAb9pVkSTNM/ydqxFO5sEmXMxBkDr/FKPf
IHW1bYw6FsJ9L3+A3cGz2rvbtbx8K9ggiVCczN2rRsbsTa6AC9wSba0BYjX7W6ge
kItxTNbqCa/HXzJvXZPtkXIFu8/dWneSSr5US1x1B5B31eoMabiK91HcQbDh9/in
nDkqkwSB/tWpgMISKDviGC4eoVAsubopJwn7TGk064lLTPN5/xZjMqev9Nz7mkU/
xNeGWKr4uHksrGN2rzaSDU/C2AOU7yXFa9Dvxldh2F2JgRpdRahkAVBtggrPZtfZ
xctjBACxFDZpWEGYVSo29/+GobNPb4jIWE217dNEoXV4m6kVjGEiA5URJLQVer/t
9OtT9kpHvNbM8vbkj98AAgnttaIz9q3sNZtynuWWpk2r6b3qB597P1kkFE/sLeIh
lIJVusoENKpUZBwyxgtcUIi6J3I5AtIwh1dbM6LTalKAqh8kykz2PJpMFRoiNQW7
EtqsKBKEUK27ij4tqPWcx+uMQjXX5hT5bdYgJk1fWsQF2GnCpiBOKY/sGNJEe02Z
OtvHIEYaxRERp7/1OpBeKJ9FIz774gxPLArr9JhG38OSf1MmARdm3Oqo3d5fbGO7
/P5P2/1fCkK2EHgsdGy2JlSwOk6Q+GZRbLwAGwZqNHWper9NJ+qNDbfsOBI+uMst
fu4YbUurPCENwKl3EzYRkDh8/jtMq7MHi/yzj74ZnoX2DB9joKepo0UoLXkc9X3y
DRmMmPoABDEke89iA4O1ihh+joMNp6hpw/MkGB4D69kzsuGBJEFLeqzNlS8HxQaO
DWCBB0nEul3LFMTDt2b/WY8Tc0mD72mTUmL3yD4o9RPU+Mbj1WmFjhleGItGSVeO
YJzjNm1XUN/LC3N33gixQaBqwEKBHajdSgGE+JRjRIXBrdJtUb+Zg2nnue0I/MKV
Dlav45+yEnTOByH86EC4tq1LY8qhGSFRsBHXorTU49Noaybe702mjryJsr+cpbrV
INzI2WWA5j7HrJaa1E7zh/RaHcRompvM8LS/luaHfKexyJlxzJYW6tJY6YKr9F+J
tuHlYe9rdq95htTsYLKur++3QITQ8ciTEqwR6eOdmhYB0OjxCOkKpVJ6XE4PaWQt
Jss5sAz8xYDHDsipiZMxzupvTu84Zip33sq1mBSSl9yAproQqIXJmMLfFP3ddLf7
e1dyrOaSpooT1FPQmOeOuzRNVoFji0bVs5UzgF72l/AVCNvDaalO1rOeUc4fakB0
AGkl+TlWQGZ9/hvx4nt/Oy9HLpTZl53kMFR0i92q919+9OcmhBd2vwQc89skOpjq
it54isW3AdBxhd871PuZzVvGoyzplx5a65V0HaLRHAgSjkDzOomPuf3u1cH4i3Mt
8Y1nerNCNSuQbBNdWYvhVHAAKRFldYepRWWvlvY5Cgv8Z0ZyYBzFmj1i+ekWH2wl
MYjflQqHvVILUSNwFlRinG/aqJBSU0TF5Xxx+sGJcdU8bSxTG5LuS0EKKBn1XTi8
ESJrR+ADsj29EbTV3HGZ1LZQeb8cp5SDQqWOU/cFXcmNSTB8EhCGUx6ddyjp41uq
3Vorl/Zi91LrtDAWROkR++2ol/5zwqDG48ZcSGeqphMmyP+rEl30Fl8vlEFNp2LX
mOYcAgy7B3fe19vCZmSbZi9n4HOAbuEY7bE8BRowQIzK301zidhXx4SKcUzuGutL
WQwwlLxK6k9lbeQV0tIRbAkOBTEjodz9ta3MHwc3LjNxxTaq7Dtkdh5riXCdFVR0
gUJPSFKTEh+8OgJdsw0akns0nQDdyrScjIbvzKiIJa2o+mtAFyKHwmCwE3U+4jAq
EuEa5lCQTlP0YgzKzb9A6nDX/iFPYS+N3BVC+iFtVvTN2QS/dmnHSDCrtuVXCS27
M6pIkFcEknWRyG6Z5OEzFwsPZnaKxIY1ps0UdCH+aOD6X+Dr4Mz0w9sFX2Zq0kmt
xRmRZpHtNan8z5jG4AP9fois9r4czfdPs81kIcqQXf+plKguUrQHG7PzBgjAo2SM
UT7ujLxo8I0atNm4J1JuhqlvNAJqTT/Bh0j3lOQnk3E89tj+GVhcG/Z9xS7qfUlU
BqaqOqNrDG4wPoKt0PWXgXm5zA3ff4iHSqvieOwRc619T5CrwsOORY00hM7fmVtK
RNK3J+ZlRxcLsunfO0nBRzoSseWK6NCDbmWl7ddH7/TuxlSzju1nLUeCF6kD2mXY
THVdz7xtbi1iCDgHNhAJcHxjG4mG9FhGMrwNHp5159VxJmtAoUtL8XPfJ+SSDODj
p5UXTgus331A2SMrR1HJHF9VL8lFcK1r++uDwHPiLNtf4KHEgebevzon+6LOwiG4
4rWQUr7I6oOw34K8SfNrThuJZieLLMz4dOpX7R2zhCH6d5yyu9MpwQwblHC05zmJ
C9WRS5kwMorfwDxzBejbuMsYi5ZFjWR0A+5f4uBSRHhS/8VxGqS+DNdmAGVDPa39
agUKBtGRI+Ngd7HnsExdjT2Mp5GkIAHGJBJj4a7SlQPr5A5wTyUJvOwmQRGOmAFF
P9TklS9WYOGoN2+Y4YmoBjKlwG31x2BP2PgFYVMNkdZ9FFWcgXFU8l3ndq2Zb2UX
FwuEwpEzWyaoUF7GIGnSizKYCcoseSODL1VqLzmmluFNwLaCMeYxnonoBeLTBMkj
XxbPRb1YtFDlOBSO3lkUwONi5y0YFCpeHYrOaDVlq7ErggqzaHxIE79HEqYDVuWY
cAtLry2nKG1Cd1z+N1ftk36t0nVde2t2UwziH+bKQSbWVSJNGChD2n1sLDbu6roq
bXuSco2hKGaQhkNV5e1OAA/OnnLxC3awcYgilhgiLgCF2puVWvohB4BE0vyTAAVS
7yOLX9G7yT4syeMJM2sE0zW3mFmy0cXIS86cU8iccSS0MxfH2JNO7Pf9JcbvTvwB
1NAAINJOTQ8w6lpc+ZpDau6rhEzC/rR/5UGvdfj8topxBOW9DAN+i5r7tzAuMDTW
adbtEL5VY3zfx3N2RXN+MCqbqGpq9AZDfj6D93q2YVv8jJTDwzdMveE2y0eGKP/V
NYwartn/TesoPwVNRId3xpjRMWr5EyyR/RLKv9AsqBrihdOMBrqboKai+SjTA6Z7
gjyDAHuWHqu+f3HfqGkElz+unlJtjMGQR/qa6BrSPqOVwkoj7AUB5iYwSe+h83wY
Bv4j5NxypRsi0W9cxU3zYWIlqY+7xoShnsmRYvByNzklG7umMFVuVNhycgMWMLgx
XKa8nKtukeR+/am2bSDMUsUjxzMaIXN2VVCS3ZUARNOjW4dlFnlrY/L6APx0p05K
fAzMWOYY8LwQUV4I0WONPpuFjsA2m9GrdY2eKOBU/QD66guiN1ZXC0ydfgJYtkan
B8b4Nm/EPV8wSfzk4NnTMpsVnwzqXYjLNrrWCivtrXVPdZ55Ig80338FllPxsQzi
FTDQF49PE4KGYGC/pFvhhndvcCf5YcETnifpYBBPoyNMO0XcUdi2JBQi5Q7UX8M4
oYw48mAY9EwQcncIJFv5H2z19JaebdOqZi1GKmF41HGQqKHGFO68sAabHFoG52fR
j/OcCC2FXsHBaR72n5ukPCoEuu9WK3cR+J1x87T1LY1sZwm27Nsg5Gj/ko6I3mlI
SGOnrHXmV85iCK9yfFmIDQVxQ8A5ssiws/YTtoIV1qNX7fijvYcsNNYTAaqGr5qY
3oHEmIISgIQ7mPtLjalGLl74d/Dv59vFwRoKWcrw/vXmWzIaOXi6JACbCq2Y7zgh
hBSF9BKzQTDR+k3pbtDcxJxvYOVG+sengJQaEh1xQsdc26kYTRZ1qvrYeDay3xlV
wgePwWdiwXSkEWQ64ka4ryD7fq7R5AOQTQBxRYfrn+15OKUMPOswXw8b41PmIRHu
O0r7bDQ/xV1vQdSSOrle8OAuCd7Fxt/ah1w8zvvaX8UtMLgjjGPqTnHt/N/1efWX
s7WeXD54L3VJ7T6W2a7tpLHn6z/RvP/lAaKpIZcpu31egyWhYWTdOLektKFcynEq
Mj0gfuOMueG889uLfvD4uJIzW8yvSVT0j0BqU0YY8WLQo/5HQWPGKWAMWs5RCWSz
fx7vJKzfktzJs8UY93yAPV7ZnFBIOBNIBTJzdRGeSYk+rnUrWteh6xRShswLX3SY
U92CyS85J92NzX8wiv7pDPBwrUDVJsVzM5BqdVOXMl8rNMlIk+SK71/Xke1MV6LH
KTRIoyBxGdHnfbgIniAQ8wiv2tGgfPzMc4kchLGjazVnS7nHMoGQbZPC41A3l+r4
8FDbLdaNhhsBBFo0SLBr0L1VodRiwe/VgNPLMb8iPPfc/yD5CVXO6jY++CLPZV/5
kIEU9fACWyG2Q2IXY8dQNIXe+LiHnF2FbIlZrIrGxi4/XzwXI/GO0JdjfBNbPfJu
wFNIgfEKdpN+jH+PntEnNOIn8z2N74sijK/ZO0fOcubfJIUZGrucP7gdu+54Vb9m
HYfzSUD3Pu7C2c+6c2y6KhKD5fvhvthGTmMVoLs0x+rS2uF/XumOrKjR2Ebhpw4x
xGHcxxA0s72xgtFxoBBsIPdv9nd1gkFgVey+pBo3LgmDwJUJAzdgtFNkFxdGOvjq
BPeqNkGA6+ohUE4ecnKxG0NKjPum09Jzw7SavjwtSvhTzOPC5Eo/v1mvleIY6dak
YOTngOA+7+wsXkYGKNGJ6i/SYd13CxGMbvZv60Atz6J/rCTpx9TV7YEaGVyHTOpl
ICHR3ZCYTRFoMm6KtomrTEZzwBMAO/nhnXNZ5S2eEIIbL09Z3ikMfVDO0/DiaV3H
O508NgbBiGRVOgcPl5ReXwBgnFiffiGL+su3fII5zDiFiHDV3A/2Gsvn29uN8Gpw
YQhhkTDPYjs3CCTDoKbWWtGzqFmOeoBL/J8F7eQsUu17M9rn7MGa6qBFYuR9ZZe/
jfZL0rjiaP/bVWcAS/DrRvVpP79XEAgu6JbVjCZjMHJBK5LaJsIUw4FeaOI+RZkk
9o33xvPvr55cPNvAeenTAEV+EHmXB/RXc58/ZIuqyqw1cT94i53ODd5NSECXYvEY
zE3FB8Ag8OFt4Vvxlfx57kV9UANe+82e7oCQJIGGBG299fIKn+uKG6ltdZzI67u3
8p+C0xtpqvNDleC1agoQvFz6s2zjlXLdejp0KTstCep3siVh3sbNQ3lBhBt5XrBy
dXGPPwYa/vELXdRIXyxHbMdDoCLj98AvXnPJfAF+hR8zwlww1m8kdeJMko5cbM+k
cLLJe5kZQROseFtFavn8VMNRgvLDIawxTGEa2YoD3rR6ZOghr/FN6xF1SuY3RCjn
oSzKKWsrNVCH9KLeQ6CbrSGtjHLceP5YHFQYui8gOh+79O+Dv8A6lT2N5gl6mH9f
BL65D5QUVn/DJNM2oxUmL0wKfe1NtsihywjXSFGDKCRqms/p248AR0LOEo/M1sDc
oR6V1xDmbL5oR6ukpdg+NdrtOoO95eJDSzW+xltvlrvzpEv3FNm5jihLapf+XvEL
aPbGI930xyhaDIK5Ge5mrxZgf1WlKcgnRX1L9jvU03oAf/J3awD9rbNZJ3G9umFz
JNDYmpQFDFxcA3Qii2qCtzEXT+MIaHZEf8wOj50tvXlzu9N7NWeqEN4WSvchacCB
6LyYpMc8v6uexuzG83lUg0npQwXCNo7gHO7YIrSzTNXVeCEg3y3l0vohuqpiAmsL
BW13aI2/O8JzbY0z0Dc2U28/KV+lGBnDrc2nWyHWVWiqVk/F53MH+SSpY9PvxVXq
euiEbFUvNf3tMY3TEltd7+cjiGgBO+YWDiXMAUSlencZGYzxEX3fi9E3CPMGNEBw
Lr+v8eID4peXONM6aD7gTxVWQIKdg5Q1kXuNGiFJyv5WOSY74xj6NX23fxC5hsTv
Bf2imyJwVB/b5hhWffQWc1jxuUdAlf5AUlTxCGXggwIYefpor5UMe9ZtBB6V5qoD
6Fb+q9cTTJNINVN7y9Whd/I0YFfFdJheHoUIFrGKvun3B1sutowYn456aEXsfbZb
fW0iqfoCvDhOz8Mv0z5P/GHJghQb4W6hyrCFkUXxU6e6LT4k1CK9+XqG925u4hLS
qASRHED76CVjE2mNZ11RuX5Zw9yKhoXsHLadrCC16i+ftNDZtHS5eBK0PMWqCck7
GnOV3884K6Ey0nCHSXqZhV1H1mmTyVmqprNx/URHAgstoa1RLvv618v5zCYINqTT
A4tACdpd9HPA1oC7E8BeEPdg3r2x5AbQ9QlxPqJPWhycShbuH0Vo19SIqmuTakIP
UQXjifybV9D0OECNEQhaI1K6+702gCMjCRULbnNrBkAPyI9MbmomH3w2yGPbw1vx
GGgbokaWxavBCeYxCtycpbF1UDKTwZSghxvmmqXkz1giwwZdP8I27Xdz3l9IvGD/
6dIyTfPM4OCVLyOVMe1EHCHr9h3lhme/EVmYWO9g7VCF3kiLk35va3tKDS3VHeap
Gi6d5lyBP30QzxejSmt29a9GEVBio6o4ObXqGvspJDzgKh0Fc1xwKFRq8k5C8Edw
Xcp6orc6/zxSWVdac3ewCrLPn7PnRj4FnJVuy6/IZMmc1udMrQqKPiRVbIhlK8N1
sjg5+nTMPOFh5gdgSdHmECIWPzNmKtXyxpn0dnTta55lfCddIPUbd23QqMyHBP1h
C4F2LuI1WpMtCbN+Iz98C2IPuK0DqMP1pBC0qjY+ibS4Wl2AcAUFIIjJZwU2Nrbj
VouyS7aNkGU9q2E6/IGux8+gfGwGLpokwgmRl7bU0+VcxxVqDgwXhscm2TTj96Jx
L7eEeG1NBt3KruVrq9VusoQzYR3qPJqL70y6TwRnuYRwQs5KRfD7lbdYOQmsBCpn
pfYgTH2HI8QCu6QREfAhTOeWrjxhh4WbFuhIDGSbFRkjeKq6IS8Vs80TATmcIWTo
UgODKp+Yo9fz6qqD8QJ8aR293JVorv4mUrjmYyhW4e8EnylNaAA0sxbOadYxdwL2
KQVnomB46vyRVDxCLYhUkodbM7parOAw9GaFjvGWYKgcHDgzV9mjHEZ+1JXO1i6Z
urCj6ijnTh1YbC0ALJdxHa0rypQi7Kk3nRrT+yXtCCX3rytrRZNLu/ZoUEuq7Ltz
rgKQ2gIqeW9NRcFTpclqxayfBtVMsaAs7APunOxzR27eTX2PUPRyt6fYzBrAZ7/Z
g7+BfxOKpNsPfBAUwnqZN7qn9c5fZQ14Gczr7qVtKKivJe56pUXw+nU5D1o9vxfJ
Vw6F/A/3FypP0+fFoUjw2q3/sbLjtpQqn1Nb5F00ezNcDkqa0SBUmqp7NJjeB5SD
2T8IqD88JD5+wc2DuLzWU3Vj0IYaakjisBpJsmM6ammqtZVfXz8YPZTA1aLRopyh
2DcPTUniqW69lM0H3sSSXaSsUT5W1Id4ceurzKy4iYX7FG7wRrXgZjtQFCcnaqC1
3UXaEFD36S7YIA/JkmfKtyAVv/RskCdjiSAzu+MOx1d3O5b7O2snETWOJNWLXxoH
GlHTJWL98qWVQifIyIqwtWZSqupRAsTCjDZYbQL0ppH0JGEbwiSFtPKyDLeuHEYK
lx4Fnyj7Ts4cBAZhF6igmiGgxU4gJoa+qcsYEnvXn+tpB6oDjO4+3s7uTUNR8qwD
ckrEftTdWuDQgXu1wY9uCmmCtGgn27go1M95vBl+o3Z0supRrEZwRlQuUZbX8ZGq
QjC+EwcxHnWrVAY51pH4Kb64ntF2TAFd2TgnRH9QuidCkgzhs119KYIeEfG8HrVe
GNMWVFaiM5t1IVYk/MD/H7pyYSaxK7hzRsudt14JpVGDVL/r45p9qNyaPXiyZw2w
1F9RSd8h66fOs3EIAXHcgS2RsihTeaOg2RDGS/9k5SQD8fNwwpfNOFqsE/pFqJh+
vmigW/PpG7oUicetYYi2nV1kuvxba9SfXno8s2cnQQAbDAXdGCjjYxc5zSTDZLsp
k4NHANM/wmeCo1TeuPwZerF2gaV74kbPcEFitoSymi2rgtiLSUqfghGIugBOiSFl
m/kDC57t2u6SBdun0ve90dfpJUKRBcBS7egUDYreIbI1LRiaqdtxwW5ok60l/r+D
nfLvxp2L5Ua13q24r1z7PpJaiUnI+4cz/GbT27uWy9TYWeR5K4DuLfXqEvv2p/Qt
z909dX8PUdyn9FobU7ribQ5a5CCzF304cIvqZLJMKIlqfeEeQvpahKASrD7qXgAt
3HMAFk5A27vAlIvkZE+muUdjx4dN5FQLjVq+kkF4wB/JfLan7WjGSQgZFy9bh7x4
wrQXo1DCHxClhh1mfUSCXhOG9iCWZtSoSQwEvo54P8TaA2JXdlogLFJOVtGCjvvS
yTwbia6BHoadp4c9dzS5XbnLAhZ6Ui9CLKA3kj0ABT0k4n2q9pkQ4SGPV3g7yO8r
H7E7A5VK24CnrxAwoacItpPZmildFBbrHcLQ2A7y8vv44FBNBVNbFnw2KUsJrZ62
0tGart+QYmH5kix7fkbHV59U3E1XhYqS1GtiXotEXSpV5AiqJ0cITzp2dSELGf4c
g7+exK9mrUukIvz6l/SF7pUqhUYKz/4inhRdrznJlGK0XIvmZDJdJm9au1ta261g
zugGk0EuldRMOmSiCEUpkFNUfeEXU2NmZZIrQx8muripqLHWcEzumiPW/sEr8ENW
dGTuygp4OgAVOd9DO/0D7CbGewZ5+BNo9NfuqD/DrIB54IwCmH9YCu6R7E1YyydX
qwwIS2xfEwaMOs4eV+JYTPEv/Xd6oHxAxvWzhCzX25SoFU6i6kAdRJindOG3egWV
dV/pHVMS3rKgQojynBYdUh2O+fLYSws59LUspOeiA6VdwuSipXT0k+Rj9ROeYON3
U9TiujmQTI/tacK7IuyeDDwc+iaj4RHI3ft4MgXnOAwlBQM0VVN3vrmPgE4gp8D0
d0GzhpWucSwwNgEwRyh7jRxaCxCAk3f6bYz9rflqx2ebAAYrUj8TzvKGwpzQXw39
bpaqygZslLu9cAchoFay0+H36Ktf16ZzXrsAlTun+ik6aGONhH20+4yyudmM4Vf+
wUgMo1LrvTxYAFzvvRGIxpq516S+4rNfXrlYCwoHz5ekJ70voCj1hP8dc5VoxLNA
zLJ/4CbL5wyXRmH5B95IK8R7m9VYqikG62F3om/tr8Q4+A3GfdH9mz1Qh7rzfn5R
99MtsUW3pH3wiOxElzbLYyBfNhuxgqDF/x34lMIDhNtipGdOosbQLUe8WqlVVUlR
1dqz7jGMykRktXBMRBBPA85n+EnnWkGFiZr1UQK2w3kyrUX38HJJksCLHI2SivRn
KalTBgxq30fUzOGeouws/A5Hg+c/xglwSzI/c0jfWX7bT4spOuckaQ0fv5eKHSWD
Pb+nf/smaFxhWny7b4pf7v5h/hPrpSxiFY8JTnlVyORv46fXt/7BtjiV+b24l+6k
9MPlWvV/xGIfNuuPzDEMXghzVvV4E2jElJycWxRIEnZYIsL/qxie1fyEaz258VBm
xDxKceOiRiAckJSwduQLVK8/qkCbbCGUfwcxTjl4DfgP+IV9iojXsnsaGTXjHH/c
WDWXCD+wZygu+pTyO8nvPadiRNs6KC/qT35I+ckRszrO8YKeKN4DEbPDbcddixsm
3ka8Z4bLSNQ/WAOoiI8d1AB4bgZJcqRqaAHKFsZyQtoQoz2kakaAKmfQ6S7296ak
mFoDDNeFounORUHNc+PCQ+4TW3blEbwnyNHoBo0WJC953jMzx2FhT7l8RqAny8ra
EKR41xvOsYbQ8wvWNMTkby/NtXnWjvy7zS8dmhaBFKtsReFrMw/z01M1VFrL91CJ
Gavp1/9ohePsgIoJKt+uB97v+480sIwxHJ8rWGfN8bV1/mZch66M1/sOhnh0BHg1
795n0TuPeElnzGFoFVSqwJWvKPh847onbN0hQgErIHXkROMV5XHSmrCXmn9iMHRA
Jqv7mt0to4Zh9aR/YlYzuJDv13vMkyLnoQSqNLsE5t3cnp9HUQK41qQXzWpp6hL8
7+6Kf+2QD24NBPTOas5fUFcj3MdEQeG0l1Op4bbT1bOcQ4phNQw39GXlNlLIMSCg
qtQ1ZDbWJOvmkpNKM3Ls9v2Lvks0ba1QZsY+SrKKWlIGP3zdVRIdm06Ltb4uTYBt
sQ5y2NKQWZFJGQhzlVvYbY1ZDIBGKfocBVPgLErtKIWF9YzWgI0HWQ03VJTbIbom
WyaQ319vNsDh4+vYy5EqhOLep82rWNPjPS2MKxmsyB6qVHCJfjarrZNbCaduHrLJ
GmqLAmx4GNQL1lwp5hbWuOM4TTnLomtzB8cfctik7pH0UMFi0WSSsDKbTWjlURrI
bVSeHOk/NSr8CquTQXBP2yGPrKSebDvQGdQxs6WKEbbyR6/GxIhw3toEFmQG3TB3
RZKcNmP4o8yKsqv5cb0wObnynuDvmDiVubSHwHVzO9ZpvZUCmcEeorsAUaxdSxC7
90vZhUKAsjrOEGcCqrH9WEf/DJug3J7XzXfbWjUIgxgdEWa9T58SI1NqPx+TPQzD
Z9iYn7J7nLKWYdLbJy2DHUJpT0Cpmz/M9TvqD5C71IuxzNFO373DmlKCam8v5SnY
SnIqH3FDEi0bP4h827UdpZBL5dhuubEJWyBAqWEAVKYH5Q0EK/EjYiFjfOiNYZHK
Q//M6j9PJ++bVmV3ZO1t3qXnrbkX1XSagj/lAv5JDdKdLRjaspmgiVPRg/bBvNQp
0k/51V9WhJO8hnp+6oohgnkScd09aYCVaacsVh42G6Fx40St23QkRs0sIHsIHpRH
lCPX+h+BxZ9Z8EA/+00X5x8QpZQkUNW79mxyPULxDA5MYlePCI8Ko9aVmHqBc42I
v8CpCddzUxGID2eDrVzYI59u9E2TPd/jvNP73Qib/ELWmTSadkaEt0Q+UpGjk4Ez
GwN/MjCr9gcUqlEfiIuhwlz+gu0/Fh9T1IRuSZ5T8QthsFfRb7lCBqaVkbArrgR0
hqCtKDGBcH5YJ9eLhbSNHOslGsf3IVGF1Zi5FuuPbcbkUvUTCFN6rLeSewHfCJyv
5BKneKfkIYETqZahTn38GYUXSCLynANtWaw0qOj2K7GnyuUZ4eLNWKUZk1vv16vu
2eRnlJ4XSuzJ7g43+Ra8lUXrO2klJgTXYWM9dMeU23LArWFw+Z5/O1FwnziOcTNh
5uZ2dPNCaCDv4jsu/vIAo1G+fxzfrnIS2UZ6H2lZ9sXwTPf9vvZbagc+6Y3iFLnK
2NmIHHo+d0Y0GZyyFlLof6ERbhVGo42TXytXciuAT+gbfSEqqDn1vc7gmMtNSqmj
eRJAN+P97NbvNLYUb1e+O/ISkbF+sOK6oVxoFVnJqr6PpgRNxDKKTFWlXmlnD/VS
AyZOgBI5XRe+yhG2JFGG4iy6Kyy7vvxfrUzh07W1gIFjF8iXAUxRACL/yUf8xTn/
WdOhOHyVw7WO7JN2rP51rIrGNVNRLZDarLwn8cEn9SEaFsMi37mBlOZKOV+W8btB
K/2ops1SOVx3CkOHeXSf3s/RAJ27BoHKco5f/GiHlK0AMhemcluyoCYjrucuVBmC
DLPIgEQmTu7ZIsR4ZwbZPrms7dVRl/D8nmRI/602RXeKBgB5H9vOlLQXIabJX9gj
vMzPb8li+E0FgNS6oiYLCPP4ATwic6j98Y4Mg0KEgAejRSrAap1DdY66u8Gwfbm0
06yGgy+2WTZXBKZ9p0t8S/amNZ29Swkw/E28KJgDCyFnMLrSixcbLVQmyObzcioS
Ji8bU0cZsFLjp62od6j8jnhUoIz6pioFwRu6Rvuu+nLelbo82pgSIOqaxt973BkI
qd63ZJ/fcA2nMbLAVpQ0r4id+6GUgiqCt43GyC+IXKOobW7b3AevNRsE1gHbEGsL
RRGNAV793uvTUxmAyl8I1GYQqUwdz+oxQJnjwW096ip+Ya1IQV8iP4t2uFq7eQWT
vsZdJpZvgxGao6ud+3U9TSDFpVKY6OermOriaYP/02h+Mif54+lYGNRE7A8P+w+7
wDecXHbWEQIEpcv7LjzYp7qs6eTKBweM+PNmVojj82ejJZTvQ3hEeeZ4mLVpP+6v
MrNhv7TICHkkIiyOEwKBMcE2HbBc92Qx7X8P1bf1uNiMoPNHvLWYVko8QDqJpAzG
lelUwig1kZWrI1GGF1rdi+Z3kUcJbZrYM9Vaizfnc451Vv7HT16kd2RTCNbJ4b3/
czjEqLzvnruVNDx4vmxSKK0quC99sZGW5YFf0LLC9d9nnHEymDwNWm8dt7ys08fV
bgXS65pZuu/xhPpzNQD46s2UV9vMUouVqHifMXFTQrDh4hsY2dEiKWEoOeQMEzoq
hc8NPDcl05nLW5e/W9yi4HgltxkJspZagZuIxfkzYHdmkHA5jivJhq2vniA5CgBg
j70UlrwbLPWd7C5pSHDHPYWEKyCIds4C0RkMpz8CEtVB75Ii8HqEGpURd89pUu9n
weuWP05kl6lsPqVXlvQuj2gB60PGntVUk8/qQ9uU6yBCCxF12TE7sIYNhliCp7HG
9ogBTQaIzZQsTewhBQueI/sfg/3T18ez/cCDl/a4/MT7m4ssZa5YsIdyLHs8xXaX
7NWmiRDraxWL4/4Eb9N2mJyDWHp7TS636izPDMk2Y1kV8H+qNIPYEQhAhM1YgA5J
omqslM4+iAqt8rt3PKIKSoYT+7aZXKN2loavKyFu19ix+aQWSEr3+t8BmI9XlL8E
UIuklzqYHJ9STbjo4yuq321yHykQ24yCU5TSXq4iP4axwNAmYt317zTVxCxEW11k
zzG5thwplc9prayJxdhSaXpqDlxlMyfm7NVwLcrPGKqwMKuEO+Hfh7iNgguW19ps
7ZhZ/jDfEbqcUh0l+6l2y3tJBVXKeXDMNOXVY9dCwTz72rf/XabfpTTXdeH0Xppb
c7K6hi3dPciAx5sbEy24/ElOgItDqJ73Zp0N4ueOTdpr2TILDXaHV+0wOc5r+B58
g0vjbRB+gZpJCXhdMa9XDH/v6u9nzyYePeURbTpTG08Y5HCqtDibSyJDUE7E+aOL
xUc7xDmPHTCksh5y+Q8taYsJKhLtdAw5671TjSJiDlGr4VOBPl56Wp13ZeGMU+W3
pn9I3/7PWoF6CRSknthvIVuN6SCnn0VQyywFF8g11n0udjZN0DtgIS+ezuqXsrYU
eIxiA2w5KerCRg2jLCb9YH7adOFYQx0Ycol2v49260gQ3gOneHQowcS2Y/9163f+
0Hr7vwctQoCWcaB/gGsQFQDTHMEWzSh4/gMStG9Wo//591IBEylYOLlaLisaqz03
fULJXQIe0yLTjaiihR/66jZQhhWjhXBgWQAvVC+LlsFx0zHspQyDHK7066QSUSkx
qDpLPEsni8semz1CKco2pRmIkJWLxutnVuhK+v6d3u1a485npSc97oMrS0M6QWlO
gVlRUqRaDNFqJVt2G+IK6es0+cipqxBBfK9GT5N6EP5kZD+lPyziBa5vEBkrk62d
AID2xoIHCAfdgXcmGRGisXDkmpi4AFjL0yPZ5tnyTvcPZF6UrFZNyvQacrlkVOsQ
WKeFFhg4uuqhS/EBcbkMZPe1r1+T5Gww0rQafYHmZkomGIWKaFMWNqrFuy1P9Yca
gfGsu9fmo0Oi+dW9OIEt4LEXbNznXmxCZH9tATloQv9ONYPmGcfxlT3KSPVl1pPK
kLjfi5eDOK8PYPv2YaYkhhJI74QbUSAnaUwRyck6jgfi7yYmMDx/Gh0i/qMndkgD
B0yO3ohRReqtWd+6R4kBH+pvaBajlH8xwXPj8T2gT+MtCit/3QS1b0X3Jdu4KkQi
24gaAIe6JrmBBx5RzyMvVj9ZMJfRYw+xoZNkLdz7u2RLVEAyUZkftP3gsY8OTXYI
tBiZPX59mzbPSYdHEGa22dikSUUoCeE34ntXxkLTbBAoogoimq7IN6HmJ+H/dvLZ
lwFOnm36yO1lA1mRRO6dkzdR2EbeXwSHhr+1Hn6Rzd9/Y/rGWbW7P/Dve0br0PdT
d3Vjz5AOgyx+lHaKnHpUmOxbz7NsCLmJnfzBNhMgwS82nQ7v2y1GgumTj+syJ9mg
Azze4QQh7EzgdiOYNa9dbWRTDoMOgxZ5xjstkoFbDSF18IQ0alL3KE/wh7qZ1JxY
ZWWrGWZDHCp3xFMNdbL8jc+iZ1VAdwZU6tuyhdB1iceIVMjXGCbOrHZ9dBrIXO7c
fIpSsSfgQ8SRWX9hfySXysYldQXgq2Lv+BOlZZMScw9Rk4PUJR/NP6QYSQulDGOm
4kvkx1haBbgS068MvBYe8DiLslvX7oyT2QBQhLFwsSTfecOG5wxB3Zc4i260zrS7
3oBu4Mi+TlW3rwduEO+3mc59JFuUlwsoVuE109dKX/sraKA9nU8ghkVROnk6SIEz
j54zbox42PVt6T2amU1mfMiRVB3AJgTxgS3ac8ciotEcRIisP4Zphd0Xf6twbL3t
jmu2sQRs+LIHK53Hkuy5IZwolnw2VpYhGWVpmtYfuYiDjkGCNOVuxggon0p9547V
6kFiOPraB9Qs2TNYhE1lQ730gxem0h9JaJ48ASz/sEn3KnoZYWThWAc8bOorJ/pw
GX4l+kzPS1RnR3YNcKycJbCSmQowIGq45QkamsC5yI/IwNoHKCzqV/n7F8AIxOtu
TOsEm/I2GYDxCX0JpdvAu2+9rICyF5tzy/pFsC1t2d3DOGWCLjBpyKGhryDhoulc
vvghf9+bHtlhCKrLN2Z6J7LYn6sOP3Bm+2CrFxaIIbx1Z7+ylLpVfgUcu4oF96vt
qXzFjhLhq3XGjeZ8mDiO1PldHHIezhYUlXtAmK4RC/O+lsAqlPS0Bn6Pcs7uctR5
PI3mBi9yxJwqxY1NflIgoQ3Eh8wF/5fSI7Fk+4GzZOckBj3WtaJo3miQvF+OZbGj
wtBtcfqdr/mvzkS3NlXsbSWorPrraIN/BFk7Hi4bc9CB0u9icYKtzeFcBduSTAmW
UVYwFS/LPR4TM8dsZlJBvo4KLLa3Dy8aEMoUr2RwXrJUEkby+yPY2xV35w/8b68S
qLudptuuy/iRyx5U+hmh/zI2M9v8H2jqDMJeHGNtGTGgjE88ddZGbR/atC9sL1TX
ahnNKnslRgsN/X9oeMJZ90jTGFFqdwuV/TkvX2pCaSQNdaimGK0yrdhfZZBbotdu
qXMcfHRvBk7DobaYEkjtZkYi0NukLS0ErVgGZfxC3/VmoMwZN4sdZl1KCwNjUhtR
D/1Wl0+Ta+JiNg0kX8yTY6V0+ulHBfVinCWqUpVGt5tbpNuIf9laRHG+NMeo4o+L
GNSBJ70sH2ljJuo042WBKVbdvCEjcMQSpBkdSIh1Z8AjzsEjl0yj6KI9EnR7xoPm
ZZ4feV9b13fg3dy2tuiOURIIMSmF+z4EfYlu/lTPIqbZVncfM3DLa/JOV8PdYE5O
9M+SpfBWA/xTsKVedKsa1h0rluSNdB/pULzn/mmxwvI7D4jDVSsfzG7dHWQAZ7+j
AsPlM0gShhR4SVehXQaPd7igwxpG6v5mhm/c7bkSPPvvKhSWPj/sfSkJGojTFMKr
2vqhyjzWATpgt4r6IzTy768werhPK0lc9UeyfCFKZrR5dCqL5qRI8zLPX1t/vG1c
NAQiaTZ25hruvwC2925o9m7SKYdtl6qByxGPMSVrAg804WOOge/3rY2pUKncmJyo
msbxo6qtZ/wymJjkYeaI+7iMdNbWSOzwEzU5xzA6UdBliTnML73JbqKx2LHqyJNb
jE0rfuyJpZLZ+/cBpvYcU962q4GNIne4rx+MQo5bgeq9nZbpwV8Gh/P+JLSxNuoK
oP1jAlB9m+u1AizEIJnky/bpErQ3n8iZtw07w9t+d1T16c3DQHQ8ZeYqYpavIYPt
oZTISEhCntOd3Ho6TtM3f8WQtuYZAlDQbJKmF/h0xxZ4k+kF+r3tJx961isdLxlZ
nU3lvk0MvyZ7RWlzHU7DKYVHPSc6+4fZrPZcgdC2be+TcZShzuiWlla2Mw6WkJod
uQMW3AwkM/efuMt3JdeErK4ZA4acWyQgVnOlOPGa03bhyZMIcItgxHxVf+tZzoAJ
knznjWFwIzRmZpk8FKDZCx6IpTWdYy7J9GCw6iro7dvBxOpZCLvcrKUag13GrEkX
s1NaJTMSsmLnNPf0LnRwRfG02otNcxZW8tRXLVmznu2heDGwj1/EGfv8K+w09dd3
U1x7MoE11RingjjK4LvB5b8D8JFeXLtrtSCqshnHuFCPa35rJ7bIq2Y0xfvco6Ae
5+slUGSz1GsdO6RFWJLh8XiraAGp0iJbuVVMvJ07efalNqbWIaM5BDRCZqHJ/M2N
1wkBbV5odaYPKY8K9TywRXhQDYQWXhQSCllQ2ZGVhFZ839v3fhKEYyCT+QRioR5b
9sDFem5ZFBZbjvxHfWYXcVey5+Q84P9hPpXMveYsY6Vz6lWMkrkrk7PgbG6q/yXm
WpwKiZZKE0a+BFIMM6iprdzKGFeX6BwMFLSvyBMmJzeypLT04k0CmCqgtMZmRW5l
SMZuDauzMzAkXPvaXh6ER8gITEjBvx73ruzq2ZaTJ/U87znxySIqTnm0Rqkg9Q36
T1qqq80Gva9CBcR9NxnjsJEWO2pkLu0yqhQOAdYFrEkz0bOEXPl7ldmUyBnyBQqY
6iyA/vqO41bHXCUFmfcUqvRxvTMW5uHEuV5lbmKbwOfmx5YPIcuy0qHkW7qOcWQ0
R8vx+pRDsSVPMsxrfoS08W3WhmJ+Wdxecgi5G+PitCtWSUu+PrWxVbZwNj2CvkrL
j2woUcivZhGNn7qeF39X05E979NQs1X5L/qoGTVeyur0JdCeYXEk22ESd9IEEWyO
3g8u5uu8S+sq58akxJGiO/8+auwmiWPFE0qKD/SFLNGU472N8Y8dOSR7qii9TTNx
cPhEleBC9+HLVhqsoB629pS+GOIHbYdCxQPc5gDA5HFQ4rPRU6vAzsRqWJW9oYmF
Kem1PwS4MetHCQn0eBt3jzSPiG/geI3AkId7PMEOWc8Z8AF5DkHUx2XoDuEjd4Ee
CULWXsS147FNZj79TXqF8fTvwP/jM80cny+3mtiJ80UcAudPgX9GA877TL/Oiv/n
jQ2oweTkKJgTUD4Ua9CTcWjUBy6SotLEqbTO5RqzM3pKg+RHdgMZmZAvmYXA4bG5
SK/VWqxD+RLJlLzravh0vTHKF2n/l4kuP9DDkNX2fsHPvg3Cr1jAJBVyfBp49Zo7
`pragma protect end_protected
