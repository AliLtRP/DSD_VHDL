// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:33:03 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
bbmhERa5j2zAQtCBbWL9V9GomBaqnmPIAjxYaxQnxCu5XMDaROVu7Xfo0MLXQ5al
87vplAzdTcY+SQBv9O/k68C6/XF/NqmnfeVulweA5K1wew0ZMg1HQ5YbifW68yv6
+AOOpGYtKwYk2cE0caJVAyMRmRB6AvrCPRrc80XHmMk=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 6016)
Q2v90iT4eWs5tUAyvDIuhRSbly6obESnRaMyaxt6GcgNdNSbhsv/PbTUXLPwKpZb
nxnurJiMsLz/W9ck+rzpvFH4q5QCTSEyS3Du8MRDyj+fi3IkGVI8OiOaMx9W8Ix/
2JpU0j7LL4vWe70noUbMhNOVXLYEaIZA/KGloeUexTkHlQ3W+M3N1xYcta/cX647
kIxafKaC1MF71SlQTRdU0SJJB23bmejpqFY32d/DznOEGay5mnoxRPZgkRsEpdfN
fvEDMAQ2rfLfalBUFhJNVLeSsjspdpBMvgY34Co5wJx/Nnfw3PBmEgqBIjC7wEyR
da/R3fCz7sthX02FMLmP5BQig5ZWSXnP+QXtSJ09fy/IOHZO4jNG43DuWNfKvwiH
IG9EGU16PN6Fc3ejmX8ZlwBzkagux0faz0dZ7CJW5lW5E700uCA4dqbjevhmyeBb
wtBH+J0yARee/SvyYPOdlSiN/4NH5/uZz8h8V1OCT0AM7bI9SS+v0E9QqArmNK6W
QD+x1XTdJXE9sZhMjoP/pyIt6o+X0yjPtq4rIOu7TpKb1bj5KKxazsqSfu06f3F9
Yx7pShXH5vAmTpboTEAOwBktOQ+ePN+WT+VVEKbiHUAal9SYxKYY1MdkOALfRR1s
r7KAGwIT84m8g3AwJO8+3uR/Xz1c53BjipzBuk5+UrHcMVVIj2FNvhHMGlKa7Hfv
UCCrS9ES0Pr047w+NV9/MXdA3SEAzlRdOE9cflNtR0BM8dlKcT548KrefY6rQeYi
Abgyny2SiaobWoAgNiwl/nTi2TKd8suGy7YiIe7RCs80r9ezEaJn7g0IteBekfja
xG//CTl4IEXCZKUeGsdaxq3bCp2OcKAPnzEJV6w3ZiZGRgTaE35/ny+FLuW7HBAx
eCTymNZ2oWfPtKq+xmgg2eSDbnXa/uJVZmLQGYXU+XREDcPmB7xqbTlYP2W3wrTK
dnkb3pKQKPqS/Nl3oTVIDdNxK2PNkbryo8vuoIkJSxqO8vVWXRDVjMMGaemxbC+7
Qp7YayVPqQoVhcNIsibrUQbgZ1rBEpDc+oPWWEeS3AmvgD3lKLDqObli94TS5/sh
5u0hL/XFrIbg8W7MOgZ+IiZ1oOMrKvK5IAUeggXCQrZquinaDHnfpKIpORRKgJDo
VlK7eYBuT25LVSe6J0SuZ4mgH1pez1PNdgwx/VXRzO9UA19eGhfQQBO44BpWM04J
pfeOEA15OWeNv3+h/xX7oFhNV90n34ZPof1e39IwU3r27KYwSUm1HRR/XBbP9quO
2BBYeMRsLSFw8fCR0pZW1GGwgY12KAMoMvD9rtSJnas3AUuyTqR/njhkMPddVwma
nIb3mQLwyWw7jpY0AYvY5ZIYXnND3XKSPq0oytWtNFlauMRsn3+JkA5ngNNzC6b4
cHa+MeVNMJSOYTzhGFbuCL++1SOhPrpJu80OpO7mXBu7dNoiJrDyDPp6IyZnqhsZ
mpWqPTvKIphImFBSYxixEwbCmBFyUVoxsOp+5d5MeWyKIIRt2ZVd6h2vr92rUPxU
B5oWbwv4UcvgyHabOb6DRJQ8QX5oV/lZZo5EMlZwwc5WLsKBNbzzthyhwqnbrmT0
kFxbTNC7ksEb/HYoM0hgeGpSbuwJYdaWgFKb55YymwxcfSQvJT6gOnJgh4nHvHH+
GgeOJrVZu94jgfY1ZqfS93wMMnymGQHQekhRZeEEc6b1zq8Q4wVUUNDfPnwUIzNK
2TA/BpmExEo+zHQgH+FtP4CP7N24bG0EDUsU7iDbWCScCwM4eO37Viem+fuXCJTn
fZaN1/r+K89cBSjiE9Szu9iQxke8Xn0s/XpiBpL0dyNkJxlWLz/TZYp4IdrV0DxK
DRz/Et44M1Ha0fnwyM8eJ8KRyc2p08or8davw0B2L96Nguaz5GMHymGGouTJBqms
5wyvyoSOlXV9UmfieU5jfMePtQjroNZXw3vjJ5W/BIyaVjWfuidL2m17/Z4u1Vf5
jtdSBrAawsA1ZoQSOdECHiY90afRG3eKwTGyTUPeLlmD9o33gUfEUbRaC3XaTG77
YnJLKHLZ0FY9neTwvNzlNB7FNoO/lkzA0N5VvY5OYyTRjv0uyxQ/8w02AJpW+An0
xlc/gP404J3SGfRozimzduybHp5nMQR4map3utrOUOkX8fstRBBI/plahdGjLr2h
yUqS8rdUJXFX3hLHiL7q/7+ghyRfcS+QzosQAd+NSRbwJjqSm+L/r4a+XMlSArVI
TCRQlJpo6Ym3uUAh7KWNDTTLjfMnQRgg0GWx0JGrZer0IrkL10rXk0rrebxNLrQ6
eCo9pESmbn9rt/JRxPaifD8NtXWkOvHKkDbrJBCYNvT59kfbwi3m9WAqKQr08KTO
IwkGcL2jQU+63mltY+DWtAyDyYukwxf5N1yfrUtKt45BUFFnnNRdOrBSOXr2Vj3c
lcZsqcHcyV5tFuJxNooXdI/T3qqUqzXCoBZk7PFZWigbq0TnNXAcS5FTppNAoxEV
77QFqgGeZ5VZalpw0wH67HG5CKYtqupAc9Yg9i7xdm1sMwjfR2pRlz+noLWU+sCV
mNFgasaOo5FDp/E54wABDiJAMPF4u+Ac8tfFf2FzYYdlx/18991Q6B6/fThZ1wNs
QNNhFCXsj2ZVFPAsfNeX9d/q+Uy4dWtGuP61EyXM849/rYX1UkniMPesfF5Qtyok
k87SIZX2GHp1XPUQ5Ea2PkqwhS6GdHzVtLSQGzzBDq8o2sXcIBZSSzwel+Fc4heI
SjtzJPRdkXs8zKkuOKV1MSN2q/tUb5/JXFiAibFsTxdSQxMC7XDbp7E1K3+CRViS
W9HveovfITaLx9qVebg/j4rJnNTr8r/6/lJKrHRkciGyDkJemEGtr5HMf7NPb59d
Qhme2BZaZNeYBQrFbLzrYraemTUlNKO5t0aPDk5SVpwyqI1muVRkAK4m4CxPQvud
uT9E+Nc08pq0KTHTPLErGrdO3zzfc7b6AjEVd6uvtlg3S6AVxDQIGoXqtvbQBLbJ
sdqLljDSsveMTjbTRtzYvBSD+kqgV7NsBb7jnIZs2U1vqbEEpAo7A0UjSucWKBsV
E/mMpondXH6tJuwRQMc8hMGksyxT3Mkq83uC0m2pOGb0/UlPaeHTrzFbIwhjQOOX
aU9gmLfqRDW1GN+wmavVC3czMr5PuvICajrdRLfVYsgvOYfUdcHeD3evZLmd4CAm
AJRPzSBNvb39xZI5Ah2Xc8RPo/I9Pj6QrIGe6BsDuGO4jzWn1pkmTyRLUpjm20Vw
vZ5jYVmCbH4r44s+mgAcbGDm095Q5QANc1RcCjVwgYWU/zXy0y9baozoz94zkFip
1sboWK2HzBsMXvoFDES4TeNUV+kd/c4L5k0bsev9L/OghZQkYRci/2OvvRXBWUTs
+nAVYMF6YhXRmbcrpD3dtLBVX2ZDgQesPjkX7zAPiNonEUIZwNHDSIUYUj4mEt76
j1xG31cEId/2POu26s/jN4VAuOz80Qk+jxYVUv7Y+sJ674TTa0EHcPYLhe948qG5
EVBWvM6Lcc57fdWgpfbC8hK0sqwfj3EbSjx1MI9vYwyJQPGEluCjp8h9glnzMbO0
EArf3LIGZhFRYuvOdUe2w8mPlmFvkkPAIN1kULcUYu/uNXuiMfhkmH+koqWNm8mq
fPVIlugMi1kJ8gMTBaEDXsEgXZ8nCv1aZ6BIdioCFXqQyWR5Uaf/KYADw05sig1A
gcgtLPnltmHRpPXG3uaABTOGYQxawabeXsUHEiS3MDfBoKSJ3hLyzofnf45/mJAh
e+hjj2Zg0iezZyC+FaWit+ErrP27Nor3O4RB0al+tnhpIsBMG/74ntVdGZUkCfsZ
dOA+kKhkDW9t7KY/SA79JmqPky2E7B86jhRVu4ssW2utQCIGudn6VTrVc/WKm5WY
a8jmGo0+ZOPdJtC/iPL2qjSb9EOyVJbX2x5XNCxaDaK6nKuKHGReI0EL3qSwNv7C
CxxV0QZbsob8c/S38Uz0a6QERfk9xjvfscvHNpIxvKtTGvZisrhByZtLEYpBfPkA
FKdaSsdNKYcoOOLJfxERblBXRkG2I85zFmPYN3Y5wPThxrfFh64ZpZk0tLeRubAY
ViJMgab4OVG0WAPM554y2sk0yfORrTZ8tOAzA/f08N8xDL7mFW4PIu3K4YqnoiEa
jf/ILCmCRfkHKXHX1L9evcVK/qlfaf4Q4b97x3z1rygaQVi9Kx/v7mTuGnCcSv6S
MJ85vnWr7HJ9tH+wx7PxIT7XZUGMBTImHcqEI/D6uEBEuWbBipspvnbotmLNAOtI
3uGsuXq3hbeB8Qan0sdWpXdcrG6tNcUD6MXEj/YRlDUmb+vZfVJWepMTMNpXNfqd
jqsoL5XotxMBjD1lUu5CTZJ6uCvstUc+B3iiM9/7apoXc/az2M9MFsEVuYma208W
6zyQXziBFkxPk8NHzVoPKvQwZW0PNLQenJHbLr418LwrITvm19evp7Rg6PFySCvE
9luiKWgd5eARbnywXQa0ajiGr5TqK034OYfFhbdqVAefnDWvim715cWucUAyrE9c
3Ne+v0fmSxz17bl+/GZ6XsOPny6DhVMycihHV69ChnRfiWbljRyZPbjlhbbgnvGW
AG20YIazOjKB6rPWcNHaVQ7WqjQg7oerLTBXI7mDiEzjYEEBCB0U68OQQPyo7SK3
0o2oJHKuWX7X+txH+cK7qfMt/7MImXYl5C9om5fK/CCNUqv+VuWC3PBHKfNqy7Sq
N+PkezaU7+wc0QfkSnK/NZXo1DvdzC0PUtHpfY4iiGUgShtKqlsmn+MuEPjsNarr
iwHC3e3E+C0apL++sJqm95ja/wsHXy/hp5xNVpeo+LfBTgra4LsIrh2I9IyEVxZV
QslZ3qrEfK12gGk1mW3Oz9m9ntDM3Q/o2lLSuMrdLiT4XqdxG0zVXX48TBOA77cy
Ly72xWY1H0SdWQlzzk6RJ4JOt7O7nqFsu8FUreey7F7AwXbWX6R77lwFFekwc3Un
18tA8bVNxaKMCLKtCp0ZoQHKOrdI+ZX1YAGD9ir5bEKjuN98zRCOFbVq0zggxt7W
njXFcoCBT6fFW1lfaUW/2NPi/CVwBUfvl6rwqFyNXQNiqwhI9XrCVcHDT+C6WW1L
H46gtgnnvDaQ3BAbt46IXdQxwDN4NB6sHBaATrIZejwPg5Jb8TiUZfBk/+OSKbGG
Smn/4q+d/4XY+XTO+ZrhIpRe4WhyaOWTSHn1vcnkrz6bobQPWvSF+j1VML7+Hfxq
5jQ9ggYMpPNkwQ/OzaUIiORnYwv9trX4GHtE4xHOAT7YFcEqtzWUzyyopkHfzy7D
ctx96nvieF5dhhIE2X8qtgyyNX7vdWYju6ptbweJDfgpB4SSNkQvuBFwfMI3gyyD
JPt7Ny/vGwPFjmKI7Lx+wo2S0Z3cBkcaAgZDjMP8fmOOMTofYO90hNG148DVq3yr
fOr3kOmZsFlODA/sPdrPWbdQhTIaIp3awz2CzII7kx+G1GS/7MBW/8ZH5szkUh1W
xe/JdZnVNYIF3TjFMFsKLSctE4msbcqPlqEX+jto6Ch3KRLpJhs2OzL6r4sm5sWx
Q1kXOTiBg5sKgXyDjUDuAd2Ag1M6gTOe7nLh0SJLeSQqjxFR6Uq86q+0uV9uu0Db
0YjHjqrFM4GVfkkODpE8RuWftmcbhzl/IvQisvvzwOTlhHyr+hZEBo/fbAQDw2i3
QS1PPla0Ff50eEScolk/lrA+sABqSgUvqO0nVi0J9mYOGXoAubB+GgoevEqxujxZ
U268ug98fRzY1Q1T2VcJ3rg6Dn2VnZmfFBCJkQXFhHMkUhoDFsF2y+8FHIcwkVFI
rVpApRWSXIui8YFSPbF9zk8So8sjrUpBcvEDzg730Z3k4stMCdnO+haMfJHekmwY
WTI+0jt55w7Eg2tyraa2cfsYonNaZ5N1VBuAIPKmRV+GMUso1OtsOoPCQcd9PPNG
VTC4e+4GcfJ44c+uNIpIIZeLrhNmw4t5rskzgMjU7qjEiiNH5DcD1msToUv2dxJA
D9jvQ4W7guP/9J3vaICWek5Wjrsuyt0/o5sWQlvBvHS3iGK/SyiuopwuvbMkEHPg
aQRUX8UNgcOoteDjR5fCi8WF+2YR3+49yBA4XbOGyiuLHTq5vlA7h6vf3rHYZHxf
PJVDEvO6QqVKKJi/yl3g0Iy6v3vcpH/Qg/AVda3VipYvPF9QEagO2KxvouuhnsAa
4h+Y+Wg3v6aNrsJKcWYxOpnV/o1bSz4df7Cx/m8/+NBNiuAvbCs+77g6mtt5qKBF
68QfgtxNOOVA+0ag+FscdbfY6enjmtCeO530NXUxdS2zAb4xhytkW5qdTJKIb1Hk
Vf46stmQlI8fwR9GOZumGILdxx+XpGhOl/6bUMTJZSyvpDV2+EmuaMifR823RPOV
LztZTPzzKRXkF/NNP+04XWB7eH3HW3Njgtc07weInL1EOyYXRi8rE2E59sKtr12B
7KAu5DysfsXAShA6Q9YK+DvWq6UX7OvJby0xIsiTtT9WrZXoSmxx19xCZzZrGOPd
USfSCoSUM3YBxu2ZNJbb7BlYdWXDwGiX/lQ+7ZtnW/iRPQ6GSSVtBz0l75+ptU0w
tpH5IVAiEaq0BfpmZ2vdGOqy8mG/H0s3hU8TcJ19TJvRc8FZHRAcne0DIk8tZ2CS
VrWTDlOj8BL4a4p6Dam1OCK9ZkAB85NAVeS5SPcLE9fm/Kgc4e9nXsCk95Yb1o3a
syk3IIR/Z0H+3zR12dcg9+uQNsUm2BzZiKfvG4zRD23pM1ne548Mpsj0PL3Qlt1/
K9BsGpNw4tCmFEuzPWzFOlVQIVm8wT5QJtf/Bimrvj8VhBThYXzJOb48rzZoMhus
+VuKxPOCHvpdj+x0+LYMy8IQhgAmIzAJBpS1impuvafEMb+gCQ88ZPzVI1MSoMr8
fLC8kSLm2h8nVyT0A0qbO6kdke5oBz57aflYxEnskIyulKwd1sdmpkBa8g9nkeVB
Tr9rR3cxcBTkxVEks3PMI5AjQ7xcFoO7YYjXz8GQBsJzT8jNS3gsSDv9aHm5rR1N
DpNc6Oa75dlOToyUeNCgPenF49S2V+wruSXFcJd3ZVcUmkIOa4VLTZQ19uWuBBpX
fMpXUNYTmyb4SmWG8epbKe3XtBg1D7T2DW2GQF+GjwzRRHB5zF10zohtrQB1zbFZ
8g0xpsGwQXieUuXA+M9a9Qk6XdZOBNdqXjBqFjIVydftUq+iP02kIOqi/OLGdUdc
NHY76HN5w2ZS+jXSBckS7CDQcRC7CGLYf1xn6907JsYmWAzRF0G4+b4xkcvyYF2X
t19svqS4TaTnGp4VIo29UjsDqZPoAm7wlMsZBhV4cIReSbOmwmGuMgm+tkb7BpJ5
Qv9URUKqa4kegPOIfvQhJ0Q+zFVOScM82rgLEOgoJkBZJUHwwwcUNA+JZTUKCG0q
PmKtUTy7524tryjbcENscqwQBP/q//M1fjFoqIFaFOwtkAUDrAaDw0uThQ8LQKQA
/B8mM/wKRuGvK+vbHqG3j2Rb0CybH7KDk3ElEEA/uwhCX3i8IGx9qr90NOblvU5k
c/fC6zRwHa3jpDgfiux0oUjQgF9XVqa42DfFYDmwZU4eGdKv94owyQe5b5TSuJNo
HvYGWQ6aHdvSiuJXA4x8Gz1UnKbaf2tDUN/yNlQ0aKqUMVwCLIkkO5PBEhJir7k5
Mky5ok6xMK5v41Es/pg61ZZZgnftQ7MZaI6JsQheQSPia5rD9HTIiuDzgQcYZoIn
PK0eg3t7R/VmneZccM84N/wAbW5LMZpkMfGzrg2h6Bv12dNEKFfCuxYMzgwt51+6
zX5cgDp+tyPiE8XA3ZHkOM6NyJL1ePChNd/lxNC7QJJx8FjEkpT6hIFv5zE7v6Kq
wIPaak4vlJJi3e5PH2kz/mclyJgRnJPhPOCPd2J447BjCTl6zbxVQ27aRS7r6Jpw
iMTPEAA3vsQH/rfCiHsoOCa9mzGPrKFF4ePTUHpkw7QpkdPNyZ4CMOJcBsVQNIq0
uoGdeckZe7u5FeEi+0GykQ==
`pragma protect end_protected
