// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:28 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
I6AE1XRhRdIFfiXq8ZhbK/1tXZL9ECCwM2LY+8YaLrKt8JMajzsmCIt1oCThhb8a
ogAfl+ZQKe/+bqB8mLByuCs8R1VVBn2p+j1s44K/zDuQpxa8tVN4Rn7d1c4FhNNC
r1s7tTw5/C1E6OUYw8wANPfBXhGNuOFnYu/vNkXyoTQ=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5712)
GllMt+2SJQmOTGYxm1gJKyRSSu9szHpZUxhhsVhXSw1D+J7QSfCLfYbZQxEoDcH2
kzAq0J5OAFgY03zt8zAWSKl3e20OwbB+S3hY8rFr8bWx3r7qlCZBQHTrHJr4BGkP
lYCH7xYoc5MdFkU89qEA7VNOeXDlIZ71ZTOWRKfvU1q1Gqfr/mWhVeslC6Ld3PTg
stGispNnAb4/l/Ci8QjqerAKhdEZqPc1mc/HW7R8murlKLOBpJKP1XeI5RXgZJ5T
1zkYxv3XtHJDgPyiNI9p2nWwHIsQYemZUwehU5QqH/AOt8Qj7/QIouieFe2D0M3c
uK0QyGfGgus8ECd3RhGS8/IhYqHjKTiuElUxD89jdys5XvW5xvdKaAqF3jNjPrmk
LXtaxpzFs+mPABoj9cesiv/Pc/3gVwger3fq1fjdtY+bm46vXsNPc3YRzuuI4UnP
x2fZlQcBZ6bLLGX1R4bKdxu1vbyjjxmwBbmVI+cpCJeCKNQ7W8C+2j5mTlgq6Bji
mGwKta+ysjwisTehWpNSGyd+3y4/gtvws11/AXTHfZytUER9NlhF8CuVammN7B9d
Y9G9CsQceNP6N20+Zq0qtnXTju8DujWULqhhfVatpMZFW2jcqptnGMC7nBQcT0VC
Teo9qYsx9Bn5Jd8GhUa0MlCqci6G4cP+wLy3TSzGm9DwM/SXUeXkhLhl3s5Tfnjw
qqatD7GlPXOmHZ6wnGjJ/WHzO+fUm/25Wj6LNOGEZg0B7FxLbkVefLTboh4Nf6mV
3A9U45iolKrQcUEFFhuaurCwXuGn8Ice8htlu5IpVXBGzYHLOhDmc45tBzIdXR7y
Evx9ltbZzfaTuEvz/O7llS64E3B/5jHhfVQWNB41Ub4x5H10f/bFCB0L4UWRu1D3
l08hVKt0iZrQvl2IgFmI9eUEAv+L0cKM4DZshDdtB/tf7yj5VmFtWQ02mc+ixsDB
XhZl4YwOJKruN7AsVpATOOplLzrYvkihseTY4q7Ls69ncr+wgOSdH+UvWYxFWfOk
znbX0uzDScY43IDUyIL2AroFCmuOoZkmMZR0YYFc+EdaJOWGtxyl3VuEfzQVGgbY
6xzCy9BRv32Gv8IiYJQrTZsfPy59oSSc8DX28crHsMhxKyR7MmREfVxeKtNDJk+E
idOe29xIqS5KT6+IhmRPpr8gnsp3mDshUViKpxzXAmsquRDFsOcjm6TuHSIs258b
0t6o6dFEPj1Tz7s4Ts2hlxEx038QeMPKK6o+eZmXeGxBYzPGK4VRa6yTx18Bq+2L
oSdseZmMnvyQj8idA1u8HuZomSPf7U/ruo6DLFDj7rMIRQOZi1+VQjMRFpfMuzs3
fW8TcrpSl8Xy/pr1SbgJ6B5zV322T57S0DwjUADC75TWVCWXrSTOO05YMwegrBix
uf5FFjBz27blDUtEK+Ny80R8ANr0mTy7YCVdgiNTgL/V4ACAaKs/a2rHuBXkHend
CYLRuFCQgmzvXE1U1y5vkTe4I4w25y66IuTMpVAprVSRifVadzUSdEOpjxbor6Ua
8IFS6IFNer+R9Ekp1SrKPATUuxeLjFObC02X7YxACwS6DdReTvYr8iAanT3+s/Ky
6wWirN8W4exX/zIrXmwp6g7saC8Z4gzX318hUWcctjwvo8JBvAHKcPhcxuRjq65Z
dHrDgsMzN9yIaYyQIiT4xoZbMmCEzw+4UN2bJ9DoIThZmuf/svFsUZBw0IlDd8g+
NH8o5XW/ajY6lCTbAx5SJacuSFj1dOaSUmCbFWigQR8xQBeGK+pnBiIJL+WC8VXO
ZS/Vl/0q8geRG0zJz0YGW15ODt7l1K5DD3KNEPh0VHnyEvp0x8yAH0TMeXLgn/tv
nHckYMW/uPCClMx3j6JDP2b4MR4bANl8MASkhhDDy9c1czr988Il6+rtq1zBoW1S
U7VH3UfgkoVmeAYCYVecCChtQ1HAtACGkz7R6f6wJcWyLQUnyREfE2aOmvdFSJUd
fnzv9riLsniuMLq1vtP891O+b3p4Juhar2Un/Qy+fabK6MDSgSTo0ENJwNEhGoEo
STFEt8UMyKQQkkYDNPcOQCDWWgeXfcvwNXZUljga7ZxEoo2d4juehQkFVDTFAI6h
oJpz2hooiDt8v2BFXVMXNcNVHuEGvXuEAqc8c3AD8LiCU0Ya8Zdt0sSBmiJAXBb9
jWufkLNkWzJWlJWQaToYVSFJ/lDhWbpeq7kyEVSyenb4EyukliJq7savlygBa4Hq
B3Ev15BBW9kJwDMWME5iNKCUCE6TxAtEOjCFMUDcprhrKvUynvKJmVXr+rPfpa0e
gOmKqxSB5UbnFcPnQOfWXqNq49a0D2wfUcUssrXOqLHMq7TsRAcFfCzrPHaCYM3T
IZgXJil6tvgOCZy82ADrzT7f1qKZushM6xWUPwngIn1IO1XqX452I3TL7ZgNET/g
IcP3k2cwFZWvVfojS1xuJx/AEajthMlTENC4rRNm1U7Hvo1XFYUhz/y5Zmc/AUEl
pYnE5SVtITYJV/iegDenwXd28lCcxtYk45nILRKATNrUoGaVvw90+4JuF+H7s9CI
WKlsZREsZupSeJhu6yR3sku1pCdWfmnBUJxYsjh3mcqIboh6zZU6RQfrYmymrwpa
7mIVz/PTa5hSjIDZZsh5dgWz8sVyGY8Vncaj1o1e63euofinCu8RTBZOX2qtwJWz
w3xkeEhHphtBgCw5iq+fr/A5C9kivZ/06gHzG1Ag2DbViKR4n3ZEXP2Y0TYSHrJp
uBBEM4kURvqUotCfEVcMUMBSurA/k3bkdQi6DeXTElegzYDfzDHamDVDsf7VyILI
yYfMFm8s4UhF3IJJnC1T8qhX18FXbByFgZWccMxfi+CB287c+9cX5upR9TLdpyX9
nJsGVGfJkWoZ2TSVbcvypkB3PPA1hwJpTfJYc7LJlbeBmebKv5yRgkW3YI3QN5oQ
N+2nil0mufTTMjiCqkqFrenQgse1FsBNUeRYTFQ8dTwvsFkAg02jn3f6IV/rXMGl
Yv8OwiBLk9EJ9Kr1DWStI+q9aFhqPenrUlN5YX0Yprqji2B8+FSc8ym2l/JEP1li
GpqR2lTWb1pY4tFz2/N9zGIEPTywTbeAWcJaFQT0H2WDqa3scaDlYHDtXb8m5pYF
0ZrcEoyFkNyC8Z8R+tbvqoNHB3FkvVWEbCbQHfo2xrA+xszB6hGnybhyWZFquN/+
L7meUOffhDBG+fzMOJgw9MOoxqRezXwhE1EFxqKRnpT16Fz85N4v7IVexcm6wMPT
cA+SCdIKt1BZuZa2Eks5GpHEQDg+LQ9hEQAr9jNPd3g2I9EWFL98BDrevIQ9Pl2a
GrPnB7gpfJzyrZ74U7ImN4M3qyyw38z8hjLwezH/sU8NwVbyZ6QkCuiqk7EwqHdK
jOVrYkJlLFCfc8cBXot/zH/mNkBchlPtJHf9Ee7KvcLu+dLsm9e+7xGimVFcB+1s
pMejMNl0DW6WPLhdlqpw7KuDnooiZs5TvY2+FDKICDJgPCH1UeHLpqSb4Ys/syKX
gKrkX1k0Fb4r3ziKAOonzarbO7PT5DAayBsX4aSWHvBe7HzKXNs5tB1d2Ggkz8tS
lLCz1refEjzFNhz07rBqOIb95c06k8obUY/Z7LE/TEzzUX97IHCl5HyQujOGnHbH
cjdJ8ILtTkWjpWMGnqc7F54NjWo01rfWG9Lt3+hOT1GBb9IHacRQ81uP72E3P/8K
XFg3uPf4H6Emg3lsWv88OiA0Dn3JZSa5T7ypYlxm6RfxFOXZIPWDyqYjkZazHPlX
m8wDpFUCMgOmQZAmXdJKzc3si3qjMpAi0jMgKLF7OWWgCP9aFIHestYgXrC26YUd
4FhyLIAdiWgvUEPoRXX24x4CXeRfemfUqBY4xJvjtxa7sW7JmxPl8JjlDjpE8v9S
RvQzdZsrs6Rxy0wtDTFDcux/lGO/oWKXfzp8IxcBEjrHUp/YOqP/NICt0e7HU0y8
iXuMAE/I+zYEItfUOXgcbAxVxLgADDWWm6dZex70IRXXpqSGbc54s2z/7cAOTmE2
ONplExg9xbm+GAoVYXCnYEfO/dcix179sWXloHfk78KXeYqLcNBhZD++s2EzUA6e
drPolEhxuNVlRFFfLPaXLop0XhFXEXiz3xpw8CXsFw63kP7b9bPwBRXgCX0n4L98
J0F9CBLupyjCFqu+8eS/vP9jnhKCGSL18SETaJaP1HrvHeL7IfhCHOpyaks/lVpx
Vl+9fTusDzPrRrxw8H16Z6So06Yp0Nuun40GaEBuIYiM0oQuv5bCBnsk1tZ8ws9G
HUWRaHLRoP3CgGfVJdBIImX3tyoD6pisZoKKAQShzRiW+ilwidpw7liqREIuJTSR
jRQhLLpLsKpuvDUBrhEP6UR7TlmqpT3UNM4rJly2pV3N+sauH2J9Z62whs4xXgVV
DvtNJXhfv69g157QCbMqERxfp/8DKx303UuNg7EWcf5kLk7y1F63hFY9sKzr3+09
0pKpjMrJ4U8RPT35P7a0henElu1XsRLYXTWYjTX2tiNd+F97i38GDMZioGILKTuY
d/u2ADNVVBKBD63qe8kFR71WkViGiiz7Ytg6HEeIXHFp1VXzCpJeOQsjmgrgpdSk
oCAc7B8hiKKVZR6MEKnOpgcCClKW6XAZYSjeLMuo6IJb2/n4pVDP/NoPNxQbZVxY
w1FllNJ8kOUfuu2BfGzl/FR5Cce8PziUgtn2XzgRNmgZ7V793duxmWRaQooVzY/H
iH649nIvp/zH+NrdNPl8WDTKWGYvlCVJwmH4aVVPuagNCzmElmGTkmz+f0r2Iaa3
TBsMb+Dp8pEp/8lUqMRQm9iV/pNuUlq2YYbEJv9SWvyf8BSRhi1McKSEbtkLNKjX
QKZMcTX29R4xwB/JTAex5jDBqKygilBJuPilAtvxiVADmFavqzVS0DCh0i+bleDB
MWf/IGyxJUHEfdQ/NgLdBP/rEVfcleBwXXtLxO/lCP7pPUKFWWGpJxlzLIfoR2+6
F6WmSUaBFCPnKD2mrX/hKsJQgCK1nU4+D/06wZ49sZo24/8Sn2sUy77QwwyAGyW+
LT3pJHoygNAwlK62hws+kD5g39YCeGReiouAEC1HxC0aPNtiTX5ebr+L4Zh2k1f3
KD7eKh0L800Iiy3HwG1JivF8AWsLsBxSdHUg6ra+CPJH42KsAcJ9fWCnBiO4Z6jG
R/MFhL8vRS7hnePHJ31XRnE9VkDDhiGs/EGD4zF6H8fZ0o+nKtZ2Vsv1sAubr1Nx
fMxFSTcJiF8iNrMjS9TA4y/F9EVmayw7o6j4W9CF2E24uqxSJ43+DOVVadchWYma
dvTWff3pDya0UfLFxQSnvQBXozeSupYIJq6h0hicsldkSzLx+b/pu40bLQpCDpr8
1/shQO9ioZcL5M2HZEkXVw1ZPM7JCvp8ig/LQtB8p6Zt4pWY1dM8VVyNwSMTYkfR
uBgygXgsL6XkFMaXe3RDtBf+7YvcBMhAvhrom7IipPXOLQWhp1i7w0Od5et3hKPe
MOgTSgxemB9Yf04OlMMIbxsSRhRW0TA1AE9tj6cqlUN6sHR4C5JgesbgMcZuznMa
kLH0Q6fwc8h+A8ynXI0hkCJFQcl67160eSufDGxkc5KC3Mr7on9aePvVL4QPsLtO
Wc83Alxxs6K9R8VSrZJb9F/mi17M4Ao6buJ2ibPyLto/Xf5QskztE5gSp7P+7X1p
7bUf45mwF2Dg0eQBGYDK7GHWoQPgqw9zMjTX1aKMs8UZqB2W4yBFFImH38OatQkj
60oBcZJBXfXA9NgAk/7QFfXp9EkSTdJxiQr5ZDtQwiuHeX4dSB0kBYUrKycpX1j5
9KkCgb3nQ9EwpvkhakuFRMIcyGQVEWXWua0APCKLba7XJXoUg6GVN83X9Jn/YBnx
FlOdC4Fl4Gw4JrJoYFty2HuBPvGZxx9JbO+BwHspG07rEvyichipspNa4XbhX+Bt
BOKN4f3Juf8hLZwwMndOIu3z/T4P9w9X948ZoJSHbYt+zA8ICbSdj5eOIkAQG5dz
hpekxCj1XRIb6t9+J8G8fio0KhYXrFZNlZvKeXYuEJ4w1PEs4NlHtmVV7KRfleq3
A3Dx/OEA8wJQzTyGB5W4fVbolHjiqDU0vSG3XV7OdxSW6piKie1fIWpHKCUW3jTW
1//FBEnr/yjDPZqH46BOPdcu9qtgsZJe0IULd+OC8m24WuVLtXkSgJsDqeigvzf3
1zJZvDpRy33eaXNHHC5dgL8MPIL6woEYz1ITs9BwqGakaHjOb5zysP2B1HtNwdmi
xqqWE3mLDxBOiKZ8lEz2j5lAERkpwvlpyiywzip3nCYkfyIk/Nm0LTLvW5EawLMl
6ynToygAVvtif6Je7Is8wwrBmB4SoqNPX4hOAbMc9GVHprQKjlvM/aRXlvLbgolg
TapfWSecxvXvT1oHIdcjf7TG/PCzW2WXns/JbOdkGMNOOhR/PPcUD7p9P+nkKqvr
/7r/bKCaEZfwl9smlxZ2dy95EMnW+Iszfcb2/tU66k7nhSxb2hm4KF1NrpgrB0zF
mRWap7oyqAA0wp14U/+Z1E75hEyEuWvAF4W1ivawuphQaBmNGqVBpN40alasaZPy
sMV3AyFjeSWQqp2uQJ8ZvzkqQ8uw850d1IkcPQfxqbRoevwhdEgQmVc/e5s01oiM
WwsHmP737zNSiMtvAMbMruU7FEWooncoNbaEf+b6/EwxmmEirEhE3tri9f5lunSh
pWOl5bxxRoThOGq49BA27+yrVsZopu2DxJkdc/kl2InoQuXjamwQz+buIVF20/Dv
ZHlLV2Rh6R6MXfFNDYieULxEwY/ZpqvIt9xc1jlTNhDX0x5wPlsaggxGDJn16PYr
tvkB0i5t/1O9ZYJg3hAgLwcCoukhGFvkCK9nTgO3rjcxPWYWsRauudcNgp5u0WiG
XBGe0WcuYd0HlK+J/R4tNKFWTWT2ooqW/QgYzFVAJ/Nzb12IjdPk5eFPRdkJZr+o
k4NraWt+7ceZW9uzjeKzN13dimgZ+bCT0GBN2aO0tnCBPQkXL62L+CPtFtFaStD7
MXDCsz4rDkX4NT1+Qeh1l1WH7X+gscv08E2nh+SP0baXah/ZSc2wlnX887SBIk5G
b7IQ2Bp1/q8t5Azr/scBB4P4ddqVMPk+Bl+QW8xDAHu4Vdkx7zMDkrbA7LWDqi1V
DbznR6X530Ghp+rFJpoN1vBg7cYqU5V2gXXPSAMh8zhYuDG+cpiv3N2Cng2q/y9D
yXnqlPmfWa3QSX7xrJvM47bHox2iCMoUPB4tzoHDyLxU8TvOUikX3roF91eLLN53
FAomVYFSQ4IhrTETPt9+xdUb/wwrUcT+dpzG0KZT+Id8p6UVDvoVY5a9oZica029
cPGSxcmuTqoNEuQ0sdyOjq1nZovSijeMPjo9IG5hwlYsXll2X1R26jpVEhhZzDvi
AAb4KxQEIUpzdNx5+QXcnfcALUGQKXUw1dnncjZaxQAuaWuYEFzLEH1dfHZcZ29i
q/xJPV5jI2DiKHkyYllZhSIgKXopKIOJocQ2r23XuD8DVMu+ZsTRyRZVdq5l/1OT
7mikSqTZpvdPlytl+/cx8ueQSzNT+bhJfwH5weFmTW0hsz8FR3gorxDCho8xNyGk
`pragma protect end_protected
