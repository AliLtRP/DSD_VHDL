// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:31:39 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
bjT2Dg658UQBRdEuDWsObCTq8msvqdbh2nWVtYNsEMW4gBzwiFkvVyQnXb0WZ1Xw
8uGPA+tU2dWIYxAq4AACdvG91FbcPC8qu9PPfNBAGlzTUCiod7u6+JKoDr7003QL
h5rfkzK8ki1mNC7i0Y1hX8IC08lv9Jb+x5sczF4WdOI=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 13072)
eQkotTiHL9QY035+flz35JRYWzx4PSaLy7FC881wQv6hQEH8Mp+iAwE5CrJiFUw/
HiDt6gw4P2XXfS7QAE0uGbpClm51nfjxY8zVK4T9bR2/jQ2FHxgC2La/EvW0y5RO
pUxC4VXqbnHU376CcOYJxSsWFHJokEixUlt8SbYrCsuNTeFy1wxmlLKQGivA5x1n
2cjWpFXYoBniRvnbcjROnc0iEE3xAmQSCBzleSVAMY74sPAPFXCFWSBSn0TtdZs+
NzP3/4/YyWlXn36q2gSR0UH4yB6/rkVYLm82OFc2hNiEyEePbrNSxSVReYpS98oS
S+FnvV2OANFrOE/WHiOY6rB++Jaa5lRSdPTf/qTOa+ncAN+KVtuvgjkmdQG9Uoun
pEtLn0g/CFxwBIpgECh4I81d+ZjQkn8OvxSnNxwghBPpmp1Y4HUEq410n67/Xd3T
hmCPH8Ou4Hi95w9yG4Y3BQOO6skHEdgChrEr7Dzki5CCCIDx94v9gXkgAPhum2qm
7tnBZ/J3k54jDkuJxL6y/ffKaQsLqYVKTz9mJVBMC6Ay9tBwwd3C2DwovdTUq2hB
xhq7LhICzrlsrT2E2BN8URYxe0sf80SL6JumcO7jrdjssYTpJIhJf6UcFouZCOot
5iPBjemt7zyXqkr23d0bs+7uhlnHMdE909HH2qpQhilj/zJHH9z/Pu+huctcDaFz
NcZ7m/Yw68J4xBYEF08JhlexGOVmSS3rSPnwvyo/iolhYvzukg6qiXZWdHUnBe4q
KPM7dH9cQqCD0onBHRyvQMSYip59DC3ESgjNReF1YYb4Mr4Loelund/wCJFeUq+D
TihbNfJx3UO80PyH4dDmswxnl//BS4XzG+9DBXkXeyRZBxSlTFftw7ggi/qCFHMn
xTxKq9CMHC+XVZK2qKKTyYcJnL0PXHqyHumGB7MLXglaf+SasMB4A9u5kbLecBXb
wZ96a8Pm9nyupX9/KN40tEVAPUGNNSFSkmhqdeL1BGPCN1bxo9jQl8ATyGmHO8aV
vzXUEVlkrGECdntbS3u2jfbTAAnuxEQS3zJaIxc6jBVledaolO/XL3aiscxzPRMA
J0Fx6W9ZI69V3DPjYg81tZoyj9282eYWR0eIkz1GOb8D/tZcCb28OXsl45ihOq5e
vfP99pszYAOL3FAgkRktrRwziWvzbfITub8w+eN+VIF/M0Q2Wu530vN3EIPzLaxQ
ejr/zaNjrzMCnZ9yGMDxKbfRgj9lica+rJnxG8us2AlKxqTGLjqHngr7zJR9rh1u
+gh0qzxJeuntkosKJMQl19l4CtBrk5F8BUKWE7x79Fe1pTQ08Sora5UaWLnoZGmG
TpgTluXBWzfetjUJJFTZXvFa0sWuqoDwjHNaWgs9p9RAOGqJEGwCVqgwuazJmNAz
eR7lTCytDFp1pYeRiIkmQ8uET9QkiqGGpYX/Ya5nl12xg4nOzcbhfjdsJ08zNepN
1z6Js1q0QZ1HfYKgqJwvV7YnsvKJulOBn7wDdgj7uUQEih1C7RMkNIfaO/8i8j0h
F1wmX8Kb04tKIEZigBdrRkTYgnIslwHzWw9octht9d6ozi5IHYHOG8q4QZr2OEBG
hTnQN2uTa2vxqDyf8AfR5sxuQoYcvO2sOHRNznUx+kWEbQmQdTex8h7s1jc9R7AX
wRwaEGsHFGLmRqrJHzJgwZebQqoApG+ujrfoolz1xOJT+HFkAG5EtJ7XvgsW5QGv
tnadzXbKamNYNtpyl/ry+LRr8BqzMX2WhHdvkP3wjf+vnZqfYQwfItyYhnxmqbwB
hGiq9gnB4ptlj+dOkXjY0PsN/tuzlWdD7bBxcIJNlC6FTueMA+CE/amVzfwAjcB7
gB17vZ6um0skWcu2VF530CHPaPsNz2IjefA2OONadkz+03dcjf/tPvmt7w1c3mmS
bQosrmBReEW28Z/jr+AY3RC7UC/3umF2DnVjgUqFBr9AgXvtiTvIGvm27u8MDG/J
ftGwt6a4HeJR8IuWjykKvokOMGu3YAb+ai5lfZnjG9B5xcegT+W5XOtfGZYJnI3V
2qZKTfvE6KO9qvkG49OKk0bMycBylvESbpouvU7cziFLuumlUonTm+Qo1tg3iVfO
f3o9rIBuOD/GzwAhROSiLzyI3GYUhdfBIkzVVcfo1l7kfBSLprjMJB2ABOCRZA/L
Hin35bFrXYWYHbO0Ie9+AKa+6TAQB56EOvJ+GiMwrD2rCin3Pw6oxBVFzrvLGTGd
QHA2NY607vI3EVv2rs8Xu1id5k69lv3B+6Glh/AW4bdW0378HypW7W9EdIAZEzEC
vAu1b5yJveqJ0Kyi3SHaVrAE5mYC6jMFNXO3aPzFr+yjAJDmZHXlcjLM+WY2+nsk
WrVKML209BDIdDphCVocyvn/0G29poyq01sX2bWwUiZiL0dolZdCiGzUdJRtylAi
jznLrI2lerPTsNPQJ/kYsULheQAKXfE+4tn8JM+Glwsh4PQsOSvXpjq2uB86beXB
UfPvr6LBLFjFGWRmdbPi5yzOVvavgzlNyahgYlSbkRUh5mNa1pOpPGfvyA339dyw
UmiMtDhNQuDJP4h2hQEgha8PxjROUe6UEILUvyntO9HeczULloEE97IqPJ+RDefg
VyDU4SDFdSg5PxY6LCjHt2oL8i8+Oxw0QTVSg6+2dHnpSlX1bcaBPhVcJMeUN4km
W5Dylyffn1nAlzxg14ZAHeSNKJMy3cwSl+KdNEZ/qRkkRLA+hOoLhDnsaahrRU/1
HjAodeX8H5lq0rbp2Z8wHfTxJJYm23v+VwJSiR/dtSk/yX3f6J/ukDXLWlEkvCtx
4r5gCnswvLI31rLPIJkJDbu2eF1UzA0BrD+E5KCwvpu2NNL4Z9PlhUZl9WSlxp3Z
9VMdES7vyQS1VrikK1mPVPVCCZuDJfrUGU2jaacTOro3Z7XFA/A/aJVwgbu2Bucu
eTJPwszFTBFaYVPxa1VXrxERPN30GbwIdO4JphxE86YlfIgNQNvteI0279DeVx6J
/VsDyCfXZWzl0rf54p7T2ZluE2VZrRjVQrWELbMefLC6ADAyo1YqMz4n0tEnNAaA
AfWqWYxfOTjFQWJOy9zqqEVl+kjzJlIlNlLBtp5xRUnE3oRq8R4F49IIvXf2ESXw
qGsjY/8G3SUhckIM81NMiO1sAFyO2CS/7LwvsZl4kG1Obrkjtg8lyYMuwYEewpR3
8bvqzMokHGGIM4LT9wQxTcLEjmqheymX96LSdukKxnb3vQXMrF0uTetpu2jP5O4n
MIgS/FURQisHkrl4tD0hypGFDEOIFxoZLKnjQO4BfNvNFIeLRhiWnaS1k6uP9bwj
/xymzkhrtNwUr98GEYpPZcluGp/uVGt7CU0VUXn3eI/apo29atIbXJrD6CFq3Jzs
TWzG17RBf2wADWZfLzgHLL2mKGdZgxxV2G6QobeuPbXCsUh8KpHiZT5IYy6LkPSC
nu/n/L3ImVMiyoxYHgsscKoPbjW4S376ejkT4KaRuRS+WQb6ALnO1VZtpY0oeL2B
kf0r65Tmc+Wq9Si2yaL2Vxgb8+6DVgga4qJcSaDJkUFxYg0WgvkiBl8shceddSuF
1kCOPvOdrhqDOaI+tUuLmeAdJw0nEnHgFA+SxTj0WgyTja3pHIzsn5YE6SCaaFGq
EIZpqd/+PriYroB3zcGQnkvQQ5Sau+aJsh5xgMXX420VsOZPwWCz+PSQHghDbQGt
zrGrqmHyG3KqOMHsTjvBfxMWegvdDLkvd3oOVZQ9XHZgEbybQcanR5a8Ngc733yY
a9Ixr4BDdvKe4pJADnv7batIzHwlkEAb74VxPaGIgwuhRDdREfeyj8Dzt91uJbN8
8/PhaUWmukaHAFUmRFsVNhC/qr9go4zPrDiWfMOqtYSVGv2vkYuB73mNzgP1ZVsi
YbG9e5ptRiTl/YUydgcOdvXoFR0x8B8+S3zKuOA4xQrkV24SvJOHNojaxrlQ20z/
UDfkk7Gk6oH6H57U+wX3+ujrvXLp+mKJ+O3sJVHWqJhRMAqVX1jNTX94HiFVjhYF
fgeft9UzpGF1vVvUrESsac/NssrBOFAjScjuccf171RqhPRh36bTFADqOLEch1Mj
oVcWZAsO8pP+/0XhvmgrHzbLzvFerQVmzdne1m2JK9oeKDrgHN21c2yQ3MYo4I6I
+/IiVSKTtKsl2VCBAiKIlbKyL9T2HLjnCSrD8/GdiywEKHgM970taY30pd3AIq+c
I+0xfGdtHrZ8JjIQ6ebgWtnfw+4mfJgLA8IxyCKsS0QfWr1GMpay0dlw/dIs0jRA
g56QSh906o1YvOW4SayJmdPlQnaZsAop45ZPX2Fxkhva9BCRiasTmFe0ZtDDstPL
5UJOl0cqdF/y6nPml+XF2QOI26MNaqWZYvGnbCVUfyK6XMUW1/raZQnLQBHk9WoS
9ih7u1O/j58ZiFZSXWJ4p+LYctg5AAglg2PAWLobEg/kDMar6pWPCtcp8O6WoIH2
ckxu9MY1Y83LJzA+r6U30ATLfYTXkbF0eUI/gKypDR8n/8C40zfwHX62HsynrwEX
VMmEBhBROXibkGczYNrD7DtFPWFghhfyKtU7nsyWCDe3JJ2VrR/OF0+UZk0hEHoB
WiqnLXp5Rab2MzPalNPBPFpyWKu/S4UycZoXlpDdqDAD5Xt3mpPlLXXaqdMHaYEh
nDgywDHO6pikF18YDFxjH5Sftwa/HOwIZWXXQuFA/rgclcP9jhx5mZ226+xyQTLW
7rtNGjcPuW+sz/E3P98U4LmNkkaCB/jr+K5eamTAgul1fVAh0dxtLF84pPdMoDXM
2hsfriSlBzsmL1B4j1MGB3MlcixskUPVxUEhoFRRjY9guvYu1PqVk62Ti/KRfL1u
7MbDCJLPBmhtd88L5et4mQ7BJi3tFSuL54pmU343ZoUSdXxJ6hnvJICWuiwADjO+
uisa0vCa07/vKZxbkmwQJI44OAs5gtQDEnDmitfCIuWJUnepJstE+ffOThsSZICT
zZ/ZE0qOAFtrWhi8VjJkIw7+VApyafyP3DBrj0g+rVMWmVMwgFzBUPDWfn+9jiGm
GPqnyQqBfplWwTB5UEFNNqhlf+vEVv4AECi4dHgnLQoPglt1XvdUt18qRL6ZW5Tw
rT+D6cqmFZfXCdbEF5TrCFBXT0llJtBTKqqDbYqPNOxqBqT6+CHeNHDy2rL6eR+C
QQS4TJ4+KUZPSBZUVB9+NrOhY4pybPBGd7hv8XJeBvLD6aLENvKMJQUMpZHLJYAJ
+veN+CnBdRJ4s5VRuJlSiflXwEvtHvLuz/bCSa7Jpk4lsKGDL74BqaqFMrnY84hu
389tdAoY5xQqrA+X8LsP+6wmy5PYMAOTDL8ev1OC6GLfh6YbeRgUfS0ZxngQ19n2
RQHTxeLg4feu8qZQ3ugXwZjEw95mmr54ooUg8HJ20lhh3CoUibikUCRt3RUx3wnx
pAaokTofymtrB4tZugxWuV4ARkWQIj7RoorK1/xN/m/pFBuR58oWlxF218cucgfe
wNniCWCXL3nN3SZFZDEK6PTMoAKCyQSnS/nW7iJvCoCgsMbI2XmwG1Ymle196lwh
A4v9aj/WzAsUMJi6lpfUb11HDtyLel+GaFUQJzhcoMEK+UfqZQQN/nELUsY6asXn
JoccjefYinSjBQxsimidOssZ9y5Tz8HlOShoLHNLYb2izQ+KAy/4b307SJiDzXdR
DomJVJInEGT+DabxmaxA+h6Cg2Bba3dr6oMksOuXJ0jRikjCMlgS/wLkeuRObpCM
JXyjRXlBs9z5VG2foFhX85LuExTsFGVJ6YV+T5FyYJd9h1ccpGt7TOemvtdEm8ce
l5DsV7IRPMHZI4fWKeFrtF2M87A2El/I/MPWsVccB8yCbKTPv3R5aESen8dcd05o
OjvaYFTEdcMHz5HGSh6CaZ2mhZ+t3vHdYkfK2LhvnHHHw3fRtJWRQF3jxYGwZCYd
2F0LbVA3llN1ZIniQGsi4T0+kSND8cGUiwcxEjarRBCxkG+T60/7P8mo+TZvsGQK
UWLjITfJHk9fZZROO19MeKfF8arHD2ddT7qKnjBrhm4MhOzzGe4wztFzhDYuX7cW
jvTLCEBoaWcjloJtlj88364ejAprPMaq5v5PiA6jnOnY25f1CSY7jQzzTFKOxqhd
dp4L3rsTUhGnd3/15yg6cyZB47wWFv1OnFK4Fi3d+qC7ah5rLUAZXpSP2BPQRXm6
dzWrmrVcNJU+NXXRlUYyJZUF+uJjEAiW3BpTpBVw56gqoXz/ZikA3ouvhwGIroAs
49KrZCdz5mp9aB+sVuMvaM0jrUf/VWLu5J4+9kbPAloSVjaBIJLAvHRp+0q9tdtQ
X9p5IZb32fy7G1V27y/DwAFLkWst0BnSD8SN/bYJxNPTRkc2tTAgMDfGnT4aNgDW
vz9pA/MKiMjvXDsjlkV9I0Ak3aHi1Uow8VdHRdRPbPpjfWwBChHSWJLjPtJn86pK
O1X/9iNlH7Bs8fJPM1cgDAYZ53pfTZx5L/pgfF3Bo3yPtX0xw5lgT5S6K+hSwrLj
z/uffMFssA0V3HguQO8LLnNSutPe90sRDv8IXh6ULU7mXbr0nG/6/e3hUO5ezryY
DXY0yzmkxSScIE+CYM+Ia/sWOm0Z8DiDC/dz1Y61erh2OVRZCKiAASygeD5DvvcL
/5VLso3SBTrwepIb7uGd9Ep3JYj1bUuzinz3hjcJAFzxFOCoXb6lzQNM+gFi0HOH
/2CwBXoa5CUN4vJWbqxSLMpOMWvMiStKvWKcoMhs2+1Gc/sBdGiLhLLbke7TO5GK
2Zr1mKGl3l4FyRmZ18CvzTCOVR3Cm/V413QUdC1/mDL5OUnh4s+Gu0cYQoURbjpN
RLR/fVmHHmgSbJUaGw0XciSuxHMNtvsZCvW36uPSUxP1O/X1oWpD7B/Kx/1Qys3B
/olUaVC26TE0rBzknsB0qSmzRxgA+9LRHgXpmSszfTlHHJd/HenrDLp8k0Iz0/Gj
XyveNY2/VxNyYihfMUpFfUwnOpYPcUvCDFd96t1ifN1P/YU4vSuRUVa3+WQrSWuP
m2bW0nqdqZpqi+SjDQ6wrOqmMbrK/hTGl4h5O/q4axjwKmUIKlrmPqRSgNQEHwQa
lFihLjev1lG5JJETs12cm51xleBGYU9/DQ7yJa/IdILiNVoHG4PwzfL+bZw4sOoE
lvSwLmE56tdbfV0LryEBWX1a7o88rqjR3HpDT93Mv0pn3lCLNl/QeZx5tgUtxisU
aRk9ezB0NlYL+TMdv3wxl1YfC7LnRqb1m774dz0gECCkAoK+dfkwrhthRBwVPNO7
sOgWaqUKVD5im30u3DFvXc80oqE9XysDvLeRdShrA5fChqoa5W+0sdIe0sc3oqbu
EB6K2MXlon2iyGGXkbkBbGjpVMq/pZLmdyKp1PXwaMnDgHvLpcHN4bUzEd9IZHBx
UhqDh5hdHlV1aAkgxqKZSW/0MHa2wq/dj63cKIODg9KMFIRAh7p4rsZ8um7hXcVT
EZV9/NgEMyR4hxbr1HlauXL6yN709LUkl6Htq5d7D5InMnj+/yvAVgToA9EH8zeV
bCSN+43oS4e/J5wf1TZ1T/akisyk4eiGTnG/Y0DS+3Jl3Q3UUGusMQQ+naahzXa9
YrYOSG73l58taeOBtq5/BuW2zZ66aOWlwcno4cctuJ7ZS4w65oLqjCqkOX6B09D4
qw3/NimMe97pT9m+msXR/zSPrkpJTRULpgo430PBP2oz6RqT5+RZItPGXaPtd8uj
DiChrWdUHq2qFo/9dnkYMz/++fMTa5pDASOHt+e4slkBhR5dmxDytBFqLKdXU36A
VlSPM711r9fc7ZRpZPIQ/RaY+7XHqjif8AHiNwJ+AwHcTsBxdpJAcwjZ1VppdDwn
zbo4ijxEWK5rIn+MoeRwWZZrykxjwx4ZT5lMbGbB8eieQJ596GgZZvRe3pa00hXy
YtMMPHsUOyDc48L259SxlnYp5tt8ETNcAhhwWUGcV+Z2kdPgHKqsCjkbqw9BFu8s
Gqs3iSMkQQibk3vCIEyQYvIa1TWtCUOX2ShGtIk6JAwJB4Zqmssfs7xgz+znEhF9
SrO6BV/CZtGB7XyECy4IKCIZm9AFJxLwL7f3/bt/2EZUiZ0Qba+JYXMpdykBu4xp
h33FFObfTJJMQRcNCdcli3aBcw50g+2tUIR8XUr9ruc1BYxeWoKLaYzHpMqrrJaS
XJnJk1EY6YQrER+iTND8m+11G3EPJ6Jw3FCUxwK75HTR446VT2Zht75eqTtU2TsL
NNol2/BgS6ADFiOQfGtRcHPH2sQUPzy7g6mU6u4rV3dBMw4qgpkcF8C4wU/HFg7p
lWBgOb/eEXFIqrGWSQqbhX1hD0h8SFCvuAeHYwxKaClANbojaw73uqsWF4M5TidV
Qo4dNNBdod7nsdOcUzTpu49nuEU8q5Oyi/9EnVicZKEOxM3NlcdT1AR98cdQL8k7
1ujGwIbZDtmVyqCPT+v9U2iXWfmmnq38Jfg0vJnX9sTYTgE9FBOEBY6X9kGHwYEt
bZg6nZiPkXi35Y7NYjTqN7fKzwnVfl7I0VfCaRAiZx1sbAGe5z45QT+6tk/rHO/v
+FVqwMiWKnaJiLbKh92pNIZChzlPi/hOaf3yRx2JtmPrnH+e7e56c7UiA+1S9KRO
cGozuGwdxqMJM6NoVy/DKBv39qum5YJKTBTjOCZJjSGt8eALJOelbOzE/7GEujqx
cqOeNA90L0ylcFstUr8PvtAt2Oxog+NEjZZN4InflsHBgvkwYA/hHZvClYHSyuAc
pJk66J0i3Pm+U0xwh+rEiu2UnpQb0W82dbBjeptwccvrA/0gkUDJM4tRvDRi/r4L
4RUq1d5MbrAdbOf3d/Hsb1ptRKsBXVa6KkCmhVwiwCEjD374xKP/XiEtcztJW9tC
eOTBB97wGxlbc2Rq0/vRn3chAPviLm3erwu4BpZ7qceJz1Wj5zV9l5L9L0lsGpEO
8HBXFrmZQoX88LtRdhnQT7rpiyq2TLnTB4WiT7I4wXKsyjKVSAVd5ZS8zJUnA2ts
mzPPWFYHc6/G/+c2L4k2qaywwmR8lBmsvfpKAiMXQ/k3oVexgReJFJCTCjybY/fF
G3KefcfJAwnlvYysMt87fwzbAopzh77GpZpQjSHN0Qk08kifMdLfrC1C2aEryM56
EowDs4NuChQi0ZST8SB/15uPz38nAlUWsAN7Vsv0FhQ7FVcnDDXXdNI+qraaaD0Z
eWSEk6MUWpoOVWAbsFy2Mj4cjNMVw0fU9hOaEhtRp8Z1h7FgcQymjZAhA4It7GP4
BJXAmXInIBS4CrFvSuzZkWiEb7G6E4TS4Hz2R56x5OlY3tT4f9rZ9XrfT811VJXz
hWizWf4o8kidYEF/JC4D7FaZ41lp5CaJJu6fuqIet30za2M+3NwKbJTpxqAVyFlz
eq5szD0j4zBFJJpF0evHV8XHHP9339SqvpwGRXhhVRbGwTxUQgdIIg3IQaISWrJk
UFsDq3l1h2V/m61XzZIQuw6rGRzP8DF5dsQsQKo1juwHI4nqKQXsdA5ix2kuZXJa
1nTq2MpHxPiKQ0U0teVMW1bhVkQtsx4Zrf39vff3jeQggz2RfG5OQddik4zVDnw3
PJJ0/1m0L6P3cORamTrYjCMRZUMVPb7GlHdBYzISD2Yc4EPkAS+r2pLoK4gZ+0qh
VgMq1g3IoJ0rwZzyW70hW6a1u2SxZ+dpVhr5IenG90sYaZT3OJb3XveEV9jJKluK
Gm+FNFfeUGcdXxuK6KH8FMP8xzwYEkCE2pG7AGyjZoZE80Wnr5HrkbmBXk6koVmY
IHxAB47Ihgg25ws4UStNOl5jYZSenrg2f5GG0tHImM2GLGVOLRIac96Og8ibxvkd
Z5WW4KDrICoE7VE1XWmUBjOTPY0wuoY6T5dbXm3lRLlc/jH9q2s8Hoj7mPwbE4wO
Q/x8c1N5Vl7wBB49YpvF8f6HfWcJ/XrHylmTk7GXQObAzSJYWOTL5qjPBP2Dllmx
BybV2+tqw4acFUDhYgEsa7Ri+A6Uj7un+31ScvrnwW7SbQef18tNqYCUYIRe2dSH
pK+PnwWXbHVL2a8RNl5k9zeXL56P+Vo1CCC5b5+AI7FpAIKMLLZKUecUAjfr6INi
AjVk8rbppeWaPEe2sddyyYJE8MgNMeRM4gKNFhdh76Agsl0clppTNNmVELj1GhON
XSh7FEpUOq38jgpM510RWrnm5bmUebGAfghTNaO2JFEKbpXbQF8i7RZY11YyJMMt
eGyGRpaK7jjJTT4aShDNG0Fv4RjC+QyHs2xUM3ZL200afKOYbzAeJatWs8DQLUYl
bR4bsWU9LaXhmgCSk9i+2jCnAhhgkL+iKnrYi1KwN1jq/kQeNL5+NB081yKkGlYy
xqZy7dcE0L2DW0pLDLurT/NszpHMapp1Ag4T3jRRu2eya3wZTkWnIc54D6y9t+OP
E54s6ejUJP9rRUc8dFf1AOux7B1qxQXmPZJBMukii43TZy2jFPmMbD7CgL5OBwfV
a5PeckPa8A0C9F0NKS/3tk62DQBnNYxiwhVKCEONj8h5qkWsymUwACxKjkJYFDGL
kpTrADnaxxqpT+62DHr3jse4K8HIZ/N1vy/Fr62CuEUg3SmZUo1x/mP/vEIfXJhQ
XGzxxSEXSaHxWt90vdBThPVluL/LmJnkvf1IiLYoIoUTvYBqn+LHoEt21uF0j2kR
kAEXXceSNGlD3u5nvGXvUYDb3sWhaIF3eBXJVNpayuVWivJa6TE3+sxuPcAFO/mf
1FONTsbd2McKawNddcu0Ih4Wk9kXxNBTfllcFh9Kp47f6KOWTXc38QLfx16YIjtT
bReiOryxYKnoRw5BcWKhrQZsu+Rd4NZjVckLAkV0ieSVv32B0PniHBjF4pV4/w0q
WW80wTCZiks6FW7IPEV7wL+de0NcCXY4Gbi81c0vJD62Kp/aUsIRK3n5iKeonOK/
wX+horHVgiub3VawK04pL7nHuoY2lBba2AjvlDUoAGVgT8bj5+I5QHj6X+o7RBNc
cXLptHblsp4JkkUQ4Qumgy7bJmQjVRXQBZv6y4I4grpZ8Y1yvMFNf+EIDwbvJalt
a+IVaAY3y/NVogoAvZ1X61KO6tfV9uS+mgAFqPBn0Ag0q81KC68+GD1JsGSG+LVD
gbyC8No0hWLwOPuZHyoNdoH+GDxKU/yk1g/aakQpYyLfP1ISpy4w2SvnsTXeSxii
Meu/73fqeoNNoVPohJnpDTwp+iamr1JJm5ppx/uTATBLWffcpQx+5ecvOdGZpF4F
GCh7q/HE1E1LW5Tsm4v4Lm8pta56bRjM/E3zuaWKByFnvP0N2ezEXi85qxWPrRQg
/0f5F7xpYFUCglVCIcK5JdTGQkE/Xfqmtn9JlxpJBBY4TWkdUbqeLDPnl9W5q48A
G6PAN9tX3zeSGtUzGoJMcXveyp7xbPQkY+fSx/azZ3buLLBj68D2gJgrabYUbclD
kmMI7z2iasWN/36OgQjpUeVUdR1Qp0IOGfxA5SaERjUFgNNWWiFz3fmUxTvj9mc/
68G7Ith/CSXHcRrDt6DgOWYiC9p3RipXNhZhrqnr0J751ohhbY6YGkIJCHjrAY/0
hX0gQD1iKxbxRCDGhpHUcATBIk54KHsrWgv1eXD2dcSsXtxmX5a8F2Y6R4mk6Mtm
HlcUt83KB0/LcFNDYYN2QsOPrIFjMrSACS+1UW21MXRF6VwBaSOhkMjrvTGa3PQp
b/ap3GnpA58GRCmhbr/+Zc05t7UxV9BTJd+Sy+1B3lUPDWy7bUMLVmpw0E/BVQ3h
i2kNoniwgL+62sdFv4dAUXFsADkUDf6ZRWaB4bwlbRJYkvPJxaHSSKRyLd7hEIYM
q3uHXvFEobj9G0v+NzRXq90bQFffC02xBu290weQB2v6E0wAUvuuipIqBuSvLklo
4pNJ8iMKzIGHF8oUnGqgtfTYOnmXGI5peVWXpvMkHPbekoe3/ZMhxwPRAC7GYegE
kOYnnLVr1EhrDgPHCvwxbpph7AV3N+g8tzgOrb/BlVzVZXU2BXNV/GNK6j7xBVMI
XmVTG7rdgNj3KyFiJj2NBzPrlFo/LcFux4S2uzk0ySXSM8CiDAtRCA1ZYiOzt+Hp
Pc8NFdZhz69rmqRQ75UjN76pMiqmsi79/83byh3Vt5uJE6L9gADkaM0IYD2SaFLC
urqlCbeYK+tpTUwV8u1jZ2KMie4mzPjGJ5XOOE9mtyda5+PDwI7KekjJgFfhqQtm
BuZmYgU5tpBsuZUA4o8ebPpfvXl7CzhE+2ctGUX2VgIodnJsfhq8KO4MuXDrUeCi
24XkfddqP9M9iy5i5v7AQb/krcLETVY76cOecMi882AMdBhzMK336dSLLluDGYyq
w79NYvE0IBoYZdFUVJvz5jJHswhcRVfHBkoyOPJG34NeWyNkkeJmUHdrgeAgV+HR
kURqeD2/WLIeX/Qs/n/WFAN7KT7Y7/i3+AP6HfP9xhURbZQM4UI801wAXdv/iH8O
0YBP0CCr+EAVZZ3R2eO3ZBShfIQqU9Z6DyU+Z1iaA7F3PHJFLBCSrbBBipC5mxJ3
M0igZFBpI8NjuM5b87RmkekpFaW2UdU6Jnzy5JmWivFAq/5FRq9hwF88JHFM98sr
lLNoMAUXca0P3IMH1OPSMrC+1k0+dY///yKvdoh6IsfTYXDB3by22x3wXUnfyATI
BgvV+W/AXD5oF9kvwNIP3kGROEGixUNPG5z8xDs+mSPyeWrwYiqXlPEl7rLcehCk
AAP7j9y/0nVDPQ+ViQ3k0R5hM2ykdWOksMKb6Vs5ER7eirWS7mMI2cZxGQkyZC0H
v4KE4mIe3I9rSyXKGKdDv3Cg6eADPublvrhBPPaCb4XJE0fjsP/yd8vdmGa8AXzP
fKXRrf1cMoOKjFxnQIRtABMHj3QkUslRkly9G3nvtDrs8zHDm8nQgPatMYCv9h9n
Rgqf7S+6k0oSVhKRw28U8zK/36eXQUpg9aJL9DoPuguQTZkGxQcBlEHK1yzJ/MrZ
ghmZS3bMzUdaggCrKVU4X1M9qEFzus2q0M+6qTqU576t0Wvv4N4JJKkHFRAFFP3n
gJVcr6bH38urU0/a7qpFT7OKefjtqcnSCHYdH+pUNz20+/eb3HuxDC5Y6umeloX4
IYgMb8ku0K9lu2QjWJh1oiNTipY0S/avvUiNncWVymDHH7ooY339YUZuTCP6/jh6
p3oVBc9GVLuVHPglkCnMF622dk1pmsm+wmsg0cp3U8R0AnGo8mDZhnpLo6xCeyna
qz5+H3N4gBpZ5ALwfMKmVxsv/7hmZT7GUNap4k/si3Rn94vyXvlE87Li0NrEPCGQ
O/QprkW5teDqDZ5fl5Cb/N/fV9obRIBkF0iXpBgliH/rFFwte8w4SvclOyZnDB3s
2KCUKSUXjqgnVq0o6XLnPgyQvP2cvRcFEeSrGuQf12O9zoxwwF/JiG5puJp5qmiz
/mc7HcuCHOO3HW5FATN+5JOoGvlWvzvq65/Xzh0X+7va9aLE0IA+gEuWivMFASlK
lgunIGoJmtrVPLm5yhJUQCx7yN0hS2ZNZAGw+BDzEXvEv289+Ot69SAuBOH4u5qQ
DXLiiTgrVWvSBzLZT+xlRb8q52Bw52q6l+zbKBgR7dUXNy6cV6hGcIfrkYjWeHwc
Q1TfgsqqRWTksgFt4BuuFQV1U2jXcjQsY0WmO3xHVsg6ETnru7YLykQC8izV87/j
bAk5d2tXnhdp8+QZEImzBZ4kC8a+sejJi1uyZRLS1JUCGSDUFsCK+d3Sgu754mqp
7BoPAiIZbsqEJ4htNyr6OOt9ZsyFwE8WwgwrTqp82XhzhLdSZLMTF6g4mWVxBN66
RDq9kgx37sGrIgDf/W0Wx0IYu68ieGvlbIJgsuXyqhY9my+f0l8EA+xzQ+X8fnCC
m7ScPAb9tb2V7uDSbdSRe6xdt8Y4uZjsSnSbXyQUqQ1oApp8FDf8W1xtCpVKh2OQ
q9S2GocGZXbUEAnCA91dlGuia/r5tYLwwyvg460ra+4TJ7sn8HwBrWNAUvjKiilm
1+bWEfYfT5+GY87NmBsMETId8GNxfyoRVU0sF4b+XefrujlI+nkDvxofP55RcJLe
22RUC8ndbWzX1rZXjsVA5WZSq4TEhzUPoUE1SCh26vtLka1z5TJa9+wtB0vPk7ko
YiKhIUnPvrbWPyM3oYUSq6gpuUzJPanm9OAIsbQahr19pdyQOdp4U05JmB2FK0XR
OkS+I9wTpqc8xMKBUKn0Z2/H+Xu03uWquwoVf9Ui5JzbLwgoT/ivkxkBEKv65BrK
prB5AOplMDKPQaMtMMHBC2x1k8A39o0zoo+jOXom29++I5lG4SVN/Va0y1MXkoCK
GO6EyXe9Tg1ctr4RrFik/Oic3V2Gy8a/4+4U86Ua12fVieqCuBE1GO5IenZEHh/N
/xEKXEa/cne4Ailr/DiZP/GXLrZejPO/ECZ2Z2Uliw9llVvYjLTxfUb48AxMjQVw
if6pf18u5HP02x406yd8B1mUz7yNLtjTfC73dUEYskZlhoTggT0ChfOM2OK8K5jk
oGXei7EBGSr4Dbr1Oy9VIJW00mYkhYLwMRM95MbFm5HSDk628i7TFjjfZDIlaEFZ
/+iKr61xR9+atzcbOgQabxy8CRkGb3pSSA4CUc490K4OMf3adx+qCNLOLBAmEGAm
D5Y1aspXlu7sMkOs4WVaqNCaf2ZsyFuA7GEsf3S/uw556N9+oo/DAoFffpRFU/C4
sJGs3xb6jzp8N941hB69Ru86VmKL2Z7R39uBF5RvNMZ57sVi+JtN73SSWqSZcbST
uqBZVHzWEHKl8GaooG++FncY7hc5eD0jIkE+WBSwr2NDuXlT+x57janH38ZslTy+
m4v66WgEGTz/qLt8I3Kj5Jo00TwvFRH3fl+7k/BD5f29d99i9hWiVagzreF32a0g
iUcFWATBI3INMRzsHcJk1mblOW+hxUydmej0x+EbAhPxCRxFEd+pfV2r3tpyog4G
5huH+EeLhfUBy8CHsOEcas/rK1258MkMxHeR/n3ozxlRqhA57njn11Q+s80uyjx5
9wNu1DJKXY+lsK5JH6lTsUrCC45rszTFblTR6eWS21yePqm5jbXISJUB41rZmynN
9h1Syu041mPC+7bsF1+1iJ+ZVaQd8CNUgjj4WrfbzLp7NSo3evoOW/CzGsdwfqHG
PgEoUNqDFSVMlMaa+aPEjRHzccvgZZxuxEfZT8qlT1cXr2DbC/DZ2D2HGXPN+ZVC
g8ddaeqro0eEHGV+eneGE7lkjNfeZDR5oHEeYG9F4c8HbXRYY9TPZ9lredc+feFY
OwrupWPHIg9G7lH1ZYRXGBvpVZtVDoLovHDyhar0ynexmiCm5d3X5fx8Ke5lbdyR
hnQAgeGqwdTDfhUpfeGEg4L+aCn/ywnx4GJN8kuh0SKo+hIIS6x2UWg7rW0go/Db
PnJiDFC4YcOdN3lzHQzJMG8JSExPqlrRPmfEl7zod9F1W6vHo+y9XxfPgBXN9HxM
QskBmfA1UZ0IOpIQOMNJ9GKoKk+10UMra8aw2FSuN5FlsKG0qBl4Pz3N9rGOtq0q
cGDgm0WWIJARaINCCFcwpbJSZ4ZveRu78C7tduAkRa8UmYicJIWgmYsiJBueM8Rj
K3qewucUHyjhWqoZahaTkHZ4D/AnwVLKnS0tg5lL71Nj36Bu1kH1uaP41uGJifRv
FRU2DAwZw/fh4sROYUAAlpVkPHNT8/B9dSfL8X+COGrNU/ZUVvqxLvZtVnZVDRMQ
SsrtvXmDmyRwcTOdTp9L5g+VSQBp5KkF9y8z84By6a80qhUJqPH0Uy1Y2DqZFSi8
HSXXAd3KhAfpyQLKKFhfMc99sZZ68Ofy8hPN0oP9twhjhyDKT3cV3mvX4451m82a
bXdrGnV29OjjKJMlqDhFQllek04H/HqewTsLEsUb8hAJjAJcWlnUBR5THqwUValX
XD0WNn4Rk60CjklyZDMz2JajTKyhkk7Si3XmyQmouu2niLYZzMXAFxw9M7CxKjd2
+3twmbiE2uftLBS1RKuJjC1sXZYyzm6h/0F4MnxQjwF/rZEu6l8Olu8lwOqMeC3c
nnp3377b7lFszUoITr/tNTa4pdED7CKXtkNBZsaUbYjA+MbzHOvWNlTeW69Menv/
PuxiUaiZ4/wWPX6b9ja+r1uM7ymT+7QZJ2Mxl2w0PnuwdkHjYbve1P+by8SwoZHC
m9Wd04XUR0XpVPD3ge+/aGiMypcqvMwgQOZKyPQ1Cx9yMtzV2UDsR07hw8CoujqI
C6kSihQmINLbhjZm0+zaSLUHuHYghW4NfdNwC0ua4vxjpcHtL/Vu8GAwFD42zy+e
OId/YnxvqpC/4TMb5HpJTnihL73gUFs1UHJEiUf+Re0yfVREHrBRYSvd75dOsmiL
WeA0ubRtxx6HJjhh2m4QL6cgFoDEPeukp0rOpQr4MVWHt5HgFSOQ5ldja8kGOLRs
y5XEonvrjsI+nFwjNsHYUHtxWY21ZRKIx1NuoaND7E43+sYyjTpIcSsmT4LSA/4Y
070qw12/00KDjjxVy/XzhQ610P62uv+SAfmWicq/IbH4nPkWHLpyGTHhSTrD90bh
7gT/1T3PWALUhs37Sq1XVcdrFXcODqmgkSHxNzSTqqgGBVbp2HaTOZfDp7q0/aGL
JNHJItcN9+/dpkVj/4IU70f3vPBrKgR4wa2uWyXaZdNK/+dOjTud25wQat4eRQJf
Q06hX0yBst5hL8V5x+pmF8SGuPSq0YS2GFusoF8bVyX/YL32X+tVGSzFt+O4lCGo
u99X1yVvyXkzp6Pt7sOWu0Ln5icvw1s4ZHoRBudv2wiORE96bB7TahVFnINZRYQp
95SJ3nSBZkHIIaVRswabZf2ztxMFUeT3L8hgY522PNXE6QyDSTWAXCljm/eQgt5l
9pWcrQykcbk7/56qRL/F7t+BFn1/e7pRVPwSxWvq0RhQtrqV9+axUQKY7D4UmRFS
xIuQloi7aah+uHhkVjFDIkYWkxDJUQnKiH3h09zqIj4jWMnBYslJzdAGr7AY10NQ
OTN4yttHP34sHIXIOHeSm90xkN53q2Eb2AnAJxcPHaAfwIQHkmg8ol+/rKZd0g8z
QSUobvHHAgn+ECge4Q0RjePE3hWgLEZE3hU1yOA6r0ytf5UO3piOYChlB01osNEW
bRf+FVuUvqSFuAgzIcuvA3Q91cTxEBuyOZZ1jszgKBLn14dUc0rUuEICCVAJWg0P
nQoW9OyZanPYPMcVvABfsigvMQPJh1UQmiYj2sD6GMArZz2lXu9Cl3tMqYHU4KAz
cEulszm+pUZ9VZPYL3x8HeSeWy/8bmbcYs4phHLUmTwPOLbiuDX8SqEZrN2ps9s3
1Wa9jEUAlPPq2OwaNG6yzS+gq1T2D0Z5I8FMmRv+F1yTD+fFGJR2yU/46Eytum91
62cvCpghiNWUcjK2EWwGnQ==
`pragma protect end_protected
