// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
YMN2CWbMzaHd2xYxQItgou+wHHFCVaBgTpMGjNBIIkhNGzmqrA40Z33y6/Bj5RuvXlOMwz4OiDgb
x6YNKX/v38+Wrf81I1bv4wnfX8UfzqZYC2fIZ++o+VwC0t8r5iXSxNPseC+yvi1atoq1bLjBsPvY
7ror5DrcwyXeoI4rLH+op5kxjSUHjmxKDkliVyCTBQZN1sjEMEIHlF9PkMV0s5iWiJa8UenH8pDJ
TIBLIEgWG8O87TXq8c2dbw1DT8rL8GMGkArY4Rmsg1r8oNxNJ67RvZpY5JOjFqI+vIt+id/ndaJK
R2PFmS3YxF76bJMxFeI1wzBtQBC6VA3hinQngg==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
E7ZYBUh+pBfes27Acy0nYfflEzP76lw7oPEMui4vCHnTU/iJrbMfTfHb/wU4vYn2sORnFvO/c3DP
pbwDCwtRQ5wIpOprvtbYC70gadLmm2ij5D/Ktr7kNzHPquzjmvk7vVVOLbQBPUqwlFLFLU51rlWI
rcNzuo2xj4fftPgtPlMyr0kz4qIcX82h4YkpTyUMYXnsr3s0cSVYjsuUVLMt/w76YhgEP/rE6MFL
anVW8WABSXk4ie4H8MzxOtrm6mio0thYa0D1JJScUOQq3M6cp8uPO9wrH+QDdl7z1GvJ27eJHfCe
ozRyeWkaeYFLzpKqQWDsKuvrtmbtv7utVWpOVvd/bFr4AR9bI0VYBdJKD9iQg9CqQMA41j0X69DK
MWi74PQ3kGrLK3LS37LwlklGbC7BWnjpSmlWGZcKRkHAgrXcBoIkJB+FOK544YWcjZtJqw1ias4F
OXAVeSy8YmMnjzQjjvQWkK8+0iFw1u9lDHLuiFDZuqR+zT32tR9PO4r4gZfLGCx1ZQrwsXTvTZO7
gv8aEYBzMfyEdsADVhGcHtB7HlGW6TbvAJuHNd6/btoHtoHmZiWEiAqWlyrgsxD9CWze2ev6qeh9
+zQhlWiunKV4uSi+0nKOxQZ5swyEVN5iTvNUjzrEtB5PT8VL6DV8syu1JIEjMFM8Il7tRL08m8sp
3MQPcvEc0iB+S3aedkWLU7D0sXEXpUe0Kb9jlP5VSrSRyYrONZs/N2i6FN14xaTAI57W7voH9oMT
lbtNVeKMD0ccOFGk/EWlGIsYO0SfD7/S2FAvgHdxPogs4m1O5SK6Yre92BMfYObrDcityvf56hsS
BE4ADMREhERamFq+IZov6R7Pf3oUqET9/BWISBFQQFwSg42crls+9MUDx4Z3sOlE8d+uae9DcsaD
JoLg8W+caN3huZA4DO0Yq0Va+xSuq/3885bOkw8ay0Ca18YoO9uIw25ULTVleDiJHzSM6U3g96pC
XgmNvJKzc50iW3LgFXgfhlfNlW1okRxozUiqPA00Y+JIza+mxBn5aPD0bX2C3IQp6nbArineI2lg
hzKM8dBse8SANl+/Tez4nTBetnCOX6CKeU545gjyjY2NZGiJN+tVUWhvDkFCuxgwTeDx0ZL/iekR
Ti9X6hWv7jT1RXF4l0cD/sKO9hYzgWzdvoTSCcjMBat0mv6auzsJN5P3AJTwfcx3Ua1yFwmOXLQb
MfBhumZz2h08MSotIB4KwfHkPC+H0kiCjxt2eiOzGtYteT6wVoeFHVHbDMKChchuuXrdUKwzLQtX
OJ43SuTZ1gl24Pg+YoPt3g8xZIFbshBYGoDzhJZmJzGh62yICoGato9YwTNsQ6k3FsiWV49d7uJ1
c0+6OItkhR0niUif/9e09XPJ0GMPNMn0K54TUdKtadKRzGcT5wwnN0E5q5gOXRwxyEqc2SK2dP5z
9DysAzi1A+sq61U9kZTRjev+IVd0jornc1iRweTv4QdKDUFmgs6JRcc8uFVYN9TI3FqDe6UaySM1
C/+P2vuKMSiq2c6a1OcgVfpmILTu7ZWJO7Dqf0zjSpAVzJQptBezebkX9B1VmMDQac3PHIEFdPhS
/mSpk8xxRf0sKinbf8WxaIywC1hFk1s+Ed/NAedDezg9R/LAqPSiJ8h4spFaW8c70nj6p+nqvJxk
r/2SfiWjNyW/KTxNahejG6EQ7mdN13g84fGU66OvMewaC8TismxL1jG1YENfbwmwGiWsNLQRZl3a
ckNCgf7I40ndHO350lUwt7kmleXTHrvrjtXOOWK33jH8+EVq9gZE+Wb+XtPw2EZVs5oa+7l/0L9i
fM8cm/aK0RILVvsQg+0ehKznB/Ds+ur9e0qqSfbGdEk7kS+dCBV1YNygXPya8bpPsXn11//CjvrM
0nWZ9eOl4q4D5emf1vWL7LOO3HXomq8zJfS5pJ9OgGmNBrQ3xloRX05LdUng/n4qioV2/sYhlzCd
vWE5+eHCXX3Y4YAUYFi14oRRWvbCe65AjVNz+iDCGr8N/9b+3yqS5O+elfacDEy6sQohiRuU/HyG
6LbY0dGmaI9YAmbFkxTfzC/zqABLdjuq8jKJH47B9QpEjVyfeJfL0jllPTjOy3iEwlBVX4MvLhDZ
CWZniYkHz5FH0ZrIWTbC/AFy8DzaRvrXLFqTHEli+SRxZd4hcrAiU8uNX6mnErctE4Xtah0r2sbL
YufWRABGbus8MuT/91v3CUikgsAGoym0aLeUAt1V3jLNsxsN8WKsVVw+YUIyQEKzZEWSDjbDfxu4
OP7mN391dzHzCHCIdBheojhHwCoJhub8yoi4uLhE8vqj/x4JFYcsHAco5/Ca9T1f6ecaJGST4mPZ
nqZj3Ne/PxUmb9n0UChdchdGfW+xGHUoKuKFap6PnLyRHbD2uoRHHjttEzb3HeXGWILwuYl5HhgI
Ap+sAOfjLpkwdx8wQmWDRrqYgirFHhAVSfU8IGRsChfJJNcvuUFSbJLNJaEpBu29hOXrMicmkCXj
3efpGyecyDgOZ4XPXL5FrbawKogcoGXmp0jZSgLxLASPRjp9Zy2txhPL2+9KJBsUFtbz0T4z9Ebi
mg2AvxxjKB+uaYec53APk9FagzOz75c38iSaw+IUtQkVuw+CPeK4YnweBDsQb4tEQI5BtkT4idoV
fnXcNN+voSgmaP/jSIYrjd0XJkNaIhTaZyL9rHXjlCR4adHYV2WYDEKA4+uf0POfNgP2DXx8vZRS
QWoeJK83tlI7gL3FhnGi4krd8l8mHxJTBgypIRe+hD+jmqe+/dTfRBRnNxZRxPoQcee4H8DJ4lWm
GLVaaKTydRaq8TyGS5PzK7Z8+Wm23U/eTP52M5zzGFmU8ttyoxU9ThNBM2Q+YpcdX7SCr/RtnuWj
/KWJ6wDI40LZBmk98HjE5J6obMAC1GXQNm0/A1nPGb9ztHHOn41QD5d8qctCLP6loXPGR3FitWWl
3KNecqqdfCmoyHfSMCzoKDoRI1X11xlMuz8z3N0rhXfgSchNGQtoRT4ApVdXoqtIH0hvETjqdeib
n9jDQK+rPTfAWykVS4w/IIeJ+bTdN2750k9Iq25CWHyboM//KJnDUKRJjtQlk+DfAuklzeu2t04W
W2tJriEZE3lF4/0AbljBtc8WdJtzK+QHj8TsNHMM71Ob/aeBDpSBul+1NtdHSBtcqcsBetToL+nL
BaB9NFO3sxM6jzxRL17hIVMqqqScVUHcpjr8xtVftytX8nZXRAZSWXfLYXyxyOBAY7n2gPm6dMKQ
jdWugNNoCz7OF6BhioSeuG/Y+fgkrgPZhh/2/UeDbPZ3a5g+jmc6DsVSe23Kxnk0ecWet6YM7FfF
AY1E9WS8uRppOYHNWmyDIBk6E+Fuv1f4quikUKv+1wjfmR0U0oFMAy+PdVwsLUpXqc4TYh5YWdHS
JXZ1g/F+PqxN8+IURzFs7xwnV32P9qEqs1e4OVGbAW76/xI5V9RfqnOfQx0yzp1LbJWAUi3hq4Mj
AspNVjWtlZHzwm4JI3zSbT26ZFOJ0Et2xDX7vYg0095exrnrKFnYfGJsF2DvEHEEKJQEob2iFqf0
/A0r2ULnUJyoiu9aeZpMrGduv1aWMVy1QZbMMJpj67zDQVPDPUkMZ4QGi0cgwnbqrxRdkqxnXYNu
IIJHn6SkjbXD5l3sr9RxTzddDAtK2HE8BKeTzIsUSCnJFrRHWWHlAVQp5xib5uaNlkXaetf1kDgA
+NJjHHvlqRLS79Pfq98olzvAPz4Gq9YvjW0k+qAnzmn4+l1LVE2qRda1gtA271gruGYNGFDk8ajp
QFMKP9cFSK1qsilvtBu57ERfo1BJFPyvxsv2GG2u61uvKVd58O7pTVyvJHReLHqFB/RQ9mk+R8KL
WGAu4Vq5RUlJFP0vLUut3G32NPdyDM870KYZFssUesD5xVz9X8xHyLX0xCYpY/burCUtGjATSHWf
UKq9oArZwJ0j1UDTr0BY68oDNqoMq54j5+cpPKHKiKSDb5MGRs31E9/BU2eAE3V+UL+yTKwZks8n
c0ASrCOcUMsbnO+VNQJvG5Fj2JL9geLwskk5nveXxAlviqU45mVeBgp12nus/GMTwpXyCRI5DLmG
AR7DtZUHGERgsvX6aWBhicI8WMeB55ECd+Knt0484rZ4zijCTBpuLB/s++rA/VWvHG1qgZwjHkyD
vj2hNuI8puZjTMfnxCayqTAA3+0m47SwBKQEaNPTO4qEkGM726UeeOwI59c1AZDtg22jKH9AhuHl
LqLlccGyNxuHwFEcd1B9yKbKh6J/v5a+KasikSGF4j6q4pOkMFyK04xX7r6amD+NvcWcn1gFZDVL
Vo59HZq9FltTuZ0CsWK+26LGBjjKagB9eLFcYtDGh8w++W9QZLUOHHlOYUYArDHIhEOPyfi78n4l
sve9SJavFHmGOsIja65h94ZfdgXRBYT2yzqUBPk1+DhF66FzVjecTPxtH7mPenpzk/XkLDPp9Hyp
qLStV8yqPG8NKUREm0gYLnxsqiDXgHjfaYZNMeKfXdsbGh0XQEsr8cVafEtX+/DJ0teWDIropdL7
kxGoKWJEcNbQBx/IRJJO4fDpkDAo1JIA7sBGLP4ds3EQHR3qw2YYkJWHswCapvTeJ+w766jp/qZJ
y7AofU/IwHyUuKc5A2oa2xttQgDaIq7fGPGThMH0X1hYNbMYUhGxBcW28osU3la7EBEe4YghBMSz
qDHB+z069lC5HU21lFsgab2KAsn3ZVc4e8+CVgZd0n6fZEP+ujb9ICepKh5erUNc5XEbFNWtijnc
Qw4Gx8V/90ReEGpM4sbjLjycXIlCrExhv1EwYhRHVFT/Nt4jGmDEEj0OWGNRFSpdceMkAqIBbSTn
lNxBkwwZGsywk4BuCZ9III5JLyBjTDeM9rTDog6SXpMdqXww0+axKhnpBJqZmhxdQhat7fOUR9VE
AHHvSokxPZAhnI3hFxLg0XetAYs1ak47moyS2xnwtVRZgiMoeHsMwQ+Qs3tP9nqWZKbrpOvMfNjP
krCj6xzaTHScu/8M5Twjl+NaIEWa/iLDHUYU1FlBX4jZouBG8pF2h2SD0oN4zEh2UN99DtMm47IC
0oycaSHXd9zv+QlgQypoyrRKWFHEu5CFspfLcuNlliCp7NuxR49t5LgEQ5jraKYN6ULngUKpvP26
riOY5kCIjSO1YwfB4yu7ForVDgTA2mFSIkd+ybro13EH76Oh5Xank1hp9mbDRSIobEXce1qhuynp
8J6+h3TS98oR8gJgyhfKpEi2B8sb6Z6a/+5W76P9H/Ao/IEyAnPkBuvNdVg4Oz9oWHhosWfafyqo
BNgvQLBwJgdAUu2PhtmGTWBP/CW4TSLWZCVMaU/RCsWSLKHqmgZNRn4IkQhdheMNHJOY/TYmsKiI
Gje99am+jxSVU85867Nqed87gyuQpk/pupSi2WXkSQXmyxBy6MmGisoZiAEYK0nzxaolDc9XqQsQ
2aXKYf6ymiBBx5GfHFrgGYDNhqilfCN4ev/rpNVzKGla2jbSKPPtlNJ34txur+MZRZkPKdzyCYKf
YP4ayVCRzi/4NIhQZs4Le63O1fqV1+Fsp+u7FcdNsaXM56vER4vR56/3O6IJUrQif+V7g2RuG9Ob
gwA2tdN0l6yNlzzEwg0ZNXH11yYJEuQ6CyI3qHOs73/7onZjz1FM4DWIfLcR5bQj+v5TaAoKYTK5
Z156nSYBKiriy0S6k5gzcWcZSHKiLhpBBY3KugtHiETl/LYJzFY0QcgAbkDO0cJs/v7IXciAzsqB
QVvbaJGkL/cOiP0YhJwdiIfgqVlsQ/+6b0nljFAG1hUgCsVcVLhyVfO6BbhD2P+WhtUbFuCahjku
zQ1jgTCR4JPE5/kAapC21d53hr/lCRtpB+HUNdG8soNtQda8RIqG8kxFLe/qaUMMs/s5rtd5/uNk
Pso6Lpsy7kkbh9qZXZxOtKk0XgbAIRN0aeeIutjvoVoJ/F6DVLwLngVWXVjcInRxPYRylEGCToGk
ZAIwGhp3hmk55ul0gxj6QoweB4ULlqd6L6FFUTWO3GG5FaQvFQiNRP8A8fBnCCmYggmK3/TdPnpr
rMblvh+4nvNN5pLaJd6wyFDtdjdOFaaChzEqMNwfERcXkZFp49NfdgAFPHp1k8OJ4PWHOWc/i14a
xKw4CXyT6cVk9hW5PF+gMNuHMkam355d9DeSI06hZ/orKzcntp+EP4gVbMQOQ7RmJiynD1xsaJDg
m6E2NJ+hqiMuQ6yWYNIQPycSBAj/E5TyBmfm9+X26kCXbhgYKfSNyUoWSTFQwR0vFAEIWUyJRm+0
tjaN9IFvdIFpM72vt3WF1fuRLoQNP3Umd1rRcFKp2b5H/Sk5lf34v2aFLwRhnE28MN8FsME2t3VN
OJNs1dGgWftE2dOv31YcRZiIRpsyNgYw+pjxBq79Sv2zZQBMPs25jt2bNoPWkgkecbfSyRijRB6F
Obklj7DiTXxUSecXusbxbPTEnqt98YYHx9jzhxitRVPzV3Nh9Jv/Ali/duqFexLzP6DJBPObfo01
eotwDrHi2MAur3HUopEdOhBKsbpBlyMGZtgJ0Ad7AORhnfv+XdWNvrxODBK+jRHUyTfRwyAxCcth
Epps6AgWr1tu6OQlttDGkj3umLcRk01/qyxdqtXbrobjOQ2/OlsTLRKqDQHwQ/iRZfPP3axV9TvG
hi1jqcmhFv8gcF3yqvkXytBoT3etL3k4TqWpJYG80J/fBarXXSxNWk7SpdQOyVOS3PwHU3rzu7GR
BK3bdxwilJzpCXrPuLMH5p1PolxcWB7O47zeOZ+jWmejzalAKY9iweq2sMzjxy31ByAtWJ4OII5/
uCH10BvzAudAEQX8iYL9juw+dmgVM4oqXzanqQKdcCyix6A76v1MfmL6imRW2thiSPnMqjFpLzkn
vARBj6fIPaPEMSpo2fFJDQpewL06jsLFUn2fJ1Hh6ttr+sAv639DJaITOPR0fnwfpfRGt58EFgFo
mriv6rJGghv5+D66CLGfbwoBUYP2ElxTtBdM2s8UCIE/Exclfw5OwcbU4lLQfB8E/o5oKdfaV/R4
qsrnqP3zbyuBGJN/Kdl9QY1p/iH89qQOAErOaX3ZeqPb5fQMeISY9UIhHu9nKuemuH9A3bHbKLVh
wqb9ZZ8CCDJOJ2cykKHZqXo4atYX0+jtjK3TI3apA3Zm0dkD32J7OIWvuCzYa6qw3CFtZ6gOQ9mB
ZBXbEnhy0MykD69lwnlIsO42QfHOR0n/4ArSKzrw/d/WZqj1fjijdg2tFms06YJ+Ib8EMY04kkGk
Lqe6FieDqQ6gQETCRQw2kjviUZlxYXGaq9NFcMJF2W1WiwShWLgxNJAOiVguqpmiS6j3wX2/RiYA
vciUazj19SvGiQiDF2k5X80YZTvzzv3wB2Gdp1P2NfDtow6oUWcyKoR8wZcbRgfHXNw4mEXcF4Jx
dO5JAZ58tPtsXewyBqK7eH3Ew47hORRwLFBegSJEK/HU8xJjQ/XDQm02IdAMVcITgD5RSrBjZjHG
V6EekQmh5m9X2dzp77F8mvxNPQnmFI412yga+u7lwVYiGrPayaSboDeQitPgi/2jbJumS9ny60xT
tFlrIW/I74Hz1a7lFx0B+f3hg3YmRpMyPDOT+975i/j3OCp/JXiA50aeKhUz2yjoIi3wzTWIjYpl
niCcSPvSJZZfJUY73e8lIMZEK6DvSYXuiipDaE5ctTAsn+qfGqNgh7aYr2z8f1nAIxWB/x55tS3s
afC2TkToRQoog3MehAcjvadwrOQo5SrYZFE5tvzsOoz6u2CWQzobADgNn23sxQF35TILu/cT31fV
5WQBJt6M1TCBa+3DnpKzlTvUyJdHlL9QCgH00rkBvetuyvC3jT1K3tbRdxNUaP+S1k8e9e06x3qg
plb6Xl/SaZZP9CMAPGXLy5z9HnUbRz8aYrsfa3WaFa6pwsg4saTVzlGCogf26hdEyvK0COwPFUNL
G/Gf4gIs35xF/b46a2D7oUJOCvZ2BtLTKi7LpFtuFgP+key8mN70/CoKKVfkut2nEgk0MtYWHXCH
JIpN0H7rAE6yRAsYZgh2WPxorJdTKsnp7UIDe5D0rB3ZpGu/st6v7SvnsjhqrxM7ImWy4q/KGtN4
EwOclQxD0rBEMOPfHVTaQ4/Ox2mERXXlgud0BdtW8QjSkTmWaM6kYCE8SHh5XZq1h2l2f3XzovPM
1G12k+38CupbKMvQVocEtJbXWafhGpAl7HT2FjK50bwsRbsn8wzvNzMg0vJydqH/jOg+IfIsef9S
HbsB0ByY0gUGxnob0O1pMu+vsS/kBVrfBKPKzNLWnn65wqC9EHleztXxTG5jOkjG1DV7YPLAg3f+
VlmbTh1jgC5Q9AxwJbbR8D1SW+rwGI32e6UnDjv7fD4LnoGDPben2ArKTRBosYSsPgrF3UgbKs5t
kBtoGGiFvubQVkzPrG2xxvVUapHaFcQjce0xmbrQUHrhkEQKOXvHrn46W2beKZYHhmajB3gSKljr
6i9onwx6Bx7uLUzza5N4dUJgJv9CPDiHVKCTmStU1u/3a9SU0T9kuFDXofUJ4681qVcxQmFdYq/s
3xnuX1+MkGKJUrswjIH1ai93d0UmndXGLM6e+Ro3y2Z63wDQG3zZWlIJryeuFv95wW6hxzlUarXY
LG91p+7aNqRkVuyIKj6QyKRUwjJyds97UqjFQJpo6WUZRCNKdvlskcthwQKNb21Um4Efav6iOW4O
UlbKO2smaR94syMbpzez2366xjGY2XMRQUNwf0RqgjVJPFhzay3+QSG16Vd3d5xwvWe0Hr2zcXuh
wqLLwRADOgwc+mK5hrKx4hF/B2NHlg+fbV4tUtBHmUD8FiMWRnLQ3Fy+AKfivKAnLLuV4Yy+sfFN
r0Sknsc2bnSDmV+SjUt4w4uylGRWqubegfleKzQfR7LcuAB8uJ4zCnB55fwsuOjQAZQv/4LgCicH
lh0y/jHTvL+pzb2dd809S15+/bwz/lew+VnWTb9zw4X9RS/80yfbcvBh+Zs2yTNyx18HAaJG7FVf
XdVfeZ8u+VEJvz5kL1Kwhtc+SMH7oy+k5jq0EIvoggHmR7wQm6v0CfkFOcsa3p9uKUbfj7IRnL+X
rqIUbsy3Q/aCLE09WOcOfsBWX6tuNeML2p7v+icTNQdFFxgkVucJ53OG8dPvk8vIHfcv6I6iHPGb
dcb5UJFbOHlrPMSG3LKU8wvL1Na5X/Ug36OK9rs+u0OPS7X3rKIgDNmpcbADOucSYyNdXAgnKLq9
C/cfIuQ27bnTLqJD84yzGihaD/b32dIr74bB4xU2fqb9JJmhZjVxHLze8JIOhbwgBWzsyt14N/Ny
n+Jvl0M8TX6dL9BIfk9NokymhsOIqRLky2imJD69998+dTj9WYhq7weHi1uRjIgIZskbK+9ZI4dv
sDGun6u40ggIni9Coq72OdOdfcKXo2UxJGZcSnHxkEESCfcmB1KO/hbSGqyvRtR/G7sh5DSsoe8Z
17h3nvmAsV17+HealXJ2QNP3BKOdHcaIUQb5aCCU9qvtFv7hNwCUy394eKS5gzreNtuxKe3UYsfF
NIhJZOBebENMTLZj5sO9+v8KL7oy8TTofI15B+GIDvnUWxV8AJSvamxVLwXJqL07zDhRykfX8p6o
OeUCz7J/N4un0rXSHcZRHBAJPTtpdTZPeY4865cpb6OXRgfB2A+B7RFIM99TaqiRJLeyR82lscVz
mIt/873ypRfwx6WufFvC3yLSl1RlJGq3C1dYhtprexUIchJoasRC8cGBM3cDRiBmzk3TojebHJzL
S84qxWpjA/cr+ID2HSY5nQMBvyqj51/m16oqF5+GAfIM8nu5AJmqBytEHgLLmuE6dd3rP3asx00m
7Z4+0zHXUM9jWceiKkOz+PgN2PrhHro8rHNeMq0coJD4lZITS+0feN9vdPfPp3Wtcg7yhBDVJ0qM
erg6PzAdPYbLuOmHOMl1EQRuAGvn8RT6ibevdbgyXcppU354so27Hh6konnw+m1h0cgrOXUSY/zW
9l4hx9Jr24rnk/48a4f5jc6l44NsUB1aqipr3bH0bN7M5owOHaeqCIW7CLgRXOarFTZqRSFG8YJk
YeDfDZYQh9JP1aWhUzEkq5VoDXDpMD82iiU7l3UA+7uqabQl/DFLjCPGgby0Sd362lE+dLoaK3xd
3qdONu5yvwMMm6xvUY3UDFYrjD6B12x1zIIVSAb7ilxXzm8LuAm9aEsBk+GhU+ZQji3psSOAnocX
aIPlJB0j13h8NFAXpnIdAkhr5I+rC+paZUiblABx8ztBsfr6TwDy33jgE7nudOwXTH2PWT+9uxZ2
W6VzdwYboTYd5viN34gsljDc+sxia9Wcs+GDC4C7dyRyfwmkaB4AuZBK9iodefZ5XwbUv226NZTe
vUaf1tSwzvxobOJUF9d/qggwQo6N4wnLt1lTmNJJNUsQSPwuVPx72WQ4IRPeoIFykYipmmcR4j9n
KMmGUklBWblE2NSkA/FEQ/m7q5k5PeqqsUvRt56daPJuKlNzQQ1fS7hlSLLyvDcF0QiTS7fk3G0q
sNbzWsMVN3+qVBuVahdt5SCIoivaTKkJOyfeytN5nP75SFoTG+QVm2e4cAE+6T2FX8VmHN0riXKb
O5Or4s3fYQsr4O49T8lvLQAQQHzypGv0oh3rEuMLA+Va7htDJmyp7+5a3SvvIyo5lq3z5L055EOP
RaILFSZWVjIpkPNE5/4cUOKn4SZ6LOXUun6NUbV3bXgXEcFatMBmt0cxqD9Pi05474lKCUTD7Z5/
CByiRuF/7Vdbyfd2wcpdxikZBbwfNbaToLMBvIUesk0SXi1JRzdz3J5eTmL4LYrCGRGmLlue9p+D
MYr8q1aDocqs2bS0F3lufd3fUAq69GoWimZVXIXBPLew+niOJ8DVVpuFj6/7MEGcBfAhbVkKbe0+
1rvWybkKYB8XnjMkfAuaPRjMl/D+5y4IxANiPHX+Xt3gST3uCkVWcIAUOfPTqhQs0LuZ+6PLXAAa
MNmNQBHCHvWNEGnqKx3DpNCVMF/2sdEwbitkzxgIk9DDlcdoXlaBIxD7v11h/PGK6r4c8Mr29Fge
5xBz3RPTFFRAVJ0fYHg=
`pragma protect end_protected
