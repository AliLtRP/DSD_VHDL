// megafunction wizard: %ALTGX%
// GENERATION: STANDARD
// VERSION: WM1.0
// MODULE: alt4gxb 

// ============================================================
// File Name: rc_s4gxb_rx.v
// Megafunction Name(s):
// 			alt4gxb
//
// Simulation Library Files(s):
// 			
// ============================================================
// ************************************************************
// THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
//
// 10.1 Build 153 11/29/2010 SJ Full Version
// ************************************************************


//Copyright (C) 1991-2010 Altera Corporation
//Your use of Altera Corporation's design tools, logic functions 
//and other software and tools, and its AMPP partner logic 
//functions, and any output files from any of the foregoing 
//(including device programming or simulation files), and any 
//associated documentation or information are expressly subject 
//to the terms and conditions of the Altera Program License 
//Subscription Agreement, Altera MegaCore Function License 
//Agreement, or other applicable license agreement, including, 
//without limitation, that your use is for the sole purpose of 
//programming logic devices manufactured by Altera and sold by 
//Altera or its authorized distributors.  Please refer to the 
//applicable agreement for further details.


// synopsys translate_off
`timescale 1 ps / 1 ps
// synopsys translate_on
module rc_s4gxb_rx (
	cal_blk_clk,
	reconfig_clk,
	reconfig_togxb,
    gxb_powerdown,
	rx_analogreset,
	rx_bitslip,
	rx_cruclk,
	rx_datain,
	rx_digitalreset,
	rx_locktodata,
	rx_locktorefclk,
	reconfig_fromgxb,
	rx_clkout,
	rx_dataout,
	rx_pll_locked);

	input	  cal_blk_clk;
	input	  reconfig_clk;
	input	[3:0]  reconfig_togxb;
    input[0:0]  gxb_powerdown;
	input	[0:0]  rx_analogreset;
	input	[0:0]  rx_bitslip;
	input	[0:0]  rx_cruclk;
	input	[0:0]  rx_datain;
	input	[0:0]  rx_digitalreset;
	input	[0:0]  rx_locktodata;
	input	[0:0]  rx_locktorefclk;
	output	[16:0]  reconfig_fromgxb;
	output	[0:0]  rx_clkout;
	output	[19:0]  rx_dataout;
	output	[0:0]  rx_pll_locked;

	parameter	starting_channel_number = 4;
    parameter   rx_cru_inclock0_period = 6734;
    parameter   rx_data_rate = 1485;   
	parameter 	effective_data_rate = "1485 Mbps";  
	parameter 	input_clock_frequency = "148.50MHz"; 
 
	
	wire [0:0] sub_wire0;
	wire [0:0] sub_wire1;
	wire [19:0] sub_wire2;
	wire [0:0] sub_wire3 = 1'h0;
	wire [0:0] rx_pll_locked = sub_wire0[0:0];
	wire [0:0] rx_clkout = sub_wire1[0:0];
	wire [19:0] rx_dataout = sub_wire2[19:0];

	alt4gxb	alt4gxb_component (
				.rx_locktorefclk (rx_locktorefclk),
				.rx_revbitorderwa (sub_wire3),
				.rx_cruclk (rx_cruclk),
				.cal_blk_clk (cal_blk_clk),
				.reconfig_clk (reconfig_clk),
				.rx_locktodata (rx_locktodata),
				.rx_datain (rx_datain),
				.reconfig_togxb (reconfig_togxb),
                .gxb_powerdown (gxb_powerdown),
				.rx_bitslip (rx_bitslip),
				.rx_analogreset (rx_analogreset),
				.rx_digitalreset (rx_digitalreset),
				.reconfig_fromgxb (reconfig_fromgxb),
				.rx_pll_locked (sub_wire0),
				.rx_clkout (sub_wire1),
				.rx_dataout (sub_wire2)
				// synopsys translate_off
				,
				.aeq_fromgxb (),
				.aeq_togxb (),
				.cal_blk_calibrationstatus (),
				.cal_blk_powerdown (),
				.coreclkout (),
				.fixedclk (),
				.hip_tx_clkout (),
				.pipe8b10binvpolarity (),
				.pipedatavalid (),
				.pipeelecidle (),
				.pipephydonestatus (),
				.pipestatus (),
				.pll_inclk (),
				.pll_locked (),
				.pll_powerdown (),
				.powerdn (),
				.rateswitch (),
				.rateswitchbaseclock (),
				.reconfig_fromgxb_oe (),
				.rx_a1a2size (),
				.rx_a1a2sizeout (),
				.rx_a1detect (),
				.rx_a2detect (),
				.rx_bistdone (),
				.rx_bisterr (),
				.rx_byteorderalignstatus (),
				.rx_channelaligned (),
				.rx_coreclk (),
				.rx_ctrldetect (),
				.rx_dataoutfull (),
				.rx_disperr (),
				.rx_elecidleinfersel (),
				.rx_enabyteord (),
				.rx_enapatternalign (),
				.rx_errdetect (),
				.rx_freqlocked (),
				.rx_invpolarity (),
				.rx_k1detect (),
				.rx_k2detect (),
				.rx_patterndetect (),
				.rx_phase_comp_fifo_error (),
				.rx_phfifooverflow (),
				.rx_phfifordenable (),
				.rx_phfiforeset (),
				.rx_phfifounderflow (),
				.rx_phfifowrdisable (),
				.rx_pipebufferstat (),
				.rx_powerdown (),
				.rx_prbscidenable (),
				.rx_recovclkout (),
				.rx_revbyteorderwa (),
				.rx_rlv (),
				.rx_rmfifoalmostempty (),
				.rx_rmfifoalmostfull (),
				.rx_rmfifodatadeleted (),
				.rx_rmfifodatainserted (),
				.rx_rmfifoempty (),
				.rx_rmfifofull (),
				.rx_rmfifordena (),
				.rx_rmfiforeset (),
				.rx_rmfifowrena (),
				.rx_runningdisp (),
				.rx_seriallpbken (),
				.rx_signaldetect (),
				.rx_syncstatus (),
				.scanclk (),
				.scanin (),
				.scanmode (),
				.scanshift (),
				.testin (),
				.tx_clkout (),
				.tx_coreclk (),
				.tx_ctrlenable (),
				.tx_datain (),
				.tx_datainfull (),
				.tx_dataout (),
				.tx_detectrxloop (),
				.tx_digitalreset (),
				.tx_dispval (),
				.tx_forcedisp (),
				.tx_forcedispcompliance (),
				.tx_forceelecidle (),
				.tx_invpolarity (),
				.tx_phase_comp_fifo_error (),
				.tx_phfifooverflow (),
				.tx_phfiforeset (),
				.tx_phfifounderflow (),
				.tx_pipedeemph (),
				.tx_pipemargin (),
				.tx_pipeswing (),
				.tx_pllreset (),
				.tx_revparallellpbken ()
				// synopsys translate_on
				);
	defparam
		alt4gxb_component.input_clock_frequency = input_clock_frequency,
		alt4gxb_component.equalizer_ctrl_a_setting = 0,
		alt4gxb_component.equalizer_ctrl_b_setting = 0,
		alt4gxb_component.equalizer_ctrl_c_setting = 0,
		alt4gxb_component.equalizer_ctrl_d_setting = 0,
		alt4gxb_component.equalizer_ctrl_v_setting = 0,
		alt4gxb_component.equalizer_dcgain_setting = 0,
		alt4gxb_component.intended_device_family = "Stratix IV",
		alt4gxb_component.loopback_mode = "none",
		alt4gxb_component.lpm_hint = "CBX_HDL_LANGUAGE=Verilog",
		alt4gxb_component.lpm_type = "alt4gxb",
		alt4gxb_component.number_of_channels = 1,
		alt4gxb_component.operation_mode = "rx",
		alt4gxb_component.protocol = "basic",
		alt4gxb_component.receiver_termination = "oct_100_ohms",
		alt4gxb_component.reconfig_dprio_mode = 2,
		alt4gxb_component.rx_8b_10b_compatibility_mode = "true",
		alt4gxb_component.rx_8b_10b_mode = "none",
		alt4gxb_component.rx_align_pattern = "0101111100",
		alt4gxb_component.rx_align_pattern_length = 10,
		alt4gxb_component.rx_allow_align_polarity_inversion = "false",
		alt4gxb_component.rx_allow_pipe_polarity_inversion = "false",
		alt4gxb_component.rx_bitslip_enable = "true",
		alt4gxb_component.rx_byte_ordering_mode = "NONE",
		alt4gxb_component.rx_channel_width = 20,
		alt4gxb_component.rx_common_mode = "0.82v",
		alt4gxb_component.rx_cru_bandwidth_type = "Medium",
		alt4gxb_component.rx_cru_inclock0_period = rx_cru_inclock0_period,
		alt4gxb_component.rx_datapath_low_latency_mode = "false",
		alt4gxb_component.rx_datapath_protocol = "basic",
		alt4gxb_component.rx_data_rate = rx_data_rate,
		alt4gxb_component.effective_data_rate = effective_data_rate,
		alt4gxb_component.rx_data_rate_remainder = 0,
		alt4gxb_component.rx_digitalreset_port_width = 1,
		alt4gxb_component.rx_disable_auto_idle_insertion = "false",
		alt4gxb_component.rx_enable_bit_reversal = "false",
		alt4gxb_component.rx_enable_deep_align_byte_swap = "false",
		alt4gxb_component.rx_enable_lock_to_data_sig = "true",
		alt4gxb_component.rx_enable_lock_to_refclk_sig = "true",
		alt4gxb_component.rx_enable_true_complement_match_in_word_align = "false",
		alt4gxb_component.rx_flip_rx_out = "false",
		alt4gxb_component.rx_force_signal_detect = "true",
		alt4gxb_component.rx_ppmselect = 32,
		alt4gxb_component.rx_rate_match_fifo_mode = "none",
		alt4gxb_component.rx_run_length = 40,
		alt4gxb_component.rx_run_length_enable = "true",
		alt4gxb_component.rx_signal_detect_threshold = 2,
		alt4gxb_component.rx_use_align_state_machine = "false",
		alt4gxb_component.rx_use_clkout = "true",
		alt4gxb_component.rx_use_coreclk = "false",
		alt4gxb_component.rx_use_cruclk = "true",
		alt4gxb_component.rx_use_deserializer_double_data_mode = "false",
		alt4gxb_component.rx_use_deskew_fifo = "false",
		alt4gxb_component.rx_use_double_data_mode = "true",
		alt4gxb_component.use_calibration_block = "true",
		alt4gxb_component.gxb_analog_power = "AUTO",
		alt4gxb_component.gxb_powerdown_width = 1,
		alt4gxb_component.number_of_quads = 1,
		alt4gxb_component.rx_cru_data_rate = 673,
		alt4gxb_component.rx_cru_divide_by = 1,
		alt4gxb_component.rx_cru_m_divider = 0,
		alt4gxb_component.rx_cru_multiply_by = 10,
		alt4gxb_component.rx_cru_n_divider = 1,
		alt4gxb_component.rx_cru_pfd_clk_select = 0,
		alt4gxb_component.rx_cru_vco_post_scale_divider = 2,
		alt4gxb_component.rx_dwidth_factor = 2,
		alt4gxb_component.rx_reconfig_clk_scheme = "indv_clk_source",
		alt4gxb_component.rx_word_aligner_num_byte = 1,
		alt4gxb_component.reconfig_calibration = "true", 
		alt4gxb_component.reconfig_fromgxb_port_width = 17, 
		alt4gxb_component.reconfig_togxb_port_width = 4,
		alt4gxb_component.starting_channel_number = starting_channel_number;


endmodule

// ============================================================
// CNX file retrieval info
// ============================================================
// Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Stratix IV"
// Retrieval info: PRIVATE: NUM_KEYS NUMERIC "70"
// Retrieval info: PRIVATE: RECONFIG_PROTOCOL STRING "Basic"
// Retrieval info: PRIVATE: RECONFIG_SUBPROTOCOL STRING "none"
// Retrieval info: PRIVATE: RX_ENABLE_DC_COUPLING STRING "false"
// Retrieval info: PRIVATE: SYNTH_WRAPPER_GEN_POSTFIX STRING "0"
// Retrieval info: PRIVATE: WIZ_BASE_DATA_RATE STRING "2970.00"
// Retrieval info: PRIVATE: WIZ_BASE_DATA_RATE_ENABLE STRING "0"
// Retrieval info: PRIVATE: WIZ_DATA_RATE STRING "2970"
// Retrieval info: PRIVATE: WIZ_DPRIO_INCLK_FREQ_ARRAY STRING "312.500000 250.000000 156.250000 125.000000 312.500000 250.000000 156.250000 125.000000"
// Retrieval info: PRIVATE: WIZ_DPRIO_INPUT_A STRING "2500"
// Retrieval info: PRIVATE: WIZ_DPRIO_INPUT_A_UNIT STRING "Mbps"
// Retrieval info: PRIVATE: WIZ_DPRIO_INPUT_B STRING "312.500000"
// Retrieval info: PRIVATE: WIZ_DPRIO_INPUT_B_UNIT STRING "MHz"
// Retrieval info: PRIVATE: WIZ_DPRIO_INPUT_SELECTION NUMERIC "0"
// Retrieval info: PRIVATE: WIZ_DPRIO_REF_CLK0_FREQ STRING "371.25"
// Retrieval info: PRIVATE: WIZ_DPRIO_REF_CLK0_PROTOCOL STRING "Basic"
// Retrieval info: PRIVATE: WIZ_DPRIO_REF_CLK1_FREQ STRING "250"
// Retrieval info: PRIVATE: WIZ_DPRIO_REF_CLK1_PROTOCOL STRING "Basic"
// Retrieval info: PRIVATE: WIZ_DPRIO_REF_CLK2_FREQ STRING "250"
// Retrieval info: PRIVATE: WIZ_DPRIO_REF_CLK2_PROTOCOL STRING "Basic"
// Retrieval info: PRIVATE: WIZ_DPRIO_REF_CLK3_FREQ STRING "250"
// Retrieval info: PRIVATE: WIZ_DPRIO_REF_CLK3_PROTOCOL STRING "Basic"
// Retrieval info: PRIVATE: WIZ_DPRIO_REF_CLK4_FREQ STRING "250"
// Retrieval info: PRIVATE: WIZ_DPRIO_REF_CLK4_PROTOCOL STRING "Basic"
// Retrieval info: PRIVATE: WIZ_DPRIO_REF_CLK5_FREQ STRING "250"
// Retrieval info: PRIVATE: WIZ_DPRIO_REF_CLK5_PROTOCOL STRING "Basic"
// Retrieval info: PRIVATE: WIZ_DPRIO_REF_CLK6_FREQ STRING "250"
// Retrieval info: PRIVATE: WIZ_DPRIO_REF_CLK6_PROTOCOL STRING "Basic"
// Retrieval info: PRIVATE: WIZ_ENABLE_EQUALIZER_CTRL NUMERIC "0"
// Retrieval info: PRIVATE: WIZ_EQUALIZER_CTRL_SETTING NUMERIC "0"
// Retrieval info: PRIVATE: WIZ_FORCE_DEFAULT_SETTINGS NUMERIC "0"
// Retrieval info: PRIVATE: WIZ_INCLK_FREQ STRING "148.50"
// Retrieval info: PRIVATE: WIZ_INCLK_FREQ_ARRAY STRING "59.40 74.25 92.81 118.80 148.50 185.625 237.60 297.00 371.25 475.20 594.00"
// Retrieval info: PRIVATE: WIZ_INPUT_A STRING "2970"
// Retrieval info: PRIVATE: WIZ_INPUT_A_UNIT STRING "Mbps"
// Retrieval info: PRIVATE: WIZ_INPUT_B STRING "148.50"
// Retrieval info: PRIVATE: WIZ_INPUT_B_UNIT STRING "MHz"
// Retrieval info: PRIVATE: WIZ_INPUT_SELECTION NUMERIC "0"
// Retrieval info: PRIVATE: WIZ_PROTOCOL STRING "Basic"
// Retrieval info: PRIVATE: WIZ_RX_VCM STRING "0.82"
// Retrieval info: PRIVATE: WIZ_SUBPROTOCOL STRING "None"
// Retrieval info: PRIVATE: WIZ_TX_VCM STRING "0.6"
// Retrieval info: PRIVATE: WIZ_VCCHTX STRING "1.4"
// Retrieval info: PRIVATE: WIZ_WORD_ALIGN_FLIP_PATTERN STRING "0"
// Retrieval info: PRIVATE: wiz_speed_grade STRING "2"
// Retrieval info: CONSTANT: EQUALIZER_CTRL_A_SETTING NUMERIC "0"
// Retrieval info: CONSTANT: EQUALIZER_CTRL_B_SETTING NUMERIC "0"
// Retrieval info: CONSTANT: EQUALIZER_CTRL_C_SETTING NUMERIC "0"
// Retrieval info: CONSTANT: EQUALIZER_CTRL_D_SETTING NUMERIC "0"
// Retrieval info: CONSTANT: EQUALIZER_CTRL_V_SETTING NUMERIC "0"
// Retrieval info: CONSTANT: EQUALIZER_DCGAIN_SETTING NUMERIC "0"
// Retrieval info: CONSTANT: INTENDED_DEVICE_FAMILY STRING "Stratix IV"
// Retrieval info: CONSTANT: LOOPBACK_MODE STRING "none"
// Retrieval info: CONSTANT: LPM_TYPE STRING "alt4gxb"
// Retrieval info: CONSTANT: NUMBER_OF_CHANNELS NUMERIC "1"
// Retrieval info: CONSTANT: OPERATION_MODE STRING "rx"
// Retrieval info: CONSTANT: PROTOCOL STRING "basic"
// Retrieval info: CONSTANT: RECEIVER_TERMINATION STRING "oct_100_ohms"
// Retrieval info: CONSTANT: RECONFIG_DPRIO_MODE NUMERIC "0"
// Retrieval info: CONSTANT: RX_8B_10B_COMPATIBILITY_MODE STRING "true"
// Retrieval info: CONSTANT: RX_8B_10B_MODE STRING "none"
// Retrieval info: CONSTANT: RX_ALIGN_PATTERN STRING "0101111100"
// Retrieval info: CONSTANT: RX_ALIGN_PATTERN_LENGTH NUMERIC "10"
// Retrieval info: CONSTANT: RX_ALLOW_ALIGN_POLARITY_INVERSION STRING "false"
// Retrieval info: CONSTANT: RX_ALLOW_PIPE_POLARITY_INVERSION STRING "false"
// Retrieval info: CONSTANT: RX_BITSLIP_ENABLE STRING "true"
// Retrieval info: CONSTANT: RX_BYTE_ORDERING_MODE STRING "NONE"
// Retrieval info: CONSTANT: RX_CHANNEL_WIDTH NUMERIC "20"
// Retrieval info: CONSTANT: RX_COMMON_MODE STRING "0.82v"
// Retrieval info: CONSTANT: RX_CRU_BANDWIDTH_TYPE STRING "Medium"
// Retrieval info: CONSTANT: RX_CRU_INCLOCK0_PERIOD NUMERIC "6734"
// Retrieval info: CONSTANT: RX_DATAPATH_LOW_LATENCY_MODE STRING "false"
// Retrieval info: CONSTANT: RX_DATAPATH_PROTOCOL STRING "basic"
// Retrieval info: CONSTANT: RX_DATA_RATE NUMERIC "2970"
// Retrieval info: CONSTANT: EFFECTIVE_DATA_RATE NUMERIC "2970 Mbps"
// Retrieval info: CONSTANT: RX_DATA_RATE_REMAINDER NUMERIC "0"
// Retrieval info: CONSTANT: RX_DIGITALRESET_PORT_WIDTH NUMERIC "1"
// Retrieval info: CONSTANT: RX_DISABLE_AUTO_IDLE_INSERTION STRING "false"
// Retrieval info: CONSTANT: RX_ENABLE_BIT_REVERSAL STRING "false"
// Retrieval info: CONSTANT: RX_ENABLE_DEEP_ALIGN_BYTE_SWAP STRING "false"
// Retrieval info: CONSTANT: RX_ENABLE_LOCK_TO_DATA_SIG STRING "true"
// Retrieval info: CONSTANT: RX_ENABLE_LOCK_TO_REFCLK_SIG STRING "true"
// Retrieval info: CONSTANT: RX_ENABLE_TRUE_COMPLEMENT_MATCH_IN_WORD_ALIGN STRING "false"
// Retrieval info: CONSTANT: RX_FLIP_RX_OUT STRING "false"
// Retrieval info: CONSTANT: RX_FORCE_SIGNAL_DETECT STRING "true"
// Retrieval info: CONSTANT: RX_PPMSELECT NUMERIC "32"
// Retrieval info: CONSTANT: RX_RATE_MATCH_FIFO_MODE STRING "none"
// Retrieval info: CONSTANT: RX_RUN_LENGTH NUMERIC "40"
// Retrieval info: CONSTANT: RX_RUN_LENGTH_ENABLE STRING "true"
// Retrieval info: CONSTANT: RX_SIGNAL_DETECT_THRESHOLD NUMERIC "2"
// Retrieval info: CONSTANT: RX_USE_ALIGN_STATE_MACHINE STRING "false"
// Retrieval info: CONSTANT: RX_USE_CLKOUT STRING "true"
// Retrieval info: CONSTANT: RX_USE_CORECLK STRING "false"
// Retrieval info: CONSTANT: RX_USE_CRUCLK STRING "true"
// Retrieval info: CONSTANT: RX_USE_DESERIALIZER_DOUBLE_DATA_MODE STRING "false"
// Retrieval info: CONSTANT: RX_USE_DESKEW_FIFO STRING "false"
// Retrieval info: CONSTANT: RX_USE_DOUBLE_DATA_MODE STRING "true"
// Retrieval info: CONSTANT: USE_CALIBRATION_BLOCK STRING "true"
// Retrieval info: CONSTANT: gxb_analog_power STRING "AUTO"
// Retrieval info: CONSTANT: gxb_powerdown_width NUMERIC "1"
// Retrieval info: CONSTANT: number_of_quads NUMERIC "1"
// Retrieval info: CONSTANT: rx_cru_data_rate NUMERIC "673"
// Retrieval info: CONSTANT: rx_cru_divide_by NUMERIC "1"
// Retrieval info: CONSTANT: rx_cru_m_divider NUMERIC "10"
// Retrieval info: CONSTANT: rx_cru_multiply_by NUMERIC "10"
// Retrieval info: CONSTANT: rx_cru_n_divider NUMERIC "1"
// Retrieval info: CONSTANT: rx_cru_pfd_clk_select NUMERIC "0"
// Retrieval info: CONSTANT: rx_cru_vco_post_scale_divider NUMERIC "2"
// Retrieval info: CONSTANT: rx_dwidth_factor NUMERIC "2"
// Retrieval info: CONSTANT: rx_word_aligner_num_byte NUMERIC "1"
// Retrieval info: CONSTANT: reconfig_calibration STRING "true"
// Retrieval info: CONSTANT: reconfig_fromgxb_port_width NUMERIC "17"
// Retrieval info: CONSTANT: reconfig_togxb_port_width NUMERIC "4"
// Retrieval info: USED_PORT: cal_blk_clk 0 0 0 0 INPUT NODEFVAL "cal_blk_clk"
// Retrieval info: USED_PORT: rx_analogreset 0 0 1 0 INPUT NODEFVAL "rx_analogreset[0..0]"
// Retrieval info: USED_PORT: rx_bitslip 0 0 1 0 INPUT NODEFVAL "rx_bitslip[0..0]"
// Retrieval info: USED_PORT: rx_clkout 0 0 1 0 OUTPUT NODEFVAL "rx_clkout[0..0]"
// Retrieval info: USED_PORT: rx_cruclk 0 0 1 0 INPUT GND "rx_cruclk[0..0]"
// Retrieval info: USED_PORT: rx_datain 0 0 1 0 INPUT NODEFVAL "rx_datain[0..0]"
// Retrieval info: USED_PORT: rx_dataout 0 0 20 0 OUTPUT NODEFVAL "rx_dataout[19..0]"
// Retrieval info: USED_PORT: rx_digitalreset 0 0 1 0 INPUT NODEFVAL "rx_digitalreset[0..0]"
// Retrieval info: USED_PORT: rx_locktodata 0 0 1 0 INPUT NODEFVAL "rx_locktodata[0..0]"
// Retrieval info: USED_PORT: rx_locktorefclk 0 0 1 0 INPUT NODEFVAL "rx_locktorefclk[0..0]"
// Retrieval info: USED_PORT: rx_pll_locked 0 0 1 0 OUTPUT NODEFVAL "rx_pll_locked[0..0]"
// Retrieval info: CONNECT: @rx_locktorefclk 0 0 1 0 rx_locktorefclk 0 0 1 0
// Retrieval info: CONNECT: @rx_analogreset 0 0 1 0 rx_analogreset 0 0 1 0
// Retrieval info: CONNECT: rx_dataout 0 0 20 0 @rx_dataout 0 0 20 0
// Retrieval info: CONNECT: @cal_blk_clk 0 0 0 0 cal_blk_clk 0 0 0 0
// Retrieval info: CONNECT: rx_pll_locked 0 0 1 0 @rx_pll_locked 0 0 1 0
// Retrieval info: CONNECT: @rx_revbitorderwa 0 0 1 0 GND 0 0 1 0
// Retrieval info: CONNECT: rx_clkout 0 0 1 0 @rx_clkout 0 0 1 0
// Retrieval info: CONNECT: @rx_digitalreset 0 0 1 0 rx_digitalreset 0 0 1 0
// Retrieval info: CONNECT: @rx_cruclk 0 0 1 0 rx_cruclk 0 0 1 0
// Retrieval info: CONNECT: @rx_bitslip 0 0 1 0 rx_bitslip 0 0 1 0
// Retrieval info: CONNECT: @rx_locktodata 0 0 1 0 rx_locktodata 0 0 1 0
// Retrieval info: CONNECT: @rx_datain 0 0 1 0 rx_datain 0 0 1 0
// Retrieval info: GEN_FILE: TYPE_NORMAL rc_gxb_rx.v TRUE FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL rc_gxb_rx.inc FALSE FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL rc_gxb_rx.cmp FALSE FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL rc_gxb_rx.bsf FALSE FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL rc_gxb_rx_inst.v FALSE FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL rc_gxb_rx_bb.v FALSE FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL rc_s4gxb_rx.v TRUE FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL rc_s4gxb_rx.ppf TRUE FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL rc_s4gxb_rx.inc FALSE FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL rc_s4gxb_rx.cmp FALSE FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL rc_s4gxb_rx.bsf FALSE FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL rc_s4gxb_rx_inst.v FALSE FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL rc_s4gxb_rx_bb.v TRUE FALSE
// Retrieval info: LIB_FILE: stratixiv_hssi
