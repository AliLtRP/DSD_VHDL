// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:54 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
lClDhPnZ8IloBEqpR4SbEKQJ4v/4NF+la029a29saYOzQl5QbbWbD5q15FAA6SwG
G+PQr0qqI7Qd5PO81zR/E7nag/ifCAJOVWkNv65Y8bJgnKI62gZCCBh7NhUUwAwv
+pOFE+CYf8WpA8jTg2MU5Uzne62yHLFAkaGcJ1zNqY4=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 19424)
xzzjutQzF/mpvFZPgUqtNu0ya9TLcwKSGLcK6Llhv0po3chY6juyXEG0pU1FFo75
8q3pY3slEHgp0XVmB6aWye+3El/JOmMKOmJm9D0P02eB9MsugzofToeVypOtlSpQ
5uD6sCdL3V/eeAs8Adrdce/3X3klb6jLrSyvr2GLHrf1d+E1Q9lo/wJRntvCTI8O
++1p/F1ywYOqU+qN8B/Q6xiUJ+ZbWh7fe+5ImY7/4DfvAed9KZrz4FpftePNO8Ht
Hip+1pQJB77v6Cbv1SqB7l7sJUccQv09WxyOnnU5f6hyMUC1jK590Z/D1S9S5Mpo
c8eiD1Iq1BQsA/g7UV/sF3X61tyfO9/fTzhnGFinNvM+L3RBcAMAaOIXUNHRMKVU
ux2Wt4eAKl9lDzemXlYsntvIHIIIMkUJJ/wx6AQtCgOk0k4ac8uiff+DeD8Wzt6T
e7Z3iildKJ4BhOpxdvP6nZ4SL9nv8RaNbWj9je8Fqz2b+sckS0rH+wHrwzT9Gcvs
TUVOKB5i6IxJHyS54+uGzqySFvZ31VJyveg+oeo3mDbtmbXefrvPEGtDMnnTDXf4
EUW9b/2tiA8dLs6SQu2dw3ZioEVivc7p975rMfc22I7OK5ytVh/MY++rnB/Azz1U
KpZ/neIvStDJt6HSlsDCZRfM1+0/JFINN0BTsO/s+1+284PsvxaU68Gu5yO2kDE8
W2M/l9UbicJqVmgw6Od3hts6bmt9AQ7Ks8Px298RYSnP60s/RPPrpnszkC0mgiSG
+rf56amD4P+IW3yvlMzUb+nBVeiF8asMcQQVnutFuw//wCreoNaGzVL/bNoASKME
bZhPeRj/TotUWPj9W7hPqR95NxF48h8R8cWUUbZHE6K832knRyVt4VJ8dku+/VYE
L7zCytGEL3/B3gIxzzLSeO6qWR8YRT4rvXXTfpzukKSsGJGD7q1rfRoy/aMRo8cf
G4v+nO8iR29wOS9bpMJDzhFW+CVYusQWd+h5inLIawc+/Dcccx6aKUzO8x4VV4Wr
35GvsqwDmIMkoC308kB30nnjkTMjGvSpwuLeP9td3uiNp+DqrBKBvl6oJVI586ut
iJv747XydQZoEFton2XdOaQBwuv4Deju9uh/M/kXAeKoG2bdA00hZ4lYYlSKoXvf
bm6Mh/KjmkQJ3miU+7wzTV+sIm2zcYUeFvnA6Vmb96lbwIwbvQgoPFEEhIJwo42R
qdw5nMqyPNoKj9b2bTc+tHCynO+dcOEee9Fu48ktZlebCWwRDShyzLoNOgEKbp5a
VCS8HxYYweetB+Lh4vqackPpZ1KP7saIup66RJb0llx9HdATnUJ2vB5NIj9hM9JY
+5+MBPxd05EYLZ9LWVj0efkm2BWI5KUCTemxjL4HkqoJmQwl23E6NKZHvZjQ7T5N
GRt+zxVIg5CejX/dkPB/dXbXTbAL2zxfIWi4tbKDVsGo0oYyCD27y/2Jf1BfhJwV
ciQ3YY0lsQMdw5LA+IJ3mRffDtZUXD1XbznCPtgY8/pTzLQsHONNgrMUGmSzI23Z
2W/n1lFOtz8mX0ZPCJltzeAdUYgxXO4F4Ghc6Hzl5tEBDkNA7VsW4FlH/I2ph8vn
vOpvrn52AwrXuXLuoH6YPQbezBhwYJ6RNa5yr5GHl+twl+LeLn3dsiVnBP7o6mRF
8x9i2EDkrnia3cnO/898y+sXMx5+eQkDwR8qiB2yNLlMWKSJqr+XIdhZOUgYnWD6
MHBTRsEBbN9hF5FOI8fQOlb8CKdHjT64d532PfvtiPprS3aXFV7fYWf0GR4m64jE
2YdayHdnTwYLr32gpdpIOVfOfIihMUdpF8fnem+JrYJ5LVxx2MkiW1QGwMXxQmce
BTYvju72+h34exNFtbFnlBsrEOf+2qMPkt3uPtdSifcZn8L+13Rhnk5hjw93kbHu
Tt8fdukCv4X/oJC+/Du0pb7p3st8kFbEfqzJEqPW+4P6t9PX1NL6wTepsT5Zlb/6
gBM400vlNhKGpmrYxXpK/F1LdKE8yOKr3wShLxgi2UmpTF+k/zNtvqBCjqboKH7R
5eEZGOuQ+OG23TzgYXMTCs9236CfM18/m4tVPhKAf5xNfZMCJzuBh2l6SIq7fLdL
PU08Xu6Po1e0Ny0labElc+H9KgaY2vyBNN6mlj+UzRIj18efxpUDp2BNSSST1w4r
M5QtDixUMFZtW09T3gl2aUJVSViLtK1Td09o14yjx52Pwuf4spoQwgs68uydtmWr
r0CKUyKTdh5y96/+nPO4G/+VajxsGEmrQkOTmu3+x5n35is5+FJ8ZcyKvJAvdXZB
DSmFRsHr+HcKcByrkIYEKgG3ED6oY1qllpjc/j/pVfIEVTRCWhqPltdFDJXWAeLZ
zx8AiXJ92UgPCxOWNvbrwdq36RlBSqcUiKGEQWlQ7HdkQ57E3x8JIbiG97oKXcvt
KB6hsQKxcniTdcYIJyJz4Oravr1h7JMOzb/JlA5fOPZK5zgX49NNwbAJBDEakaun
rIyURv35JMZJRrQQCJnnT16h4Vk0S0YS76WVLiprYmtfAaFaPU5HDnWLpe+xyOdU
kbni7FVaCKsjQ+Yal/RT7whYSorISmYZ10ES9pr9iHuvb9Qaj6TrU+i5Dbr+Clem
4FYk8SV6apFSODMDUgmONhAv9tK9D5akDpF4ZWUVRACcJZHxMynE7n7HSEpVzyqy
v3rZBj6BKgu9jW1f8yhEPlsUoAwT2IxW0ldlZIXsHtKTfNufahuEFF9PvvnNg7J0
4o1uSDP3YoU8OTaxQAtxjHR17FyVMqupl4SFEkR5qjvNWkYt/t0zgVZFLiE8XnDo
zacEVrEyyNIZUNZXKnuh3ijxvha8xvGdmZZAWcSKBxExriRfqu6Yh1xjH8qDVFYw
JsspzEw7yM70EXzVkhhbeXFx9rTBFWYLOLuRhI3SA12fZdzaS6MHeQWq6rHnzOwh
ZuWeTuDzz0d+8Tbwq1ZDDIa1dtxr+rBaoACvUfsBj6oDMnkGAZpBCAje84wAW4Ci
hv7bal9FEG4T9NcHLhy0TtIFMmTkMi/vZeTnlYwIBZUdytHjC8gxbDslwJxBf0rW
PCxpoH9aq4v0T93BymW2/jJYmQZsRDQpwZvUfRTwnzZW7iJ5YyIssPpGuLuOWNgZ
reHyg4ftEE391znxRMMdvIgn90TPnBUEX9pGeHD1q5Jk4yTEt8CHsnh30Oj2rw4v
TpCaw/Vy9R0NGYs+D5wrBktoE1F8oXzZd5IVueGobijphVSI1TyY8h6pD5KA/+e1
xkfFl2B9qv9dpEFeWe11Fm2FxkFaqcEZVRIFySrSO5GH1DvJ5ho653+fHVzicg1P
UEOlvnEprDcBIqpqGwv7NfYG/ePyUB1zgJtcVE3r0lWinCxONohfM34gW1+mRmce
iNWm/CeuIeM+5J9piwCkhucp2vfu1/KyeJbiqqm/jJTckxUUw6AG/cs8y7Hm7N79
RM3rQ1LRscvWjyJ0Wd/9GH9e5uv8XM0NPA6J7LfpIlQo8+3cTzL1KvmqC9K8I6AH
vSBc7JLwIUrxsgsUMaK51GzA5UqvFbj9E4nVe10WeqjbLiZqK7DAiJ49+n2copMc
z5IQw+K1baw1PTy6zRDNEzV70Uth3KmOEzYmqy6GmdX6O/1+AHUJKrUQaKXjycn7
vqkqOicL26vdUbY1ZZe/ojYy+4iSQi5U9TcV9kRFV/VvzzQqfNm+6QLg/xWyTM5S
VNSQ4kgZRyhpmZBcRNSbuwkTvkBkUN7pTcyvoBPvzUzcXwTbAmpUwfGffAyDkSiE
f5VrTI8k++TxdvJFk6VuojNYSLZ0Dzmftfv1RQJbt+mLzcKdMsuXjQsND0Uqrmr1
AcDGjULAM8BobYQWiapOM63y1VRMRw/8uV0oniR7omc6u3bPc+5f17qmCnFzAINF
fohA6GUWKogkafr2KhD/ARDDD5HMZ4VAq4mv3wOxFaRdZ1bkzC502p+jqQbjKKQ6
2G1IoJNtA3I2+dimXtxnyk0Kh3wh9m2x+xetbR08U16ncU/Yk0Hd/7Da1f6f9nbg
33zax/NDu9fLPNhG3+E9v/DGOPzNCR2ZOI8asJjtCslabksbkADPYhpWNrGLKN7S
FvNzKtOh30XaCCZKy7d2SN6BdGAlYtxkDmz3oLkfS1L0QXfI6GR5ZQZzoPpArWp8
2b6qJHgRcb3/IbeNpzbHbfwgwrOKcjsDbRmGpGkMJbhPQiXEnQ5lXfom0n6C/R+t
J+8riGAfIBOvYIFYZe7HYKKUwyKylWde4kbaxJGjRuc9LWV7y0NLUDI2ZDri0IWw
6SOocn7ZLf0czWxa1/imxiXKb6LZWUCARhPKP4T1sVpTqVwz61Ee9sp39xN1FRdz
xVA/Epi+8KPA56zi9j00+eCun+4uj3hI2TXjxdOlJU/otbZnFiOLG2KEzcjy9ACu
DX3Oj34RoT4vMXVymiLryDAwSP5MO4ZDu+b33eia1auYPN2ZQnUYPJNSPaPrBEDF
GkK8ideXdjV4NOHgaC4qDbP0tzb3hF9e1Em1MmL5Ly4Y2vKVLdFcU/KkvFW4DZjg
4jnUf1ia1gyoVr7MEgp11diczy8lQmWCQO4HzKZKYGbvR1RyApPovj4Xw8GVJSra
CROLpn4/K9D6qKEeW16doZD5eeNWy2uqCS5s5QdI1oK76rU5/Fo2oQoZF2TQ/HPw
Y/PSfZKLr6vuaME1orDUVdOYylkaeZKC8m+1z6XyC9FeZd0Mq1S+74IrNvYznnXC
ePJdsgFe1A3oMc5IAez6nxkhp/H6keucqn/i4HFw/tutBuXxx0XwVJwUzgFXiOUu
Nt2HJKhQSowrJZTTSKinw/a7kkFi9JqGd3yOGznUdENzfi3BA8tQqRH5ahJe5eEl
ocDaZsY0GdA3UmiufBAfiXBSPR4F3LoPRJmcjPUZZ8bIw490781nGeXfeGmyv2yr
Za1K00MhAL09Pah/hvvcN7ueSKt6jWrGCtd8k2oOBX/yuG4GTLe/r1S9mHnqDOq5
tuM1Xu3Q3b33D/zL8VE4lfC/XYcWCJK+1BOZp124X1pyfWnhSwHuynAMwrfFA189
9ckmMb/UIIIagAWsy8tZ7E7ndldfuEuHbxAr229pWQmpXfhkjkwVxuAINjD+d+7j
tOmCTm22XCfUmHNbQgJ2JshGqbajBe4ABfSUWuATFF1WtYOfR2L344kfaqw5LGZX
+qoLPqMilOlRK31QaKz0a4CZDAFaTqCmOo2TU3VtPISvMx2A/H915t5QxLo2xx+L
cxbc43O+zknfJ6kItdwnoeuMTEbKjVoso78qAKMZu6nRxnDA4zzCjqEFQaW4L/s6
pnBDyLqvIqBxlqB4OEHrrMXEAjEZdhG3h8uuKBFtDEs60sCTcsxopuRGRUZX+bbX
HyRC65VvBpBh5CwRsFvYYpywZt+liDJv3aUuUbzVOBYtVkAHnSlFa4/728CrF7xs
9SoFzaSG/ffAprwrslk4KjHLfhxNc6MXC3VRgt3qiz0aF6v3qOcvxBVkQL+OYKwS
tZoybJKGGpiGSlI5rFiniaaKYnZ1Jdx5ter7uNi9UdU18c1NwvrO56MVi0leUaB4
nZRpdoCJ8Rqve7Gq1blMDB+g/DUSLHrsaE4Zwh7f75vvbwarJ/lc669i6cY7Cavj
Xh/xho/zC8vuGdTdhyCwor15aeJGKOqAfK1dA7QCTWfd02lnx24ZQ/M2P8simpeb
0xq9puor72wB9MWe3qSPWohyaowNQfbn/zrwJbvQ1MuFBDt+dv2lzIiPHqT5Pri0
PRbsZxuabceJyohT+0/18D11TSAUgC2WmtN6XT0Fb5nRDGrUenxYRBsKA8Xyu4WV
2mx3YGYOfZbnvEcvhmDNd8KUcq/Liixtcb51bkYNWQ/IrnaeU5OWBGhxrIR6C1PI
aReIYBlo3YOx3CCtjxcKjqbF1geaBu3SuE28DvQOGNRwdVIJGgKHNM8ordeSRWI3
U+UN67ilWsNIaAyFUpmf5vrqMDpK7TAKoq8WTFZ+GbAgWm3sKRqniHFg/NOHrw7U
m7/3minPDivmoBTUZFUzyLLrnzM9Zis5Uy99BuLna6JjeomSKL3kVdZegZ5Nd0Kl
TQU+7ZoGqxtt3vrtQU9IMMqRdEkUVCNn7eLlZbzeu3dqV/wpR+7viwz8yNXH6rri
mZzfD22I59W6eA5INe7OCTYfjQ5wxjgkso+1opDRXyIkB2Wt4BiuGS145FqRBseo
lS1QRNhA+ZbnhNoE6KqOn1RiU16LerD1+36guEkJfVBpR+eCVMMqLacS4GbTSngN
RXT9Fr2dPV3tLc0bnAyqj9lhlgEfCy55ba6i2NB9OiCTq4BROR1dvq8LKPUsiMh8
FsDKM7WnJuJQg/pTN6Omcwjjj/gcD1+FmGenvd5Pe1pdhBvKCcV3VTSuf0gD++sN
9FOVoZzMtZop/JnCaO+hROWL2Y3iJN79/3yUn8wj/uABsKswJIyimI7L4sJcxc7B
MW2coRiw6DQAZ7xibezLT59VXGktaQJ1spf2smsW/Em8jIQOIP82j9q1djiOoHTC
nKR4rieZOOVCXrcHuw1TbmBqmJkVkKfGCainoV/Pgz3N5G2qIzttn/iTJ3cSpHix
k2uFzxvlcIHIEVR1j9nhmoW59Ni+7aJobC8USu/egP9PbmdqGo6d1ANQirAkggN/
Ax+qJ2JdWUwc0fJ2s90B5VgTbDQCwrBCemK/j8Ag/Khc/1VIkqwXg+ETBNO05EzH
fzJMiQg32WBOQQ66l67f7XYq2E/EzsMbaYR7mm3OIQtRXOhV/tiU08pBf9bg8fH/
rHCkIjTw/YqKh2I1lqkqVWfAA/sZQ6+8kMdrPQVqEoCMJ2ilpB6qKM4huxSKMv9d
GWrtYu7zSRdId8BTGk7JUH8wwZl0TsNVwn4C+B/zwiwUGr+6N8f66Imxj5cxAuYK
+N4RvLlUSdT+BN1HyyaNNwIZKTLUsxwhiY6GHpnBa4cqE/uS8qtzS5CXxa/Hj8dp
krcxFIAvf5PvoPjKAO3nxzJmc2ohx4qETp6CT7wpS2HqugSSQRvnsjq4NxPyQAKU
5aUh3LLD1TteWI1dbQgqdv85bwO2iyzNMQDx9p62Ty8YEOMIOuQm0Zz2ZqsiZugf
0i+VsPJ9JDsLB16ol72ElQBwri+ZXlYil9DZdzQOYjqnEtby8mPc1aW3lF6GLzg4
O4fG/8KSLBr2RA8PknKedEm4QsIFqe64gugVUUbr8AOYJ6UP14rIuB2bWnN2gQeC
qlL2oGU2ROeJpIAa0OQUA8syjz4/x8EjLa87P3d0tzdeErYaceK8itY66GOxDIcq
BSGt9r4E5fSUvOYu3ByEe616cY/2ZzJkeFsmAdZ0pqAHkM9Ab4gbTGY1qeTYZpyi
94dv+LycAcrQmSitHmJ+HzR65cIBI4+AL+mBhpC4J8efc/3+vNfXANTQSJefzgV1
aieX9HPZakrbDlEsFh0uuukYTT0MilcQ7YpuyS91iCWrUeVYhB6/g9FoZkhnhPR4
UE8DzGJmmyd/t6k1OiUaH1KmuVjh/6xpQpJmRwZQncH6Aef2+Qi2SPulK0ph4ATO
gA7nGzGSqtyL4kWqlvL6fR0eRtxCRJDZqPF1ADLfpVpEuZwNEh9SGN6XKIS0TwnO
b/LOpUm3DQ6minYXiae6Ci9CvLgn4ByETQpgraBS7bfjyKXbBy7qyBJyK3eZdPdu
gMA0m76J4DztqYxm58rFFLrYiLavF1gA6TVCAHYNDUU+AFAiVwKiOgI4IE6LBqkh
V0asalkZ2s9C66O7mfgzYsIsJPAdRGTUQTIcDCbexaj8E2U9ZyKtXjbM7AOZsSvJ
vpCPCnigTB5hCyYZOYM4brZ7qvAjuHF6tn6MLeaWJniWonhlQh43UbNWEwUan9CA
noCKNTKRnl0rHiNSO88WGnDAhppuMcyD/BGuj1nCkbMuqg01P3rAbbtnyU2qFg2t
0rhWzRcGedO4109IBfvPhnzQwboBrK63IBWkKZrKzdQUjuueWenlQoT1FQDc4v6A
HzZaXXJ2OzhKRdGlKpe04JGPUwRaCKY/zKzBeszAItyjz+wlKXS5K8aKiF12p1xD
Gc+w0P11AhkNXh8nm3tkRwa3DzYs9C4dOagPv7dkyEYirksMAfuB0Nea7lZWgshl
4df6UFuCPy0JUfoFXT+9caV7IBqJpQejmeNdd9l2+2Loy6vHZIUElXXnF4j27bsL
pPk/FHlBWRxYY9IA9LBlkQuZldG1wGkXWoz8gT8dUoOBiUqc3X5gH1KOECUnLSrP
D/V/DRHqbCXbpGyetd0yoh4l10vYDfzBCAhTEzNLckHA96NqUteli5d6VL5AKPMe
w6NWE+pok9mCoGoFsnKnaKpKyTgqyFAPeIrgrhaLdqzMV96xJ+ir9P7r2fcZSzD8
coom4fWere68mCFzq3ijvpglebQdTcNQwKTxqhEVdHlxHxc74QnHJlVPPYfh/FOF
gR87xakW+4ysJUXL5Nm+M6BwNuDI9wFflXmjsbuS2iwBrcrPB0uINx2z6aBpcQVx
oCLYMFThg4T4PusRATcjwRXOhRR3P3F8IqBfXzlUb4T6QpNQPNLwK+s4dYvkE9rW
ac4NIWT7vb78khBxC92PDT0EHCdMHaeq9181YokHNKdLdS5FkDACFX+77A0MBvE5
ssckmgRPfvKjGxV6L3hsz1ImhpBF6SqlT2wEbOdA5jIqUV1081eNAZ7eL4IuKnQo
+mKGO0dqFiIdVhCvYywuX8mXKZFSVEMiMB6iIQBqgc/GyoaRldWy11vD9MOHe5Ed
Cqe5NqyAdxv4kQqi0ZqjvlxKrCSnh6EqcgY52Lsjce2ovHHcpd7Wk7rI29EwkI7U
qQvsXf6Gv3W+hSngvSxB4+9yrHSGsP83iaENx6tyGzEtH1R1btA5UP978Q+uZW/i
NTVUdw3OTFMkH1CF2Giy/5Ie0XdQKRKbCHPv9wlnFpJ6FZ/AikyGYODPnOJ1Hdlb
/WiWtSbYzNSkJIPs3z/TlO3NiJ/y+G3MXpswOyqKtKBFe1aR8G/q3aE2oAjqCEUF
6ukz9bG28+A8Ssfc6jV3HejcrgU1qoY152mjIBdX8wIfvb0C1E00nkLobuSTQixM
OqeSnwSwF/jOBk48yShynq/1qKINki/89/JKlIDeEfe+0GaqbJYS5ooJNc9qbig9
8kcPaoUnqozUbHHrbC0BglQ3QsYHoK2xA8Gd8FlnC9d7ItN2uqDl+HLd7IKmrtuq
bn93Ax+gQ9eus88jMD/Oa27S1Nr3R9VhrdjKuwu8I+ZS1KrZcp+NTlLIRb1IrT0L
l+NAyR005psMrhdNlX7t+xoQPgLMJYTAVbbjwqb7TrZFeZZftEgk+jJJhgarP7Sa
uS3cI+oLpchJMDWNV3XfY7Mrk1LlnUP9JBwsbnS/6Sbtt3glAwAnkbW8D4oBdtHd
LKYD8lC1ZLgjoIrE1CyM3HxFOFa4d84J95/y7l/ZRdi5QsacwbYdswodbR3NhDwJ
I2Z6tZpAntsLsbQB5iIpEXCMYYPzNQng31gzh9R6y64Y5JeJux9wuyUos+1cb612
dZfsp4K6NFSXQYGXS7kYhLABpju7qiiYibyv0rLXeu8kNc407YguNpeW1WEJTbaD
TvG+avn5JToFuWSEYFnkdGaTbh6TKqxA2gpmFbfclRK79J8ZgDSo6mxU6wjuWqeM
YDVVpzBWLDsWSd+LCWBPAQHJ5LkzctFdIFGmRfxgf4tpMjQwtq4ge2/QzNZbVLuB
8WUo1xX1i2bwlQXPaUY67Vl7okWDR+dD0Fb/78bARmegiRJdUGozXaK+3xygtfzR
OxTwYsm+tynTy05T6jcoI2FOsBOLIA+ExPf3uyOFUNg1sVBQh5nSvU3FHyrUckhD
DMcaMMenUobxOXryqjBas0ubixfkgx966RjNwly66DYnE0b7Dj1kSFL9/ZIb0L9P
zACrLi5MD1LTM4Dhtvx337kLAq6aMj8imrmMlup5BOpmkybe9xMOYiYNYYzoojGF
OkFjxdrGttrrGbD01tn2zSitGPZdrBaFK053V2h9J+RFiowq/ymn1mBbgLccAF9Y
HnYSZBeMbeMlGFs4sZySgWnHte7AUFhK281m+iFckdOf4mkHrIMA8lUoCzN+Af5a
4mqbC2PPfKjVq/jO3zIJnMFedMhec2vWcJljIiMYzZDcIvK1MqVi4tLYXR/2e8O4
xUNA6dsm5VlULCB4/rrq4OkjAjcApaqh1JhoRT3ppLvaUCqKjOEj70/0bIkuRkXa
MO+dSz3hlr32nF56XR992srffAN8yYY7KmcZ7GxHbLWzp5pydpz9Oi9g4bIPno8I
krV+Z/lbvXFUZws52DV2N8PZoglxEhRPwHRF3kDFWgH48eJmXKN84yn/9uME08xa
eX22vTN2pwfoRWpRX0zIwsQZGbo1qhnV/8fa2Lcgh+kM/+xoLXJZCKdTiHFV9pXu
JJFTLcRgnDjgUIZW85qQWqb57mQHwuv9siPA5OmyHAirhXXXw/1P2G6dBWhoNNg0
pZeJIQaFCisa1XWl+m5agSI0MyUp8j81ilrJak7L5ZqMdNb5u26l7L1eiXtwYzgj
lxwjYtpmXOcAPVjbFKhUhRSVKJtxWOQanCrG49GTDDPSYJbvzUavL/FwMb3NAVWm
YJJ7POP188DO0I6B+iTTd3Tt6tRvkN6P/4C8OzhkE4k+d3fFLZXMPcVTo7+H8CVU
o8xWEPzsqf85kkeGVPZhK33CsDut40YuMKpfURSCeqAaLf457YHfxm17Ot/k6ysv
1HqT/9kYXvs3SEURKQaFqHX60x+4nYya/898gUMOD6xq/j4bWLd0x4IbLP+/AVuz
LptgNEuidZ69I3lS44V9V6+n0L5yLpI+djggn2ngcmAou2SAq4ZxxrypZAmL6BKT
1djwiBEHEVgs9QkTF5RRCMJUxbKp5CLbV6Uq1SfA8G+eNMRVH/1ivWQpBQomgAQu
SLtO2007N7KrLLpFKczMWDaqyE9oSiShUwxodCLd5RLDNcZY+Zfr3Z0AmrXe+J5A
U1kLzbhRK0VdouyXOzMc7vltCWdxHnbU1xfchAnc/eEoUwuCzj9gjo3cd5XCi5EV
UhuKfZISKzoYO53LBjox5isnHnhDB+g35wGGY4GMcjcDD4UcurxN0oElwnqwxM0Q
5YEe1flL7UTpEKZbmPsbeueWLh6Ru7fjjaki68kI7ijOHhe0F8favVrjgi/qZhTx
kqYVp+4IYFMEtYAqmq5g68unDdJs4+9FQICbj5IEOYtAHJQ9vZoeYrRi9rNJwr3E
OyyB++ZsLFPt6ewgJwEyUKUoOOXPtqB8174HhVf3OfNcUcf414e8TxvRcvGwsMwT
rryWLS9HFjYb3co2xxDRqyXLPcs6iKBVYGVGO/tdb48LTucz35hpm3jLzwLntkrG
48VUAbs9I83rwWQ1K9HoNOFUASO/+tkl6YGRbWUWs39kC/QmoCjOLEQWu+Q9ycDr
vzA5heiv4AgBFlwdZ5/cHh9rewtcmriDk0TysEl5qmtN2XGGJmZ6OGoFQSupNXG7
7DVRefrFetDTO6mYUZpIefRuAAroA7fDXM7EyAvKOEJjSlvj1OIJvzqyVhG8mp+1
Mn2k/rCCOponVFqgmobn0yOVsSF+ugHZLDCh7t1pK+ybwvGYOBu2BrH9+Qxyg4Dl
XUoEDWVBZGxOQ+xk/H/1JXsmz9hEYGdFGMQMoqFwhQoZN+jWt5N6lCiiZFSXXyoy
CvIO5QKETK7HHjtn3gOKtq3vRdXLhSQ7E6+m3GNjsL5fZZ2nsJU6OWszFj0We6iY
3JF9NzJMcKzbhR65WIyC6G9WHP8Toivdayw6P3g2NsE357/1DIdw6+Yv6CYAK2dB
Wez6+okrALlYkniKztPHZVsOFpDB8B62VcLgzlmB2G2Ymfbi8LmkO1lBcHM00Kr0
0vipzw/vb3LXODb/fKAo2Q0DCc4+I0gBYiFZA67wxDjAuYUGnFg1xPbBB+hzScD4
yOYqPBKJ5+8mRTZ8B6f6HMrMvg6o5StHneJhjs2VkXjYeT2HRzMwjaU6vXIQgvJY
JhMo0z1tdvCUczKLIyXlFEFuI3MQoNeNYBGxt1RBv7p7SYoepiiWhGyT5eDSoEDe
JjcefTOlWbQ0JOsjfEsAi3acBihTs2AgKrOkO+/XercVuuI3QOnqYh4qhEur0P2G
6jo5WL4i20/+S2esj39UFFWKmWDuQiWagUQexrMo7oY94VXSdhesqymLkhaOQSpf
o4pA744vIWCk/LADkpcdmjRERrUDVvR3PsCbIWo/ahxsZycR5SUJG1elyLkxNVOE
c5V113dlLf0f9reJQzyTXOJWQH0SjPbIBPO/o74m7u5T73C5RwfIfGH7ovUoOkcO
iJM1ScPwLaMKr/Zb3Xq8bAjiVpY6IQ6YBX2hFd71tBVe3Hv1HxcTnp00xMsBwZB1
+7cGIH27JXbyTknnJ51Wikd1otiOsdsaafY5mJLyUoxhIRv9QIy/3+99is9dx1eY
pNB2aqWANRExsPct4Io/ufKDvDvX/AJshWYro8XlOlp54UDcI7E9nq1Ju+XhIzGJ
VfMn88CTsJucA0rc0MujN2DxFx2YjWXUbmqV4cQkGhcowh/KImhyHEFU8ncjIH6i
F9AjAAmXCBr6wTXAFGOj+7xCZzAi0eWqAVC+JsWCBPyBap00dCXRioTsaX3p+xA4
SbhjjTuR15gRV2FRWb80+EpkCUT5hjsZ8HP6lc8fBxP0zmw2wvEg/ZEGY3HE2NgN
hru+VjSPI0jeAMWvjv9ERlJ+kNU9iIRTlDkZFeJGp49vnd+JDqcbS4ZKVdhW5dH6
s/0Xh13pqcLQnmmpw3OqTfBHQOWbmkzwuQBNwWFiZzUx6Y0A/8s6lixDU675YbeR
IwPBqW3b+CrndE7IJZylNipmnqMX9L3Dp3OFzUxIotakQYAJwycbumanDuGVrKYs
Lmh+1EeRE5Z6+WAab3SXZn8OSfwpN1E+FtQXHvCEQtUB4i/PFf0DZUwMxFhDtIsu
cm+M5dmApmHvBuRirOYINsshhJIkMSquzdCbf6+JML1xLdg09JGDykJ+HDYp0Ckp
jY3MXMCw24mtdCQvI0HzeE2Furs5duLGiPODdhglM7pklr6k0QCJJVv6yn/dIG56
zFdmjTA2sE82M8WOIA0iGNF7KT8T1/F1ANVjL8ge6RaVuzZNeKkq/5hZWT/Ctaqo
fPv2wKpQJZWA4yADv1tps+GLAO2OJyNJZAofllEqyG6IpNpU2CCBl/Q+yRHCD4Q4
EcAbcdnvWM4l3fpeJ+oHafIoZzxOyl3ZVXfmmsK4uTT8opvhW7C5sxHONKFOhkFQ
pKH6JAJt9bqVVhZ2k8jtzlxAmur6yKQ7nFVaM5Rm1yPi2FlEfW0HbLeGsX+oKpNS
m9D5eppQ1V2rnAXKzvPmE39cDaArnlJ6imO4pmlayIsAmTQCP/O4L1KDlk7cH/3O
PqF7NXLcMqbP9Qwjlh0OKIhKAyxNjzoAaaGBD+TB9qvyHsmxkRnZrsUdWb5dIpD+
M9tlBJx52JmaDnbA8PleICiYdt81PZAGIV5UkxJAUzgLjrkK+PjJ4y+LkXejyl1B
5JWf6dAuxZzTdZg0cuukJ4XgCzLgu2VrEeb4bSNoI5qFkIa2o8FiH5+ouyZ6To/8
YsErhIAGkyFgF8G/ocFi+nFk8vyd5QiFwtxGiB+qqcG+N2wSmLPUollbmp1vImzB
pH4G1qtgwdbm6Hl3qBJ5Q+ABvxzmj35knaJtVkGDsdJlUQxexQXLlQlj3DJ+aiQf
d615jdfQKTg4cjCrx9GLQndRi4IZPOShFMLkiX7Xn4VhaUwjz4PcKm/5U7F938d5
c34ezw5ZGC1WxrHFERKFeYCAZArUaFJ44G/BLDxOoHExAG00gC2wlNSLWHShNGkU
juhqnSjMqRTVkoGKcvTI3v3hvxgKKi5VrOQ9c86Evo1sq7iHB+WgOOMrVta3t9Nd
4PSa/9k6eY8/8JwPTxM0bGu+WRYzi2RUS81WO4T5lEaWNeQvLMzDhRPx365NoUWr
8Z8Z72h7J5r/7L7T4JuAN1x9k+Vf6a5iKXAO933NUatkjwjWziLTEY5QCLdUYRSw
4pZZob7q8Q1DyprQWAgsGraQfWkyFnlAYSHtVR+yI9eoZrvECfLDprhukfkEfBsC
Vfm14i3S8nyGZJEqvDCqUonoCi0WOm40Aa3LIwd5vF9oKVtzDwdIY2Qdg55T4QSt
b2hRg0sul7DXnDhNm3pyBHSxSwNzxDjTAG24+AYPx3j8a/rL+SdzR/94r4PoDORD
7vFDl6rXup03WuY8KAuopY8npRCxDvJ2dfcscg53SL11qUbVOO1Urt52k/6zBiRU
xw1qmR67ppXj5yaV9fOe4kRmD7lv8VLFLiTCQwMGUIi8qeJR3MpsIFY14fEj/e2A
Xq4KTOXvryHF/LQq4j5OIcsz5eCC4PkpIVloJ5l4uZ1zXLNjJJW/RpcQNd0mBMi7
1HTEbZkw55gMgtmDFA2IAf15Gu0clBimWruXrNZCqUbaYlQMHiTPYJ2JY9SZ3J+8
Tje4fEcWS6RM+jTe3S/ttRuxccEbdgzjnaxJiQtmACmT1FJ27oWG2LwmwRL3NpOm
wA2wO5bbpXCY010ugRL6g9Tioyo4lSgH/ziHt0rDwYibJIw6K/UWlBirFaGV/YUq
NDZXvTGnwChjW442EAm3mMWiy3V9T1EOHoD6khwew0LC0XM3TXyxi9NDEuW+KMlz
/ZaMeSqLBBUr0Z4aB54YH4GCbAbMq/+tXHgbeJfJBc5HgvZJfH8x221GS338c3E9
yOv5RQynwsM7J+t0RDPG7k1WKv1PDt0bFDqe2uVN0WO59xik13AbsCCTQaCxrU8H
ZmLynBCtIk29TjDGTfB1FEg167TbfI+6SogJouG0+hItlXdVoFqab+7bl59KwbdP
1DUno2eqi+8/mQdPBD5ScPZYHnjHrumOusWhyy0t/UZtPAwpEPf033ZeM09uNOMO
1p2nbIeh+2vQXK7T53BM7oucy8IvoUjTMxcMKD8UvyhCkqNbORYMiamJUkUcBnN9
dnzc/dXVmsa+N2605TPuKOTjwX4V9tfAUg4KPm1kefbX/VHi9KTZI4RwIpPJtPc5
ifGwEna92R6G6UCsmS+yKdR6WFe6P9A2e4SSxU/y5utn7GqFBlZeV8O4Yqoi7AL3
7x8LPnwsNlTqAMH1plRKpqH0E0GZ7+mdSxoQEQ058/HHBktnz0eyBOsiSYmUbS05
V9zGYekesS2ZsAdhfOAVL70DxmMaajtjxkKXMgCxYshU1bdGm8MsMfa89erpZ09B
ANVf1yfi1auhIVCmbbN5xttNbkTmsxEYdoS4pISz011znZc62e93oDRn+VUSgSA5
Go763O1MiZC7T96Tb8b90fUWWQhGkg3DbFtmGh2tuKNYb2adrcxJt7xpyNY9+EXe
A9YR94sGqqS/sT/pjLxrgvEj/EmQMKWjyHa622XIrTiX2hmt0qhAoW/nZEni1s2A
Bu5TlAbKI2rxCV+8PYGfJC7YWSnDCjb4FF1vBzQjgD43Jpt8S5u2alxklla9RUgo
kkNLc0YNUSlpAB6o+Dy63anRH0gdGtwk0O7VUjKcIUGs3nOvWQe8utzWIfUv5tj4
ae5pkvju8k9ZD4rym0wzJ39KP9Uf72M4+4mnO8enLF/9bQyYuexAC1ZEWKibmCrP
ab5lxzAAd7GX3dqZ0SuMnmOEJdO+iW7HzDPTxdkKF+53k82qPQn0GFL2mNisfuOT
LVJ8zjVka48f15jdnQcFKPWnQ/ymKs7uPdtl9USFw7mCiXIRrZ3womy1EXP0zpwD
7cXjp0tqg1DG1X72ruxEUgwEC+J3DVGEBG2XaRA4mwEawtJlaDX0B0Ibu2HpfZaH
3X309IpANhuPgjXQ4g5YmExTSam3NSqPr76mb2pA50FpGaFHGssnYnc9v8I+qfWx
v2AaNPVqC8zOBOqpdiem1l16f/lLz3r+RV+sma/v4bQYJlO8nzlHRieSkxnVaz0u
4E1U3qvU8I6nsS9jT0jlPhkBg6Ar0Vq9g04hTxuYC3fMB0pBioB9YK02yyORluRv
NUBAe0YuoT5gPE0iE51Poa+hQpEAi9hZJrHlZgXuCVqUPuqEQ7KgYuxSVuNWAYfN
SMh+EMMCrBQRpCpTSdH7KMxqQfQnLLTKETZYOFcgU36vHKB8ZE/M7R8OhMnFFlVd
AFFIRYUVARwZw/rnXRO7O852+Tf1r6LLjm/6lwUz2BPKWaYClLQ1RkC9Qa2vVVO3
TaplLWIflzL0A0Nc0OTAEM7LPd5gauFqQF7gnRfnQDTSUdlNG70EJbFSs48d6pi+
5c2e+DLxFMNqVX5m2J5O0oyLZQbepaOSl7elnomfxZNprndTAV4QVanOgwjOk21W
RbHEtBpUw/A46cpBOLivVQsF0dpqJqls9J4chkPnJJ24Rcukbu+De7coa7/lb2OE
JCE0kwWDrg4jxCz4wWxMk2AUCiECseg76KCAqZ+jo3+o451wpZACvy72WcqNSzJ/
hMohqUJECzKoKZHduJfvj6Wplxv3JJ2hkW5sA6vi7LHz5+8kg398dtjxfuUAfw0z
zeGKr1Adyb9PMVZBEhrN1fOkbBlHs1SK/Y0I10B1I68U5iV3ox2vJZAyOerUtpTx
bkiXZVpjcB6ejJ+EGQkrDRDpt+w6hrMlKFowe5oABPDzUktbMhUzPt2a8syAqQ61
dxruakp6PrOZ/hzdnfVTheFi1N6i64c2W4HTzNRD1k1wVwpc5S8lR00ZtSUmc0/g
hKVsGaKeF4frwDxXeEd4gbmGCkMokpg9BpuQfUHeRXW0ceh1jwXzFJt0AlfJo/bw
OTamTHrGm4nErCDimIALoE8z6RgMbIV60hIW4R1Z3OFpyW4wmswjwjaDHPIDUR5e
HpMZDESTBHZ3DYYPBSrfkbTVxH5NUrAIOPRYEoSVEKGVJGT/hcLA2l54yggIJ7Xj
WRvAYYhNs2fQ/6PK1zOx8quETNLdIsd1StM89tOFrUcUPDCQ+eXpY+zDhSX6l3Sk
9QYPjEw25tlk8OUmXjGRN3Q8jJGRb0cts1yJkuSva4ASMNxANa0aJYKYP6YQTCuJ
VZXPXidTqOvXwOGMkQoldcvyBDVlsOqgNBfAaN2iF2t06LGm9Mr2KSbVqiFKQn6w
Bsk8RnV7sq0VTPCap8J4SIafOG5ObmyiqjDbpkr/SFwU31Eoz1vvWXmtzHWPwxc7
baoCoeGkmQmYI6eIA7rmUGZ3OW9j26gSa7hBf1ddzh+KArJBEjs1Y19g9uEK/5Sr
fA1tywarwbkOSbxr0TJGSA9mP50s4V8UdAhjGfJA1tPNe65ViXcyEmunjD6qH9A8
UYXahZbn8LLjNd2XQtNEfTJnTxBgVvF4fJKmO6njw+dYGIEpehKy0JSIf+1UlWB0
gxyxznF7aHnL4x1dr9w453OvodHrV4ww8JudS2jZ8GBBaftatVzttDqLsN4THefk
LAjEmzh/0YUVW4Fqj/riaAgy1bfYJ3vyEECg33dMmmJV1cVuTRY/R4BUaulOaqGn
B6wONHuRTvUGDLXGlX9nTHvzfNJroKtThKmvN7z7B66ce+qViE8mB5hNIVJtSSEW
UBTUqm7u/ASlBmA0XIGGLDk2+V5PIn4TEx+lIivB+kOZcSBVUT2LQg+9+HS7SlGX
0ueorb8BaZ66QqKX+ZgR8QfjS98UWyi8HO9cNDkCQ3aTwQUqXbsZjTp8SgOn49vA
FryRA/Q0OEkAJYVQVn8wlNWcavLKA7x3WeIvikDiKjuVVngABYqIC6miJV+q7UOX
9C+lo8+kf/RfCHh8OZUo+sfCAj9vcB1TDgCOpU6HPA1ids+/yjRl192wOcaKUOdQ
VkPYDfeCRcosfxAiJvARvSRCCLXmN3lhCGy9jxxvwJYPzzxlMnAvkaIyVNBWi9n5
Q3BlREHe/Q2APD3wWdyzWUFAl5LcM0NwLa1RvqPMXdqkLCob3X73VMKo7QkuZVDS
2ZygDN6tr6vgULvVvqF++qFLTS2fym1VaABq5TOv0Dbh8RVjxD4MtXAORAgyilcB
74FNSpqQWpaLFAHvObn6vWoBYVeT75ni4mjr/XhD0mv+IKW346qcTn9DIpRZqUbY
ff6MaoysmbiLcn6ezlyRhlq0WsyaGAra049g/sFj76FVypJiye8+ooENDW/bc/QJ
jhqSc7rulwCST0Cm9K5NSyuB7Thu2cTrGQhdh/AbXP+WKS0dPOHmKwYdvhq3TGj6
x7HSwgmylZbNJ6XNFUJsww4CuCVlY1DnsTfoh5+I6hVT/+DAnrc5OX+ki22TsSiQ
PYyEhjs/8PrJmdiSqFPgCTB/bV3EhoY66Mu6TiGUW/iAcNFz0PrpCXn/USwD1Il7
NGRf6VA06LgfHmqE8et+1Ph4aWwNl3CDo1RA3oHaGjIzhNHWKqziKD9UE3av8CsU
IjYiJfsJlOSKQkOtX0viudUnbxr62TbZLfbvtfyR8A9QWrZAlkDo4vhA4ybg06nQ
IKRYyVH3teueusvNvJJXy32R84CgDCBRTmrYLkLEOz/1m68b+agnS62n5z62+bQ0
vCcDSWidXdcySijy3iWwSpnJL4sSjJEP8hvBrHsy776Cq7AgZFCShfi0WBYtIcph
sKaRmSu746Ai0YEdTcGhVc07oFeJ6h7WdcGpbgPd52VDoZwOQLX/HM68+JX2BP3w
sR3Yi9ISmaI4hXtWunlTDdUIW4LKLaqL4Qe//a09hY5eodP8m2kCbWacMzpx2pMI
cnzGFNX7ZMDZoC76JzayoF47CcgXJsfkNkPO/7KRiOI3Ds6X+y2GpICcYNA63WL2
udO9hIpUZ6jamkB293kx2iQzp0lbshLtzQIMVBG4SQfTnTOfLbT6fzzB7f4l+HwJ
6rfUCPEv6q9n6tpF8GPHDDld2ZyK4+ysBCFQ1GiBnFGqW7n/tbdx89m93japDs3i
AMnSoPz7uHc60qRfiCRL20v4aA9Ukk6d9/TZB0zGVFWUIhBHqTp0lfR6KAFm5Hr7
XA39BWsb5BxbXeBbtY/LnWaChCvowDm5U3XdnKQonrgE6PamELFLPIhyrTpu2HT/
FbwpMtgY4SUT5tQ59YaT1GscCTuZgWVY4qY33Ea0JZZs+Elf8neKk3AKMBHKUaTx
D2Uh/klXSo1S55gM98au7V4zEegcXO7wyO4HTNSTc38dqpYb6p/oY4trhgo9qezC
feqkgdTfWhLbOpYrQV+UsepOJ5xmTfunXfZtPUM+if0ZKraunCuLhQylmnplCfB+
goGcSYq1qtPMiAuCuWVRqWbuq8YTc5yrg/MfaX8q8OWGEg3WNyGfgvstZR50bjRV
n/7PQwvGmEcsB5LFCIeiGas/rJRmBUtBJ9Q7goR7XipUbIyjQvq7IrDgvfUXLXoi
PuTix1ra14DUxbmi5VV874YvDlNScFARQrm1SojH/vheoZoMxpNM7cRbMk2g4nGT
W5YA5/iRGQ2p/at5qmH1bF+v/1JlGneDGLT7JZd3ICyETr+LDG0DrHwQg988ZoKp
ca0ISmz1vZ0Hywx194WHiPvva3e+DhDy8+6OXkSW9W0uNt16ltYPJ7N42OYv8jZ0
GF3a54LQjmT6OGv6WNcPJeQaR5ToVmL1N2QmIKavYzMdbrmFTY9dAEhXapmKZLYp
ep91YVk65xHYwnP985n0oP3AOrZ78+I7SgPXAU221/OxoUcpaNPqCwIH7JDJ8woe
6PjtYR86Uwj1yWtalozt6heF/POq2sab9gubkiMopp9DFqmWay1nerCmIfAvfz36
tPL20aGVSapYY/kpHEIsBXi7M+23IhQCNVDHN3hRismARuTEQM9EPqTLph1cWPpf
JJRQqy2Zr7IwmVk2oHSfyEPz4pGD/V+UrQGgH2+Jiwco4rLDEjXgGSzXWP9AMwML
3CjDHu2v7wHzsbmQWU0cd3UKK44fpbLeixYomaH+HrNXe2cZoSTrdipqzhOPgObe
3zXiU1bgXDhq3WWW3XnhMlXt+zZVlr30S8ghaHzRY2cYVdTD9IT56TV9nZoN56C7
C2oUDiFaOTT2z+8WdcN1vPBVVdUtee0DABQ1gND0z3DFa/ZNEWDrbVj3tzJoxtS5
x8J3kWWaqOJDtysvPV+EVsQ1p3d8nhH4joRLQ5MU1PGxDV42gwxl5OmNljgrkhq5
4H2uFzpTfpb0C04Uo8P8NaZxl/jHb4bzyZIxt1JT+4xk+A8Y1Hg9IA60tTynhUSS
lW42RgSMC8ZcTMP/EymFGPLoo5alPb3RSRTfCYF1SaEV6mBUfxrxS/dEE4hPnsn1
PDhLaPNYIX1wePjUTCPA1YKjK5fQX5NbQj+vNzS/eERtQ+vy/ZI6rGMxsOwhHFZN
PjwRL7ZmJHNbI0/kUBU+ZsqwSJunD1AYM09cZgS3JNMW9FmG+jPacesIu6JBBwZs
1mqgbegUwLd4fDAmfWVTxg7yU/VwkO2pG9uo8J75qMzcEhSbxcQWxc+8xGyj1N7b
blSS4oYQzLm1F2Ircox7ZgSAGWUZAF/fvagwGetgvpLEWWwyxby2vhkgUxtp1sBf
q6ioVt5Q8aDVEE8rOc4zgC0qjBrBJ1+8fo9YHhgTEu9pejdx6dT2eEr5ZNCLzkQT
/aezXL043Siksy6tz/p5ZVJqEotrJ3OCGs+TC+FJLKzHi9lZcfmKBsiMfTdaszqn
PeV7COcIcHhe80Xbhg11Lu2sPFKfW58wyKlt80TvjSS4IPvTI/z4EqNcheemAzcc
ns9iKtLGzJJ+u62N169byTRu6kknNQrOtXDNWZFr+g3ax3i0aAL65mLNjyoTRUvn
gFz7vab703Na4faVkZVuYObLGmpEGMO0PVoLtJcWtpc5ujYTeLixkRMX4QGXsBtT
mbsHu284JEYOEEapaLW7a8G49RP63OioMclMFwAtG+cCtI7VQsqX2+vHTy5LCk5V
iBy/v28tvkt3QR3nM1J4gNZRxi1I0T20R5EnzfdzJTDer3vmZ0TPAgHfMxa8mm7H
vVbGrj+UvRJ/yTv6M1WUCS/1Yp1DchFWVSc2A+zH3bDw2P71g3+89ZZuXdspvoWm
8KR1aHQ82o7VzVmBaEfjoaCuDlk+SOcqShtTvreS4HXd7gkp5yMuwT+D16ARUer9
AcwQ5aNOeqBWyMhcB5iHKYkM/zes3vpjQUo4+ALqahE+PQxYKC4Y7A+OruEOhM/r
PpYL8GdnhSCb3JMf+U8p7tU6LTNZ+7VM1OU9iABcBKV2tqcoPgKcPQ7dVepw6TFn
XHa8EPouuWn8KShNwj/W1qmrkV6WmAu3M8q3+R1QtGX8IHbImUenyE+qT2eiwLMd
3aCKl6YuQa+eJwH0uJahOrSmznGy5gcwRvBPnGKH6ETK2whRp3xQbKydJ2v/T3qB
xOToS+owO+MxgeC6n3q7wvDvhqM04Hkc9Uko2yFs/5XFT7oiFTWG2OF/+Sxi6eYr
ZcoWREM3Neqa4dRBomegsN2hhCcGFEOUCRe8UBv7d6DmNPS2+/hLJOqxspj0m+tS
jNKGt+gDHXGiKx9ov1po61RB8PTyABOOrDc0ZzEGgNzjFfDxhnBPApYb/MnXsq8t
nUFWnGEuSSV5IRKNPQ8rTJR7+1fiWrqAUZXwnubHcyyvb8828SwInLoREXEwIJJ3
RfJ/HTOkomCNJXmVMnn4hja9nZMEKFLHsMidvUTSrAtLm2pxDgGaOfoZn2+y7wCV
7ux17e3LrqxuIUZZj/asidXTMDAKah+mbaYy+J/YQLRSoAMIBDpOO4/AbFNm90OV
7I7qFPTKbct9slt+umSP7OjKyHeDVaxVeDxSRjr0K9JM4sm2OsoXBdyj83DmSC75
FsLWYvrDqdtz9duJjPUjYEyvqMv9MXHLAvUTkBbVqxz7UBZdrzgFiAPdg6MqbGZ/
6BcW7gWLb2IPu6KSwA1mSGmvTGsCG7Qe2bw7quHEuZCpLcqhoNAn2BD6UmVZMZl1
5N+/90+x0qiv82uV/+EdCUIV93b/R/4fWo+xUwcTrNC2c/PsLysBrhTIIl/ySqyo
xdGfK5svPrXqXMrYwufdbazxG0FjQx6EIAl/2n6COGbNKh2Wzo4dkg/4Yh8JkvuS
CqeGsnhitqNrhwe3z/GkKTKw3PWSHmIF/WHTGkRVmKy9UrVQ/6q4cV+szs2wFvTX
YxUriVcZullqiH7s0AJm9dky2/gCnryPmZoS4ydZuH/Mqv5apTxnJdtUBtSKB348
A+P+8LY2yDVGmuFayPVmXYl1rAxf6toRrOmc/DvATKunSpfFMKoQcKmdPLHNxUxx
BRVgXn/sM4Zk7VfmROpohRkXQSQMeczgaFxcbMsOBnoHYCf4/l46tsft3ig/h52/
KB61YQE24cgJd5a5RS+eI+8UTrnSetdJ+QtrVCzl/+245xSl7SBbCwkawm2Eed7w
OVlNTBKraEHkrIk2J+EsJXcUBZFbIrs658rDafL0JCqr820bQsXqW+T4JKTi/tN/
4ddMVf9Va0FMffMK67N3NzzXbXBJTyDl7rtutC6StJYNcb78aiLEyZFjzr+/6pfA
GMBt9D5Ov3M0eLFF0HaY9qexa2kRc9qxYleE4kNTcYZsKhiRHNFWs/Uk9hlX0pLW
vc9nTNZDAGQEMEB17+jyY0c0H5vfDg7McAlDSUdFKPMquXtwf607w1UXAFbF59pd
b+kqzwgVKotkGZ0d/Kf+laIzEiHNapg3qNGaVtJiywmhLn1FKw22vubfcaUfPxVU
8tiJjla8n4SQ9iJQs+cQFzxPkAV1CCu5D29X3jzpORfdBwXuzMwBe5smds4yHLby
esNBuFzRp9msrUHCBMp+nM0NFQh6mqCPUIoKp2KY0ldAYYfVIfnZWHmU8jCoDMEf
zLDQUEdvzsceYJUfHAWJXfQFpoWtvYNI78feNZbRXTgmIcf8aObmAXfDKwjdpXa7
3FiZvFTKRmKMUBMisyTi4y+zRsCFczIQJooJy80f/6ZmLkq4m5W5uFnsgJ9HF9Q6
My0gxX1oRojc8+Lz7UpoD4dol4W06kAyQd495bXsB9kmvi49bWTYmrKrac+jgU0J
xz425zV7gIII1LpXLBZFmjZK6MM67IMxogG37j2WytF1o1XiZhp14O9s6osflEbp
Ym18Mp4IuVtUc9nixDniCTcY1DTXbF1cQf/Bo7WfAcKGHVQPkwpxn9iHqXZR8MlV
G7W3kTNS4yr40hWQbJOABjyxMbJcJfU9csI5u7UYwqDzja15g55B4H7Tz6i4oYrl
H/KrRyM81pY4/mPuoluLEJyfRNWG4YRc6Ay9lHnUuB/2cp7BW5L1/OFBJdGlMocK
kNxAqAMA9cpswLqNF6JxyLTbB/UsB3nkkMtgtwKqf6pjWZl2RONZPDPD41zvVrP2
rmdCY1jXKrBkZ5T5sYqLrM5tbfxBMOGqmwsVVdNNRI1M0JRsEeFZ5pV74L+dZfq9
ptu3Bcmg73ElpJ3c1IOe9kYSQZp1GLfnDf+Aiii8H/mvDKgkl7f8nDVIik4eviY3
KyiqfD9oa6x7jGx+t1lxA9ufegLKB/RURo3hYVQXzH/KShZCCCoqotvBK68BCTlO
OYdr/4QMRcLg0oPFocJWGTnZjbTtadaDrCoTPirrYI0r69IhExYn+5u4vv6tKVLc
hW2EQTLFgI0IhyhgVf7p3fl8yzT7wss1YZLiDhGqa1/4BaKLOtwnJvBaxTbSZNo7
TGzuXLBlqq4aOHJRFj9ZoDjzRtj1ltIQQk7CHEtoepknup/eZezmrjSDCnnAzbU2
bG7aOddtljOf0F5Q4Z3mUK/jP9RGR/BWsb+t8dtzMSEAw+lgFuqVbS8Vu9hiPjUu
qb2uemDtfyrYT99KZA6dHurgRVi5EcSqTGBTzWK5q7pB3syVjwHQN1fD9rTQeoj8
Aj9K2OhZ5X15eh+iSyhxAQk3SsVYSYxknmJZQokU66QzLWROff0JuQNIGTFskE7D
hrxbvXwJAmJoomu4NwXGbqQGRRwRurSNoYxDWtzxu+eTxVf719MU8HgrMIMVw7eN
3gs3GqnWmxbF/TFj+ll4jI1kpNOswb0B32nGSLMC1Zk0JJPrmTRJCoLeVkEaLiL0
VfxMcx15tCk5OlaGHOGq7U0Ot3xY6AJ7Nxw9lKF4Ex8KhmX8fZqB3yNLui54ugxm
xjPUMaP+6aB/cEEK59+8PaTrd4PZ5DkC2djIWlJ4gWzVSzlq5WqOvJfDQFDR8u0W
Antd5hxsxMsYzhTz8kGgt9PIelzzgW0h3b/gFNwcxQpwv+IvjbCPB6ujQx3pQNIO
Np2bZIBYCPRSG5TyZAQ/P3o/pNZagNLvEoZCx/0yIVMoouOoy7sJufJSi5wUTPtX
hxlRSVxJxFu9LvAp/pbbJMg7KdyrLQ1wvksLCUQvF4hw5Ll/kvZb5sCr42M1LycC
4wIKs6zak2UqyMaDhDef1doIEO5EYBnyp1Ld6UHNxp7h1yCxhrNon5qL0AHWHGDV
dH8HJMnBHOfLNLPUaIHM3GifslxBn8sFZEh3dVeA2aeJQzu/xwVycrRZ6u0da05x
d6HTh/2duP9yBaQ7/Rk0DoXQM7vwUhJlWgPZ8BVpT0u3viZp3tSkK26v2U87moBn
idusKv3A09EIJl0o2YU8R3wAGNDMy3fct+bH+2qOpjU5fy1N59BwYApvGbPIqVMd
lxyVgXHG+xcZjfHlerkTKVN7hU0bV5D9qMh/AI1Mo4uxuj+Qk/duUDkteKMwZ3Ou
Eilu9PkoWryqd33IttzT5cLppTR6K9h6+UmyTKJ9elgWylePVo3iL6muMuRSTSWC
5lNejCLY23vbreWDwtD/UsZdhphzyDHkU/qGcg4eoMhHChd7iRVuGWz1pw72Vqvh
KwVU6gy/GLgOOOz61coHeTm4uBozof/c79vn7kbllB070vZfyMIbSOyU3VZYRWlH
5+wTvLWFB8BtMLs8oM/aYpqNFPknec4on8vsEvuNXHijY+THep0cdc8fSzPqVsKE
G/Oxy7k99LH4s+u/ZMhHyFjXbeoLZe5kfFEo8zGDPviXdxDmV6dJI24G6WLNNkVK
60C4AoGV6stmFb0afSVe8UgHkJQDoyvZMRvbR+/X1HBS8sXmMx/eo31rb8xoEnYx
2NSLdhZ15oSnsY4TVJzBF5FKxKxBoGr/iCRQPGaXukjL+oBuKZ7kwbyz2MJWxFS9
18Jn4lx4tx9JxBeTEXca5uM41MP020E3sixivz/pTCfPHTOkpsh/tlha4dYzWrOl
d5VsxRrDMN3S1IL9HQkRwlvGVe1dQiUe9MMYZ6mCnUwBrj+1AEtnf7+rZBPbSVMG
9QSsWhgxkgbkyFOAru7dD+J08zm84UxazH3gXwYE5AJT8azCXGda6V9uh574SBWI
M/kmHXJTVU88n5zs6IjQrXfkRrZyKhRGLJrZm0uGCUCMVSmgZGWGk7f6e/x5FPoJ
7WLmRCJ8lQjp3FgX34twDo/iFkKDCDCsA/pcpjC8IzzM9cYk/coGpSUVl4R4YbZu
SFd0eVA3J0cLEw+37ypepL/eYNepUvq8zvkuPGSiCMApix3WVG/uES8W9Vj4jCps
OL0yowjig6chJeh2Rl6DVp5h31j+2D3+A7PMstKovStg3I411Equ21Tjjgb86IAF
aEmeFIxLbQy3zERn7qj53NegdHbPdI3gEJXkGH+O1NLeTYJUN3/JzBmT+A561iP5
NkfmgUrzZ8TG6s10sytTN56+7uY+T14vfkyD45w510Kz4ti5u0LuXVxXpxBFAKNb
W69GnWxtv80dySPGMZVYd8bc2ggzMUc8yeZ7A2Jp/I9pk91FejTrnpmcsrOTUI9g
z5doPwBL1RV6z9+E812PKn1HJp3H5kG4jXFNglms2wT4V1aB7u6LjcDDwKzIcbkm
AewfSQ8EaZvqInnbtgXLUgNIoE4a5txIQzu2JiZ31bU=
`pragma protect end_protected
