// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:35:40 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
RZocEN1buGPkVNB45v9CCbFOrH2pc8XzfvRlIRUE3TUnTj6C9Hvv81nHYWjoXUTE
75oOM+72BDDJRVhfMd7AZG7eHIqwJhi1PLPx0arB3wdIfbd0kMAIH9SeR4Qj6WJs
wqxUI6Klb5yrp8hqCHQHm/ehh1VTHZLK387s1AXh2ck=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 4016)
i9ZrHoQLzabat/qfI4vcvQLowm+Grhh3T9qQGVKSNTC6C7nF0bR4tg0dxh0LstCT
evad5HjRmn+I+WUPph0yel2lcCcSct4GBO0Lf5R+82DFUjp+peM/zF+pCf62hTBn
F3zzdSU499rbAew7UI8dwX5GSsH3yBW/oCLMHCwikICfDG7b9XszcBADcqk70SPj
1AktlFELF3Tt4RCjwjl5Pcnjsmail089GYKys/QlAgK3J3dh6k3yIz9StqT8iWAZ
4SWyTMgs5AWjwEp554YIP6KxfSWd8S6crvIxN+jmNDKBbpuc2mN1bczKfyLbne0M
uIC0++/ymENEes/RRXr6sUdagnOeifEGkGXp4s+2ffbaS5tWD3wNMwYmi654wKm8
wGgNOMFci6I1UoO+wvKnx0wYYQJVKoaaOfYIUS35kl67JZpGeJEZBdXNjnRki6hm
qxFlWozyCivtMeEp8EcFHp5rPiPFYYTlN4XJ99RwfPHC9MSaVLE2cPdnpCHyzXkJ
zPmGOkWPXxIxtVYyx/SbOJOnhwSI5FR1MTqaCge/dV0QlEZtlvvKVSwvxf3wpGmh
rtw/PdbZV37V2DiU807LXhx/EpKyXaxtwkT9ei26p/3xlfikyGK8AV3erYcFbaQM
uGmdrnfh1kEHCTXYC4t8+zGheIPjCaRSFJo9c9Kt2ydD+iZptnyj9jz8DGuNlIeU
hK0qeXZ4s17aBZ67p1TdRusSYEQQJL/kBqxAhw1b8Uqn7KJ6T4YmJALILkb6ZSOI
fMhHTC68tC3ROH9bmoSaJoEFelX6RtNiUBkFxu1ldzl2PdKbI1X+1prfHlehVubi
TYQgy3oYO4NRze49G+jsVMCDzkox6vNSqvrp/6B3E3dxkWxnNbxvJKX7naWGokmX
3j8wb9f1bWOrhLaP1GiRCJNfgmAaYk1eK52hvNgn5P+Xq5stD2avRGxiePxdpPhD
E4NQvANsZ11oIxJxxPdGhCL+yiScj4nEAQEp7aIYT7+1cSON+BAzB0na/WJxK4GQ
Pns5yvVSANmjmN52S1JCk+KKKSqezc+/X4nyRKqgdNgUafObz/d4wBKn/IJlsTli
bgZ+gNxgH5FrR1hcv+TCZMQxBpdXUYcCb43fC51UJI1alQU0z7Bgs8MPQ2rtBtK1
dVUsH3Dk1ZgtcMR14bHdKbgnFHLXK9iRWFUfuM2nmJH8L1nWsmfcdOjQy0Upl5UJ
RID4qyyYV9F81Lg27e7QNkxPa6xWd+P5Ua632fxjFAbttHgRxVpiHcyS/f2uyDMq
LICyO0rBtPPmPnnMCq2xow4hM358GcKDyp009nHxDPhOvEvgnz2gedzmTgfTKF0x
UTlYLJBSDnn+tqRn5G6+pW4Jh/jC0luF17OFTMF98y3KZUmpFwUNSe3zcCr61ZP9
SPDt2mpFBexchts3+jEb+X8DX6il6l34iC+ADkJ3TwqO4RICNTq3fo2O6pJsAbZW
7+n8gPteq16hMwSa0m2oBPo99tlKf7TYK0curWPvroxIaangov/sMLwF0kx9OsJ0
78QzOMNiHhU/t3VVAAGaJTPJ9aCvUnQZmSL3QbiuGQWz82f15UlgWBJeH1bJcrD+
veFyTvsnp4fqvHZNfXB2bEFyT4mpM0XkX5fwzAHMaJQaH0LMfhcCZn8kD+HCZUui
8X2QniY+9fhNFGX2vj4q/Ua++opA8mosWX1sUoCXUYZsYaInH/LtV1u6eFUVMX9V
vTaVYpYb2SR0qXinzivLO8IL605VR2G6WiD1n83EezXqbV2xHJN8mqiyPPLU/pqH
gW2qAZ9koTf5TIcbfEkZNYsDz1anhdsHGRTz1qx+jRLUIK+eyyaAp8MCJlmmTpZe
j1BpgfURiV0S/XEI3ojZLvdRueCSHLbZimmCqBFDGVORiDv5fSQJ+63R2CVxDwi+
jdMeCgB1Zg9Q4p//wTRzYvWTdckdrW0xhCNtDW2y2NcW2GLGBfTrDdklxbR7oBGc
xQGHsbXOtV+wTrJQBZ5r02h39Cuv0rGd+ac/Jw2p0aigp+KK83RxZ4OMI/aVCtnk
5xmzErmmkuIEOL+reCjnvrVJJh1CVqpsF1lCf16mU0Er/EQiuTPMSvZDyI1+M3a6
rtFaj0y/8OBrEiJv+lWn0Y7XltZFLiUufN/jhGNZmK2Hmxk/kLSf4fpJBDT/5/Ll
ikvWvX7DLwfmMmKgUMyEsksisxfWoFESjV+SiIToX5/W+grui31xxdi9VR9o3LWN
yUA5Osn8vQWn9dA29zKZUAshEtcRhEyl6hhb7PjCUsp0k0iBo0MRo/M62CU2KOp0
07FEywKQSsENYqVA6sgnBabgk+CD6FxhHWv3nuN4tm+Qra6RQRG9ZazCIOSWSgnq
S0sYqVRWpUs0SbqSqMd94vXfmfFJBICaEcpS+X0WBgcav0rOkUWlJyCSnxTiqy/2
7PbVkCx+Kn6Xh9N2q7qknqQ/Pvu8rX4/OHiQ1mDIr2EAM1zDAKyxheOYfafc+gva
GJk4zYpKcTnuQHyxd/u1vmoziVkcrFX3uFxvDYefcfcUNZh6qOUfhPQMxjKoEzUR
QHOq2eN2b18YcqxLeqtyQJxm0qNJxhXWJ32s7299sh3E4kNYpggMwh7Ss2kLFJWq
vwWccvtcUlIhJAoXpBEoEVt9R6BI8BaNw4ihTmu31o0JyZeYACzFHWG3E0neiNtz
BZLK5Es8YjCXgtp9eLHJeewf3qsqpPdyYYYc+XA1r2SEB5Bmyc9YlK+o/cPH4Lx6
mH77qrhwP2NxhodTMgPWG1sRkMLdeoI8CdHG87Lhgdn4RvfMXSdiNr5HeambXSAX
fO4jjzBUWYqrEKeQAjtiWhJ6MLatqdyXzbQI69gbARADhiaQXanmX5M/dB1mrEWW
+UpVp168a8v+rEMGCuKaODO5eSq/h6iNmk0W+5Hi3wJdbxYOkgT+lgCxffP6aj9w
UqSTVvTWT0w/iUgcLUy/uNj/mvspB1NxMo0ZtqeVl950SBedlYrYloftJ2RDAsbA
hCzVUG5uz0GeMZB435LSWRbamJADzytP8F1E8GJSce3fxRCOzE9T12OlvQ2ydgXq
BY67faVEJ6CTmX53lwK/lXqs7BkQjwnjI2BVoP2SXeBLFsHQ7w5B+nBoTf3a/IHq
wpuofhLefcGgwn4akcnvjw0+MyT/Ne8ibaV6b0rdwT6JmWUE17Jk12lud2X0vnal
BQQ0jg/r2ztE51aIM26Ng/glui5NBPhe20N1kYBkedM00QTWRQbCJtgrgGs8/Z9A
kluWy3A6/lUKVWfjwp6yLaSz/M3Ri5Hho1QnJ26w+yGa3y+T6FD0tK5dvZhKd394
9HH8mgHf/i+e/k4pJyRjDw77+rMJQ0u5fR0MFikyOmd5rxUbZ+MwitfB6MrA12fj
QdnmEI0lMWmH/DOMh/ZfN/cB88PA6pN8f/6go9qnhXtaQpvaBWdvI3xPB0IWFcuG
q8wGrQJOvjqrga/EE4YlGHyj9ON2vaRuJOQtfparxDdM/muforjLHBjuejepy/4r
m0A5pCbQJIXDgmRXSR6KZ67fpisEUahHt7qJw6Mq63ViFGeIkiBigCr3g3vctfit
D/xTH59+4sP/w3UWuKT6NkBHIJK8cwCZUtES+3MLWB+0U6MZdTh8M4W575z8OCfG
VL0XPHwBmP6avBHw8dmcCBVr6YdFpQGkZfjPqReOz1tzktWl1jwvKHO8HUMxxQqL
lIkaw14LMflpfgswhgHA/rUxhjKvXGJWm0SA/IoiPFSDMUZ2hRmbNyOpZIomz9u3
80cRryZuLJSgPW/cnjoSROMUu6ly6kquY0C3HnhMBQJV285LpBu6/RcjSjVo7kuw
RWmJQfEudnPi6D0d725B5HDZZb/8fL0pybh083DHXY17w8ugbFe6cBYaXQpzX7HY
EAquZzTFyyoeItbmMuSPX3Vam7NUDeFr0jck2Pm6NMAtC8m33jXk4ZUnB/YY4B1N
wN9sEFF/FbOAp2pzRGEOCKxaphb+GsrZPRsSRgNmbr2XYmsaXifO3lW9HKahOOHE
uDuNoUrel0TJwlQGnLBq+SpSJno01dIogEmgdNptuAA05/6rLmWwc/a0LaRzQVnO
vOPuTzgt7G56SCEvtKZ1F3hcKx1m79npvp6nZ6XVT7KbBkp8QstJ04ymA5WJAoox
qtWwYtWFqJb5WD3qbvWstrg9q0mwXsrrt2kpR/BeU8VgnAie1AFp5j+7v21yB3b+
OdBTPz6n9AEU192Rs9w8c0zS2jfGQ86tfGOk4L5a4Y+0GQ2UE6mkgLL9nIlpKI1q
AaWrD7yr0t6Tct4e9Ml0hlB0ofF8XWjaqBehDPceXMgC5RwGtl54zOQNfmwXq6QP
F33F6eqopZqBNBRgsnMGRxgWPgHqevvdJajBAwFBVVw13dXjYhkGXnRT5jsqwqbX
U7OQQda6QuY7CrZc5GRvW6BLeM1THUuOxdfD3SGEBAeaJ/fnlZTU6Hwg8480qfqN
ELKbiKHsCdeAxhV+Yi5Ric6rP4CxBnxP7I+MUgv9WsnLyBDFlrWajRforOkNu9ik
UqPOu+ZhlhZosLBvYJ3ctRfojE3G6iGYxo+RL9AMNld0yPO/RnCJJz5jsCAjWw9h
V6WBoMa2MWyMyBH8oew2bfxzpO5MzvMscqIcJOU3HGKv9z+sw6+/NUMScOxtIw2f
nLXPNaTY+KIHhyJofF4RM3w4GgHhDZQgZwMK5hyHig5f/1yGJ0HTyVzUh9X7wZk/
vCx+dMkrJ9ApyFj5ql06uw66BH5MYNNWcKY6t39kOnWHrnv2XY1G1aOGnx/iKY0q
ptLy/ouTrTDfjh8RFDnXZ+LqYukmRn+vZLBFPW25nXLEhnqhoRoB2KIshIGr0rTd
UQZJ4p48qFXm7ivz1rMLBWIyFWj+UMgZrwi58hgse0udDOo1O+iBPAC5PDnm8vZ7
J4Gdb3siBfPJqh7y+jANZMVb8Mjn69D/u9dEkOU+6aA8JCIwy0BoNnLXZojxtclj
kbJ/kmLe+IKenhjjwlvjQ9yNWbkkFYxKwbHauqP0DcKbtB8DbI3rR7sr+eydhcjM
lCe1jsqfE2DRFxV811/8HqwAaKEnF43uzBXxcvb5HHRc2i3yJV5zt7my+sqYHK5Y
wMsxA3Tv/QWXZFQ6JJ3mo8QqkeZN14m0s9zoEl58ZiHwHLj7YjTFKmLn3ecL4N7s
+yMhnrnKY74yCk1G6GuA/H4zgHjUizfEJdniko84O3VAlWCBHhfHCfvlSHgY+Y6m
3MbqaDIDhctOpVbTTqSGmacB+ag1wQo98UOK84klvElIj/xloUbUy0chdbxUwnGA
NX/CkgBuJ15Dc7tIVfNKWS0GCWT99MahZjrmovQCI6o=
`pragma protect end_protected
