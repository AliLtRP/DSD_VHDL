// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
qIL9RxrDG7ULKGX/GO0QC0CLqa2q2ij1F+UdaJdSiXrwNtkaZjUIsfoc5dBot3G2db2miGBmd5qf
tPWDnzdqYC9QS7B/5GS26lnDD6Lx26aJpb/75/hLtQ+85VwuXD6VCey2gGQjw+IfJ8dZcI1w9kxX
0B/PYNA1HzBhBdlIm2UPd5OSzwQvTlgQ/wA8dWT0Z3OoGkuiZKN+ZqQ/tnFYJCbt5tFM8MxS+Pyq
Td4CfJf7WbbGL2sz3ZmH2WfsXoIUXwSlkeK4TxsOcsVJlmb89GOOXgvtxUP63vQkY6LSeJA7J4vQ
mfqjP+ueqa9U/BTw/k3VmBzLC8fIvZL8zIE1Ug==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
05zCLV9LYAflkiKyEe5wkEc/KYvIls0be5hXe+ZAr0rsxW6EQ51PidcuTSLpXzcjw6oFmJvTkWaG
E4bUW1Hm9KfrbMVZk+STTvvPdmXTXE54kvuyaobayvxBZasQisf5dJ0IWM+pMSkg+ATkm5UWMAm/
OrzD+o2zLNDtziObg3koNInxqMaDWt1tGovhCjv7uRXlkSTL79HIOsN6xVayuKBoHLdSBm0iG0DU
YspwSXy1Hx+S4Or5TDYaViLFRxN8kDoHmypB8ghOhXU7LXaBmyI+BNGRQfBYMbSyxgSjsfXVpIEf
cBx/MtrwW1CrskEun/8j3rCRYfXa2hAq9oawPzP3f0eDH05ie6WJNm8Gm1uy2mDQfkaRji7Z/YmC
hvlXKh6OLSXyGzjP5qS8CfmzTKFY9Ol1DtPEXeE25kAA//2OYxyRZuL7UOXLeHeNRQJQG4+G3ltM
rNgv2LLIbMBOI52EeC1/jqR5DI0ToYQfy0mhIq3qOO7E/rLi4X5rsVi/bz0m0VcgToeHx46zHt7U
iyb1I7gexD/9x8skutrnRwTXCGEaoTyWxoDFh6d516gvEtew6p1oLtUkGGfOlJ/AxU+zNfC10rnD
Ws3yUrKzvTqZOX0SGY7wxYvMOx2ux5PYpjXzfQaHa4XQ3h6+LoQKBeSUT6+n2vSbZiHU7VCaJRqs
KC5lkocYkna8ZiA8AqQc2QsjHct4hbyyn6R9KBb2ddaliZDag7m3s0+aS5Zxp+5LAZGMG000eoiE
jWeJ1A8EiFcejbxHn8p/v5pc1LjBLxI4dSSHJ9AgEULby8uOSz6f6ezoXfTUvMoYCtr2vYbuncjq
79d3QiAAt5RMdlVEZXX9CqiUMHkD2FFfS7lR3NF89YOu0jN/wBBbApw9jhRFIXbV1+lzaKxxVBtF
T0l5Q710QkD5qnCAK+jYle1cxwND9jb/O/SFAHqfm3K0yEaYdPV1V6QOEiP9zvTtV8MVOpx5WjIt
PYyoMf0SMwPih/00mn66GoJNg19O6+pKnzwcWl1WQPUyDWb7x8jyW3GciAYMm8J0tt1GrLu3D2BL
a2Hmk4XvI4i4+myp2o3X0eVhv/prnX0EHy1UZYx4NPIwwyWn+nyd+VmIxECkQ3F67YVuf/ORYUfl
2yW4jpdtxEuGMLI0Ro2Ur7xwaxdx1azS5hv1iinWOH3HAAGJ//Ro1pFGYQouYkDDgDRMohi0kqoi
0+uoKZGtKEk4ygXaSXgMJ+AxR3shFCVcyBouMbvWE9uH4FHWolQexFxI0vuqne5vWprNvmI7eObW
pmtO5PsDcLdH8hudgOUbMHYdm3tXg3LZFCjBmIBJIiImeZJDBWOmHOC+DKoT/PAvOlbP8TTzocs/
kNft6pkI2aEJJ5spV5khYsmww/JgfOJZW21Pumo1irfpZIbkPoJNV2oys0RpTQr5Fs0tBq1jA4oS
1s3ZRo0MqWksx7gLeOuig0bLspL94jaeCqNjn7clXt8NASAfMulIAq9q0Vzt0QS0E+mCaUs0526d
RqA23L7Fxm9y8Y4vUz7Bh6NTazMprsqeXG67nirxd+79upsvut+J5Jswlb0Lakn4w4UCyDXB5lf4
0BP3vjwyt1TNJT+XY1Bq0Fz416ZD6RW7FT+CiXglO+GY/rFp8QDpVY+Ux9rnhpN0Xu1xey8L1ZEy
wfYMQXwYv+mjfdn8SOnjn3djdQnr0BUkph5mZrxPVD/2UPtab3AG8WKbhLIzzaU8iCoChVUuBG3J
S0wxc+yZoC2Lxh1LzgzTtTlqEWT9cAJpFUOuuKZg5uNh29P053n1HBHl1+YlPKDLtgjlAM0sqoqx
PWcepppkJ9eDEENV6f+IvS/kJdqJLFcYdGFRZ6YITLXVNRKK9DnbVHxoJ1V8e57Ph5AFgX0SjYTO
zyFlyfMsZNn+4VfJXBoU0RiaRkTKva934goSFtaQ2OplMTmvdtwS30sX4GcNRRFqAP1Zg660Udnc
obwFG+OcbnuGHmqaj0S+lmTAjiQx/Z35joTgKv+WNK4j1cPI4ZXRkbOYls5ZUjXszcYhZdMpv+Dj
vabCKdA3r/xJOCynLsplN+peQa5mujJb2d6r91YnU62N0+pt5YRdgktqDlPLrhfCsipK9uzYmiWH
cR/byl6HoIgw99nGkRCZvYzfz7X0UooXtfSox+kO7F/kwU5XjOG0i2nt4Wc6FKuGik9VvO1yKjsc
9hvLtK9dZdayoye4JYxeitaBQAFyHxhZZ5BZTDwjY5Vmr/tDY1Ql0MpPc+SW7fITVnnXDpNs3Ily
W+s92R61E5L7HCudAxjU/WdL+TkqTiQgLD3lfMG7HTmXyFMGjli1AnkUvyS/3STuNNk43RRib5LC
4AGvb2QsqpTyTieqDfRVDxrwAJb12dMHSRUETHUg8m05cleVaG0B49na3c1nAaWTDYwM8eVNfBNm
FipVs8MUrjaG88h08VS0BJWw4KAkunEnnvMbZRfWfosc42BPgWdp/bdeehgilQD5oftCGq74nTk4
L0vsMYBGZLFzWmmefmRK50wpP6cLvKqPCyFL3yDj081ECqqoyx4CCHhrlukPTFstFYY72oQQwWRJ
30FZV+VjaFJ3bh5fo37CUNGJU1HrpRXzqX4NkL2L7SitkFX6yPI/A9iJBg8ofmGOPiFQCxvsH3xF
1bd6cHPjWMpy6XKOIwEofyQBnnU3NhQIhDL/HDRQqXF/BrPg3lSSnX7rIUlPFT4xaJFIDP4PVuu0
CYKnLhMeC5LSQYC39QKCtjXicQJqq6kJ2D31FuDH6jK2Uj1LeJCEnQATXcjk8ciq04N4593Zim7A
PokS7kCQA9zHmqdQsnDqONXa9pzU3jO2t2HswLJUhCzKynWOuau3HzbEIYvx/3FC8FUCo8gaC20a
4WZF49B6HZyekxrYvSIG1q9q3e62GAawJsCE9nXH+HE1vkP9rryJANZcoSSL8cHHGs62CKPSxjtW
pH4WRziJSe7+HVTRbSl+mxtsb2pq9MlW+zuU7U3d1ufV9g3JzdtZpcWsVa0PZu2+b/E5zvIGbkAS
fhAfefM3IrkWm5CPcBsc2/i8MhtBskZlO0VLkyQK87s4HO9rgRo+ULIt9s8DiJBfvyt30b2E+idL
ZgyTtTH8Py/BJ99ewyr26dUUWTSH+z7BgxT8I/wwr3FHGV7tL6eNK8yJyan2Y8GYiRrDWZnFSLJn
DHJQmdKcborKUqjuyACZEpsZDA25MwidupD24zC70tVczX+2W/+SrVVrJVeuXtPZTGR1/oXUkGY2
vXIYPH0I9x5VeG+/d76EVYfazQ0eAXimmvnD/Sig8wIpHR53fY4Ll36MyEQlH+XY8fqRKe4m4YoM
V7MUo5rZcijuNzzdPQuDpq2vwB1e8C8RWtn4tgvMCmz5ZZiWOq0ZRLOMuKtbW/LPAYhFAq50CfPI
Wrt3RvZwQW5wTh+RL+Cs7p9e7KJHm09QXHxzkq957FJs85u8T8cwyWLObh80XzeivQVw16/t6WQK
4s22IHBQuAyHC7gM+ev66FKnh9/KQh4C5QeyqRCIQdJc0Xl+9DJGyYVtMARvVY9oFzPbjrh2UXLe
0skLZLMoXnxfoBO6tc1RMaoBAVSb2sVmRAkp6NWNEI+w93BaO9merHhn2nc0H5Q8W9MzmBiQK7dv
yXw/BqDq+1sIEQNStQHu02N2gpQ1/J0BqCivp9UylbVFXL0jIDQIfK1fE8xDBvcP5HqdpjwsUcwm
1wq8V4a9GOGhO43EJ+bx0pacZmnjGTBebFDA0WbeCDlExpUUJcrhLaB4ZvR/0B7ER/pmybdpKYwF
WYdhHPv/x6uLnnpqOsm2e2aZCalClDziWkOuZS1VFfyehn3u+WBh2akDU82E4XFHyghmrhJlI2DW
EKy1kXOrebINyjLKnSQLOerW0V1oerzxTxTcHwPbrVCmo/3V70TyI9QbPyEMrIfnShF6aD6zaE3f
SemV59iKPfwyvQWiGE4BiWE7yv4l1GczvHFe/W11EanQI+/Oigxw+84fZEvT8WCb+vYor4I6m6Av
9bnOmWjJihgTfXlTlai7pU7NYhRQFsSFMMj2na5DeFg6T0MhsYCRuCvKT/yUEkzduthp+oMxSA6B
NZos86roSMN+YXdWTP6fBpxM4jZwECs9ynfgBkmni9xP0avZ548UYMWhmdDNO3bHTCfcgdB7Sxlw
oSWg6OyNEyGUKOzf00CeI1iyS/s6+fAUs5W4WLMXP3xlwB5YiY2OTvpsf/fGRlV2ovl32hE1Wo9w
OBob/00PN10BjkLsEQZGrAYbMT7sXx2v0CW7HxtdE+fULsyD64pMLmVxjhrQkbAU6340SNtQOPTB
749dTOcQStL3kXWGf3BiiUM54yYbUvjPJ4M7/WC6nYvl1LRd39UU/AcukN9MWvY3D+qjZ6ojrSIs
U3TL+p7kklV5euZW2tzpmd4znZIRyFFSw3nbJCmAjHmAfT8IZEW9rqOfT42MnMOuSv8yljg7uR+O
AW7Wgq+cxiALJ5HTlq8clOWW5TMFzKGukm2BRDOjsbjQJNu9lJbhvmeYnH/AcF8Vhwh5eqLtDIsq
nCN9BtkP7c6hUdPwLeKxAmsaAEooj79lcjQTJ/7taGwtlzo8JqGUtci6gW0alXLwuPI9bUsJo4Bd
Qa//chZ0LpYtAsKsn0sfalXcuhqcZtHuKund5EO1Di0XtyjALnB93EocfUf4vlzF/ZhSj4Y59uqM
jNW0JrBBJrch2Mp58fTrQ1uMDCPZmOqE/+WsBUrq8QDX4AWKjKEN8jHdM+SPOsmklyM2aVCmTG5r
GnLgDbtmI846gWae5R+/hxhouwDGJrd5eJeTFmAKMC4fnGtPO7o3+4bOfCuDqdrk8fbK0pxL0dNb
RV/dch+jmgwVApDQzF9pXLJrW8tMeF3kWVJUhykIVGPLKtHqDVTc0iqzZ91hnUJD5s3rTwPW00h7
AFQVBF/IA7CL1A89vfPP1XVo6LmIa7QQn0ab6hPPzqLs2+MWjNVg4cIGWkUqDuBsfpZvXy2G5dnb
dmsc5DUlI3Mz2efObzfNSfDdDBaowGJRZ5OVQLQAVoHO7yEfRA6G9EMAeMuO9/thaWvoE0/34Cjp
p86/JeCQV9JGxKqkkvvyHpXlDfpEeGAsUBGsx7vV/tn+7yetCkDaglvnmWhzfleFdZQ2aDaiVgpX
mNzpPy15kUpS/ibMO37U11eitELpv8aLSZIvIGhxGCGE+3SBzhoNwPXpoc2eq7HYiGhz+he4nC9f
xIVAM8/4CmzRlm5Z927qDNxT5+4qUKtPaNGQbTdaZLPDYVdtCLtrj84DpsmyYhxboDIx2CcZtjfw
opWsFjHtLIzKEd30SZpdUMcyVrT7sjMcBL3m8OFL6GU1FueSyDhjHkRKLLxn8Pi8atOiOU0QQkFq
IgNhg1Q4NhHHVYHkkad1Fe9zT5Lrp8MAxlSiiW5iTZPIxVBvrMcQhqyfDToIc66y6EQujMpHxjt5
dE/BVpkTWLeHsNVStGStanKy+VxC1FwhktIMZvVofNT6JmIL9pKLo1M1+Nvnd6QIjqjdJw+hf0bq
W2GwhxbKz7ZEdkFycyTCiXL1XZzNDAK5VuxBUBoWhH4uo+LkAnGIKQf+Xgrv7PM+QkM1R12LPV9t
35T/1SCZR0ceWytyLLvgwQzs3aphYEMN9BvyzS4lKsBf2BiTMKY+CXqHOHFD5y+wZJ8DDBb8ffH2
+C1YgMdVw0GHn7+ESdedw6S4IwTflQC4sndR6iSNKanQTt6ALLYEc0yHMC7KrH0VeOVymqm9Mx1Q
XO5Yww==
`pragma protect end_protected
