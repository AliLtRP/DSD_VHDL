// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:19 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
biUOipx8JkaZy8bA6NEnugQBjAbgX57UvgbVveAwzydZH2lS18z3PmRNTYvkTcta
j/kb06ZkCxhEVoPHCOYakOb24LcC8ajDN09Hm9lHHwO2W0StvI9wJC9ROn7noSjB
wgT+ikBsoE/UT3tUK7wuquUJMPa7iY1H3IKwdxpZoCk=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 42064)
ZcnqM6Is2fTDCzxWUQP2e6gEg+Ym2quORdtXrpgBpJ6mEinCL/UcPMBQMT1ZdpGd
OP3/5gYjLb2T94Mse443cuIc9Mw9kMmlUc9qmMffbUZY9eQvhCnvyPCved3t/5sd
+DWA9XMLvOaBnqBuNNWpX6xjbSB4yUBh8wKQ6P7jvkta5zObgn7cxmCjO2E+GRAH
Nm47qMTgupLcnIDZXgKhI2INyHb9YnGooiHieyLSukhIuidrIjr9bMG6VJKAB4IB
mAXemektLLtf6fwVepojC6ZiuiqSKftUVQxg6PHGC3jBYwUFLAQl99GRCEezRgYp
08jkcPnKNFUCm93Oh6NYK4JvPL0a4/P6Uz8zZ2vfD9TaA0pZNDVoaHRfLfB64lVR
KU4+8ugq9azoBnovTTdXoIwE2mLx4GEjRLGpdyDBGa7jFpdg+sJegbf9HEs7sy65
LWCq/plP6dj8GWwsRCy3sfJo+lgH77JWyEVAJywy2sAc0rg8q2Tf8DkblyfcJKX/
4Waw+kArXo29hQUewZPkihCIlxCzICwDtKvljeqp60xwJm2oPUDA5i4KJRGPNhFz
o1jJYgTBX71hdw05DwYH+hbhMyYumrZ8Ht619VAxHZr9ED8CmeYgQO+J5Z6t2VWZ
UCK8jhFO425P2dNA8BjykzhbKcRayGcm7JLyEKyMHx/Yj4DVyyjduldAwtO1H2uV
MGWt+dH0ucvSGlm3FOiuyrM3ZXWQz7O3fIoGdtZBFbJB1Ayo2g2KdnulK53ZtIjS
U/2ebF6bM4ZTwvbVq8iBfQfAOA0MyE5DLFtYabwvDwluWnQjeBdn54s1Htz3V2ef
qulInvkJqA9cppGr/zesYpg4JTwk8Zo0O2kz9Ho+90bBlepjvef/KCZ9B4TFcQgM
EH/YoVXheITMd/SG1kDfzKb9VpgW10BIMZT/F0i893MOG3DHnkdWHPi/UnRQ7pUs
aguDKXvu+5ab0mNY2mn6n//cYP91N+7ZnosoIQq3YW//jHzxFBNBvuleVF+1Tf+n
FtjTSYeECifMKPAYycdgAKfysGX2BzhaJB4NZ+IUQy62+JKdBfAuB+Ia9T2n/KjC
HbwKpS9JvpAxbivLyg+6vYR++xVdQ2rOqBfgGwUo5q0f4DRIa/Juip9g9og7mahe
neb+QjICBYkFOOd5cgOYSAi8v5rfjSJlKUFC+gZMc+O6/VJ5maS/3Pv3QP7cOWPE
kvAbXQIlK7nWNbhTCNVIlOI4ZwAx+02Xo0zk6tfEOfV29CMQj/WTZY3OWt28Omjm
v5ItKi2c0Bp9IMCxSBRzyNN3HcJ29lBy4MgFB7lzZCbpiuNlOqnfxEpHIXw8SxRI
M4vb8sVrnzxnR72yfNwfQOPAK2Atsq8jk85YMVXRLDF0i4nDJ2X3mgIEEgyXL+l3
es83DDM3/xxwx0OdDhnQoaRiILrzkjXzNR/DJpCRFJafO9/lZnAhVulaEwtVY81i
DR+1g2o9W/gJIqbOL/fczECPsT71+G/96H5rXDlHwLx1dt4iAXpPTX+OzdTC1F+Q
e/8lcNJ8e6gROM9yNbfhd3oaR+Hm01HXcV+6dOcMhYUE/6plM6fgj+tz8Mi+gqff
Sbsw0GkC1mr1kx4HoixwvPN5tefxxPyK+jZ3ZG4gDxDznJl+/caJIu0B1dGFDHZi
q4NFEmYOSheRVwj0YQcxITVPatYRaa1/K4quvBWPxaIGLMuLJ6JL1yg73DN+YD+W
00iKXgiXLGA1qb0MqxW/T8RLctAxCUkEM/Nn7SOyIvWv24SuRe/fvS8NNJ5PWBZA
YaWLWMdPtxU3cp2YVzolHpivEOfBcFo0GiR0Bah3/RSRiisnrEIyOIYRb0x+3JLB
XSZ+/t+E5AKM7g4Dc3jpTzFFgDwAFY8wjpuCJwyXuKK4maKjzY9hhyWaj8MXxTFr
Q71LqOEG3SYe7D5PCxopP/ORrGlUhOBM36e9az86dkRdOhA5MahZ2VyC5W0AIZ2U
3vS97nD4qtWZZGH82L3ImVjBpctSjqu9VnUW1uazCdiK2alSCrauUT/QAb8CFWQo
zLmNEP+j97+H0nrLmiW2sy/1YCCupLrB5/uOJ0BFBMFF0CtJ2fbkAYzyQdSIVSit
GPOI5825DwJspfuiV8ogsFCdW6Q9l5otFi8dTXPS2XuhFyKzk1vlnHm3BD1VGf/N
XZrS2NWFQcGJScX1u8hEgXRd+WrcNC3NBTuAaRIQyqM1m70WIrLfb8j8GvZa849m
uTRpZtBnzySfYqnL+VbF0KVCyiNCGTb9USnuF2z0gqSo32S42iIR83rJuGPRZziw
OrsHr9USpeOAh0EF2x2jmxLIhJohQcBi0fGX8YAEFPcMkQPnzdYHBOs25cNtevyz
tAL406L9sNsce3UJeAYiZiSGC9u6FOAIXpIvsu2y04zXzgJ84VEiDw/ONbCCO8Ny
Fu+NOFgty8XlXAfRId8pBcRhDcXVo8wWxkTGXb8f1xcSeKK+8UgpZf0/jzywpVF6
B1jZAXwCh2njH5WajS9tD8n3CdiNeLVV1I3uKHBEHNFgJmvorVVXL0woB/EtBO2B
xCyZ0kyqwXDGhrRDxFQ5WM1lOc/aRKbKp29WrA8BxK1es/KVk0D6awMqb+DW2wiT
49gLoWxcsAxnit0Qq2JHE6sIp3ZMnr0Rfurleg+vfTEhG1bGDI+h/a3Ovhhp6WXD
zE1nS4sjVslcXxKdToTMnPxTUQUVS6sDGdLy+q7XPFaHrN8ZF7qaGaWB25u3ogvY
qyaJKdO/t5tFS0bpjYJ5t+4N773A69t7lyEaPlu0Wj4waybpiHGjqZu6Pn6u4yep
MLwiEf5zQQXwrPL1IY+H9XYKId2lWK55+CnAFxr9Iv97tFVF1sXlpNH/go+NSQux
tyw+mitAR+aDvuFBMxnotbFc2Fvw+Sk5GADoQ7JpvgH1TMpGh0WI+zZImWgrP+9U
DfKBYTdDsxChi+fyIqYBR08bBVxvAEnztYRNaMhX2fDGnBy++fL+DUy8OJX4BVLe
oPtYtJWeXBd4l3vnoDxvigvji0cvFGIad3E2lyHhHmpUv399JCtbsDTRv+ZVyJe8
UArOhiHrYv0BHzOV2K4Hb/H5gxZe5zIh6s+0k3ThjgTEd1Rn4/Geptlf+NMc6CFZ
YiPTod/XHC1/RiMqeHk4J6kFhHbagvcRE5I+leKnFn2CxTUy8w9CbAdDqcYU/Jpo
39EjucWe2s8mvrwCb4kHDQ35S1ximPhzPWmjBplU+Z6kAwklFQcGFjRAJnqQLZgH
hd9BOgkVzV5/cCNHlKFbY7cD5rGPDVmTBwaiXFQnRdk8TpJIe5VTlbXcl+rqZ57D
SvrZEG8qes7tYnmuVFnFVSAb8zjzKPYTRPWCriIIOsnlLjhue3oniYp2CtGn0ENm
P8pLWiIFJ2kBM2vtk+D6/GFDXeoOzIL/b//77UmGJhWweP8/q34jtT0Yqst7A58C
HZf1TQ1Z4Tcp6mkYnY8RyqgQIsLvjpiJ1M/Fdy7CcMD0Tmgo4VCVm5Vw5O6NKJtn
z19a4Q1lgF/0UrQudRgi6z/gtwrqNrVv7lBtlXtS3uuIDQ3AK6FrQ20L1LEJKRfe
OQZdQUqBp/bmPClT8tTGgphmel6rR1OYVQctYnWk7RCmiGYHCQTpQR8x47iRWBFB
yhjCd/c83DLkHhQA2CTLEEmqKePvVrq2bHxnBeBe85sdos2Zl+6/yUgfVvh2/nCm
Yh79uhj+qNRXDrvAankcxGKvvENQr5VJ2cV5q2MYz/zggIL0Xu6ajNyyZ0/CoRmY
0Py3M8X2/mhu8Af64VwteMxPaHfCuQqK9WFFhB+K601RwPOmeuTZJiuVokeaUlkU
x/dwFU7jVONFkbfxq3TT1tWZtIgcsx/nOT5+3Z3XP7Yb8TGWYyM8E4cLSAl+LOCc
kqHabWoFO0ckp1z4VT8fL6WTJ4CXMG4LxF5UBFtp9j+9g8ven+wbKgrEEZZe7TPV
PqoegQ8kjNm9+hn8x2uGn+2a3UeAU17DWK0uwIPMf4XPespKpaSrATCzaby0sv0v
vETV95MjfrG/jZh6nW0Em9LJcuhgCRS/35sU+5A6oke6VTnUZM8x6tJB2NZHa81i
yc5B4TMrmeKGvaDOCYDCm8HCelJK8ALWL0com3WXF4Yxwfm4ZfBIbzWEV7A3qEud
vIsJ+SUgjqtYTVQBunQ5uKpFSEa6KS9zMEXZZlVCGZdznIPrAVM4zy0t7SfajR/e
9f7qREg9OtlPZ9bPsnL4fLAhWm6ApkTSDZe4eqd/D1H07ubhDNEg+UwHMXDR0kjL
zp28HWfpRcE+6hnTq+/SB0TQ0LHedUlCpuXLufPSQhE7S4+0Vy8t6pAHurIDMQ8X
Yn4HfxafiR0tx0etoS3RC3MsvOPtBxdDAB6CMqwVXDDanHGNZaNmc4tOvxaielcC
qckr5IJlCrKEBcj/G7MLoBktxz+o2CHwF2MzNbHqAc1bE9MkKEQqs4UTJ4MfOCy3
nqpx9IESylffcnPXgkHlNnEGgRGf1ZaQzpU3Nz66ux1KQUb5KbLXqi3muS8wQ8Eq
Q/lSgjP+ug8aSMvDWlM887cWKDTcg8L39KsWKVClSgWL1A7ci9qUbq2KAIQFwC8J
l5r10UZX0A6UYfJfGyA9RmgW6KvaAo7siintnnjUIoxSlkWM9cKeD7ygVXvhIprs
Biw+HTRROQG7PxblPdP86pn5c+c2BaZ+u4cp8KtbdqB2JV3qgDGkQ6IvddCG+MR6
bhSv+nxy3TourMrbbBAaTzlx1s3e6Zulzm3B+Ors8IrwN2a7OMi3wq1i4K8rmjv0
Awx7Cf+y+01g2533WfdH0j3ah20zWlc+cBcO8BDkP+VRj3qBIhas43AxMvEf/2Ba
sMOAJgD44FarXqlzuzg7prFF3xvGe1IyF4oqBuZOxf2FxdYpTqgwEQo9s92K2kNu
u5RXEBK2bOtv800XOx0dtLIaDrOnQgC+SWW4gjEH5du6RpSNGtIgNoSe6CvnWnjm
ItwiHlQ3xSsPXwaP3Gl/j+hyJsLra7ypF2iooy2r+9xOn40yDhiBr7rql63rlIDl
fnRlAWFbKzKOYjggMc3baXVGkC0L/SvPzxkUC6zoTWFtvp9N+C6PkFzRwtxluCQ4
I6zSQ6dIkQabMXZpCym5DhX459TLbE48R7X+ZpWhtJw5ts5hDtlUo8Ir8LUpy8b2
h1zv7dJJbuDTYMMoKJMgB0QJES4CuNVteUVD8kmwNVQDSh3ATYDP8pt+kOq4lYSO
8kZVoDiOo4E7oA+qcoOKnSSozvioVjwT2EVZ329leq6xvlm0fM5D0upkTKzHZ1wp
3BkaMZ9QOzoDCSV+5AKWsLU+sWAAVRTF7MQya4+LLsOv0ZAWCK6EV/dbq/2wSFsV
BmFB67qrcLqIBTdvzWf2NxnMSqg8B6kejZgvAQxxz6QcImHQ/twTVbTltt3rRhbr
LIon3sdXRdqHk+6X2qAPS6qbIcctwZS6iK/Ny/IVm+RtPCUkfqco03J2mvBq9qw3
x2UHT1WnopxbwmhgZW0Sw5QkU2MP5FC0/yXzN+0aat4eyPFyowQUJXUrmLkKiyHY
87n8nxF8RHD3rqvncBMvi+dCoznuQa5Wy+9LGTEx4ROlKHgtT7l31v15n0/5PANF
hzs805vLuxfw1Ww75sHOZ4WyP5zRKPcAZRnactk1zMcrFpwV5054hHKjUE6H37aO
eLce6p4RPjqsulh72klbHfD4CUzTEhcngkB2NcS6VMwPolY1C87Z7d4E9iJbyJE8
Dhsn8tP+Tb7hEfaTw7Zl2c4Bt74BQLUIyW7+1lvBztHIns9bjEokiaRC17HMADnb
QM3JrX7u9jB7033ams0VVMAs+2SUM7Eqxde+G6Y8kzWoGLXSyYmhTvWVME3W1ves
JcvSpKGzdi1rtR7uMoPU+OXhPdZReBw0aw2L6gIX30eJbSFUHCGZ6dE7wCsBjrZB
qx6/lYKhbrq5QhjX89HgkRPHXNA3BZEOCytGRf3Hy9f43fR3yKTZVEa317CKwWiU
hgMWRSmCjkylTEx6jIKR3zjsntaPvhDfvoj6X6co3eCKt0UbxkHHvEfdkDIZHDQU
HIvIn2PVJhVmdSDQDkeOoPZUb5PRBlUEXKuPfNFHMfJ+Ng+EGGJ7PrgNwvQT4/c9
OVt9Enk+ttlcfjkRSfnbkqr1ZhldLYP476RjYm6lRQShOUosD1xGdiQA+Pp9C4ui
kr1ABkvH5vsJL1Np5x1ChxfOYw4S063f1M3YMUygUYQvt9knrFhyi3K5yiekRCqv
+vDdpcIN7I49e71rO5WpgJpP3DxwrKJIDoevdkS0fcEAGf35/p6Jo3euJ6pKBRJ+
tjBI2wRfu2Wgt4jHZqEAsk/gB+n5vKQlpZ0J/tzaLCyWP/jJgXxROwa0IlBVXTeH
/whQ3ocPhdKIVj35b1l2DMrOMbr29EtCkoE69Ufm/S4HA8WmjP2oBztDQh2i852A
gmhIbLPp3L3SIRkKr2kOUAmWFRP/4DFDCSDQwSU/wL1E+frLsmZVgrKwXm4XavD3
dYBkfPfWK27DNcYD8IoO4HTmYtHdlTyMo453IjK3iUagYEA5Y1rqbqT3h9f7FssD
gMwRYFwx156qjWbKGwFn3w8rSfWfhe+uN1O2q13PQsAv1GU2RH6gFQSrDyjziwu4
Q6DoMOWn57jf+zEjve+LaGN+tnM+GGsfmAcgFzQW2PtnzpAA2D991nJBvs0/6GZ8
F9VCMtmraedd+zsCdDugSMBdMc8PCYKyhHGpLfJ19fxLfMPlma1Vxp9KPwQUFYpi
FPltR/G8PffFypYH9ACQ3pUzxk85Fdy91pa0oW1dI4g6U9ZKvXdmywI0ozTU7Np1
9nHF9JeW95/Xj3Pl0K0CII8r+7mroEZo6MhI4btKOUB3e0Y5vC2B/AYfyULSy0Rt
oUhSqkNCZe22z4szNldlFNV5Rf2/qY6Tjb4A0tXy4LdGtVjwUUzhVp4S3fMbvVzo
p/j3vH591bdfPjvApxt0llgm0J8kx8RTKFAYC/6fKm5SSVT2VCbVPuxtObU/5cze
EgaXT4HKgiLEBEsLnwzCv121jksdNFurzHVPmDtFSq5bkj0k2rSTPZoFuXybv0aY
X4j19lQck7HnHLeyTPR5T1TlU8vByZlCPy3ldc+G6srT5qkEFIqBetDaiXRPGukt
DBJsvsjcyOjJhJRxSN4Xtr08QVKCJXuos3zq2CPW8NNbG4A1We2Gy0EBYDkXibYu
pxUYUfLuWPBw5XoaKaIp+m+4aswRDQa6JF6kR2w/f7AeWqCP4c9CPatanY0Ow4B+
JM6x2O993iwLygNDP3Z7cuixw3s1D5WydBLpBDOCnuwLQHx47ZcLh77S+7YMd+ci
XMtIXO6aHv4AmtPWYiZExExR9ExLU8xm7+/PzzaUnd43sM5BiXhXWOMU4zTH3V2j
V+QBBWMlLfsCIV8tWmHLTzkIzOUNOdhBmy3ydpVLVJyZJWv+dGIVN3eBXYm9I1HC
1ruiF/iLoWiWTqGA2JlIxfvKBASOp5M5yBlX2BQWGuolXtXgSTlgEN0k/MmkcEbd
vUlOwfx2MwjEcmgYNgsxDNN2Kfj2eF3D3WyE5xmc0oLWxuvMTSZwfp3c0F/FxPkI
EOsCu0fHfA23RLkQBJxZ2ILNG3PPnro2Hviuc1bRJFqx+9vHb6F0v2gVyXPA63nN
CHLS1zQrj2PODkTHQVabstYaGWj+t4mDTq2pDjjNdWjzlrkwWmOToT/T2OaJzyWs
EQoIF/gGg3bYaO01XH7nxRtYmF0KSZLy6az9q1ClKeoQQ28/W/KuFMycuiw38Xxu
Tbnv1qpFGhSq7h45IJ5JB1pnP6mIHToVspoxoSBfLx7SUJ34ehuCL09wmxEJ8ImK
NzSg4Q01ikEaeBJsPHFVF5iIUkyTMel2VtteflsDPYH3sxn6X73tlv0RDbyiKFG2
ozcB8A4LqGunZjBp2WXdMq0YRUOiuUObB2YJJYZDu1z3BMhxrjA+neG5sozXKgfK
8lTw2ivc7CddLFzn+dU/UhFmZvitRutTDYpsEGUKLvaYRvr48mUKjdDdB2NCOrWY
lGvFrm3uO9RZn8vRhrkvgZt7PEj3sKUWehJbd23bdgrjF8i/kpCY3MDt6aDvn73p
+NqIuFl+uZ2EJdnQIEwUkpw1qgbv8xtJTXFJrVzWxGjTO3KzwZ2B5krf/lNKG1oY
nQjA/DIrIf6FYeRImW5Hqmm07LhvLDFiY1WHgPfKzNl0QfCl/r5Fa52fkCl5llNz
5TF3mcToAEd8mweHmFD5iAtVZ/0nMn0JjY84yPuRHXGEAW/Aw5yhWxsf30y6ahBD
8R4Im+I3fjDK+gaSnF/Tif2MPDR3Jwj010mVvB5wrdADP99tgyPijYCmf+hlrXrr
9Ppvh7kdn0BLVwAavgS8z4DWIioxON4JMsRmpH6lBrW7wc2fsBq2nJ+P1DlG8/47
f4N2+Vc7cvPHbSIYCZ2LRjkJgBtKgStvFncS6vdIqkDQua8KuUZMRQ7n4hXisoPv
kVuhhvib0TAo6m8gUGiv2wP86vRDkIz36GTPEpySQxBy7J4lshspPg9iMNNQX5Wp
tSUG/T1BCUWzdwRinCYiSku/CPId6XJy9MrhjwZwwUfh7ocTIpdSnXlpGeeZoHY6
Xkdr3rAtpOFUX8elhPEXRH/qjVANBH01IkqV3ibmBHqoKpu3lR2R1UdkY+eOO7tx
1OEDTUIMrJeDFnNViyHAgjehtGcZUzpU1gqoo08MsrMWJYO19pg+ZKPSH5Vy0JhO
sW9+RaEO6YRgB8eruOv9NhlnKwgEJJhFL3vCPBx5KABf7UxsDvDa8KfFylqNcm7y
a+RJ6rSf8/KrfStZbmNDbDmM4xeQ7j/E1lMBUwQdWGX/0Hae/aPiHhlFUG9vYBFb
ko3bIHwrf3Q+B58mV7RbeXKs7zJfyvU9IawCBfyuFQYg5pZSlUaXUYYQg9El80on
lWsY31R9NWrpv+CXuweYPL0Huhg+j79ralDLGFIfYEDX3O30bO1LdqxZpTQ/8pkt
/3TNzHiF3KONhzWAL7icEtJkssBJhtpLMGY9juqXYyAkWStQyf1g+Jp66H5yqKbZ
erybMF8AQ5BHNAS5UO3vUT3GqhnaMMCrbyT/PZ2KfLnzc1O4nvsIChSaWTka54+r
gZKLbwiuhj3l4EQ6R57NlgwcfhTBTdA/DmCS3Y4aOIOnugiXVvsLAg/4QNVfVA5O
F52kxJPu2AfDs85IDVCFg57+szLDeIcYnm2uTOVZwCkzxPx65cz4y6+LgubJoq2t
oJjag9zTSz0Fh9t+TrY5o/Y+lseHmQ6bEVjalqzg3hFPPevxPyDnQ3feoX+MW1X0
8C30NENUhzhd41bfFkJJke1JR1JX1LM6KV3PPNJUztg3wPaI225T45TwzP4jsYag
Bqb8u9OQs64rvGqWTB/rsL35R3lduHImgm5jxtd3meyvlUVVFCrwL0VhoB5u1lJA
AaZAy1NS8VujXPJlQRX/xUUgIp7QRYhNsm6B5EVXwF9nuanDRyut8a6jmzu+7OQ6
fgSQnQrXxKi0peBGp5PJOpPy4xpgufUKOZYIhi1AOGUAuIMLjWQQChNvUpbIM/ML
X8JX7muxyCY3Sx77fw7mmR0dZ+3F2oopSdVVPMeJdQFJBDQu+ia9+MMGtTGZK+jS
oUb0BJ8AY8opbiLReWMQYfCfDwvoJ4wzDsfrO9KI2bQWyV375UWoBtNrj+HbB59+
NjmSKAVXUEklSVG0GYfoVJREROYiEq7Zy4349wxdomepaKVQ3RAkgaKvZThmbda3
ALUUJbnOoeer4JZI/GsB0RE/PN3mN8LfQfzn2qMbZmSzBEclCMFVOXgdA+702/TF
gA+7V9nJNKFGhA0TR3ak6X8+FMAxMcrKmyKThQBGvCoXIIWFc5gdbSjjHoG9/880
YVu3hJN9pwZHR1kIwy2HoHBG82Fy7HtHz1HtUeV7r1p24DG59mPYuNay3EfxRg+f
NNilsRGzVMEeJEF8ukbC54++8HnHUDm6Xs426Pj2ZPf8BvOWkj7IxHeeueJIf6lr
lv0SKHT71jbIciHF5BeWOz2uaxpLczRN7WlMYiZ92zuS75Tvd4MP3jL8xqSTZk/p
dROodwr7PnT/DR+lBJ3vo1Zb+/wullsbxwXbcWLGBZP4AiHvjl4tqfjNblw4srGy
iiqpHMOnW3iw97JSj/sMBt6je/74LnmR7xe2T8NX3tmgTBmye5fzlQLcqqBW9jmi
Evo1IQ9d93J1lTyRPp8owymrdY3Svd6bqGSOK4JDYMjlGNIagDLA+KsxuJx+8MnM
Hy+eubfUSieQsYsJ7cmHKCPBadcM06RZKA1PuQXcxdqGj+kQkJNkKFejwenS++1u
oJYAZsxG7oquTDgdGoOtTIKKu3yYtGML/wltmglrP+PCSSrTI0ASeFDzvGVTN3h0
zLhYutf5KFKNpzRahoxuJMn8Dq7yVoaN13aK+i1mIgApSXnDPC9PTaXocxQ7Dmbr
FF6wsadrGG1xiaJqeKokPceUfEK70/oSuoN0B56meKcdBrlbVc4K30x6Rm06YNNy
6XDAuUCEubjJjn2/PRFLpElsIAc6kESo86Qm+UAhFc4MhJnna8xy8ulJJWv1gG9e
TwSIpURxLLomGoH4OzL8JU1BKjbTLVJM8gY7Somi+7/39CPzFxhmbWKMZ3/BeY2n
nUnjAaPPoK8FYVD9YEu+YRM0u5ihuq3TpBX1QF1KGjo2MMhojVmX6pE7Dl/gi6gV
IIyscxWLttO8wR6N1p0VSypLM0re9GZY9NSeVh4vJ5zbl7H6osjz/jB7n/zU4RaB
gUDadXpM3SaEKbqOeKfuIq6KYgKKMICU85T9ZZ8RWX6PVcz8FDzrEY9mIn1ImUz0
H0JNLEAaxsmNiUw9Km8AUTXNGNuugVVVFhNcMGTsJ2+16AH9j+OQhKkvps4pWwb8
2CS/7qeN/AiMs46h9Q5ZUr2ZIs71XD69YHslCq5IdPc7v9DB2QNk21WqTVirQE+/
4P9YXaKJffcIexcWCaq3ZDgz80eEIbuXrcmBArqYx1m54jW8m/EBHQoP5ygHwQq3
r2w43EtoZ+vX7F29rXIXXDoNCed4vgfaWO3eXg7jCIjb/SacHR/GP8DwP4xlhgn0
X5MzCwCYHzT2djkyGroJSDPuuIIKjsPPebSdZLpIbfaEgsKl3qRypDwL66nFvxgq
nUM3P95qvaEpvjIqVYw7joRL7VWKjzgU8g2wyLD6TIaaMJ05tGN2EgUF2a+0EL5K
ETPg3MLr8xQD9CQ11P9jNOj3h1A0Bf3ASzusKN2JbLPg9/0v8rMdu2g7VWfXXXrW
0NEAh+U2WU/Ko5tYiTzo+tAL4kqlZUHuUOAgi7aQfBA1Z6jTiJSP25rbLzzDAucz
TkLi7eSmLjK8RoEmecG519WLQuGfeCT6r92Fc/7C7nfy8/MmWIyjAWtLXrqksOeK
JwiiPL5jTrbs617KABUt9Niwjy/DHwrH1Jkpc6ZKUCsIQuthSHhB4KKYXTu1KKyF
TBZK1zLIrf3Gpcg7pzg3fIEKs3uEa9dPUjWLZTKiWm3mnssGEGxSr/TB5KyeMkz7
h8WQBBvNLfABe7YL0lcQmtPUhaYFqtGZW4Hw8h8QjJif9bYQJU72PD4PBDQqjKXl
rxISz66HIV1eNASWks0z66ckVcGrHBGTEtVW4oZWlc9Kmo9aJeCrQq0zU59QR9WY
I4bzJarNaifKesd/bzCh7uPuYDfEcyXw9XvW2ZdOywr7ZZLBZ3vMovTSr9lXbjtk
eAtWAURaOJgiYy1ygWS49gkjQ22sP59bQoUkkVmdop8r8HC3L9444t+qdGvR1Ibw
IiFlDyFJ4+b+Sfj0Yyt3MP10Bu6hvG1pLV0ZNUT/55SLF9jUfPY80rAjMPF/IIaL
Itg8hU2nsfudd76qtkxVrmqdHA2IXcoVuDQEP6KoDOe7Nyid6m8eDJzgx8PPiMwf
DFgHnM6WVp9DW08+3Xejf4Ao5T5C11sdSeDQr8Ee/0dnM/h6voQjhu9gxA5YvPiD
+jAaTDOJZ9cjGALlw1Gdc8gEZgZQapXZH9Z3aSfHwiXVimmCo2xG7Ijj8U6F6Nas
fyp8uVKlp0Vf+79+swrI4Eozz12jxSAqQuMC2aFX8n1feZczR301mLF09byAgzFB
y0NH2u1lawKQdC8cxCUz1RSWbnm7EaoD35WGI14H/NwiCPvVqzMljsqMtX9pkp2+
N/bguR5043kxxfZzFllkLyqfa5qrh7TFUDkZivohsywbZjZvOcYwTN0CiRUAiWDq
zjyu0Fi3AQgpWWdbcbhrBiPjji50yA1lWLS8tHhFepgD4j0FZds0CnqKSt7cz6yo
GVT3Yo+/jb4KPUchA/dUPK8c+If9cpd+4FW0CZBEYfoIEWOlXn4n91GH+BkRKLTu
Iolc/keemRbTRv9MaxvSBYKN4gxdHSrL6UDO0pfggwF6/BhtYI+WOiDWqX51sOCR
Nqx5UYi+JYxMcOUTR+n43xk/1JTFPyV26IuoZQEBzLE+AFsxN3jOsSDatuAkLBRr
3T0T8Ju2UIOGu49JoMphWABw0Wbt+suP8hUdSVmymW6y07zo6tIgp8oFSLvb8arU
qp2/3rWLuW0cfwgkZc3f6VvuMMNSYW2UolPm/BC/9MCtLtjAFqt+A2aH5Bj2q/ZT
Pbt/UIxdDrbGBf5LKfDNIkD2CrOzv4AXRahRDgcEUrTMIY35Zy3dmiMQuTM0Ejl3
EAs2bTkxCL02dYa6gosXb+JjJVTi5E0LXfVyNaPRt5EdPSDjT8xFWIZm0HnObyJs
W4mTRdoyO11h231CMyY3pzcJubehFm9mWgo4uhVAibTxRbLL2UtJ2PqQpe1LXLID
x/SVR6IDhzRG0lYRupqxmzI3Z8pPLizeo2qQ3kmvtjgpCC4pY7YpHDEa0JElNw7g
zuvuOWDgfFIbQsv4WwEpPirtpSTJ4Eq/wmRQOrnPa/7GtZ46A+DxYFJ9Zn2Dm5L1
9jrf6LJSNTYI5d/IQmCvYfxH9x+a0WPuXiOxgrlt08hCidZC/F4+gDWnM14LjBQ0
LK4tZwcwdYWciewfXKWuM+rkZXgOyPKPzKdCMZf6IQVMHKk+zKhzOcJXJR3KRkPT
Rk+dSSOrzFdONO7+dgFsVWlohnaab/5NzGL+2oBlS7nzqICcEHWj4dq0nT2h058q
uUqvLjxliX2ThGbC2U39zW31GdHTRQvdHyGIyQnD/AtpxmuFWbxQ/TOX7nHcNXpG
rVB3yeb/2hWvJSjYJ9V1pT9n3vesLBaNBxnYUXwGuT0gKZpu9YN5i89wDqQFFIDB
UTqhLi9skW8KGUkE8za/xOtQW5U65d1RDVbrKXmWAujfMcW+u4lPhRHBNzTw0MYb
zOJMp3+uOrARVA4b9Y1ELglWSWesZ9X5+TQYcbGYFPWFema2J++cLHvwGpbHQg01
U3Y2bN+c2qSy5MmKa3Oihjy6gM8vZIjxOBAqBctcUSzphwTLtotskBH0WLFADJQp
ym/DT+Qui1SOBO+9a6e81Syc4oDSzZTOLQ1QtYvYJ2cuEELw+cAvI3uUNE+2LNVm
Et9dVlJkYOUPqGgIo2M4+rx49yo1yYybE0rr3aOsqA8cKy0MiDYBz89Wo0bBQuu7
qiXrPZNm+Ldo0m1cSM6XVRPX/2Vx2zVqhKt33B90n2W0iiJtRxPmV8yx8Duw/XbB
noz89z238C5cf46rUQFheLAEe1WkIfGhvM9TiRN/KEvQFGk3Wy8GYL96NWEunvOX
RW8nVDXL2BOl+E2S3JNgkpDFWH9zgQXp+0K4YwsUdIYixP6o1Vk8+xqL+2wH+hTI
GMi38ZFqgeQsM6oluduCoGKKnNdU0WlhxrFbFEPuqryp1rOStPI8sD1Pl1fGaqUs
Ac/WNAj2aT7AEDIqxA6oZXMvktxza5kzpH+gFGqjkAlah+24fW27KCW4Y0G05dsl
9Cdgo9OZ/Qo/MVUIhToTsrikkojC1dr70D81kZWlYJEGZiHHbxuUeOOqzNTlTJro
ZhA4iw6SKxBiz5sGPe65b0CH50V8EAn1RH9yuH/GIUufzbY/UgJjGi3jmljgqjLJ
KJxl5upghyStXKSlWycYEoM9o1rcWzaSrzN3ZcCm0TiQYWIuOpa+/368C/BX1bfY
5C0xVV/MiUwL6uiZ51PkFgXGG6xI5ngD4/GYAmxc+14bKBZDQuuw1MNcOCqUCcic
Ea+noax6gVXZ7dyFze1SQ8cu9HpWpQR6eQh+Vq1mAttz1W45SbMFJY9SlCfKYmXK
2kC/AiH1Eg5wVhUqbLXYppzAR8WeIuXDfB3mHROzoZ1i/0iVL+NUbFxjTNUG/s00
ofrW7vPJtdU9H8P9Pa6SlQhuCXEArqVKdLZ8xi/9MNz44qW6OsizC65hvwnFPLkC
QCti5wuTpC7ouzz7WnWCSS7IBmAmGvzYUQHleo/2U1LiYmCvAw+/0lCcXSxptFah
THh1Bgnj7+hCJXaq7vmjx8Adtk7ly7OKBldlTuQIxQiKBLzldqIt5WsSOs9MwJsm
wY4vVFmmUcDlawX9jYrEtgxFKcVj+jTxWIu1Mpfkm/RZTp/N2nT8EJS7k5c4Jg4+
tYwakssdwfoX1pVYeIHbX4A9SMHSnbsPMu9x2krOLd6+5ga4TcAUrtyL9RnNoQTu
0/6GilLZ0crFk4174VHip/njpp2N6LNW2mc7vDBMuq5pIOSKO7F+NbJOGTlwjvdF
aC+Xt1XiR45Y9oChAUI5uaxH9Wx0diAarL0tfNr1kgZ0Y2gxkT5Lwu6ZAUj5LqvP
UctZD5eA47asSpF7xOxwvuobX//168n2SK7LsgM/VWr77LpW+JtnLpIS4XH6z5d3
MQZeu36J5X1NSc3c8Cghsq6qu5ceczTqQejjyypcV1pSHVevW7loVT1VW8HgHS+V
0B5IVSLmY7kmdeenzNTotjqrEQ6lA1xhVAKCZGZpB5+mEQkKBMBzvW0pl1dfRznV
bGVxoVU0h6AOP7XiGLBUnN8zEgDfHZFc3//+vnOXrpbLdGdeUZg+Rivjo61/wIVX
0fqr8EGSi2RDySHbhRrsNf0Ag64RuHzsz7Km0oRKG2bSzpE0YTYsFffgfodmqSN8
6wBhwcPm+6cF/zEfs5HzY2FDWtgmxoZ3BjllV9YCPEzyjTcfFtqm0uk37oVyNdNZ
BG/oJjSHOy7a4HaesfPkIJFf1mAsXOz9C+0Q3RN8LwQ+xBgv8mjbqQYi3BXvv/tS
3lmaz1rign58l49ta9wsWFz6KMlN/XCKe4CTW2m/1BKsKbQuzGHSvCsDQR6vuUAB
61PuvpxvJWUwyYiuy1rnbdOQnpWmsyp57xv9xfkBjuJ6IivCrDukgHhBcqln8Frk
X1Tv3hJIUAUUp7p88A5sgFDEd+QR2GUX21OjrQVHaVQovwm2hE5fBc7cEq3mg9E9
3Hd1mleX9BwdCI71omw1YJIg3Y1cJ5xGwXscuexHYP84c0C+VQvlJko8z6/rIymA
zB1Zh8pKnNVM4M8XsSBpiM0KuUiPmxk3hYAh9s0+bweQggIvgxEBBb8c4P8A/l60
WWUZphrYJvu89STATLGOeSw52PayA/rIbBAdhaEx/1uG+JHqkF64OAOrPP5Jw9pD
OapdQg3WFuUvlPaTpxLFMd92zGbuc4kbltammIOAb3zUXQk9NC4VNs5fDIW2Mrue
Qak4HYBsfHkZxSU9eZ5Z/Qw5sm+Ucujv7qJxK37efFgFt+UpMAvaL+iWweKhhDlN
g596qd7sKZnpFAD2XtCRs/sMlX3x63j/3B3Clu/X1umkCjSksCFR9mtgapm5FPDB
s9A+vobMsKalwhCG5mfRZ0jFPd/6CMiAvjI64q4Jw3djRRVA3NiE8DriTYsXGhOS
0rAnSEL0uf5I/H7JNqVUokoQ4Qpy/1tf058+jQ/0h8zgZvgWSe9r12Nauee0vxPW
00/nO1Xzv/aR402o9ZtD3BFktJJGqSsMetXV0FJwDTqy9NiXPp+sUfpIQdgTA1YP
cXtVRPzmiLfsK6sdSC7YNnUIUSBBqMty7SjeaLVGW6iDRcLwuXtOWb1wW7/chDha
nuycxDgfgkPqJA1HouUujfHeESdgSvo08ELvny/qrBQ0+MCOP9pjuefM67iKD5xY
8AhRlLbOHcMP0s3KbbRKmLhTdwN/7pWKW8mivjNmqQrIMoilYzs4JZxrNBrZLtUL
NdOhyeYB/3Hp60+5KyvSVzkBPWDecRRV1rmcqxwtoZe09e34vw7n/lRM96urc2Z2
nxkVHk/946Kv+vFffOB6ftmqv6nIP8ZpQqYHg9Zx4Mql4AuBeAagTxkqk1SUbXir
cOXEuHX35vOTXeL2EIdfUOEmP2B/7h0zUtVT2dsIG+Xx52uJvnTBn5EJizdc1/yz
3XbZeb0b8DVIQd9dZuecKifmp/KF0azg5CQXL+7Axw1/ZYC5ABHUT7uLfsJQN7mW
a+LFbIVvTAqpBiXMU7Y8yOFqg2v+co3ROZDY9mcoWkSvwc7KT2mXPCp2s7DD06Td
hUmB46SrUjOwOQEOGUT1UMYz92TzYzKvlH2+qzS1lT7XKK3Ljcy+tQiFq7hlm/sB
zDwj+C/HzkGiedemCbM+me7RNSrbjUGSrRP4sWG9D3HTh+2THNPvtkA537gty1Bb
OyGKX/MJ47ELjY22NlOBUKmO3qd3UOmTTwFRqLoK5yfnlyhnHMUzHlZzRbu2Xb0r
1dTKBVDqaheBp7F34AaY/2gStrX4c4PNrffjXFFo/Ag56EKdeanQ9KsaPiL5jnpi
BAN3+I9fp1P3PbE2dspQxT7f1SN1DTyXrKp/xN8mwYM7l46QQJR5f0AAwWWNiUQW
sG+I3/RNywk7eP8XLVss7RbCsp5DygA8FXGF0Nt8PzrLJpFxz9fEGgcZ3+VGpT+1
T7GrViUzMWpJzU6+bMLXtCGYiYbt2YZNRkOhUswsennRGOODKgCKSs9nNp+hNiT4
J4R+U2tKz/YHorLkZLlLUm3G+b2uLaW/jxnTY4B/n8PUuEFNiy/AmvIpTfvUEbWD
eigXyzbKLWSmkYrx7YT4HkszZpy0KMljbIwRGRl3JgcwgG37PIkoyEtLTLZFIvec
0iMcGLeLoDFlEigT0Sc+qfvmjLyCZd/LyCvioz0W1wRYw7HI+llkhLrsVo+VGU1+
Vun36vn4d1tMAlNxYYLXWPxosX9R9ZpSJis0hBCNCUnuoQNQDSlfPhtSx3ZTHJRh
M/n4/f9lT/tnwwLNUx4fsIs4d/XUTqZ2pbHyVP9XqcOdxUV/219kkE2+MGKM7L/Y
hGv0AquwmzwPk6hCjCc17ISBnXcDfAzxitUlOQpzO/uMcae5HjzPuz3o29gtLPWK
irjb/IrKiKGZ37h4Vmkdfsbmqh2zdSRbaxs9tzXuseLG5p0ZAzAqh4xsz4FwQx4B
WWpSPrGSzAg/S7983ssso+HNcJEEqi+i9tvK6mx4mIjV5tyGcuHyHB2ure1j80m0
s39qBig8pzb8tfyldfNaAAnLmcUq52SSSQyioH+yX3lXTitwH0fNhf8eFHLu9fyl
rrISgxewMbqFLsNj6Rf6EtASvUk0oP+5N4gLLkHra2C8AlSkjezknVG3Y1tnhDK3
RhkGZyiZ9v5rkQZ35+ivlZcAF9ijdPssMUY26Z+VYuWUooBMxBg66a6WvK65G6AA
9qCT7jVIcrniKjxKuBG0RgbOx756EQo6IriXkf7KT+rFQ+PQVuy97ulpv8Fdwzo5
rHNao43kqlLdoSZCNqgz7/ZTux4I+YWkU1JBVxoOi/Qffu5Z05l0dgq1gcyNvZkh
4GtPzLIIouxxfbJBEWuE6z+ZJrTcPGJ7XL97kDhD824dAdhaNkY5M1TD1WW69f9P
RPLAxUgzIeIUkxQNFWQDu5Nr0xPeBJfFF1Bc8Pw+Sc/JF2l2yAIOlJ/XMPiH/DL7
H9ATVEq4j4QZD3avPkl7sDxHHootw/dNu4M7rN4j1rO3Ms4SuyWfl50Zg4YPdSc8
7peD++vg0N5l4UkmEJh83FlIL5AT6xiIkRiEiyTTodoEPdMSHnKHudVU9G0s6lRL
+Nn/OoveqedWh28nsuXPQgL8sHnIogeARYIaBFeLtGTpO59ujMJnIyG6L88EpC/7
dGiq30/hrb2gfi6clhS9IxnTvkU/xE5wP1IZ6ixb1GmXox1lRPcwv4xV3S8tbtw6
jK8LwOi2Ub/8CApTWcbMypd0JS6uXF7oCZRa2B//F+1d1Xx5gGSe6E8gthGk2pPh
ZYpmfsqye3J8EWXs+vYB7P+ecBpyOJXDoRkEqTl3K8mVT//ORAKUmt7Fks8Yz7Hn
2DWOV/NTNclyssh3txc8sC04i0hVPFxAAaghPYnCuMPND4Ys/uc33+Or8yoRxU8x
wFRQxz9edePikWW57dbxV25s5wuvxPapXV1q80qSIBmqlo92cNPKEhOvTOxm8KSg
HRZ/gYu26V7XKeAGvv8e6crYzOYiixkTvS5pgwTO4wnQ11j8AGYgZWY/qWIiWcAf
1OqtILd9/t8aksRCMhdBmfiiuxR9bD1BZo4iPg90XHwBbW1tLg0rZjeRKF++AiXn
1JiGbL19Vy5W93/YRzGEqFVC0fIKwiW3fgmN+rj2rlYq/Qe2zTvZ7aDuAJSLVBf7
l6HbGtaQdn+m3zd+X6cgwToXoWIUC6lIoS++3Nr0bLL23b63yQCoorg1oQ/kYTEW
U8kuvXvksM7q6je+GMtDmZegZ2c1i9NJ3w/ZwHrbyYiaUt8GdFLN2X0Bvy3RWJMp
DjMIrJL+CvPyv2m30LHVhPKOgNx0F900YtOnh/7aRTQhIMMjodWqFgJv3UnrM8Ki
CXD5ZyC0owVDaf5UU8loZgw1YvfBas9BDW6ZJIs8v73f/7dm+FGTVjDjcMr3qge0
iYq1ZvaZbWHz7gCpKem4dOUm1HrfgdOeZ05AUSsBkU0QOoIcS+qWsU9NjENrnfHu
y3Lt1GVabRLlVk4CEoZA2K776KMgtfHdmsFESwK570wrxC8stLWixE+q9dnJOvtL
vBCCWvw4cv/HUlpdPTIfi4zHnoA0+d3x3GmIz+JHYSRhBdXGTqn2NE/l4s7Ez7Jk
fIPGzkR3y1ndup5ZPsKYPoHAW9EGyOmiiqLa/bAvy7A6e2z7Tg7MYVCXIwMmH+AC
MEgQiqnrxcN3V5xyXlx8+oG/81gKVK8E6WDjSW3cUbYp0hSZSpc0umdBqn24+XMa
bgLV0v57CJhGFCiuajS8kvU/36YqW9oPpbEQtI7yIU++kmtOzlNSavkFFGXsQWdG
9cxmwyITUeNDAtG7mfeNzTKKtgumJ1p8zqGjLnxQ4uGMfBXi5I2ohtF4eNrN6YYq
aigAtV7RNTx4Hi0enGBn1hlAQz7+Dm5SNsChw3gZAyE3yiaRZMy5qU3IfOreuj6Q
6NqE1msWZgOqqYTGBVg1yyI4h2e5vZmIbXMc5SGEtifhmwXuL3Gu04CnKrdjRw5S
5vRT2fNpCdoUvnUeN+PZEs/jbr1rdYvRTps4sUNWqqsWSmDn9/LL8pKExO907rVd
lChZF5RH6LfaLjeaW0CjkMevDvdiauomJNKPHkEZud7mS6lfqzKkiV4EHK5kuuZL
sWH8Kd274vOs1jFiFMY9xwwGyf+sQyOXcvaTojNb4EdcTYjm/7AR2GlY9QbOWfFR
esAHoIc3HcVKiqa/bTJNtyApGIMLzqlZCP+pMcZa0e0N9mc+Y5UJ6XsVoM+A7/j0
rpyRBgmFI6ioPuxiyrVO7tJmjtLWTT2M8eLsUTw/TfkdS9RVVx9GeOaEpP7qn12v
oQwKNLexCUEW/zzsnZxip/K2/pO/xOW/Px9drObUXFXq8MH3WIaDXZyRQOa7y0rG
L8kNHiPsZ5I188c3anYQ7YN8zz2/E97vTNR5+2mC/13JnvVoNtkbXzXYdYl/iAdT
AJySZngDVTxp03Wp2ncHvbQ3msyYSO00ftrtdTOpzyyicVPkayu0xEdgONZpExwT
7KLruJejpgq0L6yRO/HkWs+AKgZoUj4vJddBHH0IaCAAgJ+LGIwn+EWiWuR50/z6
pZbqmDsDNuPdy/zUpVlixCzU6xtl8Vch19kK7RZ7VtkAWgsq4qkUcvuK6w3fEm/k
4iZtiVAT3BqXniMkE2QLAYc0DKJ5s0hQgCJ4GMYHZyoJSAeVq+BhnIIK+HngXhNM
g6FWGXCCpYab7fPEaF0vPNUIMNFf3LGtLlAv2VFmbIylk9RoGZMlpg0DRbSzatZz
YFdu5dF7bgr/KmbEczEtwuim83BrTjgGODF6MAUAtjuMFZpCTsvs44Se4kZzaxKq
nDbjvlpcJC6MHEMOEQUEUyK+nng5Ltz1yLxMpxDHZ3YAbmjSXvBknnMQzrr1RmzK
qwnRchwMLCpz4R7nNSz8raT9inS+9QX0rbDI91bpyr+UPvr4gqmU7yh9lASK8P4l
SE0uwjdedZS3zXa2Tv4PKTPLaYL+5vaN/VKf6qLJQ8bJxziFnMSlBBVZklzmsVOs
HvoqOGapVn5DyLhBpK0maIdO/OOKtTTt1Bx6vQOfNtuXsm5kHfDs+eR65jGk3u/f
RLb0uhreVbTg37NYI8qjc+YoSFve1iaq4SzyMxWK22Xuq8XBAkzi1GCkdkZGZyaM
EMfOXzErbRrQ+BAVjuh98gPXDSNWDXKhuUxfZxpHZsbBVPYf3kDrVE49GMtYYHm5
MSpPrV/URaX/K2FXjSKkLS7czY1hi8LrSRR/I69w5IIzoT6++f+00FedV7SExshe
bXnyn052sWeabwTzzdSVhQSP/5hNSDq63cGlVLF14wArCZPQd7JIqOcqF8zDX9+r
q+xNXYRMDtQUXV7O+cjSOKYfOkQpg9pEUPgv4OJA029HkG99UExAQE8yhfj4XGtb
K1ui1pkFDmTaXKV3uS6X2weNVnVSO73513CihM78yqMLl73rqOl8nUXIz7+GXw9S
YpANx3qa0iEf40Pf5gfgfMZOJajmJZ5SNuXFjej01y95qAjW4o5tw2XOi8Mk6h14
9XqyC6N+AneLNX7EGlRULDw9YBWvyP9tCreuowbc8oIW0P6fxZtZrCgGdxCWz9fL
56iBZvkRUQsl1DoOwpmV3/UCi03kIeD8U0D3Bcnb5Rc2X8bq2OHsnf2wCWbd57zX
a1YWwxyzSzARHO/T8QM/jdode4u7FLR1T4DCXLA49L7/7rYqHmY4gJqqu0sFgs9U
xbIdYh7YEuIl5VTaAGQ0q1Rv95dfuyN0YgSeEtDyXU+ytvq8LJ8z0k5skWSWZfI1
DXbn78lnJSP1zjq4GnojEYlycAOXdPie1cF28+SNW/7CCIVzixxhGjBGFxf3ULua
cFIxH202FH2Tb7kL7LngJeUe6iXVmz3js8/xQo0eKQvpo5Ko3tM9XKNKIVJXWow6
qJkkmL9fXQjsZGkcc4eSeeTTSaUc5C2yjDH35vWncCu1OjDe104FMDRbi/S1MDep
VfYAebIIz7FCOxd0Yv3dgF/QvdacwoNVgrj2l2k6Rhb77rg86sFr/tGU9CNIFMe4
zV71rE6o4OCKt1WmX6TrUsrI1tBPUE0ds3rtXxzOpw3XSwdY2F4vTisF4tJQrRsK
tsrPX/JJlPnoIgjc9Hx1eykIqVOuLOC90Px5eSROxOdPUgV7VbB1shiaDgcL+WVK
WkjyNUUCl/c8PN4mJM5v5sIEJ+0lzYqHH1dgarDuHAaUuPtZQ1kzct5cqKRdSURS
qwXDD3a0myxmA3WRb8rsx94C9GNqW6qZR3WlNvkdArCnIpCgxaDIEQQ954SzDzjr
pNbHo4Rw8rFS/G6VirCsW4SEZ1/o0qjYuf4J8GKA32XPqtCEviuKTgDHXSmzslxq
EpCOPMSrYk0ecaSmu12yfAuvl30o3cakBNIabwVpmZCdlibQR7g1OQMsjgQqmHGF
9kxB1Snjyu9U9gOTS76qLz4QYKYdFEU+oksGIYBWEY4H2WmNtBqCexJSEAMqzzCz
7t81dpmmfo9VF6sMvmJ8mKgvrMNI4gOEVtrFq5VoRGZOdGeq6S8a4Ntlq8eHtpcg
eujWX5yWaXKwOpFAJzkrkQpBTHa2la205IOnDDFPItjHNFdlTRqhFoOs5b2aik1C
+8yWsPXusCfV2vBcGapgFW+jT2wFm7ZRnQg+gtp/MEFfQynlh9bhm+TxSc5MuD9w
3NTkMwWQfmYpA2qtqXcwzWzZgSe8zug9bZzjpKjF1WNzgP48DCzMGCadhQRJkKFx
9rNnKI2vUCuR6NgL7dCfpFyC4ap4+19TCB4HH7eCPY4oSXSaTEL4gCzq2mXzrNpd
/z02dole7OWntjNib4J3sWhVqLylf6bLfjaLBnpXxdUSX9uCKWyxTuXjxnwE76j0
XWo0fug06ONY4fC0Zn+ntjrAjFPuX5m6/Np/iIxZSs5dfklNNUm5fTSYewUXDAE/
BvzcSThWN2evKZeMHTDpN7c8Pq+6zmsZ6qrEPZt56d4GzMFC+Ng2Peng1crv2+t0
2gmWRbbBqi4YmzHVhKlYPs7NtchTWwatzMuFY8LEKWHzL2kSdWWH7rhEsUXGVhiI
9aZ7MqUMjlnjPZPJ8WNfL0LVQ5WlS/ue4pgfUGUVUKUowYd5Zf9WaaKVxcel8mul
PMxd21tw8crjpsttZteCEHfu4Eu8EeF1stAhbueJtEB8enU1YwwVADjDehtp1kmD
cBcufRKw1zIlzXQfaHRH5f/qCcEpxsY5vMGTx8kSWnmWmko3lCqrIHRrXrHbmuA+
iSXj6/kb8+Mhtz3n9lVoiNVT5jQMv/Y7cxGbvj8w94l45zK6op9zekCDUHelPmVc
uZSGRNbgxl1kEI8VuL7TOqvGdELE9hF5Ufo8dYzYKdEErt1/+6c+Oq8MeKUVf7Ne
pToZtMqxqgtFnyA1YxBvWnXCh97myBM+Wf9yV8ud0tsv9h6vhtNFm4S6QvVtuuKI
Wp6T63/91Y1KOPqfnu2tl/K9eS2rMxtiNbouvaQa61mdYymnrkIqL5xcAEG3Kn1o
8W2Xj4o/Kz3HRD7RYtqFFKjKgTeyHSSkDW58O2xdEliSX1rXqbO9N0AjlDH85hKc
+DPAAvD8EWvru9GNfGHto9Zqt0gWdqE7QyTUmbXDrQjRf6PGaZznVWQTZ6CyeFH5
tjrsKHes6qw8p7CYFBM4brJ9eMQMjiov0Qnd9rpX4EpBv2ewiU2LgbchmNgSulK+
hjK3PE6G7mDSQgHoQMgjIlIPZCv3Yf9ijeguG2PezaFreGty+7N4APFDLFIaEJKZ
IyEF/GTsEVPqA65k/GZeHSPy31Mhl8g2Ogpso+n4JslEW4qXO8jYcQqYXZdl6a4l
CJ50I8DMPxefzCksljcJ+M2Xt45CXIkOSNUSSsJmM5udtYHtmOLK4QNhp28qVBpi
TXmd739cRL+freO+KOm1uXEJ5khhXDgr83R29lZ667d7tecUyvybe/9EXpL2wvqw
jRkYdFgWbdWR4xQE+MiTfBd7AL5Pb5735YrjdCtVHtsKfvnvXemjnm450PBGzolC
b0qVwYAR7I3j8yz2zMKgWQQmZb65cWnsjmt+RoZj/lyb2WqYjesz8Ei4hLlDZ3wE
TtJz6ESgSUVBOdCCEx39yolTDObCfzyOtdPmITL0SJQQoXikHZWwMz7ZEEY3SzpP
Ps0e3aE9X1O6I5SCMZAMUmPkJllEGnCeuxFbkza4qNC7rSAF+n4cxUx3V0Pel/jx
XvUw485u7ODxd7L9fsk1JOUbwpo0t7Yt6CCpK5eZsxyTe/PoPyabdANgO4frq/mN
yrfXEKc9GKbhxcRKo6osGoxnADBs9uIHKO4DNdzQ3PxnMGKzez3BgqKuXSfdzH1Q
QIiFrygAtiuTpyDg60k/rI9+18nuayFBBoHDWNvsIwNGGAbqYjMYeJYTESNzsBuo
ZZ7SbI0/dVqa5ut+IfR6lby/yOX9UlX8YMKmT4IYtqBm5i/dzWGab9CQ8PG5pnC3
ZCHROkAO9BPFMn5o4f7PqvsGObaiQAp9v4mcfNgyt7i6PVIbC57VHZl8Dkwk34K2
k4XlkBKpYVJMLdxGZ1sHxWyBDhIfwLvnd1NbTzS+W8k+zfq7F/ah7Ul6lflMJJ5R
6dWFJnC0JjLVb3owHmK4qaZYLzSAD5N4Jaf1mrRhSHrAQ523ZRA0N+KRCIseuK1R
L2evlVET/v322yCohbuxmGw/iLD+F79sBahAxU90VKH3XU/BeE4V+xQyIjKyOSYb
QTryojcN3AWim/g5Iz8l1wiuciFmGDfLAvouMNf7fbcPuRGP5J2wXoDLqDrO9YMQ
e2ShTjfmuZRGoha7sDPL6PjHcVwSiHa3QyK/1X2la+0DUuifIwmEfrrp0VNcYWLX
JORfjc+jLYy2Avah1h6kQZlaIyiOhQAGpWWhNe6vQMfP62zwiMN4rh1M8IOCYJWX
9AhKQaBa2QwvAJ7jfieTu5KUuazTRh7R7oUCUZkV7swukHfT1TGYPHsHNcfzNjMh
vjPi7s7oP7f65ezPVztjVzqjo5x4fPLPHsNE05q3TEfCVZAitpcS+gFJ6Aa76V0o
rrdeJZzbkXTd2W9uIJ4V8IJaTwlu/fzH83JTZaSILPDBlfcLDtktYfBCXYjfSg/H
bddDZHQ80Sw13+dcVerLAIsRTfTAN0Qw0U7ioxj2MMo/d1eujkpuWtta576aBLru
+w+HJHx1IXjLWKugprLZe3QinfD3t6PQBkNiYdKNAn5ugQxxJXm8ccRitxo3dHig
VOjZNgrClbF+0kwtFmE7nI8GfemF0l5uZoJcq7DSleYHsne24ajX7t+59EOPFHh/
yQufOC9QHhNWosUMK0LCrkt+ascE951hHcopYQuMHAzKxn18bt+WMand7iNOmwCK
d5+1LfNnWyHN+AZ5GUZ/NHJfxwEHh9g8ommH7gtPvAPC2afNSo9UJUZXJzg7AB2u
8mOMaVrsEuXjJ9tdZ2gsubcPX/x7wDgTxgVMWUFXLUDl7q+lMNxfKlXxX/dJHHUB
3yc0rStmE/RgTfSTN1c1d9QGaDBY2zjCpARTwT/l2J4XQ5sdyrDme6W1Em0sW0kb
dlj4zMRbRsDKPVXlfvmJtXOpDBHxRWUGJaAOSDbWiiM0MbN+8xzrFpZ0k+tymjPS
asSPMFbYL+g5JQ83rlYo2NTQFhO/o42vN2BXdl3Rv8PJotAWU+uBYEqWLp1tSkoc
WDlj53Y5LiIQNDfm9Qdhdchdd/TeQA3UDc5MGiCWdtZrK2+1AqhOqOdNufmu7mjA
Itp7UiVWzgSzV7r83hhkmtF868jUIM0pL1/pG3Vj/T+w1/93rOgXHxrfm1ELjdkG
ls34muQD2k+uRXfbl2vVLkcH4D4DjJ++2ep8t/7kgjC4+o6vL/AGej/oVjP9rL9Y
Q+xGn4UzabC6J6dBd7C3LPQesBDo/ZI/0d7IVLNP830w3niq/hDcHKBtKiPSAyQd
8GdUaVwe7C9YY6TRdQcJFaC3iO7mGniQmRcwGBdASSQXfZs2b73sDa6WFqaQB4cU
TN7gSRofCFGN6a6LjyMSG5ZS1yrqhZafPVed3AXsnAW+h+UB9ozQnoRbCGYDWfxM
L/yjAQuATwOpKJoum7xbJA5I8Mk7wT6o9tZuFC/+WFRZQi1x54raXPHAg62xwyGt
19xtZl2JOeZ9mak/bGQ1Qp59Ia1GqFsH6FvqaGzvWCOLzuzWZaxkKjGHmEsbf88y
vLYmVv15WjpepN8+1vtsqhzsl6JMa4c3EICNnR4sD/ge4/XNoAhzGWPaCmcvtwzW
SWK3D21URDGbfCify+zYsVW9ne+dzibDkvrNEcoEqscA9h3oFZyWyqhkYqRM5Uci
AeKiPZ6BljcOHjShNd2XqhQ9PyBbVF0MV+kaT8BmOfU8QX/ye+w78cKPvFXGIvcL
qV6Dn9fQjWmmc30lypaNaSwbA9FLaVED3Uzyr6t/WwP6duXbQsqc/FvBNgKxbnZO
jmrNskXNLsKzsIk4u9Qu6Zn+IzEwJwfQjpCJVqnxtu1TsA2mZmfWsjEYurAx8/jz
06BovNG9Ax39rA65YwZJJqaI4p9tj4oHeVAoXv7NTstKl5yenDfmJ1TlFSL3dSLv
CdgZcGrBgudB2aIjWoEHp5+qk8PNsx+9KMIwQklpuQxRB5YBUCAkiwUOejGZIX4G
qnPGM3FxakHQRwf+3ZUPW2di4kcoDF1iFPZ1I39I+/ahibr+abeGhV466cmnlSI1
+4DCgiVnFljaMbz9ZqqKks7XN3milCy+e85XJ0KkS2DNvK2nc6Gv26kO4kRstCaE
L/T85mevXI4MKwSnr+fj97Wpr9TONczbbjTI1gwj+YrgC0gSnaWl4hNYvb8l4xbh
EEE31cTVYrJkvCZlzYgjKbA51EqMRCoLAJyhuVUQuKyIhIljDFiz3wmfNHMhhMdB
xDIkSR4ZqgSGA+RpbRBYnMqfjEIMAKBQTe7kEizaW+ItYrGUx4GpJpQKHooE56WC
HvWctLIwzxaLiFb+QgJ9d5w3297ykKM3QUn+pvXU2lUBTbYGyWE4p6cBL9buRDCT
lPblsI/IPp5iRnCFWPJW8vdQV/41+4q3JWJhaLpw68n8A/FtlP2op1UZwXXDK6h5
o89MsFm28KZ+uIHyrimSllW6/HfSJDsN2ltZKChQwwRto2vjVyQul1mNnXST3nR8
bzj9FBFfMLOth+WkvKeRoLxfHmkKqhmf0xUVI+8eJ2ShOpDiX+N1ChwyXvr5CNhn
3VPSNwW4RpGLK8vN+qtfdChHeRlFJbTNtwrdax7rhaaa4wNFpRMir52X8wVSCGmg
ObI3B/T7AdoG7XsH2qy1QjPlZ6E0N+JtDtXp6CgUHg6Xu0bgrnjGwe78JS2DVMvr
jg8ZqU0McUqIk0GT6bdpnhllVG/kZivPIMXmMcADR4SZh2HMBVCLam6BAIicKsEM
1JjWpEhsokKwmp0ODAGYhuqBgAxvQDmNAHRsfn3cNeLSdRb+icKy2ws8+LTpLo+k
EI8nZN5ug25FRBxK72qXrJcmTMR93WQGdabxVqHEIEAjtsAmkYlAHuM4lNQVnVPE
FdJEdeCrga+9i+00xKRoVVJhLvr6mUNgtS5iUra2m2ifS1L6YmpovLPw+ku8sOG0
2QSFPn+BMDr//7jls2GT34OIg4lmDkEoWiL2roUP6Ee5OV8B9AIqJC2/sa6Hm9jt
oIwqTzcUTc2oRe5t+e65GZ+aN3URw9Z9qmrWUHh4PskkNKR3r+oK/vKptPUNH+9k
alXddYNLDav3w/ALcXiQ8YpWDBASUzgdLsivsqBCBpau7Cuef+qNBjrCzuOCjiWk
KQKm4ihhhNFRFPNXqqEaxGLV8uQ1obhB8L0WWnxje9xrZU9tBYeyj22p28rV/ft5
vCRx6p5InlUYJ4zfACQhzbNYgFgHQCu5SSRjkFwupk1Pq9//0fbFk4Oxkl6IYSfY
pseR94iIihsAg+bxgHOQLZpKwuOHPU9NXpM0eIWVN6FvcRrwC40e4lQGQAMPbNje
lK2uG7G1X3yTFeAkw9dEomcmlzPgG0UU56AOyEpL3Ly8LX+bmzSDK61XYr1qSdJb
hx0tfgtffjCTVB0iRmsvr+GC5vNwDP6gjsn1U5K9/PbknMsQPr/iW6/tkwVcYPlv
xvWQtwKvcRmmT1bAlLy7I8fOt2PJ602NFUuGVSfJc4xbmDscw5vJyqO/GZ6CWEBo
/y+L70lSlHoPked62kJO2b6k5AHItAGBWyXyi+55Q+OU8anXf2gqSrwFsdpxuFQK
6FJ3fWerZasFh4rYSHq/uXanFjNzM5Uz3KX1i4kgm2frUIrN9fySc0GSLKTcL9Bz
RRjkMvdDadP6JKjCVDdjXFmwU90ftK4ahHI2b8QDL6MlYKi9eMpWdEhUC0D8cguh
qIy3JDbXUd06R3Z9hhsqQhCBbE0LSM7IiTj/tkadSLU4ukOKDYGJJ1eqhMlYp+Am
0Cv64kS9fJXw2UTn/hxCRcXikGcXSfM9AReBg39qftHq+f2l2rVWWzNyoH6o4XMG
pFUHslTKvOoNyhn4anuqf3h8goSMO+teyY1FsYsHAImjgossaAbdC9LpzclKH1Zu
SusHJgDEwfKpWpM9/B/z8fTgAVoPkFl5gel8+31xvHY3kBcOz3K1syCCpLtx0SjH
XIHVvd2N9/spElYind+PLtBBruGcBFwjgxF5tPyorxyCEevP9+6GCjOuU3d7qJW7
T2vOLA0rEXTKla6EYR7Y/GZ7l2i3pk3ZwVGqPwccfUjGx+z/hZri5YvjLwAFvtyo
RTS2Qqyiu4T6ScTGp0bvwfjXMoD33NElEi6kG4PD83W1Zhm6IMX+D3IO7QOxDtA0
Naika5u04eUUOlU2Rf5A7UsW87ogcfX/WWEsYJ8RQJjoiFYLzy/JqzZZhl0GxqbW
Eyn/9IDe6Mmf9NFZuQH0w97Ceh8TgPmBWYDHufxV9b1Bb/7sulKeHaPH/jijFLTp
HKsSrNqFNRScHm5+ybNBTkEoA29HyaRLkfchoFd7IcM4B8Kf6qO8OrlKVQQhjQJd
cZgcwWy0LJyyHW6U//6M0NOkaA7iICraIGqAcpATv327is2AsTyFiCpyfO7AehLy
74C7EnoQqiu+bUcOLZLkiDe9jfvHhVdfk5JR2mXRPklz1BvCVPUmyIUlFROal1iH
E5Lyx9Kd6m4IbXOLJbEWgMJBL3imk/Ha3jFBKuJTULug1xcfYdiBoAX+Z3LH3SP8
Djcl9h0Lo38DkoStflYq/QFXp4ljf7jw9Q5PsojPUGReeXM20Ninj06TPcLxxEfJ
QMKxm0Ibwoc5DpRkGfV5pIu93glz7Y1tYySIwYyt1ucbsrw3iy5dMSng7fFBPixb
hKdr4xFZ7udbyXeH57NvirVdwxMbxZRPhcCSKVnKCpSD0cTUW9nj7KVVy2X3yorg
sG+C7MUjt3JLjk6WgU5o48AHotcy7u8zfW4NBfry8/mbUGJDecx3PZ4No8yWiQDP
x4iyDg5BrgNWoJmwZhPMN9erDJj0+0CcjcTckCm7HClB1ehix2LqCmeGQ/TaJ/CT
5InJWVAPhSrsDyHOZ/MQdnI6CO/sCtAqZPtPt/5ixSgYWLcYuovlMm2mkQxb21tj
I6aiuEkmAZFTuWCmF2y0NendNMed11mBnATFb39+iSZnY1/0/Nxm6mCZQCgXIojr
WsTxkjybA/a5Mb76x7YR71kAeSRwgfYNEnUAk/iAm5eo/2meSx8p7Az6wifA/1Se
06OgrFZoFOwrwNwsHhZEHrunoIU9QicK5AzHhpmlOyf+z7tLCmWFFETuVc1Fyh6b
YIK4XyN8z2DehKv5G0Pjyml21fGVbTkwoyh0Djg4akx5IAP+yQAk5NaLAMnWaLA8
f6ysm1TiS2PbxLoO17vmfRUY7OmBqFf5lkuPoVrnL/33seIpFTkGuG3kPUgjBiBt
mJmv/U7jyjkpT9AwaQelo2ghl5iOyDKG7kZVt9xcrDhOe8olA4kxjgVIs2w9ZcRo
/ObbqY0xoLgqkf6M/zNyR9lAlUjJMRl68DpA03eTt24MUaEtq/ulS/vebeajTGZE
ysx8Y4ytSIL98zLPECIgUCToBHyZjsSitLlklzSSQv+jrdrcwn/TZwWRLe/Cj3N1
6E36O3bsXTbx5zIjcNynVo4cLwz/X/qlVcqX0bOBzU1dnYhaid3rc1/G68YiQuHd
ZeNwV8Vu2RVQbNqnvhthDP9jqE5NQUBWh+FG4l07JkuWs56okijQhsnTATB0EOFB
g4MnVd4zaGUvOeu6eWn6/UJ0qcPS/kg+2V5PZJAkodsrFd7ScLE1BRW2ar/1rWDP
PdeSwCIStlNMCuFySkzz93bP21V4QvO39SMu7eGCRxRtaG12bXwRv38d3Xyeoa33
mFAzIfWE+/qISZjPZVxwJZlrEi12w4VSEkxbCNkqLVKqtJKivWY8mgJC4REwEmXK
H3hh46idac6MB57dejNNBnSJdzH2mgYfwEU9srCiRA0pYBKsdOXp/A2aJimyb6rs
eitOCnG67RZpR/k47WLJJnD3GwtbllzJglBsgETVJl6PYW0QpxsTZki7Qj9yUrXj
oUHb73z0Kyv2t7WNhvLADbXamUXaSt7nzmqsWCtDebCieJgbMxE+2usbUKTJFE4e
Guo2poqx850nir03SHJGEfwNJhXLHOW/UEsOkbr0tNXEsGh2GbcQpHW6YdREJDce
vaB+MKOAvNJFC2atccv1/vrmaIlhrtfP6P2tcUvTwnKKrzf/K07i7Mpu+ANffAtf
k4HBuF3eT9NXLfqfp+EBGjkG34ig41pVqO6sBbwUzKzqzh2Cy47pHJJdGRC3OC9g
asEcSa4BqZYHH1bKfLiFpo15htCVGuhLUXSvj531Ij7yCk+18nOZTjslNFs25o1D
k4SygPE2PC/JBBc8lhBPf/AmfCNHlmyx5HXo0typ7c//RCf1fmK172fJqcaU7Qbp
70DLs47Jka9P+jlHYU0SKLdiEziiWLiD44Q238piSAkRNG49d39CNgHrgF+QtYLi
hHLwmzOsVp7MqEHkYJzpTaQzYsI2ztkLlCkbva6KqTx1hKkKPHgfn/P0xx7rXBci
+B571s9u3MscbLlJdi/qH4FfV2/Jjt2W/65TfMNf4MBC2qdSWMdv1jNJwDIVb+K5
8bhkjZWRSz1AVvRsR1SCxadfTiT+bgfFmwYi7h/4IxWQZwNYb5wdgFQVlhhfjmh+
/w+O4XGgrIfFtgU5le5h1Nnc2sO3Uk2UsvAvfySXh/liKOSw9eCZpvU6v/srWcwg
0PkPBUyEmYROZagUKmOmuPRXbGAFeaoS2Cyvy/NBMjyfhuPL64pRpfqHeKZG8s5J
t4P5r77ZKQ4byJpX1b2snwt5vTaATQKjUWYXBblWP/XIRZFkZUDfwpCPs2PMFj1m
ZfZofE5anYguuDobL8KmwnpyTHkEzxDeTKIW7X8i0pjOTEAIk3oz/JrZYIzf7hUa
xWuiTgPVcyfDcHPnjhMj3tYJQdsAfhkoue6xB+jbVBef4O/8jpsVzFaIcfsM9M/z
8MJ01gXdI9n45AdI4HsJ3T2WI61xHQFlsVykhoTTi/+8X28tcpnP3aXNXx+SJeE4
yneaVD8p3YeCFU0TAym0WnsHHlNH0prKfOJji5gXAxqZBxcvz6t06I1ykmXfEq7p
+SbVsnKMAfL2wRwNQ7PG/bFv7sO49KZN67auzsHIq0Bi5l7U929w5VPJD767kZzY
INBChEulkCNydtc+ZUKxqqiYV2gbwhJYUNBhWW9hFMRrND2HooSMc2iQsl1nWZ4C
vY/je+74fZFWagWQkcxhMQqQIZh15gMv+3rixpwWQhy9LVd0qhsYtne2YhbtG3cl
oGoMtU3kt5qb8/BmvmrHqH4k/SMhY0DSvifORPjveTosqP7IcCcIgPqMA4llKLOK
vdkb1BkXcntJetwkPeGrIbzySoGyleXIXpHbMHxR75xii6ehhUbyrH+87iKuCUgW
WOcJhq4z1fg5bQnQE/9SJTAAkZoR8ax9lVdNIy1TXrdUD1Zvo7kjfKLCNLrXBiy1
FbTnhIUP+IDGtGFUZFjXdZowOynUNsL/iT6W7GCOuFTeTxGrGygaWo44otsJaIwK
fCsKP0A2GfnODqQ0U2HvqRYlCuHWXR/CB5bbAVqJON67ICIOsUeBBniFUZED3Bhe
Dhq9mSHgWxm3B/mrkMwsYcLOPAFzU2vAeulKOH1mu480kyQClAkP+JOnoeVlm+mL
pj5yAAP1n8TkSTaHVFK9+1GrxouhgEl7G6eyJ/sFJ2+U0K/DLRx5/2W43zNwfVfe
/R0DUoNybxSoW733ifS5HvYkpXTPEekVSktP0OC+qQRjTuLRGfMr4JbaS2tkSOFF
77Jd/hXl13q8mVowW/+rBxtwSEkBngyQhvXOsyT79WmiuB2GK7lxET9OG3D61bqU
cgQ52NZldLm1dgHIzwExgRjWmABGJCNhPA6vb1q/ETeUrUjFwU0IYWg85IufEq7q
UOlu89idsiO9WTLxb79dbnatWB/PZoJDJiT1YkLgRkw07OKhnxoiYdLn8Y0SM5E5
ZKuVXZAF5aRGTtTrrZ6fV7umab6mrzWKI6u73sGX7bOnTwGIKR4htYqd/RbzysjG
Ea2I7wP4WPNOCMAGbW/WPPWlEcqmb5w7Fp+SP6VfPJ/xo4Rn5S4xIU65/nknHQc0
MOLoDrRjPZ16hQJNtaMAiI/zZJsr6cUzKRBeMiYQxbKypoJlVP7uAPdG7qV1pmJS
KmsRrhJFR3C99xykTih9gufbkxhY9gpqKGrhoqt0+VU9urovRMUQ3RRyyEAtABte
JTRsk21tjyNBW/wTEG7ak9QM2rBra6oXkFJcORLOgnwYb4lO8T/1fch8olHZ+9fz
g5lOFwOXyWcNzrrMJ3GkCgo9cc4vgV+UPDukMjc/Vis7U1XJNj02wNtncxTJlQH3
E/uG0GCnSF6hRphge3+7tN5dpO1bEildoc5KFG5k/Gp9lcEouUubFHz+o1Xb5ign
Al8T5wzXCxWvIsJoTS1dkOHppJ/Uz2FHNbQmoxx+wS0lQsxjo80U30pj6A7hVfyj
WoV2jp+02nJn6Us48Gfe5/DdxzbtrElmfEYUXfTJFiCfjTxvbhbF05QDQ7v1M7iY
7j7bGUpemqLarOAwEm6Gm3vkc9JNeAbSuXVsqMrwFfbyC6Ezt/2xShy/mzwhMrGO
p3WA6r+m6MB4Z52vf/+i4Chq2DByxuAq6non8pfFBBuzUoK5TvGUwEkvZ7irSW0o
2AkHo0AwNL5RQWUil1s8pqckalUfOBKFe6TnENfqal7M6v01EghDfcvaLn2HvahX
Oft4hqSf56NI/e+4wfczQLC69xHYciuCffMIvA10Qmuj94skB4P5PmFOpF55+MrE
jgM0Oz7BZi0Q1AofSQmIU5AdgdAWG9XEF0wpTr9KJ6sEx7hC742UBKEjc/6VWemK
M+BKPiau/SBUQNvDfweb50s1MsIjtVv33kRl4+zxgzQQSjghdUIwut8GdKkJ547e
15scOJ/Fsy/reTz9mx0XlsDJT/qd6Ic+qQfLeHhuyb+lEMZs+AqfXcTvJR2npR+E
Gyee2FKUZ1/WfYb6DpXQnxWfsdJgYj9/6FFNLjnw1qqGB/rGBaYnBLhPvU1NBh1M
f+wrceCRbRGcd/sinAsf4zFf1U1otRaqna1X9nsHQiLymL8mU2DkK+jkB8zpNXv8
BTwcVgOpYf2gnCP//60wpzjI72adPoCRZ47dZvVHjAxXEQJLNDv9caiw75DFJPjq
Zy6aElndVkKEj0CrLXjUUIWE9R6GzzrC1WUEjJiLsIY/TMLDPLmcjNDb8LTPTyxL
6w46nqGuAicw1CS8akLqQku8zEBQ95YZeC2AWLJppG8+YQxYOkqaReewgX1EWbdh
9Ufs8b7WT8SJKavQk6XeF1xVSW9re3rjf449lllT2++dyukLjTtiXSpCub1n4He5
jlOGoGRk8yfDdfy2qBDt0D+Ak98syMmVxR5KGFXKU+ufEx6qzeBD9vXnnRwiIYtk
aB3o4ywOQyu0AKlzHLITDlegCbmZvMEV8fvpSpcJ3R3nR6lOoh2XACQrSD8TCoDR
8x7dsTx1gq8vEfIpG0dKSTSUMnyNb1Tb4XlDnJYKb/p3QlF5iqyd0VERDAhHL10W
+4ACpAUm8iXcrytpJ/5DwLwAlp01PtChEKqj5/A9XAueiKf9n9AXcur6P/1ooeaG
MdrupzKboRiNjMrleNyFa8IbQXo9TUxhjSXl6zUW1kR/aorLEMw09xMsJVsKjiiU
fb7TRmw4e49UUjksnYzwEFwBE7fSTLM04sveDSHz8LQGhdOsorJt13GZewKki9ql
bb3aI9DPGUqWCzTUCgBjLUQkStvJuJfXAvpzrz4KCLyaKRDkt0moAOjJh2N6k5ae
xLlthC8bJhzhZNU6H6Nt0+RYfLSpqwVuSIr8upU6H50IJyUjEa4r2tpnOp0+YEPC
9kRTTkgrhHlY+IqZfD5TPYsdAduutW5LMswYPE/vfcklmj8lnDpIMR0F6M9nI1NS
EJOiwu6EOJ2dtR8Mn2Fb2jMxihYqLl1mp+ilG1P/YCnWeSUpTPC5O/Vv1s8DCWc4
ndrojRln6lHx96crbYFovvEHXUQxZcxXLCva4orjJV/72xNAtZKsG1s0TrNsf9iE
7w5gY0Mj1/zTkON+dD818wayUTO9JKmf6sKhHJiK6SzgxDXxFuQDEV3fxYTd1jVv
kqkTzJsHORI0oHRzp+eeSLVg3DDxTWVJJbXxN6MBynKHO8ESRguaaroWTV4woq0O
Mour7BJGh4dgVXnzYb3Fc0X4aOVP15/1KbyPOdFfrJxLUMOJ/qo06jzhVnnB38pZ
4IglcMLWCI/uK0iU3WmzRwv9BL4wFp+0eeCFUiDBYHSzWWhvQ1gOWrTrfQowmUd/
SS1bgZhZ9ZYgNc697nNWdtWrLJ9TU2S9CjelgMm/aIQVWkiohYj7cMXkB5V55+fg
0TmNwBlEtwwx12+wUoYAX2wcqnO7sjKeDclI55Dx4xfHq8X0hCJ+jeY0o/myOgpG
kM9XljAYRVVZgaClwEoHDQM/cjNbQnk0IotAW8RHZX3zOh3O21NRzm7Hlg0vFxy0
6qpQDUTb3522hxoLTgTR2rpjTjTANDOzGwtz7WMc49S3L1zE9mDL77p46yxLM82p
s0W+xF0cPguR/ibnoXw9XOZrzrpcoHNn8dSGwQQuCg0rTfOYdShWr2KGk9AbIhPo
ehl7LpQQjYD0I19IYesfEZgn2j6MvGRCUKbC+lRJ/vD6wwQJQCMu2uHWxhqlGB93
juuvvdDEws5WOdo6+tlLpd15flsSm69oau+1IQI6wN97KykWGYoodMVYicQaGUKE
FTovn2evfyF93Q0aeAcveaE9aWOEtichuJbBh3o/pXjUAs2sPctezZZqjoNcMcyJ
x6tRqkD0JVKNq/DwvW97Xe5houdajmTzwCxXWwQl8D/itRVEIYF4fP0JF8ZMX1OD
riX6D66MFpCwtszspboH3n0hJkn1mbKUc6Q1trB43WKZ8XeIUf7jiCkbIuAj2mjb
FK59uahx7W9oNIvjYuRxsvA9SSXNI8SEfDVZDa9HHf6c7IiiziLX1jaKrQSAC/uT
Qui9Rthn6yVNmYW8t5en901MnVJH1227nnh6YBHmNZnp6xJl/E7mLSZjuBLu4QZj
BKm9ixkfmAleUDElaA2vVnwLoYfvo/+RMcMMyRM8Mvr/tS3wWAKboCzFBUHsY7XO
6mTVXV7jms+nnAGUXz/nktz+gTKoat6dCT6XGt1/kpniwHmdYELPVJCvZIxNIXK5
J4ppJZNt6ODIbSm1+4zdhE4RICOub6PNiwBfPRESUpLMP8BNfAh/Kg9qiYXNUw9w
TO4GrHV6I58mofeEaatqs3CPtJTLifpXiIhAGZIjTyeyWXPyd8pMytnbtD2RPC+p
bRCVqWjNW2zp/JfZ0ZwJCfaM4Y+GbcVrhy0Ch8kcv2hPJmDGaIP8htXy6gGGaiOe
yDnM7s5BLXS1P0kWE6Ak+iLvXLY0XQkHmi1Di440NztBVw0aDnucKSP6o1j+D9fr
xsHy3TfuPGu3EP5/vomggFcGC5SyZwNsoZihDxNx5IDVANo7AfYV3d5YqWQLRbea
Ss49uep5l4oL1FWAoKdwFH3me4pHCBC1ThqylY4jA9gNx8pR4mxIoOj6BlijMlC2
qEuMWA8T95GM7oWPdBb6TdIzZsNF1SbCYHrxWJ+8Vp5eOXPUJx5DYakWwPVIevOi
vRdmOjRwEuPHAN2qjQ02QxwuBTwTxo+MPf+t7JG4Y76Z4gJ0nrrcRJHDGprzn1+E
o1dcEeSuHahmeYEq+Wt2JKo2HCqyBILAZ4cb23yzAJ+gTUtWwMocZ9MWKxkcMJWp
HkG9FbSEfNbEdZzhPMQTbpmNt/e00iEVhdZIAUQhSXmYTAfFVX6jjMEvEx8vmjyp
QV7rDrOqK9sOOtRHbaiyD8T4GGfEYgUgTQqyHtPAGLcn9GI9l64aww5JLERXkQ4C
HjKZKD2GwhlD62UnPXquSBwIoe3HmKnpKMvUHg5m4seS5jDEmaz/LYaBsGnuINql
EpDAdEfy8JoFjZp/2aG2TW8xTHAOYsCg4Zzam0zh4YojPPMpCvydHfJuCgRJuAmx
Cws3Ep+RxvdkW8MLPh1Dpz5jjrQenyI3eBX+SXjT5A2r6olWc5c3c22UUfMibjvf
AjZR5esV8kgfo5lJsaLQH/nELT4VpxM8zaQzKTR2I0/CgD3Bjr1O/P8PySCbXrkz
80k9Jx9skQXft3hPFtz4qtetEDSMtZBKeSu3Jq2d6d2X2RkqfrOCfY9Pu6XZuiQn
b1KcEG5Pbm+jxkVCouEoN6lNQUuEgPyeg4vPTlk4hypt9TuQB5rSn/OQdzaKGvGS
9KzTwVv4rFYNFK/bVN10IRuqvYKJbagTEg4zxBbhnDwsa9yGjfcvs7+JProrjVbU
Oe1lO3LhFWB2T2GQG8FQ9INcBncZXFkNV2OT/OnOsjoZXGZ/T/4R9+teFLo2sN1X
7HUF2o05ojj1pyWb0v25r4c3X8+grpoGLKytShBExiYPKeFZATn5jrTbM2kNyGKk
MGoZxlet/HVHhlGPax4sxE61H6Uyfu63E9stP6n50wUdiiJSM99WAi6wSasPoFJ+
/MiDNuhcIkvgexPrmB1Tw8aIUoSqDseukKJsoj30GwYU+/XaNOEaTn0vI/qExp4e
1zt7uZZ/N/2rIAF4ZxDVxEt72PCd+AR6Jpof3gG8+ixBkbqtV8TMMkfAQ+D75/r6
jtgPYsLATVg0+btXHrQKOpa8+o1FmDR1JtVx+uL4zjCYTnfOsaLAS9pfG7P3dzUb
PMuCL0r7MMnCyKUZSoKbI6a/cQpPzsXFxVcSr0uTT8oqbMzD/y7hNqAiy+QrtHga
4roGxdh+8S/kYIJMTywO3IuI1k2VoIVzaQgyPbtomdZop/ptZLK3AjPMRaKFmK+m
HBGGEmGO7TdNIEhFlkCnYmG8Tho931wMGLh2BaOq0L2Iyl8nxmpoGqbu8KdGoyjW
oq7fY3ZoOTQvc8eMnaRN8WH5G3dAAjsVVrsMVwDm6M24IP6TB20v7Q7AI3044/JC
Q9+gYPvcdNGl2AxtSQL264pqd/+3i4RmCIkM9y9wUYcmWkTHwCFCvkP0aAZIflcr
60r3beOqqACtITaIIteeay4J+yXuGgMs/aOmihMayYbFobU+/yq5kBbo6VtPNjrs
gRWDnAgn21q2/gFQkGDMAP8VAN2+WkuSf4PvoyJZGNUhfuya5ZHoDUHwyfGQDj2J
2wEG2PN6qMGMwQ4VY6JsQPCF4e2DZvcF8BkJrJHwc7Ahd1iDGiNcwm5Wac4JDN4Q
hS+0VBCOvrqDbc7woNSYY5GVRnxROUcJWpXpuTBhxEk4qe8y4dlICy5GiU4UxBwL
T4vm9HGJVLmF90CMyDKWVytmxD0ORIwXhYj3xduJXSfNDKTAlyIjg5m0ffdcqtDr
K7yP9D8lgdW7DAfhOU3lbJQQCPKZtb+pa29VKQd1f/b5vCh8ANrKpKVyenBvcjcP
9grq7ccJeDF8FDxbsDJrTqvbPUpPLUquNo277utkbCy8wvJp/S++cLhGxu6QK4J6
AylNPCBoBxf4S1DLOyCpAoGdGGA7Q3bKCEc6gNLh9DA7IgQBGslvhifCRJKFOwrL
uaJuwSCyTL/+NRMehur9Vi2WdRsqHsp2kpKrKcq6Qe2/djVqqPpSQMy0BwjrnEYR
AjAihE0JVFRwqGEspBYBdIB2zwPnaHz6auUWA9A5QZSMLs68gEIvfjNA5oQShGiq
0o2YpVj+d7wPMJw4XTPVXZc5VgVLvbAkHpX1QhspbnbYDs1CH4QRLClAzO3dM10I
dCaIjyojXBIk0XXZUmENIe3/XqdQvZ87O0WXybvOiL/muuxwF+1eau3Kx2fPYbjW
5R8bn5cKEZ8qzVL7cPNT1JzUUQ9kjiBSPt/d9tpY1QSD/niJGhO/Hr+jXo3nw0lN
PclZBdMuI29Lh+AkDXQ6PlsbeAa6edqytSSF6auP5639ZTQfCE3g8V9uCAyyKkYG
FO3fS/4RyByVtDkZQ6hLr9QJkjkszlmb/MY2BK64NUJnnEFy4HkM+XqnzQUOyiWJ
G5KuVlHSymnMok3LGT1PzzCG3ry2OcDdnullMHaRgWqilclQB7ekY+4evRmf1u7h
iyy6ChPQ1zQiQHwXy4dQhCDZ+gndxuEyjsMxak0ZXUWWnbFwfxpiQIlZ0910SHHz
O1h09o/vRgcgawnbrTsmyTWMTs9RFuqlllBqzLGoEhVsx1Gvwb2sxNyvMS9y25Bn
lfaZhpkVlPZTcL3O3ndreAG8Em8FNEdAL5HXpgETYdqDACCRrcIkLGBdOnJrAwCu
uLTHAmOmIv3SvUpjXOYwsfyHb/eTLYkrzJyle3z9ZkS0D9mfGb1Bbr7xCwHKL68L
xvb+ZDmi/j2uoI0+ZCkxFyOeQowhwaFm9alFe+waPOrwUNNTm2pVGJi1Z6fHxalv
xzirVs7myykbJ2eScTyF/wJkB8DUXW85F6rKZSQzreIaW7Z78jCstTcS4ujbto5P
lt1LdTdto/rld9Bypt1ts/Baz88NipjD4poXnpetlhPMjr/zH9hOzVJsg9Nt12es
VEIVHVafcAPl/q/pyBieA07I/VVTpYhJ8oDByvldM2XDn2NRO7n6PtujeB5UfekR
wTn3TxYWmoHgeCzHhiXti7x6X8lbi4tZjLpnc8SZl7pMc7ZIkmp0oNoXTnV/FBgI
zq0FSGx/Tm1RfaEwyL184FnFXzrEpf1vp/r/8uP98lll4Kr0NdRgp91Ic7qpoBXM
kCq4cTUISWkONfHroqMIksW9tEGmbz0OOup0ZNQrbNPP2myY3VqIaoP1JM/rPZSg
i4f9YL05Pygfu/NRZ4w/OriZrGvgTH8mu7DG9ZczyUNa2t+RQnHZf6OyQ6Eyy4JD
qjaa1X72/GhKgqXT1t/lvICNDfagJVDs0dKASboQW9QP51bcWf4EgFARoiDx9QWa
da0tbxhwAVTO8FQrCJwlWF8UXqOgf4Uz1o5m8qRbbFLkA8sL8vg88Aa4ytgHhNdK
ouBbp5ChTYQ/Inj9I+2anxvRPKI8VaEg38zZJUM1pe2Z2DOgpX6EDghWtf4+PWVR
FFaYPhZDc0uoZduL7/w2PZTWyW29I03lKmCBi9uiQB0hJ1+eqTG534jSPmHjdTFx
DFJ073K1kyUjwdbWcxzkKl5tjY/GKQ/pVSBFSlR+Z8jvElkzPz/a8QvwHlvCFixp
gYzlu18XdU3OCK8L6SE3slc6haLwZHvTSWYi8pVV6UybAq0dH8KCDiwaHIlbMz+F
lPwZyIQNHxeRX1PY5UBNWHaZuzvHd3ZtsjcaDUh92y9bLpz618puXj8OH5h8OHSa
91WvmHFH+5EVmPRvOU5uug7wEYmS+Wy15h/ALWG31zHkDzyIDTHsCrogn6enaZQ+
JWsuW6rAYqg/9d+Ro6oigal5Ye5OkHsRC12wZ1c04ll8XIxjnq+CRKAUPj7a+exo
5d81A1/AcFslvjCyE8DiwDplrkb0+bPuaIVDfvi2GM3kenMyaMDQDKU/fTGrV/wy
5cEQU0M2JJf00Ieh41uSbACcnCjYfztIz8OpQZjS+rU5eFArvMjE0X0ADSce7Qjp
U/8j4WwgvEMT5tftkrBd5B4mxPmFq9ue2kIfzjP/wLpXD5il85we2c8tfQhopa3a
2tnpXCvi9NDBWyhTQzRWMvGCekvItoKLouo40zup2tAuVntmu1mklZnyW3DqLAKY
erh6rdkYso3+Re1lHmYQDWkQzyZYJ0Gn23P45zcBjNZj3ncppKafqpUvSNuHTM2n
LjkBJ8vxBSm2hey4ymzIaPEXRgRmQRvToi/PitSatVnikgZ59F6uantVFInLssRK
R6IQKeXXzJsYpFSNSUJ4pa89PTv9ahOqghyS9kj9CkHgmSvwL+IW5vdPRIe9IoQS
hrQ42Cg17T6TdqE8JPB0VBEJfKEz8XIFQBe15LPLEND/pBYCZRx8lUxaQ0tr9hkv
FxZmbLxNeVqsogLWgbEJfRZkW+lLiDx1fnN/YlwrxaVav5P+p2WLCMbRBUfZ5dXn
jXTbrsRE6UR5baV7BfSLfNLDRcd8jN6m1XkpbGdBXzg1ldNrmfAydwe2eF15lRpT
o2SBYEx9EiHy6S+zauReYStvFfFsSFSPWQYa33iV5bTkeGFFWQSutKw7o3zI5frX
Cv9lD8BhDtvPnRaJDO+d2IWuNh5ceHDHDu98oaAU7gZ4N/xMIzRtS0bMHz25phAS
4NaU1g1xjs0Yrf79h0ppiIUVT1atMttzoBvEVHTifMxLLabQ1QgAzzSTGaaFFd3W
tERf0uI2VxhQh4serlMqsd35v9JTDYYBn9paOWNObH27MyJyOA6+ZmxE7TbBFxR0
ICsmWapUDXoKkEakJdB0OyqW9Ac7rYnI5OX/yvLYMM7RAzjjoB0ESv2rGDlSDRhN
H7FGKcBI13TABGwlKZC2SU8YHhkJmuT6i7UeATLnBNfvjFsfkapOxuSh72FgNNMz
kyCMXSVmuJDeC4MUrzqcZZz6IyzS6MgBSgiPIQtUrcg/1wK2EsMIgDD8QEjoSbmW
IcoNGaHD0FQYRrQxb1u3Y0ZZjdKeI72wooWx/YMUPJyvmmiFWu6ytbSUaUKHg0+m
bNo0d085ATwhzgLqD0r9f8GmBszIAK873OzcSY1cnUurCd2y24cLRUyEDJCMhNmJ
6V3eEyUsQsOL3LP8+cbaPBaFkwKl0vHuCuFuBhRk3Pa595cn3RH6xohiQReE9u8v
xnryjPbhnDiM9BoW+xQeimQClIT0suinXhoq767AyuALiuD0fMlsiTl4u8u4R7z4
bxbsT9WUDxMZWWXHUQMcHmcIA9sKINy7tnZd/uWLaJGYz/UMv9y78OeeY9ewaXp4
vTUgKUVmiZ6y1GNbP778AvC+Noyz1mnAhG4VxdzEf1mqZ+NjmTvKC8RJOveTXAe+
BRtzo1UjLXChju+3STyF1L8+tUYLgH0nrxt627NATIWERVayUnv2KAS/HDDpFAJy
fZbZfc5b1fxgNzqOn7qWXJM7xjGam07+fbUSnsVkxrNTg0mSgWpLUDJgz3EFZRzK
oWU2IuNWOyU3VlY149mws+YpYoC7Z/jCCpPjwKvh6a9fqYcm4oHFPz1E0kTWGl/A
ooeZYVo9ZGysPi2aOZbqO8zGy7K/jGvRt/3lALwWu6nfnU9b97Ee/w6K8YdXoiSI
UdzYfES6ZhfuC2uIv4vl8Brj35T+7jbzpOOUm4aIBRzup3b2VBQyEkIpyC5zUXI1
CJwkd2EWJDo36PmlLPwXCo2tPrHF3BbHt/Wb28fIwrQdKRtI3MIHebM3RftfB09E
zt/APHcKXQPp5YTna3dwv8fCiIbx8DW7/0wRhme6gvrRWZ38addI2Qc3pc37qD7X
4M0mCGmofGrTt3eB8kn4Doeyu28BUla2clkqlMsWrgqAZUbdy+pvXPcFu+ypiqgY
mKkKCGzfJoSj5HwYWjJcb2jL9sALIkBISjC6cgMkAREEDuKBcmmZ1hCP7smmKcKO
+hzqiRcQOHyU6y75A6lE0LM/LxOxCsAIiElFpz/HKh9mRzYvoKX3kiIkJXSSt0D4
r0PxQAXjzjOUFXC6uvsvqGrmoFXlhmXA5/NPpdORgq0kkftf2q2oHzyBTxTysyLN
BYmdJqFE8Cazugj0FwBki5kb7Cv9ssSYAvxjbuBoEak0VqwKyjmUYcuQpHInhHhD
2T45i0sm8vaOvKe09fIiEkC2kam8+mXdTaLBxFyp8fetgdY1WZDOq/jzKatatqLC
0HBeV/U3xoiwIKFpd6By2a1B9f8azVWiVorxJUrRM1w44xhVpz9LJm6fRuJHBDAv
YrSM7xQ+TGcwkYTXEr8qnAyfPQg6dX0OApiOUPh02d2AJTO4VLBSMMKHsaWNw/K0
A1h5R2dh6cKo+Agw1gNCxwJ1ZNVd79aDTnTizgqd23uZhWxERyZZNrYr4i91ZdqP
Oom0V1Ih2d2qCpLzKEWB7jyATju0kBrncNEwto+pF4hdUh5/olnUnCTPOlc5XhoK
VyAKaTA14kOg/dq0i86AldQXn5EehrmcqvZIcPI44gjLS538DVIMvA0gxMufn2Fx
3DL1MBn5qSC5SW3wS14xa13O6RAK2O4HjA7+tqsAx3I+hnSFrZkKyHtNtgCwWUE7
21/zgUVxqOfNqhNeJVPLVPDhYKkWD4oZz6d0rw7UoO5poQqBQ1lsz5u2grSrVHeM
ksI4yese/9uL8MP76DviDkmL9n7hrcmwDpME2iLfob64hyjKHEIq7NVw86VBxYzG
goMNXHt4yiI5rMuxVKQvsKHzQQI1xkb9OBE90fLT6Erv7mx6evcm1FukakAsuTaW
BacjtD9CH5QLaVnwgiUovQWOIWIR5k4nKQZDqK8mhkFR1g++TSkcxvqm5Gzvu2Ta
1MBt/FDWRmkXlOR8ZdvqclEZm3xK+akglw9KAZZhWlYqkM+OyboZvo7l7ZmHsr+C
3AoJIqAweO2WYRgK24zKAa1Uwkl+kjrhAFhklbeELGksM2h/jHcJYv4BdBveOldp
CbeG8C0E2WycuIuvpyi/cju2qNnsOIF78x7AlWKZFbKZjsvrNkf+tpxndKqp63Kv
oVqI+fLuxN++9f8XnhgRfM4zp3ctBQNnYZbYr1NeUrrBzksCxQVe4IDw0jRYalBe
sNPPW4yfUsjWnsYgnAUUtFeJCzuALrTKwUG0dOz8Hd8mfDdljUyKG9PXt5OaaUDd
6slpsfE270M6r0IiBaPdIAUZ1pvYf2fKntsaRqnb4a4alZwbMrKLRlYxQbQNRBej
SS+SUo+Uf0m+/JxjJ1CHzRX1iPO72bg9CnZWVdsCOAL8k0NwgzUGzeSeL7licLJ2
ik2RoXgy3IGQVPR6Yer0HpLHo5m6lxtd6dqsZfDM+ET0DD9L3lEotNPJ/NB69jk0
lUtblzmtx4LPFHZyU2gI8PYjy9V0sNsp/S6Rbtfl8wexImkDmixIwfHXN/Ytms4h
sPTd7O2IU2nh3IoUd89TDiSeLJBWpcu1Er9I2YXAwhcoxFY9lbUM4ZLxwCJ48/Pa
XoIt1DZls9ChOgZQf1Lvz3vm8TQQl4G42WBARBCzAbuxt47QaEybftrZfPN+1Ced
Q4YlIMTfVbSkiILcW1EOSUGH249Jq4TRKdp7xn5wgrfME2L078WfwD727DEGyWPl
W5hNHiaeC2RVTXBUYHfYXAXa4SKChtwkx5VU0iLA7ueDTnNOJjvYXjRZwnWqLEi9
h+tJWbK3Lyn3/q57yzwii0SNRcEoX35RTDBznbls15KUfUgLSvDTDIGEeD079DTo
v82a+00XrEmr3zkWVRpETV6Urz/xPsDTEyzwXBTAj0HPYCLiXzGWRQdKsk1m5OPa
gsN/mlsW9/oqrmNBQLzxujGUgqVsMKzddFfw/tGLWwBpQvYA3e+sFMRjcUSUIwMs
resEC2wryLwFu0pkp52fs1njOnHEmeOt/kAFZw0THBOlLNcqJgIsHkY0HPLVIgTb
aAHKtcS2GVKE34FwfaGbM480DlCi9ae2qOBi8jEqBrhh2E2dknAJfMVZMjtTBIN2
IVN5iImM/bRzLvJNuh+qBODzUWIEFiCEtpJNScoGakxpLaHfEVekROA5cIXQosXn
H4QiXU791hN8bVbwDlT/OLlYMo8Bq+JkQZYsA3CGFcwt7zQEAGST+xZdF7/7vTW5
cEq/LosP5LR1nAtKfVDrG+uxCk5HZ9qCxzAIWjy5hqEMsWhDr5wR9+riWZC4OHte
IeW+QlvOvaRZ7o5QJfoazlh6lVVBwFVx3u79TU8lKPBdDSva7wQnJiMXemLuZK/0
dFi9wEDy4ArZbzFXqfYiGa4IeHDinXUXt3ahL7b1STS4kdX+Bwifb00zZt65rAPm
wUfgIK37wc+CDgBo/F5FsgBhrd9A71ldSMBFxHTDjM5SvYsztkbWtmRXYLSdFnhW
PPmbrPcd4a90aclgMyLvBOmJ3cNajLfLOq/R7wHO0rPcQApBpt5OsD9JpxvB67Vr
7F6ACIOVigImbPiu9cgkd+0B/pztefNfPmLh0L5guBmB+S4NxM6nngzxTJ8ATiBL
jIeIVHXrkdvPKgeioi8PzqbInmLT0jiS+NSSgqjKqjYwaEtdtELomQ8I5MrVgj4o
DnFplpMA7u8ngIWMLOUOMZFtLkkqqh+aZyO6tSTRWR6lKE0OQ5iZCp/3iMgjmOe2
PeTLpiDgP1TSQcra9driFjtvFsikaUovbRXAtlqoRI6i+rnaukEOnPPgGm6GskqB
e964wmVl24Uzxkc6HvwRzWtwHBsJhKfuOON2pBNXWfGhxT/q/v11I6JwUJCP5yVV
AT6zKC3t/WPOhaY9yvHmIqmreLLb+9n2vuoKVGKWAnz3HA7Ar9hBEeLwgUstT0Gl
u3/FH9sgNgkmqfKj6B4DxDVMWt/5hFVjFT1Ty73C66i3UHmdhmwI6+nnTHVDtZlz
jvYU5NxcQcI+hBJNlBcvdv4rtnsOdm+xb+fwkXlmZgC6DaPEylCljKDgLczqQq3B
gWX6580alHGOPP7JaDQMPm7anVnn5MYgfukkO19FqD08jCJIZ+QO1biSp87ZKTSX
z3kxLYzLIflrfgv14DDRqaGcgVcsOHUU0jnEAEM0qusWRCz/JWjf87DYo2uG54Kt
k8xJWiLPSpOG7G8aUA3/sDZ2Rwa4ZVenxx4jIrEecSBDCqOM8mDKH2TpvBt7/EKC
SzHdlXxZWzwLRO69Uw6ejvhoik51XL3AO+TXLlVMYBX/SIX6ijoD1dhMI9CqQyRZ
Ih2F+mFbURoa4C7H+Ikdfjn8zFsftLV77xr0mj6fQtyuIQfzvxkJlpE6ctZUnXI9
3SARQrORTF6mM/SkxlwzNWDz57KQJ1P3YdMOf5QswTRFxE5xJ4d3Rf0ViohsSWFO
I3uTvVBiWNfKRXIYL7woVL8N/sbe922ZLa6SwYuxdqZNOGQwoGgUJiVGSG9Yc5Xm
3iVyqEqCETcmn6KnQI1qGNC4K3T7plg1Bn4ljfVgdchbRoC3yGa5AStNVrxEbYdD
+TtGAvUcr0xKab+roruURqosle3Y2c7yx/4d0crnTjaQZX6amBnnuau3XIPZiXtF
GDzmwzgzMGeECCt61ZGkOE5I6JZFLIjJWHPh08srpwMIPMcNQTUlg0sEc045q6nu
xyzbJZn5EGAofyBsiy84eqHh35jWI4f9D2k7AGZTwNqftGJ7ccxRrFrd7tPTlbyj
DwbFqD7EJ6V8vkl0mxKg/UQab0HaxiN4nWIfCsiAyjzmEl0nS+wVfatgLSPOnSvB
XyiwwEU53hi7+evV3phq3bSoUiKmc1uheYAaS8/dG9Wo2ZlgI5+zs+bbZeRL3OJ1
c2WRXUQl+D19k6mmIJBAmyTEKU0NFK0AsnAdcoEUtCUGZJ0RIULC56y6RjAM74k3
LcmcOx8AYgnwUwISVHzvQIlKZo7evQYybrBiDG8VWWBxt3JMvuEMzbM+9xXX/qlQ
5NNjz4jvH2bXXn1xrk86Xh5d0I7PI5cJKGmmdlDCi9uEnJbgPbSbSb/CSkmlR7UR
ZJXnwXTfIWcDasQL5fh3SEJxT6igmODCFL3SeI98qXT4lDSNphk/kUQigSjNXUfQ
Mbcf/Z1s9g+Th9aBlaxa4N2G04DpSulUe5nfeNDndwdPgiUggQsV2orMwPg2NgKd
YwBcViyGMatVYnqYfNjwKBZM8UJHl7seS3JUsKLEjlNvIYPlyM55aohXY/q4cq5d
rXeIpm5gC/nfiNPXdBBwBS6F+Sl4Mea0XIKq3BVytnQYkL7rbp+38J/P7k825fbr
LOpU0/KTrItQQqXaLAZ19Mac0Fj4knV0N7zKRoxbPWD1H5Fe5nzsMh+6Dn1d32er
psTlXTgFsP6FMdq6QhUtWYxEQAh9tLuSD01s04Etov9ab5+UUhpltcw+9YF+w7Gx
Soc/fk2p+Un0aYiQxVJViBvw2PisqbWq1tmMocKCimhOoyLqi5Hmc3T9RgoWYGwu
TzM8YKzF/UE2uYpTUXYjT0Xh9kaJsda5k0u5NaWY6Tlk/9QmkJOnD3jq/8rSHmHq
EHOIQidppx4yUgfRA1v3s8FeX5dqDLU7MDaUe/Bj28lg5FHAgvUUZ/QjIwnrrPF9
BiWBi7Us1xzU2X0uSx0+w2HJy49H7uPNdrGVSETfDiFUVJIqSldHuoBoyOwHP8HC
TJrYdQGZ6oakzHWgSlR2faWxqIUA1+4pxd5daTseSDZwmk4+qeyYIv2antf+5Hty
t+diD0m/HlJssBicNQKirg3P4yojtz28nKSGDIfGEzA8soHihsD8+hw5oJ3t7d8Z
V/Ex9Nd2TpBUODiMYvWr3JOnsmX4IrViayNQfmmyN43SZykHzWa9rP1yOfuPf1Om
ycy0TO+Nd78xjpjMjrGLap7/iylH8GhXfRzA50hpTyMw+CIXlOB0NuJUKuqTjaHH
pzN/yNwquxZpw7SSjWveFw9RMbr6LN0c7VAK+X87WH0WKXnsVQLPe4uu+k2LQyya
QGe9T0yjLEeKhl/77Hx/QIiSe+aI1LnePzdlSJU0JOnjRF49atPJn3/gi8+/IZkT
a8aYRW3JiUqBucRh25qECqBqnEhOtPvTa+5SULGaLUBxpfGMSapRND4bdJknswku
rztpNUwYUovTvmniZ/9YQLuAnMnwpybd9MMnUAamEfVJDNAUh1+wYOj4a+720+xO
KWyYElTLXkPrwgCJ1oOj+eiPX7swF1+HWsCoipfLivBcoibicfGWPaBy5J0FZkdy
51DrA0k+0Yg+Cc4NHS/JYLFAeqb1woxH63opMZmo3q1M0CIr0/1BcFcq/YBZkXR3
6g41B2Jy6etynooo+NdU90kqIqlvvirXsoY5rvGSo1w1dh+i2gvbyUB/vsXmzcBT
Ow6y4/JUJyyh+Y5J1Vou4emRWkUhraAEo7DuBjmDXrAm2weM8wWd+UbZnv2kx+5b
nEAytyBwOrKdjdlEo2kljXkOzvO90FGvnH0rn+CUv7ThsOspD808TQL1V2zjIgF+
FjxNqQ/IMLMHqlbehBPPtuYsIT80DzavI+ZPr6BKZjk86w+Geg7Ayi63Xv8zkxvU
mvlGkff2MyS0Yz83o8J2rwyNXa9NqTu9MBL+vqGVx898JAneJH8IfjA58xaCjemT
L92sG1hv6KiIihGvRkk377OLdVH08g57rAYBWLNMtEDgqyVF267uWfHlg2XI9hMu
fv8oc8S9TOUawP+60dbaVA6B58bCknfGOwl8+1bP/AYtzkVxpFMiNaNucwgBjl5E
AbfhDbrdqgpQiTPyenAg9iaz+M/osyoMCd8KdbZCWBPbRGwDmjRB0gY//SUuuRdU
rbcp+8jTMCAeCfc/pwKR3pvQ6XNqFS9uz6mfQCRGTiBP2uDZaHgq/1OgU5lD4owU
qYk3TZqhXLtynxmLpNddTftxWpRHXOedMp1co6SFv34rycKWkT+upqmYb4/PuErB
8H97WKhscAIwozGXZVkOl3Amn63XIlUZb6S6E2piGS8oCHVm1niu0GppL/C1NN/w
KsdjmrJazYM4ByG9NcaKhzS7O9OFl5RfHXek5LnhjkK8+Xgz0nizBI+NM+YJE18n
V87sANGwMGs6kSk/UaUmcQK+wbpm6QWarBAGf3NNTjpHfZE7Y4hkLTmu90jTnKEc
hG635HopVzjCZs6OwkPjCYgx9A3JdlgBDJv6qiC0VML7WECn2bqAJZCtaqh5AoWI
SQMD6kgZHNDUNvhEnyGYwmQg8FdhmtUniaAkqR+QLsmROui02jVyI/xHIEOYwvbv
LVIGWYB7coJ0NDPwDS7Ybr9vt8TmFaTAqYa/cM1bJBASoqTLdGsPWSgsnus1CJ1c
7oSnrFI2yOHCGpYz8KSGOLU8lDQk1q09GkXdPaeaj6TutulwWEcPtJp249g+EfVX
+DhHVztIy9WepUavraKbaV2HYLU5KxD0DOo3YvuOZRJRKcoVztdPe20t+Syar039
g7VP9ahPTtV7nLNPkOxe8N1TG/NgOx10xNNCodItrtP/ngd+pmYyImjpDPEQ4sqx
a7dS+R5ZQ7MCx5gr2Llg6ubYtwWp265wDCPrV13QaGZXDKt9nlnZCOZTS4dylVLT
FsLPzp8KqGTBDgRaO5Bjumb45N8I74FYRbYgABqIrdC6L5STXDMd6E5AiAVPLrW8
u5reZXDCgP+SXq+P2uXkieTuX5pBzJTg0arIx38TMUj1fBGNREyzKsSI3YBnG6Z7
JABCPJoX+V6l1nasHUHkkM3aPICGCPmkVjEEPTtgBOUUTPmQEbCAWOcriPeELwCH
2uwOF6mbjf2nADa35zfraX0GyzQEwKTLjPfUm60xOU0qc69B0xSUDtKEfdW0wVjP
zMP6eMi3uDrJYpzSfjY41OHQAEb8Be4maIvLTxBZtfcO/gepzZwVTjjzUx1qy7nt
VHX5PmIMuwPpVbz8LeoA/CK86OwdvZ623zRMnAF0VXHiMDJfQOFfNac2xhkLsEjK
PpE6Bp1V19vBOtBMUbPEuwgBX3QRmi43MJGqSqvF/z3uEqowXYhdqku54hKLNeJ2
cv1m/TXSXFbHgxxM9Ip+yVxUCT81OX0pGSTJRO++6uS+IFAOAxGQnPU9ttTFwR2A
UzBUKSJPT85ab1BZGOhFSz42Jch8H55FhPaKpB6PmtjhntojdwTjYNuBKamtRlyy
RvHMk+AyLHJ3qmQcqVXje8mGWZjfkxkTi3snX7FRUPM6BHHm5Kpzzu11K6cZgGEA
3giO72BHO1hmi0pTnFzjX6IO3xqsNPuv58PL7NTZ6d+AP17wa4CAzcnRvaNHsXP0
pIGg7fM/1j2YinrSj81Ea5bTMKx96/GxP3Mbio4UXKw6IkYStM9MumL6ftsnSafL
9deWRvA0UsfcrfoGg6bI3M4YLEvCon/Hyq02gbxh+2YrXE4ad3bR3SK2/0vRi/58
OkfMt3cTD7R+Vw7iDkFL3/uo+HV46cUFVGm3ddPVSUifwNtR9ABRNv5hq89DjBW2
rb7D1Sbkbk3bTZ80Bv2JsBec2mMGO0IWsiI0rt/I97tFXQWB+OJ3NZhkPtLWRqO7
MetyDIUz6UB9jW56PpKJETP+UJIhbaP1Aks6YmyFcnpHrwEXLLIzbpGwBuorLc1j
mP5vVTPI+hTCIv0/kgdD0R8H41D5z4s20wmnS9GchbkggYnFM6a1pGwFFs+5ikmb
ApUJBuEl/iYx9WGJd8nX/g1XZyQwNw7pRgTFa6BcnphDyDLEP1CVZnscQlHSoYgt
m/Cc63HJpYiY3cEUENEWRB1JQ/x2DckuNiAXy4AYNM/BtlpbLDH7V1kzq1HVhN/S
IQYUtzNl2TgXavzIWqilV2yWQZsZUekmyyOSugy2hNNNusSBtMNdSql2WFAVzT5F
92reiJzoCXTFXtyn2Osuch+GORGooY2EuJYE18dl1NIU3b9bDvvp1u1RMKTckX0F
b8jtwBqhwFrxKnW0LF76l3XD0dfNBvJh3Cytu7M3rdPAQVtCOZK/vkqO75ZmSQVW
cDKIT8jQO4IkKQUmpw8ppMP0WgYOCrmrlPFBsWuegA6H98LhLqpfkDJm/SyL7PMm
GkLMtOPag5MOmdwJ3u55e4ql2nbkNFZdgGqh7KD4nh+X1AEbaGoRr/Rwyarcu9vW
vwlQwjYO0mNw7WcDVJuzOT66pa+V01GbiDK4zk9cLRalDbFqrwUl5IGI9qGN5LOg
/60dF1ngv9TM0wZgSGgqj1YR48yPFlmmhN0E/MiTG2cbGMtCvOWNWbcoKOsjzZPR
JxVPo429zl1m4zrTIidHpSdM343MuXVI8EvyUKyX8FtM0iV+wYBBkQ16Q4LtnUlP
Q/NojhRt2Qc0My/SNa7nRg/V3xjePuS4bv0OFAffGQ3tG8EASV3wg8OPOmhwSIW1
HaJEAGMFSMU/WTkDvnI0vVNQtHAFD2cuSBEBjFL2oeoEAfqa7x89RPyVnvAZLFi/
V7EpJoHIAy10TSZwLov4lHdNeEbfm10Qp6G/PkiZkzbmZxcoVrmJl/EHoCwmyTCX
dAzkT5KYhZtbJGTw9Xm2/9YqQxk5SIx6TxJNHG0SI4/raabZ0JwGOjcUC8vFuYtC
wqUECO2kMVICVgVWVoJr9KHOwfX1XBvOKjgyya6C44CDcLOu/rF6MUmMvq+QJVRp
V/agHuNzcI3CEkr8PP5ZQXG4IxTweC32wvMBdeH71+kS/Uwd1T5ZwIjcAEfbVBPB
UZ45ZPuZch91ojdHOpLz4vlzsf4ZkoQYO8F9M1Om4jjH9MQm1V13qWm1a1YJ7cXi
24woyrYjvImUrsvRd0coV/WFtEB+blf9yGkavRG/6d4BjG/p9Xx+p2OJwJRsyZDe
ePsaqAH2SXxGhUHgn/6SJZY7eMQTgovPXIHPiFDkg2mpd2xHZdqau1PUJ83SpMRE
uTbExwG8T8+OJ/Ylycw7j1FA5iPcxwOTpn3zb1QyWBrz91ivjhKFGiuZIqoTcsAb
7dVTdkfKbRBraiLGx8K3dfdHaa1h/b/Z4EzUP7m+kwQGyJOKemD6v6cgsAaZLTl5
a6WW+F6ZM8LW5g64Ys5Z3gsE88X8M+I5FPJGGKmw1Ik8stZ5UfY18tjiJccTTNOw
GPuJEgffEyNFSpoGrBEqXIXVDd7fO56mkk72cE0+N75PQbibHUgb95e9tCuE0HKZ
a9vq4kEUd1JBhNtOKoyM+2Gq3NbeN2aScVT7+z2nRUmKYcdSHfBOK2lzHq7V4WTz
OF1FLj4GIAGamZsS0HAHTjhDkQNoopUkZI/LRvglDmn/PzyU7S4NGJ5tJsNILR33
TVTH4SQ6WdsTPum7Q/dw1fgq1WE4pq2FTiWELEjmaRphmMaZuENzpR8OqHgxgG/c
/ttazwdTpjUYnM4HiAe2XlyFQ/FVskpYP75YwJ8yf49soDrDmd0bDc+ChVjXOy4D
5RHSyut4+qdtOH3cu0z/hToqDn7cwZNzIgvfNU2iRg4CzxhckFjNCpcdCkuUByDh
FtrXpYFqLVw0Jj6F1jxsdPkxlOT9k3gjT7e5l+XX09ZB0omrcMZAB4RVZHbq26r+
zFxkOYnIeNzrdbOHoKQdzfNc+7+oBmnI4kOV4rvxMoEDyYVBJt511iMU4rJFqh9v
QnOSKFuB6TCSJOTgUCQuR3NlsdLCD6uaLqRgNNu6WENynoFO8MuuKqSWlB26rld8
edOE0ajQIjOEfVL/ep8alovUYZJ0dg9p1ajvoMzYofnGQi96bnLGlMxSi1B3aUn0
yr/WFC+d37RULeFVTSaL1T29az7+JlgOH+qyG5k1Ll45eXLFiMc9kLIo6SnT3I9e
EykNV6mIX3Fol/JSXks1qIGeg6Q9Iy3coNIHC7S5hmZNKIpfV6RED5bGsBjG2j5S
MhwqkuvkqLtL/ViLsyLHgxzjtPQMTc3ioZKBheul2lhsf67aAgBFK/j47ttDBlEQ
abTlFgtvFZaxw8tdUXxOKSlpYijXvVnqmOhbyDk0sDkYLzfQgZPF3S6ZHwMsXEr9
HU3WZoSLurMxhGvi3saYRmFiJBOW/d7ifnqFupfHOSlUN6a+nB0bPipiFZWU8xEO
EGEf37lhb/b5+NJAZZ+J1z7meIHaLDCkWpaMgOT+bYPFL2jyvON3Zj6oqOABjIJe
m1jPNd8Z92+MgP26zOmAXZLX1LNd8RG0ALo0YhFK18OcjBFm9npsT7cHG8rctGXA
562fK3yJTHdfWfDEnSGul/qAKIA26X3HyQuR+3KWj6ia1GnqlWEg6/4zs83Sem7s
NwsQjhdfVK2NrH8UFN+ppcvf6P1PGY3iYXiEDOPVjeKNud9VUGLf+1/c9DXdEvKk
l+lIINTY10s9u3A1RF2zU7txut8+vM24aJWnFmorg+I4xl1o9GsjfnW/013f0GTe
J76fO4+8i3wiQCJiUzSwGJs+lERksqXmhw42qJUPnYJHrlio28JxoNJl7p+ge8+m
zz+PFnvKKx03Q9VsyPBssNIgDVg+BFpG1zkSeXObGoroK3zon8yT///al0UoPWv2
vW5LFHC2aUKnFoA4GiGxhyX6Bn5O1TlbXUTq9dLgxDbPMzagoYx89AQAQ5uVGTdQ
k0MKf2ZwSMHF3TrDjRZROdBXZAGlBFDGT5sdVRei+/wewGWsV5POrvuqA7RKDXn3
N0LCkoaRGG9yLeZEmB7z/6ky5xBmYNUNFmCq1JS2RPs2+SiSmImJ4kSnF4IJO8X5
r29tFN6oCNEO2LTipjKBWNBt3E540PGL0znoRFoAVq5PNWWOO8foJVERHw347yXF
scIb8vq6xlamUVjX+j9CinS/TiP+kn5dGHGgOygUoB15FH4Zz8UjqijtetqAAHBV
HBj7ioK14LxtPr5D8UG498Fn76+NLqI7Ivl3TEX+Fdn+nha/j5fU2F5jOKK3abmo
ULXIhLaaSd4i3WZ2t8dVYvyYg5O8GGuUZgPp1+MLBvoWO29cxRpsGBkVShMz20nt
yPtopdfPx+bBfvgXQAZPGiieTlKq4iWGwqpQHycrHtdJzUQqTEZIJ1WZXrw3qE0p
PwbKylI+1Eum3Z7eFCZVqyD+n/BKQhbcbXp5piWVPtYXspF8cz1VAVYUIWETbAVp
iuS5HJhJvBLqVYIwDR3nyJylyWhxJwl74no6Oqzfw91D6BQda2LP1R+GZ9t2360c
YigjeAUQ33joFR0msavZyZmSWwJsqEddgz/11uzoVIniUDyUbGuWAh/7IZ/EPD5l
1qKjtHViQ2pV+8WHDgkVswwSPbjl1u8AzUsyeUBZOba3fw9n9zG1+lgKQeBnobxK
3ByJ04kRp+WrkH8HTP3Sq04Uix3YpybC37Ylx0E/66OQDHJQ0sVJwd2TC3/B+lC9
amGWxYgFb7NlHT8R2Yxp+WMvmy7bFsM45Yojp2tM3+pN3M9X0Nk5iZRAvDQRNEXn
WTVVqoTUNmKaIs7rY/ZNT3nBJVlTsQgOb4VCn3pN/F/Br6xfXHMTcKJp7HirSH6I
XDf51WKTUtu4wwOggq4JWQIwkQPb12nSIxbSrGLBEFpUXJTSHnAOdfva9BYv9dSE
qXjUCioYQ5TIZVDmoHDUlwvb0E6bmotfP7D6s96xj8R54MhdrO16poTL+WSeV5Yx
C1DYbAiSsUzSc8vjjFG6hjNTXODqcgeeIbVkHvAxqrLsaAzIb9MDDL3R8mhhJJuc
5aS2yGZNZMrLgPYGyjBSlMLV7PuZTaoMARt8wdft1WA7gBtXQpemBFtxAWaXCFaj
70FLsJoNqTEbOws4GDGljpfavQrgzvES53Ea9zYTksPqC5P25WcevVX3lLOikhn2
JQpI4xrnYewsu5sX83Jg+l0WVKkmi/K5Nm5lc0dhqxVcu+0dGsTj3A9rZEwk8SXE
a3Ks67BzDn/IyXZBsHJztzh8IlNB4xnP2Q173GsJFZvwVKfpDb4dfvcYTs0jK03M
N+Q3fpIhhvOdS7bUgWZOiX+vRP/OyT7M797gtnvSN47sILZ4PjS9KjqrnQAeZCn/
SSq1ZImfJ+4G93a+hypExyGRkm4t//BDG1ePm9PxxInmW5wl5Bt3x8I9xYgAMe03
MxwPX2fRDvslRqCe3sPBFGwv67pLdBhVeEW7KIWiBTTUqdK6zwXU1wpR1zicadcP
A6gbf4yVtbAtFF7wUVkfsafB4H4CGuuFrOlWOmc9yWBAdNWv5lRTYIho0rA1McrH
XZlJdEL//ChwH23WxawJDjOZOkd46EShUV4lpeIDqs5HFvtlht6jbH9SAuL3gghj
ze/M8wqPAsmcB7Mj8dTPzoHj00IrI0I0Axtg7yCQLvvSdLHiAMr9DhU2DxcGasEJ
SrNZjugI4KPEkt/2JLcWpdJIfxbiPkXNZxZgwUOnUnlwKwrQfT5095q/NMVO1NgG
1718jb9FaCSSpFVsBRqTkzzUsN8cQVpRRhg/pgLroggvF6/qWA0028wqFbB/WGM9
l5XBAnlj6r5ODLWJQpYF83EFJBD6H+VeMr3IdACJncgvdpOBthFhFKN/gKM7NOmX
Ix2MXX6wkNPEXRGInIQchpZRKsPXtrfOeOWYsWU1dU8s3rn7rAQVM7e8vL2685CH
SMcInILLzE5j6uigGM/yyTBDUntXxu0IhL728jFRbBg2NP5G22opkgj95lWnDCAO
VthHXDTucDzUCvv573TrsDELrt157RaTxUlb3UH5nMKYgJ+Uz7hJeGZIH3K8qHsl
8xhJB55Owm7Zm7vtqDetvKPyiIGEUzaB/FYKv7HXA8VsxnOrKj5ZDrTGICRETUC4
Y06i/Rytc9BnHDS7HktbJ5P7qXiUU/PdII8tr8WvGEHoBR59khD+QpWT7eGztLfZ
KCJccUvZa7rK09ogYf2iAUyckYz9JOeOYPbny1Qs0ZqMAvJO4MSLOGUhpNW/JfMF
QOCLyYB1BFG4A/asCz99irPzZEY3niyfZWWuFFs7M00/h7P9/D3rfd70U9OWCyaD
0fkQUvZHjgt9UOZCVe8uo5wzpqg28AK3YaKiErhiRerZMZigywLNiPeD5qj7jmEM
3FsrZbQ/8DIORZWE9pd/fkj3KzX0W0jTFv9jupp5ClATnhhzIunTssl2y2BMwTa9
hl3IIlLfZWPuG/UEaEywAgUao7PEZNxhQFCnaPSov3mNtt7E+YTFWswAdwgqHosX
tPH68J4pXlGqLYuARXrzJ43S9NqZDLYA/0Zf+RQ+4IGzf0qYpgIqFFxTc4aCtFIM
cMMCgTrvdiaa2a1mp5JhxOjyD047nVQe+bZMINGy3wYTbuBJ4JEAcHm7AyvGuw6+
DjPT9GlH7Nr0aTWR+5/zZpOLowvaaLZJHvgCW3Qi5zu+lgYR3EQ0aVuVxoMH/oFF
Nchma0wvTSRP1I3mAixelHQvK6eXWJj7qblqej160an/+QI9Q4Z9Ekt8uNyK9XfK
BDxP6KhYWuFh6/6Lan7ScmOo7/7aKrgcGsg8EB/VhqEdBXE2DkjS0Als6bZQRgMp
u/dZZ0RBBFLUK/K/pBrNBOhFu7PfC3kbOdnAjnCEPsa9lmmFIyATBJzoJclPCcZ0
x/O6QFyel2KVgam5CbRo3a06FBEqDIZ6XGj99THB8qFgCXPovpcDqXOZy9oelnjD
XmEY4GOg7Pb0v3H4gETOFftiOc69J4PaY2jTlXWObV30R1XyynS9AyM0RhCWBVYS
OfnqalyJOG0H5YtyaWGicU1MwxNHcqL6BaqCR7UFN0USzvu/cpa8smqsYI3Qi2Fi
NXzM7G6X+LyRMBX+8kXXYTlcLgaiIYirbHyAQ/5R76nMh/U1HF2EwZqkaxdxgPYI
hhcysTsOAMjl2EOk8M5gFOU0iyOZoN7NDwM2LtGT6mGJUmLKosV12hmFzOz7Wfet
z8Cnp3A5AjqitREwb1DufjIu9BT5c9jvHc0q/4ps8G9mKFUiR07rALFg7raaEDct
EejU0tB9fN+wui6HaK2O1X+WkqsPNeQLdV0QNEyDXkhX8Lp6X2n5SEneC01xFyTU
Kfv3UnpI3gCHzwXgPUnlpICADekMqi3uNTMYvMIVPOwQfmUL13AurY5gdid9GvSr
6/mWRDxYNYPqjxeusmW4VvppOGBsjOn28nA3H/HyGxhS6f+Yeh59sHqU/BM26pT6
7dwI9dk7YWNbMNoq31Y2WmT2QaywAtOcv3oF5O6TKZL4utb3usAd1rP5UApY1uwd
S4syMCtRLUloyu4s2eCHQEdu52aVc8jW4D/90PbFMFmGQd1NT8x91gvGgWguJyEF
Aa0apYEBCW7cZg+a2a+1ZuzpejtSQsM4IDyDiCROdXXzs84TPPqxqzPNkg200ZVf
OtHO2gTM7VcKN7ctPXBEw+gxMCgxKwCSM4RYSoHqnGvtyCcleEu9AZtnESliAeAO
oIhYZcQRp3hrT9h/D85RTJqKgid6ZLqT1Js5ibmRKO3PeFaPwtLquI1TRTTFeYxk
0VdNJ9rzI2qt/D5vlnrCt0V1CYuqHRKUvhMB7oB4iEzOph9391Ut7/LH3/dQgUY4
C5nxb8nhotpKj+W0FyqdC9wVc/9A+7RVAcgiY+VlrHX6q7l5F2MezErcPNm+awWc
wvZjZxEu4HDMK3hsxxrKbA==
`pragma protect end_protected
