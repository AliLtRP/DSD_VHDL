// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
Oy2Tg4fvLzEA9RhvQM+Rb09RvBpVzyKbT4ZySBSawIKiyQlMvxPWttW/bH2uy/C4gAXZ5LsUb5fa
2fMWKmp6XPr+rRqqR2qg/W892pMinwW/xPQ6vrliaFuo41gp2vWopPkFq9NaQpgvgmqjLurt4Jbd
SM5ZjqN16U9qwi77NbGy+i1NI4Xyjq3rV3t1cUfM9cWLYeTUoIFR/hIkOkpfFeksE1WugMrI+dnf
QDt+CG3V6rCeLHzS4sksKV+fzF7d8rKxUvpDmcd8t8XYNeavXNcOzdpVxYpSrRmQX7qT0/Zj8CVE
Vnu8Wr/MkGGRIUgIaFKsY4iZzE//pLp1ZddE0A==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
uYLT0I6I/BKi6r9TDPqYt0Zsl4Y3d60R38Rug4spEupvtwhY94ZfHTkVCktA+hEmt0JePI3fMfFZ
pYg2iNdpx7dFmNerMkpp7ntxSxrrG1+QtPD7S36+g/ypfcRTKg4s7HW/AoAcjOpEFQBA+bd+eAQ5
3OAVOpxILYip1yVEYF7oF79DzSgzc+p6eWj0rx9D9HagxNqgV9a9hQ529LdkROOYiChGawPBGy4w
tqHCArSFAqRnSF+OZVka0hBojywfd1uoh59m2P9r23kdj/MyxqTn1gUNDfM37Dc1Qb1O7zxYaDml
sGJkdq0zNe2V4WjUiDnT/0DODaT7O4lqsyHBR0xpVQSyKr721gxyhjQ4M1KE7f5viDF6zGc90RC7
v6Qc0TIAw3IABhYuyq8qAWIV+2N2e9FjqubZ0jdL4Cq1NyYWPQhMhwX/TqmgVmZ5ht2mR1lf7EoL
hjsNA926UwMHVnjLPrqSNvI8K6xYy7UP4+qtnZP2qb8FhxKPAiHa9Lvz0ueuxzwl4odKWLZxrvgX
O69dYdHrjidiK+CbadRGoCh+hGvuuzrvTxXvGcc+INS5Ule9dh8Nd2/TWEHlmOwY9Ba7yy0EzlFg
zM6sJD9oRcJDpe0o0z0Zhp0pwwzopXcjTj6r0J31BnUTwqGxokwAksamYfcWkJzRL/8uoKJ9EYea
TMhs3+2xmUKOSedPwMQraqeVCLedPm3sUxeRSUjdbzGmjxQlBm/t+LxWRzBR0zLYGp83+qRYPuXh
8pvWlsyXWPXTjFC7+FQfGCdsTH1XTS0MMBTzZbORoz3DEEd4QN/zftbiUfzume+2RvnB6U9h3Shf
RyWpVQrEkrbwFaMDa86CcwZXVwLtRMd1s1A/Bvs/oC/zVh7P2Eiip1XrQNQU02CvrjRzEQzROU99
gmsFWFcJpIGnQigO97NvlM2ywk2IEzi83GjeJIPUqvQbvrDxTLDBV75STqe9Wa0RaqkoEPOeL/mM
QiuiU2Sz80RxlW0KOBV7dLa4TtR27BRUqAsCgFVa/sDRZAfretqSsSqfRvklDqr6iZaKnRZDb57z
ZfOOBiKmwfAVUP20DXM6fsU4Iqqsz/q0xs8b3Jd2hBb2FZhYiJZ1FQh1w07k6dcmoeLAIvZrF8j7
0ljejyEDFE4DbzNPMGiKl0zu7YEqA8RjihU8Xgbt1bXzeO0m+qkmyrP7Up3QtNzzvpL/DycPVLRH
a09535tWnZHIXG9vKNZEnB5+OvOg/NxlZQi1f/k0+JSqoDgl/168yJMmSCX8mOqHvIgCKtgBQ+m2
oYyrALbinEVCmMQaVx/TmRxB/WYzYdMw4pYxyY1AAq/YI4xUt3u5PIIa+BI3AKJnCsGZbr66SDHG
folGBwlAJc1TSF7eHUUZXQLJj3pGJON+Z0GQdLH+Mv5jtptgn4sMui2TF7FcrdItCWu2EFLTVKHM
Vz8Wx80Jkn0407FGrYy8O9OEQqRvC/JhuN1aHtRQ2ycSR4YZ1qfpI2zBfp6Wy5UGIOTyK8ji494O
0GpEwo1QjkCk5ddmrU3OMA28WgDleqYSQv2j5Hyd+k2S0uxku46WclXBCfTGi96mGsqAjSfUmY+b
t93bcEMr7JoTWj/NFRFhX+HQ9Jo9Ob+dnJQ9kj65+em8A10SCbY7UdXsQE1LDUF8HDi2O69IoscW
7R3sH5ID69mghwgVW6334NqnHxNJFpk+pYspr9i03Rvt9zLma6sV/nWM96q2F6gH5Rkcp3ZYDdGW
GzabHLuaEQtNcRGZJPWpm7dcvi2YN/9IETLazPk844TpeHEq+bA63bQR8jFgkkETMqEXFU+8YOmV
5J2AoDPZZINS0F7u4HxLn6s1klEDZUpNFu3pepZX/FYGXR2mkwfSsDzTPrUKe/voVln64/hWL5oY
t3uc29I9XnwA9g80UWFgutIJuk6P6N3Q3mBWtdJJnh0kteLlSVBZx4jYCCJe1GV3rlAul9lkxR6Z
WsITVn9FbpomhX61jYju7mUxeoHu81mHJcLCoHwd40rMkgRQGB0PXohu5B6V2trxO9KtrXV521UV
QX2WOx7571y62CF0jQ85OTmwtC/LPXPf1RA8VLTeXSOJ5I/fSvVS8CNB1I22lAbfM3mykr4tDGBA
lDW32i9dqkKJPakT1/uFtW1e35h1lC8t5mKujRIpADwU4Qq0qaHrVtgXfXJfYKHgd4W6O3tIsF02
Atc1UZ/KoeSSk2Ga9zNzXmHjkrEVSMYs2TdOAgua6DacBTAvsEr8cr3wdI/a+dFD7lXDjfA5opMG
SiI3N+W+3JglpLqiHPCb70HrhFas8T2gxrvzNm2MWolNN4U8ByvPNJv1Lz/HIehGBRdFRpisLF8C
7mrR+LtUZEGbVGrtV3BYB9yJcB3J1KVBhsL6SUJOZ3zPN7RmPpV5ZqTX2x8v4lbZp43Hr7oXgzXW
QhRGoKwFcOkoc3pPmWvW4Y3DYDZfIjl5WENu1FoTAk1mBfN3wcykGYcSvWXIQWvsE7/pq9A2sXKG
n8xrcIbqEJ/pBEsaVNH5iMTIHwnr5j7q5OA0PaXtJTMy9IehxAl28B2VpPL4jiGe89fitIJ5Bpuu
RhLvjmEa5zhlDEWwwF8bAPIJZh/mPOxM8MYZLeGmjYcq9wOn/sdtyIiIinJh61wEvhx8CVCx58Mw
sb8fPTyqkucDJSbeNEqPshQubFVUREPAlE79deAzuUzRMyYyngh9SDFT1T9R1ED82Q5dGlvLFGmx
H60UUJD1Dy2hPcNbm9xnp8LdaFCnmW5xbAAx1fRfDKWqKVqF1qZQQPgGOZlsiwdEEJC4mUkiebc8
6M3sl7wln6IEyzAJXuVy5/JXCq+YMartDZ9pXSuPTVfBpvWkz5aFZHvqqTn6D943lhfZOVEHf5TM
mNoZMKasQxIgtGu4AqDtpn6rkfdH5yeLGwPeKNdVrkMtfhqAjCMygERzZWQzrEd0ZF4vHr1J72bG
HjxivCFRvnqfyCDsJmAJMq0FpL+MKLf/coVoe7JJHy7+uPTmd8GpSU3kqZLML0eJ5aznqvnDSxZS
8g+6ng431o7LiGzM12fx/85MP3aRAeH4EOV01Na/q4J8y1qxYUcUbKQXvMEkDNZZBOMW9LJIHtxC
9A76BgeVn+CQr4aFMeoir3tWV1RPGi6u7vTu35A8dNAsHMW9rW5wPX/k7+OizGFdgQ0I88y3jo5w
pzYOQt+4vt01MuYlvql/YyEo/PmoRT0/VzxPwqU2eptW4Y+7XWQBcH4cKUKaODSvaaSniB1tanNG
rhuN88Z6kpmrZ9raOMqYQuWZtdgCn7KgLdsHsdTO1NmYCzLG5WXZinMhcXRuDq5p42gD2c5G6eZ+
2vzU//9kDN/CzQowrZPzE2wpwfhJZ+UdhnDpOSyCoUU0WYgKexYJ2YZh0z7ylgRJtSNt977IgAoh
Eh1Dgtv14xLJqJ8CkMj4fyc5WMGzax42XiTmqaOLoAkIKEKTHLhxENSSpZ2QdeaYebyY8eAsI5L7
+qjV6A6PylwPb2+a0gc1FaOMbHFVmtyhfYAyOJ029GDZYIFt/57yaSmgLqoyb08dx06aAfWl7n3a
hbDJQmwocq6YVjQOl5UecmIHhjcBkpByKaJtKBeZRqMs5S3t8lA958n1axLR9HUX4oc6zPRg6PKB
zF7khEzkgCuqwfmL+A7ATcFrfPhynakiFAMSK6vhoDVvkl1OJujbZyCBFHHOmMDCpoMhtmqjQPtA
saxhK25FWIoxZsEH30vOeHXLpTAJpQWvRTeXMKXcebEWFkLmILgJjcZvLOrJvveF8T5zQ9A6PVMF
n+6SID8PNwe3xUIpVisMhurT0TRVyLV8D/ax/GA5kVukd4rVY4xNdCXT4lUIfg3+eGAxHd6Ekl54
+IU0/b7T21sV8T1V79Hu4Y3gU1OhtfBTWgfL0SDvswOpGJuPX2WIHkc3KL2AXh9wjKCElqhJ+nO6
1XFtHEIA0NEfMdZxx6hAPOI1IvTzKSdT+BnVZ2uw6JoeUNG4We6yN2zqM0hYdLblBoqzv8siU0vg
41ov1TWGB/YyxoWKwwoLN8AJKKv8QESu4d06k7yZPw2qo4Y7Lg5M0AtaAjeBvmoT1rqJcDVfIWMG
Sp0M9Ud2YbXWcQ3fmVjvh77EdkNVN0t2VSsqIWoYQzxpsHgTQz/JvpDUs8Xk9fMlR2NaH8COgIQd
OLnBFOxh5yUSzKLIM1gPytesJo4mrfLsVPEOj5oTgoJQ3831gwemgC7vc2J9VWRXfN13tbxv4/vb
ZF7T+/+QP/bBI3QIFB0FV0jzf/O4VkyUFcIMRpI6/f3K6VNhlM6U66jGnZ9mKOONefqK7Jgb3x/u
VPZ10R+XDDWzqlgagA4QLiVThVvODAvTgiwNmpROmCN65wP7QmW9EtDgG5T0Khl99nHGnbp2cvmG
7o9qVYWdn7cxJxy3+UihAs0U2k8TJ6kxrPTEcp7oWmGUSke4BPMWvqNaOTWTC+PKXSaoeLe8+gT6
9spCCs6FEZclj1DBXrh8yYVRpSjABFtgqOnmt/F9igEumwcS4l99VeMSqEqQ9KUEkkrC1HLOw2br
wM/buMA3D+X4BzGmg8cNj8yJ128+v8QY6UVWzn9SX8+2eenLcasG7RvF3R/7vaiGFn4X4rBfEI8+
T9du7zfERaB1M+qxsnaV34hgVepFY6my4+cPjbaTR9rnW8Nxsx21hDfbFqcsv6ygho4/H1kte0Tw
eX2v4N8WHguPBIyQJMXfTSXMA/D7k3kZfH+vVD4em5P1oiwG17u1CzltsBskA5vNSXKSJFA5LyrM
w5xbpSzLW9imkth2CrRQ0E/nsdsPJyDQuujNn+J8T4JG8Z1SUNUqrrWuw9nQhPuBZuJeVVROecr7
IBzrE5ojlp1SXc1eAGzMl+gOT4Hqh0yEnOrSJZyx3gqYe5F7nC8/YbIKj9LKr/DoHGs0e3mV6TRL
r3skjOf3U1+YClAL1uRtd0OeeWhpm+S3IfJd6Y/56ImIqDLOrYv4Ck0FpmrXdApkNJyPdYRVfviK
fyRtywXKdf1L04KqRJy0mh3nfFQa7zTayNc8S0MBK4VT9DqX05m7nq8qhuNg+lwycC2GYGPxLxC0
GVJxyhuUzegIFg5TVsNTLsJTi9gmGrZlFSSA/geu3kKwU1pVn4HqqPCf8IA1gXJtr1IOblMvrkw7
36LgbE7NftxGV7LXdDTUteDqJeteYxSoWcaeY5IeqPamQSQmMWAP0CoybeoF2JyDuxLvsWGDsv36
8B3JYWKdOg4LWe42yREcXU7gqHzJjr36SEaB33cqFET1gmJBH9eBJQ8tj8x1C2lK0JF3BRNGDguJ
JdgsnRt/j3LaIJ7J2+dB0Wjp2rSiK9m6G6kHRmjJqG4ylmFTQg4kDRSJWMNUx39M8VU0j3jHctM0
l+Eh2jwCgPkug/YvyXnZxthI/3MwNCl8ZnJ/aHy7WyjxN18UouBO6VailaSR45YwYmwZmK6sKC6n
CxNEFGYy/mPRZTt69UwQPMhWmpRm09KsZUfBiRYVlVdlKfi7lwF3m8lLaEOdQGez6QpPK8Cxie9B
IK2neIMoZrKqoQIT8CcfocVAntquMy54SvieGzAyvzEIkk4bVxPbJG2pbaFHonDEfmlIvRZRRCeA
Z5pldSlSInzjChQlphSmam64I12rU2d7r+U+LPspckP10gGQGEb/sQKrFpI9KzlJXyVWyzLrLa/m
5HlzF3QoSZ+cZvSZuoOXDCTiiA0kG1Lt0/c+acoZI9A8iYMosngKfQRXKZoTeXuB8fqBykIeWS/m
1NoSUqiVE0lsYIw8Dw6RmTzfHue+jtzdUAooR+zJ+LyUULhrKQc/FxFDxsZ9gNawBB6ylkEF8/Dc
wVoLjwml60PAhsBtQP5BxC5MqGKfdsH7feM2cHCpXbPmRzGw0V73nsKtU9HLg0gpcrDRE9vU+uyd
VaiDyp2dzAZpj0tu9pBZZOy/TGm8KjVLHDZ8b6/108UClbLohGtjfz8ZX5QGhlUwAH10sCL12NWx
L74j6Z5/BleT/Hmx8Q+UhhZVepMbbpnsxPgcoXVtuphttg/MQ57LwXGc0gxCOpwHt9qtuOK4yjdR
+Lj9dL2AvwHvUnqlYv4hYElVOnxuYeDwj1SffO4RXAw8n0rJwnsspDCkGQ8J7cFFs4PMCzN4q2uJ
Ee5QXa5TxTB/VcHnn+sGomOQbsGnmtPlry6Muj+ZN62VEx72V7mSp522pCTuhwYgBlEoS92ZDfER
zLAEUsKVfirHP3GSY0EfxTp2p+X7ACQWM0PnKYLFNZuyN2vtN33Uc+yacyyR6sFGQjIW6Hh43yZt
aRQZDYRHh8KYxCddKuw1LhE/ChKLSIM3dIjak+9xecc6/iftiKqyUvSp7rpPqigAUgBHSJsFQ/w4
yF90iIEzlagdwAWXpZB9KKt/78FrBCU6fK9tpJy5WIhvrgvDoYYw1OOHsEBctV2qF5jrlJqESXG5
6JplXNHdYAYSJAnMNozNPBMbmfe42GLnGhSTVKtBCXCMhTChNk/dSXiQOILeNWuXIc5bF8z5rC8d
hGS4hpUzvTsYnfres17ksz2L7967ZmaVeo/P7N/ryTiJhFG9OfnNZ4skxvk951jnXmji+FsnlJxr
oRHggICIrCt/64582xNX/45MeHhOS/zjtj+7zZ9igrZho6Cb+2xBCUzAB9GkkKgKniab9DTYI6zu
ANQ4Udhlbm0bmm2D1wyPzEj1rxGppEkl+1nkeTjW1uDNkZrL77m6ZfSNEnTJHG+XJun9VnLVgFay
PMwP22WcxIkNwE/SrW/5dNxOd4bIVRbwVy0jbhFOMMG+N1W901Qbis8C5lva9c2PoHcCjb35YwHp
/SpGjjlYxbl1vhmAxTwMUzTzakFi55IBbZnYmY+dOHcpFdIropgPU1lyKJbf6if5nGE2vdGYcf12
7saWZnPNApGiVixYSAVy68HMoqcumK+nXD2QZxPru2ghHZabhjp33Udk0VW5qJRUgh76W1yutumf
HPgha1NhSDfIu7b562DzKBanjA15STqVCG0BAxQ1ti5DX0SM/0uJ0GK2X66AGTKoV/00BVw8kAjh
U7hAVqCk82cLR+JP2ylW5oWQ9Qz5ZLQy+dcBTOEq3P+8ApCFZtv0ZC9vZP2NSyjSw8FDa7h5diTd
MC70EQYeQzbW+ksFX8JwICGr8EBfjG523b1ZgooLOT5iJP1bqVriAL7EUIZouBNkO0LjF84XAolv
Soqd/1OIiph23NkhMPLeZfHLuUWD9HHSd/qjY1YMODMmcH4J6MZ8am4tqzLsgwuh9wJMZ7ESj6/W
rSexFohPZ1pN6cjHL1v+ZIjvy+Zo0WsLY1y401X/qjYJqvaQ06kCW5SmZMjmhFjKp/a75WA+ktfT
PJiJaxxUDGMVhx0yXAVwARjnKW986FFJ5FT5VLqe3DHyn+Q9z8oe+/wZbQJlbCIOvFpU9AWL/yKe
JsHTInQ0gJ1/8jLSRSik7HSV0uQcTMeoTOastB4ID6ETIDA5/+PPKAjpUqJiyLeOTubE7f3rMOkS
LGxucyavDkQ3/RFbR6iNmSp4JfkZ3oJn6kCefecpFzgKXqCzax1VZTAJaE1eiWmWlAkYENvKMnyu
14oV1L7DC7rbO4k6lklu2zOI7d+F9S8Qr9kEufw5/8U7mMC2hMYcK142DP/zKPfRUVba7JL4Auag
3w3rwhd5fi1EOdrk7r2qdVM54kfpphIeYMg30IVDaZW2WN/VNY7YSCrtFDl5CDkYNkZXumoFEi8g
A2bllJSCQUwpd9ZmMGmLNeaPYI3bcq281uoQ2ynLQ2R0VwAalDzNE9PoOEtl960h74wXVg7RHdfu
0qJVbKE3EROKi46GNpc2ro7l9ozOOgWJZ5ztIDaytaqw8qX9KzR1XdkA7+fMBCYAsfG5QyXzfdN6
JcZi7BjPUvC/HCW/LasalI3HjgFLryjoDdgPp6AChxp8oG29DlbS1/yRP3Zzpj54qQXEImUcykiw
5DPL35tjhmDyN/aAZv82UhRD5lw3gGBKYjcE8hp6gXwBKJrwXIJ38+QgT4JlU0/0hyXRIsvyob3F
bhe27iv/pDc7joaC5+lsvK4XHCcD9+6TZgsLeUGaLuQjRd1Dm3kaI1HIHW6zhIjykV76Qk7RHvoN
bVI602y157i0Fp6gZJ75FduhwybEiZHo/uc1tCFbgZYBlt9DSOtUxV4ahFWfOmyw93gfgB0dbpsS
NqVYoBorZ4WRy0h6VwyIwFyKIDxKL0v8vXqE0akV5ZTlStYIfkxxXQqglRI/0lMSCp3i0bNu+tqM
ZbIk5YZS+b3RWQJ0Jv4tXUsL92Iil25Znh3NCKU/XXJ3qY3hPman4E20fiLtvAe5Mf1ZpvzTg+uM
XQc4athluID5xyk/mY5hPywZpwvzinbvsySh1328ZoOMLn3Z2yP46PZCn7O2xl0EdQGCLMmYSPIu
mP5SJghpB0XHwdG0DYiNTGV06LhOsctjPmzXiV3AdHn1gfojAQYbr8oS36DclU2gwpuSIEAOJ8Mc
OPX3bba7svBOIoTZcEZk1EX5tMjiUFc+2rVO5dF594zuNvgueZsQzI6riJT+PV1PAiC7yc4nEiI8
x4aQIWXHR8rERpfke9QdYTZvpMEr/QTQ5E4wd+KeKCjiAvJnH6dUQhexyRCY/+tZTqEcx1GvnAbE
DugQ4KS0HsXFHvwmDR6TFGNNHWyzNuZ4uVlXcCeTwLGbWpzC8nUbx+6kb6n9rzI9fOlkVVgC+HyD
ynhX4dNSoLkwpV0igb7DXRIneI0cX0z6/dXLgQPVzIHPxbfdHMmzJ2ftd2Us7L0eoEHYy6AonqET
/rhQrMsqihFSOmH2F6muepjlL7RSsImyz6oG99H2YXZdsOj2nnlqu/8f6dkdl/td7bX0CckIV+vG
4n+Zmz4LvISAD10d89OsMGlEzuU4Gz/h8KnCQJoUHOXkar02PiD1Ld34QatV6Wy6lFy9j8yqcr1Y
YgN8stMlGYh4ooPvlxyXjJZWu1IbVlYO2vWw2h4DqJKgX4l7Q1NmEDwxkvB8wIxRhV8fKSq6KehD
d1zKqAaifNzjLkWHdrWhE/+46IwIokkejv7rG/EqgEq4DeLyHylU69D344teu6H5Km3jgtinklRj
85ppWYgcvbEshEX4DunXqWNDyocskZtjMS09zhDTpaPf3TCOG4TpAXx2FxfGmYGGy5egCthLa73o
n2dVE45qncquEmhknt2QR8V3VpvDlKN0Tit4SIJaZVH8qdhtGLULiR1ajuWquwa5Ewj6+2wGdRjX
1ZMTBScnVBRCnbURoJ4HMwmNijHmk3fZQoqZl/iSmwE6nBWrB542jji6HgidxAYmuw1RhHw/ayHo
CTtBK1IOn2WWURlJY1GAZEf/Zlztp9mlBv0p3BstwF+cnc+bMKVLU+XRIoEPTUbRPPrCIAw+Al0y
Va33vLTFEiwgvUxBiQhurOI4IS9ah/WO3azyN9OFCZB2d99P3XQk3z4eZva4upQVAm3JXY3H9Ov4
4gY9h9Gj/BT59rA6rrfs5qIwQJo+xAKUVNiQRIqnPaRdItqu/uZ62lyIpjEPlin+21TLCyfbnY+V
z6O8dCCLeIp0GxVzTukbUhDRjiQ0/UZtMFfwiJ6KqyiOCexoD4rVuQ6Bvgpsvu0nJl7HWMHglNLm
f+gZXy6PMqB/WkrD8yxnO6rEDe/VPOLX6W4aOfBbwLoSFSvzfg3LW6crdgnuz/l4IU4SM0pVpNIu
N3+hnQxWm11ianoY9/gVeH78JSKdQFa2q91uuguuffCCrctt3ft23jIkLO+Ws24l0NGXEHZ2kHK2
6uuLVFc6IMZZHC3osw1tqCYPVkdbVi4o1oD2n/UntBYmA/lM4665+tuI1ec94knTQ0bsihsIofaO
klPdKwuxQUac28td7ul27MSD/IevC8hbu77i68JoNnNGojwNRnjRm2Nsb7vtKlmfvt5hp7BjD7qz
fu0vUbv71sB3/aAB4FikpLBKavZ7NzvzPeVZd5VxphHAGtmmdv2aIKkKBVdG5e2HoyrbnEqIo4TV
WE0DJR2Y7D7/j0w+YWigR8CnJVuAaLCmpXjkhKqN5Bn6vonGfKPksyGSIZn4UzTp8NJBcFdmx4bL
5oHpKAyxp/R3Y0hC44aDzR9Yia7/O2Vp70smBtLKx6dA+1fptBAxCzC5Kox3EzarGqZCj6vTAeww
Y4TkrD+RljzI5kwxZ6rZqPExnO/sRySagksXMeN+2VNtoUaKyBLIf1OYlJ4JdZtEw7X+SfV2hacT
w/glVxXqxjmPmq8gmw6SqWl9vRWiiYd1tmg1tZaq9SaBi1MXyEWeb68aFXxUGxllcsCArZMkzFCf
ehIaamU5kH8yMkrXGvQ/5/zxsbGgP8R/w9Sm67UiNVlFNXpiDjEtrcNIkMo0FEI+WKsEcfkbY4Ar
Vh61dmuNP5JBfYRWyaK1j3KHBRElJVN6uZ8G/Q3arN+L2qmLpW5B4HXKJTUGgpywIg5kDcC84UlT
E2kgMydLeLiGzPkF3jJKO90s59ahkShoiMf/WVe/btmzBlS3MwHdAs6/WdfYFjMqEpJ8ocALc+Fq
x/cLHznD1d9AkswaBe5PMtwMDXJEx9iZc8+s1KSm27YL4/aJLtOlb47R+QwXF4fME+U7g6HP4utr
ZJFg20Oiuq7lW1mQreDO3WMSh4Ip6kQpy1U9I3f0bj88m23eEiRBDXKPLTPF4hVlqptS3nFQAH44
13VkOCrt5hb/ofojsyxlQ33v/XwvAtIkofkWCOWbGNHpvghvznGbe0UM9OLOBob5t/9DzRuK7QhF
i9ATxuBGFUa12A69Qfg/ChG5S1Jp7yRXdiXVUQQS45HsNn480I1KoiHt8bCK5/IjtblJbZ8ZX6EV
NsSymgWr6x46W2NVgcBW+vorH5bvemFDr2ZhRxjsLyaER401oNvk4L15iFj4p0F5hv05qb1u+JP+
MEaF3yc2JTzHlNtmGRXO3q5j9hvvvgOTDnHkwa4j1P2KnfF2mk7xxtMfR/D+z0n5KilNP0Ewoeoe
A+JO6NacNheNvhlYSjtfDhg5ldw7VXO3f04DITzdh0bspQPCXYoTDJlaQSOZNBbhWKUcYYldfeu7
HLO1OXOtvH5OKQClbTsCGSl75QsWjgAac4uY/u+SUDz3ZwIVP853mYA2SUbkm79rF29dPapR+pkx
B5ura2O3ZVXd18MjNpom7YEFVO68pLpyYhXTzJ/HnyXFt028BtqY0z20zpd5291mA2vwWx2dBRCu
9IsHNSl1EE1PxQ97nljK62sLM6wdOoVa/LNL/uUtWw6iZ2tRyXlShGXSN+/3sfTkfRh+Uzu+9lqu
X7b1kskZYlvCQ2OhAHlcfr10Dmc8nnswtuioTv05ywKK49BLJlW6H6/3vHwkHyGWLHUBxh7DBfsZ
DfE+lLUOW+4o3304soDpHF6J7MwM9Wm43ujY6bqM4ZijL25IDJ1sLhMJP+ChPBFuVqhU84j75YhJ
FG3vOruWSXEUdk5ZjEZqDyPXrD3dqNGyYcDxD6gcybm4iwXeDrHl4finSWOTNzIFZ4qikPpgHNha
bOhcMdd1VWmstSsY9O8saktnh4fjwRqXXmWw2SIHCdpCwBHeftCd5B12WoqKd4x92olp8lwc0bOs
xC9X2Xiczm/9cXvz4CryI87NOJjNES6glLspiRz6S31mXtMBIrEcz5r/yyGQBkDRvj09LhYkr40I
bl75Q5ctLitngPU29F4zzAxMd/dbGRTzCbCYk7lQb9Tw0Dgtdf7GQxFUJnP5jlxE7kG9Lyh1xGf5
DrsqGjiM4L/rD2oMQ9sUFV2gImWTN+/YqQyjIhgqEIbWiUbdQcxLarFzdfzBR8hvUGrVREmVlQ4u
F/cPC0k7iLraz9wcw3JC6hCTzCGqUGhMtoD59l7u+zc2f2KnB38HZZRnViMt/bCCuyYP4gNXK75I
KOGx5dEYuthapTloZ4Vruhu2PzAbarPQMzdANqZcvyXkEkOczeem8vPpXisMoBbbC6uc1jeqYlDk
uNDiRPmUuGfQ3VQNT9T46uFAGP2z+XAgyPxeBFbK0M28SMNcxZTAm82eatSUEDkuheiBPtBbugXB
2FAP9VCVkGjR9vKLHG+7yjFLdaow93YTJELNmAs8mdnuXZo9LTPat/RgUPurxn++p7fJ+Uf3zM8e
6Nj8duvl3+GIxj9wdQw9HazlrG42V/Lhps1IpgO+y4riyIp4LZyIF4PwZicKaN7sUWhhtBhGqrEh
EVOCVLFpn6y+7GpWQbIzp4JiibP9bKXHZK3Z6/r5yet3kjqt2lRMstfKMq4MASpWBpFTbDTJrmwP
3/BCoXp7vzYqLBBym3UwktjtZBR4mFa5nJ93ZhczyfY90VY6terWaVoJwZVqE2b5Q2uXgv0lmZ8k
ZwT7Qy2y6lG6sKqXiqyqYQqjXjVPKYDva8xD5b1b97qXk8M+EO8tONOpyW4UC7Tvb0HY5bK/OipP
kAOemngS8tLHwPly9yi1lEFJX/TaouDIsaYXvPL6QRPtZitZ/8dJ7CVtJyJqYaXPHUFx5WadJYRc
N1qib2x4murUH35sXeyPWU3e+UllbLneNo6axYNKlBoOtgQXevxgR84acRRYX3jFo8cPa0UW/qek
PE7tgev4dyQZDU2r5VgxImpKIvh4b1YHshHmvhcZwJj6wdO+ubE8xGomGK1xbY1cnGEfrVlfS6WI
IXk8J8uRf/oX6Zs68d41WTGR757iDFmIZrtSvq0dPTUKiy1UTJS/x2JdhEG0DuBa5bcjP5wxkQq0
9l/5hEo35aFf/tH4NxKeM88o/h5fvaQpoFhPEakipHLF5E6uX9PlN5ZTMEqLBHEhsame8ii7SulY
gxrCgytNskzr8u9h0z7DzxGpcrNAsx4VPAhF2s6ifVE72+nH5NAE/7ur+n0ZICtAPDGkq5mN/ERe
cj7jKlF6PvjFhyY2lHbOie67BiSLClNMjF7GS1tk6JY9xoKKPeXofkcA4Y/NGiDnSSAU2K9es27j
TqsC+9a/iPpUI11IRkBEawDi07iL3AR2q7WnBRXH/qdkpP7C6OVzQ3XX1kd1uX8PYGKtacV3Ckvf
LllEhULNjM7SNikAJ2ul6N1Z5afGVIL5YKrJiZpsnwDAmxomQvo6Q9xGtq7ibIRra0m/VTLbxTvD
PFGrPITJKD2c5XiKFLpPJtZXCW19pjVKGao2D0X+xyzeXntPaRXDd/GrEpapsjUriwP3emOkam83
kMZYJgjocSrK3l/bTyzdNw5P345AiQTmW/RMuP3wWJ6SfO6BbWpNVrxe467ALuRrSTUiyiGnKqQ9
UAxih1S8G9mgKtc1uagRI92WMkl8h7Y1MM/BxINsYNJYccUSZlrI7K/Nd4s1Amfmk4ORVU8uu5r+
VMPj/ZkPqEWzbnrj5mYWlrgZkhNyKPjU/IOY0S2IJ/q/jR8FEhQqTWacostp4d6DQNw4sIP1VO76
JNDU/yQRtaFBdNgonbVKd8+A49UcYIEuVWjbtv+l/pyswntVpdTp04rsicc/jWxT0T5j7Mt+Nbmx
a7vI82oCarteubztjXa5pOXhNS4bnvAEt58JF7UooAJyOtUMkowlbKyMdfK2rqN/sn2AGo+wBs/o
pp4+kvTsNVffwP1FSSDqo5+u1I8AG0+IQC0BGW1VT+vNjn3iCXCHlKg8UYgRGaulFXqiZEytwQXf
XXYq97B1zC2XnDcIeApK75JHGMR5b1S41x0+Ge7vlG0rmxXelEXNafgKx70xT4kz4LWvvMCi/iWs
+BFzTQJDt1pFPX/GQPCP7BaqCFBYLfNTQYaykJQgl7qhcAutD0MXXhxHwijdmmDNTg0dMADwFoPG
c5mRVXQ8GyJvkc4SQuNlwNJdBNtErZcFszacEt9Q+MmyPtm3R8qVhB+x2Y9Pdwk8HbuKTw4RUacw
Ljia2sSCuCkv2iA7Re2WspoEFlj/oOhNGori55IFyhv4UvdYZr4tcZGLIgnNVcj+WUMDbmo+3iha
mhQjvixJimqyNNPFPRA+NRPzfYwrSuFqV35oxAv057e4OP9kJ9awhfsPmqQVirQeWEtxD0DdJrTG
tA6QTHrDbgx0llb5EuZRlGr0Ajj+Qo7ro6QqhylrLWGQ2zJxhVQfxjdv1piwKW1GVPzgoZui75su
eoXBLYSWrpHhYnPrJPTFzXBJ/72esAkuVG6e0a2kTFR2pXEh95CrQAKsp04uM0RvBwk6D9XklVjM
T4Hk3zZVBnjYYkdyN4lDDQ2fBuhcJ1piy8Dyn2tJlTl8ahuh5u62Tpmtg7RGmx8s7O2q2wor/uqC
06376LqM4bhk56CjCHXjbhNG5W9gIxr1oGmv8duULpONZsqHoD+WP7bpzc9hWFz3sPgksSuUhhVZ
Q3ZdPUtsOVpGKtogR2Ea9h+U+1v/MpHg1Q39TzxCTU8MfxwB7V5BXqHDl5Lbx2PuNW8MFfy7h7rt
164e5d+bVnmhHTtLIASjgOwouB8tlAAkww1x6y/lcUuIEkaPDzfWP9tjDrrpu+MBfu/j65KNY/ag
naELwPwA0sy1Bh874yZ1EocaxJoLVvi79Nr6vIZGgssNF/huQs7m8nshb3cdWzloinEJZtJiVNwp
TvatL9WGbwlhz4bEMvjQs4q+d4VHfOrgkF2EJH65swjxrPB+Pt7EzS5nd3Eo5mbiRCCVnHlYnpR2
ABNALot3Mch45Shb8GLLSPlYPlPXXSROX3VuBIbixJoSXhATbWFyy3LZlQHzbFT2MosKwqBqwMFf
0cQLcRcDD7rA2lav0WKmoMs9jeCD/FTkjZLQpglbZmgP3TxIIFHn8r1hd6/TtCi+DjOWvXP8IUIC
pcgyrBtTyELHNeNpqAKU3mkL83jv7Mc44Btg6k3L4UR1VHpo2Sx9t8mvFpsQoVYfee9GzaSdzFOc
U3fLjUdWqNXYm7A620n/6pl/zriCS2AJMmk1mgRb6uYck3/v3x/xYgbKd/DomJwURsjJgwpNTqg0
CfwDtT53N1Bkoyv6vcbq2HBswKNdlF6spBcY6c/SNdznv9Bxm+9YwcelTgzUBUa31tOVPJ6x2vZ7
+fLC4qPYdgZ/7zf5Iz8xlNDpJJj0Ynb+AoOPqdGc19GukRDK6m1g/Pz537H7bZFcYJ/vd0oZ8rh2
iUrgPdQ6YkZ6MIQk5QIEIi8VokQOrmc+cBr1fhRAgljMSRZQ+p4FxDbDrj2n4+o280J+Kr6Mxhla
3pKAtJC4/mGp5oevKHhI/zHW0W4X3l3ZhFb7v1Fvb2dKFdm0FsR0arWj+TSbHXj2uKLQJNaj7TQT
lkMufJM5w6VcR7Js+NXeRSDQ2irk+fsIvQrcWPUibf6hFvqMNME2hlv2MWjBdA76riU3XoythMOv
nePa+LLyEW0bC1QUalsw66NXGUx4Bq2cPtLnsfIhr3VlEbSdxCMNgO3SuXHVC8R1AuDkOIqb+DLd
9sA1zn1RRzPt2Lu9yQkx4Wll5fXh92TPjxbZwPPlQmS9XComW19EfFIdYq+eA91yT+xBAt8Z7jG8
tZsaPTfPLg1CbI1D2SJgH6saj1ycsfbGscUOxHRovyQi7/lPaPkUAjv/uxCCq1XJFQ7rDe3D65N0
dM4a4AINM77V3XeeiPMPH/WzgRZT6WhTokUdIh/RwNr3qefRoa/vDmEoSqW3KrADscs8Yyk9cWf9
OX58NhGNYXiIoBz8CjWM4ro7rTfnlxWljk48p06Lkdv0KOPhgg93y/NithQxk9Mh0pycYsvh+qj5
z2oBdz9dvZXru0ebPnzvdhsW/rYdGtNkMlEJXy9ow6NzsDoxMWGW5t0e15FkIJ90cNduNb5FIjZx
10LbwJjVWLP9kgscwOoED4UYrQy/rS+J6UWjIOgVOw4WdEVKYpGaXGL0fiJDVQ8h2wuHfRi+MsKE
ZK61Vqi9/jSpKTmt60rbxgDybb/6T/rkan7cPlzRDeiGQS2TCDoNxDzrn/qk54YmGUdynsK1POek
vaovIEeuE+9dhzLcsb6GNrvDIiFDNdIJFHUqy4mJSiBV9bCw/viqC8Ow5eqZQXcemm7sGhZyR4YJ
/DNv0Wj8oFWFvdfgNj3FWs08HpdHEJ33kv+GvzSrjrkxixv/itzL9Iz+4235AmdxPCC20Ai8ITxU
Jz1Uazb9/bBGvxXaW+BoTr7PbzvEr3++pIshykMQ+o/XaD0Q6Rg5iiT+kJldtaiLyT/b6EpIK8Ie
WbUsbkwekc1d0UCBm1lZXqJ+AxrZ+YN94kLWohO0Mb1MouZtEzdBlurKVpgeQ7Z7aYxr+dXTa6k/
1GUZ8AksUhJ8bOGuHfXhnfWCaQov8JkrwM75eYB2AVfh5XuOiiD0Pryh05LfxZgl+OHW3t+5j75Z
YNURcI0r1r90mmXBVaAnq56iws6lwb6GDQEfK1vPm7X2seOA8Fu1nBu2KsLe760I2SZCA+81ah/i
UuFpfNKQLbV65IhaeFCe6Ln2K6dCqdNEvImPvoOAoD8t4uZNWlRvxv7qjYjR8D5iu1+DYnTRw8SE
t1Eb+s83B38TtlUxzUDzQDzdspNog5I6nG5l0u4JYEqSncOeu00skokZEbjzjp1HWs5SI7Ls8TDh
PMxn04jYsWh9QEKLJIqzbDSzg6k+/J8uypi2au5/Ru/fCH6eV4F1xAboWYXgLoIe2Fe4ncq9snMu
6jwMP4XafytOPmAzHfdy6+4YnypRpiM4YrZGvspalwcVdm4dnCsoWA518awabCR6nuVwL0pYvS8Z
Hx6yHvcbSVGstsM+njRzrVIeO0ukmCqJi4EOIDAK8rfLWE1hu/r6tO5q4q3EexVj8L/DqvXVspbI
E2aIiD/uLXtMK11OXZySKV6gpTnUITLOADv13djjwDcjbbTwtdkuCfdID2j3cML9hIITbfzBFwMu
1bciG/c7aSorABtOkPQ/6Yus4unYHmEVWv8I051GTb2oKdR6plY1jCy3JhNpvkyfvE3RK9J76euB
dIK7ELQLS9DTo13N7T+JIR2BOl77lmX2VXjuf/yt64depam8TMm3hRVtFwOhiNRvTgVtYxbWIEl+
rhzUYLrT4L/r0k2e9hCDbOWgXTzbxt6uDZXOx9y3jimy/9KRofJqHOBPi12x1Yyb3iW3Bp64AY7u
4fbd/JSoAzJE6W9vYRuEddp/6fW3Py8h8C/YKqbjnk/dC94SoTwYtPDSHB0T0YYbcP8Mu7paEP3B
Jj7dYVu8D2V7zb0cMhtU6EGRqg62Wfg7mE4KK0ypLZL/VTAhJw9Ug6s75Z6Z/tV2IDRAcSjW9BYX
Ri6rhfo43c0C8/qbpk5MQXaUxhm3QjJ8sViDwfEYKBk9uBoPZFy4AfWdBl0o1s4YdJZuFwgYtcov
z9Sm2IZiBwu4lRS/65SsMYHrYLBOi17wQG0nBRY/3+4T/SEDa1fJFl4B6Yt0HeaW8IMOcDKRZyvt
aJMBdexpitvWimBhW5kwIQrd33LLn9D/h0TCu8lZB+YYewAd4PDrEB8Xqu62qi8/SxgrPfeccJ6g
RuDHj/7RpRNxsnEOD8aPZ/PH2xG5k7ZV57MWOmmVayNezNkxSLbTqFtkXbDMdw35LaAAd/XYBMQ7
wcy9x15KnbAfRcMRP/28arDukGsqJhP3uhpIbzo+H+YD5flRnV/zplwtFBbXk3xXF/BrhAqek/WA
AlscGBnQID/v8ETP2ZnciVfbAXTiuX9hYZgjeIIyoA+mBdQpF8fk/AU+hDYozztrDjtNM8eNGSkF
hoQO+lOyRUDZInzuU8+VSNgc66JsY1q/dAvJyMwJGA5QnIZ6EI46dexx2YFxjoP/uJWebs/MGmVi
cjJuLg0xGxQboewcvXWhxVKaLiTZmVaiNuYW5Pck7OM+dm9ynaOAm2uvwLn7Ljuvs2v77NRoFK3n
UBZSb2ZvLWm3+jCQCiywNotgsk0nldIpr/wrxSmGbnz7uAGhA3iB8hD/d4eKKNQ4dIYSonczXnqZ
MtCNICNBIXZ8u2ZyhAia7E9NI5murZtAO3m1LthCSD5e8RW19uclKXfxaHgQsit6LGJd3Wbj5fRG
6lGWxlZmybinXc7EyF2uaUEiP7cwphDdZSfk4fshjuve/yvgdLB6j0eDnkOEmyTtbv0q1+XVLdts
yHDqOeXjH109rki6j46so/Kdsp+cgECtofrj1v9AUOYeA8IZH5l+8xzFaYl4775HLNpQ9ZknOues
k9H4lJ//sYnaVRio9BnnTotFCY4JM1tXg2vicwKFhrKy6cvu79S5sXMAa9bT5mlDRE0tysZUnWqT
Rlvhkj5vN2hHmWVO+bAKn2IWnEZL2bM/7QZ+/eXTXLSQ1gtTfe9Q69IwUdxLJgAXsrevJlVcTafo
KiP6aCvya1kjzcVi0qIC+vhFiR8mhpABE8Kq+aLUPO90l6FL53FpklPm9wlGJ8lC4cuQrmrUQ+9Z
NQn4R1MK/Ve5EwkCFV73gzavOm2V0du87uZz9V46IxaWH1p7PhWofmb4ZSC9fbuCWvenjtLhrESO
LeUqndJ+hUQgiuCvmwQinkl1y4RPaXkbg+Wvs6z96FOiGM0yn0MBlkHzOzpvgoFA1Idxy0wm2hgh
4MFH5XNXdjOIka8nnBpd2WRL9fshCrjav51sNd4XEvmlu7puVRdEsPHLKO00aViJU7hg8/+uSQY8
TMuLxMTJbp2SQ8QH1b3nXihBAevhkilU9SJXw/S6qOnbi2ft1kfF03fiHcL37G6trwh8EYkMgRHT
z6AUcjxJ8YVI9cbG+hacb21wTBP6BkUQcYXG9UH6nL1RBH5MGF8+MfwSbhF4flcW9aMztsIEsGPV
avx87Mb5ogd0Nlr0X6NSfaeWZXfCdAK5RrAGxFwnLUWRDeL6t2jpgtBHy1GB4jF5RzyXnEXpJrGS
gp16oAJ9a5Ufx4toSBy8rO5Lbfb+NUpnvVqvod0X6DQtiv505IPpx+Nd2IYuXfWucY1NSB04v2IE
7JIFmHtFd81la5kmO1oKEph84DHRsLe9hiLOZNjjwJ0tcYCN+0byA3S/AnBKycujAF+6A6lUWfHq
jwo8jlXBF+UpRHJCjpXZiJuJQ0CdCP0qX9J3Dxsea7ngJ7vEuNUNDIBQ0FgLXlUVD1leBzepw/fd
oxbjZUa5rwplO8PbZpOHNRffwHhJiFSopVUmFbPLg12CNkwexf1kN1oxzJnDblb4NL+BWQ4BS921
qMcP3Im/R1qP01JxJY1obKDKPpy+n2qytRIyixyDdoVrNBZ0moZebJqQPebmXilOU/6xAocjzSPi
dYcrs+a6JJG1SqlaNgQ0OMJBQeCbGw3dVdm53XDqji8QufOUPirxHfXiMYEbHBrgoTtFhKpAXPA+
wby9MnvpBSSfJj5nVAyHWCWAHXoH+qi93/ZWohVEqBjiuNKpn4Atr6bqbr1iIwexgPQU9RK2lD7y
aHDyrb3N7g4w+N1ggBhmQujfZQ44Os/QZhNeJYSL4sHIx4o0UE6IAsYNjNAW9gXU0Qr6+2JGHN2e
aMVtKXyXU5DwIn2Ca6kNaCVRqm085LjTQfDZEQA6k1bPkpHZvxJxAZ5l46T9PJzqsnSs4lapptwq
bcHzJyvi4EICWe7hKyikrIeV6Nym8pIXT9UW0Qnv8CoqTduEPu4h3Hyz5D/XoSWZcslZGz9Oq8rM
2aUVvVEaB8zeaaeFy+90g/CZkY2rxkv4cZzgYC5t7GRwJWRoYWnjdCRCF1UmBcZWxyk7Yl8blHt1
uHnN0e3OQ4H4GtJZx6/05CHsbSqnvGJUg2k1+0fRiKvkoFOrPwevyhwOowhqvlJ7hK2mGzbrydsW
C6jyi4hqYHyEe6rGzirivhBNV9fpxbtz+Gt1pxfZoWRVB/ZlDXUID3GIBl2HmEnD3TzccLeRVEDt
p45BonfLw3yxEsNHPhQqH2+B804TDqNvygABkmGrlxaEUytYlvCHcsb6PZATWGXCcLQMU/9W++MQ
dVmHRQAkWza1kXYM8/2h4U9zMweYRJ9yoEwD6DL7LcSuSszvkjSb0RNWj3GYbSn6lHCZpLC/L8wW
8SXii6plEsl/fqd+99dtNUQG10lttFis3IkYSIssiU8N2w6hxNZTy92G7i8ThTAJKvE06C7VcyTZ
2fVEYurhXB8cbggqLE/3ptHglA0ic8phKEoQrJTyP5ioAQdPDua1YRro2iQeERqS3rQcBUZ9zUEQ
CGF9HMJrUaQE0WjlvOEMA/HC4wR3FxS8NPMlQo5Vjj7U30ujPeoLBO9kqUePs3wWOAjRbapnGmN5
n8BsTduZwn9SPbsDku2SOMxNMit2OhIlpHpiaeIFt+LVioosLD1fvwOM2NPKAuao49UOqEZBs3tv
7JC3oaKTQKf2qz9z5m25RQ1g6l/U/z08B8RbW2qHHk5EzVf6qvGHJjNVz/wvOmgTX/gvSE2/3Za+
1YKzULLGhPWVy6EG9Mzi4L2jKs0kWMij4wMcd15zK6IWtFuTRksLjiftBVetB8flWXUGi8QKAUnH
e4Zg1V+Vg2AqM5RgRQNKLpiKzLa//WN7Eo0YhtKB9dTaIdW5zMKRnt4csOef8Wsv5tYjngGx67tm
oh592AfHx5mFpJXaXgCS3eespv3qfRwmrPVK1/PtFcpj/JQOIUP2Zso/daKt1h79RHmRRBzeuB8U
ZIrJeWgwzRlaZhrWhdGgoqRopKSapHKvTeLYkenGpiVa3WiH130R2YrXcUeuENgO5fe/cAU+3ITu
qNEd+kyuqYlnzj2GS2EpAZFOnCTafKWz+1lORvgcscn7hZtfQxSZeu38UHifp2xCkYwHFdBs9h5H
NYKkl7DjvM5FzKYrtbRCFWnowtar9O8/4OhVli8goYQAXkESVMVu8RhrKGd6MEavNWpXZfEaQpJ8
R/ut2lBDFksyONCPjXYENLbbbHEJjINAOKCtZZVdJ72MEuD5AnX2uu9JAQQgqPZuOJgnFEqsCcCi
3Hbfm6MF7HxzMcrVFfx2fNpztq1x3W8J0IpIpvqXSIzm6qeeHTRVxi6wmB0TOGXyFZ/eB5+oiBau
N0F2Z40DbJ/zcH7JQduWNbQSZjYAEJnvHkrokOYPxPqn6vbRvnVIZPYOpH7eE+fQo9K7vxNvzji4
BLgP7eUDvC7w/4+BdDD8ggA+1kIQRG0ZuOyxDNhJQpCYse8EoBFdSvDFe/2yTIdgcAMDkgVVc1gy
g4EpfbqUGpTro5fttphYEmP23v7UGis45jUuiEl+rYpHkY4qxZF9l+ysTQi0L7MzlzzD4/V2pg94
Z2CeUZiq7jZguNp8JSr9VG6RieXQ/ugIrMjFUQoaJfU97Vl8ae0sS7Hm2BOiuTfSDLZMpuJMBGIZ
yBvWGfMBbJK4U7m9CaKqUHPGWzq85XDzMEFUob3qdrj3pfQZ2UQVDuk2ATFOzGk59Q3Pold+UW2c
0bzgzIq7yVYjS6hVzCDywQsT3bvpHBkRYgmbnf9wMWVEXZZJnhspLqScKhE8YJ9cBrMPrzBYNWx3
DHgTX998wLNRj0U88bqtmaJWFMKibo8DwzYaKQHYakj1ubz75xfUvppsgbkRajrrz0MF4CINkJII
ck9eTKZLWBEjq4wR8/eIOX9ZrWGekDcljatfnOZa1Vgv9AlK8I3epgn315jlEkSrSY893ZPExljS
e/QFXlgSLacx8ojwcnFZ9eB0mVEPFpkRjaWohOTgZmSpMVWSoqXo5//7obkiCKjlm6Pl6uQOcjaC
6P9BT9zm0QJ6FszEVieiExFWhiRnM/AvENXiZ2sfEnFt0gKea/68sNTG544Dl+rJlhfc4VfmWPKX
qCnm9YC+icr1IQuqT1uysqOZkGfHbr+DxKFIumuYEst+cEV2nRVDG7OgG41IlaH1od1ZChrMRR/v
07j0tbqIYZxAa3VY7RbT486HpZUaWLejovYr4x6EYZbIPlE074CT6BygYoqiDjcCyglApFqU4sfr
Fu/zoSzCwHAzugZvRZeV1prF1J3IjMzMlp9PL6gbrJLyPr+S9XYGYRPEx52cVWZbd54PekhM/+fh
rRgq+EuYPm+8sNEUBimHIwIX8HBH2d50dGNLqVYei8Is5y1mZKT6Nr39yKhQOok234Uyxy8R+2Hj
uCXcR+YgsAscJvw14yHd1l9yOJikc8wgyB6ljkEmu1hOFmb5PveTQ3RxpHzVLUAOpaHrIB8VKs4P
1PxISzyMLKfG1jQQtmSkE25E6uZrD/mhW0KQv8CO8D9LUWZktPJtgS6HPMO/t35swK3a+IXToLuh
FRaIxNm6OjcqMGQ06+IEUU/5Kt/jXSjVjccmO1Xf25q3Bpmya640Mw6DNp0HStywl3gaj2eCATq0
2IJnl3nQ7cyD7BkYop9CK0Lx4Knp/x4IYAPGAGzQL7Vj+RYrjN1NSRAFZykozYksZe7LCXGLj197
JbQEMsq+pWRLE9wWyatiTFbHf4gkF56hHmtLFrs2cAMypTbIrosvU86NugxZuskSsSVKxFlpsVXI
LKmKjwAjZHxXCx+stJVPxnGmt0B6ZSwKqv0r3AZs86YS721LoMxAHlRfGRN/Uooc0xWN71MMt7rx
ligKrBdpn2G1qUqNGlqigPBC02TaeMtTuGfkBGSYteKeq2LWtxanFGj5kRYLALaTBcKyKAP2AoWQ
4jeM+9OwUiTKHvVx1NOhCv99EPd5WcUaCdO9YMz/3+2vEMfZMRhT/dUOualLEh8YMCVKDdllFzwj
srHjRC0x4qZwxCxTTCOjrNRgrDDucnbkpSH1chCqSUVK5HWxtdCzA3AYfS4NdslPbsgOM7ddSnEy
WfyAQphVbbYFRBwJUUhrLA+bWENd05sFz/XbbXn83myP5XcVsdP2s9lpcNP8Rj892t9JH/gGM4h/
i+td6eizXjHBJB0nLnqQJwbFFHcxscnJq0wvdJpYxrW+VcOrhR6FlYTih140jGU/Hz6Wff+Cw6sx
J2+qNYZtSQSQcD3PUad7r0ETQSBXcxRsVcNC9BCyQCgI28lks5ii9quPIv0soK93xJB1cSeB3vOb
oWIM/8zu01kY0eXJZIL/CAWARRFjjzaE+F+uBi6HIqvh0yed4YRw2A+IUMSoflkDd909Roy92KUM
7AXhPQ9cYijjkpwGnZoKAeecadFHTDKu/sWIFy4k0UppjTFML3yEeSEIog51g3L90G6NEXibXSPu
X9UVv5LadNwOYgjgXNhlyYZQSvdfeJrUwYxbux2JOx+gYW4uQbYnGAZSdImmXQNe22EQN+M1Ejpg
fcHY3zja3ip1oHfwRqoI+52jZhhIfgC7OZf9/D6mAZEmw7N1RdKV8P8BPa62AYLHIDGz9vo95ZE9
FpBPca7rsEY05IV6mDYEubMibEprIu52+03zzH1/Fycf/tURjF01D6QrWCGjPYjhMOOY1H1oqi7q
lz6inmncuuWB0JQ275aHtRYd20chFBBX7ekA6uzj7IFRT8UwXkSqf+0ZmZO+hzqI02d6MjW86UsY
nfm7Ly1DYGa0U0o4ILbORJCduJpyEUgspxONoYiuW6/bP364GZdPH6icKZINpbbKr/2BTNkee6Wh
MFe34025Djtdz+4bdpcxaoj0CZkg9bzd6hlpPBDyUFWRquExjr22o+Y5rJf1af4DVqNAKACw8Ulj
VPIHDf53MnuazVrE+RNuEhW3rgy3GUqUINNfgCcdCwXC4BAZ19/Ks7RUZMHECgHe9qCUNbA6sF8L
WF8MNEBnlK7C0kaIZUoR/CtWyJSGat8wHVZYWcjfOI7PjUZUyNkYKt6pQg//dmOl0eMC5+Bq6XyC
ViCmF0TfFrLoRLOjIhs2twD0UdlgBWn0t/S8i5Grp1GN4xPrwV8yFUfTOwFqryhzVTSj9S6HxEz6
Eun49HF0YUImLDvjiRm0FEZmG8TEg8GJeRSIFPc44bsV8vkM8xLiMXUvI/o7il3lfAirxbNepdKf
h0IJc15SZM1matysoIdcTXUWGd0WjrHE/qvaBWhRZymyJMcInzs/DdRafZhNvPJLCeefS9Jy43Gj
0kRKHL++7/XvCgzzCSEoPv3kzqWUNEI+wrGrOt6eTENKljDgjwAfyjM+l+XxChlcpnzzds69c1gt
g67Jg2lX/fLhGcVprFWofm9xCI6pqrcBHTGIhk9lcKO6ORUwCg2RYnSm0pEcdlhcHxJSg26zf7wV
tRtV/BlewcXOu1Ogf1v6d0tQR8V+VoWOH2Q44ZmWGfsiuxGaDokeM+WWmWYeVdCtxAiQTrUQRwnb
HScf1X/GkzTF6gEl/I5GCCYBN7aTZD2Z577/SXcRo1atG+GYOVIhDJhqgJqAJN05ERwSAEJTxcjc
AiFViQz4ngOVfCJnc0iSqjC0SpH4K2T1AkbljZwHfmNhs2D4w0HFz0tOKUKqLeNyEJZttKIdiIww
muyA0Dsy139sVRMzSzt6/BO5SvEMRRQSCa83avgm00CC2S5s5aliueNvg+HqaJalIk+waWD/BNGk
px7TWs4+K4+b9arpzrxmfTfae3l3Dgbd07GnplDIn9b4190g51oAGjuLi+AmWjmmvbbIDOgBP8Lm
l+VluKN4UkerSkfFsdMG//VkdBqlwOpn5F8PCEb8Bn4RNGIHBKI/roixihV80Nyri1rdtzyllCJI
d/mcsM0UqTfkDYNTTLIbzZ8F1lvpAGhHzCWoXrrYRDZOVSK8XXlYgpN2JNH+3eVBgFMDUQIYn5xE
/B6/J0C78axv4x/8EsZNX2kjmvwa3T9wRZmyQch3zWuLic1el3Utdjn6EiMxHjv3qZmfvXpjRDmg
uyIFrFo3L9jULAI3qtt7D6zO82XBq6lzlihMKA25kLMCTzZ+JRsvJRIS7uT0WC8jinpUcyJZLeyB
t1s1PipiS24znp3owIPUr08D26EIJBBFIkw8jdHyAld4FNIDm5Aqafu51lUPqF02oIPbWMpwVKpi
ORQ3GtzRhcP4TMz4XJfkIUQoGxbXf0I0oe9iS85AG81X0QkgAkIh8w5i5rB+nEy0uN1y+cLfAl3A
Vxg3ic0LurY3M27AObpjsBK9+IKkUepR0XCph2gn5NGm49ZCOsK/fIh6TC1eYVhHZ5qJ/lIIvqRR
fN1LuS0FEBLvbHPUIfdNZvjbm5N+2Ct33aS9JqflENwRo4chqqoK7VU96HHk8/Ccxz9Qsl/A7+wm
caVsYvgPHR0FS47aSxYtcKkKeYrJZUB3S4K/7MNbPkICKaLjPwPHoJeWbitLs88Guh28+7q7cL1g
J8zjN0LzqkNSGLd0zFRtMiBAPNJuiaEv8L2pdrSGASdvjRJBwBK+RlLDImyI+upQU/3Sbo0SnIXn
lJLOb5a/DaBE0omvfzpVowspEb3fJPK2sNvFiI1RONECEWHXzac4UZc+WI8TM+Tb7mKZFJ6D7V79
O308Bu0O5amUIUt3LbUsnQKZ/bLZsJWD6BHkI8Rm8SXvE+fTcOmpp/Kl//7WsI+pkZYRlcTNNbrX
nlxst//w4lanCcJigFIu2S25bolJHaGv5jHbtKKxtnJ0Dyh1dOu6K1iBldpHLijwfgIP9wkJw/5g
ZpHspAwl2GVy/hg88VJyQaZdeX2tQfIZzvourkH0vjd/aenzc9OAJb2nFxWIiqTTkHMRxPxzljJF
t4JEb5A6PyQIQa6XX6bH0wuiYiPRFZ9wE4BorjD5if55RlzHVIWlNnbmWa5F2JS2IEabwzB9/NNy
uHTFuTqX9/KIX3vS1ppzyWPFuNWqvcwBD1EZlz753yY85optErB4DR1l8An3zQLZTTEw+gTUs53i
ES2pP2l4HRL6Jn3fbGX4ydROCKSOoXE0Oyb/NVorGGDZf5zW2V0TSKgeMJQziuJmflp8AFo8Vz7C
rfrZHOrEVp3BZ7Tq+B1az0UyPSYwRAKulifUMeiYcbb+Ou6Hs1nlNb/iVwpLXhZd5Pmvwm4yBp3O
q9buXQoP3Vv9mZl1h3YsYarKDGhLG3e9DZ0uyBM/O2+mrAuydptf+3ViPO0kfOXTER2PI+/fSAxA
BYquQ5F0P1b9sHjjpVcjAV8GNs3qmGwFUIFAbvKUhkinoV8b7qYrccvV3VvkkQ7dfnzFy4gB2EC7
WX7RtDG8FKgZxAzBCRvORTJ+KWZ2L/C38pMwEgBn+1JS9Kp68F/YON6AHcR4a1yIyfJA4w7M0CmN
sv+in27WGlB+I7MFI1Ft56bvA5zv3w6MVecnzlv87SWrz3UVbc/K4ehjR0o7yWHXRy+lyi+RbbO7
g0Ytta+EvtdMxLHHsb1W3wp2/AKdDjzAiM/cvuPlR4EK8dvWLmOKktlyev99xIQEv9WVDO7omcW8
cWGAsAujuGIVNHI5BQNnPicXtsMaBiakOsbCdCziWLMmsqlT8gw1coKynw9bSrgXVqYXzxJVbrnV
uEdbbfranNRgwIkMaz4CPE38IeTuqiXo6qlidhiobk1epZO25OzIf4xO7GNVU0shn8CURHz/Nhby
9LsfWpcioq8CcsVIWPz7IfY6BGvHxa/xyJujEOthbkTBFeXn++AqU3mGfl9VDGvVPIYdbs6JeyCR
HDMT8YbrdJYziHxjhEcHMt6d9xT87ykaU4OvaoP8PBEtT7DBtL11vr9AeCCfAXBqocrtRARXnwgR
P6OU6WxE7aU0PUwN2m7yWCkyk15+BtxsQv4KZD2R3L0kF0SyX6tx+JqhYiCGpc0ro3MVPdd4W+9Y
Xwh+ik0UEUEU5WbsWYbOHTBc3MlnIsd+sYS763mFuEbAN7tZkQt9AnHWxyX9HBHztgQZFw4Zx1GA
B1DY0uGhcn3NEXBGNUiiEO3ZMmWXMnTEb0A5sGSDSl8fmkWJTqzTPXb87wK0lPtoQZ5l60Fg0xv1
1iJ1h4ghEgfsyZEU0373zokFW0LxW83qu8y4fsiyBjFqxpTawRJrGQEmXSGL5XJ5/IwuZKvqupnx
kVfqMNCdtVajus+PYJ2uh9QRnZoWYy7ZvT/cfWXoTtUYpiVYzleKef90zotx/7X/eYjLRc+YuPP9
vFLykNa6etpXu2E9Zf/xv6LUifCHljVjuE5Aw4lTfaWrpYhPOEKQM4bO0Y+FmANtXFU+Hmm/9XI1
tJaEkqva3ASv38bi1wEpY7KesAINq5F6PFa4dd1yczh0tyZ3654xbiAxBbWR02RJ1KXxQ+E4TYgP
uIanZxFbUOyW2f1VviCnTNwBsouC0yf624vZgB/WWlRk4uHkuac/eVnLliXrq1+GpxN07BqbMokt
haJZGLN685ayyYlE7S4Wru4AejsoSO6Bmf3N3KbR8Vx3csNBRyk+adxVh68GkgdVYoY4o0/7jGau
+ymIxAZNMrGjeRYC7WHYH+ZtAR5go4eaLHXlnGsr1xMXT17mC7lYNBdRHFJzq+GuJjtVBt/L8nxc
UYYXkiQlVtJcCg/MOg3jCwWitHivtcMj8H22Ire9ta4+kf1c2Xc7WnsZrw4V35HeGvfFTdHombse
+RcER1fnRyBAtLoanHlYhwnQBSavfHAML4+HIrdEggVBoNRdCLwcO1XEoPERCAz7+yajXsycbULF
Zh0RE7zM4MOnPH2xt8m+4ce9Wi8UQ56jqRwiyQc7yNbi/f/EY3/WTECsXvwAPpRteWWvBqexjMDt
/P6rGwSnnPF/r8Wl+iSXlWH3mrD5K12PQwchC6cPYJlOMeyin/zDraKBOcpv8d2UpsCqZOycoK8z
6daTQ9rm4Ym0RVBa1gXieZseREZFW8jKjV9ucwI4CpvhcZyb6YmDoN7RYoOWWnP9AEue+X2UPLDT
mk7Zww3OelBHuPMcnuvegz+EdFlUGCFtxVb7jgQFYksmMP6fof917GYMDAFW082VuaZ42fTO/xxs
Tz2ySyLny55IhKDXopQKjYR+qzBU+T1JtlnOAb+VyHQg1I2CH9By+BOSfC2VZndTTFbFJYtFEv59
jt98NU5x4uLIIffzS4hkDZYhG2vXgIaefGIEu0CgIfn3W1cLE3CrRGj9nCbN6eiE0tJvxOgr2rKD
+8QZh8TWB9xVDecXXbAZqO3YiyGCkHM8Vobq2QEXUypl8nCFUL2tNx6kzS+8tGo6tPxDvugupokb
pS+1hvEDS5F5VZwcPCawjZaZZvliYS8ycZLjAkhikrUGILkcVsVtPGMPao1x++wuMXjSgkkX3+gE
l3X0193Z7N7ENxOK+5DM6p/i80JsEpcRn+ZjnNgmNBEsicMEjXVoPkO1hR3H9zRBya08pkROy7sR
XRbHr0ROuVuFiSn38Km/u2Tb/UbfW+iyD/02Sq5cyWtbp34AT8vhYzuXOrPI1PZ6PChaotD40HON
egXQJOG1WnKSN5vTkk6/rRvkAaC42ypyjCGlMYDS9Ygrv05J+f9waHQv/t8HyQNGETecLXOMAicO
bND4t1kCNalTp3AD5iN6B0wAJObKnOBM5UGp3wJi4knxfgxX1kndgGzEfgflsc/1BZCu8twYIVdn
qNDLN5svJiIRRuGfyqonR0fWjQn+OsTsBg9BIk1DnMAA89wx4usjo1ay6PmiuTLA5jkTgoTVgHqs
85OVd1+f4jxNY5ECdf2vOkES1oczLzSHDa4VVA6m3/Qm3DIJrzT3QLK/cnF5HAfBugfHu2qxs4XI
ZwtZp2rxZtOA2G8KXGIlqBEL6dmsbA1r2Z/j8W9OJIJkvQ+em4124fKJsqF4uJgNZiODZAYr5F4P
T68iWYMRC6Jm5SlFTHazA/ushJ/v5dz+NujoJsKvwBOOiPtXlcd0QSDjnAOqpozZYc+GtC1rVk0n
kO3QzcHrHY2RLp7kvGj9/xGbQLdhhZ9P4EPb/RQ2dyqy4D/mpp415bZ0Y7AqzTRbgIvKdOGTg2UI
8TfwkmlLtnO6cksNdZmUHv03uJoyn6zGu3Ziz1gkDDa4z5/9ELGSVrQ/lGXtCyr1gGGe377tx6EV
6G58BcpdueZkC1FDehCxcIbDYt+7az4ca91RWz7QrqEawanpgatsQDPXwbF5EoomHgpMQomYe1MZ
STrKNl0oWUZp9LJ7z74YX0zdeUB/9FtKQ9NYjuozlRZhRDE9shWQ3KD2VmIBhJtxy4qmyqnGSiRH
vSMy99ZP8fCDIiLkBklSGKMy+oHTnCVlR6IvidviiAzQaC+hqpc7oCyiB/4QgK8azNQbBns3e4+r
n23XOgUVzoX1UcosFTKu8dw4/bGxpLiNnjJj7wZTFQ9VT1WGeZlZupmwdf6IehCADamktuHYyJHt
OYbZkWH7i1F2eC0kkqfIi7edWFezQaA92DcmMuUF7FGMQanDpoQQiS5xvljVgU8bdirjU5byj84K
dH1D/EemMfPtKVSKlbqmScLjPbVTVp/m4Gx3wuHyT+OZJJTGEONl2fTQHB2wbMww4wWTh+vCFW7M
SyLOT9YyYK6Ao0sI9qj1yw2tvoeefYyO12mwxVIP1SS5n+SVKLGGgiq2ujMFILGBIrD9Ha/h9748
IPD8z9M4gKcbDdZgDPEC+g46ZgSX6tsQ/B0/ityq2wr7oAQAVfDkn+jhiugbpgXtgLL+ZAS3FPIE
2VxYq0DFRhJmK9JlJTIXRMqYjlRI1OlH0q8F9y7oV4F3KxnKDeFHcQSWnMe2LVQAUehRPd8RJ6ij
Ymvp1MTmAm/pDjcIy0/+B7xsXBTPfqy6Wzu41v9uIIlRBS0I6bUNQpILoGHyiZoe4ZyU/oqqUCaL
HYmvOsNNvH2HuAx2qQc+F5Gju9Wx2oXDgta/Vqg4dpVhmHR7S8n/BZLYWHVoG19enE6mZFcDqTe9
wkzLL5Uf/vMBDpMYU0cEkvVsxKZI9wH/9n/Ci3aB6O4PFg8qRZTpl/BpEoD7HHHUj3C1bV8CGdM9
kiew8Zs7ggvc7JkGoZ3MRwwgbrLroosaWqQS4qy4pPJ3kRNY28DeiNrlf1fIy6Vz7OtybPKBujC9
N+PCGQZYy57wTTlOF1hy7uWibB4w2eMKjXYnG4yvwZak4pr0fUVn2nDvT5LNF2G4nUxDEzJ3ZE/v
a0Yn8mru4us4Kvn+hIR4gVOFY0ru8zy/tPusNXiUZCW9N65JiT7jZkSD9F6avflLWX1dmfA+0pMe
Noj4P4Nc4DZ33i55RKVe2eg2wfz6+mLGJYYdFKeFg1dxVxNtES5e7yNyLamN+p0lLxMy1nP+SWC7
v1lfFR/p+3eD9xwwKCYu88PrkC8iRnfkvpqZBSpZr/MURyPtobdyDGS9sW5xx++H0xPxqLyRtVP4
8Ol0CvxACJvznCgYJGOjjKDhw6IsgPpb6uurmTxMZUiwndkNFCTVIjArp+JRxoaF2TQQ4WzwjbTm
d1IFWIxYdhivKyYqZD+dVWvPgWYa3OKwEOmM/QKpXNFgC0DNrKB7ZDyQWEGW9KvAOoMw6iZOjjxs
0pYy9Bb33Cu06xxM+p+RAZ1Hr+eq/ISwGNW4t8ARRAYp7TYEHoQj0ADHM5A0lRcRd0aAXRNmchqh
pc+LieFec1TCrmdyyyx/UreGwJeWnfRdLZxfcz6Vh88X9o0t7w04RfHa8iO8kaUiV3Eq81EauVZ3
aQ7KHqtkmXgZUB+1+IDklpubMzK+vVDpP7Z8zF04I6lqYJeALlaU2N7tizaySrUyhYL6mF8Z3K0F
AE4z65LkYvKzOsF8sF+wFF7ltHx5v23jLnpE197TQWnDM9WXiwrPwhtgOLaZ8rg9i+ucGGzb9S5I
2QWXKQvXk4AoytemQUBj4L81rN/x/jYuX4ZxfQBGeqau+rwQn3iUg2nxl2OfYdEh630+oNy4gIYC
A88Wck4/1fZ4pVi6oR4Hn3Fvl0WrDCi1h/fNvdCUZIKTCzOzBy8Av5BibmExWNXUe8baj4ilN0Bg
bt1xLW2tIxfamhciDkRIO5uZtsmq57HUnQk4QEE6KHxNDEdLR1F5uSBGt2WhK0Ox8qEaMG5AcTt3
n3GYAgu/o7Sd5VqKG+wnNml4gWy2QqZ0244i+UqbPgx+2vztEKSyJR5eqJR5bonx2r5AAtqdGwfe
fbXgzNSXKp8yumwHoZzomueqakrJhVHuSZ/tMi2Tc8DC+8QPWmTi4p1lHQAvpjI5gY0k+R9yA36v
iiw9j9rIUHAzYr93e5o32j1tCSMZmouREi7lr4Sanegj62BWEsCtPv70t0sjSzRzjERUadXlbgdB
6/uoltbLaZikbFMYlXMyBjYvGasEqY7GhY9a3cd8aeoxD3AhkxVsHDB7dRS4JndlKbCAfphripPO
JTOItlYCjlOlDOUarfB2SgDXefRQdpWTR65EJqa70dTQtPnRLnGxGUnVBU7c9eBkY/pmAZMabCDi
fMA4jLvnsm6miOb5WEDT+BNrBzCb/5hxysc4fbp6dYcVzg0rCs1XR9AHVXx92SpE4dzytx+PgmGX
c7aN7sgG07NsySvH/j9FK35Jkh6EbKade1BZS/ljkj0siCTOprv5O++f9wXWYujfS2iCd5QkC4Wi
3B53CtYemeqyTC6eb2qgOWZx1loM+BpcxTO9XKO0PmiM9GpyVuIkrf4rNzs4cgaflUSdt+lWfdld
VQdKpaHRqATdq+TpfYAtpDcS0yJ3lLzOkYamSDqn9DDtIuQo60G9rDtOa9VrYeL/7LgfK7LR35cl
Ttew49BGAPMfm1ShopSG/UesUPVjZFDiQW2Y9mbq30WjcWV+xvL+UywMZidWtfvj/wYZAlvir6/G
4vyj6nWO6Rlyo2MLrPqr7MvRIoItTzJwEMmH/8pIvV+W7nlA1nvfekR5xtuasRCXQ1UJAU4tS8e+
fWUpdQgcGSYCwq/f0qkImbN/xsvPRfjwNYDoNnmkobYLs5bhELXNmZ5iLwdCbR3SsBuX/RD008OC
weWV0/6ix2yuj9FbD5NUWk1rr1ZpVfFBv3IsyQXh2jmN8648sqbU0o5RNR9fxSJmacTudE8dLYvW
S4kr6Oqve5IW52XeZY1Nx/cJKEwc/6iBWH2QT+HV58VBgZFjAHVSVNSy8z+ocDL71q+YZ3o3EXYf
JRt/8q7TPVANE4dmAd5fT6FEBg/+TAr4Yy6rZIzNSmEfWiNLkkVR46cRMRyBpc1v6D9aZyGsBGYw
A/YbbccINJAQPhdjVc4POXsdyiC5c6v8Vk0S6Aj/aitTxpGGrgPSid+r8E3B0UPA8rm7xfk14YGs
IpzyTKhC9JgmMUSVYaaAhqZTdv0vqVO0VHlLJOIEluXtX7r52kObii0KaN9oDu8tzi/gvaKcZxNU
+IvimWD0Fs60HqKi3ThSE7Jik0n7COdIpJ/tbtBC1hI2FV2goUNIBD2lKExSAIaear/+VEZMxI1w
CVkLCRqemnbpK1Zvm8HlTNFi1ByonAPkBdnBDfv4+ySmSYk2Dk4EBhvaZetgCZVajZKiWjnpnI3j
5hnZt+b/B3hpfxP8v0ec5Nj8X6GUODpGxiLJ0I7dDy/gXZzPr+JVV+BuJXOIb/0PVWOq3nvewMAP
5neU5KqtNv7KlcJw55U2Uj1TgVZfjG3JL79RlySWfZmMPxMwNW1ERZgOAfRlTmHw9sJbTn0rMUFt
JzJyfs0oDzTPSYZgFv32aF2aWUabNYMxz9mFvEL2rSKCizLncylig8RRmJ2//+b9DdCe/ZZw0ALg
MoDeQqh36EjY+eDv72ryI+DTmLEfcYAJ1YhhCbp4PpiqtnHbEbcBATSar5mtmSM2yJzOVHXHD5Ez
OfKJOLyARYDyAt3QmvpuvwLiKQ4P9VR9Hrha3rFnY8nLtN/a3Kt2KisgVjA4+xD6fZPSBQ+DLXCr
VU2UhqIKDvl+sMuCl93Zq3Ecza6wsRMyYrgTTNwVFfzlOiWwmxgwJ8GDg9sYVa8cJ5UOQQFSr1t1
heACwnvhCI+/OgOIEqvEDHESOmv+HXyxy6BMY1mUGVR05bf0oq5yMNxKeHDXeMjQUii1jc3pbc3k
ceOHrJ0ERVxl5ziMQszkTF8GF11vb4RD1S7WRiUXq6nF4Lcsb6Qd9m4nTjfrdBkCUFlv/2zcNeUX
b6snsPOV7vTo+dBGEawco1sZMGyNrS13MLwM+rsafsKmm1W3NUw+7441O1Z3boKYN9QZ+/QJO0hg
aBTRw6zLSSj6+V28NdXWGfSrDQp+/ng/UfPUFb5++7ZtEFcoZGhyAKTV8dMkZ0GAPb9BX2UJFmaY
X/oLFvu3NlV2kpBF06LCjqQLsjzbdFS1yisRktMWl5A9h24SDxK7aKad1KSpgmOWnW8DHFiUPj/A
c3i3ZQrzVDrIq/V4iO6PCNMVcYThmlb0UnPcb9UITKXVlS+WAbBiBP64UAWMRFdyK6YaHvr0msRZ
n03CB1OVIm2mlZGRncjXFowQ9d8k0Xv7E+yZONe/JMsMa+7AgflZTi6I+bMNqLvbUmDJMMEbs9IG
YEtrQuvp2kNd624JXdKGttgR8Phslc4UJWFEAJZxU+RlAC4yHb63nTvLwjDWdsYZ9lSRelyqp/F0
hu5rolAcLK5e3L/1JRQS/ENZPZ7LNGv/D2Mr52LW2wwCmiqNUjD0Sl+5LELAZcyb5lhXFlcc6R4+
ohVsvXLU3QLijU2xMzkwbSELGlFxMDcEohCiTuw261xiVuDqD0RWASDTQrAU5cnE+z8qjQ1cW425
AKJHSooSa7tCkN1QldtTcwpOoI35eElYC4o0oXkiS+ujzc5dU5BRGP9wJDeBSEzZRX2oLr8EF6ig
3/W7pIhXzFgyLGP1ufIP1Zs4DBSQpOf+7/ndTd+Hi2O1nr3slWepBDK4TMaITUro0xdgCz4Awg02
6S6f8Zvd3WGsXPjGJupjMQa/bkPVSBbvp0Hw7s5iu9wnN3iSdlrXgYEH9UXySSG2VQL7tgFfOQaP
w7FRGgDURxFRUcwGiJ5Ar1Lyhl9iYENzB2E0JfDv4N505s1RrYYQaDoV/0KK9HCaHdFd35X1waxD
w2IhUrAwDNgpuKntL0DZjgxWRIily6dPTq+x0IUHwLmJeP4jXpIcCc2zXDGsqW/rJFiN/2q1YGVj
K1hPi+WjlTlcCEJWKK9sZ95PXv+sWeIuj3YHxOHqY9b+cW//ukHhOxmDNHKlHscCt9abBuoDq/L5
HhQA9qswu8CDBacrhzEIMdZth8zW3Q3at/UXxAWt8YpgDrp1s699yZrmMo9U4O3hiXQ345kZTWP8
+JHXL54hwFhU52mVSqViVTfLP5WecgU+tNz3st7yklE0v5RuyJ8267eyhaa0Xx6AWfBon2cFisWR
wF6llXMTPptP/zNk43W2oVpgXiRyos91wYDH2jS05JN0q+bFETHRkR7RRC3KwYe8K6OPwVhLVxSP
Gz/H7LT18pYHKFFDdPOFu1hHcFtQnKm6YU0f7jeHfZN5WWg6cupzPMILRcobhSzXJgIkutEUQU98
ILXGja+NtOEHQSejBpEKHyhkJgny19rlhsnjbmPlcREnNVsYiBXJfJDlNBfIQWrPh9RTQWrQisXT
TUuWMiOXjSdbl1uOW78QKBFxwmVRxAOkfwqppyiCYkWs9lfsY97yTE2GQmpiAlqKP/kblCM7lPAD
Bzy1CPQOxGT/7i1fvmGF7ARkGrfaMWL/2d0Q/5GIt/iZQiKICRgm7NbwBlMBW8Mq/Wc7ZmoZy+dH
IFzcatEL4rOYpQLunj6FuZPbxufd4wrPC4Jmt6qTUd8WZoAo6888f2MSKG/QBqklr1Pon6Fk8VGQ
EbEZ/3JLZZlvISsWR7m/0xQ9naDs5s+cQwfdq9RbSjbubbi+3Q4HEfKCSTT5nvvazRwJb52h1OKm
7gROQP0WN03kLIKIv/dtbtRYYipq21XOuaUfaI7FI/WkSS0qx8QvL9ClryfO/RPYrYjpn52v0Gfg
/fCTrb10nIRItI8sRtGufcOf1X0/gYHzceU/8ujko8wSTGyvaQzOJ4owycKZccZRtXf8XGe03ALk
QUXsNV1dJImtS43cQOQzCTvYqEqtwxvxdWTvuLaZU9tA7/SvLzCwwF/mruL+D8W3ZRzGqHp70+iN
AjR0faeuH6/DC9AL1yKzx32b5hEFQRXqSUZAaRohkPGnUiRWWiGHNSmewmva9vgo6OC8Ni6qi85D
bow/04ZhcHiT6uyOrJS4DyEjjy/0TxStMgWLoT2ZE+f/bSpF9hN/fV9AYcGjAYPvJ8fgj2NX+IST
qZcuWOR3NfAfo+yui4Ooq5D6sPow0v5gDWXPSaTT1DqM/aKg29EQyn86S5hZ/0CBPbz5MXl77JVX
BnoFwepNWWnIPxKJA4R9a8fW4fVF86i5P8Wcm/d2NvY93LE4g+l7jdEiVX/lRgogooykDD/KicdV
Hzooz8lGIk4Tbm3C6f6AjhkNZfIBQoxV3LF2urPtfrTUVWgjcUbly5JJgzNga6eBzxIFiRk6PggS
53dDpyXLE7oGPA5g3EVjsV22nxj0iY5epDVIA+UjYeIySxMomDX3PJKIafOt3e6cp9a+aiZFmm8t
FUGwzrcIjlweWphF22AmPzCpAzmeWepLmWdIyYdGurLGqYR5iYGIPI4Z/4k2V3Q+7YkfVW4HpGao
CPFHOsjTJUlUv1OhZsfPITQVembtd3sOhF0RHqXSXk1BS4wFB5DfOh/qaVWtJteMGHKMtSmQlb14
WxZFas0ujHkq9nXxnYBX+lubHfuNBdgbpiFsm7Wnwty6SQrGKJs2QciS/z6LHmv4qyOeymRVKhTy
2JXn+9cfs4fnJUwGE6vGo41n7VC48cMn++9gigP5ZUzVqY6h93fbadCKt9QGDar+jgFnkJQVPLyF
NCFGtela4T+zKD3c2OpRCel9hCpGQhhuyLuqFqhf96D8h1SJwW6ryHJKVeys5t1EgScpmjWLtqnm
SXdo0rUqre80HDF8OxoiMK+ZzmeAavlltKPnYBgLuxIPr+grSSrZotmoQBQ+3Pae7xYqAqzL/ill
ddzmw6bbrIwwo6TZNo8PMf4CZpd5mJdcPfCOuQJOJ/jREM91w0JAZ6tCMv/Na2DR4tnGUeT0fvVM
qYer5u+DKHpx59TCL8BeO6ORbolqyM8jkv9Rhyn1NF/S31owjqzsU5JzGUPIXg1fGfMvnNG5BOpr
qXplZbBRFbV1oGwnKeuV564Qt+pJPoq5W+LoQptwOKE9JyyFACIxdg26Tb8XR8DAHYRFVmsnuuXK
0M3IxOKBRK05ndD97pyQtbJwgtr96OTUXkrWkEcRpN/OJaGZgQxi4xsOUmNNXR33JG85ZI0InS8n
RISKlzMluuI42F/r+7gYDZ9N/TKg7HRcAU/tVw4y8p+btIwz2QFNCdV8vY513MAwPx7PhQqmWUkk
KqtMdCY0bQnsqqCHMUqoyOvJfLb/5gl3uArFdemjc/QxnLdSkIWH6Ew3Sk2OpPYtBk71gt0+pb/s
AScQXc2B8JVoE2DXNR3RVAWIBF51wW3ZUE1s11mDSWC45ebG4Yk3CpCmRCKa+MPT9eNV0oNuKeAR
r68jN4S86YYKvz3kGUAKhzQKlK+wGu8BkykSQNWWPoTFky296B0oklLvYnxZTpkYsFzfVEpvSVms
9Aj12mv7RrKCvmt8chnY5Lv3x/sxMczkRklnfnT2dye9sTlbQsal6YH2T9Qw7wmpBSYr2QH6w/bA
jm7XzVOJxYIuaM//1iTy0Hm8aLIQduNG0B+YojmYJDmW45mrsZbU5mp65mnqZaZ0DNsAWYHwnMTX
OE8omjG92n7diq3wW28NwQz25EwbXGXq8qt5GYIZtv6pwjII5QS5WtVyAME8P2DsuPDvWm+ji3SR
2mD9tFh/hY96YF6LX5s5VyKn3alXgRFjcmh7oM7RHyMAdgTwqX8qVv/3bE0M2aKJsqr6HQhkcxex
ieSVlPDhOnGJbUhPmOdrIzLXDmOk6uq8IX+CXjm9cCbcSZKxbSbXF/IinjyOlCChqkpRIc/QumfK
8M1rcNvxpjIsxhEqiUnKbukAxT8rh1JMRRsSLwXMXI4lU/QKaqJNSto2YdWaCwpn0NHbCVNPsiMP
fslsDFM8eVVPOe9smJk+385AfkkFn4eIQr0DXyyHT5ZeQfVFkD9OfnsGybSMJf2l3o2Q/F82k3LE
3oiewu5TE0OzmLYHe1xbf85DTYfb48B2AfcBAJzuxru/fR5B4GCpQpHpw7z2w1dDalWFNpjXzMxu
qNkqsb3GXj/Q16BXU4L5n608qZvgbJ3hMBg+LTx0Ad/vhSU/ZbYp+M40yki/ccABrSChjZKFWqBB
fX+V5Jb6OAVp2AJxtNlh6tIoCrX6KDVd4UGFNSkWtgAwiY7fSJh3d9YJUGJtz/ii9gJbmQ6axba8
tiIJTqLGO0/UT6CzG8vVaR7Mh2RCv7XhGt4B9r0FDT92Qcakgo6V6POW7mcRhwmN4pzz6zSqlqIR
XfdYeyHGhDMk59VJoJDTg+7BD8yDvJZh2d96OpkfGBExwh5npSGSV9Z+O0gcznNYVtfgs2K6kqC0
c2fU6WziMi+nZfGJoN7nT8tDA2inMOBYfnhtSb+as/KdMZYArTm6PrkGOVMkakqnaoDxo2XxGoKn
FpkY7HUYTMZRxk1mK+e3auwUGpCVfZEwj7y+G/LTBsjtUFWRQJlPP/mS7twN2AXO+z2LYqB0f7r5
Pqve3kMOZEj/Bx3TrOz654286SMb3ejEMX9s8AGIhvv/7X9c7TUe58fVm/qRJV9p3oGaUgHo0Gkt
E+uUJOWgBV6yH9iRaATZ64gvBd4tylnHegaYeCWBanEM+UfZmlEHD/AqlJdC9Geg44nkuu2FG/un
y6suSJVGN9DLE0GhLsGL8O3T+vv50JW3/yIn2wPeSU+1Ncu4bjz/ubqz7sVP8g284teXCM35B55T
bCYF8RDFfF6b5he/CkKN9YNyIZirpDuf80yp/W+z2vSkA7mvd0SWS/GykRzsvmGTYKio9vA/minA
TfEsEytXfi8NOQbikxeceqNXrDZaCOLZQilxxQhIG/Ux8wRN3wJ5Y5jBaIPfrKCuFiKHg1lXd9su
4wSg1apHivUwIHkh11rBXjIl1Tr9o1YRB56Lp9qviGidgzY5RLFRJh6GgGArs5AVN3ctjgG7WBGJ
kMIr5pxF4gVNYmFSUwCJChaWTnwsO0xOFg2TxiK3C8sfe9GZf4QdOfMkhjcdPFxk9mt6e/j3xJiM
9YeMwg+4BikT3cRLtpvG3gycyCG/P2cjE0nWCM6RaPyFNmqWMTcKpKDI61xd9J1IMn3eyrCrVjlM
EIk+Qd9/i/t5qc4nYr76VjjxOA2T9skFZen0Wcpyo1vX9Za2T3geurrPI3b/ON5fubaDZCpj0Ndn
eUWSktEHp8QurbUP38glI+2q6BkvgZAGiijxevwYSrp82WNt5p7t9SAeDPBqrWyeZWFTTZFXyk3O
Ty+VE77AvHOayzfpzRzwrHvb6lBedZLUnWEj34wOgrj4dLVF5vvZOSmMLv5juzswWe13pb5Sl5Xk
FlvH2/WYhD9LPXsq9L3X8bMPrm1m1UvgHjTH0TKujjcJB5NpNJK9sXP0bEVht+mA72sXei6lPMaI
2WIryi+Z4RiyPby7embMv4qmGyIR1d0M96BAm8Rxbt9+Nh16ksRRIM6aKjyifyOb1BrIraA+AKZX
42OWKveoY1+YHvGEyxs5H7cK7bx1UlDJCPZ8pGMjkB0+ZExaz4TU7jomaV7z/MhQ9DNYz6bJVx1r
IB/pq9ASCF59VskNp7mJxSXLnz46ZBSGGSkVI4VubvHayU06EkiJUaKTe1cRjm7cmwv22+DA1+6a
2Ob1y25oPoBjBPHnXBjUuqy04t0jR0ub5KhvycM4b61AOaRy8pklOAttsF89fr4DqWzLoGpU2hNV
13lFKtevBnqrt03Uvw4cfs5iZOaQPrAZR7yELYaD91CQy6nmI8lfmhMStUuAuCTrT9t2rWAdhOhl
bTEIrImXdSc8ZlSqfXYKJRklA0DdpWPeC7/RYzoJeKYZwAlkyHF65ajR+M0W4G3G5gWVDKRBN3Mm
rS6Odp/bjxwf4j6g1MnKvKpYunu2wP81JmPsNQWQ/eQwfa5551AxU1aQm0hLcnW9Czzsfe2yQiTe
7G0LBImv0X/sRTF/QaNZbhEYW/IGPpHV6qni6S23jJifUS9YJq8bwzlbv9hnWRnIROt976J2XsgL
zWxJaLDOasuL7qz/+ZPvw+lalDVERIzh8k2YsIaEQTZk5zF5f5O6TfkAGamPeRaUPpRGwHARnLlk
NV8Nu9qlE6tXn2XtcJ4zEAiHo2tSbVsLN4+WVlzZ2lSmqwSC/LRfMAYPw/La9oC6HfJ6hHxXLCuj
9U8dmdLUZKom4JqYLz9VJy5DExfU+eK795jnwX0I6G1ECalPmSLWZDW3KzgKy7O111EYh+cCsLtF
5KgISYkNY3lQbpIqXdXZJMzqvtDStGdndvElGti0rDSfC0TlhSgzl2MBBWkvO4WTTJoiy2Om0LHx
K3pVsXo+uNktIopgt0KwFQmjnhj5qOCZUnIInD0v+YeEYX2gwNrFyhR68/FHob8EVjjSjABG+AB6
wvNNrrhnaUBvDUoFulkEV5Xv0YUzv2wye2D7OoiBYzWyZYM6Im5UMj73ReSIOBSbbybcMfsNVx/U
mdUcwyQUWrYRvnfSSxDDUO8TG9hCOIn1e61utLcWLCr0ai1kmHRE+NIdG0RBp3W5E5BqFaojZ5vY
BSIKuxAdNpHBaM1hpO3/JXgzYPxWzmNGZ5vyZUR8aJ5qqTeIG5xvX1W4u/cVTkjC4TlaKc83bD3B
IUqdl3y1n5Vj/fRCphzk86iEqRJBMjzsMhvbMx7aTJROfiYfzbOCmhxnPuJ+us3GRtbuvLngnf8V
limT6wTTyqgqayzO5hoR7xtngITQaTocDSpxSr55/reCDTA3HEvKhWH3tW0Tc9BuzN0WmDfDf195
hAA6/3KcHdiInZmoFirvLHEPubfeSZ7a+ZxAb2LYyVa/LpU4Rc+GehLvVinY6BOu9IkSK9orj9W6
WAiKIKpsTCDUyfVToiNcNCQ877n0aN13z44TN4Py6pLdTOlea8bKpyp+3CKP9VYbJMLGNmPPTAdm
U54ziV1ewtyy6itUMD7TtAxMnwhA59YXUBb78FMUAvrJamoKJgldvBKaruwxthH4RSou6D+l6ayi
i3gfewFZAcwyRqyzcZbA8GV3cdzEAZ+tUA0uRtOwR2P9C51LJ3XZ1Uooow63V+v+LhDSQIXs5QJl
iEL+rIauxRmaOJ0Wzxa7qaeogZ+YlWJqR5Pw0x8jyRm/dJ+0c2h1S9+LKyaxDtS2VUiW2g065tZ8
akpi1UUiFXSP4RXpxcIy2hH5AVwfC1Jhf4vQnS4J7ITpsLUMwk2K6RIpHBSCcFFE0hXHdoUAOLAR
qTDVHM0h0ZyKuBPNIJUBGGQvyV4tMrOVYEu81GXftgpL/mlDpCasjkGVfzEqougXlePANmgtO3kz
09HpwbklWjV24+jKnvsBuH3ZLXGtyEszWBQTTbX+U5wRCg6dSXrEY/95bEhQUM1Cc8BbvCGR/ROU
AgOo/RRixoART3R72fFwcgaq8ExQCdDYNpHVIhJzPrs91ws/q4YgqIdF5qzw1J7PxBmSO7cPwrnz
vsqw4+ZmbpmzKDeMlZsFsPrnGJ1lkYbNuq5pw1ZBYO2vAxTBd4dR8B9a3BLWqazuzeTamZh41Sn/
4zGzDOTV+OrUte5+7HS5PMRMpv6RSw4oGa+XF9JzUZxum/akZB+6sBaaqLotZdEzSeR/yN8SbxoX
JwFxKGKaH43inF1lHBvDOjpC1Q00bAOogUQzhJQOc6Vy+WdsvM9qTsGa+4Fw5+pDUWpdtOYyoPI1
KwdTIVZylpH0o1wFDnxYEeKF11Lh/uWHVxdcoLZJScCb3hzD588vW0CyQ0p5SWfFvhWA3iYaLz4F
R2+ANwFjtmUfsLQMVoJD1tlJT2naj3PdCGGpXnO/E2Scc6V2OuHzCQfpwM2AAM0uLfvcpsJO2dVl
jHGUDZ4mCJ9AfRt0m6OPVhK4ESO5AESp0SzLmgIY/4wSMdXFuGk15Kb/tq8w3jJUD9BiSoMGHSLS
3hoM+M4btix+zBTIgA4AwANz10AKSazNNHExBbmtYls/RYE7mpfJWDJglMFmWLzT+eNukLY3i8SM
XRPYmb5Nt7PKuuhTI8/vpvjT8na5OEKNMD3fsMmt/BHDvdbXpJE7Pg71pkhv+vyLj9/UtxFdLVNp
qfl66g1lRSUyXa8c398FSS6+EPH6Z/nH+/VLKcGwoNqQUO2h8ciyGKpaVe444m+qC9N7vKH/l0SB
vjeYeJTrSNa1Hnvq2Eia/0+/0M1J9p2vmJjkWUoscHN3Nh1mIthD0a562Phb0CKI+kEgHN4KDTR+
IADuQcwXG188s5+b1aMAY6+diwWiA5+rB1UZB/LfzhgFRwaF+goqRKw18oKsEYzAJ1MJPF+JOcfc
IDm+AlDH47GWWUxqBroOQFldJQ7qAHkkbp2eXuI3n84+Oyrm/6+s9JZCJu4oym7Lq8WBd6iJKD3V
knIIBVz018e6joPtk87S3t8Y/EjJ50YPR7/BtOHGoGdgjUEqDzrjBiet//9G9W2LhgqfTazlickq
O5urCI0we+9ngrICKcUyLLqF8DatLqOG5N6FeSLwx53eYxij/jt1PbrYbP/54PjxCSUpLkqDWujX
H1btKMThFDwkeWqNBtFqJpMOvtVekWkOoU4zLeK4b0HHvd3R7xZAmUoNzdqh+Kmfr2H8XfHx/AD1
zCjXFjULVdQVbUCmazVDO/2pmW/UqMyEj1b9a/q+cZjakCrcsVZBgIFQcJ2auZakDW+QnvI3oo8P
ro2Yk6Kr2eOKfeTG0dI68zjzfSprYqyWYY3n8eVuxSmldhOHSd+WIOkOnmG5gY38tw9bNuYhW5I0
aOjcAzKMwNf9rQGJQo8jDJgjJ9m3fChbK4aOJz3mFkhdGcVYQJyYADSIfbDc6WoRba6C5VwGKPns
HaYNnp9PH8uWZ6DVcFwOaneJ5yXPfk0EF50/sSg6Me1zxQwRVSkbh6DVlegSlXPzWoMYoFRTeyf2
bxcHQ9z7E0pCZ7ETAFvY6K/By4NEJCY6RpUKFQM13Tilxx8805rjDriiDzkYfr+6Q00qQNc/uGIH
0lk55k1tWc2BFC84EM8QY9aI9t5HxCCwm5syp9W6rWFc4yKr+Nr75xEKt1nSvcC9l+hFbfiA1WSL
Z6KIGBbRc0e8MEy45CAZJVZfKkO925dJ9uBsSmV34fJlJi02j2g7fablxGAQIvijU8cTky23f0QS
cDUoatQRRepcw/tOCkx9qQf3aVNUtYs7oT+/J1pWOzR7Lktd/lX+TFq/iVc7G6B9o2hkqDXhTHyv
kFsuf6BmzZfhr3kx6rbw9qAB+F8qq9jI58vkoJ1R9VJDz4CLTMfmk6SkJRMkM1PZbWl7+EdFKuDv
b0ld1RBMpbEFTtf+VSdA8MXPXALyP3atZKWVFhJ7Yiy45fLk//1GWpD6Y017suB6PGJImPaZN0Es
9ZY8Ni0BleSjb6wet5z5iCVFLdW3UC1W66v3XJGy3R09QDgcbIc9GJQw0WawmNSbfQB0UvV5qA6U
bAkNeTHi8RUfKHm4OKkOKbOwQkGc/6GDfuaa8OcBLOBoOqsm+vRgtGyWR2+5YeEyhpneQc3HXS8k
RbdQoxsaFC2XAci66+EKNS+nZ97nULG1L2nBpROr0oAg5fXn2oCHxGTaS7UhZ/1hCxek/zUfQBrk
1UO8IE45QxpmCb69OJ0nZrDzjxFzaApDCss4BWdMo3xMgme1FM8mhoxoKGJGnxLp7qb3aIG37fDW
7ML6w9EVoOlmkNQWSRAtxHZSphZKG2VdsOJGD70FJjRnx3/ZFU4SPUA+zjkU90rzm6mF2x2Iy964
pvhzLmIKw2A57zX67PYAoJd1Uxk8sEen4iN12tZPOUWn1ZVbYi2sPExtLN8GEPQ6wTKnyRx6Es/J
9aNHMeC6GQhfU8QVrC+pSTvV5r2CsWqXSFwvJd+Y8WKOq7azweurTlDYoqaN+XmS/Ypu86iaJrS1
pErjdc8kQJSt6wA8knMCjb/1I5qOmsz5xqVrPo3DG6T1GB92DMMWf9sRZMLmodt+2jt5mDULRcqg
SfuK1z00jD3eRKtJZQ2P4w7lnXCOZT61gBslpSVZhuNbqPjGtc5OiQzfnlB9jsVrmjhrecfj0Zjv
t1ae3PbSRQYE+Z9Gp5f3M+DBnn5ukNIsSGog6n4dmJaBetAiH6pC7BydsDZQwWz5BA6pc1dB3Wnp
AN+ds/Q2ZEZ0yk8dhXn+DoUoLlM31NVD/5gMXG+V3tq5TdlSOolxx96hFkJRBL8o1Y6zNaRkVIlo
MeL0JOBUoURXOoGnZJm1NSpdfGHvXWSDTVJcrBHEZFh0h3xeZ5BPIR1XpJxLsgMkpWgrHiutKZho
+JKkqp8iatGmCwbomACPKnv413vxtwbTsEZyQX+nroQ+rSRKSDBHo4+jeb9ftU/rml3NqOmY8mH/
Uk+EKYap1kS7jMhEAXQhle1t/7kWEoOuDEyo+zWAFxUjjUIfqZq2toUeWB8fLxLRCnPiL6WF0KLO
oN1WRCqfAHl1z8xLsMauaWuMlM6GOvoTOI5J5VGzWClQsVNwmVbaOcSY2fuJeF8L70CHmf6081TO
qvEydm/qe7CuvR/X8D31oREu/Cw8/0npIemonIxYTRZMYnt/r9MFy4CKe+LVKmTnajIDIFDWTBbr
tb2NrGFZIwGvfFtLvCBsGi+w352b7q9KZ4cJz/F6zp4HGBu5nHK+NcBCyJn2p9iu9nVcnmZSoliN
KALjzDgdz5RMWZvxyhjhwDP7V1WTg2b0DKM3lZQkAgajHoobT72e4i7433nBC/wm6guSEQPz0Wqi
L6Ez/GaAO3NWxaET8Q7eMOndtgeCDSGbzSXjNdYF35rJKXpLDynNMgfZ2Oc1Q7cdYoEHGytNzPoB
lGIkivYOo4bZhJsFGtqSx7Mq8uWWr4bfxy934dfvNfKvE+XvB+DbO19ZFlNVyIUR63WVh5IcxneA
39Iz+A/Oa6l7yYUP1HyN1Ruts1yQ3k2OO2a2WhxfhHgpiqWmw15Z7HipgZopLoppBCijdXxyPfQh
6tMpORJCO00md/knL6Lp1eDwNO/yS6GpHtEj8Ii4P7LKJhoJZS7V21NPngPujgECOEsYBrL+54Ak
nnJbf6i6iW/1jwkkrQYk0Zvb9A63xA3Z1JDpQQvKnr97cLUZ0E7Esjg8s5lQ61PRFleCxwmK2uL3
ErERQgKXW+ldgtgT6165k2amm/CQUnTYf3SGAyz60YlFn5GuZ8iE17TWCEbgub5iFXffMyuy1f+O
I+9CxteMdMwITMINa0iyUTKDdfazmKIzolvc/l2k9gqNNiBojzi1U4ta/wJqqHvP837udtUtmuB0
bWUtfsVeqBBIyAMANm9piTzicZjksnWOBlkneX2s5qJ1guU8x5pQ964TUn//zWh6f/fbs5YwbtyN
4uWyjgrcyZk23r6/3u4W6pelnmYoWSSUCjJ5F8WLY2quQSB/zYJx6Qfgd/KCUk5gLLXIwS3F3CVu
Oo0phm/vO1zTQ6p/ujHYgbmnU3J7+a0IARbcZJOtOv+MtQpZYlrK0ec1ANHA1aQZ+1k9jx1OD/Ul
5uLBuacc8VVEk0LzqkwA3D4cg6jiexS/xRoGi0aOUIQOjmFF22ikYDXDhQi5P/2/OkZUbvORQ3Ah
eNYVpbGwbraoFAcqzfVsRWuunuwUX+10if9Ss7RRGOvVZ7L1kum7kPIt9dHYygjk7+7uiaWFzONE
vN4pNZCiRToiRAyHPZULM2hqaE8HUmjoYXB2mhOT1eZazgOhBngxVxzQzM4MM9XfL0Ws3XOQ3Gal
Lif9kePWdVr95v09huILs3txBOn7z7m86yxGf/xL0ZDBrW3ouIN0ux/vmV9EButMVQpN4WiY5E8Z
6bdInJi89NGH1nKehKED/nCVZyY94z8+6NUlaQq6QU5xWM1qibcAIelnGHKeaLT4ihUJWEB4ZixI
GA2vrd6xDaQR4EUpPBIhOjD/Hj9Bdm9ZCF7NROqVbSiQMZ+YgCB8ARlh5BYkPCvWxkoapGYaLyPo
ZCPnHaDhXglaQvDPzBQSlKQEaeTv7XvNzCEKccuzQu/KQZeuGW/mffMwYbWZGyF3IRLkjPo96zdL
NbnbWpBYoGvEFeHcA0I3fgdKpv2oOaUoVMjU1AS6PVod4Z1PXmr1hUOQytQQp/p2X8zaZT2yrRuS
wxyovX4YMBKUZ44fKjzHyE0Zdg/kC90YBdMjJyC5eOsA0vzY45QPbbNsfbg1oVVIcRyNBk5dsejh
Av45THCOJZa7b6DKKs2YhnA6FmSucjitQ8piCnCnL+YtPzkGjBu+f780XVxJyozO323mTdX2Z8Sr
MWPDbL9f1ypjyyTbBJU75bZ2caKa+YSXJqKkTrozp1s1LJYnzzfKVaVMjUVHuTQSf2Oc+VwFDDnI
o1GRnIaoWEhYbeuWIkjdwEqyuaudjhhNeaNTeyRxiD3Kfi99b1Q4fgxWkZghISdc5os6zKT0Ci5c
niNAG/WLxY3LYjzlfdAf9S7iE3ZSGD5F8lNM0w1HN8wem+X48DQpVm9gXEetsJbmTfCyaWuByzIK
31XeeVtCWBJD/00JcIEweCNKxJ2IeMu8Gk1arCq3Z0nwgON3zHybKCQFJ2IdB8U8WsxGFqDffHga
N8JWEmzPtSv+5AjVm5sW1DGsJwFJdto2UEOJ7AnN4K4Ik6TEYkJMfSEsHBqF+oCiOL10qfFle7oa
8Z0gmlsm98eZ1e4/rFJM3Ux2IDECwCsCKpMSxcXrTZ02wEGe+5WHykFDt6i8XTLgjFMsXsW0qxLl
l8tefyZskTwfjuKBPBfDFuUR1MbmGAsc3cjbxWEvSVzQe7n5T4XISEGsa5bYzwu/nEVM7ws/BUWb
89VbMyWZFRMtuhQru7R8fuPUNlVmOm2nuyC8RB3lWuCs3VIjqHjXGcrLBYFCjNR//wWhdPlKQGBd
OsuxhHo1t2Z/k75uFolmINoeCKpe48YpUOy3MEM5b64omKtBF+V/k0lY5ZAzExyF2kYGSq5VSG/r
1tS+DQKCzEy8P8wANWx8LxOW0Y91k0sPXky+xf5SHMMGL1OLhbC+Jj4elZAsVL9eLuPOMJXSVMVm
1/+nzMNk/LSO/5iZ/+8j8hSMi834kfFhIiJ+KDiqnS7HgObg5wsN2+BO8eM6FLfxbziSMlc61hV8
irVzQzPoLptTIudeNjxoBEw/BG1hi7+63lNkvgtq2fGFMTRMcVp23+2wQw00iR+kjerrKS65D2JA
xhpmwmeKRfn1mGYXdVTH0O16mY0LJfLKph5qsDD6tctD5ue3theYq3+W3ANh8i3PIBUyFqdvmoAA
o/fu0NFiez+RzeVQ8peWX19292ogWxskX7F40sxWpds2UJmazJxb2onq19xE1QGYpk5dmU9gdH6M
hqDyqMztN3nw9PntimIJ9EyRRryfC4L8mVvnt5G7EuDcM5nnTdQPMYByDWTfg/AW1GRWXXnuNdWb
CubQmd+kYyUo2zFtXgwzrLCGqekl1Lsl8bUn6MZjz4hv3/WZt90Wwp4Lr5aC9woPScMxGZY+3v+8
C+xrltHKcfzFWBn+8dWGtS0WZsQKjg9Lenws8P/K6s9YgEBso3XakuI1x7tuOG1NS1wBbiqYcxti
VAcugEeQdAnWBEt0K6MXG2z07R9tt8f5UjVjeyRVR6RMZxX1gv3EQV9l2qD8UoBZnX3rfWfzBAeO
UgsmxBlxjdsB6Ad/3u38xcK9VcUsRexcY9ZMZZMyviDawpg/0kZCP8sAZ/2sqKfvCOlnnGiTqMYh
L5ii9Qm9VPo1bcjTln/JnxfLXgaW+1mtwSDuKEoYEhcLT5GEzqn+x2AiwncS0VnWj2Pp2A/zwW78
OuUtrCdgz5NEPbLHms3ET3+IXSp3SUOUTjVqPnEwgi6jqnXV4Iwx/UzCL4ZP1mX5JiMSBVBI0EMK
71otWVAVdPHXbGz1gMBFxmGGnCoKIqo5g1QeYi8zfF7qjN2knP6hhYmFHSIHUeWXdpQ1O2NjI3CG
lhkG170L6Yxuc2DgOQmogoFvcJ3GJ3lJLFxl/QnJE0UrfiihEkAYIbOryL9xy/sBIRiWJddzVcH6
KpQB4kxntVV6TpQryNeiz363bn1D4szA0pOjQXxPSZbxQ7MTaSL1V8am2inZWsuPXM7mqK+OYNqN
r3B/ok62DEvyRNPDvNjb2gGLIqgyQ6FJ93SJm6KG+LX/TD7X37I10Tsgl86ZFzwJIQTz1Jjs6UfK
AnzyLfUF6rkw5LIXdHZMeGW8wrzZl9xhWnOa+SZn4NigPM3XOp7rbMCFiDLqn1JGTql55S+2MqTH
Ejg+/HWv9l24iLMMIcUMlPCsnzTULhgT6oQp5AHpnCpb8SkH35ePH8gu5HwqMD4EySiZvaoEJ/Hi
EbWt5ZSSPu2WWdhsqZLyZzVtumR4N+GlPa6H/4g3zi8Td0QGMAQRodH57+FbsJO7EtPzbUTc6YK/
nYXZdZHfSM+Xk/F27MXyzqh183I0yP2zZSuZMpYXVZH3idJw5QhlPuxpe6xzQ59k7AN/CdOM87iQ
T6tb+dzBK89R5Gjlv1gsC8Czg9aiuuDNhihETXz+maDw6rOGI0ZmVnGog/VPJEbOILTmFzyJNbm3
+SQAMi0BbLdAp5/JkaHDBfYFxUw1vHl80rnU139QAcZfJw/UFOA34l6Ik0rM7zfaWoAytf8l4/qZ
mYVQlNaedM/cuVjrxlL8BCcIy0u5qYle1H6JnHCUsrJoouz1tlWUt4TtKrZG3o9Wdp6qJ2ZaYV7Y
LRoc3VSfzH8tjQ+Tn39UWQW70vOkEMSH+MVWBZO9wfq6z5kNsemHW+Qk0eotlNr5sLHs3gSNSYr/
/kR4I5hbU4cb+ahWuPcrb54DxV1XmuCCFQdarb4jOKig/UDB5VhEse+AhEM7j7HQkleX+O+1LEyK
HMjfkxQZKPFuu0jWL5pgHKbFF0C/IpbKaShYa1MMYZRqnmMcV7yurcK9hivWzqTaU/59Exhh++a2
+U9TB2wu/axsf0+oVEn+YpTfdYxyQkaAKhrd4zhwIRot/GOqaiBVOxY7QVCxaBq8du+9PaSDQZif
Eh7X4Qic0OZZ4kiGUPqXTwSy9Goab68SbFNcQYDkJ6XzLW0tMlmOxSoJtInWUlm+dSzS8prl8gdI
fB6knO0c6yTkEBBns5ZIOjSuZKjHnnqD/Hh9xhG9yDRvsrEmTEAsXgfhWZWNqEUPBET+z2/VYzrN
nylWAC4D8Lldqb8ayKyMjb5JtqY9bA7VPEZjGRXjEXuAYFbXOJJDKBFZFeglCJiCaP/kP5EznXlC
0ZXcIR2exvC4UaDrA0pJJFlKuHeJBtZK992uwyixXQIEjBez0ZCoERZWQ+xVDa/zmwD+SvpihwHh
FVByI6yhkxI4TpZcW7tXa+0wtHzJpgM7oWIuVj3xztnQcNlKUxgcXtrY+ls9IcDJ4QERuQgdlFGw
teYL3utzz5KmCT8ZRzzkRxxypOYUSCyIFwyS1Iwnep4L8ZKoPFeyvVzoqmzCd30kx8Solbb2gjaU
IXd/oeUZA/lFOm+lv1zmqSAbAa9nj8eVio0RrUZcMhjNrzpUbffx5Kpsh210qUZbNbjEvW39mSDH
jfZKj+bwXqynUvJ2ewFExzp02IomDj7/Kpg9npSnR8SWUKNIGft63fVeDPTww9alTZy2ImJJoJZy
n4PzuLafDtb9UrEeORltFrW/y/+KKlRKOCIX3L4S+1h0qPkoQ7YLeegGW/37ELMECmN6ajLfMnuA
wgQkVHWNxyCbs6yNl9SAK1anbPPZqD8JIT+irk8gLB2EaJfbsut+61mkfj0aoJbJwQ55oeDPkG0b
xHxYqj/vp3fP9zPhw3grnKesU7z4Gqi53ZK8DPrZ5WJ5zCQyuIt4SxN+Cl0VjeGPNeAJWCKmDlEv
R1q/xg+/vYarbCiqLnWoxjQmOjUHKhX+lQw5M2irFptz97Vt18GvKozEoLPMAehoP+dQoyCEYQux
8un45xanp/j9h6ynxe2yHcWUTovCg6jk3s8AeyDqcw0mTqT12/UqYCdjTyj6kyb96De/YNZi+UiL
2loUZjIRQHbh2yiggj8NV1pZ7oHLOk1GB6NStMqJX+WQBxsfdl5uZ+L2Nz/6ilTQDOaVbNECeE0C
osUTdEHb2+KWzQnvOE4pOAlmYeEJ6ZPiiZg3svG7Je6kt8t1vjCoO8TzlXDxulEz8ihdJdnL3FcY
q+72uY5m5paddlT4r0y9R6leat196vcser4VBB2m6hEHzoC1VPgxg+xX899rMSRw/davv/RcPre1
mXqPg6/cpOJCsQNR9P75EQeoSDohZPzFsVSdu+kI+FFhTQyxGSKafEUHBJLUpuwpo0ls5y9cG0KT
M3SJvsXkKG+95g+tFC2Gyn0b2+Qjz6GmqGRvrbek4LlK2PTrXVZcodyBK3dPELblbvKouLBPo2b8
vpZzmGQLbxMYgcM7Kv4wnnsajGPaCiovroJ/dG3qiQcgkzM5hRIfm90pun5ayK0plErn8UpgwLAv
x5OXCEjymXDmp/xfBQPK8L60wtTEilpkdD1meybL4dQ02hP/APoyf7nRBhIDRYSg51cMI3iOcRww
S8rOpOD1Lg/WPWPoVELYLtZlD0FS0Og5pxjMG884eCdjl1Wb80VPfYc7htyUaI6HiJK95KrT9w85
z6WFNePwy7B7iw/qOs/z9ghiul+Gni8/H383y3G9eg6N4M0ofIfsr2A/dttbr9ecqkt5vxfHdIQI
XzxHiW23+ZMKYdY7TycqR1nHsQLx54RimfDJj0ZnlOiXsc05V6bl9D41QZDyFVvW4gU6qHB7/nOR
/2AS/I/B3GQoVdId3sqNX6oLo+6VQepWI6+Yes4Rhh2v/4UAbB8+WBGFPkK7TJ1AWCVjwDoZkKgk
ajYW/PKzJy59l+POU7pi/JelRP3iRxZsRDcPKRA/7C5+Dpnd8XaQAag4Wb5r6+feWolIizY/h7PB
NjySpfZHuzcZtvUbUN5Ax7Ur5P3BY05kD/HifnBUqyno0+rWYTjbeTM5BX/TH+OGw5x60wMQpkZL
xGc3FPa7dZgwuyCrPHsBRMBKSUvtRwNJGXihaTBigiLx/fpXw0mOkXq8E4J8sV1YBmrnRh7ViQTy
rx3xoJeqOxPLRDgPhokohF8ft8MjBYYEG8H/tbFRmOd9lPD8ESk9gdXQZJGORqnRuJd7MZ5PUKx6
BismeQ8qTwAqPZIAdox2Z419q0oKCCR2VlcSuL0FhQc/SdttNSlFS0Cl6f852CYIBHKQ/RCCq2+q
af3iRfdn++dMbskp77mx8rHLdH8XSMqeyZgwWhrxJqaPaJsEjmd/dURilsQ2XGzxF5ecJPIlB1/s
wobs2LtNOMLYjGSw/NPysPKH1Rz52cJXvRN+ebS9iMuQAqrAArD8uHLCxYWWdScyqxQyMQD+KBgb
tHFZ67MSFPhD0bmT/8Kr8Jv5DQYWN8Kfx8vbDuANeLPyqyWU4DsUq1kx5anOc0aqEUmsvoBCHftO
CW8TbD0wkUlei5nyn6VK9R9Kg0pLOgQip2DQQZXBlqFq383zvXzkEfDsJXaBjyA5JCEWqSA/Q4Gn
8tBg6Xhi7ry+vLoAW32La9I274NYMwEBapz3dfico/OmLsIEey7GLo3TozM98TE4RXgQkEHC1VkF
CfI8wqh7A/f7n8UePLzMyMxLbY01bo26MnvFQXYixWZtnF/dyJ/rJno2WNpBAx4lWeaP92G7vunc
vKCUk3XDmikabpDJquj8TwpnLDozoQWOGhiD1kETxgXd2vUkRsJZLt2UbA/3cIKRdgKfRlAwB+t6
gxzq2EGeU3pS/OnPG/FoUw/DVkqsUn02yLhVuKze2rl8zZSsnctFpTzXjbCTR5orvjgXdzeAiI2o
AO0JtwYJv15dCK3zEb1TxNQeMnpYvlex2GHzkMCXvSde4CIA8Uj7v+WjFYLxGGM9b0+uBVrYNKRR
5d6dhNvu38tg+FzHsusyKhhrVyw2uyFsYx09bng58MwqXCAl2fGcw5TnqVw7xzdt+zD3GCj3NLG8
A11hZVoGi8BJnHyHOkRxxpw52Moi6LSSgCBqJVaikeef/VWZ2nwIXq6SfRm+xzZO9ZkAm3taK0dC
fC6yjjdbDIANwNPc4Dcqtb/8sP1GxpmMyHCdyktcNrfVxLzmAQusiCn4LF+1s+0WLQb4ZqOd3aeQ
RNOb42eWkqGGvoZUpyfsLZRFK1HdoXTPMyWC5YNEiQr9HEpNq+KIUyEmh5Z9BGQW9bYrIx7u+x2f
Y+uLvoviuCnsOmdVxjhLTqxWePvj63aKg3n/uSo52vDyW+kF2Wgt9faDQVWlG5nfatNWp9YLrE+A
KxPhyZ/3/jutLuDporZRhqgg9EhXSds4sLDYNuEsL8VtPrUBjYOteeuShQn+ubxexTfhvNacTIVW
I0/nJmaj2zgtj1qBuPcA3kmFvaWPHsE0psSBddm+govrdOfvjtF6d/Z8TKgTONE9eEK3QEFch1Xa
VXImeI2Z5LKsFltWB4CHQO0N3F9t4anylNuJOVxRCVJ3qNgmJCpo1M5r6MJio1WLzZVLJHKPaQ/c
wevNWHP7YxpGIKWSzb3mkS68FAFHuNHy0jxUm8JFhMOhiRVBwBsBNgipnJubydoJw9uRRj9XN1Bw
ab0+ZNn+m5x2Xa+OY1AkBA6htUP15w12N7g1TY8xJFzADhrMnmTHRZ6zmlIU1VQx89jz2uvIpAde
lhjKUDCAOeJeiRY1hR6sUlpP9mnUnxrE67TphkHFBPLDLLmeWuo/JBm7bpnOhpNV6OMIM9Dmdlcm
8avF6rBskHun0aX8pZZSJI41sOTZhnLikMyrYluFQJ9RGodXW9fz+B0AnB8XoCpYcDfSK0jeWgGm
OTHgDp6J/JTy213uNNY6HcY/azVXN3/rX3HqWwq88QVPxbvbjHYw92vhdszoFzH8cNZALjcggnh5
soacmg9fh4tjYdEZN3xnkijye40IBiHS/l94PiCJK3JvFVPDqMHtnG29Nigd34AEs4RYqL4uA/G/
Ad+mtlB5q1ZprV8QcqsgfKROfNfY6GIYQ8f7vL6BQ+4Ha427WkBoRv9Z+bJsuhZe7hCLpmAwWnfF
6Lu6k503IQIFJZdFywCxUh1LobOTN6TW408VuL86Af7FTYvdTKK/XkStHiyVjuAXChYcX45Xg+D1
g9jdCp5AtLdMoR4MXoYPOYVGQA0LZBPv+rIcL5Jbj58BV271ttvu6VtHvUZr/Kht/kuQlayQEPfT
TUVxJ9YFrCGeN5LIxUJnfjwLksyM/oyjGIlP7itqFNcHE/9MjRRlPJzdzO+U1td3QQ4n5HWy/6bf
1tIN5yEz7DtMX4LShFwaNS6V3IJS2r+jwjK9VuT/rdRuoJCaNF038FFIzhLsXFbCUkNM+/5yzYdk
E9ZniJeH/fihHOB/zGslhHumvpVta0HVOl5NmyNjlmHP2nFLogj9xDMuX4Ks8kVf/4INpfI+kM87
E9RHeTqs9JlSjiS7H83X5nxqVLYYiPqIZBbukhtXOEpnnVI+ng8G/7sQ1k68dgcgh0YusxjQksA/
LSEwqHNAZFS//PYvBktD3mD0Uo4IfKhvDrfyv9DpZv2MczYkQFVKa9Agq44NJWyfFIW+QcjApbRB
nr5tcud/5idDCCBQIQyMAHasJqQw0hglFaZgcfvLRRy65DmvRHBbivGmJFGsC/iJKxY6+IaLiRE/
FqK19pi7siYJeJrI3yHGj2P+BnIz2AQiXQxsKx8pdSfH87F/PhRsCQAflf8aJQv89OERS4EZi2tU
fXr7PcIvYXfc/bWvKSfQ6ykfC8jaPLmC0Z2XcQmVwUDuQ6J+/+QihimW/EJ+jBBnBW770Mb8g0Ig
ha6PTZruvJJpgGDBn1V5RONBPOBy8HmuwD7LNA19VA8gd8qw396Yq1CzM77QzmxpmT4l5P9+V4W9
zGV4aqL71ot1D0R6YyY7crqPkgi7H8lTieAmF1hGan3pQpJOnN6Ncd0NY7sPXfJYVvC2Dy63OvaZ
6ZDLixLtpLb9CSuWbBgbbV2AaRfUsfInLvohTYI8tIxj4V+zcGVMTJRpxyQ4rPwnX0s2q3zrXcey
5AVv8RnydOseBcFMi9Fz84VrFk1JiW9aMBfD7kWNcOoktrb34eAMrEBn+iecHSGkzbjcgoXMAKau
v/MKtMX7FQpC8cKQZTcL/N01wDnvwWePAQAgh4eg3BtZQ3MQZS0o0a6vrTkcVRrgSHsU9dpu5H2n
hzTRCwUoBCSr85ZP4L/pcbkYWjEZngL5bdeoT9cp9MwDjpRk8XOyHO1UBOhpkcD4pvst57+jYvXA
WLP5JO49P5DwKBn4xXeCzLUyiZgx9l/z/Mz1p4rDp4cn0S+WuW6AMqyqgos89+TkhO9AfcF4yNBf
QroLXOFcfFs+W9Y4Sa/t2Bj7l0OAebngkJIJD7EYbSxwAx1ZgMSCcbDGxvO4lsVFZXHeF/8Ezbcx
/TIGJr+i+imAes6aOJCcWReYYInyirvNL1jILWMXXw2mDtez5ASAVqk5pSDX9OXmrcdTkecNFm/u
PR/OrVT6vTRCzjKu21MnTtl2UzDaONSuzjEL/4PohCHgzSwzuYBxBX21r5x6suyuIoc/HQdUJBkQ
6JRoRJKL7/lYRjdzqoEbKVnlzoAXRYjQnqF0Fp/+u9+vkDNC2Yc2ELEKVgXaMPybhSLcvXey7J9c
XLhEp/hCDEtt2BwZHusWKT2Fl/ssvNTg2EmkMJy6sL8OPjhdDLzOYr0tC6S3NjMETqO4H1jrys0L
SInNeBD87fRCn05yuHFksCRrZAMERr1Ovj8Z/GfpYCYieYcuiMkxUNGnk0Sw/q0GKaCN0aiRT6Um
UWSk83wT0cumsarxoTdDFGtzjvbfL1vufPmFmqWX9XNjdohSdklmdiuLKzksttVp3qToZygcDVjj
3u+/IADWyITveaWSH9XBEmo13jGjg7XMOqtW04m/1syveA27GOO45UKuU8/f0wldRtLf4d9eaQkM
Bl4DPBaP5IBL2c4DvcFgTefexIiLTTtKnusre4ctWmPG+JFqcSP2PoJFZfbEVlQH/knSlGAs7+Vq
LL7x6r5BnuKb2tKt2OyAf+5TH6DhF1CwabWHzrlYboRzB29vJsFbGC79ZiNCZp6tqkpucKpYPy8k
fLBZa6Hmjl4CTTgtl+3LUZw+f7maafGnir8rw3rne3TN+NPya3WFDT7ODDWc5VE9Xldif5xixUyK
MDBBmpucISORtYWQ3uVGvSZxb10AmIKgOIld1kqmgc0s6eZr8b7r43Q0Oge3tVAyuuWWpk0y4VAQ
xRx5Lb73jiWIvjkmXAgYtCU/L+0GLe8fiFQoaGG1S1xRzjde3O2fjcIsctJPwVa0Wjb4wY41UwM7
6ImOmYX8CstUMWw8c5GKE2oRI7e7G48EdT/VchZ3vHIklTyQij0/s5aVTcHUNZp5Y86L7UKOjR5E
94U+xiwM2NivNb1EUPlmXqZD3oaq40XEW9nYfeHsH9q8OwcuMZJjifbnCH7W5sVmVX6WLSWgrrGe
49J5/qPaynKrAO9gK1A9VzuKiGNs2xo1mpW1tC4GQhaBDMXCGWZKt3VL6V+bPZXR2cG0NPummRbN
RE9p8F7IzZS9y28hM9QU+RIRSqvdZuSsiL5a6DC4157YHCiQEIlzCwqc6sFopkk0hwv3MMgsaOex
+nMdS2Vzb+we9mvPczFLsTLHByTer4v9tsthPxEYzagiYL/rPhMG7zNzPv3qMNbv2KfGQ1XuacOB
6xcIPybzQxep5WkapVtMLnd83mmcuKAktjECAvQp7WxzyOy2aO1+AfQJvdUXHGhE+NRIkIEe7ozM
gK48cYV2rx3wPVlYU7GmYJpVh7csQOnNwflUoyulCtiPFrenHTwctDtYPFCQwS30rCCdEnHNMPeR
swhL3/mw+gf0ZCbxOL4sTxvbmlhme4yrk6tnZUm6g4cykBOdFGHZjhs+to3OKFrjZRptXN4sybC1
FOf6w3lQYPi6fLpxpzHjKEE0jmh206pmZ4LZvKd3ZRRqXr7MU0MITjV/XnMY7Zi+nE0fQ0p/F5aA
+JVOxlTKPjLfgsstHVMf+ujWbjJSzGKGVtq8Ih41yPAoOAzqmydGDaG6bBCK+XG4jLYJ5Qp/92IM
T95HEegApUlqn1JzGnmVkhpoU2diqxKSreLoOrbq80OnE0wo8nfcoj6wVEQTxCMPxvLprEEz9cZN
ezO29NqxABRSPwuTWM1XWGcTiO1pJtzFF9hVTTh+pMUfy2wJ9wvXPfga6eUEVVPX8c43JxBCP6wG
SUbVjROA7/AQNcQlsWnpHQqv3S9revTNyIpuqjaAEMMzb/SL4EFa0e1IPgHTJdAThzYKazaZ8akB
60yXHUCLTsPHsQ==
`pragma protect end_protected
