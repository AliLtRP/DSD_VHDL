// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:40 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
hbKkzWs0Vw4rpWYYC85zdWvljKRe/tlV5AOaalYzf0tUe85n66AWBhQ5ACvE1YXA
XWLfIRiuTBYfhbXxlv03bpzgff6TgsNv8RabDeenBBGiUhn0UFUprmiZWrLFuTnR
MxACk0M5z9JrDa7uhI6IviW6KQpMxGodtVBZQcCeYV0=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 12976)
QHcAYp9vGwKratfncRtl0urBvpQoFMTDxWVpt44TfbAdysQ9C4+BQxiNWJz8WAWq
SBsdoaWIZpuDMhUJ5aPY/1qxQ06omGb1RMA9R3FjSOJ2TF9cm0TvJtr+370eGa2O
BRkZ+ICaNbxniEF194oExGMQsig01PWAZSO91tFMph6gRNIx/JWMsBEJe6F9u3sE
wTcfb2i4GsZqrwl/arXK5w+YUadR+nhqAgJBr5hC6uZh6Uh4O8cbG3CNozmDZCEf
AldYz3DTHKPuXFgn3TNn4oP9Q1qgLibqiovjh/TqdpCjyAMHFfgOoHa4dl5I1G8X
TVumCTmypWwsQNSG9UdTqdgKOKZLM1bxaxXHAsWK82+K3/iq3IcrnLsfz+itYSia
eFQ647c6hG+OUZoWJY/nq2Xp0CTZtHLg8w38ebgSrG5AWMEIs2azkQgDSvs0GYeO
T+IE0TXGmdKRgWHgciNNuK3ihtmypuV03cBjhohX3+Q6hh/n+NrapHa3W0fA6t0Z
aDZarpUUwBZKpSC+GnnrQ+Al+4jS1tSjJ8pzZBaLtTefrjj8+VpB3ptT7QKQxZMN
iyKs1DcyLfuDh7jZKm7U4HchqGJiGRRG4DMeFAag7I4Y6cyxl1GwWFs+ShYTAy2t
1PB4VKKhwUeKDp9q6wLy2yrPusLH1qZHWCFWijvjEar7CtLRyQ8yZNADYao/Sz16
uujySR+/l1xenDM971Go/kRZhWWgBXhsRO7dVr70H0uQaPJFaQv4ciMmFWIs0zhr
yEknN6JPFy7fyfeQ7AEzzDFgYT/ag/1yzBh31q40Pyxf+HZqy4UsHKBhmeJ5YMzr
/8B2ayDCF13h0ukALqx4UxIcrNGZvKl5kgXMs2QSnx/01SyV16+obMw+77ndUvhu
KBAQ4gMoeT9UGE/R29ZsJjN3gBYNfvyj0IAFQatV8NCcreNtppTsk5ZT6+UoxkVc
KWMKw5QsD4I8v9LBN3AQIM22iCWZsp/8CwvJ76WdMHRF0kz9cCW8rAtHDLvrranc
HsJiSVtKz3khDa1LLSQGXOAb/Cw4SpLteDL/ZjusV7Hwk4UxDn4VrNlc+W8ob0Sk
wyPuy3Fz6cFLTDRz0HVMoJx0I5pbjyz/94IVFa0JWDoudDth3dvHcdTTt4x0ET4b
p7QMlhoyBApUO2C3Zm9Kd5100/ug0nzsTnKT0K3Lp0ZVyjq+OEXALDurw2SR6/53
rlBQv3L1HUzpwoi7wRopagftMvG+ZfCHivQT65HBc7CstuKDfIOaDDvLdABJzCPR
ctMrfEIjmJdm3QeONOV+twJ+JLtd68QaEHP5uKmSc6wpYJrayzUKCUvlarCXW2QJ
C1s1q1aQ9mvxiA4js/QQmzwf2jrVYxZMiYlrfpah3Px1sbFkmaCq9zjFKDL+hKt4
14OL/HJIczlXjarxJciucVbWKx9R/YM0kg0Uwyo1cBuLXTiJNNmqA54nKKkSCgET
phn0TOGtxIWwz+TvctsHTJ+b2S2d127s4S1G0yKcsB1873Zi/1Vg+Ym9TU6RKHZo
b3lB/K60EX0Vw5cNRvrlKpx9NIj/gc2wYyWBOE59SkYVd/ytwVTKc6zEZlYrsN6J
DqagqM19ObiVWOaEgZX1VwkGjywmMV1W9ZXY1BOFCk+EZBgBOwBRx6pgO8mg9URr
RtWRNE3FLpYO6jYfsA8q2OKk3CYLbU/29d2yiytmL5TzGbgxglTZ76zTVFBsFHFV
2/nr7smmS0eJnglxQWfURrJUYAXrUL+NH7bTzfgWCYyeZ+ABtAAqNa3LcI6/fu4X
IAxfknGuZLMdhA31/4+8AtHqET1NVnNk0VxUkX1FmWIBTZyfj78qHq0W1S/Rdwel
J0I26mxyUu8MauCd3kTfmtnw5T+KzMPPv6OBFP3KmyHgd6rKPS3GOEo5lLJstjvn
h1K2PkhpcJkMr0aCxdtnQarXmdQ1vhR1GTJ8qWUsqF7ZX2SzDBIY3TRSFdrZzirp
6VCpARM+6hbIVhBiJwQ3AFu9fJJlAfobDYhP48VH5CJDqAQgh5UsdbYfR07/UUsm
mgHFkKEyPZWIXLEz6L65awzS57y+yYD+6OaFgZNozPi6mEpnwOFU80MlUnpF1fEk
NL72PuXP/q7yreg/sL8wJy7Q79Brq6NXY3Y1vJvjoPd6dVyVfrtiYlL0CSZjrLKC
q9oC8yc1X6AQqRHfw3udmnI0wa6XbGyJBBZAqXU1eeG3XMBsixQ8HHsxohHLE4AD
LJzLBFMQvdUeEAvZjfqotQTPECAzmHZYQCJErpH6CaAnG9UXpqmWAp6IrzRiruX3
c03wkkE1xObzVQWhGR5xH+GL5RLW87I3gQNs3jgW/o1LDtvG7XM++5xVOxmP4GV6
jOfTPnBKMEpseTOXk3ZmkXjVICOIffjrb8r5iasyhSPASmWZ7m5J1YX5wK3EW4Ft
AmlCBS0tr2BpAmdPZmUjw6z5KwS12f2ZzA5IJJel4hO4oDHQ/YMD3isPQEwoKc37
M2iXgu0W9pysWsz1gDWGLd1P1ZPY6rZn36+d8SmJkv1FMMAgR66QXXco3Ka4s8jQ
ZR6aqGmyktI8EJiZJBxvx+CGba8BXcBpj0EfjJJHCw7GHfcN4c1u0tcylMsHN82g
QAApE3SD5Mw4/otMID3jH5twx3m0jt9Ec4TsQ609+DO+Z/W+xLU0i3TZpZIMnHxw
fJ87+VXzudAUXBRQgc2KhWQvVMsActKd1qv5w4XKJ8ZqBPS5kM7cQMpEA6UVOK2n
NrzLRnLCMcHAEQiSmpas7qigquZ6gwd8kyZUwNxlnxvQ4Iomnb2lgB1sO038xE28
y9p7nqu1QQQsQot5WuPCIzYlHad1zOq5vXNexWmhEID8VB8pF8Y+inFBfk3H6EED
gFF49Zk5NAiNin+roHqKZta+3RIYaObkAwYQB88MrA/Ww2/IvaSOmxx1/hvk17mX
GBbpy/tnwQdVRVE0nb+Tri1E/kwTJAh6tcVuyioel+XUEOfllSSenvGiaHOeZxYX
Mvg+8Wlaep2lOkhnjUyBgrp4+mB7iQLhhe85CRqIEw2In+M4Gt2VOfg4ctdXGSW7
0F7dwzjmu56fBQgeXY+2sSDKRMvq8HRnZx5xiD4VxiU3WH7d4coDu97w9v4QqiT3
SLfrrLDx0W/4ikNgM1xV0Y2gi/kodhn7qV7PIyCeru799Pw1pIW+A4TUsiCCDX19
qBFmmFX+/Uo5A+8TMhrkeAIh+JtgfozChddyvDZnYECBc7/spG2VODivDfAsBmH/
sm2H2qdTX4AeTfhFT9gBvqfJincG9XZ+zdAg+qEPPAmqEXsskmJ1z5eTwbqJ0fvz
DkIgsPEGe8VdQD2JuXKddMzUMFSnmuCgtpeKDI8gGMoOtPwm40VA/a79+uVAixYp
AMABULsX1EpV3zSwejsVa9Lctk0awktMUMuUYuneOkbGMW182ZI8v1sjqSHUyg9p
6WMTN05BrPBHTBlKEtJ/vhKzCGpJlMHbwjMRXJLc20Tjoa2Iv8An4EDqu8VCrpJo
bv77n3PBf+S41TdCQgGdwBVAi6j8nzd2dkN7J8k76ZSMRz1b9v0dPG4Q4h38V7s1
yLAEwi3U4DF38Zb51BNKcm+MYj0SuNBKQxARX2lIcwvd6DyLaEbTwI2wC1J3jzpr
qGYXINBLgvlKNdY7I+GccE9GAaIn1nNvdz7pZ13s2aLYCEepCmvWYUcvoQItGJe2
FnHztIGRv04wG0rV7+RKCRoUahB9nclKcNM3JXGLdT4zFU6pumB/HhEUIjO7zA1c
Gtrbb2wsxYe1nzJuJtDI6Ng28tRiOXNsx8fEXLyWpmTp7pCGlast+87h8xbc1MJg
0k6GKve/bndzicAMPBkuA/+wLsSWr/76BKboGMfLeTXUH0lPq+/AwOOrvPoRMBV/
X9rZ54cs+bs5NL0LsI1EWcjHY5hUDEwjf+EHDGrDF/BjEBGUQ+9FEn3M4eCY4YGt
4/CGTuNfgRyNTIAh6PlgzCL/T5DJ3oTu53VjbRHhurs148Shdmbt9uHrHUW3HMdV
8lkImcnqwuDe+V0uCuRPnfZIDj6vYp6dOucN6YFWsTfTjT5cPXlHNm2UuJmi4mr5
5REG1kTFQ2EgSTkpBQZWhtFS2vUUtCxLaYXDzDMf/7RsKhGvZHjvnGYK06TJw7Z3
xCwZDQ2Qupbt5sSdC/B3Tg16tcO9ocETcdMcEtlA/11iYldjgglO+TVMUc0bL/aX
uVzd/cvDvy2RTVyiWFfjuDAm7lywbF62MZoFB11vRQp0lj0UcFymS8NM/Cvfyklj
4cWYlh+48AdpY9VsPLtuI26gzL1sJSvk0T7uttDoHUJOmiSdz8ucDpF/KLEMN8c6
2QeqUGx3NNorRzNwjMrx8ZxQ94SOJPEXujv4gIocPH6shoE8MMZyacewNH0cKcx0
T9/GuB94UC8NhnjDl6wxonIgzPKaNg8B90gWx/m6y10vJRKypmQLuUg6PHJe0Bsz
Btj1Pphq5kHh0cfw5eKW2PeWBY3238P0i1RykE6VogOVJqFTeLtZQs6xgQHCOG5V
H3fJvi6GfTmuAXGW6/PCOB2gGDPHxRzVNxkjZqvyFbYT8cl4JVUuuDRpXn9+SNlb
61bU3J4MBiwd7KT1wYcZNLWsWjACn9ClXvKzPkuMcEaBsbmopx5e1apwlbnvNJBl
gFbEWWGg8oH39qqAO0hF9jqpE1SZtAC63SXKGzdwfvUT5iH0cselhR8Pq8iB6+YT
EPp1f+XjTJweCqQjk2RzVxlDlLK0819MEUZAD8c3LHX04YKeyW+OEEnEfRNo7goO
GVcEK/FkbNBNfejc/ZHLAWCVFQicqpw21iUSZ8uYtYYp1ZT8JdfJtpHlYiG4eLWg
RymWpB+sZc6uQrTC/co6NgaQGem5EjrYfXxz2xG3r5HcLD0v6WWhtJravJKrunWx
DYnQDawrgCG5Dal9KjRbRM9qilsV/vgWe1geRkSzZQf2Dd+3J7OngAP4xcF9cLdm
X1ff1f7QIlsuOFyAANTXqccwuZSgQI+ly/s0CkNUT6VPvixuMt9dQDZ+rYB3nZfm
mv6mWjsQ9pq+acZy3CfmxAb2UasRzDs1ti2n2GQDa+YaDjGyf1RBtfIGx9b3LFAo
NBFkuhTMGnvq9gpwPEGvoF5tpJwPCuR8QYtsa9uJW+bMTCR3PDPrPC1KfRC4gVZt
BoiptE/Gv2naPkzFUnF9lDtx4Ph0YbhtzDSrNJvUuRLBavrKpv2a+wcCoBGre7C4
x/PN3XvnW0yikrmuedTlq3I1Iaz3+974xuVGdxqsa9Z0AshDisnq0WDSN2ktI7pa
tISwhH6npXP6dvmPQRRozKZ6BK3AfYdTDssaQvfo2L5z1f155otVftNiOtaokFVq
Aa0FNrJtTLndddyLvgy7XHXB8AILPnywVM6Pi2eKQL8tBy03/rAew0LxZ8OXD86E
z3p6ruIsF+SHIWynoDGOnpl6qhpFd6Xsq2tNvh+pkd3twOnwC1ecGQCD/ibKYwLM
nH8AQERDZ/pP3bj1+hfk3sqxPtyj2yX3LNcP23snqjgvPmxGFwwDeEXUGiZUZ9Uc
BgJ5haT9zOgpb2SVdwRyUWNwlAtJ+o1zv+30IU5NImAYKzHsRMWwQhUzQ5U3/ppq
ujqRBaywhHohusLoQrKcwLdYQuca+KrLJtCq8WLwTfw1pBwIC9TC/Q0UtoKFigLP
Kbd+MfppuJLwD5G6nBY2v4ZlHhbSgjeXDdJTO+CjnCfX2dYrZgbIt2UALZAF2R32
1RoGUSNHUBFMEP8VKuTzHSFE0ozBReBaj4atWH93OujO4Xzn8XCc9HMtPUL23vyP
hitx98rusjOKz1Nd8xkzRTCdsDhX49/l/RUpl45Ty386x6M987s7MwjLkyP/7sv6
XGi8vkp4W8m7591bgyhbtef/sVDNiyNQFoEZ2FibIqdvLSi8EyH0D3rUavIwAOyT
uaXFnLg2XCPsqZIGZNiv1x0SGXKbpzDdR07sLn88kYuLkcaQtpiO+BmHxb+5XCsW
zPlB+Dxo9viaO2jPc8LSk6gw3RMkQoqmvWK0vJhLCWWCMo9RnKiElgYk+3HJbgS7
ZTwY10SweswVh03asivANGbkYMwiutTXPZQ7SabpJL+cIXtYHaPz8eCJ89WiNN+/
Fq1Yphv+cDj+asgs45t1G4+qJxrDF7QV8I4H+cVSF9bDCnF7m2cOtqkjnxG74Tju
n0YXj2VzcaztGB0ZpPRtscpITtlrpWHF7eVarQsN7cwLF5ERheFxJj6dMSVBR+wK
FwuYv7dC660yRY2L7T2WSNzPEaEurvKonANCgHyyj3DVkYH2W6LIyZ9f7muhzX5k
5VIf+f+P6JIFAcx6P+soIOyqp34Qjg9e74Gaike0o7sg4VZxXwxS5f13CF8UzICJ
wXq70fYaooXKbnkaiXN8HrIc3JvGOwayuTckXNCVPhcjmw9XIMMc53mjHZpu7Sck
Prn7GrqxadIjAAGfnJq9v7gh8fPVxlMooau+EbUi92CgqsFZ9yCMSEUgCpuVBdBs
uRVuJs+akgTvhF2O11pJB44iCD7uzSmr9P0sXREXvQ9YgJYyfn8pJI86mgpBK7qE
cTYcHe5aQ00RsxRCiSVEE+WrTmTYjnZRyBj7mC7vMVZLy2qNdAgVhWwutlZVXoPf
oXb1HyariI2ogEaLPPgUMlYDOa2xiEjZTkvZOdBF8L1ewFC2iItRTNdVIu+kN3Wm
MWFKbVkiuuJpu9KkblHd2f8q1I//sxYyii3ZeGJVPWSBKF7XiFjOfYegPid1wENA
AVNkUo9OA/fWZMdvKLruqFn6P6uaI9MVxr8vd1f+yFuoGdYjEsZaPQabnkrwTtZQ
xS2uy2aXXSJ570OYIvlc7rKKLN8NrLjaTWZ9uDkkukiGPOgvjzcjXBqJ6/o6G49/
7IYrT0YTzZEs3JYEhrXomoxHSHPZHntbO2elLvl+UQGVmMSWQZsSfheAyXhsmLIW
Z2spRMOhICdbSx/jDdCNnD57T6+cltMYSMNvKiL8RMxJeufsDVm+YyahMgRkU7pb
dpekp26VzgeuVa4b2GlrR7bBbUcqpnlOcAb/AzGbLlC/vGW/Nh99/olhXJ08Pp0O
SU7udd6Q9wlIIlBRXwD2bLK5fD0XcpluUpaZMAAysDMtNKfAEhX0G5YCg0MoFdlg
aW4WtRE4nKE7fHaGaDiMXMUNqdv63TB+ghBLbR8WEjYe7n8pYi4lbMuNRS66kO01
5/ceX1ewCdycTNa7z3JHq7EQVbVH6Jj7CoPHLDxpAG5m9EchlkFts8VnheKMOh2x
HNIWu8yKCGZNT16hZfRecy6ZWTMjh6PztZLJIrY6cgb9xVv5r0jEBiswVO+3zhlr
VY0+eXctbwILgdhzp2HlXxSkSFBK8RZkFpZB7dh93ZbJkGBl6p7jJQjr3m2ZK+w9
2qgobFwNjV1gaf+XHPPKkeDpyFBEXRrEe8pxROjm8/fzA1IUstXruhFRDfU+7fh4
kNFRrPHLSIDHe8jBl3XhiZNVF9Ssn/bi/4fqm2zF6HI5iS/ZVmwo6uu45tbCC+af
IIzO/wvTxMz6aINKEAdxmrc+T9uvxDYlq3voCS1C3Urmpih2JmvjQu5FMmOnXbuo
RhLyt36Kaa5/6tU9DzKNZ4JSN9e1giJgzFUp1wz1MEFXWXvGQKlb5aeMjsHy/gLL
QpIQYIPleBglNXCIOw2r0dDYkIb6QLAi5J4OcKHzh/CSTH5IVVuzTHjv7VjFZuKZ
13fBftLrGVBXIHrf9PYea/iY7/ptYnY7HxK7x0QjEA/Puq4u89hTFL7dq5kvySU2
U5CSqRut3Ellm0acqfbQkAdNTpEH3Elyr1cv0Al01PYtcVgU6gjHP1ZMNjaIQPxV
ADaP9g9wiPHSoA9g9QoLBoTJPaSxSV3xGJH/uI/STfa6poNfti350hZGeyf1htTk
7xRpAmb1lnkbJvR/xkDqpeoQ3yimMuzIGnohK61Ihx+wBKAD84d6thJmGR3ElRW8
hpJuuuPGKZ3sj/x/iFK0GKa84W5b6p0VKdRlQnQbAYgfr4084Ei7X8j37yEi5FZk
UZ7XdBOkety1uwGlp5dBDcgArJZCYtwc+AbW5WmZ/uz3KDLCow6NwF9BAtMlXAGj
JbjojcdLIRqSpnJxG+GIEMhKL6LLhNMh181nFNdCF4ume6kJTNGQ44JePe2rn+hf
1u0sXDruRC4gKCi6FFkEG/pDcDEqZwunB43br+RlNj04E85tvBwStVvuIUdP62l0
VaYYjPjAOi3AEQcuTe0ZEl7U7eRWk8auj9rNTQvpx7LILt1Ts5pd62YnZQvWSqni
N7g8VhqpqDAl6Gx8rlEirshs5nfHHvIfR/sDlcFiIZuKZLsxHsCiekAsWjrthLo0
WOFIJolMVKmuc1K74lDJ6hEE1LafZo118sI0fvOGRdk5+2G3tpvfSoQMKE3RP3h1
i3r5QNnjHGhD2dak05pr3YK0exISP8J6WgtRL8plFSEkaOV0cQRiVQ2WEW275KpR
aiAqTfHmpDnKrGhWoLR/06kAlly7TQkaeAJzGx66Pf9sNsaL3/Qg5lzLkt83oDIn
PU0wVnxCZJmJoIx3GynkSw1APrlrxMMJxjTSh9BpETYzdGEx3Raezau7zFnIRwZs
uzsBGiVSSII3tMfJAApeJJ8yxh/lHBlR0ZQ4qUjAr1UuwPZAU1/XadiKs+SOUHqO
GulrVhFf4HuOLqFQBT8kB2PhhfjaHnTc12HoOE2bm0dZ78yhPVIA2hx2/EjFZd7a
BbE2uhPOw33eqcQx5JaL3evgzKypPoA191Bjb+v4fmo0LpfcSL/wqe9E3lyJVgG9
RbtxmqyJyacNN/dQ8u+eNyv8fdGK6TcN5I9LMYxOb/wTiF4IP5e/nkO1xQA0S+1a
3Ksvn5kQkdVrqFioHYCYRldTh9/3jqgnTiYXV94mgkBtF5tQ2KmtPD+NjBg2XNUy
wzZtDqaa+qbQz+oX6d2+TLoCKy51bqwq/XjrCQYOm9eWJLSeoV50sH6VWMTzZ0VB
KXUBc8c2TVXWLpa9jjhWaO3EAQ/Hmio3w1qrpq4nvNRf1lFSEnryJVMl1eJONdLM
QUDeeLv0goEQ4CQC9pM5CJ0BVfss8ukLioLg6v2g23rCZKdm34bz1RCc0Gol6Wlj
topBosHDLVIabln29xHzxCSOudN6ceh8oznwPjkaLGHK00neWblCOj77FfUp3xPU
sFoOfUD8GdWLrYD7jlBb7cc6mxgKV7c1Kx2jOxFKh0K+R3ABZU3kTGPvyHklLGjQ
NOEErIXbbDPCsz9RviXhyjEiWO13i5EDiGy0AW0V1QTKVx8F6SgK6rI50nyHEbuh
ei9v61k7Mp8GARQXyxFYr/XC0EqTrCZD2pOrvZ4f2zvK7fXiUNvDvRK5MeSOLUwZ
kNKsO9YIGed4ReeAIpAKWl+slMXd9hYDvJLbPs8O0V7F215rJvGrdAHhZwW5f70S
njFHX/g7JWqFRoLhex8ONKxT3R4dg7DUPJ7/gVvW6ucOvr9tBrYNsKRcIoaehTdK
KjxVZAUUyOd6rfLXHXTjnkZkt4IC3TklrSMb961Ch3zVMAhy0b5h4xQB2palGuGP
pFwXlGZUNgLukwkcsj99XiTfVa63rJb6FIGg3z937jeBNSX/k361XfG2FFU1qmJ/
SMtioPrye+QLvx4vvgitwJPunZDBtoDNIrJn55KqART/sJACytOS8cLYWN4KoAiI
B3WQu+W5tYB7TJ26Ydgk/wNNzk6i7HjuFYGkGq0rVX4G3d1QyeCkIsCTk+dwFOh3
3Eckd9UdU2ZnV20SaI7i0kjXM06siY1h/+b8skwXwj7emOZhniYUatWkKdpAGYQf
SQdwZOH5NRO1zJeooEZMEHsHTaR5F1FBg6ZOh3hG7rwImKGtNyBsPbuYQieK5tpT
zLPYxl+ZXeNBUGC2AqW1Y0Ry+YB2wzjCej8tiDsl9y+Rn2Eek2o9RaqGAHV5YBv/
oP7PbH17EUAdmA5EL78CFUNZ3R0g8SltKHcmWOQTzrek+uiHW76cl7Y8kusp2RDH
+rRJGCUW9JUUBJGodIFqHK65Voxh59EZp20ikzzw69bIKM2+myuupjseVyaBxf/P
BXJmdkb9wvSJ2otfr8OManIAsXwVzZZDozDKXn29a3Y31l74CKoZWWH/0x+/WfES
TyuKtB91kKgwwS8Dp6pLhpdO9QPH/Lcg+AlpUsBbtFP3QX1YAqJv5DpQQBQcHtTL
WPNnRyjqwoyj8u5kW3J3qYA7dSlqb9/QD6hBipQnhBaSt3JPD+vUwgP1Afz9L/6c
i8OnHBjgQC/1YUAOqLsHYoFneNdPwnraDdvJ0SnXmtSxEr0/LnOrAroFGrWO9Z/o
aG9NzbonGVSB7PhMjnEQSes63OPI7EM+4TH3yQFF6jfKt/gFzmC1pRyHlVebroxz
i35X03YcQWq8yPgI1a/qBK0b+yzm5sozhakyCr1pYKfGxd+7+zQDlnT5ySbNzR5d
rw0ZDLuCfnwibWmd+Em5OV9G1+MSKz7w0NbrOf7iJmZx4rDJXuP0VQP7qbfSAIuh
q/o1f0LqT7OpDObw0M8fWyQRaaXE14zjaREqYpLeQkD/+nnz0Tsc/3kMq4gK/D5c
RkHPVRSjNxHnNLatcCuE6wX2E7OYxwm91uGNl9d9GDTtTHxbQUnQc1FSt2v4yOq2
hHZUNEWTpT3N04PP3MDCrK0Fpu0U5FzYROUsXYQvUghsZL6uBl0AIZdqZ+JUHOy8
/YGxZZSEue992Dh5QB1GINlLmlO26Wk/gFH//Qcs1PEu7xwyS7CNrpOB0Ov6YxjP
Uuyi4f48NEWkN/VQOlvrQ35wpYPvaXMhtyUEC5R8obVo94dkhTVgyeZwKhoclOt3
wUEJBCc1GUhzaScBYEjtvqcakvRpgVsae0L60Jm/rXgWyTmmeb1fRPvx2lpcY4az
02dZeIolLQwTmUTbPeV0ZySMEx8eR+Jpv6bYaxFSTATqK3f/lBa0/Zmdu9TLEa6P
O8EKL3RClQgbJ8o7+OlvSFQu5Wx67mrVxjZT5UcZ4lW96iBdWXqYXi0spP2waMQz
juKIfpZX9O6zURkNQi04+DcJWpR86L66XXbxDGIYxjPLAKX5QxDhejNixUAjcfb+
YylCIPm3B+KzxSU0UaKdEIBCvlXhscP4dh39JVbOIBcJX+xPXx2X/f4re/mkh3kh
7SXck6Bw16rWZR2sir9ljo/FTKKumJtxbglprsmmywd/E811LVOZr0Pj6jjj3vYU
qe6IIAaYpu+eKpWf7o4bpcou69XiNquHkKYhY2tQYlzzk7AR8MVql8GK5JJMuGro
EizAC5tvIV7jWBqfhvohQe0uZ4K1BJSUNRppPSEdaXbdb0tOBcF+vaRsuC/lD6mJ
rJo7QaLdbyclx0ZCA3U+wQ6uTZ/1kSaQX0tjxCQBEu5nKkjN080C2A/3S27LjOVs
SJGxjDOUiNexhfPFpwYBJ1/tN+AKm6w/MEgSFhZuMhP2Oprf7gzvFMxZH6BuYRrg
G2FHMNW7mKzmJgVr6MTmi7RW9vvY8oO0J3bfoo9i+FdUmPAmRjxrRwC2QpBV3Uj8
UFk4pEY4RbxqRiijAiRhGTM/qIEr3XxGATivj9Zs3ZgIVKQJIWej/Pha1CQMXnhL
xf+g4mTm8d/HHkUcxHwHpqiLt5aMi4yLMIGka6hV9CTzOIdD05TYNPv5FtocZtaP
YTYV/K9KRw37aPD7acNi1tYDE44tTMdrbWFZa2MxSZDymTgU52IDB59xZu+LcifI
HNtFFK+WOkDUy/YUokYvs7NBVpXmiHDQSSTxhmQkClbBBLuwq7JCygXi6IbpoILk
NqoDp6yuPRofTzvDUjQbvczFJCq9sfkw9pya/4B/kHS5uqVohqsoAdU/ZCJn+rlL
px8Ee+H6HNakfw1tRaKQ1GlyN4sIpZuzdVff9LBxyr/ap/yUeU+xXq1gggWuPjlx
PyOw64U1ii8Q2CO7gJVn/i5RHaS8qwT5hi/bQPEdjCKJHAKYpoZCwtTAE3zjXQ7A
CEcCWVAoH6aUiAJNN1dxZiKhB4VAH4gesAF8YOg1IXJ27LMlm6zm0sep5ruZZ+Y6
wzX2dMJqI8e6uljhcZjTasJeM9/eZ58AahpNY9+GpBe45+s3AM6knl8kkLTi9MC5
gY+Fc+YZ2idqfHUNXXbAmfI5PQXjfY1z+vtRXqfvvPvbhceWyBGuFrRD1rs5pnvg
tap7h6wYTuLhOvM3f0S4nH2iESzrID0ZGdqmgRB3+u3ugY3+FnCZYzU1qbcySIFz
B3VXRscoWMNp/nPtSMLExrw1GgKFNp4rg3UJWVbubz+YyphBFE4jN+ne020skPE3
phBn4WrQPkQ37wQ28706QX97zHk5dYuUD5YfXczBoafhD2+4b8o+rYeiRz9da5iP
qJuKz3YAfOiLKijoDMh3m4s9uK8xdtwTFLtnlbBpIlM23IbsZFsguhJyRNnIvyrP
DB03C9xdfKrIZ6HJTTqmOWPOc1l0cKy3PyJRWi6e8cZqHRZpzEHIG8NeWciaffrd
qem6ec9JHKeetSxIZhk1nIs1rCcab9If3waEeaGgfc/ypXGl6NIjVmDcdpBYqwie
N3sBsMc/Y7Cw/UB3M/kMAS7KdhGWVwSHnSpBAsdMxP9vl8syyri8d2VLkcKey0ig
20lwfYQtbXD5m8gZfXEpQ/yoga/kXImPEa7gDeiJjhBle48GCM4+6h+qzknT50sb
E9Yt32ONlzINsJwuA/fdxHOuHp5WeQ5zpa4HTi0Y+htPxe8D8dHSK6vf0ZVMyKLJ
sp4lRPBf+Wcr3X0rEG3nIpJDson3VvF0mvq+f4WJNoP4GaB4TWoK4EPqXd0ze+of
hXa6OHRLgBxKZjwgj/SN4z3J1q7LXRnOW0AEdP01lGVdl9P3M91bJD9Lx5gouCeL
6Et3NE49wqa5yKpgtDAJxOfagHLy0TveatbqKuHzKxBv5u59EtKFTWOcb94TaWXG
yOr2ZXS6ZEsyvtUiRPJ5nkMBjbG3yAUde7pnLkdfHoZDlbrUFsKcDLxo5/dlfsMj
vGDf+9JAgZ/yFCuib0DNTCh3+6s9iKgAzFOhExNE2jbwh9JeUDkLwQyedX7qewi/
Y2L2OPyldD9FfJdf80V/RAfIOKhMxwizOTHBC5VzKH6GyIuU23xlPK90C8oR/kDk
IKhchxgsnfS3Rwz9Bvvgw8XC+7+4fXtglxTcB5kyaKQdM6AL3CDVPpbxAEzDJcbT
2JOzdiXbk5mmXO6GjjyYNkzlf+ASSfJSMBhHc6iLLmORp5KFSSgT9R7B6RviioPh
tlzGqE4jA4FYEwEC9cbztBpq64pHBk4nnvtIbNx4mE0YQW3RlSzxutZ1iIVy6yps
Qw6DZMjr0iOUSNHJVr5EvOZnC2qBSCWzKgHzy+jnXRpZ/8Sj4CsdXR7P4lSxRq5d
ox/HjaUcVQu9qlHGtwKNAmuFurqa8vDKDX5P/yIdZKkZ+B8Fo+bOdhzG+iqb+wQy
GNKDGLxDqO2aqRulglyw7wi6QZU5Xfmj9qPW5CY0t9vlKfbF4vsuU27hlPJfrcUd
I+jeDn4dCCMtsr7cotTGXGpzv1q/c4i1mMYLPRSWwGNsLuGiLCt1x2ATyI8KvFvw
IUqfzB+03pNREcClNQbodhaE4VUt57noJPjyx6gg96nnJySLIrjR8wWeeUyRgg1N
ZsQ4uqjygFeke8oX2X5TV0Cd3ZDLrILThIwl3ek68RBOvYhsvTQdBazoSfXRYxh7
1xCUUBfSWZ6GLM9fLbdmGBj+icQNyuTfW4m8Bi6mX3WX0uIiAbGZ4jxNS+kxLUWu
p+S4CvSPPS7q3Kfncl0FMwU/YcPhggbTBlB/Wiu8elTvEMr3mI8TO0v0WXnW+Q21
mKOWlM4KvQ0ix9HWSr0YtdyClJFoCuCRzUUJv5pDEEhOeGRDIjEn+aN0CURsNM/5
01bMR+VAkn3fGdpw1QksNyEMIHUsABzaVRzsAZiYW24Cx14fjlEmdH9Tm7TtINK4
ZdD6FQYRZjRXA5Zps2687Mqq1f+dj8UsevcR0KcR5O9lGUIPh2Y4sgpXr99k6P/E
oc6d5AcDt7svpWUobQ3iuMM6yLGh6XMongjKZmRZS2IoX6NYygcU82U6Jxh6Mgoz
ltFFtjmw8/YbD5fYckzJwqIL0Xz8q3R+6mDOZTgFCuuHaE7yFuSh6MIKOtQzqCIB
cOCnIIJ1eWh/i5CCMoBeIdghaKkPLP9BJb0TqLUGr1Zhu0BiRguCYV2CY9DhQ9PL
350OvOWIg3k5AeHInTTVO1mYLe2HiAChYQrTIM5pVT7dspLLmSJAfZvP4AUrgkut
iKwyzl/wHxGSE3wL7SkYhl4rUzssR5m8n0AVFnXCQ13nCUbH/oAcbBGLrW+ABLJV
TsleVGwzJUYDHr0MJltBIllyv09LUmYJEoR7NFGdpG+zkeSRpWz7smhUh2FgQhat
NQTgioW7yc9p0Xl0kiuEm/4KUOFLbO3P/MtUjBi6DDPo32R4WwZoJwTP6s+85k0W
3qj5BUueSr2cr/2otPw1/bORGkTQz/zTaVzwR5T3yNKH+PMBH30Ns5rVIe7lgGNJ
xUkD3kR7AeiT17KmorljRYZB7llJM3N/7ROL53g7Kl/UlUhk9UH2RZ0780tfiEK+
vm3TBvzuKL62Fnw5c6jjhbTO1V/XRAJisRyjptqoOi025bUbBlsTpWBvOTTuo/da
ZFtphB2gZYDVfamqPw3g6dM7Ayqoa7GNysztdI++A99LJwgnm0938V44Jd+U68lF
KhuC84mL36D/3Ns5U04zqqa+lKEtMBBCNC05xTzBmd/3xu7EJIWHkteT2rCRh8/K
b+xb1qjms/cSY1gWeQ2YBlLi725jBmBzOVAyORJ6J7vgtr7fgxV3DSEyFvJATtcG
4KkN99yToNwrBCvFd/Ec5HNPC5A3WEWVm2KmGASppqO89qUMlTgoKuQyK4OYBHLs
0MjDPwdggWMhXo8ADOsqzuqCZefSNyixdW+Hy39XBdNMbiMqxfTC6Di40NbWcMTj
4BaD+cgksTxQ5JCj6I8zmufEPLHvG2uZQwm6MBFcCLl0/4Ttai9nqmc9pPyHZl8a
xwwYcfGehwF9lBn7ByGHwCDHWOs2/ABTtBcELV1ZAVC0E28+yEqluf9w59Uvt+Vm
2VS9UF4VwUkRvc76aDGcvHcWKJr2HZh2ZSI9ujAUt3PSwxif9AU6PcMaDcp4Y48b
JPvFao2ATKif7eIu7wQtROoWOrODoNiB10zZvJ33ZK6OgHv/L36xWHjgK2ADV9/w
iOWQ4Jnbs6UJ/biNTeEb7XW1J//EL5M/pixOXudBtTh/7Xn2odOyp/Y1YQGipDBs
te8qXX7Wt/cEPHvuujD3GI0A2nc7U1N4FwEnGD7itGgJfCi6Hl0KijrnS33IRsCL
/klW3uzd1pCWT4n8TepBvBzKeTfAqa1UEVR/t5KiFOHYnkvg/KtXHdrZcFNfz8LY
XWvwGjECyBeVEXBO/5SGikONsItA8pHNYJeDtbC9FW3HGLCbeJG+Ee0p5EoDoaDe
1Os/DgmrHp4docGqdIs6KStIbqcG+PZLn1oVJvcfBayUCC/7DeQu26Xj7+qXoESF
XdS7WFOQFFFI8kNUkgx1rAcXh+vHeY5+V+1vzsSufZdc62rFGn5mGmTYJVQUm+FL
L/xeiP7b8rxgNyafpF6r/b9YfxYz/Js6etVP8RenWCm24XmHqehc58UCF7nNJmdP
Cvop7kM2yFZCTpxnENaU3BCk9/aVo/+N7CWnn8u1VHjtfoRgusRfneAqjliSxRuN
BWjfcmzSkNeTwqrXPzbgbXbcrLU8prGvMWp01h7o6Bp4aEiX421i38PB75paWYNO
v3kQrIhIpe2RkaAC3pysM1mqDpeXCSC/AhEb5HovAEtYOSsjL6uvUd4SkCvbfJQI
7GJPlNxrvu2cNlV6P7aEvgkhUqa9/G2o0/+TPmprEHFsvYSbnRZrOmPZG1pUS64B
Z5XCHD8QOcDWfbXsHx8d/XCQ+b+aKArhtQuJx9gA2HQ0ureBUEWyBZ3d83agshVe
ZTVENc6/pZI2644EobxlbeVXoIsO7g3Dn7wYiMO9fZHpUmGMqeq2eRQ3pS03ub9C
MuPvb2QbhtjFnjr0jbLQpIkykDMvONWfufyj0J8i1HYkAybEiHosgSt9FV4E3g5v
wPEubdq29GdagheYDCIIn4M2SpfQeq08uXR0X6IsBhMR7zm5vzRcEcVj+ZNvyGnL
IrZylRiKLMU4HezxjzHGqfmgSxvVuANILzqoQrAoQgTY9aC7tDZoL2zrY81dvkk2
dB2Nhmpfo9PDU/u89oO4efb4NGCeXbBCEj8R6m0tN8TQqFjFVI9lXOT9akqDHGJn
VBqYJ3hekSGipI1LQd3eve/vLRCtU851Szgi7CUDb6Hf0ND1miYoNOLtdSGdQo7X
FPL7KjRyFCB21IXPH8pwdeBt3Zkly8y5Mpk31Zxgg5jJA7sZAvEuEcniRSwD53XO
u538docMVTeSCsPr06ZPvY/GDoC5A4rXcWe7BeG7NtPJSi6F2w49IXgnAnsTl1ny
K0dOcSFu64ZK4wAsabomHIcoBlJP3Rk24p4rDALwRrq30+gY4ZnbRYvITh+MHOKX
0s+Eq7cCcpH9JwGdpmTiBZyVaOGulve6xU0sSy70d4DtKVEStsQGPj2MgEhasPif
aznfPUqoKXzGLXrE48lGBbPpaijlBUxEwKS1k0LNo13Ms9Jd+N6ch3AzbyWEaltu
tR4xKBRK8jNXJvurUMTPS20bcXzBjMwXNl/kGcT68pouyMknNiJduKU2hP2yrxGF
DP940Jp7zYxYx1vnhQOQibs9GlNwOZ3cCqloS7d4orElcbhHsKiaqUlkAf9pn2Na
KlvK9X/alJHl1l8Hrq15C9nEWFCjYLkRAhMh8GHjAUJvyNBXud47ZJvtqqvB1jgl
sE/EKOiWtY/d9h5jm8v5slhElz3TOIpqRvqg59RZNwNPYR5MQKLKUkq8i4TIzEWL
Bf4/5PTGgBmk2uoSW3TaageEi/ZSe/8sBg2JlVUlRKEUEoOpp+uPiXJ8pCyrNpE+
J+g/BCX+PeB79xB0YPf5GBbSJiXHWQTbeUzPXr7YnLxitlnir0uEjgYL10ysjuZt
6LpBtnJ4CGMonJw+YT8AynGT6Z4bnpg7g4qdPqT1bg0nfBcSMABJqrQ3yfDnKaBZ
N/wq36lhEJt3AQ3MHb3IyVFzO7EPvg/jkukm4Y2WOVKsjDQ0JYJlJDIbAUmsl1KQ
ZafgkrDbC89fJXwFLS/efg==
`pragma protect end_protected
