// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:31:31 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
pr3MNCquv3cq1T9tDRygIcqWlk+bmBLB3TTHh4qqSeiBuUR5CfpX06UaJ43eM77d
PVecfOfAs7F5qDf4wYUvWulOLt70bUdQ2c9I1+oN1Tyh/UEMzdDmSuAH+Iw5FP8D
oKqLKmDGlu2v+GKh4aXWX8vhJCjkH0LY7feGtl3NOvQ=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 85952)
9Dv20NAj1vHjtek/mSWn4yp8Z7gymaN1VyD/3tsttqGOVVTM6H2bm7JqEhiX6m9u
9NW57YleEXcSib+unHBlnQlfH5gRzdZJUfYaD4IJC4y8/C4U3DkIm4aPAF5JcLA+
8yio1mYoJaKKtGUVqqBh4mUtQSIr6krcALrMsMQlQXiSdKEOrkSLO3KSs3wvdRhu
mrqPVwNSswoA1TlATbgRnoJnTaL4prseAW5haZF7AZZoAmXxBBKC0FJaiOy6fM8O
wnRTgfHkxKGsjnVG5Ciy5pvdJRs22AHaFRqiIwWhlX3dJVeFKF11RFkVJsys6fAN
/rRVFHiOWehSAcgU6pKqHl04LbhDwI6THIxzq0VOSvtC8gZxzolib5GBkMzJ6OgO
EHER70YzWDBFJOrTlA66rXIV7xOKZud+xmbCVCf4y54QgmQncvA286jyRMpf88bb
N3IMWHJgNeMq3lP8JDqah3pEuilq7Gn7jBWXRXfHHN3tMA7/wN5tDCrDpNiAr7D4
AkNq1H8sMXMpmkHfeNWieESQzgoqUMmPOZyA6l/5fTyVu5rCKtmgzhBAHU4nxDJ1
8yPo7IMODXlkL6gh0B7N+NChZzanVwOaBKUx+oJukOus3WxZTK4SWWoujtjzyecZ
KTxpFSblOScYC6+CysQXdJYYrTORxQFjy/zEgUVNzwkeEdwiTyJz2aHepQO9OYUS
VHpXk3Jpm+yakdvV/EAC2x5+iBfuKKS0iyP3DTtulQTMTPsEI4tet0Xv21rCSyIC
c8GpQqZoiKp72kXNy5BtzwJOXuJby/2wIzbc5Dphk+tmOaSOwF88ndWfn2Nveyvz
E+Jk8I5Kn4E4k/pdjseuT/QxnoqO6PRCSEvtJTUazLOWrQO3zZev4vc9qajY92Z9
GlnR6Q+1fVLG2YaFYKAi93N1VUNXDIUz9jKEjkZpr2ZOKyCBDatA0dlraq5GPIvZ
RzcJCui4Fwlo/l01QXWOWoK2en7qyXwqhHocwx70MO/YY7Ci3UImgXHYdHzOCZSQ
MJ3ySEha/tzWBUbMZn9r/aFb/qPgraVnWXNnoI0V8gUVvVdUNfRGtqLfpJG/l8rp
bgCD+Vv9V80JpYMj/RUH0Zfm6cOkS0GjWfLdEniqBItjQGk92VAiQb7BM1WjF3Nu
ocuFdAgbWFfQqHHDaaH882vCH4X0KSSJcmGFUGDbcXE+Jym5DcwX/K6BQZhDJy9P
SfRmRm3v4+kGohsTzeiim+htg9e1EfFq1m6+HJ6zexnMiJzRRuIZVUge0SmIjSCh
tQOQHlRajgOzB72ea2wriRj8gftedOHIw9ehK71I3sYBBOHVBDCLo+Z/Ag5BvKJU
4nzbhODgeLbRm4RQN6fN8QoQNepYCPdCUNpcn7Y3o8thmXRqJ0yNtJ9yNRjAWKIj
8l0GIldnvGfPkNBBdXPjgTB9WVRTTHknYORCVFsAEsGjP+YoQC8G+Tg1pmS5PC25
9Y4B+9jaxfj0W3wL6zCvHGd/9nXJDs+VW3IrsNa8rU42Rog21TOHF21vQKpeEmGj
xTJinoRLsx7NPzwiWx/1O0q7NXntaOhekP/CqRp/k1AF8DLHQ1LfOGbqm2uLfryR
QYnzAKcraRED792alFJFLowM9KNhQ1VTGBiiN1p2OPSZpEei4JNY2vpvD5U225fm
eUWeCH5KLZGARKrCrOBrVVGiWD5rfQGKeXJC44hrMcBHso1I+/gGbJxJzZmKt/rI
fI94E/0pmNZQAlnB5kIxGZR4zvC6kl6i7lqyakMgUlIUk37fe6Th5S3aKvuFfFf+
PyawH3LAU1WD1KyHqoSBVezvkhlfERs0fXeo93yWXeB2pVmIlWN3acvAwxdCcDy0
sMz/GcrRl+Xa8ZiDcLk6MvCx2zRKs9J+flxCnWWlTp6lEkAIijJ8N51bzyMZjpIz
kCAcvLDy1PjS6jehXNwgOKCccaqWVQlurI0abV1L8ry8pBCnxdGetfZ5TxbZzJYV
TChV+H4mM5NJRS/Kyh3x3etyoWGno+ntcNQ4jAIrKrlW0Racrr6Noc6g4d+bk9vy
8rOtBwMxxLEQY9n5GpmqzFI5IJSEN4Eixdu93J6Hpr4bxMMIMUYfgZID1MlTk4Gw
BlDmF7ZrASi0JoEmuha8P3lhmeUTJsdmJA6VlgsM/uJb/sfA2nu70qETU2DxIf6+
aOcgCPL81OGIPIxPPssssQPR2OpIX/BjtOh9oU3NEc63H6uvzGX7Wj3gBfY1CIJW
drH6rFbX95uufy1SMOYqLJqCCM6YqpfVcHk1B4QZbOwKNGX5aTOgEBAKJMDIu3OR
xnov+lMLt9anLEJx4s/r60fQwblNe98pqETUG2JMFkJ0YddTcF+Je6rRM3sbJkWu
+P7OyHhL2CfhSgpzK3Hyb07uGjB/zvMLnu7+LQhGWEwjz4cjUXxl08JAYksPzYcE
WduS2gOfyDzs0AW1Z2q0LIYmUEZWVDc1bBzXBp8RM5OSrFkuIDcDPyxYpwEovXHv
1cTDdPYeferCnrcSXJxYOJCYxcsYUe9B/Kaw6rIImrXQtdqKkkvFn77rbkSRI2zR
t5nFlZ27rXLf8JUOITUzcJCoOLACczAxWdEF50fBLbWQKQOo1FEN22tfmwtkKYcT
JhsKY7Ner8rZH7WKj6J7+x9xVtoMwecDjFT7bs4uRQWFnyhosSXzNT9PtRDkriRg
GH1R7jej8E1Spr47T8g0+h+gqH8Uf6WtRVV6956p8WW6Pm64ijexcuSYwWR5tNrN
FM4xn9iE0sP5G4D+E5HZo+OmCd3fszYnLk1vloTeigjGlFzEsIUC5ysEb7SIlk0V
oEtTIxZIJ22X6/D9zzR+75yY+BUIyDJdcS59CYYGFLJkuFhQ8hJGf5hc4LywhbH+
qfUFl86kaewtT70kcTZwtJoCWbi+HK3+zZTCNn5nasKGvoneCXgzoLnESJ4SDcb2
JL5wpshRVvkRK2crszNaHvBxv3PplqpAA+sM+wbDxCjYPliBPmmAk/y/p13ayNKg
Bru0dQvOXDOhzxz6SI9mz8vJWijxvJdBhMjfVzq8R5zLAImnuvespG1wPp5l7zoh
lScSeAHIo1vBZgxCgCWXNwK49kCxvNA/7fPYwcOrbvB1AdiIV7MvubMsNdpEL03u
9//APwVB/+NjVVJfToFZ8hURACGje9Pt6TFiF91x88QQnHOvNUg+hbUiI+QKKm3g
aVoDPGPTfN0CWkkKk7+KryXOstBVqwV4uvoTM3vopfSIeMtOjBbRaI/X2p4oWv02
BV8v3P0Uee3xe34lD1R2jSCyXPIPrw9XxTHOatZd49HIywC+MWVLAptgukvU9K3Y
dK6eU8mOlAmkJRhAFspAJV4mCVEW8wmtDxzYdmK4kAG7SnY8WEqjrHTsuS9zXSBr
PZ1EHXcKuodmKYY7SW6SfkyPm+iYtqiNpd5utVYqzcHPFBneq5SQMh2NdGtws2rv
AdIXIgK9f7oRc0SRSDgEMA0QBIWl+3pbr4paiIHHSJE9LvH5FLQZboXWz8dgQ8ez
c9tljtoVe2fMEvFyKyQQ7+m7kHXIA4NtxNsGmBN34aq3APpoiB0ielJB75DYwyR0
6nNvdjA0KRdoiS77zBtEOf0itTOFD4NHriO1/aPJxtl4LTr11CAPEs74pnIvT2Gh
Eo/FJBxTGHPYnIj+8Gh0fckmpTNBMgNWRGes5eakjK4R+88cAmQJ2Dg/rz4eO2zU
DL6+twPhkMvR6NmBJI28gHh3cu+loiGP/68BRLy39iRcftNYbGik/FgUjeu5Ydlq
yXXQpawYsBOF6+7hFyOwh0ruUnv6NesIjZUB2LumKRWQ8W1Ap18gnE44Zs9lF+F8
ZKY9Uv4SsX78KY85Dbw/5Ng8x4rto+k9gE2Z1cJGRFuHHeyqpFZPUwvIr0ilfg40
qLJkPPyOPqUrQ0bYZ5SgRjju1uNX31xuv+yu6r117VUZH+uIOjHcz0YypBjgU+fU
I2Wwtzp6Ri6t/icGVEvb1aAbiPsrlr+Rkla7PwCbCXwxyY/VXTfQ3dloWHALVEmr
bX2w4OEQNdngi8jEGN84lG7kdNl6aKZ5lmTqxi1UC3K3EW6serIefkW/JNT8RrNt
5ktN32C0iAt/kGCest2zQFldtmqp0uWuGvbHgnYQOw9L2KOZGOFW9k4UZs3S2PQU
7psaNHuUrkF/8/hycKlx7soRnCDy3HBw2p1DmIgJI3IMxy8xU15T9gcIA2hue2VW
gC8AAEqqfXkhn7uE+PvwaGdK3bUDX+GXt6qpm7bxdM6pu+3cNGPlLiCuP8SSu7e/
4kPUsehtqfojuvTKgDbzL7RQkDXi+SJ7m5uyPy1vxD7WICxn07AjQFdbcQsMZEFr
eZ1FDzYR4+RtkKd7ZWtELT5DmvKis6w4GFSo0qNq3UiJTjSt+vyj/gK1YbJiZbTJ
C3vQhEBMyYgODZIGroCrI8IkCIHHbxscSku0lL0IE/ARqlfnP15UPsNuok6Q1zJl
+8nBQRIpJaq9wG7NHSZFjhKsieQveIEJAiilij7kA13NuqS73pcZO34ZjSpf0TBg
vTMra+OUNnVp6BuaPT9XRCuCclVFhjsb+IfF1Cu4VV7RR6zghkuVeqbKgmWRNjsV
m98XdmWezgY0XlYpUkODCdtv4PRPwBpXnyeKpsdn2aQY92N0BoxJPqn0YJFR6sqL
Ew5BJP7/xHv4g3hD1sSRLQNFMUAveKL1g5v6vJk7cCn0/0JDaTp3x7WRp84Mycye
I8rvuJkW5TXoQ8dFGFJG57Z5UIRLANrmNu+hctRxVO7dqfcbfuDMXXv2S9wk3bs4
rlioZsgo1Huvg8Bhh/V09w8NwWZFoTUrLKF628RtdGhFqMvKX0sqaTFPr/V+whqI
DYG8TF0VGYlN5sxMxu8fq+Jv+HlXlCI9sbIr+PCwNssYVirh75MBkzpSI5fYQ7cG
1PIDNJObUrE0TdBONZOGJ3C/qX2k+gwsoyjCD/bv1GdfW65Lr/x9/qTyHV5GgnaS
Sv5ktjrXe4KkbUXFHocIjFhmCSaYEWvRUbpbzhTslAt+j5eodhTVay0DVU6Je1s8
cyhlPmUr7NH4tgKiuoBSXYjyCS6GeXivR5QvrIjQIilJzEIxQTYEh/MI/64CFapi
Ks4QW5nK28/jHE0VsFsldFZcZSQGmY0fxkYrV6jEZ1wNzb4vDnORG3WCLeEVoLCB
IHzg9N4UVh7U1BNeHDJE6xDjDc+yje3yfJsmI/40P+Lce45XQpZxeq+suf7ottRu
o542oveb+yGqPOS68Cc3fePcpTtVfX45tWAA4w9LcKrIa7H5W+4+mAa8GByQoV1M
mag65ztJpuK0oPZjcpg9kIlMW/V7k+r37AcSlkvvtwQqEmXcr/vAxyc2SYjp2DbJ
2mZaK8FaPHHc9JD5QNutfOJaierJkjv966ujb8W63e7LzOz4EJD0137x67tlcfLu
TAD712GDHDzvP1pPvBwQjwxyNzPgS9Dtuv+RInHEC6UIVHP1DnFPJn8CRyPX0PCC
8AaKyWKavwvi3p4I0gtnIq/kToIX8h9DFuuvtNInYVT7iqIa7BinSDayAd/iJSRp
JyA1McJPUDhQ6q6cYtEvuHfnAT8ykcQizyb3rvuWpkUaiCcPPrDbujv1FhMeLrL7
AJyD72tpq9O4klQoDO5Jie1reeotFowZDuOWwNCVAoGKFJBTL6fsF03B7cYc2CES
SHknldjuxi9c0EBydsM1r8ZNPFtYyodGFkxdWcwpBAdGcVg3chZW0GJGCeAERcZS
+fx25fDeMFx2pa+byvCNNytfCXLRimpCngd+91n+rRkIMt8o24UgDiyQhOoHUUSq
zDNgD44XaqZTA/GuZzRSTL7sLyirRFwUuEln5UU87e4zg9aM9zCX6N8NdHu762lC
XrjGKSn1tJc51kbU0ZXY23kvQoXzUtFKbC+b8h31WTB9Fwpuc9vOzNMuBNTcTk3J
wWMeey0ZixZVpr2o178d/EqeU0BPvElTTDqh4sNxquJRoLUzMkqE9WOMTuyogIN1
yaIC0UBLIai6c2XlC7bLOK6Q1SWvuOjoVa8zbP/UWweqk2QiQdtxRi2LEH7hVVkk
N/mVCuGGhCut9HPZWCJuUB/5FwjYTl6O9Wk+xhuAG6letcX6dsBj2ClBRc+pJI1T
Iyx+rpTc0Wuozk5sPsX3ohElzDgKckTfi10oV7znPmyxuQwVOOUcs0BnyB/hn0aI
LVxoUYFYHyYR1yfSFBiCAXPf9d5Yuz5LqAel2AYiIvQ8vF7f5mcpZS/ePSpxoftW
JPIDKleKPOo/Ztq6ZA6mk/uFtb32HzA8CbCtKU4OwhM/F/e7gw1ub5UmlK06l/CZ
At7SQcDt5jngupRJ2nyHMpb4KLEUymbi5hgt3BhSIlg6FxeeplgKX13L6ZAIoncp
/jdbFEfmgjFydsLNr6imrBW1rjJs2NCLkl+MKbzHIRML2tfcByEMBMmwXNhWZ2Mi
90E1pLYdBF7J4Rv/uBiFgeb897qSr7jMhiEBaKOcKGQc4l1Oemy0X6Hss1Mvjll6
Ecy4tiKwG6olqkzVrW8QgC8a2bL5WJtdPF//C2cx3AXbcvUTHsWdOvyGsonh+FPT
6HZrbJVmRfO0oIqXcQHZFfK6c1whbRtwNX7LtZCTCnxl3H9lOIF42QiTCEGMiEo3
Ex9jbflf/kUSGa+XJjLjDOIYFhxHpAmdcsTpmWyMSy0X/FQw7dLY21FiyejK/H3/
fwlK+UQGflzs/dJDQxYTR6+UTK+C3mqZ7dqh1vQ8SxOguqjhltOpb913XJ2JyxCl
BhSUG2Scy5byzPXyM2d3K2Mv04rEAAshFl4Bqe7z9QB8oQy6lmuw96aUiRgKlcyn
SFhCwbuuV11LYgJB7+R7NRfVZjv9u4IT+7bLbvKSFYXhOcLDCv6oSZJi1EWs0GoV
qVlQfDLHRoDuzy/Qe1A2ueDd7p8kkAbH1OEjXqe7qlKZ+u/MqCMei+Huj3PM8yuh
9+TOybRoGtxK9NbR/4uH+RWXh+KujOXKynKCQ6qsypbMTSrQ/Z5fNYIJIr0NGihy
ZBaJAda8UiARfJWlFXnHR1mA5tKbS2GDEvnqCruRQ6sbwF5s0fnplKJ/hA3pmQaT
KOQsbCiM1k7nKbS2q6YP9CujijI4pz1emAHl/LCHxz6Xlq3Dqe3Y2ZfVNheUNoSH
Wl2caNSM1/a3Gtf4zcFx4SZ2OS93zyyRmO9g0uApo9tUyHh0rUs8pOCDia3eq5i2
V6o57N02sak+10blDN6Wenei82DdKGAwHTyjSEblShqcvhzcVZ+k84jz9Z6gph0X
kZ30Pc83FJn501GcMbIob+LWWtFEx7ybw9f2rThlmiK0S89Ky9N5AtascdiinUEZ
L+Z5EUXYNVfbIUX6KMqSaEKYZZpYQFyRiGG+lBuSLUo3Lo7kUg/RI2vAjhs6mPPo
Exqtux0iqY0CkgyJYn1z2G08Y7qJmLD3+uLs5qRGewrhu/mZx05PkibGVMI1pa4m
Uc+thH9eKkFTACiPv23xz9UDDtBp1J+GKsl0ib23steRruuUrwNkCrf439fp6Kvf
BThIqJyiIVtc4Q90yDfMr+AXqwl9DeWGAbdKgE5TvQ0rhOfyRq8OaTNzBzcM3KyP
0vlqdybT62bSbJOOVQpRX0OUH7iJ5zFeJZJ+j+w0jMnoEx9trzIJg8NJuYKotdod
wDxf42lLc7e2bmjLi4LzP8K2AvwYj8WR5YMuBllZ2CfYOh2x1tCvIk14rxHKjmTy
m20fmhICf45BuejFIWogdH5AbsgoHkxYuYtPNEp/z3Sh0s30GkZ0ECY28PeNhKeh
qrsqGPzr6JgxGYNI/qpATFnPN9WgjEum0h2WNR3GhRh0Xo4U8ao8kUZY1vkUCqht
t2nXyyPxvvSYdX58X+adRu/sEkPnzcc06u37TbIX3nZTM4E5plZPgTdZQ3HotYlW
yxVDBJLflX7DI8ZhODTGtQk+LhosHlNCmcBHns4j/RvF9DpY7jL4fn6EY2KgnWWv
9Gm6eWTzoWGqyVSMzb1KwtHHtecbjbXzOsEJrYa1C2LuuKueX3cK8CulK4DjasyB
5HokkrcAWc8BchaNMdpLr2VytZ53PPl0Ni9XrlRkt0/Lt/dBh2aoOsxHtFOYnPK1
wY6XPVDtlVw5GJYaqXK/rIr7ggIykQBlEXiq7OT8Cjl/MdP8Y21e5xylHxFzBpaz
IbQsqh9oVIZh37zIIAY5Xq9DReG7RC4yJS53ZNX9zAb4q+XL3Io/cOzs8AisVexf
Pz0oGXaAV2yqBiol//PhTSy+oMKvdggpuRvjb5hNRf1McftBYeUWyCDCfyu0kWZ5
GJG77sfbiTSbWxnbvwZia4BJ2znglUp3cw9nSzyfzHYvXW/eIHKesutUy6Rfvce/
ozh0KdZHdHNIL/PcP6oalKhb2sCuf+LMiRxRAwVvKXN52u8PMR29eb4epbGPWcfG
FZigEQT7Jukx4Qn0yZUOOw41lfTbduIYmdRQ+U2uLBFLRszXmW/sj7ISUo5PxoXX
LaRptfKGUkgMU4q6RtNw/i75rOo0ylWvY+B4tJpaQK9QZLVC1H81RTtWgYFLFxJL
NnZTDFNqoPbkpvEYuvs3KNOpDtymWLxu0QAl+ByGvpLgfeuDFG3xPVIIheZ7AQ8N
CJ/1p+y4EJ292zEgJ4gZ8Dv/DsfKfvoR6tsCGfJqdloxaKwh9WIf40hTu/bZ52cq
D7gmWwO2SZovkIn8UWTmmFRSiH49XFeKGgaBvoU1ql68BFo0ImbmjDFVOlJWGWaL
qhNOT8nn0t3TXkDjUOk/XKwPPbp5TSCRkg4Q7eL6hML6EybFf0HI/H6FY4VGbYPd
hYwi82MSptcc1Cw/Ixwy07LrT/MkJO5FUNq/bO+yL8IMkqESnwHnKPfySPBO4lmF
fiZ2F3Xvds9rA4Q2SGvRSsh7s/3EbkfmYHsIHPvbSVkHVEhtaWI/SamyKS75lhbN
WLJydOnHzLopThyrhIBqwlNFwJDJh9QUyQ0BK+QgxPh2HKPbP5QooNXsvWX8f5X+
VAjX8ppkNegdM2IKvl9e/w+qagU0RZ9uZrkXIW5UK1COMXoTjGXuolsC/lMTuJHm
P5WLUa9u345o103YLRRbKPMgx3fSLjOPXe6118D80k6hw6kd4R6N1NG6lBYmEmMX
jUFE25VNGq7t4xRJC/birK29PMzv2fJTTCOr2ZHq1QLaH1sj1UrcI3tqpjHC9TTd
VbzlUYQNScRutISWFUn/yfjRB4yAdo6Ulu/UbNLSMHceb9XfGUOFuGp0h5SzTvMx
jQqxF8rzwQQtNjFP4CgGVHJrJ2klInRCD0r3wXx8y9dUd2HtHsg4ZNmafu739NIF
LKAszmnxYzEUbO+NHQV02HUWPo5jw3x9ZPvQnsSsXsIfum0nkpJn1kbFHD1Komo6
MKU+DKJ5B4QgqKRZyw866Sa5NLejNaBrz6X4FRV0ydKU2NoGVMFXoQf8HrgEuAy2
K3Y917a/Xnu0W/L+6sgyRqvGF/NQvVmrkUfKEalsx1ImHwIan8AzGzOjqkVXRJ3+
1mmeuk4ULiIdx1+EdscsIHoSeZRMMTz48tjnMdw+GU0isqWyJE9I6XA9sRxAffxr
eNIOGnpqRyGIeWUnDQzLQ/UgreRQVDRct3KGW73dOzz8uumKM1yHChi600kFc7MD
Y4d8njO/rGHxNSb4OR2QhUsyoN8pBqrW11Pum0+doMUQafXXnVedH75nP5UNzFA1
5vl02tJ7teI0YgFTN2+wy20WbpVeHXoYdEwgn/rFOCZ17Fim1W3x9dQ7nunlF6nn
5vRQjLkNscgY6eRxglCv0N/RZ+Kt00N8V2R+jahDeUHDOyo4yWCapS6uBPjD2moa
aQunyERrSued4cf6enyggTI2TusMy1680CsfiM1wIdRirFUlCBAEW3HkG9J1N6Sd
cST7RhnartNFm1ln2Lx4b4UqUSSur4yPbmjDeDPGJrEtEY/hnuBBWHSB+EVhwzfL
YAQXyKxEpHuiZl1gghlsO78oSKf69CfsfH54OrIek1czxanulNvi3/jALQ7NPcuk
nqM5m7M5tzmnV+RLI2BeCbFPxfj5BtwEXUpn/TdJwIkk12XdJmSSCMEQwMzMFwP3
21zHLNOb3swOBSrTMCkxUP+oPyPIP5nox9cEfDYK/S5/AULFStelvAcggWSBX2fF
+SsRljO4HnKd+EuliyhK83EEMWl15S3GLcI7nRyUdsT60ulxZ0tTEmpHxTpJ/SA1
gLXS3zZXgZyLF/WYM5PYzdlwDPkP22aP4ZWSP1CyeW9mfO6y8FAv0gbwHGQ/l++b
V4I7zijc2uLYtIGhGcF8eVC7YQJmc18HxVRqeYZ4HVcCYOA5xSipWxseQ7KQz8xu
Zu223R/adYsZLeULI9f3u/RhRpkdjCVaKvacC2aojy03pTUCbYgZgCk7Gg+N/HUh
AZ66I7msLw3CluytxZ3dZoqrGQFDiRgXqcH+1V3WFUaZeoK8VpHPmMGyOqBIqnVN
wZCfQSKNHLO/PWNKsHK99mwd8y1YCOXJ0KqMUPsZ9B6SsKMk4RtdyIc4XTRyAmQV
jEE9niznwoqkvpVbAi7LEG+i6TA4/iSbY+uQp2K+N00/DyvQkRgk0pjAEcas9u8l
ZFFXine469z0fJx0cheInghXeFugEnORLClW9XU3i/OxMk1T0ciSlgZ32D29QSCI
SUXzq1PPhBvSYfrDbB77XB+KC1gVqeArSKBozsP/Oy4G620yuhp9Ozf4y0H5aSjQ
vpDfUtYYXHaoZgIqDtvpX5+Co+mEfWW02ruVqO3SOhyzLtzEsRq5iCqxMLabiAiV
7PQSrlPdRp2icUfjtT8ScoVNVp83uYQgvMnYR1zFDxuliwPUEJYEQrCfnMaLoaK0
ZPAEdo7xfnb5oxq4NFmH4gto8dwSZXJwLe2s93DVGBLxw89pmAqdfK4hQnrlofHI
Z4UprTLHmUAX1jRcJTE6UPHtpoLYKQFlAwkUiGjZ9oGtWowEQNvyNo4GuYI1YkUY
i5j+MP1KxjqljtDJC3P24l79U1Hv867ydT4GEPGub/niu3eRQtHbj5GOMkmyftDL
d9OQwr75L+CdzcuaYatF6w9rIZkaPF7WqhLxDY7LCQdychh7hIoOTsFvzzkco5JR
500AdLpQOY8yWkBl9pf7B+1UOk93mALiHhrYpKjlgRtT1h61gKJptKdWyfSZ9JJg
IHLUNpazMMf3C6JaA990VC+gmlfds1Gf9manX7pVQhI++lTwZeP97FpDTRaGdTG6
tXzWIYv6DZKmRCfMJqGNeTlO3SMPJgH2+9Ush0cw/ZucplE5Tg/HwlHPdsdgy99G
F6LNFisY2+cks/2yhujJJYCULzo2AC3rZJmk7yqy0/kH8SRR2TPIdJqnHzuxsXSO
N02AjZ46D4Z/yGZPOTjnrcBjSvmrW20+APm39K44rFz5t56blZr+9oPpr3EQ6vZT
8Gq6lBmGG2vacICH7BEgzd6bzw8w4LhDTybWU0ehbAqhLpZnY3gnQbTegwKHYqPL
tgcUUiV74mth+7PQSulepiWhjgap65PQyeoo1QidR8t2QJZSYM/T+rtYt2KkKFsL
WJ3aGqCrPdCH3M0s1V/IJTYlErWxjeVzlE4GM65kCRNaVA1881a1qeldc5RoJlNH
9fUPPvds2Pm45359JUikyS+htzxgKxSAeHfsWcvrf2uYC/cEhjp552X/gYJbSArM
YYMxWgVz10hMqWLLaQsxsm2J+hDQqjA5DZnYPEo9huMpBZXYwZzqUyAHdDCAeqGs
01BmBhrfyeBMqgzzzOu51Z7vjAfwOw6+masXuWiIfIwkJSSfuqulBD9VKabnd4sP
A53UJ+BncEXKyCtMsM43iDKz/dJtxvhuTKEniSbCt/7A6hjUj8tPBRxh+6IoCk47
i7qZH8xlkhqv53VqJHbxAqPP+UAtM0hKLgr8MpA6ts/qcs9Cvlc/natczd+lbFZw
XmSQ6AzjWo4rMCzd2Xx4U++b8XXkT2qNVmKZoO56TpyPzzRm5/L+gTQ8wP82bL3E
hLyEQYxS5OUy2bTaht9+Q0f7SYEnhYZL6u76n/Lm/aKFq23yAK1gGw6xPvkxNQKj
j39/WG1qT/HMHceYQjkMjgXaMvksvP/V1M2PhoeG3ZaGiJfQy2F4u2ly9kmLHPP6
kr2FIk8jakZbStbbEsEfSuhVeNyeFnP+RytMhd5Whd5de6oE1JZ8rcJtUE2Pdpc8
+dFJJWLmbYGUQWTIPfXGdQxMUqbMzrVChr1WgE3HbPpkXLQMBB/Uu+Y1Pfrp/XRg
bj0jeKyQ9Egyr8wtqavQ6Ildbt5Ojoff4xKpLQVsGrZgBIb0cSJU4YYN6aaFGdMm
g5J2Am3hm5SiZRgME7iTx+y5/QkGwiOU03hnjnwekvVU4AdtxtsdX2WZ41F7tkRy
M8hZ0cIdgKgD8uWMxbAA1MEhIEF9IRLGOmUXh+d5HSkgAjLr+W4erDB/jq1v1cuU
xOKWaI+vgqhwPBX6KbypSou2El4boBmQsFHIzdOYpb8LFvLligr1Z4TU4oIFM7yx
ghWc8c74bGdnte7kNODthmG/cZ7XMEUuDeHgV2yxP19Ro8HfXhplUUDymnhcfQP/
gEsmj4xJnOOOrj6GFSEl0+Lw/XgTiPopJjE7nd+ejv0R1Jf5sPkQxZHzwVq5Fj4l
7IU1u6EIOeYOBe70PB62xXTdaFVAqQv0RAvi1Zhk5ndZfazCneaJDpBPjPoOfj0m
ePmEaUo33JPa1kjd+qiYwYCTwyzV2LkfPffw+YWJiGhy+7pXPnGvQTExkz8tIZvE
hPd0ML2rnrn6qoRlU/LT7/G9wA0c2d1dUnnESJS1El+WhVABkozKGznBg0P/MpRA
1NAMRzZnmdM1sSCtULeMFzK2xK7UPTYVXUob/QvjAukUWIIeEXq1AHo6eM6gknEi
L0GFd5hdL0x08JhzZm+03H9UsO6fQ9/2rylBe6n67A8c9xyB7LqDu4fpxERBUClX
6ECkagS6qJmtliSzYSx06GKQI7yS5hrT8JrUk0Z7CmN2IfWrynJII+v7RBnpjpZ1
UWarXff3es0oLEp4+8SQ8ZNU2J9EvHi8imu38CDC5P6JbU57eVTajKiq/ik5aKVt
XROSfdnyaFJ/UAVS/RWHI4ZfVkHBPcD3X6oj2xZzGuBLIoyzikCBaQsyzqwDQLBT
JKR5fN6k/zYw3+EWtbKsf+JDv1Zm9PPqOexDhKH4PxrQJifslrdLAdzSC/N4iLcY
AElMMCvgQhxhbsmK9NBsFMbqFZUDCtD09wSwS9nUNvdfsi0GdgBErrguWcGHQ/a7
NdjyVDNC+AXhZRjMHZMw4fWQCnFSWoayQqhtCcHns+A+hljQEUV/nmnTv8DIf9Ed
oN8xsyJcDgAGutFfnS6+zr53Uo8DVyfQva4BEu/i9FUeFw+01w3EgrRNbFq6XaP1
qkk5t60iWobax7bu0ef2didOiOrf5ZvNvWW+yF9nDrzrhwNfJfNOloD6gy4mvDg9
rO/AEBv+HNhVMoHIRvGCXIla3dAgUtQffJ5MgSH5Z/Rt+YHIYCFIyq2C22NPy0rh
JpY2FnErkIBJS+pilAIB8rD/y5qr4tsnPDN9g/6i2EC0AuGPucI59/+vBo8F6X2Z
UtoTWYMEAusXuuZT+wVAMIBr266kriktfl+TbMq/wobZv/pM9RTWAe4Ps7R2CX6u
NFzM4Rhs6tAbF6Co+iwVzRQeXgrmAXyniV4PsIw9xoC8dkOVvUg37Qa9NneGZCUF
N7A2QaZvkcGaazrYaNz4ljf0/SFnvuFsN71tE6mhlMLqVchPWfa/LcTvKw4kJlyy
K80uuBpaNBLHn2xBlCtXES/WnZ5IHF28T6qPzy9yl8kHyMjadEUjaMjYL5/OpM6h
NixqJwPx+xVqxp96lrcXH5uRCG9haq9t09F5iAflETWC4uDx4Sq1lvu6+6stZLWv
Y3n9hVURTCQNDHbyZU09gYonjvMquDsyV6eabOTw5ZhpRmmcMwnpK0k93FyMSwe+
669WNdWluljAdGJIcDbOBwNfsrhY/kXsVziaPcBi82jqUpntaAhGsnJbHe+81DoS
YlQcvJQhR4hawjpas33j3eRjiPJ+0yfEYWGkeMBIiVxc/TrVlt0dOBl+rx6gxQy2
sZBeo4liDVWGsenhXgmRF4++b5ntUd2XZO83AoZbjD7l8frjDtilM01aV0hz9UU5
gISEQ4PlOoiptHn3FAu41eXYGi9Xp7mOkIl7Y7u2uXgysL1e0Nm+ASlBICatZePY
futXmsWuLkUgwpcU+DbJmh6MI6/CUxRt4ds542q7vPvxprRC7r8YGAZ0Um3A+B5o
jdUiiq+j9SYXyFJGj7fSCGY812fCkgxjUA/ttN6/H5nu7E8HxQriIfxJeEr3SNGy
rlgGUeTeb5Y1KQwVSSMH9Ho/PqsapSQ54ZdE85xAPVbj8bzZhtGyQiqrYRdK0Wql
ouGuMLI+kiqXWpvp/HkImr7rQ+12QEMrmHeT1QjYAcTo/T1XPIcz7dY6YQma3gEQ
dyF2lVQnjhyRsTDktFMQafhSbk0W3zylm+d/R3JSw6kERDF/T8Rm8c7mAO3z1/pw
gEhHwXeD+Xp0ZldP85VNLRGBbTPZure90gZx9p50e9G/RcC0DM/XIgWy3ur0/tcd
Mr1rbFvpnvLubqN+WCtq7sSJ4HyGp48gWUyCdXUTnc46U9r5RV6KZWPiSvrBViPI
DhSWUFljyAE72x4SBH/+Fn8Lp0UKZZi+bhaggcosRnkXjBXDY01N5/sO6fcOFv5a
mTOZQtJJ8E6BxQeZ1rwo9hst0Juvqf5+zslVCTdmlyxzsHVChnBOZbW7Kqi3sMVE
xzmwbl1NnSZXQkGRwFjLSIzKnfUiVxdaPWsHypK4KUXx0BtgUL5KrPGLQDfjGjGp
DJ6Ph/hcMR+AxgqRcGzSv6UZ2AW+MapRiOI0MtIRqb9qfpWeVMaUNR6nXB8vI3Z3
NpJCiI4x6jO4IpQzljxSNegahOA4gQhbcrnrB1uVWsYQjBrBR/A/Hv1eUJUS/M89
r2PFqbCQ2R70k1c3UR/d0TgcrbsHjQN9SenkUR01oyUmWO1pFIfp9gfMleGX1YI1
tm7nNvlB00ULuXSvbRNH3SPeux/2bKjIWc9tOzx5VfeiHqHgy1xnsdgFltxcaS8V
hyxM9bJzmxevPsucIvtlldx3sEU6sutSYz4ASl66YidY7YgrliBT5zSLhsBYLDaR
bXUfBxcgdp8/KQWVrQS+YAlMqbxsqhYAQkLbGgz7Ilb9Bmc4YD3VjLr14mpBzMgx
zt6AAJKDKwyqaZZyEsFHByPDNvpwHg/uZUv6eyknYieYPMxUzC3fdpQgIPIsrfvz
zyZLuVgtlM5ykoLMaWZVtoq0VVIZQwGyP14ABezDIu11tEotsv07ISWg4dg4bF7s
qf312vBMG9BL4+7pbANQ+/WaVzalqh4qgGJlK4GYhLmZmGnwG+cxSU5rxDWzqJ7R
/+L+qThCoy5QBxQRKnTNoDQOHd7aqMJL62/8hWCiIPeynLwXpATQgBzhLOdlJB0E
HsuaoVn735d5drIRmiOjGlyKr/9PIhPKkGiKqcE1hcWMrizRm1+JZWsQ4BT3GFks
MytRxtfhqtOeG5PVPacHsh3NAhdLaXefD+3ob5V8erBG9doXYX06pLec+nNV/l9H
T1gddUhNeF0YSmmx/ghtRaL05zgv3y9YIzyBW1sCN2aFGbiYLjH2ZHgNwePViWRu
BHAifJfiFeGk2efWOrV9jwAZ19Z/NlyZOXI8XNa63LNOloP/NRJzdGKLe367R/UZ
Jug49uCd9hQ8cHiJqZ+nDQWLHIKsWK/ejPr6BfSSi9N8ix+NtaL3Q3WNx3wjrFYw
g+9ZU2eebg778bTp+H8Cfh3FPl5f9lBxQ63IDY1JRy93S3xRtvB1ZJO4ahH2cWnl
/+ScSmhcd1PsM/Xfad4qcmaUh5pXi3q/E3z5E4somF2X9zF7SFKDNugsAhvRcDb+
/hAPuNt3txY0Hl5vU+8y+/Q1gylN64CEts9o2QlgZ604pJaz/j262AsZzM3QtFvi
8orr3dPUob6Mu+TyoHKLUmWpkk0zpj0sl1fKz4JFnMuk3FcO0cONVNkvoIxh1OmA
B0TPHmWVwAahSc+ZxLDBNflYF8UiCR2USjLwcEP6HsHD7sXqv74Y5MUmlqVh18ze
zRrdC0FVXEGAK52xdHIaNgC6Z08CUxFs7cS44x6/KLnA7Ql9EgEyteKB3xGWZvJN
p1XgQgC5IrVrKrzB6Fm3yzOMT4Zb9Ig5DEVGIbJXT4z8hK/ER6wAbzunP0AYMI4z
n+qMd2UGzFHwpiD4uU7xakZmZbwwHr66jpTU0Jejkg4G96F3z5bd0loeCEpuJF0z
oB2LNUZFBw5Ls3tWf0xORB6nVcmKFKK8k5al6YFQ45OBGVeF6LvU6cyUK9mFBPN6
0+wSlDLZ7CtDwwcUQDuJsHWiHqcEf/NbmUTDJrzYdD1LPwy0bb+6N2mEK4oq0NBT
hZmSAPLojkywxWjwvgG29zoC0Kp2hxL1qgmYIY1mtHvEEZgyl1rCajvZ5LZ+4tcZ
Jr9EzFfPZfCvsFufIw5ko7m0QkxiBLMEfVOk8zsWkuTRrKrIMjnNNIIpK5GAraT7
98H2b4eScc1lWRHgCLUL4WZwC/tEiclxbT5BPOVdni9SkdmthQ8rE80Y5idmPVse
biOJKih92igADEIBDZFKz5PuD9IDOmh+eBCWPjmxSENwRh3YF3kCoh3k0VJIB95L
aMx1EPV6+34kb4pR6Hinfi0BD3nE44XETxvsuyIMUkf+mCiSZtzB+VJfN6vME0k4
02PhurT1zf/qaoI+sGXnwzBxUTrTr5G87dfH+Tb4zAkL2k4iIbqkP//QUHrWKUEm
Ju+KZigN5IwAYjB+vht+62hYYSvhbBHduJGxD6D/F9M4GxLP99Reg2dJYFZ6SDaW
QcaoVH+OnGV7LbyMA15SynNQ1baAQgC3t3nF0OU74Hbsmb8gRlKgPkBIYR6ttdbG
U690Iy/10+PijDF6NkriOtOMCwr/MHaka12LOd9LdpywfWEkiwWlV/9HfhamjJ9d
+o3t1xyotGT72G+SNAg/VGdVKETtcezyIptaJgOBNtzcAPpoxJctsyNwJ0cZB2BJ
0do754SUkFRUCf1zbY+WX6vmrOJAoxVjngsEoudJrpqwzcIX2hDxLy3zupoUTD9E
/yzpHOQgTEoG/wCWlZ2ZP+MI8vLYPihsigeZoE2YXdnMWYq+uWegDpCR32JQMLCQ
2NOKbJszltHy3GY4zTpPO0x6NSDCJOHEuYyL07saurwV3eNJIkDAsm2mo5ug3Fo2
Jj7Rmx5dzWxkxRR89T2wdR7J2QLATVNGf8REVgzG+rrr5ThDXnkxutpYXnI2qm/g
XOLbFxsw/7ewcok8oAHlR1Kh+3xmCdDBI8CQDxR0BkT0NU1c2DyF3/gb75vf8Aqx
f5uezmCrmW2C2mKPDWejRTtxUkVmxTuxJgCe/4sRjIkEl+QQRgXBGqjRyk5XX3SW
Yx5kHkw75c0GQt2ZwO+MXWMuQwMeZiXXWiiecv/Ov/DQAgE5aYixd2i/Umz0+TIe
QF/stbl/sNLhrw91IJjxzZOAuitOrIZXk/4UCb8xKzt1Nd0fgKZS5qCcSraZGejQ
BP6l9AJ0UzXPBplbZGHJKPhpJ/eF7KYPkIE5rwVO9Ifh6/qMTP3bwawsFXB0YFSN
07qZTsNGssIZNmyTEEPD7XSRB6xQ/4xQiEaa8Yz6JjsQCeICPDwyEMt2G79VR8bB
SgeP9n9iBnJrUnhS+XaF0P7EwDsQYV9JirnEkaWDzf6Uj1sfdw5u8+jX7ZS76F2Q
9uaiUUZmhT/sZUoSX7pl2vjoEUF+ckNy9sIfJf9R2g/3K67EUFk+HUpkO2/ElftT
zmYKyOJcq70CRoXpi+jW2g7+3Goov/kPP+Wb6lDQ34gGAUL7Ayqd77XJrZk1PtJ/
IBHs8aPv6tUrPe6Bd8hySx5qnHTK3CSO3iYAHE6d1BdAEa894+8B3x2VnlgT91t8
Y37m7Gug8ulesrXOjv2fLQe9V/iSvuMFSx4zr9mLTZLoxKGp+8TxWoLtCEbYdTa5
3on0RYe9sA828gfHOQgjttPF85pLr3RVU/i4GSvW+ZaYacN4Jxy7v7LBQZw/AKS0
Y1mKndrxUQ/cRoFsX6DHKkIQPk1SvK7KISADJqpQFaJ5p3UfZmHpr/hv/dtTu46e
H/17j4unveVfjn86ZY/WyeGIONK9uOqXi0TLKpAwHaP//W7kHsNqt/jCyXNpmcOF
+GXuIkcLyc1xoOWXVtSI9svdCsUY1byC8CzTNmyuJ6Ca2VNxqIxnJKdnVUqYv8fl
UZVS2xgjQUibAU8DMvh3vpzQEVe7BY0CZpUUidvuoKx1E4IIKFzT6Qam2dXoAAc8
LE5L1Zl5icTyieyKHlqFvukl52jksFCDw/5DDAc7MrEkrey4545ijuMCDrRDXrxf
aXlswTNqDIObFNBQIxQPr92Eq6wAdXd4f1YmNOOavIjRxZrbv9GDD20fKWnDBvx6
OL8FLvY/mn9R+fNoi0OUdENTjbx+Tv5KfWGnL/f7DJurOVwhEG9nL6xDztt+SFXX
43X+phn1xpqoj/9inijUhGqB8D5feBgpj6FwCOtkyWeVZenLmxM+W16E9ACleiv8
J96T0xSE7L6ZyJbzzFV7VDlZwy6Cbgv5WURfFCNYyUXxFLvLTxlYCUhBKyZw3hvT
hcJr0E8q6wjjqBwcWEOynURzzCWpjEFNbs4FyIyEOOYG4QjxhFBD5WIUqDAkuw3g
MPNP4QQ1S3JSxNIy8t+fQuqoBBXBQ50la8SAy1mGRCHbXKBDhNzq+yAIkni7+Py/
ZMwKprVIYmF9dK8ah1ZhhfeQvxg45dqrAE1UyH5wPHMiuHAeVl5y7Ay2wcwsqeqU
khTad/lx4XhmpwhmnJYi8de135fyYFoCCjJu2qrFJKLllwG0wAI1SrusKWj7pgtz
V5BT1LRkiAOVnC49RJLFIBGzS/ByyTxBOKIUW6erycaMdPJ/3pT70C8PXgqfdbeO
SxnPAh9JpAjcBujfBRYJpYwpMVQ8SNWuUwXkegngu9Y25ueuhaJHDftLToYWDe40
8SNgUmKKiaY0n2gd4FQlD8KgyBh90+ws8ML744bQJ6q5gypru7bPg+de2d3a8cga
e6Zt0am3JNzVMCMaUlD0IEo5wlJ2oZDj42WYByVvMuJS2YsYm8t6SH1bmw8LNIed
+gXt8aI/HMG1mo9o8Iw+cHOQtlcEsDKNjDx3e6FyOWKU1LZDcGfz/F1VI4ubFOi9
ztPcEsl0m2OGdcLFtfaN49nQIxvlmom4XTrFIylYtPbHCxCaCcZtLHRO12XLNma4
dQ+tt244aWXtgmk+TUK3D3JAoDziBK1psyQyDVpKzbi3YsYfsVxe8yHT++DY9TX/
CrsUFhXzhbjBHlDvNBzn9gNyLCcRwMoUScDhBp2+Qbm6q1sr4WsdfrhX+u9q9VUm
RUWSmeVQysrH7TrQybSvfM/HLSetnIYkeD9sHKF6O1llAt03RCAnYlDUUB8mAgrV
KJ5SleXxCraJOJ5qNiejpQBku2qZU0Hpq7WdEQP85I/vtrB9HpGjr+o6oGN2Q0KD
hjd0xwSqMSJ1NS2+rshu5Dd4WmdIn4Ex21rZb3fVHAXPit7/JenUKl7TMB6yHEgu
8jjfNfHHADg5dMfIL1AhhvJM63FB4aY2RkKlsphmlzD4EuAIqY5zy0M1xTsLvDRA
vzt2Eub7XwLEiCSUdHpjkK19KxBPfkixJHFisg4nNhX021z4ihr1D7/Z8hj+av6w
0G7qOo6VfQiPLjvlZ2pg1iybGHZBD9q2yqA11RAJpcOvtt6tTOPHM3nzRpU9bPBr
fk5hYBnw13OhJY8Fx/lxly+x+Xb2spuHHr7BL8URbN9WrTABVa/heii97Zqs+MdA
xpZGE3hlADiZUXz67SELjqEnUiQpSGz4vZDjLBPjmc4T4FITXomllMh1SXhZSS0p
QYsavHmLVoFd+szMNN/yxmrenrCQvDe9qI6l7GrTtw3t/Yhib/6sEPiGQlOf2s0P
6OJKah5/zcSrqZ9bY+z+e4gJYSY/OTdtdEQGzV+H/E8gHf/ZJHxz2mJhb7KQ2JLS
k2WyWk87fdt05jC9wSWWsiKrm76ptywn5qrt0W/YlAFQmYjC1ZoMOwSLtAk8uraR
bkvI9jVxQIC6SguS+IuL3v95jcpVK9sz4ACFprr074ZK3jB6rfRNaHH6zPuGI7o1
0bf7uBXgiAECyBAVgCUOchBaHTq4FHBGQchhRFpeWXhGyQmvVIY9hpLwwMNdd0uZ
Co0W5T8yvNnUTdwk86FviWRyaQNzNRGi43Xvll60JNBEwOOoe70Xr29JVs1XdFPS
oM22PDELtZgYdJs+sdkY38ZRC6v+nYMwg9fMFP7M92l7IviNzeRLlXWfFPqHkkj4
BndfW8qvEYDCa0YBOEW9UN+Th9HEaTimL3R1t4LCN3/JQudyc6djLTmymrDQlb3m
EV1QJe4n+v8eEnOhKlTwSZV1+1L1y1I94oLt5Tm4yoVkL4iwJdUz2X4NMW4KDu7l
cnS0kWl+5uSosEbAFElExkksYnOMKV+iOgALeSXXm0iYdD6qNAV5G/EpVToNmB2H
6mFLd/vuTrrEW1OtJC0D0sfAUX9JN7+gwqI6DYvkyJrs0wy77FHC68QU64+9Q1QM
d1FS3BitFIegVkxujW5TbUqIcGO3+cB3VNlH4EXuLxUcWCGn+cyS6+E0oZENkHeI
HNz9WnQn1fp309zOCI7yzhNsZg9TPfMpIzy2nIyEhZ5WZOMYk3hAfFHsubZ12wlO
XG/XpIwtZz4sMa9fGSrEwRHYEO/mkjPxKAvqkuI7cNLXLbVZ31n11ryLrgt0Gs/d
wNfyoXV0k9TpUR+ZMK23UADc6Z8KhiwMDG0WGCvmXRhyB/V9Vx3X2Dpe4CDOkgnT
jozglb7flOvr9oWTZ+FfiuQoWQJ3T/EAVzP2Sic1cGkVIQrSYSRWtLRWwu/DyaH/
3J5Nkpyo/WJYySIKrUOiasAeLHv6t4BDVYJTzhtql57fcPEVfeJrwtMLUaL5hLO3
4m8temxkO9gwH/f8yzvtjfoCR0lbW6eFYgef5ZyToneyOH4nnmXrvtZLpYvhbcjO
1Dc2Y64c4DrC3Z4/LjA2mlY15hmzp+1EVlk3YkgGQh5sv880kUTIxNtIkMsKulO3
TzSvQBH9F/hjbHy0W7HLZ/LLoxL0lABmhTte4LTEj23V3h5nc04HEdanoGSxVLGp
NwtaJ+xlpYo20Mcvae8+8TNlJQlzJN6b5AigFGqEerEEKUETEqIiUOdpKfZxyY4d
2lkCQGHY4HrNuOxWYSSlBfranHjqudkf3pmWSFwBMDf8H8pin8vWpeglE6Ym2ixK
wbz4DwmYhXMvQXxGfnXV3wXVYD7CT8oC/yvLNj4UcD3qNx6ERkYhUtNIIz37CYXu
J4Vu/m4jKlXII9E6CYlbd8bHYwgi7E0lA40xT97sBzFvEbh9h80KUcMtCGPrbkWo
n2nBoOqHDsJVo2BNg0BPmeQ6bn/6RNIbX9+ITinFgR4m3+ddsq1qfgcCQblrIIRz
3uuNtcOVPYfpwZ+OMgdQn+tZdez0DRG1riPKdSHclKdBBvcAnGDl1DbYhQS4yGOi
K/xs68xAXTlzi0AVIlb5d52eQDgzOcc7DShJH5yq1+UBlw9lZsvXtaI4lJ3UbgzE
eiYJ0WWfvJA/b+35Zbk6ZGy7S/LDyaa0oxdGAKx+xjwnDDc1fuambUOvUzmwMRnV
/GPmHFMyk1qmkAnidlOwEMDsrIGKSLrCo9Y+sBD//okoOueCuxrQybFDwH8qH6oA
oPLePHF3TIeVUXxoADcU0O4F4tIfFXKK2+bgXTfYi74V32yi6H7aWI0ipZo/2eh5
uS+Cv9zsLkAHOJDshiIaYLCYb6NHV0h0IDaGolD8goO/RtRydL8t5KnhVH2Zf4l4
snIhIZwBcGRbq7zFGng5xJdQuYifxsYbhn7C1aiK33d75A9rFVbJiEP9W0x33C6V
LonAc3UBrHpH+6nalh7S+AJpBHbCHzPv0gZky+mXhoxotCxEvLSmuNKtcR4gePn9
dhHimMRLOpRGvFKKMpoiFyIK9SQgzWwai8rn4FACeqmZopv1hgqn5kfkw8Jat0z1
cGcsP2Uw1g1tZQ5kG2G/STOPbnGJV2CADexuSSir9YjOQJqNMtIul5w9Syj2pABh
AeA+kRmEjJPV6IZv6VQ1OUljH8/HQBGl7MQI3VRoKUzM45WKFfuJBresnqGSezjQ
ZDeZBW7SDkNKqsRojkICAxFogWeQKPvtgqv5iQpcE3SpRw/XWEUADDUIJ9PcsDTc
b+uB5oq2HYSEfRNysRVNQO5mJxgIqIt7G7JrTrGoYxomiT2Q/sLI3D9k/yKqpz7l
Uj7uLW945vOkO4/Nam0M3Ba9MeOI8HNgDyBSmZB+qIxOKrMYJQ03gheZOa9KTyC6
1QsSkQZIus6jvgsAT9qpbpMc3y7YDMPuh1Oelg+t2Uxeko16/ozsmijk+nwx5i/o
2vGCmtEdLCntvqJumQwCudbvzrUxOr24SdrGydCFIyTs65FZ1LfkmpqIrXn3EVtM
LID7myza99MhnVRNKsZoS1Uznps40+ZTSi+YKd/QWg5aKBaleUvLlt0EK+2OlOJF
l/Mwn0r1gEWlOgV3SAw/ULu9UZaTyGfKtqSd1EMUh7/0f4q1eq52kNdzoG6r7xGG
P4aChcoZ0zmr3gJ01zXnJEnc6UyWe2vdrvzWDUaPVV1dL06pERh616wpXMgYj8mS
bCh7zk7AOAeru9qIgG9n6aE06HkKw3MouMzS8pHHkJ1Kl8YaX8G0v91LL9ND8OWk
cck8GArU8JGmMDgeXERfiHcPJPbUJVnhjYiVLOJMCFVnEGQo4Z4RRVTRuCa2m3pT
j2HldhnfFRAP+GNMCtdUt/oAIrfysIaPYKLAB5kGP0syCM+C0neknz4RGOKO5FQu
gEV/drfhW5Lbh197VEo90nBxIKg6T8WoutDvDFv6Rzkd3hS8botW438p4tFOsf9L
wxtW/DZ7HOkyQA4KczoBQ9pOLXB8N3avgyDZTY0C1C+pkLCRze5CN1xC/jy2/jM0
XPrgr7vBqzR+B7WdwO2ytVo0UCZD7oulj8TpLoYZADiEvbX/SYToWck1xrtmNWzW
eKd4ubuYKxiLUDV5TPU0xkVpZzFMw0DGip0aeepSPXaD8ULramDfytaCgktgDbbW
QAxj5eSqx6NidA6rTfFjlSVZKY+A/yjlqiYlIcZCcpYH21/oj/N95vZlG8dEumTV
d31m9+U/kWsggkGgv6UAwFrSNTvs3kc6eplJq0eaPOZsIGeIEvHsSYJhfdk1S6lu
tR1eGu4vv0hCnaEP422kmsr2dCgZyV/cwEnRqEhLWw1aDKGOZvhCnXeD+DoHs7gl
Q1/23Q2ejUDKBJyQycpg7kDVzeTwNvZSxe09rlaoT/2l18p+thxBwjPZotZ71pTk
/PfkyfKaH6oRZO0P005pAYAVx0BBkM/J3nB+bTydm0jNEB7RiZPDvoe2VKUXYFAk
qnI9uu9Je8VknsU7m1ef41ZRdqO531vYobEoF9KBQNZ3dmy5JdK7352ZEmAho2m7
7alHsuHUv747W4IvFmr3fFpwzRIeeLt9VXkPPOZN3IJYFnWRW6zo7+gt9WicFZaR
VwZNCowQqzxfNzVAMKz6aIC4kz/x7ZE2phXr0FsPdQWemiYFBAByVjceky78RPvj
6hJECfThI8x5GF4xTM97j4kG1lxiLFv0rVFNlptwhQR8Uf4y3KLRc0lrW/TCwYK+
R+VRrRhu8Wmx7TT5qRElAw54JZ6j2cTq8KQFq/FGmiiJz0X4f+pEK1NtgvwNUD9M
l0Zoi7rxpMZ8lcaWAz5ohpIoPAZJt8wUdw22tNKAZL0AGh7gQx5ZbmGSpdpNaWlr
JUK43uu5Xc2XTwfLh7qoZhskP3dIu0zxJspb/HNRXKzTZ3x5X2o9t2WIHmyGOHf2
U1Cn7zAzM+XqzuAaewgzvo0i6Eg7wqA8d/NZn55e9DgsCD+fBz0iptUw2q6zi0DT
7xyb5bCwKhpmPLaJASpw5upKuJdfa6LKERUEsfkYE1vBQL8REjegLokzwER65R9P
ZWS/ckcGrJFqUCRf6YGAOoYiirO1fZOKlUwFrA0PmWLxU8hQ6cpG4IutK33ol6qK
0cuq2udVz1cwgc6dJRUy7uD42ceHOtbBOnxROAC7O2u0VhSoeuMxacG9mvqvA5Fb
rpheNMOzLPfiuvKr7f/ZYGSyYnVr+TWR23X2dZeorAV1JWvot6Fa7c07YMoZSep1
dZLksFS/cJnsPWOMd0CkBnX/L+Np3NQmxro88jxOH6WhpXZpH5pdIX7v/yBvyJii
MDenM0S2qrXdT6x+4UvqYtW24GGZYFpl7OMl8XVZ0DHw4zrZkNOWdQbtfLymgwoB
/bkTGnpCTtwdh62Id3Apqeq8WqnwQFo1HJTTNwC0CisePainz6HRqYipqoQnWyCz
/G73jxK9tGd/lFQxNADH+s9D+rSfnFPo4d00s9ffvoZs80Z0cdqqoaCvYBUoY7qn
mwdHRHcBdN1z6x1bNTiW5NW4ZIEu1JxL/sxiUYMnUHpjmOEm6RdWDmKfg8ZzNMx7
SCWvWA4otC5lP59ZtkZIcOTg0X96LLdRuEyI48lozex0EL7wlUNbEnx+f2W6u94y
9vEV6WZuY4OgCBs6AbKIs7NEax0n0mcPjWfB2hMdaAlKQbDVw21/1n4X6L6Pku9I
r9rq6z4tLX7W5kkfzjrzbuVVt6lHFVKjpM4FLjENxrRUkdsuVCKgKt6flPFWSUF0
JXjuCD9PMNlQAsUTQZJkWYyoRzJsdBXaAqxWnKQqmtFCY6uLxX+UvgRHOxf88z9U
LtTZF4SqmB3HSW3TQKc1MUEORt9byZUL/1eBWVJj23cxW4JepxK7oKeJQGVX+6nR
MMFcWd+uPjNaBlPvzcTaUlWwf8OlljzIVx48LpvGcMOfv2tkm2TFdISKne/Wo3xd
u0lZWJc3VK0SA3Lbkg19xFeR9+S6qKaNDJtijT3PmWY4ARyDfm+qPp+87PMR27Z3
xTfTxbXWsUcLhJnrA8F4xB3HYUEKinYemFvPvCo6HSm+Hl8JparCO8RyBHt7Pu86
olH/2/ltslDFjsXQIpLLp6mktMbV7WvNvFWwmxj2nSD6CxAg4HlSDcoOfm2QhPyV
MA2NUMV1se4fFcERN6g4Au6IJ+xFUGMdwrP75nF6qTXFyWxb64ykBfI6ba9aJvil
+jEbyZ3wx1dxNz0QEuqhfR4QVFuG97j1wfXlZ6zbHANckBit5+j4JJI68I2rp2AX
LnV4+JZ4tqgB3T97KeRFpYR+Jw0Hhh8gfpKMI/Ec+sM2Ij9jm8n2PId5qiJnutpR
1jtf25HntNjQCQp0BL4CZ4EuEU1SJTTlv4aPeh0sLh5lb9OVQzLMD+plViktdAl1
tiKXII9vVqG8Koo1LK3Y9g0rNXa1JvvzHUWi2Mw6t3+WwJ0+Oy6oOJxB6DTolHJ9
AJ7I42YN8B6cdNgDsFD9QZNH+VEF633G0N27FGWrnXF/HrpVDFn66P1ECTMwlW+r
kYrS5hA+loeWxils3zONhAj+bTfXn+JhOtTLGCP3+ZMEC335bAzsioSEVOfudR1E
5Y0WMhFYxxvQ/qIVx0eo/EoCq3HJ5exeluhg+p/c17TosZgYBi2HTEWdF71D6mFx
HxAPu6fVsE+XnNm3MJHE/J6fiMnOwdOS48WGAmCaejBs2RuOCEdT5EAHVtwjenK0
hhX4d1Qn1jzo3Hlhag3KpLUIfO/KNVz4f2O5QbNoXsoB8VDy/KZ6U+SXgDnLZISD
nPf19P+LBISVflwnxQdev8+KHl5WtrndgjM8FwQ5bOb5GcuKBVtFCj29NHfJq/+n
XKZzPk/MbIppwRUubF+cNUBGV6/+NEeY1I+w/o0kPdJn4Oen4UkGGEBkJ8YIagRG
tKy8A6iY5XfliZ0zbACEr1xC5o4NdraxSpeODMWs+mXaC5/W5TOEA15mb9++CZrA
kkA/MqshojpWsBEkMCkYazWM6Y79Y+R3lMjQERUNP03+Y374Rx6PlPv1HDhuUq1H
Qp+8s3X4RMKHAGuDxyFMY/nKNJPXo1O6tGmQbwAVWVR6qTSyEAkYcF6gjR68xuRn
oRgLe1tubbhz8c1BNAC4nbYJyep6LnooNi0PT+ySll9vOQpfZDqyOtUfS1m+YOWb
vXD1Uq1Me5f8yYRV6FbRL5n9Hu7ru5SVY0rW8DUgUl+w7mGkLJy3zjoia4UT30Mx
iFtQfrHJ6G1jbRZHBfZ0GamGiM0hL1wWPqTneN9yNbuQehA1eLDHFydmdlywxMpn
CpKn5fVLZK1m/Kk4yrsrqso3eEt0oeFoV01snF+EBXQBXw/Ko1fv8sMBvRZ3i6ee
7R2TlhMFTwETOy9Mc4I2104bQhsYLWWgsqjEnz7IeXY+B+nGekBbD6CCRbs5g+jO
Ibhz/i/PlNupZisbhJ0NDrv2xTQ7u7Ewt3NCvxRk+R1KcqlTs5dFCyeSmMMvNfko
+oyOiV3r6GjczSS9CTJME13ABw+PGXSBQ/KdnhGQjCClruth1SlXDFRhdNh/auqB
q3LugVV9pZtj4WIDgGF52iActFQUgLr6zxzqaJKT0y8D/sIQ0ghf7LLH4BKYDv4O
P8evz75GUpyGySxawvTyJSDmw30g+dNYUCIh8PETIXang7KYI1IBmANNxQtBk+os
ONhYsS4aJJfh1hxEkYpqEbShUibbWkHGnLWweAtf0Lz0iM/Lpia/U3hNKBMvMsLC
+mr1MCUA/ATjcE9b8wAocoq9yIae7H+jXbtdmoGAXfNgTb021ONVKMqk6lPMWZ3R
CjqQDFB+SW6qk7Zj5dqu4524kVIuyhQfQXQcExBMEw2gPZnm+UKshJYSxnBWmivj
m4VbXzYL82nfN2rxWXG5kblXbKxnZvth/rK7KLKrOAX677jJ9oArosVZzeEUO3Lf
51a0KSYOwnDFObWmQ6y9liyF3S6TpAlGNxZN5oFFhVM084MwtoFNisi8bm3MrOyw
WABPpK6Ch0xVqlOQ1ipPdS1XMwfs/D7mY3aVCDAdqESzgGcqPRkYfv/hTENcj8r7
hSaw0a4rmkWjvKbzsKti6UiJ15GADUBWzJvgS3Cd+pd/tiDie8PPb1YYTguLg+BW
Nx1D6hMeXN9flOjK54KulCcLNDOqYMiIWj5jeAHv6r6sVqYudHyuw8km61gzKAMb
vm3CAQ+Es3WxfeRWwBaGZnSm+0gYfrjes+lKT4Ag6sDO+KG4puLkkfC61hlGIetr
6DDQIMd/FACdwm3TXV43EanVfz8ZoJJ/wtR/dcd682dhmmcJBfOxmvuvJQPX8nVG
x7mtJDQgxvOPujGWfd5iRuGgWOUbowoIEOrRwn74VM9gC5vInUHcpx8SUGRrt8RH
GEod/tKewkfe+uO7IsrlAiqUm7DkPcM5lEZA1DwuTd5we+IbWMNjIAevZ4bZBmzq
3cs1bTIjBptxmbN5dUJG79Gy3ZWbq4ccjhPVHRJNFKHgJXCSpPQjkoHMjYyO07uh
g9YhiDYZBd79dHpEo3FZpTwfGt80CwqEnK/M+4LZUrG/7ioNVUTVIBrulLs6/B1y
U1Hi4PX+n69ogUzIkSPQWh5qntufuu/dIYckhM6fJlgAWWYkx0eBbIfaNzEuRcDy
vRmHqOkelJFzkWGjrzsn1Lzw0kQRZNJxMv0z8W1PdZ8EURSIpTTxf42KcOaoD7Ez
3eQErH4IJsf0iry8prc546Opy1lN/rpjPErBaOR7xV83r1xL/Pv7rAgHl7zTgtJa
2+GxjxLkfPMW3wJWCsINh/SGf6ZvFnJ5RxhHGtCbjoFcPqlWGTYy/b35hoPK/DY2
/ttNc3pPb1GSqmxf6R57eELKYp3TJo47xhfEM3V+DUuL3cqB8r6M+igow8neiHEi
sm1GdbN07LUmIGAtcVNN3/YMmyFnAiHYHKkF7WhTL2b+Xf0CYhqYt4CKy4efzfPm
PHltU11Dt7EJNAN+TfdSreGGy6M8YNFyy1oeUfzPNoryZ+TgH25UEht59kAlYFVG
hT9czu+O8TZIF9Jba5e6hqwXKn8Ldq7i4AYIXM6hncXCWhmpsx0DpShxz9c9CXx+
wE2sx/o5ldJxAsF4CjtJ1u2SMCS1FnAADCt3VlZlmJ/32xj44jQ+WHDHzSfKK2zI
f8C7cE/nqPhFS/bDblTXZ8Wq5du5t0s2QBZEcR9NLjZYW20Y/TU4fENykNza7v3z
G9wfknJyt2I1RHzdqYiIrydIbp2TbehOLMdiXs/4y54kf8CR7YkWDp8/GK+nvfyb
iBIzJlSTBBoaheDTdi4FY9qyzPMzWpoyfkROhx0OXCfOBSymbirnn1YKMP/1s00S
Vm8deh3OEAngXzkgM675kA2knDS2Yh/UDk2xJuJFdz0OzJMHi4Cnk3mwUJhkCGMP
IFE/xckCwhDyoU+PULvBHZOGfo2VoJXhVdUhI4SY6imAdcdkCWn+jCDtJFYPfTxH
ummw9TDQjCRGmDw9dNrvUzHoSEdrP7JribNn3wqMwfF5Vk5gRlejbGkye9aucpFV
8G+hpp7+pSlnnllRgMlLInFMHohhVzTOG41NL5N128fPHdYuKQzvGgfYVhZRNFEa
P+Y//8wXotvYY0csjjowrjTQ4fU3m5+VATjzCAy8uZ9cJjs5+7cS6D9RJREzwMdt
n+OJ/Q13osDVfI/br8YP/aM8k5+lAHQQYH0z4ko+hWwBa5HIMLrLWin9mT9a0bHn
SwqaVIA9O3rlW6eysb3iIb4yFAYY9fHDCQ0hm3nK0iMvun89znR4a/PReuoSRzEq
Rpw3R8xE7IdIVOeuRptEGdm091Lc6Ck0/6WHn/DxazWD7iZE+bTLT23CtC6NMk4V
TrP2qHfS15QSTco4SF5aOcmg9YWm/AF+zxeZ4MLhS+TRquUcTUTyfLYw0UBzh4jI
rjYzFFiO1/AYcN2JEDVWRQZdJFmqFFhAk9lxeAajdtWveR3302FdPrOpx0xWl1pF
VbsRXt2Ze48C6tmwZ1Raed5MmnoCvQnF+IsGFxQ4IctWO/zOZJcSUXcgsE4zPE5Z
Ul/sXVE6/s1/a+iABmszMLupNkQKdC/R3qNdvTfxw2fCa2Jvp/JQfZXejZbxg0GU
7sR61TOeXubZrLYD63WczHTbeG/m7g7El1L5+oxEvw5KATDytyzX7tS38j+KVAtK
2wtlEv2weMQuxe7JTKepcspEIScWymeekd8+zWRv9NGJ9dPk3/3tk5F4JCArDkci
BZ0GAxFpioUSfihjSAGDhOab6q75Le6syD3X1s7Mnc0n6YYqewvNUpd2Lr9Z2+BV
NXs+kCSgkxa8FW1+GWNY74NTx1Hz5RN6kKllUAesOFb3+NDX3i56cOo0FP0M37BI
27rwiU9S6O4CRArza+pzcC5CgHwgoAK7LdmQlyoAwsDuy5FF3958xZ8f80QZSfeJ
OuM8Z/s2Z+BrJLwbyYhxEBtAWQezV7lZiFkT4iCjEeSF9NoNy9Ofs17RO888FKtj
7PueDQITJgjxLd9dhuTtj5ZTZcxQepcYD87ungiglMyy6VHD7gC3KXO8/SogrTiM
awXQUM7iAhi0fR/nqK3PIi6bUagMNySFlADjDglyaw4lw9M3srlM/wvXUcG5Rrqp
L8pBHpmVOQxYE392sC9cDg5J9oLW0puglNZ5m+zkWfRAaSsXgAxpDkWwpFWVHV38
irZd3siR9dcJ82dBS65LiCIU1qZR7OcwWmovsZ/VKg6jcUfsCaqv+965O4LZoW5L
8T9wxlpXsTeUteW2VvTMcIya/LH5QM35O5Vhbafs98xR2dOfYQLa3dhssXYV/DTr
l9GpgCyg92vt9Dly+di2ySPciQCZUE8UThnTv/7JhIbgP5YlbDU/C+2ddjbQVt5B
HzKidS7Qg1QvTXr7Oh94ndKp/5Hcd7O78q/sYmEeiGEhBl5OKYwep8CAV3NJKBsF
Twzo3DqEAdOVT6xq+LbLHw5j4G4Xl3bvwfgdPUJ8JP0TvEUHd/C5B0oM2NVilBCN
xY6phVps82Sn+hgjfqXGuPAEfMsknLDd2TJjNUVQO15abVFxN/KDjqGEZstEzZRS
E43Mw1z+Vbx4MzW3NUysZpNqaCODaVlcrd7+9HIQmfc3MIRhbYACWKnv8DW8X98+
KJ7srAenbwU82tSks96gCyeCsr9w3QDaBxbWCHUHgc8HBp+I4VaRWuA++RkhXH6Z
nbawzHS80uJuqHYfv73TrK8hLZpER7614bbbIiFF+GAdFk1N/+TSpSU8i7MCbK0r
8S8kUJlVqYY422KmfAXBLREfKABrobNK73W0PafB4O8ZXrz5LRk8h67iEJSODc5v
1Icce3Ix8uUY29K+vqkGuFQIY1HY9WzUj/+D7gbQ82PEarNhJGtBZg03f6l4siNB
q3s7dS6iqZbGOtIQLGCIUDjbMMrnoi7RBsrr+Cu7PHInSdFKlhDLOVsV+97bFWlO
MP4VLQQpbe3XhwRLA951J/Ok6YKQOyzNeedP+T3vuocbqAhI6+2tVnJvw/hjUg9g
F0fLXsqX+vC0ZzNghFjgh2p6PiAFYzKUo1KBALWmnff7vkAvsgg9ZpYCCg85QHr7
mIuWvKEUUhtLA1yykdFISwuV5b1o486sSqeFSH43M+NemzIrZxXPlGg2ZjUaJCAy
WzJ0+M1roeok0g6hiryuL3HgWitOP2oWkouJRyLXrBmOJdPTciIJF+d6/j2vXl4r
gshJzdc+AmpDq/zApUghEi3+LaNe0jaxoHRuZ/iNxNrdQ4fjIMcucnNEzk/zx9g0
JUmBEu35Seu3fBtRTaeCWMVjhMs69wN1tmi9q67jZtGJFLQR0Pz7HORX2RsKzFjR
bGATfeH10tYqw2HTPmYkEWFs+vXaea7sapNAfrWCQYtO08DJE5kO0i2Uu2wAOMEb
m6a2nmDx5S5WMj+80g3FhunWMYQ2R6CxDUKXev5mg34cAHddB/qcXbWW44vmd9Zm
ptBwO6I0grdlVTKd/V5oOvxz5viG6p/3gLbdL3fbV1i8dw3sD81lg1w/y9/nJi5o
xHEgs3Zx7Atsbm9M4vorfDNOQKccUimh+fvWX19XONsWwwxTqNjiJjRF69VfG3HD
34jbio9ZEWjLo/Hwkzv+qDv9ANdTB6p6gUD49FHPjikie/sJQUu0Pr8V4/ox/8L8
RWRffY7P0cjHXamykkjo5KqzntvKK0QKqS0I0plYVVBJZP/gWR8OXEAQObbC2wr2
m3wJx0ECpkB4jMVenp8D5dX5JnFqRhLbB0MKJcvglmOMQIbi6mso9hwoCUP7f97s
65kCv5JCycb2O9tOGpkt8rHc/fvPmv47JJKB5eO+xXNpreN3pT2c5w0ftf0qwb6B
Jt7u19hjWN/CBOg9EvQ1QUF2odY1GGdvhGic4f3CPuhtXU6LmPHpy+DhiBnfctEq
RwxN/9uAyYlPcuwhNVfP3oJKkmkfaHgY3ehTYG4s2nHmO6rLLDYU2hV2Mv0kDNJG
d4ZJL9RH4uXgmWIVlOfGxcTnuCXN9oCUkmjZmhxm4qDFAZ8ZnlTDWQOBf8n4Yp44
qzrX/cLz353CrqjfrCmjnDS5IL/4+Ueh5LLSp7+jZ+nNJPmYsHdyHTmTsea0i5t6
H3eppZOKsg4rUH9lY0FhbzbDr1wsRnNvyIG5h0jJTWV0B8zaGMXWnEzWogN+8+pY
r5kfFcBqdCFXCHm8lvZvGk3Ro+XGDsH8veh9WZ9WHm2zYqMsPUDz7vPplXKDNxm0
yDeIDrz7ASyTA/pacpmd9pNe74RH42FKsbkN7MIZI9SjXCRm2a8cthY/nnK3h1HM
ebne+H/8nPxidmcYoogYlK4pZKuMoqTpkTG7hpU7+gXgwkW5wwM0SrnPFmMvRvwS
wjlYJ8HnsKMELV2wV5rGNn2Kl9B+1/PUNJ19xB2NWdKg2Hj91Yb02+fMAPuANfPY
gBN5jsBSoJ0F/JJCv+iLBmgXQNPE2ePleaVfGqJ3mUmOTBDcgM+2J4fhjDWOrKUE
kF2vdyVLSQAxo07kpytek/fEkkEJ1HSS8b5jJzfLKkN5p+b5t9MskC5fcCSfv15W
bGwf06HwPAry509vVJgeTi9tKQSvkW+JqBfrOdfSv/Iv6wG/MpWhqNL2NOvntARq
RHCMLdlcpQ5SYiTpwkYAVgTqxWwSfrm9a6b90uVbCVCLNzri2ZaQY8/lraHdq+GJ
QkeGCdz6FzPXXJIui6cr2Zr8sFLm39zTRRokopeccxwpvaDbNV4EEf1tA5vEJAq1
RZeX+AVFUbzTDDgvcA9lpl/r2267Bw/baolYJ8WzhKQfDabKAxiSl6/1IGkhxpn9
XY88pGbhJackgK7yExBeJHGoSUJC1eSKz9zVx41HbciteOCFnNpL3ZYPWK9ikj9u
q0tm5vYt7iXnBbBCtaNJKS5y3D1QM3mv+SzmTx9e7vbydE8u5NUfQsyQ2ZxtQdPz
tpSf7+KhpUkpm1Mb0Y7yWBJwTTE75qGGa4hUJvmF+k3C0ol83AXQZzvcFuFe5rSX
0fu/MTWylzf8y1x/aplw6KHOC1RVFfeL4Meb90Wc5qoqf3+nSHhFgyJ3MCjwly1p
5Ok5utT6phQGN711+vL24Gjc8Mj2jCBPreoZDsWfFI5yCvRmH06bogYtsc0tBXqW
WPgtKKwBDeRFw8ATREJwgABmmwUEUc3uAwZhmlaohFx0MbqY8bCtauiUto/eGh+W
jDC5pzYQAJD9pTMDG4ZR6sdO/Q7AdWo8WuWzJNaNalVd4doG7AL2nOvD2hCaubap
ZHcggHac1ILDKGiZAzAnj36UzZCbFvwku4xf3ugXYEAl5HEGXAS9KI+Xv6xCnmhD
UzmFlSQ6x5XN7z8orBcPoUcsOIvB/u8yA+3PUHhl1wRqTgfq46pY4BkRFqVdn9cG
+b7xjwBea/b9cg7tnwtdYaENuZQ3Gg0+++ex4llXYBtt/+WsDju1hcR1twKhJ/p8
0xAFIlihEfRSpRtCWzrH8OMtKXtCo+DabIR+fM2vI0/YZNfF3FeqAXopt0RCjujK
0OJaW3ErWVMDll6Hsf86fnZof+GAM6v2mN6tbKrTDHwZnHYslzeRwd791WhyafD3
WgINZ4ZZqe7jymM9XADPZbh9FK/amrgP58lUeEdk6bWagjagaKj57yP1Vj/mLiLX
cZ82ChLKkkmT+Uggv0hm4fTy3MOQnzHcar2d/3vRF+3E5dGsdV8+BC75F8G3fiPU
8WXw25meW6/YqdsHOXOMCmJlZ7POE0ILTJ54tRznirXCDhX8ztAf/fTZEPsHGqTn
qZBmQ3zjbYNVIwFFkMWqVAWm0NIMFm4z6RcuVHyOUHxyqPuRWrhStTXb6er69gh6
dFD3rWuw6f3/tQZbbtrI7K3sK2z98cxAlggfBhq2NfdIUXWD1RI2z3mZOVqlwM/C
MEnMuhTu16Ap8R7R8lkKoBF0iogJ/F75w6rLK1NE9JuvbpTFUGADpPOQ3na7WIyu
+UHdHpao3O0YLjaYklGXnOGlANBoZikCdy0HtVDG2LZl2u5hzM4X0/RMTbSZtEJq
3RK9wbV8vljJ/kja30tc1S7XINYg9Hkarusvsu3f/9bAatBF5bFa0FPqTOsFWnjG
cRyWBrBqKbk3F5grBLbjG9Fz1bjblLCJA0OXBrEIVRr1yJlkwxpG5aRhL6f/N0QG
1pf73RSyNJzy1R0gZE6619/MhoJqvKLtVyFoBhDbUZCJJ61gDdpawCGCUga3V9sK
NuPxqP6YdcYwfF0EU0ghvjuNJf5SnzoX5h0HlfOknSB/4l6WVpabAvYNxIXZXl/y
YeGY7rGi9jb3cUTYVEEp9qDa2Jx1iqqrtRmNPPy95EYjdebIrPjlv9OvPYUXQX6r
oO4WaSkk3QqL9ZhHLChEsy8jQJtwHjdLJG7RXf+WwYtbyXDGoKPXp3u50apeFofx
nBq6PhiFnoUNUgPELO5aJRBvxWxvYOvIh9DaUK5iJlyTBoQaeQ4PiAKxLXYZXCMq
KuPEV60fXcyFBFY3MLIjqqn1f0skY3g1e927mZ0DEn8XBjnIufCwyiYV9AFj7sGc
hcbfsbT/1jdvF4JD0iQ7lJLR8kyjs+TCQhtN1mK5K0e4G3RwLr89UCmVsKD+/Bb7
7D+DqGBQekQ/GXkZeMFHIPkzKNU1guMWf+XioKzx+arRbaoVyZBosjltDbTjLVZZ
f8kZG6KbVJo+CFd5xH+WCAdr6HHg2m1+nWYYfAssmWKjEVdH5+kP5b/cAw0So67X
oRLarVx9Ad5uz5GcY0BGJM323H3TvjGnMqgfK/PiXpWlwws/P1XKF803N0mwLpHC
wri8teG3o0kehMfBnpz34w0UTsVzFOoqB+vobf6TsMN2i+qB7VfNlFUG32MnpH+a
nn+EQ6aTkXnD0g1U412SOZbZnQFPRBpHtNMCzxz75u21Cgx4oHnAwoIPZNKOajqE
VFwUbKhp8swQchWAD4Jn11hfDrkiUZAymFZPJyrOAvTBWCkYjNUczk/UHHKURZJv
anXoVz0V6YUuLHdw5n1zGXEU6vz/oNt3lzPkkoVHjFgnKk3wDwQ0K7ZhwM1eyTZo
iNqjX/lWMY9L7uyBfKiCYQZsEcPO6yIfS3JiwNELRj0Qjjy8iyVbV6+EiZaqU2A0
2zzGXE6XQ9feDX3d1xzg3fJUt3+L0hy/BmUdkUmK9RBEQvo/mprY9A4p1WHLQnW8
jQ6RtcTyMz4ZBoHvv8pxG99Lue8oiOFAE/Pq60QE7lDwFw2GpklZV58KeWXvw2v8
OGr85+u84NGErdN47l8daYRI7UbFnyM7MsJ5CANOrYmF8603/CCoEAkW9ywwe3+m
nOpud8zWN46nqvKxACap3K3n1Eob4LYAoiFzlMq0ZyyATNvvW6WvvHwsbrcNR84A
mcduSQ0/3wnxSKSAFVUIQSzCUXI2E9BENxXM9glPf93BsiKzGq+taK5dn+CvZOgs
CUJXDpak4Of6jBdPZh+ATivJ5NkSYKwn17Pz+enJD210DzmteY425/Pqe7jGPVzp
J3UdSqFAxGRhtbuhSfMfBoXh+lj7qq7dCEc7eFZfmtXc05rTSpCgG3dyoiCx+Vr8
glYiOi6MveqOT2LJmN0i7HjxujWi0eya842IDNL6GR0tegPmujtXISpHGpCI72f2
t8DumOmTrHQnpFyUb3cz3ImlUEdMrbfwSlLzo4ZnFI+XDA/PGEtahQXikceTwnlG
01UouTtVZfr6/rxVwVtZunJctOxGP0Reuq+HyRNnkXCZCjzE1rH8Jv9XFGDojL+G
kxRpGz+MrZ1ZMv1CYkeb5IxUvpOoJQEq8/QYxy0ElKZ40fjTV/NHTSNuV/GkQ+/Q
IpJ4/1OPeOaFdrv5QFtSXVntOWPFJHsKzRCKxCySqUL8Mak31dFl2J7e2J25iFYJ
5FvQiCPfKN6FjVOjA5dHQotDDM74tSgIo/z1zLhh0exi0q4tD1T/xmmO5JW+HWQX
Xs+v6R3nGeVRNDvhW0A4oRRZMeDiHPErSyG0pScM8oCDQV4qyDxDcGhrxo9IqluO
UTjl/vW/fODfSsbzMOBU3MzcwLXqv87z7cE/Q9gYxghR9Rjfm0r7r6lEuimx2xbo
4KvGCKSp9jwqjY2XuUUgcggrHES078U2fX9S5SusQ3FDAvAWk0afWEhpW6uqTrht
+pOOEWRjFWKCOdKIrV+9RjwvOP61JpeLA6zEhHoZre9YhWZ9hcKTMFgAOUDH7K1s
fHsQQDgzKS9h8v/2xl6RrBqa8xpMwGkkJlhNDv7SCpkiI8aTIwsazVPoFOh3evi3
6ir5sFI5lOdK14YFSfStM+VUlLzHiLDyZIGCGCqvNO6CwWcbwx+RZcHJybMfOD9G
ypsn9Gu4H/Wb//QX5scvnsA2AfR3cxjf/+HvONs4fotxJgKmte5O000z5iNPLFMa
hp9wloL2D+zX5rgKXOiG+HacKlCVJXH+U77dWUN0LQ7eioQrsW5sctyCkm61CkvY
HgDhPWJSn9TE4FalFGxjTMmqnDExZOfAW1g0nHTQiBIm2mzrADUS8VBg2prjmTHl
nAuu2+gVvnOx+UXY69zGllVIAbSh+XsVV4IZo/NdFNRUZoEqe451G1/tBfH5tRgC
GTd2XwPFRm428jtdQm1GzaODZ6CNF8PbBkJQpD7gmV5f9Di4PBfScRAaCdw7awQw
a93djjyKE3SQbyAZrCXld1jSV0nO2E/8MG9MTWP0M3uizvTpBDU/QsEkXzNJxXCN
o9wcHRcN1x+Ila9GsU+SEeyBzbmDA2Ly+wOBkOvQWr/bpAve+ZYaxMvhxpisLoB6
qkF4fus9cvwzzsvvVuy5SlzIZayVPXw4FJI4ipVwkFW1JFpcEUjxKXBfs/Zh5B8X
/oTyGB/wB3czKP5IYCOFtfydq3CguCU3ClRCwmTVuXsS59wTfX8oF+hx0/ByI30i
Xy0cAadUhoLpiAqGfntv8ahe/WFVcrvX2e0+IIVIH9bMtP7FZdqVB7qVoiZXgSwS
K+cwWepxjpk1hFrKOrOr6W9kLLca7Uv1ErCRhxvJdJbxj8A1oKMdLO+2ZeBAO1l5
9Lcz/fO7tPVgUEryrM91KiUAnETbyP8r/u+wjMInd8KjFusQFDFsg8zb655wXWkX
UPaGJMwpa52nZCIvuDepY5cqNLLQb4dKbPe0trTEBtt2lj9YNDJUeom+3FqEFpji
YJk3eSDVTbpf6zgp3kuH0DyRZgjmCqPhvQBggeh3lOgsb/d5Ts1zEu5zoPGqxZ3U
HjFrFRBhX89ZoNkxCsafKfqyXik5ysDQN8dvAMzr0A2xznYfMg2rHJ5AsUVccwDN
2bqL8nPiqA4RzjzkSlvE4xHBIllVHw3Ktiz3NtiCQ5eQ8OxfToNN3ozzKmSN2iAA
g+T2cK0t5OTvi09DY2BmcsuhnCXSfjRfeBMv0eZp5ukQFPvMiP8X67EJoxvQ3Sxe
d4xpetUL2sNPWXSHsgrglv/mMepldEqDlnghxVX8HQF4shWxpBxHY+OBU/gQjk70
6+yyowYZRdTBrPSxxIVolFGe3kiH5BDtBQ7bf8/fdGyiq8ftbU1J6QLwBP2vmrYK
ufAP3eX5R5XlWMo2PZvqSec3lLs8PrViKPhQu8l9X3KZ7kWI198Pbz7/HGWYDyJw
nsBptvjdn6xGGNv6qh0U7lUEmEGHT9a9yoe1tABR21TIhAdlmJ4/VKRthPqeDGNW
7iKjRZ4KVXkEC06VlcALrFtEdYc4GQXStouUH8tuigxSg9rf2q9uGg+82t/hQRqj
PuNaAvKgGAuaNpnUgSFfVyhajVGOnu5ExyqV7ZWpykWn2UIuYkXoETic+KN3OcZV
nWuH8/d9aLNE+E3HXauxmZ/oSiT+X5H8Fi+p/725YBxYkxwVQMUj1nfJOA1yKWyV
+JjyfY2ANRdjVRG3KLtVoalh9zxmFVCwfjTcHJmVa8GsBBhxjUtAXnB/b+vGEico
+U29+jQl94JzvOGxD6VEE/Oiq/q9IRn3049XJYx4yXVV53zQr7SZ2wvSnA1Tf9ou
wKkLSjS3ybNA2/pwsfMW0qOCA7u+uEHCfqH5js0ovdGMhi7wRDhMuA5b4XV0jmu6
St942/COBLhUBfgQTm0T1OS/nFo7ljQvFpmyLTMcNKpSkVMaJZ+O3rpukSy1Wlea
iQ1Tp/YhsBxLL0WOnTX2PVjCcvZF95BqN0uTZIBQxE6iHMSFfuaLzJeLi5jysccu
Bf8BCBi2YRU7wdqvjhqZFjb+0EW0zSSDqQxqwpkz1XTwO3IDel8lsiV97jyIulfC
FZjB6SFzBXdcc9sYbhu1p+Ym6wUSN+/C95eVaiuO2JJyPzCeBxmKUKGGijUhGSwd
9h4LBTh9giPsS8kp2MRhxwOetUhlzJ2aQ8rGPMN0D8+nhz458zg3DXGJwmP/+RDN
fLu7ZO2+T348Qs4emlzG6rKI3MIMVpNNZ/dQQRo+8zxmB/cWQaVIZ2txXYwCcE9D
O0RfebSd7+62Babya34mquIrt81uFlx0Gma2sYLouHt7X4C47FcdPfTS4PILIBNC
eua57AFmEwTjAgw/pgLxQonRgBpvFJgB8dLkBdiQ4BpIU96vrxcIzwkLh9sEoCL3
v0kgdz50tcmT12iUaCnpi74AZOVEYqd1gqRXgt4+ycXw5sGlDxa0gc/t217u/4Zq
Ac4vOa0H7xpHoGX1KtCUhX3zqvcpdy28bi2eGh5AKjUvtya0il3HNGPRnvt9k0cJ
FvyWJe/ZPTCcFiC+bRjg2qBD4TzlzmixrwC8sI4UKAVcsiY51BjKmrFypp4sDPpY
Tls/R0631CT7OvLJYqBE7+8hSCYE/SMuVEee1+dJWdPknzAAlHtrOUh/AGgav7WV
nioMzqBJB/DIbEyXGuxsCuAAvu6fz9KEtn8vvZfPZSbIPJIfKpOMokWIJFzQCRLX
VUjh8ZrmB8FH1dFiL2fTn6oxSeOWMnPattyf2SGza8ymeFPKox5CuS920ZXasM1F
5frjftfYaVNMqrKM2HUz8mBcYR7sEKbT/gvY1MwEiuq8IcOE4ROKzN4yvkohYNRL
gwktWLxNFDbh3xr/1HRoFjAYEOlatghkBty28ZCk0byfkNHqPiJOKItuRn08cAK+
/jeq4NQ9UijhKrjMa5Co3dVucFlGJw+snAsGNn0hzOJ82V4pNto5WqKii6TXH+oH
EcYM/P+K0M8bRKGrtbC0z7MvBxb9xLF1evFrudq2Fft4EmE8KYsmVpByk9nRvYGa
X3CGCooC1QWaRxZTfcVeyojSIPDFOYrYheIblofhzkOOiIQSUtgcxJKzYPac72CY
PfFeAC5vlUpcxaMZS0lKP6vaAPVEw8mf1drtEEFO12KWX0V7Kr5AYjoyTeRCDMhS
45gn18kIqiFuzy5IElAYJlijUycYtW7T/rMmEXfJfWWB0VqWJB9e5PZ3uWJjmE+l
FPufg6xxptfiIkwf3HKb4rAgIocU4sdNreYV8dUY/MiBwOaEzgjkxTkiCIAsu2L7
kzpaY0ySSST2Sg5qwqsFHo5Z8rVcLDbSB1XmLtJeBarg7r8SVYL9fZWy7smrCAFw
lCIVq7a0PSRxkUxTcY/qTef+isFOJxz5tXpi/R88Cy01N9jFYbb5Cgly/rI2LauM
h0qqLsbhi5n45HvS7uhGRqxRqirB4oLPIG6c7qMhYgrZS7X9WccWQwSTMG/AiqWf
0rsSqY4nQvfKkUhWmqwTAcT3SXBXK+b4AoU8C4Jp6uKvxD5Oso5fCj4qTpuOuwXC
gKk3kU8mvvLHyoBZqPpYqp8SZIFOs+NaAx9qhs+mewwc+tTaC99vAWskEwWGAFaL
FPypaExUMmu2FJER8bphy8dWyRfPXEfE0wFiVpqL6U8ypXiB1hSrx1ZiXfnWGVhd
3APNiyD2dc6wWsRPpVyl/akWUweiwSOTtmTOawabLM7eOSugkP+SomksWL9cvv9v
NUMuAptoBXMAd+X1xrZ9rUE3z2DiPDws7yIc2E5wWsB796CwhnPA9TibjiMknCPX
x9t1hxCh3V9JqBDQRwcV8TXN/oLgAgFa7j3VtBI75Bmp8WOfUXhTzqbzbyEeDxWY
BwJhLbiOCPJ1s5zrkhhqqNAM41dQTs8c0qCSGiAM0Y/25QUmNc8f1WtkDsFaOS3/
LCz/rrOKVcyUUKdgM7ZUxF1jf4pMCgePeAV8iCqNs1Zy1jtgA06IvDokJYABKwh1
cKZmWqmI+NlVYvBKOYZgJTXB0qYlLdr/FGGcG+w5zMcbg/sxUcT9pDjsepYZMzk3
WB2150NuaF2McdhQ/nFcGv6Q6RNprNHLPqcQHFEuVwh8STikZuRZ543uFyIx0zjX
I3yR1HyhVhY/G0sEQRlD7f8akeEfpLSflmPH7YiIcl0/Oqk+sPFLD0Q+Np7vva1a
rK6BRsNZJurCHoET7+WZWLiV9x5u7cVlYpgvcMnW+FaTrUkamMkAHjT75z0oOPH+
JAPGOGHrq/kAGNeOt3MFB/KxQdlipikMmz1JwQ04vWwhqRmeWFkIai+6BMW+wyx9
AXazj1zusvM9U/41nQ+t7ifWNxa0EJ/dNCwk1v5SoWDtSCOduaEADG3QiYBoXL4q
6BcBOHZNe47ZRA10lwDsF67ANtqTQ+Qwzq5w25V3Lgm+nutQfHalGDhDXRWiEO3g
1k5yp98Cr7n4lJdMi9jVKsAMCmv3WWGSNCNXcaZXns4+N40Mz0oOSOZrlFpaPCIa
mK+XfV0+fklZoU5zJ57/2kl7YwpprbXCAEINPQ7Airtkpt0VJxzjS8/nGzZz0ja3
WrcixGtyMLt1r+s7DC6yvrlHSzoZxNTX4gYGX3TT9TO7TMw31l7X/lTeiFwkFliI
Wo3Zpo0iPhbVUrQpJjH7fPNgDXNmu7Iy/E/UghG6LcnNt3u+C/bUr+lxh+8kF0MQ
YC7b85p0/qiolrEU0IgUG919M+Khb2tVYkFkc9XhApJ7pvsPR1Z7TOQgj+w+pOtr
kICauPQ6wFc8gD4Xu7NphSYZdKgkn8y5PP9ULEs/kQ1VReF3mQWxWrqsVVfxvHKK
n+T0/hahLPvgWxwWu47pXnStpVKbNRt1sZje9iUsnGBlcRjvl/wr2ukaWFBzf8zL
8EfPnuYxxRp0lK90VTdKFPzKveAhYJ1Rg+54DbWQnTf0FNJoxZeUjUJx2Mz5h7rt
+Iemy+ApgzFOwxKrvssTdEhT1iORa7MVkl0hD4WF9gYLuWSctYzxqTjoVQ7dig59
inAuAKmkwvmKRl8sf/BG4PkdrhEoBVBbhni0WM6mBsAtz8ymPbfFGvLd+fd/runq
HsVV/dbu8tC+cyFbva6QbYnSwiBEgE3DGJZf8BC3DlDCisk1qsPKsNGU5ow5p15b
DU2IC/v0cqGt+MsR7FSNZal955jw/oSRIJud0oIapnbMfO0uFvccqYqAaX4RwYpu
kL3XlLjE0p0jDXMIF1Bj72JamXYk1LB703VWLrufFVpx3S+6Ro57zNI7SEkMGRhQ
z+AAgsfU0gVxw6qQf2wPUf4OT6nHTY2NcCttdW5Yg37OrjF0TT9WSz3+DmQEo+xM
HtTq0Z81mkbF80Bir4drIBO/32xCFTs7CmiGzgqHHgM2OsSdl4KYFfXIlY+L5InC
KiSUZzwwvtPcKzihh2BbTmrIJ51UUIuv0CnMkzV4C+SOQnF/dArIAvG3/MedawBT
IScV/+1sX9mbevcAlrHlOJVTLq7L+/7bO2Z2TZ3DblOH+AfhxoMDne50GhaNeH+m
BlgJd2/kcjg3UpZEmpcd3rsCWgE2XyOrRQ7krmFRoUO16bgcLEZyP299k/fQFpzi
Stvl9B0NAxU7TZ5gY/ntVSQZLtawHAf2vLIU7mOvsnuLPj4diRtx/cCDJ7CdbC2b
Fzha+rl2qd/gX6canCI4Rtm5LQMPF7gbLF0aT/41m4VtZZlPTbdR8MvKvGDvX8dx
4j8bYfXDCZdyniAoq52y3Zx4FBNjPYLIL99yoUS6ABrPjLIRscEVolDAaHAEFDwd
EncPX0fFVMYVU/Rp2jfn0xx/+EKAWfAV2oxAxXJn0HMXyAL5nKGuyeBU3YqBxsU3
oOvuI/nREU9dxR3N8LT5xFlIz3+Eu9banprLiDhTSwazOPpbdgJx/MfWksYEyUS6
68FDIkwYIULoaomHp++rQEpWpo9xRT4CLYAmx/VGKdTcqhrEj8rkUBYA+PoRaACh
ITPJA6tpTiu4HYExuZjEBKyMEmqOI0Uzv2Sndx2sg/2GU+judTiQj/yXYqFrrgQP
WUvfEqsxFJNGpPs1zhPpb5eHadQFUDWtzrRZuSp06KVJixWjlsR/jWODP3yea0uS
eyot3ykDR6gqSRqhuOM69hAnE/DsaAj4oW8lWByPS4rDyjZNriyGgHgk9NfPU1w1
s10n2XZtNJMAZH2Kk3cdhVABSA+z9GTQdDqfDQWABUeNcxwHMM5eaDrwjERHQoDW
HGOCiXV68Jeb5sd4xIGPvG8ShdL9mIn4oyjdXjJRHwQ3Ul1eUuNPFGWEbR1DiJ8V
tkGXJNPapdwawvtzry3WG5bLa5eg8IYlxdwwlmKEMwGjQxQocIqDdoujstz7zUzO
MwvE+kkaNkvcDxq4A7hiH0vi0czi1dtFjJ7xwO/wj4hgyFCnm4WWxnGF+g0zi4kZ
ApbRsuocuZ3nhPOmg0CuiPgwr7pSjQNQn9zAtM8fM6hTijl0mnHseBUG8OZhhS0U
4xw0uOjCbl9etnSAQHfzbcrp/H+TsjBq1xwbVV1JNzK+Ijm6pgRVZeYLRZz758AF
qzLP4tMmmTORQlKfclwedSFmmD+Tz6X2yF+h6HH2M3OLw/NNZTEuGuxwsvTgd3f8
l14//Ddv1d1HrI0LlIP01+/vK5VwC06IZRH+Xu4lbxb6EJWSpP+4M5gFPTfxZLBq
DVOfEzaT8Jg4zpUbTcOcrphGKcTuuNA2N44YSHxQgQuDkubHIQ62FT6J7UVN5hng
SXlsVIxoFzfigRMSxiABQ5srl1o3tTFNAp5umBez2fP+XOCdBoRBGbiTEk/aJ/3f
oZmoyQni44IheR9RG4EYhqs36B1ii8/3Z22gKSfJ3NeNOPMdXgtzGKfRpsCAvS3k
G3I3p1kXresV1Q5MSd9StFU9bQo/xLfjyLYUQ/ZMVghBc3EXOVdR533RwddfjnYr
JX3wNf3l0c5ZPSW/Dj+OjZw14EKdxIpDUa7ErEX339W2PkZkSNJcANFHmTRm+ME3
nIvccUuaMPa7fKVlTiGxQsXQwA/9MIjeLAneW+oH6gau8M6oMT2E83iHLhRTx5Ty
UqWAng4Yn/RfQQUgvENC7Cc9R0QmYGDShx825wK7qj9vVMTdz7copTezpvlGnyxx
o5svIejf2b3WznAyIZ4CK8TZhbzqH6NqRMlwTmqd1/MCUU3J5he+n/SZFQfinJAF
+WBGLUn6CRO7qZXUWRm/2xeCgiUBnXVXUjwrXXba0U9z/aEnVL5a4fapIDO6B04h
14eWIhD/Xdraolr1qnmwMwDuskW4BeyDH+TSJytriFIQsqL1cVPBghea/VUhZWZi
4Qkp0BFWcJFFtrv6LveTWloKM3QzMzdKkhMrVx++3msnVkGeyMEfQtzoOsQRNIlN
oyqkN4OIPeW2ekLF5Zq89J1hcpAEZwZevQ9JJiYlLCLjIVgEAeGPK1lKeRybIglw
hGHdaBBvKtmRfFwAOTUTO/3jXbrmzyIOD/dP+yy8WjnhFAp0r4cpJOn7x3vPO9Fq
+d5ws0KFcbqQEYgYptR4wHvIjsPm/012sFgV/i49ahJHxQEEQjmMnEkZZ1cN8YGL
tHy/Pv/Sx6a8xzhmmOIaiETzszSDb+O1UGqZZk62A6b6bcxbZJt+801f9wHI9U3c
1dTW8Zw/zrFrUfN37+zWBL5SJ3fEES1K3j4+rexsfR5PyjfzPhp6rIjVRAVnSeUD
vWBN3z/G8+n1vAXhpL8cqATjaKojj48EpSoned1hEfx2uR5AnYeu8aO7lJFEvAdI
g0yJBfpDcUWavBQa/i4s46iC00xfuZTu9lWl41095TSQ8suTENDPSjyZAVoinCMs
cpCqTV/g+taxtWyARF/X2hu8oQz44z4pHb2pnm4xjBpfbQ4mN8n+UjlLtRRCj8qc
ed/1Fjs1/ihlgxbTd2LjWeC7LIR+IeY3V42BtYjhTRvWPuteQDgZrpnQWFmDyoSv
esPOTGf0ds0ote5FAx/bdq/+f1UIAn3AogI/KA9pPn8hY+IaiuQJCSnNuNXUMJwB
DuRP4D1UACAxoHu38NRy5FOtjH9I5Yec4T2VG2rBKhI8V5PWgiSHrtuWdIeF78f/
iey8/ytsLYdsyWN1VITHqo0ypwt+Zm7YVNcWfWhcSjKPo9+kxGuurkIeSFoR3dz6
xZf9Y8iZdNX16pECOZA3K2uUXRyYPh6+eNb53m3jgPT/qNFU2utTfckmZivq1mg9
tx/DlxkXX5qGO6C9nfBtjaULFUd9VsHKyfgKEtHbHJ/qOmhn+t8ak6ndQBrjumXZ
mWlZqiJt/5wZcDyIcPB9TI1DIgZ/B2zRcoJHbuS3/zugVnqdwJblVBTlXMcyQYU1
vKoBrwH7zUCzG697CAvomOxysP0jqIUrQmUA0fErkejq/spe7yjvNGrIeTeHhuuo
ICLwkVSrm/1W+PAz0R0uszF8Zp2/kRTHkr16pCDn4IsFoIbkGE6PTgJIFo4kqP2T
d0/qsnkHXQo1VvgsKjVekkabj/Usj2FmsJhFuVYSK83cGzfDfvSdN+/JgWLoz12Y
U9M3fMjP5a/0QOvigdRif3gOXdboytnloMf3TlXVJwyeX2hR2QwmaIawxfKIaS0L
k9lHf8eq58LiljSbVwqvDqyqGhYprHGzns2mw4oPv0GxZipAw5+OOxQqXvmhkiZF
aposldAyHxTB/mEOJs+hWW8C0OD2gr14CRxPgaZu5HeSkDnM0KqeZobmjdsIUDed
8B/Pij1iug/XaLaR9PbQiTL/8rV0rxf8qHfxf5cA3Cxs1qPP3TUZepSX81/g1Du5
D2Kh7Miho1SYE1jCFjDGJpLIDY5HsWiUFrNQgcTAzvcJ2RPkYc/tDLa0Sqnv7TNg
vd5lBRU1VoftE1sUW8CRlJOC2ftJCDnkcSUnsEjHMWQmAHbXoAuARg1EtTRsTE4d
w+LQh801SrrqYGQ3bs47WNXyeO5d1MhxA2DrsMHXwwuO9m9MZ5izSim7IP+CAoKQ
N6SmuvhM3/sR4kVI25ndxbv5IShag2MjFULtLVo9X9OzSSzfNr+laogmNIiiUsRy
Rf4SpyUjdaNGkGuRDe9lFLXdhRHZ2Qlhdi+Vb8tWm2XOYl6l1ce3hs9xuBIlFImq
WUta1EuIzd+4+JXGjNU+Q+PkEfKvxjrO+IDM/o9sGJGajrwwUlvmql23z6ByzfSN
h+xJpxFKctzOB/sseNSvhulF//T2AuJ2pTsnFQ67dZmk/MFc4lU5qekXD3vLEcmd
twLuZEA0Y/kLVgGrDIjJxYG9o58U2Ru+DeCky9fZFfj2/KGGf1HIAZ6ooZieOo//
N1xoi7FNtMZuJfFHiorINPs37q3aFSGP9AddynmrmJj1HTurUxb25L1zxUsizDVk
9KOBFWKw6kfRbx3+L3GxJOxFAX/tOORpgowREC10L/KVR+b1DMqAUa/aVqxRY8Ui
AbImfLhpfLVIu3hdlVoQSqI4vEPdmw8pZcv4m4JXAfrHY3Bgwdtg+HqDQtR+5blb
luSI/M3/WQxi6bWLAZKydMyN3H+w3BnzBDe5JacG4HL3oRpb3w2trIcRqPCR0EUb
NJRhdKUoVPxeW2DAh2VJLXilc6dnfTdhGCWyHz9puZQu6UgBvyKEr8kJJLXIx46K
uxfNVGy3QZtz9WOFiAmcmF7DF5qxlrc12XH7xbF/uwcsBuJoPyd9XmQM5gm31EDA
RsTefxnTZ0pjb2MKWqvISWqwOJ1M3s/LYoQojzf/+iTrKkvHVPz8+1y6whGZ/ISc
WJVjYv1E632bKWjvLoBbZedq0qaENCdM8m4pvUV4oI7XX8sx2etA/yP3LDP7AxfV
s/mMqjzPHlu3dSQ/6q3pM9oJ+x0PDqeCiaDMJNAH4/JpFWkrB9sb+Aj5wc1GzGhu
+uymhotBmqznZXs4qafi/0/o79j4typlMfOibV7HNLVJuRoH8FSPAQnWw5fcf0Qp
UcwmW2xYOLr++KItRIZQjn0XylU/E/TBI+aUnhhHRd1h6sz738iWvGVj7NPa6lgi
s5WxYSJKRsdJlP7/U/q9GTSu1Sps8fNyTuT5oVoBK8cHgulPkeTTpWyTo1RkkOqP
GPljeamUc3BI4q26fUX6n+Z42TMlqUzKfocwf02yU/LiRUNGmkaynIbmgD7E7rKp
Zf929ApMRCFc6Xwl++XGzkoKp5Kgi6YWCrtFdMOslAyZWI9zdlHP0K9Ocl4vDMR2
Y1rJwivHtlV4N6KM8TnUN9oHJF8S2OuTPJ6cHlmfkFjPU4J+IRj+jUk1TKWVkHRo
2ykCrIQ3RiL8VQjU4hpyqqLY5etmWKbeYoeoozpd86vi/vbbzY4p7jWr/fPfkLJt
//dn65REfu2cGedm0/lTfxIs9h30Rvcih1RHxUaREDX60JE90VNxn/jlRGINfAS1
fsdg/UqCtQRXdLLNyQKLvgqsN6vwsQ7vYTudJteSXkgUnfqLF0AlEHnW9kv4bugx
gAN1hdCekGPnZ2izLfbdOC3jYbK9VaU9wXTyrDONYbMzBJsQ/DEHNXDQBdPkSRFd
HRS9F0UWapB+G/R2ztNHOBSeyYN99dbDgggDX0L2/0jxITocD2+Rwr9XGZso5gu4
e4c3l6vbX0rMlVil6SiYfUHaGukt+99X3UFvrzaw4Kmldyjvq2mithQYMrM+womG
r33zRGConeTf4vFlM7/qSNCJNxJroYIuBE1sn2ZuuRbSedzbnR2W4m55AZi+YOaX
HGgvuzWUfrZed77rEJ0U4LiV5VyYnIj417pK6KevHICbmlP1aq8291nuFqG+IKMZ
Yflcm+lp83lyu1DTe5Z05alQU9gUsZXxDRYqN8AJBtqjRLCWdZ9v5zeKyUGywchU
mm6L8axcVptpv3hITeBwxxMfd2jrYYvQ+gfCTr8YfJiVNB8oMSTEuGTZ776qH+DW
Qlv6Wi4mZmBd6PjaRJtIifIbyu/oTdxUB6gsnp5JzvlgAS9La/MLchN4TYax1+4F
hGrWJ9OZOgMiZClgeevsowCguqCJFFvHpufLs5XIGDP77lukE+PRY6KNko8pF627
aI8QFbcsOLujLraOOtE0SzZ5AzsuKvqYyBLXKQ3FR9qb6Wtn+PRr+iwZdXgcq94Y
Ypb2uOi10VwvRAH4a9lARSL5QikqtMObaR34xaYN88krX1worucCNhE41msqE4Lf
GWzK5G634MTxCyeLcMKpue8LZ5MEMJ43O+eLEWFfurSTyFP51xvAG7doJkKvgNZL
mo/7PVvNnPRliLDgIs7pc/C29tf12pfGW9Z+6oUefV+YNePRmtTqjyUrvrsQ9e86
N7jZi/GXPdqax7Jv096TkiievA9pguP1SGRTAonl4I0W3+2K7R8bSC4+LNoujzwv
sT5ScAM1GGlPbrvM0xSnwcUmeIxJA05L2hv1XqPZzij4v9i3w2XTkWWtsQyQr2qT
MYcTHh2YwJYbLqDz8U++c+LI8LfNWCzgJnrfPwnccKidi4yMyARiBTCWVLBXiUSY
9dRiKGYqcKt5jLtZtRukHH4W8UWknDDhVNqOC65/W4YotdDkPxTAS8dPbCqZQDIW
Xm2HfosgB+mjX5Wvlub6uceuQgmCw3VV/+fWMCxH6DExq8k7KZx/aXCkMZokbWnC
+ZcHYt8J0EmjkOwaMxokCCUiiCYZWsc5FAXH+nCfJ0lJS51ZP5BPFwIAhKAxEoeA
9Me0sqwFx5rIzSXtiAwTeEoTCljGjEA/x+rlDcoJ3LDQMl8wk4iAklDBhT2NM2CP
bvzyeAQFi0VuZFc+h720NCPA7SgTBRZjfjIvzjTPRwrAI9qwORTy2QagH7Tliwvg
W//lY1LkhUhKKe/LqaNRiFSBymFo6HDeQOSF9seTqgrn5meoL1AEltb4J2m6ll8a
wvno6nJwx9OKNHcUgKjGG4XMtdkINRMZ5hOxV9bJO4rZfVKk3TFDx/eWszLp7kOj
Iji9649NwPB+ZB9StHaclAf82GIJn5rQ0MNkzGYNnY+ccsKvr3G04MaFm9xrY61Z
RCJ5VftXkGii2SwFTi9uFwOCApVX92LMGjPkQJvO3J4CxcuVvtC2aqQgZUfRg69D
I7Lzlh/VupZG1GMZGqE3fwt90AcvorZQjSG8PXKhg91vNBBOYZH/l/v8ZmuQKvnV
ijdrI3UHeSae99oGEVxrL5ME1YwOq9KG5obuEmTMlzHPVIXXx6I91D5ciZe7Dir/
9/nliccl9a1oq1oTBd507lnbUILmqr/xsko9Sv/UvLlkR5zD+/9AMCgMjOs+fU9t
UNfU3R/vwFomONRUuV4rW0p/LQ6Mg21xccnVOPRwaVOxj0AcLucgoXp+gLGy+LTC
tNaZKPfutVt3Ynbrnqig+yqtgJEcH/TsLIGvGnGuzY665LMpPrcqKIcycKDkGVLr
MaskARAN5yfgv3ytr5//1hAFy+WoY2w5yDlwHhddUNnojjDiG/ZW1Q8scsd9UckV
stBNI8OEkuYdFslgKmdswa6jRa/+2mJ66s/LNszUk03on0n3CjR74RLvJhaY31ct
Q7o0V2Lrnc6k0E89Cijx+OIx/IdalEVnswhwlyiesb4ELkrfRq4DrOkfz+8QDJUz
0IP/JnPTRi8pEp+wBQ4mjzcMDlb6ATikdBO2VCgMp8QdGBtlLRyLuWmS2Ah4JWjm
UDTOupIbrX7nzx/rw8L2GC+UkGCKCja0ULVbTSF4SAgCgluL61ALKNwtj1aR8C2I
8UPvyA6+ka1Z5bdxsrcwoQbL301u6HIR6d4r+tLDovh8P/w+sYziwj3C2DmydFIk
ZS4be2KAAxLcmddsV5qEdsgPEm/M5PDp1G1u62JY8r4rHy5Gt+uFpr1TcYMOxmyr
zDvagBeyRb24+UqLf+envsBHnIwdVXBLFtmMuD97lx2/sHGCa7sUB+44b6iaPyan
ikHbt8O+l5QIhcOvdZ3SsqRd0c8Yifs8WnwA6GvGdoSoWcKsyhRjV2pLiisN39V/
g87P7+FU64eZ55egxhHzh2ef19AYNrD18xQFHaJEdQAaMVt7L2s86XBlDVlz1Exl
teo4zq2sxCRBmcXSEAfyHlPZXOY3o1e0PbpuJ2idjc89XtdLtlAU18fgqVdupBuh
SDFHuhzrmKTB8OHm8kMzaBpsqvF/ssWc8tpzSW20S94gJPJ6jq1ViAnRItPi0npL
tXtzwWDBgiJWe6Co9LvbYAjtIoORyVHxfyTWTiAcsh+z+WaUcXIPaS3b1K6XlQn+
kJlm49VwPzjEphjaASS7aA07sQEwOTC+yZO9gb8s4cSJ2sWh/fInROtjL+HuusFD
GJA1GYANyd43d6Tz1A2KnKT2pH6nr/3h56TCOmxBeVHBsF/QNHYNLTTTYXTdwwlZ
SUJY8uOjkjtGOXmPM891liQqLCMEkHJa+4FZH9u8r+KxDttPBeyOkf+QuYEGrsrj
/DUF6EKYgWIHz8u+c79Kbpr/cHrPMl8LxpziM2ctRqe2omg3aZcrLXPWPonBOcE8
V2qAzo2T/yGdV+IWlhqeK7YXaoQ/5lTmB1H9Kfkvi/Mxq5ONUxFoe8S/IVnr4S+G
yNHP3aE8Y+X+xyJcC26OaKKwDM871whkujpDYH95cQ2ZioI4GWGe+SR7WHHAZOj/
nkCrtWLC1pCpx6YEhB6Hg3L0wUkPEe/czkXZ+MtAySw4P7GXdAQ9hgB5hlh/L2Cd
8fnJUnrAIoJpRywgLBEAxwZaKEC+KzhNEiqvekjc9FMzpOsBV1kKm3Yi0f/CBpLt
/E+758ypU4476clY6YUUdIdTj2MAw7v5XhCZQjf7GIRSaaN7cnfobbvdVFmM8K4J
zSGGGWgeLGJLRyh7+DHhdPJGTx45G9EKyNtZ1E0HajDZRvMp+mvLjWg7GJizOUva
4f2dvIKN5kHGGVAG7qKxM+59VuMp5aGFEchV1Ok3sF4N1eOzu9D8E2xu17nraLVq
W8G+GNZ6Dv5L6UYUg19Yr5npfaaCb4LyfG6J7cqSyLnwFl4Glt/gMhovI+gP9bvj
LwWvK8Jj4r9Ibzf4ZwS416k9OaQ0gWL+WVLDUKb387U7vMwHWDDttUApGCbQkJx9
9j8rPjFvpeLj8mOyFD1w0yM0ydjRu4TZeYRY7wb8K+FM8TzTag4AcJCs9RJZ7caS
IGVuLM4Oi3koxGfStpdH2M1UggU5Ia6+mItStqZndoUulifWsX3UgopzP+rSmF4T
6Uji1qlP8YStJ4NNMDkqYgTdF3mVvukjGO6GxDMFlRkSzmNz4Ymp9b7YDu0Nb/d9
5IOcnJ7/fvaNYiP25RiNmPhf/pW+TCfnNxTn44yH7axPAoLrsqxvAINA0T09SAMA
6l5N1FmK/w8Yw23OurtWAQjG3CCrq0Fq7gUS2yUqqZ5fcddh1p4NvfdbNxizTEnH
+lK1j7BZqfqTXwP2PgQsa8FrjrIUM05aSK5SXDC97TE464zBE91CEhEf6Y9WfsyJ
B5U3IReBM0YOCpEE79kQY2KYkrqAHz0GBBuI0+gXM8oY38N8Ed+ymEAbUMEpbmfd
kXuShMQ277PmDH7MsrAZKlSxlQ32kJejycUfhFbGcBudMIIUWzpesYO0WGLbn0qS
hCjCSj2Nb6vJlrOtOTj0syccE0q+BTE2C+SUeyehYhefJs5sl9dBy+8ZwaO3oSc0
5c6BjQqvvnfvaiLkjizFJ5507nhOluBoQ7r6ub7Kpw5JHRvjyicX8SaM7EHqoYmI
z0Obqkyd/ny7ja8KDB71Y63M9jIH577BrXKZFA7yFP5kmvlduyewpRVZC8hY5m+H
Dr/S2jbpe3Y+i1AE9fKlp7Iw+E8qVi9lNZRCsw+reMKvdqGK4wMDviw1FQ+EYnCx
uF4Hbax9jQm0vyALO8g34ewKnwRtmyyvzuRhDvv6p6tT9B4mTfcyx0WVTaGTXpZ5
UIiIVIBmBPtVhVO+Dj24b11yIcnyPxQl2cNB0+fxrr3OUykU0gCosIILuV9kXTPr
b/RQNJj3ScQcpE/6NFYNCuMFGSdH1ApCACH1wfxtviK8B+5vrO36XgUYRlXWuGZU
PQSTfRLZRZX7KZk6nGaxNhmioppK27NWiVExbE19pc+ad+zwWhcPcp+KTOEBo4+h
G4+mKWUtvxuYldip/eHBXZifHjWTRM4yrdh3gej7uyxEAnMNZ8ValDhn5tDMeYwL
SGHjB8wkBBzTDewpIV6e7/VGG9tQ4RMQKKwMpAeDCf5y3N8Rzl6WPdrDyKZZHKQl
uDZKfJRvY0gDZUiDxdSpXuYtSw16nSOqusLjZ9JhqNR7GZr7Qkynba39v/oDpq4s
OkjnaNb+7U9SAd/Y1mC3OsclnOptntbpLx1cABo2+mvANyLBnThugVF1GClzoZh0
sEV/Frg7Kk1Deg6CbOY5BPUXykO6qIpOYFVTCL+/Xhq6DkobrRt5sDzQyZKHhjbH
Re95qCZsNEhfmfPprM/pjBUuGb4c1/VGDORnb+x+JIi3F0AMLQA4+4OP/Qdob2C/
yTch/qcO+kYbkLd6c6Q47g18dPqA3XPn1ZsC2H22StQkmj1Yl6gcOW4MepJmE3Jc
7kKwgW+v0qZLzsl0u/Gnc7ecWH0UQT8eJ8Z/kjnM6K6qzAibvbSFIqTQEuWQb/vl
wZatKi33ln7a7JmNTCfufQ85IVvJq6fedSNmJ49o2MCWvogASzh2A7DY2mnnsO6i
XVv/TNDTRa3wP8U1YiceW+h9DH0tdcYyhBSo7c0i+ynz9JZ/PwkZ7lTjjZgegIGB
3T2aYtojICXXMOxQopTagI9R+Mm1qDgasQOQfjD1zqGlkr5nZHOcW8+Mzq1ZJwDH
/agFs8NKmbumjV//+dOW0rbycu9wH4AcX0qTZA6rDKghiksxW3vu+S5b3rz2PG4G
udZ5GQxZTYxpBfXHChFTsmPlVrYAUwThGgXAbTxG6ILlrwPCxu+EAfTeJ7Rzl5H+
c4F+EOFQKKV9DE7FTzq34ypu25jQAT3ZZs2fRNQwBIPZ/dt0TokXBsKagaMmGwfl
KJxGkVJlzL+F7r9jhoiS+yFizaaQMZwu2EvdyQpFPKGxTTUWl5+Du9rw/BjRXQEM
WeeNY6w7l/VP0GB4mP0u2YgO3PFIMiEFowhVhdkSnAnIIpdwVKjkcXmb1Y4Auom2
0ricePNVlFrVEuv+4v7P7MIMTr5Z4STjKrPQAAd5DkHi+bxDUQZu5Vr7nbDvIlwc
yX6ZTwN8pNGlb7iEfNf4HXoyzfyIlC+mZedmhzvgfkZNriEfzPaLRFBdtxUuDc+E
9MZQUYUCi7IC9L44nnsjGRFBqICeZmQ8oq9LLmm/cTh422n6vQlthpaqIiNXQHlP
ofn43PpKekuVulqt0BD4FSyEPxfsEN9/ToG9zKEJomLaYnftQCmzNTdwCAq7V+mU
qO3nM6ZNL/UB3FX/F3w2nEKjm4XviPFbqOPRQ7kybfmNacRmPDDQ2b77hH7eED5a
QtkVHZhIbF0G4Togtr7g3CCIBQtZwPDfAFEWMBTQw6vIBxdDwm8pGDrTzbjYUEUC
MlJwVQEIhZYAy4/hZCOW+lesB+Lx70jHhzLcPuXf2Jsh7ZXZsWsR2U2iilq93+XA
7/SWHYxV85cxujh0AhQ9qdo92JzvCyHlX/pLzRnBkFNsax20G0iJ7wOByJzv2IFr
JL18pqUGfJuuS1brN7lpNC2n3yA9tR7V9FKypux5/JumeKufP0dKrz/0O0wWx0ZU
mMuGwWvPU+TAII1LaGD1kYns+xbzVY6obeMlDPogpwq8cfqj6MNwcXYeeMkPsrot
t1MgFhvOFAI1Q1d7+aK5o3a6BxACc0vFuLv9daphj4qK8ibhYKlLaJOvoablZaqE
zTe+pTENd3ZepaERl+rWDh+hiAB0vRXr4zbWBRFNROetXfCW9bzUaZQhHVzv7fya
R/FUg0uG4lMvha4UIKSws/PYPGzFvzS5IAmG6NT4ojpgN5h7Pb6stY1kylOzztZr
GD2yx1Zw8XDZzSEteY91Ncz62IU0rIRJgtvKQk1WrR9mo9Aykqd3Vufkpxa7kTjq
/rEa0d5jsxabGW3o5dlH8+EG55SgwidphP/Lrf555/8PSRaS8qT6RnZ5wga80pUw
EiysgMe2umYpfXvwV0fm8NUEHP07z6on5XT81rw/qa+djbBi6mo/beg6tyIJP+Kr
N15GphvXp4/6+jxPvRTqjCnzvmpmuZXSpcUklEXxauNE89EoOynkfar3rydzOVmT
NBCnmRiEhMQoH7gU4LT2Venfk7fxt62nGFu98vXxeN1jGkQuyZ/ORLM2VyJ1Ty1r
B2/ZQnwPV9jMtWNTD+Hkt4hO/2diLalxKMyrLOuSghK0xE54ME8JP17NlsT7qeD+
LBkIYPi3GZRt2TtI/+6wEAuk8HP+9pkzYBaM9VBP3FUbY87WG++go0U5pPALijBF
YwCprGqZfl7So+lcU72azFRfxsCAhXnkivqgZtNR1JCULSNCs4XyPKawAJVyT45D
RDsdFIQA529SoxBpy8tDINW+swl8AVCzy+F0zfF1bW/M4WmhGcKej4+1cmcwL1QT
Vp6++tL/d1+RfIc2VakPuNbo0no9/D1k7i0pkfjNL8yueIJ2TCZ88+6M0yXZ/n/Q
kZwwyVRhgytr3+lGQm+gXF+2XjazKpI5OHJQ/r9PET2AXbgAIIBeNlhECW61LC1m
LxsHEGaAeojghD3nTU5M6321OtKyAFbehiRqU2xsa0abY3bBQqcqwIYf3MMv3Ijj
r/xpvVvlr8Rwit7OqAfqlm1Btkqq1CdUScRSk56FEFu5aMcEm6LaYYTEC7OhJAGs
6ovb1fs5EItth7sMw/MHzNTX1rzTeC3xknGE96WKYqfBSRzcZ4PY/aV0tVLn4bxW
zAlL3zf+GVLDItxJC/EnTeGRyvh30Etu0M6/djhdETOZgEFOjE59mEEmuYYpTSHB
aES7Tyia1ghr1K5BhmXbTXM0/WXxphEBFhf3N8tP8F1nwLJ7TF0r5fwxLj5p1yum
Pxa0yZHcssm+AsNmfkPgyhyVPOuUZr5rdJ32nWWkZAzU5YSaf+v0yBLw7Kv47ZBl
skDl7F+2MMKv8aAujW6p77EFiNJoJTbygdjnrY/SwHWILxvacCD4Ck/pcQm5WRLV
cR1hOttfI8sth+hpUf2ksuqrAb+pF0QCFuefTREb0zwUrYaRnuvydCmTgNsDsgZZ
qQ80cTOXM3fOCb2F26u4msHWP7qaghLOttSxZL5vG/BloX9uqswkWz57nyVQmQtk
kfUlT7bR6tMSKb1gI0wMFmejKW5I3h/rV0w/vAPa8wotxPVRtSp/hF6mpmmPhIzP
MpjTU9g0reY/DJyIdOnoYLV9uA+C3scqJa50KV8HV37NMM4zkuTyOnS3kf1kuktG
C5r9/169adXiNvGDpJ427DH2FzM9skByNENRxFvaJ5RCXHjH+0kJF1q4Ko44Nr5E
057AfLonfwr+tfa22p4impCq+rQ4UffXhPRwX55ret0xXtPeygLRvLLzT5ZiTbhP
2trYR/qVHOoIXxTsOwl4vjPNjf/uCvverYFXD/iytJ3EhI0xBfXeJFz3TvOdgAFG
PbIherirVpqET9lZbyd4pB5Zz7Kg9vjKFpEPh/ZxSzpdf4vJkh82bIaJOZqrRIfK
69lEBgygZ5mhfqzXQFoxtVMrIN5+TgpkLZ+oANY+K+N5R42hirua4+yQbuZdu786
dBi9gHHQdoJfSq+XJhF7EjL106e5C6nFjOZ5A+bGiEfE/zgUR+YAtPS3/pR9wqwc
fJ773XlUe0jOwMzuP4T4OsaB1Mg1b1A8G9I5W9i8LKiaQUXSM2gYx/dh/iOnHzBM
7ldC5tfJPiK83CmktqKzz/w1VqUKxAMi3bw23DzukoLfqn7xOpYUvme7Vagky5oF
VZyAhq6LIQwQJHMMOl3E2sUdI9enl7QBC05CLcblG3x3yDMbAy9dG1V+qRSVFwt6
FmIx5NZFgLwK3EW2NUMKRKMqEJNfb18HlFNiUT+i2VHWSA+91xg+/5FbLAFDOsp0
KHcnixlZh410JnwLs+hIhpCuRCI+Ecyq3gg4FGyCAqhrU1iHrgXV/D2tuXZMX+m3
b24h0ik4eXmOPxFgR6SWgQqXT61iB5mMQvvSpRJ/p+ZU3KuGJNX2FBlxRVsfikM4
tgbbLKTBT2I+/ie5sHgSYBtKDCIIJ7fc74Z1j8/4FJ/o+J95pmplJmdfgDIVU80t
pouvkFQMJDdyanBtBOndfWLOi+J9kHiq60p8Y5shtma0uroZavo9qH8SGoF46erO
R5TFqNd41VAessAV4NtLxX+R7hJtigQ6z45pY9JAiH7djY/+vacpDlGhOC++WOXo
pHdK9PxBgo/X0csDNAk6Wg/6ejIeKPk/VeFgGQQEGvJOiUPA4U580EBCWO0la1Qj
bxp7Z7x31toeGlyrjaIdxxMMTTv9/xugGBVB2YqPlGObvRRtnp8wkLvCNg+Ai1fN
C6vsGWa/YIweE4wAnh3K+mzm574poAu3Y1lv5lk7fArHicTRkDIKVbA4eGQBIMJH
6ajNzzcL5pyLPnNMMXhuHiFkKfGSlp29UEoTHlOhDMqEqAbEJLNMlqLqBD93kiX2
T6DHf6h6WAiMf/wiegqEpjLQTHtP6EWlCIVxvWs518bEKTV3sqqoA3Rt1WdlsbOJ
2ssKeIO1Lf2BPWrf+qlewHGmnXLY/d/YJhkjuM9eH/XeUtKo61sIdXVmYP5N9Np7
o+Uh7XlXJaTE8DsaYD2rcjHmlvfdHrx5kioXfYkNIB91rz9RhKDNtnjH121DEBiZ
RNfpyGwDP8RcOPZ9cs6Vwy2l0fr6Ca8iwEhIPbXC3HoCRym1ZszuH/q+i8Ie7Qpm
RXUYMWGhCP9xbh87BSyMfoABeKZ+NpQAbbwKHt3CMDCH7Bzohq5g7D/XvkgIUeyW
zYx5+0BkxVPAsE8Op6yfhCaWJPnllzqts84CQciNkFCjGW+72WUKNfmhgoVDSATU
SRFf4uwfLz1HM6zIW6FklVVNkavP7r96eYy/42Jr5daqOQrNRGg/T+wzHbk+JYJn
3reImrnEsbjua7N0wdgnNG58Y596sSqtRAIjBgXwI+AYQ+CFYMs6d0MrOCTrxmOZ
qLQONAv9m0uTmGgzB3RFw3KTCI1xd6h3ApurdHWsrbx0G0k2qEzkiV3es9DNLcJW
/wC4rpLf/5Bf4VIxDF4L+0ZHIW3zQuuUzBV2Etd4O7Z+obm7nlBP+36DYz9gWImZ
RlXQP0OiFMCYiDB7R7/AyLxGxXSc/3qkG/UpGqW2uqvquae4O5XY+m9rxpu4mZqL
apAog1wZauYQu4ehUgwaHVBzcynczb84uvWk4uSKGzqHbvdvZr0fQoMUD5h9Qkw7
LAd7u3YAKDHwze/mMVLFnWR1fsM3GsiTWOu4tp5RAGbeDghEq2w4F65N3Hob5684
kiwb9nEoUntp7Weuf+unxV/NtuZVoLfqePfnpohsh6xVMm4nZpOCwtIpyiWJxq9e
xY0DT0Pu58OKnks2D8TSH5Mq0EmZXHd63tqv1Te+XpTrSJ05glVtVKMo+0HCXAvO
Q/j4JMinUrCD/b9Uu0JySsVSNIYe2a8PpGpIR2KfYuhlFXv0KnDdYTD0y8WDzJ1V
TUHEmvxSuKLywwPs33+BvnLFyVRpHdmQR2SZn35BuLIcfvaJSB4hx+EkbyNrwXiU
0D7QyVX3buMkD5BwG7+AZAV/ec3DVqxhN3uC6j/0l3uNTKjCbhLLKDFjLJCaf0C8
Ajbtycaijsru4UCLbsipipFz19whbORkvh6NISXUyxtIaPBPwvVGPvW/I2omAD/F
9PaEua1TpbTP+PRF7QaRSkjIYMMPnZKp1PUDSrJREYt8Mg1sdicHEaUjJhmlCOPi
BElv76F6BtFbrqL54YG8FzDLyVFD3BnPzIPwq1Qds8wGBQpCJrW1rQjOUvUxyyaS
hmgqdTDCVMy/OIQuMjLFmAn44cNTivsqMEgibkXlFC6rvpToMlMbcQ7lVYtsfbzc
JNRofKEIoGe85U++L/L9nkqN/Gp74Q5rXEpH7b4sdXyf+TeTqtJsbJMAnj5equ3E
H2syoaBmpSng7Qp6GFWc0Mm3HvRt04rWAW0s4HXcIf5z5eRTLD1xEAJXe03eQBJX
/m3auT3GxcJvgMl/1yifIUkV/oBT0WZf4+RYicrEjNkED5855Wt4SCx4PGEunzBY
Ov+R+xDvV+mtq8szGF5eV9jLB7/p5+CvvtFqfqb3wf0peo1pkmNwId4Z/mDuQ2kx
JVze7E5lUtlYNjjrOgKVmq47YbNQBJWKXYGwhBExif8kumbogAIqPkNXnSnUxQAn
s5oe6TQTtPQMDmhn/ZCCtYJji3uppwUJpQaZLTHhUhMv1T6cjOb1ECW3nlyf+hYQ
90nBUIHISY80jDmfasDBpQvX0DyLVMzldcipVnJSMtzNsJ8yKlC2shguaszxUHeU
H6FSHHk3Z9iEnAbu09iZDj/sM1/4a5fKTLebeIYELxrk83RU/SOzLeUs0Qden7hO
VMEDhdTTnt03ExQsK9y9g2WRiV7T7TfezySXyEnT68a3mRI/ejgw3CfFj3Z/seab
n0WfvetUDG7d/DNaNAoFs4+IcUmHr4sne+HMRWTbkaTymjqKChfZ/MdHNlqMMjYd
sX4CBlbYGIIlhwqR7iWRwp4u9mH89ZtlWi8BP4ve1iV2E6wakeB/BnlJWmOSL3o+
HJHkVGH6cmfLWqNcDbGZizTBCInwU3zjda7917sZPNozUXOPdk2b8cbWXOBc4KXn
EueXdbeElZWXiKA6aHN/pWJbZ/Nf4ZuUojxcDsGFUOiv1mh8pvwBJZg8W8XfURj/
bH2J/kAzaGwOh2ESZL4AD23cscj0Y4uwDOJWsSrFawHCqLXRM4usv3M7kC8Q2hCo
iDlEMXTYVwbXkIAk++a/NDydvmwLN/W2ktX35NaeQ/gQnLoMDi/RfGyi5EGj5AHv
UIwxw/wxQ+EXNs8bipLtDSlPfHgHusVN8ToUgMSLSSxynaSnPk2n6vgizud8g9QF
w4h5jtUpw86GWIJBcoGvmkjGvoz6AL2WOkHr5KbCi0R3igqGeoTa14lfvQ8WRdCn
1p/8j2okh52StIOM8PduUNWPQHnkdtGAWdqLL3wgaw5AM/ydi5tMwnpXxLroSW0h
uUO6vS9FIeGBlmBJ2uNWSWAEdJ0c6XTZOogzYkv0Dt+ATxq/Ky4I0dGzsiWiRs9h
6p/bm+z8Ty57xpH00IIv3PsMm1v7TVy2nS7MTmfe07b041MdhNjinehb7V2G/WRt
Zpx2ICMGjafCHb3Q0BHvBVEoZpk/oCvyb/F9EUqQGELwjqxZXn3zEIXPZW4s6t8n
ICZyoqbYpiuZ9yOx9XgBPOyxKwRofsPVe8yYnKyFey1vGtZfMalZrB11Zks8uxrl
2wZTqV43xpVozaHnkIv7wgCUVcSsxy4uyInmJzhRqJrwGyNJa1qAniYKKw/Y7ZCd
gNSh52kxUUa0G3Vqotidicwnb659r+92HfOsGhMZy6I8rywdkHNfLYVnvTFOc3pP
/y/HkiMwqR0OVBWDw637IXt4a7sxgYKNM1zy16qE32qPwpqvClEnkdhLNRji75g3
fwR6dCTtupttPJk9/87K3va6qWwqHAbV1YDa1xvi56JUPwWgABkl8IFFckdYZH1R
iZBfnLXfCeQ19H2mP8tX5M7sA3XsxfECr7bJcQmsV/VGMe45aD6JndMmsusJo26X
KecXCmWrPxNDdYNp8EMTTXExh8gVWeFJlNZgtHGvu6swSHbqMDYSICXt4ega89V5
OnHdJPgp7Ta/GPHKAAB4nBzPW65cVYSqJoVXxsBUU07d9XhOdZaV4IXGN5mfPrjs
wB3Bsu6Koxw7/EbBFYatpL6HXn7twXHAKyfDaZpxPeo/049YE7ojThpA6sUxYEbz
XyjlNusd7b7uKg8t9HGDqjJyEciJb4YaFZhHKcVLgYfDuSr+Gqr13dFBQYW9T/Ns
QgmyZrYUDT19CGXbHvPMdhe6SDCTiiY8WwoNQcxfYI9qSFoE2UCwloTJz9ck65/c
9uMWpQng6xCTCld7CbynqycvDXy62tbjG6Af/5cGlR919t0iiZ88fY8nlKVabFOo
bXUZuyf9aJcDxZVvxEBy4Ge8Q+S27yKcfXJ4RWtrx5TE1DYkn2ZL4ju0uKSzTpg4
tKP3f4jN3iwlIPEpOl8KxuW8L3YMyDpbYKC9lGa+n7v4QV0gJQML5wVTUycshWRr
ZIuICXWX/niJ941dloB71YOwpyvjDCe5FSzacSWFXpYiGSPUCyQI+qAApqABNL5D
QuKjVAPdpm0PTgsidNv+z64KbgNaWg/wtx/FiE7SJh8EjJArPkkpIb2gdc7mUG1h
X43u2MSDaye7LCLATbKXatugUO3DiPNcRXRJ4Hrg8QN0bDErntyVnSIyjlOAK/Ry
SOFCOOsMDqGVRqINbtBsmr4DfL2MyCnb6kdDyEJ6bCMuHG8c89JjMgLHJQwuw3Gk
BNS2nQobQ8HgoDk6ueyPebsBgm/iXdGAqltGdiSpTiFxXufuDihFDqqxqyJ3PWf3
LiCDqkP6f0Vn9yNeb/0RorRL6nm7ftuPFm+Q0Jvk9jW/H2WWhaQwn/1GW8GMMkAZ
NoSRbG45Lag0mxlAMFFt+H5XLCZDPSvmpw1EWRavOkwnSgDnLY9JHbV1T1ERe2zJ
sAgcWySy8jWJNrdXeFKVeyX7NOenldd4BD03RLMyk8++VrMn+9BzTe1dE1nN/TE0
GiSS9qxGVA9wN/DhWtoRt9OXRs8ytUMzy5qiusqQYcP2d2plNjGnkB+C2Tj4D0ag
r0dmnec3BTnmvhGf+Ue4XHXBkd9WRlEmXG9MB1k8tX5WOZpQ5LkYNhzIs4pPzJ5G
xeFixhHZniucKkmiTK6JdZND8h+E1X8O/YdXxIZaBf4sSDQhgkj6JLjHa8n+m8ed
9dZXV6+GIccHhCNdtoXrV2umQEPsFxYZDaR8GwSvIf3hn6RjdKbYUUlWRBwcGnW4
6YKihZREo8+SnvQOSUkq7slJmonEpZk/84HArjgiJcQZJVl4MjIOLgnGtiZIhpQ9
tRQeGlroHCoCav7AfhvYmE24HNciONU9Mq0gvwH6Gd9Zk44PclNMOhiZKTqPY3Bp
lU1tDw2rq7qwOZA5hwrwCP11E/iivzpZNIY7opU5tj13ePhJWQdeiVnT+c/V17w8
uxDcsXgmMBhRyvuFYmrKSLM6nCixofXK8Lw7Dff5dT654hOkhN5b3upSLNLbvQzT
PhSFd5TWlTKfsrCNOmMnT7XHz3ulvfzkVQnjQIGrIAnEmKiqyW/hd3YO2iz3+xeL
zsZImFm6XSP2KLOVznqvrJTVCcmPNu+T5DaepNIqCAqe+PBbf291iRV2ro20WaZ7
Ovph3t5BtopM2RpbQYnhtUq0ngxUTGeDLc+R01HJvov4Y5jPVHVgtdR7ws6WX9l4
GjmWrNieEVgYRwfnRM56omLh+Eyd2Uq3v3IBsdwBdOr392mt7Htc8HqO4u7n5Nsg
9yG25nMb2I+1O5e0kgplLYg8VqOzvHLpUPSHoE5k7LZ36UgMCLvZM8chi9lNf2vY
5O2S0pYI1dolXSNFamWCitFwZvwlCZ+8qdUfDEuzhPtIIRltrSzQ4PVBhzr/V4jB
YvXSb0SOKD1o8piiPM4vs8YBWLQC1Bmzvg2CRepIvbu5t3QCoAZ4aTdIe00r/zja
LgQ4n5dLgGiwtoskAZ5w6+Ul74fWHyNH/dIdqI5fzxZaRD5KKPGvHjPW/og6k8mL
mo2smW79KKxk8i5z2c3fUjoOxD+pA7aKbTP1Vv5kQq7UHOa8uc5sWjJaStNzfDL1
I0AqLcXBvhnEhIDOH7FhtmFnrIDNcsuOW45FwlplwJdvN3kP/WgphWE2queNHQm6
cn0mjFCKLCvKb3SjxXaYkIwhyymVGH3MF8nCK9bM6z1Xk7YcZGdqqXkKUVN4VxgV
aXm/XpIFB5DkVdtad9z+xWcnD+HasxqarbS68d7E9PTVJmYg3FdsFKsmUCF8pvNh
tbs68ljh/bgsUIgN224bW14JKiPNfMFIcr4zCQmO/zTF68kuM2Q0Ls1FkuOgl/ds
7G+LwFFX2h2L10wGmmfUzmmqZ2OT/PmQYMqUOtJsLEVenvAr6+BBT1L6HCEHs917
dC8O3VrGJdJLGVtkqNRpPaayKZ6VGOQ5SgzkDM4ZoAPNVWYMUxYt4DPtEL8rOUWl
PaD73e2CLL/qPaH5rzUrKsY5ygctcpu/eK6SKhEHXWIHfrffCr/m1IgTM58LLKxt
JKP2i0mXHnB4KpXB3Je4mD/igUsIlohm08GeT4P03n5XU9f0t0jozaA+bXUYYs9d
Xc6eqjVd/cCduWkuQs7k+fFTx6yf+owbSGQC7WhEMF5AYSEb/vP+A7o1TM8So839
8PwDbGOb0tdn0SJz4o1zkkt6H0mQ5gacKITXrHXz9LCSImAei8Bs9ci0ulAoMqR4
BhK3vgAQsC+tEfYF6nX2N+Tyupma7eUc0jpUwNNRQ6XY+VnUrIhxmDRKfzsBCm9G
BSl/Lcm7yT/FORrOz5RidWE4lGhtmyvR3dBmv43KhYecEu822lwkDsz+ZDgpC8Xj
lPZMEj2Vaky1BIDyJYO0Kbol0oNtGXvsLDFq64F7m6iF0QdGDO45oGyGtGUovJpu
0xZfcuK78eHdrIrua8Ve3L+Y81zgjJ37y1vc5Jp5CKzRvCgE67AJQbBrUyKZd5ls
v+k0iSSldJA/9Rta60lME12S1mXlkcEmuR9ZXc/IlmHYeoW+KMLJbQ8SNM9JUXdO
n3Y21PqtO8TsXJ+yd9y3bPYagbvcG3Ab2OaId4/JwbxbBs7DI0Y5srF9kT47jPl+
qU45Nki6tktkLO238nBt+23+BaIn/tTvhoKO/tMAwiz7f7QAS9/9sV5Nw2yIVYEG
p5MwdY/v6fgtw0LHeNoXmVDE0z33BnSpLlr7oJ9Grm4FLAAzXysFzWU+R+XN79es
5XPQzrbiQAGIyOnIKLiDBTn0sW+CmdZyFWYfANW3gzoWjLIJNBXBoI1WuZccwCZW
WIYQDuTetDprA4W7o0+cSgpyy+bIZdMZcK6xpo/E/IKxMq73giLu7D/rH4fPi9Aq
7UAJKTAB7vCjhgLDJJcBMK8doJFdYHG4kxdMuZ9uLbp/dkiRlHC/PBwsh3BxQuiD
SVqvv+8voKpC8+GpCfXbKnzpva4Hqhqij9spMCna5NhLuIwMQxsv6vlDQa78VtOA
GzndpMGpq0GeheBhcIjBdfOMdE1xoYLj1tdJspZTLV2bh+OHExicjC3dL8D1sYpN
cpwpHtBYET5ONIMz12wQ2SYpcrYuEfodTGZBTgt6otkk04JDBkFkS0FFA2FCBMaz
QLcd2jc2fvrqBCsG79djElpUW1vLvPJpHnlNPeURnusr4pTXiuLWyf1hw4TOxaHj
DrLH2gGN+4mcaDLThZ71O+50aYNDsr2hup0K2nGMfLQoYh3/Kyw959cO9T9tuAW1
4b/QYqILF4ZhhmZhD1pM3tUK8ETzASOEgSPtXBxt99HUFtI9ONVE91TPovyrhHE9
QjCUJPxA/hueaEVWOz7iL1C0j5VNmgXBKvDQhd/bM5kYx6/qoaE4hpjfR/w+pdaC
tMUBtM5KqG36KJ7G8HA3FAFz27Q2VOGNO3EffprbmUsQvaChUnvsfec/l0tEfd5/
l3zmc4qUvzzBYobjy71K7nYPwoR3TczxV0vncvknX3Cs5CVzJxFyn5gP83Y/npyH
vrVhNJzf6eiqGx8XGWjDVgWm5l6r3xoAtsaMiqB9H4SZpOfit5Sc26gxOlmtEe5Q
lSvvT2wN3TFqY/0iRlBoUjCOwCeYkkp8HKBce3Ig8LGq3qkvj/DMJrnduXYTUXcx
SZ60KCc/zzVXTmvbAXGMehfEZokekDBu8l1MLhMBg6/TrKvvMJUKwiijaUuTNhvU
Hsf9FngAuD/wM9JD/ehR11sdzRUMBDMk/UKB2qo4EvvD9tnztN9W/MDYU5EJW45/
5P76zZFfVu7hZmSZ5UB+2Xj3JjoqEIo3XItzI0zYlBDS8MW2orSHloaqrUJnzU+m
q2O3CvuYURoz/GNflkSH8XmG7lnhr9KTOaqfOe4frf5BwJda/7ruItQ3qBIh7VIA
UccR2IzA+/0oq1yFXLkVnI5vSw7g9ZRxv6jKOZ20scxDbcFpuaZkvrObhu1tSZ67
m0aGpwUAwZR4JoWLl6dzSFzjPRAPdjIFItMbxcGoKy3LFDIe/eQKnPNox2bZsI7V
fL9V+owLfulgjo317y+4o5TelC0J5X8ea4mw+oQcRUbOCWrX7zluwlVBEAfL3rjE
AS1y+H9nnwKm6jzO/TSbhEeulreFQVUfE5qbYXKcp5BrBD2Ll7TUHRdIXEZcYWHi
38EFouufuqRshS9U+pfYWX6adgFcYuB3Jxg9VjKMLiNx3q4ZccYmDdmH7djFulh3
DbdPBe99o7XxhAmcEJArDLe8vke2p8joyK/vCJ/NnfNfzP1e6uN1B2iyorr+I5fv
whxByRSDODt5KQwIk3hM2lUNP8VFb+yy4TiYmOh7yA0HMa405J/1ec1tJ+Uslve5
fQmalPigpWskbLex0nc2QaYLwSCt8Tpk25R1eVygyfgPjVdsPayGnOuRYisax2eW
HemHiaTqSdlzqmV0dULF2pwvdhI/5YEvbdH6JUV8Ma3RQmGSRKTbTQH896lcpund
wzIbhRrW/89+eGwn2jf5yR8ZmSm37xNt4CgzVQnekSgusS1aOLjD2zXmf1PvDBF2
QcF7Tb6V7SVkomozHYhKUukNMbJAxkRNoQbccRLQAm1DK74EXHbPGK6sYOMS5PnK
edZsW2+JbbM8EPQMSZTAnSGve0I4Sj4jJ+dt3naJ+vsM7C5N1m60o970XjiPGK5L
9Lzl4SBL80ziTwavw7QKtbn20s5kFii/HL6cfUkZt/nlRMxPihsvZ80eCliFmpa7
TIzqNUytbQRB/uWAyulTWB/sG/5sVVXeSOLzC1ttoCLa0L8ULiS3vguCzLGeni7I
IFX+fM+GbD2IVrIrEjXpPjsP271lK7vpozVCzRrPquXZDhwrIttpu34bT8hjvm2X
WFZlIcE3ToEHCQ4TmOvqXnZYAP1yewHemvuGQ864DTavIvQJabMC08jV6+cMzRyr
Bp/Y+DTGK1v00lqritJYqV/9b7a45gf8KZg0pMNP7AoXltJIxxzZW4Po9x3l7X/G
wAP6oQrLaqgAm8kvN9I9umtLRNqT2KkVFGdehnBvdDter5RjEz2Cbri9UT2l+EHe
xPdQCTUOexjs+yW3BAHPYh/rKkjQvJb9bUKRe32zTvpbXizyUU0oxtCsR/XGaago
VRtGf1w0ha72ifjSrK7dV/7VCSUdIbBWYhI2nsEPSGtP0VXu2DuKOp/hg+VYlswu
UqvSKXRRZ6Az/FVTP4oKda78Nod3F/T5qDduymSs8jwLer9iOM9nZPMqww5/GZma
jeYg05kVd/JGexQegjjeDaK/oKQNQC1afNg8KG7imaN0SVURpL/M0XuEBwHCfPiQ
gFTFrJCMj1whvhkK7sHqDQeOmEEKDGFJ1R8SONFJT0IxX+C9jDCnw/whYGcttYuP
8ANHicFtyoM3cZxvDsbA3EQvhlJPVYmvBNNC8D45ODUsqWM6vhMlaX54snOTfvBV
BtIoUl7+X2nynLaHzI8P9a3824kc3DkLNIx/pM9+lZ+Q+3WTa6/ZLmGCICfLeU5V
KaIzsyM2fIDQWdiYQp2s1oVJec/2cYcRT39EFLXAYVuLLAMlM56pP+3OfREoRNiu
cnEVQ0bymSrSCeFsMju62iHBWTfNwEbbPDJobk7eXq022Hm5ycy3dbk7JuyJ/Ube
ErmsfXgoU4MRT11jT0zNGKqn26x2wY8UTI6eesUP3LDpGxx9R0de/xHanBuOwBUZ
Emtbr57efRkEb67llNTdS16hISyMK/WYMNIxhwUz3/abi1RBWOwqIU/2XqVCmDA1
m3CUmOM9XH/KA1sDnTMpObgXvl8O/et6l4LrJQIg2atglURbzJV1h3waX//WtFe5
u9I6EuVpZpw1T5tb2q6LvUSJkbyImYDcsXcg52H1eqzBqZq/IvVN8tuVco4LFXqN
cYJBUAre/cMBBmC9xgD3ixwk7OfO4SGlSjpfnPxXXZxWkf3m04HHN9ZoYKzAqPQJ
K682v/zAZya1X1E+N4me7ta7lUIAsod8sXULZWBnXGNW8MADabJYuEHOLoplA7uA
9UfmiDuT+G58KzSLTNhSLfEUqQak+Dn1GfDpGdK9xAdDXJO9QML4RfPMqPO7MMwE
SWY/TdRMGw15DSWjPMuG1JXcVLn+rrhKUajYyK2dY6Cfl0LtStkUczaKadmSERpc
QDi5gpxlNsx48X57KJrPAkbNtFEqIKI/qltm45mXKlys+CKxfkh1a9UZJeZPWh8b
7T0bCGLYLXdHBMeUsJLElflC5CxBrXZiI/p7H/ejZjywBfIRLoXoXkfjThxyAhIl
P2jLMe055PThc5XrwO+Z88j/tqGW5HFeAgVL1dJBZ5Plyj69rBnVKD5286j9b2ao
McBJ29cn5k4idCqY5zmO1HI9ErYvR9Dy610xXYMlnU3fSHXqWCinIYbKMf5xnyBF
+fd9dTnnvpHc+9vD+VQcOtLaA4JUxF2G5laHDAW4g6++N8YFmm6iQVHfvcIyuMa7
QYshTm3aRlIiBAvP9TKQC204xzZY5odb0v+njjYQCYUd0AfvEHnCTFzy9gSptEE+
ewO1jVOT9UeGWwWO/KjUD22Ve3Dn2zXck36AZO+cxpm5k87F4LxPCE7/bwEr7z+t
16qpFj97Y+jqFDx5cT2Vpt4My6NpnKiUL+p2yidq2v8svphq2QdOhCpYeqN6PrQj
q3ei9t6bv4Jj/dMf5f49Fgd4ieuPbi2aOGwmtE8RTjNvaZlm8h/3tau3Pam3O9Hf
rPM1y80W+kOa/4VyBCs0OliaCb5t4svRINueqiO2ixps5zBUnQUafOHgRaTuT2u3
2qG0GkKG571PlucRuGeyhFBCt3lE+LMMLToIcPFOwQdkVdwFASZxWK+qt4TIJBZ7
dKWmXCKQLXgT9GWggm68I3CunsBdgvz906LDzkF/JjJHkL79Pb+zwAXx1oI+3jJn
QTOyBMiIhDZo2D3OSm/twsA9MPFV4wHmIKbzUXC4i7AWrYuWb5VvIG8iFuzozMvu
+fK8fCQ/7X7FF8JdrprzfYkwZ3fwfxwkr/8kgi4DdXyFWniIwqI0T2AX9G1xzH1Y
VfVc4CEWJ/WtCXflgo65wETaIwauxoq/wQdT8t89vgcWRhB+Z3XOoVgxV/lKw+Jg
ynf0kPgn7p0F/HlK41D60CCrTra/MfNZX7RPpI9vFDCb1ic6w8uawvcoAi6/7Qbh
bnWqVUadmUPT0CgUyEEkwnR8QiAKdMR+IHdmq9MK+dAvsIAsjbyyzGXG9kvsjl3u
Kub3hiRVoyLZO1KRUGf+EpmtL0n333TecLtjx/wqhoasENILkcjaCsdkRPLdeNS2
C87JUNeUKf4miEfIhLrbp8jj9KBPu0ZR96prGcNFlBeKvaynjJhHON7kwgZnN9+2
yiHx4KaxTkW1iBCOii4qnf94FWUPKmNDDiP7dYpH2bW6Hwl4RR6Gv/ez8X3tGpx8
0VRHWGNglB9h/7CdulnfoK1ycdLbV1/EFcU336Myym0IyTZSL0gAX97e8yX4/b2w
yMPKSV9j8KJqG9g7KDFwpp8hqvLhUmFp3IXeHlKxr4x5MTWFN1YRz0nsWPuf+V5V
lN4UimPWZff5Sfa8XRKj/mJr3LxADzc3R1yC3DNCmYsR+d07yURTl7e3KyCkCEUR
BKFKcFxTQUrBtDeA3mwGW/lps4bNL40G+2sVAzGP221py1BPLpZ5F4znKZJRJe+v
xakclchD5AzWQYY/k2Ef3610A52F8nNO5WThRGf7EW8fdVJgPBdSXft0gYE2uecw
qyWyXTEnpottBqCbTr4faVPV/Y2NgOCY8wrd0nRxHYKmuSDpOeg9ou6DixzngrDK
R58De+nFncxryANzqRW0fY7tSBXRT5MeJ/CvRcBzvGIBA9L2BeoYOi7q38PTzIgX
Vh2oOuLz7I1DZYTDEljWcbxzISTEDxXhh4io4a6ae6jDt1VQ2pMhD6MeD8zpOj5q
3+tzCYfw7lAybp7uZqCl4tuzP2r0zKEaxJ0dccJSi4sN8Y5Q9xHtQ781G7TwRyMW
uM85211XwusAriHVtuMAm/H5XP3itxgHJ3Or2OpBKM/U0Wy6/KReHoRt2WkCC6Su
bU5ASeKGvfEHQ5hjAS8ba4uOq3Foa7CxLtfPxdVcRqHyjYRd/yrYrIyQkoZ8Z8T8
l7fxOU8XSrzJh/xnCZi4u/rMw8+Wf3dpRldjGGNuWAScSn3wQCx/wLKfU8YsYNDj
0xl7UKOY3EM06VsOS2BkL3WIgGmJj2o4IS1CvkKxXU1KTFykgQeU/NVSMW8XuBJV
Ga3x/Pg8PQ/uQXyS9osIgZHlfPcPZH+tJcIWH473ibZqJvrLhKeW1FvRMF52cT5E
ne030U5CEL7j7PT1QS/TGemdJybETCuhK8lk6Kx/sgDAadCBiBkzwzaUJvj2VqhH
xr/+1JZ3qFV896CovOMB7teNkDG9v+ET/QVJ5sjqewl9AROoyvgT+6Tu6dDcgu3P
VNQhh/e+qcb+cHfaZlWIJ9VDloxijYT3SHwmvp4KRaPdQdMVDhM++N0jVCGw/ho3
ILl47Jdz/T3mJHs6AY6NUNOa7AxZY4gEGpq4PAGQv/adX+Xmpip7+kYjpp9jAjk1
C+2aUit3m3XTdF4XrRKJclQahcdGu4Tv4SE4BaoF3eNtM+U2jm0XZ47b6IXXrL3M
+KWTzRB7cbQ1wGfrMJwEKPwoohlymHZ8xyTkYnRHn113Z10DIzgtTAqyxKAon5qg
k2JifmxtK78RcJTCA2IwhwowSfVwlemfgaWwgaL/GVGavDqIuGnnQYjIXCklfgNv
sTJdUU+qG5hD8xa9UXsWJDr2QeKXKm+VodkYPAcNl0eYgx60bV5f9rGvGpbNWdH+
TUIHWEIMIj6wdMnqtI1FqIx1yHsm2lJzLiSyR14gTEpwKo/3C/5450I/hcegYKSB
BCFXIYKsxBzbr/DHso5dcTkzgNl1HY+Znd1VOtyYgmoW59ZlOR3jSmdn6PDaTPL7
z72EwznWlDaUIKG2uy8TQpuqMXoeM3vaAsQsZy6UUkYbTchkFsPXAILu8Qj2DyyR
ciLqJs/LuTra/P/GoSaCn1eEHZVPpIyj6RpEknlUWr7b+xZMO2Uq6cHvz8MztCdX
S4MbQAazrNh5+i7PT249xFt6amAEqm1GQfScBTaiMR2hodn4+NIZ088SU/XIq00m
WuKZr7wZdI0P2PUP5lzezAHLEBei1nCK3dHzXsp0f86gLSIpyeRbjjG96cC6gifP
DaMO4Ccb6/ZN47zFXDPytWy7l7HX18awZq+l/oISaWD2LhUXnpXD04YVK3TGRBOC
4YgSu/o8TcTLvtasMx0SkhcoH79uiuh4g9OAYSzGBABi+jzJeqXiKQnMZfs+Wlkd
KEyvXBPL6K2FdHF8iuPy1ft7OZUmjuXUi0npftD94aOVmGrQLSIlIywNLREfmcYQ
5uqubgfLDC4vRd+usutgp6OXHXqUMDJiZLgkzcucwQJQk3rO6gA08LyKYd0hX6eQ
v3QNOMjNB2J2wPuGA3FKHVfNY+ASyc54gB4RoHx6G2liOP3yPMWqLCTb9bDuby3c
Kuvw74ZSH+2HhCgEavCKPm5e7R5j56wntphB7sRU4h+pHLWoN7eMTmXn8Jpzg1O9
kvBtX5xmUIvKq6JSqXNu3ySsnpfrYVYNRKabZqMUuWRraCOU+XFO7uvlUphzmgyI
MTXlA4buVZqU4My9EY5ZgFvzpnVVV/mCyl6IryUI0s/os30hLW844XgnXBtf37F/
pdMT6gscK2IoW44pkx8Kbc3e8Cph6LMV8KZ6uh9R+K0JppYpjUxFxELxJoQC+zMW
ZuPeNSZ57ykQk4740G3JkRzagv6sqcwKj7F3EI9jDd1iwrXwVH3gOLKgx8eiS6XV
tjvFkhw8D6ZCv6eKKF5JVhOjj6lONgNZDYE05Kaa6lnqKRXmwh4r32AAQTAms62C
IaKcEgpsVO4VKsBovtv0ICf/oRikZhroSi2VaMRauVypPDcLltGSXQhVIJHj+Maw
DIpuxzz7Fb7VdZfjceJBLala8gR5diUmuzrPuWmJFGBehmBVseLWA/Wv3mWB1ke7
lSPkqgLtouyvUuf/EFaHiZYanXC5Lu6KAUQ0tWg58zQRa3O8SxwO/A1Rdt5aLfCZ
+p+f/oZXtgikJP4+HW5oSyxXAC/6C7GVlq3rCfP/C7XhVzOX1/4bkigFBj+myZIu
95o7W8y1Vc1kUdszQF2qCo+31LZcINwBsu28plsIhmyELTDTPDc2bsbjKS6ybSoc
aMFM8UeZDG18pg+LJMxw9GbcfhrQrGoXRo4SX50HIPSJUaxsxQWNsNf+Di7FlLH8
XUeUrx3DEYetAlhZGRY11oxyrvd1cMMefJF2pYOatXXiBtu9Vl1wZrXgH+i9Ve6O
uIBkB9FwWJ2wt620M7EzcT2MPLdwR7VytOzcBhxZPjgdHFgWgvZvGjMio6+ohjfy
a11GSYB1smlHseqaYy7/ODa+UeOaUdE8TpECA89dcI7O6Ddc8uN9eqDssdozGxne
Ssai/4ECFKznAVh1MAJm31cPvmgYuXVCskFJXDQJbJ8KjOFmxNBwOkJ8YJb03rKL
qDD9J/L8l5C28K5i7fTA9KNsr9sUBp7yd1UqzyZHvbICD7tiHQimfviqPgYoTIDS
JJ/r1W1fMuqvw+lPyCWw7hjLcu0QNMye2P8uTbe7OEqTaweDE6tJxi8xcDPrKZjk
QsrjnJ2ZNQDxGZbfuYAJl4hrVly9jgURBV2khJvu3XsuX7pdyVkdJGvujxPL7wAv
+h2k2lzpnpMxK0vy+AmiYtWI5XIs0D/Clw6prwjCm2UgGShyJKEFNj/R0f2UM9tP
VKgkKeHKSv15RiLw5DzXesLIiiP+eQwLhCociS2I5hJCnjRry5MriUrDfj76iEut
en82fJe/13wmppTz+TPIZNF5k/OUMdaonJUm9x5w+88WggN+mQxF7Cg4sW0OizJH
1fri10YWmBJtJvXTTbg6SZ2p1IW9+8v2paWW3DkWHVmCTiyHGbRIKrvohTjLt7SJ
Z9c9BULXu7SOSVjPxkv/Szc1VCtRSqHnnDo7SXMgSGjJZ7MLo6iDwryu7hVz7+hE
rlX8AX7S2GwWhbI/0nABhZZwdFDOjTId7mgHN4UPmcip4Geegs+zuwBVK1H5YrT3
bOY6yuoR64ArKGVXgvYff4fJAtfvS5a1dDmX98vHGzGb6L6R9jpkhjDfg7T/pTFf
hvNTFAJ6d7yDkePNb7pqFPHJmPQe21DUZrXj7Vid0cxE5yaYvskxAYOdOkBCJTiI
TH2PY2m9RyKYzNoeRxQ3StF8cyf2Kbu8lTaopWcGDaZrk72TIJMFJwTiXHn7bi8V
emcoh3zNoeWOzbCrU6nPubFUd/RSf5bB5LnMGdeEVMfIkoGzTztUS4xObkAgbBv7
eJ7zchhFQIq9ByQKxwyePXmx2aKqSwlIXfos0IPdA7a7zfI16AiFqUyOuk5DauK1
+NJLL8sNOkYoG7UXSdatJpifK54KoSaZFdsofdeyD1h5hlPA5Ok+QZnVzm1EiJJO
d7dPOQrPyuTCUcE6S++4omA74VkZoIfqpNxllCTVGHjGn5otSbu6169x2CFgZA1I
Bhog+Vy+XeUsUZY7Okw7+Z0dK/K3kl/3nWmvIrlr9LUkrLLgxcQHvqkK8ShoOerq
DsB+lBgau9enZjK155ENEpP2TVNrYbyS8zIni+rL9P+TvlUd8sM1jLLduHZlK6f1
cO/4PC4rxrLKnRdZwx7To+PdxfdpOQ0iTbtwkXmnzpyol//oKTPsFVVkoUlJ7aDX
aCDvHXbGpOtlCAPu5Ire4B1SA3JyeO/eqDzd12MXGgE9vhgGxPy5SKwR7a0xAREm
eOsHv/T6vUz92wUUUHCwvukgoePqVb3D7O6sZDAu3ZiYXa3FbxW31vKewHRqtU7G
uEEI02Fb9wlkMwq3XWLWYNX1IZ97QlKmIWs1D0eguMy+3Zp3V1vIj+JJtFvFYtUR
68wR8tz9piDGQWPmfnW4p/nBFDFAfWWiAtYaa/0UfTsnfnIIR/zqKzeoNGlNLFC+
a7RilyO+/p3b50MZsZuqLpIsLzvc+gmH/NukaQTtV1Cs4QH83qYY6jd5yagkr0L4
yNJJArKRavuEkp+Gjrh9Xk/yK6pAbwQks64WCJiCZjMw2Q6pc7xfCkeIbcgSoeE6
XHLpH5ul2tAGB93v4yMzDOMeXCJa9t/I7fXLQ5axpV54DeCxb91yZQ80BXx3fcwn
vABzZM16R/x09AL+x7VIKTvnuTuywbm/cnWO5ryYaZ0oB441OEobeT68kX8j19+0
YVJcilI5mvSWfv6BO3/CKFpeky6DNSf+H/+PkbkjXdR2i6UUGuh8X5KCoqMx0NZa
WN2PXEvC8xH8NdDR2VWbzZrR5NH5Hkla6xxppFrTRLhe4JPXFEQ0feHIkMsPtHfX
V0hPyGWQKS7CTeFsNyGQHf1wchLS04nHZSwuoesXF4z2ktaIYXeAjEOrOFok6txS
ybR9lUHBuUv0YnsISZmDkFngYeyO//PlCeVIsdYi/TnmzFMxEdu9BOhPyKnUUDPN
LhzyHEbEx13zpB9uC/rIQ+cA9yJPKx9rQUOCcD4HlJulHQR5ny3LhRRjXMhFBlKd
uyVjTmVUygVWMLnMrrRCM3v+88OF7Y72kQ/aaduuWJk/jVLe4cAln/t5Gxnp0giE
NdHYRlVqHuIxpudz+PUYbsqG6mp3KrHGJmGI+jrsVLyk+BatOH3Lccoctg5f+PzZ
8WxqWKZKU61Q+hkbAI413CwQ+0aVCrdv6vtoNFNL4BM6fY7HvSje3z7H0twGcocN
AOnIQQqG9Cu061gwj2RhUHfNw3AdEiI29tfpmfD1FQEJ9IP+Q134MVArQNQyw3eK
jlTJ3M++nzs2Z2fq6Ft+hmRgZAxgi8OIQiYZRAWrOm7CzBVKJnwzt/pesOrFBTb5
E0k/EJRE4XIZJRKyiB9+yR2R5DuS2G0JHnHQzcweC/NuX87JVitsdczcPe+BNxr5
yVPkUygZvaB/BBXxAJp0ZAznXrPMXMRVhs+ry0BoaYEmXCO0xc9ZbZBD/cYpzg/H
K18+1DfUA2DJi/wWis3D3krFZEmnVO2AAEw6le5uG7Bt8dYFtHg9AlbwXgDN8It5
4PwqNaqC8uSY25QrA2+YhabXPuAWVJopOKEfo1hayqGtwLmM61To5dA/y9trOs6v
MGNc6wxh990p4q1hg0JdqAMGidAfdMESuEBiw1ee/x3XiHuiVUreXJWdyqObIYA6
EdcSYy4PohR9g7UZ2EgBIqFIW7iAa888kFIP1L1RMX+JX9T4vWhPj8CNBzSAy/bH
DaAzkWOps70guk6tyJnNrGb+D3Vcu4KCEy/jeUK2sQZtZsi2lhE7j4XaTrRnowTr
rZCeUdU9deUF7UuFoypuWhbZh0FYAaN3j2k1vF4X1Neg2IekTJJQD6XJ3w4F3tWA
uHF/X5vrtdKRTbskvBAdDSszEP4QFT5KJmbuKZ8jpvuqnvBR01uvRmmncCg4Mqq2
6ZY+WNNrvRqO9FK1E7l6YqNjebdR8p9K55itnV6eXCJ2NATjdrRc9Qx/M1bVgNfM
G4ZE/EIZpT0VRCsQlxNX09QKFNeyMglMciR1ODJPBPiwMl2NvohvIDPd3FisqZu1
Lk0Naf/4mPJGJgCiqC8StSS3gePiRG3SDchRNX62E52TvsS+HKVzo1GzHB/hpOFh
A+3PxXUSlyoCaXVPIdYBm7A8eMlYWDrsuL6weRRe2SGRyY4pQXPofZ1Y/a6t15h4
s4ElTbqmdIN+VbSYMOPg3hdp4lx7qNZ6u/2bpD44xUw6U7WG9ZtuRJ2xF5qsIMS3
NKcJB/+AAiSfY9keaOaT6XepA2L2LW7KkgkqzU7NHp6bUzav/aJBv4CXzQWSV85Z
c3/zpm01kIAkkqMgRxJ9SPR/88MSs/6aRqfV/DqDaOBgkt/dxYPnnxs+n7jwDUkX
4c/nULERK5hAyrTfcKgbp5QKBkKoN2E7v3ubJnp9kGoxkOOSES2BOzHvCq4+A1Py
etIsw1a+0iOzoJIUuijMaUNxOWD81QJbH/7rSMZ6Ypa8Q7GhMRAggDR2+tm9rRqP
K+I8LBOu6Wj7yeTzHd2T4sUdcnFlgjw5gS9dhTvSZ6A4blEeHl2OcbiO1mIZN7xE
0oZ7m39sTrLr4J3S/y19c604bf8baC1KKrtNfODfRFpAgmEcBivKETJTKlmA+ZDM
hCHeMbVP6X2vJUkRYcUG2n7B5CWQ8Avy05Lf/N8yoiAk24S9UuUY4miIwATLXPfv
AdaJsTevnu9rmoJFzz8ElDrCHZm6QmqgyX+EJB+FMD4aeBzH34uEAKIdmlCGYySn
l+czLQZ7CEOL3WawcgKx3KjSS93hDrDSSgf6SFuSYZc/WEDSThSGaoaqMIBQYRW9
rmWhLSbbWUD0vCDyEUf23IPBSUVFxUztzl8hNSttuMpglE5lTbkZX37S9KgXhLI0
BuZatS5YgY+E4nahJzxqr00GtgaDaEpjfgmF2O7gpPxgMkmoq/VX7+7E0CDTD4yJ
zGUcQnQmaxzvAdDgGflQ9i9FWFplaO6p+jvCAYynjIQ/VJXSkWZhKIBiLZ8oE1fj
GPAyI0cKFONNid+kj4wuBQvmt8DGEn/c6VVVplLQXuWDtjnQVxkoPFtdRAESZHQn
LHmd+UKHj+6Ps6UaDOZfTDynw+rib+2Wvq7Ske9YZfK0hGutCe2lqU3IRndhIBQm
LRRKjYxjtlYVtXbKbm0QgtlQP/ppzdrQQF3Q9hoYds3safPY7iio8wYU3oTu4M01
+Bku+NUqsywAPRkcnt3KgjYYGdhU2hPhS8RXCeZA53ZZL+Jk++Yaxuj1TThDSpAJ
m2+mav+UhesTqwGSqC9pNfOs/I2pP98TCQZUkB/RjSpdOjPhfW67pzLdZqa+2cYO
YvVUkaX+6zOTj4sk/eLENs7nEeF2GXstKj1+aaipRcNnXVUjjgtgpgTDznZt05jY
czoccf023pkyzaz7wFbWpDpKRMDXlzJ0zJdBBeu5Yn7KXxJtIVLQHo/zzbendei+
lFoUHu80qhdSsuhtG4o5XhHxZOnUeI1f399LvHFji5gd4xMNoja0sg5VnbSypvoh
CA3ysWZDHqRVlNv23H4FBlX9/uihmvItottDWykQ4DkAhyIG2gm5TADd1gj9jRwD
JKjv53I8rAN/wlTtU9880l/H4PU+3FABJAk8DyH4Ix8oheZ1N2cWRKGDSihb23Mo
1ToAaLKcVS8Do3uOWGxSM116xgS5djsvEK+y0OxvuhUlj3dhEcaTIKKkNLsCocGF
7ZryF4M7jMh/c1ujePkUg8cPI7jUoZJ5RFKZ0IXaXsiljZMoPDxYzWNobHRQCmq8
1PsrgO7MLuPTS9n7o7LV8ve60Q923nFIQ4ZCraWGXBjXmUW62h8lXAz+8ZsuSnsN
fL+FqUbfiMi2j1W/7c1CN6/f65GfTsmvcHPvbgDk4OOe+iHsXx0t9agORIf3WL4C
wqFaSqc9Kmiad1Pc/9hTJjxkFUKVUwkP4q0EHJznsxsGHWYqa7EVmr/KA00ijuLj
7Zf/KGIpmHjsYcv3rU4EEdskpixU1I9Ce4ZN2RlS2G41S6+Uo9t4WIW/UazrV+9i
l0uKAtTWESqIvBjw+f3GUNg3Q87rI4ncHQLqUSL9aS4eNAkuf/C6XN9OFs0NuCrz
RlgvcqmCtH085ZHJAh1Ufu9khEI6PkMzSzUMUrK4sEko1CO2HPYIREE9UXtEZHfT
wyPdCPSWJqwKpXsK2m+wOjEACgpS+GNERdhSZZHOheypsyFqzHVlU0ON0lz7ksZM
eWokxGTD7v09h4cv7Ra12PJI+3RhVZnsKjnTiz+L/6/c5qZRdgtQgVknzGPCfgPt
h4Z6ilV0WrzPMuL8mjOGDEydJp9SOAvra8gfMJuaglKQJivy6ZzCmbsJcIYAe/jQ
Vebm/Tl209r3eOAjzg/0pK/fAqDbzVZiJYf9ncsa/1zg3+j+eZ1KzRNxnBVf3jx5
u7ZN37NnjZRpAhmzSmUAbnZc5AAG+ZhbZ/jEFaIjPe1hebRCtulLEUyJqZ+FGZtb
IeCVTRxrcpZdMmQo9+BGc1pWEkzC5cU4WlMBwatu9CHKBsSuAH/DhE4UF5JlChH6
vYUX5buFTTDfWoJP1LE1M60Q1EAW7hMW5RrpZP3z8ikpNI7RmpmmucQ4fEpxHTsA
5n1KYytzaJcMV4Ew7K3RtStxL5zHfuksH+VM4pOpeksSozMjFTyw1wZelXXmgU2S
b1O3dB7OVu5tTxYLsdSY2KNVBl7zwUTuNT2IgBg+dXI0f+NF4b8faoFF4SYjtVUY
jprYDYis1DqRHY/ZENRSU6/gYUUpjEthUXfDaT+MCGUiVXj4tYzlOQRDrxtWg8tl
dj6EEFAs1dLNY5Wq4BoH7mYh5aYAuIluqRpShtCD/zpSX7GaGCSbfZW5mRI6bK3f
nopP7a4a39n3s8utZ7TAd0Gvv0ZMvieIiHnTIy61NMnV/B04mVgq44hn45zanWnJ
Tu9UlCqG2Ar1Wa76GKp32vRmcD9GSYkAioCU+1+H167KX00AxGAEZvJz9qUZs/GH
5L21Ol/KfgKwDXEk3iI2TjcRR243bML8nXYYjNvj5Et5gKPtwfCerO9JzVr4HcXi
MhWFQgT0MfWb2Xf4Y9ZVBTX2IBxkxkmoUKWMGpZFT/qow/046j0w3kn74jTKR9AI
3BozvOcVLpjGQcVK6kEJZP7TcKH1SHpem19zWyJboShf0coSURopwiafm43IbHiY
+R0rdd+jsRTdsVEddbWyLbisAEHe0ceMIeXIrco8/bT73YA2ZdESk2aiBcvr8Jpq
lQcG61Zg36/WctYV4TmCwTCpALeGuJrK82jXN2n1D+gKwHesCIiN3LTU0LwyQviS
6VQ0855mSuPPPXpmXfbYILRFoR5uxp5Bc6ArEq3bHWbcG1LpoT2cCiAzSkdlaEQ0
Igr78rrdB8y8h0hZ6Qg6upzHTMIqpmXjnmkNQFbZ+KoeI9hBwPkDMlU7NgHBJmfY
4YL/kkxUBD55s6iKFy8h+jcTk6HZwYG7pTvnNQKApTFVQn89wbC1VAhZZuaehc1M
oWuiCntsIcDwYk0pI+U3LNvFh6Bb7Nq9vPy5nyxwwbWpGmPUrT79l4HZEz3/eqHl
X4YsktVY2lNa4GrEKicmFo4hV/Vww8nH53CCSktRWSjazkXMoyAY+SCipx/A8xVw
2t/aFJu1H0VnT6EFZUb6Ur/dFJlPUGYqgqQ8rOdC21u3OFQBY7yypzFM3C6d8QMz
1uUqo9U2pMgnUyPipn2qOm5bCSArqgIQ/jQg6YErngnaviqe9BYbNO7UjbZd2jO/
xgYmvVPZ6cmJA2SBYMqKhGNGFpJSZrecAKQKcn0SWSHlZAFi8U4uSfOxY7r+dk+s
A5Fdy87vAD/0zqpjkRD2VX+yjvKtU/T25jc67f7YJAnJ+e+B6mOqKwkpYpkKom4p
GBPlg5HbVTWjjAwrkiznVrDGxwdCXA9c16/vBzW+CXhLDc30GnH83VKUtj6ntcH6
bo8CIbsvbsNhzZLdXD81sp2ooZiH8W3m+X+rkQOdWXxchOllDeKUY973QpJhAkyv
trTdWH/CLeyxMDaOyD6ikLj2CCOAukXg/QEQdgFrCC2dnO9sXNAwTzGrB9AOAh9X
9I7IbCMvcOWDcfaFwycNsuoPHamqcF9q9hUTud0nSs1YuFIvi09mDIE+wSUD5xU1
h4OB8+xkQjnmtU3SQAtbRyHFOJTRGYxvWv5WGiAJKmNfgmPFX1zKqv3JYENO+QrY
k6T3LSxK7oQ3CobbMSpzaKTiaZ2sQ7C6VdeCppCwL1FlKRBmvAWuu+s5lMSdTGyL
dTwD9EJF1X+km25VuxzVjCWv2DX+VsBVM3V3/tiow7rcj4GxubTf8V9GeqCxNF9d
dSo3jzthg1n/h5+r424KlENNMsAudMatBNOriUK9tVI3ZDveYd1k9ELreE+3/J2h
MiYmTHvGddIO7+a04wYg6PD+x1+PWQlpmX/vPmBT10VM3rDsTrg3AX/Shd6FmzKG
qVixXgVb99glct5luTiX5fEi75F0YOmfosLWErGgyO347X/pPRzEtBowjhf2D+Jg
HRpk3ZBKqrnPi/LGZQ7u8fUugESZQnXEk+gnFPPill5VGKQo134y/bfb6FyX7zjj
3MghFBAKYgaI0dqFeTezyOw8KlP4xZbcgnMqugnpOxFtexaQUL/XAa0SVkLLOUzx
p0C+kPjJVXDFc4rFgYDO3SjvumZcKO9wglOep8x/JfOGCca74tPaEXyRrLHO5b43
tN+YPUf+NRxKtPGbY/AyMxpDAHf9c9FzbMeo0DMzgLfJXbx47bvafieemBq2mbLP
JTYvyo0nci7fnrZSk+Nas4nHE4O6foe9wg9/XK9ydHcD8Wk1+WyXim3ajy9B66RE
9UJyxwYL8GfEPyVno32N5+udmw+iJhBkwyA62fnhc3xWSIsgPjSG+QcIsnwRUOX0
iSDfCCDmGBMjj9GIV0NNWlVj4U4Dlae2SU/VV3vxwAQ1bTAXMr3r/JN2hRB8QyzU
+fogfvlKL+PjTLqcyxttNxptxV1UI5YSxg5zbqA0Vib6PjtrlGWlCvbIwRCwhM0X
5XgzxdQzqMaxyUafS8XNKUwZKc6kfuW+6sm7Mqch7RqF11BpbmU+uT4IJFoSprjp
vCiW0UgL2bIplt/D0dXEMWHZC9h0h7DMbBK/2MPOdgdHiSBV4hqI1suIOsK/3cAp
WV5k+5wTt1COvryvd8lKSAZ5OGfH2ay+f9B0Lzng4Y1n/8Pr7Q6Ws99Bvy+d/wL5
nMG5nB9qcCNI5LiO2qlHoqVgRIO5Rfmr3JXNYKVdV/lLavPxGsBF++B7nz1MEIxL
borega6EGeZC7OrpRP+G35NKipWN/bqlOO4QzTLzoi8ODhzdENym5JOWPF7gYHKZ
LzHGZYdCUVXuht+G1kpF5t+ZwTG6hcP4tI9LrPDLvls4AGdgjTubeU9iL5b1a151
DfEQEvWaT3eL7+ADwIspaQnlevW+GizTpzA4L+y+slyLrRVG+DAWlSKptlnxnd17
3RnkQ+vl5YbP3d3SOuGlRwDKO7xFbLED3grKVRhZys2qYR+9u0ttgu7YvJML1N0x
6VwuLgxoeTKzhuGs0oZX3cuYUxA29ZFvsUOrIlw4PKnPHHbh7xkMgCjsBJxm5YVZ
Ryh3BzRAEP5aJT+fvfMy9GNfLXFFElygQ/YdsLKfuL5mFNjeexrs0USCpA46fWzs
7r6WTEBZet12KJ7NJ7hK376InZGH1xfgmZEAMJVxJldIRQOtqcOENpE7Nnt+aydy
AuSKpietUKoS3zv0Ouvc+AGD0OPxhtNN+xldaRnaUTYYnQaUmYkW0XIkoPaIkBCL
VDBGkWcCwuQ3tKzVV45uptsApcVZbJDiS/FpXKRDKZwyIHW2tutZBk5fcv4K0mi0
hHzcprpZ9IiFx0dcnuBr4PAH429Bj/mTvIgPISgEwkN1U71C0XbfCDmp9NvdHtxd
jBTHEX9fsrLYQ9UEQ/r2811nMZ8YHf28kcFcWWjwGBA+HaGGJI3A7hBVRfP4PIxC
UubO/9mKIsgfCDTw4XsMV6Ap7qW4UEW6j9VSOj3YQIdVUH2urQL2pAZFlboDd3pg
nlV2bRxUsk645FB72Rlohk7kA4HwngNi91/nBr3CBvM3rBMDI8XbhpDV3zwrl2GZ
/YWHzzMLv3886U74b2pJ/G3YBomdKL/K2F169mUrK/sysXhEa9GKxsFJui+VXQpU
2KvRcl9Al8pmXbTUEHSPaoZj9tE+AmTpdY5oN0PyGkiUElL6o66JDFuxYIxExrsx
sswis/bk+rNL3xhaAeja83NqiePgbbsVhx0N3nLpdFhYVb2TAD2JIidZB9uR4n2r
1cMO1OfSRnO1HaUHrdqKxS+ZpLDzMzbY6DfaQmTJH4+nkIym6wTjxyuygFi9tID3
HNX07WCSCGdSGBjAyG1AiU7eT36TKBDZsetL4NR5CGLcKpKY8UWVzUDtWk8cLZH/
zdqW8konOuVnZDGdbEt4hzsJqntjjTCOKJSn3RiXwd6mLl4pkcq0llvSMPsffXx8
sSBUhm8807IzMnjgRQcfTzIst2sh0KglVaapwD1e8jQJ0uTiiguZcOj2POd21lZG
IZsRzJgxj74SdYoTKBeMtAv6CM5CejIyq15FXVcEUXPo0ohuNC1mHsvG1rA1Fyqd
HtqqoAXaaR54p6/a32kXfAPm963Yxu9vDdP/3Fwz+XrdMiGqL9rXT5mPnbKiSrsc
f74CgDCo0Zm301UpKwOq524zhX9+NOF+1gh6/yVL879SiGTFYIa+C4qsF1BrDl1Y
Hc1Rtj2xNHzww3CcXCvmjQ9e9Q6uDbX/1Qxp6ZSqdMX/yOWu2fGeSAkxGM4T9g8w
NcOrlGmzeHwvOS1zqhI3dFiENhtJvQMkUt+1vxZfv6w49dnRDUKTMa/FJqc6I/BS
PM85R+8lSfj3MPL2SngsVPAEax62aU9S5TgEz3+UqZd6JzrfEztuTo23cLFQgcXk
RMJ20fncdBWQyw/7B6bWTwsKURVX6s2Gkfw5xNjef5YQrFMHo8QetNF14b1tfvuP
w7+vivPFLbmX3zLmFuoxiBrO//RwnhVAnh+QHSKI6g1fGVaFjYU2AKNewiySwDra
D/9o+kErcY8otgMjEou0linkSueeijGB7R/bsaaWWTlRh1U8yi/EnVfpnHLOVF6Z
LfsYmilns/ZQP5rTwGv1SSiNK49KgMmmWpAo7K8S3XC8hDfOe7zpHuRkayIDAITO
XQ2rkKke9EcT5IiF7KYUjehlnuqyTavv+tXQsaXkgHSpmYVC67Ih8k9dnpF0Ziqx
4+nmvq38bdRbhctnn9l7EiFZbels6wy9cAjoXIUDMW38MWbMRj668vJ6uq2XdLfY
QgYeoqZExBGHDrK0lHp7lcykQamN2kmbsg6WarCnQMu/HljETBkCpttSQTWrEy4E
cSQpj3cXF2cRDk+EhE5zQQ3rSt1nF2uUFi0CEtQY21OhB1p1WkfAP5IPiklKCY/D
U+PmUzERoy9SsD06zriBeb0I/MN1bK5u+76NBvcDRwHS18Eh0KHeb+2srnai85Fe
4SzyBe41My1vbM444MkFCq8xqwUKo0omLuCkRHzjgzXVCYhzk8cx6kvycgzPpyLA
xerL/1QcqtXV163AQh29uBzPp5/2lDz2LuVvcAGQrNTuR0JUHgzSKrTmsI1shMhC
lssM9s6kBdy1zGXtR9Xw7aBjroTI9SyTaMPcvdo+K0evGk2BwHrsDaiNpUeCHa5t
FfpLVK0wqagp6RD9G9jsUoteMVNvCZeZLhUOBKr8RwcX3nfKXaL4MPdrpcqjvNrJ
pmlw+KkSiohESwBmvEKXDMLQJQN8Qm4izysPI5Q9E8WrNFdgiMhBGd93YfmNPYSb
Hq0n9K4yRfNPyOyfX4TmUmyZYFW9gIeB101pEwN9Kq5voplYpOsmn7GHREaLwC0R
yh9uTtEsKBi7iwYH85CHobQQ2EkiRjnm4/zvEMzchZrhhJKrnHeHHSXsg72Rv3a5
Ja3KaNWgIV/g19AaYopBdUpfuJ132rwN4bAaz4Pwwh6LiGpLNqXkeEo5KpiRRWzg
EDANwGw4qsvwAqqJc7JokplFj0jqgePu0qdCYYAcA2FKpoIXTpDsPkOIZwQvzEUD
M2Kn9lTZxlbq+yx82bmDr2Pt4y1r2AiQNorLVGicus3+glOz+r2IsTXM09R60MnB
QCcsCrsHvuwAPK+erwSWEeX3Oa7pKwljmYn9clsGakdhtsdkB26TRlOJBDxupGqy
5aolSWK1WGi6UHuztm2PEDayXkt6w3L03JThKWP0oVyDEY1NErXVjqOUEBoa2z8C
DOmxN+zMfB/el7PVu5Tb02SmBxLYJSK3wvzlgRQsIn8PmDal9ad1wf2okKCPdGiT
haQP/9B4FKGQtW7K/umpAXwdZxyszq9UX0iAzoDjlqymsJPsX+Y8zZJEF3Fzr1RF
hRFc4yBh4yN1M6pDpTj7yRlAy1UWkGWPJa06LsALaefFw6A2PxUUEAJCHjGdYvR7
0XJOtIkwHyfTSQWiNur1YfhIUjMFN1Aen6SeuHjluXLXFBxT/Oo3gS6jBzli08Y1
q8nrG5rN89yey+1QYx1ASAa5SjzyOxJh1A/5C212u9N7DT/rn1j+d0jinPxyd8oA
YSLoTRHPKpDhgBb4MLwxxepkZo+JxKHUp0BWP3Dret6dZOZxgaauwNo/yquOW7BX
59iQrpJmWSSFDgQKsy2/Fu7w6SnI89s9vrFBPJ5NIT7EyBxzP11sWqoVrjZZOoNj
dAajKf+4IKyWAf1RKmbA7FQs2R4gYUUnN8N1dlOyt0kTjPLVUmckKMqhgJ1wc2tv
NEdvYN9holWohUAC5EL652yUAkoYH7Uz+6dxeeeYjwAkDAaNHgKu34eSbIAOV5xi
p0TFJbgkouWnBaHJyEB+A4kBD1k1hKfk5mLR2q5hkEBaICFchVVsDYDWhgGT7w1H
0EUCFZFRiud6bTcO/JU8r84ke71leS3HyduYQ6IyUNJetIE4eOeMzN17R5b/VYo6
a/5MxVaz6lmAz0es8QQjD1GK/Av764CjSXFI2CgUZcpYRRi9CbaYeXinAlMsgl4a
lanmkeXkB7Ug4KmQvaxFkhRfUKdhr3BOJ5d57VliqGfelX3waXv+qluyzdgYdi+g
f1AS1iQCJsjOiZ2UwVTWe85i2JhAjFnu6OdYDsKDW80k4VxAubkYCzwGDSTi8mmo
j5Y9I1v53tfJvozm1IjoiB5O1/HofryBEKAt15IUf5n190JEAWE47/5ALex9NFVY
zCu3GkQGRw9ZHHHZ1l64m8JUJXLmBYshRzDEk4bbqjlYAENbs3HADeV9c16UXrCJ
MbNDyT7OnhVukZNoRbVFi/roC8e6cnQVegS+df7ClK1Tav0Ln0E5M59zSx2VDqhH
Zd7+ANYqNh1fevdEbeS7fIcWUsT63Y6bFut7qhxPpMbhyirc/cJ1oNWhKssjiU8O
k/6VrIMRHTzyq/leQhEkI5MM+RCHHmlwEJ6qEmYbMTgI+Xvrtr1xuT+2C8Zh36xM
lUGGMPNDvc5oLbTT2qwjEaitjsMtiyhKyixUahvUfQEsOHDzEHyinO6rKKWNUMJo
6+rL98zqXRY68rZuwNEAjGbukbgTQNHB6QgZm3cw9mcJ5CoUBiFjt+4YEBdA95fQ
v8Ffnaj7zmCqxtQgz8PtLDuX9G490JxvIv2sv8ZoCV3sWQKdz/Dycn+Qn40mKozR
l+09+9SbOK4uCvbZ/3uPtDUMVCvCYFaCFMizJZY9X0wRcqUHGAfDCZEiCChtp7Ad
MDrgQ5VlkHAGT50POhoHPz8OFGbusNcenx48IFGIvymiTYbG1B7cmiwvWe+y+4EJ
FsHhZK7SF5sSytuhk+DjZPHzum95GYMe8wurhPdXmRP6QyqVahfkKGwtkHIQ63sK
4Hts9yyDR9TCQPEOnPmO5lqaCQwKaNPEal2Xza57qIS+lWrphA4WG/64Q40XJvDg
A6KtSMebJ+wUMNGEUUXGQzmJ9e0KTzTrJQPFuUr5cBNVloqR8fZD+i46IKN6KZOs
ensaGZSWM5RQMfRR2NZjg28ZTXNWuFKnbhDCjflikX6qMJBBoxe41Foxf2Bue5Sf
sAHz2wqNZl1rEiMpvVH2OTBKkAyPdqOwKdlbCMtDkSmBwkRNyn4o5o61YdYxHOUM
zGEgpLzlgPyhPp5hGJK7ekkJ7X+rmw9oEl2pPc+X6UoXHgNnE/v2y8Efk0di2Kq/
rPVhy/ty8HbiA72i1o5xZcJiKXz36gS6QhcG3atUFh5NdRXhJvkCk1P++x8hDl0/
ojgQKbywRyWxquTDfEoo8o0MaYW7nIHh7ybcG5P7vSaTNGHw3zIyaV9o0xUCoGHJ
sbSA9TjEpiBifz02UEq9QIEdeiG6rtR76sL0CCd7N53MzJnNocCvMjBFvB8Iqpjo
ul/1ccwRAIZ+A0x3AmO7QfFI9khTnKF6rWEsgIR7d+HBp//Fcn4BNKZDeevvZfOc
2mPPK6WVHknnJgO3h41X6ah/gmnWZOl1ky+H1hNErP/zFSoF3CNWSkdtroinnhXS
ixof9ftOjbj4w55z1ivRjEcpJc7mmwgF8IzL5S4u1aaYh561nZ+BOww8JTjidcUj
FY9h6dRecvBA31/I0fvJ1M7PMMZe9B0hEfjnIgdt72NNzeZPj4wNX1iYV4O3mra7
RGMMbTFRwbDFxN5AMgXsGyclJQdjv7YGGS57tXvLfZkBqUOC2YknhEiYw6L30jAB
tnU6MU6sbV04Xlxg+k9bvnOR5+zIL3MpsawQFQQ8MGx21RSwY6a1gCSIxNOOfNqf
4AiokZxw5EC+/PApFc4aEy2Wr+ZdP+3xcrEdW1DgocAoUa7ZBkQ/xmxfgPpnNokY
9DrSgQpSVqsVdBELOsvmmjNnou6FEDS6EkwqCUjWMjanN92645HGP9oDSzs/P0PX
VVKvH3y6r8PPR58TuyhTuNOOjOFWGdY+8QRlXeVYJUlR1RYugZcRbxrYvlPcD5wg
ZkI+MgDhWFaRjx2TObLqjLMK4xQTDb0j3F77FNOLTnfc1fo3vMkMNn6vI8vDo9xb
SZ4NxH88GH3Qno95S7tEt4Rq40VXj8i85q99B5Vz4QQs3D+t54M90dfxdMXEiEJl
O4Ke7Xp0B5/Qvd7XheXhtB5X0vaQtE3uHQTy6Equt86nqgghM8ckiP0gc8roZ3JJ
S3UbbEYtXGl29Zeoc83cHjBuswgQYzWorq1wWLdDM5yK6gvVtnBkVMz4yUTpdXf9
/S42vbQ64jNPjjM5cY30/QPMcneGPMQE9szc4GLyLmSZqs0gqgCwXcvUu3JSxZ7I
US7NXe1ru9mXwPnU06Bef/Pwg04OEja2rRw8CbFrh71IP0zZKJAYl/yW4GWz7ZR+
n7O9hhBZccL+FLIN5zigpeZ3inPLoek6TNzl45mzg2Znbn6eQc6AnROhrn9BdJSj
vxVa8d5dSjCn0VltfY2NY0C4IZVLhjhUmislYUOS6C/nW/tCU1E+z59/d+j6qrJp
PT/rpQj2zpYD9mgHo5PMZdlkxqfaljiQE/C51sT3QczjeT6NiEQbqEOVXUN6bjkL
S8qUTZ+XcL+A0xZGUoF9eJlHeg7Z15XGBWMZkrpifTgHvWfkrLVru4QCf3V+mY/U
khKMXJTZ7P2+ZG62+OX9z2SZIMohEhfmtU5oMSXAt/FLleEM6zvuX0eJz/mtb1rX
LUpE+fPDdmEN0uDGaDN1aeUOKzdxaHrSSb9L05or+WmopSdJ9Hjj9prWJQEj82PE
kJrxejHAHEFGQR7a9wUq15A9EkkOTD4t+xnBVUCQCRGpzbAD/qyo4UUtBPBIZOe6
oSm3DqyIcsKDjtKL905WYhrz6yvdUJaAAIGx5ZmSX0RFZn9CPx+rWGQAkYNt60F0
BidP5canBbRPYcdqruFwehT3KJkHWICz0BFug7YKfiQluKqnGet3L3dP+OQrJNSU
4KOMTCDAFkVd5tiSYUh6fAGaHctDmpBITqTHnsP6n0RZVwjS22XGLzNCPuZfF0O0
RmQhaQXsc1BFef4XMkwYQgEccRD2cXuBdsHnEVZ3qhDq33b6UVcl6KxDCAIZrp8s
bfjXz7+iIVBDIsQ9HFYceTZvzC14s5C2gPJ5dbrv6NBVqHO6q1XGWMOMW561AORb
KhF57LqngQPd253Vz4sT58kydgiamHUnqNbil/P7qZPREZgcRTHItT/hTcoQA0xZ
BXPEt2gB0wmpRPAkB9ioZt9YZkHYtH/SBPH3aFGWDuIepjeg7z+keKF8YA+cwLvf
YHKdnzDDO+JskGyXDJSmXwP3ZiIX4KGXr7jHKW+qn7b5mUTuGndg9Wt0EmtD0YK/
XoHQJyYBwuWrnRRbAk58z3wjTB8/cCorQMInh4B7doMyfmdMygtbmqJBwZkQlhJJ
w0P1IGzKYpBIIl337gnTBnmXuY3tkEbm3idn/1j7lIqMfRlqZJu8gX5GjpK/zEx5
3IaN3DJoVzMF6hq5vrtCQk1DXJKMEfjf9VSVdYnK80Sx4P6bhigCX/G7zPRZYCbH
FTETlpNFbblXD6XtPbdHKiDy4oW7GkfqCuLRDhom+VHfvbXBTkeS0EJTP4r5D5vf
ErjEoq3tSnC9K1BWy1spQhD15MaXJ+BLmkNJVnG+pGsuGTPZIKsl0cS2xJPD6t6X
3cspFbaQh/mZRRJJP+b/vHMKPkeh/9pMF8pP48RP1svhLae8+ue7BKtT2s3CNzc/
rfvu9pADXewn27Lqkh11Pnjc6dA2pWjxMNGGW1F2N2ORiF5KKxPacTy234DuznPh
8XrjWuNrSmTcQqE3nYOvgVI063wkE/FkzCb7T9yEAlAxVvZjYGGochwTJ6W+Sxwr
7HTEoCwTunAfMklyvFSdikflNZWzTNWkF/KDVLr6ppo+910Xv/Ug0iU6d24suO5q
x9T9Vdtb/PKaCchJjSuWujnnes+ZHSg+A1y0JPWn2V2A/5HrIPtAbvAnFtW2tYF9
N4hrzcdfevdeV7Fs9LTp3kY2T7l3xtNHsJH+Neg2xFC3zgWDmzSXP3rL1YsrtoAq
pOK9pIO6LP2KrLetiBvnPpS2wWXZwRweuvzhXUwzhlvs71o2fYc54POy7vMsC6I6
Q5cb+nU0xklQwAF7mmDkH/OolzQcz7tvKDemWXXieetkLDL7k+pNAoK/gAFxgz3x
16GG0kX4Fi4igxROQqZ94XW8HTrL4ZBT55jr+e8MvDEle90+hK8U/bDvIlMQUZxb
DPb+/asDKGATNqaO4GkOsA6m8p/CRXAefpdsLCbuIslff8jNaWLs0d5/eiaDS/2W
zPgfgSHYuyUKOjHo7N6Z6pzZmLsQ2/vJIhqP3c6VAgX6wxQvPrMCKhQqqET/isDv
+bpZocN1YvU/Jh9K1YSIYtMr0864TJcPpTMOzeImJ/paktwnJY8m8uRfWMSxAdmH
wicMlprph/I1kHtJd0inzVZdR6cKqonM+CtDU0Am92jwfYQ/+kLfoRrEsn1QzC6j
A53GnN017VgQxIta7kSfw8XAMD70hDXnGTLFGQpzCC3d2b181F537Cq1texDwH//
fd6wmoRq+ID4OTrZ00+za1+OtlWElv6eFAvKM7YTKMluUgMS5+Uz8jM5pXOaD/1G
HjU9gByOfJ37AxzjlJA/BOYGGaKzU9IWMSjQ516wjbZgrq38ENJ5+lSJlE+VYS6V
84Qs982F2NRzU66VnPm+RhcdxLK3amohhmAlGvYspJ70997jaWzLTJ7NZCBz03ov
7GrY1mXQdPIRXG67VuiP7oIP4ka4XmXSf7tyvCdgiPi9OcKhhaSJ0mRLP/ljIH8q
DybxUy6gogzVWCsezwiRL+DmnLd+HNPtaBymHhC4/NFZaxNcZB8hTMKhdEw1Bd4q
s4+FQHu4xJeDguE9Wcqc7ks/GWFgQoJPq9GvEvnDIB7oEBdQhINpZkP3qpENx1Ei
PHm8EPmL5CB0mUvbToo/U2oQNg66ZJ/HgI79GOL3GMIzWyRFyzU9EEL9h9UChQdu
vkyhef6q1QEeADiq45DeOD3khr9LBKYoiVGyOxVCSlGqsTB1vkD5PX7WrgjmqNCj
p6V3Wigvj01ZlovXyzgD1h02WQ/CcQV7blduYvTR6CGxpXIv75bqeCKsEwCLAvIL
z25g0vBHPvUCBSDQsDsgXtJnaY7VNiiaPa8NKl6MaXjK9OtUegB5vt1/am9GM/wB
zIa0Qk1Zmx4bPMUw93y4jVlaLobXNgv/35RA2202oRdgMf4O+DTWlcmZ1M2NdPBA
uqsnhgISqBOd98N6jZI6/NSwI+ilin+6vVBGuJ14BFMul+t2jhF9u4nGiTMNVz/X
Q10lQq+vVWpxcHyJ4uChWb95+Ykk1rAv/+u/15IB2N2Ysm+7fsaYA2w+06vl0foe
XRhQ41BKF0vGNihkKT21LE0bcjRBLoE+LXzviqvWQWA3oHpgSZJ/Vp5CeGtMANXR
qcx6s2Wb86YwHcQYTdXRZgbHhrLRzZYblqv1bANv3TuD4WiWDKSy9WOYNd5t1G1M
UH9o2oaNJzTo6IazrCwToYNt6Z4yu9Ni0m3Z6WXZeXucXv03+94aixnlkn/VTKni
1JRHri5RFbh3iBQK9uEQMit8x1N4aGxIG8nU/iPWHqO5twlpJBDTHNP9pyOx1IYf
gzeTX/v+VIVCqEwPS/+8rG2DyDW3/vAfuDTL6nvX0Eh6Z3i0YE408Gy3ZaeMHgYP
MjYvo2oMRbuzJKsgAVUfsHrg7aUkd3lcD7BU/w86BhvrfMRLv05xxOlZTcr+4tBM
Gy8wCQNNUuWs2Dqb7KBXQYX0iCeHjxLqKvP1mFLj2BcSFbj0A+PCZd+jh92yZU3s
P0rx+CUprnui0IOziB4+fKDr6fDr90gPppCu8ozKrLmE3UT+qjsKQJaeIyPXiIY8
9w3T86+iBJhV1VrpK9nsZHSEr9Z0TvCWyGplO768c1h0pPMGAxnJAbH5DbP/ce4d
DyeQSHFIgJVKfNFjNRBASlcI1evD9gqgnF7dau72RH9wLh8b3wHPx9IPYAAJvA3o
IYf9ETd3fMpctvgFy41wlcwo4ld1BQy8h4elRkNHZogWzc8YOXm7fNzqEhIlzweR
MLIi44Uo2k/EbetJSi75KluGIamqSsP98UIIlacJZaIwfahFexBwbSGGNzaqx3Oy
dMRzUOkw96Kv8JQI2EQEJekwteOsDg6yXNbJtej+ANXeZMbVPp48RR9KQJycZQE/
HhDCUnJZ6QvF+8OCm/wOuvVuxR9Xj5btjLdKR00Dq4w5OzmRWugLKqnMZxnpqxlP
lq5N0AgyMVRkm67QAR96+/wMWv9c4R868RZS4H7n5sDkKGtQm4i/EFwoJbQQ4JpH
2hB9YLzX3fWXEvcUlwtDaod94w+UjJLOsuk0KFbQ6zOXUTTvRrgIYxx9RB5iHMJ8
Z0DKBOuXNULZDXW4ztQq8JCtVXVXyBEAaYv5zhRvIEF6r1yL88+ZAqI7BD80yAyd
wjDrP3vvbHyQLthMT+fSgrIqcIDsYQBGFw1YuMwiI/L4sijgyYK1R1LHmjawn94E
Rz0zcHhubYM2KDMBwpcR4Aw6saINhTNspvcbdg2N19ttiL6EZpOXko8uq0o/Px8E
Qisg93x5SXaCsZam8/kWG1aEN2fsrHjAhq+erocHpM6kyCB9J2o0egpM84ZlkGph
NEe9mRz0AwvhtoUZODTPIgGph2dWc00x93SFkbsZllUqpv9XNmLe6B5fVI0pfYg5
dcx15Hrj1IT77LU9JeLdo+2H4psbnOSRwBUSiCR5D3xm0OLe5DGtiHLtvFUI43jJ
4k/BfBMtWmCIPQZANtAmb6av7Tpc12Cs2BmBQLesfpGyfxHYfL11JaMS2FYmYZ24
55Ch0piAU4I9jD5wjx1k+TcG/1cZfqQDHv9gRjpUrsyj+14YAt9s+1KB9mQf8hUL
YimKEaG2bKJ6j+sBgMn2W/foeUJy5mWChlS1xBdvkltV/joZQhWF1HgA96F37t6a
RB3FV76MiZuQtJ6fpliI/9TjhIXK3eRa7hInS5j87//Yxng92YvRFzNWq/H9ivb0
Jm9Jrfqh5Uzm7EURfL2FxVMqT7X+RqOK+2Ywn3pXHd3Z3sALxCGRJXQZdQXwK9rb
1gbQRuOuHqRTzK8fli29SB01TG0fQ4+8McenuC0mzVOEiKm3Ki78YfqrqKKN1X8c
xe4fKWvLRl50ju2iUJL/9kHBLFUJrqa4Fywu+K48VjuYx2U88KAo9T+t2AfjUAXD
u1oqUoNpYlc/WksDyYwSQi2AdjBvswaQdvUPZ0bTNEcp8SCVK9fXOTtEI5XLtrpH
itI25VF32c2bOI1patC8TAjCflg6C40+0MG8yqrJUmtH8zhyvTC47FyAxeU2Gwr8
yvKj0CSQ3Qs5IyPgV4Wyk6lTMYIJCBtum2LoyIWbATUxi7OUZuAh69xm8HVthH9q
mdnKb40w+fNpaAlYPHlJGQHO4kAckHvNNd26frIEpt/jJlGDxNZbiAfObk0Khnau
1HyCIyvY5PzPhPelaHGs+efmtfwXp76w8G3ADI28fqeriZtpNNei4XMEuqPGLtYZ
94FJJE2jlcxMDATVw1s2uGjXIFuiKhInSHYqLXrfapVzRlCDG69k86sDhko2nVzv
fjK8QkHEW7hI4+PmvLB37tfr6LYkrhztvdHLBx1SHW9GRS464T+O7ZG/iIwqiFDA
miaN8BF8/xzPakgiybb9p1qw7xDYTqaXKhfuPdFbYtir0Ewir6juc+egKRxLmz91
bBSMCyg4YCls5EJeln757+5Q+O9J/HZZB/qdrVASK6BU5y3CrOYQIxb3FJEdDWHD
NaPJ7v+cne3TCHlNflYIrvBeqLC/iex0NvZNnyxRFrkxk1q1TYT49SxjLnBgP/mL
8ptRNH6HSkuw0C+yuYldKIJuSqdHB/NKblXaym5TaicikvevEADG5Bnz4vpNXbf7
lmbFHH9d6RXpj52rBd3cfB2rsFDf+chbg10iTUS02dlztuK4jsHunmXmqol9Dk88
UPGANAeJAXzoRybOAuINIxoV3YojCVSoCumQAVGbhJz2ZIRyWaTZiwELCis14T9z
Yku5mFLLZr8CNnx4+Vkca7xD2rPiEX8IDJlTglLd4IpnhTqdksUNnYqCPqupBrrw
3Op2B4DhvRRMTGfozKi3kjwn2faf4NrIY2r0n+JIPpqfxq6x1VJjpd2wyRP80Yuz
MD/otNYNF0km6+pnGvRiVVySYkpZaFlh5McAT5t6PrpGP4XizOgY4wN5gwEjBz7U
iRjhSDAZhQqeSbJ/LYJcMf0+0mWBmpYVgfO8xs0t+Kvm0a9fdie7HmuIgQON2gbX
31KSr9znd21uCyCzMHxxzJO/Ho0yb/tN2Tf96yC78sHb/CrdYSCpGTLhXbdVURDZ
/DEJzM3gAY6RvVai4y4zHgAbrn/hDe0Cds9DC4RwO52fseeSPhcQ5YfWt69DFVl0
AhhlqvZnO2PjbQP94obwl3WRpjxxpB0HNwjsptjjU+xaVHl48wUbCO4lKAoHqFFG
VyrWzxRz5ZTn2RjTlhmidJTf8MDJhkNnhLvB3D+0NnRgGBaKd9wYyPdoTkY6GubD
LYnFKCI4G2qclB6E8F8K73TcUdnq53txS6ONwjRq2aXNQ+g74nCMjBDrhaQQ8iFX
jVnOIfhOnx5x4J4eVZ1IRbqoPX8Wuh5/yTISVEMpO25YICe+wlqnn8QOGeTBQQMx
1nFYgGTQUMQ60APQVGX/IehC2fnHOlD0xBippliHKaudwz6v053nsUX97XOHjpDy
ZaMwesbuz1AYB+JA9GICNF2gKj04tYXYtuE0txHiuSpjvnJrrzaDXiLGAlZfS5yo
k+Rc5Lby48y6i5Db5c+HfrDpGZC358BPWDeN1xNVWjnawrEl02czU69pcsFs9HWO
Be6SAsDymqiuIW1ki8xxX4chCMl50AeQUeGekiFeokP9eFQ+RjfRXrxz6XapNxzq
/5s5PsyZ3DjSatlEI3TLSygR7HjC4SoR1AoyN/23hHs87kaK0VQ/qdVVv16D2BV7
Bfur22Yoczv+IvwZYL+ZBfTm7VfR6asBc3fmFJL7OV9gI9oy5e4m7wi227TncW0l
rqdVo452nEC1CUXXzGzH459PfZAjAfzPU8yN2go1rBZ+YJjY3ch/3DYImtVLHlee
HmjqO2qAQoHJjG1644Qlf3ypiAuBNFHWmna7ZIZC+2RT8n/IzSXC2RH/NK+G7yEq
4qJ/oFe81ClCbvgyeXJ53FDcHV0LqTaY0qSl30JYMbAzM0O8cVkfx80vD2c8CGII
sYOvqOWzTGSohl75txqC4BcbermsIXQWj6ZaYvM8omk9lYES+Il+n4YXfwxuez3O
5Qr129Om1Xf0G0igs8YqLbujHq7cVNk0qpEnEa/v5udo9Vrd55mqSUWXrjztK+vn
VTJeW/OGMEdmEoqm/vKR62OtckLnTBUzWGB69GuLr7cbWZ623s3OgFYI/gUle7H1
rhxpTlcqnqQlKEXI7UcBe5ILcMsIGD34v+ABMVq01sA+sSz2w73uJxz713/R4I9h
d7l2O9dDLvSk+fwNywxDji21rVFMuvamjFfdy7xMu0dVKlR6vgVd3NX4fvO8tqGq
iJ9C+DLY2yQa18zypOq/p0/oDe7dodEgJcsMpBGB7Un6Vz/+Cvamihh6x250jnm0
4QYfWlXeonyclqZYme79TaDZmBJBLeEb8ibGF2/MdZv8ovHsUKe928+d0unaCXNO
dyAXwePV6Y6B1L+9DaR02icOgro2DKDTZz4vo8b+Y3Ru/1JwwSobO7PaSZX8FSIh
YKeGPrqtovnbPgLZmjxBISTdwFo/QeQ/OVJqtnt3qM2XESgBOjguuqHXxb/0jB7T
ccbMXnLsF/YlF+vInWYayej4LpeVWTxoGjpkmGp72+VefRdH3Cow775gU/owukz0
P3tTLgGchLsXx1pelKJxXDM2FQtT8yZf7YxQgwLoRi8QT2mNdxf7+/zsO15nT1H6
kQ1yDjjpa8V3JFpIziP8zRCGe/fbGZbPALaeXUUSOnKXxMEoGhGxsLAUnF3CuMgI
a9inOynRQpxJufNMp8Wwy3Z/cGmzu1j9rZfNt7BCOSFyZ3JVfhv6oeU0tRlz4Y1F
S4GuUlQSuDfZrztDfaqMxnPRbik9sOH1ixoktxX7nmxRDcHYs4h2rIhXyPdMMyNW
e1DpuRI8Vgdex7gWxzqx19euzmcuE++T91tJgIeKw9qMbleN+REe7UvlEodtkNWE
bOgPd8X3ZLuyFNxm9N+S8E/JqtGCOcOx4uLVd3eGSRp1INQ/L3NSPxgIq7koReiT
TZo+AAf/HB1t3PEceelGivcNzGX1ZfwyimhqvTWVIqC+MYD5E3B3py4H4DlnKHy8
Ay5fMY7Q2fkzkt2nRhzvFo8f3i102wyn5z6DBH3CvTp9S2lOJHG88sMDBgzoxaco
e8N8HVlfAM/sclqD+HIjfzstrjD8Cx32i5e8NjVQP7tMeaH8dCVIaqYPFNcqWCsU
9NqMCPMkWBjXWn8XT81+fEYFoh7+nsA9a7JyrsboY810lfwk2HLV9baQYHUpHazv
dtttXlM6P3HI3+Ft/RTIIkfvwNlAOTAl9mfEU3oA8t2Zh+tGVUGSMTfAyFg1V4De
/I5A97WrWLrk1dme1on0hJAZC3KIlV7HS9FzqQIICSBPvs9sHSytcIxpO9S/hYiZ
X58h1+MsODNr6geZ2rPHu8UHbDwnFzold0VopUgtTodG4rDyDvsYFx/QjY+ck3xr
alARddqoY/DuYk/YDqijmCKi5OofSANHcxD2/HrV7M9JsogNA3sZA/BwgA58BY5R
CGa+jEuFms6C/bqyp9C80pV5bT2ziATCJaN+/Nj4Zqa0ilmzL3VYKRGEvRdSXDm/
pTVdVC/06n0K/2hbGPG2a7P2FqXXTwccdTYAStDc7ukkbBX5dcwEkuAZfT16JBOy
sMJOhdIY109lDkUI0ZzaTUBPC0YUrj9F4+nYdNTkb4xE8lOIrlXksZUTFe5nljKq
z9lExuiP52FIyWPccdpOiEHb0hnXH/n4rnrVc9XtgGajVtpT84ExIgZjQ+1bcF+7
VMOO8qd062RNYrCdtlzSAEETeXp+TcVtD789oI3c1/BcVPWjwuvimWL2y2oZjRpz
XVKkmTBOBPKV5Rww9n1bk7+EE+zn6lyEByjDrn0f7WPYFT+V2v00vLNe7SN2AE5O
qPBbW0xMU4XjyOSbd2GnuNw3L8mRiWQdHiTB7jLol5oIteSL0v6+33W6b9nbSAgN
brg27Pc625wkXbhy1UsfDCvlO44QuGkbV/spX9K7gYql1GGlaAhfl8A7MSGPs4Fe
CJJ9d+KKQD8fZvrVSI/KvOM8z5AsfTSZXhffY2AI9zxChiWXzq4UaZVKuU/9wcDU
Qc/TAFVCAhl34K/Gaqrmz0Es5Au3qx0LPoQ14wfng44SN0GBdUFRTprp4HBrZr2r
p4vpW44JX5hW+reZIm/i8cHqGvAmPH5Uv0p7Pm/mYl6cugxZ2Ufet1/b7TXE+HLy
PHopCC1vs2bOUFlF+WICgV/pgZlweA07HaSUCl51DSQKKYyhI+NK7XBzOXlkXRAs
F4oJ+3ll6mthbQZhlJPnzbbB+n/gIWDO4v2r34D1LW1KH4YomW1V+rAtkELZxLOT
yNjR5LCaWQFNh3PvpYhsttM+6RSEpGBhXKYSsgye9LfcvTh5zHLzgUew3hTHt7yO
wRS9eWeBslcXa54JN4mNR2qgM9nAMdsLDdw/leUUn9nTmvhXXbnY+vB6XGJ+rddU
AYiPXFmzyAs9HWjg/k6oMjSvFH7yLJwp4vg1g2Yp6cU3b+Li+WpisZrqlrzxqiS+
6jA3XjhI4k1glchu7pgjRtEUlZkCmHh9ma1LD82apt1UGljBn0m3JGyh9TNIywpx
3ySCvYPEcENh2IMTjLPKGaRPqQVnpkFdCq4u0oSr5JtQsFpdIDUdccsAIbbWk0t3
k0KrB3yCyihsSpXnPBejz1+URYJ3b+CSUgDRdh6Mdw6ZNh3GzA2jkEz8JEtnFTv9
sCNrrA8rTMNmfZ0T3fhOAWgG+7t7/EwWBOpWst9z4vxMODIWtBwpf6BT/AjuuERf
EGpYGGB+epc+U1umoEDLZU3Jh8W9wZp/iBMjGcvZHV7wKEmTx/pz2KyDerpahKVz
Jrf4sUYnwwgLUnb5cZX+uD30JSWuPTzrCCWC7djc1UXoNUcHceOH40Kz8BjHlybm
mpcjwUZ6G2LNUC5mgqu4gxdLErB1104EiAnteud9m+/q/VABnVhVcPFF5kk6Z37O
5dl+HUC1S2UNt3S4tb9mDoBCSJnUPjKELlnjMFJsoMlKFWU31+DKuKAntWyozpKN
DCDn4NRlONJVaGWaEzN9DTBlY797GuOPuKk5ORO5uYwOdnoy2OwrZSq+xLvzHDq9
254y4G4R+tBxpra/CEZsPRhnSHYtswouiRSY6qGLxDEWPJ/THxFuQPR+VHIMZtk/
8Iyr7ORuAqB4aU9utNNNXR5UONwk0nDN8wMRTzyDHvxA/1tQUdvHghFG1qcZukM+
VjBqGrxUqDK8ciy7F0+w/32gcEWAQAllGaZJ/MqvLNTf+UvJDymkdRLeiZ8zr8oE
jh64/55xnZRsae3aFw/GOP6Vy0M0yXf5rBSHO0GC6RR/hZIr7CnzqCBccdd8NiMx
VA5TwnQlEoH0Tgz+ZCuOlme3ckNDw7+pAbbTBD+acKwk6IFDUv/ftx+OKyhLtzbR
TMKHqFRIdfex8usLiGXaf43FfW/jQbvk0TsmamE1o1Lsuru+vjJlLpgdy22cuh7e
k3li8Jcja0KrfPx9aoW5x1mC6Fr0ZfN0sPTLmujxw+XhF2HmVBfcWT6wIRvNori0
NYwzAq+GgcAT5uVdLGesT91pOKOR2kwZ2PkOOeZojkROV2rdZ3pFFu4zO8ga2gEh
qAuwrOVXYBPGyCv1dkhDgUnWD8Aaic2ggh2JW0jN21jVplSs/cvVhKN416UF22F6
gsXJDgROUTw/M117jXPQwyT0ElDbib9Jwim6DEWW7J1qIIsxjuPMfIqL4bsgf4/f
5jeiAv0haWM8g+oc7wvNEghJFGxTAGywGh6yzU/yi9aWxTCiRmIsENnUCYB87Qxv
+L3/QYpd6oLqX7SxHFTFjCYD7hlk37Bl6O9pJb0Lw6f89DUbDGgLW4PaALSo5R+9
u0FPqQ/cuRFEWQEOcYmhs8UCXlvelvcAEOlUvAe2FlpzHBWr4XsTuE/HKFB4hB63
OtqkoDjEx/uqaX6yEsPn1CqlmXZoMqhbo99stm2SruU3E7FNJQYsIOQBlCT1fsLx
miSBE7yME9qqA+sgalBphxtjqQBOuzM5xlxuQMwZHQkohn2FV4PFIkeVy/gKVjhI
qLCpZXpT/zk+NG7WGHBnQ6uOKj3rX/nQyJVuyaSdllRPzhC4h6wCjDlKtpiNRjdC
tt7xeEeEGPHHWamHWbv1r7KzX97nViP1vFYlaEWEXKH5Xc7OJQ/mhOuQGrKlPJU3
Y6zXVkkNVEDbb24HF6TFsrhiqKq0/6hwvSH0iJRnQb5CZfgJsVKOOoeEU+rv6Bly
h5wRLK/vSCCSSZqCJtB9hRrT1RQWqrN8ipVBbxAYMIofpV8G5nyWsgGD0A1YR+t7
FyZ7Jd7K0B8DweHtm0xa9jPFnZpeCJorYkoNiqVSniG8A/QWqLVu6ckwnGkL0EvM
K7256xzxv0hog0I9fFcNr7tN0VwkSIntAuS00oJlIgID8WEVugWKitT4Q6dQW8md
+1al3rd8g/Z5Jf9lFBw98f/OwMK1Q4lgWK50lZhHBrCrhOsWz+XoUunvFwb4sYKD
9MJnrEDGqbiPussTVQEFOGRd0Yv2Zb01n5a4GdmtGVGNBGv0Jct+iD1ULFITbdIc
ZioY1DnDmNrkSChUklFvQk0plrqKM8BpVuSpqGsvm4Jyrg6ZWPy3QedeNXOfg7CS
MYf3MThUdb63OtdYG8gMgrIiTPafXfJdLqcK0dxZW7JQgXej+oEvBaQ1DfGapBJM
wKFfEHy9bH6diQh8F6tCK1CzW+hAOb5UBzuw95KCZDjrPuxbqki8DLXWgAKBIDwz
hZ5K1bTc+mSMUlwe07ZO8AK+KqmBEF4REx1vULPK/l8BY3f7DLJNHHCLTP/5Ljev
/c32nWjnR9D+tMWZkJ6Fnlmi1PvyMMVj20GE3XR/9BX3Q71UO+mhoqhsiZ75FB4T
Br50haUeeLr1aUXznSq1vTyMd9KRftzbASFrGlD8Kjsehal1RXizKANQPVyzngiU
AKtYAJdp4BXobhszUePxMJL+ejOX+UyS9lnQFPLa1ncwyyhzpP3Iv/AeIqwrojYY
g/ag6P4NKOcQLOebM1sh3hyCGyFCFVxIJxSaYZ8w8jJ4AYg+8tB+t6AVDvUohdlx
HsUlSc/9jbQXGZBEgBg8Mfa/qCye+Hc4BWuY1vxFfVxjYw4ZaeABICqNDpIa7QmV
b/Ewwsg6qvDN851GBKXFQ1qBavYGBHwjuDarE0HmOetD66KrbyrUi3DfxQfwwlFh
BD7cRwjmL3ehFmohFqhU5R6aDsLyQGDMcyW13ydoknewfmd4l7dcwa/5ZxyPEAX0
sf5pgT+gxR3Rt4yWtMJEEbrIjLTiSUlBaxvlKiw3zm2A6kl4/ATwzWDKUqNrfOkj
KfZAdfYRoXGqe5OCraECanmDATJvo8yQ5l7PXU04woRU0PYJqYRT0PK3hJc4WT1/
sDKMY4triZUET/N105ozU5ULZ5YheidWPNlhqWrFncZ2X0DYPZIEokzLFx0WAZe+
ThQZ6rb8YQZZbLP17ETYP+xOyNJFgpU8vnf//zqu0oTE4y3cP4NfT0IQYHMGSKej
p6pFzNemggyVYGrFcvCkrGm/W2YwD7vlelq9Cpkgdf4AuXkDiFYFPvx8tDO9fQPn
8sdeelrYAEV+XXDynjc34ylcdti/XFN/dV1jiaVI+KMTys2uYurGbc9aDh0icTum
rWvzRi91FbDTx8D/wpao2+JaJRqdWl+uAwh3dUDUt34yjJP6nBG2G9M1I1O/7h+g
0MrUGL3BmAywu9UKJprTiSBg/igD/NEogRO+KGQ64uuEG5ukIyMCefRpKpsT43De
IwEXg4ZVYj2u4CXkVkrfCeKGa/MKmWtkpGGpAHsUti5Jird06vkZSYyfv6WMhuPC
xJ0kUZf8g0qq04ToDakZduGt1+znG6xYYdB1IrIbtw9xnWgOWGoDUCSPPcMxjt9x
TwlYkq8FEFLP0eO+cR94NQkBqRXnUs+LvcK5CubdwulrqFV/ic+KaL05ztZjFKKH
Q8gkB+BoEoaPzkygxzCqOcaeXJjfLe5S4egxnSHSMdlw2DocJtm+mrT+S6FZHOTi
VBClaCqxaqoGhUysjo/9PPmx3O9H+kdw6MfxQpgf2dx8WU7BPeJu6iWpmykW5QhF
rUQXqiN8T2IU9o0LvlyrTgnbZutwTLD9fUcp8HP6OMVOhNmmzzIv0ivdiIo9sARm
d0i1HlK+YHthiIjM+/+CP5/X8IOtGv2GU3FEblN+jIvCJcv4yWJotLIaI+4kcYDe
WkieqR+49nyKVFXFPNcCIfoVif9KA3dFsbjKIrqp5BxOIH4Dj7qxRATegqFwp9Xj
E/ppC42gmaeBPCw9YB4ffB9CaF7iEE9trR1DMkhhYKUy4uDXW7yjHcaa1YJVcBaz
QLa1nhuX8qJAkxFUcC0UGfufDtiybBWmxwUoHjO6Le9+2lfbr19H6IUpDC3B/m5K
QHYuc1sAUmFFMWdau8rtdvGP4Kj9ag0MMrdqrVh1xJsIuRYvBWGUXKkqHITy/FIk
Y+fw/XKyzDELzac/9jZ8aE+y67DtdXYv68JYWBwSoN4jCc7u5wkAEDSGQ1TlkkOw
+LqbUwK2jO0iONTv2xIQnmLAIujv6YgKOHpA9DwuwtnC+1UG12cXDQWbbKTezVK1
x4Cfyls93bSmKocwUmOHKKwXuDsGfge79LHrigneE1yQOPjfyzJCPOXkI1JhEfpS
k3416GkEP9vDjj+pqtlaXJzFDspaBXx+xTlb/h55VvfiYwvML4J5WBnD0T3EgXZS
KWEOQqCKcybR5LCmekwyxFqpTQHuJ2yd88tGKvBdNhTPIhhC433YX7bcRRykI0Zo
rZEBDcqPZ8DHtEE3WJ+J+uzaH9g+G7veJsknKHZqDBl7Uy3BytE8bVu+gnYO5nah
BA0SZp9G5mEeOeXGGpVo9WwAdC1BWkr6TgnBe+3bSkafn9FY6Z2GXzGSeiV7Nufa
PanrWeZ5oEPM50f8U+kSTisP5UFkUX6IC85z8czN4PLAzE93Q1ZLib9h04gH4AB7
lIQ0wWIjEpIkpbwfLHB1ZxjisP6s2di5THQhH0tdyrKqVB77wzFhaIFzecz1f1h5
egjRTjHRTdI+GKYYs/iadez5FhPhxECcug2izqHAYhwjfwrAcEUtTprrIeWvKfXW
f2NMvFg8pcKEHif6GroW2D89mWjYtJnmpYUGMr930cNlANwLWKLlhMAcllOWVsgV
B8E1yTSATGu1noEEoIXzdyhyRiocYCu/zmS+c7L+Fod4wufJf6oylB5DZus/79a3
vKj7gGckz1PcwGDW+5pLnaf0WQ0jstAKDm6roFIsyCgCTblEwePeN0D694pqeC/W
nBlOW+t7ai794fjl/CA6Jbpxv14VvlI6h76r/B81JUFcGa21Zo4ku/33MOpi81No
76hT0RkTBldcRciFD9BcIJuTNwjqLUkSUbY8obRmQ1FQRmzDpxOZzueETUs4ajhW
FDLei4akqZiCFNGCn3emIWmErICWEfdiMGSjaQVCneGWWhoSgyhE+57/wNnYD9+l
2r53H/+l3/iTY/N1NtEybYipOHDvmaVBAb0lY3ZLZ0LZRNeoDqa4IF6tOjR1/HbC
CXxMLcESXJTgBKVdgg0eoDO9xcEn1JzwJGU1oGA64b6CS6vzpy1jfHj78iGruGso
IzIxZ1LxU2JGGdJqwIW5V5boQrJcyuV5hWd1Rug1aQFFSnt1QDNYk6DMAlDn/3HW
/sYfq5Vz5ckivmgbON04GVqOx3RcNdlhCXPBbsCUPJ+XSprtWuRz0hygt4JtBb6h
4D97eJ6kv3vSkJuC9Gp/Cvi8U8sEAS3a+9sRSGU8a79UcZjeEQO3KPfcAFA0U/Ku
KmQB22G0uoC0ClqaDZRvMYPWIn7CqcLNWyQhtBTtIMePejDcYtY5z0M4zCNOXhS7
R89EAEqpGt482s6IVdqQ988iym+vvYH1dovAvPU2VfrcsK+XwRAVb4v/HJBjTbYV
Zh4e2VvcboebEk61cRLlG8DDHwADd21iS7g5tKFz7FugFfoLLVBXPdHTT/+QavxN
mmCGF4c3BnSkItVuAGJLnZS4HM1yy4AWdnTNRKBGee0d5mLMhTeK2Y1njFzwuWjf
8OrBmgswYFRwmJ9hUoNLydp4xm1DTrkYOoumxYeZOUpZiSJjpohxPSk0PGSnZavA
zYybO4+nWyVHrQBFvRhnhDyHMkDKUp3Z0aqFQ3ojTiiYVi265OnGenZNPW0QxSx6
ZDtjq8bf+ZDpMI6dDuncYnm/HRsMbHn9pAigBwODkrETlgl5m5PylwMJ5phwA86f
+H8KkmZeDFn/rNYawjV/FQnaKP8viGbFrbYdmdhihqBNJo0opPfUuUfvMxsvT18T
WZNP9fAlkKrjlhZXGFygdjAmYyUUk5fPNXWKYda3Oh5bGfILmVG3YRsoDe+GuLWA
Nf9qCztiekqbAopfEH8LYQPE6N2JRv+pKaLwiO1zmCr78Ko8raKAsV3HCsbu+AJk
VXehuopEpbENmbLPEXgRHrZyOuvo8El91HnOPzuSCQu3UG1Q2N52+JDZ7sdSEeuL
BcmMivEgX3+tD00vDGJFBP50H4SvPDvEJkhGpSddhXrFxhVbwOx2TRQsqglG1MY5
K5nq2jG287YtoMhnBJibvvgC742yngwZqJCs0wCdmzU00hi6IHg51sR9PWds5RaK
+gOs6p5oVjWKKjjw08lARC1uOh7lpfegFUnuDO+Pyidz6t8eYC2rqdRF8D6rjWsx
HpRHWLRvkBatEiq1cY6ALZbre4AFE2ndK1BJJxgAjK9q2ErABqJFYSMEiH8mA6D1
F9G98O1A/UAUmVwYfwHQzFtZxR2itQ3JdGtNz5NE/FTn/xrk/y/mFH7dO9RgOUx5
WIzrnVXd42m9He8M/tiLVmygAooWnio9z9G5xEMcwaHE/zUhi9L6LhlgqqZS9YAf
PYvUoKaciiYot4VbUnmQiH0AmdgFZLrFoYijyfOr9PbHLiIK9HPU1KPLIhMAvk6f
3oydtfZrhwl6kEUttFZWwSHE9HILOrl7D4uESbwvwVLAyAouSP6YGH4LYQy301Yb
b2tbPnVW1gqh/N6GQK5hfoM5zzFUk70Lwex3My8yOMwkzhj9Abcqlwda+qsJF4BX
HsUdhWkT637FTDha/gVBw/40u7kbb+3TCrvQQYdwIrolbf1eCeZ74c7gNZ4OiMoy
xZVsyGNWrZWz4uvr8hcAvMQtLRRqY0f5zXf26xa4240CoOsJobDRysP4D1gKb3hc
SRYwp/i/HDUWyT5fNT1yjt8uEhp9lAGZiuDClGu8zGqYBCU5/Fxt37R6dMgr6F85
17g4Bmun3VuKlGrZoxu/qB/Qf0ydELlBmeHXEXXn3JRSKj/773aVHEWJC7RhF+7c
WPjDJBgjqWOiv/Qr+PSoEKEBWPNdjemS64AB+cIr5iAzgdGm3ZamNv5WrVJIxx3V
3hhTwgUt929U8sn94kdbiPLG1hPIO8jBCLRHjp50t0Fy9MLNksC371Ir0kzQ5Uyt
UrdtWb2cDQgeUkAjLzhjjA/CIt/77A8NrxW28e2IzDH3RbFjoYB9fJs85fqRzkmE
+rjrxNYS6o6NMAz1j6jI7oW/Gkx7Zbvq78C+yAH82eLau+6X5DVe8u5iCS2bmuib
ON3cIqpq1fqu7qdCXtTWr2kDgMp5Cvo+wQrpd3IDg/hTG/FR//Htwsg7VDu66OPr
4gBdVMnWFm+xacd3yZAZvNjvW7rA1WxbqnXOYaqM4PPI+o+Z37P9huZc1yzz8vHx
6DzaBA+ItEzoZgRikGTTGbkpQd7VnjTZQwIYbaD3was5ARw6G1mfi86wck+Kh7k/
DNKvT672r4YokOTJZU49unB+Tp7MJxOmEfkGeS9DkwweV1unwLw5+zAoFdzrsMv4
k8sJGUjmIk3pmzmj405QU2gbgBcX6DnaH+R3JOD8XPH89pErd4g5cKeb0ywB1EL9
KoH6OILjuI/jL0mArfWHWgxmfBrL48TbfGB6LkuMpre3lEUnxP8FvNKUtpia7HQ2
PlzovvJxajASlKn3pHsl5z2/y9tsmCEzk3HX56J5gj2u+KjVh87Mqgc22Av42UDQ
aqAT3LwSW7buM5TXzE+Wn9CTqv1aJcVfJg9iv/ca2zd9c0iHZoK3KULTiq5g4u9G
xmfCstLbIN7hNoLCdg7HLhhd8Pbr5bupA2k9Vh8Y9rtOt1cAQg7Ipoo+4S0MAeHW
5yJChVZ8NyoOhlQHt+R8zSWZaiV+SP/6gqCL7pEzj7/vDl6PL2NMsq4nCGJE/jFM
VazY7Fa4YHjIckpL69PrIfs/5uEAgeIqHClZjxu08aKevP9h5vuFTUgyGJEfa276
R4xjCn1ELAhjq/fv4BvfQM6Dm4t6za1MtzR9CjoeMaeNiC8mr1w3MOc6/S86zUZ7
ZrMBL2/8FhImXQD21TE7ecaSSrBEgZQCidtAJcLIgNGDuEYi5gGUECHZD5cU57Lk
ju/84AaLJXkPcAe/oQVMkT0ovkoojWqRiHvdlRuCAh3vtIXq1dMJZGrGBhUh0qYg
2dU2gODvkfD2oXWjv2QTsvOZOaLLJuiOPidzhtpDWZFSo9RVh2LKaMjDSvtuDWPo
1yhpfQDa+XdI1KUA0ZDhikIN1S6d98xVFU5Y8eXNFPIPnJKx8t6Gq3YCthf9MGml
f9WDZVymqn+7N+9oZsaGhjWOG0d4KpuT6bZK/0YbtnPxfVmxd93jJ2oOVYzjD0cq
osRUT6y4r9ll+7AMsNQ5B3y//I2MNrnBaQBTUCHPg+0ykwsge6uHETI4YQgCd9aM
8qdMtM39uxogch72DtF32w8f3EgNZ3fAvErn2a61sKUZFCUL+r0GRQAD1JBHLuUr
19KtY49C8AIHfPn1CKK1uyoA0+B9rhe2fq3yo4HjRY0aQToKG+/fAXZ5jdPCaeuU
q7TRltPx/KQtscGqtOD5Yxql7FsQRJC/N66ZKBp2IBaEzHPD06YS7rGLAJzFZXEK
Fp/kskB3GvloCInQlyDlKEH2ErNx7JDoqjfov9AS0NB94qDcKatWEB5UbLZpU3g7
z8VR4i255WHtfGTc5aOefOfbdY90/xvjXqC/dDaRvzntNzH5zA9o41/FcReS/1jN
Wc1sbUDT8fAkXhS8YyPDqr34v5B78cuvjJqPuQE3DLtIDU1x23vsRbe3F8ut4WRk
FhfNZTDScC0nkyZN0313W+pL6wSRzth4DO7IeOCQw7enPLQC3DeUtieWoqLWx+WK
O34ue5DjkSEg7Dj1CbXhTqw+qu7A4nHGxs5gxU61Wk7Ny6iV+29bxoh7LMG0fi9V
ugdTi7Kxnz48NcEx72htUowv33hQtf6mH1Qkxp/5c0rGOJV2mKcyv3xRZpTpd/FE
3LwgDtM6WUwFb7DOiOnq4H8+vMCRvp2sFoYwMDgEvKM8jX7IFiLByhOrLXrTn0Dr
zTzZW4BbHehKkcyoY+huiDOuZsH7WgAWbcRx8l0TDpRcc1bbGtBAzcTrG6yxnFKK
eW6uCV0Hsu2LJVCzTnZFb/kFO0Qn7W1k1JkK34xvnmMXwKcLImWCnloCs/GKY9Wz
sWRQSrp8ozL+JFRg7IIH+Zl0iTYHs0JbEMLB+do+uYfoKFiyIFa5c6xnC0m7RcEu
gG71wYkjTW5T+GAWbFr8+PC64kbdxOs5Trx8m1tI+3bETIPPwgdGTMr4htweUjeD
hDYxcwEVY9Kn8bGWjvdWv5OaZJyuCceuioV1pO67tKw2FOgRQT9CtH7+BvqYSeB/
gCDTgxg16hVY9WxrPVBLfkwyUB+TNc036rz1aGRlrxOikPkxml+4hR1+EVq2xuay
iPnY+jC+EqpjN1tU/8QoaLSIrojoP5+7gJxdD7FqmD5OtaPZgJqJ0BleMdRGfIDD
4EBB9PbtDn7CMIpb/VB+kwy0hOpSrp05EuoTqDlsY1bJP42Xetk0fsERkDOIt/F/
OUpnjm0LVR1VUnyhnylPZJbpmD6sl2vvwhAc+Ow0NVcIPt7ourDn+Zqx7CDqr9j3
ZdL5sre76XDQHgdyWNdy28sWPWi36oB3xOuJDNsW6tlaS9DHedkHcPEvMolI1B5/
4BTnFfG9iKDZRJyKbiWZjiTTNldeMBIch2RbzoWMUDKWDQGnKGTvXzrMAXs0L1Ez
KtHdoHgIY6aAuReOJE9XzmuDb8xyG6lUGHOxj6SyDb47CmHXPGNZRMDikI2qQK0d
ou21/a7xeaMcCo6HBeNQ3P6hwyNHxmWRUpgKUBXGcrDR4lKFOIDO9/9rdJJfTiZP
r6cYDsaj5uzgeJwbMWtFm1NMSzd+4vOgcJgbnNYbUIajK7AafrX8N3zmBc4O4bU+
n5tASFgOQ2oI2k+srH66F4rDXGRWONJYiZ2AD3S/TqkJwMa7ywH5dT44Bu4kgcz8
7FgOuLQnTjNsReHCa246rAoUrdNr1qubU4wDi6NDG1zesAzJ14lf5QQY4gBzmcOC
/RH15cDLe3V3OR9b4NAfo7EKN6mtWd9ePUferjl/61l/952BL9xEFJbqKAv8NS+6
hMZcSHz5cEPKXYMvYvGeakibpyQQ5qHRV/o1o/PZZ5buhbcaR18fRyz0ORs5xthd
f4BSi0kx8W/WIlWox3IfXBwhrOLONZjRHu3QXiBPEFQGtgQUz0cB/4lFN6Kkbw2G
X3Ts2OgAt7Javc/aFTKchT6TvfcLQCE69Phn5x6WVUWf/L2GskmYurUaLgfb0EqJ
sNr9o+dL5GVaiWJfJJ+kgvJOYeKtYpy14OxFUDg+U3raIkmVwiF9AzPPe0b9KLa8
IRxE95GQLwt8+gWTcgvO4IeO8uNpi9gLKo1LARnVPUhWMnZWc5qwg91DSPUp3p5M
ghblBbglxESIREyyG8XxiIWNVDI8bBKC+grJ3be3NCQBZTovuvuDdRxaVpTXVh+C
MVr/MEmOtTnUR01WgPsoMQShFoOU5doW9dV+N2YXRenJFc4KlyNvroEM64/SHYQ3
YUMYniO14rLoXT0oAAMsmNAwM4MlZCtAnpIr1PyYDWzDJ6rFvMfpcu1w4kN0IJhR
Hhfw5y9ZlBycxrkN6n1yBGdUGgTbxEMM6f4trlHHxSBZqDmibBcBmJe+/5Jsm/Au
JaeXa5ihxDppYlt1dqDB1H5vEHyORdxbnQawRFCAulbbKu+wt4STK7tYi3pCGary
olKgqMhs9T0aUdtP38M3PQG1FLrG46ht2kFs8NkyOi7MVMkZibsH8niXgHLIuBh4
IONhjOdKiguqXUs138waUaDJ079qi23CbNszSJFzRiNsWoWBM5QUb6dCi7eGrTXa
gFlL/HriKNr0r54Jn01l/Hehz2f+DMudt03/OAUxpiKSEjlDTYTAxu/p8WbPLWBK
guJx07Iiaq4JFPSisARr/UqPCygXFn42oPrzsN53voBtN2yv8sSahECKZDGJAQvQ
zZ0edj+ohUYR4lGvNj330sekNsc6RsQAw+vr+x1ZuGyJYGcnkxMD1AR+itzz39/9
CJaER/bClZQuPPlHbzHo8hPU3sjRrTbCQf4zW6QeJV5gtcJlbR5QGZa1c7ZBEJY+
gcF7VBpMFmwWyf+40MrmqjLdQbCcoeuSIypn6d2TbdHJhZu2lP7kQt1qvCbbVLib
Xltq5J2OkxN+IbdH1tZ0XEYNLA7vLUyCKLWTo5RgzEtoHKt9vB7fSrae3q/KrpTj
bmiMlUBIPULo72TgPbGjJyNbF3Kp7ea4KwA/UQ11yvwu0S56LGNy1Ti0SZ7ko77j
BEnD0vd7h0qRZqZ1uYy2o/v2XC+obqPrmGQiKhGjDlIBxsAmhjWYiP7B9oAOw4tM
BdftaKnlFjEeEIChCQbTmK/V9ONJmwps4RuJbPE8xrFOl/i27IrR7DM6DTPA7E40
U7U+0nqWQocuqKiURvsaZzBwHE5uyZv3zn7++v4DOAuIr4/tQ7hfxFihFd/P8/5z
C4ry4HiHbyxVVh3JdNMc05JqRDl9k3B87jT85JE5o+v8QJczpVL/XhMndQR1+7UI
SFOxJBi2XrwHsSKiqTjM0utTekIzdcKSlLcheuJ5Qtm0KoBmjedlvmu/aLEwpbXY
tKu5tVAMIdblRqA6BNLvAFfoUzY81AOhWta8nPJhL1CjR9TrsAOVUIgNbeyusl1h
9acckYhE9kJAm7nDG1mP/hup7dE+yPMlm5wSvFjK/2t5CGGnRtqb5AyFCBK15VyW
PmI7bRAp/QDVyo8XjPpO+vxKuWcbxmORguWErJJywGwkWB46DqaXF7caoz+a2xd/
J0EaWzAg4hldd5tA1JWnzZ0RVGXUByeGzU8deJ2xqiSQsz6t/Dyw+rEVyvg7E1Sf
25+lPiFjzcq3rWmxlUTOeCnhJuDPMvPAPB3QRItvxDZXHVo5SvYdAxfNcUj0hBJV
nV8/Yng9K9lOyYtct+cLp6aRrr8db8yXJdJ0CEedkbs/aN1Exvf1OhoP/2+hHrt/
h5L0VdH5rzA3prxKnyz5tS/uJci5p7MUNDUpXafRIauBoDszHlPrKR4alt7j64EY
jwQIfZiKa8Hcq+BZiWkBUEGNrteK0XwNOIJ7ieWnZ8QTY6JKTdWrGiBq0MUb8NK5
Hc0BWqhxk6EHmsXS40/MLXMShQWru1+1do/6bHoDlmmnJz9aXRKFiKuYidbPdimJ
ohPsDL+aJ4zgytIB7QvabIK5d7rEeCk/EKnxvjPCz6iqHvSx24el7VSHeLFsCXO6
gPzB/fSTgg4ztSX+kuZVPdYR2/f0EljLKXvP6l8uAgbHexo1BmxIBzpwfWuoIAQP
JtbKfjySLSCgW43WsyiPmmee7KumS8YktEsUIrADtFTlmbFlEKS83ZPQojW+rJt/
bC8dJJYOepS0BaqO9ib8JhQkFhB4jRsZXUAYcnkBGYRRi+eBu+kTqaOaJDfVyxo0
LwN+0UdxJ5dVcG5ENTHsHnDGnPRdoN6/+KMbvM/GrEhbgMocQhPz/0NPRHJqcjri
uEwY6ZuLofCPU16dA9H6FbBAxO9jCLsjiGEyk/2Zm1QTmuOWZ4+x1672XB0n3R+i
KS+HaWr2ydZbJaa3ImLV71SFiFAm5xIu6PcZy5DfJbERe26Au8ttdS2gej7kVfWv
GdeJu7Qsezii50cxydUrXq7IO8MFfNuNnuOYktZ5pWBe8heHIiM0+gOAVHMPv0EM
vHNHMSZjxa1gHul5v4OY08Pn8345z/sG2OkYa2v8h7SiEvIc1BqFSOHUxqU6cOI5
WLVKz4FID5AdWMUDMYf3P1ISW6/A7fJHsvzHjCOtgawPYBH8DLdhs6+riRZ91vni
DfJA63/aKQx3roM5JLFsrhB6nC8WUTwdf1FfSxpfgRjOUkWHXFNsuKrJlWLhfWtj
+BAIDz0FeoIWcCoGX/uZiXl0t6j5PnHWw9QjqkhS4t11lCCfQECSGhQbn78xyCoG
rjtj0q8iNpCWohGEaoiQnJiTEwu1U8dArxMyj6aDWT91ynn9mhokbu3aY1UiMzii
Ci1V9j3dYlOa/tcnAH7zbdNccanlDfwOcFJluDK8si7/tQsTO7s9rnI4riUBu12W
ou9Mi5WF4r7rTvHjkrleor80xrh1pMeW0INBko5l0RJaLSJbm52hv276crEDbcEg
iRn9dykMrE9F10keDEw7nUgt8i5sILCF1tfLki9JVHVftNHB6hKcaZtkhkK2Y3ph
q6V29In61Bkg0bEsm2vgs0t9KGjwMZS2FDZWEW4f64XmVdJea4u/TwYcvrOzgSou
yXDrNzpX7YzzPSyLZpPf0nSR+MV0CKjLYRZjmoVXpNvYPZPVqPk6xRTuYLoL1kMx
u3TFzcGEH3gma0ArM3rmU0G4e2xUiqNFNQ91WV/Xhce5Jev4izeLJiC3LuWQevFw
XDKD7xRDiKPRpCU89pgLvJt8eiSIXTl7VNunCH2YXMLJPwcpQWxV0NzVYycXLrgy
2DHl+M29KbdP+NS1HbpbsIalq7Z0EdUFPP0ZxurBAOn4gtLUtHpAWif27J22MvWp
uoknU/AeoVyKEq+He25WGIvGPuwfsvlD+vwuFKQ/uQ3C69zam8DaxQqDVYUUvkTY
kQ/wW/QNpRnodA/QE1FqBjqVYmdrxLpenEEeVHpKUidAKYqANQ0RDA1sYITa4h1X
Flnii28qQzUjxlDbAvN4hGpNdH5x9nrSFylHe+ttYJZd3c1GKpOjhk7aLu3tiz7L
6HlcIVjOMD0D/aEk632EMQE6ZAINVYwIg/KDsb4OYLcLzCSsav6dD2zVu2LOKH4h
fG3NlRm6ujhCpzIbxLHH+4bG7OJ7lEhXzgk+o/MQEaWWPzQEjSL6zphg0hZe6OPF
eoJQoUTZGjMG5wboCSFn5OO2UW9wEalBlI75OVcJTAZo1K3+aw6QpKAKPXn2LtC0
XjlVZpkyK455h3v7GJ8myDSvLhXIBEMX7K8aqD20oIZY+6rSGHHiLhcGTEslAl1f
zWEGMPo9orVATmjVOrONGJrj8ul3nQeTQwPJhQ6bvscQym0AHYQn+4hN9DboZjNf
+GfbDEwIGGPNh9SQNjk/k5QQk1mXHlBWbK0Qm3RWuKgDuVklXHmcIqOrv/DgUjMW
/UfGVJ5y7WdqYcD6c4fay1Bsut9+xubOPIJM13uCoQ5xPrlo/zWQnREZ4+NZ84Sz
H5xlYcNpMl5YkjSd9Zx3rvf4njzE8MYrc3xeF4QmYn6MghbSEVgmLuYQ+5TUikI4
+bz0zDkqFMdhPSi7gfRn51TTNom2MUPlRrbCIoeiLJ455+NgqnxXJmvn5SHZ0L35
aKYLl9bpQ+TfnR76VT0PHuC48rlAAgSIRJwfMiDRsXKmjB9DzJggRIkVg+FzJ79N
0su9ArO0zxsiOqw6Qu7crTmD4G029x2IcAPsWi9vc/3ajkrbovJKEUNYkcIhEHhT
7vYgvIT4fse+1PyGTn/Ow5kWf3d2jt25ce32Ca2ABV2L1vvQrDhwXTG+wLI8lNQE
XV38RrOKKUEaRpJCPZY7G9fhRMEXY1ysaoJIDcYsq3t5EsPf1E4diWSD5zXyvdu3
xMgVnylNDhDpniRQH4x0D2YAzQzZgkYkhAgA+8Ow2bWHkNFUXnJ4nUFVpY551aMH
K1oq8MxLlqSzNhNSZlNxrr2fsPVVGkvRMIweUHca2AqaFYV0RPl8GJV1KHtC1DSC
cZMvpUgELoBBkNoo/OMcDhOmKxVYLCWJ0lRXOLJ4l+bO3NizCOe+8/caVGOgwEVo
c162XKgaLFqxG16KIjdKsqmLRqn3pZAw9H+BTDoEw/KnsgiAEKFjVwxT21CH0ECB
HJ+uKOzPSLSiXb/NOVq1rGG336hbiIqnaJybFgeE8iF9o5prbsmshotAALNWz9Aj
/LO2DoMsEmo1nUkZ9UdVvnIN4QFMN0KNqWpU9aL8EamKM40AshBm7NbQifGS1ACz
A2b+hO37HfpTXCcrc17rlWpV9pFJAam9v7JrGPpdwL2xIEOspo3rC+8idD19VkiG
qZQSb0wgUBo4IpLHVX8H+Wc4/wnGiFQJAIMTFTVr8D7NZG3szJlvIXak60d/8ApJ
Iv5F7VOsU+sjOgJrvuiFlcpKd/80bHuMFTd9pql+s7zfk8cW7MjzrYB7a+XqXPko
jFKIwwbWKg7BmRrP++hTTjYMoel+PwViAt+C0ePlPzC0tUenG5XKZibgaF9ORK/a
FfWdnTIQhG9/v2zfNYZb1+4BMJZIlTElYru88yuTvaJI9oPcgXxhy7Mi+0xLVu++
ZkRHsI3VPYlFGl+GnOaB+SorjbzN/xut3iQC2zp6DhyoQnBXOeDj1EypwwwKuvc2
oL189GCFeMQYYUpVbCtDepTyv4RosM1zMJy52CkV58SfU7pdVDjHAcHtIlC7/eJC
S+eLNpdOG2c1jSk42NfH7BSVrTPQ1syQ8Mc13fcaTxMqbx+J7LPva16z6je+zLPP
gEuIwxU9vfWpb1ww4KafpuuiaGPNieVRmHpyXf5LrEPC69uOU6ck/en78MRrZNEe
HlhbWLjfelhdkQ5nHkZ+9ymQ7LUezaUC40e5t3kpLhRVBTJ2eLhM8DUA4eDU9IsD
bLypk0UXTL+OpXeUyFtaMULyUajEg+yuv5Vbe1hhbi+S/vmULaFqpu5M/tcIK4wg
nOYBxXxqdXTJ/E0N2Uncs/shz1HuPhVA9OV59C/JT9/nLkNxHGTCa/TJxemvJ8CU
zsvDHIfdqeZ2Wz6RdXGmikbzbkbXvzMkPxCRKkbFSqYZbx1hcCVrO/ve6g4LEFtG
s29cVjiEx/RGVB1HyWjpq9ZGY++3sKTeAfoTRVA6uNAFLeAaNTx9NEMdLasc+mO+
t1y4yG/i2t+E5sno75ZR3lH1hVEwfjlJKMbICeJReR6AtX+F9hk+Y/Ll1LTAR3ja
ixoLbQQw3kidxIOKxgCA2UffFy2x3ZwxJajaYIO0phd0c5ODonBS6gvSgSmGqVKk
AAOK+r3tkNC5FvG1FQegRxXPHHmtrXS9UvfUIO5Xdomdj2dqzihYnYr0H3uLXiaV
ZjGYQSzoCmsS3W8cRAo1gw9fsyqKlkQxh9JvmxLeTaYDxal4MUlsBERwNsZov/OV
wWHyc8/WJgTZXKibzNGebhtW/ri8Ao7Mtw2B40wWaP8JIv/rzYNRpbwsK08uXgBK
h9jb9NrCy913NtnjKyJ3QhRXXCf2A5jcn605Ows7UWep/UWJySkUJS5uc33QHeC4
ECQQXukvG2oerrIQJ2Ci32bjFYUAMTzP6NwegZH4PMHtNdxIqCNuk1Ak8JwdReqi
8lHCoHtiQ/sS3Wfi7Edn8+ZAJm1mmNfInFHsHGxb5vPjVkEfgMZpG5CXOCjPsF+Q
fXO6iY/JmxRHnGLFY78i3O3WyiHga4e9WkNzfB7d/7RZ+AU6f+JxDTBgaraaOHc8
JOVjt0saFCWMjIayzqB3l6u3eZNDrzQmQl0a9z/Y+44zmh+4ZUWspfk+x+r9LbsK
VRXWiSOmSHZPzOTZEGBz3XInaGyqxpNUiORZJMSdrJWrF3O4vf7BIlKbcSaCsBuL
kvN+TkFiaxhL3p4fMiAcXyUEuaCYGMVMyqc1X5euIGW4mhkJUcyS5L577Lp0btSx
db2LUtrJt2h83nS6r2pISV1r9AJwyu1sDfyzhHsUdl88RuzzJdTXF8CaUukOHMpD
bDg3Ug2WED5T9HytnK5xRmrk0htMuD+jfy0dbzk3qCRW7SwxPq0ZMVMsZqlUO6bp
2PZNU55O/2oVhZaMo3cR/1W7H+5qusgbxBBfyJl9ewtEB+2DtYDKBg8NH4Toio66
zWWGsugbTBfLUOSf/m5kKK44ua/r85abvdYoGXcvgHr6YYMX7i08MPBgHKz6EP4h
SHS6h19it4ZRlhp2xCvOA/QlB4+sCjGrrTNfrRcr7WkvVrpC69wZT74XtkpLBBAD
vPcf1nIuw3XAoWf3h1kh6/LA7aSv4hp/7u8Bguf+xuQ185numOAWK9DSz39AQiyu
EX1Yh0TdJfB3qw4me3R3ZOQqim4j4/1KPLeukymEmdsnjiFmj9AWt1Kf5nYZTdmF
wpciF0sR7T2otU9VsJ/1JQDPRFLA+ejyFhkYMhFOj0y4kESS6z6wiXroBbT8fC0N
AEeZrvlA0SSzeX3w9TUDKLMudTr2dtpxHrGphuccZt+TzyY0eZpTzrEl90Kh2x2C
l6lATPC/H+rPYOcGDqMMK253oZDcSSEyJrbKAIMEPgrZuyqAL8JAZUYr6YbTo/EV
mgqMAXyYc8iicct6BylFvhq10SOZO7pIXuQ6rHEPNJWdgMYI5a/+kke4ZdTfIlUP
qgC0RSHfKozsoDNI7FlyUHHLki/TYkW5NVEGRi/O4H+yc85LDjgwHZElZqDr1H2w
E87YqI+CpZMUVU0/L1Jdbu+MY44IMhdE+2Qq6g5AtPmVopsmh/wAx+ztnRvWMsGW
aVeNQJWm9UHA5AJ3h83Z/LnQobJ+m/qXhIwsTMXow+ftFs1QI3YdaJkIA8C1JFZv
06mNdU1pG0KCvj13pspoUYuYpvyocpaFZ2frw5LY/BHzgJW3VWP1/3WfKNVd8T2h
RboiaLq8r18atcQRnjk6nN5cZiEN1hB8QaQeD7XWESewvPrVBsVZfzSAPY8ieZqo
0NDQrr0kLkgDGu6JuZoRyvCO+lZno47upVk12Mg5brfAiZ7Adrp6bwFtmgxs00ll
fjeDrAcqWIa9Fd0jt7OaHYKdWSOgrNLEb0lulZP+vZyC/eKMTuD4TX/et1BhaNzP
o5iVSC2AFOapPix/4bYtcOrk685NeubinZ3Yzpv7K/mW40QchCaqT79dCzX2mRuG
gikeSmUfsw9CJBaUeTMU0spLExSTP1RY4GrD/abrB0bvG4VxnaH/tTRvLCVutxlf
cPSMMf/S8sLRbMC5HPNtEI7UP5vJ2yQKkBxR9Xn+iWfc3RrqIGAyW7GSULgjxMpo
r75zkjfWtz5r27GEoqu6ZOKBH3kMqaapoVDAkPmsWZaKvmsW/lbzrVIXUE9uaN27
VqvuW7dPeoS1gnb7nYUfHmCZ+iDUXv1uZAz26Je22wpboYt0rj8FVsyPhiMfkjXp
X54ZstRqZjcATyN7smuNotVK07+4ny2c4MXqnjobO8YnGVUXZFIDuMGRbXGv4nKZ
39r3r8VUfLxE9fo2mWEIR1H74vGEnML0kezu/ZIX4AgXrOfwostg1lHZRGt5fTkN
PgrEQgpMQ9n7bmLsHbNE3t5/w5hFUdF0J7LMYDsh9r9OhnB1aYjWbZ+QgV9uKl8Y
rWTb0zawbzSCI1vP2DAZlvt2dzcLU+nT76OKO9l3YEPHlSBQMo+3jE41JZ/UiRAW
shgSPhYVDA5sP6Mlh+5+o3d/BXWyAoYCR4+0CIdCl/Ljq+3eJX///sV0+t5A8/Ls
aOUUCQQY8/2r8nkDctOyETTudUqHXNhEDTsi+ZCVEXZZj9Au1AcgVvCRyAKQViz1
xLw0xtGCb59AnUrez6lS9IhCgBvCFHZGd7XbJK4+L/3v4esIQ5salEJ1fM9VD1pV
OSgqmTRZdfq6XJSMkBKE8dVb3z+gsUfX2LjmFy9FQwo8lqvzOp09VyArLG30HbGa
xrsDaDHYJ4cFyM4wdmmHjvXneNeJT0L9aCj2mFaLHuH7LP/vuZhBz9rOavY3XYTN
G5sr6hOqd0QgpNHOIDi/xMrXU6hr8ZH/tr+i+ARQqRHqTsEz8uA8ge6nYbr38QTX
AxZm2e0lZerLhmIrHseCLCfFDsNePGvH94jtVvnYI7ySp4SSp37vY+kD9PU4eVTT
2ButMXnj6sXsj0DAi9g5x0MHIVNRCj0Sze1iulcBA6wKF1WXEtQVdh8yOsNjTkU9
HGhtN++AzdOavYejHpesY3GiVV8hbwAFJnagD+3ZBZWxjA5YmL7ZtvIXMBQ86Tpm
l0enDcLOhGtG+oOQ7Wgi2aWNP8SyeNKXIHpSAzIWt/PSC8xKfqwQR0kWGQoxeeoL
oaVLja5vNTCJL0uPl/n9nPnTR3thSLH0OJ1xDt4crX6eLhFjv8FghHys5lfRlP4a
ckuMG5OTR5xp8FDyYT2wO6FYSUKKWxpnsBgIDJIdd3Sg7nDtrxMr4N9ECgsko58H
WXC0QZ3K3LggSnYwBGbiDXCkyrRXL7k+y+PvjFw4jre6uccKGKUH7zQk/msWe141
3Uq5zjbfF9cVLvU91htzK3/2aAwoM/vbxf8mizNBNXAEBMS86r4zczikpt02go5n
egD8KqhKXCkW0IOayXl/hY74iwkzrbiOxRMGEHcONq6bkUHwcQ0Lhcic9m4jlMQL
ySys1ckg78e9Lh0jUZDRmKMSAdct7KXlMhlYts/dxnpVTJvg+lfIYCiVtVvY44gK
608JCpJ4Cqzxnm8LjQY58zNPkB5z3kxPz+u9JN5rqdLwqXmcipGI1hJ3k4y04/G4
KVaAZxpAYZejiYgR9kcJLKSTuFuVPqvuMETiI8m0FNxZnf++wpIaHHMwws34TQXu
hbkFfaGl5pII674B+z4hjRRRNtXfh0qFM+WhYjaZvOUyT14G88LrXV135ht1Spw/
wltP3bDIDUSLLsPd0Gkjpb4PbZGMfXo7QqsA+MMc/AjmtLiLxxhOkz0XOZtI9gpE
fb8JgEpIcnOzlQCcEr4mqkGCTAswJMz24J+VaShz3+lZalOiXLAqxkZ48uNpP74b
x6fOoLxj1tpU8UUQWjEDfWOKAQt5EfqgVzXD5j5WzlBQqBf8ntVSOIZehonp2JiZ
fyJaY1ooA/b5BSzVaT7ASziSSF5Ot5m6TwDfNA553AKQE05DzrW9jBRVDRSqif6N
FNjMLiieOt5QMWu+jTI62WIjEndDs1PdPlmi811pNRQn66TKEuH5y/kmj1f1WGBG
mUFiU1ibxxgV9QaaeX6C6z8ZnNL98X+Bn/qD+g56kQ+RUTDMiLmL8qpgfyVNhifw
8y1mIQwwnhYMP4HxUzPyNu6b6Vxn4+oy0DxOgmS6eB7fEuItTg43QMGz5LDO2BOq
7koisQkSMrSwLg+Dr0a9DNyo+DdKL+0KCdlKvptQfwkvlSFwizNfSMwofdMbD5wu
7AltmunpbVBKOTSsHCAr8/0c9tbCGBuXgLNv33BScjyuIhPJiGlO2b60b3xNkMk3
lClU1N3wfXH5D/cSn065sHYh7u4LfZughJPFtz4FkIOw+RZQ71BTMHJawKrDZe0E
D779bCEDWLGMgexBUaT36WJWTZrJLm9ONR2RblZkSiAvvbyaEW+aDsI0Njn/VlIu
QTHhfD7SZsRYBxEetkYG8/Df3qKhcA43Vi+SrIWnaWzBxIIkNkCnBFT8AzXIYyO1
bCWS/c9ykRQUU4Hnw9aSo8gVVqKX2esiIg3ozfd9a0wGR/mVJuR2AJr3afgDtGl7
mnKyaJWwW5BU9/ik5uu8kcI3zVO52CE9m2uqPsytIjlac2Y4QePevtIuOj+0UN3k
R1/LP0zWg1edgT+B0z0rIF6aFWkZX0efBZM9Q+SwkAiV3w312rooqykMdhfCTf8C
gm1/SIzC7RdNnd9vFdi8hd/Y49XXJtpfakKEQfbdf9NBjmfArMmeJ8Z9hDHPy19M
ARI9qaeVBa2N8bOEIOrLAajcj1WPIS+yOGqKkzYS7A+DROcVytklUeq7C3ue6S1o
s/zRJZpkyvysTCGHHvIcRi7I+FFt53KnXs52UCPARAAAEcI79vD6SA8dt4EoW501
/Jrz6Bc8t7TktSa1g5xgLwrC3A5HPLl12mpCGIw7KCvyfF32Nqk9TWbyHcEOC6Cc
2+Tx0jRBmk+/M19azt0v5qTH8dEHmF4mj8EIRLy+adPCccIk65m3UCNClGu41syM
NVT4uUNkel7Fg6mC1pb0CjXPj1QWfUV7s2II9vq2Q5qHIffEj8Aow/GspRLuhYTi
pZ7os5sDtBmPxGjuEbqrEOK8EbDsmKlmldHH/7OCqkPuDipZ0TO86Ml4T7y20oSf
vMpEgvAeddkDDxgHT3ntI7QuebHvnb2tyN5HrUBnNwXjqxLUCdEAIjwzCNVZCIRr
3e4mf5iy3bkUJNpsE8hXcEHhv1OQhmHwfK1VeqDFQnOrfFAu5Sf3GJvB4M+rK6+2
jkQ++iwPHFCJ6bi0uR/fYkSJolr3OgNeB6SgtM3QtowVLpwvcErCWOYOKuTIklp4
3CoDrhI3LpeIqEeqVFL1jOX57H7Nls9PmMG4sGoHdAKjkGGTTASpiB4tyZIXTan1
328mxtekwKw+6zLUJ4VTNO/BnNFR0p+juTKSa5IOf5g=
`pragma protect end_protected
