// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:39:13 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
J2WGCC5f0Yfs8kkiG16sYeGIRyn1VW7O2m7m0nRr6FAKlwj/roPQ3zJALFQ6Q3Qn
Jy7k3Msl+D9BuiPJFQahe8ZuYa/3NvmZ+tt3uCY6C/7XzdQnuXkzJQjD2G3KmIZa
tY4Ql/69PP0T0QjVn+HPq2nnXaXbnokleoR5Ra+7U+Y=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 22144)
jki2SNnMiNln7UsyP8SD7sYcrQq+Dfoz8WzwNigNMh7yaxU5O2tUCO4OmVOPRoVw
p3/XeJAS77XCJM38USaO/8Onlbtj/4ULB0+JS1Vjo+IaQHRq+uJHuNcUnIPWOLBe
JjesbQgmDnDif9XDYxJCQWQnDuFOqOygvcUs2Nw3OsQz2GqGh9WX5jEx9oLpswms
galaKOiA4NJXbzec5sG6VToKXVH/gVdqPAneg5bhY3RzQk6TJ5Z/qcmEO4nYiv20
BqeECxjUY2SV4Y+9ely40DYeHBP/OIGAhu0pAta/VZ//ml35cm7N4EdZwwxdpJLq
GZeSBQO+ZbtcgD+oSUjB7RPI4pmasoxBx0SW7+umQC/wXH1InHkb0sh+8HYv6kvi
AN57QYG3y1Y/nLKCHD8U8x/kgqE4qJcvlBKR5zbLB01a5RZV0L1hPYWWqPjOYAlj
cBYFPUsxTUXm0VV2/+ANRwptJTVslffACtzvUP26q/FiX+IHMfIrCX7weGctyRtg
nDYzeIu53pvIFoKVOvkCEAusvbRTYlsEvnG5FxYzz3OqP+eekk+TIH8oAmFL+Jq+
mXA4JThr1Z+dHfWWRUBm+wc53zDYJUIcLcJ8lAA9VKZV9Xc4Cl8xQ0CY7Q7LA/Re
QVojO8UkM2Qb2Z6SKE75e5GBFntTlTR4JMctCh0eW39rQQbA22o0FOmCYnDQDzTr
ii2bSBp5bgti7vThxdckEz93LySl0QAIpG3Jw2E+Hk23gkVzo4s2/3z3hBQ2GtpN
6OtJGXiXUq8csC4kTQATQzD87WFZiuOATKhsMDBDop7ONmVtg3v/t6VQw7GZu7v6
drddpxV4E4bf44VgPdmzPh/M87oXrgYpf3B2k2y4cFjNUxEySEkVPsM2MTfB+D6W
OHV7R6eM33DPEJ7PEq/d9vjuSwps82v6Xmkq5EBv1JewyF5KDUNAxVNXKWxjV1Vj
N4IkIqxZD+1nxiYjC9gXKPVGV3PHvc3zxkTwgvzL0/bZmnE2EygFAa974CAfm8vx
B9UTu8Qp5pKgPCPse/jlYxDuKLi6Iuh+szR1blB/yDIzJhquH0jGUXCDfScY3R0e
iBzLGgHk/Wj4Mp8iXh2zp9DKghKvAHU2cVOhHZnRheGBhP3fB72fIQJbAMGIpIxs
njibkIk9t7921c1lWXbz6UGSnNIlr+JsTKALtYZ1zI6MI2mI+50sR0KROHLd5Ift
ZuHOkRPZ1PinTOakPg/QldZKw7eB0SOiQFDWt+34l6RhwyeBvgR7ii4q0+k04syB
GDUfYk9wYyqtyJQ6K2ytmNpkpB4NlqhZu2bF4sHQsp5Cdo1HCbfnq7qW1wW8qdkH
Yx3HdPIcdb/rfTFbdSZQKYlrfrMW89dXS4MjX0nnpOy4gQqRML1+SKNfBFne6Fd3
/RxEfuytaS70rUnbvtrfwMH8VQFrLCJpH2i3UlM2rrS3tt3lVNiXdf3I5We1CZNk
T3ofeJOr7VR76YIac1UuTvouPEQp2sQXWuSOSAizC0T7XCptm2vurXSvydcHJo+x
QRnP2RJ8A2VO0jAHrUzS3WAnpgJd0v7ihE6kPh9NwREHAhLeUBYsbsH7ENfOO5fT
caOiBpirX2mnPb/BFJf7/tXv7Z5Wr84hVPAzTiMGF5MWYV9CrK5Mxzn5tmygUTnK
FWBA+lNTcVua1+yaWwhpreZF0PPqxPmXijvlHCNmaCqbbSECAUs6nhti5piKBQKY
ffhzqcCKKDfS1GZf5D/Dpfo48FyppUzsabzZS0QjC5GSxs7UduG49YHkLQYH73C/
UbBjCiC3lJyeKr4F0fvjQANs16Mv8MHSfbZSWm392KFMS8ttK/YN2JY7jfMGNtnJ
As/9qwDYB6fRqDWPeHI0qeGQAenW0mZY0Fvyv2fO7YjTKcd3ocuLP4RlpVNXHXtm
rY3WTofTUmu2+q7dKLwO9bpYx2HgeMiz497eiA+6UFSwMZSSG6HXIKo8e8XbumVj
zWEzgvYRchXFD+c2MlLfYDJzGha55y3lerbjDeG/y1i0zZ93OK6B9JmKQcSal1Ec
gr45lMygs6Q3vbp14ZhYZEWS9j0VyE/luXLb9XIOVdPrA/IUJjQ/01WgViYUP15U
n/uN+Wa+tmmuKlzkCOgTeo+wMfdDMYhm5AcOFh7G2MOeDd/weqBWTv6w2Z1lQxy6
TcznYE19BFVGB1dUC4acZ4N8w1H2MRo296f4yd5pL6dGdWG7nsqnhU6IA8NVeaLy
WJ6YyEuX0D/zPsmt++vkdLD9DZ8QS3buT+/X4jkQpppBJUMREuoikxz3SMkiHZdQ
eX52rErqLMWpT154sWG1zxkAMxVHLEzuSkz7BHlhEuYzTcXdSQSmtm4JLNqF7Cbg
cyQoKg/MCZVsgXZH5EHbbbLKjEf2YbSdUoM943TqsCdn3Som4RvoibG1Nu1fIoeW
FwpW/zk1H8605Sjh58cnz/dTh+6d/F6mYW+oorioP85VJ6m7Ot1O//CS4Dq1z2O8
Lb5+1TnNT46vKorQ0fBfQuy5dHeltqPTNLZcOdzbHpdoltlvl6vT5P5l1TN2AZ/F
qe0vdIxubMTyCTqvS4SpJxpqekBnopA8AxIXZHzlsqFi5pJIwNMRwV1jQwXrJnG/
dya9LsYTEjZBw6Vfj6HKQ0col7Mw8Jv0QkOubGYecYZgNgZinC6XE4WEWs5dO95q
6UvoI6e8S+ceNu678prhVTm0tdE7agPUltHh6H9BJpJDrO0TOM7ImmexiQ/Z1X5N
W1AGIyun0r7By1lPdvOo1E1YDvIc6nfgUYRjoGFzqZM/jXaSLxCo5ys/dxSQ4J2l
uKnv16iEfjGByYiNal/8F1j7GFqduG3jS4NKeZ3yyN85VQA9h67Qy3zm2pqqvMkd
JRyHO6E/4oCeAk22WrxEr9sMWbt/2FFoA66LHSZCi5ze0n58yu2Tn7gny5pzzf0a
LmtPeaIJyaUdginbbk+YYmyum2HusfNnTKy4QhHDcuYAPqp1TGGAOEN+HBn/t1N2
Ge5li+sd6Iv0hLME3aL/jKk6oVJpHFZuMHoP6U9vDOZGPXlpHA7vxvLStXbT+JQj
S7+FtKZL6KCNyU1Uj70LxMrhd0WGKeK+Qlqq2aqkeMaq6FtiSYOKMsSqvnfL+oaH
428AbZKZv7KBezpxPK0tnjzyZfrYBNhfQn+3CDnhLhHdDl1yt4TO81ZSbxfe5TxT
KD+ZPY0VPvutUsjtYlqK1Ptdy67Z8xeLjYTTVLWabctA6Qokczjv8PcYmEJ7btnd
5hDLYp8JIc4D4rv2wdGyb7+ehOaWghyRaOkJB3WX04terslf3gcNy1x0whyDL700
5WLivCADynaN+EYI1FtcKFhtwpRUJ6ljBqEI6xrIe9j1K5lgoEV/8l56oU0PWeTW
TP8QhfkBxYtbi5JbjckMxyBZAnvF4IRvkMQ90uRdg2ERsAeThHXXvtaUMl2MKYmX
qzpY+1/ZnjA2oWRZhHtfwsrFwSCuuSshe1emRiiRffYmZwWhB8x9ygciTcWRfrJK
xJgTpmzAsD/JaVAh86zYkSW1bjhlLsQQkJOg4wwsHK3w+R5JkGrJZ2K5D1enC7v+
u54t1gu6Dghbe2NBXD4NkliFP8v3oQ4exwTKN/VRVBhPA5iDNuxLRpp6HRkthSuY
WEH8pUzMNlGL84RT5cNK1nowGKvZoG3nW1NBKy7E+z6QzzlxFUH3Fz3Kj4AjRD1I
icxi4c4BuYY9kMM1G39k+2WLDWOhu9Qua39adtA1RKr/685/U91uZhbxdzcUu3l6
A+fRfCCUxa7e5GtekFvam6YFDwSNNHaI1i6FuS2NR75kLZ9p/0OR6qiA5sK4KI/a
V81pQ7vg8rV6pPyBrlNQRRrPo+x30PPQfqM7iwDUq5ddpeKIgoJQ3k9pONnWNeMw
TTI8U8E+NiU9TsCJAXTem8FLRh4Co9keXsVpKBtp3JoLTGxMdGrGl+Z05GCuG4pS
qtTWXzCemrrtC7awNvNb0Oc+i8/MxjR0nsI6H2PAwVuVNIiAmmppQWLabpvhWVtF
RyUvMFAX+oCs4hQJHbY92UYAY2EzuBqo8QscvONPY1LJtFLutrBYlgi8LNDPgCpK
cuNHSP3KK3sm24eA3vwNyeZTGeEX8XJoTxGpElxAeOqt4k6S0ZI7yUiiK+lGybHH
SiJ6NSBtVlmbeprqSfBvHAJ/c+bRoqw2HQ6zsox4eQ8tobp1+7XrY/y8XSGovbog
SBAow5HvoCfGWiqRUQL2Oo/PH3hLjSMP3q/bYL6u2hUye9LNZZUN7Nq/s71B/tc3
cVEMwU3gI11WAxWhDeFH+X3No/la9nA0I807n8aBOxyXPyEkrtKprTTNe7FHHVID
ubHtjwW3JuNHDwCP9c2efaVc3ecg8TYBjtHzKBLjSkkKssfbdYx4xMpfuOCN2s2j
bEPGbeYzX0oRVxZZQd0Lr8DrQnUNoe4q8Wmzg6dzMwwV+Sh+rt25aiiIgolpKKIM
OYQ0vbMYmyaqd+XVj5SujoAMpmzqHPMa5lyQeFRp1Y5oNWNUdZxdXOIpCF7g6d/I
RWiorHqs8LoGS66/0pOyI2NdTnGxcjIDRQc1mQoXTXaHPGuCtDi36bkZN5fLbOU1
tABQtnFBztCDqV96uK/FmZRrqIk7oQZE0FeOF7bQiXFif+C1vhlQEj0O7r4kJe8l
+xQpKMvfQFiRkJuPhNj30NMRCmI0edWbydKm3n/w6CCsYPVa2m0U/yRt1cPmVlYm
Sa9VY7M+ztj37vyXJ1Z7WL4lWIIihvLhjEwwuNIvzcx1m8o3m+XOfncVBnOksoAD
l0q08eDXT+aLlwT5pVIRXKqUO28IQdfPDVQnxBv2SdpQ2+iU7nxsXbt0/HS8duIn
04XOFhJVfxD2f3O8rLpeylDlyp52MR7BjLJl3nKj2ZfscqHyGsWHgdSAJWCszIaS
vrLDP/8HkYC4esHFn3a62m+KyxY+sbTNT6LGBmVsHyWpdsPw4IHgeRVfF8c8jLvI
THR1X1TLAMNJHFKLhG8Ny4i2vd9P0B5y9muN21H0o3ziyGx5C+0IjD/KatvkOYRn
3XEe2ycovwb4J9k/8xxU3enNfAA8vQXC2+PvZfh8/xabcbsGE5thAgxyDMgzvQ7r
IWlG5oiifkTF+N2lLalsoYsIRzRpLVawHKi6k+lxJ9/DL6BIPWVRwVRf7vAQeeuT
mZ97JBe4cdutMS8+WZ1ssx6myxvQYO+UuFWH/0Yla7HhYKm3fq2qvJAns61xHU1V
rHUPDgClF9vYgc6CaOMuaYcGxIa4cexQMgYiNryfR8TN3m1rjJygvw8Fp/PmNJxb
18sn9svFPSoMfKbaaLnCjPmhown0ldFrSAIKtBQQhfhGXWcFRJy+BNEmldslyu4x
6SN52imOeZ+xn+5ebeb47N8o4OmX8e+Vr3+XR3/B6te/RSjTxFKM74xYJhLBtQzX
mNQM5vtS2tALcYgguVrMsNiSoRa8YKvNhD98pDGK1J+lqmAciv3QzOaddx0hUcSG
pC5CbLocdQvPDC4DeBJZLzhMteKjDygYuVY7w17obBMmNQND2FxCOlc5ARPVH+5X
f24FG2Mf4GLlrD3hjHS6BVQPJgch1SZFmo2J+PD8JleCzo7axTjoIcIZuGPal+/J
aSkOz0TgxMFsbA6AuaDNjSk5CeCOWrGAxox8HnZKC4KWy7DMC/j77/lS8dwb0dvb
ghg75RthsdaNivpVguWGr6l5rbM2XungqeYoSk/6sCSaV121cZJS7Qo2tIJsWYGK
MbejD2RHSV6drM5gUdV36VRqWr5Th/moyMewn2QMqpCGllBKmcnUToXaSori040R
XAp8t2J2NMKr+u6br3DTb47pGHdSHo2MtFinKZPyXLK+zpoPM866tfvPke9ddS91
nRqRnnsYpMbvBcUjXdap+w/Pxu5El+4QvavPXjUsxXigWchwxBc/EppImgLCz7Y0
g/B1lY4mUgaL7riQES1Ig6J31O3oPB3gEDx/zjneovjD4wbOe6rPRj5vtmvnnTAq
uZ8vzumC1drm/9Qs5QqpvPBrIIk4qI2a0Pep9C7azWw+2f2wIUTEhHagLUe+02JA
lcw0PvqEIul6US/yMDyV0avjezKxTHCdUxAu3A1AvZx//PqAmjCCdmd5+RBmrGBd
3B7hACL76DTbFkMgv2770vd/JFvg0U3h/KzbQN17+ZVPHA01FO8wQ0/UYC94/QJ+
ANT0W343ITuMVshJE4aEj7yRx2fBGma8+fmW+g9r6IL0qRrpVDe1sKEpwOpAl1bC
j1DNaFs5D9tWfAWxOgEVcxN8VjKx2IBKL1Vimkv9Lhq2nUSFRaL2XOyU7u9b387r
PhaMqmMTv5TWcgH0Kx78D5bEiFegzUcD7lhd/v5DhpnODEqCNhW3vY0U0wbJK7IK
LOuYWuMUWAr9zJYmLGdLkxPjGEyApIkdahP26g7qm6C7Uv4z5ePmHk+Uixikv4rs
2zJM6nvonwRgexIc7Pkc17NFaryjABcT/7PAvqC3Rk3N/JSok5qeuU4SC/x/Qx3t
jx8i6eAQUd+c1yMZ1lf1DeUcon23v8nQrG9dQgcMNiNxhiwmqBn/nEUvsHKq7Cr0
zU9ITFG8tbArnQ+GrmVNVVc8r9lve14Jvgg/LUOE+B4cx6/bn5bTvVvPjIKv/D1Z
hp1tCTrWWvQyH3ayZNvC+SukqZM1Wdv7rOfSJM1eCXRoT0HqHfOPBElZvfe1Lzea
2PZaFFdW+kxWTGkM/0lz22USRCxYp0vk67LZc/ynGQZ4uJBHJnlIgprSCW1jKZ05
QWRe/UdPLeOIgXQ085fA6KRBciDqiS5EuQvkBI2x8sxn6dOGW1/pRolwWUU6TaJY
G4Qiqf5fGUuD8MkoSi+TohCmBCj1NagO2kd9ynNsKod/83P4NKW903mWAdIKM7vY
KuJklr/GwigESnJ/JrczU2WX/uhhmCI2YwSOkXMtRYSEwSCnC5ndYU6rrlSPBnxu
pevGGatmVRjX4xW+d3xFga//M3dKuqbPz5Ts0DcL4JioSp4/wJpbqKUKpPDwxEBB
ad90HtkWpDSFlyuhy9uuPyTmjncmBOApxEZnhXeg6164rdUpbrj4OpS1g0bNTYfW
zAdgAEKjAw+SW9FQ8n8S6xdqrtrtcQKzjAqzRSpi49TPk6B50r2LUdh0FZyAf3Wg
BMFNLXwAFj/3697Zq6XevNNO2UcUmzD25qiEo2sKYRQwCoPhGKJm5yr7catRyl7p
PMai95WgXrdk1ZeXJEaZuF3N5HCS4ud/TEt65w8cQRAD8cNrWiCetHao4apUjaHB
n00VRG4RiDsoICu3jDKsyfk4u+2oOj+rkT7R9bpwnpmT6z07nKBPP9v3Zyd2KaHp
Ttd7P2QhFnKW4+Sc20D5H4Gtd00QKQ7/lqb0v0YemOjef73QmSjRMXmEM8kWjPjv
b9g7ITonh661IFALO6Tc6D2Y93thUVhemxhv5bEuHLqsPBwwTLc0ckY02rKLoFmf
NrH6wZpg6znBBeD7UgS7vxFnkfh9+GZY0xu65E7uZXjehh0jrvLTa0kmdii9YIad
Xea2zf0hyoOgSJcM8C5HA7MhhhMcqdMOJ1VTbkOImI4mWk4SUDF8theIM9EcvVeO
eKj8RGLZ5Bl3rQjHuWjOLkBq6yk6wVnv3BPonGmRxSyfcrZbg51k8aqkTmH8OOIR
63bIw/IlMYvPwBoq5ylpUb6PXHCbaSNE1WIjTyvNE6Hd0rJB5Mh08+uTdQ+YCnTb
/OG7+hLCafzSy5N+t1BMzdEIxKC3zwnQmuA41ew2V6AyxIdWX8wLPy81DRONzCfY
e2MK188SYBXjbN7yob/wjyIipxVfsPCaHTsRuMweY63GWcyhH5c5NudJvu7IITx/
Rs9vMCJq2C4Z9pXtN2EDS/t4IOgpkveb/BI1aUA4B8CCkjrsA9REcdgPxa3M0Arj
PccU9Mb5MouqQXIndfPbLqP7rG9KCcUVTkgCEpctFewZghELI4l+7pFxR0PLCmvk
3E+rf0LZomjEorP3xsKwTGLbNPF94lEypF1xkgFo2r+1gCn1pVgAUgj13L2OhOsE
EudF9rELON1k/nyeZTp/OZ22LpDCTFmqzkQtlwIpkEkGIir9hsZvf8XuskvnQKz+
fL1owxsKO4mi9C0tjWmTc45Z2d/HZrDLVFKMCuQdaVQfXQAd/TAYoeGdk4phJ1Ec
pIw3OMRVvDIkwCpri7px5ZoWVG8+pOh8gJ3pkvl20cU7kuCbv2o1qwpfT12NT/Jr
TAKQC0D73sw/s6XJtQ+mXfUcgVIYZJ+YYePPqJcr3sBmUZqy7wLFH2lWk/8UNHrX
Nfog+rj3vq/pxm5KP/MxGdPeS3PEgWwIpmv+fQ+i91oNFbU64ioJrP539XV98Kd/
vY7NpwyYTBCmNahovipVxcDRBDdbNk78Vtk3wdctZnQz5cetUcn62eblV4p21g6d
HGGghnQgfqBYPbEwDFyTNqnK+j1GsE60e5vB5Jn6qU4xVt0DZHZO7a51ztQf6kSy
V+s5hS271HJYAQQIhXaIcNxBpe2KAD+2LAb6wXqgpASE/DowR4KElLYqvj6gbxty
IPiUccc8UGJm7Y7bN7jVBqygnKPLj28HMaMWtdc8Rl83f4fWdqror5lFStduw4wL
d/CF6Um+kPsysC02KPxMhvCjCIm9qAA0M7fMUeBNwE7UwpNLFqwZ/hJ1JlcIKmEz
qPdgm+mpEzB2YSi2AWEJOxRe8mY/5QohCZOktNZUTm2YhA2nh7iFdT0S7ZLXMiS+
JypBBf1BSo7GftvsUbPrkyrmh7k14Bap0dvGk37iI9YvWN/v1LW3kzacZ6cfwu2R
NorN9nLJhbwiP1PvQWOFsF0csnd7OqgaLnUGfHpUwbeVSJ/ZQLKrLapLc7yMLeAs
F14Y5CWSasy5DFwTa/ovxfzjs2rdAZLgM0auMus0ZdJjaucbB9CneV0iZgb0h8B7
Z5Jn30sWL4U3GoakeG1s56STp/A3BiVy+j/NeGcGfw7vdqK63kwiQZzFIaxrhTM9
+mWxewBjCkHjdxVnYkrhrbRspXBIMZ9zJ88E/yHJuRAGDu2FHSKEPSP2Z3oQPt/u
U18nSM9sM0iPYWyfwceA8rJDEfVjQZp8P3u5anli4NN+trdviDz4i83Z9x/ISZ5N
z/TMSRJ6gXw4YA0DeRQPadnXaqBWtpA+SqMCJEUoLkONggnvSnsDACiChwZ/ZziJ
ggxif62+qlG8D8u6fSyDi/lPqBMvG2QCrgZKnESiLtbgjU3Yb8vxEQ2oPIjn7vuJ
MgXXCr55ForzBOSwSsx4WARhQe56X11hPW5DOdo9puNX1RU/hAqUrUETOuE0oxSQ
pf6Fl7c+uFc0MytuGmj//kjY12Zp1WQQYyevA9s0QwmplOT1RoHKIjkPRckdZ2mJ
qML3sJ6wDPcOP6up3JxPtF1sfydPCwaPw5Tk5eq3WvCXIXtmAIsHYIIcbnvEcyLW
+oyBs1W8aFUaTnLqFhXLlJ3iRtsgqksHw01PTygi1MWPgnY5UaYzyhmQbUWJgywP
zccfHkVC60c0YQAhLZYjrYaAqsOwPV6qbIP3Kcrrss2AwoXyUbHnyw+eRgje3KV7
gYdrUxjCyb5rSQMCz9Y4sHln+FzOkdld5cvDuKc+sRFdCAAf4T2TuTOfH9aimWy9
FD9+HLlLL3/VX3rQYT16LRBS1tTMA1f14pG8G4jSZPSvASwnJ7+qLzsd1ANn2T8o
DWeOk0KB6eR9yQ4vYF63ZKPnoE/Wbt3QVZnQV3I8M5giU0miyrNrr3SzrOO2l2qP
YC0quYwaLk9HgGww0piM6VOJsk5lPFP6AmK4J4j/8PIey/R1hRONaOA5DlR9eMqe
IvgZknoT6xxzHMxhfdjOL4DmYc0OfefkimEeUnLLdpI4zVN+P8G6dxS5PW5cIMLo
u5yZVIHExV9tm3PU+nbbrC/CWfOIbuvIerjVjnGRhbY7Aa2wwFDcccHqNEPigJXU
DI2vxZTzd8nt+b8Eu3qLAG5g2yfe8mZVtus6gwy/WAIx0XeQltnJJryO38hiV4O1
K7bLfzPmML9N7UoEOUrY9cfc+3k89N1WjND86jRJwUD0I+a8sRRO7XRvjY96SSKQ
i98m+YYkslxkfxRS2DHef6niljVTcFpAvIweVpINLtucC+2ZsH0QL0yxMagXhtQE
qggLViYmBY96DpwHJqtuNlV4GuGWGD6zfcMEMUA/DsBik8ZSHJnnClu57uAihIU2
r/ClzrLfP/G3LBl8bwXnLydK1rQl/Sj8Rw3L9hQUb3dMvcbhShTAumZMRAYJ8TNj
m+x8d8aEwbz20PoxZxEEiIPmKrs8gZaVfo8eXzdP5b/FW3Vj/B3cgrhkJWQZQWrI
16R05jzyg3EFdU1eduf6eDOAcHsgZ2R1de/5aZ2w5xuI2mUpwAMjq1nEdnKEAgOl
RcGCpwHw9TgQEPbSzGwqbOxI1s6jR80ee7+s3hfZCO6lRg4jfFX+Nbj1jQ/t4K5G
M4H7+jsF+DwnBqczrklvpVyHfFpOwBizoo/aFg84mC/ewqeldzHKhbUvwFrMgiyo
2/ggIv6HA/OyPLmhPgJA0wqE5Zxgg+TlTK1t5dXEW/XkfM6Lw7bTossNwbuZyNRL
mdKrsZ++44VyLg113F05NszzkOHTF88dbyuTeP+S2H6tfU+s/IKHw4tBatyuZ+zu
AUB1X9Qg5BCvwkiPlEGdGntd0pMexHRRMpbyi666PJxJEJsNcCZ//xVLPn9zO6Zx
9gzCFlc6HonLaR0SKXRI/fv+7GvMBe9jE9nRgGSHkhvgJYewJjz/NZgVVCyePUC7
We2vUss9cVFOc2t2aoNVAyEEDlBVIpYWvtsVBDdwzH1D92DuU10n+qdQX5U1mTsA
qDGNT83EOtD2Ghd3PqVdUmEUt/tYygOXnZWGI8sOvB7L5H3uw64sbDvaVXzUVwg5
A8WOaJdgaGRdiOs0Wd/zDRDmNl1eCt+rytgf7MzQEILzRs4JfWn10dOfbqEubPk1
YeP/RRtW6HCMqsCSeHEitwABqTU4eNxhE8fZAxl1CJA/6zkrtUHf0w4ICoP1fuIS
mwd8bmTK4M4G1cUvcbqe8vPNKA64YuffmlU1uCvDPK6Z/elq0v83oAZL2OwT+RFu
9lyyDzQvF1pmPpEEALy7N1Y1qghhiP/2yH3swwiFf6NfH/6pRPrH4+xFPrhfh84L
rd/oCxVitBmTUDz9q96CEVNU4TbpaQ5Iz+3xZj+OgOmO+3Su8dQW7LdXGr3m76dl
CnnLKBvqyeXOZjdtq8XFEvW0EEVVMIu98pNp0kSwjuucXUxAsfECZ5CBrveolFaY
mHvXaLNO+lem84fDhg5pyFAWuFGgJvEsDa3+nVAiB+5C0XFJhcn0khNJISmJY/5d
1YrvX3zQ2D1iTtuODw8S+U2OoBzfd1yRNWCelUVGWS6rS9VpWl0T22IETbJZ2ccw
bpDz+SEVPg6uE4FCPGKhsNdPvSlvcomLhLV+b0mwvJD3KB39t47faEZVG43vraSQ
guj8pxGsrC63seAivgVB7k/DT6Y/NX20fdvY97JZ3qaEEeDp5dMZHqedfi36UdTr
cGnh1tqGhhzt/RU7V7XKKtG/O5D1zy1wL4avojmTqz4hAT1e84+NYD0qyof1UFNG
szjPgjAmqoI0GwIEZU9JR52f/CpQlAXuE9meMmAkOCG1P78ABPXuzI5+M/VaJwa4
7PIlPIa1D9xV3ITlBN0C6JK5GLYqEDgrEbZB5QFbZCRsC1iPmfaGi4O1yEdiuu7o
5ICOMZfHhXGZWcAYv1uXGIFDGmRAht7Zv9oQnxYS68QOu+J8NUKsjW5tsgIMWhFc
Td3JmXZSLEzxjfyB8Oex0QQOHzBnt1f33WL9j3pUI1/t/XzEJq/0tMYPJMGvFVeD
KQhMu5VRbq56ZjMxKN6/w0L5rgH21ZAIha7rHBAHAvleESQr6bVOMi0ULbXCRcM0
5nywyYNQcVjjBcmI9SXnVYfYA1cfGSha1C/Eiamwx/kOJX0IagapqjGGrSYFClKc
T6aQCQ3PIHPhWKcstWnEZsFdYSNS5rvDr6W5SfugUKSXUSFmW9WLAotE50BHkooy
CLSX4i7MDCZuxc+pyUh9+PYbh+CiNDhWRseurosIFfmR8p7GtoNZMtRRAztEbeyy
fve1TZjDBcjkQHIxG4F8QJn5Wh8Nx2VozGSPg5NwHyKFOXOMe/1BOuinbdlLvtd7
2hTFSFQMdGBUriED0PA76/XA02IZclNGuS9XhObI9chK7wEZprvg5tG567xo+a99
nHHKxspuAZbPhWP7+rldU21SLAL5l2+ooGJh3XWjD/Hb+Vb0G1Kzn2vfOpEzzFj1
qhaUUyh2xJE3sTMZaQ4KGmhkgwaz5/eoJN2vHnhJ7x6JZajPDv86/M391K5fzs5F
5d+2pkssXddkWNHT5PNZUgvnWYDXohFXKCqBLEI8ikNmjsgKLq85RYDDSGHk/mSn
h/JRoKQ1NJJvWkuxrFm1RoEuUAqwO1bd+nnpIDpxEk92bvzfXRrpUn1VhQ9lMqDb
qPAbbXx5xBJEkbfiNhzbfEml7ar23ssVRqiW7rICG92pxJUy1GaRMfpRRh8LsLP3
L+PzmYB4GFWK1tFPVIsyMzN3wpc6yEC6J5QEmmmOpytWKAFCVq5O7f0kjEoWYCHD
qxBan8Rupmr7DDPaVzQHs+9JPKOKt/t+FwvBclo3UaIRgkz1JpvnN16gWFN+Aq4j
V/8V0AL2WPcILIcCwOlrhCOKXRtjx91BIn/QztFu7ZZdJ5fHjidi23LU54yYn2X0
zR6uZhT+noEeIz6MmsSrMAkwkWSRmi/+Da+A0T8NjQBewi3R37uXFCfN2IJ5+jZ7
OEk1ymOYuBGzNBP8dMrymFZA5tdnwhOwddyO/Yn7UrqtUDypiW14IaMAlTix9heA
9nv5BZ1bcm/0sxVK3rldFddUhF2gAdidOspD2J8r90Sl//6j+n/ehLcn40T2wxga
YZNbpUepZjCIDI0VNXIg/id2WYwivifJ3Eb5yb0ipoRDTj3qudQYuZOg5FDjSFck
apu5PJKAXKbdgpWdKbIm9/ktykRo0uzBFpFZXUumL5b7Jz3pdtQUcEa1jkZPhSUR
8lQ+9O3vTEMXv17X+NJS0oQZA87IfaMF4Z9i/xlW5isuQotlGe4TjJj7W+SVuqMK
dOy1zJL/mkS49542cdRFziONkLR65BV1Os6pUySDuwu/zxijQmK+5GBxhuHzRHe9
nib9c1orZjkTKdy0y0J5Aw4m5wLxCpBgM4cezboC+ntcdsJZQqq7Wz5rOdbQNnZ+
KcYH6JB52R0Og2DcSddzCnUYmuF2fsRDSp3n6+rk08AT9cadYSn5Ugh6hTFkfboe
GXQSN/CQHx8/u1P29zNQvt6GJHdb0YkpCW6bCg4GY+rqRiSD19BBg/7nvH5jOIkz
t8/VwEtiwNJqaZCXG5j5kOkIMHNS56Ms3sNIK+tNNsyWxE9eHQfEwn8ivIcgJyQA
SdK4EFddDv2edzuv8Ex2l2DRnpdr/+VDfbbGQ1tE4ZqTiktBU5VzQJF/G95kewhQ
3EigmkgiRhqCc5GDQ74GN+zhsCxfdKFNXvyu2Eo22p/Ih1QlFw7+xfknI2LPdMlP
u2LV/zz5eRx7yjyxX56/W1RPudR/hordrM9dzOXqdxhg3k7XlAvtEDSm9Z6ZYay2
XtqTv3ZeWLAuaAp+ZAvwgb4u5qKTyZrsi3WkOaii77unhxPxfYFojJ4MYbqPTLM/
cx9fc1fntch+pKvDW/mwGY5Jq2lpbMBVPlxr5PawfJqxXLGAEtPHEeNs1AcAUOCP
Jou9U8os5quN8IMGxGnOpcvXPzwLwt2S3eZOEjV3WuIZypcUp8v4bzrfHEkxfeHX
YcogS5sKvN20l+MsKz18dtgDyPpDkYZ1TtnyBSxb0aEQIiDUnJjxw3iV1JcN1KQa
ZSrNLgyHEjJjYUdP+hj3Lh3Qxen5+O24wrOacFrFworKikz6XOApA0KFO2z3jfID
vQiBDJkGmtT7BK/LkzNMN/l6t/jExR7f91OClzANc5wsXUnwaRyia+4d785I9/B/
yK6mJWXIwYba+3q2ZQK5gfj+EL0BJOR0AGIWcW0YYrppk1pbMEuUIhEC07wqbW3N
rrW6WBhX/cG/P+4eaPuUyFL19gMRif7/XMJkcYmFuTtI+FBSkK1nbIy7sOE0mZgL
NWa2s0tPY9GfG8xA6/BcK9yCwze6nSj3uwcFnccuN6F3FDCemewrU+k6dHriU7HK
PpUiFlTOoN4N1ubHQ9brhKQNbGao1yXR6z7CCl8vHpDlpB1qxR37x+PZz8UOvIw8
W+ztWNIkAJwkMDUtQIfi22pWxfm1iZuaqpTEWg4NJwU3qvyx4HAZMqoVtrcM5uR5
zO5U2xpo65fisKanYebV+5mjOOXqKgW6zAjWSAddeSdMS5F9Zw8D3OY6gvZkFSfo
34VsGMWYgrd6E4ij+cZMMmB+Dz3oyeZYQFDAqvldlBOHLWvetTbiG4IGxnyI4KUp
h0v1jeTZrxxewOA18FWux6Mf9hsBJ5wSYZ65FjKAazwpDTZpsx6vstu/NPzeAVNm
guI0Zzfegx85ym0uaIdlYDSnfD1VYnAok4CZ0pieIygDY+UvtvN6fWs+GHFgw8Li
txmqsuAS00BnQglWYg414smEynd1knteeFyzBa4JP1R75MZUu36I1fxI9/2cGEOD
4LhE0Te31NclJ10fUCQiyJ5wDQqJO7B5vJGZNJIC/WYmWg6uGIQ//UgU7EY1y4lr
u01eyi4dGKcftNyb91Tsc+aiSY+mL9LoBj7zNwQ9H4/dxF/TbpAPaM+KVaeIgNeA
ISqlXIeTFzZNfCNwHPdQO/dlOGTGSViM0JEvY/1xpoqBEih01qmQ833XsPuEiOVQ
6rSWlA3yf7kaVJE9MZnsMa2/yQlzDqbOo1+uhZ4I/Eg7YnNTZxPb2iPoG8U0kiux
vgnYkLsR5aWdAk+cM/x9q0TbwxKFt/DInJMWN0mRu4kcqtCGlNW62RH3SpuLBOBB
q9FMI7BxONImYHN/5iW8cXyO9t/+27nps3ZcDiHvctJex/OItE3Ggm8ydQeZlnEv
OU0R0M61bX2MLJIOgP3D3oDZlOdJh6ZOJqk+Dnptb4aWwOztjOimpSQ9pfD1IFaK
qMmavIayajkYYsHCi06V84OztjcltzZiMNzfhYJNSkDBpffHbw9zvNLltMzalZu5
axBq3gAADq+05FsEJChSPSXElPogRbVuZHI0qJb53gik/qoyxu9+F1DDu9DIfMh+
KivFR+cVzVmQC0V3fSUWy86n/O4ewaywNiv9d6UHwBWxTeiS8744br87zcnEHrgF
n6XNR/FWtcurQDnyiB0TCuo7tcPmW6vQx096mfAIOhOciIFgA0qc6I1LzY9jMeV7
FCYRv52dcYUZM4PHBVblts0r384dw3f2WMgZoHO/0vj5TaGTrXN+aQBBJgyYSVRV
rtHhZ23hbXT9ua8OgIsD+/86OyqoFxAkmZOEtCC7fF5JV0aR2fVw6PmN7XY/pUt7
zBO4Jdh2TEKNshBiCuu7QutcGxwpO8tTphYUSCP/wlMLL7aBhbNV0gBdiVX1ViZX
PZzj1Q5c+UN42flkMnm03nOM7W50t2kV9fjOHPAA/zIpdnAWLf646mAJZFwtl30N
obpjtICHzPDE241EeDw5Bk6IKkTXa3sw0KCsdsyi/8oum9w0Q6UZCFQfYALUQgwl
8ojERZcOHjHJg9Xc8ZYOpE2+aSpTHy4uiv03JmunCPwE1ow/9OqAmnm5pdoXwOwI
/LXCOdJsewFzf1vXLyoRRJ266vLB5FVxRoBKV7PLUn/SGxqOlpA5kcXieiDnYGfP
RA+BKeAPgCRNMyrTPjTMZD9vQGYKB9No14Ultaz32siDndbJEBqjLVavKZK7InnO
IuFnGRZ0wrLrKOEgK5cOZh0l/aG3wq+ydYlhDHQBLddS5hhLfMsTLCNmcWed2OOx
xgjWRYzm3BbMQUQBZMRehCHwfYEfYQMOMZ6ZpW1/yujYc67Nn6jb9vq77BRqpw3d
Je7Icj44xkN8fyWuJv+YXo4gKlxYA/qYjmRQmvfX7kZRNAyzp9VJznJVcnfHI3/J
7t1iSd4MPKBkVFNp/U2TlrvI2PpPr1iqArYXt7m461bWCIV+f8mQ0x4dbAc2IJuf
GBSaAS9FSgoNzzgI3SiMJYUgEn7nzJ/OeeJ/a9/oooVbnbANdEPW3Q6vrznI9QS+
47d54oaeIBeXzpbN5EkKGOWq9Ag30IBcYuaGivXiN8uz9X46mkThapBGM7loqGFi
wzv+rAP4cWSL+TM07elPe/7aZdIOUfisHBZj6H/byZridvo1zUHMz/+Pj9igiy0d
kluzp69x4AzOg4C0Mvp1cKe6PAKfo/Ewm8FMd7Qu8VqWxIgsE85ZoGpfofE6IHjQ
HDj+jUkd6bawivYQd38l6adYGGx7YNi0gZjhLeR1AtKvJ2k+WfTxBA/3eCI9KtHs
PDF5h5zQHWBtaXKdXqliGpnJslJ85cml+ZlvUtwmdohCwfAi6UPVz8IMdAQH2g3L
gDyoJl0wGMswDXmY2FSjJI/xPdqh3mg0GxuG0hvPiP6IR0OEpVQyPxF5RuFuaktS
6Ny84oYbMJDnyd3+TRapyW5PdRqS8xEOrlbsTGT5YUf0elgUuy1fG+kwpEyt1j/T
IWdhAZZBMDXIb980Qk3pvTeoADZWoAyJiasILW9bIb7Tv/RIi7S7MjdHH9lljanV
us7KKgfhk7kQAprsuFTaM8W7GFOMNquR2zjpqnL6NVTS4j3JeyMDq/lU0r974h83
XZzNMTj0hed8VsiUEqxgILPUUAWBGin1Gdj/+rL3f21bvyf1cBvxIKHGibTiRbRX
yufPzWaG6Ru6id5VoKejIO4NvCKDKF1G0ZHs6Xu3v+mGBaaB4JemH64CeI460bbd
aV28hsUbBqfhbdCoOc1+ehnu5efe/booUrbIAACsPta0fXoVvcGBWnbWiTwlAVWP
FOYoY+2oFVjLEAauECV0zwAfbjI9MUV4vMSDpYaVzhZhO8Z4iz9pIKcRf3HELIPR
rQZBFaBz7MAnV9BF8MvYzbqnJybUgWjV3uKDsbNXOXpSo+52wpMR6c3M3e5YRjCH
SF0Qu6sJxlKKFiblQp4cFuQ66tYS1ce/NwBjd8cXtP19F6wD5j6AVy7X9sNWgXig
SdnxvRQ7TyY/KgYhlaKvPACMZZDY2vG+QGgUZA9JxrA1yHStgbS5pzesZTqG/Bok
7YRMcJWSwIdyp4u2Ecx9uXZZ8tclBzGtuum7g0GYY9hRRnErwbacrurp1LaXwqN6
Vp36sY9kCIDZZKWOHl3slbjtsrKvpzlu1SB1VvxgUhyWavNKPjso6xdt2dtqSfU2
NnPy6p8uV0jInp36qghuBNpdzYJE2GHFxyJKWc3HZ0wEL6KWYGpvPfd6Oc1juEPp
wR/ABCE22KCnVB8CkqpTTl30biQjgqkhpJoMxqZlr0afA/ZIHI3eB8Je1w+gsoaa
/qmZLsyPmlQJUdHHyGFFZ0KHG5ON+FSsgkTsmE7Lad7tKTGIMgJT4+ACBbsf8Tt9
6atOTv7mBXt1CnuzuqvL9p+DjUgw5WMojrtDhPrHjxDBIG0fj7KpUVdGSEtz6P4q
Mg2VRkquuAxqPUaYuyWpVavFyhx3pCfdGeK+yZUTrw6Qg+X0J3R4eFBqUpb3F9j8
2uXjyTNTmmEmEPdwYJ86+kijQmIS15fpOFBUna+LLWik27oxW/sflYVPRrgOxiKv
WnNRCnafYWc03W7P3ObwU/o3K6a6IrKJZAI5GPClJqlKYDIhXHe4oJ6Bhd77f30w
wSI3xbyLJXaPoXOXW2pFOr8vJyp1LKrII0MzPB/jynee5SXSoQFrF+bmcK+j8+3I
2Te7y98/QyEh9F4DOHP3yPyY/AP8dlAzECC4Z/GNC7fOvrHKmRBo+c7iUbQPfic+
bPySr4UERahSalYRMLRsXV31RW4QUUqkKHnJrZkgW/nHsMpf1cykyach5fwkbK/A
xwXxZRXR/61aRyjoV9zM/Ci73IhrLv1gPQZsMIeFtRIPOB4TgHzltPjKCgx6qVwO
L1eWE4pU8GLLkExyeZDrRLeteeiZb8zMZJ8SUDMPWTZjn2ffPX6xlJgOtiNYOmgY
lws5z+/57qFU3w8oQBhbgWkvlNLdKgHQBni+QnCSQNr3tQW0sH9GJy1UEKD+xBh0
WiON/uhNYX8nSZ5rBKhdlxG1fVVAYJyf9QVHuWsTsKmLsoUqCTW+KuzW+xYoHunU
Xp+pcwhR81OZSXcSWsuRCbYi48saGgePZlcND6XkvyTl0VFquFALKsccwE9qmhoz
Vt4sO186uqbe9U9bBG+vR1r40iyEC1K/QUMUNUxfOxxmLFzQYxak3uAxU3dRgJMB
8CwFf6CkEAiZxOX3JYf1ECsYZYI/Ogihza5uOGvuOIUbstuIAW3vYecNCfEgAw5q
oiEooFNgvMhzNI1GNi4roSFcWZHMi66+SpLddnjbK5afDb7Clc8QwyRbYe3QyO0R
S1VtwVDluUAWzVppsyJ+gJhW31nomHSfTGKDhsP5oLhxECIdKd9hLzeeaGO9YWa2
ajZgjNqO6bCCPtznxZKUokyDiwckQiO0UaTqD0mBpaIkKWluSjtlVcTMJIoj9de5
EfPlK7I8RWN9DLaC60vFZUh9IiZ2fyKyaIpbzOJ8z1fT2Ys/kDtS0jDthJ1cNT6e
0oIY0evpmR2K8NnW1ktSQ44LO9MxaE6VtzPAdeR9pfFg/EPX83ZD97q93bzKxAeg
Hh6zrJ2b8hvpL0nDhlUYM8gbEa+cATnYVk40tYMy8oJzh3JKHGy7bHColh6WkVjZ
TbEpnfuX+Mai6vWdAauKkrxQ3HMLOWa4xSXFF5AJiA8WrIueOfIkEwPwhaapw4vz
JCNQW+12vD5KTRYVTH/qn5EOQMeWiOxz1Dkl/EhdYV4m1F+HDerRh/IbAnc/CAI0
jL2lW8KEEFzxJ5vcBxTjP6VOepDoginVwrI2tYd4ZjQ7wkIqZIkSoTwIHzAs9ObW
kBKBdIysnTTAXKYGD0u08s5DI8m9GTjJPQ7q56Qnm0DSixsvHALdXO/Kimz1EzbJ
S6S5hBngNDc3oLoiB2lFCQTjvB+2oCJe1I9uRshyrz9EmPEejofynpLiSrYQIbHq
nYoqJNKvZKVKJWT5Q3acH4TJotehDlbqq4lPY48L/T93jTMqN2JVce9Br2TVI5lU
DGbCyYmjCDWoELPtcF94lgBvnA6q0ib+gQMBBCmp0q7TleU4tAMVeuUDWYRKOvmZ
oST/eYLaQklwb18Le4UUdp+sh+dEsSF4Mp+yJ0ZsVozVY46jood/0uGf7PUktxHH
aavy6gEPognoT60oDSFfI4Hyfl8QUqzDvjUITbN6IJd2UZm7T13Ru126+KdUmASn
T3ZND2bLzNfyoIJanUro0Bde25+rcnESDod8fxcxFG6G3kTizZf5n68euLc2Btkz
az1X3xyzKLL/LRBtvwZ5gnXuaAoDWcMiEoaq8xTAMQFVQvC26xAPtxADZD2YzkmS
mPCLxEIyPqJmQC/wKwDg7BwUQGufm5XElZSsz0lZvgfxYMG2bW5T9zVE7yzQdk9C
vLTkyF19jf05UruEaj77B8S/MR7UOvZPDDBol6+lDjLiJZE/ha01TMjo6+ePt9WK
BM4qCVdqJlbZuIFS2V8DYzRybRvmmm1wK+n0pywpkoWJ1/u4b1tn6iYNUSHSHitI
TYoIxEwwqCP+JmldAuR1/qdjqp5DWAotijfb18+cijgft/OU2D7qePIlX3OxLrAY
WkNOLXhoxZRkvucnzpYnQS5RaJ1rGdD7X96bpl6rx5c2KLo4HbvVvAYgc4gU5kZC
/Nw0nsCn8ugUe2AkVIQP4apKKEoxgqLkBLqAH4DcBHLaaXcDwbITsKLNYGhGofWW
b+IpEJlOJGN2vq+a2Aqw3XAcT4Cb2rVUsw0HEEGawJZD9tz8X2cXVrThhk4vZAnG
/bpXXbS2rXEqd6U6xfZJ1nV/FYgWDNs+biWOhsWjzQn9Ly7Rg89CVLgZErm26n21
SwYeRKSHTrIzXy0JgisXmtvPpgGoIsGbPthYw6cXuVt8dQkxkQeRgQ+07cP4/iHU
zRgJbhcY9icBejjwT03Vwg6miv76v5sZADS7YkrpVb1uIrAzDQ2HMPPeUrHK9GrM
+m9BwCNuPVyVnu3hRs9ELK/RHuF+ug+/ULKoOov7+ugHparvogbSRRNsbVXySHtL
V+fbrk8EMaatGkntHZ9WQQthf9/49tyltr05kf5sfcz/YqeLTadCCyCF7HuN8vRM
HwtUh2JQpgCail9HR39MlcT2zFTUH/A+tiHXM/l6SLYMX9+oyUfX96CIdUjyrHw9
Z8E0Yc3OZJvikrRTltoqvasL8GyKEtEsvHl0tWdEHorMWoxvqwqsmmgrAq5tx7kL
5AsvU0IocHaa3ssFydkwE46srxjjTVEEP0JB0k426Pk79XRnrtjm+zBbGFjZ7TF8
tslKLp5vVNde+tfbcl0njco4X2tYTnfw1smadh7GM0bhJwt+GikadOThZ5Zbz2H+
NvWJosmQFZF/G8oefxbCd/y4N8YuyLYcwDQ9RZwX/B3QlJVk0svcb9+imugABWtU
0ttQE5OiZ5uUelfI8v3chsvDZsP/2LnaO6ZBOrWDYXBSUzYEMcp204csCK5ZjXuR
mXE4taf6ufSHg5Emz7NN81ToSCs4T78cj0bdpSLmm7Tl6k9KJr59nUVbXdW8fsqI
8N3WA4En7NfjwFWhZxHe8p2qTLwVbVz0iEntwj9mCbpDubOvExVVomq90r2zcVV6
00gDN5H8yCf88nYmkl+1+M4r9aFW5b3rugvBS5YzwzKjic5FGZwFkQMXmi1H3cT4
Wj3841CZv+tAj6umrg/HUtjtiI0JDwyp1D3GecspctefdHIHTDfTFwnuvZY+Dc/A
9iFHIljgI3t/nKRZUZbYo3TpKqXkV0pY/SmZNP/3fst1gtT8E4J/x3IjudyAWuVl
eS8URW+IOTyHoaomwyQ5C7mk68P+cp3bIuXbv4kq9DzSjWlMGo4DFtC4cDMR8u5V
1tOmhHVhHFLnFR/3Ok5nw0R/oXTDU/jSbYZ4e1meUaduQzRnIZW21x2H1srMMxZy
s1G6f+HQtA9FuAjUI3GDx/sYn+gpY/qd6rYRb/RpfVlinc9vVUmq0/6HPnBNh3Fs
VsOyqdQxeRUJoRCoRbMPnpWiYuggWHgFW7s3qIA90tHjBJ1RWYyP5E30GfLWW8ac
1Y7o8zbkbIDrN2YBLcfPTL84Sp3e44Rmn21H7rRXTDCdeKQzrhO5GEgNQqHoPY/b
pja4Y7bcwsgnbn4luT2zfQHNHXo6eKwtLFdXDpJYIkS1sXjrraEwx4pjxtq/LkXB
QI0BwAXNO3oiha/8M5DL2EAYFmdUAebg/731Mtm1Y6uehk2d9UP5U2jRsmWY57W0
X+MalXQW8Cf1KR0P7Eg22QiwjvUcS/21mrCaZpXuJdjYp2n9Fvys8vZTt6Ijj8qM
95Ji4slcRSCdyL6IdjZpW2lCyIQB1zEc3beDkHof6WIvGgN8bNKj44PMfqLjMSNP
gJrKaWYOXrMxFL+01ZH8mtYaNCyMYvJTJ+1KTj9zE2BO/cMN29YBypp+ixRgnHaf
GJ/hau2UXsSk/QXQ/pWJAY1WO7vsJHass5YDbacshrZ3Ch3hLgbzH1cbAViqN7bP
4aChT8OE2meiuG0h0T7j28u/1pSaLWjj2JTgPhAbwRHjppt+aXCDTxf9CNWA7zay
NJPa6pGf1wQO8h7ivOYobegfmvBM+CWxGyZScFOtYKDa/aLdxsQS8jc29NDfLTXV
PFFYXErtZ5eY9y6O2ZSHnvaMTaAfugrb1fTsBYUr8T34gyOH83OE2IAT9CIUfe+a
BXA/VmdnvCMBS4WkW8un3UFBnEBhM3ATmcjtTkhBKASmiGJJo/+GDAFvykplg/HT
X07qguut0NsPwHEL8GQ5xUAtLh2RsKpxD5JJmWLPt4+/kuApoR+drDdigLcijg2z
Rrc7UHfCzhh78bwNk919AjOjLCT23AiFjKEr8VAgDHnAiVwJpTnHhWI/OHwX5HAc
QhkoCIlP6RiU64PSc+K9tWS2KHwbilsTE7435wagieoD2piU6hEP2XVPItQm89ur
iMxgAWSp1DGvoLg1Yu7m9+QmecXGt+IdX45pU/DYZwRGTuj0kp8pf/MziU8zxlmO
Xy0xmgl/b99bRnxTND2Tv34gRRwN0OtxsJxvLwCZ4FsbJnUsIFIXOdUn05CJmDhd
vhK1eTuip07IoAlptlCIkicLAwO8/eDnJJkeK9Yzf548658xMIRKt4UbWsFApha3
ecpO6KJgdMugfwJtD44glcSx0KffeuRcf3//X6K18G17moXZXNOuds5qp48oiN1I
WNplNqnPBQ5lD+lucgwn7PYGfHIGeJ6e++FoxtsFHtGgqZ/lhIqmrjjtxGQIIfEa
Pe29PEOxi+7RKO/vZ5JLMK8iDjXKBZUl3b2op5qsUqFfWRAamwqkmKWiS6Ndmu/K
rEwaMePVjUa1b3mpRz0TzGGDRkl/yFmP46wkOTH1A6lsDLul8p9uxWiEf489JlWd
IL2xRZS8oTs79I11zhKy5hbVLh+cuYtVmfTHU/3a9CmxfBKqFvHihW5t/7j7ZEbD
d5ecXWKbtjX8oaFX2ucmLgkVAA4IRxoDS0VueDfm7OKkEhJuhFYWbGH1xwYEvkO8
ng6r83mX9PeEope9PKTaXMs7+5buoxzeTlhpSK/Y4UCV2HuURKtDfhOCUojcXLea
uRoXGKNyf8zEOHhvbq4vFmRWEzrSUUpd1rP9ghrGVKpPRXLp28n+4kq80ONQjG4D
Wie7ye/ggGJT5vdpehraxzq5mPUQd4KTHuG2k3zlHPMcQ1DJhDA3ofJOY8g6XBfI
ihfQfdEZqwBU4TbV0ovvtou04+XFZpKskeMyELDTUWs4ISyVZt0r6GRBiTw2awK+
KQM+dWudIkbZq140rtXl7rXFf6N4Y6vHy9ghpwisBavjhToW8Slr30cWXlnoKXb0
/07nwWD/EYLpv8fV/T38owG9AclGgT1ZxgmpnuE2fQAp4X8ARFjbX8EyDwC84Iip
HgKMYITmRtsEF8sbhQiraZr654GE/oXtJCTGqlkw2NvXLA8xchNvav/eLtFcEGkG
EeKZpiy3mdYighv2GEM4iuJR9/T+XXWeZ0/JQaLkQ5l9BHO0BaVX7j5hWFH2sRQE
yTMPytmIPQBSKre8UP+DoaBQ8PWP4Jq3Tl70po+Gw42uXa/XsfdRJHWn+Yw11ilY
fg3lHRorGCDkgJGnyu8h0x4w1oN6PlrOkRETa5NnzkZwBAUg60dmfU67yVt/dMHF
HIEIjz8eFGyy0/h2iL+2XS/GzODl43WdhzrNLVXz3mMv6qw42W8u3qMofyX4Cb3V
bEXaDLrkR+9MsN+wxyGnEzMq/1Kzzd5vpOyVOvk5pHOa5BKzeCoekVnzRrRb1SDu
C5JxR2ktkKIlHhuL5tgIlFFGS/4elN+2oBDxB0Ebq9xL1yqQovb6dM/pYhS9KhH2
8dW/tD7nZeg1d/HtsIBwg54MbMzfYy4kAokGvDuBMqfbZaWz6AVlK7NDfpfvD+aH
j9TT3ARtbZwP3SL+HiYJ+iO2nESMKNwGr4bCi/hntPRIMxlQmgavct5UKjY61tAY
mRnE1U3G2Zmr+Ym7lnM5dHwbsJ99cR9/oCLHGsOlQlrY2cxdtStbzQ/3ky6SpF6q
c3n49QO74IqIRLCK0W+mu2dBmJQ6q/4A3WPiZu+01vsjbqs57kxgLjJIKCxfHXcf
l7FpKv1f80BdtCPI0tuzomC/mI26T2dcB/yO8sdSTMnzQApKUnrocaycKFrhQx3t
0urIXC5c0iiyazxdf++L4EXdM5J7MNdno7Cd98U5L1AAVBJ0paYjZjrpt8TAnuDV
TEq5qwqMd4W9fnPfyZYyg3vnxPbEKschK1t8LzoDGEctpCX/bb/m4nZi8iG8rQ71
XwLGA81YFUMwtikUY3BEqw1OhEDkYuicDjfxCB4yCKcmCANH4nxz+SHgY3l06KFi
IWxytw6u3/PHyKhhF7D4OUdlK4KPiy4dR7w2hEvPleFhfd5p9LgzssQhT67sBTFn
KcnEIq/Q+VciYPpIQbqkXf1P1djzvRPmJXtMtuKnEbJUlz8E7lvXFfLfnf+dLyK+
OuHOPfXCoZ/Wc5r5DenBTu37nwB0V8f8EaXGveSKQ5KVrpWM4d8X0qUIY6gcIXZL
+weVxoG7OICAZNZHq0DRhq63XQCjIpIrEdTYY4cemmvhTezTI1+pjVYlQ4IyqeFQ
vi4z4Rk4QFjEEbh5CF+eon5G+mvdY0VDNDZJlDeiErIbE57iklGIujbznY6+F5Kb
QtK4DqZ/W1TeXfDC4JFkprOnWaUzMGFsctaS8kGJhIq5McJMmp/kQC8Tvjh/cMeE
4B1LAjkG3F+See2fRmEt+fuFzkLoloHAWDq+SjX36Ud660QbfzJYjmTd4IL68AyH
zlI3kciENiRxEN64nqXJwO2jfNv6UJYEG3uFxE/yYVJnywDx1pAaSQcZnx2Cal4O
cacmWztPcKQGg3z28IgoisQA65+byFJzwbdR5WgtaGinebO8RqeDxK0veVOdRBKR
0dSICNqK2/ez0Wrpi+Et/tHbNL1ZI2fskdTN30xQmopWWoHsNHkF3aNFZcZVU+0L
w1L21KU6WAP2frqbAu8MNITJ8dUZFsrFIqWRCynPSvRONVC31nJIkDXbhV2sxHCQ
7rgxyZ2k/hywjM5eNYaqbREsWKTRHELsxDKyV1FopOUqP+DsU5OpdGKJ52x45cvH
WPtUoSUh58UycO/f/a1qGpCK7MR+DS8QRVZzm6Y3vZGr5zsA2VjzTYXQ1k73El71
DwkvyF4fjwZVdxK5dNyAHId0Ql8NJ4k5gMNPj66pTuVYuLQMO+2ca+VJs7krxY5p
+0cwBBlo6Ca9PM36mK69ha4tsDS2gMNdJuhC+WwR1ZJDC7AFrSumobe4ZAD2hn6A
1Kgm65Qwf93DfNWk1Z90ZSjAa1BAQCCQ8W/dEGwyGfi1z1cRMDzmuEh7tWlGSNa7
huNoslb/IuKZ3y1XeYPWI1f95e7gfSZmQXQkMnhKQfnPSnlTqS9XyRf4Ca1zwPaR
RlJKHElE0aZAMGFHM1KbXg7zObrAZwnMi9EpLHOcN1HLOG1PvOwswgFt1FtbW3Uu
rPdhAxHwMDRk9Y5RQy/N+5jHI0aMQdU9BKPGNa1gJDxLnOSWRulooMq+okdqRwcv
xyTBjjIk70HkSvThzfAqLCaKD0DiuLIZFeFHF/jmqnGCNnG6rsdXK5iOtGx6xZUC
BerA7H5nl42wG2IwHFuCl2iIXP9O0WfWI3FGR/A027DLHZrouZ6gwifL3FmEoo2Z
9k4dv3+IbkFE9GFCvRxp7eSrEX3WRpKBIvaSU2Z0/TLw2VehbK2QBOgMLYp/2Qp2
SiZgbMfF0wchLrGY5XD+eKkmIkE5CkhO09cY3a3b16Q8D2vq+GUck6rZR4wyYsLs
uFjcsYAY3GwbkX5Fw0a/N84nyF5I2soqzSN9sLbzxokWKC82VLCmQaqRtnlmoL+k
0Yaqcy2bw9pe2QhOkjosB5WwHOy/gJuuWb9yvcMb9Utp6AXA7W3g//pOIGVYpcpJ
g2lEtOFoKH/qEmaKhHk+zWzbsK5Z11PVYJ1YkHdaVIPtCfjofZZEG6CzE/b5GSJ2
nD0Han0Eeo+IC9QOrVUAVhFCLYcIDbsfWCBjzMxwmAINc9qdfod/X6yAUmY/Wqiu
r2URqP6xfeHqIUOixmMGlRYuTT1spNEcWHv84m7AwyC/Heqrp4n1iiO/bi30kcMz
Oz0kzBFc3Hy69j/YsPi9pGioXQImlxQHqAkhGX66C+fA4hvpWHKcreSTa+6p/yzj
e0zRTK0CtMCfZPYq+hTpHV/1t4kRWwv2jbUDKvrOOMArrQTOOa9DhwmY23SDe3RR
6bn/SVcj1exG7bNZNJBjS+QJePlZT0EwNYSgHqpRyPvhgiJKZZsRZJz5TIlF6UYw
5QbwY3FLCJpn8h8g5+/eWlLaotvq1UYwC9ysww1dzgsKDdnlLBlJEreR340SORkq
vRrTPLygnVZV+SbgFklC3zee49O7jZYCCdzJaCBWFzSAaeP6kbyli9nPsiXkrqPJ
u5GZ0tvcSlCU5JfDykYSJQwSUTdRG8HUM43NejSGcIauaoON6pQ55yVWZ2u0n5XO
8CzfAGb8nwsAeqyaFZlwTfzsl/5Fw2XbOOY42gMK2rOSrLiW4uGX+YsMGrDSiede
VYU4nMPNHBC39nZLHMlBM+V01evT28chFaQhj7E4tPuNSReWfsB6RB0lioaoIi2V
YEkXx7GFsvfw4+e+1simyOvGg7t3XdcQ+MmZVLdCM2qH7oG0gDu3GIOt0zeuvNAL
qeM3QuFTBK9imQ4tllA9kuwKuVGOUS9DK6bxOEMGL12mKu+p48sTAldZxWM/+FLp
5DU5VZG1dNbHNkWaDhBZrZO6hoNUGw94tCy15TEdBu8bS6bHQo6QjIgMzVod/7UV
1BlIHrrnf4raRxBUe/pKMGd93IcJdmi0qH8dI6zBaierl7hVqoXNe6RqblnllOec
sHChIyg36VsOZnUmezwk+PtNfb4b2KSvMA+GMp9Q/olrmUo4nj9ATNhsQQ5S/Ile
rlAWHg1xWzHt2siqO2nYxjOzwyzLGa5fBbrvhNxgM0jSWQDutqIDVSdu4IBpREy7
bNgwOfBGeKFYY+FSW/eHjfZYCyyRsGLCQU+i+blaYVSs3J0Llp9bag5wZ9kuEiDO
crT+r2dtwKOiIwv3mjSfaFJwdhlVNvUQ6xCzv2eO3W6lneHWJ3pa1fZWCOKWrgYQ
C5G577JqV1xNKjE3QwRjteTd9qryO6VrQpzlTVexuBUH6JhG7NlDiDp6NmwLiJ5j
jnd3MHGc1shPfWsYCgXvuh80X8prK5Mf6hxlp1rkZI1BeVMAIWT0fDeTOdkMkjFQ
wQnaJ4J+OWi5rsoz6/CZGu3o8XZit3pBjKxgBAfXF64Yj9yE13bEGKTdBMyqkVMI
ITTZJR/sp05PzOjWRbmPVPFHcNNhArvlIFovPbNtClzlqVARRyNduovcoCfCxc8f
qwtzMU1Cf0RCDE42WuHWl3CJO9Ad62oP5ek1j4HLw4Mwpp7FHl3FVW5wboRVQ2TB
7ALfdHeGvyByyHrPbaPzUYoAuVIy42/fr/qB3pTIzSpgszfUq33xH+u3hc9jI/9p
Urqo+O1GYawSBMtBZePmGJocsyRrYlBo4YNwK7C6lmm1ClzFHWKQbLglPW3fQ/0o
mM8RiTpCIwWy0BIhtTsqfTlbPPD+08qVYLjCmXjn0s33xoKDkZFRSNWxltnwt7ae
PJbjZBoxCcRqFnosE96mcjjus3NQs/JfnEJIJ0/Tx7QKbdLBNHncCiJajwcswuug
LwZ+GcXL9wXIJnMT3Qx7BmaH3AQ7t/9IaeSWRiFSfbCMY+h7uk+/HmRkPDndT3wy
Y3s3RJuATWB0reD5S8sxwxjSV7ktorZ5UXAxUOoIDHM7MVVvXSpWBpWlR1gjz5Tn
kXlsYx/OqW8ryVFy3cPZpst5swSn4eaXfNEA5UIS3+ltUkR6QXVsI0xVqC7NXflu
JHsG7taybHSBranXlBijd8pILnhwTCOO+SBScCny0eZWyo6Q8ms20T6qWOHkvHDJ
/KcnNt6znb9ClfgJFGQRsf4IYA9rx29J3Zr8ikc9nqX8qDFiIjHj8aHsR0C9IJkB
jqbrrONQNlnSrtoVPfzuTBU1pxJT3FgLIKfxYQbRMURgcuzCiz3xOXZhPShNewgY
sa3acyLLEpUxt9Daqouvb8VaE704os/bpJwB3KJ3nnY5+9974AcXI0kCaDfqz+3v
2g5xZc4FDrjxNXZ2sW+yC6xhqoaLmV9/sS1K68RR69apDcJYWklZhoKHXueaP8Fm
x8Qt0iwA34fTVr8P/sDygJ43Q60BrgNfBOHTsL6r3PXxcpf12MJ+UsFg3pgLkR3O
hc011MTLuVyeAPkjhP8K/mB73ec6C75kEYgCAHrOdw2jU8/CYWRaWwvu16uOl9Hd
DCYUVn5LlHbC7twymdmpwe/jZl+bt5gxCk2qAt3EkEFXTzbBO5xg4szttn/292tS
wCEn92Pa6ShfMP9gWrFVRHSI0qtaNKBZ9NKlX+vltCPPbPfMJ/voPPjmcPyh71p6
Jzpp3bKFuCUKJWGF7b0XEqY9A3336i17t5UIhuJPUibj7yI8fInPAfw7qg+EvnxH
hwJ9tgfWXl2bYB7vT5ykSsPbtJNfCSE3gX29XfvH8ymybmx0/aGnA42nNMseTj6/
6Xfw3L8kNRTwwLqLg97NB4WPTfLrrNYm22nKIgyba7DgEcOqbIwJzUhvQ/sQ+rhY
OOBc+2z4zk+mcHDy6b20Hu0WJQGelP4quA3d2PXZfUy3Qci3/41tlwFp/XKRB2A0
OyTl7cPp037mubGPwYEztn7XBvDtQqi+YdD3nf4A/T/ld1wuTG4ZONoNt8ADs9rk
VDantOcJyTH+zj6nPp2mkMM5upRIy9TmJNGp23uTpo/nCPPWzFZj3Q5PjRY+9Bm7
fHf5ORof/f1rmfMFQyEjipFDoPKRnBioqMWnG2Ukizk1BCdw1a9+OYj2soxkd2Rd
wCui8RcB/LVEzcvyRPOrCyEOfCtxayKJrMDa/Onea8t8xd+qVLGKN6Bp6CkSCIcM
rY9EAqDirNOYhpqOckDCAG6udsdNEev8N4i1QOQ+mxt+J2p9oRfabosGMKFY20BU
nA7zOMXp1ypITIrhKr60ONwtZqyRiV88+BNgXJ4XHmGnI2VTQVB9Q7+3USAHbN1r
ZiUHBG2FkDYLY4aKHqT3m5CUvWmzR3+zs8bYluWxUpbocz+JIZcJZIk2e+lR30pE
OdULzBRSIkmX5DX240t/9LjWVqd4QDgihzRdOAk+2JdFkuZndEs7EHR3rjNZNztB
G24Cjxf1AKHJlu0HD+Zn5+YoJLW1jtgQ5731ACSRB+tkOKkcZOBbDZmPa50LTmWN
FVaKf88rPF/y+P/5v/mUEHuF7lWd0Igk8apbTVEJpC1bLbSavK7kfe4e7L+HDJ4a
AXYwQEPhruiO6QXEFB0kcxvoE7x41uFL+b5esLpINBOq4elUCJg9OGiZMW49du4S
gW2sMXieH5SNTbD0ssGhnIvjik+ywpZVEFVQClsOysgsPaqO2DRhNou5J8SAY8nV
AMwosiX9SLVyfgwbu1c+ShM9T+cW2pmNGfGiWfsT/xAbEM+PKQJr3K6IJLZ0Zvxf
HpjZMnxliW1+GEAnYXqffU8Sw8DwFvRsvbQ+42rPsqJ6A6fOSn+fkPHBaRd/2275
pUr/cCencuFshkCygFx27NIHUowUz2dI3Z2090F4ZJH573HhHDN7jy+ak53Dx/lH
yEnsX/Ej5Fsx3eWtQ3vFJg==
`pragma protect end_protected
