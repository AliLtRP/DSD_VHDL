// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
AWferLalEKxJ1j+wfnynBSo+17yuJh90jWw2MGyji34ezu1LIjswma/IFe0u+g4C8EmlcWP4UOGC
+xN6255SJ+BO29ILvu8dqspeN1esLIpTHLHuTBRyUSLqFbPONgF72JqhWtSjWtKj9MGFp2Nu4k9L
To7cLbvxdovWhM8RBToo5gmmO59w0BUi2FhLEZ37YZKYVffKB9bq8lupG+H3gBARFwMtWbNh/b7m
YRt7Fr18nsCWi9C0q41URhauOdVcCIg60aM415kaSShxRq+7x44fjA5t+0AKSqKnyMLU4mOoYK0q
T050kEvpaKtHuJbOe+qBQjlwjIS/TxWCDVJwiQ==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
IwHHc+FGJtdoyy11OXkUPoSDmvlFLCmM5nv9HBzkuHMIJeGwvTubN6UAUaQ+I6cNklVUeMysXDqB
Y/YD07qIpzPpfw0RAiaA5jcK+qJ/iCJgd/3ggLU0qq5yc0+hQja9bPs5uHRV2eoJ1jDzPSA1ymhK
5YCZVDaJZ32t8UJ94kyxIcgdTO1K97duEtiS4zcRXspkMjfWiZAYgolVtrSqMVDfV6hPPnZH+IeA
kC3Hukg6+wogwoqlPLZqhgtiIfIq812cseFN+MQRV89fM5J/mCbxQ0ZGVEeVucA55adJokQ7bMvw
d6VbN01M2ga/eKOWGRYbTV440pNXIexIF7/yCxxYXiDS2pU5zg74VQZ7v5O6LozZDKUk16qpGGlb
EbaG2u4o8LtArEjrGTm7Jph4nUa4lyRe5ppCxmykM+cK3Lct/YYxgYkx5lnrqA6Cx6TDooFe5oka
JniubfLQ53MhPeEWcDV/2nCZlmEcsr8ZtzC6KrnWzAm2luIVjLdeQ0RHecSBJj0hB4r8yqyTu/HV
+NtMfW3lMcrl//KxMM0JaTMibrWeMdGw/v3t2GUHDSFaOIc7nsnXHGRmxoIhctOVwUH7tqS/3xzg
905hqeaE/qaVNQqlAIBadtRSvy1mJuAe3mCTQ8gEhBgOnmE3B1zb9xgA70nm+1M5ajDZpM2PY/ip
TWBv+N/7QUzRFvfZha2lhx7sHF/n5R+cVONgznHKyp5FoA6cRqwbtdedVVSqUIuJngdxw18aTpFS
IPdJzwzmzIQC9C59OG6ZYatf0Oq4bNrMHGtTdChK4rcugrdkEaHWUONKzDGGKGsvnfrCb14gI5hd
uLOoe2vG/BMqQH4znPwpj+M9BGt0UBq+9c1sBHlSQk5HfYo7Ti2KnOtvRVWY06K0c/3y949aRNqL
0w1UnywenZEJBMIH9ySps64gdBW1A5HqGUA9aqq7Yc+sf2RKw2BBr3OnGwLgKHOMjRmazBTPIC6z
9xgGle6HcKekBNVGjDP7kZtyCnsTsExp+oGmQKoS+hPQNVOO/VDemsKJvq1dbVi36Q4yZqzo1dg3
IMWfux1udyB9HwoRqTpL1s1MX91qNuAs8eWfjsFYR9dl3+H1BQjsdshk07x2gZpl1WXELlRhLoS0
9J+oly2ZuxPx+Tisp1QH4mOmpxCAFugFr/yQgbId72zyPsRBsT365nzZM9j3d1wtoTFH295/hoSW
+2OrgTXq+TG5cjr1LusMw+vtZc1lpXsP43omG3brryuePQVZ7g8QfXaRH0aB4CXNiNOltflBAFvh
64jTroGifDG2/hGgJ2V68BhtNFiUjASZKpIrZX5f3zbK5sV8+Hs13gbXqX7t5+J5o6WmsVYNmhMm
wHRAF1AP5eBgxvDptwa8AENcSsfJmmahhl8LuB7+5+nyokDeZ3xjxbbqfGxGVo99Mv3zaTLnHR3r
NsUb3812H3veXqbsuPFikdSR0wDDES9zeICI6pG+QyGpoBHlKpDHXI2N7943i3FaVw7jgyBY+cIW
/qKdriPf6JlHEziHNfC1FjYHHGTxdODMkEK0QmNMi7QOdHaxiAAWc+gV/W/SsSBqbgFDVRSA9yao
Juxn8R1PzcPk/FnIxsVodhMgSirIldKhntiS+UCmJbS6dcNAS1epxiukiJvG313rzU2UGglEyFFk
XKclXtcAgwxM6upNxy8hemonN/n90jKZQnWvwIvZlCIJWh4vRO5z1GGCJW6/2skZRI547+r7h9y2
vZGM7C7i81eTYWhzQfYlPcRjAv+1tVhOS79DKgKK1FtsJxcOPJxLM951kov2ApnWEJhgM2BxrzL2
m+f5nLFDhQqpCTvMtTiy5AQ3RqeI5xzXabInQ7/7yxeOcxUZX1xsM+F8VMsL2PR7rz59sFRd9pZm
Wy7gtpdDH8MY5o8fKnVfT2WmbdYMoUzqCjvGAhjqF/RhKzIY64cnUD/PTL5ym0UJV8UgLFT2AIuc
bSJsfM0e7Fscjo0ckQ8kiBbBPIizSKBHtGiQXnoV8H4vVCcyyGvWiZ84fnHlntVaMJI04vJ5xkPr
LnDIYTYH90aLOCL8655NOuLfBHLu0K9B9ezA6zSC+ZDBoR6Lu1C0Y3OKnASVj6oU4EQ8m21K696c
Vh+rmaVuQ2pRfj8irlY5RsI1F6rf2l9HRgPDfhNZH7aaqTNQJ1POqPsAvVjCQIJItJq8U7UDXyI6
U8i1oifUJqTfGMxFBz1wLp/+u2xiyzpkN0E53y/IlKdwUtJKjefFwbfgjBJ3G2njizNEpxBmIKEX
uTkJfFblmE9INl8EpR4zyGII1+Ag3c3/Lan1L8I7YnZNvDlQO1lKx4cmuZdc8a5l8gXzQcRTgvry
J4Xn3eX3iiBTXZ8h+AA+f4HNEsFxC3j2EibAVLG865UbjiEUREfJOjP0GTN2pmHeow15Cyw6Mh0C
bUbFCEIGOG5xN6sBh2isGRmCMjEvyor6Y1xON6CCzIxJBDy1qQa0QyJZoy37GQiSalROdWD6Bq/8
QXrWrw+pwTBHvIzcEX2dks9rbq2qM//wGSnBOTeozfD/qytnChw08codu/tM6Gdt8cj+OyCZKofY
OdjUC58nSBoxIz6NULyGCuuBwvmWmFgk4AyV2jV1M/X60cj3kPorzcQADG7agTsc25LmqgwayHcU
YdULXB0T8dOs7QyHpW4jFu+GwbAsMWwQN+fJR1SnEDMRLYe0DLHSDV3+Ierp+dKiSkt9RgqCH3+W
2f8b+mWN666AeJ2+EyIjnsHrRHAY8EB+iUbJTZxE+bCazpAR0adY1RDwm5a9sUtqsDFrnewR7A3E
5NVlDSNq6FZMglZKN3d0Ly0KXyrYlRj85tYgPvEWr9sTas9WBQMD4qRYBCAmrGUsogmucYHNgr4x
McyiG/34jc/EJss6LLdj4kCTE+6ulZubHQwOOaLBY8v//lQkPLNGHi6/hYMIWS3J29THyGDv8uhw
B4aybFKMYSFBgxA81P2st2QYmyCZSDbyUCOdC1kKALZXf9rSpd/UWsSkSf5RZXl2w36s94kcMDya
eVzB17CJC/UXzmb0c3Z2b5J08+nrBP3AtLUgQT6UdBzxlmozjm4z73PHF3yElylltcJsSKWPahv6
h3PPPjPXp1+MhhQk6v427BGL4OVe+j2Z5KHJiQs9+NaJ1AeMpVjd6F8GZGKGDx1BP+TlP8Fo2e1q
NCa9IXpBTJuC4UoGDXYntrg8LxjZUI7hcV9PzKHsxyWRKuTetFgrSFp0Zu37VucdC3j6r6QaHaYJ
f8klWA63u/lfo+1lZiZqvziGSEr7rKZMUQAAJdUeZl0De3dln/qzh7SGATblTTmWpNDbWaxLFyg5
sUVZpPnRdDa8U9MSy0fjLCj9zzSz5tLuraAEO6UbpOzZXnHZQIp10f7VKQEytm8DMCvaZxJqjcqP
YHqk4JBa7Cg5p/kxy4EoUju3JS+CZjSkaIPcMnP7JbR8Bcel2WMWFoBUBDCC+LFScM52+9msEshi
gLD5TA1CauYIchLSf0n19qfrkQTUVTkQG/0AxcVZqdtwd/EHpLfbEAOPR0jT1Wk3QQQIkAgTixzh
83lokpAECs3otMrXKf4O0mlA5dGXU8uyd5iGX+p4Yg6TnpCb2BIStz0eMo0AMe/aMXoM1cPivN9P
K4OF2FYjoE9OAHFjSVCx6Fwbj1nqAagWKktYXeVgNGoV+xJJFiffXIc5hZqwIYe6n0MUMp1o3AbQ
MaIkFNaSdsoR9163ae9iSWDfC7CjgRyIm05mKRCO+IFzd1ez/ACRKdFWfW2roQaij27iPAbwIY8C
GTMer3a3NmjtOz6BNstnJ7Xvhx79KGt3tLzFB4sBTvJmN4xJ3HT1GMwnmiJ7nGzQ7pO6JEpBu+tm
XmpAgqMITn61HIAhPk0vf99JSShB+0/VhxaC/Y4GmQPL6DE6N2J7s1hu8xxwo7cIp/+GwF1zi7T1
uyvFZudsCkwJjBRZIYGIsp6AYxgZu/wI0zRGI7yGG8fS2eJGtc6tuZ8jp9o996S4Cp9WQFfTDt8W
ywbH2dXBjolEDy/WSUr3bjipM5NA8JFJ6tpPOGyex7WwQd9iRmUvc8ZWBVNsKaznziIDDIwOcg/c
Oh/JfVJCXcsr4fswlMqam6C1rXEdDKL6YUqnRl+oHB7+AvGLbCxFo564QDP6hAdPdiQgq6HkHb2K
Sfj+7BdC2PTG0Ch0WTNrGIjjFSS9wuxyTk8uqjXOwqi96tNcmgXYqPUEQyX8YGRSwgkXKiTgeQJc
DjWnphZAJj2MG3eu5Yt8LX52l/VOyZr7kgKabaIcTl5XpPCmepGDKr2Xc2oVjWvkMKBofhYzO3Nt
MxVoSoAxsJdv4708cqvZYJKQderDmiKvj8kBs+JH3HgTesp4XVlVQ9ABGZUrtYgOBIoxfndF+CeN
poCSqyN3HM4mgiUsKVfKqezyah0iZ4b+RwxOpQV4mzp1s/c4GbuX34ndzeY/kpAN7aqXe+5Ru7wT
Ut0FiUB3M7IGpW/gHNr2d9AkmY1A5Jm6mW7P+8f2YR/zB3t1WhTAKSRhrEOsVO/zkcBnQLdsTCup
b6TZnJ4ek0iJsYypi7mcs5btswbu2+xSTgYZbFGhScTxXSR+oAALjLwWpltoH0lVA6GcMqQug+XM
9hsI4y4/EuRo1vNxzBlUSs34Xzh1g8TLvklF3kpEBPTiMsJZbVqEpNWhD1yZmlig3UbV9f0ULyTB
HXp0cZbW2ILniwxRGQBYkBu4kLdsF7dpw+PutY3wnnv3QhSBhpI3UP69i7kbEquLDU/gaDyzn+Jh
7AfpcAbu5TP8IHGkbAwRNMvJmUX3U17QynQw83VtgXw7gkZ6sAQxOPCsHk+TwKfa+HyAwFLLWxRp
AoZ4cGCqNr5blYjopAMoHYN+hqlczg7iogQ/TXLWPfZyf0tZoIleGF/Tyuvlu6MO8Z06yIvrECxB
zcbeB90VxjAcUPyDr//6ZfCQu9RnrvFokP3PbUEpCvspcWFRLXIOQBQyzX8btIYn+s+eU1okJWC6
VSWhMWg3vCUjxl7wU3lpBOaiBBEsXrdIVKUYbBDsFtGhA28SjfI6totgsCQx3TgmMTALmJpxuy2g
oEKq8foZ4Jl/N2SDUnJrs/HnU/jGduCXUWITJ72Tldz6G2EYlCWs2a9p+spWKji9OwYfDM6YJl7n
aCuhNdAhJDDsdCO90pJSon5gojyySS7lVCmCM0Hu4tvpEp64raecQnJQCgh2kWqevSsKDMriQ3DI
zgoWTGX8uYMFod3TT5M41Qv3Ve3xnzxihiBzV4Yk2uDQzj+YuuNPAgGnCg74uxfSolkVpXKDnxe4
mCLs8BjIVzJjede95eBMqDA2FBiCTesehGFHvXK2njHE+wRFKOXC4FJmENfKuLDkPXtlqxQ3wD7D
ocaeC0qeemwiMtPeozG/+NCckD7QxY5iCI2niDVzZdOxphR3QYsBLTQFOV6SBlFOHa1/3mfl5JyP
fUEYM7TmYFUo+P+RtufaKHXsO1eq072iLT8+o5pMS3J0TF+GpVBP+wEdWctNXmXlWyICwQU+FY1X
hat2cCQjdK2FC122CvTJkpndKYnQtfp8TRe4mHZFKTqUZH2gGTyfEaAa/+H5wncKbzePTfxpCPYw
Z/Vnpuyh6TBtUhA8+SPFM7C+Jm8DV6h3QB9lwQx6bqkTQL8WLsCSwg6T9JFLXNjrlGesaO55E7iB
q3To+o3/WH0yfa4k4LVvLVY75lf4XpuH0E4k3vTSEho2EN2qhavR2YkbrHlksloW/bwt9OZ3D2be
Eh7afbxTSFTxzdkphoNJ48ymKCJgyVLLZD+e50SaC25CseQRZx63AwGxy4vLk5A48UzzxRfJhBo5
ddOCHo2Moc8tVoYlebeukBahK/fvvvp0/OfI3XvZhSGU9hMiehIivGYWrIUKj/ThneInskRN/tE2
MoQN4UorG5c69a+2KSTpG0iItrUiqItcpp7xddr7EwniviXY0/skS3gadEKgAO1JdRg8/V/GuKXl
MrSZ/y2e3/VvM5+/72sDl194xiSvi7745Tas320XASmqIcqXkHJclTIm6tt7snzlrPGYs1JAY65b
MCryvFK3d9KnWlZbJeDih9DMujZzanOqOR4v0rxLrnAf2tTdBnVTSKekUTgQ0LjbzQ7SYYnRGadz
1gmx8w9NI4jf1yD/M9dxilkAYY1gWX9PsXDKcdAQMlVY4IrFqrud7iQ6fSUBjgBRaMuAfplly8aa
uppPol29pZvDpyPzadcsKafuiQnuE8uj75I3Lr8ENTY7KU8Z2eLHU5Ap0jXCdBE4vTPLv/lzSDBl
UrdZD2k4fUB7XX6zK845Z32yFAEwz4yW9jczfkmTa0ppnPvq6o2BRJ7dvHBlX7uGXspswIKr/CKU
Rm/0rdTnYKbMx/tjVpzKeO1kCvzPXHdgVOy1lvpxPArxfUfq7jXLm25DlMQK0tbh2jClOJUzxP/q
k+euSEEw3kWQrgVp93TPYJZD2vTqll5qcj/Dm5gRn2/aN/4JfH0ahRWIJ85kCj5aK/EobkSrXQDT
W6BQQn1oW/CRe4V25mupE13cfFn2LPZrnzZVB5ucVuFiO8GNfB6dVhH0au2waGRR1NbYTnO7sfLC
esclnsZj56ddRj5/fELWhlXAsvDUGgxAZ2pLqMnojI+IYF1OcwlJz4EwgKya6TJN6agbmD8gHvXC
nnLTgk3lLxdlRyJOquTDAFDA3pfYUktLkjL2/LgEwX5FNFnVUFJi6VFNPpB6WhL+5FfuzBFsnzrw
s1y4+xEgX6PX4NGd9yrjjbcHlVzJ+j97zXER9JWcBZ+eXN+cLvEbTEIRS/mQ5EGKPb+o7m5PYgNr
bMOnrEdjrg7m+iwKNxBorO/B8DgzRv08hs9cY+oKpehE7RbvEXPQRKqgrWDDRME0dJtXn1tx7MKT
tHMrGxn/Sq8oXg/a8yWPUEM1gGwxpHs1ncMGlM91R1+mrf73IBKlEPWQeBePGwgKXGKlzQuxgwMc
pGp6YaOA5XLQ+fehAnnup4UNxtHRMeDrx8eKw6KSMU2rejONv9sdQADTzgFpAyJCjaT5Qp8LriA8
rLqGRtpg4iezsXc7ACx8XoI1tQssVvNp2GTAEsstn8aTo0lDjmc0S1YAB8q0J28YAHQ0PT9DU7FA
2KCiI5/6tjS03MNlWkpKniFCCL4G8jVTIIm3DQtrP8QEgCfhTDzZhgZmwYEFB2zGa7R1m/z8p1f5
bO9ZplF1uyXlgo9x9qiQJjv6lyflHXN9mx0zm7OchkqW4ZKetEZvJt+SxuVynfwkI+ciYeyei6Jh
1xVNup5FTFYE4yF2Y+3063aAbvhp2UJ+aS8bG1QDNh4MQkb27y7UbeaExfPT+t6/Mpur/u7a8oQm
Wsu+uWf8CA77LXdnJQKMqUAaqyAwnMpmX2B8i2u/JvUjHL/yA3Oi5jwoFUcyJHRe9WumdcU2SP+m
CwkrAEOCyfGiADKod7TroN5goPgWiLKzKvYDRy7/Utabad38JXTc3ANN9A3fNiE9KY3NeZ4rBmnG
b3F9zRlrDsUiEhhA7yzt2RcCYSL1bf/dpTQ/nOgzLr5w8bLfkGMZeCF2BOYJxtmEgi16RQnWRH82
A59/Jjoxhhd51QmkyivdnVAKsaFgDWKuZQLYdzlq1+DOJMoHgVtix1DlzIFSk5TTlvHP/Yr2my0Y
aQocDXNvJ8v30RqK0zdKafYY5o/Nia9A/EQJYo6RBeR0sf1+Vmrp9kLGJln3FHXf6g0sdYyZ0s6B
jloASC6WOJ69t6l+utYEREFWGhfXMcMfGd++L+7ylpMNbgZI8fL7lcMKv64qzl2NCYGXhDnsXTvP
1UAWX0Twe+R4/Etvz5JvpEadlDQ+pB2c6mPCbEiIbLMFVlrzijnnWYj8KxF+peMM8PbLuy1xY2Np
zMGyLqXVJ9IpWqbEi5yfNjxyNm/ilaa2etiAkmTcEpK2HFyXOf2dV9cwlUEVTOsNJyapYcSH1jJL
7eZGU80N97kuqCpZvU/5qmMF5TaMHFusT3nfm4lOX6W9bKkTRcT9ERX4MXHRpef/sgcePxQtuBOR
N3Nh+TOKFGguXZMHDqi9EuMO/qtE8fN0bLAYAA8IDmWnCSzxH7BuYyOwF+jq8Hds3A6fZV3H8RWP
/4gBnqkwK+Ve9B+lU8ZGimSWDSDJ7rSN7hhlA+pG4m7tSC5+N/RwaBynj6C4/CSKAtpxipDMrVkM
nJJ4eK4MO0ZJJs7ZZYiLOoEGmm0iJITHlN45cme2Rhj993pD84dzmIc+xdWyv5WiYqYhhNa6b8RF
0AucDbbFrYekZXIf2RH/9yniBr1QKWaphUP/1XYTEdgt84YiWxeEDw5MPhYy3ffS1v09jG/vLSKa
7IHUg7j0xe12tAhKGyYNNG0zu/qNj5yb7sGqAv8JgydnWkTlQKo0qKMgl9DM8waS+lEWfllCLB9W
UEYBWVWiKNVKRy+a1f7nrS4S3F4MfYEGtcfdgYKkO1oSnXqjkG1P4efYKimo+JY0KJMT+wYq6mvc
7B2Jq97YlycRLOgusY31HmOx5nGFkdzdpdDDX7TlMJMXJLZhTDDjKMMHsXur/dSHn/jtwHKXgd9a
5R4p46FDfKc0GRIIlC/ZNRB8PUh6xJcomlZuVMNUPqNgTVOptaqvG+6jg0FnQ2mIqQVDi3JNzDE7
PphP6xQPApNXxsKbJ9xJOMZXcMtRrCBsH3W5icaHwt4D9IG/sL4yqGNJn4/RmHuk9MOTQlYlPeao
L324pAV/5J26CtVYy4YjQXO0V4fE9y5HIVfIdziV1AC4JC9ogukbmc+x5PBc+5Ix3CEQvymxsugs
2afTAG5usvNNkNeh4Jcs8CTrqAIkDXUlc1p/Ej/wqaInfJit6quopegKW7RAsnw3OGL33fSXwU3a
XNXwB3uf41uiwfZ0Yqt9uIn3tUzmsMIAi0f39ZWGbrVtGIU=
`pragma protect end_protected
