library verilog;
use verilog.vl_types.all;
entity and_3_vlg_vec_tst is
end and_3_vlg_vec_tst;
