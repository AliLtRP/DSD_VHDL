// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:35:32 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
G8yAIVhGsniV/Ik77BiyXZq8gr3R9ZQE1EqE8TNBftreOVsc38KxvoRH2oRPIipM
GOS6KM36RNZdgJ067JhGjbMxENXwZntUbueecWJE9mHQ/t+z5rsFusLC8Pfx3LlZ
wM2XsdhOczWq/mfRhbW5Bs5GhgYLU0mbfUlJPFh8XUI=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5776)
YEfvMvlyUNXTZTPA4/EyAu+P0735ham6Az/VIXuf37o0zdpBJReJlaZZC+PGBG9H
REfQizboKBwVCs33H8685sJCV59rZZlzwy+zwMef/6EX1BfGQmEYYVcF/yiCvqeu
WRtO6fOO8y7k7TWOIrLWl4K0aO0+OxB/pWTdBmc7x0Mpks+kFZ3Id2v0DEsNvbDn
NIHjRqZZBj7q6weHSDz5KWKGvBW979APeaMiPOeO3hQr9mC1gGNZccc6HH1WoZJv
5Y0YcntWv9zWM7DIerxcM9mfmj3HA+xjafXIRrEtVtZhqnduMiuQRRxM7hE53k5l
BJKCP1jJkhHBCocNseQb3QMXgJNwoZuR61NxXS9nE/NIV294EIhm21b6MAa71a+L
S+Njf+sYzp60nL8WT68KPvty8TInOy6aHu0uV7QuE+wIgr9Emfw0LNpGQrBPzWOa
I5MBPqvsrRxkJ29ryTlHaFHJq9h50H7Q0GXmjPDrkziy+jNTyhSUEsn0awlJV3RV
m75FkDJf6hCLaEBZx2paxXV1iqA5IjC02RYjFvxQaQ9knbW1qKsn9xojCf+rtSqG
MlHc+saRxq5A0dGe9Fm0rl8IMVOeO8QXRL96Je66/FbHPfL54qDX7Sd+bBZ3+dKS
cQzu5/u+AFIgsWYw5YnV5n5JPbYpcK/KRDQxh+8+nMmKwwuXzl7bbrKtaiBQvRUR
8sUyahAWsMGXDGv9xvXS1iyuVYWABxPzYNsbbbWKZu6fgS07UHXCPy4/fksPf4i9
hi2mZbLb/6deRqKgyy0PnR71GjH0NILSZtGJye6BHoZuVllhzux/zsY4Z0nC6ORU
XXVaPjTzR+UtXFWFLygLQZCSMzQDRUHowtOs5wzh3Zl2TpvMVMYdKYplVSTO7oWL
ouc+2bNN677PzkLP499IOwd3AZORgy05qAppiNxLh5Ti97id/gP7hQEzYuJrcUFC
75enct8KhkVXcVx2JV00DNtfDb0UtnIZ0bH4xpLv7j1x/e4wovGFksTh7lyVo2R2
3Xk6uGr4i31BErBm7Pgia3N8h8C/rPG7O7xQsbtWK/jbOGYnyK+8kFd7o5Nh/ZK+
UTOKr2O0suzD72Qh73aFDCVc22DnGcSjotTXDqvLlbc1uapcMiax3SlPckmX0UKd
/WAYIyS3f0QK1JT5aLeJ7QUYpOQqodWvubFbbqZ1mt2uoa+Pw/sbZVsdkt6/tBuO
l+ZQLHc+jHJPiDQ38TA64jDUHQA02KPRgInqZ8LVK5iU8ijYJVX3bu/6da/s7NRW
kSbRKpLdkJgvMNxWKObqIvrdEizH5gNT5gnrqm5udjLp5ZLZzhgotOlYHeVig5K1
fTP73skcRJMDviIfSH+sE6HQMViFw3INFCYIsiMaQPwLWIEAbEIymhbKdRK4PPin
188ieaz2sGHjFBkoAQNfdUFGHb5nkoobf/yFmCOAKsoqF/zbiRoOkwzxvPI4aalR
VdeKpuG/Uq/LUeU2Pnbmu/kkbK3HpkHk8FoyL+X9L1MFNo7uIszdXa+CSwLTTsJL
1qgLEP+aapk2jZewVoOw9IdWZf6+PRP16ooPry7Jes50jTLaTpXKKk+MQus8MCki
ObfnvNuPvsDiVwafQrdON3A+amsUpldHoz6bBuDw4Ch84QgiONm+DNYNFRcbylAo
7EjwjQfl9jxqLhG/eiJJzJkUSHZkK3ljH9qPNroXsXi8N6/Y3IUfxqzpOLQDMk7E
Igz1Gx63njdCWuzG3vHIP/5QmvG8MLbbQH0IdpNRyreERbAqqpe1VwSLaKdTL06s
oGkNU7B8SaqJNFD+MWzLdWzPwd5AW2MOveAkrpTZfjTVWyW1RXjY6NYlgk4HXKE+
2KpIqYds+LDHEfWUzJfhlAG3Fi/FAXGobksMYh6I9/JVBNwm74szafE6KsmPBTtM
HKlnfRP9TbZI+TOUX6fsScd0DLd9smRFfL0sv9/pQOcTBbAj3Kwemn2hV0Igoel6
xJ6V1zQkOiekqJj/a5L2a4W6qgsKh0GdLC0jQC4topy0Si4m1PBwPjdKZuBM+3wA
jgOXKapOHnF/MajW10uj4EkUUDXm1crUWr9lvKnFXD6gSotYQtGfWMrOSi3hRvAi
frc2BUqXRU9eEK7jyk+7YD6h8Nuvc2/8gubuBBYHrPj1lS8hGm9vo2GuepoSjFYu
wvS1NdTfVmY2eai8Puoso0f70Z54ilyiH91yJOHvVh4mfu9hVU29Qdz+ywWrF1hR
0Qs2Onxzst32bdQq/TTs+e+5ikcR68yRYCG3uNNmAr9WjVxGKiEACFVrxEO3rgo/
opomluI7DjoTkvfczlRJoHdVty+Ak6NsFT6AU1t9704+X7/0rTtt0wLkUGfKqinr
S/lytUIdDeMaZg44oUCee8ix+Je0vCT/15qD1xhhfINJbk10jg0pCJ2prgpxCiqc
+a5kKCBjW8LRDPZc0gTw3X2Kji+mC1SDZb98r+byMBgXCyOPlffmHpAP3UM5Ernl
Sx6VoaNDPiiSf8WhxdOhNamu3GJv/scPle8qgOGbPSaFCcz3IO07/vq9E/q2QGw1
jVFC1g7jmIge5sSPr5cv9l/nNkXzVtmNPy+U1Prj13OS1k/Cmo4838jpcOOcyLYK
Jn1DKHXKLW8TFEg7pnosqTozUuPxu2x1Hny9H8DAnEGtB9TQeToasumkr7fEXRyY
rFNBx9GDqHU48riks2lW9n8UYG10AW0OKseDtFCjXjIDr9SL8L4w4+HTTnXWzQmY
+PzT9xZWRkEB0qUKI+A0ucoGoryYSpyYQPetXRYrXEtdaHEmBv+U8YHwt78SxzUh
VRDn7CVGrZT04pARxIp95pbu1Ty2rk/hTYGOPjUYzmq9Y2+iSjhqIkkCCnw4jBMf
1qIvxQ60WOTQDCdaA6C5phAqMPgS+sF4P/McJ7XrPTx1vCPixkV6UhVYv7nS9pTx
lQ2ohlbn5z1yWEPYNqC2k/Bs841soDJaFvKlSufvO9q+sOVhS8ya8UjoMHkeIj94
KbWZynypVyM8mkEZ7G6jR1hVascamD8Z61J7FeK1gMNDyyCT2aatbZyxbYRLVOBt
QaSGcU2jarJJgxVPfd7zAzxGfX6ZCRleiU7jocWrk3f+54tWi6ZyQ/IxvPzGDU5E
tKHnrOTNgAc1VK2eSDEp45vqP6mw7nuwG5v3eRZYM+2tQw4aLui84IxYmAhAUay8
Jdt10vnkxKlf21trfhfXLqOv1EoSoRrUsfCQ73IrkQ1qdCLqIR0h1GvnkBrK4KMs
KryGFQP9N1aA4wK+AMYvhJEm7F7bcEgVs7oEMFjbWRA9lnfuJxRuIl7IRPsbM6jB
lwzyUbe3dKfTMW+grdDSb3cLNif86NSJBp+ils31b+sHmS0cghVmg/dQgnF2Rdmb
SOcTgWXoCsr3VSBWefV5yp3TREcyauQ/nFUvHjvWu7EZ5XJ4nsiSVcPSKuveZgUn
uckucRXB7IZH1y3i//C+2QqYChQFpsjobr8vj+jFWKTz32kas3g8S4eyWNZmsObv
jt1QF86op0bcs7zhDZ2VNc4wo2m7HKxJtd3cpvI+/iT6ZydTdcMJWO5BdC9PLwXg
II+rqvx/fMB14XNSzgv3PWSyLL99ZsPdfcmDmhjjdH5L2W5f8aQuvZn+QaBJIfDI
T5KZOkZWzHgC2wNFGOM6b3CEjQ3eYB7P35Uq0d59c83TnQqkI6aIpCoHHiu+UuHo
oRwkmPpdikSFsZ8+or6hgA/W1xzvIr+ivfNboeFbTnCgJzGWWCeD87Xy8T1/tmxN
ChHwENN8LvB/MmnzWyRpycLw1/HcBfYmMgfwj1FI/XM09q4VBXjjqPzmRPxRkHGh
VzYjdNYtY4+/ed7xbUMwH2qSFaoFPa5Ok1E3Ma47F/Pqs9D70Z1aLuGjds/OhrQg
SXsvBNadik5ByIYecDXZPUfh1pyzQ3E00qVz1jys8IevfqJ0Nbexd3hl6aS6tFUx
6TeSedYCtPANT7oTLBLDcmlDm3/E7gbdJ0hGrB2LD+Uib2AbOJ02Y3u2yQg79N1g
mL+4MaCyhBCjiptLsoIV+DP2CNy+ah1lQOZVWRpKZspM1BdAGiBnYEtmWRNM2jw1
Xl3VuqXXHmURDhYXwouLwbXFOtryDcRH4syFjfXFIAXDLuW155ToBppcmvIk0k0m
9Jl/XblHJn2Qs+gId1FYb0HaIDQiQTuNeHuDpgLpJRLzFE4DtNcvY4z3WSsogUC1
XTxiqlW/khMbB8UmqbSna082ZKNn/sZt0zEN/jVoNfdxBL+RkTB8YoBRvtwLkPt9
/NfxO0P/PAmAd3kUXp9WAM6OMolWQNUJbdNuMEFFYaJ7bQhqg0ia/VbxHGFXUerK
iBSgCQp8MCPKdJs/bORZbkzoc2yrG37Yb5U7dwoXY7f7EmafMgD/xh0uc6uAUvib
g2jPSWhPQUh9bSB0lAlGKUGO2f4rUKfdgI6kqQa7HXorXmgTfDhYUpn1YAqibvB+
9kLReUs0+eHV5cbs1GbsFYBmwsQZNx/09RWDvyJzEkZMQYf+yeOrNX+zpp1YMbXa
Y10OX//C63MXOIftv363Dzst1AFRPnGjgiMamKk3Q3ghrs4+qws87OcaEH5fb5nP
GGmpxqXIZIvwPu9d3F+GVF0yNqejUBXORfuZKupXUFLXy9ZMkS4RWC3i2dhFUtsz
AGBarct6tGiAYMCyxN/R2M23fCsGim9QgZLTQGVIxCNbRJ+ADw7E88SVJHA2Td1w
qtdaaiOeDF9eZhb9wbjxTa+ylessiK9jhQRIJP97eLP8c5jzufGfQ5qg26GQNsrY
tTCBpiwb+1C4lqkfOfVzP969KPICC8QNMK8ADt3V//1g7UTbWykzPZd2rCA5A1Fn
B8AQlyNSTSLPxRRVY+xQbvnFVmxVSppnzlcdbZQMCI3X248H7FycOPRcSKSGrwXN
Vluvz7fs200k9tr7YH/HZhLA03is3KIO/knssYUVzlxiHQoip5UFmZ1PjqNTayT3
XS3tImvuZT3sT8bOTsOB5KaSVrF9t9qvyxNJqAwsvwJcRLHefFDapJhhDyY2TXaL
iOOD7zewNXKqM7bEF83L8Fq1CsJe+dhXbx3mY7bfov9pOu+22s2J3WZrHvyCT/h9
acqTg4YRTfbslf2smAEAEXgJBSj1b10Rqb3H6OBLtF5k2a8cdSvi4d1a1Ue7d8lm
fPHGBtP8Wd+eDV6ztZjDKrLrgx0ipq4U5qNhC4iAD77UEY3dn4M1hqStmihUbuXW
te9d3L2yMNN7S51LaG87y/oMr+ReWlpwDVrVojkOBXZLxKsapc6IyoLAZdN2Lk6j
iGzv5RVu5JmeJP2rW+nwSwpwYy2P3NGdW3y8SAYEImkVlBmEgdMspVvn/hDBrXCo
AYhciCK5G+Xmp5u2oJORNiyLaCJE1AxX98p0Je8UHbnuCNvaQplfo+e7Xj1wDIPc
ggjIxBbQH4mOTTob1r8yLiFLzOspPLqKdUNOZPtN6DmkJ9org6f/LVMpm1wCV8go
nYsAI10fmUJVG/knLqT7I2Q6v0nk+jQ53O3ryxRVC7AHgUTikwAhDOGIM+j6gQyD
xmegU2xIahl5v4WMrJLLA0pYlbTRngbTh9uKW12Ez0uAvKkFgQzOhfbaBXmnTA0u
jb+55a7B4r8ioqKQIeC6DkCAMEj/AP0Etz0+FE9eaf2LP9X7z1RRVVAOsLryYIwJ
f6B9fLye7pdPHhRm3EETzqx6dF687hMsMByQJOFOImh4BAyIKsN9vTAi9m7OTElf
pHhE9uuOEkj7qGBfTX+vrT6vmVKfJlXfTB320MXlETIr3cj5q3bfrowsLfcb3hjI
QdCcbF36ALmNPyUyKZMsjsVSTZMcBI1/jTnyUGp86/43UlDC16kx7CI5N+aXlsjn
doYFq9ptOlJQmYYeppqk+df4qJs3fcMiCYJ3twuXk0VL9MwrC3UNp10d0prw6iSX
zDQ5FFp8PONfDeWwxAwahOV/uSi5ES2UQPVnuu003DGHDBofpSxGnPNKD7UeIX2g
dm5HCUxXNvUxPj3QunziKD8SA/pATU1yCE5DgXCzNi6mzeBWmD3q1I0B52L3N8R9
3Bes4mL7ZLCEkLhYYHYiDJP6eFP3+BnYK8HtBNcNOHnuAKB+QviObpdJ/1vGJcsf
edtIZOV5wiNiKwjrj4HzPkgLlvjbjz1Dak7dJ9MqPmJBr8xOEnqz4pMYpMKLMZhj
TL1Ee/BJekDv9IxSqigc5Afzz7TLDKahCekpJ7U/cGwXKr3pTphNj5ltGHaKTRak
voTAFrJa0+WjxgwbVrsCB2/ZtRy1wXbexBRGv4JRPvGUhS+r6ERuv8ewsFfAITVE
CLULFDjoZZDmatZ+l0/eFmeOs4jz5dczNFguZpoTAYjx4Vav1E/LUK9dyq9y255s
zvX3OlKL0VmuY6mA1r835XKQNU8f768ka10En8gBiylRnFW5fUmvT53cVEgwWsA+
So2wc6vZS5AD1J/Mg3SdEhTqCnq/Xw0Xq0H/pp5qGrjIdmIjSNuVyVLImZ3LXZAK
1FLRxHsPw5LRFLAec3Tnn7IUl4V9KrZAnvE5lNwyvRLqZaTrfaZgzRhTQfhdxVAY
G5e+njG0RJoAtXW6HUVzgKyaenttlSFMA/Wa3CKvGed12uHHIjBFGZyUU4ZCncIk
Bke5X0tFiy2Ln5PqWSDoVb6zo++0XtXgJHNFXA8FigysUZ643A8d55FhyibBoldA
HtI/e8CJcTaM+fpA6bY+9Dip6ylZgWhIFZ01n138GOHfg0GMFcv0x+9rcrI9J1gk
8s4ztyyCnPiquY6qyRGCxsPEpT3pVJuZzxH7Q9Qi5atZ2SotYgc1i3TfjLEMZdVQ
XbhvZFCLusm+4f/iMRoVaL8xxQ6Hhk+eHCErHzIxtwaHsoXRBHP9PleM3B9XeABG
a8NDVlOp+oezgF3glh1//VddDdu2L/x0s64tZfjkViDQcbcQohLo29M4WSPWlk4R
99rft07DG8iZnzuOGQcUFQCIiX0HXpdud8GRq2CYTFdbO0ivvRilCKGzYRly5XcD
bnpmYyz5Yv74lU5NpIwBm/m4am5jRuAbOmRehViyxlnVi5YcYj0vJSTqhNYa+p6q
K9M1v4OVedFmUcxu3lnEfdj2WEl6Dw+VEXoIFUNB1vSuyprCfqqzFFPSF3mplgg1
CV/jqM6pyzQtaynsEe3Zq07aZaOQXLrMLrTs0kJtY8Yut+XEfBP58dnP43pceD6W
/FZjFa4KqwXXJNMGjtTjsutpQdCtAwFyvcwXLYaNA2t2sCnWxUS8MUVt/6R4H/ji
PUgM42zdaw1fijfHfHQqzYTSGBbc3GlvViz02IJouXefY5W5BNyvR3z6S6fzzCJd
bxtGWTVT8kqqyQjrHWiTajQZycHpBHOdCHGx8Yx7ddpWjNpqvcHTMODfNsyxQbdQ
uAYDPkbvWSBuseUeoLmHSld9YnVajLiiY6VTzM3ec7Cixvfg7ImCYKLcLrPEEBsT
EigmFNFrihYEZe5RP6dqQwZxLho2EhTvbo41bLi8dRQLu9yKBLpC58nPBmDuLY5Y
VvzlhZ6414pbMxMN4BAiGL4vHmdilffi+FAn03LTvf8zz+HJHSvfTNhQ8Ckjdora
ZIfWpAu+m3gYy13GUU4gE2GCNgAMrsgLs/c3sLav5I41QGCRws8bJ9YPZGrp2F1K
gcvjSc/pjSVr+sZBkueNwQ==
`pragma protect end_protected
