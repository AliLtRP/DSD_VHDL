// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:35:50 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
OPB3NiA5Z5MXgN2S9Dr9OFFItfCFwAuTdR4jJbllLEmeyUSeR9CeD3SqOsgJBWze
+3Niad/0cxKv7KA/RAHFQf2TjPJohTsrvMb0P7bY8z0pM7dPKjQg/BtTBNC2q38Q
5okq6VzzU0xOCB9XGSJv2hrBG0/dnTBSK2zb4LhlF0g=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 3488)
rPwISon1WKJodT4ZZQbF0MBAkvL7BIsiA2bJZpeHAjFnMlv4mA097x0MZXfsMaL0
cWj7HEez4XZbPihIkWhiMqF1vKN5sAHuSsGJNftGONe5wuS4+M/B4g13B5+YUrYO
4Ln1TEoWTFmT5WDYLItkjFpzkDsADp0/zI5rcTGK/kVO4cBSVMSutx6EyYbkDBi+
p4ubqiIfTGg3an1KcEXrIho2BkWe8Vy7Q3L32rLyn8uyL7JtfyHlK/YWIdX1H9jy
vgpkJSZPVyZ+xnCfV7qCmd3lEpNo1vahGddSLW8NYqyjmj17+6CHigI5qGZdYp1d
k33vVSlU9Ik9chp/0zmPigEiOO/z09/hbQcGLFteOnPkniJo64WeW5DZ4RfGhJMT
RMGyCo/zjXygXbs+hQV0kuldbaNt1DqQzfM2eJy/SBtxwW3K4faMiruD6eZBNRbX
qV4J09Fv+U1ZNM+rVVn0vsZk8LDAerblD7421GavoONwnRs+AnwI0sNJpU0c0itK
7wQ6llfKH8nc1aI+p+aC6xTaXYpoH0ixusr5fcvAl6yOm2X2gX0vW5hvlcAxlk7A
Ryh+gDqhETR3ywv9MS1KADEXj3cOt0tFdyj4LqfyuZQQMmnmV/Muc9vQ0Eauexop
BshOOzGFcZyGr7RTKC/pbmXnox9ZPDUGFW5boJwhri5rBsdFhs0vPwec1NOdeNNt
aGGMNLqwp1ncHZKympncfxSSzA1HQCpJBayE20/unDry70yDDWWGBzMdiIwYWc5g
g2Mf6Ogtc9ekzW1MTnfud3ULmSsVMwLaZDd7pIpJHMQMGHpCkFYY1eZbWjCRbuGq
I9cXbZ0o3DBt7HbDuL//hiqRKsYYgXtWiFqBcIWVqIn1RKMYA8i4F0FuZ0MSri88
jDTDiz5O2WN8kuTts19gSdZ4079J7j4wbpRseLFLT14xfWRMmMxg5Gjs8QEX3D1D
PTyiLz3uNcVvqLsLZh1U0AHPjsKlzO95MA1zb6f8oOKOzpBxd0B/bQGsYAWZSo+A
dvLXyYsXdPC6EbFrTIfQveyCLsQzs/ZA5YnnkMqozcWUrTwwR7ABFI2pS21Kc5tQ
2m9qe/vDvIVbzstBrCZv46nxgGX607rc4Ov9xy9qKvhyRmfkyidn52HJlGX15C9X
R/p7sRbS2gybqb6ZSdGRUvIrg26yZDrMWIvu1EgGUSVZ+J19wj8iv6G4CtzGuu1k
MaALvd6cSQrnjFnb9adobf7pE7PjiC9FAAxpaGgYSjhZ8nDtNQlvY7SbFM/P/nAi
bvTdx2RKN9nVKR8rA/m6qdPiPBHlihdsPsiICeDsCF46lDVBV9TCFUWecep7Whx+
yxmlvZV9ErTu/+hJ0XwHVEYXXcarufG/6Dnoh//T0rQdQa3WGRkPf13RGMRWSq/c
1waIe8X/IaUg3V/E7c25qxet+4L7YgWKtI+HHWxZW+JUqOaHeg65lCZBgJzBgsH9
WMMsV6XP/6nNHIBabkMo5/+F7UrqmOrvK/ntFuRKjRaNjnwZBgiWsRAGcxtEQ/cY
MBrpbeALorb0oLE9YNhc9BeP9+YRVZO4IVWygg3mPvIKq4EXRGZjqu/2dlmdnu0r
7nGB9MqgkSltv6hFLem7dG/xHEfwsI4kYsSa7qIkcRbkIQUHImZ5rwWKODIRzX9n
GTNFJzsl+o3QFxDd5Jb66r3VUh43T9/MUV4SLG/u7CkSD4GSbFzZxa+flD2GCCOq
Ol95qZi5YEkkFGBurKTFIRCQl8UmVKYQgZj71lj3T0pUN3o7Fc82mVdowcm7k8Na
sIfsraC1bcKEaNKof77hQsAE/tYiiF+m9pRqMrbrUHBJe0SkGGwDNKJyhIcJmynJ
kYnN1F7wIYBRJL+30kPbDtY52HKVZIe/sZkl+8sqN6O3yi00ixbgItjsmTZK1mwy
waJVoIWLfOyGHUZVSNV78Wr7gWYqmtxXvgTHglEwZ3ufMWfPeozP3SdC7aDqWbgl
U8pmu9cvA6pzH3JU/jP4zAYmwKOErrrxW9p2+GnZYVsJ86RP6r8IBRPThcM51GPv
Cd9T/AQ9Ov9EhuxT7zNp5SokJPUAkgcK/D8YZHurBBECgc2rCVvFmsh/04oyHoh+
qsHlV2qSg6MNq6/Qv+kN0GYR6TQ1zWsSORvey7yJ1yxFYcQ6TajksWWphaUWu2JP
NJubANLF2KyVSe+c7xctx4gRnnZM4VAPSZlQANyzWYT+py7VltdfbH3mImy2ZpyC
hit7/99RL/P1amwYBtJFgAg9vyN15sn+WhyHle717j1NaF0fSviHz57Wu3qQQy5O
a2mdcK8CbHTgCx59OeGdLWhabd69UBWLha4xN9q72aY0SCTUbGHZhsXJiYuokn2N
uKCC13olv73bvvITk2SA70cy0qsrLXcK84t0MaAk6dVNBhWf8fKtdwRZtIfpZjh5
DwQqESHzWPJI+Dsip5yFgPicohpYGQFtl3r3AS4eNN7OMSEUel05wLmRs4cj0ADn
0UFgNmkUtpdmPojifrGzmXvdkaDv4p5M8166OYVVtyDZWyQSK6IgOmYqqTwj0RyE
ya7sgriomOS3oW2I79mEB1cigiw0Glx2RxJ0F3RoqYR/G7HGjlbNsC64fnFS28oV
OQz8iyhnEjxRHK1bj63HBX2Eh7eeE4KHoZxvga9lr2FB2sRrOYX5oa9Dq3rFhgLH
VicCVgeUuZ4t2xj2Q4WpuQMLtrmigmjMVRdspF0m4SFD2GdB1aT5DTxv92RAml12
4+eNAOaDb764AA108VfIP12GBN7TQGEuSx08qVbT9qRJBZDIXX1Nae20lK9v6qSa
VzLkushKq/AANJLjP9t0EMFmYcL6HQx10BpnjV30MV0+kBogizVUVvS0f347aGVa
dtCzsq0jsOVGpA0QnPNcNRWMCrXN6IB93dTSMHRnm8sHfz9EsJ3aT3JpRVgIbSDf
Z71YZ6e8rowHKZ4vVuYZJbAucpYr3bLIUsfTfU27KSgKQapM3pC0JanxtM8tgLkS
OCaE6ppvRwmsi9Z2uoKbN/JOcaxxI2hcQn9wY+ZhDGULSRIQ4sLZHiOWfILqeHxa
nMM4t0nFvH9cW3HjI8PAeuvTN0hx4ScpGYtTdtMpx04vxbQ4qenfQeU+nL9wTOTd
YrQlmI1nMoYRvA6cF5iybyp9LBiU64ll4eolVueRbXlrH+6vUdm0JXotc03rB4S1
7LGp/iVjEnY7tALyQUZHbcPm4RSoY35WG7aPYz0dVuOYFQxopN5kv99y6KB7GxHM
wN3BD4dEyDaH5tnksNu1gcHo9MbppbY9uqmdEIMsZn4UjqAlK5ZEgnphjuAp+OSc
IbqFGMtJxO/6ym4jI+VLPb9DMkNoUYAyARL+7K69rKgtji9wafopSYkfXuP7syBv
FKyZzfv6qJtd3Z1GvdY/A8iUe+oedB3jUGK7qVsXhEYK6eIjAqVEW4na6JDKsk9f
VoDpzC6/I6odY4bhG106HRDkdTOzEVCXDvTF9K3geTCv4EDbYXbJt8dsWYhZyt7+
DdgBBvR6rgp1p4cp2BsfVeS803Q5iHZFPJVbfbXmollnLQA1e3LTtWvJJiDXCYFO
dPyIOON0DQL6w7zLBX021I8Fq27CaA5KuLp0nQkMWsvcrJGvgv+QL1ySsOjaQExN
9oDoYJgUQuToOwf6uX5q/2Q5rSMTUJn0qy6yk/yEHB084dAGTJz2L8JAtCylLYN5
NzxAzqzoFdO4SQiSiOgEhqdyqE2K9N95GJryl8FlrT60+skeApb5vp1ATQI7yzI2
mlEKDa5ucctBuox4z1OcBmys/seDrryoILtmM0aKgON9BIqgOWCNP+D/ibAS7uDC
alMIEfsaolaS2W84SzjZy40ViBNd/AucoXCStEb3u8MklBpVWYYqx2dmCRuoHnKA
68njyKmNC8Zv/ehswBlk60xyzr6yTKuG+42aowa+jmcX8pPlyGZmGFjQ2oTlPiM+
2le0cuDNIAb+kGcXB3zPLd99A/CPufYsaUX9wQ3a52fkm2cGoZGb1D/kxyQOZgmL
EFXD9OPmpUibjH7AB7hoRkt7aHvZRPIoQZm1MrIBFdYR94WljOY2BrQbblB8H6XB
bGYQ4A0TG0/vbznA+8vFVTogsyzBCSGSUoBsEV5/ju239PFiJonf4kwSAd6tOxuk
Pw1cg8KGWrc8vOhF6ysl2YUfAq/oqTaWgKSCl4Q9QRdSvjgH2WXdiVPMbgqMqHTF
T7QI6AreEWkwazVZjdtzYJ34TEoDDtfV+YkgID5V/vk+FUalrwH9MJu/bkJ2fASB
i/y2sEj2vivqPsa4AQEk/01yI8ACPH/kaYF103p603O0QE0Cj+odFCa/ghfSuDls
pl1hEuxeSx11ilas/BUSJQmHGu2e3pBWjRBRIzpSSNARy1PD7ubF+0y0QklxHTUX
SzQA+A+/ODK8rlDFFUkurwz2w3Kw9FXFr4Xyue66BWfNth1RxCCTRmWDPf8suOcl
VYRsPP/BspxxsEb+9UC3zdFPN0dTdUVs76ddJGknjfWz2sgZerNASXj0EYx3HL6B
WEJkMowXY5zykpzt/7HRohJz9X8jLhW8C68J8ddOWnOx+DVq8oukk7MXjc2+wMlX
1QayTltjg2h7HP5Qy2dqEelVjDPbNMGPlegbOVJySRM=
`pragma protect end_protected
