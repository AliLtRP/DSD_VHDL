// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:35:23 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
C+4qK7NHo347SG1iwOeYrzDz7C7oR5+cpkCzyunOmJi2HI60+k4LQGF6l+gKI9x7
dkIy1fhwTC7z//tK957+i0FVtQUfMbt2NM3oSILdx+XmDbXLBU9omxiavc2nNtlc
tmXUJvt+dxZkMx8FkKqEQHi9PHTz94YumcVkFDGbKsI=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 3264)
Zd4Val4T08mBKP6u87dcTwr4UnbmOxwv2YOf+bUznHvUW3+2FbNDXiZxjqxsJ68r
MMwvpuYDkgfbYRW3OP0KFpmf1zxPgHgBOVRW3GkUXcTU3ZAXzxZ5pk1sBuUTig0c
phtjSVRLEbf3kvrK+tMRK13KkMf6k2PseBc0qCAhAQOYsQtCLiVqKdewhtoHcECt
C8Sx/y7IOG7TC7mHQq9kiq1Ij/bIAiNYdHOz1kUvMpHdcDmkVzAtNJ2eNFmERIaf
R7450ldnKwM9p5SsD6BxvunWLH+xQt+gzrLS4h72siTqvUqKII+fywdzyBNpDhJ7
Jy+es09ESZcogKsLbKSlEzBsGF8eL9kYbX4y1D9tE1o11//cZxMA5txJ2qLLriMW
Jy0JrHjgEOCNf2yqwUB3WpeflsaR6cyeQRg9nZgESX8eb7STINGhP/C7yTN11ifF
48TwOX8c9OH0g/KCkfRfkx2CSEY37KzH4X5yDS0WWBB5lhngnkiueOWLDxF7cVYG
bQS/r7VZ1iYrMLkkMYTYeg52pfH7OaT65aFQ3OOe72tnPJeN+EtaLu2CS3MeMQrV
GITFyz7B1qr3KLgvs3LYE2NxMIKb4mZekzy0ahEz01FJbgUa3pubQnFjZ8I+T3T5
wlHKVl5qO/58LY8q8U4vCLd1YSBZC7iNsBZN0S3R9uimGB4QrZUsc6oY3bUBVR7p
dTcGMsFuDDIyWrDP8cTKeWpWdfQ5PRANA58YrM2Pr3V2Lex8CXIo+SEQRgYxm1SM
jCeI6K81X4d/DyizldWfr/vosfXd+pa416iBLq7Zxjbc4vuuWJZaz2vhu9mNYorX
0Z+H5t48XIXHskmYF38VkHX/0TxsLZwgWgjF/gcIrBhQBTccBYE44gOWMelQu4l3
XGTd6PLaA+YH/W87HtTCI6AcMARbEMWgRudXYZlgjxV9rUPFrSNh9frnfTl/umcN
3Tb8Yt7Dt9T5+n5hcVmmErTXjFJAjAW93kV7zXx+BQKkfSyRbnC7EToFrRsfR+c4
Nc7fvcj7awHYtZkHiifDhDDz8YLajinbMzcRJ4EZPd0JfUqmJmfGBiSf+wWtOWSs
vibNHkyVa6e9dDVT2iklH0/qxfti/4Bi1GzLKRiDHXpmhGJTxdrAhOWOqQseUpD2
T0SLFM2zRk9tzikEbqY8KFDpKQWLlaTMhO+CYZmHwYMHRCSdm54zHmSu6//lg2X9
OdtfUCmXSNIdek6rrqONlQRMbc0LqePFGcyzF8L3gpAHxKYhsIJtsSmXgM0hn7GL
PUw61s+AnuyAYJPyRaXSKTm08K3bjaSz1cuYr7HIwOr0zvtWRCn4zn16GQLoKPvC
QPSVFHj0TGINeBtkr0M99gKuHUNkRAd5/vfhCD3n9aXpqEnZ+G9wIvVEQ1iZZwSp
+u8zxsLSuMrJyMnr3Iu2SSEV43ofwYdtka4bjRN4mG3dkf0LTOyjQ0LvO5mvk1DX
njLoKKP7n8u5pEN3VWHyD2ELF4sEPgNnjMDXyumaIRHCQuFoVgNOMWsc5MAWci+9
hPi8psli5THOoPVSSZezBJUcFS/MaNncERUNpFFbYLM4Ifj3j9Hq3rcCdhmoF5Yj
AOdTLPDDVehTbNz/BY1jg2uPj5B1XSPJhXAighyyXOzvd336VodL/dBEto5yy65o
Y599T7U/kWGzcCfnAjJh48T9w4dQ7LAFWxIoh3BbvTEPJvSzsRhKZ1OmFIyXNCER
f3NwuOcV5mUM2oOAz9JSHu/ZHAI/pzmnQG0q+l+O4IGuzuqLPklOONm/Tnk7PbQv
+mtXYDVU86cjpumvYUxwE0iufP4+v7FIO5xAgG9Ob9zWvK+fU5dRXC+0v23GZkTg
tIW41HvsQSv9R3k+k5b/NmoJa5mdkjptaGejiGDyhwn/uNVxYWiOLleZpAY8043L
9OidMUGMAqnO6xpO/OnKLOH0PNKywu/Xz+fSk/xYuRdyrutfWBDjx5Q8wWoPRUxT
lPp4Iin32pHRNjVAzVAvN5KTPizYZfFAAI/5zY533mLbJKwlmyGwpKiXKRoPi8QZ
VOlFFziWz2nusHOmQWE2Jq7DWhb/ve/r2ULFCxaSX5UZIFGOsnjoB/0UXfsMCx2O
PyC6/DxjB+cgwvys/vukGX7Dq5YqYs3gcAlvQ1AhZcEdh1h8RDzYNOnBOa5v0lVp
Va5jEnGQgAvHSS8zCEwvvVcaXsbopsdoYAXc4X7YFoGZIFw40RiqeojgmMYlg3Bz
21FIHMO6OUyVm5mCcnN9aEgPuEX3DAgEkUiyb5lNJ6o9VZ79H+0TfltUvitkCgtQ
xQFUezfO2zjrMXspHCcmMEO7tmuL3uXr4B8dMa6KQEaz6pmo56FZg3YTiP4xGVqU
H6yaTosRA086xbHEnk3kqkr+SQyM0WYxzXPXHZgmby0AEO86+EHhR13cjyDJW9qf
m+7Z5cVO+Wd1/yi1qet62brDPognK2ZBTLl7pMEhoyD+lF7DTrV/dHq3D30q76HN
BmEL8BjKFipL1q7cicgT274s4sJgS84LhSrUTM32O8TkY5KcCpXXVRW/pKu8EiLL
fy15eE12mzgvpMBDs4VcZH+b3fCGPVws46cgXlEY17SWDUCON73ebAf3BObev6OY
tUYOT0e1Ls2nGmgfd5ZpbJoOnxd0SCSJsbp2HQwFxV3uM943Ug4dJ4g9C4SKsHQo
Gu91PVn6AM2lUm2XqjBFoE/Ita1A53boxa/qWwVD8isiFTuD1M81MZFUkrg2I+uB
ihhSJYkNSz59vM2Mmp9R4l8Abe2ss/p1yVUoF4uLhAIo8r85JbKzRWd8XrJRMU9B
v5F6z8lVYCqdg844lxaRhTq/qsrqdMOzyD35UAHin4FTb2xjTtR6Dept/IDalvf/
iJ0lhZZ7Q63HxwE+Lzl38Fhp310TK6ZAhtMVeGkA1wmttEvxy5TFOTp1b9+pmaGa
OvN8M5Egq2aWG5Z3sG/BnrUC6IK1owS0E1Ps+Lxdj3YYcT4uLPJDsDw0Jl9k77Cm
9HEkizzOnlBrxxGwUFCF9w4IOnuDd7+ONKtwF2HM3vr3yAPGUhn7MtnUQtfnPfvY
iq7lifXH5btjQzaJaUadJ9l7r16Xa9r3iSp+IigDfEfEbdI5Jg5UJL3xGEB/k3pK
QOOF2mznKYpWU5SZ64b688fUDkRmF8GlKc7qsCJUiV1BxSIQ0btdzmjIUqhwp1Jx
UMiTo1ElZ6hwL26E1A2QB9n9SOW+HTayBHX1RduAV5or0m1jt2rWdFEqnOtz1yg9
FxnWqzOKrJHSBMqeYplZoF7Vmlkdu1AGMvCFSyThmRSSOvGrLh9kwem6J6audvXM
Q3x8gw6t7eaQynAICeH/aNZ+wy8HvmoT7fNp9ZefdI1xivEItRAL5YJJDUqtLeYK
olpFRL0exoCt0s7BFWRlMD0itcAqpfBTTf2M0LvkowxyCiXwruk4kQgb3/1+HGLC
7iSnA1X2g8GB+q14fSBM/oPU53IaxuieiQXfWpuR9eLBYb17RZtd8SqAE9Ked4Tm
HjGvxgSzEvb92sAwHjloliY/+7SSqy4UV1cYbttWXlnoUlzmmznuNx7Kf9nJy8Ul
eebQTybvxrm/92jQUQQD8tPycZ2NQlpyUVP3aJPFD/wKQZ9nQvNWbs2u1O+ngk4D
JVNYljIzSR+EHPZb7ihCJ5K02J7oZ9PhS/wigP/4vw9DwNsTXk/CmdyERT5H4Y3Y
StKXrE5zkMYs5zFtT2Tfqw0d4EiTxmRtg04vDVyA53YoMFexwxeC7faVPHjp+I/q
rzJLkoJNK5okjPQS0LsHq1m/oPyzd9gbog9s+YqVuUkX+j5/92AIwCV5Nh8Z0GPA
Ng16cJ6agXB43IPkwW9T0YBg7fJH5mAhhvaeAKLn8Wj5f9eg9Sg7XpCJxio/lgxy
cANWk/UktTJuWMZMH9shqd54AMDmeyap+qPFcbu/YZggiIYtPRdaIc11iErFhLIg
exlWEMPA9hjfD3f/gpVjhP7eCCaa5560p0nzRxxfMtT+pSzczAKCHavCZ/ck12R5
z43QKQYv2sGbESm0EXYEgAWgUduSfX8fv+CqlzCfiHQN5MCPyrGBKSHe2wHI2nw0
dNMaKPuE3FA5YMvjmAZ2Lqep1IaFX0BFpcKsnn60gPPZlVD74j9FN5HkLyVKnqBm
nXxDgR3OH0mfCAsap+u1+EKDflyfjtNpKJTncFiFyR6NXENsBHfipcHILqKiV7XE
t6YtO9nWajP0SM6Z0OLZxfTlbrkAa8Wij8zFbKPkBTqxvlGqCVdLWjZU1/SMNsBf
u0FFw+fBo6mQFIArtQSMsulfzlvcLHrnhi6mePi4V9s9wpF+x4uQSyVi4fNdOlIo
`pragma protect end_protected
