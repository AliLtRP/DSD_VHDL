// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:33:01 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
HyTtWhQ/hZPw+jIDRtIfCyv/xE/rYuq4sp+NerN+YZBxTc4jdlwzh2tvQBkBEPYI
4HocJGSl5j8lYk2iJk3Y6qN3vu49a1qu+ZvxMo+LJd7CNS3eVqRl/zx1CZeDl7oL
NQL2kaZ94Gk/xRISXvAZW1/HMOokgIAhctnWh3bSXEk=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 18320)
0zkKJq93v7W0M5xIbKEs3AJBXOleDwC3kuRhUuoKXXYbO1PKElx24HfaoHWtZ1bj
8PT03Ko1Az5drPSIugqQ+KcP2cB829veZXx9ZHGorR45CaLR64Gf8/8RDeKKdVim
5dEqeULQ/q+Fmu3k9ZaJTOfgbtFkFWLwX7WaGMl+UnFCIU5knBpXJMnVhNiGK6Hx
W+5YXdUy0lApJqaEu96Cnq2N/EKkrX5Tjmx+nO0bLk/7P3UwPCpgL4YGtyVV1Z09
KahB9PfrYKPpfUULpXLlFgrWAdQ6kbIGSrjDbL4PemuA0V8ps/hPz6kc06oZypP/
cjf4FfpKMFYUotykUtORxMHfpcatrJhtRBlkETJPOasabFfMvFRakKZ6oyFZKECf
aAydByKldeJZvyjjLAiGXD+a6/kVGTzdaQtC0sVG27a04Ecd6MKnwTWbQYKorFR6
jjKvrijFwHuO+HVTrlzajaqrcsmZc2rUOGwBWeMcWlGDZ7N/Ncwgdf0CX6VSnCYJ
2JbWL9ubXma9P7//H2W2hLDw9FjEIcgwbPm7D8ifqiw5lnPcsQ/zYZh3xS/mplf4
ypk5WzIanZwFKlMEjne6uPwUSs5EBzdk2UhO6T+4Ug33YVOyEzOzi0VgwUMshc7u
mzQBPy2CjyXk4NXajn9xPr/Z7FSkC3zxtk471PqOhe5Sop8SAClTLplOxNnCEKUF
1WAVTZeK1wZb8VXi/jQtpluW2G3zM/MKKb9/QYaJmXufao6164/dGjyI+k3Rwjmy
sI9IHTOCb2YzwfTqN8GH540gw776ynsoucHH9+/mcTwqzeB1KDjIhMSJIzUcJ7q7
9aVaGICrmmqCj0BI4iWh28GxmDeWofZ/i+nFkEdEyWZ1EuRkoKtugxkMTMCSc6NJ
yk0J0L9Nb64g25u1l+ztaaspbeX0eZ9H+AljMfGpEXwAPzUaGUmKzd/ffcKKC2rc
ipDwgcE3OpxN1ff7vM8x6NIaz5mZi2WMiJ1jQs1Cr8VOgHmTVKWWnGbxe6RRulAu
QWQOhI2Q2Xl33fuuHvw9H50oWxg0LL+8PoAgN2O2M/SW4bPLigdpwuE9Gn1HigP6
K4geeuZ5wpqNOB8P3fZFxn3QO5Do01u9WC6VMVaxXmWAOATWIlZ3YLXWODVVNnP3
xK59x8A3QCtlh5e+Zz4a+8EIe9nkVh+GyKAvDSU+fo9w01hwrXNUFzMRWtL2stmH
0N3PjJeJ/GrR9z9mQC6HqZJrIZaoU47wXPD73JtmoBe9Wp7+wux8WKUHjHhhfcYR
ocAFy/AtqaOOjbJmHUE3gX3YWG7VLt5WSCRtaaAZryWjPro1Hmxz9HyqGHJpKxd+
kIk3NXfqD/ziJZALpXHJKm/QSpJYwllcfR3+f3tNpyOmQikBz+heqVzpJnfBP8WI
32epnAHQKlGPeJ3y7jlFt6eltqJ/zfzbpW1JcYohd8nWdjIaVGpBVkbRMQm2wKM0
DKiX5ngJC1Y6GtALlvYby5bsiZEhWRrctpGEAG772zJsuHKssMg1uCfTUqZ0o04Y
hrg68hbIqBkAFuvNc/FhMZHUcw7iP0iTQD5ve7or88im8uVdLae7XXwaua9foTzi
JDmfRTt8ETH+ctfNYO9vCSi2srvZC7s1b++NTxipU1owiFvgub7uEcjTuRz3IhbJ
/otcHkjx2HFZt/+x75fSfXMYCgIkANOFK9ksPBIcCgZ2OSuVNBoiDiyiEzLBdcbH
T1hrc0xpCyWEPq/6U7zSL4j0vbfIiUZWnumeF1GCyc3jVpW6YpmbQ8vMqrfhOAfU
Sv1bzAOrp71HsLpeBtFtWIYxD/yvjHPMbocUhtAVpsSGVWwauS1rYq2Dp7mXVevr
r8vzH21k1+V/hjE+t8HY1J5yYQovXOrpVZRQutlufH3chV90t0N7jntb9QxVzyq9
sxoXwaxt6zlBX5IZhoHaJaB7NLinP9CwWsHN9okTspx/3l1+ICDm3cEau/e4v1gj
8er7q9L8UihAeDkRbbAGs7RPVfM0omqIZUHvUFFbUsMUSwQC5q0QLHEUb/GDedzA
Kr10SY8IkmNixiYCdf/I26bhPtIbk5E1K9ypcMYjYRPQEZuPrdppL2jBenZ5P6/N
wFEmRrsYVnaT6I5vvjSHzN86PymYoXeAX7ZPpw8hCT6mQ7SxBmipMHaCvFpYkmjA
3rG3McSA1LSez8/fZSQe1eQXmVFKly1718ILt9rL1ujaRqAP/3kLEsZgm2f8OreT
ms+Ihyq1m5KUZ3SHD9OKMm3hDuTKYW3xGAkAHrut69ymdTspJZnNE1TohtYTQB9S
YnOSK3M06LU4tw8mfOUtNXu9nei3pKd1jKcEgzJPmrYbjwI/8suszd7MG7VefM8x
WtXpgzHZ3mxKQctPAeRIg3dhCfDB3dD8PSO+JunFQ0DHihNDTAKU4HkI3uOOgXkI
mwSkJ3lxG8S7Dhx8ovUDrKYEkcm7SjSOX6d+lQjNojPvu4eBlLLMV3/ORjV35drc
kGvPWpySsd7y4TVUyMZL/fLf6dsARcki6Ogcma6fvWiVT4xwj6HzFyZhvvQKgFF8
sXe4Wbo7lSzrawzqlzQAC5A9ttYL/jcEtonSoiJAR9pnTMNcyQWF6e3p63Ut7Nhv
BEKTB4h3nyef+qeo4Ek1DphTZrGzRFmKTWGQ/MuAEmAbjJ6dLKgq88CtfZTF3pg5
52+dqY4Pxs30PkSpj6cDSYxEhOtBMgqwFF4heC7iQCUsXxVwKitMuCaLYnUToRgQ
cNe8v+g8o9qOutkzic6u/xu7YKvyFgdazE5ptI/15VtMuwLExHJSCliMB+TResR0
rM/8Wmm7DTUYOJ3Qoh4jwlMzQOgcCQUlXIB1k1s+wrfeCKzVh976ZN2Gk6RLdy1V
H9CRudrJvlGwFYB0IScRojrYlFsUQlmZ76Z9TzdloFo9Kq9N9NmVUjNKaC412KOi
pWEiKrkg09/njjZd56gq6JjeQD0zjopCLJrHMIVLceMZCrFE6CVtRrRr8G+kdXij
IQlvpUcQS5UdPDgQYyDatC/OgHJthbQDxVXvey6TmkHgzH7G+kG21E7ZFnR4s2JF
W+RiMl5iAVxTpHiZQVksMM0hlvwj5tBB0V6/nmrlRr5k4TnVseqSjdfNpfRyrO7N
6iqo9j9/KCsiIhYSNWl9lfKXWFpZ/2Q5FNUpUvpGkK122sxfzqatU2l/mL8xKtXZ
XobvysKbHHjXQ0BOd9XXGE7oO98XLbzZnx8zMziZjNx2Wy2smbqYVa8MWG0Zqcfi
hfoV6Lp+uzGO8f+CNtIxptLjpHNcoFbIrpjFpWVylS6DxaPB1qMC3q67NzxDBeqk
elyaZof5PUwy78q8DbUgLxSwqEcK1mSUVxz98MOCQEBnnwln1ayMhQGImc0R4eNJ
r0LBmOylDPwBsRlYy56+tnC7/0kFRFTUwaVgeeBWAO01Nr23sFeR/23eDLIX9oiN
it4M5/4pohmfQpYbexVVv+M6m5vVSjCwkQyP6Ag6KB1fZRCRXA2QSRc38MD5GPSS
ziBLFC/uIFClm184ZRjyFovVExhfO0PlCVu/+k8xX2M4K7P7H06GwsA/C71449dx
woApEozDki6xe5tfdccMVKZKiWdmi46WQ5rA0Y13vsON92wS8/QTG5rjUqEhaNgN
3QKI+0OWry4jEgXksa7aGZYfhtasnyFL+Y+lipaxxqGkxTi5fRiH3vGpzfUwRdqh
SdcAtDM19gkcwo29qjyqtAFwZkBsfPh1k/jfRqipgjPWRVfSnvfXfp4pAQVqCQKe
FShu5giTTDpKMX3lKvHktwS560lWjJxdEQrs80DGPtSj8DQzCVkr+f9qZoPyZ8xK
1KeX8eLPmdn3IjrWPyzF+TE7TTonBTAaVMPik2ezLu3Ql1JnQ+rgbosYXpK0cz72
YBmDvtgVuPpd0vg0uHiHid0lOgSCLCfbnLLaxExgrfYDEHO3fpwEHmfGi+P/6dJC
RBuRZvjkib76lxrvoK89EbB8h11k8CSXOIkahwbCNFoteIyxwjwxid7fjXznyQja
Hm7NbtDlKO+asxT+Nh2CtvXomLOyqt1/BVV72BoBy70PZJMg50oNyiFkxtl4NuTj
OnvzSJJ+MRjQDYh13q9vQur1R/BTNt0+JNnHAbRKPl4k0/JAbKAqpM0Z2qedc8m7
abmoskCm01q29JxI2DlK3TqHEPCihlRyI+T2kJrSq1d9SRJEnSEms96+iljcqu6Q
/GfYiJnLdkiI01A4vuJGgBYODa7DW6i0XXQCHwV/1YdUQCdiI7buh5USEZE59jAO
RT2jYErxoq6cooq43pVosgilAYw6T3akyVKZOiNFTldaT1WzQ8VeZXGGJZK6VIkg
5l8Vakj9cA8q5GIS7mDlVPj2v3lW7UQy5ln9KVUH8moabweKGGorNsHjTGQEK+tl
B825krP43YP5vlSG1ZXatP/lt2kib4RKVy4urJHA2s3WzYIF1wCQJLfMlsgTsz9N
bVgNTApNMBOXXkCT6XijeLiAh29vfllINT9w8RdvDadd63yyz9WUAdxI/ysqDXGH
+hSndOK363bijdwrOdy0iIJ7M7qFQeVas632eAt66w/f0yNZi5H+uvv69wa18zIS
gu4DtxY8+h6/6KI2UbZSZq+D92aHx0S1e50JCRSkkZJGtD2VeGuiZVPR9EwdRkVV
3UgjJxKukTdagYVqErxZxuYcbGKxqlOKxRhZaLX5I9sQCQHMbI7ofMhKOb7e343o
LRTYNK5F6k2GI+A5Er9yTto4kwRZDXhQfJ4+TtOfK38iI1mOGh6FU/SGdW+Kyxk6
4mXSv3WYoMwCfWSb/zYK8G+KH7OkfT7JmAa17X2x1OnGwf8/c2GOxlsIp/MhI95i
7BqeK2VdNEpCnDk31unt3GtTL8SNxKaOepGoWeL6QjzF0g2MILvgemvizr3b+5rF
0nVLU3OdKnfUHERm8cIHuHrKhIvpDrq/aHQjZkS4jSgywZNNK2fSYuDCAfhCARf5
Rag5ePKweWg9EFWGdm8mj0B9AO1Qob4EgHRcITnbPE8eUEUBRi115bNS+QU3xS/3
OFrMFVyA1fZnHVvGIDOBNQ0yVeNeZjaUHjWwO0CxHcP/AZe9o6rDL1vnR4dEeSx3
44sZ0WB5RqSiTqo3iKYyP4i7RkkiNtJk7o5+6sUQ7yKe14WK5mpeNBZnsGEGHUc/
1mgmZt6nh02/q5jT+3ZUXUtIw8GbbdomG2Sen1IZUu0jLbMJTwBtkwVU4Bg9RMSS
wNE2DojT+enjoGLHiiIdbpkLB5Ig3Zw8GW4cRu6CB+F4i7h7sSPZM3XM3X9jVQZh
KIKP/Dds+RUugruhX+Y3GFF5xgnCNzFhtdcpuA0BB6gtXzQI40g5QA33vVQ3w+3O
UrkVa2bkBjptXMPdwE8MBkJ+F1MNHszFmjKnv/TVvrnTliCsZ1HdnzMaEk5iK/Eg
03dcd/MLNZZXQeLqyH+gDiCvuaXvTO4yI96EtiIkd31zJv60xf6qvoCufV16fxjf
LK2o6VXVTUL8LCzlzg/OpW5rLHbAOElCJWQSex4vmA/UhQ8Yd9I1nSumLQ8Pa2nx
um/Rche2LFtOeOHp2Lb4DxsZcPrwy/QA1tnF4AABrZKRVDxrFZGGAaFMWl9svEJI
ro3WBnRr5c5rBr8YCY6LXtcXddgjJOEQYn5k5WV+gF1TM0ZgKPVhSg/IaGRk1roy
cbd40AdLf3UNuwiKKvRwo9b6RGD19CKTaNogpPaBjk6w1ZiQ7jymo2WrpQYvvy74
z3Ryi66JlEDoJfNGgfSPXLwRV8YD/11ku+fjVKufI27aXFK/vbFDDCDlaW08ARC3
a2c53pc7CBgL7emYfCD1GE8xtZYJmAHgIa4jV1GNGBe3lK3PU7EpwUdgLgu8xaXX
fUqvHyqR0FcQb6BqbueC/rEPljxtSAKVOwas0zeIp/XVzlArlTB4CMv5GIY5+NsH
XW1C14VLEPl8fUtV6ut4vmC39/EK0IpQ2hJK6qXSNpJNSijuqcmEnlyVYjw1NBZp
EmQr5is8epzRnMFNq5DiKemhz8zj0wZBXgWHgEsXk2CSM/pK2fAddeTxUTAwswO5
J/BFMTC52MXUBOFN1ouQJ+LJN3EGI6PS3sVPbVu/1QsyLhwvNiY2pWTPm8lYjXLb
Pvl8EQGEySMfGMdG+OVZr72OBR/HH7c/hmvXyL2pb7paq1ZNClpXdsDEN0fezg1z
5CQbwK0ELvTIdCkxRuVTwtYxcDfOQtp/H+bVKQx6ER2h9DGgA49ITTEGd23cxP7/
i4SvMDF9kSpKyTJykn918NyK+3jhf2Z7S83I2cAW2tFAon5m+VOgQTgpv4CjqjwS
lJvGwFENFV5kMzCme8zV3hhah180XdebMgjuJgqB0O76NM6w3cgqmQGOEZHV+vBe
PbjCXMS8nRHTFY6lGYr4sMw9qAW11z1Dd4+DVRKGOJhn79a0Hd8q/im9XoY1FImH
GzR+EUv1lB16Td3qyM6Z9LhQ5/N2akjb6P0BIevL14JXjpCzdklJlgCidEtr8VxF
W9M5Nth3LpAQGUyhREbNCk0c/fE7DcL3UKn5llzD7UxZPq0ZqPX/vsK8sTWDjj49
GFFq2SfZPu5eEURYcHls0Hy7MK/cg6ZeaoaIcvuyxqbSAzx32cilSAvws1Iug5tu
eMeIZb+L17G+cPsE7gxyN/IjWAXEokUZLS/f27FRK51GV+hEVXnPxnxS87EfzGvB
ZjYmZlG/blAHqZaDQFlsi0mEzxqPZmHiQOGSpKU4bOz7pGz1CHWfB0bmz3HNPOwC
O5G6Y5k3LOcC2R+PrStVpWfzNq0zlqmqqn8vjaww5O4nnxXJhPQbOsX6bhc4/7LI
inegfHgbveFkUqX+2fMsfh5M/ivhN7OhjivcUulC4zfYdmQuNR9fqKknK0+Oj/Qt
RKNM9qROvQwyWkAi7MNOPCkuC80ba960Wp8I0xPu83T4V4eSYm5aOXPyKG+Wj8ed
jaR5C+AYhn7RDtyjXN2W+h/9ycOrMavHo/s04kNYIG3Q8KJk4jSnRv0m08sH9zQq
PhNBOyOuLDx5M0v0quAWECvEboFegkpwiiy+lmF8Uqb4XC3wB3OnttSJnJbRp/Zv
HlYoEfuiGxfq21d/HRIq5CW1xpSOmWIsa1UM/MLkkd8u29NJzG0TFJIdxkfegFSA
KDfrtkQAH55/YTvTKnEbd5CKZsVsJqHIS8wOQ6VnS58dNJYdtOTxVg9lga7BaB0K
X8hjPBQfptWjSLOqm7kqk2lm/3lark1ZiDo5ARjMbiwxbI8wJHkGxRo99E/CTfon
VkNYYANvnCR32r1PlVfvOJocUuRgKQuTzLr3IYY4kQprnAWAIhh+W7NrQa7Y58VX
g6hvbgPD7KgqG1Xl1hOaVjHt4m3qAj5ihvZH6g7X1t12dxUUKLpI2+0fsg+GSqEG
8Y/jap5xI93tAW/Tv9yKb5jhOkOt5HZN0hRkvuUrypD2tYV1meIklObP6ttQyZhv
ozb050WD11lzDyyafQZ8fksED0dgIwlmKpNQIaN/4mb0lkaZb1lZwxVLe8/9Y0oX
LjY9DOaS4nVOz3HEKwuEiOUdcH2JfecuHMuVgl0f6JKjnyWwS0mSgUuwC4XUN0ev
WXCdeZiHk2p/G7PRh7GjvUad+B88jzpBWDtU+TaIZUuYOaVeb7kswJkxOkoy2b21
1iN5AIuLhx7eOSzfkUoCVvwybgi+A11vrcrbeGZehj/lbGeQXCK0nCDT669iC1P6
W2Ck0cgRY9CloHkfHyPEZDYtZ7hnEj/2bHv6UeXsgiSpcbDdTqsm7VbEX9pYZVwM
yvNVEjXwNYqr+xdygGT/WcEBjQgMAva514EltSUNYpOGeFFI2l5+j8pcQ8djoDUS
dahMnEQPEEznLMYlG4/bhaH9SlyeWf8LT09mkS0EYrRU4xKiNgo4OnqVewzDHhLY
WRORug15dYLRjGSyPeu88q/MhzhzRtkdxDgkeMCLHZtqv7N3M40s/Zs1pEUVOGAK
uOZP+w+aMATX08KoQZP8jflSy40e/hSGZEPKWlIYF07o85BV5QJUZYvpkkKqMZ2N
eQ90jtRw5BNVQPat7CNfcmuH3N74hNAjnWJ+NyEVmzv4UdmdskKdOUhFpSwwggPJ
zZ5cNNLgMiayBxKUHVb81SPUdFVZiXqIuQGNWuZLufrCFrJT5wMvyEMAscAKeRTE
7rOc5PpSYKUCZ8N6poG/xsa+u7b9LDhkmAuITx+TlMExWa/6lBZ/zxzL5sLTmD9K
2owrIC0ja0OCKtEpQVkgGv1kOf7IR3yYh+FKRwGCv1HXZaBQjtkG7VLad7C2EyQb
lmAemlgMJ+hegeOrz1rALE7Wn404c0Bkb0lZ8yLUTGljvHOKkjj7qqvYIeiM+AZP
91rwbFMN/u4gMhpbGdtgSUMHT+mHvrLWGu1GDuA7BltL8RCi13TqdbpbBbhPNlsV
1eW99p7Nt0oEDkWAndudHAIyBkMFAexQh63FG59f8Cxadzn8zmJsqU0z0pDdaP63
dTr77sMqvBpSw4rZnG2iVSzTfAKTj4srot4lLRlMAps1H5uK+ufz2KGgdFBm4eRN
X18Aj9p8Ksq1BZZ29lr9gsbnytyiuvMY2TZQY0NdrASTWA+na+oTyR77GMZBBw3A
uVFcZIfpH6bmwQE/uPenmHX8st4AJWBDd9jppjoOodeNv4fyQFl7yAWld7Ql8NDw
41w9jD/1J1I1sOt/0Y/A+RapimPb5kixfUzNg5IWF6er85rkNigL1W1JxlpGPA8p
MMlKivCY64mjw5Cy06ufVAwmZkmb6xp3ce/ti734/n9ylTjhIYJzm3JeN+vasBAT
zIbb7Mm2Llqs3u4+oeaQ7mtUvpehpx3vT3fZcPbGqe1eXAaNdnk3nLGlLpGAvfkG
Tt6+iRzmaXFKGC9AaleQwXwiXCcF3f6B2HNWRxxyU4N3B9rEEIIsL22KK/6Aeoap
UiV1oZlW/7QHCYFoyTgW6IUXWtOP+DapxyAFi/OuFsLA0dKhN0zveFQSuQAR/1yz
o2U1mefnReI+q8gvmboVNMnhQYuTpTP9/8XK/j8ltHCIkg3+Mcr7ZEoPIKkgW9ML
eymYYVq1JhNxcbGf0tEfPc3eIyDa63NKXqkenDXJa0bKXC6DmNYtASQf8XGIrcdp
r+9Rtp5P65dXgBiz/5Q6zjl1ggQXRPs4zaY7Et+D0Mv4zbFpgQ0x7AMFH9mKhNjF
p7XG/TwgwqJ4z8z7A33mo7v+hnd6Dn74Ji/2KquP5TuPI4Bzm3MkIyTAkhFAQ70p
nnBVKyWOKf94QHiVq86raDqdm/qolgXq1ku68oyq8J0ASNYqdrsuRjs2jQSqEYup
tHnw8/f+ZLmUlzBoFb1LS94nGbkKggvTHJf3dDzk61T69sWfcbwmJZ+bKJJ8fwjN
HI/fnme0BY2NBpLnO24j0qMXAGoF3y485kORqFYbPqUdjQjNna+FVcFqGbNVlhIZ
y5/4Etc7IHF/29/PYOHR75n2Zx+x//WN1+46dCMg3tuismnLl+ItVjBiISmg6md4
i0RI5zXcK/Nvjg5jug7uk0GzPvynbDFRNdv7IQcBPRjtw+MEmqOPDzpe4IqdeWVW
KOeBvXLHYOAxiDGA1NfIxaK/C8QDR23AqYnraqhVXtjz4o0OcJEPbk3zs/SXJjfb
5wF61DW7/vNzVd55XSeXEzjr9OMnDKz+Nklb+UA1cbiWGyWXjEib15gJkLfJRBwZ
VC6z4vimyAWDc4kGH+o33AxuUw/cVsA0pmDXxoNrcfBWfWI+T3UYpuKVzK1qMRS+
pfIoPesfSj8wEa+tw3kzcQ+CN49TluVbJlixKvTf1q7RG+in34qlNXcXcfQpMpKP
ym9sad8m7CcSmm5jN+qFpkt0L3mTzsrBsx6llqqeT/GqB7Tp9b+x2biE4ZC7Dg/G
QC34Mt92IJrcRk3ytOCdzy5vJQXgV4zjp1JQqR0s3U6j2ZopIIMRT15KCtt3DdaO
wxto3h0b5mgTIOg8Gj/5+/GR697kuo5OiU6Q8iEoKp0e7zOZkV0RdeljSRfyLlv0
in8YyBDRSNkWJLJcp1KqnFsoSjrF4gZmlImOzuN8W8g8FTUHkHOxiV92qRtzuk2U
3onr8tCtdF/mz+jOzrFhs9YRUQuUn7dkRGv0oxvCLeXEOFxuwQQt2PvDAgdBVW2X
JV5/bFVcJz6h+CnX5Oq1nxOin3kXIY3n3Kwl11BGpRKFxLwAYMmYeOkJE4lJ9TIe
MFhNaD5LSeeuyVISBEHB05Gjnhi7bGNGb9Ok13rAA+HqfQijZt+Q6drJGsY0hApo
VcxdNMxeV/Ml4KneuztiGxbflgjpuQLlT4s6hYRus+AiYB0Fc7uAoFbCtwUhzfGP
Drhxab8y9L/VGYNsXx3BQ8b4I6JSvhc0VJ2p3qnVuHFtNJ5M4fAXPpydi1zYblTb
1vcHm1I4MP9w70VL6Zngr70SgoX9SpjZMAlVzDiB3r8lsi3UrIailOdVcEs5ICjf
W9NZPtcfb7GkbvTtySdQOGqG1f6NfwICVfhBIfQRa+D5k8cZ/zIRNoPQxU9DdnRS
tsxMi+4x3uJRzLPVsTnrIjGbrSNyeLXtHoMOjYzoPyVd2X/KOcimzL0D8bznkLkw
gngI7wYNzbsbcNf+p1LHwLT66P3EciBq/tTaaE2luE3f04Vk53ABdhiductByO/y
WCFVbDn+zqao9h3Ij9Nx6VJolomdeDlbr0Vkbdh8eA50KelHs2MT9uTNN3uojZK4
618oFPKyZhqmjfs/OxahW/K5UkCCWVUwv6C9U69qOIWaFiHMRw0bFjwFhXIqcV7H
qSndcnhFmBrGPhYcZFPVZdtuf9wsQEXFOeBmWYNF0Zam1x9AJVrcKmVlE3Hfnv0S
T0M7AZW9wjycF2rpguzU7zfocixzfTI/fWFBUP45ZAvAdIf+ZpGpUtGARVBZ070V
jkgwa7ubZ5snKGlrpW1/Vs2Pg83ae0P1ie7CS4DEAtayWS+drY8TRJQifQ3+/bUd
YQYHRKFBJZ+NO6oI9m3tSlnMsyqO7QkrQg+D3bZFxNN3WOHTMvqfxGm/Le2+s/l9
iTZneWmWsnUdgBv5hOBgEulfdKKHreFROCQ5fVDr0VtHnZM9CDvraP6cLZP6jWdB
RcPdnlCy6jhtKJUfX780h5KGDs9W+yb3yoEHqWnFF4+iYCk1CG0bAEq5Tj3biBuH
IR1M2iDLZ0NohFPGDo2pJ47lCnzTEa8oHWQqupqQPqzk5FcJwM0QxpboThxLtO3m
DDJCP4dewaXNl+6m1Vs25EfH3o/eiHLPlVnmm607ofQa3sjtE4rs4tyHp88cmAQ+
+RiOpX7DyqlOBU8nwXkDv2NWS4wRd0ehyEGBEXxNSVU/khk3V5Zqqu+/1CYvPBvc
AWeSGrwVGKOg14FZJQm4NP9AgAYEyt/IuKE/pN6OErW9z5XFcgJLYSnfxaA43Kcf
X0m22voEwV5UEIvgx7QO4FlyoctokYW/tjAIfTBVdFJCELLB1vkEw0huOv3AHVG3
v6P1Tb6JYulIncq1AYFgieHH7f/ZaaiTgLiDRonO7G02V6oIYpvgsMsP6jGkbUwN
Lfu4NaHcCZIKAChuMbJKou+LtARLwndKJu5NDHI4OiCxUedy4BXoqZ39B0+99l9q
RidcMrF8IGMvkBweAewKlj7dzbISdkD7W5hd5OQeNN8u6xk50t9wyooSnRghAb2j
YqOaD/VXan4FWjquGzffSkErr82QCvlOYC7PaAWdXh3RTPGAc5U8Hfent/c52AFG
HoZQbuUay7WSyYn8RBTI9xs8M4T3STEeLxTodFg7eOguXWKbIou78TsXXc1vHE4+
2ZW/XxuZGJ/WvJ0GdS2iHdyz/BzVqmAcejq2xAXPdgCvStV5T5h14Lnpa2wODsbE
cTxtAgom3nS8lH+i8qacOJ1qZPJw0uKVhyDQyvmE4RljITAOnYMfry091CxUKQs8
71cP0fjw1J9+a6PFMmnEO1tR0tHeJRXbmq8VlBLXm2kZ4l+isXPteQtKdFe5/LK0
4nKlJcyMnXem+xe2vbuhACY6xR+8emogMvhM7IuAW+MxFYsMtB9Dbkah25V3agPB
foDzkcmT5hzM1OFVGoHDLlJFsnxGnsm21VGBnFDEpBRhaWOz8BhMDfpPCMXtavr0
OUFQ5e8miWDxUbY+EKR5GugJ8QthbQPzQsGG/xKg9vMW45iJOdC26fPo9eRdicLm
leiHL5qsPEniSXhWicwHbGf3Qx6iyr2iFXDagEQFhSFI9npyqnmkw+huUnXLtJNg
k4X3g5KDZfSn4/DYyA8XWKnuWF559XU9rNe+k/IVi/LAFbprBjsw4AwPIeLI7cq6
Sz3hKnkkq56D2BM55Vl+FYYpa2hvipdj7+DbXj1LMyck+uYVgvdREeIrGCwH+uGk
aJl/8KYFPMDJFK7fxSxrf7ghQ6kJgva4Y39VU47Gq9TYLC/d5d7jVQwL7r4yQtRI
/TDm8j1CgLVZ5dSXQrLGoU+tZ0pn/cJR5ARfC8Ps3yNYQZn33RRWkqazyd2XZXoh
qmPg7s4hGcbW1yYS8lvPaEBBH8a0FguRquS5h8USpnzrOeSdRyIC5kNALliz4sED
KTIOM9Aik4kqxHDmv+XCs7PYin7NpThBpGAJlqCRKrVFPkkOURWuJgUidZSDAKhj
xFGtEhtEli9kM0t+V1JLjiEt2LXkoqEXneMbx4uRg+v2VYoMkp8uFSxuwQkQBafQ
LBo4IR0VFGAO+NPJrd8/70LAsMW7i493l/naOGrAx+SN9jjG9xx49M0PzzoeHcHX
miPe3wRtRVBfD08gI0HpawHorcZbxOViUmWAuOiyfIpuY77keoWl6udydm6xe96M
eRNzqfoE9EpxTGfs6mgGdDEru7bsOQTU7NFEGAZDqWA/DkNJ/IsRQUrwmkA0GvfY
QzTEGvXnue9bZfv8uw/+1FZ+TzwvhtgQ0dQV+JGktq7ydPfLqqQWZhg4iRSU6AkI
Hc2GX/kwmdLDHiDveUZucr0Cj7htZeBShYTI3SpZkFIavbbRZnkOCY9zMzhPy8W3
4Ji4XokO4qrLYGfPb55tZmceCkh0gQYgVm5HbF9lZ93spzG0ymGja9qxJrzPBLuI
C0e8Qq/SIV355iQ4O/kCljlKpLIpTL6Zm2ua1YB+oea55Uym+FDJjl4Dgy8NxfLu
gWg4W3SrMG1X7Zvx/uK3u8K/w4QkE79mUI1nMsHwOHp6g5UjV9mW4HOLlepr49s6
oOOXdfE/A3vQ2tc544LS76Ah7ICzs92AoFsKutR/JKuEdLWRbmqMdYjob+3xpWYq
i4Kl1/L1piPv+ejEOkybk0EZq+BtQ5V+FLzeIJ8KkUd2JnUfPR/pA/0PR2xE6IHD
AY12Xj456lZpjzPQh0JYZGUaaqWVM3z8OauPDO/mUERAzUe6TtZaZMEkKk0TvX5g
TWC8rs5tyIH1fH3pbPayN1nKRAM7WxBiLkLH9FJs5kDIjoaVLrXrrqdfueIq5uQk
3uUbW1zD/jlQMTZl1frIsas4Y5qbFBtBvA8BLkEmMG0p9nM/yLXM7HRjQyA806gy
L2XJTd8SPGq9cE+Zd0i+Zn1n/tCU0f7bpguGk3u36Narj7rdf+o80OzfE8icDEAi
/BCwjS/Ik6uSMOTuSl4CsEXmT114QUCKdBcAZStqZ6tf4awAlNXAk0LEyHZH6HkF
3NOFqnPhkaNDd/N2NR661qoxrwOfCmJIXyKpHNVuqDQDPkCQR9vfgRpaEis2GWjM
Az6ftn3wtXCVQ3XTlE3/EDdzTVuQ8VkdyORmQTw1Q5uwR6iqxrBS0OMFIphFpG2k
5fP1Mzk/4YkVdxRGStz3NefSUMJDKWIrlBUL7SJTgsLdRDEeP3VUR/Ev2nLdMI50
GWT2gmlxiQqlQuViz5D8ezOeBdm1fATpZeCWWzXkL+YP3HicFeMRfeE7YgCjuMa0
YwHnm8J8GLIvm75niVS8TIadL/O65t93JMfiUrPxEKgfKTVHeHeR0JJ9zwHfu6ge
QYuy0KjVAeU9sC5ib0RN7N8AdBO8wejxYLiezbturGpQHihxcSMwXABkdNp1Mkhq
LGYQEFyRCqO84UHdhGNfbVVqoSeRUTqkUIj8umt8rKjJIvBP/5D/6CXB5C4c96W5
K7fH4hjaff4TkvjdwCufNkdH0CmtvdrZMBytnEQbMAlGcLQdlZ0agbOQaH5hBevI
ZqEAtWzlAoIjLjp/T1NE2opstL/LKk0ZmcDkYLXfnO07mEn6VtWKTuSV6fBqgaRm
UZCRlhIEzlm+Yc2uOa9NM23lWej6WioqkwAsxzmI8pwsNVAUYMgW6HW0GGENA89b
JSzrGsiALB6h+JKetuXC5D0mh+MMl4zhL5l9ejsF4wdxxRwv060XMPedHONZPQAl
9Ed14uDXYazFUW/8RjkVDHXJlWyZ8oKbIqoGSojyl7NEZwjxZDHu1+11Fdto168v
HiuCkFfuo78JsKCpW1vxLNqfrMut2xYoOM7XN2DfF2xPzhmxdy8M8dvTVZ9NiyPE
3w2mPA08Jhu1vkS2KVWTKssDAl0hW12lGnktF4hrOjQwOLbOkCD3rSFFZwGG+or1
rkYe1BAJScyxcWBZzHiHeKR4gWop6GEKyc6I5vvYD+GlPrDo5WgnJAT+lFPfm6Oa
rt7Xxqo17iQFm3aiXD9HXYHXRqEhj6UQENU9JbtMn9/fPMmBkomoz506I8AWKf9p
+Rsu3aQkb7zzDoW17l4/1Z8cPOtzIFDOENJ9lbgHFCyoWGegMHeiSnDYO9TUzPIS
Z9KyGC51LZoMA+DW3stQLVtM5YFsjzo4d4Ig87u5LsTuPy8Yh/NgtUxC3qzglC+F
NmOMJdGi4o2sSMfHPCJus01adxb1ZBWoG6F99jcV+EtWv0NYwKk1krFoQ7hRzU8k
73SP21OQDRcxbLTwNgeQhi9R10GQivw+SdpuQgVxg/myOIwDSiTu1WaYNyRmHxQD
an3VV9LswJF77XikRXyNC8dFqHuWiftT2D6GExw9CCc0jA9cfwDB+EPCZ4b/pDDN
+BOnyckRuUcU7g7rWlE4WX0S33zh2jDIVR3VThsU5CkkSuMPhXZ0XLcyR8+BnF93
IN3wBM5WFtLqgPHlzbqQgblrvZ+Gvokfp2Twf1oXcqkXs97uOAFgsA7zx93k5AAH
Z1HKc0N1ZKwSvI+hDgooFolR/GV3EQqD79CCHVqM5rdWYDTeN3cjAIrPCUUHLH6U
OL2a+ZG7C7Ckt3cCdHUz0JKCKPxKNYozWJu6Arx2VO0KkG22hLWczidEaYENzSlr
WRm3kgOpFCv72z5cSa/tmlQJwINSMLgBwdaGe3QKp2wrZAXNWekj2/j6XGxjmHrX
o5pRz1eDa+8vU6I+zehpGo1q3J9YdX8Y+Up4ZcUGAhAdowuWT1FKhPSX8TtMJNk4
uNNFg605W39hpQTlT0YzjIDm0DYAwQYO6Fg/s1k/M7cWXId9gpDfVrGy5GdB8R/h
XiZ6nGOvjNo4bkg6lJgn4fx7exMpoqXVmC+YxiE9vObJnlgx8kB9EnVIK4c2zZJP
cyEdO528EQS6j5gL9p/z8/0f6TFMcYwqnTfxXPZ0+Ft1qjPFvzG3szdZQJ8cBbkR
BFOJLDaXFURo36vizm5Q/9tbMk52mIjshHFW7IhnNKakeYxR2QCQDGaZbAnuwQ1y
AcWIKxNa2b4KY72qRhjlIKp9cFluVLfzC8xVwkAqHUluQaQH0SveuJjOGSmYiFm7
boB45+QREImnq8L50Eh3vUvEQAUSIq5poDJAKM1tgNQ+8viUTEBdTZ1jy7QGPJQr
FqqvWQtYfP07vJTFdg24mqeQtPSBRabSirafMAlywT7j9FOK5JOxGaQQnFVXpK58
4mclrf8T8tRaJVsFeK3K/XDn1QVheMs3j5etaeNqFvrSCZFACse6e3SI7m3Z5DMS
RE/CGDe+0YNF2f9VjEw+BytjS71lb3QoXXcJ5C3iNKwO0lYUI/ONPDi1k02/z4BO
lgasWdH2LJmsxYwrFvSd05vgszF8gdvl2rtf65p5juUziIc01br7ZgMifxs0TFlX
601rKazdIVKFNZx5HSKcArQHLwxVfcSalkYI2vTA0f9MZoYq4IfoR1BWBLqACgmP
wOMvtfnehqJc077QhJwyDp8aE2mLombY5E5rOaMw7YL65ii+/VXgtdecnzv3BzB4
GcE9XbQkX821m7VwpsPXDU54AHzVlz6YnYVKI6EC01gghrZ98alEVSDjlWkAmAIO
+UqThwUUYtVSoatPvorWhgvwwlCV5Bevd0613LikwxCLF+R9OXFysjrpapSMkJN2
h8Cj1i2CY3r576Pk+qXvZLNPjZnYTPI+4EPfPZJU6rBqzg5NGct7rQ5gwUV+zEvc
Ir2aodqO+5Wby8BUjnAUUIMFeIssGRFRlDAiwxgfN71Am2LtcQzr7ri0M20eF25n
dtJWJGVktwb0R8B2R9cGYjHD7Vs8YG37QsFjBuuLg+dMQViqUqFIgSi84xDg2m6F
vXgfDM/rSkewo4sRjpqY9qGZnGxFiiG5drOM/TEv6Ke31iGBOaghvMR82J82zTby
3deO5DoJ0jNdlTiI8JJjdawu+0GSmJhgZwKD/eZhpjxM1HwDoi2RN32zMNvlfMYn
bh9Fhqdlbhb0n/wJYELOOjVBKzTAdU2pXD5DLvUbtryFf05RmiofJ5u7vqA8DLR1
pPcFK4SK3s+XQZhLWRJX528sH7Ai1SHUEfvlhbOsIuVOaX+D83L4a/YQzFlvjBV9
czdiVpYIEL5I88jKPefcI/i+fU8JMiz7BAzyTsyqea9+1Z2qNdvNV92qcq2iHI/A
UR++imiDDxRqk76dNnzODQ23ZEytcbZe3df3+wLTLsExNCa+KXZ++14sg2jnWHY2
CRgiqfchaWYDm3WpRW7xJzkltvAtONJFMjWdG3fhuKK9Qv8ywoBIfQFBEdaZY/j1
zv6iGV3sxwVGM1Zu5PlI1zshHBvKVDxi+xWJyDjxypsuV/pf39P8WeUMqrKxzrnt
gcyS6ec1LE2nornk9rIu/HBh6W6CYKo8NAki+OAoQm4h/IjQ4vLwEt0/4zptjp2V
o74INx0zAqUGnEZraagjtlOyoUfeb5UzwEwnH4E1hfLAXG/XhFhmVr58J7TLyEJp
BchKUJePUrQvH4PGSG0/YDqRgcpPFAo00xUuvfkjjsQLYpzC74LQRaJc17jwhkzP
3Y5z/SYwcyKCIQDxTLOeLWLVSKkbUiYZnx7s+fEh+7I30O0X5GSa0uTlnva42j5t
SX6vM0/w/sale337Jjcnwdv+OveGbO1bNDMJuEOMrb6xQYcYZdV+s4aURnF0IZxm
AT+vFrv8FLlCj/X9d9MoE5t7+Cxomz5ERe2GhryWASY1bqXLUS84srY/9XGqWRlw
5AMF1kuhx2SMnonOXlh8IcitoxWy0dniKBrehXxc5Ed/KzXGoBGNXS7I3lT24ZvK
hH5j4zzoLs4rHlbE/LB+WOcgCKllzyGtjT97e5zFGgMxUBevnihzirEnnCyK3k0Q
cmyhQVIsUgLg+yCuup+pFPl6+gF1jnQhf9a91gNz+sHCkGeWStPEVctp7Tgoxh/7
SADLa4TaHr56dHQbvHHQCAgtBTKfSi7UDN7ZEE6ngcKkJo/oaBnDmIDYTr1FkQ2U
bBLu6XCYo+JVr0chj6Pz103GKvJQ5hsRVrm5A6W10NwiTDETMBRum2UuMeIBGJNv
ENq9Iroq7Fjo2Hrs8zVNgZwK9MhSuR5GH0AxtHTRIgumk3p2YUOBDLVZw8iUNj+J
Jr5UmpwsiHMv63OcvKVb4PUe7yKzwDDz4LVXKkW7xQ+3lRp9pTGqYJpU/qxaVyER
pewK8k/6B17pd/BW6vNR0/kOUth9gVfOoCmsH/WLBt2WWXIIf/kNLu17G6SwsceY
lCYeOtl+SeQjjXJlDyiEmagyR+g5y01r86eOoF9OhBl8JiuiNo5HcdexGoNWKffC
du8jB0QKTAooo4B8wJC86pBtESTihgjH2gGGOOHHIYztg9Lk1f+xlDThdvcL0Y3j
rG87cSVJntAKwSjQ83uIiDBw4rqRsrKDecJ+UE0AdUWY4urBfiMuxeAjThnPtahJ
3ohcdX57hrjpEcHPAzw5kc7junmgj3h74NbKF09oCjoVug04R1ufmnAxLlcQOzpb
IO4YpjNmTgOJJCLqbPDseMyZxgFJ61WJk2tI4ujYt1u8hbQuvfbu/2OKsHM89Fp6
g6dnt3FVAeY3EqGXmJS8b0VlFd9a2jhQUlomy6aPcZ7En2pggA5q4YSd2ey8VY65
XkNezyb1ejTI7jSmzSbKLJbq+7hRpb1IyQRLoOt6nREngIYgQ1z4bNLYIWvjPwJz
E8NBK4CH96K+BSjVDBVZLKjLBexAUsRx8LojOYyA4RHsojLUhpkj/ip3enuB6P+/
kkf4cMQRnDWKR5gxv9afuOajRDY5+RYj4VgP89uzNJeG2JbDcCZcY9o6KbpDjf0h
OO0I8z4RU52fFU52YaP+3WlX4CVlQCdCAsUs9G4onxFb/s6iWmoU6RTpztow/8TA
4ZnAWkcsnRtV2snVmPWxoUZtLF2D/TIawMYR6AZRWflgNRwt+2b17GdOn9QnziTQ
d7o74VBtQg1m8XFe+HJJZe2OizfoaL7u/5GVuQNrd32uHYS5KdCq6JzMTKVoYSda
PX1Yq60hXsDFwhkXua+oKqgJq13/Hb4a9Kjx9dSRltxsWziCqWZHL1RRxw0cEN11
zy1XCeXiHxppxJ8xjf9qGWNyfuZI/D6bQBI9rA5AAN9O+u6G7NE29DufuI1cgXv4
RQAuAImvB11yWM0SBgF7W9h1R8Pg99wjy1mQeifaxArfX4WrOdX+l+YjWd6HAXiD
Nbl1rxVYub+uCZsNsKn5aOA0sfneLLbUn1JnsIAh+vyxfN3v8zK+JIyvSWXl4gau
3gbVyKISB6Igchiv4h98+khRzN8Ky4xe464/4C3XUmbGejass+pCpANK8t+8BBu2
GAhqE/UDtIZO36aFrHw5DhM+S9eHfpQSjuKF7slnNiinaEcBMHV6bhibVC9bInLV
cbWmmHYNH8p6mJpS+1F6mXUN+xrU4sXW8SslIQZzwtXy6VYZk1w8AktevVr6FLSC
TsXtrJreDp9GCKkdaCQn5LHRDbDT4L6FacWO8hmz1IJtCedHEcvwC1nugcXgocho
h0HIys4dTE5orH19tFrwvC9YxLTyF8QjrJ4kEC1zpep+WDxcDlM2ROye0u/kdhnF
vCC3PoNWo4Xptsvn4brxwQG9FuktPk48mEq9blR9klLhmhSWypuiqxAPadqRnrgz
CjBfFmRepC/sFHTg6duS3YEK4OJc9IuvK/22B+muUnM5YTRj7NS4mTB/WYeuw/Gx
N312RRMwI+m/WDfkI5JPaAo3OCQrHhbXoY5xyso+aD2zCyIRBKxsA2MxwV3kBWeV
eW3QJCY7E3f+Pxq+8gTfX7Gt+vZEC22VCdhkiwMGIRNqlvMhqQvqNiewEI2g3VEM
DbBBDdandwmDXJlb0S1jRtVUrdkYzoilK5gbgUoIJ/TmjYk4UkwSW46iO3/FWnis
fzOZOrRB6ZbqON9tAhtyJ86p0HHQfl0Xfs0flMrKEtaHr+T4ef6MdbvEJ2GX1HOU
vFgt5lNemZ/QSeZWhVK7zl+dECto38Ppw1DQGLnPGrfs9Lfpf1TArV6C7joYVuuB
SxJjXixlLsxNgs7qU/AX+YFacVY/ZqU8O7lHyQzb6CydVJpT0cgjA3C2iT3hUQug
mI/G54o8WrU15mlLvYksRP8+a0CYchlYHBfEYCarsrYjlS148M9nY0sSp3eL6EQ5
t6honOG0f9M4l1Cuc31cckLRpCdsfkEf7LoAXY3MGnhjOPWXmLTrSw8YT8jQCfFx
SpZ2NAKafM36Dgc0BthK8XPsNdiFO4WAS1mjx4qCjpiCUeHceZoDerypKM22Z27Q
BZK12tHFgB6AmScpSw2myPQIIZYgXxOcX2ALMfX+tvvZHePS/Dxihq2QqWfvN0Xt
XK2siMHTDIiOpWCZ4Wd5mSNzHq80Hh7BKFqhzKsLDGMrKKIy7/Y9ErqNadeNP5+p
tWJKiGCQRD+nb9yovlmDdH5xYOVdfOE6auP9/IoCIp6uqxFLqpntKM/5b77yvQQc
V326kIyOMN1UB9Su4QJoeyKeRXKX+puFq+qJ5IeeNiehR1ZAx3UqpAanYYWDKfzN
sejf6stXWT2VkLsW3VNk2BbnA0W26z15FhdOCDz7DiJWeN31S9/5x9HSmLy9RWMb
TBVeQuYiE+4+lrBVjoIa2zGtIJhflFzhu5qlBq2Yl6xbytqRetxnz93d/FudQnRV
taFFIpeMRD42HhZm/l87qibh1VudwAWViPGveXc+Yn/BPWjkExpGMX7EXpovOrk8
4oLoTkw/t+7BNrEnMgG3iCl9ernYrT9MPBDjUFnUjmNeW9CFWeDSoG/4yu42aTBV
dxPWwwQZ14Bgp38o66dqrI5HFKVlZA1+fRXKkWLJxcdSltifsFA/txOauz3R3ER9
iR48YIONdXltoe3XDpWNOZNRh3LuozayK+0VRw7/5C6piwfaneMQ0XHOb2s/9Z+A
QLW4lSaufLLAmZmcOIeq9p9EFNYwCDlCL/hNK9DTbzanqmn7+k5yFsB+NO1cdWtw
9ktw2DKsOs7fij1o/bpo058eI7tJ4F7eOxYPyXv9SXX1sicpYy0m9YEYy1g9/HgY
T4A4hQaZebQTm1udX92gF5wWsEOV7V1RAh+1QHIrDuybRtk55FhDGYGmEVttGrmr
wg54IHOmmur3phY7tMln4P0qy89amJwTJsjEHemnyXZd+8RQ67kc1q8MXM2N2xnr
h04HSKlH1nCQOlppPpe5ifQoJGhRieoCILcIY4/iJU/tblVddbSxGuMX1Moil8yv
xmVVarHXKbWLq/H22X1Ijc842NkkgDXuvYhlkDNqeLgGPfGJ5oRclJDJc7esheve
ys1yZPPx728VweEbmn4riPcy3HacE7yRaYZbzsFhYbueaoMAH14WwFyAKYT36i7k
0TIqc89dv9LLTm3Zi3we1ImC2BsylcSAZynwKwrw0RftXpExb0gthwZUA/7BQRpu
JF1Suw859Z/8rMs+yrfLAwX5hV7cYfkLB7oBB5vfYMzItqz6zGbBc/Y+2xwrlpK+
R124fhxz/QZFVsTr5wX5GypPGWK7rwHaXwtieiYuhWcl0FyCwtlXghB58uqd50iB
ljepPor6wRmiUQaNEqFb66orN3MZiKkwj11B8bk4Mr91zjIq6SYWfxP5GgBRNF9F
WLJUZ3PRtoXxAG+scE61mMkD5b6lHIvhWlhXSngYSssGei1pJCluO3HAtYGceNoK
HbE3ERq0iBAAosbV1tmrvX3efpWhoWqF+qPJSOpNW8nhZn7h25EWccgVkR8kkbFy
vWhshpJ/oDDC22b+HRYGX91sVB8ATTj9j9TXz88ys6NeZ+fWuQFsO2lIXxxB0qcU
WJJiJl3ode4smWDQc7NrR+uywYEnBldY3NhVBXQSnLxUSdgNOmN5LWqWR3Sfb9Xa
jL4IKJcv79PGIO6fPcWHFnwcEiKFtA0baByvgBgxQ9IhifrD7WXCXDjUNMxnEGjg
dcEPVCEHDyGxCYj66+BGDNWzdE4HreehaTbLRP+kAV94Jel5PmsgYpbT2INtdtdO
jJEeQsRWj6GpUyc8Vc8TQ/vGnMZS3wZ7dzlCQFmJK1DEJPrGrAEfpBPt8U5vmAqN
NjV0zZreB6HHU3sc7HtQf4uDCvdE1YGcmXhxByMnGXd5ekEsjjfHTGpI5ylahFkf
GFgCvuZI2bGFDP5ftOkoThlj0I3XQfaA8dYtidXJxw4PDMWlCcJbUfbW5SVbegO2
oCWkyALLKtLBXfNoCSZ+XcUGAI47ihrRmu4zp26fZcRGM4WVP5GkdC3cNx+tlnln
6PqqVlhzVAJOVx681aOMIDMnrXksHiL1E0Ea7JRkTuVD5+V2wZUt7+m9BaMiUvjg
51YKHoOC6X4pHwGcSXV5/QMxEGBVulXcj18EUqGrEkTuTOvUt3kbrOFdJJACKX+f
w0y5QdvC7saP3a1duETNIo5NQXpHLq2ZwJNBU0IiU2ExHd54Aqn0cuLeSje7r7Dw
zSD2m11TQdYQip/6fm6704+ICBc7wAZpC0qrCGC+SATLd+0J6Xjr2vSBHPEVfkwi
AlOKVb6y25DtdS3Aj2qe0GLtgkA1MdIikKAu7MKFPXOCZ/uKtCFh55MdgQCvWFyu
/Kl+2CYdAYYVNxvW0kpDP4OJux1HqXDFYkAExld8GWEZQpstDfNdJj8YvxFb66xM
/Qubkx/c799VruYcc6oEcjQ40JHjsLvXzbGub72Ynxq5jevhmbkcUg4hPY6MZAUH
Xq2oGoefjZGW1Ow2n/YYKcod2Vnub3baPy63mwS0frZduv+4Z35r+LkyA/JO5Ali
+rWLUAtk6bHDfkkRu36OgQId2SD19uuqOgdM87QIoUM8qJanI6QjBJ+N0dPefB4m
ibuH78hebSnByCccsaLd1w9qTLsN+f0rq4zCtuCZwqTQB7l5bH5ho+71rpaWJ5Dy
TM2gaKLMFfQzUQQjK63ki0lcnPQAwUcpWemhHOvDo9JL9RsntMiq85GoqMyy4SIC
zEvpzD1sxxZg177gpWiKhtcbLgs5RhGKRe+hflwkKFw0xeFHO0drPp5dS9UV2XZf
69uEm+3I8ajXgIceMtq9XBsrrgXY0PZm3kMIPD3OzlLf+bncej4enP1joJpjwGvD
4DPMwwuz+4apX6OMzQo1qsb1ewyH10OokYD5GUHJu9zikGSCSKvkW+Mjj5sb4TSo
vl98j6swx4QYBfe514fH7R44CQLtDY8HrqrUjNhySk4iqzXDyeZJpbePUvvrHF1z
WQUU5Xc4rp5VJrb2gOqEjAGljWBMV1pZ3K+3M7vjPbEJUfnmq0vspodPvKS8g2fW
Wnu0ymwA2D3eqeQ7jJPeFfSpoKx8P1ed4GSgQqGEjJjUUDFMCBni9fWQdpqteYbE
cGSpFUmlksm3goxUNdqdp45phw2ZWAdHzT70rAAXsdt0asY+ZFkd/KNqshMTYaHO
cw9Irt0tClN1kL8EJtAjilUErJEddGS5fC8w8cODlPJvcOBYX1gfn8vCRfs9Y5L2
cWwV1ItrVxlptBleuqHvHq53aCWuhsR9H1rW3yF1F2lmzDpSCApusYl4B7h25g6Z
p5A820o9PqY8vvfGMB1wtY9RuwC9U5HaNgB0jqk7JfMC61qu7W+42nXRocrdPftN
eNFVpM1wF+nshx7v71SijwGpeixoB3X4P9PRr+7GWy9TXkdU8aa/BCDZpYABEMtF
X+GfMx3AdribVAFoWNNH6gqJpcgMfsU5eMopeEDkEdF6jssaOsv45Gx5BXCEkb0w
igNP0XQSbtIPrn8mXq5EgJu+H/HOQVV4fYgwmMhzJ0YKRV9d95OOARkhwUcmuM58
OD5b5/XjYrw8+/qO8lmsdzsXQhxmW5s7rwj0eTxZTf46U/iaoYAM8ltj3+69vOY8
VlJ+/2qBcvfWyLb2vdkmbBo1xgl+9d4LtzoOFd7MNLav+0qBch7fHd2q6yBC8lKx
KIYl6nONaa2bbSOE34BoOZb+JSAe3Zvz9LW8sshhlYDhpodXec9Ga3rcRLRHYtU9
rPtUTNvtUcl7vJKf1EkqWZTaH3n1h3AFF8Fz5kNargrrmkjrhnibCgP4ZLR7FTo+
qHhwXzJRW9TqViF5yYal9Ko+/Y/WzCtkin7h8y5/r750YS7UgoGcGipV8RUgEdeJ
44GjyTBkx6HbP3w39rI6oRP7k1JsCHnqEyASfHmONWRSjLzq+TuDnFP6UjuzaAph
gxBbaNJTfnMqvz6+epXoZ0zzr1hrVdxKUoHU7OaXH2Rhg0EC6Pf9ocqXfYTzPmcU
uXrj4QV116K/vdtMeFrfNjl49SCxq8hV9K97VAZ8vKkOB/tOrG8B6o0yy8fM/Ry2
Y+uSye/4V39OTKuP+NsdnjEDfF4YF6Njj1LuLJNZHgUbUBiNl1L74rW5GMfqc0tv
L93+mPod1QWJg+E59oLmMUlgtJP3Wi8c1BekCmg89R8+OpBUNK+To0NtT+34Yq9w
aCBNFgIi4MrZN6tXzd5PikvcuEe2mSbmEMW/8qbezZE+u0c2Xnm/Io5f/f4/HkvF
3krf3ulYuv6lBFGAcgKqisYKBh/RSUBB4TorUWSqH9R0swh34rzB4Z6i22bdHZtx
LFxiYh3X6W0uRNmwXeBJhtxViI7ajV1yN7g71E2TUqlkvKnwg1veQshfYjv2dGM/
XKpx05/SmKPlSnwiarVsIaHZnUSW0uC810b+UPGBHjX9c0FTZ91BCyZK4P28p0zN
wTmgTKmTL0qzpuGrQ9FNG7a92V2f+OF5mB9wF6BZYGM=
`pragma protect end_protected
