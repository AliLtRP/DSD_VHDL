// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:31 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
p6hVBJ3S8UAPXcinP15Az+EmRc9AoeBEaxyKOiJOr3BMyiFL9g/eWbkP1NKbtpeL
h2o3Z/m7PXWcsrHqQzUJBZvgNcv28JnHjKskxWHX4iRwEARy1vLvn4IPid4tfQYr
pfgmbuo0+5i8mYgFF9KDpZYWABaKB8tkcfP2fmhbuh4=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 24128)
WJRGmITPrNWYrFE9WUVOZ4sCgUYa6eNN/6RcJHlwEL8nr9W5dW7qEaHMmeAJs8UF
0pCU3rq43VKkk72SuCo6HFsZxoV0TQNsmlTvRa2bjt4xoiIA+g+lG9/J+5wif+a+
i7wdcg5Dk4YzwFUv0YdQjaV07EDSCrkawlnjsfW2KEX6JI2OKIF2kz3NYksDZ3WJ
5iXMybYBb8Az6JnYU+vgapDEcyTCDyKfOoicMEg4iJFFfocAgYbgEN3xBHMbeGcw
648u/vebm5Fkg5pZB58wTCBYdtJSeEPvMKxuWgJVv0wHAwVGiVXgr5o0gcWQBaqz
iUfOuCIML8pft6oFg3iprTuIodbUsGckX0EltKK3w33tsvbYDOkKCcV8WAD7Emut
L31Xsw+e/QgHv5we3VEmbrvib/dKjL2dnpyAJByFsdMSsHtuinKWkd032gLbMe1z
u4DF8IODp1eFzY0ipCNbvr/wXrF7f6WFkzMnhecKIERiWoPq9pndHDbfFYciyu/L
lzGaTyb/VU9eYSqB++FCJjOphvRrTBYlaK1pfD/kdn1rlcaFllB+mHWSwa4NntMu
OBFyMRnalUZF4BFSeFkkjddcYUAJHa1jci96u2U+Te46wlCZFCfqcilqotLP2t7S
XmJsV4Fp5jF/Y/oUAUOHwUkT5en6gSKobS3MmfgzTlDUE2b1e41yZR+Yx1TF2LZg
ToWig64tIBdvXMk7699c2XpaanchiD6Ii65Jbu/3zNA+9iWzwOJ2Gc/bvV0xTL2Z
emL5vrdpNgganMX7ZkZHcGA+qw0txeuApRtphMonLzFAkHCWmb+gwPSdYF0aHc7K
rKEZbr3R6YD/OG+jqc432fLCuv3wo3kdZBRAoEbO4IMCv5P1KMuD2GpzE+SGoSVT
SedZQpSLnKnnDcZ5g9A275s1rR/9H7xy8mkQyvfTdzkTNaC87081ESOfD+pRbbZ9
hua52cGS/mrA6TeA6DwhupKJA0YRyHRBh/Alm4U19MB1xHIHWs9AYpo+ITXRnW0A
iKafv6PwiHK5XJ34DzcXvS5lqiF5Q6COP033hGBFGu5NxYdAyaDI4AuXTxS8xWeq
4Dan6frGpXhpULYuJH3V0fXvNdlndn1hl2dh3kF3jIvGD/m5kAsRtrghN6YjIyM7
OaVtw+Vnux1GBa/yJRKwQx93dZrcxsPZDvTPsyYAAbIu2tzkvGrxrsFBnfeijw9I
ffNPWXsyMyYaWVmFSti5mF4CeKvLaH2YB27wVf1QavVuDj2a2/VYN9nL7g8/TqXl
EXQu4awHTw1LI4BT2EPvpOuiXp256CygE4ngaK9+I1RlFXxSynm9Altlk8hSkqJN
+oNtyYlY+sqTsocT8bdtnrG4IHolmqBSboRfxSHPWLlFl84vrtzlnQs0lOyQg60s
0E3Gz/XgmkVo1NYjbbrINpfkVKg1WimtB+nLdi9g4KyifPV1WjIkaH3pztoPtofg
rG1yVYzfJRlQEcrUIxr7+fZLH4NThznsEaFmB83xGhKGW9eKkV0p1LINWldSRCLk
0Hb8lXqt7XpU1ZPB60WyAy/BTMbY409yQpHUpte32k3W0eVUiNrAjCuWdyGqkFgO
oMQw8neom/a6iIyGDXu/1GGPo6fQm8+koVbzkX7iaRd/40LuMSaDAZUD205CM5sj
yEmRtPU8HZZlveI26ZqkSd8QFM9XdPNplED1JX7JdxrxdxYuYxTOgBnQdA4smStM
ZMsIWto/8fFxRpO2zuLOEPDHlpv71bk0nqWPFdU06E/8apb+RTipY4CUxnqBSq07
YdJiyZV7xDccMcQtE2SBVe4g0gkuIY3ynVd0Gu7bbFbZqQLS0S4szTWDJoLFW8Tb
pqR6pJMAzHP2aBo4XHKXNSmpsNr6VPZEx0JIZeTrue1oKa5zI2sHhkIGbQLvGEHL
TcARDg+V37dzc1AxEAAjYaA0MpqbsrOpF6E+NGkTZz16LGkNi4IRm5zyv8etKSde
vr2hB4YsSvou5QvV67WYHOINzOl572BxOUtW0Z+RG7/qDgHR/f2kcV5lS/0Kajl8
/VY2A5obiR+qqOdaD0TpB2yYgx7k4a56Oy9uZ6Aq00p47OPhOy4S658f64LRkMYs
RN470U88TVmtGig6QyrhA6QKHUYN3ZRQDnNvzpbjxxmkrf9cNtsC6khwm+jZf9Lf
dSyz4q6u4JFsRaS5u3Zb/VOBECrjwBgC1d5kTvsqARQiqJP5BZPKBC4S7YrhEOUV
SEUI4d2mJU/5jdXabwVianO5AB0sexgLKlKz16ZXgmxwx2NRXxihOMP4OCtZHFD5
whlicQ+KxiYj8OmKng6hn1eijOjUy/BnneRzdK5qZfmNztkjTk8UbAlvVZFQYLfp
oKlZl94duCsaIh8A+/AEQN13j4S3n27fsBJETJeOhizNJKVaGk2fFB6V8VU5zDSC
n5OcviNcCX13QPUXwczAXMo/QhBiNQocSIZLEtoGlTw+dVkYTYdWmHegpneUzIhZ
k/WQaY4CzBvXy5e9BUX/OpQTK3q5ABT4RPzLZFLUKVkSpeSsgDeaBYlRMCST20Vd
cst4fs086X4UGrvSymC1hshLInSw3i0cJ8e9gqol2Ik9lPbAjob1sOZaooJCaSd+
qv3ZV7xSf+irvigPI4cCb2uXxDz5gBbmWBOoN+Hwp3FWHdAkx1Heh5NCTYC/A2wJ
RKCde0AxWi7wl2OlVlCOu3lKBFcEgdW8YkbvCPnFn5QW+zCARTfZiLwh9ytH7dmY
I4Uy3MGPw0Kw8fa2RVHvk4WWGAYHKV6k86GviTEjJ+p0Q/EPrVT9CyUP5q0cacOt
DcbtUF4w5DyTwOcqKr5mPk8DVBqpCEYvUwdBRlPVW/nxnoQqqEm5gEc+Q1w402v5
EN7cW48ET+i7t+yOlYsNU3Ktrrp5mZwBdK+omGflElh4J+Wrv2h8unGdAC3mXtjd
+4JuHUi18msG5TibUFStzPHX988a7JsU2iWvRL3VW4GPwHZdZSuPf2f1tUqywdPe
561FKJY3ejONNMHDGOjukZ/Ot53VtKdUeCuw99Ye2JGfPW7hxoJvTDOh00gkEjhu
pbMET4n4U+EdG1DnBtkm0pDufUCdml7GdUw8wsuD8Q8DqeJk0wqH4esmODAL1fUG
RmGI3Bn3L6cFC7KEm5MkST7NvNFDUlGGIWocDLthzbzPgkfcH1+pakAfuRpWhjBr
2pr6RDy06HrwGk5yC26v06nUek6KS47GAJ2nMBX9avJxXuTef8O29C1IBe8n1LFA
t0mxxEljl9dAOU1ZSFyMuSUH+waFwXpDZIXf2qflhY74RXrIaLo/rfV4GC57EPiG
rAHxYZq2E+oSlYps8leFqF49/8VQ3kt+57Vd+Xvv88AC7o3P45p21padSiHKh/b2
X5aGyTgw84+/qDtqxI7XYP21UTmo83wCSjXMEtxU3nItcCFZXI+5xWAqYygh74zo
qONoCcZVTD5/SN1NumbctHm2em3niTrx3MvamYcbhk9QA/XKZvzkfDfKnjBXqxMj
4rBOs/duRRRJbM3exL9xVm7IdYFpYUKouq4WUzRssmTFmHqR+PT1ygipvh9KEB/y
nTN0heLtnaJLETKwRg/PaJ41RfyOpCAjmCkzvOAHUT56n2AkzIaRqMDNMMAf2yP0
ITqfT+2oPdd56ExNqBng00PJcFoBtCbO/kl7iJECZ7g/W5HJJhZXB5xGmWH8x+0s
Ydof9fh6mYOOc2lG9DKmNMhXaJ5BcvCB38ZLtF54G5qhYv//kSGXun9o2H/N0kth
Pd7VMNva7U0o7mtgeG4OGukscMZfaabhjdo8F9nTiWfmTG55yDsXq3qlLe9SwBBv
NSPNY++k40T0JQTxI1qLR4L5s31vguKtLLsfGPqCedzgBUo/wLQ/vDotYqB61DiN
v2xESRvJHTA8I7yKMouaDk0diAoNWNTE5QLK6AzI7/DZSNAvRrhOVFZTi7C+NpXj
PgQBECrHdeT09I3Gwm0Alusl4Bs/M1gfPgTTKdLDVCN9EuwOspesqY9Cg2JD1llT
m0yQJwZQbuk6YhihZjNxFvCR025yHA3+LRJcFZxj0phafx8DXDhWzjbP8Dp3llCI
BAKd/9XKNiz6t4hb6YJn/AxsksA+gPnAxxWNekrpnk3JGEG8HI/DBEGMRlqABwpl
v+yxhrZyfU8QUOHAjeKH4aF4zL6NHuD3V/MBoez2AKQPPZbFVbYNPQekjoA51Imo
cMwUCgyWoi7WD8wJcardIqYzwHmp3a8VQm0TcYiWLHr2QBGrtpapH5yyz44NlGc4
PsOYSk6D+JqopfStFw+N0O+VSzPXDpkw0UHVJIBC5RatPXhiAop2eaYgu6FRjaIW
In6sxfUZ3rA0JoVaft02zTuktMlbZ8KcGoWvIgFb8wbtgWm1KYrCR1j5c0dMEZ3s
bJ5zf5DDL+/Wv+OVXLiZgik/csapH5j2SDgohFDbxfhE1FKopw6MlZ+V487TvuvX
/gwRq059doVKfYQHW25Q8fuJDowPUWjzV0sCK9pyhNPzPckbp2udvjVoRj04rW/l
72t3KBF5U54Q+yxj+80Xd0EfBmE2Y+Ouy6De1jaHWVX+V1/u8XhBlsWjzlKGzx5C
0yekSCtNWxhpZCltZMotRujEFlqa1qRh0KToKfYftHiKj51gXy1WQvaqFTDnOcmz
TVnamSWHZnVJ9+aexIsthkBtE6QfPD+V0VSl4DrhP65Y2JUaig3oehc9yT8JJ3su
7IkFlBAvIVsjzBGlESeNX4qSOKE3oJs26/wLEaAZKZSjN5dG5UvNM4G6AL/ArxZD
HELXM6UfX8YyEfQl8vxfRzzny876cQbjkOayrPmoZDY+lb7xa9eKLzKTAXQhQlqb
5sWGEQcI9LrDMCRxRuQAgcqxYjdCLQQEyktJmADvK6q42fPX971O8K7a35CijRep
/AYFVNhnnnt829Iyd7npV6jqLo8ss6bmj79sHzctB/iXNHLkOZd9hJTuhLkkyE1Q
HAJxUMEnO4OjUl6parX4PXR9vL/AJL/QK1ur3nUPsIO4yQklixzPgm0iW0HHA6r6
SsZnbqFwPg44zEow+rZfgLP3jeoJ2yz+5MB5CZnnLE/tEediYf30uohfmI7sty3g
bMU/Dy9ujmS+VD1k8LymSQXxMjtIWgWLVYABy66TLHa70buynTmcAbl+2hVkOGCI
+OFYEjSaqOM9gOGWhryBOkUEjWYywRtqtnu1zOU7jPrxRiFmnKLQF2T6rJf0ryfO
PJQz/oKRDNNmauD44QnAklIwBOdWzuU56Ah6Tiz2sz/e4TgnzjUEBPfrdBQXf8iW
YTdxtT/+tFOClHQNUVfDBcqTcZUfY+cgp9d2U8XkUmnLfM4YpU8LDr2ufbVWD/NR
tlmHg7qDmenbwG1/OPBBB/MqLx9t1YPBfgkBst8wARqhn3Vo5jX+DOcFpo/G5h1N
GhVeo5/5GB7MODK6zxSbnFt/4m6BfowB7yCf5Ncxm3kKtMD5ORXusLyYcr9ir0Z3
1VNq+LcyAxM+loKlI4Z8gw4cye9HM02elGX/YtXEyJn6iF4aLm5US/8rsf2iwmlj
cmVfGL26BJWRffB0chpJfaS2v0OhUxFOZ6GaTAewjhvYIC+yvc7+uh19Hd5Pbc8h
oLfQGVYKwAS0roxTmL0yBbhZ+dAeo796jtBYUbZWdMZp65XLX4xMbjyaaZyx0Lm3
vCu7gTQ6K0v+cnI2m6zYsrkNvdzXMgHR0DE73EQgkMqbcLgsD24TLNNKQcqlUPbD
9K7vCN/6RpTcyho3akRkCRraQnlgeGVJZQEV1BJnMWhU1Nyngh4GqRMQzQx+6Rqn
RgD5DpIVtiTsDeHt43zNS/L4IqeYmcInsyY+oHzVKoN5z1bLCIALM7FQYV3N3A55
eZdBBJxf1T7JlVHwHnnXH4t4toAm8gtO9zlA2Wo9xy7cwTOR2xzEP1OCkH5Hhvdb
PRewLzgTAScVbMdDJZ8Y70EsnhQH780GmirQ9dYRTg26F0s1z4sd4ZkDBDvvIwCJ
I2oLKVYXUE83ITCcwNC0RwGlZDkbm8xSvrezR6n4930ahkIU8mORvYk1NXIA2vng
0TVST919zwE+eGw7pPSSqofbJ66BA7Xk5TAdKD52xlQERyxI7QgaxMjyVXr3qayT
ETOCllQseojdbTsbA7YaBJ+v/bjkB1EUAQRRwgOskSe80eP9uPLqNWAzs6YxTIxC
JtCfEZU0EgaBP9WEtsxwv5/flDW8whVKmG8WWPEztwdi86UW6ptSgE2baM+DeMAX
vzzoSjcpYmU4vrmzQVjjzjFvD8Bl0JJnIkDl30d2SgH1X2tKzrqOGQhCvS67mnJR
uAD3Ysl2a/CbXqqEINTWGzgQ+jtEa7Bw0oLpPQi/j68grqFKFF3spt47zqllmNML
dx4uo2TNbfo6VJ8bGlrkHtJ4uCNW/kAzljisSaddEY+hTh7oM3DQ4OCIkPYjAW6d
1xMzg8TFqtfxOYK60Qzy0MG1hJ1f7AjDNCYWampIgzvdaRpdY2n07SpfWgsO4lXt
9Zfqvp0p15+MOZrF5AdjJwA9SyDF3PBYy4d89godJvAOPjbRX5K89AEpa965TC/L
QqArg33R9ZA7EV2/QaoFnRthdRdLHyN2X/v9D/BWAeHY9qPPFeYktL88usG39mR5
4KSbbSfPZZQIpxX6cHryCQIeE6v4or5SXh5wYVJLG27QvOGau0YO1RRLlZrERJkB
2m+gyteKEqXh2Ui4BFi8dSKdepeD2p2UJX0Nopd+K6vqEocdWpToj4FTcggFpJRL
ibqEGDWqAAGNUiSYj5IGF80aP8p9nGuliu0KMUcTwwnKXWNjBNuuliemR1SQlMz6
aXQzSwjkS7mddBKqL9uOgK/qcsOdUITYfUvrS8w1lGWdAOQn2mgMU9Mu5LyWhcWx
Ih4YFkPE0h/aLcpEQf/xpSdd+vhD1Z3Hj33H8cYJ3w829nU4X9gnKTHa1IQ6sZZa
op08KiTvPsRajvJCqOuOC+wSE4bcZAri4i+6D9ETTTR/c5cA5zsN1J994M65IoXF
yYNG5IABbawyPm5dW9KYAZ91Y9fjrZ26kFFcnI1mkUkzuQeDQqUBjaAlP1J4y1rl
MDQOBt9e+RJq1bB6YtIJK6IFIY9v20iJdBjSMByhAcSWwgur9vKk5/Fp50Ve8CqZ
mHSTjn2KC78aF5y4xzl3i6fj3A291AzsGK3vgF1bnxygkHmx1nDJ97gqMwKyCT8z
RqA3qRpelaAnyZy6dmvUBDShsaBr2SfyV45VLyCTFxHRds8u+kuHLSGyHdFNbX7F
ZYtDz9Hb8EmlLHRGaDkrak7A8S9M+ZrExdQSQQ69bNdRYPFkRd0Wc26JXI67bVVY
bV6AP0ibZ89TiCIQrAud86fAhVygcUmdy5yYfXUvI+zLZ0bPgKkH8LIvJ7ursBxZ
DEalcqXGXmu9gLAvKB4ntyFbDl0yZlavabcdK8cnFnWjwnw36dzJ5BC93VYhu4Zp
XCjw1491wv+ZlpCtEZGZxbxpttYGeBhVPDzusapjMR7t6zCSUuP4TqyFxbCvHOzD
/RBR1n99nwDx7zx0zzHgNEfmcnAHPo9YiKPKpOZlqYxPRx3a5ksSipZB4lDLs5Rm
cjjpiIdRK5K78cr6H7Htfy8ztzE2pTKajFIbU9+Kyi0EjK2yFztMDgAWAgZojKbA
RoquVFdP2T19nePJDYEyUzetKdPHqhJMngeuYraTxj2NUD7696dEE9Cg7nOWKE9K
V4JULcxjDwWZk7Zve91hnujHd3q4nf7/I/nltx6rjv7kwgcJx7Zk8ZhPamBRz04v
zmEcNLdHRWqrXttu2IjcMHNeC1eIoJFSxMomuQVu3KYPKzbIq6SRKYA1N4lUe918
ZbQJMHvTlTyfi+/ZWpYlx2Q9Q3DkboyAENndgZDfu7zSq8S3z5Zy2YvQwO/WI+AW
nmDnfqPSZIU/VqnTT5OMYyHKKDD3CdtwzyH1gCswc0xeEqwJuMWmKrpdG2Et/N54
rfbuB7YqO0TI342MB8GbcETd2XYsIWE8n4tFr4PJWRNGmxbBfikUhE9ziEN8a2r8
4mprYRHgZDEFjzVYaiNKbDHHOWzgrkJ+MitfXNq7pAuVs4M5gSYByXCrZJQh6Ox9
wMMxACNk7ROdO8ij/rl0ceEtbLRWpTVD7ZRR6Cuh2ESJRAOabau1cYf34fjZ9vTu
IsnOAIYlhSUr1y9S5+j50lfhDcrVvXRFnyPkiKc8Ymhgvgu2w5dSkPN/1fCt6wdB
Kk91NguADL7M9bIoPqsWaVQekD3Km6mT6sCMm617nvso3xeqzCmn9MByvkBIRgvd
PtozLqWtlAvVEHVxCzVlOrVhxwD/YCGCcSrmRP0PxvaifZfBd7RQlwy+LDIrRHoQ
NP/zs/RMLQDi38/vFFgRBNXEQ5Nn695n/fyOV94yaiv8ToUg8fbW24QDYwXDtfwz
giGi7Mn+h/RtXMuC+Ch+sD7UV6oJ532lMXKKHNGxRNUbx9pPjsz44TQKbIilW5T0
GLZcV2bKL9OYN6IoGLS71Efv3pmrvkOy7YnonUbnFj7fMnRED7fr5bRXuTgMR+13
1fx7Ml2NraIpGQTARA2RrQL1V/4fLJBDpu+QIy8d6LIXqHuMLp6sQxZIc/LYpQCb
9ZuB5jANvsj6mxYht0UMGmCSwNC2FIi406/8jNGZ0SV3d4+JxD0tN+wtliKCk587
DwVWUuMde5Gewl/h7m7JzkxAddrJnxRXncXS0RLDRa5LPcnS/I6S5dXsTpYGtWjm
Jny14y/4+3us4fpPxEaBWpCcMKfwNN0O02gCnbURWm4/16C1MFYVjQTXeN4DodH/
yN1HFyVOZm2YQbarfpRy5IURXg4KEAKgpNwFx6eINmOExQROj/icZv12C2VRdZPl
2ItUL/NYXsRu0aqKGeeDzz2DR7kZ1cBu2kV36hgr0fH13HAWxB5RJhpnFSoUoXfW
4pGcGBtdCbeC5QxxaStmfzOIGUMuxXzWebwPdGlGiveedkE8vn/26buy/RQR91qu
2ZDNqAeA1Q1JGOgIQY1sxjUCCxyFhQBfRcUfK7RPPUbLCPXELqMLDgKlFbOiRFfR
4B0E0VTrGS6mMB0V4uYpZby0h6+B2PmoN/kjaqQcT9GBv/6apqrffVM8VbsvM4OF
cTDUsUaUD0e2WligQMUtgK2tfPEyWV7Yc9eeQkqeqkjsYFDRiv0NLn+OUWi26VM1
W9HHlixJIjF8onUJUEqATTgyqxTZEoJCYujhJplkseWrOsaoerCA3zmtLw+iXpoW
vOIUyFG+W3FP2aOPr8TML+CNTIjRQZcdYDdSdw5PjccLgQzygeEl0ydSuF/WSn7T
J2o7GfDuyRc9yNPKBACD2ZriyebtHhHYjOyfW2UYTeO2gBdIE8D6U5HUy4yyDpZp
WfrBWmrHiNsyjLSt5C4EoIvfmK3FOrNxjZXRVA4FOYC1nBKL0O9oSjHk8kw74nin
E29rM2EmpC9gslMHF+FbbGnRAyRwPMvyyux3EQbRWJb4AzsDthddTBOOvVKu5gUF
9yV6sibMS+RxTFqlQgBwfbZlih37YEAckgWFYrC9bXpo0dfYzBeRO5ChGj2rnc0i
REY1bgIGIduEcIrwnTKHN6Cev7iKb2oofy4iO6ZncfIGjv92oMFPpYA1wRLPX3/2
D2QQvofjHHhyj5OtJQuYS1UwcM1FJAm1VENF95sIdBDXNn62Bq+LLAmHoLu2/zsU
8kmfBPBZIKiTrNNJK+Phst0aqA2nrDIhNruW20CDajNYalrsZG4jIhajzoSz2rpY
nAwj4964uCCMsbc1SGRRqVKE6Y6XHxeOSEnp4HsIdpZcRkCJkAOwjSCcINH69fAA
gnGUkYIRylXg7dlo+0KBptP0PyF0qY7x27h8pT3BafkwSu1cYjzewc2wzcsdNmEJ
hzsxiRJKyqS9FztBIyetHA9AjtL0ePqWeDpzKbb2OiVZnSmOXXiyszwGyFpk2lKk
gmK5LYcXLASi7KWptK2PaslO79t2ET3tQ6vRlGX95j6EzlZj540vUlAv7xSwguol
dZeA3vaTW5R8Wl3ZsuNYnLNt3lP52K7EFQmijzzdnght7w2S10wKtNYUK9Zf4Znf
AiFuDGcegDZNdHrS/YkUpKYwI1HyrcO78axP5twoQTx/9zQRtHzcZ+/FYqZhVbcq
UeHP/9l8cFaKKCtfCV7YiyI3X1RolcPhWBq9AdIvMhbIPHCo26lp/75o8Lq14/3Z
kl9cyGiXTma6f5nGIglt71Aw8tuTXHIzk/ohqONxC2lMqn2PpLqZotFkvDOoDCcX
HcTgnSRbMjobfAq5V+2Kxmfhiii11OmiPalJhAhRwMu043zhyyHkqWUlNeLq7umI
Q9/CaC3MyH4RkAhOG/ZMjbTbk8J8zGATbjfWR5WAniT7/tYqtFyTEo2SCxAQgAuz
fHXykaorkKib284Z1eSlAViqYiy2CR8h4AXwWc1kZufV+mIAqWFzmFkTcJQILVVn
k6yowzOAKDidN0N4pDml+xkYRHblOPUQYJJD6yRYt4UeCPp7rX/6njDSXdQ0NV7s
A+Jwk7a9LRRQzvvsGre8pN+eYVMLhYLCM880OYn568Wf4GdKQUZa3OhmP/xI43/X
bszuaezKUqVpQByiNYCyG+gby/n5TIBsWWY0Zng8RIOi7G5/XHIawKh0HB8eK0Q1
dhZjt81L3QQ4mE1mz4ZID7gFA8BjjmMZzm0BFlv72PsXlwpixJlhGEHto+FFPASo
HcjBWb7gVuMSDbRx40b2ygtq8s1KpKtbX77UuWMAgap1OR/ZVvuNQ6UH+pic882z
ElJReD40NZ/vTU44aDZRev8dWju5/EfKHgtjndBoHBczTDg4kkPIEFNEblMrkc3x
AlrStzdVzjwnWhv4ihDjILWMN6DuiBUJAB5o42zcLzfEu1YL49ggwDP7nJKdL1F7
ZzBqD/6MwVHtUZgaY+99LOQz2kkKNzxm1k/UIrSn13tYCYIdrOQy7VMEagpYgTzA
wZuBEWKYImc47IchOgMCI3s7u2ciqv9YejFYRdy0kaT+maAs09GEJzKFo/6CCx5m
4D+w+MhqNjyHS50Mg2ItRESXckuhcZniHALz9KiilNgtfAlwtrE7OvoV8jrgq5bI
jjZK3mFBcZkHLK+8SpBGHtNnAxcebB/V+mWKQ5YNSulaKQwJO9YHR4mBNE9MaGzf
lmmHnYN66uK35msg/gh2AOWrXg2OVWMcdaliccCQ6jr7HDyAovbwXoyqKRzYg0Rp
+QiHd7duyLSbNRmW7WZKFsX+OWwavtX+ID7IBl0XaUJQPLOwF+dVySQsvDEb5Oa2
J1IPtQ4zbkLwDrj/NQpV+KzQtCR954gvbb/ErxpFtHTM83E3hORih0tRq3rtIfvk
2BXOjQQprTSXmTSH1/lgDpo/Poz6Hm2P2eYxfumgO5mZui+9zdaCQ+TWdGIuE2c2
5Vy8Mg3995W8XnZQGLySlACd98ZHL46bpX6TtaSdN4iQ5Vw5Zgpo3GYaXJAYWXjs
jOoddnMx+TzE0i07mwYkJPWeNvEJGQnI3UDLR0exKWFPKhDh1gDrvoBvF5cxY0WC
+G/yg7pZhbwXQX+1X2taOCVu9d5SP5/bYv4gp01DcMzhKZ1l7NM7oBxTF29En8ra
amvcZjJMeJq5fO2Wv73ngt8daFVwcwvpiVGdjLjkQrM0XtmeTBw20SbQnDavCr8Q
j3TS/P6WWW/35cNz/xlqhvQcMbbTP9Rn+p2hdZnJSsULROu6GRaAQqLuHYEu2i2e
RfuQrg6bag8x2pzevyiVE4UfC58mciPFByPN1U9FBoFC1OhBetRhoah8MMmhmSDZ
VD3UdmsKyHEtiAwXytrAf3FZOGmcqCTt8zIVrY5oMnnnNAkKiG+1z1etJA1BAJ6N
/DoB8qxb2BgOAWoICCgI7wBbSpWiA0vgIuuUYUzeQuW/2opcVctAvI7eI8EJQUwe
CbGoc2CDafWT6ozOM1lsBoUQlnlxAm1o5KLMWJ+pDECWCzHl4XHUwIl9cu4BXetT
zmtata54Gw5HA+vi95vGgkpkUVE/vLKKWueMFul0IHPAu0G4L77aRJi7XIcL6Hce
u4ewjQcwk68iZBXPWIht9kqPO6eZX3PNsaYOmMHcvTKs8dDXjlM4xr/1BvQ55Dvl
3fPuf3Nr4HUv2aNrwzr5k09Sfp1iljhK2rLqWkAMfY36GQ903NxDCcF+ZEFhrIvK
ru/+e5f/cnl0dppli6lQIKVfYkZkoSwQ9+BHDQhTLKdTnDRrw/7ycjnTc3rLxCcp
E5dpDRqQAoQcE2apWh7KDWG1kNDP8u6rpJw47uJTc6rQEVQtvu3/ANlMGYKEse7k
HB83EsZytDkPAqJ8o71mkXOl6ULlZbezfufgLLQmKIIh1awk9kDwpYWTbwVVsrlK
2nPxUuhw333Uk/1ySxkxCqVR3Cu8coHUazDtPNP7Q/N9TrVHKv6A/R36uxTiIG5Y
sTCNaunhISCUQF2X8TIgc1bL/cQviws1GgiLa+2HEeml5y1j2CtV8K9QyVTLVipH
AfesMzNOYbNBqTSwxXfjvwD9fnX1qcTJjJ1W7xjif5sE0p+gAoyvoUNxsMNpF/cA
A5HF0cT8H6hFu9D6k/OSns/iSUpZmJAs6IZpJm2CYU41czH+Plw4Dfq1ZcHCiEJA
Bbu8xZHOBRFT9PYggMvadl+cd1WR5TZyawL1uBN3ZiTYd4tT4I74VT0mkt8nDl9J
8YWACbIowslTuMa3L4WCdOty5ohvpx35iUDLqxVgyPya1Ug8GS1AfuS1lBoLsGPP
u8W5ausYmpgeNSJOkY270BYklnR0A243vyE1DR7/0oV5e8qPAZmgnO8WL7JQ113Y
elLJVFp2gxygv5rqjgmvwug8Kt/Wjq2XK5RFcPOyFkhaXE3I1/fxslqn5HhZw9x+
4Z/F2OD1YXMRp5LenGeQkNuEUzis2JB4nRvX32+8TDiZMAjCH/SM8Tpr3KEcS/2r
gj8qORIp0mOCyeBn9CMPONbx4Dj0fvqZIKxW8pTO7hoBZcCNVob9gPbegHrX/hFI
s2x7O4/5b4I/gQqF6nAjOlaOVAfoFc0AVvo47eAnO2V3VflwOoL68L8gNY1pNshG
LFW3jYf7yt0um3/FflokwuIO5YA64jhz+36F0D2bFxzPWpDm6ukfb0PT+8jSZwyY
9+P4cPMtopJQe9la+dKmjxO6c1v1CDc9l7xCO2cZlZixyeBSMWVHVljkePFvDHGj
hNWZ49bMdMymIRCcLLq3AKBTm6diMEK1DhA0oLMkI8eIljcP7/GLvX714bMhtfGr
9rnHOsonBCZrQzzrGIkTfSJPapZjCw4wbkTN6ulQYl3Vc4s7jZqj9Emwu7bgO1T2
Vb3G0CfHRdnVXHZ6P46YUP2CdoErfxtzcZPEYManztaTkVO0aRy7i0h9tpCY2CVZ
qK5ah8pj+fG3GHN+0e0lB10bNEILrc69WadMNBlnNPlYC3/EKkv6s67KcwcLu/v3
QM04xuVXOWHeV9Vg3TBZZhCP6V0VHB9ynaDTd0h/aqAIVwaw1LwoZLe5EVqjzBKB
WHT+VjcoyTyJVYsz/59YFwzas7UNYOPyuBx2l+rBLwN8fEZBwQD8f1H6R3DirSTu
dgzXNe3kji4GCCjSi6tJONle8XHdN0DfBUe4ruJN82CUGke9msGm37FsIZOYzAR8
O0Z8AYcXCtX1yZfcDyKwFnqOegjszcBlB8soggWhfjSrTdaV83EHvAvL+mVLV61D
bSlhbOA+5u5rj7uaBVJ5je3VvGXlqbNLpfR5mjQvr0reckbqkbav6NPxvAGa9G2Y
3x5STTLygKgserIvg/0Y9zugXxSFAUqeLPFBl9lEuACk4bmgZB/IeaVAY8MS20E5
RhSNslIKWSirEzm45bCaoNIyXWtHVTsXGPhZCAYdPx0/aSXNzLvyQOxKhOGVNiIn
C2s4e8hInb3hW7sUE8LhntlWf92kWgHcljUjWLwZGnzJ37tPxdvsrgWmetgguf/n
8swoCBrKVyFPNDF18Wyw+oVk7bdQmxJSsAei+E9SEfSnJYsl7odtKU3j4msONRx7
5LnjTNyahVBKPvQm8PfznXCTRRN0gHv8BMRkZzsMtXi0iKENCZK2adSCfXYoBzOL
Lqil2nAPue8sh2S7LtB4W+kz8tr15/LpWt8svjlwausFs8bw/IQKOD7gHxfvsXrN
yAJ/AWAXRzzdWVyJtkvBiLF61cSEym702gK0c/k9Qmh2AszYBesGSNUA5eH+XwDs
jclXh57XsIMWY6E3DhcHAONnc0sxsJX3ZtqAvSFNJZ015KYHcQentPWVJR06dDnj
aBvIA/C8cGANvU0Cyr2Do4/VSKi14Plt3hpIseVSUHaqr+p3OtFOf8gcfS1PUMqX
S0izyXn8LYhuYIsl5r4stYOPSWSX2pfASp/wd1tz0prgZB3cayKVmKpAMCT4xTzS
2TJObQSzj2NQcA1ZtDhcxas7bZNpDlgNByptCPgpCpqut1M9Z4vTKMAzOktGKxyo
4NDEpoapW8pkDvqfvbmzI3qk+TMoFgXpXu5zubFrTWyu0VSxC+uycGunaSi2Vope
9qvCfWtIT0z6a8xtdLURRvkUHasx/zfGL46ZSBPNda69H1KQTtHDWTGw2xtRL2zX
o7log7iPRNdmjsoR0LMCd/4sw1yk1GA6stJy25zioK1B1wMV6ioicUN7YrR8AtTu
59i0FnGoSoYx3SUQjZMRxHKv8hlmHg6haPkxQXdRmTsgUeo3qAT9p7uVYSxCj3HZ
EwmphMdQN/pnch0K9Zn8MD+rvQKy2yiGg2W13DBEF+C4f0u9bKVgrFZjLf5hW9VR
d5S5Pe5porqEVPGUYggxsRKGTn8Eg8UgPrewqOpIl/dDQeGWHaZkcTfO3eehocvy
qcsjeQBJSUYyvSdFcSpMlBxGBIqlCx6CbuHWKO40sVU8ti0MUovtx/v4TivGcoV9
ZJC/3fNe7LgJgnUFYY9tTGc5B8S9eOmlQSYhjLz6BSZum+VQBJcf2/+V1IIwW1m2
7KaHwlc2p4Dl7KcSvKb7xsd4AEV4omlHQ9tKOLnOLsZX0oHCrA/rhM0ouyNyf1rG
ygMgUYlFYBWCH6IQn3s0ptBOVol8wu/8YF0qh0MI/2oSMQg370ckDvh0HT0cghCy
wmhzubBZ2cVzq+iY2WaFzciPzqf9ZInkmRPfI67lNJqBDYKkAf8tY02o8Lux0D05
iDsyEkdWNsXhe5tLc3kfSGwJ8piJb1O+XmdZppVVS2TJZg6sl+uk+ytcL948Lkiu
NfIlwDHNe/THalGpWp4gN976l6EXIjLjofDyq8Me+W5z1LnfEjzPOA5fKHcOpHy9
aSra0cGLSGXTOYA/v92GG1skLDwhA6iOO0I9QoaERMPrkUZhHMVrOPZMxE9kW8E6
XhLv/KO+uIU/uMjAaAW1SGXVz7jLPdhuoxw1dgmKtLp0QtsI1EnV/ii65KZJztIW
ANoUFfB5aDlWUHIu/Nw0u/r/sdoChf9TjsFYpbyQwLmAH0Va3E64Sim6sSUG1Afd
ZCGHqzdvXwmaWuO4Sgsgf1uaC2PyYB/ySQ9hGsPpwabpCvAE/jcVqQQ0Dr6Rh5vn
uVzRzxGpe6R5eL78rbL4L4YaJc7ciQFvZ2ogFWCIZyGjQ/OdgXT92pafSc9QuvmB
u5rXhPevkBdCB7Z7K4vCD0qCEkJPuFAF0o1vhoy1gTwRwejDA9VBqSwwLCNaZtvP
t4o8tuJIy4tbA07MZhuWH8CzHnUL7YXyPpv1OCFxgS7ZbQK4zpPpXVNgd+7/+tLy
ImgVCrFqGLVFgfR8iHuFOXC97jqynB+ZpYdQgDBgepz47hVW9zwmGAqrZKVnnMqy
1P5E+ibuDHdxixYgJcT9o3Moc5+9yzbgquBiGzy8RRJdkoOlo4xg5awWvbocfiIW
wJJbNtT3rdfn5NIijcwLuEd1a9Dpwt9aa8UdzjJG3AX2sR/jdx+ksOTxL3mynAoH
G2/uzykhPsXUSDDQvW6bG5mH1L3dE8olSB+asg2m0/ZGH1qEFrI1PbCg/rpyXmtG
idRzBtX35LmPqusTitX1N9GMA/EEzPBRcBhNjZenIdoTTQsA7yIeWSXYeoUnaxbm
S4FjIs7sGZXyhZGhzx88BWd1F+zDwlrAij3w5mAUM9i57c3M/5yu+nx8eFkuqLLG
PNmgraQnvU/EJueDlmXIXa7WtB3+I7yqcP2tGk4p3ht6R7XT5Nnf0O7yjJXWBNrW
obautcQrmGaCUhK8DvJLwzatDufSolUKR44bbJcE+R0/bYmF4JkQf1rJLbXpIBzz
tAxRTR+mQBqOn7iUrIHtI+MajMzinU9x7RGeBVWhD/8FS0WwRM8iAGR9DhQJN09q
Q0ZNtw0ZGLOVtKcMU63NUn8iat6pKjAZQsjGn6WN1qvMLg08kSYovhseubHKM53o
qIKjDqBMcZLuE+bO0qo0iVOpTON0vWeBKwlICZd3rbjFb2A4aTFz6FxLgwKYctGf
EEmPSs8o4pjVxgfVJV3COv1YQ+3HacvoO3n7Rs1EqxbzXCgUWVlh8OM9i9N+1InL
ZOirEdlLOsQRDWg3+qKUnGMV/1Ybc+Pn/R0M1frGcNQNDDxrqCBDxQY+E8m4WC0S
qSFaEDdko20e6tTabZPNP27VDCEoO8rHkrtQheuK5L4dhF7JcTCxgszIHGED1ACr
f3vR0Hy3FTceycWVXjQp80R32k2mr6FhJNdQFUOIfxbzp+ZgDPrXzzmEH9aTNbmK
elHndhqKQPywXVMyFzvw28+HhP4HRdG43Lw0aAQgqaMLuEhCteBfl9MeV0mBa39U
2TibxkzpXSkyiJ86Nebj3hkIh4vYEXVq8nQDI6opsP1l3i8bwZr/ogrvz9plydeW
30ltAhiEhlsKZ9q+zTaKveHj5pghwuUoyXyFg0mHOfcmVDEvO0lhxGv2aogXB4di
LRVav2fxQYzUkO6v1fNw4Om9OfNk8qwnbGKjfXc4RL+SVP+sjVCLXh2dZ6zsZjfW
z2V1m50cldwPYdbtGU3g6HLWqMi3uQrJllORvZ4S0wKXr3VYOb1Yw5v9qMbSCvCi
1JENRgI5GJXF8KcmfeCT6K7XCY8sM8jXgftL1wVb5F63AveyiWkUY3E2CpcSw3kd
mb8GnMgCy1YTjQ30Q5jWZsHlXrmrkbzHLurjM5SQCE1b1Tl8uXxlAY2iraUUmn1u
fA5fDGi419kf7/0KZxdkqTlw8KPVCdEFunGmXo94QbQZeFDQEXwIdAKMyMxnwRlA
vXcDL3szhYrdXGwQHD1kArbwDLFnpNAhLQFnIr0i/EgLGHLnHTI1l0Czu5mPEm9w
JNRvNl/7ro1+Qj/dIcToE/hVv71rkmME0sdnl58cgIBKOxfKJGZpP85mYjfFbUOJ
hT/YXtH/D23M6lLv0jUOyCYTBY0GKdM1JgMUw8m2kmGobygkJLAp9EZV168vypH+
6Ytj9B8hS9GyEUmHYlayf+uRAk27j5vAqqzEh1BFpb7IjxFS8un9rnhWxOZ79Oos
76gaC+b2sRWD3zicZ0u7lOSRHFTBKgSJTSZiH2HqH5b2IZAO/hW9SgDs0naiM0Qd
MuDggMcSWxdPV9IkIP+Ko0AYuh65gyKcCfpfQ+/p/01s1eIIaLyBBl/d6xfkIMwS
G6DjeQ9GChwPcRTuMXvtjcjZ49GeuLeKjJl/c4jSJOhwSO0rVm/+0nov59+qlblH
q8/ewfd1xuoi6CscVmPjSqyHTdv2Xv3soavga6jgMp+s8GEoJ5a1479AdcKsRN1a
krwU3Vjg+T7fBtn++NNd5EZGGXQcpHoY9clvGWvqcmhFZ9ZtP5ULkLiaej9CBXuK
GJwj7NtfOaKYLhhiR713d/3l/zVejjXwLAyuCVwRVkGwedXOUsmJqfzFK+5N9HGi
+8Xo18pGKspOjbLy12WZ/907xlNCXkFig+yQSYx8tsyPw59f7mrIqhk8gw4BKnWP
VM5Doa1qWghR3psIj0iBtBUS+qOwznYaYXvF/0pLujrwsrqvMg6ukfsErUSfmIQR
C6Ozp5M1/1qUicIIOwixKQo2F5M9p4wZEzW4GhdgLDVEt4ZmgFtuRJCVNPeapHcI
zEM2h1gUKXQK/WPs/DR6/vB+O1APBfyeIypzKp3oD782AD4IbIvPjEsIePc9knno
X1RaSSik8LUoymhN5pGMEr2a9sfIDYqV/elfjWKG4M/m2FaDnh9TADUWWpTtTwju
qcBVtIrajdVBYSMNwNUhf9vHnn9TvBHVwMAQHtO/DN74G3lRcni0mI4uTqun8z+M
5gverP0wC5kHb/z+ptjtWwUW7XrYqF/Oq9DG5bCga46vq2oUZahVKnTssIzEpHEb
OggGKEVKLbwGT9ilwqra4i4nw+//o/HH7bGgzA8oXUI7syTBPrN8eXwvde8+itWC
a7B9XY2dEEBUrI8N2zsI07EJ5oYErzoHblLl1O69CJ/tPbZySJvFi1uZIRTl0NwC
MllTCr9ISew2Vje6/StyiznO80KKGF5wiqrjb2S3jd4xSzLjgaKhQoL9nIsFN8Yq
r18Z9feJMIT7fpzE9WW7p7O114TOWx3lPXsYvFWXvST1oUcwOBvsYhQA42I64P4D
KRzDy5X58CNFZnDwh5P1Az5Mwh4VB+ztO+5Td9aPvHusRfEJ3j9126Y2z0TFOADx
2Jj5+oKMleSidBVd+Tjue/yBT9MCSNJJIPQBZ4VS294rxhLA/eWDZNUm/PiJN5oj
OC4mIUg0uaiV0VN8b2dhMICnT7KW3E1rDfj8ei+903iWIIsR1/lZx8WPAzbjj8hh
zBz5ZY/h+d4y/X/eUJngSeHRCkMuC266l9fA/2e/MtsdY/zvkKmQW+sJl99l3Ch0
ECvTPv+eN+FEkAyJAxLNbzQMgmLxNLYzDY/1sQinIgg5YHxVM4mHUchAfprQT1HZ
hLonn8qAb+/NuM07veMAv6HOLaqrFpSGL6FvJS/b94+DXllaj6+O56mR9MyU9m+r
gzXyyQ6fGooRZXGcT/ZPFLgRkyCs4Ij4G5B2iP2fYvbOcwc9CkqgomO56ejvEwww
WZ3Q5P3nxbmQTpMQKNlkaEcdgRGBUHLhUgEZ2VTCR0028K94eUpMpocq+aw+zpSs
x5DonOPX3lK1i8BXk4zI8A/q2ZWRSm2uz8fSO2pYBlsHAsiYOWDSpjf2s0a6e2F8
OB9fQOZ4K1BSnB0YStgeCb9oMVbgnuBoVJrZK5dMAhL35hh8/2YlCy1OOSTMYPmm
Hd9qkSI8kU28iwFR3zcyubkbFycUhNYbBpIitoyaKjVI64uDJ1qKFLMcEn8it79j
apXzjMTXevQyGs7MUOHwYyUZALgbPx11g6nkkS3rD2mA9Mgc8Tw0suHy8kwPhSbO
l2WZyijPchFUp1Umc8zQ6jjql1zZ2E4DKxhEWtFZm9oQHTN8iZoUrSugFBTzPDsg
6VWeNrORLSzP67kliUAJts9M71nioXlKeH3sUAYjrL9+tHnnopv7mmJBKo1mILfe
/15RUj5C6HLS3FnQiVIGjBiUv0RhFeECWllpWOybJLJudBppFbEHGulUSrK7FAUa
FnEbyvzNddUN2tiIBAxpD2uvjkStDQ5zRGfBw2r0j2lD+KjrGfXzckhdO+QJ+rgK
hQxRJaB7UUr/4CUBxPuJ4bMwOoTvVA7Y7EF9Xe7H2HPwne7o0NGIlNLF6oC7S6qR
mXkANzN1yLBwMlLNQfLuAN90yVGm0/fXNiZuKghXgWd5rCptEp08Nhy/64gkH+L5
4EmQ5FZ5DcGUfNDi6YfB2BjbJQevs3x461MmC9x5zmRzlLHDwIxcl+qzXfh/VMfT
/HTiy95QUVMLXv4nYSHJRKX6Jf3wR4CA4KxuAb6DREolPSp+lZwYv/jR5YXkGyqo
tm+FDJRuJMMIvO1Qj5sh06bRvVIAjks5tZ0852AlsLQCEqBI0gU2BeVwYxnUTitO
sCYVALRDeXzU4kfslxr1M7eyRSJs/t5g7hw0bboeBCYC+jeVCznSzzNZYj/mE8FV
9ly4bapyIhpwNwmgE5kWOrVw757sCAFMHlUF+/iIvZJnZp1/hdK5RjRktocA9hxC
beI302M8gImH/76NpDWY1mSfPfDB+36ZG33Z+UT6n6xhl8caRGIalG0ZH2m+TB2e
8Oupgc/+LWnltcia0VrIGmJgOQfuihls6cw1ZKrK96ppSLqy8Yp+lzGchQLr/q3c
EWEi1Ih0iY+a0kCouJ64QGDjIxlhHo/dYuu7T9ej3weOe+28Iw8Pjs1G39YCfma3
Lht59Bq/052Vi+PqXpHWEBbaXN1AM8KScPJmkl7Gi0khBQkfEEqd7ib9Fk/ZkTL7
m5M35QOnNvKcvj1rQOt2lFdLA2Ci9FKfV+jKvblR5axY3fRg1Uhhce51bXjuvP1i
2iNSd+Ry4QzZCV3UjepbJhZXAQ9NYDpksBXQ7X+Nuqjr5qoGf1EC8rimQJIbtKhs
Q90J8Ek/22IR/lRaY1dxKEV8IyVKGgKDmDh6tgHLTsXXoWqaXp42PcxOttDNVa1C
QIQVvywibuLAwTolAo3YphdeqJCUpw2e1OK5u4u3FjEHkT3ATTdHF1v33gf4v82d
BtAdIbd2hRXKXARI/VVfBECxjX9WQFjyKPm8cr5vSN0237hf2OtLHbmdY5ND1uMf
lZ9CL3rFMMTC8LjqUCdzf9SnAydn4uf7/5d/MbPykjiiphKLd4a7SGCY+Bwaj7Yp
TOGzu4FinJgv9Typi6b2acK4LjBN9L7lU235yIOKP0LZcU0fx31vFuv5bSPWMiQX
ftR8Yyxct8dsWrBvVndyausXw9T7u6BX1fv3Zg3X2chwVVCZHnWdjRphc9kDfWpo
a9s/Jug2h49WXXQth+FJ6m6joLGEZvpwvKLUoxpoXyh9jdDSO54FRlcFVFRErp2p
1Gxp0K4n4BqsskFoJS8fY0PH09AkBjIrNSHmmGqg3k4dXpI2a+aZEkZ+yL23VHKR
q4sgfNzOo3QShfuzkbg1HIYrB/MWF6O/9bzbVy7K3jeyrQ63YC9qibpjhYQuFA3b
2Pxtmkrl96Mc2SAK9uVaDNPfjHQPwLaSl/3kXsKmr2N4qynI5XhiQWuADS9Jba+6
uTVAcnvE7Lh5qCuPlrxm+eM2ZXdOZL/s8X3Dl5pNZJPKzoEF9XAKIdpwdvaA+Q46
Em6KiLfKVCSsLnSc3B9fRWO9408vBt6KB38jRsVSasQmGTJmi6snNb8JaXMvUeXX
EesMDY2ovW9iYT2TSB9X/YWtHA6F/ZFddPw3UAEDhYBT/0cO9cNwgOZ5KjzTlWL5
VupupYvjYusS1Y874CGbCCIfvsZaEMm1q4z5GbXOVUSRrOp4mGuCmpI8yWcflkiY
NXDwD/ZbK8ZeEJ2Y5bT/QZHN864vqVghWs83anBxirPuKBznlSOFAKciZhCwQnO+
omefz9ialn7BTSkXpsAQRQRga9COgmAD/Vcy96CcDdguB2+Ie3T25gN1Luf7htSF
8N5j1FF3Uvuj630kp5EQXlccTGDm+ApQvGhajNt35VyTMPqGeAOjb4oGxxYbW8d9
xoCR5sXJewi/RbjhVQ6ZjZ3je2nJCx76Vrx6ogl591H4WPSodvJQvApq0yxr39RN
MInj2cB9ZVZJNkJ5AoODVj8QGgmniGS5/fgCLRPgeWpgzYgKAgVe0vdTVUlkHGdW
+ovxTuGJ1gYmFEfMVdPi+YjfzbZMVpO5qaswBkGqOeBD+9O4TMDl2yT/GEluFAFO
NoEAurvh9N0a+QNtRe4Nzzbbyrr3v3cXCE1v8UYF/v6zO9rDxORKi32WhGDK21cX
X3t2Ix5CoAIrsNmZT99r2nhTrxZrXWhbGPLBGLmwljIddth6NDXTF9UUcJNXAf65
uhsrD6d6CvG7vsZQTNYB6aNsgusqsY+sWeaZe8Xvca1dNo3jwskdfqLCiTA+ec+r
oKDHI0yjRqzBBpOe/1zAFSYQ5uxPImd9n1KS0LFG4byolMGbldQTLVRDZJH5qrGF
f4zDN8V2REXM+b+0awSJg1206wUFoeFvZjNPOwgu4DOyOAakEwbjz/h4ME48T6Kt
yjci9AeNPkCwCLSH4P00uc38jY4jO2Z2vMMNvkq0mY/uh6PL/MVGnbF+ePu5Z9Nx
KjXe9wgChTXLSOmL8f2sKwdebsIyYj4Bt1K2uKFNTfKdkqXxV8a342+zY7DDU0OV
ILvPRq6iiRTeI/T3h+u0ENjlf8b2BXPLVsav2WR99zXbAoRuAFIGEg1ghgCu2Tff
1cTZR2Hfr+FUpcdnrytGwTHDAYZczlDymKTkUTMNz2eb+O/OqXJlBFr3E4xDGh5V
7pA595GFEllid4ajIGuCDZj0eZQeN7CcITEtLJBOA8sP0pmLhOoPm4kIHXfPPP8r
OEkLq1puEd7mvLOyfobDHbSj/6NgKS8DCdMFSsszWlzZKy303ZluWJlJDcFI22bF
qkVCmE8iVm0PD900ZdvoSc9ESSTPTBrFB2GgZSPh6Sx591tuDyHPO502eZdLwJB1
SuDFr2UEha8554vzTp0lgMQwb/SFIF9dphdhAHdDmzfcAMNlHGukw6yaMAVux/aK
q7tZLWB4wZSvXrMt0L+4YdauH4uTw/Blz0ULpdujKR1NOX8mBGdOD5jq3Nc1v4gi
NSvPpRBA837fv1sho0zOTZfUev9B/sXd0gNa7eNLkTtbjqpSoe6BUaJPBAeQ5czD
dMKbP4cYX+/Ibgz2eYZC7GCRLXV3TazqSIh/KzqM8k4LSkwoIpbAEk9WGfYJ2atP
FG6ISBadAOgSs89ND2EvPQGfQ17BFCB3EZecD8k4Delq0FegmfEf8ycAIng15Qbz
J2G52XhHQ+CIcMLKZGqzJxCieDuVlRQWD1XYep4puMOFLENpcI4dlM3MaGveXhzI
XZLEQ+1391ZCMvJ/sm3MBUfNZqCVY476+ZMninJh0R7Gh4F+TUzAb7NB5t0q1Hyh
T4kaSeEa68OUYvqtY2I7hU7jeoc+AMj2CC0dkw+td4Hj1FJzKihlVycTS8w3Dl1b
XP4coZZXV49aohAprzJmEh8YbkRp93HIeTuia+j27No6E9ws1GbicLNadC6GQMW5
ucM/Zuro3/Tlx6O1aIz6MfQgxwjiFaOenhc0KE7h0pEguLk6TwT75roU4L6ScArW
cg7kUPpvm0j2IQcwrUPKRQW4+lZ9/V05S0pXt3rJLInlHGRNr+PEQR3ZkxkzhL/e
cSakZyjLAn4lRFi6cVTrZ23dC21Det8gmXCB0mdP7dL3Mb0oW5V4/hgm4xsOr0BQ
DzaXOoN2kho0wnW1DKRPaZ8h+/Xah383JzJZ0zLIibtKX8q+XeE6FwPW4K5bODAi
Z61tu81zvFl89m7RK4a2Dj4+bTSj5Tw1tp+3Y2YkPd181yCIKAX/0TB1NnqhJQk3
p5RUDlLgZAAZRox+SqXwYAd5xm6DuC+xB08MnZ+WBmkSES08Wk+LxUTrbumJRwju
tl6lA9G9wSWhdrou4beJwEWrjeHJtP5cijcSDXMPK/lf27GTJW3hd6OExZfcR2Z4
+NmUJ0B1fpIt7PzwnPdlGq6/9Wf2olZl/CRZazaJhnIQz6FJkBNuesTjPm0MslUA
waJ55sOy4edR3JKMr2LKb8U5xkxZGNgoq077/fJuDVCDUZw/MVMzCNTqtPBI2yF6
yJyyQIr7zh6NXi3UDpIicytrafKPha7foVuuA09m8sEXc6w5kL62aHWy4IgXqpfN
p93zvvMad+eQttGKoJr0VrWM4IndlrcTogCK8spg9aBNCY7jVQqP4deQNUXIOGwO
xzSafjDFGd5p/dpg0pHVY0DfQxsJEyza0cYYXnMz2GjOUxAhRyf2hpJJqs1WMpMK
GeNdxFtMKrkD7rJ1QPMCpEh0H/ctIXu/aQX9quREvlYcfP7xbiKdiCj6dvRQz3FH
ZxWLuvPht5tnjwuqPttG2C+yWxojK4kRcGdUzD0nGH3ku3nFH4m+JR9AtN0XOUrR
HONLUZYgjJY/qgsT8WcCnheEut5xhkAaevx2HRYtXzv7oUjNXZ15tteoqwSD32ew
55GHzApepmbi4iO1TAnlZl10VPcHffbjKwnZgH71M954dGmxbb8He6bOkhqreGbI
tNX3eoukjASMcrAFibppPpz0DciuSMd8MhPY0P1pdwtXX8Qt/yXokdVsXzADi6Ot
K6w6TDSzeULs9+I7gytPGqr89xCmFCm7t4P0AzqJGkORZQ7nVrYsJUql29DnCOTK
KXAynvogQzQ+cCqT6msU43y+CrC7dIQ72NxI6w27ER9iQGfzRgxd5IcghSH4/4+m
4RNg7AINRCnjZtkN6nS/KdqBV/9PxjmZLcs8NoO1QPFTXcf1+2qLPghj0LgKLMXD
g5/YvN1JEpSWG1LPgb2STNx8+Crm/Gfni7tvZ6MBFcNy9TayLPbjg+dfnJ+mORju
HHWWvOOcHVjvu1IZzFmqCbGWojdjJoyGqSya9nmFtUR9u6JvXm/wTElE1jIWHxHL
cDQDPC3eqqFvln32C6M5LqW2fn6eNsMux5gHepypeT4lES4roAmKci9dCTviPdUf
0mjkT2ortOpThszdbzu+LDQv0iamulNVEDFOqxTZp/A8ML+Sw8NhBiLSAP+sW/Yj
JRmidOT1h/tYLJ6G1fMxs2CdQ1690rm4FXLzfODsC5/AnZ+iobsgwLOyeY8J7mnA
eZYM57vpAhBT5Pw+FpzOT3A9ZDalYLOzaV2/GXyvInLsONzCe8vWE+XobWryzTRr
qn/1eoKe9pmfCrOgb9lVBAQ8G69sDnX39QQ/sXe0WjG05Y2R8GSChQtkgaLUD/xw
jzb7u3Yxdh8fWUbZINd1SoI7w4QD4SDSoc8B8WriyRdHspXWXkdPyyuJ9dioPidH
hQZdzaMtEN28pH3bWbUD1IVB/GcHI9cKAYlv2yUsngZa9BDo7Ma4Ck1L0JhAxaZ9
BthfbP8uFX6NaK49zCVxatCNxLLSSbf1zf1fYU7VHGmAyHISqrOLQRmhSJ0a/PUJ
qpmcpz1Ph7OpKcGLGzWNqzlsprYKCokkOuEXth8sqwYDXGUnEp9zz10db34h0qf0
zbzGdF04xgEOvtBx6yNuSDq2xiZRymwxn2a68btkKY8VjxBiJmb+KCjTUkxRGcP3
Q1cu5sPpws594tKcCR9xme/IkvQ5o7d5JUClUP3JaE/zP6SZytn2XVG6qyUDSGBC
cf9HmZYN/2iT1Q7DwtQ9K65y0pwt8dnhHT/xKNwUYm9Aw6FQaJb4TYhg90KMZ6Wg
ZsOHrvlRrH5aWZpQnzeEGMNWPDIcFekalnV8ksZbsao4qsc8OnORsVatq9nGZB++
VvaUWT3dbx7E6Izh/7iTtjvE4rBnJMOEhkpS6phxA4NyPz90+ItC8Q/VB8WHiGMD
W9PZ2Msp4LjZExrkBtEiYtnlfX/0iTGMnXg8ufvyqw+9aYQOuBfX8blKBYA8s31g
f8Id/D1exm8wIkqNnEf8Orhr/kEDmoScVD6gogBYdFi9iARmAjqjkXg3ylqDRvCy
2FIGp5mRpZpzfDTEhe00DkMXmZ3xfGUPK3lDL3FSiJJMZPRXQtgAWiofgJJK/fFu
XN0pu1fjolOJT/jaHSq8VN4ug4NixugGZPiUj7ihs7hKADp/CWLKsKyeRBCZU5Bf
EBu6KTeZRdnLr9oPnV30A2c2fqAvFvP2vUF2qVpXfFSEMWiX/R67s5DaE8zcGcFh
6sIIIvf1e8CHyjgD8sVnLOwEhzZP70wOxpd/UWpnWz+/+wLs3JaNtaMBhPGVV5yY
brtHU3u1cjFHfHEsICobups2Sx0LJOEH54EDGsWfECPkmwfk+Dt1KNJmMmE+fn31
cLzrzfaQIeSJBbvGE4vYHrZCWD9ER8E/n6qQBIWEbzIaMKBTWUORQwGWMUl+B066
2aIVjFWk3go4ejQp4jCUOOoX6QbwlKaKnAZ/KJugkgI+asqKXj7IcS0BEjHZE3I/
e+z3dkDDY4cpx7qLUF3CXBhR5aAOd6XsHc8EeGVr17++zN1pyzn7T0wSRY6AG5or
LvT0C5aU39abi8cOLqFm94vucW/qDvwmk2LPnnZrsK6FE+qm8VW7YHvEGXR1keYK
UN4EVipB5PVlRDArbm4eg6GaLCDty/ctFw2btp+LhxHk6xBa2I3ClelOkdFCJjrG
aJxC+GoWXVk2darCjB4mLhOPP2D1qEL4smhtT1jFYnvUkwLeXx+a39PwjlcYMiUA
LVFDz4UVDJz7PCj6W6Zj6cG2+8wDARkb9rJX2ydqn6mhff8uJEZeIQKyyp1CoS4x
80AmxKSPm5HJvUigMOvnw9JILmeGNDe/TCUBuDcfF0oAhJMAKo3hsKDfN8M96Grh
vDKSqoLVqOhikKXkfXAurC8Hjl71XLkOV2NewshTAYXCUQyl5XhtCa+SapdclXHf
1RaIA2onwc7w8EXgQ68X8moTNhgTQrx0GX7qI7wsRJQ2nsKEOHrMfhg3ZfPddZSo
+mpoc38lW+5pUCZplJ0+oMacRxxes5czRTjmkHOnWdy+weDnmE8kdeIsM3x6kHfR
Bb3uvdwDjZKZLFVDxA+I2rF361WxZLPgpOIk0smbQ8GgRVsA3uji5rvmd/1UsQ2g
PYzubA6izw7uGK2umiLz4VpKw0ozEQlgi8+m2GCjRdq4J8yMcg2WotdpxgROtM0C
n1+aIz+8759XwTSoDdQkJ7RB6ESiqcy6x9tdhkXGm6842eduoBrFqHhGw1vNngp1
KAuJTmbCjCd0l1RiLzL+eiuk8NVTdEgnvJ6zYKzHYSvkh46vrOpQjaqwrbICtyqn
fudTXmUe3ebMnMyqVurpZpA1rulYENIuSmvTfq3ysQARaMWCfbDSYceIGbWxAtTU
sZ6pQB6i69YMnZ63H7OT9LJCThRSDhiN7bCpRKckHw/jEk3QjAErnKRM8oui+7z3
CoCwCeoKkVv96UAcHgbdz7jW1D99LtoaJ3xs4bvD2un2Ojp1yJK90JCQQxSuMPTi
YdHt86iZFELznjtxxnTSMUjrS56iVfxMeKGMpu6rKEVn6H9s23/0Iuz8gmuBsmx0
EezBL/cb0G593L+DQWlNCoV4DEMmVBJFbM5sm0eXQjZ4ln3Z0PPL5Tqp8Q1ab1MX
DF2hbus3Rkp2NQJC1WhHa4RmbcYhvx2gvthkbGHKebVWnXRaVeS8GD061AnvRXJk
j4kTd8ndwnPuIpwX6xg49o6ykb6jKokOydx6aY/A68zMYonQdEZB8oSbA9zjRTKc
IkCi32C6oOkZNkp77I92LOImg1BEd1PeO02JrD5kKq91fc+zplFrXGopGR7YtIiS
10RoxWweErvPEsBt3IwD8Eqv0bA0jUx/C98FM++ELrp1sKheI5fd5eOaVu45FWZz
i/adr1XHeCvRV7TjT1nHAy/SnEB1A3gyGPp+2O5VVCKxxYKYy9OWGO1rd0a541jF
9nU7dd5BhSEELtDRXD8lsd6aDCUqNavY6jHbasOvDfcJ/UOe/jUXgQMuKxYf+XwS
rVADz5zaQdDugQm6F6ubGFi7RXqBWUAs3mzMyiVrq+cxYLIIQqmJ/q9OgAnzGTQU
RoAClFdc2Ql8vyLIogdCqgmJR/7qry71tj8HeGWjcibaCxKThg3KYTPaka6sw95n
rXh/qTQQog0ky0BsSUk9OWrEpoTMlA6OkO/9IPpuUH98SzGU/J+NRl/pq5MzpEkq
ZB4jrV19JHNXfHNny5eIpcVFaBnCk0wSV1EIzdEpXC7+VqPaa1RzqRAN1HQUqP5d
09TiCbJJEccDImWLG7ggPk3c0SzMZoIj7zRnDYX/gvpmB/jRfAQELUD8NQ/KsPLd
P/+3uFOUaH6ueQebZdambivgjLABuCkEZ4mG45Vfd0Z3wMZ22KjIwKrlm+0HN1e8
6ySN4BznwzHrLLVztgnccR8JjWsNiZqnb+UBDqroeEnUkhC5v/tJtYj5XzCDyB25
oyOCVvGiTQx0dJu0iPD4UxQEXTmMoVtz3vE064yy2QEjjp8mmZkZ+ZSQKSVag0me
pqqjCDrS/DvBeHEJIbtHjec3lVRIk2S/W6SeLZjUWNQIUoCk6Qx2S21zYLvlswwV
/oe6n8+I1n5em/Ntqp+OOsc7pUrX+FruL0kuA1Xd3l2jvbZVMlw2gQjXOPiM2EtS
OUBMFYeW52l0uiuuvEpJn8YyAFlQWb0X5QR1TYTtBvSNq0ayVIjXl1HSGgesY3AN
H/HePfkIdOHGjj4RF3ChjHTWAAxdaM9No1+EQf9/JQe+vZtKTTE5YJc7KdelvZ5J
WSXbNPYoL8qJST1g3Zkt7/PSPOchiqhCmdmgw6NuHTm2mqhwsVsn071k/1AVmCxp
NnuNlyF69T22UKBs4iEXwiXd/02nct4YMDayovfZL7q2VtGzIEL42MlkIJIpVN+g
BHFkfaarbbQsjbsS15VfvZHd4uGOlALlmFJwXMrSXCO+Q/L8Z3/2/hzVqTMhKdQ4
pwY7QVxEyQ6PGemgtrozcEwR7imn4Kqpq23E4xqofFV9sQsi5qx5rvWmgomSrvVh
A6+bLDL3i/BaNb1+Z15WziDqQ88Z5x/CMGAaZD0rJdyIuDqFTchndXA7foj40I6o
YNDN2R2MT1Sj3uZgFFy6hHjwcAzpKiuJOXmFPrPH4LqQwOsmPGGnLw49qEaEMyi+
rFaqMlsdRpr20KCzmqY+bF+0F29fCXr7XjVSzQnBvjYFq2SzYr50WfaS9K/iI2dQ
/rvaXpJcADTHKjXLACDqp8tcZLsuSKoHGnGwippOVzXbzfJj7tE3KSbGNHy4JGfy
ZyOBIVDYCWYUXQrsdOyn3i2aTM8hW/aadqDOSC5Sh72g5mSogwf8GWdZJiBXrEjz
pOb/jmAy/xB0GHIHS26KtJ51idm84ISiv8t1HYa102Ksxi4fHqVMXPwyOiSv+1ki
swVhVqQht3eFIbJkwucTjlZG+4+J2wUPvkNxqslo0aUMm7npxekc+pE6wy5TrnWE
FSHdN6tF9UNS8AgTGSmdKUai/lAWdTW4Mioxw99kKS4U/SoXd9jgzSSpjuIGdGIw
Kk+pusVJNx9br88RIXJtdEmymH3eOvDhGRXVtRi5W6goAoEdVdcK+6mI8i/FzYHf
xliM8x3IIDpvh3td1b5hT+/ZwI063DfObQe0rvjD/Zp/Wvl5aqnfYs4aaf0RQ4yL
RryYkfcADH86CWdEVjmFwdxBojTMxfXFb5GQfo83jYV/XYO+J2k7Zn36miETxkN7
G+/ZYESLcO5Wk9dtwQEckzLQAk0tEjHXBZw+by7INAUnaeyMt1M0l64l395ccD1x
1lx28W4nDWnRcVrVHXi3A5cCVk1onFr2cKYCZM6up/RiXNxPL6lAe/I2m5wHMykB
pwzpqBSuCHKh/OtXW/xw+hbAuQB5UtZrIKgqzbbP8GXlDa3VpqRAxCA02kBZsN2C
6AqR7kSbD3r9IwSBqBYs/NXphO5g5za7DF1iYte07qZNiaHVoSwf+BXu/vlRVhfF
9SfQnprIsK/4CNsRFHb04ManLd809UYlbT0fLlx6xtoeGzKM5mUmbmPnvuR3N37p
5NuAjBbHwA13wyQyQuMJFdtPvLO4hObWDFGR0Qcy2lmGP3JX0jJ+gHEYEJWerk/F
wYJo7g/VGo1+/gW4MtJ/tVo4GqTN5oHUbSzumASODf4+HnvkD7/ETxXsqyYuZG5p
I/o7CDgaV4331XzdH1yZ9TLfVG6bTzDB46ULQf3C0KX6iuA+xdlfB9L3Kw49X89D
MPI0svhs2scBIQRamzvNCeB2dfV67+Tk0LS3meE01AMQlz+Gs1OwKsS+R68CV1Zy
/gbLiiEqlkSQR017MAsykvUOECvcw7RvwX/mQakPur/eadh+Fck0cktWS9IMMi1l
DopbPzi4pvhz4rPoeUViOAHAl7U4p1D8R+g70vUT+gUfZtgL+/E1fsceUkx3SmwI
teJoFmjkxUxSsHywxikvS31TUtshqINC7CSx181i2hE0m+++Ddet5ZRv+fheYUl/
USrP3fZYJYY7nzRuSFV262Tv42P6M9Ihygg/F+diJ6m4Vp8qWPyaG6YhJ7pyKulc
u6Dl0xkybz8qI/JZ5LHGz+siHbXrUuyX4Y+pxtMANTQOYR+CdRxYD7+LthkgxVLV
xF9Uxf6d0RBYom0RRuOZCj1lUqUt/q3aPav2keVToLAAVMB8Zd0TOaWsF5CCBl+b
H+B+Td2Skn1tUacuIf7pdnWS8KOJ9jhgADB0U21gauhueQG3tdjj/GwO1XbL/mKw
7cuHeFBacOZbMybGF40Z6j4TnJFetlKLq3a9zjebpCYfA2k93Ukukb8eFxvKwxTH
ecbmsdM0YgQ2fQfaB6wSBBDx7IbI5zarsUVign0uzfDpyegF6jhe443nu+AKMIzB
inSdruUDS9GZQoYDnmpNTxD5Pf3A1XRiS4mhzLQioW3Qn/zc4buG9tfbj2MFifM1
z3MkBkV7lIUQS/zVW1RXyBtj9QyiXAJABHb7zuO996O3ApMHtrAIhlmhreQbGy+7
hFqb0W4+BI4kFZu8vqEq+sDoN6M1Qgz//MRnbrvVKxIOAVyWKeZE/F2cfRTyPh54
xbcSXHdfe9Z/aUKox60pNzWtmLFLnpT//NS+sttzh/WPPA4ycR/ZrrJ7ZrdZX7n0
Jlnu/2jKti3tPtUVk4lHbs9W/HKsE6Zk+5cT+AZTKvG0g9jofeq/Q+XHFvHfWOc6
xyVXeSkXZT134w4YV1s42pgLsvrP9qDlp93DWaXN2/POAM8JbikoPlDOBtcEk7ti
xwpye+w9njLkF5qQ100SCZUCe4pTwIrBQ+B68IeGxPRwgICVETO+lY2Xdi1GY5HH
JnzctltqN6hNBPnJ2trp/BQjAejyzYk/hc1ivyX6OfHoIGYV9sN1hTtdwaPKOyfP
B8Sro8vEmbU1Mg5wd8qbBF+WcC7nUYX4EBfe1zZq4NBIwLDTZK9DZ07kw5KDTF9j
ughayPnDIGUq08trth6HZtBziQ64kpSSCTbKwMqb83FQWXnIz1bLbI3/H6KCyteU
/facBqMKxCDXO9p639B/CBi8MxliuRcqg5MNve8BHiE6pX5YlZmznYYdLwevQnlG
xOcq79atdD0prjrv+BLLAd0rIClozsQlRgQdtCh3OI+OuknFyb94B3TatPx2hbqD
h0MxJlGSEaE0/r9B3Hq24Ueox32QO5VbRIVCH+xoXFSugDoQAA7s/m2kAZiWEYTk
9QEUF9IXbwzxMoS1S/zC94aWTd+XpcNXPEC2YZt9lNVr7NS3dC260kkMxK/k83AG
ang1HQ3eUc/8xLA4wp93UBsXJasMHsQsIybxtli8WNcA6LNIpKOd1E1y+TLGjOnK
OajRq4tUZ2lx9Q4cruTNf6K38jcViACJB/7TiNSMA7+MruZE1TGIQuLXw2jAhyp6
FZgUihF5LIJhZAVcfXofre4myagLmavINT4ip2EsnI4AsYyFvPF+tbmjQxqSaC6x
RyTBZGhurgu4RNd2H1XNGTfX/qfXWhh1d6AfskrZICi+2Th6FPeVGz3VolOepNeT
t95/x9UHOVHqKJUYXlaJS5ZMw9NCMBbLOznfojfAou+YkSZoYQCgYucMFnQdYtMU
VFy4dLzug7rrfeQ1rY+mjjIc8S1+CK4MMq9WrM04BJPbstpQtS2KUm9uFsZd5R+g
qxBjp1MJQJCk4svTCWnydwoHzHxNyoOcgoeCkhB0xyJfi9x60X6768jCjpzv7SwK
MQvqGQB7eY6jeWAZl9T9z86u1T0EaUjX3N8oM4LrNRQ45kObBfHQvSMJWEeKNHBL
D6YEM+C661iRcabhxdLiRNUhsDSp9o/ue9MpIo8pQGaHTLJ4W/MfQX7mH5rQK9Sl
9ODBER1T7Q97Tex5RG6TsUbmPMQWdMRNvrap4NW2qrQ3kK41zBxZqxO2hsAhpPSg
mWPhiuwJhRcxOnoykT/K0W59RBGS55UfkTJ+loMKUryKU1xAlY5SpBemgMEwgXbV
yXP7Wd5IHB5jzfqT2nRs/9xT8oz4qxi1SodSDBzgNsOxWCIGWrfbaJSftxzzXQv5
5jeanfOpVmhsfybe5Z8iPyIueot77/q2Ji2w9Gwe50P+fQQy4ZZ+xWIZh89DAG2l
hbCAL424mI/t6f0+S393BmbZeLePRoI54PXMGjYk6bo=
`pragma protect end_protected
