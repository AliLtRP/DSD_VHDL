// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:40 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
iZgPUKmocPA3Xp0VqHQ0n7jPC0TrzXI7xPBr/ecQgeluX2IXdYT/Fjo/0Gj3InbE
xtIX7rXzZ22KvyHHDeB+xqj66yfdDhEStoCOqfNn+ghy78FqWSMjQ06uBP9yWwCV
7WOYjsRNmk1oNQOCANFoHM1jWJCEIpWZnZq9SiQYi70=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 8304)
+OJVciUpfbdFKbofZIs1b9TR1nx0DM/zSghabJ54HdTq7H4XjdNGF2gN1kxhx/Dx
7cPVbHIJ7BRn4BLklYr8QPJQGVyVpZcwlGtk7Hb+8pAamS9OJpmHJzb7tlwSUwK+
L7sKbL+Xh3POkhTGGLodeIINyQ+h68BvedgG1DTDrzIppvnh6kz/5+JYIXqhoX3x
B2Up+7kO75IiBmQp5TSXtKE7y0Yk3e+S/TwTAipMZiFq5DszmWwub2V9SpL5v/sI
1uDlkN9uThEERx8T35k+1hStHwa7h1FrZeKCeZ9za79cRdlpI7l7O/slHvoQRD9B
Ld2Ax0oB/qrOBPs6z2jLUZqjAyayAbWBFgIha/5FuD8TO4vz4XFAoRZqr8EZ+JqZ
7Ys8GSiRU5ixEJVbENaYf3OEIfh9k71DelH+Q7Bgma7W8hyHiiBblu3ZHVT35L9q
jNYpXsiNSarZjlnyObVhYPD0Muzk8jJBauVbxBzClkhofDcMHLFZmZHMxNuIQH7b
o3uhSiVq2tCrR5T6u7SDfPUErNmzwGz41hNXjEaBSusmtx1+Du8e2N/wKwjbtMzA
mH9BCtA2zCYUcsUGDQImNIe05+NxqqTz2quKP0gi+jlJHAocPidEOGnQSBYWUubL
bm2/FOR/oH+XMnK2zgCBN2IofdnGDrTrGXlkJFeXccAMvyaelPnsrGHtMyQR7oeG
cr6D2vDK5q8KVM5bUM0pCwQES829H/cy15qIKBpUAQ9gNnLXt9I/LjtRHJRoUQxO
3TZjihfSr2L4y+VVtd57AxC5sd6R73pyFdEnIH2dmIztjCoTA4zeofhejmxVO/Xy
lA2UDzDy5VfzQ4/wVK1K0be+8gojYZ7bGy3sTFQu1nqOI+Dog9AvxR2HI6XerbAJ
b3v3KC1vrwOUOqSznPGWCAC26YTIxwAaCseprSrEj0QHOAOf4ZgDVO0SZid7q4S+
xoUZttydQiboF8mZcUzDPMbl3lJ2PJf2YlZuSA268H7WBGOsFexpiKdzDEESTsvX
7oxNqXu5fjtA0eJ0hqvQdNBtiHvAQoihbpycUHC0wN1CKaEAZrviQZH7TYKwe0h2
CnI7XFs5ZOSqg/o8M9NtlyieCh7WxrYkBYKRqafJF+X9fVGc4UnrQNw6iQdhTR3C
oeLNjT0PKFpuKovgKH3tH6zJcL7Nv9N0/LC1K+gKU9fmd4iVQYaCdrvDwZedTpR0
i001ltNd3FWo6S/rv5M7QhlM4LO35RN2r0LEeWChw2QOOsDB31x3zZKW4auZooCc
lNzDOO0eSd0NW9wGQCMs+4AqG2y9a1uFWWtGYQhcsxIZFsifEmSxqoap6pp0hnBw
HE1ba5FvNsz9UKVCw96mz+ac9qmS9QwGfy6qz45zLBwq87I+Yk44E66YpcAbOo6I
7vOLaTBO8xiNF7iyg2Hpv6D7EUmEHWZzK4Swtwlm1xdNX0e7pH45zO1FaBwiOmT0
PKLwuBmkkNPJHpkYpgs8VEkq0WM1T8bo2FmYTPt/CQzc6cNC4ELr+RUM3FOE33ZT
nqGjHv/QdV14pyRsKWTzPIXjtcpK6KCptOC7YPZMP0RqXDhGTNmCHelBib+n6pS9
iJLm1ixG7pQrs4AyGAS//YZZWltrv5s2hasj4ejlUFWKqb5I6NxlhwxGxSaB1BBg
7EjGntSFZjC1nOaEWc3GFdLAG+YjU7FmEhnzUHg30bWA8Pv70ydekNj1dXpvLQzm
XKO5DSoBbW5KTojxn97rT59v/iZ+3AocUOzT7h3z/CV5BtlDW2tntPLnMpDvaSgC
v8/iQ2aGMOXllWOF/o0gbLRjlmdbpb8uvO70UW1QiOjvqgIk82v9z+YN+TgBSSrV
xi8DMKDfCcShkKoWgrtuXOWbijcQBpCpsiabHu7gAzDTfHA9zYj/bexPukUzl0yD
OiPChAYeXs6c52hTvCNgEgCsxH4z4JBYDOBzVLvrLd9xKdi2BAv74+n+QOGTkZXE
iggGSTaM2xSHgup21XOVjFGsqsOjL0A81QkVI46OHq0McEjzIBo5ByWOcms73qTL
WBjqAAi+6iUNGoAL5BeBqA180u7F0zy6YU9SLhnYIAtPVps6U1UeJjO0wwaUXgtE
Nj0w58x+V/i7AYLiIoR+Vgl9Eq0hqrobOp8RTh1UbdUHtVeQdWRf1xxc4ANK5XcB
1PxbMwImkuKcFof8hisL39XqvWsyPLxThBMe+Xp1xHM0eTwFSFmgChg+OOpAc0ay
QSCF352LzRI0bcRxNs1rzISOnz0G6tFkVYfMs42bZzFAFXq1qv9it17jd+oOx8QZ
6s8K1X4D7jUEKLgliOL73ui3LESL5VAWblGH4YQ3wbe+X+4LYoibgM/BKEZcU88w
mI3zDmpoRRpM8iE6NZj7KKvMHJRZI0unw21dXTILa5a9reIDlLgSQMLC6gNKV8Sh
5bssWOoI2+WheW8YPdhZl4BUEQTR2NYuBPHcGNq3oXOFOBlkOTV0vT9N39xOpGwe
iG4PxzXsxEZTLZeaFeq/IzjRdWBVMRyqR/jYZ7HGJRm8sQMcd9VTFjJw6aDBEhyF
ANgFt+58IrBKxDAXvVXVOSui0lEgH5ORbwPeD0jaPxQX+mT6Msgn3t/8LDCE9qwq
yVw7LQBmyo+GbKrBCfJE4QJE/Y8aHhafxDyMMh104TJPv1YSyiE5ksVWlAHktpZL
HnVCNI5auOdC153x68hhQqBFHd48qHS0RPve8omHqFtUmUey+6VJE+REeDe29lCt
WS9d1Hfr1oez3AdSfHQC0TAAAy1itfTvAIfeFjRtsQt8+zmJQdHhHf4dK8gqnWWg
7Ns4waXhxWGYnpfX40fl2NtR5mpKqKnPIcookFJnNMfwSxVGigytO2crp/LLkVLw
XsWQkq+9fQepzYGorlYk9xzc8oShk8HbLMjgme4zrWw7yKki1DE9M+un/hPHdLST
JZH73AO6GJUNfN5HMwnXPXeqgDn7bbb7dBnbkr8861zPd4TGjAFtrXDnvR+MHVDL
pVxmj1IB03saKIThhRKyiGlY3wyzPGHJLJixAjSY2fppkTeKJCiZZ3JyF88kXop7
J13XzcJXKeoGJ8nggB6fISCl8vw1QxumA7Vbo09UXeQwpyzweDr7+KWQd+mv8xjH
KfaZUY9BeuXt1NUaE6axbMjSR68cS7V0skkh+XHogwByAsQtA7g4VlZWHuW0IoTa
Fjvct80Hfgpz6DprlOjS3aGVEAVDIipe9xSTJOOqpEpQgpsIpQzF4e7ThUxKLfos
aCnCbKeN2olxe2Gd8PWnpPp8pHbbVA6IqrNDcAlaRoHmLl6PO95983AShPpT8mIf
k0AC3VqtSW64OrErPwUsHXuSmCSw/vtwva6SlE59q++hwmc8JxhEeIpZK26XrNke
UmLsUKziSXkG9QuxiHKhxuhUyAT5K1Ng+8iu1RseKxYKs47FYBgjA4X7HwWyTnzI
4fN257WBkZXQwogAU/24hDhQyhp0xzCcqoaiw2VF9Gk3U2CJb2Dsip6ZcJ8ndH+F
cz6+p3d3MDFfgA51oF9ZK4H3nouUEgGv0V0QIXiJnAtHRTzs/RCoFOI9agOuVehq
ji+SamY1a04z8sIjIaGkWzmqQzX1jmCta1uQoGbBaTJHWl68VjOpiYs6IHb/qGtO
6b8Ic0HD5tk5P5ZkKBdRyQCmCN21b7g16Q+QSlZg62xJMFJYgseYyGowX9B7WSZd
nLUFHcy9d37BwtJgv5ONSdYXGeJyf4F1FdL5Ebb/EIJbWS3JZHiUzLkU6ucyCkq+
WKEllomA33Bts79Uep/E6FC4hMI5r61oD0nVhUdzCuyeflOkmR5bmdY34+CMaeBi
st35maU1prr2Vjdn0LJvhcps9ifDC5wgV8DZF6D1lbGgbj/txphdsBitRyf/MfWS
sEFkL8z4z9v2IDISYYmeXkJ35w7Df6SNgoGL9W5jYSyTeC8V+M9QARGWFE5EZ5kp
tTdSUtJEYddlb5d6VxPk5AbV+4JOU9a87UHhSbRFDTCz4rwe3/IA9zTqpCR7gml2
Y0geU8aP+vd7204FWU1VCxot+difRRK1lZS4hXd3Wf+5pj7SGBFmF0CU/1qBBGg+
llcnvf9Y3DwJPTQeQnbFTSLz53kzlfRbNovpzMmYyQO/2IVfG5TRZAdsMhKDWBmx
0+mosrkBloc/x08c/gVQDrluv+bKB4ALHJ4MFxgk+orYmOtut6/WHxrCwupsI1x8
+cxDwALHwtyqssmumwolK1cgye7fOP+DIaZtUvuevJADlfI1Pcy0+znOyZg5FApb
qy6Ak4Seazv/+2aypLrGNhkmj3I4pCw4UYOiPrhptth4e/xqOUWxOYyrKlJyQ4yN
uD2dZqWMm+7CH6j7gL+u40KNLuGrFwrv7iYYTrcwEj9ciAu3+tDw+hKtJwFAZscM
w1quru7VcbBlhxLfSiYsiYgOJEQj8H5TVvb8slbfEd+x09WiawX833kCT7I3m1wj
hcSGEyplAejAYN014vsvGB2HFBBtOB1K1zcF2agk3NovxyqSdQdR33sM7RM9mq/6
TJ45EU3cTB3FeotngKEKWNkJD/Q5Cd9qMuq5VT74UhFWxZdWLD7AqXNCmq8LJKtY
AvDKlygF6CSt7xP4o7UHhTbjXo+PgdCraYCdJlK4fQ7BomRGJUW6n+yso91faPKi
63IApI/ANNonteFiUWtkgPUy+lI3E7XxggwlgdViPa5WPFdcPtbkekJXRqHPoqU7
CDEUhHg0Xo/2huXbDaehVWuf/DcH+lW82oaLqj3WIyspDK/PT6diOy/JZ1QlI9OJ
nWQ1JlQ/erWdHkGWWfcEOeDMuzEnukKEfnY1ntQxbHuq8tx5xFdSXMHqtz0yyN0X
QooGDBVwps8AK/gZ2Aiye5gwLmLFVnwG4WD9P3Lz9uKrtNmun8MjEfPJXG47Z7gd
FTNdZozDlPyRQMmyHKhE08P+mS33YPnF4XUqggpU1foEvypG8OfHdxDZxv7j9jXb
QPTgOgt2TUsj+KElMh0ds2rGF6l+hZ8gjCycUei018w4GhbcZDocfWP2qBCIUKdP
tmUQ7SboAAxWitJDQquHZsks/E0getTe/2vrNnJ8DplGIJlkXO/eLZHPLlJmJ9Zh
ixharN3x/QeCh2o5jVKs5yuW5dhQlo59Cq7D4cfBjAArTSLemJG0tinFf04OHVCF
xJwiurmfWbX0b3HW1L4VQtjOXAsMu584HVE8Px5Gt9eke5cM+eD3XkgDKW9sfKWQ
Ai9XSZ859ED9614QwTxTfDb4UIeK3vdC56Mi5WNR+6myGoy9520c6K7KmmfZr10T
gI4rmmQ1PVA1+jr250PEKOVO/jX2FOMcGX4jhlY+pxBMsy/xyzvik8vAeFKcIuoH
36L2MJyxSV1kStnW/HPSfJhdIogcMCLk91pCeUrWlK3VfQbeUjp677RnjAnS/1AQ
mqj7qW/WCZNnH7abUx1b6mjQ5p246hZIAYUjcZNwGPBfF5SsUFrEeU7TEh5qk1L4
+8/fby89OT1FUTeWmeJImUv6uUjlMEc77QhoT6buuC8bpFHmtrXKJ17AhXw+a2Zq
6IDDdmGdChsw58Wd/8gOl2YvaxttYbm3G01DPZ/GYGBww1UMDnwFuPlW/9CUgCq8
nZtK85Ur1Nt8XgOqfW0DoRZ95thGmYA70Ol9sbNjVkhl2+VSLGD+3R65SGJpV46Q
gq5uREfwWd2Qohj5YFrU3o1+jGLI+BViwAwpoNfUXgKCZHkP+7RJwCHCezPXJNSV
LcAwy2LujUJq4eZn6fPi7knArGM3JoFAHjXv8Hxz5VD6UQspBqsQbycKtxb7g+4W
HIs9b4jzL7LiGQqPzOqYzFz5EuXZkQE1Arq51ZIq0QlnqvbzkpPbh7vvtOUqUai2
5nlQfTQ4jyZE02StvS8qUd1gfFN63ZO1yi+LJgmBlE+I6oSlXyQutBBq5W34FGRF
479XSoiwkVFhELRSV3PrxVnXBn3jgTDwOemQTDq9k5YnLTYbOl/HxE5kBBuc1KaF
heNcyxLYN+U2KhvBw4C6548rvnpGsfV+WEf2rcGCmDxxPM++K38g60nwc5th3rS6
s6Cl7P0ddEcDKFkdTWMa8sAnmiTcLcFat7tVCbfjlOxn14D+i4/lfGxNTE+yrnbU
EdmlbHz+drw6BMncadO7fQhkWIgHs/NQnTGdRqSLP0C7j2T1AUhqeSSHYcG01MjL
MQjbe+YIrCBbKtouFRZBMSfDUzzfNzfINW8fwkKiHXWNFGlcwTx7RdWyorLVrAem
I2fK8LOh9SIHLZm6R/q58GIcKBIjrImjz33jURDil4YENiT/AVMhoGpZZQFdSzIA
XtX3R4HtV58uMLUsWh9KUhYWEisfHPN+zjMmy70VWzPBz44eahjQqFfyywP9X49F
cFR0QCE/LEV70xXTsOn9R5QRQyVndMAXJUaD3Hlu30p4o9rPgC6WBnscSaKNn5kv
6a793OnDlNu1BXIDtQSDErg8qbUpQGglZ8eKDxEpLFnL7pvII2JH2DVEK8lnPTcS
wM3BGbNUUCI6JmXkwlAMA1ma46838La0J6hu0ehPUDiNbW0wb1czrMSif/njWe7x
Bx5YatHm1dzfYlihVTvaKo4FtSdWnSG+kBueNdvrMFXkPUjOiLrviVMO+zuqOKmt
DiqXNDTwhGuDTjIZnkvm7xDHoWT0AEiT765tM5sE4ZEzHAV7f0iEe3NZLXgNXJFv
46D04PsPIziye6LLow8hYGSVsyMEXV4S4xs9GZE32stH46PMZhWgi34HUopCsyo/
G5Ij0DpJaXnWQY3aBXBclMsFE/FhJzxv9nS/fr/manDg03WMiIBqDOdu6tKmzeEM
4Wkk8UL+hhWmkkhANmzQA9J/kniKuQU3vbkyZG4JfVM2Ro2g1NKR8vA8CmbUWbFP
/sdyp7uLj56z+fotQWxHwW9Uk+6pTJmHm1gkINzkHsm3WMer7jLFa1GSpXX9Co9P
an/5MUK+UlYqbiuz1/wSZWcnPAGw+LCG17KzKNgebbwTZJZZTBJd7RNNNsCQgeLg
Lw+ymd4BnzKGkKyb3AFXV+A1rx4WA6PjGTX5lE7fwPSpiCRn3mAzmKVtmgbu0tkg
cvO1Px8GzRA2V9d11GqHWycsc1KnORbW8Q5Rmz2K0JBOzIflZUVoo+y4Oq+Dmi9W
2shmGEWsRC6Ls4ACVcLVNOkARaTIM5fv0CbhEbj6j/OzXrFzxBOAFyOfF4Ztwote
FzFVeYBX2aF6e3Naw4ALTPBbFBZfKaFJARfgjOiGE9tCEuQZ9+xPMSHQeNC5/CaT
n/CyAUJeIMzWo9sd24OJPvuCvW7jNSdg5DJ+TIxepusUs1aZyridX2WqRLvEKuR5
gaVC14nChTcyvB5w1ft4UN/9fdyP50p882H6ZASHwHtAc/SbbYYNVKqjTpv4/0v0
6PMUT5UK/oe4t4pW1Sei+1mfhjzYI8afKDBhKm9DRlXmcIDdqsDlZxg7CoTkBb01
2SajL9p6FCQGNLveM7AY4hNIZekfCFS+I3uLfs1wc+DE7r7ROmYfMKtCf+UviVhn
NBtBrgG80DSiKauVl9toHJvVSvo0BL4qzhDdHhUqw8bMHAZLJVHaB2gmCwaNLhNi
F13V5/GHP0WPWLpc2nV5FbTQTU0BSzhRzhq+9hfIq+0RgmP5BtqDbetA6W9o8q4k
sxlSDoW2yMzSie2nNltbs+PhwhLhOesyCFb3a2ZooWzGXoOjaeD8/rnnDaa3inor
ZaSK4tn5nOXsc5gHzYCQ2gBjG6t9ddQJiFfZ9DeGTcGDEjPTQWqtWvyJoTYPYkOD
xAuMK/je1Ot1MxMgLUozkgkc4yfgogPaUHKjfB20VhTuTbRW+aunKQLvKvzEYAhy
rIZaWeVLyY9XIFz39QCPu2JAscW1axWAOONMZObX94ALsVpQg2Bn23SViaBKqZ9o
2OKMHG14kX28NgKcHIqdrstb3a/XftFeiPj0zGUyrMM6YpmeNHdG/z4fmSaEEJme
nfOQ/oy4QvkrbppI1IDW1PSN2Gb5KnHYnGfUgLFSBV4j79MSV9swA+EVCplBCa/Z
8IbWYuwJyuHU9LpiUG/iPR1+Z4GWIOaTAHJ/eegsoCXXVXeFbMOvWbwpk8pfzYtU
Bga0LQJGWjGm04PCa1w8s1KM4yCZWXGy1EfoW2FrOG4f+SysVK4G/4ouFU08o5aD
tXuy5lFvH1HX4giqAYHvjLKwVVxXhVrcE1WQVI7Llvh6IZy/QVzSZHMF+HF1tH1N
zD5AsGHv4DapeU63xjshGc0p/S1CtC/rluQFKVkoiiNc1Tu2ttxCn8QdDGExMtGn
mxWpx7H2Rr/sddDHngTJjxv73wN++a2L45Qhuy9q6frjjuEgIdPa+x5yfmHHtxWp
5FDDhrgxH6HURbYWGXDitRcO3UqpmDr5u+b7jXkq+2e2jtO58LR40fcSAjnjVFq7
P/EGu5eAi3ka/di+PBmtGKHctGOwkOEoxYxy4WI40QoExComk/adGjA2RQWlqB2W
4s7PEkFqdgK1/bi/HD9lGsCBlvlciwzjStGdBG2pHlNt6XNazwP7NZuyq/T5Gael
ZSCwBnoB93Uri1HpXdDsYXbP25Hg68LDtjUU4SnoPPXQ5+dVE61kAVqTt8tRQR+l
/IlGBJmla2K/XcT6VfUCvGf0Ry4WHXqqdaVo8CrszX59YM1KgWhWH2MfN8k9OGxE
8Pcq2TvAgNQz11enHMluXWqPBfqyKqHIIBvJLQqqoAB8lJlQvg34/ETz3bze8vKz
68alPI1jiY9axJ/Y5YDeCtnFxHNcBXx3K9HkYwYoifQhjlGS3MvneojAhJXxO/Ji
Xt9A4HIP8j/1o75S9ftYxGTYKNm5rm0Trf2dGm2Z8sY7qlVZaQiHJ+gwmpcOkSGJ
WR+01kB/rBElPB7c2PdXOgzKGivhizIcObWvEAcqPrLChq3jAsDQlbtFmOYa6O1n
cmwbcKaHP3mlL6SwsVAIT76rX0BWi1usEEb3UkOgy0DletSDqTmjgfZ9vk6RWKey
W0bcs/fA7OhGZaPn9DfPlMdkL8gCZQlYJmOttxTDMySuEXAGSoNDkWJLr1Dt2gE/
2kbu7E2EHNbeJP3AWdcjcxMNYu8GtVYHB4OASDq/r04aVuflSs+kPIuEf0yyQr0y
kt6HRvL6SC19NAn5dN4nV+grY4K4aXsjkRTIjyItBut6/Xn5d5gOm0pxCYOvJFpP
L+mQa8PQ1ChhodnRRFKNNClrFzAvqOuQeXG3egIWS9+08FoQKDMwK4rRVvaUct+I
bCE8rfxuxv8x/NKSB+BJYA/MJZUOampyF7QbXHVCYYPFrtmWrOoxsSnCypfEVsW1
uNTXIVcGHo+2jb3LgusBbohacxUUfoS30xf0G/+VXe8uXFduDgSLdaOFPzS5P/0b
bNOos8SRIzazeY8CJBYRrwx4Nfw31LiBhGNrl7RddsCMf/+Fh/SKGN78FBwfCdHq
VK3hEm9TqLyQYTyGdXTU2qbhUQFxh6knsvPetEOAPtOONqwr08ZInUGriceVHwmY
pFuAb8X+5gydCTu6zRblrWTQ8DFs7vQf/dq+ZdhbeohdwtzhkwZ9VvSwNjfJepB4
J1gP8nLTRVyGTYz22FgeVFBMPTWOi+OXG40JQ8nb/Gx+NeJpvgpGzHKF4cK3xwhZ
B0op+KBlJSXMLLsWiTz3azeGgFmxeKcUlryK2oYL+bUnEPX8sPVWiJnlUx2z70rJ
rgzshlrgtDpT1MUzVzxyo+enjOXhFIHWtqBbV3Dr9whPOPZ8gpyRgIVwTlVQqmHA
9SYBYVXpZwb4RvgGGxpeXXnGgVTEY4s3xW0jrTRtJdSb+MC10SCu9cOAXV7eEx54
ULVx85yQDgaEwRDW6hPzOoaOj5H5RVl0PGaHZ1JRN6uUZWfcmtI2WoDhAQEEl8LV
CLZjAcqRms6PzlAAhSSHW+1ADXde8+umWNOoUXuEP+VQcweBJBMV/rIOh9z67/U6
3/FJjg46UlEGM7fFZLMdz6eF3qtS0RjYYyo6TnR/G6L0p0RkUcqgmG5YWWof43NV
ZUBYalXA+q7s97dgyYayhp24ffUWcI3ywQNoPVri/QUdnzc5JEX9SnBCdilW5rl4
htieQko0jS27QqFOXf+9K++p9wmgevEkAxa9rjoex6ynYvlto6Z3ahb1fgrhvS+q
4p5q5JRhM424BCkxSeAc2EWlVG4cplNDcugNwvtIrLLDllITZzhlD08qQBRrgBK9
EH5lFSqc7JKqn89brKDMYrLSDc+lMs57N9Rt1W/wngZHkzFKx/7RQbYN8MISkiEj
jkCwNSkB4tXcJGVTpjlxVdbqME+OxWtO52vV5rBkJKRd+drVX0Oi0j3L1r97VHUc
juExoCVSGhsk4Lyp25QJE+NDDA0wvF6AYV/mdSKWjTHLOmICRWViWKKE8jXYDHnd
ktwYAemAH7QYuAaYwJlac89RUvRGUt7OuFGeSfNaN++bde06eL25Y5nIEM9sPoIw
ZGUcSTmWKmR8/sQq+z1dRqJYZDCa0FSrUxB2R8bFCjNcx4t2AAQ0EGFqwGLmeCaB
zDFCRjMwVo5GNs6TXTHvPifhy8vzO5wFhjmqeR7gMCLTMaMxwHIFmVchtcP0SCjH
1K4y2BNPumy/a3c2F0D6tdZ8K1otr6Y4t3cBeL8q2YmSucAmsh8OS0GzymeFqkp9
fh4DlLBIceAcL7ry+SbdqGREWvQME7aBATdh8/7vLa4Vfrwia7XQznTPymqjxwzJ
PFOvncVpECah9c+Km37wZ1/OJ8OuMXWA0Jbv8Rf8wMK82aGGeUQpCD91aIij5j48
pZN9URvEzwQsGLP72rPC2obWefhrXxdkpoPaP80DxHsBPUdC3bXxWE1BqYJ3Mj2K
dOt/k3MyFYA8EQhjMx9h3GQD9Rv8WgBfvhDzpWhaKwZeluXBCfYIapg4CTsXZo3W
auX2rm7wUfLCJ252wNYcif6Gm1LU7j3/gDkuXuNFN+cPtUydvBGEN0R+YnidetY7
ncww5XEpqTA9v+8ZSdfd+f5OkXA4UxEd+t8VyQgJxqkMbAXb0yVKZ9D8Z8X1f03r
`pragma protect end_protected
