// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
CSmod6nHYtImwtIzPgl6BgJAYyFVcNjvSEvIrOjnpEpZ9nmUwPQXSfHbVKz07gIqSIku2EtgzTKp
ZjBETdnS35DIK7766iwPcL2LAU5Z/bvlo7U/wgzXWoE1/dGrwHKOP1cFOM2H563M8p76HYMRVPhu
X8+0Uo6WMPhPGHGipirnN3cVM+Q1Uv+s3PTiufP3gmzmYNpPiPhsyHMuJM3/8pYDpCVd/qmNZauV
XKO9QoG6XnTPqG/rxJYdnwOBB5C/OiYJ7YjfnHhUVGdO1gWCAL15PmqT2mFLEZa1Fa+jzUwuLVNX
6QEFFV7mNBRb5MpmsJqv6zcc+JPP6hRwgTxmGA==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
1c94x/hGzN5ilRH83HxlFt4nrRfV+qvdTSssBkDt9rORT6KC3OQydL409WGG0DCKgp6Xr065/adu
EjKJGR2+Nd1sAbqmavXMfb//i0sqT5U/aBVaG4FmQSFj+W+W5uDzlqC6pClEBC4b+NLzNjpr2D5N
rSTSqBy8elqP2ST9RQh2GdSszgT5CpY99Unq/CgWWRertgai24xOX5sRq4BnmLsVGI+VcbMuarL0
ze4bCNyQhOPgzGQ4rEdnIFV6uoiqxXljcF/E8F5oD9UKPc9nPJDN8vAB8UudFzS7k1CAePSAmy9B
A23ltNQvm7AnlSsN9+OrYXNqjjkEldvfK1s/PPsEkno5XJ9gcy9W+WD5VL38GbJlKlngxrcsr3UT
UmMHTH9jiNr9e3BNmDyUTAIri7+z9dT7bEzq2pNahRiv+jRDewg9LwN0h/FkzYD2rRc26ASd5F8f
taa2Tae+J+MTk4bTldTfcJ4udY5LP9xR4anwc9OOc69B1Na9PXbKAZLSRyKRb8zHzo9ONec+ZeGV
Y1O4o8NCI8l2wOKUDXE8wAaCqvGlATL88TN2vHdTu46pvibJUT1PGU4CoAhkLMvzP8PsDEDw1/Rf
nsQHf+AwePA6FvYCgBs9UFQYVYQk1XXKjMfl6VGiKUFp0+C+QUWymEfePaBf+JFec7h8RontKHMx
7i0CgithrUYMxRWGkeo1uvkGDAlVhqlnI/EIcqV2ILKMkZ4PAKzVz1Eodv1XRG68i4cZjjSLnDoh
Gjm00vlaZN/FU8tmK/3NeAuau1rGD1zZTwjNIk+7AR+S+Vp1oU39cH0k3fwZT7pCgqPeWFnbJabb
ZLyy8nGqEcloGUAcuxlBG3hrsF93yEd4lfqCtRSM1QtMwjQzs0JDiKsThg3EubbND6tSVQsc47t4
obpKQWJUaLM4jjl4Lx9nIGPlfdIEOs1Pyr7MnFpJ1exZJkwzG4+45sI1wCI+1yjoLwlCMfHfnSKw
O2CQ3AQ5jUU/DFfygvZcY68Zt9C5uc/P8hhV9MDsqc9oUV4oKCLSu1MGZGQSi454oTCj2c3nPUcs
0neVHsr7i3joCc2qpB7DXJqNcII/raBmtmiGCCqAsbtcPts0U9OjIcBAWtukVsaZa7uLoz6EfIQq
4HDtF/AlEa7D8I4+6uukDDv4X5O3ZEupgXAcJWD8URzrFyTKXRaZyMZsxc1RtJ3Cj6gbJ/iXOtqH
1c/5AU+e2m/xlBtf59IrKltM6K1KsVlaPT5OyEZrbWFrv+mzfvq7XQc3jgJVqwrjjcf1u8NqIY1O
/yX6D7nXS2Sjz7hFlqmOqLmIb7GghTlv8zR4OYug/3PZ+Qo5JgYAT/Sfd9S3V7k5taWroqyD7gjT
1+vWXB9SI12sxlZxIH1XkFStLD+LAcn3hj/MtmK2rZ78FCGQ2d4NmZBXPbaywwurXOBgMtuu+zvx
3LGVWAN5LsEZ8nkmAtSNadd4eYqZmtpylYVXslmzxmQGXQ663txklhs0rZhPrm5PECLcTId7JxRp
VvoFackBYg+Bpz4g+XQgYj01QB0xamjoWzOI0p1vsaI848s/JHpZYUf3fFCHL5wE7XQDqGxhcd58
NpSEM3Xyeq3E8gl2+u6olWtyWBVOtdws4MB4zZrtu8F0mzzm+Kxdm9JGXqTVLLAdohsPpn2HDWyn
os9D9XqpDboriudXkCHyinwqBITrSlIL1UCNeqefIRhMzJVwQYgfHre2ZEJcKjHEmPAXpSv5v7eg
FWNJFR7zw3lXPXCwnuZ3Gg4uBgBR76cvuI0mg3/eusNx6s1VNj09Wtcq0dvdpcU42UtKWJjVBDJ7
ezTvjE77sOn7OPXd41Id3qw6XVhkeeQqTRNqVsFnpOvU5HLmSqrzCsAykdycuE2rMmesWk7KMAi/
2b0aAgXvHNSiJLoqzesnwQTqSrjIGD4st0Bffx5H533HhcJ1QWyj09XEgmHu5ZAuNxcooNg1ZVm0
Ibd6x94AGDmMTLGOAb+c01BW3BLTAB/0f2Ll64Huy6lCCqNUTk8YBFRyeTZzcWDM0qWkTcrjIbjY
HNiyTI19VB7W+uJHNrMZOs0GM2fzPPCInXSC1IbPrbt3DsYYfR44CmckSepgcUeQI4gEaGqosqaR
2RnrmyeHKaFsWAempRsVKRxYNFPbQsE5Fi4lRgTTGKwch2zmezIMyrDEQU4NKUPTOXr0PF7hFOYN
IFjZCZ/kiEF6OO6CNbq1Q1np91Fz1o0pcn+1+q0jlgw7BRETAlYN7Psn9Txe/ugEv1yAoLcrq930
+FYYBI8acc3NEwKOJuv7TVK0h3oxtxeGLt80Dxea3OxrXIJA8st+6OEsvbnL3oPEsZz4PdQlVGEh
cNrLmCjr3KXR6C79qk1pAw/dqQKpEk4AMBwNv5pAUXFlJdCd7K59vWl93wnZWZ8uqWqFUPP1DmB8
VDibfuxAL5ApItkD1x2HIBt8R4OjWoDlb9Fy8ETMppupyIzVk62Nb1oWys3RzjE7zNbIJIoCC3RL
UOl5x/jm5EsKikuFAJlY+yvPY2H+B4XTS8ySf1UnsXH0wFvB3WHMTYaNm/Pit/C/czg7kQYlGkVO
uG1be2i9KvgNcb5E9UCRVZLz7wwNuyAcsb0+u82Xk73AHVdpMqS9zS/hJBp8jiZguvJi1Om/i/Hm
0lRPCzPYp1ciog499ebdTAYFOpN4gJA0UL4wnaR43OETP1reVbZo4W4RyhHeG5v2jSNi+FfbWdZu
N2Wj5kuxqI7zXwRDeMIfK68W90Ks5VIUI519FFo8LfhBhD7NUOGwE25yHXDl8akMdp3Uk2dpjjpC
FpZLuoVDXDS6LVjOprs0/gfPWdp1cC09m2ud2r0Tc4UeIm0rCAMJ/gndBbBXIhDZB3AWaCbP+2wb
vjt5pu9tV+qpfVeiv4fLAPV9ItgdsYtQPpyos/Z1WihPqxPCksV7s193aOKklaBiFXuq7g9sQpYt
Ttyeo7u0QeSMwyNjU/qhVftIFQVPQlGuSzqpd1agEBkQbu+cxmnKaC2WOi/9k/cyalcTWzaWLLGa
a6Ubzgs+dFWqwe1G0tPdVBXyX401SMNsIIghFDioi/yKqYDG7hgwmLKf2ATE60jcUSIBUoH9f8l/
IwxIiiS0LTWXXaHD3ltFpU0Xv34fId6VVWxewtwULplF06s0+/HCNYTRJsYAtUpVwh0SiNG7z4FO
/rerlrQXMfjRS4oqbAySE/OuIhh+u+2Q1l44qShLQCgbkHRWspacA770uXnoUccB9hzHCGKHCZDS
jxQoQ6N6B7QjiHBmAZdtA/YGT9rAhyHBprQJS+DW7g0AWyGfTJwLFpkkUr2atwDysl1ilqzjPuHF
A7AjQrGPLBu/swiYRwkusqNw4nerBdagmNRFL9EyixeCqj3zMyhZYqhQMVJNzkdniYKOfuz8MmnD
HhRY2gpEgaeoFgAA58Y7Pj9NItkViQKM5mFk9xTjnDRBQczMNLWaMm+LQjDe5YteLIl+Vf6x88kt
J4uIcQ8DUcLLlSqE548bf7Fx76zgMHb4jOvWygQYBwo2yeDLNBzGvs/0OyNEMIFsez8zkMi4x0r1
wvyIS3nrLujF/HfJQWTML7ioMYoVEzrOQZAANvB1mWKtdLC6wcKvhEG2+7rUs+IxhJosmH1zt4bv
RmbLRo6FLqkJuBVh6yyVbXpZ69/CVkD9ZocvSWOiHxrMvkRpn9a54dHj2dHCCM/I+MMfRC8dX0ss
f8gzbxEbmkmCbsFM4owb6OpfKdb/eb6OThqhBPh/tKxp8NlQFUKkGrtUsxzGmyY3Dbq8q0VTfoLQ
74X1EVdvNSZ1oBYGyTErqSKlalzwuTC4bpgkDYAk/APz8khGI2alYhBC/8Y+32AW9n6zGrdz50Ii
mmxA+mtKpNoFsrQXVTBii9jqHw7tt8gP4bqW/iKB0czaZZltIy6uvKjiTo8eMuge11egiGwF9nu7
qp4DDcr/J4n+QGLTe5NysgMI3qBX5OkwFOd/nvgIvIqkSNsvIhLmMnN6Aoo7oNznKudGKxRALwLf
UvbFemRuzO0svJqOFjncE5tyoM5xMUAsax9i9BZZ3+znVSFUd53VIW+PLsx5yx1WmYjiKgl+niMD
3xaAPKgjvqJnv3hc+6aFfU1hDfHxgtBqma68Xc/f+92qd19/jGpZetPdfyjqOVfC5tMrJUaorzCP
ghZ7JpiKvU8X+XXrVVxo6uemt1HiXDmXWuKHacXNljomPLcfgEhSXWGt6MIAuLzirTEeUAFh5d90
rJNxChvB4AfJY8ZJSsSTPy9w+aQfJX19z04Hph1dJHrxOZnET9d1CxpMLogKXWpofLDh9YUaJJMk
RwiouNkZ0qBooEjKsIieSSYudJUwup+iAN3FRM+a8HdZwCyTp3Co0/rkGB1G/EN1nJ/6vEAvsRqK
st8vi6HhIHBgo+mWSz1AABOw9NmBfVs5LgrTUTkrRTz52Ld/7Ls7AqZ04nL/9FKMjWWy8BEjfUJ5
K5m28MhuNoOH3le06Ywcjmlg3J86XQ9diebylSZnzKa0XoiCwtN3HS4itWWWcHQtPkXWeI/iStcg
YexuOoYQEk40xjKmJ2JmQ90wVo2ThnM/981FuioJ9YXJLx5gueIXTdavHLye2BTN8hItTFDkPBDR
ybwTr1uV/30aBCpdAAzlI9XoRjd9Z4V2tth+EZ/U3joZEuGRzOOx7hXoOGhbfGJnzqJIrM9CukGW
b9WrHywUDFIgpdpwjSJeKwc8q9pfMoUozITjiKmPp0GEacYHJBKFISA1U7MzxwaojI9ZfJLHI1pE
q5uyyFz291EtvVEigykr/tRdr4DKzPVbE/GCheWJHew/N6UgUXsfvPM71OhF7uAbzZz5PBMyEfcM
tbfV9a2AI7AzZeGBj9Qur9K+liM534RnBFvL3+5dcjf/aKmTEUw9ujoQP3XXfS4tRGpcLY2Bl54m
Hy/u1v/s7bzG/c7A0lEnQ4RKq1s+NNSsbfGdjmUFS55Frc4diyI10Qs7f+im/rDoj0X1fEy09s8A
tG97WU3QC0XYiEtbwrbgJc/Y9DoMRogXHYpSMdmhOYZr/48efuvYoT8eVlKKcl23I1FdgeQyDaKs
yYvWpD67H/i65rpuEtJaRSAp/p96CejdEPVGRWoHHOASic/CSYw0ONCbWUGs0WDQRaigr0n5Rkgb
U+xYF0wxI5wR4VMLLw9+PsB4igpjY9775oWK0Nke7O+5DHXzUzK45vc1Bx699agKtb41NERw733m
vaXVjI3TZJgambeH6yO1shECQKE0sSwLXm7m0iooibev4UGqzcRGcUco8EIeE1o4GzK1bsXPBLtC
N65lJUs/83QOlEuxcInB4hKGRKKnelBL+RJ+JV1zRfk0I8veTdd4TALQgAaSxf61sbCoidfPrS10
4GAHsb3GS1jBXsVCXM3TZZc0E767RSUMRd0ZidPh5bKYGTHF5d5JtV4RLvsg4G4wAzE933NNA4kN
1xSjCskaUbSi8SlTCoyTTtA6RYmZULCujBpoZXYsYp9JgYlKNsAPiAiSnYfiY/yP9joy20eaIKSG
mM8LBvfunMDYmGsfXyJaE5pnFPNlZSPbLYgBLFgk/J0IElUlTYEV8XwM3+QQ2IpkGtezfe2UPI48
lRnY/kJG9EU/S3iMqMQXyNfq0oVWCWFC/YB+MGZzPBolj8bEkvzMZYYecVDMtdl6SZPW7Yg9XnS4
D2AHWj42ZQbCo5Ogxy1fJUtYWmYESP+fi6zlMRu64b0jj87iXC28MDXUdQvvMfFTsUPpnSnjk+4R
zNIBJdDmdhSS0ZMY9KNnXDb5E3pEqDWc75/RBR2BUGf8YtDApQR5Alha3U6wTdJXbKU/nkBbm0J6
ikBhwm8wS8QP6bM9DjhCmx0MM2hMCHo4+Q2X3R12df07iMc83nF9fotNHsrqmEQ7SjwDRY7xDl/1
JhyJCnfIJmvaSw8rxIVPWfrHIUEqELWpycOAFTV0Drw+nvpDxTw6kf5CrcoA6H5xgitwDmHum+Yb
dq2HdPLw4s0Q/Qmr9+uytM0EcOhGS+sPJo+0RIicL8UVco6Ot7UylDomwaivwmzLozIRgjkBzZ3x
bBTf9mowa4dKZyWXwxONVpK9vH5gD7cLOlSBg3KAJDA/cOraBjiJLstw4sf/U6LflAX8owz/9J0u
kfVm4+xs4ngrYMEwt+MsjPuEIb/wE2seuI3SyUVmLpGHUmVFiUrd8c+P/he4EXqV5UPTbKmk9/ke
Mc4yBOU6R8hOGgMmD/KiK8Wawj6qBN4DCmwKlKsvUIgL1UbMZ3GQ5z0GzLZWi1TPz1BDNgX2aLPE
HoZcF4M47URxRAoMhQZv/7eqLWmCR3bLZngSE8LQ55IttHtq0H9umIQ+Rw2BPb7zYaUBiKD6c+af
P0jwRPq4L8u0bKD32EVJwNkbP4jISKYqHLXO+FNkzBUFOvCwQgFbn4v7fWbudGOLpG0buUE38zdF
ZbCY0MG/VUYQ6IwPNuX/oA6c2PC1sPUevT1ckVxsTUPlvBWMS6rocRHGsXhzJZEOQW+B8Y9E4eu5
tzFA70p2VOTZyGT2pv/1n7+M5RJShAVDcXaRALVtm+dN/3EIn+eSWptBwZmFCq64qyQ6wUnkxODq
bOA8BCRDgGqwnpZ+LhYpmFFCMlDqIn4xu2zE3/lkMuRSW0XTBAvSI5en7VQsHR8pVUyN9CfHivJ6
b+799q/k9/hCzEsurx4gW5sitPCx3/0Whx4yPpX7UojwbnGsrv8pJnJzE9iUYJY7gGrp/WCA/jkC
+xDuJDeYv17ClQ3vHja649dGBJK5eYL1GdXVaYU6BZ3tjYQO77+RbeR5sMjE3HsFkcRnC0aIzH+y
sJxkSnVxwCNWyJvTBDflwpbcnsFklowSvzDDlzExu13hP/3DrLp+K+0hZCpqTh6Ig5SoxKt5MOQA
1EiPGIgP+r4xmIlhAJ996HW2nFiW5FTWarAZZZHY2EcSEN0kG7+VqFFfGe6mAuFVzNSesmwovpPe
DRLOtEBWnc/SzzwsWnErVYz4a4Ery98XObrdtaL1uHSXeBjRumAYLo/7TU04EQwGlCQ3Q7JC1/KB
aqxtQag4IZBEWtRl1Pt4e3kl3Pjcyg9fnNoB+KjAIliFBKKcLRNJM+6Y1NNYSG85F8htqtwsc1MW
fewADdZct9mJK/ec84bOcxTGFReDJpVFMtNvA5EGFHd5nE9UrGtidanb8veiD3qdv/BKBfoQVyug
Hleb12FAdYrllaK3giKdNzfTCT6VUcsZc18c3cVNQVJOtvkl73xRGVc7Za8T3+xC3upM5p9OP8cX
v4csxoh7giHjZiLxJt26fdRLB8W51/K/nuIkF/Gxd64QUBJLoRTxS9XI1jVRhP6alzZ832FpOgrG
YQZByRDfFgMgKaVU55wBUcyO8pxh+CZg9rB+o7PTZ2o874ScxBnsEir8LLme4I47c8LvUZejvqEs
RFaIQgfmL6K+3vCqS6dfKXK9cp1yWXE+jFwyAefEf7ADYPoR+TIr/XoPyLCtyIwAbFOq2h7S1zU0
3Y/xzeivFHedH+/TL34ERmMCWQbbYkBcl7OaaYnTouxFEET4ufQe9I5LspLjiyCEKZTKw4ieW9XA
uWAhIXFDkkRt9BVR+bhN9kuwJg5gOu8M58Z9tijAGLFRlJCiA7DgN7KQHRE389NhNIH60Cl3bag7
b6cvJBqPEjOJyP/JfDdOIY49Lpi5vqBk1rOwz7CxJKiONJM8fEOVDrTAbckq53S9J396jZAWaEOP
HwMBlFDnVbpb2brLQNfPo8Wv3VHO4EoSOAG2/u8bd692KrwoGUYO+0vSx3FGopPDCwfgssl/8G92
3zfJWzAx2V5eO2xRk0PhDNJ+k44lJ72W6YtP2ctax55g9+zhX3rhsruOBNZbRaFIdnK2Fw6C2Qme
pvhWDIRAtSfVElZy0Ekp6OC/HJ10P0qN7nq4+ieoRuDVxxXhRS9yLShtPYjzwfI56+mJ2LJsVt1e
uC8Y1CjWpRD1gcg1rLzsASjtP7hJDfCrR6FFn1R2UeRS/nbDRZUOPo5Hh0w8ynjI8dT1KnG6djf2
eRwj6cAcL1HMZvs6zSorrMdEHNlXQEWvH/hK3qTXmVN+iS5xD+ByqRJjOeLkaAaJfOysFQcPtWSj
ZHXtWAAZ+EmtSeM0V0si8iws63oXAcpg/lMtLDAILwcIpI1tUwAP9vGPvFXqlfG4nHobRi7Bw6Vx
O5lhd11tZAtH1chIzkpITgQOvV4V5xs4kCSOh6YkxcvVYRwJfalo4XxdpkgkT5ZKIm/ur8HceOm4
BVmtjA2+yfK0i8Gy7pWrVzH2y7TSGqMrH5hacRjJX+P3EYsw1lcAd99/o9blwsiOs0oeiLM9RNQk
24zrySt9CHKUTVsIC7wGn14nmZkS0q73pKf7k9tiWE/SO0suaiZYKV4u24romciNQbtmSN4jCcR2
LqZK/PYHDIq9oFl82zWziRzMT8URLJdptYcUNQOca6eIDEcBD6/gEfoFN7HLgJKj+uqi6Jyokr7M
xM/ZlELLG8E5+moE7Je9ZQqa9o74DWFMD5zKpB/dxH/v6MxM8Fff/y7zmzTl98Ixqw2Aew7ioZE0
XUQZzGJN20Zwv3h3SLcTV1NOu7TqYTX2fP2Q0R2dbDqrNiq3pcYEwrW875hYqamIeGhYtglhCAJy
++ky+OcYRu7t5O/3xfk696pq237SnIi/OADEcfEvd05q78EiOXkdxfvQi7WS6uK7BlKY8PSIhBvm
1Zarm27MRNDRguN/7BtsTXbYOjWm1LCvw+0ZqIgoAbtgghliBRd5OT5LAy/GYvwuzyS7eZj/657X
8+2KpgDF/QPBW7e2zjYz9BMrQBXcbgLQohyNmidDXmjsv8oW+WUrwUHq3NyOkqROzwYs2Cxh/cA9
yV1WZXIUGYhGuds85o9wk5ODNPiImduaWIRzCNdTmvI4LtCDAdDH6R3pRMV+f5ZQEfhDpGNG6jfn
nrp2IivJHZ1dw2DX8m9ASHFw/LCZsbE64Wh/t+6AZt9AvwDeiy37ftTrfVrIWPL0OB5QL89+ehlR
CjQ+8g70Jqy2Gzwr4pY08RXbtS4zx1FBzpaT133Nj0z0um6qOZ6gGDus6RBARXoVVmfoBjLdakgz
87axgwftxnXJYboMrMZeuqTHib260ySslc0Ui7bsu/QtHWswysTVoeZjRFtfA6OcICF+Sw+BeO1b
QE16McFrBvQUsDOxUZp45ifYeCheH4xFHj5PmLPP6KtEOKz1s4ViSYEHHudUUFApSuaPGdyCd4Jt
M6i3eMEB2ChSyV4jpIOKCiCI3I/Nr8oobZTc2kjmGaxT4bs3WYdSI88oVRLSMinEq9XL49sqE4+m
eVoFx0RV4EMXAe1dNl81KQZ9pS/NBETC0ZRF7HweEp+Ew8pgTtVzl6+GVWSI3C1YJO9u2kbRxNTN
gsDHsCpM9WuPoET1iR38enMIOpEe/7EB2FPuTjiq3vjYeNlNw/AZjsiAuaVxJIvmeJrIOJDyUw+f
szeWTtyPyVGRGY7EsX747GwpDXhfUEoZJ4nLLX4bEULIW4Eg+XfyQo+3IqRIs2nIxIOkFkq+cuZB
vT7EIhZg55OT2HhNpN/AndZMqoCl0bivXBgDTFVOe/vnGlFH4/IyJKzAYJQPYX74s/QOWRDboSNk
cNpszPGTo2MuZLsEZfguJDWorUyXpmDgeRmEmzo3GrAZQJiUSnupqU0T8CqrnYNb5mXMIZPODleg
9YL6XGoVyT9t4ZwnYhfDSnHvCMgX0CHz73vsSgVDtDfH/AMi4KGDyPpMuMoDLS4XwuKkYOBSQxI+
12p+ndDyaFGDlOzX0MXpc89prNuFoHq0Ul/dGMd0vRYPe8wCWcV6VC5cs4SwI6xvrO+Lve0aExC7
T8w9jnxM82zpVVjfvPfJrivr83ghp5ztlL4DDIlISVM0/NY8QJWssJ9rFYarWKw1MMo4PYiF3Pfy
0PsjLbbC+F9yE2WS9HMYqZrZzsua9xhyHsJJ+LTaW7gholBI8erKVu0ajgZ/81a9OocOtYhpk6lv
RKkmIcKQGSMJswriDxjfnQj+a0X6pnsX2AQyYjID7VhywJ2l1BHMak6+vE6zxahN1c8BrWf24pBA
4CbENHgPOHPOlOTTfNgCyiXA/DrLn0pBbpLI539uZpVHekv6dGgbAz+ArWIP7fd/JS6gTGFPA8bn
GEjRIx3llLJ/N7SxrU3ZTggllgJua/HSay94zjLtNrhD3exNRZ3QFk9XEM79HSRU53n7De6hP21b
FnK6L20gr8VuTabWEFDAOHBBlB7R1KygApD+l9pY5meICRYCUrmwzyvW3H79Kt7zEVD6ohvGZ7qM
4Jj2Koh0+i0g1C693Dd1+Cva/bSFRJ6N1XnQvRlMd1alcXPSxZ6ZdIH0+W3/UO1NloV+iYrBbf9e
grdtNJ/LA67R0iUinvR5+9p8oifPkoLx7TQDrLLrouso/4+zcQz4UnH16+dhuE8PD22IqKSXZ+N0
mVUCQcBpF9NjH+S3ccVBdofbXtg/86/nvVp/OeFtNXOsGX/n6FeEstXf3HraUHgxJqIv1lTVTjkP
/PH/0MaHO7AG4Op46fn+LRib37qvs9zzcnXmOZHZNz/5Zf7KnbohTYbsjQ4giJW/ljbB3jKuHYvb
q8kOWwt30KcfLe5HE7Z912i5xJ141T1sFhtgJwwubcb0Y5PBjTqFajb23DHx0m9j0SpUfRutZtuq
ABDBG4+QCVFe5ZBlRYCoV/eaNZVsj+XWH1n/A7k8pb8Ftn9dcpQD5EImR5V4JVOxsuc5/I74DUA9
t50Sfi2Le3hI4aNeaiuhzX4wBWTdxom8bHpz8JOkDwsLlzLhLgSNAkNshiWdO0EuI5vi6Hzr2BCD
K35Vf1D9HzipWbNEtgDjU+cg+STGXjocTRWinjni/8aVy+ZLut+ZQuGdeGNnZygG7gseQckO5CKE
lpyOnzd5hCNYKyKPPoDPgy+l5OXnbmNVF929W2m7XsWWVI15hBZWEKsvzYBNMiDVwfQPsqA1aZcw
qVyy+qnTLAzn7JmaElh52KtlcPrWo/VSKVDowvQ4kNxXcP6lmLrjyblxNRNBI4gqUeyexngJZbAe
VOtt+/EQDhe/4KjjQzyw7NEQn8EJs8ag6AhZU2+ge79iC5b2Tr9geMnO0cYVnpS77dJiDAtIV62o
kHI049ghe4Z5jUI8PadSgWuzqNOLwAjiATCZtUjgiNAC0IAZVvOGnJKTrDqW+SEgHNGUlvBpSwAr
y6ca7dBXtcjz4QT9I7MoheRku2lWV+/Am+TeKlLyI4M791a0U1r8DoDuwBD4XVRSORj+ijQbenug
djYjOU38NzPT6jl9V+VjH1ubeSPa8jft3AAdpK7UIMmA0e/7k9mgCWURD3t5ds9DukpaBZ4E4Iff
V9eJRt4G6CXuX2Cr47YOTHC2EAwNhFIZ0TUPGar1GrhIQcLsXrZVVoeQqllVAZicv9haplqzo9Ih
nrFt7nfR7HQauT/mUMhVi0XEdS85TupAUrbjOsocCqJH3ZGiDgXxCFsfdZ5McyyTZERplLXZI4TB
vca/HGJn4TvLodJZccqPBKqiKOUPIXKyvCafyXU9Bd3beKbcVezOzc7x9yuieSLuTo3+kcnvuBj4
2Mvo9G1ftcGtjeORcyuPAOpQ/eeIELlCebla4qy+LvNbl9Vg9kj3yd3ML9tMxkX2qDm0+/aHkM4z
JiPMYdXomIAXbjUw7iBAztKoM0zRhlfQopjF5Mkj3AurS0zT86/+vRQXyGl4sVNZgIVlFYZRQXqk
DdLvq9+x41sWU+Ato411W8b+aRJNzvXSBoGYVzEgBC2vCnncbxMzrqXPUXqyV1nSXaFf6PbgBgl2
uklIbu35otNMxcwSGlUEZiuWL85qSm5/A96zGyVwRfd4HdSn39cDkxJIlucg7u5ly97RJjQ2IK4h
BEVZ4Dwzfb6pTltfvddv9GlNhQczSzzOU0lKO8nXdD+LdHcUnuJouMVv+rHMrikE1VTD4TXHpbWt
eCqnh3OzQwTUUK/KsFWBrLF+ykpZ1yFEdC0hxUdGT/PhCTUnQhyuLZMS+SezLF77CLHa3w30Nz3g
slEiN0jpJvcyzmlV9eCwlegnXCiiul4qKXFXs/2kqbwZkp1GkUPyRTNd58krI6HQPtRl1I4C3EiT
4+vfTlWYQeQNH/R0e25y5j/GIi1WPiTz9QgBnYGksocHQ36DxkKzB/gMgi4K+RqQD9c32G+utchj
aMLMVsCzlyBvtZ1Y3cJAT0SvpvYb4/JJhBTUFfiJYHv68pZ8no12GVXR3tv+uuvYDdAoANcxb4rh
igzwLdJ1Up4d+74EpP4ddSyxlF0UqRoxrkIVS+JQzyZOx7HsS8zpwXDK1yXn00B7s9wIfKIdxwsa
RKQekKPlo3PT5AdKvtDWDZkfORnSl/3Y1wV6BmZVkh/yAd/3SUrrzUzOtadvZZ7M/HXauueC6Qi1
0ec/nJ9ssIE2sBfSyLcBg11lQDL08ROQD1qeROFiiNMsNhRVqTrYT3XzFc4K5vHmhRmTFAz36c1o
Wf7SfGsb9EZhRgifE1z5w6+rdqZW32ZIQJEwGLFfBKf9X7XvHlrWty//C+aMs3PpYwmZnQFQqpm8
0oz3klRoCkpsTT6iJZ+0bdVxhvoFY1UiZbFCTijL9W7S8iY39ASEAMcL/8FI/GoneZjOMubjVZRQ
ByI5XCewF+yUL3vCEw6IMA6y6zuNevfTndg2koTP4P+90F6suNjet6HXmVigLaofMJtIltbRECZk
dE39bAdRDgM+2FmzvZ6IzILLnesmgzdGW2i/C6ki5ri25NbttXrg4KPQv5BYsnednZSn8m/vnPAh
+StqKswduqY2iYgWHHZ7bx06oohhfbuIVwEa6cipA78MIPAHomsTAA3IDOw+yFNo3S4GxVRv1Cy+
vxEZ1sx4BTVPec/yoKtXWjZxd7swCpe9MXmWXfzhOlSJ7//whgLAQ3EQXwBUJWThXACsW2HH4afE
8S0vVg/bo1xktGhxfUe2e009wBCexdbo/2AhTKGk8R5rhAMRH7rtL+WFSrN/jccq2aGxqwQkoS1G
4Di8J5mRhrtiYSLGZ0mFoE2enplU0yC6oDnNGFv3WNnd1o2u5M2qJa2+NwHQ8Msu4mnsEDwRMwtK
kGpg3Bd8C4wpmsEiQ5/WhqY71+5Fbo3Z0ZTJuZSHtTNV/y5Z710yK1/1ZqkNSwpViMRisV0kixHN
jpB7Y75DDaeo9cBGhHpE2QHKPCA+Y00dge73cOVhFtFDpwkL+oTUWXr3MZHoiOV8jWjfmrMhdHpn
TyHi2ZjJca3s77bM/l8/4hosRI/9w9bcbwyv2tKcD6GkttRir/QuLUnDQYMXdgveEaH376CUeqOI
i0R6uDdGUDjTkjvc+0Y6Asi+2y6sROhPCvAWHugWExzwNl3of+lbV8f7+72Rl4aFpSaqvjEnanAO
sYCsvLrXOpOmG/pTvvxefLoO/pEacc73FRaRA4S7W0mh4rpfNsZfZ4AlKonc6g/Xlu8AY/HrYQeA
m7zsM/YUZIbvmTJeMgDt73TSMKBcf3NK3rpsAZ0hplktoUwKoLoRWABmNYq+fcvs1IF9VzIpNwPy
23KBN3Yzl/I/p0qIeVBhj9GVrYs6pLVwa7cEYwEwduSfCHxadmVfDinnsjzkLDRv5+9qEikTo/EJ
7ANqUPElkmgZgy/AJOQeKtxotO0Gh9M7W8hNxrHio1MEp/H1yQMNFaWF7/8a1LNqOGwkBxtA+LB0
Q78evKmprowlw4nuYvu+htG3sEszzgGAvoUar5aCLIYGNmCza+OuxTP6Suvqg1DSxkl2ZRO/iwyZ
3e8ItGT7ae27eWwZ6kT9v7EFFZr+5qrQhrFIduwXEcc6YWVe2jkw3MBuAVesBaXkwk4XthiSoWhU
rnIko7ihKop2+aFnHtqRAmQq3FVUMjr/w6cIbay6tyr7t/UC+VnWEOC+CmcFe2eU2uMMBk5H/gr/
bKrVymUhBKLWKknmCSRc1xoVhuRziPTcEbiW9Sk801VKo53Hp2bJIl7aTxvYl/cODW5kxcMDuLf1
lnOIems2++ueL7PCBvmHCNfAtBY+f2QAn2qPKrBc8Eg3JsqCEmpUBJVSStZOFauc9m8opi4DBRc3
G7UUygHB6DvuJrVOZrIa00hKCKU7V4yWQz2d7mbgshfHLcA91m+WsoLrDh0tRbNT9Vq90LbomvMy
K+qS5EeDh6Ydbfkv1z1Rjtsxxai9vpDHkOde+qt1xzgVDPuduD6UQ1sm+eUEQmv0Rl91Y0Qs4T4v
j6CIVh29vJ3w/7czBLhAMHgwVhJUngsQ6YAZ3mZ8K//Yv8NyU9+c0CwBYrsESeR6j3lfnPzrADHU
Jtz5SCNjOpVntt4FbIOMC2yDFLZY3o7Lz7Lu2BIjgc7qNnU6InD2p+RIWoGqd3W8F0ydgBj8Ps95
jahgAc7DGk5g7axrVLiY1r0gH8qNy7gtJeeAzPNAepRl6xohK1o4eTbVw3caO2COft8ldXl/6ZI8
7U2exZizJk1IGqyC5djAty8y4jJNtXJ14yxnx4C8litGa4WVQRPRBpBpnBYFHKbwLeNgbt5Hus8b
2Wv7uw0xosIyFBJ656/8RJFHqX8HvdMwlrcOBZndwmvq2ksKB0QoZ+5lpZ3IX1xJpG8AEz1xDRVx
GPyHe2PLWnNug8/GyFm+sdxeZAE/l0j+HNbMEGm/qwX7FoJ/c8M2J+UtO5IEDnmaZPdErRYpImZ1
w7MMcCmwTq+F0aH42VcFyz8vNUS1O+ZW7CwhSivQ2dJ65idW0v5jPhCFmw2PeI9wzUw6i7MDjbp6
cnPfdrekQkwcFPiWQoTEhvmsw8m3Rw0j+mNKsfU7DYOXryso1dApOTq1z5jHz3wiCeEFB2FFvYcg
Bpphm3FYXgJkKA8NfbdZ+U1VE+G0kWvP1GXe9OKdigvPP9kiYNys4nH8K/2kECCN8mr4RDJaEbIl
3jxsA6ExbA8AKSzUWKf8m6rRl0ZfJyGUaBe9aPcqgYBiW6dURLUT17DWdqeWMBnvsFIw4f2vMMFK
Upm6HPbV61npKWgquRU8sAunOspdYaa1YkLvdouknQxmg0WNHPL9c5LiBVTDNLm18RTLalFPmzk2
e0NXwmQwrRs+ztPdieHc9zh+ZG4cm5uvgyjLLCflWNETpR/AWcijUMhBozIM2CS8aQ+yVukhHwIg
GVGM+yLfIXFjf0RKbmXNihZqDjX1Wdk48wPtyH+jhCzyNW3dRvkgJRzLqP/dEI56SS3x+l3aialU
O7pZA4ZRxVwnAZImFGHoatV0lp72YPHs+t5oN5VfG4Mjc891RNYKpBCYCxaqyObnfN8zahVfUSzv
ajxZo0NT9C0QVubeTekHM838Mw+7UWNCDWo/Df9CuHdtEX3BbnF8+Kv6uAPR4joRQWHEqcnNIExU
gyTegdX1flKTedKjXf6X0D6k66RUDuLehH68fMPff3CXsQQgEQfpy4cu0p60pCOvELhWzu3BJZIT
5u1elUK90mLvBvU+2odSmnJ8LqAVAzGMR6Zwpo4Bu9UG79qReQ+7lwn1QLN1UqiqFfC2VfMzUU2k
ExJsVyqV/emrR74cbO0Xz7EwKiaNZt32OSll+mp/tJ+4wc0lpYm7L+oNGN68cOtQ7HaKi6aSN54V
eBohfG7joinSupxQKG9kNBFp5iGGl/akSRs3QoD3JjuHimNej4FbpuJpN4iMapScGGKF4OMlv8vn
u+hTXgY+lOdA91Z+1EUAsAVCPOKVCfnzz6LgheBSHulUcOKQoeJHq0RQcmLAk9OOxAS/WlZCbh1M
hYvwGHDQBE1QJpbCWy+p0Xdwab2h9ikyLGHzWNXN1SMnJUS0Tsk0IumBcJ8VGTDbo8hAEZckxb4s
oZxgZCkSmmAJ7EM7BkYLc7ofIXDwwZBZfFSMR1zqwtHt42l+80o+0TtPGD7ZOjKdqmEDiRp0o3r0
xLGQ+CuqShlzyfTFHjR5S2It8bFKf6wSp9iYbpxlqD5bEXEoqhpDaTWuzj5BXQw99Ud7DQ6D/0DN
ar9oHpKxQHVB6i7h38T4VUBzVnnPzGspMRlrOZN+eUe2eqhkFcKeZA/KNfkBT6Tco2lqlvcaWQXl
WobUbN7fR57TEsmR+tqAkG6HKf6WLOuxw7iGmr8tF7e5UuMeMcaDc3ia0eJxBFORGt1TA8up1bwG
st8zPTa8TQng3m/xMV1XTy9YPx/FS1REV5cuLaSVnO6WxKz80WlIm8LE8vZl52TXu4Q1HPwPjpu7
0VIVX8d2vO8fi/oCC7/7nlOg00sA5NP8Ve9WpgclI9mq4EeylttJaP1QEpB6cKQT8KfP+QtQ9P9E
d8llCNQjwAsGjhIQTiQfjzhiyzCJMb/BQ11f9gT/b079dl9Vnsxp5RZKDq5Phlu7/F3c2sTP90yh
d1MA1YTphETH2WYpKqDXTlQBbIifygur49fo0W0Wexnu36B1V6jkwW5skihCD8W7bBmXzZpzZOZe
YXWi83N+fD/ixjxd5UkYGQwd1PJTjN2QKkOb7RZ6KVrRJ5vzosRNVNMOf5K5PyOEHF/f/VIfv6Sq
MvvYgFGIeRNDILTPvLbhHX5NE0uAwZycH1oQLPdNqSpwuI7Ii5e2dSTkR73bdMDMFnU6VztpzPld
ghZ2/teFu4Vt9ct/prUJ0p1LsMucqloeaSYEhMO8R4GLCrho48Z9PSUnXIeIo/eJYLanjoBTCm0l
D0OTe2KFlkum2Toy/1du+cmaRVfVfi9nnjmmvZfR9Gd6/cDqF3jw6AWE5vNbg/BRxljXAN/2UrCT
wb6A49W72ogfiUl7yPDxtFLzG5042HE8YSHdEKdGmgmp9z5E1ycg6+yPskE48bZF1FXtfcC54BaK
rwwsOPtEQ4qTdPeZPLNwB6PQ6+0LBOzXRGXZtZyU8XW7gIOWojgBG42m+yzLNi9LbIbaJLEiMP97
hzTdf+4Sz0nL+9RsUlMPlECu1fRkTUMdOq2tzbl8nnzS+KoSrI4Z55dktdbQknsrei0EEoO0o1KH
JMRChK635+MR+dBwntDVK/c0eYACr9wy8oKRS6OAxrDgiH0SFsv9iJeSVD+L3iPJA27LjyRs/flZ
Kxh0KoeKienYJJ2TJ9dvYdnqp9SzdaJRUQm+xry3e3EYvaty/+iOXkcD/pBVY3mn0g78/IBLhBUi
kO1WUs1RmorghyMwlV7qEu1OR6EsTrefijMK35Wf9Y7TQpFLnzzhJ7iaTe1HFq9nxCriKtp1ZODg
kMb0hV1EloakZaWRqPrDP1OI2z+80xZQnamyynmrSRLo1WCqXSB9iX2dME5gCuZsKQMzYz4SjCGE
EtUlsY2NoZNP+9IDVFxsO8usAAnx0Uv5veDdMA3SSXuCQVNGQqdHnFGBERVU1YiU9XGgYglXsnEY
L0NlQmYHwbqblpcbjAkzWjSmfvNWD0oYMw9O28LkTo3dRTu9WB1JJPm2Qmr8WCn/dH1yHV686eXa
dhfUlJl1p1xlYCN9tMGKLRtA1qxlvhMLrQOEU5P7m0j5J/zI8XEk6aCp5h45x8pvCCmc30nbjCKV
dHhOSw/WX+coZavl1JXaMhEwyHrQ4T/rcjU62u5Z7QbIkrvtX8EIzpCw1ih77bfIPWdDcsWe/cJR
7jYOcv2ZwEnH8XImPwuSLWxC/BkEBf9390q9mQxpWHmdIX0nwQfPPrBXCgN7v1dGTGI3exy5QlUa
MNbpUpphnprGt3N1UTX+R7qCi5zWHS/EO6RY9jcuVRLvV4Z5XVrzYNyOEa67w1DaE3iIHFsgNB+I
sPKJjpk4LDmYtG+KzC9JSNs2MA0EgNS64C1LrnoNok/18RfLFV0dNWU+rnuawc8v7foIEr8srGkJ
LoumkT1PMFfLwP+YZKpZHPPbdgsdGJg5Oh9uvuW7wOBMp5ltUOGfUW++KU/lVQpmWGXXcJCAdKa4
t8pymVytZlsg159xvTj0yL/tpaQhGrgUlEEwWrGzgqWdTyuDqdCH10GzkYut/krMhtjDrBb3BkGA
cGRHnDXz1+ZZPVKvT3Nu7ZFfqxrZFg4/rBy7ArxxTt11KFKgb3tfpqtZqs+7WHxx3ryNUmqthcgx
NKBvh6g8lJFCE81x8QQqXTS2FrmGSxgX2V6JNBz4lpAo6848VWu9UDMfiNNDmK6Ffzaixl8NR6od
Y3Tb0sc5AEgObJYT7ImGCtB0EEw9QNSS6V6z1LT3Z+xwxb5uT6cH8DMM2K6TJjf/Ag5CE9Bvzbpm
UqSzaO834Tu93JV647ZCEUcTzIAnQxv1npuadEe98jDoBPl9YcmNGm7r1OaUi17H8ktgC4y12M8l
1grP5dl9tn9E4n54T9q3QppMP/3exqSerqnFQdaWxw5nQh0B59pjonFaAjrMGfOAkm/BNkRdLlco
SddQJ0QV7ettoFtFoHw9vb0bG4+/0CvCTnQngF5NejndyVbvUCURY/1vC+ZecWB5p3qbY3l+2dUa
tLxO+Kzn0zlrwuJ90B2IlI5Z1HNv9XkvFi1iO2eQ1SxPu9H2E+Vfl/0QUtArudNe0ON0RfcRy62K
FMFmwno91sau9D5iaeMqBciVPhex5GllYq1jPvuM+VWgV0etqw6Cc2vcOiczI5xP3eIdXOzPryZO
wV+zWkJKY61QsyYKe/Wv1haD5iETH0ZmyQFwNExpN1axvM1/eSEbwEnGc4nER9pWhfLuixjZpsHg
82zwHkFOLxh34Q/BZY59Iw6XsroFowNK+HY/4gcWhMOU3CEphee3DcfhieL6w0lo8tsO97IwJMoZ
5EY7O9fOcWQ0HPGCfDw3i67LogitB1S4cy+vNSfu7/g2gqDu++aTti1ORXt10j+696KXNehr+cDo
AaHB5+e6vptFLtni5dLYC+TmY4atQ1svfoGdPXtkAJ451CXSQihX/oqzOh6ZEJTHB7vB0Z1qeuvU
Ui9VJg0y2ELW9SdsGU7U2I0qiJd69bW+4JNMezFEQZJ5sXLBcbAS67mzWMOimbgBIMyXyz4fs7JE
DWvqQ51TvDzaygcobKIil8sJBisIjCcxysavXbavdTw2wGHXoIwmla757JqX6mwtkyET4auTywuy
LWaH7XQLeEx7EQH8IXVq5CYvBmaOizjk/ZsEJveR09Z16BUfjEEznP7+Y/GzNYwI/ocDAXFz+hVk
epfekfwqEFnSjFXuxQ1lzxkkN+QoQ5KGBzagCZqnztjzR4RiT20G1GMnf6R8yuBh5Gce9QViYBEM
7NCs0pyvdkmyOed9SaOOr9klDEUInFJ0AkqHRrCTm+v+HU2SdFg5bYWBAyM+KjgaNNpF7sR1IItP
SYQvCn547PpWrBAcjP+7geqZ39WL1voSyX3+bQhvVmHQ2tVgl9/xUBmkM0fyXHeOpOXB9+VN1ais
usJFaP4d3+oXsAtlPa/0Rs8fTuRQkhRucZdvDQwm+yFnpwD8fXU3iCt3PNOEhBk/8+v7gG2dJOp0
azhlONj8lHQr0uj/idkIAbd+NxMQzVyBCqecePzOhfwCtwFYRuAwVGmFm04dM4hsy/CjVp+HXf3F
8SoT0P9PBSLTKHrwiOKb+P9JSnCnajCc2qxxgsnyNrMWHXeI3bM+7ODKgMW4fjlkMFhZ7EpIyT3D
Rk34tfyld1Z5AlyKOyM/OvFoYJhri0e/43wsX04Vt599AlWZBZ7Uu2gIzUBe4bxk405qo7V6kV8J
fjgZPevYNh9P0GsGyhm7B1Zqj3wVGwZ9nU8VD04EoUt4+YteMzMwdr8ReS1oKYrpY+nmb0Qj3Zth
9YZ+H5V3/6JW2gbwizb/H7TKqmU8mb36zwkZHZmkK8lfN2c7Af2sgFC51wxPwhsckhxUemSt0ZPt
QAhw1Dt/PfaUAajdGaIbXpvD7wlTBbQ062Xw4X5Zk5s+x2LPAFrB87SkMiIJGY5DN9V76knGTK9O
G9WjdznzdHtZ3dKEBhWtZWPavft0MoR/IRS2FyE6BLwG5VPyOuXxQbPK9juosf9TyA8/kgZuwHRa
pTHgT59KNNVvDlCvjyGJwRY14MC4gkp84A1EfGJoZjq3GzK1eDt4KKJxgFyyQ+4t+uwNrNML1Jqt
PtDejE1U/LktUMuod+BqTxouZ5AtMkC/xJAJ4CUDuKaywn9YkQRuEsGW/Gl9t4sbQGs6P2cecmJc
EzJD0MA7wfQCmZNNuWrrBn9puERPc8cm6+N1xE0tayMkziIHV3JBQAqV2jf9fZXekLTBGhXzhXaA
/Rf6A7RPB/OzKtNME7mQ6eFEQKiNfe8O5g5KjhpDNrIi6mo1QXn1wWXq6wQIBpDkDCo392KU6mNA
HiHJaiLFtXm8DDoo6YqdI54V0pyxL3e4garBkAyc7WHMycpKSXTjYFoyUWmMoW7zSSY4JZ6i7EUK
OvfG4uj+kA6Vkl+B5HvFHcKrcfeSBqJEoqkAs5g3NTOwO0f7e1qIelMHhJanXOwHzTIazm4fmiM6
ztEIrIInKiktbwdvXvbNvYncA79qBfUTAAlBkpnJjDc56JsQZ4Tt8PxDl7f8v5F1D6t6jfJlkrUL
AO7D5BzqwcUNLJkqU/L4xlDU89YOYiihHwQUQISjA5PXE0AWY8mOqk/LEU8gWymvABLt0ZYKT5vY
u8XzoyOHuEUhO8cXvLUwg/aFUL75bdBM1018dCot475pAaorOfD56inh1wThwtQ80kaCV/OT44i0
WswxIGoczRPZZhrkrftFVfCrAxXjV9HMeSgxkuv6N3d9LzfrlWGXfI29i4FfWBlBNa3IH4daIxwk
uZ64E3tI2m9rumnHmfpeYiMVrcxhznmqh2I7e0DmS/Pd8RNo1UQTuOK+kBDlP7W2RJ8IFdbgAehf
ZywKxx7c1c3cjNmH+eqQ6EGaxAp341IK4oWVkR5G/LHGWp+s1k1Fmv0d5w4N+KcwbfzVkLuGomSH
LAlsxKrFpYG7mvLzWID4m5PV1QrO2jeUsIGeOYEZKv3IUoZJkJDxizez78VjrQ87J75lld7KrizW
htJO5Xt1BYnoxJO0N3MuDXrdM1mspLVzM1DanBZRzZhiA/JdD2c/C6dd//NkLGEiUBh1ZzgBI+sv
hEYUAe6n45eBC6bBh8lwgwUxG4SRnlgRSrmQDC/A2GG2ZAnh0kpsq6dvLMotUyYcNHRMFR+ufldl
1C5W8ttx4bZpzTAJS5ouFUobF+pmsGSeZpRa7xmyizDkAhpTI4IjFG807HaUpiyInhzYwuh7MT3f
ulAfy/2SRZbiDJXxCeOQxYtSVbPZf3DkB3/7UF3YAEeQlFT3we/KMkNk0eVJNxgEbuCZhuzqWsan
dHKqE2gbm+cRg8b4lnnlPxV5LhxnXdKiqPapz9h0PEzuFDNQ7xYiWa06ZmOXFzPWXqQoBlXrM21m
SF1jFfkUQ9Lv8E4OgrO8vGWSaLqg7ThpeGilVGxrmXIKbo6Okt1NjkuLWxlERkXZZ8hfN+RfmTg2
Ewrq10GNUpZ8rqHHRQTj6FPxg+yK+nT016QDcTZmzGoG6I1VQRkpQFcz9eDFRon7l6ehhn4FKDu0
oY+7isTZ8+WWfPYveQczb+EgRMjbCYNLkPzZQVQ+ctj8ZYdsn3k3hvaoL91NSU3cYCXE4yOWtW/w
LqhUBbxw0rPdu1SHkkFM8bNeY6Msy/LGKXLGLsqygI7EdBIDzwa5t1XEgtaE8TVYy2MCGAQx8T88
DFRBLb6nVUrPALNIizi/tNKefbEGWHYnjWN80GRg56vXfDyO1ZcBWlfGQlO6xaqeOGc5nJ9lL3DZ
XTC0/s57g5hPkw/dQHIM1sRAMqb7U2cQhZS6KVQXTyzLQk+Zj20saF2hlCHsT4QaqQT1D6HIpvTA
6+IM+5w0LkElVbT0bUA4gq6uGrtZGWyAykij7cFrCjufLZmu8c7haDmSOzbkLg0sbWHAB5D+kHM8
LSKoxfEYj5hieuSs+8fIaSowbFnnYJXd1lqWtEGcVVyl7DjCV+3510lD9+N2FkdzctPOkcQMWR1A
2WeD3F+lsONzlrm2O/uP6ekU2OtpB4DklBkii6rjsi41417E8ewhz8bqjQezHomt8rSn2mj0bEXz
C65+zE2aYFAHf4/tMSPGI4fzpgMkLVTBiz7HzN80sfjHbqNleLIcoaDMATVgY9v2lmx0Z4kmWVxX
1jp//TqDNTgMyNtFkKDxEJ+oBRk0ZstGVWnRuEQRSpoPoAnlQYdFuKnK/kxDt6+4uJA8b5usJRwP
xZZn2vNCeNl31ejHFrvSyF1CIaj1iicsjedPWuTEp204NPWiuhcESW26sl2rIN4NLmtO4xrK9TVv
UBoTEm20CR+OD42WsXRw185ZWTukw515ZDWoFk12VmM3nEX3VaVCXF3mPaIDmghglkKGqtOVrJ6Y
Pa9XIkMV2JIbzyErv1h1ye/iDomEkUtx81g0TLQwCCaHYDoJzFlB6PNMOwzCEeKoJwMsZmZX3RDI
CFnLCPtE2hDqOWS3eq6cxEjtbqxAFd4tlguprG12HHsGgaUh416XvHAocko+wrUVePSVMmNAVrkT
jy469RPsruqFhDCqeU1rBsTHxdOI31SPw1+THL97MGrvwz9se7UdwI4wEnz5LlTz6uBcWXWqzHdu
H4DQXKEh4mTfr4mMMQHaOtNCcWAgWzXYflJB39JxUOHZY+Qoiy/RBlXh8gHl18sSlbdWjKPqioz7
p+7D7eDzCNITaVfI2s+1bXpnvBCqIbtrzpVbRUDOZnTiAHcJJ8SuYeo687yissG78bUr5gHTkKlz
WERAaJKQw+EEy6AEJ87eH5bQXanN+q51MdJqylW+jvA+ULA9rBJL9EGv0OW8JEXYOddeHwM5EZz3
Ju+93S84zPyF4qh6VXgRS4spbk8ehP411LPPYZXDBdPZG0GniZH+iingNgGKtxu9IhZx43YUDvDp
zHsCtszYwEPbdCrytOYSLssTgEWdjryz7JZigzYYNlynw3Niqk9PUxtlC1fjn2VNxo8wIIIZHIxX
CLQiGFOFki6M5gajAXhTv4Fyw7Mz1hkJzCXkVOqTADLExR9NuwaMEyM+GRmt4MGgdPxU2JXy2I0g
fobHdqvFK80xn8y37yAI2N1szy9AoNE7YjVsvg0Eprj4a4IJ7lzoNC4el0DhG5B6Yrj2o4c2WKWN
elFp12C3Y8ZyQwpt7/2l3/b66mIMppAEiDXCqW2DD7G6eQtF+19/0MtGWxCODIgkz48HlHINKhgI
wzzUEPMiett+PbQQDrnrnG46IRxAUepTvkP1QnB9zmVM7BnOTZGtxkZBFB0bnEjK9IRf0DrcGHZZ
X2tH9szqkHmWFuatv7mM8UMn0VySDnwAziyxKswhs5xEUanQfx1PMwllmfPXEcyRSMMhUpkjJIrF
MeQAzgQVHWqj2DXbGmAMD0lDo3RGMGDJIFrOQF5OzqaPCzwgNulNY0lEVHwon1COzKqOl8IORp7F
qSLJjC8S51nEZfKt7yYzmznJZ+XHAHVlOlVjL3Aa4NSvNNO4Nw6JmSn2Q8x7xjlj1tzMu9otSf6F
hJtY3Anr8NRURZNa8KFSw7Q8airkBnqjZTpWdFJ3PPoCjECs3ogyLa4C3aq7GOsXWClu7OXYrANH
AECKg4jL4D333ImbsKOgrLoo2cjwBS2CEF7N0Y8z2Q2+VJ1D/O4FNjV45EeNiBXPic7RVJEUobFf
nkpggV3hbyGM7Bu9iPaQqzlNOwkK+jpPBWzaFAbVFei5uQb5Zc8UV8DjbtEslm+mKitef8Ylw7m8
wbNYw6fp9c3oQggi43e9OHZMwAB8pEy+Fnyg1Su4Wn9yWjDYo2jQFVAQDJO6swxRd8/KYsxTqjeA
yfTvOEh1UvvbLmhktwG2QERpXqBevgZe6mWdYWBAWvjtT6u7BEJORGbJC5AeUlD6jGyoL2k8JCUY
hDqo5LFCqSgIilDve/WjdB80UZp1GJAI0uO0QPIk7a0OfGDZToHu/1Jnivg52GnIO4lfmgjyacR3
EjAA+AUl7U+GwnKQdcd/WxzPu6n5BwVJfxImmYQzZN9yb0tuE3jv2GiQYxzxhm23px/NMXen6Qsa
zMZgUoR+qzCitLk5iTcxHocSltWv4cyRTqExoI7tCy6aI1NBtH0dHamCsqL6yvEDJh+KTBXw1cbj
SQJ76NzOZgaKR4DGjsCdQV7sUKjmRZTpFkGhWI/f5My+s8rbKLN+yfbQoJc75D9gWSFhRWupKRqu
JqL/Jgshmx2x3GVmPiTqeCYUXP6iG+qinWUK39d4Wb/KK2zBREqicfRc6dhfMd29DTot0rkQ9PPr
OPcQtPXAD6MqMIMGPE5xRE2Ep/jXit7F7AkZuOeu7lA3QzG5XOFqdOtDgMZKVD3iwjCTMo+F0U0Q
2a9dYt2hO7BbYXpdNT9hYKrzoXT6kThXWWa0zDECrOPyA1gzKpbJKyTjfyO7S/GUcuFkdNhm953o
3hokm7oIBOL31jl2KrdLw8knOEUaUFxZcw97HdHO6P3Io1id2xcEms6RthiWQgu2L/H3VRRxJYvM
4wxRBn7haPU1fN/WyjBtlvwCaTj0CAChl0dYxu1pUh10LE5Y2WuDIJ/g8Jn2YJRnnX8kX4k61l43
OTl1Ndc3A7lJwJKqc4qe9X55ibEZC4ckghBIjIDLdBTg0k3XKcPQVzxHLeYS5I0AD6aL84PLBH3u
7nLfrUhnxa4qUN1y9BNQN5OADJ6hMX+l4nKW8IdbmU3i4AFYLJXTm/kkbVJUY8bFA74wl5a7Jats
rLqA1yY3uV8DoVV3J4AxOCrQiSzNFXs31OoPmQqjd1/6DMg0CN9aTaV9JQL3eGeaztR2VVvrSpCc
gb2MGWtWAloNe56Gn6gAbqiq1EBxmxMQanh7387OU2nCHFodLjHhtJeBHbguvCqulQIKlLpjpQyo
BiiDs8N+xyrNuHXW9Vb+ZYkPxVZlQHxdVY8wxlvykARU6WnD7V0eWvsNVio84k2EyjaVVw0ulAEI
tBNK0hGw3Ae9gM9JwH29Tfya38kkQOGDQGFY7MNNfio1uL/H7kjFb/sroUxMy83p+5EP8NlUwnxd
fyzjCcpXFDr9IhTrkmDaKH06SrOU3+BWN6/aU9Zz3MnDo9zPA7mU1aRXINaBvpUTpAyeFD7a1h++
e34Rs2JEJwNMY5M4nK3It1lgigdYCUsBNSMzma1b1VSkafB9QRiKOzx+MTGJt+qwVwO+JZnGayZi
qcKAvQ4NYsVY8ZwPDHkMnRI9BhkJTkJ5kCjGcwbyXb5Uh0WhFvS12L/xu/O/3dGeusbKUZid/2q/
dgLoia7EiacN3c4zmN4JC7jGWnuZDzrx7EFJ7iU3EXwk8zGuH9/0WyydRx0pkgeBUkeAmuD87JoN
5QV2bZCZLFmmmeZV1zfNCoiK4DgCufWxui6C9HOKq/3/MXa877CzrxJEr1ctFwXMwZGTJEwGhmE3
MSfukxZf0o0QTJmfcIF9sEI88z9Fcg96ZylkUxHDu7/Tsu5CgnDwbhhD09aBgJ8IxHzPaXgyzKAD
7GeZMTbiay9zJjIrbLXk15c/y86T4rLnL4DNb0eYeUZaoU+qlcVfbg4r4H5viHBekF3O3n+KLA57
UKWZGYrxBXxDjeusUAMO2ij7+j2M7c8/bzzzkuavEvmvYmxqPFgz+YhDiYIGSPInnu6XAWvMVkFi
NtqCKHvut06OO/vajZYp9qOd3fXpuQ6FoUj8OKjdum1bhDqEn37e4HQyJ0Xf++6FEpyHq+Eg84D7
P2AwsKxj0EtAG6QrlJseqINXX+qR+2LQ7lSlwPRw7njnTfiSTXy/pZxEw+g+jbnq/Scxt95ua0fl
r/NbOStlGW6ky906CL7jgwo4rNqEUQRkRv6TLfByJp5Mu3z5914UgJRtJZN0qoJd1aNnR5bTlI8x
0jnVvY2G3OnE9adeDeGYA1yxI1Rd+oNv7R/1iecrON2rEb9ssDI/S//YSKzJuh+3CtcBPHhJFRcI
N/zE3Kg2o3yslaMXoKxhwE5ibt2XIucuu3U9FM4c1euMxL8Fu14w/8wa+4l6ZO8/KRFTeV5eO0pi
cOq8CdXl6/7DyLWcynUqiUvJ2mGhHteYIoFdWgBVAgPpzqhJCEp4syRpUp4m05BNU8KXOKwsfAeu
mA+HG0c+aovdJshauADA3kApFtm3R9bEwADkhXFPfilDyS4PENmoXi6vtslByEjmWnY8GYC+ljpQ
BW56K4Eilj15XBRvWKkAPl7lDSE9g/EzlHxZN9xGyWNTXUwSpyze/p12ZzobSr93rdIEkk8qA4Kt
VKjawDeyDpwOySJ5C2Rq7aX8avGkreXFvwEWkmtzf7EKCbG1EuEl0GSMj1BaWsdhhrpQjtWrvTI6
NyBW5mTC60P6+vu1ctiriDant96enznS8rikfQyCUVDcxgi2xmjLuYmA7hFTb0CQ1hW9PlNLLis5
K1gurg0CJvaa2SqkSJ49g/cEwVLdhVuEu7Pfmr6JeqcBxFGz40LGPh2qOh9kkoG2X+hrx69k1Pa4
/WAFxF/uOIqjuPOcFTzIrH60hja7c+GcaqoxRIIzA9Ztwub49x8eshi3ehvch0o45+MqmQzeMxXY
gFcQUCdEa6DbDvVL+skV1Xv1iAAbxFzaWJyAbzIMMJGwax/OL0I8rPtNuaQHBTYUBD/mfWe1S8Of
42Zv5k+Sq7tuSR8zIxSybQh9GDHpk2P6CBIMirNaB+5TivrZGnUlOoH5DZG4MLwMHwOrcZ78mB+5
DM9pNSGdT3FnnvogRh3h/xNPdl7/sid2tJpAkdC0qHHr7q99gXjmIZArlMleaQJ8ACoNVYKb9nMD
HVIEO4d2NgpypuJGtRs2nEJbBMWKiH/Mq7GdzO+uXVWB1dVpCl3QFuAI+gVJL+c8LdUpPP02AbcD
ORXjItvRR/0/e2Fn6POeknLMRp/gsFNQVXAJpt2+nfV05EOXEBiDGHTOMATz+tSoEdC3CwJvCeED
0lOpTWkC9pQ2wRK6I9Qhc+aQdQ/2ml9K4X9srwPHSWlqdi4Pv66QnxUTy90yLOwPQqOsFrqPY1bt
vTV5pdJx4FC3wH1JWfCo4cPxZfW4ABDcBJ/wjhxJR/I86gMhtX5/OtksolmUbV/oG4tSSDlaUZ3c
IeVekkouyV54DOu79V2epdljW0fB5zisYp3bOp8rYUbp5byqBYm2iEhi9Wvc3BgZZpRmDKrwRGX9
ctkOMe6b8BE950JHM8LaJkYsagWt99nmEjJ1CK8ZQoRwLCEscPh4HIKDwJrshNNoKqMCUY167iAi
yW+yW7sgp9JA+NJI9S3zj9xksD3/LJr1LBAnNzYnDjJiqgxwapAacaeczkZgBiDLhtmR+BQHuyKc
tYVHt62n5N+TCG4FK41Gz5hjpkT1d4BmKVLkDHJgjLoMSuUhQAJSFswh6dpbsW1Tru0N1ivt6twS
J/46EVVrCxtIRoRKadprKz9uB+WHMSmbv3VI38S+jSXvgVd2Rn6YBPg3jOwRAqqEPK0gXhtqFIpw
KiPsYf5ZYFvSEEGFMzKh8g9usNMe7Jl8mdOu0WHoLoquM6y8fO1Obxx/zm6UL7W84ffTEqfJDxEa
0Vcqmg6C2wJInFXD0EFihnjzBdsgv2QzjcM0XJEsZWFZSQ0NK03RbYH3+8BRYK5C0P/5ZgVjfG6M
9ui+2CsTVge8yR9U7789zvvdiCgipmQsnyqPR2rL4hM4lQf63MljhEbzRYesaCuaW2Mdm+fuCh8K
nDr+2AbqrZKfo9U2fQdW44dRNJ1emgAGrK20oWpf/mU6ohlY1qTE2NsLEG7Xn5NWfJCKrPCppiNA
9J88Dqri7EchkWI77IURFPI9vdhO9ErDY92qbsz98e2Jp4pUeysAxKAnk2c2TMG4mrZVG15IgLoN
gbDth7YiEV9AYW9aOGcGTTss+leICq2n4kmWQWsUvXSYpv7sXNChNmOx54mXvstVo2cypAasKy1x
OHcph2zRP08HTAJgO+AbwIOemZh5xSNPh1B+7673d9rPPS7ObTXQ0l3E1fhbK4grgCY/AQ9VK4HQ
J9pVI9N2KykQPytPaiZLF8qnINjiXc1MxRVIZL0lSDdX6AxPQbw3HYkww2zsxHC1xE+1ZYLkwSr0
c525d+OWkZ8ZpWAGvSsYzR5r7aOdc+q1B7uy2BlY8DvrT5/kDZalKAahvkX9xzdqiKcT3PlOEQnE
MGgrnOYlSrZueEwr8ASnE3sle16l+JbXp74yIA9+XRVnqQ8VwpZx05+cNyVACUeAxSAkLzkEAwfz
jo59Z2Xq8ZdPKZuySanfg5Ah1f/NtzxE5nQj9Rau+xnwQDPV52m/cHqFqUkHLBp/O061opTwP9US
Jrh+uf7gISnY+xR3pAH53sjFoidsEEQ/TjjzshYLaU/hh8mdP6Rq+tHqAty7sEO0sbxvkOuvD0Ow
aD0zWgKgQ8Mt14keJm9Sff0G+vpt069phG0/2GXHIiZHj4UFrqu5GbcgOncCmIOvP9y4QvY9WglU
DM2XdEq0SmoaElvx5os2jW21rO5gCCSMUQGJz75c1klY+TBvA6S4bUwLK9J9AqVCytkDRY11VzP5
HR0X2MMnDV9Fe0VYydmyAT8A1r/wC18ayVhI0SvnJ0v1WNpo3XKsztsiE/WBrU2IuS7E2D1Co+pR
+Y1Lr+OF05JhSmOAcHWePhkcZXLHGiEb7rtpgsMhrSSNFDVCD55q9yeErBqWSX0Hvj/ovQGdreIo
X4J83qwjXmBqVd/Vf2BXOkhGti0ZoI0cP38nqYS8mcSyTXh3FNq1I+g6zZNyIOdK27G+8pblmxpp
NgZEHxBpXx5yFPxNwlwjSCzPIUKqKGPOFXhMt3lu5JPDeKyAfgSXzNdfXWSXw9RzH/qAMU3Fn4hY
5ZZhVRRwweE/putrmbjt3iuFIyyw3r43pOnWOL3VRLUK8A3f+rNkUrkWp0kPDDmGSVBGkiiobp17
W8ifeXmFt9T9663H2hbuROBbJdagf9HrMqTh2tZtHhHaIYXPljie15cUGKqSEQNdBlbXOnJja0Ut
cZRa6VfPGMgksjSWyVCUwEAhijZDTsKGFerHIfVF+BwRzisyO8Vq1GgdyNrWuGaMZl3B7C+2T8ie
w2Dav303HntOk+hsAOYQMfcCmBi/Dp/NJ5HbB30Quf5tgYdcHeCQ65NUNMj5YKqp2MID0zdtn5q7
UguePIrl3eF5rc6g2JUaZk3J8w14Tpm5SO4YanOsqfQitkIrPXou+f4aAGyIe/FmsBJlIKPbDjE7
UgMxogZQbcjewJP19Zp7gM99HakdrZsJdZ7311t34WroSICM0bkh1r0iG8Qh31cgctlnghgA1T5D
ftvEyiWRvO1h7Vu5d9baSCzopKF9QTlzU4Od2Ej4rVWoVUCC3VQE0uIVVAOMPo3gZvBkYRE3DAe8
vUGFVYQynI/AWDput1jg+tsfXMJSMg/siGlFIcnm2RmqiDIlvdsf9PGHneN4E7LrY5bOVqo/pZlw
GCGlk1MdvQe+o9jAclSJ/yOywTX+E2ve1SepNYKtCA/MhTNGqfDvCF9EawIOOlCxtEDHV1KFsKO5
B1OPTV8OPUy11bUmnOrcnzIpemYRHTs9mWBVYRklibvXDaDYABtYxTJnXKdB02Qz9ftLnoZCsbiM
aBCOfoWeLjMMOyOG0UPd4WuFrojNKllgJ5hpdZo3VUTVmLr+JHfl9nrTSOKZ+xtMDV7BHRla6CKt
/4IkDrsb1MlGs+sViY9Psbb39InPT1qKMKrYhAg49IgHHGiHtrdybgvvHCkXzHUFn2U1jFvRpFY6
SmIVR2ninpPvIMOSD4sHersqOdH44Hvjndh0WxriAEHUPH05UJ2rB0YBFv2FyarQga7O1zIop5WF
8raFMC34iin/rUcn0SpG5F1QoQJ6QhJo867CxtvuOrrvp/kWDo6gE/zv55IeYH4AAcETE03ueAdZ
qMM5csp/B3xqyIakL+zxmAfkNH6ykPmxptoQ2701pTu16ccLFitQrA4XBjSV2yfWRQh2pCYThmFC
RqKrIGW6nKbP7TbMo6WobT4KV4rosl0okk3unja+a5EoiJt52GaRqxfdx/91Tj2zEUURFAMFi4X9
eN4gdsG8zJfGELgmgpuMEftJFYQtlQRkh+kEdJpsFSPdm4/zvsw+6gakqzli6UHsgOaqLn7tWYLr
JcZCP0FFtkDgV5xbu0bWPByPXSfDC95L+tDOmAeNXcstRUPXy7762zsbXj+VLiIs6DtaDcsbIaBH
P82QdIwUcBlEUZvSFgxaG8Rc/Cq2ZJI8HmXcrr6wanXIB/46ViIRyBMt11kZVmIQuBXlrFxE06ng
6o/2ceURaFtFKL4h4C1bzsDweyiWfWi6Q3SW2p9VYepUBpK6i1XHzOtmKr2/mJlzWlcMWVeYsb6P
eNp23BozWFS5j6MCWx2Rxv+fHPX9Ft8Dhu/3NEaDkQwpPGNx4NTZOoH7IvFi5DWoNSKaBbX/UxfW
4bdg3YFZmZwQXZJpE/6uI8MV5qB/tr1YWVagK5u+kngwmSSKPrgBhwfRGQztGuiPzV5C5OPCumY3
jatwFAym/rQ14gA7b7Xn0Mx21exZMUAbNtnS0pOtWhQLBD50yUKeAEx0bncyNI/JWCu9QZfVZsGA
j2ZNMyyy3MkjbGdwMLWVmo1Ve1lVXnSSzmOYVipa3LVarGjzzCOH+DrhZubUopVJFfDxfrlvn09s
pSwLV8JJ/2emjGnetGVFVbMJ4lV0aUyjM2m6XTfNMy+DP615BUrWccShVYg/d2oTSh5zqq9XHhex
tX4790oOdQPXbvgQcke1lbBHsFRs8yZcYDgJ23OiQDvA9+mOWcvIUaaEeUR/1WMXEtmBWxC52gFI
AJED7n41cJXScOK0ZNwe3zCFOrwI9dC37lTArUW6oCTQQRfS1btU8cIw7C5OXv3+c5nJytm5Gbv3
HaEj5ZDI+bUStaY6WuRPGQAf5yqu7apkRf5sigE/lh7njiYL9X+In/UgyPO23QiL2BciU/2cUrFM
8mh2qIYtQAyFcpE7FYYDFRkwcQKNvvkD2qbAJQmTl5ckquELwObH9SnUCW1SRE3aQXGAqIhEJl7G
+w3fdZ5cukVB6nfl6jVP2aCeyDe3Tbmxjb7flCNrxz301ATKEttEtaGbKm4uG9k2dz6g2yhqZHRV
Z/Cz1eeAIMHbXyxkwungBQk+3KbCpuyyKUlInGQGUSK3QIi0OIa38JfJF6zjJpWas4KZzBm+7PdX
BEdZ7OQuav+d6xpWqjsFe7sudQU/vd6ENPTP5YODPzMWUMG2ecxGjYHjwbhUV5ogRcN50k9di+FZ
tARP1uOhVlEkaUv1Y8iFL52L7ThMDORfseTEQl7X9l0mFYHGemHt4tItk0drDGND2yqodX/TnqU7
RTU4QDXzo1JltViyKeCyUQX6MEQ6EXt7kW0W7JJsF5+wel/J13n/iRK8dkVEO/X4A6tut7hg06NT
wBzp4+OcQozZRTF8SBQtOYrH/XzfNPYUXNaTsjwQvw6ZqQNGT29Bg6HbxB9tMZVWFoOe8vKgpOoQ
eSwkbd7DHXzmETrzOc+Lu0ZQ9Dj83WIUNiNy9hmcRGDdESXUKoxBXmbLUR5GGux8+7wqTQMJs+nq
vzXxIzMulxbmw/jr1zvI1+chf6zaaJr/zwt6I6EojObyv9r9xteqXCUCGnbgyQp1QIU67wh6+eDa
GX5LjZymPJJGDxJ4o4Kh+94rg9g0IkPA3ACylQnQAFi6T9e6Hs+A5AaR3uL3Zj5Z6ZZYHdOUkIvo
TZHZ1L03/z2YdshynJpA57SXslUCQQJ8sZlnYpwcsTEGsbQJuOdAhPbiFz+fnOZM5WnDqZWM08Lj
79dqQ/QP6mbaPGieL7LoFZK4jkpDYqnJQVG+h7gsgnwiPT56hCdn+hvnm6ehE+ynJ4x9SPIm/0I0
hs3beRcxriLPhUhpP29SOoUUwsu94Md1FK3D/iCcbL4rL/EhNyUcHgn1rOxePILmNB1iNO/lB9po
rKVFOlos2b92mf8EB82agypJJFptNKlKvf39WAfRtV/UjbHl55CrOzFSSK8A9KklR60GvS1jK3xT
b9rMQ8jXx/O7fzmlLVqpk7DZl7DoPpUKXKcQOG8mvOkjFVkXRoN4DE3hRV2sNx9Xz8/XS9WoChSk
8GY4TX09Xy/I6bNsmW6bXVX08gZqUemFSQtlQEuGNA9xYGaHw3lQleQD9xSKyk8BlnwqgEAph9Qg
SwxUTIYGn3gr7FlbqnjboceXR4hL3No8TrXPawgtRGHGVLv+Il2tj9aq0PkVJzksw1D55hB8t9R8
DGAYmiOZBQniLdPyKMHbg+ZDA2NS38BexVNkfwppzoYIS2HwNKHjD/4n7rvztxctnmeECTLTtSSj
Jgb5V/YVzWELHMN+zFCGgUSwLc5/6/tFmAZRefSqk1u6pteUxhPxdCvuxF3BF3ZKDnT6Mn49ygZy
EdhFrGL7Nz2OBrH1mT/m5dbI9T8Iyt7DfI3EHE+Hq38ATGcVDX0KDOpRVhB+X/hQ82gSRWR8QcBU
/3Zs8yEZ1AUIzFFnMkt6IADTZiDHHl9K4Pf2mSFyZEnNRWeaph+oIJi5Qs9PRqCBYmwKau6+2Obx
g8dJEbvMTHWRjm4iPlN4hFLBgYWYA6HRAtCFzwkg1GmIbGW268D6/ahU38U2weirNw3wBrkvwe2p
wDSRMcr0cqqgnxd6Ocplycays4Qfb6WvtNIH8t5sxdxfHgGSbamThpbSntZxjuYFKXDR1/YBB11N
TmxLEXk3HR1dmkuOQz3C+YBikherWPTdaLNSQaMQi8WaRYV+udjpnd8I4XPMHbvzYf4gZvBl6iKO
SLtyifY3hUkA9vH3UAZnSpaauXdEavCmYOrEVv3biHuUK7lGG0foxsw0eGA2+r3GiSFImpisL+W7
yBMKsFqMhomM/hnQtMtWZWnju7viYnwr3utV/5HDVV0ZkNZUDjGwRpP4UjsH5xpyxrrtESfmHhkN
YIOKo/Qjqz9G8aBswaQYBrdm+T1EVKZ8/S0mCY5oG5Ovw3NpWAnSfZ8oSBxU9Wmcj/5pLZhMOr6t
iWYX4zXlM5EHaIWVn4NnPiNSIp1B0miP9Z4LEKznR4j181CWxvruk6Y6xKc02eSq3IYGlYaP7Du1
JGrhLmVrKd3XR/vxmdvwLb6lNYpdmfQuzeTqS+xo8gTy6LHq29zRwqcA2nAIF2i36EmpCIHEC2Bg
S6aFpMcow/m6+xMRDq8xyDBKmhdnbM3MSla1LikGKLFOvKJZaGiXEnD5iTxIdhlehNjxikgEJj9/
n0m0/x6n+3AvDe/SSxpwHmAzgBKGh2T2+qe8Pky5ovTD/75vA2sb/lDvF+KQzbpaYtt3QXnOld3M
JQAG2OZ/IbHkXX5LNS7+CU+vpTzalDnGmW6LdqDtAE7TaAZe8jGzckV9XWhE0z5wbL1PwKnCaSPc
ioql3D7My9SPehgDXWzQ2lJMA62LKrux2/jw1goxu2laHIXk4uZmDcFC2ZysrB8+11yiLe25hk+q
FP3RF12dg8sOk30HWPAxJPCtnc6d1S7RGhw8rzymWCRcpXfHMAblkb4FOUlopRr6lA8sf7hXsELw
tksf00BE8WqRAYmMrgCgY1js+lYH7VjkleVR4liFePEltSce5Y3Vpxc9eLjj2HjZLkJrT/wv+GUa
d6H1KhfIZqvsfX/2ZYhsRj53uSafObt5/LnBwxvbVLlwMyqqosicvk9HrhyN86MLdfr9gcWHvR4A
EjB0uZ995zdiufONodoyFiDBbGQ9GRXCCVvSIMAKUjVD0D2dxCs7w03wXIYV/nNb5z9u5vXbnQpm
oMNHNu7UYZ9fp6TecjsGEIhcBR7PQScd5CYRlykQMqS3xqolfoLeCx+Leg7k/0dXbcMq9eW93z8a
4neG1gZTjyB9fS/K3IipZTcsky9d18YIO6Xnktbt0QOa3MMVC+n3PkWpq15sSSqi1JuBlyIbEIrO
97m7d2fXPftC2nCLZlCk14tOcIYPht60vttLlwhuSm0azDYEUdMdCnlOZGwZ5bMgpvvtoR9pyK1Y
nb5rnuT9fpTI6dWtx0UplbOkEuuOxMn2T74lgYG9EsT5MZG6/4JDbBnWoT7p5s7yalG87IqIludL
tuLnPWXEU8myjE0LogO+3Bf8LOyOfLSBp0ZGr93QamS+plxAGz9OoV3MIuHG4GQj9mBa/MkziJ6M
yJ/f07CJysVy5NCRsZM/Vb0y18W/5+3LGLcrW8iMcF/5I/cym1tJF8NAWZhhsuJ75yjZL4jx/mTe
5yoOvMmW+ylktGttflGYP2kP3EQatPCLz4WBMb2PPJzNR5GYawnCOUSXqY2tsoK9/meQhm/Q0GL1
m+JLDaDfPWldtoXkfJX2UTwIHU297OTTERT4eejax65LIWjnBIKTVnRf2x0/TndR8LEjr5MiaU4U
sexc2/BXxiz+nLzlQcWR1eVlAZtZ6yMEzAx3x2i481Z5AcpqqGbM9OrHf58geYB2R6RYGM4VcYXm
bh9W0u+MuTUPGEHZkuNt7g5detHGwCS3Fzau6/jY773IXz6IhMLe09OxXnmmeW188dxcinGma/gJ
s94AkFKW0I8mbJG0zeuvOBFjVM0nC2HbqxWOVz7jsGr/vRB+QuyXDqAySgG7imOuVgxwJxQ414oI
xmgKTtSNB2B7moXwQ7b8baTYEo6yRKAdumZGKD3xJ8BjFaFPDFT3qckeQmX+AuIMwPtMSjjW9chK
PN3gIYXp/lfs5sBh01iQ83wJ4lGdaEqVwVoWRZjElDJU8vo//uRzKZV47cOFtZNi8GSU8oBW/gKq
WllrFb0ulrs4jyWKBm+FbQ3dAj95H4CGjMc1haqv+/YV4r4cIkXlsPXdwkCJS/18pSOkTpcS59hp
baq63yaf7ROgUF+ZVMWp9OwI+VTDxAChGjIesBjVFZEne56rqzfG1RcPd5HpBrBeli7/Z2qPXV+e
KWmqesh8brME5l2rgBQgo9cHQbaqE41hYjPKbCF+SZ0dgNkAAPOdOFF3q9Et8iLk2uuXiCW/J9xB
NO9LFtxvHnkmi/nO5SAcivAUe4HORX1kCvFWYKogv1scQegGNmDUHePWpygyo9Bb5Vp7FvvDeUU5
SqrnQyX2fveACkvecLuTmuzyf/wn/YqNMn9TXJ8DwXAVGCO4wg8IALvY1ZoiPeBTw444na4K/YGq
WV/77BpUn3oFDNuXwSXVwUTzTET0epcgw16yarr3aZVEaKu/WgtkG8GfSoqn+pGmKuDjFn5I0tRF
MTRvVHiB/XMqko+6VTJPXAxXmH0M4vR5mAlo1j9ZSo2WI9+AfklfGaOWKm3yHUFqbmsjllf1FS2+
96dW1IQB6lzaitXUqVBFRqz5XwzGiBsuVu+TQF7ZSI+eWNqK7m6cxKUB0QfkN7NklGiN2GdmjNck
KCQj8twy0mS0k/0TzP+Ei4lZdRoVCJ07zoNMX+YyY4irMmoktCog/XceRs1KEfVLh95NUT0cCprN
B6CC8pCtqgmQpz8EszbahGc5s6IruhCbOxFTwXew5qfEhUlj/eH1BHJ7LAQhQLdOSp+U3mjuphMi
wGTBX5E8cayz08mhYtuBRJ7VUZrRUkwoewbR8XRnMbOrxpCwEHeBzMknPiKsQTHVy4Fg8Gythj44
Fi45zfbGUNedgL2ovCgqF/aez5qpSVCnm4qPjjf+OF3XvIv4CLPSEE3I8FegqC25FfObN67WqLms
DN6ZO+3Ld3XbZ9o0RJdAN37BIJKqyi1VNLMMJFUz3kRgntV1WOg0DUD980uTT8Wq8EIlunu/sCmu
5Gnr3G79iYcjr61S/leLlX5pyCKakgvnp3UDZ8stViZEPvQ/cz89F7VLv/e4+KkkgJIJn3YweyIc
R7g5NmVvzMaZYqFrU9BMWZ2JoNqwurbyEEmCPJQQYdnHT6VsauUbxZB2PXOLosYSZJg8IoHqjl14
jHgomaRsNNSi4FD6e73/FR/VRaGeUUY7oOCO/MWt3uDKhJEt3A1fgYDeg+VSJ2Qx69lNfDJsNmip
KD7F2uv10mAAVRqZeRZBq/x95Fc0idfdWn30Vf66Iij9kBmsPIMhvWnYwxI34hgJdkcac8X1xOcb
9rL9kl9FP0XcHiV6Kuw9S+ZS2PalWB7jIUTzH5W1CbqEdtHHuIiAS+D2v2jkVpqDY/Z0aj0ynH0q
3ztgHHxEIHNW6Ew7Csu5/PZN5yjHRStwE2Ah+hooNzPH1ZU1J7xadKjUo4FS3XIjwQWvqDlVrYRY
dsmTo0rAu8mE66i31R4myy2X5c4+BezYmGqHIa/C4CBcovrOrlpOgtNia3xV0RBDrWpnhKKuh0Wt
Qnmotm7GPPLo+mykf8UjDMDP5pk0eNY7vRwczs8p0s9wV6xwD6gvTVO+vYORyGgolcUZlVIZSMDB
u4k7roXlekKfbKn4HY4D8oStgcZjhZ8dWR1ibsXT2LusWMc+N8q22S5cpbAhzc3a20lEuBqSZJcd
N01mtgv434Agr+QZkPU3nvaanDp8BGFtEguXMKZgs8GcY2zQ6dGTKKB9T/w4W3O9+AInQl4JWUbc
LB7XWpbRPyG8E5Yfx2+hs/kA5iOMXMAOexNkGOgEeMcgUx2KaZuxj77r8dEB0EU0J5SAmJod7ihy
ZtbVBctsGjG1YSYM3Ttq0fxiU8tKCFvpOrcJLTdoU2TRckPnw2bUaNlzbZfTjBD8rSEt/806Dlcs
22Y3fgCxO00a6sUED/h6T+GW5gm/uZUpJER41RjKG6QqWGxbGlqlqab+zFQVMqR4FjO0FUoZJmaL
r/h5wMPVlzo/qYFcjYReq892I1tLOQPTFNkOmy2cxMhPgojlGjwZmRGBXBCNjALC9+QvLnmgSZUp
kLGSejiBJ9fQLayPjgi5a+RHVN/U3jR6KGTGCZBP7OrrbwyOs9zw5tE7brvS+OQVr4T6hPWoiq0A
IrCRyCILhrq7HN7KYfTdr67+PkD+SmIeqCG7vEdX8/MtSeI9K9Jcsyu/aS3bJ0P813SqHJiVvqjj
LG2Fg+Q1CzsRxH62ZhENUTHfHXBPM08NRqZZyz71v6g2rPEG0nmEorYQTg2Vykq9xVeQ3zCnPmad
67tTzoXId7aGgfFT90n8EGY/Wga3t/DSBriJ/Fxru90zA8nXbMbSqjQKOR2H6oArOtKssqf5BhQZ
gKlbmFMU25IUtJDx8jUTrpbF8CBl/wHvY14LRK787gQfUI+NP9lIWgRvxjkhEDrjBlQwlPNPoeWc
wbm4RJWzFoXJZ7V9pqS5Ub62e/Mi9PJV8+n30+PUgRwp1MXex39ioHLjPDmyQZnz7mHixNnAvH7b
JOQRci2ehBLtkFZTVYHsC+NcSAnSRLXC0YI4y7M2rJU9vrfbvdxEjMn4SFjZ0397ShMFDUduPG+M
jFzZmKS8RwkmqYAFPrP93aYMH3ye/Q9d2xsKWe0K7XsoqZVMTsJUr3zQF+j7TGTiMvLumxeyQ1bo
kdYcs9MGWe5PUxyoVjhfRu+ig8ufLY+DA65CaE4wQQpKMm1ekSMmgD5VSkRQIauQyf47a0XhE2V6
3s83dmpqiiL/KUzRxPL37a27GDMvzM5hnEvtt6TTwZqEvRxMWJ3q2V3tLiNyJfXnVMWpzoeP0MCm
yevP4EL0QRk7CeLSolA+iAIrpb47ZiNqoS8KW8BQqvx9oWX7qJXQXEfCn+VE+7aptDLRDFOOQEfb
W1lQplyTgX2NeKc3eB8Yfn9J9qKaPHajnZwLhQekKV2KxacbHTdCjeFbNubro+VwQUcKwdsYiZI1
JjqOvKeWajqxBGud2/tsac3yASRDxl2m8p6ZhNd7IZDcTaIc1j8Ev2t8n8rxshmQIvhzI9gQrvkl
LQ4g4vDh2p6e6W3RnHB68ViqEE1/53u/FqqKlhzHK+cshP8f9QlF3J8hLQIQs2RywbOHNbHHR7ag
3K3So5G9cJXfF2cWidF+0GTAJMy8oIpBNa7P6RLqlgowi5hwEgY8P4Olk98ZIH7i+6LZl1r/naLn
oOQR94bxvWK+WQtVd/ee1ioHbOQFRh7yhB84XhvOIiAUkqkdtTXicto1Qof6dcqMY3CskueDKTq8
Lhh9R17QKLaK5KHx++hRurIqMTu7rWH4hxTYMhh1WQfvu4PituMxN52l41Ayl+zkHH0E0RClXN02
E+dObmZeAA+gNTxdEax05Uhq8d7l9hIsDw7Ey4txIY+33Epah4wUJK5lDo4ZrjtqWaOCvF4H01wY
Xua3IwWxAU4T7trXJNvGFh0KOdFlG/XCXaa8vH2U3WWW960rB8zlERIp7zloOSYJMIyqNBasAj6i
qLCoDooTMY2QgUSr8ul0v+MqTHW6yZvkm4Xo4gedtqsDp2NyQPREoJS6xoV29NNp5q4j6EASKV8E
1rUwOk6MVRSHI1EcixVK/odNrW2bYER2p78e1jZQNnP2vb2CaZ6Wemu961DNsjYoAh9pL2p55NV3
81hEe0ly9Vp05Nq9ecbKSlVZkLYooijUxwX0Xu9CPUpiSSahk7xBN9xckJRjmY+Us1Bep/u0wB2n
/J+GDozei2shtw1IT3bfmRNw7fXVGBILFyHv0I8+NjE1OH9XvQm2tple1uA3ZOJA/vXr6Y/Da7t0
fztLgHQpl3cCQ9TNBRn+AUh1IfSK1rVo2jT+qvlpL1FgJmbmrw0QjBJK2T0L9mFWnamBgR0v3qK3
kDUEvCTx5MEMj+J8/DxnKOUhUMNwA61SOqU9gg9GNRuEJUolOfE4MVC3Vm7xJUe/dINyV0ci3C7y
k0yBglRwOuqDtqawDXhhM90S41MSDZq3TYWP6BNiFaVKGXLa8NCD10GTc6v9Ymvg0O2gO8IppxLA
O+ykmE1zj44MFgwtVwEH0X4tiSQffNkTC6xJjDBTVVQiqy+Tr3Ebgl5ovWPCpbisOhT1TCEbVrvv
nXJDPNHtfxsuhgulmv62/Wp7ahfTTZ5AL2h6NKCRWbJ2um1rto1jiWPVvAxHirgnKPS/lLIvzp7i
EHyVinqfnuD3Pvd42W225gLy0b6705Ko6klWGbeDqbqQSkxeLJiqA2RhYGWIb/lEwfsoR1HzS9el
1gGC4GdkoW8iN4dV+PhtYORbFQz2H7vjZSdbgWbAZ8kriQNFuXz/D0fKnr64f+H8s2jjz/Lo77Hk
4z6dd8rUtQKpdyxKX9HA1Yj2Q8qQ/Lunluvj4T9Gn/f8qiyMsuHSo6lrACDWTm6O7BBupPIqV49N
5Ulg28TIVgnjd2fEekzYOwhzdEOcfR/PiGhZCtw1kt2xArb4VGf6c6WHVzCQH0glfcb7t6biIPH6
hjm+BhGpC+pNf3OBnFDxehDSfNQIhL4dEbHgWT5svkC30lGxNZdgOY72s5usPhoWOJYKtkC++JjD
WXW7pg0sEOBxg/E3+XdTL24y3XzK8xFg/r2p8wE1rEkJEwMwooOYLnpUw2QMNARGyD9qhOSmCvKC
b/7m0T/7H1Z+blVUSnghOM9dNESJTpfjLi8G2DrAJHgtOp4569DRp8BYqS5L03Nmrfat45fX5XeA
b7RmO0RAtSypnq/KPy1AJ5JgZC4Yp1PnlD0x1nsyUJ+diHXI535onsaLqncH648XfF+bT33dchpI
0aKbqeHT45tevq7Z+X41fO/SCH5LADebRSEPcZTlfKI8H38h3rz/txtM3gEBh8h45uUCNcQjtDYv
3s9/utUaiSZkOPvX7kznC7upEDyL2sAZqCW6M0TJG2yKPwdBKqgEkjV6f/E00xCQifeCFwFDcMmS
mnkyLMxtIkc7HfhsNeVsAixaR1szAmS2NwYe/+9JEtX67iwr8e81WrPpGGlyYbW2zPxGX+lCKg8T
2kDI90/+AQAL8uqY7GQkSy9Ztp0RYjdIw96vckXSGL0Vh03f0athETyB2faVpAq3ZDMAH7OxW6T6
JIZ+Ct7h2aYa++MV4vN6IP/XmLrBQmBCt9ZK8lp5/yeaEzk8klN5ltSXb6QgMB3LhOsjWU7L86iz
kfIDz68Dz5RbOplsOSOv2gUeCeHO/NyNzByzF6ZJhhxA0eUEUtf5eluKytugfPsoqFJDFms2uppc
EzNi8oXLAIVVAz4Z5s/N9dknnODtcI9KaB8a4AGrKJMomb26ezVy7KeZY2vm04GcwFhE7ugSjAwU
862AsyCYO3VCGZBkG/sBCPT/cikxeg+2XNQMA9ohzLPfe6ROqrXBwnpPoUl76p4eTIQPvr9dFnBT
djAFI9cOIXSMqJMkBoPhUwiUQqzW1UScJjSD7fkMJI+WV3ElY0XRadJdv7zorWzTlLsNmiynghJJ
qh2UKwz+0RIkeDGEe/cBhpA+TNNqeBszbVPFO8abC72WHsVUwmktHnPXdaW4cise2940QWbBpiCD
eFJ1Qc7IO1wTGHB7DF2GzOIZY/GSpi6nEd/w3Isas3UBXd5lWszxDx6ehmpT5oaWbmZxZK7joOf3
JwJjmJ+UPg4JY1wjUeqkPrkpEsXjCqR8Ue8T1xxBD1rN4Ka1+lEpRNI9Rki/knzYmvN+hwWZiCfC
8BQDok/RGaohCRh8SR9hGVatBv+zOOTJvESK9+BlaxcekAZGPuj4tUss6hdI5PHAREzyfTRDA2He
LmjOYrrDDp9FpMOlM5IdcO5/dQdh+VWDE4HUb7fA7Hbu4T/Jxn+Q9kOgTLLVFwlCR6WGPh88pTIM
TenwfGRMW4l3oTg+V/IhAkjizGtoS5LVYeLiI/7i267hQS5qfEGzx0Afd6dOFiq6dQyJ73+z7DGI
H41xiBak2jezHmNGeS/wwdeFiuPoHKLy6Poz608FTIO6+m2nIQ+9NnhDqX90v8oNEq4tHE4EIw46
wZsfy0eNirkpbCi/va/o7Ox7c2PohsSyUaMeF5zeBeJPPJJYPUIaz5UAS/lqeGhTrqUKS2kGcYnb
jvaRig9vzl3MxcDhxawF0hWNfbtqkEG9+aS4DXC3ES5G77tQcatctgpp2uMKpGzmDH4KHGfy+pYo
2i1MRgoJlji4sY4iGEyMCqV3YqSUnj2nZOpvpfYFnlnvlXc+RJH7e0KYbHDDcgQqXFOsy+LGm2z8
Bo9nHQXBns27aeKVqvszQRb0TPY2VR2227QpGNouPEfU72yncD7Sj8B5doAbpCDFlsGQr/sGJlxD
ZIwJAG18jd8v6yu/XCFCmS81edgKwCbnivN2I/o0ZaJC82PcnWhbG4eZIJ+jaRbLVGev1uDypEjk
gg443dbQNUI3kdUOACBYu+Jh25VeMZlJTJB0Z/wp9CIbYfWaB/TLX2Ntufv16/pmraY2ph57Wzzo
nYguP8P1ikqwmwI50aAyGNuTB2PiBj4y5i4wmlrsHJVGYJOUlcD16N0p0zcOiQR+7NAC68PJtXn9
ZNWQkDsnb3TUUoa2THdWkB0K3Wh6BhBFnVvgkF5f3gpfcimQk9Vz7NsUw+XuOEwONftxBiC5v4KL
9qUtDMIuqZ5pPSYLknLRLHFKQ3mZ9oZIVy/v+khww7LP5VP9E/Gk/XvuZRNMfv9EwgQuRnvWQCMW
v8wUmF90opm70KmbeRNFEiXzdC3XS0TbeIdMzlQkChqhCoLAefsiuSauw5HexXh2UOK6BLO6Taty
sERdS5YFt5zQfB/Cz6JiT2hhiA33pr8AV631H5hYeoIWhUO0MOmXNzyvJOr9/3j9IjJoslwR511s
wkpngqmAav5l3Po9hiDkt+CJgwbKiftcaiQwFaNJetx72gnLr/FzN0IxLn67ymuLryJj1ctu0r6w
gFXR8FIbcsgYQTkWr6WQGG5beGO5Ew68qEeX8Yyb9E8FGJoEVUXR2ZxoVTZ3JBstwjrLcIlqlEWF
OaDR2ErOTnK/97RNXW6jGZopqOzrZMmpHQnvhI1gz6uizmmRAmBwfyrqQYhlt9N1WI1p7Mbjh7RB
nImShq/iiUCsNBrh1L+75xDV76MKsYliTZa8sW/WikLAt8KIW9UfHGg4g+n060yCC5VMRESG1z+L
CVRIepby/VZYWiSaXnv1rOpSf1rFBImEqi1D/i9Z6YtNap9jNr5pE0Dl5kijU+XvHdffuYHAreXg
14KBSyELHYAIAIYTLxCCUbkFJK212bK7oEhzAqLKwQE5k9jL+xGZ6j29EBvmCqqXCaJ07csnQqsE
Sjx+g1vN79M21TvDTL3T3tX+abhYMfkTEnwd7U0KAZUpVAtzZL4FG1KxR/epsDZhJNwqQXTGWN5c
ij8tduHkF+I9MM/MV3UQfj8PgLiGpnkIqQDpiq0YIqvSNQxn/D+jvrSRl8JGTdVuFbc5TGwJe8Iy
PByYO+jWraSZQ9+ruz3Xb98nPuqN0ccsJEidLy8Y98Wm0xTFzlaFHosYje+oHYtBmSpJqIpBE3FH
7hvbW5U3c+pkftuZd0jxFXMVor08DYRb9cyj+z7OWuoYH5aGy+iKoe+YOcH+wuWb5iK7ebvJ9ZZ9
+L82Pm05voH8D/BDnDh9cHauQvW6IoZcstK46467A2jwz6VVF6uJlum6xqxUMtvisPQp0So/84BJ
OCls6tkJNUPPbp2P0aIcJu+7mo8tPtOkMiDU/qWKcT6U45VzWkBJLM81qvvskmqAWcIss870CmKn
7xqoto+6yEKpf/0osXNnCsHixF1/xdw8Li6188LelYq8gLi5YgIgVa2Jeqt6Pa7TdWSNdPwE90ma
GEnFBShaghoTwtW6sP5wWnymYT/1JGrWmwtf+MMbwciQBWdY+rrXsX6+28AGFcPBwWn4ehk0Iq6p
YEax3bzf/GrVmn6J9rwGV+oCk0nuekr8wZWYi8UKgkjMxIEX2twaWje/0tkjLVG9ngWbTxdPHG4m
veqRyGJXqNFRE5xzBAfv0zRJfd/EBe0b2lNF1rhJigj8Q/rCb2YgCWo+2svUdVXvKv+EMA08Uw6R
lqkYdYnO+210prWU26hmEEg+sqTZs4phZQxWtFIzSgMvpr7/nK+rcGVcjpC2+w/Vs8ToRUT0oDYh
RkoIahmOyq1Dzo+lj3WU/2p+A5mDQrm1TPSzH5kFjyosNoXG+Q6NA1q0YyW8bp/1Vdu2ujlCkRAq
OccZ8tNUU/iiDQqb6L5YpIs91mY/Q90/VVo9ke6loPl7YnMXm05MU/kefwI+qEdbnz6Qm3UV33Jn
4+FWz1A/7pog7M+HmQcHmJaCwESjNzdfHJhHAjcg3AH2gIa3/E60/VUMSu+Pr1LkzfHtJUYNDMtZ
5frFzvvdKwLj4P/zauexQa3FU7mKCKu6SyL0XE3q274NScmStB3v36pzHM7FlpGi172e4qAz2WRL
D4AekrNDW7XKYdGoMa6JoMc4/U34AXLG5TCGlWFjO5zEakq0M0jnUp3eljByLabAKUocYsVlSzhG
sRLamj0FL6apzgJDo88X/UsDYbpXZl8ue1QUz9gDQIviPENfkWsonJUohkl7OqzSiA7ascWPujGw
BR5NofxA0YxkRBYWsKlD6ExdQ5aX8IY2bdeNFEOAkycu6ZMJRXc5EV9w9fX8KxHjSpmBuCQZBrWt
0mgZmgEqNRBpFtPwFl8XY20+mtZOPvTyJc162qRnWCmRTxNFGoPFpqKrGHGkeGd9R2aGr3bV6A1i
fjXyEdLRnE2QTQ+WiazRRpSzYHDp3M1MkUVerUtG9W4VJirwVCWZWFHIJoyOWPQlxn0kLtct0z7F
sK4E9XdQNHtbTXZiVWASG0RjF25ORKp1r/IvagTSWVNaIgvPp4QawY9Bt77YZ++UOxuvwb/JE/0H
UzGxBroNtE5uGhJM1+d+mbk39DCJOJZSPN41upVX9GqK98I9bXV85VpHhUqwanwzWJ3Dw64gdXU2
xvWNyqSSBbbW1/U6FloTStWGwJrcxIE4K/tjV3nO/+D0ClTd+fXqLRqyj2DDrpm6J8fRak6tR+vT
gRUoas6Pv0addpBEjxjRkzhwvQrzdkeapap6jsbvHUyAxizVNiZHNUXQpEvlZXQy+OqhbHKUhG+A
NcQGIBk2HmXK3AN/KLEUOK5f8SclPW1XBlJ13U5s7rC8pwNgYnxoV1k3zUdFJNLYVgP1VMvSmLqn
DxcklncXdY1zPXPXvBLNvHPnQ/0SxGHFUJbLDYBG0UEHbeDjd1wxn9MLXOusA2MQptpvU7Vhsz80
AQKtnqTexffPVcAxRpDg1C7Y7Np0pEtDR2hXEi2Otqo7VD1ocQoIVePPn5ls4wJ2JPzdLGhjbwGm
k16e1HeZeSGiejNFonUzbyiF6QJ8AOKl9IaIMUEvwgi0xI1tlN1gfNZtFaD+u7sjLXjau/X79cTO
xW3H4Bd5ihO3SKwjLLZw2HlqiYYJj2e/DRXtHYJ46Sypia7pcJlNYgl/EVgP4cIeukylotVi5pMw
y53otBFRse4WwmjBZ4d685YC61bxtHff4aPX9LwoBF/fM4RGhcPgOuMUfeDROvxUYZ4jvzfGcsSu
xOwIds5W02FcET6jNFlzKZmUzGUhD1yUNZVelB+YXTmPhGMCajuYL7eaECTwrwhSf0RSDkjoB2HH
zRZNtnHJuPob2rn6bQP58D1kG7ayhWfTKDuJRDxOP9YgR07G9fMOL0GGbb5O/0q+DtTnJggDX7Rt
o7J5kBq7UgvBrZRA8FHHY9cGaG+X0Khwsc0UMRjW8nJny5GcLb9R8MsEVNoenwYkC0k88awy3MHw
up6eNj2ruvCz7eGiOTh2G+6gHNjBZwfWZySQy8YWA6/ua83dDkRqbOSvbWBGiangQxQ4maAk2mE4
ky1SGcVyrQ38KZ+8IXAVTYx4Mb5ILN9+LzpPxVZ/hJQgFtU1NrRtnHXuOWQwXnz0rOC0S9zIWm3k
Yhw3kQi/Msbod63eL0BQIXW6ih3xXj94BTb4SQ2kgX/D3qbfVDlmwcPJynS9xXn7DygGrUE+eBDt
9gcNybvw95QWNv8OM9WYWTcu6SDeExnVIiN+SzaJdoUIHCHeuG1kZIkgRAOmOL4Yf46ZWaCh8zLV
THnUiBM2CW9k1bHcw6VQUdjihvms39XV+4dQWJFl+wb6apGVi3b/cspYI6jG00MtJmGiQidDYhSL
MptIF9pb8fDB4MsgpGhZU8nozWENsGwT3yJuVIO5GA40hh8SGJWRA3C/o1AVQezZymnV1EkO5VUU
zmaKrS2zf2YtknZ0m34vnPSx4AlMOngsd9Nb5N7sl0QnhBEgug3d0Kxr0aXwDQnRRMcQnWdFJGUi
YdjQDZ5dtZ4xKtmOgHKpVBDPEpQjDHKsc730i3T4FLu+KuyBxtKL6aLWmgdMzqWQS5zqyl7LCgPQ
9nkkYNxWnAP/KAR3pJxo2IMFI7UnCG/XttwstSy/wLLm/i+rZzQxNavGeQxLDzrIam3Hpm/GYPdK
73GxwWW6643f0nxhR1vFKHJj0/CIJuPfaaURNU4IKyntQKbgR4OmOyMEJfM6LtN6Ba1KgfsuUN7A
vtqvxpNaV94O4r7y6zAg63BOZ1FmgR1tvOsxvfW0V4B+C9EMWynvvGRiNnH6PT/GS0OyINjyxjVD
SN6LuyOF1WiKlgFWCyqAdMdRLqNbX1sBogwmgP+j16NOhSe7k77C+FQ/JfOc6oWuIq9LPu3Oq9Yu
1dMxHKJUMMxoZwICCaXsxB/wV2nvmsrW+mIQ50zSdaSS2YhGStDFoY5PfTZfQobIEZfsPvZaLe3H
nGaFu0NFPCzP/rgmh9gk0IMCz1EyZvWrDyL4qiQCOMokse7xZF5LB6jYnz3RObFfym12QXCr7c13
sG1TdgpDyqVJ2a6i0jO/OjO/Qlf7YjulXQAmXvU90d8L308skymhwEwdp0jUiQ+VTfPVegJUH/C6
HD6Mx0QP8Bp0VTmRSUs3vLBLDmiP++cAp62JNEIQ+1G9kiA4w2sK+JSu3ngT48I18U6CFiufueT1
XzjerIxV4FMdt+mLscG9d+K/esyqzaUmwCKSFrA2nWXE2YK9rP4Nl19DdMPdRxzxWPpM1GxW9gWn
cCt5NTXe5GzIj2/wRwLVDMrzM2zxSjWcZGFGEnGYwLYkZaFZbVapYVUS+68FIcd4IU951lNnjuFY
kQHPFngLIHqQTc0B2d8YHBBSe1GuICqhSz58QRpXgJqam9xg6bFv6wcSCVPWWyvGGidsEjebsRe4
6/uY+G1gb9gUbIKngVkCgQLW8Lnt8vE95Y6fqJkpSAWruaUsAzg3xF4vkn1G+11ZiEScaFpCcMOu
rXRvFMBJyHup8HlMLN5USXtd+FVLKvGNVnSo2PGFfphTyre0zgQAsDEFh00HachT8IVKz6qPDhW9
KvPJT9XRJ/7wUHc/775RiHmZgPVZGJZchfdqPYznDzTjcJnGb8unw8V+ThUppKGi4ivVT2pc+wL+
SWdENzjSO4/LJ/968G5RWrxwcVhsoE38zmX8Z/swDViE85nse/A2mEelYW+LjGJauPWZ/vCTm06P
Xoo/Y6aWuYqemRGjyxub4a6QP9HwcL6avEmq4V9F6f0Ul4eBnzYCoaUCjduf/5rNDmmsnwdy8WNt
evvvAPyMHpb5va7OybiDYjW13Od1GsBXhCsVZ1DoKV/Zrh2yTi1EihNqJtpMQB3q1cdHaP8/7HVM
TpBSwqhxSUCpcf0Cg6WVNi2y07t47xJijd7JrBNxd9wi2do8hfwtRf15GrmoyvijtYns859qFmBa
RbZiAKOvMXout06Ni8ybU3f7iVJj9GbVb8eCkI0smUU7K2veMxMW5Q28oK2bYECl19Umg08Tw6R6
B4bXFefUAol2gGD05483vJ35uRQiNwGTYgMMY170uzNEsO1FVPHvuQY3mfGXn2aXMzd9VeXNUU8z
tU6tJrkj+5rssxEL3DfufXiWS5g5V6ceP6lQoyg/qpTVM+9h5uWIkzz7MTvC5H5nGv7JQQ2buLIF
Jg6XYcydnL0wlnocU5soxNmw0vqhQkvB+lX/3SC1ejLbgDX4QoHABWAhMEaLah5JAkCxUf8JYUlW
8MHxvNEJYhZqZnKh8UVJijlZbj1tQ7yZ8hkkv5BXgnF+N/nwOR9Q8PKBhE3WHAUrhMMJ4FiqVYTp
Q3SpNqkziugWBrlL2iEPeIOhFvVw8CD9yDbjF1ddGroCURB577EAqVZrn3Es4Ij6iRmupVnogZpA
WHMX0DMoGktmaJSzBJJk5rjvBhXiI5TUpnhGE/VAfFTlcbfSiUC0yuPpgPaKyt/6l1y45dEh5ldi
EqhssCCraRKgC4CPiydn5Nk1rOBjisF9Kil2Y1Uy8Ye9YTGol4CGmmilzBif4JawEcETK6VPdCiX
VuQf0HUEV8gKndet1GanN8KEq9Ex8QAg/xcaGL2fmBn9yJeSo4M15y/pInnd8FBXDUVcDRIPOEbg
3n8QmGqZ42hlgvJOUlX1P7K1NBcZ/Wq3XAxjvrQsZh5/Ik1gCxuiWIe90et/OaELUIYFSTH0wdDK
av6mZf1JCdMefty0+mvLlMV+OVkWwlCoBxe/CMs6AB3ENDrvZgjKGWccoe7zmTR1/0u9U9F3mU0l
6lZL/9LeoVP+vien6+Wt3hLR23zzSG/etz6gd3uwEfSeKiNg4a/xZT6zjUIbaoiB9fnQKAgxO2Dn
l336RNYEdybhXrGl5hzlriELAD9aHO3eNmvHuHHtLvRvd58IfWlh4M27YBFeBRGiTTOm3FA3PEKW
RliT1vZThKh6gdpziqfOuo69jelhYvAwmXe+/ey/bUTbCvGoKXa0mK7PR94ply4FNbo0XNJDHAhX
Q27M4+dj2EOibevXO5cWBPHwVEMCZPFoYSxYbJxzEryfgjjlqfQD4ERp1bmGbX5k8kJKezY/GWfT
MJcDTGWDlRcnSQHIo7Iw6iHMxAEBlBK8QeIh8o8EMNuLzpCPx0JuJHikBOx9iuFKa4qs3GRtbRww
u3W5cO7C0jIUeEgI5OLQIVXnvdL3rz0BoP0kc+fZXlRE3eymFvb5rAR1myOW+idvs2RKjikTgMFA
UFhz/WtYCufSryTPpw9fQcK4Rahjihe3elOdePt9WkcEA5ooChkvbkj72fnAl8VoPxjx+MuIJMjJ
7eq9GlWXZsw5StWkKQSrm2jTOK9aHZNVvSalY7zZieEYvOPMgWytT3sF/tMgjC/mhOkfVBEJn+sv
TlbDFobhk53AYFxAeew27qyw0SZeBZ3bDZD7hoOCIUULf8NRm5BBfdYJ0IXcHxmFauHLKkpv3x3Q
Y0LhxBd/vEwY2SWD4Kw+xIY/n20bRQ/eXVWyGX2o52Zm2u8RnoSj4EG8uRAvHZv1/STirXjl9Epf
dUnpJygQnEBVYsId5ZLWrdOq4YQCDbRvf9PUfEiQY2RmFA8TImhzHLTF9r8zGOCyDiunaYTz2wHL
qYoOxKc5la4GEO6zr86zfEq/UQAB07QIZZMlV5Z81BGtnwOffscbynYB/Tv+Tt66W3cDeehfGZb/
3XtU5aApHZ+ae0UB40aNhfd5KcgsWT82C5AeKn/l4bcppz9lIMoKF9l56+DUKsUQurXy51T0+CTK
znddAXLTILnFrIZJtOjHQzm0vOshf0DFJt6hNaYJcx1mYi+ztQKa7ocmX7XnAXj2sgMP8gWERMWJ
oc0XpNSTKGuAhFaCOc7/M+R6BHVuEvgVzn2c9t/AJoi1wiJtN79AkCigBYXd2540FhC5vLI3wQCF
CSyrNCx0qtdQLMJsDGrVjJo/o3kTpBzJyc3M4tneRo2fcHrdIzqReiQJ0oa1ldAfTMnW5EztJihG
nOnXyX1txDvr7zYWBvNZ1l5KMJI+ZAObdPOV/zQLE27yuqlk+73ac48wQXYIkpJEjlIri4gsl3aY
tgSijY3qDsJwH6Dlbw+fEbPNpvauhwSlfxspwWyY5l4tPvDrqohPhovXebDMF/TEKbgpm2ULwWw7
9O4fzoK6sIekHsI5wGiNYZHLc1QTo45OgMKGU9DxVCYNs0mzx6+ovG//ApQzNF2t2sIcbcIW7Nnu
y9hxOsJo1EhYL0NuJzodcDNcCKg3vapwzH9VIY7jwzTmifgh13GgKleaiW6Jwyw4Bjn4jn8X6ge3
xVM9LpL7pKbNH/YyGb2wQylCuCHcm0V3I+RKH+S/5jDalUbIUKtkph1s+uZYTyfyBgfOiep1hAoJ
Q4QoVdtn9pZMpjdQX3CTMmYrixvGlFYAQDxH6j6oNIAI+ZAq9Ksvr3okvZ9CM60BQAcZSrcuzGXN
IDaSXl+AXaKdj9pc2j94pEv07ErVneiesNvwevNDBqUQbHglSVC3BEbrV5trMUQBss/CRpQIHc3q
UKkB41bWo6cly91w8A4MTkvGmu0fP3pzN466JyjDB/y0om2WOdN93OuiKVZfEpqCKSYhJJl63OUi
h39877EHqhozvZPKrGHWZ03hzjrhM8MoAwrPn0e+ShlNbWO0+anxEvs2pfpADmYpWVhhrLEAVnZC
EQi/2Vviti35YBRu4Bnl5wXpAZeq0QYB4nyGacc2NkcrTc7bGYLOSMUt5cDIF53reo29igrt1nPH
Zeg9T8sHdijo18Us77lDUjjS0FHKeNjEOJy81jwoqHJxlYe84swH/wTE8arRk/OUfo/BhDNbFTTk
sqse1yYOikyO6XIXLBF0G+ejbjHSNbbqKyQw28H3dcSKfk9PHJyrWJWdxD6A6XcIICbUuZ76jwum
6sUBOzDuUMF0j3S2HFxrjKDpfDZCZAfd1qhaKkglxplGNIHA/G7MDnoWiytDia3ML30106iSdfRk
uRvhEhuLYn6TzQYmbZ2LeHl/4lvAbq8Uj6uLKnsI707yk1QnPMhV+MEzro+TYb6yBufMCPLFNsV1
Jw+b18D88waJKGmT08NyW11Ar6lKGIkJtFKLqQ90iCxySA0ubB8jMPkDpaI7ZryxssiH4VDDzeee
MSFtV18DTy2xaumzAH/QXbaeKifSID78pmE18mBdVdfYVtDXr+ymnfhzfqVAljLweXahmPJNFkzN
OSmDU6+zaBVA0WusZA5jZlMkWCJjnP/viJ0otrHn2fBdRYQXnZR6NlyMc9uyUnM9ilgYz5OQgkl1
BDyAFq7hY/tFh8Dbpc67FhZmXny6Ke3j2A5xc6/I3Whray1ln/Rf6sBAZaBJ5PZGo/fYlyhapTew
oguAHlPo6YEJ8mQysJL8gAPXDvU1egwHCC+YhN24fR5jO0MUtYJfv8lGMZuXQLDXvN59CQOI2vKz
Rm82zvzwC+I2pA4e18AO3JbsEdNN2x8iVgPhhcQ0Tx0vS5kzzQai6pTtGpDYLMf12M6hfebpnpv9
nvTFGYvwUK+yg6x0xF0pGOixKWeI2Yr89UXpsO5Btdw78E+VysPWRauTcwm8V4ENpjAaV3cRk4zS
D35a6cPAlmRETezNYrWDB51emeZKnqxHIn2XQN1a+DZi/4AmIRm1s7Fvmnho2mjAJSy4/Zurxl5L
NbrebsMgtktaFoq6ZcxUviAekVDMlSQV2SGnlGznz0/PzAYksVlnQEm2csmQGZ1eJCqn/d+N77ak
qbkCt57fHclJ01Oq97Rxgs5ETktmskYcpCjwk8QcmOK155HYaviYH6Hvmp6sXZvaSrFZuYzaEx5p
Y9xTWNwt1YikRRTlLnfMNbhxXYaoWUd/xTgPaUHx9AcqapFtqLA2VzTrZRGRszJrYFvFHJVkj+B4
PtimZNe4b5AKLeDhrf0tCCW/1a8x97uFC4vqQzyVLw46mHXnEznZ/k4KYINMmzCBSRr3MrFZBBfS
ftlBpa+yBR1+9uh2V7+0DygA2UKp047St4iozzQ4QwxkGj0UiOVxIZ/cSKJD9FzC1hBsBVZ0cOwo
5I9umjrF9bvBd92qLgHPeuAaGxEkKrhJ87OovgpQajx2hsZ+I6lF+8bwaK8bekf8Um035D5og+YV
0CHbh2/uYyFG69DI7hd0+mFBEm/P9NK3mx5PMyWxaq7nZlSIqMQVUM+V6zq34JJ0Mx9FysiOecn4
ZLQXfOVrnJSdHb0JkI23Nr3fS5rlITZJRl5oKrzd2YgJjHgCXGIFG+UBygzuOsXld4rb82shLBlV
OykLQ6yl4M1npNDwqVSVqQspOzQJ1B5/A9UcZMq4weLESGav/BzrsAr6mhQtbVW114prLn3mt7i7
amzkE0kMTho6z+MHkXTDWeN1S7l6TiecS9SjnssSs6MlJ6Le51yR5/wLD9kAgBRh9FtDgLX/4mof
Z4QOEMxy1qEs8sBARza6m7wY7/ou1dnOPIK0zrVNdu739G0hmG7exNikfPr5K69NkPhZ/XbjHUbU
zTeYMlcZ6bLrz3JrCwoZfk339l1vcQpRBJ8lkpiHpwWVZhRNNVEU0W95xpG+zWO3RcagUYNvWVI2
dmIHYDUGuue8kt3Ggg1sKaPNeCHggniJJCFZhTazdx33/Ktu9fKexOB2CpYPXO8P+mO/uNFJLuv1
sGhJk32sJEjHPr7pXHaeW8USOmMwT+F9q+FQEtp/ijnWAl6G7dFU/rFYCICG0hXrylgdGso2IrC7
w0ekURFWBW88YPlOT2NpFKLukfJuz+NSlkeSYWZyGY1BB2vX/m+WEPzU1XHHqNWaDY1cWtRNuw/E
kOGQ0HupjINWXV3EPfRpBxN8JS6dUZL2804rPK0mmtQFq9Bwv9THSWnkNRSuZtGPxsTbNaemSqD4
vy+oCDKnfhAE5RiZIWlKPqrQi92txRFw5xn33YYiGITPsC/oXRZKJhJq/gMmUm1RM9R3hqz//DRs
Ul+qPQCnLFiocnRA9OahG8W+qYBgTqOFROriiqiAvaIWTnWn6+m57wuaGn+4rdZgSbA8+X5xNLuW
InvBhR78ZkD51GXt6Y3X/qx19Xbor2/D3eKL/suWYwkffhvaSlbFNo4/+nUSNSnOgnY/N1rVjwvr
BAjI+rr+10+gZ8CRyQYWYClNSHNuhluFn4ctjwXhM8k694Sd3qS5/5l0LgJwB8/FUYp+7HoY91lw
cdv23pNjSAaB+/fS00D76Ydmryr6Kl3J8342ebxdnw05+mFSr9ut61HuFVto0AIPKbcUt3h/jm25
POGVfxojUdc5jLwhOIj/s1bi/I0Qh3HFO3FnVfpF2Nu69kQ21ze4aWLLPzfiT2KWT4yBrLkK+J1M
xyJn7QGE7Ru2rYApU6VF2d8gwE/fMrGyeukW+YA08SQoDO9X8FFrUgMzlr+jDarIlZ+C0SOCXN+3
SGYeNCfheHe5VmalyLSZsspK01fNb22bVoYy9GEfvBrvXyakEFZbE/9prKpSq3SVF69GPSg9Y5G2
qJY4sE7Wt9LrMION70pX3CugNRUTjVCsjuI2LIdmfDI2DlUWQAnnbTO9tySykc3CeOuuDN3agjdh
BGr4ovNPVq/1tBPDgWX6kXs+N/hNvErpuLeV6ILDNeuvzZ2EGtBuclV6K+ELBlPrN4Xk9pX1D0X0
ma1Wo/eOFUK1rqMA7nAsDOfBYmHylW4zvu7EDpZ5OnzA6zldmpNArcZ4Pl18/JSOkLeSjYcDNutb
6/lEt+yHT/oVD7g9K4K3snHNE+ZdEdiD/smeyshlVfuY7Lz5CZ7RQknS4CpVLhWzBP8vz7kpP0K4
FHAGpyjMLipkOtglMd34XNC8LcrMuyWXgo91a8uvAlef9ui49QpxIHUGDG5ZJVhs2D0ccoYls5BQ
BYrnb1quTGc2cMYbxA7oJLOYB24g990eJsxvVuA+q1oVix/sEMKhNo1PbNS4nyvWonLHi5BgNWL9
tKDlLn+uXWn0h8arXQK/VNyXS0X7ZrCzQzvKGKQMwpbF4b3dlh9BwhiGtB/MehZmq/gKc4rhMQ7L
qHhtw0DbQA0hnqNNzerXcLg63mbb4tMusfK9chP9AuE+d3t4s1SpD4cLRSAfNLISsa88JSD954O/
4PrIwDSBc03Y3CiIWNRSbswBmmGy8BNm3kZWROyZu0wmW1f378E3NItGsuHpdELsazJMHThdoHDu
JcO52Dghye/P3dJfAC4u+yVqfOSMgDiWTqcs1AEMwCtxf64pf+Il6Y0JifeKSql5qGTjXNgK/4mr
Ja0OWN6t0cCE0TAV5Abm+nr3n9ZA0nNb/TjUiAhs4ars5KU8jRVBv52ALLDDjO79iamcnpgTAO9/
llvGaUnExwN75gkFMVhRikGx2QFqznePZVxARhg12WlYVZ1a2qfbCVfbBqVCO624x50cwrVAVG4c
pjwPiOC1bstgaW3fYXE4FxavAOKgIXZlqol3rqPaXJK6JRYGAGhTemqoKADvwheVyo2LSusB589i
+EtLpjsPypol1yyW6m3eXegzhLdKu3O9xKw+eut4c1BW6OgUhOxjIzmDZpO/1QJM53DnsIu3QEtU
IDX6h5eY4GFG/khX4NBEuoJ7CcHX03FV0daEpBQfYCJjJMMuZseyTJBwNJGz1zKGT+47tiS0Gs2Y
9BM9h16uRDzt0Z299s03Kl9qpxqr2e5EB6dR5aAUdFVxboYuM9jiZnSO+tX9MLpGaUrDY3UHgvpv
o1n9hsQZRvzkR5yoahvW/lJFQp9CIH9BViiUyRvqIiLOIr+Jz4jInxWaDItSQaUN06QSLltD+QIF
F9UYGLBpGjmtc+IsGPnswbrwq3SZGH8GKtISDXRGLMJWd/YQMdN14JfVMl/DKpJIn5CZg3Fcc2yg
RCO1iDBXGeqzilFGn3uNSwVC3WhZNDW6zxZmWwYDy0TlD8JTU0kKqgu1gRPCcCUXdarHokVUAapt
3GKi3XpBlS9zTDR3Tudj7oYyjAAJBFC2hUng2hOyQnpxp1sSfy6dM6sHySA5pbq/sTz7Wh4yj6WP
dFQTWXF197/kJ3eo46s0mD51NpuPguVlDP9oKYEMbFWgCb0yVShhPueQ4Az1Qd70zjmbjNm04adc
1YGz5Yqw7TVPo4Jip7H8Hu7qJuJWTodcIpuUevgJAwF8fozjxel780KuDkjQxM9g9M1lxiDtPx46
BgKvcbTKJtgp+UMB2kydYoPIt/RwoG1BypLXRJmstNDhJ7ZYtmzCgBFUZ1qPcC4Ouvj5C3sqnCNv
CkO1ScHK0dAYEYNSRYGZFwzGn7CfI2bQW9oub1MMJVjBmVCVJIEsAY6+si1ipyR2wi1nyrYFk5kn
Htp9CroKRBgyIj7k3AGR3P1u9Kc0Qe+j3qupjE2Rzcn+PcVdNtKiLiSNTyQnjXxOQxN3UYHJPAaC
iASaeVjaVHvsJXT0I+Jp431JP1BwVCYF7vD19lTRtCfIDAFtH0BTHx7wPBrGrWlFPKW7waUU0seK
1qI40NGWX1dDlZe0nkGwFmNOWLUe5mOse/jcAS3P016Z0NaTHKrdxge7TrYK7qVW1FsEh8AmooOb
TlJDkBx6gQ3OUAZTtzmRXT+s1B/JHcHOf70EN9HJzQ7rBmLUll+ZinQzP2M+TzkFHI8gqL6x+rnz
atHuue5+PI8MAS3qRWIJ7CZ8IY+inLdVLw9KGLuyrzFgxIKPTCVzYFCebxwk2oyXOoYjc+jHH9yI
56atAGKecQ94iesEe+kjv/lbzqgWua0nszlK/YZNZi84X0cgvK4S/w2TzPWHh5QqueZNRedr9qLP
29ATDPHMIwzD1xQKVAvsil0Us41lyxbb0UZ/A1M9FIPkfeNHAeDR6UGVwQtm7E4d8+tFFm/QzgPD
5dqAYeEPsZu/ObQIe9qD+fNj4v20ittsU5sHglfmHXUpU9lza9DtW+s8iffuNfG0Kxo3eQAWongM
tVpyWn8F57Yx16b2hc/8cgHdmNyY6xAUYd5qqaGkdv8EJlJv0+r4m8VmW8NEJn63Z3ydR1yGvx7K
2x4aEK3K/eFODOmlYgzzyN1aTo6sPVUd1M9Kw1svED7iKp/r4ij6gHjJimK40NVAEjNNPziYvX7E
POhPRnNg5Xt7tCbGkkn+jBCyVkDN0OKPl6DaQxFny044pcilwCQZhdH67F8o1U2oYygPWmLQicS5
0le9rEIHNWDGSSWsWIhud2ZrSwoOCfZyAUulHnez9RSA//cD5DpZjA8qJVo6AF2zP1xsKtVHqRvW
ck2m2gX8TSDTlx2BJH8z4Wk8SrGJWxDAeJeqVOXON2PuEBTkZDAs0ipAqUlUZVHnEhJXkrK6n7MI
FHYv7b7YyMg8PYpbRD9QyT0Dj4LQRxVvZLEJNu4rRhp4cn1y11WeQjBnMkCIXglH7OabKnAJVnTX
W3/t7qBhkojcRilZibBipojNGFhNFsGsICEqnYfbzFOBZBj09g/WiITzmhb6+ZVYXvEmcaZ33qNi
c20JRxGOgglw2/7hLK1jyNiPGKrYgZ6wZLdm2YF4pD5xorTnoaYhkcwAYSJEHKJkEGn1SbdnlI4g
ZS4C9a7RcOSiE4/Pf9LczY6aNjCer7XAMmbNJeCKLnPiBFpk05RjVGtg0oXgztmRAjIu11tq7ejf
stnXsY0XUUq8i/anJ4jlvsarsElDgEpxZwpf46WX/WHK28/Je7zw7NxExGJ6i57h02yiaXPcMrsA
n2SDE114M8I0F5tr7/PRXDclS13N6DUcttdmn2gpbnfKXmBNI7BWSTxER1HYhmjRABi2QLUKApl7
HK58ML7YPluTVKl7lJ0kDy80jopuk0bJz9aBxTPzkegebMGI3cLjS+Ju5/txMyJpHKMAiVQEUWfs
8lMUZKYDY5AcJ5Pn8zp29cow8ZJggs0LHViwjWXPrd+QvzBj67h/ee0ukNhxB9lBlZBjxEFO2XKH
1OhtHNEMOC/6FABw8YVDjD5S+6b3Pw70rZSv/ci3h2umhXSKuB3XRbBGcR7OEexeTOCj+jQw8Fkd
ULa8JZ4aq4X+m/qnn3Uzl2X8IXr4pMeJIhXsF5/eAuYt4hpOspIdJFIFyPbCcsB2eIJjgsIwEaes
y5YVezT3ok0UAGZ71dCL0Bk5isTp848Y0H/Vs8pOSQ4Dhx58IpKfBy12AmIL+MCfxixl1wEGqPx8
vhI32l4D1vlrZtdb0HrJDQegDvJs5IHhhxQwSQW7p9ZOWPWvl/TuzRZIM2792iKManqYF4hUh6EA
rjviDtxva2Y9q3zYs9xNtaeseVI95FLadRMN23bkrIzP9n604aAZEyJm8J/coyYSVwxWrIaOjHpj
fsFZBBlDGvNsK3rwYEdXINhuEhlmnNd3A1Yk9p2mFsJLiqtEUbmBgZyWQdKY4tSkDFZRHqPMC09d
s1Vpjo0O8L3oKkaU+hZke6jG71rm+87MdfqTcmguDBKhBWuC5qWX8MBlQNhesdbCx92DQwY1SneH
yqbRMFPwgHHg2ASGzekDshBgDTnh66pf1EBUM/D9eO6ukLObOX0hCO+65v05t6AExImO184+M/w/
Aaw3XcHhROwFl+dGSHTLn6q7ihkA/U5hPCkh9Ay/aGvubdNwSiEMt9HJDPZScgoHzBWEvLeHWfK8
7XnqmbLHsc5A7HBfzVWxRDFIfLvUcwo7RPUSIYwOxk6XnIhHv87n0v4pxNV2JO7Hgdm/LhIFHax7
OdG9vKLqP/0wWFGTPnNd0FlJg+dKAo4tq/VBfmFbXUD2GmayiIaWNKm/RSfFQQ5RC8pIXB/Y90X4
oFdJn9SflVIADPxfd2lOhpPgGQByd9yWGTAWPR5MTd8vjcXCfRfltEF3i9cvpy4c6PgEgqqO10Tm
quzKM80MlalQo3munM3xbsUtoplyRmpD4+VWpb4hwzgNRu15cpR5UDg3gmFQMnDVjW2zRbGv+PR2
Ti15K/jh1AqYMViagCEXzz+rwIFgOGlEnX1wh88ehyIyTYnRGgppa4trARGO/zzN/iq1RYgXFBwX
Fg7mxwBsobgA9SSx4qtZC6ND5axKpFBGV6VsElmjjM07+5mJ2qBavqbbI3Fa5OhvPmY7UdBRMFyZ
RTh/HC//7rmr6PPvtZnYEVG4VRYVrFPjLhKniaoBj75/wyWl82y6v+PuMGYyLsSaKjePPXqU9t3c
IWyIlddy24gvetwJCglMrf1frMjR1qkdb6wW2IIWfVAggXJAuYgqPxeWDJDMAzLC80g1QxzuTjNW
37AEGe9o6yc/0ovBhx8kFm86xQFA0PuldT/RifvpJcN5XnB/lgvC9uXy3iDsqJfgYqjQ7rES/dw6
g1p6NwucUkm1IMF0v5iQt3z/9RbrrtunfRZYZTaYI1dnPzyrN1dyZk2EoGVcOvYYtb7F47KJ6VOy
r9XtbkPh1lEcBcXibV7y2Zfy+vXRFiCb38qrVdUhUEtpHBSLsqV8ItTyhV5URJKWrgZ8fVWKSHs2
flRaotMzy7b63ejJb9mAACCEOhp5VcwY2bduuyQWN+XTDkNAA8bQRTC5bWe+vI966gr1mg9Mm/Th
9orEjdDGwUUx0kPxrjFcQCqPuRUmxKyB0S9zyb4IHuPtEYczcLRmwj6+KN5TTyrjRuP13Je3iWuA
0mN2zbYLB8alaAvM5JGlzRQbv5LGhsUgPD8JHF8pZGKJ8mutltqy9MoUl+YufAO9IcUwP5s0xpzB
3bxAuK6bat/sq2HL6k4X/7ecsXHrtgVWOvqcE79te1KUey+1uOKxnGXMNIKbKitHJs5Ybs8Nfrrg
fLMp4NkUrQqpugoTnFV1FE5399XypR5vTZ2eo49+LClTkb03zIM7KR27c/Du7H/oIJhBH8xqk/jr
QFOzozoakoGLk6ZGswVuqwdY9/jxQGNKNr1Kf1s6vuV0Mag806b5DGwfNgFj767pPiez3iHnyzbx
fqhHcY4QAzBD7949omkEh8fhHqfbTDiYqM8BYVFGkUrBkN7c8ytlv3Q0NikWo/ch63S6Mc+FD3mz
ZRgOs3eylOz2W3q9FMbfDUwL71XINhjQ1oLg6YtwCmmh4HxiqcOMDvMnpB8IT5SCG9Yz3Slx6Jj9
XUE6vtGKoi3YjKpsOpIQj7kvB4iUM6nPWg4saBgQgqCUsbXOTThHuyfeurqqTRktjzXblBXcENsg
pyRtTC9GsFgjkJUTJTeabfAEg46l8d3MIR9delQnv1HZBZ9BtWsEArfgY7Ovlzlc5kk7zuESH0Sd
lheGHbgve7QXQQ1DrLd/FzkqbUgJSdUqlfkBtS9azpsfr7G3RU9AZ/FXDzKe1NUDuXTDW0j/7wZh
95uikjGyQZNezl+hgk9bw4BYzn0pMEVM+JsghTPv8FBcrfuveeM7CTEBkEfSQ2EUgHsIInQatb05
Pm1PujlZ/HdIxetOz9Fq5ulW9OuBvCl8q3Pn02xcA9BA6cPs2KSoLl5JyWKc8JW9scBs3e+BJqMU
uZoZGf0c4w2cY9RahcVJcACt5vvfC1ErfcuTnmu5vsUYIotshVZbC8IgO/+jOENmFNLPbHeS6Fqi
Js4XgQHzvj0oJ8uDa/D5330gIpgQRwu7R7PE6dR160dIF+i2FDsNrZnXqMvXeEfh7PnfuIriKxAy
7CPZAHxCLBpLslrw7MmtBfTEZqIatocgkVLMBV6kZa2Dd5QE3WaI30xCG4Ycf4KC5vc0MZ/PxIu4
MXxGwlLf51DvHpMmL4hYKngr8wLThu+9vzKybAyqoxUGBKgXFc/ebAirK6QaBLtzya908qdA8K/2
oMb9iQI6TDqLa+hL4tIh+Yb4mJQdOlL1LVaT5425dkN1w0Tb0ksTrwY9B25Q/cvcgbEGb+rwKk4K
HMbXJoeiBml7o+CV3XldFf1WqJykAxWhuokZ0fzlRJ3ZmTOCGTIGQMMPA6wzlVPbUAM2ohyE7svT
0WUbAPS4/TARLpWxf4t45dUQ5WlspktrO3JqVchbdrK5bdC8abhTNS+MFKjPYPWF21NMXTkcRu0d
qXeRGhw/DcBDfccYWoIihVpugQ7DrdMiDbP+cKx73ThhuanHtqxMXakwDTPQROjAlkiO5WJ8eIfl
ieQhYKDzmrHJ83aP0UaLeFFV75fiN6U98uSQ/a7ts3OzReBN3isuyESHx8JLpPeN3rnbIWugZqAu
yb70bCM3zCNQKvJ3tQ5l3AGI1GnxlZLLtQnDWGYPt1OI8WRngNavMh7orVNz4Gj4oNK54M1mbR0k
42OpPeIlSrYBwPI5qmnaIXBXI+R7l6Rwc9roXiNGaQm+mGUyi45xP0ZxOHAJZBqd8ni4rwnKkBGU
pAOs511YmAh6DBaJE5CH8SYw85dmwh1WhZDu34TT9mjPzUMvrC2eUxDoxMDeFlbxj7mwvrhxX/O9
OIFHO1/qaG99afMyQSkVE0vtyizOKT6Cmu5e6L6unD49yRu7tLsxBO0inbGyL98QcP3vOCJ3cmED
TaIHvcPVKCeaT6/0XL0ndqEMjuJK3+2XhGdPGRwO5812lxFwUoosU2f6ycuvcYY1NwiGJYxocwUH
AVt63Td1J38EehVc1ZSlX6mBlbP0EdQG6vPJHT8eSVh7mnu4rY1uGBVWhqVTT+LVB8SMISgQvYch
EGFjPYzqFmX9Qpk7gjYOdCnTod/mtPOhiFjn5ubuHAB0TKS2QGY7oJt0oiQI/YMZnGc8KLZgDSSV
q/+EWYlUToyLpQhaQW98w2BymkV/L+Wz9KwZYayErHhPeTxssejUbNe5vPlIAdfwEYVwnn0fo871
V3UlCDUwzEtkCkhhwmfdbMJEVlgPhfCNH6rsHHKC6IuCDujTHx9iXYjeVrJXAePINuYrk9DJTjUU
4yyVLsehpKwB9ATSFAi0fHig7gGU2XSspYmbaggrsEc1CJtkCI+/0Ud62NkMADOiLzXcTZb//gXa
GF/EQazJk/uwAY6FMNBd7o6qtTN3cXLE1sOHdKOHimUf0OY9ZqmvjgrIOIVsBe8Jn3W7gkNQTL4t
L43yzo2LDiXdzzAJvgLdahlTfvAzODUIyY+N8sez0OukSn7tXnEv5NtBia7eMSL5Ryzbt3C7RmW0
RgfKW+UwMvHy7ThgjBxIWs4cyg44A2yNivngzt7hVvrnOmPR2TCHdpiTR6tKwTvQvV44KasvU0LV
EdypVz+lkPao+7B9jEfOqp5jzn2g3kJY//sDzJ0iXvKL683EZtviHZWk4Ax4JmSIe5wU9bhKxmzo
0iOKI+i1PIm2BeZzqnekeLTM91FxvAEf+snpzXQjzWvon+MGgo4uXWHVuobsjW/CyGMB1ODHreVk
nH4ngMAXdDGDQ/uSFSOgxCOVMo86uqQuI4yOYlgfXUnRmO+zRn9wQZukmXbIJmzLDqW2Ss6Aez8v
mX7FCho3uDjxwr9xxSwTN7rDFD6XMTdlwxqSuQD6y4DT3LW+/rc5mWsFhGeTNQKPRkuD7RnGDn2E
/ictx6uceSxAfXEbYPGyk/9HrWHU855z6jdPFDkRICNRLoZsSFTDaZv/tVFBK4XzJ57zeYjVTn0B
ISx57aJ7fRydC9Cn+zDl2wQUt3aevDYBO8J2+zNkp1JacQ18YmarObMgu6INRkqoskB8JryFw5Y/
n4yJay6LyJcLv46TGOlqCF6M1y4Rjcwz9YbQ/UUuzfXJxfQg72xrJUnZCuyvoRPZmr/3KT4BS28p
QQSSar7Utlt7IOLWxfHr1vFFQtuF3iwFV+LnsLio8Tlhk0Cga9aHfBZVVKu1ZDaThcWUzJRQfCrh
H/2vj05QqDMkWlC4TCwpjD5bu8fztP2MSPzOQXxMpfNd3bRGmPZMocuPGMnIOMiKNyAWvAJd9fKo
+B+yd9jwwyU/yRiqkVEv3hI2J272KF37b/+9V7t6LfDIglpD3GYwKKC8SOGFbg1/2ZRN6U/UzJ7r
8XYa2eGWFupKr0dTcfQzBOccwpD59KT6ZX1C7Ngx59WVd2qF1qf5IZuAkaHun3RgSTQwdSWFdpOp
tbNglbZMjSs8GCVyyILGqSrz39hmLDEMN7E8eBpEiTyQfZS+3bRqKx6Cb4gNoWBBrQQvpBRvXEqU
JGlKLMxlPl4meuFv18tdRWkm3RWKB0m/DpXgtjccWM7p3VrvLRvwM4/sTOP43WaraLn480bHGuLR
xUTkYaG6A6SjipD3dlGuurWZhJ5lQrrXFbnoKN6E+6hahHmwz7KCKzrPFBTft+KRtOfQysQUWKKU
Br093+6s/sWwxy+eICwKNsZi6CfW7VuKFucE/YLuz0dORHAyJPSBLZnWyftxp5eoZhqTC54A9QNa
kaM+HluyOGyhp+zYsNGnVnLPAmRgtYgaI688/anweC9ctmDgdcjTiFsmYNsroJozDGRJSrSczECI
PGfXZoHxxur8fOfgnMe8U//kMB0HMztCm/dXvTy21o2jst6AKAsybo6S9wP3YkChW5yW5FvJwDMf
INnCxcNGjSK5kSXJ9RPPkaCO1xi3Axo1dFVMi9xuCXbco+B96Zi7rojwIPJrk3suu/wBveWLn8JQ
sr6FYVKAtGzzWml10s7BITWOT7KmwI/JXT1eqrolfc9u9OGGlQG30ZMgJQjWn1f71llEi39j6dKB
mDbF9q9S8XGcYJcwd8SSbZWol3vsJwUh2vs1ONUbNcCW5UgeL7rATyfUESjkd8u6Wl6Y/sa5Kueh
6rUU2a363SUP47/Dz9Xni70joZnbT9vvsJ2KRrqAx5Yx0QPkSQaPdLjjYYBTv01SOBGPQEDI9N3N
+QY6uSGLNW2pJ9seZ+kPGDwCzlCp7FYj8ySwb90XhDuBnDvH+uG3o8ByTjRJz+vtnZ8G/KCQCP0h
AuOmAQ0V1o8hV1UoQvKSIXulQ+BR0ejDWLzQXg5FMXpehNejAZ2HTgmSITGsLO/5uqPlgTgM6IRD
QaGgGCd7V9kG38ge2vsXwDjhttYb+h0y063HZDGgO63KpmjkKbeSpTj1AXt0HdMVqmf/cqO00+aL
VC82gotxJR/8QdeFtX/s6FDsVcGQ9/SdxcNtbzSNsh/3INrgoBMIqi8+gQntiS2aPsQq1RVv2peY
24rooHSlgkSv6LjVoTmxNATxe1vf6ElX7L9eeb44+WL+RuPs3Hh4BKazLZgIowL7MqQ8IuC+tz1Q
Ne1XE2mvRlgiAIePu6QjHwiqrCKIcxfUqrJ1VMS3ngxlsqeo87hRK9ND9pQCmvZdSkvIWn+PkpCY
rNilz1DfMlBjKfSK01lHBsX4jYuoZbhKFHTAhg83jGg1bvyzGhlsXSZtFdYqw6RlJuVZ69dESKCs
u1rwzb+gLwA+rFCc4SWphwO8SxAXiyGHFqBJRtTN5e/O3AvdtEsBgOuKh8+oaX0rsBvUTeI8+Wof
jURXyy1zsqq42ZSZgIcEwOCyPd1odTX5fGFT5/lvHAdS1oVwNy6XPYZU9eW0fwmBxnCqnBeDIIWA
gD28iagcjwr8/YcG9q3XIKCe0FGwdNY0GZesqsJRiIBACnQSCjCJZZpYrSE/eIdxmwPfPlNopA6Y
PaNSEwQ5128B3Bi7nk4kZiOHEGgnHnrMM7dYiIAXR5AS38EXYSmjNQPmeAhBn1WSaclF8I5h3HlD
g03rQvvu4PjAWxNAfCNd0xmtpGFCZXcO4mrVyUaepQDt56Kh+BDeZL8ZdX/o3qNBiq+F3kRfwVJU
NxrGddbcrdQ3Q1uMaRnIKalDeNCTJibGfmHL64WmsNVe+D8O0RbgNK1JunX1d5BBt5+y/UEdyp9w
DX4j1FMKGaXQol+XDDDwBkSVnka05WWt7DrhMgQGQO0jFOZZobUm9TqvFf+4qRKdeYX487PsY4O+
jaXa43EU/ehXHIlRw1feEJdIFg5NyqlLykqChn6wzP8JuyQTH3GARFYogLooBr+jCchOuW7QAv43
GPp/mpnReWlZ8P6Qcpj7yOSgOb/Sm1l3tAkbZ/l59/ASA2GtVBB2A9li5SBE86tnfMYCpHWCydH9
sWY3DMCyE3uzZv3w8Prqj40JrUosEEwUqWGB6XeYfQXDDDf1bB0t+BRvM3GDc9gGyOp9AntdDgbV
m8DgkpmPO1e2PPaEgRWB6gCczAeAVkposMVIWbcMxoJvyHnn56KnCWskobrKxqzb/YR5AAClP3aI
bc6f+E4hoK6+K5GMCAsoub7oEFaCY0HpZnq/dhxKki0xQa5RoxBUNL3rLqLKYy8UYNx9MqA6wXCd
lXctHoKjEkBd2F4iEvGZsjq0fHmDoV5N4CfkcPxe8ybc2oBoTYYMhN9O3cUGJQNpz+fAV9x5l1WC
Jz3FDwGPwYyowGQ2o7/qnRAGy+0+tQBuc73oXIndh/zK3Fn4a+lBJIxoC6eSJFaUA91yDYVmgMUb
dgv45ooeo3tr75YjC/q8r7POizDZRv7nBQP05NaA9AcUEGzvIDph/bvnfBymS5AHBl7RbW6ph1VV
Xp97HZZPd1qU7GLybx4AbMj2JSNW6SAksuVcss9FNDFotkXMbxuXI+eGN+5+fr3lo7oCSgQ1Ggw4
1pNyiFAjpgprWh/11+KhFR7z8OQW/Vw5kQdIu6AMQ+KK9xeAG8HJngE5CLmdvvkVcP3Vny2uUSkh
ehDrxYGeEZ2tBoVMHCafpgH8qPaSVl00LbVUe4uUQd4RxxXruo/FF+EU00lOW64dnUG1EhSnCNyY
/cefwQv5sDN1gAr/UFjIhxUEZ1OrtQl0KE8nt2jHk1/60hYNgziZs6WJieC6Ef2yvtGjxi+W32JX
M0yS3iC1KdVgdsMp5z7YAc+OACWTWIq1Za8/La/vnVEseAPWIdLlHX7nqlLlQP/0LCmvPDb+0MDZ
9G8t396yTWvzxzvJEizH5EMu+km2T2a3g7tUEJBupS4fC6SGO7VaRgAVJVZ4SNFTmLJkcUP7Dvdu
g+kQ+ollQIS6WDw/X1YfSh+lsmh0kmcF6l4H/Tz5+7mvn1qShltvkNQtJ9HvIIk73TkcldWqljoj
fUCtninFVQ60uBICYbNkchZgN2H5UTh8m7nAjbPZhpNy+pwZ6qBKUQniFQuMYKZw/g0G1P9zeyIR
Vmu37ogGAMJ2LviI5HZ2/nS9VsuzIYZj5uPlSovOTfz4Ptjidc+Nrd+rUmhwEqLCTdqBJ8CUoVPV
A4pNH8ihCHCjMljTS5s+L1i5RZgAySetOAx0oFQnd9hVRFDn6DPeI2I64BNWhlVSS3j2OS0HoIpj
T56DZAOcM6kffSwh1pNmp2JUoS4QtQduVqZmiOBrmUjk2y3bd1PVBVWIositFhUkV/OSxtHNYM+O
Dn9EJmKNEueV7SC7VzcB4Y0dExqEVo1rkuWDPF3uuitgIHZfAFFCmlUBBqQNFF/dhx03OkrZe4qt
yFivvHey4YyywaoE0UbBDaWiDQSThIAb6YYhw8bcITXYIhzVxMihp6sCoiw0Q3ZBFAfF4FOjwRvb
kCMqjStAZzfjolUbdo7soWa1pkcK72Vt6sHvHmHmdDLdnjX47XfE1bVnMufq99HBQpyJPbL1+Olh
4JRVG8nvrPqpR9JvobCAkySwsyhJyrS/8DX0ab5H8U+j8xf2kxCkMLKQbYMBnVpXFe7e1Zng22m9
thMiQvmHosm9HRL5mkq3xpiNF1ZZ/ERdBSJMRDDvcLS4Qf4zDvnPh9rOnwkqJT6uBRiamvtK56kH
+ur4R7Z/1+EzWzyoDAwI0O8h0TltMRtvGT6jzsDbUj0HQtDsZbQpIgp75i3ht7J1ItNPCkr+BVX/
cCYEfTRYnxzsZwS0k/Cr+oOr1UHv8t5snlsB7IvcWRC1Ve4bFU4S7HUi4cMOtGEOvN3yIBLaIvGp
gbtADoeDc9WscYuG1PhetGRh7navVNwjrL0CqZCE0ntUk3CpXnkd2HEXacdn0X/kz94o3wzxeT/q
s6zxdNKkG6rMSjxXBLqMO0JLGPcglfhXSttjwnGZGYJkgjta6IQ7ZnlIhWBDnx3lyR+5lt2JyF+i
CbDIrf3+mMUsG0/KnyruLEOjR2ja50Q5PP2trkur6rDXTMgmpOf/3F3d/2YcZoI/q21gNNXfR+CT
RcpsoGRwyLGRu3wxScdGCWZdxSzIn5yh82AY2RekhePv8D7IvlJ99JzVJBoe4EjFjm44pDTH2wa2
G4LSHJG8kPXvoCdfZeGUjCUod3IlNjCfZ5zfeP470NHsP/wjByu80wRqroAFzjarCO2DPZB76VLf
qQvds1lrokzgUv7cJww1E7hjZs8YHDf7eG3jSx7Pa+3ATC9Ozd2+DXgRPMbCthrUtAZbZamNdh0i
Ne+1abOgc31JdcASxpAVY8awumgfILzy36211Ix0GrD7oH7B5CAXyEMkQMweCKRXMQFgrwEKFmvW
XYREgqt08zwNM2AEdmYtMoaQYDWHcc6N08xAkTMunBfKeFZPU08IEjxAQXqS+Kx/6EPTG5bk6dY9
kpXl1juR4sgZAF9l5JNbZ59z8O9HSt1YcdaUntX/dYm36je4lx3qJNj16fW1gMK7dpjt2RiT4X3L
TkBoQpcjTXfkGktSE8XBSVh1do/Ge+bFiwhoDK3om6IEwLkFGXr5mfM8x8wkRcedhd1N5gddWHg6
hUbjhps5P9HrrricSQLdpo3RuIv+o53WX/PtzWD2CnMyGnmz2Las4Lz3vBc9wHxNskPEQWJHxqGd
6yIjoDVs2sNCzEv2LQZNI39bUcX2jdrMnzgXijFYQV7zMfv60P11gwHJRZTx2L0cAwNmfScVYDDc
1ay0dJ3E7kem0wtcVaGMXwx0qeUi6oQxtKbhwPhjShno+jHRoZlT3c1im0lkXpm527/BWY/SNq1J
ifGZewCNOFp4ReOCK1g4tPIUfUdNIf1lf4D4/L/DqJoRDVYG0g2wtnkG9aoDWElitKVSFEroDmwV
sf+WXJXLQ5AQGBsPPNhgvl3y7NWAJY0dWcfh7oYBxhxJ/v8A8AW8hzqg2o4VZneILXNQt0LK4TDe
njmb5va5pG5ofgeZD+KbCGNSmqumCjaEEOMB55Rmj9IC/bLbpgYzL4VwekSnglmYSbgp4ZSvlW8l
bBt07Bo5x1UkFChNDLuak4cq3WMNmK3XWqp0f/i7KeXHqD9EiP8PDDIoz5VaywZC53rITtVS2cAP
PPZQHAC/LVie9Ff+AKAQdYMdhRlLZQTsfZQZb7aKqE+F+9tqgia9sgVMd2kNVT1XWs+rIfaL9lSs
1IsIq5tnGs+AP704zkFOgMEbbmASiU4ZK/NgYFfXFIEdgxwa6TP7yIW3TqW8BkSmEwd0sge12ux/
48UdNLCOhmAJClmS6dcEQAT1Qx6AEtYUoOvSeAPwt76UVf0hfVhfoe8tIMvAf1JcHPTep5Elc8k4
EaKGwoaCxSCgwE0MdUGT+MaEcJb6X54IMmGHnmadEnRSjxfqoziyP3VLMxtgLWpJCnFw0yikh6Yk
fR2QHPwOdyK+baizrYUlpxWCuFs0EgEKjbkPAe3o/RudLntpnTl6eiuajb+Lw6WgpgnZw4JwvH2j
TbFTItQN3+YFxD71LaGRRncpe7jjvKP3zfDsg+E9f6r52NjFU0IwLlYIRIKQYUBEi4cRHDzGQfgY
R8bDFOImz+9XckHxwXKblBTxUEeu77eEYIFXkjt2Uj5s3mS2Pkho8Q3IVZAVe/xZas53/uehvYgD
HerFaijsf49Yz81jhr08tOhyCjr7a64AGekodyWUOSoQRehwKDurGzK3DyM4SrU5DTybyBjopSk9
RJfSCgSmcFg1RQUpZyWxaCBMYeFW3L+BwN22wi1G6lD6lK6KBoJStpB+a5PrEGV2WW9Q2kG8h/li
yPwg/LWPhhoA12Rg+dayq6r66/fnG1NJ58GAh9y5BiNMSqJ3+mGE6aD+x2yx9cXuyDXQARRs+BnS
DobU+jEJwdkoenVMK8LGc0C4zSFf1d/SKEYssGSFto4ZaKMPN7ljPpd8cNVORs4VyncAZACgrkJO
mWuT1ifTceHNzvc2HvEZvv2T8S7ueq19LiVVeYgXYQjqcBWFyRF8K2ZOS5mtXaINOsjH0Mb8CTS5
V0UMZ3TGhv1Ka6VL4SCEG1Lfnnfi827/bZojVR9XjoDtMm9EETLpPqkcQlklhczB60mLn5EMgtSr
1sk9KVD7dBz8l0JloP43JxOmp7REzyPrOohbVZ8VU4J6PUQbjmpWi24KaK+Veo7oSZ0BP2eOU1a3
96qFjfliAeMOPiaGyMPL65gioSWTNMphzdtEiv5umeClhlZcl1/1yeHO65LXYw/JQqADZnpQr+XD
03Ru5LE6wye8T2L6sDW3N+kf5MmKoGowqVKd9FklODacddgcr1OFYky2DoUJembv8D+Zjq/qEphY
YGwftrwXUckbJH4IS3JD6sdG2L8GQo8LW9GC2owRl4Mns2Nqx+FpXL6ZnbFn1E2ZHOJ1MVZLoVog
Nff0L/vQXRk6mYBSxSpdeNOqVmDn/JtWhUwyMT1kwXT+ZRTzKm46PPLtIk1xDUMMqahggYhfSkcg
bWTO4vzG6P4dYc7vPaAp9u8qq5d73BUPqA2oo8hMbgN6jzAno+eD3XOlC7X078FVvm0Sbbanugs4
Fiq4jj0pAEoQ+KCARIKsC33k9HVqlutD6bUd6QrGLqmhzbeHS60hj1ni3qK11Yd+YnhocUvHHDLQ
2bnJDFLhD0nnsnwy4WAc30VDnoagjBU8vurXv/pZyB/Y+WXrWN5UynGvCLfxu5YgeUMAD30+/pp6
qIKD2BCYslu9bI70EHQqBSryRaUqSWpve5zDkC6nh+fKAedUk2GsZC5Mr4Hg+/8+bb3XZz3rdFhS
6QAE47EhfQl1hJmixQZfeXDL+Gat4QwbEa0G6QZuFsS1dbLBJ0kFvPOrQoKhsyEhfeSXsGu0Ebwa
IOCCRcwi1+luMMggy4trVJ1X2EDgbCoIlfLmNG5EaiDlSvIvNf11VVvR8qiFGQM1jF8Z1UJsSGq0
1J5//xSn3fXbmbGsbkY5p7mv3fproQfmet1p8OPBjI1bgLk1UlBZ5a+zgLARslszHQdD8Pfnwizm
ntxj66qxMxee36/DdqSck/ilxluC/0dB/CSTMaTbhc5qoiXGwBifBt7fa3abWSTBlVH8jMtmAQkc
gZigAERLW1IUWfXdZvYG7RvxtfHLpqzYVZ5ZhR/Vx5k9dQ0Y3m6DQ/rWLBd7xwj8GM/PY3SKajLf
bWdhVUUh4Ibgb3otpH6t9IC0cdAywhJywKelWEVKCUr2tCUD2Hs201vZVdlgufZ2hmCPhe5n/xmG
v5k/GO/Mfd5lcocc38quB27HIFhrOzvDMpi+eCt8SI85OBR73my+1RwJI6krf03sk8ARjjsyLyil
lZF/PyagA35jqh4mQDKErZt9MmFJESK+n6J833hdVZeuk+jTzCuRfW9nlZGc1/mJCz2gyYkpjBqN
H9Kw/VA2JL0gTXiHuNukRWYqPxdVaE/OvkiqfOyvuwMKv9oN8E0j0PIkqR4owXAcLe4cSa92iu3d
VQ8pJt5kblz6T0XlQO5fQFwovtiquzL6mDsBpyUSSu1YP5Lool6o8j0L2K7xmES5hgCGYzmNJhyX
3BRML3wyAANZj6sr55C7xVSDQTmC5GqLUlYdGCuCW1UaAYF5SLN5NL2vY+uM8eDq14khNSbQDVCz
9RwtDAC2ae7UZd2doaGmdvMZKUOwto0bCvV2viwfh6D3LV6YewQH3XnEQLicmM4V9mEJKWTPnV6e
CcPkSuko3rqncn5U62KJbKLiw54OGOJ2sbX3gkj369uWhm3fTc22e7IohmWAA6o0swGpq3Fa5XvM
EjQMYUgp0OEqsOzgEaQtYutXi1CJ7RrkgPc9WG1hTZ7Z6S+GCRWi0W+FaDvXWRU4/3ijZwHdxTiR
pvyMIQzaHaufWuvE+KRbsClyd6PvoCiZOIv4yDVWpZpv15YzK2Q+fNpoPx3GdX/jiCO/1BxMj5Vg
1TmzCUZ+6kp4sEcqUGbAGBni1xWtm5yq+sCdZj1iMVqYQmzWryGgA+wCJLmOOagpCr2K3ffuKo5d
iCxZUXWfowkL5ElMlvm7ZTzGvG6yutdb+H35ortyDy3j5jHE3pMx+ykJkO346bjRYXW6beu2X6Hb
tnohBPQ4OhDyE/kW2+qcEbDOg+RpPGB+Vj9BKAOfGh2ajnk/1UJgOPbRw9Ic/M9j6KEbCJk72q0o
f/cy+0SQ1H2/nEbXDXpXVdU6P/shcKzCsES8mBt5mQUYhNbe3hVgjPiHx6VzJoO3D+dXjuaxGlk/
DjnfbmuE9u4BCiBRTXXd/y+kVWgCLDHV/pSONbSedREosom+kVc1rstk9TPAzU/x7S6xp9Od2Sp/
2GNpOwuTZbYdm/0cy953/lHhyqp/B/TgzHr+gUd1W9P7utRvhul/HnYOdOPCWAi825z/Sim8YmnS
z0N9t3Eb4IcZ3jwhQ8gdFMInDlLhoJJMGtsfiSvIQ24KW3ZOpOr87W/LK1CjdXJJHVsmY236In2w
ywJIBqt5/LEirT7DJjWg7ROkKGyf9vyRoFZBE/tN+vXbo/0PN9gAp2QVD+n6fwRQmjb1lGpMzD5o
bZs8omx+2TqjZcrulzxEwE+h67+KnXN0K2dOhEORzz5tNhhFftjNmtju5iFH0/dnwhno0OHJlO+R
S7h/rFv62xppDKsXe8ry5ll497+rx6OX1/HUdhmf4jmyhrKbglXgvxIXVL7HfvhKjMpGNFRj66KQ
LimvK3sJLfwEMPvqCOBg0tA/Kxlvw3ppuoOcu6eZ4f35BRoJVAqYXYfZdZbFX4TZ87dMGGgP3bl1
pgtmqiiBH5/N5z18e1UMS0/z2XzGml0Y0TSzB7LKopPIjkRWqM2JzB3hR51fJtQViYrBFc6MzERZ
qrNh4D37LtyxgCGou5DKq1UEe349Ys7hvhK7ca6flE979UAqnU3G3t3WtwtRtFF1AodW5RPQyUrX
wzNxrz1cvIU0uyI7SL4rEvaRGfn09b4KuGAB5icN8vRb6yDoGNbmumAy+C3kBzWOPfC/1qk/UIUT
agRbfK1vmORIzmJldBgP3QvVk1tGzOhlW+UsvKw0BwmMeVy2B957J8PXQNn5YZ88NpHiHr75G94c
A1nPVziPQRvPieKh7V2gzWrX2hD/NWlR4t3GiGzhhkzHKWkdIlGH2rI/dJd0bPS2U/Z3OwU4+AL8
kdupMSxDWJldAIjQC8GOvrdAKuyUPxazPF2y2AO0ZCFw8vambfD3O6KQH+Jn+ONqdBl9kcmiqPwK
eD5yAiKssarYxfmIGlq4G56D7bBklfRKrusQRBKfLPijFiDWANcvJBT0y3vYp5BSwfREmvRsNQCg
SyFWFrtU3LiMyOKd4L0rooyFJlMJZupV420DME8pjIiPgmZlXNaIz0NItl5uGDPtzCRWp0M8/2lI
bqbvNiRxU/ppyaPIZIo6crhpJpTp/1qAQFhl/5a2MEU49rkvyE1VGOox+rUEAVtrPyBv85UGMGKt
RhgYN56DkPw36W/T8sjRB4dODMEQPZ9rAAzndLTT9bsLsNKMMmjtscq4kgvpzeWOO/eP6gM2ze7J
4qffFJ9dFTYaf7mmlG+NS9jPL9ieIfhHVQWEJoSz7KJnN1ig+sDfQxGs2OaK284CF9m8fLGOMIPk
m++3gNYT2kJsr326gfrOaeKBsoof4e5Vi0m0zEx2fUZ9xcFg7/XTsK9rPSrgODj2O4tjh3C/6Wr/
Z81zaxpkV5VwJfzJZQAKTPeOBnqm2vJZabBnTWJ/OGl77XrZ7OBiW2fPZYqB0qQb92qn+OsK4rfm
FGBBF0KyK0M8+DJAMzYEfLTyk1mpbrEad7B/pH5doBjC4ImCxSb2eJOKHubp9EJUEd+0K+zdz4jM
ixgLEhRD7Jb9T96zQ8LO4BjLoezaFFrgANdDrzAzO6Na5fRTSxDDKSY651wUGkWoIQrvYOmMZeOR
Gb+FeJFEeoGq914q49BzgKINCHSe/sUi84Bqj6IRxuJqyLwDijplxNUwHDaFFGNESj01tUR6gCn8
K1mx9a/eOKiGudKXSc6dERKvcFDUK/5Ask3NwhVZep7yo8SvObqbOzWiAzj9qfMbIBkPN83SAZXA
W8E8j6JAgNqmgLAxJbKJibdlJ4eeEqzkdIpUmnwWDVP0rKgH5T7A9spTmO2rKh2oaEWbvN7XKI93
ZwhFv5egjMvDFrKYXb21kE76ERkx+uJlaVGk9uK+NWzfM8vBjDpdt12ebAwLypu7i/IlBDl9zKep
gpQVM66r5Sux1ToAzY8mCQaHlkk6iyclMeO/ixNJq2anMpOi5CXM1iI1swojhQNFqQXqtfGEcwpc
HjwE4two2Rjab7XaERSxLPwdekdKj74osEY3PE1BDJPBcTxHKIjAQinuThgCAJST3Cl7lqtohhCy
Exb7C52RQkRsRg3jpX/2UpyP1UoYSdA/VbVMPmn4pmfsHgOgjeiI7PD7MfKk+osWDSJsugpJqoVY
3CBAqOMyA97SvL0EXvsZKkBNVSAKPy2nj8GN+mlILJBA9rReyxiKX4XWYMimNWDPVW4cuXUfYSC0
gqIJCH50r8NWvHtKKsgFFNWdVKO09G0nLcuzErsguSzRYuVawOGxznNW6hy8Pjhyonzp2xPQXniW
wz0wpVSRJTzh4XMND3BGup0A6MAuF2bnXOJmGDfgJIBLRQPBQy2blxlOfJALT2G9PdhV3U54sXur
z7et+I5MZxuwmx1yAKmazXzPDNeaWsm8UV7g1xBn2wkUEi7iWKBKRHX9xMtAgfTMwVSO0oAJWE8N
qnV1d/utf0mKSkRAyTQjsuPDCgEh4r9zzk25xPgxR2VcMguPWMBOUdTJqA/NmRXVYGJfozXeREmL
CF9G30AWoHf5ZmZoH28NXM5t9e3GtD/rFSZHdmExU+xUy6aIS9c7s3NtOuhmJ8ZQFWpJ4gV1FclE
Msl372iA7djgk+zOpgE3RGUlLc6d94WVLimClERBmYqqgLFgJhgLBwNZ29ifIZSlPgGfyHceRgew
ArnlnT3+pfgpJJAZuprJjMNBsRk8QmubXFCVDG5S4sL5smzOnZ7WxeUN2VipppassCgdVMzSeJYt
6jD+UVU31A2xUO3hxtBldqeulusBTYdEFHHJ0Z0y8wTFZSsqHvsXXCXKqxwhu7tMGhj79LuMQrOF
yROPasdeqSuKwyKHZPPw24zLAP2qoHxXmWj3n9eK+1T+WtGz24LJjv/nqn83EgPYwkuoeaGaesFG
FL3a7/Dj3QaYgFft2M8ezoqPsJxeguVcxC002cqiFgXP0uBr3gpEQD7Ksy6QzRh1GiI5UdmS/Jo3
eooxFKHe7CyC37tJYkqTKKOFMpxC7rh2sskrsIjBjI5+XonoTC3zJ3lTR7OnooiTCgHSOba4PG+j
++gPJp0vhjYpZoS4mhrPH3y2+LPtC9kw1Dj9h00jOlSAcJcn9EovUIXufFuJhaAP5OAcWOArcWj0
WAedQsR5UHYdT9JuVj596In/xolhceCS1PwcVp/Rc/RxtOPkmvLXXXdPXGaovweC5Z3kanlwGz7k
nzM6bD5b3ZNDV+iAMghx+QH/TC/L1DaAUCCLx2ghNlFYy+N/NO/oOH9aMplacsOyuCVzizRqQRm6
Q6j/wxp7698n3oaJXpy4hgfkZi9APgVcg/YZx2WewqLlMQEnlr+CJLV2Q2UZQ64zEFzn0Cg/nZq3
HnQtvDa8iHTdD5ltHFbheCSICLa6n31Q0Np8NCv/N8KLE0pmv41uiSO3X1eMwmbIsxPUnv6Jjvee
dNPTrA9Ee/E1w7Wdo0egVXaAKKZ1jzQnfBJ4EJTMcO0LE5owHnE7I1STx+bgleSZnVK0+6GEuAaK
atTErqdTBZDfG0Rwu4QtwVNvYiPfsVDnFkLWGW4kqv/cMKyNv9G12Ya7EuolwesmW2FmSQBz5G3i
tzxovnUL0opIvTFhSaTlauIUhjMWJZ+vFeXO0YkHOoEIAZB3lF4xkrjDnW1RwEtdMn0FPKjHxwE2
6BgSDWpArxEAypS7HtUR+LqpR3IBIWJSUO0fFUTD0xfi/kd4udesKvhnZSltIppKlRodFLee3Zec
EzeBn9k9o1XIemYr3W4re3jP/YqLEo0sNvtqyT6GfPJiJFxIS2Liyjud7nQIm23FTB/HCwsZXpdx
3oDdHYiJcjk0LJ2K9+C8z4tFXedVYbbAiYdu0NuRU7X4l0c7hkCqrr6fJDlHQ22/kLxI8mcJ9lxe
Kft1DlO1YADWAWYN9AynJl6VohblDIzCmrRTC2tDEV+AQTuB5Vuccko7N7dYHChgdWJ851yVxlC9
sNGjc46kwFYP/XTr0gQ+rdDD4t4f4+rz65vTT6KokdRmJ9/N7eeyPFBX2tIgJ/6PudzfVeUcIjFW
oSYayZVN6CyIBQQqwPoq0d8R+t1xn0+Me9dqvfNksoJki4G+IXvTYFaEVMJkIOmb2T+eXv060rNr
yBAEBP5OAjKeKgwr0qTKdK+RTTK7lXsmJFdlA9njTNrHQHiRG0qLu/743upmc8dale9RQn27dxnQ
Lalm2Xs/TGxGRG3xkwQMAZm5mquKgO7xyZqpv0//NbDDk07K7MAOw8ywp/MXIbJL3laBEXAyPhgM
bWF4H9+XGIwtYm88ETv1vytc0LLt/L/a4b2UYaJX1TSFfXjUV35Rj5bIqPBiK7+1MSOkTAoZTc58
4cKXVOxJ75Huh4NFf+hRNg3OAU75IbgoyOEIKvBAJpK6asvbDJMLPAueCrXC/C9h8tduY3moyPyB
yHxpmetGAAahKYN35kZdyISWkgAbXc+cTb2Z3P80hX1XnG4fARbKU3wGtlHUOYm4xGtV5IeTlYgL
InWKQP0aQGN+k/RI1Bnzuo8DZDDtBoqpDJ22oDmX/KchMiEIQLwbENSnBlGZQIFGuD1sCNmAc7WX
kjCH/L0CAN9/t571Ni/hmhvd17P0Z4EHUKm5Ul2oB8EOP1iwtCWTckSlspNJXaZdrq/xQ28CZgi2
rOxIOLbTMFqA1V9LzoVuBu6r3QUb3VXGOfGmUPE+b31O7TuTQcQOaLWaU5fmY9H/+1pqQrjQrAYJ
R8Ljx3MpWnzvlgPp61CEgTE6ynvHobpJAPB2OaZOgzfSbnAX8856OIfxBbo+vwP3/Z4CoJWI1WeA
y3MHSo6YG30Owk/DP/Plzntof2sn53ZL72U7uaP1bAYW5EBDBc4lAJ94LwtZONWoyTEouXwMbL4H
aOFG6h7w5R6cqnlDHAVfQo0ZyCUauodcNkSpD3AMAhiONtYASP+2Juta8RlmG5Hj3NFDOh3gBKIl
ZwXPJOP3VvdZna/4tFjn7wKMjXERT0v3zyMsjsHp6Ujhlrse4a9eOrcvyL91yZepY3XSJoyI8E2+
xIBTAmoaKYI+z1OSVG248hlURBXrIDJQqWnr+O0laLbqwxxbKufhDC4V1Ay8ddRqeUzZrgutn7ys
/aJOyoWl9LwwqlZke7ELZgXqJiKn9OQTlYmN5jEBZBUWesThjROAaoQCZIF4BAHpvZcEgp9eLut2
6BsqiEsy02V87e6RFY/KB2gBSOiBZDvrvC3FlplHpWnMvhxkblURjS+Djq+Hezk/0UqWJD9fioPV
y/hTqhTVrmaBEqHpiIl/KpYeOYE0SnlYgZiabr1HOxU8cactDQi7KyoHVdyeICfv3ysFlX6sb+S9
qK8P8kBrC6FtdPJLkm8X4ShZ6o5CYulIOqCfoDDOoi68k4u5iHoKjN3HvuiVH+d1xdN/m4XpiVQC
xOH5cjNVyCqCdeZBc+LCoxl4tWzyi9rs3Y+qwYhuJkcQUebEijbHXWfrrq6UWZG/3cJEQjw8x0+d
WNUx3FAlFWeM110pma3e7pWry2Oi6eXCEzSedkchSj1NCCi5NItkbAhi8RMUhi11AwlYkOjFp+XQ
Wj9WodP/L5Ws6WQ1AC8AXl+cy/flB+GFwkzOizYbSSJT1XC5HUVkx52sv5wlgN1c6wA5iKUVfHnJ
kyX/rJ4fRJG+Q7xDisE9/DX8B4WeHbY4DTmcSYIOgmRjoT+l54pmtrb2vwrhrbMwVBjqR68zw/cA
YOHW/8PRCBY3VK/l6VhXWg7EMKMA+PkDdKNYzENCH3Ch2B+9H4Par36AVZCnTeo5IhcMdCx2vR6o
YSLqMKJfLr1Z3XcwDKlwnzv9DRr1VmyjSJJfgZxgfBi7+hAhuRKzOT1JRJmfpVYRq9dbzv4w8LUc
mczskFHpTjWPeReLxqVyeNNypBSu74QrKZhGb3gId7NsCb5nm6CRQ0kt5ekXTHlHMYK1cXQX87lc
wneO0JwBYLDAblSp6cQemhoh+0OiqtKKCzidhhIOjJ1qrKy5RCAMTnFAP8XYnvZwQzANLaFbEjNe
E3fDMhDFW57vb3BkrIosE2Rv4e70ZDKueu4DgFbletbs4N4eloQ+qfv4nCUV15Q0wiBWohTLZlc8
DLPIQE4Ww10eY5QdR/8NiT47jAuh8XtqzyyRET9LxvdQK9SD6Y8mgm+VTWbEPMb/SBKkzPemOfbm
OQrLqLO0ptMYhLBCTiQyw6XwniEVOEIu/Pj5llmfWTsgoJm1wXZipbMtCNV4OWQ9286o4gEmZ6pK
KOQNldaWcI60bLRyI+nr7tXccU4pRblMAedhuOu4NipmxDWL6U5jpR5Al5MDOev0m8ANpQCH5wku
kmuUF64LUJacoHUsglnItqOCdrIL3ry6dwSleo8ZiHcpBv+a6CnXkHom6z0DRD642Cg9/7Ccjm/R
oKUhrmYbTPLm7vNtt62MN5Wjx0co/TL8bGs+IHJ3rBycZIctJNuYnoDZK6J9m41N9jDMiJwN9vjI
MctOb4cic3imkCMouVitsQGimfFyjxPW1+qRg/6EwP4035QFWQ+gsLCG6aLdc0d/Wjm/8IyhSejQ
Asd1QO/98vnQzsyLQhXGHW3P1wR3abLgk2T5MOj/KLfcFDPRInHynwB6p30OPSVLdvGoNrFO30G9
bwkc/k9IkkQ9F45HiU3GqK8wTpzH4KG2ukG6efQYYtfk2t650nASpAPZtgenSczCorRYab+pxwIE
akM+UV0WRBpbNcDxCbaH5J4MqHRcsNZMx8z/y7mBlZsQOwYMabXFqIr2CF+p7CP/8RwL8rL9xLp+
K4IGJq0FDQph4mql4QDs+lbBk+cdT8DiFJ/A66RqlwKWS+upa00P94J71VEgcMDY7/LhjUIgNdOY
4/cuQy17oe9PJwydSlvYyyDjHYEgUaDyVtrmmIbl26kTPLKKIwT8ZMWCL8rHvN/Cz3N4DFLVJN99
C4LoxhflCtv7EEXX7UFr9ovdWfZpeOI8Jhr7mwkzFKHdo8YYm2Yae8bgLIUY6xph3MqpVs3kMiRp
zcNMm3OLPz3hPIVe9zdBGm4FQrlv+xZ0xcNaQDzdJui+aWiYckV3mUYkglwTlu1ipfhjOEBz2+jG
6U9nOJZdKBEPk8GrtGol6yAcoa0LYZamAXhsysVpgeA9vJFLqq4sJurJfngLraKgAyV0E4C63q+9
6M7QmvwDaF2keBkBHAHbTrv25LtUpa4N9xNOxv8vJjcY/bdRsZGq0VqqC07IBpfIzMfi3YcNsaXs
pbbmFLOLxYEDwC73uUlsNabd9otrkxz1TpTGY2XLrbivVFYoswVOeB9hfIQHjR1NlDIXYsUnpg+t
eaDBYRvak80UkaacPuE3cm5ghwBJdX7En0g81j+4rhDqb7fHYyKiFuZMdBfVuQJPINt+vJGHsVcl
L9DBfTRyv5pQMf/BIjtGJhbuisDpAVyIjsi2uulXpPDrpe5Cc8dYsn1uLZymIwGsYRYzFJL7g2Kj
B7M//XIqGbgmOx43Uh5zeyLEBNI0GUK+LiqG0ySEvEls3MF3cCU8RmEIC3f8n5wuXH6V7zwVR38A
eNKdPsshDQrmI+HZHPagcrYpIp1aYb8cNlmjUrzJFS1zHyB8k0sL+exCbxt7qQYJlUaKb9pVqNHe
Qbg+qigKnT74aw+KgER5am0/6tVJ61B8StIui8z94Re6fvV2kgcPFTPuw+5zCGJp/OL3nLYSj40o
G1/dMIYSXa/EZfOhAxmKjBsDZM7IImnaF0qjgqW5AYaB26dCxa95hQ0LejV5s6TUVsBtRK2zxLxO
wDlW4VM3x0uqCyf2VsDrwYWO94MLY2PvMR3j71rz+L5rOShUZg6yODMaWNjrYJoCtPH5xnPt8VVO
1Zp9C/uLemAQNhvwnIr0MRYK0APmKOCc4tPG7QVIHIdXa/qoPnpT4/LQlp3IQOyNy8v6dVIbP2va
CYh/nCe0you1NhLbuxqyFk1dGNNnsxKeIQZLftqY5daBbpudi5JOIjWfTqcgKISCQlVOa06oU1zo
UBjVsb3w6EoQUwtyiA4xS1OT+SIrfFlj06PQ3AxgAqmspARdgo3zVQoXhBfAGQuLgk+HE1VHewyE
VxOIvsAG7MIfol8DYPef6WtZGVprNr8+afkqOY94KbnpkYpx6XiwbyrIfl7bc86rG7s/UnB98Tfk
OdrNxgtfSaFc0UsVTrikGbbyyRkzrc+yDearuRxZs3DBzdiSvfA6qmvJnvAWj9t89e1Jc7ZNm/Nt
v3ciZn6iKt4OAa4/Y4c++LN+0TPszknCxHTMRltmdzgOuQqHf1w+jABO5P1rb3Viwk3nZjFmCNc8
YJI34H+xoZF2BO+Qa02lFhHkXD84ZR1pm3lfRrhieJtPa/TpELArRxh5R3tTqUwylw7xjc8Tkux/
kplwmsOljXq0RCiJZWYkhMZ88DpVmQc7DlOoOrGwputWm2Omb6yuULeUZz00P+vya4iAONMVvTOU
8We8YWthqe7otf0CwqckCZmUZ0SKg+TuxKTXmTk2RClOJPJuw30uNpwdL71JSVwJl6+isx9l4sz5
AUgUoxvC5Me2RuqRWTUpNbe70sUFxdRNvrWca1s0CKko+LQ/F5DBWdvpiNz4Gs4v4fXC/ubJ5VgS
RJstBQdhbEEAb7jfiLijwNqPMtQkj1ppblZ30n1YULhrMb1fmHjKFSC/MyN6Z07Dwq4Q4zaKUcZw
rGRLrlX7INfLyXa9IlZbSI5M1TQ5mclP+uYKGlBnG+LnWOyP0TXGRclmQr4LcJFqF9F0OkwuyW7t
tBYLtFM0O/9eZJ9jzD8G5ksfVilP1EBcMEKLu5UPEyj+LJsAjNnQiyen3zJGk6ViUxx7+N335BBV
DDaZbFZB2pfNDmJBUlgb6/qmiE+4dMN3HmsNGS3YwxEovbHXLeVbf+kO+HVMZXHgOf53vjaPYFvO
LV4T4CFqu5hsrhNNQb+PAhZuJtvlzhr3uSZ+fCgIKgAAcNHNSNx0VGExCWhc3W+6g8YCYjLsjH5N
s7VLREijrYBFrA8MvYCGlAVw0zfMiHPIjTtCxNMETtf6ofuJkHFk1hlQxs5CmDsfHp+SOCzub4No
qLuL+EKb71T4niUm3DC8LJDBErBUVdx45CR7ulDpoTYXixU3SaRyPE/XfPdErgzjLJeYWo59/fM8
/WIdplO3ugX1St8TS2AG6jVk6stGNFS3mmooi1NyuBusrJIdRUpWTQrhQNDDYOrjgC+bEmIPnYqd
FP6u4VOYmvuUpOruyMWt2fwihWmBKqKxgY007DTFzo/T9J8VBh8WYil9cIgoUQf41dBj7yCV34ko
Pf16jPf9JppiIsekCei4tlvz+oz6kHsZ7ByjKF7aVInkju2r4EPL5Gwy8a6inqDYYhwWENmo2tQJ
tkw/B1dOLHf6dzK6hWj+F2tVH8fqx7GiWqKm+qlzGd2CZUjj54boHEx0GdX4dTJHVUHqRk0+Ne1j
5qft4NbPPuRpWQSqmcyR1gvYobIQZAkp3K/2ev3z+r2q5IuUW2wrN15m1oFEDBe1z/TvZer11Un9
MjonXsYEmXqnd9gXvEmMq46e+P95MQ9+XaMO9rMSDvJzE653tz3V5df8NyQdYxJYbRWBEmrVOSdD
IV6Dn4QuMIqnjtAPp6azDxWvGIOoSOkln/HhQNbL9mMgnj2axJzQuBqe0cd+DVl9Jy1KwBGZJfgi
qH2UBKMtU5ix1rQ9t49m6yk3KHNLMWJqf/4YtGjiv74kxrR0HUHe0v/dNvPRKAm8kuleokgE8vo7
y2HN/2Wq58KqpFJ9K7KYvvEaN3P01U8XfCSTJol+sTo/Wg/j7iNl+e1cmwKa6BHsWb59RR4P0eAZ
GiTdvR9RYuzVUEpOYtzQpANaYaQl9BZx89kkX1RtBK0e0PsCMYr4RYEcbjNhjmqQa9JP+zHApdbx
ZWbLbBlToDD+d5Z3f4iuPo2ffJzMUuPHig8BzGzoTUUUYZEIF3zmNx9TD12KLZVGZ1Azy8Gakh2c
IX/NWGjYM2JBWEUJHCo0VLPCmSrgeTF0vVNhd1TuZA5Pph/WjmLlRMoKG9y3mtfnwfhM0FcqR0AQ
E9DK8Pjjw2l245LQOIYtuk+pb9u700Fuv73KkkelvR5YDxFJ1F1Toar4LWFt+U/YMwpABpTiu1A9
0KjXbXC2Ht1HzLYcHPLL9IBYWZMOSx8FaHhjfALKi7s8ra7nwsE4OjYCBMx1I9XuRC0i9U4yg9Jb
6QcDxvu4/rFCJbewptgx5LixO5u0T7CcgnX9vz730mU+q0eHzlkDl458CSCkoBBYKYOfjLmY+RdS
eyiWEbidUw3N+cZAF5GuM8iB1q4FdzjqNiyhz8/VDq9sWQ1VYbbA+A2yg02GBRlBl2WqJWWsHsKy
v0bGBDmtMeQY4lsIPfFFso8DkWl2HrOfvh28P55o38I2zG8JJXCq+Z1KZTI0qXqIZ6BGnaYBZZP8
NNsiOlSuebBR1MC0ThATp4501XgKqiTo2q/iVf/5ZNbcyTznnhowePfT9hcbkPz3eSwMgCmxM6t6
UjdJdW19tiCTUeqLfYNjXCVWV/Yy3eVBRZuX8/cU3VH97hfCbFPLRSBjhnVADB+9LtQJw8vNYjDQ
bywS4Rlfh95Tu3U6oEdN6b6A5loZEVpIC1GStiZPli68iSFu3Zl2VSMRlYwvs1fWtPzQdsK8FiD3
lgr2vVoeuuw3cOknaRBr0MEAsJPgxS683KTvcJtGYqaCkyOlX5bt9xiyKNDpBB7Oeb7+llI4pcb9
xDXYNbgqAf6FeayhCErgIiYhOxIabQ2+RFcKbozazpEQtom4jihUnh43vPAUzauC8BLq5//75t/x
yuA8o5M+hdCQ8+tOt6JxTq2Z6FDGJs1DfrzPdGtGDXmm6tKiB2Kc5WgWOEjGsyQfcotCxcgJ6XRs
qYOM9163QvQAZ9i1qJwaiLVmBgT+4eIipDKYJ8AMg8e4kPW8z2SwfHnMI/BHfVrt6GGmcsrwwXOp
ny1sZGEls6sICO1Ss7gpv2W+8pVMQ5QfN6zy46libayOS6pO4vArFiVsMnRjMPjh7uWFqy8P2Zpg
BT+jU0QPRINYF/C/up+NlBdEaNkgERV7vPcrHco+NICkvqlwVdM7klAi916mPU5xHA8ySruubSV4
PTuKqNDhr2LcYU93KjB97LgmkxZE8U1yXixOPjzkHS6/V0PNGb7WlP8TpFqReYfjU8Hl0VkAdPMS
F2RwQNCHZuLV9QeYK0rd7w0ENDP0JeQgcJuN43spWbtxY0qp81hMQlxaI99q37MGDdRMSHCC4E0l
rw0wKmtfSc5M/lLMflKxGOfro/UI+hDdG3z6qYEDok90QZNrbFd340FAiPB3rdgrXmosJOtYEgJm
hIp4+J/AyjRCv0X8CEfHcPYknfgv82U5kiPQhuTinprPjxW/PN+moDdqo0CG1Gqo6ahK6X8UtpJw
AMg+djDwcO1oyIfGpr8/eCHtOAxktwmwIywHEYX3ZW4exQj57maoLQCmPg6rHQ4Bur/o4lrO9KIy
Atfe+h5C/VzhvEVPHtflOQpspibjGqbJz0UIDX4B4pZHRFJkTyIkXhw9il4JoKmndv5oN1bv4YpQ
2fppXmjvK89qSPB6fzvTERYNApnpJijjlUde19Oz6jI4CkY6uj35QINDQiFP2OjxjBw7nEBx9+xU
SreTP++DXeYZLAEzs+tCbdAbHUMFosWBpn3JN+SyMRfissmDOIJnA6YSyAWZMkYnOkBdDyZfzRVd
2khf4qF9pQ/mjwBsRB9aIHG/nORwkGfZltgARQqUMhlUIj8Z79Hi0lYGpjM4TWKTmDZkCYKuPw8Z
nn44jwWckZD2/9UFUBhRw1lNN2Ls4q3mMfCvVwL/A0QXUCPQByhO9CGkj7qBi1ppdIvEAfzIyevO
526kc3C/fli2axuEY4rEVVbXe2mwWRNogG3fLC3l0nZ5Opi8Jn2zrT6XhTe94XqiqgLFg0BxDVzQ
b/xLGzbbnZP/+iQsV4p1hk8WWp9Wuspy+T7/H1diQYzp/6pLBP0meTumnfSjXxOBDgzeUtP3FLDJ
XIuAFArZmqXCEH6CQg2dZDr7xR2jp2dyQDqZzUiIu8qwSkWbBv+bOVwlKH/MsWvzhMJU9QyqwHzN
Gq3Aag4ROpOIW44VkUK9saV/8dajf48gcr9Wq1KNiIZrKAifStawqUXNFCC97QhQp6ISpbPkFEAw
730DDDGiJqtcgv8c5yOljbSMHXoymQE28vemNH0Kl2DykxEVdtm51Qb25cP2hCu65C9jBgxJmEpb
pB8q6YQi5M165Qnxo/PsYuMvarH4y2DPPaX35zi0K+kzLd9URs6E57jGyZh3qj8UxrYQ4bUp5rhG
1YzrcsBUmUaRiXV0c0jKB2iQaLEwzXzftsJdLw8fnWxswUylRGr88+cOFd4urxwmV/nC2uLh/vHa
LZtRMleUTGBfQTxsljbTwarvho0IqKdK2EA0IBHGrxw6tNYV1uhZu2dphr13L9JmE+jrOKDTkmts
FhLbPyVuLfAMJyhHIYVUB8mplnDp+gtSG7Bc3o5Ahb53r8ELVmavPWPDgsXzW1d3vRsRLwoQuyNs
Q+w/iOZdggNvMh283p6eHk0OdZ6FS+luLTLqpM0rZ3bCgJxqDkx6y17S/QbyIKi1wYlU7h6BJBrE
rJOp10ZJlJXo8Kb/+Hoevjn1E5n/Efuww8HDNeyc3Ij6sU2WpItg3Al+Za5+xI8iKpfGVapnyeQe
9EJGcLin8DPpZbHxXuGIXV9DcfaYlbKDuS8p2niyC6GNk4Yy3dwOi1pPyJVVVcHRCBOfJjwnypVo
b7KJvS1shwSd3zd8zhMU1wbPkGFaq1v7WyeY4AFPm3ZmeSMelJcIsZYezptC6sSLul5gN2CAYRwd
JtEq0LWuNY5FWJlDSiKaNDGec1KSnApu6qcMIEa37GQ5ONiavIu4TrNzBxleTMf04XCmSs3u35ge
NJgTCHmVmq0/1pxRpHAgnSVxmrBBUl4yigeny/vXnz0gMZEEDv/kLUSGG/LKp9xJuQmO/cxOCQXZ
SMeCR5zP+nuRLdBhsQgElSpDeKVOf6EMlbJYQeu7E3SXCsQ+PcZr2xIM91QvBWTJr73Tx+6datMu
fOSkSlSLuyKyXIeL+qvtMNhrnWLuLj8Cr/10o0xexHF0HD0n0kWyltzIN+9V/AnH0Ssu/HgTXX1K
Zn39qdbRRckaXh8zrDxn6jJg4zM7pRzdIduX6F6E5PA/zfSMGc38DoBHaX85wAgGBhF2tfv/4Ova
boBcZbYsIMnuBl32d5FJQwqSB5Ix8VtmOhsa2Se0O0K4LFxYZWKPIXWDHSlSCBGQ+iPmM3gUyOAx
ZfQ9Gkj1AWUKBG01ax3lYBibC55GsWUwnZNa76hBfiOFUcuVv0D9QQcSnWBMaBZpY/JW6OUM888U
x2yRC6DiNkP8UnKR4VDdYE0ssnNC4sAJ8CKygN0XgOT0TEQEUKc+AmnmyjYcRZ1NAt52SMOE9Gn1
zOjP0Uc6KydCOYiMVxLP9wohL/D0IExgAtoBT9rGiRYPKtc1G924eLuGp/rHNoZd1F4lthR5oVTX
sHjVMtFDtKbRYuAILd/L09rta6ATgl5C/px1aRlreoaMIFGctyKfYUqg0dC9zDCLetVLVLAEbXNK
d5+Esqq9jgFeI06ldfEU9Nx+2g88V6WRRFmYZCdtGScyDIxIymsjb9dlhL/Y9P0cl8g/SFS0gEg9
K3Id7//zyhtbgkYGl9xmejjyXnBczfgpImBaJBf1tJIbxBpPNySDfIp8Oj0XU2/l/NYJAPvAFiE1
R3433AQnRJt54SgUnKYok9GtDc+U0ubhHaNcI4I+CBVWXwX+JMI55sebFo8AVmLIwjZbv99JuuKb
S4kG/bYEoQXWwLi4sFGu8MWm3Dr24paFK0fGXAg/7cDkVIxhFcG6Jwvu7Q+eFmyXsea9+X2NVKNS
X5NSBb9T3SP7UaovB5GVGJI9Ys58jWSNF/ZZovi0ArxCJqc7LUUSJ+/90IZeD3H3mKVGFMnzZgeg
/DF7W0dtmpCwi2CATgPIaxi02HASz4xXt0XGZSqSMa3SlGpYr6NspZNcBhl78AJx/uIiku9Ocxpk
ecb8Ob5shpDanrLLoFZpN5coeHpiWszxKWy28ISs6z3oX4/A59lNg+Z8AXWE7MDFM4SB305WpYfr
5U6O4ZpZZh7bl2RZC3/YXX4o7OSum1+E5Q9JPjTIf/Qj3upJZxQalxeGLbaGwfzjoEx8s0jJB6Vv
rk1N1g8MDZH8K9ag0WZfrQx8gHxM/heIpLbCUpfM8h90DoiXo8MdK0jcPKLj+Yo/LyDbr7YiT6Wt
/PFqDzxmSmJjin730nVCPQPi/sMZtNGoN9PPsopjmqSsts/lsasdtgWIFJ4lLSkiTtOvS2LS9rPs
wj/KkbB/roX71gt9+K64Src/XAOePiRdL/oVUSrFURr6frXUEvzQ0vGRR7GUHCXJvg/xhTcm+Y1W
p3pPAaNbojBlpi3bVJokBirX/Fzun6X7FIIYIGW28zB5anN2u9hxn8MbvZpPMJava/1kvrl2Dq/O
mWVrzTKSvxwO7YOh4JvNzL/2h2cHBTDbqKY6VuxTTmMBR3nEOR5ObG4jRX4Rv3WcTaHPUaDgYpYg
OFI2rrdy+4+hf2nLBiTpbIBruuFuw1Ctbq5y3+XA6p3ApcZeyN6xRLo52rQyAGbSuJJKQkL0C8L8
cweVPFgtfFTLY6P7pIjQC/bOt3LhqjS5hwqzelWCPXhP7mKEFjHkvAfifxQAiNX0u4pHaOx4sT2S
QjAWhgGGEhjhsE6ioW7WGE+N8E69a3KP3puQKhrQsQJBk/PlFdJv8vEKlkEyUxFPINg2Krf4CRYk
V5RzPTjXAAREhv+OMjtDtHm4B9JX7/ALth7vbCL6CneVi3IWC/HJ2TWQkj9th70g73SfCF4qX9Gs
YmJ7jZ8FLJIDOxKFjU/16gwGoSendDT0H+a2QbPcz/4/AjVLcH92+7ktG0CuyHR7//4/P3dqld5k
3SQahK5XQl9PFKqt+iKb53qIlir6GbGLWyxn0WEbn3JRYePH1PDVjHgrUDAXwYYz+6UNoDi5Uxz2
rySBfMzNwN+P8UQjDh2oWVEkX5E7e7xxpqQgDw4P82R5dRkz54OJBeG81jaIPcFAbalCSowt3mFz
dSxO4FZuEOw2TaPWS3KDgoPaakAfJGGKCaRzqOGFAwVLFloAVsCFH7GwxOs2CtoqKA62JYc70pas
qIkstkpOGsByM6NmBz6ihxh82UPUQcps5pXV8NEgFA7mUyn4Wa88GzbH/mZAqqvgZZFZCGyAy70X
rt/Q7CE9ONlDu+hoQGa64b9npKpsjwCiJoHO3lZv15wa/Emul/eG3eHjV3YfFNX75i/UovMd5DeS
OeoWIefxREe77U0bkOBc/q4Pz+iZBI13V6Od6DJemb59pFVlPCPi06bP2VFkr9dACGqbE/EWiSH2
jE/m7X0oVbOQwNcyl6IPePU0/6CaqIQfxv/C3Xm6ShTCPEjiKBEi05bA/Q0I9JPVvl0KDwZyR8O7
sbIDqrB2Iqf4OUxGEeGChVfO9QRmyjLT70G8XQG27CRyx38O5RrR8AKhPN77D+dQT3byId4VOeUD
keD/BaVVGBT+x5TuT/rO6n+xDDlcEL4z7SNCzzrxzv4wDRW18O0QH+EO2K+peAn696MN/rUH6DGC
aJoQP1ptw7ttRSCJg4DBrWq1cmEpYmgpTUZgizVNSFDU+6A5FsOi9KWBgZfem7WITpLq/WqaXbvc
diRgdkB7kZyfOc7wcvW6n1Ogs02q/xaDrvuweZvNfGx5Dm+erK0RDJb/VZv6Y37pDyt3TAOtf46M
Uu26CQo9wi/z8TXvDc1NXrFhwear8smB+Pn7cVy+WQgvk6/gup8idnjQlz7U4lW7VonGTu2mq34l
9ANq3Ry08y5ugJh6QNlfNA3G07IP0wkCN/8PPECVjj3SHNi41u2hUilzAPuq2eW0/55Dl4DlH5+A
K4LD7XcM8NOk/8It/mTw0UGBDxExF0HgUtESMVTzwfLJTwdzVG5Wqq5I6hf+qirdWPGqr+DJUEEl
FkZjbxZV3AmVCAVgP68TquPFYrfiy02xBuVW47Q1Gvyj9ET0g0ff9CO25tJFc1U3+MlXPAXjk3zT
LJBt0bfX/BS1HsiWW5Y3E8nRokEI1O162ywxLA+BMip+r0MjYIO4f0bMAynHs/UH6XNbztyNNe6v
wDs5YrLzV9fPAiJfRa+tqG5qXR8TNiP9LhGK8iq8dJKFAX1joHB0aAXJtUyqlCto234UsO0xJaml
gO6C1B6HQzd+ZTSmKk0y0aLUZRUV5ywDkZJiVhDIq69iaytBTHzkq26jPRGyAHK05QkH5v7yARzv
/Vw5i5qw5lzDckeI6KBGDuAyZXzDlSZdXoYMAvdT7tHRVaC4SuiSUyG07h0zp43Dz9MmObO2N7iV
5kUzxnTLqKinhN5ZZqzFClzdVGt3lV0PicyQDOjS2+FHnChuWFvL7BxMRsfSsC1nbostZKnXi5Fb
Wi45c3AW2PnMCAwDvhsxOGvtlUdg7Tq1Nw996fofZsxvnXXTUZyrOAOtWlfM/1z1gHDSNvPn+q0V
XipDeATfR6coToVV2wSdUDvo3YRv3mOhAcGTZqMG4fl3ZaW7rW8S5VkqByyqcmJKcAa0pA+CRVQ3
l69FW3YwrrWoqBc5ONp6uWncCjictiEiYa/n//zLMT4U23JnIzwj5DiJJ2VUhUDn97d0TeC/4LDI
KhVi3uzIY7c6k4EC+KG2ezvdqt7QLAbWOf3TJhj+wenP+96dO1twBl2wbtDJfTcYi3HWflQGv8Oh
tUt0csMYFPc52jrzzE6M28TfybGMthD98UhgeJKiY6TQCAcNbXcOysd2tzr6KNfeeoNPyEQ9qWio
juqXp2owGLqwbAN5kZuMj4lKVApFbfQAXDerk+y9svzMGv9X+sg4rxZ0AJY678gcGQXnwbLe1jNn
1qS/WeByz4fVd9qvKFECAa2PvIiTkBQLHJuMxpEU2KB9KUqgvYQroJeWtNMnI/TY2alAaAlz/usD
Lpg31EX5zS3xLqhNK+3YTWGdov5KlEKTHZoluF7b9SsL1StNly+KO4zcXX4phCLZoqja0T2OrgZt
Hcfr5hruDQ0vGkB7Gi8Qalecldxsn9Sl81i2IWHz3a/zJG6btF59ZAx5L3tAPHa2xEKFWnIWQPE8
WViCHjAIr9FRqNfnN7c0Y4g8PsJmNdti+p5N3gnNYkD8YS5CsHWtVF7gvRka8q1qasPfSkjlZ3Ui
blQ8H1sEJc29kI5+fFC013Agr4IzU5O7eFGxkZ2afOPDUd828S2wu7nYFM4LYzXkdxJOc36chDdY
9DQSfSimMFfz/xXyMe1+/ZYWPT4Swvpca1+b7Bfij2uYLDYdEaNVj7fZ8wJNbPSB664wjf0Q5l1P
1JFtdDXT6O2c3uLm93UPFB/H621ojgGQy50DywKTFS3VBv+LuxOZ0JT8i+ZGscD8kuMDPrpilAlM
PC0e35z4sGa73RprX/m16z4YsU6ldBCzoKkHqWauxvyQuGxQxsr0KQsT+py9/qPS7eAMcXb0WgMh
P2l1yRX/eB1pcnkmSM/mO/16r/77J7Q0NAFZ/XG7HdnamucTOOtae2N3T2GTzLfZ5uzyuS9qk8zD
ImRWvnZoi/HwJn6c8F0XoR44IAqjznv0yZ2kArpQ4daHRP7j+mOwO8pzGHl/HuF6XaE21VgA83mS
BVLgzEiR/915gnrt6D17exPf4p+QCqTHz0qZ+hBt1eUsfPi887aa5sz7jjM+WmmYNQ8j6mH4PcmY
KgrsmqXG/HjXl/PpXNpYGrv9TkUSSdid+fhfNhy1Lbe5XXnMwVaw1dBkrHm4VQtUU/DYWtF2TIkJ
crdjmfhfR4oDQbwC6coG7Z7LUnowAssK6dehJG/W43s9kN+5XzIVDp/ML0c6++VvUJGXM5Xd3pSp
ODlFS6ZF+iT8p6GOIJek8I4I/mP6TqUIxMH6kKwujlEW7GDxicSAyW191Gfo4qW8b+hYvNMtQ263
hSjx8IPjq1TNe9n668hvFygv/rrzajYbz3wK73GZ0CqIlnu7a82fegQ/RN//sajM2qOzSdAWsMLo
QU/a5h7oHXPxLnSqhCor/0jwqd2QUIUC6AXmCpzpfmDYHX/N/n2iIPzF8Py/DCHL5xzg2/8VJyvn
6wE0mJtntaVMnl8jjMdOGVMQleg67AiNT2mxQub6jbcvBtfA41pfEfUPU2n8pUXjFPmfOtqFiQLb
u3kSj50FW00afxxoR+w+WPYXnWEsPks+Mz1SSlq8G4HN04wCNoBFS+GGtC28yQZPLkoD8W5iwz5j
cxXOdnSoaD3xOO2HsMVUg41dHoMXQVn0URBI7BbPO6/W7h4n7OeU79SXHOU1hsGSJadMz5ytXOOS
p0fOsBUhF+FyZDKnNHB+3c3vJ8Lpso6k2ChEjGz/FmRRQYq1J66fD2iSSP15XElu9GTfed7TBdep
J2k9kzaAkF37iVcmLcx77Brph0WmVBYxxZ5cILP+hxEJe2OmFBa/jt7bqaS9TH/1TrNws2bFf60D
865Lw+Aq9f2CRUOvFcpbp/r08U12ch2ZuuBrKpyPjk1bVKkfdrzeo7nScp7n0HmJ4v+eYn9zpi1x
I12QjftYhyOuXZtuIvP1eCllFPEEkptUAE7AsH3CkewPE5MrNzzVFQJWOqXjtVGwrzSEVT+XTokp
QJgrMaGuduRq7ZSu0cKffsfVmzTNbJMO/8xyveKh901/r4aafnKaLuFbKkXpebk2as+PS2dXvUOR
OwtQuBbphD/nAMdFUsvuEdbWYQ5GkJVpuiVzlGdS5yEtf10kZwNCTMIBLUL4h/Mse87DzNuvKpuW
MbTgvkAVqF/KV4pjU9LnEUqBl6O7Z4kzewIAaOkv9OilisRcai9Hx45bX4Ucj80QexcPJ9C2g8a8
/zO5Bg+yHogFn8YKzoiPbZhn37WsRYL+tIWNK+TkGkXxU8EXXiWDE1gQVn/hNsyRM4U4PjwTnITI
j5owOa2ltAB4D9LfL+9Qf4SISJW1o7CTPJKrkNRm8WSJoiKZmKzpeaAU5MUJ04aQiadBtxsd+A7c
bIoDGk5cDAl84YsHBKB4qzWdB7iAJ9GKCfrnYeLfjTguIfUZbWt3OZoneGS80vtuSgCVq+SEjPc5
Dnlhi0Dlcf030O2Icte6XEdWZmP/+usvKRZRjeYsi+r+ByaOvG7yuWx79OIiAELK7pKBhOrznjld
oLwbQ9/Co0R/OMZ3+b5GUaDCz8dUzp6OxJiM2yOi0TkS0WnQK+1k1kAwkQbqZSEFv/u36xnr/vZG
6CWDFrAZJkp8BnFc5mHI0mVWtOrJnDy1Dr8yWAsyEDPB+t14RbKm4GhXf06WqWpYvOKG7Rlje0uN
EaitqCHb9yx9wqJFdjOtHj+ivq1jyYWlN5qHLj8X8KWx+fHP1S6lhwwL62hA8rA5wJ0i+Jvji+ii
4uufc56luhoOZOyDw792Y6LPiBljQCJayj2l3Wlo4PkFm3XUxfp7/sKdzrfKGrXSHmo6/37+HX5k
VVyM+3qF9Sof2jd7ePU5hg6QBgwcsriQKUR06/uGjUfVUp2nujc1fvu3Njo1Kmsvzv3PXmFUL5qq
uTkN4/TPE4c4XM0D5lgxm24Z/fLX1TR65awPLUlheRPqqib2aggH9JygxOkLrnpKBehNWR2jiLYY
UvA8PDC/SwCcNOalBotSxMytdU+dlnEvkaiYm0ocMPZFu/t+RhqQJPmGdRPhA1BQIIMTTg6S6MXW
CWeR+m/ZxYwIJ6eCLslh6UlVHbzEc47gXyobX4J4ZhpdpeW7yWK6vsti6qoyl8s9h+jtf9clZb8T
Qd0C6eT72pw5z2EhS4peaF4Rl/GiLEGKv2P0p7jIq4xAWqPKAOlTTG/rwShY9RkvNoKE7ecUjqAn
zFyVQJSqbYpRKtzcxIQwnhVdw4d+c05QN7DYnMGS18xhINhpFrHoo3xm1xAittlkpM/XDFSW3HKU
2NFJJrrToZSt656ZLyDRvmfOZCNnGQhEYeY1lTohF6Jmo3LDHTf1ByJbuv6m0dZlhphKD9xUB+vh
hxMiW0Ou+IVy7eIqC7mjpJF8QkERYgR2sTbwNqaZ2Jy7KwIT7fMezQ3fhq1nxj3sFdijH/tC4J4F
8U72xZr91H929La5ZWYvHySgUU58hGd8TPWyO/7m1pkznElleCjmS0M1xsp7tthSQ5QXgWcsKClF
AEEe2VKU1n6lF6fqKaSCtvpGaAP9GvfxOiMG1XvyAcpi4QZHgjUaRemNK8I5sx4pNdBxFm5ZjVUV
Sdth9wXjemTXH/hTmAiWEnCCk/nQfkrCW9YuzAKXPbW+8AXpozy1db80784SRUrFoOJyrqcRU7cH
zMA8Poa6mgjJ+aDPPOyD28Ep1zvz5a8n7OfTuS66+eNI7ZQ75w+ISJt8MS/5SRvX26536Qz7L0Fz
H3laomSyXJTib4m6PAxNOyAvNpMBicWkstrh+fN46UILfm9KnQnDq98Ji8iI9eKXrwSsjdyfNOpM
Mt5nWt3V7ZyHBIjUtyWpatCic8vuQKfpwNaJqG4uc/1ew602iYmgEkj3A2Zz3EwBIPQb6empbwwj
nnKm/lYUi6cSv6EGEs0Eb+TsEj/NbUrwC32kWkeocgtJZ28fw+B4rfJz4oecEny1fV0QjmEMrtgR
fpYd2M0eE3wJshuiK26JBIgoxFUcccCDb/AiMac9C58RfoZxKR2G4fo1HSxi5Bwwlnrl65jwkAiI
tqmwK2guMhLHklrGta2UHt6AT8Wt7TrvH5s/VhOwClDd/kRWJwZibicp++t33ecouSX7KnSOh+4Z
cYnBH9XG0UUd/3nyRmTgooNTgwDsx4dHQHUhCD1mAnPOdw94vfRToiME+Mmnh8DsHm6oXiPBomFc
0RBSyd/P+Y5zPWWPykbSxC0BtdpEuZ1YGVHMrTtte5So72oZK86s8PgxmpoC2eQ/EQHdlDLp5oNO
9wERkdvSgTPxDzsog5vcQjheeyenkblvHOe1QOHxDvcIz4wqUx997waWrTJtnbxy3cuPhfRqQttX
mBRObbqN3yKcUYQitvmME4c2N8MDxTTi+8bUPobWsEY/ZUUvDz7IX7pN5JnFjIMG+O05us6IXetX
tkwonhV2yLGKyLAWhPLA4B28/Z0d8htF/+Q6j+y8pQIadPRoYSJAyyIy7en+cDeKxcScaBxcxJOc
vid59yLpxgHk5ARhA21YFUNa6PeIL3mLqLCFkqXcWJUbeSgs+2bGpALKHc/zwl9/qiEEN7kw/dxr
TB7lUWpqugs+0uALTgYLdi9yTcohIuE4hrmkcdf9W8yANZV5ntIAgFfPqbqJq5CdnzLqu5J09DN7
8bfibv518thuun4oEb6XiJxNpm43M73Kg/6iEASTuUNBERSNiNCv0fid6ZSK2YhVZm8SM19QYlIB
QHVPQRc=
`pragma protect end_protected
