// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
ZklKG0B/IWEMHy+I8isNPetIMIL8IpuZZ/gr5cV5+NaxExDCFbKDykd8TUa5OJ7LohRHBJSnPgZ0
6mEMmZlWkvZZ+kIiUMtWuYZkzzSHdcwQGKXXdFaz9ScPuuS6ii/KVyrzs9UrubwTj9Xe9vXy20k+
FzwiA97PJam6Vhp5Q7eXV7qbR+kPF0S3FpHFMKbQJXCnmZ8SA4qZJJpweoTaW7kp8xkdaIwD/sam
z8k4vCQu4lZJcFE/HD651F8EhQXjbpxdjvm7peXC9nEUt15o35qW2zjKq7d4J9i89wSFuDPSHwrr
QvWQ+DUh4RybsUdswJACFJq8V9fZt/2wzQQbbQ==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
nBJEKvjYY2fPaGKCtjXYcntFa/JhOLl8xx0WjtCG9pPvQsfAq9oDiJoyBiX3dcngJ5f2XErVKlx4
3LGvk15Lz+276mC+NZvycAEY8GfswYqQE0Wtn/Euts/u4FBPcLoWW+dJ/SiEJ4l4p8LJdsqqkgkv
0/tj5YL61ccGUxvNTnRczFjC5rT+2idJ5BpxRaQG2sLfs4YQ4VnrZrGkMc3Htqsrw5098yyFlZ7O
rqimzyIyo3K43MGcd9UgvCZbgbT/euURrOg4PPwsikhTSd9RXGKdKx2m3h62XPPHtrwMZyLWZMxM
gyTF+DuIOo9yJGMPJdAg/BjvJT60rNB+k4bAwgJ1IPPYQUZl38A9ay4d5tEbtr5DDXTg36XTsq/F
aRKgFkQhImqcC4uaPOE2LBEY86fplOO4QcM4eEd4YAo5UYu1kUlvKNOTgibXhTBjwxG5x5LyMbMZ
D+ZEkzNfKXnsfwXv4LizJWH2T+l9fI/4Z+PIY8aYij5Gi5e5z/D3esqt/b/bZ80z64jxiF3GOq9x
cGyZ7e2pzuXDCaBhV1fyL10tKxmOtVdWKi3tjM1n6zZemeur6vxiQdCvRRBM8oovolSiC/YINTmT
jdEQzsZyPWDvDWKVapZTS37HlXdzwztxYtLD5jeeqPYEU7UutVaK8qG+1IuBC3tP7u8IGbhiuvfj
0z1BWcAFUsfKU08vUZJutBj+jlWrt8vWr80qI3YV3GvyZ2fBhs6fn+OqptK7c7SH4ni8hA+VD+9n
snfHma9i2nleu4cyGQwgXe3nswcWCiCtfEyLwHdDWKBsDNaa5w7rblyn5VNoyik+3bGUsmorXMhr
DpAirsQtYu8bgoaD+DFHJvU/mj2kL3F2aEWiHPLomLaUQW+Q9mj/HlK5Uqq0d7X9Uj1UDgMUPUOE
3jAfPTO2grvNj+OL8vlEdITRpUI/CT6CAbNeFa9JuOuoT1kmSwZ8wWGizsdhaeqFS+RLrJUeexgm
cb42MVykeOEUTQ1NdaZNP2UqsWTySY1teX/gYns5RrZLEwDzhNHX8Tw9aWHXEombV1KyRsNpJr1G
AproxPWMalrO+s9x42JvRzBIP3OO9oLpgLD1o4r99UHCfEPhEcOGwrkHfNV7nnvDvD0jT2UbGTj8
pvlgp5okx8vxvnLB7LUadjL+zmHMzYY+zrJDkkQ2UQu72ImlwQ9CMAzH2KH631Dugl+oA5b1crBS
hSduEP1dsLGxhm3KCcidBap+RIXHRUH0g7FfI3ht3rQf9RZlAi99naJgVUsFBgzO5oZFYsvbTyd5
7ydqbjoLIl6rORxq+Kl7MhyDofYCUus7VyE0I0i3if92q8Bie55GAmM262k9aN09xObYzYcSsOdp
IDinFVdVRVPMO+V/bENk75FxJH7OE/tscsZE9qLXlx3kMuewiBPHp1I6fdO+UWdQOLcGDyL28JYF
pDlwL9KKtfUlHqx9IeL+tHtHOkFx2TYQOIIOlX7CSHRt4IQ/DikExuMS+tgN+UVKpRA7c0rauSHY
pU2KTYjjcwLbsdMV/+xvSJb1vWxnsIN/A+xtE8GCNYZRdJ5lFrIZt2bOPplCB09YNsmhYbZ1uEls
KBUbBER3iNDztNrGyjycApshe8vDGcdAZFIzx2bLC8+mUMmiGxH8lz8yD/Mc3uk3lxme6PQ5E4U2
m2AZ7e+wBrL/yhdOmP28sjIsGufQCNH/mGh3BTkLCkYHUaBw69hDsfsA/vGvYY2u+0ByZfvz/wyZ
4wXZx6N4BEFbgiLEvtMo9FxKREGK8jSz7CyUx2678EomUMHtRMXteGKGa1WbxgQ45B2H8VuEJYpQ
fTeUsVYARrXoyofwIKg3z3eXXU2xoFWOILjyosh6xhvrCOeW6tiACq1nn7OEohO2YTXWDc3UGTUq
dlMyNth3OKxt2PysAgJr8ftYef5yWBYzmgMROdMQ+3rqIGWaOv8xMbYWQ0FnQLcE8hifhUEuF+Vt
e8yJRju7dUDoAfxFzF3pzmL08HGOUjuiLgSOrKVaddLoJ0OMSlKJn9ij6fLBafqnK+VIbyvJOJ9D
MT/Gxw/NKVWVIdY2+kl3rfWtaIyaepENhV76aZ6ikIefaKBcpHkBCkafxkifnfURyUVfA7znOwHO
wDhZ0P/hXe+4Qy3KU4wdkTZ7VnQVphqt3T1ZkhkeLhwVmyRUyZZpJLe9gQ8ZxTNA7ehju/z+2vxh
RkCiZmSTS10gHn5wnZwbvoMy5aoK+ubGs9U8lrhR3VSau/PydJKLNbC9qjWz9JdIhHQ3mEYCGtSG
T6sn+9fjSGTxt7sK6EJiLzvW+MCjIjGS3XCPg/nA5myOjM4TA45BoZ2PRXE4xz0LS77pOtRqs+f8
6ojF8H+bCDguhv/rVQm9JDf7BOuaJWB7nAKxYcgOBG5UO6WCa9rO6/58ZDIi7XcpqGPW1HxjtF7V
qBna8PM7aV5SIvdOGkHgBmz1CjGmIi9K9tln6lkmzczgA6f/XDUE8/bHjRmDDZpiEwbtpQ8h6BMb
L+mi9sayH1F4O07HT1ppZ57jGIOlIiJri7nzBjibwGtOUrBVPc2QmRMsFlBW9Sp5FhcZvWfVA1Ke
zEU7+lGMOUZ7C4yKf+PgkdvaWVcdo7+A/Lq7wiDal/5e8j43p0axrGlUvZXygvJ4HGrLZw7zKfbP
bZ6CE12GZXOGvDlTCkXLRR1W0q6Fn5aSSXk1Gd/+moeNGzuvnmePnOiHt9JT1qW0McN6oozfzqA0
nnx3HzP8Ev1S8w7GJYcWEknJ92bcZs/7WTWy5i/1NvpmjMRQetCbYd0Lz7nIHNF+g/ei/maQXuKL
LdnyCjB+47JtO7Tdir6TI2Z0SIIfm+fzA8tGuU48qwVjFYqzCjBb85+zg2oJioYSEnjNb66+tk0x
YfBv2Mws5eUbSqi8XYb3vmcAJIh0XujIUZxXMtiWxI2O7/bnaPGhcUhak2xlNLDBOD1JyOyfc8ER
itKM5F7jS2K0PV3knqNOM7Na9DgseYH1BDWFjkxtQ01VfLn8JNiRqbnkqCYKpqg8tJk/MQJURThG
5mb9th9P8SVYFC3d3lAua+VgW8YPW+zquHXrYx3v3pdo/iH2QpSaHyfZY+E8Y8Y3Sqp/kuyK0Ff9
wllRfJlZh7Z0miSfbVCaNEsP6gadog7EdeXYLRhjhjAoDEnr/8dJTpkhDAJ/jS7Ic9kcpoDIBv4v
43JyoVxBdRAtX/WBjEOn+KSAOXDNMvOq3iJ/Uad7GfdtktXmVg0hE2mQKw3Z1qFKwA4k7NsjYRPk
epSmVZg6AW0VIqEKjRvJYfyYezxCzIcFJulcyJTXixwRADn+aprw0KX/2FG0cQuh2/NKpDbB8PLf
YVjLYGsXXzwpEBXZeRUUGGirKFQOxwN6AbtvDUDckiVfaoUv9TDGYSc/VkjX/3b6gVN7bfWaEyUE
yQzxMGD2ckSzJyNT5/IWBH8f0p3M6facIvXfGHNQOzHdsa96GTDGT6LT25fcXoZ8LgsU8QYSN5IU
TrLFWwKFkeSBKmKeWh8YOW47bFIzuze4U3yVEKwLPQgglqpAzXm9qy9Nh9Gg7/31mC9jTPkmz+iQ
tgy94lSN9QYKyOjNd2sKDjJl5FC4nvusDrnr/PGnZYba4m/nZZZD7CQNjJeAY8/jK6dgmqdfQzUs
rlOaeDSmNK6nfMx02cpwM7wy5pIU/vyMqUsoF24+PHMvcSrb/qCo5Zy2WDa/RUBB/BXrS7aGoaEe
Gm/DLvbapEQ+e2zV0yKNAzV/zgo4pIT3jeSH8S1KWSykH0xXiiVywTfL3tWctamnOiQu9cSQlnNw
wuerY0TEopOksB6vZB2cxXXCEI162TQ34flvbHxBYqaPGc+rY2im6TtgoPlKmbE7euIzXuLzPUaF
qh+F2OCZBCPW222OnysmbVHe/ZP9tio4Q68K29NXxB5twXw8ogWmR0elIAbBhjgibsi6FrPVF5rw
EbLzoZmpy2tlxpCEeRiZmasfPTFrb6OTP5qq0/Qfx2WMjHkm20GS5jAAYhtZvIOeTwEBfNHh2FeF
ETgoz98uahQQ38Lgx2ShFIyYagaLB5c/Vz445azhvMKTyKrKoSwnnqsJh3d7LemlID67W4yg9R2p
KEuNfiEquULymGdei/aKK4J+9gOqYb7mYquiyml69McTe9KK2MuyjgCcZLtfQRCMU+aWW44Qd5Na
O/l0eCkEVfNGLnMONk2NoN93lPYjYeS5XkLCVVJv0Br1M5qqgymnIZzqk3aJs+A484YbWT5nkqLy
RY4jCl2Z2NSK39OKfAcecWml+WmDywUNZZpB5zWLFOeBSJwGfxJht2IRBugDdY6jpfdeefs7uXMm
eJGpK4mkm/tYaA5DwPPdUnKWp0MbgVaNNb7sOMpkeZcOZodYbKi5fi2UIeFMQUAsfifw1rUw2kcq
JynXLPvKAChAYn1LD673iY9uXJk8F7O5xDoSzbTMQ4nwIEpEZAYblLAFPq5cpBg+zNLzNnnJDXqC
jFBaS51gMFYVQUhToXSPakcKWPIwhO6Xwl+3I1C1fKLY0mg/W7w74P0P+0R4I1WiGS2htUKQx5X5
XhYpl3AH94NEYVrMP9Fvtul6VG5m/efPCgg+B1AFWJFe19H0OsYwbWdTGvqbfV4EQ4Zrbxe8VwHn
SSfo9n6Cdky51IwCIWG7YyGMe/uaz/suTv6BiwiKGoVQqCPI6D5AqjPemeuAybo3mLSiiX1mQbuW
LxoFK98UB6140xb1OikmvHqyS+CAZbKgBBwU2shY9HwCnnuyNpKNMhCUgGVrtvoV0GDmv3XeOje/
4ljApqUswnRstWJZ84JKHNfZZdLroORc+jjwNsnUuUcXeiIzaMhl0wAinfAEIDTiVqWFxRxe+1Ml
DsL0TdpqF4/5kXicZ72xnHgW1t8hlrV7RcSCtDLXiafiIC2OntKpEkkgDFLb4SVP714eluDPx8YE
XF3UeLZlP7OEvXH6Ar78gppz/BWQ8AgiLeCxQRVeWlyv+bhOnF7i2ZaULdLA71hwagtE6oD5esjv
fRbdfXJVgyBaGmnhU1imC4L9WY4eXDbUd6qC5WIJRa5zskIJy2xZt39xcNi93qnUCDsQLz/kLPBx
sWDy//dt0EGbMRqSgSbwydVEU/63eLHYGIr2r83WpvoLYws9KHdspMzZAulvLnhevm1M1cnX2E4H
jxk81GK57No6W2wtzCQg1OGtiE6D0WsNchYyk2YFOfkRYLdOMZFb/lUTc1quTDMe0IcELQe6pOB0
gcP6Bvg2lTe1hCY6sEQKhw6/tGKlGLryUW9DgKjpEkWxAPb5N0+k7uZKfejRaHtK7wYV3Ok/MbF3
ND0SN3Z6AdlF0xHeq1pNv6T/6X0tA8SWbSOrNjMJccwyekKUgDg5dtZS2Cp+jMrOSU4G+6pcJQyY
fUKtno6Wo+ByQ91k0DgDxFZYTjl+PMMss5FM2ywhUmN4NQM1FHR3bG0uuCJNZDs8L2UnQc91zJ6p
PNyBx1ob97/HadYqW7+1PK/ZXexAEfQs3JNSTxB9IT/72TgDdg9XW8sTgplRxtF3UcRcl0fY36Sc
DA7Y4QsJp5EljnaTqBqkskmXRyM/I55xwWbBHAMPpRi5y/Hg+6gkrRjjdsZ6juf6dl3v7UTv8S+k
HchMmy1tshQGrFlHXfS+Cd8NU0GDxKTxF40fdsnjkZiOoBM6w690Ea1M2u7BEJQhyXthRS+wqBpB
wTpkpp7hf3nZlaKmZJxBDy3b9tEssE8xlrMdOMvSZHKaHT1sUIWn+eADZfBOmaQAzgY/qoXzWqiS
VTg4JXqQd/Lv6EhLW+hbOLPNJEOJEJKL3V1VPyIsDaSyfGSQLwIirnNxKDqvoDXMf+NEb9Btrgkf
KXx2ZTzs/7mTIDyzFf8IcAiG0d//j1M01s33VK/T+Zj4FKk9MGuIKfsGgA7ub3etZT0xk8VINe37
pWSnIkkROidWy8ywsHMEn3SksCrutE7ksLtCzJBZ78oqGOxY3L3Z7qEMnFoyM3pluLPfqZg9og/q
CQ4hAiyrxUD1rEul1wF4Lu173PcsgLp6+fOWCHjC7pOpFvCsu6ny2bvGBsvVNDBjCHn+NSgtZbIc
BCzKHQJDiE6l45GqDLq9fg59010BmLvCaincHLNyJ/uL/+KuYP+OnE6qt5gZHdJBychvJ6Q8SplI
8yYPuy3drdFa9EHX06gcEaKzoY5fH1RQuXLqcjGR48QqSa48wad0f5LqMkjl/HZ9EG8jwFn7b2UY
WIsXQKuAdDic2cBl9UsftgmyCJimjf3i3+U5MjVgyiTlqpdPXdnjtx82hLrzxFuWhGWUzUi/ngTB
cKVK16i4GsNdPfyjB6b+feY5/evQTcuL4vxrqcY+1TJJJBLAKYV3eiZZCl4qYvEA5do46DIGNbH4
vDZvaYtFF7hEI2PKyqReyb4xUo+01HRDCRK9nqJre/eiByBKC4TXTn1CP5996HFFvk7r552eSPcK
Ot+BpRm0K5e2+niTwOLllTCMEPdIBTXh3BVs4pNY6fQmYS8UKht+dUEAokiJjaJNcwbTwnFrWZWF
PxSc9kGSMH/iScRJ/AkAlGv7Rr88aKCrkQWsZnJKqKC/pb+7f77Vg8wvSaRXyJUHAIq/1XvLHin9
Z2Z8SsoWYVHQPTnASrIJsVzdqT510aCdmssGxydbthkk06SQjr7yP0BRbtzUS9zVmmOE4xWLaI3x
pfCOcASzt7gbtGBZIRArlR7hYVhl93iM0ODXAJxEn7XjSm/o34jgCjgoMGc6b7K9jvCeEciXkF0o
2BZfef8ynTwbs/AhiHeiSi9fzt9jpoSGUn77aUA0yj4xVe+Qxf4vhXeCn7cKGgRFilQV1GgIX1vL
N7iieE28KQ6VpkLLpBq1aLy1WnOYdtVkwphz6UF3UeTWAKAcMFwTKqK11a5/lBKVIG8Hm8ioDijY
MQ6CzkGif37igmVtFahbuSPiAsiiLBwGl97NXlHP25bXshz44lKnDMy1BdiO6R1xC91i8yYaQFUp
/pkDOw==
`pragma protect end_protected
