// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
pqWykOXkoqEzJ0KOSE3bvWpabiz/46NlwJZUSl4OT2xXpNTCCU1ramII3QTc5yg+d7tOJaVcHE5o
gp0gx6mkxyPkGY6iqB9s6eFWoGr2qvX94yCwSMPf5hEmjDA/HI0glcoO0lfrvqQH/AfUMtPEhuyT
V65TX8uXHD0JM2b/LFV5k9HkQ+ijyUVDrTHv6iUe0QxpzhXPxMqsP8F8OjtmySx21VukdNukYmLw
W82XiSNXlKSDo9taW7WZSPLRcVMdKYaqaQ40vUrL1mnfc4a6M1o6mVSoLMAXqQwpn5j0Mt5LbN+O
rE9qfdZcIElRA6a3Rb9li7FsVFnAf+XZ+tbvSQ==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
EU0UyVDX14kBvJnu1RC5x+iZ0A3sjsyAt4dCvg7nadj8nhrxc5pY0epSigFFKDcQVJWMPArtDJk9
KU7K6DoHvnA2IDsx80UVQS+x3aBnZ7dzrNwYYp0jA+6+yc9/euDTnYQDgX6bf8IAQF/IxjLS/27Y
reDQx9Ls+tzL03kfRkU05lq1y6voEqvJ/iLonpgnZTcxzKCBO+uSxL/Uo6nOJbFyRosvtWKV8VWC
pktC8Zn+dLTWS8OU6VP5YY5fDVbK36Rc9jhnhgQtt6enYpJeHjHFGcgKoEqY/I5qx10Z5lxYk4U5
xyhG6ejosg+LfASkLUMeLWLDvnpwA935IGA+VxG2DCX04woJXAQ/fPKyuH5E3lh/93X/L8sAOSeh
NX1IWwpQQxMJAzqD7ugcFIVQAii0JlbN84aqmrEJYPYykbwDtODYIbqMDu8SYjxi4UbGQlOOCnV4
0vpckvWFgl49nstqyEwfMJbajjHnoWPlCBNn1D/HuC1w8ETPMRVP0NUv74IVmgUZRzopUIi5kLMp
IdCP3/jHHRsZpmGI/xJTTuG0M2NYUkJaItrh9UwTsr62D4WlTSMRwobGmgFJJcToIZm/EKVcUsRR
NnisgqegWMsG6AZadtMc1mUP+Qgl5/BS9YeEnUzw1pBUSZFgH+HquPNeIAohbOXOOpLK8yAbsWUt
ssL5TNvPPBMxOkfE0rxZ46jBK5WMrgIFK9/siqbZPSLC+nP+zefxJ77ECwbrog+Ab2t5IKBKarnV
sGsGgmhbyAHPlTQDkPD23Kp3nuBtoUNy1uCjksS6G7P7YN/Rv401wNG0twv2y8DvwjO6d6LTBIkQ
1jE7Z6mAxd6XHstOLnQOm5JGQcxQFzLuFiHAtEH8nrx5q6/yG+tBzrmBli0jRpEuUSWdrqoBuhx+
hcstgj3tFqTBb0nY9MpBDQGRIRFzG/B9aYa9539YK8XGhW1yJ2MtvkKD/ScYthX99dz9eZkLhED3
zmEujiLrr9LIsVuF7QmG6YFoX881xh+6LBe2eNY1hIjTppmq1CRZrrd+bkMnNpRlgI2bRCClecBg
JCc/KKqFL0LoiEZzDR+Yxugl4AGuWUc1H8+AKRoyUMb1u6JWtNL8/KC8Od98VDATyLoWmkkqgez8
GHcp/3O8Nk9I0wDSr2s3Tx8noUuz8Ojl6wIfT+63IGBp1N9SWIUnfizcsYjfaDewRHb5qbl59KFN
nVV2yKnVuAvN96UlXc3TI9+WX72jsqIkMg4UVl3Er1KHpBDaTIAitn9V7skY53PgtVvW9iVsIUIM
zkFBc4Zjcsz9iJGSgIIm6Qt8k9Fn52IkOX8ZQvhx5y7QWNOgrNOzW6ggwTpCrBcqciTNChOWSJSV
SyGyUVf+FYgRXRFYo/PVRTNg2Osqv0TmFbGTMq8ng7dI2nLlQfm7GOGWqVBwuq6ox4wrOTih1CfB
sJoTtGXpOGVBDegdpfY5IdsChB62twuMJB9+LtA9tNfuoJMfqur88gMmuDjiktJHFx+ztwxNIDrl
qmKkT3U0hQ1u0l8QjpOYGbtZjePT5N3gIqWTjqTkfmoDuwskhVkeuKtzbjLZqwxnqLrHJO3WKuOK
/acYMmeO3Y3YVwP8GJ6rVBuMD01WAafRpahbtxKkwbO+dbU/gNRfPXGnIJpN9IXPEIVIX6rjgvci
j/pioKMfT7VKIsE3lyKfxDts0iT9Ah45il+pbLmpCgZqihJ+fN+lSQ/e5FRHBmkp7VbWvjH26nBy
EYr08kKFLuTXDZh0KNDTViWRZbM7Fk3HLWEzeD5noH5oihTc4aAwGfUokNk/1BUpVN0LA6+MGi59
h9cQjfxcQpl5QVnfCPOytuNnDNTtt2d7cQKdopVhjUVtSsB8btcnQ4IN21Toi7Yx6FmRBgRsjOzG
4D+9tmtgYLSFqM/8fjYD9A0Av6+yHNiXqQlQEmsaGG/rUNI7zIyJj6aRNN+4pM4ITGJZhwH1autH
XwawpUR6D7NLDsfTVzj+sD14aqK9vYQlVahzqmLWHQ9Js7pZymigOj5tPZ1RIORqDc1AWH5gslT4
SXp+0kaF9ECDyd2q8+YgxA4EvL33Ss1XpTCgGcOulBWKz2agi1dNSqXe1fiWnY5XGS2G5YltV9vS
hDOC8v65QUq+jpNVVHUk4wAaRoUPh2LAUvOkVPJgnw1B4uysyyyAzzSokkn+KQB1E0yDihlyA15E
7Q6zH99JOj/h3Lf52glli+eYoI9TiOu1ivyHZeIn1EyMLETS5s2R0P3pSNEuPW/ng5KJ8G266Epv
bfGiDW65RSHv0nCVqlfpihO5fbRt4wEyF5+MXz5SKO8SZINs9V8MSmH8u2r0ZSiDuZT8P3yKbato
w6Hb4c7r3hHAMJF/w5jxsINWzifSCVYSMTVFJkV2Zeex8kfg4Yvy4rN0TISP37tRPnGzCmLknwaE
mO2lxyfsyrn9zwS17Q+RJq0sXUEqSwN9UnYAb4XjI7GtfKs+XId9SpbwgUDc8Q1uUtUQmiZ22M00
yLSvYXKuwb/phLus1iGBRB1/ZjyLidgS+9OuVRTRixit+o1mhS3xro1t/RjK+CWZt3Y3mPotfmyb
flcZ6C7lxi6yI84ogoyHDi2GE2GY6imYmY18Ksu53rUbPl0ROqOMQJ7kClp38EiWSe0uu23gUlnT
N+QbH9DByAb7qhFemCEVvdHn0aOrUY/dvti6idw0klF4Y/MGbrg0TkwzLnv37TzagX8kyz7+FLEb
rfw2YbC1WvKNjzrlVZ0/dTdSaYLnjA9g+9TO9HInbpqXGd0d45NT101uiXH3/UY/rIeVQTwA4rbC
BVBF8i8in9yqTvpFvDhT4CKaQhAIt6YhwQS6Xu4ObvLkr9ktXiLbbL3LefCV/BfgkoWbXyLNGjOt
o7cMKOQubIF5HKAO7DqOETX/0/o8QDGSAbuFmeFbllaTNhikWdX4IKyCCl+rHp7+gOVmvdmOQIvm
EqhuMPITZ/F1tt5aIwTUrmrUpML7OicuFzbHZpTMVlI0KGAOBa5NBWKN2TpBSl67IjOaOouh7iNY
p6V/iekrw8X8eKTycc7bN3pXEhv4fCwMdKg3vxD7ii+ux8kUNC89NT88Mchq24+4fmj9/wI/iUE8
fvl6+rTLUbN1cJuULrxthv3XfKH+4cKFt/gs2mVZNvo5fuUthWsq3OmxFRb4IF0YL7hDYwHYyf4R
2+kxiBWp6CfcRcITOi5W19O51AdMy48kbw23/q0ON1RaO7ZBPW5hMJ+8uRV+UQfLTxxjDKhpSHNk
R3jCC0+eAIGuUF+ISolEG68aWZqjOfhcfhAqB/5dCxiLK8UZbvrqUb8F3xllc6DDTFF+hAHfCvQ1
TKcWk/2MvDsY2mSIUL5iaS743Gca9hczUF5uE5S3JljnzhwjzOdR5UdHfebfawolgOTqRmqP5mSU
5HCWOQ3EWP/fIVmreT2uEbY/PUFD6yCwp+E1JRLpYAOPDOmsxbvF23UdazNe80/j5wNikQzQs21v
x1+/rBkhcby+kMfC1BO+t/D7B123eq+iGW2iUwLGYOAKQRlbg/odZyeKT6MMBGwLkP9R+CRea4up
zluereXnUxoqGGGCNnGBav74oLxrnYNOPq9rDENYB22aBH70M0z1+upp4OMz+/Z12pegS+0cIV2+
nZDf6XBz5R8lY69tvjFvmWdO1DTXmbwM/ustDvhHInTq3X0NJIDIEobcE6Hvmd9rHORvOG5Ud9hZ
Y7Yn+RDpLEgBj64j9KhE/IdATQkDOCBdxXpM/ADmV6AAFK3cRugXwn5rSNmdWbg1XoWJaAkOxT0Y
5GMfUGf8zshdjYjLDg3yI56a2c2Ckofe4fdsq+iTzdilA+UjHMYXkPvHsk7rGAN6qMdIpCGG3uhW
7sIB9TYMMe384/qifoCYMrwBpGl1SVTKVvtpBn+w9AcdLz3ZcdTfVavYtKRFfRag+7ixS8aAX3Bk
ve/aT4aFlCSh4XIhdfstHzrInBk7HdrNOeOWxcPmdPf2AGWr01v5sNHOUL2iC5l0W9jjpIC9uNJ4
TT/5vHrhyMzm2whnfwIwnXMsMlWBGqh8yWuzz+zCM4L+gqjhPUiLTnCKWZrjRYFaligHc8m5V8d9
I4XMNb5SD8HpCW7J6vYXUnt5J/3deKXd57YddXWUQr44pEPerGTeIUnSsVICG2Le1ln41H9IlZht
jk3vH+RIG4yWFQBHiGtHv8fvjIdBqGta7hdoDwRru+RcR0t0kvCBTGGIHiVfsDXW6VHK1JmVyY7K
Xza2k8+2rMjbIyKW+kVPHfjQEDV0YvSbMQzm0XPK5hzeplln/j/dt7aqZZGtnb0PGQwh/maZQpww
70YeEoV6Djf5KHSGORqA+TJMvDb9ltsywQPe5ppiBcYGauLR0qbXNAh3zkQs9B3NutYhmTVU5V9R
w03GnrJEQ+aW7d43EPMuLb3FvOdrS5QkFF0AAo8vj1Ka9YCMyAneBOq72TbzGrlhICmWhp3fPV6R
0VmrLlbbL82blc71jHI0S9cC2bNNV1VE90hXPgqyx/o8g4Hgfh3nYUmWT2UWH0HbqPIUWK1RzQ2Q
YCEVtKPY20oyKRXgKdYceNfb+Smig7d6XSpM8Y6C+Qm6PMHFELANnRhaQUfpdVKTWCx9wrPMwHw2
pE3xHfbOQroPzp1/2DBALN1FNsjt3fsR4yU1iwzCakSs+SHyFk8F8gPfAE5KuID3/PQ4q3Om/PCA
DkWwWi6ho+iDDL/9FmjDP6re8+cGAkuxb8Z/Qnx9e5ABw1DEVjULUCb2kp7U4GSJ0frHsxiDOXYU
CKLRjVrQyKKB6b7qGQFGYF70KjR2r4gz28nGkzfi2U+RRKYZfMQgiYx0+bZVj8fQc6cjI9I2zC5Y
FvLu5+tvHqUXINMG9wpoHtobL7kjHyZT0ZUBCXC0G1oiaoGPWDkCvjdjmzF6Srgn+XUL9NVfg2kO
s/7aQRMzcHI8+/O8GHwAAKtLSLq2c54/qcimPBPhqCcFIvn3SPorom73oLpcVVobgJQY6XARoCQs
QIaEFIscPobxSK8wRYoSRRO6L2UnMb0k4WShDQ2P+wp/yulJPoX7CagceLcnFovocbbzqtj+XWRE
cxKZHQYekgneVRys5X0eDMaCmvtovobUNqiMel48xvOvp9KnLFsuerokZc7uFpzOgNwhH2C77YYV
SkSekvdSg8LT6WSVY14AhBQ/GYjZN4hdPH2D5KQH+gzxPNdTXjrMttu60gqvEgc46cInHoS73eMT
pmZFZXog7KLJ6lZ7MpqrQ3jmC51Xxbc6rI7wBio0firQedg0khKjT7zFdu3wf3z7PM72rHJIqQ2n
XP4lLcrMwr8gFBv2STbrXGuR/PlfszvEfkp+PLVgm8dFCYM2O0UQ+WggfQV/thOEzqDbREsR1/ib
rPbVQSCqanwCcjT9XFZ4No4iIRrOHUjK6YfT4pedmTWCZJoc+v8nV2CK01mH18E/lp9R1/ySFHpd
FdTQ6U4evp4x/HiuJiFDJpBfNhLnCrjXQPTr8S592L6z2q4jtMcm3GePa+g/LneowFlYivbK0h07
NF91uzOUNGVQY4Tg4IAWuBPw9zWg5cNLmYeU1vlRSwgbGTZ6W95RszVBoOEX1/SBt8VLArQ0bfm7
f34wRnaCZm241jU0qgOMhdaoKG2ZPXRrbhZpRTOQRmOa678+j82Z7m4/nE7vFqzmlxIf8zYLpjzR
PK5nQWZRP/BuiI9uqxOeeZRXHCotSrelgq+jCXqQOzuntsfjfJ2V9kFmnCyY9JeZsaC9chRx60X2
lSF/UTmnDc4pysDUYdlNJar6LO9z5n5KzBULmwdeLRLpMOVcFAKn0DSmdsUq2U6P42rPDksM9F2U
e+c7N0svkEjzD0RH6G8VrTGpXOpbDNNuUzfvIxT1bmckmOHyGXtHqsk15L4EQlXHun9Nx5rKWjwQ
NIyiHfGjdGQqlXIgQTfhBqsDK7gzLmu7ExZ6gK1QTGjDRjviofEm916UQRSNI1Rjy3qTN6XofaP6
uBNlOK4E9qXVvAgHELvSiqjbsf9cZbMoHvoMIdMVA2+pdpnqtvm/gEdmxiHnU+BicmOSY2Kdq9Gs
iEX2BqwiLp26CYSDdK/w/JLzKE7ZrJ3cE1xNj6MxW0QHaUzcb3DucpWm6J9HGArqY7ibRwtreGs2
5+VPFwrC+5MG9SzJY3Dw2NcC0buDMJVAoyewfg3VBf4ZTHWcVJz6L9PiVKS7kKfX6wubbnwbF0pt
ScOa51XE2OnZQ32r75CDPOUD9RxgcKrXObjfOY92ZvcDmVoqGyY5tu11AQMLZGmFg5ysKO5uHZrb
OVU+prhTugkVNbVTt5kEDcatMLK8qmqiFmO1ypmseoyyDdmWrodAo8Ef66pZ0FZbroF79nQ/o2YQ
FdgAzQMfqurrF/n7YUyEbRboEJEtgtUr6oPn4n0ROS9EgPA3ZwFfnkBkAkl6BirekaZ9CZVUuS5+
9oBVuNRb9B18KcwpQMNhKhBO/EwBwBTo+1lR8D/WlfHGNxRK/+TEGUYR1ltci+jpeoB+LTpPNz0T
MJu9IQK9GBCZ7LlbKEt+kRz1Q6Zj06mhWkqDwLjwedHo1SlV6lwy5rnBY3D6KXgU+0p0oWcIsG2Q
Qn77O1rIVpIdycT3Lz5YZuVqVMsoClcrXwe9HCgRibNaG5RO60YtFayA5zPWijmLPENypwkil26w
p1ExTobusZDPl46QIHs2e0LRCufTPHTbn8MV/mtDkvBsOyAQ3OMCqu7jYPjtB0st1t/ldUw7HijM
gCSKm8QT9oRVylYkWph8zvwmjK5JnOmqu0JcAZfNq9zVCrq/7pC3/Ck2hP/8HZACU2kQxRrkpYPA
QRHFrQ04LgoPapxd1wynwd/X0CVte3wtuu2T6u3szMXRBzs6zC8p+OkRduTOsBdfKKiIkcQ0ilxO
lumwmqdA06JSZuRbRoE2m2DU9b8OkYG3YYzrl7CKMLYmHGtSeS/UxoqBXcl+ZHnaZupZ2aooJVxZ
Juf0a7672F2LyJGsjGk76slorGi7fiM3pWm3qy1iC/iAKIClej9c3YW95odhjiGqQWZPyCDWVyMJ
nn2nvtfgP1N3VlAK4GkfILnsf6sq6ATmgim5rITw/dDZa3uT3j2kTKheUsd+sCS4ovoNMoig8bKx
3LA4gfkHW7VNyPvhLoLRr5tFUaJ1N4d5MSgOXUdai3q1YER9X2hr8jHReU/1sK6Yqme2IPXd6YTp
x73BSiBSTOz96XaYypxriloXpGvvai+2lEP5p59W3JS74XNxFXlBpyMosgfzOTdX2H0KtLVZ8rSn
w9eSEPpFUGG9tmsn29d8jc9j88KAwzjm84dPofn6dk4kgT5MpQ002TtOHc8wk5DEYJs807Yl1QEt
a1NslY6lvBIa1CzDkMVD/RRKomJmTmLe34XUmgCVV/8ULEq3BYHXbvv8F2QAyY1HLO38hZmGL7XD
WA4Tbw3U7rP/RH+uIX9awp30wj+02GIwSW8sFY1SjHTU/Xuuqjr/zAbxv0SPzfdjbB/tRoBhuOro
1gYNUoVjGwcAJzGMUrOKtbS0566Hi+szy+2RpehDiTlGcgpoAaruc49fLviDqIt86oSruHjMKDdi
TYKlv0HGZ/dJhFLbFWPMqLDoCAQmR4iwdXt9KgM20ka8Pt1HfzFOe7eQxwmQNgT0wJcfpvxXzASx
1hm2whZAsnhnLyzLynu/8MF9kPhcwWdUw4MhjVpD7xxEBt1WO8LelRZTn3XrXgy+DyjXaO/58+W2
ZwuvYqVB4csTADzfeaz8u7yt06cX3FqU42GaJdJJql7Nxh9ypldxmTt55g2WLr88EozPOk1IRmIY
Ar/1P01NkLav5x97O+T3aJbpF49aeMGWERpGlZ8XiaIIWkgmcS6BjpGP3UzhDAF4YDRPScvs9jxj
tj0vA066accItsHbfqW0b0u+LErmO50el9mOk2GMYgMbrxAy0T2XEoJZI1M5++A6jL8ihoewXNZV
exl/Y1sqjY9+tzOHETeNrl8QkpqlDHotKXnrKRrOGpty8yT8wuDfyVx2DcsgGOgcqwTnhw7SzBNn
hOLFpmEL7sfbNopa2MPY99s5pe08cwfVORcVgmo02ZmX1mTEBVRkou+6vDcgAhyHZgNGDp/DrIlp
uTUJAPzD2AMP47YpgH80hXxy3V8vHfvgs3ykMfvUTJqgfUxRvH8YrsaraVIlzUK/p4MVA0T4PwoI
zI2cXdGk/HsUNo50PAP7MU++AHfn1s6ptS+6uIXlKkJJyuqODYuJbwP10HaLVrsRQozWp+t4/dX+
eq5dkB8UlJYOXL3wbDq1aANSWPWq4ErbAmLfw0CNpfjhKbbLp2KQbqngHGcSN1HynGZiefJ3kNgj
nnRqqr5aUeO3qU0VhOxztWd8Im4sPAWZvQom+pkuHAqbioKgYMLSQveMIKUJOn5480lUDRudk5Bk
qvZ0OZdg6Sde3ZJSO56z4x1DNAR0c02M/gjH2/d599D8ZNkMziIp73lcg0oi0aBq68ZlyFM8T0W1
FYZRSpt9HAbxKf+STVw0E9pFdud7ct71PCvFL5rW0ZYVTyDW6sicl1M6Yu9UmAS1Qv3RqnoMH/gc
N/gvbhJqEtM0VT0WsMqq5kHVF2C4P69youBdDBVmmChRNvsM1P8Fp8BEhwv6nQB2WF7daZD0g0tH
7sQFC9WCEcXXHeizjX2D4/wNN36o+z+IWSmLuvjNmIeLtzLV5MNW8nfviYjSxHYVnWi/ZhNx1l5E
eSNaC4hFSNdV1eESJm5JNY9gp1jFAIPocxXsy/bvVZ5T7jrzsQrs70cTAEBrqbA/jLpXf7N7JsTP
6wPHHLAaz1921iLO5HnIeptogWhY6V7TJh16wXww24UWbRHEiahq+rWthAGZ5agvx9uzBjLLtiTI
FPoc/lWV31UjFOQ9JRUztU2801J3V86tgwuIE/LYPntqa3FzDs92JAh5Af0mHjolQasQEvrWOKJ2
Gz6ooZSLYqzh8RWy5JucNEMqbRO0m1CWtKwYhpASpmGjKskJN5MEzm7ZmYwhdgt45ejW7gonjJAg
nUIG0w6ANaU90VIi8VGnlC3VdPh0Lt3vE62ugqjJMw4tG2BbuqFHxhcYbPR20b2zYfDbzFlNgGNw
3uHc/yWV3xuJXCxIA1bnjGvZqDdWBuGQL3nallemQMbRUGy4p3XOOCU+FcPkzU8nR8CH6zNbGqPF
WgdJ+NQHdXzILGsEbqB7DLmo+Lirr+IRXNmIOOHgjsehkeA4vHD3T3s4aKAw3HGECpQvfB0lDSg4
7HQloZV7L7K8B85RdwxxrVcqQDss4RLJOthy7ai6qeOs6H+f/moIh1hjonlLGD3F/fgQcRAmY+/f
qY2SYXO1vycZsmY+a5XKddgsIB/5v9rjhZgbyOU5zg8bN1A2GvyC18kzAljI4+Q8IiTRywWeGMqb
8328xT5isXsrkbxtQe/z3K2kXoPFFxWCY8Ge0+2NP7jB5tsmMfPr7dY9humX3vPG0TcynkgWVh9M
0FTeJhoEWWlQ3JWQLcp1y1qvEgq2VBtdJfJVaKXg5FK2ljl0iAj1waZ13rEx/kAsnMvNwpSyZYsQ
Qt5qMNLLrPiQAR3MvM3/oFw0ikLlPAFdtRIDYiwMfvuP58gvW7UDNufY1JehjHlXDnng/oXwjT7y
Rz5WG+QNLp0jQaD+zWLvuLd3Wa5/DtFwQwhIGY/5GjldBboRNNmpv3Vz+CB9bqJO5MprIxExsuBQ
rkI7Vnd0JjGg4QOUf9YYppNLQNaxrREiKV+UJw7t8iz6WkupvIBUUjvOLV8TL3y+6+6sVqOYW9RO
ezBYlpaTu5jjw73cY7y2H0C+0CQB+3GrKBI9bca3O0KutUBpRY8G4wxzKfvzdfUeujP0d7rAWqeg
zgc8S11nhh6wrZLsICV8MdczR2CWfb0oK/Qcl0/mjpIDfDn9nSXjHUAbRYDdfVLS+VMKxqWY7wkj
LHiISfaY1C14P5czITqK7vvZReZkPKa0jk9Vi3PFy39uxtd3AhjUtq28JBeEznCXmAum56H3uwsC
QNNHd7u6C4XTIozz4T1/PgqgTkrgCSCQz7cJq7F51CFt3UDEYtsBApcdvTMMjZ6Iw6W9ba+HMhtB
5/GhSSP7aGRHYHN7T8lu4kF+AZfq7dS4hVCaPtOOOBnDs8+KOGZ7U5MU46Gx4FXUuBGm7PiyFpQ1
veTj1LW8bUiMxR9gYBeFyykC3M8sKnBp+SYw8ohehwZNz7Z0u1hh84yZs6zVRh3NEetbiF05/3xa
gaH9lnx2Yf77LKywqfcbeSYBCXFsjUmQto89I4kT0YRNxSwbYWZydWpxoyOjxuJd2RaZjZ2wmj2+
V6iQqvS+G0T2m1pRmsPpJsqWEh/EhCcMy6YUxpzY29xYimYwZ74KL0FD0AajhrEa84lrH4tdt/al
F3b194/1yVe2vxfImePB8RVJi4jpG5PoFDcC5gXlTiHvqk+G1vvDkgAyP2D3G4DN2/bsYCAJ7B03
SRO0Zua2EZjJJu8qXZvTuhXtXn1+lSlJXsZIuqwepVoJEsxHvRK51lZehW3AP6B2T9eKdWXMh3z5
BTlYv2Gq5T5I/Rv5SGTompMkgqJ6VKSc0CEaMW664IVwK8yhDLLkbv+ptLVpcsKuUi4XN/kA/4V1
eXd2nCVPBx6VAXJNeTN9p9HCD5dRLhZXJt99h9LdUupZkrI6WDHV41Cj6XVDZXykbN9Qe9VC42BQ
PjzfPT1zrGBDnSo7Rf6ZOrn0lwfotXAI//qSjS2UbgQLwL77tKAfFnsJkSHCqP33xU5pa9Lzicjz
3GoKjSYwaEZJrEnSFG7caCXa4cjNY03Nf0mFqh0SCd/TXA8fNprRAoyEYqN1YFd4ugCqc2o+UPtW
0OVA2hCfEfFZM7Ep/peHBAgftetTZnSKPFfExYEmrVK03XRA96CQKE9+z4kAwPUwVRXm92kYx26v
rP4Bwachqn5RHYgoJN7S9t0il+GDW+RjJ4djXTr5/regkFBArCxJfthbleP5EubjwvqCe7NFLTq4
9CzzmMU8u0dSWQ52OtqGhWmnNwthKWhpCVk11a6+/CWMGKUdXU6BnLtVTdQ7GY+GVBgJvS+ooB0h
nCq0qT9jCBtO7GzfFdLcxY9VdJH8YKrga+m0ZLl6n565+Bg1yTzdjd441Bk2T52+/cGy0CDAs09N
sdlV4aQzR6fygLMkEevTG+ILFYz/hSYD96yvoUdB1n0aUbWUCZcPMAj4zdKqZKpQqgzZWIEZFfj5
xgofA2djB3m6cEIorT02dWXTcXpcrPYj0WWVHpNQUsKINpi95uXY3RXKTpRDEhOl1zqJc7OFFlmC
11rr5yP7+yccwZhcYNBJyWkPHAqfLFNbdx+ALwT79u/EBE6HRGMLsJlmAr0hs2F3+IA5HH2yZ4DN
UW7gOp57qUaV9qnJMT+hmw6i+nMOmJ4aDZZekZHSzwa39MCnmyOu6fdqpEJ8h31fBQwDqoXw/Pxo
yI+e4/0iaogGlsaUWUTAOgKsvf6bCGrEBIt3NXVgBEvVuDeAaTy5FI/yeIcRDB7VXNLlnhpdYI4X
iYQ4JhrLBopdiruJDoV22WaLmjKdIfAen6DfHOJnhoqk85lQo7ZZ/kDBuHQ9D4G0Kj5X7CYeOGmn
Zi7WsjbecdhosoSif6qheW9MZNo2pTrZvH3+EHFaXT0n72kTvXk39uPxWf1KhyVQD9SJUh9b9Qc6
Jc3X26B4VJ5ZzwkyAiBl2YY1Et42ZL7XvwSmJzk1ygwLv44fm6BuGsz+SM/rMpAsT8Lm+NxaTPtx
GesUK+bAwnXbHqnIclJWW4MKLxch8B4XdtYxgOmVSLD9+CrB/WrepHxmgPGkhshkPLtIFMoX6NXL
EpFaTka3PiCU5zvlkGYkfnm58276nQ/aawMNybCqwA8gYE8Zad0oQ0BTCgUKqNFUtMoMTbSrZ5UT
LzJUXGhnxIhYJw0uAcxKgaqtZN+9szsQO+E9bg9ftAkw6vDAIyrouQtkA5IQ+sPyIWmcbaWYTLwC
q49zTyrk8Bzalno9ls3sVJcH9jDlUbwHNn4HHvpQQpTs9F5LE1e7771gS3aNZPr6buVdSTYtVXWT
hhfMdFgoidhv3ODRLtCQ+J1IjbW2utk/3W9Q4Obd2XoBlNMG8SuC94Mj/pyIY19oLyYFV0dc4wbg
cyEfUXYngLXPpW0pY11YTx619X8lnuqU3OuqM/384BCyf0pCUitzraLIIo36O9yN4GNweJXf+tbe
Hwugq8x0cjdoYXzyur6wCfUxPN6i34W8Y6pby03uz1P/Z91Ms/63xjF539++Lcqwg/T/6EHae4MT
yII6wLiCYviP9vKw9NhlQmdl25rcfYqpj0AEc2WUfbiykPFk/sqkoqfAIJYXUFdMRA1fVhKENmZ8
yE0Do/+cRTSpOPfO0z3p4MX+NxiOZi8b3aTrVFC/rctWeNhBwRoRRh2uCFbT/odp+kBmxxwyxIxg
HqQKmjQ/08o4a0iAZaU1zypv22HZt1K9B3kbGcdSp3weHUcHWFgsxU5L5F4RHejTyVeTdtwyr9O+
9bQBmYA+2agv/Q9IemsdBiRwRY0PUJSSH6Umv/OlsBzAt8yk2FyZq4AGWnsE/4DY8A/1JTgNZBOG
rA+QjIik55DM9Rw3C2xACrMxonakYjD2nK6x7Le4WF00LhenQCjbReUgf6BKbC98bO0zlB+hVVYm
NpphbqeDuGASUxGgBB5m92FOTjigpDDCyJ0TtkOJ0BrPo+zzEkt/fR+junph/A4bLS5nCD4g3U0/
6odqalB/MxfdGXkXVxYMThgGSREIVoyli3/ApWI+JyP0R8D4qfuajbc+rvrIy6oYv1zKdwzIQOzg
Lrknyz6S6KPn0GKnit1mEgXy57EVHCYfUxAHgvqxHCUdPDHmlSLn7PP0sJFE5XRlKz0IIyzTfzHf
qqgKNs1L9wjj9gYOnVFLRiCZKyCNC2RoBPzdkZXyKM1VFevKwKzJhFvpbe4lpERJuv+RijSnSWMh
x9f9kZ41LmAskk5uGbaVAYwDXC0YvHNcC4Y6kwDvQDI34D5nbdL6ezBWFOww+0JKIXgUCjmNhZiQ
I2vmPbiaNb1npX0seJakKjNvoZ2U07txLFQHCKXghKJ2uR2KnJwIntaUA7BZMvgbm3CUOVAfYT0E
/IyWdtwjbCEs0mj4V4x6+iMtkUVRG7F5IdxvHJ133iWlR+oTcPeaLXTA8L648cHIeFG+uSdRk8mN
fqOna0LUEvrRPf7FPKBrIdmNpLjdL1mEjiUvBu6hlUJg+7JrqxoVt9EdqWmEGaZhCWiTW2a7sagl
IPqJ0zRmUcKqlewiHGP/vY1IgH3jB1VUfTg+BqC+pwegjgJpZyxHvMNoy73DMRqvpCoeVBRRG611
ouSx4lLOk7oqCBzgWjRobjtQtMN6PymQmAcuD9EZgdY3p90zXuER7JEYpvE1W94VNC/hZQXDpntf
dM/b/K/NrvErt4m05WF7PL2W0teHriZRrCmivdl3nyLDWtUqKvJNhT0ijUORqheWkbljf9hOA/g8
vB3zGMiXO8VloqC4tDf5ooHW0U9PJ/HyOkK++5O+feTEi9rVzuvoUlIhZhpFlbdS64sW3RhZMBiW
NTeVjWg2XeJWsqebcVKRCnSs3OljST3jS2i1JqX3GXBpey+TnkRf3a0f9yimokhCbLEcz4JMH1xs
Pa0sEtGaE5TDTKIcGLsuG/lqKaB9pijuDz0t8QtdE/Gpq+RDn7ArdqomoZaelLRsflrgUtHKJqw2
HFxEOcCGmTOG80rUA1hGy3uhbaM7RpVtykbLmfH5B7QgVG2qSG+7o7atjh7juIIquyr4HJ1BdZI3
/e4jTWZThtMdjMyzn3XFxuq5a47rHSOrDA9it/Ygw/RoEPdXRzWhHQiEUHXiMACdSijZQ9VhTOXW
qBb9LDNEi8MJH66MEu/7JuQgpoEw6WvnH9nUWB7Zm2pGifo7/m2z51JgAHFuCcnlNGdsqzhA7aza
i2b6983EsypbRUGBAbqxCPr7vLr6KUqQiE3g/gXELR0RNT3Uu4zl3es5pT8qXef3AJP15ol2FP0z
N7qoljBaosFe6MeTXPzasd3mCHkhk+R2MhnnZqT17PHjtLYxQiEhddiPzgu2q9Q7qgyaxERwa3BY
KoS0Q3ZW1nnRz0EAAcyJSBGb5ESi6Z+GJPnRDjsn3Z2N0GTmBQF944d6e5KG8sK5IXd8GvkP/I60
8PXufz6UP6mUfvzj7uVuUYmqucfcB/UTwX/nGeS74+L4EmUd9TjcMdwe801vKN2pAEiR8StwZds4
5JG6ruXO92FBgt8eM47eUPzuFmWRb9xiWckNCJs5QPGmtYcDqEUZJ1nimb0Wa22Cezv7wAkbMHoN
bg6SHI0/QobVWnDPQlkNUw6PwFRp8DJZwYHe+CQYCcvu1gFdEfdxgiPFMa119BRdEkxNGIumKc3f
bbsfDmlGR+4IR3YRkSrUwMFYHR2UUF1NanGQmsA2vnMX/pP3vPmw2a5a+CRIWKTQ4dV/HKLxrmqB
sIu5yz10DxCxSYTMM4YyKEE1Ag6cr7p8Sq3npLXdgvqDT7/mOPCxeFOCORvTZYYOHyXdcavgiftG
YpzCaVMDzZhJmOZZWgw2Yrmofl6RVGKkvM1f6zT6GGsf9+mGVk0SVX6ZQpue+fMpqSJDfJ0Cicii
+7YPJXWMikxLTmxqDL4ktALRWQYlhQkrKB8P4njyVwopDqr6AgCrl4X8oItK/hLKUAl4p8siNfpw
k/ltaZUyT7ppUYE9wGT7vacs+wDMhQv0gkXKKG60T9YDeyEJ6CfkzcbwG/pHjihP3NB2oJSEyRv2
+CPplrA7OgTDuKHP2/wM2X0Pf53n7iVibHZUp65fCzcCSnDWt+HWtWi79nUDqjkbKu76RZM0QgRo
lxNiChBvVY9xfJQyzoar0W6dEu25Tq2driL05qshFDzw2osjuXuyH1jAB8QJKuQ50M+h2KpxjUkT
0eQ3oz9/kBOU5r5/wP8sF0OYAgAfdhO1E+pRHlmVonawVlBL7CmOnCz6+2Uayh8lY45cMSsbgH8W
jjPjxCl7Q9GJXeg1c39j5wqttVDsKuDtqDw8mr8PU7wJ/DweUU83CDpnBkOjyznAZPBznMPNLmua
LFikHcQLofzKgiy4NfvS511KA5XLtudPqyxi4UFOsY9t5FL7dMRBbTLsO4OwN49LlZNtI8lEv58k
Hqi9uuEuQsTYwzTwHYiLTGwQpvctFERX8vWMERbXyBC3oBaMlhiLq2+vlkhBJRDKYr2encb5Nn8n
jZL8g/GFW55qaMWlD93mk7baLAwiTXURmKOMJeiiyc/QUP0Cze20VWg8/NdODm9EW6F2JgqrEYge
RUCIt2UrTQwvinPV3YifAreV2xFEYikxef7ZM7K7sYP46HKkcpN6fQjFXAq8yzq7QpsFSRVkaJlW
aRsFPWJgr6xcdhKIZ7/1xocgTiluXorR7w56hFouk+pqQKOsp+dBNkRz18FEIhT8R+zZgVNvlHgc
SAhrFZ8TMlr0en39twcbK1+EjGLhwiIrJJyG81pPWQCrxMqp8HrjIz/fn7l4CySG0mNGjZf5o7Fe
SR5Z0FGEy8RvDEqie2WwCY7pO3qo55ibAZHTOr/al+iQwy25zpOq4lzYrkwgpdsfPBFflfRqzPk8
chWV/417kDXUrM16pBBAmqZ2MNtAT+cmZv0uQqhcVa4UqEpDxtEILoQ2aeQpoEf5AdiN0sG7jcsZ
YGFvzr8kIK3qY9cnxwGCqSfBaZNrzbZ68JHZa+6/uHiMsrm4qQiqx/q2Uk6uuM0DgEvseh2mTZWf
3c5+Z6RdgUc4LIFiLk0oYTpP66C/3UgR8JHrtpsJmZsZ7lPy7fQC4o5YCs9Lnk6bAklVLa2uKcA9
7ZJTjVEmKXGiOeJdG2MPOidiBXspUNfpUCZH51rInp9SAl8fFg5olRPf1voiYGQkM5WQYYDLndyu
s4zriDoe47VDJD8abYVgn5SQvmMtou+jbiYNU690xhpDKYAZ5HG8k2VGWM9/qNScZTU1ZBNje1TP
tYlDz2lAQL7x0JN+aJW6XtHkBmN6KXilx/xCfvy9cTY1lw/zHQcGy0Nl2Z4gi/aIQgpTpBRnDNw4
rNIuhSrb2YTrOumB3w8VWS9S48rBUtdNHfqgdrupCvSSAX3cxqKq8WYXuqHnNA/6LcPTJqOiYC51
GVNe+3IS3cYuMkgT1MTuMdvyHoAf0qHRWgpGzoTdKRt90n9j0Wi+DEYdDOk97iYXrnprwxZ4H8K6
Nk7Bzc8l8eDrBcqlUVvF5RgW+WXoTHNAALFK2bKdoTMJfk2bKOliERy4ntYwU2/meS6r3doe/hNR
FXnyKfR8xeNGORbDuZ/tJrCAmPSXana52eDY8hV/kNN9evQvLakoS4EY1uzerAxPApI+Y+7uLAEp
Kk+P+z14F3za83odoz6lFUP0NXxYwfcfmfoTNIi39JckO+iPQ0R4BKMsCL8km7xavvyuFwHvvgPQ
8DlJYDWfFzmt8cp6xkJ4HqxjUsoUSgjq2xrTLNiINhhSOvNI13lnW8Suhst+8VL4Jurcdm2U7xEa
0tZBwJtLPp8RFJi6LGCl5/rGAWp70qUhjUeetprdU/cNykkMVx8FqBgLHIIVg3gmXERvynLo8sV5
dUJL5nM3BYmKwrUfR6MHDxtSU4HYemAwAg6kIO2U9Cq42NmqNcHasXEQ+jSZUaxO65JN+rdxrG7o
jYn+en4a29SFmMIhl/8ngG6p+hkrYFfShysGQRS3IzIebasbfossOfwS77QjGHaW24DEUNrFbpWY
x0oc1dGC/vriwAEbsKcMGthMK5E+6DQlSPf7G9SpvtuAnf9qor7miUjvLOsCzpaFUUT7Aiz5xoVQ
RwHqA1lCU825Vibe3bC/e+ZXkE9OuRmIAYrOjUVK63aLhCG6OF1uAMqdjXMpqSx6A4KFj66ISUVG
yNfhkFr3tvo6vtl7bN/7aIS2XXbi9K4IskDkWfFE+nzuPwMW6LRyDqPfxvcMAMw0D40tZYfiE4Yz
CCuASy5ptpKDE6JhQVY8nCCFKP37TRaxNd3D6qJd5ZdW+fRzVh1grRFxbcbYR+a3+RrNX2Tk8Tl3
/VMm/hYdRwzusQBM/9eqTRuYDFSAZlV7JBRdCnnmnF1GwG1OLJxn4SjsS+3KMgTsjL9mXP5fH4qy
UVtUxar2EL0hwce/RKAWHqZk4PmftAcet0EmH8S37iMi5FoCZpeiNFGE+2bLConAvtjvzPWVJfAI
11rD6hU7UB+JaldSdYcvG6TItPJWoK9G/2Oi+NbTW787ual4rwwAcZkIBas4Sxo00LgD6CVHc+wC
61hHEdLeLif44O/VexNOd+gKAXqpDcakOEYS9deNdebXvZtGgghUw82BqBYNA35xpw8UvCgFvgxb
KYlqVooS909hsPYdRcp2y7Ope3KSDm/vm3B9oJcwrol1AGhO3hTSCUrac7mJBrMGJYr3R5htZGH8
nLzQx4BLL86HU7nQse6odSb/qL6D7NT7QVIfXsVjg3x1yv3pigkg6XnkCRzQC+Z0CozZQc3zMWHR
J6W84gaE5D8lb6Jj7Z6CdPj7J0n6vVQyVUeYBWYkSyVb3L/CBcyn74hFsR6+07/KftdI86AYS7ym
QcuxCQefDKyrIxzDX1vLmI5rCwyU0rH37aeXTbii9vWTy9+K55IIFFf2+B8K8NJGuSdB92qYVE0L
H0AFkQa/OCLzbzlQZuSKd1sQ/OiXTGyQAVxehKIv2nmI1PPBinKlzLFrYj1lkII4XzjF4BGN37sq
fBA6WKehEwLcRJC4/AGKcYTHbez5Pn7opMCUr6z+smb8CSKL0AmZsBJYS8w7iYbZ8kyBiIDAbrrJ
jnaTZ2iSauMcCxs9LYIViI8g4kJrB5PD3R0f7xom5sP+P8e/ozKeIjsvYgkuCTbN71HDpfGTEFMH
WNfu33YFcHJQMHFmWOkE1S7dntCw3YU0HKrNihC9dBU6Hm3xZPlFNLJ+rcyPiOm2A89UHHQmLd7v
SKZy5SqDaSwVhAZblsvOXg9xUQV58unNdpl8kbRF8ylyqcLYEyN7QU3P45s7at9PGKdhIkiCNya7
T9zMrx33pgpV4IFUx+NbBk22YnZdNEufFUd92OQuz3n+JWVMTGNmB2Nsl4WFrg8a3F6Yakmt9B70
lTvWRgvyGaRaQSKqrnUdIqvreY8/4p1iSAWyTA5gZPmv7XP2Wim0ducCLKIq+AO+yLZ2nw2BQNHb
x/LQMqhvW1BH7KX66KwsoWELAflaWb1HNSGjA7/gmIbhyLiQBj62TXa2z25Fh1WGOa6dJePUYKsM
m+hLfHF4Ay141mE6WqzM1ZW+zJLEEPlaoGaIsSSvty78iuhtvS01G+1bsnNKZLxlKxgNuVyOBgpD
nT3/GS4ZrXoqVtwgf2VDU9UvkyACZhstsGmOXakGxgeFUWjgfxGsqo+3XrxFJhzsYv8mpGP83tO5
ZIwBf+YKEQXh3tqMSidrpWl1bfsVKBeSWsdsum8Mjota2UPRGpkEsrPck9oajF3hrTADiwq2yE0G
DyHOtK0EpK6emYs2Y+ZQN6zcSWzRHUMY0gFoKfXN8IZ6r5cf+9VRUK69SrwI2Y/SW9FQ+G0BxKRw
pFbBkSlDKMqHKa6quZ3qbenJHqtpbkh9i8DGG9b8TdqKxQc/U+aVESlZHzXCEc0lTNnzMv1X6Jth
J/e1PNJu3unAaP4rbWY+oRBEGPt+69PFy5N/4LvE0/Ycvv6soeguY3x5uZc14OYQ+Xfq7p0xVS2k
9ZySl6iIerEG0SGCW+O3zZ416+EKGlNfM9JsyTu1TRjSQgzQj06VURMf8ecL7uRmd2xuTCGqL2Yv
i3Fscdg2aJImfZc8YqqHplXsb3si3EA/IeCYsfhkFWq3Sgd7HYE1/V9dp1NUzNWga41lxyJxR3oD
O8WM0tDImIO/TmImhRbvQepFkkh/M/uMch3kJQreMFCAEfiY9sjg8/lA/UV8B0KcXVuBijzUMKjj
ghotFoOvaaac6Nmnj/9/1M+0T+lQQAjn8/yk77nSkankyk6JB6RpTJJEMMYGGc70KvyQ5yRWJktp
sonHeHp8NMoEaupX8n6Ot0pSwn73FRcBSqlE84MmcT4pMK6EUtxGrHrmwV3Fe7OFrPizbajt8gAM
DfAeo85QZkUnF/f/eyubtqSJgYNoaFWb2GoSbAugRi06e677DkHsU6gndabeONwETBUnhw2EWHRX
45+yBkGibKPBeX2jHi4aeKxdncqlWEENKI9leBO0xMDXz2basL0SPpn2cRJPPDlaB8J5AmNA+ncu
bj47Jok7bU2nCzk5qpOzney7fLAnYX1RQrpOBBd0DAUXpMnB7WNimIrUfJWUwWKXEnDvT0Mlrh1t
ADpSXs9ckT++7/LKhstkkl4jZXoDzT94HdopISAVLav5oGWhQJZs02OgByb9qxnqUxP4VBcYc8qE
gB496r3fW5lcCO46umYpBwL7HVEQcHg1HIT0SIydNwt3rBVPxuyVviTOHOSVkUOg5UpAMw4PNxHA
hK0z1YPfbiFT1eVG8EDblbELLE0CpezLvWqhiKO3odTgZI89uNaTEGEPK4Bb/1JD93ITo+da077/
YPqzbiwrazV4quSR+MlEt4cC2G46bC2cgNdl9pzp7XUVAAQLDezKrjJOaMxKty+AWf5rozMvu5FP
yyNgvJadSJPCBmIuygm01Zlj6eHYUaaqIcztTN0VG8jS/PkhIZYoFTK707HTwGs768G10ielDvtz
K89gnNypu8fhAefRR8g/b7WFP8In13KGRKOBo6EOc1P6RF6p95NEcMwyB2LqVyyFLYF1l5wM/CYf
SwdLVr+oLEzmaXWeQaoI28SA9p8my7QMQr8HD+wiFkgQAEROzIQyi9icnO856kjZnnVghQOf2flK
OHQ7XGyHx9ZcZ7EiA2Mcftsyu0NzitusvrjvP6gQTQ2rMSrcQjiNDQS5NqVafUhbUocZbwJt1zWy
VsKT2Odp5pf0PkF7H3HA8JN3EcJef4RnDJII2yP58CK8DC1dEwAtdQMGNThDaGGC9Vwhnx4JYJ0g
5uQKY/Nd3fos7rWih4hNTWb6PapQGLsffdLUUh104TjAQ2JIBb6p34yJVUliIGkUJBDPVAzgfYKs
g5X1kGqvbFo2Bx3IicstA9dboUyT926lSijECyRTKRk9XjEgaeVVs8fpyvbdH5XmOMlKHkKDDAk9
L7utYCs3cGdzbpcTETD9sr+CRsYL2q4ibJ3mLHuh/0YuLDX+msOoJmt0cw6ntm6BX92/1IwNTnTM
M3yw4nwFv399c5MKcCz2u3dVQbtzkbylWRQlBPdfxkkgfhZXSfP0iNfDkwtlIC6/sjGeyptBIQ8m
/s/zKYuxwq6zkGWAuE4o2gs4KVpEcQU9EA728iWn3TZh8soBev9fU5qUBwdQgSTY1Q6VagoieQMy
KU5fOIm1iydUWXYyDhr7t/eROkw7D023hmyPyzJ9wzT1Uzai8LGzuTc59cmKRBgteBMKo15ExpAe
58cAJg9kahWNA8lQwNoPfT9cyYU5m+hoTY3ulZC7HRiB3H8LQejuUHcfHtUBxzhnRiXYY5sTNx3A
UxMDYiTZQAHN9llFloNoU+LUfVCgH5hLBmQ1aWOC19L8DyK0J4dBaDVbD+ikQR7Hk1S/NQqvzRIk
f8pw9cWVm+PBBaEExzJhDShGFMELKrGsz1VGJVXWEtB289JgpLqW5rfbiQPqIBll5QLd3zuJyAoU
+PpcIeTC1XrbDi7AHD3LR8dLWti90FzymWwYJj+ZYYAiXeUY7OAH1SEwdhpPpKHpm+YzTA8YFP4R
qraDveeMcYt6Trusu7G2pkHp7e94htUhrbDzrS8higI7uTCh/p/Yd6EGjiPlUe2e1MC9EDHZyVR8
RUGQw4bAryVGBThrOqX5522ClYyqdMeEV0KLeVN1t2WcdMbv1H5eJDs0BsaYpsfPaHevUdY8KeFH
O5QkPzjyo/CWSKmU/t8Ezysq/JVxPhLMCF8rj+ATUr6azL55gahhEmVUSF2/75Lq1eDzEXjtn5lV
gDOMJ+/6oMqBQo5cFtMs9uvu4RT9IM4hvBTou8sdd/AWIVcrwNKt03oepeGhuOWR6wcvA0g19ql7
MSOOnahyW9YGDfp9JIG9HpXxsBB7UGGSaIht0L7m+Adzv/1zkhFbUXnouolo+GG0S1jXVtdSohde
nTvdCGFZ5Yq0ombSgTyWtbio7VE0u/sx+lBBfQGkf9UkX5v5pqdTly47ZgG40uYo5s4ERfiPuGSz
rIghudjqa0nOWc7ywE+khoXfadBO3FdhZEauhViWWZUdgCH6zmh4C4D5yAKmq99TkzX9gZioR84u
fC1P8WcCCokh2haJhyvzrCyNKqopIYoV9WKoUSdKLKSOdvunjJS+J8SFCCHFEGK8JNPso38APjht
cJJEKuiy6Hmrj2VHJkQJhsYvpicWOd+dLZBRgImLdnwiFvZyedFxx0vF3rXmMnk5DdISycHShYr4
kIPh3YWP0xGz/ae5QY9cna0bOFLe5QMe6xMIIQudn4v3cRzGUU00TMRoU4K0mDbNdzS7o2UTtqtP
GOiJzZQ4xuQQYPFlJuvQBiNmEKJgK92L/7n/8bHIvDQz4txqYaCPzxysblqmAoBf6DKVDNXoOtZP
jlZneVvsoqAKwFM3Ni98ZolHJ4bmZD5ktz3yI8Coyp6lePgct3zNxro4o9YpecB82jcO9euiVwEp
968t5cCcQOWoJPJH0+Wjtv3O1PYwcuEBKPpFoIfLreiWgZr1A9gUHz3dPnumTjjIBWVbXfin2KNj
LgKXV1INDdB2q4vST4t757AY3/iPxkSlEifzcL9BmOgFN8lyPhG+CmFELLmSrHZVfLK/ocOgAvoD
SwemobJ80yiwyO787L8orqfEOMg9sgkIWgiUuvBP9CMVt/7jHOv5QyxmUOT7IbSuHPA4zW6l1KxW
wkm/olbwVEVFoUCOvjwiHRG7m/tgOanriTFE7NhW9SJhAjls3DVCbHaLhSNfaKBhR6L44wYpwxt6
iK6EUxA8wky3TMImvsgkVTd/XzeT7zkgS3hUOM60Lhn4lPuDiFTR2J1Gwm8B/tKnfk6B+aogZsm1
IkNnIqmYKNk8Y79uqOXBFE2lQ8YxCB/6ehS2RYWdJf7VBv8tuOwQAN8PIeMiN8QXJ94AddGjePXt
Z2xW4jwajlTunixOaIVpC74CGPTik9pgT+Hqu9Ek5JgRRoTb1d7IUsiVdC6L2iilH5qqigmI3nrI
C2YYDZ2bcR0mHLNIa/XHKR7ixfBIbZUc4hV3Y/4GPJv5/sjS/KoTUAoN06y2/yWik6lh0BQ76hjT
FbiSTG4qkKOF+7+gTFWkgpDB/6wH8uWhQdYxJ8V8lS75sVB1JYAb10mKjaRjbw4j4XTnCzm+ZwHx
sXD/p7xrlQ5ISoY2tvzUF4XOwZ2MUBaotXoRegJ7gz5LDtx1KYYYprsJv5AFznTGP34GuqrbzTic
1pmNIiH9TPC1ihJPPgkRU6NR70uK7Mwq7A+I0DUoL05caE4e8Bzcl4Rx9hSLY6+pHnlF54c6cOHI
bURWHXSY/GDobhiRXSKOvqAS1CsZRFdddFKLz6DqoH+rzXCseWZ57wAWQakR8i4ZzQJ8HNv5C6QL
FYVqSPPfeyzyr9mT5GEoKOynYT7wINiPzuhqIDaIR0wwCG1lIeYyjcA7w2iHBR1JwcB9Y7ycf0EW
49dYLoz/I2y4JdRzfogpeBgt8QxCtXSnxI78yrXGpfpf3W70PMc8dhzuwS6jmqbQ0YMxUv/ftEFz
kcSht9er7eQGEdMzgc9SbyxVuw54nTKeFWStF1Rph2sIynb9Nt9iBS6xIHODMVK8XXQ3U/Q/4+p3
UrdDujoWd9owsaK+BVpTAdwXjk0hjbJ5N4JPL5pz9TUTTBDYhxiPY9QGykprsd8Ucc6dvqVlR2Iu
P0221xndgNZz4VAHsuMvjixWeGM1+6KpTj4xd9CsJoxqQrfzt2gIVGP4J0TriX4Anbv2JGaLE46C
a6qNJ9yeterF7ZbfqwKAfTMNCQF7LTq+AlVNcgM64TfmvJqDK76rDAW16mT/SNCWvVQ3lTLF+7y5
UoczwTUUzHFlUZYvDsH/m4wWF6vTG+JIcLBM9wrk6pFUgkzpRoxZUPAE71hhanovtRmiU2n/sC5e
QmdDEqgpnAl3VoRdvEXtXlNZyoY0Dr3tcsamG06ZydJp+KVvRtWAkw9mUskPLO+bin/IaV6PaKc7
CwARVB2jrhM5KOLh79kqZckw5wb62F14218MpHyEr6WwE3kzIm5z0lNRGqAwlVoqa7LyFmZ8Z5LF
oOc0LVw+ucK1iNeAwjiFfau1qIapNTGQJzWjqw//Xf2FaZPs88wCsZrec7NmJrD3fvzr43Xc9dEz
B4JdCQz+ZwWFrb2ZGSmQ57xC/l96mkdv3CU9kJSuwxpkyctDQjuqSzNOXiRSRDR0P0rgB+rZImAo
qpiWTjAW+IjKHTs0W8cpGmUEMPRC3sgwH4YidJf9anVIde0Mbvg2Kn83n8Q5+3JoemrmGwxccm2c
2oqTavqrfs9glDTz/tHfJPVs/NzutVI+UsLaj+IV1JUZk56UJQ92NOiulIHxvhx+1KcLKWp98ra5
GmhQGxkc0+T/QAQZTJ+eucsC0hCaSNwn2qSjMAqR2JNTqhD6/lodLJC3jIU2JRgCzbVTg8pyqm/o
P6xqyq0v302jq2jPfmz3ZrqYKXdn7XTMDqc9eLDVK2etPx3VLmBwit8VWGPmYu+v4Q/BBxBvIcqm
OUXZn81bOghYZH0TIGmOR+H0F97DkdIY4hkcq7OCmDSi3FBYnSRwcAli7hSkMmx2RuXhYa81MClP
erYXvi2OECCCMZ8JLtCavxq7gpa5shMeTy+PHghJcd6H/F/gcDbJQcLvD/TbSu88/UPJjfJJRNwF
PPDA7PMuRpTexavGNlJ5sHYe9KM9/Yx6QFbwK+CSM+1mEwgoGAYa0N+wxQzdtuwJYFkDmpEkO1Df
64woBi5L8V4OzKn/TJbvlC5do6kuj71PnUnd0MdHEza8iFsRPSyVHaC06XBoTLpI9F3LsvleCrDd
ySBQO8PCNDynmfe7YUsmSAHtInxFVaYl/eMiBGDGw7+j3IfnUzsCy5uamqIIqe9s/LdPhKFTai2H
UfQi6V4N1j5vzVolQ0+j9ERYTD+P8FB0y/6wC2NUafLzeg2Nqb7I9c+YsR7I4sAqZgNMlgKIH3dZ
3jGpnocpkPwtG78ONJgqSyoI+kOrHSMe64XBbw/cBqMuu0g/FMXIpHqmfT44xl4EGc52LplZO/uV
W7S8+2dzwfZDJa9cO2av4yiZVCwsmxTK5ZcwUIdbjDu8EfIlKtlkua6Hid03E/7GfX5K3iICtW9s
FQnjVt9tDSZVA3xWTKbgHGUryJfZY11PinViqzmA1zZSl2tmwNc8Oh/WPYCgLFsicXL8Y1IwKgyg
jJTSXFbvmDpJrsmuOvhx2DP0/21+7JhJsH8dq9xyxCDq3N0j746b/x90S20qJhcyEuOkDBW5aOEz
9FqIf7GeL1a7tGeZA87RoUEkr/NuLMqV7AmmBF7fiuF8239H0lFZ4uTVz/wgTAwYf/W5A/RGWpP0
xNeOH+6j5yQDQnc3JY17aalhUWFoxTGYn/QjLqVenHd4+xa1aQ1SwdgXUq1dRZLBvKr0D+/JN/vo
FzxQA359YyaHrz3xwzE2yabWh1wXkP5emLShmBYCLnGi0wl6fVfVCuX4/keqfN3Rz12pyvBCAYjD
EitLGzAbDmmJC06c69PJYll3/+sEntSVYEYMkW1b/CsUDMPmTl4GD3WNl7lyrZ4NKf4LBWSEUsR7
R5s7XiJL617xbmIh3yWhDE+5AzUO6riCmAUDFy89LS8pYggjGxSV5Vkh2wWKg7J111S6HEiIXIQ4
1IR47M2pqCfisqojkwDDatRUXrG/e8rv1JbxLVZlAxoh4aTTkLw1WRMTxKlKuIRhOdtzY9sg6u8g
dmRNDonIXoCS18QX997PUdRc6lVRCi4RIxNvAmpIV6FazIQyINpn6/CIS1fZxFT5kjrA115D029v
0/l99xH3wtDUCPnbKqvVhQkGQRSMuSYeI7iZetJP+CUn62oAQiIjofcHtoB6qXBL9tVO5Oo6HW1o
cWNG9FtVBmBJaukH4NrMIx+1PfAH3mgO3z3SedzDWpHVkCFNWMs19efQejDzDK/QDn+NI+XhM3Tk
dpEtX5PqRSjwU1VJbI25O6P5XOqpBdWQfK7f6DnOKL42k1gw/vzPtssGNJpoFJIVK4frkIouomwy
LrUAdBhIvrS5ub3kdDBb4t8nTQxdMygui/qxMLthp7GNvU9qB+wMOsd9cMrmuKuG1eAApA8ZOWmf
WYwvXZK+xTIiw2vgVKoasURMs0Qe3b4BJ0Xff2Z2BD9L5sB9asU9xrFbGbvrmPYf9dMFQhK9V1uW
wG9zdWG+kvbOS4k6D1xT9lV9fSB7Tj2XkTxlK2NN2jc+PFFvbgsjemFHocRJmFQIvJ8b1342TQ0D
aj2FJbWHuIDTpxxPS+/EPnlXi4/pkK9VM8rXPtkTrM+H0r9epJLI8NrwckuLZMyyaYSlgnusg1C9
X4ueKsIkP0kUS8dC4CADpq7CriFeYnPaoGVSPx3+SlOa0CW6/V7BYZrLu6XMDx1+vHU6UE/n2+p/
KDQGpOuSvnaP0RKXqxu+LMxENNNapBkeYKXow0VusZinWFXHflI7HvT9c0TqcwYRSW8c5AL22Q3w
JE5zi3nJvBsFC5ynjKPY1VvMfPRykL7YLh/sh48BttB7R1ZvyINze1qrRUnq6F60luPcUJ87nrq9
XnhCj3zF0Rh6vKoR4hKCpfi1b6Z78d17RGAYr1QKGSWQJ7lZLh9XmAoTYsTJEpssggXOU3KdD2cr
ruGNrENgSsa82JPlctl61xv2ycfvcserRHES4HJMeiHNlMPVy4fw+i8vxfInaGcOhwedyVMnUE+/
GdVQVJc6mk3AyTQLOUf1gT/EI/a3EVN1F9jDy035ptSuIDKUySka39NXBWu9izu3iQoSqCzSWCiY
ohR9Xx0qxOmsrjiP/vInMwdL+aHxPQWPGLnJBz1vVFlA2vdffZzPLeN4wtTcLO6ABi6pkv9BlhGN
C+mBtivxhpZYck5R+oE9BBQvuPy1eJ9MGjr2PiKaRY+Aue7zhzQIDaYoesyWx5CTFLQNoWg/Jy+n
zGxuSHh6SW2tUc1UtSwDHxjzRzPz8S60Cmh3yy4ZEPrT8uKP3BnIZJqpGahHamDv1MnfPLb5OmJv
dW3T3UAABN2/hqzJyH0CIme96ICDoBf+M3tdMV+MAjscY9aUTkoQfCqofQj7IxuLIzomis1YSlGS
42DJa270k5SySM82bV3Ni9NXCAa3p/pWVhA/sa8FYNgrswz+elYLEg6A76ocmi78s32SaGHZVezg
v1mVB2jUx2YY6i6nVh2rDFVzMjQBGS0N/5PdvuxAd4iuv1/exqDbROXukqqqkO2ZdxyLzAyFvTuS
4lAWv8fQiZZ9cgI5wY1HQZPDAzjqxqN3NQHWVQGrJTCPFW25olxZpqBN/D9bCOJwolJOH6M5S2b/
z2ndUiDpBTlEfyuL/TfbeZWPCzG7eMMGroNaJgYpG4oVCdMF1/8mgQww0FaEf5yxIC28GcCJUCTu
Q+TNxvF2nfIDzs7o6fDXLk2VZK9d/URBhCfrV8+HHzL2PuwsRi88IfOr2mF4rj64uAUVhGnyJuew
Tu+xK/tbR9YPp95owOtNVNNMEcjXIZRUzrIJ/qUvt+9Utz9rdc92MJZOfGaL46AU8r1lWlUCn06n
4JVNxWA1aL1Nad31Bn6t3hI26vi9s5hHqGfz+6uT8XqfR+bndFDNyhJlXNgTHV6NQcM1jS+OpcLW
ZXZXc1bwwF873baWNyL4S+YvalKbrO3Bx4u+obt5Gb7cfaNUpdZAocxCdJkuFH3+Zv4JOJnzxr8a
3wtKn1IhdnxqnnZywHEQWH/zLvOye0CjD8ebPyci4mSkxh7JU5JloAbrvEsWeRGgONHOWbYettFU
h0cmAfxKjZBcd6bneICpps5U6RdlZAWK4wSo44CTEVEgECSJQDnCW1QE1kP+j0g8CIcnn+WMnPxY
nJp45lioUXxtTb0bMHTab7QDVeNYqOtSSHCRjkMvE7mwwwUNbO9lXeJZZErdz8Xbwfx6p8mHz5EI
Owxy6BQ021CKkCxPogQ8tN077hEzcCahgtzJdq5NT5AEz/UxN8Ac9e97DITnDm63nUFcm5cLOYjn
HARj+HX2w61Ytq0tU7Fa3B7Ewd3JVy/eANllzUQ0G+WkLKIZUVf3oYKlez/hn7rTAG0S8X1tfrOB
ISAWOdMvozV1BMMTgCpK9fZ1s3hB3q7XfoUuVOPYpZ57QVxX89IFD9qjeSJKHH8lt4p/vo1vp5ey
o+yGOkgC2quv6fEXjC3wlqG9jhe6HnqyToZoTHPeDESHaLl2+usMuQPHyv9812/Nn0MID9vcjzBj
55hXiauhzoW6DAtdzEXeNG/9Xi8Y+IIQxX8SqeZLSNo9VVkt/DS6QaYuOzO/HV+ZHwyROffUj0OG
3qJ9Hv0xvkQ2XSj9IRLSOnzGsLQ9UYa9xcey8C+MvAnpcfgkFZ+RY23lYZ/XY3OoNGOEnwIeyNLy
fU8jS/qhSHSsh0kqjnFb5bUMgbg8ZwdIPgcFPcYc+xhaoVkTlqwlNXMNqAnM6TIoSfsm6SPIKtlt
VTA45U+AVYVkPxUINLYm1VBQnY5qgc/PkGZsq81kYvKkTf677DxPbWVxyueSno7F2jsNy3/UVJLQ
RxGNFyBXkT8Sfuy4OFpy6OPopHDDVkXERi6BVoYRBD2bnQUZRRBYPLRvkx2pvLLroRQk+5qEKONQ
UGYbuuEmEDG1NE8dC/Sx/A5y8j8ewuukndTI2iDKQ4n2fVJL++MUtj0am5p+N6KX8YJ0dMRkuTBN
udg1R1Ia+I6GsyZAN9N/rjyJsHNHqAwXmKkZRHnWxNkuQAKIrLJUracllkXQh7aSnzVdojTqKT6i
kWE8LTWeH+o4Mr5RDmlWb/j+fE7hEtGd3eY3+VA/E/8xbFpdKhZMVobSkxdK5ZgklueVo2V4ejlM
QVO/sUrjWT6tyiswOCUim534YvcLAF9fe79Y59aZwsbcdACUyewdfv0g8ZAuj2G61ZaJsIAuav/B
btSCuO1aIGfSH/PrMBPAKDuanZ678+NedZtDuYx+CSEfxylc3PIsm5QWZYbNsJInmYDXFRkhktyC
1+uzWTTF0KyqW1PZrAZT0lnFXKG5XStVcRxWg5QziAbhmGp1nUawfQ/X5Jn9ifvqV6KXLcVh9M3o
hYYLJPtfN6hLlDzYQLMTXbP9MMsKDi9xFd0VrUsm2bES/8ZUe3alwovxDcy7jFeggb5EKqZpltPF
sSqj9glHhLEhN+PYZXC62PvhexWaewXbKJ9f8fePacNHX+s7GGhkdm7hG11KBEbmlE636/4zlIiZ
GTRjJHdW23BjagNCy3KU+SKzsD5e3MZ8bDyMEPqAzIZMyhc1G8Prb/JIYH8aI6WSTD8+hmz5WPn+
AGi22Kts3jF25acdpU+UXFAox8r9jLfLaCjLtOyr8LLuDP6mqZCw6VE8zUtOs3Z28bIud5XGeUpD
gAAapm0E9j3weiJzTtwC2w+DXHu1BjfUWw3BFl4kg40bIVdWAf/VBnodNNE9o/lGr9tNuRO6nWPC
ETu5Sa7QG+7KQrNYt8/O0dpcAQ5FeZUHDkzUBTb8mYiozxR19HEWvW07jyWwXySmZMhAPE6ny+FG
yNEE/4VpyEjCINXYN/5GIIvXOpMDGPexfnfKhwje2m4EUdas/amYKoVFgviRBR9Xtcmiod0n2nT+
JIU58E2727L2Cob0nJ19NSi0wpVTe7Qj4+KMt+EX8WsasGUfvWX9xRGl8s9K8AWGcQZwM4O++DVH
LvI8sMadZg7kNd2KzgZntBPKm/fyfYTMDjo7k5tn5YsIdvO26itQCTuOFtOAZYIpe5zupPj39RVM
pVgPOezoLeCo0e3DQho8ipf74EIDODJD49tsT1Ys6t89YlSQgH5KdeWw3DiqHjlQQ6b4EYRukrzb
0chwMJL1A9+6ZLhy3u7rOivFHOTa0Ty9hUknXV5tQtpjivYeQhu/qOIDAa/rIUOhBlgJAAf44/+g
Ghtx4QQazSMsO4tWfCI8H45yClOfmivf/Xc8oIwJadobSjcxvQY6EW9SqrBwKRaedyx+iKX+EKyZ
J32UCf8LPlSwrbIlp29w5gxeDA9ESpp+uRHoUSCP3Kzg1zuaEJVH5DBGSM1qxx5b05ALo2rMzWih
hXVa+51/0QP8dMQ0dtCjw8d0uDzlyljChNNYi+uRDCwXvYxrWZ8rEqryWjO/K72yib/yvJ9FlInO
log5jsXzcFnEco02I0bwTmDTJw1uS3G2E/tTONj/hsrcw6mwvYrEwccgx+64cCkBbZOo+gwD928n
6HVD5unxKT4AWhNxaSmYnxK2U2Y1rDEV6iZxVXVrxIVUc5GdsYOzfRlr3/5nEs9Aym6bnTEVKDDR
lmKYAeESZCN8TbGextU6p1B7pCEEbxg6Aaq5OyRWnxZlRaxGDejxTwLeRmfB8Go/0JvrR7z+ODDt
F+qgfeptqO6NHQuUaB0S445evRunm9cY7QmAI44ao7WYThjrUdwepXehKmyblTKJY6Htwef1jUzs
RyHYcTXRDtsz7jsLLG/16e7Qbl5SFvWYIo/OOpeZsoYpJtQ7xkigEe930o3EhkuJlYMrFl9Cm1HK
ovpD8/vCYWZcA+Mc89Lhc+QH0wnBd0+gLGS8PjJ7tNSUCtGxYKDw3XZYjxaSARfjFj3q4dJ622CR
2ZSNVLgEhs5NNzkxV6RaFBpMRM376Rqq9p5y57MjGnzv6dWP47/K5MI1iJMwc/JpYsAYQTv01BME
CRVKt/XsG0v+gm3jvcSmMVsDgzCE8w/gdwDbZTmpdQfI7zvs0tzMobeJKJyhrI1o5J7O/eYvZLcD
DXX/G4vAvrVzSr9yWVPGoC+cMkNnZLmZreuu2G09cR/w+4eq19xllKYvZ7WGgYASkHsCRjZue/IM
q86+7EvxSiUuNbZsPFLDC02CI1EYtwma8b9vmZrREA1iLaIpS2G4Q+uvSSX5o8OhLOOKNO5dcdhX
jbgohK9Am0eH8njQkQ3vTYeA1RQWbynujTu3IyTQqj4aon2jgpR4PWlwiBIATtI+cCGFiTs0gjqK
l5ggwFW5iiF4wclY7dDKVrhqql3mo61hUdglf9K2wY20rrFXjMMHAJrdduSAbdsaEYg6+JfKVhnl
i0mAp3PDN/NceX0mgc/5T4RHwItPJ9n0VMGAEK3tfAXNnQUlJVn3DvggfCdfd7UDtSvixv/NfE8D
z1ukap6Ocb3OotK+1Alhv7jTpRIlCVjSRcuxAIoDlsiKeyl048q3NxIygQ/gpJX40MyosXFLOKQe
pCMf2iX+5YgN79MZrPiwoK6rERK4cKGYXwGXM+pF57UZ5NUYFHlEgVIJYddabh3KdbWDP2vjMdIw
AoV1QWIzSqX4hhKrJAgZfb7g2VbjtN3R8dlKjnca+8dCtykb4qP/yH3MvcnuN0ttby2hDXIzO6cR
fS4B1+MY4jfM/fIaq95EowfSjPtImIht82UY6YXd4c/OMBVrSfUzNQ4kSWeP9nEssP/CfazBlJlh
9iqJOrAlbY3oDGIIl2IRURYGyh2g0vjQkPBAIYn2jJJjCS6asjOyKTCMNHEtK246ayUSJsmIuKmx
SzEZHr3jgs5cX4SLqwwOe7F4r3MZR70alhYduZaO8p6PIseocVUAJfKZ2NDIqUibueD36FNH8SZa
slWurGp9kadOMJwe+69Ho1i3+iGcdv/1s+7Fp2ZFzgV8ORb5GvlP0hH+ksq8vXujoLhmL+F3fCEt
ylNmd5u1bhmgE27qFNNHPBlyJlQhyVu8twNfmPVFvJBxaI3fckIz4wvtrlvBeUaySq6aIGBt/k9+
WjzkoYQe06Q8xZC16oWTxoRqEOSMnwqwA3REVEvlfqNWnKaKtZTcOzqS+H8H4enO29ah2TpCunLt
8mlytxky9b5CbizQTV6w9sgOkGmXSI07T4YGlha2Vo2yjbiwDbbPL750hoE6e2P7V+gRxEngRZ20
aDIJ2YalhG+p2mAT7ckvIcbmGrhz6NKy8lFXFBVzKebfq2jCISGTnps8vXPDc7EOXINrOMykeO+l
0aVa1nEw4y+U6v5gMr5ISi07rgHl9ccqKbH1MsAQNS18ted8ZBV2KnXgAdoJ/22Mvez8KG1dvXnC
pAIV3gzbTNgDuQypAvb7vfl5MA2UeKHGyG7Fl/LAxKN0QCDOhpNMgFf8u6uE/BSwvNSQ1ynG3fbW
ZHueIXkdcwAibFkLfqyPOve+sccrADi6wj14Xy7oblBk5yvT1Je4PX0rnYj3UYfMgjU9eDlhQiqS
Pj6QeMhLNJO05w1EAzP1D+oRMQ2TmF+SEog2I8b6BQkfjqF9o+v9pMSDsmfCCESvz+zWXzjIfv9C
xP0z3IOUGj2OA12Sz3ZTUXaVVqvGxzLfo/rWxuyA4WFTF+oDNfpkHDxuCaLVomUYtYUFuYj9lqSo
CosRqHx9aUAJW8JTLlKgM6dUMP2aMgKEU/B/pxrx+ZTJwgrGJCnDXigHPGIh/RfUtaLQbekUoWvm
/T0koCUvvZWNU+cwjfeRxGGGb/kBAx+8VSLZivVxbIvK3uryxPWJO20zRXdJcWIE9/FFMeScf39+
WzZJ4VmcoX5OX+xzjNp2WlWz4v+pohdSWujt2LLCE08XztxoUD8LSTy2YAfYfWB7b2PWfY0/c9EA
NTZhF7+6FcvrmkEQCcqWEv1hLL/ORlsYlkaht038N0VSfT9AQFxPfN3DhAs2cY2M52Gh7uR5SvT+
3nVzWur+DOSCLRRF+rH19HK+RfEokiNSQvC+2K/NgqBT8Z5dKIolJnN5a6GEE7Dz/SIabiBMnJPZ
GjZ1lnEkWUqfjLyuZtmDJfvVyiD+paXff8D+WFMl5OvwtK2x8W2/aUytI09Z3wLx7uQC2D7DZigB
dSsNhYBuaV77CAzo/U2Zc+S6M+S6UG15uwGTkyDLSkKk4HreKhKsuNgvQcp2Ey5LzSGSMY6nbudu
Pa7vGUyFLBpoDS60LTUxrLbu+ZlFJaEMrdyZ47Vjzi81EPzFrqJ6dO/dfiljL+jha/O7FV2cV5bm
voeqSVl/+HC8w9Vl0+Wd/jzy55yKZKufaagnVPiLNq//uk0flwWcT046A8Da+DcjPMxFgIERs6NI
LJjU7hhr27caaCl401fBjMhSDfxf+wcUjfW+yO+BsTk2nnBZymgrK3ZRTmCEwXUSKZoTKMtKWEIc
9lYvXNmsG6L7hr6FTkjel7j5W+lpvPCjgGfoEcKbFIvWiJW/EkfXs+h18z3gDat2gPEr+QLtDNh7
/gvetp1RGc35TaEmIwlCmUXPM2K6hmuolHq7dsjqfsYmRWmZLAQaOWPj32nFygUa7YDEY6HFxKe1
6s4x5LwrRJiqkLFLa8ixJGKFdZzvCxXZgECu72HZvJc8mr8KcdsPGJiYxEl42W8QwVaI2VloHuDl
7kBcXsOnqMtpMpUnxCA4cQED2GAGrmra6BChJH9zSRMVsA/JsYs1VM+HBMF8zNGjzEPhTAAPWS/S
riboUAoPPjRY5v+0e8atRgW/+MM9q4Q99yzVEvYm2O/ZmljHxMhTmimgXWN3/tkDjQxmSjmvlbCR
5Yy7ssvaI0eP1vhwgOOz0tl1u80ka5F3AxId7w28hfXgQ83jHGgG8BgJDaAUFOp9u0LGYi6uoptU
/jOfE9qjKXeHRzinAW452CdVvDqu+wlp+wk3Ajo4ue+1opw0Z4QKyxs+WsEX+Oi1jjPxvV1zRDcW
lNaqR5fCETorqiaNODGJcM72AvPt28F6o8MKeNBPWVce1UuH9bJIH850P4PcdHk3pUobItrVQLhs
z9rSOrwwEOZd54yjO+q6U2SOw5NhHR0+7dm1itMElxNoCX7Kgq/q16YJT/IIS/HYP38K7gF0wf+l
uEMw+0SPlQ2OFpiRDKMe6KHxirkn82ra/W139jQXlmN1tpbq02i+UDUeuiCMSwenodrxy50yaMsi
+WRApWdnXNeZsnMlUSvMBNGk51bbKsT+CCWXNg6pv7gqSRBMYM+vTBmXa4LJGjMX415/ma2jt+4t
2rwXCSf7T0bz1MvWCjAoJkUwzlndkugM5jccKCTZYSBbXi+kZTLOOmeZBWJ20z0435lPXaHi/wQp
qeRFIhp44HMlFlk0bTTiZie4GpFM9Z6Hj9D9rQPZSFy3Q/qBJmztjYxxsEkbrRSgZ0ryRWSlc7pt
JqqmvXGIuPoKhZGjYnjMQMufSDpc6p7aU/QXl2SnwpgtXi5A/43/nXXIbT/aW4iV8zEpa1Z4hrx9
+rFyOzwjXc7d+i8AZcKVpN8O2RkOuSP1xswhC0xNwi8jmxJroTvUKqtRs25B6ccC7PdHt2NcaGzn
HL4Kd0aZC2d8BMGX58EtxRlkTcisgmesZ9VgF7Y9m45y4HX+ouYAOGH+7qxE6yvAmmR5byY6tscO
M/QCmMEpkYr5F7JmaiIu7hQsHUGk0j4nmnoayf1ipvIvQvTOtRr9tgKf91/YXRqOSgKSQrBj4mJD
rPY/QVmrFpZNBkx1/J8FMytuuUnLfl9WNwEFV1OsUh101CyQH9x/TxYfUj4zRe+WY116Z/waxyCk
r6QfMDoppntkBOgJGlwe1Dq6dMRHHjcO5vMro0sYHMNPnXkcbyVI+BugMQncS3NFVmRISokEV4ej
j5I2PQzR6R7JtHv8cCfYPcGSY1BjR4hW7fIJ4UJOblaDxsbPxqKzezseTwYtn5DD5hBJnsE691rI
x/frYQnQc2Zjqn4O2kdqXHZoF4dhclm2PNNBaQvUk5dSDd3hLNYW/jhPvj8XWdILZTIXr05WsFfq
e1kehcAZpVSC74mLqzP1pdm0N0qT0+yWHL511wWRbSnHpx4AZMojzI6wJQ6FsEfDHaz11laE4C1A
iHbHCIN6jiUSSnrrTiYECLESp3uJ8v7N4ZN5xwLgP3Rakkkc//BB/VARWQ8vMe+8t9caxdutAzMO
yHe7tGcA4MlUqutSuZyAr8dgMOpDVCTAazpSSfL7qGRzE6KSHc5ka8B5x4dSRYA0VEvsHcfsxcb/
YgI5a2MFtTzF3ie9LrSAIt0OozY32We9aPDVa1TEECzEOpDjK6PuT6GMWkfXT1KZPvfTMzDEcsii
uhSMwtjW+q+tE7jxtZvvcfjKcZo44MRl7QlbipaFoWiGynzBtc4QSSNmbSmivw0pMq6KK8Z+0hLi
LAOQniVDZuuPtCji+bvkg77QeTlOKXXvAIQoWTLalpePOeHNc8CDLHmXVLFdt+dqIreFspbj9j4A
arqBniHtDxpmUPXtHQ14UKuLFG5XMBhz1CEd46sDvi/l7mSI0ow7prfpg/x8vDThL6MSmwRDIkWc
wEei2qzN/zi4KfqFfGR+ZkN6BajmH0NvVtc83sTHqRErqwmyhnmKDRqPgmgdO8CaBX0fFmH0L+bu
Q3yl+/sZB+YnCuN1tSFk986IRCIQWy4RNY1LHlabyRELAESbUJpsEm+MXhfF8SXl8ZgRHt4xaJMO
BdbgGFiqcE/XjcddTsi9c2+whZNikLdNAUopTJEeb8usdsydFni0XCKuVE4IGhkXsXI/7rfufLtR
PQ2xlNewkKd22mT6QKPcRev+qgCpb5oM8H7ZD+UU1yU8UOOmrna0AawCOz2+gZmKamSZsURJT209
MufpglgSJ4qffi46CyghZ77Z7bF2NRk6M/guZWuwZh63uYkDsRfPi9Z8CztYp1J2aen+OpDO1Ype
mh566pjAB6o90wEaboBY/B9K4sHJZ+dW1pJh2hHcLStbSGZTqL/Im0xAo+c+H7VslqQqIlT9BeFG
4UzK0x8TWSOmF8h8VV7rsDbNeSF2tDtVs4DDURskSE10OABrdOXMcGfEerxD10E1qkPyNGN0eKHm
VHaRpSnr3yo1G+Tz5eI5M60OboW2MRpK91vRBhObS8z6ijAd0M0eBy6NOxMNqvKNlGwTCv+tQDip
PAEGuZB0vL+hmyNHP0EC/neUlH4/uwJKU+ZVtwyNqd0Bjv3Nu1GUpzhQ9tCyLap8rdhkV/SxJjDh
Z5RzKE2hfRmuTvoqV+qALCJXyInuVutiZfuBqoj8ntgbmSj1sMfmHAEGDn+bdRxEpZ1duQBDSMwl
3eoHztn5moyp95Oy/E5a7gSlOiJXo8HGYr0do42r92zINf14prS/kdp+4xYBteY1+dPMhoXW3MC+
SJ0OMM4UYUlVeySV7lo1ocoDwKkli5OSbUOg5dPFyfrpVFsKExtxv2yCE7gfNCHfqtSFIerpbx2b
lASJ240vx4HIk5u3eoyMSOO9PjJjZjR9459VDIQpqtAtqlQFZmCOTs0VA1lBpnZ/8q1Fy5ednnms
04sq2rFWMSYTseXlmjs6IpH9dU6qygRvBxqe0dCiMJpsMLG92eLvEfmtUBDgo4JJo8g4trtaWTJr
NKW+DSqIcApIUx6iinQaVy9OKcL6MbrehIrryJBveurDDhocOvNavvJACxFxBjciVPlCK9AahJox
+0FumRR1IqNdQQ93A/D2QjfVqS76dMUKZERDMbUoV7VP1UZryYzbG/mh/w/bRz4PWXepqfJubqw8
bQvSv3xZdKv6n+WfWwAqItxfFrO9zp2ChevaZqNZdvBhbE9+oBYpq4MQKisGACTsbutWo0YinUoi
XCW29XvgGcIgZ4LPWegruMAidoUM4NnYy//eePDpZM7Kucsa+SUpzPeVui9ck1hDc/oWLCsnnBzT
MzhY1lUUzVx7SFdFbuCVzvyKqgx4ie8FJh0hdQYOoqLlmGd3Q2Yx5MohC7axtpgOIFJqzf4tw/dD
I14xQhh10O+Fk8tTuA4b2c6sUxv2YJZNMB1gcTnOjRv93i3gZe07u8rXyUxLorKXWjcoNZFgnQMS
f+p4Ml4R4wWqGbrx36AiBlgCQ7PqZcAswgEgx7RBJMeYWSTkk4ksd97Ei6tlZfYHX8ZgupCU49+m
8JbNg8AqZU7gzlX/vaBjB6GCEFkJU+yqNlNTizYJ5RwL4z+Re9/ozTAC1CL/j5dxcBdak5h9otSZ
Y11ModKGNu7rWkwdhflXANvGVrIf/QJ7DUlp0AX8SE2G+lOQoFmGtf6TMRPD/2cjmIyPG1Bhaa3F
KXqdcRdYDO4DvN090Ks2ypYbGxmeSGZO1pZKTxCjGPtF8jCYCD5o1myFHtnVMDSe08/HkJlRD8mr
tJuEAzycYU788bvkOl4vRp6kT12btv8ujS9dE075prYP+x6PJkRdPifX8dfMin8ABtzMySn+4D5m
z3qTQg3lN66ons+80fJbowYU5777gJOGg1n95/uOkXu7qZFr+1IFrbzttDqfhh1i0ZrpJKpnEwZj
NSlFDRlNL2CPMV+SVipn0bG1ky3JFTEygztD6I9BEjmQje432Hni8nEEDoZz5WnAot/76JNZXKwG
JQRGI36mDr63LH9qIAoNOaN4RUKX5TlTI2asZ2B07f/Cr/0w8OCvF2jb7VbWrrw0QwL9wab/tPMz
1JsUfaq7tn0GHfTXXEtEezPCSAjlQxwdcamkgdQ/Yt0lIJTy9Oa6ms94yPw+l+7KQnAVlBAMxMGB
Ynl0juM227z2+Hahcxx5WVcPNrnqNKsvct+eRt6Ad6TFa4rek8CgQMd3H9k6Cwr3absZYrU6nIQY
8C+BaiBrdJQjqCZW00NVO8Qcfscrr3C0NZJEUNeM9FWDIR+3Od2W66rKKZoHdw50bGC9fOOY4n3+
R4DeeSjDxaWXQQtbSEDc40qE4CdqipwIE4sCHtTrYquR43jc5WpHLTrsbpuY2MAP+P2ON0B+B4nv
LGgMSgbl1vYkeTh6hZAryNS8eybQ7egYkDkSRTAuuRk2331/WoDu10AAs/d83G69y8o8CTaBtCrG
OVKoIvD2cq5zgHLfvvFB5bO0IHGYUcSZEZ52CAzywQMbE15VAwfoD8Qsv0pKGmQwQVQaWM3JX4c7
bk/GwIfoXxVah1H0iEYA0v76E19vIbN4MXF9vK7cLKuDHFYX7WhsNzCwHWtnBmUjD1lkAEV5xpA3
9jNjlFzNtth7NiXdxB02N1GEURjA8l9UXA+g9po6y/yTDbemszBfajtvZsqB7ZRRL4/OQKtS6bfb
/oo/T92E/hiXaxku7dcEWWXPMEmClapSPgJt8LiCa0weC0T16gJCt4W2ol+p5Xtwb6YKZ3bUIFfb
O4N2H3gBnWJqbBjsL7iSXLOMRGF0PK2lesKATmMFKx+0wJX9svcblt3d/DYeDifwHnBi0zMoAoFE
+hAS3U/hImLflV+JcwW7XZqHcT9abV1u54YKam6awy7fTR+1/CLz8f3gz5W/b+xoTdpcIKRhTkFI
aUYMv6GWa8pRLDYJlh03gUFDVIbrNFor8JKwOMfU1DGjA+YwHvNV/yp2eTLn3Nl5P3ifwHWJ4lVb
eIC4XP85V1r5XxyCi7xqDeYXyjf5Y0U048nreLRIO7/GyVifh7MZQpFEi1k0lkoqb3FPVxkxtE2e
1Rcne1spIQsLoWWHoNVbfYHLMXaEAmx4GSW7/TfC/zpqN7qzg5oH6ElnVZB5ycigoZFY9Zs2xots
AcAiLNpFNCqk3pYIBA8MXMgTtA72oE1epUjSrdYcZ5meIMh+d+Tf5DsAVU+ZQ2XzYkGbH9Gq6bNR
VpScatyVMa4laz0esuaPegPl1t4pwIIocJW6MTwZngo2Pt8swRcjP/Q76SEcS8bRhQImuwRhnvmC
Y2RDe5YCE5Z5D37xUAdoImJp48/5FB9BkLL35U7Wb3frnWdk5n5V4W5G0/xKi+B1wyDL6YZUBiu+
nLnTYbe29ELd/r5QzpW8qIJeuQJWwZYVYmrbkh52VToQCqU2jlnYwm8cYOwqYDqTmCGaUL99FwH4
hQ2BDieOyMUB8cI6RLickKBoBF+sMj//SmFl6LpKzROIKSTPIWLDBDMv60ErG76NZa/A4M7p0jQt
IBArEVaB3p2c4jau2Kv5kpBRYge8gd+L8HpSUh6JqCkSbWfhj8eeKkLgLIecT2XmQaU8riRtzcmv
hf0Hi4aGyPH5a7gK9RkWfr+Eiok/JdpoXBE4aoRHen1BUa/GAJr1ycCnCJweIG6tCRFSCgctruq5
gYYuXcv73KjuRYCqukQ9m1wAGitVZKHQUrDU+0qOE3yAkuIXLqG6SWYSX/OY175od5llEVZziH1/
ldKj58O3wnY3ger2UPlqNTHAaJj891Mpf3aA8IU3QZiUfEEWybbcDwK1g/Gf2nKqZj6l0WvosZ+n
0DpO/8wKA4fGs8kQmjMgOIO9StJwrBMyUHguUcuZJ0FGbYSl5RVFWNrhBLqckGB/GzYl2XcGdVh7
qmro4E4Mnh0KWs4NLtudi/+X6TB1n+BVrwlHq+0UQeJL/7PIlSFjVjpfq7QIolvL9wDT2l7DPE92
K8gWG+g8Ax0sCAstPu9QckHwk5oREeqUVn/kDHZo31S6+ZVm/BZGMlLt8rZvftb07l9BgSphQjnl
Yb1qBIXS8TfbUCzvLM1NOe7/s6PeRc8pS1ZtzZ9EhUbXJYPA968kZtIWdmqmvFfbo02pVQavKnJl
59hVg16sJ7i7CRy1f8PwSDM8ucK5duFBIVe07JUm1LGtGsi9xhUss/D4Vpw9Ax1M/ljCsnTrcPrJ
pk9ONJcxNJTKXvKJ5iQgHbEDrCCNhtZYJCMT/DoNkrI5GkBoqdDv2KL+iBtZzI5CGi+ujfHDCTpB
BkhKozCHCSrSYOpEYSJjMbHRt2b+mQuctZaQE+9/9nrqeMPMeYBQkfB0UKxtr4n1gNodT39k+Hdy
mCthUvG6pcIA7tdXxrRAIrTyCUpm4I0IZ3FzS1AESoozve0aQAM8XyycxxAUznCiKCeE2lF0t7jO
6WlnVSbdjJjWGmbTcSUXrxiQrnQqr1Vxm6DyjvjzGAMQE+twI+dSM3i8LlaYWIA8pcQGKGrinPj4
5z7JrQrpfH7Lak7YyJmSUB7LKiT+PF6hqlNcZc6pSEKJWdHxifKUjgPY1fAh29RwXBYCSg1iDevU
Lv0N0KgHAvC3XEGs5z+AS/r3Ue8koBPq18shSa7pV+qLpnLZLgiCql3wT24Pt02O1MnLU2MrTP7B
wt76zys79dlu5hdDFIV8VAhzYxsdBdZaA7aI2E2RNGygh/0ssdNB44e/xN98h54f9smsiuzD/9+3
KkrHaJ6tlanK1VScoTv+eolQU5aoMqArFMMkLMloTExwz5DJcAWVRAYjrXsS+B4d/sOHSCe5uT00
T6IeWbruSZfxmU7cfmtTuJsQothnzDHajT0mA4rhmbcKULD9jmCxqNHEXJgsJVLBqFRWymoG56d7
QDbB6FVj7gGiTAn4xrCmxVaOjaOPraoQ1LE7kNrRcf4AELkbqyNaOVVbu29HPqtg7WnoaDUPg+vN
F1lUK411Wq49gzKiOh2p356TIQ6jLdy6xKFIorVoILl3G1AWo4vPHQQsGFPDzENx+TAqW6eMDu0e
Yy+2yxTv8HDniwfkaK11WIoAcCsG85FzVTBsUvQ4S1yMKyCc31qd7TTrX7HiuTUXOYXf3Ylh/2xN
lpJjqhSScE/e6QICceK4HEnKZ265eY9v8xrkFZspZVYPhw75zlP2FWcYWVBd+F+iMF8RmKnALqf5
pjT7bEsLnyZJ2T6OLu3O3NgP5wT9isZXaS5eDfzV+CAZmC5pOGmziy0bL+wX4DL5HZ0cls+RByJx
fnwRU6FKuREozF2eLpEGGhbDDlWC5CGXyDbC+J0t6CKE2+43Sg4WrtCG9hVeCRk3MB9nJkEoI6eX
vYAnCtpzNt2Epaie5mMJUmo5gI7wMCs7HH18zNnArISsz60HcxX4CvPjtiumLNIIXarhbwBdhQXo
zxEg1JRjZoy8XlpRnRdGFGzh5CuMQzrg2YYPIBmhDNjA3HJvWS7bpCGNWcokcYrt5uuuEWNvJilc
uAvn+Jo+rqVJKWyfGjSPKNvyUDh+ET3JzAzVZOhy1gFGE4BxN6g8k/z6zxTnuuHxXw7O6d6sW5HP
G+PoOHrdUtDcaXaHVESAI776MPw2MnMXN8PnEPTQo7A+tQ26FCiO1MG3r7X2IJt7nG1g6jRMmtob
DPlVhS2lJHbgcsLZVI7gxH8ICf78dTg=
`pragma protect end_protected
