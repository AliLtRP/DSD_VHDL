// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:36 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
K+Jm7TUZZp8dEZvF3DVqIelOfpxJnfkisCzMcryuNBKtlaHJqTMgO0upn6jSmWH0
zrBlFcShR42zDuuxc3UkvSVtXFdKqhGEvIDDmFHr/gwWWEek5b8/JNK8MhMFmrzV
v+vQBc27zOLYtntn2udTQx0Pe2Pbcu8alUm417uXE1A=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 3200)
s5eojcSLLu/cQ+EmxVt1KfG8Y0Yh0nFjN/IRqEMZU4v3x6N/6rSnspIVSPnnGlss
1uZvI4pwFdT9dLBJ+UQSMA6zIUpoP/Zc1mN0lAbB+ckF6OO3LyH6g0DFmRVB5M/v
y588S5WileFICCnGQidnGXtuZCzIHITS5hx3uJogdpPfLxxADvZDbgi16vlfXPXs
UoG1JV46q8BahodVhmNmdAR1ym0tJFT0gS4XTkU62Kl0Ge1pYSh4Tm+V+OJwoRO/
1TmR9l4Bsj0T2Asv3bV62f6HPT0XBPin1lyRqgLJ8hCYTLLmRmy9VE1pLPVWNSNP
/f9VESQKnH/h9x1Q8diaKf71hgsVYgvzkQR40uFLyWM0cLziF66FHx2vdSPAgXj4
xUwb47aV2bYg3V9e0RuziSPwlj7GBCdUqgybAKdoguEVny5lMXOapplfIBS36c7D
239bHvLcOBnIO28IeQs4xFjlf/AwEw2B25nl0UJ5zDtGeOwSjERv0jkFkFbbo29j
xp3l1h7XIPjSMGu3mzzLYfvw27RgS2wrMaRUfEbMiXRuaZAdCS1r3S/0vXzBsKvt
hqjbo3i9a/S79c6X/hDfWxoJMOdmdSMxJRtdTnJtfvn4ogwuSGAOVPMNqA6huZ2H
NJmlOI+OZb8MrHjcOyhVWJ1LmbFeqE0nYSejMZLR/2PapSwZBRB0/TW3aYdOK4n8
dI2ZmW9WRfcDGp6cmPPM3RgmYnHKWTvVOYoxu8M+oG9JzSZIpfzMB7Q/XhMu9QcJ
0Cz3EbkEPGiTATEVBI4vT7BETjYfsWl0ByqamsIGCPDokVkd8SX7OY+bp11aToIF
O3TulWlO0QhW2KC2/yiL0BoE6fR3B6gx84wPBXxZ4yemZCX27rZ+ixKSWtpjcbJm
eAU0odDQ7MHi556AXyCQ4uFBVsstfZxeTqfdD+meoiSRO/EueEMvWR7mYIVZFMM8
J3Xv7nUx9ZizGddYizGda44a0Q3h6X4kayzll6cX35lWoEAkt1Dz/lureRzXEiPy
ab/Avte8foGRGxMFqfByRsWyXGGvjviBLeU6+ZLL+f7bEjDdLB5Yt12vddFVCzo6
U4E49Oov0S9Zt2f2QKT5inTGhFlF0DMFPsL5o02Vf4iu5fKRpjlMQlp8yEyTYhMt
F63Fs3PFK4apsAW1nPcyZeIJfdbOvB4ydAxHZ32WpWKREQfI7gFD3cpxQZ7cXnIu
jw4BcUfBuYTlRam4yDw/mn2ne5K3jnn7o2Hbird9qsNLeWVhXKSNjoSGevx3Fsxk
yHe7kKDPXRlYpTbkZM/B6wCV02CS7/fv41+VqJxB+xYoKsQynbqkxoE21W5nBJPy
t2ggHJFCdgiERwm91pHykxfhnX9CDv1+uFdWge3aOzvuNHkWvdY3k5e4U3ofqFng
zePC/WybLwkb40WmDcxjYgfkHqp2C9gEE7UL1P18J1FbDgH1YHn/FSPR9Kcjb5Hc
JzPFp7WziMA6lTF7V1Mqf1BvPzHH5qbkFbk8m0xuM5mX6wk2sa8uqVwGUtqjsu6W
/nuxGd6byI1LB5SWCvfqkNllWo+gpmC2VS0ohweRen5n8wfdlYDabcr9UkCdqZry
CPB/rftRgoYIlGbitTtIgQ+cRrAhCbBtz0SyDPRv0F0Q9wXfxlFBxNeWPKgIRPz4
JJx6Xu3xlv63mBZyhOx1OPfai4teGDsYRhgplpCdB/KWv0Zq53nehXTs8Pc2jbdI
+jfvB3OSIAJaDvx4KHed5t83Tzeg0BhYITPzqKBPNTU/eZiRIg7wIzqvSIynPwQG
lTyVW1pKzZrD/E0Up6sq6G70aTryv8BMlGaKMElZW0ChrR/vlaNQTQtBZzmMJXdF
wD8P9ym53MS7YZZLcaP3lWQ8SjyMtkeai1FHk6zt8FZd1mN9OiujRQtOyYY4kS+W
w8o5Kcf3PG/UWxTzwuF/cDSqwX+UR3iGdqev68o7qbLji9aEbgtuAkj8jHMQCxwj
8xr7SkWpQKE4lVMyaZDtC+FzJ2HDgtcIbyXkVLslxw8kV8PqYjolDGPMH0jDAA06
oWyJcNRJ6/NxjJ63abPiTeqIXuvGnx6/l8P+1xKEuE07XAL++/2ok9efcTNcGGIh
JfTqQfngdn0YA9R8IPd55xDV81bwIKdulFels7H0BkAAryYA2hpudd5jbii06+wk
MkGbK53o6PG/jR5AqwJltI0O4OMo30hWyBb8mMAetQc9srFBBccvebXrCppBb4K/
Xd3QRz1Gio8VCUzz3oVGxsk8wF66n+YYT1CiUtPW3t1S9TBOJeKgivNddjOn/VSV
fEIuEj11MzQX2a/kanAAqqt9Y8lcn0W/MDbTIu5DaHhTNPsk0WJQ6AcXqPQveLXM
3F72wjqpb6hpW+SjyolxKMsdQt2FG/QaZyne6UHgTSQhrdB7khbLSYGpJCrKbl2L
tmvYh3Gj/WZQ6CFIsaWicxbDhSEFtHS3bWMrg6tyg7VDNRdomMLbSOOJ0+kKUjSN
zR7mQx1hJACWtpulGU8GHk+LPvYVIEghhpT4SSzmcBSbDfk1LT6OrwQQ2zWCyKVf
xlyn9gwIWSdAhe+SZ2Yh0KpJnrOX84myWmJ7u1NIU8CDHYwUKmtIvYYsHHnFUxk/
q0lMFKP7pBGgQpguFvGZQr3g2T8s1doX4Ij/kj2SlRh3AjGIFZe296pCZca9ktud
nSEY18f6Pii0BZXtzBK66rKYcl335I+O1Ty4lw1NuxHCZCTcPbIS7PJIf0z4krak
iPRl75Wv2REHkAw8gNgvtoulPcG3EvCi1oT/bLUVSSEntEmXZrGQUtHJeKqYoqCP
3f5U/Jwu9CkpSQDMpOiztz1SkH2+mgQRuD9HU5kdFbOtotk2uqSNSHU5pV1BD/6o
WKOnYsir8jpN33OT9R1U3qjKMlszhM9IwJ2mlgajK++zFRnuFsi6Ui7zkmzuM3VX
JH3aii3K88tvEsVXJZWDDB1NktqbZWqiRj8ae3n2k3HtRcWF0cAuc7r85tiiqAup
aBelqMlDayhP4d23iR2u6vCL8OpnUGw1Rla74eIiHr/k5Wu6zTydvE3fRn94CmjA
YfpTcPTyhlKW1zhw2IZZY48BablcJkimQ6eN39hbi3Kmyh28Kh4No5B9KRhZ2teK
qoT/max03IVNFE7yOFhYc2PxZ/rimcSpCflVJzEGIlUxJA1hQ2nzNU+a+JH1r4rQ
Jyx17VDpI5tht5AOz+6OtgVrT48Wpi/LAvRzUv9B0jaXFcf+Duu+j6LI0HdTXTKl
UmZ61l6ATO5o3yaI4/W/rwiOT0btcmt2pUWx4Za8fyxKb7hpr2HT+gYC3AHUnbXv
h0+82k0vDyUWUiPy0M/Egm9ZOHQirhAejzzxJOinUuHLja3fOEqFyukNy5xxY26k
1+bIdB6cjsHC1emRChvJdXHT/Tk+tAjqi2hDmuKyiqtErCwXJ2bCL8JAxYUbdrFd
60AdJu0iIIBpjtBywUj21/bwvGBoaBU7s/SYPt9FaSXeEitO3v/n6EF2Wj42pYsx
ZT+/CasvUQsPcncKW7JjxSt2CVMG5qQVP4KDq9tH+MYee1kawdJu9Dy0TLuKI6LW
6f41/NIHKFayZrCDnYUa7GQL2IJA/sSYFmDWbk7/fUYIxuGiVqfAVzJ/B/y5iStn
93JrbIqc8Tz+7D9FAdV9zW4dQODV/dk4BM6OxVt/UjFTRs2ZkpIIK3FyKkSEn395
wqBkQgsONVSZLp8+J6S3rppwzbAlEgd0QtvNbZwBf15C9BC3jvrbqCsdoBxEyuSe
rpcscymqAlXZuFBYpsYRzBk6f8xWlz2R80joCMvC9hDgU2AazRJGRQx7jS1RBrFO
Q09odp9WN9/C3fzv8Xl8vQje7L5ESfrRTsTrW9s10oCQ75Orw0i88RaHwtwIH7Jd
y94ZjGkKbI5E+WLj7My3n7GLD00M62j2e5zpI6DpkDgZmWjvM5nXkArXnko3xBBn
j3Dg25o3TGAO3qLf72Cw8RFMIJWz3hoDiMsmwuVej+BBM22zwWPWQNqgQoYq7cvf
JglORcZdM4+5v8p2ltcbwTYFAyhvp4Qqrs8bf0Qs9Las1gRajQBMCZvYrbxtMzCm
vfQUHTtCnbXDr05Bgt1JfYh6dXC6PP2JcnDoKydPVV/oLldwh7k8CRbDbAzRGOx3
jfxyVNK1obLo4Eqsc9Ai3VIIB102S//In0Mh9szzkHSE/CNQPtgfubo22WPaCdV4
EbM+FSqOICrotztrgyiy5YlCc5gp7EsJ5Kb0iA4IKL0=
`pragma protect end_protected
