// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:31:30 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
VsWJSfl5IdasMojKZKEWlAxtMc9JqJTs+dC0objnSDSErCfz6F5qKJeq/e4YR5AS
RZCYkbNDNSs0tVR53DS70FsXjUcHcUdd1bYI5W7EH7Dx0fz0QidqmvrEXk81sop0
3efiof089SORsDvwnkzTDWUS0DnVda6BY5PdOURngKY=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 63232)
8rys5DhsBpq1+rwYMENdzo3QAu/+fq3SNdGU4gqwX3yxI05MQhyEFOPJyiHjINLy
fZfg02G/L/HUYfkxPU7ohClsXOb6IjQ5GV8gxojjjnpQ4XcZbKdqXb2RX5r5KsR5
xVAIyqBslVOMnl/ppXhNuKHH54suwpSgm0U1hFY12vaI5GPtof7dWWvTwIf0y0KB
5cQKqv3zr5518nmIdNPGwJ3DvjUMFdVhi0xh1D3oeeG7eSJNNiNvl+7LQ5f3p0tV
OapkVaeCmznDa7yHVR1RpXKshQYJG3FBtG7p2RMhrCdbG+2F/5I9qORYQEhjHwfM
K8aE17huXe2y4DmlsgT7SUJ+SrEDBvfwU2HpHnZe9TwGfY6/QKaMu12ydlwkoitz
Mw0nqUeYVejuX3MaHXDVhCvP4F71MAyzWFPhgqDBcPdkCYQk1bpcZf6he7ZlziXG
UH+UIA9UlppOzlJ4jjWX1Vl3QNdf2CUrfttNNqrZtt3njdPyQBwyy2RaDiZAwtTO
TDGAme478Bkcw1Y+0WsHGMk3G0iEv3mceqEQGFpacyAPbp4YDHe9Rn2XcQAL99HD
495Xp4oK6z7TFDRs57//MGW7oaE0CkrsQBx9zHMBj9UPhtKbVVhp5qdywHuZ+HL9
Djmvq2cX3AMWKcVoniOplN21LmuyNdqlmRSjv/B6tpv3WdOgW/j97i28NLxt7mTP
gHwIJR3yb3xFr1CsXpFrL+NOFiE3IuRlD7D6EVw820IKMPMgQGMQzB1Ih+b6uXEC
A4A0E1nOIHWgM1IVEDeorpRe8RpIFjskqtLNvvO/5VMqhy5e5W28zzr6n1bezkKn
PwjCdvD3xMgE3ztS6n11PYfnxo3Qkg+wgtqgiZD7sT4tknF3QDtEH/ikufngPtOU
al+yEXG1BKYcCJytUeHYn0S3QnlZL8a7ArHv5NohXIPnqoowtSj01kb7psGQy5pL
A8qIkhSAL4DLpLkK+YcEfO/PpxnUbxe/G3vUsdcn1b8speuXnSVFmVUjQc21zFiq
eHksL06mDzBxlBUcInnhYAhTRoIdSoG4Peo0dPBfht+a+dZDxNslpcNam3GjUAXY
+FPjLG085y+m2L5ZR7Dsf6MLjX2mtOygOukQRB1Bdi0V+TjlsaaCzj/MTUaMvTfL
LVzV3cNHPtA95JqOpqk9NWnqhqCGmxPTyXOaNUjKxksYXmT5uB3i8CiX8vRmmcOG
S/Tw7g+6EfRutZqagWGDSttLmK2Scxw452xZxBkRyF549W1ZKeM3oBkzIK28zSu9
OriOMfCvkIyvNxhtEoZZPSbZBmqdnUAwRyUpBBFsYuqdtm9CCOq6zaIT/RNKoBry
b/HlDIB1f949KM3+8OAJODJ6G8AWqun3ZhvYKBGuzIiatoMBbL43Ulljzv268GI8
60Ibj6/WlJJ67AWv+OZoKK1CTiBSqNfR0+LzKKe/wHlPJpBznL1V1y1bhOOvm5tK
1NMIcXiv8TSfGKqxbac+X1vtKVUEAVaD8QP+KDtgzyBHkf5MzeG1jMnC0pIzs/gf
Lzn8Py5B380ZkiomMXr+bADjxggtqz9hPRcVSv5zJLbg7cOdLiVbYgkwxwppYSPh
EkIiPzBFfdx9FRy3Ft5M5WyIEBpxPwxWFCq1INvLT6R3ASTrhGOsWgIxj7tO5Fnr
/JlgbGDzFeSSwpwp0LXWV02AVCQE1pMvgv90c4X7/2NfuV3XF1M5zHz9/0RVGurW
YeQ3mJE/SfWKg64YCGk73kvN2grNYrYdZydu3aQ1Bh11n4Eh+GoW0nvdl4AWiksP
CkSt9x2DIiKnGiTVXglIZ36TU52rJnk/ncHNVufY2+6NAExUrMO1ZR/BhTU5Kr9i
xeaHgBBsoJJ6j2no4V8re569mY6bVjE7m1c7zzUWVqj/DbcMHR1TRm0G8G3tHZOm
t7QEj3IVR6vtmAgUX1tSURd67dKhSlK8ZJPzv6VnwZxnDOUI4cc9+qukyo10eN0n
fpXbO+pmGxwAmSmtBz28LduMOiIfPKMGIseTlRNN0ENSP5fJ7uPZxMNdGMxURHaN
SenHevxtYuxs8hdQby4lijspPCwPYO/ozfTrmdDfyrbOIwSadEbDs3n4Y6u+Wxlh
HNrQLSADM2gRTKF4jaqPGre0kXc2jbgdaptEpMCF0VL6hGdVdbij9Du3rb1gr6UO
asr1dfeXUTgeJkRxEZCtmERE9B/gcWhB7WDH4Vn+6PMj34BsGRO1JINewVNk63FK
8R1aWd+KO2g7JSBGvdHHRL506SUHQ4+OEiapof6sD3UF+6EoMVrGWaLOdenSjwDQ
GcdogeSBmjMOxerxSgdZynJzmMj7+zKBdm8TOdlRmZJUpPbvJ2Gb3S/N7Zp2ULMl
aqdleFmRe0CjvKsRI0A56XizPrKrQ147Qg5x5SJMAVPmbklLR6+SKDKoMOdnwW5/
Oey4LHs4esCTZ1wBCk9chbW1aPxmxxcmYtudRkcgvIHsz5Y+PMrTVlczOUbGdiQt
w8dOLkoj86XZJ7EQIWvgXYVgpkiSOjeTwY5xKtnUWX34MswBmPPeT+uvQ/Q/Swbz
fGqeHtzGiDXsHvqXLfH0MM7OFitmcMDQvuhUtmVnr6GHbcY/wVO37JxGYQcOxrMl
6RJRP2ZnXpxxhVxe95gqkTju+EgZgtHr1uZrI1ok3qvzAdI2ItMSzbUMPW1gCZ4t
869PYs/IYsL41oxHWUtARSyM27U/uu5qUtwJdyiS3DL+qswrqxa3wpqoHruaM8gG
wQJmYUDGBwctBS6epiDyk0BnlzZkQkFnLDTvIiyWkaym0R5ToIOzG31elw9TDlAL
vCvDTR32dKQioxpxAb8lncRjGp7f3G5O37IpwA3/RhGrJdD4tZLXm2fWdbK7+42k
6+0P6h140qvNo44q+DUMlX7N00wkarznHSxlgM4YEqMJ4zDN4eENxTKESLSbXz1Z
M7U9Loc9uU+HCY7Kha8k2FJ3S87a/iv4wspxZunrj1tVF5cqsSHSGNywPp/DCQZT
Cbzooz1mZEAhystVyQQEHOGjrSvxt+UgKcHtXa26Gy5kSTqWZc/5qkaA1ZwCY0v8
CYDV3BD2MKabbhg2WFEIDdLCN4OoxJjxstspISV4bH2Sg4KQdkoVCYseZN5bDABx
W1usxDJNfjO0T6KphBeuKP+dAO/Yxxl7utyPHXhgWdCNAy4o69q9QJDI3oyEMx0T
nk9Jv0dNpMwzGKd30d7p7iED9RG33gMHW91q3IfrEKKGX+AbAV3f9fIWIFsViZ5W
oMK5C3qCdMeUQMwCE4Lwvybwx8UqDpuTSZQ64pfZvQE1qnxma8ECt4tcaaeY3/n3
T41/BWZK+lLH9iYOV7s9C23G3N4JAVcPINoe8VXkAYHFjPFUwaCWpr4gS04SE3Jj
/UlBauDk7kgRvRMrTvlIzXVsT4ZuQYnsnxX4uv5w7CbgIn8MkSXpQRuCt7Fadum6
CR5iMAbhmQdysjv/8FtZ4zqqJPXrB4mdHgyuvq0I+O8RNJoroF0tMpHCDNcHo9CE
hbg9X6N6sAPwWS9fhtFxVBt+KNI47+mCaZgndZCNrGjd4IY9SVRRCvtSXKYWxUnI
ySvU9QGL3+owiuWJZIcAyEpvAF+/Lj7fQTdR2bhE75+KfnHgP/L0umN3AsJIy16C
qnr2qzgrsXcuaOJKIXTeb4l/p0ZgMtnpBClf24GnBCwTPQlS04stShDqvQnFtNMN
H130LlMTb9XX+R9dquiqT56z/2lYfzQ62WWfeF6/qTARq+JXjOVb+ilM+YCraZ6+
blozAQRS+r8S4mkhSSdEbIpVuxyYt8j38ffrBXhcqoi51JTQabQJQT0N98bvZhYC
QccaVN9m1w7JRJCUbrMffYYCFyoK1WuJU7/hgkffzFNo9TO5frhI2JRWVDlLezTF
y7ictHVqyLVbBg9jm+Ommnif1otgNGA7qEAdcCF/LZbLmN/8Ov1nucoCeK86C345
EGM5JKSi/qQsbD+R0it3UMhHbPl0h9f+5O58MCy2d7hiwoW8sM04dc5SSkbwD6bT
BzBE/EbTqIX4WMz3RpRZjGcSFnC8coECfUkx/OMIif3SEx6QCuV2cxyhCHxGp3lh
tTwv7wdIT8cI4nhTUBoUQIl4fFH1grXLjfJhSb04C5PIllJrk5Fn1SvbijYqagnA
3TWQkr1A3A3PRpbkYwnyI9173YTpK6KjiXcFxCVGFIUjJx+P93Q1tWjGW/Z8AEsy
vxvW9fODlWhrZC3EYBHHEz7s6naf2XatVTmpyP7y1VnCL5LTu5oTJ19VrBZi9b4j
M86wRW7OdBngpSwCm8+DhhwsWRpCZy2LZU4iX1+9KeFet6G2ytPt0Rits6Ux0wf+
XNPBKHQk5O4RjWh5lLLjCmB6h1LbNL9x19h3jahnTScuw27OwvxhCAJ/yf4pMckd
FX6Fva06+xoGEummjaPMxhzY8/O004j/PRjWNmPndSEtuPM6ZFLLpBvU3bemZO4g
MC/d7O27cbbkhOLxNUyz0Rm+rz6YiEo11NUvHtSK42bHrJsyZbOmpv9ZpL9Xew/2
efeDo+UD95i9nlGl4eCC3TiZJGQJzM2XD8rpbUy8YIxXsOdL5RHFrLmy+4yYmKsM
W0vxvXjrnc4XxlqYersJMtMqHBa2y+nGpZ6xcdQLaIJJzhIJSdAzQXeT9uYSCRNk
wOrbH7jjOIBkt2LnRxrOcilxdtEq9k5sRI3E5bSvZuBMQly9/vO8iJhK4etJ4R13
PYXiE+e9Kg3BYJv4/N/EhWf5BYdCJJwIYvEzVOPpA0vUhX2qplfpHfeLbEFSmiM9
sYaqtLs3rvd5HwRsC0Wv6xQb9Hu+0lb1l8o/B0JDvNzV8hKJgrX3dBvHSfcyhMov
3mR62r/Uq9hTQm8j6zzRPXxJGzDkM1CLyjrMeNlfLmblps2MOZns4EQRDVgs9jrY
Tl3T7IlEg88JJCm3403BuglOFjtPfmJMpr4zJ7JyaqV5bG1QRaiwdDWhryp1qrIC
vEcBL2DzlL1nZlpUD5PFd8jSVqzT6YlA3sqVVebKD3XzfGppa9rGygaXckSaoDis
xzLN0EmvPW7o2ekbLDzwFkz/1OdMkxiilItbTqwhoBFiwQiLyfTKRQts3f28TiMB
Y3W6qwzEOjf3k1DfcaQI4QbsAxtlM8jDUGU7hhdKzW2V0vrFw60riy05NdOqaUyU
/8k32dHe/9W2m24Cif5CNR2JZADqoVVti62yWskRQ1Ubd53rISiYPnwhKzQcnOPE
Q1t4Kd+vkNZF87NwBWRzw0Jx7BUKmGKG0VtjYH1e19gCx9qG2e4/ckjchjMkT6+I
FGjAmc/kVRVAHFJhx04It6uzWOHP6NzV6RmHIf83LOJCTn81bCZVpkTwgdzb4uKk
Lv24yawKcGUM6/YreWv0g/7kLEFUFuroimRr5eB1+IcVz3pRKi5k5KARAG2HVg+8
wWbfdQFLJmnCkcWwIC+odB9t0zQ9ZqZcmWooCz0FHKZ/HEFjOu/NbzmNPE0JHQ9d
OpQ/T3KG4cP8OZc0Ebf8AFngkwl5X5I3outiPUqDmk6lpEHPzzyuzyBR436cU8FD
SH+EM4qV5kOzV90mWTA5JQtOAYaEBjqDN7MOsKOLJeafRSxkoAKb7wlDIxq0uhDE
uXzKL7vscvsSDPJp2sWr49+AocIvoDJ3RsB2U3WB4QIpeVYkE+lhjsO4jsPxtdpy
KYHrhkxHMJyiAmpL0x5HB4+AfTmI/pYiKci4qk7rBiPEscuZWu+eLFKBSHcN2h1U
Gm5lE8ylynfutkjD03XvTw5h9wPcjTCEXGpzj5sAxUSAZHhgSAX86X3KLcuZb/M/
ydur6HD4xJ9QQC9pKlslCH3hAwfmjVtaUe18D3B3XZvlB5KNs3MQkPdCZrv0iKMW
brxR3mZ7pHHVdEmuI7223p1z8bpe8HkQdJ9lmSQ4rDg6oiOt/VNADxoc5dWyHoHD
Y8ORBXSeukrR7pfQtN+nYSAarQ6VAvD6HDopgNNZ8RmpzfmkZgLvERwLW1m1/67N
Lg3oD9cpPcajJVJglGqgvIz1i7WRZ56O9falC9RVoX/G7j8OU6XHPrqTKnA1AyYF
IxxXr7XGFcrYkW1jvPqzKCJUJpElgx2SZe85tKUvXUp7VOBoeJeFaA4l4g3xt0+A
USpRzeEPmpne9aTHiZf1I6cUVAOpkkYJJRBvuJhyr7qqtFGsQMkELseoFN90ITus
DhHpZN4kFBoKX63Mw4uzQ1mvytlAhpKuVoStTD7ystjcPCl9ol442HbpsaYLSU85
j0ItflInzxIVGS6DRn8sTpRW64mITgzKwuTJsfOaRAkreeYJsJriRepiLi3JfOzd
mTndNHZRTHxFMAxzJnsJzIpnfgqD+3ok9bMQXihXHiYxLe4M0gYWReolUXb4aqEE
CDFBcZQjfslHoXJIzgN1Xb/ASH308NI4OS7ezLEDsUGFA+TS6TTOU22VpEfKpcsE
H+zuaSnP1HlNnJa8c8mNe5SUCwa/wYkw9l+g880eqrauJSoSjEqHsor2+dhGOOrt
yVaGVMryJ57mrTud4oyq5m9XkFQdW9aQAtqMQ5/NtWHP273Zt7z8APsjMLB0FEIW
rqLZokb9vVe1XYWq2uTmF8x2gzRozGyfMdlDjcatYrkzsHB2vWDgCnRtys7G3QKg
E9z++7Bkfs/+6SytiU2Ug7RYsCyN/SNd3HEYTnhrtrNqx2fuJAScfGPwZ7dZ8uUZ
Osy3es7O0guv82fdb5NTtBzOPi+ajjl8sJR1nwPpP0UtQgB2wdtL2ZYnWrrJPIBG
wbSllV9xe6tfN5g9CQw94m/lvY8LgCwvDblgwp4i9tQwYemCDCxzQXYRueKEbdAR
6lN7atuQpKArpBovhEh1w8nUj3zP3ZkSkVlvvkYWb6v/eM2hKvfellTxJCwnC7AP
kRGppUXZPwsdRCDzEn67GE22FD2vlTFj9dEnmumBiGYL/pER/o1R34RPzRPaqbEr
DGpxski4QAYU8cnMbsqND3a5UqS9OOAvya8mJOsYmvlVvGVyiqaglXgkzEA0bzyi
Y5MZUOVAnybuHf4iSQCZnulcRzTFndt+cTT1BvcK3IJb7utspp1ZVQPsBNYZ7gmJ
CVNYI3Axhk7fERKOLFwCq32abnZLgKuxsZ1Ou78ncY8y8ZCZPhT3DpyoL4rB2i2d
ik686g6vX1nYSl2+Tok/RGlM7WtHdLmZgI22b+Wx2MttLue1BNC7YoF2uH3ppjlH
vzKMOBHK9YmaT65wO+YKR36K24ogmO5MTvNO9vaq1Wp5sRJtN9jvGcZsGAxQH0eX
FOl5eqgNMzqaWuK5nTZ5WtYeU/qZMKPw8kOczpR9DWcVVSv0DYUuO8E8gzWi2I8a
BUuG75FGFGeqmElH5Llh9oHG4YhIGtlnTIl+VLDYFcp5jms9yLbHKRgQFeDOfuam
6Wtfs5Rv41AC58o0jQUVxVgXL8YcTTaE94lCJ1lcG+2wBnNIaTCbAmixbSjcqjwx
/Ilddm0R7Dtd0qMB9HzGTRoKwDf5ZQ0DYJhc4gfQZNix3jAC8Z9Q5kmn+JoJpRDx
aS/QI+MAqFbZ80Se3Yd/1MdS+n9zY/smAcOVxl/TnpHcuw2/tAn0sohEwn3qIM9A
N3hNjneAo+Ksn2jJjf4iQw5YfTbS4LY3XQjp/v4s3CXbDi5GNhRPmHCx7GBuypHS
t1JO1f6VhK8EhipdOGJtvAN/DA/oXelPKKZ3BRmiPup41SdgPDzOe1If3GtD7Yty
WkGFrP4wcMmJfOODhgJeGMXena3V4pGB6sII5OgAqVwX/E+zY69HRgJ20kW+1Vla
tw8uyPI6V/OfAYL/6Nyn11J711G07e326O9LpVbpy2aI1w4u5zchh8ahkHIoRcAX
l7d5Bh1/p/Kl/CT1bX3+U7hv8xHD2Ws1nTboGFomJBDD8pLqQLWZSoA7UGoULolC
j91T1seK4vxitb6RHwX1X1HiRlVP+NShmQmFTgCSUEzNGBh8ZsgQOtkcN1TXWXkN
nnhvvmvvACxUsOqnHl7In0HorwiGYSCtCJ8pSXS861YCe2qEkkiv+tsbkGsPtMbi
tYejRlqoNlxj7GQP6Ufhj2Qhf7IOTziY+XlIvNNJBc2pWa6QEtZvi6568BMjrM/y
omrMQT2ONU51gRsz6Iy90BSjb6Wd6PjmbZf5OhHrQSCBeIp27WR1auu5aWVvCgss
UnZswXd4cr3Owtenez6Si+eaXrm6382guC2qxqhbiTb2gLJz66CoH+C1QPJsJc09
uBj+up5HDAbb7kDcdAKIeatu6kh8I4SJEpw23Hubtnnpkd4wTBMTQjUxOI5toyyj
p7xbXjRNO6vOYVMDcPP5L6Enk+VMPhvNf9HQR53GceFbioaFTJPukFTowy1fSTBv
eSukIT3sA5xDGJRNSIiq18ijSnZ7+/JLmTLH9thtkhVJ2+F12EAQAz1+GXHKPIWT
0fyb/2o5EFIWtMOoYkhakP8G1W0euz3D1obIUSsVmIequLptByvpuqwfCUM3BbhC
Nv0Pem1V7z1MfxzxULuqFbhtXB21Qr14kZQqElrkEzw4TNrAD2VsaJfngXoOdscF
Dxb1Bq3K/apdLpjMm5w1qYtdmOhVA/UBtF9+96DS+AK9Dkbfst3VjrBIDObSnUKg
SyHKX/fhztutlaasty7xPA8kuuNgUt+nK+P6Xo7hzFg0pTgFDIHLqdLXZNjrmQ4J
38zKmDNtT9wP+ge0FhwNlDhSxxmr/Sb7H/k1/xNFq0nbRq10zzaFkwfNDim4bS+Q
lvVivNsEGEMgmoBlQSVLE1J6vxDPFMXjv+eDjDb8CuFEPTwrz4CioQVgAWT7Gzp+
ThPFyFY1xjsNRnxku6/vqWCWGN+db+X5xxcKxEKKrhDe4zfAP1AgeGur9ukMAHbL
Fx99keYU5FilPFpw81ECuPdJT1npVf70obUeuRgRM9pZBpqsrjTo2hcbw9Zios3B
mPl2j6hCexzcvE59AHroR8JstJJu+ijS3VlUtHCQFqJTHad7WlzEGTvFOSjtI2ys
qfhJBA51m1DSVbN22Fh9QyX1oHC54tWPWrauuJABUGfmG2JnCOg8o5xvO1a4j5cx
jzz9H+KoSYriBd4kJv7m4nypiUs5sPvGkTqHaxWAalinDTu5KXnbSqsuY6R5aHXo
X3IYDLJiqKZDBYWVvMEfFzr0uo4sPOpwZB9SS6WoN+kT1+6BG+unpEpfKcETueCi
iq1SfdybTcTQwQrY1O01GR8iU9bA0pLD1BkZ70FYnOzQxB9KZe8t3LuEzSaD/ha+
TaQ8zoQSfL9q5ovfSfrEIJdFNKKeyjfCMkURG5zYaQvesasBrKGBjzFWKJ+2+ejV
qz0moRZKd73X5h5wGFUDoE6qtUN+hdgVazpvetgtiM84SPzC+noZxlfdia1xHqUY
gyO0JsdK0IdC/yMegLKztJfgjlgELiRJzUxNLyB1C2z0bFemhTL35AuA4EaNVA4Z
fVYPqFML7399Kj27dvkdyRl/8z9sXhSfckjXmpEmeo/b7z4q/mFPvcyAppHdPlRB
frwfbtFk99oR1WF0BadMRBdvU4N4QYCXAubd/1qIg7o0nbQdUSIoUwKY/35WWUtE
4OVbZrTmHOTVZRunk+bhepKr4x+7y4IjJ/x7S2S0Dc/YKYFxBRe1C4zXlQ6bjVL9
SMhaA6F77VV9RlufHuXZRiUpMMqSFukpvE2KNy5FP6JSc6NAHsj1xqjqyzqydUTv
9PHWLQijf2JzQ65xTcVDksLNvDV+i6AnWJWxaF4wz6yZv3Ln+1IgU8EbaPs750Th
tq0IcddtV1UbQXFJwYmoxfcLttXvTF2kKJGyIDa3wUGZlFoJTlV6yNckpaPupC9Y
JU8BbV0Ak+07IFLBIBlwe39mfTqwLSUrEsJXlHedwb2WNRQIXrpIs+4OHUTPOplS
sSKI0HI4de3Mjb7i4R9P5/vprsqXTF/DqXL+tnzdi4iukvwWeGzA66aCHSNuJmRl
x3z8yvNcEaXR2ew0RPW3rLOIu/ogUFldXRTRgekRkahfXUxXrbsSIFecVcYYefkO
b4mlxtZtler87RFNtVgL6Wj+1/p84A/s0EmqmPIlU9N4Xx/EbaJFMOoC3hyt6PSA
vVqxcZhL+8DwJjf3ASTvvM8GfWm4Ljx31ohsIATFOciBBatWITJi5U8c5VNJW07S
pjR8AHEWXpFfsU4nkrLlZvxayKkEjZjfez3K2jMW1Xm+mDopVAxk56537TA6oEOK
NEa8YF857MiCoEYmr+YYcyMud/jdKDjUiS2+GNU9HqU55DEBdBCQwfBFPJCMDUWm
IAjBSJmw/aTIOZ+3wiUer07zlx/I5xVmU6odNuJVGOVoGAPzTxVxlZCgwIukAn4O
4ECOWOLwZ0J9WTqOUyyysPxF3UglCk6M5uJkk8FFDNEkfJPvzfcp2gOXpo3HZhbH
90LnKe4KdAgHSxMyr9WIK3h5rVWmpYP/YU+lBsi2dmMzL+kkcjItwIYmz0hPI1jx
UBgq2NiEY9gnMBBahUnrZbWW9u9Axrzym0S5BZ3YIuCgwE/Ube6XHzo58H4iiMKA
DutKvRMil0GS3PrZZq/XzeuNbTsEps+cSX1g6sP3YvBnFZKK80W2Y7rvMYbOF2NS
FF7046ocDCauaMtXpMhEoishAy1IOIfNCfz1vQEv3kLoC5yH2X/J02wxyb9kYxv8
M86vBWSIRQzV94xgfBO59lJiHfL6JMxAXdUKyF4WLMbvFPL36eiva/ks3cUyAyQJ
4Cofvnt4K4amazn5LXyurjhdIprZjD/Jc1+t0/yMbpKUP3aKaS5bwXkXS0+LRIYe
jwJmz+kFGujXsQ1HEk2JdAKUe7oWQbdgNV11jUhrO0tolIQ2GMGuKLrpbnFnnVKi
t/7F+Nd18BNXk4ZFhmt2HV7IfjXocqnDcSHNFHYiyVlvV31tm72sahlCzCpAzPE+
xeFc75sqw7/Px06Xi7i937Sfcxpsi9V8alFnApUwyyPqWH4/mDaP26jln606CJRU
rD8YLfTH+RXrkow4qNuQRN/X0P3RSfLFWLMs1tRzKXFvD/P7U4EqnfgWX0peOEXN
OAzYfYa33Y1GQcv/uouKjoIF1cxSuWvsY8M9VTM803PvYCSP5X6RCZi1aBP75+5d
199gGZ4p86wgqOXrvdJP393udk8NDa7rbDdmA652fIYJknj7D5a2sQfvahoSLUg4
SCNy3gqZ2PWTG7LxvcuvvsV3R9ZT2ikx2K7ORcfyHbMmjehvte9VjfkrjxutaVGJ
irKAurvNGaEMw5ZqWkdB2FLmUYwHc9DMpDTTqHOZ9pB321kg0A5gk3qIICvjhbyI
gp9eSYI18QNtmCvMAmw7YBf7lW0ZzPCu6+fNe8Quk4gUL+v3SDfufcjGjALs5Hy6
Rut7C/t0o0V0aGCPhipA4Q9dshRfAG8TtkviSiE5K3CpO9w3lUANbVFx9qL/8VQZ
S4oum/xzt8xhGcjDHBrt73iB+l0Nq/u46iANLRkppnwTBWPevSFdw/HBZVnezO2l
oADCvOi4C0xUa1vKx2p5EPdwknp6Qa2mTiCiorASw4SLG6XnoCPMXBbdRSTl4+LI
45eCVTfQkbl7rVVeSjp7PgtMRemaFtGEJ7Upq0EH8OudD0cdLr/CQDKmEMqU5ODL
U/60xSNHAHrxz8s7JHQMplsFnHuCdmgvYRsVZq8zLRkPG/S+kc6mVzBsNb1TvFQW
RzQCaD+sa2Hjk/QyDwLxIYsdp+g8hMjveTpgwO6mXMbWwLGxZghDHzGnZ2QVvXjz
rQ1Sw94u8sWmbkpJOWpU+wFUTLqnaVHebtFpAxDKv0KD405UOYFfQpn9pOPqHRai
cVXE4lCLr4ewS4dGze27MFS5YAC6QG1jxgTaVe4g07N7ctbgBqDyZWXLcInrxZW/
8+UE0JRdO+/AYEWXvKeAV8G427D6fLiKpgK3ityIJ9mSwRHOyHzDHrQx9sDgot5l
tuBN0ngsMKnCjOEiRedlmFhoB9mtbrQjyJs76G/0O0hf5QuE0cJvIf8NyCnODX8e
6m+/hqPMf3nC8VTAAkrSW0IZHBy3X/pgqYsSCXsmNqBNIA+Q8KRo9rqwB63Z0TBA
/dNsuYFyJw9VZN3zt1m9fxzqgF+HXjUsZ081PjKQp2+X3bzMot3ItojcFaneZ2Ij
5vw7XtL3rcxCkumqHjNqWCd9HFvS7Ylps6WkvvjM8wAW2cuxrQvuDcCs+XjC9yDT
+QHaY3WyIWQC+tgGaXi76pmZvJFN2khNUbtEQT250/QsS0FxcLk3RBd2/2nhlUtH
HFgGqHq2Q6c7SB/6ZZGKzhX+IDTBnQHVBZs9dy/2QlvxBfXr609mbWWPFtMOmySm
cZEkPXZLlIQphj/fO4vISy8uBCL+tlORJp9D95Z1CZPQIW7lKvK71eqJ6ReUqm2G
shWOwQbSsol8RxGGHAlfza9aXM7oyyVhSEVfde2SKkLuTnBnN5E8q3cW88olLALb
ypWY8Nl5VnHXENoIHfMe7xscdNB2Eyye7RwnsyP43t4DSmL+uLlSLgp35FjbbM8e
u2PF3XZyXsvR7j6NHVEQC8EZBK8gj619Foe5R4WHEnUyYe+Ba+LrmnXQQIhpEUH0
9D1riVPmZVn2IcfzaG47rTlijsxhDCDPQkhVjfJY/B0uI5vkja63AwTO8/SGcrIk
hjvqg/zdMdMR/n+2j0w6AtfAOHcTE2JVtTsrm0qMew1jvJD+K5KtD31XO34fiPYR
pCeRsTsVVmenGb+NxKKys1Ks9WM0CwYAvnL+w6EsAVYUwTKZrPn/f6qfFqFmLjjW
9tXp5HmsEQnOpL+oi5k1CUv/wGJk6XKL0RxbOKp+euPL/uXJIuBqotMTS8TylVFu
io68TdEPu/aRPS8c433yd/eJsbh8izOxjnLk6w40h8gZH7eZ+fKldTMjP4mNgsd5
l4Fa588xQHz0mdHXepFj6//h2/gUYL8LX6sv7TQ9wGe7p0bqPHuz2ZUBDii9Nbcm
v2yKqFMQECdO5cbvGLaIwpYUdBBljG0fVA3qAazBU3vHbAPyVd6c5G1YMq3Bd+4F
w3q9Wk5ItqGEUmsglyaTqjlHXIfpkrGYrZP7/YUWFvw/1Hv1TDtBCwtM9B8OpHTq
EaSBuLqCnxDFMFoyoGHa5mnuSKrikxaDu3T2txPS7nmx1NfZAYBEuMXBVtXdRTkB
cMjvcIiNvoyjkBjAIspDefKj2D9kFIN+Qpp0AKhcphGK4IBjdd7SRrzdkCOs+s5E
sFQJeigpLRx9EdGPNWJ93Vsxez54NWeyiWLAX7noHXQuX/W/IOJraDFyIL3k79Uq
/8ReR4dV8tu5vwnwctG57XL0MPtKfBefNPt6V5BW1Yf49qFgPIEc9dU47dT/ZWFV
L+rbZvk31+5CB+/pzQfy7ojSIyvbSmtDfyFRMOjKJvZyXfm7T9kd0JMxhLle9tcs
64zb713rPp5B3N7GmZZFfAGKWO7VLD9IgAS6C1/YvkMOx/l6gGjdRSREU/FL/u9I
lo1bFweoTUl2qrjxvWxro967CW6EP1/lug0rEKFDskjKRLgjxGP7vhiIH3c7+j3l
+K3SrUhpW0EULyziINaF831Op2mOGwQ63u4Mq0jN9It4X47lXseHaKiPTZZ07O1u
KFq6fg82lKbHyItGGFdkctWa6CsorHXx1a+d4diRtIJsHM4ugsBDjbC5EkYcNSkC
BllNpG8AvWfj9QQW3MnpcU4/OBIzB6nZWAUjknYeubNShXXLFS73nTrkZheN8RVo
CByDlb3K3y7TXyGw+1BIBBB/DyCSWIHHSBkEj83P+oQEBJp4U0wc5XiyW8SOH02v
6N2tgfCzO/8ivV7JL32w1x2RkSCzUubCv5v9LuNdgzx3BBXZL5mMotkAgvELUYgx
YYYIWjuUyDGWoIbEOsvCtf7ifp/mJO3c+YVlkYzNvqjL6faFAmPuy5N5tjZRM6o7
WXK537Gb23EPGQE5w99kdixCaJzVw+T64Zb5t/GLQTdkDeJLeo0SHTVdzLscsLeT
dnk52MybwlsqhssPlD6SGFFwzUgjsNxYyAvykLD/lKWzoqCbtHeFqZFdc+KkXLx2
GOEJVVzoibejdaNRDuysWFEV1bDD+4XC/l20nEVSDRqG8jJYuKXjtk38ljma0RKs
9SFMrWFkQo71zCzIZf3SdXJI/F1FN5lkoJuVY/tEiUnpjz7hCEYwxBDkbGckSGPO
vJjDGyQ2hrTgB5/6R63yd6szeNGi6/HkWp1RfrXjPsPEyVlLd63s6NYCzErFaIC9
iGXBQd3LudiXUT3umGHXlIX+CYckl05GQRrU+Q3LPhH5StaI95mi52jMWF6U3Y9c
RfX70nvLkqwNgIiu3GTXVGr+t1ixOQROihVeKfmxo/H7gE80xGllnluZjgcwNcsn
wktak+BljucB0YoFj7Ig8TbbYXC7nTsjiLE3uLDyhqwKLzMoa+TDd7I3pZ3j/L11
RqOV+JLhUeMdaH1QpBYWrxfFVkTDoOTkbh1XsYqn3FQvVcV5qBtZgfr98kwlyIjO
wjB2CmPZz7SoHcpPNXCcukvxO/2x2B4cPY1maNnS2FVC206TXGw75pfdrgQ8y8mZ
tF53tME0/LtrplihBMhJWMg+zE0llY4Gsu9qZa7TEHPloDf7UWFfcaqCZQm3gzK/
DbE5lCHbt37YKV0L6BbKFwFiSLsP9XPB+VIHZEUUqopuHeJQxoki/bMltRFvCQ9b
z7ELw0Y+WFN3utLhdtg+9LwS2AF3Kq3FDXGx483EJRidErLjchIPeOojv/BJLp5P
GtDnPOtBrip/ZKnMdlNVXl6lYtraZ+qr/UrNClMmfu/KY+Y/znA/DM8r0n8ZItH6
oUucz0RPDodKzNotJY8kXsFhVBJLRah+zwyEiWyziP9CZuSJ1l0Gbh1eDqts6Crt
nVNuOy5cSmRGYOpeWRPaIgMNMMC209+kav1EvKzI1OCdeTCcs3e9JbVezmDH7izJ
fm4wfjzbfWxp20MDGq5aM+kgFojPNnDashOAFvMwG7gkhsapwpuc8udI6J1wdOtF
fbtU10qgBo8qVEJwncFfFh7GtR2wSUQ3EluRGHTBfXpPT3eKDlaFJcCDS272RLS2
9Ad9x2hE9zb/BON7n9dUwwCsl2bfTfOjOHp2sWeRVfAVyhY9Vtq+K2unirtejVpD
rO/nK94wrdVCYq0cZEI3YyXuCAV5cGJKLdpYKtYqOhkVdCkDrC/mlcz0XeEQZE0x
SdmShrCq47qfMiI7wzBx8Sr8BNWxavYxyHE9QUF/QV+bgOmLeT1ksdMjIRDqF0Sq
RIPb2JnwJoK3s1mDHXFKo0a3eVAql7J8wTD7qcydyKb/C1wiqlB4jPOOUDdlAR76
8IVzgItbX+DXXPSWK3Hu9JKyUpqNyf2c9HP2l6iKF+idmbORD38lFcZfz5nVwLC6
zSotakXlg9unH/GDeqFwHvnWdNP0hHvMDrdqkLo2fzu26LdXqsNH4iuzy9YBNkbj
SnnYAaXKdr22DJY5RY/YukicH8mEROpOC7nz8PBBiEbrW2D8fyTq06DW1vx3ySJB
NW8j4w/vvaP9SL3HABCXQuN6DdtD8Dp0JIfVFaDoQe4MNFk/WRKOZbLOWa9zUU41
JlydSI1SpiRxgZGCblCJhTX7AKbn9vWCfNzaci5jWRargvXwegytn2uV2EdeqjlD
nTEpgk2ETCMovbgi7CyGglTAHm1VIeNSTaxCWT/TjacmdXdyqt2PEB8XQ5ig6hHu
2QQPGodt6Hf12R59Q6ISFOZGLTceiFZcO1m1VQon/WDyMqpVtVwNwKTEqGS2YdFb
gblS6jtjsA7T0S8Pazaukzgv+9AW/MFLuRMaJ9cmxk6XBUTg+qB2Zt/PKD3DDqpm
kKT6zB97do6hMMS+3JYUDcb6CeW0IFWPnjoOVYzBzryXMfE1s5+Ks6+f4GaKFxBu
w1iXbPNDQ5NcJaoxDpCO0VDhmycnmFb2D8h+1PUC/gsWYw2zTfhBHbp2otkNQrYR
0JYg8X0BIRWycz0aFd3R1Z9VWhaYy/dAJqG59pOAz4YffZwb9uZQPCkawDvK3z+g
t2s3gcZPi0xfeMjUsQW9IfC9V3tj+WHHpJLW38g8pZxNuo8HQk4zrrUSJbBqce/W
a7BIKyfp5p6dHp5++L//+Xal8Spi/VYffZiEozzZn1a78Z4/V3SwQHSPA6F0IftW
jc14EaXpzHSc24euR1Ydb2RxLi8Azbaxlpu7eoCLo+7SdPvruocJIvPo7VMKNGaV
Uv/2ynaqK4P94ffqSprd86annSOaYWCMBGPOAcuOMPgDZ1weiUwcxsIbEZUrf36d
lM4q3rRrgjgWltqHAyba6a9t6aqkDWap0LzuAKcaVaX821mjVkyy/2/n6ZbAy/5a
xmt5yls8ftbNjiFBKdrPPA04+cCXlXQvhUsOHzJZHWVch61DFYdFzt5qPjZmc6AR
9t//NCdTPt/rJ5fogSdYOi+ts50zOAdtEB4fs96RR2UziDLBUFH2osqki6JtIMrz
utLls2r5PC88QWLVWnpufsZe8ZlISsXyTvCl13Nv1RvVF7+exNg0nkuLaqvX93ME
jk9wHtJu+vJ1cCC0jjjvPciLDkv60MQCPrTiUANVE5/lsr4ZSvgLt6iemf6Q3BMn
LUXusybM9x946FKhGGHFOQJzPaHSOCoUoLQLZR5R/BNZBr9UrMXTItJvAySsG1I+
oQjgufpFOMeAfQSS/shT3itXiSpRvKX8FkfUuhyH+4MsMNrvVD3ox/3h/ff7f6C2
TPRpA2rZvtplIzdN0vSEoMEtswo5GWTK+YE580WmXNq7xpw/MPF4nFrasbl1PaR3
RdNJY/Fc9YDomlSWgSzAr8EaqJPI2tIZnkcb+jxmpsn0nxgnQV+Wv2Z/8IVdx2l9
JmoHsnQD36USd94lQB3PszEijgQBVPRI2wnVWZkEXG14jBm8gS3OORXgCm+iiVU1
zWGFEVvQz0OmlSaYkNDRsbpzN15/PVZ/Yis69Z5GhcbLhwuLQq1GzfU88PwXbFl7
vIi7YDZs45MwoB5EMyoxYufC5pilLfurG1paia0GucdUQFe0+jFEe178SuSf8UXT
X9LGlbtpZwXfjoNBnxcytOxwwX25+mjguzEqBPrrgn+LcVwWlQn6xW5uePt4lijx
YXcawLZh/1rXhwSbj8GuUnh/D7rQLwumo6RtiDDKm6jdfV2VYqm3M8oowE75gXSh
MOIWTOUrxzcWBvkbHPE9vDHaqGYyJYK+l5c9O79VsjvkuQysesgXjhSd1wwT4owi
nP0eBADI5L2az64uUAssowUChSb6neGiQRJ0Px6PIU+1yrbiLtumWiuHMrrWJhVj
vPnWNuIy1ijPAeBt3SfS0Oy/p0+Z0iIOOgeP4PDbgycbLPclyKTZnaYJJjK6PYY2
6QdyyIM62ecwdMqyA1XPU2pEloQ80W40joObHY4mP7kuEXRWvWyBHErliKeCoAl6
Mk/I7kTGAwS7wfBlvH6wTDtGJNKXf61rBmyObhvsdk8e5SG7tZvrU7aJ7UNfPA5a
4F6bXro1sVWimhdKH1JjqbhoL5+D262+Q66ui47vKo9ZzdI0UYUw4KjN2eYGQidf
BNR3ZLi02kXxdtfaLFmMooC7+kW0N/uYxx7jBLaJnVdZp1zQd72gfk939MFM8rUV
gf+S87ZVbopn+rlkE2jmFfRYdL0nIYY06lhfJTcq36VlF7PzuU1fRT2nfZKuHtGv
Zj60cTAjzIq5BiHd9f6/VmT9ZocN66m7fQhprFc2dkqMnK65Xr+HLqi3tLiwd7Vi
B8mv4MESpVquRfmWNExf79FZWGdKItS47F4/ZTiUQTFItQn2030tBJdmPXet2m0M
wuitbkEBf8hudCxPsraJRqVpToGSLyxDS19HDvFLAVBcKanBFEOCF+jcKOEpzmFM
5aaKop8yRQ5qc8d/aU8yOK9nA1O3OiogtukAiSK3mKrmtsI+a555Co+wkZXBZaHk
po+wZEZh90FRERzhwnsCRPvNumZzccH8edn1ckwzC30TOxGLpzqtYLtnJKTqfPzR
TQZmAYWWIPqbN0J6k7ft8LcR+O7Uo0iRHVf0Q4ugGtdYBKK6gucd+8sMdqRqb9XY
cWU05KqpdRf+BqJgdPZtSSY32Ed6otvwjlioKMwtQV4AArfznza0YvUGURTv5zFS
zjtfeaOvJbpsJp2mcx2By7z29bUd1tAq89YYzGZx2P+AG3Qg92OL7PUMASVqfnxW
2OrT1URbgdGR/i4LBW4uO+vfl/XQNjftMl2ggLuQqLen4yEszR18Pmmc44+sK1PX
FLPsGIRHxhVAvBlOLKrAJWAtHevRAkU7KR/o1PUrtY0sQ2GG2LXJVX1UVVCsJ4Kz
8IUSo7k/WlCRGJGCi/yh/twoe85Urlnibksd9nbKSFnxOQ7kMl/8ZSduVXHEHZ/L
OcpXIjdUyxDBfu13vbXFW4rm9eNs4YHkWesAEqBPYgCYsK9zV3iMEdv4WtZkUjpC
Rl6hlYDlM8+9OE23B8ha5DcudG7YSzwwoC0GRMN3Ror9jXEykGEr5Xa68T9hvol/
KC01F5BNEaAOLwtxMcXl8n7zgrbr8bTAOczvMxwYVKifFFRLznQ6YAHFsxGUSWiQ
BOOTazYE7WC1dFym6oFCCaEQ/itUm0gJczQiwD4FY/2Skga9djgMY2FhP8Ec+gYi
2Q/hqeYh6VTKH2UJfak8/mZpcfyC+lqkv7kvdSh8TlHN9QZod7352VmgWQVESeAY
AKOtGoD32Yb115y+Yu5GPsuIFPvAbdK4UaraP1d4JcBUff2Ecux55Snl0a5rvA0u
uyP+IptpsDrvTIOHBE7h/5e3ik3dtSZWuQ5SsQhs0iiwpYPNXSBfmIHhiOHL/lmS
PiztXPKy46WeW7vB7yDntoh+hd1FmL7AFNTp114OUFLt17A/qMYDKSJ1o6IZv5yI
6FZfc+s/EL2Dh6wkhANqOjrBzovZosGB8p7cqYXCS4BH7Zzi9U8bS68fUxK7RH9Y
9AY2XgHr273I4dwhOy0pJaiR/zxwVDtAs2r1IcSKnTcXyLxmD/KViVMSU7MM3PZf
bkdaalfWMAQv0kNwNJEZFUZe03eax+LRVY6DfQZ8xl7WW1F46/FhZIXE+Ct/Qd0L
+DIEf2S5Lj0EUzqEYb5yk+2BDHvdLLiL7VmSfLA+XaxzSpPt7r5V0smz12zsBOVK
9/vUOcnN63dMbdcjuD7u8Se7CFt83gdH+gn8NCLla0uGQiu0iTx8Gxh0+i4Pr0eY
KQXduSRcW89uREx5WkkOvJaIS5pFaoAsds9dZ0Hpg81bowLWjrCizbBtXk+f+EWV
HVdE04b6HC4UhBvjVDz/C9vDXbcbzdnAPybJtNiI5X+ybAoa8ToAw/9mAAEnSbLW
0JLyTqsAt8173t0OvbZugQdrxdPgZlSgpZIerR4e29u4soPspkjtMSTbeYPwG+j4
szhNBqMKXKxw9aedhJy4AOpLImkhNoHpAT//DEt9wRo8uUy5BzixVzfrIz9alGEN
NpW070UTOqHrLt5YtotHBOFNaaAB6SrBUBIhIeyLMdQX4q+5dXM7Ml011No0U87t
sT+aqL7BjLI/EL/ZL/tVRyv07XEMS9s+G8Pn0LvTPFrLyjXBQzfrRbBxs2Qdfu33
s66VAATbhNnFewTZH7+Pt7rw67sDQzq7kfEnJ6ZRnGSj2woV/3G/thmsNz6YP8kJ
UQbBrO6n7SBnGNn6wK7mC35Ry9vy+hWiF0w5z//tAYQY+ksTyGIu/LdES+JXDKT0
U8XLkyus6SKCHBo6VTxZZxrRBEm63Z3JpZoK7obQ3W0Vpjt4dJZl6JG2xYcN8apA
3S88+NWHlMDqeZ55x/xKzsrU6PjBiJD7xNnvndB1GTD09lp8XNCnToJlho9tr1IP
pC7HVmNy2c/F3nX3U0Sae+ET+0Zny0Y8XNXCwOEgjH/3fkFs299nMODsLkew5QiB
BXFnKvpoErKr4m8Rwo3DB0edP6ZtGB7pRhIk1HZG6k0EqNjQTK6LntArjWD6Qb0i
2jq1xwUo4GSusBUxfg5f8fsegWB/kRU2auuaaHJhkYHTDVgRXcF7G8WMmKaWg7ur
X5akPT5frvslLRBiDIRZjbfdZ22VSrpdJA6WKH+yD+ragJmYCawt3w2tsotl3+Bd
5CazgYZ5m8AWfWfnHDVfcalHuQWMahR/rNvmhg/o0CmENcNMegyRwPtQoTbRNfCI
4fXthCC8QZwASSJVuX++KkoXjMG+HUC61U8tfjys3dM5WwUF0bomu+Z0wc4tG8uR
fxRuVAeKsxVVbcy+lMH4/fvB1oKlTBe3uBg1f6w0bqNTJQ4GLMAbDs5qq8mFkosz
Hj4f5GKbLk31NMOFoSg8lNtVqfsmQLk5EQ2RVm+QyGibujKkHwM51tR5fMCSiymo
xFeWxOUWY4141fmYleCivbJCHppWVIDAUuC9lzrpTKGPnCcJnyVcWkOszxW1Qj/a
ed2UbPLHRgofjKlfhCUC03HqInXIrVqE69CXEi2TTxYGhyOdOy5XN3h2xkQ9XkW0
8wFDtXARuNy4i/UD0lDWaGUUDU4T0yHMbJiDe7otMpJG4FxV3hCCPBlux4+rgx3M
LiUCYzRgCgvhnf3wsG58LoUWBW2LDxTKYquiaK7kDsqTR3tsnk2B7sVubq5lpu4g
qnGRTS2Jx1LqmRHs72neu7XXy5IbqpVn9YC8RFGNK5sDmKyh/eYvq52xJJdaeWJI
Ucf5vi5RJok/nFQbwr3dhdP9qPZ8na/IzCMIqembQn1lEZ5TK0B8M+TehnOeb//a
vxV5vR7OYHa9OuCP9IzH0IImKYw4CqzddKsnRFEeJan1eF3OW6a6kBO8kJs5fXBE
RwbKCqDCWHWeZQprORQl85GsHPFvX8ListWenB98juWzqVAEOAKxZB6I4hBxKo8A
9VlhUFlbmCNAygjlXtrkaooY25cJeY6FC7yA0R1aQKWK0Ko1ztD8qW+h04vF6/NY
YnNi3XP2qiwNKpr0WI7DGx4YHtD6q/jzagWKQvOK1MYEtT64cT5r0MHgX2vLlcBl
Lhv4Or0M3dn3Xk0WfR41tle72aM/LSaA0oRYkrcnYNtmoLbwcDGFvT+v6wy06kRq
0m0lTdVjyQjoZL/+MkWGpPKfjNLvRpb89QYSOE83/7yLtNCBTtRKVt59CBRe0Z3K
5jlybfLAXknihmohLPt+jY3BbIi+8Gf9AZ37RT3iGVpJxsUnd+SIG9dptBqDWmY6
jUXd+ZQ+5Er3a9e6n+j2AxAriwwiBabjs7ra+jgj4y50bdvMR1b2Cr81Eyrye0aD
3/ABObVBsIIAycZTVizOj2TaUe+qr+AoVRugAso65hrAKcUi4NExVhoPj8ZknUYj
WdnW3Ze1MOPw2YGGge2Q5lm8onWcXvXmCpRAWJd9iOKZtpMtTx58Cq8wDf78hJWW
kDTSEmHw3hc/GJZRDj9J5GOvK/mYr6atrXFsR8U52ybxiq9ekMakFWqdE0CjGg6G
ntfS60ajS2fNe5jgSI02qvThsU6xxe2+ABKE56RX/caz5R3ogoHjD6ac8f57U3Ol
yt7UncE3/iCcondT+GgM5yo6MoqVW9VRCCAl48DUMA1gpurqpV0ycSrf4DZMfDNO
+nJVoaSlabuSvs6cehW/oussOuJ40V7Rf1UpMdjsyo0ucGo+0HCatunbAfNligSX
7Dkqa8xQiIYAvFrzf3lkS5WFkST38WYxEc9PERPMx00vnTSk+j/5IYHY4441i5ys
BcmmLqHLisEU0wXMptdGtLn99uPbb9QalfYKg4k5AJ9w3uBUOepFVuJ/CUG8zsg1
h45+yVAoBnK9qFtEEmAtANCepxJSiZLudgYYsmqAaM1M/kICQpqzSzQEj5kIDdBl
scf0dUSZ9ZClZbm9Fe5LTh2nV4v5PauOUszMobE3KE1Iz7Y3lABjSK5sqaXXRU3a
DI9uchQjwXRp62mlBebYP0vwNLGVaysBKTahjfM/j4vO7s7So/a2cDRByI9pbXSy
flgwl1sgum1JSpIveBPgY1XPRjxDObCVcJhnErQJtE2o5iZp8r/sx871Cui2L6PF
rNowE3IzTeHg2c/b9MUoJRUcvuFsB4KS/rlB9uR0C8q7WijjYbZtbDSHlw+FieAi
LBbkvyOwpuNwO+wsejOQ1Ei0IYQthZZQTsmrmJD6ddoskRMgahyuytwYY8fq8Okp
oNBAp/g/P/H/dHKh2XFoL0076IjNB1xoKvfaoiViObZyFxY59A/yMesYu/AW0awX
dXtGX4lZaqae1JJub9XCbDw1gIji9ckKSJeH6MfQVratPoIPyXfb4oLi8DnSLwua
O+Srgg1olnIINCEvee2D2sIHtpFYEEwDkw3qBBOIJ3cq7tAo7Mua6plh3Ipfocel
UIRh5cNIleMm2GJr3r9+NvOQNnC61sABL3MoAXkz/r1AeQxaQfVoCqD8X2kl2Mft
TEY6HkC/iyCn0lWionTR95XS3xzgedue08HTsltm3o5lBhb+ZPtkIceW7/315jN8
AK0sO97wVWcESDOIzEOfnSNMFyvImAA4Gw5+7Gcpz6WpXCdOhoF5g24wiO/8yeII
b3PFzMrgkzhAk2rjeMSApvVQ83QbYXz9m7qAgz1CVYwLGlP7CzoOGibd+pQnfKLW
bH0xLeAVoMwS/2zJj8odScK7UvCgn+r/gjeTqwDg3rurgZqoreV1qFx+HW4O392r
3z7Px+IEq1hvznkw6rPx9+Ff1MOwjpFtASa/I66Zm1ByIxEN91KolKdoPr9QpiVR
UX4WV1mCUDpVEyNNrRdDdeffp7HrOdbi6Og81xFNPJnPCjp15FJ8DikhZR7XGu8Y
j4B/kAm3X4aPAIFtJ5Zj+lOt9sP7MY4La1CT/DAdTxgORcH24k/mBYqNeENGxydJ
hG7GJIs+zAzwjR0wkQe7W8W/bn9bwotG9U5yM+IHYd+sdx7WOjbt1Rl6E9tIs2X3
SG2mWuQIFnmj5YeMJLNHjyTaLSIL5a/J/8XqKQ1feIuHyo28UBXrXINkRxFsOCt2
wq6KF9szISnTcgX02gNxscIO2BnfpZQ0faLCgOwTt/Lfb/zDoeHJM7pgQQCpCDMF
IA2d/T+KIw10Cphc7rQzn/7ozdsfxRRypj1iC2J4p+Nx0Yu4FAMtOJagHHlsiwkf
HFMshBlQkP5P/Ks1iUnzbH0+iLM22XWRh8qQSO+Nw+MAwbgvsiFMNcFoTqTip4Ra
oBuD/7L+ApLkfIVBrggFeDU3Vs7FwQQQuKM444lz0oHI+k9NKwWqjCgsVJEPLoLU
q64JZ//YXPiIWS+04IgDvYWNdjXF7TmAvVo1BXa3tRzYfkervG1kh+i6eUnQn+O5
OHwf4mOYiTGklINjtB+Y6wNWVY60S4Od7dmdVqhLgdo3nmA8LKYdpKHataOEVuJh
sVrbZvYIM6Uctkm2pmNjF6rtL+/V5DErCnXUiEGrTM8aXieqPagYm9y3Tz3q6x0k
oewXf80P0nmcqBsvTCpfAwgLAIps+2MrHmv+zmcED7y+IFLUpfOY78oRx/6KhqOC
sDjHaMtIsKTK0eaaPp3VGJ3BkZv8js6L55eXK55B4IA5RjP35x/Aj/hxpVB2YncG
FkbZles3J05fQHIJFJ1Jr3YcwHXK71gcmb9iOZLmj6C9K0+5NxPWd7b8VQMbOM8K
mQu8ut+Y3bIdf1VsP4FlhJUCOHeFxKvdK7riSn5J9tsTvh4RK0oXLGRFt/fdnJqm
xjAwuIF5UXEtf5RGZhDwQSIoNcmKOdvlQhV71ArsbM4JvZWU7L8QHcbEJdZnaONS
7J4TTsJyxgX4ccCVhTLsgcqwqfV765QsTz2IyORqo0PDuJINxQ2kzFDeECcg5Wgn
xdOuyDvf2YT7dYSxPz8Kn3WVVa7kJ9LSy8gxqmlAIP5Cn/FQu3WARCuPx55HbS5U
IDfAlct1Thv8Nj7oPS1lV1Ouwv6tLezgLXLryIUJisTVI/XXg23wLPP7hJp3SDuS
iXWIXBjqImBbwpK9+zI8VW8RSmz94ZSlK6Mix+E1ljcyjBfGmMnQpQe+m+D3Syt9
8ll+yGqMbJeR0zpc4T9V00rtFvhjeIXkRpHakj5qpvX/QH7DxFszZuvL+IZUIcSp
L/w2rJfKnngs435YvMteFCuF4MHut7yfPWjskTETmmGr5h0+FctpweKQIb7t1Dl7
6cB7Z69rwdHmO5Y4lGDFRYP/r2KTj4V4rqhnlAw6ueUFM2Z6CAxEqhhYQ70XuihE
EP1PFtt5wxbDs1ArkOkEqOqbvjAyva0odcG5jf0EbASQWcPxYyszCwwJ3qBAUOcm
gyBGX+TWqB+gKCy8bTW/WwTrVEgHYfYS1ucn45Dce9cB5nOzHELUMOK5jmYX9WI5
/mALB4BGe76Z2d2qkJ/01QERaLuc169cDrwGcA9lED5GxkvvNmLCDOVhGONbxFmP
COJ0pa8J3VP/TFTsUOmZlCGAF//bM+HSwX1YbDGL3r5G43bERR9YhWJ/7Bb8VDOy
q1eJnnKw8sN/8iuMn4ZTpuK4hrid2VmcU+jDRYuQahR2AgRM6t68A4vzfQJhKrgR
sGYy6tBJxJSqbbfpDQPIh5HNy82Ox3JITqr92+ubDAcel4TdP68jxEcC/mSH4jKH
nRZ8LiMlHtRVKGC18eMoQ8beCT5b09neEJFqOQC50+AkDX9JesDojBAwH5jR4GIb
A0raBvvqQAl4GiSBDaKF0TRFeUL9pveiaCGfYyQke3E6qEUplTmrR4/JUc0OMiQt
JfE6cwl0mW/IY4a9b73ct6+3jfiyWOrpMBvS1UBLxouKbABAoedPNPwt72dMrpuA
nmITeWSz56jbOsvF4/YMHsEkWS8g2pzWFEFX9J0rW7wL56SzPZCMbg4rX03cxtKP
CK9gTDlauIevzz7b+IjMqrsTNO0HPXfjwbBjZPIOWdoRMSF8h/6KE28J6VnF5L38
xQKX4sT4RcxSYBdQ1Vs8CWapS5RT1UVvRoqf/F7VgPtiXHrw1PruIPCsMFpXdKb/
gUAfcT93lt9C+50Ikdy++Ozusx+123B0C55d5EY8CDeTtELvWnvgB9JW/RySayPB
4X4427f4z7C2bSamgxe+7ADxcpNQWLIdTgGfiHvGG+HlgOn0bvhR1WQKajbmfPmI
pKbDurgTY7nLEAgJywIEoxWqnKsZcB/UYASbY4QQFn+T/iL/5PNpcGOw6L5l54wj
k7YD6+ccuh2FDwcO8VTLtS92lO92wdG31DYyZKQBYLBPI4eWjEv8HI3zKhLaQEAm
ZWjZN/AdrFYVSuIstvhhmkfPbAnQW9fCintkCSJ32SdtqIQaRVaJnXH44yD5vnQz
7cUkLIH4Wnv3YaU1a7+q/QbpYk6jivVD/9VwGZcnxVwXI/RFj6Jhsb38X4dGBI5z
XyUVK7cKY1KTZkWFv+Lsg9CGnJLjXF7oJpvxnsUcc62+/fDjyPbO9gJzZ/8k43D5
HlPwema1qOFT25U6gxOT91/kyJcs5haUliMZTkszi7BCFUQZkD7ffEqlnxvkLQpH
Or3Bchx2XAxZ0D31Wr1ZeS+qBJeyzgRg1SJ/GDNtH1hCYdSVY/LLpY+rZ85ypj8P
lFuDoAQzgrvKVniqKOBq40oIac/RvFEk/JP9fHcjdFMtGh2Vb7kGqMs67kIl7W5q
xCjttnG9d4b0np9SJMnCbcP1NGAWh8GfGMKLvotlhcTlQeM4B9F8Zp7vIPJzbIK3
s/g8ubBsZEcyzOy4E0ueEaxX7XXUsE58KoIHoHuLAZRjGXwGDFspshLg6ZFxEJS5
P/Ij18OH+fO2ezv8X1mh7TR8+7dPN8sH4qhDLaB9utbhC5rmDvaNwmDXtqNcHu1W
rP+wZqw3eAv7YXMI0uFJRQkU2ht51Ff9ck2admtO+3IVA7HzdFP5R+CzXu5Hlye3
27eHud6ylt7MXu2HfRojXSByGQvBbbicF3W36m3oiosfjZHH3ZYgyCaWkOQnX3ky
Q+xgTLfII4EHMFMoPNVcITKJeGI/cT7IXzVS+vebsd9+hbLn5aPhwP6Tu4et6q0w
+NzxNj2IqZLCR6NwOu+qXURjfeOuvijwJtAUnznugamBGwZKB0nVD/QoyWFB9buS
/ipEVVmQHQVJUHyhNAUv+PmsbB910WoKfFCXakkM/t1PieA1EFXVlvb20+pHx/2v
6xIdeVG0ww1tqNNiQvdMzNW2wFZ4VeTayqNjs+R3I7XPeJBrzcZk/U7mutYuwNoZ
ulQhdPZ1cru4TbAgsVEr3WWZGDYJh4ac7t7fbvOoHe1rNrD+ZpJ3PXqlCZn6VWYa
MWNvpB8tKQ/J88P0YjnhlgHRsQe53LzulH5vrNKBX2zBBO/V3B+eB8jXRaJus8py
KHGjeYqhjD5ZQz00/8+k8ZDQhmBP22BTV0Lg63jNRmtD+P4gklC5/zd78M4JYgnt
X5Lhc1fKdKA3445PQFNrCVqEy+Xeg2GuKJCdd+6RND4fxAoTyNvnBohBIUx02ppD
XVyi8jgsIojiuXn1S5tx2vvDudlP7LWq3tX8JfPyV3O8HiBlqSd1aBMMBENG2mkE
zIrrzP9oecFcq+O99/DXhZu+jzdyNiUPUj6kUw/BoNnKjfwkAaCVaQEjJtnZ2Gu/
TPgRqM+0efZ+EPiC16B/sernzB/Z+Kr/b1NtqEdzkUrNjkhZe1YMD612l6gQZpLx
mmtpDLYsM4/aNzIfvdPGC2rTLp/sgV0COIU+uFtPzmtddBwgSISyA6e1o25rS2g+
F4us+4fVlPp3h4u64QLdHfLuxh1XQqas3kx1wiU3M3YTmXDzewVwmAQ0xkLafbha
PoktHmhiJUmxEIRSH5s7WZ6NEakpGYlxeBG+KYpLVYNBvN+2c3X9zYqz7mMmP4B3
Wsev0mGf6M99rF3WMe/Z5VlUxQn9psaK9p7UP24764ghBpMKpQ+MlWnX0hxr2NQE
pp2O8m0n6qPVNMk7vjgBbhBtpyoWaKwkXKw9DjMjSOjOJJI2WdbwNiSCdkwc0bur
NUhw2iPoZiYuRNykybjZLQ5Uh2sLi0XN2AlImZnb/v4cb0piEuP4Z2NF8oh1koD5
vBXJcViPT2UUojWmrTmA18BL3UEbNYlJBQDKBk+NR2JwrAG+3WnvsqjFPFTdW1mr
WIwH+tXKgjYef/Xn+B3CSbH3eRdM9CnVg+0IPoAj1viCNBDGEZTAiCUgXZ+7rg2I
SnTFPh+I8e9DaIiphmVNpeuRMc8O1Hw8K8o4Jjs7NitfbPGmMZIbbfJYyfyHzSTM
OoxW6l+/GtpdCgiHzxaCMSWE/JDNJhrViVWu6HprPQdB61mas9Bx7Ouw3LFty+Y0
XWplbguYbcJUvUPD40ixA32Kx84m9eIxwl9Zw+VbQG/Qmf3wMhW3oMteDywgQfTb
dubza22X16MMfLg/GzckyPLSWti5MsVr/eDfxdfouWV3n1WXQ85jBqIKMPyEehTt
BzUcHQd08jcfypsQGJ2pMvNnMdbfllJ67/75J1l5EQ9eXI40BcLTGR3ZeFaqUe0L
0LMVZBnLDajFiUF4OyZlymNEWHkLVeKFjptjvLp25UyEfcmt5VOlsFOsy6jdItkU
L/eX26uIqVnSDaU2MoaJd6rzUUMTdTCgmJMw2XPsrXcm/sACaowpmF9V46aDy+pQ
yr2qFUxi2oe5AFsOBCltWFE0dUav6ozr+ueGA61rpCIjiXF5Wt+2ClJ2TN6qrIA9
HpPNBHzkWvq21rnljIyBcewJSqDx3ZRTWhLO5+D0BUaq48Q1UGUBFkGwWHTxMnn3
1KDD3iuax2X0MGEH5QVg5VcpQYd7hAVLJx3wz0TISGSU7b0EDaxxv67DGTOEUDN9
N8JL1Tad3OrjFQkgzjsyNwqQPZXgMde7nciFD4OLvXa0vl9CrpNndZEBiKzolOKa
zWa9pgL2zYE9p4yARzFmS/CHU+lWyndqfx80Ml88n+HyKDlg2YimE+hpesVF0cWJ
cFKNw0SxRqi6ZxyJNghpF1Bagwld/V3zwwuiunZ3/LbaOsFct96+pxXrdFKDSRt9
EvqLUa5Hpxii/RsOp5q0Zwj1gT5jWqsicW1n7VZkMdJ5MjCvK4BafKD0CHKl94cI
w1mbIhXuhLGtyJWWyGVypWn+mZnKBX7/a/fR0/4OO819MNuCoKkxZ7L2lgm5iWds
MA8oGkmMDQxuMTaZ9fOWt9wk9+VjV5j8bpbjim7Rnn8bMA/uTn6TdubHee6QNzPS
/UYNX1hr3vKai7MNursKn6tBqOITpjZaVxAIDVZiGiXry3csMu8V2WQ7FWP4MVoG
s+IMyg18d6KOvoM4tnBxjlLgRJc3HfJ6VNeAP14R3rI/WM22ZZ+8+Xv0GdBNNgfu
l5bj5vExqTHWN0FZdM6Kt6yNoS3+25jkV45NK0YB4dG0nYK+6FUNOfxyjFYLetHD
n/LOiCPfPgZK02OGM+p42bVo3eFqo6n72/TEoX7879s8CXe+HBM7NBj2v02SUap3
7C7EkNwwKkOnkpbsv+hHO8fa8HTFFKTmi9uJhNX8RozYAyICQFSY1TH/UJYBaTy5
C5FZcC/Q3x36VWffScPXzep+Kz+dpvbVOC8ra9kGgfTI473VzJJEigBtMyGV3HXI
hTcFfJ1H4ddBaAt1SFhLMJVZvQnNLCU0iMETVe57/D8as/1IXpQkT/6dvT/l6/Ar
S+JFsJstiKIdJQPtegGLV4iDc2cVL+kkA9Em0ZL7iieG43siJOCEKfT+XnV0kS/+
8DtjnTQ/UIfV4ZLUoqebMvTyc9fzOSF/pIyWXI1RPBbTPleKN7P05Huj6SD2yN7a
zbRzGL7w1wjKWfGtjmq0deJlHQXpSXeA8iEOIUsmxOxaB/nlFTw8sk5IoDdory4d
zPgZUAp5+zP9bq33mryPangLdo024iJ4lh5jD8f7XU7384zC6t+G7vNfifhUrAx1
uI5tMqujPEtLDVIVkmV9ljNiURa8nQSW95yNcBSEXHq29K6+zslbLabbK+yDcbkg
EUkQ7dZqt9S57WZ+1NgDm5wjd3aRGaBWjAzC7YY2HTKV4gZzM8Jm2wEJ2gWSM08Q
cnFw3eT7aBDs3w1354Vczdxy38QtC7pCqWCm5T1XQaX6WzjcripVmzflhoWxyyHj
7w7HS7MQp9gTc70Kuutjn8MS8c9rFn2Qkf9lIapxyg2o5jMRWYPYVcP4S53Pa1sO
claHMpsHnyS8ofuQXdNiuzT+xvqKc3Ckc/Qmkk+HN95RxurvtGGe9OAqCB7YZYI5
yrawz395K91BUjOPp0cMI3USMg+YwbhlThgaI7mMZ4UBbI+mODH9nLrovXALcOtU
yH27g0CajP0zdvX32LEK0Ds7Ef+itV7Tx0TTuXdG1z914yWE36/+RKYT+B2Jsv2J
iYuduW9rf80ACojAjmUR+WtLWPK63WrkS8d2Sdg8QG0CHK28pcXo0mGp2RlYarhe
W97GWaTvMBIU9DLNwOYDJKUahpx6dChP6N92F7msJsdl1IXlii9NT9UkeRGQ2iuS
JgFR2TXOPiYkmavp0V7sRy5I3H0CzvCoHy7vKQCfP004nFea1m/EUipsDK+tpPMQ
kqY9B21f+zSyDWezteOjbubG6yMC7A5Rqk0sSeQZi8l2g/bqFN7Jt3pjiGk5Gc3u
kxVEmOlD+ghX4499CuokddAsLS65IfeiV+jmzI2M8Yg0koYeYeFOE45cBtBGyHJE
SQHvEKM+f9aug7/D+V8cCiDgrSlsJC6mOEJaMehwS4cdrg8+DyqhoGPMPlXJt7hf
KQO8kxCMtbLx2KeIylKu3y7zUTaPKtfzOdzviCH9tOgiqjaZBmdJXWFVORra8RUL
6O/bkHwm/RjviTJOgYRAgXukXoanYNp33ElLEp+Ol8bd52kD2PhLS9KEeHJ2PVzI
loxa30bvIFKhe33Spj2uwFXJ2duylzrXYpcdfGCmGbCr9zgjcexPSjGU50HMLu/Q
s39meiXYakGf6ZenxaPB42AOpm304MGcm8v6qpIaRJ18mHUAaVFyfPDiB+Yp3yJT
dqjYNP5G3la/zqQc/K4x0ErwhEjz1f0KAWltlCjfT46KJT4m0ZpULcL0jOdZPV/+
2C0jjHE//7VtQ/uU0J6/hYU2f9NMhJk8Y93TJGjZJ4LXcsVYKL6cU3/z9gJo3S9s
wL8ES24I8Vej32l2sXF++nOYPZt7T680A+QceXgoX+FyE7pnO5Q8KhRkFfEH6Xcf
ZLZYzm3rPHM3+HexR8RFN9TFYCZROQK/MeI+NfAvwCENt8bLGZrgs4Xq/j5/y7Pe
o3Th5ZAdLVjxbCUnS2+4kAPPvU4uqTnV1Xqozhf/WoXaSAJXaDGlB7onHfM2nWOE
etc8DW0aDnIdfQojqfSzDecyGHZHlZjtncX1ShYVu53pdbTfRGgGnRjd89jwuYSG
lHvIbBvlVf5pBEFqIxve6pgKbr61dw/vc0jJE+/kFHsWUqygDDIUAYTlWSFSQYzt
ZQILxRp70QoQbNFRbAEElAEMLLzL0+THz9SnXGzi56Q1lWrJwHMqS93uysvEabJ+
jLh7UA+zrYvExzZ216+iJsyKf37vlbmULLUrEfmtRUnCWmfsK1fclrOBqGHCipcz
6m40MFwE2ToytYRF6husDneLXRgVYgvAGHnKdK27aHl8emoYZAKIWUiPttpU7YFb
m0xd/oDEG2lR9udrsui2gLbuzemvXQJcbqoVoJreH79EFiZKKGqJgD11ysflq+RH
oRtHr8TiD5w1/6x0E4q7cvz7b7d2vNxZc8gSaMRgfzeudDuQZjEgA+3Fks064v21
GWAsgl78KPZE7EJjX5xgVTb+WP5W2t42mBKi5SPNUO23nMc2qEWKAh0UToVfSqQT
tNpLRANfEWXkwFwzLTSg8StaDl65k2BegjAnXWUl5VFQPKo3PobTsQLU8z1G3QKu
cB/CYVTZPKRZm+Fn4VDwu6BbhTifY6AB5VS0VZCUl/c+eEqk5ekMcMKULFLAP7GD
nJiJVQAduu7iG67GtW8y8UMS3HzfNc6J1a1/bFalQ7CH/m6F6jVHHNTAQoU2lOXQ
Y0Yn+2tLqa5lqMKOPTAtOqCUN4i/lEQY6qOxFup6GMLTjcW8FT72MVOxnfKNqZZ5
VZhPJ5DdhYr8Az/6+ZTtVpP8EJcQQIGpyPHVsnuvhYOYiFXSdFPjUD48s03dZafW
QJ3Sy1ZbMUIC8uxI5E4sqX8WAtubDiW58YBJ3cxHZc0JzRc/je8wlET8tQKbixzk
4YUWTrVBAlI02k7b7TJ+Sp2QbtWCiznZ3NUGGk0kzJ7ttRmbcGWMdqPDVKEzyE3z
oh8F8c0vpiCKUy3o31+ut5QpDUHMNvlLk2U5dg5lAVk1aVW2iu/0I5ZKqayGIrSm
VbWP9IE8pNxY2NES6/oX5Xowry3HfZ+SQmXPDlP1s3VnoZhv+Sz81AODHCGrykb/
DwyD5M73OkGY+oDS434WZWJxoW9vnyXYPLdCKm99guoSg4sMhkB3jJGSQB+si+6d
LuNLjUbmW2hv5ULfocTc0YTy1FfnuO+0K85X2f5d86yvkxfZbMW9RNwKK1+UntvF
se2Ee5TWZDzHNe/glmgm43Fe8AHYqOL3l6cM7DsHq3NZGMflurI/rqhPTtPa97zI
ZMaKnhaTP0W28NCKlJDJUv71PW+Ezq7dSRij8/q2xoF2U0OlR4M60vKf55pY6/7N
9iED4pehfYWqx6sbQvxF3PRikMHjDfrq/BHALlORsNTiaSlXhqIre9p4MSWocqOe
bqERj6mNg2A9S3ULOKG5PajwHBmpNLggiveXinGkob/JkK3nibxLP9DY8NaH4+nf
cHar+LRucCnUo2BKcLOekwnlU7601ZD9K9Ik5tguydTgW0Y7QqJqdNaBLJu4X6au
PJS0kG95MhJVyy+sPJGE/iha2yQ6dGHZZ2N2IEfnegtFAnPfHY08pBKCcKJ+7M4y
pEbeW+TBnIMgth1yAQnXIYt2XsJe2cjWwbuqoRH8UPuijAiKANajbSwWxib3vtuY
7PA//qFZPwZrZo7U8Ioo4SKIxIzmh7nRP/pa5IgwrFW4gVIwe5ogxs9yNgkAr+AO
Xdtc5T39CQ4Lkjzzr62vVJ8eJY6Efjtylg5Dc40BOZfoCmnZ31yETrjKu6Oy6DD2
m1qX2M2OxYtAo4RlvYi+dwXFD23ubAfnACoMDSZoBnzr+cZVj8TcS8Rzb1vNX7CR
Vnx1rgRohremHqIH7/81OyNefgQ+MiRxkZdcDBt6QuSvYlCdEHwza3rZL475noaF
zdvWc4xE1GLSQeVwhzOQ4JMxZySloFqo9XMUFzfyT7iBr2dH5aive8wJfj6Ww778
O7JWG5qJMHsZZIFI+cUvYacipGxrlSMUpjKVBT1i3Te4z6PRwnyidTNadS7eXvAJ
A8EHBMY7geyhBwww9nyPBvtxBPAG2nPw+ZqfYCtXKYzKI+lWS+yOSn1g8z+sQB1L
mkiL34T5hwDNm5dYHnlI3l/wDWf6dp96I9+syYMEkMpihxDy1JQzzKnOtONdUbjZ
ZbKgVShwW+mhKzfXYYsxvOg2gMAYm6aFaECVDENqP20XarzXChUk1G16IASCNVzq
d8aDQwEfhftJErqElfgW67p/hFSkiuDQbTz5CccsZnl4QTPJSNUyjJ0kpLM3rDgV
7f7R+c6Eh5F9qEsvxdRS6n806wNWvXuanunrLVOJob4VowQmHfo3MiVLxjD1Bttd
Kuj78RKB7H80FAWID1DEZ+cWPFZ5WKrchiZMldaprg3HCn6LP0ynlcN2FNuXtJBM
d/SKa3D86JOJZkaJ0RQssCFqb/rDRsAe3ZQDJJ2nmiU1RlG5p9ZPu95sTKsqMc2h
W5fkikhvUpmwRqgiUxUn+DIV3sM+xNaXukmSsDZ1Ak/euoM4bAPy+/0Gw05Sgyc9
3q0G6d7xd5jue5S4ZmbaDKhcCP41sJMQ2Pk6g+Fs+Df9g0PKCwQSQQ/f7gX68nbc
ow6+hSwakmxLsG5BmhdahnKk37zYYgBwvk5iUJSt4P/exXwup1aiecntrhzTxnuP
z1A1ZnaTyFGsx23VwcT/9d4hgQXN4/FPLHtQZK7S8c64v8mLvyuTEAFOPpnYXlF0
0j9g166+riEqlXsDuC2U9qTSDu9H3LjG44VT/I3HcXmVxCEMuucuIIn4OiVFJ8fE
MfXhuWNgAlnOBz8qtx3bPV3eAAGOobirUsz1bKO7Y8y6ftBRfwbzkxm89AOpsDgQ
aVYay036eA7r6WDKEOirtxRn7RrpMTSaScP27kcLTRr4+wR7IykM7QuhhHIgtzWG
CvhlQxlD1YUBXFh7BEhXi63d2U28ut3DT/Vl1zdkCxAl/jBx6z//GiZ3W0sTJN72
pAnWOgDRtM98nB4YsKCUDX2YdAMvUUsFrMW0Ej4yDz0eQBIi5jDuSGn42ka9knx7
8yU3OHZYDlw0dsVwLJiqaX0CyOooH/CzgtVfNJk5OXxB3fWO/6xV0lvcm06VMlEG
EgyoTM3t6d8bsOK5cxY+yOr8ECspyZYHKmBh89mSmNx0Sva8b4/AHWxA4f05did7
OLqAfO27C+uS3UczTU84zSdf5DNhhEulfvJYVpuH3PWCf/pN/1Xn3rFl8NxW8mWl
7sf7CkmOanAL0Qeb6xRb68rVZlgeNeTR+1yiz2FNdQyAIlpkGkjpUlUDLl9iMGs2
NVqUKB6kLO9bc45h3MoJeBXtQmvjHX/lbIjc+sNk5oA8zDTLdHY8APtVMqVUR3lK
ZyMQzsBva0b+BKKTgNptS50tQiE/Wcd5bFoC5SAQt6Oab8/oZixNUkll4+D/8mtd
qA35at/2VTA99acue1ic2bkZVhfi0w2vyv+bZtX/mZp/UTsFDEKr6v40xs2UEYzr
SAdY9hmNnWjgeBsKsG1O8z/Ys4BFN2ynieYU2RFn00tqHJCaTA6YPSZNiOs93tjr
xubQCzLmzqiqfBs5WqJ4NH7dSDlOgfybfCur8pnclRBPimGE1O1WTr06JD/RViGm
g2X6S6mrNiiziLjZjniI4IR2ZL6ARwyA7FvPq3rKJCqrKREz6BkkE48kNaq5wu/s
j996i3ctgaIqT3lZ/wkvFntRSkhtLI8KaNzwmL8ymZRIYMFU/8dNT22+bqkUJscz
kmfDNBLv4KxiXY05YH/VPRvaVf15oB4poOfGvt/EzvSv4vRw88nTukPcmaUjqshb
UXvk/sPzplSgccBwpbdDnBbrHbmSi0vacjx7OgpsEfoRhSJg02cpPNIOED+RLkFk
oMklyv56ag/gKnK9GV8v6IkgPK2BEQVkE1ZmPl4AC/L8oSh0aZNiSuln9owNAvLE
5JoOWKmqzyQljKAv8JW2fYMeqPHrBLmtl/xcZkzBFiYNysl8tUbiFkC1UQWhLBbs
PNqFPNL5Kov44rtDJCYFsDctMadcUZrIZhJ6afc+phvMet1YpHabdReQCw9IM9Iw
tizMyXevRh2ouiD3C6GGgXAx3yUn3gXU3lN6q6GuJXYtYrgPjtJip7C5kTH7KRRO
giFafK656sv7LYQcdQwXNY7LPh7pcdupSgpNCzIRRQ7Mx1jexE1SiqgLtm6lW0WO
Z7GgVi9CCdxCGhsF44qdK3XsCECozwh/cXNknnYQjl0nVTOvsnVHRuGalYKVkEHz
1sqtBYZdYXaD8oJ23hdef1wphSZSeWjklcfbEfA7Zzy7b9sby0vKG1RRCKp/2+og
B7TdtGMcLza+avRBF8Ma2g5q604Yu4r5+1ChgSyl+OGav21O3N6yiL8AHx7lfys6
wIvNsUkjTRUO4DHlfsgEYYx4axh4KqZzxsrWyYynbhi/ustF0NaeWsA+KukVQwPJ
sCXNssSwSHF69EWaeCAv8OmGnyXsrErnNbNCEcGDO7RESRmiKm/ulNbWrhht33P1
SHyahUov8bq59UWIerOiLjPxF2yJSSVfe36p12TSfi/umTXX8HrnSWF5PlYwg2zl
pB1exSYi/RbfhaRxuApLABywRZ0hfQwMxP1tmU0cxYDOLFyENqWljXPB1DBhPI+F
B7sCR0UbHRRG9CAsYJiYt8z001fEf7nQ7qYUW1jDb1ROxOThHV5rMJgr1iCNpJyZ
f58RQ+GZWvntla4pLCkgUfZUW7Dx5IqxtMFqDr1yz1dsvyMhmCF+hsNKVeD9NjFn
QVdw2Mk8xGFKJnRiGExmL7F1O7TJSujWFwK43/5JCSWYaQMpWQpvTygIn2PHMaG/
nLaSyYyvGKvT0kSytjs/AUsa5Xl56xLtdPdilAyT8kw+arR84rG2INOwlsvrJ71r
+mrAcoeXzl3U4HyKxbeNF7mj5Ki03HKP1SAB6inHpUGWyGM1bcDiOHOAbkOZReiK
0IF6gi5p8CcGZ4heD4WCZyqO7ka8EYUHBxx5Tfwv1aqiCR+L91Oz6qs0bVSJJQSm
cYDFILxcrRlsvK51ty21FIJTZCIVpgXJDor6YJlA5czxTWol9ITzILgoTbImx8zp
C/r4WQewG72Hu1mExkinaU27wmTJ/hBZZsbvLJZXN77GQQxDwc/II6BBwpR2HbWw
zH7V8IQplo577VrRNM5Ju6j8eHObgbUho/YlXHOBhncduDS5G881lf3dgsoFtaJe
UYzv1MGF1P4gab1pObEuk1TwbYqD0Y73QT27U27os6UGpAHhPG35M2CAhPweZ8N+
y6bTBa6rn2cUMaHVrhtN+IKvkj7LLkdPa+/jqJAMyhlOCDi3+9OMW4//5HZyF9Wb
zMhiOwb86FrZvR4HLE7JcAtH5AsxYlhu5QOFcB5EBIkmaS+YqWPXhs9J2cE75dDL
K/3JmXt1zPUfiB0eULWfJPhRRwp7g7lQn3kmLEpiLCTK3AarndfS5yZATi6wx3K+
iVthvEpbtWGCOJzCTNRiE4swzyZ6LsmGyGYhWdvyHTaIh+2H3p0XAyVAbuZEOB4j
WuCJXxqCIwv/dqlrnKLc4ihXY41thdPjOXhaEL0Ke7Q17JdJfdKAFgYHf2xJIqG5
YILN7ZmxM+SLbuu5hb3Os+kgKnvV6dBJfEKcqzGuMXC7DRkyQVlPlL6o4Hhdzv6x
oCtTGSWyE3P6xqCbNi1Ju0ovlUDxmc1ImrOzqCD/NXS/u9yZ23jrC02Ln09LI1PC
sOfZjXuA/6vpmnWsrMzjbs0S2z0fEaNSUeMfwcAr8XkyqoOaRHKpBgsF/jQeBm95
KJZ52ulLcv5x346cEMVIxjsN0nTip0zo/F1wtAE6vZS+yNAaJgmdTCMbW3ZQZtDe
8qQuTEGr7XITw5z2vWO9PWjlWsvnheAWmkS0Lq4VgPBFf5AXxrInp5QvMkLPWtEY
VxUIc1YDzDf16U0sl8l4SGWenyXdiF/7/ia22ZhRFF7raEpmKMldKzb+TE+UfxwF
SHLfvh4jpv7b7UQuIU94W7ZEyLhfH1c7szNwYto6JEnBjqH1K+5qvQbHs17v4cBM
U3EVCw5cV6Ci3oyo2ySPqehjbmdVhlQUKIcP/Gfv4NK7iCTY4paZsLafnaetp4ai
0cD4oF+FWOC1BVOuts2jBnYYL8msN268RS8384Ydx6xiuGjAPo9webwtlixrAjBl
7fbLcwJpHIMYjDUiKb+exVRZEAnBjKpNmvh87XXd/jxXgRmgLVMHrDaSgAiZbo72
8Zn2fGkduBBnoB68t9bHM7otbnQ6xkWVGbRU4L2Jzj2LopjmrNPYZ1gAK6Fyxmr5
WuI0t7etGS+12cVOj55jtzl4HtLX/JuLXOdsDEyWyhNIPVmW/vChpbRNBhaTZJQ2
8kBsBKBck0nlAF0sWw95NTnEKU3X15lpF3xRBX5kM2vMNQIRlddJSAqjQusdJC8X
v9Ymw7l6xNQ73IOTLaCOh/BffsYQNEmZdGEBwzUV82HciEhjoicYfqHNHW+74alf
oytgNVNPxTv8RJGKondLp6x8ZilRe3fvL+AvywHanmn54vxoDY0je2bYxaIgVV1S
vjmxkKVE84YgjLMdZUTflMc5ezXMxGnGCQEYw8RKOmQ32ysgv7EU5iLiv737cAp3
jXnmX5Wuc3508dGKtVYKLHyN0tBhW3U+i/TUTnIMhNZOdCpoho2Vy2ODJtfDp4wy
wBIeU1RtW11ABNHBoqFvfsUqbJGkXTjTylYc5P2KXpYcL8447JOcFPt9FffXYSTg
GxJvOjMHRAbGWroFYqrLZlSKr8YpPf0liUU1FabNfZDVq3t2l7U2VFkZtGkViVRR
OZvVg995dhZjslnJ8Itiab/lPhaIuBhmMVViXcV2SgjnjoD8FD323bZFrtb3HIAi
K9L/A/W2Vjpx3GEptAlM+6aq87NDWhcV7qVC3uYG/N2lUKqV6P3UAWAJ4qvmqDtI
PJgfGh4GxoX6Ce/FKC8myr6eHsLq0Nv47N+lKcm0DiYZNNkkV0EPBd5J3Tp+evXz
hwnwTf72b9yr9NF5dbORZsJi6IunBwg6O2dPvqTAIusZ+5hdPQHhD0VKdM9kcBfk
tsTq6AgAwljltRZdnhDUJOCAeKcWppwSjZOg+36xyk2T1c+QsV3eXrFVP2oz+op5
v2ZP7VPSPjhWsH34z+J7oY8aoKumwRGLVLk9A5LJkVf2askvyu2bdS7sZwb//kMD
sQuNLCBc6332mRftFu/FdCp7b2lYzxUApvBF4xvgPrqjddOg2P4JDgKQbWjcN0Hi
LjyVqnZ2FuCGtRI3SPS18kTSsob2ALwHNgEIhdyZU8bMb6ZybT/FzR9D2r86SWRW
TpVMWE/9DUC/maIdpxsHfkZ0lumixXOXzmkij/g4i8cAKcdbKo32KwaG8UxYTBk+
ucS5azTntaDpvhEomSTmFRavFnjpk9NP7XzlkY6vtzOL/dOSFsfFLlPNnHakpS4r
24bLrNzw3oCw5WU7d548zfoeEhuR9vLmlbsGkqB/HRZ62cuVSSpUzNPHSICSBcPx
1sbsxoeKF8FOVOfwj6+ar0jFFTTJy8ZZroMm7L/zNiT6xxQgujGXU/M2gjQ8EIyX
4jN/LAVC63/z+ii1lhIkPm+yi7PA1z60RZy7+gujYz5s/259eKD1TxriyzJxVG4I
lhMncjpijxmZIJZmXzMSFHdk731PKlehWQd7UhcHrE2rKzWqVAboEcOpNlfpCDKj
8OpJDFsa5JvtFbX2VQ24Kp6OzQw1U76d92hEpNyuR37YuKyMf4QOKEnsKC8zDoYJ
jTwGhmt2BKwlinSBfAwEsr4TMqbg2yMGfS67QsKc/imz2u001m2F6sqHkDLNRgzB
YeQuyXQ52vkR/Dc9tUAnuRTSeiSsgVmObgE1XuHofBHK1pdW3B07AKEPUL4uR3wF
pr2L/UZ1d8Aj3m5na1wtK7+VQ+6SheVkp+EpNEhLc6c2uSdfDK5It+iiDFe948Jy
h4w13vaUQgZVBK4VQFFFg6BSTFiR2e4VbqXeYtvbn6GIWWgR2809SJCjTj1silbM
jDO9ZGfuEsOEs93PU1OTlkhVZnD2h9kAaGz2GaMWUlK83+pJn3gzjUK0x8grGYBv
TYxvS6n1mlFmX+CdB/JgsgAdv2pPGxL2p5u6v9yBgCmNj30S8H6OQcn4cBn7z2Xq
7u71eLsf2yp1MXJ7KTtI1XSrFiRgalfWPWsPpis9SWp/5umv1x/eJG13lP0pJxIn
TYeZpJozNDqbj7pk86V/lI2LMzamKv3X0gMqd3UoahLcJFMYLkAt/0uJ3pvSbOOe
2OrR9oyXVpU/xBdz1wCE9F9X3835q9d2k+KCVcIu4fqi9POEM4uh436HPUR4uyyF
mAA+sXaXzv9IuflHALfth7Mi1OsslXjUOO+3WZvaaYTe+5JwmMQSawcy42fsHARJ
S4hF1SZuHIGIgKbDNaShuPZj6euCUBUFtF+i80tT3s926mffatgl4FLHpuXVuzpJ
2FMgJTW4l+nZiAJPQR2DMJIlxm4oAdd0xzOPOywCpjbG1F85QN116Ibpl53I1rjl
Ivk/jfJdq8NLxjaOQO7RSSP8T+wrbhsclN2pQm2/xlNJEmogtoD3oiZ/7FAkMzw+
eDHnxO40v0cyebzIkx+BFGuncBjS93tL4S8MRCt29JKXR5+ymVVj0EhuLlDpjb/e
zAJDMg9EVUrrARJgQJGv/uPN1P4dvoN7ubWXSoHq57FZ3xCbL9HkkCfZQMJ4mxms
8UACs9KbuB+UQNl3OwoxG0V28OLy2ClO9iWn3/pmpiWP3JPiwvn9Q/8TMnfNQvOS
F+3cwfTAX3BhHSfXL+lt3OXAQKmdywRYf8l0SLiDDeb9NybXEDOKXV2YXfBFa06X
yA6MqwmYjlJiBEJ2uKZdwvu+OGVE+0lBXDZvpLox3VpOXlI59DGThcrF/smx0Wya
vWccjW/oZOtggu8kHorOxTwMAOkpg3vgbSROkOJyc2qsZmnLwktq/YTpJMQd3zRS
kE+9/Dv/zFXEBiyP4WLBWbrkcj7ifsApUZWpEkUFwuMLaxqVhKFC13sV/jelft2M
k3+uVNswlq3tjf8dvq1a90KUOaJksZnvUGkSr5cQNTD53pm/dNsc0Omk1rG7Lkoq
EG3VqkB1qSKbMlL8P0CAfwC2g8+2Fz2BidUl0GoqFm0u8PJskbyh004ej5d4VlVB
EoCfYYqYdoeVMPXJPtX2UgBAZ6ZSzLEmqm9ypq7KAfFEWSctnmpDRWNPcykYdFlY
MSSlQnIRBzcZQ9vx5RT0FivTitYKQXpeRroRBCyzo20sDnOUBFiu3wHUmfj5CP+z
BnN+tb/+e0rncHDgBaCfNyjh5YW+hFI7gQDGJMszem8ss4ZQCVGjQRVY1+5yHWOT
6oV2pukjL0IjYnmm2+b+JlyWbw+8F69ci/ZrD455MEPs8CNvoo/tYGYCWohYEFpL
X+PXUwRuUSaRJEHKHCc4L33l0qBpr7SopgJO8MjH1JvLQ4ncBcoL1wrfc+PlD12r
PLC0xcz4JNRXnX5k4C4qbcWj05oqfvXMOZuC7d0N6sMx3k5AWKfuGg/onUvOskUo
WOvzEDP8pJt9I7GD53Q5BrfQuzdHZNPLvMhThI1MR/6hD3pN0Kh4eO6sfQMR1biv
er73Ezab0uEYw5cSnijsPiZ8GgQjSTgZcKcI7nLsHVuvXaZseisHZnca378SPZvO
77VYNuRdl+Kfg+srb2U+S7er9BHCNcuXOSfSDGbhS9BMo2ZHnx9VFp91bnpq2l4q
U2savH2EESwXNDBKY+QVi7dQ2eSuj8cqAlsweQhby8mwST3K1nrnqmP7CtjzHVMg
KnYHu73Xk+ap5UKpoTWXoUKt5jUGqfQr706d5ZOd5iArhHdDibTBzGuXIlVJUg8X
D2pOnYF+CnbTH1qxYOYPdwKnqo2/LcCxXS8flMyDMe43M3PkZgbuOUArqeWaEw8X
XAZLcfMlORRz6rYLBGxq1al1nKM9Kz4fYkfmkf11k8q0+JGPwFnIUIcrs5dul+QC
+HBCj6zsIAUFfDIaRdwe5MA7MIdkBkznrFlLab011fJGnTJqUQqPh8csYsFL+XA7
cJ3Hblj1YjqpWWSWKDdtPh0zalBPC5tBjZaDq7HMrfQFPB9hV1S1IxelT/O/tZG3
CQeHQ+cyh/qJdS80XWJieDsMP3xgnxqW5ePp9rxhKqb+aRpbdBYm7mDACYbINM8u
cHkQ/J3NbrAoX0FxT4I3oYsNnFRHkWKlWH7WG2doG5VaH+rBsJ+mv4IQc277/8xX
SqA9FlbXCu3PijCvaXGDcG+vBnLUEA8PRIvVAWOgorg7ZmU25JYQ30JucuXP8AHA
y8pLavbDHoxznxqh9ErpwhufyLJ8pGBUt+yXg0Ygygm48/3r4H9ZjKAzd0hnqMQ9
9tgfvN6ekAXdE6fDS4TWoiqjnRjgqmkV4zizAw9svvSCTpL1tI3Fy/Ku/TGa6gM/
mnhDyzmjA0ETG65tC5CfdvZDUUogbICiEeg5x4tgfhTHmHcEfj4lYdl43AigL6N/
YQjIz/29ZnpIyAM/zxqUSp4s6zyRMSCEmQPVxMrB11ZYixaC7IIVu9VGjfdmPtpC
A0Dtt+eMGBX6CVKM2w9HXncuFVGEGabSOECX96oK9MoS4BtnuLBhpPa9/GYb0T6k
N4MsodlubhkMVxROZRIPz3aSCnpAwgnlQucivoBQ/l0I5QLP9r7Xx+S93N6I5Iyr
6UgYlVv+caH59kuX4DaKuH16oAHHyGjL5DsII38424mIcIWWwbl5MNWG4/lRUmdT
uiS+M3KAYSzSw7jXwO49xHZMKsIafgZQxNNVjQi0WiVPQL72k130LKbdCGJkgqjq
fHhYMSOXeCayJDl2BPpxgyy2UKAAl860gp7D6NcaqMxxo6eKRlTtoPSzCq+DMVZr
7lFo5jqAvcHRB+dqDuY+YJtAW1+R1/5zkzeO1gLn+B2QU7bgWNPMlSjh0S0Jr3lv
/UEullBS0BetQ7G3iOkVFgQfeUiIzAiri9HfnrFcaKfWs5VRApGDFUVI5J7omg4d
PEB9QWw441G46DkYRVZT0hn8sfR9GdynH3CFXbJMBKECSexI9AkP9dQXevaKBZl/
M2tyKCdf8xkjD4phXpjT5FFeT57/40XWkJJVWipjQ4kumJRPxak2uxpJp0fsRQNG
D4sguaKkNr2ZPKYV2tdHwsKyk8w1Hj3jWzHx0qWyPCJpH8RbQsbma1Qbm8ExFKc5
4vnf2WcKA7RbIPk7X8n9LYO42rU9VRMTZPSqVXuSIhUFZ2co593TiCMu7NuXWUYr
yEk59nOgIeNR4n0FaYvXjr5tqXssm9CFYagw2pAecSosfezuEzTvePl/ffZlSHFV
qDIxyh5n2094wNtbFFS+Q3lGODDqno/2FYcZ2LX4GKTGXVxdSJw0oXhL9uRCzI28
0/4oqIPPpen+AFAYKmF1NTW2OCfavAQTg+5mOx3Mj/qPwWfbI5OMZgwOirRqiath
xwuC048ZRIfTN1yyQnOD6RCtmynlFFhioxuUfxya/+OLMEaQyrKilBCV7LX57na5
pxc2nGYkg+o3b0idPHsiXYWrgbx5tXQInp2RaFU8maFyO7N0crmhVulxC9yHOBFl
mSBUw+kev2LHeRscPyQYAuLRYC0ykvECUVUWfuWY8hdPgy6eQ42zocdSKVtECtFG
Wc/b8XnU2zmqq1hFaEzj/X/k4uTC9hEOsDOYUqCadScXx9+2Eo2BYVlxOuHiG1zP
NzJeLiLfv7tPmqS95fBv8NmgWX1sgpetiea7+eKpEivvF1wPx2Fb9ygk/9uWVxpc
pU0xSq2D742dJ4zDIalqDbj2PZgPnPuYoQGoU34As0avABezpaGHb7ddvTgBxlNN
z2MzJlELeZ3gAnLdeY4zfUYkp5VeieiKM5dNbdH5TK+IvlfBNWqwP98XJhpIGE4U
KZ4KFfALwZwN9iC61wH/mQFfholT22T4D3xWcudHdWSqA6Sn8fjJS+MXjv6ckugm
k7lFB1sCr4aD7/1CcenykA8YZbsk/iwo72gOolw/v4bI7nFR3gh6Rpm6721uAp7L
1k17ZUP2TgETPEJUdTEJm7AgJGs5CpokrAj1PHgEX6Y6dQfzSXN5KvjoYEWnK2OV
Dh3YtUrpiLo6QXa/sIa4EcC5RByJB3jx2RD1JR+o+57gqWvCJWZCdqREJDLRABd/
votLO5vj2iwVKIPKAZ5IQDv6BfC254jjLTOgS6ryVZgIyiKtAE5r0Kz5XOqRHMM1
UTFR+p8xWnn4jMSAYnVWG9LHzC5xeOPn7wGBg8krV4UgsPkRNsrBAWETaNwymri7
ZTVOjXfrugJpxDu69ZiLFqjXYJFOHmpvJQrUAHWqBhtQb9eKDJZYPwaTFp7dsppE
7duoJ62PlvD63Be7Pa1tp4U6mM4H11xrNlRqsMagjLq0TTr5u6obgNPhaG0fmTpo
O8PLQ+QqONkoXE1/Mi7YiCOQHGZ8kwDikt3iqpgeOIbG+GMbQzmZDEqTXqukhLjL
6bRKeQr6oPRoRj2oiKE8PlVx2JolMSCjmuIsm51rc/iHPtejFRza4UQvNelIMZ9V
DYbNku9r3KugJky1w2IrgJFgww1ZV+i99VVJ7BJ6P3ncyAQ30x6tGV4HlPN4yUHB
cNhoir6JDYcNdrWY9QadCa1mu6y71A6a2DvJNH/YGxHHVQGnGTSoaHcsfHs7vNpU
8ZC6J10vpMeuPf1mmiGSV7Tv9DfBRS+QIEAtcRIH9SZTLSN06Ba77EVycjQSYzC0
huAb/EUVqRFcwDSUQpU4Ds/NTw0YcYQdymM1NulxRMuYSmmUG1u+/AOL6LDLWiBB
PWoBCKHYZa1U5spF5CKLzEVVmJtZyka2gPLNJmahffY3KCW9ZDmm+p727AaNTgAm
ovMDlAEKtojbot5J9RwBXor7DoXF7aB4Fa10L13tzO/hdVNIZzlWIg7Vj80hyJpt
9Pi7i6xQxESOKbWQBSuBETXrDi5tDkGQ5BVW5ZWJhWY7yISiwXVsnHeUWfDgKnW4
C9QJNdS8EI1H5psLgSyMHcjEIQ0WsaGgeJUN+OuonSk7jY55xsBqvCbNZDaqJz2C
55fdcSncSkDsGYdITaFMYsINJqbqqrK5K55c7gNhY4hCTtaIIRIQ7pmyt/00Ekj+
F8ZLCRQAxhHQn2mkr2cnGGUhQhia+tvTXAGHVndJeFWT+pUfXd//hRviuI2UZ7x3
4NIwGTk3+z5wwA8AjLrJ2LYdrLu4GdQOcivCT9xo2D8/3UiL0R+rnEzaaXKE3zTD
3KA2fuUOlB9HXsrvRgaoHTOP+g97oaPlh7b3H/XWSLPKck2M/1heOsHXZ7wH16uB
UdFhx8FxDXCdRC/4QkKRDXDTgCmpv+trkSHOF4STL8TW3NvsFxpN+LTHG0TGD674
ZPZjvO1wOerXvHb3tztI6iai2c/VK96eWBE75mBDl9/+7GWqYCWlZXsR7c/5V0Tv
4rFe9mKvtQ5dz4HsZJUg5fyDpSNrq2gTZ39B2caWEvXgMFkVL1hPmzgmfjuIiSOU
55dERVjq77z/khPUN8anDlbRa3jc34zpKRDMzoQTLdTcUGcqK9bQC2UbRM4sYY/0
bD0MVdg8h9x79DfwcXgd+54NuGzKwiarvIlk+AO4n6HDW3VdLaAdloGKOcT96HGh
XJxeoeU+4nHhQFtDZC4RDnYXylkYs31VUkPC8aiIQXhop+TLPwOeIqDkJrTQxapR
s8Z5ypgLlg8JJqnm5NgqAWZkW18UZVE5bDS8vDpeRc2DrgowXgksqTmhVfjR9o8L
0KQIibANgHzTRxR75g5zL735T+lxrvytAmpo8dLQq7Ia6UEvVoXlHgZ8yMCS5jdx
znMRoe7lQyFSciLXeToIRBKeyseYE5rMiBBvdwjxpWj5rSteBdA+j5JcohfV+M1o
zVhJaQKflgfUGJT8wcD/2JlrVCE00GLuT4Pl79DkhUTSgk/WWC32WFzxz7rbF/jr
LmOoJDq+SaGKvy3EaqGTb4epyJ5SXBq+P1sAe9Thf63wI3Rw6R22jxUEWbCdz4du
EZBO8BPl6cqr3Ll4G6h10uIH/xd3jSU6vK1gwgIs8rTgPemUIPL+VSfvpzEcCt8t
YzTePf3U91JyyP7udFKz2o1oFBVSB1Wdexlplg/sWL5YGalSCr2qhpRJibjbCwLb
zN8x24THKSrCALKrsPWQDfr6+sz/wwwGhomFWA+x+hUhEuHqHeXghfLedSCsGSOF
ypyRB2Wn1bD+3bn+dgtegmjeM+PFqAnJGTfj3lX89S/AZ7VfKL5cqtrcLptetdSm
ad2neeQRG3OtkzAapf1D7um9ZkAZGVAQQ1CIUV9jnxsmWyppHHJVqceMm7VNo6Cl
q4a2CumUJc+aNX01ASzQ5KOoDPVX8lQlAPDz0jalxvfSK6cuDBkQqpa+ZU3Kj0SF
mivdQqYgYX0D5+0i254tms9jKEk9p7Pw03e1QvDhImxzpTVb3/sGTySii2GOSlWz
fqQ+4BaDplrIjpaGniAB8o/UbAk993zLHogdu+dt0s2ld7nWAwPXFQSjS0aOmBv+
QfxpH3mTI9WLuqLJ0BliokOGxq0CIPFUP159KZPvFwhUTcZXniE5ib0ReoruC8Om
H5hSQt3jymhU6X/BPZ3geMuxPZttWq87kT/auVf/TMMMxuENCNII4gkWVrIolC94
pNHTvVDQl7jitCTBzP682hkgtUqxd8JW30Fdh3Otomp8AfJ7ICe3Lv7Ww3wSARJz
9lqRATITYSVQVaYF+wNxgoE9G2v/DUv+LSqIGqy/I3qK/3GfJm+wy9LEf11fQ2My
9gb8YYlT4fyv+Wt4JGEWmt0wV2x65QZAlrT92uV4v1/eX6krvuJzvgGQIOtNt7UF
nx391gFSZcmLDWQvSUhIflbqjWt4KjfI3TxSRwTx0uhUy8ZVVClCOVuGfKa9pVll
Rqaxi1rSJ8pozTRxQPgQ7tm3phfaYrTvGAPmGPpEtnZPKyMQctavU3pZ1xft0NTI
42Ajsr2FLPNqqr6/ljRPZQ46poVYaqkW8FzsBJ+MSPabtvzlZEw9tYzyQY1A8QKR
2xokSAncZVDTwrdwMOOBwAbJdS19cAKmpiRVkovRqE+3mLdI7WCvBWhWxzuMvM6J
aKDNpsbxkI//C4EZF0d3u8oyF2P3lRGbO0QxoEevSGJrLq2qkFOhTfmKYyFXupe5
xLFCd9j2JDgqWJmjswM1hqkhjjkpKHBZQ0XxkF5tfPtMOfTKliFUnhRtRIVGfnQ9
cSztz8IFeohOXNwr2/aoM7L3gEKC3qlX/V76q1SqZn/FFvQV9qkdzbn79y07jSzB
zQb3VwsDlhG57naAAo4IB3+Oo8oPudPV9EZlaeguY5w++eWv2zhC/CVL1qAVw9Sn
DHzwtN1j6fmKn8iYC1/+LGFT0eINtUKtM0IbfU9OPhjq4WMrs507vYlmTwj52/53
fuV1jlhq81RPHHyQDXdVbtuVtSR2Pfhid7rBTSJQygsd1+getJF29fUKZmuzLGug
lmjz6kjgi/2h1qYiJrB94H6vB7Bc6H9eUIGpNcty7aitABw6vn52DrLqXaBZfE7q
ZaGWmTAgyXV+NIREg2yM9O/mp4Vs6T+3v+58QsuSyTdk/PkGVGu+V2AgRkgMw5Qq
rFSuW7ie0C/PqAo2JIwaBFc2wGgxCdiA9E6jKYsNh1inWMlg7Ohrro+Q/1hP+uxx
E3MLHyxf9S+0/eUkdvNpLMnd2wi34k4+mKUhgf+fkBW+A65bDqjxYzYVAdPiVbZZ
TaVMtuv+bWbT/0HiZT3OlAl/Hk2MKyItC1WXvGlAQac8fTYOrWrBqaK40CMWdj7R
f8zXallppfbtL3wKSjy1/ZJw3quwlFnN4OF17bGhWGGo8XLTwoRVIS648kowAzWX
cMzC0KK6uNglyyJdLacvWNQJJPXfgcoU4bODnXck3l4fsDZnM/G75dMsG8rZIE1g
2ZJoqHChPL9DrTN4D9HgM048a0z/F07yeE6UbqTxHBhOElJZ6J9ZN+nvr1UWT9BI
uRILlfqYtvYud6QYUk1G1llY3qZyxr/d3NoLarBSzEIZzqQ07a9xEEdUvz46L3xG
ATMvSaYCcuV+UQgImsTAu3MgQlN1dG++8LyRbKs4AkJ+gLoeInlDYYes4kooz3Yx
wYsHkZ+Pva8DT6kWYbJpMNfmkhlkToYd6ZeQlECk19LNpxXdjUsJ2x6C26wBjnlM
P/Bbx9P1GHADgIjtN2NyYwsmWxzkCrN/rqF0ROPSt6xtduYOXTyN2ty+3tplB+HD
Cd69JAIe0yaWm0PgOwhL0ljrLZI2UWqC2Lj6wyzGxhEoX6YwYP7jnsYk2zKxQlJW
NQ1G69nR9dlMOjy3JvDM/TZHLCINzYk2SxA5xZ1EY6oYbAMjhUt4CeRMvGjioPja
ugUZi0OThThhmsGe8bb5WNYFVrqDL2booa2NDcHhkNYaHkgZ953y+tL1AvFAzY/Y
Ub8dA72V0I/4rlYz8fbz/So2IXztHffzN61Rap9mYM+a6NVpTysPRiXG6LWH4Y6s
k4MpO7D6UguHPw/8ouPwJzfFjXqZ26YJBmYcsm17etV/8GA2r3OLFpEanb+01keo
Q1oajIEY3r8ZOWn0H37xrMFDrx3X1cl3yMLp/xJBddbEffneEjStoVbc6shha8is
IC5PxuAJKRXjQJrBRn8FPmTTLRpgJy8L9TFG6zZeZaXRsuMPU5X5yDZ3tAHNZJA3
VwIchVohWCJQQjyXAIrJy0unFPZM+5G9Y2ZK4FVY9PI+pJ3p0tEw/o8arLyODEJG
xysvrlBpi8ii6zJlDyDdzi2B9rKXrS/Lu5zekzg/3OS1dzmYJuYcEjLCYlfH9UXW
kO5oGV1ErjW5bVhg70YKITwLXMJWEdtErg+6DI6TCBH1BH8rSNZ+3Uu4bz+jaj+r
ITo4+IPsvWYtI7alVq6BCciy4KiFVCQXDzR6pFLxab7o0tthxt+uoUetSeCPUTq8
/nd4pWuZxhT2v76cGpkpaAllfbagTNIRhJFXakp8slKNiZfLm8nj24r5ryTrf9x3
yt5iDjBshVOxavjheAQRZi+V/psazgXr1G8iYpFcRZAZDvqa6GC+RzlwOxx3Ssnk
2K6nD6jq1ijzczzeJrtsLwVA/GTryfa0Is8keOkkJQPUQzzVviBknsTezRel3uSX
QvK7KITC+B7M7VUdM6KaJqECV8eyFGG72ai09vLFTDsVtr6Co7BcMwwfxsa5QXPX
z1PRc+Jqalk9lvMrnyOv3k99+ZqzXRYVA11Z5tUK9UTS/skNU9R4wpEfKPDf2rXU
/xVcmKiSaPxyQ2QEwk8cIbIgVl/WJlJoZ/caLFaigrC3Ahy2HyUjiZqXRJB4xif4
5XpuaqPZZsaHxTBdSes/d34+TBJSalQQqXuojDX6mfoQk+mjDV1jcgQuI7OeGwGh
beF+mPLB8vcPs2r+LZtegu3criX1zK9M8gXw9Rt1+dbsZlQCu2cpCY5oooOuf4c3
S6YhsvBDo15Y3AFybVUGe8opEOucJpCb6JasfJrSC7sfNlzWtKZYAY/PNeSef1vf
NRfrp9hdw7uMGmA5o5vOE+csBC/u798+cYGkVn+A9fNb5HuSEyARVnH1nm1D7ic4
9VegdVSE03TmriY1z9vNRMoUCkwieUTvhU/yGmbZw+HwBhMBSj+iEVnRDlS/1YyG
MdeW+prsR+VNepX+lwL2Kt8WLJjwKeEetv8d+4BAI+gp2boU70IBw4PVZsFrA27r
RsMKYqatxTgYOyBg7ufPBXsKTLjfKxQ/G8jWonG+pO9rT+QHfNoJVj7gfo3r1toQ
j4csuOI/GcW5veLcUBwpPa5IAKxBWV6EsCHyPxfVq1EDJAolqzxLeHv3VjGpJFLg
ox4ubs/HjVZCFI57pwhPrDTJsO6ZPNUm7uQ/j0/kWl2ExHFggjEzqqAM6rs8oYGp
xJDfJQ8+2DbKdDspXJhajXV/iNc2vhnyvcU7+ChPrC1y6Bb8LCVdDbrHWuL9ULzA
rgksU2n3dsoDZ0OlDSBOWdLnGAhKWNYnYNC/4g5Msstu58MHv1mQHVe2G6TL7nE1
j7oD/Lknc6aMfv03PQDoRLgyz6R12OlrbmXhk5nfxrHXz1/Z/WUK+u0dGyjH5nLc
VvKcVyTcSdATWwOQxh3LJ+5baMjd/Pu4Li+ZggaIc13XF9vGeZ/KoDtBz39Ik7i2
fkVRaViTQOKdUedRKHXAQlHSL61wOTKPuUtAjgWx0FlRqzKTyvcPfhFw+xMt/s5o
6xEjl7vyq5R1BCk4ZDiYDLOOafJwxU54ZBzPl6/2nc6HIROZU3t8FMhFYw8mVyKi
pDkv+1TOF8Yg10eCGPM4JLiTLFq4FCf0rzWNPat3sQTOgQagDCLjzOnjbU+B4ugm
ia+Hla1zr7zEJJPDefkfBIsKNwKKZWZunKqkXfHDP5+GPCd4Pn7KmcMo5R5o6ptH
th6V50WcDuUg3NmydKpQL4R+bjvqV7Qj7PzGigpEAH4JN7bIy7LtDKssWrnCBP5V
padqVIViTh6YuDSsYNNJBZtQdFgHJX/EG2IBPK27JwTHB2p4gVrT9PW+yXbGkjJT
+o1piLUSqxA3z3S+G0oxGydJkcadF6PDVkn8ABJOxuvMzOyAwXosRxp3nOKkIN4D
6McfgqbzpGbi036lqJ08s0hbid1AToBOXb2UtTCdVLPR4+FQ1I3b/0hly5oK7wxM
le7m9+yJFC+jfV1lmuVNSklvUklina/1LX9InFviI57+3e6XFDeEg0IZ+ZxU4Ihm
JkTrvuzyVPZ00+DeGrRvz5prFXLk+TufHYJ1+iOjIMqVf2hNQ9Okzi0+7mvNPcLE
BZgIi6psqfEh8kLmky0KWI2uqcMWmFJKC4S8Fx497r7JJmxEBcGmvtZ+1a4t89fS
KvjIoNJk997Br63BhHd6JUIcVDNvK+g9+sBTMNB7dsNFl2i0fJ3ZSLNF6MmDcZSO
ApsByrv9oGSl972N7AXyIDoDSenOiw8vPsgEA9mBBDEpVeJQ3VRgTI9ghvezQotz
xVj43cOm7VZXgdaC3VdlQJWX/pzRdmiES8Masv3CgOO/kZ/1YwXP9Y0dvdjvGCPQ
4wEXTJqV3zmNwJa250qfRAoFClyAdJP+qh9yIAt3sVDLCMHB1QC/s4GSEjVPxaJT
DzYfFxE8qbQFhhF7Drj8HOsFpu0zaW09G47ouLXWhDaKgiJXlLpDTqMl8trJTxdx
Z9/0w+6du5MS9HK5qyOuMVQB4KMsV7JkxSLnI8O7Qo+BDbYzxlDNT47mwgp/3CJh
t3MzKaHe3RDj3Alv7kumSzsqBK/RL2YjzwWNKkVa0NV0cMfv4OW8ULlnh6Sxa9KN
0h15pvqhDY94w7lR4jJ59Vms8LysbfjTR/nwaeXoiB7njLNbTP4iUBBvXtVZUl+T
ydi/QY/lyBwNNqwv+TdpVtzzmVt5YDeu9PepEcRsRqXkj45Yy7z+AZbXi/Mrw0tZ
nAr6p+xLeBfgOBmNq0ptce4XpGyUYmD2RTY07FmiaX6AsqgEf2HDabdIoEuV06OH
8eMfYAQs0e2RorYJXdbAJ0pzaZAqsrVYQf7RoQ3WKAnoi/IKtYTANMzN6ChCIZ+f
gB2kV0DlrRHz0xuRlFiop5bJoc3S2dj4Z+IR1Hh6y5KvMA/dmlJpGBWf8csXu+of
m9AJxvjNWSbebXe+j28F94RQNc/0XnPl9PJz3BmdV2tolJPSEfLt3TdqEW0ByiIx
6GPSFTtu2qShJPRShiDOpNc4oJ5Oxv7cBcgn8UhsGTPt9LxjJIhv1ZizoL5yn9G+
bsImz3X3gNwoB6++ez7PpDphKr301g8iqB91R7EbwYsuVgI9oAPenIy+wTWpd6+P
94cmIorEzT2im/35fmnDnLgZLXZXSp0WQAsHq8v3LkxO/ZyQ/deC64dCntfJps74
pc/TBqqK9zHwLwhcw2YUWASDzvQRZLkvo9gcZk9lc/gpVkCbYTKmaEfpV1S7pf1T
iZ4AY7J2XisMtln7LZwgHR0WnUnFN/Z3jBLBVKzmeLKY3LikuETy5mItnmUv1dw3
fLMgJIDjvygGDP1SXCil8QiO53xvnv+SAJLFvJ91/yx4iGt6E0nDFYGxZFHS71B1
RAz1cn36QB1yNrSPiDOycbiSz1PUEAimMe8iFr55H1d3vp31wwql/mEHKqz8ll3s
ku5LjGlhlf75et1dl4b3Oz5762R4AkdEOu5cSk6NJgz4/gxCGAeqgc99PsozVcsJ
0IcrxtRpy+1/+DeOfNA07Y9JZ8E9vuDpBuZrzRdyXAnsNU5ZhYuowzG2Id5xNJjo
hHazwiW7/zcqHVikEr1JuJqwXOhPgjqucBtbC4fuvkyGW872aAs4nx232DHS+tdS
lfL8A3WxzXFuzi2WxUAlrtVBa/UUCLEFTCo81MChxtmZptz2NzTVlvSOJGKZqazI
mIhTfajM1BwNWuZZ9VMT2gyR+sW7P8WMbWy6JmticiufiPeDrvDcfrJcx170z87l
BfGkFqzOlE6VzQ8sO+F2pvtDjIebLl4DjN3fZYR6rr7Mm1pFqUlnmpl4U7EViaDw
O5MctqBpm4tjm3gcpn2yINwdXcQZKjPIiVnHRE0jHkGZTy/YMFR176oBwPldEbZj
u+Wh0TM4LMLPuOAG1XCjz3CCUtxNJ9JP+yEkkDRIXe6f3kkf/fQV4uvu+tUjz0Eb
KWT6IF3KcqeUpFLuVmYIlf5N6ykYdxnvK3uwYpqxGYX5mv5//R7mQoPktCKw7n6r
nBWBW0QDtm0iXW6LDsE9t3SPvzl2yJvFmDRFCQO8Wlbp+yX8y+E8beoPARSXbxoe
+JvScbvZ1yPSbiF/vF4wXNLEJpLIV3Cnvw69aWj4nVAU8xHHSZurygs2UPLhItnV
3YHG2mfHS4u8ur53h0XGIOSC+dMd3ReueGNy8QWb1FpmzTpEkY5biOV8/GI3jJB3
s67VvgLT0Jz2BzRd54nl9MdrJJOwcSJau6s6xqOd8OEfVxpSXw7f5xk9HpAasQ2G
hbPe4PnyhfVsRxTqRwFMRdu8qS8L9GjzBzDLE/+jNg8yNcEo7KKrsBsJI7wWU/gn
hERNQn7cNVUU+k5qpUaB82eYl5SYF29tqaCddNxRGCB7W4JsXDCQ+GItA/lvJgIt
kvmeHUivdzd2G6HQvb9dj4UEmZvCGEag7h0OrvPwHwfbYrqaX62x9yW5jNjDGq/2
dZw4oUH1SREo8u0R6ywL5Bh2d0yCvqLP7hA1m9hcohLhGHfZSGOI/ZDogOLC9h+p
MUp8Qg70dXMbmYV1fGglsTmotT3vVv/V8cK5EmdoZBMfjj5Ogza4viAzHDOHZGB1
3W+slq5q/bzGkzKzv53Di8x5IFlQ6z/TU74KBdLVQDvLka6eRqPxWhDfK0e7KAca
KBMaTXn5Vi9IxYyrbvXATSruR/n5WLojST0ZtOXgYK8yNh8hmlVBVSOGf1f8Rx2G
lwmMa3gzZKI847P1eSC0ORAmXm+neKdt17nG3AglS2z4AmHaHRB8dOLxywp3GJLr
s59e/NbdM4GGcBUKgr4PVXc0r3AuIdEfeBfgY8jnG4mMnFJW3yuEq+SuDkLGO4NO
f/+ge/Mirfun7mhmFlJwgR77+uGNSiIJ/yY6iPICcRuqGYvi4/KxHvQV/UfLATsT
VCRO5JUtkLOOc5+hjxUSQBqHeZwqAEw13hHgN3OFZnGol3vtWMODeD3K4jtPwDLy
AdmoU7HCcgKZ5mnUBHK4eYRxCLwysg3cFUv1KyE4qXYghZDjPyUb2bYFGuxUi/fs
K/GBdjmv+l6EQGXnZvCGYV9k0av52FVYC4KIwcCujV+W34sqIXBArJBTiPsp8d2j
+WV/cRRSWOdekiBiMBMQuq3G04cWop9efqDcJKy1tmneV7LjjpBWcHQ4H3cPt+kq
U9ZT12GCHIrTkgeX/GXPS1JKpEANkKdqOT7RZ38IbySF4jwZLZ6NoMhuLnZzbAT2
biRnhVIizjYOFXMHU0s7kSddPzpd5jwqPHZ+EPXU1Nv/LAAQC1RHePh8bH32nIe/
i5CPw0L1EeUyk5zCzVu9n0xTaFWazldV/9mz9Gzkag6zPFjCzPYBDHjbkkP8jCFW
DzvtwisNa03R3ko1en3N67elGnTdizaEDb0hLttLE0tCyQqKrz4bD9R/4a64n3oC
fqHsJZWFOGsDnhyC1/AKEMY8esnN/QZSWpButqGJ3fPc0axb2RTaNbhsYExddTSh
wDdGJF4Vo5LW6W9UG/pidEeTDGNKTlIW0FxGo0iQStfWElo8srt/VbwdxdRZTV3i
yhfBO1RMD1pYmlWkAD0fJ2ecea/O1bqlxJMwVxlpHeUYI1SxsbnAvif+U2QgncVy
Ey1JcLHD+i57DJfbkW4WXQ0ZmX28FUn8HPcXZiHewZpDoRC2kIeOA0xbE30X2uAD
kK1Cfgme8mFG+DfFAo1fxhZw0D9EzT5oUCJVOletNbpHwwBRF9gHxylPj2hEt4Y6
QENkYV+Kx24DgflYy/ouCi/LzaP4gtFko5EDLzP3k10mi+FgeflhixPMERENwqzD
60VjaOkBjQBVNHD7SKybO4cL4z9qzrfRYvugrNlPS9hWhG4ghJuux2G9vUTu6Anr
qAmhD1njm2go9TiwPhRQ3udU3UyNH08y1nDGqFiUf4c6//93zh4UkZZgWiZosq/m
JHgjsaLrKkCU20lqiQekpxKzGl7aFzcuPbCgOdjn/vZFof/TMAHE9srtq16cHp1v
AyIfhwcZmYDogPNimi7TlEMBKXTo5f8wRoIkKyCDGYOwYTJ+3QxXSnV2tg7fwnQo
QL1DkT7Hxqe598EF3k3WYcg0Acj5ZLbApYACtEt9CShEz75GP7BsK8/R71KXBzhI
aw8jFRKhhDH5YIo+LUKzCLvmgxANYIEIyq3kIkWFp/M/008hG2V5HoWh6pVwrZMC
zlafsWRmi6y1DxaYXP+rKVOcG3TpqNqWhx2NiItUAXkKqPMCt22QWd7AB72j7dYi
Cfo1BrLTNHewCM6XkeqVBMjwREs3FlYdkkRlQ0tDZVNN7gKlyHR4lMqxHYbvy/Ar
vfVdSGY43GMxGbJjenEtxXvUpF/hXuxLebehk6R1/eidiNkGfllEAztUsZsy0fRz
qtCalro7Jc37wbBZ0bPw/47y7LVsJ2sQw1hcTSZl5n02jn4YkgIWsXZ6mOz6gdlp
gzH+6Gi8xWX8O53JflNV/3aTd0waSu8ExFxpTGJxkgBirAPN+ydDllLT4IvWwH3A
4ItxtNrIfIkunGZ4vy6xNny/PS/ttJknn8e99CViRDUg47LLdGEeBjAJEUUDxL9h
lN9hIbQNKv5dTDbkico2o73gOgs90YZbqDrKgi/GHPS9DhcVeDAxkv3qVGtGJDlt
6KjC5sga5LqDxs9vaPU3Rq7VUjDxmT3wO/4ogZ3b99XQhUyXYC5xI/Oxqvfbn25j
sMDACJs+aBmfaOOnSCC1Gd6zydt22KCZKQjUVrrlCLhGEUg+J2DQdlSiax7SOg6C
Zor17ky8cvVhnUv7HMtQ6r4XP7oOS4bFMQFuJN7fv5w51KqPWrXSJhOSlY1UMkHx
sKRUEAADGasEdurvMaAXfuqUTOSDOL6BlNDrMMAL/nSQHAeri5NB+LqnlH0WeQ9K
jfmFCn1JEDzT7iOl87KXT9+hbv/XJj74c01UQ44mXNEAyDQVA8JzZPkP8p9SxfCY
XfIOCyYK77BAeoLQ/47Kml4rmsn917oOXYc67DJ0f2W3P9N8vGj5xV4pAXiyLRw4
r2O4Imc1QUgOl6mp9KqLcSUkl5vYjR/EVIabEwLClhYHpsf138ch2WHGRVlYJ9Nn
ty7XBs0bUa1V4Qy1WYx05HCQDkQNlkbSXtY6LscnVQcUTMmbg9j00noLo8OPHExb
YfzI7RuhpQylVVg4/BVCKj6uPTVataD/8RCeB62pKthjQ9lRizZN7F/OpSaLxpe/
Owd9Br6tNRDBofbIdHN5GwCI+xkttswm92zBuAJGlZBVHfswhRh8H6LxGNEwaU/h
0ptqJ4n7V8weIqsLPSqcxClMWLRx9VuR68s5sdm2PXUdU9Zv1qAT72dbxuRZlBOC
XbvTy5tSqaBrAFx78EZtOfon0WYFqtMp34Wv5raKShH7CpMq9bVznETfCTNZExWd
cnmvfC76wXRb/5qFkT+WSkCxymT82e8nADkbCb21GaynM7oB8Mko/xI2yxZmu4/z
V3/8z0fZZprIK3RT8gFGKx3vP9LlvlC11KJSlLLttrhfqqLjqElwhY9EwB+ioIt2
8PUHmkgDHMeyaj03PPeqvz9WuCN73+e+DHmDGOgKuXDSTpMsaK4RfD1NoxnrYPDD
Q12G/+2XNPr0cxbHwkkafjjvcsgFJFY6BnLn9aMJCP2Nz0lKxiFMlKCpMqO0gihC
sZQysYJfpMx+RVA5HVxrNW9cuDC8zqZVwA/HgeiiY/QHQgIl9UC/w8zCypF6P65t
WVNVL7JU+vn4idLl1Aya/fJSotDg37LZgzHa4l1n6nkUIDcNXlWFj3JGAVvVi0XE
NenQqfJU099HmYTjeuhgsO/exD/spGcxJYdXWdD/R96Dg9M8F0CNMf0ddGjEgC/s
sfGzOla2m8npZS+etaAPNvVR63kIxYXMRFdjAe71Jg6HK0fYMqKIK6AwPJtKI9uv
3rmgDmtmE+fr3NiP3Ba3bCeL57yA9F3E3Q4AXxFfFGTRDp7uBhD9POQSFa9kL2nr
5pdDCLtyt8T02WoeDlbLyx1GftMhNx18u3Z9Nba+UJiThPrHYVEnP7hd36h7uaEL
cQ9vrO7R0/R+6ZDuqtnATp32/AzNA7mKp+L7tWVV5/eqCUZtH1OIEFyoO1wcstx+
VT84slsM0ae+aayQLxg3nJAS4J0ylDylEvJ4+U1vDjtFfZIiOw7OXAP/k4F29bfh
ezM2mgCI0jMynmSfF47YhURUy+7KSqJLZ6Bp7PTK9adcRWcmuwMsqO2Y7HIm/Qls
nnal+yLal4l7QpdjMPUh9Ukw+Qk3cBMx+5+aTtN0Ee3HZINEIxYpmUqPLUlxnxL8
ItUk5kUhbpBxlbtQ+VcIHotpImC1S1PyK6ksCruHRPq5Ea12Z5Y74HLiACoM/J/D
CoQJi9DHTaRW/H3OfFUgljs/S6PG5ymVfsC2+2Pd6lz7/FxqQG8TFLxMCFsfwkfA
tLyhKBsv/0bR8dYqwVDrO8PuLr6ECZuAJVlSihfVsA8Ke7/ZD1EBwj1SgozY2CV2
xaM/sKm9MK9m3NpCx9V79avVMAuHBILbQfWFsJCEW37vjY3MuqjdXDXuzlx2a82R
2Jy6lbT4A8YZ8vRp3c0aFfBIjWzRKxCfDZxb+L25+z8WesdxJjKKBDTENsPOfGrt
Zkuswcl2LiWaprv37BQ8RAHZKTXPGlyDEBVZMq/YbtA5X9OfOCOtlSbwqchf61Lb
hhTLt3/SR3I6fOLZx7Ij87RXNkPFKfQg89ISuCuOEruFPwy5QjK+g2R/rK35txQH
HS0OfLJDp2YGd5PbWCC/+tdYwwXzNqe/0nHUfPUm5Xb1qjWaK/plHHlXzO/rqPA1
z+2wDL4y8cxnqitJ90iek2SVF6mKjN/9RhdZIUSptG6yC9zFwOXreA2+lecDy3y4
KuwhJ4HCQUKCvio0T9b/bMfTHIxCGNRgM1hBSrFYJpthUNUcQr6DkoFLpzLsiZbm
3YJ7039HXaEd3ocMgkn/wnnifYUXExT6Ala+2ncU4nebKF9zU0TUDS9wgMPjsAim
rkSCdy9oqndVA6aUS8UvLsjcvq7rzQnlIvjGNmzhCM8OIM1uMHViIpP3M84tFh9y
taGFmukX7L11uMnZ3YtCASWxk1M9xxxWI0VlG8aDZTcG6QR7J5DD/xnAiFW2Evpt
V8gMS1/NS4+BIKK3mQWYuR/jVp8V3fZYIuWkaCLcfHb6XY8UdoFKMpN8YnXGz3Bt
q/OqEpOXJ6ngIPieXO9qjnsSIMr/gBT/GX36bwbbo3jW7+77I14bd9NzE1oabBOe
k2AzYS0GX+3BfhAtWQ0ggX+4jC1u5RBiUWxHqrP8Ezi8GTJPfjkhJXbAlkNm5GT5
Nsj1B7HJ6Y2p+srwOOg5T3TzKFDGf6X7DS8gVBzAHMaWxintKT8uebDC///wEfFv
MO3XPtyT/X7wcaOIBZew8Wm9bixeQQG3z0nprN8usyA+pr3Afv5iDsyfpz632a/f
FM+ZOikcYx893xZm/AhBOD4k9lnbe3BGMfbV/fOra6cwBgw/tspPfnkT+Dl5oe9B
bZCoDdj2wgtthvdsrdEvppUy71BhioTla3/gHbWJRW2a80vmDcrrbCa1w2gGxJtC
nJGlcRgxXaYK/fJyZK/wjfx+5W0fgSXEts7ftGL45MhJQWt9KAoeMJj99h0ukEYy
noi2IOPRMXIL1RQBSNti8nMHZdAJfdZCP1HdIr9/fiVrbgHHEKe8Rn5yKG9ad5iT
2mGGNCH3wfKtJx1MpvGDjpIZ6LMz4ZFeOPolXWdY5dkdjG+Ck0gg0fv6CbaieTeZ
K/bOG5GJg3OJeAG1mlWKqs8+N8lFHT8MhuiwKET9t9UEz38k0jnCnA8FEW9Qsx5G
QBGyPeq58RHddH01w8hhZxexCdFRkKX0kBSvOEXIzn7dUdgCR33/p8lnKzGmaSXO
C86POwywoctyZ6bcIZdNYwf1rQBVEJhnKv1jzemdTQAyyQc0jPyI/hCS91HnK4y/
E9jkkDXeG+OdQWYptW4I7ChGwwOgqCKHTlg0ffznbu0SC0q91s3RArl8IFt09xiu
VrGhdPzmQkiiNNctITrk6HyYv3mfbv9GppvkBSgQx1aLf30GMiFMZ0yEOr8dFO6O
Xt1b/digS56RIFobdQLnT8czgDkPtNTENv+sxJfB73q2IKQldPw0zkyy30rq8oQh
XdZIkKXF5emmdS87HEh/0CfkiIXIVsrIQu9hZ+f9qfHNnFYfrxGdb2cOD8bpRvwr
tt42eJklEUBKhyHpYHwpDqFntu9AdondGLGh2CiVDTvbOFoGNnYxntLrwFoNp2pX
0O6SuojebkFcfGgOQYsYQT4fEWLtkRmnyd+3b0xbnoLtGT5BIcqce/o6Jxc6XsRz
FPPDvKATVEmkpvK4Yx2FOEmHeST24mjpO/8py6GL3pS7nooOnGzv/Fqf/Rqd9pqN
/52cL3e9KSVvXzXBlSJqScgnkueFIdwMN20t9cJ0FUZ+PC/hFnT8DbGXp52GaXfr
/fSkGPT8fxFaQVgj4sQ38dnKZBAK3UaxvEX+GQZgv0en0JqXj3MULdl2LJe2eC2D
8M+cxStNTfhtPPEC2MCQ1VQCG4/eLVhZStKCJO9XOReP8gr2bV6pcOZYdLjjhZxA
9O+wfnXPm83s0/qscUqnI/T3PnOEQBM7ijgQPxiCIhWkN4SHP/1GaeRn7FpFj9ry
xhc9gMuHWQmCRzN4U1rpdsBfaMsq082/We0OZAJaY8zDY5v9OKQFAaBHXladK18c
f8nz4WIgiGMjs8lcE88i+JLTZI03fDB4sCLL25kPlcTD5015tpXGA2E0PX0TgeNS
O0I795SAcHa/C40keKrXTaeChAUNIg/i5z5PIN0nHy66T/2BTvJDpWIcJDTiYf+W
xdlBdduRbeeYwHJgGongm3OVQxWRNUdxGQUK8MVony8742FbC/O2xKd0CNOcugL+
D8IocK8DgTKa93sCfQS3OPF289d8pcgdlQRolJSi7Z8otO8W9RNnZ8i3VwBdOzGr
qDmg/GbhpWEZhfMbOrNtaKu3Q8r3YjTVEH31DTOH1QH8BPWq3WrGWWJ8pb+m04l3
rNdU7ckQPUuepYHh2ca+fi5jVZOauYrW2jZKvSnX+liZikNfkrrRMr3/pi2K62tK
y/dXBv7NHFXWUElrKyoRCTE6IdJqfL5nvrStHvDneSUYC93TPC+lA6Ayb9q7CzHC
p/zWwQdxtQqLTNmDo9beNQebofaXbPbHQt6xWjXs5VlfSzQgm5QyJei8nkHEHhuD
vtoFnHnmcCIxRcaceyys1ShS0ye76l9hyJ4ngd6AXpKKxD+XjNKh5hq8RqSh5JzP
D19K6ofjNOZTgMVmqv1O1ull7ulbZfeuP9IOByTg0vEfQL/bLj/7LgdcceOcM7nU
cNnWaWtEa+I/MIFQTlPoQw9vJ816UHlvRnz+ABWFBF5MplLVyB2KsMbpdpeNm90g
zM91ga8cj7yVN/eHMyf2vnaMR6afsMUERYJkyuWWVM22+1KdJRJ1pofPWmbMGNlX
qGhW3/Ebv8BLcyEBUdqY6H1lm5Nz1mN4/1qdt2//Rt29gyBSe3GxEMoI18Azcyo8
aVh5i+KC88g385OHHmkxGv24PsqbZXhW+z3sVKgyHKEZXq1QihVrlsEba1krBUkp
HAhJbYH5chyvI1uIZioQmrpB+KAJ41ZzR68IksLXR55HG24sDfv7oReqhR4Ttyk3
6m7/zEFpyeUkwL+5BmneASpkMPn1lT+iAKFhWHwItd73iRuhDJSTjWuPii2vM47Z
WWB3gvwBOgMWJucVFBrb4BealRLS2dokVbNzzbLN6Pv/Vd/BDzRexbBZ3yQOtr+q
gnwEAhVoUGYCviEYtwYS622+xop/66JklRJa/iQrN3mptSBsbyCcYrqZdN1ya6tM
JcOfnItea0X3dy7RUFjrmd1RuEvZYl4I6Befg9/bMWRIr7xrKvtGc+ll7mZ+Kl9K
qFMc2cBFoox7sdmbCSPqEuIk3wI7NEaqxH3h3fokJDzBBSd+TFwoz3t3WzWwLJ7i
CDHy85B0HFKjEiDoeikV6p5GjkYH5haN2QUV/RqYf2FBXG/QF+L4e7kjFBLI+mzT
fOh3C9/9ArvoNGI230hXpGFY0OOFdrjJOsVBsAFACPOITNSsUBdDbUjd4p7kTDpV
hM1K5/mG3hicLCPPBBa3uwVM/4Vgh6bTkcI2sxJv00JLwsylQ8axI3eEJuHUuOB5
F+MZRkdaXyrfkvHDbF0wpKNhn2CAEyODvu1+N2wvSSxeQnNWfmCkUOcXoOIYaqCd
CTdhHnM2JdHQRdUfc+vAGlMFGYsgtOS2W6Wsls8tzn31M59bMnKAmFfNaTxba8Nd
s025Tq6ffpnF+5+6xTUC+abmORAgCQ7dH1GJGOQeqLtk9c4gV6LQwMC+R16X+r3t
UIv2aD75QmTVmnlkNgWqVHGtsmv4RntYHfUoQzpoIwcuqoWEK6S2x0Ug/Cb0dPwF
JL47SBaqhnf6jqsCok54v1Ad0CJMopTemCJVAMBTd28jLdSAf2WCK7sP3Xe2QwB/
PxSDuTbFdyyoMDETErfJmaiN+opFbBUiE795HGvcpj6rB8tI5trVgKXxBv3rZ8/h
gd0J+rESz5xyAaHKWR3v8NYqWjHmg2T6nFNTNs4uMb3cv6kMJsUrM08MLNtX4xWJ
/+LpbmkTjwSVQb53jv0+KVzWHfAoTZHTbfTOzfTuI6kqXcF7A5PBmew0KVXWsfxF
iRTq2+wBRW3SW3WqepnWmE3Sd3Kdm0eN5w5bMuWwa10Fz8CUaC4B4D7iBMY31Ktt
74lX1P8IGu1NbVA4APqMo8sL0aOixbvmIv+6c3x+mXxTIooC75P6C6tKdhWe4PJZ
ATFThuZlsbA9DAnxACXTCdLvtLJg/TuMncZUYBT38X7zUxoTYNLqtGzx/WpxoO4R
/rldCVpx74ZMj4cHvXS643rtt2SQ75wXbsvnB0gaisLXcauGSUW0p5nDYByHqV0K
uw6wwOQdS/u6/L6Q09MZUAvVqGiwJ7GMducGtu/sS+wcokpf2FX/xe0EiApWiH6e
W2LCvwKw6Nilbz4yVl1moIAV3smvM/UgHkyn4lw3Mi9hvJF78eXYN8dlWLly1/XJ
pGg1uNq03Wcp7fvx71ynYbNVD4RlflVAmz9lEvnAj1wk8ZBbdlsCK4eUcMU6sX8+
KRoHmrIMU6qwSlwasbeYuo1yj6jWkdrLgW9EP2So0udONAduHGhmrMGV1z4YTvvx
AkF0swOVNugUvP3HufzDOwuN0CSkjyevJay2lZI3tEWkEqALqRhMsfj0NzrDWvxv
mpamXgIafyUOgQeUDXs5yXkaXr7iqhQs2Kw18HeNEPlRqnmpJpzk1uaJ9YOTeeKx
7OMGptxToJiKf91Vcr1Oz3gvVHYMbH2HAcOEnXF4oeB3dCv8wNz87bH9vZXxOShQ
a2oAqRnNuJj0DQOQWmt6tyQGk0EG8bsk3SbtzJhw+Aa69uydyJWH7Bt5R7/bgqTd
YhLBV1Je5ismAokLeilRi3v6dyv41eRQZ/Fxyzm/5AH28rlIvtTqpvIQR35oveQ/
xjzd+qONxN9YHEQ/PUzeAMJAGhlE+LfRWGxUFUXUEtBSdidL5b9VLEmuntMCYT06
kzcFWOzogNPZc/qavpzVSXn7TqixhRCXJbE3zFmO625wjvwb9MiV4fwNMO/n7hp3
u6pVJsij4dyOMtvuw2ulZAdgm19TCrYx6yxd1SB57ljRPBbYy5fYFvGMThG4EXRN
psg15fgjQTr6nxKPjWcmdj8Hu2IUC2lWfUIrrYKwSzPdwM+18pPhHTZcDcQH/IwV
XEkTJlxpFqMQ3TAhctBc+FMP/my8oAArR95WIfuQGXXgfWN+WCvBScFfX9ic1xqG
/gB6dRrARFVXTsOq1MbRoEJdKM0tptdWbJO5kicxn5QnSAaVBa0wH1HljGHuCGQy
Ytll63/SguHmumqwPwA6TEsKzUCJMc8C/HYA8Pc/8rciKae3M42s6RR1AuZQtm9q
yD61TskJ/A25iiTnI42q/qC1WW8Um2oZN6aPPcCTnWYbNpNuKAD0H2jTXirYW6W9
L+8l+47Vog64OmhsM0uGPuGFqSEvDvjn9UDtzcDtyRQvxj7QNbVrq4PmIhQLgpK2
p1c32UqkOhdKpmMgJijhHT3yIUj4xiq40XagjbDInT/GwHJEao25Nybibo+15EQ8
cZ7+zEjADLcaPah8t5DT4Fingtw/KHuoEDt8yjIJXlqav25SSYsr1Jw5QA8iZlEf
YHTSqacg1bLeYjJSTkP5qiBDs1nheEFoBroBoIz1z2wxQ4wfGW2yoSErH2yUuVuG
nHOlCqY16x0zTGphZTNziiwYO1nHZAhJd9pqab3S0oEKQA1gOcQkb22vo/bvriCr
90WaMQ2B43jrC+LDZWxeUVPaVn+gSnsU9cWvfk/RZIgAcCclHNN2+NSRzNnTYnkw
ldFTNMP0428aQvQJugzUbM3kkAwmGNGzQ1s82MGUIZSvYoUbYcb8TQ6wBQA1fHVX
jcUgl6Bs/R2t1sUNNQB82NtJ3xrwGY/vX+1JwkKHPIItgL35kuUczDXEAtthzbA1
i6mQ9T5iX4dwNlZBK2n4g7XLpC2zVwq9d7SqIQuBHeX2W36Rlow4rfBhQRGLL5+P
tzrutgYDx78EDYAxtbvUeNiDt83fPqNAJRW6Sc5VivvQ4pCHT+S6e/riDgDf2qjB
nKxcvD4nLRoFdI9IrRRQDRm4x18KLrOxYb1QSjnBcBHYe1i95KrLrDH/T/tisEeV
c//VEGNhfwKWdf2O/ts+/T3lnL01UVdLBcQvJvACh12ZCPrawZOfHs95rIibZ46X
7+s8kcjpna+VKCi1DV4TM6swxVhTfvNl7t2y0uHPOchqnXYXP+4ZNwU1KtZ7nCUs
yqBpKHfaPm5TRUZCzX8iFRr9FxbU519XTCcTNPZcbJdhlVBjsBXUwvPWQf9O6mEP
vjvnJAFehSRPZY7SVdaQxrPvBA6bztNCxyX52vF97YNdSeqgT2sL1Ay+qP0HmRc/
JjFLXXWRqiFgcw+sAhxNw5mi0HQucjJi8Mdexsa18luubON6NFauF6B0smOW+BNI
+mH+ioq4AdwmPB1ih2Qnj9VEnaCQssVMoq7Oo8rFJtomQorB5Dd2Fx/7ermKK/OP
GlyXdzSLfsr+2ko87ulDJeuEyOeXcP/vTgXmeuPT/PAb79Frc5OW/3CLHj4mxFmb
/H/mKF8Wq9vxw3iZnVRmS7QPuwp/Pd0r317qv8pIEGLwL5d56F6XwAB1sT/jauts
uqXnT/2LbTrMzJO37P4Y39ig3lDfiMMCOAxnivEsRspEeALIWKmQyWk1WQ5xk9JB
C3BnfdCtLAwfIjMISbyJx2J4/dQr8PsNXSCXaTMXIn0JAL7R/u1P2avEPgq7STYq
MjOi3GoIT1TcwTJ01414K3bx3/d7in4s4ovK3+aIj7x7IUMc9GpIIhv1TizAuKbq
gkTdHRhdIQ+1UVU/Xrh+0tXYODQyF92c4Bhfp+4kQX14+JAd3/7yvu3aIfe79+u9
Cc+RScNrhzO4soyGqNOptkZSgbCHekqzQjuHaUZ8Sxfod5EC2elViDqjjqIJ6MSi
q3S8KGoe6dGzLVb2K60sK4oY4bx7yL+oV1vVHOz6+LBMLHRQvGZZnddPBCBbWupC
s7lWj0EqlKj0xKa4IR6hRq+8njNwdZhAYW2xCkdkncTRRx+UinGDGhHUVLrPrWxB
pPNcDpGyz9mCRP8oLKh1ngRnFmzya34TQNVhTH5LIjV4ylDF6oQxHkjTPgUCLR9C
lrlcQkbor8tQasw+jz/yofdss7M3V8N8gO31QMcF3GovQT9248V3kvQ4iEMAcB/2
ZA5bczzZfUFery4KfK8t0/Y6MWBW41TsivFh1j4auaKOtCBa1JXxFmPRYMAP88TC
3uAMSFV1Ah1JDv05noXPNixKNJkVqh7OWEdg3TmJjBY6w/97Jn6q0TgrCK4ioUKf
htOCBdEvP/vlM9QjC6OoMw4VFE/mu+tXUfWQ8SyAtRG8mv8BTo2Y4k/YuAwD46lZ
a0aZzFOY+dIXE62/IkuI7XL5iPKOnbxnrgDg/W7bRcZcl33YKaZcF5Vn0cQgk7J/
bMADV58xzj6g0S7Nx6eW4dH2SjYMKHVmbUyUOczkW51nkfZko8PgemNdQYf2Hcdg
NNX0CjfyEtQ9RPbfHoKuh0FKV/ILajzLLvYz4a6FXSLCvsQS8XoebvR3h/ivyWWd
9R0ZUiiSzoHuniZOhFj+CZZK3c/TAf99Y2uX9vUEn/oiQ3XXo6MnWieBw8CEXKCn
x2DbSrONcFm2RreJm9ESAlqLLU2ufQoYCwYgoWIuxIIqeEPuiHugOyuHJLgQPJYS
3ckdHuF57suA1xrGxau/ZAr57PKxptwyS0Xd070Ez588dQ/MGtW5qfo9mIevIZ3F
izIq5VFQAHuA4mQvd8stdt/MDylE4u9v5CfmoOelIgBjSPH3YMhojnwn376jUH9p
0g4+eDvr53LwYMfqvl06EMRav0r4rJRfZxfJk0Ci1eAvKwoswisBEF4qdW9V/dhI
YBCKl3w4BLBW0hiFKXx/2JjirMlPF6Hcvtecwg4NyAzmdguNygeWuGNZl8w0YH6O
ZEnUVbYp3WX4nkHlokmHwQqvb148i5Q+I9p9dd/DV+hO8IOFCDFkIP1Nhy/bhGFs
ZtbqBpql58juklkscC1vRJgp4DSBC5IAWESiud6IeIhJhfYIVdQHGue9a0GdCpg4
QaepHoPhXj4nfUAlJ0c0gH9x/CpRS3toJ1qQ9iKXwcrmOnbzcyctzyAuraoAxITy
ImoBh+PUWIpCxOO5by+unAx1oFJspSj5tzeGMyri6ZaOA7xmnDH0AE5LhKvjrYW2
OM6BputVBg8XtG1++mAS0qrgazjPIU8bNWJJQZGd3A5oPRIcvtr8HP2Kwh6DCZ3K
08FkezeUTzV4qoSap6ICtYRkymAsfh8MDZ284d+qqlIFuHWY4xVixao7lfdlCP5O
xmvBPAc2YAfQKoVm4Srlf6z2JrXjmAD91Fhxvp9Vi3+z5dyVP+3ytfUkzly3APKS
+HWzOhA1iSTqI6jxNJBR21aJ0PWVG26fqGi+34CIE5uTtJEv1DZDAft73iQuPXmo
0Ue7AEKIcmtfjRc0ujYLzIjR8nJfhdbj2u17uYTZAGfNb14rWzSxv2BAOeX8MOlr
gsGMnlY//IrnyfS9Kkik+/zUs773zXwAGVO48VFQyimU+7V3pp4Ic4tkdivro0dI
rd8GPg71yk9/frreS9yaHAuRY12VDtgwTKqTH6yd16f6529O9IP4Xr441MWmFrTu
THvPnMM+lKyzHm93Wa3rHNMyh4qFlLzSspiBFOlsunVlGuWpeRYCFapF+MvACjMy
A9fKCHl1maiDLsebAfEnflOU3h+yNOqhw7U+bPKhj1tGRDNkelaPfHy2TQQ9Pbhr
5kYzT0VG2KlRyrFvUrnzB/CjVWP8bucYlgcIyI2oiH+GiF1v0lsjkBbzRXDaGCZk
5REVmkQ6TThTeVoBCPeQxs2YLD7yGuuHazjPsLDc13nrHQiN7mFAU1uM0iM2VJSS
ADJo0HI/8UBGhHm1PLk1Hzo9pmDftxH3n/IoAAX836zDfmm1BEpjZk8jjRaWqZ9r
B2bkkcFqTnj5lI3wCx4o3/Dcr+DbUQdckIFIQQfzaTxpCaQxN8PELzcbcqhtvmgw
U94AIlxXAwe9MUaUNl+2dg/MkfGLKNb7Q/DICmh4XhRlDaTZAIhnwjXwmw2xK0dp
+n2+iSynLPvLVW5CJhyXlOesMyFlM2gT2TnbVtqfTfpwGRHWTOriE0DT+2ebVfj5
kfW+/bURi2+YmX1hbaeMsVqKIM//z7aQa3tZuFbgWFpCpfQ4QNVhF8nKTBZkWeil
P1hJ1WC2LIRncYKl5VEy7yrQ2xlJNt31lmY+PknYVG78O6xfFT7jJR47YcPjPcTD
62gJK4ZWymtr8sFZwXvsAnMsHrjpWWexWSkeRCBIH1Q8gssJFTWUWue4KegTXXrK
u5dS/RwHTVYTaPDERvq+SQE3YZnw5ZkKG1wv0IGnhBAOxppU/GvUOIlwYfeO/zfa
QpIvB6T8I/u7s6kVDJbqCXp6tADy7nZlZigjpxAhSAN2VjT+KRmE8jFvT25gJhsy
CbBoxA8OdiTWOmX2XrEEFu5hwws8DvlIWBe2O+oeOdfDEUAxRJrURzx7LF+PgrOF
ugEqpAvuuZ9NBtWlFQYazRMUdKj3LhwScBjPatb0C9RTqP+k+HS4M9JjgH/UQByp
kDTSfiaoAy4dtFJolwRjZ80wpPw2+1axx32G4LQK2ntKnQunpppgQtXrJDxCgVgg
BPNj7EXmhC7GX72i86NBwEFFY2Yeg0h64VlL3r+bqss2IyYsYthOqO/o71ciwS8i
AUVH2dzu40SnjNHLSVCdAaLyVTJYY6Ns6Vq1y5tN8wKXe7BXYeKgAk/o2WahMOYd
LVPORYgn4R+FU3dXyH5iDppou3Q3eOpXvn4Q2qeVbEK3dPIMYrXdnFfzd/9fSaFM
waKMTahj+yGGTiF1MxfULRmeMFGM/clkjlBb+L0Ba9UN0r67Mkrq1R9OuACuhVnJ
zIWfxnMBkcWAT/qg7+RnRIkGmT6pRwlhYpEUMvW0OBB/4yh247m4VuBsy+IeF4Wx
Vt76EhEzTbJGqCOlZGslmyZRYLq7eiySvDnYVCer/oVWtWMZwVACLrkIGs+JR/2A
BLrbRPrJe/JuGjY6KH5nIbsF167tynBAndHoqVMafRdEAQC06U1DqFIW+WPLX1Lw
whlctkx7Iprmmk3jJNyagqjBNte4VGZHAqZtTH7eBYBLANsuOqLRtpAwLs3o6Gxf
JSAb8YCSvwx+UoXrRtGBWVIxhkWKitJRYhOv649vWnebi35o323N6/y+hkP2NSXg
wiQ/SjvPtTflAqwYKBc6nhLYEtgf8TSVbMV5FreuUxy++bx6zO2r9j+UgN06hu0S
+8BiTsSE/9XP1gW6TLDxB5PqGuIkH1eP8LhKhC1cLLtfU6+ng9HoET9My0P5Oc14
+bFd5X1xWnQw6hXBs0D1zDj/2UKF8Imzg9mtWbbZ0MaBGYbGm1DByA1ivNShsXk2
01kADk/SRizR4pgavKv7wxwJnW0PE2rJnKXTwprsksiqxNy5IKAkUvx/abn/79ci
YQ+sTMdT6ICinBXx4TKf10ooNgUooIfBgRB9FH8YClTu7cXY/fgz4zDkVO6pOHNs
p0qLKI2MXPiRR518syF4kWp09VDOeArGqzkKrk3ivtLXn1xp9nbK8F/fLML7GVq+
GSAYSrRbB0TMEA9sRdRrpxFFBRolq/GwI+S1Ny52XJ5USSIHawzXcF/XH8pzThH3
Nz+Evj8qis5zHeKeQ/wvS6xZVAVkTpx5qDdzuhpwgHwfuwnXodZc/sLccHQPr2i4
vfqpHMrAv5hcwXKD8wAf3szE710GxvpuaNUdaE4w4n54L+C9npzWtTmms5CHxnSI
DPbYZUZ5nTyhlDKSKQVRmfC8m+dVPEfScNttAiA/13PG8PzICchF9dsVMv62Tz2K
JZlNRJnQLA8aR5ffJQACKlKNQcTqmzQgoRzlLkmvutBJ8Wic4ZcuczP11dg1NTvB
RmN9eoFzMtix6pP/1suk+tZB6TwYgAgHL2mhUkdEtgJ3A6aBa3T1P+ORnRRbBdv6
ke7bYfWtRO03UbBaooU8eQLBYFe1F+NXMQY0P+xL1PI48mC2m7JQ5JgVTQhGNabW
pZy5TSBqivultNy6C1WBTBq1l4zNAOgKMQBrHhWkOwGHaJH7Aq3fpmQUEOcTrIoE
t7kqYDodKjYGZYeonoDJAIjxNb2cBJj9tB+aHl/htw6WxBOI9kDg7aRF+eIAYn+6
SYWaJnT9vlGcMQaaV49Oh0FUSvhNkPV0amN8x5Hkj8+268GjQSVsRI3ayhXScSs+
5oh1V9AFk7ag4MiAGCpmOJ1yZ/yk+H6teaR+1MphhDosElA8xvIv5dfsW0Bo9+tQ
OSJCg9LGb4zBSV5MpF5kh39PHzGi6961j7jUw4dtTv8E9kqXNGILI7OoynUfKJko
OWRZDx/uPsaKqU3o94opUPe9+liXqfOItE4S4RgSEhrQOUYDsOm31UbYphfuId4V
xkKnQVK6xlvD0Wb3m0sWZSq1kT+zci1ofey8Mb2RlzSbDzJXES73wkn93BTcfwK6
c9JEBhthtdfCnokxZ6rYf9yET5awyzlW3Vk/NGUqGoP66eG/ehnL/hejeYeyrkVf
82c1l/EXyIld5O6bXDmTfoX+W7pAXfPobQATOlV1cmMd/BtFmcOP0+HdfBfKE7yF
zZETGVBCHkFIMYFJqsWCEf3sRdBYcVfrPUo1kFXpMZ6wsNZbY5iRsQrtZaw1AreG
huBHGDY/AcTAAOcv95ZI2JxCWwQySW68RCDcF2TYmw5kVFZztpRRgIvP1dx7TunV
gg1V45Eq1l+O91jXkFeQnf4MN/+G4hUp98gPvSUKy7JlJRanAqXC+D/AK/dKclw0
J5kOui6q07xZKPT47HYUlEbmpA/LK6u8fDgsUeL1mHI8RIT29MFn+NEdpwAt2el0
DzSyebMAJNm9FKIF+FPXRN64hqaghlIE2OAndQ/WH9q5F6GxBtW19Dl6QRf0vJyH
7PyUkVHabU+TOl3WQINzZAVAGejCpie5bg7hdvxyJLcgHAmMZT3Asjzfbp97EFYX
aUtuGLurDphtxsKtEZgzDTSDJbkGBti2sI6a2iZlP755UBBtIICgQr40JkEgKk1D
08Tlzdap0kV0qpn64pIkmcUmgu+aBcLir+utLgw6OAdpRdwBL17O0DVu309gqxfs
fSbb6TASW1c7AYXrL1ydAR+tw4eQxQsvtGSrd+8OHPNKeXueNZL3kTg2BYSZu/rn
GlTEgLJo3y4dKMYaeE/1ECmNtluEVPjjc40YMWcbJzpYHGlqc0b4Hs6weZ1gRHAK
yOs9z3aSpA9jM6p/v+RXyukvHYBuDQDBsHAji24YsT7m9C4w+G1CeaM4EKpouY/t
Hgi9QdtCTI1Z+LuXnYqBm34h6dc8+W+hyJ67ioPJOqkfPYB8Sn/hyFnjqvtVMFjZ
XBn9ERtBqUW6expu0nlVX928r2K7BmQtU0Oio95ryChi8a7LMNq8n7HMAQF8Aw2l
nxHIkMP5n5G0xohm/UKULBMWCNhnSN5+dsy/GyRn7/eRn5xE1/FQ/OGQsuYYKPmX
gHdybsiSlZWsaWbhufEnW7BDbkrvASO4H2J8PNupZVGy/pLt2zjUHjrP8KtAlzbb
87+1k2O7T9MkGdGL00iW3H1JLLi/vq6bAFFlkcKRGlANhV2uCrWSvTR5QEMQJmJd
HJsWqvO8zozTBXkUltLgZFVpb4lVUH2xhk9hesHHkrImeIrDSjSsdAooWaza0oCi
LOgTct33zBctkS560y/bezNu/IbaBj+sid/f6go4zfJ4zrVL/t3L9A8zlVwPHfUu
9xmMExeH0QRYrqHh9AM1wpaMlLGoMPXjX3Becy4H4i+AwR4Kj8FpjZQcDuvfUFrz
FqM6sSn5VJzDZQqCUU50eCYCgD5eJ8h2YMsOxWRzn18yKHJNVK/yUVeUg8266BLC
D2aVj3m3rk9KFvw55Zc5JCGK40lih4uuRcPlhK0AiwJoYhYxZ7YXMwzNKohH8O94
5Ik9wCuNBwrMsdHxTVrdpzzY5Sbj87sh+jz/8fb1Zv5uiJzZqsS5ljJ5egCVPRSB
RYdOUBb8OzRn5P9ewKTtwVEDsXzACR7K5jgjWlhV5shS1e9aqImeTWijSUk2gW62
SfDGrhIe9vCcXH2LaAYFNdctxkVXgV3IVEQyk6TR5Ikgu9z7t8cVtdNS4Y7JAlN0
49aNDn/A5OnPLzL1Tv2RdlXTPaevyharetBk+FsrvPyKGHCOS+u8n9el5HZb7kAm
wuvFO3YyZqXAVM8ssWOIVFjqy1SVyI7spm0Z+i7av0ATmyK/lpslddD0bcZgINSo
CnTS5Gkb+a8jJO6uFT4Q0srY1Jg9oCD+WDUW84QaYMQamaGtsQZYErYzGXn6gzBy
M+zB90nlC9UMriJVABXRj1USjUaQ3tVpQIslfjfCyvGWRBJhRRjV9XfwAT5YeyjO
S4bzkAFtXzGFJ9NprrHuq5+NIgnKN04tHIiniR1Cie5m/awbtoCnwrxbQqxAYJaw
1YDnRJ2MZGAdGrb1XOZ3Dj5VMfBq8TfC+0rxUoolCiVnORXjVeyAzrBl/JbmU22w
TQDJ8sRoilZCkIGv40iD3UCBkM74UXmWuGlWVMlXz++RsKy4mdqEX5DNU2TeTbJ0
OqZs63sinX3PRzLPK0jBr4Kw53pGNvR9swGXXSi4oW7zPYGimip+lMM4bwMqQKyM
UGmE31a1bm1pGQX+NU4LIMzY8wEaH3wJ54PogNX6UrVKnU3jGIcQmVCkESndLRmI
duq/9JDn5nV5G6XXwpFPuA5tVKUBxPrfvZP6nV3XHQQD0z2NCOX3IhHs6t48suY2
k7JwtoG8ipbIsOXGyMzTZwJMtgdwY7D2JBSPy910TyLyagBrc1AvIwj5fvdY+7Jx
g3mAkTTuGgA4BAVxa1sjU6s9+CDtCYGUpW9qQmypbDMLnEVtBBgSVU27epMKhBzW
E+NrIf23lCY+Y/P6OoZQICZE9Hop/Dpu/iqge0DUvPt2CehsOBzgzNxXYUsnfdgj
QfdBTaVqjbv1ULLjsP6BDc/7oYzyMFhaCjPL6xV6abod6s106R/QcIcj7w/NXOxM
hNIG90mb2mIQgWO9oxq3EWWlUH111kQvyLNxVWAYuKNIH1K7Hz/Z1EYv1jF4BpTB
S1u6YiyDoDphb+Uz6E3HAHgOd5qHRZTbDOtWE/x/L6l45TAxhyfFmbIO8VThxVjf
jk0+Ad0qWX9tnWErAN+2f1ozIpOK1AnI0Qbtd1Hym/pgfN7UBdb48TlLzeVkiuY/
gc11zFzJckIXA6hDZKVPka+gUWPxj+aTCE/AFFpL4RcbzH/KHY44YmbvJj1Kq6O2
R2GNBr/mh+p3RTBtvn7iiQC2H9j2hPxcy0TSC6g7pXZelehgN0UfRkmXF1LziqAr
nglwz9LfbLsUvXPRJvGK6l3K2rFmsnEYNGOpWkODMVn+CsGh3oW2Mbp+LZb8q/sd
G+wTXL63dQiXA+C0HWCrIKtQuSZET2ey7HI9yiZ/6cnllYnZU539Ole0f9scBfRG
XHURxtNrsGR5oU0SdlKefQWSn55tWcJVjfS7Lpbsw3K5P2bGrCioUGclCAVshU39
yMumgUYTGZvcs4DCgtlk3BeA3cVDPWl/0lyr8rVe7IFsVKFqkrT3+PgxPN4gEI7o
4OdIj9OY+snETxePG1toomjwB3xEDsBk3P+gY2lBGCiGqe+8QZ5Tfp8W3SIJaRk6
ljXHR3bPODTdcHA8ccKBgeH3HSAZRFbnE/X2c/8lYv6gMJtVQHdiocSafB1SW12i
lgEmTyGle7lKpQvPVfwmxad6g5IfQajaEydj0OHnm23MhKEh3S2+p0Mh93KcQcfw
ZEknP8NgCj7G6jX5OLplJJ95KyAm8XhgIx/A1xDCCthMdY8SPRTNHVAFg+y+01U0
Kx13tH6GjKZpHh/2jQYFEWP4ipnWPbbXZT7jZ1zmyX85m66ydzLiIoISDuluN+qN
n/NKJjdXmmj2WfNk3vM3sQecGkg3ggUCqLVtA3UNdRDTjgaUQtlYY3UAwaEjKtis
pM7mdbW5Gqif0w7gTvDq5wnIAIxruYA+NHSzzX4XA1+Ca44WzlxSRKcDjYkN+S5C
1kuQAc/U68n4jCvIddwTFCvs0SUZriKJCaLwVsF3xEF2slqbUbrRSHau7fkxpapf
is4fYn6qcMkcGwcTBkC6WxJxCtQQejelp69iZL4mSOFTzz86p0/Vq9BkIaSdAroP
5Sh/o+DodQsSKWgp8XMU0fEh3LGJvaMf0q3TqDBFwvPI0Gxfv3ssM30W+vHNvaZA
DE+JjGxuIE+poxif4Xk3jC96Vyz7ZfNGI1DiaVBqxETp2jnmWf12SJimwt839n/a
E559MDRnm58JdAt2JVvmE0i+/LMjyLZuOOklNaLklnK17+X92d1KH/5Lv9Opitf9
ja/Fp8XujfqFt01Pu11qSV4GT3R/wgAZ+kIC3lh5+5ZHES7cAiGZZu9EPkb4vNX4
X9ZooLBBd2dbDeQ8pHhHNcGqDMnTB/pr5vg0NMJtH4N5TRTzmAPlL5oMsaCFC7iy
raOx2ay+Hc/4Iwmd88zPAf5r09Z5TRCDIpFTsnSPIemlWq1RNZHrZqBNEV9LhekN
nVDitefke3flQu95A/T66Bmb6rpIkK6TJTiJo98vm72sMCW0U1xLJoDUYq2XG0++
o2hv58hrTwllR0RN8phOQ4r6hDSXom0X6YSwtwGaUfd15uLqvJhipv11iGeOgqJx
bn0hT+WHn2DPqIvh2yxSFBN7czFQ0/jTTARkEEldoNrq7BrX0CzWnvvFFvbzjoMl
7qibOuKjM164F8rN+Aj5xgh7t/uM0BA2DTrk03j5cfO5ni4jOKLvlzi5uz8gL0nF
X8Qwgr3DOWNLNojWFusnwv1W91zLBZOjNARvhMp1juHhJvW6uOlKRsv20qgG/0ZL
YlxnM4ZnzC5jc+NUK14io4eTcf4c88V4erjS2O24DU4LS63H44S1y1pQRfHQAida
TvWTlOrhMOmsXCoxRZXHq2kVcvfLNGhZnhMvBOvNAVF1Z8inHOf38eR0y3D6jAk/
o9fzhRVvw8GcK2OvK/YI75KpNyjQduZGGcdzv8fmeds52Lbm85UzjZWfl/83zG5z
/OTf/Skc7UsQ49VTeFJ4lonOOH19pUi/33TrwOcMuLZyQtAAldej9ReXkgSxZHH6
a62dpPxHPjkPvS3ufsYEMY0oWINZeLOIi4J4qZd5biBCioL3y7mk5nEe+o1oqpSd
FU5Ox3C/Tn9RMqg5KaHdrnBBEn5ImiQ01rK//YOMrk7uGqDvB+iD6XinszHuyL82
qkQczqDhqe5wBgn/pNyNOgJJN0asZy1uqHaVg0T0OWW5K1HP8h0ZeThqHC3iTMJQ
FIM3roUqhTusFM1tBaMzn6s9mk9ViZuSHdCcVvVDeFQS87HgchNg9/FrNeP0Lpjy
Zd59eANTKSKwdU4v/aj5Tvf4jIqjaonP46qF4DSBVYYuWR5x6xaVX+D/k4Y7sXZi
vBoontMdeG1PcAz6v7bI/t7b2nOz6BjCvqfNhtECNP5vA3JCLC3cdt04hwIk5yIz
DfccwtBGOutgXMZykMaHO7HoYSawpFny/+MC5Ux1hIwZQ14K+TCyLGX9p30GiU/6
1ZmEvryytc2EDjJG3PWpX9CRM+NFOMpE/0EtXQeEnPv3VDuBMoKXT4KiGzmHqvlo
C44VURkKrvHnW19ZduhX2xTx0/xXE02GMtdZtsJL6oxRmPiT8M1WNdQaeX4Bmdkm
JWBGpdSKWLgWRe+foYGvXhZZE9b97gsyb+KdkLynBz2ZOEH0dLnwKD58VjYmTrYC
FKAQ1QmefDe1rhYC/MXGXuGMG0Nll45nCDmXsWNmuhiW+WXkIZUztOd4afKxg74C
g6rsObNH/pc69Ix8267hGxtgB3BX70SY+s4mxFS4TjypzzZEUprqJAnAzwbeP2hP
6GKeuinvp3fVMR2ypUrzdpYof6o7qfON021Z0V+Rfhn3LsED1Iifm2lmFUWmH6xl
l7MrGOgCZKrURSmrdl1uyjUQM5G4l5fEsOzshLBkIl4SZxl1UbBdppQ6ZhvgOGD6
DfBf+IE/z6+hGRDKgUHsSsXUZRcGBhnK+kqtZwtqgvByoKKMJ7udxzmeP7MHXWdD
xNygW6cd8su3ELYC9d1F36ZilYsn1Q9Se16HmiVJkWgvpQc0B0SxTsOkupvhIaCt
CBQcguGdAoP+Isvxur4oxq70b710XQO4gAZy12yvCNac+3Fqof9I+BqDlXNHn31y
aB3nUC2mt2hmpaDE6izPJjT/Vad1gkgGYqlfClCyAZWESkcX1T+kA2TqlZO/72Xs
qD2zkhrcKkeduDj2LwJX8oV5Vj6pYRG8f6aY16ebl1PxgqNMnPWc+U0Db3qZCAT6
qdcqkli4iJ7B+VxDhgMEQzfc2+K6e8pwH6CNE7I5ukh+lyge1uWBgXdNJAuzawEx
bk1S0NpkE4vO6mwrtg6eXZ53blt4MATHz6M1Sr81hXmMNf+80FUb7tfRhXvJ0QAN
/U7JB0mM0tJ4qo4J2CpcRJqYFQgzjESZFXoqkqII4fn9rC1qxGJiCbIamSeZKGO3
/YIbdgaMhgEGSXwlb0qJFwhJTvDHgwHCKJdinjFU7qqP8vwdeGJdr5oCpL1jdOys
7KuVJHWy51byMIIbfMbyX9NNm01XGnAXSmdQ8Cem8pyPdqFAjoap5RF4CixCs/zx
ngPSQkvVvXBCuvlBL8nwih1QyZoIhbr/2lIFABJ7Xoese9cYlcI1RBm11KoaKJLj
KXU2XPZrtK+bSyi5ItuiE+zIzCmY5FHholBLdpHl3laZaHplCKHWWEVp9tamWxNO
Phtqd3GvCaO7gXxg2INGS0cDDqt9cORzOCw0UeYsDsM2xsC5ndoSE8aACPsr2B1n
xoDl/q1w94ooxI+ZHcCzIl2/zuXyMWIcVDbFQaR4paMTbJ8wGuvUxSP+l9sZG64H
41uWRLROtUkITLUhmFDYooqvz63jKHZT2ZtNbtDtqScT28FyNHBU4gF4MWxftZ5Q
54y9ZRrIFizo2HJBIEg00BJTYCMaDq/+g1FTdjN0mMVPoCRDjLRoFywoZylhb/ud
+grPDT966//L9d9tCNzXmVb5VqN0i4KQwaj3HW4g8LT99m3H4zB5R11G4EuVy3YC
EgzoT1dgsjB8T/u9QxXXltjLlSJqdGcZ9gwzNvUqf5bUGr8L4i/0fmJQM2cwSVOs
KaM2nLYDXOR3WblRUd4J0SOLYkd7jstq3y3Hnh3aQPG6iBUxKHX4rp0K5XCTOzT2
izPRzvCRSW5DMPyr/dCNGW7LRAAE3zdlus6IY+rFscUGFk1JPqXHbBWuRxPLkJgU
LXvA772wd+dVL4ZewTYudQYDjaBNCHykGwfQsjKqofJ01NpiuoOeHI5Td3NOh/Ct
FssIYGoh/ckN6G+e6bF0krT2XMZe20GmT5R0FRE1jxxMSkECXOkthPH+B4J3W+Ch
dDFJ61YKgc3MDIpYWnrqCkne0i1Gj4ec+3f39PyJ6oUk9Bdhhu8HWHrasfLfNWdy
GQt5DfQDE90OvRL3aY1JGgXI+TBOIIJm1cX51J8kHPr9q8YyOY3T3/PjSAyjiWnF
EW73MKUeGqgKPMja6W9oaOR6bCnWcOmdnL2UXHK4mxFK3NX/M9/LZ6RzEvYT1x1u
aQBIJcPxzQehml8Ujx4KBqqz8OgnGSdIZ2QKesmJd5QJ+HrFMgTja0hfguGD0jmA
HJC6YBkLgEnYXj2gKVQ/9u6Jll38TmvnBskhh1ee53z1GN6q4uotAAia2CZ+nQHX
plI2aPN8AJBAO1/ZZZPgPDw9YH5BUXVg3bQYe3vIcVRViM1RfqJV65kTKHkqxQje
i6tUzgkWpkzXPgYsE7GgWrz2cEgryXnb91LFTz8Cds2Dy6MdO7/43i1ZrtmIDOil
BSdoZOuORlBlepyO2W6zCC82mFKPKLNm0ZfSXkumx1OoKZT9zJLvyx4hf0JtKo05
UbkNsWLIishxo7c9PesbnXWeazZtPUCSfiwbbcHpcyAYqNjey5iRdCK5lq2jGS7j
Ljllhn7KnH/T+Mw4TFvLDYpusZhRIJbMsTufUB7DbSxgVUT+w9i64aapra/LS5Q7
xYwMhV6bNCrFz9KC4t+OmIr/7jAr4h6VX4Wnd/8dXHd5WohumqwMpP9hwuyC2Wkt
/uBjT/3xb717x0ho9B5U5yXMkU+y+iAaVmtY37Zy+Qca/xKy1PTi9yr3n+/o5Wdx
T7MMPIy6idGxD/1LrFLXVj1tEQOgCeRswD/5wC/VmOkP1QPWclns8xFnbk9AVNcv
Jludyk0tqAdr+NSHUVBNcqgHU8DzXbJe5P2ueqqFjtuRE8IJ/EH87+0Kekj2kk/S
zfhwR7kKhpM2yT5HGmTm7vYFo8ftCpQdRWY3c7TkABmVvUwFTd8D1lKABOwOCJ9Y
a2uM0SGfzy5NHDkyl0yZHfY/pnNYuLx6GCw/xly2nGnA3J13u6HF+8wLgBhAQfWE
+RXNGA4Brldi8ZwKYN8dtb9MDIhxhtppza5MWI41jagZHwz2WKUa17oOPaX6Ns2h
ZBcKdi7BKU3vVuVqHiOnlBevQVyDhIsEqdnxu1oCAZ4B3CElsS29iklmTDXks0mC
yyEY1BhKv9EARBSCE4zn9mqvBdEwNV2+wLK574A/DlLoTdq1Onp4ImV/TWV/qP1s
JH00abtQ3ySZm6stl9ConlnCwMNT3o5bq/G3wrTX1VGQLg94/x8A6lKU2GLCAsYu
Y97I6Gpso/C/4hFRWyhI063InKkyqbgMUWldBqhqPo04EUb7E0Udq29kwuR8LLFT
lyazW32+aLBb9lFTsMGChKSAi259OgEWc63LSw/RZex9Yh4leWMcVvRbivHeDw+3
8MjLn6zb6uwrnNBoTMnd5icXWOeTInWc0mi0hDARkv32VTF+Xm9rXMzivgRAZH4H
3o/iVIq0HmfMI+oyCacqZLbph1o82Pbtf0WzOZ+p/LQc8sY1BIZTTuYba4t/nBZW
edXxsqzZQYLgkCrllsTDZ1o30lD2k2KolwkTYeSqaR23YCxPQxZu1/zzLkDdhEI+
Bopc/nRzZC1f2P6y7ONNv8iFKrfHmfeM2gsqcKY7iHAHdGeLrpNKmLRzjJtrKWU0
NNfILjqJDeqUJGVWHJ/SQuOoDrx09ug1oj8HqxKc97RxwcYoXFKM9dU8byf+3PE+
8DiX3Wa2tSDuh5bNpyTSNKCQ34xclIOTBI/sTJ16pvmq9SqVLPAi1RmGuXmjZXSF
zbefUM411zHnHoOqokWYexv8M+swkyMSPyyqQrvluPYYAWFHWa96o25W8zaoMUrJ
i/ydX8bUJOQ4T+535PrQzC2KQGSZRfWxZYo7uCWhatu67iAl81v7tafEgioMNLlY
3OLDjwNrAuwJA9EMSdFcHAMOFrx32ya6kwlP8W7cJeH+psfq8tJtCWojIBw0rooG
iprG/JwYTy/W6xg0BkwzwOUQRbfzNhoparN7im6aO0VsyFvTV3lREZs4XW3cXpyX
wx6IoSZfK6mWT7eN872HjN1jTJ0QIwcpSmdYxfWD0JW5dN/5Lgf8RvdjDMkr6CNP
XxnrStejcjJlaWQxACdNvqbJicG+wZJHoVyNyQkAkroNCaeGi+ncWJ6n7nUU+5lJ
mXB3aPX2sDsGjbLZPe6tiuCwPQba91MNubD9qc7ly8f+bhE9uSCJhP/KViXdhnmm
3WJ3A3E8ObjkD7Fa8J7thpqCBcatjQ+zSv1AkghT1fqVGkj+VX/XlMz57rZXkOUF
QQ2BqkitGHsjIUi4hj8FVAmGCl5mZJPL7cfAUl0f2YIkj9T0TCk/nzplKO3yV8xs
AN1rhsTcy9PRgRDG5gxgme9tZJwSn0wdrsWYPoCOzZ1Zo1m7m8Y8muawU1x3hpXC
N1egwM1AMNaoI1zgXDG3UWrpJ5ooZaJyLlotbZjrDShKC3iEVb4pTA0SFeKL75Dy
gD6+q/kXsGGbhW6YLF7uri5um6Cl65PhIHt284Vvzn2KZfqIN6w1SEx1+KTZgAx7
FSYM+5TaVHmqPO59r2o35aHrE4eN+4d4XxhKNrjFHenmK7KPOKTmz38JmnUH2eN0
2ITo0uh41mpGLPIu1iTeghdctEUhQgTvizPP4e7/ifIKybcTYLAHG6lmuzEHVMAC
yKeRAw7AZZFjzUylT6bPCo+3klFHLoRiZYCaKrHF8zyY0rS5crf5/rYyxp/TgXW0
Verj44/+FjAmnWchmzvi1TunTI9VCmXTsSIQTi1pXlWfIAmILAphMPBlVJtGsD57
1kw9jO+r3J0JxC0D82U5OF6SFen+ZJjtkp8HccY17+kqrjmZQwb+GoTVIVt7Epce
nvgEBUedeHQAjt4p3AIGionlsy9SKLtrCPiS0qhsbJdMdDd345KSSMcyGzTt7+1h
IDC7U5raZcj13FOz2itlBi7b9cHDa9WSSPfhlYg8xn4cZPF4jXZucJlCKHvx6Abj
mZH+lZT/BdR4gIS3HnUzU/3CsKqlgvPxF+1aRG595ePpLs1mPmLboqIURIb0rzyr
UNWFLU0AN5UhnywwD6VtpRt2oN3BuWM+FaZEeUCISH4V5T2NSdNDenFl2tt1TOPI
O2FDpnQKz3PjDppXVVwEnEUGIDLarfln9tm9jNnzgsD+JJFUhVG/vh+Aw0gZbFcF
fBEj0kKACRFi9uFapqha3plfPiQygWv/2w7SmgxyuDoCqgw70bkfiTtANTYbBmT8
T9/5JZ1FW+UFwYI/tjEsAiqd+OXwOtn0vg/GCi/KK0+921MU8ln283i0CuWQAuTp
2sBKZ2v2MZ2MRmWO/uwWMiyUe+67TcA3VzRYeF86Ujy+9OYBvalD7K9yDa7NlG1q
NUCRcbcJmip51Qe9He2sa9aSRIXEsNnIu/vcefOMEg+XwXgxpbWN3wr+w3zr6RM/
I1xrOp+EZR7q58mcj7SrdoKi+moTlKH9PFXUVSOb8QhSDJXLkuRY5vT9nOk2xvMy
LGFAdod1KeyvQ/l0iE9f3wWbocuiMTz+02vEuF/PJYOSofSpBWHxbwj4apcUjkkf
YlaadNqhVuOXgnnMEYnLfJ67Qzi/N1O9ys2PWmseOuXQUK6oeWIDMMWwGJPJAbe1
T1CHLrBCbIJ0snq8upeRu+oD7xhexAj1VlmAgb1jWJ+Xc/GhxovGAGj/iel6JT7n
5sUhW+v27dARHVhJcY4EZCJRzwRjb72fjK2RAI4/5Cd1AlqXeGxYL7FjW4y2zU0P
mCv5EERn5pxALExGfAo5Brf7b+2Nu3jLyYvI384s57LDbvKf1+ZQLndYRQvcIl+2
qubpXehd00mn5DOddn60Qfio6oJ0q0GdjrAv3CIBCE+kuM0HH2RetvoeTYBZHCiP
3MpU81dQqK41ltYwaR6cXPQo0VB/+oYYNc3N5UzWNINjLG5zMZpiDZtw4/PZjFSH
DK1v3SjlwA+MEXhXgQ5bUo4/Mw0Tx+xeRG03+aN4kHydjmZOy3Rtvvao7eJ/KOPZ
54LLY5VDNp5ROUoOelx2nHzjy8jZJhrOlMoT378P1zNj5cytsztjYUwLaM4qg28s
kIGzKQTlyKUBA2zpLMBYPNRgDpuNVFoznX+jn0q6lsI2zar5Xj3B9cE6YBne1FnJ
B5L7GN0OMoqUSUHksdkuuhSU1iUtG8ojWuFfKCagoaXr7KipSpSQvjKU4XAsKyJW
2ceLRYLbf82hKZv9bkmEs/peoWBG2AfQiqPP+AhP+Pth6UYmWhOL4BGRJGShXddz
efXFYqGkM6k7oWig9Y3J2YytB6ofDCh3MIOvGUkjsZq/g5P64FTXHB6BjiJPncf7
7OufOM77ZC+OuLtTJnoFWAbqMQag+4p2dEqXbQN/nQOZeKNJl2mkv5OxBDkd7zKu
shrfyAwDQtjWHp0w8pO0GeJ9SxpLHMqdwlsksil35vdRqHFXNHezo+1n6Lya9EoG
/K2WSmMCzUPHTNVDblHFCC/qzN8JH8imCba/9M1HYV13BZUBiU7G5ErUH2Ky8n3p
YJbqUFcECTJhDkczg8gwxcoGCUDPpRSAbg+7CEiEaSt2lvgnMXipxQDfkFQYlWfB
uLuPDN3qkbUcd+ZHkdzJqz0vDJgqlaOKPQMHSxXM9M8lmW5k7MkZviIGOuz59J5m
JbZC9MoBfQ0Ec2dv8uDtIYmChtMtE5QVxbPKD4iPQzAtaXrZddV5GXH25pPEx70/
Yx1iJCxgKJSfllj1MOqiISixudswrjsscB3r60cO6JrKiZvZAq/Ts7ZrfdFsFA10
cCWYBjkwXYgiT1m9ToXqSqJ6/o9ASELG+OUHswH9QmDm2I+GTS4JUXpdqfQSm1bs
gKOr5JdrAbqmP6XxVooeCEl58kPbHf0gBo9/pftWbPNmQfDdyTKsPaRjIEQhZFAt
wdg8VYFQCqEqnbug1VRMl3Ciev1Hr43kzXg9M7Y1+ixK6mmfZElkwapqSC5tTrXt
KhucRh7VM7koAp5xxtwesUtUi57zsBl9BOJErfKCJBC+u1EqdYtjHcBGzCdGSqa7
stfKXQW0FH0Pa5QFM2Teuq8sYBw1wcNG3wN2alZdXfnV8r05iuBK1JMp1qeh8eug
SE8u2ybFt+sxaVcpMy9J8rHK3TFL6SSW2p/+Q8bAvUzR4LbmNY1G3t7/o6AbldcK
22HO9Gn1YjVW6XTDUWFXP92O6hF/TYtGxxBrszqwmKyg+2JltdIeHkNXsmWjIaws
5zCbLHwXJ7xYONLVYUERVlRio6hqwh8VO9iwOZw4s/QdtvIQ9lQMSdVrOABNOWq0
vZ1sX9s1ZhBojmO+SBouF6XZXU7Z463BiWH3cEvFe5gQV9/XZkZ6iTnbAqj75Cv/
Fm0s6fhPIPiWNkN485opDSPA9BD+jb6XTtkP88ir32/cXmyD79VUPcoc9N0aisrK
nr5qOSAkBoCr9ZmzdfAaGP4efsRQjIiOx9xyk+QkWj78PyqRtyLBb8JDuob22bY1
N/crzPKut3nZvdyuVnKknxNSpuPtfRwsOEtBnJpry9dccuaG4lH69kvcG4v32zk3
oLURbyFxelHLgUmP41+RDGAEtNfC9K2nEBQ55a/Srb6Df53/0LNs4iNnFzefUbVS
KycPbCHXogni7Umy8ezCcwWwR/dItArjCInPZrcqhgriMpkKnZeU2kOWsssthOJm
JH7XJ11zH5jaj4+mczOkD1yN1w45oJEWq6ZbRgp5IScOg4rIVX97BJ5yFjeGss3s
39AwoFFXBOWVLGdTSxbtXhdltFjRFq+wZ4438iuzORXcNbBeI4LRCNxWmzLDVPc5
uaFwv6IeQDG5r/QCy6kmIy/hw5zNXtqup5jwJPv2TkemgdY+atckvclXF0TGFs3o
rWcyRh3Eq3XQ8QwBwkx2xD4baCYwdMxuAZCiQTNpNzgcwJzTLEtzwmtK25V9QF3A
RZOdwfzWkzQDe/DlFjfvP4pDCsCRdW5AVBkVOgIAZA6GiIpnfB0lHcoxlthzPjjc
rqk7cmxY/fQD5SUxqw4MZ/vGIAd/twDQglZci/WKdKIKC1oCQTSzSFxNw5E4DfA/
a57v9EqZ1qEliyLQwe5sFZZqotPfVL2OHNimU94o+4PG0MfIwbSoNwXwXDehe/0P
aS4cuexkiNGolgFonLpnHu2oYP+/IEc1CsOwE9lW1GQmmqRg6GvrBCEXbyttRqbQ
bQh0me8LdKx3v2nPpHAYieS4VVZExYdCq4BlSyinNRF+1E9WaOqCUyN4JtL0bgn2
D4vHi3Wu2dC/IxJ7onzL4PnZSOJLdiFSk26bptNYsR9WGgo/tZ4wXn71AgKUm43H
6Oq5mRVr92l1zS5SXWLl0Kxbvx8keLneNHJ4xWoTLMFWbw6Tx5HX+PQDZVoT38Jd
bm+SeZdc4Md6h+LAn1b3O9PT2lvhV6Rb1/aJYPQ9oSjH46uVk4/JlFzO1+PNOpCU
fBKyzupHL+s5QGHmQ9ZzDF8CmuHwi521aX0VAPIpQs0c9HAXQVkuwwqpKDbXNots
oMdH/wrFSnCe0BlsdxwZxfb0Srh3vzMJ9AN0zQSswwbMwe1wnrGZsa6HAoScs9qH
lMd0h5jWILWOsIn3Rqm2SEtGGGlFiFelFrdJEvzYlqlPHz8Duo92ABxgImsLvvNW
zJKn3v0JXurczxR65ssW/1Hi/ohoBw3W9PCmNEcNjKu13UiJ8SukwNvs4Kzb2vXi
qPcWs0MxAUmS3gw7QTSukRLqauGe1/wswtVxcMZ18LRQdojFehwLQt497T2uGu2/
3L7uFrIMjbCCfvHYuPiPpXGlwtTHFzze0Pxzj+S+a/6OePlmEF3ns91acZh18Tpr
y/BlylkJZAWj3dwhQL5WT81OQdV1HKGBATqOaFEwJgfhHD0G5jneBhEV+H8saXZ+
ocSkT22HOBI/f9RUneTot1UhkV8MYbJ10Fu2k1ILOKKALh52x8jLQ75jwOKeWs/5
+UU683TeFiJxVu1TJ2HH8msLdI2kAVwGbK6au0xa6SMZZgvD4xlTQ5Vgw68xWT+x
uxJOHJUsCLXE9T3J0Gk+a8vg2Nz0D3wJD7WFJPQGkEzVqVx+A93s57TGgSu686UI
g280O8hOUVHfZL6kYPwpVXcumaOIJhPEWETcSZMRqXbgJ1lxX1gKojW6dtv54IUt
eLGLscWCHkMw5LNjodC3ZAmpAt/jkG4WO2ZN2GpitJMSQLmOFSobCRkAQD9/5cNH
SCw0l9XmQWRJtY1OADMTi7vhJTD+RpuKT9Yw8IQybbZ5lNfXsmqKs5xuQXwE2DQn
B3M99fErzbzGDvnGifIjWF8jgj+qvLaJjqyXC9hQ6QY08nabClmanWxjYbb0LVqV
qQ9JKZ5QI9GoZc417ONcbte26ZXx1szt8cRTEu1x3SfbAWOECuFuAHTLTeFhkoli
sc1oqhrvqDSGrenamg7T6UZMsSuTxMBl2eKJy/eOBNYleOtcP9RWbewu30WcJZnn
Zm4lltza0GCXGCm6LTEMHjNmuO6BCXisKiQu+Z5JUbe94zohuGHdL5pMBLx8+4OA
IkZD6boJ9q5jh7i6sIoJtAXGk00+KqvClU8BvgQ0d+DBwgyeup9iCzkXHGHAg/xa
GHXf94ytoPz/BSotiewGm9kJA3kMv/dsHrr4MaAWndoblxdq5MBmm+qGkTqgIkd0
sWYPve/3Jj+azHRszMkwxTYiAH2gX/32mj4PkxVJMP134KikZTKWlkil56XT/M9V
Riiw7eeVMposG1hcUr6ygqEh4n31qDtffDSPoSE0r7K5xrVrbehSq/fT+THOukfn
T9LrUj4iVMnFxMRR1H4W5SrMHjSL5B9Cc282uZDAp3do5Yp6GHzBUmEpK91jj3EN
SBa1fW7tXza5NbQhfq7MCUH5n6rK7OCoD1ih+DXoFfQhOt4ruuIrrf5Mx50RQ2zp
pnSLxHV324jmSYUx/AkO4VhQEIiFsBdINFeK6ibaPkhK09CSyHAIlsWQXGJ3q9ik
jIzbZPDh4656A9KsHJGfnfkOysT1QwGHTWYQi1dQEjsou44/kkIwLDoMl7P/XqrP
QvevF3XjzwaqIVu0M0gkI64qHZJaagSG+HylTZkCFwcm9ZeSJlmVk/NfBw7Q5A+Q
okxSsLFzJQ6szb9BcOk4xtWU8B7pLXVMoMXLVqiNa2sSry/21tfGwYPApsTr5r36
cCVp2BBwUxtDzA7+3Sw2vgvETIk2jjkmob7slE5s58MpyDqTmnJOJa2Q79M3jLgN
HobpB0OlHjxlFHgOJeSIn3BY41PL8jRJoI25Ql+Ns0LyQ8zZ/c8LWgppIbYMresN
2mWURfWadWPGofw/zTyjDYLRb55I1OLmuP10FWioK/18ihvw7Nlu9wD7TWOiWNoI
v3ZsYAo+ix+2Tur0nYtWFVYh6BlBlcwCH8A7OXIp8maGWhaAPw0vbw/nhbEQlDX/
tWZ7gzCLtz2xPrJQtnC+LhZXG8BKeRXwQ+C3+nQkD1usnxdhggDTzm6tTDIuFle2
8oK8a2lgb/v3UqoosuoY72Cmj0DYV+gMB3l0o1Ejlq6eVKwjhu9ouVpO7mAbYqMj
h0G/mAurzj39iDO84Ki8d59oIl4d2n6o437S8B8Vmf9TB3xeSwkuCe9NHixfz2mc
ekElRsXq4N4dA/xUNfvrQETp6ajheQPF2sWPCb0Asx1kYC7Xm+Tp+GTw5tu7qScB
Gxnf1nClP2AcMe4MoFQGSjlDQaT2tXp1r4MA6wy05d67phvI/uNcCvw5p66OfqJk
ETvZoz/vL/FdQtLRvGzKGkSw9U0oQArEBNwTDwj6eza/mRdDuriwlDLx65wpr9Y5
BiNLqrS7DIeU86YQjp0U8eRrGFNsk4FlT239Y1TWwZvO3pqWGRBk7cp4kf9X9ykW
UcFCD1g4izWGT39exqRp7s1u+I7Jsac8t9WgKm9EgZ6TdikBDPkfoU1Ano7Xfivk
x+MtZ19b1LmhSztLn9L2DLdqIlIM77378PLphb1Sq79pV/gnJTJCYNprhH/mhufd
4PqUrQIuQA1WzzNUqRHDiELITqEH9+vZDw7LDwRLhkOuH9YF8zVAYiw8sZFyzvX8
RLwAegIg1nbVGrzIkaTErkEzXb9mViZyzZPiDtLSjnPXOe87W/nY0/7hm0jibAic
Z3Ncl9DR6TNsVuIrOAAMTS33FFjbSCP3uuekJ9lGoV5iD594hc/ghhTOYpe2a9AT
h1OZBm4wGseq++aXQ49vqMednWOCmK+wOvTaRWoa59qKBNS797gI+0GS0/fZ+Ff8
GS0OXkK5Uglr3OBssZmteNau7QoXngmipIScc2rkyZtf/Lj4T4hgNBilicVBXEaQ
qurCXTT+lF8a0ZYBy27K2wtu1K0uCzbow5BLc+wfMddNr9AkPI29H6NNGLOH4xA2
05WdhNRJCPU+Ba/1qzBO+e6swShDpxWUpU7ig9oxOx9TdV+4rrvHeheyMVhcZWCa
whVt98/xBYh9cgvnzi+IGZeHxmmxVCWPPIZkH0lKP47jC+yQ+njxN6d+YrG7MO8t
8uIQNq5F9jIY4L02sgroV30E9y0fxxJmnDNrdBDBzaIVcshwkfH9AlfCAcFqgi4J
uQwz5OJD/UxbnWTTL5uIj3Rsdj+tfMe3p3H+GSnM5wsIi7pKyafhtYO5nWaM1wqX
MZH9KZ7cgL4CDUPtvf0aEZYR5Zw8hxDXFnWUpFIHTLD5CQUfVvoGJ+PxTwMcHfCy
Px9Tl3eB0+KUqg5WLWP/keHbQzeX+dK4eJ9tIZupmA1LIimwKKUCRo9U/lGdFkZt
j2CaR7iOwKtVTU1uSqxGL3NpHJl+HlLxRC31M2plxjJBVkKDcCoB4qX7P87XZHUW
yX8LKb6mZoQxoqUkmFGDXBIsJKcLKKvfVJ96YCjpzygHY8oJkiJKINTZfw9zSZt4
VZIdcDilQFqhQa87nU/6B2LqWY7TjUkQK/ytBR8FCjPYSwNMRcIJ75PFB5E1C1jo
D4P4zyUEL5FDsjY8c7BozA==
`pragma protect end_protected
