// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:50 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
rK3LWLcW/rh6i4A2wf+a+BszvJ1dztZHwbhPq4yHU6OVL6OGFaiatfw8akejg+nx
pa7QdXVKQFKJPJLpQrCFxPJuF0ju6CGmWdo+wMu2TO2MJBYanFQrj+3R9Mp5V076
crsohQS1FUydIjhGXX5juBQf57Dg/sEJY07MCICijF4=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 29040)
l0SZunJlFmaNMicCF3d6N4S9aa5Nd19NOsPyNFCz7pZX8j6tuBtrMoha7rOPjW/6
9pEMd7F+TFVdEEtazZdwwrtA8NzRBQguo9t405ugEgj7+OjRHpV21E7RxatZEenR
jPyhUfEOO7F5ruPKEkQ3aiFLE1XGp29LmnOk84/4dtiLfMgc9EVicoT22KhKiWHr
cnLV0TjzY3h40JY7dsakKeawTOHfjkPlNzrlodA9cQcV+dmbF+rmJaPAXs4onvgx
yoaxjeYgCnpAc/0e1sqNf6jP3Gi7PlfcPpiuZLZBnBTGYvG2aEJt+fLaPkRQJwFw
8rfqe3gG3T491YGSa5SBaquV9er4y9pCFn4rhnj/6wef2Of8dtTP8MhagmQoEXad
UCZy7bRL2nAB2xWazjfLtuWlJZLqVE2tmBxaEWITzV3vnV55G76zR4KAor3nY+g8
EJhEw7rjcKnBtiJpwIcW20hw/3rOqo1lfZYfku2qnqayHCbzuPWcrXgDmdVhSU0x
h25hu0YRzpcDnUsGvK4mLU3MY7lTQMuEwnMUMkLtN0r0uwxuYv3DeNQJ0PDpaXK8
ySLRDjvzDxxpLl3qUagGRy1s1gP+Sc45DEJttqV2V/ekOckjt3/o8BwL/EqddDVG
ctpLsowvxwh6sHmYw/3VNGztDleVWJAX0PmD6eJn1m+1LmRlt3N1k5pCvNbDSFU4
7Z6MdlihCmV3Z2VSpH8yuVIThdWxd8aawoZGhfCS1CqCD6ReiCHDqI2Wl13XhSxI
lWenL7g5Kv2GlbsLUAi/86R99B4AhD57fQZXGYHIDNTfz6pykmNanWwAjax2qcJI
sHn06tDW00dpzVPKYEaXBOi/RpXKR2+nCahBO/E0ZFHqkTeOpFLWKD+0Pxq2xyZF
qTQoUHTton8d6XZH2LS9PSa3OUTt65K+AW2MXsYOS10FkmJdE8UaRTGgCYQhCWEj
vmXrCq2Og0nuBCi9qEOxsRSK42nKQT++busuFCcTWavlMoimfHizn6n3/DmW4xbF
N36H65EV3RoQrOHwyz/VWWvZYAVe50eliIk6s2qdjxM97k42SwHICO+FjIK8IpKD
58tZ1uhEzKHa3iBz1buqIzFuE+U12igOF0pb0XxfK7pZyeDra1os0Ia81JP/j+OH
hEtsajWZa1CGfTOXbMTSmnxTmDbCCRWzXkkZ2om1xanQb/Y9CCnvhehiNGMRpqau
n4Ru8FNYU1kl+YwLUYnwdl19DsLDKXXQyn6E0V81UIT+QbX3CSbfxKrGVHdf53aC
JuAHzSCweYnzmlReJ6g3A8J6stXIZr/3T15QHwT/x6EBxSBz93Rv/yod3i9GaWAs
1jHfIdQJuGEAjv6+rmFhLrP+4tTfTPadCWwXUwhYud+Y7rtEV3/NoaGsyUsajcAJ
DgqlV6BhAD1N33sjVplhYoX/OACAhPUGovPkwJOQy+swf3l6W0Lt4WFEB1GBFNOx
umU+fKycu4ho4cBPw/PZJe9pzMEtXyJ7erp66BwwW11FuJRd6L92XjX5xvZvrSE9
t73yKqSUafbwyZWtCyQmWw9kKXq4lwIau8fMfNe5i8jke/Fgf8+EIqScnbDsTkxz
OBTHiYxITL5qGCDOGesZbch4GVjq3MkvHxlctPihZL8nLYkyR5+KkoW2Hf5XuTDr
LSlTZAGAHvQOR/dL2w+eES2vS7p8q0LXOQDg7Wx9LGi0HDP2jCKriZEPqMn79F+k
uehcUbNRRsKeeDx4TqExvxCZrDTeBWrTpsOoB3XUxqEZZjiQw7EqWqS+7Oy6GdXE
fo/Ge9foF12uVFdBdjBA8Cmwkjqmm0MqV7M7yidyF4q25MdaR5+GtOetEfa4xsiG
2yKtJjTszDY078JuJjergKXO6/fo69UILs2mOnfm4oskN2xwbs+NhbvASQOqvnwB
bOkWlXgtIjGPD/pVxp/m8agu2PuP0JoUPC5Ma2KbVv1axSggWT+zVplByXE+YXKk
losHj8j4ncLRAYVxxZL0mR7gcJQUMIVwfvUMq4MTlc53sfQeiCpw73VLLCZjBPFu
romtiAXRgCSN/Nf8/Onvi7UClH3pUK3p8asDlgvyR8fHDtHzpHw1S1YTNGVG11hS
RrmJoTCQ3myVKQVHtnr5Tn5teebrGKVnkLP1UNjMjhDLEgVGqE8uDam6dVSwB8U3
A5iYqo2EHBije+LgYM020N3eREed8FFcUy8bQXORqIdwI6nXW63XeeLpQp5/6+H5
a9DVxjEvnl3SqUeMQWoZ28AtYFsU1h85dsg8VE5tEquvOpJzTO2aqu2QtTM5EQKk
f43b501/R9b264Udm4iXcrMP4sfIPViIpDOlPUIXdj39LqUZLfnqTGbDWwVGMK8B
u2xdFaBMBNX4Ov61n+MljbPguT8lurJALxQJEfEiPBIN7S6yxacVt2ymQgCYkrM2
J7m+GHPcoZMVWgFLWV7wF8Es4NZY9oCcrcMYpzf7TWC2z7nDkjesiyjnJZRXJBUH
U5svN9Q9NOxBA+pgosYjjEJZKIXIEjx6oDULgXHxrYBrPRA/ySz0QGVLT8nXCAGP
wqgAidxEcMU6kko7hWv/V83rSRGXMqSe87Z/xWVm5BrxsYivq9g2OWozr6WRphJy
FX8ezkx/HYUfDJN/di/oPWucNwnNXZfba9ln+vGuXrR+nhHuBUsE0ITklxZoV31A
cD3MCJrzwWPLcS9Cs/bffaFuTFuGz+L2iabjLzxs73ROjN+I1LKMupt1/fggaO8J
lAzRx16QlYbZqomzng5FG66ABwwpoyrqX2jQLFvu+248cR1tPW6bJ23Xp6+wLTG8
DkyiH6dXGYb+EKEmM+q0qHpnwK/J8oFuDbbJznnPwMQ655I3OaIQQPTCnq8hSCvU
CEuaB953ZkcznKFMIzXaktwENyTXVcN7X/hzuKkydsmt3shmiB/zRmkLT0tsyG45
fY/xap0NIj11WD4a5FKUOjwS0RV1UZJ6xsi6tX4k19mGNp/XHDlPIsocX7A40zNu
YFeU5RK9jaI6jNVnxhLY3w/rlz0sBWCEHejOeFXCroaAmm0t83y6aJ0CdQHngaOj
/QNTiIcWyLd3AVfv4fbmNeiKNDl8327eYcklNJv4OqHm9gMa15cnAIQZGLyEdPJk
AEBBvW8vYqiTgPTbtYR5ia9yVx9RlBgc/jGbvRCmihaoHoTNNarpZtAO6CIL/+vb
dvIjxruD3GJ6XX0vnsG0CvaxiXQhOv8DhWZZwJsNwcA7WNWUFz1IBXXECj3Nzx3v
tDmlkj+ATRsOgxoQG4+W9IOKIcCqrmo9qzt9yVLOgHsErMp4nflrpf2Rsf+/qomt
rRJSfkK4yTGMZ/u/hxGWRGTHTV1MkhrUwdzza0byas1FnisKLeBjOdKwtzQ74A2n
o8TiMsa1nsFOVC9X9VMy2oE3iQnsWFgnF2qx+cpgI4RFGmGsZR7oZrrGLoQV024v
D9jOcxK48Mw4TQMDS7+0Fxw9iFWnoX3VVlWZyCGb70UJI8mqE5DEXfmjLzj8o2dZ
f3Nt4zSWs2eNy1O3qywWSu9zLO08C4FeB4gxtd204o9c431blP0O2mBkMorO16iL
z0YHfpxHsSErsqBdvpaj3JF+7mpy7XR0bmXFnQ81BLfmN5IZslSw/Ib8Um7hyfC5
q1kdrbtl6qmFWRTyo7xO2oXd1M5GRTSagMs0roOPWkclGnhZwKXooohuw0Lxdrws
Bq8PL14MoV9mKfPj8c1X7iyz65mpELK03dRTJUhu5fWBQBQmGP/smt/FRVRbqZzE
isLXV8pSzgtuX/yXdXiYCaWhsRnrxZc1SpMxuRdvPZeIXYi91qQQ/sytu5Hc4ebI
3/0VySgWXEECI8TBUdYsrDkrmWcwSJoHfxwoQJyzv05xuQG7Q9HNAc7ZvAJUx1Fn
xHn5797kLocfmVSvDNOjo+qBQE6EkN6D2MiOefy7p0g0NUczJ4rf3Eav0KD6MYyd
LNQ1IxUhYqQvP35nD4rrv8lEngd/pO7Zmw6+hkLLVQuTsia03OG0og64fK4uhGV4
mTfYVXnJ5ITMa5evq1S1z5elGBZ5e3i+Dqv/wbfVnckKeaIEzRglq1NZczyU+izU
N0vpMcF0/NxwND/DIqUjRxmfS2hGPSZCtWNIXysjbxLOUvaw6hdzGF3cQSok+IiC
K52164aed4Y0BOsWCHiN5NWsBzLYKqJi/YAXYLys2kic3MALgXR0mqnCMXcRcjfk
mZB/1kaZdmL1Idw+AkPWZqgS8MAsTQzUgTsiPFWYKXeNDoGc/bbssvaMMTahQdLu
pJDNJ0Z+oIF8AH/f7ydQ9md5DvT758Ubf2QcnDAdXW7f6voCO1jU2/Om/BaehgBB
HUi1qQv1eF3d03Ownc+UMAEupAj4APy1jbRDVrM0JTXrB3lwibgP5G901tmLWmZG
hFsD03kuidV+hZ8YJWnxF4axXYOjDNbkaM8LKzNxL3Hye6Zdn+JRcroxed1HpT/F
c7GSQM+/HLjFFY/LJoUAYOC/2/oNM7JpwfNe9vz46kEbdoZyYrY9/KoZzecILalO
lDZGlcMW4Vpg9ldJCS/bAFlPJFwI0w//Eva3ymkGrISzkPvzJjaMirfAb++XmXdo
ngSyahWPPJ1GMv800p4oCeMDLnDsp6Cn9XLitidWcdNtT5bVCh/XzJiiQkB+1CRo
LofH+psmnyMQMmmRik6+WW+mSAzuDaG/N67DOoMmU7cyMFha2MIf1YGZGE8OI3/S
bU8NIHvi2XHVgUri4GkbIArq1yynd1Hsk667p14QD09fjb8q5ecbA3KYH4GimPwh
xtiZnlf7yEUxBa5g3ZkM7XyDMMfWwHFKWj3NEJ6GflDL0gFey4xEICNXOuQkVPVl
Wz+KiekNNG3FpKmCqwF9uxk1tZCPf2d2BSrKwosdBO2whhOBPHDtuaZMRL4oC3pm
BpcUPgOMgerDVemSR0snYSViFgM+qCChxMXN5NYOg65jhpKGG1L2OzUbhIhfk7vP
yZRHqSOgn1ZSbVnQ5Fwx6xLw+DHm4SFUA0hZTs629zvtrqZPmcT8BeR+6EPzwA1Y
O0hH+O/35fXM+6XoOvz9w5pqIpawx0m7neFrH9FD+rGOHUjrYkNB+DOzqaZMJYEA
DmGheoxutXmtTG/oB9iNgkarZUEAAy9CzhiOXFSrZWkJp689ySECwjh7uFSq/+Jq
mm4k1rY14PMZ8WanC2GSKXka0vFweY1bHjPiLlIZteLcTY3YA2A9nT9vivowyV52
FeQM1Hcg4O1VcKQ5wh94MWRgFME0IRw0fzn9GIMtA4y0CM2mqq7ggCQumMVBqXYY
+1MgRuf19/yemcA/yffDxQ6xNgwCr1aI1xsXNRI1mOYUKf/Jhjeb3Qcj/q+HMjbN
69RdwhSr882bBZ/KxgKF0FqauNlsRuhBYeI0/ZT/vNss4qg2kcCAkdUPdh5i2fCk
zYJwf73sg2TW0m3KX6oHSOrM0QZId0LycqnQAMCLsLOQpc+MqjU3YyV0YrepMsVU
WY3vQ1j1hm0YlBKCcFLNNPZuZw5VFH3WTjgm9YhLqSFSqt0ZVxtpUJ625Sn8RvnR
2xz+ennVP0vLM8AIOGfnGxJn1aU+hBdse3SBJkM8MIbWyUO+85tBOYz37hI/fz1n
gDG7D0AMGy0klDjFAVsjnXDX9fAAXO/amdgHg6ARsvg8T48x9lVm7NsDn/B+xW0F
L9lfemafZDuu5JFYv2J4gwVGeo1N+VttcR+VIO4XdpQfaY7pZPc420DY4mD+QDVu
zfjtIarEbb9Yez+JeYHDcDz48kQOoDaQXktjQr4+q6VbHGEwGFwu2JJm5AgZyYp1
BleJDD701m0wGpG2ARnk/hcNf7wPV5Bdg/PymNok2W6mUtMNE8fVLxp8jgf7uVau
SFnIK1zAfDCNbSNeZ1g7bFw2A+LQvLGgel7f+DsXwhB1+YY1+Uq0t0DHvTSwH5bP
qFqcC6ao/n5DnpaLFILKTMtcP1fqZloCvycad1T32irPU2Y+smkj/c/PmqoJbis6
4UacagrCb+2kFCndW04cOlM2aUEBWPfXxVBntURO76EvnYhpzSsvwv6WssoYFzIg
v24uvjJNIprvtZYG3Uq1fEaDOTEhJqBSX2aZjvNxHaHlfeiYYZnp3xWFY4TWQu17
H74I5QRAG4U1l389pBcH2/K+vCVcMYI3USxXbWRGt+C1YALc8SAwtPDcE2iox1us
y2AUj/SW1EFRYfCp0iChcZbRZ3tu4hSxwr1IxfXk1MFbSDv/plmuYHfqSIurzu8g
CNO1D22v6Pmog13RmjsbD+4Hu8oCguSUv29qZu99WQ7wOoCzYKm6EOwOf+Oyd/1t
gxmp+g4cZWRQIO/5b2ZYUTJTHXZNYFLJPTiwirglLfxyQ7VZ8QNNm2VfgvOP7VYQ
8dLGuyjR+zE0Kyp3zkdUo3iPcNV8jHZsfMxRG0aDdLdJCd7qlm5S16sPpZ3GRIRb
JYyoXkrMrrGEleI9uHW39E+47TqpJR9pGyAOUxhyakCCdtMnOOM0ZNi9oRcDgAjZ
LUZaObCM4yiIuYK+rtJm+w9IcnFhRuP/dSd3gmeCQFeXuJHnM7xrgGt3gAhedcQt
GWl8lzis6brkTpvqnMPDLgzJ/i4QkRboQKzzp4W61DUcoTBLx2/zCJRxFb7H461f
GNz0Qt6B3u9d2Q9Vi/7U/Hk1oJfWs/KplaInXVl0e/xVCk09KAzhULq6cDPbpBVh
KasQt6t/vkkfpmz2BkMcvAZBdOiB3A9hNbzvKrkgtsDOkXZ3wNVMtGUSUxX1rySG
BwdJgZx5GAHHTqIGlpwgPJ3vPlRKAyyUR3fv0qJzlGrZHFRLkjgNEgh41pctYTKA
EGDYjb4TfG2yOCBOSJ2u7gdGKqF5rRPGUY4hUu4IDey733jXzjIlA2+dzJF+8/7X
6rzGwFZXoj2k85eW2YaBpGF+z5vXCwuQ34oEF+0nCFmN3DMHw9+sfDYKXK0mNlm1
Huvwi+cdMleQ75Bfy+sll0CqXZUyOV5XE5s3f8RfTjHkVnZIjHW6ssB3ozh9GKKw
xBSwU48qUyVCXeMlWTDtEK17QH8CAnytCiuY7bmuwagWi7+2dk85tF0vyvtkmxue
uk+UxFxLU+vKlFnlEOYfYYWfFHBF+tRcZoC7smHFY96Wexr0W5fREfzbADLnL+Te
ZqmT7INAK7hkAJ8g3bTj+fPCZWQL8wwFYAds7UzqunVANk3ie05gNXrp4Ou4sox7
jbuJOj3mf7pTRFdMnQ19llkld4tWPY0oWRjr9hTtGKhsnMqBWyClF9GL4W/rb74G
Ap+xgqb9LhPS1fEq1AahcBJ/mDA1bT3HF39DGV8LJUCfRNrr9DZVojpvnC+nWJ+V
zUziMyqMJmVQi4f3Y78rMu8bwfe+dRkL2+/sde9QkPtlaXnzPInZYFx7gbgPbSaI
+uXCGvhx4E6mt0DgittOeytfPt132ZhxCQ0qQj8BBf0Y7qloM7Dd3+cBZXgocNAW
ekZRDkWZO06QDCPe9pqPWEKE4RUpmtVO4tENUOHSnMfa7QEuu08kwQb8kz+AYzRm
7TYx2+kSEFL8iy7ERyfrX1RYjSrMFBiVJVxj34g1zHo28IlpHOIoRH+DvXd/z/yL
Vhv43jsyBu2dwvvIo50VLycxAbNuafq9ifHFiQfGy/m3arDqaNWb/vvy607O/hW7
otp50X/G8zgMIs9SdllE61OBqKvU5ljnsxq1MqYASx4VUUt98QoQgY/FGeArmRUz
2FFqKM+l01todF61w8VqAWS5F9WIKYlMyGZBkQeztVzCsbjWI/s4/ohPJyPETcMP
zIdLH5Gy2vkAOujniwwVseZ5w5W5PqJYoXG0VTqBfZOiqefh0bWlKOeQ1yybCzxs
4/NPcA9vgPW2T6ouITF6x+ibXGcBfjTiaoujjglJw7Mcpj0iBMMCCobYdA/IDuXY
GkDBCtGfBLNMn62z1KT7FZYX9Zg7T1eGP4Vd5V1AmtToxSc9BfrS7qFXlRszOT/P
EjIB4Lxi9ShadWhX2WJZHqkvgbMIwvV5DWL85qXjcL0h5ulClqCzbgbt/ah4//0e
Qq+WC/++qo09nJ3FfcbAnWb1JJVZG1MdWrmBWmF7s8PpUZpT96ACUf0goYbPCzYa
oxQGPJNbmJi9GNHTd6K6rpI5DiE0RKufkFkKBjT55izm2sQtmBlzU/yfNMp6OCA6
tO4tZOdzdPNBlRYgSCP27SeTtJ8AMI6wdSVB7Y8sZxm/HD3I0ed93LUXzipNjsX0
SSSEYu/9SaBmnwC3ct0UwPo/uYwyz8SjZXT2URli/cBe0MDH4OH1EF57CCPPTysg
FDhKI/j5eU/kLi2s5jirZaYBbWkGoGpuhg6mWUu2UYAU32j3hvb2j3WjI+nhgsGE
OTzata0+hxoI+uiCsmAWmkcj/TDs2T1qChB/byi/OBWV9/UP/v2dD+m+Yrnh6/Ru
Q2azCI4vEISstA2e5D1FKyF2XlcVJ9guiJ+YuoGVSdhyKSf2NEVN7lbBn9f06uF4
EkFX3FdzNLBAdIIg/l1/3VyGHkgFhsuGigbXv9iwAKqe8HTgihdXIytICYe15hOn
/rxPy6AXlp6wN/f6Nap93Sd7/ZMIJcaOCbqpwEONoTwfBew8fTEtHNYDPHTWagCm
rt2vHh39h+RtJ0biZCw5nzdhBAd43G+2vx0+vEhp/QFr9TIg8w6gXoWvpT3S7gUJ
oUxURI+xcW9ZydJjnx9obfGCt0mld7/3CwLmvJYz2QKlyZGKlr/BPl5mWD3laTpS
NHBGGgS7lHGo7c0hvNCPdEtvtSqjcc+hv1iaqG0EEptUTGvCRyPNvOX5uMXVX4HI
Wxd9e4JhmP4oiNJkvosCuNLBDDb5gBOd3YbhWIyoEULX/EyXbasgYBV+bE9prEhE
RMvM/WdFrQDRxpX+Le1ZMN1EeOSw1jiZz69rqQONNKl7dfvBKDp/EjHIKn7G2iZs
WTPmMZ0l3LqYAayEXtBxAOF9ys+PVWBzVD2KE/PUYPeq1IphdMG+p64wMp5wy/38
dECLY0sD2yFgEWciPdfhF8j6xm3hVvyi6OvEAyG8nuA+8Aa6uJxaMt9YLmLVEG9e
sH+qO8W8NHRJfyshxLJZKUVhqM+O46Iz0PvOgu3szlw73KeTJEvrxxksbPipmV1d
M/6COTXMTRD1SlVFt+eZktrOA+aLPb/6j2HMs8UpxeIX51/Qav4be2n7KrYeV4a+
+qQTpA8rhQx7ml6ihvclStvv33oNONWprTe3i6xWqWseOME1Z2ucEJ+NOtKxxADQ
X0Sp5PVya4BvMJ6hD3yuN3LEeo54a3wrJqbRh8a9hgVVECbdldxuPn0RXHTkP8fo
jnQwQ/eCUIEfr3TlGYJfHd2cFK1je8E2fyQic2C4Pfeo03JY7e4igiSNXGPiuHT+
16Ni8VxeLSB/3DAJ+a5H8TMCRws6FtyYRXBi3YPxvIoJVI0zvlD22E6Cw6tNyIQh
bMkNUhXD8DhSax/0Xn6YsGRilbGtDBpuAxJoOPbVnhCppSSULKNKlsofUNKCvucH
vm4tbFZvk5Itdgc1cy45Uf4FO0k5zWX5hrUbYv4pkIvgt6PAX12IcUdIZrLjdxMP
xsXlf3peC7IJv8EvDez/lqSBLZ+THVfzEHGW85HsUo1lXrtOY/G4IP+rEF9zN12Q
YMOtfUWyjuDO6VzSmcczGIxkVYFRAYSSaqluV/2qzuL6LBbaGvgg3LUSlwHn5FSo
I5iFzKqIr7hIW4+5HEmy9lSmSrCBKmwXHRIvp5pPiRSFASHZxcWyjaBigWWKxYxv
xKupUhJ3hTTO0EXG0XYwo19a/nUojnZn7o1hxfqTL7cYShy69F8sh5ZcvRgNMPKj
/EzFyF6WLlGXY4Gdra78uyGE0jnFvQ6Qyc0zTnGzCUoerPmzwrt1ooXKQ3eW1R/g
mEnQ64vBupFEtYsXwirCRFq6yId46SrR1+QAi4yN25fQ2JT45XR93OhTqvVLWkkE
wesNjkpoLljjIEWVlhIasF3xtbiIPyOC7Uc6DrgP7JK5ikHizRN6zyOpMBWn20af
qJzf2/IJ1YGXC19522IGH3uc3qaALkwYeKvSo2yEgzzugPyINLkcz7TmMZWPio+u
KpRY7XQguJ6zj4PEBSuqmRvvpdf2Tu1Kq8CUgr1iemCfQJUro4JH1c0G6gzJ1qjk
NlVUkFkvqtUtPqqs/qKFld6x3RRQa0gDYR5fSIjf19A2uVBZfDPxJJaeM8/xZMEm
llc7+H6l9+Sn1LABedOm+1tvC5EsmKZx6o/9DM1JFV5sXyvJXtf/8IVqAjzErBT0
BLSKQB5t86V7BEA4VO+wMpApoKwOvMEZjBkgUItlp1GmqXqJ31wdPy72NmnH6vyC
p1Vc/sljpU9lWdullMGtR2e6LL+aFreRBQ4/uGk3VhW1QS4P1mbadzdb6DttkJ3n
C2e7o1zvdpxBTJP8lGRCUayZcbaTkls4sNz4yqy/YapmCiveFnuA203rZbbmq/gi
vQxLcfxTLSAPISy0hRi6PlzXiuVGddlMWF3wXdzPSqe5NSgFyLUOdeYcQFrWaBj9
VmWXZio144gbadSdYkw+gfaJDvuA8CQpPk1WTyLqYcoIpZJ4w8Fd+yrM4J2JrVBm
5IAnqLap5kEpy905VnQA6v3Q82I51KekNs8DzCtDyZ9XssxUvmEUxwr4uN/Qo80j
QwrQPhK2afl5gHnqKCLwBBwmKY5iHVrVJ1olXe2/N8G/9MufoqoUict17UvlZ5MO
HufSn4FFLImkyoBxr2sCVLthK/uH57poyc1lhp2cEmDrcMf69u/hsUuCaD17lJUZ
hxW3UYijE4s8mvI7O/H+cvHwmcDpYK7dvFutuvl9QLZtOymrmI6oiZ05IWgWKpYj
65Bie/4Un21+37B+nGV+AEWoVrQcv4JABZDULNFyHq9R77LngTxT1WERdKfYkEH7
mQcZK4wj6W/0uZdK9rPXu6VaI5iChFQGRxEaaBMhGLF3iVnZnwlTTptuovQ03HtA
h+vp0kLEPWwM45neZaAqn731KQrwWQ4jC9u/FYJKLxs9RnKeMFcYaGRwKVZFXGe/
Miz2ZsJXOBxE+i9W6R2PVY102/Be/VYpBbvLjmb17N6eoeeCHyp0Tswq7NQzR9b1
8ZyJ47vNBF1hXUmP60Ch+KqyrbPleJ8sVGzWXx4kmPLhPWeSzb7swcHPTBXOE1va
A0OfmjrW1rn7mN05stJGlZUhgeCvnzrrmUdmJiwyNvtOlL9LW+zNMY/ss7CTwec9
cEqV0cwiUdYfD5Br3pat4Y9M0qm/Jk/RHyJRueYTvLQz8xOqZqIlQ14nQmb1uCzw
uYk4H8O4RiJoaDY4BJk+sj2p2HnU62dF6Na2HNISV4aOzXNyU/JcqPZbmE6dYR3i
TfqSFCJIGrIGOrbTAiC94eoEZ7AwbtOODN200bDru7W7thMeky2PU0BmRbPPNERf
rZdsHRDBRmgNX18LKMy4tHOel84bfG4DYrEX456OwYr6PTJhE0pBglfxqkocVcTW
1Cc9jDVr9VNAJHtTH/bWfDPaVwpH9ZFisN98XuWpnPaj1anXMpUFCAKBgXrxhoEV
Wf2/SxgOkslkEIEJ4dbPB0QzfI94h4YlMIM+a0penMhS47rSQ553Q0hL6z7FIUx3
jJcdahKFVikJqyfOFHIO6e0wXfe5C3O6//VxD/li7s2E/yaAtWyoQlVVYc1OR98T
++jGIQ+U+jVX/KkejP8Y9SKVLJ/vreUjHPgl4CmmgSRdrrhpGD6Jcd0gr+3MQ/GY
z5TgOZObWB865Xb1/w139iiuyTxx0bge2BsQ6t4BI8FgI85le2cWZe2nxCiCgav+
MDLBVIyapYTxxN6iP9lb6vcJZNUyzib2n4NVBjntZ6bdJKZEU7YlKa7HPMgCBBOX
Cjia0TLOrJHgLZFVhTb7h/GocPMZzYEiNa2C/YWnGSkcGyENszLV5eyHRhb9jSCh
sbFxd1OyhM27u/48k90+A7K8maoZeErT+Ko1CfciRgCOK+JNOfWbrsl8kboZjyhY
Ht7/5CCYKbs1jqYBr/UeKQ5hsSZDnyUcPpGcFBThAwRfXuVD+8JmuzwpfnGrzD91
j/OTfJWoaKQ7UYPI5Lslq88G10X4lUBpYfmtBsx2LXWmVzY2NdgSVfvcw8WzFVC8
N1hnF49XWbaYRJPwrYBGyZ+TureYWJN9az/SDlYggpVqVV3Kaovk4jfndNyG+e2Y
qSdKfiutkG1N3fi3F/qNNxrSlamUcxRMgw0OYjCDFHImllsgF/r6JFhIWjoziopL
Rh0rITbMyCry93ZzHi5vf11AF5abAPIPKCp9LuuioCiRjNmWcF2L1fZxNmke/Hgo
8b3iz5tp4W8mKTgAWYZJCfiKicT/3ZCZxhpiibtFzhrGRN21gpqJpqEZbEFOV9up
Zk+YLkMGoXtSLP5DIcAf54D13jdT3IC4VLfe/9GwUb9+vO6/eXGIHceLspOXwkwu
WvYBfCsJC7c7PDC9cat4Y5ExCz2rj3BI8a2rTwqsbYfeYDwgNdTjNiJRqrbMzteA
NWLF1BKkkzBwTo8zvPjiN4tFf5hTyLju3gdxp1/582UHKfwMOZOoD8/xKOEmNyU8
+ojhGJzWTfURdnxQhy6Q7tRri62IQg36eDhYWZfa1yscKBv7OAK7ulIOs7lptzwQ
6xuO3/OBq1R9JbGYrQGq05qoOs5i7B/dWfIVA+KLcgTyEHrEr4bcBfmhHWLaDABX
PQh9a0aN4YcDTigSFCFJGWfmRl4Bep62vXBgZRI0HR111XBZZFcPqHq6WNjYqwxZ
JVY2SOW52Ox3+GROwoShyyCj/mauoa5SMK8XOpjq2AgzPfBhNsl9Vz36t0Ti9JWD
zEt4D4h8q4sj1glh4KAicYqzx57dnA1ulVsfN12g8pNtVF68Q1my5bY9gobp1Wfp
yOSdG0xM60Vx5ra0V8HDYpY+bhtB+01svM/8e8yjSNeDYykFLG3Bp1Xlya4MOM2D
s8+dH6xNHyySnrvaGwzk+Z+KXkBgE/2HiwZjA1aKUNj6VLfP9Y9uT5UFKlxSf5L9
MSCtBBDXAR6myXNn3n68NeTNgFJ0ddfLbxE1D3n7mOkvQfuPjY5yDgaYmG1OkIyC
0u9IjL4Qc1GiglfLvekamMpuoCjeNK/7y0JQMmyF3r8AsoLTjRJs3Y9Qizd3IB/1
NDn/jvKNybIaOZaHatbrUCkVRZbkQVejMi9PfHkLTcLoptMPgRFNRvrawR2iY8JB
myybiS2RIgx0t4WNZVp/l9tfumuXP5GTVu4CmPonHxamTQ2gQ30B3U9GKjfn7q/U
UJhaaJmhcIraLNZv0X2YrK59qqkqxkcCFpnjErLChpr/DYCBb/tPOiLGU10evLBZ
5KCm8Swv/or+cc+onBuYTCSoCqQr6GjPGAgOzczNccTObBV2CBNvH9AgOKxy8Dr7
LZxreAhonvk0Rd3eyO7RtrCfAwTkY4OTPKnMLKMAoke6VMIfnll868k+/02wzms/
gRXlWG+qXikF/In09GvyVt18QLH6volAIYZAAcNnTWelzE7naHTjAIoouCRTUI4B
nLFxJvkXiq+uabQ57Gb0/9LqTEUAfgOS5dk5h/uFKvpST0BqEWAQMxEAxWtWSOBS
c0EWv6mvU7T+2Miv9hCY656TUvMOSz/OF39ipiSCsclkUeeRtG2mvZWNx+VO1TLJ
t3qjAXWZSnlxugLfixuFkF86p5hMlgZaGzy76fbw853nKsul/GI4r8XfKk0ptwGb
lN9cU/8Qh12vs4+oMP0guoTpHrxrhXV5jtQE21hd9P0qwC7+1N+Q/rlhyz7zw81f
J+EK+QgJzWmELhaf4xjJzPMxeG2LvEG6Rd3X4+GX7CheG9kPNcyfwluBwQa7l8Q+
K1Jw6Kgk3umY5Md2tks0STS9WRELqYA1xrIVZ3QLk1kXZrQV+kcdZBxjgQknAGZN
kW41kmO/MxiRdRBLzLzQoOmAkDFvKLP+dAqcU7aFB/+Vmc0tbw7/Gl5Xc312Nx6N
NbJZgnGaDkJhGwiYj0uXsRtucsiEimOup0/2BLVUdJ3dcWx5DDBT2u4oJM1A0Z+e
cfwoeGzd5fN/R6Uv8GSaHHDM/hNQhXxJ2qcPIU2S8ITy100dnkxfRRZ3zqErcBfh
XPLHuOEbme2NYyS9dSgIfELLgGNoWuKmV8ENSB/tf5GzEwUPNbD6nCY+YBxpe05V
ndPRfhHz71kxr58m83/d2LMhPZhDNYXWIfAMfhguEJ9k3dEotn9PGL8m2eyYwYAu
k9BX5mSdePUh6VAnaxsHGL+Kk1Ux5nx39e75VbSliLjtKvPIJW5N6Yf79R35Co4f
bo69fy2tCI0BLvoIwLhfwV/15xvaP447a33mkBvpErtTIwaEqDg85wY19uv/4XPL
Y25LEodQc4t6601mkAzbaFozwEOrL9OM11lTvlHU19cyD4khRk8M62wCGEapRYv6
J0BNuy5S/Jev9ivd7rYCakwFRLFno27FMAdV13PhUl9bn3F2tvP9+RCrLhMDOKbx
Fi0GLJK2yXLBPFu9noB1vH5qwKfXCarx1L3AUBTB6xJ9URMRi/0ez57F9YkUq5w7
lLQq05Xr8KWeE86DcsjxshVh2EkvQClrQpHepRbAjvqOSLYK4XrjxxK6qiqir2Kj
7Z7CTuqh1s8ss7fRcewD2tmUHwH6CHGt9G583LM31qhoCw2FqqxzhWK/NUeTiHPt
4sWxl8Wl97ucCQtppvxSKSw54rOEpJHdjKdYuliwLH+GmEbsqQSnif9yjVkB8P6J
o8DbjTx8hY5pt8dK92I6M5ueqZjgp86q9oLlflXLKBNMQydkBa7ma8ajFhX+M2a3
8T2YvQpubRP8xjAGzBaZCBbko+wyPiKOknDOlJ1nEKub9u/WMoSORsU0OBitJzUG
xe6usiYuW0qHkQsQuLZ9i/H7/ptcgoMcdWycOETecxsPg8yyIt5umiTNu0HctyZI
3YNWJahHDcwpOp7aYdJTwoOQHo7dO9cBhNRlcVmYkCCCda2OlURdAxNyS6tzASYB
jeiwKYP1343C5eXwbQI7XkLInIfXGhntOuNBLit6srab9BxBmTLfo1R6U4IjcKHT
XSk2u+QaFbXrBvK25MRzjvcx7JcxGUunNf5QGIRXeOB6TcSalGabuG8RYLJPwM2G
mMJ87b6riyAhUwIFFFVj2plIxa0qYm1m+Sm/B0pfeq5lX7KpyZFc3zVJSeJFrYVS
eeHYL9PovzoUcIHmzS0kYx/Z4UZzEtIoDa3lchVFEvS4iXVBUFecP4sh+4WCqT1/
z1cxYUKpZvpWM9cxHex9v1LMO/8I6AdfRnCY9E/iszCH20tOnlvDxbqFuFWD4gwb
HS//d6iIVU3fS4sNQP1JJsb0A714FhgAMDbhCv1SxUbNw+mmOzETW7kpDIWFVrwr
3dYqJVH0ivrFvn2yc9/JbqmmxSvwL6XIBINvgu4QJt+O50xR/bJal6TR/FkXAJtH
puEiJM+gwYggPJ2ORMpuRr37OI44+cs2tqj/CgH0kNrnf03UbzWhNxoXbcfuB7R/
jHN4VOw52wzC/qeEKrBkJFO3XFsMrD8V377CDTdGlPVRpbTBJIydkaBWOEA5IDiu
PHItWOchHI9vhsvGidSSJ8a3NQZjj8xcMXHNoAHzg2DfmZnvLj8+oqWbTUNnAk5K
KopYuVW8ULd//amt7YOeDMOPQIYlaznjZfqH8ZmCWYzlRb8B8IZ+pOq15ZXZROuS
XElh0ZXoQanpC6paRov+dQ7RgH4a78alquIDeKL+sSEeuZRvRbTxQgc++uZ5Q5zv
HUW0LZ85JNb3l5zDAYOOlPFfmu4qEFaNia81W+z/5yjesVsxZ/bC3BKRsIWUDOY5
cgLZxphCFVdKrycan37F2E7nrcTki9oCPLzZFaEDOXVVffsRKTp888ewMQ/qXwNB
K1QDbRLGmP/eCnJXa5TZN8DfxosZ4JW8v/pkXUAtCe2pmO6EO15gWFcD0xCLxdrz
2egB+nHFTNnVQ5qvpbS5+9m/9s35R/Qg7UUomLSBGZXMJpnAhdxQqnrTyo9oqs44
r4wkfvBILDEQZmTm1j57d+A6C7RdthqWbXYU4JKf7aDdJV7N3d8TrTyqbAzuY523
AbShtf9Usy+QGFu5HM0j9oHcCmfTVSPuGgKe+0Ta+QMs5B+WT4sO4mF2PntpkW7M
uTFxxCUMsAezj6YrP6z1BFiG4XRIk7sReHDTY+0aeCnnKpUz9nwo0fPdl9C/WHhR
YgddVH2FqtbWTEFDF5QlW3q4Id8sIUTp5CSovt9qvA8/bfu84M63+eYrDrPNC9C2
0FJl1OBksmRicrsVNEqbY8RGLu8em8X8xWvH0vNOfuV36jpuMFXlRWHtEh5wxWJu
Rb+7vl6kGD1Xv1W+TIOtHL6i2NPQosnITWFirArIdkJFwjE17tjytxgjtsJFGlKn
iXtkwsfikg9hyLzt3D6TeFMwr0xVaFyvAGHJGDBc6Ihgvv2tBrLL5y3GDMDdiBPD
emDe/qBCcWW0I1eNqvlDNW7xJUBBq6EMhDG8OaIgKQzUZd+F5lF5fMKJTne4XXu1
kZjJNgRbTwo/W6IXK6w7Xm90Ou1rQR81tFAUy39IzSpF6TI5tSAk1yJEpTreRdPP
lFeTGm4sm9tunAgfLb96pfL+iG0ly3tHa2ZWgZOnOWxw2GiStkLFlL4X0DEB7dDD
+IyHJe6Qpt7ZJk+IQMZ/UW0GZ8JzrIETXzGvDE8Il6ZUwXeY7Woc/VPHINXmtmz0
OlQ7SO1/CMpRAkX3euz/6Vrf8okdacXd9G4pCL8MahZ3FQSy8GzqSh9QP9LvFj4F
cIs3+uGwpwWksBAXjvDr9WRQKb6TfuafB70R7CZvV60ufir3qrGLUD0GXmafYHqu
zrproTVTFYvOMPEqqiWyQ/f8dTrerBjgAgmS+JM/7PfaIuzl+nw9o/5euG+CMr8T
CJpBo3g0ucH8dctk3S1+h4+CuQ/pus/UGYCMrUxXtRd4yhHI77D+qliR61bQeU83
xbFGiwu/PmXyqsVVDJFQE6RIQkni+J/AaNk5qfZH2uPXu066y8L44Qi6cUdAHetk
EqWolOF5stqDuunfcIgwll7QhmW3t9VLemClHBVNNY2Qv1TlEmxGmidb2Bh3D5OZ
iGIixfbA8jh7bSypySjTbq8vlHsyJgROcvSEvXP/KXs30Pq6FQ0KAM5fcclxhF6x
/dnGlwB+bSe/qG64YmVVoi9D4ji0Ig++paAsJccrvSUjjbV70cVPNSo8n9x6r0uO
gtQ9Uvn368QKbkPCvZAwtFCH5TayYdURSBsDPMul/DkPWA78FXcqshsI1A5ZQKMR
DaJAxN+lKdC69RQ3M0HZLgLt0Ujt9EgarzTBghx8+tF+GmIZ0BBwYCcFJVswmhkS
X0FwyxHrXEJ9wSlpvnfXO5k4BV+MB69dpvZAGIBjKQIRXa9zwWv/DTPny+21gI7q
4rRqGQRuG4Rub9ZnIxvPY2xlxPmkb/40Bve8gcYTqotBPlDDagXTNr/eTXyHyB7y
WNxfePpQN7TT01eOwVl07hwsVfWGQUfP0PtVkt1Y3R3fnHF17pt5vDckTloGk83V
YOWNkRuVpnsGQlYH0kRkjt/nvK0DyKuKEBlHRVKLWzvs13dPlxQCoOmlGswZJ/UX
BjxXbJ3hnWQsVFdIj3XZnSmmEXpGumIgsWN7FoRyyiZdF67nm1azY/jbpK8/xDYh
l+TJ7gF8BxxoQaIm20i7Kmz7anzl+AMU7X1GSeTIUeX9Jc6gciERip1SaeNjDTWk
grUgznXx/VgSHG9JBOIQPa9kiQsWCZJjW3oHE3nmwQePzaUCeULscwp8O/GXhEvW
2eczKnkzF0aFKkzoTRsip7w0Y0SXnpW45rzVsJVJ/fu2saH/WlS1lM4ENp6d1O1z
U7HFgrZPXIfSlGjzpIxEJhdPN98IXkj6yi6/wjW4fANkPx/TRtV8jCPDt00F80/f
azFnTUvmMGFFfnsC/YsZilEHbOH/YnRZLQjxsWw+iNynxbI49xTy0DGIRE6bLrIr
Fjl+XKIGJe/A/bGN21a8Qomthb1dnTNgPLllNSQTEUc1rTSiuwM+BbFknair1Qgl
ihE9V7H5WxW+Y0eFw4z7iLw0GKFYAn0Zn9ovLuwl+YnUzZeTciTAATTzI0MdSSz3
fM4ZtYNNtL8ySsorRdpipJ1zyQ+u1VTq7M1XqJZREmA6GgP1vwgzD5Cv/yGyQZcp
jFWTJp2QcoIPE7GCnE7bUzAu+EzKj1PiSnSDPFN3a1j1OFneBAVmbjvB+eE7kFaJ
/1655MHUvk6l4Zj6tD682Hb+yU8mfx+Q+wmOhTXTVhpCjXCd4gkqpqVS/jKCdUNO
eUcBEU011tYB9mUZOffB58XV+w/Ru8zjnuNk08aHyAJmozotV8fdIcR6WLDeMQQR
F+oKIoo4dY3pbcexxF53/miTmAbNZemLm97r1pT/6OOKzcpk4/54mK7MyEl5Qm0o
0TOEbZ3X7VKACYX8bUprF5plCWD22X7TlcsFnAOk8ogM14f9Y8x/1mbhIrGdGPv9
/T8kNTW1N37M6boPeHU6sNgDDYxuqfHx8UXVCDKwX6VvRrkJHDyuPbJE7ZqHd1Gg
E80DjJ8mug3ZXNJ15s6JMRVWz19Q0k9EvpcGmJWT/MWwX4ZdPzw7upUXNDv2OLc+
N25kRl/oVVbuNchdbJb44FzJt46EVKSI13a2IAur7affcfRQTaIDvSZYZ2CXF0YP
BXmZRYyGt28lDbxNGPdoOE0MsZoVK9kWZf0dRU8TBT7pVD1bDXsH9b8p9tjNMdaN
nLnKj35Q0AaxOA3jYp5t4g/Va9oZtzZDxGwFMEjQURFEWZ1mhUTMNvsELsaRZYbN
hfK5S3VjYIYrr0oeUMEgPysODNk7/S9zvtyKPzoi49qefq5O7QNY/muLLDVBQ5Tv
omEILJeuoGV2MEpClyXlgd5i8GE9jN5icoMnu/V93DJ8QAJNTyNyq64w06EISIt8
mRG8a/hODbeMjLFrD4hBEz59zea9/Id7Mcyr8akWnyKhm0eqrv2prf3pzFU+1FFs
F7LYdeb1KcHM8lRRZpygxsnLELD3TRmk3xyGTv8WwVIGVhu0t6fnyo4lMnZIOSYp
ZSA5cVU/moB5TxfALa8Ei6tF0Do+EGO9+HeNIwCXsmt1nvNsA+ZlhuaaTcXhndZc
M6QCzUS/1OMF4rSxsvNbRKXlgvcU2+hRb/B0LsJhcC/B5KR5GGrH4cqf8p1AYPOC
wQnNNIzm2dA6sU0mAWt85Gea5eUek01tMd0kBLaq782uLDxxOVOzjWgpMbOUqc5h
SSrzGCZrU/+jen1fI/AOFi8x51lRw19oiOk5VRUFtSg+jHe1WIGOGHSMIavCgRyk
edrblHaQZVloiuQe/vKHpTwZGQfxHKdfwp0s7PrIqLVzP+w5/Dkcnj7NrJYzH/Ar
ff1h7lFASukS/tXF5zGFH+awA6WirFXPcAXgbg+tDtuw9kSQbNQ8ZQLnmiz5COuH
QulRGy/ELjaMKjdLPO57BkjidwCxAEUezFSPgtNbZGilrQHz6MXVu4NiZYuEjoEb
OQJpyzY2cuJ3GcnN6U+cAPRHA3PqDBQkTaJCd42CAzYVpEz/A1k/afENZP5EskFQ
b3JWp++U7rS1oJIZ+H2Do4jJI14l2JgB7W8Jm1lL4Rae877NadIQnEMVEeu6IGH+
OFmYHVqfzOsYavSVEqe+8PlJ/TptnP8UHz03fdL2PfnWZxsVh8TJiXgWcrLdfsyy
hehut/M3YL38PFmagxq+MHDoC7Tsymdo99UgEJ6RshEMXcASoh9JBDveluzLpCdt
BO/bSeLwzKGT2Zl1tqrfbR07gM243S5E9b7W8csC5ha/EjVjHWCuXmSTSQWUAIxm
3n+njhMnrmFrcZqM3Eb1LgPXCBw3HnUatTxfhBZrwprhGfb4HChHFwAtKeIChd0j
XdPsa1Ki4QQAFAY0Ew0Wx9OEezkQOArZcPwqErTYWExikCj119WpnTAMXOMQSLht
vzP2955WS9rI9tCN3xjnF820eBRRxCOlxnda7AaGz47cIlcyNig4Lrj6C++QfGlt
QSiJ5b6n0skm1wLPDPHQgQJ27jGxaLdpkWkTyNPuqa8DBWNGWsrqVY6bt/M4PDbd
UnAFQnuqIOTl6pSus4Mf16pt5zv8R6fCw7RYs0ttlVMloHw8ebmP3w4k5Pyv+yx9
tVE27fwRiiIJOQPhdyw6gMmMwLsIW7IxfdzSzDlWSjbLTKUYkDwr8IQOHqyuh3D3
vicOB3eaaiV3mxI1l44G+PRhdWvU8BP+BXf75Fve1pY6C1cP1LME4YbZX3s1HKN1
a1kjqbyFhT6u3eiDY52m2MD2gygzKTCkfIvchHQmyi4AID8JB94+BkZVKhp/aey0
XD+iS1u/oho3XeF0JXIZJ8rHZw37p+VwrpyXMoMC5+w8BcfQDlXV1EYsdvV0z7hu
/98hYbpt6AM4ErYnyCGunEuf6dWYzlZOMqZVzARwK7V/Vzbyi8sN/l1/6+OAdz6H
Nr0Dj4Be0mLA4AIXNexTcSjbACIr9XQfsh6VCUQpXIa78COU7z0cWuV6RJteeGte
6nTiwzlUu7XADxK6xi4FwfcoZQsepoF4iGJY462AoyfVUooz6LeqyIDFkxs4rbKZ
c7FGclNhPMuRYB9+eG+NYNJxmXLb/+8UEIcEbOh18ROnBOCOfpt4a/el0yYhNkJz
Bxr/kybIXxbEn0GdCB2zV4wBLtUbX8ML+PlyH08PKxhMzGqUTm0zbDPuem0/5XOE
kF79XuG0P9ekn7NMf2M8vaoTJ2DDm++GAKVtno1HTKg5F9ZYQKB3oEFXbZsfnMxX
4bL0vp4PeuFCH8qA4qQgZNmFIo85OpXhUmdmzAgdKUkWEwfc+G5YSWngR0w6r0mT
rOWyudcY8jaNlGnLAXbrnZuPLFWtk3u8Ja8KV2pa6yc0gxkI8yhczcacLwGZ/IuC
BO/j9XtEK/5dQsXlIYGyi3dPMGKe8OjtguogDj7O8YTUHaMOP+D3IS409gUanSGz
I0etIwhIeBb6xoNP4vEV9nHrFoBYO0WFc4rNnVbd3Zq2D09EAwwiy2cxtOaA7NYu
JHqpBgZz3vOgu+b5LTFQ+U6z3ukHRe923mUYSl2PSW+a4YMeaPBgumtRDgoLyyPn
89pNdQzswC3eF1NEmpHfQSAvB+gwzUmo/RwpH95uc7SO5NaTBDW1r/6mytnS16B0
b+tv0UQGa5C+Blsx0mNdMyvL8tkueQE2PoI+IYFBcNLhP140Y69f+DJg6ODKibbJ
hF+b3fb7ygR+XmjXY0SsHnLBrf726qE7nZfqpFUzXADQRWGh0aTrMlNcAONMVgsH
86+w+8WHZENzikkRwYsfClGyitfpag4ARPNlCVH9P2kxgCyUtSKJxEO0YQM/oQMM
cEN/GlSIhug8Hki4AZdlupW+I7Ui1UBf3Km51JFmbstPRV3l2eZ5/oSS+E4cAGgo
o/VNZRtcFGZSIc+4TN/RB0x7zbWsP9s4ihqjQ0jVHzvR2O3566wU4aLk9FrBzzxB
9X7KIjyZA1RkcRdviy88IHd21vKxMwO+iXTIXbB17+OKpYoAUQTwt+M8leau4adi
vvB9qZ+vcdD49wuK6HLWu1VczRyg0IXLgGYIxUYoEUy4+LH1MqPd7AtORHulQ8JL
n/h90CHO5O1m24Voetf5jVnVnatFFY8TDhwMLJA/rFAqFBMH0ep1/sugcM5uwG/1
2rnI7IKMEkii+2Dy9xx75DwsI4RL+DE7ihLLCpSRagqT3K0Rpf5L9gNZaIoG0VxW
cvLU5fIkBOu7sPvg7ONlqFclBKpFs6GEpVRrqmGBHiMaR5mAb3P28+/qnFbZw2Vb
jurCf5s9HN5CEDL7t9oWJ5TZRjMPXNr9VJNVQoTTFqtFnKj9+JyoakHWX+6ZRi4a
/t480ns4QO3q2y6pfc4sl+iseuQs0Z9ivZARuwSS3zS5G4Y+yV4FJtzO7aagkWX5
891UA6vmunYj5bc9XziCUUCXUVu4h9VrDYN9elZpp34wS+YLDdkOuGfIP9FL7ldk
4L4vqFHJNAb/awkKNWvbbb03ej+QLepNliI83AA/5MhCDMMWfodIjanumkyNKqRV
nbY9nUeQI88LlRomUFBkIDunrms03nbuCuz7dfyE9Y8kT2Y4C4pp5BfYj8vZHs+e
5erztK6112n+grq+VZVatN9kLewD23YdbleIAA9FFbnarl2eA4yB4/WpeWSusT1B
R7+95SwObfpm8LuFdWu54g3zn4KEgJN2oQUZnAvE61lZTPrmYp65fdrCBhIT2LC8
BcrgDCWJXDP4WtNi63QZ+PmRrXWToet2NHCj5ZC+ckK3V5hLK+j3R3P/0BUhqb17
aWQZlpKO5uldVl3mXoenHkWPkXgQWaY1LbhDoEm26kUAiwirXwQgz2iBeDYqmgEO
ZNvf5xAdRygKjFq7C1LsJVEwBWPdn74hS+3azWtXoE5a+Fg89bA6vshsLKsMplyj
QZYtgr0PqaChfIpbP711X0eni066bt0JLbnEH3sNlPZnFv26COL583if4MBm3/O5
HvZ7Q1naYYnN5Gcug3JECkM4RdwBy9CDVZlNKtyvJHG6pWQVAzUscVj85zVKnJCV
nfNPe7SOCiaRJfP0KWvh8G1GfzG/mrJl8nM7wWr+O+/FZbUtPPcT3NYGRKD4+ID+
B+eGxvXP89S9dF7bTuhn9XuQfuxR5Z17nUbtAFgMHZh8OHdLa7oS+Bmk/0Wmm6JO
xqeLarBV96dTLiyaeFdLkKh7WJKGck3m0pDrdwAf9E/MlkBNLd9DiNrT+P3r502I
bZbCZEyT5fTr6WpLsWX2RuxbEKuBaylklKgY+IzzwFFXV/SXNzLaGvDpxZUyk910
RkVogHKwJWM8AZ4l/Ej5a5mmgtpM/TrHeim6xpsw1KM3u+QOSHwxRA+BAr/MTBbY
OXKaEIXEr9MfpS5hfYD7FyeZHiCGznsIFs9BTTXoJaUBU333EuEPDODUhN9L/pat
38+iPdqteczcsPNYhvwMEg5xAlZ/P/TxIBy11QWzjuSMeqs7DpCuZ+6f4OZdOiwB
CARJGnZ2vHWtGE861gr7wzKOgLAm1CG7BmNYZN/w4QeX86ET7RFGDfkI42dmbfyi
iWu8Y4NL6R+DV+UWbpe5AwyqRLihLSMIT/cyxL20QdsMzs2Z/GSIX1XgCHmto5iQ
EwG5hzoCTe0iHMJRw/cItFweYnkIKNcEbQ8xb0zvilArGgL0L2SiRbxnV5GQR8QJ
mv5Ooi7veFBGk8yFs0X5m6M+/aQQr3CDjpcn2Wxh0yAe2CsRPvnYxDjDmj5Rwm0V
IdhKHSl8hPu+r9DINQO0X8w778IsqWRhT1HGFMOgg9ndbw0tZo7pHPOA5HxiGirv
J7zyP7ltmFdneWR0SlqKQgfSg4AZmNSdI392z8B7dOSPbkzrd8eHNRv1nlUqoIUy
7D+VwsW1+jUr5PMWPrOoEbugycgGXJfRh1SlNjcXgVX0pNQl1UqEb2awViv+cJDv
E4jqYBLGmHx++p3mm4svW1uhBgmTLMAam00ySwX2UbIX+DkkkKhRfnitWocB5qXG
CEbJZvnl2FfJTJos/iTudFlwZ+OznyIAksEfD5enf8AuscCQdNOEKWk+Rvj288WO
aFr4Qd9ogWfk68IdSD3cN+y9+l7LaYYf77qti6K0cIzhmKvyUJ6pfsNKca2yZoCM
Iyd+jz2Q9nOQnXmK3fTHW4qMYcevhyQNwNCykHjRughSlsZRyFC5hP7CbsIZUswb
5qoks7/jzAHudoRyb67+PGMhngabF/yX2qBxyPJBShfXcOMh/cOmS5PTwPjzK9S2
ZaAbvL3MqCrjnHVcEcZ/ohSwkZJrNI4S+slsfgPSIlWyLDfqS4B4Ejn3fz8vjZ4J
4bM1kv316DVq/O49Uy5yDmf+IBUtJwrodSWDOlYnqz5dcxP6l5OdvshCqg2te+M3
OCe4VoN8UGrOxFWYzVjtKp/jJkHvLRCmRaSmvZW8NV4tMyJnS/Z8MsJQW1cjxnCK
d2dGiTyt4GlNcFnN3ZaUCkG1uupVFsk6w7p/B7sYYvRGBE6GYRQ3JSMvdQqZ/xnu
/KNj5tiZFquD4l81VcwvFuXpHytVTKRSUR92lVrxN4Gbj+GaWq7nQrdN/3lw0zaL
tRE4vsEEd3BlnpIf/nVioTzJ3tXvSB5A8eN2F7Y0ZIXUBIdDr3Tj1PxuxV1F+Mqx
/H1WeMYAamgK15zwVVxmYQhlit2KnTBLAIi4jYzkmxBcoysvLLVjK4I6BeHRrlmZ
1aFd3Mx/prWgHh1/AuwSsse2drviFjxdz5exHn5HuLVe899z2ARMCYcra5XMQm5E
ZsrPvQp64H0FvhzvlUr+TM3lmZ0gS3ZrA+9TnYvMq/1+/Y/jLO++O5QupM+OU9vg
9LnOiy2iEYzdcoxd5oVQDJgFbF1bIDHwHCCKCRwfAAuedtlPyf8Xwp1DNtaqPCmX
WhmMbQZtyrUb/abEsnO0VgI9wPQKWDxwLbAxznhoMfi8wCnpN5Hw9z9XAHWfzMJx
3r0U9TRY5iAyqJ2Gg2sfK0vwp7pnFgYDI++25fOQe+RzGUX49ipkolQ6f1R08DbM
Uwqv0PQ41OaIrTgsepDS4Nc/B43+xaa/kEEnIKP+gd5R2+uas4ToV7s5yuS4afC3
Iu/dWIw9+jc+v6ptW6YuFkxD5ZT+pKcdjWe2pITSH40gf7EwgW9ccTT4F94VeKFH
RDacfV7K1xkECehv3HjswoZhIS281HstttqLhSJvaFppMoIZbfm4kj8rlBr7b9lf
vIZaxnURk2EqCJBevuz61SmAL9RYOi7wTGc4xZtFwJeYQEUk8ZycJPDVRoVcO4Ce
XKTlrxGgaTrZXgUXXDbYSaVbSpgWpBQgjJ+VtzEtpf4EZjqa5/LANl6dyuGCNAl0
Wbpz9GtVC7fam8nAOulMYAgTqei5yRNLmwBhABeJ3FqEOQXrBSJXUR5thGMLIeWk
E0c5gUXv6driACw/fJG6gYfe8LMpwaLfxTz95hPDBprIhisWnms3YrPcXSTSY8Y4
TpqMlKz8kKRxSibU+eG7pn+qmWZGhaGdJrHZcl2/w7USRa4JRBhLkON+lxaDUOux
MXSyIV/vmlPZcMx5SMpK9YReWLS4ksOT8/y/IcehH9e0JeR814OA4uUPsIphu3Tn
/sddjY76MoOoTjxu2iHk4GzTXDBevU/2CMLa5Chp9+GgQnqZTCF32yTGorkAERVy
sO+z6tYNmC6p8RV1sJRqPrlsB5TrDXe4XRjLN6Yje4OdywHoR67y6E95exf1dotr
o3UxrRx/zbwvp5Y5aKqHUnfuS8pl5I4EHDm5UoE7G4Il03WFBJhdeXgOjzHrglEb
8FfpRf2vq6kXy4+xRWmNYZArDVXNGrj7FbE2RkxAbIKP1uVhru5VBvVL9MQiwf92
Yy8IgIkiw3bRhTuonJzZQEwrAwgsU0g4kP2YZBa591QNvOPBeL/9EX6G/wHb/oVX
CT4eIQxEnAG4jZngF0DIE12OeHdVCySxock9VVjYpnuOV8DREFa1h8l94KjA7QYJ
w+5Zc7wSsY4inN9sDTpncZ9nDbZY8EWdj6plmU8s9BDYfPnaH7xmBUlM4CqXZPl1
RFr0j5SUwewSoe3c9qou9RoU6EMQLl0k/yNr8pxKiV+B8u1yqqGgdw7c/Rz16kw9
8R6NKy975U8YrMpnZ+/f9VcnTP+4tGwoXyJYuWFN55981M5AWdz0odUtir19nPwB
w4Dw3MVjmTyf6St7+sia4E3+3CSEviKLPb0w8V/jD1OZV15jzM075eX9v4VfaLpv
XIgStYNYZBu6SAG4wk/9VQFrQoZOH/h1x2QW6Ayl3zPJyrSctV5d4qHRXrFrzfwd
Bz6FwW/zSToAz9+kHYBqD/7eLgNWA8OtaU3jIfk04wUV/VqlbkJ9YEkQ7yD4mww2
0HbOzB0D9C+I+I9FwLm8hF/pKX17xdjb+oWhtQ6H3d6Z1ujClZOYgGpD6xAvj2Gp
uY/RTasNy4ejYSu8N6OmXHnezoIBWeqSs/mArxMMn8UBY7s8Bfz54n8027e9dz3v
t2LFrO3LHzffYa4/4dWxz/yjEpRbwC7VXqpquOLBhtFLm8vpgjIOq4+u24oo8i4y
j2kyLrwH7bPDX4pz4M+wpA+1aHblbAcYh5JgBXTZSnRg4NriGV4aZivF7HYUQZLM
37qgfuda+auIXDvcgVKe/3HMS1HyDR3BysSqdDEfPtURG8+cxh6cqkeYOh9SQYd8
glMN62Mt5SEDKPVepQY7XPqajoYNdHBm5Abd4EAEiEAwOE4S3/Wpv2JCUwM2Ogty
6gdBYnWu+vwazR8LR7Kr4Db63U/ZbXmwzHEDVqUxjBn1gotDgUsBrC0IR0qu8uk2
VOghuFVwOg0il9HI6UPgkpA+cJuxGVqARprTGd48kzEowrQ/zGvDV93Y1E6iJjDo
BmZAwSQUrGW4GHjywzXZeq2vchkaj2RHm4kt8yMYWg8xGMHnEyPo4NGjRMSGtLgO
V4/Dc/3HoCgz0FLPVHh20EISlF0giT7apVUfyCiNZCpclacL7CI7j8L5fRCGxJeI
blWgcX4ECyLyUI/zpG3wZDAQuxy49hK3mipuVDpOkmAVSHQGxA4lSKYTH4g12ihC
b2TmIubL7qx+c98SjY3OzGzeIAFZITbb/VidgM0JMsRT4UaYIiLBG4G8/TQQuaPr
hxB9+hQFsYhZAdym6vZt3L6KYePBTGwC7HXyY7p0ihKf9fAZqqeCc/PV7zB6A2nR
jCfMYKEInHxIL9XSiw+IkQa+b6y2qLOtNeGsxNr0/MjTvH7ECMEeNZGzire+aWVX
SucUc+HyXftKwpEuHWMFQX8B3J2EXVkGCYRwsE+fSJZP9Ul3wLB4+DNTiH4HSc37
MBreLztYAdGqgqmt5DJoX1MSjhOz8ZJGZ+ntTi5+S8F5D8h1NWigFudOPsWGUUrc
UZPuIwlu0dGIBI+ZNrruiLjlypwjiUoQ5iAlr3TMtJsWonY19kqBMUi3Jl+FlzqM
IDD0t9Vak9HmA6WCYpTP0ywMu178nbWSYAws9aSgmhSBCW7ABoy2A8hIsS1oO4CL
KKj6p20LJdupLGZFNUJDfacMff9KXC7CfLfjnUORY6RJIYupmTEps0sS/oxCJ2+T
yOTqUi3hNmb0+sCoT4UfIL40NjgIuQ9g7NlvogffHxqIn0IGb7eClf5PYhevz4SO
PUb63Zoo/RSQOXFVc+BtKUnoA/B/SU6ORqtvy4I4e2k/LFY8eiEArHv4m/77I1dY
uwLgKwbMkXKaVtChC+pTcHLcNsnpnCsP7SaoHWSbSWECFl2NotQ58ur29nlmf5VK
8Z6V0qpbjf7+5UlcZI3utDgJOtuMSMEg9dplza84VFlwRz9LpK02IyYPo/iGY1wj
TfJ7H0Pz6lghWXl9zGKVSNNvaShY40qWDjk2Ng5ZzJrfURGOIpANOAk3CfBRUDw9
L1MbQ+IE1d8LrmSl/t+rDmdtHUZWj/eS6L1dG4+4WhG9ULAiVNY/W2KV6GuXe243
jWC4+WnfP5dcSeEZWz1sVv1YBBuUkepZvL7MNf/B7NmPU1ggIl6RYgn+kjcsKPZ1
nJ0hcD7D9f1b2ZDHEZ23aYQcZZPVihGC/Ee7jT0iGmL0PlUJhUJ+dmuKRHsqtbbj
q0S7YHcgxfU5NbgPIraePeArKFTc0hWeTSh7xdezHp7eeWBzL3taYRwBhdFU4pBQ
BU19lm5lABXkLkRlf9ymFlN4/8ZhxTP9E8KHc5YDEMGnc8anzsW4wyTGK3P+VrYO
/t3OsbKJX62ExzTOQjObOJS8Z7ZzTO4hslCvOgcm109HMb8eXpmJHyS7W3N3SEJ8
CZDDsCp77obKPQ3Hg9ZFtWthNtAaWZb3zWwOkUyQYGs3OUpi42NB3IBGK0vpUhSL
iN35222DvhSr9W8TRKW5Tn/ejz+sGlp3EzCJx5/K9vb6enZ+oMQeWDSZTH9AiY9u
T4lEEm+y0AxMUKqRrIUjXJ+PgTpH5i2gAmr+fqAfMdckwi1jibyVjrPA14QiJerz
hfsccVNyDfRz4MCak3qlatE1/6y7ZKpkbmqJzHMaw51X1hcS73Y/J/5uPm2qnTIU
hamGjVgiTp2txiu000IhrHyPFscjTghcphUWVnG3rpyieTdAZCEZ0ApK9SK2EWVZ
L3rOk+7bUNADoKyl/xbHbSeA5JNR21jUPl1hqb1OpTP4N5+L/pq5HfkIUkoOwBFT
jvO9QO1VwXJqheCdHPBs9opaNcBQHdp8i5hXdfi3yj0gfl9RmquXnCoA4TadBE9V
WNSU/4yIJZJTxB5aaHrVsd/qHoQJTf3Vm0UBPvbOOvsP2CyOAxuweLCZ9Kwm6gSL
9H3XFqUVRU6VOEjf5qVv00vzDmg1jOHjP+3X//Uw+bzq5Tw3QnhEwRPcqh0K0Dnz
HzMFluji+2lyw6rzAOE9DOKkVdPjpQB0d94VN7uhUp5LezO+Lrrngw3TwLcipuG0
W4WBL7gRKztMNXVjMhDdCp1cDSxK/UVCL2Vs0k1yljxjn6DLDfRw12/3kiVQNzFX
0Jp3f/44FwRSnC9NqIkUCwFzUeGfQPLbnUUYGFtnFGPB8FHygqLZHpaPcMwAn7dg
V3bIpYCHRnOUYNbLIW9MeXKKlZplVFLkeeMiLEN4+v3oeug+EtBi+9243dKFMCaB
eZYSYlf77BaysFa643CYgmugVXowX/dqKhLLbotg/A3a5ZpjcxhM4MHjyh5bFqiF
SNSxoDaEawJSomizM3rock6Lw+nFG6vk6ki4SQc5h2PzNpCxxET7B5S9w5gawFen
9oPTjes2zidS5FQcKhSlFV/PeLeht06u4V6Cd4bKbSjWqq7CUGKMo2IQTzjm8LWf
HbTaq51nDfqf/Z7Msc0Ok7J/WsCw6jw3JQkElmBd9IxByTWx5JuA3Nkg2JXNt0fF
8qDEmLo/svZoFTXjHJwDmeJl4PQdd8e+50idInIJ5PMYXikU1Xo7Ud04cuRMvtbM
CX+RiHSG0ZGwbtXf/DQoFu0XXRi0OZqdVLe9LX1ctBunHpYCL7evP8FWxrsqJ+tt
erHZwrquVhLikXxF//s4dhD8kI7ytMMYPhID5Kjub6qkhNmkgOrve843hlQWxZMZ
+8rLIc09r9PUnxOEWU3fbY2FPsk+paFjVw8GDuEElYG6XtksFlRJfWk6T2sqRn4X
PL4B3zDETlwGlK3IQiMxV9tfdldutrpnKvOa1hl0tzWO4avgk89ZDeuLEb1N+c/b
6IrP/xaDBxmT5f7qs0uMxkcpHcmg6GFORZBX6Rk7VDG+dtYdanDMedbmm4pYFZKx
id098o9tRqyfr3FxTFKvEUcn/3KQdUJ/fd6lN+Sv5Dk5aumpwoOXBC7ggbtLlKR+
IHUaz75FGN7MU/L6uIKG5/uugISrbfsFmR0QHCQsD65kQnwbhXUiPP2Mv77A2vs3
hAghgKWf+A5jv03BlFDqXNj2UJcdgrYBkJtWt574RlyVF3uCMLlbCH8sIoRRXxV2
zCLO2aEy3ad1K1VIk4JsFyrI8SpJQyx+dJ5R719WP2KzP4dpFZFO3gwozS52vfYh
/8eoKnt3QUaY30QmHSsCPQKAdU+2QvqhM5jnYMgLeu6ngTp6F0VSOXPlY/LzgKlw
2U2FUU14RWYxG8Vo2W94/6LkQyRGtxZMPKfWpicKIE0h11hEPEpMdNmbSDCibC8Z
oheDEGVndFy1LVRZ5lxtD8ipyFRG56oA3B4tfLfSa6Z6r4bF9YArN3x2kAIX1WNv
j1hqWY2df3csJ6RNY9V89/P1Wj2BCS9PO/D7JkWSOSZyWVCJJAzSm2hQdaCExOXw
QUzpRv1OrRAwAeBKgRkFnQBZe8eYuu7rxFwl0OY41MI0mjlmp2zDUKfhWLjXEmX1
nIegyhYrk0vw3yMSJussiRVXDFdcdUW+/o4+gTsLaqQHhJmiIQkczpqnQ4YlHRAh
MvUNiRZDwLv156OgTxAe2fODdE+DB6qN6el6SYO4+h+JxFjfKCQ5Ht7UXm7ziAOe
+tnlldjvkvmqZDiXQXZQGw98bEGrR2UymNVDBrPnZnIYx5rjNFNCjnpVja7TJDgu
Wa6yMLZCuouEVzEVK2eedElOtEvcVX/CuEDV8pA0/rwIPZBd0kXm1nyWsyKY+wUD
oh8JNKyzLE+2kwSXoZKxzbJ9HT+n6oTux3hYnVs7h3nNtgaMR2TMZHpARvZ1711A
kX9e/hU3yjGcUmjE/2QwOlobNbGKzUIf1swb498VoRQycgZYHzLNyyO+FD3pNTfo
QGJN9xH885tR711M7x8d8VTIuAbp9Oe9Vcge+xNasFKUzzJrXyf55jn3zH/54WZ7
lETfvAC0zJUP60M87LLrc8HleUPE3GIKjo9RCCftWYgkCvIf+xSi6WBVlS9fkRS1
OzBauhx59g3YnCalW3Y91sP2Rz6UhmjNZBYXvHiLRlFXCm7gEBZVO2mrP8JEQmjE
r6AOsz9PP3UEK9zx5f/jIsB4i0z9QUk3CDBiNdCJtuVBkxNMBwWUnpdkyfyMm0fT
V+pjjqcQsZI4N5bGm4ahxUkhDq3nIuLbmwmtAip+emqlk9BBpJUvFn0ZUxUxzT1t
LOOGJt7/BKaCN+x9c5GaDdf1mNbzg7NAnYR9ntpw/WkoBn41K9xZ41m6fYlteXxZ
VAws5XZ8ijYRCm7Mvc04y0jhXRahoOi3zZn7kjIF/Wbdhy5StCCoDwaRa7m81WDE
EfPsmgjUQV288AQrqE/nK8WYe2S+PDOBcuL00jQ+vCPLFDugQhmy423XTfXUOezB
98Y7NxU1ZpPbqyCZD/inHyzAPmeW4ED2+AQkGsaoMOP624PvTRRNl7uN9xt+pimR
8ZgOLI2ttegxRWPYAcNtPIaiFtzFKYkNNXIatPlHBJ9aAjIidSHPbxicKIBK1yup
AlnbghkeZeWbxHRvQZ6qMpcPG7XFWEaaWruskrEUrGiUO6Q7XRcgUU7ZjZxmqCFT
VKwpzqHp6GbNBx14hAodaKVwPOzJpVsYVVvsGGR5Qqqp7KmLOFdXCLEpvDWLO7Se
TCV/G+nONpnxgIeQiSUVGOXODOmH3fN0BO4ydm5S+pE2YdnZoGaA7327RCh99/Js
zrvyVJEHCXRY01lllUrSoZ+5UgRR82UXOUoofEh2gC5IpnX9q9zh/y1fYXHH329D
DXOVYcz2HYOjufdrbWjIb8mfECtiP8hQ9C5yPmHc1jcp/7Dxch4k9gWr3m4jUIck
dSmuIfMPvuOVWD4JyvZbIvp6z6ATC3aSeiJwWGfSJoY/Y2TudWPVO7rcTQpnwDMT
W5IFHAzYGDOcrKx7cPpqjj1hv43qEGh2Fqw6YeWk33kQTbuMTHqVpRdprXY7UES0
2zE9BkQ3hLRTzg0wKKkb1qJyQ7aUTMr5tl7+G1PhUNKdpFiiBE3kXsZL0/0vVVAA
fyEA3+TpRpHmQ8CeGActFdF9iLK5KelgnQA3vJvdHtpGir3vVzMoLQyswAjh+XDP
yRsJWtGjfzXhQqcXlpK4EgU57WTQPt9L6pLPI23WiFVfQvSYOSk6wB9S5Vc96GgZ
Ibzre2nBsXMZJJf0fL9UbQoqGTNJpYjC3iMVbRSeEMIl4rCzMgJnvAvZx7WZLuKX
nsGqjLojT4N2YKceUdg9iOYxjzxez15+FiFN2d5JE6sCAdrufnt9/Io5aEC3xr8V
2OJEtKC7m21x80C+E6qI/Hfttq2kVSSYygQgsp/Cm6jEZptk7znHnqSpgjq2i/G4
cm/Py9oNOGALzMpcCvunXvn+Lz9DPQGaE7Ipf8UNs5211xZEK5/rJEDdwghoOKBV
NCwKZ438qQxygy2PXlb6aB6pEz+IbtTdSJ3Z9fL8dwMk1rdZxJEpkPrE6WIcq8zB
/xS5R163fH4ZshyhI3kQyFOJojJhgvxN8ERr9wurnoU4Yk8V/nW8eYyPbrTBdnJy
brQ3amLEJLPDj+13jVB96NTuLUmHrrpaWLEpuXiW3rVG5f2KuOVbYJGz5uuvrUvI
DQlAvnIRkXdOsUddF9sZmfoWgrj8OGhalH4CgxEcG16++90xwYr14DFsjg+zD4ig
EWTlAI1egxznCRs4gkJC/cQdUmyRMyETuQMBFwN7476WgQtgtOM54UqgQ7N7uN87
IiXCu7Uy2qDhi6OeWtAvR9W+od97/T83ZUT/H9C+fS04+ft05LPggHcCE7H8wJUU
zuOtDF6l+EHmV9XV+8XkU72S+jQD6zqN4ge13PK47dCAUZ2NC+dGC2JgfUug8B3a
56dsHMy0AWIcEYBwZ2luBHyEuT+hcEESLLhutpBTDEogDyAxG1lOAfjkVOfPolHD
1xVCeq4Fg+ZsQHYNQp/tM8OPZfe1qtfHBBJGFMMyrS0P4G4OOJCv9gWFex+yle4u
5utWe8KSpa9DTSEioi+sRsU4YMMSQtI9gM5LCcM9hWqgaq/6MF1PwFUO2eeOh6lU
fpgpx+hO1yF2FHs0jElkLXGm3ExGx44iaKAsJ9vqrdj0MKJvtcouN8sXBiIHNGSm
tarD691hcLwB85D2eAkIgByk8gqYB92040RuIQGby6iWGCocmp3RTGHHAhJON5hm
pxDL0BS/JA9Yz6jwSJkh3j6k/xh9ICzdZWEQ58DgG17Xa6CLgUDxfvqg5QKxwYYN
CR7PO7yMWSDthfYU4BCQh6wpnocKYxJ8SHKUc3m5ni+4wcWsIob+CXp/oJc7tufr
Yh14fJN5Dtg9FAexifySFbAC2yx8g7MSPwSqQTOVhzMO8qeIPERlFInhhcRn8hs+
qNr8Ii74slmozAPtm7AUud419faWQgf4mdTZUMWlwkki8dVCQ+QIF49aw/nGe43Z
le+Rbt7g39MQBHji+OHBdsSPAN4HGlWQd0X0LsfIU4muHLAGelIQ7q6ZE3QTsHb1
zugwh9cZEsEa07vegn16ZTiGdoc12zN7lsilNOrJ+UPwNfBcYJHx5laPFBrZMF4p
dbvXx8Dzol5n9iCXUH9Bne8hIhLCQDA0U++AIEHfyBWBZpA4XUmXLuIAsvq8XQ8P
CcpM/IniS968rEaALO3PxWHRSJtr3xAfWe9fZbMVbdD4nOHRXF22KNmVrFvFj7o+
J2vCicbVOjat9y3MfmE6VKMpdyWYva04r/VwFfuuLuBi1qBKYkGPivzC30uSOkOv
utg0FCcIc+a0rlFVndY4gp+OsSXakDxaaC0JIaZgAPwuK2Jqn2Ok2ISBHfbiF/gK
M7BAz49A+YAxqdr/tB3ibpC5M2WBS7iWUhM20QXdiOk5Wd85NP1eUr91Kw9KPljl
QQRpkswxjvShxDPHseRUGvvjn2vZqstoMt11L4zQMPHWMCkHjD6TY0TVr9CZkPDo
BNc1S8FDt7G0w5VxG4HWiInpx4Ba1iHuZH1RaGiHVtrQUGpAW4Z/+cEi2J85f3LC
vxE4EB+oorVDWRIeMLN+cifpy84pGQQq9Q9V5XqEJnflntDWxtegH+zLPKbPBzee
AzS8URYZEgx2IRKjQRKheq2PNdygPOUpydkfDuUqgmm8nSre5jzqpjrxsBPoX1FE
+BdzqY9+0h/zOaiQsoxU4RCNQv2d94xRr/7ZClHLjYDyX//V1aEaDUaLAEv5cQ0Z
6hhF+XAmynwBlIgFIhBRjg65y79KdDq7jS/J7eRAd9HDXaudSNIZ9rjahoRuqnay
9C1myot/9Qi0V3vEWs43EHBWZULhifzF2S6oVokCeiiQWgIcPU76+OabjINfVqRH
UbGphxHEOriZ//oABIWGwTm8uobU/pOjdvrCqBY0oqPgWqzJHC8Z7kWoAuYUtkb9
IMa0vj3imgIjf9M0k5NAVzTzOpYYv0gPZoiLeYNl3/5hmIvBZ9/idwraCiQAxcq0
PwytzO85w/icP24RdcNNswr6cn8/Lx7Zh8Exaa/jFunPq0khsIzsSk4c+LKTkJ2G
tzZgE13U9nDDkFNQBpjrLxOMbmRdUqTqq/zcrgLw9X633Z5gVSbdK0nryHnbgqQo
YOazB+zS0diZDFap6cg7mShLODoGlTCCUm7BjRXgYUsXcCmZfVRXRc1RUqpnZ380
RrxMhR+EFKj+1I4vvoame2N9Ddy8jaQ9m6A7ak8p4xKhT7mmc/+ad45vNvltBSMt
Kzb/47Mc72aGt3dFVNRUzruX2bKSuqsA+M7c7tRjmLofIUJwrGJRELEj8dZavXho
cQ08CzQ6+TfBZBbZtKuPWRgrbiKm+quzgmHqFQZc3mduM75QrqetTUkveIuVTMiB
7MXGdVURDnzaya/dDMaxPaBYkgVIGPFoouDm8YKIUU9kjqlThdMhf6lYP0ei0WaY
/YusLH4hi6Bux2mrp9hh1f7eTLQZnwV57g7aLD+aIJofxZGWbxs8ad0fl0rbMeq4
/SKMG9Zvt8nT72/rLaSAB4MP1XGSqIdlTkOvbxpqY8KY7sFsGu6g9v4xyeuf/3kq
I85qaVAUxwW3D1UPNDBJ76qQ+kEo4EIu7gR7MyNIOO1+JiBmpx8nGoso+cm8s7Wx
vU6M+HBhbEDNeBS5VyIm/I8TbRexFVNd/du8X0b2rPNKJSka8uJwDsB/4PhPw97n
qy2sX1H6HJpu+d8e3APj7odcrBekD2GfyxU84ebidmnkdEyIWBvVUjLtnyc85W/e
wShDwGjFKJ68laidEzTSViKF18sKv5f/ex0bzlaTbFs3B4beZOSf2i+vgTHEJMos
U+Ufoz0XamaQhcaxF3WVXW1tsY29GPtDu0IKAzXxhRJH2EduFUM8WfPdi0d09gfr
usEhj77de2r5YbGc7d6LSM0kbBCp97rwzS+QKh7vtq/5ultLxlK9lSh6QZ+bWlGw
7wUi52lYSp43J8nS1qmkwe6P8OseLKjILZaO6KzyQjXemw5QMww/UvaisNoRhSwh
Z0ie9LWe0jmvNezIkoqR5jk6EmDsgguLW4341pc+jm2kazvtnD5NrShDVRYuzLLe
Doz3XHxUVxxg2+t4uN6/4YeDrSM1X0RSrQOFjw13PaNHlVlgAllrMSp3nyXDgd0P
WKWDWowUAuG16ssYtTaXTHvvSMtPk+cMT+rnsXHojr8M9DPjyyJSAlNBuIJA9CaY
A7B/DUTRlWogOBzJXGCBLnEopalITQ33rSl5palv2EWODIz25o+Jcxi+tNp1UNNF
g4AQHKclDM9jqKNMd4cjxnvAqiQqxYZ7djf7g6Vmw7jGoZg0g2bajuctn3uvhOa+
Pdhg7GpMOTUsI+on/wNi5YbUhbjw4HCqdM2OMOehs89biXU7mjMo+0DTWUMZEJVx
ICqC/sRjxyEsKylHTZsENVmdgeVMyTaXr2xhfjnZbJh1cTtGi5DGKEwCuknujPyl
RvtUwKE4gyMpX5KajdBPHkw2TE/ssiDZykkUShDwNiBhTeS6lv7vA/LLD2kAVUla
ThJbFbNvGL6W83RZjsHQeR2TjEVO9F+jGRmIcPR3nver0sno/lq2GpJ1apl7S40X
5Ayz83F7qtdL3Zd1keYxpMEY8pDuO7EKgFkZo3KRA5eFxGK6flAWmeXkYJdq7TOH
jMUt+EMqMEmb7IybJBzNqSmxSrExePP4wPQedRaV3f8Y93BAOtCk9JtW5BeTF9IZ
bIZWc6MVkCHi6J5YhO8L33IHDtBjJr/8cSSkovXuyIFPS5U3qROkvfyVX5M4y/7w
5IEqZByRhb4hsir1BzZnxCUT2AI+sJY3YjwhyktJGrtEjkTPGj8Al7FLfvMlk7DS
2nqb/j1fJ2EZGKEjDwx4kp7JnjPZwINbi+4SqAc3YQo1vSQ77Css7hhJnjXdZqFU
/QhJ7FD90Kp0qOuv2cQ1eN9gfAwZ+EeTAgIqqK5ULmhnNJ4sZkZMKnBdkgbbVJgx
cM3wJJnWw3tCE4Z52cV//aLfL+30JuTk82bEetf439lT09K9LuxTga1YzJ9eopS0
8E/2EeTiseYELMTLcWwCePuAg7YwsyCzISWGTiditdsh9boPF7ReADn1TsM6uzzm
c3GdaCFs8X+4n+OKO3Xit/nQnL0mHTi8LgmTvPWrCxolRpJMs5Hhl+L/aXr7eM/F
wTY/AqRvMntszT7NXvx8ilrzcSc1PM8d3X9FaIHKve0CCnAsHZL7usgWjJS1UVNy
GEDzrYUVig0qREOEIxNmkt0M73kA0XuwM1HTelz+RHMChJkJwCfITtwI0fVwj4IK
k8tzBYs+PwrDZNdp3DMoe4CX+ZvZn6sDyKDLuBiMfRogvMgcvOUbV8lLC9UxhTJE
iuH7Nlglhz0htucSX5GccWw9ZuwrkhNSqqU7K9pNwqb9FL68ptR5na3gWpJLf/Ti
2F9gGJasRl3hf2HrszQtRGe92XUtyEHihtqqUKAPPEjLa/3mm/XTQ4DF+cmHI4mC
9etgHCLGRcJBiAPGB0N853yXhiYpNwM6BmxBFmRzc+alwV6IstwmQRpOr5M3XbO5
81P7VDF0pRQX+zgOa8EsJ+DyWPPOAsN7+yQGo7a1JenwRL2CCFVQkyiHBEoy+8Sk
ZhQk8rxiAVK7ya/XzKKcQuFieHvo9GilAJn3Phsq2Zgu6kFipt6QOgU/a47F5VZB
pXOuQo0QxLFSFa6XMwb9H4CT42sHaizH8MXV89zbkq8+AvR7tCZzeBCLqDoJXTK4
p37RqEzcSkSHIUzpcL0f7S22TDzcEwhQ9mh614yG9s98OfY0AS90kru1GzC1r98Z
/pCP32aFXpxvR2Mi0en3bhV509E/N4XaeJKpZNvBsT8xgKr0TXHtgFWFf0NfE6QA
XMyX1XpxQjGwuSmuwZFGGw0g/1shaKwiZtk130ueoZ/9OxB8vKacjpJjNwNiY0TT
U+6fEQa408OiogWJr7n3BHHfh+vOLqZnCamKaUlYzXrF3yRg26pvMzCM8slOKFaw
KKHPqzx8G32HgeKpwKunLcl2lJqcAexzTK1LNE05KANcXuyAnTmLwyDK5Qo9W+Pl
XQpgEQSt+/f5zaOwRe6HFfIiYvM2nFHGBED93t64rjb3LSEwyzQ3CsEZNiT64Aaz
G3yxSfErOtICPsd3BIrl04zLWgg7qVpGLhchNht8NudqIeFvmi4vLW9edzfSd19v
GVhyjI9B5OhkgepvPbUbQR7SIRjUmsdT88djV77G0SdcIkl5Pgg9R8JoptMRJWfZ
1tdySDUzlYiRa2imih1o1qz+BSieKHcFTLTMSLoy8hqn7INzd7PUqcygK+cUkgS+
WAYlcKRWZIjQC1Tp3XfgeJRxGKwg6vQBYRwVzf9xAOPGpCqMaS2bfamIRFTjt6sV
muZJ+RncZQNAfORPajBZE7Krq07SpbpmW7ruFDuZNl+UfdQuOU0ucxPvIeHLK/ob
Yo0iwq3nDjYqrxqgX+5jAfCJjPsVZjONfDvompHRFoHEMIOh6WU7uJpG3PFpLmas
oIry4Gb4fgo+2ZhohZWTi2oGYZ5Hffc9xZLnKOwKYioBPbNY3dAJj2iY1uZZMYBW
Re3DD22kBLccL1VSYsXaQcI80Nzxh2e7Uyag6LQpjH6gtqL23NJaWW5Iqeab7KZE
iiACI8vogv3Rze6vlP23glJacoxoEMF/cOIM3VOCcpjVs0NjMmFMHixs75GKu4T1
PjWlDYLESSiE1boXmNMUUL98/0l87LC1mE9vQSB3A2q5rDI5F9XkaAujM9Z5IWA9
AeUouqgwPXtuOc+RpD0hapVjjO9eplZF6nIQobJYYeW0S5yDkZE4QThG2JyEPy/f
ixrfD2pN7f2ACNmGi2uVKvFhIhXJdpGcyMYXbw7TVBSIfhIMuy/sHgU4BYyHfq4L
vY9fNJtWdRoGXESHNMNjrkuYxJq7gypHYznxA4zbumGO7ZFGUVEI0VD/pOOzSnfn
kRvcU89PHs3ew5NGHGWBUd6uqKn9Ob+P4dSPptvCtpY9On41FPT/77nHLWCK4Lkw
n6YIetpeRTnE5fa7ICMM4PXYSyV8EXS1zn4kQ8bPDwTBMtP4dT1Qh6SCWFT9T4/8
xySrs3J6+f9e8r8D4Sc4tAkCA/mVBdSk6dP4jjcMischI1mAbErvT7Lwm6129O7M
RcGpbQ/QYNvy9R5vEoS7ucHwSScbtwfvY6lMTpot0P5t+uR5nHmls+11FBEbv5WP
4rbFxjPUNMocrO0Tety99zynsgmW5Ro8L3pPT+I5xUe550NUkvvvTrSpTx0K12wi
eGsSwa1jiIxsi75QF2NaVIqwVCMYxy/mef9xwhiqFqyl+hSj/cVLroeGYWUjVV+w
PRbatziwDeHsTkNUMPURwIR8xAvd+rCUq2zGZW105v2ERhD06ql5PF1TKqMiSEn2
bQ2dZgbR4IIc0GAYM6gVI0lQzBAWbcJBBe52tDl6oxYwiNAqoQKBkI1m6kZrH0ic
t7m4ckRxRL2FGaHiMVWKAwaFspbamGGUQzTY2gxB0aRhZVUvcvB6pDCUionivnz1
5u0Z0I2qPh6Qvp3mxxgbXScC+fd75AcPH71QmUjOd2lNnjCBvwrLeFspFTl0IHLG
QUL+cJEfB8DNONvJQLlb/yUAtyjyT6A+qcriKlc3fzG+Vv34lZwK1brXnJZk+X7U
sVLrceu2d6o5eIlDswjiZI4C1dxjzupiJE0Kow2l1KrE+Sl/zr/5ErZV0lvsGPWk
xheRTmnTTYebDHZHyqgL7Y7JFM2EnJ5qnobWPLigsIntDkBGH54DLLJDanyyty2P
`pragma protect end_protected
