// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:49 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
obTUJQB9MWShuT4VBK0BwSwcOF2njs0PG2NPCx6UsGGc+bUs6KnZF0szNZaaxEMC
rJYIxUY4UnAShlvMrGGipHc55fM1TZVvEkP4gEomrg7plFb/T8fz9aCdKqRM1Hqg
3GBpr13hKgkfRSIo8SLQ8Vfe0KGWF6f3XA2Oi/gwcEo=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 29056)
aMjaR+RphM3digIkeq7slOvN+nDbRlSeeYW94kQ7NvuwTxfNTaLl88+1CiOGBhGU
KwhzRYevbehEJwMir+lnMtw+paPtKGg2nHMe0OY79LkzK/rRmcPHGD8gUUA/O1I5
bKH6vRFcKGzkG2wn8qTpVHdydcnnAm7KwGJrSc5/WlMJwr9ZnWPCkXWNwJZc13We
ty1TxxvMzRMFr4EdG92zKzwelhq1aQrf+gn0ZSF0Clqwe98jG1vjIzmI5msM8lKT
zNNmotiR6Weg8N2vwY3sNk/wnQmNWRI8bp1nDkZoBaRoAFk+CVfY3EnY57xoOqCa
FjC7pamcFwtKL2Y2RxFZhA7pDe028vHQf/R9Rqj21HmTKLvcjFALWHuIoUempgDg
hkFgnL8b3duhPkp39uLtbF+QsN626DVW99+rqKrzTv69rEUaPKKJ4/459IkryLC4
K1oSmWpqRiefLo6RhxIkkZuilTZiIxteTZnRVMKEjgZ6EuOj6j5T5+fUM4ABvaOk
3ye439+lhMRlrB7KeMAA//p1dzGE3gY5WmWfAiF5GDCowZSBdK9+YbH1Wu1ti2h5
w3FFAjHQEBe/cUqFhR2H00kXdtNxOPKsAHmdo8SJ5lWxKcG/Do65B8UWxgDiToQE
mUyGVwhp1mGS9Q1I/EZ9yxbgQ5Qj2ij/B1C7IvVbmmPlgTcWM2IQvOsTSX1PfdW5
QHdE/pw4KPui17TlqU7x6PB8uafNFQ7uFv4QfUlWQOcCDorVA7FQ3MpEbD+lsWJt
KUM3fqVZNhh7r3QsOSD9lqtNxdEKcZwgflRWQcanOivmnH1qYkm/ojqz64Gy3Phz
AYBQBPPUZegj/a2FSdHYlIEll9lUuFylFiHT0Hfw64YBdIGBOPVtBLDix1idHerl
qMugBcb2aHt2IPkOPjiF5Vptzx4DlMfpXZpFZroRi/J5zOioI7/fOyHVa7lLU0hz
xvrbCxSWJhy40hiQRBSQDG2H+sRej4Nrw+es276lR0F0ilDjJvvaBKq8681TIP5s
zW6GE0WaZxNTzdKmpy8z95lncdl8Gd8kMgD/29s/H7141i7hukiD+pyBfHWxs+DB
TSNQtwJBYx/WN6MN+bvCdwNhBPflxNHX8d6hVntWu+byKOqvDQVicw9NmcC0QXch
kDIwICYAfOWulaSl6c27H3J2bdMGSMlKVdH6fxbhEb6GGFfLjwEtoIfkpevAexLg
9Ar4n90GyrOQ0io2BBSkmtJM2K3OVdta3l3oPlDZGjnCTSx0ICUSyaAgmIzqxYH0
WaO5R9g9BYSzlSqaB78qoLlOSvPkQksbBsrnE9pVGFHen66eiceud+yTRA6SqmUZ
9+8G2spKFTVXjxJ6XkhPl8sjSdjSCx+h/E1djNgwf61nmFKmbM1jfT3tPLYRNI65
ih3Q+LE0srxK7V1O90EbSiX3eMsmlxYUcXNMHnHszfEOxUTomDVM4oVOpWJ0lZCv
TaxhZL2LCe0coT7lUAErrrdbsKL34tJVZBePOyrXNmravlMhNA7WKJDuALtEx2Vs
45joy6Tv0KCYyv+dKoILDKq2iAI1rCuSOlKfzgkn7czoSFyimWIgMUofpJnVKgnH
edtRFD5eoRWfUaBUPCZ4rbXv4u5YIrslP3R/7xyrjthE42Co3Cn74Gduh1kQL9NW
r43/jJsPEMYvlYf36nqaRyJEX4fbSdobgIiAacHpfZPJWGzj+5/QUbN5dDlGH7hV
pm9kYUmaFVN8tcnGpsYLslp1CxHEV0DNhWU1PTRCCPHKHQ9xKdhT2IxYH7YExz54
gM65GFYO10zy1yRJRieUv8gaCcHbLx1i5KZG7R17oIxNbokFWmLcyI/9n1c7WHYA
2KHsEmsuiSDhygN5zjz1FqUtzqXHcr4TXEMJHd4x3OWtZNjqljeZTkrEr4jE6avZ
hmnAnykB7cZX8BRxXi5asAnjElMDIlCNs0DTeJ7QNspTFIdXc5sEpmTIt/6nKj+8
rUKLQnRF8KXnAM9ohdMXAQEW3DYeQccwPvHQltJuCWoEADZpnLow0YuBbJgns+Hu
Xno7pAM4ba8TpJ2Ue/bqVGEIqxpS7tyo7oX6WUV14iz2uyjkJfVH84i4ArF4Oo84
2CgIeqpa1MppBbXv6BlC6i10LPdCpq1Vn9lr4bNJtCgLlf0+hUwgh+C3cZp6/LsO
cHcRPgD82mm1uhbcQ7REcjE1PDXJWvpIVNKxrtUPfacD0Uhwh5Zu4PRMUCnNvUGL
fRCC9c4CxRjJ1bYDO1BKXGIgt9I85p8iVsNsZyrBpv4oEztRwUhoZFuCJn3vL61r
EvyEMvJdj99jSGJePxPtKvxCCnyrRcV5vuGLoP1Qny3Qdx14uOY92NWYx1esSX4t
kTQAg8tQQwD1I6RUseLnMxAVESCexj19I441y7VK/U6zYzckyfwSCvvPHE8wZXhc
aanA7EgF8C5yeLRhMJEsJgsqiH7bgc4bZXGQTFNo3cUj55hkjslVOrJzj8OOJEe1
YAYYSafFrPyiivZ506M7Ku6Csu9o9lD2YucjS/Cwcpg5DaNLgn8bUdTq7KjP/Ffe
7P5e7I1vUGMG/xq6shBLd0P6RsNdhi9opqiXYg5racEEXKXJ1Clm3lIjPmdru8i6
bWPyM1+gjcQF3rjFFuU4PaWtd7NZp/geHzg9hQL1lr3YvTr+f+IQhIEvn/E6JvHt
EvyEZ82kYimKutQGWQiAz/TXp5uTCwb9XHhPlF+28rg44m5gBumZnL5S3vL4az7u
sll2cfu5lMGtin3zSnQU2/y0wKGadHFLSB5cY+n+g2D+FgzIgCCSLdaOLBUsSzIA
48OfRVb0rXi4R+Wn6bLtClbTldiIS0755zpSKVvSLTPUXFXOEqg/g6EvWdGJ9f3F
9mNIYCtNlrR34rKr/tKpCD2FebCUoBPOzGgbd6vA9SogYGFiYX1JZqZFBicW0yHZ
hN2v9Rk+LbFMbiWuOisRJgvqk+JMJVpb8LLUlBA8syRnsqwUwx1uZfHlgRxWPUTT
xCUsI4OKzRhUWzUTHR5N1gkATfU/lisuAc3JiuMCG6pTMFUq94oPHm101tCOYcfg
+6ctg65xDqmU5FVWtmIVd4vVfnID1pLpoUL+t28nMdnE86WpMXgjiF77r8YJGLbi
voir81gjHPx7Rl+jpc5pzgBJ4sHsx+p6Zr01jO0BZIW0diVOyg4BZhAaCRsWOPEQ
0PfhxE1XmEoZ9CR0/WK5LVCcR8RGWvTgArqrNv+rDDiYKBpLI1eAzB07Zm/FvEPG
eRHsVAGt9F+fQu4FOZ8S8wpHh90HExVgbiacMw3Iifr594ahT9BPDqjz7y+GqVhS
YEDsAFfzNHPojOlOHcXWBugMfC7dk4Vd1eVBi9zK165/eEJ0oJeY/46mK+7aQGf7
J8Uyl6TVUWM2zj3e6aGQgCCiYpW7PVRYX34QtO495EMc1CNTpIj+ezhbu5qmTH9f
BEobOlH+PzJcIrQINDHDnYUgbk74ae2DVVGiPO9kKdBX8v8JmWDzrFdI8+eMsuz0
n2BV2gKVrbk3V/qVQyN20kDSDToTZLw9CjTcWhkzAf87HwWMWkLUVdbsj8D6+pi0
o+UO1ta/lRV+dBl7ms6RRa0xk97MQK0y+9podOECciKi49ylRqLeW2zHwVbxpiBl
2ILoSTOUyPrljL2QQl7YgyjGn0d5BBE5QaEFMSgEPE+qSanRDchTObLtfPl31W49
rdG8eA5ucdIAeT3dJZeUw5vqNhl/5wD/Hw25nv82FATvPvCDvN8XuOYFQSg/tTE1
PsR6/03USLI5kic+POuJOThFFPRx5biUiVuB9PTiEC036h0qvTVskkjTAhA96BQB
c9CHoh616WV8XIA3aJ/W9b0wzGCrz2Ed4of4gQt5vDsE81SoBJp5vH2f0u53WNs8
spZRyS15hwGEOLQb8U5moKVBwJUiDmauTMBuL3FXqKXt7BY0nAxTmJBOIsxgyin6
otb2z7BygE8+tpo9zs5uAII/P+qdeXakaB2QAqlB+WIh/xDmCfjpy9PhlhSAKn5H
yLzheUYTl/1Cget00H3HlKjKBYd7UtYqXQl3LLawXoZPgcX3AqwPw4QNeMqZyUZh
+B8xgzz9R/aT4UvmJ5BQfmtmQw9qx9siT0jmo0sNNqz9WWHI0HW+KX2HFvHjU48r
7RfcOI+J/2ZIx7zLt4rqG0y4pf/UXV6uQOTsTtRSjmvm15jZUX4VAoL0QN1uMMyG
kgHGb39KXN9R2C7muxOliiVSk0wstdHnIN1Tuh/02bdUHlQkl/yxl8WKgG5xQx8A
OwPlwsPY97sh+lQUfirejVaoiclrjPOsJeBJnic/saNI1hreGk8o7ff5v8hss8fV
5K5nmodDjsWSoWA2eZPLgQZ/HMDbotwiRlGEo2U8/tlpzBhP4uR4TqVVYDZU9EgL
l+X1nQqWPPBg1BRlCC7U5JnnI4tCCEtj7sOQUN7yMscWNplW72Jvyvwb7Hrtp5Xo
es3I4eeHQ0suW4ri4qkYrlPQ4MNwCgw1g2d7qx+eAWKGbWUiPlTARbDkA6CUiKcR
O3XU/fwpKRaN0TfCbsJS1mvtBpQQXPJSW5M+HOxJSxWdSf3ianOByd1YiB2NBdgW
WdyzoOSmtjN9BJsdvCcpw+4Jf1/+GAJN3t9UGANXpjszNv+ObFQ2Wv7abMsA98ab
M6D4B/2ioop6s+qpMV5xqhXur3h7g0JSH5jg73F0uStpZ1tEq1h62kbGVjy5AmtS
IjzXB8SFTZKeb/iRIoTXgsU0X5YkNF7HBl2/Q11QwpX/zNHE/i4Jyd3UKYfDuiEv
ejzrw8pZGAc67xw4RRxgFNslGwIFeFPSE0iaqCrIHR78qyuLqvXO7KpjHr+zsntA
424GP0ekf9yL3NdC8pdHabZJd3pyXpQIf3zbLXDX/k/HX6T43sxIBsdfmfolz8cp
MZIk4fKjP1EoFNhvOGdZIH8zbZ0p99UnGYqCQUmlYvXu/+X+9IXj0mkFYC/Uvh2j
AgkDPe3cXnTZnwnDLpFe5KaQViuv5r8n18QmNkvyVKPMZKtQutKG/VBAh6+QzG2n
yO9KFSZSFqCyel7f5FwMHEJ3Gx2PqZ5OXSuREc3Iz5WOYQaK3gM2yD7BnE7rV99N
JGFO6dIcCApmLKgR+ieUxK6gU6VqLaOiQCDCQ0fWr5nZHi+3sSZEiVr7nArhzMsI
Fz77exhqCw6RQnqOm720kw3MK8oDlfMt2RPYoOqcT6Fa1s3zqd4G7RykqF5V+k5y
94mGxOBs2rPe5fknOnaJ1ATQTcnwbhVQ4830Ya3P+Z9jHTthD8VIfDEB8vZSkBS3
6D5D3QK1wO9F1ckwnsWd1saTbEY0uxJ2CbGCz1Xm5eiXbPwm2eHc5mOf7/i8bvWO
LbizC8RJuv08SzlBvbl+jYC+x2DtP/RPHf7IfpGWmAqGXGPwJ3amj7iMqMYtsN99
+FeAUt43jzwdJsTC6oUYDyVHg4/B26kNcOIozTQiFCLBcw0I5eNIr4Jhwt6cEgwV
yhhj2xoHDnkrOJRXuiOuSRnM2Jj4IjFzj62r5glBR70NtnHIsPlYHXAfpwWRBJgt
A93amqhVpP0IGeiStZ+zoTeJkswVtGk13psL3klSPFjhwa8GvPkm7CTDnJejQBSI
lND99T2ZcJrz7/3kWUWM1ioetjX0Dqgu3DHlNgaIzk+UPEdwOSzyJp+Oy/DlxjW+
HFOYPXJEzYEFOXwmNUfIS+VAy/eR+GmUdiS+KYttA1VWd/ug/4BDSKI8W3glqJis
GEZ0Ygh8YA1GPLhKfkId5jr6V1prdkX0pwspeL5/Ow3GPhF5Cq8v37SJvxysUyK/
pOTLJiqqm6yU3TeD/c2J2xomLapd6LF4j/0nAVfGmkBVnrfmGBUxaXOwNPu7KkA5
cBLVzum/q2m/7FmsTqzoQ7nV1CIAAso0azi90AunfomLH9SGS0Tck7wk60BXkJ9v
rnqctGHgbSJV0KKgHZAbZY4rygFeXUEHBzJm810QoOq0QDGVp4lIVwqaTRdo21CE
w6SxP0qEIzpN14F8/J+k4leVr4dZLFQOt5k55m9KFOTcW+4SUbkQbUEtLgHHEJsK
zp2rkxH9UU1YzUZR0zSrIcqzfERMS0DQv0m5sQ1zDG/4+KdUgClt29sBuyJM5Wsx
47FDQdeigCFBnoJCq6fDljG5cO1JI0Z6aS3/meqOoemYaPBjsSXJ13IguaHD9Our
2kX1DO+bXb3J2e0IHBiu3VuDbBISXBwA7rmaiHFYmnNA4nE2YoghrgygN96MFGDT
YzWtr4QVXnxN3GqPMkTQ2WEe5n5FsqLK52mWkKG2WunB+2iRrM/zktPPCY0Mpje1
rQ19XXhmPTzert5i60AkHLdwZOTshWi//Pt7KphUmIDnKLX4Q/l2uBNNqzFkWgbg
pAgSx9b11ADsd9SQln5fNkeM+KPfb/1iGLVHCG99tBAFcopeTwb8K1ZigsDXLoIP
l42/th2P5FW+kRvlRHdac41BB01qbGaf/jE1bnWan0UdF8YffQI4PcHT9ESC2Rhu
sUzg3G3b2L00EMTJPkqdHkBLdnAr4+dO4FhhySSddtNKj4I7F0DtXRAfbyQvD3Am
ElldCAacuWNWk8j2I4NnJEoy5iHNiPX2TJq+8vCfGov7rvdjc/QAr1MQbbztqS17
A4Ybbp9ubDy5gFUA2bH6X+VACa7h72vrtPyeJCpKxeoly2HUbdfFax2ILW3F5vme
eNqDYkNnccH/BnQCfwy/S3n9j9cGCmCZXKK1H5+QaWagVkCHI3IWyI6iOM0k9Mcf
Vc6lfrbOs1EhSdJtRlFzWFUFWQQzvGdPIHkSDoBk5capGUsOYxubBfwahl0aD4zn
dz9lcI/nTpXc/CLfy9PG9gfC9DnnaDQRkH2L/fU4BNOm+59wyhlU09w6glleerhv
8+e7q6ij2chuwvFGdUnWJkmu4q6F+DW10ScNTn2mG5WP0s4dLl+tk2KRmfWgxHKi
oEcjIh7O8CVXuIKsXX3Tf0jZPCqTs95A+6es/thUhqEsEzHi4N9i8VQaouILA6a0
FrZBJvfAmwggzmN75BGqUtLhGe+5hVaJzl66U0yRbEf8u4dVDfb5xsQ+8li+owcU
qhA7iuNDG9YF1Yah4qSBOLouJUJlIZGRcrthaQDyxeGfMuL68xUKaJHuA6nzRts5
a5LJcSF1clEIkhQKwNHgZSKYe0Rztj6YcBUNSQ5RC3Fejh60g6hY8MLSLoIXUwG0
Mt+gvIH129oe8mfdV30nKiaOewztzlHvrJGx7CnQNqZqLF4g/pR1Pwk0iRTNmr5V
dtMpTWLBp8tZ6H4zg68QREL+oKyfCKjQktGQNrDC06NlLC5wkIX4pHZeCih5RjAF
cijjs9E1NheEDrjFXEQqgL/1l8BOZV7H9D6gWbUu1DRrgXuuLQHrgZ9YEAmqH45I
wGt5rTOIq34+Zq39blVNFiOoSy+1FTkd5xRNpWTPoe3akKPc4jGkE8WNWBPcZist
rWVT1RsvN7p4TbefHJf48whBLVVzHMaGbMEtcIXKgTZZItmuOJj410a8h9rEOBfs
5mxdEi5xIObMvYCaYDimnpKGlTy1JUosJR9uVD2p2FEy8wcc/cT5K7zjI2AEikK6
TT/UeWFrTDrrk/FOhDInXcol7hHtW0w30tvTGaSnTzOfnL4OmBAw+mySDLOD9yaZ
wcSiJbINDKRv16hVv7KM/xL0X9nf/6pZ7LwXqa9G16Vx50urtxlQFe6nOwP72uC6
khs849QXuZb1luiO91arY0vTF87t/vW6/8jHF38o++wKKZLOPGs5iFTZOp3OUJG+
O09OuHgIJSSZ4cASyWSRVLLdxgfsT4Y8mfuJcB9K4IeXH88mq9unt6pvb10vhgfd
E5wYv9FhdNMblCprZU8z521svqFjsMSXcvYIm+cqK6bvBCq9/Lktev33dkPUMjyA
c96fhm+IxdhCPRdwnuU4aEHVHKniiWibmjsqdhaePXhsJEIQGqmVgLfL4q1TYJbm
a254yRc8gxY4Q0i4FoNz0c8K7LLhFreA9IzJ+RRn5P3wdHc2gjbxTsxCcCDAP+O3
/26ggbAd9blx6XdEA//AbWGgPO6DY5iMd47pLkkx7m1d6634LVOpmPWppGzmr7b/
IjOg1/QPPjSD7aTskfALF+oS8W94ydXVkoGmhd9/R67457rknwn79JrwM2RazIHR
GMrTNVEtu+mwfS5FNqkAHt/noXXUyHcfUp5BpJ5ArmitP8tf2hvjyTFdQQZAxkBP
rLpd2ywP9GyUb6yQjWyIMJx6dBX3LEiRS9I0BlUtDoBRktOCC4AizbStuhl/Gx0M
DeEF8HNEiz96An0j6LJ/uh7iWPwxI8y5TJUeR8V1zx1reZJ/yCRinsBHAfa/vk1G
5jXz+PJXdRRvcleoPgKB1TiVNyYik/js6zCoa/ubVk5+HMrJvIlOfScI0cxxGDPO
64anMBSfD5In4X0h/mExkQfnL3WsX6elppZX/pjOlcC5WraRobHFhpA01uMTuxVV
ucVJ1ad4zwH6O+UBalMFQoIIn3pJuVIpJkkdCaRiQpjlsRLlkvY/LKTQ3UlZ67LA
rWITVkXJqUaM3x2LZ2M5YIBO/6EAHvTiEgSMBpKO2BxnLc7FfkQYEW+LetanxNJB
bszUIlPzjGH/Lz+0F/6Fm7cUB+l0d3el1i/n8j9eiY49ilXsf6YMIR3v3IONjIht
wYjY6lYCmKFLQrZPHyzoMTAGGSrZUT5FLH99yaKXQMV51nefDqpfh8WWnhJaM7Gd
WueTE41HLGTG0813faI9WcljyDnxk2I3rnD0y6ysy+Db+XZdgRNQxUC+3DDNaOE0
b6VJdEKYHDYABkhqdUbIwpcNtsOOgRcB79yINYAbctD9/LrdY8alveDyPjM5N/Gu
sQtlLFXq/ITTjIF8xAjh7ELg7mb7p6Xcekpe+cf/U0Hria+RY6v3/4I2OVCy3bZl
k8A/tw4Vhgpk01exhHLbfeUmGfZLCixWw+98psmvzBXrFJjY/yzPJpjzTmoEzvXY
C2OPAqISKy1WZjiphHoMBvTg9cQmuDIRivtLUXVlBUqca6zmmg/WNGZbDNjnjQPF
Bq3vB/f2NOYKaAuzoEoomprs2IpO9ddmeOoE9C79EETb6KC6HlfM0TYyDNRntJ93
IwwxJKBORWx2nyR3/90CaimpjVrBOc6fc1S/zhK2w1nikVf5yA9/M/IdteaHs2sc
bqidzL0igwll3GVV1KXRItPhWcFI1vtC2Rv3mUyla/g7weZmCfirGfDpoRlbvDWb
b/6b8rf1a/+7XAfsQT6sOzVsvFGeNQ/EbnAA+ib/6a2UKdAbGqzgUN9tY9nEigDq
yHv3jFIdUckxzB8aIfArTpgo0IiYbqQTGsa/b6xM62C9u9+f2qWm6Te7A7WpHxuj
xuEzSJerJUxVsHWdde577KXFYHx3ggvY9RSSGbWZRlyDGFLrMMbEONf3pr5YvcQa
mL8sK2hsqS0f5Z8q5odn21xoRP1dSRc9Goaof8fyiC+hWTmli2in2lJqwlpmGSVi
BSr6twSfS1DhugFf6ygc7GIBzqiHLWE4mQT8lYcgSirgHc5/xMjgf8VDH+oElg2y
87lGnvzxk5+2+nCRJ5BcdmcYrWVZWH+vK4DusW4vx2gjv1tz9tR6+38oSJGI8/tX
NRuB+8zDLsIhJnHtAW7BoMhupta/a/GoENlOrkcLba08EfT76lNunJBKnQuMKOTs
Lfh5MKBhuF2N0b0Aa75PPNKnfRUhDJnkD1PKohYm46M9qZt80hc6MMrcq976FYE3
PTg1uxo7Hj0jSqiQnchFHz168qfd7W5JynlzNDkzN54YB8pnzisDWVyOGiDJgaJ9
AmtBLxwY72q/hsyOUFFxTS3hssO4dIOGI/ccNg8Z+cH6vAPqhDBoEYmFrTGRfwMW
XsJWx0PAlBD2YUMBvDk9udhsA0MBXBqT8/+zrABMUtMg+PkerjyTkRPP+zurY7gV
swsOvvWKWPhSmnBsPVKYHUgE3poh8/4SlcVXvVGYZpJlKdsTdhQH4rajBv5qtdgR
roWUNgHcRLd0MXUUiZXGqKFkYcHdOUzWtDEHgiQikVpLSQ5y5BuFWfx1d3dS326x
aKjXTRIF5Ml4ua0E0Z2pxFaTRrpXBQ4E2WyPNPSs3+Kw4X9O5lnwxMYmtLoL3T0o
/S1nRoeH8X0wongpU/jsuanfavgDyUEd379eUdzS2jveOwSOUcRHdqsknFf8BSjm
SLzWw8BSj0qZ8kqb5DIH7agckjrlRvTJnpSe8FEyvUPIxZEM8cti7hF2rdVRbzAi
whMsiOjf9TJJ8VigolLUiBXP1M8+CWXgQc2z2bweEvaw7/n1Jh/Ha7gh/8HZAJgX
AD3W3U/dmc3btxcp7aT0W27W6lGMIysnxevaYgmULFn/xVaqkZ4k6yBGeeQRizLn
4K21LlmF2xZcAyY/2mrUfNnt+rgP2R40k4qlShI+tUFWljlCdLtWukhEYRU+Rh8m
g56w/mICO3qTs3zBZyOyNwg+sNOYzks9yvbX4ndmawgqSt5jsEOTMFm7fBQeEwJM
jkAE2gO7a6ywdTAUBqJMugDJDpH1qnl1ykdcevHRJZMdLfRy9XEZ0dmSdCRsP6O3
ypEyTHH4ZV/iVb7zp1OVyFU1XKHxLR2Pefl9GSq/EwKyhhfZvvVM0TlN7sSNX6eT
dsXmPkxjGQurko0pyBrdYRnYFYKjFm+OFTXNFeR2OOSHYszzkiEaWf2Sn/xgBU6o
EWxJgJu6mViZVoJTBq5C06KOEfiLpJpz/XUdsSNHYvf7o/Nr4cXM9ZO9ca9WN0G5
TnjHBmoxRNjjXLkLyk6iiT6bZUfhxUvzTkJ3ttfnXjjItmQmE06C33YYR4YpZIjG
z4V5CeTOPy5UncdCxNnvr4JTwISotMjYktxH7T7mrsW9l+CloPg4qQb3YWPUBQ5H
wfQTt4HZwOlElOP98sThY+MVN6iNn/cBVifC2x7wbJ6b4hPLE+7BQxCoASTJ9utu
fqpq1Lu7Hhngp4kJgNtMj8SaO0Fv6sHYvka8urXoC6CMpRjF1+zTFbKhZvhybOsx
bl7iZUG3ubm9VeM1seL4DUDfIjgOwzbzDI2RlCrTQVMqo0BtYcGK3tw6XpMV7/8q
UF5AJwnFQEvj3o94yRKWKcV58CV31ppEBXYDZoDiqjojvoWCaFnopWbRKNxwk8yD
yN2QbG0rkHjvnzhCYP1CNH/jhNhurbuQzh7cAa7NCyaIcAPPOOs5ApYDwXtqrXFV
19/T4NM9/lGXJqDb+YP/gkCF4SJv5iLWuJDEPvcKzwfUHuTG4RUh3NTLRK97o+8f
dL4Cb0RiIRelL9PEIbVHqVcXPGn29FvMAU7E/hHtUpqHuuuM6Z09jZviCWbXZuxM
c/+6t7pC7X3Q/g3dPnajKD9hX98vH5cRlCekBh1fK6rgLRMRTXBP17S7616muyKO
XDFwjOVXj+01HCr5OwM5PkCBkeb0R+yIDC0bJvJ3AlgbBQkXEDkIgJ3XdSJw/I5Y
qis5G0OltnBg0qtSJ+dNB2+Ys4nEvYEtt4HnYNfDCUjDeO/SueqCD99er3YS03XX
iCB+kobvBLagWjENl6Wu4MWqWV7Bv4aEroaGHa9aBrLobcFMieIRQtuLNMGWNpXd
LVOVLlsmM/Q+IG3aRfnjvQOowubx1mb6xksiTFOnHSoK2iNRJM7g7sBI1ivI+WLf
TUYvzBmHL13Fv4sVj7BpCWmU3JbgOe56QTYCfPUvqZYnw7n43NG71i0lR4YxxR/O
nYCxFhgrL5rdOMr4VrYy39G18SZqS15pr6V3RNvNUP0RecAlgAtZiDFIAlXXz3X/
wWQJYeWFkzOuRGiI97eQ9C9RsCNE8ansXNh/h9cyQPW51jx5G70ZFCGKVlEjFi0O
eXGFebL98hS1vmeEWAIvJ676XYIe4Oc1LeNvec9XWgQ4dQRHtEEx62KZHwsI2bDR
qYspDX6bRibCLfNFowZmfKVYodyaxh7bfCd9s9Mvgc/woLLHeLdf4SuYzo5jgghW
cYOaa+TAMytjo4y8go6Vzd+LZzXzcuH+7aNPbYEm6ec/oh5ay8sC/Ysmq31hJ270
EAuLu3En0UOU79Dx9EMxb0bb+lsx39Ygzqwecb+/yaXsXdBTjFTs3zcB7NXNlNDJ
qSu5vcvfTcaNJrFx1AEFr/XHodwenbLbAT7g+u22wBoG2cV6GF6ZKoUfmCLrXVTQ
Lgu8ShSce8YBpuiAE56Z8WvAk6HnQnZosViZ7uZLHztfzsUnNX2eidy134r70P/E
pol8Iyi7t6A3t2gNLrRRZd8SnfieZCbfk7CwecQFZffI8gLzw+O9cJ/f+unAHgHG
wsEyaQVClxbSKqtBwj2E2FYWau2c8nroX6aRQ72E5CSgbOJZJO40/UQDn/YA09Po
+aCRPxkNrsSXxIFp05AnQejs13WZCMEux2kmNFCPV4t+EnWbkDqGiMJsY0YQo6Vz
p+xzdXzyoxEBf+mO2e5ccwje06RaOBn8F8KzEanAdf1V2V0eKCUKDoM8lfsQzRY/
XxL+1+xVRz4d+cThr9jkUlu1hL3P50FM7BzXodEjEXlHmrCutedUc4mLq60S29eb
BSFnb0a8v1LTzht5Efv0nGXAkOlUoisBQpndGgtO6KVT3WHrCNuDkrL6k87wp55Q
TK4CaorGG/2NBnMBJ3sm2dWNxaTCAS05/guUUIi1vtcZIhprjwe9jlpRObh50v9K
nIbFYRLt4nlmPyWbKCJ5qhsbDFaN/CZi1HrKpdxvpFKbuUvYxjwIobd/BPty2XwX
+DQtWOkwcwPcMv3hcYx0Yi36m4DRw05l388GPWwNEDYq3V8FJkp9JSAELogfM61k
A1iG3a5ZOS2iLvzFe7cNZLLGlvMOpUrnyHvE0RQKKOHzIoUbNviyPOfXGgB9zZt7
1ycq3SI30WzwJ/J2POkhP3MurAswpA5hxOXXvR3BWmZ5xNx+7QCQPedzW9ArI3z/
h+CWvDK1hXCjvEYULv0EBU8gnMUnKI6uTpiHm/CALt0XUMtvUkTzppAj2WXfpEWB
pL/4z76abkTNQN/+VjGsYv06750DBUXHMqmhWUJt8XDGb121xpFsbX5Cwthh+2DT
OCmUFb+XZkP7A0fMmiAOE0wsTqR7GwP7OKDWOEUGdeZfIDmdF35l5ETuxpIvcIN9
NNLd6mafbxxhSlfrtqfQu7OMItb81EIYX/6UYDasvkQzsoMRUYHoBcG2Q17GJdsw
OpQEd//uBKaNmB3jV53UjkOGgp+PbBOZP/xrlWMmfKJUhpyd+fe9wtnHXqMLSfU4
5AZcM0dBYK3MlSL/vI5e4lQGXinVvw6mUwtkKAArjo0N8LRMJbOuIk6DcaK+tIni
l+7hjtR4rHjI0xVJQ2+63wDGufF7DwittLRWqBxnm0n9WUfnhy6BixogF+CScZnS
wlSW3nUI4j/gPI1wg0ekgIMNiLYQAdnewbEoy3sVHl/G7YPZzNo39atcPz2bSUxV
9ONadfDIU7R8qENIjn6ptH1IGLlJaCIPv/tZoGggh5jvJLAzGuBB6dh4ZuvSyX3v
9zYGUpASGp+osPwPwXWe9g/kNQ5RuMC5KxaDz8DBgMjR5WjS2lrM/t1+zMcxL6y8
A/x9Vef0B26TV8WCrnXHRBQqP2sAVppDS2wBrhTbKmmkzcw2m4lpNls6Vh8s2yKS
Fx4lJXHo8e0Af/EJi4En+DHh3EKSuX20pf6Qlm5Vx4g+zqEejjrKIxxVdk1c0r/r
wsifGN4aXBmrdZc/zLSysPC5WowpWrt+jS6QTX1nz2pD4KblapFRftqBkCwlsiU4
96CO8uT6C1GqcTGj9W1/d9u8+KA33lnIt2NOj7dOprGgiDlTan+y1ZIEDzWOPEzG
0x/HIMT7pPLAViD9Y75zkDeXKerm8J5IEZbeD2vIxcqxYFmZ6YBjBlEPo5i9CZCY
HseRGBGNpK3WRR+AHEi+3nfAIobyH13xC7bTJWCEvdTEJ84LKhWy4QXaywWSjBM7
f2T6oo1nRR1IjOknqDU/KjrVgqTnQiOvUOvIgV6jPvPgzeMwKvkiKSESd9upT27S
KFA9lno3qfNIDezCnC6XCgAd8W66JaL33UYsvJs8CKOUhV0UWk2zbWUbyLAf0yj2
KNbQR7UVmjutq/TAomsOnIvXikve7J7q76v2PvMY5gSSROpeFjFWvApgGKZlRwkz
LEPr1rtjMf/U2wRQmOm4Ib2mbQkrEwaBY8M058vrmOT2yJR7iy9/RAVHiPkvfGmG
/WbM2LAlLNC98h24jI/oh1QBdvSmPojqgq3VouFewa0jjG+R9JtpIL8x9JTC80rN
yiI0oO8AflPNrLT4lXiXjX+r9nLTvHGuQfdBka4k+/dlvNQ4i9AvitpgwGTcvOx1
Xl+Z0nrgwEh7S8L+iO6r30xRRwKDJErNiSQ2/c3JmtBCoKBfFjSFSXaqqPdv4jaP
s0djRGvgKBQgF7tfz+mGwvHwW3HVnloPR5s115idO1hW6jPFR05ZTb62c9YkBidz
AdJAHTN5S3h26MsV6fyGAauTPTk1k0Lr+hv+RtcBblmNVEaZXWG3kKhE6rWeht2i
cNNVB/66OapUuyCr8YHwPdbQTHvkqLmwGlR/9lpGd1uiPnp3HUh6ztUhsZn5HZAn
RlSBWo+rN7pBPO9NQHIGemnKCpQqkUjEAmdrhWpRC1q60Q0ndS1jtwzFBz1Xhf+f
NkXAE2g2vW/L/DNnMHcxphVrGSEUwggpI3FYzFzTGeLVR9Iqu/zKhVnAwUD6RKOd
Y96OaENgxPuiSLZgUCYRHIGIP5PaVo2a7kvqP66PpGQ+LOn/19qlz6xfrGMbDHfl
M81P8ESuLmhq3mmZiua3rNpqP1TKrtVwBX9JeDWlc3y9G386koCcjuQolTzx1ykD
yQt3Ovz49bjLgrRGn5KogxfwhjaQ81ELG4KBc2FgDFBtbV7I7ERdhQth258RgLfn
yJaDHXNcrYPfOThimrB/tMpFhz72aTA/n726xtrXfQ798SINmYEsihl2TpfgM2tF
Vacx35VO3rgWtmskJ4ybrlwyuW2qoQWgxbvmpH2yg/4StMQZrv2BM4mt21GI+lPe
KRlCISNgrTo/QSbipNXD+QjU12KPX4LHKYJ94EctUzEUMecZaBIgSb0tEvXJxtk3
o/eO6czBQSgTkEdcN9wUU0JuavYepGz9W+zUH/ByoQEZKgMjmHiQU23XDhhHVs9y
KdjDA5GnK4N8k3k+5Nzo1Jn/Fnx6uj8+yQBFChtf2VMN91RmH0O0g9yiYR7rtjvX
aVdHwkdRGUExVibQcR3iDlcnmXtyJXh1L9MKyA4KNoWUWzpzaDQbmzhVANik2XA0
W87VYUQdEzNPy/rvSC/hSl6QTgA6sKxsoYV1erlATktZfEmkRNLJKk4obg5dCgLc
dbHqSTdEtPnRvG9lnQJBp3zW2Is8j9TI4aKEeZfuvQIfYwf2Gw5vOOo5js6W0ZHV
cHY4RqJF+Oqz7Rb4RV8zduESRDGJktGYi22+WdVNsPa3cBUe9jC0b/KCWvUI2kQl
NT2nTQrCI/WSucjOJF9IZ06HISY+J4zQyCcM8K2kKmIdoe5uDiSVegPuNBqhqhU0
CWCgzt3W0+Q+7l3SAgyzgg7FJdIZ1V3JXZyukEccD597aHUkA4fyJOvygfeQC289
iilCeoi7hQ4as22kQLIZQl9B65NAkWgbCObqxsPqB79a55NJ0wd+iWB3zxqSPqQ8
NPYsoGUtcryAOSbBno+3wSfzK6MqsvoRug5BOnScJwXWwKVcZoVQ8+uFovmF9z+Q
94aJlqhGzP0y84WT4oIejwtO64b9AH4anUXKcRRkhm7oZMJp+2ilYboFYyf2rMpw
JEtBbqj6PxC7zuuCsALsFRSZXxWVM2AJ/qln6Se0z/bgkoYNiYxC0kuCm8iGZtU2
kHgWo4q8KZyShut9jfhlKJ+r2vPfz6uvRiVyiephxA85Z+15GsIAqCE0ywSA7UL8
0EDPiaRk8sixvRNNL1ITTBLafnIqAbQzaDxyRKrc0an1+tNjHlThIjIIeoCdnaJH
DuF8BANtGI3HazUxcS/7iY5iKvvPDnWNWVhvb3M7cTIYcCLuiUj5DW0x5UusumAV
c87iEkG0TeIFnM++sG0/wErqpe/qBQnx3RQJi+Rg4xc8PodwsARKwIIcgyjUUFGp
nsoJW9t0zltZaNTdnTxKebirkpYR4El2fCjAN9VATx/rjJ4BVUEEuq00fOqeYCxL
qapvPjZ1zSNXygM0B0crCzgfj2NFG4DQBhGUHLM2/T22+GApSuwYx0VKyc8Z6y+I
IXeTG40xfX1MCtoTYMM1qYmVfSjTAT2K64l2cPRHWkerw2XnLhXw3iQW4Map9T2K
rHJgAyvgIzk5riIBKMATDFGWup9rxTXXRxVRZqoRkPVPDJ03eBz04wja7aGDKUr3
QYVwyNMSEG2ZjzA1K2ovhJ9eHEms4xQUZlYXYvb1LPf1OcXmjnZp2rgvfHLJZwwx
L1ZdPK9g/IHwKVi1bw+x2AE76k/4CveyUHqvZqCrf3wfHeNjVKE5Fu3imw7AZVMZ
dJ9Z5r0UfOSCzBKzsdGrHhzc/er525HIuL3AGvOklEri+v+IxEPr22DzUp/PDmcZ
N9o+cGOG2Ivvz6tEJTrhMveWD2eC/CFI4VwFfXI2CLAoqiYUzugD2CxKpL65V9/5
xn5Skzkn5yBpY1w8sE3BFYhLhlVx71T/jHKAvaCHfgidWC/UlIT1VI6LNVse27Uc
10wQCle/Dr1ivmP24ucfJMCBybI79eSgzCUOcQvyLPk0DAckxxp2ePozNFUm309L
XiQsJ/HvXpR5GnMAqTUtFBkNAYOZQ8o81+pqqGMvUi7JxITo0GwWeylj+hgtrwuk
eSqnn+EAWdnusEzy9I1/NzC25TTbYh5snNTrRVr4PDRjgfxL5emGmuEnLmsBGpI1
uhaBbvrhClHD5OxcBzELbtJULaoFCHD9xtAkYB11+G1dqx1ItTYFX+ImFOkSwgw7
Byb30MdXfmpCpOMmZAw8hOQ8h3rSHRkmZuFJ4R6pDkQBsvSozbgITMtLjxYdRCPn
tzG7rZyxbl3sQOTBoQfDRGBPXKEWslPv2t6yJyLqDU7pfjR33wRgtdzlcz4Wcgg7
xWYrzYalnqcuLGDktlbVFfaKZd8qri/W06GunY+/JXs0YdA4INFan7C52fLanaWv
avoVmICPB8KjhrMC8mrT3KqIhK+38xwxR73dQyG2mqPyDfa7Jie3vHANodO5mxH5
ZvKlcrdC/CyhP35dA/YUKJCrFEscVkE51mNxspGMJhG0Eli4a/5tNtviRfzKjOxT
OrkrvA5UtwT14x8yxVSNYJ58ILVHh7Ypgva8Oe949RAtT8t/YekRunxo51aWZLtj
FKU6R83QJjdcOaQOaxf3203JqRSyiLMJn8GKoqNbB57MntC5zNNVy42hbqbuRn2i
dNSCGy5AUeJdZdQR8U/cN06aif1/fB3stflVCi5JLoh3LMga6Dsj+1WL+HGTWUEM
dzZz5Tbdfx8pL5rt6YqdGGc3tNU4o1Gm/PEpFAIdtriRrsoPY8hmMXqFvJgATky/
VW1a3fgRZvhf/EtGFPVea7uji2EvC0OpISWHKCEJsVY/9xHwOHrN3eCI3zs6vUap
MZnfn1u+fyOKAEU9lX5DJupOYOasDScyKhBI7yO/4VAF3JEmp6nv+cjspolpp3tX
YpJzl6th9K4omz3CEsjzKmeinibO/r9aWUgT9/TbZTLY0EjXpHxbCuqarz1yKheX
EyGkAYb1fzxslOq/ryUv5w6lKzfZ3j7IQXyItTvCeVbjP0ZXJiGRu4Sksz7xevP5
VPeLgXvyNt5fhRC2sjTRn7HgTJKqfhtOIj9kJFnyXPH2sgCqcZ+83YTW3bWLGaHK
jsQgOxJao+zR69RjlAjyBEkX5xV4VBzFeI5Qkk2LBjnqud5DdYVgb25BWC8Es8Ab
QV3f99AacCONNi3cNycnKLyKyaUeKppUcEYlGwnH/dB8zEYakdKNuYR3u9AEIytt
Jf11sBdpIhS8Dhculrxm0lYo7vh34KCiKPMG/+RuGAup/sUmASyWmJ4C2b0cw/Zh
hJs5WPPDmJA2zT5QbEnFc+3hgUdaNsoTEeh6L7pcnGQtaGdCkDnMsZVpbePlSCPB
LUxYiRKhRSlcb9KKbkFyI/0kJZSXuq9Hdg7NTywvW28/JYKLHpplP4tzH7r4FdzY
6sFHludPaWQq7F1P12P+BpU+wO+mboMlzgUX9OF2biq/rkqdv+6wPxTWIoVyJsNO
J01T8UU+0ZAOP9IT2enfaiJadaWp36a2356HtWxqgF6LneTXi0Zt79DJTrKJ788e
hN2f+E481K2V7oorJ1buPkQ32HqCgs6+bMp2YakilsTlU4nkRpFBbxq3pllBvW4a
J6TbHhn4QC7d8PpeHsobUwvUjD7nGOk4cltVvz+lyQbijKDvjP9L6toRdUHKFAbt
pDUdR+aUAjn8Zu0zzUCdX6DClEgtbdf3bmrb4wG197oSOEkaTrXcLKuU25Fc3fDT
CdCu6gXXheGBUU+r0l3PZ++6v42fGWlUSixBm2+5utaswe4uc8BaDVrhOTv5A10R
ZCMoKpaE6YDkO8P2GmJOIqAEAcFZmkMGeNuOiPknXyhshpEfOKkxj6ulFvsSq8Vt
pXXhAaXLP+nJTxy4jv24p11ISZbpfVERxsVC/QdXnuyl3TKA5+5/FQLuivH647Zm
MFjTDfRRdltWKEo1Bd65AbM0eFR+6QdBFR6TXjl4DllYJ+nSOaGg6GG9pqf45fwQ
XajOZ4N8yS1HX0kh3bP05mmZ/37i0gAib23HGhHLkZrkCcIQpaRsO0ohEjbRUC3j
v+01jExYgsIKUz47KMD1+rf/EE+uB43hNTkYGVts/GgetbLVhFa0zCF9yEMMC0ze
PeBoi+hYF0P11m2IZjB202ToUdT9HFybzXVgipz190CqhkE5h6KU96Z8EHnrDIs9
IfITEkJqY+McxnhdkkEL+MldIJ9iEY6eoYsn+UcfkNGJV+GGuxF+7McCmXAUIqeI
niacd56Qb8zIqI8/gq9EtjYlhS1wuOq2t5GfBFJS+qnALXJTF8l5XjbShVik1+N+
dPYvncBc+yYAoEEw8bdUnZxJB2C2JhuIpEQIagpHtCqqJia2iILq2u15eLVQoM+W
+R5/qh65hlkonv1GV/y1X/5dObZNVaRLj4VVtB+MgGkC3ZJoY8IHkUB6GwbSrUDD
Vay2920JEVD7B9jY/Q3egKjLVwWjcMAXHBzlEIiPXjLt6KL9OhCayf3YYFMP8SPS
yOtXyBhyJbOBqmRPU4FEt7V6kJOAl5oIkGKFZHKgP/ohupkFsJZkTPeJfkN007zk
w0RPYzqshhvBQPAZKOj14Ms/mtWyQymgMlIxhn++yB4dY24rfjIbSFW7lQURIn+r
zobn5KSyb56FVye0s5R4syVoiN2tOmUZz8V5X2fkn23S4AmawumJFebDaXMD07cE
1BxyB9ud7DqhAmpThKL/MBSe8B6b8MqMLJQHuQvzxb7+3WPLzWB2P8FC5qwMZsTO
5KRIwjZIrFqcoH2qsUIehGwt+XxnDWzBrLM3fMSpvuP9DSTfRv9sIF/EBlo4qR5X
pN9uRruAO+8fZLryVuwo5BUgvqA/qbLJML0eoRVma7gEEfcF64j+/WPJfTdF8Jx2
EsTTL6VBx6gzEMcBFXWoHKfAvifdamt/81H3dSy6gnlOR8RnVeNhH93k8ZT1qWl3
M9bAKGn7OfT2+dc/5os3cJIkMnH/Jq2PIAu4FsvO7PxgvFmkyGJpUtJ8SzuLysyU
oUsFyKwCmZV2AsB2s93vhlmg2Ej7/6wyPMWml2fnWN6bF8Zjr6NfkMPSylMckya1
WdpBCJ3jX7QKOzNL7hUKof6mv0VZnRtLsUqkkvXaPYZZhqkTMZMxhH8Tmly5hf6l
OVY+d6Lmt1j2wxSK/ilbT614W6BdwnXTUomZbXuCAGDUF80E9b+n2Xb8Qez5pPUS
HMiC3Dl8RhZ9MuKWNMc4V7xVo1OWuirCM/U1o+CSwsUruPyXyS/Jke6TENWxtEy3
+idjXkF4pdutCzZaSTo+iMswnA5K+rReDbk9E99+VIEl2Q/gm1pAJkg2p37cvr8M
vsra6oKfY797azrMA+/71C+QTlHnrR33EHJniYjUdR8rOfAQlidHl39g0bDiDGgB
PqFoJJ3lzXuVYYVgujrnbPqQD5QapW/w5D9P61qNnMUgY/7Q+kgn9bdlqO2+ciU0
kSOaXk4c+ag9JMKwPFxIvuCMJLZe0/kZIm72IGK41sKFefzR4Z/yN4vDOEoIvJq7
pE0IyuW93IswXlGPjZK8hgto4LHt/0mVsZttJlb+dlEUBYYW5gcyHES9UgcAkw8i
5erUeTzhtnYqnD4tNWkIw7DgvWlqbupGAkgmqPG6YPqP+MoA98dChr87M4RtTICU
RxSFrFb3oh0w6Xe0h40B6uCdNCnHV1r3RjXuWIEHlYpJ6wfdHTFZLTvE1Afl1Sr1
VaA80iOTCF7WQixnti1f+Phd0rJ7RY/y+HnIVVJfztFx2GKZfLot6i+3jd6XVT6P
SZULhWx8KUPzg3z84GN258zvzagSrwytvie/Og7wDBnya+unkeYHtCuYaBW71me1
HrWQoO27ff9O+ezzDk+Eqgsk+DbM+ihnvbBi38mYFfUkMq8mE4rf6TUOVNph3m2J
PN+mOFrXvc+z29c9ThXSi1N0yuJzU14jVoVRI6n/3k21/ZwBbUL/xm8Pbd57UZcl
1+I4FpVgvgOspXRm3qXi5K6n9XdIR3a/n0Gw3Pi53Nf96zm8VWnFbKhYT+NlhL3Y
hDDMfzsv8nfqveoTijmmEwWp9fUpshPQy1P7dJCwIO7tSkkl08qnNX7QmGmy42Mv
hyIluBtkfyrNPM/ZaIIY8KJMJZRsY5bxapFAfnLmIOlkEInNF4Cn73CA3+m0AmB+
0KCHGbJwvM5AKiRJTan++k41fJNWeL3xKVhVzlYQDe95J8a3Hasn0r1oCp2c5SwU
u6sh2rN14zcpUpSuZpWGTz9fbKZvjJ4QvWuM2ZUe7Z9WjDYJF6i00ViG7F4X//hy
9iyzjw55GEkL+Hf/PkoMcFpVoMNqJ8xoiG1kOl1nbviHDtZn18PYshd1AF/KNoIh
YlDqkXE8nckIUcVB7ndsN2oWvelbj7eNQq4X4KldFfdxZQwUQSrfEmrp7/ZWVtQ3
keIhNav591KSVdquNync76SQrfOl9DeML9tK3nOWyPp+kYvnJ07jHE2UN1PIyfaS
7L+q+yclP+2iNvmlibpSIOnWk4eOVyvC6BTGc88ktE/7jabHRWnKE7COjY/x3AH3
UdXn3Wk2vYTWja51iCLrYESDR47JQOEvQazJKu5vmaG6Zykc5MRFxhyLDY79mHOB
SUjZpSjiOou588ZiB+dvlo04hXpFmgOOThK5hAwhkHqky/xfGM+CSBMYECSxyY9e
tkS2iae9xCQI61sahRAIK1X8LS6Q5or2/NZKSr+dDR1n6IUW21yOxBPa9xw8p49t
9wsEFzJxX2VfQQF3yAk2hLTipuO6Hld6aq30lDaow44OiMl6LJZNaPWrHUXZMNpL
Sb2EoOqeR1BIPgvAETwp0mLWZnIXpXdri9qoUfsEUpiU1djtq3vdyPU8bF6SzRqy
slpIMHcX0Ah5zUUHn+to7KHaE+/iUiB+lqjgmkaHFu1o/OZFbrhayZ50f5qwMQ7b
tEsLZhtEFZpM0B/xqrjyyTv3HvMoCM0pb7qerYaXeQioAM62AU1LHpys4mrMA0Ui
blk6w2fiQKJTxNsCcSAG73J2igqsP4xMh5S6OyoAQsPHrEOAAHnJg0HybnDHwVe8
UKiiR2pR5nMPM+xAn2XDRPwTd+iQDKoo1m6dAGY6QfUIeEuSXgdxEAXYz0fOqYH8
eEnsdk6QtKPGLBx0VWq5wINk9NXYupdN3qJ75b9BPyuNhy/pq9aarUDZ6W8lX+60
t0CV6EMPyLGKAyfLL3TmhSRYeWWZmfPFh+3WZRjqwcEs222Uln5iQCyY42HazLAU
vlsxp2SMmu2OKkhv1xNEZXaMNv2E7tBnl0jeWxU+7AX5o/ZEGgI5kMVhT+iVWz5q
44GYK1DLzShAKoodLtoks+VGVq/Ql9NluDOGbMF12Koucw1WjNoB7NqYbcop0jtt
zqm7xJanaQY4ZU8HLKbmsTVGH0319dUSGnEqDf81lzjE1Xon5qHWfyw/q11pX3X/
J29/cAe0nL2azMZkrNjlDS/aTJlSrP1+w3kMueydi+9+zRXF9ZYEWN8vJVzGCEHC
LGuTTMk/9M+4TkijIfTEpCLYrs/MVkaGyrGfc4oCSfYyKI/lowFdeUStAqVUewrd
bX53SecsJGOccr37oHgxHZZBgYyMCXFp6WvO9gU/krjEetaclRkyS7CnhxfQEFUl
6S+h6RJvYfS6m6kpjngl2GMtlE0VR/R1fHiqOlK1qR03eZrMUFZhe7QxvGkJU0ok
N82Q6bBIv/OGmv+EcJUz6Dc6UzVYchu3r4vRD8UWYjYXfQW66c3LYQuuXpKx6/RN
fB2bGtTG/zxXci1E3oXDLMwkOPS7frVh8xSj0BiLEqbrJnWtzhXBPkpiol+oPNCb
vmMQSyU8o5z9C0sUOz+N3Yu/IBnpnVIe5K2e/iZNhzGDr8IHfjpVW+wjtr96DH3+
79nHF4hc55zD5eMr/7zigJ6qbC4Ws8MfjC9QR+D9cpPwvQJDBhJndGSkEj0+OwWv
ncxykeEnEz20I/K+ssiBNIxQTQb3u8CC9ktkpsytMlf3do+lLtDc7yQD4Fx3qXuG
EWhCf7oNHPPw1mIHuZne/Y/C8SHXGcxX5BXzY0T+Y0+VPSQVrdRSXZJQArlKO8H7
5gbmwaPvtdbVs1gAgc1mX9HtpVEU3ZvUUrlwtNXRKJ0PkdBxCFNIezr+wRZEZ+5h
ZAICoJwEJsQk+QNyctw23IGn2IhA4xABGg6GbNCMuMk32UCCh6D3ntZVCqdxSIPq
gS6GOuZXl02oWf4crVwLXTniictxV6r02uKUeZmlNnicgsL9IR5hIk7Roo9fLOMY
tQF14QMnplX3ePkM7+DmAZVHD4Yun/CAdGblXX/fY0yMj5ifVmROH2LZPAZhi08K
Ih0/vwLjcRD1igVJF00wl34WHb9wnV79LC0i7lJRBUarZlbMiqijG4S9eQj9rWqE
shEMlroa59v3M9lMoPqUy0EIzPwBxoLzQ5oTvrBjJ57UY95zZ2yFvbvvg6a9YlMx
qqWcel2CkTEUr8JR3Usi/FXc4cnyCKXENxu15piP6282JHXTqPEcxyCp1TOOWhC3
ZVUPQ+huAkOyePW4XVP4fS4Ig18DUd7az+YZ772tFVVWKmVlFX5WZjAX8UynuCTP
bSHsgAqPbUlPWORqC/8hjIlrceyUSB/qRf2GJ9UThkSxShsjmsjTDT5pbEaa8Mxn
Gv/ETupJhprVmAj3SDvktVwwoNcxa+JZKfm/JllhfAPaL7ola/SxtR8W/e34tnb4
1EtWBSblRj+WHhh/5VdUD5/rZN9ZzPhkT+GprU7mA52Yqr7/m0/ZJa0d2f9AOuIL
9cww910CZPe8lRZTN7KDIJ9MBkE6oMx0YVHV7cVNuBwBvZegdsNLa1BBztdXgKlA
C3A6cRhDDFWpeAKjkzQi4idosCucrYpzdFJYjZNVv4mnXPy6BiUU6jbakwMSMSif
e07ew/ejV5xv1eiVO7V33Ox+ToOadjtxqnUaECrQjyb3KCBXuPsb+6zFENq6n1bS
c2BnbTS909oH8PLJ/WbuTUQVlNbrDjWd4ePEg55KZ74iZMMh6s5HmI2Lh6xZJS9d
WNOOYb7kCjDp6Ke7ATuMJCWtiYqecW+t5jC8cyn95pWCyGIUB8R6ceDFG8faAXo9
pAZq9mPWN48t93NwfRAxBlIYjtaDZy7R5LnP32NaKXiLp1IiQFequ69gsFqtaOZg
sk8xjZaEgmWe8fL2ZQbR+w0PszhqV9kR//RWi1iO0VV0WtcvZobLX+zJ00Z9bNbG
iJcClxt9I3eVC0kxUktTZsTKW4NDmnPW27qX9uJoMeANT9jCH5z+7RvOy8JYC7Cd
xikaPv/Jpxo5aZfd0ElPptO03PpE2VyfmWiJzd2OGcARaHXYnWYWIDYqDEaSPvC1
L/nG3V2e9gD5tHyQEA+Zr5B6DKEWEx7v/RaFlYPJkea54AhE4e5p9Xhwqiu2OFRC
ZNHjzzp46OYdzotYedsyxJaCU1VZw9NUd8SB0QNhjFv4T8TDeRkvUGH1wJnAP+jB
cAojtCag22CadNlAHQhjleQw03eKxdD4v1SJ/ezKe1EWX9mX473RMGEd97Jjejcq
eruo1wY9oalMft0qYYtwi4X6C3RXQzDx3r7Uk9fcu+eZOgrYvIfbZxY4vkU5VSiD
N4lJp2Gf6GWPjUKbxMlgpkz6zxFkLPlX+JlejXjmB0utww1rFydqBEjy7PjgjCGV
wRkzuODtuhm252gH7QeBQ+g9iKdhstjx9+XdQ8nK7PQG6VqM1I2fRkeW4HrS15oG
X1zUcwHpgPKn8K7PG52LMVpco9H3ic1A/1V2HhYx5tYLGFUf6GolCKdk4a7W13sq
XlP8/BTTl/cMWp+fqrcSibSi+89uajvzpDWpTd+LXGjvn6uJYHX9CNVuOdUMCy7D
XABJLW6GqfEM4SCu1xnfuHDQvBie7EakG05D7yZ9H34sUKneZPpOcbmcPwDO2Veg
/RfSYmt2Mc7jdTvKJv65a+j8H/XpVSftwsKlI0YGNuLSX8Yz9MnUzZ+V1lshBWod
YmEmSGk+SHyyO9CVKZfcAw9Hc8Qbx2f1xSZZUW1zIdnw6WPLinmjNfqfGEKPjdbv
HqMerO4kg6ovVoQ6jO8QFL7j4me1wS5CaH2PxoM0QKt5+Xu1zs5xUJIS8N6Zh0ZN
WOR/RITv2gjz9fltgJi+MbFliqjRzHb+xMsRs3CJOrtTjH67vkk5SyQxf/Au7spy
ovZRY9ukhIV+DT8XO6/gj4l9szKmYT+KhAM2YLZu6NTFFGszsMR7JaV2B6cp2SKp
hftgc7tPIWEWYX2IPsY9REUJXYD1TIGpTOFkHaM3HaUG0yKgfwBcfpIb9SH/BHXO
WXuRoC3DQqdr2VsvJDrj0SxFzyegoZxgEPPg4hk0LLBzWAbQPiEGNej26qFlyEnt
QUYDX9qQARW8Dmyo6Gw3aa3l9+ypH148I8Tu7YTAPMNh+SUVJ9XHqyN//3ppIhcC
R2U4nY65lSoGPTUTPkty138AOiWDyM4i01feEnBJ3qIcDviPwd9lMq0xLPwxq6mP
Tqn1MdWLaGxDyDMB+LMe26Gm3OHW7UZJ3YXoTmeF4UWxcvX3DaxJ8HM6jFQYL965
loZyA6fyn2uY+JG5WQLF6S8RxwAu4sR6IjfLXDMjtUsluY6rOd3oP1HZJvBAsP72
FEf5AtnZICROI3YyUcMU2oLKBwqXKGw8ZQ71MvUlKVpLBaZkuGebr6lOWLJeEOc9
LcDfaPOmZvBMyq6SUO5vRxJgvjQjPMtqxPu6uxpZvW3x0F7E+XZF5FSPq9yFNYbb
cFQDwgetjh+R5K47Z+Qj9X4F77giAWh7dn75GSiB6diA/BurtFnYaXsEvXlHrZ3K
bjkjJFHAnck9uHYYBtuw6wFIcHGCy8Z/GBVJNZ3vzcaOWYmier/+A7aBD28G97yV
sq9Vbc/4BWAHtDEoB0+IvncjhX3a+YTxMUMOy8C+cTcNjkCPoNHAu0OLFTGYq2VA
1FvYmtTuhbHbTWvPnd7Lpqcn5VgIk34LZmcM7Npkm/yA4OMeUH+HAaZ1KcqCXODh
Vqitn5vNNT09KxGKnpkDww1MM4LrvztUn92Tbb9Xekc/Co1RnR44QXgUwTeSzUOR
SHmSe5LUpLUe8RO5rD3L9LimfYMGAPnAVP3MWysF8Qqp3D3Qor4RtcxzIF5GZGSg
/Ltpyh8Tvzt4jLe8LwCoFbegCDOT1ovk63tyeCeP0HaQiYjuCuwmVqGqI2/7qza0
PMDHmeLxpEuF9tsJmxGqSxs8qu9CbVDZeGZ4KTnlz83U7qEng8b+YKyVHhVByHsi
kfo1JG9g5Os/dwVtc9vbvrVXZmq/Nsc0eXAcV/PbrANDq2jWjzNu4F1JCrDOv007
SIfUikg7DrWdQ2uE27SR11LM/9O2WmnRFA2JZbRTNME/I/toPK8kMMvtsE2TkCRq
lGAmj0Pj/HeIiUs+uYUJe/evM74ylxD75cO8j4TgBSDG0f1IM7fL9OfBvv/vUAsv
1G7H+Wf7mO9aXJd25KaMY29299syvBPEa3uMOCdhsDW57ykYRaJFS/e9wCne6BjH
4d1sIpSEoRh9jDHCh73++p4JjjjKR1qE65pJaFt3f98o4OE4Vaxyl9h1e4mkRd/J
Cdbvj0y0tVAaxEyNlGj1MCxCFYj43VJZbyhEzQ61oqon613wWNwpkr/E9m/B1YrT
FMrxNHuCjh69jrdHvUY9gBykry7JtqShiA5j1p/JdAq2imlO0l6hwrcmWAeu92Wm
3dy3lZ9F6W7rnzk8Ns1cWsBGYwjJ63R0H2fdXVL+JVTtlMtt53itAAsSog3W6hDa
7ZzuAeRNnBTw2SQllaajXXR/+X9WufKLDgP7O2x8ZS1Cu7hb/hxO80X4tmu+aODh
oWHb+Roow+mUhuqZo4vkR9Guh3Dxl9+zMDv8WIXrpopij+1XvZqZ+zZNJzPv583S
S/riqtLDz73vZc2LKOEfnHZKLWyT2aFvXec+qjwd1+6O2xqEYjloAtm3An1xlalP
cU6/NLKF95B1W558zAk7+06xuaQBG2xFSops3uF54w9lsstxWZb79AW+Zr8k6QlQ
XgBnH7gaUnSnMMg46lYOcgipWrBuLlE+XG8QdhRcuvcb8EiVh+Od9ZPJ3AIYOdmy
Q+7iyp8ysXIolGOKKc7+Uu1hflY63N3ILVkJUV7Q8CLXwP082iUAbi0bszAJHfLT
2NjroNHsbyhFngCv02iwzw2vA2qn8KEYCR3ju8IDlu5EwVoyXUopOEGPQTZMPh58
sHwN5OhrzZCFvES3an3DB1j7w7NuJ5Gdige63QKwL+wzg2kugTSMWd2oPPp1onj7
D3cbZvjNQgqLnSzKE/PfcGbK9J8pW0MMzPjuN59cOcqL68Rb8o5CHKZzQ1Uq1P9C
5lFOFXERrBUaLblRdLtIKacqyqfEjpO2em9VyFJ7f7WTkQ+idJKED8dqIckJgDT7
a3GdSJrGKuketcX8kWN5l2VVMVm32m7NkgBGptVp6tGRHCyOd0HuTcI422rNFhNt
Fc8428YkU09bpOgBG0v9M6o8uklh5eTKm2E/B6BRT9ixf+pilXofkyqP5fxID71/
zXaiarj6sVE0NBLrkslhoEMiTF/KF9RfQfPQpwSePYpqcZx3qn+Fj8tBXpjsI4Fg
p0rG8qnnIkE2YUUxZRRSs1UBUWEWABDj71bY0KBq0drHoqEoF5nO9W1cMUHG+Xrj
hFLeuZ34wVYL0moW5Bvgs5EfWXCzY0Z3K3K9OnyU4HoJNXPM+8p9fzdwzOBCjaiY
OrUAn2Y1H2CbVHvqzQFHGioqnVlU2lDbrUVbv37aM4Jzjn3vm0bGdJ4xfHB7OEXT
kKgKQMILA9QKVwSFWTJsdvPpzIPelQpo0xur6NwYWgg8IOSOmEzkFyMY5D495WJo
qPAcT7vImkixOZrgcscgFXsxPwNu/6AcqcWz8J2FkVvXOvZpAqCcoyc0hNGfW0aT
iWfS63rjDqlncyAW2Is5IuEHUJsBCkS4yMEqsEiXu5Zsx9eRlcn7lFqhHjj3p2dY
ttfAe69rEYb0YuJE/vq264cQ39K2qGTPSxnXkPNRHxGYO2DOlXCpMt6G1Q8E88Pv
G/KeiiXwsywWvj0PzQlkwQxHjeOdwBiE1zundau8zma+ZBKOiqZoyOe5GTX0HtJ5
NcAtsc3v5sJUGTSg8GNaFXrTybrgIP2TmJvPFInJHr4Gvw9uCmmgfNShFVv+XFKf
KYtSfp85DE1D82y4+H8fkKZ3h4D3o0kYjTLNneBmWaAZ7AMwDQV8fHUVHjtERFmH
3VmRYAw6247CV+z/6VqCkKdqmH8l/5oaPWKDoWcslQwd3wVWbkCx5c8YOJi6vTZS
zp7mbUPJemv4anaZNgJEHQjipssus8+q/CaFZAHcQ5nbHhsM+Xy0vhmA5U67HHAY
ujrceCDQx4HC6y6ZFa5Ypr+RUBSVf+9GrHwf4kbxdwQjOrZuaV3KfYegsiHFuhJV
9rnJrm9ONIV9XGIcM98eKADpY4UncPecq9dqfdkFiEFWONmFyp4HjzIPRC9e9rbM
YHG+MNY9djU69Pz92HbNJVsDO9iM9NN8+TzU/Er6Jh9cSc+our+w2Y2UJpG3popS
os8j/ZYvIlI05foX3bz9WWH9/Ub4b6cKELgJsvkGPn0d0XJYS/0YLHsWlAXBcPxD
eY774vmOiAqb3UVjAcLdxSURsZrvGyZxxuAGYDp8EBhUjBuz8pEmlhilll0YoU8u
P6cWmX0YpSUd7Z/yM+tlEsIdG+OxS9c7M66MljLx7zU7CY7D5U867WDDnTntZnS3
79bZnV9zuJEQKgdrqQUoD+w6eC32Wk76uiDZQoBrX6lClV0Pj8n/dSTwBXURSyN5
5mpFKmiZm6xTwfsnAoLRXI2+j4FBxKX2DjtxlML6+UuBLf6rHk+4cAq5q5fXwy7j
NAQOwaugZkh33sPPHmGq6RoiNSLtJlaGLZkeTUdi2VKT5OmV1y6fFt2ezUZH170a
YiCwWzhb1afNHypz7qr97+jtkAtqqhVc3+AbM3CdyLYUi237ir+ULvbtDcoMDzx7
DQKQI004Sm9B38JKfdhm7UX94krO2wxWg5VDNwNQ2cmu/fMBXMDm64zFloLG7v/g
ddNwjGCkJlJO7Vjk3qwnl2krxzDaimlNqiAQk8y0srBONCE2aIjzZe3IuUCHQo5p
FsU4h3t9WiXPIUXO5pxaB7+JH6gqDgAq0nD5guetOgxcZqmCJy1A74REA7Bo6rAn
uonxGHRRKGg/N9Q5kJdN2+ANgZU8DPxswOI3gV+CFea6Nt/09tk0sl75YhkJrBPP
7WpUs7vhI1y/774ms9K2/3xLmbYl5+obbLaVRQFqB28q9sw07MIxdH94Q0OUy4Vr
LEzPIWcxlJANNCzLTQVpeoxR87UWT99A2rhZTBil5Fnh7g7z6/67yWDtRFRdDJdo
6AON4txiFYF47ziURrMI8aUL4kHL/9tYqsoGkmDTz0J6sHLQBzvkKuc1oDXHtJV2
vtT0Arm/YiTOYnT2SDHYTZAr4UKFIinm/oY6UibA0R+inaAMY8XreZu9kLW4BGas
Gk4RoHcvPGEKGmPPawslRgRUl+Y3RwD0pfJOjImDId/ytg8vi9NkTpOzMVovsEks
rYSEdsTDib6VkyaBks1D/pRhAst2NmR3u7bCn2VjI7b9QJmXQD4sb5b5qTa2CXjn
VdNxlZ5IweFHfRULM73ROuEkWVQgpMIquvTL1PeIWpL/q1DQ3h3kQl+0Fomz/AAx
WwHYS0r6UYdF4iCgXNIXCtLJXjBbJu4ZpDTmZm3VnGHxXqI03AODxCh19xVidldl
jfTPze9pqXCCqX3euCTWkxHHB7OQ1P27dd2rp4UlvEqoWpajmpt8AKU0kBtKGCoO
22fYSgqlo+YfASTZ50N5CY1Z/ZKyKsm9i2vr1Iib84nJdR6y8pD5v4PBc9Vku49v
ZW4PTRDrxoqeh4ieqbDMEu6uean8M14+pq+w4MNdgtrKUFh/JgI6O37oRfWJjQcr
5BlDOG1Ak2d4yhjH8v3v29maFhjeygnxsTRuHJN/jLbgmYA21M9rqmuPDyitGJ5a
qouZisMrJ0CEhlg3w15cXagPWZkgC8LSZCCs7PxzBojZw0kD8CkDqRy0tsE2HZbt
HEcSuMdo8k/ttLMn79Q4RBnmaPPYGpqGjmUpjRk7wo97BMJ1mYGI0YcLEzKlKnTO
0/N2L6PLeBkutlca7Uh4uS/ZHUuWQ8FAZrUskB1/9UA3HrxvHC9aXU2Y1lcINGfW
KbJndWI7uzyfNdo808sCr7+ku1scYot49Wy+Q2oHAWy2SfGGNIvXfAZhdGhX+fL2
4Ha0+h82RGl3gB9Rzca+u4CO8iz8Uz/jgd8Ilp47/cmbExAxj5rddo+KxdSKjA+l
1ZT3GklykL0XWEmUoi+golfd+ovPdbRpxoEQDZbnNxozmMCQATld0P22/3tPAckp
W0cFgB3eZhmbHvhDWz2YowXvjRCp2PKHESi0Phr2AeMUWZNteaxFX+KbPVHfuOgR
rotucsAHih4MDwxy7Wx1T6VCA91Ujjal0achiWb4S18bq+ceYn4sPooiRiTqYFL1
ZYzpJS/CHKITGJT8p5/tOwN8s3EarXtIpQP3AY7IznU1HmKF1PkhfmXYrYD+qeW8
TcAVLqdhIkCj6uv4kY4dOcvtXrxiFg7GQUXxtbCfZP03X2Q13rspP8ZLYjBce21N
Vo7Xo22HEbNt91RKOptmRRgbIx9JdDQNKrjGfJ3u7uQQHyUvgOimKaqBqhA8zUg6
jCwyBWkEutvnLlRTqFDbfwvIVx/gBEh6RaLHjx0NqVMONBTp2+Qbj7MsQR+aAduo
vl4eGK3DX6Umo+ITY9VSJhAO/alHofJSkFAsYyqSCRYwCjPSdmIC6tvTMEc46PrJ
DmLn7CoxrOFxz8upAVaSe/zV0wwMDTGvk16Ogyq5jYSs7czLSgZq2CqluALo965x
VyO2Zs3wbHcerRrOrmXU96UU4NsEcca8H0XPbJU5N8GhMySxYR99Rbh9m6M3aV+0
ZJMx3o/Sh/81vXAGN5iXpV43pQwgS48gj5nEPwGoyJFIo+yHeqIsJ5Ix/mU8OPqN
i+WoKpf34P6GIjz6/xYAR1lP9lHQyq1u2Ms5zCoe0HTCOkwZEJcLVLguAeijmV9h
vqhfN/lzSbbyy9+UTyuVqIq+6PRFQoSm+TCYaxD2taVhS2sXxCBZ+bgmNktsgNEm
EVpzmEDgJMYQaHUQzgIpgwvJSOMu6pWY5vfL4+3drJON0OBRAm0Qs0PR4SW/87Id
umRU8CzuTMDiMOO7rb3M623ey6yoOwrTGOW9/ymAdp3LxWmVUggTkoJoeJBT+Jsg
84h65l+fzN5Q5JfDpdvgE10Rh97tC31dzr0VmRi6RD8pBlqdceIV0hGal+yjYx0p
GNdopM1IsBV9WvPyReRbhVLHzM3XfPOgSJ+AHRBh6R6ash79d5uIpZlW+d7WJFn4
p7KoOCwD53T97GSUbu7oPftBLT/N3VK2E6Raov25qklFB5Um68ERBDfIOryxc/QT
aO2NsiL5YOXfOgxJBCHNQAJZehhE3FjLt5jTC76kzWAQqjra2FQNPqXU9sAg2HCq
gdVLuEi29xWRh3PcL87qrYDUe38yDc21A3serrvDH1IiUYbPXUoUYXGvr7XSXMdB
2KbKQJAMSuMTBWEkAw6Xtp271TPMBieSxXvF3Z/GVuxUlfzvA/F6DQ+S/toLeT6m
2TVLRsi8cyggvKpoxbeYBEMMzGrF1hjO6DlncIydySp5LwAzJ3m1gxXBaCVgiQrU
AaczXeizso8sP7tfE5YPWW3+L4O2+mdp6P1FmWByHtnblgrqYOHBRHKIQ2jRjTXw
bxgLjDQFgrrN+UtrQT8r5CTiO5a+KKApd4MwseYhXcp1cQvunTsWUVd/RGMAKmTB
KNq7z1jBOtGUK1OjqeZ3YG7apGkIIREcSPXkrV3ygW3B32Dh95qwaCNQqOuBLBrm
L7aAOjOmZPiDwxkgk/Fp28SaloD1X70S8b644z6q3eDpgo0NPmKcJ3E8LsT9QMcd
F7Q2YvdMPvCnwxMuNdNXeiiKtQSY4G3QwAxTTHVkk17G7kDazc/epuscAAV5/T7m
xY8S98bD6f9pkRRYLkSFu3fJ12hPwciUv5aIz6MPJ5Xg3KVLkooco0i30pK3oAQ3
gHxRSEHBdLwwx+DX4XJLJnLAp2aSUm+BeV8NuAAQ1uOMs8nHznGewSU8Ydhz1hXh
gLMvxikmPm5M9KZMkGALm98iVjXdFi+2PsfT/JWjydIiwp+CLZHsQZjf3iKgKuE6
WOwxW2/+RRWcaiMw42haNjPiZEygzFjO7qlffMW3QzSHn7ntzWv88oqGc43u4HKH
9ydrB2QZE3FFjV0X0VySA522k5+htiEiv7B8CMf80L/ysHO6rlOHpaADmFdgawgR
Rt/M3XilGYCZh7hf+sR5DfyvHdhfuv6zgKQbdQx4CnVdWoROoIv+b2y+/GOuQH3s
vqj0OaODbQKJPdEIDrLSIVuaNFkuymgwz3tKSnv/X3mtNOMtSd5qohZxiMRl1l5x
9ZnQxXUQUSVHBxO8eQ8yjdoQwDst7snSO7yJOgcl15igimT5FQXH6amEFetuQloj
Y8vG29D570mFMZjC43G3xyOzdczcQng5lNmZ185CDyCEaoRiG2HA+r8UCuzzbjCs
TmWPCHBSvEkAFyV5FSifSCmzIujndvsg/NzD2DKktSx/b2lW4TXzOzwshs4Dfnur
c7l0uESvF/rAXub0RvW8WJVSHxbrgsbDZVS/TBKGVYi6uPfDtZds+nBeos69Gu2k
g6ohhLDuziXX1sIi1Cw9rXnzB9wSGlFIaSrF+5dxqGK+T5qeLaO4YB+Zn7H9QxNR
gXCsgsR3ckaraUJXNrVZTiJ9zOQkgw8f7Z0JZk3TYe4+VYUHBm/5BTTbScvoK6jD
bduyIAEHDa5O/d+z9xGkl8bi7SFtLYDCo0KLLRQ86PaOaoZDhQbboOw+gL9kxGmG
HmC3qUkdWY6cmcn40s87GesJwb7S9Wqd1BCH/FDHSYW3LJa2XvOv0C2UgYGWqsSC
QTljMQJ6HIDXWY6GuICk8/TT6dCpH3Z0J49S/L9GjM029enFu8jy7pwwB3EefCZo
2KU9msyuxSzOo2Tteuo3gEuuyg9eFGp3oKD7zdF8IUZ7ntmx1WVwQ19r19ftsOPe
51JJeBiOkMX2Vy/8E5FHLv2kMtXuOabIvq2iVVQLoXa2PsT8JhpXHWa4JrpP7PUt
lYYM/+IUXUXSNUybXQEvdZAvhMkQvpbu3fPA6X330AnCQEVQHt/l9z3KkxiEjObE
4T/X3CWkzjPw3YPOLwE5EBgLaXBsFQXAqEzSs87IJfXPzmCaUkitm3rkQPVPteu2
vxVTjWdCc51P+FyYsNCtiKURWECWmKe4zCf/7j3cKfDgBaiIHiSoZvEwWRKFUKoM
7yn9yKN9ulTlB9c0eX1Ns2ZMIKvzJQV7cvDlcEkzdC5Ldv5h1A5e92l4Wx5fIBNk
c5N6Ld2OHkHVFEp4UijoEjoLBJjI9o35o7HydHStsFcHnz4bzwofEnktKoAWEtq9
P2W5oR9jqYeUvAelsobO5oG5aH6IHey7Tlmp6AQoUAKpFCA68X29QxZWbpFRnWN1
YLUlDg2cZflmURRCHED3vgBglF54ScLky74QOVHDJxvgbG7JI7vlJxLxsewPkzkG
Z8eHb4QWRnVshgIVAYhHj+E3G9Z6JWR5BO47NCRcuxjGMmXF9qbf7Bs9cs5TX/tQ
PxF2EoRhyeRcfmTMH2cFRo4qypsMLSKIrual/n+iLpC296xZZDlXJT9DTImcLN6/
WLJ67ns4Ag/Qm1V1hsWH0J0HGgv+OsqiljrpiXKIbc4Im7tmd7Z2BDqYNREsVycI
R5kq8kGUtlVoPaVb1JmhGT/3dNaw95T36P3hdCKU2DcEdQMo/EzemNwadtKaDtLB
sXB1OagFRi6OczJQSI8J9ZDcGEWMGKqOczb5s1GFgLUHn28k3i81oigq/J63uaoI
b+/OKyf3VpI+xoyqWvJisJbxtP1rCus5AjS+rP59BgCwLow33ILq0ZLKlpWZdBQx
shgmlB5K/SZjSRx+Qst8DFC+j4YpPU61uRAYcTTSasGDjxK6G8jYXRTJ+ekl1aGr
bodGjf6kskBR+uXCWjIiaKfKX2X3bAIfvljRo+9sWbLgwGZH7oesa4o0fsEf4zbp
yxYc9yRvJz0o4b1BFFlnUrvaJHTScABeAFsIEnIztjfkU/RNJMPQSqrhFMWgWIZN
IzWnzGdK+ahbhm/ABSpcgvT4/JmswNkrFT2ToP0EgFBJzaVW5OUzHSXL0n/4Z/ur
FuojkuadB8vC4wPLwzpOkDqWUcFZKCiyePkZOlo77ghIY0itF0Be4mNerjdZtky0
1hBIh2TwgxvEJDUd/zs8aPqMdF/eT2YfBUoY7BVZCKo7atD5akM8k4XZauKckqxJ
wyGQ8E0gfcJkTqKIKWdGmm9T3VxymsfrrWuUOlHLOQWTZapqYXyoxjiEL6dhwrFX
ZeyEhmGqzws6zr6m+iHRKgdwa0g7ivncclvwxsKZ9AYXoLaJNeUA1ZfmdyOS7WuI
WiFASfoZXVvak71uI84VNZj07Wl/idB96SXdFc9nfRaSyctoIpJ4quiAI0RtbS5t
8vvDdDJ8W0ry1DKSpcHrwirEX8Ssk40uwGpLeWR7K0cspI1ks2/8jfouWz+h+rbK
ehncbrSXCgZJDZtOXohVP2nX9vjFKLFXcOX6JoM4dERTjz5AmfHbnC44KReeFlNN
lJ26lT4ZDlPuxl6OBXy/wAGBgV6p2nsqhZbM9oPfQBgjVokSKMMjdo4ZtY90U2Gw
a+zVvWyiR3uQfKp+H3jeBr2O76QxRkF/bQquhAL72mlJea/aVBeER1KEp0L2Ib1Y
FUin4acNKWHV06+8TYBvVPqWyjFfbF3/ifuRLVUxMmQ/LDTdEFB1f6I10Zq8Gfop
AM+UIV6eIazqJeEts3bKDBBHN0A3DMHtsyaBo8Gk+ni5KD9SAQ4TqdLo659h4myN
GSU4yFtsNk+52YW6Kg1wGO7qmvYmvqrW+H3AcWHaVbBncye++BclOodnV0NQeIZC
RWf8ZB/SqFGEZtMhQzk1Ju67XVMOMxpGQjoXXHquHCECJHsBh0P5+Of/8jf8HHsJ
KBUPDPci7nsdmTLlhaiwm/FHKgxhp/47cqIj4nWJRSu1KFETHCUtFKdDpl9n5qYe
pPXY5MhSmnrcgFOW2D8geeMMDkYydrqeSNhImVLic0I3LRzYucvEvvyVbQ3tZaTX
6c5QsTsjb3LN57E0zp4OqPkpSRaDVd1MEb6Sp3cdd9NxqIHP7y2jvapyuQHE3geT
2WEb2OAJpjUQWigKSrwxcIooKTilL8N5D9XQ6bKetp7k/IM0IfNdmcu8Sbp/wOtl
X1W23G/hnkAdBTs5OlNI+Ry36oK9oYWadQzoiz3ur+ttAoV2YrsuaTFoqJuMk+/s
a9qgM/Hy2/m0Em18S2YVY+XM58tjyKgH1t+m7idt6OwCQfNJQgHNBvfx/PSVYcu+
bru9AgyWfWx2uPRy/lHLVR0sVrsRrKosTufl64aeHVRxivXLksobVAFnKFoRJjsK
XCPnt7QpHhRRNt0skD0Csxwpru0rXfjSD+s3peg6u8OGUbSMbFHT7pYqaDgrFv5S
e4+yMAZWitm3btojy4USF2TxpjbbcTnzoKOjfrYR3S+2ATPzEfMqv+iFGEkhz5j/
bHNB9Z9Qazb1mU3J9LkisvZPQ54HDJYARuDs6ivn0JTnRg8G+y1fAfouIeD3y/d8
3BUZ9Sorcb1w0lBFu5mqPU21npyKVhOkbcMsK6dP+oMhQ3ekS+EawfRnU9ZNh5hq
6UbUD/+fEiKcMI1fv8Zvwu0VXkma2sHEUYICzeiqHRSGSj2LbM34xOJZvUS8gkin
oRCZ6L/IY7Zd5CRIgRTyvgklroiwhbQrAO8KC7fwIfinyb7e7N1qeb4XHq8XoNgF
mn07yANilW7mJjeS6szv/4kEEbw21ekwtJW6sBURGtXPzYQfFaAQIeNAfZrAnxZJ
37pI/4t1g3ZleYlb3l1oRNKp14GwpxdSxdimV5ta5pk2Iq9PK7gxDGcxQ/NjfPU+
Yh3uId5lyu9o806ZuDlfzibxu2DLU4p7pibGIMVyiSSZIWrEbp1Qbbl00tuPEgze
PFYVlmxIWZOkkvwm4Ad6Gswe7AycO6VORZSxsZn0mI8ar1Z2/l+XRTiamMdX94B/
Zf5mc5W6OD3vL+8u1jlkXxBhbOW7uvPguDRUXmwMYakNpZ/pwBRwEanc2bA0eNQX
J+GaOFqh9TQdsjT2tPH2kYJdXGX1xnjFIpFSlOc2P73qY6qZr7GQm5OZbj7odQCp
mesefr3ouaCq9XOG0Md81ZcZHJeE3BVBwm25dPePO8f3OeuB82z/UsEJMDQqe2kY
qbGGrJkwieS/thon4wbPco8T1G1DdGPF6lK1GASZj76QjNJzwQpHxIhkJlfmumlz
RorHQfsG/64cADGzFsuOV3VRitIuqdJP8MAsILKpnHQolZWx98N1fu3rqEFzEJYh
FDBpvlDDUZK+3uO7SWHaLdQYiVwLF0StBV3+l/Ls+Kt+a4wfKs/rZUlFAAnACJId
w6jQ2Y9luoaYqWXM6Ko6ckMjKOwLgZYonFk7/N/Nk6SMmT3ZlinghcbBM8VLnB0X
glm7R2EfiTaYZTtZuViJTAgvvn/pkPEo7trQeDbVHaAcsotctAa2gBVo1JkPf/mJ
rGdMsrFGJs9IUijVUNhSQstWr/9uARWSEw9LT9UiBeAhSdjIstAZqNDfhAcdAcPI
wSDW52o4dwvaAPl68KN9hm1Vth3iEa9kmRJewQy5BfVUAU7jRIeLdqZoteMPWOFq
a5mvyCQg0VwdVJw2aI1vK5GqJvXuJdHbUYBF9wQ1babyUkfcWe5/CnKBFKbFVCXo
W0P9hS5fPgTe5isCuIjE8VqZBJ8AFzWDQjqf5fzpCCN+1bsZetmtetdvznOpTGYx
2pu8ANULH0KGbWtVSUMb9IU678zUVFVTGK0ARSfQF9YAfom+kD1Ei6lv5IV6k6cj
ThX5VzIK8vbu+kKd65wDVa4R2xRvZdeNKyYMNNN6maMLcSWsdLk1heE1aUdwy8X5
KwhElbzkx7BHxWDY68M7FXcwnBnVHv+pVv3dKd3ASFKu3mP3FDtwYMECiWRamtbC
iQJ0KPmiWmTC5xHSUsdsL5dAsdk/d2PfrTlrv8te8C7VETmJl0rV++Fvh1DU0oew
k7gjwtZs3etaqFUAEzTKYM68kJrMzDO4U725jdyigyREIRECIy5NXuUL2g2k8EIK
Kba2Kl9zgfM4333ckifrIkpaStCCW41YEN/jmwzFJpDELfx4FQXFVQluRTey7U16
jcLyADZSLrURdNRmX9x6bEXmAW2K5NJ24NC5XrY5tdo5iCgf49y9Xb5lYTXITa8T
IhlTYtwNQ+xJsc2h9GmKEw6Rw4du5jR7mk5fcyIzh/SQTviZBapsCIH4mtgQVji9
lkcAjq3f9YhFkQYoTdfswrbkA+K4KjnTqvWZsZYqndDgJXWbYiJhv0O9A0VEhZDi
5RWeNe0C4FDGNamjKPS3KKJru6zqONdFQuO/b9mAuHZxHMMj7pLIDs0CExWP3bMi
xbzB4IRyENs5YAD4LHRPoCO5RMypCDkM6omuyKYvp8P76F5802u2mCJj7E7Gelgu
idznJICvj8V3m5TGH/uHLyosP6IG96wCIrxce/TOfArJFhIkt9doZErEKHqmRgTu
nM6F69apOYhzNnZ00mcX8CVjN6z6yp599n4HCPekKtX8wwHm1eEJKUr+7If5mQvW
8oCtVK/4Jm6mPusQKlz0pTyxpMD4IRalATcxvqGOJTyurJCPI909U3TTNA2xuEGk
TlKwXxyojFaAIioBPaO8TtYdsHUJaEiN4BW4vev0dGcF4Jz0vPvYO2GDogjlAo0j
C7ajjePQPROdCXPLmMxzUPPW6D944cMNbKwpUZSmUpjjAGJK9q0M/Am6nIOYBnSj
JXZwtjT2Gwt2l+Tk67Ifn1kQDRUUwqCaY3E6jaFQE7qeTBC7BdTqL3Tsa8jr/vQq
R+B50D4Ln72kMQmne+724p72anjMWPrMtb5uVqphh5GT5iQwWcRLc8krHxAJpf+7
IzIDIV4c7naW5dHLAT0LbiDsP0L4dYOuxw/Lgf0M2WjrhpFpydaupAy32HeHEH64
tutCNZs5tmSQMVYZcEognt430svWnxwIhm3aFLBgU9Wng5v8QnCv4AbWXvoeyW46
ZYQ2cIRyoJrXXG2pus8GbPFwEb0c09MdwIMGuUx+Ys0uvW8odlFl0xfoPVK57Sy8
B5MwKPMdAfpKfpDdelViKrlsCqcl68XppOtFxeo5JIwipqTzW5bqbf44t7QRdz0a
lbn8uygn/BNls09PORgF27mA52ODFbm9Iq8LFhnSIjofizDRCcFh4wI73JN1WwkC
8/9vw/AQRZf9KPwgg355EH3qf/6RZDH94jYRZqT5faU9xLGjXsJpYc4Jyw8eA1gJ
Q74LGRQkaZeDennKJGmZy07FS+F6fzroTuafMlD3Zs5ZhPXzkqKWWJuXBejGhQX8
aU5XvAs6H8zaYTxo0mvtgD2c38HRVQXQU9xGz3RSKCDYwwP+8rNtxm6vYgDZGcQh
o9/+/zCtJLGC/YVu6quLiSmsLIOXHnczhkRh3tWQf09JhamYK9XQ0RbTh8fD6tda
0luT8LI/Kwuik39gO9j7CMl/QhsQhUTy6mTZB1dDqeE7wWArVbApICl0vUvPMv3+
zKqRQzutwCmqDm49TN8F//qmf9PbMzkaUY2Ih6kn9zo3ZOj9vkMOT4n6mcnIDtPf
nswL70eSpMks3gQcTWGbeA==
`pragma protect end_protected
