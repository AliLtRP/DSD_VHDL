// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:31 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Bqvo+iKIvMWa6gPIcWYjC1YlwN3SVetPkGdDTgweL9vUx1Bbupdv8cbRD97FqAtz
YAtmYvqEqlb8Lk+QPuKDL1nkCP4m491tUj1bI9MY61Npno0zTpyTnEienUsqXBnd
WUoNGIPdIT349kdCzoZtsYNm9XZDVak5LkQc2rkUUbY=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 19360)
+2Wbgk5vD/xwqQcab3kf4QA4eV43HksdffpXcH8D4VJ1s63KMmrc92vnXAl5gg4p
CZgAuKRzNcZoAOwREUb2gIDj9YJ645y9Xi5gxASgnbKAhn7i0XT9ewRhGnPOTygn
qyWaVgWWrTLjBTCBauDcujhg3yv8srJMxn6cbxcCDFwThFwLaOzscryWZoXcwj86
S7pH+yF61UYEnMmjBd/FPk7rbS7Vq/4GGdKt9y+KfFhUaWDKhRThapFV0xlrApBQ
lCYt3EmyG/FWGtDh/IE8UhtIo78T23nGUIFqjFiHjt4ATAvS74BjkgV64tbUIv5J
VZABp6LmY6kjYgS5N1QrMvp3IWq+Vrd+KXIZJ4dTs4nENvLGiRT/ocWORSVdk11J
IrI7xrVfqQCSfQgi/oDQK+f3KHhMlP8pcT7ttb6s6pslHmDnQo31QUwDE62VRyDv
i4gddmWl/UcwK8kTk8Bqjta8ceL7QtglabPq6Yon7jRoiPCM+rxqGR4cxq0aileE
DF+Ss8lHraiEiKCLydIICW32cW2VXCdI/jAhuIz2jkU6fuZ2GPomdttEodFjy/Xv
gQALfw6RO9aRF1o1tGCQhe0hvCF5nFd519L8aQXYj+MBsEPr8GWnktyn7YC0BMaT
V/T5LOw9BOK4RmzIiAlOzATZiwvpoAjOCBSibk/RktwCZvUdHCqZthOgYW1KHp6r
Cx10oReR4ephCA6S5r9P0KHEDA2aPdNRLil+TsSRvwBgBOmgiky5kwxnwi9Dyy6a
aKR+pCDzfNFGFCB9vVHxFhKIfH0Zo3PvmK9hi4j/JNfb2KaHBP9xHBtiYafX3sA7
YjlE3Dwczvsg4pWESVIPty2rgMeBkrrb5AE4QglieaZHBFqUH92N4c4tOJrNH5sZ
JysKJyz98WzlsLjOfoOo5u6IzyB4zqjqBX3FnBw6diMk/fYQew94Et7M6oadw/uC
Rx9z4dzEomC5iSCiAZXrM9EcuVXM/nPy88CglnEcWh4fgyOB5udcngb+E5Pl+hHe
BOFymZfw5slfe7BKBc34NGdxFyeC5Z51xu1NQ33GpdmqkYxGclWt7apQWm086W58
lCXW56mNlvq1eeC2rQElFVjABGE7XK4rSr+2DXa3vk1gSdR9flbSPU3zvPJ3VyA0
i0yRGZ4uPjwOUjFmzj9ZTVAaDQnnDqh5kth8D3u4hk8DH0Gr2HxjpXWrISWWMubJ
4OS05qg3Pjprvluh4Aa+J9gZRCfdoE+lctF9UFBOWxpkbgkO/WrdyqbpzRdUvDlg
kgLr3/6h34uIFccG9PySYAv1lEdGYQYGxbN/+R/e9Ut2h45Zm5+krT8sme6EySZx
HkHo7CU7GvpNSTbptprPii8+h21KzD/gATXG+MpNR8DCRmhu1B0SVqBreog51Gv3
PxkKUuiLxER8IdGC3AgpB3qLKvh6lHhgry3IIhzdci6maQYhHEcGv7d/8MNIVbX7
ChDPskxjxzeu+Sk2iJVEFe4Octx7ADvQIsHP1J5tYDd5MHlKpH4QD2p3mqANQpkt
c1Vb/VKyvYjTEhdvOyhb0M1rCazIsDJ3wHNpO0fAhnxYzzReL/CCI+wMfQPXHgLp
saH+gG43rTMMbxN8+PgnhqiJpuCynwZX0QP0QUNqGEgeDJfJCBDY+EOhaTHrEpmU
bakjKAce8GzmgXGgkn1KTtm0BkmDGmmM/yFPMxHe9dIoTnuwi2nMclX3XSYzuS03
WjNpyvgTKDuqjCFj8SjqzKGNedvd1uJ6rp7Ap2Ax7blO/9GLBG6SNMp11jQoAeVW
R8l1MMxFoRb86KVg6EX6FIyCcSDSVZot/g/n7E1zFG2yRjZG+sgmC7WEz9bzOwTm
M/0yVHHEhK+KR9IqZWjEiHADQU43Ntr+IcxRhWTxAp7vypKcLnCDKTSE6dVkT9kO
mdtJLXaXsHCDCAgFaEn9hYx7N9+Bl/1OSq8f3epSruEMsho0dp9boteUaBiEmDG0
zRmxgXVjgR2RPG8CndqiZVJV3qcIlmHasrMzZmF/lXdotF+Q/dDV98NULzownF/B
Dt63ht3ALu+Ck6OjPyg69fwRTbhTa3fu4eHSaGGlvpzxUeF7SYkzFJSm+vHZfXZh
+pHe4d/b7cGOt3SnEDbTrr4Yq5L9YCbCYuRCin+sviR6VclKNsZ0ILVxGtciK6cx
lGVv3SnJEYxMf3bueEfV1skh0lI9v+/pRv53OBp56fqTOFHFK+bfqytqRSzm/Fq2
Uq39sNRVEKG7YYeNM+uPRx8ZhOr96tplBdt5NbkmGFuHAGtkG42/poczdZNZzI0l
a2+oawjAQceHvcUDQWjFJ9IfCJ82gniLs6L08PbNnDGpcUQmZYsYfX/58scC5CYI
L20pv5Vgc2FOpYdH3ixIPKtThqmzQR+JIIqZbfwwZJw1wUroYh00zKVmCAxJa4Hi
VnDH2UVKAQNsIWA3xTKL8Hg1mx8HdI1C/2xkLM3H2Zw49QnVbPZblLXOcWdka2iO
8ercC5hEW6OcWkOmMX5uPPDUiM48xL3Y0xLpevBGDBKD2J6PF8sKefygfl+bnUtI
fx6XOs6XiIydp2HRdMg7iamMHTqCaB8wqbEgJYH90NqLh6l5HofdMYrAAB5bA5qk
eF7OdySjNHw4hNcHHanEWf8ryiiFIU8+Doiz5+yuWufd8JTd52UVhcRty8mUgPki
RflzmpO/woh23JZGwDwE4Q0O4YgEw9YDN90mguWHAUCiymyWdUFlJ2OL3KWMVvAO
+DiR1KOCCCtS9QCVr4v114+s+X7oG/SrmKyfjUS42rez6RjlXDK7+9LkoERU/i7j
/yFZnOL5/T/3ogkwmOTvFXpbkJZRRjkD4qkt+pLVrmZZ829K0FYZNQCJy0NZ/45U
/klOM1ai41QRoolecfr3QCZ4SxRkVoaKzF8rHJ34idKszXuds1Zppd6Ac42QLeYU
UyCjcQrn51leS3NebH6HH6Nj1UngrjB+2LukosIfWIe2ObD2VMQMGE+xxJBPLAJz
uySrejtQk1bWCy1hmNfH4lHjEef+8RQ5ARcWv0gOXYtw+fYRpuW8wYu6zmjfCnbi
pjyqROMeciiigJgRSIl7NYgniJr6+O3AjYuTun7IM9eATorg2fiKpUZUyFLtaycf
DnYM2D1og9kgWNSdY/yJIIfCmKBh8v1uDpFXrK4KNQ03Kp3WtNM8KJ+uP3r4OKy3
WkVpn0n52LVDV0w6uGkZ+6153X5wjO4D4xBAY60zprBmT+u/mxdjHcDCgFWkpZ2O
6gggzkD5v1WH7QmNNmDpLQS3J205LHQOlLISaHi2aE3miZYDdmg4TIwNIt64oZSH
D7Ho8dmXo7FoRljNoFeOPPo1V1cQa345ZYbfvZ0KBVqZnB3Ww4o3fxHep/rxeKej
iR7tNBNbfIXPA3DSrWCs2v4gjbJ2O8xKzbeocFukXGUiGsSdNFM17gYGv/4kqnCk
rzFEnTRYplLS1JhD0wOrQ3/l0/bywsBsq9Lt/9er0SG+TKVYXbfkiFq1WTgE+Eye
5Tl3Tc19uMalnoqw4euYcUBo8JBvUwgDYi7NpA622/IRCe967v4ON6K2CGlqte5L
Hcs/gfLvlNaZT+eBYiWriD3GlqfMCfQrD5iJBUCUafDHg4rVl5UytMPD8tBN0LPJ
AlzxK+8bQIs00NrAbbdKnevGmNNcVoy+G9/W3uyRDQBOlQa5DJr9cx38I7gNNR1m
kmn9QA20WHIxPYn+3VoMpOMvuuQVqgk0Zc+HNVEVF3LShJ4gh5Aa5+vyJMpNYazF
wx0WcalbSjGISSxfalyioqKxfPyhfFlRd2CBlgXJmQJ5CsCwZSVNdPKXo29T+8vk
kDXeskdF0o1gxnysbajkZXb4so+MO3KaQNbPvDvy7i6YRyXuqTIbrrGXVoQgHm5B
wX8JmQXnYaL707vDImlKHMZVZDREXdafQ9+oPoruY9bE3MX9KjHqW+aYZgR3p8TW
5WZdndKPpVSSyW6p/Mg85+4NKEjy8kWUhtj56JK/ELEGr6kHAlPXqgIJmqhQbbXi
Hemun7warVzAULY60gMWGJdWFBP9wb9TEyxr17NTIRMlXYh8YXOCVF9ze0XkA4i9
z9Z01Zb8c91kCXt3B/4qmN6b1uiznh6g4KUtG3Nj7Ymx8hxRmIVCOTbzhIaNBpxp
ePRHA2k3BiGndlWdrU9/vSYIRtQ32G8w2zBNDO8jv9PzyXr8wKFwJE6fGRrrOMkG
een3hfF4IWeszKagQmvtrxF5OtOeP7rWukoahoHlVmGRk4MzIaGJUX0dUVg5Nn6G
wQgr6ztTsnVb1/GvcJyDV2eGyQF6nfs3DMTEfThoxzoRDLXbYvR/k8DiDR+l/e3f
2TYOZ/0fb0OHWIe95strp3jq0y1bDOD9b7FLl2YZxAKWaFZlbc1FT06hoF8NB880
g/mxUWWGhC4+lhNpH5h2KURtnSdtENZlJtLAq5djhSLTTIBaRS7lpCOfqUoepNYB
zKK4uH+A3R+wvSNwiTu52paw8Dq4PXqmcnh0WC8Xb8C1hzT9oS55OjvlM3iKNGGy
Ztm3+lE3+InDP8N+nHH2cbKauwDlwuVWnmd3B1iFkHIvPGVWh09pomQht3/8o2Ry
NM5rUrjuhzCf8/5FiNs7uKkpUSzyITNUgGRf5cu+07AvvAQv7O+6mutxyBwQkrXw
NAjlqBnsJspKuVuZH2Y9IibTSZ6y/mRjRrWowj2vcZl6HS3TfV9HpwV13LTG8uPa
VjbHTijjv5UGpHzC+FhT+fbGZvsMbBKjpqgGCVpgIJXPXnCyCZ7peLJ37wAG9aWF
A4Is1ZheJgYnKJ7LKF3V7RkG+j3/YCeInG4j8YCZgOMCv+kjAanzJjhRbQbuTG16
cYBzioOFrsPq4rA/btJzGLWTHHycK+Eh3rzP/sZOvn5LHCHlWERJqZZoozk/Izkg
eB1t8bzgeYEXafWY8kedy9CforeYfGpy7w/EWsxlPgNbaoKgwR4lDpWyv+Td3oy3
IBgAVhShY3u5NRjkl7LaYBhLxF7u1tnSQiotLYeg3rQS/RSEzIY6MJJBVKGLCVD4
HJf9//7Zct2ivDcG+xVwo6J7/OhB7fAyK1eaUcfuQX3fVmXYyG34bNUHd/ETYUw+
FtjuUQIvPvMryo1Sgy/63bcB/Nf1bDmMxdzPytBv03HgWKsgv0yaqYFH/ntHYyOt
5ESpSmqZ+gMH1nOMMAWZqP4LSWyepDeh5rPUrLysDl9EVDHZeTWskCOYJK7rNzdD
hjCzz2rTuTTbjgFE7/lVF4ORWCGHjsWbJuAOvfpFEiGBQJtdrHtElfDlKv2KLfTg
29Vbe7m6JLH6iH79Jp4aKyv7lTCHQzTChzRiBszhp3bBEu5zlNXBnQszEDenhjfz
Y83pSoypWlSMaGOs6xF9/3K/35fhwC560PrbNgo1siQvB7nuqwtdK5FsvRwwYdEe
Af9KS3jnV9Rx0nsDXfrSV+ZYpxqtLrgAk8vbCgu7dphEBe3+rhwPVFAJ8KQ29+Xg
jtLofGK7vj+Bi3yqd80TCFxPyC8hgROE8RrbfCLWpixukAQudFsYOCSkYf/2N8aX
N8i2rCu8hzg4I3DOjPSxjQKYZDOXoND5i60kDIpyK4FeQ+F7Amk8TJiy0rrlW4xe
GsVtk+yvTnHUSEe46zwzal4at40G7PjRpe+CZtHEUAVvYJho6SOz2kvTvEjVeGwp
3j2hBqNWO3+0se4ukT62fTRY+yfVnHwsfowQ8UaO0pWqsziyHEHoxjPG1Lh51U0X
MlEdTAflO8uCsYxpJT1pof/f/cGF76Z8NOtru2RZoGP386WjME5WCjqRznQPqM64
1DlTOdgLsCR1SkxnTEbrZlGG/vLJYv7ORizdPEBGSMBqgjg9R/UloQgUcbtqp/ZQ
Teh6O1hE86EittXsMzs6X2gF6qp/zGGGAF+LO6WOh9TkLZ6nRP+0NHPhkHkwCNKx
KHt+AY73RFHMAdqVt4Pq+GluVWjR1umxEVKWXLdr3jFawkY4WjxYO8PGQF0qbDpO
uW45cPpH8K3z3iA+HdE+AoaIBTBHvER+j7CjgE6zI1H/Suj03zhCakwy4+ODM6+8
3E4RrnxqvTq+58T73osKr0YFwIXKsbhOJ7BFAzt7euM5rE8y+xl97WeewY3scAbh
okvC4nV3/0haBA69dL/x2PSM9dSzt6FjkLM6Oqav4RblQInR29aTKAGgokqHauTW
5SFU1/kq2WWMw+V4WuhKfH033lSV9wLynyUOvVLpjP7/M22wLv4cIGuDFbC1O001
TQgiDwGqqUlNnj9T8f2+Ch1J4dUZVW65SE+s0cw57CYBWbdwXRh8riLJOnozNBpi
xLOLx4vwa7Dd5/JtrDGeyLNi8Iq/8a8XNHO/u7fsY9XwqkhupbUxuljUtIuHGaUS
9vCLmodDHpvTvNKJIU1YnSQ6+gofnLYF8yLGSp5CPmEptBDwHPSZEtrcNKQXNTvL
KkyzzjzctiIHOjd9jJRauSgvgV6tVaRXiWxOHpbTuOuF4YQASsSQsCsYIrNjZfcd
bWxdInpX/PxeFGT8dLu1uorJ9RPJWwwKroh463TRQ0bibiq45WT8YTvPsP3cNlO0
lofZ0/Jy0WyBweibGJ6ZOqOoPwfTxiYzXho8b7tuEmG4z81sWCjI6KLyigbZxf4U
wKN5iwxjL46MZOAn+bmEyoJ1vFy6JEQQT2Ej83haGGEmb2Fu+uSBg1r8tnB9nikB
m7il4SJHxpMXjnvY/fPspmEfMgjxjUYMxPjrix6o0/9ZaS/63xvld3rTz0XaWT6U
5L77pOLLdWpD1htsCVNznkTDQazwUjzonELUs29JIcg7Rq3VbgBuKWkQDAmoR3Hy
1mFYh+yKws9Z1JAK0/kH6A/T7gVGzoVohJBD2Z2RogCCCZW7oxgeoklwfuG/wMUL
vBWE7eViNwuKqQzNmtcb/6Cbh0LwV1jkcdxY4OEL0D6oT+RIi9UQxOa9NkCNgmvF
a1bB9KcIp6nq0CzSO1dOClcDjNb4Gb2lLDQ0YTOJ7ihcDp0N8bi5OHTHKHG/vRDb
PbxO7po2mEcPWRgG0+NsZuBREuKAKzQnAQhSBUDR5V4nOlVNd0Rs8FnuJhI9QA+k
gUQnFpc+bJDkV+vIGOcaA812IYSDVs5GAr0V2ISCb/ArDldTgJx584U5ZH19Wtrz
RR/Log2nhWVfDZ6qicymcZx5aN2Lyajm9KtygnrvOIc9cl73ocmqlW1HfJkJgqPW
2vGzyl0WOm011qfBmXfhY74KY+EVcGZcEFo4AiXNvPRPQ3MkhUiTgXoL7v1Z9pZx
QvQDaBtZ1kSnozsjeOnAMGxX9jUOb1W4J6Bic8nmDjYB4HjwILnnZxQmWHlmctbw
AGtr4BMCvP98aZzzk7YgJzbQdkUI+LDaqFvh/sN0mFmIxdQ+WZWwZE8PAV8d5AuE
eD3jIuwxwbU0UGLTI09K6EcTr2zxv5czecNg3k6hvt2f1jSwtV3cqcd57olQv/1C
c+GJg0Hfu073Q5ftM2gkPNGJyPxYg2G9dcDE2g7wDpGRH4E4dAPkuS1DW90DKaBo
heKqlu2/BTkIAuat6syJqY1fgjRWxdLMLZV+jPDy1dUDEBQ3SFmO85LZ4C+Y9zHu
no9H5AQeBPI1JRHZhi8Uudrj/VLC3sD9FAxvfYScPj4VVNtBGXSGfXZuHSrkKk0Y
PEQoaBIhvGrgALi08uuXXuRyOoSJGsq9DnyR00FQO7ABWEPMbG2ueoVeOCuOCl9t
9kDF/kK3s+U4PwJVamtBKJDivjMPGQ7l1qU5jgOdY0W6Y1scwmlb3iARLVSgnJDK
HMKDS/JatMJRJyeEn0qNo7UPxTTF1Q0bsTi7TNShX25YMQ3eKyzxpNT67TdhuU/v
jPQPrE7aPcsGY3q2UElelhF3krGT82d1bizTq8hHyHhYQGgfQXS8dFUNPJviR4LH
778i4vLtMd/EtmidBivdQoAZvil635DlELOD7zg5xQLmcl2G9LVL0WYjF3qfoLql
2zNwN/TQN57YogzABffMLEiNuih2sj8pokYqunSsjdiiIcYOm7ozOtLxXVXGGJ8F
GSlNs/i22v2cQjtmY25Jj6LIXFiJ7Ih2i+fSNgzMNr1fffWatpijy63lbz1ArDtD
16xk73VPqBBNwfqJzyWCXiIdgTdn7Y1+WMFKu8BSE55+kS9bDZPnY/qRp2DAhdt/
C6zd0dVzQFsSTbjVJmSz72EeEtgtgKRMMuiE5EzVthq0OOLa1NZRwNM5dDz5XwQx
6p+TdeQ3dHeMJCtFW9YTrjEaG2+4FFvIwk2F71e1qcZWlPRrMRITSHEjsj96HOrs
d703eKrgijpe5oMH7optxuZ0RcpmSnJi775vZ8VmMWSsZMq7uiaJkX+z9H8HNpCu
X/WJECHWjV8Ribyub+bsKTDY9rKak8qoVi+pbCT5OkbSy2kQdLrMn7NGVJzhlyDK
gr0GrDLqQo26wurbJhYZ6nuV9Y0IsLCMgRTWgLMHDFxxEUY3fAamKdUCGg+YXJfJ
brGmTzJ1w+7hs1xkV1GoeZjH663/bxlMCVik2K7jKQfZbkc0DsEGLq7ScLv0G1ri
IaXnKtVDyM8QP/BBj4Iv7HgsAbW96s6EMEyWBapXu/YUL+Ymqi1gbKhv/6skVpc+
3YEynOmwK5v6zK7Hpz/x+PZ4ahKlze3MPKjoipfcPPiIp18AXB95aPw+VFTadbgi
bnJUb/59QVtZ/7jiwsqXjxlphHgMBOxedsdmktG9GoGXglzCOw+IrQaFlRFMN7Ek
W+RpgGNoSgfuQxv9Aa9dU89hNx5A173VFJyV8F22O+R9CaYKxq5iyPsWrWKuCTE1
qOSKgxBmZONz+iqK6lPQorQtpCvkREjsmmrH6AWvXbVM9uGgY4OmdDZsmk4282Jq
NkBDFX4Rs6b9RsJVEx961CSgtxTkR9MkTfAK8Hh9lrv0c5p1xNOg701zdUG8TN9D
rl99CmOUoA5fi2PlhaM1O0BdO5Nd8kEzkep6FDR4Cgfts/XXSZtuf/YuuXVW/Igw
wNselbjzz3Sh0YMtV9EVr14qzVw12arBvp7ApJe6gRAuwbh1FHy1uubyABgED6PQ
aktfRr7U9+xwhrxdwnuv6GNHYO9/ZxL9klrYpYcu4RlZwokiHdFTUjtwzngup7wB
A2OQFnEEFdxoB/GEle7wX3a/18lvcKAy4g8mYhRD1zQEB1fkXWUaDgwNHB3JlHWi
LcQfi4dyqX1OfRftpoMxhNJovIBZM+64W2LVOXd30CjX0rRP7xkRHQNl89vGgsbk
I3ULx4P6zfpFZDalnUsUGPmhkdqj9lXQWPAqg1LS81T9lWp/Ni5QNMHuuhSx1R1R
lNj4hgzzJfiXs3pkfzzIz2VSQg8etMgxGRiHshMI9fKEzX/ZXJrGH3hHMdMiWgSm
5N743ChXqJNZeCNLfsh8j7RbsY/I2tZlXI6wI7i60EqNGZ089VtZRqheTJDfK7CO
msruSrjGmxyxGDUrIjnyl6u7Dvai1jzQfqJS4KMOlk0Bq/7U36ORqp8JAVV4vnmC
7Xa+SGyyvjz9xTRhj/ybCZExw9T0o7FmTBqdSMleJ4BSAY144XVDrUZw/IrslqrV
LyCuimxIslqpbMpEfitrg942qy8oMkOqjPgcNibt4MSIQgMapq+Rlc1anLswSNHu
m6F06ojhnLcmBRoMM9DX7ED1levsHNrZO7nDMZi8eXB5rE9N7BeF1Ar1zhfcQyld
mJVPRXTbFC6h3BCpQqJQyhtJjTFcyuXy5CT1vyw9AZsn5IwZuPgEW0etJMjaYz+P
/l4IPgZaI2Fcp7nm43Koh0PbuyFjHEn8Bz+2O6bmlZmQdWKPYO6uVmL4B5VkRIoA
L0cqLB15hnV3N5i1feagIRonDIScxJWTzFhsh5KGFtk7Qt6ixpcFJnKjTBZeG9iV
v8mAyPXbOcQmsqY9jKAS2f8X1PT8UvpSHAEy+d8Uk+6PzWP0LUGjpqSvYrQ1Wa7T
nJQaTeWTzUSsfQVcta8gqcPpzPKjDDtmDK3vw4rsjEPPd9NPMHk+Ptsq6HjECs2n
SfvSUIt43O7/aGMuijYdyL18CJwWsjz0g80BA44VGCqYmKNBQ9+tmxaUdzVhh++R
ovQJRHZZDZB38if6nd8IsMFKu00BBetZ1VroGn9m0y+2jisKc2Asy0O50ibBO9Go
Pox0yHbAaX6iEWf/Lb78TxLZKLI/VAeJ2QHnirJ0r+Qs7x5ZRQx51VTdtMb7r+Zd
Kg7O1PHEI0JWI3kX5yYW53NLSWdo67ZshCeFkigszqWViy6UJc670eNPFs6Uw/q1
/rSJdjmJ0mleuW1AFiNBZd9+h/DCKhsAAc/9JlfywRZDSkJBISacrBwwQJ4zhkgK
5fbzo2wKLEbifMBpjUPHL3VRUbwK8fVvZkrHX9fW4pFCI/prgxc0PPaDuigplat+
B0lTebCn5r2Vzkq2LWU17P/ZdRJAP2nQXa5Z5S9/CBh4Nu3J1YxCji6GjFIn40Hp
mF0fnJcO2VRPQpcMjlUMXEWA3iny3Ft9aK88gTg7K5lXfi5u0+GoIKgANB//I+iQ
CRQaJ/cUJQx+yzkyOIbisZBMsrL9WHX2AG28eABkNgDO3mBPaAv8y+uOcS9ZtSb8
hNZ+LVHAuBvEAVSedYZ1GQk9zENvBuDCgbrt6dTw+3ir/45H6WJ0p+KOfs9OSe2h
PfkxAj+a24QePfoBt7MJOwH2SPlveApShQ6ntFTvc8akcS0QzdXgm3iQ03PFx0Da
6rCLwid71790iO3nEf2dj0SlFUKXxsERbDczcq6dje/yo+0iJtxf9HwBbSPnxtyI
IVA40ThrJ5pZTXu8PX6BzAg691Nmylt+XHvpPA3DL2cf5d0+2+0ZbiBEyUSaHofq
ykCRZ73OCtHprtlbTqU3OUaMh3NoH+CTgMDdQBVX62gcRkpvpx4V7nT19ZjFii4z
EYV57joZEsuTzGSNG/BmExoZQ+h5ojWGirObFn5H2te3azvh1f3s3PhaOpxsNqfC
xMFK3vA7y28IiIGzHpdY58LV7qucdOrmYPi/wYxcPmCNxYhqy65NupPlw4IK/wNm
7O4xDlezDo1L9t6RhYr0/gQkT9KGMXoQgrre9SrHMxtPoxXSV6w0+elRHm1sTP1h
yIfYpZ9b7Y/AnDVx26tvcIfnH+roOFkw8IJ6ByshnjtdrCl01sM6Fk/J8PC8xybx
WeiSGwcgwgs4xQ2cjI6vheoaO65t9gY3j+T2MaFIjGEe2lO7lpzS6pb2kjq/Ndg8
C368rR/iZs3WXIpbsOlJP+76G25V+uDl28ODXgpWc3+K7+dApMWvaPMSoFhq/PhS
zAb7B7qL2LiibwSHGM0S1Z8wr8WEScAMxmYgwn4G7GqtIhIWo8YEiR5QJ99CdsrZ
md2CwlSWBH28cXjO7G/Lt/FUaDhH9plnEE80dS7z0HURsDqaCMz1L8nkCIpQ9dwV
yPfzp+2mHGu6oOwk+eFVjkXb3eqzYCZFNNP1QfwmD4wBj1sNUnPgbDecJ7yxMua7
bwv6F45D+9bFtGCFeHIyhjUd+QYADVFWlHBskXHwvc/DyKb6F0df5UzLYWPGUJ+4
LQoW3jyCUpHU2bn6/XgpZIx2Ta5lp12HDHmYS0psZY16upgvs7+BXQnH8nED/NgK
O6LStzCszMwE5/gO+TwOYTgpF7yuQTXTvfy75LVm5mf5CZMrCz6495+5x/YKQ7u+
uQKOETn9h+sq0j2v+e4l1kFJnxgthc9e6mnbUnvGaP3GCA9ctac4nkBMVJYZpb3I
FeBYF1YZw6b9rdEOz4CKKeeapln7iNmcsr3WctloOnx1M2eE1ByLysZitrCEKwkE
dZxD7DyHibWxLgVb4CvFK8/M5eAXes9slXAODM5ract5aow16Ph4ZSqGTy5wFYUM
Leb7GfbuN2I+RnIs76hSrHrMBmyNdi1SkmCCJiJL+LKsb+IQ0WJ1JcuTaoQh1k2/
K/bCyPG0DSFtiydHfppEb7ks2EeK8DWAq3pIdzHJ6+eACxYZeh7fb2gZw+VLlHo3
gYwoQmMuf7sIpiyQV92ohvN6Q4KleUeXMxQfW1m9ZePtOORnc2liEUdmtXw69tZI
I/dcH3pTfcT6HYCDa826WTy7BODBoUFmMVsKji0Ca1sTDIMV1+tRfds8H/XMiUpD
8G//GKxhaUlaDwpEkk+enXwG6GJgpUAOJHgPGIxqzwgzsROuQhBNUanw1IHOi1yY
gpto3PbI0s7mDcgn7lpjkt7+SPBjHcrqm3kgPVKAsP5qTKGr4qGoeE8s5yf+fvPp
ytbkR+1S0DLUW1NIrzc6dVL8J/9heYEkOtfSvtZmdpD1O5wYYFiAFmt5gmKTu3fC
+dAGE1oMPm9a8OimLSglTc1AIgk5HGgWeoapFH8C+dgDsQfM6Dqfv0jrSewatlTH
RhhNaeYFuUApJ0IyFrUG22HhlLbbmhoqN7YfvZeaTqcGcPpIh3HiFlepFxx/eLfx
g9BfxyiwS8yN6S+uQeMUwDmbTAh0mqW+8rigJPpyIYTG69STdRRc355VIoojcrKI
VtCBLUnau319+5CNu+gbsP8qp4jt0hRLQpuRowxjuLccqfsqR9+1OBlWvvntZTFo
TjH74q6SOCVH/PkCGY/aYF/NJuQ0ATlaQFA/BLQWTLOU8q1obIei3ohF5ZaNhy8Z
pp9DIFLoMqSDgyXjnKOJ+7n2/Kix8VW9iiKCsE0j8+FeEoyvEivlN+mCrKg6eXV6
IhF2wIs57E96S2e77Wba0yYLM7tIK1IyP2HeG22WYthfwhgFfeZxuQd+0gz53ubN
GbgXNru8ZCE6aHD1VuOyrU5hgTFlkA4rKaAtL5zmdK/dP74bK9KLU/HZqgCy1gxG
ERqpmLAsA2bCKTOJN+Z4aKA52yd66G64O0F0h7B5C+OBn3HlNjUSUU6K7QvQkTil
+Tllqm3d/RJbpw+li75MHFL5/yHs+6EaGQdAwXm9sSeOZvFRTLqIsBJsnNrnHHms
K4fqyUynWe+yTq2YFwnAd4b7EzftRdnjFkvCGBH7NLhoCAi7/B0scwXn2pD5eLz1
UVp52peWvrRkspKadk1ypqcQgUyMyQpoYK9XHntdK5CTCQX+DdSCtPQg3R7Zcu+2
G06HvlVx3p2v/gpPTpMka3FGeHasCHSmBqjjBt67zYenkPyQ8va2K8Xc454jp55c
xSw2vH9YLZ/0l1suJMqJgcRllu0wmHoPsEc2KJqGYhiVtLLwHEA35H4Hs3QpY3EG
eL7ccPMhOnB94OgEM4w2Xlm6DS1TdEzJm5GRGY11SuN87RrJN+ZmL+KRCROUA0pd
+fH49g+nByAd8aZvQoXcpej3e1tomK5KtYvoQFDsgpZuCYYHczvUAzNWPujY5pAW
4PjZKTxg1h2IYfLGm5BwSu0/IAPG8FAgfPONpQpPQoZRlCjGvWJbLURQxlItgjpY
vzGmFDRKKX38cffvypfe/DpNRP5TqYExpx9FrwZlAgAyhEFu6CHlkNFUoguXHXAR
YU3XVoyAPO7vKv/KX4aLc+AigodsNr5jQNxNFJ2WwVoMmv2pIhEJ24wvsZsFLc0P
dbjc0nctG+CRziD8bacao0AvzBPNAD99KIaqj9SsRFHghUW0BcP8LvRrZBetkvVR
NTgVHEBpvGpEqpa4DkgAL+cE8MDP2d/bpzJ1mz9CA3ThZ1BJnNOHtLElG9EsAcVj
Kb/rM/SOe7OksmlP+EwivUk6ZyKuUmrlwjF1mxOVpyLzCO1LUP5CVubEuQxHmfSH
lxvl9lhXrbI4qXt062rFypmLqgAye/anCSKDK3CIpVEIsx3aS+U3An0pngWUcp6k
+Onlizn5A+QuVRf193gHS2WKpYOmN6Xmxh/2eMzBy17JbkTaNfyGJnamVf1U7TgL
ueJxc9cvFyMXX0ZCHGGqSRnTSZaY3bMD08u+/JWfUfGkUx6KBWUgEuDeQT2MA9m5
EcmzVMvjck/sPiLi518IYXilpxx1EtX5wpY+y95R1c0HRQ/b2xyn9N5/HLanSpuF
LYETFu3/y9smDkaeRfhpafVaT77+/2BvjyCTDmHb91orJgO28LAN2Alp3nyhGODX
VdUYmTfChEPON+YqeVmGxLpUgEnHib+AnMlLteO4tGjZQc1dlCxNTOmlT+Oa61Dk
CnrpnYiaspvy+bJZUIZ0YCsIbayJiQp+l17+F+AgrNzX0Hq/syb1LYY4voemiJaX
l+N8dthm4cakmrsO/fjF8Bchatva0jfWJa4RO8MsLg+ZRr7KVmO6FO/rzF/Uopef
/TYYpGAB+eo1cNod9iIRInRhdu+TRh02iD/WTie4tlRU3wisZoKgZzBN1rVaoqQT
A5XY9SfZl2v4bVqT3VNecI5q7JcNyAdSuW1wu9uoN3hmuCjUv55jwSDp/iIwEmt1
n8tMzd+9odi1QQrGoyyVyZYhSG1xCV0ncQigJmh32MNi5GPm4AUZKzzWK6cDBWRZ
BOwqWa8jt6dQm11WUm8BIfnK6PcXFv+6JQ30sF75LoU/kWrGUw3qRmpZox6McIUp
QYVuqz/q/Cxy9vrADNo2Zh0DWodv4K/CooCUN2Xa1CJ9WcjbKjanK+zs7Y4xyU9h
kmGCr4KC2u0B7iZlpQRuMWzyL5d8iHwNbFcO4XfaNubnCldAC0E3IZHExRyA43a2
AHX4+nNpkvejtyCRy0l8TRCVHJ9VjjV1oWukJBjx3JjNGomBcRjf/BIM/rCxz55B
/P7h4dN5uLkcZb327FmgxpD9HWiBngBvhO8GhpAKXwfHQaxnCastwOk0YS1R/2Wa
XPMRUtWKwABHlDrTJ1zu/yj3QNn5u5wdYy7gOVPy6Bly/AZybB/IxMScuUMBlw+u
6r7KwK+kty+eUlzdSXw+Lp5WK3UhASK9mvf6QholdxdASXTGH+8/J5aeLgCcwwPL
6sHbXdWF42yV68dxl4NhDXnXfcF/wx8Q33ycgIMppMyK/IU4Aaygmr623d+hUWZL
Beh+NT9sKIud1+rDaV0w0V1zN4D4IGyEsVajYoiZIeVF23fM4NGorSWm3ol0ugUE
b+xWwjfr9BO7i2sNXF5mFdv0A8xWkV7J/rcj3CrjFR1IxWHuibY8dnba8h57e53w
etVOr/s5+HNblVtvK9saMRpq1cBl6V3vPcil5w2ObssThtQidYe7xuzzoffdWC9d
bW77Pm+LnVx5qeLUfFvYLgk5T2Qn8yKSpIyCTXL8ov4EADRbnR1IVcVPcy6Ezah/
RFzSa6l9p1keiR14cAvoP+yqAkT0e0u1VSeVKtN2fnYU8KN32GV6x6mazHKDhp2B
gXhY8efXmmGPhhBb/TdCYWlZKx1nUji3ITxTUAFtF9Co0LN5VBYZmeZUsW30XjRL
1SHBqqJ6CpiVX4YpuZGGzpVRloJ9dWN1kX2u0dgQPuhqDiOCIjbeKbeShvTU/rlx
7f/0biDSfUt808ak70+zlY8/h6GAntAeb9a/YP1HCi1C1HOUuY6ReVfUPAUYZY2V
woxl+gnsY49wkdU7k5jsnmSvGqPduk2r5Aav29IUIKfz2qn1INRuypi/j0vyRIT+
ug3zMJNWcmSIxm8epYvU6RhQ4e6Pieu7yD3Ofmk54TYKHIQqH5FR6pMU/qPzyCzk
0+T9Fvlzm34l5eH1ajut8LeLJ6nkDgFozc+VtTV9Mn4jrUztM6+edoBaPAOas0/V
mBycqH0/Tcirx76OniVgOWwImWpwb4nea7AwNOpEy8tK/GPOErd5rdCi0j+wkm0K
QQpYcfqm4o5QkbgajIBJUSMS9kIt53VYnYzr5mgwgSuJEbeJBYLt7aY7FuuOCw+Q
yrSSZ3X8Qt7DH234UFFLBhbyxIPtLe4c/bvT5TJG/GFyZsh250jw+GrsSia3vxmP
IdPUcCWIWqhZMHpYiyb1gBuFkcGufkYtDBqeCgtEkUJ4h63Zn5rBdEByI+Bo8h21
cX4sEaxU9pIhZzp4rh9hy0jRPww51S+YoHoaEcV8VBGZ9BSwvwU1sFUz7ui9dClw
WDFml8wOi8b7fHw3Vfv8CbyWJYnc1BMMrYamoBwzS85rPUVMiZATlz5C7nneH6Kd
G0aT/a6hvAdqPoNwjK38ffcrzM1te/g/QCXESqg5vollgCx8tgCN9QQZ/o/FjzVc
Nvs+xE26aFWKIE3YenPnzeImgnl4QwfGIevNLqci1IBhAjGofSqDPrSKNyoZ/Kqg
H/2vG/RNnmxEVkHzkKlWocycGTGlqMsu2zBD0gep7AssSCk1772/QdyHe9l0nywJ
uCkdyZbaGrRwBTv8fGOkYeZtKawC0o+/LVWIWQY3ae+t1k0WDsQc/BZ4VMG/CTlO
if2U9Mq9Gwfmb0ybsg+HjjoVJueg1R9ST5Ju5GxNrXWMIzy45slrmGfLlQ4Hyrni
rbyf48r90bo8Ui8cW7fc63Kw0hAFwN+icjiZ+kVI0LA3gv8mh8SakMmc8iCKUp4k
A5oie6zgTVidD7L5gjPJqMh+UAP6xeTXT/g7ABPQKf3IWY4TOBugw+x9JesotCuY
3pCV889EGPrcIKvNsas6fpEc6XE3uOOWyZd7zulAJVC+l4H4X274jYDw/a4V/ZMo
vq5QNBjCdfVEOHDYQ1TsAXeFj8rGbXDEKJVqxJGLE3XMH9Fi25+mtQxSzEsDCi53
Pyf237xvXQXY611dy79fF/EQmNf3Knts3BKCgJe5axKVI3cs4LHViQMXsMn3+9TL
dGwuJWerWYkg6hs/0MUYpscJO7V4iAaZvden14QncZXv711welH6Wp75RfEqyh9O
EloquADcEmFsNC+mDkVUUxBJ438sCRNfxTn7WwoGjEBwlBr46aVUC/yPbY7kRyIR
B8Kg5MgTu2ol2XEVuVL1QuI3bi08LpQhr+6jyNOxkSlITJ6lAtDhxqHsAMjJJlmq
N5V7fHPm8BFaIAX1PxNPwVqDOjtlQ63c7E4HpHatKIY9k9uQvgXF9zvmpp9naiUp
hs1+gYGsSZi+bfrpOFsJC2/8dF/jAPP36YsyUNQrH+vBeIVgKXB30n5GE7FJJp1J
sGoevvu1eByMF59MMaY6dnIkVecOd4a6QO5E8vkL4ukIiSPkeDI+EntBxXpEX7pB
UYcaWV5NUFqI95vlnFCPRSjvuu6clhniwg4RzIkyjePoFCx9nHDoG3VL3UIaZvEA
2AOvvdQIWTM0uL3fXmt/ecTQWKGgfRvFziSRhcVfxeJsSnkyl7I3Z7ZU7X3kZM5G
cdoFoPhsXzGoKtywE7+pTExuANOjkGDhpOFKFehKCzOJXEhktFLWCrWbRmwidCe8
KM6rusLaVTL1BCH0DjNMyC/5lpWnhmCC/5A0/3YA4Dowztlo0fieDS/7LmURtBbN
EzLOgyVDJVYlaEXUl4TD5GU47qcivJY919Rez9tIxBNq3AUQjezL3VKGBu78i9c+
gr9R530s2m5xNp97Qz1pHLYHS/rP8saHnOU63p681980yH8t0VYT6iSGBNP4pfcD
ulkvlGQIp8OALronN3AVjmMAZrHHi7XIf5Ba0YB6z0/+GkpocdL6OXmiKWodnYBM
ZrsIYLpbr7KrdCx7K3DdgRXk+zyb4Gy0U+HL7wkvCAeGmkORkRhBTPYpZsOEVohO
lRZzIHHPKDjhjtkPYt5i4KQbOx2mL3OE9HYN7PVVZ+v48q9MxyqgSOJbr5yo20uT
wGeY9byX/d+x4WN3yeVEZPdyaSz4x3W0xax14qhV5B/sBfq1PXTX+yokINptNxPg
Sc65uBGGK9II11xDK1xsjC6N5ucgWXgdYY9UO7Xvlk0PM+WsHm51bdGtO0ITPfye
lEFtU/Z7yZEuY0HfT8nBEgYN8EQJxIRZeB1pb091R8NOyuK8pJozTIZsUSv+sZmA
ZRibYRCjpm+kVEJpWZk5RD0eteE/uzZI2J8NSbdRK3xyHN+x4bJTaYVb0vudMtvP
TvkAHsvJkRRQM1U1Ve5bImPJNRP+o2NbD+AQaOKqUkuJ4yIHtT/UA7T1SBsSW/BQ
tUwMYyG28Cf0w9t/3naqt+gGKh4tAFRT7z0gbQ97v5KMWxRrVwnIQpnV5wOocEg7
3PGYN6E6Cu3iZCMToCFghEG7GGrOJAuFBGzFYqJ7/0vkIHXXgRguu+N/ncuVYjBX
jqLr3Dwfe14p6mHqxCHS8UpDNBtwZsaAJk23ypVUOsegvnip/nP+B0rbx+zj2Xvg
/W0Qg5F629rfq1dG27Wfji4TsXA2GN/igE8hZr2FOYdVaW5qd6TxjC5xjzsCjRVF
EWNC+d1cHBQm33H8SpNmlYIC+vCOuXMA+v5A/bHBi5WJwSKimq03LzYxd2ja7Jm3
JmqWICi8WLi5YgPlE1wXsYxIUUxGPSKZ4z9fTqWVGzRLpWdT+YZ1rZn0sANS6ztB
MQFUb8bU0exK2xVfxve/4H+T5KlGi67FYqoeUBiB2bFAl6Be61oDKWTxJf8tZG7k
z1oCCmvyd4pSu/kYEDy0fWhmXEVfVYtTjeuCo81oafzCB53N95OT/+w8pDhD8AgV
3L4Kxeg+AxEWtzAgWmNYeZLu472AZHu+uhb965Q1cXqDLgSm4QGnWBeV07drM3HG
N3YvE1Lrvh0lZicyhSAbYCIWQ58JMN7Q9J0SklF5psH0P5YYw9QIkGnNsT3BrIe8
NVsv3wKlJFD5MNoiKG63FZNaItD3eA5oM5laQmng8/LEYRJ9vj2IJRLPmMVsjCkQ
AG7JP9cBxMLK0wOWtfN4kC9p7bvPkQKI4WqIx2nTu5I6wBJgUTaMz5qB9AXxOpVS
at/63+Bl6KcB4UJFjgheMpyCSJX5elihiywY3FpH2145QFbiLfrfXdTjAI3hGAeS
rM19bA8G9AIxhDbG6Kd+tOCNn8JJjNohdajWrikIhmOm8Ke3+JWTOzOIY2QwQ7w4
a8hZA9Elee4q88093hqm0EswCkDVLRhaf6rQPU1R0S9I3vmGqAvuRAfQ27PFHO9D
kZxoKQloO84NutCgH8Kctc5yvD4xQx9o0xJN0gATEteEJGDdfGKecjOMr6Boo05G
PMe0Ie1BrY9kd6k0fbLhL+gHAehw/tCR4SNyQAMv/ZOHfY1CH0Mvf5fYjFUrWq0i
QL4pNZIexPgehAXTlyYPSinuRm2SA1eJvJLr3wK2bQPBgoU8KWC06zFAfyTF5Yeh
I+qHE2BN3zQEfL1+qRWQjjZ4PEVv7Q0woJ+L9eqF3Mz4lfxbeiq3HNsqxNFW9g4o
rrU3FQG8+2MPhBik2aT0fhtaB0mk3Jcj/cmLoBMM+S5bfaeL9+t3qxgDZof0T8fI
8GtC1O8TPs0Vc9OOBdB1gx5jpbL2cyEFZxyBdgZOVHoHh++kvsmBb7ki+JMuHo1l
sfr7SU4TkHqnlNuLmgX2T5Nfj2Ka9S184BUZLwRNhmgUSR4sMsq+/PhymYKn5ac5
+Qt+2ogpxH3Tu2D/pSZAw62AjmzT4VkQkCJHisHiYv+UUj8I74v6+2/0F3EnILoX
ft9r9GFcvxnbiLa62ab+MdluiTU14A1AQNgj4EKHXHWRy5Q7a32un+GQ0ufJmb/j
+bm00w79caHpicT3lnK9k+gU6RmU3nw02hsAVw82kYkeIa4RHM1QknbtZlK8v8xb
Vi4q2y5NJHgJB5dEQPdvsL/X6qOOts3cHbYpYgwKRaHOZtj4RgKM3EUUo43sM5xD
7F9IV3myZ0cVUDaWimenjG+5DCh67vbQODMisdtbIx8yf2fCqfCKAfTLXbA6e+ha
Lymb7k9sU1sCP/Z8nLd5TqAaH4J5ooRe2linrEhTIut8XF0tgnX2bXey2b3nPBkp
vX6l5wFzJaDvTDi9ri/8dV9GC/M60kzwqmtGlNGveID6i7ktUayCNqiIXy9SZ43C
u1Bhqy7Ker/8R1XaxjQZ+yH0LUwitWVK3XD6TEweN1c49CN7LFAwQcFy6zT25czw
CrWOWBYq2uxnLXaYiZOoQc7Q3jtp1ZdJQTlH2Cejsdy8kdAbm17UAVHIMr9atdBM
8DImISBSnTyWyPYvzTb/0VuI32ITSswcPFDvHdSBL+k1QfkXWb2qYfiWcv9iMvhh
GU5SdxMfuHU0sCO8egn4mpcrq50KwD/iPD/95yUX3pVAsVfiZsuQslqsn9VkQZRc
MGKz7KAOGtst5JJczijoCZ717BitatXYNy13lGC7IP8RLTsNmNnilDa9wNItNojC
v0YJoeyr8DqgkM26LfoVHBvN1HDMc7L0mR44PqZOLCiKtysheExIYE3Ty+Kmehgk
AsCzxoTRwmSMM/N5KG42lVyakpk1KQk2XwfUp+3ObcdnHBA1FjqmEma7LG3M/sf/
ogRlSS5BERA3egbaVm0mTi2cejp3jIQ0FbGDHjwFJTunUTQm6BWHK7E6YqHLua0T
StzPnbDoMn1iJ/pEvveFLmvsaI1lxi7h3JqosviX2oFey7vwyEcpYUuaO5E4BYE2
2vqEvmAhj5UWbDy6ulJbEUbAnnsUfEehnxS/5unDyU6RwgcuN6YVj+NACr0n91iP
ECqOc0QwuHfqoe7jaE8DXTukjsTxI/bktpcgyGuCBoyjDwITgAm1dmZ0ZDsQbo1p
bnV4Jb3Dq/hdI5G/yaSzLSqjcQfqThhKrJQOh2gp738e2DS6B5+uTwpRbZJUweGB
eHf33fc4iwt4ozRoBdB6pR+HJmekRNa9cUM5klgx5Ah+JoiskUF3ZursV+Bo1LlN
9gpVf9bLMhOf4e8yDOKBojrpPRA3sQ76/kfwS0s6d53sdc/223t8iN7+mSkrXa0N
xhYQe63ooIh/orib4lVOYw9gAcdAi9yg7rkJWFRzB1FCL8sbOBDMov5Upp+oQBuU
b1TYhAe82gQurICAmkze5VDnPDw/ErQcO4nH9ivMmELDBAwo2UHNDIW6aThS/a6Z
qE1iZQPcwCw2OJ/aJeatJphmP15IPnZ/3uztTet0zvBgvJ8SRyLOITrQrxxQCGqb
3H5Tg7kUBEJhELMJauKU2xnBO9cjNJQk+JxDlAVuJyrvgo8C/eLZE0nNbFzmL4RE
1yNbYWTU1z4+aszCKKcEmdH48xmTuKBlXLkSXorJXBwzNr4j36aLZ4VOaeyLwrl+
JfjRNVTDdH8Hht8I1V9sSTrL6YO8zUxULpYyeJAEXBgp9Iq7JHg+yMGanC8zeGNz
1/f5HXqKT1g+WoKi43mACySA1AnL+Gp9ZJ7DBLNxi2xDkqTPOqGSau+FsuCFbN7f
RmxfpR0YTRaLTUjHEZPJrdCIPGjZsHcoHusZQyez5gJx3/WB7FXF5vPc4SQ2naUC
eUPz7dJDhN7ATo1kfal0aKHv62K+2KugUdQZz8sEA16QUZapvJxOoCra9gjtzQ9r
vl5LVTF7CeW4YCBOJf/p/3405fSUjcWyeKkGVn7y8aZO8ri1N3Y5akGOqXw6NqQh
Iv+lp4cSYDMJCipndZ+6NQBjpBv2cCtP/JaFHfNKLyTXaDUZEJmuwIf2k50M2vRk
QBAy7YGVqQACE1WZOBa/kze96+BlnpiXRqyzheANRIn9melUEr13uWifkLdrTYKG
iFg3+VF9WFJtkEQPnf93I51g4NSon4/qtrsmZV8jVx/cPNk8+VzcQ19cla9uy0KX
CSZlSDJaFigpG4SP6iPQmFEWTIIKKou/Mi9eR31JrPbFljscRFwIFuinEasVtqV7
CsZRUsmEFHjXYhaE9KWqiREtSXCet1YqzhPAnVJ2LCoutjImGc2KDnC82mlSgw0B
EcAON22vxjctsOhdGWkhMuIAuSnz7peQwYw3qEAGKx3dlF6MhobTY+Dp0RmYUrMQ
isYJTpsKNTin89OCx4X7Fx5l+JwhnggtsZmwi5dwZWttcpJXNweise5iNlLZDfwS
Oy7PH0iyRzEBbEmLBhis4JMN77g8OnYflXtM0j3vOWRkADFQDjrd0CDDqaZMPWrR
Ho6AH5o1lYT5JbSxaJyHfmDZtLp6LmJuzQDzwcxIYppR4HsGXM0O8E3MmK6eOBW9
e9Gf6yCZf6srlInh4p0jkXPjJwbOJgdPdgEG2M+kvkWUiYNQJ+3+5SLYlLkPsgdv
R5yCibRAjExIojsfWMTa93aLqC2F9Oviy2UtDI7NgaLFcyZWq24LoUW6BE2Ro83o
/kAZbwFvjBsLE0CCVi/wK+7obVVJ42Z3Hr/c+a5FjX5vdt//smTocMwjWOtsz7JO
giq41RqUdihuBINaucAZVRwbgk8PiTrLZSNno8A5Y3NGRhzb7LZbzlEh7mmwpx+W
Q4fIOjbQA0cUrjRuCPMLtm8LjVTS2k2RRyt3uH+fZ41dvCTIX4bLi1pcYfA7+UT0
QMVy1UDIFYYCzXK3QgFo493akEB0FcvKPqjFHxTuNjROGc84lTDT8zkuNqzAzCk7
RsXECsI5kGRhPcgfs2YWvmkuuDEKknqyD2EUXoFcFuu8xXoouh2awJ3JaSCgzD0a
Tk9nP8dbD3n0xz9IjZiHYj0p+wk3FVvgQ0skhSJJm0n1uJWE4EjSyWj+rpX2OeK3
eh6tArPTM3bDJgBlgRP74s+jJ+YMtnrwPVXABmwLDiwZPT5jWetZhydWYPc3qJus
HgZeweU3mqmh0VYR/5Q/1YPZK3jAEnO5m7Itdxq5s82OqyFmlbHDbmPxOsZnBAvR
/WEgkpp6xSnF97F24iuBngKZu/q6oESar8ruMGHNAM1LlFZv3OtkYghcVhvK/s5K
gib89nAv7Z71pzjr63zMlqA5JHvoivLzi3nqRMtrPny+08c7wm4SOGmbWeCC+8L5
qMDoaEE70K+KRmg8NpBry6WOIy2mXGvUWTQ86oP8UnhjvF94QfJsnlL5DvlofiJZ
MQevluvBvWMNS4uJ7TwIwOz6csZSjXW+4mlcXHtbnYhXi7AynuE7JVehPBTLizS4
YZxEhCwHAv4O9Vye/XEC+Rvm0kCB+l8fFcrul+xBblY7UEoeaJtMcdEPbfn8GJIe
RNL1qY6G5eSAVPd3D7VsBnitrdod01HwEqTfLa5Mw49e8kE7927Xm59fnROJXkmS
VrXYn5DmeDWWbxYzfOnNshRqvJl5pxZpkZyI/Hjl/QVNvT+oAcOMwPyBY59HLPi+
SdsJsf8sbwty9QUY+ROg/5yaSC+W5bTTnmsZq5lesmbyl9RZWDh8N3fl7crlBung
XifBLmCwrt+S8gK0/HbF66gT2q+XZ4eaEdojbNFpt+7ZYCZT0tjvYTxntvRQY9Ns
nvin3mHVQQ+Z2SOAvGsG5Z1K0qRwhqHqTzCccQqDrAMOG8UTr5tWtLsTqq5Nb3Vd
AmwbK36rPyOFz4jsDg4K0np3f70+JAkZEh/wmPE142EsClA8+oUsJHxoClY7Fcde
Wyjyw6v9j+d/n2ZkfQwm8k35ovVGxdSl7jG3ywtdNGXMryCGYJnV5HkhvALX9J23
eqzkuQ1XqWYlsJuiRTMnlVR/F1UpL/wKLi6tSl9wX8sYHgyiA4Zee9U/ej0MVR1K
gMWzKH2FMPZg0gU7yOZRmLoA+phD9Lxlzy2PAam5oiDQ7RUrtjZMhsLB3K8EsSEQ
BkeTOYtdY9+O5sfCVOxgKCoVqNK49p1kK3cf34Zm+pK72nS2T9ZHzTJWo6OoH+N8
AYPnk/Fv8zfyCELB8oI6DGhpmutuwYa+GmHX84oHDdqFuSrNQ5ajC0hGiTuUfcI9
xliCiBwoPkEBfiGATgLQd+A+OBpbxVWmO1h6cySwdWdMLDgGm9mj+bnezh4ue9+w
7mSzZ2A1p5CRF6qHBjJ8g1AHGkkZJEAQTeSOrVY9IHuZvSOnpdwCd7lxLlitl5XP
U5YhCRx6pTOkckuE4l8dQmoJmJ9PlN6jefbPRxUXXNHy0t8rb3Yrun36tMlv/jjV
DTvbb9R/TPto7jHgSD0wyOTZDef1XC38BiBT2rJ7EVkg5i5KN3BSvl4hRPUfGRuo
65tN5Xjyp0xTGOEX17MtahlS9VFMSfHDOXGWITcKigHY2/o38G49dncXHeMizwMI
jgbybF8/b/8GxSY2xVzQ8EvTVIDBSFcVDh9wV6qUl93RrCAuXXrU9RRQz+6/eK2d
IGdf/w+yXAf4k4VAB0P3CBvtLiNw10Hz66A4HRQnbTLdhlenhUZgFDDfbUhwRyBl
aMbBvXHSYEVsV/2tsfB+qtYhXdNwCevugJD7o+HNHdlnK8jT5rsLxLDa9hmefcKc
ZifxdQaiVRWima0DV5Yh8bucp2jzaoqkTFTNq8PhBgzODmgNC03dc65yPdo434pM
chYXI2BGhdSfnEpHo4XQ15ZBf3HzqgcpFpiPB4jGc2tYZ5niwZEAzRPR8YIKZJaF
r6Ve/k8fCNYRLh6+DCBqvCFCAabhyDasiTqQ0LaIG61HM2bb6Su1Fg9fA9mW5vAu
zDVi0ryJU4RrYxJ3mmfudSmyfk+ZXgGt35FaNbuLQEmi2mkxPlWNabLxd+rkHtsI
SLlqVbF8Ek4LfTJoWMdPyWyv/fEjn8SMJWccJBFVIX/hXdU9rSUPTiOREFTExu0D
SeG0iOQFM1dZPCB7iMNu9f3ZgZ2F961FpXt9IXaf9BOfmq3Pvt58wza3FWf01sC5
ESx1aPR/jwV8UQCNxMqh2mPUTtmxYlyUEe1u0R44FyunSvUXWOna1lkgjz31TbFH
OrjnZymgzvC/uQ5o5pPrKmoylZlodpeO1UFfOCZ4iwi1nBnm932X2xW0XqBoSoS4
w+6yhZXxAu0JP0rjEE7icpKTb7QY0NMBWCjKoG9NaGh0LxWGUesbB6YAdZAd21ZL
3U9qhUR2/pAVZ4etfLs5y3eMzNwNIumwVNytfK1yE2yBfCe6BZa4B/+8EJ8goz97
A9adhNx8Ec12PD4iH3WdNgQLydkbW+NP2iLi5dzA4j3QfUtzjp54sRt5j3faPqKX
jdDTXwdoZ64jUcVUlX2RBXar0NanTlJJVKK95quFquIECRUy2GG8Pp+kaV8yDg7A
Y/rXkHUgnO07JwrWom7GGLOYDTz/EA2rsz9SqgBxfwzqyAglklyEcEwOI21jKRSz
UIr1lCb/BmbfhXyVMCUEGhKOqxnmNUeFeyRTEodbCo3bf8MmlTMjDoZit6fYXbLZ
tZEJczcioIzIpe/bcgzzv1M71iTgVwf7P7UB8hnxcL+AZXvNtwIDOjwwjXBJ0pzo
lpmzx7VAsj0/0IX9HZcaUTc03VtbkJdkYs8nXJf5TWxG9KtXUnnrHPKz7tZbd16B
8iEasssBOUA8eQO5xDa2PjK3UEGmLDHGZaMWfBiwPjkzJTTaM1pkFkmc13IPynqw
qk8amf2Al38yeMw3afsKDYE0xmSaqXotzcjrqzEjlb4gjb5lU6W+0RqhYeXrZfLt
kwjRwJh2ylFW9SSbFRqx+HLHWLYHwIlhtLaXoEx+OdirE5+/PMcD2/xYR+SltFoI
Sg9Srt1VUy4N/ISyEJQYtkG8GO3Cb82xXU1Jbk9ygQVuHzHT0rmYDJIjNmtM6ffi
UQVlF5jhgHh8q5hzRB6q9JUoFW+VzXp3w5dpV4UPi4CEvl5lBL5Oar8wYkm9pmvc
vP8QuDJspQqcYbILGipmyDXF8YYtJyrs7ZvGhhNm23oTog1qdTvj4yQF2asF/kdf
54hr9xvpS7xHAPmMbU8i21VX3R4qs5C0dDaut3XytZUNiBqqpN7/jTxzxCqUU+/Z
7FDf4ekRAdhrMjxy/O+NytuhByN9F1I9opFtVL2cVYzaORGuWqhMWr0VRtQzmZ6T
w6sqzaz/P645nOz4erE3P5pHFvl6FnVmnVtIID3/2fT/zB/mKKkSNqEeTa4hiI7U
lQsZBnRgcq+C9tmkSt7SaKk26odekNjJRwBwxjAmpsYH8d2LqywmIvaNkRkN/KiX
FGPNAaqa+8hsqWgrFosoug==
`pragma protect end_protected
