// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:39:03 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
etGVLstVr7CgpVd63cJZ02i6+DMEtO5kLw8pTFDpeyxiCrPsEi9+nycTGOEKSiwm
Tx3FQJT0rIzprlwKA4yOPkG0xjiiX9PGI6Fkj+N3fFZ3Y+bKc1Ww9SApp4QltvHw
pNt9AG0lLV2a5cPkKCfrHoklF4DJbDYNERFDoxWZPc0=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 15408)
zdG9/o/+/Qwd7D0s05EhCARvwpUrv4wfqnQXf5DnXCmcZkmyG+Y7Yd2vEY6ubSsT
xcw0xEUPJR3X95wh2hzNFV4OB3/L1NxSD0rzB3ba/d/syKF1Nj6CQPQOa57UaQNn
VzRev3sDbs8NsYzJjPBtjAl4lMqxRcRKnCXAvqCwz1qzlgfbIWC1rmmJc29HLTX4
eZaPCuVPZhDvojYh3u8ElxbwOzWHuXYBL3Z1tfUCpEoClGim9XH87g1oRLr0Fp+4
jm1s47pm/B1yZWmCbkpwvCSGD++j6iuHR0o1faCQYGf5XeUh+TplqFTDCid/BQIN
MqaKMNXMnJeRliyPp/nK15EaQm9sNZVJUYpuYePYxpu1NRiYo0yeg4ZM96aU+47I
ARTOX9eq6Dai4tOetWRnZ/VRqgVWf5Ks71yKcTu/QbGzL9dafwZIJyLwsKM3Cz5Q
0pDF3ndcT2Xk/974N6P+TIZifZ5WpZvY6Y7lcpchNRSX+1I1x7r0xOv4BQvxvsKR
8OQoiafRgyGseXjyzqLXMXCYv+uWRWRGg/T87xmHTnUwHr60Ri+FJFGyg2oj/OZ7
LnY5E5+swauMjiB3FxXC9ti3i9knNXgMEaQsl3Ay9e6LPLesZ1jMkBtBgTlPXYoc
4bH7mZP9Db7OfEiXYQvxxpd/WeCMfrlHP2m4XKhfYK17t5/oaItMgkVeOKkrZkQ+
FC+drTswIfIKjFCvZQYnSegp1BoDpwkXCRksvw+0b1isevOKy+AEkwht5Cj372Bd
kjgjHORsHes4g69oAjCzXtApnLwAjzctwKAIRGZM7Q7t+s/z4EPHwscAgUif6kYQ
KjWVumgslJcCerdNBte69sAoUf7ETU8qf7paCY9Zea67+UimQvjRbz9X9KfRSfx4
Nny+7lbAbYoioWtccYm+GBlPx5PtzwMG/+iQ5U9Zaxa1RzER0nffW3uY/F1pJFpj
UohO1E4TwgHoWQnYusNAUq1UMV+Fk3pzhSnWb5v2uyU0GijlC7+/M11NJFtu72yV
ybwuRJvtWBYJKKip4TTkxPwb2/0ejznirceruJGKCCHhRxN23z9WP5STNhasLUc/
uyn7obF/UzWdYdFBn+Fqb5X7L8auoUdQOEpe9CGxM9BHFWE7MaV5RLaPsLG7Ky2E
0ry0e43rVamwU7dJCN2BTN4RdDsaMXE2m6kRP/OqZ4SURyWqq/LipmkHtlVgB6dH
F+hig8muEvpEfBXzBj29nK13JtXoEDxsknlpsqIPYafiwwXLFC4zQzsRmWZl9kro
WN08TTqr8PPASfCmAi8hMiPhHteaC1G7QMzo20Wk6z61A7t+X4Uk+S181wSj+i9d
YNVbl8l+THRQpxJw4s37Mc8EkEaQ+bc4ScL5jD7bXpjhkEhhEIZTt6pe+K6di0wQ
9L+GKJGf1tu2oK2BT3qzpv6xRnxO4Rrh2P6l0WmEU6W/5oZqmjkObHc+pPIQEvGw
cDsLXT07+YkXowYkwZ8bUu1l6VpzpYCAkyp56P/4bZXbNq4tAStVMC3T/JOPRiB3
J3DxINjlVRxCpN5D9eM6QX+ZM1gKZMRL0PodAsiZfrcRommlAbJt5199/YxlRP19
oOP635FA9CgFNCP45MlaIsEOUKgptUqb+vv6zG7DpJcugKLw4bW3wQdkk5p3VLch
d1JyPwjFq9Z9XzYwTIarBgZ+ZpKCrP/vjuIxtF2v2tS43uHiFw5xtmiuoCnnplsS
3uurlSOyC3Rl7Y1O5EkXWf+JHv3T4GyeaD8h+/0VJLgofFsh9MRn4KcVKHNn+7VJ
JvqgKnnceOoterlM22CccOC76HdNL6kSEN+qOsXWIcCrEpmSoKayvitHb9Jp2LQ2
43H7k20E88I/oQTcUVtLRqmi+Q+JSraJAdF/xBa6uKKnCtSOG0DKBVu/Q2aZllJ2
bACwwvcIKsl3WgSA8E34BXH6CS2Hc9UV4caqrfuZCFfobiCsiwGGFafjFQo0UCnb
dCkE5WwwuiWVq2nIglGTGkuDmbPo+S6zhTjzYG+wLG0WP0BDcUSCzkNd6iuIVsPM
4hI/ubliExj8pKSjY60knkO+WRsYqIiZaR/HzAAw1xOYcMR8qGWQQTsWSDr9oLIW
z7UvdtFQ8Q3Y66MMh7dI8zpMhjra2mhXF4+j9ZegrhN2wEQD8uvjP4jHzJFXW73c
e2f5EzuUgal4dzfpnX8/AEf5/tUzCXqRonCxzQYASqkwhErcqP8PHFO1A6rwjiuo
RX+v76UMzSspzxJWzXr7SQJPaZQK2KLXRINiJaCzSTiemwY+ZNJNsTzb4jcvZCHR
T+om5JYphtx4eHqlY8SzUrCz78F60q1MTlyQtyvf7ySG6MnfdYgjPL5HVkYotAoZ
uf34gu3vsv3R9aI7KMShwvKus4UJKqQFz4MJLdBOIqiPO5QQLmf4lTZNnfkREjLI
NTN+JsNFT9A9SOBRWlHawTRNTbUgAOkTkzOEgZAQr+nhFQYcpQ4+6Azcr5fFY4JH
eEd0yzPw1kvGrOrere2awLolJJxl5dJqUwHnXwDume+ZFP/S0U/oMwO5g68IfMKM
2NpN0wCAZ0jaG8X1gXUvSmOwQ2NRHbTiNHtolwVViukDGT3A9RwfbCSaafITMxYv
pTsV+lggUn9Fmk+t0xgG+UGs3FMk43zIwXhLGQbEGH1/jofMjxtO+9l4gknh46Tw
PhTAiHkJxcgmT2+YmAy3Cu7sk9wMj46jx/xvYI5skpqPgKPtqJgqLMf+TBMiWvbT
NOd+mhyODX/sLBx+iNM0ckf+n4shdTF2QHVWOZuRimiWsjiAaDAeRmA6wz5aDIXI
i1TPOyt24AZ5bkKYj3IW3HXuDRdwSNQT9EMhfr/K1SE33QUl7+d5tf/8BrK1ddBP
l4Wpml0ovfA7AL/BFFMjzrSsVwWM8Urk+68R2S9rlYEbDJKH/g2ruoaSIsyGTLk+
lhtVTAmKCKHaSTP20mWMFwD3wC92vMn86DiVR4jzSLeL2o66BwAHBJXdGHFMMs81
jYAFMZVQVGh1cfTYWq4Bnx3gJdEn0Sf7weuiDmW4lsmwTS21whJL2HtBx85HRluo
L4VUIZblXKvh+Kozir2AfDK/8YqMbnCnKhC+PTuh+8E8YwI1QglpNkcsUbQFkTpD
G+IKgfds7zEUqdBoYusXH7NKbuJrbGBbmhdEQUf1Ug15Qj6Obprwr4p3DMdlAt+Q
dOu8YH/SMX+Q01Eom308/2GHFCKdT9+Wfpzh5JEA/c/OsscNTKSpYwwArUbJd8jx
ml0cJFSkHZNMeFm2hsrBB4e7XP/ZoYS34o9Oqjwu4Bn1iy80Fc4/Z1blPPd3PRUg
cS7adOxfBy1In1dERw6GwHuJjTsh6KIOAu+u3iuXDqV6KKWknne8o3RIepDc+tRN
75Zd1oOdpG+qqOdsL+gK3ZIdm0IKC9KoeN0Y3XW4IyX69oad4VbmWd/yuFSrF7PN
7q0t/mZm+6IutM52c1H2VhvKez+rInXbgeu+zU70iaH+JabVdKuVsbcZWfpNtU0M
ZkcM+R9OMG+/zUfUiyyoCyjCY3DVUxaumC76K4kNQvguhCRFccuR1UKOud8viQWe
5h3bUSq5W38zLx4+3TT9V5f+6BA+b0xhLNi+++vfn8XiZ/cMWzMmoKxiF3soHtgy
J9PLYOSEWlodONi8qZtnTzHOCPMsgRwEZLczXGFF/jjgjXIdqsaGJa8KaMeFoCNR
oOOnb5HuHcVdNQE3r5TdmOA9bx3jiu5xxUmvwzkouxtiyaC0ZprW8IhmsznuLQ9R
4otFYYeL1Xfrpnmfm515uyvzgCxSuFgiWvEqrK/orJ7BpuvaToWF2+SOxyJ1Kp8p
JjxGYeXiQ+ENZ9cvHDhmsQIAWJcRkYxjuXWIP6spJHSysvJ3U/YdOcCn6v0nsV41
KvbSeKrNXIOZSHUT7B/bqVhPQE+mTAtvbMbRz+XqSZ2I0S6Npew+vW/3WR3ehlDU
dIFIwqmChrEUxJTAzCt7LEQnvaXk1+t7DgpiKVwB1Fylo+fTb6R4GwNxOdoR8xDK
gZYl/vWRputtkSQyuhpa9oyJk0QbqJ8AiqiC6FnuC9w9ayJ5PdKCEwszeUXc/NdL
XV8+0342pckRLO1cgeGmK31ztt5P9DbPS+FKHPGuzG1C6bH+anayCUpLg/XWg5UG
/N2tZxVTAS4gVkqlB3Oyg8II+pBXq6fRhgSLjOQx4SQoNM1LenaH18S79bi4M/HD
25kmhpecLB+lXkcn3KKgqbPSQBAix5paUkay9IQBMO1I0q3VY6IAlv47PF5gNIco
DGOGt+ikDATATnVBwBMA3fbB3mX8oO5Yk0xK1WIcx30cDfKHjOmwGQWOlwdi1U5J
pumyevpcMSp3ptmDuEU0ijGM8lTYpixqXGx6MZLnYzFnpNPLRdoz9Dh9RCpyAa8u
3Ez2bmOgZ7EVwEqowPUi/6s+MBALhtZVWJq0hAgoGNuQrJnydV0NKXrVUkBWckGA
fx2DhkK8swgbgeqb1oorz2vRIs6+PdbpFEEU2ecs5sckDr+cCf92pqlk1V/+PzaQ
+U0klerXFQGWguo9roFA5ZhchlslkabmRqm0gUpNK989vwylbXI4eTMkKWCqO7s6
E+SRyhuiW7mrw67pP3wfCtDEuF4dOEK65AEL7np55+3wyQjD3ShQ4GicT6bo+DDe
kRjd9FChhFZjpZJFZEEGiq33U7hnppZv8J9O5j9A2E8oTlIOOOZpSChQFsrj+GK7
QFe3/Qom3XbTm7sLVPGXveiQ0KCAxsJO5fEZFdzwhh6yjmMBAsHP7zgvSTKuUkkl
Gv31eVPvw/fX++SsTbOf77bYwp6yKSp0aPOpaJvpSIA12Dy4OcT733gEMcFY8s0i
2ZY31/iR2rZkh25LKL86dIm5Epo2nJHem3F0zChGDHaW48UjBPxctRHBCmol819I
dMkuzZ+R6l4buFgZKVnvvdlPYO+OC5K77us6K1R/cJiheQ+d/n1KplTIfLO2fI1h
xViuQkddTc4CPFTl1qxsNbb1UNGF0AjwQ7S4pHHLyUHc7B20zcDpgLkBW4OxxDyz
dM0hbHMworqj/Ik+rNmueFUYsRAUPDLhJ7E9N1+AlA4QW6KQDowYRh30QCwILBTR
r1D+JKRC9osSjFyA0ghfxJK2+dGwGTHx1dorkq8+lzmM7bXc31QVHAyuW7B9eN14
YYxVMOr7nfr0Am3OzAJvmZQjQSlQwF+vs01HDR2f/1pel+9/VsVViawY/ihKJ6JV
nHIxmPu3RdHgp98oFqcuTxRbdA9dnFdp79afvS2HNYKHpXI4iS3T3/j/8AqdtGJz
cyrbYmEXf3EdOGKvzZj9q4mnHJO6Df88PkADW9djSvU94PDeyzurk4G1m7CB5wol
TmzSSg4Ej8RJl5WnPtdjxRz2GNN3Z5xCwzRtOrrm7fPDuuALVLpyCxF3PGmUQg8h
u1kjTBcCuzimNoHN9rBcbt5KAnFFsQsI11ore8EAamBXhr+5HD1CajDro9rPiXp4
HQp3qJ0IMtmnIG13RZdQYssN29HwR5Gi0oKPlKGYKno1TUP7OLAuVncpd3py+AU7
uUxd5T2BI5ymXyfCB1RAX2ea7HzG4PGoIMODICCUHp1ki1NLa9Zws1yz+LO3b5qS
QCr+GhapeckHTgt/cx8ycSWV1x3ypzCppY6UN9+y9qzWsbtY7MIHLx9ofQSNHiB8
Og7JgMm7LQptnskbZlvpsuSNAQ1vK1bw0PPaggwWJE2FmbNpisEyAP5gHi9hZl4c
3dLEBTcRMdHhnfnlps/2tqBMQYvxtaHnpKbHXpyRqCvVWdyCKe4wvjDSycFvB2H+
9mxWGKP1fGGpyBfCLABa+uS+W7BZYiqo/2n6B8UhxWD+DyOZtE8BEzudkonzht+M
2SYzydaCFZMMkJSvrauq8zLVpQdLe+aMpt5peF6uxoxySAp0T5f/eK8xbxegWdpc
9huggm/DrgNyFQqIU3zkwllfUBrn1TDt8wKhhwKb/J7RDpmq32a5sHlQsz733xok
9ZTWhLX5J8cqNWaLRQLwiUyiEr7ELnEMpRsD58UeBGvP574l9H+uMTcpCMoRcU4Q
aVAIuhfCoxLkNZ6V3aBWP3rGlHA/UDuPiUmkKNTCfAjVZnPiFOaQajDuh5FsFeg/
JJRR6RJ+5puUQAPDIYLhKNYfs+K59bzEUE1OiI1VD5mJ7+XyUcpwq/5mAvnfKiws
/aOGM5ZtYqzAXSiwCKnhV3TNZgN//6NpwEwjRHkalVlU24jjOWL0FUCq0JvcuaOG
N1BYouNVMIbb1oWZG6boFyssgxo1xXp+AFyWAxr5VU+FB08TQ7ywMnc5bw5WMej5
mrcQp2cadEsSbWAlPqD7DlMC9zIddR888Fme3Yb5T+JTVp0m3HINAR0mMnJDdi75
dOAzt5YfseLqy2l8qwjHPrr8F3HMen5yrqCgDrFguwnsLvgv2Ix2ovMJNPPQQ/ao
iVoYM7j6Yj5R8wti3WzE7KomkCD2AeTAFeNLmpnPS65jyMZRkBv2BGadY391w0Z2
TYJoNwxoNtkQA8bDSds4QyjgbyA1EkwyuyfDeeJBZPYKrSwCUDTDCz+h/670xO/Z
MsNlChZ707IRsS8SX+oTaf94Md83BG+BUDSpZ8W50zgVY5zyXdRS2SV70SR3nH9T
Rw/nTxgSNofBUBHqOK8NLIjHkzR0KlQNz5BASI20uwqFCq198y2tHhMdPXZCRNA8
HV4qNt60W8WLkgYJA1KcdpE9cUfzoSNQNZZzhaNIaBLL8o1bTJrPsHd0qfzWAviJ
RTk4T/ksaLJ5pf0ZPQu8QUttspDxZhhc+yVwnqdkELQCw4LLj6auPJ8eX6crPj0B
Slj2DuaIpOR3hzky5pel/+h2p50T55PARai0agjsMTtADuqenX+8pwYd2bahd+P+
TuMJXn7boVx7HRjuWGyP2XasvCpfC9MGox0xRbSy2gteFpEWpNjw1v/GWU/HXXGe
xUDTSGL/uVbguyeBtTi1P2ErBgBp3ADIU2Fy0UEU6NKfKTLZcTNIDmqlVAQUqOt+
pua1tInajPUTURV4+cCMIlXz5XxZiMu7wxP33E8D4v7XDpt1iowEIBELSwBRJNJI
rgxjU/ZNxzlENP0tsl3NXjwDw58tIKhNpF2uVPCMynJk+gcX6y6djRz4SU6hj68o
1xEF/Hy6oxJdHxj+y1/AcUCXQLrlSSMxH39uRW2WxjmTTn5r008FlC9X3PLhxM8x
OW/VoElXhKKlzC6ai03tjsyor0BJI79pO4Djs3riu2wgm+h9LGUPSL58hZUMfWbJ
fgSAlSUAR2RDolGnkrs4cCxpq0GGOvL4tp4m9Z1KnZhKeaGFKJciyFF8JUSigDeq
tPB03rmupHjhiqNOG5pAPVH6YZlZ2WH7DNntWI8F3JQ/nGUjMvFaNqPL3zKJ7dMt
++Kdbd0P2ZBF1Rhi8I8IV9agf46kp4GUlXfvKHn0TjpQ+jYsiBYw9qxSJfMX98/Y
CtXlvX8U5vDYbaRX9rdbKTfSYLkbLQoDcRiyoit2hoYiEFsDO6BOra5pj3PjAN6X
rb9OYDf+nkTc0u4C5kPOAxHJQyaGEPuHsp+kBDa94UuHDfD9gr32sdT9UaXRW9Ir
Q81pi7HlETDuLG1OTJmcZaGIfZ75xDzYFGXqUyrfA5onL6QBa9GZIz8PWLMJrlxk
MNJjEUBCvamWqd1jJ+fTONcjnYPIfBQnf72jd2F3NFNyIptU+t4bz0trgyKs1x7v
3cR0ObVY54bUHGopv042MoH/R20REAi+Mmsdiyb6nOxhoWoowz0tjonq0/UD9yE+
bC9gctessKWEvenKkCXhQnZs6gUxuzAqLibTfouYFalVBMqi28tg3jRgMcXOhjAa
9hn/KyRM5/glSWdZ/BhRcNi3Tf6OnhFlrWRFFqrK+GEgVEzjE5Qb8bGVyftUC0M2
EAxSqbqwtuexbqPqOdRgW0+zc/EpNPGhyuM6agNDKYoVJtLoWSc3Kfs2mzOFZlG8
IgyT5iVPMxez0whJwsG+s/0UZbefrMY0GyF7zuiYrtbcunFxTWs1MEbRsMiB5MAQ
94itdnvb1qfB2plXR8WFj9FHLjXZIUvRSdbCs2AYBTE/vXVJDKQlVLy09AUyF8N3
gLnKPIdy1AmFToA9cjCCV7HJGsTssTTM8Ki8fvhd9E6PgyDKJ+bi6ZtrGz4UiidF
HjkahqmoEGBikYXpLMlWRJsMvPZVc3VzCnHlZmz9K+Qmn5BIWLqTiDebzEcnd0rW
o58Z8GNdsr9tcApvbBH5HvhjtvSwYQLi4K8d5D5c3LGWiyFUF305JDrJQ5R+y3Qj
YFvd92gBtWAgBNd3TrlFLPiAJYsy14BPyj1lWVPhkvaF3cmKbaZ0L+XlcQ9N73j8
kY0sooU3zbDXlFH8T3G3bf7usl8wTbjdqEnrLGcgNnGgy/Q+yPSqtr7gWBYPEyOC
4I7pT1r/UHOXeAqx0glzQ3+xq4oaEScMemn+dAiqDMCFMnsqDTyKPAJPs7EIKvv8
+AnYOXaObSGZCIotok86jSz+wkEvE7+p4nOYzVV6brdLhvhX00O1myw3SST4kOTE
g8xh3zIWYP3NsDCrkgUX45wFIx0rBNzfX2sEVo5fDj3xoELibOpxRtuwx/3SfpKw
tKLsStZysAscMeGNZdgXEfwn/gk9A/uXH8iqJsQNbVyJZTBu4OJj2c30lwkr4ob2
Cc0eM7Rm/536kqO0D2DIzXGkW42e0YnuWHSP755lQ5NH7apTdSwt6bUifAJn/CAe
slC2nkBKMSbG6nk4SoEjEgI/dL2USHEid2aHy4pm3URlYIFNu+SzBkUshl10mwer
PoRcI4MXCIFEmokfT4mwoU8PIfsg/07qFtORreeQUYPUjOdfO1Ne8kmOxU4xV9PN
3Z+Vj91TTGeTUcJWythqZGGKtNZqv7K2RXHJVRn2LNRSjg+wkNB3UUH6SUqqAG2h
VQSYHOWVVorVWd/wPpJQUqUluHtmG+oYbrFJINaTXjpyzM18RRZefJzD86I6MN/X
lR+4zkixShsnA1SsyJs0Kkq9o2zyHlNCAnaMB9/lB4EOAJ/SvBBq3q4WHCF9c/k8
N29lAIFBETV/2ZlnsY3QrM6TNicY9tbdtU8tKGKZE8AsTy97fX+Nso+5zMIxDhwT
qTz37OtxlVxxM/j/FEFSb5gRM89Y6B4rfSavXFt/cvbSRZ6fVmmwWkxDDQGRWyMw
LJ+ETNgkQjcFqMa1/dJHo0WqVm0X3neG1Cw5KORr2P4VTGzqT1S3hHM20hitlUR8
N/Gg6dX0dF4oFX7ViSVQ1qdfDZ7uHLK2MQBh0S64E62YVCUjoyn/rvTNbhI5mqrm
DVzZJABkHSGXnk/0iK86FQ5yMmsEsjNDHPekwx/0oGcMHLi561b/VB6HNXwcTt3Z
ZKoNt5JZ7k1jJtVFzucxfa02P8ygR8DLUHz5CcOkbGxdoXdZu4UCK3NrO51TF7Jh
dduPXBECGOQv5eTypXI1iwLu/g5o73XRpvPtF+nDCR5vrm3gg+LAuFl1kYGR5eMs
5xRg7sOzhal3mplo9/P2RcDgN/aUANlnqsdNkOGDUg8u9bP2dsNb15IRBPbKr7go
jgxRK273HWLSvl9+zC/okafKs9wLqt72Azf+Hd+tADIgwGhshyWn69fUa03fOnnZ
FiZMo12zDaKpas9DmqvX1r00aNyVVaBQKXFmF2c4ObGGlXdVaXV86NyYFdaMlxLN
5oN65w882EzDH726az9P+B1JiJkY6rklhv46FSy39luBC8FKhZVjQw6smsB1Canh
f1D+RG3Kfyb2QGnnhJ4tItbs5/s+hAXXqZjlvyDdXVWTL6VLiA8fiHsA4SmZO0dG
erCBCq477xr1d3ndn5z7TKUSUuvJDrr63SqOEgOsvwyRQPG+ZAgoQK+LHlw5glGG
bNFvFTvmowXfSfqIxWcUHc3dAwCDg+U2L52Elm6m9P1ju9ujW3JRNFooCbhgZCrV
+g3joR24tWfhEZxVviokoHZJ6sYxYDQcJtsVy8urdWWNkU8n+qFE6L4lzzIkc7LY
yJrhqb3wb7ZoMh+3K6d9qR4v54f6ecnfh/uXhJSn3XlUd8z/VMxwQ9Bj1b+Ut7hP
M4jnI+ClEYhovFITUNbkW7fUkf+KrM2zjc3j8qlKmmnwzhWt3tYeB0MBf+kLDTqJ
JpHSzMSG9Te2AhVuw6HBs+mlgOeOOAfu6adAe3XWjh3hCoQbCiI/i4sBzoVaPNJc
ZfR9i1eBWZG8p2maVYKZgyMnzSEjCKcjNodaDZ+FgIr9bfas0BCJ7t+tO261R2Jh
AYF8C85lNrRqoBcW78JSzdiMpslW4kblK5VBJUgkf3CRatp+ydHo6WOutEnU7yPI
1MYltwgd+ECeb9qxw5ZZ397YepU14zbLm6CvVAVGkUj4xVcH9zaBtCIx5lsNaB+g
HqUBQY5oizwacoJxNo+rtFnglaqweR1YlrVj9HKrv7eCYng8VlgsDdSz0twJNlPx
SHDtHbJ6Babi5plSFDunAI2RtTGvWNohRwc11BhRSg0UjoA+bdF+BB6Yk3HP8Hof
Egky+wuHUY9b1RJ43LU8lrxt/Q9emVWL1+PWmOo9RX/Ju0TnldrTqPeJfw+18mPj
Tw3GZs2ngwQx+KRBmQBcdUB0rXo93rA1DpMFEtPVhS4grbyahAdIilCysqEsxY2X
7vwm9VgYAs0la13gFqGkTE9ddij5cbpgavghw/+pFbEtk6MB9v/KQDVwJBPQLwYl
BroXyP2IQm497991CnPx6REcBr7W5uX1x2/iQkW22VkBRlEHua198slak9HySy9V
rGny4hMGu38Qs7Vien+hmPWihTuQlOwAd1CG08K6HBIbIBb8TGkJEFP9rxa9gPwe
PKaB8nysgYpvVrezoIwq+jEI6q5LXS6zUa9FsL9qcSfRFiVzXEtXGLOTSTjbAF+8
aDxfU3Yv+B7T6RcDeV/ZnMWowoJrWpdZFWLVyEjjE8jnNR1E6uetqOl4Xwts+TmX
/dCA//XdMIUYPuhqqkf/khBBAq6KHu+j15uBt+9MoC9XbvyGvIvRAUpaVCybQlIX
vjWCm53BeSL4gA76ViRmayCWl/1nT3IdYkOS7pt0ymZr9IBsr/cRVgfK2zA271VV
nBHrKmxa81xsL2HY1992LrTf/m+Ha8CqjCBKnmCWqENZ2UHB2l6SPUAuMeuUJVXL
pZ/5tIBDvbQNZvWKlhH0cMXidSRp72Cr9op/UEGoE4QdMeNt8JeWRCXc725weGOa
CumAdOCNZ+pq+Ad2dB6nbwmk3wh6jL8H4/6xnKmZZc5/AKuend6A2Ew2gRagurvu
aLyqiT1cAdq68BvziKryN+lJFW5zpmFZ7ySPZ0ZAmcjPdyv8x/ldkeHs8/QcYBKR
sm8gb/AQCE5d4Qba7Sil1Dvq0EaYqPbiSpzwwtM2fX+GTRkW+8pmpn0S1GbTtvKn
PclbDpsJz2u7oTdL1LfF5Y+aIXZ+BnWnj7GgnQlo+gLZgCYUtiiSliURVVuvQhbj
uJIoHNwJvIru/UThHvUNVWFW0kMVd7Kf7ak7d3Lxnvscxd/uOZSfgZAoGnxbk5Sh
ut+sP72Wv4j2tB3g6443bG1vI+WxnsuvvR0qeJPPBjIypi2UsKCQBV8tPyG2SoHo
PgLSb7WqqJO8mD3g5nwrOErYHbhvmdX87A37AjyMnQ8dilzbwJc6R2/dhCdfN7ha
N/y/kgwiB+A792Ih2yiCHBKgKdwwZALEvhU4/b6dbpUrqVhFPwI28SZxLHxVSeS/
4EWxTbuH1TF7rF2QFxvmf5EFhFR5wqGjkUJCLgoUV0sKYBk1PaM/An6IPCLCtVkv
mUvqW7wHG6JpKEt6bcRppvakprJRetwQ4ut8IXXbFkGChkN01xRjUHIVZC/FgS4A
LEs+D/cMyMqLcE77BVDq6icQsZV6ovdWwzOATGv6q967p+aNxb0UYKjGQgn7JZpv
I98d6Ky862QNGUmdiJXrMrfzfolDnmbsDQhF4zv6qANkfonjsZH/zXGQzCRaBVfu
TuQlfp+o2DIHW15SH54QXoSHb/SQCCx/uutmRCvP0Trxvc1/1wO3YABbx3ZEZXCL
nfp+UM8X5XNI5fwBDYsQsI8Brb54jr1eg6vy1JbPncxY2oPEpjra932RoEZoCBRs
wpamqaCzWha89RKryqOEMnVdItUBOq+55uKF1CFPdoTnZKXYnEBdDF7zVBYFy9Cb
JMqkwaujuGbVEAEYGIQ6iu4rZ9c5z6SRDbdFCAqP1H8X4pK7CBBahY+vwlaYIp/d
D8RJdPYzNUfc9EU4J3OyJYYv7z815RAbq+ClG1hUOu32a4Fl0X7/41suWlBYM5HG
Pz8Zch5QBLUMe5Kf6+hI6k5TTEAPksnmQE54rsm3VlJTiKnMsYuPb2ofVgtrCoim
64NHyVWrzUUsiQgosHLH0yjJ6xSTUOxF6CgrsLY0JHMDAPh68baX8ElZkWY6eTOX
JsTesSr6soqbjq2OPjU3tA2ef0AyQLYwdJto7oSFQKDcPiSvnDTs3MSZTM9ks3FA
M+Mw8tWZRawvcgm5zGMNvEM/PGYTwIzTyku/Gmkm3l+fi1rtTJPEiUCMQW48yh+/
AEVJ82Klc/YfZmNQSCreN3kOchSK7Q7qLwnMojnIOhmshl0mPSpMIsYLzX4A9Crw
mvf1OTufuMW0lqlKvuLXYFa6y2IvexUmpXJfHE92AlMyqO00oTex6awiKsaQRngz
bxt0wT/N3egjGcpiLATLk6bKnPeROuviJXmGE7kkRDH7GCy+0hC2DlmXEFXH4wyU
Lbdl+wfKbW+f8bYiUrmaKD3Xcu94VqhGCsAl8mOQKGG4WPsesyNz57ZN0f1lARJZ
svFfQRJkI9hD9hq4im8OjSIKdgkBBLy0pmuxgBJ20DbHPZu9q1Bpe6mvB1qawzRS
ZwxcaxHa7GUrooW8FBunZwsIygpWZ1IBhOqtjiQjL3VBnrYkBkIq1g/GOpCUID2z
seIqNYb2bAF/Frp+1fEaUCfSORK0RqemLc3y5ewwUjhh+zjQ3jIFLsmCQk5817iR
DBxwpnXMqpqG+NJJ5JhRQp565Xd1xDjO2IhEFPBrdvzoUxnnXSYsqV6JvzQkfmqk
RTKTop/Gc4IlRINKOGTMuK8uEakUusZIdluALFL8GptmYZSqkRIlHNYsH4OTKjAy
QxhQvWFJNmGq/o5zgRmkiCb/m1f8P/HDiDQd254A3YfvW0k+Z3mEp0IUXMiWyfFD
wWwsHm0dk/b0jDnuXffnrWo+S0u9n1+VTLfjdA9nco9HU0uhE/BMHQCrosZNkPeg
BDLIb2tlL/iB4IhRz1x5a3r/wSaUfNB+SJ7U8/DQaKBjzOkM+F63w1rKrEhO2uqa
YzICfthDJ7Zx3FyQ5PN9p/KCbml7oM8Iy3MKzQJClNhy0mvfr5rD/FdVwUNCS9Lw
eiV8przfGus27pISBPltMtCisOVZtV2M4F26ihZadjRwFFxrB/nrohBtamRpKMuI
oluiOweCHgZnbZTwa9hlLz9v3yIh3vimDYD6mZ43QeyGi3vEP1pQOZZIVI0bNq+T
6FNA2SSN5ORaGRnStDNTfOa2ne0y5OUA43KDbySyB2Zz2IwFjGrKed/bPzyiAuTl
3+bA6UkwoYSWS1qpVdAB4o8A4uUL/D1Yq3sW64pa46FKGCFJevL6WM0xnzGv6cKL
dmd2N7P+cxidP7zMZY8N3jugv0iv89zLx31krkKdxzUVHrlnuwiM0XfH9OZNP3fD
TliQOAIJNFBWliQF8yOnTCpOV64HLFDubqPD8eFs6pQY5PycTCXpoog1SJdRUdnE
TmsCq3hZ4QN1w8Xm/lIBYZLLs9aQguN1c5/a2MexUKjUr1o0SWk6UfZ9DZqmjDrE
QNM/ulzE5aBWIApD2wjpifL5vH/plw7MiBHzcfcsSQkRBStMBpwLrsYlF+5q12xc
iUFnQYbxrslG6r6huD9Mm3NGCFRmQOcstFV50t7+/Pu4OZtT1rg9tzIZzRVDTq05
cZqsOJd3hxVpNP46cdwy5zBABpL9t+io6MGIauVdckai5lDFP6dzbZH4we5cVthU
F3BdVFS4lo49ramnk0hkaUQ07gSKJ+69qwczmH9Ouc1wklSGvXNDXSqHLFHK8UwZ
qbJyE/hzvwl5ikg9fRIVkvnXFE4jdEt2WWMk9FkKzSZtkS91qKcHcJrmV98l44w9
wAdkcd569EHrPC0QlS9Xz9pItzPTdcQ7fqFg/II6+KaHq/5t8B4aIlQdcUFqyZuL
QIGzBPD0X/Cslv0Y4m4zDnhr+V8KEEw9LSCzwuyFD6CIfoJZP3aoyKr/lvHt9eHe
E+09sh0bXmREPac9khd+LStxLUzj/e/PKRGwRHU9u++gPbXOJfvQLkKG+sHA2T/4
gTpwH4zpNuKPTJFBFXExIYXDvB9JY1qZKuyZVIdQIhL6F06uycBhLDP8qXsMXCl4
A+CpsbZkvT+aYpHqmaLNtBIYInpF/s2K7XOtsW92Gm/MMPbbCqKJ98OaIRzFrPOV
hmRODuGFiZSHuLRKTOBbdpZTtIY9QTKsecTJ+R8x7r+OgGWF5r1pinutANnLUmOj
P8u5NHW13a6Qj1+srd31D+sScbgdZez7H9ZGIwA4R7I5uLBWIMe6HwVOZEe7dan2
SbPKZWl56pgyQjYLfV0hN32qKt9kvA6UTIBK3ez+zrbvrDYyMY1lzTXQ2uLurnHr
81m0mi5TKOj0E2xZJtig6p675OgJTUEjZdzKAlRK9JMDeMLgrXvE4bs7e1ph+L9P
vQE3WLL3kCzmrpFzAniE34RFZi8vfZdEoVcIJ5fqg5Z1uy5/611NRA/T88SCL0b9
AC6nJE7t9k+qCxgmrEHKkGOmsWq17cFUpQKBreOxEmR6iRR+DR3xOBaReu1HGo86
WBfTze8ApCr1xaif2BF8X/2xceR1c3DyQ9+x8JpKQzp4CT6nIlUMWhK45fCPOyJN
G3LFE6GXJk+4z3BRh2hIHcoPwHnSb1r1vUhh3Tl2qWgUYneo59PvRDsKGnJ6ejjY
G/gbPD6DZNtMICXyQ2MlZ3U8j/I/FssQtXQcC5fLalGhB0itEYUwTe+Vgt1YZzX1
pySh+Bsqvgt479TVLrHosCA/Nv7dcMJANVd7sTzyTU8uU6eCLeHukgUd5uJ/zkb1
j/nytXb855vPVqe0cGRmFiVGNc7rvMgC+55uaO3nTmxuorHDvc4p1l+bc7YmDO8P
rmd+t33v8ontJhzfg5fONgDX4zfdtvmT3GwmK5ZpxNjzpF2EDFb0iep6YcbZ8FqW
DhyofY2vs85fMP+z6ooI9NQhhDvuFhOw2dl/jm3ovZgzbhb+rjwvLuDbv/xHt5ol
mmsua/OCXmOmtBrRBMeQ2TYzoUjB6Zl/QXHT4sb64qYA+hNZGw2kOGB7Jh250NIe
yts/lGK/nWFtr+wf2ZoDSTmQ2MRLv/Uc+fJ+MXyHaPIldnNJ8P1wyUDQczxmhCIR
jh1/AcVTAb3nVXoYz4yffVEQmzMmzUC6XceTFxSkSm2lWpPYjE2Xt5oXcS31+dVb
fSQvQs/IbWUbjPjSZTEtMWzwFX92qLh4/Sn/u3sNERR64fQaw0uySqUlVF9jQQra
B/18L8uNrvm9wB+nPT8t3XrOXIaTrZzvSB/6nZ9TQryjwSjpozt46yg79lzMDgMC
FTHJpxgRkCblEN145ezWk1Des1BIT6dqlzBEXaYy6xdKIhLclkdUFJespHhHtR3U
kNCvU1+sLrU1zHnOYKPbCygpZHGuH4wcMD8ClbaIebWZkFCs2b4DOibASIfcHfm9
Hd2zWjTiiHqahRAJmlStnCd9oPWclq3N9Sj1xEiZ5eEwypWOcWsCAGUX/R3A9TBK
S8StVY00EJ/xTKa6ZPNfajsFm8j3JCudAHH8kvLehwfiCNW4vl1sTUakxpZ/Sqy6
il91tKMvrkutl7YK4U5d+J2cNprzIuM1OM5rRVdTnpbbufZIGGl0NoaJJu8VnCvK
TIdkN7SaNjcXgPI1nbgwfaK2KDN2dxh0/QeqhIyxAwQu1t/5W5FenZTk844KQAWW
cEs9URQVB5NUGSYURiNd6Fwt5cfJePOAoljpdje3k0mIM1ompmrn8dYGzIpHThJU
kYw3P2uV5NgcVphLPH8HOakoIAddnYobNK5+AnY01h5OGruFvpgxeFoaIzf/Hhi9
6JhzVDAwrQ0y6weRk2N6ZifV2ZMPE848V3NkFbvT43xcE+3vpXLqUagh7lCUNFNJ
7P1TFv2nXDGKoWjfCySltd2j2H9UWX5gTaPuxdO59XZJI4Lht2Oe0dcGeVIOxc8n
e/vGANv4GX38eMdtH0J4ayiRCB+PWsQ4orJrGYgpnkkwEcA53cixT7pVfBuhVP6F
zHQNUwqaew8KtZ6WFHeLVYTI4s2fMgpe71C8b619XkzmmGEN3eoEK29DNyecJLwf
50ODnRz/as+GMiW4LVuuSsrVMH2NncHp8SLz3oVn3OyC4DdWEEjBYV3+0IwW7mX8
OwZbtuc+yNt1g/5mHeEDHpb+ZPOGvOLR0iMbBIkAuIq1UQamMMq3RnqD87hXi813
BLNoUB2Yc7vXDVH14v2xaPIAauz4W2/yWuZCpODjf5vRDX95WcUEoMtwp3AIYsHW
aUWbMXsEF5jCMMB+NzyRzX2ZSWimzrro+C9tHczBmaVz0ANb8pr0HQrqOD58Gy9E
gde62XXw4FS8anB4G8hj5nwimC0LRmtOYKSreGGTxZuS4JsvFYrMMxQLLlwZInXd
kwPpLlzgeEeLDMwCFUyUxhdPIhsJaKPSK+DfVnQfm8SV31N3mKlE1o8o6q5poIGZ
b622nIae4yN1aPI+EoDyHgA8wznVdqCJzoVkYm0clLIm1o3bF7XXQWvwtLPpzm8s
xtZCTtfGbZPphOS4a0y1OQElv1NpjTs7a7oTAsraqdmvXJw/23cl11SwVDa2qEQ9
8yLqGFXxt+QlVYoXKB/SnRkKYQwaraKq1KMFxXyRd8g/nudpEMCrAXTcN0hNxoCf
7X8BRI/uT+3HRVQgzpfSARYtZpWF2P+5gKGWQy8a4sTE5qbonm6un/xWN8PS0+bq
yPt+2IODi5LzhWSUxYMT+QdoxE4qszvILbGEPQDNlQIPt6I1fTv6rPaVp2zBsrr+
tfYzO7koR0GyrxmzjbAh2j+IAi/cTuRCWhlJKs9D0h+Jdy5H3NVm5iSOYqn9pAIx
UAkfcuz8SecdOV5qo3uumnDwqT6lublNZnnEUo+pXu8naNwMkEqwBy8mqWEdxIrc
ct4pu5BnWgy4LPawBTIjEE1vjsRmpukmSUhGRWfzYttzbefdscIMMznEVL7gnrTg
zhLvx+4i731lbrOGhjoSqtl6rSS16oXJZjKSREk+ec2vb4Wavn3yE012dwdJq7pU
ZtdS2xPgelhz5P04dfY1Lu9NRPkEpWqKnkyIZy7zGhdYZHeX4kK44+t1pivAlCto
ROljg5NibSHJw8/6uA9XvHVP+7I2sWbG3gv6iETqlPcO0k6PXOZpDHQbxREWLuAA
2W/limEKruyZELmy0/F3dIU06i9e9sUic+vq1FzI3LVrmffo+YtKhgVMMURrorQB
wwPYZ8l79ON9iKYa+NjSaIGCM6HSYv9pq61B40H07Vx78xx0wzJgYIaTLyHt/5zB
LaTsGjJWLGws0ZD4lEnNlMVs2bWb3xGuX1OvYvPhyerXSL6BvQx7d9KcUSDmGWef
wBZVXUCSfwJK0YLz0l8PjRf61lXbRQDph1yo0RiSztCvtYa6cEjCAFrA7LI5bgaV
xEIW84WxIGg5l/uqCKFhMt13Y24bs2ovc5qC9qkVch1S8yI5OTXWTcUsPIyLmD9F
f4s1oy4Bo3FzqpW+xb1G5LYBSIkwnCVs6Jg5jdlMjaQsmojf4Ujvo658WUC6DFMt
GBHBndWKRAirvC6fC180evFRE2TdmUxL5FeS5Lxqf7VNEft1YJ1FVhTC3vx4MUR1
/3Tla5JzN6lVwGOpJE/cf5/w6n42TZaYAlvMzb/8+VIgWNmSGhkpnaeehtwOH/DL
9vI4mCsKcgCe9+7FoTTATHwfRx6BEg8I/rzf79MPW3wwYJDOjEbzb8ssuO1RKodF
FugO77S7GJHNulvsKsd43+3ZkFOtv2ezz/XGPG9v7IA9ElEpPTxLgaYcF6SqfjIM
kDCLqiqSPQ9QL5ky/PzXP9HWbeH25nZ/dZdasu18+fNb9Xll0QseS/L4z3+qmiF3
9CXfKPh6gTSKlT7J41H0E0SCFZvMX2uFTmHjrF6ZReYkqCQLTbpWcwNTukDXXTHS
jXMPkkT+vovRGXdBbPrCsKRV0EIAT/EgKqgOf/jyjfdx1JH+k4HLy9XY604D6ma5
sJawn+g1oyPGGMFzUPR6XlZACxpAQDbW/lPUbB0EZ1MbNJuSPtEhQCfn8ID48vBf
Z0J62hVUcwflCsDuer+ESkmpiCLeXL9gXEyOb04metPjLwn+X/2kjZDHaUA154EZ
5KAlEtkqooxKLfELq5IlDW7DMbGAY7iJ/M3M95WewDZafSDfHSKSxRdsLln/yxg/
zmGZ/8nf32RXQMRqJ+WhXVJ1mmQIwftV2tqnDjYx6+m8i/VvOvqdObWokV03v3vD
XtWkuqN2jT14WeAZkkCQPntuOJ6P0Z5RcDHSTTtNKlnDwoyQOP6xqRHnR/0IlcQW
UnhMr9bUHRKr4ioz6rvF3Ij+1WVFt6Ogsy6gQeWH0lEqPDxGa36vcKo2ksCEGUWk
GMlpLOYcHHn4JeaoMtkWx2p+yYnHLqRZehuVixW0I0f1eXk1Drj6ONuJ9NEWPCea
YRVK2qCblSl4J91waTNkj8jDoxn0wbuNjNJWM0fIyr7RnZF4YmysXjDv/zMnxr31
a5Nmr8S2tV2Dyatp+k5741et2nCs+y+d1/+VybW22NqkHp2MF56gGGaips4iwiB+
84D6a1eBQn6cDmejyWTOg3BR+/lLfjqxeHsXCYac5IpDvqv6fjYonAz/tIUgXkcw
c8RhxQoyM9jVXte+uFJ60WZzFn6G7VSXvqCVtyiv9r3jPBNUt1uYlejesRBfXKEY
0E6/P4fJ1Fe1iy+Jvyz5SpUlHFljjH0VX26UEECwVqtCmbS3kuXSuknT0IIHfDL+
9vKM2XNFt07JZYV9/WgwbwJhHf6rCpWCqukTDQbhOkBtXOn5ouPuGvFbFfkIuT74
hvudshZcLSRpXiutbl0R4WWjsri2+hhUVt79fk2qjZhFseYPKAexgFN/SnyPE0+x
OPAf5uXkFVDnyA8ooNcEAIee84hXBygxf+nKJy+38LQ3PqOX5JNSlNeB+rjqqmZ5
2cVf6D/mKfIYOpAjyvXv+ey6hKsZM4kyvugWoQZ39HI2INbgH8D/9PI5TjKdFcfb
7QK70LOJeUex30+h3/xRfDOHQ3JoiJvj682qACV9Soa3ZqkGbsc3mr2rc2jYYNGO
ozVAuZ1ldU3KGJzgTF8h2+xRqQgsc2ArbPZUtWCpvd53ZucT8wfKA3h+qIPbXL/P
vWzt9FRYA8Ujm8Hw23fKlPDeeiAXGFZt2cd5u34RB1nqlaCrgMl0Bde7i0dk3i//
rA4EVIbzfPsOrKprtSgkSU+3Op83AzNaGWwNQ/jlocAzK/aVsbztpdz+qJ3P2t8i
YHFZEYF3dR7blJoL4kmDGpok1JjJlI5q78dWldNIU2KexB+sWgVRpVK6KPdYZoXG
FeyxPV28EQG5w0dQQJ8ptx4PTRyRgIcUDz66A7ce32ZAU7gbsdeFSvm0Kuqx5m+u
bx3yOda3xG2ldyXPXFdn4bKJN8vQ8bRu/7kZ9mr/COujUN4Ajf2f/Y45V4kUuFZZ
/smvg62Irm7AzqreOTQIOCvZYhXEte7JWRZSoxSBNeqi7ueMl0lEmzA8SRft6GGV
cce+NLj9KhaxQgoLZZjnQmMCCrC+j2WG5LCosX2Zim3b7J5allpCY1zJPBZDuLBi
xTpt2zYXViJz5vwmvH5PIckQdF+V87tx/LfbBnXRXxfxte32mFisxLvrdDJTHQ6K
M69SQvj4V0tGG0r86h4Mb1Q6MarAVtASURDM9hPtvjGFzmQjURDh0CDdtklIg0oz
KrpH/kueK9s6MDPXT57R9CRoEGP0PSuPHPTqd3BTTLumJiv9NepCoLgNPaa4UJxK
cc9IALFmXlizesBq53WmpBNje0XaqpRj0/P4Jni95tZ7oOQpzeMYxVQXbE8lEFPL
6ucHRA0iUMx0JlMltSwkmXLdgYnMORI+fsEXFr9qA6llzFuWP3id5F8E81T58ans
nim+aEkuVHIFK2YyFYvtjdZE4uiW0MjEbCHVP1xgmtC2Vd1lcE5gN+skkKuRpOm+
F3o3UxxcZXpnWXu1YKT5Hm+1SOfCOmsaoNDBXqStS+HttCRBQpFsDF1ZJReGgRuQ
qfebjzZ7ZPRcbXVyJA5ILIH/rPxITieBXw+XD09R3Mrgrt1gq9y1zopBJTw0gliQ
2/FMcK/e0uyeZo8RpTLC1gpO2xAArvwhl3f6FcU1N63F8W061mDHGXwcZLftmC2k
`pragma protect end_protected
