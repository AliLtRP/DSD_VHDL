// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:37:21 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
pumy3jiAuJeuuHaS7T8gPbfUGjxodQhMrQoO+tsmTtuTN1XGfvndTPBv1tJlJ4gR
op6J98VkvsSdn5ZcxbkSSetFKu/ZZDOW13xTAuoufnAIlz8KgI510flTcSee0/ld
uHnxi9zCHtpB92yy0ggCg1Tc6s9eCzgCyBt56U686PE=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 9872)
k8GHr4nJQ0M8AbqWl/M8jNiMRgj+MK/eM+I4eFZQnLjct3pdmq8I9pMHn6HRE404
D5aC7PP2J0naE+Qiz6PsSBZNv6S1SZdXEygove3TpEaiNZinq+3WuUcDRpXlsDW7
M6A563mWWmigxqNshnkEJXmT1gzsBrmqjD+QAPInisO7Ey6QbkxGIdx3D+8CrbC2
012LfEvPGsPapfZG8z/N9fxxTWHR8GstOwh0IDXA2bkOEcUeWji95JYpy69aCkxI
zITDkcbQtQmYA35+O2LArVcxAlehr1TDjZ7p7mY4SUGowqDtCAXcIKopxdiK11ut
6S+3lOAlnx9QCaNEb2E0bli86Eg0F0q88bV4Gpj0MNbTq7w8n+lOlHVLBQXkDkP1
bVZrv8k4b8/D9wtVzvR7Bj9E5RolYeqmZ7ReHvqbBfb3ociD+Um6ZsSR9OWWPhGp
4fbZurk7t7SBgzqmlw5dqsqGEUybVhke3iTLvl9JHG5iLCDsppz2RuN506xAdaMI
YiOjo5damB+Fi1a41xGcteRrAMkqUO4PuFU4tDpqp0z77QncQNk7S0gr2N+uHZhc
gAqd3DVYKEkAoZboSnZXBdOVEcfyYgGXQAwE5/sWJEX73s8S+E0QDTzU1SRpNty9
pVYq7Mypujs7hX2bL2OZ6Zxq92rJYH3de5DLAstTKhT0ZG6l3dsQYFjgNOiYiTWh
nj91psHJ1PaLXl0ZyHzyIZQqu2/GIgsDtHdHbPszoXY9OpQM3ByrAO/2fTYnNDVH
O9TH2DCgIDGPCbMG2dgSJH0rueBAA7SXSJ+a3iHFfyBGO2cg/89rzMK4U8T4z54J
GxdVS1pjf51pMrNfoUkWkcEvAyaYdv1rQB3UxSjlDU+Y+bM/okga10LwvjSphMnK
rKW43fXqenywBtQM9KMSRCOzXGsqEEyqo/oQnhc1sXG+3v5s+4LrYTJaS8vdg3LP
JVQtG27BanjEhhkFvjpE2fsBgSZDcVRtyt2S3l2gBqvQQzMUH9sN2AhkvyVyO4a5
qvprMWbaJEsan17lMoxt10LCwsx+90WjqTeMNxrvgrI64kuq3FUYBQWJcMmJXW5u
8mj5C8U9QpPh2etvg5AsBk1Yf+XyxDPIL52NMd3s5iP+hH57kJRaVD+t758HsbJ9
JRVPWbmvdEWfUjWtjGSPbyEDk8gHLAGFAbgVfDXwskWACoo7W4r0MSz1qNPp2aN+
rX9W12me7ksFQPfJ/XIPp1PqrbDMIna/glNySyjUshefz4S/PRr4ky6HOSn/IdKa
/ZsMCM7i1D7gtMaBtFRpdi6qB+RRTwzq/1qW4CmAXGKhMF+VPf38GBLfdd6Kdh/f
vyxiJ36NiYgIxivPRghyqj91Pr6HpEPYrkLfnPGFQ/C6xKsIylFkPhbdL5LfJHsy
4nd8+JWUI059Cz3ce4CO+jOZ2P0BFmjbHkSJDT0gkGIo4qriq3uPD2m0VCHdyrnb
J8s4yJ+TXOUxOc2CnYvlEjVp5V4svgz0Epd64NLMSQI3Lp2L7HXoJEqPsPQ/Zfn7
mVj1OAcv8HZ8+Rpn5WJeNOtxVMaeboNRoc7KNrqcq7uyUAtwmJ9t6zCnvatMPDXB
jAlt/yfZN1XmoBGIWntKX0EBQdpXSb1V/FqEvNyYizJNkc4G+CBDS4xdj38t2Nhj
PekAGzVdC3xpHj2IGzHFiQK7T56cqVGsP9SoYIPl1wdz+yi8AmgFQ6c1uvZ74Y6u
ySYp3Qa69a7ATboHFRfP7eZ1XUXPexobJb5KzchAATPs+RZ542pROLAG1a1ICa7N
fAF5aU8I7IKamzOUF0QdTCL9HLpR6klr9JoVKfzwd5K5zpBccw6YXxzjeiL1cTwL
tQjQ6Lkw4aCiKzKDVkYWswwJ0KjXBR6+91ablQxV5gq7ZfCMJtlxGW/klQmzatUr
aao0H9FI57OzJwJBdhT9OG7pTgNOkz8yi2rcrR6sKXesgTdWBdBam4a99CJEYp0R
yHZmPjVc7YFma2kgT/lnSG8c+qk72bXX3+gxxwOVi3zZIM3iRNuUY89p8yh0roXM
Kji88aWF+p2lNBAHakhaArcwgitmraCw+Y+GfpcWnDCTrXywHuOcqgxbqD9VruQ5
MlSqx8LLcsulRy/lBGbBGF7Ssmy8IY659Z/p+ZlnHiVIS7IZgY5Hv7D+ZKFb2tuL
j0kY/rCnrQjJ9Nwe6JyDMjnp38LZw5Uz8S0XyzUhbuSbKGppsxm9APLqdrADfTqL
jNvbGOBDhOf2yOuh5eLVynTQ4myxwKCyRzKFWdeCUAVD4D3MKaLKIuhuOJoaiQfV
dBR34e7KBZ0DYYwPDrIurYOGv8LAkBYjtGO6Rx/2z3gCRIqnfmUOcfNtqDtMinFf
SX7uDjj7GSyEKq40gffUp5hLlPGNQCr4WFzIvjq+BNbt2opC7cAqIN6p3ytPF31/
RP0O06Ke1GvJE/Kr9K2AQF+ARQBmL1wNO9yOsOU1Pkd1KMgKIJt3zi7gEecMK8iI
sMBODKpz4xdpvkkrNsMixjpV1+qVoyGYJDfFAR3wL3H33J4jTmxk7qcZEHpRivIS
o+0nFqJLL4uU6vEXP56aVClGXJmkcpYAF84GYfR8TzdR6LhTK4Eudp5QODsT/j8R
Y3x+zVd4l6aV31tJPGPAxL7Z9vIERpMU+0yjlP7LrB0xynTsBUXM6n9hJJPPCxta
+OTF8XHy5PvJIIgYlSkJb3Suj+0CHRocDNV34a1TtFwMYXbdpd/b/R8JYV9tGHK6
fiMz2MOKeivdG0CoRO51YTzoWNlH9Div20h7XjVlF21JRWN+6Gj/0pNK6JA7SVZ1
GQ+QDndx1tC+sfsZd6azAIWjvaDPyCpcOGBUG6DAzpnQORNH7VmhMooNkxjD4yJy
yg86Sw3BnG2SSKmdDYYfrg5QqatAmaHrb1p3KKBOxSNtBbXA+B4SHXrxMLp7wVW7
ygpmKNF8dRHtf66vDj7ZI39dzTgyJIaK0WlGQN4Bl1PwL/2Utx8DB6triLE0Vt1l
tUQxEEzjNISGAcJdsCZVAy75exlFD1Cnkt//5JfhHNuMsEWXhlpreCYAmLvrem9O
gwRY1H1WSEnvc81vKpejOvjPW0N0XDn/KsHpy8f3JE2xlGMGrBF3r7B4A7/tnR/9
H4VcG/nxIM/zrVnPqkR5Wc7NJjAyy3utJbF8iT2L37l3iZ7zOwg2/dfvZpy6Ocvd
Mx2Ww2udmcyVSqqW/WMfnCv6Fb07jx0l/pbuihCf8Ec/XcC4zIRAngtqwhEuFxU+
l18Q290rHig8ORNASNrcKFfEXmUdj131T/3odCfKp1sGeDzIMCVMhNrFPUcbeV6e
mxRd31BsYd/KmX9S7ewxWTF8NKTG6QHXiaAibgg3hf1xJvHrNftV1uhCO4enIL0A
r8OxLPLGcRyQrFX5m2L2quvEB/H3ECtcEvlW7rD2OD5qYhzqO51j2meQut0Vk6T2
HtH9W5X+unJtCjR+CKAueukW/1bdbfoz7sVZSiMHjkP1YSU4JDh3KLeQngnlafG1
xB6WHmpVilgfYotgWMcmkG+ff0hFo0COw5VVZ+o6VlbDjNz4n1lWmSKqlUaWeYYg
pmC/maBsafAT+k9DWDuNnntSSBbyD850sde/YryM4Y8h9Bj92kmpTOiHMtMkRfDf
1XXzD9FHU9E2G8QkqSt/TXMsToMZdhObDGJ7wgUyoG12d3Mzm6sBJruuPJcYsX5z
ZOOwf8qCa1hNu5YgrGfQE6T/h3Rd/rgU0I0soizc4nkID5UoUjdEnzfceQjSi2e3
g95/1xi9MW8UJvWVR27VZ0XkyhHkrd3Cmp1IPn6bhxxuMVprqDATwg1QQaaoCcLm
KXNbWM/7CMEfPUo5ncwbFQlyhy9N7hsv8jlEPNZLauR65wXuGrXPHNACHLAcXjFs
/BbQI0J3bRCZJ29sXsxp849XPXA4zPeisqhvzbgZlVEJPj9LSVxgwRdUZRiBGBBD
fGxKLt4mWcqLnc4+yk/oUvbQdGrCdERGuSgaUX/pgeVZ4Dv0b5IOJWfSckvrjze2
Q9DEkccpzKljDcHcJBmEGcqKW2HBLxWqcyC3deO4FvWki5ztswTgvEW/9B7+973u
L/vjeP7OuX4yW94Lp5MThT2uq4uS+W1/zzMqnZiUMJwKdkVFjugIbxOQtvVG+5at
2Axb4bm6UkvaHl2LHQkN12YHUt7PS5kLawnIPedWojgYQhH6YdXjL8H4bsQfjpsg
IheTUoN1Li2x26iQ27mx+uqxL1lCVVObaRWH13WVNJecm0kpe+7aoHN0ivSUahuU
srlkR14uAmi7jlgd0XGxlDc9Gn6LGT06gjwFgI9Ex/J4vxp8J8NtHqRASI5eDscx
2dB3/Mi/TgJWZrIKtuMXZjCMMLADmTbBJfvpm5LX5Wz8qbXrZBm3iCxQ32kbICfy
6OmymLJPodtYox+i/egsVp9ZQWljaXjOo2j5OI8Mz0YkuLyscA0NOqGxfx5snTrv
4mFTjUUCUfUgaKmGnRdlSVl2XmxaoesZG2y7WtTU/53+tQZd5KN2aLTMSjvDWAl0
TlWatjAy+rYwxdVGIJEUfm/NQhCNsnowM4/TpCZ9YwMoE3lgfgNXaHMDks/9+dkX
BgDVHGagupLtX20w+4NUDj1OEwNmNwokuzHch3BRiyLzeGJEJM/AiSXP9kabNZYZ
lB+LrtjA2oHukDeMJp53QzhaclQMSq5w88Y54faJ7IgqZM/wT0qnR+ucH9zTzY2w
5piLnmSRcd5I7cmOpCMuJVEdTlxMuiAw3z+5FEMSUbROHWWVVFgMbEp7PdVP9S/I
IOR9DgD37gwxHPXnbJ3ugz7gXQrr0tbVHcvTUWx8PKE0XttzmUedz4hziv6ELxS7
OnTVykiha5SrKcpC94ydng60+Qg8fcQceDjGL3bzQi1j4nnQVsYCf806dkEUNE3y
a4qR2HTVLLxzWKCi+5KwmoIx4ZjvW+mIkDF1ePlno3ep181JdOBeARqo2XwvNYMe
eGcSFRVcWtXJe0lJqgYiPCoZT77c9uwmK3R2YIHccZFwj9tynl2Cm3qJTMejLZd2
A4nveWEvUa/50MKLQ4u4rgz9eqWgfEJpUgwOYunimZwB5ixAKjcbNE8vffce1ABd
hIyL5n8CfG2w0RsgkS6mqJRP4THTeqbPdltY3oNlH3IFYzA9vPiG4YqOlH7T8sXh
8o7dwwNVAzplp/ye9YdPRp+AMBhyJGOzNtVlfywEAL8ROIh/5d2HDSnvuLcVglLB
Rsmrnxih7Pathz7AVkaRkfCrK63W57iylYGeeB4og7HZn1Zlw04zOiDpKLe/Rh3w
YEe6dTS1V7Ep+UbF2XLQBzv5o3Aj/vuO0GqVVq/cvtStsaHZ2i+kF3uuRaHQIQZp
rD7ijCgvy01AWv9EA9qnRQhPovtta4YbyDdNXtMCsZjN/P+wRFSDZ4kQkepyJeEb
U2REugty2Pgg+Fg54wSV3TEs6UdfNlRViXA1XcUj6gVysSi0IZtdRSgNvWYyrwB9
RJ/r+Z6RUtk68AKK6DCgB9KVWfaviPTRB96XF9sAw1sfpIcKh6h3NLHbaX8waJSv
Sw2+UW22D8roAtNq7p/JamsnsEClyYR+e7y1yG2/GajJLgfFLItx3DEuyI3Z1AaM
+KXn0bQQAJw/PNGzMNX2rn4g7qLGigmy3G2oQRPXFgdUf2r1K2mk61safkz63fTO
hLFjivxPRpt2kPtVFbMG+eQDXnEoeGgTnUWAKj9emZI6xeL1WFEQhoLBBAO5Bjyl
Uusn85YtlD+vsnmBnVLjXMTkk3Sw00HmoAQzeepm0MGZ5u3q3NubPYD5lHqE0KdE
qXj7J+VDJydWQQIXD2NNYW6e5etramB4sM0XWsbyzYymN57UNTZxzwOvNHaGJgnG
mm02ZbTcUWitK8N+gwcRlPUp6cjxOCkEoDgiNSmGr5WueQbr0YuIRzCq4Rqvnwk/
btc6HzM5wgdr8BuTJUDf0D+AWnKIYPUL0YPUJHxxY4hJx4W9KdVMAYL9MezxPzHF
tziU0UjP9O6Ss5Nxcjq+3LMDNGsqWBwyy6UJgow4bdxQF/LC/1Z6Ywn5ihzDyvhs
mHGjoFOHW6SxzvodVhEdV4e+NdZAbYxeJTqxAQbtvxYz67JXtAKlPZjQ5Aov3IjN
CLE1thHRn6HPZ6Jeoq/HLHUE7KturYFjTOxTdMDezOxLGTw9kykADAuRPHMnkOby
mEc0UV8Ai1uIeEWMvZA2NT7HmNrbPKXEOPrUuFobFq8hfbNs85+T+aZm+fM4Gj0F
8EQ1boKyRbdKTEkNTDY2REiI51fD8DRSwpwQDW9XyEHdypCr0/GZKkOyRYQIHCbg
g97d4BmIxWUB9QNgIQR+YAeZKaiuY4EHgS0nY/HbSptuw7L0OQdHdFw6n3K/f69b
FnhT8Wc1zx5t+MOVmcJLGVfgJzEsYn8nbRQ9I/hP3ubSDiuF77yRsqWCwVbeIkED
gjzA9zEtqKi/Jp1vmHCjq1FnokhqOUeBHVRPPwglIFvZQtJFR5SSIyGkiJKuAauR
cLKUeinsAlMTkGCkwWtgxdfsNiNGdw0+79wDgd531lhtjLnORe7E8CiBy8IWqb7p
gA1u1vCViqjmqyhbchKUyohHl1Q/FMxZBnRclGPpgFCkmy0JSeNGpCWLXvSKyijG
qast6tgCABTzChcWFeqpew2F7Gd41z5Hq3eUepRjPiW66NpjZ1rx6UyHJ58XEmwi
w0KL8u0xUvt+oTNuCPOOAs0HhNyzqbXpobNTNOFQtJT89ln3R3LQ8kwWlPzR5JeJ
timQc11RQshsXRtnrEPkFswpX+5CKxEza3atIHoK3IWN3wAVBJZQWIuIIjK5yHMS
SEQ4MzdjyXa0W/RK9rq1gaiCgti2+63PU7wo7pKTqwm1v0bzr3MwWLpZuiLVuL+W
Km8d/K75cb63NM/pyyck2Ad+sCkprn10gYWdRok8MhKwLH5kRrR94mQVd/o0rCKV
rzBByvvZfmMQ/PjwHXhb45yKjbtl9FPdw97f1OzKqaU2EXVDoV1LmtdSgFzvBkpY
6J8FsIAUeV7sAj64G+xbSzcy1FOg5pckx1W79dYGuGN7Pxpir/W/DA/BQgvDBBsV
jJK6NtnKhZ+oKm0YhsIYOR7eju9dNba3722Uw387M2pxBO8JcyNDsjuuGC2OlhG5
utIG4K3p4C7VknBf8BYwpEEUb40r/2BPCF61HaF1yxn+eGYclnE3xCfs4kMU7xzq
gH7skFh1zVwowy/RIc/QEt0BN1pWU6DEUjgHVGIOYgOBIRxWlrc+1C5kQELDnQKD
lMHTxx2PQprKSG4qi4kdSd5eR7yxG03k8ZuKloBkXDB/JwPxm4hiFZfFJ6MDNtmT
/BuBPueA5XxtqQ5Fu74n8FNEdal+QwGDYTtYaC/wTQhTFgkqyebMj6mZp9AicqP8
g9GFmuphDs8NatYY1w0JtIVjfWX0mnKz1zXunUPgZMBEb4uc7xGe2Wx0JV2dOmAD
j1a21xPBuQ7aHwIpAiOxfujq7vdAefhrJCy1Uw2yj+IbvFjXGcUsDsBU9ZJwzGnB
WCCVVQeRv0rSxqOXYil1LReswKRLoauthDEpq8HYDlJH6NqstPtBGiRH9XLiZSBW
CaJbhyM2AYf7cBgB12zQLGBB2SmJX2pNvJd6AaRNqU23tMMDjr6Z65YVaRckltPL
jRHStASmOERgIvCrE7oZjWEBUaQR7QauprRYUo23tKLYKlcFQOLNWX5wbCuLuNgz
gyQsbG7Q7rZmB96jNdoF54FYhnBu4oBAXwSUos1AIq0uDHm7vtMLb4yu7an2e5vB
gCWNOdeGtztgYqmr4O0p3MJbFJdvCYeKrG35oYFM9Vq6XfMeQ/9j9y0vWpId+3BI
u50yOLViTS1PVzxUl8ZmrsZz4C+A33XEUGx83wkjlEcU4VGY/dy+Dsq3gcVH2E2x
skgCyovjAVIQ+dQnhw8MxGJbmhstTEjJCAVk5coZ7OZsba7vcdtQV8dTq3R/VTYZ
FpzA2Tv/HAzkHVSDmokTZNy48cgEdNsXioq7o/jlvJaM+30TwW68taLJsmN3yCoY
pG91lpnPXjdWwdIZq0DprctrwTZOGt1rLjqPBvg1+bh//pObYpUvVHURIR43eLTR
aUVAdaEdQ1BOOKqzyoeCpGevLJn/MkaiS+TAQW3VneE0OIxc8sH/+NvoGrELG9db
R51ydc9XeAYDglPyX8vuRK3q66cX7CUHLHw8NAwsw3JJRN2AaNz6lv6d7LyDcHDY
yU++5+/j12LsPM/qIDsgRFpLTot10QRyVCE7Ai5VxmXHvHl3/DXstx7mhEq5TBKj
9YC3VKtj16/MkdFvKoxV8QDcuRYwQJZgyD7dpmTiUxPg+BrL7IGLAnSoOvsRObF5
nbWHa8UtxiJ35HdR2dIdV7otVgs5HIGgk1ZQVGeNjGmS0sHsyiJJkKlIzHBE+msy
MY30YRJF+zugQjlXbwrcobxlMkGbi2d3+4LTTJBLrc0h8/YkMjkV0kAtGQsNZtkW
ET/o7IVvAV31Lu+LIFTQkMltPwvfixkQceQzAnnaUERNmBsEDSPb4Xt0JMM8PPUC
SR9wpI0ARFKug1OgjdXXYeSMC1YI8kxQgHm1nNIEb3Udz0qdSQd2R8Yhsi/4KI62
KmlxQoUC9ZhGztT8DQ1hmukM7bmruDpWtOa33HG32Qx34XKzD+RqlvbgF8HZCwAQ
g3aTmyzFIb3zswuonO+fSLiJGUlDonra60Vo6zXmVbywG0Bc1VOmLicJT3I+jlU+
Z/NCRk+AbLS+o0qLcjA8o1Wvg7LAPRPjRorf69RHFpERvbx7ldJTrJVE8CxGz4j5
e+4BcEcqW5u+JgfFNHRv7Q1nzHz/MiQdXkcgyhkcqnewa1+LUTvv10izJdlEes76
7vLTnT2uoDteBNcYl5FrHwud+4gHgGbaac7nS3hLIqodoA5gZkvvW5ZkDreV58UK
WChVmu7/M4OjJiD998HZcHO4vwLQbLuRLuhM6WqcjavtQH29wEmbKEDyedvuylu4
P+GS829KUlEb4i5HdvRhGb9cV4qrTh0PoxPL+JvEl8kQdDSkzrAfwNnTLmWrpDA5
MR02XdmCy68MzDP4wwhbp7TZpEByJduZk85ejgyGdqKqgRi4kzSZQs9FRJ0bUI8L
9J+AHc7aHe/rGax27A7EMEGLZznJYTaUZHI3FcoAqSefaCMpXu58OVnmLZSxeKCb
Po+YL5sGkIrQpmMsrQ0Wi5BxiE7kMiYxpog01PN5cqhwnWDOVqNAWJ3HBL7ICUoK
QkTSFvDXRhhx/YU1SEuQUojmnSnQ3Vd6DNtL2Uv/K+U8U9Vi0lbesNum5ZknryyU
Mg21w0SmaU5y2ktxstbZvGIGEssRQFyXDCp1f5bjywUYHxT9tfYvZl1zb37rHyMp
ee2bA9Q99sqQ7xNCrIYd/nnTsoz4UhrEdbGcbqMeh4a1Ou0Se+Wr5oANt1owzcYw
LKK5C7NnwGbNOjISX9dcfAoFziG+q+as6KAWIWje1al/xfAjsSAdLqi8/QSQSvPd
Vkdk8VY62M8H/ojENXlspe0Pq9OzGdpXjipQcx6dKBO8w1mD9ykAO4NAavFIRHf+
Yp3WzmjycZmxDsOFw06MWQ08mGjSX5yvDobY8JW6TGH4oMoBfY14O5h942DH32Y4
RafjGjC3uwMQReABjVoNdHmjGJlJMrccJPWd+5o5t1Yx5U2oaoLV/nCuxb8+BkZW
KmzHyO23499EwCOH8ItE/L6nvjlKixEZuZZ29YOO3Vj5yk/YiH99Is/vuE/hfGbV
htdedUC/F0jak+HhGvYwex+uhLqOgy2XWbVALyPvTquthQZEauiZXk0IfFqBb+cn
DpPQJ+h6LUU3b2LWd9xGCerdaz1a0kbZD/hDThgJDsydfBQW9CbZiGLf6pnwMt2j
hNt1g1U5kA6XOY3S27WcGwpby7kHtcJ8RVv6xM4wGxFntBOkt3oBowmo5La/nknH
RUcrVOPgo+huQ06GJ7Kv8kv5Ae5wgTEN2tPLNXq1iRk2JvPAazrmYrF6e11rCk0U
/oYdfUq58cl2CXxDuz/fzEmS4wc4hcQ+06meT0hoV0D+atyW1akHhVu4jDECtgdz
XDSrDUqRVYMP2WqamR30MONrrsC2dLd1TV1QhRvQndkuUCtYuBnVco1NIgdKbjno
lN+JNDZomH4ni5zUTVSGST+Ut4yzOzzTxHX6jH706A2KcYX050AM3TmtZqEdJ1Cu
0xO7VSINSpkGOKeZMsFm/5R5aJf7JjJiWLhgZ9AlXpdZDPG/e0PH3muJzX0Oroa5
sQMC8pBGedJEEJ2s1sImOxw/n70N+CjRebsrskO60MwCdqSn5+WqZ8/I5667BSXs
hJtL/whCWS0DrJLrnctWigg8koLJflwfUUGcoiBRaKAb7OqPrBhPUmBqvUbLm4vc
vnStI7PXk+6S5eEw7pYY99wFhpmFJRyydmnHrjFwA3+BKLEDXdK7ZylTtZH+hRtE
o4+1uVJ9uOuZ04AZv+2wc5cn2/zrq3Q+M2zFDG67h0TvSW2ROLCo4oDB5jtvjGs9
HkXmaEXmKyLjmvAzO+Zogp7AQfcPA7K6RhMTdGjlq08eBpqw8o2hrJG+Xwo18ZWA
5NCABj59FIFJSTQbADukQlTwtPs5kgHe1pDTMjNcetHi3bXAekEGoZzZl+J33uOg
THwPL/1Kmor++0yMTgXPjYfA1JPEbtRGuYORWqsYGPL/HdbE5lzo6GjvQDTYHBjd
hvhxeyt4etUqzCibhUUS1TVUuUZ+GeqHFPF8VLHdE65/e2DYW5RCdl4ZQhq16GV8
xanaZDiC29xVBoswIZCdBp5rs0gGrwepWqkP5fXmXA6NseeiSFPdL+GOY7OoyGAL
h6xm72Niv8Em9eO2PkRGwwAGvyBSFh7EaW/vH9cYjBYnbxKCwLx9gcPrAsbo8khF
c6J/kfuTZWbfzBYQu46fT2VadBCRP16HkA2nlY0ghupCVudj44Wl2L0B/SA5hg2G
bzfffwghszJdm5B2TMr+PDoox8mPBmjdElvNcwrczFJEoO/FO1cw/Ai9rVvSuf43
1YfzIKV/f+09TY0YWSqaiS7rQXsI3FIuJA9s2IRSuMRqzk5zJT+UZGxsnd3OQ/7M
uANzkIkJE3RDbqPbsrmCWS7ZJGDLdhvrmQGZaNIhHPVlJMb6bwe23HOZoBusBMHg
SnqLyzOmfK26V4jzf3oQy/d8zd3M1V4Dl01FYaTmpnphWjhKOG6Sb/o/Qf6u6JBZ
EQ8AuwdjPQLG6zFR3nBjbTigwpw50O3Bm3ZqBKFLrLYzfQ60zMtODTuA2f/eH9NG
C9hMAu+ODO75I9XCfGO+2mkqhM6ZrYghRIW3SQqPwNpwaocHJ5fVzig2uea7vuLe
g+NSTZuvQsTdlbEwpbJw4QnI9aYSfiVk8I8EiBSNT2RI3vGH6uLfoCvidA2cvi8V
fQARPhwox25Ju7reNeb2PcvfJ3B7cK4akF3MUgFHPK0bLahmGIYcKsHTgX8Kk4FU
Qj5MqWT4dDPn1H4IOlMgtCq+h3g9QG1OHxSP6ZJ963uTy5nmPU5+rOhbRd4AMMby
srcker5tdJIGoCoStKJWLpxq6ojalmjuknwtPixl2DEZpt8bcoFmtyKiJJQ08ija
k97YvWXFjinI2bdkGrVYceK2TQWz+B1CyhpnJNWvjHg7Zdn7/LJprgYeDe3tUJDS
NfuMLBj95x78XMMcHYxoQrF5SCaYwI2NbcHQexdyAixZAGlTIOTggAdQ5YHmoQvL
WHHSp7M+HNMtu/zZzvB9TnviBcnwlslDJWfzyT0Z+x9Ly/qQ0jLnQg5WCsLyrfGg
7fbvDqcTO7UFDdES7INsPI3felTIlahR5Ec9PHydNmoJph15t6pDGpTPK2d+w4xq
Une2StnR/vd5xqxtkqRNX3j8GL20GW8amcIj/+QFfdnsDM4i3Mr/0w3NZGwrI8j7
yFZrJaA4RO1xNmnmlE3dGYsgkFmnVEDWHFewMV5oM7QzcTZnujCFD2QkPtFPtQau
xIMcFvcJqaOq8P6VP+oDC/gAW4k2GxtH5JRD29g1Ag58dKt3RHn1ZObhakIRsh2L
4L4CObkqu4N7LNzLwOR1cW68sPF0eCYauZ2uEuYU9JvVu/N5dBPEQUaj3cVnMacQ
JVklGIDR6PIrmX2CEtKsD3gg19+GjAhlVthn/BC3oq7bSlCmYqdvBA6l/PNUtDBd
RIn4W6evaKvm7n7y6Qo4s1036K2THpIgnKJG3jeDwG9UzfvjUN82nbU9R4/1avuH
vJQB1r6q/A90CWAvQF02W8SmK+rKbsGYujUUGV0mLaPh79yRiMjkmjfeuO+CQ5Z8
CcCtEDAbhSYGEMHnrbMOmlapAFkQ9S/xO30NnkN2U0mZ9LXl5CbX1JluQZXScRin
eMadDUUUMsYfXlSuC4OmQJf98cFGmebDKbYPkZLcuJlkM81VCJ6O1Wx7p0zRXt9F
rp83F20uO9njx/ulK4MalVWxH+dB76EdkH69K9l2ySAVqqB0jA5b/te3KM3vh7lq
IrxS3g3vLOBRBB1Wz2omDQfMx6G6rHlZV4rMT/et39QrstHyxtOxmOWany5zCsB3
LdGX156Qnap2o8zZmz1blCHolyXLmXHcEeBakuEnGXNZy0yoKl++zz7ykc8lFMvR
KGCJ6OkSUioazRY4sG+pvzUfztC60Mh6t8oRSeM+/GADf2ZFR8jDbT5YkSkNYpTE
kAkFd4hiYLlXg8TRs3+aLf72WVaa1dVmI1lAOSP/EdrkxI9X0IQZM/COfRkZGBDy
L86KNtd//+tx/Uzooq8tQxrnM5ixgdU9Rgys6kucGmdRo/dP7lMshg76xgT+pnWT
k7XWS8JbiBj9//4fk/JLRKpu9R2chlA8yO+3sQi76rtWw8/UGbaUUBaHzGMctLAa
C5Wm2INhTrnLRpjAqiG7Hvh1PUJp4uh4lCm+nHohchAILR4esYodmlldLp199nFu
iOojViS9koiaZhACCN1i86dZcfgEAXh3KeJaaAWDmQv1+lmdryDvmtCkDltdQjQ8
B6/TbGF90vlEGzn8vzZtF0Pmm9FBy1gvQF/KM9ctccyOFeoKrSEvqozG3yCXzWic
tNP4dCQYBBPIV/+ZdNj5uCMNhP6oT80H2UVvGQZo2C4=
`pragma protect end_protected
