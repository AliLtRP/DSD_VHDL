// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
Eus68bYCG//znkYLM+FqOWGEAqVzk8+d08mgFIGFwB3nxsDPxx5BQ42+zFU5PLea2BiMxRBHo75x
dn/tavkQZ6mCwnh6ifvC1gJJ4mFyz7jlPZleLxKlnwjkhSX9JMMKOXVNqkSDk3XCM/Gp0KvCd613
w4YrnEmPBvWJA5tdyts1aHQUOXB8CgY9NDvcQ9Vn1I0/ePWcZ5d5/j+TKTRDg+eJDV2WKM34zC7T
GEeyytyQTyHxqI78I12g5sW9ODsoyi/xI0THOFjZYWNPdGFY6nAP8EkAyLekE5WWFXJwAdyGox3V
KGl2ob9FYTcfE/Ua+jxvZBQ6tWJ1Vf8EZ0RUug==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
P1RQTvCtQ0p/TzUezDya315L03+ixGcXdN3nhzSv4LdpYJkowqcxiZZyltgP2nafyVOYYXtAFIel
qD49mdkw+yph3rJx/hh68Yk39e2c8cu31r8mCDynLUESzOHCRZfeXSw4yw80BrX/gLTCD2Wf54XM
FPCl19JTQezb31MSaJ4yOs5OZ8m1RoKIOw6oHohdGnT+rVO8/AN6o0KDoIh1w5CEy+/KUPalL27z
tFHwttcw8ffVUpLoGN5LTBftpKRwDXnc2yXFtxDXA87s+YkkWD7LBZ+9+KTdd8hYhgIvZKWgWWij
Bcg9HXLVULMbYc8hGORiV64qrNaPjA6Jwbxxi4C8BJL00Iyc5ru1sqQNtg/OFOgdqx1KNQtl3Kv4
T7f80XW5Gn4ryc1xJxne9uVoxuXesWeYJAp1z3859rY6cwNeCttaqs2j/z0F3d/8uKWET0rxxJ/N
McS5Ezpp/GDlB/EWln3lJTrpuzyDT57OKC4y+L+9at2UtPEct8d91eG+GD3P0MNiq9H6jw4oeCvB
XWBMYngOepZHK7UnCDZfxFGExaY65KCG6LaX+TbOFx/z9Kw7kOw8dQUk+fs0313IQjmiE5zCmKiB
VLpsBRH/BGUI7uhZHSEy0X1PNzRJFLQprjksq+5X56x6pjklhVaG7UH/pSQ1OFviZL+uhYSuMDDR
zVmn6fFHFpaf91BMqIItUbppIAt24XKvPEE3N7UD1gFBT8eaFOts2yKwOFb9iVVpxz3whILxwuS2
7PTvVp4lvUUHaKBLsPDwYqtAF8ckLVMvb12zcMhyty824EvUFqFPL+ca18UmziwMgwfwGegxAlzL
YFvuSYqHYP2su34hpSbEVFq3mVr5jIoqjohsYxc8IR/0poeCLGC0E2+rID0PnHKdU8G8oryaMblK
XZEcxtQh404E6B2HxChP/fTT1GYOXHKzXp002ECLl/MEKtn3d45iwBSm280UWnItSTzlkFMiOkSF
Weo2+cLN0YDeAzQi8OWt7+yQr/92nzLb6riEZyK/DrSK7o0HksMqgJtrYLBxTKQPJcLsDUzGvui+
QikUhv6oZ2rBGCDHg6rsmGmpX7ihl8ezJSwVQz3Dm5wNbu3CEfy/HHY/25Wl3lX3FcJzY3w0w+qV
of5UnH1NN2D+JedLgSsdUr1mRNSu3gEPELoPGIPVvShwZ7eov7q9LcrGOXDO76u5GIExDYIFc+3E
iJ8DyMiJF5M5Il8PdfAkuAy2MmXmSMrFRpiEH+mxmiDwMM136LGb7bM7FtdRwNwLWk7kWozwLvz8
P38G4OKIt9reb5Rt0WEI2KPDiDixi2qig8UvO4IfYUya19f6g+QKSeMGGWM7IQtgOxHuqI5/GcKC
BWoGdWFl9Mig+x6bVb2bFy5SUrXO9busCnB5Bd4uJHHUNhoZoMNUJZ6+cUIStTmg3jE4+qhqmU2N
LOFOk4SZuVkQ9lelvnpQKDLqrShhtRyzUh4wBvqt/memfTss/dH7vNlMAAy77yOsJ7NoU7++jdjk
MqmRiwycjovpprFML3CeD0oQAf0vGB9M/9DvNtXIEbIXQjzN5B3Bb0G8hOjzpL0LY88EfK1vkmX0
ezK4pnXk/OXAMaUIqv0RzuRIconVxJ1+UMW3ZThp3AMn2IV9M4ecow2z7wG1XIkqDqB/VO3mv/Yx
gIlHXLzaJtqRH+rJoNowjzAm0o3Bo65WjJqRq9YAcELSWzZG4CEshE8EhkQhMpm8OL15cnOCGKLu
LcnbSHA1+o/aI4ReqdgDrnVrn8aBJL+X1XsB4hNBIGwoxo3eciHA7eP+iUibWl/ZAv1QU6aZUKtM
jMMGN0TIGeqnzlUGHPX/p99+G4Hy7qD0FKlzvyfAjYgIhBY6O4jFtQpoES2E+ImRh1ZZXAqhBDT2
lCe+mtgNydrv6gft0Qqty/ac8SEvIFu+axK8DCl85NTOjCk3fsNkTIbIrjrUSxAxa+ec6PLKEWSu
sZyfOdY9DoWt+saxmm4yzUD9VpjsjJ3Fx5nWia2qmLRPLHXCYuZ44R3xeQPRjtXYP6KmbhmAKB/T
pHjiJax8pes9zIfzy3EL2fnvxQi6q+W1vBwF/n/cgC7yKRh/zvNnpixgT37d6qtx2rGwV04gbNZe
Y+ugPrwhpsi4U6w11Ibbw3ilmZ5BD+J9aZzqJZq8ksS0baJD7Iglrny898E8knvKthxGDsYPYzZ+
FjcRXKij5/HXfheNCnaKMqquRIoAgZ5Ie6Iwqo/a1ZgfRnSomf6wD0L42QUXF48VLuwj2AOwoS3G
XXIVC3p2+jGPgiGG8SeAA12rIgPRdkdc8UQm6/ECSPeK2uJLV9TNpfh/mHAw8Y08ALIBWsjJOzss
J92eGjom+aJezFEKVRbibZ/WgFqOGOpNum1KIoBOSYuWMkYKckjkL1xqAX8dDb3jlumMZTpDAOgi
pmXl1mTOBQKw9s63g6uyqYE+baalOuMvUITjMBtxYK9U/8vFBdxhKXAdOA370sikNwpBCnh1PFP8
HONvCX/mYQ4k9HoKg814zccJY/E32G3m9f3D7JsBdA4rxtlf1MFsabiSwHNEssUnDmDCjY98W8fC
kUsOymBDeSapAOMxp0t+bUePSD/Sw7m5oSNaQBeiX50WqlelpoBtvY36YlbkFurC10/jcPRcC6fY
T18TiI6SKi16dpvEm69tCVIL+/jl3xws6N06sErLKGf9Egckf0s7sVnQajhtf7KFpu7E571ZTRK6
GwSNiBFCPshZG9+ick4V40ltukKetBA+d+1mQNnoy7Ro41Sz5a9H2sBdTfY4HxMg9h52JgBqzCd9
nLxjpCKknQ9ynko/cVou3mrU7bnTxqberONxZXeyOqVXSqtVFC4TDCpVpjXufa8CW9x0Pfy5vNVJ
KLie3Gs6lqvXWn66Uc6YVzdKAwAMgwH1drEAvKFXWDKvPUNdrQgKvuNjMRwZkjKzL7UkRLQkaAzw
oOEjz0Oxiib871JdNMJpWzrE+gWiutiPs8etFNiHZQ0cw7LcuubH+9+z5fqGIR5GLgPIEeCBmJRA
tamliHNc4yiOTaWn254VSQx7vYOTprSCmMMQ2EfvgZvhJ69RJwS9evM+Zg+uthrHfxW/svP+bmyn
9eVR6QJKVDwHZu4czeHjxZMtiCUS8hNnndMPDWjizwGyAbC5L0BbZszl+898UTaLZ8cUJ0D3dRMe
vyb113d4M7qZHFHsj3tPMmteMGmHI1s3kWQ7tUvL0uYd1nle6tak6OeSCBkfdWfNPpXd2IlRdFrX
dG5kvvod4ekc761D/U/Fonxa8D3Z+ace4KwscQ0H7gHRbzHAjlFWF8oLtbIgMI74YM1RtYGzkfNi
6FYs3DM0tUphst97WMDzLe+u8bfLutKgH3D6nmXnar7d+5k23fSQl0XJsQxEGWXfi4JFu5ZhsG5J
nt5wCoC4kpnACigkret9LnkLOVJTo136VvlrjrkU3+AaiVi9RU6K4kQH157BeHKirZuwUPREZcf6
hNf6n5RH+eNp0eSmvUb1aHivSIW+vCGSvuDwbpWnh4Rs2H7mXjPEi4hPB1Gq0QB2Xf8yMYmKe2H/
E4qpdmt4ZSYrPw5FHAAJMLSUWXGoUBpr4rJ3IHAzg1OckLd3JhnV3MmuBeh38PNoNLB0grm70/Om
HfHI6X2xs0bOSJtEs7pVnhDMw81GmHc4FmUEQ6zAyxuW0WHQa++7Fz1L60FQjRN3tqsPol9uSqPc
AWvKFmFD3kvU13J0n/HU3Mudc2fuvFfu82ohKRC7fq3FqoeauNc5Gyi8qJar7/XgJFaA623A0UBG
USa7zfYsgPA0+kja1BWcUVALZodxaLGA19Aib+VfU5djXrSNGNBYQp6XRzQvNxGAC46cib4Mw2DW
Fv1hCxsakp2f+flRqoT1kC1JCCuMCbqvIGH6BmDM+Jmld21oc7/pKw3ePMZ1cL9/5Hk9LG3Asamr
p8gJgt2BVYdzpvJkCzMDpVA8B+ajUWT2h7vCm9Vdr1uy8nqiYw6j+G3o7+NqRNfHp8v4LkwCw+IK
HwQvOzVMSelIBnCRcPpfvmbB96vDH5FRsdEDblv9UgoKZJtJo5yiSx0mq50vAbXE0kS9g4Kwunkf
7gBrUCAdDBMc6zoflMoFHMXYlKsn9qpiRiAmxMIZWw+Wt/NJ++kdcwMAltC9+G/wq+hHja9qKwJ0
pequW0vRnvP7VcV8PGzLKXyWr6kX0Hs0hdiAVVIIl6YAmUlUROWaTihGpCPehqCpZ6r4GVG/y11u
EpYVrvViYuWkO/NzJFYEMUWEFvdwUHv8DyuryWWRZmdwGZu9nkzAy3gEF1MzGWrcGxQRwypfWKg6
26lqmZhygQKNmDtuW5M0rPUDe9wyFJ4kVvfwXTtuuaMVLKcYIOLHAU3/1rVurn0jgUceycNvY61a
ddg4gCoApWj2sIOzLg+uDT6SNtl4PRaTS/HCgpwpKliI6WPv4rou27Ao6CFO1OyO6zgVwBJKwPcJ
plcgj3SxNyiiUJVa9bLvnc+D5oQ5xWFbTkmpWvyUfHFY9SSTWsGWL1hY/zKywYxWW2l8JyHK7rSF
wfDtA5nNIjIBRehxw7sDS4Ds7ilwGPBp3CWHb0fPSScb+6hLkShOqtfn9pchp2rgcP9PPJGZXmLP
Zobg0iRJRzpOEMO1f2/maHV5AKycqKLMuR50RcOFb3QYfIkUkUPRahtMjM+HA7AoEnWmE9j+Ukiq
PFWyAfBM27EXic8nJQqVkqGkKYJ4r/SsJgJjHxEdbxFYe9aPRE7+1UWQ4vVWkNHZ/vsdYcGLLS1/
0AmTCWP4B1Hs0m4xU28lTJtOLZ05IgiYbsfrz5XirV6lugSr9IiPdQDnwnVP4OdnOHOmnmOlX95S
mu2uNDWH2Hrc1NHrIfWm5RqpKoTwCmTyaR9t5SNvK9FBqlHOSon3FAbR7p6fy7RUDwXDvwHeJEoT
ckHnuRFrHrayWhVXvTxW/W9thWKwrLWpL/8/n5wO3/yiGA0U5X/hWgWPDFCc9oQI/TG1gn3SeX8C
CSRcYQOEhKavKvGWGbPgS/dlLZsao+rq4yPXQuz08Gt6i9ywBqpXcPUaE4qBXETKee4yg4rqNZv5
xM/szcyj3IZa/1qOBcHsmBcDve8Nqcr0k13VVrE8XydkdHOZqCKSk20hPivx+bStTgwifXb9r/kB
tMjD0y3Vsft9KbpBnZvB2b33AkCHOYYABPZ2CYznqSKQCp0kA7jjK7bf3nd3p7q1E6IVxWaASsZ7
Y32kORNVx9BQpbShwxIhZGfDbSmAKOgOWlhpbpglbbtuIcx2BMu+1omaNS8+V0Vy/ygzsDuGdHhe
KzhWDcb4pkxTlSf3FWE5kZtQM8z06bQM0Z17ttHLuTC2eLF0osb2Hf/m6uNsD4wGxu98MGr03sGD
zUR2SQ0vxO4imK+c8bkEeoBOMCEX+Mu/lPIRpWRKNSwqF/hEsDEZDCc5V9XSE6AUwPkUwP24XUgb
ZgzUBn6D0slwZzNAMVKAgpDQo+YDLadL+IeawcylNs8y/mz/qSbY5ygdRVArraP8LYLk4Y0mwJoK
SIhDj4A9yYLnqjh2cnIz7rRSAlsl4axbgQGV+n5D93FQcrXm3Ix2Wx4uspnxo0qlwUk+9XZtWBeX
3/YEdgdK1xK3iDhfCTnDNp4Kq3L7HHYKYLJ5tX8UaGKKIVKr+9FBD/BRdU6UOBXblBhCDfT1T6d8
BLmB6cjToCajDay9WIytckqpT4k8HIYc1995bLm7vfOylkUMcei1593rRoxEemlL7TxUOQnGCGYZ
/ejQxPfv6iEy3sKRk8ttKN9U3nX9W6znQVuyWsji89Seetj2YjSYJytRZm+l8BH2vY+uRC0YU55A
H7b/2fA3L30yyP41T0iHcFecauY5dEomYV6gtUsNJWS3/FLyS0z6OV/mwupLj+gWn+0Dk5vP1VSz
RtqaRDpdwBm07vqbMQHaySIclZ2hurbcjYkQuroUqrTqA0ev4BB0UzTNeIM2uCYE0vxoZsKLr3nN
K+7HI7MY5oslwNM3G18Gj7MBiw5CgVoGzrPsCJMA1ibj920T/JqhUSuXlaE0gex9BAIS1+2tNpnz
s9eNC/S/r0r2kYC03C+3c8d+3Y3PoZlWp0WDMt5bp4lyzUZFDMMpPMnr4FvX1dBpVawzsI9rg80a
6QrO7X0EtdyIja7jtBVkfDASaNen9w8H8XZ1VzUaHwI+sbrWYeNm2OxI6ZS4KhUNxFh3Mtsaee74
W0rJCqu60xfQeFW+9HhSEiqXiFID8aIzgm0l/5vawqLzyCsAHf9V1QFAYP234nQI7EM/qR5c2Pd1
w/+4zSMN2d3PkfqEWm7jw1wfkQzPBQHK7L1XHM6OPFjwUubXb4P6aBjUy9kdRXEUiOJmjwP7YwUU
E6BPqk5D8iKztOpRLHN0F62F1ARTei4GMP/K+YDqm4mQ3acU0UuO2/VZ4qe5L8k8KJzYoBa9SdUS
sSsN97gsHV/4Pu1Ce4EDKiEIde01vxp8CRGS6pScKKPdT9sUk7QgP8mSJUTHTfRXZ5Cwk01Zi4ZG
r6hkXsrvHJ75ZyUJP7FFJd5Q3VkAcSH6JbBbNSL/8oI5LqBPcgcAJLOZOBoPglGQ5u+nuU8aPK9h
HmLkUqjdMCQu1vGm/EfzCG4TZg6IhzNQsS7yqIDUl6czf6pf+6HO2YEAfGVzEYwms4GcZ7em/w2q
U5Jp9dzCAr0N1Yk7V7/B9RrvjZofMkLFjJq6+xz4CmrcfKpV7AbIoMWWw+V9CqgJc4ZOPleRrC9W
I6RlxzRdDXA5hKkqDchFD5a38QuCld66nHsSU/cGE/m4KbeD80u3nWtFp9rLebzrXdOS9RvpU5SZ
5SRKXpRDFcem8/vZk0oW0GZPS9y1EJC0HLzQFVtam0CmRmDbc08Wgdb0eSreSJnK4sG1/aN4kv9p
C4OnSQBlrnRurm0LlBEzoHCXjtzuB9ITOMSECs5PhGKJdPntCpxYdF/CMLe8Q4Qcyo4go2TyDItE
x4m3fSWSZhbTKODnCodMYxjwefKyM0rfu7Istwilut0jpFm4UAQa+DGdfeaOoSSzmZdSdGm2v2yN
FrW8xDCwdjSAqYoI+aHaNbNikyHRbXgmeG7s0CAO4tYyUOiO+2xNCcUVr0lndZ0ZAlkBc23aCfoG
QMPjFjwUIuzsHZkcvM0w2dHXnrDeeB1jGIbPyGQwzcmylyFfhLsPHpTQBpBElreuKwrulroZ3Dkb
YzH7vd6tXbx/vTuC1FBU9xuyDYw7EkuoI4wDnhhlS5m9ynAmMxEes1pKp4A8imNCPBsWvP5zinvv
ucn3EmqxFxnAn6bc5RbiAd6XEr1/+EUOQRZ4sKXaJ7IO/2mkgTxx0WtXI+OoYiLLuVuMjyHVvLsO
UXEtKKuOqxJSl+ONNsdFmcHhOEYOUDN0asjTX+nCy1yK3qKxsyHu7hOoR4qp1Q0ZELmk4QFbaNHp
MVQxzuKHafJ4dm5nP+iu/TeGBm89z5Xtr++EH95wpAgu1EGsaD324DNPtTKHAjfKVOrA9BgdEm4T
EzdiAVg/MdMhgqJtO7HPAxDA8PV0HojN5qB/cfe1GT9K3JMhRRYr0rZ2HTzXdWzi1L3PNJ0oP1V4
NESDgJNbb1OpJ5UQGjZDZ9FvUBJyEM1M//y+WrQPBxxjaXbYjCajN5giKIgREJowpgUibVd/rwHX
4pvTzfn14aim4HbIEUDSMkv79WPEUKuwp+VeX95bgRXSL6h10+MaeTt7wsywcs5FscFZ6wP1EfCk
qUWHNpMxCZfnbnh6qmPmmeOc9K3g4rtDGzEEtjXahCXrb8ErPndu3BS6oOcHSWSogpECbn67f2NZ
S1IzE7YaAKIN5IWvzBIUv5z2xPLMMvTi9D/Tbb/DFx0a9u6fJrQuez0NYrs8V7HQCWMwr9dlWRp7
ua+XMPIWB7HGq3LCkxB0WjLM1JUoviCAmLjyZzlJ2skymXNW6DbslY65tD97lbwVWVimsF70HIvM
i+o0Th8nxnCUWFCGa+tDWfS4dS2xmSM/nEzlHjXciPv68ON6gYmPKGVUysyHjpsyddDxo43/cWAR
b7MC5svNnwvK+BoRHB8dbZobmAJYN+XFakNzZwN4eUMlKoOFZs3m1UoZ2IcVc79pEc29dAEUfx21
8cnCY+CexIjU09T6Dwhqz+IiN4OjrwAJ1+jplRs4tsGw2OgdzIvzAAFSTPj0/k8sInprJrw4CDML
f03L3MN0eTIhlTqQ5hqQBff89xA8jSrH159aPZA/WjJv9tB2fMHKikdHVMbETbGZuE5RGDQ2SZ+e
9/bmtGxR+9tmZRRhkZ1A720OuhRPWzDy7HD9zcoJVf4iUZkV/JtO+cKaT77Rr9VIRndRPh4wWGfj
Ln752vY274Us1AqPjYY+0X8lStqmFKTsQjqXvtRH3oaegYe3VTHXTlsi7bPBlp/b7/xP0nAyrLWK
LmixbbKJuWyaRChvJQpbMGNl+iUdnSCm71Tcl4uI1hLQHa+ZW3G+6HK9+CnZ8vZWMTrbjWx/VN/1
Gu+oMiHMfU82Rm0JWVUtsz8OoBjM3kw4u4FhbzLRSxotp7Lt6wydSepnCJqEREGaI74nb4c8ioA5
Totib0zIk/5aiG6QrwG3KhYZ7f5NUtEgW8U1ZvRQRPlteMwUKHZSeBFNSumTh3f7s8ulBr0F0k8G
1kstCeAIwPKFCAp8o18ziJViUgo2nebkseokmII+4jXDMTPsiOHf648KNvR0x6TAVN0XcPp3Vi4l
Yrv8jcog2nj3EpEtKiJTTRtJzn4LElDQdEm9TAzU6gHG3kibXuckPe1Uxoc8tK/+hSZ8QpGSfZsz
Qsl5pw2eLmujwUV6O0C3OHKhjoGietnWVpAP/VtxN1/RKsKEhmEy/UVPAoZf8BrqaOUi1MlzX3Fq
mvyw3Sdacqjag26/l9Hy3emNdmf76H5NvUUK16vSQyE1tmV1vHWnRB6GvwS0loYIVr/x80uhgRrD
druqK+Vw67ZMur4Ll5rCvlOZgSg9AIY1B07Ktl5cT/7UFz8Mymkj8oDzoG3L8WOOHyXuk1qfyHmi
B99J3PiSsV5BzabAdGpA7Gn6V6TWPBRnwLmsoCnCV1UhKtxMRznrTDR+IKI7tz33rOaHXSfP0Y+O
n0X3XCjZfHC6wfLEXWFUWUZCSi513xxj1sPWZSQSdGz4qPbCAYnwECPqYvmo/ZC88otYOQnS+TxH
GJNvCa0lBW8r1G9l82VKEwNcwVQ/MPRoFY3Ai57WLj+ojZaZcDGUsQpK9vlwRSkN7+OADJkCeBmO
y8MI3tNvIJ4v+Db1EFJXh6GALArzj/nioarhgRImgX58JSyGGB5LERXGx8D5keOkVDUqspvuMzsg
F87vNYxmZoq54v4Rsi0RsVhpQBeIN7QiRVP15Cit0Owu3UEydM2ODnaCnM5Bfbmi9C21+pNNVtHA
no6aWMb8q73gLIqKJCs45jL4TXOj4KzqCyVARYZE/2+qANSrxjv7aMOwDwLV6WZC3pxMPLiXeD8p
UrjBMBo57xIMQNKdGxHBOiA8HDg6UzCBBrhWxqeq+ugzOkJuITpz9Xjc+bgnkWKV+o3WW89vNVwK
nVzuIn/VOMQodMThp7oCi3EevoZXFvIWkuJpg110+MuUzzW7nSWx+siw1vjXgcRudtWj940OCD/h
5KBbAQAaDXyYHn131t1DwvBy9RRGAQLESM6u6HrsDb8s9YVOd3cjhGG3ZKuiN5F9S73xv9R92jqB
Vox5rEtVFknuhOsGvIIHcYF+Ck9Tc64IMqSougQmcFK6KbhAR3EcEJHoRAucJ6J2GeMnSALoQGiD
dkKoC7ESyk5cO+8dJL3vyti8AFcXeX6X86CbXqJA5abLQ/ww3HV2mdgS6zc/9pCN27chFtJXj1gP
3zptQyhJfCWw1UrtV2NVyHzeiBVJZ7DJj5WeqburKlnvoWCesRtmRxzj9MLpsZiEF1X0Wy4MZyhh
q1+7UrLbii4eGX0tvyoPAUozSW/abdxIyPOTKo3BsGJfN8eHNefj05vc5zfzdFFR1aLpZ2hCNfBB
DJYsy1r6VkTbNhCb30MOiZaifEiWHERSqZxGM0z7n2q2DfDTGWVqsQ+Kv9oHLFeHGMfWiek9Uxi4
lrDJbWhhtG+N7yTOmdDqVczflwJ1OnN8823YiryJbYnyUJcg8lV1chK+2zWLz/Kv9KXR3YV1b3ow
dmiDiejCdOAhP6g0KxXewHeE1FoBpU64+QcP3PxAZs8PsllJEFE199p7R/emVSDJkScGICp5Ux62
XwKJIxcbFatbppuJSwGkGfk=
`pragma protect end_protected
