// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:35 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
aAR9WMSED30gtgg/2Mm1J/WBzFzKVzrOqqJn8xhsFpCkSvoZtkGM9XfvAA+JwQ8c
pyJUXhe14p08D1wBVcPpNLH73jwoHwG1BkmngizDLc0mxwOAhIOYhnmhimjoPLYZ
EuzW8k8sYFlg/w3C/hYE9tUMf5BNut3ssccR2epI0cs=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 35152)
cBqV0LAvHSepGi7SvTVKwEwkRqzu76M6hZIwFQPN0k+u6QoZwZS6VccDn23GJkDl
dv64dGvg7zlrri1UZxM6b/IsRUgoPsA8E/oUQMWsz82YFW0EI32LGnZzgD9H2V7f
mRVzcU9ggMKoenHwcv37d/WtERSeYY45dAZNaw6xNyvnEZhGFVGV/2YIzMBvXjxq
StGDnHBDuVaFfjKGLQzFaFR3umgtyo+CAN4kZyEdTNuct3zeJCcAqjDiSMkZv9vC
6ZduZXKiFnxPLduptSE9ETWVg33MZacuhHoyx+/f7glhpGRht1A3fZfg/C+X1Buq
0f5cSyWWWZCvzTpBmBX5mz4Xxg7D4RQol86GMVtTazkgHdUlVngG7Ss0IVvczrpm
jHFh6w+AvIp2Wt4IJmhN57eRHhQU6yrVOvZapvw5K+GXV1nOQ3TIppWX0vB7VSbc
Feb+3Ji9g9EGRYBvOlodIwUPH9xcFadUyclHni3o48lsbLlEmty6pXzW5t/y0zUG
Re110DNrTZQ8ZikHZieaemSBUlYRkjRHEp/Plo/ipg3muXGG0I7Pp1XkARJfHee9
gSpv7N0PuTUukuJa47BLyQREnr7BA7Nf1MdRzOXtdjo9P3pqQhhh/l392vyMfPIb
ncHW/KFO7OhKB3w3oz2F0ly5ohhODR/f7nkD+REXBkixpBLq5+bVPIRppcxz9QzX
bk0ML9NN8RCVhV6/GUraPNCrWY8/0VfZpd1rWgLKjCNvK3NAEpPkbW/mhe+M/SzQ
8KnlfnG3IQ5rjbxCaQjlcHvtSQ8fLaD4mqWdaMNwq5FQN2UHl6DtKpAta/BE8Zg3
2Yi9a098RafbxCZiWpANnhbOdz+zAE+5/v4X++bq6eXcKrkM/QFPnZ7z9XAh48n0
CHg1AoGyVui7MPi/G6kKnprB8uGK2V6sxdpQxmFDEK7BXuWCtXccw3qr8i42EAbW
P0Uf6jV9/Bao9DD3I40hbFFru3hv6lI+Y4fDP9aLKBKXcoZiDNzyjTn6RpcRRxlo
d9UfU125SuSm0JB303bPgzsnSpLcUnoh3HC+68DaZ2vDgwzE9pqlgtrEXfwcGEap
z5AmjSGM2nIY+t8VtZXdw9ephk8i2VSUzlRlGnuwHWyj5f70tSd6r+L0DEd4KZiy
ZjDAC20rosqsNfF+UPPZLA/pzYFkUyAa/1pU0nrS5rRgT6Oof/Y1iUu2C+OpvHf2
LyVIfaO/13vpPhLPLda0IJrEPchRHg6e462g4FPw7staQrewAof8FER0TTgj/R4k
j+K7MVYPTPnY32xfTtqSqnQ5wiCFtHFx3uATeIxrfksFm6CZGGn2hnq3qrun7gRR
rLx7H0bEUz9jnkKXGQC04BXVomDUBsqjHPbMs+xwo7JBN4H4NBcF3LznlUvANKMt
Xn+yJ2dQkkItqE0WmghwgvJBEbUju3+dD9kbGlkkyoQTLgpukyna7gEKS39+GiT/
Aw347pduFWX5pLz3Duu3LTeg+UMWuWIfvjv5on8TP3ntkoRxYQq2rn+Jg8IW3Ies
GSFsMV2NExfOO5xY4w/5yvwJE7CDcAIkgT8xStwSz3eY04RRYtrOdABzfgXMRggw
6uhrSwkhoN5x6flYq5njfqda1xpID0hyo1QEG1nftvPHKx7Y4ZKZuDnUzz3tJ+W7
iYUpwOW1hIAW8XopEJzVx6cu++VsnU/PboJYWka9IWy3YebmEVMHi+4lOkYwnuyB
w49Oc1ZHtMHDa0LPXcVSmmp0CQFIAEuT+VBdVYv09DxzFOjJdD6oj3+3JEoFvPTZ
RaWDm/+2Br2saTVeYRONzviLTdZ/Z/w0z8sAhfQi3G7X8++HXkL/Z9k3kAndpqG+
mSGMBXUeWuduL5ytzohqzgOcBJ8tWzfOF2TEvvosH1zk8Z+FPG3lTx4JlstKyfHC
oGf4ROkE4Pk6mtgYMUUdEBsqJzEkY/2+9Feftphplc/1kkmKTuVgo5Brp7sVN1Lx
ib11XwyFtLY3hulF0QhBbAEMya531YXg8WXZtqCb+IG2Cs1W8cjRwrP+NEkMO/5G
ZZ7D8WgKEw5wyn/bzIl71xh+2ub4NjOWjVGZD0774vyKhS0l0Wuy/5/wRIdO67YM
T9AkBkzthA/qfke6f4JaqyYC0h/d4TL4NNZTv4Q8OULKufigDNvIrCJEowe641Df
oDuYwegk5f40RHSaqyTWQ/R1gXS175BB9ouZDAiYCbZvjZh9SjIYDHSsVqrNEVZO
fsAM3Qj6yKgljV5ZXY+vmVtyju2wjS3C9rR2zLiI/6sDn4qE3eSBnTI8IfFpV50a
z3fD516297M0JOVCmjJR5j2SNDJZSwD5GWwKUhAtOT01ZNdp702Jw2Dj1Y6LdQ8w
WpPuxU6ecJ3zxn3cqSa/3QSnn8UJLkuThB3gsA1QkDbOrFoY2X3kRkMsoyVjZ+M9
R1WeuoQowQPprTZuCYnxacghyxOdmu8FpKl3886pKCcBFwu4GW1rFNTdJbEQXHsG
T4I5y0X6HMNZZabSdFYhE9BTkzDDHCtiu8XpmUjiQPiyUSP9MLzSYyR93+J2NIlk
tbhbyXXzEEXvAnEIJ2tMV2AKzfMleRk5iQrYgV8Gb7Xy6LsF9h/mevElV3on9m7z
dhE8nQ2QIDot4n9tQ9IOUEY8dQd5hyqS8ICYgoxQXrM04bmb2hfxDGrCoYG75XjV
7gdxiZ1/8aG1OPcBZ1f5pKHib69X8DK2CsabAche+2kd9HJUwofg6LijaG5hWxL1
GHZJPxchvp9B2wN1OdAX7o1f5oprzHdfeGhdR+MGGQdhuZdotuQEDkjRvoc2yIIj
3TV5gy5MddF1YyA7zTAYL7zM4N9SF5vvCJ7tEJCuN/i8oZPVPkvYuCFwh77gZFSK
Qq/lH463lh8K0dkO7H9Sl54kVLFBHB7Tl9Np9MzbtLIOpHyTmHjhF2a60XzetauK
cdp6ypdDBiyqgXFI9nk8/C2MrFvpc2xLhyMZ1C8m1KdT9+VtfqxPgVM2tVOJ0C55
Xi3YSBv/nKZjOZK4Zuc600I7ydHiFi9NUfDiE1fhV1rQfKEiDgveYjoJxJpL0ACz
s5Id1MZJTsPDJGnhM/rbljYXjvGIF5IYURUSL/8hbt/dbIPuNBwuvl22ANF9s6q/
I/2fIGjddDtJnjl2X7kJaYXAWl/Q37nTamL/VPtpABUkEWIGCHcw7rhq93Agooso
Ov4pZY+R/Wvkg/qCzhFTTw68j5tvidEK/Ow+WTRClWjg4XDfIenM5SWnQbLxyk56
e7odPYXlnII/B5DRkJ+1v0f3vMMQzRJ8bko/bMHmnFg7/PVTd/EGtv6R/e6i6udf
SbQTy23FMQNlrHqKEwVV9BBpeKgrrSCSxmH7YyLoSfro6n94T74yAR8hH+b/AJiP
pzkdNIgtAY5ABrcLWhFLXOC2Qau0XRVy21RBHwv3h3BPaPLewJmNYqjH1AM9O/co
xdJA18XRCTxooXsklOQmJizCgedEqhJ0+N57CxAOUKdL+x12xGVFXcwVoqZTkRsB
vQ0jCpUW2Q3Atou9Rd51r8R04UiIy5a8Acqr7w3dgEniJFMW916iQj1eS3guVws3
xeJgR7tlAUh9Rx3ZH2Al20ny+YtekjaQLmHnYrrCNPpyzL9/K3SyDIvSQqP38/d5
I7xa9g9piW7LuShmUTED0lftXfEFgr+qKlOrAN5AzKW1f77Xugb2B28LdxCn28N2
8huh9ltm35xUGuZgkKAHJC/0PW6v/yAXrzvoYLbOCBBpta4qAdZOZ6acPVEYk0hz
zX67XT2oL8bDIHBkgms9eCdv6fRQxtYpqGMfi5tWo1w1Hfbej1iX6Jko36tVFMAc
P5EpCWe58cpYw4WEG3s+uH/5qvFKamyN/6/6CrB6k/ouruvkzZmG9hkCdjjYLSO7
4P32CpRSoKsaTu4aRzhWnvoZeigIN8rvyqacn7T6UYTFXkv2eR7LqATEGbh4o7Ac
UQO1xx+dFrREyFY7M5t+RTIGhHVg0opB44jP3AApU5NTKbAi32jsNgOmalc7hE9q
8Lde/SPQy/74fPWtXwWpEhvRIWOfelSW7y6a8f5J+aZQu17jwjHuwt8Lk+hOgfiM
6Avd1CPegvXX4dJa4bx9uVOKYdsBBfOA/8jTVqNayDUn8r/3RADoI/HsJwhLd8+j
2YNrcQoXlvs0ddz/i8eOXvzs6Nx9cUnGI9Cv9hI917v6IFvQDn/mHfqtK/OJF6Sj
H06THSbgTn6X5P95t2fHpfarBjEEpn7Y7BZugrFCTOM3silhS2B4mQP2kpIM8Yyt
KA6GKu5EOayFX5TiX+ZZN4vltMrmRHukVMEx3KgA0c8RB5n49SZF3rNZdCFb7HMN
Wlx31KVW9n7QPiChHhVZeVU+R/SWOqyu1C1q8A0hz1qb/CIp7a81Q9ULMyOvjiW+
47jSZP/IL+DF6xci4At/22ZwxfaVPm2FICNVRWb/4OrbjrJT8h3pPmVrGMtH/oVb
b2OZsB+V1dD8udZMAop4Xl1Xx0Avi74GD4XTZ2s77VWnZ4pCQ/eeoHJalRKVmX6N
eu2Qbkdp5vOxkeyR0k+NL534u3KNuA7mYx/mkBZ/wLjMt26kxCndzjzh3Ikj3VMe
b53jYV3Bt7nBvF3ngJtsH3xGgf/lNJZ029tdh1rTS3roX9Z3XI5W7wgMviAumCk4
mYWtsX5cLObZw7IaOPFS+bsr9x3zQ3Dwz6X+EXelAyn1mJbMrxrLWO1Zfrept3EW
PcisHEt458hIS5qli5E/jW1wyb9F2obD8aFybZkZoUw/B4WsG3eTKsjy235xrlhS
QrvYwvnzxGpd27DLgG55kLMm3mV7hY1NCF0dxipFTzHhTeGxEJp0jKBLhQzLOnKQ
o4g1KAZ3lWZhwuvpXaAZHDLokCzCvF439QFDHbpHNRPbMybJgGiCO36+aOMO5BML
4GAwhfDCJ/MCpBVB8KNA6qqge0vOZr8QHyOkJa4+G4VQWV2meiKPq+eY15u8TY8Q
wV1K6zrF3lyeRWXZxtJ0sscqIWmwfXSoUf2ysn9zr7WOiG7B0MEQbgVOkvXSqSJ9
xMk579RVt2IRt55/O5c2HIWgqecTG7ixJyJWWgn/wrsdTvIHcYRjCqYnHdYZRi8o
MZqYEJb4kY88orXNkw5oMEbhl0jzlCvqaW3G1D87cfG4gl1iab9f1a6729xxNnw6
a5RrQOVG/MdgJ2Qoxj8w1b5T+bEhIsaqyHbKs5kI28+LTQE/Pq3Kxrt2U7vA45+4
bflTqC+Rlx2nBacZej1iEmvUSztvrwlH1SXW0OblyXpsEXCPMMjB0hmugFxsLDEC
svtipudloWUNBPBO0kx9kklQy6eL0eltl8U8ZLqpnme9p9u3Db375UXgiqphL+Gs
nO05TmMgkNqEWd3IoL0HbaGklCygxvv1CJDqyLVnlcie9V75wDIGUN1q9XZck5Nt
qr29vE5NnMB/jaGm+bSu/FCPYzA13x2OdY+YTS0WpQHwtVL98feMbdz9iZvbr6Wm
9KeDyplct3U319AG3ApS1Elgy7Zxo/eeYc0vbjJ9GU1mONHs0CKlPrkJqeMz1IqD
GqOpKvxetRIqNqCZrs/0mpu4bnNXRsbVs0MsV+LGE3yUvH+T8PIP4nyV3+XvOarj
NzMKUf0ZvVa37xMlON+ODhMW/xqOFt3LtPfwYR0LB0H0HumuCFGVfQBpTnLjB0Ir
y0r2YlaRlciUujCbST80gx87SimBxGN7Sl49Npwapp70Qp2DKKdcu3wlehzXMZih
03+i/N5LOd7mcJYChrLsJaTKC1zK8p0DYzBRdDQsu7GGig+uIQqses5e76sNsifJ
NHjJQm/IPER6XGFfR8OD6kC1czpMWAozKrLK6ueDGwMULNLQ08G9+nIlyQRCKnKo
SSa6sgCPp2W7HfEdBiIJ5QMx6/XSbByv0Z7pJDwxHbdpSE/zbemi44dWgiomp7nR
IBlBt78BmAjNVBjiUnLITYnBRlZ0y0CJyi273OhH9yBrE1SAu0IdEhSQLf269qPJ
gZRelYzQ5SgEqLIfAO2JyfYCDPKCc3q6dR3Cd4e7+f9CbNBOuqAPTzP2f8UFtJME
0P8zzQcDBvfkYUfQAvyMXMRDE69cP4niA7Vb+PryFhaMDkk+BWCFejmLi6D1ay5z
c9PW1K8jISYZMQmnpi1rOaRlp8grOiuiY3Woz2Zj3gyfORNj43SU9pmC91oAgV4A
vMDBo2i4dv4AfKfpfBMeSsy42Jc/HrXv7WdpqA5+gSSScbYn/llvT60pcvZHJ4k8
D61QqwuSPbnHsUhWqajh5YMzbfOlM2ECy351N63S1/OALDyJxWyRClZjoVsh2jkz
1zZ6RGSIQ6zEtlY+uTpjE1YV4mFcxtXfX8hBuN56Da0ksx0N4gS3IWFyzPTCgOly
9OvZGMwGmd+U3B6g4uSn74My4b/ykzpJm3sVwyo911T1iYjdkgsNJAVTEc0ymOt5
tBqyiA5Lwz5q4Kxipnh83ri8SXUZ5yBt3ec9DPdyk6NHjNkMtJqHbzzxmQIbhoq9
KUgyelK8zEkWJfA5hcmD9TK16QUwynX3gUJ2Op3cIMOG2Za2FOzQbta65qewasB3
CtY3zVqi936tmMZqEb98RPat7FZRMKTwzHyl7BYl7Q5Vx8DPaFID8I+IE1p+bEap
u5QwdGtg5aG0F+CN7VWXlJb+LGA5rU9+Pz+jGgvNENN1RbUFnkHMrJRdiD0MuuEM
z2cSH064V4jsMTUyA83zaMzCOFZCKoBtXPNYLhu0LJ15MQB0vXhI/4c+RQTxBjbs
nhoxRN1IItpIXZhM8zw2IJC/mKEzzn6+fwdQdZmSRZL/Pbs4etP+SXplburw8zb7
2fjxE504rHY1yAuEt4rFUvyF+Beid/kl22bnBOn0uCODbTfbT7mdNOPTg9MjCkuQ
lTG8lyXyvOg1fmGywAa3MVZGuK6rudf+pjM8tmrgjw0iP3BWq5oNT1mkMjiWmour
JJU1wHJcAs39n3S0DjcS2pvO0m7dq3MHyxPXPFbNbuK28QY0QWnALblQEy4zKfPv
p1AVJKVm1jRpPYOChmiF5u1HxHbXeo+FjD61BuOMJdp02SaxgX/ijFbHRiYp+Fr0
lESqChShJLIKNsVvzyhYNKsTYMgf+HIO+jOYbQIDwheUfmhjdrqt9lLSXXu9X+nm
B2lkBdXsbhfF8NJeKlAePErks/g1GLsn4FZRyeEyPeN68UWyfzFslG99hqOxV8KJ
KZbb0tf7HsNHwb9fYQdzKR9rFXk3/JcH3n9jenOCWExeoh0SiEAwJprMeo6aPXSC
pwLW+zcOzYXjYXsba8/PWeNk/OYSMzw+iz5TTYy2zI/XiBgmkkR+HqEidqrFdHU0
3LQGGJ+n1BCBeNRo/eKsLzxFQu4dfYzKRuY4Rm/ba7R/jqgVr8Gx2IBfwUyMYqWn
K52iAI1rjvZgk9pyol679CUkBpXUYG3Ew0QrkPeTOgLL4OX0+V2ud0QG1l4YdXWc
rBo8gse5nXOIUM1kDN4vX8Raegpcv47Z626sUU7cSrflmtSw1H+hK0IvJhK8kpNz
Yi9uhcyb/VL7gcassrM6Vr2yHNtJYforvlN4lq0A5387B3c8PGmGxKHJ6uDuPN6l
gG8RtclhfBPlkG2TjxxMQqFZ8WNpxmpKENh9Pg97nNS2DLXUcUp1IhZhzvLiEE/Y
fcHaURrF5IRGLh9h2rYgNGNnw0cTTzw91SwjFe1AZ8tcDgnxRr8XdYO4JJlKU9Oj
Ro9D7lOwTmEVwGcf5ykAee8RN/MrYwAN98XjIf2rELqQYUZRV9qffeOoIvE4HaoN
dwfP7z06L8oyUn/psvn81ddLYgPljxWXl2fHUut3fkt4pKy3X4/uBUheytHf3UkP
ZVjpRoJaOXA90+54npyN/7g9aoKMPdFkm6kPmGK8Dc0mG3anxGdcMreu2mcHQaz7
A9oTAEvt4dDwsi6eel7sgv5LsBkuWvXNLzAdPM+4ymy3u3RHzq8sQcZyV6NrxOP/
g0rNLwNxUXqcX9eCzwaqwUl8M31Iz43NBeSnZ46ycE+WghiSd0edN1Sse4Whgmrv
/S4zg4fkOBV7df5G0xhT7//L4Shlebt6ThZ0kjL1nHDLpsQoaY8j20/pQEOGSGCK
Egi4lnjCHhpyCrPd1KLpTw/sRfU+rQsy7SoXiY5m83ofFJvtZ9s/D2xTP6q3Q72T
RWy+SZ9I5hFU4QRVFQuniMVXKMqMnoyhsf+9FtW/QBVZSUiiHVnQKJXpZKMAlek3
Gx1fO92jkeoNT0Cs6AcAmnuXKiZsu6G3rAfMo9FFhO6PAA0nQ144eEvXOI9BNn/O
ZBpS3gn+WXqju8GERPQfXb23kukhX4MBnEURcvnzwYGfrWXA9b5c6ufS344DTNfK
xndnunXcf0UxghHJOfe7FiOK/opDFVcHOjcIOGNbH0M+USKpVM0VJlhZFtMtvpvX
pQ8Ysq+8qlJGwwRGLFLRSzB4yEXqd5/9FLzmuOw0nXedSGB8LQOAPRvj2oQazclA
Xlk3WLdR66cuwWRRfErQ4b7WopdSfjNNDLWoYXz2/gMbwE6dEi8G4GifYKWrxJss
zDbl6jTN/t0ZpKPp+bP488Ap+3HVMfqJIaLkSfui3Y6HYYYBkPuOPIPEFFPFbEY3
gOuIyb2PId88Jw3TpvWGNg/YBLxDrJOPfu9k6dzx2OtqK2TOSuhoteq3G0bSfGzc
ah+jfYkANhBf2jTOLLxNCo1AIYOAOT9M30R+JFtHGiDShBPQrzjmk2TJUBni7T/5
kzpGZC4fOOdiMQMJPYZ/jEu7ANaIhLBqyNE7AfkjQLFKb6X6UtjLAa0NXbAofXF9
jCeZMTHhV3cxSHIW3CZ7XoybZiu3YijiNaXKPxt2btlpubfBhzuNN5sqrygC/bt1
ZxRyvk2Yy8HaaF1QyhioRgAljtS4us2/nfjU30+ya7j+lWmleae4hg3/8bxz1mOZ
oZ4erDBlje7ZYPM3Ff8IO3ttV19vg0tcoyR3MWCZcMwU65GzIdZfpY32n3NarDjU
qypueu2CLWl/1VMTRjwg8Wq6Z3LxyFT+a9EVchU/7VvfNSXfPelvvxYlx2PkPCg5
jb2V+T/uAjG6KWRCpO7r9lIArSftWiLgf/RgsQ3hTplUayN2K8anlJSWPdOjP0dL
wjcBZ3CA+D7KKw6AnvpO11oXUNRkiSZ6GSojrNP+AbqL2Mo5n1SLjXv6mYcuihvB
faNNA1GZO5BLbdNl5drvgJh4RexGMxF0ghvW1fT3OYWbx6CD0WT5gP62MqjCnedy
JEy7SxCXnpjQVBDfMXqkMH+N8gbtjMS1aPjbSuFSEIwwPqF0nZ6sUq2B8DuiZLDY
/mlcUZ0jLL8458/UPK2TS3zUNP92qFJjaakYpS503D96nsIEg5zLnKjQucPwY9PE
bv14VtiQxCyBSxAl/1HTwFSxciHAzvFCxxWIfUQukEab1gc9RzNmPgiaGGazQhss
lOSlc1HdmGElrEZd1Qx+AEPGsC6pkqNykwzb0xPHtHsZJYGUChWDCtKQ7z19ORcG
sqLaWkR1Pq8idpXmERSab7pOQ8GMAbCLb8njjgVZiPBOd6pcjNC45ZPDz+vJ8Uga
jQPLDkxKAhAIwZzqpe4C0RzGQaQj7YRmFIjAoPKcbQe3WezCOP4GSmxy7mzdM1Ud
UcqBrWjPpv2mnRRpr5rzGpQOqyEoHex7JcHnNWa4aQR9R7XbcHyBkXmChkXV8mYe
AmM44P8LNnFV/nUfw8zk6uuUUfaBFORVZdrnSr1Ohk3yTQ0FLabUE/wzNL3KT4fr
DmHc9ZJXfPmvwtQnS6I9pJ7jSmAH5yUB/2i6zV1xtEHBhmlAcrC2ftAFPx3yIPh+
JyWvtLloQ7RmcnALOzStY8wKJLW6yeqSFagQE3bLdTx8dyaBRHHsKo5iKL6Ep2gR
RBxQ3ncKPY9CFPKwLH5frdhfeFZl8ryCOmLGetmyC3LLGD6I4JXGsFGD2I/QhZZ0
dJBLuwwaWWoQqx3Q56wRfA/UkywtbXZJxlv5d4ESArpkFgjzGyjU/xZA7JiH4Odq
Rw9Hl9gq/blbYXtlitcFD54i78k5JQS8mElM8+nE5BtDWLqERGFqfIjpCIaNgEgl
g5B76ndL5wtmm9+dmALP2ey8rd+5LnIJqz/4+VWm09x4sXUoAloXl1RC9KUj+ArE
WtOfI+YI0vGDRogUKWqb8H+OR7vWPrCWEythC33htqv+58kpjo7IBZ+B1zEMUW4H
mVzZhGrEggHtOe0jtJMv0Kaagq78JIvyxE11TmWqSEg0NGilxILWg+bbHvT6SvUP
AJptDoDDHq/tnL/LPSHZhi/7Bg+Q4eKv9OZMz1eRtYbRhtc7NMyByyK5HWGZapWz
4pvmGaxG5LklI+uN9HFFOOOF4PwU0lZa/yzQRpKSUvb1C9DH4F96M/4XV221NHht
oa8ZUZ9ZIiOyW8vGYIUS+5Bc1kYVYfW9jZHIlalUtLLb1B2N3u5X7JSsJ4zHYyBW
EQwGwfnKVl8GfKDrytXsmCn5Jl0lJfaUvSeG9B3oPGivxm2UY8IeflQzGqram2KZ
wNNF0qhZrLTDVyQCA7TGh/7SsBfxaCVg0KsoFEPQhJRiaD63M9TmG98cz5urbauT
yj1CnsU0SoCdqJp6n6ibiyd2ps5fjIZzuCpT4M0JTXtciUTu9w+UxEel49LEwYBg
k9YCRftZ46oxlqA0cOYs5EIegfZVwyB3ib44NYfI/mP8K4QxAYCVPaWfeop0a95H
F6tcSzjrlBXZYUNarmhqGy/SqPUnddGvZCnpKxVjnlzYY/2DmNeQqxqfo3XD4PMd
TVVdovCLtu3dGl4zFVT426ZbRAS19pV92SMNeLjb5I4/x63R9nciB7O7hXsR3mRJ
+Xev48Bv+QZ4Cc59tivasPwFyBEicJe0wbrg5y6ShJmk75c1uVUvbmDSdl62Vg45
/2KdIFn2R6YpdvNR6dK+w+CHeGywMZivlKhm1vNuU0MBf9zkgOPGJwGwMEA2hGcN
GiAlUnEjbzX2mAUcvy/YZVLMA1cHeOzo1hHMyK+JZ1fYbazX7UJf+vDexalQFVcl
nDXlHfYb4cf9dKRgAVd1j3A9rsJ/3mEdPp2qbYugo0LBrU/UgaaVjAwthbJ33jDB
X1lppER8Rx1iTVlOZjUNhK9JmJFMUL3sNbd8jtOfm3h4ExqOXa0pgkZrHia/yjN2
aOCrYDGg37VcGMH1nDA10arNcv69ivtQk3hOWLorOy5DjdueEABGVkF3wkXLuZmA
r1n7w6sUMNCzNG8lpw5TxTwtOlHpfhcmdj+gOFJR+8e3eBB742WFMN9/++x7rk+B
4lQX9aLcJNyvPx18gUmKzWMPLmERUvgvn6Nfb6klsZMdg77Pjm4Q0/dIzptWbAj6
Tf2E5uoeVFswv+T3x0T7mcHm6H1dC82gPOo8fYnIwsQubEIM5NVRtRgu1BeymiPr
JErwqCcC2UD7jHjskUC+huDGOUBKLhvnza5u0YmOtU3c9NDLczoNsU7Gr6DZMJgi
FxZ9zKxRcrhcqbFvduNnj9EX8qDAwK3J6bZlovShgXMuSiPDDw6gKzr88eUY9wZW
T30amBoIP552Qb8yqX8w3U/A/xPtF8gULjVdX2T07ly7mZr2IMFDmC4CKMfyMPqQ
Qc389n4A7Pd+2R0E6veoQqE1nun77eTnGpCR00O9qnpUedHq+bEaOKxsifwF631S
p2kF6SU9WRO+awye76cuCw10Wptl8GysrmBbtwvSR51yhD6mMB4nP30uDG66xAp5
wSQk9lcEmRqaIjrlA3k7i7VRpNHK5hRw61TJJrWg/EXqfpna44q/8CgdYzJzrsGz
oy0+pVWvI8inDsQiykuXSu/6VD7i6xzkXaTb29FKBcqenobx+W34Gf2351c3JrfF
DOe6qEkwYTWzwWLVlR6pcDq1Tc7lTbQzsfrBc52Zl9cCubvmWhHtaaK2RrHiJrz9
DlUMYoyrHwUWSOgn6uIkNSpoi4uOzZNGOdji+arUe9pFVwy0ipYznPdUBr2nPSqv
qsbuZhaJamiUUuqBRC/xe4MPgON/NlpLX2pD8TKM/rtiqV8IzfIdCeKoQJUl6jei
jEo0xaNruQ8Dr8LhAhUa94Nh68QCojOerX9dDRWUVRY6WZo3oc4Bjotxhhp5rMza
0ANvZPQ9V3j7rD6iNisg+7LZLPzAXkv3rsdJM2ffALRdt0vjyEPsJU6MUXOiuVzD
7sbiTCDNE/tqDVPLc0Y11BbaDGP4wdvu1hbArgx41kMjnLzPnu7PcePy4xOBTcRX
Mhgsxngo3FyQUndKaNi18aRx9wPnZcl7VkNr5oZYFX+bVk96gBjTIjS/Z2VPoqX6
NKrvIJVxLZND1WSYUI5QAVzjm0tCiphKFucPsbTXhRQDnDJGA730dPHTrDyye4YD
DQRjWsBAi6lk1eOU6bse+/KBLGnsvtBpxTKq3KEo5K1qpzodYYdq5WBzucU6eh8t
aleT7khZXYQIKL0yXCb7O23/y7SksQC9Rt4mC6/FRAraN0wwBSAHBwIomJmr94Ob
hzQ1VKGY6WtU8SNe+ytUottU4yrwuFl7Ht0P7JIE17xgTWjbV3CI8DhEtYZNgyTS
ulAkf89/DAg1kUHoQyxAKH7s1ENKXNo4NRCj3235gEdtNG5xNMuqax7ODVNGlxUf
NT/pP24X8saT4AYpPn7Zb9OZW/sDFYr6xxFGDnDe3fKXisvKvuSSt9rp7ynhTU/7
/5IDC+zlk5lu9TnMNBBz/ofWDkcTvrjXcK+7Nxvmigvwn3+z1dCXC6tQTSNtpNhV
jePOaMSonyFv1bHgWHZ6OFBxtn12sj/7n/9oGJw7XAEjTArstXW943NgA+OIypdt
XvdBngDXfjrG1XufV9TVZVKCo6YB0T1TQzE5GxzuRslYxZ1t66DXDZ6fj2tEiCDB
IG6NaN7wy1+nEhXsLynTlHSrpDk+ITzkX3/8eA2vP7VDYJgQGQLYvEFOYdfEsaY0
mvltDsmgfYrR0CTLM2vlDbUhQaV9Stsg1Bfnlb9EYvN0ZuzXc1pxP27tt/0xrcek
YJGr0dMbIpDFleufYVzQjZNCC83A5zb/BrQzYuH+qVO6qlRq+Fg+RaefOKFUCaBE
lRRjmpSoZCs5OIDwtSF0Kl8vmFnv2IFcm5jMfyz2VZkwdQEfmdc4uqHRSe9euzG4
UvBNtnvDGx+UooVXEWsIXGUJYzEXbX9X/Kog4PZoVlPcUpSn22OXBZvpg8Ggilf7
81s/Q4ZnFa9MuUww3swZQlH/2C+gQ2Ep2cXiaxQNifPTzBXlJiL98H7KJaFWTTQz
Me9fznUlaTDqiWQNC0r7DO1Ls4957aFkIv57briZ1lVfJh9pBkvB1KrhQErLSQ3c
gjIdgx0LmhwhEQIPRQt/FlzSyU2rclFgA9OeUWJ6XddJjz+yndMORWI+gr/z1UCR
3fmDqAz+LfQv+Xy8ZugZwr38oQZE+T+lbZYZrNtG7xKfBWNmJXFrijfAWFKuTov/
ilNM2F3J5xm/PPWNQrw+Pb/u7M2ZlVLHw/ZoocG9rvypX9lpDtcFSIwLUuxD91LB
YXTnImX3r+oQcRRFJdGXeJiVwFx4tDPKRfg0brZr6WzTpoW5EaDxf4eXyaPv8xr1
xBA4D4VhTICJARAMRWKACie17M6sLGhJkfESy3FKyxjl9bK8wMzMjPakyJHQ0aYR
j1SGSZ1zfhGC+vwukm2Kz86vmZc2YXFrFp2fNc10yRIX7fKkLEsiPaWAMtOw++dw
njw2rv53yIDP+KgOfsPrWsAMcZWq4wXekP4K6/ZwxR/NGSnZPqMtUaiIQNpyxZNA
MAZEyqCM3Gfn4S5ljGUZxuADLmNPqdqRUbwk7IJu40HjS4Zg2U8jmf9o4QkPtGtB
Y8Bhm5wlks+LtldSwlGe5fYMX3+dT+h610K1FNE3iRe6Ez8O5RDa2cDGgX+oFZxM
nZ2g0ZYkiIRPeIRZPFVxiHw6fd6IjsQYgTKm3OhGwPTqcEFt2PDE4daoWOI2VkAS
ndGZI/3Fm92hH4+m/+U1xgPU3EgRvz+RTJi2JVqduUpvTFQ60Jh2d4hGY6y1io9+
bYcaHj7Et1EHJzLYFqkxux+Mc2GKo3KAcvdYpiUnZDajnaV4iQmsVwWAuOHcGmi5
64FayPpxplY5q3s/xtsF/V2qleqeYlpJpjZ1n25bhLfA9QPzkCFOUuV/P7hc9e+P
EbCwVd8Skpb7S7EYbip93Gf/tjBJtFGnYnLP0Uw2KVX2iWMxxh64J87aiunAD2B7
e9dgLce/o0KdIAGZzs79YEfFzOq354pNsXEELPCxz4zKpUz/ZrWj1w23I6qWfGgH
tFUxT99OA7dtJ1zrwBAWbiTJJn/iG1XBqJ378JfrOocdH2kPrJHB65YSGw6ss/az
LcTbfTfLwaIDz7t69MhzyCUXkVVk0ciXCv85uFX1+rwLunD9iZr7zTBzqLsK1fXL
CuyrhbxbCJ2+0gJ3HDQBeC4pkH4CXZ1feyW1N0/1CSwTfdbw6DblaIGd/SRjCrvT
4lxhdPmCRx6Rbejgtp6E9jh0rSCL0Bh6gBAAfJLKY2cIXCcQZlZlAZ5nBMrwZWMX
u44NUZfdiyR5PA8dQ7taiiZYbRJ6vlW7gBMTQJ83wblYWmVxU1wrZ52q/IQVsI5N
YPL3v6KCJRu9k5yS82aL/AzRWg48euqu76eWuIepCtdhrYPuxH2e9UymR7loo/pz
MFkxJ+LR762Jn2Vq3lirp6tBJtLFno9t28LsH/3ahT3pmpiiltDsYU3a5ini+Pu3
zOAb2mFqY5P0lRHMTmrFhICWgqNqbRuVLfxAV0ok1lJsBIYV/OLNUjjjqrCi0TQI
uDhxLCQ/IguRAxJT7IlPS/kd2a5QXXjrpqly/GjPCGkMLKgJzgCY65IPd7RIV2F4
9U3BlRgBi6U0mDrM1VcYZtG3Qk+W35YKaOyl//v1/C1AyncwVrDBjZ8TfCTfT+ax
4kdeUcPuInAe+6yEj9NkAy0lCMHCsWtBeM+JqSGEjt3HtBl1aDxQbLRDvpPsJSav
mbgeziX8vT0AREUvqdn0o5DPzbiME/MaJg3LCteQp+R+RxuD0EkxWWpOqv03m8qL
MXzVQbyY7jlugfxk0wk6TZWDwu0oTeUs02hwWdnQo1ZEDXEjECDEJKitqa+VzRrt
Pwjh/TanKEOdw/NYz3WAXgzWEaBWGYncxcxjPqZ6gTF/FK7+FVfg4cfCm3YB+f79
LGUv35xOD4A2kiSBWQ/YJ+9L0tlcrGiyakEEsKmXSSP7+GQrt/cQMaLhuIqvj2h1
k3rPI3GHuRCqcQn8VXTUxbh3y1owhbKhKiA3BD8RrfYNQbJ9X8tBnkX0qyWtmG5j
JiiTwbjez8NRC0OxZ+uw0TXp3Z06NYlZj9uhVlE/VfU2t+Ay6ErtO5zl5m4Ve9Ix
F+CiwyEBWG7mI5tyqQGHunpRuhyh9osOS75qmpuppUS3kA4wbNbnXdqvGdkq1Tr4
d6gKHtG2ZkAXbG5JUnPB78fLmkNw0q+xyQsauIv74O5NEx9FE/B393EEzDv3bjl2
+D0PMmn6Unh8BqidK+RwVXUpQSnl+5OGAant2PkR097MXhVbYQvfdwB/WfTEryPg
+/jq0UESicju2ALpIAmXcH4JXzBtdgO/uxDI7rEOnF38XY0HYVvpBDQkfWESZ1du
u6jDywjScup/b+YVQW/4E0pN1kTlpO6vhEhkMPxD5t582mlLDCGjS95DjR9pzWNa
SPgo8m8EIah6vWA199uiQoXwyo7MllCzYX6bgDxoADu45mWCnQ2YJxeHe16BFtn8
DOpAODkI4XoGjb8BgW2c9n5YsyUMzohQrdGEAaIkSV0J2zQ0Y5IEW+P5kDPq5MVX
u/sCIGefRp5MQHsirUdIsSKi/E4pf2Ty1yL+Uj9R48LiLd4/u8h/vw9Mri6rX4hG
md7SDMZhL88pNYQoWWllQn4gHWSYUtgmUYq8GUHTZ/LmVkOmejTu9Lo9Y+R6aY0p
7yS29LULh6s5IreXaMt7jODDTgogrwKnI4Y3BVdWt01fpUPiuriek+9eH+Pyxy5o
UIIe1mvcIa324ihQFYLbeHrpoV1+fSLNblPd6Rna+ZXdRmu0rZe2ZpOlI4wzXYD8
uFQdOWbu9Z9aY8tE1f6rfaRk7XkZEd6JyyMKXGDIM18CVCsAdYDR7Ay1fy0dOEcq
dvZAR11350n1rwWnIVIlZ8Ec00NW9X38hXRFVXxXLtZ5Op7juQ7qKbB/T+RNH+OC
GQdhgtDLHrOfw2XMpIQXMpeoZUakJclsSUFKrck6IQ97Pfd+GzFw576Bt8CexMdQ
NCwDA6SUseQ0A1slOMBxu0RONV6K86uL8/dRqQFBnrj29CirXTz+13QNvkXjD38B
UHUx2Ze0ozbKNqsmEnE47K3oQYOXyc9cSFVsp7vFmvsHSuWUwtTSe2LcJN0tRGpS
RV3SdAyFQCgwzw56sqYlsYfj7UIdFqw8wanQMYJnuloez5zYFayS/SfGLaATxoMZ
QSNWLR/BfqiS1DLsrte75/oJXbvsEYHv7laP0AO8EbppdaVUGpIlmL6ATMKUP/dj
Sp1oD/X75/5gyu+9Vb6WMGOdrDNjX71pBxi2lEmxzUKkKJWB/+QpP0WTWMlVj0bI
s/cVV6npdePEtagWDVZEEYSCGGl7Jgw80HCfaLJJNVi8Jhw4M3WzXhRD9JUHFrOl
BomHjUPeJAfFef3LS2zOJ0COGghA+N1zVHzz41Wu4860+/lvNJL3eQD4XrpVDRYO
fdvcGm11Hcpx/tcxxSfwjIJreg9UHQOStKSApkX26yKYHsrc4+DG27aBMbo+5KBC
VhKbV2ygRYoBoedB+KeJCLXTWvSMmRxchmcK6P2iZX8IUnvKAl1xfZ5NLdyMYltB
dMeZWfbA+kxPqeSnoICW4oMISQsWgTiQcDtmly/xEc6QAPW8Ip5Kk5xL7/GI50fk
GxI0LhRwirB69/dg3H9Ku7F604b1UhdWLWLeVINGpsEZ0Jx7pHB+ffoO2u9Ih8XF
5mVuEvRmYhVEuiR8B3Cn+c4L1yK9J05ZPYmkOfQSpLjhQ7Y29Z5cin84wb0WfQFj
0jjQKbPrK27X3tPbsBXqwtjekm5tr6b2YBPpyf/3bLfpMvXuyMIPrO3KJrg8aP6/
DkAGIMUEL7NoURR6cs8wj77mgDvRQp151spJYANBLiChdWy6wGNdDaaHFukCd2Qk
FureHzEQjXm1Yq9htQNv3qqtPusd5JjPEg6e8jH2VvRCHUa4rwA6pcWqP/YSMU5v
7hvqf3nUPuQpaj87bHoIp00YfnisH4Z6ckN335Z/cHIrDaMCcFm6BUhoPdsWfiuX
V/1YERqVGDOZ4GuyVVkMfpmPT84ToFGFONUtCiTLf3zkqjBTC6M39jiZ+A5rA5x1
PmpEacHT4HdzCFLBrs7UkXfffYUGfabE1vEnMmhvM4983Sgf1kbda6q9m/Y9HMCa
DxZ32Od+Cj3khIm7twER8667qOwgYF/SOSSWW8nB85BMWlLwZ0MuNmLlq6S7NuMT
8FaCUFWD7q7AJp9evUe77c4ORY+f9nXarxreC6Bn7nBi4P7z5684hQqxEWdGE621
n5ayd+npvr9pun01oG0dwBefE5p4XNWxdH4b+dkCK7wqkRCEtm2oSXYkBWWrZrfq
M7XfGW8sTPh0Wdv2YBkcaLjQ46Lwr4wPADSBIBL7QD2JjOt5VrH+M5Y0PN/eITNQ
ojKiic0XYoAef/pIE0Oy9z1lYhb8OZ6mbW2xv+exOlpiFUWf4AsEWQe2MYbibmOX
+rocSvzxYsvfXUiUyOKPXpOXR5eDSzRctXjAxfF++YBgAJJNN8nu0qv4qHOjPeYs
2DwJ1U/E4RfTDgfGedBUGwweHVNJkcXqwn5WdsKem8PoLHP4qd9A88q/Ax0UBBi2
NSO+c+H7G9dgrXfSP5SnXOsKxo1G8u12n52mj3e1gTulWATPuVsH6/R8F6onE1C1
Bkf6ZMpgQ3FmCRhR6eiiNViVUrEFlMiUXlFeNST8tcDogzk7mR3qtr4mc7TuM2Gs
mmBZ+rjFGdk8pjQjrV8QDFyOiTmad8ZGiyfwuecfPWNuBVHKFqPLZAMogNQhwiVI
sagLl/D+T281ykJnewPy1jSjknG91Bo2hyV3NuFdo/MMlXO1ZlMuNU5kXYAruZQf
QZQ8EnESXaJ6S14DHqHfBqzYDJSq1smt1+klKJKfcRiVxTu0rpPLUjcH0vD8eM7M
3KGw+RP0gYjTk6G+yHmGcbSVXkWO0U1fguPYVrf6/RhsdMZUsNWTuAjinJc3oE7b
sGUJ+5hM49WsLnUMsuMWkAtY1OLGGLigpKn8gsT8FPdJ7/XR2K/X1oVnZAJWMJZx
Xx/Ccs8FfBhrV+M41ySHrM9Ocu7Mw5poC0OiXZUedO0U1f0b0HgkfPlZK/jenyx2
3XTEjvr8Y146g2/BfGRakuSLNN19oiGENP55f7PIb1TpeMHWkda15yMa85302Y/U
UhR6JlQOj5TNkLFEyaXru86J5TXEvoVT16dVNIXeFqQYw5r+IB6dCvHEr+7r9jeN
lmhZw+uQAOVpxJYsUumYisf7D7gxeZPIHgcUJ5ji6QRljG/XTSkT/CE/sulUbQLq
dY1CBJXGDiwHzEoR9MHNyOMMIh5Lrtnw3UgkmPX5LD0lgWeYz6M+B4uhYt31+8Qy
DURfVxfgYoJ57OMo75xHFgJTl+FHE52Kbmkh3SptZ4k/HKir7rgBc8e61lbe69V5
AqcO32ScNX4+H2keSkkM+/E4DJmEf2U7M+p9ZqyCD3T4QeS7hTqfYqfcUB1XlhmX
xM0lsAwK8JUpMWzpG8UTjSI1oLP8jy8+0SwWcz8R3lAoJb56vgDq23x3Ba6Gq3Ge
KnYcf2Jx0WbNT90RWHLU+mBf6+GyqtW22Da83OzLhfGs6mjVk928gNW30ZCq+upR
EO3vR6GfTddakvdssVKtJH4PVYi7coMGjs/H1iThZvFpIal3UNpBeCkS6aznutA4
fnlgo2/vP6BOZ3jgdBGX460TQ37flGbNo+TDvt038Jtef/J8QDna4ApUPZECf9ab
IcyymPJBgMurP6u6DbviK/bkZBvuzwVrPd+ExZtfFE90QLPkYa3EWcndBuJmpnuc
fSm5lKJAiDDA5K97cBa2tQgFJLEZIhaFVhujoJPQAuNS/qpYBeHiZjYlGIM38i2l
9zCt+WOCAHqs4jiCnP2FqYSnP/kW9xrsEcIMp9pClM0pxsxWNIAGyLxIspEkd1m0
gJz+7G/CruibD9qQZtkLRCzBkyoPbS3k3p3punStRPfKpORORljmY/54d/VWb9Tt
FK1nnh73o/CNFnrdNfpdAL3goO/oUMAQsqUW30rSC9ljwfd0QboL5XNgPTRBfNMI
2qNlAvywSOkRIT464wHElDBihrhmWVRHWbXQCS8TcX1Fpn5joKC/qMiM05tgWDb6
QVafvxabcPnc9x+Oy43ORWUAu/59sK4PihmU4LVrJ3aO0+vqcptIt2TXCRqhiq1z
NUYm8vhDnKWkKzTFwpiJsG6UIctn3vWITy6Stkq4X8ETJKb51c1WNP1q+6/OgiXd
HFS2kOJVc5613l1gO1NM0g436L+StBeGZLQCtFcaDglwDbnqiSdrafn1cyZbqCoz
rbuRDA4rqdt0kBVwgrdkEVdQrAJ7KLkTqpAEDaUQG9UvpenjHkgG3UdrI+4jaMQv
QYr2PECCtzK7q2ZLhk1m/6XLY98sfbfrwy04GPu4aK+CUWv2+zinobMKfCLVMchy
D2Ank6Hx2AVpLCYwVUwFcX19shZi60s7wWVHQzOlyslAaLqRlRQmg2iwPqIH9F+/
T6GmQHFkF460Gfr4C7ZZ/4qTzpPKnRQ98NjEW8kEYwDyZFkFN0CNRtyBZuyP/HcA
Lipcv6J1GFVUPvQuw2ZDNQT3/2iKigEwbOU4lQhB7X1IpFrlv3nCCjs8kQRIfKP9
FVMv37zcAP2TrNhexrXYN+DLJCcx85wJcvTf4o5WIX50ppJxBQJ+W97gDHZ99Eec
NUbvS4pOTWmRintueAfdjsWpVEEja6AAR6SIn4KZHYMhn0T2O5kiyQDCylCZAmy9
HLuBeXvdHqVFFz87D/DxsUE3EnCpH7cFmSAzG9QubZDgM+31YPMshrBtsqxD9oOk
DxRRtBH5Gm74dybJf1+6VqeqMka5aZ4O90htwBBYcAIn4u1i3DG7OX2rAuFWkS0D
pJ/CyfSNPwlYQpy/kz+EMBdX1qbSAXU6tokjp85CN9GyutLBDU4U82TH1wFwQX8F
RN5AkOuvqqHdbjDtc8HS1ck9F3YTaI4vvvtx1GICFO3kPVYJD4aBwZNkTKMiwNH0
Yy1zfAMjbJ8gPEGqNtO5VP0J5xdBwUMDqCaLnosGhlZm+u9mQvxbIUsMP1uRv3qs
CHUGLe2RwUtQwICHot/qLDdlRQgsdzyF6f2E8jfuNSf9m45bUfbv3wxTNVqzOjZ1
AponKjVHPJaHpPUhP5aqyWVIgLI8vlEfH7UDacKPZrH8vXo1jOOPQvx4a/8o9gGO
ppXorEHOf/oiH+bQu5nKN36/BOUfoQn5/xiPCov1TklIlEu8s+5DKqDEO4/YidxI
F3Sk14+qDr39L3lQ1hyZN9zTJUgXeIPEWVIm8DggH9nOCTk7PpYwBdiLid+ZnAKK
hBELLikZeSGoB3PD6V59MyCfzMDvSGqgvNkI02itdDehWTw2G0Ki1zB48oxYrVDy
tymiOq+EXK3ySXuCZHRR5qhMmn9EQ0ZLsPE62rHJ1MoTkVNbCWZMg7sHiZT49EEC
ueQ6KGlw5HYdWYxHaw/k544a3wOqCwJr5dAp/ESEd/Y4jgxysT05lp8MTO6O6zGS
5GlpSO6GWpiXUAKoTu/hREPKpc4891WmgQ2ZVesgLWo2mG+zG+eHc+74JaFYM/a9
DkyI54zlzGB9uCYfXpsXqzunOjlrONLgwy75kT6d0CAdrFaR54+4JMaCxzAza1PH
dwLIyLuJgwHsReH7Xbab0WGTIS3ugdzSQL/bzaATgROFu3fjfv7IKWCy3fUBF3dS
H/AAYVhTdR6gGT9WXrzAaEkf/MjAD0SrHReS2HsF23M1yKEaioLldTOBqn+NTpa+
LTts+0y2To3rNeNJpJG0ILf7rXaZf0ICXnKhJY5Mt2Y1aFVAJpHj1vI1ynpl2X3b
2wm6+ZsBRCdpK6JKvvKWeUmbvMivZGLRpJzI8pmvsus30EEWBRk91aknxR56avVl
MxiAIaX5jaMectGrZHdLleZY6kVdQzxCZqhvDNYCtxFlzR32PoXP+L107iVB2Sk+
/qjNnRNv4f83ZvuoUIPr4/aK+IJFrR3nhhFdDLRSH8U6Se1sCAOGHcJCc8RjPV1o
NeWZulCkYxMkyJMfbpB4zot7rhmGYVNgI1m/9emzROr3eCyk2t6Dp3iJx7OMU4co
9DfIMZXDgw1fHUkiLits2yxVfw92bpVA9W/jbA7KDaOEuXxgp3H6DZwtZnwzLoqo
gGXM+XzkbpeFQd45R+nO7CkwwtckVEbHHSu3wHpeBXSH3IJ2JdPheE0kYvbhT7MI
3Ms9x+hlIPaNJMAocDspBGm+O2hjMstCW6lC3PA0BxDuL/hsU5U5pQaWCxH2Zy6T
ZjuBEx/ClwnvQV1jHtF4/j7mTzVtQcJQT7WxGX8gjp62O2peTxYrRKrDJylfACTf
5F6FB9K9ttRP57jZ5JuEJIprIdLyhk15Izt9vRI2qZSiGllR/TCY94PPtXt3Hj/U
poHt3BB3UJ7jXcbjC3ANqnCxuE2N82XGeg+Rd6+X4yHXQPMGi9LtwLpDetYvWtWr
uLMgGjm0nqtF0b7Fxq8RczTtX1bM+mmG0WCmDkXYALwzOJvDMoxaIi6EfV+YxmT5
V1PLadLTZlC8ioBETAdBzKQzvTJGwsGNv+femeYHTb8rXHkBOcrAcpHjWsQyTwaU
UHPqDw9pfYS7hGK3lLeS7GLT6UAkF0QePzLu0z5dII65+kHi/3BzMhKBwWPpm6k/
EUXqTC2ntXRlFviEg1+98aZpullzlw1hA4wdkWXp/YY/Ivd8TGJKJWfuB6umAtj1
6yct7b0hSYJ57AzpTzpumQoaWs1pgC1AoNlGFcqSN6ryXoMZW+71pXtnEdf0VNc9
crxCLbbGyYhJ6R/2lOZbl2f72vqoVOnEEZKFulXLjESfBEwbgSVBMDqr7dp5oPQf
Q+Xb8li3xIoI7f++fvYsakuPlC7TExwzflibsdfp9NjLXhB8q13byJvS1IlcsoeU
j/OAhD4ZKGh4QuUqQPiYDHQinys0sNxYe+ccr7qIMhVyU0aBahOOho/wlWD9cX9D
75C3/MglEMqEpJKteDtHBOG/jCNsTKcciZPEFz0DC6b0L7rdixKYIo9/B3FEhBsv
MP9kLCxwFNWWJV03hQt8A1bqu17m8vdplh7L7z/MYEb02aPLOg8An/X+a+U81f2s
0xCcC23U25dmvNO6IV5x0tO8KerbkhoVP/ORJ4FKyiPBX2xzOOK32eEdScrfeO95
Y3EQ+tj5kyG7v//9br9c/Ak7h+EodrBCL1VoRJtbDoxqqNrLqymP2Bb4Lm9d/IBg
YzvKt34Q5wAcpoT3Nc2ZkCkrd6ZpOhQLihq+8QaSFNQ6TTX03ao79bAefWjdp9I+
w0Ogvm9WqXro4gZ9HPoH/UQbnGJZNcS/gI0F1/ghPBweAGAjXlotMFReWDB0U5R9
8fn1Xv6VUOramUu/bui0Rncv/4gvz/bAV/XxznmM44t22yCc/7IbheNQa99HbfXY
iEvIWo6gJUNaSgN6fm4s+IwkZ42OmSzsUL4B1pFnO+e3oO5V1GrkkTSa+y32um/C
xyyzrT3mEw8IU5yDwYhO6qFXsRmJhvRupjOKudB+90h3NbtmsDYLT/BOF76ZIrrg
rC38gverhzdMWWzMAmIS43cpXXjcfY7VzDGmpce0JJIRF+B4onsHSiGGbVBPJqjS
+OwVw/wq/IF4N/avKgFdxhlc8uRiaQDy+SX4QYh+wyJSfJDx9Zlm3O6iog3/6ney
xr7JwcrjJIEdpN7djEk0O0QA8gKL1KiwIJvFzUbPOXJC0Yn1tWk+wt6CRlQ55rZM
M1icdjpyDopjmwzfGtzpnFh6cW1ieEn5+a7YMTGhewzELJcrqx97Gx4AP6AqzMcX
YFXnhoGOPddqG6P8K1KQSkz6H338lQtBfKqRvubJm7FG7FIaIT3vkbZVCaLgmFpE
Xh8FBKbLq5ElReLOi/NJV+UroP2D9yRqjPfIy2l0y6V/mx4GRxqAhHFoMJ5C6jyL
1h/g/06TDs9qzGdjOQmxv8YltAwBTjGOEsXClWIxkW26MPeXHInct5YPdTTnM9ah
dcmEyR4w5/wZjwGraCf7b7RKGdd++/ggNXnwmwXzrJenCzGT2APd1HaHhZMViwMr
lCQ9EXUTd8TalnMF2MBLaD8qhJScmDHIcW+B6k7gkdphfdVQnIpV0oSFdsq3hNz+
IqWaeiG/aO25YSkaJvhCgnC2Dn5Hgim6O6wJhJ4mgpltap4hp/OUgrAThsnbgSnB
i626mOQgZTPrsAxNt4ONF+LvQw3kso1PflMAOQ34UtCAODbH/vdEg37DJlbejqPR
J/I0CaryEgFZjurhD5J4RpxlnfHxAdK/zCqADEv/1wz9LDYhlB1DfF6Zmi4EshYy
ZVf64/CD/1iCuq/7t1y+PduskfF2+l3yT9Sp2cF17uUywylu3rp+IlTsSWfdJD49
VlUDRgvfAvhsgAi6qVb/6jZix/L6Mc/kZ0QwCgMaJ6KHHO88wp+Mvd6Ntf1cmAmR
NPIJiKF8NUm8/uGkcyjUYf2sCaFmtE2RQjQxUAB91AvMxvmRA2usmi3HoPKTpOak
CHccYfH2olrcatqbz47J0uzYwYz6KRWTT/NyyDAjSYOozxPk++Sn9Nae1LLdkTYw
5xs+O+h4bUQ7+iXPMYicZkVHLmfvdbzM3LMgoSK1Z4hcAR7Nt/gekzLwKa39LElA
PcALM4zzqI+sV4hCJhM2T8EUi3pCbBV3bu4Zszj6EXN118G9NkIlOn3/+BA8baOb
tIciKYeHRYuY0196p35sqijre7UuQVpMe9Me+nkO/NRr276OvCcvTOdDgcv4tyrT
m1xpK4JSLAxIaJqCBoRzReFwU/FQ6BPU/b+LP59nzo0o7QzyIsqaEWlOz5x0g3Rp
U5lfvmokyeqz4h1T4QQUjeMo0ce/Ilr43HNe8h8W6CByGXXkJx9xDNzeX8DGlbPr
ikBeKXNNqiPYIdQyBL1o91/3iGOmBGPhXlVxHNjRWLYsvkG9qbsGnfVuCFB8sc/W
Pt66fOSmbM/QC2je5snufBRsS+zBDKpoQx+d7o/4ElM4e3ywuhpS65plD91Owos7
XMnaqhcLA3te8fsKIpzCcL9FEPGhftbRK319v90e+tGou9Z9x7aRjAlCbfmk9OYX
Q1TxSILmhdLiwVIveB0QN75C1jvOpmlaB0g1XIDUSoS/YhSO5TrD0kECkhoEmaOu
P04WdoK/emcAH++M128oWERs95dnS9t2NNodGguZqYTVJ3+jM3XLMxRP1nMruSjN
8OZKAbjqGsPVQqFqT3SOnCbH8x2TStTocBZ56BorqRIc8h9FZY1v4M4TtLJ14Kl7
qaSogNqWspm5NkeRkHbYT2KrTZHt1PyCL7NijPke1fhOjMJCLgU1Bh8qhneC53mD
GCA722AJLJixiyp7vDDIebp3UfDtObqHAmXvGO3FSCAxTa1F2iP31bslBkcHlrx9
RLv49veeEEfhOvHMnwHYyycDsrSBp4YTKPhxx2z+kJmVwaBk3I1pTaW2cns9XH4G
5vj7IaE06tVeB+K+dUY3TlY8aKWx+3lqXXQv2oniJPgkc9yE47FUpTX9v32xspTd
FpSgRXunr1U5yLPViN9NqgOYqpYyn8vBC7mJyfZRrvPkNE3jr58F+s1SMd9UTkGU
JFYB1p1Vr+QW0K+YkuU3uJJM4i9H86KJyPzx7hEvF5Yq/y22EXL+w3DywtsFvtsI
PFbovYefOthbFlWxNuCZyV5fIkbT5EvmqsKDu6Pszdev1DwTsDLGoe2lkdapF1Tp
rHPMUR23rNLq/zRYpDZ10sKxkRmZvC01uxifm5uC9X4+JgVZz8rUVtidZoQfW3rH
aDDX31BSpn1wGUOxh6zFX7PL+vMjRYKeT7AsnVOSGoZrPiseyiE/PKEI4ks1oup0
mcqJmSUjk26OUhoQQU7ee+rh1HPmk2MUz3eQs2OWnJXSUNIIeCkSiILFbfGOS6AP
WXfttrlT1vjAZk7pAVe5BSAVZlv0dezOyX1xdic+xcOxOv8D3VyGdwVMfXDM/oAe
QEG6MRRaG9CaEMtKeFROrkFb4/CkKaTln5pZ4yPezfA7jGWM9TiKeAoawZ4qev3W
QcwoeaRpbRJxJS/79BFZLfQ2qdtqqnUqnBZUSWTyz8Yo038s0edrMYVfH0hdB9Np
7zeZ7b7ej5VSgwqNTsuZSeZP9DQgwcbI3kZTWFwfeCGun2dQlFS0oti9f81T8ho2
gP/PhgNKLpswsJJA4ajXzQG/VCndHmYYL8eItoglSHVa6K4GNfTAoykP4eBfRThk
FOct8vr1TPOCFZnP3HiwAqeB8jt7mkDRXzEvkeMogV1ABJXr+flX83jIRr2IHhPY
vo0Ei5cCnA7764jpbB+LGySw5gLtyradOobx1qQG79u1ptSNmS3eDe7K1ZSbOAvd
jyRNPXG9Mwq5uKSXhf0K7Z6otmRzXBiuJhQNucjH2RI7bP5HT5WnJK2I1ZDH4cN8
YG+8KWbceEhRuCMmT2TMoWVSM9zumC8INbaEYmuW7ge+YBOwFp7Lac4dPu2SlUEX
sqG94FAbYD2ol6kDAlndB+83ovN8hbO1pS5QrsCLjRpq4chm2YQxFGhDmpYmxsq4
5M4LYhkwFwLaQg62YZA0Kkz8v4etev0cu0xSlMbhC6r99FotYPqI1zwkVWKf4ipd
mF+nMKhBOIn8UstVPsNRJYcAyNrBWEo3lTkoRmCphPMfi22zAmEkKTS9C36aKDhe
Yc3SK57UkYIMyV7yeg7HeAQHWG2Clhia0sUppXOfDsCOsgfGex7pWneasPWzbZMB
IDVKxxKjqLziTb3NfLoaBpiOFZwr4PR/6gGjfVmdG1sCakx6i3O9kDoj5MqPrVpS
OtIaGSWTki7AA6+RXEJaKBYrcXc8fe7QM+37IiMwH7R+EtQMzPWcfP44GL6IGtHL
YwzH3VxZNg+DjgbQ0InsYD8KRtluUisdnhVWkGyV+cuEHraJJvrzV8AuPenVcY90
NYDySgHUtmXH96zP3+t9Th+JPzK8pTZkdgwBzRsMCSondC3DQQMr94j8C6dqnsm5
clu+1K6DRvPyeKVfOkpcO//FKDPJAnARtcKt3/GK6zylqETUpS3lV2lZwMs1lkqs
CNDspmA7AkO7ZQsfwRYcyjGmdju0QR8fJ3GyZlpZPkgiHhU/CSFlvoCZRgO46GOA
S7im1urUiXnxmzikIGq41ohR6cjr+sArWa3SpvegXmfkxzJPfe3PHbbr4HWB+7XR
jbq4VdHgepssbm9gOeH05rFFwVLLDtsd+TD9NgmsVN/QGQ3c2MyXfz2wZlQ9XlXI
AL6GKB1JHXyfpeWZI826YsgFw1VCoNFRMFAdIyZSzsJp/W4aTOsLVkvBOqHdOUBq
FF65tu2Qzr//z/jZ7boiSFDRdI8V1UA386jRqkesFqIEe4AJYYeyJX9V6uLPkaJK
JtshVxfFsCS5oHYV9pihCEAnCcpJBcsF6/oLyPitO5zgIwVQCYBNF4q+253BskCU
YQICHRliU91ZWLrWfaUnZvVevH/gYrRkOw6iUMg37a4QGG6KZerM0i23Cxvqhjh1
3vW3b4Dy+i9/Jte3/ywal3FIInatTKgMt2K8dc6rONJjkqcslW2hmBEBQaziKYOc
qI17TpL/1GTYQOr0Lam5TTSpI5adcgyGQjrVvpKFigT0vyVgQpqTzlpPJ2QXOjLf
ombA1iCvFZy4uN1qpcj8+9NvtICqC/AUecXIcYUMmjE1X+CwUnvegsuceZVoSBZE
6/19vewNGJN9w1IMWn8v5Z+Nb788k/QlmLlsdKsHR9ZD25I18h2tf6tUToCBEWX9
oRsnWqzDuf27u75BLBjFtTesairk3muMZy8h3R8cse89k4EWHuulqY+KvSobykVw
UoU4kDMXQqtyj1IqTdESNw7oPIVSL3alnMUUxcrNXY7JSeW6xrpQ08uZF+1BAggl
EZQygR3K+Iqgr0czC+0OqOD4TnT/yHF0JYjfyYoU5eL0s+3aVUG6EyjReheRjIDD
vMyAo1jEw352DTZU2G2mNoLZdAxOo7fr3Gv7dsZ+2BEtSfW4FfPMZlaZqOor5yyC
Dr3aGrJFY46JQeO29GCsZ+pyza3fYfzvT9qBVt/216uWJkQ6pOrIt2bdeoIKxwJg
3kdb7MP/oeNgeWZ0vEtzkhofTGYdRErFCILtKNQAi60/SCHGGIKDO4MlbWO4+iLz
YJMiqrferXcDgZBndTH6VKP2EY6AJC7nC7heVVdEn+Uf2sq48EFWirz1mFK8m36y
1puifuIa2BppJHTn0TVkSa67h0KZL6wbmGChtVt4FzNh7B8/s57gPoO4TS1Oq1Hw
482WmWFyDQcKBOiPOCPLGk1Ga1aEbOIeNy/MfKwtIZxCUwlo5sGturxD54DaQuSg
uw0QqivJK/Jsb3Ak6cLCx1GzEK5HCKQtq1kVsKfP5JuOuKCwb4bFnjq0IZizxDzO
u9DmiMOmG22G+9g0W44mOxKZHQ5KlAqcpUD101YLXqTmRqN8JHRYfQ5uoC8zwYW5
7mZJHcANIxTj0lse7S3oZqzVZvvxxNpb2ncudBem9X8EH/e5/2gy4psbln/tmyMg
ndjPkYllI4hEruu3i3yE+iE42HOPJg6LgB4GhL44ivAVbkgfnU5umqcgsYtfqQSn
gCrdlJs2czhyigKfUnpj01+p1hnVlR8gHEW8/iBG/pmLj9A28Hd4l3gax073YcMU
fUiOWe7xG9+djlNihywW8E/uLOeHvPBxOKYSxW7ZBPs0yIyqLASgIwHKAV6YTDOi
HR36DviP1HL5CskqRX9Uq6m4X8DccQhkMZyWhoL2ReRvPcBik8xG5jYY64SglV2Q
pM1b8UZsekq/ZcjCRJOIUfLuoFol5jFS7C9da6lMXhmcoWN6daNwFI5LLEI2WyL/
aK2voH+ndK3QwKTqTNmcjq2gVsTAQTiPWczrHMT6dJkh9uEDjjPehLHDuWzoFJ2Q
gaQmYU2sFpvD+NeRSyNzHKDpOvGCehErMtXy13+HAaAoQnoo/DFtx0rmAJBkF7rX
TV8fFU2eG3OAqleB/TEyzoZgSfpF8PxjUaDTLqNyFdz1v8vsDtVpflWyOs5KOeqt
xnmj9CL+Zgj6iWmu/kwWRHF6o7U9bv7gyl5QuJSw4zM4UzK4QoXcK+NRZbPZiZYn
UXFm1J0td/K5plMKi2JmRIwAOKBAG0OmQ/zgobz6H+mM5HGmeop4rWm9ZxmbvnpM
8uP9R5Ml+QOI6O2lRQsvJ6RvR6Ko8AmbHPvf0SBNbGqH40ItGiWFmi4ZhNHnrCIU
MysMy+1SS5YGhm9t9S+Bn4mF7J2rii+MbpDPlrV0R8IwWqTGmERKa45vKKgujSXI
s9x5WZHrxtx8clgTv+NIyOn+gM4WUb8CO+NN8fUrfrxfs0Z2DlT3TUqtpI+5WQsU
BgVhVsQrsvx/SF9PkJnI4nVhWuENq4B5NGQoddDU9RVIV3g8eMMt/oUl/ctz0NpQ
QXqZsE9xfGqxLPngy34FHFnchJTTpMEczavf5KMMG2LF68hswH3n8mO6qtKsFfkI
cJW5OsLnnFA1WWDq67d7QhvmLc6TvKC/GqLRzPFDtsiEQUORBOYbdfGNp6NVvNs8
8j+ZbX5WmZOpQNEDSkLeIWWWUfbAE5RF21tV4lTdYDxTneJ3STwCAIljl/7o5/vG
LaXHHL0gCp5DCDiVyDwW05yZ7yPcxS/ZkszmYm5JDorjSdR7l2vfZzyRHIrURi4A
GY0P+8+KsFsLb8jJ5tqnqABql/UbjdLvNWO8HFRVZRv1P3P9swI+QFks8GZ7j0Cs
AEOYAeb4CCPg6Th8IXtoID8QH7OqhcxKb+s4oxsdArN9k6xbpY3K0zpEUua3L1pn
8HLjXK6aDaVkmR5wtl0hhpBfTism5Pdjx+C7IG9afkY9sZ7G/uELj1xUIru6OsRO
dTVQ9Cu+0y7uvZS4ZFHLNdYisSpqVs6WHtJEghJI9ADqTbtsDsvXKs+/IbembgWD
P5WyorUTn6F99Uk86PkyhlmnY/T920rxVb6U4pwip4r7t1YbbwNdzsM5EiRaTunM
HDKIS12zKX6+/PDlzpnbYlTSDrmQz9Q8J0DOYFi30w3ewKCnZxaraBxqcaZ9hRu9
0BtH2cNoy7Ez4JSytWd8JKxPig2NpQvQVJhvNrGwqI3h+f7sT1NTw3y2kCQmEc3E
cV6oZwUNdzcmjp36BnIDfaf7dE63GbX9pUAjbCZfrH4MGQ6zgpAuTDaVi2ac2xZo
v/LNORHOkobDo9cXtIRpvDvRZ1bb4LqEoHoyazxjq7RvGuu7mBmy9xGQR9+/k+KJ
sXV7H8Aujaj84qrl8qGC46fxIKqGZfBKdJX+X4itIQ8yt3YYZB5YvsLhTpiYjCUh
EamFp3psvssWYj8kidKPMnPVHVST7hVp7p/decIAv4fHpbKupUGM1nH4Q+9hrc90
14d/znscdXbtul1rnmf0Gw8W9R+9+l6g7wrI/wIFGM8YPEjvH75vXoBHTjghOJjP
gFqWuv/o0nDHzHtMF5pm1JcyY/AZ7bpKaw8+TJyMG1oCoR2RQIUaX/zVPBvPn1P2
Q3vDJAhMSqqg4axRiozVn4hAHf5F37D4DiYe6jDhbYMafq6VOxRV2XsfR0gs86VM
8Ar2fe/SonwXWYG6HcBpxXqARpq1Aqc+aB59YdApNZUx9JVkH1LI/9A1C8iePozO
V0D/oCdUcwqdDHPevyoLFy7hk2mPq4WeoWSCeG/7TdKS+4svcSnzL+HTOL+S2VJJ
2FVhQe3EBUwu7VZ4Zo6gW1Wy6cy1PB94K3++u/Lsku4KgKv17Rc/52h3JIbUL69B
oO+RdEDtept7ttDWfCCprvZV2pU3v0BBGwwx+1cG59U3K4L8cCzmQP5bwgAS2fBv
7NCl1EPvRhRmst+nfl8JiQgILoXTCljD9DwYuOrydYF0u6v9PBkMghXFV3jBocge
qSC1Doc24tZn6ziDDJYE1UhuwryDGLEVsLwXlfFrR0s152saICL6qDNCGLa8Ga7P
aSrQApqZO6UlTsKc1Jdk1KRw7urXO7kjJus5608jBh3eA48P13wTsYnroX7q/Rjm
dShqaTwUG5q+E6DcmSozaKTwGzA4UN/CYjGm7PPj6SQbZ5K2Q6d229lVro2Wnnu3
SWT9DS24UJBPn4fbVmcYEuwDxYHGUj4uDgiMrU/aXBfCO6x007m7NCsxBRAwy1eI
/sSNiD7Ob31zrMu40giQJPDC0B0ArACr3Sn8GPncjdz+MFv9Q/GLpbCtiiSVyZJD
R+x23NQcal45F05wUHDVHGiv6X59R65hAUlwkjBxeN/+R2yY6Y8Q4CMRLbJlKr8v
IpNVNl+BAju5sJx39Pi+Bg0MnW1Jz4IcgaNm39t3whSsvHIzXLrPzV4VmMcCOFBY
RHHTNe62tLnYOKpCtxYYGj8h8xntFMeXrIRvE6/EJEoymlgM7qoVz9N8N3K3EmGO
Rz/OQV0P70jx6UAZWswzuWbiDpxbMXExlODxAVZMALSX7iGyuRfEiRNDmVx5JqsL
YQQ+pB/he99PMHGfD09c2UErJgmZaOKBqHiQnqCAE4Lc6r14Kc42vln7vE8GDDni
EKa/yd3/DunrfO8rsavzlifwTFpODiwJS8gogSOAqTtebKufPDu0advgmXVuyvne
Xl60fOu8KoZfSHcc+Dg/MPQ64F2VwSvmChfFIt9te+HAUVrCItwxuKDUatNg/V+F
ZmfiiFxOHEIrtTQpic0aK4+1MsW8hngkxNqixhRhT4okFChMt6hczbmbXliFQwiI
CzK0f1O2253sG3mpmPQPr9ihcyx2BqNr2s5LoGfAxRVXfr4bkxZYl0RpkBs/qkEP
IeQvyC6BOoHQU1h9HKOUITaXqzoGj6Tqewy6dt3ce//moi9r7Eidwo9GWDLoGych
8gqWpEnYCQ4+1DIZ4OS5x+WTaelI2Y6ONwUxgmjGSK/zXtZYe2froQOTupJje9oo
vJBXckDZkLVQw2zmQFJQk/LbCOP3GJti/iHQs+nmr0Kp+lfS9uynKSV3c1cF21kJ
lG0moEShnmlNF/4RqIYTg0oDSVUO9Ehd5OKT2cUJWN0UQCHt/EieU6jVFFAKD45/
AzarqDsg8+nL6PSp3UG7xWeG4zO7CW2bvIFf55Uidq3he7fKx9OSyr0YCX60hHo2
jTEkW47EXKMY45oGRD3QuCl06kBAgSleiU30CrfAwwrxmG1HtbHtyQBxEz6D1vRt
HJP4ULrxub7SSZV/daAbNWp6fABsI9QMb8K3QFpXL2j2npIIyQGxVBK0MsIXDfEE
IglnSoYSLhSS1VxUzltGtSgPLhJLbB8DeskOs8TBS9hWPBdKdI4oZUTAWOZxVvfd
gEy2Am3kiiVqUouT0TcTcDIdbQLC+Ofa/21grwz7sQPN+sQ68Aq5O7u3VGKvXnPS
9kFNqOkR1PEjVnutSF/KZS2O9nD8NIZ1E7w0ipd55X6wVffL8bjbNxNrk11nEf1C
sPkgMlAuWhSUtM8PuJ9Y5SsfW1xmKQBaHOBVxh5cZ1/joDEsz0S+1cbxhIcHHgWz
GFTW02yIUr0GbT/x7G4FxgzaPUSa1j1/ccYYOnzxIvt0M18Hru2Aut+ar4pjLa8d
SVcZiVN0uh5G1pif0F4yOxgkSP89i66AjgeBTu+KUHpoJtwwbqVw3QhvC696fXlY
I7xq5xvbOx8rQ4vJ1UOPG7BczapVEJGfiDL7a42HfTfq04OQsvX8pIrOIPGQG3fu
c/CGw1WZREGAuGBe0sX5IRrNlYht9bcahomIPogxXLZrfzO2xSGC+SpKYWXjo1mO
H09OBtOjfhmbrVxufTZ2sMqMHT8KTh4I7XNQoHh4FWw7rM9dqTgxwbeP5fFrC4Lc
ArLYAyih24XcL6ohqecbEY0QFcsxcDF4lSq/8BqkaimgPPBTSe4HgvZCE62CwkDT
Z/Uy+3KyR7MdHwRO35cwL6p84u/94Af05cUXeJc/OXaesf90qBsOa5cvz0zfOjkV
mqpKpsTKKbiWyyUvJSr0EN2JhllUAd+Bl57AH3dbXBf+cHPVPBiQh9tBfT+wA05O
jcJFaq519F7Ea26w09cf7eWDLdVQSbDYpPN9wvyAsHqUiyGsUUwYy5IBCONgSDmL
/BIdyCTlChXyKNGwf+SzhlgCF9Qxr+U3nj/E4l2DhwlH8AZ3pAN9PH5tJG7oQKna
E/gloX82Cz9A8YStnxhCxhOFXu2v9B0MDbBnky1qHufHLAkvSBtKzEInieCT04Vb
pRtM0cL/uo7H8jBtH/UrUL3JRO1ZHoWUHorn9bhGSDfvu9J3o/ZUncvZ1o5IsPfR
KpbEzc/jkVmi3drWbjmaj9ZEnawc7nKM0UyOjZ8Mz0Cm93u8MqOGC7aMBvHFl61l
OP1eKXouMDA0l+XLykCXrmXNaJ9+ZaJdM61qn2UnL6g6MsNxMAy3Tb/NGPTajO3/
ILg0aEUyh6GVm5Q9QPRJNRHnwlIx+wBKkPSQnBpVbJnEvuopQuo5l3e6qsxfUMrL
v8eoy36u4Uqh10HYdZJnpbq6OZSyX1jokTDT2WVt/RfXHukZNkkVxjr5zH9grSI6
pdwN71sWDaK7DmLBXTILmuLCLOFTJqWmRTXociX1KrJXLrWySIiiezOjoSW+mnTy
lXj4aN9b6Of9cv8Vn4x3cumgKrK3Qzt+AVEIW5w6R7N0JhBLprKLLGCTr+YnSugT
cMsPBY8zaUPmODt5bHTfHEwwF7TwdYlULnDani6sgflFtWXm9ZqBh4jjd6nJ8/Jc
+IR5EcfkLpZrprAEchdTr8OaCuea+VPPg1ayWhKRkUSTjn33CkRRwroHocYdtFuv
8LshPfs0heg11eost6IqOrd5vLtDi2lNXV21FZZmhWA3mV2Ie0/EA+s1LErv3sFQ
FMmDf1k+E/5xaPMOVj3ozQB9GWbR057j/D/XKiANkjtx3OTU5xw1T+2Ua9tlHst1
VHy4B9jO4tvsizXt37ghX7CZUVZKLtzxpk8xWp6C0ZA9ouiIZnNcufiQn5mY7UpH
Pb4Po+rclFX6ip7lp+IlUkjSw0TLybyXITRyG1+2Fom6c4KlxZvkU67ejG1hZq15
xZNCuuVt++ByC0P0XhJVNw79iE8lYdLpXqre0ELkY+49XH3uStKq8OVTX37jEoju
DzWvJ6tYOA4Jur4oFSm8fNH5JokrbDMhiayJQjt0HUxzRA46iLPdpIyKlCpWVFd/
Q6zUirplr2d49KvQANVbWTQTfD1JgQx1TwhLsnrWZu0YQ08HwylPMvrnD7k2PKhT
civIWOqezzG9WOXEDsf5WuKOLCwduUQdJQpc/cl9W7Lf5XbXstQjKB0cb+EQZ4V5
mQdzUke8GSnhXsnZ3N/lSLQVx5YMZ7Yphv4+hVMoGt0qXrEQ3G1UYy1BwPiqnvPv
QfXPp4PAwbkXXqOUaQs/MoQK/hgyefYPLm4aeeDU0Zpd+rUfkqccd+xu444NcXQp
aUP9lm6RLEK/F96+jV+js7iCLUI5jQl8oq+3INiIhsKxgqBfVjMm80IM/3htze4u
g+yzhPqDOueebaXnmx2KNPDBZQhW4QlOCuw9rXWx/sLLtIm/VL6a21LPfRM/qr9h
0jJyXRtyKSSbXtiWPeXR3zuPr5TEdkF/jHkXtvsyYehxPZgX/lGc4s7/dSbeZ7LJ
f34K6faBZcnUBobaTV6DgUfgtPpVzyMcokoQt31zwhzvV7mgrOzAfXhR16vBr5X/
1/hlavkOQ+uXxwudRqbEAoeIY2oM8wa5CQEuCbaKnEotlk16N2LaBvPiWANetBKY
nzWbiYIKB1X+61O2rYNNYJggVi/9VRTdQ+LVjMAXngf0a3qIdfyhyiWCk050uHPt
hWqXOuyBNzngH7u3Xa+gw99XJYxtvt+8hN7JmYjBeBs6SV0zt55yUenDDIcn2jIj
umjP7CkN/W/rHxumlNbpZHHsxNPE8n7AxaLJpafHcbQwPadoQ+62Jiqb95SvDQC4
DKUyVoyFj1ifj+GVyP7XzNuQ7OHKxho47vmsegpwbaJ4EWftyqJ0Q/FzaJrUh7+Z
ycXvjbj1kPjj4hmrq/ZCuIzBmNQdihB6J3FcWQOFnAXRsFGpqVa4MuI4N2x13wD1
thiOmbUh6QjZLzXtO1r8ubBKAZKboibSihQ3jwGtG3ZzpeUR4QETdHdQPt43Lzq1
kWNegdr1btPfMWn+6bD7ZUBxrK5aODhLLpiNB6mxrUMRh0wUu393cUUTNgyF1WJI
MOmQ7e06MUwyYXm9vnpe3Lu7CgOR2eJ72cDaHkUDe/l6fEC2cDpwHinoAb/tXfoE
FCIMpST/qW2GoY7NtErJg6tHrPYp+tIK2Ktcoh5/3Hz2ZlyEYbkKo+reCRDalPzT
LgmM8akCfdPNP10oagLN4AK5SaWrJxVyasSOVnIq1av+Ab/wJ4belHWVxY0DTg8f
G9dhek7Qjzfkpr+/6XjUP4/IRqblyMcwjH3/QGcGBNOyg+ZvtGTi2++FcSR7WULC
p6J5rhaAnn+nInm/g7+NcPfTj2uCqCT1M3AaOH6ziTZ4UcVXDQjsveAUB6RKy+7b
FwAxKavjaYUTyA3MuQewm+5D57OZCG3XFE+2jLXoQm91mEH3zfm09DEOVLLFMze+
ZKpDvPLIfRlWIkSg2dhwPEPhS/iVms8nEn496yPPNHlxsPzcshCE69Se88jrT3/K
7WhYcrPxJVUSfpEelel9Zzsp98tR4LYvAu9ea9gzY83xVowFRFdOeY4lnjiZMV14
bO+M27woG7FQ0KlyyXGITSMiGf04MApxRB53cE/dwQYgjZfXZ2HTp8ZTfeLPDp2s
UvtcnlPQhWemcVZHaJz2k7SFoEC6fWvuuoW+WWaLlYWuzm16OGz282jVl7jtLW/r
oGWZLjghd9MCu8QvQWkjJJOVs5u+HmP4wnXzgQhYICxGqmCGlTAyG0h8SvDH5qDw
M/CwMJ5k7gMW06DZT+jLi8qSSxHprk5d3z5E6IjP51o0JWxI8Np+8d9wziVsGLxR
rShSGBpr4jv2AdmpgEHZIf7eAzbmfUgVgF6aJZA5M+kMqOEGJWK1mUUAS5G7/c5y
9c0aUfINvHTmxy/XV+jNSb0jJRor/hj01GICP4we9bSOdyYdcLWt15gCqf80k2jz
qCK2G90OdT6vOoogEwOoQYSwmkLyhz6BvyYDTEvZGx1Ly9O7tSC480ZMe12dOEN9
t6dLrKFOR5lKK/V6SLDCn2tGio+tnwCl9+TwR2gwxmdpXWLxmO9eg4j8pgOZXdFZ
ZXG/FQSR4wyaGy5Uyv/n8c/Na+AGM88p/VqdlZbWVKpALMImgTBX9jv2UDqp/Czc
XS9Z7mmdPEjt9Iu15158uA9/KoY4Tg3jY4GSyoRmNfN2UEtNprwNAtPsZATEEwmG
yskvOrKtCXL5ngq5KOfRijM+WS58Do0tDHjflqfUWa6dJjCREEW+MdmdrQL+26OB
U4vyjpnuc1hpwzicvWvPbO6kHTnCWQ+8gJXDU+x7AiKwCZQd+so01dLIlP1ixsJv
O2A7iSY3d8qKIb5UdaYR7Yzosly5whH/B4XmjP4I5h6g1aT37Rs1P7LTOSd7Ggk8
lV1Mk5RYJKUU16HBSiFqp8ruoMbZ9axvh0o5sUbQ9kHuFD2cy0V14yb2EmCHLM+W
onkmTNPlCyP6s9n67FRYfO39s+UyQgBsHWm6OSOkTylZwHCu6817Vx9f637dFhZm
rTtsWpkN6ENNgKEGnzCVhFFPJ209nRXhOYM35wzCPOyD/6nBEc8posEXzx70xwZO
zOJT2RtTMqfkMij69T2TfNcMnN7w3+ZAqhEhObA/ymYMPg09uFIA9gIaJlcp5UjL
oqfIbN+gPYES7MbWuguUSgO+2XeWuMCNe2wSDJv+gBfhQYum1i7HHQBccT2uDKow
VP0V6gFrJQu0/Hvtj7yFbQCPM8gSmJaAJV1OFSgpuKto5a7KsCB+RkW9p8448U5+
4+MGWG8fTm0RYdD/a77wi3X4XPlDYIQEXWiMCAw3kVBAHcgVSwnHh5vyji8UcEVl
ZF7bheEYXvFUFwyp1SKd6GDPq5g4TX0IQx9V2tvZ1FFKNZ6bbyYxoXLVUZi2Jk3A
AMZdcSBLYvPM0jS6DQg4We8jCnVhBhIYuLyzZfcgsmtUf/NnJg4JZ295+KsaNA1/
UViZKi8X48p0QpJoawiYRBnDfdwCJ/0CjaYIixSqWcpRxV4fT4de6hoeqyNGImi0
c9aphq4JgOcJKFlXgz2iovegpWu5FX+mDloY7MnoCoz8KpIImfo11d9c49mtsbZN
CXNE9GsubjnTmiaGFplgGsaM17zNu3w8680n7Xwo7e8ne8A6AA1CuuIKKDb+icYx
Nz8hqAFOdvrbE2JITDGq0YlykQEP6lbtzFPhWmRU41D2GVUKL7rWXNV7uzXhXa4o
F3Zrf5d2x5VdfpN7Owf/8CxkFeFKURUJGW+YlbC7/14h69OfnfgBvk0IZ1sJLA7i
yyn0WD/S9IFUAVy3nRj9MPanJD6473lkaG+8kBewKIXf6wXogqON8QuQBOMKR3kp
iKZThWRaKc6LMPFMJZhrsc8wFCr2eE4xPqyh8nuRQcpkFW14WHIn3TDYYv9IFfRr
iWYvEDyqZSZF+iwH8jgkVTYata7ZTwCkkvQbdzTwAiZ0VP7WY0Z84/dvgUYls74c
5Ta3RiskICGVDs8FasYEN0HAiQFGXwd+Y7gPdvdcj9oUDuqXHG4vqZAzs53vLE8V
Xdxr8B9H/8r2Nl5Zl2OGMWXohv+9yZNTLZSz5jzzVw8HGxpdIyH5BocJfivUo9iL
4QtmTuohSB7gZMJ4Wf0VfpUrH6I90znzXZu4fs/7glt4QdbHG5kh5XuxXSg9Hc/B
/2tIJtZh9874hN5VJG32OMIBF+98J3yCXx7lxWV/BqHSW//KpQRNYIusPzXujdMU
aDhESaQZCAWFS2XzmgHoQ2Y9b0ZDNMmcZ5DmxcOTKTOuAYLNTvjq1+3vY0BH9AGW
vipHfWcX65eU/AquJgabg1wmSLShn4ivi/4+ft6dfjgC8LWo9UOPhqhw2h/2wnzv
JdHS1l3gFJhGIufc32rjb+hqQHkYLp4c52LSdwZS3WqaGRd52YABb1gEkDbHCeQL
E0mSG6MvF5Fk8Kxg54z/eNOeL0yd/sKVxK6WYovsDtSOo0hxinMtGacx0wWbWLS1
Afnr1dJoak6i1xpg90Rqv7r0txf4usM9RNDzU+GWx/ClswG0SMF+A5RLVachmK9q
EtL/wB5N16hMBX02ixcRFIwj+Yh5nE8gDq9Luqn+5GJ/IJSWRl1jbCqnef5tJiC7
vvr2B7LOTVK6v/SeytAFMgs+vt0RWhbcwgpmSFFGsJg5XCnZHfxYY1bInDtYaCRX
wHF8vqjXMt9I91Jbgz4eF4pYb+D5sTJLmhZBBWLV0ZlE+aIwGiGLx0M6J4joAQRQ
8ejGgVF0Zyk9HwVMZEolFFpwfAfie5xWFSAMKG8OigIwYdq5A6NyagG14/xu7rY6
fvjvPg9aYFqAtYz76gGydNqcDrD5CI4+f4taS+lUuhI1yMwsAwkAF1L/K3MYEIhn
+YP+vEL1Ws222tuyEEKEEpshOPcNXDyEPuuEbwDS1P5+HcuD24C2BDd0cQFudmOU
bogeo0EFMZxwgPxzY+hLcGazOfHPPxK30fgn82iaBAKzk1Mcm2mBt7Zun0+Z9Tt0
VJ6KoCHrD9oVUDVNoJ6dFFpIohrcryDh6Ad1lh15x15VOdAURh5t4xfezpPKY0g8
Pz/YZcnRhnDaMRnElLcUV0n7E2EZRcMLDJHJkYZP2kF/B7td/N7kWzREfE4L3sWq
phtMkroREtI0soCMykUERl8j1E+umFxHmUoRTYbuNsGOTiYrWMwlEZYpuhFCq2YP
FKv35GK87IJjIX/gC3V5v4S0UZ++Ax3tm5ovCL2gSTpX5M8H+6n0nqZ9xAEw1k7u
I0/bG3xNZMii0LeEQrlTIAN0fJdPp24cHpkkZIpqRHXdyRg8C6+qe6kiTrn27R/y
wkt6dkn17aMtHjMmVoU63tYNh0rN4zmkHUR/jyxtztDOSU8ZGGNadDJqh7HnsnR3
VIWq6k+umRFaonHcrBUWGYHchgc5T1Pi9kpk+xaWSK078QMoL0mHTPt07RrGLMn8
jXeXC+CppdOQSkIXXQloQ0xYNdwsLrnNSF7VVq9uNPH1WuakjHIpT1U+ux6yaIXR
yhCp1xDinZG3eIfG85JWENIeFoCDWY1ZwcukoCDpz0TdDg0mEBnvOmeQA8cCxYon
Ozk9JfFU9muzaq6cZcDpXji6eiXq697VmHm4USAhEJUWLTfO///pfW+HHf7fKA+e
jw3fYTHyXRVVf1sWSx/1vM0kWZzCi9DXWZyj1QHjqEzjEo0FuADRURFjAldy39oD
jrw5n9YKn4TMvCkIwH5aysT6Bj4aWYOQF/1I2BDY37qtPndcoEsMLwJYtFE41nAW
Et3XDFSKq8tCWO3LL51c3mbQYePw9By0LAKnJR8U2CUs2pDvmGvaDyiewzYvcizN
fIvp4nepqIFMquucjPN2Y7bgguiRbK/02HObf2cuDySjwfzVniJJIkB3XTv3gAtf
BDjIJo8mSLbl1HqpHeDTDlYCmHjbpQBG5x3oehJM5JXhMoMhZgtgaVQ2a1dIfq4T
RLRtv0TuNEqTaBJ/4EnPgHGWocoJWSHy6MDWaoBkLJpVt5qoT5s4sh5NuqhWG91C
2jo8W2qzpejwfI5iovw1WhKCfYWKMMxtehNf0S/vWNJxOudtlHOgDaEN50Zd96A9
uUsQOUZJZsvbxqhYW0TgJpVeQMBuo24JDOStZPKS5g4Egf5U1T5qFuRWMdQPYwFW
Qvaz37R1rM5AwR+iw02GAOH4jolwl+YzR2NcHzlys3gME59o9jrQzZucfUnJfi5a
9ncS3SouCnO23fIO4izHy5Z3gY7skPD9M2Fv0R0f4KM+E/VRGZg+LomtGC6EC3/c
Z8ViSG0itEKQoBhsJrfPglO2rkY4viiutNqCqDYVW3d6GfC2F1dCzwb8VYq/s5Pv
z3KGSX/FAsi2KZxPBqdghtrFIjbUItnMlNM8ZC8P4uao/GttmfXTaXXp0isWJrfL
ME35i4IwPp8qwmm9t/in+6n4hLa2b20jxyubMvWS4QjcHNU4jP/mwtWjOx9AbIxI
RKoAdH/FtwD1f4vu7g9bNeLiTnAf8H4mvIhD3cN/5kRaJ6u5CW+dd2DXtSuK8YL+
jq5HthTsb3fgoj2ztFxrvHbT1C7gfmH47PALlfIO/3YAEeFgxU4UXnHTB9/V83LA
sxHdU1qpcxi6ehaTDMSRwIlvYfTt0ajaVhj8XlWh4K4fHLDvsrs/c5Pq6gVFxwmO
n0oJBEi0RLi7GlASZF2k3FmNguD+mol2+4/atpwWXdlYgsKdNa7T59b57n8gzj07
7dkT77jsHapUJJ8r1SVsbtjRTY02hVM6IYvl7v12pjjbxE74MhzVINBvHKXHabzL
2/Rngkx7zhvPOjWK5IIWnl6lUxmKD8DGRdlMCDQN/bmAIngxkch0fi5+aBTItrwW
GbtR1c/o6eLoM0+zZLTt1XqnKTc2Hi35glzsXI0oZslG6o7aFjBN+b4yxnzey6GQ
1MBBGCaqzbH4CNGOMJhgPzU4uY/mq/eseUV2D4JOYl/2dzqO2mMwsYG6ioqLRMkE
igWtLJTzt2K+adMYl9t/dbzuW22PYWkhOYgqoFhVYhNzdWJArCBFDpg6usaYabW0
gwW3JdUe8XCXz0ysD+RlMRXF884Ex6eHhZK0HXNPZdX6f6PDvOG+ITwfHKarem6b
d3Ww5sZGajEODmfKqf75RS+vUsTzU5hl4TTtuE5hkv/99wBrUANvq9jHXheJpTdY
fUA8QIK/P7SlA10Sjo5qwIN05wqdIVibKzKG/xgtC0rnrGAw/Q0Ec2cDh6mMj7rC
msTjcqGw+iAgfObWn6AEQzJPRYICid/TgL1j/avdboX+pQSM1+odJy2plfQ33iKp
aUgYpCsXYZaCntVNOOUL2GYmPX4Hoz+Db+yd+UOwBLmo/vxeogKnlN0tK5h/WI9J
SK2kJ6r6fujdc0L9IWuCja6Bf9tUyF8dJWMLnZaUWhaDeyYU+djUawEiRp6v93aM
CdEr8zOM5TmDl1+VSJM2cGMmVEC0ldagadDjA6+EWTgWTdSM72UbikPYBjsQpjZQ
0YKKBFzn/3rs4+4oJyfhysNXOmflzDQiMF6L7QRWA8inNnpjt4yUF4Jqu9BmOJEe
ucshISbOzoW5/DCGycadqfTfhRrHSdNxGdRqJMyKFy8b9dJzlO4XAI78DQp9X0oY
k0LYrfMa8164fpkeUYjW2snO53/ot/RrVQpsslKWPEG6qQnSTUN1V8O06HKACrgE
aSlNVHpSiN6928NNsS04eLzzTZuytsY7vqTaux+XHor43a+EkvQZ9pUKmh5Dp9Zs
ltdKoT5/tdaN1ruXvK10TgburNCaRnYVyIB8j/xYvvj7e4VQ5LMbBGc1aURalPLM
uVdXiDLrYApnsDEdxB6oltTGr+8vbKrUb4aJNlyg44/UubZ/B0C9nnEy/QnNUmBU
Fo6iAaWLIA//wNezn86mpv2osb1VemaYRhSjwnZ9U5TK9SIg7SHAfL01wHF58MR5
rr0U0FaJ8tGTY4L3zVREsCVoJcj9n2I2HWxL5hf7gdhdt5UywuyurE1bGmom17ev
dFW87xjeQll7n8Ng4KtWGHjE5O37Q2yhQMwFusAC5/9Dot1FV2ytxklWdcIS/w+R
xR1Gfh8FnBTfJxHEHc2CIZCFehr6UnNrO3gNgh47g/V4Ahn5i4dReqmCi/RbY43K
SFfoSXbqJWSwLtDsFxrRXePPvCAImEG9pW2rnK11ACurl6QYsN9pt8YZP6MphTZU
QEzd5ZkVJR8mpVF51Ouak01fPy83naZYauDNLly6N6oS64ZoGy9DY411HgyuC6Cz
+JxiWyPRfnVEijQ2Z1/vmp8CmIuwX4yBBl2yTduaYrOFDXJ3ZnvJO5/2M87sQnEK
tAFpAXmcHlhvIYu35RlVNTWWyFguvAcwzJdy25GZK6bus2SjHjYK72Zcl5XkrT2e
UzBWCg4nKmiersocniYWED9dDKdOL29IsmQ7u/amAKma1TLJH+36plydttdcqb+U
aIPBZ5RQvtOpxtwKI1ZalNapUoxM/VOryyUhOMNf28pkBW+MaXItTc2B4g4N9qIL
WzaWmi78wPpeerMS5ALQjYIweqRtl88LLki0hGLgHTwXkTjC7N7nHtqsRBFq/tK7
HD673pythz9XU1rZZeUsmreoxVkybmflUVvhBOIc0FR5u3Rwx5Sxr+xoTEtEu851
U1l9U+v51t/i0Ct9RKMvnRNUuiMGijYQAinzsvgf1eVLAmDcn850O4X/KDjxfLIY
lMUZHA2uWe2AZLKcSkSxQ72N1oHNVKMumIAxu2Uedn4dHHOFKEOwJXHtdPjxVkbi
4Bh6GzNScGUsh7LNiBFfWMlsmK4dzh828UDAi0Vt94se5THV0WFOF9VT1K1HYU5U
HdafN1wzC2KuPaaTpReB5Ev2Wt2ttbZfFlxpeoJv9iNkC/zOuKbNrkBTF1hgQGcC
9UfNL3g9HHcPl6e7tPk4TQeZz3tWnesuyhUhpFMnljDhRyLQjM9b4zT9RwjyQ63s
1BTPFzIRhugGZbd3yFHuodq1uo7xOT68wP2s71POwsD2qa7RNhBYuvDfZxW7rGLu
m6YjC57hkQi7PWh1FDe05VTbTMfhBdYIem1bXwxiu7xOsHPnPDrq1LXDwRUvaFR3
96LUyk5MO8RNFBMyA8zxtAwH4Hxbcs+ErYPddxF45IHBgRvJUxeof4L/Tn/196+Z
C/5HS7zImgarBsLCMsCKI4cC9U1jrae651IN136Xa5z5jY+lEUI3SIvS+xbBR8oK
cor0UU1LLXJ/S9KPuhtJt3QGD59+VQzEbj143mIEYHkjFF4120P9qUBAl1OyHI6x
w5NwNrMPk1GDWRUDaPX7yIY8s/hGJO73ogprfWzQAeYwhjtYUmynVvqGVmKUyj3H
CMe6tMpjstsM7h45NuGpAiwrP5mkEPPegLQYeS+Cr/kjHtV+v3nA3DYmIdDEXIDQ
o3JFaVvyiYolpPciy49gyZfxv0UI4mx44LZTjUkVvJ833rSCvtmqavp3a5n7qF4j
4OxxphJtRsqBg+BkQC/U/1NnBChbUos8HRkLyyANDIIOZyjRd73xvCpgmsl/z97A
JCWKbVB4Th86W/hzMV4YXyOelYLI8bdSg+Pmwcr8AyPM6w1KyvUozdGm2AOebmRV
wIGQm++EO1ygNcLuUl0UlvkUWeL3UkWDvWc831UdQrt6hosiMJz5c6dIdiGc1YSp
B9APpv40sxf+/TwiSqvxFE8p4O9iER4NbP00NTX6vEfx0tq3mb6R5ulo5pRkFjty
Sx7FXzTCLg9z5+Svq/jsM1FzvYPZwzMgFwdKYrFNV8VMqlJEYRnWC3La1OTyXSlG
K7IhH+jAPGR2enB+7sRQE2dP7tGK19eyQb+p7GSdvOQECMXm5t/PM79RSKsRHEY9
W7uM0h42qoEzwZlC5sGBpQITqYp31U1dB3qwZwwFDgEihnwvsbCueJfAGJCsAKSh
VO17KxgoUZNVrrS9FAuyWYw4w1F7aCCkYFK3vVKhHbrRbRrH3bEIoPDV9OS5TsMx
1MJC/qZDRwPzunIoO/j+817PDYi+WpYvyrnVGqZO/Ltwlu+L4M8CrxayAtY03l43
VBxKnv3XbhI9pn7uA1f9uYAx1XlXSPXhJWyOAb499tGEGM+uokH4cFrnQ43b/NQ5
gSAAD2P/j3sBc22AllYmHi+MsfSzwrQQid1OJgP/hkL2BtYneteNOrbg11q7bR3B
p/niYWIKQ6SMc8FSec5thLXerdAg2CffEW0PvO4EC9DVItI77SmKAE40fsevn13Z
8QtKI3S00GJ+jDHCEVObbEiQ2WCrAFkC2mxJV4BihGTk9FJDdQN5uUjuQNH/nOXj
n0vlse4RodHhK+JJqxXJ5P8LOWQJC/GYgTfOz6tDXFhlwS9SqnqTog5HV4TDx441
2C3eS3QkyehC4mFVjTq5dCjmBVU2Ws2QIx9nUfQ4V+lEOsHn2ZJ8S80OjPPzDRNY
d1Vokkic5a4Bx0oFJP4SjhXUJQBrzpUf6ayrqCd2WNd36rhzzX3w8jinJBkcRZ0S
Xzs/AurqAdePQaYIQzqbhzTccKIniWiXabGchTtd1bFwsamJ47NguDC7jmkPYIG7
DpQ0B1maj3QLO+mOfZG+b5iXXNk4c9KqXfPYXVS3ZnpazobTXMJquenvu0/T2c7L
385VDhn0JNyIpy6ryzG0GvqYj16FGsEIL3b8eIySAvDZSu4SvCoUuN8OFCveeHIh
E4qCGgfCNkHnt7M0iEp5dD+bwW8BrCADnKGKKnoQI3goYJXhXGOXmj68oGdcL0n1
1ymSuhsfl5FSXffCxmXHaIrb5KpRQdnNXqWn41HpbPV6GAJNkqS+a3ERtp0rbPc+
CylfN1XpIayPEwFIv41XkKY5nXjB3SOk9z+Yr93krf4H7He+yc8aKRSooDpD94EL
sv/4EMKPFnMZMY+wnbbMMbgGBnkPJ+SVKo1mE94IZy4owc4CAznkoI2AbYvuXPzc
E8OvzzzFyD9z9cDRLkGpwNO/XKIFoqf2PCLc3T3vo8wJ2bD+VCglCeDGmQ2nDTb8
qkW02YQz6nFccirq3BH/Fi6+REZyjuUOJxex7JODqJRKohU/soK4i1+CJz42rioM
rzkHeTwSFCPiJJiFKXCZTqedlghbMVK1RRNgUIy821u+mo5/Uev02XWCAnkv813X
8zsc1isT5vV8RFR2wKM582XBdXbvaj7EuGfg9ZUy+dhGznxcgEyvgXZWp388tpa0
J5539P7KJ8GLeUwJuHevqMgmn9ni3tvNTegXNO8KMI23V8v835eoTMBDun8LMVuv
3gNpiyGAKt9c8QPYi/KYCgQy/7ZXIFhtl69iYf78KoFPxNYolHlVbTrtYyLGtHw1
9NDqB4/qn+EAnSJEwwE+2BwEymG93NOGQ34JR9bW4KKFwVLSUS25zMd20ArJ3qgL
9gb0KbhEdej9bmU4yTdO0pacg45xfN/Rc73fRIrnaEHIQFVnjToT3bAHI5EuN8A8
ARtpLn4Foarhk5PSGDk6bDMGb62+AhhKZONn6d9nj9kxWRU4aeXBwehPOsw+ouQY
SZ/+dd4KpMW25h+NQ5DgAW4WKIVdmhM7IpRs98Kee6bU+EnpC2iFGmnNU2NE6t9T
sThRIQ+qMrBPARYn8ojh8ZfKB9FrQWByjILiyKOYGhddd0V/ThHdQD9s5XQCW9Vu
wmY83FNk+NdQI3PwPCrw/uIaYh06oMHz5NrnwuvAQDMvAxZEdJn+W23IrIdSZfWO
9+dQZ2UTLeRD+DIqnMC8jdU1SBm4bMB2tmyolbxEP7m39GxjOLF6lux8Y7Ib6KeP
PX857mwZHPcKuKOCb/eC8K6sgR5MU3PGYldmd7GW4l1L0LDQZ4+6iMuXacbTqtfb
cqT7x61IRfjY4+H0LvrQiZQ/I6EjRiHtzsAJenLW8esHhkTg9qmxSZAFM3LkyJrR
pDUOcLGSmuF6VESAtrIyBR1vQZiAWPwbMannkOlFhMBhF5/1F+bUrrv/BBBM0ZQW
6bsQN0+TZtv9SCKnTXCD6hciMdJOzfSH4PP7VCEwE0CKqDYD5JQNbH+AWOJrfdgH
P8nWqZnaYr0cGq2oF7ZgCTTVmIxwSONpQxzpLuVAUKOrfFOrH/Y3o2jiE7JMRGiE
uSLsYhWk6MijoigbfkMQyivyJugOVUr38iey+Ag7lu4jKbT0SoeJpsAB6WaR4A8d
nEUIFc21tLAqeKQTqJtopMPOtgia5a2eHY7cgCF54w2Fwe/oHNg35sb50D3nVLML
OaEIRCkA6g97Q+Lt4DlG4NGifU9PVcaMsFNhRiqBOuc2FmFaZwvZ7glBWBqMO7iM
ElIMmDjcZGK0NPxhPzmPG1pqlgqO0Bkn98HUCHcVdgb+4gv43Z7fw1aMu+SelSiF
89h0LnH4BmnILFkEZ9mEjsTdI8vyZHxKKP48nKnIoyz6jbt1iOZnH0+Qcgq+j7mV
0JS+vPQ4mRtJYVc73UdY8G3TvM/0xApiD23VYQEwj/u4rEObDjQZ+aAPBDywvzw4
Y4Rtc76BNprGotkpLObs9FrlTnC5JMIH2l2M7ZDrONcbVzyNNRquIrhyi7BRhpry
pSbK5gEB9VBD6mDp/kmLunq9pq6+/ZnmpJG86Ahmp5HxAN0FOycoaDS6av1RdKgc
ofbLxhD/ngQmpTM6DIIvs6bzO+2iAZXrvdrnNSzm5mT29Iro+MG0iRaMf/9rCYHt
ihtxj76HhKrrH5OAqAuCDtVPXeo0tpeFTmwVWg/vJZPomv7G4PHTxA5I+xBmKkhm
gutVxGaJBMdF45M48z3xb1zwMp0t85eW3Ja2J5lq3lGtC0s8QEYwSb2vRJ2fBLpR
9cQ7jDD5ZBhxiTFJ2biIX66iLTTEskm9FV/RWwjhVNTerenRoSU81jrBqVrGij8m
1GEhOtSQ9DSTOuqYmcCTQbTghlctrv+oa3NMGGEAYXArjPPyepAI3cbE2JQ9QtR9
P693XUEAlBOkfzLf9V8UZ+VZNwei8cXayyfjCEoiaZAHg+R9uTCUebjp8STJtKjb
gmFWnMna4vSh8VU3/jZx4edHaZlSBeATdY9k6uvorlXe3esezgDSyrepo4Oqnre5
UZ+3W2y+kEEGirZTmT2CkjZnbqQncFgXIfM4AaSp4Uo6fa2mMwyA/kXeGm/tEQ1V
mbRumeNs3gHiH1bA+lGgTGa++xW+D0x9Oe5/8hZiVojS9W3qE0tIRnWK+my7lrJI
ZkgPOI7ANRJJ+ZveCFYQ3L4tmLwOGalgVIrOOQrxpoP5ww4iuJinir6Kji8scr7X
9iZlOg7wrsjR9dEsdrqJvTdnFMnoP7MyX84gBeOHREDfibRLtE5kX23oNtVo3HiT
xr7RU9DmaJq5dUVsivT1IJKkt+R6KitEg/xCj+ha8JqmSm5jqrpuquFWcvfRv6AR
7eizvcMgbBoZHcpagdze/3b/jmOcWhUJUJdVAI222RE2t8oGMgWqBJZ/qxJmm+9I
5WOrLEzm7MZh80PM6wrDCEcrKeMy++xyr4JAVbM2F5Ez1X23bzeVqn1rc/tBPlZQ
ogrwqnhX75O9/QbS2Pb57hqklKhqLaIOAHlOPqZZK1yMY5g7uIVRnQwYW9akZiu7
j/NMguzTmhyyJDcQaTygq1JRT9d9dv3JepjrRGi+zaJPsuKWp5U4PvGrAm5OZlOT
mtLIy0oLe7cn4z+yY8p2lXPpXvOfADxOjoB3SB6XjA9s0ZyDY5Vk17R+99j+RdtO
UgO+zoIAlyXN0Zo9/UrhOoWRffm8XncmFI8BACVGOZoZHQkFWLnv8I+G6Hk/HCAS
8OaR2bBR3lvSkym9gy2RJ6z+y9VtbJy8RLxDigUh9NkylKr/5PDJFyf1tzeF/c63
5hJ36pC2V3RJ/kyYRrUidw==
`pragma protect end_protected
