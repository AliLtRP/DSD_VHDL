// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:33:35 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
k/ZUX+d72FmNP7NURsN5aSXqjids5ZjLdiE8rXXjEEfOPpG/i4ojC3VLt4IHl6G+
bxzAZ0xfuoh5FoOjKRINc986MZyGaP3xrr/WZxre2/isGMGzARWR7/vTtypyc0fr
wNFG/KgArL7GsCvck7Cwvve6LKvxh/qBSRSMEAlU8Ec=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 22848)
duxna4L3JLrX3hZASEC59tWxlb2YlrsHq6SKOwQws4OkL6tGi3TQPjlUdw0ExdS1
vibBbaF6TTdTIxgRRTMO6KHR5HTZeG+nIJ8Gy1i3tCsMmHOgxjP3iDZ4BF5wtCyn
IAWAkqc08no2qzYf6/1MI4UkPtr3532EyY0UYovtlCw/+24O1viBP0AQ1T/49eiW
N9S9Z+Alr/IS0fbT49cMqyKvvm0Y7MJgdqU3RFyimCZfQk+gg24IBb/vrBo5bHdV
ovh1oCMRQlDiNHq6XqDvsfBd/0F6ri/raDzM/+cwaR0uV4cVtUJCZ+r6g7DdjofG
6CKMzpogZ2Gud82+bb9/zbKjqh2XdmTFwjhxoiA0U3JfD+G7YZsGrjaqWL6O/loj
iA61eRNx63KBrBs2Tnq61FWZqRdNXqmAhycO4wfMU02E5kNBe1HmdmLcyh8pCq/M
HvdHCEpx8SD+UAVOlqzZkt5MLxuCC4eceXYnQHlRJh8vFRy2hpzUC1oXhQZ3BKzy
HQRgmCUVhbZI9bXV6N7nyxBtEolhGshXtGzS6tHUx3qoiRT9SrQ1upVinRLQlopm
BCT4G23RJdDJ2gxpPFsuWzgiQPPeLIQfFELtyJ6iF52tPl9aKXoLe0thrh15WXv2
Si+QV6w/ZnHtdEMdBXKO8p+07yTDTYHLlFsUVxTvjSCdf1bkrvdNMlN8v2SfLT0X
rJZP2h1E3JB2kLUFDQ71pTzJtN+FSbSBlkXxD82lzLbGXaN/hBkzTkePfA0VphpQ
9rA4mvBdK3IjKhN9ylyS1AfywFvWKGaIZc+Uq51G8XApWa4rgkjZnBmrMw6Tdy37
sEPp1qxd65JHvlC/2BVYfoKYXusqktdBTYXSGBHm0YkK2WDrX6lRPsMmaky/eaU2
+aTAroQki2UQUWFCT3YRc45HmtzDTftDCnz4HNmzcAE7492ktuXthWAWjAuZd+m+
Qb/vKQeyF9MBOvdmcetnbNg2yRvOHiSDqWNhxPPvv7XfTHjyhJEYvNTd4+f+tsXV
skQvYOJlj+6alIynUipWU3TP8EZdXDMnUFbxufXz7VBts55gJ/Cy8VE06PvBmkI+
R8hwFFxGR2gztC6xefw92k8f6rzbg6E/pY/+hz/88OUbyv0kw5X8W3+UHzZXnmzs
x9TTfpzar+rM0V9z/GsjgzWlxrojemhNCiXGyukNYu94sZQo9X+IXy4ZnsAdX3sq
O3aSgFu1Qg5IkfJQ2BR85kEozPjZBQw+HU9sCRzIJsMP5EI0EuE2ajRcZ+211oON
fFSqf1FwdPNAzX8mprNgqoC/KRsQcF8r+HJY36CdtKfXsvg+bo2CZZ6HwJFUALLX
K9BDvDmTn4W9VRmNEGH60IVuyUO2ogRtYiQpRaEhy+mCDCmTFIv6kJImIINnR0AV
y9UW97GkZdbg3VMZIbKrUD7JFfAYjGXPf0QjsC1BGX/k2TiwYY+aGF8GjC4jyMQG
H7obtGNKMpPgvnkNLSgJ9in0pkt6ZI7sobJlit2xpbjRCaTS5JBNB1busj+xV6Ne
pwUjA6BOKlkAVTsTTJ3Rg2qBlaGnnCZGmx/4DWmk4GExKdaVL29NFzfVDXYxaU61
rMkh4r5yFmSU3rFmWDH7htLf5fu6NHMLqqXbwGzKEa6uBFV06Uqu2h0JfIdtnKdw
RvPjsj1CSnUTK428WYKT7wYLiBCkUDmzwhV71nwuuxGWCfKDtRhco8HyCFGk2Ujt
poGAII5qy8Ga4rxT22yO2lVvPfaOZp1OWbpWKXksetY54/s91kEnBnwTvrdZY6ok
I/JybBgDawPI60BsPe7Wa6wLOsLqL6BaDyytGVmX+cSigkCzLA/YPfmIIP1VmlMZ
GDcZBQngiR69Okp/mmSw9OxCkA5ygSWbCPUxN6Ol7+1dE5KjdgdzvG6aVPm5CAmP
Rpmz9tF/zhh0RzulV852N5iXN9rC+3AaycG93UMMc6fpbuyiubBVyzirRkohigAD
enQIxedAizrsrCYz1LL4gcuB/cOIenXCanqCX4vbG3DnQCmdVhSnGzMsHfpiO9M3
dVXO3BWwMj1b44ADcuke+Yb8D9hdFC7+rqlquBIpbm90EX2xuzzA8kDp6wjOfrJl
P7ZNBHk39sEATP4T5WzHK3gS4EmFR7IIkAcmQ+VqFsK0oVpSLHRoYM3l31mquFpW
QHvq51/PLmc/tMEGEry8q4RFK1b5jDthRj84ncgsfpggZ5KFqkxWVEeo7M8Q/A+l
CSmYvF4yF2S0dr93RMjv3RTCH8ZcVG2yfZraZkRFsPwVEyZRIkTsAD1ppI3V4QdR
998C4N6dBYqnZqowsqbZsfzFbtNzsi8ewBlm5mgYE1mg1WljThxLzx7cmLUSRNtV
o2I173zuHv1BzdAUDyoMObTPK7p0+ryQtBbkbucf5gaMmwJKpniP3N8X+GvKQSZa
OuYFApaA4+LH2+y9cZW+lmtv8CaaphwinobOINkhiJq4HnYkNmF41GF/MNNaRnbg
aYJ0YHu9u1YlCumhPDCEhQYnR4RkvE+Mxc+CedHk/1bZ6vPh3uPu5Y2wKL5zpE+S
p0o7ShSdw/Ybtlbp6huU9//39+B9LzTX9BPpZFDAGC9BbT+iEm0de0lwfJQVCM9H
fqYxcclzr+1ZR+wS0iBbRNjzwYNbeekdOKr9E5Gzel5OwCqBcAirgnRQ6NEGFzvU
VSpesn5BTXHojGtFbcy8EDqj0kQUs9kwYZvmC5IlexwLXUnNAWEN6LSkMuWdLJUN
W3CbzorlwEHCOjxWSqA4xenyKh6wHp+Rc7/DCKNJUmPgw8jgQFsOlePSUoqCDemZ
7Ct++haHs9CPzbxg46WT9xB9lQccsSYltufb0UF1GwuqqHY0EAlT2NJuQEZ2i6D8
kATgeiwZ/mZeLa4BSikrWDjm5JfYB6S7lPoA3sAbapCuswxuzccx5TeDLKIkdJfy
H+exux4TkQxZbL5kjglCh5YRehhuxtcTz5NHsP59XOUnMl/oLoSJdIb/FF5bcibk
5hNvq1Qy7keiir1I7E317I1yonE3UAt1MbLzsYOj2jiiKQm2E5uxopjfAGnkVFqi
Zj6v1M55H7ytqALVs1aWtPC6zcxaaeLO3kAl75kA/LZqOwy4fyUPwQum4yDc6cHI
MHdhS4lsdhABgkC0JdMFU8ziQoAOPdpiEZxBRmx/1KtpmdY4VhdBbMtmhy3u547S
OqahckeeiTSIoDFU6tev2nt3MIvLJXjR6oATI3Q09H7YdiGhPzwuC52nwFqOjX3O
XcBWDqwxaIKiQIUuB9hD8v3zVtPnkzFmyWZFAjVN3ra81tuEll2hgwXpLd12DQd0
iqxPY9uLzb8Eg/jxwktvrWOBs+ZSRcX708fVT5pVWZ9AbkhV5UkDio10n98pBYlr
Jq+Uj7Qcv+RbAkkXup24vX4Rp7HRdXCIZho5LxzDR1298ujnYncSnRt/VDoJ3x/Q
/8x/lGed365/59iDfuDUTBsoZCPTs886qEtCOS3Gapaht9WOATsj4K4/+vvbZE8L
EzZbW1lo/CJkDLQOejxPQVFU1xiwpSBwvvieEWE8HdXnJEr8QVoqYLwOzJsYkbZG
XEPJ1lzeevomGGY5y/aFjNAKjZNTw+3LiSQ62NZFPhBnxCaXqnhk1P3X2j65A2aW
GjtXvqjtYuDLypyRw6dkq6wqf9waIKMHz1QtcVrA8kcGHbXe/W1FeuD+DvVGeYOY
NBYsfkHy9fYqHuOORLtx2yvcRqKp8CFw3H6zNbM7cRG4DaQsJpJCDuh2RnMj3y8d
Lk/Ksyizw20Gy05PFOeWacMALKF2W6S3Sn52hXiEbZREFBhLKarv0iKkolGbgIL3
kGTde7GC5FlvrfIPtDHrKwCUh6IfR8fhzoJhsOrabx4yQnIows0tQyS5NySy+U9/
iJuSvbkiRW69Hn2FBEdy+y3q/pAXIf9JKrCSYiIgD8TzbuMTfnmvTrVan2+cOFJM
4d0P+OEHHxtzD+HlLVbhoQnSVMhgRaAgXjHmgsND5MyUs4GGZA0Cx8+yBsSHsAg4
BB1g3RNlZTcVWaInBJwkJMQwSkouvaDpi0ZBbup7DCypc2YFLqmpgbrHlvjrkF6O
0ZCh23hRNuqp55Vgl/nmqCskJhXtAIIUVMfe6J6klnJGrhYn15FWpojYp7aF6Kwd
G7oAQKJaYbWeHsgqGq5DgG61cHuAfybJ8p13+d7cXzdGwhixQ863Po/Q+p9yyu4+
1Hd+2DgREP+m9Znbxg/ESrYFU/JgOlHglZXqYWtO/G/mtd8HyWK1d91QnjLDI1Gh
kO9axa+28nhPNo2f2sYz4gmLpwV/WUCeELgbY+HQ5oARNArcimQIBrw93axyYSQL
HcMpfHRSKik9ESpVpicfs+s4Zx43FfRGg/MJ4Jfbe9GaUm3aKMJHwFNKTIgsBucw
3eVzJRNKat7mClrJn2HVBu39iWU3ARI6zvB2tSRFxqQJ6U6jZkS/1oZb9B4flYYg
5I4GhrfiHwHiGc9esCGNZ4jxiZMrxGb6VqV+0BCfldrIZNW4xYOj0w0tQQWcGs1W
b/WZtJ46QpTHv+xQc3gtSQKHJRhQxKEZsj0daMZAHeGri3xblHj3GuMV0myDaI1B
QVyPnc6BKHq/hxQTzNK8ujAbqIg3MCIgaajqaKVNfd6/bxOBvWTuI/iGYZefzvp9
Zt8hinxWB0lbJ6uBK+UosHONOSwWMaJRiZSuTBGYCV9x6bfNOYQ+68WpjZU2j7sG
lZuU9WMFFWwT7YwSl0TuQhC4+4tS4AiGoPYiQ3OPBIDjkxndv1DQMVUANn7YCmZf
Oe95eJUFXADca9EGMoqypv2uGyX4mCup2czGIRaawdA/s9XUhNeOrCxYEYArl/Pe
LfxJ9ABOuIqY40uez0VxUzS17FZ6SoEegbG8PJ2hGGhZCZsacqCZ/FzJpbVgxcbI
9gO7BIJv+Si91YkQvUyy8EkPBBOSKIFaLaByf/23aTZn35vNIVFausbf4wnFve4I
Slo/eOUZQFmb479ISiPocNURgcoXX0RIalblhM9YQRtWQrTLJhQNO9wMDlbGDmyg
6ODdKg9dGOYq2G9iAMIMqsno4jf24SHTpkW5MKFzlbj+UOiZZ/yJCzBTvHNRj2h7
pzeue4QdEIXud+rxE6CYROU7FSYRh/XdBLasMhcrImnS4JBi+74okK5T9ThZd/wh
tyuqXoRw18NkDAdEXHAR+4rmfN0G6sfbCnqLu8Ggw7WTLu//oHcKhf2kT8Wbl14J
9qFrTTCp7zG9wAyyQNsMzm/GLDocJhhumJMekNUfk+W9ZHtLiN1qNjAh9NRyfAU3
ySdjUINE8UoIFARid19lcWqX8PmvGRTCP2/2KeoDQ5zYu/riU9mYv2/DVDvsE1is
GYP9YPn6AE8WVkQrgaob+eTvEJOFTMGeD3v8fdAcTa6l/sSkFfd6GslLn7nmlPYk
E0jDR21HkPLLxNMmOiZLsyLAGmAVA9XPTQhsjTY82YjJatRz62KQoPbtsKQyAhq+
2SK3HjQSJscb6ZQ86P+61Vu8lA4bNogLM5zP9VQ5J7+UYtLS/QGvvTxS9TIefeel
PltRrMX4QmHIWpnHWJbCmJl0O6G1ZvyroMZxhxYa45pqxhKlclgWtiLoyWKCM0xz
Cn2f6+zY2puZPv/7ZHqbjq+O+kBqKho/yjH/7kPmUwpiX5De6nOciTx3FRi2XvSm
hHMEUHN/WZgRke1AC/xlhFy9rl9dQ6JFNJ4VABjYYj6QRhvq/57cf4qr7xrZtGHw
o/TYUdeIqxLvOKgf/xhXNxo7Qzzfk63lod+1EAVmvCEZNRse8G85NkqYp+IoA1+b
ztFzBJWVB3Q8RH4ngrlW//iOEpIrK/W6M6OxsGgP255kkfk9ML5838a4kpGTR96h
RqHJSSZZE8QhPaMB53A0SUb5mricH604I5jMZDpI3EefBdcU56az90tutrgSCDoK
bsHONir+N9mvQe8XPUei/Yu8BawZZQN4K8zww0ymGw8Rq2NXGW0KMT48kZWUbSVE
dJDDQbY0MsvDTXBoiyX9Fki3tzpOJoBwF9Lxgtt4H5ETSwvTwQ91VGleSXWcv3bF
Zc7ZYmMLy7x6EVTY4xYQMi9MjAzdpzYbc7bZouosfgsMl6g4w87OCJtWOsCEYSAR
D3Fw1Tf67TI1PrpZECWY+gnXb2EgeT76toZnVSI7gLGSOALDn9eU7quNJuyfKqGx
FsgDwvpaGRzstpyXGxTNT3YHEmY695GyHpZ2t/mV+iZJRkT22+WLxUkxfpdYfM+s
yFiV1Cfp13TbqdKRRJwzzMOGKAtHfVRLPg9SIRgaujMTOWaM6CeSp9m6R0MURuE1
rFLIgE8g8jQhgfS1zw8w+7VUDcex8RRMF3rEZUen0jGbNqtZfB8FEWkO4Cjt05kB
YFDB5uZucOZ9xFDG/Holyk4COuAUhuZMmqz3iUR/8hrQWvnIi36aJNwqRm6iYISz
Q0a2A3YJ3ghrsjL6bC52v6fh6hcV13YMKlb4JY7s7Wpfs7QBjE+VslbzdZblCqQM
sWo+JSQwG9hHvT7vXbL8ytBMxb9DCYENtYU6cSF8VUfwk3At0jxh6j2EzNel7rag
LuhKow0ooOo0qxsfQYNZ0lASr/+gjouxz7w6kmxtZVKrcpAd5eIAToM/4mD4F/dr
Vt87W7KKDk6prsFCpzU6MnICntD4Cp2QCDnFdwkIr2mm0UKbmYxSG4AW+2OyDXNJ
BdI1qhAW+pcthf2mwaMIjL0OQ6DiEBt506w7J/qylG6w7RAvjUSHu7Osdk2dB+pF
GFkCQGEbmK7P8efMEBfTPDS1MEcIaaaKtAygHSsHwI/EEHn/dnUwOObBNqwYZp5D
4YQVgqXNaZ+3QjAaDpErWHUY/NxpmiGAVPPd1SdMgq1e6L6cGip2lXjSfHKBmUWl
/YS7GZZQtkSfsT3glD7oAzQ2sTcPp8v8xDbd2tJ4HyU+YKjt7XcaRrnEuTpkpADM
9bmUtvnUMZsWwzg89cDzElEpMSOrR9EizlSbksd09R5WgLcc4uxgm35NFJ4W1Pc/
XabPie+u2AU6kI1UpK516b8M5vYlMJmiJENee+/bDsUcpaAZVcJdJrfTlmeb1eVi
AnQLwXfhqbQecz3w2FNdVOahXdq2gUWUgsH2OJFd2raVct2uz0r13usafl74SjQN
xjcGfRS+jN83W4tq6UPtkvykjd048XOBLeId1LqnSMohVZ1dA+KN5Jx7imJ+dtoO
FFhtyI3nE+QlhHqUFXUhkBrMT2on5tH+KE/+OFjymH8fMpth/+VI+mYfWkIoFtHn
t3tVoFMpspAo7PVFWYiulDKVUnFCVmcm4Olt9eTnIcw2je6PNOFKfRJRIJe3ob/V
M9VROMwgm2Ds6/ExFS0qrO+ENulzs/GlYR8x1erYUPiFZ5wEfsbouD9xMwZ1fCeh
/vhmpTbSvvn3Pd2Z45jWoE7ntMkC8XkQBgS6Vx0JhlOA0Yq98aQ17V2Ao8fS3zQ7
oq3ojSAXT0CvfVaao316iyvkOeRgDo06m1PQZPoonrA84NzQHjTx4JMok7ePb34h
vdF6NSllwPYlddDoJP6g0W7l42QLjhaXXV4s/BOnUVkyolxOd3ghWMsKiCR2W1KD
oUhS2VGjS5+FuqYNvg+zLu6PSi/Ep3mRoYEox/Azcp2YhsGUS2LfYZutfU8HrwKP
rKRV22smg7+00wIg+KTa6FWYnv+jewcuMxWpXoWOnUhG0COx404pxo80qSEFs0RM
NocJ3mVdVbl0kMLjsfaP3M+TOvGNsjJd4Ios4wIYWWMMQOUoTnxB8yvY6EuTKrP3
a/KMPmr3Qe1rcqxD3xs9/vIRumxMK5tOWm7jU15L4uwGj7/rD2Cex4ZjoOUEbh9m
RFxbhrkrf7I1U8wjb+SxTyBMnFK6EYWhBy+O6n9luG15YZOcaaUNXsVZv1OSRtAl
tJzZtvWspSm+AkMt8oZpE+mE8SoJqBFMaJcQN9Z+s3xM8TexnZFiLxJz2Q3pXy6T
33AL4HIPSt8MFegnv9SrFxzc9OOXQLKNcv5Prof48lo8lSZdJfdiOLwRtAIDGogt
dJ0BsKgCahVhvjbacB8bNO87pFbtZlx1DxQB3MplEfMJ/AtQdvGEjT6UVx3xYkhV
pkyfnh7l5gPkdRx7xpLB/nmYpmg/c8Rd54FLEurIExI5yAJeuTkYSzQkg6FC7ylk
reS7/KT/EMdlYKT9YBrKs9jyiwhG56QzBxA0V+VT5lrWYyCLmRpEk4A3mW7tnHtK
mseTiWz0xypZf+6Il7ErPhQeaf6tRFc+wI8ndnpI+phCHxjN/Kl7/2s0hT7j6ynm
9CknppGXX/eTOjM30AMZqHMaHezDzDhXqcxRi7bdRn6px2u6PJn/6CwSWvoKKfu5
uNtAgcxP7e9TXtmTk5SWldeqg+F9epS9sXBGDOI9MD8izhnmXcy+8m2yVUbfSjd7
AC1KghlyVwJxuN3lr7J3//rIYzAgtZ6s8oNFZbAIPQlrCESpHApB4cW9DUB13rwo
HtYe/u4zLQ2+k/ZoB9e4PRQFo3uAht1MSFJcmk6fbrlQiDZlCIfN7XrKo5d3Xh/H
REW8lf+vjbWTaOWReBWqI/47hKP2xNwdZ+OyQQa4aFvN5BwxeaSUasDJqr8sPIm5
wAuhupKj28kqb1LkNYkUYJWhqr0cHd13dBJvl0VHLLzNLqF7ugGH5469OAjl5Ixm
sWMqnC6BLdsHWtYDmf0l3lXvyx/dOw+O3v0ZSVJ22eWuQgi3WssHaNdTgI4Xwtfs
TmO22IWVNIXBxVqRcPbuRHHTvEAz4CEAFrZMgD9XXRSwm3Cr4AKE/c/SSIEiSp8t
1bTrlMg81cV6GvO5thFN4PtufE2Kpm+pV+z2YygmYIL35A/uXnUlDAmUN42b6I/Q
Co5gqra3Z6ZZhiyrFhjsIk0BJ8ov0/CRPN1hnrBsu5tlz4LKUFFRHzHdCJrPmBAk
tUK7t3CN51oeOzaQPzT2F3rHsJ0Dvoe7hFDiNy4TVfXbE1WzxECKBLPsBp0FAeKZ
xRLYM1ueIv3p67uIhoaPgPDU+VPR5Vgeb2EJL/bWpE0G1Yb6n1ZKlYeXzjKn+xeI
OmwDlhQWR2L02f4uEGD4Cq2c+HDwmujhICUIMV3doahm0uCVuX4OoPQ504QQ/DMT
93JBFVA3tdYtHyz4vIx5uedd1j77Q4xsffaXSEC6NzWj5I6SsZZ2x6MCc9io/l94
RlP/MEKgTjYqfpVMdkSYp5v+TfPTBXzJj8+F5JIO8J9QFTPS0kyaX5xsz3/zjYwo
nYUeb647mOPvUY2HLFqbZ1kr8ck+DNRJTXYPmpAUaVAvxbfLAb1Ab80ECoksFM7v
VSOFSVOrXorWK+X42BMEPRBjVJIJiUXo0bkqNE7bENDmDRXd6iplSY9MqKFnLKra
7OhJejVjeo/lgRsONiMwhUEKlW7qsT09u04MOyqmMItxkgVAmu60HwQsDIKrkJA2
4qdlZ24zbBOjp1An116hBaGCiHtWgMCzFafoCQqfoqC4RmWxvEcU10lED+k+6kDJ
BUz4H7+0RvpHecU83ggfOy57boJQUw/EcUaLVGDjOYoCUmUIvloPLwEBhDkQsTNy
Nr6rXVR28jpGqAefA6kNyJT+Tp9J54RWHQQqn95x25JQB8ThG+lyfFiKfRfXG6sX
Zl+A19cYiTwjzoav90G+qF1vJX2BPzyYJaKEuCQ58syNlkEQ/qltgNU5/iIPJiV5
EXQBzgt1sSzyvfZi9PyAz8w1C6lbkQdsTiANtGwT0l7IVlGRKYeNMSK+7eGyldZE
5NKOFDCw+xMbsJl/bhG1l90wsTGwASrXU8Xtslt3X8PCB5TP+mN5Nod3pmbnF0Y1
6eBzqjpo5/IXD1VAvHnlwUoazTFe3y4X9H+U5j6RS0enkazt0DWnei5dtkR86o3k
WrH8/LfMCZQqQymdGZBGg7QGfkDrvdO1T3tIRZMpCxJcacoJUuH+mdLaFOFHXo/g
KUpSo9MkoHq7PBBYhcb4nVtQqRgmXNOiMzBmQkl6UE9fW6OiNZEgdzUTcYVM2MVF
4edxf+ettgVTFeJEukZSASHEE4X/84sSd52ugU4bUdD+rq4BnFWSyxsBxHFcRObF
Zo3e3NLPfuh0wgXGxYyM17IpLNEtDkAPJncm7dIOjrRi5yyBRJFgDWWbdvvoRZYY
ih6dBuT8/xe5pj++UmmUO5iFD53eyNBn4oSHEBGWOkEBs5MaNUU1nL7Bd4ckIugk
jTNZwwtI7ixW7TbAfKDajI4tRzLNV5h03dBGjWmStqfS9vkBxFm739sZpn+3XBoV
oHriRMGsjQeQGW2g3Avhz+wKoxGoMOyGSZmYv9Dg/zb76bmxGRrVn44FSnIjKPrH
2b0Qs42IK+FX5qq2a5N4XY9Coa/Ts0qgMmmyewV6wvWs1HWlQDhekjq2rOC+TKKM
mJe2V9IPdylxDYerH56qoq7yJl/5H20WygQorUvkk9R7lXOGuYnrwr72xCFRIP3e
DzEk9iqW2aaKvTenX1/US8TYiyTAOcBhc0OApxf5mkbDZe6JANMIqU4EViTj+Tli
dx8w0lxmcip9m5Q1AghF8A5bFLOGCvX8j0aU8lUyBtD4Qupm1Ji60eSgbQECksFA
LZc+l5xuUf0vxjE13I5Ll5OLllMM6rNYOi090GF3Rzb3OApiyQEfogF46MmDmhKH
kDhBJPzEJyZwaqKPh3DVGfTD8D6Ney9LmTwbqivag4XwSSY+6BPG+NDM8c5aC4CJ
7P8n+2QVa4yGuMBROAhu210wVwfEl4PSwPBybA6Yr7LdL12wX7/ceNSJU5l0usC5
SvyhogIdcWgimcqQBnR39zr6TVIA7PzldJ+1MzZVKNyVAQ7VgGC1uFr17iYmt2qq
MiuKCycIU+cMiJPHkEt+cTvmstj2428omequO9rSQv156+SDLyBbZNJC3OJ36zS/
u5k5p09qODW3ijOCggz1SGvvh7DE2/nZU510QwgQEiRVdo0t9416RVCNS4AXEAvo
HMMedr3LqwPNb2E1h1npRyLQldeoTquROYNxAi7uPoYcj6KKYrTtfuazzBINYRtg
gikybRklfLrCpX4mxAFdD4RF1NYLLD5nrPs7wXkdX1Loz0G7CH1nRQan5S8XznLy
UY2Ij+jzOoJmkKJp5V4B/nXqAnKAPJdDCsTAqkvF1lpDtnGWdo+B1/E2J4iwz2g0
VPniwp8KjEWl31OZhidF3CLC0oBv0HTOi/yCnn+vOUGClu9z1DTK05U2Y8T+8lxJ
1adlR5oogh+5tTLjQBOQRhbAUoB0iHN6tQPeuVUeAqXzT8xYhm9IucmUazprI2LH
i11cvgwMzXWtZCXkMILdBgothRuZ37qjY9hnEgeXb1gSHPH2Dp0cTBxWtZDKXdP2
d+OgK0uU/+/AX0I1hubdJVy5+Wox3c+XalWsvdQT9JIyc4YmSeCI5zO+rTtRScRT
mZjBnf/O8msxM1J4byHahGpHj5fnadLkFm5W4fjBqd28KwN3U/Qw6w6aWgMmAvkS
lTldZtJAMOYfYwHOpVj3izzFel+2BAoJcM4IyyuMjOv/Jxfog411Lx11gSLbfRFR
Mx9p/IFXfKwXBfbvZFCjv1vGLNmZw3SQu7PP4838cSbE/4c87Q7DnR/inV4SDL9A
lwsJaDKbYqg6j703rOfFeHo5hVjB3hqCx4vNtoN/tlq6+reQrIb+UMpnhsWM1awP
gy3awgSxd2afknoZ5MojA9kyrefAG2VBmTonR/rmJbZUHyODcDtgye5Tq4833r8E
l+jhdU3FUMorXLz7FeXog1zAvi11D7yQ/oDNufxhWQqqwUEi+o6dK8/gPH3Kfqmr
MVoAkUF7qyn6wBRcjrcJ+CBzlvGRphaOvec05TV8VPt8vr0T2IF/25JOnuv4Q2Rs
JJUDMP4KfOdIsJiB2absBO95p39YB6iv19JQdx0++CcYcAPYg/luRbqPXk58i+6w
1GjAd9UHdXq7qlVNJJegaUIcyPYY2VgHwuY0FLY4PlvM4UXF4Hrl1cvTZhWoNVR1
XSDXLepo46CaE1552X7pLpiPcqOe86EIXD4/XMG6K8kcgIeR1fjo1qCOelS+g7wN
MlaGfM+Z4phHI6ZE9b6XNEcXEo3zISZihmxApT/M6RRfQA4mZ1moMVKdXA+evp9a
vv0rEhdMHAL5igNEr9dEd7+hT7n0OGpAK4E3e8qlzmhMNGx9HXMKUDkQveve6Doc
eKae1rXbWERQVn5ANca/YYHwTcdGVmr1G3aobyqqFXvgUsCgEHLtLv4P+HW6KQx0
yfv0DeXFnrrcHIpSEc2iBVSMWFazCbgBdorFqfmRNu5j3yOFh9nnlc4N8Hzuf673
nPN+BIqQUYmCdA3faLY5MV5pePbBm9CzIUbGElKvf/1Xa3k8UnSGKbICgMJrRP/n
i+1SZhv8eov27iRgDFdxE+r+Uz04oUWLrnQdlgzhsKv03zO13zBBa5zo7RPlOOKX
793khsSmCBUpXcYWHCTIvfUNwZUaFSj9tFLooTMy6y3uauSb3ihLcz45o2CC2htD
GDcv026t4eq26jHkQGdFychPuOlMEVoxwT6+2vkgp4ErWgHxa5XikY+qJVj4JjQS
t5r2u5HLJlYnkKl469SS9Ce3V8WK8Ua09gxN4fPWl5OBDL/RFcYwhwWuv7whszwg
vWK5uVQLWFe0ziuRc4J9wF7Sz3N3sn8PCuXCF2S+36YfmP1V+yLLUKidWuu8a558
R/pQHuFqT7jtUMBfKQeP8DjtpYMJ1Dfd0ue60LHrbkCWWikpoW/kt8UTsR317ZpR
lfTswvzeUxuvhVeKVnt5dfohHqyTzOuDYFOiQppgwvxTTNI35arKh+x0AqLMRxpW
Gc51Min+WgTsMrzKbH8Wpyr34pmhGtvojRrHaeQbZnyjHOQLDgDpPYv6X1sOldLS
y3SUE9jVTkjQgRRDFNNKdI4NwbBqp26GsZV8+Ik+ezIWB1j0V8iEDR95zQo5kF6z
mOPPxmWsz1U5BBNHG0uHTt330TbeG0Va8D+Lf1MhaM8l/gpZ7ORccivgSJvybwNs
/atAVYejS9MV0IarobCYK0Ts2XSES/BUIKtJxVV8qJUtqBZj6IF1NXPW9xa/1KdY
Ys+xpr06wzoJtd+KZMgYcw8lg5SvHfNXIRDh2Djl7imuV7i7CHrCEGtmSvMgq33r
DLNy4Qr+XYJai9kq6g42VhmAq5/QO6FUDicM0dgBiVZptOBL2GOPUUoknIO2c8sp
WKDPxfX23ToSJW69akCwWrR3T2MI+8vZEJKQwYEwcIQMZzvzN3EUz6CEtXPW56b3
+zn0tRWyDepEAQQC+6HLHZWpGwagmkp8axwMCZjH/S+JfsY6WlxyM4a5mStUPyr8
fQVKSVn/bD3faUw8SbbEAUXlDH1NDPrXQlIfPPFyE3wdOn0wRI7iuSRrGjYF81mI
lCd3jnUwmcTpyMmvFy2c7gP4/vB7GypD3jCfxrYkVzSR+TgUQMgJR56kIYMV6F5m
WBmtdQM+BsEhckvdwz5dGBhCWd2K2UZg/7VKS9z38jz69oRi/0dPOMkPJ0Y1baVB
QZc8RPOqk8aT6SpQA9bZj4i18up0O6JurI9YHbIbWKN5ns7+AKsFJXyJyaxrfySk
5dN56ZjH8fdWs0Don6lk7Sk28bvcfLMrxKSNVJXtandtLh8sNBLmGDE4VA45SQM7
rZXaryw2BX0rpat3TftXlztXJEiqYCzvIsvsJzkkF3Xb1mqpOaDkz7CZTmZIJyNm
+9+yvNB3RbDKOrAvAnK0KaXx30SX6LfAlLYTHqIvY4ew4sOgyyBpq/prwBsf64YV
6MpsVUoZ/DJ6JIy3pea/rqfgLpQpkFf8AYRXDuAnqEY6ZNVxW4c7XMmS9fOUvKOc
RpcZYp77mHGgERXN5ZbPBxYITkyYGnB4y1JGaNGKlZHpKpEypYHuiLjFi+PurgL2
WAGlKTy0rATCOolpBEkiGEdN/LlNa8hczmJwOmIuFxGIDwcMi8hEc13H/4FtOL1M
etVEa5B8r4f5F4zclxuuSXT622X8neUMqNHm3g3omFdiSZu+NYUYBaDZ8bZX84XB
tRuGb4MndxfxDULCRH06+ZwR+CiEZIV4p58I0CrWkMobA9HgTi9ScqceidqM7Ggs
g6OMEsuG96BLWRSoswgLg1csUSprDUvePj4Zsmj73xWa4JCdhj1o16yI2uVs7Kns
Aczqo8RvPU0g6Jbz+6hKTdpnS/B6sOgBeYFnM2tFYMCPdUAoSVXfick6ACTREVIA
rq5O54HJ/ZX6oBJblV+a6UNqSa5F2YGZVojoV8XMgcFXdFrxd3ph1szPMTGP2CyE
rwno0XXH98z+RWvXZpslLooZm5jtbEK+MFr7s1j3xB5oXuRmXumSK5e3Wkcn25Eo
MEttLi9NVSXUj3MNN34Tk/f+962aSIvoHsIwqje+RR40A4x40cQrbLdmliSgnrik
ebxSxxbsGWR6lstfGW9qbzJCXHR6mOakil1dTCfAFSNZxYHIwFy11X5loCPaKUka
PH8jfwqKdj/MUJiWQF0e5YlyC5EqNDoeqEk11F//XLj1hLHL7kCXScBcaaPFruUs
03cqvAupdv4KufdwQiqdgGiaGEPOVcgRJ9Yl5PTarY4OgFWN5nYuJztNwswZhpPg
WSZqfCvaMiaV0oYTnra+eSnk6F4H8p1yVz6ZGWt52juJTgCLQBXD2wVKS4esOLWb
HSkok2uvFVQXhrEM+KCTB3Kr5Y8YkZ/3Ru4smL175zrf4mjIkJh0LVNBYAjBhQHJ
MOAyKdzznSyW7alOjmIFFoB11saqJgcCOSnthh+EAdCPBjHAS7/8YbKaSMQNd35W
36pKIoobZAr5HDXihmSlzcpBFDSxj83Ej1pktUDgGSPQEO/kjGtKnezrQD44KlGU
/50URidq/SDodsdwGVUB+oGtrM3Om+PMe5/WwiAjFdoA4ZbdwTYSf46bNEJ1UMow
Kyr2RwNYG1fnpsrMMLnQ6nqvHsrijPbSzBkxOdBmQicEKu/3MtDOJ6VgaIRJy81M
ddxBas7oshRLtj9C6oSGTTPhIMGjZp/QAYHfmVfSCo6AQceTu+W1ZQaLpnavUF5j
q21gliSsWrgiKjxW7tOrMXNkqR7ZxD1WWkzTZVR9WEghnTPq9qm5kn1yych8Q1VM
Zq38ZJInxuJBPYLa6k0rI3mgOyAxlSVOeXfaL3Rj0GgrHEXg8DbOdBXFFzzyVx+G
/uNSoThuXfW6I4KK4FdhzDx3II2OsCjcu7YCLyufSXQvpbGt3Ze3XJ+Jn8oAOqtH
9titjWxNLNNFMtWijhEHD84lZ86qC0G9/prDgMAJQ++dodhRgIHzbKGM+Z7/N+l7
cfamX11/2NK4cdNpoq03G3AxdiScnDUR/Ap8qf2lO54vMw2q39YuCvbUBLf698wj
PeZODFzWuWwt3i07skJReK+W0a8iAuW2wiRgrT306co9yLLmYojxzaY5vRA4tpVv
HIEoM4YIN90lDFKqTJ2oFts0McE6GA1cWbnpfdm1J8Q+CiGnHNPFHXAjED4ASGGM
1fDtjulSPsv6iDVO9hEq3r1XRwQFphY/MBE3Qut2OCxFUq2xFrtzObUN6u3qA3yk
P8wiHyCvFdkDjP6jgGhDiz3xNP4QBNuFVwMbgo1qQiktpwQ2LAYmh5HvNVHNIPKK
x/FkLSEXaW0gwUNY06oepSMjeuzl6sxAiYiK3MK8plOUh0INixYZUyXXsoAmy8T4
g6Qu84SQEImr42faMZsUMuq5vz/kIcO2fjvkPeuADOV+A1rfFptFEUDjq8IQFkDU
5q78gB2dcV9gFyUXtSMO8htrtpWd3vfeAhl4jKPeccv6fYfzVTJYjscgnkzgulCm
RglwxLeg27nJaEZ67RFOkpfzfwP65sndwxZxbJ7oj7QVGF21oXyTzl8VXLgG7hCw
7fqSYN/STgkXIkx1BULNGRmZBD2p0sXHneNsarAT2fsU1J2bvMEVF+NZcWsBRY9e
8Hc93DsBb2lYWahX4+z60Cm+85+sKrZf4CMafqNa/nh+cz/HAkajtxcuq1C2irVj
AGQyP83JtfhfoI6FQ1gRStHZAUSiLO97abW14u65cbciX1oGkz1tKv+Vu6zMY+EP
Oj2mE7ocV8dNFvp2pc2KLmEGM+cpsx1/56X4/E+iYulG4FKypzg7aTYHJa9hfe5J
PwqS8sOpw93r/d6iyjQ9rxyj5ihgps9iSoFwaliGy1t9UkGzTufTBMZDtHRcsJfD
evDHSCZ2uMZVp4GPdhj152EuAg1A+LagnhtFb0oXIpw1Z3E15lpD1ixfmvGy2nGk
KRAuKA7JD4a7e6IaEvkfjL2JIymWLSDWl8Dw+MIoQnUXykX3asU+FXGiN8MFilA2
Nz8R2eceZI7p0iEjIl3d0KwNLrtc3380HoP93dLU04NyEHj2/p66+U2RGs41v9Sy
eERz+JKFLF/TpkQmvvzsMOfDQGWTb4wyAOqPO688+ESgODIfToSbLv4Gs/zlaku0
Of6OqMSPpotwjnpKyrcHEOSQZajPMDg4grqMduGaTlw14gQ1OtQ/dzj5MNZXnFDc
TZmExDKtBBQkCrJ9pE4v0uBYzLqWhp8ego0vAsSkiS41jk6ln/9QxULyaJIpyITv
BCpEjs2TjDrlVDsNxa3nwceumdP7YaJa00WYoagFywdUgf6q5e/Q6p0NZpqhqbhh
xP/Zw5WE3aFIorQhborPy8r7wg4c1/jBrpIjvVWL7ztIHvx8OB63pFFg6IgBFIXg
NlZUmAo/30JLPOyPWPMkHnorELUpPND7dV6Vsf4CipLwq+z52Mugl/1vR2MwA2Xn
/7hsEdGl1cf1tLQxgjydekKAr9sUGjB6xbs333zAv0t/gsZbjbKyfsYcVJ5JjV3l
WrDFcDqGDXXR1aU70JIakrDXiUZlUKHKqqHE2E8fXgUDOfYTlWNjq9O5LQofm4ye
wHAf3DFxAFqma/57Vf11+AkKFqqmflM6gKo6L6WN7iV5KlJjTgaC1zSv4qzDPbPD
2wTXdWrQfyt/kXlH7yXDzqaC9Tw5cNitW4Cy89EoNh+IX41Fev609aJrpTZ11A+l
wiNGdmkH5K4P4bxT8uI1rOG6EWqLRL+FyfxnVP914Fdkdkz6i2P+iLnkURSmz3lU
3X49ShPV0LhqhxkqIjxeSDnGqGW4HzINBfClK6WRMuZtncJlgQCCHFTPPHMlvinq
oS/bULsXa8JRsibXElGjsPU5OKhHiKBNBJ/EObAb2iYGaI14Tyy4E2mP3KncVGR5
RECP/3caienhcaeoSyvjOwgSUsHwjNfQdmPwizv49wweqpYYiT6YhVUJ44okdchf
D2ZsNasPxbbIiuBhhG/vzC9WgZ98opmppIafE7Phg0rQo7swKmsjxrg/MKKfvrmH
H1vA9GRVZ+qlZehJuaNvYR6GpFvOjYSQTRg9Mp2iRKqxkvJYZ6ldOWvnQ7Lx+EVk
WSz5vhlNgiFXGDPXPy5B6lUFXNtvPTC6gScIblTL5uMzcTWPyOKU5EyVobpUku1I
CMaz2m2kiBQsTVgvU2x8HjIwhmrZe3hTvXYAkspM3iysiP6q0arn9ocUZoomHmtA
S5BkK+yu7tP8d2D8NUZM5qbn1GnnUSEujXrOE/9o5PFMu7C33L7gER2cqe5Kgimv
vv2jgVwI8vmOeIR2e/lrXd+ge2T5+fQTXivV5UoOGOqwDuzi8ftnFl+qjyjTR2Vb
C6LbXZ1ycqT+47suToIwj34xJPRx7KyG413+zMrQbrQIZ5o5VEI422MLz369b4xt
oM5wwdYwAuVf2vN79zQZMLDDg6kLvUpVZDtSry5iCsLIopNlASjxZHKGCjkd8FkX
ysqpTioOHItjmJGMh3oUaSbB9RvDwRA91ToaFRjsusgIx2l46XU0+8i+R6Iu7WCh
Lqkd+BV9mT4jm7WuDVaUwAKrHjGyamOu2pjObK0IdDNI/wNisfu5y45cXo7lLY7Q
rnPbgSRdl5Nx9T9mrUPv57IHK9dNpq+E7Se4o3cg8ab8T10SH/PKqCoAdfLqyXBT
BCcsViRjqn1o4432QgjbhBP/iszayqomJ0LLJaktYcRARdGmYfEVyx2mOw9W1Uz+
0UntXuROuFgL0NNLRNNCSjXKb0Qy9NOyNCwR0Q7g0TeCUiBSmagZaA1p601OuhKu
v2jjOQn8I3fCJo2Dwp6BUGqqJMAuBiW7XJNGc33ebiYz/M9/lcu3IqOxi0I4eC1q
SsQHvSwHnh4KwXTcUrg+w8INIYI7Q60MWrIsoHSAJXZSqxOG+Nbti+kY/PXzT2R0
loTfdXZvqA29SqmVg22W5LpiBFBFJ1Q5oIZrF7YTkLfX4WNIqxS5xgrJDzO84gM9
XxjugUilPKH3n5aGD2uWmJ0IqxJnUI48320msWAg18y/U31vo5rLeftLxJZ9tUUy
WDN1K7r316QWhvRolRfmulBxMz1KqqKrJfMVVgn9IKZBgWqInR8HFp1oAYsWIGkv
wGueW7KN97TKX0IBT2dKR8kl3rQdDEZK7rBBpp37nSAMIU4qrzmnBkgZTc/fajMF
42MelzJiUpAyqgysUyWacuHpJEpyEH8EYQgT56ZPPKcq0TAnk4TnKqrikDbaO4eW
1TZXP/HSgNQ4kNCFBIJw36D114lVS/PdQh73df+UUEeh5F8qjEO4Bn7IpRJsthU4
PI1ixYSNbkiBF3Qws4+YZK7DMZv01w8lYek/qNMISCP79M96Adf6vgT9ykfPuiXY
eyDQkEmus6frR/UdhKFpir6gvZk0q35OJeR/FpJIaVd60JN8oXo3eSEGQXMylcSu
M88+N7AbsPRCdu1yr89P6/Oqiu0jqOOg5YGjt4Uxexdj0vgq3Y1kBlQCOIAbT/9S
EkRNyjDpUzKjyUjPIa9Zr3aERRq0u1SSXeujCmxmsirhWCMzxm2aTS9rVCPFeJ8j
2S54HDlj0hjWAPU102/yITKpDJblTnPYJmgYiKLSlHSmG6dia2pzmhtQQ/wJw23i
XtC7FN/D0kErt2MDzmKj32YVpa7aop7+rXEXJ+L/Yx84mZN9wMEgKuTUNjJPm4SH
I5VL5K0xzqDMOn7rY5Bfo8BuWAUDXw0cHHksg5QhKqiNLTMWEwOA3pHmb6meATZ3
wkz3Awy2klPEOMIiCqnhQBdwEPtFSTlTtUZPrle2I4bcSdg3Ew8jAYJASeYHvziw
u/23fzpXOY2718J81OJTvOc3rGXlavwaAla2daDz27w//vBzB85qwzFIeSa0yury
e2zhccL7Sns2KZ+BQ+e2GEIX6OHGzfN6Eu7xEOGdXp9CJNOz6mZ4t2pEoclTwOfY
vixhd8mTPIakZYwC8snGa1AHdRQJY9F/poj3wIvMcrXhwLuM1MDpc7qsheT7ikul
wIpWOGEI4w0boFtcbbS1YKJ3q6MNHbBommx/UtnlGMy/lE2bI04Ov3oT/j5KJ0XN
W11p45Vxkp/X45Smw50f6Vf2dTD8Pj13ZfHZnla4KF8HpqLNpwUDIyuezFPJhUN6
uuV/BymSBYtSCDtZrzvSihm5XyYXC5pALg0onvvmbGhjdESgHN5mfd8CAzQdzoKS
Dp6JWV66H+RSM594haRFn3cIeRPiir/Qmobu1tvauCOuYjNQXLrtICS6WMSy9m0V
Ce8H77AWh4ZmZtJ2JSRaOlkYgeV2fXOko2uFQBXYg6cstBYM8OQCZZ5PkS4SdAFu
NWL8e+OiljHGT2e7/wnFz8Pd7YwFqpoUSgAZz1JXfB6ZOdV7qgJCiYPe6mcImL19
TRdIxWjYv8bCRZWShiTR2NnGQHafpW01R92rgtjUEHj9bMZ/8hQPB4gG6N9v/XjI
wqW5GWvY4kZ3eJLp3jV5Ufr9DwaHTDcGQHls2DvDyZkRMhJdCzP3e5fJsMqb+/HV
Qiq22hEOy1SYZs4S7JwG5+WslHWTmawcPjwWpLQLH5YFrUbpYmqOfAy6rfHUKAzx
X9/lPf79x0HX4sucCT9skG+ZXm/rkB/JS3WU3ga0yFkh31mmP2wYIdHW/GNif/Up
GesMLNxCjzkqiQ13Vg1wbXjMNYd4g4KU5ngG3FEhwO9Iod1ApYFPC8C5ImPuH+Bp
Inl1tr4gc+xtgBFI1mBjWWGUGqmYXgu3KRY04cfdFDpWfSTFSeZrCMdN+ySRshkk
a/gzlc8lXkrk/7FhYbhS+Lkc8TMLP1ECHAJg2YZhtklzTGVFRnfH9kCIBnaCQ8zg
+QPSWoipG6tmjlv6K4melsamSahqirRHEAxI1sSWHk1MJTeST+UK8wEMb4dP+V/2
BBd2CFisGcq185Zo0RN7xton5K1aHYvm1dw/RaatNLr25IVol+3FzBSRFUNuJCm4
p14z+B7rWUnLD+zMroTZ3Y7TeJ6HIEkIPH7qTBmdNqve1yoZVhH9fM+vFGemk274
Bvc2t5ouxT/fKzWAwVC10K++yvr+4W79PkXrkgJEJiEw4Yc++/2nTw57lzYF6A3k
MdmP+GD6PvnO35NNGYIX3bBZ1oDiOQKcM7bF8f2QxSTa7IQorIT2IlKuguHmDBy6
jnevXDWBjMpolEcQowRIyxi3tnESLQZKj1QBPeqRHA755NKd9MGV+gDCU1Zj3wyT
y2HrUDzJxkXn3jN1gaq1hBq9MBMoYx2Y+7SICviUzS//nmDrxa8RyndpFJa3rh2m
He59vR171tTUfuQQZTgZPA7Y9qVIYnIUOCRzXsTQGOmk30muQ3B/iFDyfMVJraog
9XOu+nmxRyoCPrjS0NldnNsL3XpnILgoowBtfCHl0VVR0vO3vBHfdkUQYSJNCQ4t
8XrsNKDRv82Efk08NO8hEGbrYFCkzFTnlp+zsO2VZnh1Aee9w2DSLfhNiXcpZmlb
YGEqSoDNazoYWOU1u5OQSW5Prv3mWBLZYj/MAyqyjI/zaPN5t/9+x2GCBvGLzcRo
oiYWvMJRy0/NoVKQruP5pESbuC6QQx6aBxFQlFLwzqenkFKzro5f9zX0oBAiGk29
1qQU+2uokC1YlnQkRP/E1gUpewRjSEu2glMNJqbV6zN8fzNNoYDRGurcOT8vKuYG
uDdPFCOfGF23u0jaUFeWB7zcxBrlBnOGtNIlzHBTCeNKnpK6Ir8jvtexSBErUvxg
gjcsCnPRmuyXrZjIymLIMV3popQFRzV2kjEPZ7AoO1uG27fMaDg5pSHl38dOIxiZ
/A1aKXrd/5Eb4C5UxzXbqx7jYaeeFJi0seGrC5rTbj/5pwxcU6j8UQg6LNpnOJmO
ZzxsrRMklJGWcFf3cOEyiZLR25fmgx+uT7T65g6TP9HlrcltNvmwiJTJAMxaO9eL
mHd4zBFVDTqF4xtU5Oa6hwqGwwytFa0Te9SM2cF9/5zZg37CPbF8To08SSuNtu/Q
3mwlsi89sWku414Aa+gFk7ufJTAQR47JY/HRHPQkM2RdRKPBSivIqX3G1uJDTsws
GUoLWw/fT3nDV96352pX8Q2dYRuYS4i2eDycMitGeBqbUYq+kc8mN3O1Dv9OiwoZ
5S/hFwnLPD8+MpDXh5ekHmxTC4FOTPE5+dPRDyeYCyiolS63drWhB2I6MawRQCS1
8k+AJQlcmEuGgXX4mnQ0aSozvsSIt0R5ajcJco3n40BHZFF63rgshD0CQWiAsxqu
ym0zIj+LAUxdPrITUpqVl2lSsW5G3/rCZtXNm7pdo9t7WZL9oJYQJPC6OdJCU+qu
tVAk5Mklc6tWOXB0W8sAXNuQoQ5VPpnbEFPkpEgXwK/lRp2z3EKAieQpeDLLzFAc
5Bn/o1LxHFnYeflFzy/lvF4qfe5stMylY9ASIT2yROgxglHg3MH5GJY6LpOWpX3J
RGoMew1MoVTrIIGLzs8AAIQS7OZSbR2Ev1xXe2Omm2ywFJjRs3ELOFenPNOVhGYM
ZwRNWolYmI3QYEGQtk9FZFUoYQAHz1TYQCrsaqaOAbk/JDwwoyo6nNZUAKwEgupE
YRPJGGd7DZnT3I24ZwN9lQzZBDn7mj/RMtJutmrXgVrAlReiszk8YoQM/HK9Q5uD
4anYJ37K/6B3W38lu0vMz+8SH4J7FjeJN/wLWxKwE+bgbZiyBbUiJgtPLCJsDyv2
NQO21zyjxuUPx5B4Rxs3FBWPmHMi7O9htqtRqGS+uStGzmuuHPO9K19+yWRdIfma
y/WE/BiK1NZ5YJCfkEzyinGDUazKZuBiE29hEo9Hk3kd3wSDK/QE/JbxgG0d9sei
ujtoh+qtOxhdmxq2FHHh/B7UqAL/AlJpbRNptpI8Q3c1FFcSrRxt5gh5WNX25sVW
V7cAuv1/dfqkRouN/TEy7OcyWjEegarNdf63Yhihk3S1rIAK6yA2GIYwlZT2wo+x
IJdsW01iWNQN9F1PMOgdxqP5+JkvMTCxskn9ApzL/qtOlIWitFKpOwYQkvJWZ59K
7m45Hcex7kAxFqcTtJn9KZGG8i0yivt7VjQPw4sg1c1HdR2CUd3Bt/9M6ALk2AKg
O1EZ0s4YNxfFZJavZaAn3HTVBO7ZoBT9ge+xP070GvlfhbTPY3a33xH/80kXiNNk
fIA5NK5tYHHz/+OSMmLPDR4Bjh3umdeYQ3tBWu4prYsECm+/bjiUI1yCvHbZwBJJ
VDjfgxaa0HWnegfIMoRSNwA/h1ouwaAXIzif0gca2B1PT+J7PwiR8dwOZxyCOITv
RBYfah2wO3DnM42wS1uCUi533xMdhp0weY5gnVOB7N1eWgAzo3yTxZQk/pB5kKNV
yoQJjAYBzV40mCPmeODqU/v3HC5qrrDkLlv9EpxPy0P64waAHH0t2od9pg3TV09L
BuGimk+6GWziqBQvtIIcqdDy1qnBg3ZBr2CQ514ZXlwvJoOGcLZuy1ATWZJI8tvI
9As1Mcf+wa7cn/x50QSCZEQpddfn9cz/yOFiEXZa2FZLq+Y6TGezZA/C8jA0TbXD
f1tkU+MvOid2rfSHoODChO/iuALgLlrs/cBgeh6amGEd52fng038slw4AO9F6eHL
FGI1Ovqy+fERO7o2hBmem6dG4uURWW854MEIqsI+0fiYL3eLWb9LWtEwrwvplGca
VcitVuHgk3XiFkJSV8lt//JGa5u2HDplVu1jRgLIAPOBHE41HD8xt1k5y+KtHpTz
DKyIteq4135kJP1uOJqVy0dD2Et8sN2zQM/bCloqrLSqtMrdpauyAjgjMx0ffaOl
oeIDwGDKELn3uZ0DWMJqDXlNL+ERe8Jl6ggaECpjdhfR2kR0mWvVFLcy5+ZR/IVF
/rOXrJgnV7a4MmYSV9ylQ7/0Cl2HHswqzPumeugEjXKU+hdA/MZ4Pxiqz0QMrydh
mIog4350a3Oi6nvIAfszpRwBRBqUNPnRskGKNc1TflYpIIG8VjoGC2drvL3DmJ22
jy0SMViWtScKTbMHgD/42KrnJ3SsOKayrBbjNGB0KHLxorioOE3BsHB+1PkzlXcP
nQG1n8BNtJCDV96C5z/vkVmDOuP5zzGd7xZgOhbKesuIbMwkx3uXqXKcxQlf0E0A
Hzr3QhovBin4Fs7zjRZUqlqae74o41CSlLsCJ4FfityluUny43CIy6L08uquzIqW
Hgt95PHtfPqFwHf7nvKsc4XhRsAsbhlquhpneT9RrgEet3sSPl1wUYHKwsUwxEbS
4VGU1gb8sNftnfBExKqwyhSXplWGHGkNxfYXxbJzwlrpno+WdONdsh208t2cCzG3
23TggriKg35ak32/KDG43DySrnJq7LuWKLKziH8e6C7If5I+QVtcYCcGEKyXqfxd
dYVUAwA6MOI7stRfX+CdzqodNxuO1hOt08MInDRVafJbuEg+MF7yNO25x+UiS8jL
v+aJcyYALAqnQF/w0JqVvjukbYh+YYJ+Jig9TkdlsOAi3PczAxcsCw2/TeAZoLp+
14CX8+9DtGOdDMbabwCGf/EMR27QOG45Ifei1opAu1VoUqhgqfLVw3eT/CJcPMZd
qrhycL7eVZYzJmBjPfIsLehbPadbUR0Ft/Kyh9kEaIAKoRAK9EJN1sqbk4UY1At2
fsQrVzzlSMzbwKy/GbIVJ7DeMDS5PlOtYtCMKAxujAVrs/Rr/S7E/9p/9RjZrvoY
rZiN3oNUVEqjSMNp4KmBPxASZ3jhJ8RTLCQ68AsYNpbuGLzsAtSFOgNO5B2lO4jy
zyeETqg1nvoG0ZniietuBuoRjpM9FWp8qgfM8BP2lWx0LGEURw43hv6iWh1JNNAR
Epz188M4PUZOJXfGI+rU6kM0oKuSghYsL92sMMW5j9vXYRJId1RtQyIBL3HQfNfC
GffPAv1gCdzNBKOQgJrFJxqARAFL5+Oct9PhuMK/1fg3Dfdqk7OeWGwyiwBm1RKR
Mvy0WkEQ63hIp7uwK10joF/vbgi5e3n4gjEKtX5oVN9TBCNjlwNtMajW5NJnREDL
A7jc2rRWTkQlOwQJi7ls7+NlfxC+54oeu2wwCJn7MbybPcNh1IkcKLSsvCUdTWCT
KjwfGdBzFG0t0cZoSJJzmYQXKa2n6JU7rspCyyL7q0DGOEMcX6PxxziOJGZyOBzR
ng/gGfUfgiH5CdzaQeCAdRyv/kr+2dHcCcTuK8epsJvllRIBYy34RX4D1KVP/qHl
Tl/yrJcCKjRxkG9GddwEWy0pnddRvbOC9QmWuRyAcEHs5fktPxXi5Iu9DBrNvSt5
xREu/BfH7nsyWw3cSQrZu8BOB8kX/+BDnPRziEnqD9albY5WHZqHTkzHMp16aHrp
qeRbNUhNW+oqVN/BtlDbTKymQ5NxNZgvLkoHykaDXmQqoTt3sKz4KKwAlZE6AoZd
DVikRqnkofgOHLTxmXMc1Akh5GP83W8FREQhuHkm5m46lto+denYmFyKrd+uJqem
2ohppz1eeMoGZA7W315nCmJKW/aPsP3C3XWF6Ctg1sI8PAnkxlEIw5VPA/JNNay/
Dibk1clFsJXT90ed8YLP0XlrqUIVe/OHLszQr8VbKoaXgbxsvga3InyhrhTs9mb+
u5d6mO7RmLa3XSbn1woS6gg3UyqLtTTBcWD2wdlmWI1+UhPDX4FpfnWSE4VeK5Tj
UaL1igKAgCBzPl8j1qmyhkLR3fCz8obo/L31GJCdECKNaDf+EPqNCrx3KVPYLd46
UsO4OzMegmXFS7eppoy7tPkczVmoto8JBlu9OxRMP8ZiFTmK+6LDqSiBwfcXEajL
YZkdX2Wz7sGRJgSrJa5qBvnOD79IdNhvzj0EBG96SG1MQnLrkJjuU6QdWsitSZoj
2qq+KeH/DdjHOkwDK0ZRv7fboC3uNtOPctv8BG/IfC6YD9rHOgckBiOtyLeAQSdX
xLLKO52Em5r4S+50vdhRc2BRUawUEZJIdIULVEFil+tgofi2yAhejcYYpaijbzQD
zm8SBcqeolwSUlqtGVByfKT1Q8R70vO6RBARyYZKitLKjRT2of7FqaMnPywO+HWl
RGR/OG9JubP+bI+DZQaAAwHk+MOLqrW71F0NORnKSU9DFpwu9tmHeOW5lDAASfi4
IN7h77cSx7UH/hvPReD0Uf3jnbrbuaO9NyJCI/mjPsELEGPt+hYITvmMA4Sk4vyj
iB076qVMkYJ7SNsvyAg0aULmwT5Ru5yRiqpZej6Q11BRVOoGfwE/va9T3/kIb1yE
SrNqYWdx43usvajR8bygLRfrLe7Ga0avbUTNrxe5/VLcoD5uTTCXmfT7Tkricb2Z
wWvJFwCr8z8DshCUM3zeEzpeUK80Rps9OhCVpGuJ4/LnpS/UepeCQGBfG9IAlFAj
fn59iwpkcV7ifj+E0wYYjmrFluGMr4Hv3iw7lKl3tN4boD0sycYhkZS8WrOBhMKc
W9SdQXnDT2JWDa/GVKZsrdd872RwNtUGpEvZdGypnpVSZ3wjkj2BidA1Ab6r4E5m
YGhw+EygQ4APMgMJqcm7Z+USNbfq4rGwtDmPlhKAoFeoeTnG8igot2ysq9E9oPUC
L4mYcWVVwnOrBkDcH1ZeOH9ES8XbHcardfrPGSVB8q+nTlLv5mmoXP/Uu6XDD9as
Ii5MR2XpKfYqXbjVh3xRVwauRJZe3yrssGtPj3FIdArKhO8eR7xoS3qzyHacU3V0
6++X67iztUPViBwm9+9Q0JbjlWRSUMijV3/VE1lMwvWHFNhfv4ytOXefhTdkZ/tk
3N9PXbE3t2W04GI0KLY0Uc8T1zSgll3yyB08EK8MvwkSDivdX2/gUcIRvGZCxHYm
aRdiqqogSCi9GyC4ObHxlgOl45lhQKK3hmHKe0hFWOs2PIIacdDOL1qf1XGOpcHO
q66p/yK6QPHBPf+XdKwqKk+RDwx9NBk3i4DrSfLfarVH+jUBbwgGhl6P+xaQsJcw
qgs2uEwXvgS4GuWu0EumRsmUNkR6IeuVqxdynEI3Ss9Skv7FDdKFcnUrjsY+Pifd
d4lQ4Ag25szy76ti8KgiBLBiHerA77lJyuO3HHCyoeLGhY2HVYX9Hb0h8nMW4BkB
8SZQJ2P3PRALKMcwRBh8/G5BxZ8bZHX5SWMLQfQet+uH+q/VnFzI3lYgCjHFp3fD
LpWj34hVC1hMJ8zrDY2/cGJK5Eth9rmadnoTepX/wW7Elxx4Rf3niepviQxMVjpw
4cy+whHbAM/xs7wSPmcwp3l87rWkTwDNIYQrixaTN8+NlQh7Usyb7cweqm9RSPJu
OkFAF1bpdsiYaHSm+jN4QOi6HX1s88kZuxgYIrdIVHrtfGOxpQOm3uA9FrsySYZq
JQFMmIXqo/595ntRbyZZqN8FDNS/NBeb0nFM3+2qjKmVZhZqyfTGJdLYxb/bKPLy
Tt55dzH8MNrWi0h9npga/wTRk+BwLjGV2NmQiN1Ch21anXkNpiesF+tX/mOPMjRq
IBT5tur4X1fzi1W2VZ6m9VDeYAOu0m+iDTOTdy3FTmHL73aKvfRwmxMNlID0RvU+
0NYJyF7LZ28YCyj+GvnSy4x2tmezl0TuiNHG3zp6xsWNznJVcsc8I+66/6wIP8i3
WJco4ly9B5P/Q5Cf6326fDkxj6o97FhbGy7b6PRDkWAStn7p/3r1S4K0lkpYklM9
tVQsvxDqcd9QgxtjlVf8FymtleaS7MmjGoIVTomUX29cNGc3xtmKeIrmaHUJ9J+/
8ECSvwLZvlvWl2pMI77mhrXdRhnTucTOAVcgaZLW4DgrHDsnv7qMRo93gEl5u9Eb
YEVwa9nUCYzKKColwRc+7mg2s6mwzq7FSGS9ErUcckxLBApkunP2rnhKnddJ4V3L
LTmSMWWCUXoZM+pPkPOjwqIUQytmFYTyOUFur15DnYWT43fUMJejGTAgReQIEy2P
w5bVpD1GLehDsa/DBS9CErhIC802yf+LNaCnWRndVCdvtUYn2q77IUsO3EHY3XLd
Rvc5eTGUvwrrTUYFGD5GaEmpOhTwetslUsnxInj3ivb/iwSzEnXfvTKM+OxZ5Lx+
Q3lL/PCof8/ZSAnJg0o27MwEgBxYhpw195OJkeHVzGWYxr8JFaNFayjiB4cpN0m9
PlRFovMbwKvpB92Aat85biB4TGLcd4CWVrAk+1JicJdBcyg0QU1hdD24XlDTrhju
s+DcJLbPy0hh+X0Pg5mrA4GcbfvhfOfGMDQ3Qgwq2xhFJPMJvE5zVkzdU1EFptiY
V5jI40fxZw6saftMdSSjjjiFJDJtoJsTsHFpsELEsQSpD986KVoh2Bl0njeWvwuG
AYhidzIeqIM/Z9gIa18hPqJxLPEZFcE1185arIMyxWqjObs1Go4wTIkL036tPzIA
dGyYYNz3/+tjgW3uqQbAxT7CROOCf+7iL99Mt2AbP0W9qSqxytOdHjpxDESeMt63
uAZubT1cbuN9vyVzDWgi3B9YC4KJiSyPH7nuKJNiV/Y15hQa/QrvM2muH/KTK7pw
ETLgCaKOCB+d0lh7h/xL19fWPCg1RHucDFJGqQ6yR18SyPfgFFKF50V7ocYpce9H
YjdGiLW7r3zkTzGe/P6jeGY7GkDNf5IZfvJltdL8G9dGvFXpYMUQKvkXyIXaSTdH
8qY0/Vx/mx2BsIPDGOnjfSvCycN9bwIDSoK4YiwohBX5ejSH88L8X91IOEySkDij
DGWHdIuKJnsTRzUcrBboQjlPVkoD0bpw/TXLO3/BLXbFNF+VvrBM/D7lv+VnTfzb
/ZjaIMafKHLTkt3bb1U7JjyrEfvjVHOhr/Far2wHXruIZnWjGStjzhgFretaJtwK
2HmvEuI3un9KCoCggXXrL2Bi/Tye8MEHZDRt5PyCRvq/mMJ0SuwzwVky2oODD31r
HTDYDDHTbdni2X6Vsn1+QVS91qiA+29qqQdIZzZLEvJOuVF4wacpA2s1aVp/kQn3
W0tOT5OmYuh/sjBayo6Mj+dkyCFlD4jQzyvvHQEmDtWLKsXh1n0NluAxjTaOcDLc
gHL+ptd48LPZuZ/WCSO4tkvns/nSHHe6TjU9RmNDakLoToPoANtxCE72WaP5biFQ
7gqd8/FXiofJJ38yXGAeWC3wkKDbah3rlgSD0+h6LqixcvTGhxCv8znbHx/0ey7M
zfmTW/7ImE7WjvreUgC38dRWRBPn1227IU5B5ocdAl+tUmcSbr2feLwCW7JbFKj6
DVbr5iJHqH98sDcB32BMvtGz3WMcePsYhA7vhsV8G7Tb/rSXK0PJiGfUz6vsVSIN
uGd7vcpK0Ua7PrMTbOM9EnBqxyCnUOEtQZIvZOqG96v2P57i83aW7MQGIjAojfj/
+lXZVVelMgEmv6iPz6iCwX5HQDA6wSPEnXuip02sTg7N7H7VoyrrX5fWwTN/7UR4
6Z/ofmGxLA0GN1/rXzkQVCEmVhE4+9GBCLPjI//uROq8zH7zxbcpZttwGUPZ8scd
1PKSxpSEFWqQreGW48nr2y4OxVf5G6GdQmZDf2nj9JqxtTsulxWX8Jcapm8AZjP8
HvMTF0zX0tbeQ8Vdnf0pmiUzMi63BMCOHa0StBtPROtKdjwsnZuKtJT9OtBbtgzh
qWieSNvYCOSZsKEa/1rfkkuS/P1Xssq1xTNGoWLjNxJuKYC1FMfNNdqv2YtvrgKJ
nJDrMSZcGgx0EuRYrdmAmpDNoNr11aoJGM+gtFl1PWmkcgXfxU/3p7JZbWaYsMCi
r92ixvTnSS5DYp5YyW6uJyKaBK3sUay9KrnpidTLlAJgyPWzGE8wVngs/t7UawUP
9sTgHjx/1TnK03i6NfXp7JVlTBS8PiDyWzSsfsbDjPfaW4DOcxL0YH/WuJ+7grTy
YKEdmKfQHThIylJQw/XR9aO09QmGXKupE2RLzdbHwkeqFwvv26a8UD+3qzmO48wJ
Al4RVQ++JdkuCVwY7FU19LC0hu34GXqhnoT+9KiLq00Z4luMDxxBBvHuIeR1CHdz
3S81FkOUTasziLWSupVepCmxThstovqCx0j8+SxkmYH7p+4BryLPLs+kegQvOzGR
7pZKSefIWkecKb9+7e5k+rs6F1B13YrbtKrxPZMbF7LpNIz3K2xw0WINBMP7tgf3
fEIVDkoqndrioD3RN9Uory/EfyH7USONpwNaggQBsZVLyLdmEyMs5nkdZaLi+tUk
JLpqg9eUlkQKijsMrZeZojY7grYnclG0Vnet/dJeBEv6qRKGKhH52iG8nG3oHArw
h8eKrlAmT85nNrhT/7Yv87NsVL+Befg2dabxp+2y0KjOyDKzB7wHhkxJd9zjXVCC
FM1F8+Hp6fbHaPuNywDGHMqJ01tKAelCMdUMj78buPa3duVnZjDgXHJ0n2qLClj+
z3sqR0OAWssIUf9lEQ+rYwTX0tkbZ+QeeKMlNZL1FbKs0QnRqdcpl0yDtY2OBvH1
bfqFJAXPHtb4xINtWy89DnipeWYL8B00S7eU1w1j1rD3kh0s5fjqYxIR2pIBa6Q3
ct6+VUfHK5JLVq3dJjTBfgVE4s+4I2uYjmw9xCDIBk9Ok9Rs0Yi95S4O24BTsQ31
oKFu1+TLYAQ/6BLg8DKDHd0yo9DHc6IAC2+3jBMjFxWCiuQ7Uj107VOKTe7ysWnF
1miaK579Bi6YGYaWh+odmkwN05K8dtZa5pRD54I08w88Qkb2vQV5QMMvO2FLXrvJ
JxIcP47ncgMu7bKvb8rH9b5ZOa2fmb+K/Y+VT1M5D7cHbz1h6/XHcThfKHAdesHK
kDvW/jqNSuPQizYlpc9AqNybojZ7rLYegPE0mE7NyAF9fzq6vSCrw0g8ENiX94wp
Omchc2tnfonbg6koaJ6SMB3uUF4cG36bD+KpH1yS/XQlcjxVFT4oD5r/7MWlQWL7
ylwX6h4llDXI4/9fubEUH+X8fYkPEL+HOrc/nCzGfQiCWHC7XJvLO1wbWD548VVB
vHtQvwZ57nGc5eUOfNigTmsKjt2A0vX3rHq6D9ojBVFcTMY/Ok0bKyOLa2ZUWufb
Km8VOwIkDjXp5OcjGT6psXfvPAAGSokfVC6/Y0CWIIKlOQ9QiCJMC5f+2Clfd3RI
SXZpsUkzhknZk1zCPrSeAXI38JiB/7jvXoqM78Q+wBgggVsFhhpZclzc61lKpl1n
`pragma protect end_protected
