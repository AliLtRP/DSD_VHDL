library verilog;
use verilog.vl_types.all;
entity two_vlg_check_tst is
    port(
        c               : in     vl_logic_vector(3 downto 0);
        sampler_rx      : in     vl_logic
    );
end two_vlg_check_tst;
