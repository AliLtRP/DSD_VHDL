// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:35:49 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Au5EBAzQ+ab+9+8TS7M4iiUlb6FrmwKMftgeNpjpQ4JMoYEExVzhR9U7KPXULIY1
J57/MOxjRSc5Z0bvrhfp9tCFDMxlZTQD2GlgdyFrrKeaNbvbIHICb53e4zXN7Mwz
z3X4fn4+t+/JGf/Ulmanin+kDQ2lZXJaxhqqgDAvnAE=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5600)
5U3FB3d+VBIgZUnho0lk63OZXM83tvGnPYfiQz6KQXBAbk9vJ4c5zVx8PTGisOvp
3K2N8/rPhojjnrd3Sy9HW1GyKVw+4ftm8npajxDlgSQXprWDWQiFbKBqsiTm8bfT
AMUxWmenqLq3Z0FEKTNN9sCB2AT7O5OsGCHVwCagoh7rpuIpdMwY+W4poFtucBkc
VBek7e8++qNC9Fp59umxcfZ7COyiPu4FXhBB8GMTVF4WuVnsELp3DM+klHy/YxBh
MbELOTTwE7ZnAu5ismv5iX5g2gLHGhH2qOqdMLhxSF0yNSeq3hchLHxZ6eu+YK5A
k3Uxjpzw9eqxp3CpZYdS8cwaJzcNEFpJFph0+mFhsqK6U6QhrdeIzhCouvTfP6GP
KPVlgZ1gGQbvWIN3IiICmxXF3nsEa1LnIl/5CsQpTb6oldD5lnza2bUA4DAL5lgm
n5BAP+l2gJKBg69wBE/DSW+3vHQcBz34RHsloNc3uRyRTii/Ab0flJE3OMZsuZ0W
uiMPwNxSPsjIeHKUm1vU+aEbh+phhrLQ3J9s0JGTZ2p17C4nc10HJerhTog2qOso
AXRmobxEqyD/8UyRzN/TT3tKTPsFwN29SOY29EjtlSHETTZduIOsKIPEw+ZURGEG
kkhMveqDPluJsZYVa43NqxtcVHDNqKtTqy6Te3qlLPkZMOM5kgqxalRi/Ym7MGq4
vuDPc1aX4HcT4AZ6UBBgMOmsJ20jOMqekeQOvfRuI5Y5WOerYz0uJwkoN4Gt0A4Z
TspkuoE6yyN1cQTffex6yNJkNylQoYmM4w0km1UgWdizYpPlNFlAiXJz4lgWGE2O
xawyIrVWaa/w32nvvnNcnyjviKga4sHt5OxZiIPJJGHnEO01mwGxva+/MVtiOP3l
9/Q1QqBXNRQfyIGMJfz+mvOE6zAMKZQlV/lfks/peFg1KnRSyq82NyVIQNU2s/17
kJZfhNqPIqZIqLNkFAtjRWTfohh6YmH9W0LIQ7ilLhvlgp0qNuTJj5Fo5NofOgpb
QvGYuRwYxgINFIROWzQmE+bj0J5Uob3zlWIj4NcrFT37jXDVARWuWIe+Oq3oaKQe
N+A/PW0MJO3Y9v8v3gK58hGhAwGh13rRN++l9q/aiXBjJPYb/dOcf5G0Dz2hZx48
srT/jMbdA+KfdM4mPfIm4fkcHlpWqaWjJHkKvHdYyYdcC+LGVfWhXGW3vAHjj8il
82E7uHqWlhVDWBcGlnw3RYlK/ydNwm5+qW7bEX+4e6OyNobQ2zYd6GndJVpshQ9W
qTbNWUgtqjcCrJMypsxeVw+AQio2xj8MGHCj+/Pqs0zNsnx2hfcUPAItdh3B8NKu
/32cMC1wGUUMh8tw0smiSbhpJq3R/ypZhMJMd/LSiLBy1pB3ySPM7eUcqQtSHRBN
gJ3SA0CRD7pwoPTqBgJ4DOfDcLIPxYr9OlpldoIWZ2tUqyCg1EwiggeN0nS7Ewpm
tgEfxY+rypW8bLcyUGp0qf4NhHzj82k/0ZobhQ9jKDDcfYSDBJaKal3+Q0Wfvns3
ylbylaAjygna6XtcfE87ae8cpYuzxe0TPXh479l4WsHbTq912EQFA+HBobQf7GUL
0k1gBfGdNiWWdeFJzrpb+fKrtVV5t2xtfQji+XJazwaHwYRywcbL8xKDMeQco1Js
PIMqvw7lCg+8JWOrymB0UcE/Q/QB9NGNlcuk1ZkrV3OGHQVpo46lK+tipxq+RaqU
Tf5KAGkxt4X0lOVTgCb/hJIGIZTdhOV8bxdNld//5bATTrIv797qoyS+HWQW7yth
Dy1WVBIKA5xVfiCDi2iOJdep5ZutTIWGqA/2nwftREzA7rKs7VmVXAEUlCOsfWrH
dYw37Pt/Cb3YvUFPqA3/VllYuYqHvWYORieVfoKf7NDLoBT4yYjdPeZUp7ZdKFG0
UrDKYuufrErVn5hxKGqukSNOSfyJ7BkhVVlPHRxWyDhP9UujDwoSA6Hj3o05jHCE
m0Fojqs/ysRgHeYd+3PmkNYPIu9xPCE0ixbv+1DP1AULzc1qlidLR+p/JhzMoRZq
049Imd2vuMvY4LBF3ABVsCb6KMXU7iAF68UZ3J19Wi6uhEz4SrSAW5HdAOqUFl/i
bAZ5n8JSqlk8afbTavSwCEWfdW6ltOic6AG5hPV66gIwpvbJnRq3gTP1e+VfKLwy
JX0y2aOUgcoui0f4MpihOgXbYFTNuQaRKOveXYgg7FpnDx+tljH2+VkjVzLUzB1j
tUu8I1C1EprenYmoVH/FnOUUvcvpOuFLt/qZyIA54PBDXYZFcOStRJ6BiYpQIbHf
uwsCPF65Deprbvn+WJ25tbcfbch+fhN9ROK8WuX+EKKPXdLg6qITiSj2L03jnigk
0IxHg6OpCD7gmTyxGPSx5GG99J634SSZenrUN5qThbb6NjPLFu3z6+9/CyDGR88y
vbtDya0Rr2QCfjYN1jmVVk/Tz4qfF3kcBOEVaSxIAUeOSk+372yg4AVjLwisrH9K
vwIs+qjfaBFhPQHyTGoUL3Qq1Va4hFFNL0QEogdqObK6oMWpdDH91uPZO9tx+Uhc
xFFLAhbVMHpNInzK2I+WT9a5H/vv4capkVCCtrMdkAVsVdtNWcBPT8492jGV0+2l
Tt5OezCiooisEn/dNysmiwUcZiLdTKrIaXufznDYPrAr9q2N89UzIoIfzE8mFdP3
JjPWSM4NKy5uhtVxfsQwp3HWMNOcQIlYZgGEBSDDlWIuB5nbs6a3pNk2+8oFQ13S
8MY7/2/ZOFm+3mbW8u96lbV0SXH+DI4Qw5J82diOBVjS3YDQRcxpdP1wApB5Asal
vDfUHD/LAAryrFgH5oQwnzPjLN5WhNLx2MceM6FvjWeOMj06Mtz9VzAfOk+cjsK0
W0bs4LuLOvcEeDk1ANuBI/Xq0/4t7Ltm0NH+evIrPSClsyyVcYvi0KWsSO8g4jyN
qJt52SHZxx/aTjQ2I2pv9kFGhGBI0WRgzwusZZDeiRgprYr03pLNGrkkgoZWu55k
EYs6FiG2c8Shr/awSy+ns6YttMofvPryasUk5c9R0gZpiaFDBxAWKlEBWjBULRAZ
KpZZjsUuVsuiJ8P4YH5pkj7IOR+HTHcKDsazphNXof/V+N9SQKVxI7kaHpg4vpsl
kX5YgNeLUOEfh4iqhhv+Mw0fZlA9x1A2vVanNzc+c9PcH62XinP58BRkpNG+kRQE
ciAW8aSbcl/Weavpu4J+xl4IQ3tpJSIAhjz/Pmp1iO0Xlhv5x+v1uGeiDrDPuVKB
dqkHDfRKZn74QdP3LoNBP40bFe+m8+E18EjIEpj5zO9c8DOs4T6MX6kLSZ6+Delu
ZzrrJMlHAqlBxPBqpXwNRHevfXs5QLP/0zl1KozIWx4DoNHPBLAS/+MMcloJ4rdO
rKQ0Wl0sQo3Q6a3az6HgH+hQyYCLMKKEyN4qogspypfx6W2gEDDyG0fmnBOWVSBZ
2/nmnm9KZbPTDxdtAWOhMEnRieJHw3vA9mXp6A/tMW47IWF1KxYRyHwSrUYz+GHF
4vb+l+cZL+CVeC7xAAZfh4dBq7QBmfz4zmn2hxkeLSMscXA58cmIN23dSk0q+Y9D
JYtFh9lp+ECif9cEM/AS1SnHjYXyywMZ4iTGsBLvCBrGDYX0GoUWSCOVMvFzsG6U
zZqi02WSMDNpNsplb9CNDk+TzCgSFLLx+OYuGyhAYgoduDXHo/BZB/dY45jBpRa4
895OEFkS+djAI7IA43fj+ThwHfKmrbtkPLorewnu5Jk1Ras9dLG6pdN4lI9IkBUI
CHxaFILdLzv+nkBl+5W8wWKdcmQaWV9JCT9Xz2QLEerICp+KHTuEeCdQT930Vdmv
NlvyXDc+x+My5MPXzwdJ/wuX8vxECdEhs7PNMIx1aT380UOWZodUDVAwhFWY3WoB
kCoP55tyJrlmf7kArzb1T+1UcZ+C/Pte2SWzS0cgyBczZNLzVXMydohD3tVW4uwy
7yAMP2MnA8umye74gQO9N3wusW3IhrVMZEJZooBCroHeE4V7PYHNb+6dMPufHLDC
nYR2qscUNqSEJTgcrDAzP3eEQqhDuc9xnUHTvijX6vlJAW2pevC4TwxywNMaqW+/
abhKGTYDvorkyu0eSU/0M1zQaSdAz069zl0OwIO4j/Dg3Y/ND2fN5GGdp6EC8BgU
RAukl530sq0Z9udk4ZYNx3jJI7vZFQscBGgfyiCJdV3c4MEqunjfJS6O3fjF94oP
mFr3AQZL/OcqZZ0uGKm2EH0JGvbxbwtTPILpYZQTBD/8LSF/Omvh8g0Z9a/B8Uyt
s0pZ7iJLGghwQxORVJcODG7Le0lH2uvdOCHFyMkNpGJ+C8p9K79WntmrgB27yR51
yhHFM0cHM2jZdZbn3PzGT63b97zQl3egbutwib3SMfAMx1DkFfIW8cFCDAE00exD
0jw9Bfw0oKak1+ar62kmS73boloeEUeeJjCVcmyAwt2oUsq28wvCXO/01TNElxDe
C1+N2P7W70hu2jwOqV/kSiIW+bPx6Dpd8eSLNYI6OyjcDu4mCBRY7agLD47hIep3
xOaaLFlZ1yezvig9uULQ4PggdbmS2WC6707FcEbSFaLpHKLqUjSfQj+L7bsWyb8J
yfLO/jMNLo6aFEMEx6fzEfzqM80iAvMjgX3BM9DljMW6kzuCRHYvqLEuVhy5lscI
Djq1GYapS1+CZBxKjA8/+Y3hktC2JNQrditysxbZ9Bwuyo4mqtC0Pe4/vLc4XLYh
L/TF4r0W9V8r2UxR2y26u4TRQvjLAB/p07x+JVH2Nk+Lu3eAdQ2lDVI3lixFgc+z
f2CWI1XvZz63zEqRx2QFi016Yd3X1ryQSIXpVOEbnYRqDasID4t8AtjFAPR6Q1KF
JTxIuHVr5KL5bIinFw8BVh/HYmPjeykZLVyBLb3ybMxYoINpexdHCE7l7tOXwbQS
UOIk6BDudSyugvl6nFrlTL4CwW/kcvPwcGWm1asBqUhSi84y5wf70HiTC0iM7hJ6
Fro5YC6LtbJyBbpbpvS00OKlEp/jfj+npj+nOBSS0cxJ/o/3aa4n00a8GqNw3LMH
J4jCqIh0kKSasIEyDIFkm+6kgDNMAsPsUrjtxi5HzzNM3LD7cZYqLtkiSs2Ce3x1
Qb57/+niryZibWa15FYl3nnkbJZ9ROgf40drFVGHQifl/2WxejCTH8lGBR6BJsmY
svSybKVs9LDd2nlYfhYtk44HG+wlVVpbJYhUydeoe/TOH6zV/kK0+yHNV43mlo6L
nFcy69wqYZpF+mNrVa2+u81Dea0DAEEPC8F8kU8+hzpeyrdsLilrKiqhHgN/0hLe
9I6YJfphQQtyRnxYFWVV8GNneUix59Yrm9VUMg/Yj/kWTeg77RqFQCsYkV8Cjgsm
QRp79rAPn1jFsXoGLca9TcRKbkOSJ1KB1dQcec9bFwMzVzm8/rnFLprdoL9pb0w8
mAwjYDUoY6c+RobTwhw/MKPxAn2GSajSUTCFDOTkDaulfyQhclg06iwEIR8eXeQm
2DrAeYlb8Ek3M3gPoxL4zFjYjD485qRky+ATCcBzd2brhA7bPm/NFlXAyMJS0Gr6
94TjztvD8Z9fLmNxIlQqO1lUyBuKD84bE/IJrH/3zvnYAVUbclNxv5zfuTdU5C3q
a3bVnBsdFhcibu4z/F1+CjePA41LRdSrJol+kn4pFjte8ffE5lm7ek3csBY37aPE
K64MxgTsjPUM3NWCvydRCGqh76zggX7kvGEuFN4Q3IKlSbFVuCoQdYdcHmp1byDV
7PTBq9ONPCm1t0KjR0xnSdrQdFtlFMBUVD3nSMeLogi+E64NMJSd9NlqRC/qttGV
DsVGJMjtVcx3TArJlFhNzgYCFrqjHHAO+adzmnO/kdq5Ej22XFB1kyTDcUsIwrH0
SCeao22OxpSGVo+NXwD432aE98ntuxNQXstdf+eY0Hpn8VqE/OgXRgC23p6P316i
5V6kWo9qAKQeTcgXdNukvYCp0jOYncHS2etkKdV3uhJqaAePE5E4XS6Bbyk/zZuU
qWypXxaWKUX7UWeQql9xIaFaCMVm3hmOwGZwPoF6K5isCOrIOz3BxuIIXBj8geeK
PeFXDrBU6YEVEfg1bkL89yXtdwrJrRpuRJiIMXGFCk2U5ulI7PuruYk5rzfftLOo
ME/kVTKMTHuKUed75uUbiEroRUf508+lE9Jvsmi3pE8t8kZhaqsElvKrZ2KaioKQ
fK+sLcpZh6NFwd0FrbRb1mfvmfr9Tua+vuPeXWGT517sMmhAbQ6XupQhqdjmNZ6l
2tlet6yeTLhTVM7CUcO+0yzPYacIW+p8kcCTRBwuWN3s82dZ9TMr3WHcoS5+YvR5
KFYgfCnozY6pmhz+sEqeVpl26PxflhV4m6BuArbxx04BrtFFNihiuwYQ39iSPnRJ
AAh+rcO4aASnu3ekpuaFJVOfXXna8ILoP43KVW5qOzJv8GL9qG+TPAEzj8vIHpKA
trrZPgsacoERvOIX7h4/MvfzW+Bhhv/F5L3BjIFYs++tusevJt0ANO+YoqHOLi4E
6XRZHfcKRXKlstWH2ewAZCl0LPo3NTI/HsxCCrST4ZUV3ZePR7nnCyQmXE3Dk5s1
deBdgxLAfIlg3/l6iLJEtpDW8ovu6aJGNI6QiYmhB6VwmeziI1iGDI4o1UJgNtpE
Wd2GljcjABts9YdAwLrTk+cpAiLeShQZ4kAAG05dYrSZpjVtL4HHU5BaOwa0D62C
9VRtXx/ljKqEnwxrKQp2Bl/VEz6D6FTg4Bi5007tZ+J9cWAd4KxgBmwyK9W5W28M
XIium3Z5Xnp6tXtT+PLRMLjQoRgukNP+stzW4ifS66UUrbTiWVQZDtLyvnFpWr7D
9Y3BqbytNNr2KVTzmNk/6EyNWBN0XujdoP7YqeWBPtPhteWrZ7fH9mz1E+TkWq9G
dhw5kDA6t0aZNim66Bt2uXR84hIdPeQVfcpRomPH30scXGzxzewky05jjx4k2jI1
lSb3VtoOlI/GZaJew5LJfMsXhd/eBlh/SS0+BrwAmdOdw+MZp7JB3+UdbX4SwI7z
fYMggpwXp4J1tVrqxKXwlOOuB0OQAg2ZX35ZJBaWQPARLzSMJF1RtwcyjgKMsY6v
ubQOv9z7ziwVAytN0OJlfv6hMaOKaMhQRmSk5UHB7KC0kUFmCAi57R7aM6SDrL8X
nyAZdSdHCzBBW0HYqoVRGP+FVlEp146IfUnRP8XRPd5JREsSYaKgPMmaL3ObafyU
4p7Z0KMUN/1e9ScVQJjVOzBklnvrY8/S6f6IuemqCf4+mo72Of3ShRb5zkpxFMA6
G7WEo2TOB5zdiGL1Wme8GsccHFpggAJIdG94KXKlxRl0+AlFUM5sPJGvxpod+Zvo
P5gLj95fERAGnKpABeRKN/m4hMprEEAD3EOmloKYJkbeGJANgRbeZIwEdjNeBxDC
QKX8Lpy2wj1c+pHiI/2YAG8sMU/qFYIKc2Bf5yBx3Ps=
`pragma protect end_protected
