// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:37:15 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
eHWC11YxjGMBxvT3QHkN5oCNsZ7hBK6fCd6lTv5OsPvYRXpIXuSxeWdxZzGtq0w/
wtOpi1yM4boNv830LXJnFCWMwVxEs4L953NDxEtlxBU9aPHcdHzXvC79/HWXkGwA
CPtUi8jv+U463Q0ri1GCxviNmrmMHlqhk7AwgBhE7Uc=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 12208)
j5YOb7vlM4LRgYkj0oPOpmGEEzl/0eS8eekAeK5kKKD6rD/WdvZSTC4nRLUzvYij
fINlS+EEP8Um2zG6rfDgEK/HWe3mXH1gpXS+WJwknzRCRwA3cqsxSmgR+GiDE9N8
AsXd7uxOKBywdYm6uaiXW0yTEXRA9SB8VFT+MiVqQ8aXDtNVoBz8zcPxxZeVcPM5
I9wjwwM0PSZrna+6aw6NlCq+KEbW9AacsxYAyQFR27QZa49mZ/ZPTr3h7OzaWpyO
fEWyBUA8AAbQAyVzGJ/6AYmqx60kYT0VQtYJvMqKhP40llgEocGmEIkOiRPtFKXd
Rc8NTNrhHjrIpTlsYNjIbKEoQfby9TleHZtxk7oGX16KOxaeSuop9Rx/QQAAsO+F
JBeAZve2av40xMkmS8GAoqbhhu6vUTZyDIcBBTFfjZ5mPF4MuR8iLHBpjvCh/J3M
nXLiQqky0vDl/NHQ2QdotIZ5cAO2oDgw5iH23GxWiHcTpbwUYOkXMLJUMef5N1qv
CFgf2p78LtAxnOzm/YhajJBXXAhcwPAtrkJbfnaDtojk+QAgkrTzTkYTnIOGhn0w
lGejd7fotZwyRkyVKrWLBiT6lfjHGIUqQLU7yKFnsV4wqnxw1aYtk8z9fTQ1MkzD
WH4liIrqTLg5k89ypuk098VVwaIuHCNVpQ49w213CNASwlhU945Lgy8uhkk1x+MH
pHjtEU2EWXu2DYzMx3A57I2jTtL3fqOgiwjEzb4ycJZr5PhKQU4ydkPTUDvcXZrS
6dICq8wdIcNd1mEtM0e4mf8BrXn4puvnu5icY7OEk2s6POZQ7oibUA1a7t/Ku+43
PDofN4cle25haCBF4eOysykBK2WBD8GG83+bCyF6szSrrWGCq311scjVjCU/OdBz
SPKNUJMP2sLjyR6aZbGQ0nNH6t4qc2onlSvokiIb5KJnUu3t8lhf6dmDQaPQrnDv
9Q4/KKjbhIpa1lfDRYLUSycMAS2aSnFxh7p9xhv979XYI6qMADH4egY7qx71rtIK
OHvebpZgLvD09v/Uidn/niyu7KnNamlE6DME+PXehvadk42HKfpWRPnKHX+lRYfF
cxRBep+XVCCj0JasKT9sV9pnq8CrM17XcUp6ayFArOCX1C4bF0ddv7YvrsGyhBVm
Ii4QGZfZ1TUfDu0c4eGy4d3AIxTPyk5hWx+uS6UCiVDE3ccM7nXK3t2xuWHMTxGF
P9PTTiFPWJNxtydruYMb9PQrjq40MCZ6ovT7VijcI5EpDHty6R2pckrlPfvF8yxg
0AoTX4lu4vUA2ee07sTBhRJOI/yHByLpnrlQOMic/uUAQFqzfM2waN8OjNgguWlO
xB0jBoonE0zry8zvY76lYs9o8FrNAF1fdalMoGP1SgIMs06cBxzAsK5uh2k2/03G
SDhIfoBv9ziPYi3WAmpi9JJv0CWOrhxmLOLWt4HJAp1b78w1lUvMdKXik+jB9ysJ
xtu9eG0r2D+SYNVAdMbGdtdvumboRkb5U+LozgaiPJdgX2P8W2ocqrX/0Fviqrht
AMroZpkzM7JwjS9QFQd6xRQGC1RDmr58lIgMw432vu4RIeMieIcwlJglW6GdrG1i
vE/GZloHoLRZ4qssm7uj0LkjT3BSjnLzQ19GTj6zQikoWMl2erKD4/E6Qa7Oltjj
Avy43q8A/1cHluPqtzHSNGDs0f0/o2ALjsDJ7oyJ/inOZ5taLY2n+e8xkSb7ClK8
OrsR3xeHfeJx5pH6F4SIuXgVNnYvCJ36XXYhDh3kCLj5ygHDqkNJge7J6ZwgMYXK
nXa6ZtKcd6ZlPXWx5gcMvXkTEdwwUvgrkW7C62FWzJinKrjjefQaCRoCGuUCFqe7
oPAELlE5+DqvGeBodoERghx5XQZS6MApqzmKb/f+/2XWvKZ9slIfm9qeZDD/th9F
ESrD5gXnyUhUfxFDuYncBXbPFGeqRuj9lWnMMLmxspYV2wBjfHP+USyOSbaeoD4L
pjGENpiNczi1L927L5fu7DFlG9TCHVfPMB2YNtQW+9/UiH8NVuq42Fwrj0v4Uj0h
4WI7Y8VnfBypiFAknTdUf0Uxtn31AT0bhs8+CgLTqB+r9YYJBlo2LIKT8eezMT89
sD3Y9eh7qslpoYF9tt1/PWB8f1bceuHifZDvlUuJX6DMJVhzW6sxgdRnzl1MRL+j
RrVGN94CH4f38DyciCfI2yH0GKpJMVLm/tOKuNLEUNqaUSBkBSmSuc6cDEdPyKL1
lG8MNzUt+tF7jHyFoCfB8hFZ75a2L7GFx2cWlU99tuHsDHaPYSqXZ7Ah3pHm6kfW
tUIypTodfgQsynokelIl3v5cwXYZS8/kuJ9cczpWJkK0AOUh3dckrmxvYF48zoPH
P4t7zbkk5bKcsIh7Jz8/jOlHmGbpdAIFPmKU7BV1ryddDKkZTHJSji5NA4FHXOyt
wCMq6hE92iclAyh/toHRDB9k0PGMUmMjKCzWYUGl3pZFckk55CTn/3FujcoNvvBf
RW0T04UmrUaNVEboQZ0gLTWuyEOtwSGf7YTKnV8eALcWhBYq0RMbn/I4pGW+hi37
UikIKiaTZ4kxuMZXHWEk5Th7ekvFXsgyJiLwolIJnWCYAXAQVGRJCx3ZCJ82ZIm1
4yhjrRIzdsbEZwGh2ePF3qSf9iTiTM2L7wl7I2E8XK14vkHSVrdgNs3svdU/et8f
PnNoX41GLXB2TUJlRx6nd8KSB1nwglXv5yyD6fr2bFxb+xIWx+lPFAimlqOJAk1v
TI+2KV4eMiTC30eTod06M6hmKdcbhTKcVwzwkTu8TxGdm275WpF3SEUrRR67Tf8H
+v24UvH2R+GFeeen1Rp1sWp1hPpXvlcaXW89130oQsCeWdSDfQBBZER9Xzhx9qlm
TqhqSxyPSvjYXqPnzf8RNK2HVglMEktLTaC5Gi68IuiRfRWGQqtaO1LkLh4k+qjA
EsOu6C7aNZyX2riDcF7ON/GzO00bKmawnaRh1xx+bc2gN5lK4NBQvCATI/HZXFvF
4CFmW5YRzrr3QFI6yOtmJkT2P0g/kj+vMBwcpdmn+RQuUh2gj4I11RfKRO5ll2jW
CcmcV66/J+JX+BqQLbEty5ZwoEPpHJMT0DMbYVay+fFitdpKH72ru/Qvydo+zLWn
EBiJUzWDVvkhCUzxqAvLtgATseFvKoxh3Y5nkPlKjZT3KwW3AOc8RxXcEW8EOKn+
O7lg8gTHhQEhaewc2yUD+WUDpzdZoOLwoUfG4cxk0aFrx8S+kKtEq1DLzbX7NvrK
N1rZqECtY7am+fRoakccW10TZ1G8PXVrexapK722yTIpy70m9tqvcSvCMAYpP5F4
bQw2sgJbVmUn6WgZsFZ6zvSrmHbEfXAUaboG5ZpJdlyhN5i7TV+FFNFPYnutxB6i
BiUDGul3JV34qxDniPpTgM1TD0yzAYHg3amRt3yW9Eh7Ic36pToXe9gQIVxcjpje
wH/gKEHvvN86Vj+2/Ew6M39PrfjgdhUyUadaz7Y3zIfO34wU/MkFW41ZzQLlUlM2
veGjwJAYOzak4N5gMVoMWYZ1MMj9ZomBgpvLMrFG+tECqGVhpqx0xqPDT0P/dRQX
qmLkVZQv/fxe3XRvZZ9FoG9FlNT7PmKoeFxOKLt+155n9nkCm7rIKOG1JcxptNPi
nzOmv7Ju/mrtn/ylsoAVW+Xcwq9TN7n98kNcDxBNL88sSkBcO7RPAQgoUrOuDSmz
kMMLXElxljh6EPVQjsWTFIwpvhRb1yfiScthtitRnB74gX16Y5aJVkt+HMRJMWSR
TkEEd3vwQWNjhIshPHGUiah+84Z815lnyfjXVKxs18rgL2urZcI4GzHwScjXyL/Y
l1oi85IavA+QsFd/eHbY3zri+BAKEB6NegFOiTmcpy3QXmNIR3YppSHVAcXIzZN5
IyG4ATBlF7MPca5vynZFcTGelZJrQatTYxmL1Y8XvkB2homaY0dD3iqiGH00QEZ7
KjbcGra3bj3082fwHa2Lp7t7V9umdoYvOM9ykb8k0o3fW1m3B2kQdeIaGwncoGqP
nH6W0rQoG43kYn4LJuxs82jPnQOWxF+ecPJdpzgm8qplor61LcRBYpxjCskpmv9S
Y9msCgWDhGrChme/g8sPVLajX46O5PvVCQExkA777YEN5PbkB02xflajChmbzhLy
nLJEadKCI5RWL2bXylNTAGAGpOGjrnobsu+37feJBTf4r94HXtAxsROYUwa4k8E0
Pbml1ziezc3jFE0x5WgZwBUSIxBhTzmkw3Pw6o+VmpWixYR7Q/RQvEwRjjYMPidC
OMABfZx6aqTx3pVJV9S5oOHLBWdx+lREUGe6i/H9glNYDA1124/J0bu7N65DIkm/
MmgqLbY/8YCIYGpbltAyEfNHjaYhHWYt8ZMN9arlAFJoMrrjMBXgfnvFXqreIHTR
9lVzCjC6DaSh/IcxmQ3yO2+02JHOcV+ROJ0ZUensjyThPbOdJhamr+9AiusdbJEF
SgOSouIm6z8QlJ7zk+msIiK+DIobnGfm8E57UvRrWOU/TNMFD1Ch8R0cldntcL64
cFTBZWWtK3/zeEYZvZn+2Yy8WdJun251qWfazgxWSPoVG5WGCqlAPZwV/kFIXq9d
l7q48KByv7TEnht4yixdBtpTMYpOEdIlberHv4QUjdrM0RngQjESNaEEjVGSSsYv
49FHJSMeh3eXjF3mw2xR4fzWxaE7CSrKhEs3bjM7hud1aOC7W9INisKoPZk9omGu
V0TuBVGmqX+TNWyNS9TPHXFymucpnktUJnANUKpms4ZTYeIUajKPjQbUwqxrim0D
2F70bc9dBuqWIHQS8BxiLhwkag0V+YPMdywKzJdDotXrpnzW3pckGmsMbalyol66
0+XAggnodWLUZRhLsVa0XwEPiNBdKTECBuZugCnukAws9LCH4BKGJOhg9CDcaMgw
U2avG62giemG41CvCvAOR6hUXIN/FD5XuUyYHi91OLE7hFiBbVtUXZGK2ZUcDavb
pXrRKVaHso1qtr7JRjzwLQFGNASBLQ7xeov/KZf0vPuxL7axZIlbR5mhsMyisnUE
A273D7jkqNrpkjK3IgKmxebNTQo3Ms77CPS3OSo0gRWEVU2mZGkZhTDSTepzz3R4
7QGtlTqJSC/t8+4S+QepPL0X2d6h8q9XCNqd2Aw1UCVpZHF65DxtSFq1K93XKKCM
0vezn3jCL//oN/rkWuEXF1DEH0zcuGmpBL/URVREF6OQgRLAcdYppfUurS5vr+Bl
mHOo7nNLHHHu9kHttuihjKHmb05EsZ5KXAAF//uVgmhCTzGnLowssLKD6Q3PHOr3
AULN3dm8kLIzvZahGwtL9CyBxytouUMEbzMbycJD3bNvSyCk3YeW/N+LCRPzsjgh
eIkDdYomLafuctLtLXzi8aDMGeh6tCN1do64aZ6C4kxhRfeDMW2ATwls1q8dsf3q
/468Xy71EvOfVeAZCX4DCSKHFmKIz+t93499HeR0rK8mf+41kZArak+zYWxJfOrE
a0a0/o/+vs5ukxGCBKSe0h03i6bJrMiHWVNyEpQ3TKZoKYUZ8NSwWXncn12DS6BL
UVZVLKqIGq4o4ClqqCFja2THOoTFW8vxtQW5do8DpIwB0DHwhSxmgZRFG9D2aXca
sk1U4L8jdOdY0S6GqQJwtFIqLYQ650EmROCc+2nlaqodGnqDP0cUOixJkEt1ZhOR
NEulRLVSQ+uChkKo8A6a+cHqsInIASGbZnZ4m2hZVsa+5vUfada+mECVfrZiQ5R1
0dBTIgsUyyKakE5jVuD3k/beWDIPWHLfDe7ojeU5H13gYjryrHMCzbmjQR2TivX5
9RlZc7rm2TWyQOCbkgp5ORmvjmw/uJ62Eq6zhg1wV0r4gCurlBiS1n1EXTDkiFXD
5EU/GviWlULXfTBLv99OBYJHTj/KVPwG1PpLIGRDeX4FVITd3UbKQxxps1F1TIch
ubDHQVmVwe57HiBrKzYqdkcQOe09GvOhvuNDoB1OlMMTxfSsyFeIyY3uw2WFi4Go
fYFoL2fw0zTz5XoWRP97HOEBEk6MrFpdQF3Gpg2LN/XO26ByL1CGTWBJOOW1AvDD
WY5Y6ttdfOQRuxXtynU+RU4QR0sEJ/CJPs1nT/oijG9LY8VPlHuwUo6bDbwFcn3Z
IuoageE4utxeCnok+OVJhspVHtWTiFEPoP62/HwHhp7G6GdB+ZxpQng+5gKwAHtB
Sh3w6Aej3iQ203HMbFLc7fG6RT4prJxQjmTbD6utSn+R5fwkngYNxIxq1odaaU3H
/RokMDBYtAqQhms8wJY0I3IgntA89h6Ovb4I41H5wj+2eRDVlJuJPMbWyNtII5KJ
MjggHNmwty/I9/ltprf7qp5jH9NU4QaWdrZggQuixBirelgG1zFNw22zvYC1XlXL
Yx8t6EobvEoiqyv09UN5IPxwDsTjBCQuxYy5PmXMa2aV1UY1nf4sLTsXB1MXMLvD
TGMMFWfWnUFpavu5PiYdIkbi/PhnwGgo/eInKXtlaU8GkSCz3yXrYH1OZM/9KYyK
RJSpT3gSWexIMTL+sUNiAGWbvaXeksggW/HwNgKXVv+6m6sfTGFoBI/R86+VX12K
IXHqe6DiuI86neHAhTZYJAtxMrH9wQLBJcEMhUcxKEpediYwIIzD4uWjxNfHRnIg
3WMfFCG8uEylIREoc4KoxdnzX0FEkFyawff2ycfR0baj52hxwgJWFlPlFT2t2jou
amO92vVEABD9n+f76HDxzUqf0vPIRifiIRzaUNjiljhlWkUYUvUj1ZOmoPYTb4q9
IldeZP3o6EuQ9tPtpe68elOzFUieXuqK077Yh+XWzcnp6+Ycuqn5/hkaEyRedor5
6YEVKWdOC0FTRA/YE+QdaQ5ICTfhlPRt6c2A/r496G8heE182y0TTFeknKoFCaV3
pmviLrb4SsaqY1ZtBQN2AkCXn0tQ7JurbFSmphQCMJlEW4LuWAjGKsk6Kr3vdazk
xDNuE6ocDBliNibs/3KaEDMdARqqdaATXTC21XBuEdpz7ub6bOzNiIpO9bkg/fcO
PHSh4PwYX1fa9POG85vuNXmNJurYV4BOfq0xJEKFT81jCgtwaAV242gpd0ER2D1p
VCopzx3e+Ok+Ga1vgVTDscR1G9w5Nddfp6LdppuPP1LHDiUtf9ifdiu+28WjDols
x7vEChKkFc5OtRNuqNizSsXBJWXC571n77kRA19sDCh5eYJjDg+//HN/GdYtKaVb
suD0Bfa19KhO1fUeOnEa0ZFbw8IiVInYWi7MmzeCcBQMqitK1fLBD+xc17pwmsY1
gl7Py2W1p11I6YYjQAzgqzmjMrwMOl+RMyZXpoGTdxfmsMm0JuVu7qhZtNdeXlUX
mv2ohIunIaVWfcKPvoz9YIlVKJshssqLk0qYesOsl6182OHJILwg/CLpqg/qgUYI
NMQlAtv84XtDPvgOEFcdsyjqSI4A/aQqQ9/PQFzq036Si3f+oLnOeFL5F+QK/tb3
tI7EMyS+na4o4Y6CHDkFCE2EtLFVjkUm7vwUnxe5Bn+HO2ZNztFlaPIcdWyR9/UK
SNUjGHUkcnjyLphbutVZ3U522z3ZgZKt3tODU6KQqjjiuGvORquKFwBRUesDXY+h
rdv6NOQwRfapjQcuLBF/U00ovdnj2hHVmt1wx1s088q/ZPzGR0AtlM1DSZncn6KO
Y1PG6z7B4NACQ9XAmwuK7onuHg2tt6jl/k9GJnMYFuux6Y1YidQcqXLdpi8A6bPv
nSwbCgnKcntA+xDbWxRn7LagVDN6YDSn2RJ0iAlXRBkEevMe251haDU5gesteT2J
t2NVD8GZrwv28npN/k5e2SmoqTPy8wCMkghkUSaeerceA9fONivo7Fg0ZR5eyNgt
3UoG8+Y+kk7IueDylSfMS+N0/aGRmuag1FIp1DVR6MCQKnjULuCvpmgZ9XvIUW+m
qHS4fn4TzfLRHnu5QrQ47E5jycYgATZ/9jb/n9KC0C6MBtzolKGDZWcV0F+WfWto
LBGj0m63PTE4IjY1e0n3uyihUoRC2updCmnX/sK+12KCOnczQ5D0/kAoycdRkR+z
8jZYA0n2L4kmZHSvYCqo3etNbamIaJLcxDgVD5ytuWEzT1oxdNLxXm1RqZDVtWT5
Aw+lGkWwQ3+CNEg7X/DcTIWRetcsMCAUg833iMlF2UfBfpwnuG+vtOrZoveeTov3
qGYmOcNVk8/YSr1VO+j09q8OVADUB/dAa/bO5wgYr5CMh+KIPX5VeKmx2lR/x689
k7Eo7HS8zQlfnWubr67xTodVDFFVenucVEwFFhW4lDXQWVzF/atFzdWB3PiHnEw5
Wb2nCUzhDLeByYTUuqgCjA/RV0N2RhTa3qV3utHIiVIT+M8PwK2k9n5/K8cJs+NO
k+z5gkwxEK2Gt5AVEOnGCfxs7AYiCZJz+TtP2QpWousKqnRNmKxSxwXikMYGjfF1
/54e/f+wraDQTQQjmw5N3yNVEt+Wwl3yEPLDoZ9e7MG/IxEWTNowcMNm6klxGASr
JY0ogqHwUVWZBF4OMcZvLcLBsAC1QUCHVTIs6qJhLLeyEky53uWJIVF3Z8fq5Z0W
EIoE6yrzoFywBjFDUczDnsyGqKKhx3VxNm/xFS4+B29mr/v9B3Rmeza2F1VZslGt
aFcrHnmWMo/QsMGLY1Z+SzX9bu6WXso5qhQDVewiotL3B2NO0Bu6Jec5sZe1S02J
23HjGHWl6Y/HqAw7qvziff9ryUas9OXrh8qncaOH6WdQbQM8VMX5EuNLGXoqcFBf
D7MWHaT0Qju8ZS/AP4qyYbmlwuVMnfMnWi6CqJ+Y+3FMzN7kKxvhE/WqM67l7pG+
rYfut2981iW0DS9xVCe/DLyfubQyJdqE5YIytLGm4fVWrBA4v16QFQNtyu/sQ9o7
kLMSG8uISKtl0h8gLkjE9XUgcBk5DcqEw2IFXF7DXyKN38GSBmA5XwQ67MhM9ShW
Ewz+/37yGRiTkxxjBFcWuzwSNp/719cfQkDGVkBRJr9OMtTm9+t8B579JwBoQzLP
LfxV/DqfeqdJtUnDuLz3e2ZiIJy09xW+TupQfJkzsXE9aRcbwKl+3/ci6xH4ZJAx
TCqqSe8yPmwGqJywgWmxnDc0kZdBR0Otv9JH43oMZV4ti53mGKXr2apUvzMwvgRE
QW/MBg6Z61a39gwEqG+vOPk2no5ubKWJrh0MM9HfdpGL3T8k8QUeROE3RZ67wd3y
VEyeAvinCQLxdR0y6GH4IMspRQaNanvIr5cXrmqZnEL4GIr57ik5nNP58Kj10wf5
+jERhMkhRjiSexf4ym0ELTpn14ZdftwzfYgelAW56XcnEK9+g6+Q3hP8DsDEcKsL
IgL8Mbg7PxDRfUWiHwMYCsMiXtfMwTSwwBl3lixosNlxT5wzgzhKEbVRUSGaKtG6
/Jv9+bYiQLoDSIzdrdUsqGB/zOC3W/+WWYE0aCdIhDO5UnJNgCR1tQrEW37E+S+N
R+de1numh67+lOLdABtryFiQXQkUt0gyhANx/5aQT5sIF4KV4b3LHjWtIlgzd+2G
aBDsKjgIGRo1mOk/eS2SeuK1cjGpmwIKuzWxCM35OHtsxaIenTHGaK9KBpBHV0lq
za9x4S7dpW7mQLIjDyLns8ca7lKX4v7p8/cR3aVpsqrxzgboyrEfs81b1+/ZmMTG
OgQLujuV3ReRMVksm8ZTOgiYM24RGLPyRemzX4MQHqj/060u2qKoiE5IdjgJlveU
ZhN8ZR+P1swzaPhNWC8H8SWYCyZi6YxYu5GacfmcXtBL2ORBc7KJ6lK2MXXUGQRA
uzSo0CQbS+7ho5BUe02w6i7HCkjDZUncyjeICK8mmbDlqMqWV7wT1tPwXAuhQcVG
hGt9jJKm7kaYnxggyivmXTnvI4pDVVci5iJXLmDaVBeV3uUOYUD2melYC6RfF8+M
hBViDzx3+Dpubu7f/udBdmAQkscuWaGy0B/I0Q+0e54VSxfhgN5Ys0XsLvEvE4TS
FKLZwv4ririykayRFyfJGkXwERJDKkhpuMYsMy/rgOjgTVH6eBRgulpxeojSIdvw
H5opDIEqac2H5Ixqvg2JY3/mon0EeIcCvQj4iGazHsnKQIMW+JJDz03vLYdIUOpL
RW75wnEb45g5BNMaX4yEjgPjeYnKYas6nV+HGzcvpOVRIH1I6EArMQyk79wmOFOh
QZnm1RwW06eePIUXSvl04iSU25vU8tXwhMwNW/Mpdk/qX45TNXvmE3rVdlmwdrh5
RRb0wYsOjyvb0zQ79QxFKZBA0YyAl64VpnX27k8/xVLnKiEZye4eKV3i+CAJZlZX
CgITsQUBVjByzZB4oiBMvKsyeigCEZjJboMUO4rHdcABiM4uR9iPOsb6Hd3a8GZK
9IuRnL3LU2iPo6ls5t1T9qiySqlmtBlgpANa/9pbdLulUZ8UBmhdaig7QK5+RAoN
UsQK6x8GOkmeYjY8bPj1MLKIdXUwEbrc4K2X+b6+JqigEhFYCLSbzOm/oFST2gbX
YIyh93BLu30Mbg11LRBbDjp1rZ6KT3TuobARmyz7d+LDTBDP3hVl0BjYd5O8Rd8m
zgeQkmqM45iZyW67XNZVnGr3S9U8QZdKtJl7UyjEX1aWyo6nP2/ozk+wdeaRe31l
PTek5uzeGpvN8xKxE5OHKPn7N9U6RqZABPRO/43QtMhnXZ7wjTpktvI7Z8AHJ/H7
OdeIFhP5GCLFeeEFw0zS3zdT/gNGjbKtz83VsEsT0OgkWhaosAeBXk15MNCQtxMw
LBbDz07PZDJjWUCtB/fFC/+BxnF44wSPpFwC1Z90AWxzsp5/1SiTWdYeGM8j46Z+
zOzMJ12kGDoN95Oum4xdHItBEWzqGRUjU45Fh08hUCq5ZVWY2FgMHONFzxM9GcDL
jv/TGXyzvD0j2PnIioJnWkZBATRu9w87BV4ga8BcOffib8It/EOiNJPYmGyf6OOk
BQ3T2oel9uI5N62F6pjCT4AfxbkicFZ0sMlItr51+QdBK7oQR87UZXL7wDev09QK
UmiNPMq26QiIFVe0kcG96DeLjY1z6RixOhFDzl6AzFD/OhJgvztbOcBK1F/61AIi
HYtsgIK6qwFYVFcV8MeHfGNmzrx7EnJ/XL8wLDc7WDnD/CcWlVa4U5jZLyK9KtJL
Edfxjk0yZNBPj/fFvV1eDaVAv88MgwH8P0HoKEJ2eoBSbu4GA2LYGBybAALA/wUf
74YhwTUa+Fh6Xg1roYpYPNzFW0yJbpii5+wdBS4/4o+QQ9DiVEgefXxmp64Zc5nQ
8xPepeITbYf2xEfu2N3ezEfytI5ASln7gHlsNjiATAIDTb3PoTyme7Ni+081GKjc
rUDL5jX76SRl02NrSP6lkGi7p+rPkipCAmIBwFY0m5amMPBAC5Kzh1MaUlfgz5XU
Jug7c3Xq39mEYgeMuE8NNvR+2/U/8v6WsnNwuZzEO399GoYyNZInYuKf3960aqHX
/wlubvryl3o8RvXCmSYZAuhZZ70PeaVMYyVSPYf6CJpeWf4+v9Gl2uDfimUQxm4R
5cCYZGxsj3Dthh+J/YwsZqh6hg5dv4WK+yvJBjLqBxQ5j3xeHLm7OubvrfcPpBxy
tZKbJYEwT9hv8DAWEzF1tbGVZRR4NmgeeaJ4SK3uD7cSw0tKfm37gt1cPxUYgQX+
Y5c0O2Uogx8ZkRsCqWUSlm3ZCt186xdkfz1HAGIskbDQWo5M9jt/BD5Nesrecnbd
V0396LTO+Lc1KDV0dDelsnd81l8a23UQAPR6koHXiJtxS7P6ojvWnjWi9BezFClC
pTiyrwKtcMenCciqDzEST+UyhoaZ2JrT6heAYtMJFaWAPuO6V2mRMAz5ujcb7rpZ
0XlMF9e9HoWXnWrgALdtT/sjep9CiKggfWzEBOX8oG7UZgLuU+IoK7+RV7Hb8zOX
OEDKyNSf6Elzoc6A7Vhn/sikbc7zS9QBSM4CCzobpYQzKRzZ2c4Zbkqba9wCEwXm
DFlylCLJ9VxUuLlOh33CpYz7p2TUHonbJ4BOXL4jjKcIhNM+e8oPNXVsQglkMOhK
a+Pn+gCkrcxo27Wm4+hINOiIPR/MvzG5RVrYdLR3/rSa+4obsc+QMSBI8CJ+Tw1h
nAvBLKAFiZmGWE1OwWiIN38zM1i/03ThRj2+OSQ5iNMtmxaNpbE7anfTfkHXLzhZ
JuidzIcG9kCTTbwc+9Qm5phmbaY1BpXQfsY1Va0iUPO5uNyC0w6HnJZy6XveKjVO
sLKpftvQlOMJcZSOMO4fsg6AWw9PVp2GDxrR3LqXV+KllCCMdHlgNflyBW2gOx+9
awdV8/Kja+WaXeuWZTELcVmxb08WuQrtsHY0oIZNgCGmtJ9e5CPqww2DSILRKS08
anHvMlE3Coweob8Bwn/Xro+SwrIvVKRxb4RqNscw5TU01ESl5VMPvbQSsg9+3ukF
+dvrwzDXd3FcPFvApnZYeRk05k6qNmCpTkGDIjBpAZxYGuQhMWB8g67Ibg/rVEdl
BYTwWcWxOAD96whjy+7aatIb9njbUiIEteekbHOs3++ScqyMhALBCt2AuacBVZoL
n45j3Eheuru4T3hQFl50n2UyHXL3TaZaKiQC4PzhalmR9aafGji6FqcQvdOxGmnv
kICGYV6i4becEZxXJ+SNTtQ2yoCTWOb6gcLW7Y4UYwRQDh65i+vwJeo3fIIO+0EK
T7IRy/aP6TwAXEFWOXi5nq7ZXKZfRMws++QzKtk0TLpWq3nLwPpE3Vj8x0vvv3jd
uigge/ziRtapauBxu7uEf3uXIg+FQAOe5hAj9sd1rBu/sIlu8kcOJuU9GjNRmbOH
OMPpBIDXTXur6Ti7FmtZdbsGrC4MV5EVffFSgldHKkqGNALrTTGnfAsl+KnysTIu
/8Bno6iJxH4BadYk1KyLrS0aeTj9cImHKNN+j145VGk5J2hVQWsbervRfjq9xUSs
Zd5pHdGSSJOXWR7ECf3UU6Oz1N9W19S9jTyufvleuxGGSMsarw/G3kfPwCFicna9
AXHhiL8n9dxHwUaIPDDzBYqPoFtprYbF86vJI4+TYvYlGooFgAkXMA2usHuvuKmr
pBKl91E+OQgqAxmWaBLFa7cbmFiNRVQgQYqXKxiLbxQDcVC3qBc6ytD1xXuImUGU
Irs0BemMcakXItmwQSJ6/fB0MbZer0cVfkue04K/UMes8PaB56Y9hD/QMdUGfz+8
rRjJop56KfL+x4Zkn58uDUlHq7sGiZMY68IBgSlMHWN8S60Nj2f/3H+7ctQzKSee
f/B2IYWf5k8a6YwH3kuM8hRgvqKlG1/NUVLDgP1UIFf8CCEnFkbQCdyFo68DBGJB
EwTz4NKgdbc4JQTGLwuLAHy8XNyWbxT/Fj0mk8DPikWQuyz3grLgw0g6u8DeQK/o
z/BvDHPU4fgRbvXMjxfxN9zh+NKF2V4uuWG+01RCNb3bHyfpSRWzmcEuln6tsdRQ
1NlFaTVYKcsN62MfAhWsbWkQen5E9S+yoP8p6xugwaKb/qwcFtSJ/0ifQl0ni177
UW5akkAB3JTUtCEPEG1/KrX00DnA1kn3FEfsE0ho80HBpvEKxw0Bxx79AL6Bye7Q
SW9zOB3zl6/xXLR6I99EII69HkeWnV4pl/NnTIxJ5c193XDUNGm3LhMO302TlD7y
5qDkLRf+fDuWH/AAArBuvkST56QRfxO7Q+gLN7s7M/pBVVFEFQM9qAlrsjACzT1R
KAYyxutOukFJIW6oq6w7GSIeNoUtzkSWKgvYAwJfM4asOc5ALw1bUEVsu0h+S40s
/HA00Gw1pn8m1Axq1XD5pXfkhK13QqR05jLNWEivBI2H/YgVVDPJRI3gAhYKmuzm
NX5scK2uqHcL3r24poyhayhP1b05YGrUnMBTeijwucBvcsjuRTf5gerETw7gVU98
TL0hNdZGm1rcsqS+Z0OV9cLAGBFpsqT6UZQOhvMUFl5UUstwyqINSyGVj43z36PI
olW63jAWv8es9eZDh53HOtflTgWediiWtToIlJS40mNIfPVRmd41tWysjW1NjuYJ
ePnqddzMOWPptsTjch24aPhHjJ+Gc92zhptH0NEP/04/Jn4lK9aZxiC7VkymqMU+
jo5ZRtJdOkQeT8Bt3g9HZ8a2EFY47Qa+P0H1jqRNfj2ifCqarfJzVEU75kdZk32v
Q4ShjqxNRdDqJ3iN6nZEIZTDFD+TTl53NHZYZezjV18XqCUEetDqszDIJWcPWfeL
FJhha33j9RMrxiAhQ9R7dPusIddDWbFXy2m7ZofJREEe+6zzMKIeXeNI6c8bto69
G960N5YxXJBldXgjHMseiMfwhJixw65o0eolssg5oSvCVi5aeusIkMwOF4RXhzv3
gW0HHtx24XavwEYZdlXmZmBifhD5OAd0JJROZcUIyXlknAC/Xkgp/cWUvVJQJLO6
aQwSieCcizmf5N+ufAMUf1EivgpJpJ/j7nl4eNmbGt1HAL/aphCTqgaoYf8Xhd1G
9yhwwLXbL0mMm0UlJYG0oPIzlzeOT0VDkRcElKIRX1UUZaPHK0tmZAWFbUGH6wdc
eLZAgciPCBvH9iVfHnvjsWRQcHZnbTZBaHatSIowAjghuluHHJBM1tPFmyDgU5Fi
g5CWKI/SjTFwXaq5xyTfLlrawWVrvtm4+pQJSYjl5tEs9rQVyKJu15IqpFX38BeO
v6y/K3b+MJoYoun/tCa7RqyvgI5oGrS4gODl86X2G0Ex2dHMXpfv5bdWE6DvO8RT
2FGx0c2T+Th/esu+oxg9YoGl7QuKuw+2JViH/3k+kTW3ScBRbDf+44qVudtSvTmt
t1xCl2NdXSZW8Fx6bUSKDN2WBus1OcG0ah+1+NcMD8GpAwPF6W9t6NnYug+EIhhG
YfwupvgO1qMRzLl+CmdGHQaCXkKgif6Be1znYEM1Hbl4Jm2nx7Y+ZMaXGG3Cma+2
XYBm0o42PmzoRsPqIR6wCbOf8SpswkF81d99o+GDLq/nZ0kp8d+FipjEjNWEdtDG
FnWL/aY7EB8nA3ceFCDR32vGnXMWv/YHrL7yBcCteiMWLqM4m/aczCggof0u85+G
L/7qxLyMjqV1cRWYfEZbgbDKK71uY2/ZEfudxciEy5VXj7LJYtTERSYwmwFhYtp7
Un/BNaSqOqtLoX+aAtS2Nfg5uuYezugEmeNpS+CuzjYsaFkBPc/cNBhwlKgrTZCX
OhywvVmNcP4Ax2tURYtokdwHAILBIQshN9DmS8FBAsYe8BJQnojAQ7327TpEKc4w
oZAi1wq0F9q2iMi0ivnlsRkWpktS3gR0tcEsYlqwIcqarXmtDpKL/RcsRsuR9+SF
mIVr8pLrz6pOz5hByw687RhVnwSGsxLjuS3P0XDXK2u72kcqQb1se8is719cyy/9
165MbxOtfDmfmLuN9HxpLmm4qmbFnn/KmJ5QGN8aukw9J6ljUcRI0/w6RCDxeS0K
MvrGHY+khN2NL3R044oo+qfAWX+M3iZ3ADDFRxr3U4EfwnHK+uuGRID6JdrDIU3o
fR26oogQiU1pAbGmQMLsokUB2Kboi38IvIivp4+QBKNFOMqtisiqDVV8pSfPw1oZ
5EAoUoo0JpZukW1fgITxcWAQ6FPv/5bb7qxZsDRncga0XPd7RBT73IDNQXdKMG8t
KQpTAvOOTCsyUR4G4y/RPAHq+LJ2BVcUXeyX+QAOhPF/d0NtSz7Ym9eUtfSLSwTX
Wef3Cc6bnmHHDp+ijgMlefECbftt+GEUqFy19kmWEDr1yWt/IWAtQ7oyJPRfMIKf
rrqMbc0ofWLdML2v6T8eBjb90QSYSFzNPeler3nHVBshkGzcgY8qpUxfjNEkU4R4
/tS6nb6BZo2+uKhLB0OpRG7F1WzpbULlSqRSgNOoJT0dRcrCbNKRKMBqXrTFZ1Au
C/e9QAU6weMyIIpbDxS2m3cOZWul06IOd7P1cgNAHwSc+VF/zaqwlqOaG3C/riMe
vtE4/WgyO9KukTwbLCmu6By8aTm9AJ3d805Y21qJ/3VsFYZrR/qbklp4k4TzA7vR
mXXwBo8vrIdPew4kYyxRLmCzrzvf8h1mGHgwN/8K5mMQXIpJyd2o3TxFc82x7XC1
cxQELGpjNctAfsWjM4Kzk71ALb3h9BAhXrNkAifbcXrovOtDREizY57yoECFOlNd
AvYw85Lyp+Jl9o4WlrO3p34oJNYODTSDsRGB6hIXwzPv34vM1B5tyqchApSHfe8+
QhS5WHhBjPQwBOaFepkQ+OxG9ZS/8FYrthjjOtcvFoc7l0IH5b9Ex1/PLq9NieqD
bDbgCeJEjH8OXUyRzmzcZQ==
`pragma protect end_protected
