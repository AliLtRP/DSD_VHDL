// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
XSUnbnM48k5DYKcgO0D1pJxys9rZqEDbDREenPeFh+0v+q62qWLZ/MHxV7HFMKsnU0+Bce7xHTNE
334Dvj6XNUWlrx0UdlE1+wUJJO3h3WdWSTg3Ev/I7Z3gDK7y//9vdoJlQ0IGi7OhPC8noiMH7TT/
lkt8hkYm+ze+sTm/s+XruLziys+xBUk0bum9AZZtNE6B8/6ZEN9wnrAu0khjwC8ziRZbAU/VwQTr
BSF3BjAsTx3dInr6n2KXWerI52TXfEOMTflsd/b14xv6hGSxD9grku6t528wkAJuyHpdCuw1AzPz
uKYfgwBCG9Ovww7623rMH2uH3fuyUnSUQqbjtw==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
02j+aKQGtv3m8uOD0XASRqkdY7t2UovmaFn/l+nooCmfVQKVcOVgxn2WWa7dEEgsA+rNKCgzlUeA
wdRO2QvN88XWh+VDToWjVj66sKKpiU/yiZtNP4pmSxk7SVmG7TgJJpk3ANOitkw52Jn8sfMLkngX
cv4PJWxCiX6P31bPDL90dB/EIGSmJlk2PwAEHdtw6tEWK77scgRHRC3SF0Z+tr++N9ctFALI40Jx
LmEQLjFQh/lyl22fvErJeL6S1eyP/vfDJ7BMX+nrGafszjOV7uOzSZ5Pt968J8DDd/sP9f+XIN6c
MUW6dCsq2078czt8iFmOV4jqwMLaMu1W4ZeuEJXByXAIH3bg6HC/KS1MX4G+DUiT+kEE5moTZJdM
SMD3cCpTmoaJExehw2bBOeKoqbTHnsW3zL98p6yx9+ZAeMIgozk8dVXgigV4WCjUwEYKI0YeVChZ
7cWfB0CQarL0zBmXHbtpYkl2CWbCfDLlQ1vKVNigulRNIL4BV8J2/Y+V3TCupm9qfN/TODwjZ1MB
NHdnWjd3RYd6szcnWt9HS93DfMweoUNA0rAt6VULgL64TRlV3UBKVdO0uPFANuAk92kNhSUz6X1c
WotFy94XuL9Fa8z4uPLTrGSGF95H6iyUuowYXdWq2XXrGc2f4ox9UL6IWjkY8nkMuaDbb+zZd/CK
9CKACiloLYj+TO7nHavnTvDolIu20UBFLSObioew2SoFLSEOReOFXdSavpeOdakKpCHlmn1jbKGi
1RABdXt0t+vm0rz6IAiy6GauqUC3ghjRLtUvO74ik+9HUatpZA4VA1zbdfC8hTWhNHT1IdjHEAT0
LQSZuCYWWgnXXAOKxVq8m4kVLYXBbEwLsQLuFEizZ2f5HXuYjCIqpwNMVre1t3pRdUyZuIaAwtEf
8qwKQX7glktvRB7BEglfKpqISztq9Ky0jkQFpgYGsjWMLVThsGdVyczx8rZVxn8uDa8JVAsv87mb
xSNwIlDQd3CaGQjSfv76DaW8UAnjngbTK6ZmpC8ZP53aMqe6pufrAeqVKE4Xp/X/qAPcAHgklimW
w43cLTfH6ktyvrjVI23uRypdb4fJit7HFBcsOr45DP+WsT6N5SgZrfZAOcPYc15gZMaTvw78DuCF
sEgW222Y7zNPlF/BcPv9VspqfueBYHgOd3AEgALyw0LOiL2ePw7omxm+LW+MLUUqS3zdcOV3ZpNQ
dNUFCrWfJlilzvkcFvw/HPbGrf/5VndSgxgAX+Fo3hIbs4p4lbK35HdHW0frVUxRkzp8zZwaz6Jg
QNt5VJ49vc1hFyrvDvNK58mA2FqamPR8Xg1StkZDmuO8JtqWFRjH60FbEcFRYPALa6XtGvf7ADrP
Na+MQ8GtvIEpSeB6QodxsoFRZ8pXHFr0UGzw0ZMxGpn6ehWx2eSX99GWWSCNpg1e78xNZghwWb75
IrL1OG+6RozGN2tmGII6tRiGFOvnWqn56c8Hj5cz+L2WbbZXCNidavnwFW2bCOJX8fFmmarq3vB1
PTedrpOsxvMAsj8ASvS4OES6hDAG/pqSUuD4DynCi+xu+5Crajo91ZIwVZ5q2OCDbaE1elTG2U5P
xdyY+tPfGlFoYWU5F029fihA/yra8uFGOYMjc9NM0KjlGJ2zN6iJ7I9HQVzkGDrXrQo1EMSzdOda
xrYnexzZeno7qG38rzssDc6sr4rCE6BWkK5oN2MlN+oMQJV/+/1FFfkSWb3gyDyDsjSQjhjl+sms
y8nLx7NFMizU7nH00ycFc41pwkY1t3HN01ByPlW2DTVHga9hjrJaReMy67FrrBUM6WhT054kutpv
meVP2kaDtP1uoNnCNqkwnqmYQsycxHGFOWXpWx3Yy3fAJzqeKeXdQY6Jjp8AoJ3HDcuyAXB8Mz+W
4WSJr+d3QEjKQUuZkxDswoifJmRxS6G6+x2syQs1o3Vxxrt8NcXtzgSWBMzyKcPf0DVrDscbuPWt
oVLfH4dL6Cqoo0iW5aD+WalRO8VsLgd2VpicnYm5yi98lyELN0sy8m6ZX1ZY+n2YoXn/XAmmPDJS
8Q9+rfAgmpygFQkLtU6aq2bwVgOkoY6rPz4tS5mxADJisY+iGyms9kPG/UDrOEkQ+UqDq3NnzOu0
P+B6O8tE1eU7QQHN14hRmTKRHuX9fR7JiWMrc3HnJRzWkozQbpmJtvVMCPKm3GgHSsaSZLmxiu8d
CP9Va1W4e2JbXlpc+c37SaYweBs06J6/jssd+A6mnk5RumBOt5RKIqk2QthDehW3y1kt2fjdEu4O
9jOyKcElG7Zg6PxrH7iTfCzMELU4NEtB7Q5NUzEUIdP/Twc50XraVsDN5vicAHFzioSkE0JzD7W1
nTrQeNnZxGefEGLahs7h4r9a8PL7VHgGUbVAHQAr2/8jwttWDvgfRpKpmFKk55jn/nZNeueamU64
U3We2fbMXOdmUAq266ukSCqHgyw8H/k4xuUKe8hyA2m1xzWeZ90I7e97f9FQNQXHovngGZqGIcYD
7rr2aXGIor5sJOS/ungq+V6Rl17GrYqoxpWcAGkYu7Rqzobf0glgo1VaDPBFt8EY6TD5OtfSrDd0
HpKTSNVhCGpIIvK5tnv/E8LVpAsKoAmDCs/7uAbhzp6dD90zh9sPCKmwNoUKluwpo/zD7HD1sTK0
IftUZx4vimo38hnN/Xm/asQgS46ckJZH8q+70cmJ7xZucxOaSt0cAGDKj0TqARBEf+jWCI+S/GqF
fiZVDH/yNYC3BZfK4Arch6bL3Bo55Z9TTgXa5V8TE1rOvVLW8WWFmUo40hMVoXfo/hwfw3pNwXoq
m8g2UHl3QRfGSO/WPSo2FfrK80o3QQgfUzauviVtzlKmfqMcNr4OhlWyU48a+ZYi/gmO5r+NX+P7
M7nLYP+FnNILW/7vFHK2jAJQdF8gPO9LcQv7KgJVPNB7QNQjTAGjrlFi+89job2C0FLEkByrHjgL
0F73KYGJxOhKdHhiKlcU9Q5yY3AD7UVH/lGgTj4DrMCozYGC4J4t3U9lQlz5yJ7axgUoBXlfxWFQ
LL32hOJ9GM34gDsNXzXeJ6x0B+8rBPdrvObvhbNSIRLP74Tur4ElbP/Ri19M5GKgK+6L6goDfBCi
OXUZmShvPGAipzLsy8+zeXIRxPAUDjZM9cIz9ew72IDj/sHtqfaSKPmT/F6+6vhlODyT6pv6XR++
WnFWWluaNGRR/Gq4wsILBE4SqA9kfp2Hj1mR+6OMMsSdwP5X6+hsuRID46kcrMJtsfxvWmtRN8lK
RLgCpeaAOiiZ28h1yFXdAAcySCmilN0BSG74bqibE5CFhffSBpTSDm7RySaYsremXS3z7gZtjsS0
vCXnUVWRBcQQ/3B7q90UxTXkPc3qkaZMZGF3cgHV8elQVAnHjWssufngFVHotjd0h5rpzOgQyxHI
V7AJ8p/ySIhpE/NBuVoFe24HwP6vrgrtB7ZfVKl6BpTl4EeUom2pYFW5maWhRxhJzZVu3rm2WaOG
fizEUuDVkduYjleUNEm3ZsDdm7dRXGGzS/KCUqQi/e3N1G+oDJFRBsEFRm3979tE66iBqm4cEd9o
4uBYJ6mADip1/nTcGlkz3zEK96lag4EypqXTdP7ionSBVyN8Ad3Z8K0V9mqV90umjP9aBZeMaeem
emxXyZ7Q/LWpB+ZKbnwmQTVeZQ4goVhjRtpofXkdMrBdC2mYv3/fCY0/K1HYWZtm5CRK1evnuYdU
KYd0tQiswQFTlwQ9wOuUu/BqCMJSZNTGmlBoxAvbrP6kYTYKDF8pyWbCVLcPk9u5RrBWItVXd8XD
o3QHz8ccQavfdTq/yuGGdZxkDOMhV6GHG08nCE7t2QSJ5XLE78GoMjZdd3sAI1AwsBuarFu9KND3
xhDkfnqrfDBg9qYoMhuTdd65wex5/G5ICrBCiAbOlKJ+fQoQ3uHnqduAClhC6Pgp5iuNQDlG2NW8
FG3ceNr2ygwjN57CCoOvMtTQncLQPs1WInLI9pj/0lFrlquSX4AQpwU5LLxV9Sy1ikRcI5bWXVi8
hJ2w06X+EoSEFGItL+cmV7VnAKfuxWYOICBhBFNscpFF3iHXtDZf9zjTiDWI3RykTO30LhLgspxF
7zrAr8SZ+hrEIv02gWlnvgqOTuCfBe1Op6XQT7kndlseTzvojPcit4zRBkxcQvUeO5HTeNxoF8q+
g4gqqytbh0SQcFz69GUZ3Ic5w/WAzVcu/dKS6f7RTFeGJ/VxM84cK6wtsHPoPDp3Cqis6bKZ2bVD
jt4YCVvJ4Tz6kY2LyzEl5gf8cYeqvHLU7Zt4lJ2xrgGtg3TUi6y800IhHNSczn5MVmuM8joQn2rO
tZj1j2nVTEMYu/y+C1ZSzv9JzUaRaBELsncT+2rvgWH/Zm95ElCB+ZYF6xquJk8yoy+g63KOn//v
cwKwoODaMfjBq8j4MCkjpgTuG4xIpmBoBbOscpTEmG6gGERO+fzfydDQTMkYgP70taIo4l4NYIqa
pR8/Y8Q/Fg2YODbjtCiCNMIk0FEXLgtSwSBtkNoPoLWYvVvnvDoYsOFVtcpnBz80lbIhRpYHeOMt
20Wqh+HurT1wbTSXaPMJUGkDVQeu1JdDfl4tgs7xmQ/BArHTbj4vaggpNjlwLuA6L8WKkymg9nDj
yO9Ldm6S0ZcLiw7um2K/lTBFWZGs0rgTXRYniuhW7I9TW6HTUybJdfmxbkDE2bF4tHPIe9dmTXWJ
DeQLra30B/rmPNEP2+FPMH53AaiCK1yOYRuaIAywj6I7YgteoN3ricitaff5W26XuAcJMCNEBcAV
nb4563HER1takzsU35UcRCEDiUWRxegoSYrcHiY30q59iaExcfvzJvdW4UhDssPmVxkJHJMU1ZKR
DSDwcOBjmpf5J3DAPNnT0gKdMAwiP6xSD8IGnCTv5k90I2VHdzbkz7g9T6Xe8IOvnqkWEFlnN/Sb
qy40yARGeZ73I+ozxbJHeL3HQy/80kax2w0AL7Ev6VCcU9nB2vDvKXcGJZj/6vkzNURuYZMu13/U
OhMKXd2a5tGyrzqFr78ST7bVsCHJQ73QWwrrlxAEQPMgG8yxQcp02G4Aq1l2XNdJ7zL0RFR//zpF
Frzzd28RVacZnTa36RW8PrhcE2IoldtNnB2RLQJfkQec09b3mS6TM0S6P+NmkP8DhOIIcyVY/xSd
517iRdklNks5MUq0huhDZI9S/Sbh9AIwxZf6IUZ2/GrEt54eyXQr3oqndK7WbJ3s17MSCaB+Mpbj
VPpu9+yrZBUkaYJvHJpnvQdnYT9g6RdV2pCGq4PjQB6S8jpD1GNeVoAVdZXL4Q8Ym26N89ngsa6N
QDs5e9GxxKI2jNNoOLj1YkCAHgI7hsPhubk9OQ8am30qyLYN43aKzJnI0/AF8PlXH6jufHpapGsr
pDWuYD2CyOD/geb0CSX7E2jcunNFaqRJGpU8fya+5xj15VXeZJtzYxATZmBTugHRSEjVcERrD2Xw
N2MiCTvYI6EohxkN8yylZGn0SJXERIbffrngbld4510DOt8QEDjozD8lCcqAaN+ZG/SkTCUG3f+G
J3gLxwGq6CHuzL4jAvBg17woQEGhn+dBTRbeKa/Ue8j3JXu3G2aULPXCM6h19aj1F8/6LyAH0Rzu
ffNR/ggVtdQLwzHd8Tvu44KX36NRAdQ4N2XLfKEUPx4bknt+OEfj0SU45P1alIocbL1CNOrc/sno
vMnMY2sj4FB88MdlWrwIpjKHA77LTqvpTIXQwU78m23pYqrur5F9hIcjFAniZVGLKIWm6PUdOXdV
aKsH/PHUdYCgGfbsTloHlEn64u9yYgRNAG8IbFURwf6rRl/7z+V8xiwJiSg3SkDQwKonbzP1l9pA
QmGITR/kooY8nZJhiibFiOAF11CnzCaF54hUegxhQItZbF7QAQzY8P1krinQZG3KoDWWsHWqERUX
Hmy39SS1y5o+g5iUX3bznQiSCvdPsMsOVEjc3NK1cos5fSoPdRzJTv2RAWxl0ClzinVMCfx9kC+Z
Bdke4K476eXZh78M/4CSCC20VBN27C0j95h7ufcEnWDYtKVWt5Ntj8dmUZn5Oboog28ZEDMC33lS
4v/jpfJRJAlHFtZTn08brpmvzrtAduiwLQJ6eTo2yQiuPX4AaRZHkaLAp6Q5vWAfnXz9nv8MnI8s
Ltb873OZfJ3OzErr7B7w0tcV46rAz8cP1fqndVYLMyPN+29WGGHUGxn0fXTgUZ5dbuZaTdwtQibN
6iZVOjUQy3XyOTRAqHRSBn+ao8nagLj4qXig0XR+bHA9H0sakZI7ce4Mt/gMNa5256Z5/K9/obta
awdzs7LgrffjSp/OFtnXYt7aHbjTjpA9mBPLrmdkzedoCiQaQo4PFREUdq5TSdxTJTrFJ5EQ1uBr
XlY8g38G1sC5EDThzgJ58b4y3pgMjFdKSkaYl2TsyMMYyiggrzHmahxB/KDKpIinEO4dDWmvryAm
YnWfKcUIa3SI7JyWKw87/imzz7oXZ0p3Y86gmnXNzy8y9u3obZJ1Cp/C/HKPRmTyoXSZcOsIGmiP
rvNUxZegn9Plyvx1Atlni2D7MfGT2w0tNC8SJxIICNUYjQYgamYAagy5iH5RuUOC6mr4/I3OBUs/
g3QpIowK1UXMGumoJaQF4pbvXv/NrPKQG9oUCPpFmA/MagLhwT02SKx3HrLDoFeXGtK/ecaNjhmm
YTwF0fuxxOtFBqVX76rMXyZA+ZBQOR39wZnfBrc1EDjcgpcXooeoYd4uwdvm/6gnvqWe4qYtwTNR
VpCvG9hnNYBCTYsY0PN0UFrFX5RrInAc0Sk36lVM76JGYAvNmRHj/TtRiHVagA8CHvIKBUPEv4//
U7oG99wKf31lWfdtV/7xO0tCcy4uZzlCjwJWSk0vC6Rblr94Vg6CQ4+VgDT8Nu6vyg1JN60HjVTW
K+vKZKPED2RH1+QTBnFKOwfC9InDJJU1N5krXu0lywGaFfJqRx1JayuGeu7MwRBhgFrhxjjd5EB7
z2PUAvAsDDN2LpbwEqkDiH2hiTiLmfIcdaGr8KQe/nOylbvwxBILGv+mSWaNIws/3FepG2+XjDQu
rF7c/CC4bdMTiVLckzLr5ADQKexmFnvd4+ioVMQ3Z00q+1Fk4z7XSAPvBoO72TXAkK0K3KrPMDAm
L06piDP9o4EK8iljOHCxYZ0tGfnNGj5966tUPESvrYrUD60pp0aC+S9MfiA/74t50DkONLoFZBNl
ZxNwLaS7JZXzVyFdS6LBhpa3+Cazmf1OfTG9WEjKDPxT+cHoeKAH0VZuI3e44SN0Z9Orx4PGWXjS
71g8W4bxWTWRuHm21LHSWPPyimnoD4Q3khyfE0WR1zjicVzWwXQdeckhxXPaaaVDrex361AprRTp
PBdgBmnEniCxvr/QtD/Lyjl66wf7SuUqxtLg+7+k9Zkz+Xz5QCz9m7WPS4PKIKx1X36HBobkjxd1
som+fsNzjRdlokU2134y1DFJZdF8sL3ZoJHegN9aobC+8LSibQlBUpt+bquIt5nNOr2eaTF/sdLQ
nkE3bVcjk79R3iUSoNzcduUMZApqcdIAA/u+h+e4KXIQWZxrvMI8wHRY3Fy105YuBJ+1H1EZV/lb
O58xWuE8XYpGxcBQ2TG92Enpxdyb1VRlBTVtpfPU57DISe09KKKSWEkDzAP5FNfk1bzI21M2L8d+
/4H8rsR4Rui00nZ7E41xrmLSxa+rFYGUm3VbIfGaTUA/U5xguJafBE0Zmf2uo9q30c7dGZzVPe6G
FV235DpCl54r7RVycMJLeb0nBTZuL6bFauztyqrK7ERsf8UwmCy1KPkhJF1MPjm5OvaA23H6AXEI
jsc0u1PjkR3OK7fe9UhtkgownJAdyNuWUw4H3EMUUtje1Ir3ubDxDXL3VnNLt7YBa9THyxRfkJrs
LI9yaEL3FvpHw8V29Anug+gHqVQ1oIZd0pCuQaj9qEgZ+31F53DuyiiILZoEoEwdAcNnQ5N5FUOo
rvdyQ57/JsxXaERwKThNaadnwnz5YBfuAfTUoSIaH7CJVMr7x4Vw98CS9+y1lOC9iwq0DrJqCOTH
/K8OYXXUW11UKCLbczp3hw0WA4KzRwIOcV0w2adbV4dLJ2dcVkpWcVsApaXRkKOy74uH36sa9Sm6
hRTnayidwAmiOpDnZOSrj9zLSy5JAhW6lBkAg9+xcHR/YIYMSjIY9aRBv7DmZBoVrL/7WS/1LfVJ
twn/50pWVlooG1bbV50jqAkasTX9a19dsNMQLMn32C9dVRlEnwmmlaggc0m/DqAlPd9vcF7kbzxr
TTD+Et9QJgblFY6G4cscpxswmq/jifp62nP/C3Q0K1MImEQaBCLEpQ4pJnd2EeVg+rEdGBg3zTso
wj2oF/DdJAprzC7an5n3uGiQRHVVH4eU2VsjxuAsOidWgL4UqSrQ6P/Aa3XZw99xbjDmFzOe/HbE
HdFlG3/pi1sn4OH5lLiDYp6/OvGD8K7XKMkqLS+9+uzqN6m39UndNV4qNlk02VNWM5M8js2ekSzP
Yqbc4mg2OlTBD3ZRfwSZW3OQIyitfcZthOl/2qF3q1Sp9bJC+jbn8DxSJ847uC9c849DueS161Ed
yOFtVlkqfXOXFIPSLXOqXD8FCPvQ52Ltq6aiWG4nDNBCI3s12kP2MRtFyzRHHlolGoIp4qfrHggi
OjYE/2CU7rr47rLVDnuErZ8YWqq3DpI5Kix0OhvvoTfgQoJmxEv4hTvEUSptSRJoaB6LNaIOWxTi
sg/OS2m06ggN3Db/jLrnWmQ7yPtdaK8zq4qIl91yJavUZ8V3r0AyWUZtOUuvfMEYCmW4nGm6hxlg
N6rU5QjBFWMrnENBfc60ESqPJkNfVi0YHATPYmZusj3kiyDUEs7sJjVeQ7Zn3OyH088aO3m8K+Kv
ssZVBftgTiODgLitBsj+yhiPs/rYiH0VspycvH/lEYCKItLq3MG9+kH9HqXjJn0gG1k/7mbYA4h/
ahTA+EG4wFXgf3JfN65sBpGFiX81fnmyCE4Ml9na4yfSDkyLBz9EiqXZn2wE1L5HZmPnk51gNx/E
OINCbGOgqUwMoqsoR6lZn++YqYBWIM+jcNz4cZIjLfsRpNxu5k1yYV1rn+C1RyQOhtQ787e3e55K
Deb2qPB2eR70fT5uOfdWyufMPeS3NEMUKqeurhFeIvIQs1bOlRyCM+zqUyqcNbqDSEv73wP0x4ZC
f8E8iJtQzfwRg3gz5WivI1AQOvlk9VoAYHGFCJFk0F25QDtDCAAJRekcCQbgsfYbCSfW85GEo/2p
qHBX1a1Q4G7yzCctMUhx2eYZlkGz9iMXlq87JTktZ3r/x0ytzOkAK7k/iOPAoZ6tWsHBBZv1CmbY
J+DSMySIVKiDmLMxrEN1f5aEfqyIC+ORJExdgl7XHMzOBM04LFtA+L7H3bnncSXaPdLqZmIN2SE5
CxmpWzeRNTghf2LvMs8LTSxrprB9oErrRijwwZEHKXqU8VQGO3Ef4fslU+tTEO5hiT9Vb/YuPtnp
wpufhfNrDecwJ17dy7m+zYGHf1U8pVyHi9pz/UQbmnolTjO8qWTW55FZKkQwD10PN4XTlyPD7V7S
1wCM2D/Xp/fAjC2qmI8NvcUSQDq1GUD7jc/BL8DD+FOgc7HdQ10lDCO+WjNLbvlQqqmOoFPRzw9F
ql6YUamMyWRC2UzWH+aNo/Gcp72hJ+pQWAWE8htVJM3xGp4rxiAj1Xthr/LvMsBM/8oNOOCPuvN4
rDa/iUHYr9INgvSirJGYnhgrjl3WeF7i5f7DyXuK7fWDCjLioZkeezqXbcH3A0v0uP+34f7/24Nq
2YC6/UqfUIBqR/gB0kBkRmchQuoT/F3Wv/UeoV6BV0pSvOnp0aF15YUDS77wzdiJ6ZS1/ywf6M8z
NSQEToKX9P/siMvsowdbkrs9Nc4emBBVJl2Kt014pSTEm4joba1g8Qdi5+StD2PjOo5bXy1gcKA2
fLm7vMYDnbvkrBy5zL5qA4PfkP9Izau77lyp/q6dCJhzihywrx7r6fDOyBIFtUX+IiLTAi6nGkrh
Kkr1ACXbfddL5L9II/mXWNeoxBTXS4vqLh5bnI346vD07LPIqwfLpFgx/vIN+roEMD5qOQAqJKey
ALihFVU1NZHeNMIdGN0jS62i5b9DsQnpRT2lqS4lZkhsErBYMF+JHAbOb026Kb9J+qTTIn/1CyH0
VbrAUwO+n0OE3Ugg/2fOQln8qPpcV5b7j0+rWHb1DycP6gNuahLVjmAwmVxgp1Uj74ls0CXCfeMa
gQycdmGOYS7ZqDqZ8OclPgOMY24MHzNlQKcql1tBnv/aL6WQNMWd4Z2MJhgMb4UcC/GTtz24Hu4T
XqIRxSO2/hffIbQL0cSen/3Wn2Ly/lSD1cgmsvrbWusct+2GKQu+pqBWIMf6lLCc/ePHl9cwTmOO
12fwLDIC9onc6jZFyxXIW3Os0RkCJVxVej6GBhhJi5kj4ziA1Un35ghSZhl79G8MvqcM+qvr+SHS
ZLgG99buNEUJqee7r7e0lPpGPkYwo+tIoDjroOehpowGhQRyvJY09WYeMNVP5IQPdeoRcBwYdv/3
gpkjYuGGXda1VJLa8h/vkxEZ4xWbxB73wcX6QMYkDwIYnxckNUr2UosQN8H0FXo9w1NVSnDy260P
k6xRVypiL0ppbhSkidVqr7GGV/BGoGRRQMigvv8DuOuw3BG3/vpam4szCXZSI9cwQhsGbWIVfj9e
Ny/wW032d2XC93n7Jv/XJoCCretvtIdytlTKRuCzEDGMJm5Paqv9v/PPaYoGab3fr3W2gc/4QHSr
a/h7SKqnHfKuZXOGBxrsexteCm3f2rytMBxsOPe+EjCgzhoEXo3g59KmbS8pREcn4gf07IO/LTol
roB0i49xm6U5BUIbKuAA6b3myo77voHbVyERq1MAIqM6mn47gBCIrsvEvHAc/NpFsJ7vhk8554+Q
1oKtb3SyshWLEnT4EkT++Uf1dPjazJCbaURxHvLi+iYQoWT6z8VEVaVwsy4sSFeywBU29LAIgtyp
bkJIMCIvF2baylen9BSpKRZf1Sft8v5EkmeMUpdKjpsAoYi2Xt3LGkD7f9fAN1DbUru9FPX/HAm/
dF93QdPhPweNOCceTZ1zG+DeT62oykT6Vjv/9JfYd3Na26ToG3d1pwLejztLCSSwgdYoluAGRCHS
4spW6f1CiHPd+3f07xySswEdbTGeXmK7VgTU6iCQGX2UUxD5n87aHAbyu05WPG6rrimhmX6Aa9gH
JBQArJukwJdCV+8TWEdOI50LUTOMJMlE70JWjZeWVTksJZoHgyqWkdETptJM9bLxo9E4BsqAhYS5
dJ25OFbslQgEpMMDybLNRntTSwz166wl2DZAlJvWpMqpVxEcv0Z/KuBgqjWnnrqlRaRnjSS4h6ng
2DnLFAG0QQbrivLsTflfFoz7MBfi9U8Rae8pYIk6yYVfpIPxHgke8X2tWT3Px2J+5JpyrGgKRQRU
nnIou7fDOpVOux6a9zcsLXUSigCsUq6WzbLXsCDy4DikNsEfw7KaihOB1Z4terzXDYS3oIRqZG89
QiO6cjnOJ0Xic6ILgLdTQMkA65slAwK66rQ6PXXteXlX9M6sdOAKX+TsyGm6zVDx4yTXwrJkytfU
FmJESb4XALF20g4pu0/GBE9/W3MHrmGMlUZpMF49n2AAKmc3LzVyf2qm80z2z2wAc778xfuPpcv+
o8dp22Sh31dc2XFk/oiDv5pviCwb4bKcdIRkE6kab/2zkroG8K1q+vpjsuulBHoBG+yVmCNxPElX
2haVdZLSl1l933xmy/huiZFqeg/Qw+Wgwm15JaWBA8D04jqV4kfvYGWtizRTORILu575gIeXwpwI
f7ka4E7Q1bRGA5jqjY3AhUXge9yMLGJvffLQvSFB5e4Xq7Y5npOQbFZ0QM3RLwFn5Hemf7fWmV4V
3UsV6jsQISonftitQk3d+l8DwPbo/wxOzOC/X3xydecEojdMVfg4L48L+HPUoUZnP+1ejLDlGdF7
Am8fl4MuJYLnXQ+0gHoPcJA0RERVHDPPbWVKrSiZHvfOVsCig2IevG7kteOCiFV0axtDeF7J1JCV
eli5pCh8weeKEgNZj+xD3u/e9gtR3GxD2wYe6psO63hOYch7+e0+NN8a43nxBcUhN3Be6FqHcD7c
73GO6MDGQGAOfu1cX680QaIRrLMaLrc569sL68caZQiy4y9GUAQ7o9tDdgLnBPfaiGfV80QuFm6d
/IBCOzlY2O4LTcOJt1+8O6gx1IgvhCvRnR+IZEz/DxormywlOil43ZKXscQrT2Ce/3+QPJ9wgRgT
8uJqvDNSjwAtJLZjvcBJt1kFvi/D7tpwquGjL2mLM4t/k6IVfXzTAr5waZeX6PPM6JofUuccgaSC
cR5kKCi6RTsqO/ukkh/DNDntrmFbaKSxAWHU0wpZ7qY79CRrfSGNrIRmBk3yIqc1z2HqkeOXrUJn
0RHKSszgecAqk029WANql8/q/p8kPjDAXsV/KdM4hRSWqzlTneWLvLqbdEJPtbw8eoawG1OMUtff
44Yxp7gmuz3Agu/3J3BxSi28FTxolpIB6v68Wu3H3kkOiN1zv9PeT2bonjpSc0YlGTkeHaCuyaxx
oc3WVLFhaa+KJzg7lFK/MQqYM0BzSY9G9reWbCUJkUJuWZ288KdP7hkn+lpqklgN0Is5IhO8AK6G
KQGG3O4vz3iIB0Tji/Ra7ZxNuwNwdv+VetRKb5rUBWsP/s8FiuOLUFJM4MZ/QAWkpTmyfuu6ht0B
7Ex9o+tkNZlbn2KXv7MEFrVhOC778g+2A9A65I0T7rUan2qsT8yu4lC1tikwkFrvat2fYVdgrEnu
8YmCP42lXq6QeSqkDVieDR0SwgBrC7v8IuDLF7mryoku31/qQXe0QPIHv4g8shygc8mZii1Mw5sJ
bwFYYQkjpPZ1DhqAEAXTGe+t0cUAwX8sVgykdr+p9bxjjBWbMdv2HvPYnYPx6B1gw4Ld3eJtVte9
ofSEx4VMeplRboCSYGA/PSnozYEzwIEBZTilFVD0srBVg9GPMPYrcDmrb2fyvkDEHa9/276js6Zg
IxtatjdWvztgK0ySdEhnD36G+V25MhKW59hATDgKk7WTnk/dEVFKIFPLwRcl5jCLejGe9RFYcSrC
x0CfgxFh4Y99gtliD+2LZgbl+s5WQBMIdsTk/ErvMkfIPHKjCcVDng2i895g40d24iuvw+nvm5l/
OahUJMRX+kJLewK5ZWssjz84c9yFmdSLPYClidLlu7H3LliI/pOqnUaoNIotT7ROL9kwiFIzjsMm
WgAWbEpOnKOSXh8F6tF5Y/KaJeVQF88IGtk/75Ii9VgtKk8nRCNNHXnQqYaJPRvXVBvZ4onRHqf8
qH4lmqGxPYsvZtV4IdgyWwvG5x2CCn2aNNZJDKEW0Jw67T7olFrN2PdKiXb67k2IB0c0Vi5oCqqR
mg0IqZaf9gHoFrvZcK76xg/Vk8cwMDMbxGawOKAM11i0Nnkswimk2eS1crkbVjAZXldUd+Hgftcj
LUm1od4wVy0qL2mKN1BTjYoxE9swv3QKetCBfXJnVJtvDQ1lNeHSiRpJRWoYY1p/f0MBUO/YNG60
/PeO7upbU1fiuM8Ikrp4t/MByVdBD7BDdYNklcTJmpqge+KTFkYbA6R/w/4GRDckjtEnz98kXIV4
GnJqaTIDxumAAAe9OrA5WNfby7ySnwH3f1ljK+lqEvi7EGBmFS/ptaNXI8CmljYQsgSbkmT+xPal
vERBG1voqfkdzbnC82PTkjuGhQgm4adWgMj67XobqHZhBiIhz3lxnLyxe+QtqcF3vhyBmwhsTFwG
Dg/9uzA1G7iFEMR0etoBJKqTn07t+t92EfNyTLDIZh1CmbO41mCOFpSMLdWM3ANLt7QxE6Jag+/4
0B7MDMsl2YlQjS1DBYz4P8bjqm1QJdgorYeZgakklH18nDKlAC593ZSL91jOiQ2WDjC/nRnA1K2h
eZY6r5VwudgNpLkf0OJHSrQNZsWYFxcTQzKMn8enVFySfpX358gpHFMPtYujrpHFv2mP8m7nRY0q
k5IYeiDKZzB0E7nArDxEMFqqs3pQ4RlXoycDmZlvrZoxCmUNS+/9hgy7j6IYls9qlOlXxFZrsT2T
yocBC5Dlr1K23Bqen/cdU05p32HT5IZEPdrf2/7JwToEZHWtqAXdTBFPbjwoy5JTTMef2jygy7rL
zHxTjItGe1/F5hWSkpP1tXtyAriMbB4RaUGw4lhwIdhtfwfiHAeR8ESApLArjCij+uREUuXik6n/
Z7rHXmsq+NxN8WYjmPlnE5z1reuopMT/2lTd1NZs1+I8vItyOmhgChpumjqccNzAnUmxbc0XgACa
JdNhKFycL4cR1wwmscnqwvwLL0BzNU1Rff2Gz89QBLOs6zQWfM2KWk1ogF1e+IqACUj62AV9bJGX
eGgIUkyUDV3ljplULROPd6P3TGI1l//udromDrBFPFyZq7kqlTly8aLFgZETaHnF5ejgCSo/AX2O
s2OPGHEPeaPxPbkvkhxKNnCwxVHJzcxErk5tcKtDPvXTN8A8/y1oo+z96v3mbIIkNDQ8ZTlExq/4
sWULDf/6F6SSrk1rrYJGFm3JZ+W2v+Gf99ly9Cud0Ujz7gp5I7XwLoO66KglSbJ2f+OKim/Udxub
W0oLfOG3gAJECtWADCoHks5mW+piPCwow53ht29h+xFZwMlvlggWxz7lI1D/nSf8eWgK/1qZA4LH
rSOwHwzeQsy+LrvTIbzXASFYvj8lqijscYqAN57mMvgqQVLJNBbaNrp/zV+jGx6/ssCWNVSvxWRY
Mj5sT3SMGdGYbNVPXaTEbOdxAsu7HwpxNDZYoEP4lgNtRgJaf68AJwgWPWxK+8h+AEchMXwHVoYg
UZsIQhVePGxGiAbUzHV06E7tHBVr9k45zDKIdJzU0DT9I7VLU3WZu5e3HxQhy3zawfQHwuwJLVcc
1wkZdCzSkzLbVKtX4vOpCFnKVrZCKEMn4CfeJn7Oh3Aw1rMK3ehJz8pvWhF4IOtEyrJ1Uk/orvLu
5BiWOVDBB+fcYwa9j94sGAf8MIu48Qo3XWbx+hR6GX0A0tjlK15P8DiIxYU0vBM4PQxNfigwfZ1/
Q13INyMJxqbAl0Jf2XPWKuE9dnfqSR6VjAnuRmlgLKhkiJSbLKWzzbDlOBTpWjSBRJndhlIDTC1n
3EwuyDjCUG4i7ls/jQC4P8md3H+3b/rES+fkoQ7qRRmjqzalC7jPEeDYfm29UfaMlRqTDCRpFsLz
lXxnIwa2By48C6ypcFdsaFaSvRWgi24AwrZQZeXoGqpno601tP8du5JO14PLsvTKPUOrDM7lkv43
o/tKtgfUlvAFuZYiUC2oakKGp0CINdU8ytAEp6yeBGTtZBxbi3cKCSwcYrw7Gc7pNdC6DdIDp97i
BD6WyDQ5+acnlaocfaeLYBTI8IMw/bv6y4Yjd2Ho+0O/NthJYSFsBEB/wRBVHWatWddsR4nQ427Y
wnvj3fO2bLVLTauWzPZBa6awedQaVEHwS1mhXjLGAbC3AKucYcSus8B1KP9Ddb6LVQQmUTRCxh31
pUdz4ts5QmFaM45w8JHe131s1cvBycp3PnCIB+1YdEz2g9f7/DmfNxl3MBneh9Vh2vsq8OjweVVa
bsbLqX0TYelCA1RNXM6YYmr+f9XpUEI2RS/+YUZcDKpNFKhMObgEWsFkcK+ckYV+KPqVxzQdDDxA
K4D38va+dNB5EouFhMqAYbVx3yTA6B2i/6ByFsg0OOqaaJC96fvVYso6/aUGvYBbslkDM4Mh/tpP
LXvOh5+ZebLMAjYSSoM6t4dFU9br6MS6CZBxb/Ft84qWLQ1gO99bRuqvXpGXRzw/UTtf29PD6a9c
ekEAQt6gq42wSIkdphNMYcVHSIpd5okxliCyJ5BIlQkZCRV0l91Ai+crqZPcXiyglKgh3WobeADx
Iy0kEHEL8ct4HYRBJrZf9s3ujjCE0g7kRXy+tJ2xviM43znl18mpIfFs/COLJ8fh8KTbxLgShoI3
Y87OQy07uZZtSGlbyddKZf7ueFvJsfYRpNSFN042yUjF2oP4BAU1XnY4dZM3ScPvy/znPXYpOX+Y
UOv7MID5jQ0qUucVMT4HE7DxH7l+/hyViezjXnHd6qOgfkurw69KpaCRUZkkcfLho4m4U9cRaauK
swDfNfXn1xWCPAxw0un7zlJTL7MF5U7Hf9IpES1oYTsrCBZXZ8u5GLdbM9A142qQ1Vx75ZGc1CMa
MHyLZq4ALp6Dme4832QmHx4GSnK5NItNQQ/cZHWJ3UrYOn8Irza+icMVim2qzqqeVFLVUMG4NMum
+MGUH2pVb0UhIj51XdMHJKC/clUWWbeuZ9zF8w7EGkW+1ucyve6j7i4R2gUFXGfE2l0Tu2h62Klv
VckMSi8RLu61qDAdDvq89vPG6y0c3t9y+1Xr9YtmNiqSXK0VyzHvdS566Yha7OqjLuL3z1PuHutL
iqtW6U/wyh9enM1EmqxFecNNxwHErq7kTMqRMiAII3wp1cdSwpa4nTJVGDs+pzox02lAKfLnIKMs
CEF3CEg9xFyxRi1bRqrXrH4r/sooOO6BFF5F5ec1dBqZa46J4GzaQUaLitd2lWLg3SzXcwk/4DtH
hFrHhKxMsM8rDpdkyQum23om2/LKupe2GJHOXmMQK8aUSPwxCn61ahEZrwuTSWga+gkYH/GoSnxM
Vyo9OefxM1hAd2ocosfizABi7au/GqYrpYXYrXjxIQKHCBhNLzNWJP1tnANnPS25MYfZnVl72KzI
9c0b2InYSD39Wi/fZfnKlKGSr1v3Fk9JYn216hdTqtBtzL9Vp+px38Wmq9XTcXJ/PJXCrqpkLZ3e
uxmszeQGX9MmYxiHctMDwrHBIeV184lQXzHYA8aEO2LaiZNUP22EwKhfYpUKRAwgI8R2d7TzF42S
Tb4IEqG1e2XYSxJZZan9/jWoIZSgtG3kU1v9rm0fObddbHO9tgfp8A2FFHQCnFTVHqwUYAfC/FZ+
fO1FaPO4amNk0EeflylCinX00LvdIts31vtTZRwYh5ChdHFvhDCcMSavXCilqkQb5GVWDr2f3YDf
Fw/l4SLDS4qhcHqtSPqmA4w2dXFa8hsn39yEvlI0C/eHeDurX6RicE7Md0F/NRbcP9KS5lG0eHh1
OBS+Q7soxWEfM9DMjkQcsG9X5+KUbaJNDzUKGaiDaQGorR7xgb4YQD0dr5hgm9HwW76/n2qqo4kL
+09nTPKMH2RHfluMW0RzPpDHyE/Nj88ngycX9CDBlaO3I3iNFkDf68B/vrxc+t69MbcG7goIC8+N
pfijmvX9g1X5uUd0/0UJKyHIXRowFIobqa4uBzNYfzRMbfMe0u3FckdMwxyhUdp44XAx0oa5Na3W
ONVMPuMTOE/vd+eZKkts2K06K207+KIWQANRA2nzYBTpjSV+tuvEWtpHeGQEULCm6eZwirJd4a/X
5HcM/eqkFtr6nCrefFbnUwc3ns1fsr5GvnHVQoPgYboDQXQW3G28orNL8CfRZxB9RBpKge2Ey/Pf
DGXqbddGIxfSmOCnJftUdTOxCluMCiGo/qd8fR968uWQg3AHU2LwC1PUIhkxv17X2ByzHwSO1G3i
cTN1OznJ7Hwzru20WrbpnXvLufhcUNZ36xyraf2K3DbAyf/RErYLIrxtXxoBqXR5O+0izJaYPq07
HtH3eHFmCLe5eUWKtdQa40X8ULkEqvBVrJmh4EeS4H6y5efXWHvyq8EVahFtlP9WEXYQGT2O85fM
64mMULu6T+fsgfuOAKYzMnnWR9tDmr3Bg+fM2/iQxiqxti85YgD4M8Dkad5rbnU/pGYOcgZ6ihPA
26QEC2bMiwWIPtlNDNyp2lrVXvUSzlg7/M1x2Lj9XZL8F3vrySDSa3vSdkd1qRStiXztRrKWK0bN
qVLq79TPFui8+EgZJk08qf5pmIBc7WxC/SZ3P1R7fExW+vu8VvTg8VSiTq1PrUO9A6zfKo9DSIqi
V5JE8cKYoF0+E8efIAfggXgcRjJ19LRlc6ljrsNarTeF+6I0fG7D+2Ar7BuLwatRUfHPwrqN7axR
UYkIMaZikh4oks8H0kBxVEkGFgsJq+8DZPxy1/BPaB5OaTWdi3PXDDo+eYCDuXYg4rRYuzwd8asY
2ZoqmTlMn6+662/z5Z1BKmowZs/VQb01smEr6QBfWRXzZnAcJwmgZIc6EetvPUsnkmWgy92dY08k
D9/JkLF++kyc31vgdIYOpfbJhZezNZVNOIsu09OmXyB7ywlgbwQjyFxoQIXTAAQFcKWAcnuTQ9JQ
CKaE6nrcYG7JNVKMQqKV5iRKOUnygT/x9Gc7STcTYbVnnbtaSCaXH3h9SOexCJg0noPXwHHNsybN
r08xom7fKjeBqGlahxf0e9VBHYFa6fcXIHblnudg8y+RNpzo4b30p4uFRGhTvmC2ULwFu8dsWbZ1
WgZi6H1gIjQxGb0HD4znELN+17fP0mYoUQBZoIamoPRc56eZ1Ecm80OYnCbXHbIW/ohkmxYNKMkq
K2KoRFeBc0XJt+rTv6xdHyDQJ7SHjV0jEmhod9N60mFPp/lam0bXpTk0SA7WGGUZwof3AZ9esjkv
RQhyCGzMZEm669BQAJwC6tQ4Vz27IgrH71LwomtGlilkgXA+h+ffPmuVxkz6Jv5/rOBW/8mW8fob
usVHUckKfh3dNeB5rYXpCM71OARv2Zd7EW4Z7Rg44vIP5DIxwQ4wFBFVJhyM1E3B/QNSgjSteYhK
Goy94scW76WvycuD7L1rMJAvl2xALwIF0lyG+er6eAD1yLhJkRMzRNbySJwgG4HL1S5n99Aomcgk
01zbhh55MGwpK2iVGdErji0U5a6GP6hA+wB60xYsGklyM2LD6wDGw8BJQq39iNfo8waFCxoyddbo
wmnQSBR3pKVLtMewKcb1I7/4TEuKN/8V7YJyF+CTTSBsGy/+GHek4dpvKlMMFnLqJjye+pgFxXK6
bjaN5GDtGTFBTuaVmYlqSFoXmn5ET7sfCXifr6ibrM/zu6YU0wEOcNDfA42Sb9ohVaFCBjIIum+l
IyDniBoIrkdt0lOZImWNBZD//CYYR/8jODKPxDCyCjAznR6qitMyHLj7iByTvERnS8lBK9Ff/BoC
l7V/21x1on1RYFq+pByxO1vWCSqVhyGRPkO1AJt1jBFQ/iC+PpCoAfblQEG0iLIZicHzWDqP12QP
/RmVL+lEA9yyNEo9xegSC1RQDyiiLfmKHghcKcIEhj39G1fpEYZ7TDqcX/y0BzGkR8zZsmN457lV
gD8rrzj4Sd4Ds8+o9AY0UKFDIA/mF6vZlffjo5GTJkamDM+5quuGZ0kJDF8TfHvM8FDRrOg4Jc1d
Cjba/ncJt1ntmPYPEcJU8ms1+i8lkC6FL64T7FJtuxhivOBYklxK9d2Slj51P8NpuEfe0OrKJ0wx
V3/ym+v223QWRfK7dxPOQRAojusba+OX2peYzIXG2bYetXkaqsT33qOlHA7+5Ynr10ILzwyp5Dit
cWxBKoJH/p8NDwzQNNxuDTuuaWxPghIdK2kwSPC+PFj5R0CBzKuOmiFbGeeFXw90r0NCbeRIuwLR
4FyjQr1u5BZ/pDpgpqumbHuC08+yrM+oIaLo910DejNYPnUtY5THXRb5KwLbsUDtSQe6rfFscmf4
sEnfG6QmWHyOV7QwyqMBRm2VO9f/hjAJDhOT3Ho2P4BXOsTrVw8b4rkZ/lqk13s2Va8jjs8lka6w
BDuQxK6N0R9kk4dVMIAOAk9uTAiasG+Ln+JE12+o6r2HGIE4FLZ+6Mo9WiygdDwxXLyVth+Dk26B
WhTd2smTKbzSAdHwyeREOzqR4QwdVMRVWho4ArjdhX7TSOG2tYpDUhA51GkdZykhwp26hwFMJckY
UJmr8CTa7a8guoMKOXFLwuJKk4Np3rxQycj80IvTH1X61ZtsiLMDnQtWp+luvcSd+Oc1nnuPgX44
wU3hDDUjYpq3ONeasMTE8zHJhbzRkH8BoTA0cWOiWNY1xn4gBnTy8XyrewxrkSuS2sLcK45tR6W9
vwWsNpxbdAUjtua4l4qHGbzOHZ+/5YEEqVlJnvVqERzY7GjhT56V+QK/z3q5wU9y06vB1xZmtlQY
VFOHPobzrDFEedY0/C5Y/jDMaKa5Y0RIhB8hSkqHiwjr/9lWqQBASbErTQoMslzxQwIVfrivCNp2
GKqyOTiCphqwgfotA+NyGb6T7vCf36ogEhq0y/diabbt2nJlibIsvc1VO1V6ygCE5kWl8O6OwG2c
njrfwrkDFmW3Gy78/lJ7GCOgeIrmThDDd56q9pJyh8jNpv8/dnxIHCMaJDZZX5SiarQBAwr2TFQ2
gyqmJOwbOIn0imYiJrMpUQeJrtyPjQcpM4XScrQhTlyHIgexwTA+dR/+WU0W8JrTwvnHPA8jzzXA
WUhMCD49wpQ8KeUWcQ/l/e6Kj6yBiiUiqgPjO2qb/axQ3sMFGXCTCogLa0vII1MaQNsueKwXGu10
JfbqDpX11hfpx5dq2dlmsbzBTxR5hOwBfn0bFFL9ugY7jj+mPhOGGAUJzuR+qnmH4YMiGApqQ7vD
dnVPLyljqvmj7uIjWDEkd9eS0nkpR+poDGC9TwDG5sHREkZ2SiW9hmB0LkM/kxAnOJ8eFcnmncwW
gyGlBCMlS1bVl2qKe2LyVoPzZIIvz8lfKFy9tCWY2cC6qHYG2L6sfPaQ3SWXDlLsLG0JGC62Nmo+
f6IxJQ7GFvjeNBcqkzlSOgfXm1R3R2H5cNPTYOvfUrCE8SOaG2jOZMTpyMjy5JIv8KBFmTOsdWLp
9bQk+1zk8A7tTN7Q4KW9PU5YgumiTK56wt2o5Jlp7e3bSHU3SlNljFH4CXUW/Wa7v9IDVQakcPP5
CR5TgnXjofCxUpevo+wdOxQqLvKsGpkiqZGXbdcB4vmqyjCclE6DiQSTV3+vcyUm4rjUGiAZRj1N
uM4zbChPrYFFNtYcpHKii2H/SPBQLEz/EcjQZ0F0BMGN3HYOJ9wC2dN+W++T1lLgq9s3uSKyxzld
/DUCzvXrVrAH0LkK0ePl3WWD0jBVHgAYZQ3lgaKe1R1Te0hMMqd7T4/OaS2i0r2hb55E0Pn3BZ58
GfADSLcUseAzkNt/KnpnvcPUh77B8Irc8Pww/e/P0dM+YVvLdM2e+uAeTpXGepuiEDy+KgWx8vLX
DDSPQ76ajbbookdXRE3wQ+4boTkziNcdDPpaDAzmhMU2fzX8DoVGqnhO6JhEUXucV/q/5TZhl62t
1JPvyUt/1tq0vMPRNcojxH9DTPpc/Y4pdQng5jP6s45fW6H0N6Ib6Nnha3ylyS2S+D1EaYSzNzn6
18K9aYEJAaSpzo1AiIM4nKsyHYjFfO2xgQlC3cwtJUwrkdNcpiOFobB8+gbchl9WyoCCh5RfuvBH
52ABu9uusfRferaXzU/LkXSPAykjoePAwYniPfrl8rOmyBnLUBYGRdom20ZV6SojO+ztLsUErKuF
pBxicpvFrYin8FJ6Lpu5LFxtlOoshyv4S+aHyScwTnpPV/skpKeduvuIbbizem+Euxzt2a0+cep+
3370eCfy6rb7bSHJcUaS+Y1NuMy+TrIqSxera+4GQIA0WstjkQvNn91JwxjcdHYDqmrGGkHNtCsY
PLMaqRebgc05DNhuz9EwIxSJA0f8dbImblNSsFz9X+hCYJHjSi4ihln3EGW2Wpz27YkCFP0IA/BP
E+9TM4rAX6z8sGGzG6ETTwTT1PExGISJ2GRwntuIXhvgQRdGkdKdz/4jpa7Oxj2hOz4yzzYdlWwG
UWhJsSNXAEu/yykv/hxhfzK1H6B37y6YW+yhvuFBQYqCC9JFwAn5ixc1q68s4FvKg4sEQCBpNSWK
fJO4XGXGWQuCUtUgLXo+gqyBwR/8k4cufjSQ8rQzE/YCu/jLMyQT5g0f7JxeZAare/qt7GgI+h0c
Um6EJL+qvtQm3/SMvtVzLypkEWO0DXRpznSfH7rlsHRaT6PJSoAk3wSqN65wrCl9olCVY/3QdKiQ
0LoIX8KzxDnwimPmZBwFTyZrooQZw++WTECFsPlZDx4KrXvZAFJ/IOlBPNaY/8g75cSBWw9AJAyM
jhABV9JRu1vr9n5/1nxnk5GB4FtIuVH70zD2pVlO1iXgbcecRa8s9KGtXdiLCSLE0q9J8eJtUvUx
Yc7aIo2MSIDlW/LBXXLyG0fY6MZHzmqSdjn3zO1ZtNLmCf9vTeIh5yYl8SDB8iJ/oXL0ThhZ9hmb
RascGNagvQn0QEoPuXeYpl5josoLJH1gtuW5HxVB7ySnnCJlRhbGqbxIfJSc6qB6YVkIt45DpU6m
PVqjT35NkN54gCjQt6XjDgiZ7973to1Vlsjs+RlbeLvATuz8Cmao9XFHuHhBP3luwb/9ZMFxXhGK
sQi6+AUHu53dekK5X/1x/QZEIHD9ITFKqzHuwa8ELSGOyqWyiecsoDvrMerVqWiqGXohHdd8kOun
wKGQ2by4TP8hsBj9lszQfvjvao+zuwz6n2FM1kZWBnu5tUBapiIJ3MCjLVx4iT8tkvEKql28TKYu
ID57szoL00j6b9NopNtXDUlqXJ5ie3OTZzOBEIZKQ1fcpn7DecZlACZ3XhUJbtPXTW7NSB0DKdjy
Shu9ZyzpUryIQeHdiwhAU/lLmSPFEbYF/PDoBgsHzpjHL5m9ZWJhr5yGIl+MvRZj27uV8QllbSsB
yldKB2+QkCXBJ2VNMO5mGt+o/r3PQvNBZK8lbgi1Q0Yk8hSeNz7uutPvPS9kwfH8QqeRjRfJTyBE
s/NVNMBkdnBkIWsPYJYLmNG3hUraG5bqo9HHbUkF1OpslVqYiquMLPQCKYv3Q5pSA9/qa/OiJYhK
mL81twrNzE6BGh/5UQqeY3J1M+SmaKcu2aPMwKKPOhi1CrpTQeGrsuMyYosf4jCpk25HIsKx8EoG
f4pmFD6IvLWE/fPoxs0oR+s5CzIgRufiDiKR5ItuYIgllgcLoITYV8KkQ2lFt3naa5whcW/TqyJV
KMrKhQWJxTYmhOfo/RkifVZIqVGd21GvwH84mhOz7uBumEb7AobI7RV8Geu3JMnHc/Pj8cGNHLgG
m4f3FjoEQrUT1PMdJ5WvezHNtmD4NoFnN86LJb118IslyTZT+ThVTy1FkR/wh3XpRgV81zweI2eV
mUPC4/56yCtfxkR3JJAYsFXZj5ooWx9GH/P+Uw6l4bFpc0cckRc4guBchenX7aYnjqM6sWddLLWu
NI1OuUwRl4+ePhkflsLVupBcZNJXrA+dSWbQOsH/9/DqkZhHN+mPoirHj4Am4M2YgbyP6o8aeZ5K
MJXLsEZRujhgchefMinVrAl/4NpdCIbE9emyPG32TZm9WVz4Wmu2rweFYgCwz1DRKXvICQ5Cey4D
PD6zOyw36ZVc10RrOlwgzBt0pj3B9Ix+zoXWh8CQKWZiH8FvPv/uY/ZIzYa2URfM54QnattJOc2P
y+rWwihWyhMg6cudgouQgiepsfIbGNmJdYZ18uwD9XHajI64WcUV15UPcO2aiqtKAgJXJXNnoukg
oIC5doCrUv3e4fUVHLb7Ya0BH9Rpt1NwXT/itnDVqWOU3UfLCbDplgUqC0oLcqP6qFBoV8NVFUO8
9GlPloe3gsPe5BA9zNOmlFFsx3QOqbfjsMnlN5Alt6aMeIXx7O+0nup1jJQN8/yWu8OH4ibH+kBV
3xAS2U50hs8ZXrt2FrHkFjsCJQft+P85gCpENHnxnrjXmeTQmy+7cCQ8t+xv4oB31eEOmKBSMHKC
Ng+K3+HxnHUDMxmU3MkmiAe/9hi8MIF2zYXviyUPhybBJuMaK7SEVzdGfPcDnqd8Lee01GSgIvn2
hd/8fcPj7QN5FPo+fHiwjQe6H35MG50CNr5t0SI4o9Kms+JBctRQmdoNKJiR0ZTPTQEpsT9DInqr
wyWWH0kiEIcRfCZ3U2Ov1BYhS7u7CghSSnoUsbZ8sIoXbSgWhA5lqSMzoleFGWHPKgMK6I9+ecdF
sWkIcBtsbQTjZn0oXhWDUcZHSPv50E1KeoheKrhzQBAwE9Te7chAfLZJLap/l/KBQKnl79Fi6Yio
oLNEj+aGe8Vn/mx4N3+fVc9tJ1Lqna43k1qsNFAsLbSs5et1L1w0JVbx2jfL8OFyxhDfPbWT2Edh
zidTh9VoODmSrEY27v7bD2T+RbmCMWuBgguOK101OkSwQzH9nC746UUIS+pZyo/516+gJseZj4GM
XJ4vQte7QUbygika1pOXZo7XWH1y8HOxjr242E8ay6khXYQMsfd1yZVN4D3BV61TZ+fIVHWe6duw
hGZ70ord9wDYirBkMNVSslTshP+eepj2GDcTr/molaKo+dbWXRJw2Z/u5whOTCwmXszgoL1+szQL
jsobU4sIPvGCjyYseMkgDNLyoLj7zeuf5u5bnipnQ+9WViozBRbOMTuRhcTC4YRIWdE+dutRL+1Z
XHtnpLzm3RIs+w+0PFsbLYjgqzKeWrE+9nTcC/6/mkuvCQM+f8YQWyNagMu8P/C2FKf9uRrLkDuk
Xe/jQVD747xrdK328aXYwp4PKJwYI0YHpsfyyFsAt9lPoBTMVFxuXfnBoM7hfRS6b+838s+Hv3So
To5aMKE9UOAmyFDc/J7+g3VHIEDIuDA64cCIBbNhWugGgFnW80pWh5j5vyeLBVPgXeRiHi3dd0Ad
PVOeCkq+oCi3PDj80LUf8FHuRJR0yCttNe/M+QXn7UvHsnWGrJXP5tHttdsAAj5nnIm30LZdKNUX
9aSJpB9K7LRqCJLbTZSVK7ZcrB1PsOC1p5R84UGrDcOVhmHU4aEGXPQT9+RSw1MDRQHremifSA1r
m6pDQHtAgzCHOeJKzaS+CpV4zfmbc3yWIucdidJXw50IjOGXMByySSGArZkVcfrMQaZaEXapfVlT
N8S4tTkcpwll/qe28XOwbvJfuXn8SKHaxMLLH6t816q8hpwbrQTUWkLS/KSGJyuMLpw1L0qd2Z0w
aZgbRkhVf5TFXC/ix7Ez2urBBVr9eMSW2JP0Yd9F1YQ/qviaz6Y26FaBNz6WHPaP1t7rbD00wLW1
xoiQHUYJtpQsiD6qO4f7cLrYi/ltHnSJpDmffdfaJkk7lBb8RubIBPTOR3RxJx+yiGAM6ACtgvX7
7imYjgcIbNxatEL1fTtcC1bpDf8OQCfKlYDh5ARPU+aMgRRFKjOs4wA4Pzw1BiKu+9Suvri0U1c1
Drb24CZkUDkEb3tFOadX1B1a8lqp/cpriVR6J92BD1nrzSDsgO5z9KVn8UwiM5quoUqoTyDWrwdF
5hNguszPkMbbZvhZGPFc0ra2swddyCSwerSeVkaouHlaO3mmmDT1sBk/6Jf5//NLd2mnKH7QU9Vo
Gof47iCyYLLx6cpcf/NdGozSDqsZbwpfzAtucXNO6yrrwPUfYET3tWv9GtIxDQ/+UJ0lImWWluQZ
5Kbf8xIccTQMwj8cWSXw1U0erujbYZI2jp1F9vo/SVYXsv3N68wnSJMnCDUnOFPBn6HW5oAZ/edE
B1uDbjhH4cexsGwTKDYvTzD7Y2g9tJ+0ULAdip5lDueT0mTwqOJW4syurPq3oi9LF1brIYmU1HNI
Jy+MPgnMUIVTgVCnfH9d56tBse/s2FJ+MGiv/kiJtwK/Cg7PQ0jJ1CSTW7xEMLbv9iXw8R0Htv9k
QnPDI85C/dxwlXZbtYT3VRE7Yb01ndcSs6YjGZQB7hfVNdR5P6cPtSpGWEgSYppVhp/IJirPLOtN
A3rs/pgEx6oRojBcrC6EJdtFheSv+ghcBQsB20SPVZcOWM9Oqe/DvbWN3KyFXK7HhEb+MIC6EmX2
elOAGKMexQeOFWDIQq7OGNSBOj7Ik/t8JPt0ywrohtoXBff/cvJw3WAZMCqI8SSyGn6S17u+Bj8x
IZtn116eROQlrCJPe2ChfmpQZOOuuAdICT07A9a/EbIFmjSQy+jvGOfbhjSBqLapMeCdaRTg7bnk
dwPWLLLN/M4BcSrnE0W6Mfwsq24KLVtz95WxpKNMV9ScocDL39cEeFH+JB/sOYs9GtKdviPwNNiU
I/J9qQKGkvdBJUiOup7GaSuTYVZeiPBZLtEiXWcM2AmrFFDzwpWPJham67jzf+4RJXV7VL2wS75W
yklWyEJ81HAqaZPE5wHXZ5ewDI2DaCTNJJVBTmX0zFjis0FPhxGLpNAKRCHEXiTpDmjgKlds0ECH
AqChDIy4TfWQyIl7xg+/oES2j7j7SiXsrwwm9g2vAZrjWaSUlwuniwgb8x0faPK6P4s5ra7EB0RX
OVY5kqdkJKDYOtnm76nofatftIB09w6Hqvs56SJlCDJgFD8COYxnRQs8sjGJgDcUMzIxyPVDPpFD
gQscuY3JRJjqM7poWM2SaNCmq8gCEaN9mQUuWRtwSU01gFQZTLt6qCiaNEbu3xFUJoHIFVzu3JIb
C+yNoODCJE82YvZ2CFESujGPm9MyfoquJfk7u2HpRNYTmZNuBn9SIn+tWsVRhQacCgFvvY3J/USM
ZIJCMm02Qo06fJvqK/7t5hpxFx5FRNPEsEj7Q6ZBqI2Pekn6WuENDGGOwSORFPhgfXtzettIGfNn
BQaJFcvAVRL4KFj3CODgttJwEfrxkpTBMmuETkS+u5IiSeMrvcuw6+vtBZ3NTOGEEwSXz42OOjDl
eW27Xa1dZeopPYIOuSCFSf6XI2aETfMA7WUL8OqLtIWn7StuR1R54iJ2QxVTHTrCDzalcXQzC5Su
fm9jUbSsJHOGfmXpw4o9rUj3X5OhBFV/cPDwQDcCYJGz8r1dI3N+ka44NKnJJPUPJYKHV+lVk04F
L4oexZk14vY+ea8L2CuH1D+h/i2ipaMZQJUKlWHKaZjdfdeo88g0mBh0433YLQCncwb20hFlGkU8
cOcOfK2vYe9IEaUzvV3lNw19p8GB5GUyewMtxxPBVn7lBydVJ37NygVg8ixljwtGkz7jUGO+PC9C
tHgGOT/UBijyfKhU4sR2i+eHio8Eh1iY5wOcOfoc/O5JLIzN2cnCeRS1Eppboz6gBeBKnACEIZhV
svWa52knQmbjC6L0ZW7FtjkBUvcLzWGfdCUs/MGVuHS2FaBb+tRC7FuKa80aXt39jdHpE2NyE0qT
DJmyThjM5MtnhcxvNuS+UHd6o+GEezGNMor8vgzMA6isdurOxtauV8ekPa8xQOVJrAvYyqujDtKO
CNF7n4cmNrrVzQaG3Vw2r4iE1GdtO05CZTQLvlexAi8UUb1WU6jKNRTlS7+v0uahLiFsPztfsap7
TToI9AqflyOo0ULfba6y9+6S891+DsCFvPmU+uqWDBfmtf8VECjvnLG0v2uGDhOOqdWNDBNpri58
5t2gln3IHD0lh/VQ0jsuTaRQmK0hi2EH73qdCrQ21OCVFsMGQNjRPKL1WPdidhMHaNF5oQrSnoHt
YDgxJPXuXsilsVMT3gGisZ4k1NedmafOlr2RTAnrDWPIJWGxQAeHk5puHN2HofRzvaCWnPgYvMFL
fLaoBWp4WteEj4hl+9hi9w08Q6HM1IrgUbx+51pHIpocQrCQFZW/5A+RIL3bnuzxpJio2K5ywLNb
HGd6APAOBISio1xH4a14vH9EI0wvHmP1Fg2GO33rXmeamN4EyVy9jxJuLFu4diKSdv4MLLTIsski
es3F//zIRNJ1ND90c/FlzzazbH4neiJHPjCMPqkeRwJdo8qAgQ6X9aED+AYB5ZwUnKudBbfBunep
HQQ7mwys3Nub4P+GwkGAmrDFHWVSpja9QXVtXczpztxoaF8bZ/m7R00udenn/xAHAnWzIVhfvpLW
g7RqJ0P0M9EjAFY/03F9kNRqCRFxQgNEME43iouyspl1IWOByxGGQYqMZuM6Iu7qUh1pflL4a9Ei
Yxw7nuOSpaasuQG7ft0T9Q+wnpqmx4uKLZQQirQA0YaBNzgFu0U7wxvDEv9BuSDULD/O3yJCSG45
umc4+nmIvp1yJ2cZHNYMC9pJDO846/ZZSUeDQPdHr/9czwENQMjy1zBxKhc2G9krPbqcJG5g1VZ3
YeGDnGpZJuR1QokR5Jp3Gspql5zNu3YCfgerVNO+edl+3WUR3S/rbQtdv5SUUbxtyzffB/89yOTw
JJpZfV3yOEXE3hjE8nCKfUq0ctNe4RUn5zEcRRbqmx6Km3CTXQuaFAelfmwUrzs19nfEwSrBTF9R
ELJOxDjHhZ/6w/5YW+c2lKzUpigCsgaNlUKxZW944vcDDKV/CzTKhDUlDekAGXaUauMkoRMIaMIx
zBfZgrwlOfHVneNhPIfWJXXqLFORgQx5jsjx7FpJfxAvhilGhc4o8eWZzZQDVNq5JO6dL6pEXnu7
YwIZ3VN2JBV9Kvpar5Tn5Amtmy+kBU5TsFPuVDMN2O88H6c24t6boF+kFSd3Ke7SSk9M+ancoVG8
33cAweyjEqSot/FSfr68Kj4mJIMosPchsFkZUFHjkjcqBn3jOTV2HwLGH2jP5BQX86666PW3W/R+
uoDnJcTw/GZb6Sm4+GdzVOz4og/7yoGd5jzb5aaUcHSaLXXZU/r+8Mt3j7sHBRX3fNUKRHCgKpbj
W/M8a0YPYJQqmLB7qMj6SIaNj/iGTyQ4Ibw+mH+2B/TX9O0qSKCSm+Dz77luV4bZ97Ww8XV1Gwct
3q8wVFzLmNngVc0yTKSTt9ullgAQQAsMLCYL5bfeFnAvyiT+qTS3timJf/IlxWX9B/WGVN6eKfzE
bShyOPCAtng3Jh/5Eob8GybdBjIFcSkrCZ8yibrLVcHc7BjkTMsgi0Tw6+DfY6oP7J923kngEzWR
4h9qoAXpeqXjEPkFEjwFN4F1ab5HAbOhdGjtGrJ35CmDcmBxQ82H4Qmiz4GMs28l6Z9BGGaorJ5f
nD6Ho3jqFAye0Ahh3zmxhYxXRClUc/YPKExH4za5fADuvHN6BbxLnT9VP32BPKVmokhRVFJqFFV+
vY6D73JSPjUdTA/+EX5PN+BoZbUcze+wsV0hQGdRJnYns//5ZwpIm7KpE4yTgNY/u8rG2PGJA89C
YtoR/NRrvYX3g0ZmPSJHwqU5tVwqzbEh1mJySXAxrlLJpbkKqd+SJN8AAXYvssSTZWNAEN6DrPbV
S0Fc+8LRx3F6Iaf2NncYTXSN3M58un4CtpJGvoP4K87UQ0Y/k4hCKfaLCKpw9TFdlFV82paQeybd
JGanpS1U+HoAzcuC3ynn75uBmvc/hEQ/39phJ5YgfxF+2nSjjgH30LqDZVPhwCAUIgqHfV0nUulu
MTwDVs/SKs2UVYREATvoY6F18G/A2UfGK2QkAq/Pp+ik8p1UaWC7CEMDfa0bmA8H6k1nFHofiyKJ
Kinjtz9MMybTUC6B/3laEIMM+md6rYEP+znhr9cdu5nQA23bV+EK/1FjFJWjxp0QVRfDcR/1HG60
rUCXqZu9nef73zpR9N5fARro+3FSVRS5MdzJD4n+mA4+X8aH3fi9w4je0gJRvm2clhFgIbAJqoWE
Do3ZLQ0uuXkCOQQJkWnXImJ8n73++AuJU9rzhNGg3mm2loaXwc79pSP4/oX8UcvRoveeNcjhwdo4
Wet0Rw83D2GdtHbJBtLNIcqJEhpD/OSYQDPPUKfVZL9rNtWEmwCNv7v2zR4r7RgejyafclHrLv4M
v7oInt1VIaYeBdfeLfL2bNlEBP8M5QSKtx3Vg3fyvlredzqF58jU59iI6VJ/GxlVHrXg6w/I5YgP
0S4Qa1JycCbgsRieTc9/LTZ94XyccNEFlAeKHkOpDDh4DjyBMkAkEig1Epov9Gg5IEaZOjQ/H8EQ
82bkH8FOgpcF19VTiNEmK9kGVPMgxvJqTLS2i7mxYDajUoEi2pOV8dnYcVsQ4tZvvAA850H8YTZW
WHfBeNZn6929z//phx+cXbyUiWQ5MX5rU1twMIYRN/zGSovmi8m+lyCEtNqd4K8DZqgN45HqzIov
orpOv62Lgh7BbTQVGnl4hLYvU3b2riUyOYanmVwIrDn3NHbFxIpuJqVS+Uqgs9KK4CYLXQoWugbM
QhP9biEECqG4myZCA/VZ0EqrnpWpu82mE7kJH3rdUTz77WLsd4MDlxc+duab/I2ez4n8Mwe3AeWx
MdLLrgdgJvGaMv8WvZU+MgTHTPhHCgwYriYdiX/2mQoREb87W3AYSmw/6aiOVomJ/1vpnO379ZKG
NhtfAYAxJsQBYmd5p4vVQP1xoTtQmi9XOXvbyhhjiBDFXI81QL48aqNEH3jGzoHTSJOnTXHYm0hu
+ROkH2t/wGgl7qES0hiFZPiVDhyJWi/9j/UqiezvjCdH/YOnkms79VoJzRvNgv1gvoA=
`pragma protect end_protected
