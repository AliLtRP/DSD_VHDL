// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
MFKABGnyKoq/BKALpV/22bxQ1fHeTrMGmHsiZUPrPHprCStPyMKM+boe3yqF2IfSC3ZeMGJ06KKX
75DRsvKuePsp0r7aSUqJkKmcNFzYL2IUKc3ABF/RxfCPABk2C6mf/bp3IMak1brSZwgTi91FWnp+
driVGw/VCb6//WBhQu6+SNMXVSxUXWfdY8AbkOMhZUdG1f2Lpuo6OGJM0jpvfz+uW2JaF8+dNq3K
LQViw7PC3MISZlZ9piZs+nstpHWH+3CPY8ZbkGkwQPExUHy1wwbqlHb0NlpXMcYaJk31kSsULqjH
JV6Jr2WO6c8FjTPlxQbktMinZrubENOOhcVjHQ==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
Go9Sdw/QyyXiuVwmj6TsmIWyKyWqhXVpwgviwy2mEGGfM7i8hoTbyT0QFpWg7A+AbJXn7CFSgQ30
IHuJTrEdkTzMh7cvySCQEcSfGgRSqxTrA/zhKQglTOZEfzg/JyJkQILjbrp4lNXt/NT+guK3gsAp
gwzFx9+BpfCxfP/llJaWYu4R3Q9flx7ZvQR7/OSjBhaRuU/3We3SgDzoL0Gjrvpc8nQvxOBmDj19
rdeOX/ufhM+M7PiMKlPTGL1E7rT8S6O7eXVW3LTNwKWXei+zeWCFwtM7/gFMo88u6VklEYL2Ngyr
8rMfolo+1CPG+QuqN9KExdZcCKw1fYQkmo0iuzRfjfcQyq+Y6rGJKBm8akA/D/36umnLP93Ynu7y
fh1VZnUk7rjLv+rW3oXmErKnrdQLzqiFvUH2IwJMVJWu4BDLlhz0Nw0s+hsNCD/aN8eSKALl9ONZ
U02Nml+f6WU93xA9foYC16CFODcq+lbdzTO/k/0FgjEz3l/x/n00KnSK1NMwsMZ4FGaUK+XE690m
X2haX2JwnouyfzXhjsPu7OPedr6Ms5eMvCM6QWIuEnABrgHmNQPjQTldMtygMVo9ckrvOO0T9dE/
oFGc3ipBTfTiC4edsEVUGs/WT5C8SUnDihD37CvtF+PvBDGEW0kYbUXIXza2pT+bfzbSr0gHjykt
ojgFTq8AnOkAU0xu1b37OYThp1fzSOZrrUpOAMMKOd4eDWZfdu47dd2HsP9AV6Sy8LiTC2RZ8TDU
H7lfAKREgMo8RaIvuhVbb/iG+eeDCnKpvvWPpNPnw5eZF4eiFy/igk107JoRj2KJoZh1UQy3M+Mi
c5/c5Aof2f8AF0o1ioDnba+oh04xaZm9ApkEMXsown+nTxZy5nM3IziiaplihJXUMnj8Qdi+jGik
fyR6WfCY29o9o3lfCCktHEi0xiMIZit9Rb24Q2d8nfh/D1MQNgVgKO+uPYvoeiumc66iQsJypbDf
r9MWPmLeXM3jxLSGODtKlMHV8VSexzLK+M0gUVYil7FgAoWTV2UIrSLoYs/+ylcJLB41K6tykmUv
ZuNIRAnXzwDABdA0vw/sJpgQmy5O/fHQCB4nF4ajKHEgp8U93Wz6b4V9lKrnyFEX+CC71SkhYogl
zFNU8qf3JTQUfYC1p83/CSFBQVy+3OceJZnTdUvYpt5m1lvwsksjukC3L81VnP5RBcV+5Jr/AXs5
Hv1h1QbPPBMGd/tRRpbluApoMB+EUvMwmJea4kHj7G1ghkPC2QIKpXx0ly61q0ORawWStO6+U07k
iNz3lsFwdGsPFGprRJGcAoo6unLYDWVYetaKyT55PGET9OQ0qyTwoqkNUXAjmKLRHwOfbrkczb+l
R8BG1pZG7na/k0+P72hurrvOpS0AStreYcsTvT822FbdRJD5f0SOgtf7gnssF7OtML7BXXez7ldd
hRmI+j8n10Hz/c0tTUwBQEGbQuUIIIEF/2k4KHoRJOnykj5xvQRW+2lPsORfdR14eqzShuwZnTuz
E2wqrez9WAL+XHxRp4tb6ALmV8IMwBOoaCbVuIpfhqcQXwCREZHkYmgYQrSJ45TEo0f2PqrDoxfw
MjhY/zevBq7r2p5/QM2+5JLzl6V2YIOHqOI8xoDyAtU3s422FRi7XiJHD6myj+RxhBNvamvs+P+l
7xR3LloVCjXfqhnajhAX5nklP4LzW5iR0ULE4RQLFOX+oKQzWwZl35naQw3uhXC3uLWV+MaRipJf
I7lV2f9wG2Q3Gf3/iuVbDp1SDB2OSYoaAIKX9mUUEDyImsA0H4zs07i7HPF+CRo/0cYc8QYijJw5
PNPZE40t/tl5VfP2+1rlFMoTVAanh+G516wOUv3VxbkkhqZMJkaPviB6iZtGLvYqJDBiE1i90PMz
YvUmiPdogH8HosaG1IxLddfLStzNBa4AaRxCucQKZbCeYwBpH/T0wYlmmCbboRLhTlfO1T4Spv8p
bBuhpMa1XfOk7VxKYupXvS1MPWAX/sVmrewpcTI4eCKNqopeUPGGE+BZCLCuaJl33eB1FmjKTP3m
8IBIhFyK5CTW6x3EUwFcUXbEWEZ3AZ5ttD3/guEG6vO+eJTbZAPdcisuxLdLiiOAYq8IiOwcB5RX
eJYNJSAKaFsYqRrnSCOIj7T+O4GJ347WMeqL+lrHZgtxJv2l/qc1A4SjoklT9LgV2agwBdiiaRLv
vT7ngpw9YorDPrym9Zuau8N2XWzz0+5r+DwarYZUJlxPa+SrVNUFGbHB4KFO2hhrdeCLlmqr8+zB
H06OCs3rHKi1L+ozRUxCFxuEX4vo1P4827gufPNDyEaDdsjG+XU9ANvlFlaNQE1tclE+YVO47Wv6
j0jGJTUNqZT1E6lBTZnlwOzOzbTpKQckVJ8vB3Zeum9Cs3tZz5+5LJlI1sFDHJEs21+1Gp6HgR2x
NCajWw8l9WjzQwqnx4fAPyW5fW4ZsFdgFw7zp4GU6XnViasFmQFEJkBcoF0xGKm99X5BM8W+uSZ5
66olq9TcYc6nIjCwVUkSN6U5J75lyGDQHIomk7fjlrBWFDnOYM06lzHx26+luA7HCfNhoxBXQeXA
QxHtNBY5fhij4RqCyE4BgCelOLX9gOUJsYt2vPMybXXnJcKQne+3vE8hBIVQh3Wl5FyvBI2XA8V8
vcECHiVvtXkxZXVUnr80OLB1Px8QCGN+oxh3tpzBrtDwqBCX7qsFICSDMWAArnXS0TCoGAgmhyN5
S7kpwEpzbuKzLdp6eXrbrrsjokUo0ZJSgv7MS5OCwaqhh2NGRl8jVErKBiQ7JXXIh5RUQ/CpEAOF
BBepShy5OXRmAE7N3ch+/IwpDWcAo/vIXJGPnHleqQakBHYDtRUg+1lFPd6i2oFRX2sxNNMgfxwV
N4RbQW9tfgaIRFf58DGgFYQHpR6+U1Nbhj088RuJOC1IRFYng0XT5K9WdSifh3SCYAcDPVrisNCr
KuN8NEteA4JY4nRg+wsxnej0b2IWXZ5CRyuh0O69G6RW6FHzN2uOg0jkM1Q6HGdPhlu6x3MswFP/
RnCszUxPrOw6ZTwvOpI+xv8U6g8kn1+wdm55zg1QqeE90FS1U1GaExiUwxcIzg4fPGdf0EQYzDpX
5VRbcpiurd16m/M3xp4CaR7yNn3hkT3CjmePFHCc0e5gIvwAFYeMEj4AdmrqfUhSf/52r5vcVsF+
86BkEQhr0tuvGGcMEuUN3ZIAE1P54UoUq3Dm2qgd8R8h3z1Frlbu9EPRcy6RL1oZJHkXKRqdW6DD
DbnLK3omiM1OVbDYHnEtB2sMpvrOk9XzekXpevumXizRAFmhRCQeO3vZYoaWPHVu+GrR6zt/lt1X
ueyQgJoXEgCuc3FzWkSv1H0xeN/j1lCCDG/7HasdeLSz7r98hExxWHeL+Kayvt2uqtv12ps+1s2Y
3N31NnVdSu6nzzWjJ1mG8M1yCJsq+QZOX7+m8OqdHZlk7caLSD/Ocfxeo3XXzDKAQ59S4RTA3Zsn
8oRWSy3KSbScNvsbjaWCZ6kLR62EihenlmEw7o9Dy+ElPzymTkgaO1O+wr1vsc6nN7Be2KUhbfdk
B+uNPXQIqrcmdZ3IqLF9tNaXGGPaxL0ku1NarwjQhPj5F28DahXEzorz42E4DtJUSK6HxBwPyXhK
/LmaDYnrIcmrkBEAnD/X7GLsamQEENT2uKExHk4NIY+pcpbGY/jsOxTQbK7+HSEUi7wOVGQPpyND
hMVfBaKG7CJN7D3IuGYZR5fcI5pLwi22RaVY+ZzBO6A3e/MatiXpAutm+MpCuQ0J/AWmBt96CvlN
OM0lIz5qJOFyt4AY+jahYBffNMxhOGkjFgfWXsTM9e+rNEgbI3P6aCniWxSbOdcvqQ92XXQlIXzb
8nahfuANsgeStI0Nz+AlCuv9hHnVowFTFuFmfrEYjZJBDZ9ItJ7752uQ7DZlN/vwjKS9lwKaOdjt
7EMr239dzijIVV2b9ABfLpKGu0m06DZ4l/U7De2rQJxxTTpRGmA2FPVzOw0OP4Jb038IJEhDv1ZF
JoS0+dNIFZ+nbrKyZ8L9acjM2Ge/k61xnpXLdMY8Uq65so5R0WbEXndfG0xyuFm0JVFk+jMAfzBq
KSSg/y0hSLNN1AU1NztBN/adPSEJk7YkSz804PzklbEMflMs2ZnF99ZnOenAJ2rRwKQxKelmPKsz
K8eoP5u3rWFgxcJ5HVhwfxpgR6waH3CLuJrb31bbStAymtG3DjFa9TkJY2GGeEyNYZ0FRJmy4y8U
5r1xdwE93xDdAi5eER1qeqi5CCyLLbu+WVh2nJfTneCiPMfM5rNtWRwGZHR/zT3Ta2ukBy1v6t4N
hBmiESWwBkYMEkcxOkzBtW2tm3pgW8UwKgTLVtfaE+CB4vTB5xsfGOETXUxQdZTkNoQJLgR8J9lE
J++sd4m2PqvVXLyJsbMO7Em6fksr7EWn1doD6damhEF4AbgD9iyRKj/EXbudvCNVy+Kz9BZ9wI/C
PevFIiTwYpYbVN/koZ9dUhF4aGSexE+a4/uX8xk9AoFIZ9GffAtsQOzw/7CJZzyStiVa56O3q353
gEK0ZlhSnuM2vBvHZnXB6F63OyVywvEh9gBjgjROFmAMsZvePGKfYNPdtY+0LJhBZn3k8GFd8OdT
PoG4IWSepgAyiN5CBB5u3IRwPzWGWhjzDyzYq/UuM3JikrXZr0N0Pi1rHeUQscS2HSE2kSAqAMV8
0suwvzW4byzQHM2i5PIcbY8HCy6L+ntQ/Hp0n3oA1WEutyzz4M8Jh1Ceuuy54mjKn56KfachF4bC
+WlAk0B1AxP45Ov6FSCtVYQ1PEZDelLO6ad8OEgZP9p9UzCp+Uiv14O1rpRgdagmy9yZ3M+24yLr
gFyP3L7gwtED4JhAXhqKUbWIcB7SsY9t1x6AVgxoObiXPQQzcm0Q93FyZH77ZNYCbLmLj7Ios59x
SFujGRNvN9sS114F7BbxUsuZDxmsSjs0d5XASllcLCF7iWcPiZvsTr2SOr/OFeE3zxYtv5phak2r
a4wAP9R8ehHAg6ucZtVjpIVFSOAOsDtQXG4ehx2rGCQ8ajyAbsOXISdgHEL1gWXtLisjzZTo+r/f
WMHrwRNI+5r+Ku3hkxPEtOmpsUOwMXBPv/Z7NON8mUJ7dtJxCu6mn+BMWbaCkTYiPPheT5dWCW39
03NSXWeJ6mWugT6+a3Sv6USiOf0f9LyAm8n4CQeuefNUaXNJY3T0KjMMjxLQvuSosjzxGp1Lm+JG
3hOuPDvQvyosLeSayQFxe7SPHop7Oer2FyXiWiCDmVBO3yMzTA0lnaMptxGsrCjIdl/AfyeWHORJ
K0k0mCTfJ2lEEObTDMPhzcV6Hacy+TsWlkCkloaHJPKX1Ky45w1I3nRGvKJUuLMGcw5MFbGOx7L2
ktn0ynGREOCVcGz+zqUR3JuDcuc/G2nXJLL/uCjOP+/kDxc5hFEganoSB70lqmPkU9Jh3Qol76uU
gx3fbxeqmlS55wF8VpR+dqHbPT/cd/bpkv7/JRXbARxCEHG2bC+kd3GtUulyAMbJLLQLBoOmjR9Z
sKefzfPCKqMXHj3bHaDLuMChwc9Jf2UxTkWj1HMnCwx+euG6H19sbERU9aiCKYopcQ7XV2eR9p3O
oZXTW4iUNmvt1bStn8nlm+baEV/Qf4bqCW+u+27t+x2BUyC9QqySPdcoSPYO8m04I9ADEwAU52WZ
sx53EsmuH4WBChfWnG/DqZjiKDovB99MYe0x0mf3H05PB+lmEb4PFlhQ6rKH2v8KbPAeo44Anm8M
2n+v+iTN58sYA4RBEJxVxRRZN5TMH5EpMPAGkPYAOYzj2ShDFP5mEncN7lUpCvtVhwbOL0rHJB/C
LE0u8R1GPhNuesz5MtMrLWafidDRmJAL9bSffTJsf61btH+eHGX366dDf9i4ZF8CvtlRZDSK7pYr
GX2GjCJ6x7CG60IoL/zfyYqMRZGsJSW+7t6IRkV1cZESoFSqtAFz23OMLyzYbS0WbCm8zKlG8dK7
Ip5F/SBj2+SkAUVaxlkrPzKQbi0C7l42+P7d9XWKVSmjIsTKqzkcQP6XjH/YQyLGeXcweZ2E8rCV
/xaS/LvA47ztWpWFoWB0QEIvKUEim2KhSN1FBY3+TUyZ75iVxZAFfWjFnVMpCBc4sSTGFngCPG8T
p2CfFZr90zcqMd+1QXLfHYHX2mOwXJZT+7C0VRZUXs82Vow6OjWlywK2SJ5atXgUJKvJulKtQPqI
mDPz+BsGpqj0rccif2KGa33QoczAaJv6EyivHgPpwvb71wGryJ+M+RPaMEKzJZS1kCW4ISef1LnO
Ve/M8+fg2WBhW+Psg4fLrP955DHZKi0DtK3NrlZNPk1jcQlppymwsl+Z7QqQz2Id/89G5T2UQ+Jv
JSuoMs6tbs8H6VDpT3b2/RBapu4lRJSJt9e4wc3EstTWPwVF/zsoKDRy3DhozWpuV/5fS0Svzf8z
EEVcDmTy62Nu+RWMrgz3RmHkXaePQcuzD5PF0GNKyDjL/RQdj972gWjo3A824RhzRpqpGzqv9zNY
Xs5I/sp+M56YRF+cCFYNZgr8X5Eapi4C6/sLSxa/8KCrD8MerxEE8vlvmuiGQD/usQykjqdjI1yF
dSauAwy+WDSHllY8krk4MBAxUPXPDPbnYN90+83OLh82lp8ov+NrYS1QFlcnC9gffQZja5lu+aHl
4DXtYcNJnxdFjx2a+3WxIEvO4Kwm0S9ng24uOTzxoeyDJBH1jQImiTP2ADlb6k0ahEcSAXkZNBZo
QcfGQ39Cgqxb5zHu/Tw4FqqOYmbCfME1noq9hsftGsOjXhHCWBa9zpbAYfoVPCL+2C4swyGUsdiI
diKf164RNRnqni1o6BRIU3f2FHDO9ILyOY+HEHeLX75YkGfE3ykcRaixK3ZxM3qEK+iaoRbsjxSi
LJ66vIOAanPa4LkRYdm4endzJ9cG9DiuHK+Ce80RDifFC/WFFWLyhOLo6tGgVX940hofoGu3/HU1
bB4TXjm5dMWn0XIR3V3kcVGUmJeU6bk7AGRYoRa0uwZgFfMTWwKWuITg2JbNEzEu0FKFutevapj3
dyS3+tvCqzTwOoG+68yOMoSgbHrkeFfH8kqLuEPzGtbKBvKLzKJv0tgDm7ts1Rf+TaiZfuslmdZs
99st3ser+gGuyTWH2Kbn+L7pBXX/F7A8nJ0Z2LzCj8dDshwotF6mFq84S+DRLZwn/vvFzk2rt+m9
948jaUBifKefvUQSZzLAHR7Slt/500VNpEFFN/bu7CXarl4U6kCE1y1IiyMq+t5/ctISKa7GjWUv
vGuunKjq2++/FDAeS2G/FxMUfSxw8U29WTlGPxFyoMyEXr9ZQb1GLlBC2rmrjNSzCbwD3UliWA/p
OllF+fLzc5HmTFNVftTfCGSPyD4Sz9NVgkVCf0HCkPcVPvTXAIpjpVJCom4Ev4TT+e+DsEEHKTw3
RwoBYZdiwrgeXvsy4Pl5+oL04WDaaHv+Q1xTLY/0CYuWdjx7Vp8BAPyMhqIEGhExg2KB8XBjrbq8
XfzSo9fefPD+vauPwf0YPQKOpw/3s6FXNLLGdKsSYdH5/0z/2MqiXIOGxULzuf2Ea65U5TrPK5Z9
1KaDdoi91TKizPcSoE/x9VdahDbVccP+/YYBUPjJP4g4UGtXycQIbNtpjd3OEUM0/bq80ctA6AfA
ltcmGUhQOFUr3p5fBeEOsIV2KY4BSHkpszmKAhGhh7UlMANswR52WHCLajr1srJVK5t5ylsZ0Lin
ZgrnfN5ubkRf1lToXAtSSQTrsDMtpwslONgvE0AkGWf9Iz0ntWuVFib609n54umsXwYdevFXiI0K
HOWy6S7QLpL3F0h7sR6WkROWGgWkl8siRL51bvHTl39cFXU3AsbVzuXoUCywWMamtW/XC+WHmBQb
j+O+F9WGryvCuPe+yQzgEsa8gDz6TViPzWI8YSriY41lVsPS7TOVHtD8kOnczLzDFCuuQsZ4b9Ls
MuopgKhn4EGn3dBlxeJhwHNIjiAZrqT5/MK2G0QLZscnZXS1rrwDWLLsdEggT30vSrd+4JmwS6b1
ZcolmFN8wZkBsxi/q23Npftms2m/eCxVdiCu1IfFWLh+GJG9OysNFdcJ8w2/6cY8pkCdETBeK8n2
LU/gluUApIRIqFQmNawMjsamX2dVDzgc49rSRkQ5UTXrzuvFcWlvTkF5CXG8PYP0E34P3OUI5M25
Iq2EWsuy8ztJcRhzveeoAk1H2KdbSoE2Evf5bEKwYjgtaq6llb2HvW77c+pIj4pcwfJBJEsSFFRH
Y6bzZPCT1j0kh9PgeO4ewwM1RrrTJ/4gbOyh4IcdYQIpoCfZdjj/2VAhzntswBiEpFmWUHXZVYkw
LyN5jXbe1A/jA0C2M2fiWtkikU96xpZvt3//p0wu7PLsF1mNDHzrzRxmvHhAvEDRChYfp7fxiADP
3kDZyP7NHD5R17Nun4Jo88N2/Y/FR72f3VvTLqm7JJHAz9nZuDS/ZB9Y8gYiO8susfkQWMgZcK1f
jw3kDr1HKNCdvcklEjKyRnLv3Q0kG23+Wn99dgJ4Q674himuek/QvPtysFViFckLPrdkIEwg/uAT
qTGpbOHZG3vHUJms/04HNP6Xkhb6b3MpwHWyKe8UU63Dv4/MD6z90/u4o/xCVkReAlFWn30CHOva
RlpXuoEUM/376ql9olwh3P/KTiR+wU023HfBlz8gR0E+njx8Divwh0o56NDRSgAdhtKNhPw9MLfK
3zCczrVKtz7MPaFE2N/aeS83y1wI6CYa1akf0aCIalwBAWqvpIGAoNZ3E2IRvZUlKtJ2j0bX6Atq
/hsk8by8g3Fay7jtfCuV+PLrnuAF5x/DX8MIXbSkzZ47yxiewuhbrwB9yaK5MhlJ8zwYw0OqFBr3
sf+TpmCb4z+Rvk8h4dw6GWBH4Qpi12HA+gRq8E1iAQxnUP+QjHg1C3gAu+8xryjjFZBgj600G2sR
4CtgA2l6oIyUnDWUexHzzrm+qMOfIx/9s7iJa0h4/3zHlrwvmB9Ep3dLl1Rz2vZoRec1iRZXFjZQ
zvIS1E1Zkd3es9i0r1Pc80Wa2Ti+f40tWp6gHHgDu1tgq55nV1hsW2M6p8Wrl81fnU4nF1Gfd0q7
/qL6OxZ8U6om3tWCVXuPlfE+VvLirJ9dKZFzD80WvPJVahZhJUtycNtpsMFyDJIPiRN7JgM21FcY
7gYOhx/vj0PvzL2B0II9nPUfjrpdWSKFC9r/VLu++AaslHysP4ycSBFHwGK9Kg3+DnuV1dmmGgvY
07+K1reRwnicj1cB6k+DuZCbUFj+dzkJg7zfbLLjzhZFaczAN7KKqkSW98HEzQn5b7oBHRxNJ1S3
jgLiICAQ/u2g8eIxUnNQ5T9zEnQhu3j1j8luCWhwRgBdRd5NOXFZ0kPcYBc34fZtgKdGCtnPeBuk
+1uOyJU2XQchII6fIZNHkzwcGPbLQUuSTXHKkCqBDtjIGkpB2rbRHpmAgkDqDDnw+/0708qI60Ov
+t4vLTgEdhaTkOprLu+tKhwQ9gibja+NmgBUe6M58ME/Cstwq5DbIRvFdeYJggeQPbPjYRcG0C8R
rJX9W99xvPGvZ+aFZfxrHArvbt0Z7HGZng07RXdMpTc4YyCcNrpNlAylCg2DIPv0COoDqsw/GtXr
Vrg8oPQO4wh6Q2fjG/harwSUGC37IcM5yDVu39CydZMaE4p4gyv8dVNKGXYP/Kzu/T6Adshgt75M
0MKSQ2aQIJe5XeIX4s3+NVQZ6OQARWtu6aIeJHsFaOyT+n31XFqyJ6X5sHvhbatW6hjqGtFWPTP9
U0FPnT5YAkVyRmT5ubi/sggiFzGbzWLpYbMQOJFeJ7WFek8lqDC3n62nVjIJ1NcgLLEl6t7VPeva
GWYk5/bVd17pdAOYTPBpDdQGl3rLRAEH1yrBwC6TB+AMSG2oqPtEscWVJlJKKh1F/0RzR3X46yrr
hZDRNm1UYzBy5+PsrCtmidaWAIxiwo86SzfoD0RrUh9EIhqg2VgQWIL2OhVMA2BlSte8n95LTz2R
FMMyq4IYXvsRzC6GXcoNiRHKumGWMMrQ8bkpwIYzaDH60C3k1JAsbwNgM4rHlld1TYE2v4E6q+0m
9sdGkwmlChvLq+m3TdSmlj2QRTmhHhuSbIkkJ+ZhXbdsI3e0YriyuJx58btwmTtmSiHmdMirmxcd
M22C2BpHRpXGi0FPydhZW5cX61iPf0DP3+kArXDl/WlWIbWg/N/POW4JvIkSctZXksxEDzoL7vLc
TmfzlkSh5U8v5f2SLVT5DJSyjHposh0wP8RvH7JNAr9nbPE5Yg6TW9fR+mL8O20sXw4/hIN4f32M
Uo9FTBPs9K7CckXu9Jo5w25QDpu3X50H9ksfMufSLyM8NIGu0UIEaGKjcQMeZAP9pQpBB4t7p707
XT8Ifty4LIhMYLJNlyX5P1LGkPTlQNvVsstVk2rN9jRwXKImT4bRr16/eWyt8GpqD68HD8Yp25nN
ORpjxEBekNNgJfXbf3rpuZ3rNyLsAqxS7G7KWIovG7LPqRDJmbkXu4KSBAIVBpcZisLY+B+8xUUs
87fjQERBxNKwaM9RxecYDviQmlVqU34F0IOtYQg89GqWKCO4rZ5Z6oxOBdJS5rUOvK404tphxWKA
uzS3m9F6583sJ2aUMjsS07T+GL88hBVkI5HR2Wr6R0bu4WMclzhP76HQ1qOAqi6BUAXRD7+inssN
Cvui3t4g5838DxEtm3pcQLK+kPV3wMzcLRZNs96YdjjUqaV60FD4zNgqGh24Q+CWgd4rF+yG2rnp
90KRCf8Eb1LspVK3yngmDPvQU9Tab/K7Up4FhN8RXS9cwNDuLcF38eYQZsNOmqI3Q7rofMOPbYfR
kD4+Ld66MsBxUkg3RojOHQ2lTr3PGdoT3iM0KvW4bI66kDlf1lml/dwSzOaXvS08ncP6ZvpnFM5s
5lrwZcwzfmJaGavEIl0ABt+dkUoqZj8gaMN4dC3o2LxxtCOw3HPcCBYkN4Yu7cEi58AmX9m0lwgO
xG0Atqbpbxcc0Zue+olTrDhSQMV3HekfahfVd3FyGPFaWSs1jFrYIJZrYkGtjJp9zZuZroKW1g==
`pragma protect end_protected
