// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:35:51 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
fsctRfjZOb154xvmbdLEvP0n4Un2L/e6tOCZUeIAM3Y9pTs61Mcg7FUlhzgQpftj
iJWAShXwI/H95+KSW82ruCvEzi8/Jo0TlbX7NX8VcI9sFAsTwaGpzVcpvWe/25aq
GQj+c/McCmTOqZ7HPFyYVJgRFxCryHeQDgi+nvucBts=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 3712)
dLwIDwKRwYk50ZqM+bbhW7+hBcJl9CI9udz2pqn/DxZ6Ha5RdtipqVg2JvH0qQ8w
HWlCoGIvjym+X9ZdGApDnUBE78S94xs4gw2YAjnWtssVT4EZlnI/+Y83Tkij5xEH
xH+CMYISiJ039+4YVZwpw0xLxWQPPFhDybK00AIeQIaJrIGhDArJj5vHNGr5UJbs
vp0F8l81/KbHfwRP9/kPSBlVptZMx+9IOFcAp9W5lapsOW+SH/rL2LXn/gdZtSxu
BzKFcLU52EYFAi83/qtEo1J/B5ayWOAxCLZ0pzC1giff2riV7rvIbE1W1gzkjguD
Sjo0IGnlSE+41f3aUHiFQlrkfDbNtTicHsNRDs1+MzrSY/mJ/6PmqOv25yISThga
rWUZb2KzWVJjSslxjpqaiNF7WbJvA+KWOzQKaguL7Dxii5Gm1gIZiJskEOjIKxUv
4GP8hRUKP1JKkS8SclCpoY81SnMCnOE5AMrHXcxf3evDCBw7x2mFz0bEhYzyzFXj
iY3o5hymqOaAZ32ZijbyX5Nqn5I6kbBlPv0PrnkbDWhRFrMqCD4LdBRKS8NIkhXt
4387XkPTul/6AcwIPdBlCg/i1e+2GoEmMvqCxBW58x2uEsAy14eY92hRz3thh59D
0iFByPnTGuSqnUTJPvtgu6BPLxbvUb3ZLV+w08nYZK9PF1WU7mezxNfAYtME+RxB
dQRsObafSLtC3Pl+biprv7zoqozUn7qzpJnnUsbRBQsLefNL6Qs64xlcANURY5kB
at+OnMCqnqrPgcfU3/EkluYEnoqXEF56fMaQEKHyPasPtzdlcrzIir/FODb8y7ks
reetFRme0n3gLywWBo8R1qo8qXZAbr2iO4S5OPyIlIlCvVBXbsxCqR5eBoA0bhLh
vY9JAnicV+m2wFfHLDL7b/D313zEysWUl6Nl2+fHjL/JDPGNQyCzYdNeQcvAswZ9
ef6KK7EfCdURqoY7Bm8pHAcze/O9t+B6fFcU60Ey5x1Xf+2ckouDfRuAW4YpQI9S
i+uxZzN3PRJN29g39Z6vDmq4Gpandro1B+HhtzGrvGvD0GK1S9JKGVwjg9yUY5D6
H65w+JeBKrHht7ao5ekEJeWx8MTLCA9vXRnsFmTHNEPbicRlRiLZSO1VLNKHkFr/
PcRqh/KRzunt5URoYMXg512pZu6h8VkSpOuJU5xm5zHB/gCF2VGVaqxAH06qJXjV
4VVQgMStMHuXR2/r7RBLmYSRjSn9raZ81qWScfmd7BVB8HXEKCMMhuBWi+CgvpYC
ENiSo9QD7/AFZRwz9YvpevkOe4GnR7qWYGw+4dt0ewEqyP9bJk/5/CTLN7IYSp4m
fI6h+LhwkS3Bt/0Qq83q9dEY/frlaZHxFjub8d5K7aCkBCoz0oMS/dfxrNy8UDp0
oN4+OCE89ZlfXa5+A6DYFvqpCHNVDeIZRWSFkI7Si26kycbJo2Tn9RXbEtTt9mTK
Sr9A2taHwvc4+clcPj3WUKal+y9+prQfQS/jpZ4GYu1wqQxVjE4aTWfeyhPKZZAZ
+YNL4WKx8DJAyhklllvEN4emIUWe84qgJhbTIBsnRYZrAFK/J+FpaerJ481L68xm
WFmQnD1ZD2F0tk82HavV7SX20gjCURlpvDs6JwkiwO4m+0EXsa3tHSelgXuFp6ZJ
Ws9jOYW7xzF1QK6U4riDuswzlojbnqw+CSqpkv60zV54QwJ8b6mCbLS80n0OsZ08
pXyyUdPWW3xCFelRB3tucDMDbBrDvb/RUVLEb1kSsJ5K7SBvA6K9h+tFvpMHwGq1
u20GwQTgl+o1RuxqDqj4hpOENpA0DkhPbyTNumG1XPj22NNfOe3pbsct9BsKTVtS
fkeUTY84mjmRIlylyXiH/LxK0k5oJjJqd5GsGZvATMPODaceaUbYRimxITNJkqHW
MBaFBuTzKoH5qeZ3DWgUzmrZaE7XaveknrcZGg34mKO8zItOKUyNFVpjYdnU22sb
wSEdqPohsAjpDQsAkuriguCiLW+yW+AyXUX9/QVDpjEReTDxtGDadQ2gpz8V5jpd
8fkwvFzMcp8ibDLeWQuS3rzYgn6Ly1EpiBtaBshCyZjkqJX+h+rSMoIgcD3ZDdwV
jK66xDCv0A1iOR8qimSZ5s2eWdGxhlQwPMCNcaL0DJPK6/MkHXZ8vm8hBn6Vfu1B
ptUTuvC3iealh5vMhwJ4rAIKg4vcPzya+x7ZcT7pE39DACBG2eK195jsLTJFBpMj
vuMj0wp98giNlafiqbHCkl2/rdibimzGB4HZMrSTHVbVgNO75R/7Ilu8/uxCMKUB
ASZO7RNo2E2yYfPuDe7ipSmyc90YOsYRwqf+4cvfHrqPqIVgyTG9cGN3ZsbJqPFJ
6B5buHh/Tgte057mPDvE70HwZk55uyA1IH/g8l3KWis/ieDaIASo4gJVwfAK9DHC
2F9Lr5q18DLS5j5VuoPWa0HfBnS3T2uSK1vf8TN0l8RbnMVmXwtq9z4AUgFHgGDT
WaNWhPnd/7z+sbsZ+ufw5fjXm/drSHaSpTagzdxfdZIDDexRB78fm8p6xxjbg9Hx
jg5pVa9pVviZy3PYoNh8x8g29uW6/3g/Bh85vAaL9uEFJZXiYx7Baqpx9HZDsuZE
HEd4UQs4TWnmzpYpFe2H1MczeFoX1IsWw+fbsEFg24aewUwGMMGS9RBEBNdnSsOX
qcn2IQe3s9BrDfRoQoGC7KVdb4m7lcrDniiQ0oGWbbU3GmERTn8SZpX4/NB31GyG
6j399h7XLbz1/wMCAgva3PiMzR5zH7XhD7MNZuN4/bdkq6DAVhg+f5VU/fv6tzO5
YIkZo2J+B8isYhrL6yD9zcHCPDX99XEkzVcNPRm3wUN/A7PSm2Hqzk3AGf7k58mC
wjccfHWw0fMRCo2uwMEU7hLGczECysv6/yTGa99Vn1DKlNfqUvvDNG2KU+ktC/b3
NuTWkofuWRApets1BQSwqt8dTL9uOeE7NcZolsfNNjt259EG7spR6aA3mlcAmgz8
tzUyWJjDDW0qugM2cAlrNLTac5soJ8iPiYovAYezf5oTlLjQQw8fJtEQIW0Dniyh
kZqTBm8k49+BP643zNcAuO06o11QIisFa2i3LfaYZOBE56/IvZA811AWcNiH2c/j
EtU7KNnkmL9xaTb/VOqVosqho+1UTMA8vkeI73/nzCbcG0qRaKEuKVSy1EbQn3Vc
YErhmVnQsa+ChUArYSX4FnbgERWO/d5kCFnehU8TAv7La4S42SS2wRGdM3tpemN7
GtZg4KisonHmSkFIg3jj+duWjzZU31qN039r3jqF6W6FxxbqNB0M5WfYRXoBLZHE
Zo4CBYPbGwnsyGx1a/KPvpjR6LrlABOv4tVPkgBUzJqKXjqleLJ9yrs8mh4ULkyq
TuPWinKDyg8yzHRitrXCGQsFiVk/l/C98s4EYRIs+UcuERBChKD7j2R2uNWiFRfQ
MH5/M7nHQoHAeQivOh2OnubSfO7NdVcZbBMUI34ji3JsumYd7gbT9DX5I+mcArzK
CiehLz9gOZih7MLTTKPBM2DkgA21qmPtfbcFlFldzf5ICkcNwZ7h/WWZyebXkA2X
p4H4hiG1bD2OFIerLWHzJY2lxMSi+7hrwUagEuK25ZjmkTwAhve6mN5BcHRwqAAN
TbHMgY3MEUrsNEjswumkPTu5/17FqrXuksYcuYuCHmrPNPzNij3fsNVJ/WMVclMd
DswybVPgq14bt++xWb3E4xND79cN2E4FDFxpG65GAwBsp99dtND+0jfEvWmIPpia
eJnqD8EAJ4dC5cj7fdYdGynVCxINqulC4BxwC4aXTwkj3MHfBaISQfFTGw2VCD47
DSYZuVETWtri73mPXIDyHJ1A7y/BvGVj9SwSmyIN7HurH/LH3XS3b52G6DWD1ev1
bgs7XM5MSkd5k7hegihqV8Ef/UaUv7DhRFF1RlrnOMCRRWVvTJs53MseOC8SOjDB
9zFwNtBl0uMlv+DqteqxbA5XO5XksGNyZ5s8QKCl56X6VP4YX772/R9XPTdo+lyi
WG8Lj8kfnYb7ghlfItkw4CIetWXWk9dA0AkWzrtr8ujfDEb58lVeiEjeU4ap1vOy
diFBnIvsnZ1U5GoSUEpEsEVbYyYNlQJ2f/qc9refAbtfI+5cU+qxxEGVdZoNtJQz
il+fckvjFI5azx6AW1jwlRgyMHA+xUx2yXShDvmN4NvV1G7CBUC8jwZIa165cezf
yX6SdgrKPiMCirMlS5b6E6soCfThwIXqNNLdMIh3lx09UZCHl6JhFPI2tdwuRbSX
f2VkTOt0VlI66gMpUix28yhrRQPHWV3gD4xkQHUO6jJBoCiqa13n9XeJeMl/qWb6
3cL5T7eOB5bj6nqktbusUf3KEIi7j74Fv39uWBhhgHip+6WXT0tDvj6s/NnNaUCh
wYp1IrDi58IwQJrdQ03332m/YpQuVY0hP2xDSw4Zaotm66k97BmF4IfWGRAgwXb3
y9z2Jj5yliAKgox+UlIrGjh514R2luuWLmg5XblA9LctywRLaQbHiBHbqSWQfT/9
Q1gUV16Rs7UOzlzSIN5BsmdK+iB6yCXVrZO8d5c9rY9tCOTmRZCSRvpXnL4oGDmd
2PaxojXbDXK1EuVRZ2ffjtSKRbeCl4P2iBKDD6KuHmLBNO/Tm0PuvqTcytwiL03I
oB6C9V3aNjwuDTghBMg0t5C9NbGYrxuEac41xbAqwq+hU2t1RrVe5MavnFsio2wM
pkRmTdGld83HGZNsuPBhaeKWKRlFWUfLvubFhWxK/vUxo8I8EbdidUMuDBI/ZhQ9
OpalGEZwo5/mSML3u8Dh++/814OGMP6X4MLbPMHU/462SOD8NQ4gH58uRfJDiLB6
7t2cLmtmaT1ACpLtI2TCE4P5WPBaTJRwW9Alu9H1k03FNkh8fPnsS8aberzqorB2
iK18z42dx7eb1YTKC6peSA==
`pragma protect end_protected
