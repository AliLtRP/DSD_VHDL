// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:33:05 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
p+T18dnkQXPn/a40ewXcKPUJcD5DBHZ3ByAs3HBu1aU4mrogn+tztQIzfuN8ZQO+
UTN1q+qUbcAP5eFPfVXpnlByNQGmQWoGBVe2V1Lq7v/e0CYV+cb5rbm2VzUo3wCP
QRbif3FFJIQhMoRU4JtEKrzgGZ/RqN8oz2+705nJ0Nk=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 17728)
Psf/Ow8VpZh1a4pgx7mQu8YrQYG3s2/w0LUoSR+uYj3Kum/xiyV93GxNHDGEmNmZ
JQ9FwwN9HHV6qZJHJGpgYA5f2Q3Vg8yuwvCbPx0e2egH7FwclALQRs9h3f0DBdvg
XkUAXdvHZ3LEPDZvhW0uimSRtRQ5bKnh8VDVcn92klbYMAsfQ77RRE0zLqK7Qur3
4qnMr6wNGGDrHQTb/7pzLuTPicHiEX/Bmd0md3iu8TV8TcxtmWPbuFA235upN6hG
8oLXJHRhbC1mOOJ3SRbYtqvFOke/91Y6Ow7pmqraqABxWoD6W3ro37ZZojV1rDow
TDa3SY2Vgs1AqaijX7HY53dKBCNSiw94WRGS8gyjPhzi9JSl7MlXaPGAqlpJxLUm
BfU8SQewngwCHrdyw4eUjzToWz+kAQWCfbmsP1K1LRjihI8CHqZclHJXiQsumA0y
lvdhMt07JDqBIZZVZ2Tw7aCoKaF/854vH16q+dWTSkkJ0AIUurBJKWVgO6IW5gua
SP3XV8X/xFzKCO6K9qjgbHw3k144mCbqpBvfNsFNDEOjt7gvLfX/cJjXNXgMAn2v
rT1oKFHss87btaiQ6drfPs4OAaM+4aPhn+/lesjWcFOBoxf65TpXvTR2EjIZcvub
dcRPgF8wMABy9f8Y235jZq+aIfGws7NO50GSkQDQ09kXVyMbQt2pnh92QKnsQ3qK
A11g5wk73fhtSrWgW+MTaffpMX8m0b05vFSuQO6TL85geiNp/LC9cggueoJFigcI
WJ3YNGTFupS1tD1MSKQSHuXl+kRf1KCNIgU8z03lx0vWbLfe71aM5wVnDzGQFsaM
MrqA3Sy20sdeupT0oh+Z/S68oB+zYGmQ4KB8fPTR4KgSEw/a3r9zYH5ZXH6nMGm8
guiuwMr8beACKn1Y6urwVQG5W2KbT/3/j4/M/07dlfnm6aQjIu6xatV0cs11/jOZ
HeePQ/JfrBrcnPDNF3nKuzWoxZxz1oGb9k/f9t8a4/WcyrTwZKPaASa/NCGxD98H
Tb+gouf9Qv6OvHGxEAuYxZKHUAboH95S2DDA1XxWztEjDPb0JZoUJe/LfuZ12jzk
AZFHFK+NZGbEYQF1EBjMEk/nDCJPUwIzOht0+i8i9pmMAlDbh/3YOXraJ7GAuu2Q
1XQlxyNGmBLtSs702fGEr4pCBuzUtxZKu7yYmM0Qygso1beddYQrDmhhsPqnpEXw
wlZCtWe3k7J3IOci7/8aACQ9/KrECgI7Kmc6M7f4RAVCioCyoKpk8D6ivZhGbXDl
hljc3p7cNCLAdKmmmPOueOsvfVtpRIITMoapg5DS+MhTPGYhwmTdzpHyRlwF9/a5
HdZWA2Cir5H0qa8yl7e9xcMS5atA54H6u51695C3hCy+OSPqTJ0zzDzOqO27eDAG
l32CiAI3C12YBVFGwe5OwZKD3592DGltJ6Mlwrbj335uGmCQbSGfYH/aL6SquqLu
2Ib5WtHwYTd+U4E8rtFkkVd5LLFwjzP4BGxBfyQDalBnn/B4irSaRyVYzrB6vqZT
+2SwL4kvXVRiw4o5416Tf/rvjtHpJan7IztRGhLVCCrP1AnM1WC9JsJjge+B1t0P
7qCI6h54GXBJhDJKgtp4R1D4vh/GgKCMoKMFH/HBLiug3W2LF++KI91Pk65vMIPO
yKz1Ul4fd5Y5FFbStGic+/R6knbwZDCbA62s2sCJJBp1rFII1Y4WAN3vsIssjZ4y
PeZl+a6b6vArcCIUlyIsIPiiKjKraOzZsFoeNWKNY9tSaqv3opBNV9ii1NuhRokE
l4lX/ZJOOuBdt9IRs8WodqVT+tcqWviGZc0ANXkBhBFHxeS7TCXOOlXuztqmtDwt
tWczXRJvPmHk3054AnBgHLty47LPfwpt97Qv/ogTas/+8xR6gnhqOe3JW/zIel0k
4U5dExOGhEMuee3RREXTkCiWSo/DSChFUPQ6KOjrV/OeiKLvGgKdE9SzexGLlnw8
T5UcG2kbOiK2KOM08R//IzGXg6P6+/IGz26G0QiQUGfJSJhtwYBmw6rDThoFw7iS
6UrIBSJ/s3pUozhL6P0uSYoQ6/32jQ+0FeCWL4rXxlM9K4snBzIWB4qMKcPxHouy
zeLw9PBN3qIZuyuenimbqZxaDO4+ymSd0Tj0JRtc+PPEWPNWRzEnXH1P0DLIjUkQ
zwLBQ3lUO+bwVe59TUk5PGnOsluBx4UIFUF/8WyJMirw1Ap+8LLyja5SYISTZsYT
k4wXY0+bh94dgGdLOoOcXgm10LX/pZ4L0dcW2j0Y4S4/ZW5YgdQTzQlCdnCGm6vV
T94RgWkpsdma3r3+KW6SawZ2cDddA9w+hYGQWBhw4JyaU94iTYOEmdCMWevyw0SG
rco33OtkqVnANyoln0uyqpKdzh7gfNAhiRb66+POicN3VFDcGrpaqP0NVzlWVXfS
ppAsbWRBetLpYCvSIutPhekoSHaqXv6uD/gZDq9ehiM+cgdXVB3hTuvUowXvA1Vb
F5FyiTm6Jy1BYNsP6jdVBar7GlH8Q7LuH7ZIUVzTVVc6Ah99I75IrJFNlPCVOwIN
2hBVsKTijNmVlnMaUB61w7ZgztDR1/UzZ8qZmB915qC0LruzyS7f3EivGhxWt/wd
IaE55uV89+45qMh6QG3zgL9ZfFvraJTmRXCpWBt3mTqJkPJCbFBnwqYJkxjGAUeA
hifmhqwhLRiZ+fZoe5R0ECDjbXOJCUHYQWP337krw2gVn/E9E5flQ4XtMv9oIGgY
GuUwOAMXbV6ewSJ0DLNol2b7QJmbCp3Hprm1cgDL53mjLs4C//R3+pdgSIRPNNZk
ArPMEqDtyIEA9TQXRWTopNp7X4XkBAZFr3FS+bkiO978ipxwmQOfkBgK5D6tGOxO
+jyqsjEJ3FI0GfufbHtlHx1QdCvvjuBuaPapiYNmeRFkTZN2StEP14GyWTU2gcDS
KH/74xE0E63mZXvv478Ft3XFEI3/QtfNMLh/XDx0FJQNIr3g4jGfZBDsvtV/Cj0L
6qjkRuRt/nLyj2ghKUKHyA64CtcQAusn0jL/CHJ5RUh50j2osrlSpF4Yc8C3j9wc
sk3BWrgmvlbPSaH/AjwToHO/JlbaXmSyZHNhZfZwjtdDYe/Zk0i5Q9R0bXL31BXW
xdaAaKESKL7+QZkZWZONWJ47bvGfWKArESvRgHEWF4/mGgku1jRmaGmTvfdweje1
Tzf+lniDnMDr0nE7R4mpHO8LvNFTYjz3RHERaNEikFml9yC2m5ch3Khr+Az+qctb
Tmsb89VuQT7D/aSe3oXfFrY1vcPYqBGrD48pABKXUgTQNBWrYM8/BGbWy9oql2sG
UvJMPEn7ZijHOHZ6X6MuLlMKvyYfckwQog6csTQRKIvg/p7AF0BoDuWqmOU+uDqj
9/xLCJ9VvY3y6fxjJBiar3dWkoPVnaWi6A6E+lzV1SUplrVhtq9jdaCWb7Nrbl53
ARTM4QZa3swJ4CZteBoX5JU/5sTBfmmvSTyJDNPjCWs00vDV2VBwBFLVJkJMded2
892KeoMzLA91JYtaazD0sf+XX5aida1va4rAu559opPrhwaOmqH3PeV7YfRWG5YU
9u5GwdXH8ZPAQReRP1NizULnXkWarrpo5xf7qpaGAHr+73sdRlqVDBdDz5ttUyVo
OPA1vaOqYsFeZa2JpJ2pm5WM/20315xIa1kktukKkZFlNu9E5/IJsVOaFGcyKUYT
xeHcsC9hq9SLiKgjnu0m6lPP5e7+ZPmlVo9zqCiolxYFUXDX5LfJS/xWszQAuPJ3
Ne6Ndp3onpi703NmD6EvcX0A3r/8JHOrYRPsUUt9E44bT9TyUEj0sUjP0hiNsu+4
rY3Yxf1nb/FfO/FKzQ3/ln6yYIE6NaUeijyIa0VzLelxbJuTTbr+uXTd1dzp2uo5
o/fBYDkdrQLNSSQl99zQUtyMRJ6kjBJ+r5wPw5dyMFQ3j+6nYUOzIMLFkjCBas98
ft66PsPxp7eUZHNhT7s0/5MdBllTNu+FyJ08tsdVzsyweWeSTyltxrCnOEuyvP24
TgJbcFvjgupeU2b7DVsihqctFSTSBApTrWkrqKVMNH9ajfHomemQ68OJ21z6EoPm
jwFpPtqqDSU9MXEx0jhhnCrIFAvQWHRnLymluBUQNenUnW15e1YveZcJ6k0VtIlb
hL88tH7cSTvn5RvNxKPmaz8PtgKkpqKWufo9zQR4CdTUxLIVlszWL8laTKk3w3l/
gCLr+CG4SRSH67LpxcniMN2pcH2qFo7uXi71/b4dWKDwNa6/aMEG7AM+3ZGxLEi0
0yAo5wlDf7zO+/u4RA2e1JMVMrPkvTjs9TBXae0Wm4Q8gieBzhnFZRfScwmasDAC
ifNs4icKYWsv6rfqjcEV1/XqaQZVaASOOADZgGFsik38eVtm8FmGrF1kM4oWAGgd
/MuxBxU+kCVuqEB4d+0C4BlE7XtNU/eGkb3+OdQ/sPWv75cX1B7FbgBBXC/2bDZv
+oBiHT6GAf9xQ4QgfTlRrP5MJddURjdTHwsW7oC7QobcioFfq9LXl3MR1UI4hMN5
/mUHygy9Jp+hHp0c3AKMARdkXvKpj7FNPyDzlss8ccxZmvRZYdAwxjsnoxNNBKsL
Y+W8U7MTs/+GLRWWIJzjs91kEx2DuyAvG3t03nW8A/BU/Ufl1nP8rQ3MvNdaGP9m
Zm0p9qAcnZTc+Ql33dlV4fz9+X/1JCfrstp9KG/uy/UsT2K0zou7m037VoDozK6t
06scs6LsRnyyVvXXW08O8sJrlCQ2WApFtT3OwglDE72i5mc0GFXjul3VlQ7sTSCh
SuhvqD5Yuu80/twWaV517sLfpSi6XBgJ+VxdHSAC5izG4ZQDmGE9Qwf2BiFvIge+
Q1XgubjaQBa8qHvBPulqsm/f4N+UOy2n+zTqI3yNB7tKp3VXB68T9ldMhFWofRI4
y8CoQNNsh6aVwE1I4P9Q5TqAfCGqbJs2upu4k5+TAmEcTeoS9Fi7G+fDKnszKAcM
7hbUXx13nfDmPq8sCWNBl11gfTjjfCgc4iZ3Q8ghXnRvp3A20klG8kAgPagd+nzR
xdvBAKpDdANtUD0sn3jPTDDxsFd+dtdg9gHE/yQFxPFZ2jKdZWeCbCkOXLY6KqRU
yTRqoR2eCi6nGp6tA1xSYPTvTVZ2TVbfdfkive26jwF+w2FD+2dmnKIinh1S5Clq
RRq4YRoQlBkn+o3WLEIIOKHylrVCSoWP5vOgmYNC5lCH6DiFHmKQTsOxkHX0NREs
HZ0Rp1Wf7dbE9gt6xtlWc5LtRVZf3kSjUvi818yCmA/khXYu29dXA9fBKumpTjcM
2En0kvRgq4vhupagZxvv/Wc06rSAL7cyOT19NW3w3UbAhktPmusIjZRYXMl3/L91
OkpamPateDq7cIMVlltoOx8/mgShwCSRf0oE+c6nnt+NFWRaAYaYHCj4Bx1wm9q+
9s0dHzdgEhlYAMXJ/DHJxFAyMZGG4vnclYyHmAOSpPdR+nVxmkoH7RiaCgJoUvhy
+J1WcvWA4wWesTk04eMW16Lu5wQzGkrJ8yBl9Um92DbzApOFfbE3yyEJK1w3WEoa
G511DSPmGvn7RbNH2G/QNp+aByEvclYnG0064gB56tJlcB1w53y9U8TkPPYpuCWP
NOeb61PbpLOu6aUOXu57w1oVpooB2482HJpJ7BgqY3Jy3SY+LyMpdhjPPXXu+itZ
ns6kgmvZSxu0JMnud5WBN4qgFOIYu9On3qNLUG1NvoyRdNlpvcl5S85RFpvAPdOz
hQ3f3xpTE/04/1JYkg4/yDkJFXK815re8F/S96tVtgDle928Jal+ocAEvz/NjOVX
+bC7BWFk8wFBKuWYkO3ysDMOxn0IQ1QkT5prSnkdp1KocB3oQx08LzfHke0too7c
6MoSdYm2rDVPlRxd7mxcg6M++TrDse2Jf2BIHggpbLwJCo0rDbL5Beu/kAG8ZzC8
MYB7SYeWt4ohVZS/e3tR02ObFqVnOymUGNvEDCTLW8+/f0qI3UaetxUuKYTLe6wL
cvzEcXcCh5EiZFmm8DkulLzdlPEUImzUFk+nqkTW63gxrVIq+4n8H3hnj+cqaoKB
69uqNLODyZeWkQUJncOV16RZegC+qiWF22hkhcWo4vujt0MqdTgclPF8qWFMvCGK
YWNPTbwVkZLDm6NumG0o8ceF4Bod9VskWSjC1gyNYBdmaC+luWtACzE4X6qOhr95
TfNM144BJG+uJ8wCLchXhU+vbJpVcjzS5kNATEZZvQyl2gMC7f343fzm07uf6qs+
hqynkSQ1v9iDkwqrLgakkP/RMS6vGfwu8hkbbtJWTLnnHowB4REUtnkgnuErvol2
LNeQyCYgfRRNbImBW4Os14ChxpIMubDQahRek+J1DWJl5W+rps87dRPzH2Es+tHv
WwwpTAliFS5liwCZeCPUVowQzgARFnhS6a7IhfXfQeNqwxNTKLQ8hfvhOv22ERmt
LhtyUSQ7fFmN2iFIoUmJMXa+gShmNsKj3AwNx0ia8OC1YDeXzpeJoCPHuQxuoroA
TEMU8HSU4V2N4aEFtJgnnc7EL7fcvNSlhoNwYFHp8dDEXg7wx+79mJWr0W137EDa
r/a42Zn3m5Pr+rGPnRzA9fBikTLV5j7h9t6G0hdDaCaRPdA++aK2Tr9HvWoQxJBD
8mcBUbK+KtsYFxhBLKlPokzqwPeZApZAOAZWgvQvAp6HaGc5mXHshi+b3d5AIGbp
DHLDXndrUgZHb8KocNQnr0oC6kuE7W7UdfRSI1WEDPjlS5Aa8/U3q4xEOarR5DZa
20OEtQ/mHQDlenzZlVjgdbMhEGcWgU3bUm0cfjHcFxhxzvy1Bu+GmyXo3kZorZgj
N/qmrw37ZSNN3rXaS7SY/lP8V/VFvbNXse5JKfg/pZzCPkdGXe7dgvlFIHHLEfQS
Efh0ppWZesPGRUspAoYEJKb5nZsDo+q+gP7D2GZAHWBwUTyWKYH/MQrKS9g6TYP7
eCVjeKBTWOrLqNEGe6RcLxXyxeVslx4pLRJbwaUKIgiInW1sz09cgYrbgdbS6n3j
uAJIuroiBdUTngfzn+XomEARTaIWSHd5f8pq8vvicnB5dgWNLm7t/chUDGbPA6T2
7OujOza9tFgJf8XPdDa8UR8AM5uwzhhrYSbeVE3YRlvJT5YwRG0Haj/a+B6UJuBw
+kxXA5kCmCv5qaR8tDGxguHpQK8G38qm+5VbY2M66ugAL6iq/yW1W+rthcrsodCE
zNwwmCKjkfYpV7vZwI6Hiq2u34UEv90l41IXxnfbH44raEVUf+8NR4xXmV3hNCPG
RtKPURBV1aPAGjJhj1Nv29PiI/Pq0Y150iKIxowx4zVzbyuvsngfCf+jb9mw68//
+bQY+msbFMy+bt1fEiKBmSt1akbDIt/0J2dmH7z3rYMsXmM058pruDoaWxr+/lTR
+FPKWHvPYUpr8G9VEXD3ENuc1epBFtd2dcu+nuOKg9GR9FreckV/pNQBPy296Ns1
Ivnhmvi83298PXsctPf+AP5cOw/TStTlHUvtdC6sNvnE48dftU/dkGwNMfq6B5SE
wLVsszY8pkQ8rsEDd/0BKVTejc2n+jWm9j+q0bNnoQJFIZXVSVew0PSjazXxWj54
n6na3YIfkQAGQ8p/IyQEaeXSkebmqhfAHVhavJm77XNf6O/2QCPtowxBoec8BjNH
M0Ib1MzJYLER5VbEU6sEt4OJYZuvPOsygjyZvpeM5BN84/64p2u4dhMVGwtjvRUX
uK3Jqxf0artJXMGlKMgqvfv4mFQjSURpzq5TExFNftDQr1l39snIBSXrV02sc9G5
TwWXydReWMWTKDQLP5/3yrGwXTk5dOzwbBD2qUqd5ybyoXCpXF8TELHnFmOxYRlk
RwQJ6JRTyFmu9HSy5EEvXuXWCQnFKN+reaTCGSz9KQGHip8R0oWc2o89fqa3cchF
e/XIdi+prmp+nNwdft6SV5L7qBFYh3HaIJsSfuS1NVTCHhiOfZhbCGdwPCEdaQa6
Aakl4WsD9P+6bbeXKAe1KE2er77LH0yjXSmhxlxgtTA6INAskgid4t3Mzg0qad1q
KSngh8jevePUbvIvtKR+6wIWOqFQs0XKyKaEihupVg38LwtEblbeHvrB0RB4y4xy
ZP+EIAHQ5PrScwSNE/y0UfPXD45CJj69SijsPwy9AMllxxkzkNb7QkMcbLll1BuG
3NFnxgrhDGnRCqmvuugIDpaWwKhW2FXC4+RJRa6RIQERRY53jTT4wI9usgnnIB1x
/v9jKtmRLZybOABlgAc61lzIS3AkrsNCLkGf1sD96niN8JyKOKL9BPz3oJtc3Imj
C+nzfnnpLo9dxCu2LGrLaTIOY/1e0jJ4VjXuLSSE2t6KCA6Q8dq82MvoW8NRHWwN
JERV5fENvZ79EJvk8qAgTosC1zOcHa/jBitmIqiUAPSRnlPuB24YMsNH0B1QmYcU
FY8hMlOZvVNhduKAbnxGAQSh7B6/+vql/Nngkn5okMrtFUSuK+lvWWM1VxT0SwEl
5cKKqMMnwBF8fZ9zmAmCCO01fACqgc0TVSnI8bAqdll7ElwItQqcqitau5G6oB8N
hg6EFGJEfToILOQ29weLIvVy4WtUdgRvB+TkStE5ySZf0KiSQz9Tvm6S+ULsvC49
9Drg7H6PCpgaXVV0dh0Kag0NQ1xC0uOZuaVgXK821oiH0FJMCeDg9a8iZpO164qw
yGFnVSBbcl7ATvIU81Ab2zp/0zriz1CySd81P7DlIC/Hs0SQSch8J3NvNqtHjub8
EYRC2WvxoN9LkLuvqJhYKWx/v0gQvGyPWFdjNoLgNkq4fExK8Sk1F6auQ8qVS+GQ
YpsPkMDYT79NEMt5Tc9BBjpMJO0QKNMEfgELFhkfs0js9TbR8/o6xCIViDqzXNLk
bjkI0jgvOnjt6xO4yNLRU1hLDvy8TOeCz1dp3krKbK6gVRrHfy//V91OyZuqkKcd
Rp0V27kLg5t64S68d59pqIwXLn1szbW8/uDmWoPNI8rafQfddpazK36k6Aurc4Nz
Ivl/+B5M9v0a68il5+Wa0t/hrfo8uvxHIkCfMNKCDGpY9JDVe0of/gYhB2qeEnnL
Ae9Q6RB82nEodbu8Z1e6OUncgSSFGyBf/ygvhJPo6BVpXBHklKXylAJtbW5GRcTy
GKI819VY9rZ/RZjiuBUMVwjCHKiFKWq+ye3OYMjR6DNjKJu1HsFD0Ny5ZQEWOagL
VfOTL2ST91uYKfO5rtoVBZoS/eKGfgoNpZEM06g+FfEmLy14KcMdxialXsFuUxeW
F2LEKBNZ8AVY/LrHoFAFetl2pe9hvv4l1KpuE4q0j2e/YvUb76hM925dxx7R99nO
WXh8LSwoy7ChxUg5mOMTmcoHvYzv+UsV/R4n06ddLLiYnM1n16PxdSOPSSErtk0b
IsdH4mDwLCx3peIy/IpkUbo9nW87e7J2Oj16OCXMyTQnWEyon5maBAUShNpQedZt
HSt+RktJBmGEs6M4boiUnr7LfKl7lDIak8NvP6CdENjOlmBPcXdc/NVsjBdePVH5
w/Hy0gun424rrw31nYCxx6rVWJ/DQYYe+tjRWz0JiuF/4IliQZ6AV2pFLeKU6HVS
5sPmhBvnbDyl1h6Sr0NDPnQVzB5Xn2+rZCDhSOyPl0p+XbW1xuQhAre5ea/24YB5
w3lHfEsWYcgNZhO3Um+NPJU1KtnsgGP6MeEKtNUtqTZNIO0Wm8hn7Y4er38Qtq3o
6gW779ecyMKOHBHlRAMw6B0Gq/qmJ978SEqVr/9Bzz3VIyeY2sNzCUx/u+DXXCLn
D9KiiqWp1iTxsZfwKOD/DKHKcCqfNjly0V4jIhtrEj6UbkdMTRrQ9ULoXLXM7XzR
UQSwAjkRjlUVHPfHy3d4VIs6gujHyfT0b2I7BY3fuG+VG0Ta1tQKZ/6VQZcpHf5r
V+VR85MLW1E55XpliaUf27NQJE+ccCrBYYaW8+ccwJZnUng7ySOgQ0bcDuY8LEL/
75wwBe6PP5ZTFdi10dzgBFJxDt61UUjIGcavKvAMhkppyro8SgR+QND+qOd1qkFR
c0lYQDhBujq1jVonNy/PK4ujl/WmPLttuQRjxtTUuvMPyu1aL2XBlzXcezAs18lD
8BEUYd4YV1lMqpcFqpzyZOHkeVWYR9T1qGNdSApWmKE+FKUMYfLe/6bTU7O19sFH
libKvPG8lZljF5goXUoYfGK/QNHvXyjnLhCqHM9Ai1tDqN6UvPA7eySoqDkJBm03
WEGRUInu0KK80e6TIWLYrh5TTmizXdVDrU1Ds+tJwJxUESp/iWQcQ9o1OZoOH/d+
4BkC+GNxtIcybIIO9Gpgh0YMqc54OXRPzIrs7On3NurBDvgaTNPenoAqJRQlsh74
dkhxoM8Rx3pMshpvPTUeIeYTosXW+JixJ8diXn4xiVuUqq1q77uvY4ZFreAAaUhr
M+UdBPZOlVR/dDfZcb8XfjC1HOsJgmd32UwDincjlbLdbT9ix/kOEHKi02P4QG+P
865rPMNW8oDEb9kXMKOHjSh4YeCemGbL82KOXHY83VsnRgCzbduJ5xLdIJCdzeny
TX/j38p6Vx+u5CTGP156ANd46fhpupiqT8Wv7s8yTzFRtVuAIK78PBnQrx7x+Dy7
Afw+Df937E6YEFeQgmntZEFbq/61JG6zVZpFVrRdnkTZMRgKY8l+tN2B8Tu5ypGF
2G2z2iTzWuxsW0ikQAv6Y555Sle4zuPiGqP31QUMaBnMXLa4OvH9BKsAJoGdjOGB
LTLZRWAfg0xiAjflc1PeQrK0Q76cpUG8EFF5yaI1vGpb4Nr0B4SnBy36wYl4VWRe
dWtUdWe3r4dPNqVyCu8LMAxAo0hdVxXu5/d0vdFuz2EzU7mYlDaVFTGlmDRK0oWR
UtvTWRxUOnJHB65kLOfh9tCTQ8C1+Y6UQ1N5y8q1lt190Nw97J4209oZLxd/wkWq
TBC9nkdC+gCdiIXWOE6lPODrmVHNx4D2i+DrdDIOwpwZjiz/e5no1dzSpmTMgCbD
hYEedWL6QUuspgywJn0qYcHSvU01Gq04J97tkKrhidqKSEnmEVtKJ90eUzdtfS8d
5Dw6qMAWtIea0viCnlJ81f/h3rRJM+JAIdc0fAjZG7hitm8I64FLgaEpM4DOv4Qp
grKUfk/7uk1zAC/kgZXfoX7s+c/lu6QiZcSUde/psWY9JDN64+7e5m9YCdI2b9/M
jcpdVwW9TMcI58kiYHFbCO891bNVLb2to5D2ndT/ueO6XHR2N59YMiaSc/76Bf61
1NLGie2D5C4wXhZmvCnN32GFB+lnTuotLVOUQuUd9wMts0fnltk1CevrUjlb6RjH
dAVuMbj3mz/8hxcXmy28VIs3lT2QKoQMn4Tx3YrYpcX+29axaQFN6AtrjaWoBoHm
B4HEWJlvq+9a46eksvC8aD+SV+z44Rng8pFHf7jsGP5REzeUCYvf7DKjrSZi0mBn
EcBj8oK/8SIf7BT6iy5lWCcGvgK1o8V/u5LQdNV0j1b5MW2Ep1h7bv8/lClErtho
pi4dxazyls8kIfIK5lqvj5PaarKN/gfkxaD25jbkjZ680/3JfyRMZEqn+3j7su7U
IssI3Grabj936FVf5j1pytc7sOI6RXQ64doK8KWQUOw9u6z67BBlCmrms/y/YQPL
7OLc8yDvxeN2LNBUESZSIHcHKNAVRutGe07VRYCp26b4+fKinSwOwhqbGeWZyhOM
ksN4mNZaRDQKRQq68wmtWBaNdHbmxy3Bmgyxn/RZJZ5HBTNnF8+Slmo6au1TQpq/
aiFcmclBlXpbttMBj1kAKA+5Osn/q3MxeLXa9EgsBWqFuq7Tz6ugNl+LOSKSqYJu
YS5YcOnTky+RY3orsUAHtn4n61qkLnvepQp+FBJdMD1Gi8gF5EAOgWsPOZEgg7yh
1JGO+LLvU3xwgygsP/bXe4dO6oaqjpgDhRlNmGqB3HVqiopWxcuJOtMl3eoLL+c/
WCO94gb4/7w6MLryGk+NyIpXb48nw4lZLMY/CU4h0qlkJgA8IRyzFTRYf+usVr52
K1BsIPoRiZSPTktpV6TMRkvZYWca7sEwk2LBK5qauWwLnogoYSMXhJjwyjHXG+qs
f04Tu0IAOrL5u019BvudTCSnEJG8yCgSntIJ3fOxfMRIa/4WLbWTGzOUWdxZNXVT
pqbdL9eDs0es7nbwjwgDkQvXFAAJmhNLZaj6wQ6J80EAiQRAGKj8rotHV/yCQDtP
RixGduCGlWf7NdD54VM8LWiLkrkQmVD/VX4DOLYH2lOm3cj9JUPnSUUQJAJKGsYn
oxGCzirhSeC83ru5vCujlDGdrTPVN62kM0eZ8w5iq967aJKvTIHranJb3CrS1GCy
C/M69VyqPdGzYjFgGV3mY8W6NmbgzV/2stkexAzVZyVqtBa5zRUHeRMp3XKH1UBl
kq0zT6PRuZl+0QIwM6o9fDE7OBLnRMOai/aqpg9qvD3LovUP6odhRMfCtjNefX+Q
m/a4lCtJQ11IEog5DIZw9ws81LNadgRvK4bY81LcXzZ+WXu934p3LB5m6DRtO4hd
53fs9Yggqu/eE1NYNpdeqVIBLH4CTacisNKyVqkWM1Iih/Y3PPJQJBKrKxHEzlna
rjIgy0YCRGw/2fXXhic+/+8lCk2Q1YBmleRfbDnMBwqqaoeRXCqwVVoYKxq/ib1A
TGuW/dPwhd+3OmpvfA9Fi4GBAl7HKqsYKM7/oWTqljE01++L1ZTTQ+dS7K/0/kJP
aSmfWBPhjl6XPILYUC5HnvaY10F8M7IcYYPjwYG+SzwL5g/c8cC/T/lBba5cp8xf
dun7ETjPF0vIcHlEDx7lECbcBzC+atCqdEZ9sDWmCp/wpODjmX6JP9AhKXsHzha9
BWcACu+IhoCLVCKVOwXtVhfOmJj3cNBqHQ/PPSGciELAPvoAgT8wYUELaJALgmV0
7UDdaeNUfYu1/3YGMAi9wkDicc2buZIKbInbTBgyj2QvxwnJ/rQQvDa2WazYxKpy
aDePbrx7xSuyImpN9cO7OYfzIP6PpC3N3oQBY5+E+41dcdgKYRq4Auq6327yeh04
dqeBH2VpnNm/2IIS1X2gf4Mh0aGL8fwDMJImzy0GQxAsBI/ubVWkXLPbUo3HUbhZ
ezyq6lzrR6n0gINtgKf8oQPbQh5zWRXny2WZzUWRw1/gwktYwp3df6ToJfQqzmb/
/o1w9Uc+yUJA61q5xe/kzc0IOSPqrbmTfA0hMMdeoz0z+J1Amu0FwxFBLlPE7mBZ
O20vYpWgTRGPgTYry8mGyRbSSC3ZtaOvAIQGXYBpaNqV96xh7qMAog/Rn64DMN1g
nl0A35AfP89ZuFFEL7UOmC78KoUzM75vVzawLNv7nPq3IOAwRUfUAhGHhV0svXDQ
puGIQvcZzasUzdHRx/NjrvIwxUcdNBRrNUlHp3SDn96fQrumEVrbjC1CGyYQ+yLw
zWT1bFC/Q5IB8MtnRNxOYZFJL1BaVKdiiSWibyaUy21M9bKi6Po9JJ9Acy0TTiGL
okmmxhaq6l7EKS+1gLYZGIybyU+30O7LcHvv1v+JaMC52tIdopTbUHfPVyd8ZGEZ
wgWqgkms0KsKYigkG3ctsqpxTHdmO5Ko/y5TGqqa4kmWVqZIGESawFf4FzWiPwov
1esSP3rpMt+F0ixJt+jU7DdmDtyIIbDGZqz8oywV5NdTWkTG8rWijIpSXHFvrySY
TOZ8HlMoMSQKX0KjydJIzc41Ze870+BAxC9+BiNbwTzf8uC5BRrbyx/mY1s5PsEw
qSXzPB0yG2R6BK0v4GOYpCB6P7obCCVcw1Mkw/oo2fPEorRPVANecOIz+PR/4cgV
IBQYcG0oXdTp94aC7ImjoIhyHLZy8cxOIJVtb7ecLzD1X9HmCewGr+wRktmUWDkS
aUyGWEOLLUT7JUU0a73QoG3nmRsAi1OYdx52KlUpS55e8Gj1y4y7YuEO8FiAfUAU
/1yR+r1QDBsJuqiOhLwWucpZA5ahqWLRaG5gYVIXRN7zO43PbYAUBwcH+g77TTQi
SEkksxjdU1Su9+Cd92DobGZw3cgOdKo1zoG4JXzGMk3JHBSN/l5jwRC1lEucpAGt
EkFz1xDSUNUtRJRU+vuJemrKHQKuKANrvFqPGA1682zUx22sWxaCMOTQc5O7iNfI
4yApaxNza/d2qQ8L+w88I4puchDDb2xcSFosTo/yAzJWo5GXJ//ZZZiU8ZahjlLR
CYugGXhdbTirKR3ZLbkEVWiPXiQ3kB/IzlL5eEJKG8qk4dXQgvZ5ZKBHeso8bbhJ
PYKMaBQC4xGWhNyXqTHvtJqIjqcOH6irfPshnIw/zrkHFWVAsHEWda5ZHli1nF5i
vi4Yowm0+eAcn+lnyYsLWEPymh5S/v+lNV2YRfBUaPHhtcmgulxgP4Y+WP9wDpbW
ys8hNfmenHfZZS80W53FqYUlHUFjjXHltcBnSNFPnM0ny9GxyJYeKqcTZ6L7uGO/
2W39bOwtSQLG46UxKK7Q5OidFWfRQ4J2uGcLDFbxswGyLMz9+fQw1E3eRvpCjGdr
bajUwwNL02y9RAjtp+9P3fQN6xxjGRGsmixKOai1smkhtgQH7OSYfwD9KjO5yjwd
pQYFuq4m0q5dIQ5A64jY8NmaTxB0lnHnJdWNy+gkgucF7Y0NHyBrIG8VDGezajya
AMNYFf19HfDSU4XKWhGj6rhs+qWYReeg6fJ8pWspOQxhUg9cajwSFy1WpewlWex5
RJ6KenExboF3GKqutWcZ76v+fk8E4o6Q7ImXt7L/t/tOFRO0/lTygDIb8HM2a2bV
JtR5uknarT9jOgmxpE5UhfHTubJOOIKutFxlZhdJIMU3QISwej0VIhFXbtwak9uY
brNyIUvaPkZp1vn37MIZ3HN9VPguzO6y42HElF5YMMFc66cBpAjWjlqATJ3GeSnO
qwLC9IgN8redCYyOcL2SqqcQ9YJu/U++o74XEHnz3kOfAmBTqEEkJ0Glz8qauV3t
7P+jMBGgVFI+Ei0eMiXHGSj4smO7c7XkJAmwCUQRFdjYH2A6XEm2wadFebFIhCur
JcVzY3a+LRiihUwdPJjwbpNMokO8MJqWdeaP05WCQGmJMu8vFG8t7JZXVYHA/zn0
cFzJ03/hQ/28ACMFETHO76YcVvglul7MGL/kvkBjKSPGGYZHFuESgbZQKoe8bEBO
0IaLXosQ1wutJPEr8DEi+nZ0X+/vGF5VbRhe4T/WiffvQ1wd5wT08Xp849DIM75M
d9C1GkLFXLaRa2v04nAgvyHp3TNsQjthbBm/0KLgsbpOb9XWiFyySmNCOIRgm3TK
mkzOqyphTF2NUR80k4GyZH+WLGTyeovNn45MZSchkvBT6TtVqM6UO5pVQowTItxD
tNbIs3o+/TmewCZvVJmaE/DAHpXanNbf9HrHziZZRKB0D9giVmmkop/W0lGlAzG3
tILXr2TzRmVLUN4VJFI4bAMfN9bl+J6EdkTqm/uK9kbCjb9QGZptLRWXs4+L60OB
62rpOd7eG5DtFpR/zQ/+LcPOYZjeDhTVikDlcqTXGzxycX78KmuU/xQtmNj72Zqq
SGXGJwCCne8JsixFowJQlgdRVIzCnr6dffXFy2UMthKT7eL1Y0iObOm0UTDp4c0J
OxJ5opa3UU7T/aZ+er5jUrvaq93Zvki5lCJcrtk0Y4puE37VEcz+Fp459E1p/hmW
aeTy4tdyDi8PYD7EanLJkN82OMsuHRoWHvR8wRsy9EsCNlvEQtQpSHVTPAD3JYSq
CcQBsIPT4VWBtBkKDFYCAxhN1dpDp+6e7z8EwE0hklzkN/M6Bf6mguCFdp+n2ZU2
hyvMt/wYozy5nD4jYmy4LxijwjPVcmYUZtQFJ48veY8m+xquKJPcTP0VZWrusvJT
dBi/DqBsvmbctR6JY0pIElhZOUZ0R/8ROrDJV1z+mmY1UMQAkVhATRACetCxke0X
+arMzlxTpbYw3xWer5CJ0Wex4hx3X2jGrS+/d9tvHWNa5RhpE4hnQvZaNgVvsJ0+
+JBszXiUc+aUrcIcYn996nrhu7kk2g7R9/h6zowEXK01KS+o7nz+vLkYmwpZJqiU
b2+yI5ltTNWomAIjhCnCnHwVSzHCWxmth912R1npN8mtHsxB4vc3Q22fyc/XcRnX
0Lpi4/iH/n8W5oIOmTa2WEm0/qt0oayJfS094vIPcERHV032z0rESNET9cgpbzTB
Jz9rzTYX/z6xJPneNhY1K1YTF1ZF2a6QfiTz+IG0MV6ln5GrqkOCS9zTOwRXclKT
t2/IZf1P+lu/1naf2OvKLGl+ynmNJmVRQpJo2dTE3yDYiJ2/9BSchaJCfAGJOq5v
vQMNbD1VZoIfPpYlE3Z92PW1Ce/80snX3qHXW0vp5B5Hhgt/nFfd8Bef0CudNakW
o6YdfSvqY+3u8JbdPlnhUrb0AxtPjfbVhKl9MqnKEgT7g8WDLMQMZh64LT/DIbZ/
aB+YRU040T0uGlyg3dwu87/hvaYNMSEsbB5y7L2hjDLfN79b7yUAr+ZU/NimPraH
wehaJbWFiywRc6wvLhVU2nHT17WdXexrttKS/rwdHmnsVLfQq5Ul+68WR9fnNIsR
Ja7XgTWTmH/8u28VLbV04hNQ+sMGuuSDstE/5vvmalqCvetROKbhF89uCTjl0IMF
IPJIu/zD1gNbW2w1ILD0IOtwWQlmgnXXjJXNB03zpxAXJpdnJz3cICg3dDJeUIc2
qMKIVcS3MZoQ/CuLkXuzV+wpCT1gYr0j7M9ijZaLV5HYz2dsonGurIXhqmL6pcoK
vB8D+9tvPj1SDAQRU/X2RM2ogHsKNAjQ9GXyQm90uEO7YF4Nw9T6Y8EBIk+qGa7W
yBDyivsALH3BIM/QshKLQIgKFf3dgA1bdddYWWf9sqjZDeLV6cGVM5Hdr4ge6czI
3VdwU8hTxb3Uzhm7eL/V5eOxwhCk9S4A6PSGL0QNorZl8eC2QchCxaa9rLeAiKR0
274Kt1OPSEY82HeCf0MuWJV9ZybNKNGrcPU4QGuykmf12No20n4C0T9Q6GY4lFPK
uABU0donxVzSLCi8HZb1u8ZUaNfe+df9M/Q1gg1Haf33k1XWX8DtZ1WPV+Lv+gXp
RNLoLxm2vF8vQXOX3xhhWUgxKweDEjA3M38+iQHIzeZ0VhaWnKyfm4UfmROPU1wA
Zs53Kt0QbhphCbrqSnx5f6UyC0vvZ+od2wRs5/g7yhpebw/fYQ/qDb955Wj6GPN+
qCYtmqZdNM++92kUSZn8EVn/1abNkDVJlSHblV4OYoI/zqlTNTjkEG4eZPvnJ/dp
22jIVpWyzc5tmNQonktNhr9W6EYr9faCaPbIgvELuszk/aNxEfdD1NR63dJD7RJI
IrC88iWduBYzED/CVb+9EEWFPWMFVkLfsLnl8cXj2Titd9WPJjMG0cM41PmulJet
xaJORazWn2mGwO0Q+oPr8xiX7sa5VfdA/QWQ3MFaIts296nwvdpJN16iIC96R/uB
aMhWCMDEvNjpWZO7/aRtpSwFgGkfR84CuGUByFOV4YxYcFTt6T4NbLKRojbCNA7+
fL4vwhK8eAw+LDsKlvticbd3Rz5xJh1CDyAreIjUjjFGNRllQLpec2uLVFXiPkKu
+GvA+t64gNSGgT0ssXXb8OmWknxgDyOyHQjm57nNXNxCEO5Obi4A0GQ17C/qu0aq
UjbCB2O7SuaMb4LzcSEFaL/DtI5F1XHus7ycbumgbiMgZGD5EnWDYh2NfgAH99jC
NwDezAaz3y+hSmnZEPOXUCH3CHrnWLqCBY2WdDLjPmI8QWYDrMKlFhm6TNQE9Dua
UpZcRmpBGfWr1E9Is0GQC0DVv4i2aPzZ1xUd0MgGtmpPORNVy6j9wGx44p1KUq8v
aow+Ay2vzXrPbJ1rmSKVOFolPV3vUtKBo9JUwJQbC/xZ3Ojg2V5ow5DOj1RIBuF/
HqI7thIsrOo6qBtuaWn0OY5phThQkJGNqH7dltGPusjqlrlwzBuxzE7IvBB6EY2f
45KfeA7sWoQFfEoJSx9W3pw9xbJkV8AXBifHaoZdFLKfG7sjwzOZ9jgP8t0aGt6e
hZTEvla7oYg3iA273LL59zO4f2Nif1U58CT/Aye4gjN56wxb+/R/sC+UzNcrkpSr
zZp/B22VyHr/AYC+wSHcdYEIMRFqh/syuF7+BuMyVWaV6sGoh0FnuYmp+QnIS6fp
NwbynjfnxWBDZBPbmf1DlSz5stYGJpP8SSQDahgSGdGma5xpdR4Dysr4gxsRjmHz
/Hk69NsUC/pYYZOFrA0m6ydx6m6ZoiiwvWeM2I2gCpt7Yu3HtMpOJWQ1ZuV/7Txo
0v/I28vVcmFV3zNie/G0g2bOMTeEuclSuIBk9OWdV2cFwyyc6SEl6RX2I4GcQbLF
u2QHrVuQBr/6AVdhz2fx2scCa9A6ZVFzIDdo0eDkOlPSALktYBItrh5SMFvrf5Gh
w2P6IWQ7UMEcDSv9sZLnNnArSPDbog6RyTXCULT8lFMKKPIIC8BvkezGip2NwMoC
h2tuI2N9LkBZTxOmCwnb8Puz21fSNM31II5SBVesgdf/sfevGzP9nO5NgZBNhYUH
31v/5w/koWnP1XroBBdOqr1ElgrPJnODb1RPq3PIse2pm1n0QuhkgAqo91vHfr8q
kv/p9cvWkvccF4bfLyKHEV8zwgRSd7pI3hr8sQPNg1mWgnjQ2aIPVB/wJO855b55
GIM4zglcep25NUP3iztxNl7FWO1n3L8oQJKga2wEYmlTS1efoeZm7bT9Nj7Y9qwl
bCr3r4nVHfJghesdJP54gq9tspoT5x4iwShC20CrXYWN/iDYLxzl2s+a5NR55Te7
izxODmg4R7r7uPgZcgdSGd4n96cnl7albaCIZ9HrbsRGaHx4lKgG1k9P02l2PnKy
1/mvT3WM/0o+SiNAFmeVrzyucnVG6D0A64ZS0JA07icZqffKavCBgv5l+k8PznFZ
YnVvmdXwVbFZivhu5HC08aLpWBEQYIxxTEzR6AtXFEJnnN0SkKeHxDR48l7vHEeZ
xFUrB/1Oi/6wvITgnOIKxrWV35BEIX+Ul4WDiF4+vJTR6miGUgzWPNOGTyOBYzm0
T+KNEugWGdumVtpua6VQcidUqKaMXzaACHxRmLrMFKV5LVJJ1EkbQGtnTSQNVCw2
xMF71j1BcESDGQhSDkas0EpG09YCtb/CZzfzujkXknJRxcvqH8awDRrUOaI2b0AI
l4XgZmgFkVvvhjdKgU2YMhPoszoXB9yccbdH+LEMurC7MSf34dqFjJGzTq+nd5e+
vm9DZTe1uHnmzA1OpkyquLgSegtLp44t8minwqg7BarjLPhNucT2lKf0BF7L0lLy
2a6Kmp603BTCGRL+2JHh8uiyUoV/0+PHTWJ4wD/75+52nAGmQwP7fHpNazMjYPqb
jdcMBIZy3bukoXBUnjhzTMq6m8rRkL/yFU3YBwDLH1aQ0Amn/hVJVYuogYOsy9Dl
nn6jcmMPd1gsi86mFiPCtDjfJy8AHEhie2k6ZSnAy7yhmZvUmekQdUTXDhzlR6ff
5eeVkoLCxXub6El66xh4/8ODe1emLkKnTxlKzCL5/wbibxHfKpCuRp9l5wV0NAdl
BQJ/r2xjOP5xTsIKArV6oL+DNe7yN+qdcb3Zp5ubH2z9CeXHsrRIPDKy2Kw2L/nl
zuSWGxa78z+kx3qjJtbzLBA/z870eGWmHWAJIdUl0RgpuQyL/CuHfWphUTHwMJKt
DjMrdUumK3jltYfdrFxGwojt+IUFVyTvX2mq2z37YFXMpUGPumV1dNGqifrE8R0i
5+Iq8FROtuwWNKiyaHFJJnQaDG9IEFs3gmpvVsqGtyW4ZOJjd2OuS6iA/+T4n6Nk
Fx4Mn7Xn8zh8LwaN24pjvEHB+b1Cjl8BLb4nHI2mDw6SwdvT1/5RQt7JzPo4bzfI
PDxsmLkk1VfVvgxxBcMO6nPhN7NkGsvAYqicE0z6rToip5vWqvNdUixTu7PjH07L
IaWu98+jyLbOUYKaS8wEiYb0dGOWpViwI/S+6byK16ndWwdfOfGuEweEhYBZVcvR
WOZCNO9hVB3rTvYGPB+/AM+i7V36XM0D80muFb0khJQHXWBOoD0a2ZT1Kn/s6hcz
qZZgpgLKB/cS01Zv/h3i21in0InjzGe9KSma2GXOZIed0NkOCgwEOgjnXVGrtwd4
4JEgn0VecfGJ10kRNbHbOg7Nvj7F1sfSHEgVubTkw0mQrmKY92TDp/Og3ilZj+fA
9iHzphB5MjVsbNhUPzb741kfXNnBPwq6hvshhwtDvfYtApCH7IL3N2JJLLKIcQmY
zUZhUcEbRLePWz3PhuefQ+b4CcrAgcEZeYqccAss/LHh1GBAJuiOOOx2BkUkb2Rz
RXoVUT/3dk4vpWNsK+ijPr3uSYk5rtdRCOvzgm6layyTMWe9liyX4WeBldKnM2i0
QIEb39/IrdwEZ9pF4FxxcjWbmv1NL4sGNnZ6kDbkHV7+Z1AlyTuI75V1QdTf393l
bmLWRPqrkwEus02PnQrTmaFGhNZZ0kci+HYH5mm46nqKpTp6G3TcI985iEBIj9fS
ROYRYJ30sblEaua5UBE8SzgHUEferK1jU6kNswjQZvuxW8dLWAXPETPGB7e0/+kF
s8g5jvC5JK+K8hbWikowiYpqjHAiANsk5cziF0gm+b+2xF2uLRrTnbqnlylA2qmn
FeyNfYfLQl3Sy8xEdoqyL2k8jBHf0fJ7ce90GesyEKDk01roDUxMERUYMrMGUNca
ahuMHmdlwJoE1jcUmNrB8dKHB/mAtABHd8i4lRWqkHYjxYSRmQEkti9ZOz6oVfLl
7I9zZi0zv6bRSSsfv3Y6HxQWdw8bMyJruMsV5+9O4RN5dnRxHRG+GOyA04hs9ZYb
soM5nikDu6zfGJIwVetj3ezQq5F6FHhhGr9OOeyby+gsATX4xLXFX6wmittKi52A
WGp8zgtKZiyFld2mDij+UAui4ZgYNuVPSEStDBv5Z9RmiZECWVRZG8QU0G+6F05Y
vW4XuPBP74UK8uK5IpS8TwJ5cQt9e+QjxqKiLmqobLOUee5eaY1CNqO4SgzMszH7
SJVq9vMylvTfmopuX7TjD0BNtkT7ulL4ZMOmOXuUeUDBbSdXFDpMpS/HKexQx5yC
Iuq0JMLTSm1EXzRvp1aBHUIsmr4D5nGVMHKtHaa35ETVNOgScViJ2CVV3e2St+lX
VuZjn8g8ZnLSr/NP0baqk4ePptR5ePficmwDN7DCjvtju+iPd2g1Si13IWe6s1+t
qR3pJTh8mgDLmjzfkwCEjMg1WIjS97/gqUVqaHy2ZPk+qmmMVFvdZOL+yPoh53/5
s5BF9hb2lmp9BdZmPc5wb3Ccvzlzode0IIE6pwLfjTnuc+GNzueVRYLWncsiBf2T
IobkvUnJCW5e3tHi8QyIDL1p93TCyvLgIb/PxHEvdpIiQvu8vr4E7TrUiNxdnW/i
wJbxdRD9OolCE6ea6obt4a0eqAZOJWkI1kEDsxcem/vuP/N+qOWpeLJofwwTO4LW
3jWR4vauTvWPl1yBRcnpP5XVCQg93sbYp1Kh0w6GQTo8L2I9srmsq+1xWClmzv8L
HTtFDyTX1qAMr5DFG+KlIXsrNv5FBjq38u795mCqA6rb3qG/dnnInbBxvcMgZfSt
tG2xjezhNJZb+8dTlrtBuZNi+HpGiMwHE0sti1EUxxP55Twe31XMVHNkBC/ipmv8
2JVa1W49FaXPuqOB2ZS9uKs3vSCe+w3QiVGGcQUwFc+7zmZPrgoMQVav8rvbL0wg
SNtQ3ufu0hB/d7w0DVGeQpiBizQd1DGIxwhBIcc984fgPkMnnzan2s7BLS+wPTou
w/dMO08nnNinW6tjszC3rMNl+pg9LB2L5oxx1YhDnEifWL1mmB2GDj1RQig70RgC
2/6fnonCD6Xt5ftzDlSU8I3ldDBrSNyxqPrBA8jjwX6dshcSBw5DgLSImRs7Y/yh
I+dfBOE+IJdkjN8Gtjtcvhr3e18NG0M2eMZLQ6zlCljtzBZd8oX7g89ezg7Cog+3
5jYj7yohd23NXTBktK/OqBRR2hoc1qOng0MhygHy8PO7rwGBgMWusxTezOBpQLq3
dgIIw39LkYoqZhloZzSoFhJ93tJyE7u/msv8KT3yxIdrm2ARBanjK1NlJ0MVF6l8
+BpQzHgCNMUMf9Eue8n+WoBxes7jfAZ/nh0EpnVQZ8v7v5HJM4bFqz+5hNJEb9io
vzrlWg+6HciNQh4xfA2hDSQbYxpI5e1DowBROM61PttsjiDwvWKGyRLPHRf9qHNm
jVHtFXPdo5MIffEETr3HcMHQviFRy8sCZZXfKy1/ELMlcaMwAGCK7GjrK2urmmj8
2FcJksP5OTEA2ZItdh0vqF6F/Ipw93SFc6EsZZht0zqnQ26YK4ZOE/cYHRB18nAh
AEPSrqmPWkKXfwixoTC7oa7cLydtof7q4oxpZMENPCJiXd+WkgikQC6A6VPEbgCb
AQxuytQySwyQU9EfBtswmHXnwnwk6DDogyeaT6itzR5T9T8rJ5ae7h8cB2tGguDq
w4pR8Dn48kEtcHkCUUbub2sTm4JaIQYZYiEwNYxo+YSrckfHTwmyCGNSk2W20jig
EupOlN3q+3mJaQOybUvKl8n0ORB7YkVuIbRZzFsW5vonka/GrZoqq/rwikhPqhUL
RS/AYIgTtF6Z+X3kTq6aJSj+sR840khMRhCSpETha5WBFQLVFJ/LSiMXspUvLNL1
27kvJaPEN0cx2nTDvLHopKB2lSPvp0+XwDToQpfz+0k5Nf5S1P1CmDfYg/7fAYlo
xFyUTbUMG+lzd96XZ2GScihlGjc8qrMbAw2BOcxb0Beayam3Rnf5XExcAeZ7V/Dx
udOkh+GIIidus7QsFXYrh0394QyGqSYnuHfvHac4MXkjczypYruWSjdtYQOlH+rY
JtVMnejWrd5jBZAvsqY/bPtFqtZGxq+i3njrUEhOOLyYabUqN4ELGYS/rI0YUK0h
jE0oZ1+Hrub8BZXr7hnfFXpcGRuCR7DFwj/0FngzmC88ncgUtGObKA+8Kjm9Vgct
+Oj0IpdSoZt6JlBrZW+LdxmRyZM8RJcAqp3P2NCTUQa6QxDoxDKlaRFAFMv9bAXR
hcEqP6z1WqANRh7KzqgKicJVwUIGDlBXHndqjkT+RXNqQV48r0xdfwKeqtd0tWCW
LKAudbKsEJASB2fltYOawTgaZnu6u927nKKxNkDsesuj3qrDsVFtGS44yGAxID91
OkvmTG9Il44VDG/AZoZrpoxDsT+njc97IFlegP6dz03tpCdTsWzCC+FYlnor2uK+
XvikYBFuYgsv9jDF1mj0wDiRxzWBsfOuIk1Wg+aWLOYH6hwcCdCwAchVPcf5T+9u
l1NY8fYjdUmgdaFuJnESPyfb3pCcuCk20ewcazv9zYsbWaVmyZRs4ZqNOd76R5nF
1UNR/I511Ss0UbKx9hioJ517U3pXxu4wlynsdRiRjV3CMMdIOQ5qvkhs0CqQDAYM
uPqM95k83pg6N/TLs+6qfxNu4n5rKVPZrbe262o9+0FIZtx1nJpgan3ec0t8ZLTt
rohF2+8hqIyOV0W3zIlFQB+SJCJXnjGNbISZbCvRSwi7DS9x+oHNq5fuPMhdQa/c
pgXmYrTuidpxXKB220xAJQ==
`pragma protect end_protected
