// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:29 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
KxxzjHp/Lnbij2awBtWf4HWi/ndp5nJgqIa0qR6F6hXLSO0PxWVCa+U2bCOw/qPO
9LyYrMFU1ZKh2xT0V3lYhiKIXfyK0K3a5xkhVJZaUK2i1/t6GdLzySnNjwhId8q/
B1gyMPJvtSVbUu6NqSkgWy0GbYaRe1D4rDtfaOudWJU=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5696)
oG17WwPrOH0IG2L+8e3Xb8hwyQiber3wisHLjs1i+t6jsxTeKVsRG1BGcZ0mKaF2
JnQO7oraUYt5aotoe35RooxpibMBEPJS83KYhzmM3TyRbAF5H2O+noqKhn3Tsy6C
65no7C3SSXChNYcJfeUXHXvtGZruSGavvkHtB26e+WGaZ4qsv/TgnbqAWPq/+0NF
ssdGjbLoLlpmw2tfjakHQ8IG0Ajmd+XT1i1UZKATs52xBKd8n3co1xMOFU3Tg/KE
b+LLmfycp/wSsxBJvGGJ5JHbPdyVOFDa3c4jEmXhcJyg5yQXWEAlLdiJJ5CCC/HJ
Oy1PbECzZVeMuukzln25CIrCpIYpLyzjSlJvfOCopvhTIYfW5siN8LptonS0Cebt
6wnc+HfaqvsQJPAPDqEfAnpxsLsHoPm+uKYlrZWFHeSOxbS4PoqpwOVgQBPH1BSg
X41b3oKmiHV8+4abYXdibWub6Q+8lUKRSHucJEZQ0rIE8uTIKdwk9B/o1Pe3DeAo
DDn/W2LZOWC7UMfzt++Xubrtcqs873YRvAzBjPnSdAI14+TAJSz/Hoax6gPBqhQs
l2ly4YM5a9BrC/HbN+aiOjzjnUxKn78MEc4B2SS/RWoEWn+v0A5yZRIVqTOAlzp3
T1IiDN6WxPRERbfiiSbLXuvNEwU5iE/BQh9alZhkAw5UoTWwioRztGfjA/LPw3hq
nOsyJZ88R2Ne6PE0E4MQrHTExwM31Sw3Lv2mqHFomERINZUxL1+Af3PxagbGISpe
d+tuzMn/Pw3GzgnUDEqrjsn8OVMo/ALfYvnDX7My+5aLGywspFR3YZEbr9o5S64G
+wi4XCHTiC7nr7EFweR0v9Bd6oq/8aXxjJvVX5Oiomt1xJhgxh3a78xRZLy8S+v9
h3x00WD+32Yypjg8UBNdlalgq8BCfyDMPQtW1YwcMkeTwAfumINyAXOPVmVg7jiF
Ulu9lZBwTaLSI+4+FBMRPE/yajD6K5r1U52wU4AdtETbrw2ThxBqFkaattdXVVn6
VIezZQMI6Vw/FAcF8o2BWkqcSl3B1RixU7laVMahC55wiCx2SvtALf6fyaB/sNUT
opGwQv4qmbiBhEJADpIp4ttnCkh3Y1y7whiO8lpijRY1h3vRwqFiWmbJQoFRFl7c
dXshMLZCsc4xy7ytkq8tutkSKgP/lDa/rleSxd5iE4sQqM0671MtiNimkHCezOV5
LAzwlFewPCKbUtpz/Vq4C+eXf1i3wdCa/cWa29f+AXdWvSn5Kbwbn3VNnUIHXVi0
nPiDzuEHR+J5c3xbJaIGuW9Obpus5zBW0jUZbm25ChBCknRIGmi7G7wTzdCh56WT
WKcCWuPe82hg4s2Mr3YgkvfqA49UKQoB9njNwzaq5s3orCDZk0P25pprU56HOJF2
hMKeuABeW7paa62msp7+06j4Ti4nERtSmEBv2K4NopE78oPEIeGN1ERiadP1ndbY
lfIRQ83jgd32MeksMo+h5ubZS2v8hXY3JOJdl4AEvTX+v5znBjQWuQ5QuAo57iFM
i64HQ6/N+rcWR2thv6+SsDWgMV3ip4BubdkQNOrJnfGI+mHfhngB1tcxWq6/j9ph
1SbPZC0EYR2o/IiEfeeY4l1VWLpXHjb5up1PaInI4tfBkoCUgtUVuqpncCm69dFd
fT1Efm+siBYRHmQW5TlgVrp9oWQl1cL7ZgMfoeeFy+BZEGZWvMhGqFN3jBkMc4q0
sgZ5b1q0J1tNM+bUnqxna2zgR2V0ACo8I+FC9Q9tUbKlWwwNkMUWL5Eh1IV3G0DK
hGefbu9TSTSEPZPwgG1acpKaODCFTL6onoy8O+zXt0Kzx8EeDgPN6n+vZkJIRaqs
FpRWfbzxFZFcUPPFvj1cYuhjKtSZAYAI9S2pUz3zUukwBCfJTwf72TFGdjzDDT/6
KKQrwnhrXDWavBWc4eKmkYB3GOdm7Tb+grMoMp7MqhwZbd++pWL3iZw8EzrcEZHh
QC0w4jnWZKMG2BeXQFHIkel9Nixs8RzeGlSazHvUKH8eyeeJYcQvz3TdXZKdgjid
bi14VO4JWcgfmF0k4azO+AK/n22Oz9EXhPe2A3EZ/3BM/sFP6Alq7BaQc6GFk6iR
bIVCQcadf4hSP/5NNjnkX7roEnR8UT7P2FLzCOB7L6QyZl95UolVym+SQM6zgh/5
pqNwIy4ph+3XmAOV/fIGb7fgc0nEKlaEPYsDvZgPEaSMPXP9O0o43sxnP8+JJOyu
/TSgmW/T/8N+trNgwxwS5B9+ZhWXbno3r7tu5aprOoRRcMsnPG+QBfA0uMoLQ5h9
2wqVtm+57Resxsuk2qWafsiYezIJJWlLJe0nvkYxKzZ2nEFq8Yi5n8JKBvD/Ut2z
6TpNhcKfQiEETQaADWqWTffB6/EJfQ1004u/ChUoyf7Oc+jXZHHTfPql5/61oQrt
GUG9GS4IDJexPbyVa2CZITkn+1qhszpUTWUYQI3DSZW4b5fAooOct4WbFEskcJg4
535r19IXA4GuSj1gyDaOTIveuDmp9C74GC1m94sjC0RHRIJ5/peqdDO6C8YCb906
BLRtSjw2fOFzr/JQk1WZgXbqVa4xrEf7iWXk6aijE13boguEbRJ5zSzRINIEblHB
PGtqa2BfNyBDdOGK5JrUh3Ukpf9oPqph136IkUKH/hC/lczzODo5oazsRLNY8vJO
2rXG6d2vw9fp/B+sITrIfALarMEemst5180iAttG4hxWijKNRYE8l3RuHelxVf0I
p/CpH8dZY24sntPfI4oLkmMPG01S+UaV/crbheLcPuX0Y+Lx2CifpljkMlk0z1z0
Ujj3g5dg2EqVB0isxvoALh1mnyXDyDwVTC2eLiJrGm331CRrh6vJnYDfCOuaRNAK
+7Ai2u61SvDSrcELntJMHrICKRP5vrk9fG7LwtztpoRRVaB9JXUHfkWo4cbIOUVn
IKYnnpdzOdieJI33re4YQN9rKdwHl7suSWPpLMt5yqsIQoWEDstfC/7fxI4y8OT8
HLDEpeuYfkCS4xyoJFYjTbSrtQnMB361LyaalMlVKm6MsYRbnqaUfvHhwjKKRzUj
4ID3wd23WyqNtlj0YLxydAKOea+K8FoIMOCForC1Dg0kUpRzK1i4FW45pDml8i3e
sy3xMSbloy7VSon5eGpU8mnflwRd2zvPvkdE1VNRrXoHyvstdT+5dTZ38DKCS8Io
qPJpT6NtBaXIS73fs/XQ0w9zuGMN/kZBTeapMcZSink/94dkkUjI5rgxVeR5lwIE
LVQfH7KOxRPeSK2jYOI8o9/m865izdfm7cJK7TSoiH3BNBexN5eummYn8a1t6Bgj
0d3Sb1JNRlla3g4AnYX/G6jn94hi36qSkKQJGPC9T70kX9XvTMjNwm1Y/2QO5c7I
S20GongnEHfT2VYPdOxaxtJb/InNsKSwI4k7T3B6mpOBT7Q1gMrIuUi9SMSN1QXj
jsXY1uhMm47Yg/4Rl4GhcGLEIns2VYwRAxpARquk/ymugMwAPZ1egvXytX5riSY6
l38v4udH509p1OC7VR/ShTNAeonATL8kx2ExNh294wy+cNk9xW4vdUuyyY0ETtJo
XY7rCCy+ZK5jlGJyPAHhD2Xt4UqJbXzR39qFykdBZgrVpW/Okzf0T1ngLKd43pzz
CMD5XVvXEnWIvJioIe5xf7W1iV6OVAldFpaeU+omxNoGfW6HVDv6x0h3P3woUVUK
zs8ixCibpevP7AH9iKVNJVcH5sphQUUjH+SRSLTr9JyF9FmSSjWiwEt/OiUGy2ts
MHWOVCV2/oNfT7QA8Y6FfsV/kKqp5veQmulmyd+7rME0TrL4Z7FSpFEXlIzdQd+F
t6DyVgngG4/JLmlVaDSKn6+xLq97JgkCy6PFreeC7y7jLY5Kihc2/aJIXDE3gGHO
Zi24UBIJDXwH5TU6zinJu4Hhlz3F5h99a3z7GdS23IUFpjUncxNVGL03nggtit+m
wJZ1u21md4TGYDLh+pqeoLWlUX0Jdnr67h8Nz9SXJJnG1N2b6hF/YwQB2MKQEDG8
3AJly/Ur5aGTos8j/uUxIk3oKdzUaFkxcDWZqkP7XNz5ZE4l61rwCPHz9eJP6/5/
UHnkDa59jBZvF53iDb/fxUKH+7kP7stuIL8riN0icHgtit7jWjOuUt8JbjXmKgun
v2hk8cHTVlegSWF4cI4B75bzPT9TXSKAfZOWbTb9IzGwT9MpFG2ed2ov87/2rPUt
zVC691zsVOBfiSwi0MHYcUloaalG24z0wMb5Cwp3nBemh0jJ6lJlE7IvCPZPeYaD
xs0c1WvrwQke2Ki4ajhOHQIS+dh80ozIPFA06Bh0giObPfjB5HwbZLdSmH8QY+L3
xKQvS8BlsQM7leFJ9Oe6ZDDGJig6ft2N00+8KQaS5e4ZnXjONNW5hnEZ+2Y7fbQ+
FKpxGIh3UyQ81J1iLu9IIih/bAL1HpMvsWvcre+1huwrWsVFrz/k1aD5cYu6jmY6
1IicbpYI4ynY2xDzzVBkz9288W26sA3jbncSaRGky46EuhTvRQj1UC4xfN+lb4ws
GsHVQRocdTeqFwToii0HULvy63iixDdWgS7uFDbUU25oYmtIEM4+TvLH+OsdFDb7
xIWFTT4CVmwabXmm4NSLfLqeTYCyG7jJtNHWl6w96wkHYp1AnxmRahC+lowznTx0
ozxxBf7SR+RBrDimxcx8snaOJ73M49Kp+Szwu/vM67vIuu2CAsREZP1r2d8a6jnp
AWwtIVAmBcrLdlQgJJqzP7UnHg9x5Wf0buYuf7odtcjlOdRCjYNfHvVSS4au8MRG
TDs+K68hT9dabc4OLZt/NVlhIt97/VtPvgb6TFEwvDuXcimHA7TOttbILIoH+Ymr
8qg2aXz/03QJpCJ8LJyQK4ymidSghrrqH/bsOsUCdMt9MvoHbOkHtyYdz6PJ3CkH
It0BYE3s1JvmUuQ6ogTdfzI4Ur92HdTUPsT6kN2Ej+3Ha1VoD2U0Hi6VSwtGRnyp
PrS5wBeFkg+Lt6zX/eJ9lFOsu/Hqo1+wOiQ13hRj5g5enirgkoUrdF69WVrxHKNg
I6e7/Y4a9PN4Avl38uayTC51hebngpIRjCnR6n9a5EWR5en/pLxmgpJ2r+dpaXJi
iohKv+FktZQ2NbKsK7B08E7557kHQq2JtkFca/bPwq4TA4s1AneLTVFvaLGquDZF
aiD1EXFL8GWMCIhjxCuA7Oq/lY8Nkio7YCRJXXy5oayWNJFcutmyEig1M5GqhQaf
LKCZcBX1t/CuaVPwmA3pC34TD6kymeRR65RYbXOODmf/m/MQbb2R5IVHt+1/hvno
OY3bkT2j4l9u6apu8NVlj/SZURDDQqMBCbUwh+1JEcPOR5oNOvINTka0uTdq6u5U
IRyhQyTKSrTYJjFpsErTlWuAS88AKZS2ZVpaSf+VOGkX773bAA3VjAKLusaJylM5
LXQoueAvO0QRmland0omCUyAGjBYabNJKwyxuKgqaf5cnKoSlBtXD6Gwt5nYLi98
uCP3oW9aOin+TRc4igtK2DiIH1hzmm/+1QqnydbnyA38t8xpyLbS/c5ZxpZt3vJU
gidAJb0hvyO35fUalBNLXYF9gLoubrH7RlSYz8gRHTV0GvWwKUOET8cl87rcFZwq
kJGjW2uh/1BdWVHm3HE7SGMw3yE4FlCf9qhUE1Bu6rTV0cVRizFPKxCHnOD70w7O
ndo/v+JK2rn95cy1DvXOAn89qiHpgUAUDg2flTzpIrIDUCXZIFbwKkOozN/oJwMA
X3xS1oU4F/b+m58HwWb8LXjcOWNfZISeNKsMZIIlIpS+Ro6SsjBDkSpZ5lf9FsPk
MEbmWsffzWX66sa2QM6oD/WUoSc52JSIZTK+IHj02/bhbznvG7dcPzYf9ZVb87Qm
7PlgcLJ5WibNcn9QuAuFMOHu1wvjEVtANba4mCVycu4UnQ/AvELnkG8rJIJ+v9uq
m1RDXhhksyq1ZMiKBLA3SLSIEMfPaAHeHlUlLMiNcic+xKh9zKNIkRPGd25Wg6FE
0rnYv+RC6enp+OAyODAGQBwrkhIBH6vBZpWtuf5yAlgK8tSi4wwaf8dIjbmyJj9N
zkjMHPLvhSEy3Ks1fqOALof3XchmXAnD35+6rDqTgoWMpoi1zG0GbOyupDyeeO5h
5Biu/caJicx0gftvARmb1eO5gZ6D422cTp2E9/Q+zFQncCBKMpQSda7tGxpm0jsc
7Eaw7YXkKb2iXfRqs0BVieorjx/xhkS9j5tTt8JFoEzPNf0YY2zf4KLValGkChAa
tUyhs3tWPCS87MpknFEdWS/jyDStBApC4R+Fn2bE7OAtXQOT6ud3u3F266DadCDb
SYPM6kYd7I5ygG0M3oTtgLBlTaPDhYqHbkYYJ0opQZq+Xf45TC2ikuhkQ1Bgzecm
eJvImBQ2TM2tSE5pHW0W6Paf8JiTBLe/g/8STWOhcC2B2KxdyKOl14If6uLO1/Vt
5GBpVQsCE1taSLBqqzXhxAd5qqGKsSca+Ik7JmWghjY6VlxGPLzNqOfxwoIj3OuZ
Bnvt8ytTKdGVldXUgkN0tH9Zu2OWiE2rco9uhUiJLckWiYijuA+cNXi79jaQd1Z9
jAqzr+vXjGQ4w9fQqtUjeuaP6IwQEV6PTU8bJSdRo7uIQNZRctBs8o/g4WfoeoJg
WGM0tAIyG0M39cwQhAZmt1x43MbNmwHq/VmE/K5ziGG0ey/QdaWxEJdpJ5169ZXd
O2n06VqtZ8ZDGdThUolooiNUZbMTnrdhA4XmUpCss4z3vl/dXGc2CH3Sl2suIhge
6iEPpsAQ/sk89pNVDT8g4JzpxnAwbJAOZn4aA7Hu48kLSScbPDfNegcRYxSKWZfG
WJpt9mfF43ElRCoIbQTbaeAmyWjkP7g+wQubkb/u0BNYRQp+rbi0DMn/ki+lQCca
IQ52EeQu4lOf0mclw237EcpXe6YON3+SNUYSDVpNNuIThU8fzMlqk5VAXSRmwAib
MbrvAcI5P01gtvTajQq731tfeOmq31BLwSi277xLdfT+MMgVOp1KTOYwyMstaUdG
Kiet1MKK9CFhEBvWqANriUEP3e71FPUCDLklH32oUH4CVzlvx26GA1mBvLWHc+A+
cVoz6YGiYVqLfLE51fSTmnFrYctUcgEU2Y3fWnjoYVcgPxpXi15zo6pkAG4e91KS
ERX24kN/Gq+MxEvQPZEj/gNJoyovGSyaxucI1a1D76kSptpX1uwV9tA8M/BQ8h1x
XLkL6hpYiv8vURva5Q9wT4oC9TmZPK95+F/bahl0PSW29s42lLbpq+NzUBQwUI3w
fz3kBE2W3by7b4+erBJlwj/09nJ+oWd1Z+jzjq+WRryuzzC9j3w9/Wqnqo0hkB6F
xuNCXwRBMrC7ICNMoDOWWVhhuQRY/RKb798dyutX7qOkPccDMyMzBLX2YZ7MtXxX
6t/KwumHL9DPE/c67seInjULD4qo/XSgYfPsLRdkdQ1Bi/JDxKE0LqYJpqAkPqdH
K/fh0UcJQnlzOThM9z6psAoSdQIpQHgvRufbIdhFHm6vmya66ZGnqmN4aiCQMV0x
skk4/QhO5lShsm8kbqtYnU/hY9wwYIxYWUrPcnN/Hys=
`pragma protect end_protected
