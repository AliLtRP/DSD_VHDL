// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:17 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
l84oQL/eq5Nqpy/3odS5NDbMRGVuSksN2pi4VYpVVYS9HKxDuHXQUpqPMcF8V/5d
SCUIO6EVktm3+B5klbHRE5HrplMUIa8e9nZ4nUTK9qGAVks4KMJiX08xIbObXE23
CSK8f3/ge1+Xi4zwz2yNf2Vc+Jr2K9Y1jkP22dp0COs=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 31872)
lHuSa5J9oVvzKMNpJ8zhKoWjtFL/0TTxsaJXlMXCTKueMlYOLmgaZTJuQ4uKZT7t
zNkHFNRx+mNmRqYe/+y4I5UaNrKuF+xvnPly/5Okmvw378g/ySfIvlDkhtEgcc/B
dQhhijR9ueTMVSDiY16Lxq+SgCLielOaa40lZ2yDMCfka1Hspwg5ekK5uyAHPbBL
VE7092uJo0pw8W+qm6Fang3KyKc5agO2Q9YNzfMCbq+SkoZSMlYFvm2svXGZdnJ9
k/3i9ftBiDTfZGYVSMNE9MciCToYSwkrC0+jLrD4KuICJV6SKYa8AC7KKGfrHnl4
mv7zYXv5IpiTTXjhysxT2QS03KZYBNp5EVbfBGtx6K2fT5KbHJtckRh0csxyWRh8
sGt5YXLTtn6A+Upgl3D/ZTGqQEizj2awFWC09EU6s8e5xuyUXC3spuS0sfpD/eMg
kX+PG/x4tmhR7jHemgW8jH8DLoB8HG6dF25EIHsm2stL74KyAYaKk4nzPQCP3ww8
aORZU/7TElS7pqXBaZBbd+cFUgsaZYHkfiil1Idnhg48UG4pl6Og2Bf/kENZDNht
uQFgv43ELz9wcrCd1F4QGG+l1LZHxSi/sH1BDUEf6RHqqB+DkaS0B61FUYlMf9Vv
FtdDZ395glyTvDg4+8jAsxFlNPg5N96lM5+lfFmjXtF/zX+tOrhPEd1ckocZnsRB
kSCaC++tTMIK0uZ5ne0uXdgQOPwB/Sj8uK1KMrtGsXv76Iw1KVir5FglL4mWo7/u
Mf8emN21pqjj7g5ZuEmTNC/RyiN8a+cRLDXSkGR7V50ipV1xDBIAgsZLPVvikVad
DAw94nBeeD0Jnjg7gV5M8IrqEQvqy5EhdkL3n2AnRsmS6FaUoHz8kUhdkhzKnR9D
OEStSesWBi9pHVS+V8D4/0OD8hT4P2KXELSg3B6XpPxC5sf/8lTE2987fnrRvTHf
iFKih6NeOicEEXuPW+6axiQr7Hr6Ygynrq7Y9e6T491DwcxwmDoTkW+8Me2es6m1
1o0rxWcuRT/w05+4+5yEg9e/p0yAwBvaWti6WRWvmhVBD9qEtJViA+eBE8MThB/U
Bs+oSMc/RC7wtxEMeTdZagMKTuMBaBj6msgqys5+HQ/6N4M/6SI0D9P9uq6kQ5HA
gtQW/e3K9kuiYowncgTKsXlufBWosxR8jFudmkuQPDy8mKFTjJ6YChbmjKp1yTcm
Xtc2ew/K2RTVzrVNSeIsbDLHeRQfN2AIORKVmQpZ5vBxaSK2YKAVQK3gNPh+ENYq
S09gQlPld+CWiZaJNEWucgTHL8bgSe1h8cfF1cvR7v3bGbk1j0K67pCDgavpef2L
SBGP7XHYDCn2F6odUrkD1GuUKosJd6hWVFN+XFQ9mO4BDokH9Q3B3XIImsdl1SaP
6Dgt+zuQAhHiZ0MTgvggSjFEXhWHKF7NdA10t/mtVSRfIKy9Lm8QZKeYINGOoLS9
6GBc6KibIu0TivMNthX/kl/JEHy35vqS0XuK7zw7lf0Meqgimj88d7jecvnjHMig
MGO8Bp9HWjz4pfJxhNqoWZhDW9q+zJjYc49+P//TMtSC0x3S8nHfthLuHksQUDo3
H/wMaaExZbWq6rAXdmHa9kXxHBhqZZXCAUeBWTJ5RF461YrR8wPJhgfFJ8WYRDHy
Ori1/e4/U44BNNHclKsMeWUe297NEXYadQF8S6If+RkFweCYlDlF66kX0NE073OC
0R7bijn3YqmTuJFsQyEkp7rIdkpjX9G58TFDENAoJ6FXWCILC3qQqxOyfG7SosAA
oFVmdXh5PeXdF9SP1oY97ywQjYj0TIPf0NIG7UIX8zQJZFMCagqEYP+msW8A3x1Y
4B8+q+c88LEOdYmrKc+AQCBoY2FfQu05r/yHD4HiPODOtodtRqW/vQ83X6ZIKUlJ
O2eSd6/RK6xbixILJkpF5mwoy2Hdg4CuLA5dDJHNLEBiMbuYIiuq72CTsIa72mgp
StGMkFBintmVluI3GzQIEBAep2Ntj+8iV/mAdJ0T9dRsb1Mal2Euo5LvJCRPitI8
xPjf7CVoxJtdPahMkekei3Na1MH7obXU97hrt9kLmSLjA+UP4qJn94qz/wwytv4L
qTNfPMzxAyaYSM3AxW8kkKk+MHhqFvbsJrTP/O1dE1QvdStBVvKpZa/mNDIjvbpD
u+55l6EcCD3eXMblHV0/2FuRoJd9HQPapLY0GN1v1KOvO360k/wffjhRKVLMfHn5
ZxHqXK6RsiX3ZmT8gWWvW4y9eqUh79oRyGpbR4/zG2VTmbN3B899HzjMQg8rkt9U
OrbyMdNONn9jlT7xAqoVZEBxL5aLmGIpym4v4ADI70KXx2Ej6AyIkp8MkWjoAB6t
nv5DYjfa/liodWtW+p+aWnJbYNQ9uAOKFTdwpSX0GqyhU5NqAN513GK0M0retYlU
xHkQntBOBlmf+J85scTpFky0ubuQVwMGuVtMXKLBy6u8UIdw3/oGm8maKJiUYcwh
f9Nuh+jke4Hhy4T1PwpmiJli50mhia/KR4e+A+Hnp/eBi2SnoYdXdbfa4zwfbEgU
5FcrxHlfApdJEExiGeEBts0HcBhlqUvgg/SgK6jG7O6/WeKzqQED8+y4lRDaKHNi
Z9NX1ENFKMklzl7RORCsO3UjFjMMiPQ2KYnV91ONvirFt991wsxDXrw+YQ00/zeA
m/F3oI+tKvS9mftFMCZcaH4aOw8dObY0LpFD1kRlVjBpOvswxgGZsTyNunw5YfzW
VjB+ULJ4VuPf9E1ATTWhFpbOX5woqOXLfSG5AGA6pX/fE04u0L64NGxEC6uIuM1M
pg/PTpYPcOE6WID4xWaTkGT9P7FLM5ZmANCA8zRG7UzAz7gshlP3k3EotYwaGarW
2tWPy4xOmpr9o0oWCPWaWFIN+XCguIqJyffXOvk+bvTQ+weMPXuU7AuVS7spPnga
PSKLhFAwrPt86EVFiC1jFVU4zYcYzatVLy1Y1/EFAkzXUoYkwuy2C7iPPd3aO5mc
qteAod/rTOnC0QiWwoJuX+4qLqam2MpgxcQGCPQ7CtsLi4X+rM1hzTf/379kxr2H
bLXy8eJcHKjn2viRyjJYUn96mRKHPh1VWvfV15IV4POKXGnT1QO5m7ZFKVKFdoPZ
l0PHaUxu++fWh44YIbUrU87vX99vNLLyN8Hu5bv8zQUPc52n/J3mTAGMLMguJnhF
Vsf6r2e8VK0QS1t8NuVnHbHB/ud37/CdLXEoqLGaSTwEKcN3EZ/hdGB7JuSyvDxu
03JYNxULWTMkhH48HpddIECIEPWUEialHJHANlKMI6+F4PEeBYsSd44AvMGoeFO8
5Os9Q11a9rC0hDH6X+yeBzI9CLaUtuuxFNVq2ianYcGj2m1FaIqxGgTMiGTlWQ5L
eJd0ubwM6EdAa5uG4wfpe+tbGuxldT12mUX7bCrn8MUm6ISlh3Ji+Q6Bx/Yys7xq
AsVO0A5BlbZWyOSHW4zfrTHIZD5xTyyJQxgDvqDli8cR6XAD5HCVvVUka2gu40g0
zTGPWQPxUnPvbjsZflgZFoQ4Oqg2NlUl0CCRNzAoJiugfw1a32zy34mpoe3UfBXr
nhQD9RjvMZjUj5eOvna3uzHalNp0e2fY2OS9p7g+coMCnolGfu1ZfLySUC8gMKRB
+FnQXxNHXPSLRmz2uj5obuYv1rMZk5veifgvFOfxWjUUEd0xZc4LcoxYZLQ8CZCt
KOxUmKU1GsK9SLWLY40ult7oQ/iSzlm2C2dJEEyBBN98wFO0i0kO+E8TQP7gKmv3
KZ4i7KbN+LGaQJtfFAYWHbc9/faXUNC21OWfIoVJofXGDrXv8ql1hSjfaNi2VOM3
QIGzp8Ayi0R1znCNjVwo+b6BNKmQD2UTyPQ4b2gmr5PnOxT0vyc6z15BLKfHIRBm
zhSeYtys6zTemxWVidFPKHVJ3/vhlRUktzo+A0v2eeCFqR+P+I/ujcJe8Q5cN1zX
W5WCS2SMUs3rp5yfhn4RdzHkjqL6iFDF3akOUjCp+MTW9Mo+IG/QzWXVTGZaIQ6w
ig/QqSd4CpW7oVlOnILCYgrEY9IxGu2fW9UNf9nRsSbz3NsYfbF8u9O2a4EKuGvM
eQyOWhixC+9umfOSX1pGcZbYzqqUhxKekUfI33HZAa8ZuLy3YwYx2pV2M3lD3iCl
HdRhVeZfrEksC+1/LSdfOR2Z/DtmL02FkqS3MyLSkD87+Te5uoLCyq3vIPJWiQ/a
hgoo1m/peFi1ELsVSgzwj8Bcb7pdSCeWoZJBPOEGkDGpG3X44BGjVUPotm9/m6h8
LPLOBRquL772PMFy4QrA/1Hfu3W9RfdmiG8d81zp5otr1RLNo8cvWpdSiqVZkTZY
lvg5uT9BCIIZVxiwwhqHR0ehcKk0fNQcJUrQlhUK42XqDF9QeUsChfMtHfevu1c7
2p/44LJ7YVxEjy62lRbMQSoXx8jS2V4Ozp7Dltyww29Dg/jyVP5m2jp4liv+N4ji
PhKKsIZkLJZ6kGB8rx8sjE18P5ZuTtbkwJIXtswnlv217Tkg5BcieCMclQj9SBfO
IHz3ivfpDuq1T/0hx5V5Ee6L7ALrRRr1VYj5Hx8lw8pQrH742qtF0PIcN1+rnjSR
zdcClQvdN6qwpvzteKx0nR2p127PN+syP4aiKwXUbO7LyDlAyXU/vHmSbtJcaEif
l8jYx9V4STnWVvIRqi2Jx1I1ahRZMTU/evykyluSrRS1Ze7i1L7Xd+5p7z8GHvCV
4NCXNWwf6vmeyAUzsedwqKzs93ny0v0D7dGP9DE4YFznQ+aRADoxTv6ZSZ4pkds1
V2BV4FRR5gafsuQX6V6NqPCNQ4Ue4Xaz4nhPs+ltiJLyPOOe7+mpqSSyNzZKc/g8
I+hB9PNxmpLR8Oh4zKXneXhiS0dsO6e7UzpXga8zrM9CNfLZ+hDd5fOgImhWGkC7
8Qyow1nenPLn04ftDfpgquLYSN34GAKNT9CN5MV9mhB0VNzngub4c4q1N97n8/bV
suusPELjfulj2a9QJ5Wd/Z8n8tqHPaiexDPPfxpiXUinMJalQcwAmsh+f+nwjsst
p5rwWPX7SgAVQk1gTKSFB9Smopvn8Sh/3L1LA43OkVi6qFrYzIhTNmrS7yC6N8U5
bQPMvm4y1+8qx9S4XFvMTB/wNguY/djzEGxFTgAJNIrksjUbbe1owU5rQRq0BjFh
8H+bXIlJgxsudERSMKe5U6DzOXC6DgYijscPMNso4N8kWFosZ6I99kn9teTPJH67
tZ10otxg4G5D2MK02YhZynYrax8/1FIE6MvFbB+UNZHFM4R+turRh6bffdo8axta
Yd5GocH8/sRDaNOduMVdu8aKgrso5W2Y+UD0YfK0GPMXxbbTTi4geJBve+GrNC3G
PO2y/tSbXv7xxbQBoqkLGRfScjnm8V7He6fVeRxNztCyPI9kJ9IDCl750rJ0yalc
PrTmhpqPC6TSj2XBlpxh0Ifb12OwR4kleWomA09DYAGH3FhTBHVCW8CNxcmStaRj
9J6k8Oovkm1wrzt9d/NYlISml+pphwV4dym4jZGm0tZ+ufmwKUaJCVMpA5Oj/Ycs
7dKhU+78PTYTZyq2cb2bYj9oJ57ZuPQrx4ooSow/pAmG4Ib7ImC56+UrOrIX0M3z
9IIa6xzD8OkVq99Pf/YDaIQ5JVv1us2NYAM4NlJb9bPeAfm81Gq1tTvWXanzMAM+
BkekjhNfzhg0LLa1zJodFim4HvdC+uMpiC+7JHCmgV4BHE8SWcFGLEgBaWjRdIoH
hxHw+6VjgFZaHJ6hQ++HnModcnHuRtkUHIaf4A0FvSXFGzxbE4k/5xMmhjhUXt/J
pmkJLxEoV3UeZPB9Ynl5JO6UjuhTMS857HpebNRWGcd4IyxkssteKbuiFUreRruc
nM8zZBdcFAJ4Y9SkK39Mho6xlvS9wFMTlxLfV5FLZ68HOGZ/1izdAVk6VoClgENz
FW+BfJysyerEvx1oQMxCPaiy61yoiT1iGF+/rCjZVv+MUeTiE/hgd50xEqzq1IQ2
LRrjeL2kNcScFZ9i9Iacyt3FnFwuoOcYC0SKIB+fc0HhGJ/SKwWNVvgpAKnntF3T
G01oExyFN2ZV+dSWWJtPCVraCChaCXoUciYwmE5Pb9rdS2UPlrPeQRAvLw0QPEVH
/Mcwbc8RDd4fWWx8Vuqu6nozOyDPRObZxSaDnmFZBRwcA2LxDH+0Kpi1DmMbATza
znJ+BDl+KOONwfOU6SQK1k++WHKZDFciH5Z5TfFHq9AB5dr3VdqglfgSzWwcrA0B
EzK+cN+60Ec2U/zKKa3hCWd5VRB9O7CLL4V6P23c+JV5EEranx2jGPPL0T7gCWEa
g8Az94wkaW5FEAb3Qu8e1Cxzy4wkh+mM5TZoMhn9W+F/usJtJVhXCIAAvanedHah
S/wlenZuiEhvLfBYFRs5BL2bXdq1XhLIzHlQ67bgJ3oWy89rNrKj9D56F3D5v8n2
nxOquoFZFUCRYS3sjlSsRmEaxhEZ22eYaLf3v1I/F0yDkvYkqPKzyd59rj4kBIWj
pTW/xio2kBUjJ8rbcglLkNFU6v4+dZbEIewjEUkHujm5sd6B6kgRBrdCHOxgWt/G
9VOlgJo09xMrkmmoQIz3k1X/2W3y1NN2P02jyPTmskvfWxe6xNUZC383KFdfUyTw
XD30a6uMBzOLynmcRyg+js80bNmUZwZ1jAR1RklsrCMdH68SwowedOjCS13kjqJT
pSYwuSj/sVt8k0MENlyjo7IO45yoyZtWWPg/lbdZp7mywti0aVfLcDbVOma9C/hu
PFJk5xdzj1xdguiSr7EZqIJut4/eeHy4eqEweeEppqsEZWN7IKYQRQ/N0okcQIbH
6e3i+tquSqcAcvZ+D48saukyywTIxQejVvsWJ3JJdGPifS4wdd6ZY4Sr1JmEM1i+
k7dZE5dYgnDJ25RqMPkSe0FNuthopYdL8SHEnZn+muzR7nW+hdzXFB5rGNZpedlJ
3U0OCRF4IAbcHPzvKhJWFkHkZ4qPlDh61ZKcmGbUa9LVOYDbcY3WkwiAn4Ol4R5v
pevX3GGCbqMOjwOdI36Fk2l9Lh16VZCfoA+fv+mf/sC0X+Rjg8+VEz8v9NUiU2Ku
PoLvaV6s6LAnNJIYwk1sWmJ8EsIhdjJMrO9S8FAqg2QUyEz6Az3f/yeykgPgenZs
jFXQsO9aksklZZs/4BCLBoIJkWxU0fmfwMhHIpyNF9NOsBNwQbp3VkpawuTmNdpf
GIKtqUwF112RoEL6DBpULeXocaJuoEw6tk9OOR0EPCBrpIQjtQtT2QorRlMndIas
wIlAMrz62IXAm6Ch8QHlW/9LiMQNOC1o6xDZ6kJjVSp06KQWtt2swuPzM+FQDeEa
lIFi2tZSXdoex7e9pMRiWJ+Z86EYgl8wmuC0zKgap6fxL7X/KHWIQGhvjiZP3Uze
zjRUGhhMHeT/qkgcSezQDOYOI360Wrg8NNaGNrlh0zIyC9eBSuapD2Y+nOi5gBEd
PFGz/9bMixyh0BrQCzr6g2B+rQokkK+C/2HaeytMilCpJWjytB6Y2k/GsKb7m6gt
iGzg1B31GB8KmUpWszBPjouuVXT6jBDsRnZz07z7sIPsbeXX5bsBStkOtAlmZ+ez
EKk/AmRgWOKnmnvJQhbWyiHxY4ghO7YyRne3ZnabjwlPAfRLN37v+2Z8xpfL5QzW
BpAt27hfPUNN01Ek6i0xK+X80atXSxTqT4rZsvfQV/48fqvg48/kGyngsgTGmFPW
td0byIgnXOXiDYDLY+pGQnvVefKxUPrFPJ3k1J6xK/0lOgbgfzv1MV9+f2DDuoHW
b8owm9Ey2ZvSYsPwXL5ZM2KiQypga08mhjcuUM1LWjjhvuTg7ddYqVGuRrnlXVjd
LmP5pYjZUAM2fCStWWaN+FJ34OxbPiTH1uPv2oPjVvgw+xWPSlF/J3tBdjlP/J8c
wK1wN17KT/+ehOc4wcEXBEH+IPPhNvLfHEcB8Cuisw817gXCxRbMDgZ1uzLIA/SO
s2NdMoNMhH1V7p1nPOVGLJLtPv7XnqPZGvnC6lUvlHY2Yj5h9s7qkfWuo+6r5tI3
rubSifKkNU7NL1zanxp7Mn18ynX8kxeTWOIepuVDzUEhVqWP1AjogS3HhuK04YWE
9o8xY2LG4ds9ToDWztYFYb4BMxOfKQcQIwoKRNGKGPSmeLlQ29tQHL3jbbZchEDR
0DE9GpPly8mLUxR+3XR/MRpQuRYl2v/kAllO9SaNvwlDyO5eomaoYaEHl+QQ8X72
U2heJXBjgmY2AY3Zwvm035m/Z70A9S72Z73oCRhaRR3f62bCawjv41zsT3+RINf6
8Z0TwLubCtUefGdHUs3csVCFFfqbka6pqZ6kP9X4UrQGh9mVdj3c6NJ4DU2uwatz
slVdrivp6hBT0kjKJpSCut0wO7xfZGW9eqdwiZR+gJNdPgnI2/7JBNyGSBnQcK4t
2hWfSiNm7AR7ZUUfVVvYm1ZacsexSfFY8mcAZpjAcd+Htyc+6oj1+0wJSZsFlHOe
q7cqzIWcRtKfHh8ZpOWR7j87nb5fQBH+K6+LpYxp4GhBnxptdegNaYHwWJQDawua
M7DXjsu9YSNpICOI+JBwr7TL6EiHNTzb+lXGc/nRsPzG+Z+9e+uAgvq/TSPyV6iZ
SgOyOuDv1CWRmEFYIFqCRbL7Nblv0+Qf6C50gkJ2rUcl87n6rb+rcnXP9eElZVnC
BiSlujAheU/Z6Qf0xsMP9S0XCKE2IZYNQ745kSZoSLBJ9mMuH+U2Zgt15uj0vO4b
i7K4QxlwQj+rFvHV9PeCqEbvhvurOLwO1LhXehNFVLtHcCx268w9pqAxPwdw5NOR
brb+MAqqSKX0FMkhsPU92l0qksgvh9XwlszYYVt5NsvAmPZ2NXSlIcr4UPss2rxI
dboz3Jd2a6/56JwQ+Of/gXA/OpEdH4wyJuP9ux7q0SeMLT4hBLJLSejrnqxxIs/j
XQtzBMNRYbmjb2dLoRQI1J/XDSGDxhNsRCOkno45Wnh1JWd2GFcoxhXfTypY/nlK
Z9fMLM6lyXJxVB7O+naGJ3nbqM4m0dBPA3/nEd70orJOWt05OmgIUJs2r6llTDuT
LRo/uC4RVsNbcEb4KL2nnqEdL+KmgAiGV79Z4B3THN90IdFGAlhLCuV8rIBSKBft
eResOLsMkxHDi1wztwnNfodrPUmzOPYN+CXpGLvSD0dUN9MAgnhnZ03yaResLEKC
2lPmOtjEVPXwfwKj11jfaM4uWzYIzyP09auOwgRbA53Zvb6CoWraKpvQsGYcKHO5
Iih8hmVyDppqhBYbSNXbsPlsf7CTI+F3aEQUW97wGNkF+qu96o26MZ0cfLPJ8Mo/
aDOWyLrehlnOSmMiWsR5PxolsyoPhfxUikJ9EKM0Fo+PVuzfgwkzNjCskojYVvIJ
TTSTJCLUb/8M0Hyu792XK7EfuWfuWW8vH8G0NZBzFKR1Plv5Ncjhx+ozpCUwQs17
UHXYWEr6Cdm6mK05VQNQIMzmtgLUsHzdsjDUn+9mC9+CFu4uVMr6HvPRTzvKBwFQ
OEgHZ/qmXalI7uvNp+U5ZK+jliE3xWioP7p5lyiS79SnmAq/7xRFi/ll/rIqpwl5
WGYPqLya1Fc7bRAsw9XwoCS84SR6oycmRr3VhxogeW9BVCvg7FuUm5u+P+/psJEo
PPnCLkrMmYX1+b+J7yVOBMrRuUO5rgMaxnG0XKdgxVG09HAA73sLCeHFbObXQPLH
cc84dFJlqoZAh1tgSphN4Rtddzs4Uno7wOTWT64Cy4/9XJQoryiYkhWct4rSRKkU
uWfTzzLfMPzu/mQEAuO9RgTj2R1cY3ps8Y4/imAs+LwifqxcTGmvtH2onl3N+IQL
bK4XyUSCuwjCZ2n39H9SKmbavKSdHk+I6tODsFKSf3ZRaTWVRfT72ZpzIenxQbDt
1nAXRZIRZib1jj8H/DQphAKM8sgYTnAdDNTC0dgyK+aRE8bBJFkJC/1jUCS3/Ksx
PTnaHxaYobgeMRl3dF3lDCAi8Mj6mEYLkGM+1bR58xjF5ogNxFJEKt5giscE7hEp
4SfthOWrZNJhhtEJkGqI+z815GhvoVqVFEHNHqg7TENhbQPHKpPnMm+1r41KQehn
pXL6P5EJ3RHbnWw+ZlVY1qCc5s21os+SXVNZvMHxtMeivSN7Tovc8wh84WO5PUlW
6rsab4TD9MzE7DM9FUAVjMlt7AbR2aulCr9fzBDqqAopFllkcn3rn0GcmdT8wsFW
s+ZeHuazse+6+4S5JL3SdIdheBKxSVi4Qe3VgPuRyPMkmO3d1atqAVYqRAcgaZsI
Ii603GizmApG2FuC/XR4lOFNKXuYPNBnntoaA455GTYO5H+i9yYUqGF0I4QWKcfR
aO191HEGfCzIY2zOLx3ELR3VZEK8zEK7kavC+wo4GF3hzHYkNx5fQu24nNQzZfjB
0xVC4nhmAYLnFTPx1WWMuK+jZS3nGp18tW50OYFVq+tAwsrfo34Ru8tS3zwjSqGL
D9xPaG4m/C7t/AocBmxFPnt6cZtCarZJRoHNblbWVScxfldGb5nGy+ezvCS5byC4
rPFEjPotIR469/rHGUTZLm9Tq7SvgerAjgQItQf0BBMk0uHn+LyxIc0oySgU1rXq
LcRf0tWLgv2JxFgVQ3UHFhkWIeJ2ZDvmmDc5S3hofFqf+aS3cDZfkXyu8wWXy65S
iJm3WMqhnUAbj4oaUjihSP+XpvNNC+48S3nNZL9gSxPAomI/x7yvYV2/+eTDG29K
NAsl37GQUI/iqM3AEuq5q1vgTyJu3Vh7gZxxHUY0RpdkuxxNxXU4a94UrWvYhWF8
MKBKuiKWxIkotatI+QLLN4iFlbw3M2h9ggRa5fgV3RZqzWk3m5h6UB1BdgckcjZ1
FLw48XUUmwEwkewzbBiRtjtxOAwXMOPejRgy024hVvNTv2pl9Gjvuo4OPPtdlEEt
EciLCKd3g7UQjHx/gt0fQUs3BJh3YvKEG+cGXVVt00mTZ1eO3X/ARiieWStkvcao
HiZ2usKWUzDq9AdhSIrEDyZMdKVva+5d3L7jGQxCQeiS3YW6+cGFaHwhUWNLIKY9
o6pa+8qjaPVtV4Eg+Afy6xvHKPPaw/R6BSCoAydj/vUmKOHyzVazmXt2YHoZ+cXC
RtazH0HQ3M9viRf94HaU1JWkJQGOS1LPq0zfdpqOKQUPBqLw8P0ZV+O3e+h5BVC2
43Sz3FRWUNKNzVJdslv863EpgPhhhstAHjgMapQD6F4lN0ShPuGqpgC24kfyAMMm
dc0ZS+CCD4yS75jK9sOc3NvR2T+Rtze7C1K7QYBNhUdykBQ5Eg8JDhKudGTGjEQD
nycsOjkFvzSd5CPvreZpykSLv8WRN5wJaS4ZeMXNhGCfLtbIOoRSzWODAaE0790R
nx+/pfK6dU0cbTwodR13L6TA4OZmy5NjJalJCONo3G02BIVT3LHQlgGgtKM0wH7n
3ABtwj4m+yUGYmx1yEV4ZHQpPo402woddDNbWYOtl3dp+oDcR5ejfr0KW1lZ+8YH
8nTRFwtgqLJJwRkh8MUDntGbDuMTYuKOOoAis9+R3GYfQuWYF81DMR43KyFsrSeX
gTOR8W+/SA9ZVX6w0FwQOjobvZhgLIkqF/n82OhlrywEme7urefIMK7ZsW+MprpM
dTqBdHqk83QLZkpg4MNxsJoblxn3+ylam9He7l5KUn+gqtbgvRwbSKAp5tdT6SQA
+cV93Nf0qky8WM/3iV7fRtyPG8wr2AMrjZCwWeG74Ltk/1OBtW3aJ6PSXFJ2Sypb
sj3Wqaaaj0wdPMbfnKS6OhRMaI45lr9iS39gW+DEHcYFBpJJVPh6vCzJyTROgo0W
LeLib9t04ZuNvo/xlk8Lu3ZPJJsK/SqlYSENlGcT1gg7IghVz5mBl8o/NFykGj7Z
2GPq8KRwR6G9+vtV4enlD1N9yEfZpfm2H3SAxepP0mBk/nI8Q1NZTTHeDhxpmZmw
Q9pKz+cUomYL4n73B281wvxOFmLoYN/8mQjoX+hnbyhzmR6trNFJhDx/LRQJsji8
UBUDLk1u484ozBDixoFQ4afRAUx+3U6I1ddRpsCkU3z0WqB9mAUA4jkklk1bstZW
K8ksOfdh36H5F5Vx/9xr4S6hQUwUA37CJyboZOMmwY+FtB2UmxGEQl06eB3Zqaer
CpI+C9Il2aob2cYGe9bwqQkQ51H15pRvIE7I1dJDtaQp3ylFVh69mT/13n64VY+r
7qRS+wKFgpmXr9wwP1neySE5kTC8Nmonc+iEJqhpjaLsV74F46FQ20a13aXQQ5zu
5ptBt4zu77yOM+dyKWfMYWBuCgEbLFjRI3692h/NSOYlgKYZOOJRLxmO91b5O5Ai
kt01uH355fHZjww+h2FAZHjbJSvvoctVmpMOsAOSo8uMwXDjvOT+3TFvaHFAkiiC
u0TFgF+hNKJyAbbRV8o3+eMc0Bl1h9tMnVWXOUbrzTfUux5Spoy0ys/O3XqdhXOQ
j9zzyFUq40oXhrhwlXuNhtFgdvpqHM7z4xXmiceSX6Zcfe/AcOWUOJQX2ugWXGlJ
c95qeY7k9gU89vbbU9X1lFjrGhrlamEGzJk3emFuwBcT/Bam8Y+SfLoYUibBCzfR
9B+4ztGqKZgdOkZ5AAgnwAZ3Rs/naQdS6xZCvoCkAy9ZsF4CjbVx2q4mI6IwIF7n
cXWxPQgnC//HZLkspoLbiBmtjhzsry1h2PYts4Hk02gJU1RsqLfzeIiZFimBBQLI
OHk6sQzVWk3gYabnWp4L8EiGbVKbi8ovRlWgzit72IuT5VkVrfSo8cN5DQGbsER/
XUBhUwBM+mu/jjXi6pt2ap47bnG/fSdPTjd9N/IQc5x6CBqlUhPH4NX7tbWQqoKA
AkK8S1r4UJndYhcRr577LrSqzo5nx9sfx6LPIRKLGBEXIK6PA5STFxng9Ng3uZWb
TZ8cu0nBx60YX6FnLDn4erlP3lfrU3s373SdfHzlM8RAKKvSdq59QroiSUsIx16g
FfTb6DaSsUfdLQ8H5wPbjjBfozn9lZzV+xF646QJUgGR0z5OmiDxj0idZGvsArhX
EDlV4TfKvupFhNX+hPW0AuOuP32oZ56FQtnlcBKk8LnUFsFWqckUR0NtuZuA3+xJ
3t7E5t8P07miA9ulUbUq31MhJRD16K1slY1hF3ZeWdVOqhEMa/PfMeuUwJq4NQpR
LMHWMirERZJV1F60r4mAURmJ/yVaOMZPDkFVJf0Fvp6FGbX9zI35zduclMgqUAZZ
6LOEJDXu54v+ZlXZ3lht+XN3d69LDhFp8hzL7/RC/fPsKo5jkuOQZXx0KOPKb4fK
7mzeVdGn/FPhd+Ng+S6oWD0LASp0UeXCAXJySFSiuUtjlc9QtuchgAZ/CszbyerZ
pTRHABokkFw4teWNbDEkGpr3RYn92dIAKD0f64dpy0fbbGaHqRGEaZA8NfS+zDvF
kvCYzrZD8jBCuBp1lQpq6X4i0S5mxn/mJpNE/zThdCUADATv5VPSZmMSTASTlGEm
otHMrZ5k9q8XOwYg6+PI10728LCBRqHkqhG8Pe62DWYZ3o1z6TfcTwkz09CjMZGY
ey8hPU+1a6hK28W73fmkNlGzoQQI3oQxZwxku21L470TMF+cpghzU7u2S7V6L5PL
yB+P09gUQJYQhnEdtwlw0z3dKqG2O1esLOYVb2GDDxJOFmh2Q3ahLYAG9MAKDyR1
9LTHRzpxGbxJpUJqbvZMMTj4/hS8eCHAGUwkYzgp7EMYx+dMVYUMx/MId8TSf/SO
1Y0sQUL4i/85qwEBLV6W6YEAKe2VgEXizshun8u4fXAXqN7GYjkC12etKN8bOQWz
Mqm+XvHuYeiw2oXDsm5gGuC56yRphB/CUn1Nuoki5TnyV2Gm7L5fzIR/NAJnj8Cf
IaSDqG4Ah7g4iJfyuHjDPmyGEGT02PTGba5FQ6nDoKNW5nZEvIEzRd+06Yv585xV
ssVx1TxCqa4iUEy+RsVLp3X5pl3vkcmGMWGPBUAYXmSxqfvCncwITJ+1JSQuBraK
JB8GhYwJu+F1JUdXzqQKC5ZSJBHcyyErUzi7dglycVcY0ngg7vmCBix2cQhV6HOM
a4/XZXOOu3OOGHEZB4saq3PAssjSb28fDfH+W/Eh2N/VU8JJCTnWfxB6YN8eu7w9
xYM65p0ERqIj1890mfQ499fmVABq6ABDaElp8CkT7EjT1rjZRZl/ZXrzGkA7lBaH
Tt4XWT+epJ31BnY7gzUdzRmUTFkNGRxFiPRzZQ4vz7ZWm98YbJOdkgZ/9duFrKzQ
y38e8joOlmBIH48QUG/AT6JthvRDLUTGDpW0sWDo2qVaMAKQFjvg8gRjwrcnVz6j
UX60cdUWKrjc0CZDleYzdeIRBeXJOGUBMJDQhffQd/k48dCVnUDl+QzsoixVoFBg
LJXDJlqvMrqyHdWKSybvvrT9xUlhhtm/uATg+9LR3VIvTxYgGWJSz3kI2Lg6CUOH
XeciXBMI0Uuz0VeCSVkl+qBg+hgRt+gVZ+h2pXxA49gSilry3PY7Ex5JRt7U0x5r
ILB0lC3Sjr7F2qQ5OcM6qPYjLDtSZEM3rL3c+esAutpAUiDhFmD6IJWpiikvVFtW
Pcm4mqU1dvIJIbWSToWYELFdHnuE7UeEmRJDyYAd1TTBRRu0z7m5921PMbB+bMlp
E3mYHeKHLdJkYGEgadnjM/+BztrUHf5goECOT01Tz8w/U+3VLg9CSghwvrdRwiTc
nkPBcLJO/1Oy7ll06ebOZMHLpJD8zOWHPtJrT3c5KvrqoU/AAMeGKsdPHSPS1PYG
jwjcrpbShQ3mddZBdcSSSMx1/hhffI+GrA4Q8p46WgUngI+trK3KABDGBun/gOlv
6N/75/F/8fLZI/lPod9O6lUDv2fRP8BPY7NpakqPm7oAq4Fd7uUppDkLfXFi/JlT
ozCXyfOMt3zvBSr1W21IduLgEk6ME3Gr9Hd1la3X0ZzNiRrgA6o2zMxkwJRuoEOv
ixGlEBeyDyib8xTonF8HJT2e00E3Mo2czQ/cP7wyJLWsuVNJkanR/UF7UQj3HXvV
MJAZLumUbn8T3MlsjmNraTfnUOEYGjuL3uHmydHB0U2qKgiPNDt0fkWgsNb9z7vR
pisLY4tls2PljwBHnPfm4lGYl0N/nTgr5s3O1qSvKPkl1o3+1ofBSd9MUvkXppy6
UbBdwtnlj/6V3WLrUdIP6Ha5D/PGVHFzmz5PAHJnLTkfvZgxM5d6TuuTzDUhB1IV
8LCKZm276dGHpNnCSSds3fGJm+52XuH2X/W8YXAZLvHdsJfyWZ+Qb6PHXNhCRxIM
4pKqiZbv85LZwW8oBaQouBjkzCAKKqK8+79dZU4VWXXMnrJPxvDG0i4usj64lftF
l8r2jHcHd9k1i38SAa6m2d3WVDxUXHdBNALOpLOXenHg2hl9y8SmAl8Iys/kHRSi
LjIN9n8tjXvGhX5M2CVpzYgGx9txcJJIiQ7GzN2KMoQgulpysKwPLxW7m7UJYdCn
6Mh0SB998tg/SWcv8HM9fON2tbWjZXS/yPlr6RRz5hKl6pjww6WcpnbfeBS3FQz0
fbcg49n0ZvQO/9IDhuuClOy0juBlHGgTBSDV369yLf/wEKUyXAPBHNvkHOysMa7Q
rr+B7bzlMBRgkWyM/wEttTBSPb95aZt6r5FdxmV29HS2B/V5uYbU/u9GrtGcL3Ob
2P0inSz73RLAuXaYvAdkHtfZuq3eu894qI6L35EK318iEBtOwtOxtJ9PqlDnaehD
zLjt8Bl3JFI0Ea5sfuSrDKBKhFS985NTBeomyVLv5Z4TafcJeHwzc+x/LyEQIyaV
78TdiJIwoNVucUApjskQE/U5ZG3vVbWESWu4iZRyou2Q95qmN6mCP4+6N4apNz17
eBfa4njZlARqgMbhY1iGroq8057gFiv4nZugn39tfSBP9Y4+8s9G6odLbREFcyXh
6tf1W5UsylF3dsz229lcPdMY1cb5mEMCken1hRlI3Zz41nNAoSWvaG5TCN9oLC/I
5TrCUJEffGipwaU//Doo3augiMRI1ufOZybKnvg1Mx5aJYKz41SMAWdVjvqvKzJi
pQXt4MLcWPxnxEfR2CY/SEELfFJWaC0ny8oz64ITW45IAG6wM95rPFD9cLvG1FLD
4q1REOLSBrkqAQdYq2bd3qosvq2KkEkRHpjXHe2udB9WKDP8gZ8iZehWA+PABRpm
XJd33BBVuARu9mjFVq/CD7j7R2wFq9lBPlDi2oytkcH6qCPzuA07JB4vuYk/xWd6
4s+3TwYNVoYRWCZN/EqfQFT8hIRcGgOkQRdeSrcw7RXrvCC4t8pNEkeUhRH5NMyd
4o6ag95xZySkb+GJy5oPeGDrIHUeP32z7OCKmgcoNkAjCLEB9z79VaGZqUIa95kj
WoTvCnKBht7glRqJzi7WZZyMgYpUSFL+EGdMO6HSP2wlcN2M/6B2v+0wurJcHFCR
LOCwGGRllH1r1NIJUs9qRksr2zFUQFLTjZFcX4gDF6amp5+Wirs4cCeUD33kySkQ
KAQopg2NJM3NgdzTzcnpIv7APiCa+UnXZKCW3N8R6sWJv6io0p+gMc3lBB9WNnXe
Pr/PqpRjFoPwwXeUsssfyYRwkBLfdqUGtmms2sFc7fz9++hxVJQTTzAQwAKVCw7w
2yuhCrPke6IlwZ/dR9h4EjEZxwCNqnh8VnwQtl+7IZWLmfAQU5LqCXkErAC83nXe
oxdebqG8gytVY0Kdbk6C7K83qpl57LOCVsTbYhE0DZsRRHnIKbwahQKL9goBJhqL
J7tX51nJa8wX2vfjQnS5PkUy0zhgdT276YZF79u3LhAieJwhlGJDY/A46pcZFOXq
H+u10t01aBUBXU2dWW1qcKv9UCSYnTEkv5V8/+e2THZaDKZbeUGhAKQkuRNl4F7e
XueeD7PQhjkBuygycrX7DjIr8x43b/jQGcQ6B6C6zcNZQ4Rqch+MBW6P6ag/iXwy
XFfKRL72cPRDXDb9U+0fBOFZijU2W6NAJ8bZPAEL7yBMkEWv44SbUhxyImHc9FBP
aQTPDAMrbk+cY6lA0je1W0ur9amGynxXvr0f0CgXedC9b0zEJ3uq7f6wQTSC35E4
7N9klkyaJ+y0yVpi7iON8qTePRKSAmx7auMDg3nBlhkZYxCYwQ+nFTlgJGLaKmAV
HaJPILOewh8Eph3FvVEralhvAnPJL0zNG7DsAVjp2kyn52/FtkpRH3dg/tOmOnqX
8atTzhc2FcPf+g4Zv2yHzIM/vhBdxU2QC51SCvFy8yEqUqTFTv/uJ/WGFUZ696hd
MEHcket/e2SeO2WlJ9j97dzmVvGx7Elowgrf7cSxae/c5ewiu514ctTAZ8Ezvqsd
y+B+2h6Y7Dfa+NVMxUhYsiTV9GheV6HjTHeBAlDIuOG5UE++fi0rcKUh+8NmbRJN
MhEs+33XnSqNXlt178AiP/Oynxy1w7lWV5gdwbN1C+QZ59/Jz6I5me6O/IkkrFso
HHdWqUB0MVNff+ADS8mziREj5/rzDwAK0c5anjEeqWpKF08mfc5xf6bU03wy/A8Z
EEijKaOMqP86L5B/rP4badfPXMigFXOE1VqF5HXwx4KzV3Ee/wqUnhTHFSiuQa6u
jGQlFc1SRjIeoEqLnwI2Pph/8yXEsdJBBKxOux9dG3TCBY1HYA0dATdCDBXDu1MZ
fEswAcSyrXY4STs4YfmImv+PqfZddgGHtDNTxAom89N7lcRj8YOjYHL8uVSDQhNE
OVXbjayVEHloSTNX2a4s7/a7TFUO1GXpzYt2sRV8ZA+hMI0bWielAwG2BK6snBgt
VZ0wlHR2GZtNT6VDFOxRzXcSl8QWz8abCsol/GV75YUq56x2IXJSL7N2/Zm5mX8a
WUN0Be9MGh6Ybakuf9lPn5NVjXyNsUsILdxorWJif6WXExv4zMvxqdVzx6wF4a2c
KYKyYIJyAb5/7QvRFynHfMbBYcas6indhC8vI60uh9bqRu3SMmz7ujp7XmKuXekB
/0N9y09EGgVWiaG3zFvS5UaYCBDBIcsEq0d3dK+ZoP5N+KEl9fwCkLfx19WyZsLJ
O7d/RVVKSX1Rf/j1PKpn+VJ166EiBU0ggHk7VHyaSbwH5ouAyyfQn9vylm0cf59F
eMb4VMOBxA0ZC0GZ+dDOvi+zoG0RnNd+e8em1GqKwekCPIWeBqiheh4A42qSCk0u
jjsjd5XsqzvK/XrwnpbheGgV8B+8wmJwmj6yJkP13IzAXz9l8NFX8aR2VhRKuvmQ
GZXyvqQY4ogshJwYMxaf+G9VVNKoyHKPrD5uhfbmBgdbM2+hzloML7awdh8MG2PC
Snt/JqXu975GEkQg6eHLtTHuzijGmJviVPHFgle4mk2F661qh3Cdyp5AxI8KliwW
EKve595qEXvkSpZvK6cvivVxS73P84gXl4C4TzwJLvUmTD6edPfbYdCECvH9uVaw
mej2JwwtNqPT+GlJhep5cualJDQItg/AswUjTIJr+yPzhsfBpdWMIYu1WbCp1oVt
RhYpvK7zGZeMQkunokenAQa1PE4rfaT2/fDenGz6YfLm+HZxqcvqx2ypkBlhTg9Y
YpDTFaVbjoUf2lQrnE9a50/0E11giEZ1blWG418WfEfPoNlba0/7uyTlfXkBwQRo
jiG7zKVz3rmaCkcYxKu4MW/nTdyB+A8Q2IEb1JbSEZGs2mWKwRwVWUon8kuWmsId
rxHaZ0GgMUCmBowPRMNsYFcMylRL7eHcPFxysiWvzqdynDk7H4qtR+x/kWk47y3b
+5ke6M0dERBzRI6Fx1ncSMt3Ccl7rrCMZXy+ln2vpyhvfiUhhDUxjpVgYn94ZFIa
TXlkaLPicLbULrheJRLHTeEJ8O/ZVCdKWknQ0YhcWAgqvZ7FrOxLqHHKFkBrxXRY
77PlfMML72mwQDpaHQ3gqjy16cGX3HKpFey8b9IQGNLn4Q1Ib7z7mKOBRGg2fVN+
hccQZS7+XsmuH3Kvo+OHXvjd4Uy5A+MoYNGVAPoMl9ZO2tRLYM6q5t/9MXrLnSKN
auj3HYDFm7hK+tlA0GDP09bcESgYPft7UIOdCai5sDTL1vffbQVnRV7IujqOlR4m
Ptr4/62sY0nkQ+deCJEbwu1hFx8v/xEsxRTkqbcCjj4ghYV25ro9O3zzFPvfgJn5
0hD10v6b04EVJaEafWtUMQeQHHCwq/AEkQlpg2B++WQfhLc2XDgG/bOCMuI4zgNB
/OJnc4krdclK3be/Z5u66PwOSxmg3PW6nEKgAvi7zkRsbfJro4Y46UebJK79+h/5
ZUiC9U9zYUeyT2nFQul/VPSbSMhL5B7xSgeSLmhCO1dDP4w68P6K0Pmu6AypTBHx
kiOTYWocNsgZalUWPp+oerwsLNzKjm2z3Ausc0MDIbO77iz7Uxxhu00MmT1U2PPt
YHsiGTVoHHeP6qRG9icb0oautc9yaKwm97wf4DRf4A7I/zZnoRZPzTmQaL4X2NHU
pDgZupfFdllXRWsi/16C7ErJXHo61K6s5CgaUQvwK0I8SsVxEuTnudQ8Xs315kgk
0L8DnKenuSzCr6SUw4r4+8cu8BhvYXkF+KqONVkMQWgXwkLqwKW/hO/QVKuHr7GZ
9fUFRvzEb/mb+fD/maExMZuDKtjMz5PPH8NCoAfZw9jTg9swSYeK1pHIJqqJzhOt
7HMb4+UATbdNtNJnUagPpQvisDZuPNlVN/p0J0fhf7KEVX7+eggUE/CnCIfhiIMT
DeAgBhI3Em0STteBAHfrr531q2RusQjPP8t0wWivwW9n9E8jfalS4+o05Tr6HNO7
O3nJIH3HyB0Dj8e82wrBsn+sXpY7lKfH8ZfBnG414IYLBKw3ya94xLKJTPfDvEOU
9RfqrpUyuDjCuvJbTrn5nBAIoP4wErTXelEQP6NlMM2vt1XVXdT7QZCNP6dTo+rM
Y7vbOlssBWyIiO+SY6z7be3lCtIf611GxTS5ZrGDAIMs4z1nyi0dCh7BN6QZtXb9
l5E4tkM0AfR2ImOjs7FGK4NAxyKGHloLzho68b4s6+WlswgdcWP3guA3sodGbF1R
KH58F4It+ADg8k2nxiAa8VU4xwtX0V/InNOCZV0eI+d9mFfw5okKg4q0xceTLSK4
3OZoVMPWNEc8bWWWZ7L+WFd18R6xTjbSAc6TwuusUmhyhqG6PkGXMFpPtm8n16MX
uhCww8KRRR6AEZwaSeqqwQQc7jbvV25Q+Nhh5z8QuS8BNcn3DQdel3Dd6wiZh/20
A9xTByFoqv98YUFr2/o/9fndTSwQOsenSskUzIn9huICVtOugbjVUm9ROxt+8Vad
kXxOC17L0xghQYcoyix7VwrXr/tRvBxvJJd9DuSgPqoShNMbPNlyJONHbzkY2a9H
lnGkQOrjBX29bErSSvo6Si21SlrHQsbhUiPwlG7ruDwEY4NJ12oWljmN4qWC4j1g
eq6uWysdeNYEolrYC6h8jVuZYdDeuKdxYDl3xJjAp/T4p8t6cs05rkxnBxF1ePLd
zDGwYqB3qM/0/NhbIHvnqcvIa96N2zc/ycGu9ISER3PNaOyY3CMvbMDHQquJpePv
kln4fErO/TfKveM/DSYAmNlmoHvp4vBJt1H1BA96byA/OufC/c4jif2T5cGhhm/E
qOpd5ho8MgWRuNXhTy2Q6l7kogkxXebzQtWkNFpBbZ3BCdXmmMeo/NL/mcSFlUNq
SPg9T4/YGmL+/S6D4JRtZukP+v7++1CNt4gjetNBtdkrbzsezd7Tmcb+/DPl3wKh
9svpz3gwFbd1RMHa5dGap0UKoMX4OrYHLJrSmp5pqmBzL34d6xndL2+kJUknwQco
xUoGvTjyvSKcau279BAcSqEFK8i+5JAIVVCdY/Arpnq0pxfRncHIyy+xa8eHRcDh
SfMvt9fbtstTKCZBW9W8eqIlC5jx/It5YYJT5elTVO5IYbEjB8mojIT6BRjJAboz
vRbJm/V1iCTunwH0nQerAebBAcR3LZG89v0EQfMAg4Xam7He+IYA18CkT2pytcRK
IVf2VRTVWJYOvPv7Y3FCha8tx843DPemfvgQ1S+GiuFexSGS/WokcrXFus0o9MUq
k3DDEPg/zfP0OBWHjPG87Rli0no6K20ddrWBYvUiOUTkRkIhO9a1xQcWCHO6/Ra8
V6/OuKTDwmisQsc6xeqrqqEdIvZBae7ElhkCONwDqg6Fe0P6WYqhz/g8nCdsdQ6f
KDnDnsD8dTDRQ4cht7U/qU08f9DweKWB7fsAp1hYuX5QRev445cuVF4xCBAKPIjc
WaeIDmTitZUCSwzRl0v/edKbMm22u/EhsNkk5Lg0TZusmJL+V4wnfJbirKR+OJta
XlC6ozp5H5cH1a8x3EBhYDCw5Oj6Hnm68qKNmJVWuhkYeOsd8HA08bjvbcRsx9H0
8a3OK8dESdFlG8+SO9URgkkRvqPGQffUEJcgmNoizXK3m+6CjgrTPYki9b115YMd
ev/4pBD9GcClSAuSr+Bir6c7r4IklXQ8vaLJioNPSeCLK/fZ2GMeC1YtlfTUvwhx
siqTAwXRfA+Ik4ewG1pcfsV/dsqs061d5znwXomVdAUC3xnncJxIF7qV4+JNRlCG
kHw6dGmNHYmXEF5Rqbxs0OlA2f+BI27sIU8M3+GlaB+gZpN6AFf89lmSAhABjr/V
Q3HHQnSI7rVCjCKoXDcfg1BG6sMlubMZHQ5wPCshUwEm15f0QcId3GQJJaJFXFm5
rT9G/gt6sws2Vf3VchBBNR8RTVPKE21g81h0eQy13iadS9YPmI/Un6KWulk5rtuw
L1pksjdzcOfzxnd8Y38cmiJImGKtygwEljiywzAYvR2ZTNaX9S+smTB5qoNA84wL
9oMEFbjXqMB+8Eex21/uWQI3XcI3V1wkRevjhPAxIy8xrDaz1WoJm3skhPQ7lB0x
ussIHRtb2AW1PGh5Bo1jlRa5U35Zeq0bHSVJY3pFwxwW1HMzTfCCMNGoO9zfzSM3
3EbNxfEWuNNx4eFIUm2+FYIa6fMSlzg7hxmL5xTVqipKJi4eF/AgdB1+WEofxivo
QmBiiPSooifzqD73j8RkVFrb+qG4F5Z/6nrLsqWH5SfIQ+2xX5FryUNzkJpF4L+J
wxHa62ZDFgl5/M+G5lXp9HUJX7GFpvkaJx9oJpG8TUDThVB0LiqzZpospPyZIms7
LUZBv5LLMW5H26ThUWlm2lZqWucbKJgEVEfG3wTPZc/4ADWM4snjs7hiPw7r0zaW
x0ldm1ofqihpxHVlVb4S4c6qNKIopqQmjzXLaJxDpSlQyTXFUjJTTCLNyQ8nd+yv
ZTGTbQwSPmyyoB4IqKnhkt4Z0t4eRtscPJ9jDXKaYl78FCUjyLW1YPINucGtwODm
b1RC259nKxDEO+OKcxas2YQwaCFUZpfBOtk4ud0FKr+B7l/Lz38UQ0ZQJtMg5v7N
BJJ3TC/8dtYeboDqBX6Fxd7afRMuYmoNah57+/tKTFqLCtOza9sQ3Of9PEjHy7Uy
c0PPL1dhOBGtCHDUZ2/B33visCZNO8dDWVEnaqns33/clN7sas/z4FBQPlUwtd9E
3kB6E1JnCa/H43A5NDfPfk6hm+01DvDQRV3oUmG75aMM9+3C8q1r+fNwURRPCkob
HXHcLvaIENKLZD76mXD0OffRcKDYfgpNiCXVghsGzov3B748V02VoGv5qcqqIDTt
VVMww4pMGOo1gTp3oKOO6VdaXgHquhd8ZpBryUTXVUOqyT2hqdmojsJB0lItgPVl
JH4Y15xErXaF1RCtzxJ4VkCaNaFbcejezLtwnrrgx6FPiOmtqgNLth8DemEFEZgt
xmiMs+VMxNZ0Lj/75ufMtun/bewrPPyqbMSA6QZPLc1qACuBdcpIowtBv+CL+stW
kP3B4TVKhlizyKBOxo+CECs2RSTqinrDcBZWJTCgEoi+GFdTxw90sArTZROEff1c
Hr2zIDNlzNH5XQW1C+yjgp+Yhr3WsdeCCdAgtfi6lnxwvy4vMF/jI5SJ8uAwEBVJ
XXgSS8Z9OuKmMUA4uUTYiugB8JgPfUKDcceFfgC7RgLZDUAJLueGHDzF16RodToM
XaVnkMVbPU7z5JLtkLAlZkCzKNrNmzLqB51QC7nqMJPOx2HeETVygumwLwRp3ucx
Rf/XveWrMdawJBAxFWicr/p5BUK6rEdCNmrgYQW0SlbREGfWVOvJOEE+0AZz5LcT
OqnqUM+0esHRgQbgHIhI5NB0YSRW+n5Tuh1GBTqg2K1hgNGntnHN9rVm5Z9q8eZc
kT1oY/NyfbeOpkM/qkp3L2ueuZTUm5KnaZz+SgUVvyNEYK/KvEuxOkbWGWpguLGK
maUAL2tSFjJPlCeRyVSubxhx7RqOdHVSiUeKVJKWcc57HYEy6X3dXA6xfnEPivfB
yR2IplB7gFjec6FciGw5ymh7APuwOg+FCL0ImxIiGDaZNoQw3S7auKp9RhRJ0/Sg
Y92NSrhMPwym7OpLIPO934ppXEfNKIUBhnYruJizo4OL+2Yn1C7wkSDNQEMHjZGR
ba1OxplY5/Mlm7C+/avj4WGLqcsZtSB4ckvBSVOlQZYzyXlP70gWjU865Yw+m4XU
/Nzx7MDwRzujuvxZCsC1G3Z98bmlkRRb6P5q+m31T9SgjaoTZvTbt+3AZaLxHA7F
DxnOoUeWqzi9hY9GVx8f3Dy8LIrKP2L3ztSLvWlopBMEzlSPN0/rK6UNoJxJbXgT
3RJn6K3qZqbOq0+hrsvZ2jmR/hgqDat0K/Uwis3Yqv4HefmLcN4bPTJZTgS5qE5T
Xahm1A6zZ3omUwaXhdM6GbZd/bkDzag5F6y2jukpCO9VLlTKWsDNufTJSkT1N5s6
XzhjHWAHsrd0PFlkPjjS4zgyWDM7istO76Ptqtk1OnACbFgJXtWx+k64fffi3U4n
xPYn45L0O1skDK2ZtsXr7xYxKCoTRa7eLzAHrTv+DINiDSTfGjt+JQBa2n9AwFae
Ih659bSYYtLcrh3wIFV7/jOBdqzVGgL2h4uxgHPLfto//s2RP3CJmAj81T1jrCpc
EqPhYAGRZ9IZGfRgNJv1nrYFYLEzBd6gF1KF+nCkuUEBSLWh0De7FArsjCd2ltwg
+GaDDtqEzv91Q3mOaicSCZtQJ08qosIqzXsVEAxXNMy+BIGdwDuHfYtA+jgP3d6v
igWELLA4VndVYGnyC+Zq4RotbgWjKcXKtcWFojxRW7NwlgENXLaIqPWitGJsowDM
1ULU9impqJy25CCSySbsy8UrNugGsTcexYpElhhqEMvT775ks2cBvXT48ZLlkyfC
fDygmV5qm57Xk6/xgg7qcQvSCD9/ChMf9aOJ+G4eEZBZ/BKkQccqTyJOruHtTo24
sBG5VtURmZYq9THqHKYCXhY1pOu35RE1jf3g+i3a87JH0jsAIofrNTJpvNjzDNG6
a5/zY0HbZvmulbX9NftC7b8/wgIDeuRpMgBrKY6cF8dM9br6tUFQrf+ItGTWjZe9
iD9KA0W6buK6575TKB2GbAMcBr1BFUUyP6NrOmu+6ITz/M+tK1+0ec55O+n8Vcz9
4GEydLRiKGkfTEwJq8TmhVjsUs0IEz7l9wIjjzfAYJEKl9zTkEWocDzmd41CNyWV
+gITR229STgN6m2lU216SEqv8GkvjoCZQ0FiskCFfIt4SUEVE+Ox6B2wcNKll1ZF
dfxjNRNrsADGXL2WSgDIunhAzMaC9bFVbKJlVRc/4Hp5oLP/O7HuRPbIkm621iSi
m4QcC3eXwpL3WEzCzoPjLOJwn5Tpv++GfVj7QfOdC5qk1tjf8wjpWOaYxiEoiQ+U
+0EiGSMr6o9Qt1/S/D6ISqi0HDJ0X196dpwdDYadSuSdpgnPzxDCA0ECuyD8jpea
feRRFZKxabC1yjvKJZe6iX09LXu3id98qiKVch0BdpdYVbHXVwTXbfS5XZ9nAuAs
wOtdNLMPSLvqdVQnx4W/stUacqT3tc5cPpMNtEmA2ICOqSBuN0oNKRbL4F7lNLjX
IphDnSp9v9cmepesbSw265wiYdxYU/hUDAhOOfrTqejVGc2rUHuLGrgeDZ4A4UPp
FU8i/Oq0kkRWrj1kr/jNh9DGFD2tmp4GfgRoYhEvrvN46OdIYp6/b8UPch45cFi6
QU94nYqqVejLXpLqUtaGHDDyitiffbqaS1gpJOOqKCR1DYSc0hPXjmHrOBL9d9Ej
6IkFsd+QRlhNdkuQDcgz4NkbI/JW7yh3AS5Gb5VIQyAEuaAIb6lsCxZC1ttDcxP9
e3uSE7LkVwcaItCNgTIJZ7+qyQALqEUTVaNeyMIDMg0RTWH3JzQ9+4aYwdMe3LDF
i5WAaRra5I551Fb3wmHafzl7PjdTMcPNchGp4DESxHEcFBMCVc584LVfZVRCyqi3
Dk6/LAV6xhk2qabsXi2As5T5HMDFtIDKOJljScBk8if15tWOnb/JTcQtYG2R348x
A+BTpwGfVJelboQIkCH+PK4oqNqq8fGHabZonpm6KBBttndBntnEYwmOq56Xx+vK
DzrhjsssdeNPb2imgmJTMd5C7pPiwsvJ3GP3eLGAERlQY769tO0mAsap+QyGp2zJ
8R9zdBgBoGuSNriu5udo6mxS4OwC3C+CGEwn4S36G0ZvlmsuNd69+OthS8eCLsHl
0+t0YMDZSXa1elw5dBrAbpMzeeDFC1BirOifmnaCxGLTtiNpKuNIU4FbbAdFETG7
Wv7laAmVxMxUJPIn/qgas2PIVgDDMuHiHQ/npLj6dCzv2zRh9F3Sv1oAXPvN2KiR
QOm5bGpILGBGTmE4GJonyZo+noDUhd3o1szXbw/cdcTJBL0aa+N3hNPtUX8x0Td1
4xoQOR5xD/r5INBeppQmtvl9QyKcf0BxsObxnQQFyG0ZT8Q8nmMQvLgQfUY4keb1
QPw9PHaRG8aJqrK9/hL5wkX4aYcGT18f1f02ysNwCGNe/Tc+8wqYhzK4Y3ZSLzo5
xCBjEmhED2i9OPaaFE0egMbzSNIlk2A2rCTQI5Gqm+HQ2wbqdSOLe90zzpSIGGke
eRbqrxQQnzLVrRcyuy5c8yejn/11atl53vYF8Yi3ghqjG/lakLZ74Kl2hRrbPhDc
H5344wj70Ezth1Ww8qtCPJ8qPgw9moWPTzvqZQKc7cm+0VGiwUuEIInqI+adH/Hb
GRvf0m+XdL1jnyeqeDzIO2bbV8+RAAVDMsLikDBC8gZOE8sKkddM19G9gbMuoQ7R
zXTAsWUsqd8M8Kqy28XrWdBTbnK3TJpY6UyXG4vA9eXz8xRlKv13Wy9kUoMyJRFb
RN/XRPZJgJfL6Ik29HGAfFIswig/bZfuO555gN9gE2R2nfq73es05Rx9DzwgPqLm
aVg72ST9xVXJ3HDC2MpzYcyLQlrH+SLBA8z/Yg/C7I0iJC5Ri202uGbgbZLlAoco
xwXbSrTmOSmOIMo7Jfl8u+zLtMtreOEOueDNvLR1412lzw4ry8AO9VC1vontlcSu
888zL1qArWdWpoWsrbOutZXZGmprvfKcOsBVRSQ4w/RGfLgZxaNtvHTEE0UCLHR1
kqFtmphcJ6KuLOtzGPv2Kc8OT+FAcvcOjd27/32xUEZMktv9LRBYhCxtLIXTGW2+
FuEvi+SUreL82AXK8M1NgSdoNhztLt1tYmF88ccWpbyJjko519wz/66BnoZ8w5nO
tooZPtV5/xGwpVIs4dBL/FXJH41SV995pucM1EAnbv/716pQ3GedVXakPjc9WcBM
xnbKBuMI1absIvJeX2CGeMomwqnnR+VcFoTIvTaK9gE8i5nc+6V+8gHmyWBtYC0J
1q78fgWrjgDmClaBRNm0F6RF1TXwfmEYp/aOhIREyT0jKZGfkD3A2BFRjCQnf9Yz
Zw0onFgTIbm+Fz8vs6lTJ5bgeWvKwBDwbY59MNmfM3hk6KqNmENc3UOFhDxQKgzz
Z8qXwqWiZjPJo15PhWMgpc/dVXbsXOb6Xya2l/uy09QuRbWs3NdkX/zk1pGdlhGn
0r35FAl0h9UlX+yoBshEkh0NrVv2TPRgt5fwX7FvwYQh6hOc9HxqIagzmcAfFW9u
EDa2VUCM7CCjqmbTNTsSxgPX+hxTqvq2ggum1SYbw2RErQ1yJfMkSzSHeP+kOV4q
SNB6zHbtwEA/N7+SS5/pWjmfXL4RoVycTiPbxvolKWVmYi2oH+BZAWNvnoi/D9Vn
KKFYY4QwVOIQkWqF1FaIpq+8zoboZWh8ihnlmgmncsAbzJVIkuPaOir44n/ztAFc
lKpqYIYQU1IjcHnQ04oWILHyS5ZDgnrnjvuDV/R9CFuUCFN+xdXx94NhFI/p9LcF
6in2f4o8ux6mHbqapJhnLEadiBe6L1KEjGI0UB8ef/OacSHaDNliQ9u71HHTimOu
xSxMNwGhIXPW6R7p8SXBwK4al8jmqQ1wDGVo3sIOYtnof92Iwt1OCTOqHjyMDssc
HRrI7EGmlpIi+vWs6HZp6JT0Ukw8E/f4IBUQBrrk7ee8xJUr5iXLbQ1xYVGnmDKx
EkputtgtjIRwPSLbzDiptNRsAeKZVsHnRx+f//7S6tDK+Y2EUuIcN50yQwZ5jB7P
IT8XmGIGN029Mg+MSXdE0gdcfUtR2r6CIflaxv8x/NBIkVjqu2Nf0hqoAnpqSGfZ
wnik9xAMWC2c3lyHcPtTvyOEC2QuLbgWTCaQh6SRA/ean/ZlYfahm65NSuAADz0L
UJz2nMIlhf07CymS//V+mYUtpYTK4zcXA2ls/40blQbPbnq100Dx/1N7y4heDasp
+dBRIescqYD6D/NH47TSptSPMODu2eGaLWf0SsOZhP8HwiJboZ4CdGOVjvT7zPJi
MMOYd/t5O0Q55DNzVM5tLH0FGvLUXPGrwbzYWlCzucJfPsjMafclRlSMAGXR+JWz
ZVbPe4TExaG7GUwSbBBUHaMW8mkbSHwpjcSVCn1keIVjHSYjSjQOnp7Ugx6uN9j3
XGl3ANTiBw5BqluqjuqQnz2r+fkvRlMD3bI1HSYVSR/TMlKaJGZ+0Tsk3f0g1/qZ
lxdo2aM1MbnxyEo5+qehVFvJMM0/r3qdeslny1f3XOMYdaN6Regnzr0t6/b39QVe
sPqKGSFblDrcXfTDFiiDZTFE3MomVdGgvaICVNv+j5W0pKYPy9NEHC/YUA5RoPa1
ek5P023VFZOBiVBSyrbzU/bgQGFB6CrMrhminqgbymw9NoSTXFh1mrvxf/m9gCJJ
ggHJNLwcA7YtnZ6Sfb4iZcy+ZoRGXWiJ6Klkke1weBrpt1REWE2yX9ceMWoSysy4
bAhpZDHoJ5FDuNFWPMNUP3TSD0nkKdxHmZlmyr+dUjfuFpHM403sktSzSeGPpHHq
mR3AyWoyj5UvEW6r/SkIk9M+Lrrw5Qr3EYsGnMXm+TKN4GIxOlJ2NiJsUq2lysSK
60W03bQ/9H0WcMAY218ICvH7xDxuniq73QWZaGrFZixoZlbuBTpVTDNJwQ7yQxeP
CDCZbGtoQTY6VPns0AAQb9YocwAsu8GImtAvmxGHXPqkzfjaw8j/3Hlvg6uQbQ4m
/cFss3lCLEsW5sSMwc8IHkCfQ10LftwHsDb/TjYqpmxnBFTR3zLTrHrgOsi/zzQM
XhY17q9pdZZ507qHnxg7FfZWrLWLvegSkgwhQXWK9FUD30aq9EG6MV19BNvQOu4D
l0f2n/+/YCmgF5Vxh5BC/SEzaChrCaMPSwG0FYDC73UbBkhiCR4mKQ+os8UITqHn
N49RyuCSDR230RiZ/0AYewlsmAGXlAyvh1FqkouDSsdsRelMkdvidrC6yOj08RS4
XjAEd9U0RbqfUCWIXAOPKFhaTFMbLRA3Eo7z9h6qtfqjHXVYaaSegQbmf/xQcdaH
rjYxmin69BNkxWAyrdGQaZl7EucZ9jDCnHhoMuwD3Iy8B/BXTxLd+GnERMKzcN+7
KQbyEpqDfgKzpq5eVF9ll/v7tvAEryQgi6RkKbj564NhPbYGbIjr6Eu7PzTtPLNi
j29s8t0GFCYvmVJCES5QRhglb4Qyla+gs9WxMZiA6DAaV/k0XfhREPRa3cVry0cC
KsrWXAEsy5ZujrKrQmlyAKz7IIxYOVIvK43QbrpxUXjA0qbrIe58G+JIo2z/jZQg
PATfv5tu4PlToArnWgZpWluVQbNz0AqII4mxepTm/kHEIs0QdFfADNnoLA3+9l64
M0IL4Qxjx7+t1+6SLuMogjTqTqDWkf6TJYBcE8PIJevQnprEB6FmTPHn0SWkNOII
j/U1m3XHlVX52kdqKwzZwZDCHYiAKEtx34A2/e5UOSs1A/dBumshB5IKdDD00RFa
VdixQB28xZBQcMmt49sIqwCi14EDgY7NvUm3mB5wYtpqMr7iNoyCXQSxn5XYooHY
9ty2xYsshldafkx5QZD4EcASyTJ8dbNNoRGvSZEmJFtUpFb4/ErnMHorH6ccj8/U
9f1WoJn7YEs7KpCWcCwZtRxSIbIIKYlSglq7l2IGuAkA7EHfcJZ5FHd2oMrttGtQ
NTOId4d86bIa0/CRsBN4yjKbvaCgAxjI6jIjDZSOlIyHn5em/vHGQ0eKQCgW4lGe
vnrrgr+9ix93M2oaSW9yEL+siKDMF5IM8ezfKapKWo/gtWVZ8vNdVfSil0hGkpZs
hXFW0kD6XLDvrL5qY4o1oVLTuUlwSM/WNQeoNpJO78a38EqQKAuxnEQm4OSE+h5m
gsZQXkKNRor6U+aS3w4ZL8WpBAaO37KCh42rkiyl20+oKT981jOr0oxb8s392uRr
bpAUFOGTIXIzR5udAkYIt/DL4BCRWVsjhE5EMzTHQM+n1r6FAPttZxe1TF2isxeC
AHyM0zM+o79gQQD+gwED4cSAbA/IDUtcaJpSOtU4UNlwZZc+n3Im0viCVmP69/pv
F2AaMK4E3J4L5EOoxUTazY6seSp39HaHaaJHmNM/yQO3OGWkLqNVnzGqSBKU/S3j
VfRCIZsdlB6YPoxsnRlHKjhxrzlJg229O4PNu8ZXZP+NHg7u05tKJSYtvrW2xaJu
1vfgoEtMKF7FyTO3eOWXaLFcMz57wnWRjcNMJPfAdVLL2nZJIYcFiFGYYdS7hVVD
wyBYaVUtKugx30VGQx7BBpd+0WbbOhWX/M9ZuC3O0C7vHG8WknQwNroKM/SHrdKy
oMMQ/fWFQAImWycXyrRb5sbjTcZEfKKHhzLWE2fhHUQhuqYoGnDue5CmeGLXF6Dd
EeJyBUUsXKDjiH+UUJOTGhEv3OekGc6rSwMNL/oFpXRYqAjB6Nz7UkRDNlV8uwZD
YYW7/QPTIak/uqULs4FCKKSaR6ncNfudBTuSZ8Up0ts6zeQmkAzb3y5pBdC/eIqe
/Kpu9Q4FMavMCKfjlfZdgWI/QwDmZGHt9VG7rpqCPoCnvTAqGV+VgnJms4hNibvv
b/fSR9LNE+B3ybzdRKZA9tkJ7o2AMGxbhC938Tu4aDU+0tOr6cH1jiZtA5P683iB
7LY1NEt7aGFmiebeu8HepgNQnusZisfzC9KT4KB2WLrl/ZY0nm7bX0t60JQN45oE
0/qVRLrbUCnLLEXiarfy+6gqFFRY7c+5oVeaRD30+aQNqXofnrZpqyZ4KcEof8KF
fAn85+2f9H5CocFOjmcLimDiW6s67n7VamzZCnqSsBvjk4fEcQLjoXvfLu7iUz6D
uvZF7PMgLgIIvcIIzc3bCvbUKY4La0eziq5Ic4JizpW2zZL+mDr05/03iSrv8gtx
Lu9AzGFxBbq0H4OqnWnG69eeY1PiU3AzeOx6qFgYXwcjfuwGEJIctQU/irCF27Gw
QBsDmT9WdUUGtGhdStywuqhq2XhdfTS7pYfXiZ22sivEdoT87wP2ohavXeykbrNo
UsApWy/1ytf+PDZjixjGjEsTJvePij6/q7ETBFYFTGKX+Dcekb+1k5UG+gs52XES
1DRXuQEOw9CtbT2xbUUl2WHrzV0ltvuRYs/A9m81GYXVZx978HwRS864yW5bXQMq
dpYFq1/BOC9MTRtUBSGDVtWgAj+Db+BSPwIfUPXRpcOyFH3vIXboBErCjBAQzkcA
zdAMB81lyyzX3tD5HHyLn90UrzvG+N3ejBfQnnsNg0zl/Ks5Ii7UZfo+DAQEJHau
1gJfH5r4cT6LabdFlnRJ4JTm3fZUTg9QRZn/LUqz5NkSRPLKgW2aQK5YKSaBWN88
pnrZDj8cg4Ep0fIW6I5mcIexyHpCUsUcIvFgwTSy7OjwLqqh8IlnR8Cj8djLTXC4
LSIevSu/TJUHjc+QXIWYxFO5mb3YV2/Lv5n86z940v3+pxsdiSBwmc/7NT/ffq/b
+9v/OscvAtMRVNzDhZrOq8TgiAQYJPjq+mO8ZenEHVPluGaLSoV+FrifboPgqVD0
dCYbN4DfJt2UGPNfisxgJSlSyeGYskoAyO/KQ4w/VzEgfW/nvCaosNDfwESxxNiP
gCYhIsQ3l0xdt25LUUQd37dvII0qc4Rn+pii8qgEjL+eDMW4mJNCBMNEsd3pJ03O
q9xBvcZve9RCD/DTCJ5UQUYpSe5Ftv63kqJuQE8v/IRtEauNt3wIQknkaeRlAMTw
/Bg7KPo23d8HG/8n8tAH7Smu+n/QFFg/sSlgozKf3UuTru0jB8MDC8v62JanEgdg
mHou69/h8fzrdLErPLBy4bQusSR1rKso7QTXbSfuQeijI+7JdsS8wu4mGgEBoPZX
ZYi/D2T+bAcS8FZ2o/6FD9FvRymFeBGs+iw+GU1n9YxtEoDAx9PXEfl4g7q0w1cz
pUNlitvdeBUt4RLzzTbLYzNJUeCfM3ad1z/kAk7lYmHI33fxehG8zuFhgAPRUeZg
tYahIIY8tBDioTQ1sDjWAIQM4ZLGPDNHxYJI4naKnhqw8sn98Y2r8mzNR2VnZU/I
XnrhI6l20viwPkyHA9JZLP79GghCbeYkvM+ouS7fWTihMtg3ttEpOTYRVf1vHYjO
hniht9P6g8yADz7UXoIUrIK/4Po5X5ykODq6bTKzWmWuJk6O+teHJ0KEUOxES9dF
JNsWrqkYSFVz4K5dzcVSU4CrAUrR5+Zzl6Ff10/yhHmdM8nsO6KGz3CLxWPmZl8+
DHp6uI/rFlcODE92iG/PAO1NpJ9F96qzE2shM/2UqlryVXNoQ8lcf3ez1lrqYt5f
3PEuCKejvND4l0vmgd2xzCANi3nXl/ywtjpbjLFOixass/QNoEmDyxRK0HxthVrz
17elYGQ8lstZtVltQwdwQWPV2Q+3LmSWZlCfcj8xmllNBzsCKQ9+1VRNVecghpYc
zk1GOIcVOVtO4zeHR8ucIgum5PzZu1wcGr5XGs0YY2QpAytfjx2GEo1ZwMYdbEMh
NH/5g0W1o1AyRtnymbx1cq5ZrPiDLSM7znfP5Wz6i02L76o8nsQt9fzK+gtQ2clY
5Xc6hh2i6cfhLd3yfJGYfQUqomdNqVvMoA4jwZSjmjEqvJDeuTSgNhVLcjk5fbKT
ZQn651DfR1aZTMrhrKszzR8UtEajrQaRhpXpFc/NGQfGc9TjHOtnGMKQO8mIeDNH
7spPeCjjLzeQEoegOmVxjoqMDoNGsiMXShPx8H1GFckEaapby5C/qW+cZVO2KYfD
9hOtBx/73HY1kS6FS/pX+NAr/0kxat3lmLKkJezUZKkuXeBiYdy0qX+qyxQI3H8H
Mw9Abd4CiP0UmD/UYl+7TNnlCCLU9mRadd3mjYz99TEMrVVhJWQiWbTR8fg5OiUp
dDsLiwNQxZUERXmAzmua5oKDmx2PmI+v9GnZtEXTkDkSBn3pWkil4Lp5s4gG2kyI
ZDAozd8JhcIxcR1vgikSL44CIsXVW/0hO+vwwT3mU5ADB5NGHvo+NqW0111D1Tw3
DTNvvsM9YQuV3M2wjnnURkFXSl22yq7VTUKGxIZDZSxrML0XnzhfYoag5+3PStR6
SVGW1npkZRU6jN3zkJy7ZYwkvrk8LS/UY4E+xeoJ2vev4NyFpccCnFnleexpOwWb
PEcGIEl1Ej8WJIlwHB33zo+smqP/Hp2w3HJCKwCH5u5u0gZtf9NKs+vu6Da2/+mw
TQXLV8O6CjNYd20PE9IWjX92sK+UfBRnRffKW5dv/vhz/U+3T6WpqaHk9UU79r6M
Mvz/T8pxOKr681XvJNst4oxkCiJImGPOH4ODYSoRYKlqvn1zvT7rI1dQcgYgI/VU
qLKmvMYD12Q8wQU+kPQLdGGJReNL9GPlpECWFVZoCDmTuNShkWD8asCgTwENwjkz
kkwW6OUvTokDkcHcYLOvWF06XwISp628N86Yehejg5sLja3juurNX2RW4HnQ90iY
lB1SpuV7t84NjOS2jfwPTTlGuTlsqnysrqqgkrN+XRYkz2R3AJAmKWrg053SRiIV
1Hz6664pbRYoovwCxpFLYFtg3Ud6BGF+h2WFbBr4umpCSznv8Ky3KnkjZiklqd39
vMQ6rrN6dAsUh0h75kS8yESTVut7VZl5z+IJT0mse7q/UYnibBULfPtLrNy6/uVO
KYs+jez/UhYxgxbzX9nNuva2oOuXTMewLBBHVWviFsC6DCHupI0LAPXbrbti7YRs
2Y15GBAluLsOOJxx59J9xhlfMTVuJAj5FTYKf8Ah9LYOiKiAcTByLGFnoijPd36P
d9qXdXXlXYlZIX8zTpO5Ka73q/8GRTgU4wA617l2/Y/7047wBKvn7P0fdmFgLx2m
U4fRdOfISYfidRhnarEMoGhSv59gaU/xsASZvh8n+PTS3csvTUStQRyh/GbdK0Er
tq80W1TWXj89hjLLVZhEVV+0B88qVr8gV0nCAU1KKgem3xils/5OfxKE3Z926bj6
yNPruKPXQPYVL5U83Pb80hqRyr32viIXctg+JgWXGhbwFT9eQThwfB05Acc1TVlk
ixnnpdrWuoGca5xv1CZK/ykHdz9ASaiXdUFci2wSkZrlmwISjcyWAtaO6yEj+ATA
UoI5eH513xfIOHuME7h8lrNsMtUw3ckhIFayQ+ttXIZRIaWSIjCmNfTD65STB5w/
Y3YNFZvi67eXKDZlJh7j0npyL28CZ6WSCCMxIIPsLz86K3VhiIWYjigKkbpwt7ju
J9nFJnEUFWlf3hkPkUyDdEs20Ba0swqQCd+wLdUBqczozoTQB08uaCSk0IpJkJ4C
c/MXEdI8kCGD4Ty+v4Quv7KDP23KOCTCiuYSg/+oWXlWfSDW7/L9thL/eNN1Qo6U
XmHkkxkWmW6611/oPG8fdZ5iKApjaW+nuRUvVADt1fXIzI0JqBeInE3/FSbpI0Os
PrU1PiaEDpHnE9oZUCdLrAIWAbKAbK7aATXvJBuRWqb9gTF1juj37gtyw+YnL4cr
WPqVcGXBxIe0xywxudET0ElANCnt/DjZw097KWv/t0+wX3EAm4cYLqOEq+Xz5xeP
VbWSLusZRePm7VqDYVssxxBNF5jMEN5nsZ0nhqrUH0L1Qje1mBXQBUHZuKzxLlI1
/d9LPeQCrqrC943+2qb9Q8Ll0ZZOrLaHWvZKeYVMLtqoju99bRyPBYjMy7qn44vC
ONuTZMq06BJ3EvqW/eRI1dvJLICTnZNZwL0ZNqC0Mpg7QBGXPGqplJjf2cxdsoUK
ogAM91baeC2NsyoIUvLPxlxC/cnqT/ZA09HsDbHNaziDAqhbMmvdivl7osy70aQc
3LvQMcEOjwsSgAONFOor8yb4T1e7g80DXkvQzB+bEzZN3I6+71HpuvkGMdKR4PoP
CPF7yRVi5MMkBqgYqVt6JnZwcxfEeKz8BYp6JXd1WgNyj+7dVZIwvpJPOxSZ8yRX
RVIvhTZ+klmPE9BCvtPvUzBgzpNbszcbbOP4qYnW+YN7uhASAFgaQ2yUAqkgwolj
xoq6yrheebpR73ikSFnH09mgnR4nJiSGJZb4Wml+axvh2nT7v9pWc7GLZCyE43IL
LS2NSqqi4iVbKP7FLtClqgdnEI16hXEoY2coZJT7y1JSHbJXrlK82yxIQiFFPB15
7rDxAwWrRyBEE/Rxo7mLjRUCae4dtVTERxst/U9EiVrz7kn6PUwlIJ7brl3OrBng
0QbmA3VSWUtiOgPXU5wBRV85rzUpwlGSuGJgD8wHFU+PxspHmn7nwGhsS8LFfBZA
HcmcvFE/vfDm5xM+1/Rp/qX3OhvwJzJe5WolaHq/5Jx4WicKF0eCXkXy1SUqRmhi
F6BCGTWjJTEs61rmUEz2wN9oDHQk1LsqPOlXJucHE5/jq8lPdWfa8oV7i+rygIUW
V83p7t2pK3DlPk3gSrqx0dJ7erqAyAroOEMrwgOa+GUNsMlCr4FPUgRJfirYFksw
J99sIdL6SOZQgRMvQg1h098ALH7sM9Hfml4Hg84j6aKJwACEwLlJ9hkxKnPVq9M+
af1txdfmbfyZ542EYnYz7MLiOgTg+PUsBhqxnhPzjVW/kCBGn+s564Xokf2G2R8R
V0ooVpUM0akmiEcMip7v2nHqMS+z0onGmzm6uDvxfVf3y7lWc0JRjj7T8q0VJqdt
NrCjlieSNqp044GHTvTz19Kt1hRpbB7tMtBysGQqWRPpNAQGSJFcEPmaOUcYpBTf
tKXNe2Xs0VurVhFZCJVKouwVmZUAmncj18fdHQpf4uohn5IoVwBi2eFpDQ3KEnS2
v1WuN7A9q4Hd1DXhMElxFtPLaK9bYWf6eELCiT1Qdrzgr0fzPM9ZQNeRannS4Y0L
Ho+Nbfdi4poInF1p4FyPpNqvS/KxIdy/Wk2LIMnKnuYHbRZLKAToDpcC6k/59b1O
qtp0JvdxotvbN1bFPSmLLIxFOtxtDUYqafyJv0D/YpeZ4GmwLHqeoKi5qclAVn++
xKLuaMnYvSOWrkv5UDHC53Gj0ZflJHm92kut6uRyGJvPF0z9mrz8RAJuYipJI8S7
djZL6oWQTXUk2saUJLglSvvC7zTHEbIy1cqKDh2DXRFBxL8KNtcKRbaPgr6eGsSd
o1NP6R1YXel7Xip4J/VEapiSvItR6JsiZBe9ExN9hzOLRB23OJdujgClArqR/vsJ
36mafgbEdh+4XTQ5YEIpRvXgBNCnwn7d4irZ4i15YlFUGnmBQmUpNul3vUCPu8Jf
W7kn9ieTvvzoJdemtMdE/AuwAVEbqzIxQdNMHduGpWOyJ7JfdTUzwqwO3PQ89krq
BFeLxQmsqIxPsMLjD6DK/A3IOzfanXpXe2+F/gyaPREOi/x7tzXGPXrKeAl0jyqP
jIAh3Ic3IKbSJTMiTGtGmstYmXTOe4lWXmfuDQh+G5nPG8QPafkYlqhDs6F6eJrE
OsDLPYVmdYERLHIFjY+TJnvvz8VWddJkw4AMF8OFcLIFj/+ApSK9lPtC0MdLLYRZ
g/QZfo1Y7WFHwkg3k2Kftnrf8MEhnkHZ5ENgNf2BJHckhXtwusOA/p1FzPAv9tZj
2DDv725qsDydBP1NylNwBm/JYZVyfGYkswAeCwDDE9OE8vaTkK0LIjQ4aLhW38j3
rUEQByjK5R4YLRbYWrCzlj+HILc4aaFkZRwX+GS6F0OD8cg9ZXfK2dJkL9cF07YJ
g6ERAvc0cRmvMu71/bIaFcso4xbOSNswGo6fZ9322pm+KEWb72V4gY9SrKsAJQbY
rrohJW9hfUnYRD9kIww9vW4cYDjQyn+0tPKPvEtK/VohX0+t8SQGu/bGOoqdYcbg
eDjpVdx5klgJGP1vgPk3RHLuXEV6dRv/HHhDAsiN5003eTdt/2LRDGC+/N9mE5kR
QxyRGjD5FoezsVfxDxuVTC+7vQ53EaVGOlgYPbzEp8IVX8eg6+WP+Sff7IWOe1xu
m0RWcdknx8Gub6fqiag8iJ7pTjveOmFa4F1IBEXurRcqeV0l54QUiiyCSYJ6V6Lg
/HunWTvCqn2r8M7ibPESb/2+EWTtzCn3uFAoqoQ+xj/hm3RZ+FaXSC7Q2yvWWbDV
0U+8q9girRCXB8+elv8nCAMXqe7dPqKK5NURPxXI5E+7DFzEIof7sh1tWZGr/N+h
KuYBRBg3xgN3WBthkCZFqvSRHGzngXPRffj3skDRBMvxOAVxm38O5DXe9McfwB7p
Vw8Hxk2kAhs80ZFTHSSXD7dglCpfcOVhsat0ojrDVYwHKvvg6xqi2LYfQ9AQKOuQ
brqA+37qWgCA6CS1vFBYCHbblvb8L1oVJ1KXq5G78PYO0+Zl6A2dxpVtZW+fHIiR
kuHTQm9qlG1t3OAePTpPZdxDwF0wHkZ8uhDpLpJWAsX880qgBMXjVgvodsGZ6nY/
9ZLKY3DPT+UscRt7UPBTOYcsUEqPKU/DJc2sLeR7sFb/pxakTXC+VmkIX/EgNOIH
WakcTAMKAwxUoLEK4O5i0oHVOU/G52PmTKuX7OVQWERV+9rwUJUInbvUQeml4bAl
woob8vNfBHnVYiSUPPPNVzwfOqvWuX0O6MbjqejTTOGqsfUrlvd29+F91IjNTiSB
qYiRtIkpKxBrgz08pwxpYCgZtvRmlLG1CN+xhiqEP05UJ1Df9l007iqDQjWeJhKo
09KMQgV2u4w+A8xhu+h2QGvGXqNZgLPVgHD25DJnIkqtwWIz8jp7pb4Tc+LyEFN8
MLhDjYWBkoz41BPfXd0pmkz7gpJzOrC0HPxy4YAeZ9oycCwKaOvgWFs0xAWRwULX
jEI+t9ZsFJ8Iq3Z24Phx+gFzN1BNTDsOxqH4w32cozwnlZkwcA1sDXVsHPjhgYUu
1Gr5POdG4nPehMSORWTQE0u41mf6XxjYgLvwjpCVJFYveBIsA7d7M+KPAeGajaW1
3B/yiA8FOT10jjtbEeti4DxQ/MSmBb3ZZ6cIVTFncONGScYV34exVx1a6fIXmFEO
CfIUC12o6VfaWQFR0l+OKijKbDMqL4w2dyJc22f5vdHVE5S/kBeSRKMD+7SljNh6
4qhy3DPynjm5lDimZuUPAF6I1/QAHn759jBY/N3XH+H5i93D6g1DWQG/K53lBHEN
Q8CEhPlXTizEyKINnTQwr43TMkslv6tXope7Y/M4yYQLwwVgGhNUyoc4S1CEA2n5
DE3BDj7DMAXw1/AsS3l0guE1R7xr1A8UnAzBr01kRNiZ4l0T5yveNzh/tlBkz5H7
HP930JSIyEOK4wbUT5G0vfHufF+HiA+Qmno2s3pAuG6qttb8/fg/UITTiFyZ1ASA
1QBeNTM0kiAZICD8w28clWT/r0kcxGZLDhdRKLcqQaWgM8R7Vuykf2rcY89/ZQKR
oGGMiAeclbb8eEh1JxOOaJfovHoyD9dsP/F5VWaN7zOZ1DSWfkwPbnnkD8SNafJg
e4lH9NWhpB4kf+ErXLh5TlFbTJvsQhsE17kQMU+6fbxWFnQnaepSFqG6hfhaZdBY
13Yxq5u7taIVAnfk38XvkiaT3q+7ncqG+vy4TBZF0rQFT3MLUX2fJMwW7Vft+zIT
PEAMh4wLyMS8s6O5racHZSMfqA4fHXhkbWfykaDI0lj8CqfIiSMJmfzmGElcsZj3
o60nImzYcgy4cb3g1JkG+fRztvnJGHZ6IhspHavfe/qlEj9jF5YaMQUuCtTTaiKO
mRz9ZicNh+4Wm9EgWXpjhzFlsVPFo8wDssrlkmtQv3X86HvVX6oAd/uk0xwO1FqA
/IHiMSwTWPaTxjtXpZ1STInNKC1UxFR8z0BCM7wPheWUTYcDOJ4xXTR40ZqJI3RQ
y2z64htvaRvaKxzC6xRFrezBaSt8YAJpWYnAyz7PhQEKXolXv+nZiN/ohH2pnvfP
qJo9BoM3GiFk0WxYDoClCamsmEjuuD640VcKRCWV+FLL3X9GsqFj22Jp6rlmaOKg
Y2gVX5MJeexm+g935K8kSiKBsxM3CdSV3msxcWenCcC8qUzcXK1mNSMDkybd/PF6
jr961ibaBjaAaPu0b6pMfzRCLTMph9pBqZlvRywlJkqu1uFf/6DFEUNvDa0Q1zJb
6Wpjyl8XozFB9ikt0seynqNU38u6TFhVWSXZKLL/+czeaIrz7ISeg54hhQ171neM
hXkE7knrPIM1EaZRX4bJTDE6aTuw6SY3LqQZwtWWwp9zNYEHURx7BKojDGMCIpgM
RGOEsi6wDFLi6CaqllDkcds4OLh2EjO7YiQ7x8ihT/dN5kRH5Vj++EF1POL8Sb1B
xyRYZa2pCwujzd8IB1EtK5NWEjHNMLfvTA+Ad+B4ojq1f+Z9YVCdBEmsiXwvw+Uo
i8Op7kbkCTztamWeWXiQ4BDqKP1z3j2ZEA5wc6rHjZ6+Ebeu6tr5+HvN0Q/RyHLx
h4mPnbpF95zFyVHzC+fNmAbZr7Zz4q2nNQXgbkOF1d6uceX/2jYl5rlW09k7YD40
BG2BoKVe9La844sAQI4uHlV8neWA/C0b2lzSVOSHnqF3MXS4VbZyQCcuJIYi//+c
8BXEqLUWTUBMn5TEb9pUC+aYwu0OXO6CXMN//jc5pt1o9ivbjrMO0F7n7kNkwhL9
F7vMw8wQI8rTCojqpjj5hL98T7UI9qz54l/YoAputXVqJBcHhvBA1ItbgfzbkZAN
uK0D9yNn0j3kgPkRp7E2fbygJgfQvJDHY7x2vjcu96p88ziDNLtmym4VdU09R6Vy
lxdRkUlNX7qyyhlRmaQ3itaWqgFUFTYfGqLfxYR+QqDfK3CsSeEpXsR5g6SD1RWP
rVX7ch9cJa72+GtvOiRWYNLqcynOqLY1WwlRnw6xCjGeXLoqS2he+7AG6+Pp/a0m
/ERukqRSxXIsF6YbW5N3zGxkF3wZCqY9ekwS0UsLccXkCaodziI83XOdRpuKeqO8
IkTy6F+ArWz+q/vH+SN7sGnX2j1N4GcfJDMU5A4ajV0S5SD/iDD96cojOu/leYfe
ltNmtaaGizPphyDABBWu4HutTA9boUUu57vS/A5Io4rsNqcLRxk//vxwJHA1iAH6
TkUZ1/cVFf9V7o+qjtcRjko4BuCnJVOsITsKpbTfxJjDFQkCcwiID2rySLcwkdgy
ENrYWyArlXtMGRKqu57OTEkiZQCKytjs8U7aG82lVD0k5Vl0oFtCji1UT9L8ASNv
mgbUFIutv/HkKcJnNsTRx9PzVID5WCOfscYGWRPslKRrF1Wyl1+itbxWPnNAtktg
Vh8cmKmRbjjN5WrRIYfe1wJ3QwZe0HGpC6BcHd2HXQAO7bDO8hgcQbnBndiLR7+O
ncUNQVukCypFTaEO3JshdIx+vutKR8VrdBBwYS0qMsxcQj9ObUj1wp0CPNGiS4wq
a4/QURk3xh0Mb9ozoiT+Lx8wBMnjT5EIpYUrAPcdHkJMNIvoCsHatQU/AmRUpaLE
/4RgS0MbIDW/L+MdIeYyvHYqenQAyYi4H4UvtlArJewOgYkZC3DOHtVQeoygIDPw
J1BZc4UxNLFq3pUgjB7qee9eZxx/rAfi3nWowCFXYU+O97bG+ve7bpD4SiIf3NID
QXJlXr8Xy0xA97MykvuvhIBmLp8aBHJQV+z6bwN3HaKY17BaQA1EWyTJtigNYxKf
4csrhU4ZVc2sJpTBTD/zzris4Anb41S0LGvvPX9aiyRTrPfLikifpvHne281kgf2
d5DhVRHib25XfKlfpfo+QYX0lpBdgcRlL6osOZM0VL8vnY5CsvJ+kKHrfP7uuFwG
K8Cei2AKIGS+jukf/kl3Nki4f8Y57eilFDELO0Owdz0jL7svv/2f6W07tWygOqt3
jjwNMm6bJem+yXbejwo4QBJ5zttLz+4Ein96aQUojcsQ/bh425vtcbwWwMfdfUo3
wcgS7UAMDW9TkKfgYAWxsTL52KvroK618Y1NWyOZOZMCGnSH7g6onNDN8XN3Fwyw
nM5IlwboYAdElOD0cpSns8WZVys1y69clyWJg2B+UOKTTPWAg6FDHngGPzuwJfrK
K/2b8BttgxHwpAWUwYo0nGtK3l3om/LzptPg6psdOktCbM1ZKIEj9TFYAuGSAXkh
msJjcy+mRSG0hb1fz0MRBJ65vvoXe2yVGSfGFIkNPINgK1wjjwFJa+srZZAqkl1N
hj9qD1Po2vhGd58X69v9al65DfPbK2VYpWp3+npaKkMCit1CIgbQW9UzXrepH5kI
WSOH6dLu+wAnn23sXsxH14gxhU74iIObnplDmcERETGsMYhtfA/0MEs3ijtkqhDr
0ckMpJbguJpJQckaxe7E5ZmwAYDoOOvyl3Wem1TeENzotbEgfeY6kxDAQ3Aovlmy
WkqlTYdvZouIG+ikoqm1FZ3KzMvhajMgNN74QCuS+ZaB7EisnEx9hYzEXwzH5Fxp
KTI6aTSdAJS3f6Ro2f0mZy+QJqt6sr1xrKITtf37/e0kflGWgYhVSenZkGzJa8i1
tegr3AoFT0MuV9rj7hwEv9UECu+6laJTP61PbQKwB5FNOk3rHWsf1m2dnQQFfI2t
27y48UwHxLiEORogbhSpDS2dGZ9T23HSyRRYibyz80XeuPh6yTrLMUPhAAevp0ZO
LIK5CqmTYi82mjT+HEK9pcF849iWGMjnZfRncbdCgmxGUOqW9B/siGPt6afNEKMG
EXZGKy1fOQW58GJaUJMMVMMthTZxw32nuA5c9dQDpH57nr2cvsK6MKUM7dRmC108
wgMFNWRO7HQhFLtQtj6DGLZDYnrGDQND4l2xs3F2y3p3OXhdCd6o1TqT3ni5YaJm
pjEBzVmCK+4j7xY1gJ1+x3Cpkh3bRKhx8nnQWTZrOhTFTWyuwVImvq6Gyw2cLX84
MC8GSV+vfsxAzdOYKDtqbLj94uoGRhYM/+MhiO4iCH2uqRlWZ1TrQNBd4iYagKaC
h4Amc2Lagk5V6x0s8jBbyEVGf4cMK3QOYmOlZqiYL3t2jT6lYs6z34PbJgDHeUKF
e4scvmfPLAxmTYNajkRdpFdnmQk4qx3Q2F/apvH2KJxmsIekoZvZj8vqZe6Yks1S
WkqBj7Cc4JQESbSGxNpz4GG33SDqkJI4FA2He4jY2eM/otpXmmcUEUUOGcuyaI8h
7FIXJLohQAyFLq9Dm0OBMVR64niaCDWIemYwjDOxrEkBuVu7ID1bBHbUDNdI/1WK
om1odnIQDYH2FMzrWZ/pvK+W/EjPl4KlZx6WRijXWPEV2gmJWuEQfCUyEGPlKSCI
SjgvEV4PJBCgcLiaUHHl4+y64HNtb+etIgVbvvnHD/0sGGrpn5jeNV3TIi7RPi2z
rn/gN7lR6g5d549YxJgo+u39B6+oYyiB7p4Ibmv6YfrwG1yVYIDfXrDI+GM04Szl
fzV/DB9VcKT54RSZMKOplTK4nvP36n6DTPMQTguxHLlld1cNpQx5TiCncnSlYI0D
LCH4np2o58rS+UQ1wY/VOBW6WOpO8ps/Q3DWpU9bk8rUceHnNEbQVAxk6PEY+JBj
/oVO43p+1UTWsIe6q4v0a2iGEE6YG5PKmKpFSHVmLvmqB/w/EzVgmT00v3olVwIk
u+tJYyn6jOG0chgddmMK3Urbhg47VenHbaNAztRRXSrrs4v8+IojrXj1lhUpgEy4
5QTyTxVPU5d8Gh3V+55RUq5feoIc92h5f/2ncGxDR1S95SyLrHF3k/wW8l0ZZ1DG
SwswrFXgcNk9fRzhRnD74tfJRzv8MqW+GiiM9RbzbIuHrJ3Ng4gE3R0AWDJXz1qH
jLpuquVB9zV0HF79ArQvGWMseXlgmLf3ocRmN4998j6tMxsmU91Es/NwhaNN86mI
`pragma protect end_protected
