// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:31:58 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
FADpCDZThLSvtFjN8qNKm4U4S5xjsWuAxKzJJUONs2AHMfM6qFy3AAmQfbnbN3x3
cY/EDBVg5AtH7m1g4QuaiiAkuIYDZ8rXbidyM925LVqgltWi+4pZtHpyAlRxPG9M
KYNBvRbGTKch0YWIWvdUiRyEJHgKvO5XcTpmy+a6NDg=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 23584)
BUHU2vvRt077CTTnH+1mB3o9eblBLwKxxPWlgriq53rCpLbGmGO+a9dnVkV+Jozg
TePA7qzz6tbikQJegejPir1BvweZm4j3zT94N7vLo5vAwvOeKpKxH4GSjWMhHR//
mhLshXEUwIN3osb5ZkWFlMe0lZx90HHQoMpleFJwYUSKy8I5Zd6G38YT6WUaBkgl
4lIBQFiuLkrYIslAdaRhG3u1CyV92aqtZOAMolLqUmLWIu8dO1BO2b3Yviiz/ZGH
d5atPdG9dEIB+TZDYeLyyIpnhuoJm8DEqztEDMYVwedYtYChHDaiYjECDNbpq75V
L5fcVefrdkDPD4nSPlpWwabdplqK6cXX/C1L/3XvlhNWqUx0pQxEW9ZfjCHadZ9k
bE7qUGML63bKbDVLZn0ECmNKpTEQOqcCRoE7g2FFLPJVWr6fBsKkqzGpkbVZLvPU
74f3qi1jLCJ0N2LVHgx6nyWKM2MeJzil2x8WyUAzHcLW6u4saycnfQC39YtNnqey
zqKax+PTsxbqvdUCbTOtw5ldQ56yGyZJz+IOaTl8y3KOcNUFsXm3NKbuQIASnqCe
gmRaTR2Aj5Zc4Q/igzYqy9hiBKcAFvtbSsjdqF40C6jO935oRWwn5deRjvth9M/u
61tVRWDpkpRvYPDcU8sHJLUAxxx1Yr0ipxZXeZEg/OI6mWXYpfKkEnClc2y11b+u
Izn+mORximnWIMVsQdq7zu+DBaSaOFKNxSXZNgSqJ3thdNdstrerlxqb37pJMvT3
1whIC6YcQibJLbwKVZz51ozKYkioXrHxrWpDdXnVZcNwDs7kQ1tuGzDIEm26Bwa8
q9K1xlukrYWjbIj7L5+ltoe6kM2UFy72TaNMW8x97oC+lTH2O4Mz+K8ycCC5vrc/
sX3fGjlk5g4/QJr2jgNZNLzg6aGQQ0vR1MiO+PJ4hQqKMnBZ5wwDtMoFZdp67KSV
5YAUE/WgD/ja/5W/HU2c0Jb0SA7xPiDf9I/KTfeOOIw2vLjn32qnD74C+UoYtdqo
wpBgsE300vO8OWS7R/Iij+ERZubQQlSTi9/fElIQZzIZoXDzZgPfx8225tbK6NiG
71fWHXbis5P1ABq9bMiNZTcry4KavEpVapg+xUL7Lv5Xr0WO4QwO82bNvBBgzgim
04OXgtIQAsTFEkQC8oTuaA41fSnOTlabeEDjnuueYeuiul122XoN/ArYDUynDKeh
UfHo3RaZy7DAMW0BvSE0jm6ubgBCgrgFJoU9UyKwJZsQ2euWzeWJPh8ZjUSzR6AO
o0F6/MQhR+4fzSHkO4zpf+0LTjfFoyX23ERs9Bhibm12cr8CwYDyIzX02zux99v8
cs15SPhvdIbH64MfoX4258rFmFt3GU2HtwC6PfB4ujO3yds8SF5DlPvcwzL2Vr5P
TxF72Y8WiUHqyLmj5Z5D7EndWWhyP7nqHVPYwfX8xkcBfAS078VEDjYnZxuIxtAx
k97VvqO3I1iJMzeHjtaE7rWq4K5GDOBReF/H1RhSfQtbLqv4wl+iGYZgyU7UzrmX
+EwuUDLg9R7d930Kkd+xxM0p+fKVuCm6xK3mqxMianmElqJRVfNQMVcTq8oDG/uv
3W24cK33SIQ0R7op64yQ7PJyYaNiKB8ncgTHbvMaTmghuVfsxsrgFopjCIKsG90I
9QT/2D3SGN2DpaXmb0zxmRyGwUQSwtm2s6t/M26awyPT8gl4q5nPcY/6NHuc7nw7
SaGkwT/2BFHXlygcpqBkxWoIF+L4VDfxcZP0w7mmA/tbUC4b1iYzN16KIdshHJ/J
K/4BlZ5YEtfz0MoEa59RvzHhuHaR9iKkvKt1yq30PYm6DmJnf/P3zrRZTk7J0f89
RkiMyfRfs4H1D6nixlWcOUo7DdeqE45UweH1vSftRz3D/R25R3rUQd+nGDs1at+T
ZPVzoWYphecQjiJM87LjhywetvQFXuc+w1otcv7oMQZbrK5saNpFFAsNCc8o5B3d
29DacJHldPq8azYdPiZWXZtlVwYS1DO/N1QfKEqCLriqxRY90mWzWgfUIVkk9nAt
WwJKmDU0T+xqODkOWiNanpOPcyjaXYV3pBJnfhj20fmljOrSd1jh/jj6b3GGFXb0
TdlekY6Q2ILvcOvqGqXKZSpHbKbmwO7u8ds7SP5MoqWlnXyktxiWhP9saOzzZmra
ooSP4fkxAojVd8fYcWNiIZD5F0KgxwFkgHnIFNRbaF9wdxNDCjAJFXAqaMtnfaPy
UI2hVUq6twVHeagywJpEZkbhKgdPfVjm9QpIRCSYCVgMgItLPlOXaHqgG3BthcCb
+euEHpIf38yHOLRFHdrOReUlZhyKOS4w3yuGtyKBKYxK8FW/khAMywMSUOtNUbXe
PlllPKhG74PivbJJj6Wmou3I2o9YST1X3Vwsze+OS2H1JrVkEymvNwzilb0oGs4j
LztlZAp+l8ziNhURzkCutd4epx53y79s/+laGSDq6d7Yc08fQvBXjtqU1Bsc0TD0
4luyFJx+eOv0I0/ROcH2vPqdVICUfc0RMiYFXFu2PZQZ+0zAvL5DHX6SJpCw5E5B
PKDyeX4CSSIYMQ+yEuI9lNb7h1trfwab4lx+oYCBqSEFWse/V5FFF7n2c+bibLV/
VI0SfpL+UHmFOxYqr28ljbRHx2rfEjZ5WGQ4+ZVwGy2lzB/80Fhr4Qc5KR93nma+
4ccD2C0jjhKiLPvrtHbS5R3fhqbbSLvJaM6XFDvO3aeDYPDPN1F5QWkPqMFw9GcE
dJTe4dUuvep5xa2iMzaOa30mw0JbBiNAIi1PX+QZQHRMOLWyBpU4vJmeKRFWpp+P
FNVbndrtPYE2Iy8MB2tsCJCdO7J1Xq087QAXkz7o7s/QCbq7DVnU7jYOWHkPganT
WOlJyyElfbrkGWmI5X6gWhT1X/FkBxxcWmljRwxFWQAyVqwpK+JAvX+wYMmcvhVR
pNs9xupY0L4/FohFJHvkGNh/tRsiXxEYcaaNgZBOXAEltFF1lGNvxepwp+SXaxmW
voACHhstlIHMl1pOFbYalo61F4zNl1WXutg8G96TFv3cG1zIn0EyK4bPlPzNUtZ2
unOF7wYfzmTIrIv8vWyhtFTnJLSvauwNElgNit7LzEahKzv2zZE+QbJdUQsw+O4a
1cF2MHr/8N3eA8TzfW5alZR93K4S9Ig9X8X10yTIyyrJ1Avw/PWYb92SvYLzCGms
ImA+afNGBCHpi/RWQ4A+sMxp5O7wC14M5ja2MwpSwUqr5WFUkvAPCoXbKyGc22e7
8C1hwPg8TrD5aSGXlQtLqWOg+kq0yKJyogwIS3UdLzhv26Y+rRf4JSSwKrB6OQ8Q
9AJ2lPf+cGuRSYtHg6F9kHaSJIp4h7tCfzewGKzGbdu/HRgNlGLJdod+l6UBkdqM
311aSfI2UHiyXu/JifJxe0Df0OWxeZ1jmf51wHIuV7GR0kaFf5jOnj8fPevK1p+v
L2Di8m4yKQ8qDgCVAom7kE30tjjOwO4QinWPPDN7gRGH0Ib8JjZwGsO+L8WGOujK
Nyqi5WoVEBCn/Z5Xi7Q3Z780t3eshuqxwuGOsYOE9pZHQluQySi7puZUtupNEh3g
iC+31RnSwReAYONU2/9xbH5vXux7HpbdOGsbg47cUjvJhnNI+wqE8/8CQOD9zzN3
KuqnWFqPJwT2wZpkXDc0TT+7DNv/C0/KtKyj9dSkAewj41ROyS5nL7QcJ1dZjuMO
t/E3URL6N+qeoobtWyxJ6ah9Q2beeaiyj1B78cPn4IZKieSnn5xe8UljBMutd07m
277YjplZ3LvY4rxKU3qGC6SQle+DZit2NCxUN7S8XJdHkhu7rEaqvfT5livshU1X
A087LFyqhQM3j5nDYOg0neSa5YiGHfwP5Sok8It1KnQsj6uwTx8Qhp5cD8zAWx/J
ctsW1kUBEydLzn9fOOjtK/4PWrYP7ndH+QZko1fnvb8ALXaHom6SCHOQLz9KQHZM
4oO6MCYrwXimrz6qRl6e97jhmW4ULvZlCeMK2ZWaPpnXH8UXUz/mMFeOTKB2u3b8
c31pPVKyHp3sFCWWCSxy86jUNmXLlhvv0gDMTsgnOeIx1udaEsPiW15FcBwL2on/
bS4+rDCtX+QyJmzF1rrsd8GFgPePi0oEqRH26LS/gI1Tr4hn1JSGhQCHHsatrRZS
m/zFIHJn0Amq5VubnEx9/BTAxx44+tElzarjpDLk8J8yU0mTKkzNYL/HuF7Dy0La
SxdVFEN4lQ024/wxEHbVPSRUCRUVeaZM6cl+eiMa+tBvcHtlnkXkkFW23s4UZ9Nt
0EU+d1qNh2uS8uM5mZas+4E+otKQDYy2YzUOFROOU2wBhsP+PsrpD5rs8rxOYNgY
h13raMQMMGLbUZ2LJkpSxS0ck1GkMDc+98OI35KytCWZ0Tl9eAi7C8/g+Or/YCow
F4NsMgweXiALmlERFaka1IQh9C6tbJPwO9iDn4+vHo0rmFEUlXbsTTnR+AHbukin
q8JqhZTL9OuPKlelDfiuKGak1rbBimA3kfk4Hxt8I7+zuMPp4qQsN5a7lu5St07W
1SiS/yK7Jgd9T5tjUjrafUb4vbmVep4dj6GFFsw21kna4Fg08UK9PzlfZBLT2ZwU
4hx30PoeQzuHVfXxOgIf22MfYNu75FvDubuf6LAdfjWf4abTj+nXvwVUJAUNCwMw
2jxckMHf+OwUaz6v9m+Fyo8vlEegjRMn+JoPO0vNoX+d+vZwXSHxchUXWzd4e+19
VVDjwY/fwVyGLht0wQZnc3AVJR0NBc2BSdo3VBpXile5/SHIn8GZviW9cW75dj4y
N1oyfMgt2ug+DUFxDU161aXIrtzhgdrTYg/aVprK0bRRZSl+YbkV51xHGM2tctkb
AW9CnRf47O7FlLy7oatENAhamvOadzD/gH4fRr64/dAB9bJM0ovE8dHa/hH/w3uh
v+b/DegevRl+dg9f9nVM7GZYUw+9ERlP2fhQsZ3rGFEbrxSUKE4WmsPHhWccMvkA
+Q1JxOQwRBzczIvjMywQBCp0sOEq7DHdw1Eb6ZzRZ23aLP0GGHfFYj38M2Y1IzBb
zZLC03dcTJdmbh5cawsx5+7PBoAgMB5h2hIFL4WCORbAG27mDq0zLwQZz6FGyfID
NYzsK2PQDOCuowEtIwztmn7JpJ7pI8SCBkYUP020y1treWXz5isZdwrLlgC9ixb2
EAX4FjWa02OmMsROP1EujonQEMgpUQz81Cj7bu+Yz4+ghLOuGBFNhQvdopDLR/cS
VtHtJv30mVKcYQBQARTJSNL0puShuTAN70k06wWL1bQZ+ACUi0Dd0crYTDvvjBpE
m/aAyqdLiLQTS4+tCZJwb1Y8btI0hNjMaYXq2XwG4MgLCWcqFnrr4UeDzBmq6dG8
THtNoUhlap1uWvMnvNmLphRGbcLJn44xOmq4Mr+vmV+G83/HMa7RA0SSCCTt9kWU
o18toaHX/jiUmiLIlvFa0Ouh+I/4km3TY8pAK4MuixBM0y6A3bVMhW8hMT0nyWfP
go0lcst6AdIdIPwum/U5KplSJ4avpT9hkox0saNFw3uc2dMLOzKf8NGM+tim/sio
KZ6HsWvvRQFCuZmtk9UYTWXc4JuEgJpDNClgC5mvi+6L/C2+bTa011CyKeVqkluD
FhsY9iLpebwB6/LgKFMUKBKIOe1mJQyO8yz4G3KSuHLIyhxAhp4mcoULmhnqQ/dG
zcN7Vp6U4jxmKk1PAUbr6oDBrofOXlHDTzVkKHz6LCFA+XPEuZCsrWzBWrGGtFVe
jahPOlv2tXI1is2olq5nfrNAnzsRIMao8Cv6O/iknV3NgAwRXV0PpXPvhvyTr7R8
CGMEZXXr0kN3v8ET2gkNN0vB6oYXzWtt/nLqD/F2DHmSJv7DcsNoV214pWuRyfC5
DBwJAbR+ITrtmEAtF1677ieXl/r5f6XDOZJR90Rhnqn9oO0mf51Zw38rSpo8zCiW
YNK0JzCJVNpUhbVSS2/Tubky7ZcQAGi/7EflKXokapQcK3cHqg0cphZcucJvt7PL
dmrAaqdrrmL+yC/L/JEFEquWL4Ea+MbA5qFR7IX46xXETJjyX/WbzjkA3B2RMd0y
bWyWS4lobrA3E34LMJ2+iqBYD6mdCTV9P1Jr114nzgJ/Xk/cBZMfM0JthztuJdV6
iqF8S94QVDfogiqZBtAJ9ufqYzrvfPFuIDqoaMmTys4ucqsVEcpPHH67RJmhOmy1
y7ngpuHueAZ3ZDfQ+lF4T33PWRT8FOquBcw+9W4791QEYw5AAmmnZMCcZt20u58H
ZSRDvQp9gflaDW4gdnb+EorGn8YxdMM3VnCkCpDV2DE3CnDzapQKWq6DvH0+hiKK
ZkzXq8987HAGjLIdup1qUloo8g1JlheaZwSxfBxMRrZOl0p7Ekz8cgwqE+Mf2IxB
jUttbEJ4x/G2LqbxKTj0BKnBxLWWpUQKapGMDgswdmaNo1hW4wWr7HiIahjr3aAg
ndZcArfEYZITUGif/mvos2eGNuhzh66D6wApcZgsULm9sfpxZZVJCgS8zjw64B3g
dmJYqxJMZzSYf9t/rxutNkFO+rmn3cDSgBGhhGlWXecnx1OZKSrQY7KG4fVOZZ8d
IQE6BrUmgyqK8NcDHteGq/w37D7LXmajabqmOKRaB2YwNEzlnX5CfCmpLJ9AbGK1
rr2tG13ADpuEizY+F8sX7UE5HPrf1spWBRCrdWFzvmaotrXgN4OHk8pvmeZFtGb7
WHeSs/gwG7QpqTkRfbdc+fHk4s9fKDgAD6UJ1A99U6C5iHWrozQvrS4FaA6/IuyH
h5D3TRsZ1taOdUmDf6aHJqTuqCRfiAVu2H5PdOxSR9NC/vfzt7/irwvFtkemydZu
89wWKYwtDmw/cdzZaFAbTmVCdeA9+2ROOnsObj8Zy3sdBQdsO5zW+Aq5VNFOZUcN
LAjcAyN8MtGrP6gAkTqP8//9vi+8e1Hu99+q1d25CK06R7azh2E1S4cZ7jNrPF3D
zoAadEj9M3+di8u1jSRiI2PsliJsQAfc4WXMtc0E+MuNw6OzVmy1F8gkkSRXFyrn
BzG7hn18xECUu/+helXVient8XIrxHLx+urVWC3JTv2eIS4MSlv24slHRJw5Y9Tu
V+mn0tWjPQX8HYQ87v3NOqkCvZ50zrL/natvSjrz6BlR8IzhXtQrK3vQcseERgpW
LUDC2c21n/ECU/0NifpLkdxbP5jZ9A2ixd8YqC7OhVv34ibLhChWDGMvj/XWZo6f
3Km3DiGVqT3GHmMgaE9TPpGDZ0LhthJU6rZSKnSFAIZydt14fBi+vTLM/xXVGBl/
FUW499297gSYcjd2Fsai3CfZgVX4oXfqXF7hfwrYI8dyGlfjmgi8OZAGwtLvUMqa
1EIUQ+lf8FfrgxW9xCx1677VIN7MDmb0ytB1Lkl+VAQOacbhkbk0Q5Kqz4OdXr3B
F5qN+IBoo87ZsjFYzmcL0iIo8oPrd6iMqXxCzN2dO5BeFSu262vFXl3U9OhHFwzM
yyKexCg2fMgl7oT4OVmPEod28CfHWkJ/tb9WENOaIUUsCvUAZB975rUJnTZSdPmh
R2ro1S9PtkE49O2rWvjvvEDeJqV81fX1OEvTB/iijTuQSffQlCzoolnA8Dse479y
doN6BATc7YtLrlZ+T931MMGeWqSkNy4NW91x+x7iEYRK/c87okTfY4v8TfA8qX6f
duVJC0M+N1Uhvg6v5WWLIIeFqT9boTa+4Z1eEKjwnxAuTfrJwJP9yW7uyS9wgn9+
pYS9AGgKfc3pa/foi6aYFAjBbI9EqMp5KnI2Cg75/fV3HnQN2U3UKVDq6Ly9HOlu
ZC8qM0rqFRcKm5qnZAwW/B5+fc7RMznoAgcOuMmcAtG8AHCwuyqAvFo2OrOkE3aE
8Ld01PDOpWvFuTQkzcD9mQU67JJ/5Iv2otRI0MrKxf1z7A9H9q54VumyV3giWYqb
zYGscR3ha5jjoLhOnDsFTe3p72GbvKjO70dUyNHmmmQD3PdN4TY2iEx+9bxxijMA
K0KJV9ZDE7zmSZOvG+Ksh/JGaZNlG0LFCFXEIlX2M+/kqtpJhWEVVQxXzJ/aEr2v
QogirUXPqWbQ+yw5NSngZbzDKwtOaN2Jop6OXBz9BR8t6UXcgCy6Xu2Ano27n/pB
8z7tSuVLhTTYSx2cAHo2cWdYKE1UsR3ibPU6h/nUF7KcDQs11FJcIEBSFrggYGtA
rXbS95Z7zFgtiZxyhAHSVjuf9wZ1MAYUvBS+HxLtCGQ+e7W6SpymEUS8V4hCpwLY
KgE2hzHz3rM51g0gu1lFVgf+xRzoFd9c9u2VFZJqAiJAHRkH+LwkkZDHkCT1shpA
sDN+osIbu+Yd7hJUu2G2RY1LKuZN24spBbWnD1V2dxM/zqligrnFmPFuW7GsiTuY
MIHx01Kchr4jSRuFf1AMBooqdhKOEMHRW+i0l6es/WH76H96ZDf75ih5Mm+iOJaB
h8JvTNHyS0gjx8mxBl+vnmdqVXjyEAY7v69fwU+QVMAtvragBbLZgUjazJNrDKlw
fFvQdzrt0nJOc3nUaymG3IVY6coEwagV0N0kM2Xfu/UFL8cuI5r05ojI3NUzf+3o
8PQedh9OFmqh1N0xONc+Ht3DAgeTGXI94fSVK99n+ASO4vfUbSA0ZeH2yxlpiDD/
ExGxQXcqUTYjlrzkKgDBwLV2KN457rW+fti/SdUGv5azhOPld/9jOHUzDbDSLhFl
IUanW5jA7O9FSLmDPdklSwihwE8m7vGzYuAYJQ4EyTjd5Lh+RA7pB5O7dlvMBHPG
enom+VgLOJK1z3CVmrBX+QEEhEOf+HAi5TU4HjVY7ATJU4dViDMakIPf0rBp0ket
1QfyOUMRREozuKdaApRdVeRCCcM965p9nwU2cI3xl4QnhQIPgEL1kl2smbn/d0/s
/UrAmFFkKE8mWfWjL4cCbq2z+D5IzZ6rK7bys1ANYVK0XLX0oLWqLb3+vjvWvxbf
AiNJAPAvyyCg1fnTh5zjywNdajM+v6xCpFYXQHEypoV6VUa+QkUwBgQmOpbLFg1+
5i9gHqLGZlhChSSGHE8TKzqrgvD/mwN/DLs6cAekSFQEUCBTQpuTCRLzOjRtRUQ/
6wfp/xSpK/eou+hUC7y43g8qvxIDPbNNx341jzer43Z1cRSWTbXiLhJbF4FHguZq
0AIvGehNk0ntZy8uToS4lUC0XWesvCoKZkObL7vzmWr9NmDD0fc1dbqlY7nd/7WZ
F5guxXNlpPZYHZyKv0b/jZALBt0O/OIkcz9IA3VjuV4XqI0Knq35X3faFiBVKpYV
6w+yNJyND5FIsLwsdojCBqyt4qaYNHvhYn84fFCsvJoC3Kglx90yUrqAGfXJ8x0G
CsWtARiV2ZwMdvH2DE8JV1ZK+ihpky4oCov4Vtb+lCcBTTrVAgZi8arrDDwNN7y7
Vz/XIS4VTwOnMmYOX74obVLKsk2OZrSI9GtD6y31SAsJudHv9ZAQB3XNfebdxOCn
85ymlFxxkitBD+yG/CdfDifIfug0i6ADmGkc7yDWuY/xq9QehRhTIfxPASmCcwjp
c1Y2duwvAsci2rwnxmUU+GNInW1UFFw02ehTC85WB2J/lpYNaBsmxD8vBp5zb+xA
o5sCDPL3njuZQs5TR+6cZ4TbDsj4d6dV8qXMp8Pqiy15BgN8KKjIT6cD55dxYjnu
ZxRH0RibkIXpCXAM2ilG1Hf3w+JLlmEbCYTrcHQjfMsgZKmumWDn36gX0y+X0byr
3PQeDL18UGPa4hkqh+EZlHKua42g4ETQudZJHqLlXNblTCejBZ1BMoMsc/4DBpXi
qDEFSuknTi0veEUVSHP7YnmnTG/GYV+C8HM3B28gsT+R26xNeq6T0zUgeFhFkC7K
IdMEdqf+raQMunZJaYVePEQ9er/nJMDHM0JqfU8TLuy9BbFXaAnxCI3Us3eGb2fk
lPEWHpl1riPDSM1/qPqjB5F/YGdFmo8IgESFE7i8OiVN9WIfj5T119FNP/uqolhq
GdI4WDL7OIVia02g+W9ebDhHm2R9116XOz8l/62L4MWYHKL0rsHNW+wn9sI4GFHw
3WCpPQPaJpq8H9Hrd+a3rju4HQWldBVOjoV0kwuKYRfA7uM/PIJcIIzMV5AiUZeX
fQR10DEi/dMjkNKccRxE2pIY9StPC3+IsPVHW9hupmdOOHjYcHBGXSEZB1AtSraq
RGz6nc4nC33fnKW2IXtJLzfFu6iuptzlKqwure4RsneRmPoSanZ2btQC7L5/+jqr
Q3CpXrd67PnAMBd4Eu3jJfAVVoulspRgBjztpphna5szPBu2V//g8yGtroAndLVU
WkSJ4e3ZCDSOuoH6b5XHtlDNSvu2XY9JmDyr27jBuz8Of92YneB0oCyE/c85nGEe
ZtKcTKhL/6xwYsPt9UFNcCYja+y3hhhB+ZrDFH3qYpzxZ35f1gfq2C9Ak0hYwqQ5
y9MJjonJ1q+a/uF3OmxDhoO5mFUZebmhr+fkwl/wmpImgRlMaySGT3GmkF9wZwGn
G6EaQjJpsXKaydQUtbRV6ynqjHXRh7XP3gyiQRFOloq6z3YQrK8DFNk7v/Kt3Hxb
w687WtbEKrmg7PiwfRgNjO3bDdtGKnjaf0CsPlMWdIJcEAVE23CHpkl7ttpMH39N
X7LmDP4MsSjFRzh4yI95jzxukFn9FCRD9WOjuFT5pVs10hAuKNUHGvl4CarPdK1e
mUfTgUInh+Jm/oIDAyGvNZRuZqVuReCSFaArBptf9i0sRd3aF0KHVhMezD8kl47H
9lmTJTU+TMUT7RG1kuD7L1L9EGufZouyK8UPFxuSXfF/YQZyL2W7kE8/MMSeOrFd
Cv7w6h36dd+pOkxGWI49WaZoP2AmmAHJndOnceDThR0/CisB4oaH4s+25Eeb0gOV
vR8xMwvEMZWNtyodJwsocm3/+s6m++DNcS43XpT4HAXhwjQDbc3AhLLNxZxAFeIH
gDX3ZNUvv8UEiHv3TkD9Ui+TJEQX3uVtH1rddWsM2/DWW6aCs0/1bMl6vLL/G/PK
08ScgWSgPpuz3cxxYlOMQnGeAxcEsUUSyIcSFr2AVrn3Yj+JOYOYTc/Nlzh+/Hjf
Y3bK6XA6KVP6HLn8F8dIx4D3UqG+XKR3aMyiHITQ2rkgJHD7pkihd71gwuv9sdYh
F8C8mPUWBEQplcTRRAYMRZ6ca9z8RQaRr4NcA+K82HPfELl6zSqe/gIX+Wx0ZV+d
lmWJG9rT0IC7p0oUkUapve4x/6eCQzdmcRv6PT77E2JlRDaTKu56+xizQDXOg7sN
3+Od5XCHspiR45mm+yodBTTCEYCETiw4UxK5EWhdtfLQRJjh54sh7BmaSKQ+SwGd
AT8mnkfghDTehoXsAZMf6SZn0MbdMShsUY/o9xOnUbGZFH34l9ockls5mZuY98AV
kQMNmBseQmgJiyfGalmDH41kBDDwvls3hrRDFYlB8aZ9u6Xc21+3z9RU3GN2b8T1
lpem34sYsa+3bcJj3FeMUKuwG1c3+auaOC/7TEI6/2CVZEQ3IDpTiKdiT5ax+V5j
MaxdICPXsCarcKkRzi4lVot744wzX63e7xpLZXWeUZd/BbuSvixg9QZFy5/L7tqD
A2LpDG1CYAlbQJPZpwvDgbohqpM3irhQ6oIIiD4bYe6ptcrz2xPdXe1YVgQ4i/mS
Ti4YhKQuhYxaJ5685hezPMPZrPbjkiWx1khe1aFOfFreWFVzUy4idle4Es914RGN
9I2qnwvUYM2hsGqrfTl1WMvH1cT0OOmdYCHn1t31KcP9FeaYru+38cggkL3Sha1v
BSEWVqZS5SJKvan4SgsVEhFJIXYyTslttsxCjV77oBDHzyMtaPez8Oi1vUmc7nBg
uvSUt2BP71aP6dLG1L2LkmUlpUIPXXKLGraK2JENLOYc562NRxiWOeK7UIJ+00+3
7QEA/C6V7aGX8CrQKJHyEnb2hJXl+41/8s3uV7OVAG/tYPHs54/i7eTUYQ61UzVH
7oh/f41iqrbIl1180D2JiBl0b/4YuXamyMUeiX16caTT8STw5r+uwRy7q9D4P9kU
8nSKH0AOwZ9qA8s2+dBxb9X7dTamdv9RxktJheMXrJbk9zJKcO1bu9nAGasPfJNY
zfzEkEOn/NahLQEKqz++vaN5KiX2N8DH6R67MLQabwdZnWPhv66SY0JvcIH3/Xmr
10EPi4qwNe6QvmEu0frPwxwm++1aeUPTG7OGrgY/ZZVMxz5ydJcjFU6JLtXPZQmH
BzC6JJDxC7ArCuPi9DoKL7OB1rQKj0kJPbYvSbXqokMpvwLAE6TjvPioJubYvc03
2GwwzU9K7ir8C6GIsOzBsQ7crEot1iGi/q/wFnht4GrYTXVcsSl+HkBBQHqdeFmJ
stoZ6cpc7RZTOB2xhIB5hMQvUsRUB65mHy2Wbb3VS/cItkJDWRvjz7mKwqKT2k+b
el+XYWjB1dVFS68fzETo3+40V1qVbfc5ZOcAsLOkkOuXrYnIf7vwGtJ5QHoSFfYg
16BMof8b5ybxNTjBBGGc/SbXk9SokgVWYTS58hi5r0rd8QVIrgq2kLXZjif8bu5Z
KNIr20O8YLTvPbZrupfVE8wU0Ufxnq7ex+gPN3IsXa0CFYFmyLFR4Biqe6EU5S6i
ZthtmhU3S9EVnpymmRZVECKyN1aHI7sMqN+gWyvZJGs231fldiGunFN615Anl2cL
HoxGF6ksnHGxUodboOrdKx+vinB/Xww5PXCKg9bi2FPTJj8U//lGXVf8JOM/td4L
gqPy31Mrdpx0ymPzed7gEKTy5HFoES7iwRNkWOPZBPNvB+iPixYnxUDCG26L5/MT
IzQcexohigKZ9wp+JKoybdXzJzcf9vZrVOOZXBT/YkBTFqDq0bAwnM1tIriWZf6i
I5YeEhCgkcNNsz42SRjTMq1VpfrTSh+WzDrDaurGf8Fd1KwWLlGUBAmuvaXyn2lF
cw1nwaSt1E5er5lsfXNOWObX402cuOo94Slet1kBBP2iSTLqTOSIJ1hUrLuQGeIw
g/xkXVOxAG1XOfN83yG0WV+xomjeQRYsdOtyZJuTufTfPXnINeAHylcvM9pPYS2I
YDdgx5/duorsrD2CocMqcWKHjLB5vRZOgHsa5xNdjdjyc1ixGpvIYWxtnZ/M7+iR
K5IPzcQ68YQreD89EaHUsfsdJqm9wlg7ni0xj5oLZ58BadIMZZxc2lGSCVU+8BjV
cLk7FGjMBchKubkVLVpTmv9J/6oJ4iJZDjSlNHe0q/HmtuzV+7VUD3RG4F8qgHCe
ZiAH8VVSLbwwvyotasRslERql972YauC1mvyHLIxnhxecj+fIF9EU7n5ob2WDKIb
jym9Dvg1VJrQ71rpqq2T2+flnjDLHW8fL9dVoqCN3JjYORw3b5RcZWLFw67yHBSq
Km/pcz63lKcc5/nF1AOabfr7ILq6KF3Cn3I8pTflfBy17NIhdpL1DPPQroe1v74u
0D2xIR9reLgeFgshDuR2ZyQLWvEaiUEpiM/mLORDiP/gxtJwe9KhR0YT0r+r34Z4
6hn5UoRCriCklOyfxWNjTHRiN97zzab+1SBHRQ+/nuzAU5K4jY+hUCYvTu15GEVr
nVfXaTlIcxmP9bwD227riyN2+9L6CZkcP+zyXuyu8uXYkWUM9+hZeKBdg3Eevy+u
QCyMAxL6oDPNBsXqVL1MaJp06Iky8SjmSapxZG70KmxPAlVSLQGdmVITCQH7cQXs
+W98T7HWxj0IYcARW0YGDlgRIovGtrPcQzxy5YibjRJ5Wh/V6rwwcMZhdIvhB3Zv
K7UhPfl1PCnQTlbtefqk7N9XQ+ktWgy1gqScYLKsyvF7nYX2OZvn2G18jpipARLH
jinmLdNbJcCZOBfwKXayg7J226SXxCznNnzJxzrWh9gI+t5TeFoLkAFZFl9luNOd
Gg9LRP/Ips5WHniEEoE52HcNMRCU7IeTjCCJi4sx0Q+7qaTVEUZsg85iXp5d+yiy
a0rVsdUxHNCMnSA31tU4z9SroVdxeypHH+dtfonU3GS465v0wPnarIYIQV14Tinn
6KgY1t5fOGLWsc7EQkfSxp3PhzpNtYQjqkK7BPCmbLmdmthD0BlrkuNriXa+XlZJ
UwR8fYbvdP9x2DhYRasixEiabM8pFqqYGbkIC25lNI7YNfqutjI6E3OasP6y0v57
+hEVZNTT1icD+lyPOJG6lMQrTjBcvPjcMfulDkXpxWF/66ExlQR7h1ofLjm77k2+
SSeyX1BQivoYN/Bs9m2uq2fL71xD82xHFiWyXBuoCj0QIMjmp1Ddif+eD7PBd32u
lIdArVVOiAxk2YyWEamxU4fwS3iPAI4aCQ4NZLW/Hv+MaN+P2o1lm3I8Y0SSIN/r
5rFgsIGcHHGLgSW3r8Wg277OccB8ixnj4S5qyUQH2vU4RpfRqUXQrK8Dx2O+HNKv
E11I9gehrnZH+UYwZXoSUdpjZ/RVXB+tT1LVgVB19XK6sotGEWaIIJ25CfZXh4UN
RJhxj94Gd0rndnuwnrsvRVrWNjsY4OEtHlaEIgk9RbJ+fYRrgcmtroD5X2bMNa6a
tUmdYvRi1VhAUa6PQjUZHrFuF15ZszLF0yFrptycAnER1wNodaNt0ssCMq9kSz1K
6lpAj+5fuzciMU1QVxlgdI6d9I30bxeSCvVWnADAEjAIajq7BdQ8kThTS/V46dtB
crwd+lu75Q+3t6tVGF3l6z7ZVAc4q4v2vcSAkEWCt81Kt3ZbnVMxKpO+0/1k4qFM
rlf/ae7tbWEd+ZI6HxMTzzE9SanW5aLAaTfPh3wE10jC1F1kmmO8begZfwar/ntg
Dx31wv2LJaiY+dD5YBs++A0olLcNoXmBLgIIrveaCr7BVQVNcDVUWkhvFgxoxkBo
4Tr38OidG2TH2sw1NjfAiIIGBSkUTbq8zKswFqH35Gzsg3dIcu6XXWsEEPyQjT8o
rkaTw8KdZARIHyjURQX/SF1YWVcTo08puK8P/Tsp36gwnhURzVKVGIgRWejTo0qQ
qqHiEEm6OZkwPTjQuXrGGIFeoFRHkSe6rfRo5i/PVcVU1CJcXfLI3ljE1ptce0gT
ZKx3A9zmWiKJfW2DSbqHFFXGTjz8s6a1yzl6hfdXsW/oEOrznmtpEEg7VEKOLqCa
XYU7qdDY8GQSLqYss6wX7zotSY5NBwuSVoSOOofVaV5lltuNqfVI2ORCMPm86GIB
wAv9ZW7FGx/mi2IK4Vd0QQD+scg9rp1qZwDB7eOK65hn7hoySjdWU7IFTDK/jM0c
6kdW8bONdKq5GAsz8PFPfGsiyzTlhNw136v6bdOntWdWp4+lozthDAbkLlMPZryo
yPwVG/smFv3ZlD/1JbvxjdPAsxC7wHxk9QxRm4jjkih4iTFLCNJaj8+uQAonvxAW
v6ESW0A0MOxVMK2xV976P0T1+VciLDvFtaWYL9Gk3J1s1NXub4n3mFPGaFn5/xfL
ahnzM1ZF4TQmL1NzVhnIdpSu23Vu6Qk5XlfXIMMy8E6Xbs9aHdSMLxcHPmqX568R
XS4U+U97FwKnz1zoQ57JcjytWHnZkGKWD5eGh5+trAGiSszY/6nVvMuavG0z+yjw
c15cUJGfOxYm4AgKbQd4U0qsoMGJ4r4Xrc3os9db6LsRHDc/YqNpIng27mXwacS+
Tdquyah/bcBUUry746PXEOZgdUVNDgNkyyjGUPK/6dQARjCqx/YactsUR1hlP6Tq
B9ALuywLEc4vIVN0GLwXumL49q/DcQR9O/P5UJ+HvVC6xuEx+9ETzNBfPI7nE/uV
jGNlC54tWVBO+xsEwe+vP0rkCeoVX2sxeaGqE0cuZgvEZAj3WXn4O3ZkiNVhBlAe
RAq1q2STTRN4B1yRnz31mnKbQwVpV9UD67AUn7ufr4BxaxL4dd3IUXggMVYgisF1
lRO2totB1riN59KYcqlcTlyMJfWT93JuKJsgTiPAWzyC+8pMvUfD4XcFe44MvuV1
w2c2lDFxGhS1p1hAa9g90nfBIXe/NNvm3hJzBd/IpeoeBbS+WWHcs8NFSEkauU3a
ZYwzZJRZ9kDlEVS9g0CxicsXxFTpD2t9XFtjEFp47RCoAj+7C8E264B4/xj/sSWp
NdVRvUF8dqQJLXPa6z7vd/IyV5fvOV3ckmeEYe5L8G9UgLfyy/BwnJnz/TaMkpQc
mLW1BAeMwvnObU4C2/gEBi7++u03kLYrX8BVRipjlrrBl06md9yOguPDKuBrCrfr
i1lhB6YAu3k9fr0Ul0ppgnNcmAJME7q85OWh1OcQCf1AR90/t43+TQtyFikaXNKS
kVrgVc0NUS06smqAClNLTYzWf1zN4iut7XdWefqBotvoYXwb/cNLs2brCbOiJ1i+
Svyj5TZ03xXjWLGQ7tDoJKsYap+Gd3ArOsoUWdwSAOUgtOr9hssFxrJjvw6TwgTu
Y37+K9kXLg9f3RLlbySQ2o2ONfRhfs91+BXYMH0cPPUuUa+QDMzknpObc6nT9x+Q
pshJU10ndbsYSEgNgKW3tTy5SQ2+ni/iRNtKlt8ESj8r0mEl8BNyu1HAhjI3u/Zm
cECR8Mho8hXrcwk+UrDKSXW0+ICucLTFWsm6FhPQgxq//+LUr9t72TRpA+zSPvTk
ESa60QumYT80RGmlRlHlT05T7VVwa19cAYBUseNGRc4wvyfHjvzaxFZalz6YTEF8
04T1c28KSrUqfbwZ0culu/PQN48iUvzz+9JYI5n8m6Fe/rR7uEzNHNtIpqMBIWI8
wQxdPofwchVlozLdeB2l80Gq8Pu4auUKisRbaUypROl61hXlI0pPAf8SdxJW9R1c
JB5eCQdAz3noaIPIvx0HOdNP+hm4DKhtJ5AM+eArZrndZgYbNOXGAaffy0cl3v3M
XJPIcqnkNu0QxG9FQL9MRiUXnoG2P2PoUqnaVImaPZvh3gzA9AdwAbnbRj/BgKnk
tRKBMckn93lg5Ye1s82nMevnANFfyWbnKLhSTSqjvIINfNul0ZAavboqMzpY85PP
dTKJeevoYWNAmqn7+abhjiy1yACUjAqC0WlRd2lY0qNSSJ8OOQ6b4L6RefBZ+Bhm
ziIs9JAX4+2yPlCpVAaZ69EuOrupN73d8jL4u54JejHLlTZVipFQbSJnv3FoepR3
cspBECfdfmuiTC3SlJw8KV7yaBLv/t+Coe4an7vXZL6AHvn+Phs4KlmQGD9WZvaJ
44gWGtBA7Y872s/IdS8J9c8/J3jhJ0Id7MhHFBr2j8ZK9H8/BnEVbiJxeVCDVDsk
lmHwlLy6gqfF1MhahLcOMR1F5MljeRTwRonBIaVKNbE7unIYsM4IXzIgyDdSgzJx
ZFuMCjFEpM77nq1zsuGUzAOpqBBUrfjbznyYt0mI5f4gFfhfBmQtgdg4QtzJyvwk
J7mBHalRF5IY38oENjBeER4DljdPrTIBSrc4wAJFHy3om9HdjDwZsmALWyGOG26M
Qwe+6g2pqcCRPhBWrkfNmbUJoQnIC5PpdkjZiPvf+1P8mYOiNQuPEpJZ7g+3/MOW
nT95UxY02lUPBPJGEFCgGSNzT25MK6qz+B026SIJS0ntHrjjamUA9/lPGTAHTrum
rXJH2GQWaWwQcW8sptmFcZyj9eP9EMG22Q+TqPKtbP/MhyRtntSdMjwmhJuClYUU
dJMQ5HHUzeS5ef7611rV8M4v7vgDLf5UvLkxXOs64TTqI7ee7ycNI4V/nE72GynS
fpWEXaxW00h9QB/6Mim1GsBNRmrEFU3UjMs0PrhIqmmh4rLSBzkbKA8Ct6osDTD0
yMY5t/qtt8S/Eoo65biQjxoNqkaEB8XMfi/ODEFGNMrQU9CTlHaXK+0wY3iwHUHs
SENOE6eCgXZbCxtw60GcgeGC4djQ9ks+cXv7Ocy9ZuhOz6HNOT72M/U80oY4Tgj/
MPeTB3j6Ro5qL0RN12O/4T7gGHxpL5X13WL+mRc/DEZb9dWJ22EEjr/M8FxNnirM
30WaB8V/oFvdfQQLaujcHcQC1XTOR3rZ3fSdUxTmJKSxa1PJrWoY8TS3B0iNWZnq
rF/cW2PBhdZEkw2H248/Xt6xHzSXe5cY+jQhz3Vlc6KuEBCXe9YuT6rvcVdSSLoJ
xzFa8+Lw0ZK8NMmetnPK1J+KpXvXMoEXypWxgUKGkg4jrSb4Ym+akwN7mlvSCw0o
kTimmBdp2hjokGSzKBgYBMPNMsBKEQDc5QGe0JWADEkpqcGsJBQ6vZkSz8yiHppE
GHM0q5B59JyIjz1mOBbgpEtTUprXRht+LNmReSMuYlWeXBJQ7TAsu4dI4NhuI9Vi
7z8r4IjaDXMK4T4gEJsuME6NNLm5ZTo/ngzEZ9XI5IR2+eM6jLRlKLuQMkGhly9Z
kErGiTMiIkWJDpjgGx5aMH+PsKKQnKt3Z/jhdUOSwSs/bDSQreshdp2qZttnMEE0
tFtV9OeGuU2iySN6ryyGDm3L5X4jGFzRNuDRpwF7VjlodE5YpJjVzTPo23eLYQ7w
NLj6iDdU8oTQsDPgvQiIugaBJsIiz3pWY5Z6uPEyDZnsiF5ohjctQ0J4c6gRObS4
OMFWBKWnxaurfVx8n4xieOyad5aGi0F4b9Ri1Ag86FKLDlxkGCej8rxhHtWVfsLf
mDkmlNT+xnOWIo98hVyIbB/78hhIOQF2Y3F6N2UQ3MZN48ZF+Tq7FKO9Y3n+FNF8
BCCNYgH5QCU3hIVs1fZEZhsmI5g1oS2H0hu7Znvi73UAmeAUbLuwRFW3iH2E1dAE
CHGR85pjiGNjDNd8K4JExfayCfXu9cDNL7zq+HnfqGzs6pHBybVLQ0ZBTWJX9Ord
lX8XfaVt9HkqUNl+n8juwiY3/IqeTp53dl7HIGxrifvWsbK2NPEVLwdcLz3id3wU
1GCRRmscvSFCeVIxD1t2DsHeFPHeycGA89DC0gx7D9RfIou5MTPdEEEnibipCPRR
DYSE7eyksYDWr/9WjAzohkDI0IvZ+f8RU41Nw1WJDEP+IDavAoUEJuW8C4xZZFZH
b4MDQqA1AJlq5oszB7c3bq2b5/56t2bYaSQ9kRL6ryHj2gIw3jdEJRKOsl+YkRTn
pGBBwlgcBi382+Aesw17clzWEOsCsDv2kLEiax5B/XtubJnDb+SpyG3SVycE55Mf
R2tcqm2GNggbkj1pvKpinmlpGA5Whlic3riPx2MGOcYZQSRrJ9tQZYtKlhUhAUp+
cy6MZOi25mnLftq/CELIr6Egbcvik2dkqH+ExOL/PXOxNswsraINMM5+fodN5HdV
/2rn65LFFrvHedsh9bas8DAJEYKGui82Jb9zBWf0pjfzyfjjDxzc5/JX0XRM4rxj
bd0LLjPE6xc1Dh+NYAchRDcoOfpV30G1AUP7dEfnyVWOmrOh82n74thqBaKjL+5q
n7+97ZdWoZDS4F1KxOxsWCDcmXtk+EUynPDVb0v08CmHtahfDyFkYIdo3i0bnmhE
RCqX9fSUkJnfos5mxS5GRWCJ4TC6MQqN6WkL5YkisBhtcC48IX2VbJDDDFhvxWIc
vD3m43zrXvrGvrp4tG1O19iuGPuch0V+Ia6r4Cm8rSMw6qQmlVK0FZ2jmL1f6Kvl
9bU1It7ng/x+Elo/0WAfimx2VY7ffV8w/LuYVjZMuIHljJ99hIQ2yeSP80YjyYZJ
bqNYYAlJA+yXTwnibiCI0p+YRs+1V34wbFrd9WBVsup90i+Gsj1ICzfvQ4hVo4OQ
oPWec6hw3Vgk8n4Xtx2Ik7EqhDUNveXRRF9PVkXS+ZPxUJaPznwOINBRB/PgR3Tu
wKxlGhtuPsgjKNDs4O/Q0aVAIEtI3W7vt2R7ej44QzvhtdzuHUYaHEuPua7i5A1Y
O/WbIs5z2ABp4qiEERNEpXb4sA1dyLraH3uGI2qSg+IxMqvMSRm8Qpxqdv6IwIIE
MaVYpuE9j9ch5XDDrdgRzSMUWcUpOhcvXmy6j346nc79Ip5LMN8iAC0fL9BAssOr
e2yl01B0VEDstdxaR6Xd2yK1l97YnfFPInSVQCg8RveCvHTmbbWu6+4WhgG0aPoN
LcHJSX+T69GhpCfDGbDj2eRlgV2M7kFSPoeytRQRdJtaZjC2W0HIjySJQtQfICZq
G0dYD0wtbFkmgK3fnSrGpANTsLxTOPIQGaXYjGCAgy3F6fqscsDNRThThgSKFt9u
DsZI4btUJtivtDtG1qQVVx04yDF7DsPKADgzElkUpqw2b1Vz1qD3RICLLO+WrQls
mhvLazGdbnAHNM69YmSbmb1r2GXfWf3e77K8lzDMYbYv4PhXCYlIO0f/m3tuyPNe
2xgBKAEDflaLpmPVhtnjG0AHvd828qRPcMVhO2+KiBmCb53crlYw7Wirt0wUVHyB
xCBrRv7u4rs53bSvZuDMevZA7x+u8R7qTFw99x9fvxqOuVrXGjKSauUq4+EHd9k8
dOm0u93Kk5f+54ZI3I0MOdc0G0v8TVutHzYwcatdHYvE8+oCodqBklf4sfAqoXnH
eXdjQbynWyGaRa+QOXa9XCzZ429GWqa1K+xTXWk0m5xn5dtWnPaS2bmpBh2PmD4i
I80dLlyQZ/bHzG50m/ac7g3nqMsGheqZt2+ep0pBdItRxbOhgjT/CfzHuWIRMRex
hNtA6k278RciSXXpvwg3z82urxtuZ9Sh1+568PiZZc2UgrsblwngmBfJfCZgI8J4
v7H/icuQfhmbNGbhOWLs9TSGBkmzz8Sw+IJsWRMoNbUqIv2uiAy9jvRM+qOLbuAK
GnKCTq71Zm3oYvVSrhgBSRlwsInDROax2M0xpX4683vaRUZyzeJAmSXSwf2AWnSN
mJonTK+JFc5K0BVKfs67nh/ogJQy5tcZAHHfsXr+W8wytc3uUXNXR2N0qKYWETY/
b/kYBEcQ+Pp1G+BuTKQOAS5JnYRWjKrU2s6vPrVeZd6bSHlBdsyiZZd4uJERfPvp
q/GmTb+74Y33KH5WoxGiDs+1bybiGHyixbXspmnIUZvkp9E0z5c+33+z21+RqMjh
NM6vl48ORmRM++1WPb5+GMxqrgscFbloerua8QufINsN86N+Ajov0uYACs2aX7L9
FwmJbBIWzcxq9Dayf5yQikxic9WC5icBR2U8lFpW/Wz+c3w6JjWNpkgJqUYAR3E2
vKD71pKa5nVlYZOjpsLZ9AaVIm4OqD6v9tT0fNFOpWeAse+2rOXsSrsABdNnY1JZ
utVoklo4sEwZulowFBijyaiGuShU0VxFrrd7zKRbLF7tYyPDRKd7Q5W/WQgBUbTP
IrYYFTrFEOOpEVYjPTJD+RXmbm+y4GJf5oRonmEwTM3htQxKRwjxroIYH5Yw7xmI
+nIjfpv+GnDkDLZqLCwphMQ4BD8HpELAej5mlRpSOVLseOJ77VSsRjqQ/qzJK2qH
fgekHiBZfLdQEADo0T6UvfcwErKppnlkFqZzsMyGUHqyIIJL04AmTEU+OPhUYLr1
xEeL5tL+jILdfx4D6FPXzfDpvGuxCi7RH2jfgd9N5NnLRzfd2F7/85XvN02TDezl
IGNp59XzP8/+1wusRB35zu8VhMsrctv8zTbdb26YRkLcED1Kbjgv5o1osNN6Vbfs
N4x1M1/vEgqe+7c223cvy3lCHES+YxUBRd6We+6+pbLhOkorz8g+OzCDsiDVpdiw
LmKFV7aQkuOXP2NXNfmD7n3Dlg4WTA8QA4lbqAqPl72dd7b/xzlLH5z/E2TGOIoV
pWcvqt9HsUNiw31RDtRDZQRxd2lYb6mJLFAFaQFAGKi/hxw8AdINKUh1Tam+iVLV
o7bD0E36tXdQ42VrxmkwGufjXMvrmOi9o12pALYVd4tb4jD4Ph6P4TNdOs2H956W
0JcRG5heNtnbXYY4mwQRnjSbu8h9bhobHn6BHeQz2eEAzf5Qo2dq7dAPP+hVwJ2d
EQsYfWBJtkk98f+ndrGan9m1IZup8MnQRrDsyeva2FB6J2ElCD1ciTYK9Vf4wfwT
ADr+R0obrNZs8ihKV7w0QqHaeeHtezi3d5hp+XHIaLSmtZcqfCxwlgwiFiNhdXeB
mMTjtEHEM9E6WNeEn4fXtXe3Nyrlb7Dm0SECXP8EUqS87wicBG+5hwTi7a1JKgDp
PCiWdBVct2ocywnU2BEP1zHl6PtXztl7NkkT48pC+nF8yvVW43XR19z3G4Wbu0VM
NL2lwcFHZ6pQuOGHq9iXwUEo2t417KK4wOXFNQvT0y2m+sUmG+wI2lra6+pH3bsq
mP2urIe9nh/Mywb3WpqU2jq1Ql5NYA639vnQxX+E4Sq+vHsBQdzCnLBEw5gYCz/f
eWh27IK7rGqydE3mjaNxqCyxHmnfnW7ikVxpJi4c+AOc5b2Ze3Ohsq/Ytcoz7Q9c
N4H8G+s+Lzo5JGxIwNLjqRXRuzQvg4swjoeQfPbEdSJqBUAkUZ1GVJwBbBeDxoKZ
LZXwdGWANv9s0Q/HJPmIxsuRjSGbdZvXxYb8XLBZBDwNs+ocfRfjEhlv3Ai5XrmH
8VNzWtmZ2FBFYYDikc9uGbPcceJ1iJq71tvH+5NjPmTxYZM7jpqfHbw3rDr+Zt9X
Zj3gMn02t0mQBhuQbBj+pcPXy4mwHkDBOvcPGhKfstReI/w0mhniRfeGNNHkE7CG
PH5X3RFtU4QXeM6Ly+phWat5+O9sHb6Juc5VlWWyBrqIku5yz4vyIFXRL5bRFLYW
+rr94usdhhe+CSgTkIgtjSv9dNwWIUgSGO8VeNIo5fL04DQWBraGu8KNkY83KrKq
7QdQqSIH/izgvaXJYwZhMDgw2v97J7PAKIgzd3998RMspiij4gKPqqtgufKIx7Yg
Do/8iLZeP8kzjTxtfBuyE85aRA9X0QCKd+JSM7m0L9uZlTlN+oQm8qFtlZ4OqVJT
FJAtQ8BB7wgO34Erf27wpBeFHOQ6NBi9oZP/lIA2jY9iQ85u0x+72OsnFA6Oo67v
u3+/oxBuGsuWsvrTRHIi2DSiCj+Y1+UfA6rAuct8pAC9QaL2+FSG1R3XuN/Ysr/N
BN4y/5LVlOXfvviJyS3EjFHkOfI8V1zNZZ8bsRg9spM+UrDSS48jqfVCvvBUPsuz
6nVopN7rwcSRcaZyocONBaJZ9a8Vz5b4JvRPXSpkczG7RwioxX+RzW9Fjzvn3FNP
4SNPCEmirQtgFQzW3TICly/D3uGWNoX64Ce+CEnvVuXV4FgTYYz9LWKJY1IKE/Pc
imRFjpjy1ZS/g1sbwraWPC07FNneAmkY6yWWE1+jB83VPU+2qAdatQ92/4uInOEr
jrZXHh0a1zU2mu90lmO6EAGkNMDp9Wq66ICzLF81yyuM4bhOlyIgyH5/FIfw92jE
KwIMAJ9UjDIstTCxbjBiO4ZMm06ofKvWVeerQv/P3dscrUAtJKDPRVS8lHv4+TkO
hZEq0Foz7sxkKay9pvtVZEcbWf+/dpLUpwZakD82dUxv0fGH0oRAIwrIcKp5M+w2
eIzrH3/RzImTEmeVTvanlTVuwFDJuzTkn/LDEvAnNSvTMw2MviUo/Yp3WkjbS401
39xVMd0DDatnmlSmG/c2pXuS9bXaSRDR3En+Ec3ijt11SpmGHFUu1UKd3klc7ru0
JW66w2TygGVdWcKT8ZGCHG2xftfWLKu2mVBwky4hv/7Lmud2b63wiBsg40cI40Lq
j8Rw2KhL/VO+qm5i87AGBQVxCVqMSHiR+6G8QcRABRYqYOhE8Dr6QBhBd2kO7qml
NY9B8aYFox6d+Vy01nb6k6wkejQed3WYBpMW4MbLYri13Eethf6ZklChLUoA4fLF
SvP5pSyRSOQMOBeqoAoQcrOBo68o6QeWny5rOAOWd3M98iiinZjjRp7JbhXtArox
9XEOUk2xapZMyIIrf1sCKazAgdvzf8oCsfa7KiXKnXZ+RzN7KJTLxgtE9kR974fA
2cwjLLdlEQrLd1pixERqqjXmMBbDI9s9eh7IwUCqKjDm9p8u4moGM5G+GMenxIkj
1sa75N7zXTwID1gH2btr/htE4krdAaE4kd8n7sG4PPDWsrgKiz07ciCxNMeKKXc6
22eOwsBYYEF0uFm9nilevFaZV9MHVEL2SUr3L8qoKo3yNzsFWYEv65DfitfK2KfB
sM98qL3jctev5qLzicr5jPb6SRERkGIF2ySNFpof3bDDxAi3gM0ao/3xTxA0Kh58
q7zZkPd2VrEUO5esxo81aXLE5orZVXdcRA3OhQpBll9p+8zmPnvFA4A4bYePf6kf
MUyF+c1o4Kh+31mlUyDJW0EEmCXb2IUznoZRA0x73aawEtEEGLlOsHif1hCwGSNp
Kcc9/rRkkqi0+8fKPOsyrK1UAFNuNXllYNAnq+CN1taKLztlDKff+871thCEvDAK
NReSBywgUdPjpYpn5bCpVb0GE77fldGWp90WoYq2bqCXsjhcgv8LjglqQzSt12E/
wz9f/BMvdfnjcEAgmxMepcHjpwaIcGJJ+nzzKrr8bobfJcAo5SbCIbbm8Dv9akZw
JDBnL5G+S9T+EfrAKzJdXERA0olMfm4v60/EFmdEpB2543xabraqQMmEcmSeBZ6C
rmlrNsaJ+x25ZzXgcoUgrYkLhQs0lu4TUZzsbuMn7ibEcdn4Po2d+xhP6/TvtYmK
YzZ+105ktWiZSa/PxKvK+3J+5hOeO/b2mk+40HqynSsyiaVaezmIYXiS1RqjWqNs
hvosZZQbEPZ3pDqrfg7SBXif2JAutnwmV3sO8TcDslNpQm/qGdWslM42UQLSfAP/
9qgaUBmViBgw5mJs4fK+kOFJLacclTV24OvYD1wwcbENUDZE9GuZ2+12kIVKxHNB
WLv/tkE18yOOrBwp0zLD4AvPjSDfV6NpnU718TkibYOKrMXX3nsBZQdAn2ML6Bbw
z9RNRHmtk9DIzRhVK8pYac3cCgkeXYdH3BWf1lGG9lKXdghNtgOR3n0k455OrGye
5rPWyXr2XRad5b5b5uGUEdtA/iOwAYGkeVmU6UruRhjpJGe//GC5otTe/a1MXT/v
bJ9bI88J+bTPWRVvjk122UgMWLGsIaMBtTQ3mf5VBpqmKc1Pf9MHmv75Q+w+nZSr
NgdI0BQFqyod1TPQUxepQP0/jfq/2RkxPXthfDVnQN/EOfWxsq1Ku4hfyL15JsBE
wP/gPb9FYU2q5OwobsR3gdc8uATKDeOgKotN0/hihk8WQRHJ5nETWAYgzI0AoDOe
ls4pr0K2f0uO/57oRxazbLA23z2LesZN0BkEsrGMEbM9XPMcbSFArlmSkpsuJOoJ
nuGA7dLc9izQ6v3OrpCgSSz08owpqsXTQQlZj2gDZn4s1NDp8HB463tJeoXAUDUL
vqPjUv8PiVQNy0jaaZOIf2WLtj9w3xsa5JpPq5WuCtAnjZKWliNvxoF6csWeR2Y+
m9Os2rEyiK1L4kki1yWPnWi7dbHFB3PwiwveyxsRIL+5Y8OtLwPGbKJyyeV+0auZ
mBdBUVTZv6aCeu9Rz5x2WPoOlIOlVUptam7u5lqNR6kOWS2JGzKxVW4F270QeInH
CBDkal5LONSKu0uC5A8GAo1+2Uht9fSzhAUd4ZdJefy+U3Y+T1lruIrBlPz1iGMc
du48aQEw4YeXGZU05F9YzEcXMuX4nm0FqeFrKknb0gontnJHJyKDaOxmcT3pMEz0
TnYuj2sLNRVMAjNZRv2h4cQoelq3O0BeJSwmItIBmpA6Ob0LtJld2n3oVMGswfFq
v7sC0/nxCFp0dkmv8PSibreggt0wMXAFq5J8BUxl1s5UOj5za/rBY2Nry8USbw9G
hXjjMLjiyZ7TTEAtXihVzIfu4VDqqM4DSZJTtiuaJPUWEF+rV0Qp8kT0vJN1N1v/
oozCu63lBuO/2mpipRJfHm3XFWImiDfZEJlPnlRzeYFTrIacqfljFpVrsuUGnFPO
ekH3ZkJZQT1x/GOwCUHO6xsyJYEJ5GEvhVbdQOJ3OuXnzz7d40aHGL9cezdhFJJl
jc20Z+IL7W0Grh+kZ0gNry0Z2+TvXQBE+uE0NnyN9yzrsQOINTssI8kPJ2x+x6+N
DshSVKMGjytDsWMyht+E6svdOw7KdDGYL6j+AZdJJ/iYTTEQXp60knajEWtkCimP
emOq8SURg8IQ6rpSCjZfRGp9T3juQn9R4Sy/oIMWyarl3zSA77tkJG3rYpjqdiE9
H8B0Vih4aPL9BdTJEfRwke9wyGpR/i7aK9RXYUBikXWuXRZoI2C7M57EAhBPvbPk
nllLP+udtr2Fw/EpfgRSqD9YKatWF6u3tG6CPSe5JaNgy+dHALd6AbuecTZ/zkfM
1WLJHUVgbqHw/bwd9GE0x274tigc7ewnWjwJGwB9szCQ8NnSeYlgYxj/RT2MytyQ
G3aG/4k1hGEJPHWVvPI4weSN8657KEFQonuik//NrVcDWqRiQLXHZtUftdwPBBrz
qGhWb+zl4Y0Y89gH01bhovpXQJcRGZtxbGazEh/hUV6++m0RF/KS1SdKEDs1hQjf
5TEe3NIKYEhww3AH8ZumtrWG/UCePEwht8YhbkRa7d9znEUB/9SIZ+DOB0BkDhe6
U2qv6QxCfPtZ5F1xs7Z56VfSejvmgaxHlEZq1yUEMzbVq3gNRvhUghih1TuDWk7C
RIjK945l9gut4kPWNV7iPdKtdMG56ebtydb1pZNe14qVL/wMTUOO8svgnUz0xh8/
PCcBMoFVoa5xFpopwuFZajnuM/G3EUbfqyvTur+l5n2ELmUK9PecHx51BMvlR30k
YkZStg+60FFggqwNs2/+NKyDovLgZ47wCCSH3JLOtnm+tfLDSZIYH0WaknW/ctf5
Febku3UKcMmzEw4VcCvh0txw8x84b1oHORHynSCdz/t+jo8PLtLInwCCay8Ys3Pl
2KD7FC3gsC6y88Erm/drQv81Tmg/ni68ltDH7WVnw2msuZwL/1Hw9z+aJ58qKukL
GIv6mn1ygXtIT2u7QQcbHudt1uRk0hitwmsBoFE+cevwf+z+N1v+A6+Px5qMaUxJ
410Zq6tEYNfWqUQvKVW7DcFjXbtgI/nnBVnrGkN/CFPv/r4Ylmb9K/BqjuiIMSPB
mVduIp5Nu3ySXk+pfUOFZg0HetHhdqrOmy7juT70VTqwQrK03eN/kN3mC942WZF+
UY3HfUefvll6ZV3x16MTrlJqSOO5zdEvFS2Uuz+/VBvSEhTHV/yRQXcxw+laVK14
r2fqdfUL+81VusjpsUwrUtBmTCKWpgSFCxu1muXC2S7B2K3CnaAs4df7d116ffYg
oHtRkZcSIGL2ZiWAfNoLGAb4arCQVNSVCJnHVrkCQWmfJuvC1qP2MhCpb51ABEo3
xdDAy3E5i/W8LRmYrKtHQG7PCNB2eN5Qm+9zvINpaOt+PQANZc6TxD5PCY7bVgT8
u/hwlc0QfmkBIeva5gD25MAILAhGJyZ281HFpdlOg8fn9wgm+lEIXNwvbX8bE4Qd
quOOvhOniPRbO3rnxd2qE5hjFhCV1ENd9xQS+fYaX7OAxHCaRjoPrzoWwYGG9tAN
Un4weFnCi93+jhf92kzX16GX1HZj6U6caRVpCqM8AuMydviucqSIEz15XqBW8Gjt
ENiOMs1LIV1wIRJ6pTRxDgQF7cJLqgACT3I3l2a2AIhNBiEk3s5IVmtomoOWFLgg
U2HDSn8itSYeVNlP//+XLv6bI+YTD8ZxLOZMdGjDASHIvOOtMsPGic/0m66yeY39
hlLOWeNSaXlFMwF3G42/OCaqsM3/0cQiOarXETMFCgDZ8qoEXmEQ9yB8HhOdnhw0
//XajDxOKLtc2Q32c+bjtjgGf/M93MQ8YcAHFPYII/HVh4wC5NgS0G76jPKzJGtM
5xelbxTlUtKW+6uFI+trgKMo7reVoZKbF+/omkrQIa05cl1CP9jbPbJEWNvysAn4
KvwRdk+DQR7AsNNyP2ISHLZCP6UekDxiRg7u3MBqrO3yFPjwCKMvRDYrbQJGKRCx
bXN9OYlmsylH6UENajmm9aK+koZg9i87jZK0mzm/bQ6Z/9+gD496G2RPwYw/VD/y
j5aZg5H9F/ortMQFGZvRUz7ZHmeHKWje6sttjdskbqgDFxKVXKMx0WwyfVEzMaRp
ea7rIYEHvo40C1HF9KvB249QNGHZ1ZhwDGfsEvj7vHoJKbQgqLyP8+cxT3f6XUvY
p+sKHjN3hwCarD15MCuiTvdC8Pj8cI65yUrm9wLyFdR35PYVWTbjnXANsszFq8RX
EtlpETgfeH0G5tpNPDY+xRn0Ni/Eek6e/xw3vUD2Udu5B8eB4J/5KEAzrTh+FaEQ
MY62exqO53YdDPm7tS/vRtEhq6UJH18k+j+NgJsTLTePPfjHfnI4Px9Cvq7P7plH
UoL0WqpDcQZQEevggten+lYpupT4rDC/ob16QxWdD1U5T5O7KRRDl5letY17W+GP
5Z9JQL9Py0mjA9W4Qv1Onritz74auaEC2wz7p+GmgDvibkMtnQJP8QLH0wiyiAMo
BOfzenGoyR7ftIsXTq+LJLs8veVko6HR6M7pYNpWFZEvGZBqFGCc30kaxqPl/vfT
0llp2UDnF+COMT2/OwZbiGad8J3+RUhQrBJamRkOibRJh+jr3hn/a7b3e/P9cA3j
/soIOJjwUKt3rdeMaGZwA4NDxL+nwIGAXr2Wkn+5ccYIhjLkXeDhJeHykhvM65AU
KjAFbPfR8Wc1UCs+tuoNdfOIxU5dQbEm5hGDBL+m67FWiDYzKj8O48vqk1c1/noz
jS5NelZPjExWWRTOFTsCJmDOJbSxD9XCjrozZPJq7Gt04+XMC9I+jMiRvtRfW4Q2
1LZ+uRSdXIe5uz3vh5xgekkf88NwgefgkoQD15L2eO+p/fD6My+qbrAefVwXTqLn
LeDIqS6vOP6xXKf9Xocx0ivlaCQuyjQrhLO9HbnFFs4OFJ0UnaSOVsuUjAdgI4Jq
yP7ODipHIf4uKtqYDOFpk6hEFWaFRYljFk0rEPldT8rBXXwKDWuSphye7VUJGRms
/WvvoeKG52hgLEg9cviR5V2IAzxodHpYiOGmct5SEPKBDxc8uWY0ywDbzIiqq4kU
Q8DvxSyVaIjnmFZPVnUybwNbb9r5q6+5Gza+8rDAVvKkBxYMactedAp12k7EMGwe
wMtzLp6GyVCygBeHv71oAPinPscEkQGql2kzpbK505LvUsdutBTkvAasxpVAhGvf
/ecGPKx2N1+MEes0R2VrF+Fr5Ek/9dezfTztKOfi/JBGcvtzzlQr5HNYknouwHds
7igDKcl9Cyhrmaa0Dazs06Ur4aHxcV6Zd12rJTiwy8F1S6VHjhE19m2ZoYt0KAKx
wYezXpQsxzjzxtKkMgtY4k4WGT6UukRJ8c5+w3Cx4hTQnJaA6AVOQPw3RU5kMNRa
Pl+woO7vECI7UvxG9BUK4yy3eklYtVAfsVBmJ67g0ZFfHdmtN50QMk3lNO7TyvWN
PKQ9HXvBA5/QEEUihkX2GHc0I72yHOu6Vc4WqC0LBuVifs9Lx5OABgkNP0h8NAKt
PCWnL2CA0t2qFgPUCCGy8kJWssLpv+DFg+ePVLelrXl3GhV480MssNqa0Jb/Yi62
NmgaNnG3X9sFhn4EuLX2Z0CYAMK68/1Qyl/C2Qg1/d5DSRzK+szbWFfvVexIQ+dY
Dof1J+JZ6xjL74DsN8NNqGwMKCmQuH/By+yOuBLbeI5HKLMsHDkEYWjBNgoumYkU
AClvNRsIPy2xUjxawl4OlhduAtz+qipLlk53PgfaT5PYqo+IuD5/qBAa1GZ47qvZ
jmVlQ3z4q7M4JuUJBqQH63qW3cvY6SdigeT9XbsXhAtHfDhdZqcyTzxIJ/2tKH2j
lenxNBL/EAxFyLLyh22Kflk6mG84j4aJY2qHM19DNTuMucEML4pKQ4EF5tmgheDB
mbkII4g1PhOgEsMOA8bXmoY6ECTtMIC7I+sqN+WuNWhow0zP/RyKp05eqKxqhDBH
4XnKRZBiP6kqyidVjR24fZPx8UQmyP2mYagJJHBWWjCqe+pwhMzjqQxM3OQOhYhM
ILOHAU5YtJuWQ2P7kkxemezkqpbwpMvHWesJdj2H/jympS0Ouh4PY27lmK8Mdbb8
U4nNoPYS3x9GzDjdKsYpQ0/FE9NEJaQe8r/gBSAyvisx4r3Sn1inJCVL7+zwMhhf
QfCl1xO4DHU4Yltis7IHfOnnTClg6qmDJDVEEsOwgBtPxwx9DKYW18vRV2zLMnXQ
shvl2ZdiTEnvqSB/JDRkdSSWZWwSZFRUkMR+OSGXGOeFxqyhAiilgkoITxNydibV
jCgM8yIXVbRs8i50jbMNcO1TqZJLtTBou0k5NqGKm+7KZU1wxE9+bPPgapxFgzw8
f+J7MxZ09jddvSYlWC0cLs056hvWUo78zHFHdgMjzuiW1sGWsdrEieDBqOGYXdzA
XR1hizLX0pYevj81Q56PF8oLfKCk+AkY+RCUekK8h/bK5PDFT2RhxY3Cq5IKLtPd
ERy2PzgPCfSb3JQLTTxLAgt+5kwJ20/+QVXPnaamRc8Xag2VeMBZzm8keFYt6MmW
pF8OxtOcDk63eMyYfixFI3efbg8UOUcpQR2mgu7VwscsN6JEpTT788v3Bx6JK8Cr
9fJ3jL2AAKJiws9g5oKvQv2P6i0CVJRTLT4YgCbMmllwYDzQmECNcXVvlm81dUdT
1p0WWdYXQH1/B045TIIQOkcQJYkUEYWxWXzdo2LqLwasquRAuPIMXwAnpsHGqPgJ
nNS/ksDXPPJC30+pmXt0u+HYWDePNpEFaZLazUPX4punFxDgVYaSyD6lIPFHMX/M
+zGkLxo8j+TdwwYmdb0SBv6UQtCYqVP518E2MTqwM578vbEnr+JM8D5jHd/NfXVF
H9asBkVDeQskWUqsaFLv4qi95FouTZSU7jgLJSKEkniRH/5xubs9yA1Pu33P1LLO
EOLfXNQdAKuiU0fXVH0DiIjzfZSZPyfFBLwG2iXBQjQGs5B7BxHHYlE4PCTSujJ5
zCe/xbOcw7aWIKZIJ81WVPHq/4Dgh5tkp/UEBPoy9LX9BU53+Qz/B0KC20oKOLja
0a5KhsOZtzDeWn8iPgMJ1Rbsc3wW/zZkBvsxWZm7Fx6Ye0CTWPd+HJE/67I2eDIC
dJOqBZYwjHLGg/CBOntVdJb2Ru6QqREHV03w7w6wsmiz5twilUwF8rvTlKkiWPt1
+9g6XRCD3CsoThMiGqfhDgrSmURbx3JqZbBEmMtjuycucHmlWDnMFihvr640N4O9
/9peqbwc+1/8A+3VshZypKpbueFFvWqaqgjWL3/atUlWc1wRGAmkmUwBdsfoV3Js
4+wSYWHY9or2VZAZ6Q2nOXuNc9/NO0MQ16ZsFTdVtqK2MYwKzIY8cXUFnBuit9YY
RlPtG3eH7CovsN06I7gEK+kpTBoyApXVmiXcRlllKEU19dDk7OO8ms706Ms8jd49
8puZKeiXiiKORGYNDY6lFSoQVIT/dcW0TF6m7NDjaXBTn0o3ZDYBRYLVM0pRmyDS
sORFYK/nFQf+LI/pawRiw96dYZIGucc5lcVTEwLYWLvE9jDrI8A+AjtWZu7ZDX9N
fpe+HHDIzqouzYoHHKLvSw==
`pragma protect end_protected
