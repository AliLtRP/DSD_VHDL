// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:28 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
iIAzprTCjSC1skt4EiDi4HJY0n1ePY2HrIVKFC4CXTVz5EHh0HyZa9cBTQBqeLLh
fnhlTju5EZqWBzLFhTnDzbsEgSpYd+KMPwZc8mBSDFzP9kz4x/V0TaVCSEWohMHw
OxVnTyUqWJZ+lylqEVlwzygfPQO/mllIugPG8HzH2Z8=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5712)
MtWtHbqTd2G/U3m1CubbA6darY81PIg+Mjw0KDeR8qZNjcqJ1GtYgCTNonShdgwD
5QhqUw1G/qbE8C75LTjgOP3Oz3gCcMM+xl0ECqgJ2KsLU1fxY6NWTXKPmLawJ9/K
uan6B9RTSkGMcsjIWl0fLokwvsIs1Da31nLgOHcwJ7A4YVSZJro58KrzmfprVWmy
siHHWrItcgJa+UxMkUWURQpyCAzSQ390Y/VTa8xg5sFxdOD62fC21whaoVjuUlGT
e3NNe1mRkDwytRFAsHXpIw6k8EAHoAx/7oUyAG768e6LbJf4f+5+VG2GpJ9t4Kvf
StteMQ0SuhQ3sQqqfjEY0TDr/PoSsYxCVf4mG57yMK8eG4+MvDvAS/4N4Y4MHfTD
kvylWGWpowZwlK4K2Sdnw8ELO1WjY3j36OGt6WUhspUf5g3hyDAexJq0nwmaLcCc
ZPesStQZnfWo3eXmBKXYySPL4hAchJ5oqRwFOixN5uwnHfmCssIRcTk7qY0p6sbV
uZqa1gn+FLRnzgtSeBIEgLEY/8vvcBGg2nzNF+Rt6r9dUa/nAVlDCmP49VqkXlgF
FoeX3xL4RhHRXp7ryGGvonVAR9ar3hQLX9PUCHdqnNlyBBypU219aWUCeWnAJrHW
ZEp8xCC/MBeTtZIt9MJ0x5ixO7/fSrZwHBShFyEoNIloGDxDNIj2QSHJZSlI3KbY
ivOEDBfKtHQd6If9WbszYpsvFYQ4PwJqpUFKCD/D7SYdnyjw6GOHuWRG2025ktnA
MP79fooCQkIwQ6MkWjdXqfT1zlM02Cf3r4+TTO8oku/bEJmV9gNlCRovMAC0Dcw2
EBB/9e9YFAvg+0DUTs1L9pmE9KavOx4W7nxaLalh1MQLHN4XrmiWTfy1IuxNEbcK
ML0r51QrHpD4GlSPdn7LQUTZ+ns4K04evJBw5XiBwdYI9CYtXeayxhoYAm/Sd7bt
tmEFaAiesYyj9+1N+ojr31kbwMc3q2RmWDVV0xfrWOdVYnxhlnGYE+GK2I9FtdDM
uLOhlYVLgwFMfol6f2Ih1vpop55VL4RCLnXe0NbTDOAaVVbFqIW8uLfxq7qo8ekj
PAIZf/vkTMRSkzSScy5C5oIeJ4K1pZmEutsRB/RFsww3cRykXbuME9jVpWSgO7VJ
SJl0outzEu3YBwde3gmUHAHlm7t9r3OpekBJhJlRwX9ObV5f6aIlWXLL+/b8R85Q
ZQ1OWiYgyiJB98Eg5ptP/cT1pRiBtjN9scOHxxqveKAaDf/LjHKy5yKeaXZSpWeO
gcQEUJYdzNtpmQELamtYFn9qTloiK4lSUXXZdtcmKy4IopxMdUc6LBHHhAK/erNF
u5Of1OrAzQg940gu21RJ5jX+mR9lbHW/h4zb8HjjZcRTeSJCCUmJe6/Eervw7I2d
L3VvuL/wsbYW0TI7x70RGALshP1DGzI29FvCJSTr/IDaruVgwFwo2ezCBhKvDc+P
/gRXPrv91bMM58f3rHdhXlT/TUQafgxfyBqbCfIgPmsn8/hVBS+drip0ex8q7CTq
yXHdrXzZWjjkrR4SXMgCw9zrp8A+/KB/jJmsrNijzmZn8tlwSdjmHtNPzJh5FNAj
wUbS0+AP0AKgvQGpxSB0LdHxJiHRQRylxlfmKWl946+55voChUlRGfP4fWPP/Cw4
ss1Ww027D4HX3iFfF95I62dC/RMk8mq+bOkktQcA6yNQpRqgHEnl1ItJXVzGFeJ2
2hg6qqlffOLIStStKGiVdweJRDu3KfOXiahKdNj2GPehdWKVpBKZjJsnEjEfWyxz
ZMWWwcTkgQpMZYwJV/p3LmmdVStSJLSNCdk7He5cJXAbwimcZ3iHR4DmWKfZESLY
Yw1P3dSF2AarD/+orScaaxta6R4qn0M2CAdIkYCRd8zxPQkW1MNXW+v9A1PQG/S+
UzWVzCWNF/nUGOaekzx44pwu70c0QCOgxn/vQw8hLqCZXlTDp4h+OQZmNpCbcHcg
FQfjwmvQ0A5q1KLh8dqkjeYiV5joh8I3B1sdm8Szfl022lQSq2qvT3vdehQg4ZBs
tydzOmKz7ZePppYZOzXEWB6WdIa7U/t/NytLof0b76NuvhigD2PXdaR5Wxyw/2+I
mmZ3ckJTIZjy6ri+9kBLMwoZljOo8BslP+2wh75c804ah5Hbleil8LqYf1vBWaDZ
vwVIUn/enPFdJ9vbxUxtoVRT9Fibe1XimDooYr9eddsCRStKJYkd8pok7h7j5wy7
mZ13T0DmoA+/7KKBDEk8tqfT3sb4bHR5nozKj1keVyeamIpxXEAkESsdvcBD9J5h
d1+T1EdMsxfC6kXslw5PFWjejQgvyTuXS/qY8Wkrm+1oqg8Wa/OQxl66xA87jeeL
E7Wg17QVl5LpRu9lzbxgdWgV8BxSk65ZAIqpZhiLxKMTp0Z7yVhstCXqj4lP5srU
s7JBo7GQWgOOV0ubg4tGDO1uP9oVuMN035peI/2iM+6nrprLrRWpDSEc0s2HOw0C
jMzNQ3KATDGMEZSZubFj3C9mC5lLKpPhEhBlQ80cTiNwRss/frDRp8SQIF5mVZdt
MlnW2HpZXTN7RW397nlSPCoDCoXL97VLKGjRgbdqxKWT6WbrVMMSHlAlTBEe2k6o
vtmil2SANXxagbXJZNl1SfvPonTPqH6iMcQqL3Wg23GBxTxyv/qoXOM5Y1ckkW9J
xDjDBMxFsA+wGNyJtjJnaUDdK+4imwq0iUXx+Dc9jVNf0AvLD/Kq6q8Bpr5b8JUZ
LkXoLI1dfO8+PR5hUiEUqhwIjgRbSFQynIPMDHIEwzHYgIE6dpzBctHiil0tIZkE
dBRjGtvUkIVwbxfp4WoAjpjpYcFvnva45fBjKO15MlKnEa3ac0R5XurqTT+GRl79
F/6ESISHKiMcn0qUUQdR7ApnZ7tlWoW7mTpq5JrxYcog0u+iMxgCWLG1W+481LFc
0goEH5jSHJRp7e1R/EBq3NDLy5fkuakz9Lxaw6SGpvw1OpEcF1B9d+BEFWNKkcDa
4R60hcoQzxW1lo8aq0EpDCGMKb35GWLs/cZF9NZ2tmjRQm1apvrk3UTVB594RINW
dDHpBsmC2MYdDtKTUM535qBT+TIU/SQPYoo//HnNGA6hNgOxjzFQGOrjl8A/9w60
Sxp9vH/1MxETHAty01003MEQx1A65AaKxu6bjiJbLlCQYHPz72YIEobNtaV67ZDJ
toCSbhZy6gJiwEmwebiaS/ptG3nfnUMXdzhXnAAA3mNcnZKT9RgVcrEQjm+5BtZ3
+QSXhLbILI2V5HLlr9ZKJpaj90KGrkFImHPSuVcpadLoQ2Djmq0goVfgQLp/pNdv
+6RjhdTYnC8jrHwdP4jsVJJGMMfR5JBUUT7MzMhM+2FeaIQfVly8GBx6in4YLnHl
L6Nocp4fILLn+emJ5JZyNgFqz0FAqQtS3PxWkOFvHPqE/Ps5xH4KkcRip9yK0FUh
hsxQVPB4NfbqiFzJ1uchaHHgRWv8pMkmbSMx0o7jll48gdmkjwXvxVDB+dHRP6b/
GgtTSRI9jC/NBMjBiYXciNeBpmtAN3UNiOsZVQGeMaAXFlnD+i/IMXq1Wk31+0c7
rNo0UGjVyAXHy6xNXFILNKOMyCu0KIjMdS4Ua/R571isPtHpwf9A8FKkf24Fckly
vaP8FiRbPdDkVZlCOvVrQZWrjiPYpc9yRMa9zjwUmFAUhald04qPj8UUWfeqUI2t
Hevp5WLjT9uoCnOIdMleQ4et8yCLHHxcbTQwzp8tE+iUa0R91GFGqI9ZfL1pJXGU
j8Rjss/A/7lWP/fQkwEkuFXCZbz9i8oLK95ujgPwFinALStBkp5r41oyiuo2sucw
88YoQtvEWgSWskNWCdeDN73C2FwIKUdBTBpnCXxYwOrpNwiIf8zCzmUY6LepBPjR
8qLDygNNHJBgRrUCaCw4sQnQLydDNgzNB4y1QD2pGTP+jb5SKF8dhXFHAEfikJyJ
W6TQ5OfjxYIW7d7nxCjSWEj76OWS1eWhTlbYky0kZD4q4DYiNyG2ZFAfwTLu0n6h
hmuFlwNCAJG3u/y9eY7pkbEMe9Pgk9DrI0SPDLo8cC/h898fwBdShk1eesLrzWb0
TFDQjwnNX8sA3Ut+SecJso1nX6Ehojk97ydB5H0uJt+dD2IlYH70ZPfkbIaBKavs
iqxtCqML0BmYbQDWs9XuERs5/NhQzM51vZB+ADduA9Rukfux5y0SoWaTkXDRBnuz
IHI5YZP17BygMoO/1x3rd2g8g/5jyuX7bO5CZvpuujEcDyfimV3Ggas1BFfGrCyZ
3nbkaLy2CMbefuFIZt6n2zF0RZWeIyFZAwDeKR3+mXQ8uiE1IW6wXbFUZi4bouFg
velAuWgffZ2Ls+16NGLQYzhRBj+wgDqen8GTMpOJOEoT6phYatKLVzDOxmxZcCzZ
vSW5xi59WMgEVzutwd+Ya2bhG2EmnQUi1qNocD0SG4dHL9yUfW+8NsTZsOnxpVlC
xKNXu0WowtEniLX+H33nvRUF38I6GtZL1fum0xwY+Uaxr8CwPHRSyidLoiqgaAuT
XeNyyLUjPoYyVDV01PMq3P6ah8BsIQcYdCjw6feZXEgz9Ccih99x7h+mMRdF/GG+
/aF0zOxApPwbYYYmCaACSDJyntQ8lkPD8W7W9/DWA5nbofNp0ZlBVt8Mtg0XXoqz
WYBCRcq87W/+1R/w+FAkPjE6PfPV9h/8Q3d7XbvHVrH6bksV3b8SZjjWy/jVM1lm
EfQuchFp2K5zjA3FoHQVW43CPEY4dFwmTmg3mrJ484VmCtICH47xYQG4RmzfLufN
+9FY5ExuNv/AZ7d5/nMOI7V9dXwY6gDSMTDcZzC2YqWl26fPWjfWPgJpywTzd4Mp
lYj9Y/Dsd5e6Sh20oFNCG/ozARXkhagOyxK3MyrYOvNdjMCkhNaI5zdvz3ezrcsY
yMrajIaFlpd55I/vzoYCRk9qfSf5yDZ3QhsZJ1bc6x9yN2dwmAvttw2ftzv5JpDx
LAcCBThqJ4lO41KiO8tcx5jv6sUkyYE2hnkKknO+D+SpeAGkQxP9cJ/LaP5DPsqW
AztUlpU/Dbim+8UBFuZX7IuZGcnIWMeSl042oz13PELHxFq9MDwkLeyBgAk7UvwN
PHeLQsbpE0uXY6YlM1s1CWcTAAjnp8aGOAT6Sp5cUuRTT8ytbgAq6Cx8Y31lZyp8
8sx5/I+D9egkzbRn5rzH7MCYmbIfIIYAhR7+sTMN94Jc+tGGTNYxnbGQ7AJwIO4z
MxFU6GCH73XH+ywVva8w0WyZH9QkoVv9LhER+FZjclz9I4cNsoCgoayQkSKTSA6V
DEL2cEZorCq/sOvTel/7Up9oOtT0Mh60MEtI0udyjgEjbBHM6XntMhhCa27p8Nv7
M0EU9Xb2WmqBj6BZ2tS99PRVrL2LsJ9alZJQH7XGcwSotYAbehzNHaR5Nm7xPaXl
rLWXv2q8QwOiyvOzHxZYj+Jksopc5JSoMmGJa6j6tpiHpjO2wIDLUveeyDKtyo1u
88mR6N840zBft1HGvidN35aDbBx4/0n6wg77sstL2bCipAQITsnT6aPSOHcSWxSG
MOLsDfX2z2IOz1r2twlu6mC2sEZATCG7NriFVwQgMGUGwxRtxkhrB0FmL30DOY7F
pN+CkTUQnNJCabV9r5b6LdDO4ymL/05GvRqdzJf0W+pm+pmhYwwTbtFDi33bl9mP
yunl2v27K2D6ac+Imvs3cZXtJQTe1Zg0b23DFhUa6wT0sGFbN6pg1ofDmQj74B4J
5pwCpzOlQGO4tTDRDc2iUtA6wD2g+Hdc/m8vgmY+a9djW2+8d3Fa4okbN/ADQJCl
KuqaCLHw0GvGho3lcHJngB8AeQ7A59yViOOikqzSOV3Q1/sasHOReTKONw/aKlzA
pm/8ObNnedpMRyYJL48Hd2eJciuRbREDjS9NxSIJwkGNATQZwq960oPayg53hH6Y
BiZ/jlPNivVgJZfulcIaqbobJY/HwUNz11eXH6gFFrd+UYn9bQvVx0z7omrMKFxt
BDEDZBbyrGzOuDSSq3r7/oXPYPfjhqqKPSG5ec/wfPG/7Y2IULKXKgkvNQ1sx+es
7jZZuQDdgxye91ATdKdyfeu02bsEdph6xVESsUEateMSWovLCUKEFOu6Ngwxzvx5
f7qXD9I+84nNNUCwu9izAmUqu2AU7WpmiN5ht1LztVglVfR5/Nv0vfj1NyPiFYGs
FIXAdsh5HYLN/c+2vrcwdbjrE/zuSsIcC5mAEvT1ZKJ0bsO9KeSAd/JjDdeGY0Ly
V4AugZnksANojbmO8EJs2PqNoQigNnfy1aJX7DVJ81UeYGRBMnTQpn8CHnEr11/O
Hn+03o904EOkggm2scSEAkClktZanb4kwssueh38L9zhbsqPLec+SChNDIq3wetx
jK4i6IsXOt6tm+oT1PiKkoZjxOuXkItsJhcgWkl6Tt2tWQEvaTbrWWU5JU7jcRB9
Xw2FIL8UnuhkfDynROLn2toPiYGR+SJkEMeaC3RnWdl8dY/sWswvyH01nXiNMDCh
KqOaeE7HBdMnN+wrFwurHY+Z4NUmZHXBt90wFp5Kwqz9/2OP5UqC/ge1BFnq5hEU
iUP8glh94TLquQAEefHtr+ar1v3/GHGCtsy1KI8XdPaCLhFyCiZM5DYBlDzlR000
p0AKVIfYtwgzLERYQDRE9cIuqSvW5CQ2kFI13ihBytRLI9rEqBjPnN1yg7BWfyyc
6YoZ8D4c5wlzo4ad0y19DJUIT800+so7i/oN5vFNB4arNjaJkt5jtXrnJaMiwFuA
F69MvPq2EZtsuiSV+4j44tIXd7PuhMQRpe8PKJnWfctvT+7mKK+kopFg7WwziWRX
xegiGYIHTydIkwm2UanVSrx1O58E2sUVgF8l0RhfveL2iaHN8O0kTwFFtMpL5jNJ
ijyPRuy7O6BpzV7nBTmZ9x3uUtKQNqwVx7htLTH8qo5s7wofERLJ/xRv6lxB3MDz
3Su4ul8tDb4c1oI/mT62dnXYA9vvyjP9jyIMKu7uBMHGDAoRP8eoAiY007DDUMxV
ppusQZIII5zzo8WCpWR0KQLm5+zqIhCDJcZzA8iSWEZ8rjPSGzcg8nAKXlSlnsYf
BPhn8tvmu0HdmIxblZ7ytWnPPLgspjl4QocuKfW+Kl4jnz594j5eCDkE7DDgf+ym
JK5ktXdQSLJNg/KjII9SxUiiiCF2Vod6CQhSre3kRQ2WeprRo1+m28vbH4O267z9
U0YiwaUYvq/vSGZJjk3LfrpogL5AdAQOjHYmQi8Noverv/L8P7Qq6O0hNw6ZGTC6
Y7TC98ZO9fpH7FYHhWXrCzxEEfX6edcXaxOXM3D0nobFIgTppkCoM7EK3wASqxcw
j4WjBBuGeXNaZ7+Vl4sli4WQlNHNWmMSMpVhKfiUMVRC62Ayk71h6ag5AXt5gzkR
itp38oTsC3wjhQi+2gI8aFhg4U0ZUbJ4QMEWwFeluqzkP3iZPZadZByUwxcYqXQ/
xvnwOgA5gp4qJ1hBywW4cVvYIcw4iMMdbjxY4R34Bc8aibT7JD4ZLhHgRF+8yZYi
T86Bp6iBULjQsH/ol61hmyhwuUs3LGOm8kY1V8i66uyKAr6Lqc806HF4EnuWsonl
`pragma protect end_protected
