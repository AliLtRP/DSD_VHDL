// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:56 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
eWsBNw7NAu1+PGo9MGifq3fK7ilChaV4uOl1fzQYvITxj5jDXewmTpFtCSkj4+Q1
uSBaGB0h8tSs35IYoyfD4xbaXc1Wtch3MmlyDQ312CHuUXYDDQ8A+l0xb4iQXFrZ
awH/NjuiOwoS9d1J7Bvx1+Rtkz6/435u2LO2QCle1ts=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 12976)
FmZ8vNr1bRSwnPxOmYDLUoFdp1sTmCro55Xf6NP/K7q1+Yo6koudIQJaMjugtFiT
AVTUJs+RNp1cgsZuTdoTGMM6Z7K9SgvWvtTZemn3QDhW+45gpZhALoXc9Va9PCtJ
qnwUql7+nCEPjLNp8LBOH/VOKsRGCnNX+JX0wT5Iy/wEpU03rJ9yQ4TOH6UmJus3
Y0KIhRDxmpciuEPATTASr8xiigFlrDVsQRS8TNeRAFT7YJzgs13r9cTa91votACb
Rhxy/BTVbd3sUttPSB6HzXPTVntnNh1Yo2rurfhLH/vzGICoOAGDlse7r0a0uV4/
qq14yMmsuVaJI5P0x+5iAAbSqFiyTopgeXqD6TKifeehby5X4InW7IhzUVUPWgmJ
W92zbnRJYuz4J2r2HNFV5E85duf9AyugDfOIQC69crxOCNr+wk/ehcCE/LCwM+Aa
s8MTaXWmoFwDVz5ZsrmwTnkWfCIhjPouyL5jXF/Q7MwrwU+0ebVW8gtXpixQGEwD
xN9TY0xwZdOptyO7mkbIBowm8AoaQ3bO47ic9Z07B86LAqEryixRu1WAjiWm4Bhn
pU7MxwvuwRYPCUuQ7U/h6rSUE0ctnPQEaWKaXk6wyQ4LDAiAM9KPcDHGYF5Sgg6k
7R0wbvNjT7UYTtpqfN3Oesbtjt5pTVTW26pPtDDACpbCXoOOeQwwQpgNMw7PWXCt
d/8IMPMGpvfMxQtojyZc7wXuuNGxqa/iyMThWdntzC0PEbCKh/8tnpK1Fckyokvz
+fJrfK6KG6VaNniOMxuShCRo3QvH7S0U2S6OfussEW42aeuz+hOrD4Td+Q2hdlV/
V21mBCuWlkkG145uQHtjRRzByYQvuLVhM1EtWHQoqAgBr/4EaOhkoBwjq83mFno+
4Rf91Fc7lRSi7V+xr3MK0BX5Ldo6L8CJXCMf9MCDLbkIOvuPLXmX2xeVGANp5SIB
WhDb7WFz5VoJ53rfBMda3OVspqU0jxKaqdv6LqfR2PoH7wCJkMcROITdesJZODU6
VUE/5BuC7IeDjGEJKrRK+zG42ENMDFBxouV+i48MXrxxBh1pYcHgJomaNk6U+rFI
Y9e8/y0HijI2vzZW4JdvXPBCaPYPUF68M0mZoHOfp407iTPl/GI+2GBHCl4XIGgj
nhImNyLUdPF7znAqoPqbE78JLxBHc6em6lznLf7BrpOoACnjgKxkNfTnNPjbaNkj
70uES1EgbkcaiqJyRlYJqI8vfLjrJ7uyrcu+LvbK3yASwmMK+EIvd6dNcU4W5as6
X6fD3UI5+W7MPnp2K4v+htG+DF9UWdhDf31x2J/tuIKlCjC0zJlc3FY+BndB0Ylr
wG0T7TLJFWdrH/4bbrbxUddMFO+NDs+UzWCuBq6jLPVI59XNB2dVacaZqGxiRBEq
Y2jDcHMhI7Q9BZQgfe3c6jAr1EQBgDr+mC1KpgXJIe3q6pBN1cyuamoxbvjJ175F
qe5yIo25c0qR801w6wUG3VC6+QGHuRlhV8YavCsGNG40PoK+MRcH4z2ZvRODOagy
6KojIpoK1SJNcEIRr8PI9gm2Nq8kwii8ZZ1fHEIgxUdpnli9IO+yNcQAP7jhXnfa
W6OZ0JgLK4bbMilxMEaYNYhyWbNV8iyTTYKF/Vh3A6t6JHpkX1JydRRo9wYP+Yci
4shpnmXvgj8ZY4DyvIw3mXpr628AWnhE8IVtxkV5aRN04L4KGuzldrYhVZXxxpuv
Br33MokgG618H9njaLBzaP3jfmteA/ZGduxBYUChEBcXzlRfTOJvKi4tzv2HKTfa
RR3zaS28GLqSN/r3IH6wdruffSs5iZhbqvY5JEaCNZiob5fkGgSup9xTnhwe/vuS
mtcpJgrU4tgcDOoga+pdH+3M5HgU4lPto08f+7x5ebFUbFtxUXaPfWyGhf8dw0h6
1g7DT0bHvhM/OqHz1xfBdpFddacPUKqlhvAxT6p9YII7l1h6QLBN6e/dN1bS1Hj6
/A/5OVSXTuqT8PiQchPHNNYUJmoeSBKkekTbaa3dYYbLCVFBFr3d1Nrz3FA9okEq
zdFNVFa7/onf6z3DqJNzJtaPun2P4CK67nSf+8OEG2WMr4m/hwOKscvBhn67/pU6
72/ucsQUojW3NFhBuOZtVK1BefJ1CBxiYTk9Eahj+cd41J+UzxxCd0vHn88BaQ8W
AvIObGSTPwzwCevPK68t8oQLWqNQQp2MMbliKQFwhPmOwI9hYrd0iM8m/zwVozkn
DAcMp2P6SIvFv2gIF+9Ukhicq/qAnh5TSgbH3jLtInYPFyUxV8pWfHtlyTiOW/BO
SNnbZ2hG5JSEQ7P01l9YKOWP2nSxQSWdr6gukQ1AYg4tN4eoR4iqOKoZxLYRg3vn
3yKTrBds2ReDZUlVAit88ZonXC9QVWcCLOU9FuW2BYS8Q+6VFY8aNrq2Eh+Sksgb
zJ50ZPN2wqzrgudoBaIS3Qx2uyj6sRcMOO4I9xn6khQw4N6TCzEXIdhKAY5adNK0
uu4aafTP9MtiKDd3xfr6fBappJI357agyuwyaJU4ZB3zO96GFjmaH4pdQB88BrjM
SUFfOhckTAvMl+yPuy6K8kvBJ1AkHF7SiuIYDdhrYluOwCo0KPt5BZiDl94eUoBc
pEV+bkYrbGXJRhUJshCQujVfCHde52X9zEtUEi/eDEVlUY6dsaira1QnhVwWyUof
EXch9/Nq2p21/Z9kwafDAfajUopQyp3x7v2WRk7wOJvbyyAylAuAddyufPWH/rnv
9QZTgg5nJIkuEXcHivLJKJVyWDcbLdVwSHQu70z1/S0wh5kXW1/j2akjy1+dnAQZ
/0PCvkAKG6ByW5ERpdKftvmLOWA1fjMcaYoiB78e36Xb8GrlmvM5lDPnmvPvp5YO
IRb74vZaQet5FYEpNrDyeL3VrLMbILSZNL1Pv7YbWS8DjRnVZiUtrVM1mbgBQmLK
T936QE2hXCF6iZvCrjreXHI5nbGR2r9qsu8rIYv8EVRN8BipeAT/QMrRrsXCbXhR
67NwFK8zKV2UuJFdf44QfsPM8xf06Sn4d3XIcRxUy+6Tx+But5jArxW30lvNrpHD
TM3dA0GjMNzlyYZWt0wkhHTLcJiOkPMp/gxYmu2qzG/+ohUhWqrEv09IBMIiNr72
gH8VYJgzBsjm4EGbJR13qe/MaNDE6+JMynOvSdsGzXeAWlZPr0TWAEm6aGHbqn19
4p4iMIf52m0kg6KH2ewrtAIjIR8mGAHdzP3NkUfXOC+piWOiFTK3g7Ylp3K60Eho
A5H0QVP/XAc01DkXxjrjZ1ioxQDTGgV+k7WukFcMr+qFeIhJWcx/dILiE6K48/ez
na7XesYWAlGgWLTyeBTYGnMWLdCoiTDnoVHj/ZH4IGDYMwstafBjgEi9bPrFkpa4
tLdOVUOkYs3ESVvkIUIC0g1gxG0KZt05CMBnTCFekgWDT/n9U0QOswtDUGuPkgSt
p1r3GDILmu7hRigWUIl6XW/YJYDIhCbvvNA4mxbuSjGIbJap/u2howPpl8bOWk9Z
eFBSF0jIT04l9ko+FLh4YZ73bLYAexZZMg8cHByDRXE8MtCMUInBQtA15UiGwmOH
bN4igNcrjOesw3XuUQrsY6P0BU/QHkSYYyOevFRbiq5AOy3HE5kgwBlhiL0zAcV7
M1LPg1u56ayRarP3tlq8Hd+QD+pdiL2GvBu2AHhzfTMEKpvntMoiTM3lgWNSWmOI
mD2IViNgFrsiHlXngHQHNJwuaNmGRY04V949vWmAfa/ritVXY3hRHPYrLUZxU79b
Y8z7LVtv/6K7gLYYynMUNjr7ekTbySsgDTHcSvGHo52KoqTwX0KR0Y1InF/uES45
tfcUbDTwS8Gm1LMDfWcwm4HiUnbMasDc0LQuA63MLGD/xYxW94EakZoOcV8DhkBb
mmX0P/ZRWPKl3Rxat7DwYCHtzd7ScnTkYwQNhhgiBrbjE+cOXIsEOpsVQHuP1glP
5O84O5BVrd/dvbDizFVajIVjv9ie5yCYhvP1kZzM9fTktGGfpgkKHrDafxDAoGZ0
/6BVWJ3x6bjtWlS7CcgKHlhyqTG7/nCr8N4exHmi+7QVJ0jcBsTtiAXoXZP4e53u
5+UblGJvUhtW9WHF9RO9LoqyejcSETcw0USpo1lhcJCj9I/oKewwvQ0PF5HybkxD
0EtGv9+cj9JAnRkapfhr8yH/Oy6Ps5QT0DkTEue3iIWjQBc2j10L6Z0y0KDO38oe
fS28yE0JvQ+Mia6q/tBFD5rcjJBp04lo30uJuZqPqO90am8sTclX+8p2UY3P06Wu
m+9kZApcbbR+zVP/ChctXxKK/AVQFaPoIU6QVyG5A7+bOjT3iKnXmZSsvEMOG53D
5abthNhGWVaTmqbaKnT3dCL8eiSvqUZZcyluaV/Y5cPZrFbZoufykdBjw/rFul+d
yt53cAxSvNksgSXl6ks8uJLnTa27UonH4l+Qhxx3hFgB7HBSa18TyaP8/669Gee1
1hEF/VV7OLFF9CAAdje8BpXHzwCtk7vF1Hcapq5J+ttrt4tVDHIBIj81ypj9QThg
AwsoKvfERhpItIkPml1o7HmhM5T9yYbjFp77dZsWBfPcREtVK08SEfHP2/GXdNlK
eFhep14YtcURKNuEer6gQZu6CKkZF4dbDoNTBQ7d9Rn5pIGdKofm/Z5AtrBmQsHu
OwTfZ1hm2sckwFeoeREUioJucziKyDhHeZrO0tdrekZWdpEy2ydQotXeQeqsf6w1
7p4LeVlDFnGVFp52uZl2CDHKH4+i+wp6DGTXte/A4XwHbQ5QXeVLNiizT0OXttGn
oV+y0UP3cywWlJfwHMi8rrZtnLuqzTRg9VmcxBNAo4VBgpwmyTlH7U57qAZUQh5d
jWUaCy+dBt+fn9ssaQGznDYrstioVF4TwVJemTiNRfOFGhp/8zGCYTufrRGAiu0B
fLbggKzu4FxOgWcE64j9S981PkpjLon104u4bEYaHS2vjSrWfJFMJWNWaa5nb69i
0O1npr5aqPu44Jku65noXr30+WG8lOYxVkVkJMqEbMTuaaGATX6ME6eOR2Z6Lx15
pZ+dq3/A0lemC/dJDFPWfrnTEkMYIwpOMCei5BPaGnI9jljZWDf/qAUQ2vB5btPc
0pbSGZpOSC/1HcFbqMRy9JU6dU1efMa7pvDGIgJ5w6kGDwIX8AtbM2lgewJwzd1r
uBodFkleA4H0lb9Fb4MBv2bi31pJWNMO9taRyjtIovzIR1lTcDNgrb0qtcpZquYO
cOHehucPfXY/2tzC678pYstZ6GYIpRdUCKuqkW2IgfmFr1W9MYMu13poJ/5gY2GN
cFiwyeoNe51EueRitlmE3x6JdiACRVWG/f1kdTsn9x6u7tgbVQJIyVDrRSj8imBp
vEwJS+6MagZJEUBk8om1zYlHdXeXQn87csFFGj3ElmbY5u3bv3s+m7KejM63ypdm
bQw5+eLE+uA0hiq0bkOCPbr0JwtpWeyhONWib4pU5csqSKZnwtQTGCg2hTCqf0Nt
nYHo7WfjHxjWPIa3Ph4vw4dJZUQ16TY9m+JDqSz4zaiCJVF7pCvCtQdALK/IE7T8
BZQf8Zb1bRs8hAaUH+NS0ao6jkHtOJybuh3Y8T3hCqYGDEcV83yjXGv+koIvk6ef
8CLdssc/WuKL6gHTkmVMIXiVEcvcSynK655k9opPSoWmNEUia0/twf+CkttMz61X
XG/5WWVSdkdrmlTMpWLuARhRNCrd/4q4bgLWRWiIXM9uhwOh2Vb/V52PNIgMwdr+
j3kgH54YHy/h2Th+cZrAArBeVTDP9sr9n7l/USAJFNhQ4ke8RUxShB+XZa5wISiM
FiDMou2AILVwatd4IdhKr/kA9FXrh/oQa7lum8fgJl/DNSUugOo/iNKqUYL+S2Zn
ocQ8xDWq8NhME+ZTb/XxpYxHSrysqQFrYINzhuXTLUZLo/GOLhIvefpSvO4+3e5c
f5Ji2Au+TAF5nU9y40rHkrCF++v1+utoU59Qyzn+KRQ+K4qsyGZ7ZuTDXPxCGgeR
+3PQ+JcU/6OhXZW8m8wPmJI/x+ycPuTg6iMerrLrRHsTNO11fwxA+n6gnbRqZ4Ut
W0b/FsS2oF0kLcrbCJhkehgdCJ9VxhA/QxzJ4gGZtJZhxaTm0HsRVr/3AvgHg8W8
T+m16hAWFUpikiOvwZ8FVY+pyotlbxQ5QCN94D/oZRgUIh7uUkqwwJw3au2VPPbI
KnnxjqJNFM+IabWj5zBu0RtZJSXCDuQa1ytFAOwTa20q6XQdHfkUm6GqpOvjX8ge
cs7a0uAeikFK5hWDLMETJ1aj1PfSWnReW+6bSP+cesDwJYlSbIwmZ/Gp0dOXR3tF
6qI4NBy4hCq5JZhTSHPxcUYWk0R1SJJc6EDQ1RB2fA5c5x2rLVmpEYNRpWh1vIju
rkdC3ll6UrgGsk2FZfTWxtixoffKgOSl9Kyz0In3v0fhXtGynSgEwDmKbsJfNk0x
IO9DcvgGLoepMYLTxkC49vdmcJDhaEBoCMqOUSGHlKEjN+6CwQRk5SSkvIec/A1L
KUX38DlzFcr4ovu8CWnJblOBhRg4B5neNAQNC567tGZJVA/75M52JQSdz04V4fmR
03g8vEr9GMobfVR4NAsq5ixPgihgSKlfGL8g8ulQnltB1TiXq4ioz04qVN4ZTlOZ
zPaUPcj2ydUJQ0NsAen/D6ndgr0JvgZFnAS3pO+VHWEkvgRfxZIIZ+E4jCyXU7TS
8ww1ep9vas5P/pLbN0WBdAw+bAfDeIBOKDYR2/KyGdAaNiR5iDWMz1idnCr35TIM
/oiMY63R9oyGj+4hl0dn5V76FBxE5WtFkXCZfdyZK9AMGQ7wS7BfU/fDUNs+iIA5
pVVZ5gkJRN3DI6Le8XwWNAC6z53kcjyP1iSY9XKsk1/FACV1yPCmT+wQDhpEXA2S
QOgk7r2KxMXLDGvR4ZpkocLDaFbHW6BTfmgl4SpTSm2g584evM1z7qHXgJka8v1l
ryVSAZ/6+13bc+q4zj3JhBKf9X5ZnOvyBSvFBItY+slDIBGsfwWuvhz3uczkW8A4
ve0qX8cKhdEzncuSD6NXBqXn7rSasS8jZIB4/JxpGgGZmL32SJrhrYLL2bUVgnCT
CfGMFK5+nHAXOYwVfgolAqqGUNxL0YApScMSMC/WeTbNdGjLKahsE6K7cCAFyz4O
q2E47OjP5hNvVaFWECxThxOp1Ifabc281lrxbcKhuBRYXnX594lUs/zpzCeapxI4
lQkmwafQKH691E/CifCPAMbrZ7hJi0sZLClWrcS0KIbI2jtWDXGAAYcx8U5PtiMO
lt67XaqcFI8HxjnhbLt4k4jDRttbd875REwQ+cqNj0l+z2IBOPQUtdH5NE9NjD2C
Ean9+vBNB4MFAlO2maOuqJ0dHCjfO4mAOXIXwoA2POqpRp7AQLRNHRKDhhOKQ1oF
0bdjMbEWawdQKLau80Mj7BZ+V2VgRvzd3w5KKYNvOP1hqWWZxp6WBX7Eg3qMJSjj
KsHuDLxtU6JlMJqgBcMZVKaAkLJEmdBR7kucNFdC7D84+0/sUlJ1octhx7JBStsy
N961rAbIBoh1OFBXnJ2if121xVYf7VkiYKWnAI+O+hIHyX2Cr1ox1GS6LPej/MBN
DiqE6NbvmP3LrE0Tk/xoumj5jAhKaZnuQfP4FULax2ZbnO8EZVDBc/hR582vtgsz
kxW7KsJHOKZqSAdA+HH31LScR/hNNKDawgOpwqBuPd3YD6xHSVWF1gDWOP/EJk8h
4b95K+xJzgs+14hhoBUaRRZdqZoWK0RV0IsSnKMwd6kzQEK+DrhS1asBCEvh5cpf
+H/iFwmt3ttjExUNyZRAn7Qvuo2OtdzV5r3BoCG1HENAuZ0zvHtVJKQaRrptko76
RjnjowBC7mHHPSuYraCbMk/irsj9b4iim3oFe3vSCXnRRGWmz5Y0JUzV7ubZ2qhz
nwz7lx4zT1c34RxX54Ml9YwmAL9UifLAiRpYTW8ErS95NIj6jBwV4ZZV7BBi8dl/
q0Qq48QzRj4UIk1QpRAYuriT8OWgDFRN9jNEEck2KzWHRpZU5hEkSYNJ05ArT4S7
tjkBzJ0FZePRVBRnsxqUrgxcKBcH/mobJuaMXNry4gkLYYtoEYZ0Dsc2rS5z5osK
HaJfmn1AxSXooKMmybMQzimyJ8X/oPslIt+WfryW49H6bfLwassGhBTFq5WPDz4J
Vhc3C5niRHkqtSPbm9Fdn+kcdi+nu7Dr/M0yi3whX/fHnBLH2Y1gZIVAeX3wU6dM
RIe2NHA/KsFYzJ6Y/6bPfhBWRRbW/KQmJOLj3yEigvB3rcRm54jB5uMP/FXXCwfh
jsrgvl5BOYL3fjqihRG+/dmrCdfVqLIKf74Rl4EiUB6k7VUPEoU5ofxSnyjJfIT9
HWg8xqFJp4VlGR0vEF7WpfmDAUlDyYJDIlwG4AyeTt7iK1DF/EbunQWJifHKjWht
wjIzTEmf3Mw6DK4xOBNLhGd567OL45gaYUkgHseweBcseyC6B/COwMtx2gdOPVRP
8y/vvL8BTgnmaqwd63Z4ipl9aw2LQAwe0oJz0LvOnGHmAnAXDf7h8Fz/JjarBZan
Xq0V4J7b2VIy7K56n1nydtlEtRaCokbFStziWu96NVVaY5MfheHS+wSgUp+cyP92
o9nnvt8eKf/2lNtLSNFCsH3Sa64z9TYbDlvv9DDA1/UWVfirBAWCU+9bFxKM7ctL
mvZSCCJNCW0Tzh0ViAabBJ771qVGJMCoaxerW+Mmz/H+bNGPC8kZteEGLzUCUjDx
/dwD4XYnfjG8ff4Kh/MEfNEi6OSRpO9sTHHyobKilIqaoXN3MWifcF0NYQoGvQ68
ZTISWLh9/gAVbLfGwx1ruHWbTo/NtK7yCxnRSVwhU4dK6Wp7yK8NT2oTVOPGqgKB
3WA+Ui3l5FapK6Yo6VsSYlHcMp7faOl1wV3kjawU/siBXBydI3nubwHMVk3nm82y
hDwDsTqgB8X27bJjGsCIXa9V2Tsv10JeSe4dLKF65R4tU2S1uVwEAzUoOC6SU08N
08lMyVSF0+7hcIF9oR9liUlng65dHBh6e8qPcmVJ+2iQbygw5P74cJbnoS6OIkhQ
cGrvAdQsEBB8r/36Yl3g8f4oGbm3sYKuoE6Sl/VvVfI4CCkmIBXGXtczLsBzhBbC
FxV4yIFi9ZxzLBcIYW5w9ZKgsFOtTIQkqQfsL5jriTqdbVLkchECmLPxcWvaWLAW
4RZ1aZm7zjtOYeFuP+r6vzTDqlZ+lKe+0CZvWcmzMA4Xa2qN1hDClomTiIaShszh
YQdz+9UNSbYL79lbDhfGz3sOiCPlDXpos7PanO0tTVxxHjdMWNOolWaEcxblmTSn
k7zAv5kucnFI3RP+LtXKIygX3wcdJNI03rz4gykUPGDFOuQRdEB4WhKPBpE4Lw0X
dQbU3waEqWopOR+IP1FNDgEm/ECxvvBqNXE+1H0zJgHt7OKsymdzzFT1PM6Gpf9L
Y2ozUH7V4r383AgnrToVD4WaRTtrRSre1GHsipVpFRnpQRtd0ge+Czmq2eU52VgM
MR7EFc7ozHAC6jt+xS0RAaeyUuAEBTJQBN7gx8xxcvrUDIXbO0TkAvugqJ/m1aH9
O1zxXSy3+zCn774vKUvGByCgwUkEfPNFtWlsgop6VZ8kR5wN+mq1RhX6eNQoDZqX
rGULBfEQ6s1UQfuWzSiQ26YAKwKEfn1PjVABUFMB/JWusIuRvrDQyJBMwmLVMUID
hGvLWDBPi0sTdU7xqeAFRN1zPUgiLeS8bZGYkESM92o1y8uSrtlj4DZZ08f3TQrm
HN5nMa2ARTq+ikfzMGKSuZx+hdus4ifHSmXy2Y7y/jXIVFg26mbVNmj2pRpD05/6
iWqvzsyXm4/D7Ty2ZXeiKb0COYJPehFiOdkdBnWhCtxtEY5IZ5D5erR3r4xpgXg5
unzkrJVq+uj+uUpKuuqBAxCTnFUcne+YyNmMRucFEpCavv1opyAvj8tEag+Lnpvx
gTJcq3xQzQXFeCL81YhnpQ5YHbyaeEtWbw2xoI5xSfkyxIDv67oa9ZBoZQGJnBOB
+CMSr5XTULq9RFUjUJVSGv/2iduQAzh9DaUPmresikxQTnJS222fW2v4e3Wamscd
8l1xRXFeySBY29XCpLQfV70GJ6oIIkAk8tsbNzyrqT2yUT9808eYy3zcPahVGP0D
ohvTDlyyKbx443v8KRRMB2On381wm1Wi14OrVVSvvVqCUuA3LOnnfPw3atNprIrU
D7KmTwn/Pjy+jF6EZZhUOkWI4j1D/9q4YEXGnTcNC3M0W80dPapE09PKIJT5QPp9
fgtYBuwdx9yALaWuRYhJh/cmsyepL/M4z8vdbZINN9e8xQFvObu7TrqmFeW2oMsI
5s72TmJIvH+pWqL3vexsUIZuk+9JfqbM0Sh8IcTjqHLX8E8nCBS//4Gqznn1T1ln
3KF/1B1klSKorVb9rOEy+YlU7Bgupfj9yQllrJLqW9CY17T4+JNt+p/oAeejTMsk
bmA9DBcqpPxYBXbsfuKozjM8u9KPyTogdccTKZxNkxX03mL7OrSLHPAs5UAxsas1
UGTTNjXaFvoxETIK63ZTOxAIPEnuyt+kufZOBIRUITV6a4/Zkvlj6r0wDH7CnR9x
jImLXBcnm2hDC5xElrNgnjLEgsGcndQaNVQJRmwawVqWbcXBCy3kYFdLhly1NOdE
qzjOZoXGznmNtHcCvlntAOoQJ3/Om7artXgMAZ2mLRJTnXcCC5RkDFpkBk8zhpSi
lkRmmiMAlkl7YkCRnEUeGIRoaqR+F+K4gefFsqZDiIhU8L6xZ/wj6BSBG7YFFf8Y
9cx2tOoGiIA4Xfp5bPRZfOLMbE2p5/wa/GepMjPflJZu800+9+gHdpm4F4zDy/43
jkG5ckQx80lWpfP68ha1pcD4Sh3Jj3GsmOoBpYxXpSi2CfyULg41/jzie6nt/J5z
afKd2kId3A9dghR0jhWTYq2LAWuftiGDMuiBNDRqhTeQjsS95KpyfNS0K1BaMNx1
zSW9sx8YUbgBu29Ke/yHoGwTIsBJRZm2ScesaJb5P9my+MChE9fNHGa8M5iEWjpa
DbAqYXicjv7sVuzTWr0+nrU8zsPOaIUTAFdORGTbIDxNLPkInMjRUVbSSoMD5FwZ
QpWWSWwDjtiv9cGd0Y7BUa/vGb/oCqbja4ujHFK0UE2mV/zrU88A24k01Z0xfy0p
WKbd7MUOQbwHg0xYQZHGZka0+XXL2xViLCmiiNweZ5fwWWXqOarakR3f3tFvQtWr
X3Hu6gh9q7W+pNTNHrbACf0krJFvQmhZujgOpRm5Atfs2xBUUOevxAod2XbUn+gZ
+joiZOE79cdDRhzMcs7bEZC4Rn/ecwY6OHUDp43YptJmdgRbEuyQERzuQXGB2/bv
jynaPAqxbeko5K9cZUHB1cYFJaid+m4sTVKi4D+UQ0XS+dX/2tB9KGQ7U59Ee5SO
07ldlGADx5652/HZi1MeHOu9wdkl0wji116yO/sTxhHQIEy7+mNN8ravgHFTdydC
bjCleSg7L7DdexSZ4uQlRIDhEbJRcPuHtg2/rXbNC6C4aAtii7PmMceTcVp0+nxW
YQyyYdv9wovzOvlbDGandAhZ+w3Yrplrug1Lo723MRuKEbHMySwIyn4AhPqeyx/o
mPTKOhoC/4/edE29sPJ22AL9U2n/TRppaEHRdYoFF7x7POFXMsMUAynxVQ5kL02U
CpLuunTPa6SRgp1nrxXjuBFx3NygS88zZTf7PXlUYL8Nu2BwUQqrQNGaaJVDXIFe
67KTRKXYU5DXy+2r1/8zkP5SK+gh9jk/CLOPVlNlCCLzPladom53TbmRjMnywxIc
92wTGwQTtHXqVEse4jzMBnnmE7ERc3cTnPCVKhNAa9KsJb/ZpOXTbX8EBYzx2vky
XFZSOHUPhJBOmJBPpSusyiS7r9FBv5Sh9Yr55HAArHkB77QAA//e6IQ8j93ZZ1kz
Rlpy8KNjO31KgnyAId7gmsePMGMDkKKfPwyXdXxTgCRvpKRa9cuzXOSa6ZNS6m03
OFu/Y2iP0e/cgdoqrBfeRbIK41+OcBIuO8z5mMXXd2sRepiZYMKu7pXF/SXGOGkg
od796KkduiTGo2FAfxEe0OOGcCIA1n2MOXO1kk9hkW82XUCC0uj0xlWf42443U9I
gs8R75ITPMdjtovLTytkx9aP4XTGMBM90CCtWyzfsIfT3dEXkANLahFfAK0Y6zdR
J2BdWCa74hhfvPYWoeC6pEOw+M3gpgbFYK3ZeNhem0hjby5a8e9R/FJ5pkwMe5DZ
JwOyj3PnRlOq48Px4BD887F5RBA94MlNGhKvAeCY6Oi59o5UDVrG5NMoMEFuBu7n
Msz/ClvjkYOkxk0/ecGXVKO8m3DtLVIX93GRpTvnBYfux2TlCwOPkwiej0cjzS3Q
Wly6Plc31U7Xc6mVWG+TeoOV6DT1jhUAo2AzVVCh8DkqOguVytbH1WOOTsW4qPS2
PdN+HEuRnb4USnHBI6twu2K2yDMtnf/CS071tmHxAbtO3uka/d8ZQtN2NtWupTUl
kBauErESPKhtxboMtLKMc3ILx+w/MRnj84KiPdA2NoTQIVejv38JVxFdWL0kUKs/
R0ELi17upeBeqLHd6qOBBFSNtFYUu/lEiCphTOFHK2GVHJIOUN86nFj9DbobwAtw
978VIhuWNI9DaM2V9QnaJFknTaDq0naI6EEhNIJHv26KbkKP5hZ+eCpB5rSW0qmP
DkwUrwp6pvH+BTIHI7RXIKjvRO8xT8zXzMJTdBO/cnVw60xdZrAg0S39SYetxJ0f
KfB7aDHHBbYmFpn0iHQU8c+UQakhL48j5sAvQd01BABox4Wtr2cvETGzuSB6/ZGs
NvB9dHMyB+jUJFEpkaNryvCdW4WFem2m8ZnGYahnrKvCpA7jVQeZaOwk0TpTbDOk
Wg36sxIFrKbrlftoEX+AaZ2cwUaruJHEy0QuvpoeNZJK0fMgJHwHGGCsgIFpHUXK
d3Vnaiw0LNXv5h3dlf604BJ59kPl5S5OuFNWdAhekibhfPjls38z2ZtdD1SHfsH+
ppr0XjqtteWUcoN9g9yY6LN2sM2hQzEQ6fmau7ob/DrJw/0xtxadP2Hl5k2Fu8st
noYjvZkT3ttNKkbCWfMh7B0VabIanFbZsqnH6lzVkq/GRcin9aRdXUtp2LSu/QRB
+AidVerWzW/RnpngJHPD9OoJzMfNQD7ygnbWYrQXYT3Iq3icdRVB2kDmcPl3YGU9
NVZW+Oa8KzPDDHedGiNFNdmU0oczO81dDlSzDinPH6uXNzqooDksY4XvjAyH5fbO
nCOtiM0d+8/AGSWmj+fdWoWGdeldOy/zGieOb3LtK0+u4w0jpNdUfvdxcknAKaTz
DZgp6xOfDIkcyFQY84zQp9/S+enI1PDSjyl7P7kghGGTCPArbcphAq3veo99dO2V
bgmRxEukHNywMPV5waX40KDMNNebqkX4Ua4PtlD4FgU6ajNsXhskDBqJ0fJZnqol
NvFDisLtMha3JmX/A5td2JTLdEiauNVoqlPu/YgN2DrgNpEp69wMbPxtVQtTTV4J
hl9/Do56gd/8tyHqW+xMpgpb0+q+nerF24irGbxsWUI7VUc3+n0oWC+rKd+gt+5I
MaO3BbI4cqkloK7xy3OfISg0ukIGO1uF/2KNLH3t+3sjI3NvKLRmHir7XIe45pB4
JhXaB7a6Xs5pfIKPD8MqloyDV+kRAqi4rRPLakfi5H8u2YsWnoL3vAJh0voFyKfr
Xh/NVk1Q7FIbHfmzKJUIq3kkEDoOvE1BsRUa+NRvulMDtqToS3+pOMD9wJTKol0h
9Tf8IsbUTVx7hUu74atRfY1jRZQOZ6UJp23RSuofh4mguebgCp9ALKmKNIEC80CC
GIZAg7eNVaM4wIEmPmLPe3JdE5EPEkWb51eTD+pCPv4YCjmYjwCYTUI1bByeNG+7
7vrS7GPx/N06VF5XDUg/OcI0j6TXDv4E38YRMTQgkYoGiGs53VOtI5+KYWm+/9DK
4OiOVhw6GWINU6wCz6Z5rNKW5U0j71M4X/nWtp+D+A9h+BiER1KDwIJtDBTShfsv
N9vxtCUiZYPwfpQlWqiYxlse284Fs56jRKCtvaDD3bRcwaHeCKtmHYi5RTE/Ogjw
IA0EOUn0aN4tC76kmLbZS/zuJV2PAYhMNSIy0DiGjkDf8SMiMjMS9hliGXRbVxW4
GjowXjF8pZtM2Ih2LnadsFLVnV+yj0wupmzD+p8qyk6Ow/9M4dDviPXIq7opQ76q
zNiEUPDwKfOsNKDBscD7bt2oLQJgelcEGdylI4GdtYVZO3P5ZTZQ2RE1C60mFUaY
v8EdeafcRD/dH8wRGfi5Fk/vfSoV8vLSbUIqvDQiedEQKtwto7wxKruGAfxCOybx
p7sMMzDPG55BawFRNIesVeVudL8Tc33FG4/lFlzpy9EMCzZIRFAiEW1BJ6TBOVGJ
33Z96QLMrOIMQufSIJpB+ab75jDwdk+o2axH30YWYLQhgaBlgWWJzyutXoAd2M7r
vufkJOBB/jivSYco5GT+ZBYuQlW5LigFBZPTdG03OKMM/spM00NdX9ko2vY7EYz6
3cuVxikQSH8E30XZ3zAaisjg/BnlStAUX7CO8kCuBr9eJjWsrbX8YshxtbekZR2P
Rj45fWViQoNb016FWRtoHCygPZZN1PPSLzZA1N+4dHFzihww453t90pi2UIAPpPU
QoXYVB8XGDeZDPp/YztPkenpVJZxD8UdneBYHgrPZpnFe/ZdfaJz86Jt0e7eFBIJ
lrw+T6htl8lVNSTuk2X3Os6AuA0fK6bUOHX5KAYDbzTu/HsJw3j+yChMtbdXzFUU
np2rfOpOykkPAPBoYpGZkJX1QGH5NgtIA2NjZ8GT5SW5v0ZOYBHb9OnSTUtvFY8J
Ev1BuwEmuVCTrDn2hUztPKYp4e8TEZ0vkbHcvmVgPdSTrqKylU8efB7m+PTMJodx
+fEkgU3p4WKfjWjhI13x+VSXmqtNybGI2V7dmI7zfhgbwMcSfAxQXVJgzmS/VLnp
9CZT/S5Y0jJf50Vc/oRywgNtdzu5LS6+9z9GOi1qXd0NwhM3oaH065+exOl0pOL7
NFVOShT4CCLicGWwE6a0k0AY5DnQUZDVk8VijZ/ut6SNFFw6fDx7EAI/TdKtkb+0
AHM1wQRXUv/pKSxVZkbMPSRhLOneAhmoe0SxwMr903vwNijWbxMwyJkAVQjiV7/r
ntIQSUZRTQITz3bJxyGURq3YKbngAh4BJ5eyAF9ILH0EeT95RqiJjB5jtO3gH7Za
0XOYqQOSzE1f/CEJCtMEpDXUQ4xO2oWCeRi6qqqWIqaPuWx/7CG2mz7qH5+38HWp
JTgHB2ePfiUFJyfYUIIQkrE+DQHnL0ec9QnoZBrgKb7xbWiSuZ9wHZVPPDNfS57X
xudFp1VYDMKXIzr3iHc4nJf74MF2qUu79DnM14zfgg4pevHlEG4SXHjFcjosedGd
t/DltIIlJq8/iPkUIDKWU3ICjgmlHUqId1GyTvnbGksl340wfvOEkf3MykvfVD0x
jN13Hehq6y25sUM1tZ0oseA9Xvp5hVF3rQw1GpH2hdua4QodBKenooshI8xTE6jn
aczEtrAb44Erh1Cv15eZxy3VB0LZEnGHJ0Ef4o4LpSuxX84CQUCmV5u9D6xXAhmp
M9keBJLaTASY1pt2/W/PolZCdJDYYeGTDWcSeWzbHtbuEbk3GTt8H0wGXzLaD4/O
e9izdDPPpnkuneMuUHwd1a7juEfajRbnMKcLML3LcSg0oyxBHHNFh5uc6PnPp4g1
29gtbp4fXLACF7if+GSKIMQ2zFvWVeo4TJZoGJ+Tk2MBvrd++J07NpzT7ItF2Cr4
hX/8ca1Tx5aw77fem2it2VZJtULOYL7BeIRadgjhtXQCxFRFDgP1G2p6SrmdEfv8
0mJIAL4iOQZN3iATzuSMOcNPlVtLJgEQEA9z5a5XZSoLC8jrFrtrxD2STUQVcHaH
p8YgO1wDQVrLr9rdBBmJneaUxQ6yArV8jThF4uNIS+3LDQU+Dp7+swmGpY0ONqLM
/K6U3UFMKrZmoYEDTfMyHjXLuKOJ+XoDou4dCEAkhQhE9OM8fPsbtGZyd/SGZBf1
/ZevNMuWA8p8oVVdJCi858+iYsaAmjR+1WchdB5pRyLAlolod3qA4s3e+k+2pVFN
421BGYM2dhzaxf7+Z+RSuu9OLdbEhhXF45O0fHldMSfoTXhdLl2EoyKQUSJr674y
j6xMpi2JUNhgpSFK2vJ1mWTAdz0w+DqEsmkBgn524rMs2V7NTA+RFpy2o7G+ddwr
jAltcmfvEI05MP8tpEZP49fOq+8mmz9+ooMNC5qcGXEY8C7cgJNY8GaODdt+8914
UCbVtHxuBO7wP3msLOIXmWGG4l0Prt+zKC3GlDS87x8LieE4skvc/3hpiERpZe+N
Ix2S6Zk+SKFcR7nniT25r6vuIRWsPsqQ4sBnEU6jQX2KQDtf8pHbomE5QR2Dp6G5
3fRwlU9ILGS2I+tIccIffZoA5xWs8mlkC+chCBuIUYDDW6VbMR7xdpa+pMRI99k6
U0BNWWoN8bWs+qRcz0fieTAHlfsHGeMDQZm5lCM1efQmcDNPtuVpygJxq0xGeWh1
r3GIhhRjdKemSMdwJDfQjJgDqtPlKTx0t5pNjcuI2+lMDnuQH5ZEAuQshnsy3qWP
H5k7RgXAB4fCsXBxPhGiCdAQLtqBviMAMuwezyZj+f5rcZCkXThGB6tYUpj+MBm7
bhWIzvHpAPaFyYFs0UrWbM8NdRdBXtEWEA3HrnL28Zt9fCpv7/iZ4MduY/8qBumz
9Ram2uD62eG6MUoPn1QVhYL4Qf6M+j/DOTBQC7kNl56zrijaehJaNAyq6qGo4QuM
gXttsIpYph99MBqvkO3Ay66x6qCTaEGZV+BFpHTkcjHHH7vSDHTaDSkjxdjRmTge
ApyfGF0ewuHkAKKv2o6gqd39HynfT873sPlxMJxX84ZVLQ7tV0nGflA7qVNSoTCZ
krHPPTjb67xJepJ/+OV2FEksA45pcE7IBFfd14SYyQzZ072feQ98DeVVqq9msTfr
ZqzZtPOoHkk6t6t+lSxkairT4jQL714xIg4xRdAhtiMa3cP4yoC/9VzpBL1G0Hdy
nZQqbaSijCHApr6swfXpN5GX3gXR7AdcfnPrpl/su/sH4uk5gYBJwEqc2r84DLH6
k776D0DIKlYf/sTt7pmOHowKzMCetGe+cS8FlfOXeP0qA3W42bSTSc/NGGSxI5ke
9za6fxXRFyyCc2+fj6qsqA==
`pragma protect end_protected
