// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
UnPa98K3L+GZZn6euev6tzr7wpR1Ix8hvvrmSyh3a8d51GYjJELWYeQat5scvKQ0MnrTJa5LdqLH
7K3BskgR/yEJg6gZ3b4L6X8mqYQgXqPv0A9jKnFZ9pF/aPDeDLpypIsvDfYHEBrGv67Pn8IwfufN
wJsSc33UBy1uqdGiElDoJSGKu1thamw7cGj/C3wpuMi5ppr/maeFA9QYhAySII9KX4Q33EHMnOXj
gT8/r7H+1tJSgSCDdN7Dws1pq9neyIeEJgEhdn66LF6p6+XWEfjgzrKU3WFVjnaj32rDog/ccGTa
lj0mrAhQbf2t28qAemyO5KDEW2wD1GJpi9gR0Q==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
3YcfnP7j5EbyMoTY71ZkNvCrIxxSa57k4Qt/wjvUIs1tWyjjUQBX0jMcj046GuKDKjr8yrlnQCgH
lFj4f9nyQUYgaN7ZxFGjbKMxgdnKAmVLLf5chkSnAEJDJVLtN3kov21n8vdLhImsV83CDNNKrUqq
Katdrlr5QJr64+NWZGXk/ffISCcgdGxoBYjL3LB/BR6dFheGgtpm4Ii492njJBXHwXk53jKm4cGP
EIMACT3fFVCG3pPHOzE8+BVbjcONQ1jMV+8BN1ULj39+/4OrTE/PuyYe7psdaHu/vWLouOp/J6Cy
RvZCTT/AS8BXV5LMkY2U3DqGSetVzk4uMJ1aXiiQUt9QvkdMZpb2pWoCK3ymjXbiyOUzyVZjFtL2
ASB0WpJVnO3qpFvG8zPb6X4L6M/yl2i+4dp/sifOuSjy1gUCLbRBvCl5fO12UNreyXoWwUy9Z2im
f9mnvYCDpBMcNgx+56dyioXD8upb1c6SI0ZLr7Z9fDcRfY7v0o3Tsf09T5ZDPFfMpAtDPX7k4/7x
emmCBoz85qUnrzqJa4AOaoKD5bGVA8MbJu52P+hgxzT13m1yNh01wKabPsE85KMGWPdaYV7YDebs
KECrBzjYiHvDYjsssB4/3lAlu/9udNLKUGHTDzDDOLdrmBj/TM9toUNmcSx56KwfwX1q1zMrbUo7
rhfejgwrfbimFCIocejXhOPdx2qFWeOfHp2bj+nb1AfjjqMDmQsJme2of9y/J9fCLMbiI68lEVH4
P3kiriocUMIGMpJ+21Xz/ual1j4EKxghAS5Su8Pj01zTPYsPxJKGY8eKl5DBlWw1AzkaSj8i9fQv
2/o3D40rc3xqRKS4Oqeq39Fe2sh1Kxn6r70LT2ehfFWS1sYziADZzg9twuuEnIeImWUD4R1FQwsK
7IJ137iS9Ddbtr+E0rOQJLR9x2H1V6lx1oy2fwvLuxJYhFM8dTRd7gj36yNCK6sSztPNGtbZL/z8
LDl1wTqV0bfKmVD+HxOCpjQkHDkTjJHkzLiaC9zuQc7GrNWoQYFvC4noYfa28+WYg4UeE3nCAR6q
CBsaFPilFZRFe+17+X8n8F+QrhGSAfklc3KkTXbe8VE4nye82Mqlv8Ie/9eiYe6lBQ24ZS+s2gcv
pX5t9k6CCAlnDrmdmnt/WshLMm3+TdnW73HVkofbq/UdK8QF9j/VSjcy4n2zxnTFL8ORusGlnMYQ
de5GK0RGRVGz++uxOxPEmVNPUpWHH6dxAvIFbfRSsNeqey9jAYuOkrD828kFp3m93JrpYXhZJWPG
bjgRQS2DqVM/B7CuZF3UgzY8cTCWzgjLBiH7AuccVoXJrMkVJEyOCk7RrJFEJ5UF11QefEAD7Liq
5BuMfQnY3HVlE10v9ZYbtuWgtz7T59Uke0AvhgdXlaSm3MnjZyHhSxAySiYD6vZ70CF9vrLuXyMR
ZzBiE64VjodpTJg7xL1xKXMbSDcxFbiGU5VZ/MACpVUPqf9vkGc/TyY8gooSiaD4JdCn/sgmMfw8
RgLVizjWv3huTFDgLTKvI5AJmECXyl+Ec6w5anKkpw01qn86MS3nVP9KhcG2Jn1z8s3aS8PzZMxe
guVOw8Vg2OUIa655emCNKtG/QuXVVb187Bzm65bNph4imOQQFcYu7HMVrv+7jPd4D1yFU53zMkGK
iSTxP2fpAprvDD/E4RwpJQhMHqYqjcCPorLyyDuqU9Zmsxk1ESuZByRfhMJ4CPXoMumEZSS5ZWRw
LOH8lzKPhKjZk55wMbKT+T554sxL4PzEZ04tbXl8Hv8ojJc4jqG/LcukOGmSFmqNfKDgqLyOWQJM
fHMyIgbfhMYP2QSe1AFu48W+1KYC3ugSl82sOzRiIq7XrGGtvT0RISfFr1CyrioTtPrLaBBbwbI0
4/P0QOugQypWbaT13wcOxJsAoJyYk4VCiSng+1d2Rz1tZ3UoLgRcf1HpnI0JiZgYtsXPgK7+IA+O
Dz6g/2uo/xz5jGvus7OB7VPhMGMPzNWgBY97ZCuRwSpdILmAdPDezxgeguPpQaOp4cedzJoabJ6s
WuYrMByz9PFbIYWioxPB/x1Cbq3xG0Rr+X/hCb4zAnDNMTLn4jMryCgqBV9GKaK7wBbov72NfBk9
ZTwb1fyLXev4uBPCX47rC0y3WiucrbqGEcnayyuVmnoclLoozRhADeDsX6dpWQV14O2mrBYXbwhT
aLNZKJwmrE5lSGGFeofR4HSf2yKmydZwNCHys0vzwXZNm9lMJK3CI7Zpimyij+Pnwkuwwx8NkLji
LCeNnrbw7dLDVpFbHiEnfyVToSYPpZzY+DSVGHMlmXfs1+ejAN0qJV+7FnG9FaVuRGPGvqC4f1RX
P+/0vBAwayOzfvSeaqIY+fMMhtEzscAUVanXVKOYzva5t6ef4RNGGvJ+hibNM3B2CnOziAV4ahy3
oxSPzuLKaEWY+8fsmAL28Fk+2jrDlY5yQQOsYgduL7oOS8PC1eJ9kG4BRA6LAph4MncMhOqPjI6w
zbzAhDR5TT8eGhm9Cw/vSxQbF8dZVayJv7wlQ5yTY6YKUfGOEfm9D9aBF22MWPmlen1LG09q3TZr
XsrIUKznzzlOkvTQ8VhFWPzWpJ1+cB8toqZH2zFJDybg3Ij4dVSzgBfCMlPfD5rs2B/+Ry1Ow8XD
QWwy0ZMNfqo+KROs24uDUdDCnFB/VAP7qPKCR9912+OnOjhcFz4pXk1Imv66jO1/5ptxD/SgB1wi
9A2KGc3CWLlYjlj/pJgmRzSWieOFxqecoToa2RYcssJV8eBN5hZnXZAZF2JlQGSSW2uSUFMgNpGO
v56GkPBH4uBlIDBHNfG3jOY+yGt1ZxTv8HzPzRUEYkCwzi+xPLL8lYa4u2s76vC/AwsCqLsVksIV
nWxpDswGB5P5dWvyEgPYpMM6TlAQfINmwqnRzf7PjiyzTWtjgOpLHufcNyzB4ilwExsC+lC2oFWt
vfmPBp1zxLAUB63p7OQjBn5j4L3H4bT2o3RAXvkTKJa0jsTxCQ8JIGMxJN7QUpFNriE7ApH2E0JG
3qkKAcLrGfiaHqbJrcbpp/OkgMn3lceIsEVlZFK/pWtLJzmJnE9T+oNiSdxOz7zx0I/3yrfE6/up
DW0ECgVLsjtGE8GPA8N/qHBkJ/3ezWQ4LjHUHsIhoayxB/tTwCu1i+2KsBMMCyvEnvASNgVASIky
DlB/CbwxZDU8MvSPXdNgcZXEdkFZL+GZolrLuaHRJ1xOg3wcK+LHFODhJTB95TOi+ZQBNObWpKi4
wekPWckZR+aNdsvfDgAiQqP51S7SHDaV/IZUmB4PSNYyn077JPF50nsdPM+h7z9pCHJW4w98t2aL
TFHmXUwYhk6+kv5a6wS0Hkl7WiTZHtXpJgLJNfY+5QidcMjYaW3XuYDibhj0XxXZre2yBtEKNB20
8r8gci+VAIyqqmnku+8jEWf8VKGL1AARVjRnV4ENnVVlSsCLnLnVxwqhYyxc2KPVrg9jt4YzHUf3
LWmKBsGAN/zhMarr3JLLCMX+AG/IO5VnMC+HiNLGTY3qvegBzYhu1qgMP5WYX1SLFcPkaorSqzpn
5l57Ls35DzuoJm93tTYU5uIGqzBYcZJnyYoL3zbDvP3d/QQE6yVcaZnPKTT+HKo+h89R3t7wnBmB
MehD82Fdmwjf8XR4iggjmImmB9k1hTxIaRu0hgV1IHDFds7SWVOCRWOw+RCGXD2Ff4YJhuq8c69t
xRNXCEsTELWBvXL8L+83yABGN0W6P/Pcl1WB89i7VMBzfQRZsy4LuNl6CRyvjpGhCuwNovYeGPFJ
wF4GaKMwVjSA8IhcgtNK1f+hbh6sEdyW7hegHuk1w0/XBHj2YGpAYLirpxETdQaARNk3DB1D3Wnb
gRDfgqXI5Zy6NpfiD3XHIuukPEnegGBcH/xbYP+X2zQjgHB4NpcIh05OgYI69PwtMxE7Wuydz9UO
Q4QsD2Rf++bBcioxhqTkds/qQxkp93BIS6nJnlHupCeOmQX9KchLnIi2Hd7eS3C4NezSVWeJNXak
5y4YTTAJAcTtkUnT+pnB/Kay+xiWuzLYJaoTW7e0sMlILrRxWnkcjt+mSVwmfs8awSjoa87F3Wep
S54XEBnSmEfVUotE+49hhwsh/q5hPdi/6FU/YyCJvxIACn05R8yQ0I5JCGmibe/q+d3gh6GCdDeE
csjfhpl9sE54DukWYjVaaNpvgg573c8SrJFarF95J+EyP3QrfmnnRWUl2Z6pvBpYx2dHwh6SIuYK
0Woh5Tdj0sko6fjFBS6ITb5pE6SdifYOFPwOBPOB7xAKxS3j4+zp3kLl9r1oVpohDkbn4bwwpz2T
siYi7plovPaoU0Y4QHM/mlaJ59uzXYk3YUQHy3qw79ATABPnnD31zDi8keUUfurG2EeDAL0ooxrC
K+qkuxDQp5n3Bg7lFKAguQxNQeUmdAbGumyYht07cEPGy5e+J7DkvZnSLIFZc6pdq0JfYQzHctGN
SgMlD9pAdLDm5H55ht7Do5ERd7hmhyoaLKBdfqLEZg3JQggrpTGkFmgwPT7WV5jNSgytrFAyT6W0
bB/0/SnCaqKxQfwfhhQFL8QtP+gKnJLalmz4JcjEqrgqRVQ0l1ty1H8UNOdopjFnuC4JxrZ9Cgbz
c8lezErRkm/EVREo5+l4HCVWSQo+PCoeVfuyvr4vfy1zNpgmQ+FGHcjI+D6i5KIDj9Nacrw11XWR
UgGOHa0Dv4o93RLnviQhRjntmwtXUDFGpq4KLNuZmi0qKhKG38bWfrSK457tO+MZOTdLH3VnQmE8
KK8thyAd8OX5Fj9XHtzbalAxUE0VDgtyvm6qM+8/wCNBG4FAQePBhtB/DqpU/WQBUUYxNHWy4ogz
Y+U6pif1MTy7dx4o9iWjmNosi0VkmfCks6k3fTTwI1wgIXhh9PgEq9kpkTk22RdWpeuO7XbMhYiy
Sbb8WzZGXAG9hA7ZgYJ+IzR9RaRSM/mK+00H599x+dCxf5fypzpxyH/x66sDyN9icTk+HZ8reXoc
7+4f98QGWazp1U4sAf6dKTA1iSj3vla5p+MjNcqkiEqzaQ4rOu1rvQT00TYiWAeOhJjP6AtyMEZw
+RHOVNlJAYnG1E+yUl+bVYQr8eX786bYatPmLd6rhL2KauG1U7+YYOUT+aAp84Qcib3BC9ffRdh5
2+OAClakKmmm6f4+qAPuNeH0Z68wp6Qz0mZjmTUoBe2+QNFwIwW+hyjGNValtZyNvRo0381LSyfQ
3WuWrMBRzw27tYOmcpcaY3cxiQf6Gt23IleMJYClpsUbhTiwG52uC+Jx5JYCIrsFzaWKHARFONaL
10AxOMRBlWg3u/MJrUAOZlWh8u/cWXwHv+IOZWS2XC/zmrPAtDV6kzSejrM1Ndoo8VaqVjMULlDl
2UEJOQARR7oXEWqgE2wJMVk+oK4BQXMyIelIobcjqQOLa+Mf7l5ks4oLZu1045+/LhB7+zCARkmF
QsPawSM6bT3ZkxgED6JvlWFUedXAV43YAPz1byNYjxIQJdR17Fzd3Sma0sb/eYjwISL7ale3V9oz
NXV74rIqUdbEk2qKvnJ0s9AkFC39ABEQIglL2RVJ9IsSU2zTtUroTDnX8lKMyA/a9qDZoLGwDeuj
RAWBDW72+bxRnoVGJFq7v1rbXphaH58O+nkgLb629HLka41YDVdWPQQGPw5lHUEgcm0O9YuL6JPM
XFw0AGSh38y/BmtYemYlTTsFN9IwzXCvxTyQdTsTNqQs8wvmjv7gbB/4eZ51b4HtuddWkcN8a7GS
iOpQfhihQAYqwTtbtEibibZDx7QDPBgVROGc8DBdLPlWPyyuWz2XC1SnGF+i6W5JToq3+PwgLbXq
PQRZsPbG+FxwJpJeidEV+U92jdzLrUo11TmHLXMWS9yZB5LxyagjFdf0ZUH1711EDRUPGU6+JcaY
YjTRI3zTzo0VoDUtr9j+8oeb9CJS1QSmbh+wC1tWzkZBEP89UlUKx3OjENlBDvWogu3lvykq1KSJ
VlpRcUtR7ABHfnqVoXepv5SeYbhXfzbQSjYm5caPBUWwjTxAq3eZoOAJXA6ufqG0hdJ4m/aLKm6g
p0RJ56refmFDtXcL1e3/+xn3s51OKEVfJX8KaperGh+BzuBq0Izboh4hqFvdvE6tm5CLXErAHocT
zjjG40CEv0kCKjGLS8JyxQ90NP8Alx6q11b+Jd7qH+iFVhVhFFElTk+zE+QOy0j76Cc/1926BaFG
pG+Xu8nOEO+6sHYwhxRDGh6jrNZF5Pky3Fuo2Fne0f4GECkLbByodmdgKQQX3c30WGOInOMgi6jc
mkLdPSpUyq4C9r7nX0stMbDGk7D3AniWRCMrJSHw16SrEsranjnG/8LxbwEaNKzVV52ayvTRj+2T
1JcBjnR2OKMHVXg3qEFkGGaTZmH/EIUVYAIiPRtYz7R3U2Cjl9ZH4zT+HMFpQZHYt5spRahWR/0T
z9S7N6nnVOBtFpwGZDpbwsPlKgeTyP/0VYIO7+fmGrekbmeWsPXMBzswavelpbHTSd9CpS+yC36F
enr+onODGhBdF6BKxknLLVCF4g8pyiGACPtb/u87fY7WZ8o2CUv/yrxu1ar1DptT5amqbqTGgmIi
BPBQmDC4xKAl5Hrw0Mxf0RKlC0d7nnp25N8CwQMKNN9nN1jQLuj5yPHWkj58hd/XSFU10aM0YZPu
/yQ00L0MlO9Hbd33gbndEPNG0yJmKoMNFy06kl16seh3A6zfb/Ye/tSPYkxY9InY4+GDJCgwiwTH
zNPFGsISRjHDGa8T5q8ZMmT8iGa+NuQbFH9ZB80oBIggGm+1gP4zku+m0KmwZmQW8iBzLFSrwV6L
jD64hcBVLMi9iJufE+sPH0LUG/mFAAhbOB0+mda6F4fOL/ycxqualwSWMh+RyNozop1NIgBHrj86
5FFz0boQJfcAVAOgqudfdwNFXPW1GLAmX/vr5sTEd6+Y77V2mdAfE+5sSTUu2SYymvDbq8JSp1Ny
sB9oD3XFe58/MZyW+cG0S1rBYvDLYo3InlUTTW0wETOud79jAPtly69q6OxNr/AWOOdENYRqdwna
O4e+RHGSmxYQ1zo9+ll//v7wjXDJiWBa0oZVc0UZ8WykFendfH4gYGv6uPPokwuqY8zgxaGha+mT
OjRLl1jHXL2t1fNEedk8/Z7MVyYOBQoU4LNR2r1q4XhqL5GYXfedGq3LSGid6r1/PXVNjJNA4+gd
MoJBQd6XdoXas3iMqzDIEokdDmYRNTR5d4mP4W0gyO9ioiuAv12VsqvBBrRPhoZ3n3LOGC9BUebR
btOMTED/J9tcrRPVNChrmkf1uEuQvwG63Xn7iXhCfGX3X4ST+w3i9MgMt2T7yy1pPnb2ZaO1A6t+
k7e/hHIZDzKj9m/ZxfqSWDdc1zjWf0N1eSS/gz34mTlWzM/jwpibdFIiv9JV3flY2LsViwV6Zt96
Ykchzq3yHEzagAJj1f8gxtL1DFoO8gqa+psxefrJQ1ZO/liXIJ8m9MGoJCOCdYY744AWd8qzV4PH
IRQC5eVlh18pYqlxAwPnKcWyAr45K0Q/cAAOFguiBdMDDHbVxcnDNPkv2CQ6Osk9uTMyj0jLsTJt
nCYs0+qAb9FVR0dL/l/Kp+4eygS5GyTo5BK64UbQm5RTyu53ga5MpqYb8LGQHT+8M/rDAXYc6eyh
+Hy7rrPA3uUxPb9+veZl7K72nj0HJJ7iPnrwfY5C/n56vqDpPGS5M2dsc+MY4u7KkHZMiewZA3dd
49FNoLC54ay7Z6ih2EWK0cENotHRMecArIelklIRo+xc4Uu/Qcw8zmw9n7x5giFnlSklsoHHyN8W
l1RiVst0yprJ8gwMrLuQUsf+RnUSMRjH/0+yFfTG1lUff0/e4nTgTftvxRZeXMoNS+j7WLoiUnrL
VK08HlbXvAyBENCeDEqOGTowgC/pDOOGPWqWuwpMT87X9DqNGYhx4xeLBt8kj2lIrozRZbWhVv1A
+PSQX+vN8wuQe4au/BugqiyORLpvvczzadm+KcIYm/Wid00IkoJRAF239avMvp5XzaIB9ogs2yGQ
IXI196DBJwV1uEu7X9MgePUzXDLgR8fljeBFCu61+L6wHeg1C+z0A/1hopkauayBgtIo7DLyJGf5
0cpkh7bkZpcPh1gtF1dXZRul6BNPnDbVYyz+5/6zHgOrMlOe+aioPNJSmaOHdTtkENiDbM6D1zGx
as30PtWrQZN18TN8MtcqWP3X23O7+XmQos47x4xIjKWW11xjNLK/pEONWnUjIgfb/wa8gJFXdtdq
aG+2IXZZ6PQYh9uQUEkHASEue/B5pvUXkSYw6Yj3oKH4HLLvfTezCUqv0BdB9mffLTZIqq9XX8X6
AOoaVl+dt06+dlbsdApq79agywfGXlxTa50nHJNjhVnR3f4NYlRYZFyNHdM1Yio8rbMbPos9VQ6K
z4dl9z5q4it3c5hst8hl6thJYMkdIfCfsJmNDlnFdp/yQSz+Slsghd25uHuoLjOM/ZdFL3AGAP63
zHbw+z1dsrWmAboKi5GIiFyC9Kt6jmlqgBKbJtEJHNmcLiO2t8Xd7EusVOl8HRhkQTuCAHXsDxNY
bHZ6gA4bsXCrXH7935rnV5EZDpGFJufoBPkHH7U3q+oSYwLKCqazE3rL4f9CPA65eQ1QGQlQSPPb
IF8Mwbt1jPLCQKBOyK7Jrlwz8L6Y3P/k3jW8v3OUvYUtsRpvAcIg/Du6C+I4p162DNP0HaUkx3f8
mnmoQDU7lwWypgfkRZ47dTxwoQPU8Ge28DtWNZD/KRPnHES80WSZxtN57EsuOVd5AcrrYFwXKwCg
SJtQgYpNxyT8tw1IywoszIqTlF/HvHA7aalvnxIT7Y8wcdGEYCpxfhGvZIdlT1OaSuRvFlartjq+
WpvGtDLhhIkuNdmZuNKJcOgIiCyOENDz00hTotLy1lsF90SP+M2VNC0TlCfkaTQJwYZ7eyVRDjt6
Ll0XMZv0toAzJZu/A6aVYD+GP6ZQcXjFW4fC8tviHHOWTVtj/t1b61DCksPOka0C6dwGtkdzLNXD
1Wjg5qPWMmpq2GB4JlneqWI0lsWTc6VOiPTn78t6ux/EXYZon28hdIjwPYzw4x4hbIIocTLDLnKc
510bpaFPQsopWUsVmz4yldmnywEZeuozu9ujoE/WJPdtAlZe4Pfzu2SoOPrPKTunTqXcoFqV2q/+
TLEqwYPtI8l66MiezoOtsvCYV26snQoyQSP/UIuGh8147KYzG1DA+JqQeESGCvAJs4CIDLSnZPGz
jSzPfsZrW1J3aIO8f6eNj4/oUAsNyNDiikIsOwtQcEqns8BLtVlBhYgvzj+bjwOm7DM8YZROiQ99
XA92SZrmAoHPY2fMoZW/HzpbeDBUYCcaFMg2CwuIYtI2OeEl5vCzV/ZjC4hNs/ecZm85CwcVSP9t
X7q8Es719Sn09pKREU8XfPWNylqYPbb9OheaoA3Y4aYNK9cSCRaMUBtgrT9GwOCy69GtkYbE+Crn
owoWAuXP/A6oZ5qsdQUbcjMjBLZgsC/SHhzf4ves5hdAs3KlEdRiwgjS3M2yQwDhxkKUwvA1R10B
i4tyuQsqkO3h72WDq+bk+9ItFQWiCkpg1cz68JlxiVcZQ9hLmhW2IElrhC26JqLqS2uNekDvN8/q
djZL2BZNXMf6EKqi1Z9E1bGLnAvfoeoYodXHkV0j9DvhR2wkZW+uW7Ojde7CJEUmRyTzoHl8cZ5B
wSGS9oH7CBM7aVQ6OCsgtK0Sn4+v2F87tm0ifqOwM4PnLcCXPuFow9vgQbEks6bn3djEROhT01YD
YRbKMlYXgTkfhMsR+vQtSteAbR7ACqgnc16huPOz9fD+5H9jjziMsMsr09Z2W+zhbhX+4QDM4uie
NPOPhlDc8OErnZ8toys5wXR4GsBPQzEFNt1UqSoW2rSIJ1QIvO8AbBcesxgwDnYtvAhpqan3CvMz
4RA5CF41h9mNmcD58p0PyTQ3iNZWp4TbbjsWEbQNuaZu9DTb/lmO91VCVlWFB3LjywRlmTlkpR2x
91HoJuQWbi6xa9iNqvKXBvfOzWbWoU4uWpuekGUK18p/rHkNHMjpVbYNnzSaYM0FjxjVEeaBmWKh
ehQrARCPAxz9GHt1edbWTgXRqoN9xowkjGWwkpic6UtlCfdueEJXRuKRDLAOdxg8I7WL19rd6pww
M482Zm5SdisiNOFjgZgtYy3P69DQlI+l4n5GAHtjT10nMEaTefr52bOQM+lo+BzSgQ2V62IZ8hzi
hEDUXFh4wmdrJGuDmkyHKk6uyHKmTH4T03oX6zy1ZNgBTFsQCq0yr8cPPjOQxaF0tSV+mPZcloiC
gOPGjR6Cx5QDgU367MHz8VeNIYt9igQpw9gjvEQ49VEdYuRYOYBJgz1md4bWcTgCDiAdrPjpUlTu
itv8lpJkth55WHF8mB3qJL66LbTW/V37azrHdynTcuiBMKNBrA754GT/d72rCzwe2oGxQCtzYIT7
YAFbjZwHyDuVfZMNJoEmAIlkJ3tbcjPgV1yztjXOG9xbRzxoS272idZmuSUuojzVkC1F0WKMenQI
qFZTQAurnEha420Qg+5dqqjh1bp0lJITxCJi63sRS+Z8G/VX3xeDQB4DDy4/rG/FJBoOp0fr5qzK
Bbdit0CGBztWK12HMcx0RnsE721YF0IZ3IJzENgE2bNcXu5U/OD0buAnLz1PXKMG/gCCesZpGvMG
aVSTepgtNXxaGaT3oXiG2YYR59TEmHmIMXpLdJBHMlDSmuDG96XaXGAJ7iSJoWzTeejm5VRE7AI9
OVP3ETZEOkAnJN8Dqieo0ruZJLqtalShFbSAIa9uR2Byq1LEXXA4cNTcyv/Pc6h/Vu0Xry185BP+
czfvcLG0Hk3mbgNl5827UztZrdhm7CxeZO19xwSG30VBdu65BxY3LkAo6l3nXjfm2fZfQixP7Nqj
FUHlYh9h76C5Ds51WUrdssJRRU1aLbpuneoloBV58c2MyAPVSy3hOsxhf5Dm0ZQM09bGcgK/D6oC
NXXgtQn3QEek7w7hT+y5+WuDwtv7cHK1/tnMoUB3/Pg+DfA/SeN2TS1jHwvuYrNARFBONSx4/jav
jzG0CzGvNd4XaJRVBS5X1NzWRCFraR/StBRVGnsjT7dZ5TVc5sBepxYiwgupSciLudzVisb5t2oq
XLGjdW4hfu1Q2kFkaBC5/+OHGbqINaFariRBp/8Ux3Zo1TZphWEr+pOn8xP6SNxu3XjeTfroB78N
Gkz54UlJxCRT9eMuC7TdWR7g1VujYbLduZ5tM8AHoNDe9uxo40djPWT+IxYupJHlGBseOT0zesYo
pPjBVFHgVmJVyN2px2KHNHuMEkyYB5R0+F+LEwvhe11KZyIxeBVCxmywVx97OM846FItuaiG7Hxh
6rOkvPgsR/+n9FQb4OqzR+d6empQy1bp44XPWU/2O8CeT+Ivfoq8XoEuvCi79W5v0gIW76Gj04ZF
pNSAtGILiB8ybzgvpLobdNSKHJ4+TBOux5HvwedNoAjrF0piL+FlzpMBkXSGbVyAEGqvTZQ62Caw
6CCYfkv/dUslgRrjA5z796MdeICBXihU4MJRLMVnoO5l9LzB33bbujdC+hNUFu4fBwLiSRjs9bNB
klpSKBvugW8qdcD2BbWNXz4v7Xjx0imFYBIqCR/09MC/2jYhN0/8QH1rDL2WBMVYclTU6BcZ89Qb
Kv2vDiQU+9q8QyeB4jDAU2X3vvB3dgSDagBPgY0h9kX+AEHKr/Rh4KYLbTuA5Ebqe7JwnrP0BEC7
hJTwzqSGvR/k78Eg70KGBQwXwd52pm05z4loZrPXj2QoF8Hbs1+kdaNzb5bdJvhXYZjOp3zNiht+
A0fx6SeQJxnPgm39FNq4cG+DIxoUaV4d4LuEXLMPtCc9ySolS/0f3JVSrYN67jLMmefyLF5MuzvU
XlrHYg9n4abVEwdXev7Cs5Y6aVckT4kicUeJgs0g+NI275Zf9fEtjvIsyoBToSczir91xUOiktLv
lMo5R1B8uFvMeo+04EUM/2qg1zrtAQjDGCtl4RNVGDZhbsHf1OIlFkFG2ZAyTYvn76TYfMI4ZzQM
HN2SPWKAfjKnSZ4G4ZsaFYyerKxVjl2D0mJ+ujc3+uczWfNaZH6P3YBiHGJ6MbZseLq2wPVw1ZGW
lnKzz7hcSLARETajIXClW3BUGW/ioMvIuyNL9QEOxHC1sbRWXn1ctO7irhc3V2YeIQ7tPKsAbyBH
Ui2+3/PLAFR+FZ3IvUgpUBK51ZZTCQ6WC/ACqCMmAIhQm3zMNMEW1vunKT22lDRkFw1IUahs7FRo
tmEXqSDklBEO9Vwgwx9l96dVJLfR9/k7sKg1UTwf/2DQRC7syBwyhY2sbNNayqVcqi09tMUgoY9B
yt26UV8J6c3vsMnp+c1yhAZKr5l0M+k7c/zMzGzQ9t/jliXaEwYEt/nwLtWVhjLYJNqS8XoRU+Be
dVt4YSYpOEOYKWQrZ6Ai4OSQtImZxWsm74zr+W/p+nGhAayhzgRFWheno3ky1xwMTD2QNVmEdhq+
KbfTkCAhvDeFpxuwKVtIf5qvZN1gDQD3ZUVYQXu6A5dEwLXn/HA0jBwf3iXY1dk/Qoj8Y2UJwCdF
8LuVQenFF7eqNZavDFdT8NpehZMTCmOUT33niyGIM786xm+7IL9PA9vRI4Eq1JjSxPxv05NB1rXR
Jx0SmbE+RWe5UXMrulnpXSXvPUEfZPBfOP/13L6SKBMCF8sEcLItE6JDu1fnu4wnI0rk589wa8vp
oOxblRknEns02XPOpvLSoO72r285ho9Rk9KSyP+b18Ldg6bHxq4VW9MWI/HIfEXxOm/OsrG4DznR
h/Ey+gQwqUBxsTjkmVuKndTzGtxBli4a4pu4Q9GlKGC4hMXLUb/jl7QK1JikyL9cYjkYNY2DnXoS
XWvD2lz4/pfQf7be7zSm40K4SscHjyUatCRbWZUm8+IpHp+ElrSoEKsE4qyMH43yL7FE2Wl4CuAS
tbQ1WZTJhVFIrK++YUpg1gNevgf5HSr9JcsLsjbkWmAuWhTMJP0F820fdKvTWe3dqVXwjhv/rf/X
FDafe1Ytm84xHyGpmMZvHqhBxxZWW+bh+SG61+np22eMUKHRB59I6JKsPLXh60TUsnhXlR94MTwC
urgDO75QtswfxY1IOEpYH6NkiNQ7EuWpVnabgr6PAtLjvNr9X9IJYDvvngB/BKj6yFesqPiBn/vr
KfcwKLVZUvpE1tmX7uVWTCeHqq8Ihyxdjjb5xQMRK9edBctw6rlqJ6FAes2XiVjrcrwq7Um4CzVz
e1vm4bb+G9yd/2edodG5nz7N7Bo9JeVdViEtv0sl65YRnCYrOESi8VvCfWF98ymd+pO8nw9aMiEt
zKnkLIA3cLS5O55oOtgzTi6lZaO/qcxFLoEez6ujBk9FhYuHCzstwm2KnAHegvPkOlb6Ud0BOrYZ
PPL0UwbBCmF1gLh8oOFsxTfNClr58GfPPmtEY1XSMEa8oVwpzVKcvCeReKJ9DRjJXQUzUIUDugk8
zxfBRdCvUT/1XvuTzWfrctJsWZPe/Q3nz7o/HGVb+i3QJo13ATC6hL4CFewudl88gNu/tVMEsESa
2RP5IA249e4+UnV8p15sPUvKi73WxR5SX8x/A1gUXkFdkoyfv8NoESRTa/uYiD2scY3NstLDpV7A
mohhG8Uy+eOCANdUAMjgeT7RtjOd0AMuY7W8+xA9XUQVw+UkUSr/Vz+agnIBhmdZAu83EtuQI16Q
yqm+9redqLFzRgDnQgGSYew5HMSInYB7SOB8hKabMnnIj4VcRPScbx0miceJrH2bOKCfWxkg2l7l
/GKT0WLizUGwhLQ3oNASEQqiniP92KgISI/mYn6mfSjq7YCKO9zVIfg0T5+D5JcBVwLapB5D+q66
MStqAVvfa4UchEg+O9R+z3ao0f+bxFogLuugjdnLFIXUR3czz0a+z/lJJxzXrjhT9s8bJTUTG7CM
RSmY9VPbfmbk4/NBIOZExcb9DzgHCQB+t/dxInVDX2eVX3RRc+aaTr+y7Yx/TeDNPHenHdRdNLrm
zuLKw5Mx0RN2PNNAlWGWMdFIOx8xJ9Q72y6I1o+atnHivevXXQUMrxqE+JSZ9N9yvmBSIjBEnbIn
O/6pLQXCxgjaIRe6UnY23oGFDmVk+H2SEU81uhqDs68TKzE+QnR1TPlfkXURXQCpSf5mrjyim8B4
dQ4TugIiDdKnUK7q5dpegyzg6nq+2jY5gaNfmbZou6BVCGLHLuBMC8B8AooiPaUsCeQ+bjSDX8Tc
tAovMsKNOeW7fhBiO7TD75LYpO6ZTyRmU6SNiqosS4SIe3uTTRCUaj6OH1tp4M0bAFiTniosyyAl
vvmB/KPyLPQnK6mZ3v74p/3PvDUo7c7e7qxDBTdpUPWOb42EMPLbIIvtGkvafER7Uh3Xp4mjfiQE
fPfsS3fV9E5pNBjBnEEithjF4cHR1nAazU5IN2EXUCRfoDKkV1BoDghUXhW/oqw0j940XGU0sN5u
sTxJe8DNh3sh2OF3S9zGMUzPJvlDgkefSgCyrePiH0aWZjAAXoCGrr6ktzH+9oYGKGlWqXjJef1c
M1YFAV2dZHeIhnsslrRhIgcKJkIqnLodzjpEIrQ2VTwJcwQx/q35QPueHrVxPGoy8dnHLpqLWNYp
OF0C5B7djgoiTdmd2a32urtx3LgRigIqf1+JRd827y2DBKka2ib51ZChwzioI8EtlExyPFemAmru
Vk+RASQWdkNXG7AJvo3XS2hAuJp7EGEPsBKW5JspMjVz/5ebQ6idUUVewYwKTb/zInhXo8AwF+Aj
NeY3Wc8hnGecKWcaVdW51i/n92DP6Hogo1+G9VnkHtOeOcKPTJSggGDm9+DLgUFs8Ttq0F8VjO8O
2H6M9PCeoJ6bCMepJxkpUVX/dQeeYFmuslqn9ck2CEMUPkFbh2Gc51x3FgombHP6+OIiTOgHgNiK
WSO675UOq6TJmxj9FLaMnyr+6bn9Mi59qx5UMEZjDquiThc3zV9oXQIs78vLYDiqGhTC0xV1Rj0M
TpG+V3VFDibf/5M+6dJ2/8QmeGsYyEcZeeR+g4ssg+QJ91TJl8QUr10kh5Dfj5QqaukhIGG4DKMH
F8LtgJM9DE52ZDBwbAIwRksC7RWZ75KDblzC80GFr0QbXU43vSQNXvFq0WR7sngEmNmSvraKQxn2
o/d8Wdolg1vhrTPUsup3+5+bkBaGv8nyXMB6+bJjq1JeMT3vj9afIkWtCyzFM0+2SsgTBKdSVPpO
sOvFC1qKMFCGasyWeqlZwRYK/64nd6ectdMzyJITK9TAHL+8FfYbdy1Yfuz5NrZS0IZyzvExn+AS
7eUuPZ0UEB7JIgqsdnEft4x07AUp3j+sMg5c1YH2DbkdXSt32U4Ag9OujUiFEciaqg0YlBSOB2eM
JKDYAY1hl/Wlf4q1Yro3z0mYHMx2wygJZjZlP5qSkiIAdGgM7xaeYxBup27DuVgcDvhYf+7JL2Mk
wcLIsWVgumLSbX1QBti2Bi7JC+z3GFHmVWPtdD2fUoyh7iFQeWbRFo+80thywDn2lo3KsUMbr28B
beG8qrNKFEvE1SPCiG7m3MBr4/KjkmuWFL5c+DOwQTP4qzSlyLnjJomstI7K/GSZNru6xOdgriOD
eOeouF8KicNpMlX98wUbIrcm7oXzKhgi2hC4g+Lv3j1ECtECZlOy7+ErJ+EUeLTZtko0VOE/ZV9K
gAg7EwHs75IZXUO7cEs9Li3z4SHl9oq0ipCiwK7ciyfmGWyXK0IVW5kMhMZozHZN/WMQKqdPw3Mz
TfyH03KPoF70eipSShi0VrOqk+Cdh5o6GTkPaDWPNIEzbvrZfAMKR9gRZuPCgHj9MAcHD6aoDZ9c
8WKkrGVx4CA7KzfNhhaoif1JLale8A2AWHgbV3mBhmOnDouvzpbGmxjuJUWnfSBB0p0sBsgsnKz1
GfPOL8yDyhS6PuWJGUwUfeQKEpBAO+777zH/XPV+CaiywCbF4N9iLH4y5GM8mBEebkGOWfLQJeHR
I9wJuoZEvkD7knqWnb/npL3eIGgxLW3e5CgyV8fd1CfNlu8HdNKldlieAxsAW2I5Bd001EOc8wE+
T6ZPQ+wMUmLrr7kMgu8dilFI1A1+TGxyGL0SBRT4kdUXiYHUjq+yKqfGVuEFRmcs4SvYPj8ryynd
1NYNhRikL2DU57CgOushfYlNve6ZGDpb0rlgkNCoN3WJUPauZWhL3o8jAB0oFYNUvK62HXd9LMVi
0IFHIR6Rafc2SgLRhVU3F5c47h5wkgwLNmsZxhZax7pP9WTzDbGyCqGkMaxF+eF/cZCvgJwySODB
tHRWLI2lTCkfHK+u7+CaKWB2K2Gfsa/2PmPAY7o3dsi1v3dn0MdvIJA2mqVIYKUP27EUtB37RFHE
72JE8qFGnLLhNWziiSliqbseA4HNDzEvYygfz9lYnz5TNvFuQb+tY4eAEf0IZBQ7OGkmjRvliH5k
WB3CE65ZrKGafyFHrDr+goZQwENZK02uCDFpDns4t2I4GZt8XMMzDft2aeVYKlBnWj/Lx21+1et7
D7MzR2tkXJUq8b+V/HlzuLjjGnECIp0+iM3THThQoaS3JT9e9jctKEZTXAYwQW1fKYb+NXfCfoIB
N+HZCbbJbug5BsvoK/duFCzdo0jxbPFsTsm7dR1QpPc5xxbwQJG5lt0TQvj/swvQPe4ZlAvKMu9y
ze7pv0k69ol4aGmT/2SMCABezLSic8az7yRpHjr65mD1SE/5VMjq0bHmbbosyJl8xytkT5Ou1WEe
niE3tzwe3P7WzXGE4PihHHoLUz5CAPsMxUOsANeGpIY0pp644hFbbgv16avPgoJw9KuozZUus50V
VCvNEGQJRNR0p2NgwRspXvN38/0forSzHvfrsxli1VCvffbaLv6diGFgXWjZFCbCzirIlJVuRF75
EVSzkiO4EtPfOucP0z/9zgjuH99BHMaLMsF4txhWskDru7cTPfM5GDmwsX3xTcHmDWrVujwGq7nB
HzuiWX6oALmIKjGS92I8/QiUsk8WWAZl1FgjDz1DF5TblFFz+m3PvIuOu7hdLvg51iRtNX9jrelf
0kxb97mmLCAqfvv7NoWxk6EPWxMzINCNJgbcwHzlx+vXyFDJsYDLUreWGtblge4xjYYEux3v2aa2
dJhUQtzEVTA55wn3S9tTOPGi59RXtbQF1TXiTnL/IlAAXJ8G7mA56nNmTV9Yyzpc3vujhoUUFFiT
RzeIkhqZRijrurbU5Dwt7C5zQMHYQkpyoY9IoVASgGbbHbxWOiIXP4+laTWSHd3OIYv8ZgTLqux0
JO63ahc//huBrdCfgl9kL8/mjrsREmjBXnOZk4X50lQq7YozGV6UTFFBG91uUFQVK4/t9CSLCHIb
T44fUexjyv2bi0rHJQ43/aZq6Yacxm1O9HujGFP2BKWagHjNK61c3LCAPx5GmaB6n7fQHT81++dL
FS893nFF8dSwE081Jr2BamDu/L9NEbmadRuCtkJqszU9Jr1foRjlVrQLtED3AeYZ5dU63IQEEsjI
0r0eMEsxz5I/XzwpaeEChPksy6281W/ybWzIy92A1m+pAMmjRfDbq2mzGLTsSduYqUU7kki1893N
hwz5KGUrUwSosL8wSDmIezcymMl4Y/6yuM7tMCYbJWGWbBnStaQyKPoZWR8tIkL3rCtT3rZPplum
4B1oi+MZlCDlfEmrg0aAF7ofPPdU95mRQ+2gpETQROwrypvIMH7CD+sTp1mDkkRW6rOJP1Sx+QLZ
oCTcSLXwM1cw0/9r22A1KJebYIGqXoYDwn3yBEBiKR6hXOivZ/Ku0cJs4EtT7HK7yxsbL0OsdzUo
uPe79YdwDl49EEk0Ismlc7VyPxdAXinAFhi6dBbeRU+4M40w4JtK4GIAFwyQxe4Dj0cEpTOIBkIo
c54W6R+iHoSYtUUGYcAMXsibO6l+1uaBURDi8tpZoAg1B/FBZ50fG7b8T2nTgI6sr9ba14CfAeyC
zJiIyIjADkktU3bUarIQ3/cr10Y07qq+zoGsrw1Pi2RuqKYXK3S3VX2p+3+dsOEjG8hkTNJu59iY
Fl5X3pnPXUjHPxB+LVWhiZsmZ7SwjmskOHaRzkjP7sa2Vee+wHNHk2yPM67xvEWm6jA074eEsRnq
BjwMOVTZ5IB//bTbEGdY6YigHBapUh1KvT6Pl737ZmmT2MqwF8rDWGjeAKZ3rQMOrxOUnRK9xCIu
RWKE/wfC+jrykEu5IGtki6rj44zxejkyhbA3tmFtk55Kt6isHyMGLxrA3xGxB8w7SQCzliyZ29jO
7khOCulZgfGdaMD9GIB7jf+LPnvG/NN5TPbM3D07HMpfCAuLmQHDc2akUL0shHjpU26BOp+/wr6O
JMT7fiPKw7o8iIZTC8BWmSUkGTd+uTxCP4UoF3BwebKOhOBLeSV9RWuelUJTXHihCbHxHCrDQE9u
HesaNRxZwSsvJIPN9FgFz8EhvQ1c6zgyxlY204bHDDiNSbUKjB1qstUiGsLnxn4wIXgPT/eOQ4Hb
g/ZyydX6v7L5CqQFCDkvVqh7uQRUFoOodkmFx225onPjzOydmNms4Yn/MEHFap1H/coDG1u/khVC
ix/mspPPed5J/kkkCSeAZKA1Gu6Huv64eBxClL/TBAifvdmBgA34xrbNtEPzfpM3zdh2jsBIZRYO
foN+XoSTrFaV5cmx8gMtv72FBTeBEjstV+ht5skaGpSsMwHaGWKzRuLlZ7eGD1YXfz2EiP6E+vW1
Cikk3Ld2O+IZg83Knawa+uGffsukP9fr33L0LC7yLJe++WzosIEz54wbJjKvu8PJHYneIVdX0eoW
1FZDZOk/yFd9t6Ann/cSwHC/bg0j0zMXfeS2UuUXMspijhDSwE7TBdyRib23ss4E6pK8wRTunoPK
Pv7hZLMN7hN/kleiEtJbnGjkXM8ig9BKpBl9H+5kXUxZ9QgX202TMlcfS+PvoK/8w0ZqyPbfdcag
a6QjBerxs62r5NIx8xm545MHg3XbBS7rkKYBAlIcKZ+5yD1Yo0qiwwtHIaF3qsoZweheyQ0bokJP
o2evSSZlVZY5ssAvn00qHzRpR03VDWirFTYGK+vN6HkMbUXQRvA5kWmjoyahn449xRDvdGwx/ZsI
+JckXJDHPoWcMWCt5u8ngl2OUbbTUFrm+ms5l3jdMicMepdaJo/WDNQk1vKCOSAZwwuRMfxH+2x1
NVy6RmcepkJhBHe1YrE1WsZaLdPmzcxqvD8s2fFTXIUDlWsttojfNQ24r3jIYF/beLm57mS6yokU
brnPtfqGHaIZ7dmGmZ6sk9iROFIemsLKW8UAk0v58ahfXAnqTlzwYL1cCNJBOAMPrs227SltDurd
LbpXvL+P7HtbQ8o41pE8yAYoG2GlBafD++jbxidDt2qy6iJaL4YY1IVceJClzNAhm/RPGDYTqQn9
SXDclFChXhUfjKepfnnA2Oj3B0OD9TBx3MSepqaD7t7T9A1hwwZr3uXfPJJoCeUnDutxkCe3LV4I
0ilIzOrxJbkCXUKrS4Padsc7jm8v3fNjuJJ5MHiqTDs3axwCJT40zyg6jsebWvBxTQ7dKjyIEVuS
Behj/3op2tjABIrGU3qFTYUK+cYlNhVrZilifvKHcinWOxYESIUm52lan2HqGiVnnXyRxMGcJzAG
KiGoot5jNFm/Ql2umjQXd9enozxSg3yZf9CwT+bY1KNuNcSgIiST4nOne7UsfztQtwzqi7ppMCUw
Zrjj2oqWiweMGqnEIRnlbAZrjApWjjNaqvV84FjzTmwwXrX/KKMa7TkDrIuTYM9Np0e4znP5YC8M
uCCveNtreB7Zb6fUhwQLyK1EyYcLB6aqB1UW7d3pJN3JCN9vId5Gee4MY8E1QV/sclNnFcdfduFd
SByQiWS68tuzv+nb5kPGSs1JdXY0AkLapaSGRhfk/a1iziFFTxyV6bNfNatL0gHJTIbXhKQ215mS
OgmUUWS2gkRERw5gajrDryYnUEGQH2vgLsuCCUYcRtEu6sM+FmHXe5yPvNeEIHMFnRtsbW5VIO4D
b0v0ijwCs69w8FQzocBh3vj/gE75AmH5SKXn9KjH/B4lGCkyA1F205LClxWYNWKbIeK5RBnbZP8u
dRdBAQHAHq4o96v0Qtf/zXMg/DOJMU2Hf5yEtuG3LPuTivdc5BT5zNtRtVhrfVdPdx0wd7NmEeDi
LFIoX1G7a6hifu0NUimnq6/v8cqjALGs1ey0GFB4rhCO3RfblguUpDZhLNJwePzmSiYY/YqO6s/3
6ijN6yqg6Xx4Zj/aCttkkDP2LpMdtTGq9DihTMIX5Nx1gzAUnX3aDBF5KrrVWMvgFrqS6caXwKRy
IHSYNOISy2vngCcD7kndA9HykO3sm4uHHBbP9zlPVnlwUei2lUBXgNdW+v88K6tXnLBq8OQRtGad
43DTLOMwJm1gSjKeG923FNAkAQmoQD18HdIgV4V8ynnPWVrgMOYeLYrbGydiJ8iTOisjf0f9FKrp
m8PqXXVQ1NQWDos8sx0PN3eO+op3PzOUK3ZhCOYtdmVpXmSEsUEaJ2HmSmTlIg9BDuBFiiMJJaMg
+pv3g70U7i0HNa41H6n5RmH0+GRToXuLiO0yHA4EAUGI+MWC58vaOSPjZmXo7iwN5zyf9rGacB6z
IZYnEfA2Jlv+7ES8eg/t2oazieNviPTGgZkkl+MIwXFOWAY0LdZjORyuKbQ79dmmvuDZDS0m+64U
YvQ76XV4+gY9ocnHL8opnJm+M931R6cZVAVqcQKWicakm5go5vK/4U93+D1NSufzdhQzPqTtcXD3
gzJwP4lQjHNrCrpGcIk/mF1wgd/mDzOUCcuhLYW2eNmlFCEQELtdOsvgluC+ExZ8jieLUSXGBRi6
hIvIoyR+C3qKsr7yD7AebHGY3ms+I+eyRF+qgW/SenWqKZX3zunNpx1U1Ji9God+xJV90a7mGLuD
1esssEZgjbGkOG5zVT6yE6/mTZmINxUgiXtAvYtzUygahcGJoiywpNq6M8V0B2UAJONTazkgjFR2
cv8617eqnoqDSRglfdLleQl4xFQ0boSLG4Cx+/HRTo8II7G41eRWEkQgQNOxIXKSLdymIe1HQC6Y
ux8vdY6xlflAb/6+2nkxGhcAEeS53822Z1qC4VgxS6Shdn0U1/LrfHMAn2En2EO/ogez7EGudCAo
THdIbvZYKi8vjmYkvsbdWyHdxSeA1YckBhJJOGXfIhAziAtPQUEqwz+yW+ttfcSa4tHoBA9VbAt1
c3I8RCDjjoDPa+be21+hfnZloPOF3e+XCPWr47oaHSzm8zn1ngPcaLoytWw9fJ1CWBWMmoAlFmGh
ds4C85pfharIoyfu0KY7Xr3Q9/lzT3NDwv/VmbPWYqAqZPtS9mJZt2G2hJOyGW64sqW/4Nfh3J5a
XDIgpn7Kwdl9a/lMl6/PPlnww/ARHuWH1W3bd8PRSjqDIY+IMHY5BohtnKlre0dhOb46/7l7L3nB
8mUFZ26qte0bnDIQeZ91GUL1ll1+P7rOnVOyVU+9gSuto8EYPgDZDFNAplyacqJCZI0R40guflZe
vhJ/0TNv90dpz/8I4kY367R+8za4SzIc/Pa8iyqHtLobgSMtOeu2V8P7pKk7/ZYYpKDhsbOg9fbc
VRVAAUGrcNK4ZBBs2859BBZhQaRuJlP5AfDomJbBFW4eHRGOE1Hrm1LX4uIUX4lxO0Cv3epqaN4D
KP8xKh08gvvujW47Yejyb7MUa0pEm0gx/Z+hjqGE8T7ff5rAwoDn2/ewCHxICME2oyeQJAGUOF3z
lmM1ALhCDWWuwl3to8dXndoQXZZzF+qSoSAm2w6eiE+YD1CKcwVs4lF+Z1+c7ZSnO69iocBJot+x
oxpt3R/uzVYl5NK0LOKi211DgYcAPVMV2V2aU1ChIn829rlEc6wmu/BIgtZBEhOM/ebueO8x/GfK
6kuSimFsQEvePRvMip0OgdWMKpOjthB4PeBkb/whPkKqjxdPFc9Sd1quRfCubWA78QrNn5vtXQVL
nxz3rpbLR2pYcvkUAB2/ir6SlU9n3vgBfLKRvE+wIcQjbxFvxS694V3yFHjFboBJee9yYaifaaJP
9QTpRcMdDnHOQ9Ggj5OnlfrAVxJFGaIRo7Nermxw+b8ijSp2jWarb9srlAz02+KdAVQ4u5d5eVyc
x8eHURkSe+AYwcCJBBpkeAeo5PHbxwK52zVope02RO139dZbcCD+RLthDl2aPHrqONkPhox4bMXl
qLQjw4tuBuWyNQV70YaO0XmJPb1TUziFfrwbi6CS26sXJa5cM8wQmdkBCTzJP2+SWENgn9L6agqW
ewVt1VKzVMObGTgamgvZ4zoQl8SQHidnySmqSNGBIEe3tRKAWHl9Yeq0ulF5VvBvn1Ae0v14cT2t
e3Pqcetiv1LVVxR8z5WPGON72iStCcGmGtPQxWcBAPY/XoUHT4znkzmRUjiRZOe3NeS/fANn4OKo
uCfP92zWx17DUe2F5TXOijKJrwghPRYyzOAKM7uHzx3I1G37V4UlWn1xkluone3d8mKCHb0PyEIX
oZrT9nYhqjpK4PWkufj1aw0C69NiQHmwzK/aQdagKBdbpjamJuxYjkkoWPt9NZBf2HdwlgUi2Xy/
v5op1pIFC4jTiOnwI26ZD1Jwrp2CE5s0VweTSq6Uv3AFjpg/jvgK6Y6J93n8rhAZVIoeP5ViK1+q
wPQjvaY3JwAO8hnjJEJJWkQkIt1A5YFq7pozZKNTkOYcOjPVxbDvgp+QbZd5LH3a8Y8ntxMNSQf+
B/rus3ymFsxPTKr/lL2LjExqSPfXBACNFn+zgwWgLqD8yXOYVkGAL5Bsu7qSM9nPFQ/ukbFNuCSD
4MsWHz4Ehc+VBjC3Ae4a3QCTb3d7TWWdMh2rH6tqDBLi4UB2ci6yKhX9vkir61UTN+T9a2gVexMI
T5NLGV77veLHPo2ZQujhiwmsgGgx9SsFxhd6i6cocESxQW0jtnCl6fxWajXSoc+kCdiM6sTu2aHh
aKXp/zQeToRmLamV1VIbS9/Xnh/6GW+4RlBqFO0mvaTpvwExo7ypemHOPtks4Z0UWX+XlBkBiWvR
zfpamvA8oNkUyQ35CwIsovcuenR0Eq1OOFtvsxmOiqmy0HfZjZtg3Sg5ZgiRfIYf1qKxy/qF8zz3
o54QadC/y0cLsiBN7vsDReB/f3NoMHyWrGspw0mIdj7pq0ov5HXKMu9q9pnVto2PYb09QcuvQ28l
wUsK1CJ39qNgtcFeEWq1btGyNL+6iPIki9HZEOTLjzxumtmwX6FKBLCluZPVclZpbw3acdGUYXX7
1Zha7qBBHwORi4JyhQbGNQdAXoK7JuIOhsJ/3RW/JB74mTlsmEYf5IsZnLkjM6FUIsihSLiuTgGR
t5Y2i1z850ZLOeWdj/ZWrcmTJlKiNHnkckWTK62HnorPkwI7mT30jNWNna4ebQ4WvkaVRMl0ifeX
TNd/njem9cP6O3eJ2uSbjhCM72zEnF+xxFvW3HtPR5OIA0vy4sNDO4PJVnrJarM0CHRJNhMq7laI
4diBeePSRvlKcoddP8Gptu62POWHBgTIo5K3qwrQJ6JofF0Qab+ZSclFJ43ioPq4lqGY3Ot54MmM
JqOmnelUhCoI7WC0B1keVBN+kTBGJs5Ebtc240yOXU2Osv19f+MYUj5tYj2m49kh/s5+s9/66IuW
PpwU/e0ns9JgLVcKn6NafHncOAxIQ3HSfm+92Eu2HizLEHMZmhTd5wrjSS5EV4xzqB7/GHP/TxI0
7NlvxxO3SeLhmDSk+iitEsku4ASidxyhW4uJE005q84vSqDLI28k+WvTpTwkZ+tq3ke1VRACMonX
dj3t1UkBskLE52P7QgNWEBGgoCL0c05DCtZFr/6G1QSNOSs6HwsqFMOwbwQSGr+ksZO3xMh1Tg72
gofjJrjRNaclZs+UUPJL939MctKfyOrcq9tYqPzBOgONOnJ7YDbjz3Mgibrpc29X42BQrHf8zs5v
hxMWtTLwBv3bwyXE3jbJqn9aD5jFvU81o4uIJJMS9ABvWXByK6Nyav6C1c0r90Y0LBjpbFZmoCe5
u6OHgDzEdcVUq7QXH0oXV9TISbq8Hj0dbzel5Psez0Rk+ptdnb8Ufb+08XBg7cVfCkAcZtrq9q/J
sDxWGmebZ7MMNvOmdBhwiR8Ko8nJrh70JCWqRDgPgnc9PxIt3ACNASJuMFMtxpl2eBkgpOOw9zTF
soR4DJZyAw4djIYUjp0vP1RXNrQAtyVoM1ZoPRkcJZAqKi+iF8pQmk6T7FgXn8q75VvDRHeN5TLY
LE7D/Iqrg9HBgM6Bb8wIpUex6HOhH3v62qbfgc4wqbsIXfCRGbQEgdXEvSLK09CnB+eo0kf1zhAj
ZAU1fUIBNtomOAzZ8NNWouqkdmAMMNxfzHJ/XLqfWtVfeg1TqrP8WyGtopH8VWxCkZ5FvdjzO6ki
6nKX6XAx+JnTxHzQIIHFFOYparNpRi/Oz3sVOmZHeE04TMZUDT1wBnDtruBAC8gpIiOPQJTKqW79
l4J1h+egB5USHkXO7M4aTYWZwEohYwGHGyi3aVBp+wNyZ+PstcpOS4bjc0VWTgTmNwRASILVscl+
pVx9s6Zzx002WvKdn/u0JyLEeJKqUyN+Tcti9iqkuQeBUJs7KC4stu0ZwmblLVL7qiuP3oM9tQjv
PEm2z19dsrjmSM2hJMs7SmBDjBcu1JH/0d8YNXt0Wj2jK8JrQVVP9MvWKYypzkZLTcj19v5/1x5d
qxZx8lJoUIANScQgMtluwP92ehquwBnBrGY0UlfIOV93FsHDKrd8rFaTFObRRbwoy88D3yDFJ05i
NaSyNW9B73eteYEeQSxAUwMAcxPRDkXIOKSZhRkQmcLCIwmPzZ1waftWfXpnGcrjncQyeEbsm3ZT
VdBqJeg4GUtuG3NHoxZ0I91Rlzi2C8kC2F27hgjI86OJwzxq65bUigTMg8ulStBDO6cWQiO5jdRa
wxxPfGiCr3GncRa1pcMiW0mdo1YrKOLyIMdiI+wGPPqxegWgvzbgDjPkk8bTSH0b9Kv6cyXGqeKR
V93UU37ZDP8zkx0ur6ZmMlU5cxAHuT+dR1rd57mAE1BT9nfZ5GBwCGiDIboHsoUq46Zzu45cZ9ck
sGDzMawBQl4LUHd2JjMrBce8UxNZoV44ksTJrKStmp4B7ZmrkAhnOf2V3SHQNQ61ZDWs59aQn00O
ZP7hXCPvlwRcluE05VwHZj3e/EpjgtRYnUreUYRJU2IV+ZarVe8nuvcxSFKLu2fzMoZhY9a5lk5u
GGSfd7ngNNfomdd6029rj24MDRLNzPcEUnyxqJPUaKCZR6/YM7ZGhfE7SKZ3acJxFgiF0t/iPpBU
3e7T2G0sJAOdp42Qve2nHTl7OHh8aUSsnwXpPy53GNyob10qfvkrSE12zuMQl3BW6IB6XOrFtv8O
erxojUMv9rX/NdSfNY6wpBXTQOcB7ubcTWierI+/HdiCMYA9XgMNBjL0s89F+C2iGiZf9aTsmmOV
+YbnMPbLYM9kERbMNHE+PZlhlWGDOr/sU0zXN44UtFdiy14QgJM3yjVqOPoNlHNdh4Dr0X76lLmx
OB94pZdGnq0mK/bIV5Q6YwRn3Zugt8m0X4BnF0Kke5JgLyEjl29EMFyih46as1RrTYndEl6PIJnv
ZmEhmFshdkbdnq4W1UzdOfUmHp0jOk2TBIKIAI3H9J8vMPp2zF/61IhefriZsCt2KgG6FY0/ecTJ
uRTQnc0s4qVQMcCymUAnt3PILRYlTSNgHNAFjN/z6f1FlrZePZ0/4Cc9j+rqOkKegarFM7C0Sy8d
l8EEcNA+Sp1pCa2aDuPLT37CYAAMh//l/zrJ2NJ/xMNu2WJ4ypbrC655RpQwJhmJav/MeRgmlokm
gLd749L3yDJYiCErEsQDIVy/dPNzQGNaaY3JcjTDUWrdxbqzP6InAs+KOoVe3YfyMswWrNEZj47K
A+Pfk+3lar4mxrQUKtKXcFdnjdvkHoRcnhsjAxiS/lxbnSOd6erqn8m3JTLNjUxwAXbIA0QJtWD0
ZtzMe2+BkUyyr3iqsVM+jfbgXqeSfLNoaZsYhZKzFjNJhiALiGkrtYd1Uf8K1UlKEpRY6XD/0TFJ
2MNczisi3mpn8gmpOG664ChkeV8M11R8F5ap7anLGnOsiz2snNIKSXYLYGylPaSXqCvoMavd1anr
G+JZ84Nlt5V7LnHl3XIcv/rznbFtHGXvVC8uqnCiBu/neFU3RYcKKbCI3xi6sFjy+vtHeoD14edQ
0oB9YT/raAbIBbRbl/3HR3sYCt81AKPX3SRC1bZ1H3qWQtCJSCaOF91yfM+2ndPFIZeZ4/P/SNnp
O9hSsWsIgxTZjkUz4/+fATII6dAnPliXSHIhZ2vyHwq35AOJe9UvW8MdzQ4P2NjcdAiXbj39T576
6+FPo9beplS+t1CvtfpeoZS80x1g5Q2edOACGlSeTOCWfkG6FCKDHxgkahnH8Kswl4qv4DLc94oJ
Q0JWPnPUQCyOl1ET2agn+aJhxzkmeQhJYZZP1TuYjSlQG9x0eokXXKKRrBpVLqOAPstxSUbisjYS
gye0Y4pC+hv7PgV4hdpY9s4rpOYVnOxW7TAYPXvBFAgy5rPPS6/xgqExkUQ7/H0a0xDpiq+ePjBy
yiYYgKk63wS2GkHXiXbWUIgQmkBg+qZMTC9sT1T8G338sbL9sRj1N+HQ0Oktt934whg4l+SCdxIb
YnakFast/UsiN07gTI4FeoU0f5sbCdKlqx9GLtz8pcJ+fHmQ87fCIOMLlU/HaN7pMkeu8XA9GYc/
YNgBHkZSFSJ9fXviYUcKzPIJF3wBJ42K/ksS1F4K/qwvk1P1n/buCw9ekm1uPbk8lH2xyjebpB82
xdKJo2Zpw5J97CqgXuYNtNhlT1j43LWmKj4AW9x2FUiPpUyMsQztCJXMKrOq2Lh9UboIJGJerHn+
aq+tv08iOHZmUDkJnZm1lI6iWZNx+6TgCnBF1WTBQJib692gPBQw9UzetRYHl92ECpRO2DT6ttjK
kwzg/DMut/2yM2yBB398aCJE+9+y+CvZh1KK90kHQovwvG+zeUkliu/louGlsmPgwHgYwQxyK92D
v1KBg8STUpnvbkoCHrq8EijZC0FDS6KDNme2r0Fsz68BeCuowlfrt5W/JbvcXC+ojssPqggUOUt0
3EDskWMsf3+jFWlBwhiQ7lCku7YebWIVAxC/XNBPrlyy6D8SES/fS1U77SY6YoFuhqohqNlBjF+Z
U78kyPT4t9XelWnZUct4yPo/KXqwnfRJPcIqBCPaLUYzCHs4jQ+/2kqY8OQ9OI9tXe0qrfOZeqNI
IbRDYT0Z83HJK0KNPQCXO82JofYaNd6eQnVMSLOLl/merqTVfwchuXqKOBzE2uBazFpPzqjYSXLB
kBkIw4f8bby5DY6VQu6Bpv8YSmCCVXEw+91pbfntmeepbVy+e7aFQHAARU410JKlQP4+1ZS0qjZ8
JpNawRpyIbgTkE+87JwVHIH87sZ58+sqwQcdD/S1bnxmSLLM32m5lJnWw19KC2qJjJiKTGzmMn6A
ilEjnpxRfVvsYkko4OLUzirdo/aDdhuTfD7VTrPpZs73+6RHTztyt9SEc0+o5/jRd9LYP8ZUOQzo
9cdzEgpDXI4p6TvXsxxB8GMxiU9uWI1BTe5CVimmt7thudQEHSeYcyCCCLKHIgk87OV6vTMGg1U9
lZR/+GcCuml+CZTVoM8ldTss28uBxPLJNPixT1yEVUKpqUED4kvyEMWCIiSXGdQuM1i86lkrqVfV
Vhvs87O7n9qhsOLl/LN1On/stL17LokLaPcxTLNKOqcfmTfaF8iap1X9/hyg4T/PLH06BJIux77S
RUKEdMwIwmsRaVXv970skfaV72U5TxeXrSpvRv6RTMgyFkNIFZ89kohf5GSsl2zJ5cSFNQ/GEk8O
zf9cC1/KmkKe9O/WcCSzCBuZFbai4w4BPmehuqLLtuHusfnW973e+d1aREOqC1cWwNcXppcBTh7g
DsPT+GO8eyFclsG/SOfM7FsOugxRBYPMGZuWa8Iu92U1SqqGwVMagqdNbtKLp4uC3omOM/lsI+Pt
Yh6SOGOKowC2uZ1QmiRABpIRf9g4F9yF/Vwe41TyZJXqhr4ZkvVbog+wSTIXJu272B0i6kBlVC6F
bEoJ8GfZpxetWbaeg630zfxWfhC8W+lc4bf+ZAL43xepQLzLbMRevLH5XeEwit5ZbiLaRH6X0MLu
B1D3aIIc3ZBK9HiKBc67w4ev9xSae2/vlNO3MLf/w+SEBKhzz3uvroJ5sve/Gh3pMEnDCS5CQeXP
azG5fW8oPATE10glSNyic4MG0iuk1dZe3EeZf1QukALOK/YFgmdon/pf6bTw+BxA2iQrlF7q+MYU
tx/Vx6jvizqH1Fv7CWDVeEGvUt45ZfTMT7W80BoFl824qPrQOZFf9/WdfrdCFuR0SZSiIF8vUFKx
cbi7vx93u7b15pJZtL497o0wEh9nv/RIurLx6KZFYloKkCau1Q1UqZMBSNYmLRFNMjQqurd0nmZJ
iyXoA1krBKaZnh01eLIxWWlzlarxWJdMkt86qdiRt8DhdooJ4ppIEeVfv6HqrW/aKiNedV/s9Q9W
VxAa1PjjsJ43sg+Svjsk+2eTvcpZ5JNQkE5OjfcHDnFVB0ILt6LIvJli71LijDSqjNgY/JXv8+0p
ZFuPi9ycXf1iSSLxaDSXGxn4IQknobrlJ4enDhQ7G8UOJttWELh64zlu8CR4zxtn7UUf31cUXSaC
v5tZxJeUm1f9eKvczCbaaii4eq9otxKDyXgOjsQ6UiPx93jl+ixnriNGVDHXjHzxlD2KwrnAYLlC
39Gg07tGBm/9tSOumGkoRf52AFoyDoKNiNhtPBzShLamoCX3dA8yU7K42g8ZuzEXE0pEl5xOnROd
o6hVJLEZb91Qx2icrg/Wrk41qPXg+DNGRlApeVRI8J0SHl1vvOJVtgE/dbClPh7PNK6qRdv3tN1O
4LaiBGI61rKvkFKtYeq3M5AUf6WHk8KedMw19+NzrX6c417tchogAbawHGX7y6pM36huo5/pQhsc
dhl4XnKmz1t2q7n230NYAkuqkJFSedNkcQdMbwN5SlBegsKRKJ6huF7tYhM9JDx7UZupdg63JS7K
KcqEINnSUHzQx5/r9SApxRTb8sOu6vZe7NygtgcAemL95ElVBNAF1A0v+MjLYolvYkq2Li6zugQm
7DLc2SsjJ0QO6Mtlh3/T2BLuet7i3Cw5pbc+qhsVYB2fs56qkYt2SsktgH3QKgwSxD8Y83ewtey4
epXg25aFFmdgndra2cxXLvstiZJf1ZA3NHQ+Np7jn4VwaJUyGe6GVYOfcAjO8Et2GvnUlqb+7kHs
KjFzKhuFHyDVPARdNtyNZK2hf27WCsp/815Ot3/fufs78m1MFAm4KakfBtjU1uOSZ8HPNupjXKTB
It9bWzlsNTZTNV/t+Zp6C6bFaqmFK+0AwHupOF0TSHBL8cKZ4VDFEjkCKcsHCZfSrFIgq+RSvzAE
7UmOk6NY+EPy6EtdXKPHS3FvintpUd00LYY4H7LE9/8gCjKj/AGG208q6uSKc7ptxHrDLdeoT+Cs
w2NrQpo6Jw5MUeOywXKCT2YxOro6aRQr/7gMYUrGNCU+s0pYXlBbRG/XSlVNDMA5berjCNVPHdWF
5dzVMpNTn6EDw6DnGydHSi0LHKuCZGg+6qTPgxwIdCr/q49gaISvI1jugLjBTs+ETMwvtUfHJkJQ
IESoHLatSM9tSqK7OZ2UMj1OBbrvU4U8QONwyIU4Ur5ARDTe+kjmquykAUaqndE5dqoLvvdPXQfZ
ug68KtMdtrkaJYT4tq6QJWMo+MR7RKrISsz13+KOqdg+sAI+Ti/Ie9QSI904E/EyvEN82ok8ZRQ5
hT/umLeJM6/hiWGUPoZuJ9460HPEgRcQWqML5DLlkaB3bbSyWszgHSkjybI1dJjE65v170M5IcWt
QXhd9pxFZtDAX6852CbBLVkX0iW63pSnpGwEhqa2BDomBTB2nIqpU6jrNmp1PgOIE1WURRnf/0ik
+VNeeCTqHczM1NzpwYEHe2zHJPrqsdV5EUpmN6rvICnS2xQeW3M/Jn/cFBvjxfj84KncFjuFXda2
AHAdotolbhqXkysrVQwWe0UkiOB7fB9RKb/YoTJxheaJe3rr1wLUiAO3E14RdBqpm/yq9lSpfH+2
ivRrroRXUmqJ5NgIsrLFZ/e1ElB6kpvSrpS5au9CvVF88iVKEHFtv9g0FFiDJnlrj8vYmvTiveqh
NB/+5D5YIqDKs3uCwlWfDfxu5pmCA2Xg0uaFdF+z2MJK4r4uRCSsvv6zmPBzJVTAr9+XpnamcXi8
24AC+/udONS3+WP6AjrRF18q9f+65DuUjRtD4WJkEvxwCs3/u33VGsTDRuGPn8g1VyZQGdc7fZby
TuMm/HaJYzsuXIPE43r7byi0HZg4D9nnocySIjP4UCeF9D9/I5LBBSriRSnaCk3mmSpil8rgHTAH
ZA9etWDnWgaVvFLp1nB2UapaKEat7ziGTR3l+QC0cXGPH6fZTayuOr43eWKAXnCEluwu7KOzruXT
zgOaN77Gbjb4q/LN5LlaImWHjTPw9vPs9l8DgL7Y/H+FmwB3E1+cb+yv0vppp8UWVOsM8VlbdQtz
VFCA4K7xbzOMhbPw+bIbWrhcEDfCdp2HjTMvVjCAMYtFZ1FIH9YsuPDx+c21zOngk0PTJbF39iZy
C83+rZoMcsaY7PHp3tHBt0/RIcz+kqcRQZ6P0pzM2bvmPAnQF6Y4XF/xlznL1sqCrwRKZaCJg+eA
spWOKe7yv1DlYYaWzAqDSTay+dsCykKAFlgBGTi1oi+6aV/MCzWZWWjaxjPIYHG/s9PnwBvARShS
cqou+8wxP4Sjj44jbZp1eIV/tkZcX6Te2+Y3bl+P8F/VnaPCQaFE1ZLBc0ZIkq5EWU4sE+TOpXZY
6Q6msI0J2MP9iKVbW1ncxOH9M+wblellfeR4bBdbpxQHlZbH4y/143gJBn0Em5WRBugibgL99EA/
l38P/TtgIy5tm+fetp4DOiochqHA0qIRTIyofC9w9pG0WuT+pwB+FZPqUPaYUO12o4Y539OZmLnK
xQskiosAZj6ZiZjMABmzC3RSl2/IQCXPJhZid3b8P4OxbI1XIImxNVY1bdf3ivJM0eyIPDm1Mv8t
1plGhbjqtA1HXLEElHdHMbWKU7SxbDjRMiougERscdl2z8Y+quIs108MQ4ot4YF4q4Wffr5ma550
he3AI7Vc8OMj9ZG/73t2WSy8OS31XMtdR2b2qwOAdMirQL1nujdmyodWdCp2tsUgvdaV4eIwW0dm
FwfRiUZENHbg4uwwb7/H7axVES7qUtHdoT8kIO1IwqnL6fdp7bHUkSsk2HPRHzRGnjJLy/QwpFHW
BmsvHf+y/Qpy/t/kJKomibJzSs73itxZo3G6S4rIcsgjhH9jb7Sz3iicDwabeXccM8rU97ZEe5tg
vZ3F0kNAYRXE9NMrtrCMYKvNtwHkjNECQZlIjxfY8BMYSN6fv464Y7c4wl0H+TaESVxY3UEQweS0
gxDCr9Uu8sI7wDya0MCEwL4kS+HaWtiN4G/fsjHsYVS/tJcCCWuzsucy9KSFm+RVQcvDY7R6BG7e
DSCTewu7NlwOmjjXOOtK0k/D6dY1KFg8X0ekwgz0oBEUJH5MxHbGIOIQif1ekzFWhF2zOUf6btDf
PqUTHOjwUnW+CGLP+1+GeLYc8x+6xYhaa7wnK7mNCv9Om8y0pHP4tODKwdapcIhxnVOyl4RNEUOa
2CcU6/aanFKZYjQ3hKvmNfivOmGpWMao2KUl+T/NM6BCGtynuWIXc+TH2JrLIM84E/Fdx6D2lCWA
jCGvI9rQH+gyiUwVbP4jWid0YUYy1QrTv8tj0ZxeGaVwU+LP0bcELo/bm8Jd8bvi64DFueusq4fQ
gWgr8HhkFVrKLeld7/Ay3Snvu+CnzCHsPmNOHe9ThlNF6hbPXiaAVNPwRAiDPIAb4m0runGL5ze+
wRS4tiIsN/sQBNelm3iHn9CL9mbLYvrfJaJjrE98xilQAgm5bMCKK19Zc2dSdIluxzxIrPWRChFf
X5LifGkfpJLv3VBnO/S90iQ=
`pragma protect end_protected
