// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:35:32 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
LcwN1sNLgnljEEd+3UK4KOtx0WWV206uvWPWiIjMOL9aWgMzdBPgkirdHyBl15H0
UxQCH/LF+zCRCqFWhtHjBgWItiLJRPxeT3zICMvqh4AsEnGYvaObEL9zrWilwZOQ
gVzykZcEUkq7XFyzEJ9lq64FYNK/QhczTWqTWVrFWhQ=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 4512)
I1Am2mKfE+1yp520DUtz67aFUkybYP5GiAlN0EuRjp6xe/23S2mdtBBYrRprPpeh
5mLMmxe2PkPFNu7j0wQiXaQ3ETwL84KW2hgc78i9Y95Bj+Vi6++AIl93qCzCMJSR
G6qike+l3//6dVwmQS0LW6DYlUhv8WQ1AOOoeDSgDNbKHa9ogCOnWjK06Q62mhdw
f9uzAWlVtlYezOcxNlPmaDh/PP4CBY4JpHpL5PkD629QaIgn7Q1fWcJrRGt9d8wE
qzyqZcNgB9FRNOmFbNFSFn05SnjcnThu52G1zi8sjIM1ucJgKe0R0P5Bi4HGDMgf
jNKHoSey5fgl9eC8HIPBEY03pl12nRP4JjEvzlSKqniDf54W9nJdC36fr0L3LGri
qKRJVvG/LnnzvUhDhOI+T/3h26oK2WCa3nNCyi++bS2mHO7Ub0+nbDkmCwHdgrmR
z9H0ayD/cmzO7BETAgJDjXRKhvjHPeO4k95/bQXMz8CqodVXRIgT9K7zJm9NTqze
0m3HRM0Z5Bqfi+TICfuHmWrQLjbV6fBRBuoBoW6PX8pBj9ddwkRUecZxOGkLOAU2
LS/wJBUv0mgeqBHBuEkbwImNP0V+mgZt6XYbXVvHymezBWyeYcZZobFxTD+s/hRQ
ikMRJpzrAld61rZevOrlGboH0ZE8+qSkOZeqXKZllP8vKF/j1PWtx61Qf8my/x4l
zY/BO785QahCYTJh67V0HdSThrW22KF58xXQWGqVZMNh8xl5SKSZ5aIy4vM9IqsO
/3N10GlzQCcBS0z5ZNXHBuQJfmYAMPlmHobVATSlgIgiGFnCHLy2lizXkB8R4Cru
ivTKwOlSr/6UtmyZGnwGTfxDs1jsEkbrdt3irf3wLKxvCg/7/u888IpfTEx9eB8h
ADUXMtCZcKnhpXdLxk6L2bqW8mgfrfk53sfdnAAgqOYpOh523p2KPtOhgZNbobyg
nH1l0f5MmJi2ynQ/uPiRx8J8bZtGLhPuVIc+rkf7o9KaxXJOKG+zA3DSpo8Bdr2G
DGhM4W+dQkpEiQjDTq1hfQyNeNqeYW36sMINYeA5u0ZY3NsyaQ7PoyQQVVxoKikX
UyTl06Zjn29Dqk4ZuevcLO+dYUn+nQOZkZ72n9PaA1gco6gcFY/2gmM/pPO+MIZg
qJiKInoPh4iVfOaY2Oox5dqEycAuY/uOkhkfzBxhGDb7khm3CeFSjt3KFomIff14
YieC4ABQ09dDoh/atDyJL15xMy7P8+1jdQViuJjQ6Ww+XRTW77NQ2q2L59GAw5cP
uS+Sb4zVCHlFGbXtHvfxoBwWbtHjUu2zuB/uyAQLbiCEU6MvyTyCnDUrCoXFxua7
PkGNDNypXMGvbdu8WuD7Pug8NEF0hlER+lQSx9cCkOE9hoyqy00xg4ALMKtIwYBI
aPaHFGrdBXU/O2cIaN2wI4hJSyQmUnGC1FvkBtzCTEKovU4eI3no8yIkAiPzeGKG
TSfjNtZJLD8fpcvUsE4zV3u7JEVi/TIcE+AyxrgIDuV2+CK7BVfyu2O3VRW0iEdB
1G3GvgJNRv7KxFaaE1cvNOp5Ti1Xq6NKm2kCMwgPtO5jzIm4FvoBPh0sIK7e/a6D
K6JISyp8/jYWQuoA3I2APE/AGytgLl9wHNbM5eUo0r60fpAv2JnoK5Bt7E+Lx3n/
uzDbZxTh5r8kRg282LZJcbeSbkm7qcg0fy87XNPwYMINx1MVxS7PnkM7mQm2JXUA
5DIuxT16d5HiUQOrgy4Tp0D294OBdqUlYQ+FTjZ9ocUh+C/JsrtvXzumERE8odGt
8m31q3sNpZFsSHezCUFygUOR5WfDSFMtWJDH4C+dPBP4o9HzsYjRCAZB/r1w8UH+
5QsC2ttbh9oAjFm+acI9e4hA7UO83bbDvzpYz3YHqFhh8sUNoC5DVMcTbOLsNOMh
FdfBF7xbr6ZA4iyk/iP4Py6KXu++pkPz5c6qNzHgSPCAX+22aalfwIqqHz3RVrJY
wpn5bw5IrsTkHYFp+YhgrUiuraghnDyqf67fHcxmWseXdF9PRa2bWlZ0EiXaGkml
ZgsGCpUHxMHnIiCH9ypwjKc0QPIT3SL0FxoMJRFVjeS2w3Xkrco+8t7CjuNYAWYA
hxGkOzJc5CswRc+nLg6Ta6bzjB5avv9dm9KuwVfJTZhFH5OVcYCikDVstauDQ0nA
6NVdEyXGARRh5SY+IUeUjERJliRN0KnGZkoQo5ih/govP0V1ma9h0nYOroVMm5Lp
ZXBKA93DJhwJDYZVPazE+O8k/dtH8AfaXvE+vQx71bOgyx2nUbwqIVjojutg5FN6
Fx/Q7aS6DlDZ+GoflefRtn2ypZa4HYnBsHm1EVsc7QLERoc8lbIZy5sgTRLDNhxP
+on1glmcZBM5XBXgHpZmc0AjqP8guuIl9N0eS53CwwPoJR+z1wSF9YygO//Rl3Hz
3xS/GgGOuO+STv4DzDR/6yRlX6VOiGzEQ8apkATIL/RGXsctmJSqa6GQp2OxqeAt
3GhlGOjdirSkFIdHmAMf5ByAnn9P0Q9Km1yhK/3+D4r5OltD94thRsw61pvOfRIl
zaaYSUMKJ5ZorIVM40CdqR3iXVO8+HoqWcJBoknGYr5C7w9+6YCMgI0bSeBDpegq
1RiXAW7TszygGxrtOETeTR4hhLGeoA5ZObONrA7Fxyl6i7JcPChLL7Vw6lP1qJnG
He8BhxH8wraQE48ZlzqgAf8Z5JnGEQzBfeRqzm/4ffZtpky2FW0KfXQTNflL/+Y8
dO/OrLAVt5nYnh4hhmkuECw0+8QB02XGeSezcqfDadgqbY6oyi62zNUEGQAJYNHU
o51MaoTIDQ0daTVEzz7wUCawQDBtwVaAApfzbtJ3iLaMaUT8+ni02pp7feUbme9E
+tpPeLNK1o9SW7Vs7p+VlEEKqrvTdGmdlrGsvbTA/9NGcBVNz7rYcsrJgHCnXTYn
KLl64EevSHdua3xsKfSVK30jCav/dvRQrlnkQ3dWixLrxZ7+Fo0eQfRzvNKETcTf
ITo5GrF8BhFx3wn0+VaiS7XQbdUZqr0hPsIH+07+j+jLgdU3Oa10ID+s/dWxWYpN
Q6k6s5eIH6AROhUksA5DxjySSV6YoxUjG5VyVAEzmyw6ervb8C5DEuPe9EflnTo3
FUIlolfDMymylSjFUo+TEkpwT4pB/5LD3R/MashxjsvFNsYZW9wFUddUsrIvF6st
Az9qE06WvNT7VKju/uGRs0X7UT9Ml9ezzjku9O+MiQETpBY+ov5ehuUV3hjOlAm/
tgckTJtgHDO5qfRLEc3eXboKBAZcW7SEX2X7hNfef++7UpdOZOVPctd+h862F4yK
5dCZ1DkXX+wsrKMXSgAxGGXT2mcweZI5SZEKMMCYsN5YhfHhWnAUYwjKRSpvPrkL
01udiVtJVqkAx1L43vXj8bY050Xf0FNshHEEhRVTBG0cXVxaCuV0qUuVis01eR3U
0fIf3OJ/vvATOOtsS4Z9HibqgPkOva2jZxw327iM9tzzzoO9OJvb7gXP5o6/gY+9
oLX+B6QkcI5lstmnedfVlD5ynHzGsApwePMgHyO7LWgr+XdrRd/0D556+LEQxaAW
CVjk2j+5qL2fKnEyvdQcmxwXScYjZUvEEPPQN4F+hAJngOglEXQJ/bqC7jiq0/Kk
HXoI3jEN8FxxFxV77e1zcrnmiSg8cOXJmIhbSEiuZ3F0ATa/O7KTOx34FWb5gpot
y9KqggPNWUOgD9sjoLyw/uYOuKU8KUiJ5xvu8P0SodzTTdyJmMmWMblvsYrUuVuA
8XtlNKMxQh+zDQsUABMiJ0Q7bVp4Id6YDGFGvf2B3VEFp1FmAP6aGF6phL3EDHbZ
Mw20kDji3Pep1q2L4Oe/MHYPDrY4wqy6Gu/l11zoBYzEHHxUk2rn+1wUa/HHU2uD
1wmy4p1TWdWwlkQCHRVuEPmwFCvXEZNNad3HzHso06OWwDACW9MWkQDh24ODf4tn
KmtFjeWDFiTqxYNCJcphLZ8aHuc8PO9KRMs1g6G1U8il1NM0+ooOsYWI69GE55AW
0GsTX36+m0deGrCEMBm6ncOqlSIAQg/piiPhLIxl8QbRz0e5/g7jq7lD7d1Gnd3J
8kUir5zmsg6bIgU+r9NVaaJiitoVRb2+RYVWihyOWoFYsxKMWSAXcnBr7ROFoYXh
nVUwjZroQuIdEfRCNzHueNejYDkc+gIQtvZ8C6AM+CiQ7wY1U2w0D7YgGL4yXLMI
i+cGqjstov4oVdnY3OBTxRM1jxws2gNGLZEYWT6wXHL3oRbZ3F9GXo1AlSAmpmEC
/dm7uSXsEzi8Pwp70DxI3J5dQ7fZHj/fBt3sjpXwdjGabMJBnWJqX/ZpvG8zjxOv
CTmC1tONUDTH1OYGvBh2OFSfazYZh5cdHRa0Z6kwv3MKga1pbYCLWZeH6HfAvQAA
WIOj5FUkpkgxnCD1YW6XNaJFgq+afxJvP1qS4IOkJtNF5Wk44mbhCyI9R+18dLZ6
f3KMtxNlvCzkdCnF7XCyydzvSb8g747hj1ONy7a+fY9HkIA4rvmLhoc1XPDsRsy9
oWTI5vVem8V0bFyUbJfoaEA9t1lSs0PxHvhR2L0TdShaUDEzFxuYAuZabXZeo/72
tsrD/CkBQj1yffCORAtWqE5ikfFdoKzfL4I4ANyHB88GVsR2z7AFpn9pmimyJD+P
f0je1old1tYtZnGvMxqCFTR3JOX4VmAttrflhF4UbGuTrlrzeeZaRczILG+2Mvx1
lOtf09qzpoLk3LJgjQZ9+c7Iyqfkuc/opdGoyzKMhBp9ileyQHifH8S6W7w/vKEA
cnMrkDRmztchyWg0fQp1GOVB88uPBOinVBZx5Zb2QS0PxiIHOJnmNuQq1K9MFsT6
YsyR5bDvquoQMD8Y62TRsUaIPK4jinW+Qwz4zn9W+p5VWfzcD0jw6ToTfNR+R2E0
/I35CG1eoTB/TeDXFnH2SdBi3sCU1z4CsaGUELiyoNEfnOVV+frgrg5DmdxLfsIp
mFQMyunBLWcrzvN3b+g9Ow8bya8jCHpXiyVzQ8bA8mXLVXMmj9wj3ZyY8rRbz0Wa
MyEm1BQfGz3/G8m1PI/b3qOE1oenXNYFohR3kpO41IP/54Tq80qUBRITbLr7MoKv
+FJRBftXZ0Y94iuT1waWWXLoQX3/FN/SCpbq+Jh27/+MF8ehFW6LtuH/iD4cfsK5
937AvhusYd0qblTlFDLyUeF9b90RCRDnX5/+DhYQEew5aa9w1WSXxGC4/4Dgk1PW
V8DtAf79+iz97fISTO3hBUcSynaZ08BynVHqAWbMiaxIklAlOVbyFIZ78lF9AYn2
pJGLl/+rsN7c0+sT3RkZIj3eN8esZgSu6EDuNEMjD06iVGS8h4hqwaCZb3gUi947
yVxdQxJK+6znWFGtMLstR4yhESKEjwhIquyneC6y8FawISVBoLYzPJPGnLy0l7r9
w/wpiBbpqMuD+HmJJx9glRhlW+MJ+kRdiiPPYbOoW3YQqTYlwMCSVCYPigdpnauv
Oa3zJJ40n8LlO/QnKft2etGrY9QY7kbN2hPiIE4dX9bSF6YaD96hECTPUlXlQNRu
K07iRhBlB2v1jXLkX+zvG+dIVC4LUWzF45Q3wD8G3AtAeux/oRBugsvnBtkJk9t3
aJYcYVymvCEHBXvEv5Tr7vMlIB2Ykzn4SOX4oH0w8M/5DDfesvcseEV8j2DWu0iR
2pE+v/oj3BtvnyyfzN2Hh38oGpoG9kNTdMb/ImmVkWB2Lg2C+JVAgUqvnHfjRdUu
OPCvyRfWI+kHbcdTRadzAutVbrSgNYAc7hpUE1F1++cSwaO050JT4EL3wUfQl/h2
JaDtn0HVKLhfgIj2oAqNPhz9VaAvktBkElhpyssJT9UCpKR0m1T5Y3Y+RdUBZmSQ
9vMW1MgeABbFuESMDv7NNSANqZqI0upjYFOA21d8OCnACF9P/Z5IdWhUXjd0F9lw
tBXT/dM9uqa+3sA3BTmTB1SGex/wdb24amXE4QZDqjn4dvOOgis2ekihSXgiP333
`pragma protect end_protected
