// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:35:25 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
KB8Knxqgu/TOfVgb+kT+S4aQjE/3PD/KE77w+xWW4QooppNO9xgJ4CuoSS61uysN
bfBIjR9Ro23dhCeqvupcN8p/Gr+oZKsTWtEgrtoPCpAnkGrOcD/148Q2r1HX6HZ4
vwPmhHP4TpxO7cphTPdJ98iAgVNJ/R9/Z1xRKnWsAGU=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 10288)
un0dgJhHdwVmDV9XFXwiDMi0fkOc8ksY5T1K4z4zgrWcgqQdN2N3ZD/NptZ5RLXE
nw2fXEsX8AEAx0Zf0B06WLLt8GKyZ85SWXeqQjKSZaKUuDIflMN/hDojop2yQP2I
1GOPDuLB556gxtdNqzIIbynVbssTzJOzy/zuOBEeviS/O321VVlbIjWyYmpf0Kur
bVZI2aDHokaOeFoTkY/zCHKbLo0WoHuqChifVc1zv38VnjPsCUAJX3k3BIlYvRB+
Co3dHzpA4KKN5EJQo+t76jwSn16GcEk1qFKmQ1Do8TWsMhnds49vKRryOZPpFsNj
GvbjA38ub7800YebiAOAJUvbA4qNMkkt32tLQdryV6HO3Hb4aQWyA62oeWfrTrHa
rQEMoKicfYUt/H1o27AzpDo8FNc1vhKwDh0xdDrxsWM9CZ9GafwFd/8/lzNLF3DD
Y8+sOk7IHMuJwgidWXzgEkH7VtejAxjU1ZkFoAS3Nga5dJNBynxhjYitm3yGzhPJ
phT3MV4Yb8dL4xn80o4cJrGrzPUy9AF0i2fVwv8jQGCWM1tpMmSKoGKBD22iGeVL
tcIIrfNEdiOhH8U6SUyPOFQfLeF5vkQjibPtWvmABc+kfDSqRZtA1i2e3FKmSlRf
ZNZ7uOjBsEwBG2/ZWmD+X+fx6zn36K+UxLXLYpU0yna1Y5I4yL68g8q6DaRCFIuV
IgRfzN9Engit2VWWjRyLgF2bLXB1mNMj1QTZHelpwwJDRmjyT6JHu4RNqolWZjum
k3KJoXEIWw91Xyal5ma02uIZjo4xBaQGhNZlcgdpQoPvSepZehbGWOwbZ1d2HXmm
K4ckvFXkDisnKx6jkC/EAM5KwOeMv7gPFpmwk/7Pd/HZcCIAfVlivT0rJRZucE6j
SeGrGXeap3dVxiEGjhH+NsG3YwgPzXuPR4o/D2jwtGs6E2VDBQQhC0U64F9a3J7X
pKT6Yxg/oCIgFwqwUKw0x1bQQDNwl3TrHbUOMiXc1wKJOgfMRSWgG+5Dc9FJE9iq
azipcuT8BnsSj0Bv661xC8ehj9Bn3GNyzRGUVE4xXAgzYzzfZIbS/spmPHJlKsiD
3UUnXNJ/fGqErkxWfR+rFw3rzyo9XFfy7WQK2PHvYVR+yePMepDVGOahjyFwPA0Q
eyrlnQYDQ/as9h4NyPUiFxd5sgjUzPp1ayX8ZMAq/CrCRexvR74MpKyi1rKLRlNl
cO/YDO8okHcHg5Cih9+nF3enqIdBV4PFkyARaXb2hKEuuESG9OsffrE2A4wfU/wL
W9mGG1tfnz6Q8S+MraPblkx2XPI3HLYIabVi+IzslG58GrVU0FuYwuX2/y6xVBO2
bSg+LJHbrnVd3n4gWbCYhOL7lXU9yQddGxX+OgsAO5D/SZQl5DVIC7uv7yEyvdlO
GaI9+Nd633tk2y7nueBMZVhE7ANZCyUkM5815XqMNml8pUfKcDIakVayleEsmZlX
p2v1Acp/BaR3V7aQ7kZ0gNsaAmXMDBYlMJ02NJrOBByMrfns4MZx7vIY5XHVVWDV
TwSB5B+9qBpsmF4yHlDGazTeQo7t5mw56MTbuF+mQF0tb0XHciKYABehfTZdMtTK
ZYPZPX/yf8rsog/IdKg9zOtggwwD7Lnxw+3v5yk4HtxX9Sk58VGrqGpvCVUpCtFk
aIAY7ErbmomhQ7E/rbFT3W09NZJQOzcAM6PeEHoPbfWba7XZTtZwV2xEcE1bFREl
RUi6P2VWv2TqTwYvYJb/ggSF9uw3UDcRX0v6Lx/rGtd/R1FFAFc+x/CHQ28fXgmY
40RcH6Qe5CWsd7HHQq6LOzfMXMVQS9LfO/OwXOJfD/0qLmrDZNtfvYm/5KB5oKZs
AAVO+B++peM7552MKgAODRULJwMsIuylJfqsLbjKQNaketrUsWv++3M7xb4ttQI4
fJSqRm1uk2lUboXb8/SJxZ93gcNDA/hpfFwPWmLO59KuN6xt46gbc990xtQhe61N
0Pk5qtA8faP/0oUshCe9J6BXvdY+lNfIGuT+rgYWVBbiHOrfQJFPhL2bYIj30YFd
HrJ7MI9tly0uEGtxbU2GmEvJZBL1B2ZiDh4WkYud7NvppEqTaPZTwJtfDzY6SLC5
AoIl5j1TATdefSiHyR84UDPWa2uESFyvGIseIsjwRwTOESuBpHIQHIzwNgd5vAJw
tOzD+1Q96uKg8DrIdtGOZsl8oluMrg3QOtLwSWQUU2VvhjiSTWO5HMFG47zC8haN
bDfaKzd6ZfYpHlOlQdqmBTgKI60VudDZGpbxekCSz2wRsbPzU0bWLjqCrvCA1DIR
4MObueuimlT55JfjVeYBU+njgI8b+CWRvZ5co+dLYC6YPvN8H9cwtniJWslDDDkT
6LI+xz4WlUfO37ROmYqBlLtUZH+RbCAv+BzsGlQVCVXa1wA8HNOK3Jm9Zu5Sbr3Y
iXwc1HjV81uY4O7gtHiWgh2urdOAmaqyAFEYkmr08lwaE3XxKm78W0TjviuaNq8C
3xj2P8bf08UOy6HJPc8+rnA3GJtm/DFdaWQFLWj1tIsr7J4UjGiQmdeqF7rmAesZ
dJb8y0VO57t/2M7uVeyPTEL0G/hlkfjDGspIjtwbRYcT8iIf6kDdUJ1OofxRFKRb
eQzuSj8tT5Dn1WJF2dxIJROS8nTfa0oJo7cXrdif+RAqk57tscq8G7DIndh1oU3y
Hzqr73iYv2XIbcFwcZ49TU+h6/LmSfQaz/L80efuJD5u/Yo7gOIMOG5MvkHTZtNu
bPYX1b82BLxDfCXrV7CiCHC+6d0+betXadv1IjFo4BQ5Bvm7jZnwGa7JmDGz0vED
aJiib8Ca/f1C0oDF+YezROcpWp2zIokjxgKgiLBkI5MMVzRU9LiVB3OeMDs6XNnu
E6EXQ0PUYjwQpg8WefNlrW8++V/gUfSlrkWO395Z9+9Kq+RK0kO2PZ8MHlaSR73Y
PRCYGFyiEqkf0JbNZxyCqrzsMd20zB0AMJby0qHnmTZFsV4fa6GtIm8UfwhdK3hd
xCyrb763GLBuoh+S+GPc9MIOZW4xb5globxX2VAFp3QSM4Xa1yaKO/DkC6HPCaMG
aJerGviVxOLwoDZjhScOP9/3v7ztYzodZh2F+I8fmIyRdg0L3zAZgReJLESMeY06
fhDp+RoTxDKkWcBZRrkv0iCWUxT1sLZGZVBo16g5kQdHDE39KmHxVnAuJgUe2/SE
X/sOqjiiZdV7J2Bw8t+JC3Sp9ZmDz5PiVrf7bTu6tsJnbNH/Mhx2cS6v3P9uViko
YYxGRdUvaCmS1noXPdMy2MZRY/1HUQsXy0pEMQQsF5ZBfTEDbXCaY4rkwHC40kO8
aqUTUY4s1NOD7kv5PRJPhiCwAU3yy0y64R1l8aUwWbLXJ182s0AU+lb/yk/yUq6z
OW/UUu58svNklyYAEujbVE9EQ7/xa2S/IjpOyG9tURInkGNKfbVkFSDOnBNBcxi3
Gec5Q2GHNVhorCESCSYtfE5ysg1eSnBu2sOU8DZSHmsUPPva/9W5jb2PpbI4ttwr
ghZ03qfb3B+uFV0YiTDxO4+tXNZxluO2g17ivHs3iEgIe1KgDck1JUpctQYdX90A
ocU2AyE6dEpxdy5CvnJdQ710FXrQIvglAHJQ52regJHl3RtjvlZcymf1xAE8+x1D
zqx5Hbq1v8bCvrLDU/cYTbXU5gDm1H9pxAHXkI/pvSuOapeZqF2k+j0UDeoJf/Er
21fSjc5JENx0oYOIKzBIP01yz6LsUfrozgWWWw/XCZ1Sn5ggXBpeS2cnfH9CD5Me
Q79IrKuJ55KKEz3aXnVWArY0V6oW1CQRkEDaMArRzeUMJlGw5BNXdOVmiSgYoMcn
ro951EtbZMTTh48yU0bvADZsiV9ypFeAUAa5Z+Ye6j0NrHHX571r0zk6J4JZiKTN
Zj/I0B34Lx2rGyISqRMDbjDEcIwRH+XxGoFCw/SnkgiOO9GW3MT8ZrtSNWpggS37
/TWAWT9DvqxEchId0D2zOIpY1m8ki13mfRLZ1p9WOw9RV0druFklKDYpwHbtPiIO
okr4Rh9n3I5JrvHYUE26xNotWJidRFPjMmvE34IpfaRfPG/7Yk8qb98MCBpR7Sit
T68gkLeS4rKWeRCpVxwVNQsuKbImsIl+a61n3CRzCum4TdbZvqlq28YZwpaz9SkU
zboMAoaYT7iVO1sERdbWw8yi3V7Sndg/tW6/26d20ilHuIhkz0eTdk5BAvFQ+9LB
E6646hjrIhdXP3hLdsSutTBHpIjvsqlniF44J4eCaAT99xHpYnMl5MLQJEuBlNht
vpSPpPnumS/XhYxMSIFRCA3HVgSqtgUoZmYrOZ5hqvHVGZArsu9xFKywZIT/FyGL
vqa4eM3Vijl7URoWEGlFHEfbI0P6z0wXpUBK9BkXcLMuj1mZftpcJaXE+aInnej3
8Utoi/q8jll4Xw+cqIBMUOrXxyzvCWBbsrsgDadjgnKP2SS3WRAvwtaxCBTUolbu
98qF0/wdc9AspFEpCGpfcvTttL0BIiO+lgJ0jlIslUGOHY79NKQ6iX6pY1aN1fgk
7pVtoNQthJKQG1ICp3jvdOP/4M3fX3LTHA8EJYG5S0MUN23DgR8u3jsvkLpPnTOv
1rqcpPAC+cR+rwZ5t2G+Cn3HVAUFnLVwnOQ5WVoaCUPHKthbUwSox5soYydeALZX
WtRAftSIPogGjic8DZzlT9HdHNK46uUk7YYeTyN+ELC1wo1zHhBXrj7t15RBTl7v
zXEOVGjv14OHbRz9UD1pHfUJ8dMw3ExbJ+3UwIjmu6lFeQ3Od2pnM/SA8U6QVtuD
NxKJWKVwkAGrwIFEGaoVbIidSUaXMxFZSo6SS0ROwmQY1FNRh/8MrtXugrB3EwZm
1DBzcdq5u9UVpY/+3DRko1P825fR5bs684V0D8cfkUT3t63Qrtobk+yqj27Etvr6
tPGlaTBztfSwP6TRxeq0969oRwfbAnAfhW3r07Nv9tHqj0osAYCB89iyJ1BX1ojY
9yJuNWaWo5QhLaLkkibv2irMwQX5nzDn/3yt2x94CLZB8wNkJFEexB2K/MEfTvaj
DI9Uc+nrFKEbS9puq3ZWoOZkXtgHA0LhFi6ERx7wTDq2f6lFbzZllWxzxkoYC6bu
Zn8st2ZdqyAKYdo7O4332kgj2XSk9RqgPxY8yHtg0I1UqrQBgJ9fopqFSKMTAMv4
45YqWlbS5r5eG4wO5fyaKh+sKw028MdYolC28p5lk5i0LQFQzRzsxRf+7qRkzl2D
z9VFYrF1ZSdfJ7s5HlXvlx4JRF6NMA0K5BbnFauj66mJdolRT2dI5wyOR8/s2+v3
/yHpaM7ddgFBOLRq9QkdhX1MJugDi6gCPZIm6QHD7tG8RI123na7c/GC3FPsqhwM
5uNkklA1fRUbivVZemMIpw29TVS3mk2i+LGNm0r1euDM1ECPJNk5p2ac14AKiU27
0nsIIEG7eTimwxQO5U7mLTgBWtjjFRV582mAKEA3B4oi+9FFGi/yFupQFP2tFj1g
ZGcBsf2jSdd8UFqAScmueEppiTAfOtxlpoGueFh2VB0ZtT3ykpZSgicTGri2TZcY
QVTYUdERq4cX8kjXeAPdKQn0JmQu1O+kIUQ84i0vM7JjeYtG60jD/6FNsfY+Ylh4
SwGum464MnPulBhfAqb8g1P2Qkfu9gaE1iUuyCWMuMg7JEcyXk4xt3EeMYBZlPJi
oECf9Dxzf9nczR3j6TR+4QPTiBXLEVJxE4a1taEqzgbhyOBKot8+eiMC5hKiCrjF
DD2ovkxhWwUYXQMxZI5Af9RWIanEMv3p+H25+HfsLDPv6NdUM7ZYzS/r+nDZmhSM
6oFjwMYEMROCz3v6GIPBtIZInA43NXq8syZOiI+LHvebhHjwmteZfFvQAxedjVJH
7IsNiE9y+0l+35MjgaItwIlsbSjpPznbEqI+p7ff3jJr9ZyisAkVeMyVzQSMWfpx
X/FuB7S3on89gnKCPMMmLK+seLGaK/dPerw2mvpj7jdHKbdDRGp7rN2lOBJPg3sl
1Oly92plCJ7W33Uu7mUG6oj0rn247recXQLIvDTUo9HMPl8pImyOwE2q4Xov9B+J
ZLQ7Si/96ncQYLi1fINlVEkNt5HGHzwYiu3V5UQ25vjdVkvXCQoLeZgzsRkFKdsP
uqt+uKNXM+B3CIDv40DTiq/3QmCevcp7oC+l5WACLx6ZyMk15Vx1YQeG/3yvuoa8
2cb6Oov0b1uYpiFBSks6MCe/Ncl5wFfG7larPJlIa4y/NcOGKD99J1/nX0eyE/LS
ebYMaPBgMghmgVfr7CNaYfuDyxisP4txTbzNVBfg3YENBMV927AZjvz32PfrOkAo
rseCOY+ZK00V+7dNcZVlHhqXs6c2MRHHVmXe/IHS4sUrAbwd/JN2HWbSCdlV9m5o
EMF/kanslgXR609c09TVWx2Jeq6sCbOibI047jz9ZDPp47aQOtK9hfqgWKVPKRpi
t32la+JbXF8RgSaFHQR7AjtlbvGgz7I8+t4v4M3ha4vGBruhtnQdhKsy/GwSz/Zd
2mjhcrob86/7wS42AlJ3O2X536uwq5K43qKEDhFLLoBOtirB+NRU3nh+UVdTfCJg
vDmhsSTjAY17SKmbesr4rrFSJ2c2itmno3ILi8MRiHYl66crJAtKf+FlbsZ+7tG6
rWT3duJIgkUscRF+FtsEUAM1VFY+SOl57nURvPa46v98zzQ/0m4ZgHaLXNt4onIN
bQ0XSWxp7l/9inhr8ZqY0E8eDZ2AjTv/NKHyhp2UC2SrKyZl5HeJ8FWPvT90wb40
GNa+RigHPdbI1yrPmogiBP5/182/s0wWzZ4FWgMIvP5mwQW4ttZgWgD1mRhqVmbd
UcR4qhiSTmwSbgFinrKF/s/MvHl/ULvyiki49ncTNqDa3aiLxqCx9Qvx7LO91otl
O1npVVh5dstGk9crJy+kc58Fl4XBsYrCQw8VBzhZl/zAsbrugydNXpA5Ski5kE5b
WTPwqrIUsk7DjV6dP9wijwBTIp95W9HWUf/KLNrBjUFjoa+3GgtHqYrZSlcPz0I2
7U8EZ74x6n6NCfDfhp9FdMz3JfJlcG6dzttSukOnxQniSRmvOnPC0VNlSGNAfNhO
6dFUPFDpBbAUVBPEOZf4K1xo5uzG2uFYwKjSMCtztnAhVRJpmXBaKS26rtv0ymFM
YSuwjOmVJoyvtteFmOL6lr84pvUtc/zxjr8Ke6kfCcca3+am2L0N8fBmTmzdoSjd
MIxl8j49kVYdrplr815+BdE+q1X+9t8/Po6Ex4wL+ruqLL0zyrcX0LBukQJrtgtr
BCZ5yOkjTBaf6aWQDm4CKgSYC9uXQjokiX+IqmicwMRg3iGZ4nx7TAxsNyWqh5sQ
ybo7M9No4AEbEE2yU2Fnb9qY+xTGMaspH2HgiZprSKGp2/0t4pMQ7lASaaY5m/wQ
j4UQUUz0YQe4uvQnO8RsZ/opqOpA8XQatsrUqR3QSidvR4eVLv4QRpQdHtgOLuFr
QZsa8EKrf71OkLEqlN1LUW8+yjdnCUzJ+gCxXtVtxZ0F3CwYlQCSt3yn1O6HdOsq
L6sPgFl0mCTuqRSj5fhpObYcENUpKcTmGYFCOquPCvsG+uSvjIxfYSq1CGyULaqt
VAkEzqHdGi7Nns/lj6PGHYftg+aDy4NAWHRbOFLUbC0UU5trKW2XD8TGQ63gAhDa
MrhbfoyzogrnA1Q06vPsi7sO2XAR35P2oKhJYRd136rJk6jbTWtvOZA/KkhTFYxF
nVz4yeQBiLtQ6MnyTZwybUjz4KWhRTEgt5upG4fqrUpeqJKDOBdJ/pazIBRLslKC
CrXPb2+DXhJVLvBEFUH/Cn0CgseEoWTOKNXSgzact+xFusCYkchQyN/naxTDEyZb
/Rz740ENrTHOOd14qQKjl2+TcF36O97U3fJDAQXmWoB4Yim7EJeb1DJ+4NX6Wd1d
1Fz6ckzlsYI4Q0XSqqzno7HqEXUvmyR5M72YBXA73ee6CVHAhcMFc2iHlLZqro2j
7cQTtzzxHnlaTu8kShcs5S6RyyeP4DRyNPn48QERSxZT9e9W+2eji+QmCp/s/IYl
Alz2QaQJLXxU+HrD2BZOvwoiHEG962un4nDKW+W+pjyL/Hy7qDfzG3WeCzadsRpQ
YWt6a9F3ufLfDo3bU4lopZGcEIhshjcfbeWjajcF79PKsqWvbfqp8HYftf1RF/pz
AqiUoPiSBWcrojXwBL2TngK3LhF4W0Er0clZlW8d0MIfgfEFz//POF+ya5V7rm4W
BI0fjZIdHPzI5/SFXkJWHqGxCI031FJHoBDa3cbROWyDkxMaUROtYQEz0MdohWgl
iF54JQtaq4KbkvwO2aWG8RK2YX/rHBtfGZzICl7sphl9yItQJn8IlocfrwF7P/ep
mbOADz6/V9krEq6NQTJb/R4OkhWOHaPHYV1Tmiwvv3zwFOhLsf6GwH121EgG10vG
sprA6jMpxt7Lc7flgwaDCHxv2f1GATSAY82tQESkf8nx6YvyJe5e7pxA5fszQUIX
MthNPLb6LOYiz2yJSA6ZdIqk7OwMY7jCby5X4cDOMtqV/atIgmFYOGXe4utJUdvl
qgSMw+7r+2TxeQz6AnOeB/6XBW1Rkj8mut7cq/m0hOGdXYJXIAVPY/kgb+aZucAR
IiIxHHQtZSKlegiNuPfqkuZQ0+IMNAc6jaJ8jPj7mrMQM8dY2OMrd3Mneh58lUVf
cwiCOlI050/8akhEETzHU/hBQdKcKY2eV/zhsQiqcxlcPq9Xa8rJQDVl/fJeekeN
l2G1o+5McA5hEUssjlhLOlK9M4rRagL270eBrymzijpPn1aVe+OBkJRoNp8nv8F9
PvcNMXPsxGtWJMXkBRXrLd/hjoThTtNixHinHCXwOJxChFiSpw96X9hfqzH1fU3Z
lL1CLTSKVx+vkUiKZiiBjec5TFouKr9LVjwHtufVWA5LtvFCv+p8ru2se4Ws9X+P
gsWWSg0q9c+xpm9UvkrebW+09Qa4W5xV/FXJChdjvY1Rzs4G2n5eXqLxzrSCtLbC
oAnt2KZckeeXEClSz18uRcnJpkZSHFAduZBHaEGwGh1bYerDHR8HzETMLuWDkTN9
S3ry6KcA4NKQzsYyQdkga0I2IG+nJ3rYjA6Gxuhqzpu8ugLumL736dESdQySVtf9
TtqpWqcIP+a8nzAywquXPBTOcZkDX9oezhM6qPsR3v+DatpjQCwmHGwqHsHtIr6z
DxA643x3iBDs9c8n331Rn4smnr8/t70Tpr3SVBxkV3902A2XMmNMmv0XbPghVqx5
HN27v2C04sEdceLN0Z3guX4p3NXXXFWpb66jx9+a1snJI3kwYVrR2qMosohVt8vi
qm4H99VqykFW8tDOhSKlXuYFy0eOKu9s7v4RhH9SrvtdEXV1Kb3bXwMpkDltokVV
Pw3yLBT/2rxFFCY21dkTMel2LbF208TTW/GT06DmsJPOKP+JRlKKgkhmgtsNf9cR
Q5h+MUuMSqIVHLS5uEBn+O7WeHCavjVkDieZgS5oPXWGCTNGzR9V5KJL0btCc6TS
F2dAMRaAXqOfIkaOm3UafGMQzjj1J/VBgeZRKE/0t59wE5o+gLtpycyUBC7V8J1K
R6wYnLI2dlShL7OP3ii8TXH30uDeFZI+eHFo5W92ilw/LBna4rzyGZst6WorY3vz
ArhFc0h6LQYkSfInTvVs/6ur55Uv4KrUbK5U/mvM0WEP/FH1UtQAF/3TDyyQ2iLW
j/lmbBnYg48yYcfeQ1T0nSpeHklaUBlBVOZWvBlSUg7ZNXfDf8797xzHq2a0xCf8
QKw1bF2g4UePv+0BaIv4N/1743HGwdRM8M1mYLlNmZWgDadrMVqqj4I7WyoU2O++
iXAqmE+7XH+LGjHIgbjPhgpc+SlKnYFXpxEH8V1hXJ4xd9iRM1LwsxZ+TVKq7E2Q
URVoa4A4L/g8cqYxtA5gwCb3GwWRM088uzKWIFraRfIKDTmzHPdgeVx7wamHEwTI
L7E3SB5hibotMLSO3+ZHMEnyWK8DjTV1Vno2PXLxyWu+spUkVYFk0+TBuq7Jx+5L
Wtnos5obpnDlG74GaMJ28LLOhFuBkM+dTHMtBjCDrlS9bDRa0PJRW1m+K5im0O3i
c5bXu1DCnp/LIn1+/W/7iXpVil2QZc3wFKL4Ill3a3laDPZlG3xgBctyaPd0e9Or
fBlk9O5zOvbRNVYrVyWKraG+oXdDFRpFNjMDze7pYaZfsT5GUfQk6o8ffKPPz+a6
dIloCN0q6AsdUun7r59THw9+W1RPYo8H5RlD9PGztE5oJizoI2sLVZcpC5SVijYz
+QezB29E2BE20IFHvNvKDIXeAyQvE/xZqJFBEDpdztHR4InRYta/ez650hGL3t1M
MKnunWdxrvvyR+DCXj/yWQM4JD2qsqBoK0J7KtgCg12WH9L8uwiQ0SCJFCXrJM3t
ENZwIMOb8HfA8/PfUhQiOJYMffykBNflEomXt0OgcHBTsLvq3z/DnR98d4W3pxDx
Z9Zp4EaGJxzyLHyaT2JPFaqyP0gB1iqr/nA0LS9u453a+X2lkE53QwQ1Oxd5OcQE
fpSa2MXEd9q98fz0m/6rIafwvV/tBkOSyR6X0toJzu0iVOAyT7AKQOh1S5ZjpAwy
+x9KlvTtM9qmikL85qKSmItjm8h83o/DnLCvBp12CVelLu6MqFc2ml3Z3R5y8w0D
Qkaw/mQ+dDfgN9fam1M0FmEuhCyB51wGqDm7pU6IO/1uumxCj9YZWGPnaJcaIH0r
7S56z+qJo2ANDrvAixML2e8HiNO/9z5qZAtX9q741AwwwGzPY1gu3WlUIqncyGTn
R5u9h1nep0+yWujCVFvzuTKtjY6kqAhZpPBuZDIKnV0b++ToFAbLOWLml++lJ1QR
chqPSdzAZZrXdGp6aSQ9aPK3XTXiAY6F0b4+LNFbsA+20g/a2/4mmrJ0+Gqd5THJ
/KSKiQOX4XkkJUpELsXx0M+QYNelewHufDjsosV5G6dHn7cb1kUA60we25MhXi3d
OSAMKbdXkbg3uxUgHINDN2/M9hGqA26N+dutcW5tqzZIFDGEdPXMQ6Q0DmmIl3BH
oOzGr1pA7jjDXlmnw8WqfRjSB5PzLPjGROlpsPGreE+F0D/KorOWMQAgnVeMc0eZ
qCqpysVBxy5qW/5dB2kKpWytRjWT7RNMX6ErjiQD8bL616YQ3+px/5BF/wdOF43B
IZRvIKSPuTfnhnB/Q0XWjIqEQ5YEm1ljt226rDNM7C82k+R4hEL8/NtwrSA2MRfm
QzObb1wXncbmq+/07rSOzXfOZ1/tWh6nb1ZB+fUBAgdNfFIQNyfeAPkIIyGQAWyt
WyLL/slabVvUiNCdlMyD09NZFsy7jPrbYSpoRxsMjlpLUfRB5cZa+fmQzvakqIyP
KB1JTqdjQpQIG+mO0tTZAqFvh/ZG/XY3ledcJ/RjpeZL3U9i9J7gLhuUVctWdeKT
LKkLpr2oJqB37B7qT/DowrPrIIStCif1enVxDPhtmSi+oLYDTVmVo+6okqq/lDAJ
SVPXs3EjEXYF6fm/EmxjGnbECRAACxRJER+lfZ6tGxiQhhg1gsW5cf80SmhsML1c
TkCtndPNLPRNDK4lMMbDUCFPVTdxYALdcE0Qet3uKe7UtqCQqTdiO2umgJ8pKxIG
COznCmiC/SLRx5oCl6Ar/dLJLuTHg0HZv0tVQXdHSHOyu6pBaoEvsDvDcOBAN8/j
qJVMf6lgp3mRfo41eNx80FF9EB8gdpYCMgyUOQhk2PZW3rnu0KzPtdtQHDHLddfo
UDzGpckX5OQEj/oqbDnE87wzrZaO3nmMOn/R7CWpZloo0P/fTR+XR49IROnmLaiH
aJPBojZ+49DTOVaCMF6hNDBGlll3r+WgqbGHjJkjHdDOrziBeCMOvf/DupR3NB5I
f87c9RoLrHKKSNFjRHTeNzolkzaX51juH4d6PLnNqz8qTBi86DRZB/gX47HnS3nA
8XdAVx2j/ZkdxVm4qHRTOShtaJgEtQUlptPgIkNUnGytVra6OPqZa8X+G28Rmdgb
QPe5PGviR9ze472jqXoyetyge7aVJm5V3MPs+Og2iBi2Cd0oORXFKDLhp0bsLXOq
T92kTaEkcNGxJL9kIa4B46bNYjSodSSWaMRl5q91eXOoVfTRargomCoeT5QIyawI
xqn/VYGL6J8eKfXI1XkizAyQvxs1TELh8CXy04a+k8jIy+/CTpnCe/UNLubriEb5
tsJ4pKrvsJsknQppLCdS41vFfg/ymK7gpkn7JRddh0epoy1+D0KzmPxVF2ZZASdV
qsSKI77Hsv2lYQOM1GTn/9aGAb6kc+KiGpPUkwkYEed7tzdwFz8yTVjnCaKS0+O9
lv9D8pYKRtT19ns/zqq3TNyQK6qzUXSdLR1xjCXvcMkA66tghLcsC3NViqAiEkZI
gLMsa3n0VQJdM7Ie22fBGx1gubGeT5EscrnPNZrGB5rDYgC8UiHoIXDO4FvUSDzN
oNdRRTQP4F5dUFfQugAu+qj//pjZZDhErkdaAoNLd9q0yADQtU5QaWiqDg/YSo2S
dZTrECfBotYH8oU6NV9kDqQ+M+n/WcYNNwvRMW9fEHzmbqAVnDGLg+iJekUT3Qxq
9KeDF78FKwSlrhmiNh2Vf6SqDwHmdC195qDFKoziPcdDHFu8WoL+630YrfBRNEFW
cvMPmxCMA1h+JW+1b87Q7vGjhuXPbO6LJ+CETIFbzLU99Xf7TKR5qliHmUict3Ev
0JQQADiSgnzVKm+1+itWSEw+OEq9iM6laGDUTR/E1gezJx6BN+p4K5vcuVfbHg52
JRxODk8GhTybMMTOf8LzBJq/Bg4DDnM7/8LcF0UhvmKE1pl3vnS9p+Jw2fGlxBlI
710UvAvbjcDx+FZpQ+zMzMLrWnZVNJ06F1Ut5ufBNA0zdRq3LpZ2v7DNc6vOS7Si
/J88oz4lC0DuCpQ68pZFHL83CRAPl++NFDBz/IS5EeeVYmrYUk3OfPbEXUJa/A7f
rr/+wwHGM0rz+Kx9Am6VbtC9qf48lp/agfS7eG2lslk3MoH2Zi0pSaWnC4/dkFy4
bX6d28vKyfc61ymJwS4KTHyilZJZSyplcz6H1entISqYkN0d2/MExnid0vBjF/lK
gRtEoYN2Vn0Aw8ZsMD92TEOqQlrW5b3kTAgIokMkWTSBIfFM7I8s6SjWz33gjZsE
ImDJfHUucisQgQDn/Qlx/oA5eYS1i03FMOo7B6CTLCsx9Y+pMphq91g2PtQoJxCP
oS6fpCxmoLS2bMl5A3VUopyqiG/WScm4aZ8bhWvDr0jBit1DmteKSrCH52psBCoq
FDZ1ynbLlsBH9SHYqKsGynolyErf5P9buEVRK+WJ+15pUrwRaQmm9YIPDJPjGHu/
QjcI0qNfhjsPwcBXUHRD6zD/xViubsA5+8VUGUAA9trEsE747CldVPhdN3aqIEMq
MhEeoiaHMJb6pBju/EkikXcjg9GMDncLyMntkvpucMUUPXHvY8ii3msij49R1tNZ
t4vEbXxE1mgxsxkIesHLAoYrWL6JA1vVbAdcEY4fVCg4+yqnb2vwW3QiGAJqKF93
0BrI3xVAx1y0FpEEwnhFqedHYbLV0wnoqYWkATOfyPSSSyutrAtSkvxdFPYLis3c
Pjz+r1V3XYpqDhUO9G6A6G4cAX4KPbSUnQ9mkVmgjflGpAXBTE1UX5VwEVmQ3T19
qdvSS8qFmAkqOXtq/OBusw==
`pragma protect end_protected
