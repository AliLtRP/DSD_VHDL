// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
QBlwrFerTOPZhasm2GwE13W/WIzyLDtmiepLb6qaRT6VRFsE/+T66ghvYuFdmxURTHaNROdzTRNr
3h7bPmToyAiSqnUBnmqN3ftpQsjUZpuHXpNztvRxp1f18Rie+OL2Tjw8WspZQIqVnVHGVpJseylf
EGiDZ5ZF8JLKNdaSqZPSbLHgGQxAcOgNnKqzN8Jo5sC7BcB9qW8Y7nVof1HlXNcUK620gA+/7W1i
fDjNJur9BkCBRK3armZ9ITDt3n9Rx+eMFrJcs5sa6/fkB04yOKd+hZ8D4lkKPeOVG8Lucq5CVVV3
L3hbwQONkBtkHdKIVJmJegV5xNCf636z55cgBg==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
l7qBjtEzTnelfcLwwZLPT7wT9sfobso6i3U/zcQ15UdeMywTKlggJSjiDczJYnm2Pzx+jNKt/kWQ
tFwp8HEkcXpVOeagM3keL9t4hZLN8jv/pJCHgQOo1npLPm8mkC3B4fc+6PC78d0eHhppnsdhQU/+
Lon8Tpk6o/p4imWQ0SqOTj0eNISfl/05vfGEkDK+P5+YK49pTs6SraWSnu5F8BtJiWiDukOYHeTN
jyhY6dgyB3gx/dYSlhRa9IwKSVcJTO1YbRzj/cRUOETjQV6NB0S/j5Y2J+e5TtPeV4yHQK62oOj1
lycmhmkdsbnArGG5VxcSD8jIcS3jGf1yUrcdG6RveAeUyaxC/snTd4Ab1guA5aY7qJubMhavnL+A
6BV3KKSwHKJLSzF+w7Q1kAp73OgBZAy6sJUN74xIFklGpZqTX/XwtFeKXfbYgCeMbke8kkibwI4c
nggS4Yvow2dOCyISYSsHnjv2FNaCDanGKZDkF6J8J27z58eTNmOFimP0h1hUxkrwLtAr1bug4oB9
0I6ZuhlbPWfho4ll9TBEU0zLU749oejLYqkKDIq8BxHD60PP+CPs0H2l4foreFlv7aDAbvMj1v2W
RKQlp8SivDprEn1dHdV+ee83GaVVpVnHHXgZGde3guREg6D43ISTTicryn1RITfnuRIVWrBOKS/E
kTdSDqKsQ7v1bzsVllif8jviRIi4sVDKfIAsGkPW8VaRSfuDYLfOAOV8EMEof8vUk2rZ0J6SSO8u
gzqOvIgCY8oizxQrZQdS5Tv+rWmY5i4X3FyDzFFbNINM1XvNHjQvU2PzcVPWkpfMU6Bah9zSfbw9
A7S5a+5nZqhZewYKaECmCZt+LsNnIHRnyvFrVzqsoodU32L6cVvUeT9JJG2sQXSgj2eSuu40Ug+t
qnsyDtkCJ/AfIACOlLudnL8ag11lMO4pb7wHvwEw8eW4F5PPW6lfRNVNFEmlOZD7J9w2JoeSuNaf
DWTgX9dbulIIiGcU2d1WCIaX2uH86dTYPsLk3fqUzcolXql7VZUVuYoIggMVbI373Bx6mi1ZBFAT
2qVxTIfRmIseeqAgcfJlVIb3YzVtdK9yiMg3kj358/ARXjyS+ueTOA2UEtBKicRY92LbM/+OcZPf
VEtsDVpXMbCGCT2/RmSwXMDD0T8WF96+OMqUM/RsuYJgLioz2tbb5wAVFkYaHjtmRFgwFb7rFR79
ruVSmLZnadHoQ5zmD6mi1X9QzT0D9Gh4eOvtXc47zNf2RMh4Cy4gkByin9oZr+L81rW+2ZiLsvpg
hw5FX6yTO52l9350XZ62WLCJmhzXWcChuUHyO9U0ll/3C/ScVV8Lld/uqrlQGebbl1L4dcJk3E/C
bzJBgwbntR+naM7Jniah4cYJ/to8egwVYRwYQ1CECP/XqVgDaM/odj4jJgK+FdCX7yEC0Ge9nvnr
ngEynxY2X+ByS0NYT0Rj6RzIWGxtHisBnn/wFQMrA9lVehd8ywaYB1kLvG0cmWsy8suTOQMUMcQc
7rSSaS/Jhzo8Swy/LiErare/EhtiXbwY2GOHyDupqfHCtexPk6xLsIFxIUu9a8PXS1xC9s+AcaCE
G/K9DeyeKf3yY1/f41pWMfTwb1SFxhlaYCrsBhtBe3MmkBy+ZeCD9utZXTeU0gULs1sL+Q3os29C
hxt0nNmTCpczSOO4RT/FvcgOsEgJed8iHKGkfZttRGZeW14tOUzLreDAl5okD2K2bj1wSpXAPfxh
UQK/9IVyKEs8aRe3C9M4JhtMfhy1KMuaA51ZzU0Oaanfpj0Ocwt2kpGv8PaNWx73rOezC7ckG4s4
vNON59cqSdbWReKjtpKb+Y+mtOt4d5thpfhxPo+xZgno5LPGwMZlix7se+1c0WkFx+GtsYUFHOA9
ijLCAGEeJCHxnsJ+uojsfCf5/+22V3csy/LfHAFPIUms1eHAwh9DlGJ29UuwG4UOCoNc3eDP/DUT
C18CLGoTwIrvBdJXHJzvSWixonGHkQ0IzAZHUH3pl6vh5cybgBEoNRZ2kChHSDS7MAkBXYsS37JS
m3rEEPOSlm571g1fJ9mSI6L2q8zB6JHZKxukk0nGX4v2pgzuHD9Sp3ocAv1RB+8V0XopICbgaDDw
lG2E5z34EMKf9VDnSh3e+wVlKWWDopgM3/X01MI/HdMTP38ay//D0AINWd4tF/Glq+DzbUbKOadb
gaOFEl7tS45fjD+oo7XNKItVyr/1FUGoVzQxCaUOHZ68zdSvzabJ1J6Lwo/JR07mWCOLdyaK8eba
OteaTHTwnAlk2oqhJI6KcCSt2mesKCRDJExQ4jvwLIuujzjQOO+inRjz5SmUadANl8LNXhr1lc8f
L5HLbsefAFdxdECm5WnS150EJbuy/0Gz6c8EXyC9G8ODf/IV43NGe1sXDOhl6u6njLrJ7oMOb4bQ
QMDKg7JwVVHrc695o2hMCgNMNGUKqxdxaPGYD5vZZxcq6uWMKowfeVgxk29tbS4oA5BOk98YrMdt
8o/yv4goAwmJhipr+EodY4pnTIQQAny+ArkjStsYKjO3E9Blxkoq/pR5RIeKX7kWiThhbmBXQbL/
wu+Jlh0Hn2+tzAi9m5BN4QR4d2ye23DJXLoLLCq9CNrN4tpqWyIDyTOZ5WQRfrCMyiuN5sLcDv8K
sZpf8WQNh9dl/dhE+zhtJrmVGF4PoXm4ZVmorB15UJt3gA1snDYwRaPev00nptGCZs1tcA0EPLsB
O/rBOqx5u6tErSrzKz0Il7McJ9tUdIqVIbU4k5qq1TkDuvBb1j8H/KXMHd7dAyEvzs472ymdQQ9e
k+hOdUbCn9oU/cNvot2Rj2svG9IljBBpAZYHj03SvUf9+IpYiwgJ0QAEh48wE6O0TfyZqHWA0Pyj
HmXegSlgWazKOdazp0bRWnsJzzB1wMmls3tDJT4dLjO/zfP/0nVemsX0MGm5RZGhW4/Kb7flrxMf
pdoPkNnnWH2e+IyKweJxZy80aAFtkbjmwPii/ozp8K8/Bml96v0YK/3xJTqR3ylxaOQvsNBh5Bas
JQeWuS5ZWb4o2OkHTa3yBF8Tqy+47xxvbWOBrJ2rp2z4NgTWr1Ws3/NxYUnxsEoMnZs+VsuktLgR
F6TBFeGF1iHiBruDM+gxyQgJyFQACDWLwWq7qqSeUTfarmLpe01oXf287bkNP3ExofGfq7c+ypzC
p2Mpu/0/v0a2JpaNcpLqy6MKWIPfbsVT3Oh9wbCvFvu3APjR0+svsLZ2LtJCZnLoaCqLZok7krk6
9SLuv9Ptjjx4OBMaJtvcXmeUpI7Q+p6pqHVrtsoWP67XL0TOBwyPxRRWgCP1A/8Me5Imj84giX20
XAZqPJunw+qJAR0W20eE815UObcsMegJxN9cC48Urd5HmNDwTQ9Pk9isjPOOuQi4LoevujMbFM+G
TQnAdO9TKcakBZbLORa5Rij7a5LHPScLs6/by2oy752ZSmM48+zSHvD1Dgdo3N5WJM/HYbLdzspc
gquPKl6AfnNXH7ft+ZjJrNkQKV/lQvhBbdtIK0MWU3LAYef+nBorzEJB2KrLVVx+4mUSct2MDknW
jgIfEen0YoL6ilasnfl27+HJsuX3Kt77a4tReofSU1pIpVzHgPZFelv/+CmpuNhYKjz/snUnf62j
24BDRU5PXHzMq3P8zbl24H/JEE5R1xDQMbbFD9WAqYLfZo2G8d/sjXRvhgtidM7jF88Nn1sXw5JP
/Afsmnz3qvcgcbBHfvPBLbIuKhBtl6oNkjHRwNqFLyx9fpc5yTOjYdYsxY3FXfKDke6rHH1+2qsC
8s+pgF6nge2xRCefNPHRj5ZmXQJQNuClEUSMiRB4XhuIcD5g4ByWn2Jdao6bYinYvBvs4PdO3Iev
aGiA+fQTq3EILyDGB9NdJODxw+nrhUjJNjdyr5qqKC9D+BMovG84hBcMGkVUOROhyPHLpf0ycZYs
9rAS0ZM3jziC+jCjtuKdFnd2iWOBrubC9iu+UKoksBAwxAYQYiujWkUncmAOYeynOIhRiYu3V7cw
y5Ggx/I+Ui5l0llxFEx02Eujps8OPwtd+lDC4DmmB4yaTABhKPkDHn+6ZKAZR7wA8kXQJmkEv/G+
iRnvfyT+kQVeZYy2NdUeLFI0YEe26/a/ae9kEe88lFIkImKm0Wg+J5MWT5pK6LFRCVn0acNO9MPL
Pk9/lOQzv7T7/eTVbVNBSj7loOMgBIqFyhylNnV/hq0p3zCqxJM8epKdu2D3n2OlgEL62IoqYcKu
/7BwXsRR+sZAe5S4K4yIBCFZlFb2Ej0PJOXJUfSXfmCVgI0GmNmk2N3f5t+X8bnJ7jIEdqIeyUAt
H9gDGJ0M1jLC7thav9g40KokVxZiBgv2/YaJ1ZRiGX/SUXcbLnGGMsIacRe+5xTTYUllfRB6LjBi
8Aq77wKzstvzfU1P9hJFCaONIauQf4A3f6bAoJgoIlWKZN+G0DKFfKbcK1eXBgcMBrId4AIXpgDP
HBm1Hrt5+VBLN7i5qtIr1CtObcsxu+bYGlEkcAExSYJLDE5nAhtbT63oVhkxisJaLnoEVL854sRw
Avx3+7pV/BAZEtFGn1LKGiEwkz+NMLMzzfTq2R0hr3CLc7mW8YktvuKHwgInqHNL8mg91CTgUnNY
L6pNqoS3kGrntdlPt+VGg+MFE54fw5iQpMX4lbg/cGpAx1BafO1T1Yq5vLrh9s9XsshpodpRJX8R
fO2uF2c8HnLNzJo8bML8tar9Y+BUsqOztoCZ0yLRBpxuKl+oCbNuqlcZMzu41WH3Y6z+gP5RRGBU
jYnJ1kuUXjY+syH1gnoKR0pJayICPBwHOjrixFx4ABHWuVXNsfIHlJY36P/H/5HYX9fFi3KMnq3W
4jaCazd/LYXpLuxfkiraGF91pFJtPpR6+8Xup7pN15TCDpKrGaNAi7/e2HGEJ/B6mQRY3yEPML2s
VNTvchIr4LODL84JRnxqANRMnPor4IYqYCyx4hE8p3DgaiViFRA+69fveTMXCYkjgZ7Xt/GhZpXn
lEfiUTAMEER5531jXxnVENJ0VPdecOlxuwjI6KzRt9990jlxboEqVtWdQb3Sox+OZXrpRgUrW9dh
h+TsnlOlw0SuE6dEq0q5+ugWOlWDug+ZyKEvM6V0klBVeFdHjqRMAwaZFkLeJn+9r4zzMe5L40be
/EKKSyE1GA0XAnBvn/jQul3oGLfMBepWmZ9kOm1TWzdRV4MN1IXCOMzFUzzXk5pWqwxNaqhy2Ewo
UrV8NC3l3fspGz5tQVu9pZILnXvVFSS5jMWL4aZCY3wTX+r+es9twyNrfkzw0Ira3r66Cp+mMRGs
tjVcVjnIplgDzG4pBXaxiJV4pzav3TZKLYju6X5T5ln64t7uhWVCbjFFYoHQh7cjTZRlXKjfvJhy
itLxl1GLzzajtKIrpjziyH3Wp1gVs8XxuTs+Ps9//l5LzbJtPz+1qVFjWfdQjjqt/7cgzDxIryUo
pRoEhQWMHIsP/2UbT94FXOqE1xW8LWZUQl68ZCvYnhxAhH3kn3BitlRMoZfJjeKaG2tUONS7yiSW
ijJjv0YVQTT9Pqkx/porUfcwHYLcdr0SnEfL8XcRGfWxFUuoDp7lJ2fsI6iR1yMSdcNQxap9ynKw
pLtzGZf1xJqxYrs5XycicePvlz8FmULJhRX44IbK6a1BpjiYXDvAX52Ag32WC9RghDfOuxYj5thK
bHRvtCkXMJtYViUKW+oiKpEM9km48Mhk6xlZCcFbQ6GyW+iVqtw6zVnNqSrg97vyfbfU64unwZsa
Q1QOPIm7JMa+Y7qAzqh8REQYfEdam3JgFo2nlsNIVKokuMV4R0Af5qRC89Wq9e5hi9GxvLL1Jy97
oZ6VC2UZoQIG5waCS0Yoji12aNohfsubHwMHG8r92ZZV21dqYL6ahYDpz1PnmIzx90Fsmsh3pRSF
+PMrpAnF/Ze7vdNbjLiRjaU1qQTsVyVt1gTrx0hLJ3aKH/SrIQDxlAc32m/PXxh2ZRt9N1wTutqT
S6unYRiYHMX55n/vEVMo9i+UPPwDr1tCMlBRCZYUGRl6S8nA8d5/7y7hsXubBD/Lop7iByJb62uX
o06CCT3Cq+BcrFWfAb/9QNO/cIF6tq8ViazLXP8ub5/siOXSKe1W2zYQUBxq+xPKUwW6FhckxEq/
0ro1a06nfBiVrZRpQkqWwiGJBzTN7GJPIv7ijOZybAmYnd7hV2Z2Se/wAvf+dgsvS5hhXDf+B1te
gJlLuwtjMkkYssSCeHFvc00ePG3atWcyTPMaaWtxhDPz1E0OVQBVULXHdyCDdSdJrUc2EzMZPYQR
seldsKCuvl79XwWslhcKTAK9+ROk/fhDxe9PTG5KG9LjP1uyo6M042ukVuH52Qn3l+mLNyMxLJ+d
qin6WJ9OnipZjKh4tanUu27x74lGYlphQxUGIlYMwsK9ziWcQL6VAAyg/icLRdj/MMJppJPiKvyw
MSNLr/nBuwyvEKsY/NU0jeMRvbPG5Gyac9TaiAMklr6ugGudoLFRdgJrBz5zRJlrRqd1XQLZtc1c
ZUM/1M+ZNNmf/mXuem6MVGe2mQcEH+gaWJVRASi+p+5V27tfwV37BckCs1MmZybOFFIfbHmd5clD
10BbR6AQWC8xot26clK2Y4T/HxEW2imgiGfnapM2Q8HD79i5PoKsluvrM048mOiUkTJHBfkqfTRR
q94gjFVaisiflWtF67sVjZZZFHQwBRFmYF7mNS1pbLriJp95s2og75bRpB5MylKcOm1gWFhfvKIf
rl+PQC9GC8JyI1XmoYWcGoj2ocWjcc4ogRkQDvqHkOx6onXs7UGoOweX4efMJBmRU2dE/uuliRHD
JuJ+yDjL5afv37z1lPhuyXsh8DM92+87iMGeB9XbHPlRJzgoWb1cdDza2rQ+hEUVKU/4rcdazTiu
7ix4ZhPT/TaQlrZJrwlKPZkKmASprScysPx9U/oC+sWwxEp2J+Mrzi+iNcR9O5X/1lp5o61nzgD9
DG9XoS7ADLZAMuEIymlPRUhQ2MnlGf0nBdRUHZ7jiK3Xw2jB4oGeRod/LhdiE/QpR1i2cIvnSdJA
7juKE4Y+SLCwa3ZR42FckNLKOYCShgQRozhWolzs4SPTHFmSXdeY4fMRXUEs/IJse0CR/Uxo+Sv7
F4ERhzTxmwsUftuf2EzNSmp438/V0yeE2HDmC1aKGYKKOXUPtNexD0bGhk3DC1LyMjxQ3//ld70U
h76TWSq+1y9h80c56zq7EU5f5jHs1PUS+L0ZUaGYmzh+J7S1O0R5syRygqTGkKqcRTV4UCDwO4i5
bh7bNkJ3fv6YmTJJ31iRHtfBGn5y9keTLX6zVz0ocvgS0oOPgxMnmrsHeGw8QHxzzTZsb2M93hEb
rgRTdCOWUJwc384UU5iTgneBRP2Xldabavzi48WsU6FQ/zsSKmO2KMmAdU8C40vRAffzpsEFVkU0
8EpPMwo7uk/q5+mamvPHBHnxYkirHN5Iq2q4Q8oJ6wDk0M2kZ8t0+wuE3H3jORWRrIO9XWHYCLT3
OeJzCk2dO7Mr9wTM+Vz+KwIzWvoKhPiZSga1kTlY0zUAHuKzGyPEAC6Yb/IL61Ya07m1e/igovrj
tTRJTt0zZ2oi1vp6v9C9K/eHuQ15FRHBvN/caabEELFTYe7fcuuqbusfGqovCc44o9Tn67xzhvZF
RgUr9RqDbKzfKdwCkFC8AJncSFQ2Gpq8U7vHV1btYTE0ZS1GEuWguzDpRz9sOLEoA7Cp8OcoaqX0
oxFhnFAG76L2+yT6Bq74aTkANIcT06OgIrGFCcNhPdluANEgKaygJF21POCM1d2c2g62dKtwFtdD
aNiN0mvSrgaru/cFSGiVhI/D/cpNY7JvSDHQMHOLzVlJNezQvZqrTq9RwfT74JpUqUcleF1j8jWm
StSYwqaUyWcI3NSnJ+AodHYa6IYFTN4KyYjqY0LBLMlViRQTwf0xplTWmPdDx980EGd6d719DVUc
BAeI5v4h0R2QLdEH/STpml1a64fKE13QJBw0qaH+PzYn0fc2x0FiU6TxUqZ398albDnrQPwN9dXI
gkHb7M58gNrv5GR5smFekgW/an0B9GehsL3q5gRgYoAAP2SVn4D7fuZQvI2zloxdT1QwvdFKFu58
VUagm9EdqYthpulXZNkHO6xbBFefJjacf2XhTjOLK86ehFwkJaEoGU4pr7TVx530SmSFyoYaz8L5
pXerUXfzXiBbm/gyGAQZQPwr491AV9RcTZB+1h+RdeSedovk86GI/U+nVCsgqe4M42wNFDsMYtSQ
lesKz02OXZJQX2qY5lrSqiX6vUYZR8vkjUNIY+wwkUVFFgSZpGLx/OAs8xibArcpslmAHhApMvYW
U42IVMFLDQBh0+jGJRL53biEeyYk0zWHr5stwHrwj8q1NbffW6ukiJwF4CbSWjPlukqDaFcref3s
8ZzUqEOilpL9DlnxGBNdi6gTVlyDOWX8pTwjCKe1YSbyrgBi8UpY5FurQgbQzmu49bT4itd4yfmm
neMEFyxNiEaPJoJaKQ9Z0H/OutG4Lfn5mwgRidHG93BhetTqJcC2WjUD98Zy8ETkqwlJGfeedG08
f9jre79u+XtyWJQ224I3o7EeD1UtSmRw6XqUAjpTNtNF9bekFpMptxaDeaUzD8FKX8BPfu7u91uL
WkKogu3+ESzhL5snr0ZzXpeNr3Z0DoCViM1ewX2ayYvbBHRTBQ6TT6RFQe6in5ibqtJMAeUqrIzU
VrRDA48a9ZOJrlDbz4Ah6DoQsNGvmKM8RIJQR6FUuRX6s5mrkaVA+XvFwH+wOGJbxFjtWc1dK3nL
gcFUajOKqetivW/S5DfTgYMfweR1iCe7uvgTh3p6ZRNpiWnjI7HxhORzeitimcuhLDGHFbWDE/1V
821HLQwZLwz5CPGzvTVZlefZnTFC5mNxZilIw2cWSM5spq6TH3/TqWAgxpfGw7QC79nmBdgAWQyu
E8MfkCsBpWqVUdaTRbzjm2/QyC8krrBoU4bDwJA42TaNkonMXCLXxDwfp4LpVbRUEG+pJODg26KR
Z9BSLoj3IZzsqntrl49mo61qEIMG/oUm1KUUpIi2/IE5T5zxSzrJqP0bgtVt2XuVWtfx/J3dpHBP
EV1bZsmW5S8odqLRIrqGUA7tCNwZdNteW+Oo57Br9GSZ57JYgKZevPf4vQi/iFVWuPI5lEBXH6DW
X638La3nJ7z6CY9pHx+nNQ3byKdkmfnLwOb6N8zXAyhag2eCoZ/AoKuuGvWQEbSknBAsS7LVs+E0
wJaD9iouFDrRGA+BbFb8An1G5b7s4uR+euubREHONcXu41iqaC2y0w/1QBv39rW6lvSA8oGE1p3e
g3IcmGhfSLoq4zMVI6J4PCdiv9F7Wdrwhdan2zqyLvMCMSBNvKJf03cA3d55f62ktt3lTlkLb4fJ
mcsbRwG/nylnhzYB746rWB5kPqK584h5XKemIakxFbSuBh/dy2P6zjtBwOauf9UvhbRzz93MaZxL
2dNCS6vNYnzW+SHeEglAEl6oz/3sRAj2COTirj9JgeGpCaA1PPFK3llXDT+YE1/DGZ6FCwyXYRkp
s4aWVvX+c+xKeDnxu8F+h2IMfthfTRdPJlY2yOw7P0tXAajsOKp/SAtQ+Cu8N0vazASWfJfr5akt
fud2i1wPsK9WPzUtFsBoJfja7jYVH0hRM3+P5ORTi8tO+0XU5LvYFMKBw0z/arPV1/e+qqcaf/VU
+rYF4q/R3bxbt5GG2yDjnuzLrGFTt9cvDOJzU2q1FOjC5DVfvMolwLD3GMEUR4pAOJK/9gIxJ9gJ
FrSztqSVCdVIGvcSBRhWBq3hiXMPxsZhPVq9GF0pa4wgXqu2FLOvLADD+iBjW5iqnpfMdWE4T92H
hfs1jAuQvzVgVvnvhtVaxwzBNPc2v4PwRw2oKnSGEbSjt8oepN1ZJEugBswrxxydUpBG+lz3JMrB
3KUrzrwGSKmTbcwJszmkBM/pk2+nPJEdLBpYhuo+ugpVsKZ1JY20EYZH1ZH9R5jAC7bDSyqwhJ0X
rvfQ2yI/zIi6HalpCZzE2td1JCjpnqrouHFLVevucLfbbVtJ9JDS2wb37lFSnOCBOC7RrW02TLmM
s7K4rKopTqOVgQvyPXc7xV492bM3j91/2rG0ebiCAhPQ04B6eYWzrBo5z6swssxiUK+lqSh0Cml8
kxF/A6zpnviq8ePVh6TKA7tHD6pNsRkVAsfVMHSnd7TfKVkfkRkfkibPdtL+DMvC3ZoOCQjDst+n
gaqv5pgMtQmTiut9Fe9MxMr7H2BCGi6rkG6QGNEfg66Re8vR6yQXlbCIfXmxbxcFOPvoSxHW7WcM
l2udZAPz+T545kmWaXu2o0KFhE1dJBi5PqH11u9YCzrswGRmS5t0CPO1uw8F+oMfyEBYKRLipaT+
49WK/TFls2foAiyX0jQydjngnuWcwiyH6LroOC+bIW+nGIfQIFBS2Yr/YQRkDcAfo1C60x9ANNyd
t8krSecmeyRVMyga0dAz4gTkKODUR/lvTjd3K/u734WqZTldPrMd0Oto1Vt3RlweM+QBqSycgtz7
GdwHewcG5GNpRAem8mVBOMbPF4K9zsY1wBt3Y6KRnq00SYrkDzeQuILUvtPdIVFMxleLp4dnvMsz
FIgcChMfdM30hhglPEpQ7VdWI7IsM1RbcpSJ8tDvpr9PxpqCQ3lPkE2PjfaJ3kAIaRvoo3tBo0cx
Aqk+YJ0Yh4gxcO0TvNpXkQ/Onea4MyqfZVD4ZQNH8bS9ztyuXV25T6HlDgDvRFf2g9J3A7fyJMo/
2FkgtGvTVv0Gbx3B2YTegWC4zAvbjrvwLAk24vB+gAOLt+EFWCRQlaCGfg6pzUFnxHvEgL7cN6WZ
30nigg+8X36YSI0ANiHMMKEhwQVshLj3izNILGU+uAhaoP4fNY/T2xkR5KZ/HskndP66FOOtwqVj
ra7FOwEmx+6uJSeS1yymLGWJEY2sqrYDXZtQvgLxCb8IHg67EQHajuL7C5q+w3060vzpjsLHrFU9
IV2sCoFRIku9+Z57Tnf13oFiX+F/LHRHhvm5EizfuU2C1G8PBoBXPkLJbSoYqqcQznLH6sC1Y1jY
njTxKn+xLs0V1BzVbo/4pJKqm4PtLVKfz+LcrboSqWhclWsuPVYfJ/xOzy2XSazULZNDlevclGra
UjBsMok/qBAywakcf6FCtjlaCWFSgVU8WjlKwqLh/KlFQNgXgr2FYkSFEYR/Xoex5is7WirXz/aY
iwLKj9+WNMO4OOFJY+x46yK7pv2K/fxFexEgS3fIZvKyaNlOC/zbUnabKZkQcos6copAdnLicWBJ
nDOxWfLA/wRuTKvAtw5nq7ZnMfL5pNDcym296ELruHAzQ0QdqfkE+HKctIK4SVA971D1V6ELCofJ
HWN3kEsrkh1Zrq6yxu1K6UaQSHKaPG1Vildm02ZAESWwxRwk8gT1uethIKvsb0lfqEA3sV3VnE1V
0g8QWVX5BSDCQwmv0eqIBUUyCIX/GVuZtvXZNl/KUA+fSOLDMwnqz0LUcyEYkyHK/oNN4cXXmQYG
WUkXjyunVx+9q7UrW3b8Z24U13kQtijRQGBb31aMU1W2tVon4yKVRYZDiW561GMl40x7ySsccILs
06otyyXCOVacXs8n3aArW15Xyo5nBk+4jM6j15znddakvpAJZV5iqGh3ICG70NGtrY00Z56+vekX
1OrVD1/F+kieC/4juI/dPiVotlJm6jHYuFly6TVURStUgeCrz7xlpccQ47DYx2nDkMZSzHaXC9IV
LAby/z7cRiJItOS2lEESPHao3Cgw48qYgeYg8RGYGSux5+EFe4xH9abK+Pf0pmuAmPNM167vwcuA
1Nf9Gqxwd8dI30ypR2BXhKYMlGkiBz0/dFSaDC+vKFzV02iQ2sgTKzm/UwsH4+7pfEokemZL1Kou
o8mNvtAK2w4ntaSk+eUsDM92avZODm/A1MzfaYNNbIDNiIBTMZJ891m1Cw+RK+hnSyQTMz/ZfncE
4sdT5pI146wXByuHH+JcwS6vhZ6DLlF2tOfCMhwWChwpSLfolME6lJESyimetPK6K2DzcBd72b2w
KQwxOfZhQQOYJZJPQ63YrhiqW0F1ADPW31uHkAyL3ahPHTgCGRtP0c51xmfzXTPhiIsiU7aTZCH4
/BCqBcr+RXNyKAj1rSQrfsAw/kK+W95wBwJqD3hDV9vg0de5mnIWIaN3cdVVxOXkcmk0mZroIuWo
+u0b4o69igWFe0VuTPgK1Eu6lPbtnM0zgJNiAT0gTs9PvFsFa3DrC7zcLr8skqRr+mGjn/G5GPaA
xdGOIoCcfw+AyUrtKx7eNI+ks/a+3YNmg/ciLB0ejG1NMDDoBa6DIVdrwIFENHdZUja6uCDGAY55
u0iwGlrMO7Lw5rNWzg+tIyXEZBKVc33UopoSoS2/oj9Cj9fzopQH9canqMewXYSEYglzVIBCawFv
Qx15S9vgiVTvN1Fz5R2a0cL9Sa5vEoWSZ9VHg75zNQsX4R+ZGvGRammxDQ9RjSyt1p5y/GzufFYw
LLdnmpt8OuJtnNECudiha/tIyASnCB6dBXVAjY+I5KSb/L5pKLM7HAxMsQSxwUY0Qpy7IMRo1hrr
SsQv54oR6l881a8Q9+7Lako96vjzwkPnjRbph2fwZqcIXMc0mxcN6YVWS5e3UNHmukWwdI9/W8rO
3husepb0jdqGLlw557Glfpx+1Is3sM9Jzel0tbEt0mUXcuO4HHTOnk01qe5grHokhoNro4NuPxaH
OH+4WWLMfj7u4dYXB+sYgaNeXPRuQMVor17EPAmxXJIaL5mkdjM0AXNm6TZK0exc1yiB/PM3h+9w
XAAftyjiFFEKKnTRihQOybSdhAfkj9Pejf2euAW1U8drT0xmcNFDFfTEW1VdKMPQMBKdhBcRGuRu
7SJciY88+gQf4plfZO0/UhcKFwnvaK6x8fKeLKCn17X5hlH5E5deFFNbcpAe4bE1ACp072ooLDgE
ksgg59k0Xh7i66Hg2fkaZu8dPMGGJN4O2G1D4A+GjIMctmhCfXkMwgqQkyR2mZWCpIDP/uLl/kWy
FWC8Xvwl1LOiQQ+uma50m2gP3B5CieYopis/VsU60pFbWMWyIQz/XKvRLVPwf9aDbhrME1kvTp4f
75w3yGF4/Q3AYQxYKGNpocd39i3DmbjMuKdYxpgOLsMAsifqMPY2xxtVEmOP6OOUXpp2LcVSBfLH
iJF012gmsy64aIvr4V95Fm4Av25h+EdhAgwi83U2hvh0jQwhxM2Pxt4EvlIwR4s3wK7uGSIka0ss
2eGuczAmoxpaFa51JYdYP0kqTJ8shayz+822+P5DTyZqZZW858BSenOEJgxrp832qqGGM7BT7jWY
aqo2v5+V19Kvae4K7M2kZUEmC5xhcOoydn8kSCEZKDXvft0kg8nNcNQsrAji/qNJJr1yMik2SsS8
oCY36mW5hLTFpURatwHuRaOstEofdEQ5HU8LysFzfsV2uIBgUVZZnKu5IKmD+z71ib6W/Zge7sne
q1f+HOzoFmcfFYl1eM7mGUwDRrTSNVqXgsGxAhYo999WI2tUywaCxS7g6nJrW7wpvZYBxUhseC9g
5LxH87RsrsmbYrtDrny+C5mpulMLCX8PpyzUL4wyvHHW71skM+irCGwL+QdidwdazGcuzXRqa3uP
euRuvk3r+mtL+9T0gk0xLzt9dsXuuaLfDsvoL2iwqnq3zhEuWcVT/lbXpX0JNXn0TPUHpRwMmV1I
6tWYbjloL96FlvG7DmdqrwjJbjmNY3efks1fPugBy2PvKQe0eMDxuEHKslDJ5snIjozrmIMSLKAH
T9ryS68FtgrG7LEsVGvyM1ZgTRuDKbcNNW30SrIpzcNX4HLslaAFEBS6HWdXMNpPNRnifGPIpftW
FOTbnPOmgCJyILmxC83EROmQcA3a2WuQ+HANQfRBBIKO2zIaPJeSXppMEdB0Nykh1qDqpu87MgOw
/GvSt+5aUYri7aySSN5APvaQCL17NwlskUaUxEb0HHenrYf77EnA3/kX01pe77Z8HFPxXbcCyiN2
GWjhm6xExXzTx8VkVFtv38HEEHzeDP8m0S7t1pJvqO0hG0jvKokmT5Lzb6Isr455H2ULIgha3VKF
nl3leLtzzteCnK4kOctn1/jPLVjPAvAbPUuVWVBshLw5JXUPD9L+MP3PvVQtxOoQYKsqd0HSVkaV
8YhEtC3xs067flJLgX7spw9d4rRqYEiLD54TIsB9e4HMkNqdNgF4+xyVnPoU2XItMAW9bKFefW22
UMG5GB4TWyKZl4pyNedSqzqtbUIx3X/XRv8dsn8js/cNrz+jdgoKhl83U7ArR0faJ0w6rLNXXRiV
VQ3qYqeZuwbbL0nLRQ3af7AU/DFAjpWpw3XtZGhWXWRXEMFr8kY3gbTVcTB5H5vUXaxvdlxk685g
d3HR9inaT2o36UkzpN5h0QMNSiMJSmO1AzEK7es7ZJi4qI3fE0ae/ntkGIElQWAVOznOmpASq65r
fpozyQZrlG14i+ax0K+0A14oZ6M0jPgW1wxzb2+Qs14o82yEi/J3J+G/L0AS5zpjJYTLpw1QoL5n
aHVBVDOVb+JWfsA8BydsCTyEMMObcsNhESRt9ka6B+uq42DVB7H7JKCcETZd3WLWXL+IKLnL5qh0
eKfCZWbtLkuQqQBuyQJq68ZjBJc2RgbT5PILevuI8r8MCKdvYRezTFSIEc/2xQysK55VQqGB2I5r
Gp9RLegU1bq9C9lM2Mh9ih67R3TQaq9hmE6MOdK9fpc1x+JPEDEaxB393rGuNu7RUGuxKf0yGYut
Z8NyBdGYDlscwiGKi5jmU5vfnvOiDQ+hOXT95M8d1sY/SKjW1NFo9psVQul4ro+Hr755ySjGV/fl
VGijbqKAzj4FJ7iE1eCGqWvZ8h934NL599pQdzYAgTXJIMxGk/gge+O9A0ZP2QzWOtMjVAo5M5Sf
uzibH4smOoJsyy0Vg5xLJKw+GndUZaqeNRHIl+0i7OA1TUnQRyWKQxizc7sMO1NPbvo+JW8viEkK
YSrsY/f22hppJlY0VIET423vTwa5GP9T/8oHy3rpcWGLcwKE6Edh8rZFXZBwIfdZ5GY9B84v3Bvx
cAZCdjiUun4HY5HU22ROwsDOoxqgyk7ba9mpzOCoS7CmyQjZwx2bJz2BPTM2xHtIj9gx+lkdaRDR
vCZLi4VsgizyTn3V/28yPRU7e7QwRLtKLiF8NrjJqQ/Tlxqy/5X/dxf5P62IQH2Toj+UecAoO5Nc
EWRdy43LhGbH/9f9IVPhFc7CdSMvLuWP9hgonZydwzXgtHgIyQhIPA79BAJMS/LrduIvKuJmdJU5
jjxJ+y0UMaVFUHbjqbs/gP2tJoZIeFJB9ehqmlneCKlTUeJfnoDbDhSTOfzIaiTT+5Zp+0qVZNBx
SrRk68SvnQEj5wpJSCg/mNqN1xckrtNxxQWSzSlnZV3TPPrRqohaUb7Kd8T2HoJYHePS/S1sufVk
yA9RHk68y2J8VjH2ye8nZ/IQ6GlFV8nWWBSvjlkI/m5/kmj8GwM9qKTzn9a8vWe6zhv9jevTutct
FsF+5+dehCEO2r1Mpzm6wAuJgy72KoPDCykB/jKpYW1e4S5sFBM8H2blsTO9UK+xcdBACta1rG0R
Cr8M6D0c9TiGzdCkUJ8IkxDWqNmDJJuCMcY/FM7zrXgm51DkXn3Aen3inwS404hrjvuQ0KOxKnwf
hti2tHw2+k1/YUVoCtFIyWO/wvISxwrOWPTCuMfwzBiYWdbS50g2FavmYnkGazjjEt/XLxDft1Ok
VfPgsJeXZXfsSm/feUWclEq6pRCdfOjYafys6QtONwRfIkgEkkpqo9+OtCjpwC0eoyU3HEE8UlaD
o7vr0Pn9vw7FMMrsftkA1JQKuOFjjFroz1xQ7F7YmSrk109unbFq3kWiYzrr/2Hh3187xQG/LjFT
xgA9lY4+7AMXW0zvMoB0cG1BQwvze0ZxoMQentLm8AV7DQ1ABkcq20d7vGnxWnZHacVJC1JHYfkU
sr7reSZYRGvstFJ25/TlX8ZIyfz2oxc0mxNFJYhi9OC4wCd49etHqD3DQmNxIe2SY7J950si6MAi
mKx8nzD+sRIpaN8Yj/zsRw4pRxisdmXQzXZh3pdtOlC/0ZVRVTbXrewqyHLMS3vmqpeJ+E+Mv39J
CtX7MO4pzv/lrf1OMZIdHAuexW2cLqOYIZtBL5bIMR9HfFSRS+W7MlYSorRHvukJrv/wxzh1P0SY
FWPtDQPWJW5tMCuI7yg23CNcP2JoHj6LZ8tp9TIchmO2f+wptcnQs9nThZNqwpyTKNUP9Pp76ZGe
RHY5n9VJb5WmycASbkDCFoBQ6fQ/ob7NWD40YLI5qzWTXj49TE1f1MLHRt2tmQYvtj23V5uu+pu/
BHCmr5RZYZb6c7ApHBILmwkPXbkSqVCkzvs+J22ltUjPBjH0pCFQL95vxcDPGbtSrzkO2HWae1Wm
ZsIqV59DAQH28SBqExfpWEheq87s0yPRaGogmxgeOKSFoQuCLkXpVxvC1TXv/3ZMoBvnIW1VygdE
9FwgmLbEtFavnq8oCsQoH4YsJbTL2g7nbzGFZ599thsZ8DS98kudsogpK6Ud0mzHm+DZLgzCwh/5
jXZ1Oje2X5v2ePZ9/zthzLOJCAde1C2GD6iTIt+LnSNQe0ttYfc5JKRVmvYX72IP45Or2qiXgLDw
opQEhipczjspCKvIWaYMT9HZJjfFSQOeBxXyTv4L5SzxAeVt1X9f0LXYsusXPobhR+1qouZnBlVY
xeSfzVhKc7dc5pfV8b/BluXXBsFKjTAujuQ1qnHUS4vqtR0hnyqOhb0zEX+J9D5YC8oeHsjsVj6u
ROOrdk9DUeY8khC/L92P6GszWFsUHhdl0nvIDSRAhBBZFuHQSHhLpjeoFP/leAo77BhRXf3eeCzg
mVWmVb3KU8/Ja5+2wB5l3IIvkXpAGYmzJo0Muxnkpu6M//OzRGp1WMRBmfgxS8s0u4Rs+J8ZjCBj
gtNh+IbcwXnqXr5EWOhcv+xaDIjpr4EaeqnAs21oSnV8VpAdl+YfOGTCjYsPK10o9x1bnoNaq7wP
PYVo1lTT/ZMWhmbn1jD2R/ZSiG6Tv0OH6jMI9aIT5TzOInB+4Hsce3NGetit/t8SMGbB9o6s7CkG
0mHm+alUbyXSABfxisvozVgOgCzvc7CXjyY/QgE2P135iabb+UV5eImr8gGpu0acjtFbErMG+STa
tRJY8useDDvhqZCcBmBKwvHiLH9Dle7kkFxXavy87JKAJazdhnih1Z9K1qkTKAygAL/14mIRYR4a
AoHZSbC7pcxRbpMDsdqGBfpHyhkGYuEA0poP9KR3nWCiL1FxEGf0msAxeon+RTvzDcfxpt1kBPDJ
go9Hzs748/R02l7hl4O5ySAdIrX/O+66lTIJBU2eVMKkR6hs+a2nlTqCTAk1usz/buQ8k+I2Csmy
Fs/XLxt1ZwaDB+trJgGZUL8cFU2eS8prFW6AN3LUpV7C9r05+YwgCjTQ4X/MBUagXIi6bIS/dldj
AkYz1n60LBcx+v3EtyPjAENz2tOqLxpRvG6JaBm+AN3SBFlT7NnCiLV8S6eVfBDWXoUeWP+doDVR
HZ+3ukV4m/gmwLRIC4rsSiEYnvVXpE94uRS1KdlsoXdcsPsYcmq2nRiAXv3tldi/YF0bj7PedfM5
LgzO1DhSx03Xg/AmgT+qSxaMv5xat7tsZsF/5yMTGGwyHkxqlYPq5pHUm7Xa6tFnjqCkRXlolo1L
TOJ+8MJponLND9c0KFv0v3EiGznSo2qx8mfEmTfmPjqfcO3gSEqCeuNZ3JD/3cXTLoQj7+Jq11RU
DhgzLbzGo+uFPGPpA7s8bx84oXbebmAgeOR3tLlOIbi45XxvZWLkZ/92Mbh2WlWlEKbZZpcpaSbf
qZ0xR2iromqXDkq/DR667TkoiQIV1Tw/7gBHdweETvNgTkAmkKzqzfxNyu97ijOVXmEhnyWd3iPV
bEe6i99zrTakTqEeiAZ6not90nEgHtobUzwwYHqFEpM4vvTEvBHszCiLyA9I9gTE+ZRHOvU9hLZC
il/IB/ZxYY4wSWaVjmNhTazCJ4qp7gtSOfi2j/Ko25tbmmOMzv2KhB/Mb2aI4OE0wA+EMGC3zve0
bGiiPtecJpvUaAJRESuhjf3qGGFxSEJj5Hc8+9A/vceFvRolCsyuhhYXmGNcGbuzZlB4IUXlyXk8
Gfw+1L1ucOFOU28lQ6rFHos1CzWYyjtAuax649HrtKT3Z5e+B1lZn08xKS+dWpr/aJxqfhmMbVZL
7Dj3zM+DvyWkJHDFdnXcTZZ3noeldczQ/c53WYle3d9/mMFej3/rgvvrl3uE8xxaC6z5Kqv+PlAt
JNoY2EZJhF6DKYy6N13om7I2D/ddnKp99CLtMbcxJtqHehDiQplp3qQ/dA64OKXySMpV4x8VTNam
17ZTVtPVXO2YxC0G+kg55rTRtyHPZUfFofrwVbmNd2qtZSBeIU4hiuUsIOCqT38U/pWa0c36puYL
xe72bz47QtjcCDnWwzOx+BUeGx+AVy6m9+YJPiSRSpgyO3SU1IxABNlyccFstCGt517SOOjU4zBx
F7bqAaruuyMe8pK0eim1eOGcElNA61H/qa0cpkXBATyJXb7b06Ed5rxHvBWuXGjxz81iiCCzSpjH
61WYXA0bGoX3eQzzquB0gLSP7nOoZn7REg/fGqDeGSzlu8jNppzXAe7aXHCf4ZrpgbMpGx9DAnVd
WjvUCsQSotbLIXLt8sCUFW1xEHFIOeofFwqRLWJtK0TGLX0LmjTiZPpvInfXBzN+En2EkBrofrcm
E6AFJU2kATQvafCjlt/DdIsihFpfFQ88Nxw511nfCoksBDavrv0x3Mn9qfrbo1IrP3zmnHn27dRn
k6/ixj/IkCJBYIXshq9keg/uXHchhXWFM4CQofUZuDUCWwyLmKoqs3DuBA+T6xuUDy2kYFMalH4+
VOhurOwC0d8OfKL2/96x/wHr4YKU90aYJK1VFruAW7zdw2O3W7OS1hn0IQuuSP8Y79qisFmNN4na
di49cHbl94PuWdIeUEijfjhFKEaA7TMue88AeSVsirowp6Lp+eq1ktGIe+mXC6UwjX5a9//fY0Rc
5rz+/9IyQGbmte+NDXxL4w+vtWAv9A6g6Ud+v3zfNQhm095iSetdzux4HMtqtr3jkvVpz7IPl78D
jOUWdOZ86Pf9GaMMQTxxIoU5knEYXUrpPYRdaSsZoI5CtFvgzwIaDHokh9i3Sff7DiNKaq/BYDhn
lcMCZxbPKFDYAU+IV21AKVJkR1eE1vwc1hVlNaUtVehsDEcW7wwT18Fj7KxVJ+3KI/cdQ/DFeaS5
YorItqYmn5udXHDNJhTBd5Jc4nIVVExYWISQMy71Eljpa8k9+uS7mV84tBxX4SrMrf8oHj++9Pwq
pcKFDG61y6S9UkPZ5sDv19RxpkZGDeB+yf9XQqgkLZL9HD4Xwn6tlpPykaCpljPmmPeK2c2bPvxb
QdAG6LefO8qLjxGlor81sAQMN0qu8kML+dCmLMcjF1QOOYDXCiSckhNBi8XSGBmRrlyJ9wti3usv
osGO0G/LCyFqj9RUPhHwQVYP84ZxINGmQGZRS8n1RvzL1H18kUSZBhkz0idnArxyH9XDQYMrl7m7
YaXJAGRJzqDov8dtcbwA/Zgf4XbdgcdG4jZCLlp/B8etIdFEcUFodDXbv39SLkRxt/+dFWNJbsXu
+CL9GawDAAxE8GZxZ+b4mO+xL2mNUhzVD7SJPILPzD8L7hVj0ELCOpRPfPVCJar10R1NUw5P2FmW
AcDAsJqBIA8bf2V4ck68QB6ZxQgoY7Fo8KTATGeHuPjJVs8wCRpaXBqNogyWYe1LrVLHICADExzs
H+cqiFYCe1QbUZ6rMTgqkM7sfB7fW5yOJuq4UPiKZg9t3VyzebAslBGlHJHIBlw8aHQZfhj+GTDd
AvlIXxxEcpzcXf7Ed9SvtIj5LafAHAoD91JJ8e78bK5hbfcZ3GZaSSJM+xeRa3EkpalTvOgW+duF
UfNm0UFuCsTuLPzMfKOTS63VYQnHDZ7V11CTKtmogqsypdxLGolWmOxvzeGH9koSWzHdBnclX/M+
Zru5Mfq2FTOaQrq8fgDovKn2Jamzftq+icZwFRHSGeORB0CV6quQXoaRfcCsBrPhKBDJaXBb2a+1
21dmbIdJZ9u+gbwI78JfjcPtdsX4FP2v1u3OIB6Uq7V0akKKpG47iEFgx4gl3JCk8YOUPvqi1Rww
+x2zrSfjzrmof9kDtMszw30aJdLfZF+/Sy2CBgMQGQw22snAn78sRYix4df4u2zwWXbNGEf8dnoT
lQdrzDYt5iqVY96u2bGoNwcBLQ9CsmNWTp1XpNZofDlGTQPl0pKKXoLYx141y2Yvjgr2jGd5LfNa
q+NYcSv4DgA+8xaX5XrFzky63ggCXVJuZw4XqLhFyLdLYt7T8gyEkhfZGrIWAyzjYZ6RNRNcnEz9
DKOZaveg+dSASBaCGB2zgM5pWViWh/tlm5QgZW0dSB9GcZ45h14CHtDbeA2pxCFiuFqKdhClxNNi
JGZkzKBCwCVlatiZuPOJmgHLQy5UuCmkD9A0tAdd8YqUnwfXiZ2cvHAq8fc1AdxgZZHa3ScjPtH5
xeeK/gxOHLRTsd3/UB3yFO9AK+l93WZZalHGF3fn5TsF/whAXe5G738KNjjSxqqEKaoWx6ppVXvq
dT5V8xD0jVj6tsoD7Ee23OAbfcDR/Z8mPhdL5alH2UZpi6RXuka7OtQiSKcDGZsjpwo8N7Y7xOwv
P8y881z1D4EPtTd6UYrAYcxp8CtBBTrBsfKChpTy580pJmaWXut7GCYPlCztEMhAbQtEJGb21p44
lPYZH4RPXII11197aAfBpS3TKnzOc9Duh1UZmPRgvmcP96eCBwxnRc40HEAWfH05XeC2VoTfX6lV
6H6+wiCo3sWWkeZzqSPubjSsIxE2eto9ZlytFcP4XKunDZoyrzJWLLRHoH7UlueX0nLCkNyqh6XC
Cta1JRdkfEiudx8RkAsynQCMXnB+USDjIJJAcdO0jRT3z0iH1l7gNXpGeeaMPjmS/1PpA5+Q933R
0l/cucOFVvM0p+YR2yfOG6YgZjYs2YUjMdJsgFTXksT642sfD1txcu+LE8Ou6HeAPjsTa7ige6LF
hzfGJ6VD99dwMoQaNHYJ4tcGmuTdzD/AmCcqH4MCTPzIAKS3/sLdiLGJw2szm6reAkZSbFAAViI1
OGp8uFVS5+hrIPUytSXJPf4LfNWh0fVtOQCCVPlxADqYmYap2ye2TouggDsIGu8j6eyhDlzBPMys
H2txcXK3CBjO9SpKINUIKzRV3ZOcCJqAfonq9kL6QlBzGT6VDmTYwjmX3YPi/4rPxRbLPba+k1Nv
AjLykwBIN5xNZIDGick8Z2OgAHS2VHFa1DKOAIlEM5IQCRfYESuYmnt85hk4Q4vcsZXYbrbUS9Al
85FhcAiW7QFOG49eGT0zsnyu3kX96jF+xeJWFK8r340xHCfz7AdcqmkN+HmKI83M/rR4YCRrGc6K
QYfWx4ALbgLiJ2qyjEWHOt3fDno1PfrjjG/IRoICopRVbe9y3NiYOVEl6w3GXq0JbC93aiBZLVIF
3F7wR/goO6mNOeAta31w5bGAP7BXOp/RoE+7IgIy1fSpkfF0EFknstjSDdHWkZW5f08v3L5Rc6Sb
mI5lK4xRulQtaXEJQGg40s+F/nmIJ45/+Rq+ri6NoRGSU3AtadksZ7nFvBJZoRCno1VrLsQKuP06
lXIaPifgPRKV9qOzMr1hBNrX7FiXWarfwlpPxINzaHq9a3znjY84OM7Z3bZwGdeNI157LxZzTIoj
lcWBkZQgCEyDbf44c7wAkg6Zq9XLeN3hzUwpWbgQWAeT/rXhHRoANBOK0lldFCwNy7ACOZ/vDN9J
pzysqTOOuPOiqiX6M2jB30q26eOXa3XFeone9tTF5gBPTQ5Ev3yQoVIRSJ7rXf/IN/VtDGEgFTJW
mAWWznUbkhKHIM4yCHWUsdqPc6rf16hPUfYA3KvCOkE8fkKzwGql9oYkJC/3vIH559vM646G+TlQ
PgojFJ9oSL0tPtKhHWQO/MXNDsOR9RRYspHylcV1mADG49lMC1dSE9/UVZ/oXozwpvPzPyYCQhvU
3X0zngo9TPcyKgfRP3xuW/U3Nzq4DWmAomPqH0tUqtx26Wjleb98CFBHlypuX8SnjEQYGw+Es/Gf
k/t3wHbqG8KoUgs98zqEhPKoljQ+NGjcVMCqeN/s8oLnFfbp6T70lPL4/DizPDoD9o6xxMlKVVg/
MhJYAXpElykBUsPTrXXr13hxX/xKSLOWcDdYEtSRrBUu3MVn0bhWK81G/8kII8PyRw7euIpA5VGB
FLZR/65eCDW1ReUma5OGoqdUYdlrH14zefsCiFJ0stOYvJeQU8x62AzfIzaNSIyh+zo3SUPFGzZN
B9ZSK0yErrvMkt+OE6red++DQ+yIiSrS8YQwSIDKer1oeu4tE5CQJZgPBKjQTQTxgsKOkbvJrXs6
nY37FZbKDJC41Lcv5wjxKu9kgllpXQgh68ejhQyJ5SyIH1syfVv2lbWMCK0G7v2zPm9hBQJmbYws
EsdkneENnSdMGJ9r63EFmt5gdKaROgnP/CbQSkFdZ2z2WqsB2ysvdDxhy6BIFCIT0g2mEQAJNoy+
n6nZwTwc1QRm1F41+N1gQM1orWXLxyTJnlY6fau/Pp2KdU+hNjOzmt/+aLE+rmSmJf4nZxETiK6n
SX0OSdNJEwKYQY8nSoiyEp7VQE+K5BCUdS8weyJEaT11G7CLGUbzEi/XlIP3V6+p5/2W+bvX+8Pp
2BVMahj6TIOjKYv4VjgeF9TX1nDO7EXtrdQVm1sBq0Tcateex9x24IStcCREzr61CDd5ZhqAOULd
ihso+nAPiN25cDkXbDdJ89u+DhhIoeO+fYiUhc9zWQGQJertWjc6cIdGRrb4X5VIDS76R5YrfPFc
R38rSuK8Nfl/FABu/Yg24WaK4CmDZTnJvsjuAgoDJtDDS+kNSItT0/07rPf7tupR7oEbStlX31Ju
1p5tO+NSOTO6kwvAR74BGRCUIJJtkkNUN3EUr4nCBZt/lsnALZ0ARF+PjllCbWvZKALw3qQrNWLK
yvuXeuLQpHUkwm+46BV1vFvj48PoF6U/PLv2B33Phxz0KogQCIr0MMIY6cMoyno6LS9gg4SlU7fi
2s7Ym9bDaeaXhmnamV6rbZ2Sz1pldJ/DhNKiMtxRY7nAzMmqhQ+EGT3tRG1+hMVWCaYPgElRhiV9
fcVkYvgMyaF3m4lghoqSlgL5LewKSRijlwTCGbE0yTKDjpNVFgCAIeTOeXmucBks8fMD2AOrl3dX
ZqUB27R/TTqVKFvmyazhFt/1cYGlChMZmwfwO1jRkj3erTgRz9mEhXwqECJz1xY33Jwg/opi7PMO
5w9FYog14aZWr+/s3pAOEhfNYymDmSuiCghveYWwrJb2QNkX689VZYqUoHLOmYHMqIxzo5oj694r
cTryal5W9YySNCet1F9caSgkMhp3chFc2tWCr4wsAqoLbYfFQp1BfwosZ2WLOAtwpzkw0cjsSb8V
QOVIo7QrQSQa+fDEMiJ4nZBcfJ2JSaJliCzMt1CuP/gBQA+3vgR7hS0CV01LF+ATM23msrAmAl7B
uNi7vUIAEezaRQjXHKD2qNfna7fKOePpXMF54Mb2lHG4rlncXnoBzKXrGBrb0xPHj2KBcTFyrh4z
NHbibe4LUeAjEa7lhSkh4ya663PVgvv0O73qK0+FlwPvD1V4bKUnO8TynOOqbolj7a1ocJX+EFpw
n+lfvhKtEkMb/WBJhmbxT5prvmVp6ucuyP/Gso8zJWdAV8uRrneu6CyTQ2hFpSTkiE19zz+S1V9B
Qwu4+XtJiHESkPV0gAQrF51Tc/otjOlwkgyUJBblt6tPoM/6rOijf8UeTgXhIS5pUvkeHVX8CuPz
hx3ZwOyEeA0tRFjhqX0lBNipOtlI28LjU5MuWEudDUBirdbJPPtxf54p8M+7LyldicCK5opdAMCk
S9QdgfyrCfDAsUTk3ErVjDojGLPruH13p32/8Bft3BW19NcyH7AKLP8wSPZsOgFDdThyMnlFhbDh
4YZga/JQdsF+goCYwdpRjn9LN116Y5xk48iHMB/YVCi7s+FNa7zmnVd14VWkUimRo0DlAfyF/Spf
pKovBBJME5nzfl9ziBanhEIh1IgTR2dN7rkcnMNmIVnT1w5xI3yNY5YFwYcgbZWzRs9ZNQOCGJel
VRdf3s5B1+RiRrfD3Etzl/truhviFq+FNccpRDEn17mM8K0NbxpKZLhYKG7BkpMjbpToZ8+37vkW
EupUjjMbZm3rYZYoINfBNO5I0Kr+idPuW9yWq7BqhIQD5CbvdwF2F5awOOBNnyjA9peP20iE0jZk
/Fbklfnwb0NhDHFB1PKRk11hxYaphWAoNrSgxQnpIscbl2IoOAhMm2R0NplTtC+t8uReop2HHdGU
z5dcXbSfWfrBnl2NatWh00uQ6NXIZlkPTVGfBdSUWOsyNsiCrvfHljEDr0i9IPkkFMVTJys+ll6I
KStuwyCQ4LND9Ycc+7cNuhky4Illf/B6VZCVYVUK1W3shruRJUbbQQcjXusD3RxY9SF63Tx4hiNk
C8CzmZGHoCrS3B3HP0u87s5Zc8dqGxgTHnBUJXMEMP3pUSZAoH0mDtYRIIMXuO3C1BCxWgOgxH+W
GS+1V9Oqz21Sihyk+jFUizOQtmJHBqhr9UreAuPtgcpTrfGaJWWCtsr2XyBs+uDMl1zdhmZ0jEss
CQLQi8RI15+tnbzanaj+QoHEfD47P+VC5PbQXQ4YWgXlLbQWCqhHMPuq9X/s2roIbAapO2TldBD7
KrzWUnzoXMcRXYTrGsE/PuJdkUyxwZOgPJwPay1eORzPE31W2mEmDBU1VaPgHI/jyrk42zZBpp9W
YBDBhSkKI7a5amGhzAgz1oC1NLA6/RUVJHAIE/7RCch1JfAC800nVRETG4Edb1nRkk+uLUs2aP51
zQwDQzJDiDV0YrwYBU/EcFZS8lSKPZ4OCyMWB578SO9Cgwq25R1DzbBaTVCPp/5W/tcUO6TvG/ye
0kbOpL4YtuY2mxCyYVQ9vW3SL0wu1UWipqv/SWK/7QEev8a2CB4BRLgqLNF2l6e5sTp2dy64Qmd+
eDSyqyN1OXZQzgcktY7EHKv6ZQnyJY6ps3pvI9HpwNifG0doqKKU7yzMe6RO2CIyBMuS+p6Hn8td
Xn+Iy+jtjacgo/vRk7GV5LKQqjwPUTyoRjFo1HM1n2BdbeFsl2yegF/epQ2BCOzrBPJrtNCrlqOu
ALAPlZn143sXptKEOsTvBXP02RggAxJs/0Ah5w3fPpVL0SmXmJggIrnDlMg+KCL2fhrWTGx7YrRm
01HlsuGqs6c0t+JzUjk4flE27W3v/Yp/ElC0OYSB3+JC7oW+TLA0lGwbJI/Of0bJI0VvZEkiaiXv
UOgPo68C9l7YogkEbr6Hubd+YXmXIaiKQ3y3cccyOUX2ZNEexqnI1zGMWge2V8Td2MKXLwwcP+ou
IZlsRCU90vKD4r3t7+E4Is+QS7YHkepMZBjfEVPy22/ErTxlG556TGP4rIUWUnHtTsLLE4sNozdY
VcnArIdvt2C+EeJWbQMdYUFXeQyvVog7/ku2d5jQ40lqIVAj+9GNRldc6GzjM+d4ygyyoIveHgu8
T+R33GlbLnp681kUMXXLarbKp3dHlrY3yD5eSaUtVtmLCyZpUrPNg7lnukwmxnQ8gs4LtxU4wfhQ
+5PsZfh1gY1b3VJbYRk05NmavFiGzKMxtw+Odiz1NvGqbi20Xo+EiALhklncMiHkuKsmXNemr+Yj
j0+53JesmrqUnWciz0TgHPQ5G9PwwZfKGF3V2qOGOx0wOBgMdlCxk7VmVcqadO3vVJulSCpcLpDD
sbtB0BWcJOcH2O7xnY21q9RDCeLxvsxs2rzFpe0icIdH26wfJHX1+RWPbTimU4N6q9HAuDw5Q6VP
HKty7jyt7UyutEYjmrRnWirflgyp9rN2GAeGMnQq5vbV73TEqi9G7WoZ378Vx0Onpl/ZHi3za7WA
yijmL7RQ2RRhhY1v50drDvVD3QByHa5SO2O0Kse8BVLdwEn1QT14T25enzbU13t8LKRJBoqHpZiq
WKXJIl76LOXub9oWvuv+VPeVVmXYCLUFfWDxffLRQmGeVZdoyxMsNXUD/Xu5mnekdqP1XZfEhVDc
6Yg/6RE+xRIlbZRmKj33PScY0f8a3E3t/VD7fNRbSeosqM3RHX94n13M4PYyzX2waFCPOmFO1ZIG
PiSO6BNKM74f2G+E9c33CcvFR6cnHgQzk1jTiCQCpBrDBpjjj7PxLP540q3b6R4lcgV9rz+STBQc
hgJwlKVLFEL2qBugZr7ebo9YEMvVb4ToYc4wsrbOt6nR6bBz3joG7hGMEZsMH17ajey8fHGgaYeX
6oQe0LzAL7faSDyMTlQPCq8C8wpSmyVAl6Jx6SV5Y2kPxxowqLUWEhHxFbpxOFA5Rw3wXdMsQ/ZN
YtQ1AqxvzRRV9iKJf/z/ExKeyKJgQkbhxJRfFoK52Pk89B4FPy9ffT6+i43BMTvtQqPFUSdZNqKK
eXF5rktelb5dcBJ8LhlcBH4vOi1nh26n4+ZgfzKnYtupaEFb1DZwSIfxtmRiXpXyzf5zX/zj7hml
zczmAu2toXr/Cq1UG23XPQsx7u8+tKlq6STuK/ejl6nnZEpm0A3Fu34VLGfimj3/taURyR93nFsV
bmdNynJnPrs/5QD2M/MpqOaTEhEFOt9wAQQNh7Q/gHozyzZuxNweexIwh+GERw1iOtNVFKVMRHEV
Fy1VXqmSNX5gQn432mcu60/DFX6mjhGAlca8uaDbLRbv6fWGIbey0EvaQkqZxC59bN/684mZWQkR
J9dT2Rg98rQYo+oTwQ9/G3eS3MLHYlfLAprdf6HjcSZ86nDt6DYUy8fFwwqJ0o/nLO8Pz58vti9B
S2Ds5m0Zxck2y6kkFdtTL1HoQcA4dkwfwx8deey4ex6ueb4WhxJarJT1VO8H0CPeZc9IWMmMcfWq
s3A0liQDJ4ucOR0PjZexrJ4ZxSHutje/47FmnrEqMIsFKOrZ/H8Jxwy1lZNke1xkGaIgU4z/PgVu
RjhSOzEv8fRxJKZWaffujt3mNIh6m+tsRmbEXcgTXgCnaLXvToCxil+hn7e/v4x+b0YfIPweSkSi
hEYFs5x79bMtz8+8ZaiFWy9i8kez2vuO2xXDGefIL9Wg5XgS6UythWbWAGDxLSjrJPo5MsFUWSl7
lO76QiIRBfJ7ttj0bioMHT1OgfCl+0UMzUn7TkUr2QJXoPXFNBE/LWnv/P25DSOiJOlMEqPdRtHL
s5xLGTPIFOQJfYENuk7Xvhn1XrUPmTJBSMy9opo41nGhnmZLg5ZuL7fu9AvztgwWCEiY6iGJdmv+
5ihAN4JZFdobMQUnfcJJ5X+C3/03EtNZCG/MFWoP1oBuw7ZO4mYVgcHHmRKLswD+k5k6n6K++FKP
vZkaEHdwGKGevvjR1lVHiP8f6qvypYTncu4bRjjdcowAS7G2r7HZ2fkPc5CN4xcu7/XDBx9K/R2c
9L16Ir+aSGuBHpB5SmcUNLk6pGbcF9m+g9LRAPUlLv3X1D/j5Tb3HuifXRG1hRG93IPI4ymIytdk
ch445ScxDh1Cj7PQZNzok7LI/LRvfzLvC/6JI/DQDORInVRxvo6t5cm/jodOoVA4Vnlfmk0OeDMS
9PhgAq4tyGf6j4tYV0fOVLv3kQ1bJHhKhAYLBHkrCUxNbL1FAxzKPSFr21YbINRRIBOPdWaDawaJ
d2OrE1NNpN+jLJElBg2ywbVPBdUeZYOk5surQZM70/i+iWHHy475P5OFLdu/dnjUiQKl3d7EqjZs
kweEQ53lwXQx/6MeA2r1H0LxmuAAcO69MUfqW3J0v5IfwE5oIbtkAS7m8DQd0KcJVvMOPqSyB67F
+G0cFRSzYA61oHZcTAzMLnZ6llqyofxwnnj943mfRYa2r0RohpU2fvBrzu9obTiqe1PBhSM/itvW
H+fsaRpLnd7hRkrDInEI3gUpRif3NeIDEuEuuobAoXZpjHegNPUCptF48Zs8UtHz677x8OFBUyOH
ZV6bTBDbAqTifthyBhx4HOAbPAD18s9OiG45o88f3fRdwu/6tRzSDfUc7fXtb2LxaPY1sYa4F+yX
jG94ZjlvZvmCC+/uZ0F6sv2gW+k14nBb36dzVIWoHT5uSdxJzUcfvyHirKqR+mTXupxaSD87PbE/
38lPp/XMC4mkICdw/n/S2G4BbaZDFKzOvTSVRa/RdrSKEVkQGGPGsFgduEVjwJFjhFNfd7OzYzoL
7ToPysBPnq+V5vYoBTUL9oCeVtefzmm0/svV30dv9WChrV67cLycTiOw4DfkroOJO4lAiiOPGf7M
4ODuu0s26BxMSkXXxXKaJf8x5VYAKZMCCfkbGkHAJG6PWCJ8PAXXmNpUwq7Mw7AAxQ/OeURlEzh/
kDGs3RhQlwhNgAdxP2ByjLAyw9W1Vcj4Lc685lpOVE9QB57BDXxvUilRaC3XINKrO7WxhY/hlRe8
TJjw6zVlcztImL/c76LoCgHDsgn3w/OpeSszSOw4XoQOR3yJmTNN881JRBT8hac023DXJix9HexD
GjZ4WLEgz1yTgQY5/SFox+VYf0rB7/wihby1P3jaMeRxEFq09Km5j0vREnp09DNQ+wWtrWR9MZAg
RykgxY2VAUQmOeTXaNlScGc1pFd9XkNIBVLciKtqnfP6ZD50V6MBvvfYISUh8axLXhOuy1xPT8Bv
U8E59aGXBk83J1BhpGMXY7bu5jhuu7chinm194YWdzsAh1II+0VIpM5YdkQxhJJiw4vIuGirN8cx
W/q6kzjv+9XIrkay7TcOWrKsdH0DJSDIL3tjOU9maNYnBu3dVXvUghltPXHtsbp9FvfxH6EFiSMs
8z+DEj8EPQZKdY2UeN1nWwkYyjIoClgptQxLaK9pT8mUfQcMjJQCkwLgkRN5f0TE93ef+DrW2LgB
LGoOuuKRMMfhDd/cQLcO35wgvyEfAiCAJjeUxy1Jlqqc1WLxNRyo+QpBUKSD3RBnqEavxVpY4FbG
28Ev+c87kgNn3covgTXhF4PoxYAcnSNtS0rrJn2V5zWMEeQubgghJPIORNNrpQyMJOLwk/4CVLkC
dM+fOWcCg1T+Yjk9/x0HKTB0IfhjfacfqZ2chdZGK6/IiwWNnc5+zfYy7MaP3df60ZjhrGJwePi0
ct3X7FlqDzcNXvyANaLDLbJQYnTa4rU+N4oqqQobIrgvzbtyKxT6MfcVWa5iVlQtaNPCEMJMspWB
Z3K0SKmfk20SVU7iMe8GLbjBfizwEw2f1MfUVgBygLjCB5ENfbB+Mjg+SWYxPTAf3OQZYE0IojEG
kgjGrQzbT6gGug9zpZ3XYu8NRQSD4ar2EUG2fBdB0GV3rig9sn9Zo01fdICGIZ/9qxMphKUnPCiW
xc5WohoKUhQWlrKYNpSBC0WKkUfifpUuQTxd1VlPp3TWHaLBqoQxl+6HgT1U1NMRLBaa8+sa7WT8
2DQMAnBQvhO5A1O5M2S9jyUKQa6vumDZQaob3sF8FDBJ8y35MAc2UK/okpJQJP7+t+gdH4sbWUmB
aB8/PRtFlhLAQndCW1Nn0NW7tNmPOgLcMz3YBlYxJHMyXmWyybBCIiIgqH3dF5bz/Xb/p6gdqvOC
JqZgM3hd0d8Kh7K1TtzDpyIcmET0uB7YUrrL3t0eDq8QjLD6av0p2pj+kPSCb+rsCBy0p/Ht/qxs
cKco9U6zrGl1nk/Jw8BM59DGjfDy8Uzkt80b8ttjn727A4Aiw7Pr+3qzE0QilYmtjkMJPa/t/kzh
u0qvXGMavth+MxBkLYaQPTTO7Nja8qPY93NmJgbyoOkY0DRuTsRgxvRq7HtTu4yGmUO2NOR2G0XL
FIxEwO2FdxV8Sdyl8nNj/7DKH9YSDgC9PB/ii6gSN5JTbF1pQOq24eLxJ+HmHaGQ4IJuug2VHtPp
ujAEqshzZjVMFmdpKBTwTjvFduJv2ImZuhiGoKyV5LNxICwlNwTR4MgNJoa1TPYsbSsy9louEXY9
cJWLzP8za3dAy9+V5QDWz5y7rnZgBowdKcFSAIul/WSXVN5u4xbVa9yCtCpukW7Y9XtFbAhidlRh
ZiICEgH1E/WiaMW5JzemmXa/PZCW1/UXce9kG9uEaHbrPpnNgX/uXAi3JkHGxRZl4t0JFQHnF68f
rA5JMR0ABIJMcslWqWO0tmipqcFdtRZC/6h+ERgZAPq7vphW/D0zEM7gi+/FVlLzoJBw8udIE9Sv
hXnA78/WmJphiEWY8/gz57czfx0Y5wyYuvLbRx2NOcH5vRsQn7hDuOP1cgJOm4OFUBtMz+YcY+EB
B2s1WWgMfHp+bznB6n7KcxB8fJUTah2UKZKMsXsXPTLN7SHYAKMQZPDiQoYwN8OX25UqMm5E7+by
Bmvnmpv7+B9Yj9blW0UG64qR3dUej7Bf1W1hRtGlY8dFq957lkBhGruToMnxr8SnPIZ8ZOqU8nU+
bSMH2gtuoTQtkFxEBV84y4JZ7hnzXF1+f3N3PllV/lWIRqG5fjVOJ7VP8QO0CO0qq4zN2alRqx9y
wncwVSaP5+ahnGE85N3HDQV3ibyk8B6uoMOIhxyEiYJU+vbeK3v1mmMZgYfVvPmZ5ggKTWkjqCFM
jvZcW/Mjk+3PCFFJQyNgiDb0gdqTfxCxLPj8Y88Do6ebozJBDGV6YAYav59s5BhamR5vLjEgMj/V
urmL/YBrPAkwSJ6csBpqPEQNsStkTtnI6H6S214OknXnEfwHM274FCezVfvzVj0CcNZogYPzUK0S
PUmwJ2DchZoSjlGae+jAeNVWkbOzH6VE1TDe2l9RX1q0LEaZ2VESfg4OgsXojgViHNdRDM0yG52S
lEx/BtioAOUCFH+eXw137epOcJXzw5YpWD5b3Yj1E8DdvkxmDTB3bh/sET1wiLkBIVjoVz0FOaVa
tjLUFl8KI07925sNXpjssnJL3Lfl5xp3OAsgt63+Ik+Ql9WYGPdNHe0FO+G6f6uqsVAS7/EAcFqz
L0x+QElCXMzEY6ug02SoDRLHIgR+t+U8lxx5Vfv8UuPuxnsKxAA9/txnCJKFMj2gUNSWH1yQoeO5
TH53inTboWaqcnn2vdwrA43Ay26+dKKr5UUL/Sv/2Ou0P8Itra9no9l62yR33QyivqMfD7vznPPk
t58ywuCeoRPgGVDrARrVwHTLgizyIe9ygfSpX8SsWb61WrUVtKmMiE3pq3rOScv+764H83qNq+ci
/wmsqH72nhGFAVrpj4MkH3GKbsK08iq1WalMonnDeB2gP/RYvNy7C7FFjqHoR/asPu0zYtWzDWop
0y8XdruLU7DduEJNfHon7EgvtWLe8Ej5MKGgoxtqsBEzEOfF7z4HPjELvI86MCidBHqzxrFrTtcX
aoafcM7IlMHd7ejMaPaQDchiPfeCF7I7+yG2AlZuHM3tlJ5ztAUfnxCVNAlPZfqE/dHnEzK3mRsU
e6tzFZ27PPTX/Vidft7wY0IdMyVN4Q7DF7Bwx/xoesDx7qkcQbocKvs4UDIOU36EitYNmvI3Ymnc
Be7C71xZ06CETTmLCLHQ4jzsE2ZD5jiOTyoGzv0kLiKHLUp24LkxnLok0nRinmmLNmnDiS4q/eZx
sCI09geHxX/mK4v5QMp7wfQHQJSjSOA5m9MCk95AAveW+FCqE4uEMXklmtVxpaq7RjhyhU3g9P1Z
4ipXMNL8aiNduR4hAiR9kXMkGJ0ll7do441Fd0PY4bjiwLOd+2D4kgFpJbkiVIIZJR4lieGdCl5P
iYPU9sUox8A9GweJzso4Bdk4UJwvD7g+3LsRDDbYojsfJkGW8+DGSa1j/iAuqkuw2WqobCIK8+Md
bF/8VkifEmfNvrqGBfDsji8tRczht2610tzqkGRghWKoZiw5vvWJ3Stf4vviIxfAD5ShUGUqrb71
LlVhrSlqA4PmoDwbMYHniep2yJR021+Xniyahh99la7uYSG0eSGGrh1/TXXhTyCxXBGnvu7iD3tc
y18tfyQWtllAf5h9AbrL50T+tMuJl/02OdQV76xfjvckpS9pJCC7Tj2JH9JGrS8vJXcFKVYpAoDF
7qXJOE7HGH0XPepczptphsLnH6I3vgamjm8QhDFpxVPlN48VOZ3oL8XtbRDyK1IXNf2/o7xEbZk3
wdMRoKq/y+pB6sxQtweAb0b09RtZSFpfwZC1B+qEA5jDKOIJmdnQ2dbPNLWCSOw6cLZsPu2rgPnq
m5yRbFD7QppwCakEhoj0jWXTCJIeetxXf+0bgbtbsRh30Hn0+DZ4ajPgJc0bGrm7yPjLjJXB6VIU
vraxZahDzb2dUsEIRLMSHkvc2rLyqoQJuz/xv2pfZCigwolNFy25RWoHfWM6VEUoCSvvhk1iqxYs
wzYvnFVaiodpamM1eGcx/jTI0kQqPdHVqsRnZAjSV16YeExjJlx1gy1nSm+jFT9GCvm7He/HjBtU
wVNxPOQ6mQ0T/aOTdj7RLeaY2UPNARMK9lCfs8BobA4vFWCVdmxMx2KP9nirdEr6Rq0+w07BLFy+
WBeODlCWgO54eEKDs9CwNUTU70RkfoxTmjk5q3zObaL0eGqcpv0+6snSz4G4FQ865tKSMgWaUabI
mwdNKXz1am4JC5m8zIjxcsC105twIKXVUSmKIVwixRlw7/hQzDorZu8tY1lz6hJRwtBg05zRCpOE
9jtUg495Pg0/SiWUWyQ38uANTAVw08lBRs+JMVjBJ0Uv4R+SzKiJubXkxIhhnNGtPx2WK9BkziEH
psGBu0hp+IOfch1HxLjVMidPpYE3OjID2Vhpl5N/gRU0keywnf/Ag4+sr9LXti9jlt1Q94bwrPCZ
igecj6OmiCkf6LyGjsGIoIJexEWQoOVdPbEpZsMAV14zIwtuiah3QAO3pnhkDvF5/ygH6czRIIls
TzMzHIRnjD1YOIdzysS4x3XRB7hk8oZSnL8P6yVviQ5dW1bdr7DRyzQH/fMaPqlWw+DF05PTL/os
wBNZW1RByK5Hk2KvsjheGRbe8CqGFY/UpOcOUgYrVXrS+SMwAxeT26YlY7o=
`pragma protect end_protected
