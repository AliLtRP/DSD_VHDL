// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:39:12 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
eRbmqLa1FYjC+RPc4mpUstZKRBzAwfIEdf3HP1zqWZhrpvukWsbyp8l1ruDjmwUT
pAW2TAU4ECGuTIDGp6uALFj9LRwcsS/EdYqyGOb2bvX+kGsuE55weyYG17ba7bJt
p5sUh+P4SqyM+AvYXv+KSLHynAdo50ArlcaZx5pMg1w=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 6320)
dyChU4Ritr08d4ff7z19Ojt0E2bmECoGU80XXi5g45J3QSbM3O2lStwWAUlSk58D
JcAt3++mBEfmUkBsR1AZCqT9a3wAOQLOztG9fKqhD5IaQtYvyXEjkSt/hEMC1yvt
SWozhisVKleyjP+GK7D3FM/6I/Ch9M39UotkhlnHD6iJT5DwGM8W5WhaccY+spKU
d+Kosy8DU5XXSZEgSAfiTMNhQ2B2Llyy4GNhGJgJe+mxOiIkT5fUgqQuQpJFEtx0
53lrbPrA8gZ7oTIt3yHK7EXLmV9VMtws3x4uITT81fOkwcsnfVHfqnkoPqVnxRhR
v4Q+C4PyHzZ7ZSsDPXdbaIPQXmJm1SV22c6XjIXOq0vG19EvGCmf+rXFzbUag/ug
mjGSzwCtiBap03jvoKHS9FxV9a5G8In6s70nHeQ1qaz8NoIe4AdwoWsbbrPmCk93
yvI5VOVZBBWVB5Ny+BsGuOSrrgfHM97rNC8zvUBiovo52zLEcM5cHhrJUvQ1b//f
RXCa3DNtP07dcyI8YMVCmpVLtmw3UrrxQapqFo/dfz6lqThLd4GkhLRMU5cA2wN9
mf/ksyjzz1IT/9dACL/0fwABJQNRxRkrTIuWm65V+owGIWiy7Cger2i1cmgrIaI8
GB+6SOdt8svUHDTMxpZSaH9lZvDvY2+HGrVWGfPqnVgATpIQNk0tnea0ZxNuM7lx
YBmkqdR8g8fy2+LzM7D11Ug71RlQrAmH2JFnIMhXYVWHwlCWCmK3OjRQQyNp78uN
NCnmKx20v5h6hvxwtoJfyBi6TBFPLyt6JOGLDg81F/759/8CWETg3KvccphgcYel
jHV7NXx32Uz330rMBtwepK29YNQ/YWWu6VZM9zU0R9BpLXLvcings84bdg7edR4l
ou21FkRSJSC6vShx4Mx3L/A6EAVrBzBbHJEUNrvGvUD53mOiJb7hnIJ/QnN79tL7
A2eTXBrCKTDIcJTAVpCABjC5yDq2NxDC+PPliyHmnHAjg5PzVb7q9eyBUsaSVE3G
1AmCwwHP0jz4+Gyypny3intHo8dgCSEMdsRYNBvMm0PFXGHVGyimTDQ9vKJWuwvT
qqRSa73NsvCPtrXIBgbcbTPVn190av/LbsiRXFMUWMF1QHYc3CLXzRllfsdxBKnC
FL7nhy11rV0BxzIXrNlSbvNLDOIdb9miFUYhqITjuVlpX8yPH2jWGBmEDZCQIawT
sd07oEb5KY77ennxGmgeA0zFmrIphQGJrBxTK4msnXbJCZmZCO6SGEFvFLPOxBW0
925hl2gYNqj3QRSSoezjhVIYjhJLHJRBniAu+oQ+6YwM+rMWh1CA8YxPNX4PSgrE
zhmF7ZqGJG52SlwhAEHWxNWFBUbyDFg487wvsrluCQS6DTMtWS2RnrSsePy8gITn
Q1DG5fRH2MOnknbObZ3wbLB4/FvYKlFOgRyjObkLwQtYVrnVJ4knI61gJn2c41Lx
QyzaRfty6Jy2jLESSrlbQc2FVxgR5l/DcuA3IsAGeezNcLr2YuoYUUCXaUnRBeH4
+LqZSqLGn/vXSv+SMrGktkbvbUosAf2Vb1CrSYat/lcV2OITYQp/LTLIRw+r/YEb
Z1zPHFcG4m2zS4NnmWhS+MV1gqDthJveP589QgfcwONCX6kafJ0toi5gfDm8130u
qU/4YIPo0Jmf0Y8fKoEPWr0xjooT8/isW+ZXkaa43HEXdcxRckYU+3FLZJ0VTZqT
AdqfjM5icz4YYvBvWemS2gCCNLMteeZEGrI9mV6ECKNhZ/8qZnzlmXxMgB7mWSLt
yZAJG4MCAfdUpRqJsSAWJQoXpTQPYZ59vH7sXQrJ5zKUwEt2ozkUZVhm6ZgiQu6q
39lvHKAFkrNCUidpzIFR35U9DWnkfVkjPdUTS47Ngn12jOi/RGiOaJiUbJZF7t70
5L3+BvyWkltOHyIzd1UBY/x/5Qs3+jlFwdPseXFCnOsEekNszQOZUwZaTHzXvVkE
UaqMGEQ4g9jUmFUE8vvCqNGq7uYlLrUpfmEAlMDKEM3DP+Tw39i+Pn09KlHFyZnT
6MeTwZ4rpUSjSitpsGL7GoMKB8ugG+jz45U3wj3HxvGgU0g5a6T85hT4NrtXwPt8
5xgxBzE69mjisEOPLf8KzgOK41TrTJoknFij2PFgguDQs+UlzWc4hGM9rIJvZ4Ei
uxpa51kRQ6P+9oWuLHY5jej6ekQ3nl6tXYFElHR62YXcSsZys1lU5U2EQCxVh276
lMy/4Pj6O3TsJ0ZeC3Mj1Lid6m/YmJP9jNv5WOYxbT8/ww0FTb8DQzp1E5l/qje6
mCuaJ0QF4M1vR5Exfyo1vxEjG/2tkawoEYNg4EcuaOQEBaz8oigTkGb6ts64H6EK
mI5+aOsbf0F/B0JTRB0xnlbsI2GuwoDgu0Nu3Gvo4jpFTqjbI+uAL24LDwAeUTi4
Y8wtkDbPAcvRT97HFlTXlvBBGCTBt/WtsiqXubv4mPcyXxuBPrD0fgqWbQt6Tpwe
NT1oP4Rs8NTNRF3VLAqaprHTcRxKZECAlfQ+1SETBpVLHhxvdEdQUBpjYReHZ2Xu
4tPFC5gVwm+djTa/NMAUBUnpdIDUZh5T2F67+n1Fk+KrSe1j7WTJdgUXKCRcM9Qv
yLg7PA0iU3l9D70xfKP0MHDhsCFh/Gf4jHzq/MkGPVNHSRXSxN3+7GguD8vnKzY6
CNCSOWY6lxaMufWLlLqwo00O1/3jOOlEYaJZfA5ELVNrfRitW60B+CAcANSzOA73
OmpYLEqdiB3aPx909gcP8wY1Kb1lQErkOZxOCBt+STnSAFJZIsTdNyEOrUi5BMKF
METC4Et3ci3ZC7ai+FB7n2nEBGt8k8MIDLzLehvJPV/HIji00UT49yz91OXCBXKB
RcoJwhT1MnEyqdb0E2p320hSZBY7e2j3AL4cbI8ZzEg9dJ9CL/f7kLwz2PufQR/B
MC3Wpkm58Ionduk7oagfArHtoSi+6/p/fpcRuedk84RuGL1ele0ydqsoOaNVq7vX
SLFptQtFJ523sG5PBt4fPAMB9GQOCPOV/1sCwpoJz/91VoFccPaX64DJ2enSUzeQ
kMmEvoqcDb0eLFxdox8sTDkROlmx8qEc3mgju1bpSMfJxggLsu5IP/AztnG0ME00
KNWSFhnK8LW+sV3dcpBm+KkTkI3E3QKt0Btp8UByTTmTX+EbWYwgftIpxblPkDF1
YZRRh9JZU8DFq81gnUy9p73cAeN1n/94R+5cYuw3HCiCGSMTa3U933jL9VhIk1q+
MN5ZsULqrCydn8NOxBkAqg4nC1w9/NjeiCZ+6NCUyNgP7Ce3T5DQrdD76bj1eAcs
jna5DCEB+jCOwdiCnT5Y7UVjYIC0NBaN0qF7tOPTtFHHTHvkeJ44tVBqs00hv9bx
GGnfbxVrQIavdY5iS315ohgaXeLQ0/qJtHgh9PMG5kK+3Vfy5GozO9sR3aIChKKf
AzitEIKCBhbTQ+PxrShlNJqlKGapxgRliJmz9guc0yrQCOUF9ekdoMfDd8K1bHIS
4IWKiRUAz+QNLHfTLdYkRS44YQyhTCNgkSZjA5+d180Sfz1uK+zI2k0o/M5KANN4
wF+XslK4JQYqo0ev+08jXoshocGs8J21E7PKNT0H05Sy27dLF5dXzj/yb9Sq6c4f
BSsE37IzQWe/BJ6sXvoG8DFELZrgxf8aIwHPTlouyqWB5co2c17o7sOruoYxwZir
YsArsyg3GagR1jBabht92jXNH9Ar0ZLY56OTSLfrLS133Xx5jrCdK2r+SKCeu3Rb
GrW0AHx+LcaZIZkxLnuLRWe4/762J/+eSR0rEJ0h+T6oZfhKdP5ez5W3/GoESKKE
gi0GaGfkA7KFI4gkCCPauq2VlAgqcPg4/nYtU4BASs0MGsEJZgyrIA9hVQ8iNtHm
0UEGxhReIwdF0FasNJyvWUdlV+gGPD4We4hQxS3bhSZZDCF7gdqNJCsymoWRSMx7
K58x/ktecCcfG9E62cxbF4aJpll2et8M1biXfGynKE+E7nrCTc5YvSn3GP3iKIe9
GcmesxzqcObENhvLhLCsPxbqovjWvhZOSAvBtyRU24DuAeUD9t4v+YVomMrbwIuP
xEsEJVDAMqmEdGUBc29P/v7btaev54MQ/zwNsPD4nnnvy3ZKyJgHeOjvXyqdljIo
PDEumehr8jV+sKVH6Fo/oJrA+GhVeh5Qk2izsYNSozvnrg4kJVQw6BlUf9KXqmju
F2kASp2V/zMRgdetahERbXdC7Rf4JvE00ShE+E38pAf/LF5bJqr5ryrkXN5cvcE+
S3ilXUfoVDxZRfMQq4Zbus2pJQ60dtHAExlgGDb8WL2/dnHjF1Z+4ANJAOu7eHIs
tc/fjBrwNsBu9z9ehQlOUtdu/SZwbaGXyPBJgkV6MQfZJTNGg8YEr86oIuO4tnmp
Z+mo9O8wRSA28KuPwZ4TN99t9HKReTtPoHdHO8WnrhKjyl0fU7+Mm03bmxhTzNgi
+beTlqzkFP2ep+CELjEhOCikmtsWccACTw9lYBBBQPpFbUd1Wr1EhPx6RommpW8h
AATr8ffoerepDSow5Fzis2fTvJmRJfXXBcC6kbn+DKeOpPbEOb7TkkdsjeK1KHbQ
ad3Qr9QotqAuNpHQDgwToNIb9ntvMFQTqtDoPCDC0pVH5xWZIduSbtHWo1dG4pYp
9fQ4a8DipQJizDhIALOLZsIAO2f3drEKRYr4LbyBPgW+85VRmhymI6nBg3hpizJc
O8ptzv7Iu8+C3PMUMLNncpauBKEMH/uwhYNeZ4dzdHVJAGfksBhqB1l1GTIXbMk4
5uIkoNC3jRJQnNikzpxJeNkzubrmojPcnHA/neX3NIVwhBGpkx0RGFSv7xjMSjcL
0RvYEhteUoF8lNOtKaab8QgwHPoG8nkLk0L3NQDr9c4OcI1cx6P0zYdRjBylIg+W
2cqSzRm+CYX/DBBZMQr6bBEnJrjCTFwsv//ZPiKvml0+tyyOt1Fw5u4XimE2hkEH
nC3N6fai8CfD6IwQV48obuhRMqRCbpyoz6PvgJX504TxGlpf81AQBRDe9EcmoP5G
ehjue7hgnn5yBa/59pFmdNtiSD3SthSluSWZZcbBuFy0JMeijxu38Dz7R9zXln8c
XGpfgXW6osCyw/LKwhlqKydZfaQaDHT5LNZ336J6K+RB78n7y5mHWYMJ4G+5gTcT
NoEJ890Itla1PEL1KvCDto9DSpEZ5j37Ov4g1xOYv1IySbtlsBG9GiSpxhBmLtxK
MCWTWWloiHB8Zzx+bwtdRTEvdEPBIwB3X8qnTzIcImIQ7Shl+mAQtoXubmPxA+F/
3XbaRBrnkAWX29G7ZqyaUcoUKqp+N4NIMj+M/maFrNRoXWlgj0v7B420QnJIaZbD
bf1BcaAnIYPp0tv1yytG+/xVyBGFiBRPMF9uvzqeCUqN9Si5fMFIh26XePWEcVv2
9j7mZOhjdWOdjcrRZnc+d8gCqutlL7h3KPcy2Zf/ZBs416fn+qOxGKZRW1Pf1dGM
VRHqScHI0JXnvHfXP0ggcmHcJdBOxlavqArvf+SdMyDYQpLnnPpyam/iR8z+ayfu
SU5VUG9FWtzsFYDa1OhAFILZ06wtlonkFLN+yiPEqTyWF+VW1PngnGD10nnf88l0
G+BocVit7T9/XHhp55MRT59GokqMPukdSaCIvqw7vIlOYzkpKALPBnAGS16tOCM2
DLvDHTgMXxoxN9QgfNHVja0SPSU6kRd3bvxVZfgj8K9FmYLstH5qtNYmFUpUtjpI
6MTe1LBjlQLo+8uuZRmyl51UyqlTltaZk61lygO+SZfJceolex+QyhuYwROYyem4
6Kutk+hHiQY1BUDD7NGwsW/7ES6hpe8G39UD773UsataPfb1lVTgT564Lh9VBdG+
6bKlEg5X6ey0Bm+JEvKl8v8BzwSFRxfQULw9L10zhw/OMPBdfDervx2XqVib26+1
MaRNu0JsCZxSRkG5B8bgf+/GvVZw4Ru9zTcIOlds+iddzHF2YPbOA7aMQV062phR
QObhZ68nLmYWKi3wGKCuvNZuMk7wGocqZ1tm4UYSgUUjzG0SRd2x8eY2MHe2zcip
xv9rxA9ih0Mky/XYFrJhkqUQ6Tach91wDmAPBnFQZ2V0E0vYGSAJ+4VeHQ+obNT2
4m6qoWFzXcKNxTbEIcLc7nv6PuFvsjyP8eDFDsKwoKquyege6URBUpAQQc0VRGcS
LprUpsHD+PqlIdqItgiEPBw5XIjD24onNMz3HEnYxc2gX5KcIF/9BIS37RNQz7wA
hnGuy261iIp0itmhInv+er1ZSURBvrt2KmPUSnpd3ECUraNw1B+idNnbiD0JaIRD
iOxqHgLLD2P6vi0Me08kF/x6UIlL2wxiusrZipw/bCWhiB6d4hhTlb4KhN2SZK4I
QgWRi4lDT2mJ2KPo512OQwTj4mpoFgK/5iKhuXWs2zctxZXFiJx29nOU4uP/r24k
GSgyGPcYoIGhSkEZ4ne/HxgTwcxbxTqPryykqk6lbL3YFdZpKsll0LKrpWqSpidR
ejNigbuyBgN+aqVxXXdVtd8kPq5qkloD5BQwHlghGhJoiY2ovnloUrUlvs3HzkTK
uyCIsH5eEIgrcdVdQw65ZgXByvoS8dlfwSfB7tP/JSFFBatiN5Tv+GKv3yg0Fcv6
Y0eLgwiasZAZXSGzYRrlvCOiFOt2yqI2B5obLaMHv9OHdfWWObYoRRiDSKLMtBV2
vnjE7cb//hrG8ko4R6m3f0cfL3s+DUIRrX1qEbAudQcxCSiW45CotVf2rplOVXNU
6wDR6vBmiItTJtt6CnQ8NzqzIn34FGm9Gtxzo1sXQS4K5kI2aTAGUmkANfLHGbRc
2Nycg2uhnVy/6U9ay0AoR0gD6IbQ7csqaX5DS9ITpr9T/YM43nX3xaSQOZRY2Qq4
PfdlBFrLgfWyGPH9WHNH3u0qhzh/bBPLSJVh70gFhi4Bjkn8sBCuNX7yuHIFTLX/
HbpUNdwInEkgIgVflZTky4tJ+mJqh3hFIqUNHsDySHGGtm2q0CvmyHmCH7sSyYx2
w2qHCNdcNw8YLubNkWHtsP36jXUEeCuvNxgqucSyGSn6+DOjJqPtrIhjnwufEQ4Y
OeTs9x/oXXxiNBhuUPmCTKntBefxi99zUoLkHvHAAf3GdN2BmX243itqvxHD/HD7
tYNCjCWK3sPIMbnnELx/0DC3VhVGoo5AQ5KfD73rxx9+NI7h/9aEV+RXzNSSk6t5
bLWgJ3MtjaTTlcLA5wSZ1zDhuO+AHbQS8QMsO0IHbAXJ5NeFR3LOgJuUZD7f2PXq
bwhJNwWCKg/1VPfcjpS9WdrwQ6kHBTxfwZ1axydhqE9QckYmBGxqWddo+BYfQr+C
czbx2w1PiAfTO9xB5ZzvA46TmjdayldKmf6R6UMBXtjcmBPJOC7Zyws90GadJNew
jpDJitEAAYe0ulMafCzr0EBD9ix5W7SCz2J26v4hK5RgRl7H7BhoBMbsTEkN3iB2
slntwBIDwlPUf1W5v10za5vbSpbTRTIbAScv4qCj2NlyJaxfCcpd3vnErOjBEcws
WzCTNK46rWihVOHjSf5SkrVn0koXj+em7/FSJ4VRKfpS0moV4EZT8NA3g1U9IAzL
xW5QRfp6iE0m+9+Fe14dW3w4r+fBYmZwbG5+R0e1jyMv8MtlM8Ve0RGQU1dMMBc1
WBcuwhBCCgZWkhE7KcQDQyXIZ/qZaOAYtFB8MwIFfSJvLyJKHvPtkwjQ4jKKjDgg
AZ/ZZrql15pEmmpTZPvoK3ffwY7PxbrpxMeBXzs6jx2EpOvsaTWAD8CspD+8uo3y
jcfdNzTmCjwGwgoV86TZkN3Ia1vnCvcosV2e0LWSaP0CYgSltzUphGNU0/oht2vi
kD1h05aDAu9n+zUOmjiZwh0i+U/mrjP5srIP4u7EQ6yc2/EPbTHm22tE4a8QDmOv
+CF/EYPAAJS0yE7Rl1ZRIvLm2LlSp7sQhsg/AGzZRLRrnQ9pepGBGHN4LiVPc/SJ
N49vHcJmCma6fWqEaL9O1UPOsitsKdHjQeCFxigzQvhS6JbePM8mCb4PrNx82G3x
Y8ehoOrtHUGy3PmN8he7T9+Z7goO/2a4BTeMRSVEk46w9Ibdch62NcO9+rp9Hbje
CdMc1L1gXvprQ2sviQEG1uUUmff1Uk6kNL35mBosEPkg65SslUhMEzZq3E48H1uI
cr9xCe5NA0LClzSmLyzd6t1xuo7VpYLKRGlnIA4e4KnjybiDlGDRN074lix+mykF
Nedxwn4ednxgnxNgBsaYlEKsTmGjA9zu5obP1ejZEE+IpLL/3bZqG5aiyjWjaFsq
QWlO0yPd139CwqHGaahwdEOKMUQAppU2f47BwheKw6YsP2EjfdlOC91r8pp2ejC+
mKVveMgDzpfuIR1VeFb+pMzZwI7UBAJ9tb0Yzeyz6q4=
`pragma protect end_protected
