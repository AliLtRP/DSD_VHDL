// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
stUNGsFlPIHfZU6/HWzhqILXkErMLkTzzMlsFHfE6YXztxPdY8vYxEkex0oa/9mlESfl0JrKp0Tq
110rkWifO1amcaeEPOiodFyZrC7M22Wnib1xAidJpq6rr6gM/ViYDWrdoOyTLkCohXe0yjfnfPAr
8nZLryV3IJ4fH+7JjU8wqd7VJqjT2I5mP3HXVNqH15A9tG/ahSGEVWs90rWvmnOUn+uO2flw83QG
9SeoX54x/7TLnYo8vhQewRN3lI22ms9rAAJeoGiOZEgCFu1joLblDPAOoOACMVjkp95wiuL5pUU3
3CFhJi11Dc9Ng/kwofaer6MSGrifQjzULBlhww==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
Wb1yR+KqHAwj4xzPSrLh8+CF/Aoq4ROrZdYzT2jrPhAPCf7fmStwN2EhzoPvh5MT/MkHZEcUuAdr
ZFPo1pCwx5wqm0RNgCheswVYRN+g12bW9uwkobq6i0jDfHw+xaoa/zSG35ZWitNac644To7PmJ6i
ywApUMjKN3h1aXMCVL4sUQWuYX23GpU+nc8RnLcF6RFpysR1HdbliQslqJrmnPnMsOaoTZSgSWRY
T6V5SRLdo/UYNwtoeiuUk1UdXJsRWv70WazJ/+VPEsXaKbTItjYpqHwmiBxDgdr3Ic+bO9jUcvp4
j6fkWz+rKQigqP/OrUQn/T7iz4g+qu1KF/0Gm/030tmGNB+w0enCHr1o5gh/NMBEwftLId8kzNse
I+92fhfpBE6GdlNc12Gxj/Lgz9T1/mabxLzf7zW9q++QIjAf84RgEZy4KsDCbNVmJW3nO8LgtjUA
cC+Ru6N/f2lqJwG7qOdfX7uhJVVhRH8dR8YoXNUnjjjcIX5Ph8AXgvLgDgIWWLWcjqTgYo5XkdX1
zAEOkg74lPz3LZi5wlABCLXGQQn+WGE40BA7fZl4+a8wFevQnrZhu0JOQT/Jve8goyWa9e3ML4gV
lKkmm45Kdg3LyR5QoxvU9GCzMcTTzLctfNm0nVas04qKTjXd0wO+BOWea2PA0z2Wwb3kbrq3A+vv
c6UWtIdJPDjwftVpmn695LY2S7++9/pz6cD9Sp3+HRcVl0P/lg1In+fOAltpuVuCmlcBdg0Vm8GS
dl5KTME7bK/KonMwiVbaMLoXa6Dxt3AMHag5tOGyGum5u2rP+HPLX8T/aq/fl4H0CmboHNtsPpq0
5tiJ46TAKNN2IZDIyeke6vnWRG2jc/laatvFyy5mwqJBgTlErMy6zv32NebwI2w8Lp3SD+KpnD4D
Un72Ymn+qSUQHphIxyl2M/cqg20xU8S7VRElTFO0FIn+fLGdtrdAnynBLWXPUlbwgvYG9zDuhAoF
yiliNSf1eIulNV6nBp2JtAY5LwZ0xyUc40U5XowB7vRnOeuws4AjEfj05vgF2EX23E8jLd1KeEC9
ppllBftZlFmVijSONJRwwqCCpoFKV6/h7e0Ul8eNZh6i6ayI1CIF0m4VS9VmEcJ2UvdFRrcyR2hu
og0c5fP3vba+mAzetK1jEOnS3lyUOlns0o5gR7Yimlif1UzwBj0kSBEh6JiVrIRoz1331uyHc8k9
PZHgjwBZhTEaE/gFjcLv1ff9dqNWTMupHK2vRWYsA2QqlprjsfcL4oDByOHiuNqrL9bXN99QkW3x
EuRqkkcXtkfUSQYZUkuVUQFcuaICRR99G6N9SiIldkEhH5AZED/xSP5zD9uHQcdXvfRGFcHHu/cQ
ld84dPrTan0qRRU+EAqJu3te7ZCcRI6QFY6yuQKIYBlnVz0njTBm4B36TMUMaf/Pdjw4QfiHjHnw
4BNllqn1Ii8EMyIXeO/agxGL7mjzqBBbU+eyVvTFd6eMMgF+eW7e3ug21XtX5XvJ18b1YhZMlCxO
DMDaYkLNA6UcpoiP5F74bH2psAlgrOu2gJWPUFhS26mNVxj8l7A448zihe4emwsJUZbexwI/3giw
6/SK0wF073jrGqhTfd2lW83ROjkdQmpwU5Og/KQp10yP7ksVTiORDuUfHvEAO/020X8tYzdhtks5
M0LAJT/596OaeIcmYOkSc5jXb/WUof9ecSEv+6dQGFucNRCk2wnv5CIikIFHtkA8mizDBDfqE0yM
yK0uzDDBMowTh75l/MGCmtkzTbS62LwOqBR7wvuCuXbaLIs14Xx7H66kOJWPpsxeRMR3opvfTPAP
nbPuRPpc4UASihwlP1xfqyaV9774QCtIWvMn1JrdjgllB4+oQAg3aejrykOSj4HUlFerdbkKr3Vj
8y7WUe8gWQzZ5Bl6Vq7hgqBQgzCIBYK80dm7pBrwOZOK883gocXq1Pzi1nUJj6hL7DacZ3RWpm9a
peLQCLhWgS4BlGNPftnvEoAWumE/52umwYfS/siHLbV9wyTeRpOnMZe7uVLVLNCji1ItwK+DMAzq
kgjXE9lQYg1uybMt7sPNGsiurTpwZniav//PwrwsFMsNn6QJdO/7O6ithpdSkOmQ+xUMrstcIe1e
DPkTcVqxdw9DJaNdfh4nWHPvQzGT+ajX1Sv9eoR2b7OOcauBeVFbegT1o9Fr/Oi7CDoZez4qIuo/
j4UpFQDu3h6TVvd7G6MY5KxQIFTmPmHfNNsdeTe2Vol2pSN7cf+HFAusm4/TIlmpO/co8d/GgdLe
e7o3TPIArdcS1nda/cbvFBhc0miUjZb71rZGyaCH+N1LwPjtjGyGix1P2ciEnJSfG+rEIfmacFJx
vAp00Ve/hCTr9D5sUjd9bLpvoF5xGX3I9sKZUmA1MqSOLHzKgt05xfgmdJ7X3eYnpdOKDzQFRaWX
hzY5rtyAja68Q4KberFez5R3K6KTAQ/6Cjh+UvaRYqCB2R678ULVE1YebkrGMyE1lbTVlot1GTd6
Vx3zuLUEtdya/+hKJLIi1YEQ+RFy9mrBY/0rbhtnp0ker3L1iA/qDF6TGqzODC9oO8jhj2eLsnAU
sMMnBJob1czinBzUHDlU8tsiMdVXpJ/oIN1XspdMGT8lJRKt1c2g2dCzRxmGTDDQJAZhecbq7Y0R
4qLRNJlQREiWUTLK4+T6f3BNMEtQhs0IxMav2BuO+NWr8IQu97pF4v/68vHvz2h6k+Q/AZvVyMAE
S6PBp53y4Q9E9C9Ywg8ApUQ6ixPlUEcdEOCFbs3A+DdOcNRLfybsVLnJca7VRB0blLRUWtqhgTqB
P11o3JT8Hng9aUMZvX8ume5h9HD6/03pB0G7OaWZGGdouweOxsKvzNDUg1/A6anVowsqMf2pp9XX
yJg9M0eYuL/t9sJ+25XcTH/U3XDeAmiRmXtzOthxUHrBkkWH5jTYyLJLsgjuIOOltISvTHzh+h37
DjYaXNf9LYIFm+UUiuR1/K13MIBTtGGB8ekmlJ+yKUhDutwkXhBq+dDxsQ7BdpUCYbLj6+u9BZ+v
pW2pL7Af6t1KZMOu0tBp7Od6PUM3XDE1qITmjUHkRGcogdjDJ91okIj16nShC9Pdni9WT0rKDTc5
5gFjAfkvG2PYjQdXVVSJ9R3azNl89iQlPvteGgbj2ypKXL8lfsS+6nVZ7P5xtsyf1oxGalhZOe4R
W0yYLrX8UsDQdBGPR1HoiUYiKmJg68sTW45pQNRaMdUMnc+xckZnuOB8aiLfRPSXYsJY6KIUA87C
kdMQNy8ad5FJgF+lrj7su+YaOU8MHgbsAT10KDHvxCrCcJk1mX/wTGsIqBEGV3u2bnoiqvqKg+YM
GXT3PIcbvwclIqYWTet0LQIJkO/lDRfzYAhFdFcuRDL3DcrztkRzXqUF+CbQH3SsQvoZpdR2eLJV
6YuhVsuoFyvfA/lj7w8jRZqzEhj6UUr8xOd/y2DL/D1WIgUkbjWqiQ/Jg0w3czwygRblXuApHTuZ
luTROK84c4fKHsg/6+dFR4ZvH3JP5olllF2siLWx1LLd+7+WpTU/zSvAYTCg+fZx3fGjo3ewEfPC
LxDI65hQwP06SnO6Vxc0SXv4kmTTWiBiVhF1fuC4kr0efBtaU1NQWZyMrrbHhieoRhPxwW8+mbW0
eK9V0ZB1xC0RPn4hcRQMtL8+pJdChrAjZK0rTeOiNFC/WUSktVthoMUfZgXGElQZRHzwUvto2js8
baOA50XA4NfnoYJ9kRJGyfyupu9glZbkXqvN2pFsoe3lSCq0rBJLsEu4Xe2YrY/bkG9k0Mf+bhWL
w91pHEJNkDK695BlZkCB5452wYK6UKxa8fDmwqhgKSiU9muVCbTDW9IZKaRhrORbTypAKL/4EhAG
t/nukHHveGUR2CsceAy3yM16lcbRVu3b1DgC9poBxC+9ktM0nlYZBmQpQmA1FeETs3Tgasos6TF9
wEz/ZEyp05pGrPmuSChpUyWirjSBWEZTUFfHkqufBjeYIbMwfuF34gNQ7E3je1k1WwCXboxg0LmB
JwPU3mBPMNq9nK63sud7ODIc8jCyof/+3GFWti5xoDd4x7BgF34QdfHMgroP2WzWMlbEqBYdjI/B
/nG3xBghqG4yLyPCDKGHFEiwLzsm/EPOvzOxHE126SI6yzx+g8fFoNO18mOl3q8TKaO2xuETmLgS
JhaOpraSgElC88ZVwwoDMQ9+X9uI4fV3AIbq0VTh81Ae5JZXjVBEPqS6nlLyM8U/QLOEvkJzm3Ut
OnBAtyK7yepoj65pmgX1ROMGtr0XV0kS7QIbSa039ipTD0dpxqw6rrtoJYXdJum/qCpqAMqYCXdX
SaRk4Q61QkDn/OFMdlPkdOAcszqzsT3WH/V/gcG7sZZ6YYU5m04x4HZnPjbFxHXCj+fzucf6Gll2
48zHIh/voq6PRUhWh99x2s7SrBpAzUvRStpsu36cne6moh6j/abxE39WGespYYzmriwWKz4CyFx3
pQZ5Llyval3KkXof8U2c2tA1Hs+IHSbmipc4EpCkpPjSREcLUwWEi9/WWWM0PwuoZu63khTcIW5/
jIlE05rJvXLrza46QP/CkjW6TRt6VSGr63RXGA+gsSApkRdzqonAXr7FMhdCLfcMChDPGkHhnpJS
iQ+HGIjGjksjWr9E9kYiJcqUxPYJOgyMkVoiVnm0h5scsFx1U6b0iUd1JAkeCsjlLWpFBp/NbHHZ
Cbmic/5W3gYlOQWTqKDoOrAKCMATGt5/1uhUpYjGpIiI3MvUGaMWpQs6JRRBIhhEmOiAGFUlIMK/
EFMNvaL8bebtJMVOoWBMlTrD2TkwnsJrDU50XnWhOEDzo96mQMw5p2LaMJSHH0Gz7DSdlR0tZFjU
UFWT/5Iufv88amqHxPo2QiidSrc/D1/cdTigkbC2kI2ZwTDund0fOiejDBoOorRmFurgSfcFHOJH
cJUYETI2rJyiEz4ok5UKzvof4gWFjnI6mhal7bVyw/AH+RMCNkOPj5AEcFROms5mDwmqfY+Hvz3d
q6cGILcmDcA1DFbAv1H/0mQPpICfTcf+ar5XJFdr4pI97/J8D7nbsolvkji/tg3PLIg85tuuHfnl
YEyypb3LRu/BHmYSats4zNVsnsCVMc3JS3DZhHuSIzJSTv3M90fIfJEmMXfEi7V3jjoL0npg5+Yu
i8vQulY6gYRIJ1RQJnew/+YYtO/ot6+T9IWxemXPljxsLZ2wLhqOmikU19g50r/ti0cT8A+8OjSt
tO1N+wKXQITJ9Ubgh9pt3VqxSCSKMpuFFzviw1A7Z0Ctb0PCEzv0YLO73A5SRTAI/QGdzKNPsXTY
0L8XmhCamyDEYmx8m5rKoBKe/d7kFji9M41oUB66XrHkra8pq+KOxfxczvoq77Llyo+Dz82qAUqf
IrA1+qaQThrKDjv/11sIQoRDKNo6ABKy3+l/I+h24FiKZ1b/XkNuSIY42zTeo8RCmv3W/u9h8Mzn
0FBHt4CTEbu7TDBVRQjkyl1O5XDolaTUbHodrvni/c+8QZxskiZU806ZgHyMLpYYvB8SzumqetIf
vqOIU9lIRJA5jinBZ1EEuGjQyjb3jvH82PfqCEutl0Quj+mZqs6A1YIkvgAi3p0B/MiXrIgb6F8r
Ur7zK2jWHoAV1M4pVbnGRepDpqAQNwSemS6pql677gsGxpWroH0SaIQkPt0Fli49O3Tbb/qd6fHR
5kfa2ErXc3pAf9iZoMOYudKwmKZygo8OCckpEQOIc/CqT0ATb37HhnK91vdW/vKsj9NA5hUljd1B
PZahfx1DGG8gxC3mLKpZb4zNaeVAcDruI8T4tuIe1YybT11177FVlZkYZKODoCzfTmJSh36cVwkw
HBVQHfG6aYySlPgMqtey9eOHVCyjXbewoQKILHCjF6CO8KkQ6EMOgldJrE/RbB6Mp2u2gmmwtOuS
Dlnf35n3+Y+IWv5dCBSJp7lU9zHQjx1ImfJFH8jfCnHLQrHreB45JNju0g612Nw0Y/Nz5nzgsZJC
ZEPoKRuPVmtK1pGOymtV0OLZWMHyG5XWPMqqDtKSY8HL1avKcKn5gdtP90NYKHkfgbGv2527pvST
mxPrH0Iyr6ozzJ0V7sd9YbFd4oX8v/rQEBw2th9M4CsdlCyuspM39q5qHjDW8FZSusGDp7T9HQzn
Roz8y8KQ2xf2CWjYfM+CdO0NQ/PQSNBh6+Aq5u1k98Jdj5nvMKpgC5FzR6gPi/k2Lfbig9B6kh3+
sX7oSWl9PC7pLhe6zQvES5YOUAqBqw5H8TIPhHmaVcEa7O0Ko+GWQUrsTDRck5ZIZIdm4uMZJudC
QZB21tkB5ZD5//u4ffdyxVOlwSgEF6WRduGH16l794eOeUI1atFyyDq8hXy7bS1XNNZAo7ozqtwW
41XIz++W3EYWI5/ZvsFwATsX4y7twec4FvpnWZYR0UuhIE8Q5Y7Ha+zCbQLTT1mwYO6Hj2MFAyxW
WyLNH1nhZsjAdvQLmS2sn90Ogexka1mQ4aLnirDboRMjqeKTsZ+zWwd+1zl7a5ZO+JFIbPcSDnKq
X/MtEHwrVtHoqhqKP6HxUd/M7YYiDwdfh0HVzV6SFINxFBGYbxQRWOw5/qjkB499bDI1v3hXGc5y
4mZ/GKaltDeANOASzQFPxzQvlbIZYQjkS2zmEngmgNqaxVDMHD22w+3G4BLdir/cOkSqIPX/DmRJ
eVw7T4zCXflSylm5G5I7UH9+KRLQFL1+h1TYet8CTxqHUsa2+dbSmpvoRJ1oNUlU2AOk81L95zvD
6H6dSAXBR02c0PClgnRnj3nUZhdtexQ6LKPG6jQNlof4A/D01bGK0wjul4BDmbE6Ggma9pEb7PWd
oa1YWdPn82q4HWUtj9KlbBfqIzsO8r0GnQRa7vY3U4/IeJ3Sz9YlCSlOccOtCGxo9AKVD+YALv4m
hZ6ptz0KdVLvP6INvafJLgXcB9zwKgMrxUSGo2cg5ulGfjzvMBxDnRjmDGLvIsRqymIrLFp51GNM
bAHSSeIiYE3laQfaNWXd55Dp3VvRBAZXgzfOW4NajRSYyIjUdmhfhzMiVbGnHR+/rscp7zOvwyFn
B6J1GfcMqoomPoPGuFuCar9m5P4N7ca7kQScIeLNS9KwHoVLwoOqkHk6FwRvssn4zz2deoNi6cCi
gmPknv51Zfq7FEqcPSW4N52Jvy6Nl5SvIfCqBvOtPVtCilwQbn5LWVIDhtiqlkz8+Pz6HILiZb8V
0O/yppLvn+nl0awmWh1COyHbLRY+oTFrYehbWQlgEmM0XC9rQCw6u2QIZ5aVsaYdVSuk/An2yG5y
qjDJZemKKLGK45sBcATpSizgX6lxZn5qHp5n45EI88yFm6KsB07GiqYseR4ULlcJYc94V891ihWR
1W9wkSSWYZJqK52nPjQuc2CZ8+Ub3G/PcnMyQYk3uYLPcPPBJlRlX7171KoMC4tG6FTGnjtZ9oP2
o4j0xjn6P7p1bptdIz10yZdUPNcRDVbki0TxK4peIaYdB86/2zjyPungIZx9btypXKwZmrVWDqZU
TrNRs01zkrxaPwCInH71DoaSphTAwq7AROTQD8MXFrZ+f9HyN3OZMQEz8xKpBfZA5ftix4gklcIB
NO1pWsi8HDjmHzSe4yjVEjB8ca09YgSH/5H66Fpk7tIrc72gXwgrRPeZRExkyeIxJFgSLLJtKuuO
O2IJ8xksjO8qwgh72osATCM4mY9M0aECCX/4Kxd0+V7Ue+rdw1UYlLtqgvHlX4QpuWlpETIFYNZb
4DqiiINQOtagkMaUAO87YwtJu0gc7XCIQi0ilf7GyX3dVWpXVaNdn1qP0m1TSx4cHyShCMGxAQ5k
XhcxKpIc9iryEYLIqxlXz3WuZOi9VFJwY4kKMwCqdqVkSp2sXDqNBRVjzvtCllqQwoVpHCjZf8WT
7Dmgm+N4gHhJ84Z4NVZcv6qFMlwuwkH9PWg+VNKpQbzEo5/YsrhDSB3ovD0ffI7+HuLmOiHY119f
wES93A7eI59umjXntRgClKfYgJnk0jZ8ro2768+gAahVLEhGEtu4JInO0bt0BKr9jTBqmp6afguB
+mlMWppqfSCklIn2GEHVr3Ks6392DWHMJ910hPns52oAjx08p8tW4Nq/bG81ULq5PCQ5Z1bA6yeU
lsM/KDprRiE3P2D170v+npHuF1b/UZ7RP37nxPW1kMvMxnz0EuK70j2kT2F77jupY3+5ldRe5V7i
Fk5qi3xOh5xPojXyAq/4hRj5PEJi2gTMySY4xrumzLhmMTOOqxeSnyfc4MpiHrxX9POTGZtFdmGs
DmESzYGx7hPK4ISQmakslxdUOXxw9WGrfSaPYpNG09wrknigyCIcpYEhrcKo1y81PRttIN+nTbAN
RLuT3BtcSbK45n9I7Q6a3BDQwAQ6wi2xUHV0zFaqiMEJu943Bn7llSXmjeXPbnRtQnWH29dFzU5+
/cLysL8j0e1sv47L28XpMCGx4QE62gi0B8E1iXghcxgliJE76e8G0C3BTpdetIWP3aUqDhU4ynCs
awhFQEegekhUERItdpRJVUppTlxsu0MszJvQsM7DznBWh8Ef7EQc4TpT2IOQbTe0ra7uN+PJaDJG
36PTCoE5oQnhTk+DQxl1PHXBUeWGU/2fNsQvqAIvN3cya5h6ANrHcWuPjBvIer4pPj2/YYa69JNT
0NEjjIM2M2NBLGzhTfOPE6E6oRYBWmz9eTUotulC2Z2EsjlWxfmziQnB2qEY4enGFN65iJDtqBHS
ky/VvPsAdksTBQsCNqdtBpoEz5nztxlNL8d59hmug0vO6RvN+YKkTieBfzxMuKMJb+cEXfZdJQD/
cXAwEC5Q/JjtAFmFXl1Rdsf/rrhTlAcXnHVddxPMU6bNhjFri8CdFVpRmsYktrPhPzSFQTlfUbmE
MipTxexxnVZrH7s4rBR7q6OKe3Gq3xLCVZqschJBjEW5pwNRBCArG5vARUO61ccdqLxw41T5AWuN
Cwn3salPvWuYDSEV3l/KU+Pt3Fw9Z1yhjA15iEyFARdrjn1oZUEcdo+oHDjmNFyzC4b22rRAAPnd
Xq8KfJJs7k2bZBXuAdU+P0jC06wWWNPsBAA/BBdj38s9aAJ9Csqm/s8xK6C042Fe00NJK+Z3+O9D
jeCQ62zcODu0UdHCvlwUhxxd5Pt1JNqiJWSSlugCr/ml5j/YjvQLtOhkmIV/g1YsK6WKELWYd9Tn
ChqKvk+Fr4xpTsheTo8en5JzFuc7C5cAtYaVd3YqrXDczMrY4u0MbLqciGeaCt+D9RVue21neKJt
2mXJU8lT7H3dXXQ5uV07oW2YdkMnvjrhemminWTVU0+n0AlGBXxFYrgoJMKBs3Q9W6tA2CE4vjPb
EtVT0qgAmh+CmwJdJaoQxOPBZGIDSY1423uGUmgKzzP0YOy+qQdT8q6F0QNJTxSaqcj39xM/MPcY
+vjBHF4S0qnfTx6+k8O5pYi3dfoF57+TGiEr5JunqcjadOpeCaFtioI2YAl9HHdlxCb65HpHSJAt
vM1ysRoANWh8y1/F3lWPfKjXHYi2A2lYyhEp41JtlFj0tc483yCXjpYWABRuQc/aQHqQIYXBZV1m
D4HMjRkCSEyPyuG2m+hZanrqvpzCFFCiuaaM9OILXmhXS5HxnRFDfVfCSrrOAxlGq+UGR4164Mzz
Fv44GNeT5u+Q4ttlYTtkJp2XdaxpE+1sSHjB+XogaJxiYG4Thqv9uAhVk95mX0smyezmTxI6lXto
JNkxp5vl5QUOaxurHCquQLZCgRg1jQWak40D/lKniOFZYv4r+4+HgcWRv5jQhU+/ZXTubjba4CV4
uPPzg32nNsqvUa3s7gz2ZbSBk/5Z6z+VBudYoWXJgdOYXHydKJfs+2cfHAYi8uw9doKr2LosUesE
MJpe9KDQgk6zWST8zfKxSHlJo3xhpBeqfvneMFfYNTjHmKIJNqjocGeNkfJhsodmQguhzRGf/7ie
ZM6lmmrEtXqy5eF9zGnUNMSRjjWNl8cdF2Tau23zWKUiEUNkxzpPyCrNU/KWIrk0GKgcExBaYRaL
HF2llZKCCHFWAM3sZ28v2zHKCHjbhInXzmp1IAHmfwdv9auxZT2gWJrM0bnpz2ww1MaTXszfpeJF
CEPvfDkGgdkz5n5/7Rck0Q29i5lv8kz4mAmOFG/8eJUrSbCo0iKsx/2wO9/gLnVNECjRLHS3zTJ/
AbIcBhsb3Yz9oDPOpyy10rCrz0EpLxIQHHWWqX2nW7cS/gDD6pHKdN8QGCQmp/f1Gl1346rNSoNh
z8UJREvucUUBSYa5Z4oN1Z3K9syzjrgnkxp1QaiF346JpMNodfbEzsdRVgl48K3/8qbVroTqNCJc
2icRAx1uKmzNPsKcEJJXtAR6ZEB23EmmPxQwjfLFvoHbsDR1k7I4MR0y2Fzq4iTvJXUCM1F6ftPW
K2u5EOoE4lcJgpU9MX7pjp5wYPp0IF781HYQBlDYIhgyDtjmtJ+bQzXm9mbxzoLTp4Y9bBxlLoaZ
jeZi0H0207+kLTL+vJzNtma/xTlAjKlc6LmupH/I4bpAvvPWBK5N66XrJoRqTjuymGhNDF5A997o
82WVrhDfl7rNqBpsqrgRFmcpVw1ydE8VjRC5WpObWIHv18Ec+R8CNT+NBmxDeDywAzqIz4meXdtL
wcRx1LNCPBgLrIyQZJOYbUO6CXDLGvmfSbhRphalekfLpzRZPJJFplqonStr+SQUD1kwLB9AUz+p
seQ2F/FKhnSpqsMRec6GUtUZG0oTmMlAKNQZ4XoxEj50sDswOhnJ4Rw/pClkbr8Xb5EGJ6NKCu1l
7MNGiZZpZEy1lLTCgsuCk9o6dKTTN78jruVNVTIf5/vFkAzclhznjFMYqXgclv8VRgDpoZPZrG/q
92mPhA1G8joumAzGs4R8AX9VR4hvq2Svpt6pgw+YNxw322qB9LKnPu1muhxK4vssmGFh9WiNpmoU
BkGsV8LFB0hez65mPFMloZZQqt03KLLVy6Et+7ZLieeoZoRZ+LZHpNBAmGMRUebrLnSkxx6J1FuI
uLqk9KdWB+9nL3vbqIcKutIpbFYsFhWIm1O5fWeDi6+zS+BAYY+rADvdIkmtmOqiUS6awrShQJET
mrOcujXTUT4kT9CNG1shF3E6S2SIOxXJtHejppR9I2u8mtYbQqPjbHZAmx073Qtov2SX6Kibhgbk
PKY4NPy9hVyZ1/+UTuGLSRp/U3vpRS+UeXj/gsntid0pZbLXTxPl7v4I9wa+Izd46W2uelGK86sv
jiarSvB1+b5n4pnt3hugVgZNwCtj93UEtXH9zEV4H2eXLQSUWGCscCbTJUB2jNMWpw0+EbQyaxnS
1lLh+4MCZe6v9tk5+kg7J0PviponDtYQQrZDG96sONxqHQrnI6d3T+tcXQuRChLItHDW2AgxtxfG
VtYP13vsCT0TmbzGxEtRQon1avjW/NVFgO3spcUL3LEc9uTmXRC6tccW0F5rvLxSDBhOzMH7lWGl
2JtWX8Y8/4LSxBGs8yRHEgQgTfjMiwrXTDsEhpCURL8InW3UcaqDJCw5CNlb97MgdccWZpeEgV5k
2a6JIt9PU3CfiD0IGF8Qgh7pUSU9I6/fzZw1DKcXiJcz/dQvZ2b8ZFz2hwi+TvhVD6ZE5eTX2kwz
RQMifbSaxivGhItu5Tj/cT1Ih/r0AFSqjcuhXyJcZeRAgzd99WEQh40bc9BlV+oR4SPQOcm5ENu2
PljoY0q7Cv0tkSV4DaUnaBpVY7W4iukxjOr9Q4+654Q1EiGESYf+EXJ0CNNjKPqITQdS+ilszlc+
ZAbRuSdyHhBi7VhdigqbtKeRL/aCUj0SmOZdrWPhRZOKCKMA9mbZO+F3uG9hZnabEJC/5p7cwFTY
CZl3Nzh4+d7PgpJiaVk6pv8VJNLAEeYTcw4F+Y4L24OrGI0gKs8wKi8Vvhy82iSG1QhFZxGFbi1d
CdP/dAIhEIEQyFYsc2pwfzKko6DkGKydhsREfQ7m4tmDIcoTQ9dbjmAyu/a09fN2iHiB+Ik+exkt
Y9EGb1yoct+QabJ7RIVYmRw3ncHhTioBpKsvHG7xjEeC+4+6UYeAj/lKEesmY0WW7grF0QvJWTc8
yDZMUz4OWZrk+e9mSoOsgzDyxseVMgMhITKpLH1wzVUCHuQq6xf6XGCl0Qa8Dw+HDrPOT6pw19DJ
ffolF37GkjIA5yQCYwxBRtQEtgpFZjRPdDpz1IbLT2GsMLUQx0XvHjkCnGrTAf9c7kGDD5mUZ3nW
aXqlIf1cbvonRaHdrbprCXca26l55fie9Nm2NpxOoNGBCmYyAY1IUvvb6iODtTO6lkbgJ+AwJsEA
E+SNn47iqYuWtTe8WlsjxDr0fSVUNSofjssxVRlmjgSj9rBOQC8j3z4xQrlIZ9U3jWvl/RMgD0S9
Ipx2U52KZQ/wf6j6zhBwAQpmGUpgyck5M62H/o2e1mkdUKyLDkuvYaw2FMZFPSZgcsRUELnUtQ29
q22luCXstF/LgLRALcMFaw7mEBiLLhKoO0rWvpA0K7BVv0f0tQ97GltsbTckD+SdaTA4GvTorxAQ
2Q/0+z1kUfuO6gT/xBFZFxkJShLZTtjTa3QGc2fhLVyTL0cbMyggEfMwNXcpYsR7zAmdKZQ02hdu
IOKGZBC0XPzU+VmI71J4AmTZx0x7zf5yIxJ/FlkNvbD49/AW47RdOVCeGH5VOe6hCq8iP0Va2Dx1
Aosp5+7YmaUKxxWb/lmJ6MpeSjcM8FJgZDe5N/CPT+w4mGWdpuZjJc1thv6fvDWvdDbpa0JgPT9/
5nfhTTh0ZYy8sCakv5PqeJ2UZ+a8sPsMwVB1ArtsqaeR1H2lQ0Oo2eWQrrPQN9RqDpNITcVzKtsq
PkM2f4n5covCwv7nmr/wRYp648hPW2hbjVknyS2/EzMCp6PvPMSMP1oQ8IGrpczMWm3CCQBg7C9e
ti+YZQNEZN9dSrpFYPL0Z+S3fsY8SmiTpFqcuFdH9MD/SD98oZOqjMYtHFECo7+FHIP1sNM6Ejgz
QoduI1e3fkhoiF1p9DzvboOJKGcHATvdn6YcQDUMs9gS6xHsH25KEkhKv3ABR//YmqLEIh6vDaZa
627PyEahrNBcdHuxvt9MrfyjM+hPGHN+ck334AU8f6Hj+jk1itFxXzXQsEdBy8OupWLoBqVvv0fF
BbIwq99YPfkUn0m516YdxS8MOPt0m7qwjD84n1xrNXnq8zPp6/7G0fS7yTczPLxYkbAwAHS2U9nT
WCHxO3DS8TWDUzNeNAyZ4IoPxICEcMj8yubmtQWjMUXMWxBw5sDVgkF6/jhby6UxJhaYvIQl6Z2o
+b4V4asSrkyx7VcBRY4vZV1BV0sR7Tt5633+X3U7hCbJJ5gWj5ZTYjYynTaNUR/nErHw6t9Pcim7
xvhKPgLhMy64ff6iYbOsned4gs5nhM0d3fPHunn3mxN8fPmZaty9auEgUsdGS6RJ6d6JwaS2h3es
JI5170zdB/ORF+GF/sxqumTTLNadQ1uG0dsJl6GR1EXH6wXfbfB2/VCwzB39t4jzwakpTkppOzBO
pf3iliO7bNOJDXG2QmXSlZ5mXH7XtmUhX/EZ9L8bulCaN7hZih3w1hebGdC8C3JNRQuEak488eAN
ECJHbzL9HGyXiSIihuxGcapJPh0nydgC7K34liOkgPjBe7wUnCve4aJPzNbU1lWI5sDnK+0ZKl9K
BzSzyhLeNInH9eAkUo62wRqg1wUfoXv/fAXcue3SX3+UbbvbzLvYKaa56p2bMqf3t2OO3zo8m+CY
btpqsjJh7LBhnp5A/FzIemzRYXVXRyOlf8cJj0n3PgJ1eX1ej6Wl0Mf0YBy2ywQCKlG5dntP9IzH
1N85QV7vd1k56uvkaElBNa2AzBJKaZAVPFl+hom9LaPpJvk780+s0ECPaSZFVBh9ZX/hRoy1w9YB
HbxqfZH4jvVWE/Xyyl3IrbtrD7mbECvmgwQXqWBknR5NJhH9760ghajmbP/E+86R55NIH1o96hm2
04tp+3kaenTxUY0t+up+1P1XTkDd92uATkPhFjSzN6A7A8otoohe2sJwLIrG7TAphjeqtDGGSqKL
iG75W9oHFyJzLbWaGJCh+QyZ62k20g0r6vRee9R/6O8gEZrJMyAQdc22IG/xBptJTEMinr1m/57e
3bzmeEwJM+D8RLRXUN+mkDOepHGx+JDbdwgUDldPWEC6g0d/8DktTUvdS6aXm8vBtff0pGDBdheI
a+mLC+exX1PRJsOdZMmAffZF6SCxPxbE3rpU9uPMuvFKJ8aOMFfLyKQEOUjEYT+lfQxh7FiV13P+
oJ4boq0PfiMZvqxZroV9HynDYbBsX6BUySdGTi0SYnVtU2uOcy3ughOUMoMYunyAYuLF741ikHZ/
ijn7nj3+XwKdbaXtm3s0YFcfb1OZ9tbuS3cypDJ2MUPRmHvm9jprI1wLEGDOt5BsFpGu9DURAb8Z
E4Y+s/Fm7EOl32Dmk7rLwlZfJACN+Wlg5kBxHcPl9hKtlTOOHjojd5APBmTr2pezf8OBdm+m2hie
lVecY0I3FbQ2OKBTyKBfLSs1su3nu8+cOikUmsSjgExpOSSu8kn7HvTAdRYpsygcEC+zjgw3UuKl
vjvx5bZd5S1daBKJpM4GP9hZZqW/ZMOO6xESoABcOFW7HIPbbNz81BsAtON/nytXysMW1w06Jui6
V/oaJHV10BZ1vgLMFZXLTZ2Xtmqm9Kbiv979l8QR/R0V+moRduxgQQhLZFlFPDaiUediXoq4Nb1w
emiHcWpbi5KiLQfrObm7Jo6aOdJWTnUxazjZm0ZzheTKPqEy1nEpg49ZWXhzp43isHejdNEyWQ6T
GwO03BN7s3wb2HXVtRPcfqak7z/z/e7jLHaDvir15nTO4SSuebLo3gzdKnlyhHqk6Ls66AAfsBN4
Jb4czygLMnYPuKh+R2IAMWFb+GAlhXWR8bvMAiSwBWwRjZRbmkozfMpeHEMzb2EiX/S+WLEqYIik
Lb08MZrOw+V9GBlXAiPf7e9HUgd8Eaqy9FBTEmWq+6dQqDs2x16G7HWC+KaGwsZdzcnrgOrW/6Td
wDgae7Pfv0QWPRDW7mRdin09tNKCDYZtTkqdKMFbfNiSTe44in7a9uET/O5LUT81Em7H+Q8dczYd
NEmMjBS/qUSt5TPxAWFUtlOUm4t/dB/X+AnB8RIUAFKC4gu+apDl4Ht6VmX70E/xC6iWVlAOUX2s
vXHMws3keFYYlgcRatPRKSLTuqGu/PoLOfEGDWs4JG75ovNUk2ukgfnMHFpc2eAhZmZOBReFXhxi
+SAL/WVFfD0QzjE2vqKV+3zIsRpATXC04awwOQX3OYTUEB+wKBsVc4v3OtmOPUDLxSAbWhMZrCMl
7zHW/Nb2PJAehiuRMDK4VJHyeNtF92yrij8Ldx0OUefilyhQkiU0zA/BuH+Buh0RkViYO2IDTR3c
AlyBXEdqdqlHhg94FSTzXCh+tf49Wv81UIieRDPpMWlus5bOiBAPcla3iVCubgbjeI65UFF42Kiw
ZA9LEje9pPLSMnT5Sa0//8kB4q23YXKtZ+pipVR7ax1s5Fr/oE0PeSfO9Y3rgfhdHAb0ZCwSexOh
ehH055eAuwixDECfryHUgetPGnPn9NkiHLKTh7LbMQ8bceLf8qDHTGxnrcNTs7bVJyOXD9L7noKi
vLHODmxx9I8b0Cq1rlaisvdSHCdPu2vK4HEXKBWAfYuZ3NVLrcWa82mWiGLwwFrrIPHnG93ez2pC
TEbW5t+xYu3c+rqvCn5tJMmsCN5owg6+0oahrrLWpgeGXN4+XR0+SdVnzT+O5A9oYFjVN92dTIj8
mnc/jN5YbDn7OGOGCDJG3wLDkk+H3wIjQSL1zo9SoDw0LxjLIPybVFMgBNaOktvEZlSAi9MpMTRB
g0kRMuCXs/4BKZljvtL1yhdW32UaDi8bMcis/V5c4WKW0DnUtgQ1iaU5Ot/2+VQz9TsQdCjm0uL5
X4Qm8cY9y1Ks6EDyV0OVdQo4mMpCCeYCn/Nmzd66dxUvlSaCkjFwiPcxGikuvFzIg1dOFsYm+6RO
hSnsStmGgIFpA2AY4LOLal3REpgb19FhZI63b1Lrtt90RqgqphqUjVhc3SKiFjbj3WElyWQEu/5G
RD2rwogfUUQF05Xqp+bDRsQIJj+gJdfziIr+8cywhU2bTy/VgMKH92FKhLAHRtFtCh7157xgtRCi
O2qDpCcgMVtc6LtKe7ZaLeMyu1dFSwiIpbKXU3q6KdFD60TbbkbFYnKX703waM+EN/uwUHWO4//E
G8NjhrlN1zMHXY8KKcA1hLN/I62kjb9UcnFwY3uc638NL2DuJf9Nxf9pdAMipw2G4KM7uw9YQBXa
JDjgywTtC6mHsAEddh84hPWCXDlbDJLDiEYGKbsvy1crhHhe3ATglu2UwoUDbEqJbDN6yIxSGWWH
g6IsO+cUW/AAQrMqmbS5UTIwcxygEEQlwPrmU7QdT6XqY+JNAlzKTzEmXqxPPDQg7OpsnB4v4ISd
EgCQRB0x6M29tCMqZtPzZE7+SfwrDuy9k//gHouoZm5399nGzX46mk9/u5qukBy0jwy5kNQhqjDC
yhzFgcKAWFXHiTstfq08kJ+iZbFOjVUSoiz9OmPwC6RZf+lPOJ9JDyYdRZUqrwFqmiuuFbdCf/WS
9KZR/+37ZAExf3wjlM631MuAsxbE7Qgw6FresYGk0bnwdmTVd9C+qBsaR9vPohgrD8Hs/UvMNbgO
cxwNO2hYSYjwWIDUH1n8T7chKevLBsuVDoE/lS1C4g9OdOZfmjmfYbPyUPGqCzZj82v53WzknbX9
W6SPwscFQrtuVJWgUYoJ5zu/4sbp+umel+p0S6yCiV+IZy7jQwdkT+hlMuHA95aI6EDcQAOkp+81
FWbJU/KonxXzwt/gg7p0XJfLGI3P5YIQJDvbfAiCIy01bm3r/rvu1JSrkXYUUyC+mWHFn5NDEyZQ
Q5TPXKIeRUZ6tp+Wg9HNkApyC6Bae2mks3qJFaYFhSLAzP5F03FywvZi5l9OBU+U/MUdS+Un5pVr
du0ZMQp8ceUi3XZ5rn4o69aaOjwlu/A/vo5mUoclotTVmxIRMeEKwH23YyPRwXl6+37um+xQPEOV
6ZLrqJL58otdemjzH/rVEXqMMlLJe8u11RCH96Qb1NpJWlRTo60ftXmoL5H1MSWs81hRaS5TAMxI
Ebnjm5suxSOwi9aoPcIv0wyjsROy6ACCp0lww1vlgcuiVqXE/hdb3hAL42ZiBiNeWk33M0LpjF6q
iO2WiRsMmuyPVOMmUD8Bgsat3e79jw6lDnR5C/8mhXfm0/Oj5hKenR27MQ3GACKt9/xmR3wlmnRO
wjWo8xaHteqd/Mf8TvgdfdFuvnyh8T+qWEanFNxmCZ4eD+kxeht2jsfHQBWTrTNLIOI7lN1VBIzB
QfYBDY41lpnGqAJ2026COpuaKcXB+ueShP07IgqVEin0SKrY+Feli80UIKv4gGlOJZkhHHF5aGBo
cvX96/P8ZXNPHJXmwKlCUt7hI4ckziUYVhxn42EpfM6wVrCManfv7hB6PnqtiP/BkWHxBkqppYM/
dcLmjekPrkecP+t8rjpkAoEg18g/b5HPeC2f14m4wY4M+7FHCJ4vWJQANSM19Y75n/mw1pqd7RbE
BR4bNvnubGIBXr+V/CXnux0sTn18wBHFG6SICf9j2uop6ZIwPVlcIstdM1ivNq1mJsHdEJHHNC5a
gVUO1mc/M1KYB1GdUqWPvheJ7mxw3xx4cJJ5eSk2Q7aAlPng8EWKiGU8rMQLL5bRtDxWqCf7erMa
5gf0AlJae/Yyh59Xw0kxkSiphLkoXXVGQTUjy5duYy03924jO4E4tXJyS9QXF7kRU5ytTWvsN/xu
sYNNVcU2ltXd6SKAn84vmBQ90YsD7qWeQXysES63DgwbVt7+MpqxnJvn/mfvHlETF29cW0bXe4fX
UAS9MP5jIEvnaD7qp/kxXiCwTDEfstML2YFkofkby+20RtWEKwEp/YUGjHlEUPuBl7sTujG2EMeI
RG30kH2QYc/EjGeOIF1yIRt8r/Vf3Ka5lVWRCdGEKy6q9jRZAebWUW8EsshrC3WO0+4bcHzK7HxO
FYvI6dTPE6isSee6zYum+BzUeAnvPCNtgaKqpEqetl9YXlEylHmAwS27qqNLvi4/v0kWEPhyPvfJ
h/OdCuQk8y2C3gBfd7RLmtUfgIpdJ+bxaNZySdQe4yJxkXELc4DD62VlkUcgtyrNZAcWEwuvx476
iuPaJpfoQj65/xNW/eR+PP4JWhoeZCOybAZ3Ayf4mitIU0XfWW2EJh0ePsHAJrlAV6Dzf2p4Yfx8
KVbIpxHs94zniJhf9Z1sOjVC+/eXrj3U4qL/DUdDc26lhf16uTzwYVTuHnGXbQoD8xDD1YLrrUhU
bqpTtgIzFQbAap77SI25ygIzOQ+xbgx3gwyTTk4lZJ7ffDh9lWTNex5GImA27Gk7ulDvVikWMhgq
YwZjvXUZ97VUNm1lAd7Ar7yoBMLun0oAIuTfu97cG8PEfSYXM+Y/NVOTFoJkOPIfJNnjj/uoZ0f2
K6tGIsZKNx2BH8lg9/DiD4tftgdeqKBdnXLIle+GnDkZZU56UPQ0LIfQCWKUKs7GHdpeuOx3el76
gqLnSppgOsl3g4apVY2WGhss90hhVY9U93nIe/iQwwfnHAzKeuK+ekULvs8wX+vok0WyLN/fTkO9
dX5P4Aph15MFNn9BY8iV3jut6tmVkWe+uvgc4JcCB8vi4uswM+8MCF7d27XTcqawMHx/Fkv7oOfo
tyYHemQt/L7icizsKMJbsQ0wrnVmPRMK0rX1SBPlXM6MHFwe2qTVDLQJDscu0xYrUGrWSLUDrL26
VjacM3v0NRfhH4/isw7CV+JUABOFaLOookuX5RLHKQdl0L1Gk+Fi8B6twdGPQm0P135WjnZZTwvo
8UbPIQfOkvcnBXVEc/rjFpDEZ5HCVSKZePJ6vQC4r5LMvCG5CxkB5h10+7pFa8t5A9wENOHEJ7XO
3X7DudZQgKbYKswFFEiFZP2uv1gvFqiNHqujyZ7n3+NGwp3QUHki8J8UMAUTqhnLxZYBRQRlvBDm
iaZsJgFvGEFXXvcggKVPuNCesqCNPFV/g20M3RxfaXXtgjjZMyPlwaM2udP2XhNS7o0vw0V1Jveo
cUpuPejFYgaEQqirdl9iFm9/keXTky4pBgOnCtHq2ygWonXqBXCbD9c8PMO+RkbxoDjkhEprRCFs
l1t9yur9pgl0NPc7Qh7DooJ1JMzMfKI9khllkTF+YbMIlGyePjbYCo8vsFsQpzwaDwfXXzBKOWAW
cu3K7bTT6yuMViuF6kO4CH6kuliFwTvs7IXF5liMXUgvVGiVygsJAnKulCSL/3SPUeV5e3guNqVK
73ZzIMHLM5/1Nfy0wpjXsU/WCg5AxhEdUy0CiZz4UXqlYxGICQkxOY1lRwD8RUDIEENEJtd9n9p5
mbJEkFvw8LudYV/F2dWDCFlIR+kI6DU7zHBh8VgNw4Q/MQd+CvvZNSXAHdAdUP3xYs4p/MR3/yhi
grr1zhpOSlnDwc0b9bPMWsLu/QlVcyggU2ClmW0twe2Gy5VOKFMj6qf2rXjeh7NNU1/HYqaMKqyW
c5/l+JGE56JM7I7qoS/X+qkNpIvAlcbsGbpGOPdcMw2QOHE8QgP3r/MqU0YF3s5+vhtsjjqf5Rak
EcTYtdE135CCMJgYp3mVnJS8gvTjdL8HIyWLudV4wl+AipzynRToxuUM1SO4S3J5jcGDMwjZW2qg
kUvrgJrEsP99Y8GtzIhipLz31CpiI7y3bVWWRs4BhLtiVoG84WCjRVaaj+T+l5CmDBpKIvonHxVD
XYqA92z0j05PEzRAofbcPi7yw76Cz8Y0G2dS0TZnYOgrqDhAPtNlX00itw2zqqp1+0HWMQLuagP/
LBJhl/oUE34G4pvGFWMTu70cZM7BityEMZt+kai9tBUrE/TD82q729jFbmq2iWfghPPWxbEbttRo
p8iicoh26gKGnTWa2KPJkruuSpMlx0BZ4lHo2Z6kx8arC2yavApJl6i2buxPVjKkbg9WEvlwvuWQ
nY8CXnIT3CjNQShe4T+hrSybEQTIMSHyu2jcKihRt+Ur3VV2q0oD62ocskJZYKfs4duDVjrXGWuF
LYe6WF41+4S1lga4B1CtSPX+v6Nh5cbNxbQtrIzKPyZgTdB5QngNtk3gzikgTLAUbkiZLgfk0v9E
9ri1vbtqG60dGTC5xw5eTYxZKo62u0xurzw8pw+xFEDRLznJACYjuVhjz4WDnjVUtozd5cItXhrt
E/GsbfDJFACjZ0div9Ld5ZGWmwFeeDj9CwiZDXEMnPYHGlnKAmtzPT1uneXhd4UkNq36XAQBFfu2
EmKRNOO/pl/PFBX+w1I60YiB1Ve1tAN7WI5/8smlwX5XUlmj2PlkcJekVd07AL83PZqkksxhfNkQ
lC7NXzqhLKbN/UrXmVhsP37g7nRjMl6lHDlvOmmxA7eAIi4mH0xZr6iVSXP30oSoVKPR5H+CAJo2
zYHg/2xKnfa0VfzncSq0YjMAcNl2B67JTxzwEVyMDxfCwkKkC+ynpAJngeZyuiEuVfU4CkmP/k7G
l4vkXs4MXeKIT7ClETeQ9r/7nJCLHbEk8bgfj5GgeX02u2JGmSfft7XA4ra1RCWLDBcF+3VLByJ0
TVA3PpUOd0ADMlCG/ysx2e5hg7HOCT0XYsKtEhd1k6cY/IjwwZ1YB+iwDDB9u5JRLAJE7+g3w80d
YHbiwFdBhCSrKa1HRg4rGtedKptwFCFGvc8oYwR/2wftiPZlP/Onud4Fl7ydmo6bCU/BHGsOJNh2
GM2WvhcdHXgWWl77j8J680FBynEi69sW4e5GcmW9ENxd6yW51w9gr6EBKn1UugHrWiCoNgP7iTGl
6eKHnF2JkSQYJHYPxuW8xQoMA6ZK/C+6aFZ9rnsyLtUYQ5hJetbIrcjQ76b/9euUYOIW8L/S070r
+T0fvEWiHUG0sM6pi+HL0Un+FYtEJQxjKdTQLkyxOwE3wRAEI6l88ORYr2+g8aHVDDEEInFLHSxW
2KrUnBwQBe3Djo0x0qQ9a9wpF7I0ZP2KPw7woD5iULl50sBelCgPAlmkOsDOL3+KGOE2ScL/ghpe
19cnFB5g8QaG9EV+bgDpp3JIH+zi/mlkHthEPaQ2GyG0obzQE9zQDcVPBVjXUkPzGSMkr1cgMEJA
XCDFgBgac7c4Qvld3kL1WIUdTsWGOZdIIkNZqmltJsqbVxmHYLABPtQSgBZRNraiYTCyQPRQYYuh
f5lUbmSivB2IOUKwYBf6fDyHJ7Jr/96VO1H4gf1Z+q3Y/i+h4dsHAzdM0cIeXKMdit4r7fv6p3+7
5NreCOkRD6FdZRCvPtQNXY+J3ricVhgMcJO/QCmYuCdc4LW5tpS22Afn0/R/FHNmkpwcAdsrwe48
RcPk9B7A5h3MW6dCosYkNCfkUBLkreq5X/n31V1oVrdGLhF0sfh7g82C8A8JV8fxxNdJj3qL5sAy
SqLHY4KL7OHk/kH7R6Lof6aKbIL+X4OjMb45v4wCBDgcj4O+PCw3A+9phL5gDHyFXs/EAjgFCqJU
ARHIyrGghXio2ajW99PPC0Kg5F0KUPhgp+GWentev4zpzXKyHbFAbgToBlxnJDfiB5y+znxUuAZH
6KjXlMtg1mvu/EDwfB1tCmqJXMJaGzWEM7hdeNYQMrnihC0zToaq+sfNhEjqRO+7MZLCwalq64Eo
xX2ELBA+A9HfTJRTpsdKrn60ItUh29bs1bWm2bYxRz9Abucr3q/ompb9IrBEeUwGH1ccmxZLe60q
0L/AEzbI+Y6y7tc7t0hrwFG4Pr6ag+ZaoSubEufQG2RJIwxLD6xb+yVqq5P3SlkW6UnVvwzgD/ia
OMUh1v2zFzJ5h2JsBUJA1LiPsbaJczRJCyHFoWENj1CnvrXNNtAl2f07ddNxSiWOPjbnqHl6FAyG
3cVHqQ88PgTsthiLfYfCtJiyfmb0jd04DqH8ZXAeN/ONGnJFGE4ZP0jpzjLeQrVVUGSmsEM7xIM3
/XqNQwFiS/rZa9/3/ogiOC9YyXCsFojQ44nThwB0YmO06DtLwyFh4eW16RANN0YHkKi6gnbj/Uw5
DxJQGYR/Sx7RPe0U/bx+iT+RoJCaMYGA2O6h+eqF6sdiKvkQT7jXtSZXrMImtiF0xE//55oaYG0K
5nZFhoiMER5uE+YBhwhLlp12UpZ1bvK88PidN8UpAVDTBjLoT9RZ4/keTOkyBH7mqMsSt0QgHgSA
wRr2AymhloZXsX05zYKBt9EXOZwwAJdiyLt+2ZLYPa+Tk2TmGlXIPysOCAzOTBBdm2Hwiym/w8sJ
6yOy0XtLTXFML29yl5sp7VgI3Y9jHyHd0dn8+PTwbxyaPnX2DpJv3/FlxmKsdTMqvEYDqCFVgAEl
DL4FQ3wz/jQVQUH8BkEXCgJd5QU2QW8vkIcjJ+3kDU8BlQwrNNy2yLkwWH3xHzV9Y98IQbxL5QIb
h6nE0YNCQ+aqc+QxW2JJE58rgLTbXlx5Ruf5Hh0DqjO4UXxys7ymM50B0byI0OqwO/+Yic5j62t0
4DP13QUluYzA5jibt+boEzhBOZJG40uAyvdmfbv9DMHzb6ow3QG9pBhFus/8ZPpyCVgV5E4bZ5du
DJqz2l9u1ZSfCM1M8RXbJYhMKHe7DGvdmjxUm2Wkkch1k+g71TXSyct7kIMW3zA3Ek0i3I2Wdu0h
eChGqiBOnwQfJbWmnrcyTJ79F01TtgxXqhI607HUG7bt08KzPMlRE1etrlWB14PoDaPGKbEFKFvQ
IE5x6flVbc63EpSK99pFdwLGBgjVyQq3iKe+YvVn4PeOh34L95fkJVsvcyRAsxgVVcdn4bdtfyDj
1opN5DS2HdNAknrQjIKMsqfJ75MIKt9uXzyohjyy/FanIb4dDITeePHMl5b2ys2z/brvqEEQi7rN
kCP3ck8JZQR+qM5/NYYIOYCWVTLJNanIlfvYjzTyX3N1oMLAcQKTzx4En6mPbqJN2zxmlud+d1d6
Api20lz+eR0Bg7mKCzTIcacX22cO9Uhq6H85p+GjvmcFGCUZefX7BbqHGlZfiIjhZ2IdU9XIc4DL
tPhO0d6Ts8Q2/XDLvFk0ELyY8Nue0eneWFhFE5M3EzoIPiFw67LB5V+EEgrz7W1gZ1srz2o5p7un
rUgu2i1aYlYpnBwMxvkj/n1oOtguhZ4RoX7iZG4ubS9ja0/TQMqxgJWExtDFWYwkDLM/y4IQ0ydZ
6nAQfgMJr5qVD2P/Zpg4o9XYpjgT+zPKijXYXNenRVCmB3tvVCo6q1CIXB/x4RVytq1tiLqAoxmO
gYCvcHp5M01Kt6LkYk5W7SuQQgVJK8VNRuPhdt41sU1S80OLLzg9t3slxscrzX72DXLVxU9sN9kV
P2dIPsFryCq1FRAjklhoGYvJrtlO8ZBkpuiW6r8Ax1ZNhsr+4Y39bpo0iK4rFSX7gBisLbeLMIFs
qPCYD/UyjrZCK6qyUrH2TLCUM9/udGyigyE9GUgtuM0RTMT+A7oqZwTUbMC8zcnUdQox7ez7VK3A
HdAhArzvRppfk2hDUegGkiGKMUW4f665+q7iOpg19Xq2tAhfmqfAWjcRtv2NsBdlMDAblOlbydqI
7afAgGPtdpEgIz8a1au/+fzbwpMN+BY7O2clIXbXUcqGx3N9KjiREKHhjSBwPeFZ0L4CTVNA+6BW
4opvHc5ycIXnufdfCvGA/ohQMn8Yu7RTqfGcrxgninRf/GpeulO1lH4e9CwO1LzLsRnipT6qU8nR
hQ1KnPDUhsp0QhQXB8tt+lzyueFJTisOrpahMYSv2U4j2Gu5NwiHZy8JSeomV8u5TF4kzoyNSve6
27d68Vfg2x7IBoV0lCBoJ98iY8nksIaq1X5PAmP0/8rm1dwSCXsBf73HgsMes73IH6M+X55zJdqY
0wIGE6USIs1RW7tEGVQuocUC7TGeyk5hde3Ix4GBzZqsmLujmPnoeMNFyRvqOVSxAaT6zjPXAv/e
Ws2vZ8Y8SngKFq3MYImGvInx55NdEWrRmy52TnKXWozGvw1atkZT5Xb/yVvq4w+4GFNUKK5JmrTu
QQI1JpCn4aW4IqJuTbI+xb81Ojx/EM//7YZA78bIJKB5XpkoCDWrfhW3dFrHjJd3p1qTG2j/ZTXq
TiBgHXT+E508/FkYWYINJf7pmaQCO4FTJVUi39x+yYXNUcx8mhVUSO4k4oT9ww7jOZF0O5avN0cg
CRwKQA2HH68Qv8LYuiy9VcMbXsqhmrqvAUWwsQwdR19dGZ3rJFIt6gQW873OJUsIQezHueRZ6UKn
NDGy6aVt1brHkr1bAuBkduw8IXOauuP3Kd65fWRM7DI8N+/p6ed6lof38uuFbf8pYJCOC/Tp449k
dE56kCec6Wdx+WjkFAZWPF2MuhwUrfk7Dz3PatGr1ag7vVnOT5f8yXJGcG90PqUOhc+zkSmNQ3iv
9JQD64d27ONBvizK9+T/yplasMxnnWeI7CzxMz8LyfnIayQjColfYCKZVAoQZ1uD4lHJqPdVpTtg
dabCYiVVt55S3JgCEkB1IrP63hcAn+xCaDm/dHCkZyddiWKvLmXqQ3uHd1W/HWc98G91Tc5iNZQi
1jO7F39Waf+pmWYIphYq4KkpvFNxHhzYsFlgc09vR3S0hyZTgyEd+ZOCD8NvJQzmQC05e96vgYkx
wF0HiPy6s+HnwFc93TWZmqLuzsRiFEZ4bBHPNcifc+83b9+quIIUxCP2xm9JJ8OuxUp4vQXNgwhL
txoIHs/Nsbeaf5hxLNiuYlm3vginIP0t2ue775wy7DfuEx1ffqN9GhSi+TnaiMuAWKNwd7677xkI
/G66tB/fvmsi5ymyQspqu8BVL/+y4yLzFeo5FuH2sWG7QP6ArKXRXLP0FKaytQ9AssIyLXcy7TZr
fvTNMDhpb/0ngKJi+pOChPkpnERXhSdmFhh1GprdwhmWdKlIOzPljIo3w8EzqoMZLI2djV8iebDR
Rr3+iz3Z+tpEQaNq9kfkrd1+yQyvgSQsxymHqB3JcC71ALdLNgZn7Eh5b44Rk1akSiVnbPM/kjy4
qv/CdKA+mgWfg3QC9OP+8KNtszCNYhQJZKWHCc/2bHF617IMwtePrMx2bBVNAuR2IdOiYlh1zhIm
wnx67MNeZWg9vVw5rodmY0MF4QtRG+L3g/+vxAi1y3bRj5Jmu2NlsYTHigYhKij9Yatuta009aol
oEWEWg9y5OsfdGHiPGVm5Wj9yuov3V926GjKwuagUjCFnEPrcVZ1KfwECC7n5nFHNC4pyaq1B7M8
dn2LvpNS2r4/geJGDoBKDF0AXbfv2cd+KrTxbxcbGx0CIccLTJZmyBiWaCoX93ODM6I/nbqP9CkG
vV+lTgAAkda/9iabIMvPfHGNhhLL5TsekeNYOnSzZtKy3kP7QmPSXopTy3w65Y5w7KpgeWVVqUSG
iXetyjjy7PuYH1DECu5QhLasqEPHDh7ASXuUbemWehhTaFPyUbqjAB79ISL/7rtCYrHdjtew1JQH
TWQ24TJtM/J7DcWMPiqnPbPZ/yLUuqPbtHozRIuUFkh0FgpzjiFwsvQ6rsjRis//RILvzkQKa6uH
IfCgqLVdKLDDILgaQD0KEI5tdatpMiu2gwnXOG2alm1tf16dPt4c3d3BjE8JlAZl79/ViXXjGbEm
0Ge/tZ/t9yRTuyxWDtCTdAC+a6wDKYcO0T6DdK0gRjXWHAhJ2BwJOCl7n4tMKF/OrQQRPynqVAwd
TYk6JDFdMiR2xMKlaDq4AzXSgMAqFYWHiBrrmF7xYIx+dl0QKnVqUbHh+HRaCvClQPO+MXwqVY0g
oTMM8MzGTQ/7uEWJSxCn+4GxMtuYOpawmRXzlpGvctR6ilRhas0TnQYoBiBsVDVp0Qx5eFbEkp7A
DXap/5AS8v4bQSWQINT/klbEQv4e0wO177R/gV7FA+B/1nHrFlfAtZ2K61j+EFWRG7hp4UyoXygf
S2ySeDBvxQu72sLDoJaF7cNq65b49DJ6T9kxeB58JPpfhXKyitIYqlDPoGCvxDN1BJq/qVOTEEu9
UUp0uLpQ5qxBr8aLRj0hSwBBN9Z4qLxZAXAo3Q/E3ApaMUfCGdr57Hswtf0QWioBiBZd+S5PdFQa
6Y5mm17Z3U3oK6jYFDXkz5P+Mi3d76pXYv+PTxI38m7Q/z3juteJH34A1uaT/nB/ioPGCgBIIkI4
1cmlDNgfwfxzBA/SG4F6TedLCfyKaznagyw7ob2RjiB+y/niBUt8fZitMZApzXDvOIoGqTJxrzL3
QbmAdagAPg30g2SXSgAJwi2u8jW92JSmKWIxN+PGjYOXvYbJF/y1i6QgVkWRMokWesEnPBwKlJry
nuYtKsSkillDbuHPp8Od512Kvt+IRh2VcYVXroLoQ/MiGey1F8MY0JY1U9IN2fSLeEyMZeLLd/bu
l8iBDeJQTm5bp25oNWp4EQSEYcn972qPPMuPML0aR3g0MeNw7uaAdPm6zZBbC/kl9RxAh2GQD/2+
Vvc0YIEkzB7Opry/8RMacdowLck4BdjVmcl+znSgeLWJNBGPyGKEmhjPMVZvDBPRrltqX5/ewg88
bnuktFJSn3MYdIXsrl9+6FgTR8VIjaqoYn6jrWEQoWp7ZlJ3M6eJZ5Y6O8JkoZPXiGaEmFUiVfRX
utyYUEkcuWyV6bjccr4NE1fdhdVTTHXv1MpLLcfIO0W8KR3mTjpXwhwOdGiMYybs6UtPpr9YN79S
Yw+JiisONX7eb3Hr8PL1VQqj+/wCUx3GHtNCFofpvq8wxgf/V37yTZJSeiArGcqDP1x0uNSo4Gn8
9+KWhN3kZpkg585Cf7fHXtWCcesMCiHlxbpcpRPqAK1RC0uDrngGC0BvEKWG/PK11s8WQhPwSX+G
5v91iDczFRpPfqxIEA976rQcICjN6O2pVxdFRNA+XsCTd2c1nAHs8ul6R2yn4W+haMtAP6dfc31i
l5H2j3MYvYeN1buemXbleK/49MFjnpsrPCpJNfN7gkvRHc+M7mRCe8YmobNIbcolLF+sCpuH6he0
apfzxDyqGdSwFAqz13+n0RisrPCRSS3Ns3Nzu1LMV60Ti9uXw8a6zIDtqu4knKQBLjbnytm4QXxQ
NHO/31gSs8JwA+VHIYltSnId1j9hAV5wrUWVSLUJRCroJEalW4QxIUojLz8Qbr8DpopN4pld62MI
J55PkoD2pq0Zv0PToEPaIs70bExwI/wKYn1KA7ttkidX7HZXAZbzL3RClWBd0p4CEjsjl/D96f2a
RgbYLKaGc97783rNxdKcT8sL3FKlWeC6+EoKUVEnYOxyc+ALCljomRs9kY7KY1d3gR2M5xCH+elF
cbnYM70u0gNSpNTPyUp/A3oFGXsl9/fl4qoU7BUYmqJyfoSBEYqAcN3WB0YL02L6Zxc1baC3D9v5
Gfn6rkGzrJ4IMyXFR5zoOu03Ra/29bFDtw+UhTt2y22qVe4MuZEKTCz7s0LbgQMyk2G6YLHvO4m7
lnxFed2XOdB5FP+dA9HyggsU8QhyLR3rAaS6pjNpKhamL7EVzTb55t5bffkRwOW8jxYqgOI4REN/
sIEVk12gZT0UtkXAYlsA98e/dINkw/ExTsIvkDyl3DRYjOi+g12jYfbxT2j+R7Nj3fFd0TBoUSie
RQJjoeG9b/z61FICr8bRfuxeIyHMY1qC+HlaMEXpWPfX+GVH4bHpJeZXuv3gh06Ou03qvcS17WB6
wjaImJotzoltUNq9F5pHQR77arKbShiULEg0XIJlgpuT4nQZI5uMFOCvv4wxJuPMU+C3v4TZbD+L
EiGFNbY9tMOF6FFFz+n6F14vly1Z7er/aKls2OFvbJxE0OQj7q4cLB/fH22+nw10fWdjiYYGO44+
tq38WLn07NLZfCsvqZ3OuTlueG9sA337ikSCs52cXyUWCGGtymWSVBBFt5XQ0D9xFNfAPpiQDPKm
CFUjaFoYMjoBc2tCwRny/OdDipY7x3bSXzx7cUdGaW6hC+9g2OIo3XNDaM11Dh+q0lggI9rlBZQb
/aLizFgH+p23e03PI4c12seMtzUrPRp5ttWSnDwwk5vAvKYXMsHFHgdVasHLTQA2h3hvYNhUqJ9Z
1Blzv2Tb23ecTKPsXMfZQllOnPIJyISHhyle2A/0v6w/JtxYr+YtR79tYVA8ZLQyBrqQc/WXE0x9
9RMlhg5oE9YM67OdOKFD6yIlCuxIDcRq1d8Q8kL/CZxoquKyMFxUmIwnB5jZn1Bno3r+ybsbfDY1
58fP/lYAyXcyhTKBI4qtKquTxdsuvRhmlfxEyrJ2E08bWZkZB+jjalNqbZ8idC/FSZ9ydG0lBFYF
WoSRDdkP1cy5JsnzTC+PhrBE4zm1gDqHnRmJkawZSrs1ZJSkwYBmN/zXfVpTD9P+UMn2fjUrDAcn
gEPaAVcpPd/8UjbmHAiD2fwfl12ApZzLOSQM3EHGUd2Dgl3CGx178XnrNXZZd31fWyikhLh38aOq
5A+hR2hrY6vRZQrGjQhAylvn5lxkNY4GpyftGflI6ZjGtXUUl2Wpq8HMF9h7jG1QdVYXJ2qt7wvD
8xxIYklBlYxvs6jf5uPlmcugQZYrff9gzZZSheqpNEOQYitkOzTLH7FGtn8hIQX2fAbPqjKuJi4k
bfCmetqbLPzIJ0rtrn3zi4yiN+xPYJmcnnU4ZQ59yjCKE42hJA0l2rqgrDOcjQOkdm2keWHZW+Pw
+EJqCr61u/XZ/9NYcuj0Aq47S68xz9A92zjiDA3skrqjhBY6MVaKKOrwfOXQzvpijv9Uz8U58EFS
ddOw+RKvWPNM/bOYd63IeJPH0nQtIA/095xzRUuJqF0LZP6atgKC8sBdEcmycj2BM/C0uI3aJYeI
2J6GukkBt2dhc3BzDjcxMXKnI6SnG2zTh0AudTQC8kjNo4ZOt3OP1FacdAjF0KLFBhkf44HQqMJS
UlaK6Pva4FMofZ/0FEUA2VdqLQ3d6FZDK8UqmLL9tWM/csq6rV6sRO4HZgujS3GpgcdIn92lwpzr
5npxNBY2rzGtrOWgy0/M9m74T5TZ83LboBjBlgPNpuHhSGfiH8n1WfSU58HFpspbkBv1LsdosscZ
q6lBDbQXT4Qmro/9jkNvTUWkeccU/LFaCQdnAxpnfSMGmQRarhGr6sQ8gFtQAsENLijNTBhdiNSG
BXLUn3fgcwAyi3pHPKkpNnCWixL/zx99gFpv+RDcxrXQafv2gMljYcKxPEjUGkyWdJj8Y0WKT1df
naa6JtTUF39cgiM5reWfCuTaku8BPzo+yaiQSI8AmpeJnQnewV9DZ3Kt+VWRbt/hoedAyv79YYqd
KZbZuZ2G5IFWHhIxq3kWxO1MJ4mFmWinaWW2moHtB02jUVjUWgB/RD4le29mBBqJxkB/UQMij+fU
GGWfyDhSwjozXbWqBOF0/VV3RYETijuGx4KGtxEsBQb9XlC7aj/+XDkeEi6Vj9Nivo8MH2QcDqtw
S8WXspBkfPX3ABvayB7qDLfv0rYjAiIdei9QWAjV3ymy2QKBY1qV2zhxuwPm3KT25/SFVbe9ghVd
QQgYn5Bg3aRGmbMcOIoqiLymVv4+95Urd//od07cPHa9TJLS33v0zolXK81MqgDHlnblD5OuGGnV
NR4ViEagfX2DKODbMhRDpH7O4gvxkT3xuPFSwID8YL5Aj99taKD3JoWcrMj7h3Tfe2+ctsni0tXK
lwfwXscb5EYm0TTQ2bimPAUwF3GvIDie0aqUgsbVKOz4RtfBmEkcb5EZdanWEig3wKX9MSe4Yjbk
It09Qv03i2lDylYUfJTcFxwZzFipqg+xz8okHdB/iC73S4P9mLCfFN1E4gvloyeWqPj+R3xJPzua
YN/nxJTc08KcYBxbAkVqI00yKQtMvZy1nxU4fAAXxKc3XM4RmYnHzo1XcFpXXJ9ooJxfHp6GEnD0
l0Rghg/LrFFNaQHACHkHgbJxKynxu+942RRS7AJ/gcjyaoGLKEjUrXUxSlntmxi4Yi7t72jFLION
tuf7nnRQSf0yeiI8N+AfXR2LpaLh2S47Y2W/OeXKuEhJHbrdRT+U9cfAJ2UP4dd6hYdRKvgd36Gs
kMmeW0O7YhzQDrBPmlS6IbtIRi2l/50xK7tVWqasSGb6zxkWGo4JYwZORzUSLG2mIDRbucQXdPPP
/MnVIsCaoYr2erdkbvYrlxp/XpprLrqV0/UG8aYiY5CkCojeYqVhQIchYD9mA9nHOul7QF/GS2pj
9+VpYHF1kc/oz0Lbxc4nH/9Q6xXo+j1iHer1PM9iPu7Q5T5ZS0ym14F9J5NHxJKzbiwxDfiaAXMh
vM/RRfBBSH+JCFk6+NWxF2LlJzm/3nmqtba+i07pWenQCULAa3i58T5L0w0Pj3l/L5aLJikq847Z
/vijTn8ceVL0FoM3MxZL+aUUyFbn7tKEi40e+/0WUN3T92FJsul+uZ8HFaEYn1MuKIoKp7OSqqQl
b5U9IyY22+YtmaiMgS4I0whvNc/VskSMikputTJWkthKKU+kbn++REjIBgJL7fV6m5UvxibZ2+v8
FUJB5HyOQ8zp01KFO5/Pt2hRO1c1RVIEkYiHdTvN11xh0G5lsKZ6lil36Fzes/Eh8225BIyJsiyp
0ZkS7An60O+4ozTMesthNjc9b4kTxAoAfkt8J19UKqdcu7Lk0ECEj7txbCjMDJ3jGItCPtfG8zkk
5+s1tOEeNJF+5WmcPno4hGqfXaDwBXYGMhOnGGpBrReLMaIfh1W5c13fH8Z4JZ5oA0bLHQL5cPgh
HDs4RvypWinygerYQV/cdwt0BsL2zRJpd909Ske82Jei4wsga3KzD10EnN9FVkoCgsrMK2lKdCfs
upIihodcHVLubPxuHzOvVpb7F6lVByQBgQU7MdV54k7o4Y6O840w692NCdmc49wU7JA+x0lOoEsK
uz+hIULzIEq26v0d4qwGIwae5kJRwOlzKUQJxTt1zsmVdLw9xCplsH56YFWRY+CMBvmcAMA2Wk0Z
KYORGm5CPFfoMB5qJC4+oDLH9IhdJJCqEk3gjafmNiaOdanAQmDVxKrHSK1yLHCdEQfjDYXozBVB
Az/OUVjL1ufaOvk2Fnt2O27yWJOZ4zsk1yYaPrABy08qEfdJ11fnjWsyn13+KRq/p0fbf3/nehTq
aKh7VatWH1ruN6HvmcCLwO9fpc9c+DyP4NgbeleHOK2jN9Ck9+gupPpcSkpdaVmLQUrLtXH4+b2G
OxAcCDr4mEOQSInh7m22RPbiaMHzCl96C46oR1j1Ix0rN6cqWYllqYHQN++RDUvtqEh51GiCBA/L
s8Ud4TqohoD802vpnFUZeP4pb+z6oBwKHLaePwkIkz8eC9EWPgZAMazFN6mSsLa8VkqH++J0QT4Q
VKqCm6JZl6NIxWh7VZwADIZ3Oyoi86dP4LHLlzucTEuRNVmF9Vd33xAWejZF3kEmlqPPUM57MrO4
wJX1bBXqdeofrN+E0SOX3PCEY2POL1K+0riL6G6z8Ckyd+NmgHmcZNoPZ8eVlhASrcpijulXv8zW
OH1pdho00o5LueLxCCtTqLoIPXVUpxfIWXeZpRCFCj4V8qKOjceeTYgWP/J8p92qYskosbJ/eKb/
6MAWwSaq+7+E35gieuLEZTutwoBn8T9C0K0izsjPrv56va+vaOvjwKYql7M/p/7QSC8iRGnvE05x
Iu5s1EdZqTheSeCF8F3NL5tHuFk5Q9WBRT5/l6lFkQyBIz/Qsd7zzS5eGTU2AbADDvEEqLth5nP/
fDVpR3h5SSy+M/vs8qe9UVIsD3YNJH/NrsXtdAZXm8zz2XexMp1tMts5y272lnq+jFrJpw5tuNLb
Dllc5CfDKODszmRuJqfWOuYpm9P8AUy6Cfe3kM/W6eo1b3mgM/pSMiBOxjbLB2meWNwGFAio6piH
JCyF/oB3r6TXJgD1ncmQ7QDhKgUHt/fshGyrxUOn1cDo6G5ZjkjMNsOJOEcg5op1khwRJDGZwRUC
KA0JQVIzSmMy4ppMIK2pbOxSRqAj0V/EQsPFQJgdnL0p9t7bFZN6Ei+HH7nC3Zk48th+nKylJhv/
s7JbNPdLL1mFTNS2SI0TkdVFm1BbtRNeXtnMzIFpyC4+u2abA+HcT7P24ODUVJiQGlhfWTtEz/Fq
pUgpi//LZ65RF+z9cqs3z5VdnDqALU04Y6SotneNJ19GcYoPxzPrxr8zNgetvkNlIm/c9uNHSUhH
usP9TyDqFWCMaXql7WqbiD8UDQkzK9qyM+CQvKqKde1E/OoFCO2Kj0u4v5iizI5nod24TNl6TUvX
8gB8rj4MY/FD4h7tAA/z+r87eRBj3l2bNVL1Fl8raDiB3OPcKOYulMDpgL9pMM6A2X4qvXiB6+2h
HSbaTct22i22/zhvjBRZSOugy8NbBqIydWGlpkpe9jcYxxrfooZzGhssZztaa2Hv8YMN26ovE/yU
06SP6fk9ztsmlml7tg4oyKwI5/k9s56ceqKVwC33HnDI8bsnZ3vsxgMmcjLMpHvlQSd1O/hdkfU4
1KuvmN0o/6T02rRJyIOY/DBslQ+rNqtEpVyFXfeeQcJRiTeGUcej0/c7doo5aD7Xtr6Et3CLrSC5
Sxq/aTDXI/qW7ju+W5LrTw4NDoslYJBUk3dNhueMX06zCcXTr71jMUZTz5PTk26Xx/FY9AW6/8+n
qKDgImRKrUF0PTDSDBT2ihsulXEZvf/50+SZHfc4I2B81X43t7mkDQKnwDICYkhD0BqT/KZuJbRT
gd0u1DfPQfqg7LVVDU4s2pKgl2RCYagefbcXCY6S7NozFLRQXMbacKrJSFgyT/t6osVDV1rAzRaO
mFTRYz1vwkGyymOfvLdaeT2I0ujdc4U2ub7/Ylg15QPVFcKVMumzoY/Qbo7TgVHJ6STz42LGqTAi
mrfafV0tK5flFVmKMo9PCCDmQhhCzLl+iZ9pqUkdouljAK5uuRomCaBa0Tyk502+vxc8VNDWBBst
S7My+rMR0dPXpOZiKc5hVVLn/lq9w0Mn0+Bi/ZsjqBRi6TgraYok/KpBHNnvt5UagN8OAaygkOp+
6Y1CpH2byiRSiI1gUzSQAet39qfevm7c3Hh3hZIXEFl8GVzW/wN7gyeJCG6pOW0p0towTjOrrkX+
JRNWdPLwhKtLMOn7N5PqowbDhnYISXYDTA8eAg5+OQgE4KKz5QhD+PHIQeagASRt4hLW9iLBFfFy
ATT9O/WSqSfMNYmJdXOUgqZ8uNHgKPKXoeEbuVmjr1ftlr+E0rqC46r1czAyY6maGaV7FyRhUFKu
qZVOMoa8nElpdDWtPdgbcvT6uwS+7cmgpHjxgzetXPx1XKJgVs8akEfNPPSHglARWehsqOHZwndR
CrGD3DfRX7pngaD5AGR7TTEx7a3M6p+V66TOrJjrs3KDunBy1doThQ4IzPUoBLXZ2hNDQQNiBfkC
hucNaHt0MOpfwy3R2iZgfKNlYhl9Tvx0HK991o9LWBrsp++KXeMwC1gF3V2O7bDOb1/xCwhhyOec
oprgs9OUhvDBazAG8GuifJtDx//MfTb/ruYk27PUGKYqXekDMlfFsQdc35ZBHIAtLyhp/JTPhVGN
LmlIianudhNf+cln2g+g/MzYa0RhHNW7R2cHW4gDJl63JS3bzUFZ8ppjegt3/Ubu18f2kde8DpTN
z827FmUbiwad/Ch0fcbcGbaeMNgpjNh6KqsZzfKcHKq9HPqzf8EMtiMtCZ+A9ZGDgYpDCtgxahNJ
6fEEScu6ff0hSKMu2HUhHCT/UEKUcjZueZtIoh1ao1l4GEglY1NUsPLa3yTHzBP4rCpmg2q/vEHK
yHOb1H2kmchYsYPJNNmhupQ3jklAwwXEljMD9/gGF1XjLzUyGhZ+gFTUsRoZh2lVvrMANOxL3KC9
RDTcuspABRMR4nx6NrdFSwIpd7eZBj5bVspcIsMbKK9lNgm44qBoQ3tSMPcG6TY4X3nThbnAoM4z
1z8/+d6JZAYGcH4ILWrldvFEV5ImVxgZJEzk/VcYJwDEZAINIAJU6ynH1BG5hXlCMt2otM1WAdZY
O3NA+YUYNzsRIfk0rZXUimfhuid3+b24ePfAJk6P5kDfI/GoNeQffOWxj4D7vM/i7loqSELxlxb6
giMZ0MwA0+P8CFrxzv5t0eCqciBt1copntdGheNcrlh0mVM3NwH/M8qXtA3t18nAX1XhyGjq+iBw
uql83/kIq8k83ShfQLGEYpxprUX/gWhPmMcn6PixNPioi2fGF1jxsAU20iCMLUvEKyxJWNYhsGF5
dqumz9G1ZavrcTZfcJOwMZsKi8p6WnEdLl1EbTbUIqtwrEaBy7FyMxOAcGDN4qSx9ikLGqg1/OyK
OiDFlrgRT2uSVwVSi0XngD52bhkx9lw917UhjBlzTAzxNcFh5wX3lkP5xaVBJ0icX+u7p9kaqaPt
Y3sg9cAml/ZxgxEmj8oLhobYWYWhm8kunb3XN/Q5sT36f1MUl+7UEKX1qDb2ASdqoiWR6PyqSnRp
2RSRrIzXwrtcZOA5Hk6xgfyg4pdywXg0X2XlAiT5jJCeOJMTduRnNGalD2jkcySDIIgStlzZ7XiP
abqCsk85u50Ube3g/BiH+qOxJurSFAph72s3YIbCupGPcASd1k6w7G5z1HXw7oCPRPfTxSOnT4Wd
GGbKhkUgdXUKWIWVB6kc973ek3NRL6X37I/83GHTgsEbXLS6Jg0+uOfqB7jBbKK2i/wfIZoHWWyQ
HHhH3Cr2hVYjuQgrjR6BdPCcU9oloLT6BCrIodn5IuThO5tatctLirjhAgHZ+KLwIsKwYrxZdmo0
d8TgfN+dFgJyBi/6yxiP4Hvkk89qWzCvkHsxXMPJGxp8geQbt1eqJiioIYsyH/1E6Ob/8kjshY21
Rc2B7O2Ccsyr24NA8jSvfqPMW7ckriy/pJn9gc8jWJngQX/mdSto7L3WLxNnaEkkwpPw5J9qhmQY
cauDL/QEujTWktl13XpRdEXMRijoty+gNHRXyizTTsV+sRPgLSKxf5C2xZRF1SWZxtQxSpKEBcf1
Ts/LK4uhnkYbWdnOkCgpd5yPQbqy9pDjIGxbsEMZzV3QDeLe1Dz4cf3rD7tqU7n87ja2emoNY5rg
2GVX8tQ+qx+8FAOOZzYu0j8/ELwDdAYo7a9Z2hKjJBg5XkW3xGSGP8xYjfOUiXw4/K7dsmR8De5N
6JuYXnYh+fbU3tES2Ulhp3z36jvA0D6l+vmoevyl+7Yzqkq3PJNkrbd1jPVdC3lE5Xm3nxJnFIvQ
Ryanqsn/vmISqx/NVzU5jgazBK6TmiTg/LeUDn/0+5Hc875C0Sn82Jqq3xubXmX27NobiZV2j6sO
Xl1GrChnR1FtadgrC/STO+PXKyb3m2h1niPJPUQBFlUVJpP995Ia711Zq5VsRdj9+GZBaQMwrEXQ
9hkw0ggz8BJQjKGfH9gjoyujnQAI3X50AmfQakgtGX1Tj2M1fhvZPmgtbUDDZmyld8lLt5kZvAtS
o59SaRuV08Psis5CZnu5CXdqHvyy9yMtLyauBqOEAPxeu35RQz62FJupFL8kAPeE6moVHg6FgiPS
YG7CcZoCoF/rmUXpksMnxk+CcEZTv7CftX0wzZDvyu3BdBKCW2yhcLp/fIFQKNqirpH7kHuK11GJ
TKtareueTV5MVZxZk6KlFmndzKHZ86fWFAwubHz8eXNYhSKOgpYVzoUPmDDtSKIS+0xcJd0bwrTP
+8wGHHK+MGnzqdhyE5lEbIDg8OXy1d05uoQjkU2EeKJ77d2K5EblTKHXy3f3pJpqFZ/7B3zEM8b0
sU0zrK1TvSnpm7r8Yw4TzqdEA0nbsWSYAMnoOvmAYDULZLO7Z38eGIx9wxjiO63GzB2046EwfnT2
SDr4LZe6Dp90HKSatGFEgNaKe7BAsbLqz5cGCTp/WCFKiffeN/kNhB5ButcmZcWBdwfLcF6vMMUm
85xPaP7LFRAmzU0nrFP0nQrhP1u0kQlK99eQc/vlNDHBV/MLhin+0AxKC9sNma5exIG5JVGyT8wE
qOjsdSfVLT/9Gjv55KKfm42XZ0iH7TF6YpuWVfgLXyKj1Uh9s0g8epztKF245VV8WtifGTnoSI+M
RwjCX3gPWv0SvEufOsVKUqV+wG8aKX8fE3AUV9Oz2GAnWegvedND86wMMLJzjPQuc9DuDmvTLz/Y
O4o7u/bof5IgGc6cnNQ3yXzr+aj/T1+vYoM6YcoTJbYk5ECyZ3gZpHptUgz4HHR/z6QR4hYKQSVq
QXgsfpzgx1qG7VgbG5HgJ5Y/OVYMBQ76BHZIQ37LhYJEWaoBNBxbMKrPKoWHYe5VokOstpgx7kXL
3y0GcCNgpL9beCrbtcTglehb1dRFc8zqpdFIGl0Q6+Ea78X9bKTdlz8BXmLFFcYmS5QajuU3xouk
q2mVWExiOnnlsOPWZVnam6kx2CWy5rF4h894xZtP+Nz1W5TpcBp/TTCzoF2RqlujzKk8VMivj3Yg
f23pUrbfAJp4kK5nQrbxmBSlWER1dN8hANg4pHn25WJ57Z+vn+xZxOhl8chqa0xpNCEX165zPuCj
QuHRGPT/A5qdWafyHJOjKJiV1HZ+WN1tOT7OONmgOITwLOyL2M9D3hUCIx2WM70hHeF39u4KWNY+
+4D3MMKZtCvQV0DPPKNWXrt9DETE7MV5sf8o5aeaP6IpipI9pFTtV6y+AdfahW117SFsVEOGgtGa
ZsStD7Ib5N0Rs34ZznsgbjsOyPBbMfzKWYXheyT8LdBnQ+Z+p666jrZPsIWuxklirYWEr0owTF8h
P2B0FYNEV1HXNgWvyxnXKwIAytse1U8aBhYHhnN9zPlZ+sourrm0vIaRbDSUv+SI2ldk+SlPzlJ0
fvxqY0vg/C+1yeaYWP5PA0I3hRHu6w9KC2eAynLCpFrovWXQzREWQDBiiXWbZC8vUqK8xDPzh8iC
SFLoNLgh0f/uDwgNB4c8EODXsOKwgjL2tt+kWGOdo8K2XLvqSDELsa1hDNxsRBiQ/t2MfCCqwmPG
oARy5++5/GbRGsUpIMxBkqdFLRgPiH2wn35pZiw2BKNBrpiqZ/wuSppwIQIJT2PQHnZOTy3I3tbY
hSc9bTzd3FA=
`pragma protect end_protected
