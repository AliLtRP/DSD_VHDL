// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:28 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
LyeR9sfSSvywo30bzwQGUGFChYTUg5Qk9XU0UoNsg83m7WsaA8yiWmQdnEgiPlFu
ZCecmS3cdJ8bBA6QTV+rLv7/zMxh8kymMIEoT6b/qSrTxz3WQbZRu9ugLUriSque
cr2Kgx8+TCfdyEtfOfRiQjFxY9CsqftNT2hXHM+LxOk=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5696)
QSW49xFOKHc5AORpVa9R8UaSNLu/NHjLYHa/Pv8GoNbG7Jelg6eHvxquPHkRKFLg
pZpm1uWVuo7SfvUuuTKUSKSgFWYKne9m9ZRiC0DA3Bb5S5c7GLWAxNZZxp7wM57W
uMxc3y2TKllMhDCtzgdaWO0gsD621Oyyl8L70coKszFT7bS1DL36zXYpczbtu5rx
t2Is1z+TmX42U72EdDvlETdd87tgSqw/dFcowXCXuQ+RWtfMVF/3tZ8maXHdrVmz
SHfraZCDBEQ7jF6ibaB3l92KKhKpDxBOoSwkCX38jSLmR4/8ZRpmRPRrbaWlCCgh
9VremKuEpAlZftyiWPtQoUoIlrr36iHZB/f/ge66QIpEZgZ6jk7zWYJ533TG9UpX
J411yv2Z2RUsenqCodvttO7w5FZwZffwAeusW/Ibq9HESzl9RfgxLSNAITH780X5
n13u/RIYjw+rTxtPunh3NI8pDg6V1mrhV3ajKXiY/UHmt7ulhYcHFMehw69OHOc9
G9+mTpjJzMspFxveTkQjw/zpUclMTEOUg9E8jDa1vNeDy9HJ0enDeY9KYiFxz8MR
fReV7n+Ozknpiyej3c07BM8Fg4WgVZDK+lJu5uZiTQcwNM2vU7BtxaAnJKxme/gM
uGcaMG71Ycdr4z9sp/cQO1V95lStGRNooJvOQXltAcPTkCjc+kqVQhLRpNV/m7mp
lIWiwZFLh0A7+68jLxejt20+sDqakzmXyD4zDrWZB0ag8wfEKoRWNmc/UyLulBrK
3tTAja9/UQ/sT2QG+hQBNgbj8uOdASvKAeQy31HH4m9PolNF9lo5PcYgAvNNaWaJ
lod7DUnd0HisMgKDfzAZPZaNSrttRLiM15aQo4tydk0KMW7hwZVc4dqL2p+PMsRo
zt6x9yC2fZfiSnlwwHdoeUz6bQf5JqYXN0rWRcHqfs+30YXUGA+O5YGnyk9uNC15
jyrj07sTC2xnqZuI2rnaDDwBVSyoYYrZ6k3LBrdaBk+0g6Y4iLR1CACNy4g8gnS7
/Uo3CEIgejq5/79cg/ua3a/yyeDLym97jtPZPoo+Bl0Id+eQqYYecoupBjiWPam6
LcPLQunKcZ7ctwWsLMkl32l+sM2Nlh6OLuxKTXvcmWCG/IISiP9fb8mCQdUGiI3W
hdCHcxzEbVTkXkaMmzCvZw5nqk/VnxosEn1ulO91TMopfZ4Hr6dWg2jDfCxdqODB
Imj2DWd+Ifl97XKYUpglA9nUa6ZEECixyoHMWYkvsGSwQV76RMDbDM7bbFR7H/UT
pGYNBLCJDxR3AuizYbI/SzHeSwjyffo7xCcprFtKAqCBsQg3ve7bGZTGKgzFcfvm
JRBrYspASpmN9UV8fXOtJc84KOYfWPy9BZ0I9Y2aSuBU2Y8RNRoJF+wC5k4JtCpT
ESogRJGZtgCOXiL2d7oT4UueeTjvyBKEqaPvAG1vmIyIuUWxkwv+JLUzUiWCTswQ
NSq3LEHlRlZIep9HR5wSkRBeyCkZk/O/kB0E0QxobSz7eVxnsV0FJvl1Qix+/riE
Sl0qO8cSzynBgqT02h0rOjYn9StYydoqEK5XWnNtaPB+wFilS3FVyGFBDiJwA2c0
fgZ55ElvvMLWefOF3ksQb13xIjzmtfQ6dmda7TEjCzEsmPGlU1rooNtNVpZyCmDB
EFWDhjJ0H8Dg0Um/l2U5SAffh50ljqlDV1pmdoKPCdZbB+Q2FQXveHE8ptzKRCrE
ueq/WtMdRNpRJyYfA6s5lCUXuFWOvvjk87EPAtfUD+IH1qku6lSrLPIc81fKEjeg
A8CGBf9IFAIfdq2Dgw7xMGoAaUi4A/Stxr1T+qu/G5EjdlG/mWyoFA1r+z8Fi251
FxXx87/9h5egxKL8649GOT8V1vCPDhWVDCQDS27ndXgjuV6ZPb2z2YptP9/zFgXA
7GqD/2PgEJ2f8Ia5gf+5jSnhtXLLptZSOmWAfZvKiJieXsOJ0n6FLB2KnR/xWCrv
3OrpnUaTcUN6iZEuGpF9rNsWRr7OcqzNIbr5jXcSmDysk3MvwiMqAZIENiGbHYiy
n41aiPvRcWfpjZzRRcZQaguWKQXQPSTUB0R+Orenc3CI/mJgiLnrCDVmqRtaY1fU
e4IJlm4bb1WwuGZXo/3szgMQno02OF1OhSOnFadS6vApEVZqz/aIT5aVb0vYf2/p
ZQpZ6ADV0Rmoh5s8uTnqLZlysA17cnr5Lm8B95L1mcRVydAMtBwButJpS6Q3l0lc
sda2NUTydWBDEoA6UZ7P5EadMyPg6RzmTTxzW5gLQSeoXx2EfosMVdY8bQCA6xN0
Ni20nsuf+yI62HUewoBhWZ6BsHttos3tjt5LI0z6LLWDmtEyGazkX/Uc7sQdWd4Q
GiIiFuYVs+Qtn03RiBTA4rf72i4oIlk2obqWOqYcMMTpcUCelP4zXLepQ0h/RVIo
XpDiTd95HPvsnboysLKkiABk2JbI45i14DBB4CdiRWAAi3ZRFAruJWnhFjoDrGAz
6t1at9yJ2+g8ehoOFWZjiJoPZDW1BZTT766y46mxSYcNgnDWBknBWY9Dj5deXqJE
jUGkCH1qMCeiJkjX2uS6ysFIhZV0JOdYR7ivc7Y9cZdaWxEoR6mv3A4k4o1WG2HT
FwEYSiztItXDGSvEIwPaGa2sYqDBjOsbsyxYam8U4m8QXuWkKUDKRMkNTbx8P2jp
bLXAtiuHUzW7Qr1TVOlTeNtcu1cizygaeqXLwuFZw5g1mgVXi6mSK0+51BDr+DFO
KlmS2syeY9+GTI/WJK4NUnOKjYldI8wgB8jSdFgkV36jig0LK5Ivg46M6z6Mv+7a
I0X3WPDW7TSdRLWTsqfVnIOnWN12Ud3yW3d6fw1KgHtEIgRRQg5DE1Tcsc+iZBzw
7KeOwHBr/cwI/iKCd80Z+LUf5V+1AGL17DqKhay2AiwGgcgHMWFsyJsy+KcgGSvp
LnRhuz5wYIHMqv+fte0drRU0OzouTh3WPqUQbkhWypIyc2GRZYgtJMJ3tblE4Bm0
NSEJevfNkcF0vmswwmqAnngJzN+ABtCZYuYFdYT6VJMJubrObVn4HFDGL/L2Zjj1
D/4AXSHq41mwGbFg+DT6ciA/zpF7BGo5LNYbj6x8LsSMuzkoAhqL4O0pwhiU+5SM
W9hopBvd1MTkTqhSyRdt00MYNh1wPyOi7sc1N6k4SWmnLKDFfeZgTA4DQ7S4UtMm
G00TfDlaPCFxStBNFi/gAUWId+p2EYt7BJ0hrQvvaYmU5COth+RSrKp0t8OL8PvK
L0ns1a6R1VOv9hkQenIuzPi68Wjsc9DQqGUzB6Sti8kWTclcVwNoUvjtyGqI5LTc
FPbzTrZ911WzQH163SD0O5jju4WcOmQNfCPIBigOG9PEh08llWUUJmTE3ILK0Q2f
HJFt6JCPsw1oIJaya7monpCFu8S762Y2v8YvEVToASlcfUOt1hSgnudFl56BdN7c
KKeyMUdD+vkq1DjneGI2HaQUblonTFo+3OZULt7MDPhxPLIUS5EsbfK80jhV6VGG
V+on/T+Xj+lQDOYMj65d++rHdoAUGCy+fQ0tCK4dIiSIaJNkpNlAJRTHnf5QR1R6
Ou71QRcdqc9GJVGgh0e2VHQpqOaC4f7pjpRzQJy6zDqUdhTeVYJpcfH8ctO69Egm
PnwNInmgat+QQzxamiZWmrEvmvqRa18CEG66Qztpg5OB/geS47nI6ljHUYCjy65N
4ZTr4hWLo38cjIJArI0IL8pL326adb8kfC05DTL8Ez0NBdBlFbRYJR+uUnc5EcpG
L+lrEaDg8SVFx0mCgdTOmBH/BYgU6oOtSi8UQeJxNgAjLqTV6Aw7nhwoW0iorlSy
yhxqBLARcw9rZSlAEx7odKis+Wksv6vC693hAKq/R9WKxC5BUynDeCbgVt4UjyYo
3+NLJ9OWYvlcZNaLBf0FAjWJ8HDkAdFprfcT7njXbO8RJNV4HMhgvS613yFJG71t
949i63HDyHfDWbF859BU1mfY6ewddxn7QgKqfUPd/NgL3eFjyzXwDrGXxR2TsqYt
aaG4jtDTnbeI1KTTH6nZHT48kkCjQyhZ5s3BpZ0ZIlUWwr3mf/OO1ToB3wSzPZ6v
6kSMpngBwOS/Ttm+Yb1mmGtxw9E5SSuiR9RlVsUR7caHzGRCFGuX0yG6bs+vpLLO
e3Vr01XC51MmmyNZUztowMoVVSDoRF8+wjQ1FyBDh7ZG/k0JmND6jzImKsiae9Of
Nj7Ph3ezpItoPpnaDhRCVy8FKQw0rB65Kj8lfFR/aTVTmL5fHFMFnx7+yDKIg2sQ
HNQlRpUxtArTagdkUVyxxa4pdQ6r52IhA09aEIeO5WE9eBVju40kOGSIP9M7R8V+
pplxoOhaypEyfm5WXjpmHWOCp1OtkYn69h/9J8j2gzRvso2Z7BslD3KLettkbiFZ
I6fYqQKGKMY9T9c0u+NYOHSUgq/0zyaP9m/ehIAtP3gWYrimCkmKiEuFWDwewHku
v+iGZzbHqjxXzjfIDtHHXbkCFaagCh065SoEOdNLaKuKoUqI5iUsZiqClunC96oF
/xhB8jmoiGgK6LcJ+KbibNCbO+IP8kFCi4QxfQ5FtyYUCm9b/Ryqs/lX2dL++xG6
bCypk+sw+NFlGHZA9dFsSp1mm9HWx/1G8IQgMZRGnJYSW5V8WTziRsBJ5cA216N8
cBzg6+Sd/NXzdDZ7n0Klx5L3e3mmdAlr1vFOPMTrUI3ralodm8RspiGjeMUwhTzt
72QkHmmqjDedxJYksOCKvTOM2dA75i5XyDTUb0NGG4vcCNbkpz6qymRFdJXTfM+x
QzhYFVBMkXaTtVmIY/u20FCt01GvYJA94ntTUf+VnmYR7Zvghephw51Q5bOKukh3
ukSthoK8TY4Ar5AnV+oZjkLv0eMh0XaaqkTNAY5SnZSCKuMOp1lcdcFRRV7knd5O
qSuE+hkRhtssUSykg6Hia7WDj/DpAyrhbANTKEnHiBtxRSYcn289CunXJkFUQUeN
CpQMgab2KUPy2HiDcqOr/LDgq4sO/+LFiBHEmFeGK66OkDkiaWRt2pjYBRY9/LDh
NiPTvOZN4n3fpKOYlvS6frb00EoMugWChHJEgrejdWP3PcuA1xO17CHq+NzTaAoe
Zb2BPz2SWLD1o6Y5xZ0j4j8c02vUn7hho8/P5IjtNMgszy99UwZJmk3oDPdSQrwf
TpWqMmhFut0C4jx3HNKFvgt4UuS8yuFh047Syj4chzLNIGhI9nEc/oLkOKZkqsQ0
qT72wWVIbC23rxjQIeHNRl1XBxVOxNdLg57tU6TlwEyfhbU5mp39wFAzJJBhprek
l96JZS7DGdjNClXbpkr/rZjZPWI4wsF9hhVSVO2JLC6BoHGYcvxw4z9X8/Bunqit
QLDBXHTi7onoLvK4bHOA9NVbRZVm0QE1FsYi6Bxw8UCpITee1OEnC0K3x5gs978o
0h2U3YdTnFP9s1ztoJ3DEqpaJrFQbgpC6a+wRfJpwCT/QTSryAVnCq6YFxwi2aGg
n5JuQ5a6Ui/ZLvAClWnfnpLPtJqtBUIXy12XYiOS5l+qBW4iwNSSivGtxzE9ESnK
S0Ynz80kK+3O9mssnR8eqIk32yNcvkQfm4XnjctoEad51g1zHsA8UbuLNbWMcS5b
SiVaBwP3rX7ucqohcvVWNXFTmwiYCOQAFxRyzJmj9ulSMkbnsLoUVy/6oKI2HhEF
UHaqFwouRzoz3wjDRy5fjTHdOuw1K3Yz5fXLKgXF+Z7wl0Hk0gGQVLGkS6jpX6VC
nW6wS5hSgm4nOJ+DDKz7tmOuT+cpMJdTef4FYBz2MPffxEWV5KceXkAnaTKo9EIZ
3moHo9Wgd0AycMGr6u02j/f24fnQTTCsiyEtfmA73YzQbEvQcUPFJ+fUxa3kELXH
DI0rvKoqUOytPPl0PumiT7aDvSBEdMrseP9tLw/dGkB6jcorxGKChkmbzZ0se0mN
qhjNaFIP70m5Td/bfeginO5W0WmeqcdC2A/jKxzTo8StBHhOquK9t3T/mTFR8sac
BHcoHC2nUxab+D6uAXnydOrNFDo06rQJRVkHIAFU5nkgYFIxz4tJKEjiPLIMhMY3
O5KzJovWaHS8aQDm2vja8+3OI68Uh4YvtBNXwM32/Ek3zUB/9ueP67p4nJ7mKsf9
ch0hPavILF+FHYh30+pkeCNzX9IHdd83DKVFhmZQnlLPNdONS1eghvklvySnNUE4
f+sY802ej41lSCQwf4OsA3Ir/cspvcl7Itf9uNxXyxFYBV/S/2En5kK1Q4clHfIX
NqcdkoUXmakOdT+OcaM7s42ExWEpUPPFVbKqiBDGkxuEFlTdAdm8aNaN7KPaIimJ
9D8Lt/LJRanZ8stohQK0wwS6UfqP9HfRbzQu0XMSGSmBjwg19RBGPwvQ0sSbRods
myr7EAcdTT/9bJPcHX80FIs95JgarsEzwkYNtRiC435Ct6PFqtjxFxMDeQB7rMS8
gBQ/rs90KaTzCIO7iUZbaiRwOw+Jan5HsdegwTZLTJz7MovfPM7LQU9DyIyvqk+I
oz6cFdqoNA4JmFvYdp4ti/0099tZQv+NObH8EJR0uehDAHS20+N/YoKjamKKXAeA
q6MGGfVbK2LuWPsRRI4/RwVVD0eFkiFVTpSUfdBOMXvFL9i0qc28CtRYOnrsiw2j
mGc581IJTAN7w7kyJy6nS5CHkRCeT9cNj8da1pmzlOo5sB07Umcob2VylzD8c2E1
v2xW26P2lBiAKlD65VbgXYmmcw3fdE7mdGs9R9IfGCde5oMDeEFI/X+CNjV3RBvZ
9oOv5qaZl4Z5hUG4RzgQI08bheNhefHR4OkNaGLZrAig2bNldrHemhlrLzy/7/0S
DhNgt3qNARUO34FbmKVvl2rUZHYu1YP42AAuKX8ettRvlo/twOq0mGMUlxaZYfZZ
i03G19L7PCSwha6/nkUd7jfxxXoA1/HS+/bd2Mp+qnN+pXz94PmpGwQmMMe0Cz1h
xEGGizMrKPAznGnnHCNYSbAFBrRBwyPi9TvxjiTXgrDZd9/379V4MNGPqyaavdXc
WQcXdr/ciGB8x1g/RKMZ8bnT/oFzehPT2nm/NtY92I/8XfrIobfIvwapM/GIEz0x
ainnGO5iX4icgo++iUb6DmBrWvt/H1/P1aZ3LmtkzpGdcbKvHIzqyz+boI5n1oUf
OcG9bNTCmuhvi+tvAIHdLbmD9KMNItcyKFSc1zOewNKb3MLfR5FMPu8hkuJsGI8X
iFGNiJHpPjdjlOvhd+1diWR9p+hbRTPIjMJOgIaUErw7ooallhPly+WG18EcOt8w
jekhUw4R5xWqR0CzrAoQZJc7QK3nih+wHHza3X1EekWXCtV+ICN27peHhCn7osZr
BpWqZT84+HUyAfvgM2ZYcSisC0AmyxDwIGTzyLGI3gpOIDqcVVmBZrAHlOYToR67
CrBv/EWiHrQ4bAfZ069QWwOBVV9NwIqCGPG+1W1PL5B7+Eq76VgcCxfmtiUecbKl
WmNqcpsV+iTyRzXW22F0F7Y0MlMOMA516R0GQcGjKc4Shn6ySFIv1iixm0/jDOen
SSrm8WHuMSG/GkNnbTNc5q2JWlq00rSIHfCp/a54JJA=
`pragma protect end_protected
