// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:52 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
VKdqk8ROmjmmu/Yzz6tZkxiRQGmpNuuWdbtHEy6pNhGin1AQUZnyNLzvUiuVs331
JUWsGwB5yoZXAlmXVTBmi9eXWuYkTdX/8oBe4qlwcCuMM42p0Y3FYXrFb9hMgKIb
WWTWSHYu7/gcLbYd1CusPZkPgIVQ5L7OB0bORX9zs3U=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 29024)
Va8Fy32YeVmnoo0T0FVfV40nmxNkjSRj7ij1yFRqioW/grWBSev3+2E1z6E1PLgp
w4gf7CLu0V1327Yr7Ez4kNYgmyNMqL6Kw1SEKxyh+0c452VzM3PaQLWhBsW0+e4D
6by65c9Q3FA316g5PJtwXIpC4l+sWEst44L+8P6vaiP82UZSNkE3pPOJwr0w4Wv9
P9fmMrkVpa+hutJyjATfE7fxUTTCnTKbLldaQFin42R3mRXnxXV1z0Qc6c4EAyPJ
kQqhUlye16hFuXREvdec25MrZAiwXWtARHWai4yo7ARhaCT7QEDqug40g5SDeZlk
SYnQAdIcJiC31qsRzZd1xk0iIG4WLjXNGkMaTInjmgWBJbgzyZFYImKAR51B540I
YjNO1iivCqLgCs2u0gXAKbaiat1lHAw9ti1f/3SId1zUF6t/Op6G1p3Z5xGlKQHx
E59s0sWjtUzg9mXxPN89i48/JMEosQ+t6BFdW0mxx9afoST2uIxHoPrBwkceN5yw
MteQEjYYjcFwbljWkBkJdx9CbnYon6rsNlKio/HWja5QDqLVc+6cOKt4rBiDSM9m
p8KwW/B0S+i19ExKVicmatPz10mNdycTVufNzR8JLBaDmdArZKHDi1IB+GiVg0bL
zgSy9dc/W9RSAm1I+CXNzFZGmNBLnzdrXtz8vXH67whSmZjNs0x2uaGilOmij4xv
hST2VcGgAfln0Dl3oMeO4KrzE7ZvA09Ws6so8H3YkZPeIIth+Z4rJyD0Ysaz8IMA
CxqaDI8SdxcTmPDeLqt7F4avlU4fT7ZAT2S5bn54HIC5J62PPLbFT2Z7u9AScYAf
NmVAzNsNHwiNupq3uTIIinnQS7tp6RvkqJ6+sw66V/6Y2060mwH9jOxXfP03VCgB
A9dZxHvGvDRu3JQEAD9w9smb2IXwAaFJ0byw3UJ1HcYyLseLNXLlFxkCYsNiH1ZB
ZBUkvoUt1IdoLuH23xRcie9pC2bxenKbpGNioBXwWEJ08MDrJuJsoHiVgPv5MRjF
rtu+BSBNgF3Ly2stlSGyGuFR1IRIsGz2N3lpssEGNBnxH02yHRDr8GfJlc5rQ23G
HJLmfNLJKAKdcAKzpJNCU7XwV/6LOiqvUw/VrJh0zs6GjDz7w8ixISIZqjyrt2Rp
2QsgJ6NN6F2YP/S5Rm//gOiNQ5xxWn8wpmTZY2shJgErOnnP5WutgX5Y8AFCA92w
8o/kP3JnbMZnQIrhIQN3sM8ZqDOCV/qDYNARUcunTHbYACG2sGAA9e8U0xi/0PGS
Z8J/XVy1r0y2eUTKldKLD67vBUOc/eIDM1onztsWGuRd8rqecKpYGSY0ZwtmQto8
PDVMGt6MsFRsmsi43weBnRzoYUUoABst9g4BouRgome5HJFNF2gEs6B1Dds+W5Wz
EFfW7htk/PlbUT1upvBNL+GLS6XmOJggT0Uop/urw+DMDR8HEI6Q8kFOHEa6IYS6
DocBO22XgAANNx4HEBIx62cxj4elA1ajMXR0WAQRpId9RelsD6XGjzBRfFIjQBMl
/I2Wggojil3UoRfiROjz7YZo4RSWoxPQ4CPkjEqjYgrwKW/3qWERc7+mx31VHBAY
r5ZcV2DY+gEMw9w6s6UnsdBzxtbiL8vL3pmxr0Ndg0ujg+MvNULbWEB1CSvhmIfB
IHtzXrZX8r1qjh8X5qPB1lPGDRA7a5pvQp7yTxtmGrqMa/HzRniGQXh3TcDCQGYi
6s7nBzvOqYtoAgDhP4MUJ2Y2jp6j8nTfrpanr0+PHaqpZzPkzaWe3mXMvnsgRCYL
RfFlprBpGi5DUg0EuB1ZcVS0l4LpMaSyzaThEHl7qT8Ld9eTABLHkQqxNTn8bxyJ
hUN7BHyP08AhkExq5zmFSaE4jLqK8zUtqQQ8DLNDoKw3P54e1P65NbqgXb6YMeam
D3Z4PlTQglbvLrFM49Lu3XbzjoXuwTFic0TtLm5bVPBS953bXS7zwIcKkJR1HsOh
IbcFtgwHZsnT9148g2VXLNV3PksH7jzaQXLlLbvxEx16JTi/AXLdjpJD2WsO6prF
QZcv7cPmzXoYcMcjttYVLbrl8umykxY530E04Vw8NpyKadUm141zAb3BdmHunf2u
SFCLSHnHCrm3OvzzRhvJj+IXyDEa4dSdeDbHgGlG2aQBIgjhrN/s7L4fg6B/cXPT
ElR2UIGwiakb7LUdmTNpIwNGvb1VhNpwE40Aok4MiGnAxn8uNKexN0KIFJ4KgrCY
kjimmf+nXHCr5aHJm3d0pgnYwTDOfSL5jjMlJ1csSIi6aNyGAtmBTO6FrURPw8+U
mOfxpfXc2Gr+fBDvX8x5ZDIMa/w4DwmRFFJeAMUyZbDJuRebASBe6XSDZ/a9UyT4
MKwcBhxtU3gHIXJvyVOimKXXxP5Vxg5DTcDpwUCmBP0IOOEDToD9Pp8VcoIyy1O8
DXBsCYxyRxXgOEeyQbf1Jckeh95WvnyjC4yBzhxKjKO9C896UjTrw/nUKwePPAiy
RtJqUXK9Zue9dfHIUa4nOZgvt9phHq48DGXjyiVQRfmpvJ0k4uqFw8N/ewMlVLsp
q5L2O+eL4TVbPqGBTNvo2MlBzLhk6AjQeuuldiYmO6jwD8QcLq9YZjbL2tqcPtgP
L0Pdk0HUKOJUClpsh3j4kqJskM+EADfNFCuXaNZhm+qsajGDMmZTct+2uH0IC9SB
Ut866ZAYqfZT9b6FIT2qy4+2KoySsHBbZk259ixVMgkwU3k9ymaFC9e9nU4lxxxB
lGG0l0cEZr1dHjBxm6KW3hx8+ksEMhIwqrQll4vqxBQB4/PRjaEmDQSokE3Zu7Mk
5gl3Em+QTb2Y043S8iKGK+zaMqVJlhH91JsFOZozCx87Tv58DWw1R0RrybtEyzrF
X70ixjw4XJ4pwOA8mS5uKb69T0Bmhr0XSl7qztMSbSm2eMnf6AiPVdioQ0W0msLx
rDs+gxNGo9VfrSls9oJHxAfM3ieJq67GRWUqur5kplzTzr/iVcIxX6FQwLD3KfJF
+2/EhgDpMttWVz6jds9dCVglLZAN/YpBw4UZ8Wc/7Mhpz9jYPfPpSIXDGDxiTB/3
YrIyWO6dlHMhH32Z6sySCaciW4EQjjD7SmC3m53nfbK+wHPl00l2vG3CkjVLPnv3
nRpW+broaNYu7LoGa8jDnuzhYONdjLjqyls+zjf8jKRijcwARrksuBk0YB1JdWqd
gRoWjQ9TyqQ5p108nJEf3U2tPtoswAH55U+3Z/3z16z9LjmzGsrxrfEJnkHnLSYc
nHPAlArYV+nfWS0g94QFwPMe8pUgzn9hXqwSBzaZlj5nBI4xr9rW9iS37+Cy41wW
LH6K1ermm1NARwjaWgTpWBpGMgnIRODmEsQ6u04LzknOA/gopqC0y1i9li+8g6dT
0cynSAhFoNEnBJ7aoV3R8K6IUw8y2HLYTOgg1r0aUqaiZY8GlX2Nm6cox++lgq7v
LoWnQG+VCi/0+TpYnAMA+Y6oXoMb8coAMm4qt8FsbfUj+MfGf5UhvKBAyvQggirs
kSv0rGb3r3jMGGSn0cBPlM2lGvFm11bre4DirnIvPW/8pgQfeRlScGlSVsMT1uS+
rlMBmCWEvIJgaSsmawdpkn9pxM5GRZgq1twiMINgfSSrkBJebiC96nIc18R68tAd
scD27zYBrlCNenCh9c/GGkvuqnFf2Maqu9KZ7y7yt+61UFa0RU83Rx54e5vyG56f
Tjp7Iu1ctM6PfvCAlfKrFqRHYPRmZxcwUR5Lf2mmHUk/8GIo45vXlyG6tuVX9swj
GISveh9vaJ+4G8GhQLLKI0ULt5v6xgB0JTBOnFByCaohjkqp6xhG4+cNkHCyBkMS
e+eWL29ptHwUCqNgMo0L1c55SZPRlspWr/94USJ2oE7MDKKX9xC5CPL3zJNPVtZI
qyS1KoJAfkLpQcGgSPQVm7CFUdrtrlt35eH8Qm/XmydKvvH8ib6uFW72zDM8tPlP
hfyymZjiyXwNFfhOrkOEjg8810oOTIkbO7AGGL1MW8gqvDfb2Aq47Bn8wwvgFXEt
u7mHcl+AhJszHDrM9VzSJvnPq3JgiTEkUGqovigenbTTSLCGEG9NXZqOYZMlaRrA
EmoP6jkk1m3ElhySnJLiO3lpujgilGi4sEML1QcuUI6AHA9zaZ2NCE6A2NwzI4RV
862rC/c0RMCRJJEe330/4icpXiwkQB/OAKbYg4KKSJGCo9LiNPYEHpMrfwpDgzHn
ObCgzNxn7jKOx90SmHtCyTCnwJ39zHGTaJlM1aME7wLkgdAfgzGLz/U+hxQUEVrc
YAmkXtmfGZ+hzSihrHHJKEDLIHgtzl00k8hsovgQTWvIBOD/2SR33QsdQE7S0Bj3
pEdl3SbeXFeecloeq96NNGp0ro2Kj6LKiIQvaGCd/1Endlw3caYypz/zregfbQ4z
3Y4Dbxvzs8kM9TMu0JAZT61HbclyJct2Cc8dSUVNg7uJH6GMWsZrTtxgjegQ80C/
cXgh5evovUpXUwshpj5pow7yov7ID3ggQZ5uPLstSlSQUgYdrohpm6GNaHIjPGEA
4KqaBibDyVO/nawPSVQzglhH/FHkZ3nTvMoxjp7QkB7fuC0ASewhwdu/RDVRN+pv
5CWxFFMKudKL3NZfjLj2LG2eNNQ5uBBe11MVgXpURKylsFXLQ818t7sj0kRRxYZh
ofW5WtB8U/T9wifr6lUSMIBHD3y+q4NioHkihOrtiAh2TOHzEP59nXJcmTAyV/sr
sWs5seZnwvOPchwLf5KKjQ6BtKnvIjqMU7q/nZ/Ub37+/WW1+P3TLN3u/hjAvyYH
pgCc4xirrWlGrkqGNhfCMQ4sflGkWIJMXdkbkkSjLrEAbkr5s8dH1A3o0cBlWLgx
KKwD0czcqu4zPQe+SZorSeHBagmaXU9WMa1EjQ8TjNwxcjOrcoM5kBctvVspT7WP
HK6yEApMfi+BG+tHBwJ15YvGFtQyFgKLDtc8Ohj5phU0PGxYVFdTzxJnQMVmEc/s
oMARbYGKQVR6PvreGZH7eqoNtsuBzN42ylAMIxmJk/e85FzPNnOV7bKX7VJWj2cQ
qtuucHzmVskHXF1FO46FxWVvq0yboa+7Ny+5UJB+M2m/OMTL30yl7zj18MDicU+O
ddo17yDTmp31EbZ0V2h2fGsSQN+F5Rrr6qlURUGKT4TCdC02ivpZ1fmEWUE0P5ae
0MrICIwefqyDQ1+OD52epjPxpsBqo+wmFm+M7rgOTY0st8OGGhvgnYoG6dHZ8lYH
qX1JDRepPoMtntwu1PuvE4xMUT73Ri0dTxjMVROvHXddb42ysE4aCxoSiGfBrafC
f4GId+tLOKd7BE1cUzhdvJ5HQDCtaArzEfjQis9REBlwywsQ7Gij9vChi4HUXTSs
g5KI5Y0Pl2vanmh6YLWJ7tlgPMYerAC2hS+bBMV3hLQAlOL6BfgyRXcfLhbTSmyV
YFKv9MLKLU4LU9RqCXjm1vOq3MahySiEaxzsI8rhZ+cNfdGAtw2hMzSXA71spu/3
yS4TH21QuBhATuYETAdH2WEg45/EHopThLJ1zylw+30Esbe50XSk/i1Q9HsFhPEI
xejoBoYJzF22wUA1r+1ffh/E7+d2JPwvzZukB6t70F+n2ub5cB/x2WfCKY2smHn2
I9Y0zkI4nud6d0bOoNm18AtJ++dGaqK8mwHmumGD9pv4pZ4+ZQjcDqRsIiPa8yAo
CHcpsgPvykMXH1AI3PtYham0JFocEBPOyAGwJ1Q6wZBkU+NUovieC6OztJim5ss4
Qb74e3T3E0q6SrizmiU7U6zIrn4fb86w4BH1KZ7f3BSGcrxkzPF102h0ylo20KZS
ACaPIHs0ZgDJ34Oxv3q8bracgg+75ARr3+zUBjWaXuB71dU91vS7IEctaWGfUmH0
NlmOLsOTAMwMDUbIK71Gq8wTpkh3LeTJQh8XENQylGCFO8cFXyx0auZ32fpu8CC/
f+7cmZrT7Ew0UKXW4tDAG5pPR9SfeA7y5rfriwltfFRiYCZKN+2tr2SaL7wn3VaB
tjLBjHRNHQiWDvlzjNLq2vv7tEFQWykOfe9fWA2du4NsqrLptmEDDxLrw3dBOZvL
ne7hx9qDlCpC3Q7eOWfJjfiL6Dr8zw7zs++hzcaRP2gnjWIAXV5ZfRdyEQQM2YEn
S9Bd6dVcYcVGXRUj2+b9NylnzwUhP3i1RVpv947Ztd+F/NEEoPGFXRn0AcBwoLHH
KD346nu5cRyAJVsCRPHWM9tX8yjFe/JTObp/Uz9875tUzA+oG/40NvD6guGMaeTs
R6RC7J0THjUiPLpzs5VagDexz2NIj9sfYWPWmU05DCJ0QP30akBoFcv3EYpjRZ5m
OS3IB6uIoT626VK3e8sExptBG54xEtbiXC6/LwzULqRoA3oj2TdlzyKJq23KiMHh
ahojButAIwtd/1lIGw8Mh/ufgt41uB3n7RDudgVWfnbl/T2ysGjulqORBj4JQCEe
FrDfvwQ3nccShyi2oDwiFCwRY7oBGwLC0W8rQYBVD2JABjq17tB/WgUsy+pUUju9
rmTYPbAc0brbSkaQpf3+Ar5ms+9m2/CG2r+ujni4PF0hySChs1IhHp4xc7CXBxmN
GfKfE8KQRz9lP2UY5QKgH/YpOJbABBqOA20qIKhwcnZzoWpf6eRqJeD/GDOtG+55
Pwm8c692a6902OLEYEqSQ8h70t7pt1q5Qbd5cpEaJeAIMtWjTylyeWQgM/k3fK2d
IHeNul5OkWWOTKD/ReQg+yDyY7vWdiiNb0dw+elQnRoW9yHMAVgPOR+iKCvYLugh
ZWR5A3FI/1JuL+j0S/dE4BgULUVAHqdViKgRrgDaH0rjI1GK23e2etkObeGuXQUS
LCjNNPeGwK2rcTZ+p3UP9Du6wPI9NT7MOdo7pfgSjHxgNG/ouYAFLV2LSPqKriF6
ApxT+sU7qJRtOG7KNuAHZmwQY9HyG1MdDDESWghtLEI+4wwKHSXBMKVKfAF8s8kg
TWqbQtl4gRxLtsimklQ3CIcLyrWD/9GqJypEYNH2H+l7vbK+SIZkFMfW3gv+AOzw
7BExF3sTyX7f/2GV45r+KiSSlQSBt87Y8Gw6Xcwlitpdea7uEUPbMK7P2zL2TQIa
8QnRPiHtVGOoNy/xGIR39yfXpHE+oPT9SiWU2C2Jofs/Y3JuDx0v3jbNvDf1v7ip
Sg6Hjesoi9sTa1Qo5R1zuECTLiLPmIsCaQyv2/DKzaKkrMThDMNpUuakEUZcPy6P
3QX/CAbfa8QPC38jS6tfQK7GCR8QU6V8wdb7hKLypjMcC8rLKapmU7juBM4tLIYO
kyFURfES8XcMaJmRCCiqzPjCBkDODVXEbGVGe5YiqUbqvY7DpvnWl1keMHPvmjPx
RDiNxhLza8zEbHbpjNzQUQvWGYOKldRCARHcWst6YSjMt3m8P3oImhwTSLq6P5r3
HvKXRlS5ZM0CLNLuTxti+SKUxf/VlxrDAFU8fo64NTD/ACv2ha/WvIkPsEhq77Bj
UkkbPYKDawChxWUDlliWxfjYH3tO0WUjlZNNEAggAylC+pAQzpnLfdSbP6em2xl8
KHgD4GHbEOxdNTj52a46qXic3HME5tAus4jRNRzO+oX0MSqi3Jp3YdjnrO8zjnox
Y8lXk7jZmT40IIVvrH566D7OVYKODZwWfRee0ik5pvoVE2yxTPlBJDbaQdDSw/WZ
2WMKterz/wj4lOzJLVoUu+tcOtPHQ1UKaKzplEds8gicP1t4QQr7qUj60J94yGz8
TbezIl7Q3njPahVdB4ECz3QXtqu0KA0pHOdQupdvOK0COX4AidcXDLWPPIyBNZkG
A90vKvooyWfoBFANfwkQ8ZldamkeV8kGr2MweKxuRj46dX4s1MWEMbDCCJ1YdXjd
L9qmSOYk4J+shtDk3OGRhs90jVZN4VvtPgTJjKBxf2LKPaXP4vQgKCxsTJUBND7q
fe9ehg8tLNIG7OzAXIUels+zpCd5xg9x7k6cUJZMxLea1PRJUtMfQ6M+LekxPg7Y
L+S/d7Asvn3A23hcuvCrXlyvBbdbd4lxfScd7S37weBI1NK/qy3/EPRtEhnCTAl8
q3/zRd0juUpMRu30S0dPmSDmt6F1sA39nMkQYhoafHL3WJKybFqIsoXsrGbbe76G
43IbQkR3IqaJ5+ihhfppzDR7si/ODcbYzpZNh+elJRzyHwR104FZXO5tVR5CztmA
/+YwzLL4m1OxJqA+0fhXAA9qfUkaMoCkQ/3Flecf5BScpf3Se+0ZknB/DyLgzz2n
iNSe3+0jeuKANDh5CDpiMfew3n9VLJA3PWSSTF8I+tGZA7xMbqQwCM2p7RHHDqBX
FIgV5ex/8Ih5mRLeDfEhhb0aQrVg6etrrid58F4mkMGT6996VhshFmI0NkN8fyxq
NLWiGp1SMKtV23Hx2/ZtX3eDuk1x2FXgA5jczX4MhO+ipPpjMb2CpwZkSnWugjuR
0BOOdem34LMkFW9IhClxPLf5wUKliuIp4xlOTyKEuaIC3piYXrui7D85c6Z2fStU
2Nxch3LvnCkWPoN2jAH4egvmdvnJWKOXSqeUOtN1C8oQyZbj88h2ZxjOQo+9ESqK
unwPSXnbqsuY8LECJ/YU1nr5KX9C82hHby6oCHd4V+Ah9ZJEUoptZm16401I4pko
gUR1TW79zeaTICozcP2S+g5fw4ogdfLmk+eAhxtlEIdv0tRPgAgHxCXGZ0TCUR2b
whTDoSBGbpBV2k/NFVd1OcqrCJdzpHCTpj+JvzpgShaKWxga0HytsdTeALkD6HCw
DM37KZHws6AVtvmKqg3l35BjfybPT365+pwtYvYDT0I6IW6JYdT/cz39jEl+zwXh
HrYKrp1T8aY2LduAiHqPhUfO9sF82ViuDZVNxruoSg6C0Se/f1UJdpi09S+mNjC6
+sgzPXZ7+F+ELcZQHNoVCHXSu77DNbVdIVGqYoWeovKts3aXpZD01TAa120pCAr6
7hpsevXE9l9u2/PkUCxvmaWGeS9oUCjrtUO6Jp8HoIxFMsi2u9TX1gSlib+oYmk9
LVhibZ65pDGjpZoxKCz/HjfsdwbtH+YpI9LH62UKOhvk104jFyaQ/HEY2P/LaNYK
aryWjd5m57dKFHsWtpUdhazUMW9+US60VBPdlDP7Q2wiJmcfLflp9Tz2OMpglipR
oZvySYVI1RbbUEoTF7nBJGsf5tiBkrmaDmPpdq0rOssqrZ1Mztz1LfWeWo2vXdzv
NEwaKucSjpbTD680kwsjAtsFrUOklPQRuNUIDXTakUDxzyL8gQoYVGi2b+ERVE9L
U5bA+NBeB1CugjvhQ4+AVu0uD/rnrz6KeE8x/Av2vMYImCim2CcysD9r9awkVFi4
d55Q/MuFvz1lAgiJ58sVE7ps5hrNthqbsw28gQpxD65hCZqJf8M+3jSYsZ6hX+TH
i18J7qOnQaM6ZMjpJLr8o5xd4eQYG/Z25iF89YnjZDeN+3gLX9c/fpdF8bk4jckM
OIVQBX1P3Hg4TkAkYl9e6Nj5qc3FMavFsORW0vFbLjG3Ciyh872YZHvnuLO7XjW9
3ZK1nFkwdIX6lpiLkrBW+ZG5D9tCNTFuTLtieupD6b5ednvaTmmZocZWOp//rZEW
XSoiH0Hn2iT/A2mIj3xhF82MpkEM6hlna0XeMnPyhgpJkaVv9cPhOQFagxCEBW/S
Xq0OMxU1qsQyOPycDJmyJPCPfpXl+QvhHRlWDIJZzCxkTnfN2iCKxmmnpdjVMmR0
Hj2HRMWq3fTjsPl+50El1a6pOA1eMpmWoIsP1RGoPtCCQ/QcAud8jvILYUI5VF5c
8BrmmfWz7ud8dfXeQadSRXDpzSD34n9TxCi28fdd1mTVlKLcCUgHdtIG1/WovCog
Akxfd//ON6EKVMHh2OVAocahN5UeeHAZ42/TfiBGa0PY0V0AKP6UnYk6aETNkZcZ
XilmxRokNQRHs0CjP5kcwClctk5sG4u8nydppd5RpPa4Fa5qIDvObyRQqWIEgAfX
JCyXybgiBMgaVWg5mBE0hXS4f28FsseEgkocnLXS8+mJnf1klqBSKMkwmdigJlag
k667bU18SIJhnBSoQ/BlKoUz1mDNKq2lftIMeQiglvCkrDEYpa6PcN83quMZmD9x
Bjq88LwpT3sp3QIN8hry+F1sYoGWB3g1wVSdijvc5Xn5eTDY8BjllK7cCHirHb++
td77u65eoj6aYh4j1G6l1Jg2tnVK+CC9hrV9FiFQ8Dj7nCZCgSAB/qX4SOMS2slV
G+Uod0t/sTqc+WIvXFLaxiAe4ZA6yFqrbzjtA5vm+H9K0JYWXKQ/9KaqznazpXss
bfVb1j6v9nkuM125vyoaxkIgPsWncU3LPF3lZx149zIQMQ1WAtJVmQAzrPv2s2jK
GkZvLY6l77+nTEH2uoqLmQW0zDxzRohJiDj8J/O5jue2tykoL2JGEnapmv77Hh2M
oQH0YIf1q/pxaYdlUgf6DEegRS74ELHwviRBYg0vJwQjSk7v/i/g071fGP+TQaT/
nYO3CwxsENyIh3lDpJw29/vX9SN0Hc1IGA0/6pe94nUqUQ8xJmLOwenafSeXwzwR
bJds01mkyqHidz2X0k3AqQLLuGiPsfTT0XMEBG5O4/Hl1nGpcHY/bGK0Qt0VLY2v
pWzsYUPA5ONUvtV/8kEotQDWN6eVdUZvF7yKthsYKXtlDKbhkOrCaWrMRhYWbpui
NyZGCrL8UPKC60DLcI5aK+FMBH+uGSfyPf/Vk9YPAk3YfLJ1FMyN1Fc25TJlHjoH
ZnKFrWvZN8fJpbNehqd9oL6HBgxk9jvgHsMaSZE0r0xQF4SjxNxwytUXRBuE7O3h
vxDlpIgVCThR4lEM0VXK1A9D2aHXuDZeCHxYEKzgdxV3DUWgXfhAPVS78WHloUAJ
0QnwNMyRe8YqzCes2MLLgO1cUkVKSKy3pnOjuIQ3ISJ/VjixZ8AvmaIhZ1rhqj8H
QEf3fBXtfbkWddGepIn4U8FgkYe0/Fshz0o8Rj19N4CfUtWoCUN9oAZxP1mwjI39
8lIhNwIzdkmmWpA6F/orlzH5j8tHYnsiFGaxx1NieZu1Pao/CgL3BST+B4EGrc3d
xvdWVGOVia5kSw7equs7r5I3DsrUiWBTanrk+X9/tC1dmXQN3KlH0OLhlwA11fVb
u+xgRffml/awKg/oyoowf7bjHatfxlAF5grMX3+xj1/vqgreoFvbK2ma/J8/7k/j
8RvPaqxOM7TWSK6tNMUsqHAAH6cCNfXjHGOJV7vT0uUa/uavOQNDvqb6aOi90cUE
ccs/2tw1yz/T1lSj+JZKbp9j4LPbjsiP3Hgj0cgvyJD036mpilxswdB2mDFqmW/p
di7lC1Dapvx73qyrZNEoKrMp9WdoGHP3+JBloj5Wk2iRY0IVVwrIb3n1l/uaVc9H
TeZGITfmYf/lD1WmcM0j8hj9H54rA0e8BIFFfkCAt+BxWzpvNt00KLRJsmIsT8T8
i+MKheoV37rcdCnQnlcIeAARhMNlwoT9yivlraBj6osCfaPDIixK4LMz+OnD31iT
juysKtkaReg/QLg0hVGboQV3d13le8C8kyyi2G00LyRCDoF7K2yUO0WcCvVwAX7T
+eXpZaHa7Y0FgD8/8U8pXT+41OZxqF9oY5Kk6zXPokj8R68PIRqiYQZf20XeuSsV
2e8f0aZ+GlH3X1AWdrCMdRHI0TgVx3H8/CXW3lS/90YIVocidlKei//DrvMeyCO+
7FlnO5H0ArAf2unr/nHkErGksmj/w3jafv9UBfdk961ywXaFgo44F86y7KnIrVJ0
N03EeQVGrQXamUfqt6oGMdLUtvwZx7srcYVd2ciTLsIay95xRwIUHhJTGKSjnkao
g8rVPyqt+IC3Uadw7eJZZTnV4guiZ8X6Us+WE6bWkhOjOnea8d7PO6YN1VwSyH6S
yFt0/IfDTcrmoCgaEbRMO0CQW+a6ElUIZKWjMdF+ibmgkNCzRKFAfl1FHOD9LsaH
QtKMro2WyYDoasgkLOr8/2q62geP4+D7lYZyecXNn0xUVwPVSH9ZfAPKaUUhmy9X
ANt9xxTrir6GSBEG76xI1eUJcUcSHiDf5avUJCjlPkqck97hMXKMHaVmXlV7zyWm
UfFiz4F+dNXDOUhUZhR0re7VD4JBOdQdZops6PZn4VBPx/ikrzhoRzTvITrxiQCD
NqzoeQmKuK0KNJ7x4v624tcCGnRhRzmmDxW/VOu1fJIJur1d3kpbxpeptmkdL470
g5L56b66lvnKxjaChYKQLauiKMVuDvrEOJ6iSYJ+pm4prmbQYI5GZsAKcr2mFqSu
n18lmb69RHanQqlx614QvnC83W0zdChOPNRTgR7EAvFMPNxv9urHZ5Q16DbdHtlA
hl08zKXcNcjf+YwYXXgvOyX8uu2xMiCNU1qg7VKFEW6eHxvh7L72wip7BXx2DmZI
qvidlhrNg3TV5jTjD02HXQb5w+81vxhLQyRDUaVvHDI3rZPT1+cImdhxHOGAwmpC
xqBdQO/fTFya4hVEh+NRYt/mUDpLypUJTHw8be4vg8MHSV2yAV/7jeNZS9Fm9F2+
HPA0yz5yrykvbHTZF5hASkCz5LuDmXFNxpZn+fN6ayN2f1RjTqoiKPeV5mKSeA7Q
r/q8A1JqVdXOko1scAuVKgPynEp5QXOUj4AjRGGQAWBDu3Cv9Yt09sqM4HWDFbLT
0sHWWkxF6z3H7/ToatRqEV7wW1qG8kIujPG8wXU/L585kYdsX+uOOgHP6nqESly1
bmL2LKyVN8HlnBzG94fesW7tcyuwfiYWqQ0312WfT0UYEU7UVfmlW59TjM2vi6N4
TQvgM/sJq/c8HI6X3DvQCDznOHx9s0Sx96nlCJXI7PIuYuQMdz+mTMuONU1J4eP0
1YT1+0QWN/O80QuKihWDTSxj/r+hpfD6nZshMrGkiwExcgYRSyHdZsXxg7mGkTjz
1Ksaw8xOuwoQYfLueqTuy/Iy8i2DeS3ozKU31wk4WJpDeAs7YOZR1OnGQQRNGppo
pWJ1VvSZS8tFlD8Yn1LsfmHeMapOjz3/h078WcTYvraNAM4danXGuezNk9C5O0r3
AvFco6eaL+V9+uGTNLZpShNFzVOA5KBL4aX+E8+J4X3jzaHvysfaUXoMXnCO9n59
UswlRosXwNlm0oLSS0UHXdqBsRQR8T9N4u4Vd2DEEehUTm44PWEcqmyk2Xjyb0km
6o1KmwlTnT+Q2mY/0GwZbO9DhV57XuX0OTKhX8uX6uwwtGoeT8xTOWTTvKX3uEnw
9qqZUYSvyWr0CDTWwYibuybJkRtDDyGLsNJvRga6nh7JMRk1gMuC54kTyeyZGepF
YKJdOt0JvUSVTybcVFwyv7NW0jbpF++f9EN8M/G9lJsb2QdJ1LizqcpzFNOQGo0L
WGHRUsPIChfxs5ob96H344uSL/hNTdpk0x6RMXDNfkwPUJwa0EPWPCxRkrTGCk+c
UZWSb14/mXtxW1STIE6fAU8FC1IhegnTgdbblsvNmSgV7Dqu3Os6WAzqPJ5CUHLW
xdnLoKXWBN8KHsEDrGqXe6zyv6dv0n8D8jsO/B0cg8LGMxm+ITVWdqDUB65F9syt
JTarrm7oa6T3+RZzEJA1Hu+wy4caBcHGXg72N5qHSQCvLv4wssRzc6byUmjPcWox
8/kZ9g7RO5PJ16lcOvJXjQcInLIS+L6OjROdlTAE20Hfdyrv1H5bIsOsonQX4FZZ
O4ot669FngPc5W+2ej/FkP14suldAi9kDHT3npp6/0qWM8afIaHEf78nJaEMYET3
TTNfNkC46jsCSRzlTWR17y88H1k5b/8KqnyWqX7bQ+O6ldJFvLbJ7+PPbLzVjI1a
+agi408EjgfBpxt68PLiSAoKvomqPtXt6AQzMg6N2Q9NBpxLNxhhB8eBkSFTM5jZ
OA7wJkR1g6mBZNmjbULn/NVsg1fHtnbhuFNYeVAlaRWvftVkXuXG2e9XG/SkFQVo
wrMihoLmTrtGTpjkAbcaotpiAJE4ixugUM1L9Oe1zLOdgehCTgAJbZULsFZpyHGT
EJeZwThtfhX3lPU5YN8ecZ3szt77FzjxasF4a6y6d4tooJrfIZtNelpS/q8n5+H+
svXjqEQ40blJDIESEXHJPGhBMv7TUqXr0Rj+SHU2+eVp9QhbWYPY5zYi6qmw5+rr
nVXo9fshbW/U846x+rHBWmQZf6Y3R6EgCmO+pbeQZhlK2+p2CBOe6BDwtP4Ph97H
9xNStbvFP/5YwC/SqNoKnpr8+S0856Wpp8CEoiOnAcoe7VUns85lI+iqnmGWPD+W
YeU/ZQd6PoCEE5+hanY/lqJNQRqAOzt5xCaGHYZEWqS07J/mPjCLJZOwbw5N7i4L
y9qi1zBtFOdeEU+yLQLY2+LTk1xUVg2qj5lM2HLjCHgVT6biQZGbwAyfsjqvqA/V
XCtDPOC9kJo5vCCm3ru0hx3exjgpnB4DEnztvHn5JkW1YnVnfZdFqAPUNnzkyePp
fVgeG74dqm/NqLOi4we/S9pOvjBBuy9riisH0lojYrF1rKGxOn0hJDeUzF+B8J92
E3UnGBe+/0rJr52UTtWLPR2ygm0bMD2lw8QbGmJ5u1M9tn8jw+tVlQZoYzPUXW9h
OpOi1DOQaThr4vPg2fnLLmvrOuKHtEDiQQ3Zx3kyC3T8sxyKcubZ0ou82OFAebjQ
rKsX/ukRiqyeKlFx+5auYmgWb7V1aoyixb/wVtr9p+T7kVEXk2TRHG5yxzfEHwHR
q41DxuN4Oz7VCB110Gt6XVeqzxyKezBqa7PoCR3diavE6GcQjn6mOpY5DNC3TetL
uUKrjKM9ctclX6tyC6PM+Gv3Zw2+ImjGI5zBUqvvOS/4NqDa6u0vZhQMG+nHxAga
JWW3O1QeyGmHScF7tBXgdV4cRZDOHBGOcAPgiKcIalznl5sQSt+DBJX0Q3Aijt60
xP0ZL4yFSlJITH+aR+/TiFlPk/gIIl3lBsK1f/V1C4a7TkoMB6pXeWYx6nS4ZHra
XTAjzwhHz0KXtisoki0M/ghuof66N1JEvCpMiO+zpl1M1mGibHSdRIunh9Hm90Az
srN6qkHbqPss2w5D1F6/Qq7l0bN0lX8F4PMLVpWHwqCu2XK8wh6FCUWCIPejX+w9
3RTon2wCBK6lK/1VnMP0dFEuIpIXIwlfVTUcIEniP7e7B/dlh5bG7sw9iM0Kyo9T
grTefW508g1pghVIOXCERIwpv/ExCmByl0vBH6R3HLKa39ABmDvHMWIeC8RtRHeq
UjBUWdwZaAZxVt2EZ71ipz+DOhuHMgvBiRtUn8igrBGQ2ZLmmB4+KCHQ/ecXrIlR
LhIbV+Y/ToKbpbrGs2HIuon6kr/5Z0OdstXkZsbVDlqHPP2phflYX4QCwQMIvtKI
SUDnPFOyfwQ2U8eHOOqsBk/+7f7dj9pZqmSRB9lie/L74avVYhSD3OtyhHWp/ZCl
iZfSuaCeI+DwFfBrqR/uW25piAEDXAKPll+iB8Puq+znNQKn+wJUW13iG+Ox6prB
q9lC/BhiTCwJT46cnzFH0b+sSD0TKKRitOKudbgxm4InM5qo5b5UOtWHL5sOigAP
l8nDdv8QiGQXn69buspV43RHuli14XWj6/c5JNzIRR0Ucwf4S6Ep9qezTXq1RbxA
mBFuLj6PTMTMHAJI4a0XQgR8FkYvi0aSIlGzgDwERd0FpM1KuoOyGCgFobLtW+cv
OqOe/6wmrpn/GTf1aBjQanbJmlT+JfYdu+vqwyxnTKKg9pDg4bf6mqr4CHHMt850
pSYlvAdP71guv+kEf6liOFeimAHPLKVZ1hYkROKOi9mTD9bo58jDW8Bg6BgKkP4B
0NCaU7cDn+NmWnCA+I3P5lqA0GpSpjfYuxL6RiYv4/SaKdy1Og2+VrSnXvu8I5Kv
F0386v5HfT/hkgl69GiEbx/LeEXUmL1/yXRkWei03xMpSoaGPlFYmoxN/MvlWl8W
4/0tiokVB4+lP0r95j9hz/KPrb9z+YVVHmrG8Fh82/hcK3LMzOAI1Un60hMmnQxZ
IzHaQri5Ak4gCzG7XCeuygxZtwmgJ+5oH/wB/Bv8td6gspxT0i87hak1XMsFYZHf
JIdFHG+imqYmOv0rmWhE7fbI+9YGKvh0p0r1GTNjXXsK7LezEugleX/QswKozrrQ
R4/+Nc+jo+9u0+rXADruee/MBKHuzIMQ6xxWKV0vMMEtR4BfJDBYkdMQjnBYvXPr
kf7iTlpon4oXWMWm16SZjQGZAdB4MK+82CVxajmXVvOK2oqg1xufDsHcbKaTrDc4
cxUx2N6TMqlfws6IbsZ0y9rTIXi3qBffO16BEbZ0VZ992CFVRfu9mtQTnx+o5itj
M3diWdEEqMJLYJzoRpvUalHDaiUXtQtkhWtn+dFPlO3LTjs55xmToSajJM6My2Ot
1h/jELRwhV94dPSAEpzD4Zh0/TCHfJ0NStRVhKxocsl4xzsvt2UT8+o4nJ/AKYTJ
rVkZqVXBoAX1Mkf9qR/uLEEE+5cWNMA1EvZ2jmQVvrDfzXWCjl+ZonQ58GxzEkkl
hOSsGmEhSi7PcTpG54QOJCb77Ug24MztUycaclnLMbVHVALYb0IixZ5Gidq3QpC6
7vxUeSgWfGEyxt7ypR8oept71muwatpdJHj0ovMAh+iN+0lL4jL130MXsHhNfMsH
a+6Zgy4F9WuYVc3bN4XYP62qIW2YerA1XeV1907r9qU7r4jdqLpmcMm0DDjVrsJq
2CU6dg70Bs2dmlIPqvyF+RmuPUnOztNhcZZKuuTixxgLzKyVq7fpNaZnt2PqU1mL
CzagKr2Jdy0lQBQ7IbWWBr8sU7OkPqPDC+ZF7LthiBsJfyg94dhl4WBGBE58tDtI
H7HgGy3dM8uEVRDit2XtbPechWhByo22QQtVhL7Udy4NmuwqEV4/IoGpMoBfdtME
flmGS2cOZxa3iri3icy1o8SWvoP9F+syhs//M6ZfI2GTskUsEhUZGAXGnGZV1B2A
teliUTsGh9kjY+qMEZbE6IYtsXU0WIg2DABH7kH1WfgGKESEXyTLKcFnhlSBLfgI
l5gFjkyoPgJ86tOOsdXNI9lP7tBdjctGaqD8OirKxeya+1eq8zAC41M1b6egXavd
5dRrakrIdq8CYClxpp2pSNeeDHHURODbicfKgFVJtKvkVQbnRFUNqj3XAYQVFMuS
ctGeWKRggc0RIq1T8bqBlN/pOSLHCpCAV+kI5//rRXIsS93scO4qEB4+gWAhPUKm
Nsffy0SWQ3Z7T5+iO9yftBB4FRCtvTOSEDYlPRn5beKXGtz5R/1kIT/gjpNTQ3wx
9eM6GxAyZgEdbPzho7FkNYEntvetjS6RX6qt+vWWDX+hZcAmsz9mwzCOAh15C903
Xf4FN8+cHCnhlUymPyDF6JP0Z7tgMJFiXfZAlDRXlqMM1QNFdRB26ULWF4svnT02
bvE5G7wq/MTwqIuFi/TQ84OotlaAIk2mn815hGBADaWpxNNvCwfKWf4M1tvegAlm
aXOA6DE+zCcBWVqoyshhNI1UL3yYDU5N+djtlUjbe9zHNof5l8PloFGZe2lndM/K
IAv8s0JL2JjeB1X5X3aB5lr3pAFFs/fu+XjgHOcLIRcIdVGXTXqSUh9/x/D02rvc
IxwKuRJ0Z60urq1tIL9XOI+3QNQzKzqQbdOWf4uwwFn0elrxDpUkXdltyuIm721V
exEG/T4nC4terdLCm2ny+Al1MjAekGps0VZj/QywYlPidkeL7hZ2iEWPsplus5ET
T1LyYxAGi4GdQn9U6hxwNsOQACXEvvVrbwGHGi6/8c7leAdexR6s2sHotGXPPZRH
HefsuUwjdtizI2HRXJdp4CiqK13Kl1GWrGBzMHEO3UCb/dCSpBKMw7WQrJ73KfVh
vfPCN3HXzlX2xb0vnr6h98zzVyJ+dGn20/kO0zEmYHO5BkY/zMs8UKvKc35aTGwB
xUsHFH8ArJSZD5FEVU3UnMgHCXshKW9Rr8pOS5q4ktoA9k3/HLpA73VqIQU2+Zj4
DM5EjdY0HoMgXn9jMLX7Mq1zoXqd9PFKpeDMwG25rC05LteJ5gPDmD6lcEuU1Ccq
G6npMf6NDty1uJov6fHxohXn5OkTR9OGdbfSaghhaLr+nZpl5ucnG2gTGhMFUXEY
aJVExojh6pWgGKIlD8sxjHPJ/Z3fsPxLOElgHqt2YSBchxK54zQopVfEZUU/52S3
iFrSH7Xo8bX8858ZmB9O+E+WaGbKaw2qAyQ1nZvpXvx5CcxqUCBk8ABQG/y+b2uw
prCJEwF/Y7f+v1kqGAQGkefPiKd5NCo0OHFx19mirNxNi6DJnjVWrSpG19SniBk8
bRVviIc5GKDlZ0uE9Xq/DUE1EjXHZxYKK3s+9CctV8cm0l7B9UnPACxsjykhaoOJ
5N4visz7k5kYiZzJdRGwMoL85HNOctM47OG46Qgm7YukyAuvF2zywXC6uvRP8/Ik
Z5XNeV6W2HDoOBG0dJv33IUJGllmlS9lhjdckzl2yCpdcEtop8/hHRWzYSxMbaGi
DgrpxWzbNHzviclQqWRj0zBEDQtocURVDuE6vhEH9YixEPXB05mmgqhW+OZs/nmw
0DRKPhY3++m+y3Ymb7I68UIvoOvyFwq+fOM5prRLRedQBuTOa/IPOvYdqHo3Ypc7
xylzC1CLIBXmhlIHoe21y4Tm6NfhVLYm8g4k1hV3DEL0AhH6xPDknX4ykzn2SnK/
vowoYJudG2/xZoeN/CWvmx+hc0llX9wBy9Z49shIkTuRDKn/k+odbrmC+46B/L5J
8bh4vUrgz/F5ANQzLeKadpC9q0inpBGfmTz1aosxxHs0xzQcm/aPs/YWIpjgXvqH
60eKQGMv3xcerXZPbZnnVAn0tJh9+3ZCplLg0aMbVLNVOzWYntQ2s5TH5Z07bb92
5CpTMBlzNckKdvF/RCLXJMqrfrdMTJRR3wyG52y4NYguQXOKoSw3xFQoC8QbQyJJ
HUzwh0IhMDzGE/Jn2i8uqyjQ9wrTfbj2PR2jJlLVqfi0sZgzjKVG4twKLC5vCam9
UP+5sEgRiMS6/gVb1E6fZxqiq28MOpgG/tq6DxLkwzeGgP4QLSpNaW9RVlvJ2H2x
dutNDxakFpnzqxGLH8oakQ8oVpe8juPu+SZU0PiZ9ju5nchLVRB+cDDwBlDXqKDr
vV/3nhrMYXhwZWTH3nLf597Pg+5CVPum+CjrTQWeyFrZPIVHjviBGAAVpgQcNPMA
QDRal7H/cF/r5zoukRG4dk2q23qRYHDud0UL40seCUcqqm3k5QFPAPs0+SRlpUVm
PTP1Nq8D/kYiYy45y4Bxyxh2DRLUQn0+xdMFRqrkrkcvk0121EkrPhDg4iOlGkXM
wvdAeOeRKEaiDz05DwOCUc1IzTWOOJtbqd77M3Flip1/brZoA8PwFmOjhHAOky1N
PdHQp+B8JWZvbvJZ9TD6EY7EXuU3X/1i4TASONC92tedae+cAPovXXJ2NFFLBTiK
SJgCkYcz/13mdXr/SbgD/1nq77QpfjZCGmh8je/+L7OqDaVZWieC42FcWrH0I9G2
9dDZJzI6N00/6BDfky+HlqaNJTiFpzAhYNNWw9VEg1g8G1zY3tzRR47AXHag6/cg
zEEMhK1RJyh+5ZvNBXs4ZUjPfpaF+zgpvW8Gad9in3yNvcxOyMYGHNuNiMBa4h9h
/YLnnrtZ6UNmpAvR7/v5ZDmp2l7EhsRCXCCcdl3AAHOErqWg8+hfL8NsyAkc8BMJ
uppWmmKFaHKxFxW2wF0HZzyLXWQnlfZqaO1wVb3xbRG5obgyITR0VR3xGP8ZAfzO
baLcj7NnCoPwAJ+SR6e/AEeSIw6hJT6wVCs66AxH2X1SqZwDap+XSljsw9igXf5n
dziRqyEzIuc5Bf4mMI10DGv9KTxSTBsV0235p4QfkyrI4giBQeJsrVpfI31FIxuU
1g0t492EAKZeJDYdzVQ9auIl88Pmdv0MmBblCyDAtzyjNV7YrRnfqRvYDVa3oTea
VAw3QiI9V2bCslV6+Xh6/ZP2YITL+8Lx1IGyqrKIlp3Dgw8AmevG3S7iBO/No2yQ
c/FAneHAYXF4QXttKkIuX0y3g9dmGCTCoDE0i45n5f4jGelJ0+3C+E3FDHCkkCHk
JmmLLma3msxqsMuYKt+80VqI5E89Rp7fEjMP/EMY0iFKqH269xsv2SDb2tyGVZJE
oti5BrxK6NjS/TXGv9vaDxcwpw5m5+GKLmcuKX1Tlu9mSt3QXaejjCiI5YY8gVzJ
iSqR/eIAsilWhqJe870gEW4LIdHFNug1XmKbguYVyzowiX2+HL5TSn1Bp3+3Nss6
OZplbBci62SBtviZniMzkXJY4iCxRzZJ3jkq5Ji5caryRSF4nPXG+uFwk9j8Iare
PwZs0G0I8sXr0kqPdZSwcNK1Y5QFGR900V94wq91meK4DInyZdadvsVP8tAEN1yw
XgoNBL5ra5E9LVWhct7GqLG3WHOW1+rBaPwcRnNHQ40+6d9mF/cWjCb03psSBPOW
d5UxpJ6Scre/wFwxsTt/uPckS30nSPltPltiMjoTfKUXdNhin6xPhPqFzNgbvRet
6XeAqq8epG16OhaX2veQZv3xReVj1ef6W8jPvi1hnth+yf5+Ae2cZ5rtXc8OzqL7
5ENOnGTXWPkiJiOR0HFEYeJDcUU8ot+A/+4tfMyEDFO0LoopfglXirrtcckDZsvw
X1RUdEpmk2mHawzckaG3iRodOa7jo6tywHYBD5CBCWQSOLlSLWvkVYWAhVRqyvyy
kubOJk0XS3maWvE6qIfMPjazjQLi0RWd9NSEgEJk1xlgZxzoR2tXTKNbgG1Q4hp+
a3fqN4+i02BXMeDENBSa4/qN1HihqDbs7UlP4Rarp78GPFLSJ+DIXESlANHuJuQO
e82pDxPKDny9xzCX9G83eF+47em+TeYPYUVNuKjgyrnRhB+ELr6oyf5uPgWklWNx
oQPwwgrTag+glB7c0/7aC02T4LeJkIaRDdv6YlsSVvCOakpAG6U1WLxTf0pLHSqc
5GozrSdGqNAXcT8lMXd/NNgMQ8x9sjx3FwCgmx7P74HkYh7jOKGututuT69OeJ/W
9SoV/9QOF0Wc+/0tQmIT+OQRyiUg1UdbvWlnT/LUPNzPqtlnT4s2vXi5usi8RCaw
CH7gnJVO8ZmfPLgvuDA0Yxr+dDAyQI6eyamULkinXtKKa8yIoDD1Xl/tTwdyu+QJ
51G85/Cj0aMSlzHoCqbNeRC3c4KFH4hYOtWUUzxbXJkXbxKOUbnJgf139Vlv9n9V
zIFZqU6Cv+WonmhDTYKomcpzV3Ett81inX3peEVLSUa177WBio07qItzbwwQYQP0
Am5jteGx2UAcmo5st2qYNfaEoRTRrl8bMF2GKuDW8krbdpX1/XR1TeJmSYhd8nka
fpBSZJcVMm3qnLWrDfnwZat4qwW0ZqNBrSgneX2J8Rrnyamp6R3eZlO6aKNulD6h
umqwaPEn5XnlLZqBhlBtTTA1d7t3NWLUlSgL09OxHvUYL4Elit5fs9p9psx98zLS
w00M8MruOaFr9IEB6k6X5WfTgtDCHZMIfipUEt4w8bSPqc01/dyk5e/m4pEdp/6N
3akjC7VOsGbBRa6qSHOfnubsInqUKfZOwnZQkXq90dKYmYOTmPOMLVD6bUlsEnME
8cHCxmMV5nn+e4c62aoDsxCLI9VBzlYmJ6JQqZErC8jkE/FKC/LJdNohzWrunW0y
Aa67uuabyvsDytQQLgUP2+T/Cv+JmVdV9vo5zU8rZPfgGqJGfdwZ/IsSjFAaEie2
lId5DaSnYbKmIO8143TKQArTJbbjpPRNPphEL5Jv5BYzfjUrLDiNr3/aifn3lcI3
TG7y4xCCGd4xJsiuLKAFjLPboGRxnopMNzAPZYU5FDKhKkBsbr/q1t0jxI+Zs2U/
axfh5nt9Fkj+SJhUNOqWOTSskw69MHfS3Ki2NZfFB4AzJeeLzYptMvQxTSXKIY18
5SaTtptz9U3ebHP+0FS7uW86VOZf+BVIj8H5y0FBorRkqpmQHLZuRvUFtEXntMWf
Ij4UpPhm8Y0FIgeZqGOLn1sUqddAa+iQ5JXG7K5skMIlkQ7NqFM4C3tgi4euk8IL
mMKMV96e7rw84xkvdLJflWu6GtctxRvg6xWN2L4FAdtViuko8Gu7oyDQyUXoudCE
M4vUiv2NQIn2ivxMOzgFsot0ioWDSLnvWPtHky4H5pVb7Cm7VAE0L/bBxBhCaUH6
oaNcqigsD+h4L7ZaRu8NOL072h262j5OKBB28eqZfDBwm8QgjPBXT7K8QY40Wms8
CPRPPius0bM24Vb/fM4LxfrOxR5YKHheVlBpNrHl2XUcNGVSeTS/5rgmrBPNTCMO
5h1DzAT3oCY5Z7vm7Z71o7Ed0DEe49fAY11R4RkpLYyB0oz8HuIdGgUCjmo8nNHb
WViwXv+/OuX/xlKLMZiaIeVKvygw9MfPiVYSr3yYYsTQucylgpf76haNdYI8t1v7
TunRRba6Ng7PB8qdLKFUPGRrpYYJQuNJsk/raI0DgFtUceIH1HCdBI25dE35ou+0
wbN9I8Lrmku4VQ8l3ngxu/cwA1D6dFDb370GVeZxsGizQUL3OMtMJMzZJDm28aQi
4ZxxUFz925EoZv8wlDQWtRjgKN5i6ytayFGg+2zZp4/PGE/RxgZI/g70YZzOFwhn
CJfbo4/JKet990iUUuKeh5iqlxLct6lBUy+qhfcvJur3OAEIOef2Ht4XoNE28lhh
VMukbt1wo17ivFt+Gek8JbxzG2ux3GKBAYp20fPMOl36q5nJMphEqSVG6AWODcWZ
LhmnFY4Ak0TlI1ywyx8J7WIzxSb6BvkM8j0VrOqni3C6Np9ya4Ht39FYo69FNtDp
uugcrP4sKlPqoqEX17h3tM4s+s0+VBeiS0W2LAbAqCZzl5rKx5bUWP/y5Os8uQs0
f9PY4uzeYYIODmqoLje/C9/+4Hz8lOfXI5wNMTI4AsgJDbeXCz96zziZRhrNbv4w
9hpL4MSZEfo/70RUjQ6W5/5yHoXxwOiVKt6DVUo2WP8HQvESClH78O23A0nxIlgo
97PrxSUbvmbRw7AeO9k1yG1Ydp8GtD4oy6bnUghElwtqwhe/7N7ITgl09U97cTp6
qFdauXeIQeyGgwS9KhIIvSnNwHfWApdAIm8DutTDccOV5VhSFYXgipyGmXmmSg5Q
cvVfDuf3w1I4lBqyl36fV+RQg+yMmrIoNz/2YQyizpFfgYg9G1LNl845S++UUIS7
aVvUnFKOZ7Nur0BMjLY/RjxY3mex65ax5nd0tsKSeWCdbovii8p6kYmiwcFr44PC
De+bsYpFTouQ/JcgOCRd8xtkC1E4Fb2WGddRj8AGKWjQNk84NyOJDZ8k8Do6TqG/
ItO0es9D+S5qv5vte5YDkFWJTWzhOWFyvJNFkX4Q1LAoshvCDSNTbuGVc8iyR6zY
LKtVIZ0QNg0aiUSd2DfTGSRcpzM2L/QOpQQ2aALR8ZWlb80cV2vOg14ncS6R1PEM
z4kpxenbUMBF19AIGo9uJ7rmSgcsSjRPX+KU+SSPR904Rk40UEw3eHPjZoTCoHlm
pJb8pfAfBY5HvH4M08cTc00KMlmHDPAPzorwwlso8gNbeOsw5d8K5JJ6Nke7Ex7V
DL038HPHYAYlnX5+R/WPzdPCEgKFzJyFL0QKdhnnqe4jGVOd53zll55mduuM9k0f
QZxBJqe27eFhnVmyQ8SY8UOH36/eJkVsFUz9Lh5eb0J5QYER+2ZZujac11XWcdrt
zLC+Nn8Yw/zbl4LDZ98+OxgZ6O4xMmlikygjFl5bislvsDEKX9CVVd1GGGmWPAjw
Vm+25DnXR4m5AL00/48bwAGjYbjZsMXGFYz5g9BZZ12aHJmS0SmClgVFjvn2snuk
1BxIYYmo+4xlyGlpIUo7KInIAZs0e8iIqhYEkyngHimxJkMm+XhxbbdiR+auiQTY
ShaX+kxQO2jscAMuJMnS916YG5/DcadNLPfglXIh+Oi/dzJ3DTqYVUohjWmrW2u8
5MKqnMdBLMPvpRPtasjAU10p0CeOXAp+PawX4iCHElUJ/h6ivLE/dWo/LX7BLxNl
UXGUTkstpt1iZlTAFGKZiWdtjOiLeqy/gU70/rClk2SNWEiS3pq41QK7W4z4CUy6
bd3djV3Ioff6lI+vGD1l6HbSll6KStW6lABCpeky51aL3V1hM1fR+VwtVDtFqeff
mmBklQkxF9QU3xdDw1WGQ6Jl6zEP8bHRRF4A03FFn48l+nrZdIl61paLYvMS1TLM
LMHDvGUyFXDCmTYDU2O/1+rYLYgQlMJZYP0CVt9w56v+0W7xMbpCIM8b+Dnp2dts
3RaQCehcfgB01B4gHzRUtKF8URJLVgfm4GS8CONtDFCI+E+uAWANzxcpGchtX+Um
c6ORThSNetEAJvVPd1JC15kRoM/hXldjSFkOJ03AGptmOT3pgpPZ7Fk3hcL5Y7BS
VUnf1PrIrhZxz8WvHaiXlSopC9f85sH+m3fb1GMKxdKhJY+rfcIfWZvLcbSS2a4m
DnZY1pf2z/UZIvI1V79nfySApBvKlhxKdKr9aok+VLj2qJ4CEGX1ooueY6bNj2pi
1L630mZHYjc4wm2h+ukVH1+hIkDvO+g+NLWHI7QU3G6gXdLT3MHNEwXbDgfP1zWm
voVA54bssVBKHpbOuM1GdW0Q6R9lPw1/wyU/uHkwOwOdl6L/oIs+RHYk6oAL75/8
rSrycPEy+FpKiaPXPu25aeEtnlkSFap3uxKPALmJPRjL5FPpv7/nj+cBj55Ty9NK
XVjOYmqVqduB5jOvqLPsIGLOLsTJC8xb0IjE/HD+Tg6x+hGqhM63vry/P3qAy0/F
5P5oy4p/cm+niV1VsLbetNeiDenwwctTQQbAL5K6UBFRx61i3r2TRCL9F5A3PrLm
NnxtSrjh+Zmd8U0q5G1FZSQtw3OR4j6u39kjO7Y9y18uYPJI0euHZI3PizYm1lyl
RCQO+M5iymLqYGX3SpTvkMetl26WjZ/oGYpD7Ot9o+uPnI73mTHzCnN7bM1zLngs
5T8Z+UDSKp3FBSCrfZJ+u5n14UjLPLyKV54So3vS9tzXrYoILHxY46K6KkONzLCI
hjTvDyW4xEwGNczUni2HhDH9yfulUaow4bf2aUOBw6tlh3lycMl7942IrTb+HiRj
lVDApHk/+NtM/1UIv8vGXzD1Bk6Ksk+zYgE0rD+4fZ9EHxIuKfUzNP1DdBRXdNdi
Vux+8vroxMzTK7xqAIMr98qSRrZURF7vKBj9NzpiVdZ2HLLV5lLZxHQWp2DnXj8+
hr4eRClqDoXBT3pAXuhLK/68UulaeykuhFX6MNRVfbPSt7BFJPte9W90wMQY/j/W
hA2ZI4RVNwZ7fgm4nLuKGPZDpIL3WapBWg05EzwqoWg8acwD7cutY22g2u30RWIz
DorMMCUD/ZisDN3U7NDOHemsMrwy4kEInafTBUtHKjlKgHd5KTXkJg3ECbG4ku/J
NKkNpjvlr8TOVzt8ANNLVpXgIMLlvEWAjfDAX/6PPqogo7rdglK3EMs1Io4JmfYn
jJqYHhebLJX5zKRwgAJX1VwreiPvePr5fUpaF8jPHNAL40uVN9bVyHo1lcp6ZnCU
mP44XXN3llsJxEMsc7QQgFr0HtoT4JIYBoOz1pu/hxKBeQvPNQ83XaBfW7dFxDBF
ojhXKF9skpBxa11juHuZh7ePDDD/TTwI+uQ1H7jDvNc+x3tCJwQywCtUGXfQdi1I
hJejnQCFLPzQrZw+QFAEgtl048XV7p0X9+itC0DNLjGN+NaMIu6Uq1ESiF1pYn32
Ul60ShAgiWeMjmfA5FjRCrmxgJVfXRVEfpQerNojkuuc8/tg37gO8GwXU2+GgX8O
j+QwmOpexIl7o+Bp4hkGOeI2Ir4r765NhSbOtv0Ec1c300Rqdj2fX0cXLxj7GUAS
UVWt5+PTS+68cqZwqciBWdjUNAPIJE4vvNW16LrhbhRXOfuLlyx0VFc9Bn48/1In
D87iRLIVUYGQiH2cT0er/v65/vVAwn0FGVvVVYPj+j0k3Tvho8MYwQmAOFWa8yhg
k4ZjTjfJnTG+J/DZ5bkB1oYsWtSGjQa76d2knFnfX5dMjRuQL6tNOrDD2yovpswq
yxEtvlWbRfq7NyOBAGYCRNF9w4Zt23yeTnTKN/3kxv8pxlCLDMLxZRkSkiSQ0pRQ
03i/w7L4X8/wAxPb3NJy6/tTqYaLXkDfYikRCgCk1Ayz8guZGNOb+e/PdgZ5iatt
ihIJ6Igo2kvG1pSt1f10u/mkDPTpCMfGkm1pSHDnlwPUKylfQ25XS4ZL5w0EIhMG
aVDAeLQ4hs9oe0CsDRevfn4L4mb/GVHIIcmDA3zjMppGx94p4nuab+MZGmNVpd5N
p853dbwV5lgpfd9kB/7oSXum/114W9akYRzgj+EFAVB49Vnze6/D0BwhQ8oFv5Im
/luM8SKTwT1vCxrNylEo5E4dqZgCRTA7cNCQ3ScfGG3cffHHtagVLS6iDHyv4erg
nP2RTZr3Dp22N+SINktg1DfB/4JinZLs/hCRtdr6rcqzsEV5AmSueMwAjNzeoPsc
lblKL9gJhVO0WUN70C/7icyLoWdYC5EaftO/HHPLZ3XQ5izXRwBc2/o74A/CZMCd
X6KYojl3mR7lEzmgpx5QNaySuzDKdZK52dIopO8q3UTKeeI+vpBrC4TD9AFatT0V
U59w0IgveVmeQ46dJ/0/rbSS4Sb3szGeb42mTvPS2jChvnrextQ9CX33TE1FX9yE
TKUPsMu+LO2ObymO5UTFQoSa+mWNwUsnz4dzWwZzuBvjtdLY7gcNEHL86KFlAUc5
5Umbx0UzhbhlvEYpzYBo2A8NXPZYWveCRC9yHKTHkh939hP4ZM67neyEQW5jh9Zr
yLsmOWcHK83Vc4FbMeC14EQnKDU2GXfbq53bvc5LzUte4SiuLOlJfdZHvnH2HzuD
/3AAzt+im1dcpkkx/tfznFChmjd0fDy6MuWuqiS3ooleRmsgOTkI5rOYsd3khp+A
VgWMb903dJCoL0i/QjQJiS3DgFEadQ2+mAfNb5oJpA9ja9Z1MGd4FQVwi07JdFqN
bJqo0shqOKjymKuucj1m/0ZouGGcEqXgnxQavejZcGOevZ8BHDtzPcQ19E0kvhEJ
ofyTANJNp957CUmKdAaX9MPKe3P4rBebazPcj1N6WO2ISYRu0dCqALlwWPSXavzX
CPuqeQake2FWxOzQ0EaU/HNZ0PuFyZwCP6FJNnrA5bZPrENfA7eURpMKx3Xai9nc
S83Pg9n3nh0TMFTHT0KdMhCW7RWFFHZlyb48q6u+uuiCrFE9m8nQfM8xCQP5ikRS
5mZsVH0CfConqKhRPUQUQlbQKkBDAqW9K/HWVsrwTMW6BqQtsBk8Hh56vKnQSYBg
07jwW4Zba15ltoL8jvq81OVkuPag+oxLHhGWZALK4/UeiaK4rz8wVlfFBOvtljXy
z2u5VYMvxxF6cDhcIr1KcNRB0Coh4Up0lYRn1j8jdAAD1pUyF7ya2QqPv+IwDxfQ
PzBVMQoaYEHnAgp/3UDf156YJonBaT13schE0+OO7IMxdtpUOIwHQkHPcwfZQg17
syfybRvInNWHS9BQSnT3VahBSd2rftmdcKN4wBn9Vl3nKDPPA9sVMk+ZdT38p0kG
DN924pg4yb4fjZDYurT6AKhf8l3lHpdvi5+UjzWabysniKLrQNCUWP9q9P4wuCN0
Of5XSmZzuus6sVnUZ1+y4TpczMjklVk/I2dCVvZi7LbSjPBL1vR/vPkMP1rXcB4X
JVH92CHsgA8mBVxyTqX+GQBqQTVu9pvP2EmjVteYqXwExsqYQ//XoDjbk3S1/czv
5zGO3lBhV/jowM+qPMe7jJOO4Q/mmmTF6xM4nfhzqou+XSr7hJBgwdS2wEAS73Yr
KRGcw63nVfxqAaOLGYZoW9MSiGs1/hV4QrjB33J7/oMc17s8G8DTOicM30XGTN5t
Q2LX6PiiYu/UOm6iHN7FerS4V4ewWicMznKor6EFDPLgFVexljUTWsA+I/h84NT/
ku2vtQwIjEhkSixHWMav8tvzMIEktzSbAvMXcnAYMXk7V2+F5UZ908fykkPXnrr4
E8Ajfqi0vfYMtFaUsZePCAIoqGpm3WqeigsIbBaxQeSH1SVwaWM1xq4WqqgxQ4yS
fVoBNl3braSgDqjMnXEKxPGL5S2/Pd354c4MmIz0Ct99ugwnGmM3AqaW4CP4zHVd
8LRRTzZIUu5bEWqNOCkWOysThnMv0aysTyoWX9iO6ZAE85PPAV3381oMnAxLm78b
oKzK8im0+d4zo+SW0UxnSrNOUq6UpOF5kWRQS5gJipPfBl6iNPeYDiMptmGU82yN
EYOVNL/IXGv+1ClfNSi/yYR953av2Lo9u3LXh0e+MgiK7j+q9p1xFb3ocevDA3Qf
heFXD10QuTAeudApp16Md+dsjVYLTt0kAsqkwVc5aLurIVOxpVL4hAArcEzmBowE
gjQsgYL/baWHo8UKg+GKjKo9DPCkFgEMHVEM45tyB7vtY1OkGvJXLRNAUB0faaF5
yslzcU5dknAhdfplXHI09zSKY3LCGkADPASmnIr5URQzIPZy7Z9zKCut1RV8b0pq
kKf6fVgXyKYDRJ1xRulTrWGWKOuLEzQbaotO/9zbiyjvyH9B72b/ISAQ9bZvidey
kt0gjwej2sYaPfOf1BpZdwUQ9Q9R7JuoXcnuAAnWgTO52m+qmUyLnhDrM+zFRUPl
DjdZEa9XBT13/9AGA5TZjtSERiQ0p0QQJO7CVel4EFTObHNdRhc/r8FagwZ8WPBA
XeOAOULTDHUmTrXXW0CzpL9gIF2/bPbeDPIipTmTSyzJkIiZNgG3+YkJHWxgFTiK
WHgwY3s9uaFN94Mwj8v/fJuCS4mWD0eE0twa12bqjxeKio/Uc2tQ+SM6fNigBCPh
eqDT1Vjo2Ff9bWBg0xtuXg9JMo8dTmgu4MfJePtW2k/Z3Py7u0lp+Qn4DdkwSMz5
afMePqBkHzls4nt7pStmxRd5hZ7AV/Xx7XlsTTRiZzIRDZzlKRVqg+YkQ0ZyxvAP
f0QjKy9Z4KF8k/SmZA+7gvsUbERRZcuygg7/gJWV0hmg86JGHI2+scIX5v3z7+Yj
7OyC23yLvOAGFMlvRZJyQKJ/an7VcyBQ87zyPLbMxBWYcolYLqH72KPHsr3PK5qJ
+O5B6SzqaMW/Ol3p+XZGLxYAiKfJkXg+u2iZoVdgLFEPoXGcNW+TB77a3yDgOln9
wfPMIEc85MLNWjPS/gX/2MtBmku53ec3hsHwNEVa/QWVwB0bS/CEO7LFZHBVsWDB
7KnWkrz0eRd4PNUjAxtW0xA/8TAaw5lhRIlTC2J/4GUG78jZLx+KBqZvRMTFsUn0
COTwOBigEDXp+jI0poi8dNiCafsmdWNo0LoOdK8IpKk8oe4g13efM5e1NCa2lOZ1
MhRmhq08uaDI6a2EwpEFq3qiEcaTJ4b8tyChT+QrHyMl84w056hT8uIGPOsLCA7l
y6Bke54yfLjErZv2AOOeTCU0kYVNvf3ZqI3rxGIaN4VHh8wAu84bzeL/5MRz8aD+
QAKiiIGFxfboSXJicOJlHFAc8pOisFG/azAlBxBSQHjMzs3vjgAsEfogc1dXE5F3
weeosrytKZsP9yoXjk+8FI2APoPsSm2wsjimUhAdPUimWWvvB+LNN2jPMXCh8crz
baZtl9I+71JfMRUsWMXfd7GsSc4a0KEDx4BOrqZxAQR8T06Jfzuys7t2h+Tqujf8
H/cPYc2cgUZWrQtIClgYrxPgfw9MTJ7nEj4HO7UsXbAPxtsJ7rA0WNBjlsX83FC/
IaoaBZ/LAm8GxCua3Y1cBZz2lggULkOdoNgJQ4GiYleOhxU5BQ3Je52NrJbaEPpH
DBNlMj0M98UXc69/TXqFkLLKfahFn4Zpz4SQQ2lQCFYEenGh1M6bH0DbEaDzDw51
DomF/V1NltklHGKEO69rfltuHyHfuqj3pXH/LgfqfZ+qYgEV2ONdy8iB0Dj8rDuF
upraW2ja8EZj/P2VxqNRpq77doxxg2WIsDH5CQhCdJXF/2GfG/aBplIeIFVZojBj
oHR+eGZ3HwE/jc1d9JqPwNiwMqVAVsFXaCYScLCjDiqmTuGD+4hd6ElpeBXULrFt
jQfLFxMuek/qVYSO+rm0JsW9/iotsR5vA1DqYsLF0Qu5Tct9eQv2vJDRlNfY1mUH
049wdKnws3thoBMzbVUnSQNnr/LPugdKyFv6lYdnmhU0BKcZZbwWNfE3qjwof9fz
HOn63JVf3ex6MyoXlUyw/WDaFT0EgmYJAPgkLQWBHERLFx0URS1SyZK+jYSeR5no
1cX2zQJocptOWaV9xO7f0+y8kGEQ+44azj2U9YsH9MwmqbdjC1BK25WAUs23ax5C
BmTkfBjXrQ/iWGHTYvmzflEIdlLNDPN099cP3gOPCM/CEMs0g/94q8FBqOJdwSob
u3kfArd8Sk6kodcZkhtwsFmU9u998YkEp71zaPBo3suOefGeeqgeuuNTRR4cJdUA
+Fg+i5Fiv11WprHy9WvBZfkcEMwjInpaLYjjo5Smg1dGXYShxg+37vryqXNcAOLJ
gmOHH+448c8ewPJceAvIY3Nfrzx+6JajOuPGx1QOOo0l1ramY/7u5l2L3pCmGuLi
pp671+OnpLYeV/yZ7aJQvNEdbR7aF5udGkab7FxaVNrWwHW7EOWVQJpfWCt+4AVl
QTus9Rw6t4xe+EhKyR1+lWXg0wOvFGGJIrHwPiud8vtqwdr1lMkatSCmy/fbPb0c
zU4VrxazrXfFhppH+JnLN+VR32I0zOkK49kWAI6Uk0fwmVhLi4amtxgSc13mv6r0
eOoTF7rxI+b/gOwBfFVL5Py6m5pOYfK4nsV0gfvXD0C/MC59LcegaAJIJ4xQ2uBm
XtQLBrvQ1zhmbo2+crdULJUS6M4U9FGrPoU59ds82cS3ZkWFTZTGrLeXuOFbwVVW
Dr0zxAARgXfHhg+FhhHrQe6+4rIqdSz5tplp3gPbHLyHx1KWHD94zrntWAv3T2FX
vJwM9bHBaAqefwKy4f1IcCaQh8gtCKe1XDrggBa7LcXtrgufIzxdt37ylbFGJ04U
4M0HoXHkf+IDdoI5LbRAYURFI4PZiJpkL0NT8zZeFqsvZqZKrJB1Ff7G0UH77nmx
KfmHj48//W+HGTf7YAFtrS9zoxXW9R0IpfjvHZjnNZ9YMue9DLe+CY4GI1woU7bo
JAWRNE5T0mdrk9YkyvaBz/+uK04ARfel4Rz6KgVwKyPmwHQT1YdRuGX6YgR5m78M
+TZsH5MtJ5ke66zqcIAevLGkMTPQ81zhUwwmujBOdNEB7uDhMnWoeU1YnJGtKBLE
kmmlPR+0yMvQbqI1WrBCTH3c2wsRdWngxyxQaJ64douKGQOSonS776krYsfn1t6s
FYPcgpL/HERpJiyt1pm+XruAJEqN4oj1efJKzyQhGJb/oMy8fZv/hT2Kzg0fUzV9
lbNZVSGAY84uUGhrBT4RVParEI2U0VyACQXguTt6L2S+PyV0JQr3//qP4WLhpZqd
UhzsWBEGKsLwbJwiSrrPCjntdHfscube1PVZQdAhehYuVAnbh7nNcLy2xRMSDhSv
1YcNdeEIPp/rW+3xOsFNvP18fL/IrpPPwkSoykcryFLLQnMW7mz7Gur6h784h9R7
jNeftQ2ltUydFCcWVzewTh+lKpjUl8dRlgNLEFAzQ8D3/zIaqO94Q5bnSlTfcVVG
06qCb/2mRPQFUeLP4wQHs+B7iGwXRqxyU5tBJxQfcVUtMnbELwPlkUN+m1Vy/Xnl
pcAeNHWi/8U2io5g52LAQbIizsLUgR7DYpJbsZAhogR/uED78eJi02s89R0clzca
V7T/O7xmznkMKN3QpZJve9wb87+MEPLxLDClFqnvsIaL25a1wrmJm2sDApUpN9f2
J1/ZqK52OoChmHP+kW+i2P1TNPrjcn3maDP+RuEUrrvaEGBoMUcD5f2IyUq1R7Yw
4dqW53fMEdrH/FwJFacyvUH5XGu/Po/PmZkca8pjQdzVM/GZmMdi9+Ya9K+dRCdg
Ucp1SB/Bl+KsF4O3QrbNpQDl3Pd+EQJRFiqrRj4Em20D4YOXtXrQdSYHPRNoA9rm
eKh4WKJxctuE+hntP/vphIbIMLiUNVRuyDVHYyLH+5+uGrT4FDDaBVu/yYh9JeJ4
vN2ueiBdli3h7HZq7zZnJjcew/Fzy/RKidvpdPlgrINh0L9eZ+pYrHZhlamwjDOf
73NrXBS1fJAS6khjvx4yB21Oz/2YqT2JiAEUQQuPLFuKGuqj/cjgHauY3s/oHVnt
VuvpVMsP/NqDkHj5S1vAXrmeA97/vvfDGp2BE6iyn4fC/eiVT9mB+wWpDB4bWIeE
Q9xPE0wKBYBuNhKd13DyQypbwcqm7tGkThLi7XO0eVKLuC5EGHrio/DFN90wgqkM
lludKrpXY5ZePVnhMjLa4NXGMAubktqiMp5r8vyHKwZYcJ5s9QjvIU19KDmPiIjS
MInPgTJWeUKYMrP1hyyGZaRAj9XpE6dyUGcHN318eU5AElubs/xjHs1Ydv5Ndm4w
V3BvogNJg1ALMAJofrLnEJr7PxTvX+EUoUBYuwnXQKI2z46yL/ijB0Oob6C0kxyO
r38JwGuqA4ZhZqfCJs9tdiBZ2Ob+F1Z0DvthPTckrUaLvy25P1ZSBdlT7PubrhEh
SjqgoVarNFXAaXe0i5LBoVz4M3WmGKt85MgEra7CyUrM2fbANzRixPLK7WkkrLMM
8WEXZnUTMSPdVd4uAhAB1SrFIGz7oSDN8tJjSMr7HS80KpMZJYpMhOnXF/5fb+hQ
l0YjDyldsAVAt6DHZ4C30KS15TaHRJgJYWcRsgq/HmdSa3GWZ0JZVs1EjATjVX7+
Oe6VLoTO4GaTIaGEs/4BtzHeNWTK6p6PZh9BUsn6WVQzlt1EG6+MS1XisDtA4AD2
0ZHkCloG1OzNZqIrf9y6l1qGIX43Du51HY12+tA7bCShhITDXpe8xoQWWDcnRJZ6
orJDymFrDmwbilzPl80YNt8UKNDNLxc4pjChHEN43mSmwCIPQt6UKSlf14u9nAzU
iPwKWpCmIKwtnOwB/6MsG8EjhmT3TPH5kQPLV4Wi8rPwskSkNzjLeA2k2GcyLuCV
B2w7d5GkvnRzDMnzYvOITkTmhebqRkXnbnQSzTaRoGL2hS/MriMyUHAPPy7nFPt9
M4diSa9cnL+Suv3wGeggdE9Ow3DkePHU3UDsu5eRZcDXeAWURnAHYn7l4dQObMD8
uyMZPLyoIIcgOCjkIGDT46+231WXA6QL1c+7Dzoj/XtrkcGxbvzqKh69aUX2o4oh
NmHiG8ydxSWWPioul6BAzx9/SaCd13qODvw6B3NlwRrExxcBHfHwV9JifLezZvnP
AidYprxIs/db98TtaaBW3YicHNIig4Vp47NXwhsHNWFGuYFhGLjbhw+aYfkIy7j2
I5/QJqyCEca30imhYjftREceQktwswUl4MVflpGP39IK11Vh5P2inMsQVtelIVB6
mh4XChSOqgbqmkIrScqALogYYgJZN4zI24x+xFuLalQ9JAeu0KOnluSrhcJW5Sn8
D0pU/K4jklpUAgIcp4e1Wec4tmM0jDFNYYxa4YdsNud7rIHW5bpEX+ZilUZtIqPv
Wxmi+6aEigLsWalcvKrqOvrQmInXd87tx0VLOXvpSOSRZ/zGrcBRtUnGag4zW9x7
/GMd9+l9Wplmal0vbGPaHOdXjTCZxvDgvlH+oAVli7b2mGr1sRF+0EZWDsudD1k8
zvKQ+NUPQAybIG0HvjprnpqHepDXD5Aijw7AkkyctmEeQjZmVJ3dXNFlLkD4e86p
UjYjD1Y3W4zE/tlIlyB2ZRmm6uHfLzh0gYqLD4RQzwxO0IzyrYL0fg+zx/K1p8G/
6/YJlMW6rUXmLhEVKscdTK5OL7/dQZm5XFoS/AxwcX5fsAldeYBCderJrrUwM3Wr
LvgY/9ap89kLqmObeIW7W8V1TdGMrpwyWiUby0ep+QdgJ5sr7xWf4p3gx5+hh1kh
X5WXL1Nv9HU2GSUiM2BxB0lkQJCZpbe/qYPYni1dy194AIa+VsKKVXKDnmOA3qzF
FGyLYPYTCyOLDYk/Fx71bJiFe98Nr/v4kkdrQucJRjCCUKSCOqeW+bu1C95IcFNY
2UvlwQLGM4m0XEXsWJs8D6hhwT07Xo3HZ3hyfROTt2nCayPR/D1Ta9BPvN/N+rR8
FpIFmkbISU4yOMfhRRZtviWm0bWOBmeqZj5vJKfFYYA43Mnjrn4A5/m3SVT1eshu
MydUNiTGXzlzm7nA6+UEuGsW14DviX0GGN8lWezEQp0EYBbsDMd8w/mp9JIsp0LU
U7tcosxgzNDbWARVxd3KPyeYpk0ttd7W8ApRR0e0r4QFoekYK9MApN9j4m10C/MM
NWUqB6XeTk60ugGvL37HrqqtcUdhc4QBg3Gq8EiBjrriBmjcdQMuYaXb96zKnfIz
qdZRmp/5pAsxGsgL8atxiPhY/DJYgafbWGDCtmyL2pSV+yNBeTf6xZ7lvU+aboSV
sALCqxQb091QItd2p4zt+KwN7k8G3t2PXsvGVQDBbDSlbM7p2sexIoTerkLKdI6L
4boYFPXpLa/IOOlvYcu5Qheb3U9wzC0ECOajXfKwgNmtaDh/UkEJEstFznboEjjR
jteqD42ih+Z3tgeGE+Lai7vnlI5u5kRJ47UrU92enenQgK4JzESDY9c59RyTwatX
aJ6Tl+hW9M5xiRBU5i/+VyN/YZLhdwaIb1Ly0ehadd3c7UxhfBMP5zKU6p3JjV85
Bt9af4ruIdVf8p1+90mTkpxaXqH03aO67qU5pbvMp+8gVpXJsDS0nB1g+xT9yQw+
3vypzZVNnRurVgMcLjWWxdMOCG59uwa26xpH37m4m+C3s/VwV1jdtt/nttKz/trq
BbbZ3/Y+uUG8UYXLcXnqYfncgkOIVWBuDDD6BBzPKbasT9ct1hAbxKR3qOnSZRdy
cAR73iUygY590jsdlz+Obfuuw6Ps2FTT5JNp0UrVoSL81697Hw7FwNOWB0hkChlx
92w591SdkxZ3ZnXFyYLtq0ZRTCjmPq1iRZ9Z4ehrYHEe/NISgNgoN4uNmSXDSCz3
Nve6Np58u9iQxFKuRzNMKiDfzsU0t/7eyZlkaLBm65EtDSmUg/2xaUFi61DvTgRO
0VLcoBksZsoy/kvDiHpFxWZp3HL7i1c7XrMSBpIlXO2D+7sVlgkTR6YCgAmzpEh4
3cM3Hm1fnVI5yO8RT9pFum+1HhqSynMhsBqVa963xEPW7fhLxBbrEAnnaAnJPO3n
Lo7Wntc6R+3WvXonHupgNsuu+AKPnLzVJQTzK1ZQuVE1SqjEpM6MQzEMWAYoyZuV
vs1iOoROmYGGqlf0d5cBvWRRe5O5BxjwUv0ghR6oWRILllUzWFaHcGXxS0LdZzPx
d/hIatwDJ+MkXiajiebRadgyC+tpN3aLQ6ewuJnxtJDwiGfcwPNcih3Oh8byUEKl
x2JQ9Uf8VEqS1NK0j+nljQnnnfoldLVLIlL0xjQ1bwhx5uApRHLHQXXSlUjI0I2N
cH+I0WyPbSOQHlSQNOwdBPz2Ki2Ee57i9k6J0VGhhgoC0ENIVIVpCYLthCIjO6FM
4QZcYNiPibD/vdAhwMHEuBgkForbVR/e+T5D2mGhSgyLi+CWTWdzNIPwApODRC7u
iF2cINQqLKQeXZ5VIQk5QDv+6XcBwNBvxDBhPYEG6s82vHdlVM5EkrHZT5+pfM5m
S5+FO8pH1AOwqHEoreUf92/xTl16MePMPHPJ5O4MHvbcty3w6GK1659c3Gdpxbdr
o6isFsKilnBVHY+dizVJFbY8E+Pwzor2Hh93zY6mH3qCU5hsHfx8TboK5D6wSSXE
naI4BdTKZAGfV6mYXnLo4c8P7MTqOTXbQc5eDgjHU4y0c8yZuQfxZGT4a4etZbpS
k7xTEl27s0V5hJNt3+LVZx0EjM/FZ00v6oAhCMPTrYZ1ZJOggI3isG8Gfomv+hxK
Qo6ZyLDCQk829D7c0CupCPNi3yReNjBzzjAajLHXe92YHh88URI8rIpBoZF8syGO
Ej8BMHBuvdXAfz3XT1lmrpeQso6M15yeOlWHa63mM8XFPbQg25RMHjc26Gn4VxmB
HayP0zjntLfP9+5yClNIMPRaXF4QI2MUP0mOYUs5jCaUsc0cbJPKiUuRoPl5vuFP
3bdUXizUwhnUhIuUapdBnDlzTE8dRFrnbQYbWq2rViIVlDzszexy7Qid+kOce3M9
g59HoX+hFiygP3tuY5CDV6I4Om0kvBbzX3fQZi9jXJbl3jC6A5UYkpDhMhn6+sA7
EocPK2KOwWtM6jSLwWkZmEp1QvNEeV/v2cBikH/kMTnH9bGlwsMRuj5J/1W0wxP/
91lgfODfu2gyG71h/ldsKz0XUcbT6+6TWWOaXvxYcDp1s+jB8d28s4zltzJhFo1T
3tMCnx3GSAA3cIXpJuWGlxlV6dDRTATw7arWbh2qAgNLXfTMnCznK6DyOfFvDPv/
vdou+65Q3Oc342qoTgHvNmssDvbZu87Vq8r0SWbAevJFn9FFcuF13NcKSj45K/mp
+TE3OQN5v74L3ARf95co1nADZqXU+f/7y/iByUPK7NP8wlK0fjVCVsoq0NABzXYa
g2d/p0uZqQ7uEAjSib8/1QjyOtnVYE/QjHw8RgsFSJYa80tYUkw1eFiZeXNRGemI
pj8NdPN5xTsFwkV7zcPS2SNOp/0lb+etJGu8LT1sE5yNsg7KveWXFEwsRy2wWGn6
SPReQSltmb3xrx/8cqVLHxBM60d8CXhEE0WQ9Fxmvrfk51qIbeP1j1LeYhQ9MraL
uyd9Sm7CCRdriURehw+/9hfaMtMmzGr86YPmWo1DZGPlSjQ/gYIIr01mUS5XZkh+
uJPf+V8ObHmx9lLD43c/U7WmgqlNdWbZ73P/YZkz1ArViQgEDVtNnTo+x/dakvQW
ceGt47s9Gr4Eel64NuysT3dtbjkv1JXQ1JZAX1o6c/s5sbSKhmlv8b9aZMxyB/kg
42gMhqdfcZGZqouApkr1WkXi1MkO+8RiQ2sU5yysrTBsa6ewOM4WT20ftIMcAj4N
Pt9Z3mTgfOKEdFcFY4eXVtyGsM59zenyulRaUVSlzmuTLRvNKwATzDS528Iv8SId
lMVTJ22q4cFpB+ggpTvqAbhqqXwb7qtjqr2qxtrpzN1jj11Trrp4fz0zi6LZsKUW
O324KgNIDQ/QoOnL2z428PYdEqTdENncfpObLBtd8jc+l9F9wEbOwNnAWhDOKnbg
FOAiv5hP+J+LbmFd01acyN8OPssftn9kVDyj0G758TAQLoDnGxTLW/Q3y9ION9RZ
LJANlVXARb6qc/rgDuQEy/J1h3eLzO04VRG8a9cD++GkERaRjcZTuVXhV31JP1H8
qopkyw/BisGWjXj/N/IQOwAr+wRjgmE5QaZIrDPX1202WHZnSLnooRruny/f/p0/
85vbPYOz/0P7mMFIP8EFo5Y3j+5R3za6+vRyeiouf5Lwkc628eDTB2Cbk9uqm5Cr
tEucOSSnK5kZ9l6WzVdK0Du0l5auOJI+Ikq7mb/j84Di9CS8wd9YdHXS2LPJC7Ar
8a1TVM854M4ppGLk1INtXGeP68zzhi+esGksKSxgh+KgZB5Kx+gGXiKe9FB9oCUF
YKGYv+OYmQGkpHy2cPWij4aH7v6t3c/FNV4PMRYboL7yBtCDMt8t2WVaQ2ssO+hJ
CoBaki8+i18Zo07hP/rTSLD8fIcAdMb1rSeh+NB4wt88CUD/VATBJIsVNAhKaKQ9
t0Jqus80ElacrZJFdu1sLL/hreW7g9IBYJ6pUkC+OBNtEMXR0K6nXjbOKl98uQOX
/VPe9AonYf2KVURDh/EcQ5Q5b7eS8WlkmoPsBfZA4WXlxY/zL4QsdjdjxDLwwewl
fo+XRHNCS/PbP/swvzrkMFqJvgP7byTMogyPrWTMnx9oMn0yc8gG2mKYRoNQthoq
Z5TJmvjI49fY0i3Ik3ILbA/+9DENynHnnfNdi1KvfHIVDuy547Fu0Q+UeLo/7Zyy
W6izBEvpR/aynnR1YDJxv9DoyP3cI6DB2c4slRRPljPQhBCj9JX99z5m29CcpPXI
NjD8pMmmN18cCafynDC/dwrt3MsQKytTZV6S6U/uRfPtTpLcD2z6Cn+30AoqIcDu
1AvBv24mXHjgNztRXtINWj20U5KpCWylCb/akHaqOVHaX4iU1NiXOaFD8uVNL+hd
kaAokCxJhaxElQGkJkv6gnS6Jrw1sad99hjSOyo5GzNMDrthmfC/Gi9Q2pay+Th6
Z1Jj3X18c0E0z66Wr5pycSfyyWUs6P5mxWLZWWy+t/heK54D1nS/VVloeEZd1EoP
EnObie25LIE8kEkpIapxJeRiq5Um32jXYhyqiOsh9TFTRfiiNFnvvoqh83AergeB
dypr/dyjk4W2iIZHKZbGGaekUmmgSK6WFKQPARWRa+qc7DzqANj+zDZ/oOFpzIL3
pGO8IF4YDp/TNNoYLcEmib9JtHH9ZPwWddaRW0LLiukyOFXSgxhEScfmA7F+Lwsj
RsYCC6yiSQspIQE8QDJxoWFVMs/k28VZmyKbuaWVFwlcmQ8OEzsjCsMmOU4J6PAa
qn360xobWILqFDc+/110ZQC8xB+W8cJ2i5Wd7O+C3q8=
`pragma protect end_protected
