// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
cd6/1SmhLtGZNFkf9+SrlGmFdLFG+8WERXxxL9RuB1Ajt25PNVc5OAEcoUUPoGhEnGeiCbhVUZXS
RYzD0VaV9Qcq8upfSh6TTiSGDGoiA2GGKRT9Kemlx0QGZ1rgrkk0gUo/rTz3O43YdYj+844M5FcV
DM0veWwXaMtvElbQPlRbh4bayM7/QGWVgZVI8RSnPObyrI4iuqdGPNZ1FYMJNCkcLhgV1upNjglw
OPmh2TbmSPZfEmEkxiihK/Z+g9di67V7qxROBi+kVyr2U62ZXWBKuXBVGisyAxCXzf8N8jC71EAK
3Z9Zv7oZwVJE4AnSIcWlVA94fkT0belodXiCKg==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
TwCG8DTMG1B/Mgy48s5b4iIi1VAAAXZi0ZQyfP+32XIrs0PEK+Zbwzg4kCqNOsVN73iYZvMXML57
f1S54/D01Ke1z+vhz64c1/fi4j7AvSeMfVHokUoyc3USDEakba+M+j5fuJjB6FTiLINSC95smZdk
dNrLXDEXMfmp1NHFmOOcEjpUIEvYRD2WK5OIrSdIO2FweNhsez04AY6UI9xvEutXU9Lpy1aIagzZ
1Yq4CQBt5OFmFR+/aU2A67VRP8h/+dmkjfpUbTZpL0Aydcb7AVaBBbdvC4Ecx0xPIcB0CrC9wlCs
xbw2q2FDLDBKu+HOBCtcr55hfcDR02k5iHY+l38M6R16ABzByhQxIy1ssxEi6k3Q5djb2918OMoq
srcUtEd0b4BQKXYLwpHuuvciOVkYLN4rrGCQndYW/LmKlvFj6H2Oftl6l0sBG85BzHX+tpVPtylN
0Jzuwg3B08jqGjN4L11MDSImp7kQR3ioOirZi9B/7yKztuZkp2iXTpTMHIuq/TRNdJyteURdByX0
nFt7+FQ1jwFD7Ng9tHCwHIFrih7hCbgAKqc1q3CvPHdQjFXp2HQpVhDdhCxFGTdgMpS3IYBYh6Ql
KySnKI2Zf/9ANoFXVdKalLTqbcgeoMvDSBWXqzUR3rU8CDRYKV+sCX0oxylC4rN2YYxeldzjjNsm
o+c44XZ5xA7LL6spb2PlSvk8LEkgBG+Tu4aacCX6G40/uHk6vvQJDtPiRhyJ3V4S3ALMigTkKDaO
p8/DOWLU9HeMKxfKLyGI5pUq1/NZ7YdU3EXTVzH8MSkGEGemvoAAcHXoJJJriwU45fN/0yYbGVai
oUzU2h//H5jU+ojXlWaXwEj/60PtIlMlTL0jS735Kg2jE72j77by5gvtxL4sh3Ok1rbLPaUP6mAI
B36CHsoNR+V0/CG5KBPMmgtgjHMk8dziGWrc+TBE4siGt1eBlEccHsb0f1LRW+A/2PKSLoSHWRpM
D1YS+K/COdTGm71fDpFemHCFwEGlem0fh7KUFubcGTEWfI3Gz93SIHdXsP0PRGIhQMiL+fWNRDtW
HgwPc/lJVG9tfDqFw/RjkW62hGi1M7WPPrgEcfllwHFsJLMYk7uStSPumTJ/hDKL4j9/uyz0tkIC
6hSLF3zGtwzeS4elm8+AwAQn/znVkdCdEa6deXZow2hFacrnUo8D6PS9Zj8ZPagX7D/9QRs4Rlwq
uyescgFurxXIjhQ4h/gp4skgjFpSx4YgLjXbjl7522FRQirPnt1pkKhwfsJTcogucmfs2Tz1HGvz
pfxZ2vzW2CkJJxQ3QIycjN8ZiiezvVRUQu/S2oCQWecusbiVKaVVm9AQw98TBpnSNU09NEvMvKlf
GKDagEk9JW+pL+sFkhUmMfbStzbLKM2GXcFSp4m+8IE3aYlj1kqzf4//MYeA3RgmAEZTu6eVvVbV
FWphsqT1iDqxhGHlblZSnu82tPFf/nDPvhbYx284D7E+XgfXnF1mU12pskIDnd2Edxsxi1PheV+o
hknXWNC1LGT3BLdT9c9eE5dnX1iF7zjR8gFj/jLH+V9DivQSwA1lpOfb2A+i914MpOHwR0I4fKpc
VjSFxdjC9sN52JJdpusHWiR0bNkEpsSGno1JfegdXgtii+DqeDweQKJxfm6ZSx79x2rOAyxb2Rel
FrZfLgPYXjocmQJM0wG8b0lwEEBlMqaDx3+h2OtnLdCG+4HqUsKe75RtZVR+Jl3VEnNbAlzJydAb
xTrJ2KxvsWlUlsSPvp9oGGwMugQG3uO7qqORakkPHnRH+FuumWWJHv4T4aaHsJAqy13A5elnGzTD
dNbCMVIRGtPU6VkhhKuCT9qciPmfiWhGvoeOTXmHpems4HlRB5l8QZI+Tx9LRM1mndDBMQ9Arlkj
AXPS0rr9CftOUIv1k8P2PQ791qMo81g7iiNIPa5q6SYNKfoxk5BUmfS2/PcuzyMtrCGN4ru9ncsZ
Ar/fCJnlCS0zbmVNnbP7WBxLXI61BKjwU0+XrQSuVAO4qcnSRghyMp//5DiaksluEGOTqrmslOIM
cHWToFSP4FHU7NgmoWzunOFQ7Vl03/6Uzrkq8Xyq3gN1IzmcfByEKshr6OSRItR6E3jjjU6P1l1Z
tENN4VEyFLPW06cgiuxlQ0L6DvS6enxBtYMm4DlIgNIYDWUmpC497GKSyfX92UMhGCXl17M2JB5q
L1rimuY4EspX78IGchPQSdvbmHt8Juhb+wNAfOXyIpLrVU9YPBohLI12SvZTZJVs4rYjqPtKelXl
Y0fPO2BHMEr/rQHcvpqpXX1y7oT/Yhg4nFKTQgFR+h3+Uk49QbyCmwRvLkMa+o1hSPvMMfnCWYvc
Zb6RHHhd4CzQzgkkFbk0Gjz00qtrV67VrKd4rQWJQUCfjwI425pwDxR/VBkymHLxXEuO4wGK2Q0T
r768v9ks7KGDm4cxLdN1CRRsruA5G5C3BESl4YlUuB+06ELc/SiYNp2Gh7DLpFRa5QErKBzIHAh5
/bfW86k/FypafjTa9u49LnXcYfixmkh0vV9lxzxk1cdqhDI/30QIAJjM9Spn2Jzai6GnG8dXWCoJ
ww8oBGlYVwnnr2ashtxxvdBfeSuqAoPby3KCZEIeTTI2RU/Oh31ixtxUbxliEvxxh19QSAW7T4Ga
7nDO+gl39xiNIpm5M40/2rGkvE3eupg6QLKtZ2y+6nXZZ1/CRqRXmYZu5/KWR4eTrvKTM505wCK6
7Zu9CrW71pGUA5ed/RVnGER43jw58m8uuAWKB+kDTkq3mQhSAVVf7vtKW9aDJlNzStiHQhAM+ggI
QJXIgSRpNfxa2EHFtM4ETrlKI5npVdTuJ3Jyb0VmfsbOOkywxXnPLwJ8DEXcrKEG0I+g4iuAcXgm
uuNz25wsOP1/cBQ0cC9NrSTQLRsp+9Epc40iqopbcZu9gZEssIRlMfKOiAJVQI0tWJIf1sLumKWx
AvbvVf1yypiO+r0fAJCfX+3j8x+FHIJp6MJRlBXtgcqo3cocNNROgn95JaUjlWGtrgJDXpNlnB/K
dMrxMOIuOlPk06iFQzQ4Hmv3+TINyyXcEthqbtt1MQ4NKS6f/wcLzlw5qoFFVaaLRB4ocqFFQ9A9
GJdWaehQrpq0bh9nXJWvR5t7DpH51DY8MfCqtoSEOb2OFCABjdxX9if56I4Za2qUSf+4zy2dxwxf
sef12IdE/zXVAatxrZ7MG5XMHY02yVY2E1173Ny2U852Sf609vAkf6/4paUY2WW7ygqSueohDepl
EHgHnnHLA0HskLbpN6xgK+L5LrZUBIG5+4CoC051Ne06M8tCz6APXKl1hI0C4MHiYVjKbBxeR1iY
hojWBW3hU2J05ln51GJFWNfCWRa6R5oWY32v7lyNhf4iE38sbZTyRYsrhZaaHs1m1XBqKAOQMUWa
Skdh/cEtEHOjj2gYwZuq8EJhgy91XBaPKlMrRE8FQ3wI6boY/hsBLHNyKVnIHIEmP5AVksYcII8q
GCOj6m9grmer2sE9kvfRh+4rs9Twbc7Bwamv3XoQx45H4Ld3tSFtuQ3Z2Ws6yeFrbrrbMQLcCvv6
PDi9ilDONgB2hlDgNyXI5+Wlb3IvI0OkYlJ/srt0us9oAt8bmdXdoS3zGgURDON/2TYkkENz33dD
BGzTpzw9BtDWrnWxF5XOjtNzP99nGN2Xrv2Hq/FSLV7UIU4wHnAlHgV6AqSBeQQmynFFmK8LDK0f
NyNLCmYRblcK5Db0CoxZh6+45/m6blS9VidR/R9BXoGn3AK2XnttyD/yXKLsI8KusNXlx1KGOuia
i2RqUAl3n0CQZ407Evs3yUKQ85E0pd3NQpI88YnlNVpx9VAvt2oB8uOGVt8eDn/vfrcU4I7YgLwc
jl1+QtqeX9IXrOf+lLLeecshtWwYFcVG7RweqcMJ0FIQVMaAHruMBoZXAsWQR4gX1CQjeWLkqwHc
Y8dUOskaZmaUx+xxSdVrZe2eIE1TCR5DE/GUqDEPQx7c/qdqCMOMCETI2bdXhA0MIQZ+MvHsL6gU
cI5zrUCLW7Punbdz+l18AGkEw4ElLUsyQ7fv0ty9p+g/ndWAqanPoZ1SbsaIrXOYlRR/d2X4XrpI
n4SWxoM6CBsploiM7n1/gqxEi0D2XreXYqu+P9m0P2Z3JZBW/HrUkC3rPEcFHq6iFeHCsVOlS5Ug
tT6XfrJqmWS/yM4X113y0WWDt0ye69yxPtIwfyEXzME+/Abf8MMZvvNYg7bZCT9CAZo0WVQAQOyC
UJPgXwOJYjH+E8DjF9Go6GzeSOWlPANePovS2pf/xbwvM4uvXXQovhHA1RGoYUTRMBnLlfGptBtx
0yZyE2a5lN4FqAw8dvP2hm2TIO/dk0aBJ5TJWZV9p/5jd1tcShSxQ4SdtY7PUqUflwt8OEDe7Lbo
T/eu5xDts1WmYDmaWfaX6w82osCgYqLRswToHj9CtAgBfhtH+rqYa512HHhhauwrIqnS0qG2PPU5
eILpJ2z4tEwZCiSgPob8ZTJPItsUDE3+f0SwA2Cocl94474tE7G29kLnfhjV6kwc6U6xmx1jpK8B
lUVyMayZqp0w4Mp2xM+e2Hv+iYRWwspwRVo7mT6jNhWWIcW4PhChxllk9pTF/2Hz0EqvidgzoW/g
jXeKnHBLhTob2W1UHpU270vCK1Z9fdJWiyych6ovrlmz7hotyl9VFZPJCnLYbwke9KTK1kbAqJB8
2XTVdUl1j4i8aMNLLaKbqa27P4RZW0k9gRf5QQ84dckYPapKY1qLHT96g8n8C9srA+LpQ6SBw0a6
VeLAL8IZCB4KhyBX5MzLNpO6JhoAaFFgal0HS365Oy/a2VsGQ92JG1ypWbEAgt06QnRvkQYJcESz
b3EZSp/z03aLZNqeK7kPMRxsYWLWt+uK7MbmVuFHFBpRjZ6oihi9eAwz7+Aicopib6XY9P6laTKX
soFg+ItUwnx3DOyoQDHTQBPI4S/TcZaWYfuGuLsWLnR89ypmMVYcWN0F9OVy3KHKIs31yF7qticw
7GkWzrDkvzo8VGL4shQPmsfhxJhhhMi/UeQVRZzxdNovOpnDbkQg2MRXrC+fpVq9rGGaPIomhiJE
vfJ5DEddP214BwIVh39D/RRz6exUx9t11Qybm+pTu/Obc4sncJMHWh0ccFZsCBVOdxTOqGE6+P9I
s//dr68qJxBr/HrC2L8Vlzi8Pg3AXtyFDTJaMtCa5gt2l3YnCP3oivCwgudlWRKuigdK5V0bvYSu
pMyFcIHTSSDom1sZc/coY9mR78MIKFHn5pZT9WakIGWt9XA3QupL1xPX9NqnWgKdn4w29z5ew9A+
y7o0rzfa563UpzPKOvCtOnOyj3nzszGWdRV3i4gC9NbAkB8NGq2iDbTcawUjlN1vsAwXF+jKDrQJ
TtLM1l4XxzWoBpcMSsVVQ4PruwFQDazHo1EWIGMAzzSSIN4eKeoYF6nfD0AH/d2REImonTtPuf3K
WWBuue30TwWA2S+aYE0lFux+K+ZZ637Bf46m/bZlnPPNhZOTJP5vgE8gGIrpev9njI/R5HLgtWk3
TKsgP1J2CGxx+AZrQthZ3M26nBeaiZ/cYG6GX8ypye+3K1hYm2uIT+nQNgge/mBu/JzsNfsM7izm
NT/bA2CVdo50pijsdmlXjRk8qHrxHGwcxXR3FJ4Wn2a9jK9fCJWxD50Gc4y+ryb7eeSluzplWPnx
bOEZhF2ARtCUAWlPdN7N+lyEeSo6j1kk6GoF7W4u50U3YkV7QYP/uuTARlGm6Po05w6sV3PTGg1e
jdDSnaZ1kKhNVJhIbQUSeUlNn4v6wKFKjg6PR2hi0RAHCuE39aFjKfU2zIqSwqCa9EFyNuDUVihG
p7IRFM6ALnXE2bQrM6x8Yrt3+IhTbGRMQ8c5SQTkrqD1FpMpQ6+2XJtEfZs1sfLHUhTTkWNkV/pW
jle+BsH/AfNn/Ni3PFm90ltUtC7NGXBK/3kK78KizIRpZT7XN3gb42BSiQn/x40MNL1JUT7yomHk
EwfBQcDbXP1izSmDOxdHFI9HI8JCxgAki5g+xuwPOLghwYY8uhc8AGcOiU3Aq/xlMGsWdOeiO8IM
lJhzpH1QZbZHqc18Rlkk5Sw0wIOzZlTuigOx9JIYcuBQ/OSvMudKdoSODQ0nDZubSfXTBDtjWmgW
mqyhZouEgqgWpclWlHF/o0kB/H4WS9IDBbi0QXE3TnDwd4hvzaCkld34MxatU2CAlG/Lzu0fylBy
GqWBmQ1SsSpqOjBVp230aeCDaDqyYab9iMTfLIGROQqJ7MB4KWRi8IVhvHre3IwFAzBYNr0eqXaG
1BX+hSJNku6ZjCZ/wFOAcHiZMk0gC7pjrEWuLxQqyuD5iSF/n/7YhvjLnRCuhBF+TXMa/3A8YGC7
mUsItdbIcNmcYSp35CXeyMHSbST0mWwFdXGbWEHRc8AlY4i/lxqj7phZZWRI7Zn2R/xh0A+boILs
+L0IFUJkIO4umKD4xfQTdJsrk+uy6j+CSjCoPxiLl9TRT7Gq820BEwzRYkzeC56QZXRtEIpDKriG
y+9fyOXdLMuS3/jP/A43eO7yk/OMn6oN3ame5tTTB8EaNWDbuGHGiTVbK/9Gk7Y8iP/wxEXYKpbY
Vj+2pHwYV5L8J4Igm38K6hJrCRQ32lXJpjeU59A17rMact4agdfZsDFEAXuumLG254Gb1/B8EK1x
6OQ+X8aGvh5fsZML7WpNNbLKJFIMOg3E/qmDxn2elDGcgHlyFz6jG3Db13AXycOaYmACOAoFS+9E
qq3HbnjaYUj3I/GE752UeCtpmsG7IxoVeULADmFt390Ai/qwKsXetmWUDza4jqFToXrjlzJZYyYD
FWjynp9nIo6j1DQLO6ykow8HVfQDI+L/RCmxjYc8AQ7QySaz0gGbb9KDDGdSgPDv0rqCkx8adpLp
pT9nKarv1nCa07znOmiITnfxTH7FxG9TMQGKlw56SlXlmyo17bx+gaNso7tDpzUNhF4yQGEr+pMV
h8NTrt3etKlgviXiRJXr/kg3yNfkDIPonDmR9Ns3PltfIv6MA2PGmqpmUQrQ8Mu5Os1FQn08LVnY
niDe7iyNWnvurT3AAt0y8zuk4BkkIEKhqUY1uDGEqVrRUOqImCtnTvjZ+X4FxfWUa3qK+NUGBdS3
RFOHJuiKqCja8DiBtUCrxJizPvZcyzfZ1OKP5kcAJ53I0TnBTFMQBrigliGJKIoCF3dshUSu4OxJ
GsKwDDLEZ4+rlPChRJBQjJCXeaHdp9qPBEo2rndbLVQbksAO5dxzhThmrTMlCPS7OJs8OWj2QR7x
otIlBDJdgCkxPAYXfFu6LB7iyuPmBzsRTzJT9I7I4ZN48SD1q/xSVaw/ryECvVKJMk3IQ19fE0/6
NICtiGkBrmf8PQ68gE2C+RgBoYXBgsY926QsYoc5NEuE/V3bR246EwCRC1ndGTppFT1IkHSXHpyt
hv51FKDhS0RWMYFKCGhHK034l4CdN3EYJr27NhHxIEhY+eMdR91I1zLtAhCfLcz5zzUzWgjcI9vZ
5JootDHzWsp0Sm2Vsdvp/CQViZ7i0Edsfb+R9zF53Ns7G3sWpv2J56t/8qKG3iiCVuVNARLNnXHT
9DbCznXkzyOe1vlYS6if9qYCL6b5zjYb42F6wMD+iDbhYZm1kvkocBulpwcgDBRaA+9oFl224/Sm
VdMCNSWXPkxzKIx2xVTTGx6D7uWIiIbSdkhffvGrSWOG24BzpAgTSw8/P363Y7KDPoDajfK8BLMl
Zr0mQXO37VOpKeSkZyv8PYL024xvhM/DCSBMY3u0FPexLB71eqnDiDjEAynXaIh6915DhPhGkaHj
rQH5QXL424JfPNSOGgRxRVWbq/Bb3RZosojqVSIo/i/9fN4Ow5U+27au+C4hjHBRNRkRxDvRNevR
bt6uWi1xK9xm13wf52otu6N1kFARBBkxCe+BBTFfUs/uQJ5YrPwutZxZZKBsjoO2DGlB3FQ12DTU
WTVX4OaA8v1XgvUpZErdda6Vmi9BmtoFfXmYTSTnEs4Vc9fuXUgjOgCRTycEtjgfvjt9jHAjEr5a
Op7oSqINzMLFNgzdysLDH3/mkZmD04PrEolgiRgaBHDfsBqjPQ+/bpC6Y0l12RtlzH8ZR2kJnKvA
Zg+6kAc6Sqz6GQlK6LUYFMDPcCf9yac/OuVTtJ4QoAdYKgplQCHxgFAo1rHmw22a3ZX3z+9I4Hac
R5TfTm2GD3ETNhoMn2JTLiNq2OgUxFKZuhYgq8sYaZfHwGlXzV7SB0gTbVztIf0WMbW5yMTNj7AF
tsTHoAePnxYCoEyTJpOfKN2EehDAimSLjb0IvVyD1eDH+Y9kBvYj0ePz9l1+GXt8GiNGmB2XByNd
+T/6h/4tPxHh7ZY8yH/MV3pSNSasQYK9hK42Ejzs1CP0Qnp0TRdkINClVAFT4nc/XsK+bMGOcrbA
HOjU9qfU87nTadLcGIypO+CFexvan3Pa39+imUUjpY3pXVDWbZ+57lEvLQ0hGfvNJllP7DuoX8xa
9eliPpM/f5hGfg/SdT673uyazRSHsJbZ0io5AY8kDCyFmEG+NfTFJkT7cNqzj4FK9tYUVnpwKxbV
jS6HfqQMe1KQ4rp/x//3D9lpH20KLekDPsOWZFH0gRVRkQP48j5mwcWW2HYBJuHWkbSFoKNACyME
4wJfcFbC7rZ0ioSmhP/5II9KpnutdSRmCs8RWwafTb88l9y3DYbHHdsNtE2epl5miMRjIjkkK8XF
qo0PNb+iVMoIRQ/S8IkTzOzWu56Or8fG2jQ+VDQUGOkJxPq+tITPwqGMrn0n4UltLCYMh1sUvD7E
CQ2HaRPO6CsrZ3tyhKA5BSDrZtQmIHSDdOvq4yHGfKjxaG0leb+w3WIlT5DlzeWYzMfuX3i18FDA
mIpvnTdAdNf416JtJyD7XEbekIlfjMWeZyQYzb4xhAJeGzukUPqkMiqKhP5vozJDOvvFXcyyHx8Q
h7PF0BgWiR9N77dnyu3bezGUIy5lzwhIXDoOuNUIAk32BrBED4kdHvxe32onGizme3SCophGTNI7
VzsCbSAWtAMPYhVfWO+UvixdxsHrLFHDe1tf6bMW/lnX4+Ed1xJ3TSSkxMEiMcKvJnTPN09xM4Pj
Y7AwRkB3aWdXPQ5fqJFdcwnpvnjrs9nAo0iM4OA7hdTbc55xF7YsdT4Yh0y2EWHTKQTtxvZwiWWK
jvTSUn6K4Bn2XO1ft525RI9Cjchf1Z9BYHNRBj+tE61qjhXktSePcDB6+Lpzs5wX04Ir9XQUtTsG
IsPTaPFYQnCs+E17FIzW7DBJ6/ia5qqvoVj54KvJv/+voBQVQqFAa4rSI2JoNLSajI//wab0DULN
b21/8zE/+lRcz/GJuDcUOPIuweDQcLRMm17NpqO9TIvGMnNlijncK8EMuTSYu5ZcCnnBtBq8XINf
FNbp6XbTLWsqxXjX/3tmGqhLEp7uSqbCjamvxCXtINdMWw2IsiBJ+xQheKX8uGfG6bk5vHXwm71x
LjThRO6IBsBke4G4pknFueRCxwRXomjeH721OwHSo/YyTumqoJR7+6nqpPLnFNVzVOZz99v33/5R
HHB9CwNP8NgRS1s1bZfDq7Nc3wqRNoqN/0h7KWFfm7fhak65At/6yNwFP/onCMwQYgYD1RkLYqqO
bT07IskwVB9RZSnjhJNOtU2WHJQ2VcP9sByE29Px1HCqHMHb3D247DxeTjR3WgMmXjuVQJQx8s0V
Vsc2s0Dj8aLAFWGIV3dmqA8XhFU+EBmJuOftaOrrUr1HI3QWp9g/6hEQINUxaNMlvedsxRF/z4ev
9zfSACSDxQSbgPh+F4mitSj4Et6EweciHDr6u83NyATle2Uha7eyRjfGuwlo6VvfPjaZey/aJAL/
uHQNVOsoFl/k2Y5rmw3gIFdcNCE2sUo8PT1sRcli2Ca3bFBpbycMxt1OrXjHGtVIGGEnsFwbSFQe
P2e9vh+RzrFh0eMQoYmFTpfyFGqC22cQOu63Ku7N0P9k43oUupMbtWECzoMjlsJT5SqYkYonblLt
b20K18vKvBKw2Sw0Np2Nx2LV+dgo2pTpOlaGf+hTSxPvECYYhhOgvucwbKB51xaZ/w1kdrBrhnc+
hwRA91b5dBNdnLtUXuuGHPoQO0ohmh0OJKby/oHWbB6dhoRlTP4uytELQRwWG3dKh0/xIsF6fxdQ
Uc8YPOcwFFoTRhI+FeXU7IZzHpuPbGWJJSyFhfKCtzbKDJBE/04CzdyGdLWcDG1SePnQZ0DF5Gy5
DMu9bh0hxrnfamft391wFI22em7D1I17jNasFzUBJ4KEkRFCNySFaazubuRsILR8fk1GcvSR01NB
PNI8HE7zoK1SKs9G5Xy+UccI/ihXd7OcdRAvW7YJHlDh/2mAAlB/Xjc0pqp6aQXtPt4ovBD9yO75
Ci1eqDGyQ3IwE7LrTvAI7j2M3vjiFt7094/3aNQCT4M1j7Uw59ekaTdHrd8fY40/+n/kN08S+k9B
iwhiOTbBt9Dyh5v9D/SN7iu0uyqGDBX3MMjCVGb/V8vvP0J3s2fnZDxMcq5GxoXGBiLBeTPt6Ifo
5D5KkdGavl25oI1P5oBWRHdTwReVg4JJC2s0mltoeLrxOIGyMo0NECKXVvXUX4BEqRjxYbfNuhd1
2svB+nwpPowHKehoAP9pMyheevfy4/aYZC73WBdAGKGyOpyRpxLwoqqHsx2OY6VRXSf6HSGFgtDA
o0rR7bJ31S4/dB54thHEPNyP9JF1ZqbUSAthhSdjNl4ZiInGq8Epb+tyWuJMKdHS3K2Mghusa1PN
yFuQuiG6b4FptUXstEjyWKeGrbaKVXT38ndi4acsPqli30+ZEVoW9/+2EZg1Wx+z/OXnBDxwW1mu
+G3I5dhdWUubryh5kB5hWRQ3nxkwSuYt5yDoIB8L4SgfIqlEV6Z5X4hasDLtQpQuTU2S+drkgBEe
I6K9P+6XC3NSQV86gChbjxg8Bq7ALhY/qQeoA/Owxg/xjfAIW0QEwmxc8wtrwQuBE6+hBrpK+3JX
DUJAlHcbl371VrPI7ojjF55+luap1luPiY7wtDwVOnjlRjhEyWMOfyd+Nsi1TjTldqkgdMyfRQGQ
K+4KUu4vJK1oUNSw7oY49I6JVBbTU3dff4sorvCFXSm2934yFJkFitANfO8YovIaFdTHGE1g9n0/
+7JFLOVkY9AD/ciHWdPMS9W0tM55T4YRLeDl5odGL+o0QVkVpsyvdKJTnVjwaQR3c/bDLNPjuMVD
KSruxiz9s83C5LLKB6Fq5nqlR4VWz9BXVF6SS8/44mm4YlzMD2QesfqOrDt3eS9boxScfCv4O8eJ
PWLV0xxMdjkOBaGPNMO52rRlJbVxl6YzG0PyEV4Y0mP35O/xzfgCKqcFjDXQFKp+HGeFs0jrRiOr
9NnicMyOtcZlzNHk/xbopBfudcVZ4W3aj+O9592zZtnh1EDbjn8Q5vsxJbd0PSkLSYT2/gYYUHlM
Wkupzsw2PX3oG/I+jWbMo8rdJnb5GgJe3mYtyXsvGZhQ88jneKP1iqv+Vzb68Jva4JYmYqTEARax
Z4SMcK7FdMpCekRtaFGUIApwjBBfwhBHmHozzzw2VKBTkjGIyrvKD2NDTtqKOcytTrpBV/0xjUYc
LNvnCQb8WJi1YS3xHuEj+Me2smE5a0lMxTme3jWCDU4fWviFgSfz+z/QmKI4+ozmI/qmUxRsww8X
anLi6+5iZMY/GXhiLRrot3Fr3Oj7vkdhb2M2VlLyFzp7lFD7GmDKWCRummiDQoX8F0aZk8lMts9L
ocxjYS5wg/n93h24lgh2sXPhENo0ZqjyUadzuXy8MErRtkHKB3ZtXPjbstkkmC1GkfEzNC3/+f5p
xXYW1AA5utFFnSE3NNPtoiwm3YGgc5bsI0l7ZLU1W2H6YG5X9MlfkL1UhZfp3Eysa6hKHEch+4Oe
Sa6cmyk2p9T1YWOzToNcDKpsIm+Uhcquq2nSF4TZ/1QglMLqhnfQZ6/TMkDDIfhZOntT0uYx6cFH
CXJKWmI5HopCbbUgIEpkMqIqDLdI1Xx1tiS+ymAD6u/1CberstnHwcyX//wAOqdfelMHsZe+QNdP
GrItRO1ppVOdYAuWErCFpvc4EFCDxQ5kbnt7KgjfT3B/wE0uA4DgMLZoCiOgaPdV6M4lWFWBhHUL
rOn0xHLiRd541dqIKEm2lLf6GZhL4Tj0ROAoMRWnm16/AJUVyF0cBm7F4iodvumzJfUpS2RYwwis
EMMEBF/gDQbH+Ejnv6yn9UR78MHqdBPn/MlF1M3JhBA5Jl7rrDjZza3+oynoCAWy7HMxaB9wg0uM
e3XyYYFzQEcNjokj8bovrgMnS56eSPacbC9e35BFvcGPUC4zii1LCJo1Wz8WeGnQwQOQ3MD0QTDy
96qM9T9Mn4p21t0fSxFcJc3jmIq/dVfU7WgqL+3mgon5dvAto30hg17Sm1wLcTRtPYwHFHx4L6ss
dPsfuAVHVWa3iYOpA/l0OhtGJGpQOVAebdOHttfVAmYFyvsi/BzDj3EOf/jY8zqCG/xSbIzKAT1p
eF3R4PGnW/CLJRGQmq8AKk3TiUYDvo1cVxBhfQSrOFzDvRU9Ud8F8739XoQgL0Q20zeSiuxRqhey
3kmJck6xuD0luL2BTsEqercQppkCAR8P6UXUw2zs0QsF1i5E7CdGBNJqAOFXipqhqrhVh48lBEWC
HJKbTsS9mOspLc8Gw0TiAW0Tm0bpE/wqDprg+fTJxkT6Z+bbmYeyotJDDVrg5o9HSIIY8ccAnI8k
PKSeFOYM0bmN2gN2rti3naN6XwNWVZAR9PcKC1VO9NwXX0XOX6W5vP29QcD49MH4a4/L+qUBaRvs
8Bpm9St7OGwEeGXJL3LzOR6UVV+MndzzGsTquLNdZbK7nv15w8VdOC2KRsnBT3zpvpXPEVX+UyMO
vrShATkcha62hFT/kiB02QmHfdtRHrW/a9jBmJUIvxv2Bqhf00x4m12gPHtrNKRGc8E3zLRW75Cu
yf2usPUcAc5R42tZ0oVM2pUlCUdM9TZLzwainZo2r2+Pe5ol7fdiT7D+0l8Z2a/ukS/+4h8xUle1
6JZrK6uISsGDKUry8+BjKwfoQL7PHpjlSTzW++ma9MDy1g/dRyj6M98GKYMluLed5BPI/T+rv+ZN
QiSFbYIZoVjmBQ3BQ3+PbB8anG1OrN7scG/DQViQ7CxTDOb36ECFxn23dywWUno19USUEkVFJl/5
vRHTYSIw9uCKewIFvT+LBgX1LbkTl7TYTgbyzwS4RtGkbOyTMntTV5AUvHIppmfzglns4D3xepTq
LNSube0fpZ834Mlq8GV3O3T9RtlxtEzGXft6k+MhFGyI3VE74GP/iwpXVJFEKQX2YS5a7U484ixo
57S2cJ/KuOrkFhgIX0y6KFp6qRJmYu79LGhcEa3hq/N2qbtoDOD2zMs23ZWOawLLUlZI5Oj9ON0r
x+7V7KTNwxeNQmxrcFm1Mnyzd3vOwq2RwjG+GzJOROJCOS7tJ+ZaDo2wh4E6cIHwF3LCScIJy5Nt
x8Puf2LBCGja+Cflgu6oiCYdF1kzqjLX/k2Uybh7jn23tQlSufG4tGNXH2xRwAS58cCwuoGLjzTu
OyAuJes9Opzin3mpBHz8P73+wRCKbIlp7O5QZIpZyMK9SPTFfx0sVaQdyVQiJUPxF4/drlVaB9by
vAC4Rs/7KQ2CkhDozU1lKfgQ2XJpNtUsWTeikzfTuIPXb6ffK2Wsct7p9Xdc/KgqE5rsyxd/ts8C
PnNG0Vm4WZReWUfwxCznhI9BNeXaILt0V1E2h7nlQTUoH28M7lyuj6pzW3Ghg+xH3JrOrcPlxlZD
AgcyM3PGHhyDvDJsDjiLTfHftdRRc9KWhNu5YacEqRbd9KpcbELTLpIQG9APCVgAjFaiV8mMQdhf
fOav6vZecprxGQZ17U+bfivyIPPfDkdMSgj2c59P973Tbhv7rkaxx9Yz8ThxGfKpRDbQ6aRjU20Y
hDIzc8gsothzG0SmnuSwO4+VrWmIuEnS4d9eNPVuz7IldNZF5P1S+3oWfgWYuJBy4DeJs2hFK67p
HX+wSL9YA9bhfxNWgeb+X0zlVwScJPz2pQEBFg+Qp5EycCbST9X4W7A/BMSrv4oS+SkUQcmRxBvR
AKQEp2X0UyypHy+EqbLfpPlRCegcVam1FrhBR1OZ7PGb7Rs0qC6gw5hBkD9Fkf53lLmRsSu4lsMT
26B1/rxhnQ7jHPKQyTcejo4G/ERuPgslhuj0mMHGDVkKL2QEXgFx42L2m2pR25e1wtLfpNd+VYZN
IV2jIdpCkJBMpMB0XDJWqT3Cr1+9y/a1N1CqNptIf5vf/6B42+wYJCPZH0G2q5YRPITArOrKz0S/
4D3yXY7SNhrtxHPbJQpk+3O1D5feQQmRbZPA9+10EeHhG3S//B6jKRClxpWM+xKGOEKFYDmH+aVL
D76DyZvIuiWzHRRdIrEb/Qz95U6mzqdhX6aMLdnY+kYN4xVR8+XXz9KTv484pw3U4tnw3eWt5Gfq
A9FevSB3pPki4htS/yzvGWzavvGZh1L0yS2hkD1XNVxNWcxccUcpWsZBb04BLGW5um9mz7cmeZ0J
UGQrSX4ajUraX/xAgoMCXbM14fzgKhl7Eh+typXckfifkcUzmKZHB92+gLmcSvB2uPi2F033/6Mq
0z+euG4hD0zNsEqstqU/VWuVOys35vZOqzInHiwsw2aAuHkXmqgcHX7UO6mjpcVKV6/KCURC99g/
wi+ubIjZBMOipUvtCSJvZSnnCbcVW5J8XR53+dvv/OhmHRYhOWmMPKa0HXbynL+c9dG7GRSqnpqA
lGwr4q4VX0SVG8S0mPh+CqgYgL+i91DVbfkhcGXSo1JRsob9v+Gopa87178e5t2OudIbUfQc1F+d
rSY8dyQdwkixU7jaCeQw7CbM4X9LILQ2EYV2joizgCSRyeUtyCaafY6BV05fFoydAzIkSKP42B7U
Cs4nfHD2+ZNGSOO0OLgcfk4QRXZmoJo0xgzj71G9weFSkL/zZyXpxqOdrdZJYmaWNgYfjdjZtjuZ
jL9eT/xLOk+MxJQ6Wf/qqvmQjn6ZI3CbjJawb59ui9964KEIgpfLL/LkF36whnRlacO4ACDfEKi+
/4p7Jk6OcnORRV2e0rjuWsPCJdMo0EHowNvWEDXTe5tlzavh1gqd17X93TpEscsm6cd8q9yDEBom
DTwwaALfNnEVkYcKkC6QrbcT06V375y5dn0wxsKXovJDaNf3ebmUWVcx1xDpnIDpsyesRXdug83R
/l1XPwLg0eB78Owc5qn8u2xhxGnnv062TvROTpSi7JHAY+LC8qK9khbqLoVHAzapQpwXExEhRkB6
msFMPanNOkvUeHDplOytqGtA5Hppa+W1EBTzegB3pyiH7UwaIo4zyfNj+hwnqRXZb2dsTFC6kU5Z
dK+Te5zwWsnye9VgXEW97nUn+C3tVpaHkjZYOlzu3zxNXH2Yae0ONrTqKR1FDvTD3FilFYHMgR9i
yMibeAi2U/pyCu4SkrjAJ2LHR2D+bS1kDQvtqJFIUY6X2r5fwFQJgtImrMuKHMk0VQb02ooDL67+
7revWJGHGyho8+l88kKuJVrSYM4GLmgElA0/nq999YLwZQSOs1yyqZ6PaASjMG6/1uPS3q+F8Xsl
vBduw5tIb5y4bOdXUBzrzjc1aWqRiPF4rPplS68COx0+hNphRi7XzEV5/UBVyUAVelEw5fgsdiQq
q0Yu6Wo40RqM3qPPEtjeDGBF5KQbyI0/e1Xn6Zvx85kTOSpS61efAL2XkMZnonQTadvoz2JzKsX/
n0UetxakWaC1zTqDvHR+aTww14hYJWRX1jNfN+jJAryy5ZBNRSf3gbOO7dOKOCBRnWEOLJlxIXiW
71sW9oh/qwr9H8fOmEm36V3iaJOVGt71gZTwjWOh7Ah/HQGbwckHAOswvkMlZVVjaZe9JvnHmCsk
A7JfrqIFpw83p299lxxor/ZkyXt7XRfs70PCvT9lL7lXcf5s3QCP4i5/m9/0OOmNFeGKh7uXXlkA
6Pdhf+vrr7Pwg1SWCkynNMJyB8HkSCv5FuppzkpE14nGGSI+9hXlDrl5TqTyrdSOti686wvLdCGJ
6Q71u/ARqUPFKx/HiaGcAxswT+usRKLAFJ7zD8Og0WU713DDpQybh6o2Ou/dnrf/Mknkdc0cLDaU
+tKzUEZUZ9yjcrf/EP+Msnw4o5UdLH0bonZy8d/bqxhx3xjXmeqszuR5EdS5tMOxJbAC1Zauj1dH
P3Ne2WDxSVpwGxMHM6I4Gqj4edDJGlbqvb1XRGhPVhErduy7dcY3DtY03Zrbsetu3UzkCbRa1aV0
rAAy8F9Kf0/yM58L2vhpWBakSDPRxL9eB4FA45C/FoWgR4rjvwF97wB0o8dMtm4HpjguNdcN4ITx
RiAD3Bl6V4mQADb+9QU//yxL4IvBAO6pSyeTWk8zCtUi0hubPwVkIp066tU7xz8hv7ofiifbM/Xy
QWxjAgIrInT0MhrGUyJWErkPXBGrMHHNpRykdYbOGCy5Y2A+jUR/42CULS6uU8nRSzA0kD9D83tW
otKeTV+/P+FInMTZZtQ9fYLjcEUce/p2yeddrzuX6L00KBJf0oLAOu5EEwGlvU4t6o8B5pw+bG/1
pm+R5DuNp9iAhxzljW0CUTQQrvItK2hr57rvWvxENWgleXdWad20sDUDdX66ODOUid10g/KEwVXL
yWvM5c+pXSMFIlIlAZcF00w5czsCf3K8Uf4p1GRu9HXiWQvPdCAFpyc210bDwaCuxivw/DhU9HmQ
PJtCELVQHZVWdRNaD0p4rpgjWmfTQ7GrgiSDUwYKqzqWI6gtTl73t7F3147oUo72ajDPKK2Pqrlv
SYGzUjs+03rfLOu0f6i82rhHyPHYEtyIrdE72pvshN8z2SRwz0AhRMdQGrBx+vZdm8i8hMVnClch
t6NliBx6aVncCAYxnbVVIKEOHhvfLBqruexngwtHuPdyuAl/GJauEf4HeBed0cs9k7e0XXacNqZc
4uPyti7PuThtxjJVig6bxIzUPLdzhuSDaVMg9UJ/XUWn3wtB3RXtyOvB8IqbIEFNo7TqugI1LEIj
YcZ29AS26sW+KFw1QcDxs02pnTx56xBrLRlK+APoHGOLToDfmvDj2eOuyE/0jS8mFo/UB0KNvR6/
dvIdbnvuMnVYFWyj49fx3jYnV8kQ+Oee5IAqdGtv3YZ8eI794gkocbOgo6z5PiSwXUbf3OqTRTRe
sb2C4zQEm4e4/pM0CLS4/21RVfJbUjWY7ypsNVzoRigv1IAC1/0b6FTmbBUNjJ0YP8+0arV3oQnp
bqs5nfs7deVbVU3k/4PzxmUo6VYdlpUblXAdhTQoNUKj4dFpv3gYCT4o1CJjA0rifcQtlula2m6C
kaxQKSgeXY2CNomeSugJC1NSctMVCg54WprroX79eAbfrJ7QxEx+692hhlDME8xZoz09mXUpOHJf
ctlK8IRskHr7wstE4ulV4fgQENogcoKkbLLr74V5qrGg7fII2JPF3OsgBBDAJKEn2gYIYF4jxgsb
TVlK/kjLG0PEcdJSHywE3yxpKKPlv0CZIpeUIiP+VErGNjOcd0169zpPlUvIHoxaE3+8AUbp9WPL
9Ik5QQIGTlCEQ4a+N5/tOVhC221ksgEUKEODar8cgy/f3UIL78kRi2jq5P6LkBIxFVpwPuSlqXwK
SIm9U/cc4G01JLBtWJbDSEKX2ewP8pzPMlAwTsxqBZ0b4jCJtSABUFLv1oPplT5zJM7dQwcPraa6
XU6JagLdz8BUNSr4si+csa/7iTB5DUhXU+otQEv8Yb4NZrXWpyhkcXcKhmxD2aF0d12atQ1rovmq
6GDH1nn82lr0w0IBQIkpr26A8ZcBLJNMQFFj/LBXzIng/u4xxRLibiEsOz2bkqD/YJLwFkSPhm0g
avloiNVP3vmYpcXvUbIV8YfnWfpUmYuuoDPvgt2pQxacPI0Xqz7oMN5SCVyhiiCnRbU2T6EpV2er
Ri/9/UMMOQRxPRoehHjhp01e6XdzyABQ3XGbvKDAHSXG2nYLgPRgYaGBYw6P8EUHAVlasmxurgxU
J1Y74RUkQomSLaPKzCp/DfoL2RNBsC40dpZMpEOcMdJfNDjLMSgZHm2dmrUZRiJPCOVOX3PkE2uq
fJOxt+OCqTMQTH/HWYVuvzDAU5snwGMjEI49bPmmibakOzDgZ4fJLU40+QzGLvLUZ505RLSv6bgJ
CayrNzL0u6GDCeu4+sgENEVwMtcKgB2++nksVSXpPK9oJ366IfQcWmvYBVtTz2TZFtKpaqwpekYk
g5qwstbX4P2L8emap+xBQ1ZXvRFK1Me6EmZKaN8vY9yiwa5n1eT4n5VjVDdx/67YAP7qUh1hGGOS
P7cY+lygkJRWuDYtsTKlGLoyjodUZuCS58GSMNQLsLSRJIA7k6V+1SYZHvomthQ+Q+arNohOB80T
7TCAkfXhDz63jIyH7PrZxZF+4/eVzYieIJ5PspONfs4UkgBrbBlOO4mwVSH7PaLOl9Q3WByuGg+1
G/2mNlw09KioVcDIMzgOn29slw6eECt48+trJM1Ueygbmjs3YrRoiqhLHQTEcpf3ZTQV02MtGT9N
kpCzUgBM9e3Fk+Fh1l6ns9mPRHD1ETibClpvFVvi+QUK30x0ON11/m1zYJZCYATk/6Qzn8efkMAh
J5H/D0L7rkievMr/02Ea2QPIQZAqUOvhwjD5HbnDPoZUaVwUuOpuSlAUi5zDlWCZrr08zgDsyrjR
aX9Jxn05tU/B5Q/gd2X1foEdDTHzRGloGX8lSAQqLxTWA8PtB69+LbYCvc2eAc+q3QJHGr92CZpu
EFP9LAEZtbHU8GZknHHakiKZXYszMbTNZ8vwlId+1d5fLegJ1CRKU+gWHJxUFQfxr2nNZMdzyrpI
cqLC307ajAfeWiVeSxR+4Qs81kaWT9r1b1Z0heddSsfV8hz6C2GFM/hXXsBEBx5bVLvlC7Nccxcx
QG2ihabACgSqvtmh2s7CCoXYY4IBkq+EAhl91NJ/Z5jxyOE7GBkFMmSqWsxW/LvRgcjy3rXXnfov
GapPNKAIaNmh3PUmsL1CncEiKi8fGQCc/XmqdnVl0xnzvXh0GrZeWsznIIQD2QUrZK1h+5LFh03E
kiPTKOoLNbyhsJsAnevbZgUD3NO+uNInJAQsheH32Y6smmL3QsC0cH6grOa0BWG6q4Bbnm/SyTSv
65/sIF91PuDnk6p42uYy4kS/rtigi2xmosmQHm4S30ucQDSLHM2NjQlHcyWtgeltwNV1G0Gk6W4V
dOUH8uY8yMOxnT36mRNH7eGpg48hYF78bhQYlj1u7lQ1JijnMl/h3JAyImzBlOlkYr00fOi/sSZR
xvKpDSBynYZsgtWraFf6Ie4wZFIK68sZanpS8gqFHI9LJrNKdgzsL8jCZP1DsQhnCkqBDZ8VieUF
mhY59eKDIVzgNHVqP59P6aD2BmjPZlJWZTBmwQBrB7BDEp0VF65n9H/Uq4C58GKeXdn2+Sz+tVor
PJUNdWDUNan2v5kP7f20lGxgjnHq7RdRjRxfJjtXXjbELQb5p7xjkPbpSATY6LZng7Wa6MDXghjG
TAOpmNHWMlDIQ6VomQX7RN9FjOU+QvkswDukU0nbpDeE+s8wpa2ROaJ00L/CsetI6zct4kYE17UW
5AJBzjmHZYMRhUtXT7XJ/ZiRnCxY4/6HxxgReX/beczFRbT3NJivKd0ArG68kWfmhR4XVWiyMaMo
IKqZ1bAB/FPx+7Bb8++jL4btjt/77uHQywAddsKZBj48md2Gta9ex8MDnhxyBOtnbaOUlWkLLOX+
/OkrrJT20JBHRV79sJQXcYXR7ccXOUwz4JxoE61kwX1rkvkdB0heCXyg1kZQ6fx/+2yt9v+50/pq
ObFXwzaUFh5bKTiML0jOIk64YSvQZexdl5AWItACCH/+c6PHo6QYFD+4M+UL1Ns5vG5F4T+pnOq7
IwaN1AgfSeRWYKrLTPWq7t4DHTanVz5X0Q54OyiaY/amqLmOKug9xtzFSY2TU3WBoNWL3bqseA4U
VdI9oJ7yHVK5jf8hQS3z1YvbAvN0CV2flTLASCZ6rMujmdtYwKFEGV5xBGJOxwPkKCeOResY0Qy6
ddYPFkP307ql1So3P5HRmqwfC6WsUbfWt6CRGKMArl2yvUW4MNxdglrbgbVVyk6WG0mVLm9ciXKF
nmIjdaS14HCMDQVkmHQwzS7+IfkKOHfXggh6C7t90uqahwU5QffjY9JqqeQfgAXn2auJX+4xX9d9
5N5otUjwuz9ptMKF6nkILWa+zapYrrQkuLR5LZ5/gPXWecBa1bkrgdtQmB/oTrDj9A0OZkzlFW9L
nDaweoGRRIhTwhgnBCns4qb1yIubwUipfSZDPn2Qvr14T8qO84H8CBcgYm7s6mwApyJxnQfHznu7
Yp9+cYPOU4HFurpPm+vOagAVv/vuym6EfV/NkH7RHy9qgAgrXHtG/Wpc2wSsGPkPwySbOnPifT2Y
v8pGlD5/tD4nbA21AVXGBnRHx1/1HudaYi6ozt9OyXKVqeRiBeUTlWKpA2cvDwlm3F1vTpbQK4CI
7pCmXcmJbGf1ULKc2/flNyinLn1jhaih/jGTBbvKncw/MFXaiElONQMWUEWOqLZRctY1GR0WvjeP
3slEBSPnPXTeCRvd6a99gFTfPxZHvAMyLKGsr2vYomMZmblvLi4MC8LoeiQdXTLjxPc6OcTw0OMB
gssngdLk6aaU1W4MyZU7xys9idXCd6KD1n0QIBNWd1NQgyThN4g5n8sc7JBof8hNCnfHlozXAU4m
yj4D31jb4XAsQny/20xuhPuQUWIHzT+FdKMTNJMtLFHlwsHiligppYqSC2heqDsMijnJY/gSfeqj
w8E/ejNlOt2oBk/4KaUNruo/pOd3KEVgOcuIWezHWnz9EkswZHaQ4EipCfKGh0XGa4abqMvXwez5
H+65EKpM3AiVltrNR+lAm2HZ74FHXYNDj0WlVesmrW3jg/lBKPynQnvFuS54YGHWNav1dUK9Pg5y
7YjLOMLLCa4DMGCzshyiy9BkxEX1vrbNyectVZi/P9W/dp57ghfe83KLXprxOO0VLlIOAq+CyNX0
Ad9pPedM0trh7xEjnrRtw5kSHI9HB1TCJmA+/kWyzRB/ja/WE7aTzqHu07R/khniPgUvsIvSdwuQ
j1WQF4t6m8nMMkoo5bJMuTICig1DoWMMwnzBq3EAedX9hL/VeMeYF24GYa5m9+oZAIDe1KYW6QnS
w+lOn5IBNH0W8fRCo4TIzET+cYioH0htNeiJcxfwTubNPLtdSMdblhUv4r35vyX8ppvu27ozvq8q
/14w0i8F2YdJaZmE52sOtiMZlM2q69BKS05H0Oiy5YAqcHMaGLguDm2gnRIMGUAEFVvEzpP6mrU0
o8X7adgH/8WKWPYc3MnNiX/2DUCOKVyHavJjMJVXOwP1+nEuPtlwpXYbVn+jghIxYHgoLBKJqep4
36X1+DPG+EsqGyw4kXNnmSs4VOEXFh10NOBdxleYKzMYYBFt2akdspT8s9fhGFMKBfROhkXEW4Br
whGSIK/1usKMwrIBFumkxIEDLRMaKLOlFOvZ3TTzz/YJi3G5pUSEKqcXTcg/OmekZEh6OwzXW1U/
G9xPSzRgO9H1l5Fbvoiqda1/gvTrk4osLXsTUYpf+9vt3frooM8LC1JEo9v/OfDEo3S83Kq2Tssm
L/OkrAkgISBAjr7e6X/tJsmr3hojhRoRCYVExnPx9OHUx2Wt0nLg+kx+wC65w8cHRYW25QoJaHaU
pAp8egnrpxdDD72q7HEesr9hvV3Nnkv8TwYojpQwaTr9QfZktRhztqkjNmkDJoiYulGKZN+Y1XEc
WUq+EbdjyYkF7ctyd+SJ9CVsyDOQsrc7Vu6NU4UyJ7B2ADkSaxbhrlyblUCcIYErUpYLwHc8UxTL
/pni/0WtlC8jxz+3iYvqlf/pTtSwZMqvfZyJPChVdngKsZOVeOnMI1ng064sR83pRjedIGLk69Te
8RulvUyHyTa5CYUKSlFNMBfpMcKvhi8beqMQymITz3Obe4NU7W5987egQTomuzncS70mdkbI/Loy
cw3fEY3uawWAdRdyAx2A0R6SnXTpr0/W4y6lPdyOZ894wnQxSct2Oe/iEBWoFMjib46o+ACLRd/s
GHqyK8F6KSUQ/OGoUbZhlesenquMM+2zHKLVBGS+j7/e+165epEWWfnVGmyvAyoFuWJsxXKRSqSL
6wMgl2TJx9t/8nyN1HPZiK6o0t0xnTHk+ne+Wm7k138lJr7xr8REUpVgX7R49L1Hy+ECqmvx7qdN
LfPbphv5UyAeJ++0psNXnx+jysPpecVfDQiUFjlwpDia9IonWr3VCO4NqVDIRpa/ihWA1qPR/qQi
JivwaEHTdeu4q8aoOasiqb3ce8tN2k8mmoBE+M7fLFmm6j/98r25K9DxbzEijjOhLN6EaI2m8ujs
51DClM53TFaQNRNRZux2dI7ATkRbxaMKVGPwoK14+hvlN346l9trrOuVH2erVr8OQ04aKkIqz7ih
UT39WFvKNqvObw4uUHVC4obHHZerIe1ZjxMiu0c86cqH/MuPdjOiBaqw6LJFBYHWINaLFyGItbdh
o5mcfmskV8JB2qkXXsKUDeXHiBRwf1zbaS2tGh+643oXezq6opiS1Vwk9pakNsqfrG4s5X1c17tW
c6h7xdVuia2w+I8rhpYCUSxQTz3rKvpU3XIKA/7uCOklRm7OsdCHAjcv2+OzETWZHnOyEFvFbjuk
9loyFFSraQqmR4a1zxUifCNq+ASezTsPZJLfmdfCrV8yw5by7ozkrpF+uA4p5jbh19TydfbL61VY
cQM3bgK5IdCmdX83CpUGYUMts64y/yFpIMSiVFacwzTWRxA4aJ+/W38zvFvCUoHNinc0N4DFynd+
ezcr01WsaYJkEkQH1toVuaia+q3VmABa26nj0meA1tpNj3Pi/nMDHecGOiiJxiJ+Xs2alcXW+Wef
y8yLMlDtLPgJwz66onGPPXXVJxFegMSYLrWIFVcYetMvlxKjKLYLar4EDwHaDAc6M+x2lUOcevYq
immXqmOtGd2QeJnPvXNvUvkeOjHQOzB6OtdmMpEINUWnEPlBT9kgCkKKVLTZK2BR7NowtMePJ53H
9gKuWINXv48A/hwsmuohhN0/1twjrAnrsqB8dt3Fl4kuAW/JbTZJy5p7fKptHe+nqSfoJqDmzmZu
xuasQkSNe7YRE5TjpsZbIeQ7jnYp9+kXLjPTjjt0o11NPtSYkxMC2wxbtcr/Ap3lBUeb33jLK4dT
qw1qLT5L5/Lx6i2iTmwvNnsfqarLFuyHDxkyHLPxVuW1dZfZUMcig+aIrvjxRER567keqhOrTURk
/PuIPPyad/YMF+VrPe9jtY+f7p5N+pYFY3eAw8MDx/OAC09MBHOJtH+bMGPpZMgc6H9tzObJp1Za
hTLoROTu8MCbAUG8AWOqd1WyvwA9qhmibr7m8JURdNI0+jdE1yYnwDBZ/ImqmgplaXTh+HX0R9jD
s3QpDUtvSHnOUUCVKhZ2Dr2OVjMjPCfFRxTTY03wnlkjmo0OL6WHBuRevNBBGrxPj//3Zix+Sdu/
Zs8e8sJI9DZ0hDy9t4zGpPIdjzSU6Kf8sEqGtLkkmBeRvF/ka0BZB7YIamlv/VwDHHD5zr+/e87S
jgbh0HN2QpUzmK8tIAac2v+iQhMhTAod/pCIlxggKQ74f4Y8mjgCQwoT2o5fOR3Crr4rcuC5qvCa
jspgNz22cVHoH5n+pSv3IHW/Ib8+9rQbUmZjLlCOd0zPGhKNBnDJkrhQGvnKtS0BebiETlcG/1IY
ECfE5mOn6Do0ClksPkgvFv8YoQVln6HoZcEjwJbqzR3kyDy0mrJlMwo/YvStW8UnGw842RbpQYHg
eyJr0AYnKpdw1rAEoNIgodwL2BF1GlcqgJNtuxg/+k6wR22Z/au4HCgn7Rd70R2FcGPfl9T3dVDn
K660o2dMkG1SU1APRQEe1a9eltZIjZLzVbOeT4Fi3oglWhOxHf0tkWE1inIgMJT0bICcXwUoas97
Lu3UYEgGAF7gv2ikvMDL5XYjOH2mTnWx1kedueUvGSdDqaNwZR48YgTbWMNctkt6UyNfbAbMxcce
yepYLjHYJr3bAcZVgZKRNhZtHLb0jXo7rMMzzM1Fl4QqSfYn5WpYIetHX17q0Y/FrTCOIjQ2N6KI
NHVIc6I9P4doTxfLMgV7k0e+7bZbavFGhtSp4SsExeilLO4pWXrgXKJ4UizrOHq7iAK6WwF4Vkvh
g61TPn+n6+FSo4giir4QN1B990QU3mCh0vJvCUWFhwAm7+O8vnSEgfUpXx7mMME3ogsrkDpljIWI
aY6dE1FqEiNEXKNIRcEkRHjyTS3dQ3fWHl74C46sMDhw1PeD0OnT9YkA/qQTN+f62P8MrN7HaHoA
+gGRBw+HeW92sIfgJFr86glL5mFGiyFDqjkWpkqKCo9gWlH2JcCc5Ug+3ACZrgMgCo4VtYUhbodc
d/qebWbS48XviyYbL4q3ZCinWd4sVPXEgWMWCgFuy8r0tNoULt4XCQNjPHFMe5aMSpeXOWOTiJ+3
SYwxN5+mu0IQtJO+SFnEPUH1iVX7dt0X/NJrobPpjiDGgQ4We5HQOuKb1FPDhlgCGOJphTlBemPc
XTnP3U5GYK/qcc7n2n/9rbZfKken8Dt1yA0/JQbajhDnQK1I4p+LzFY08y8Z1zzrSVesggFkEMh7
ckh4NjLOqSC8zTAXMsX3S5CJ0gviHc/ZOLVaBnoX1vHj1kDeLz4GwfWBunG7LCeLO5f0bQMPvXzB
2M9XNvAuJyVA/AXEibNRYctg+dvZkDQwGfunnvsLessoweyCxhzDZmFjXDfGbbfhnRH7DNBBdo6w
DXfJ988tJQjp+xhERHk5IQNdqintGM/tf0gcOuqgmS6cbRBBsbmUQiXO0XlL5zwsBo9OBPB2I5W6
K218gxgrImJWXiGIL6K6g2Bt6wI20pjehQmNdXA4zhWqkgBr6G9b8CUAGhsUYLk9BZg4fyEMCetE
Vq3nDyNWOPQSy6ZZHqhJGRf4E8CJiUHEUQmF30DOIw047xTCMmae5hyMEvwfnIhZR2IgCy1swarR
1mKAdpCPrJJofPKtWUZCzwfY14mKNMrCiyVnv38E7jXDZlyAggTQgXU1xXIWqcDkctyVlbl+97Rf
Pgkt/3EamSLhqVqkvpgMYzbhpmmknSjgcLO4z7VtUnrnvaF1p6Vn5wVkT36lMQdyOWyk4cTmyAJX
tH58+FhjzyLBL5av9D0vdUybghSzOu2RouxX0fMzJ1CequSYMLWBXK6wQtW90bTTGwoucS8CNYrJ
P/pdpBY6QrfptwWJzMhIjGUI47IbGofwcgsXzDaLpqqNj931zl3DMd154R3BXVXyVLvCiteYMfX8
OM+Tx7W83o2nrmuhzCWvqswO4KEtyvldywZhgoPkWW9eS3l5kOLxKsmymAngljj5upZznB1KpKxC
+sb6SV8nBENe82iBX2l5gqLACtMcWhjb4EWeGRIodb9UlxtdbQxD7UkO/pxSlva0ajeQUs/cy+bS
HXodUsvAcmkGpjvu2okH1FxFcrYO3d/EZzXDrBqcnZh7la9J75AipmHEROwYHR8wl9Up6OIS8FxF
/ZQsarhMVKCFkSz7Lhdj7dbtIlVAO5pMaHTG60Ypcg8hbet2Ans8z9Rui/jLPOTP5JmiXhMPwgJK
hy0Ia8kbGIfs8+BTP7SuNuevYD9WrlFWSJfeaVG3NDANRPpiFlAyqnMeX2X/eRuITCw477j5Oo97
mNK6g6U5bWAtIbLGrZGvoDedNMP/AWnzTOQ8KoxYopuszqav2lKvRDsVeGPr5NH0qL7BIKPsAvnN
UU+jXF4r6oV9yRP6XWGJ+lHDmRPxt2VEdNWfTyrR9DjAO2ZcPteFgbcTWlyh4FqN1RtNJpLWagSq
6ny1VMfyHP90PxP8e8jZ2xwaAyphtwdR5FKhbTAyMdt/6cDINZrGCUy+OrlxB8H8ZYn+iz8DeEhk
bD0cJb1N/twotiL5NLuLvvTiyEbZVt87LDFOzmX3faN4wf5hFlS7c66WukOPz07LdlLkwQY5cAc2
E3ojJmQSn1+VHISaS+JJWeSNmaUopG5Q+H0cC7UypypKhBw5IhMXw+puys58bPHMi9T0DeJKv/YW
BBtJyeI52xdxop/Y4zdL2AucY6k95F8RQ8+oLOfTiNYkSwhi1jpl986ckbOb3aETvOHwKM3n06s7
yN7/wOwuLOlHhJ2CoDZ8cpiG8YlSomYSKvD+P46uH4mT50nhUhdhjeS4lJkKuoDiw6Y9nINiZU2O
S0w2dl/Nuav0YRIuFjFthJfZTZCnEnHrW+qDvBOMcTWblQ3HWWRVX/t7+tD9MM5uNZ/h0bKT0D/s
EF7Ukio7lFFh8cZdYJ8MX24C2IRnt+SdQLb0J3/ETAT3LcLL/v+i4EDJqEEB2GHRbBG4Jl7+3h5g
4knGz5xClAat6cHi8XXQ1V2h2UeVpD1J48Rf9IIVGD65QhYIwfnIqsJfZHlAmFZ9bHiRuzSk6Tfc
0CINItaNh1T/KCfimNp164g+0M6Qo8TYT5+wHzys9fvnSeunN2Uu8yIXfA2s5dFRsr9GpYF1O0UN
HzSKyN16l5yrmvk10wMg+4BPIAEUhM5+Pl6V91760iYA9gtLI6eiRYaM0dh+Zo+PbjwERwmhOdSC
fNQrh6x/jOyOjJJDU8dP5nUTrgQJORPG5gRkfKQsza6iLZQV/pDALDupB7JfxmForyXsPgC6/3Wv
cjk2WPcq7fS7Fv7VkdVeRG4uaH4irTq1LJ8o6U/cfXf2PFdIQaJE6l6Qc5Yb7FgWBYuEeN651+T+
/fkvCPuW876mvRN8OIc4syuiJZspuGC8x1+S7d3Tu7kdmHZHv9gEnuwVNkawI3wu1eMdAS1Juz2V
A98ueE83j7evovKetm+9Sz1D75APn/5YkTP8UEvWvkpIG9y/3ZEDQTUxvIryntFOPk+E1cWHCNF9
0IbLXZ5n4yTr6utK+BVLXStrS6cBKkblbLeWVw+muqNRed9mRKljoSGEjvMccLRhZplu+Tm5QxOA
ZJbapZN04X3XG+csysJepcHZG/CgRm84vbWyd0zV368Sa65E9RDoPc9d4am3T1EFbr0gpBvGwk60
w5ZpGEc8gtrVdOpUgQgTlxDu4ahTpodIOclVTdsIwBvod2RWTLwtGnRmDCTrCiVLXaswg+YuMxi1
AVuTEJkD3m1bbbENyyWiSBIVDE9eFQhWQqqS5tzHa4wo8UI1d4R/SJEmZsTTmYdY0ST0QsP5B843
kfdvy3Pg142yMvT1eUW4uPg+Tb3ClGgMvUpcykPnOWThhyg9HuCaDKlUibmGQaTWMaHbeAfHYkRE
h+gfD8rG76uVpGNqsiL2ihbej2I45FdBqmONSuBbQPhkhGh99h7b4HQSy7DJWB89y2tiNCLEiWzV
/i4dnbpI0pnG3m6UxTPbX277WdJ2ULEVdxuW3zfjrFI5GOEouv7Cjx3rbL2g6+adzd64uoJwKkZD
FJ8KfhFCnCU3JfbAqttZvGWqVvkq2PZAruswDm3g8lP8/ArqNVktYs44EUSx4e+aj2wYyljd+CHz
NdgLirin2J5ltJvg0SJf0TQzNElM2yFwkjC5pW4o9FcTk56xWn5u9kCWcIzxvyrirE4YDeCRHFfK
rAV0GtKhcFiN2HUaZeX0IJawuTfwTX+NzT18VPpMhLzxysRFRlRVroDPSIFtwGdcB8+MFiuCVCet
uFaYRr5Z9P3ihlVvSgCwuv1p6Ws5a0VTOj69cj6YwCQ5yEEgRxfQRWvY1wzYCwnBNHQMzXyL7HKf
BbecvUTsw0vQBWNwPosIe+HeuE4jdy+6G+bVVfF0/UHO03BZkygbHARpIRiq01N1dZmY/Mndbt+X
q3O8tt/yQuPE/NNT0BVNUacrNwxIU9FXXSEhRaWYAc3p5Yl1LlTo13lhgsEtxvXcGyk3a076hOES
c8Ki0DY4db/J6idqbN+zI7TlioKL96ZoYALG6N8yiht2lvZ/DpTGFAjS90tg65gZCtgBzMr+4sK2
DHJ/kUBC1w01R6FUAxlCwZt42Co9DUZHFFVqK9mfaNpvS/b7Gg9KExp+Oji6SM3OvEzzXE5iI56N
j0RgcuJlPv8H3G/LnlzXFboXdLVChhY3yqaRMpWYr2X0yJspk+GPKrJWfrBxDnPqagUwceC87S8I
wuNGz/glupy/ZhyAC64PMhtft2/x/GB2n9haV6H6UzFdQECFgWMXZEofgwLOOzyku0Q8BOq/GMaK
sw8mTvMTzipHtSgyjgR8c+pjU9c/A7CuVYMmlvj+WKJT3CnxxT5lDZ5B1w6rtUh3YizPOmbLmSY5
lSGR+FNA3XTMAuxJGKH7IpQCEs5s1IwbRxbNpq47TRpxnt5Hp4jBOIRfWTAZwNEIHWL1b80BHdRB
LmTOZMOXMj1SBZTDJVPDYxC/p42fqtSdLnd/RCqXXOj22ZG3HX5ZI4++IQ+bVZy08W/1pKYFE8/U
wWrq9LwF40BOJYF+/WQj/DusFua6y8lovqdXkZZjS1S4ci9q5ZMgzZZVvtWvvkh+1EWscXMap7QL
/s8jtcNHYMfBVgaSCc+pP1RamUludzS4rvwBQppMU+i/QC81hjTo/C47D7ytSF8ktdmNoOIgc2Tk
X6fl5HIsQIXOMjwHuWAi3vqjY+FM/hAhrS3bL3RPeWHS7KxTsynwONd2JjYAz1TGXlAsObmaZ+or
optPxsh5C5nmoPxZ2dgK7CKVVtIKN6JBa9VAQrNyE9kbcDtDxKZpiBnC0q2P7cHwGO3oOoOQCUxa
odHAmvWSshB4fGjldp3V0Kku8pKxeSVkHlJaxXSTWeVt3GRdR8pVndL0RafjyIr60QWCthYOldjc
PtOxrvYYWMucN5hzUtXmDK2gRKpUyCx+1cd42bM1PEhmffrEZRA2RIv/0/DiO4NhALul2aTjkUq5
XHcUn84mDzMbLtGMHtSorTlE6cWrm6J3838cgOKgEOageXDh/ytiuq75h+GhSf5mLAfbowmtynwk
Cj+dlX+lj49vKaU9dZJ0tDHn93+TL3P9P/PoRJvY4KcJv44uZzE76P2GP5pswasqHeg208kVOCmG
rATd0ZIetpHZPjS07IcZWBciQzcI2cJmoTDXKzEZfrgNdL68M5EaEH/8oFm4W8jTGG6mjSL8AJ2Y
ZtGusQgfi2J0OL8sPJiQaThcnQR/pTU6GzSi72mH6p+wGiu7NLxnrYIZcMq7SVyA3cBq99wZ0wmp
V4XWl5CpYufYu7zqec4W0ciI7fuutYu5uIpmY23J/QrZM75EHRXQNO40VQz2LqFVNspGdxGcrzgV
yzcW3TM6qFEW7clivp+2UZf+4rgtbMvj/NG2bmDbqoTupOPc0aj51uDQZZHOyj+apWShzlkRYfey
vXxVv7kYzwNiolph0lPwD2XARZxJlaZzlcJA/wsbEYcklw0P4fTd8leM2XypcnyI1R6JXRxq2bZD
SRk0MigfhLRxO94OJwsmZIcQDqf2mKv0AfD+xSPmoV69knjIjp7TqAfwesPKK3/cjFpWRPCTc8Dz
hGH4qFKVF/BzIi/aZFdH0oc6TLinEFbC6qzo+rElghN1L3lFBcFc0GaMkJSfL8YwTcpUJE3H7oFU
zcM/p4JWGZCcgDzecknn9zTOGEIhUz/baW2FAi4ALnT/AyV2SR+dptvh7a8fUHDlwed+Ia0FlBGI
R4/YqeAa701JsS1avfD7DUdLMChJTfiaWNvbtpYG8n87tH+O5OXhnepGO81SRxc0itC7tHQZXZhi
7Ua8yQtF7d5ZOsLnf4CHWGoJjl0/nQxCJwZ2wK3e6pUgowFt/Hb0Ig2ZepRQA9MUaAwj0N2Q0duj
ssXc9aAwHqZWaox50cQp74TfVe1uDhjCFwXjdPrRqpue6p7xTzpKbJUpv4mxiW5NlglMv5qOoFbI
8MP75zkBrUDOVidkoWWXDHgN4A+sJTHdzcUK3x/iJ2BsfA3pUTnVEYtjqMb0bYP1tXbIErDMdRDq
8jLy9u8lmh0eo9s87jdvY1hfS6EP5rMjbi+2FR05WahWIEhsrkRppvnzZynqudo21HIWC1gD3oG8
parintb7RnEf4pBWDF6dCjTp0sf9YCEOvjg7SEUQsPZoDR5QywGd6ky+x3f97ouJQeFCEvh/LZLZ
U79qXLGcZPJ5A2e+1h+rYblAqwfY4ViAFEVSlmTHonx7lG1qnLof2+Jk6qhcLCS7v5XQndAVHXoD
9Vf7Y2My5MspKMijiLwRv3RwTL5JTulrk475SSWKKGGnF1HJh06XXTAr0wHZnWC7K2oSXN3imvlN
t/QOFu4C0q1DKM55o1kv/VUEPnlPXhQhYANwCTbFG3KEHaRNoQuEFdqoW71WTSbin97XzFuBRXcK
sJnJgs+tJgtsCaEqgZ2lubNRTf9HD1VG3cEOkGbhBZCYnfbQX3/XzcRvaLK8VCgqKqTdhzDlRAcA
TygVUHrJMqJGm4Xzsrgw3lyetrZu6oZjoCtvcWMK56Lw9c8juayLxREDSWQ8gdRgcJHXJz3mNX6j
+eZZnGFdzfkyYGPs3rWNjoGA7/S5YZjhINzST+heWuph5bPZpB5omo4zUy0Tk7C/oDfs71q1o9ID
rRguEvYt5Dae/NUy6zCxyrUdEx5F6G6qlxlU1LYbAZuw6tRBMo1o+FV8Yg22+eF893wjgpzn+R49
Ll7QfKiNUKnCAjbfxLsZq48a5kXbfWS7BZuxnLJRQSPF4x8cJspncLzmePx6EFLLRs/fASeNSyl5
nauPbF2jNbQLc/u7SKINwN9xtbrvU1b8qykgcyjdf3lTTxyoyDDkywyPxZM8LOVjIVtpfuo/nW4V
bNDDAps6+Y4jYxjbkhLPVqWnsc34Iwqfdub225qJHVWbnYheIBUqCLsOHTUlkPik7NVzgY7kdWOA
Nt0qwJKCG1wBiQeXHAClDBz31ULPFYxkfQOghXP6KoH89B7uY1w8bdSyIVCBSLbFfb6yfABhyONU
NfM5uEna9EtmGBdXTALZbPT1pFpbrFl/aTU5hd/Xu4Z4O9H+/9DccQVo740eUoiScSdJtItpqdho
fGL2mouV6mniDUN/B0LzmI0P4j76IUNnuHEwd5kBRHH4VILcv3G+rU2fmbtZjG7Gk5FsXlsGvQgq
cU0uq7qnDSJimWrJhCk6cpefqYqDgmqQO51/nWqbC7x+FZomEDoGjCSvYf+wMvsa4F8Doj+wMkjR
z/ktCsIFXJkW6e3ph2SWocuoAbAY02yg/xYH0p8XKdCuoiS1PkHUOvzE8S+KwsbQ/CQhDc2lhO8/
WC8Snqe4PYm9A2iC69YrexqV9l+IeCDSipwsISSFdZI991Nl21KUxEIvx0Xzq7pTf9P0j0PS9p7b
QDBqg2XQVA5FN03w8q7Z64KKAjTFfyAfcsEvZO8htLnVe+WB9dq6CauNSqMZgKEiBJMPIESokaUn
u1+qV0lNc2oQpuNRlRNDeaB55l5YmuPl0VyItEuu8GJkOvE0gEpzxn/Bki5opyjoGVnGbkSobp1V
wzUqSPa6wWxLJAKw0yaw+WzOZn5lTpBHj1MOEShPAiC2XWfOSrJHlQvWM3qQTWyRJZxkZAUEBRCU
+A9K1GdPA2kzEqg+BF/AyCDK91fE3EwayyvQFlbKZw1K4iGD+f9WZ0Pv3NR1ghBonVCuCwBUTFi6
Ly8cQax2i/Qtbu5uJ6/V15CVGkR1Wp8SwbF29uICJO+hsx1F8mc1oEqdp9etsDi2yrC0+J8EP3zh
4OolQHXETlYMQYJ9FMRWnsklw4cu+wRKYH5MXVIaVLfvvT9jRjyxu3wxuZkfPr2m7iMgaDcjPhe5
Q79ojQiyJ/qMT+j7OK+B+rPNFQZ36j50L5X7E7njRlJLuMcRs310soFrsqy8l9nq6AkVmhXuL946
q7xrOvvMaaAsaGT34ZaeiVRnDOnIV5qJudKcUZQvmEUygs3Eu/FuwYKWvWT2UzGzrGbsHpIxjgJW
TY5QYxiCyWSegpL10t3VK5NOIufIn3NbYYZvOZwUU+0QP+qQnK5/jmjUBcq3rhhN/I3aqaKVO+HH
e1v4t3j2JA8NMCtuZ3pNsBICzyrOn/n6uvFmRH5j4r5S215oLdngFW/fE+Ot32+PMP0En3+rOu+L
9ZLowgT3GesPd2MmxzI5b7giUpUgZfOltIbNZOuWY5ntCJBxkjjJv3rYl5H7yt6psOpmv3IwBc4W
molTov3m1KVyu3z+UQnlsSiefmvPR5yd3BZXS6DlbrGGPbWbr7BgHxNgV/nyr5WJmG48t9puOQPx
VJXwtSxCO2rWvB4e0s86XI9Q8Zn3uQupCKAn17V2psv4u9miRmToVGOHj1uyMqyvS08LZL7XNxec
yFVf34UtJhjxrjXB/gRC+r9YmohDjXf+c7FCmsxcwgDAeglvuvwe79VGjLgl6G9SWLSGIuzfEk3g
O6G9/GadMaxbhf+lYl9SfwIWJ4hmkxcKpjJE59PphqXZBq9tPDo3MSr0qvpIbSYNYmu8GFRx2qG2
4FWPoOMBeEKGKSn7kc/LHQGLV6WnLB1Sy3/txiNF7weba5FgfMvA6uQLEB38QxquirhLBy96AQts
6w0Whs3LQzUmAyd48jrgdALgbzH9TwwPg5/w0fTniWTEkoXemzj5+D7aLUw39Wsmk0wUdZbi8c+v
qCxe+M9JK7hNf2TUPpHzVPwMkb2RtPT/0Dk6gA1OhWAUTgq+myOEebJod4EIHjWkCCjveAnh7e7e
ArvP8PKSx1RFaeh2mBZ8C7LO+cC/cdVvff9SzqYJ2DSeL82IS9ktlOPGy56fXlMZx5KWH94DHpxp
wmDOSxS48MaVIXctKMck5dVK7uZSYjsc4gPQiZx1j5ymltXzPvMPPttVSa9FRduKwMLvWr0uSzOP
9DIgwj0bBZXtOvWSU5k+CEqF+pHfoCgm5hkBQYUIK6Z7AuwFeeRYkJ20U4LZOYc3Ys7XN8d3PPHX
K/fHQOwPjfwefUWHzbHKqsykGx7kJ+5TgX1Zzq2AYDKxtpzTD5GUG99fkPaCbA+kanlrJBE9tGVn
cehScG7sG6ufG8Iuv5KI5WJRjW/lhNNngQk7P9jfj2mArVXu2Ib5+97xLok5S3UrOrvYY+18QBR0
GwPNIB4lq0fTwkNyqvf6ENyLFCgesHO1SaA/9XJTGpAYP9b4m79Cn2sPoFg6qLjD/67W6rozi2ad
El1muXgL3+9LtUasg7oquaLkZ9Lsh7hrw6n57bJ4grRF193RPJdCA/4ZtJHBTwYGqL226Cbly+Cy
2srvLiUqrOhaZE3bTL8cPOPXjgIZWw3lGNY+MwI+cGPw3Od7+dJCzSlW+kKNIusRpTElwjXMsfgc
hv8Mms1LT/Hc2bhIX/05rtHOu1N9qNCMXiZrK36FQwAGad8gs0OunV0e/Qpx2/elK9VJObhw84TE
b0gTvz/7mzofOpmieXDkYofmzEI+bz+cpNBadBE1RhpLKp32LOll7rz82qv+A1b7bEu90cwAjSWQ
JWcxpRKTiinKzICsw0j3m1IpaTPp3kOpzin4xDUvnBEKmfXE5H0+MRU95+p2G1IqBbxqL4xi0r4J
E/OWRyMVG6oI457qL2eCpl9DpUyjbOEnL7Z3y0GyiDhvL/PrTzRqjKa5TISozzO6ng5NGBDnFKWa
40l2YNZKudlVV5YfoqmdgmukkzW+tCL9w/Ih8sg1uyont4GpdJIWXO/D1Fv40Nq0oIq7VitVxho3
3WrQaBv9BDKEGR08+Bj8PJTF0rsKgOUxTPBAVJfguUZ8ppVL7AmeHASHn+z526XngOPGN4ayKKN2
I8U+2nTbRKDrVLfWIFVAw8e97BE+oje0MpyCgOhGZDQZvZJhGC9ZbYsjibTkBz8doW8MHoUBo6t9
31vCMG/YNgFvQivbOoLW5BAQl4nj2JEtK3W7Py1ryZhCdKC7phYeS5GiCmxCVMpJCpEmglxIgqRp
nTD9rRlLgg2dm0UXfSQDDaHlJ8fAt/SQylJP6PLrWGuxg34R4A2hNVQoj/GCHf3WrGHkNw54v+Or
HfZf6x3BWhvLQaBh2jds5ax81UeEeHtSqHY5+IgRWoOYoQrjIRiQuwjlwP9vo+i75dL2uYO7dNsP
i3jWoEr7CKagLDU9shh/3ZrnUunzNFb8aVBqvDfKhIXDDNzDWMGecTAZ4bb7ujpEN4BTkylA668K
tc9w9AxrpsuHqIFjA8Y7jzyZjO0oB01c4FbqX8tvZZ5rTDXv6d+ZFeuonaTg9oISEXNcfUPSPkHf
jCMtSG2gjFzSf88aC/YSlLIGAghZw5lMb5jUsE6u8kmW+ndqABhNp82P9bEu9IyFJBQnVhccRpgc
/6+dsVkuZPIrmuT/57ngPXwApfMYez8iWOn0qhLISP6SZytUL51V6Gl0d4jeIsiehRuTdIdjadJc
CjaGy88719FXJohKU7C0qKL5JvGjnNuIx5elTOzD4oix5HOYRaVBkfGTXBYyudMF3lnnHwR4rxNq
4iHcRV2Udwpp/fxPAcBWDiY=
`pragma protect end_protected
