// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:39:19 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
asX4DohEHacKlNUkpuo0YM4bXJaVHMHjW0i85XQXT5hTGuhvPbog8iwidFeLzeun
Z4fUP3REimqVb9NSH1q+Exzy6edxJPB53kOBUxXzxShWq8NZ8u1D7F4pGydX5BT8
MogbTYHBI8uiPTge/LexWLtdzDrupjdcA5MsF8/sN80=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 42576)
oTX4ntjjt99lA6zPxA2G3gYVv60uG1ZEZPzfScLmKK6bWZXkYnIx3dkN4dA1yF+q
HWeUabbSqshgDtBztOJBpr+twF1zXZGMvkiIFDntCz1m9gjmt4bluxIRpkEVvhsP
XW3FzM8z3eSJBV1+CiMD2fwgz6JnRDb/cFpGFzhVTbvhq4w2yB7ewtGGcvpihf7X
hI83KTW6gxIZE9e/UqzLLPhgFy+YBpurCB9mG2+Wpuuhc3EuwqaNDib5eMe1wz4S
2KnGm1Li7AIbnRlb2mp1EnlXQA8WB3QNwtXH7Fo0h5zV/Qa0Vje1dHmptJwBItQQ
f3QiGHZzm7wsmgLw1Sw4GOXdfcgm1HUGgPJW3Q9lwHSf0Pfj0xCww6tzugf4wAcj
i7LWSdBYhTbTLapUUwd4C8IOa1NQob9meIvT3orDdBhlgywCkOryUBNTYBlIqETI
Unoi952jkyhYrPd+SnKEaNIpbWSIlCX27V9eSwCGJCLgosmE0eI++Sj9ObmpOCLr
lpEruJWXfQ2JcnH7xDyna2YUVOGAzTTJso/N4IxCrzrz7KOqfL0EpumROYscKOhC
XBBRDJtMQlvFSM1pYuIDCPn0JS3o27oa7tdJ3qGRfFbupcGfHy4D7ZDUuyoULARt
PGAKZ2bbn8wBPXg3tY5PPUpZfoWBaK9uU1VMsU3/gBLCQkDFVa2unlHM/t/yPkb8
VA7ZvFzD7DTlQPeI6BgO4MAkJKOLZXkJozi/C/cHoy+Xu0oZxk2rYuJHARvoSDS1
pNM3UyzpbFXs9cOMMNIaRIaCxU7mnIXIjtlpYcQAhPxZ1NVeOTsfFchop9cMMY5g
Fc3aawJSY7yiD9Jf1nheRLMLziKBafbvYkX9JeRWdwW5g5uJjuYWCw1ZSuKPfeWY
9sE9VnqWeFB3KeFBAchAJtCTd6csqKzjZrZL375RuEpnvW2A6z7LGTvw9y7+0iTf
wrE6LZVffTEqHT5aYdYoxg2WWVwrd87fOMCuOgzJGpntEEmDEIasZKDzzBa3PyVd
DH67Joalkb/Es8Y/z5e+QLYkHCSU1BhZvX1TNpOclEpGj5N4wGqeS7FNC7hBkuT7
/PhFMO8jBZHN33mpbvEmvjRdTXSREXXqdLpgb1h1YgxL7blLCLA58Rf/AM15GouX
RpJCEtmVc4LpM3QI+b8ZkZn7QkktBMty9bxGh0SlwJUGh1KIRtuqzrQTy+Q1xpbg
BZz/pBNpol0sR6sXOL0xqTaziYOx6xAdxuEuU0lX5Izv3nTD+9zdgvPZcdDw3NI3
awFBVlUuu5XY+PnV5XgrEl3YgCdep8ub0wc+dD2KqKXNc9AYkdTMOcwtsbCN22ig
SsbhI5uj1jtgRMDlj0KfovW3hwRZ00RMtgyC4yKiBldJFrqyvWZ1mWw8WNeWsTT/
kV3s3dMibqdr8TE/4IeZD7wtR0YksroDY83VOa7bj9tSG/3eLxJyskh2kfepGnEe
31IxVJAvapZQW7i2CuQRZUjjDcH7Tc5TTTzX8LgYC1soPWse7XPFHft8drHCnEcQ
ZVKSxjqFvW9NAZQUMrsCJLOMnuW67tNBn+9Gf3jhbNjzJtGvYbawEKbo/KJS1cFI
wP7Y5wYv84uYW1uh2DrQ1T3l2vwROKN8CqyGuFLarsUKnC4PO9DqN4Ls5rxC7+9i
MRmEvfV76EJc7eUwRp6lfJXnBuL1lFo2ROiMNabYjAy/NLvdXbFzcHwTT2XMi2we
ZUYTkDinjesSr2Zb9/o1yJN440TejzsyNF8pU+J0hEdp7Jvfo+LI+nOAqcM1Mmzc
svNsuMGFOO7CYvCJ1/llL6bDvzS8zUC/M7lojevYOXnL61jiRyJOj/uJ76SClhu9
bLofzbNa1yQgT5jhrP5V7Bg3fdvr5HYddW9b3twCwQzkComhTp7kY+bwMoEYbOZS
r4j1nwi/uJhOqWKXntlrqcM/zNNu0WlVbTF5EKyIoB3JojcAZkl/VxCurswQ7ljw
Q40vqKXGO4av/TM8jMxt6MHdrSV9i+VqhgRFvtXj/RHpsjfjv2QRZeefiqldBvsb
gBBALYhdvfU/SlAK/Rlgq+yisrI7QZR/S7zFC84L6H1FGzE+iSGEe7zN0CbvqBiP
15e2k5tdnDNoJrWFFWJjsZlLvFdcSZGsWZIRXGX+ZaWnY3IylvBPcE9soLc0Eulj
P2wX63mWj17V3ao550FAuhhPu7BCWZup+EQk+qPaSTzg8wBUGzyE5xzJDbo+233h
+GKyC40s331QPifQssEtnZtNC516DkYl/AERcigbRjiiEyzvpGOsGsqVISogT2ZF
MULBnRtbXByIFBlLsfsJV7vPc/aKfBGJYS7snX/HYGuEfb/mcZ1ae/BGScFS9ASg
Oggq+OCPXfctozdauzqCWw8duLYrGLyAyyCUOA960PRcH7t+eGko3CGJDj7cvnCN
FzDKQlnVltG+MjkV2ZTxpSfcQ4iKNBAUe+QALaZIMmblUzIT0jSUN1WRlylfIMKH
kXQYB9sDPlin6qoaHcdUXmXtwBnJ1DvVK1EWCL3iB2ycnNML3hgHGOr8IWfyHQ/A
gNaE+q7L7ZbIjr2sEd7qKCZDmnDb1Mc+rRH2Ol/ZT99fhfotzCkQdDO/mQaxGEtx
hVaCqT/MFZyDiVhRYeSFZ9Ys5OBOvtrfAutbzMFGUpeg/6m7Zb/LcPQM0uvvJcEL
CF0KeCUUvt1FeRJldcvcgfkry5kt+keCzRDgX0Ib0kAK1cSTcFIya/y3KpII8wAq
Cwkj1AIJ3pnSQtwfHzQUHb3KJifNfmRwxAVuSBvUwXfG+YJToRJ6/Kb06HPxKisV
IYfFOP7lSBxprJyo8JYN+e64OGO7zUeSh5Viuf+OhaMANGsHTs4BRKEKf0g8CcrJ
aGy69lId3NYwbz9+1tmC8hQwAjAZxXpV061RD/YbHIW1M2a79z9kUybCUEb1lByQ
qv8b8TT1TLvO7bAPVPM8vLRQIzaKNNYunR0TOvevyD9h+tk9E2j/mRyP0soEuGvk
4d9wb8gX2KECi29UwEt0ZRRvuIyzGa6wPTle4YAlAkXDbpjuqFwNslML4z5k8ipb
1ypPjC2vo8uySVV44UZb3VoPpo74XOKsB+y0+yJTxVNNwi2rFT8/0o1i2em6OkM2
zGp1rpBybOiyW6HvSCXfu5xlAqAc0jpZwMGwLdLEQN+R+q7MzPrtf28OCS99bzdT
aU2vFyoPfmcWYPXih8DGY/P1XzvXLRt83YpfqsuMN9LBH0beClZ9OSoUfzpDz3Q8
ms4T4Sxb4iM93jKFLE10XfLuk6JL4y4U82y3390TF684UZK4RVtq4cseIsgAX2oq
zXBMfnLFh+1bCF8UsHN6xE4sDO4FtGTsa+nRM+0R8fwAQwVWQH9qUvFEmqfBWIXY
ZfCsHxPA/q3Z8hVrv71g1quvY60bjyAfY4C5ap7NsrQjzSVBzuvXSKQ7bL+dFLae
VQB7/E+nDFrV9JtJt6GwXK5nevF4Bjlx/pQUOXMLS5WD0wq2jPxUj83hWilcZ2Ow
Z79qKXviz9wc0wHGtvNhrgQf8/ioHL+WdKtFnnuyVakBdSBg0PRz3qAsvlNKbzBm
YHR25jbIld5ybhgAZxjqm39JfAAzHujemoVEOqr18piOZzfBbb8Wbe1xZnZJPhxx
Kdmhby3C2HOUHAufNgW9Jg2BtjPKHZccyRYqK1Zfr+hpQ873LL9Bb7waSJ8CBrIh
jKKdOkVoJl1jJh0YoibDKsF/8/kdloa3gVqmiC1/1waEiAP4/0sf4grJcB95qu3D
9Ab3ydQIDUZrbaCtrEsQdOcQsG4IjjxyzDkW18Xx8E3pXUBkMjXgTiRRnxrzUAHY
fd0Fmnwnp29f4bbio+AYZ3083ZWITF6Tm2QYoOI+w+nV1niXO0QFRVq1xrgy45G9
7femboT1at1/QuFBs0Jltyriv60kfBKN7pgXYhbx64NLfFkpZ5uTeK6uB3Gg/ImN
3NMzKqbY182j6BlargqbOjtzdKtZOAUqr+hP1jH6siKEoixVpUoasrKfY2ljpssg
ocGPPeXSC5CClzygj0b60bqmAUKnG3nqP9fsw6E0CAKwcRzUkNtrzZ8UchcPIpMt
kcj794fUezOZ+5Z1vHe+4DsUXDc6tY3eC7Vm5BDTD5DeunSINNhRLiHF3b4/fW9X
Kwoib1V79QX1lZH2ZbehhV3h1egK9/QIJSWM2ZcJ5aXdNv23aomCFB8lTkn4S5iA
Q4Hz3UHs7n+1JkyQbcDJfMuXkBdjxnXh0O6yBTOcmiSeWsSJStZnIne6MMRLcCFs
eSeQEVICsJ3Vvnn0buG4t3Abr8dAzdY2pggqSYb8MjWcC7RAUPAzXFH/89Rw+Ytl
5xRSWdsNTa6MVu9BCGzIpnOCUp6Pbeevmc98kYjgsoqCSzYOMxw2HKcQeWLmDFk2
cwrd+M09Mo8R/vYtaQdkUXVJ71lwZcyR2nLHq/DDOqZIOx52SXuJ2xVRwSkmPemR
MWbm1dT09QzeSQWX4X1hdbJlGSYMMJb09W9oX6k9hiu+M4XZAgxmm7D0wUXs/6Nz
k5my9AT2OAdB5pcRL0npQDJ0QmnoZFYI4sif46P9Dx/X5k4yxw6kPm8f+F7WzXun
WDcs9UuP1VcBXQL0zN595RfhUqpRLX9zoqO3yecRBL4eInbpu+teSc5y1bZePQVt
ogSLUayti0mM+AjZr8Wmt9E9wcDoG53SZR9q8YhoJKWmhvSbcYaPzzMopZNaafH7
nRsuO099876AHynDfm4WgV3MYGVit4ceQ1Pju6SkD01kFCyKIe/siG+tBDjPHAoj
i5+Xiwrm1tvwBnadNG9dwzKPOX3lPbvFJClPd3ONDBllXuAlh8TGbPkgb2eqh/kO
JogdK947Au8fLqarm2Dl+qrjFU2Ao36UhZ8wfbDgvsRqFYoA6AwcxvNA0TPr3a2g
QRbpKHihJk1hF9yOWzgTEPjjq/kfqG7b1NAh+LoJlqiZol0vrrS+wuIWylFfJpXC
uDGFeDVNC4xN990/jkwjXt1csxjvfLXVfSYrzNwqtehXUMhPckDmiVLZ6j0zmM7T
SbQhNQAyD7x3dEJxN/3DClqiOL3FJy9OLSka2kiCS/CMC5st5rFBoDTPMMf7mAeA
G9f8knMTOi0Fq0sNwIlmGlEmrIOpxTUJTLd7WQq2eY6VZXkCP9LVxi4dNy+/It3Z
YEOV7obiZed68Lba7DSXruhYLpbSGZiCfb9+bgKpQ0i1HFoMzFoez6xHLq6O4w5T
MyIozWbcuMdFOKvO/elhXPQiOHuu6YVplO7mMyzv+F+/tBzX0d50FcACGqT7G3Rn
9FgfyDPDPNEDYbEFy0Q3U0EpweuncGJG7qjNlp6zahQp8DI5fadhV6fLC9sX2kPp
VUGoshq8sEAu63+NCvGay9dYgWW4EaEySBWAkKvPh02oOjjTM/10blGNIIsUH+QE
vxUf4Z4QQ3nfBKsnd9nI6IvtEw7Nm7zel/D1dlCpQS4ezAt0t3m0FRX+y8TTMMIB
OdxgMTzw2pZ2ktxakwJe0KPztHmWIRPOcuEAarlWS9LJFHiawZkUIlsWs2gofRfW
uwvfCoPe8D3+1gzVarpgcbUeWSiclsBBwjllkmGXIzA0zwldOYZjvIx6uUNdBfve
mE4Dz60cc6KbVTLT00zrA+fhCzybR6aBKRMmVvI6PKplIZTCTkl9S9o1RF7tfbpT
UU3qj0KHVnB/eiF8PnrO93au8YDkkjSVhHdznBNAa2fSg9cCPPWJMCOcE/fXRpI0
SJNUcE/hys2QBjoCtGWa9175cg0791xuiqxfkBgmXLzV+jG6XWXfjhpemdcfBJj+
ioPHtHtq/NDMsiCgyL82WEtFDM5Rto7106N1ZF1dhy2QOsCDGjzWa1xSdZXbD+ac
UDaO9KwIrdoShN25XRw0ryuYAZJqnPjgBzCqflfPP6QoghBHZd6dMYDr8dMvD2N8
xZ8T15SInG8fofgCom5wpMbYittDubrGELAIMKbbOoIXcnbMyP/6bYGcML2oyliH
kDa4wi5KC1uoam/Pp1IrUlRFOVOj6/SAZKtruxe9jgfiEWZMUrcUkJ2pezGOP5QQ
aYcLDYUOQxUQUcGNNdKzwAEEFKMR2sjSBi35yKlc5+yjUO3XkCpZ9TgQBwJRV0Rh
ad4Wl5aF8agi+3FQ7wu2elXuL8SLcGRKCZ06cL0fI8alk3OPl0GulqgVIMyy1F7K
HWzjOv6N6uHDnCnnn+CcKKbTIZI8gYZqzeEylXUmxddRTnhagx3hZxgSrBmQmdjD
tsB61rwTSmd/nrfD39fr2c7dx+/BrtYxNiSH+c6LtdmX1JfCf+NJttW9DNxnjjFC
Je4MqFM0ajnKC9TxxM0RQ3lIxomO08SFMnIzwdv0lny6+PRnCk/sGk50SRE8i3IO
AdfFW5KV37iFF5MxArLCHhQKfYSjkG8eZEqfoflozOoduraGniuRhaDgj7GPrztW
8/CbeC1zybeVX+Nzj9+qBdE5eqVF1KaGfRU8Pu9LTxibpQs8X4vD/nahSFP5Ty1M
U8Snqt1DhAi61qLBg192NTkabnBmgLQ+h/2EQGuIBaCSSRdWtmUSzLu4lFTcmTmn
WjM07ww50e3N/oJ8PpddDFtOjX/UDAw+AjEWMbhz1XJVPvRHq+7jtC1CuCShIwOv
ajtqOfCIqe4kzzW+Rht8ymRuJyzvg3Au2iJeRcFr3EvMwXJ5vSUgg6SS2TWFxs/0
4CixAzaZD1GRJZkUwE6nfcZljFlvCzXk31wS7IZEwPXVnyBFFDXrQ6J0GQeZFVYL
uE0nTr9HKjRLNHSlyb6ROxH4J3NEka0EmhcKD7P6oerPAjuQwW/2dYEC8q1v5P+z
1GiJyS33E4gQNXX0A6vF/e8NRdqG8OK6sLjtEyt59kJ/TQCfu0Nwihu6UohjyJu2
mUZDWuIXBeLH2gB9nI8D9LD8PqroX1OYKbhG7FCTfy9qYTTCgpPGqpduVbWWAd8+
qTI+bNOK74efhrSvPauiIvQRK/ScdxlYcelKmEjaemRE17/JceLyxCSr1hXPC16C
705c1f9/Id7eCs33BkU/47cNJj3W4At93bIH3XA5QBPfd8PmC7ulKZM326pI/Nqg
6NWIHmVqeAaq3D8QP3xgpcYJl2SCGWi+uD0qgf6DIeq2Dnra7p6wQ5slZS45V1HA
kJDYF8HyCX4+2KdgmstPpI56HcKZMXYfwreh21gRzpWpxkT9+Bvc0uFmPZMLF9l+
XL8KxSsY22KrOJbvnH0h/hJeP4dWETRvZiqInry6pmOd2PGn3b3z2/NGf1XPphEW
8BzUkEGK47x/5XbgNh3k2Snywgjr6H5XxI+gH1v0i7ISTRojlVvDx83gZ4Z+7v7b
fuFbKUPjrq2+nDqER6WbSD2dHHmKhJujs5cmqcyqrZcq3lfDNKoxf8kgAcCyVGgZ
KrgtBBU4svqrRtQfDsqkjZsw3AuuYqWK5bkhM5m4v0wAtu36y/5U++UYDJxJN2iT
Yizsz99iexu24FmOJepq/NYIhQc6NaNVp0qrGqKAHESOzkpP8+BLNZBOIyOiWujr
xXCj+DN6cBi43fiBpIysFOaWbxxB4r7raWpXK5MZVMNdw5898U3gUUQUCbsx9oZI
4jUTmrK5z0spyavzxz4xU444Xxin/PqhoWhbuqv1ngEIhjGlVoHbAgiFaKwBvjj+
ghr9KgQJ6Lu93etRjIrgQyMPDn35u96t+fl0YgQ/6qVpmvt11rRy13dWEweW70R3
DKzpgnkLuC39TNEFWr86SiKI8v1GGdjnCK111hvZ38aJMwurDht/PZxeD/MuFfj4
hT03TMEF7GgkaxjY1vrXkGcTsB1vX/ds3/Xd9cN7+z6F2YoMLcvARqD/4Xnsb+Lj
m6CeAsH7n/gE8PDu86iVtyFrdYO1Md3pBX1RcacyjEmDBvOdCtrv71HMvP8iyjFW
aE2Df04WDgSJz+nS5ZF/SJLsXk7BNE4eMkufx9vLd6G8haN3H/nutRrbVNzKArkv
6/qSWovjiqNuoRL1PIJ/yR824muTeARWkxDGi+bAGpZHbAzKk0DuGOlZc0DyMyS3
kHuRIoaZiXLFKtQmeM0HcGg2NUVmTUyfskgx6BIHvzoNWK/NBvmXEgl/4o5LxZYH
vjSxhg9V/LqHXauygoQ30IRh1HauZF6Rdf1rk1DIgBW8PkFMyQRPY4eR8aKGvgwC
lUvVl21slhEdaj9W94vLBfa0MY8PzrsCqhQ2pXBeYaLVoFL6cET2s/3r5sg5MyYH
bBbIbRuzogxGWHr/k0D+dTpEFPu6abbnoqeLFn1D9uRO81lhvh4pxI+mqac+98+D
/fVTOdtACeKPWHswu9Gvn+rp8L8eI9kWSwLF8hGwABe1QYOq58xby51C/KTgsuY0
1nkiHt5lhskeArZJikO2d+rxsQANNWkFMiqoDicL1gCrqgzKdxdRYdX3CMHZ7BCe
9tXMTKhnV0SJU+m86W2IezFQ3cU23R8hWgFYCASd25Q5t7ODvM1sWSlGo9HwpbKz
ZkaTG5JGfaDZem9pV21NzdL9Xa7fPFHao530+WGdvTjTm12e4rLKMzT6qD0bhRyO
coxUbxZamnESz9Xc6Q9mV+sZ6ybEgs6tDX57T1x60vIR7chytZJf31/MQWtRJ2gA
y//I+fGLTZ7jvljSvdjlwsNlUUsjv5y5wMxg2xTxan9ebAo89Zl7iloi0chpOITR
Y4gfUeQ18dProsi3Tp4uXNO9qnYbPZ0KDQ6A0XcVi/igXh5OQVW+RdyAZHu12x/M
U3czWi5CRhNpDuwP6xELwRkbf2iKdN4SxQ83QvqAiK/5tyom/a75WFwMmAwgWN8a
UGtCbWFBHoU7utroBZJeufgawjVeq54TRWn02FM8Kw9thixBWYC44Jxctn8vUmRT
pVupE/k8Dhl/7D6NBhIai2H078Pi6NbpWA9OKxgEn8nVyneo3B+ruQxFdljTP8CX
OtRqOGhDoetiD+fHLb5JRfC1nGMKn3kDSBuoRjA0fDPD0Xx6ROZt9w4KNeBzLaaE
mS+395DWyMcK4OnEWahNeQPeNLWpRn8MWJ/l5O0bpPTRy+kLCFwytpY87xv57YFc
yqb+y9cFtjIsMCx81Ey3rV5vlAR7i8anGvspCgtbZuxVsx4ScNyOwt3tFWFS2ph+
lPSmpL5YZ8CfKCRIapvgtZphFJDBMrKk4CdaL5Z1mR58K/tHiVIF+fabvGX/p6Io
krBXak8sbQ/o+1MtfMV5TfTiPjlrEW5kw79+5FmDd6hde17xDANkyZ5L+NU44OFD
owx2q7ZAIA4DzYjpT4HCzG3EEPALWdyeIVRZ4H+ScNddLmdKUh1XQM+/AweZX6+Y
DK6p6q9f7/dnx8qDcuyPrOCnnKLULIISszxniN91EDqNOrfWtX5a3MzbaYSNwU++
2VwgR4ZLQrAcYE4vUj9f3aJg7d4LTFmUoSgOJgBzsiePhQL7ddv6gcNEeDIsr6uL
z9yPUzJ/l/TQ1GN+heFzhWoHC/sb/sH8B5fjP5T/8EsuH00KwXjFFI1W7jLinfXr
zsJBAEyqaaL+oSoByYVSOP5dhc8Us75OqR7B6uBwUhC2g7Nrz/Z4jseGkagcH2EB
BxHXn8tqotIEfiwAlMm1GG5qrGCpPFjQPxzkUFYUl5dkZvqQ1dFLxr+xy/y7ThKz
6hMXq4fZVcRzE3YFUshTr81WXFEvB8BTsdiB2f+A0ebteF/fMjFaVDWHsrC4nxaa
kBgYOFGjre8GriluJW3sycKSOtrbQnW/PUQsqgkTm7jYPQjPPDa7EE1w9IlIPkdU
E9ixfua5rrMkv+2LzMgDYHrNlqk1rm2TXo3s3nwW61M6V8ZgsDukvBKgZbaQ5zAI
DzxqRckleQy/x6PCCbbfLOJk/WoxpLBJ9kl9610ikMUyytl54LtTlr1atGLZ0JzF
HzfMDM9/9OC5yHZQgSJArZ5/vuha3MW+OpbpUO/rIzWxAl6v1spqMQQoBK1cCykt
AsO+9m/vsPxe0wbFB1wjclW9kjxohnOWQyoxK4QPFZP/e5s4h+D8wneZyygTDnnx
iAlY+dxihazYrLa/BYs9jvIqawjK5uopUr+LeFylk6S58sQx2Gp/cwouZM82MKm/
RbYZMu0YWy6AdtOtINMhdV5Q283/QM2Nlj6QDOapaQynGQm4cmeT+WZyDt7YpEVQ
SZOxnKc14yBHfDpHqodp2ZimZUxqbQpOhmL9HR2lPb4A0m+uy54lVIGwwjd+MnwI
RmuSHhMrbMce+0FpXHYf62uCYi6CCjJAq2fVB7j1+6XK19TBfAFKdEXq6IM4lMKQ
SnrH7o9PEePWCqjWBVwgLLV4tMXPZ2aKnteagGLhErUWOTwi+Rl1BJJIZdt8Ucv+
pxcDk5E5QgzJEQX4Y1Bu6hedXidI7eAZAQUDC+wSzcZyp+wi90MGRnR7HwNCDXLW
oJrgC3XG+vatlkP3X9cYbTQ51VKaPMLAv0hJc8ap5ODPBChCn5lAVUyEpVevVGpe
2WYCsLjr9s+oX+Ya2x8ztOGL8v4+EEGa/EgRP4EvYCUNBqDGE1xktd3ou5sXmoCs
Y6MrnqyxiJPaMBZ6BBfO1n2YbF5r7ez3Ua0TEjccpzwChn7Ffa1kdscPWkI12Epd
7DhiU8en1Ip3NFNudlmBfOd+78PDJvrfnSpK8VkyngwPJR27byawcUpdvIi1gEnD
KkJRq+3dLUOkcFUVOlTjG+ZEKZYMmsvzaedQw66duGHpmpWqu+5n+qhe2JTS/WjQ
QH7MS/b7hb9wbYj7h1OXwUvzhvYcZUlX3jCjnUACEB+AWqFyBDWGRuOXjolQvJUI
DDLWxYrVizPhibBkavVGOzwWxo2Ru43IivyAqG4TSrBUka3O4awqFomet1D4IWij
oU+Hrq/2lA1fLc9TqezQvKc3vSPZAW4hjL6D3G+Uanlqzn6QNc7C2C1HDlJEzsFk
fQuNHAYyCrAKEBAQOfRdbsjzJLsIFinp+TN+HXcxZ1BCZa3RIi5o6zu4/aKqaQqT
Z1pXq4PXi6akyW2wS9rXpQaXVql4BqlGysX50jdDsMVamX0TOItM3k/lddFBb+20
2kjeizvfbpM48aJhnCWcmbL6f1u1/Tv7+mqxTw+dQA2x2799UbI/PwpLFgDf/Qdh
BxQC+GFnmNu5iAzBlCFuBwezKv4nVYElKMQ2ZHYyYoBjGDeV8z3b8SJF7NoF9qB5
6iBuMr1wzZeaEr4/D70KMhdDyMfcOH4yhuKzHp6VmFoEFTcKudyRWTWSqGlCQnSF
l+Mf/y7UES6DQqygyZqUzWQE+AOXjMe3RDBa9T1vfCHZveF1EeHNAGRrs1tLtZBQ
fL5ERaIkhIZotBe91mlYmLYfFhawv8kUsNYqK7AzYthx3Uvvnt4z1Ol13G7fzE7f
YvsuEouGKB+4od53Ga4LDqohYJgY5wD2a2xgtAbCylzZeZ6EKh/8FbhJqRJ82ITf
wjiWEFJpy5Mn0qT3kjqSL8oZrygrhCrkLHD8CvY6CgmM8MnTfUX1J8ag5+JH+wsz
Uz1MOwK+jPLz3pskWuoA0gD/bSYLb/oTGCKGsUwTQZp8MY3XFy7wCIHPTbt3U9u6
nQ36lS2R1iE9KVswyXHZIr1k8KX9tgWKASFtnHyNsy5BP1j/tDWbZoRxJNf6uKsJ
r5gWuUIpYM/o8EHZMqKyoBIAgOJdUNeTf1TslvJFIdjMDHGGYfnT/g2igsO+9LfZ
g5u184eJqK5wJbijt1SHbBEG3IdCSZxX4TVjUw+UJsh+wyJdp4GgHbOJUKl9Vp52
R8g3wBCnR7ZAvaXkme8ej7vDbnQqvvQIsN4bgh764cxPC0TpW02Eh69puqrnCUV3
2TquQmDKTzLle/XQCC5xYIgkNwg6LJkCMalAxXqTnQhvbuZd1gytqqaQ1uIfwG52
IJIYkjTfpknY0cBcaWltwNPtHGaGZEMHGvtWgC/oF11OCVN6CO3RB8hwGPJiDMxR
B95QW5/ztp4v91/hXC3A8X7k7PEsyEVZVKcEQuwBvmKCD7U459uaZeO7+bandeVB
tchuzfntu5ac5NjRWfip+f2fLP27mDLgdj2yRe2YuOZU//F8ZNAuoD33wKQrk7cD
YYezbVUm2k0RZMI0yKpcyQPSai+B2l6ZzYXY7aoHIKctT0qI/TmxIVsFeWUKmZNo
uATtV2AaqyQMMf/J8+poG0JRVUt0IvnJ2aUvrYDEm0Q9blv1RIstbkRFb5Vn/U0K
tQIr2F69qWxuRjxU2DCF+l8OsFoUYB0Xfm15y0SE0zxGiS+I6Pae0dGLspA39O5/
s4sX9KxOSvCYI5L6qf85DBk2iEW1VSwpkFddJa+oW984aPie6E/eE+M2YxVtzvAy
KnydFPSOg5dWvYm2L0Mp9k//9l7mbqmKFTxcLIWzpAi9FEYY8KSZicMfHhXA/B9x
OaN502BRJWZcqu2kF0Sew5iEO2Put6HeSDKKV0P2y6uJe3nCLvbpk5K4ggz6ijTw
GBom/3riybj3MsDVXC3JMAb/T67IYRd4jwD45Du4lFVLllgbL9wF3jlC0CwoDS9R
99WMhuN4606PMZVVP8dBs89UMeCckWDx3C+NKCWUMEBlFPKr8zuDmbDr+JX4z4TY
VfKqNPJOddAL4G2ruYJa1tWgrzYMZlXm5R2UjsLJsltYYiXfCJepyjb3KrewZbtL
MqG4jaacNcYTAPDImJM9RARzNRzte6qxvA8eh9zGJzaoM01YXVqH13xblY1kPrWy
+/mucYld62vkp6jeRzEV+CH9t1yGtyfkdMYxmCpklNJErFRgIytbqrVIlvYqqsYz
/Xk0QvRYYaU7J3pfSY0K1yyLFLZ3r5E1YFtLqrsSFcjnGRW6itwJsTb+qyVhInaM
o6J9QBI7krxR7JWxAGFbgC2bp6Q6eggG5b2tRPFGMudH6zOF4I5vL6En/y6TcEUM
EpLpi3coe0iuAZQGjtqZOILV5+Qpu2IOdBrZaUVNlEQekLdiCg/xAM/LGOZbwXGH
IAWoaKwsAtUBBsDz84+rgwZ26jtp2PrnLPZmfRedcIp5GeHQdtiFe+i4+bJkzZ9y
raJMIYnP7eg2Zxbtk2SGGWnenI4I1KPzZEdvRUZMXL9HYkybkE+nEHLrtgxVGc31
+k7hobkKVh1Dzg1J0MME6QSZBEHOjXsUrpkOKpZBeJqPXnJeojpJOSJMSj9DEDx7
cmhkWcpL3q4GR29oPBLrRTTzmVfCq1PioxZb/VcX/FL0d3/OfhUHhK2VxJgmx6Hu
G272OBsnA3NkNkyIwmmgIeUFM5WkVeEEsme47Nr/buHWFwZdgm9s5pKnw3r5ijjM
Y0+qAvDO1mQnfG56PGGm6N5SZbpHL7+VAC3QmebwEye7tvUCE+qLo9VuNw0XbAp2
4S3SaOpjrKpdeSuY5okU+e7RxltJZQ6pgi/WlCpp4YhMzLy22A9Wys7CUe5Pkr5a
WGOq1jWSDOsAY8psuXkQkLTJf43+Y2wQBCO+h1SuxPpK1n5FX/xmL6pxEoB+gzAF
h+Uz/XvGPFc0FRUamtZI6yA+xwcz7Y0lAjvOlAvDAqk6Z/L3GQ6Wp6Hf89BtZWua
5WGU8ml8L8Sc/TvqJSL0wj281fOI9u7e51iwp3LzaWnqRXmNXInEDTSSEXeK7RdB
m5z+nXSd8p9uqujUTTzzMH1l/fWzpHt/Erj/j+lmAS4x8qZmQmwW+KzPOOD5P3z9
6xODp6brUwlSotdfpGlzHrqVMrOrSMEbXO1X1mhlkXmi2+yj90WNnWjMgnksPSEM
MDhM7+j+3HVlY2lOAlDoTa/aZMlscSxla8hEli0lNarIOcAE/q5fqA0beeqbAF0q
7lFXV4J/UwkMUwGLlj75baJPxL1QjvvYUgJfx3H+VVaajLQYuDmbDGwNI0QKoUai
rCor3Jon2M8mSNGobZBrKwG7SxGQwulo5Plzx60NMskE9GNZpEos+1JxbRuwGF1u
SzRwRtKZWvwQLa8KzVYxiN2TPqP+5lPt1VMcvw1J3vdalHAdXZCDKl8xLvlDjahh
F7ELnwRe5GyVSIHNsw3EJ9lVo9OPRsQgxcyqK+EC+wM1LJjGRw3yUvHmKabqXw/t
vp3NHJ++1NH3ZHiG/qarfyEbDeUKLOFmRUTo5BBB9zKV2H7e9/YE7pf2jEcBc2YA
uGwE4ZZRoa69LRQbnfGDooga4lPQDT7QEwk0OZAoYqQg3ABK+BgnmROoVVffa3XA
qxkfoEV7DFBXey20fQ3dVWIwIZyG6BjYqcPUld+yxBxiWlY8U9sPPTMpVxZjyTu7
hxwFRkDrgquM2mwR5v0igLBzv1XtYU5o/aI+EY1fMaHn8UaDKGIelLUe2ZvZ47MK
WVi05qxj8YSGn9AAnucHqxcDctIThUcOBmysFBivX83nDU3OTWtrrWhS+7DZMP+4
v3t967+5FSuv8h3gmteHfDctkQMvcyv4SgQw2cMBf6JGo3c1mgYmuSVfq0W46zsi
6m0Eusjg4XX9tuZTDL6hhEZXxfAdOgAhIKaqWO6Wb5oS9MWWoo6GDmyl7PFJgl2g
e9j7R6tiudKRnnJbC35Lcr91OVfmbqR5L/Xub1UjgGvuKbPhnrCVw/Zb2Dvy1Jc+
9V4SB07dNahzRZ+0WYpdQpBZt+XDtoeUdNToi5AgRfftcH2ifWyzkoKlCuypnPTC
H8Kr9OulOnglTUtCvgmPEzd5DoJZ3psSp4gDht6FeRIqhtWT5ySfLuMPUellxn0l
fH5cD2ZBarGDEjU2Zl3hKNSITxISNzhbDFHGVMS87FxN2VIjqcewTpd6Zvf+M88Y
cDbMiyiAqZ/PlVUf2eTlK3qcfPq2xfm/MT+fNrzEdinp/gTFEgxTHemNc1ZAf+nI
IrZCEmDzSxkGVkOyBYhOuH2+5AMgoT1/QfK/JXImBunw2RqwzD53igZu7KJcrxy0
ckyTiDV6EbmLRoecidMzkXR9frNihvmyM5hJarhrXuCXGFmzRrcVr6y3VaB32Alb
3lIfvSw1PpsCnZ7MN4vxkHljZ92+u254y4Ulc4DfkXQvmH9XkLoI9vFnpw4JSPnz
fQoN8deSXYztamgK9uRfi561dLB5iRd3DorvGHgitnG6UsjrAkpfSSzAzRA7xbYg
03jIif+n4D4xkA0UQ0xml6WAgzIP7MIoYqRk0d9oMDaFYZwBQIQEhbgVRGCGOugN
3mA9RYIOrUkBpIND+46xakQvmMbHUB9UZbhWqfChTBtXyLTw+qcevda0Q0tRHHew
3NDjTYyQkB4Mux0Tn6+1PYdgmlQcjutH2pWNPeMDs2+nlneIUHUajzaa5xAFnw3L
E8L0O33U7YUWyHYjML8sEfGoKJZ3u7uti4/a/ZsgKi5HPcEpomMD2c25uRgJlRJU
XsQpuy/y6WYqlbwcqxbnipLL2tnB9jk760V+xWgqqxPst6G4zvsYBxj5awENlK+e
iobx5G/IAaQxvaFb9eRPH5hVJRqsLugfU444Ugcc9z69eDv7EjB9JG2GHxXnYqaI
1871Y8FRKkSETIfPDuYjjYJaOJtuLuHvG4Cg4AH0REfclALA1pr8oO3JyWUlsxak
M3za706slxLgo8Nv/JaTd6xxe+j8z8/A1TkJQNYROT4wa4Civqej9weBhdiN52qX
tOEYM/VJTaPtR+pPTnvGG0QT7/ruNEBkxBumivw4fOqGdQSLTgY/6XWyWCgcGbCW
y9rFBtYPUJXbS/mmCLVj0yiPPqqOStK1QZ7WGYafVxgJqrE660KlIDzbMORc4HAY
KMjep9I+WBzoB/d7IG83vm0hiAbEjrbFTlnRbIOGtbF4PmMEGcZFB/p7WZFHgTCg
qlZRD1hMQ3TNhCKA2aK2P3fDIk36q+f8el9bRnsAH6qnLB5m+H6CwFCfMi9JUl5h
wqX5JxMvSpAohuUOVFIR7JqwJeY/7RoY2uleMM7aJE7EEMrdVUzSm/nQ9ew9C4xE
/zPFYWc5lbXj89VQcWGI5hznuJeC36Ic3M0A9hVvY/wxIWuB/cY7rYK/3DhTl8iB
R8nO2ihSHJ+6DCWODYxo6tXwRqWkqdThN+G4Omt4bk+D8vTZRAeJO4Fp9R9RCCzz
/1gHSEF22Vab9MN25qgH6A2iFJ+S+BMROuUL1f24FxbFG54IeoB8iAjzCKsi2DxW
hYMcEjPGgh2AygcEZ1ozWkX6H9FTCPTX5SvUAIr4Bm+N/cKTTrmTt7e5TIQXxQcH
aUS2lpDrPgLARrxnqB4GE01efrJ6o3YfRSs1EJQRFihGYUXq/Kq5jcwPeGDDgtnK
mYwsksZBriXSIyH6rbGzSf9F+cZykmY0yJWywJXbrNS/iotZXyej+hbZy0NlZF1t
XH19oqoPLLJtYj94+Dq6H7zfdtEl6qgap2tZYYisma5bJkAZoEJ6I0XgN9BsLOeP
pGezvMCT0dyuOSJBsxI69Bo310QcZAD3Zmzu4mecfLJWVXIpWnUCiuk4Y02/Wtc6
NEWDxZ2npZk/+OIMhLWuywvT0gq0VSMgwKQuCbOvUXEMPqCjfMgUd0ribEyCrLAU
ZZTEyLHBxWrd6ShM/wd9p88pnIa87t7fkuNufZoAF/5nXp+P4XIZDpuOG09bAFyD
frzhVlcW0XlMt2U1hP1jef7B1tnluRiC2Ve8KoufRG0xOzPUuJJMCXbohfVzNT/l
/wK1syi2q70Bg/RKS2C2GnB9u5FYy7NCczf8OOIXcgcUeZ3Scx8iQhZPqZD3x1uS
1DEekZtbzr6rRrYUauuMySBagkV2HF67Cw2pxJidlytYE+35Q2quviJe+QoFwkUL
OBV4fcknOzMQcXmPH2+1DUEp3lFUXOik27hlr+OD9FZjKD36FI3vtLRoCz/pfiM9
b91nGB1/fVyrFEEJkldwNmdSeAraiRCJW6ystsXTSqd2Jsn0we+nvE9mSmCmX5ju
opNQ51x2NihbToyUhbrq9URhxK+jupZfCjkNAl4RsEHVazlDIDif6XOXupprCpPR
c5FsZJKbtTfsZvHGv8gXH+ngpIvL2JR/x6jbeXA2GLXCSfMO9tIX9S2Fg6+CB3Zm
V8a8wjQ5TmsIh7yP9qxzwIKYCzu8jm4b95PHK8bxrBfLWKyWZl/fY54Hfl9IFSCR
zF2ECx5jCYM28DsSn73Ajkb9k85O/lLAEc6hTalBzHLcdzksVIrfAzMEMwHaXrx9
MfYI6gXJ2tQqkNkeFnKc3ouludnWMSHbSb6Bpr5oHLEbsztK5VUv2yjDV7JlTBoc
cYVbcR3+ZZAtzhXDKZwrITlEOxJeKi5VE78kwGeXnpZ2ZZcO1b1hLPYXQNUE22cL
IwsK9sxIVjm35dn6ieUvW6XskwsXoM1mbQjDuWLeeCFD6Utw4cunquapDTxJ5wga
c12SfswZGcThnk6ZuWmLlrJyy41i4stpVwLk4bHrh24wc/GZQ4BTVR3SKBqluuuY
GT8FVpzAY/3aSuqSenb19EZXYY7WtqLm+bnn5aG3y3FG8VywnW/SwIWvLxm1oRCV
Pqi6cChJv6W3bcjKPyI4bH6oFqg9ro4PfgK4WEFgdLSOIOS4oKQomQf+KlMBY/m3
8HqOV7ZFvOIFmp4KmRLyIuFvr2LZIN97v+y6pxD9n3WPhkm4KBZV1+4uN7a3yay7
VTsF0GqGgL3O0cjIDM5qtvzlgyaH9Q3VZ6SvNSIoDWbK2t5+HkK53YPzsBYuh4gy
LXywqZGDe+iQh9aebVsIFDw31FRTsAnIXBe8rIJNQielUv0OWNUE8JD/BxzOP3vw
FKTUv8dWrKXE5alTlBithvaCmtbDeRljZYX9mFXZOHCLo2cDCkKET3v/w41GqK78
h+o9Nm6t2Yp9WXrhvIVCK1gqZ3hz2QH7E1W6G+e1n28w1d3v/+pnuGLBdx/dUltl
0wu3OY9St1gJ0y1ad809HA8QNra4FYVKbd8Rbo6nwUI4sjGhhxCIf59P7fZ9O6+B
EM0HhxS5I281Zafk7GOSWV131yurgldcaRO/RZyMuLfeeEbDNJ4S7vSlVddzx1WS
WYaak8sAn4VIU9Up7P1HD2nIGxSYIRBjgWY00G+tWJ2bVmoyofw4PwoQPVLzahTz
yGdYzExwHh6WTpiMoEAZyuKbWMVjNBpMiqjvAuTBZ6/nVrbT5/w25m425IPqYlJT
7vkhGGFsDJ59PAMR5iwuYF68aMdOtvsuD5EQo/DLjtJR56+k9RP6mJZS6X70cs7w
xm7gT583HUBYnhQy12XJEERhvWP8iRxSGEHZ2b3SubkJlfPXQkhjdhDBkRXS+k6T
VImmSieZgyEKBZBGT5KnJZ0tOK8jrm4f86E3gKroncpmvqLlKJ8qup4IMTA1n46P
fAEnIfIp8vMrBSA3F+s/WbwtBrnO3sScHmo3QlNUWcaQYXi8+OnfBdz2ZsXJGvNz
176BMji61f+ckh6509EXV2Yynit1vLWa2TERbIMKuKxCTji1LxyifylH+b+/2V0K
Y9Cssq7HJPwnDQMPuIpJBr9+rafKH4w/LWe8GzsLq3NEV1dNsboncyoZ9SnFzAfV
qG3MKSCJ9K6NSiDDSdFhWvzjpeWaanWhzruRcW2JLSTCaZCLOZM4QJLddCmw+fJ/
NsQRz2u3glhEvTFDYGHXP2rjSEZ3gvUTH/7ikDhaw0WzGhlP3e7VcVLDtcNq1H3M
kGNkwIMNUq89i6b2NUeY4M/WYLp0ItRcsL8lYuXQ394TuGDZVBXe6GhxF9NezfZA
MzVYUw2vK5P+vmCHGEHTwkSTUms3MlX82A1YjNAMa0DqPbhbTns4pViE0aLJ+v4Y
av3TsCu3wb2uQsK7RGM6y/guD14no52aswCWbVBc8axjrqlyPOXlJxdEYwKbifYO
xtYdyGkCaN/Pe8e0Viv5gTb0FMHTj6U6MqX1ksKFwOr7WBUDRG3qGSNcoBaPQ+y1
lLj2QCFMyVK0kbbzHXgCgjRZKk2sTHowzmokltZpQY0ic5wCJcMDe5pte4LSCJ/v
clCUGLuNzFnJwSGZEl2pnqGU95dqgQgbQ0DUshMH3ej4dRnGOf5zRIeciea+2HWm
rhDp5SYQDO4+uxfBPIpXrM/Syz2157YS83ISit6TuzO4CWjv8kMyZnvMttIQzQIY
x8hfxqOaJMn0hIo1zgIIiwRDpWEOzdN+Ck1ByGdEyTJCJ3q8Sh1nHngvFzewoVLY
s9f6hHzoe/gpZDBmX3IjTcQG2MHu+6PD2NWIXHmuHUvYYHEh3nbcVny/ioPP3Ct/
4AuNeER5yjLwRb8HqrBlP6XfCwbVBFRhxXJh1tPVzrPC+2aOeI9OHozNkEhP9g18
skfP/Nf/gDD1fX+/Hv5+mQF1bn0d0WDD4dVPXG+1nyujrvKCSYDKfZto3KEkXPPY
Jn1sNS3TMU/qAfeEXpFfn93d4zWO/6YED0zfynfs3gjxGG7iK1GmHjIP0QWDujRy
0NBlrgknBOuU0W2PjvbHoZAzd+embgxKPRlxVn79oZCdpnBYB/JGluMjBKgQKUVt
tU2YDCjkki2DrUXmmeROOMhVUmYVT6hdn/eYBfB+0qzzZzsealIvKFYHd6+Jt4kU
j05bVLL5GuOZaZSOBbnIGDO35cuuAbJ/HqOjntwVwtpN5L1+4Kbrsy3CplW/YcU5
DufEk+9jURtIFqsHa1CGqvfSVctdSVp7P/YiL6P4LYfro1D63PmBZefSMn+t7coE
zkUAwEzWk2mgCf5CZ9RvSUHAWc8rxekyemBwGSjPwgAwVBMJUc82uA2Sh4Fg1wNo
IFzFpL5KJGpcxzVZrGWzVl2NS+4eByW3JObDmPwEKEK4ZVycctulzqSGwLwZ1G9m
FuK1dYCQPtHQzyOsj+HTtruzQdBsNOgswnfj+XoPcS+L8i1tGazjQ23iP1b7pkaR
3D1IXzqQARW0bPuz1yFFioNlqHT7zBCzh41QsiOtUQiQXBcRnXQnoRBMKtwx0m2M
E8lNjZVpoA44PL7QeaCESzjQ0HY1RGkdNBb4bF1QyaQV2R433Jk5PAhDp0Ha5ts5
vJKG+lap2dTb2wRLhOF8P4BaN9RwVg5g++bWGVT0GICzIV+i7VDn+cS4yZrldoVj
JZTGKtFDh4UW35JX4v251L3ZcMRdd7AP0BcOpbkIG/W+5xb7dGt9PSyfNCLN6tCG
mV99V2yLdZa8uZ2RFIFcI4ZxU0dinkHhqDUAvVUI5k0W4eYQXb2CBkNf0zT8GOxy
D38g+6SNq/rPhDNxyRAgaElDV62aInIF8SlisYsm7WtgA3QpteUusXhHIGxvk2lI
80VykaqtIluiYoi4z9JPZvKwCGFn+QWcaeQe7rhhL1fLomH9r+YmteaGk5HzdLUl
uJmxELOyOVjA4MMxfG/8ZUXGJeFUwnF6KVI3RZwEb3op263v5qA1JYxhDEjO4e9A
G4zNzX1DFA3MLTZjBEGaVlC+V9lwfHrJT9/1WfB/SZBzt3qQsqT+0VSak2mqWkf+
o71e0AbpBGP6bw3UK2d/xPeFDSoUeJbapzU04WsP9Srcxzcjs8Ch/52Q1gCVGYST
LT9ze8x+BZKX7CLSUWswNG5gvFht9kA8rhzs59nFxDyghnfxA7cjyRBVSdWiAktf
oIJZOa3J+qBbpHzhJszj4H1q24r2xG8xq2mDykj4Vq+e0akQI7myiJ+lyUlKF5MU
SelScB5Q4EpZF6GcLfcxDnMYvKbrhcLwWVEL2F5bnSkgDFwHAWdt+2S8Ac0jkuPa
CfboCoAJgAJUqr83LvnUVCN3Ausfz3tMjNChOvQELDVE1eFl/p6lN71lZ0vkjAP+
L8H76/ScvBlbJ0E2OVoF6Dam1sq7o8Bt/lCpC85Fj1Hj1HGNFoSdLENSBNVvMxZ3
nRSYl3RqwrKKG+pvu7U1DcNG1tpxYTzeX2EFPU4jqJtwC9y+TDmQiJKbRqExKc7n
qG4SXvp224V9oAa+LmGSC49SxJPqyksZOUxESv/01gsAlv0kF1cehKpxT6TTccu8
cz/D+x76Ier6weAwSrp4LJ7BrsRsxaomFjekNvLlsz1A3gcZNvbx56593h6uG0Kq
a8VhoxLmpnU57Qe8PbAuWDCN6G9JK/2/lHAaOLhNkR86qgJ45psO9/19YtZVLIKL
9d4LA8AcjcV/RTRMmkWqLy4n83qm6ABOiOUBMMfdg+LGyzAOaAdwBCiSoRxi4YvR
7frwmXdi43DkZNHvhJNHzRAUA/y05Xw8R8+hqSUv+vl1pHNRLGxHGdV0HOzNCoRp
G1yHHf0JaR8oOnoECMk0/+/6FZnoHE09a6MczodyG4r/gu80J3FMEDwOqMtv+ZCK
xxuejqDlm8ZAaYqzbQNbrtrSVyOcC9TnbRFB4ftA+ZfSBbHbNIVHSU00LUeQpAJN
oSFOc21xvWyHOVyXNjFCqN6zS5eHlBV3lyrTGc1kW2JEwIkS/0I0RWBiCekjW1xj
DK8pljIVR95yVYxFbIFUuEwd38xyVtnI0Vakdhg4jWN3JvM09AHQVvfk+K2RWY4X
3ynnz8gn5b890c0L5vjefiWOnjJvdniR+AZCL7StxFsdVxshtLdMfyoZriZmZFck
o/vEvaehDhdT6cQvl6CoCKVUF6Q6v6v8PNWoY/RIvp7HLsG4PpTfWwJawg1Qd7DH
Aar0uDnCCWTqon3N8hr9QGrB5GS9MnLvB5L0Fx/qgz1T3nLVGBaIZLGNBXKh9BDJ
+61fVP1Dvh3ILJe3CtbcGXWicZ3DyAugIYkQtPutAhRZAH0ycsL3IyEkbArPvA6t
rUZoPM9gDtTIxtEMilDbPWIST5RJWtaL0rnOrYrWpFb/m5MwTNkRpy5UKPhenMAU
YzxiqN3hCUgdTAAobdLUFScyaQIbSYI6tKuahprTGEsm3xyWZ/0PSrEb/yq27bzk
QDaaKZ/S0WVmMa+b0UVn62pO1QmlYI1FU7FQavW75/0mwij/fLFvB1NwX0kAtsWw
ox8hZuoyoDTBMf7emi4JZaUgI94EBq0SBnVQgKhGOc6cw4BHBtpQo8qjwG/6NZb+
K2fM+avcbxZyLSOiMPDVE4Eqr0ry+pabVhBrXODlyeWELBMawINw8oUjrDVmK5nS
rxYlNNn8ipGlPnXWqVAIUa10f0HcBWkutzqAIJ6hiURvOtoI4Bk2Lh+KDxJRQGyT
hShB6OtChTnkRlR9OEhAYvN/rE1xuMrU7Vl6a7Zl5J3oPb/xwg5/p7NErmWgtlpZ
wePNVB/d9JJh8lSg4eUuPP33qzEFDqF8d4/dKvLBGmnCw3qL7VnXudLQc+ZfUMq6
2HQ1eC9brsD9YbmOdp8Hc5EdHfGyZGOPV+ktmcAbdvobmClu8Axw/7AFUkoDo3vv
nbJs1BhIWiJTCHeH9OgK+wep9NpGySmwvrivzxSvTvxQH3xdtyMuSabbChB0yuvc
BzWpj7+ELnnrddx6P1K0hN2P3T5RBxD5NxXMt691RQbwU0tAT1CoUW6i11rQJmZg
uFUE9qVmQGYwnFZL6y0MyE7/q2qv6dP0opgotwHQ+cimw9qXMFlNAyxunEKnaQD/
/ypIzolGci7BxM6J0SmLa004kldovFqZoi5UWST+09dl/Un6Ibu0M2i1TPqU9YnV
+F6amzis2OgwKVEPw+m4Ox7Qzx+rhtV/BEMV8qj6oO0IlTmDpmeQ0HZQeyJB1uUe
wIsvDEOyISy+1lcGDYNNorX1mMLqoLX4lYsqy78ryVnIHsjHl0b/SPXMqxJMLdk3
DSagr/F46z3MqENcetDl0aLiTmpIfFcxj/s+hsYqKwnSt2/0VKXNPscCbuMNXNxB
d9qnTW6MkcNWJx8UUn1n+QQDFPYRQF/pJeojjXmxJQ+PnG3qpuIY/U5dJyrgPH8M
9hIY3T/nRDQ94LZN0uL3fkebfz++515YvbnyzfgOzdiiecEzyd2FWWrnliPdRXpC
xMkXJPsxeP7wDGQ/xObSSfKFUxtwgfLUKDTUEhPv48uOHuBgwsjECb2yJoyJ+T7o
NwFZvSPpd1+DIsRhRrFkVqXMk5+3WhNyFpUS7BrNR1tKvNwVjYJGBk9LcR7Mg10A
we8rCgNpYiUuxp26iFnsFI/vZWBkvzXl/k2KqCohZIzqCJH52TTQtYHcOGJD0dVc
PDORNB2P6kVSVCzQlYw7y/BWuxg0jY1wI7YNPWSl8oyAKWzqfeq1EztZF5jOnPsH
pU2xt+58V6Fktz5x3dT+1OfTfEJUvGtPVnI39x06hnwJMsFvfuJ/VmxMtyBFVu4g
APaEvN7ErC7QF7k8tGRptjWywAIlJAY+QwJniObCVC+IzZm1xa9uPfArzrVFRzN5
+cLMODRiMFM+TYK4gGpeRBYj9MJGHcVpQojxr1930jJOJ3KCpfm6en8qrABFQ+3B
s3Z/S+NPATUEzAU58hqWQh02Q/EzrTGc/bpEc9W1FOeDAjZjEaiEU+LA349oO5vB
+o2b4uRh+tunn0mDrI2DauHg9/AtIpjSz0/cyLD7RofYypOsyg+3Mh9ONFc+enyY
F1eFzCw6uWt7/kjd4AVdFR90mseC5ZZvftPf5ToUmkZNLs1MNh9Kwj9653OSlIdI
OP5Om+8ZD8hcA6TjCc2zcWjQ11ghKN/0d6BPqdksfsNVLtaolHP2Llm0eKfjYxvw
R3cVlhYA2Ajt8mD5ySEOxO8FFTRD8d0jacFGu8JJ9WXnNUaMr2rZaMq8tCnPQsTF
+BJIOn6w0MFQK3NVN0eKwRc/itiC8tg3Gepne1+mYkavFEJXk9bqePNK2pi+3WIS
WfAy/HqbNnEDOP8dlpfyYtXy5r+KugnyqVszs7Xl89bXTPURZo2AsMRIMOhpHCRj
ODfr+0tjqPctzRgLKIIsG8HJVHwiJYPm/iksCaXgKRVyOBokRhXnOtCrPAmldFPf
sm744PK/ohGXaBI8TUD13GJbGCpsA3nZ9/7sNH7NxpsOhc4D0SAht+nQjuguIbPO
0at2zUgwhkCgsGz2nvLFpHJ2mrAhbAIhuCxLOEYdQlsENBx80c3+7tQ05wq6VXsI
EbjNxuAd3x/9VlGDFg+y6gxxD5XNgj9hk0V7e25SD8VervoEdHFzTYCBBY6xRphg
qzzUBMyjtvSm6HnUGy9xFFV25DuCijm29LSazPn3Szgnzup1UIDrABSho6xt2+Jk
9vISflH+mVCSq6YkPRUWgjUgrjEbJza5uf2sMlRHySQ0n02wnVXTRyHreserLIGh
th4Vmxb6dmxKZErc0D1UwJsqF/6Uhn/1a/K3LBxE7YhOKKSfZQbbarNo4dsP9MHS
UF7r77iiHHqwKbNRILcEf02w/SxtlFUZt5UJ3rcf+iOG8E3DOg4vHSkx+PVK+L89
LS36+G5q+c+P9IYgC2lICmZiecNBzTAvsuNsJGk4fRQ92qT9TdHPwJA+uHIHwuyF
T3kiSMAfrxNjpkg5j1Yl0stR/zXP59bPMSo5soVzpDRlzP8nl/O1y8OVaX+75uBf
aDyO5KamwaD+YP3SBDFmYlos2RdurFdqc9hgEsHvQ05sAg5BAPiFUa1pBieITdWZ
gYUUU0lymjvNXfPYTwMOOyNRLE5dQax2LHDDrDNhUVpZcag2XtIc98Yg204cRM+Z
chlYNzXHknDCoq1bWcInXSOcXtKb2W8wU+aUqaR326hKHxiq3SIYwVOt7020lQG6
wUPhFhrdyZ1YGPAVbWg6/3DM/4DqMyrAOuvCQ0a53hBDPVwDzd0zwpK7dOlHOgXI
Ex7K5YGRseY2QS6QpqqLekINrbS+VnL5TcXnpfbWNk8NngoOM6W96sSGYpyGbwn4
kCpGwZXbfNMIdFmOhyW7zpByisgrAdOnccjnieMQRMXUV6CARkz8mG0MzWsi4vXx
I9uRDU1oAMEYF1jLmtd5hUlEXeq+hwWtxRPStuP/nkxfMqDswY9wVBryKnB6KpeM
LBX5ZdNi0GvrKy2K18jJrmiu610pCj9yfYgaqJNGYh3sy5vC76DhMaxaz/7za2XE
bb9qHAY4+SKRrNyuCyujVW6bKeYIhHHHikFHBOLqEmqwtdP3wbSmwIFUwAtEQEUh
VcQPNihROws9gvTz480TbAdfW0mT7xT31qUtupyw49q6vb8bQdVKh9IfV17IiH72
iMhpEEijrl80iIPhoW4Wq1XNpT7QvRTbbbFvPLy2awGjIEuqEROPD540H+uVPnzM
MRxjfbSGROEwcbS5t2xnUcpl9Em+TZPQl/0WC+nc8dMOT6AaA8MDUL+hf2BebgGR
xnsYn6joIhov91NJTEGf1QVHWVrOpVnMBExWuMd3wr2iTUu1mo3P4EA+1Ym82xc5
39c8ygJGO1XVWxW5F0BqGR12OAk00irXh0j08kiksV3J7k8QoDI4I+32n8GZ1HOm
Ucr7K/v5WRv92RWvU5NIv5AF9RWikdjjAXiLA6x/mJTOhhZs5l3HKKRT8xm8YKM4
DwwjFd7wFuBKZzeHNmZ31aB7sSqWOUfHHSbcYm0LlD56REK2hG6erR50JrjBrZXp
9DlPa6LEYi7e5vkHF7ZGe9SzvQQZvB54ga+Exqjx3BMNpVuzm2xFpAkHldJzfI1u
5AjtDvJ+vbGiG5vU4bHcsVew6o6C6QS5bS6uIUCLsRaOXyp6hP4/0AIuxyGP/qnU
AXOqxBKjmnyPdz6EMYOPuT/rrwSA2QxoT5h0TmjNGmmXo824ywbKEGHNWG02iWLT
l6qD+2cpXqmZn59BCphxdv1Q5PxF92+Yut6lddBukFgUzRYXDlq900S2KizU5t51
Lt9QhiEo5G0bFii2fTd+kWHzskFrzmtsNz2GI7PofBtK2GZZAj5jCHc4SrT+V/FX
Jpkni0TnHDlx185uX5NeV8EInAsLAQZ/tNk1d7BPwzeba2KLd+2Why4N5eBoMwOa
6SbUL4IFN2scezDlr0kybe24FUhmyk+V1k9iWBYcSqRCPkma+vGSk/54nvKflSZA
43/tj+JqRgkIOMVanYFlQl2OsyuMwn/7Zus0mg8dd1fpNiaU31HqpSc4OJNcnVUt
LFw6KIDJIso8E3RUNb2EZ+Fatbix6EYsdYLDIaEe68zziz2Oq50Wq0mWbi71ZXIY
dN/EDEJIT8QZBngZFRj8Yym94BlrD8FxU85QpbFs5YthyRQj6aDuv1B78mwRgKax
a7eJVHjR1V974yLHEiDUxtNaHGpayFVgXMs+jHLsELqHApXejYzWLwH0jNNKfANg
ScJ5eSQSQlwP7i1byOgnGlib0duRflN/3+3WIhFda/EOav5gyHwqRinFrQKjJdQv
hS3jpd1Ndk03EFYfwxabaS++9S78ATT2gW6KgxAfeHFEHsXJRJ7FRpZvOQMf2kv8
yutwqPMghAFFoPlav+Khy/gVIz+uykjBdzduC4Og8osngj4rQAU8Eguf5W3D7B0G
ySnmnZeUtXkTxyElyxrDUg65pmyd9s74PZjBtY2p1EGJm4S3BN9bKihIShSFD8vg
zMAoL5HHJQKXxhFEFMt1a06k5WAAxz0PGtMNewxLDX+3u8MqcGX/pfFNjqbmV1HA
Pw6WMstVZmyBMGS65/P2dBczfIVCdTtcJnTbWF1uxjs31ZiAPRV1jNdnfUcE5sry
CFdMwHcwBh3wZ14e+vb6MtCgULRlMwnlLmY9h8aXAiBLSVGIS73oYhdZ56RqFjfv
ZF83Uh0vD27hAgCRkyRDLQ93/CkeGjqntnreI+FPbsQ4U/TtMbuZQtqofMGe4UaP
ovDuThNvWRu4ufuNIsM/cNdF5WO/Re9dEoFvUvxzySySaoMwzizZB44I8b2Trtsv
l7uv00gmh4d/erMCcUbtGKwK1Guc1uEllaDkkKn3wrUlPFMnvX2p9tEKMJ/MlZAH
XSD0OqXLdVCM/zsuX6sJpqphlTcN8h39dQSxmPIodxGJ9OgJ3PDDqu7RQJeVRSSR
Pinhm+qD0z+rlL3uITpkgzb3z2oKgPSDmmT8+cHKvxLMNZ1L/pr9QKrbBadTLTBU
NvBVz9ltMpiy1SWAHKHjl7bfa90D1xoYjJBCY3nIFIOZv5ttnuT5VDZc/7nYbg0d
7AZhja6qpvqTV6F4GDmP/Qfqml0ozDRDAsryIb5qFx1HB7TFah7OHbWnlKTPsTqk
B/t/2XecLLu+IxZcQ/XbEFAdRIgpf9YIb1QCio9x9xGB8l9rMqnEcfKzEvw3S3Fo
yh/FLvvgGkTpa7Iyllrs4v5ERLKGU03opoRct8Tgu0crfYP0ObarMCoJv1WO/Dad
Augx5V8U1tOrdKoPX3GXFDr1kbgRHmd6ZrDUTW8KJHppi3+RA6X8hp4Ud65oo1ND
9F4WHlkUaC2WLuXhmOnlchWLR375fOZLPxyFXMGjZtK80an/+7RFAxLruNoIQzdr
PTH+OxXX02FKW7kBErw0hQgw9FmXDqEYM6yLbjgGRQByo+fFYE19JbGRDCrDA+ZJ
yKNS3326stk7cdipsS60xM+x7efhYAVyZZfEybMNQeLkeRtTGxvAMbF2JpkwLTdb
81Wpz21ioSm+iF2zw8olW83cXJolLSpiOqX9nFZvAfMeS+vQ9yWmQs0rJlR4FYPM
hsWvoRAmcchQNGFhCkaxigV/HVNDkaDuC6m6pdPLl/Y1EwNv/FEJu77VrEE+eE4e
F0sTSOQn9HVCBFvxctHvx41sIb7sRpIqZ6X1gzRFR0HBrkblFfHmFV4M1xrdA09B
2Ha+yi1eRlNmGozi9qYp8YC38EQ3c/Wr5huXcgnYVzxyb0s0Q/LmNhMaGWwGILC5
7fcETxRDKMS61P5/6hsMIsuR+U4IzjuaOcfQK/pe7i2z3DO3fNg7B8mYOpt0FYmT
8lzKvlAYulguTgBKogvBkvAuUg6Oo28s3dttgACdt8Fv9qzuZ6IrY1bnq1hiLrcQ
bfVeVd0SzuamDAkZY0VECgCIpUOfjxj4QFQLAYlDEYzruIuHzt1E2Yv7Bb67/eKG
CrUUXy08e+l+GdTQhY0mPzEmNrKS9Q5ZgPGUuF09umIZfYxSC6vWd7a0RX8WuvGz
2eSb5vngADqj/q7njAITPtvhPz5Zuy2UIf1YxYfWFN6XkQHwHFLyYYy7H8ZyJGkx
OgA50N1ePW1nikiH2R0PvegGtRYvd+FplVfBFml9Ee8Tz15wLBAuQHhyEvbUSOT0
fWjF8r0b4EB2GqzrHFZJ3aiP9axwVNwpIBQikHtd2YWD7lnpcCnK1OXF83P38A8x
xmwxxJmZbzmgwCTZ5uypG2lDAQ5/LfpFK3xE6eElyDsDrvfAwhlnbOWzd1j39SFl
uD+WFO1ksu0X4fmL0UlNuCVa9OxPbUDg2IUi4rOElXhJosyk32YidMfOD+0Ze7qn
sT132UovemIaTcC/XZ6kux1PRda+uYn6QVvA67eIoIslOipnctVnAyFeoQlAjJU3
vgaI3E5tdr/mFFGewYs9pXLatt0HMcxcZRu8WuYrI6tAIjxQj6dzO40O24jQgGqT
edhqWYlB7WR8/igS+9o/W/asqXzEJYHQBZ62pC9hRT6jn5OPazdlVfJujnTTrXZ+
+p8v+ivOBhinIQyPwlU0govwYgCU3uGw+7zCAzkIPHHcB+xi8G46n8xELCyQLIpR
Zr2hJTJTvXgMx3Jss2EVRiH5gjP7be3Z2du4I7E/JuzeXjA4NGvG4iuhws2Gd4YZ
ZWda+sugwmmqtb5eS7HJvLugr7HG5qBkVcZlrvE7C8faPAB1I5y6NiwBjSruXu7t
s0Xd1dUayKwfO/vwWX18bTqWHq8Pkz/CKXcy5utNX1ZP0aiudEfECwhtEo2mu0IS
usRK+kWvTcetL+X0YnttthC4NUtvGCvQfSqIXyOCqv7sFYIUDdk172irAEGBhmDD
gx+vN9p3aEQ9j2/RktgtneAQE1kSKaASrf2lyTG8LG3iRMHvp0pZxtIpzWkDGn7L
TMNFzn4QH73iEoPELstYwu/3md1Uqh/lT8i48cJDImo69QFDJZlxmwvKXkrhFmA+
WqPhZ1rVPWlwrbUx7YpVDtVqnZf3sbeW+Bvyf6/OQCVZzeP3eRn47xfArfBido5G
eSo8sFn80p2xTzVEUvenVMagmIj8o2AaxifRKtHYY3lWZOPUaU6KH9fH+SlDnhtq
9XPzCfb7wXUMS+KnBHzAu8sDdZcuMDDp4Vl4/07WfjRpuoPJkokjwrpnWCUWo2Kr
fFx0KfQfkBhx0vkoh9o8KxEyb8galeeAlE0xbp4V4xW/72K1gPC3SD8f9D7QhpBD
6ggAtj/EsqW5Vmidx0gaBArTx1Vg38YUOj94fHF9YCA3yrkjxE+fDHdwimtS/v1F
xlsYR0mAZQ0Tp/IWUMYqb+zFnN79rb9qsOAN40x2jO9mssTgo5og2MqNtRq5v1mt
a6HM8piuVCx+fGcGJRNEB7C1PxvBGqdqHJcSKlGA5YX8A1MCKqLpw2oKnx6noyIV
NmU6Ut2//1jVYVDsg4jli/Xufr+4h3krZFZF9rSdAeRLZR5faIHt2b0JsHgplOPF
UP/jskeb6pkVSiszOaeVom9c++ZNxFEeeIWZM46Q/AoCLbvAC1aLkok5vRTtw5Ca
eQdco7I70OMIp5kgm8ThgBCoAWZf/EHCPTHRPjOvbZgteWk8HZXZcWfwKhcb0GEf
Rj4cKxr++NeKGBnve/liXcYU/muXmTsUhGJ8yZDjFZI9rC7XlN29eFNiXWY3qO2D
eApJqPaVtKMKRV5nkbfN7TuobPUo3yS/JR3qUGxNLbNLlbMYOtDcidQ6I+zR3HDB
KPJnA0GnkLH57wepzSSiZWUYWV4npFoH41/eFl+MssFO2XRxMa65N1vyGdFMd3tx
1vsyHBKY4xzICl8adXx2+1dESQChw6inzP/h1exPaJ9pf6fotX9svy81EZZoTcw6
7juzzawHic2o76Bc36WSGVNsAGVKdyqanxLA+nSb0Z9GLeVUnXrFmCOJL7/MstZ9
57ZmYxevKLbzZVaQ6AIv+i3iDKtTyQVqPG6FN7xZ/eZHXShR00hJZH1SSVNFVJFm
LcoZQl+mW4o4VAmRFARwE/WlqZuAIvF8VsHEDufBkUFvzAU09XWeTLFgTL3pexgP
xmNGxCEj/3gtUr9KIgBsM/baInjpOeQOfsk3aBZaj64PIMvC4cbpdBSsY+xiNK5t
u6bLUGjU6tPMRYHRZn00d2XZ96mqynObAKAN93+fJwBDZnixFvhQdEm7NmuDWATR
J5EEQARPPSRTMVmelFoNmo9iM7uPLGWj+0aPuHoigEkDk8vLwqZcQ+YC3WAyIaqb
yFIJ8kPwtIkeHrpSiuDioILLrIGihdvsWH44KKOultD96vxU5VrFSuevk/E+D67y
Ymo4ovyOedOBvWXrO/l5kfKsl9Vzra/+ReRg1L4UBsdMJcpq3MF5iDPh9LyPXPkr
ObbBGZUHuxN3PFHabavlwar25WXXh5qfgxEWbefd9b+vc756W5Rk8EOOaYfPmvB+
p8uW7auohjQB0CKnnmAq5EfgSlVtcxberKv+pN54FIxYpxrcm+7sfrSKuYhziEc7
NOw1oQgWmxDERoKNHIiFmfBTYR4aJ5oE/ip8YKzuLTtKqFC1WsuEXzPs5EaTHGu2
rOqrjF+Vl7u7KZoHuP7GJab62bJ6ym/3dLlqA1mvmzUpP72yWA/gvB7U9+vSOb4p
4vahyK2rlfhTy4aiFBN9wYm//bDqu0XUUg9K5mdNd5V1IvLPtPeTHNg3MkmaPYW4
Yatjzro87wgskztOykhibWdco/h7TqUVnuoeZVkoWxSEdg1RXhXj+l29LUC/8ZWb
hj9x9dUUDa0zk3tpI0wRUTLm32JNG9TbaeT4D6S+XZ+iVTk3izcHOsxHv2ljaB3b
lJq9rOqWjJ7Urz7HfjEM0PP0aybE6kMspHE7/CMJgrjerFVHDB15j4ls8xqPh+dv
3zMnlXnOZjLP/1OtZNu7IbJG90znJolPFL/gLjbQsbmLbXcH2vwYtLtkS77pE/7t
LAwbiygmG15Oeo5jzDtfbTT0O5YnzqKXWb9zXPz9LoJlQYgKcXQozX+jHtaTspch
WbVfLrEo0pTIGMiyQlcivP97lx06oAljtGvSwi7BFnE7a8eFt+a8J9RGd6Eu7fz6
oxjUbE00e7faH2N34PqIhEL19+M/zG033KdpP0HyVxqFE8I59n6njKBF4jiAFUix
u0sA3ldwxvJSiCYqfekM5OmzKwArdr5jDHTRmtkRXg+1R/df3A8dU7nKcig1hado
6tjQKym0GcbHTD9cg6HcalpvlE5ttVTfypFSFsRIGOT99nQyremq6+zSKq8lLKtD
3enwiwsF03LwDZBftt4kzJ1SiUFp49Do8cRo40gPN5nokp6k5sUrfsmCcUTdQDsH
Ii89H3ZQ5hFTRvUO9jPaXXRdiwDzqbMbWQ/gBc0+hubYdqUShyi7u3HwMwU0qH6m
yVlefK8gCLMjjG3Srm1XHudLq+kt8T4O9MPBWRJQOrwG3fzd/MfbVIrEdFx8HEdu
xbnmY04j5IIw1ZQmCg0oWgo9few8RPLsh0+zDlVADQlQ+er52f7CnwIF3+YQQ5u4
S5YuCxSeK7jEvklMhVxmViNUDY7tbgif/wjGmNADRymKM/R2hPT1CF4LcmbgRiky
y7I04lyvYm33xX0rZzaK+4B9cYragNK27uTcoJvdWSBO4Hu92nMa0Q0ObEufgtJv
9/unQT/NmcDoiV9wjWllxfZ8SHJjgzvCEmZSLkpov/rr4GeiZjEZG1fHIjdW7V+4
u7db4aO2OUvUMByf+x2w9+bzRCb4aOKHCBewzVDGOyY+yvpBYPAiwZt7txrVaH5a
mUs85q5tTbbyPpw6LJw4BmUqyxj5VGAWIQHxaLUfOW91112KKGecQxv+Lhqs9Oje
grdCpnzkrVO1AMSYnLE0AGJvyhtMfN4ylPKO6EA4qenMTyyNzFlr3qdqpxjTtbdC
7zgVWUwcZoFuEJHm/OjcjqNzWDDhlNKQTGCD1kWaHtkjyrlyn0ePbZG8zD8hPCKF
urPOcWy4eLrT9nhJH1DG0qw+Xi0HDoeacWgjBFOaksp5u9mr7aokLLJPUQVRQdob
3LxWZ6YalhjFeiCPDTt53qcoOedshHiFo6QPuoLZj+aX8AvXf4GGQsYmUDZPaJId
ksC4yguWCTH5zSVk1ohs1APdHlBekhjhRhnBaPWGuwL/z2vuGkfpWZY52lkdgeG8
Zwlhzv0IsAFSMnmD8Tt04NieHvR0nJDsOp40HQ17AhIkoubz4s/fiZS6oEj48QMK
ItGhqCw9ko8dr3dVSoTLdUO4S/IheCuGbaw7mWfB6Truel4ZzQJEy1QQ+nIxrPd3
pxaMPCv3rvmduJtIddvsDyI2qdwFl/EPeQsS+z23zgLdf6A2qmhvJfPGdJT4nk9A
fJdBhbVW6jbjm4Y7JlG5pa5CftqZThpCSvxw0pJlfG7VOWlKG7oSoxxvRWEmxULh
AAMuSFqWeLwaMywkhOEtw8bKIHdwNTQTAyoB4SleyDKr2DJiSxLW44Pw8sknQGcK
n7somN//iMiAT40JrizSmHCGoo+A6v1NpduFTmlXc18tFLERyx16D9Vgf9K4FA8C
oWRwPlF8dgopkEED0PSLcmG0XmpfVfvGlsipdLJ3kLRRr8FRdffDzLcBlg+2kRxR
EY+eHW9qnPeIrWvzNhedV9GLQ6JjJDSIgRElHWrurh+UyzovTAj7AYMHP1cW0t0S
o5cPwCMSh6q/ItZpVpFMnfUVc6LfCIHaCsBVcmom6AobZQ0ZXjBoHUx8fQVZ6Yaw
cYYGm71VbtThUaTb81M4/Jyn9HN+085sClD5Fia9wnytWRv1DKSHLQLCm/klDadH
3dD7Ud6gmQJk7ZMk2479xVKJbEUw3x5Do7sB+T9byzpwM71xBtTk7XHteaWAHNPx
5RmyDVaWJxS3QOqWBOo9T1j4A+Sz6DGclbIULehR4FPQsTvSWCK4XC2fk/aZ5/ox
FWYMl1xJKmM2E8HnlukVAbc28Rf4DdjZRP3rU7ZVNzhiF36hJRMdqhApmOgnll70
Q0J4vxX6Zva+lEf1hNOzbrAwSc/bptDS1ou61f9L49MmPm4QNvpmYgCA+A0EH6kS
5HZoSPll/+ZpqCt1RKXjJqHSdS7HcJJ9lG2TakUw0RP8lRqb7rJuZv6rZzpdheJs
BQrs2k8Bjjsl5hXgamICXxl4R3EGatXXy1TmahA5RkhuEiOJEjtBYvSQvIbAnFR/
1M47Oz4xkVLvXf6hycJkfloMRPwM+lhQ0sclngPADkFPq71OupmCrSfjeiwsJFz9
+GEuZkM466TzHDOwIDrke0XBotxYjabSGKQKqRyjLY6WWKkhqdLzxHdnCBaUi4XJ
EAUScDiL9waXopYU6LEbD6jTfF3lV/PFGKpLx/UY5qz3d3fNPI73S+eAm57S0pAd
i9QHnBwFSABuQZsLtNsOxqKRvwiH3ZfXjrUrHgmQW8QoysREyJUCpLYpFh2RkrIc
2kakVvxjPd4yceXbVlPgmo94pFXIwKdsq+mgTx4ULMc0IB6X+DOVL1bdqw1/EuPx
oZ8kaLQKggM/WaKy0EYMy5bB3ceGX867HOu8oDgPFeCyFU1uqx2c3rivv6b60w8R
ZRotbX2zTR25wLIeY5O+d5WKjsPJfKXchQ4QOXOLMi8hVRbIUXxjsH5JBNONDas7
RrXgj2Xq6MJatBEUU9X51dwDzJtNqYcmUDQ/2kF3EvbFHGodfM4wsfJxtyGG+xJG
JzjUKCqSBpRc1BlVjv1B1mozPU6kpuL57uR9IiGqPWxLd3Ol+lQeSeuG50JDmOYG
QLveptd3u+1DBV8Nys0VGmgsRDP8LAgC1K6L/+XVIxYhDXETYx4Tbi7yoUvMvuDf
u0qUztax3bpEwYzHWHOvzpY3X9mTteDynAl+TP/L6oRAO+XgIBjQ/a0yKEAdCZiI
mxP6A8mM9HtCzU/kVCVTd9mdqiyKlXuyTa+Gyob5pmZN/0C/dzASkig2PUtEIpm7
B5UKOYRYSi0rfY9cidkd1/RrQlC9tRTTYuO1U6O2TqFVvNWNcLwZEQ3O3tMikzIo
2o0MOh3iGo5P5zB7katSbiXRZes6uIVe06yk4CPhla4wjXI07E4Euo5sHlIJKwM5
teE3WTG1uqHOgotqLjj4/lpSgEXy4syYE07iHA8+ATE49AK9aEs6otcdsB6mI2tQ
rCLZcQJVTTX3pk/nLIqkfBbZiY3+VMvxfJem1h5XNHq8kfk59qFAZGiwDw0zrx/w
KNgt06HO9LtUb0tVWt0jxVSmvgtCuI4fTCLaa20PsdfjFs08tWlIBsGHBpL5aVr+
S9knoap2JPyRAcJVW6z+LZSGriZDIqNXDH+E41tPK3hsz7m6lHj3CeSgRHEVWHvo
3Z2l+cSIGagXy+AhL+Z1iHWJFFGTgjruvveHaFvm6AVCLDrVzujAh7DE9/aW4Zi/
9DKPrGUC0f8n+KaLzfLl/cWKA2a36RgR4UnmMFUqSLDb1iNAStyluR+NWdL4cD/H
XASVtlGZesO6UpSvJeU8GNaz6fxla3ginUtdOFHrMzOnFDHOwyQ+rCUBPb6xJ/kJ
muzYXK7hqzNJSOCtSs7ZXW/qm5aRDRvgZlzC4eBAz6ve63yANaTC6c/F+coqBS87
bzX09ZjodfE/8ogARBKQqbQQyk7NIzX0zd1gKNDbIDnOOOqlLQUP3SqdqQMjLCXc
2KxqfnYLeJceP32xL52ifSUpDRFr425FSbovJA/YYS6P8iaBAmLB93aE/4YNcpqE
ZIlSHXmo3XM5Mo5J+4Az7EfPk3iqtZB1wWS4eljMRrDBUWLnGEaQ0fuGBQrwYksK
yIPP6n0RqI/IBAC475oPS/7S01gihyNIi9UzDf8flCs632LG8qyDbxM5ztF2nS1z
AOlMF8yQ6C7RKXuLHX8YIlXHbzZUF0YUfV3gUCsu4ls9T8R6BKrYEQkA82JU49ri
JkgdeM8TqRKrF+II1HKL5HuD4l7sxIiSfnYB2GvGn7JJcHjC2HWtJp6C7p7jP+6J
Cgcy95dkxxn7N34ovYJAXcPHJLVgruBjTNCujQJ6LyEwzr4/WpMXRwrmIKuS8boj
ESRMManm2H+Pp8POZUNWK2vsqX7BmU2J5QiFFW6YGb50nZELHt/JCgXPpZLJztGH
lqIZaM2D5JGvyUVVKlzW64Nz8TEcMNRhDgGf4M3HDNveKaJjyxYXXSODNcjSoAYF
dUQ2r1WLpiF43E2ihEobUsuR0YQW0jqmL+Ke2i69mhglqUX0njPB0ciGHSY8aPnO
fw4OjUZW+ow9TjtYDzdWrB/LyZTmMN9U56I4XuLDhan/zhtcoYQqlix8Pv1pjDYl
dShU7mnMjPYSj1QuwRPXd+256PUn9eOVrzK3J3Xq0SkDQ2GHV+wkRfXGBmJQYDQW
15a0O9weOhXEFXkyXHweEWmhop3a4Z+gEOcxesFbGm/YWebpRMDefTdoXHuusmVQ
TSn/kb13Gux7oCMUWs/l9v0FgVA2lOoP6Hw6K4+f+Mf5gcJTaSb88J/Ke1BsnGNj
P+Cd4T82FPQEFOwypGeb2IqKgEJpgl7LzLgIC2iSg9YL9MlmLZ9s3cQSmJh7tf2s
3R9O3qHGvnwWv7Fq1yzK3Q7Ya+ripntqHBIUBICHiQyhfjmOmU4zMDxe3KPcQmWD
YQXnYKuV7ddNdbiAd9mUmpvKNNAD7SlPusuBzR7ZdCBAEcVgzqwxYVs5LqMFyQjo
H3lttS6i9d1cQfINzavLEF/xaBIguS5vY0H1xCS3TD86KrG4fnv6/io7sOrmdovY
5vsXxZn8LsztgZqm2k6y+5Ze2jMM/bjH4gDjjvsINkBJBE4uTflKfxEzdC0CzTY1
oYkxym5vVVI+jLIW/zVtbnSen57pnNxsHkyXRXTfzVPhLF0v1rpbc3Uzf+1V6CYQ
dUS9UVsYQ6+IbN0JFmrn5lKYAjxOeJZe9+GBO4DfNiSVnWke26ism3m3i2Eq7b+p
+/sWamaH5N7yaJkmzBqguGjHe4grRAvu9d9O1MSKbfT5oHqcWRh05v275ngjE56u
qHrHoZXgIuiQjf7FHA/Cwu/WaLN1T9nXH9xxp/r/DeSwQVLIlVsRn60jRiSgTR3l
SewOFzXlNlE70LELXVTBR3CdZl5I3KVE49+KRp8RtjDviNuU8QcUTTmD1oMUgbgf
mpW42XMszxTa3BblX7nkskAwf9KFtGExjSWk+HOqn8ygsMV1ELO4f9mgQvR9208F
GJTfQ33fxl2633vzFcvnyZUIlE65JcnvUBWrRtxQoR5Vu1jRemq9rJJf0oXWKHbl
SXOl+xf0ANZGZmcUtDU8ymCj5qys1xGNZ0YWxQ0suPbiQrToNsc+CD0hFRQ2qCBq
pWpP+KTGVIRxgWY2TY16M28cCDWFi1tlIHDH5SKdQI8HlsO/gCTmrM3/KdU3zKvc
RLOMPmMycjEjEAJeSTSNqpFY3hgYKLx0GB7/B0YrvpChfLa60SoZabQR7aAotk9G
t45ZIbr/ewxxSzml0LXTHY6rgkWzAk6n4iuLVlCScMHqdEzCyJx7q6Pp8GFOe3Ef
jcJQnc7wU8aWH2UVkAzYh0ny/VlJ2SbjooXRD+1T+YhxGOuuAC1JOrISmxQ5le/c
zoJXxcRe7ZFX+85REOOactjwihpZA2ZfBmtNOPsa4Jr1cze2VmpIp5Xlp9RfpXNE
dzXInELW93lYx5+oS0SDI0OB7Hc3jvbPuid3uzEQExtiddTUgJR8NPPy/o6PCgQ9
G+5JgTmPINHUPWY7HrVeefQ28ErYz1xHzvpqCFqePxo7vGCA6JchWfzGu9Ed/9n7
cWz52SQtzyfRI+e19GYlREa5fiUDA2odMpYI/JJZ6g/nenww4+HjsnLcMcadwj7e
EgLcaCoZPIQj26kNFB/GYVDkrhiIPPaJmZC7siYitIHRlWGzKPLhNcyuTk8bgsgF
NoE3neQRBc7M02oUaMpJbTINAeR3HDvxSQ1dZgMA2qT4avZ/m/p+nVBsKeC2g/YV
TqKbVUESoBz60vYH1AiNM0PzA7LEIEl1AK0M0g3Jqg0haF2EeYgrUerqJnttywdd
DGoskUeIL2rSanqwBgNwYJGTzUEeiJYnoP6bgQza1PnS7xhMA/3pAEPj0hT+E1NX
1onctYXgN8phUnDWypWqcrbJ1pr+f6Fwnz81n5gUtp7M0oQZUPPHAx/vtnMt3ErL
GtGXJcMAeQKW/ZJHEJds1JgAo+SpeQ5LNRW1qpqr+LHuOblvyvQSqgJCU90rs566
wtsLZSclWChRNY36u81mqZDeWxVytrN9IvbuBH/+Oqw+pcwJMjMa2zFoKGeTwPJJ
cxQ8u9Gm6wca0lFRWJRsH1BGp4J2XJ7SZvb1yt96oBGc6Z5eFzCBaSz9dLvXwLwf
w/GtkJu4ua48zDcvYBdL70Y8wga1AlHh+3ZyZOM5CQj2EAxJCO7aiALJdBNhwU1a
qK+V319yfFVLBRM/8qBlHWQDCO/Yy5oGmcW+IFn6QZg82nsH9zvhQ6R/kFo13pGj
x0n/smpgmIiOXtEpIWq6kzP3e5HWDJNCm1XU5Mzsw9Ma9y9Dz2fRzgSxbQv5C7N8
h34jvvtn9YFDPWyfYa4vJgepWPCssxRTjal+ktm18TUsWP3reFP2Au7lFMAsFOA8
ng8w1tOoa31WOLPY/zCqHa6Lwa2q9WBnxFNWKJ5ML5r7EwTvq6d8aB/JByeJrW32
t87MlRn4FdqPGLUmNTdiVkT8jvLvY5Fhb/o9ZPEXJdIDc3JLd8R0jnnaZlI6PR3e
0ULiDK6hk51sbNQDn1K2vOoMIIY8gIMBBgrj9h3bjBVw0GHtuXux4wl+Ena45vw3
8g8t3ovKTcjGh9H7RLlEl14bDHSkYHKxF5BHs8IJeCCcgZPs94Dk+7OW3TdweOnP
Q5lt1mZznJYwe8kIlAJEwJrB8OUGJRXypK5gJlGU+GIL0PHYwqTMExsHIH/JPudq
SyVb3JmXVrS+fyf1vBOhNMzOUTrxfXFUDnCXu2+JxM+jbTaZhiL5UBkWCjum1T2K
f2W8H6RUvzE5HQrUOqPHF8ITNku8HjupNgME0SMW2c65TgZEKBXw3DLHuZdy+ex2
H8juUiYor4JARbu2PqMEWfDIEhBrhROJNQxKO/8gynl2txfS4qsIoDfEmkjHTj1y
B2Ty1Wl5yX1t6zDbx6FUqiUz27xDb6YXdq4+VhNA+Ck5CoD8Kdr+Dzh96DlOn+QL
EDrMeKN31UFplhmesfs7sX+4yxhtGw7kZqV7+/C/nKkokv4T/8c3BCWOjrLQnLZK
8LNEb7rO5tnGmXTLjB8yxOByP1CHimYMVkWZDUhTdtEfqnJYEiejpZEBmCcM+x3u
LpIR9KE4UYNEibbWMMC0T6Su3eJffhllvBkgcfncv5Keem1fX+YsXQfG5sU0dGWp
ZP5WvhHCdgKbWIub1sHk/01DBNSqsooGL9M6AZRg/IgUl6BtXKFAo/MxXOOC8KlC
GaWtLBmYqBJp13WUAJOgAIrgwOcKcx2bue1Z11N+wzjrM5d0vz0LK01//qT5TnoC
6+pOLZipSgCwMpczMqNYTfR5Z1wi3I13xVgZdhXYm/n30mAQE7S9MOEKhv4kVnhz
+wbyawBzsfFEH6A9Ohv/0HvJJ5Nch0D9QpAXs/Vbgjz9kNYWeiGDt9ErLwRc27Mg
H6MeEAef5h3xasuNg/bvCPY2k0SxBhuSpQbc21qtcmHutcdVeEq+7wtkwq4y2TuS
D7WX4Ce4EYR2SIDHY3QbnS+0V1zIzXAVokU9FRQ7ue1Y0iXJM5BSIOEMCjXwmF2z
xXWFi2IUPC0Y8SUdUZYQ2KH7Ip11pEufePJvRI0iTOPncZ0GfIl6nkr0FcbrM2oa
aWSglBDnkaR3SmbIKOni54hz/wsYXHxe+kWLb1BJuBT7pN57ZQvJj1nei8TsrBRJ
Fm/BNVqKqHRu7AHMswtF82lzvpYAjfi9Oh9OUP16lcWBJ/Bk5aJgt7/NHTQkFiQN
au/88LPlLj39DvF6Bb1y8rw6Hzs+MoNqgr8ZSbp8fA3cJ+BJF4ByAri1V7XhRsCz
dxBiXMHO+IgRZfTLl7EM2CtRaTnVGnNTP9J7UqmO1UQJjfQK37b/p+y8fATsd+T6
7PpU5PTiMttQYFjB0L3b5EW4jA85SPzmpa5+SWrogAeg1nrDEkXvXs0jEYF4MJIN
tcf1xSX6jDBxVcqCICMCll8gHd9n45xstYzhkg3KDgnrQO2FeUvXhA8xt3yQ+Qi7
D17qyCy7UNOdOjhuEg7iJkqAXhfA07V3SdfY657v7lVa7YyozVAb0z3FaOGv/aOc
OU3ST8cvhX+SLs1esFlbFVaZd6FC2jEGIrdQv+4JoJxNWYWYNNuUWLSZLisjJT1A
CRCdZoY2Oy3Hl3lObPcgdTUpy+RdmllR/s0AAxbBrNAkNvikH8EacBCrWwUhFJcG
yEXBAaLesRo74/HrxiHWFC4lmzG8jnwzymUd8jQrqyPs397fD7evVfb2/OWNqB+U
oSUHpYtV1YFGIpkTc8xeIF/JiVmrzMrsb1IC/Q46ayLOoPx64VrWzD0euf2jQLuk
jfp7aMYGxV436qoi2iuuE3cMdhb19QBkSoPoADrFSXNpfVh/9ThSZB53/s7bhqDs
NfOWjifgqfudklbX0MBPkIOTrrad/57fAG0t48S8XEHk0mo9dFlLAsMS/VVcZE4f
KVHigOscxRWeRUZlPhAJYcpjZIwKpKVTVyXxjdDN25YiS/nZrhuGoi00Pv5ysQL6
UtHui6sa4OqveOnb5+c3FbTSCMApdsY6o4akUrQ8Ec8x4z0r+sJDxrvL9hobpxZm
gLgm8bfaOikLJLCNTEwrlEt3EIYBWxQDTBMyrXYXcvnFfIlP23569ZDJXKrgdCf2
ufh91WFF7U99DpXJPSKKrVSYN3W0+DHLX21YW3//mG7ddPAF020WqIccJsEOecpd
mhgGVXuYEilsbtkHq3VvujwF1/ijxwW+cLvpXUahF35/wLXHwN2KSakCxL9P0IiW
Ni6J9xqGWtjUytPt/1w9WyW7Kn6hatVQFZwIHykx7jGV+XtIFJkSVGwBuuMRPDB+
sV1c7K7S3Dxa59BhphpUvXig+xaK1byKbYZ9BY8z+dxxs/BBOexHA87B+kSUZvH0
k/jtiToe4iVAUL1hHO+WKDXT4YvIEdT3cEAD0Wr3ltHZawKPM7QSQyiR4mPgLPt4
hXZ5lU59Pt6tnuLBSyD9ALSN8GTI9Tl93fghRYF9sL62W2lRvZDJi5LGniecwNBq
gKPDqFz07K6B+22b9Yh+9jICK01rScMdXKkCAI45bQTgPAuXd+v93Rakk9eb4Zyi
RDMaBg1GIiRbFtRMfFpttIMdgGCCAvVa3raF6TBHV9sZpCsbvvDt9U2bLYVwMG9X
v/+3EI1QRiHbVE5j1nzsovkBGvpVkjClhFm1ifJEj6dBgASs0FqK7Jfm65FgNt1I
mV9Ec3Qvh4RfUB99ST430aCHMRn2IdeeQ8+vsQAVq6suNkp+F4yo427nOzXIjar7
0ATNKQDXdpvSdpMqCO7/IBrh0p3Cb4GzEkVw2VXzlhfWuniwaBnJXxqgMKEygCgq
Wtw0tmiGTbZwqyMhvxse2bc5LmjGkaF+7b2bt3UWwSJygr41qJ5B7xySPCzCzZ3G
6SxZpGLeUnk45R4+QEWdmKMum36T0fDu2kLhQt67m3/TDl8yhGJRtXGjcnBs2oDy
tGR8rVkELO3MPFNqVw8SWEDQgfCjoGll7irAIPoqepRuPq0vC4zMvh0OUkHEdYBh
FP5RQlYV7LfOUwAvWbBNAiB9p5B+GRZVv6Etwq+tg9h3I+wyvKigN4aULfoxYI87
hcjWHrIs3Xg+qYTIfTuwfYMngDyEh5irOPCuWtIkO7k/lqOSafIYgQ1wUwk+a1kR
FSD19V4aP62SSm/SZ48rNURmTNi4oLLqQ5gW6b9QFdTI49ZGIyKCxrEGmjTbQH41
22l0FyGJ480Y5DNWt/8y/yVl+h1MMF0i+VbsGveW15TsmpUo7ANIopbJ1OZEYZla
PMGPq7uXcb8q1fPslB7fzKjr6b2gcG1dzHPFs0NLIsnsK8RYAuSUZG/iblMC+DiC
Ac8fsF82+3yc+/dMQfl+LVWiyfjcsMADBc1g4KFI5I5xb5ZirAYc8wuVAdARXtSS
sEXeWJrvHoh8V/0hNBY69QiELoEEDY1+2YLE5X+vqMCiChzD3p36WENmuKvDL1/P
kTb8sCyqp9uOnT5TLrlfYg6TaDNs9OpzVx18w8YfdpEjRAJuUmq/T1pyUgcMxYCm
6wA8/04G8nI37TgdoMv8YMneTW/KNm447/V4zysIi655RLemYM2SDfmTb1SXNwmC
LBsThgLywnOzthWYAivS8rxF+OvWmCYmiirLN8MKZ4Qj5QjjZXnAPOv4z8rv8GF6
GN/pbQus+ENCOnhBGzNPj0b/eTeQjzAG7KCVKNtdVO5kXYM09/u3zQXYiP4M+qF6
a1edVvo+/fDKd1r1wKo2DnTAs3eG9gKR+2SvpQ65sNiojA2YOJ+ACPQK/9uoj/wZ
vGOCKfQsztBg+S5XjFLQkc8NgG/i4PZYHkQ+ku1HGKrv2Ijb6HQiPFmtgRsNKp67
oODem/t/UzaqmwT3Ejzy61AKB2Kodhg2EUEAvQsJ1fFhytQdYu2nLgpKhGLv3q1N
gB34VYQ9WL2Do0VBdWYEhdn7s+xLzkSz7fstN0XAjJyV8nMvoVOeZsqxCTgLA/JZ
Z+DKXC6uxFvS18UlponBVGVfSc1MtSiMMvdxfTCa1cDbBMYJdYRLnGE0bI4I5yts
7zS8FWTA+Gj288WG2dpphNgstSwFDjiPhyY15174y2f3dxelvIxvZJrqdJqaDpqs
OGRVet4+kQJ5RnKo3b/0cO/FDF02fOIhV+Q3K5DN8yJHIR2ca9HZh8xNYXHfvhCy
xS8sXtA3QG9AdrXo4kWP/4fn3mv/c97WhbIODPKefADFnBEXLo/yC1QOcvA8tGgX
ys2KefBqlPW21xoLdJ63Dx0CNUBEAC1aZuqqv2D9W1imMvfn2qXkL6PuQmAsj+uM
XmyfmPYYjMx8UL+Tk32sYypPdWZE3N44kXkPkwJJRrYRTnEBvjwsVaMo9f+zXccX
6k1wiLCpFnPW0R20dH5qPE+lEuFW0GdDVatjSAHg2oQvU3vfah9mMVtl9DRBAs3P
u461AiEgRyLlC5kM/3haC+0P5sU+mNVYs9/Bv87T+DpcPbKINCAhoZfOfKVfo+TN
Z01gM7E2iWpCw3AdaWWxKjlrSohZi/qVrFxUWqsvgqtRIX1Ng4dAw3sTiAbTzuke
YuVwIjT3yC6Ga/WzYR9oXovQKAmtUxGNdnFonVJN2hph1GfB/+HVByZn4rF4cEKE
tNA37j+IghAJ/NieoBqHRQTUd1/CghTMrhfJfjYhvUFopbrIgQkTj8hXhY5fNG7w
wY6XxT969fFYy4f2vRdDl5+xYBpt2T8oVCQZp4tP/NsSizB+fvJWW3kFMQAMK2Un
SC5GXKVQnEKXjPZU4eCXBUq0z9XofjnezjAzaL92znggYUfrilOe16yf4Up4M93p
Q0SzAnzWkS8VfM4nHhlM9M4GBZ59RuVuRQhS+FkP2c1DFFI+dAag52hk9Sv1nLIv
l+KXkwz9Wnhl98o9j2pMnXnpDeVN0mSJ/HCAoqTwB2AD5ZRhWjozzzq+3cbBLLg1
ELO+F71PXLTv/MqBFONtUv8YpYuy2idGkAoh9wqm7MS2dJBVtzi4tmjmhW//fZlx
W4lC0XXi9wjkvIULJjWLc1deThvmHp/L1Q8ivwyzeLflDoHQzXOohVcPDntjceY4
ur303VO+fcRKytQ9UuQ9ViLWEzQcouJyoClc24HLODale/f60JZ6a6gATICAVosI
h6LGRbTJeX9I9PC22VDsscqU1kouu3UuhdHbB/EWQB0a/7gY/1Zdxk2XwgsdTPTT
bHXY7nqdDO0Q723PJS6mL0yhS3RQ8Bv0yVKtoLTDMXdYhvypWqIw2lBzfO+tUAS4
/B6f5QoNjYG1pi9EwxgPemKPIYeubAkJqW6tHuJWP2kVJu75G2ApDbGKeBjp2iKa
MhI/hiVK3QTgg9BhHjztuv6sLpaiuANNbgBz3e10sHa8Dra6lhQGCmD5Au+34xxa
d6uE/+vT1KsncMmR5YwaaM1f6jKnReGVjHBarZkCNWpev0BR44/FyJdmhiXbA+XE
lzrMPWU8rgX5edmKe3pXXxzRYDt88SloYPK5pIACJddOODlkd9k5APIxey3755uW
xhNk44UNR9ldavCFtaI7kh4xzEJ9dEq9KTBKzXG9bRvba60dzIaR+MoqSKCKUojY
OLO8+jgN2RCb1YVDymQchFLRXUiFrDXlA8KIyz3aKX6vuXGzQ9lrjutRL8xH1Y9v
vwCPv6/qRTe6OhQyBJVsjROw7g/0PHg1MP/8x43TJkiVRSdIOI2lSchGr7oo1iP5
MMPRSN4ocTeb42AVxhx71U1LuiiNI8dyDk4iteoI9hl1nP+eCOMNDi7s8US7G4C2
fDr9mOnU0k2v7LJRwKbnpUJ1kjrz1vytDlLiiYPc52+QXu+o3zd/n/0DWi3ANWbm
q442nfYFWpOhFGVi/mvPDkI9rc4ye5BXoXQGPS5Y2m0DoplbOn9XHVaa2dRHee6o
9DHrWjdKenh03lQ1PCMYehbCRAHjboHs/DtSCzlnCaKA2RsjlkjDVFZI7BsS0p5F
n0JjQ8Xzcj+F9PuOHNbUcG5qbCyl3RjoGE7sM27AUkEJDxixy3ZX/4DntCaUSaio
nqH21/uS/k+fTY9HVkSmC2Xh3QBYjm5c2kbTLQsA2SGIK5wSkMJGuB3MR9YnFcIv
HtKMBvItmPlyPEYvtFvIw1seyl1+ADeV0t1lPt8BeLhNz1xpGqLSJmD4jA7AVqsw
LttQHTK67bLtnDUQCS5l8aoHjE42oLS+EEkW9UiJJRc2inBDPfOEvX/xMhxTNkXf
UL8Xx7QcAslswZqkRMcgxRfBuOVkBx/uUmDb4hbfELCG8344CosQRWLsvq7rpq5A
yQp2RpD69HC8reVQ13ZA3gVMQD90Tb4t8uzQzOttXLvGqpTHEH14IQdoPJPMz3jv
S4M8s0BYxPPcO+g42cS/NiehxYmuVZp+P5jshvazFPuQ2Rd344BmHViOLQnMV9qP
VSq11e1xGnapBa8wH3X2q/puOyoU8/vz/xRgvKfwr/ISgJlbLVw/YxLAgN7v1DXn
vBUpEGNcuuE6cNRdg0pmCU97Gi4zKVz7eALm3e0DpysUuiJO0KjFn4zgLpYa3TLM
DYZ/rwaiU1Y+TP1kxkq8OfxPCX5EhGnBfy3kb+Qcol9FIqckNROKdloKLAxcGw4j
vQVGWaEZrW0jw8DKD4NE3X/XJ67xsZBmmleZ0TEXDlqiCfjoeqWl3UZuGgNdqEhm
ypuMSBfJleY1R2fr6FkWaCcHlvult762THZLivQ0b4B9HYWscznAk1vfIgmqLO2P
9FN1VKy1csscKQbGXrY1T4JNjXY9uZLNMNRb61INxYU7xQwqoqpo8yHHfqJQTOe1
VJlQM8sHKXUXWB+OhTpj6IkglusOexF+280kWodKbUlESfFn8jdllaLCTDtZG4MG
Ug4dN+3O6B0zbCUEsWaB/Qova7nbiIDRBRtk4R+v6NifLFUNUShhd9fF0dgGCDs1
2t3YyuzT80X3Nxm2Qy1pW1KXDP7GBmsUstVRMtEFa9BY9gSXg2zpW7OeBxgj8N0U
WKAcg9z/9lDssF7HxGFsXUNRW/mYtRWKXzgp+jLK5Lcjl0X9dUv0X7gyHQgOIqKQ
LBgGp6MM/fPuA8lXX4C9JA5DC0GvV3ZByErhTaFz8ASe2cMu/nN2FE1rUuZyHAbe
nlc0XDZRqMLMj0liV2/HVnXLraamrYxZjX4dVcBqTkHuF+snE178Al5159qpRqUf
twQiJ3kjaUzNCxj8xKfQ+M4BBaSYv1v3e2b9ovrGrvAonxn8vGDL0XesJPKV1SZg
eFujulVIP7vYlmvfrbCLHIEcrQ6r7rrvP2CcEQBlGuehWySpDgy1ZwnBEI2ZoQ+k
qw/yEX31f1M+PTGiG0hhpf7FQbXGbr/cGp7U/M8FlzwqugJRYY9KdHYnN7lE4MkQ
Ut1RI/EYFnK4yGR6gXsFx9Et8mlb9dzBNHe0Xqw6fVLRr/wEdecAaAqu/+lkAlks
2gDzOg+hEAHv7X6BLvNGpLNSMjy3qjOcMZMPuiRtcx55BV+QaDA1N97qCWJEu/dY
teb0vLtlAXVNM/S+yZ8Z+E1TkZIy7xHTMBCfjEQJBHF5G6O9IvPb1hGqixj7L+N/
UuzimeUbbUolNbvDAc4Xihnd+CguWdFy85eDZ5RAfFhXVRxUo5bKPbIinFvRgi7e
woaoym8/Q025lPlCICECYzZ4kCGatU/svNXUYiGj6Rp/axco9pt90yPJnttOnTcQ
igSmN0XctMO7gXgvEDdIb2vc7sIf8OKHv01z8oNz8KqO1ipwDeSFe84UmxrGi9a2
1bp3SN/qZ+P9ydr3Hh27xkDX+yAfYl/5mQlcS+8ErT9FiU+9KZ44hGwM22vjj8HX
OUWIyjNtwr11imn16krvJ0usnGfpWt/p8h1lkgVdUdWa00x2K3D/Q0oKqNVsQzLV
Kw8aAvinwXntW66YysrJahwfTepuqG8Pot9A0nml+KADSjn8DsvhPCUiliqdsDJV
ZiXKFTUemrke0uh/Xwoms/c4R3NzYoPiQ4Im0YZona8DByhfkJ5OKpzinFssNWBs
+47Uri+yTUvzVnuvxPzRtL9MAxUsisp+4RS2nD31z1fEfzyg4Z6cPI1g7x/O6Smm
eDNr1Olj+Um0qR+hWEVrECTlIEN1m02eNfTGzNYBFirUgYshGMoQmMHBs0tW9GXB
SKZuXU8unANHxV9nNwWehGKwZYowsr51DopIzs7jK7vaA48UM788ZNH/j0dLAX91
02aPSS+zsBGGEO/x+WCTW1L5nLJEmj6HOmpQ0gtui2RoH6+hKi1S8a5PJuHAqZXg
tknvQ1riQZbsqics5+ipP2laK0AjV8L944kPWsR4wnddQs5LNfNZ2aHG0zesz2NS
J6h7guYUUvSw8UmmVFq7b9smW66s1ciDhYYsRi+lbZpALczcXsClEPbeVYQeMsOg
nfAUCFULTUnKFK+qp/CTiJET2EDzzyAMMUZwhuO09xxjdNXarnTVM29aWop48vNj
GWgHFy91h8u3Ab0j0XbVjyITqBQj8JyWHUHLkMZXP6ZUCsL0/3LuEF+znOSFGmOD
DuPvaGDWi6EjE8mJJie2Fv6oghv4RlJGIXuZLLs8lY6Iq96oGTqWhCjcFeDJv6B6
ZdFNORlFfucZWkrj8hx9WZV4NMeL0wYc/3tAb9j9nMZa20MRbMWhRJS4ACyWf0/5
C7rbDBnOAgh7B7KRKX/G3p6O6I9qMK7DnqTwKmUWMH3bAw/trAEoOD3m9vrk5MNm
v0FeDfqL2AQpj0uaKAwv32z6YCkbvR/ehq12xBIXX61hii1cKivnW0Zaq9FkKE9z
qy/vyJPYt3EplWQAG5v5NgIv7UjLNlSf+kDi2Soh2CSNGCWIdQNeasiSW3sxf7la
GlcfcWxATZwCbyl+N/JTC9gC008m4TNWL5A6Nh2PyenLesV9iuqkFI+cj1XpcCqD
i0gUy3F/DNVuTawsBpqswXvMonsxRqBpCMu9ZGFG8qQBfnl+ATKBZqSmioySavRF
65O25RfUoeA5Fpwd9q+aMGSzd/aPe7JaK7YoTmyMNs+zqC9IgIb6ASJdZam6TEYy
UsSY2eT7Z3QJxoNb4ESt2n1TJdlSmGJ67Jr7oETJIHLCYjpbbBJLlISKr+97gria
k0Jzav5xPZD7PQA4HEW26YDwLJBwfoHmVRxE6rgSfAfVQPGi42gXBJmHi62hDjPy
PFQ9zLaRiEsXLCZfydGiqqDvKUHZmuZcpQpq9tW6NlVUHBBmNb3z4rZs1ppgZQ0N
znI6m//FGSk4aTWJaAKopgLqSOJ+dP0VNMKIAtW5NyebDpXStPxTKFh0jDOJ9kms
Y6vs7ZJZ6Uvz7hOL/z3bbSS8ECWoojS1Vzk0UJ2sMJWB2avY75//WXvx2qz2TDZo
BtU40u3pn446APraWLr34nDVTtaU7+Stogv2exx+kO6Ng92EzpdHf/8zoaXmGfkZ
LrSgA802VfSsmq2/8QWXPwfY4RlNrvp0KSaoDxifNJLQwxommz64CMo/UrnNmBs1
FQyKaLkKN7KKVYTd5N1iDoYnw0IpErkgMPACigUIgxHYZjSmZ8BvtHHU6wsZ9nfN
HKOFmnUSoFQx6QHnLOHH1eN/FFt7uZFeHfKLZz8laCB0PlHYeCkcmwuYnsypUvq8
f0rYGg/5BXqLwGRPvPQNswqi1fELN6TGT+ybtwxZ218LOiohN06S1Fcgs/ocyegF
HyGiEPgj/cwI+M4TC8zoXMqNWMLdefg3NerSd8KfH6NAEFQ5m1rfJjD2D8vm9gu5
Qq+tNvzuWgfwNS4x7Ii1eICTrbS4fBqUXPRVgq00miDyp8QajqAVFu5yrevCpbPv
sWy50uGxs2rCIyTLny8qmWrpt5BCdITEor+PkBS8VzgRzafuADS+gQuBlcRZfWl2
mf11BjdqUQxKwZvwJXkIZ9K4ILC48BOEooBD97Tp+CiGYCXdRhBVN7CJ57Nqd+tt
f41ozUaJcgm2ScM1XCA7ay+RAJYeCmkXQ1uJcOskQuQeZ67pID5FxrguR470v4pj
WJ4vIwEV4CZfouBEPxh01gFptYvF1+j5FTMVPiPXunpwnGsPIImcCtJa3V9MmHyp
qmR+XO9YteNAYYbaeQArq14sL7/cRdG1NNE7x6l2yATgDx9aUY8dN3YvUhh8ss8J
HNG6Yd6dRTcfJ69ZOFPqVFvyYCBAV8wAtcrNb44EQUwLOsFF1ASylHoeUI7+0H+B
40zp8Tr8h+yoz8iwZesYaf4LuWp2ZvzviYP5jWEO579zx8PJ2CiQCKftMJrQkF5L
2hq18vAOMmwispUF3zyJGMxTY5UvBrhWqSC1N4EbMdeNP6Az2YbPPvpqpyRF7Jc0
bxzA+RXKJBOeWYMvLhnquNbO3MPXYxa1wTK1AmCKOUMdncgdxQx3Q1Ar1igm6COt
hxgKo7kWk324UKxdlKAt3EZfIy9yanRRgFCO0T2W4NYZ1aK9FLsNNj0N794HhBrs
x9BOveOXb64M7doNtVLSp8tInmt1N8UkCwujZ5gJmnBIacq3csQQQf9CTDhrNczC
k8uNJ90SLhF3jlQVPeNIAUXmxIgktnLMGdo1sj7K1sfLyZSoYrw0mWDKybrOaC14
LgffFzoyV8TPyTwm9o2SygnwZ+zxe2J4lC88ZCm5L0UAueO922W67IG5G5zApFAH
X9Lsp0NBF5NTWreVCrS6XKXwuKu3UqWKc+k0YjALzxp5UiYKz1DaXn92aOHrKTYc
iphO4iI5Go1q4IwgZuI0yad32iamHsPRLW9HSTNVYMpvnxkfCSqdLyc7KB4+pjAS
/sDrc7QhXBYQSgftMQUyfavYUEBdux22ICfkM2IgLzwNOT4smvxH7SzzFescc6aW
1vbjiQ0xvolKaIW8mp2wIAQeuAJRM4CMllNrrihTQZ2KKmFlxC/IMjzLKlvUBRt3
aEkL9zhItw69MNGpbpHGdW0q2/7pJtl06aJgHyBFcf+9sE5S3LpvzJiBrpoljlIC
QZ0SmC6KpA4q5SZ4r3qZDfKa46I5xWEzo+2OUoKtFsSQgovkBXPa5Wbz5DwLOUag
oAX1C6qX7U6XlG7A6z6K2FQK7XlH6OaUBhV7CES3oe1/N61Pp0oK4xDr+ttcI9Lo
nhOagsrMbx7mfMIFugUIGXMK5b8/HBix8t5GhSjl6URmwjyh3/uLNfF/Xwq7sthx
hQwCnMJJHcxomN1qEq+t8ntXOQDJ04qvbUkgaNuZWti+c455KcVhnk3B4bYdVpl5
jEACoaQmcHAckti7UXAoW2KfpXt43JhRCe5Bt8Cy4XFnz9g0NbQSiusE0o0z+9OY
rO7mkmbnugQYDf56qGDUiGkHlcxSYXAzcatgXER0/c5Y9ZLi0wLm9bYWwiJyi6bV
yfjqa8MdWsgN5XyIPRUJmNon7x44LMMbWhFAs78VbxFWR4HO9ead0Z9d4UNJsS0c
wZBq/kSWf2XVDK1x97iOgX0wk/ThMMfPAW9MnY8kanqmBZvlYUAb32e1T5P3tXpY
9lLuUzFoCUvVplWpXAhfO4kMAbl2Q1VLdRilpDK3WIJOcMsPPBUJVZpDB/rNosuF
/3KrHKRiG7jcfWnxeoSKaJ5dF+4dX5DO+kKW8TTbeYO15eOPjW6fN14fxBSoogjy
E82FxXoLswdiAGGs79JqItMB+avX1peKDsmzdRu3FDp4hFk1Y0qq7JrQ9VcFNblc
o25fwYzOSMdSTZMYB6F+lhgQ1OFPUOzXswWZo0n4+229352td1/oICxnVmcwldIl
w0RPyBXY9StQeCG2uG5cpkVgGdZvFi0fX9qVBa1kHLIFC+rsf8gBwWrcY+5YKdTF
rvzcdB35ky12+6RNdjXjDoBIJ5a/DpmmB3M2Zavpl3ankjT2cHODEhSsOQeSDu1c
joyj1QUrkjhw2I79wUWVAc+/wDsj4295JbD4SXmoXOvZHTimkPnsxDxwNy8phfEy
q0ms8pjZjxBcBryuUxYkMhEQWKBpfzu4NSjkY9FhZnOnwRZEixyH2FjuaCCqNSAB
0t0nX84AkiZqeTzBtwSNbPkVtZFLC+qtkiEm/0T3op+TeJQxc2TBx9c+joUguUTI
BlkqiocAYNtHKMj/X1IjtGAFdp0EVNxHJIbTQQfaXvcsmmznBPtvATOsdM1mHchs
+xaCFNY9zcnG2fXuiF/SqeF7J54NtM8RCXBZ5m7aEbDLequgvCHSmRGZqwwiGsDM
+JQ4DRWdgm1n/Zf4EYTSmR/mi8Juy3XlGgNUcRUekkY/h3EYLiu/xXIpriyiLNK9
aggXk+FYlKye7lZBy4/JOKka+FTk1mnZksxjcredpdCxsA57D4v2KVM9AC0qTRVl
Y+wk2KCyLbKs/dcFMdz6g9tCREmYxDYiZI9WRPe5RAyt+eAEy2iRXvsA7Lwkb6C7
eON54Dw1NpX1FIlsvncyRXHgQYLIikdlF2xQEh44MjMjb/GhxhClA79+0dK3qMNK
VueoX7pPsSjb6xeF8ONbUq7gLP/iSZsDlPNcJMepIgCXPksDuMeRxFz5B5/AqJSc
oOJqOZ6ZF1w6Ti+QJUPQyAxP1cWq5cDKX5Dauv8PGRmilvek6Qyp05dLUH6mV5xE
6k3pjRBX16kqJ4kD0mk2MOpKXol3dXrtBXWm7RB2dhy8B9Bn7XsCMRar/nSd27jJ
6RW3z3hPycYoMUYHbKnOKYO5mzyEbmHBlEcZwMuLYmQjs1yFmLNmH3ceC6rFiaGR
zVF+aJhgDUsCw09ZbdRNbQ0lzmh862U5V5O86zUaEzUxQEsEQ8v1NqbVHyr7vEZr
wP7gjPLjTGlSAz8I9bDZOvnYOZc8nBHkkmL6DggEL/5T1bV1urDLwbf1I8SzxRaw
whHk8pDbxMwNJt8r/IfdjVlI/HKoCghdO73kIxOhuTfR+gcOFx66lHVE2hVQFPIm
tGYcrI/VCXiOfdCUX4iGKbfh0A7lpj3H9ZWATU3EOqYnX6UAJTqNDMFtjeDNtfKH
5jmbTYpvpkcd/UpH/75mnPJIrfhy9gYF4CibO7dZJv9dY3k+RKFxYFtb6aa2Zgqw
vJ4xJGDT6tAGJHbJ8kCGT9O+X9V9dwkZ8z4xo9v794hJCc50T6iy+E7Zz9NYCsAr
LlbUNyWdfvVzMsqyNYiXmSS1fsqH583t/JMVaMz8kobEyd4T2jZPxHUYAZ54syQS
ov3w5bjwUowwmBfrSa40aa1LiieV0zSPWwp0g7fDW1mQ4wGgQ4Fv8LGqxglZM/bR
jhiYAYkN9s5cfzrwRYhPAWueXuxQ+ZOjciq7OlYTrTJudozu4tKW5LmK+GDMaehm
5uq0IsIslmSlXoglmqXCBsIteAjGwt1UUExrRkaERPAROXvTwj2yWJmdMBD5+rMp
jceBtLP5WeFAvyDTln17E9oBiix5gJOmjY8AHqaoHWPc23wOGyrVUf2ldnpVGEre
pRi9Y519S5TD2wSGe7PilYP6IXcy+GqM8TgmT3Nq2CN3EptV8nDxdIwDRZDBQeMY
u9wARPzB65z9yW3zo+E2WS7LbXA/VaHBRy6fw5kuSOACbmXSH+etcjKBfeBZyR7M
vt3HhT686wkD7tRSfr3q5H/4RIDwbFJRU5nG3TbyXFrE5iCfwb/AqXO71OHBGlEz
0rIXjFlyxT6RXZ+40C0MyOVyFsdmYrBde5AMNODCv9lCLHhDT/hLcsQ5Mh2ilHTD
9yQZ9Rj9ZO2vbru+0faBUEIHn8brPkYzhhSmcIdf6me29vRd5GUUvjA+EERvsXz8
yOjABMb4Y9YB3V1eLBeCsN6xZMWmZb97zP/V+NlUdyekgXbEk5k9e37dZZ0JTm7Y
Ey5aKJfTr5zoW43PI0+Nnag/6Fip2E38FTIdwrYXG2+F4LetVg1iDyoFOUmWw0kL
bX0gT3ZhnQgKJxD4hnxIbovsiIi7BNacODgUx70SUOwCvTzV0Uw6xH88JuR5r/xO
SJ9/35X+lzwhTBTJbnc1c028QDRSCGbbMFuzInIUXlnigmF0GAYWXZgwSgYPutlx
Wcrsa3GlTofgrpFxRLH0kM1pXYX4QNgBe/Syms96BwTvHLWC057myaeRSDFh+ovv
hbfnfSXwroEBqn/PvQ+rjP9DSt1wqC50SwMRRa7BEtxbOIwmKgkq7WR9yVdRvaqP
yDkcGo0aoQLjBO+o/2T9FUfy30kFO2hktHS4HSV1noFnQQFLPySmocj/0I8aGS4C
oNfJtX5UEoJ+C4wo+mxyVQgOzJuBqm9uyS+OYz646hmh8pllyyc1kfXVkw6RldWy
7ieOoTk4aUo8SkSSXbJfEGYYQu4xZcSQb/P6l69u47i0FSuMXxRuMbCWmt9YZQ5D
Q68j4MU98Sqalmwt/kvlAwMLba+lJazynJtALONx6geiYnXoyitbgLhLdQgyeAXN
UEXLzHld8dmFl3bQ949gUbkXN2Dfs8N3OdacLY81LSAJRHl03t/NErlLVWDp30jw
KVaAYvsj+vZ6IpqyzkD3pTHZsmG7+MMevnKrkCydHWX3+hyBegBEEJnh/pA101qZ
mvujRZqVyf+x5SGQGavWxWMZ9xp+9tJJJWUqiqUZiS0GqzPgU+buoh2Qth9666n/
gnOXJZ7VCSFlaQoIr9LJYwBWreVh7pgr91WCyB18QKGjVCS4zSQta30w4XPENxNL
8LF67tkVBgHrEtKchKSh8XXt9fRUkWlIlI4miXtdvhypCB3KWH1LtlMKzYcYBUTB
J8vbm/VVWFM9RV5iJfkYRa9MjnGzciX3d5JoJ2csiebZrU70B9S1FJU36yGX7ns6
moTLmQ0YMet3pDlRJ6ouOLWgLKJixTxlHWB5EXfKXWZEFgu11C1di+8w6Kc2xzP8
ajkx5kPZEVIK25oXrQeZnKGyXB09DwvHZJTPqswVSzeGKHasxgd1DzB8rhUM7d/L
C1xKuc/uxU8Hq8/VpDr9Vyn2CYjsmledXmPzbK05tiW9oA6V+yVG8BInX8MGSVg7
2GnH4/5awBuGCgykz2/Xtc1dTIsR20jaXJMYNGK0/Sn0qA6YdonEtHbVOKyxlj8q
PkAWimNoab4SOE8l0dCXoqHUXP8v8LA6o5BHjb42TQtifQfCBoxD7nj6JfC63r8d
YMRf3hOV8LLOzdLh9Rt3O7l5ELZTJLC44UZTzaOCSWkWL8GbhZ2DMhZGprenxp+d
JgY0nThylwQMzsNPnldoNwDSbbE3cXv3HlvFcMjGXOIQQriNHhsrQyRmfTOUbDOO
G9i61bcL/Vz5aYmRPbCOy8aGWZQipEHXAsv/cHBCJmwtaD49ULitswbis6KQMJs0
vUS84ao/BcCnLLz8QmLFj/3VnhuAn/1PAJt2YNuvZFO7DzQ6vskkusHGuE1bdMqz
CB+UdDn3AxotM8V67tKcHi7D4HEgPe9hhDg6hwukU9nPwSLHD8NAicI6aZ7kn5Y7
4cpEPQneaiTgTpvF4cM2DsfAHK4oQdGZ7fx6PcwtUvUyao/gVsOdtOTviLprioHA
O39r3eQzGJ0K0dvMKp53E4ZPFWU3//3Peadq1XKaN+jdk93QVhq8f8usuv+wXNYN
iXo6NbLEDV2ciTV7cX+fS0osD+sS6XKvBaz/XHRy1Ph3iC8CXfWsN/z+ZM8AgbI0
LnogjtyYY748XJcNf6Igh9EMgGL9gh3k/7BatvwS0WJrdxYoFPMrksew+BN1ocLC
ZKCTIpR+iEVxubmTf3ET4v30GLKTPzZNJcVzmljBMUkc4NO1iG52ucG1QiKRJZZg
BbHsLUDHRJP9qqF5Tr0myT92GMaDXBJK40hUiVjkwxLl2lTT13et/GDvf0x1LMMR
WnLE4Zk62S0H6r1hfiMzQOYmDsywho+M1u0puVYv7N6R+GlZ0x/DMvamn3Pw97Kp
+YmUGRkg22SIfFfllKdq9yoWkZQDKmbjFKT+dBeY6LZsQQbpY5r6jTYgo+u9odfB
PBkm2NOB0lMKpB2RYfMPdOIuF4RXU9Eu3/qxTxt29ZI/f42jBWl9CBETlS+9t65M
UAyLgZ/E9k8HFiNBIzLp6p2ecpX/lHqo45GMHVoLR+uFNBv8fIK0c2KxIF1HH4nD
7K6fhookgXMNyKLqd6KxYQJ352FGFF7bz11kKPeAAuXdhTLk0sy+qaiK/1iw/OOY
7FUpQDo30E2xatUQJm/TcUVN6seG6O2FEWllz1ORheAetGVZDdQByalSHDhKbwQl
SGv4NU/AzmePRYM2n7PZbMIUfakMr8K73hBuISH2nc26B16LqiFPPcSjTaXxPALK
W1wy+8SsHd0asgojb+0FJARSRK3etyt2vY4bd7AFESXMZOQ7k/KyblVv561VxsYH
5huw6qViX3735TAkdIIKDmGP6iFiYhVOLFgqwd+HNLEgmHs/seBYg1NV0939ZhYd
d7aZm/WcD69TToqeifOoyFmtoUrEInfN/fktdyiUxLe3j6ldYfrlCBBJPhpsi0xv
uxaBT4cJ6/MFwd+DwnUnjGVYG2DEpkVemsWiKUESk16ldtEyG8Mwut2P8UsQ+ZiF
Pf4n3JqUgAwKNKE3dwehPGScraGlBhvSI4EW7aH4F78I5cHrhoLitOkuyapqn2RL
/8hkQPhFoPmAK934mwZ0evP7iFrL3ISqRCLu298OgyfUsK+HRA97OHPbUfL+TE9K
1kfMTG6kUk2Hi9t+0bV5XWomARecYwCLsYaJmgskqPZ2d9PYwpltQI8efzLaWDnl
t/Zyms3SQgJiJxHlbuPK8mg24sKMgDl4STeD6j6R4+XiFMyo4Ri0jHmY49asN1Gt
pGCJ52zOlN0zbVRiolccB2sPaba3G37d8WHkPDTHuacJd9PycHnv7rLZZ3dWmHX/
101Zdqq372NN/ovN0Ctx/orOb8+Q8cSjnqk6Qp4HQE8VNCXwFfCrvRQyri3GPXmW
czuazDzs80hoWrcPJ0ebFn07XwoTGRaD3FfpBrrHpLQsPyhrg+wuVF1iEpj1R4gL
I8vv+oqV+MwTUkA+V2Xd+rVeEflHGPIsqZWcUi1N0uCUe5o3Ui+tpJsRhDOIqP4x
M8RCb0WOsXHGDwe655ujLcIl7MOl8q3k6rQCTelXa8UxHuuyYPVvq7i8pQOyKvTI
SRaQvEBpzq/TWlxfPj4jGU++65EVcisMHy3LChOFXFjzHui4LXhQSoEVfkuA06Jn
1HUO0jtAhOUEQH+j79TpE6xNhV2aMp9hFrOn3LvCxJK/frkUPYxFlgO+xWCIXx7O
M1PbabhnkNxrSb+EIrZA3r9AHjiZ4d/x9/1IDuSiFCfb2nK0QMJAznTpwbdhq4qy
32r2ZfPbm8UaDG/pk/8NunPfRzHA7k1S45bQOqiUCs4mqyVgZuBry2wRKrmcOY+b
/cmKZp/Uscr7mfskc4gS7BVXKzFM5lz3zwn5IM9ML1gOxrYXYu2cAwHN6q2HyIWK
FebKtbMfYFgdXzElJ6CP3IUs6REULbQjLi9tqR++h0UPZoMhzwur5TFm18Izh+ff
E347MwXHKEWAEgGsw2Rgr6WrXL33cL3+vKY+Ew17DFZpMQHQkzv9jd6WlSE1J7Nb
LDm0mPDJcXdvTFGNiShjKzrnuzPdCUu+mcrMOYz6f3Nn2rA7dAmmwXlMAvLQpOtk
qCzzFJjXMDIRw77tmjOo6utKukEQGTZDr8+BmBxvDo8VEbIM3c6HsUK3t8Z/8fZl
pmzBuc3Q5HfvR+STVxl09c0vXVo1GHQwcXtU1KCT/eB/uxL1R4WPRoePHooHGF+k
Ga9vEvzYQIcBd6dFWOtVNhepxbkDp3S0SwPs3H0FDVRy0+Bjh7YYFb7peLGQ6/wi
Mxx67Bn1gpFrBkKoMo2rAQkrzbq6yTFIVvzlh+3Djls//ptP07rhOwO+CP2aFlmS
vKj0FHBNAmrL9njZZj7+76f4v9aIPovZv1vAx4QkercKzqDqWXyC0dih0UQUVfuT
ZD7IPJBeUW2HgfoDZef68qpxA1uJgORPcriQTivSbsfdhn4fu68d5qK+R0XgBqwA
9kwB/4pylRAjqbJA34CtTBlFs2j0XWohFsI+fzvpKBfWJR3Yvhnng1ZGjTF07qHm
Si8orJAXezJ0o/rfgAuOrH84xSmZgYFVB15Wu92/yHSadSfzYsNZWRzWX2lgn4Bf
QoUnb+ua0vOt3wvxs2pgJjIOxHQCq+ot+gk7UEy2LB8+ib1dTaQTsjI+QUo+rqcs
IasyHuD9ubDZMrsFevqQsk3xpHli5+g/m/V6Pixzn09SKXb2Hp86y4z3i4jMAvWK
RJXYCwQSvMxCx1cjpTH026KobKpeWaUPPDsJJDEELKsKLDXp8yJ+AIm4y2AJHD1h
wuhHvttIq8bVkooHbHXWRL975emfzw7OsMTF6kqz+pef1Eu7rI/mfXt6gpR1yVKv
exG2Ynbob5Q+pnIKVxdr0xm6uuZOraRjJdx3Z2TQnxgajpoWroJIYAF9kCEHB7qo
gODi3PSy+Gs6p3EL1ez7lpISk5tKODc+lK9AROFzxq4aVqbugs4n35bY6ktV1XRR
XWzj/NFj3frynyd6tUMpUHoTv+wV+zMSrixEHtiHbNzgrO9vZcqLaxCUCoUxaAiv
wM/QrwLq0COrF6ZjkKT5w7/sW/pq41Fx2vAQNP47MJZV1ip4eHwoMgOckVuyB3IN
MXgd1yoTYWYdAf1m/WUHTQhlYPW6Q8iRu4oeSmNZYejR5x9fyYzC/rk+OOuMaOyV
GQArPqxpUPLeTWxcKmz4ZMZW2qP5ea7JnCaEecmzFJSGKkZDq34KJQbTPxx1vq1a
O/s/qgSdErp32UtOfZj8pyGasajpzJXWCdjhMLNms3flrvQXMKCbRScRTN/3/sTR
dAqpEbMomC3csWV58NrTSTY9892rdR9kPnTAtW1U5q6GBiDg34345GO+s0raSCUl
E1g484nPyul1pXu4GtdciN95r5AtnOGPYS4NByg3pP977jbbhm3gHVaTqUDyuYdN
SeSFR/e/cUSqOTBN36s5efMQQJBrwF1jKY5cfslZ3W3U8I7z40/FIpbQ9r+YPOsc
0LXnZ6xzjtUDKL8eCgGZHZpvnnrM41Ydw3rBDS2n9K63QkIBuiFYcibXtSB4cRoN
fvxdBuRDzBELdwYAmmDy3jfStPb24s5VaqilU+TbqdEVfAyzyY3n8Qo0E7am5Gz0
Pue4957S5UIq/ahvGVt650F9SGQBq/I7RdM7BuVrZOEVjNIbO0I6qvjZv+zl6HQy
`pragma protect end_protected
