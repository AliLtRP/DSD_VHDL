// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:35:41 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
l2oLOK6pe+J1b7OjcDnzZbbZbVG4PEakcmMt0fSHF/0aSNBdT5tsixjBMVoSDTL6
VzxU0YFupu12whl6KXlThkO5RYltYgbmhO7MTe1yuQZDtTtiYtP6csZinIgAesAn
lPix1e9F8mVLIX+KC6SKYAqIpJVEYJM604+wteH82Es=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 7152)
QoXhw0xoO04a0xaA4lERrJUjCN3mVV1PnQ4Nlokks++LxWzaQ+5aVbR/vVCTUudH
zfqYNwwwuxO0ByoCP2w3Dl3T9oO987DvKcW4fw2E/xVlfno4Z/y1Fm64BmXJ5VnM
PvR0dRQEhlfMjZSVRp60QVt4oGKXOkyikzM9h6MfP9xGT01LGs/RHYBEtFiHLQ+k
BdsClrAzttmaXqhMW+G7h5LDGgrNaem5k0iyK55iE/BlPzZ7ciGUdhzXGAgnRpbR
DQT0G/E+BOgDjtKOG85YS+YcUSwzKzh/v35Nrm34PG7la0Lk1hP2LsdQW6CAxjS1
gG/M/fAmsepe9nYd7HJZNI72WCf808AZXAN6yfpWNp9raF1hqCcGhiRbuNHY4jJn
LIto2lxM2rBzHXNRm495ChbO2GN3yg1MO8cEqt8Wiq8mIYuOPnL7Gtu3lOFRYsKQ
zMlDPGGW6pgpmOdEb9MEOzZGYHfqwypDVFgN05dVBTjC+/wKwRas1+xoYZU9nwXZ
QCHFHk0Xqlevm+TUNO5NWh3wbh4CLxX/PNA2HcLYqFREk5RwZSZplhrQ4+mE+X8x
IBiIcoB0nXk1j65dgjji5x+GQOgdUuDu710avGqPORHvmkl90Dm3PBPh5xE/Kx8E
9EFRpLADTSJ3ryDjKU4IU48luOlsKyMIOc6C5KVne/DTz6Tcavv8eYx/jPcqKjAK
3A0rtMyV3SgM387lE4Stan8MXksgnG67C/mD5HsqqGhSODH6S7DNrXoJWoy//agv
8klGidh6TSZgWJ//xuMkKmRY2b2r1juoSn+DF6bmMpLMmiWAumsf1HCnDKcMSm64
3YWEl2boO1fQ2fMXHVfsG0n4BYPPKV5CFZUhnyCmQ4p+uHtjqtAN7tZ53oxCbHEy
9a1vI5UdC6/t4SZqE3jaIq10/fA5Frsszlmn0yzc+gBWWJscr+MVgWUs4O+TX0ei
WJpF//vTtqUQSOFKhoxFhnP3N8zY3qDqtM5k8IBGoSUo4OIUwSrQb3fRYQvPFUQL
gt3ihsUlqHAeh0chmxBxO0A7dlXwmzASmidE1OFK+NLpYgbCHT3PdVs/DHP1/Snj
gTHDC97gTPh0kVBB/kegEPK8v73bTjPcfC/kgiVP83csRgqvOAPFn42a78Xg9Wpt
jD0WosrjK4KT1QlPniokum1rTc8OfFM4Xb+x8y6RONqCBdVbIDKLKC1APaw+Y403
vhVyYzmvuSiLjKbidFyNfq3Zc3Rta+HDOCTeswhQruzRXDW8jWULoTyD/JlSY+vF
+5fpv0W8ihCY6FGISlWn9Kvj25niGDVbKpeW0g1YevKsyXQ5xzEwJBNLimh6DZq4
HUoxb5JHCoe/+BZVLQVDb5wWt98TwjMNIB+QgtekkmCGsOGDTXNkRi9mhXKweDqf
I+JJct3MUFrvvtsEx3BNqHGkcSYn0kWMiaWnrxy8OMDSquAR6l33KKzRdAVFYSVF
cIKdseMjx0zTGOt6T2zwwbe8BvY4+Is2YdR9wkoad4mbKZf4w2KJ14bVpRY7sC7+
0Bz6Y22MtJlo7FtqaL9KFGqpM/UY0jn1R45vostfDCBMg9OLgr3vg32r6VNRDCUl
i9Z1sO09OfZ8g0e/Zv4COJ//+QcdFfyEQSYlvURXk6IXnXMzn8WE8STLpNrAHX28
1OaTOayCEeiDgd0OqVGTfS+B1bM1bJR2YrNKUfFKteMdMlXZDJb3zAPlkCz8Gp1D
KUa6f1YcwmDXd5Bormb9jpg+bKwSiunlntoE8AKB1G4tnjwjbivKyq3Qr9SUyCZg
XXtez+YJEW+b5/XomXf7zemNim8yYd7iO408M9ABvt0dqCG4GFDyi+hvdo/6vnzA
H9ajc3330KEVv70S9fUmVeTvqsq11F7Um92LZmffmcQkA1PvFMe2ApBBDX4sdt1U
PYhcBMuP0pD9GjNC1Hw5//dlWK6ad4NN1uhig8Gmu8EZ4/Z0BWD8vx0Km4q9DaFN
Tzt4zOEYUtepBbA2GK/kdwbjOMgHSNIiR6h35nZgcPjt6vrB64o7v8RJZbCqnNyF
qbN4iyecscbjm6Ry50W0CvJNegteqUCBf+H8Nq9ngqyi1VyKr9J0+q9oUE7XRPeL
b5PzBoeZ7hLEw1a43Qu/AoxjUyGOA/w//B773jZ48BfTpqa76zMFGpVNPAToOth6
OMmfIeTs4gaaan/txFuc/0LEkjoDLLPhlI+7wdcYihTlWLKLHjSKofZjadLXro6s
GzwXowgKLK/Bcz7Frt6lEWMLHUKUYdlwhI4ae2ayiipKTzjY+jMN+2wN2/9Ba6ub
CejcnXvRLQ5UcgG0PKcx66QS/QEw/NjB/sKeeTPdg21ht//lbDfjyXaGLAOrk/7D
L9Hs3YAX9GpvfHOCa8wk1zYhAQKqz8UO/osRp3mqBMqFFMFyypDpnTd3T090JzxF
kAPYfNuYNDtkb2tCSb31jCZHk7xekaFqr37UL005/y02s3g9m9nynnNkYis4ASnm
BmL2iNn8gl8qsj3uzMDwn1S6rKdXBO3oJTSLMBTdOLpgISrLPAJvcxaPko16Ip6w
JwwoVF6FunSbiljuwo/wDjWil4NB66K5roDN3OdFng1+bhk6Om5p4YCZD/F3zIx3
tnBWeo2DT+ygIrHuQ2uhAx5w28cI4AIqF6AOVcNxbZyCXJaYVPBkGGOmg6ASZy6n
Q7/7US/tIlNw0g6F1zRrgsM0iFTAAG2DJfLY5hHUpTwgLArhdec3e3ycPq6rXmF8
uCh6wU9eVl0buiQN6WACMEhSeIE6ErRN4oqjV2em9+c1wuWL6eoSQf8EaZ2bcequ
kSix9cWG126Qg808Y//VWRjXHdZZV2iYqf+AiWR2Oya+wsy9EfUIuLf/fUzNyQfJ
hilJrvAmB1X+MwMjO/rFSNv31UAXrBtPTHXDMeSb0NobO4mhmZOySngAIj0MEjaR
DqvcRBrkQVob8AMMRemAeOvf9nBQ2xHODJaKV2EW1rosPHDnpuBmoul/qu7bOOW8
xKjoinajv61rTGlvfoihSh66taiooWcOtFJTMxdg9VUYYWbgjb5t92YczZETVps0
dltawC9zi6Sr7dZQmnOmbvZiXjora7/0Cb9rqetyC6fB4Bb5eSFwu/sBg5ILDWui
DsZJKqVjRrOXFzIN325SII8SO+L0tWz01FoAo6d+EpGU0Rh4W8UQnNkQp6Xnq0Bt
7YO4Weus4fcPXP8d7hcIBvIEApfxrAyRiGQKTqJpltxkeP50Q9Hmj27xNJpA43dN
CbN1Ow1hb4S7C8ZGN2ofS5MG9Q26SvFRCJGQhqEFU5WnRRFDpxW6zUuUh0tSkpRX
3Nat1PDsGmEbTyOqm48M60q1FGxuhWP3/G+ZD+FZm0CG0dlsQtOsgTUEYJVIN/Wl
TRuroHRkcLlKKuf5Vc8/m8Pu9swazDLjS3380TLJUx+6jNaIjxCmnNZnXFbs1HK7
jPw3H3wa5qbBU71x8dxATrP9zcx7K4JevTa/piqGHCZS1IRiniHoDoz8DpjFKa0t
rU/f2+E0ZLDo69oTZOfQls+NobDOXWrrHm2lU+AI6ySTq2sp5D107uKljVVIc6Tg
oQ8XJylMy62EKcNXmDUmui5zgygtJUDHwYPQ9nk/BsfC5LX4c2dDdNsY2qf1OBPX
1zq8/mx6506NILYBW322tnjvsTEHS+Vo0Zzi3ecdKDdcJtAo1oiHwPhihQxufKK2
zlwqIDNmr5jnI5YjBhHqC7Znp9XYAB7PhkTIzNe7KYeWGWW1G43eqinK9U1aHe1Y
7pWBY6JfTPg7Nqodqw2PQz4NaCrZkpI4/XXG/4HkIdqBvzz32IaHD0gGrdTMGyGz
7J2x3P2jRwI+EK8gEdgb4hi/K3Fz5eR/W8xS7YNMa9N8QDRcImC/gPZra8hwPZAQ
yVqbnMbL/PfTIZdomXQ6sOPlvQqLHLYxGGlQpbfngEtc42O1aOPj0m2HDexBt9Nn
IlckC7Mb0uRf7nmfq1iSLU5PH+L59XK/tAo38p55MhWN+vHbAAOp6nuX8WJyeozP
Le+hDBdCiAp9ZdoZ3YpqcRTaTk8RQjgg+/YOD072xB926lLZi+eeeJKSsOBTeUlL
YJTkvX4Y3T56P3xjz+d78sLZ0lwnSj3MfSzScy7JuRxKT4jSW5ElxvYu5ZxzCzQH
wNtTBgvXKPR5Zfs6KGY5Rr3BEkmO/9HFKAGA2S6PVp0MHdzyUgpBaTh0abkWKLlY
wID87QOYV+b8TbCV1+skgJSLLw9Xy3gy8sSnHAzlALbSexqBL4DhkzlDyK8vEEx+
KcoUmCLVJGvg6A0Csll9E+4FWeaPAnukfawKfelbkjEJaMvq1zc1WkVpnIaJ53uZ
VQiXFScJPlh6yDWlMQTgk/i487Bsa8rABR91YFRSJXzil2wUUl0KyTR/pXLCQ2Uq
691PZlciqmoaPS8Hzq57B3oKqHbOtj5Jnm69bER6N7epP5RSbO7ji6JN2g5ieKKM
NyHpqCQs9q+D1S0sjJHKiqDQKhmENR1gKTbh9DJOaeivgKbz94KrRLWMSbbQ6kC2
0THxFyADBpAG+Ehfqc5Blnz0bZdsgKwu9vfA6qLocLcFgPnXC11sPMiNbW8Sxy41
+WSBtW9XDmWkLBJl6ZkOImppOJJXxIlUlBOedQNVAZjpOFgh8yI2rhuB8SC/+VuJ
H15jx0RbKw4V6l47y6CrPZj3op+XD8A/qD66HCsFRIIHbWflwlnPrNilRNDZpB6u
ZPnUSUBEPePXxTcAZMfc8qLQZ1QlnfbVcY4+1lhedA82ibcwhVTB/Cwe+nMc3V/p
Atb8S4mNi+PF00v1cnKKIBOJDUimZqeiKR24CRVeN8wBNCpB6iumppZG8SLWikk6
Doj8CRpOHypGKRXnVQkMLdbP20Pgn66MYIOSnJJvUi+/IcbY86nBHTu0X+GtPEti
IBhy2k2D0GMrMglg8PDs4MGSJtRPdrSVr8YW7RBkXaKmnr5iyQ2fzfO2f50OSduP
IbwfIYmFD9YDirp/AqyZVaTq2XBp7CgOzzdnY0TCT0Y6lriTGabg3gO50WeucbMe
NIe10wqofHK3L5g9g3ZjMiGGJf4/rSbpBJghljo0uX1Ohps+05GQSB7rYONviltV
oq61l+VjhOgnJbLeaWH8OCWOhwAs+9s77fzgUEtiOAq+MxhEF9uAUTRRjaEatoEU
rN+qD+zAjPgQmRpw6tdSmJ85Hr+l5JGkyds9s8IQ+zgXmFgnOpl14ad9K7QWHW1r
orbrzi4CLuCm3RMJL1//Xl3acFDRP7AVjtuxLkq7dVkYsBlXHEYxinGstEL0J8iB
JbiTrBmBvu86Ez1aXwdb+r2ofRFXkEpBVFgyWDCC7voYx7ZPDqC7cd3zYv0//zOQ
jgMcTa8CwqlFgrHG9Dnv2A6oa7c217xYhiOws8F5JdEqh2KHO96DQKUx1coJittI
uJKQaNS8m8nrIkmL5cfhN6IhmYTMd8H5NLyoiJk0HL+Kq/YdjP+zdxDddAAf7Bpc
VESD7SLCmLxm2RSA5P+11p0Sptc+8sVjPWgWRC17ldgS8LxmsduHgqCuGpXzHjrm
tPFLtXx/4wtFvI8a+3ELexmQzPpiusIUUK9KqUGAWF6RxcAZ/vSixE6Kl08x3wmD
rEgcIRb8Jt3MYgTvu/QTi9Dgks7ZUcJvZE1tM0+WJw63zDJRwpoYtxlRL3EhQgNO
lY6VcMD0KszUoYr3LBFn2wRXw+EumsBWw57iFO307Px2E3hEIzhZYYU3Du3Q9nZ6
VPq/vrlqSKcGe1tInU4z0ZzqHvoKLnQlhZ25D4cAD2Y98P+Ar0xbgud8C4Obzgb5
+gHwVQyPnZNGGJjv/NYdiTpk9vKhzHXqaDw4vav+IcsiSCHgn4Cir4KPAJ+Qi12T
9mjl6NqJz9ZDd5teLY06kCqPaNsmNKwiUTB32r9LNf9jBPGHAWxjcEqjla9L+Gju
qfjaxyK4U5DkMVExXtkK+it8A7HkWPDtEth9Zgka0motTnRCNqv6th3SnQpwsKTN
EHOsU91SgTHLNkPHI5FPnK2dBQJ7Tts+SRpA57mQGR8CtHqCHj60IoRYnuljep/I
1Cf21SZYXmWGs9q1QJXybVwiDRPIYFNpWiJOqVCUhT4t/b2XgmFkxBYzNR143NLg
qy+ngzSMh+ATzv5V7wTr2/PEcW9gQVaLJO9IYIReu8wVXhRZ5dktd/hsv8KkgbsK
GNGu/aKqO3L78Zc4fuSk5zdxV+ZH7IyvcRkwQkvIxxVL4thBZEYxybXH/kSubx5y
i/0i3jedQbnim9ft5jVurITUd0AKYD48PVeEBtPmRXDnfAPALVc487r7Ex7tJxnl
U83ur7IyFSLse3SbHQ/EgglipHICJVBKfTSdg+4BFmj7U//1GtLy7/sGftjQyHKp
8sKeOjuou+IOjEvq2oXdQcEcZYHfI6pZvRCrJVLslFOkDMX8pKQdhN542+CIyRC6
Im4gyzUitskI6pTm4ZkrUc3qpcv2VNesgtxu6Yl+nhQ0NL7kbhoFuzw2jHwIuL1c
x8upUtqnk5NtR62tTSX4vtjdYsZNcVmPf01xtxNdjNMZfSQ6KJp6aqyl/+p3UF79
dZN6FHa80ACQyfYkcazC7OSa7SCPusP2/9nn73yCQVuKvMV+w4p17KXw1xv7Jy5y
Oq0gDRwGS5VZ5o2ubjFkzUVU3PHEY7LBWtJXxfhWSmEATqWwg9UTLQ2gbj/rizzV
a6b8uZ0z24aP9hwjvCAq3emmizF6QRTvFhzXLQPKD9Vfrc7lxX/lgQNOmf6IDZKN
GjEf7bGLPxbHVcjKY2NMhT3UbK+tPG11+Ug2NVQ5IiX28HpN7NHe+anx/f7uRo19
Zaa9IQMxSk0PYEr5iImWWfx64Gw+P/EbcXJreUalM458UMCpQoBNEcaE5FkacMKD
4YfuLHh37UBHW7XhZ/wEH+L0m0wnAkZlBYDdu9eg1/ngxnhinfjS7eNROSfg6FyO
MqH6l0hUkWKqJ2/wRU6W0P4P5ToFiu3LxYp97BXFwoUEZZmAvljJoxGqZpJEKPmy
wbv1vTdU3PnpLvPUnf5slg4d9Ad5zpC08oUWZ9jQycZIUyNI09TDg6SAWPzeqdDr
3Z4vC5P8dBL/+9LUcghS3yJGr6KAMqHNKrjtzQEwwnKtbFsNUf2KGvViCYljqMw/
IKdmiHkUeK6Isb/o8tb6wtaJ5NMDu8VD5ldk4pbmxkhKDYy0Yegb2i6l4RZ7sWPZ
45RX9Bn/VgbJmojq6bWfG3HA5p2iooQEpmjUvP98koTl97dVFMDaNG2ua3UK9yh9
0GlaFueiuc1jKxs8IJ8c4hr/kSoCB8pMkXyc8wxUQG8k6d2S+nfZV8dSH85vTbJx
kxVU/rxlyEu0oj8IQQae1Pdm3cQOI8FqNenmkLm1FANTxGEHs/P2hAD1fMpRFgBw
BXt/CAf7iNM4m4BiuzKH5am3pI1iwPw/1eOxlILdcwp13Mfg+j+UgqCsl7qMKIdi
40dCJmcNfkTC+zrlCJ30RIB9hW/c42YeM8kWDyMeJo74/tQ2lDzqV+aqy9qORcJ/
NLBGSOyB3URQenuf3YOvpUvRiMqjqU7SF0dGvzSlcsH4bl4tjzSe3pid4K79xUjc
I9HvnWUOH3AEKtF+LxY1Cqp9m5oEhPsU8q7U/ovWXt4tKEJ3JDdC3QdRvJgkjm/5
nMsRVSikb7H6FpLV/cfd0vhhAjpkyn7fctPc5fBjc2hnvrPvJwZh7r8O19d64iID
C3PKyosVAncXC4D/bJ2ORYljTLRxSmLSkY4pSZwlQKhE6F+aDcCK82F21MuwHOEt
ZnmHsSl3eOPb5FvPgzgLoj4lQtgTWb1AdoHU9QGcDYnw03Vvb1cbLHLIUNnUNvCU
79pKxOTjYnrpXFbKwKoY7xhGAjvojkf9V7fONkg+/64llGZeGl5zAr6iZe87EqHu
9lNJAJHxIrY+RXTTjy0Y9icvT4hw46HkcNFx89GaB/rOz2LY9lB6910pyYU1hV3Q
7C/wzYnu9rtjoLCgqK+jFx99NvW1qmjmYSplqX26VCbBfMMUwwevYbWNV7gyco3r
N9zg4jHE4CizwgEmkoYrHOdmR6ooIiLtmYy+ZvwQctPNpIznuwznH9rP3niZfOpT
gEGNr7F5JDz3pxjRIcQO0e6B+ApvHz4rk4/BkxhhbE4z/DndFxQlOGUypk/cvSep
xG/PxSpY0ZvqxeBr22Jg3aqmpDEnckx/avKk9BwqEtsxs28xUsq/OabDYUuUflOE
LGc6q5aH4RJLJJ9eKKET3xvcT2cRwul89rjx9zGVZaqKjpa+sI8/iR+L9NR5b5ff
eDciSHBaf2QblkZxrhccmUa64xdC8J34VuK3PWrOqoLe1PfXUwvu+eAs5zPCWjvV
31CuS4GgNkScYUu9a+J6cjgu/UL2A0PxUgQ4KZofDq7CiKeQ5DswuFeZ3uAt7/so
InFSfNYxJY8YCiLclU50tQif9Tl+8NLlpKGqRZ3AiDo0AcirvgPQCAT2hy6WqroY
di/i3Y3TU5Fou/sLSIuqcM6KvAeOz+z1C57lhbd/37YRvqb0d9gpgRIVATa41nsB
C1AphEfQt0xy3MDjfKb/G8ojXUPC9y4qavELuucy4p6yfILhwIgjpbuWVhPp1CnY
plo8PB+HGxebc7s/nykfLzHmdRMkH+rdcRzya46r3Z6LR77GckpgzSDw1S8M9nFx
Q7E6jRqrlBHCofU32Z+xZDd4+RziFZ56TbUQxC9h56zkRAJhTmbWICnJge/v+nH7
VkNUJHxxLubWbml5bmtv4LEs45mbULM7gSgXqlkOYglCwy+y/8hZt86SQ4Un4LkW
IsIJg4ZcCyr21tIkDQEoBrYlcS4ww80pFWMROnE3Gepny2SkGHo055UmUvuYQ9qb
HF6cCh/CGJqGInflnkSPofQBFh3EKO/H0cNZdbpS8Bx4nJg+BLIFg1RQIOBjZM9i
Q0OToX4suLEslZfIyRss0jhr8bfUr6CPFXrpdV0to+3OgPKfE/ZiZKa9TCbg4wbt
CWzYXEGuFBEsb3FMSLXAD8dSsGpzGMjAC/M/7qjbDQ4wUPMxQLN4AX089/KBpk9x
ixRwo3HJa0phOdE+wLXxbQmtRNYo0mDNLdr4aHmF+QBn7OEXiER+LTnfz55gboqK
yPTi00NKzNTm3iZ6vvechNAOdMjNHH7KUCH1N9xTG2/eIqe8UjzNxUWYFnYIieC3
Ico6xPgUvhuXXc6jE5bvocWsr48HY8zVViCoznK0msbrQtdwtfqud9/sBb8tZUS/
fHV2aQgqJQAvUSWZJvrVbsGxudlLhtaUi/fBWB1CbX7sUFGhggT93bFm/8zFSVKx
34qZUlzbLvJLpDpAwo+uOs7wOZ+3Mt3Ro5ncbdhiASwHVwxqSF7uNhR+JLhJWzDd
yede+A9s9oU5Pwv6G2nh4VR+Lbngm2aUYvbXg9hsotvtz15rVDUiTz1V/OQ7dUYl
yWS2HOCdA4qFy2c6tIX00UtwV38chnS3tPIpq5N+aRm4YjtZv6gQqUg1ihbSFhFY
`pragma protect end_protected
