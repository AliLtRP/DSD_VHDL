// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
BNaQ5f5+JpbcAwglbxu8fYplsNKe3aLAPh1x0M/Tbu0jMrTqTIkv1rsiY0n/qf+14Fux+KwTNa7D
a+xack1+c4FkMrtco0k8qui2bQtx/QsPxymj7xeR24MoKhsbp6dbuNyOzmXT/htB4Z1kuLeqT2ZA
BnlWPmw1YvEWey1ImhVj+a3Q2w5vuKF76FdmicXG5W1sQJdQZSzLEx+r8JLLowxledrKznUdDBOK
mo67pzneaMpc0TRIeWrRxK9xOqNTFykVKgpXw0I8SciNkwkkepv+mfzHcASDReNnJwr4ZyUdzGzL
dt/BWrzlA/4lWksHEgwuQAL+ztxlhLgb3Rdv/A==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
SWtgAIuRNcCEq6PigpTtvF7yAI5FOfzyQZ9LV7RDsE+HwMfytAdpZyrekwDlckScJFJdB7RttFek
h8SGFSM1q46suoX2qkwh714DDWV4EzXKcTWPuzFTVNYi5DFI5+WaA5ryObY1Mtf1ti5WR0s4yLp6
Bmec/8QNCNf/s+LOH+G2FVp9S01zyNPs94pDow/m/aHv2CsSX53WeAZkJsN9Aqslx8OC6uPc8oup
9vSgJ7a1w9enoopM1fmhz1jhzzZ1sQqCszd4crh7ZmxVEAkifD3+KxuGogWfpdj0TEdRNGvHXTjx
PYc95L6qKvGL7D4/xTtMVpIheWecx3U2R/ui4FUZV/M0u2xzZx1uS5vwrKAjJkVWn9rE+s5fuaZm
E0UbLI75iRGR7ykV58vdgpxe4x74eQt7IOsA+iyc3v4pq/0Vgh+VkntVyjKYDdJp4Egs6AL2WWsa
THM5Afaz73TJnmOCbPKnMMVbhvulMlCkRse2AA8LRr38BBnUbIJBVzDvkOlizzM64HW4AHi0Z4mS
7O7rw2+/CPbbMNtH00/L2vqTSGJPy0jtq0nlW2CSVr/Eot+gINSWdvbpiXiXqkiB8BxW27kh5+2+
WKiVELNCYLJhzE2K3/wPWtjvSgEGwTEOHbzi6u3EngsveLoH88ncA9XU2UzgtttcyCDfPmWfSoRq
n9TAEJGGVQtASPaSte1j8MnvDp4L9Nr01Mse+/oB/0VvfUK3Kv7WEe9Lm6wda8I3nu1yURxJZ/MI
Q0BBIx5WdX4XA/l3x7Su86jb6BBTJEZEV7oy1DI8jcRUowciCoY4jqbQ2qafjjLF/ZMhGwm4k+PN
xzYVvqq22Tw9IjTZ4oHEO24N1KxhhSwwFhJhxOsY14jRzQ/+CUz0TAXUH00zGvylC4HY+o8pEHkg
8iEV5YhI3LbeaqL7dgNpeIGKZn6Rok3NZycBcg/Q1aEnlDzNFagclsEyejpp+D5Wj9oyY8vxb3Qn
0IqRSl2/aOgsjRKkXXwRJcFexBtN+NZiE4vvcYWj5nUdTcDIAEvIv26yEWTyyzxDOpY3d6ytNBG1
527YDG4Aw1f2NBaHwl35iieV8A9tRmWE1Va5m4eUJzB0bPixcuUKPCtzAOu+aNZW8EwNMr2IfjOy
P0NIw3FgsuTlnlQiHYdSEf/lBREMlc9ECO2zMgc3g3trpcn8mYIoFIrhAeiqttfgyRpieO3QHgwR
CdttSkdKefCXwDdyrBpg2HF9KBnDe+MnWzj434kHkLhFNaV3uIeTBHFOO0g6hxnDa1tXZhiR+xJS
DLf6lviz/txrMYAvVhlquV6YRWUJZSeV1jNuPF8nCywfMjJlpr9q/kWmLWld0P6IJwXOzK0VD/pR
haM98FhdYOmANYUpo5osta7iSLJhIWdisPmXgZto537MVF4oRceO2GzJ1ydoNwGNMiHmkynfcH3n
wEjWbHJZov/847E/hzza1ZY5tyyE4oVQXVztbwl5P9OtZ27uBzS1iMeswssbC0vp4WMYsqyMVeN3
3wTsCd5F61WuQ8pQ60Lw5Nym+UjCfFgS/3SHtCANs7j0nkHcxUG9nZlOwTMJtqHVsAFZBCh/Zw+H
WVGVVFzgbf1KyPu+hlNCKtpSgiZpKb5+W1sPVQx7QM+1m74loTPg52n50BT7U7zd1+CT0GAKo/G7
eSKdBkKu3HanJbYc77vLlRnGB+6QdDtv8Vh79Scb6mF2p2aFdDTdcaY4eGO1i8u78b6LncVcdbH4
NsRj9yF8VLR8vfTbJs8vkre9yVihEIGIJCJsNUFQDZkRjjbbYEIAMso+pk0uVaj0hhsEmac8NP3E
D0uvF7CYDEhZxHWJeWGICOzc0Z7emm3E8s25gKpWQwJNIQRktLpJCqUtadlz7HhenehAZ9aj3c91
ztByKo75+zLp8gtK05CysIH36jrUv/pAkYWKagGwzdNPGi/BAJUkGhIda+wSsz9RQNR7SJcEvB8h
ZoiGfF63CMsP+cfBnuFxzXUsScRoA6h+dMApIJgpl8WLqsnscqXyApXGjrmVXP/dJWAbA6FMCciV
6fwPJcwQjgE8h2iWTLgSMljEdEGqGs1D+WdWbnrWGIuGPnv+atJ/CSn6GLeLWce20PRnu6PI1JZ1
UsiiS9jpyzn292Nie49uhP9YUra6RQbhR8Uz7tWWjS0nYE0a3X3PDxqwzwHkrguXBIRomD8mGCIg
0WV/G48DJ19dsy6WWPLBQdC0OGDD0whliC+u1mLS6Tfpg9b/mkM9oDQi5Azzg+1zGpfs+QW6lfsQ
bdU4fc7ZFGFmLglVNozYIaBG74MVkMLPicsNfzvisZE9lfnV0u3xtEFBu/CAhM/iM7n0QWGgZAQg
DOH7Kf6SvN0A8/NfwcHRKBuU2xL5Vgw/LHcq6jco5lPAORPcszOsBBGG5d1Uf2BeRbb+sY+qURN8
vDYdidTXiZuR1jjkg87/fjUE+8QX2IrMTXFmaMfz13QSEezgGcpAD+gLqz3pgfCPSAPcJszEgfyC
ygTTAOBrSaOH29iFvgu1BhyiK6layf7KEaB6gerw6uNj4HwWwi3ZguwGVyCahBdTONrVBzBgR7SS
RbPMAiTIdYkizAXeIR1RIUWP3wnmP926wLZBquZsei4xJoDv7jJ6G8gZoFha6XLjAXFoI0hltDbm
ikzuSJA7MCoV4UmXE2XzSqDEyqfZjXE0nUizUqgCZmdCn2YppaglD85BiTTS5hJXMnKJMDJzGbX1
PxqInlk+tcjkzw5Ez5S6gtJGM8znp8vdQNDqhzc6iSZi3EaDJl3mXBEszls5gsPyAdtWDU1J5f51
EPIcst1WRdpxzVKInVcafkefIGS2NjVTAbk/1EOAeo9DpNsdEQE/2QPkFKBxq8EJWLakII9A6TTC
qz5M/F+gyCjCKWiLVHsEn4A9PMZ3rw7qQt4hrqs5CGaVsqQVumGrwmDQmB3xhtbtylzvg38b7HYS
Cqhz4ixs1fBPzQPapVUyjNnQ8JE6OPNmtSKWKAAm/skJsZ5+gq7iGFR++2nypDHxWkGY1V3vEIwy
sW1tbC1lEGLUWGI6IkeHddcnNKUUH4IBx+7Ge5I994asIIbiMyKUgvZFmqQWJCajJKfDyG0ZkvPG
C9EmoP7gGqkiCmLFghSKLswiNH2r542W0Y/puiTJPN6ezkDR7if+hLpfkS6c1zjTSRJn+kWaSEyI
1Qss0rdbKV4lhwV4nzH/Hwt9k5bdwnyvuUzEEqNMPZKdqn62r8NUmGpe6q4Z9XtgkDzowEsGeSj+
BSzs8//usVHudhxn+MmZXGmucYEqBNTd0b3zp076DbDY5PWwjsn0ObhJgMQhI3J8aIVjZtVGB6Os
4Mlz3zvTQaIoze3KkqGJzbJ7K2F4ReQiuQumwjwtvkI5h3TfgZroaxz5powfppDKtaFIZ+Qu3U+q
QrHUeUNxFhuaMBp1pmjNGsNn30vlV3zihi+0w0+kGvPtVAXRE4KHRlES9tUTTKva174CQ872nmYU
yCH7XftDEGW34tMV6zKl1f6ZZc9xVDGa+vle4GmDNezAk4ErB9buxzQqbugEtWeC4FqX9Ub6owy7
p9Y0UbyZHadZZcUSB870lkDANpAm1i50vEF60BQKNEO1r1lvzwHk1eTAhzTSUsjEDHb7/mWt1Inl
z+6Nw1cS26Tpd0xq+rx9G+VpvS77C9HAxYsvP93qVYn6zJVU9U6MU33nJVkfvUWmVDCb7hXwUEgR
2qe1lCc6CFT1WaR2Jp/qSHO7w0JDDJREPEfftQNVuafTvGowc/oQOaHKP8LTjG0KZ5ZzdY3E0sIV
SECpVGr+C0E5jUCStAzZ59CxDO8OO5bPW9+bK+hvGRkWp914d2qbEsq9KRDEVRs4Y+vjRoBtCj4i
Jfa8KfK2n6oL3h+XIUyd3zoCven+7SFV17bMApY8KRV8jMXc/k2ItDxVCPWPal3G/s6zE4cHMl2I
6Oz8qKbukYQg3GVIv+9ab5AExVVmhpztV/nxSt69stHquPNK7dnsJscLW5nQlWcc15YxusUqF94e
uFHlCNKN74hiM31CFssUIxxFLY73WWkezPbBmLU1JcdCiJCnmCF0X+G9AvHbgRGfJ+ce9ZQp4jhM
qSRVbUZbwSRiUQ6D5NrJuJz+o8TqIgV6B6cmKVVFPOe7vcQG219MyM1TFBWB5I1R7wE96rt60rxG
skxq3xkoS2VTDzG0Pl0tyPwnsq5AE715m91xn+gYR1o/RjRDX7Bb1BQWGJ6EK3VZNBOIgc5eLuna
mZH2jznWVdJ4I1ylOpauGXBz2e5h6+WgudEjo/x1C3nbvMIG7hKFrEi2g1hJYldB4udCzvy1IlUO
z2MuZ2mv0Wo9fDMYGaXZee7Ae2pjb1n4XX/naWK/K17du4AraTdXSYV3cismCA7ZYrhpPkkc/xsL
W06xj3LkYJRR76pM4SyAlzYkbWFUxVoYxVxk2zEjwGpmOpakQYwbYVYnoysUqtEve1fQrpnsv+CF
HIcifbvWnS0T6kA5R4d9rrqbLJ1c+vA/12aQdz+4+/i4CvqP+Afpe/cRPdqwm5uuLta+F1BrMPvS
EPJhB8uTcWNFVtXX7ioYFAxaolnURQpDj9Hpr7dOMkyQ8jBQHPryBhIPi946udc1ZdE8UvqMoTyK
6JZypfHyJYvZnO3kVHlRge2zFKnrdmnLPtXbwAODmiiVWtYW6ISE4LzsL3ybkwa4fyVN9pQvKH0t
HbAm10ohZf/H95Wi4Ex4AijYrcvr+wmDhyMiODGLZ7s8GEUKsxE7XOLUyHujqDqcXlOcT8eSIAMY
fCHgR0Q2wzsdz7aMmRNqy8ebnCIiDLJGchi63dWc8kAGv3lKNaBN5KiMqP0m7g3OUwuFG1jgCegI
6Q0bR5AiGhCoryCfq0f2ZOPiV6lIZSDeLlwuAwlmIl8WQCtQGFNWITkLrx2JOkDJQ7c6pmOMXOKp
bnUUQ/pQWCGklnz27qlwR+eSjCa5ctER85De3XODw5XpZoHHwEwuMNlcxYKv6/QIigil3wTHEQqS
rSyyqKb/HESKCjt9h3xSiWaTBPZaRWroCBgPWWnj1UwwWvF0+H8nZzetZHc4amUPClZKrIJHpPsy
AEV1NtunR/vkVKAy9BtI4ctkZ2Zzt7UxS3Qrm01HlWjpkUW4uKft8Agwj08M4vz5cYJb7qP+NzsJ
Pd+wUBBEFnalgCUgRmwZ0ChtJrn1eMy99k2ozRgGPVV7FCNPMT6ZMdRYA9eqBT5f5ykiPaoGXud4
e1uh5S/rM6gctFM/JXlqLa+wUHS76BlHGGdnNk4qkV/62Pd70E5Ff6hawjeUQffkoiMuDpF+HwfJ
TMrS0JZ45BAA38QIbeADkHIqdnB5C6fPL9DYcJ6HA0sVfhUGj+KsglUxbdEJMb7PoxCOnq5n/oZi
zTBSCMglqciA4v305/WunIkJL4+uwCz3SQS7MrP7WrC/Xq4+7jWwC6v+sA4y+v846a1hgyPNvtoS
VclAzF8ddSZUe0SqLaZdtQpUeWrE0+uHd0ieaLJLYeOFOhmABn6O4rhyKYaL3Tow4Yu5xJw0lIfx
qiSTs1+ZHRRuwuTo1ifX38GCayi76A71gIePIRsQbdp2zygmmXTByPeHiSLYYL6NlWhTwNGSkG+Z
K5B74XGVjNyjgTC8ejtWHTC12FAi+5cU3NyPcDWbNIWKfgZHR2wibON2jElxxg0gL6YXRFXW9njB
BaXBZkoIHTItLykxmSAMovGDiOhI2YLbqx14g5zYXBosKgYCBZsFTJBD6idMnALCnNZ4eNR5eZ5N
SP7Kbe5Qtz7lLSONlfnZDCBdFQ2iGciaSDsiWc4GKsbnB+C44UcJimdIL5k7gkh8mJ7dGBsqCP1S
nFEpafouwdEJ++W69VhfkQWMXQ3HYp+Zi6MTf/HNEBc4Q7wsRm4Ebph7Ec+NszjZ1JyHo7pQnSV4
ZJ2SotSyHwa29OnNZymopDxtODuKWccTY4A6eLnPMsQSINWOVrcbv2joGJzYw5jFAhdpy5zqeJK1
G2XZ7Wa130ECJdlhRXmz000mSa4bqUn29WYgPMv61s2tQHNcEI0zfsNh/bGYWIMxNniwYowytXIJ
syhdlhBGlkm+detns7ttHIUpzbLIdW5JY8dLGRM8XPcSpdRrpUmGeAXH/sk07ch83vf3/ENfM6fu
KCSsiUjO1q7HA8/CsjMHltldUleVuezX9n1x403fzIpWwGjEIn/ME5I4PHnUNCv/mMXkt4q+89pl
SMnRbFASfjkmZ4I7CN29VBZX8zmpxE9rKeMUqoxNkeIu0pX8bAJvUVA0dwY01OK6x9WpNz1IzIoz
SBL0976+GIC95hjkr8QaBQ8Czjl6qwlZ2cyY/WQ6BEJoT+rn2LzuWvZGt4DpyFCJNH72fa785mRl
t2zjPq4fimAMwxMzvvMP0bjf3ClCsvdtKBuHwj2mbkNjxcRA56XZY/uYQmI5WRcDtfzUV3DFAEKY
F9DOIJgY6CpsMNAgzITt+qpm8iwNzWP7RVkpX9r5sQZWmPiZ1zk+RpyzCcKvkyjjhQ3JKUxCpzda
qyFP1+k/y5g3Uvkt4M2e97iPOH3y9+Vx61Ms9VPMegUCagyuwVO9pPpMlYUuStKvFj7SE1ioGoRU
GwVikA+8scETj1Q+hl5ESgmhu1V103dQII9UllY1ox9BpuS5PiGuZiu5kS/kM5AqUt15iVWB+loB
4iK+ic6716WPIJSBaKLqQS//jxBkJNCvxOnVvrZeAXixPp1S3luuwPg+kCviQxj0zSgUXfwNUC6z
GzVmnTfOjLQ9qBTniPGj/jfHUsnyJ1xvzr1lb3R3Lm+9knvAu1Vo4MI9n+t91Lf/Sx8jvwVq3KXE
0wLGYkXEDwkBxEw8R/ZRNC+klBL4vrgump/ybn6IMAdZuxQBGfBgJxdlhxVSjGRpMj4SDwAH2jWG
6jxa/K+kV2hmQskHgaSwkav5wg2Ge45QDVRveQ2Ox6eZ449vet23MKES81ALTNPinO8IDsY1PpFH
+o1LI3CiWiC430cd9UIoAGOcAyFoEgcLlFbKKO7WSAgQuuMbflsMwAQpes55/JBvdB+8PnmxpLoZ
Xw68XK3wYpq9FpEKclCEsiLJOlz4Q/IM3saNsWc3C+wVn1sfjuMQf2mJzp9orchO6BQKX6Ac6Ng5
rK1t3OZ6wzZzrgW5rRaXmRJ9/CmttQyXjONYfd3eKT2iagCzppAeHsqjykdRDrhm4zOhGZtn7vsJ
wIYvOhMdPe3QKVCQcnUOP16fS6yxl8SmOluoIp3mJ0k4pfn2I1FlDwyBMI2mtA/bfgZdRD77fJUB
Ea3crmYXMAoNtMoq1BWCSBQLHq/kz8ZoZk+4fZlVxJbcFp+34JIF6Iw+v55Brr20Rdd3UTCdWNzO
J8nZR969N/1kUrgbgMNVcE6Jp0q33sdjeD90FX1AeG+VNkp7gCl20TfiAz+sQkCzfz9xJHVF2dQc
uznrZ0eiGT2cwqC7I6tbcGYxENvkmSAoVgwaBIxYK9of0JJbInLVLlzNQBpIo2V01/TkXhRPuCsp
PKEhL5qI8JJVz8fDZPqnMVDzhgtkkRFlP+q1hr42LmugbOROiotdknkv+VZa3VVPMHulif8OJVwW
zIBtM+e6FOQo/C1Lz5MW+5bb5zfkMtPLOAY/9PPsSRrlon/QJ138ujoUbM7JNUNWYn64DoUoMEl3
wlS5LcNnd3H51SJnTAvuboUMzmIgglkAvV5FrKXODrC+k9hpWfjuoXXabEx9ZX6liXTKQ7er9lAf
7zqz4Y3ZFuu9fEwIA9QZmIIcwHCbIDjV60W4mjHKSXS5uBakYUE9VpgPLZIht3KDwzFMhRmb9DFM
8sGKf7ZtEQzRjbVTv0gNBmOjDTR7B/EPT9cOxZQJUSqLo3Cb0OBmuSolHrF09RrD0J+8lAfzc9hp
hEopwgiUjLZ010TbhWSJUS/OQov+SUTewFRipJm+1z5zKThAeESHHS0X6WRUKwoZOeUj4y5jOC4W
SJSWRai0zWGnOw2Sk2jLl8WXwbTQjNjBancEGWLcKClYyxTS7CEGmNXRTOQdQInTevEc6gXdQh0j
/MfriRI3bIuYWfVNQiRAPwmWPWxwp6NeeBte6gAVIMuvHch4NLvofwhEYSQQCz2650zyyM02MvS3
n5D7aD2fFfic0uVgafMzfnm1WYV26k5ZIAiKH8gKCSg282plzRk5UKgdBAHq2OhzRAGsrtiYYnfU
HOFde2YkcVcAzYGuOF8nQR6ZCbo=
`pragma protect end_protected
