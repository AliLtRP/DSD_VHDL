// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
sGuXpu0JVY5DeamLAx9hZzVo4+h2JgLEsr9GX+V8O3wnWbFglaRcM9On82czQX4MEaaW3K9NCvyQ
EXDC8A71a5Sb7Ia9Ky9vOPYUv3wCLKHurm8DbWpr4qTn+xIl0Qkz5zXk8TqA3P6EfljijIr7TNj1
RYHRGySw1nK6y9/U5eWOmCcrt7m6ZndPbhY9dE7RmiHoWeabkIuUjNZ+y++O+PSl7xATP3/HvYpV
QvpvDXCYBlIwUN8+u3qTkIRJPHiq/lfOTorzvdLUZvq5A8VHaaMHKzM8lVxwvRXH5rv2LSFW1NmB
L48CTlKCZm/bOkoMnEk4egdyQH2UHmbxAXttrQ==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
A6Kd0avHDTq9DWiJHR7siRh/k9A3Q+SBQ2p+lOj/3wDaSmwb4FauTWNA+0QQXh3ooK9qB1WoBnIX
3T5o/CtRfln1MHg2l48ISMOFy81n+pcTqc6d3DKBQRuFNzmWW2r0orQJc86SLoiwBM4OAVcfM4Nh
0gGf3rkN/FGv3yJd1MeHWWlG3KRVlCnct6RRWuTy/biqOsoaPY94IgLXVFQHebUOffp4OysLFYh1
/OpvOnz5W622xRu61zRl+WUxw0MDyGZmLfQgMgf50iCj95DArsLaob4mya/PThM5BhnFTd8SDaDP
JdV1cXK8NaxbJsnWYoMihpaNh3kOYzXp31phvriUgb0S7jMuTMkbeieV8TfsLA9lMr6TF4fKWPIa
XdLr/jWzusBCITfnnbydD19t7/MRKuFjNB9yCvqMh8Dypldb5IVkGYCH3/Pz+sv72UtQQi2NiODj
Nfjc1GrjZwoC4RczBegKcqyMhKhHocEkSr+fzbAl9G9GpwqrazMv6PdIEB8qUztw/lsEck+p+ISS
0C4QyqdmKpkGjdJQ1f3+WTlXAsStdaAhXeLAFV1VOeAvkgQc8GK35xkwkvkVMHjQGlYTVsysTiCG
F0n6ZdjZvGYHcYSRsC4Q8z1Q4pEhEu4ut8rTglZ9np2j1lQj9oX7rde4O/xD62dHKWLLKKl/f/mf
kTWUJQWLVeAEa6zvAYC5V7u4OVUdtqE7pPl8gLPDz/iy8BNDLsy4BP6oXQHj3R6xvw4u7aYUrrX7
f0yUJdrfE5j2OSXoQahfZ5Nqs+r/qWo40/DWmqyMzu2yxb/9wXwm1I5DAJNG0e2pd3yoeKqtgFZF
KB9WW3S1MLrdpdQMg1jrcYisCJwKMfsePuOzG02aCxmaKZtofDk64dwo8Dr57BQdeAbreheBE3/d
HkxK67hNUK2zUuzlAKTTnNw3gZVQWIW34tpL1w4rYX9ExLPxutmVCdq1mQhnNfIgeaCnUbtxSwYH
czVuPWUU+WPtCcimywgEZdmjJn11BNQssiRDiul9+lkLfhIGbUPiPoAdQdvbE53vsAKWnV8kgySo
zJdCasaxGYlblzvvsg06WbTL/raGU9UtV58uuUDua2oyJ4qC6uyJ0N/Ku4ofWptU5PHD3h3MtmzZ
7g5sw/QmDyZMZE152vJENsld9RB9NU6xPeDxJBC4KtJplrSA7AQ3/qyFdC17dS24t6Vy9gVcjpDA
2pCtXYZWIc0cu0noaOlQgtulFTH2U5ZEGJzC7Jr5czuIwRFt6IDftrp+tKKuSB9hB0k9WLH0Vfdj
hWZGC0jw2Jywi0Bp8tTN4I8zEs8nwmDrclicw8PNOSTRS5JQX66/xB9S6wrLdLhRzXq3ve+/ezQM
yhQmBsvH771DQ0RsOp5Q5qU9wGvMH4geiMWug8kphvylr0k2SiTBNhZRWkmCzCni3sGSTCU34P6P
4EXSsGN690NEZgUmH7cURi9kn50Fm6f4cv2Ew81s1ju+u6bsbSD3KO/7Kdg180rZNvjlOkPEgHI1
/xOFZY4TXvljVhKaZ/uOp5BQ8wG4D2Zk/GgGpjBFSZD6DIUczkTrxk70Ux4BNfSsb2DkFQTcLRym
kYhOb29D63srYQJN20Ozg17ICBt8rbxg/CUkA+bTm3a/ZcKPDiLdEotjsC7YUTZv7garWfZxjHAJ
kSjvSIqlaES+40LPCsOvYAAcpnhF9kcf9vWaXAy83gfWlBXmO2zYYKtT3THNtMeOmJM2uzUxLlpf
M2RHBz/0GHDZspNC+YaVdPsmQz6pdVbrR4qj2oh0gb4V+oHc9iDfAGK7M0VrrFapKjA+rylOMdjQ
CEvWm4AI0hla7AcoDCtgF7uft+RBnmc/V0HDcIAXkyflKVSzdv2RdN0zECVR9hSPJHQCbfzdasH2
Br4UMbGENs2BEdvvZuZSs8jieOCTkev5zd8QQHVPqsUlfjQ6Zf4gIR2htwUx8Hd/IxJAEryOfXYm
L5jR4sWLuS4Rex+rZO+5z1V7vqKDvZtLbfwDyZ6qXxn5qDnzwWIgXEEW5L02bkQGXx0rdhkh4tdf
0vWMBBjLav8WF3xhf8nwwTBGHBAR3REb7uWPEfHzuX0fYBt43+Dq4nalSWa3KgiSCVERzrsC6GMl
DMOuXRNM9HmmKQGTSq1lEfG3XWpkbCa76orFdIHuoXTHFMA8P9Rs9HF82Cj3+kiI/Ymp+6eeyX/R
k4wpuNatsiISg7bt8HxeMsYrJhAiZfSYaFgkGho9GcolfxjaRSN7iCpoYLm1nbpx+6LtTQjRyTFB
EoOTUEpYS857AEnGvvNNvLzeXIIMa96iavB0qkpoXsTAakLN62I17asRGKhDQRalPN14dkxd+sF4
NQtca8xiFiGPh9U6pecOcPDXr4RUTeZ+Liszl6Ql7wgmo2GQCBCr8haK/XD7g5F/26xRK5U/UBCY
d1ush8keEf71QPZ0kSokVlMiBADXvfflDWAmc8FFltc5GpIs9B0RsjMjsRVbWq4pGm8bdqH4Cskk
sNPia3/ixQPK4U1/MRJmNoEd5zpDGK4JbzhdkrrxYEtVpnfRcd2PL1JUZGpeCCiczaHRymgF1RMZ
/KDO5fxUFA05QmsRGAc7ilHrOsgoynfXtLpV9KNtvjgGf+LWuJ/mNrkLsuJSNV9j64kO5gqN40ax
UvddRD0xlhF0huNClVhAKICYyAFX+nosnn6wljL1QZjPbBwl3ntLPCbqBTO5QlGh4keMgtKWTRsi
MlFQue5bk8UivnRweQ6btcKRZ09AKRcn+L+TGVmPbfY9VGjzH5kO3ZhcYavEgMSLToTM0VB42/Fj
NUJW9O6ZPSxvwmonl30cUlmML0QU5huoAVDMBMdC9R+cJ6WfjX2MbkrhJgYnRa8pKCi1TkWCGrR1
wLafx5ahN+PbE0r966V1q3pPQgPUMbJgrJb8j/qI3nh0VZ/R2JdRdA4+hkgNyeca92H6pLYel4va
/w/3ygTphMl2/Qbz47gKCDaUNM/VVtywycj6evBjB6sGSfl63eNvxk9HnEXqLs95KneiK3V1fm5p
tIeAHMWdOWr9YUmzkAv+mKdV64vEBGUdk1IObIewK8laOaejOgUHR2ndb1lSx0b5mbfSUimWPZKQ
oVvphGCCuvvb+O2ppzBnPkz+G4uldxETKtWgut9oh/lyEEBQ95bRWbkQAaeDK7d9qn56n6X/xrl2
GdbtuVMRosWWxKLAXmn7TkOKclvEcUMkNfKdW2rT9AH6G+p9Vo+5RIILgZI1MU0qa1UjURl+Q5iO
ew6I7lN+q3OH2iMGKQhe1DmWi6kQtuLycwjBT+sye9wE2ECw0teab7LWHQWQD05VUA4EtLnIkLkv
Y/3uwzENMdD2hc70zsJTU5YQlgpWScji36Y0OH+fqfqb6w2uQYeuRu5tNB7OHXzHexJwMbJWiqZ8
jE94mLGqfgOUf3cbpXy/QAeAkVMXMJ0shRHD9HATzBk9P/pS3FSLcJd3gFiU02ejg77lANR0WfsC
k/SrKPvRGkDcYvN0LYRDNDGFJfl7RvPEAh4FknRJER1lVyHuWgqPrRD90dfXz+swogn8W+7qkw5b
lZYVuw8RURUjcD8waiP2yRC1vJib9f/kEF2erLbbuQWwf1Wr9y63/KafoMtw446BtYp/2lrCqdHu
3K3xD0/ahmoaPF0AdCXaVcqmTNQoReCw3+BdeWU/vPjOKutddtoHCi9Uj+x20CHZd8h8fM13PyHB
DLBpYCGP38sFqdlGoXzBBRopuSfRIlMmETjUoWUNGUWCgx8C9CMz5N4qlRjA6lDWkX5+WPdd9Oq0
DZv0UQjepCMZIinAsBABEswxIgRkMOilbrFEgkOLen5uL0vPchg9ZF/dnF7XJUisHR1CZ2QZLz13
AOad/H9Y9MATtOFw/SbpIid3kRGe4SXyRpA9UJ14B9R1PigZS6nxL4eYPYn6F6BPgEgE9/aCx1Z4
AWzTZkA+2Dbt3Uy6lk32GmwxVBpSMm1UMXNXnroPXhqlAAzcvTbG3Rf8ycDdk9l2AgHrCP04Zj5k
yRqx3KeFbm4QpKVHNeaBplsAS7rgzC8zgR6SZAk/s6z3lbQnLDokiiIBSadv7sabgxDd+0Gp5qLf
3IRmn8wDStvmOFGATpWccXVyu5nXOwngcsFQd7o667bTjSZTC+KMSGqX8rjSY6j/H3NfIciox7iH
zA4ziJD5f1V7o48VktJr9txK6OxcMh2FWLOINKjs/vciwzXIArQcuXOncrAPlr7KeGuwlhoUVIKG
K6oRbF4ITatWY0+N2vKsxJWzsCW96c8JmQEbJLgMn7zoyUdikUSraUl3O3+pXkWyh42SVX0TC/st
mBymHrmtOSR3mMEaXUkZJvizPoIuRpu7xhC0UJSYGPWcKeLoQ7gNLp7KOS8ovqOXE+0tojFH0/4U
qhZNQb/Uh8YReISvIhvGXMELoN7OBgh927l/c/SEkGeIDtrOyOwAW4eXK6oCvrpVVvROkM1n9EAd
ZfuvloUyruKipsTwc2NNE8nRhD60oJNv7XnSm3MaDnUgGk1SYDW2eDtbvS2jUirINy7nADlX6Y0X
lepPNGGrl+Gcs/LjXrgBUhtvmFJbCkSEunheWMzsswXpLJg4AFTDqeJpeUr7lY/Vr5mUoKfH4DjM
JM0NTrG52PYcMqIVzyCXUVDRWnyunwYzPH4toYxhI168IuJS7fGrmwqbcDppSPxNh5zdcPTmjix7
sZyxNA52QzZ+wPDAjBtTZ4YKKIOlheSUvz8pAlsfx1rk0g30DMK64lFRJu45qw1guMuvVmxMKJSA
/GVSerdhFZnozusOWXmJUdysMvgirruDGQysWG4KOAVaueglsuhhPu5Vl6VbDK7B7eJD6Ft0w9I0
QyhWQC9FqtpmrT+cVODPUPs6xmUFWZqdm7bUWe8AU/JK8eoLVRPLLcKU3kxqjVPFyzJZfHgHZUt7
vRZgtMFU1L8rwEXFfQkGsmyJoZYaWL+cQRe2ulCe+VHbajNT7PU+QqdJ6mYg/ctq5Fm5HK/GdA5j
HzC89W5TTTt2gtbbMHXgwXM+CT3vglyJ6tON9nNz5UJuwwX+qPlAYZYKLYN0NjRK1HHsVgpv/l+j
Ts49ScrNkRHh+9YMPZZ+2xHF/SHqEQ9JJ/+vY+ZFUFZM+cQ/E2ppDyOWBIr2HUFK6Z/0ZdeAX9gX
uA5aRr7crTbsDEOO6H5ERqHxgemW0EHZshXMqMtKjoJk1rrDfgKW0oxILkUag9fd6eJWRT2LHo7E
4Gf5Xb7HgYO854cxOJb4AEBXauxfXAmzc8QH5o6H6EL7JI/RXka3geK9AfgbN26oOLfXN967Tz7Y
f/FWMWh5E4G9g0TFHOeHa5IDui0uNDsp79M57fr4TA/9GBBtWA5T+A5kwV0rQ2LNPylmrkTf2ZNM
bkFOl7rOClmwBhMUdxVUI1zbvIJxgFmDkQjtmFQ3pjLLNcBk/hg+SwOi/LdSWLrc/QN+RkooZsIi
wbUgJ0/dOYxxD19TZwQEUCQTqpRvxwvqpPfbYmgOj5UAc3sxWcatadHUkDJpzhP+U9cHRLt+h0Ij
7ExJoj+ZWA6sxHqA67/XYHpBFkjRME9z/7x95WCWcfzo4dfQYHUriZWPGh6cxZyjMFlRPom0mt7R
ENPGp3StE/ozqtY2Q4O+4pOPHCCcUxnVvT6jdO8DIa96IGIlXiHn8AdMkQ0wJOr7uma/b5Z6s3Yk
Qk2NrNFUG11vzOdudUh4y0RI9lVItniZahW/ODTvUV7c+eiuUZSdy9EiajZEp+6WTwIoIoycIeH8
cxGxkGLKouG1OIGERaef9A775reKGFeRcTyiBG3esVHWw8BluNmL8xSlT6oEoYMCq6LwvOCi4dhP
Cg9nxu7iJkn99mQh+kb3I/VOd1FqE5Jvjj/VpfV8Fo27f2IgyurYOJK+JR9rNrybz3y6aRq4Ct2k
OIF3xzPl9cNTNodNDMrLY4fKZDNWjK7fniDTh4ii4LlqSgvQ4EX6ovWCE/p2vESN7mSe7594fDbz
2p6mCheBWqcTaOFcaoom8SIGFo5sGu+gBl2ylKu60ZNdjITcEeLfJiFJ41xohKO5PNFQeKIT8z1c
qhWLJkPIE7j2Mvk5j7aYc5qGeP5i0OxrYBhQmB0IvzbWjzY1j3AednnjonF69Ga9hV7uKwiFkZ+z
qhF0F1PgeLkzO9gqsHzZ3MWXIgbJNrt419gYtFfk2WcHn2MeNdlZ8ELbMbky+S2l0mard/viQhZf
nZmReYsA+QUDDNNfSwz9eLkagMCQlcqGLutt6GcpL1am2NpkpUQNqHfpyKww5NxMv6Wwjl0lag1K
oMwodOfzAhceJVaz1SE8RWxl88ndgqPBomToNtM8kMsfmewqivKSv1fC/ItNu2fowDtyhtS9jlVi
SUzM+qN4YjkhQ+rHlfk2kL3fdJFd59qjkbWw1vEEzEyI/t1tkya4i+4zBc+Hh1YzKdnGQFdp9oo0
ztydkqNoG7r6KLkCHLuZfbtYV1gFXrjjVSklAL0EP5noICihWoNqQUoFgIW89VhN6tTskU/aWELp
KxBNjdl46zt6KzacDKpYpK4OP4iWbUmUWsIKZ2E4D7YHI04jMmun4yO+AR93KLPNaZ6v27+jmRdk
/WpxwmArt78I2wlH/XbwcNz55b7W8jLGCmW2q/PArXnhHmedpnEHiWl+oZYWmVylVqIl1hXnVeRN
e6VLFM3zNiJQNq2JKLsu040NARosnzeTo2eXe69VYq/HlX4PuKEJryL0qYKHmN7TdCYz3P3LdjHh
iUFWXzg9W67cgGj8n6AkJuVam6VYy+YZp/dueucprWRt27SSA/nTQEJsCCVihz3i3Cf4vPV7lPzl
YKqGLdMZZXUhzdibYzAYd1GlBXLwfrdvY7/JVgkmAJTOSPPuXEers+868iOb+CQDlG44JEkhf7Ne
8YU7RsoOVWCMRGgmwwe9HEXYLyjEQEbupzYHYLDd/ckkWx91xTDOkwtOGVsch77IXUkx+GsYcVtv
tszKBQOappl+DiwuwvDToKWCXFcK0Q4BVIU2kphwKwv/1Hf7lT/iatHcbIgJcueKHjv6BCtwyIRh
2z/OPQiLw0LcygtsHV+VILpxPtksuJSO9TNVDA5M9vHVSZ/mJiCmyaX23oo7lK5njSYhULZm7TGG
FpINbx4GEtyWcmRi499z+056KczoSjsYj5uC1lwoBN27Voh++mOA+n+DFodQlKyEvLcd4EcpdAXB
7rP5hqzE+dhDyCL7w/F3ovzpwDaeKyBvieB59GPL1KGfNi8KX2o9anUwHAi7ZqtiDzWyAmLQaPIW
xiTWDEp3zv8HZ4RKbSkUGKSfpjGfIPsYovwLjJzaHzlleSMP96KzwaqAA8mpvDUe6MshFyFEpiIK
tHmVAmMorBYTnreQ9zR6/O1YaODAl8AkehgFq27dJHoe9E0MQ9LdkNUK8RjayHAS4N7Q4xlJgtha
Ia8Hr1XOq49JV0duAcAaoCeapuzjTE38nOLPySs2ItMJ9juhVo8qtaJ6qDx2P7p+6RxrzgHzfboI
5RL3ymRMyYb8P/Kk2nnHZekVRPEzqu2fbzcHKSkjWctvMPwsZ7D5Sc8Zl2lqk1TNcD7UcD+YS0r5
3KEH9clOU6YpmKKe3PzmmfFqXJRB2YZ4a/a1CalLY7xKBF+5r+ygErV1lVfnx+12goykRhy5hwSN
jkBzuXByCX2AfjVZYKQ2g70W5auKgWYTykck69AES9Kbg1QwqvaCN/x6hyQ7t77a3qFdQ4lqTC4T
/HWJwRQ5DRxoSjyjwYZHMz85STkzwjFFUuNlTyQFDJvlIliyntt1omt4Xno6BJY5863C3O0hjnsj
HQxABv61r67tmRgFekcJaEvrphoy6iRWIiuM18ZD1Ox56Gfa52Qr/11BL56JxRONrwXm8YmNLeCk
I6E+2ljBdT9T4BAO9t7FDh2Ya59xXbPaWtMtkIpjLkmCcuuC0ptFjDsqpIuN9kyJQEDFTU+aSp5j
YOf1aIXUs77ZuZvnsDQWxGXhywumwutkl6JlPmMlnSKS1HxwozPR/I7Dif1DUmMxoJAZ+zR7rVPj
08qx3EN1XEy6snJN8URWLRzhx5bVQC5g8vFgnMBT+ex6IPEJPT4QGGrWFMSEq5cNZoZ3ZYiKyS8g
0+b67a7cBpCd77pQBOlCS10GCoTPa/y2UqAgLIOdDKIGUR/8RrvCLs/9ofeYV2sjBzEY0CGzPMnm
/xWSjzXIVNCk8TSTYRBAH87GOE4Z5lC3EgHNdeuCqkE1wRkNFZUI9waKvUTFoFJt1tZ2m0qQZdZk
mAiVniqsrajbLfcWO+9wavBTvbz3zQnbw/mNLEPEbJRnwo+WasoGgbw9YzEHIUIRQXGD/IkzvEEK
HIGTXi588Tl4CWUebhiOLiNwFhUSZWkoIePpguXAdZK+Jkddy5z0kx6tXVXjUCUcW8qSk5jsx0Rw
vOWaJ6+cLecu
`pragma protect end_protected
