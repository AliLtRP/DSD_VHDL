// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:54 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
SV91bcVROswrl3/8Jf8EGP5sdSGfrCTYHqFE0v7+HwAJFqAy99rXuzUiqRDJYeyF
H9rijvF3hWpQz6TAj5VeHjcFygbYJteCh9qfMl1YmxD+YCsXpX0rLSZwduhdaMrM
35uPeNwe+MdhjftZl0/5zKvlanw/6k9YCJtS2RjL72M=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 4256)
BFQ6E7e9QvVJwcmL8C3B4ggEZaXRtA6P5fSbUpHfW4lm0Q0T7bhdgYNd99YEVWSe
T5Xm5AuFW5GP/f35hoCnLo5tdu3GSK80mBZmgQbnNQgR9uDdKu19ZCvrMAb/GAh3
xZxjXmqaB64SuIqVt0YZHXXrbvwFjrm/IWlyj7n0pjWN4Kj81NLGAOqWik1MhO7w
x1f2Epe8EkFJ2K1R8pThn9fQ4GxVCBfdGmX2EemruuL7NGQ25a1e63gnEwwZzj22
j7PvTA8dQVOWTOj7gwVvHf7Vc/JTeJjfbnSH9Ga5/4cGE5mMWh0hto8WqbVwQdxM
t3ffqYH9MUtuZAHlf8tZ2Pd5UTHejiSHxGLkXdrVB6sgPC/fJrKaJnIvaHxraBSj
sYQYHzpHiZVH0RljkCZpUvbNZUWR7v02xY/D7UB1ShPcOcs8BalmamU9/AIC41rD
tyj5K5xLyEITV6TvyrfKOIwOoY1Vw03LyMxnpe3MltFEepr8s/NvWexlwYEKRgoZ
mUcvX7HNi172KNss0DDLfuw/uG7TeFG+4RGXfZD24upM2lXg7A54H1ystiHAml0R
/vb+eOa2VReQ+exsl537F8P7Y5h05ZHVc8X8oHOhyaWIK4G3my0HSNek2fPndLz3
xkkYkoWkbTclXzeL2Sgie/8fyp17xieFwAIyG5864XxnveB00AwkE2Xpp2tcf0Qz
5/SQBqjO9oN/Xy9YKibhAfg0zMjZRs867fvQhXPBuNd0O+P+2lwgidMkHS3zMN2i
8Kkqo5faQAdSIwvzpjfr+hj+QbBi0hpRun0MLvEyFEC9AEjOSjL9XkG1gmC6Grl5
OR1Bjmc3cpitt4OgOImWU5RzA51ePeXU0kjtD0gwEr90hb+CuoTxrb6j0NEfP6Mi
VVkboGR9ZDmbfFRKpmyXu9pHkfcKCs2Zkr++5W9fmF3fpMy+nne3AdTT4DZFUwZ/
GS1mmRC6IB1xM6NiQnMyy8xG2PbMi7+7S+7+v8XGZGh1++kWI9fXtPMICNWpUuYR
ouVxd/ekaEdBNTi12hVIy6H+MdrW2ytwbWgOItpNhLDsj6zOz+WiQAEPszt8Oj32
p7iaNuR7eTeXb11ROjkpEAphAMhGWo8oMaodllm56/j2lwTmp3PYK4YQSBwlb1mh
Kqv+SnJ3fZS6hqp7/ig4KZ5BtMiKnPQ8bod5vAHGUmw9+ASWdehOAdt59jiFjZqJ
3XJZYRrlQipJAvQc2t6lzbSeEZBBtWOUAmqZHgWcuf26qu3a7mO+JGjkTBvmzL1p
4FnN4cIdX+XcxlUiUOT2nYa1Q9iVcZsGl0kygi8tGUVG5VsNlVNXpmwQOEGcts3L
/aXoGvbKi3+mIxC7kYG4q3AO8j2w0yzIpfExMtAheJhFqRtF2nOaVbCTaEdMcoyo
/8BIZsD0ayobVMCRZcEFEiMBWg4lcPJgT8nXUSSLKj4VeyKKPJ3E3xGFpIKSjFg1
dBTZVEmU1Ya/1+66QieB6K8Rt0DUOo6wqr/i7UGz5+82yOCRLkSwp4X7Em5Lsc5i
1yxk/wmDQ4B+5ZtrSBOlidycpbPNVx6UcXLoYSUCryltqjY9SEQfgPSPlp6IonX/
KRxe8bo4WiUUPGPJJ0MMM578rLeHKjjm8Y59XWJnHyIbVwG51nBRudjdt6S123gZ
9IHI0zxI18k/PtAxr3EkIcbDBjwQw4+cJzH3feZ4CfBJ1xtubt5+aAd/YxF6NE9Y
YvCqmuJsdClgFhSEoLw0Tzsui0EQswvun1avJ/DvqDhPCdivsI76C2pewV0cB1wy
YWwOemJxxLgVmLhn8Uv0wLUFIvpUL0cLaEqfZlq5OhwXeVj8UtcKT92O8+xVNS4f
1vLuCv/TO9VEEyo8wesKsRGZ9epiE31Kv86zAF0MpTUZAVWw/PtVM9xBKURd5ybL
2sstJJ91uSeNKQL4h53zXhcpVwtAQq8/EXF0SugCGf4wLxafDwH01mh3GioBV3Sa
OLCy4BHU5nbo83i4EbJoAYqJwgytFBUQpNZqE6G43C9WVYgJlpw7rSo67Dco04wf
3pWelxleC2W6gNscJ2mhQVNG5kDLf6icPhm59Qlh6GVthMtPcs2j8U2MGknTzMit
tq+uc6B2nvbpFN4PtrKng+s3TpskVNoQAiVL4VOf8mZ8dgvez9ufbes5Gb26bUer
LFac7Oo1YZTShRsOZOiOMYP0tBNbix/KQu692pl9XrMaCa0a+AiupJCxtgUMkOeS
cmk+gkD+QBO4p0+OY0vaX438WijkhPtMY8oVXYKKO5FdPJZ4gJa8JM4+O6fWiRpn
qQyY0FPsG5PJ7vagcQH0S5CmfpmoUYSlyCP/JQwqyixa7nzwEJoT+voWMSeFuUMI
1HnW8ROH2dd6GdCP2grCLobVjmqtJ0rAUe9LJgLp7msSGz+cSqLhIq0/TDSr+cHn
yAYk14YstCsxNaOhijA9n9TmysTt1FIZPoF7rT/PxgEhnkLpP4VxcKjk8Hpd8Swo
Inh5AW/zDVBdk84jwaU6/eTFEh8RoLc+NXMyGw7E4h5t7nAyL/yOmpKdDGnM8/XZ
W/8SLziVbJ5JWUXI2Avji2b7z915ynN7aV+e2AcSw96Tmwm4KaExbO5Zn1NjUm/S
LMQ/kVr48bdTOQm2TFsfFeliul6wxJevJjHNvPpoR1A/OggZvgzI6JAGXpvGA2fJ
oECoP701RGVu5mcDkHm7Fw973kPIb9oZyl4vC+ZoC9lw2FaNcw1n4S45fvQQAdbZ
CEl9/nFe222vY5mcWEUxUurlNrNKexySEzSbs5jXh6F4mWp92VB7cOYV23aeu3We
xCkUNGPs++3Q7Kc5KZGU7T4ar6gP1tf4ODDfAJt86bGHnrzoKOFLlCEqvH20pg4g
gZjg5+fmsN8XOF5NrERAFaXfUH9/CVHtshg2wt6UGOSTpERcZwcJy5r5qLD09umw
sWzK1HYoqxrojgsxKxKnxQ5Jo67sKbe63bntE9juYPziPGw2QquP9tcxrbmtXxzf
4671pn2RiWXw+4PRbLp02aZ7G+m9SSD6/XG8cuQhLFLARABHFFsd47hjg9a0jh9H
vcmfuZS/7tDJMifFlzfv6HS6XPGuJD3LOCdwF/ldQPP6OwQpxb1tjBRDXboqeL3n
Na24PlR0101EbFUWw2VHmzLBLHss47xxh671LcmxPdYZsS77JZaHeT4qaPRPFQak
XMQJbuix44u3lHX+1Cd02L6PQ5f/3Klm4OQwm8O6q9DG4Hbk2HbI83zsQ0SbkQjV
Ps8iDv/rE0PfoaW9Uj9qY0G/SQAY3TtIRbbPWAVyr76WBEZNhzX1NyNSTkcG5+q/
mR/KpkUb2tazK8b1XScZDMJcE8qgV6OqsmH3O0yAOcAwoIQNFmEwqlIjlGF5GLqm
OpjKPmiEAsaWuCNlOEYfwXsg+CNsyMQhaSxmBjtWVz8qUyFTbwniRivlbYfPzG5K
wHgDrkAWftUY//MU6PyUkYHsKzmBluEgEuYD3wr+6dZy9SvLha7tvscVx3UkeRx2
z7Bsk6ZdqAdm5GAo/LLoIPg0KCQY3WywnHUUjO7f6fUOU+kh4yFE0b+YN9MfJ2yG
mIUEx3bqi7b4GuEo25Nx1AQOEAmVLifPRIpBfzXmcN0IxgjoLPKE9EGyOK38hbSR
68wKE1q536feqAMvAP9/UeC93PbY5IJDieLBugen3v61wQE1wquQcY0qdppeAdKw
LeRVVFUJGxccA+P5AC+jMLr1HwFo+u1yM/RxP0mvWnmc6agULjwmISQBnXahKnAi
doeEna/fiepxgpBbCWhlhlWAxw63k26wL0KuctFoQoSIacBFzLeKrLFJlVh71rj4
p0kpsKuaeC2QTUo3co4zT4SDutNAu5IbVWWUJrnbaKNDcQr3vRepO0nSQZMLEtSQ
U90ST6I2Mwb5gg+VfFS+KLQWeVUa2zKMw7YgDY4LGpm96NV8dllST8vJxLp3vkgh
JX/DThEj0UMlZuVkMqa8QtPM/KaB0XKFbR/Z9LbcViwZLkv0WyhRNX7TUawZbv3h
CUYHlQBLQgpD2FORw4moweo+poeXD8huE15CTGTWEwDcsPI3FOpDzejr12+cISF6
DK6k9e5no4nnTxfuIgvlQuWs9ViDDz+cdLrlrh4SiiT3nSCZcnD6NpoQQDrwMQoO
CSy8tLiLGqlW6vk2yEtOLXozNI32vRM09Tk38U2tclfzK0SYicpF0sd23OOgzAny
p3ezIp6OQQo2dlCzhOCH7gR9UmRWwmty/ZyZ9xcM1FLZ0tfUD6iBzKM1H84DTpMs
DHmo0fBWtlFfFvwpw2oT0zmIjRG4ITOWIFc0jOjBtUedsofxKlqrHfvdhTBU+RSI
PJrbAC0v2y5ITnYWA51vyw5tK7ZqqZNMoNsWqxwyvT+0wqOyVlPgo62fD5HFAth7
9wE1QY23HWvN6um07vtMcp2OYPuitfy90t+O7G86mU+8F+jnV89EDrbdiCk3w7gl
vTjrQr+zbNbdwH8ysFqt80Zl0c5DaSz7EQP0FH+BIl/3+eIwBIXtGEoNxMKzloOh
08FL9/QUVuOK+GUaSHPhuTkP0KrQ/MLVHtTcosaKhEulehPPtQ5dhP4HiwYEmgyc
zQMNHVUWMJ5qhLmpUIp4MHtE7X6Gj5yGw7lYqDQhbh15/yE54iZK/IcYH34VPpsq
DL+GxeHdbF67RsGKOQ5k9zhJVhMOTS829DfSsRqIqD5aOC1nUXXgLwQ4pPKih1tj
AAc4myIJ2EkyDx23vord5ltuQEsh9TTKKIj+H4HMHYPoWbD5S3a7RKQ+2+G20EH4
tZs5SvXemM/bDRgm9HOuvIYXt/5q8w/P9DJ9yB8l1WZck/2fVLCHA34+CBsLec/Q
i3Y9IrTWbmqEOtwxyionnrlhzjBati+x6rUwrMaB//c1G9hh2Uzsr/FgJpIvW55B
9+dyzLwIERomCjiEMbkgefWbozsNO1qkxQVYX6t3TKhR/BFPmIbIKpLC0IdWJBte
lF8feuQDxnHblfCE5PZP8rM4VC84E0Rs9fIF7jpNw+E0sSBa/dwACKWtBqy7pvQB
FkkvASnll/ErYXHe4pywf1R4UDGKltZd7rgmz8Z6nmsfriJT+E99kXZ3zPqTdgkG
iMbABMsklWWmz0TDmbcdx8n4xo0noRW9h9nYpXvMGEYRmCndUS3Ov49Pg1ahbnsq
QlDGW+szPGG2qHrPWUs+fVsaCSVW4rkC3EOxEb5RgR6amO4P8EF6SJpoTWzZAV+S
vJRrqP5TiOuiN1uy98JIVFUvc8ffER+Frt8WdtOcEuQBdwcXfbxMySrlCV3rsu7E
7OzY80jxZv0Df2Jutk32aPmXE/PWvf//HZFYA5uyuqRPqqMxjiXxc6EVkjCWWib+
zZgltYn637kiVgclW8GSE7pN5bRJb8EH01wRhDmEgYE2pXAYxFoIobRUeWCGuK9e
6N8zXexX9j/UFmK8v+cwQIV1CRlvoFQ34Cmr9ZNbgqshsEXBTrnkLJJ3TcUuLRjW
7GFq8HqFkZOfbJfg93SVkLXuUnZF4csW8+CPuBMAGi7WiFfT55iM2utvnBBuvzUL
MvSxqA0lbZFGax5i6VYXFvkHXroy1HSK3fd7MAKlzTxlvuVf9Ae38MrbE/PLYATy
xbwGVX8EGSi+U65qihu3g508O6zONgZ5EGxVo3Lillk=
`pragma protect end_protected
