// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:39 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
NWW3kOpMzoxdkP25WCWHpoe3mSpuT35le5IhNqAsyuSj4aUfK7/0d3FTvdhOt93z
XZRbBtRsIPfq3y6p3ZjuaOxPCGCN9vbGGVTIQ94rCAsDv+o0r0rZQKwl/hY5jKCL
0pTI5ep5+TVCJU6M4XUKXeC2nySMis0V2CW0tJ4RW1c=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 8864)
mq7i7BRRId4xb/Z7a0Q58XZDT7jWXZb6hBM4Aw2ZdMndwS+5L7LpbAlzWJMNAfMB
XSKMZyaEzkrHF7DrHP1lgPU+GXOHGost4RX8UUAJixYhiacFRAqhGIsgxE3dmX+Q
Bt9K5IR+eAoWvVAa9uhmPXlVCue8Znz+FZgwoiVjN869ZDSGeDftBhWn2wmjaEZe
qAnBd3ZM0DmU7ql7p+rPLUHKksZcIuc+EvpNOW595uEr0BMZO70RqYPm8QLzpH3a
KfJy1Lt3x3qWuoo6IOh5VLVdFnhevcMdYVUFVuk5cMBtkquXQSqACjvc6te9ZyLt
zomdlEi7o53iWoJcchowNroU6jif5U7blJX2W9IZYTslmiwj/xKezzKQQEBbRZDB
5NXnK3h3s4PiDyjatODFEg2CZDOPd3aDvbGwwxDLwc0T1CDs+YU22yHqBwsZ9UMn
2y8UKVDPOYtQLjR5Vkk+9DNX4YXObeYZ36oVJCpH+EMZdwoCnyF63Ru62h7fd0AG
SQX+5AKcyY/ZT4vNyx/AdcUN3GbEtNmQ/LcoOlRClAnpqwqOCdVOj51qbRnfNvL+
15XTaiLo3gdsApdXEEzLAGqHK5VrHhMLXOEpX9vT79k0qQHGq6QpwrA6Fl9G0/5y
ogDLmqpMw8GoPWLty32twWtcuyoOhXtgE5l85py2MA0AeLo4AjlL6g/U7ZNo0grE
Eq5a2d9/8evSRMGomrouFygWmUfBPSD1UwOfHv1SCO3xncG/s4ZtiX13lF3Yn01g
TNMLJyH+8dXrlZHhlPVUMs2ax8uLsGYZq9ZJidl5jv9FK3m4twW27FjiAVmR59HK
Bxqwp5a9pBEEkyD0LL93SCl554nHy5LCZWUqEhdMRSUnjElbofAZ2qgAOyXlgipm
0COjYtw9G+7tCkjnAHF0EcH+lA4G9h3rtceDWpLZNkz4r5m0N2BMMgXNLH2Q4uN3
K4FgUl1XrhJ0drdtIn3DEYYnhM6W086Tc2Q5Hjuk+aBNauNpHmDF5oFzOvhlOnDG
hvAjI39EVZeLmFvkh0zdXA7LcJxqGvDrGqInqmsN7YYQR5eXrT1CuiZf9vvlkE8d
MHKiV72o65L+kMZqBfBEKRnlIk8tQq9HATa3YZ2Uh6qnTZdvgQ0mVK/uT1QZUO15
o6tKBk+ZCZxI8/XigLG3R1i4FQGQ3myZ2cIYw5lrKg0jT6pMFptg3zbL+3o0HT+I
JINJyI5mcVRiwiKR9TLtd9LOcGncIliPp/6Qcijs/tKKns2FJYzc5ujwpF/QhvyF
9rZKdqZKDmLUtCwSpqqjmEL+Vzy2SX053av4MMHYtpbvK5MUXJWkRuXaX6ldgCKz
DJ6+fV+80M6zmuFnL1kDdR0mJEudgysky/htItnHfuGZcIeo51ocrf9mTbh0IzXX
KCtcxgQHKwLSmF4eDerYD/1R/RwWQVg8FTXCCETlTwoMU5XU/VSMeXIWfwn9ZLeI
5pkh8+6cPsAxu8snpPpJ0GwaV7PQY8V4hk57jpUufpblBtModvkyNiFp8HJbvNT3
QKaqPgEOMEXj148CPF767UOkypo6NKvVV0nXXnGNXRMxD7qLOKg9s3RNXlHVZqTe
6l/V97iiK/WjB78ChvAG5nAA1TUjRCeGXID3V1lQzPhxyVp2Tz4eD0UvdFxMplyE
BlLghBH61DEZ66R/+A8dcOPYuSj4ohzqCM7TXDMqPKvPe73rtyWrcSl8bKAG/bCo
sZoZv9SMWcJnbYeMxrs608YKtqXOxqrdFpS46vFQj3pw9sZBD1Q4BjlBxAYA1HBx
hYf+5zxOeBq2mOXvhf/+bTlh/LSuyO9XR5V6pgbvdF2xHqUERgm9sD1fsSz6LXsM
QuIXaFrte4IuZ79+sQGrQPjZB9jhK8N1ufEbH3ULqmgyUjSVyIe+C/v9+avqXcR7
3KEQoUJ6zAGQFSnR1kP1xWc+/XrnZ6B+PhciBpb0BLM1S5EayesRTjVWfpd/v1Ca
ftkBZMthGAbO2QnIzTbGiuVneBaeK5BIGBns4wwvUdBJPVdPwa/Xu3KjN+QNmxu2
1gRoo1w6ppZw9h71gG+QGnyQT4cedNxxPez7JfkkjM1V8D9OdOpB9oojqaqFE76n
ZZlyFdn62ac6rGIT8ohyi/GRUvukZrH1awibJgYw7so30e8pIraTBjsLPlDhmMkq
6x8Oj4YdX8mZ1qK+5M1Q0loQlL2qyZwb0PU+NCxLyydJA+0HnLpBwIHiJGj1fn+k
b8Tc0nnn339YTwYS3h3COo3sknaQxjGdgwrj9XbDB3weLt0SrOp+7AVPlnvZOn6D
90NRyLeSucN+UFFx6P2Jc93GStMbh3JqYPXQ5sm2v5HxWmAdxQsmwf9xgYNp2H1o
5cFhz6rnw5KIHS9JXMz+oVHEPL6d/kj31Oc8Wtq8syyvnShr2LOnQDnRBLhoPAow
437PE5cI0wn/RKn47ThG5AkNibD/8G6V2BzT419YmbuRqNKghN+dCPBGwRpJkvJM
zsk/nZxGbmyQN6oGWWEdnu2RrQdR1Cm73eXdjrPNI+DmfDp4NEC8/MS/IAV8UElF
SUk4GPWz1n4j3B6jVfeYiUBAPMcTFmEx+De0GL+7h/BbLSg+DZxEaOad2qrupV+I
tzjx5YhyfvPT/rjPUPl0cb/MaSX5/FV5S3xkogS4CYVfK3WVJdfCYkjZle+c2ULu
6/r/NIjOe1x13KYdaRnsF4Zs4aH3wgyUR11hE1E8gYIvAnbrC4QyjWdMd3GCfQmi
L/1jlvDCqlmtdKlZ825Sk5w9NNsbECePkc1HaLZr9p/igalmbqn7VQkt5vqBULC2
ttIHYuGxwoVIUNZ9vXZgJ/dKIysQA0NlLb0nIJwcgLTPYh4oXikHmUz+KQI/3Svw
DZeK+b6AUTjhkHH8MwnjXrZgaUUUmAgDGZqRs/8g/WiWTbZ+CJivCFgN+xFoiPUL
CDhr4+iAjFZg2OEdyIBUTKRPg0hLId7YSVkY1TWJa5jb9aK3a2FDzGFFyOHiXQy4
5OGua2qDCJv8CAItyAHSwtcchzOzUoJJE9ees7hKRJwrBlKErL0oxlXkNyrBwKZC
zq8d0k082xAvTrYKDMt9iKxwN8bI3F0oV5Sjs0GXCNlWFMIJjz4VemxS8S7OWfTC
0JKX6UmDcb+WAt8lh+gkWoOiPFb5IhZmrt1lEDDmofbeapyHWS9fiK/d+EytPUqV
y0B1rQ67B/nzHwY6OD7rYjA2+6Yvof41Out2tnHI/ZmvoD3okRI6CgpTRVyOP7OX
dGjVArODYYp743RNjQjnyAY8lIYha7p4WZX1J3iJMHAK+OE5IeFlyyT1ISlr2kyc
yTrfQ5dtfgAFXJeBeg2i2pz5bVjqhh6ik4PyD59t7/bHcDBXiXi4GkG2F3onB5ds
5pUGf9IfXfe8s2pOP7I47ew/kae0ZfHK+XLNliyK9t94X8Ul9xSLaTuoiimokndJ
cUmg0qFCYob5hhmUIpML1iMYW4QjRsMee1VOGMkUIOzU8VeNd0w8OxYq4aPfSspe
n4JR4ei/795OiqPFbHirChGi+tenJWsBOWFJCEka88KsvMjdGpot1xAGSCfq8Mo+
qk+e6LaF5ji4ieKd/Oa0ADEG6zG+/UPSpQMdI8q/AfrUdbiJJCE2vx+/XyrU/76B
0pOxeOtOKOLORYYiHh32zLcP5JmSVbkQRqyvbZnP09j1KUJz07RyYmnrxF6BboE3
FE+ArYM1IpFdr0PSK0Vc2rnkF+nod0Pu9rp3d/SIRqRZjdmHuWgoLrA9MKkJyC9n
rQ9tdCCUl8K2CrZkZzhHXf1C9troFB0NUFU946X6uw7ufW0H4hDDY3F8i9pMaQ0a
YgjXab2Zn4Rlon3XDwY/0e5OEVclRFPOsEDYtWTmZ243PrwDew3TzDEovuD2XN3F
AKmzZ3gRkBtOBLPuPPEGYrNzR7LEqewiIySPx3kMByKJ2+gb2TMinl+oRV6WjwSA
NWor4wpjmxyrY9meUUrwJzGeXON2Iob5NWjzxEihXYELcJZNH6hlB+FlbdJcZV1N
ssIQ5PoMWivVNieKtNoox3vI/alzX8hOxOPpBJeenVhccxLLiLYEuiY7wdspikXj
tAcwLWhjdGoTu9+9CS92ywvvNkAzc0z7eHkhd7eaS/69DHE9q2vrwBqAslZ2Y5ij
UVDcmJpQtVbwlgInLCDiT2cJsDEeipDci878/74eTr7AkOLwe3hlGb2d81bEqltK
c2JX3LAYNjaGwEXpvSzihUXzx81TdIfoMxiDfIU2qRESr/RePOrcI93ZuAMGWKzy
tlrMRfUGnidS0a3OQNl2hepxSVFz4sIpKJGF+7yP3r01qHalo2Jb3vc0OiY9FAx+
/trYRr/H0kDg520zkr9qR2v0bImMSfvQG5J2ohl8oi7spXt/1xpT71zKAi0LUinK
7nIH2zb7cFQxiczyebTrFZaiRdrEB8uZ+gOQ2ZosLXD6pu1P+7qx5VfjdEQ2QK6G
kaaeg9+k6YQqU7kApQPD3NYwEDqM+g+KEEOmYdZMwNZsU2JM8f/khEGbMkfAMQLP
CfkhvDtiTQE1u1nfy9M4Wreo84z0Un8fP7Au/+tZ8xkav8ZCBde2uyjsjgo9uTiE
x0UQAZcI+S6UWKwqKrhamMjIDbyYtFHuvYyhj2AibXJhWrpTU2gmUyywifmTA2Np
a1nuWYDx9XA+zWgR18U6BtjrQ2+HPMG6Su70oVCWGbzknckIEXkFLA+klSD2eOoj
vXpSfp8vzt0mKv/RWjxuckGD2um4fCXpGg4ISZ/QvxpWZB6dvFbsfOaDezz9JEJx
RZTXC8cAreMpC1btAvlTuIuNbaIwZB3KQ8/6P7YtdG6+PdaFT+qrlG9/egqQIbFK
dpNL6mDchcPTGy/e5DCxibeTqvhurxkOcx4NH+8Z9yVMvhvit8ns3KWarJGU3SY5
RiiGeuDs94M5p1kkUXW/wjtlwKM27XnhLQ97MeEoj4JS78HM8TQ3lw0xdJPKYX7j
nAcePC36MXaKvsEuazdcUn9pss0e34S4no5NTSnTw6RWhfDJ0dlEjWC43VSlHSZq
mO54rGUUJL+BASiyPWR5l9X12qOfbaFUJW7fDQbo7D0MPVnIksbgv9jLykszRNvN
DDui2F6Fx1eWdP2zCpvmnrRBgq73ED59e7fwk6+zly5EqqLiBC9LJ4JIRMTq6ybI
S5gVdIXcLChgu3sa3xmmR3vvNDA6sNehKw+QmT0Aw0BcCON8LSU4kFZQTJKO+ddn
fersyk7R56q4pT3IVSZKGWwKMYLqxPZjE6r1Kc4gRfwzDtmnLv4gggVk0RSbQHL3
YZFT0x1FOLdDz/9GFX0mxpLw7fJEZdeFlUg6NPQmgQ4z1tBfXfF4km1kluIOBpr9
lznjDymctvc+R5zQnf8lnW+ATfV0qAdzBv+TWBqvlcLIer/xvlzB1sGfMT1h+fa5
JOSumKl7JwY+R91MXw+TrSjOhW6RiENrzFsa6hR/JgODuckLaY4VYeJWF6rftie1
EZAG/MuGLk/vgXtRMkQ6Gljsn2FWGAcaT9MBSOE5EYkrpw54XS0zGntaVFPZhLng
NHqvQuIRwTBgUCxJe5br/2SOwQihACeFovxZrnMIA1nkTmLe4L4nkORU4rQ6S3uR
kg4sf06JG1wu41z6gPyBjlftx0W+RnWT1TsKv/RowPsZJF0jqHTqtbKh+w62YxtT
DDTXjqk+PaVKR13hBBLt6IAwsLO+gu9bhNx0dE5Sf3wqKj5upamQWoydEAa7yq1p
FwVQ5Jl6SJLwh/S9xAvaUGjpih7uRLexHvmleAumRD88ITNZqupQ4W+FvM+9tqpB
NFV2zjrU3SaCWFZQ07KlWJIF6gqSDxzWatz1zZzBbTfjqwqPjuaDG1YKNUPUdK3s
xZbOpXOlymfO70F0cmRKL19UI1oV8IH+mVSyCoOTNQd1a+QKnTwaeLClUNzMYJuC
4f9cJtmb60g/Zlg5tc0LmG/fkK/aY+NxGq2K/8nwc3gU4ZBZJO7KcfqDcCcjbpRt
n2f0J1g5iiKGFqIeW9TP8Wy02cpeEBkgmdu/sglTC0C0rdJN1XyuIdRr0pi+BpHk
8o1fHEvb7abGzBxRVk1t835wUtZ0I5wECk5uK9GjBn6v8wDi2cwXtgfWPoTYCbsS
Vwv0gh0oMiEajBPPAtFYH9gP7FcM873IhgGsuB5wSurN5qDBFo8lyIhQzFSfA+1a
AQwh/kdDKy3y00TCEEbawhp9A6Cqva7TD60SYQ9+YSl5F1frTFCe848rm7xCqNkP
Vk91Ad9WfPbElQQk61OPPT0y4UHT8XjkuGBo2y5EnNQHphvWWN91ql0kPLDMWQgy
OTcUKHVpy2EpyGwO8mpG8rDBoEkT6KgoNlysUGAODhT7Q7prgOR568o5D7VJVGVD
WweuCNhsjma/RiYRd7gfCk2bdY8tOaxkfPvKtnUWLfhp68ixXmJlBZavzIa9vqiU
mG6hROKJbkwpLzO8xKZaj+9kOy0F5Re7kjlo/k00UtUsUKoHR9cwmWgYmI/mNBrY
ddtIZHLDXTpaOg6gEOE8aHrAEJ4FlzYtGGin8jNcCJ8JaXN6P4npVBu4VJ9sxWA4
nFpggigMkx1MlcPmDo4rKs5+qw+E8zcYaul5r10v1cHOUXeY4zdx0kZgCsoooxtO
UaZBIy4IIb0mvTYHPj+nx5ubds5dk0vkMHx0yQbslhLHOIeTHVo6qoIfBxoFXMDl
Dmuicla6QyIX2jreCZ+QGQhZ+oYPmfls24aVg2nLA4BEhmP8Q5ztTrLg0EEEBuXH
YtSvOT87QLemLgXSYDa5bt649cqrlVSNYEcl5jvtX1Lxba7paGpfLkYKJgf/wiQZ
W4kv7BIyN0WEQSf9fp9emXtF+apIZOx7r5YWOrklYFnyFBVxm7tcAPMnMxMuVEwk
R7nxZOUhKhE/uPHvEG5TFDQ5mOXnhFTTyJqPmyeKkIy8SdlvkTa692D+eNxeNcoC
lsawJg4mYrYV+Jd0S+xZG9aIedib/pGhEdFOhwKP36Bj3IldLzdkbWYZQKcRCbBH
Djguasn+aY1OqXUiWGvNM/SafftN+HfcADCdHFuusbmFozm9H0wPOdl6Fb47jMqm
1u15VIB5sHVhA+ESp9/d8sxLqT1EOVwS57y4oTj5QwdUchi4x56Unq3XHnND9KCQ
E1AcWCkc2e5EWiL8Vm68kpD8nks5L63eUad/5ldcSFqfcfpX4nO9zixxpiCEabru
JH+P8YBhrSGo5HWngC5EHG6/pSaP8Flkr0lgPMKrorW4iVpEUTwshwQFzybLdQHc
Kls1TxnYX8Px3Iby/TPxGjAK8Po3VGti6gppraPPiRj+ihOuefTxlDBjXQLtKTCO
0VZR+F5bFxdzg+edXvMZoJGCFKIhBzMArsZodJ2HQO1+XrG1RtYNda1RNdCZ4ion
10BI5f6revXlouGAoS1X1PFNZrsWHWIeHjq8isbyE9f/yKHuy1YNY1VgCS5EGpIO
ubfv7JxQIc7fV3XSeuHabxSZgC3MAfDR7tJ0vkTJwSn/phWldyUCE1TYZIHxJJrA
ViIzJ1N0ZffLJ608Y+rh0kTxAeaPC9A1Qknc2Xrvqy4KO1xYOjPJoVqTGcLPzsYh
1ts4Zt9UvzUzio/Lx+0qF0Abx54jh43htfVTELbAjNWJmZDysqfpVimHOzWAwblB
CMNdEBWG3aADPZrVVQa7HOEXbswT2vn4CGj1rpPSikZe8wgRV5UpMmbQpKgrO4nb
JAobZpKASLTcwXk8Jd9EkSgjp5IKmk8LcCKEGQPpFx0K61rbkKsQlPL1juj51bxw
Nw5yFsg7EAEcmHfZS6qlsJhiilZgJ2ta31QC9qm1HNtHyVx+0/N9+6nJD7PyGk8k
vEtIgqD1nbLsQnEcZch8JECIkVDjDtqAbuStwPQvnBKi5mcTPfYdkXsjAcTBBUiH
b2epyoyrmzcquXynQGYF8ZZGcNHxkvPAWDhXAy/XPJd+NiuV/g9c7SbnN3XBzQAf
nfQYP1Nktpdz59nVebXwibQ2MDvCvPXDJVRLB6dBAvruimd5dc6CqpBKqIuZ++Fr
ttk/S3rU4j+XBUVLQBH/GxraWD12exwQ4LphIEsJLFiHRL5axAmD7tmdZScLJ/xs
KIY9W4X9qSoLwIZkD11mKt0a27pdSxt55sIF2ndBti02opMrHLPcuBB6Q6ZeOFRr
u3Gm2ZPLom1bfsRl8xk6D/Mi73YEtYH7eCkN8kkUNT0LnAAt6pd0WqyoZophMIbH
nl9Xz4MrPH061lDjbPlrjWjpLdJKvLRRTaEoyvICmnLh25qFp8l/XHUZEEeFcq5V
aW9wrytuUE7LIhYZjPHjDQOCpPuz5AYjMPZJuEtUivXnvTx77CmBOeH4UFMXa0Y6
3/jK/5daRd5Q+GnSSp3hvk4DD2Xixxm/yXbDeJYx+BlnGUBjNec+OeGzdRXmiV6q
LbcEdvkIfd6sK9ZXKUPX7AFKHb8o0nBrXVw+cuKZ6fr+qEhLzn+erFKRpVPoVq2i
qkanmSJkOZcGznU44x3E6/1XFtAQSVVUqBTPxhGQPRwVMV9SbbDxDTrgsGcKGyUj
9HdsJ/rXxhVRfLpQaDLgKKBMycw17WrOwE0Efuw3jFWXPLltXXippytUTqYTGVZb
bq63RUhElo0RCUG/eUK+LH0aTsvYxMoTl2O683MDLuALQGbLID21B1sFh/KwuDS0
FQ9wtBdiili+PMo2Ocm5/qtlV411sSt+7qMwkV+fvknxTuSAzCUdvDa7xYaqbaNl
YgBvOOPIfpYaV+KihaKy8ELvyKi97PZM/MtxYpbD6rGTyKuwI4jpe4Js9AEq+fkC
XnchofUUou6jEnaQUKPYAqaswVvEy1sXZa7bAoOFZFCuf4R8PWJY0WFYhuPtiuRM
1mUYAOpJXpAvDllgSEqG2HmeC4Q9Mac27O1vVewDF8Twr5BUcDuhatb+oBXTZe7b
2vussRobq3BfahkMY8tGrBaeYiJAT6/EZbEqAeNOkM5U8oasgsTuqeAWQGeQgZIS
eEoQJAdfC2RyL9nhRc95c/WKB1WSQiVBy+8K9uUkeOL1h6l1+TAbACX7fCvXhWZF
ioxVmpWuGn/f+PISpWCDUbxIm6Q5SM68kwAZbOrCHnFP/DBQd1ECnlAb8QR8WRb7
o/78pG+ERnsrRBlaUpJBOjaGSxeZ7xC1WlYvNe9JdQuERoCJhWakIYnjl3DnNDx9
o6xezkJEWDINUufN6XxsQAmeiVlX6k9c5U9iSuS9Fz8lgCIVCmo9RuQ4dAqSMIVC
Ln6P98Pzdfwz1ZDbVBQYzHkL+Ismwo6GrSzjBS/0ukLkh0AN+pWiz5cN+XFojHKd
OE13uT7Fx01uhgseI/14kwl4JOf2pU/IeQutMw+Dr2JZvuQZJmTzayku6cTujlMq
Eo4OupVTjFpwPUmCaVrDBZM0qEn+UQYIP7drisRlugvkMibQMz4Y43XWaKst5muX
uDiDNu7K4ZhRWObby4kXSy28xJz4twI2f80uIfng1Ol8UGo1hW4RlqRpQVzi0E/l
BBEdaPjkf9Cz2cWjEKQfM74xL5pVz4Rc0lSbnqEO8iAu8BUFGkKfpmA87LZFfl27
kUWmAhIdItPfcIizO6leQ//UelE0UbpLa87BiyRZXgPnmfWl6AsS/RHUdF2JS91A
Y5Oz2sSc6uKZeFux3mCdR5zRmXbWAaf0zxWrd/5iCIA1FS999A8upvXolVBM+cEX
P+QATE2bP2+YEYKHjw86bdz20VdTgi09jdY1A1+CV+VEtGwqz8eqoCttvODnFXeQ
Xvot0boM951k5jHoCSi1WwUplo1my4oVUbuXJJdK7B8BMmFisj4mGfz18zGAMUWM
om4C47BKN2zkzllAx7xSiiIEO/gi2KnN4C8D99BTNhI197HesHNjlYTJaPCvnP+C
km8HgGL/mHfLb+UZ3rTbmJcpE4IL/dPNuG9px6JkEx+mnWtWVxE4iEt3QSEvEeeW
7Vf9eyrQC03VLDjIKyCjklOYK9qL9qE1VpcYex1sh5ELnECCPgHgOgxqt2nuNme2
9odiV+MPfvdadZUXAx/LMRHh/z225mD1UBnsoKBdiCeObgdAkY0JlXrOljMs8IXI
mqI68CAYS7IgRRXeHAJf0tyndFm8bzoK8iP5xC7FRzP4/sQ4fzWj9uuRM4XY7Eql
Edx/RQNpI2FscszAPDqS6Rv6UvpGNIiQPrQeY8Vy+sPD0JPEsShAiYR25wMPGVr4
RRPvyBYoy5Y5ITpPUTmlTCile6OuSMEyYCpZ1nmSF2WhspGt1gVzoQcmZA5zPFtY
CCKrqZ/7IE2qwGmW5lWkZc6AmtwnEG/uxMh6oTkR1tWTouD5Jh5qNOOuKKiLISpu
7slZSRjovsCiBhM6cKhaX72hmrF1aOi1vpJwKqOxsTI0FuYBJhzWT+djWduNOofH
UnOBaRFRx/imV5O9JnhITJJtC+McPheIz4jKSIccPPzvD9gNVYxsFGn2jI0ky8Wd
91N/ogNj7X5ZcWjhHUtsnkIrgitH6+IYnw2l2Y9BpvDrMFr8KZv9bj69muibdyge
RRvp8oHFcZNCdnfq+wEec5+erMINecG/Dt13rUHIoNlDxu5Cq6ySYz8qCV7Y9Cu8
AKy+fJOsCWRH+iR+gzCw5gfpFbYnDxiMfVQKXrBfo9uqH2pLvzjdbFzacTt55klc
3fXTaOuwKX9ybXwQHhj7dBHAHcI2FY3J/tRtQp1akqKriBdXbwW7JcN2X+/Sad3q
M2roamPDtXmgeOy722OOUyzkAm6Kj7JNCUWfJSNl5KJVs1Kg0HgvK6KyNuLOy5NH
ePOr7S5C7PiUlZxxaHuLT7dRE0MrfCeS9qTEeHNPtiftejn+RxkXB30NPEsbDnYe
Zr6BiouAeCH8XRQ88EkNvMfwXVgL8EptY5kfpB4f4dVB4avGniMRCblJAA6DZzro
qekK1GDR02fsaKLxsc7XEwZpXBpNeuXxvZxkxgzH6I2Z4MlvwLopepHQiCzPhf8C
uOLknZhNRIdMbEGw2Mn1LXdzC0ynW5hSy3v6JJaeh+Y6p0XAxmAPF4YSzxvy1wCn
fmaVeImn7StE/ViKbcBSPqkZwFOA8YqYTHJM1Wji9Jt/FFqjFTLyYfgZrhTNdKlB
56lG3ZOeQdt+5fgBYEj1mpShbPhSH8c7ZCCf7xNdjzEYShf0NH8Vp8cp315UNmIA
cO0eApAr2ui5dnio+QfVgux1GdIDxkgRV9WIVP27PXV41O1boldWPdDA/Fw+XdjC
Nf/S5ZnFVVOKu+9gDDNIZzoD9hULZR4Ow52BFPyCS+auwFOa2u83AoBzdmtLVjvO
n239O7pUX9Gf+g9FQHCP6g2D/oaNnNSqauB9pVrsdUmkGP+Z4v8yqwn+AA9SaYQZ
ptfSriLX2qfeQcp8y8Q7ypzQxGMNDXoCLKEW00IcxuNiySqZrLrcL8Qv1wvP6AOc
07HB9Pl/0NUZHenkcO0jRB2gj5y+oM6o8wtlQfo3hCWXCup++VPw/bYxrSjY41pn
/Ij2eQKzgaZ6lmIWQqUO3K6Fa0LPuIOYiIOVUA6UNDVwXUdvCu6arRp4qr1qNoZZ
/P0Gm5id8uClTD+doz/TibFSf8a0aVT4CJqR7fCg7rXR3V7FMaCJfoj3cdUl1lx2
BuFDugMi3KfRDLg9FpbMiQwlzViBUSeo2uCqpnZ0w19SPz2bcCUO+YHrHe7ZEaZo
xdScbXrp9qgGe3I1LH9/+Q5u5WGoft46zJlSai+FyA1PJNSy7puDKolJETl25rXh
PSARgwdZd/NTZAO3lnmfJj9wwu9lBCibj34Y/9DSsEg=
`pragma protect end_protected
