// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:35 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
OQNKp8RWc2BPKisAoAzBIUZ8GPsbyGI7MZkgGc40BttRpi8N2Pp30mlnj9J8gsmO
C79x2v3tqsOBjIWcgap4lg78H1v2AWHb/nWVyLxHFQ0/1zbF07BsEXHFsTJx/ZUl
DnGSBEdkOLvgyygbmHWeOUfdJLjWv4DbPfYwvlpT3gk=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 19584)
yPZfwqyixXeXWm3CZrh5TmpMbOmvFqPwrgUCJefU4qiioHYf7uGADIgIxGB5oowk
ftIyAGnaj1vqs3QK+265G7/sYAvXdx5oQKgajaNaOXyG1sg9oaErAR5547AeQRnp
qf4SReZeOhUZuzW4WEWPXLqRcT1IBTZg/beyKMEIoq3PRCDAzAAiA2Tmjhvo2tAy
F48CU3KX8fxWnxoQm0obYO048VRcm+igJnjAlDJbcfKJy+t9UfxztBkBxNQ7KsaI
GuNh2Dvk6RRlhln90WsZ/VnYoYnlymR9Wjs1tS/6MV0pYoaoTQWomwdy0imqLnei
NLt23eS1yxYBcTbjtd3a2u4c0atN/DfW40x+7v7/O3Pa1pKMV1Bu64Ka/j5QQcnX
RfJu65Xt9YxHL0L6ZYdUQzbFxjtbknqWMJeJ6uBP9ZNCoXydBFxVLy+cZFxijlNZ
FltruMNaRCOn++2M4qmnrHBesB0zQQ5yAik6cxbEJC7w0e4biBjSCc776zFjzji2
OTumu71ZiQRjs9UOfu4lcK9jVOGX8BY3fE1Lxoxf3SV5DdHSgZN8HQnPr41NvNxn
kEJN8jnNRnMwWVpxqKh2eDS9pk93OeWxgFJTN91dg9H+zPEKmmoNcbW+RiKDf8d8
AjPBZEtF/GHiNxTubTcv3kvfREK+/hV5C1GoJClZfh+5tsJ8N3MdaAu0iYUIU7JX
+yFDVZKaZDKEQ2lJJOpGZqheqvWQU+jUwATCRJ1YSx9DV1C55YACkqqZHfZXRSN0
UT9yy2s2ovLHrJqUpM8IOpLKs8z3fiX/aPatC9WUtToIlvXBxZo4e+/pVLT+zBRN
SXPTfrdNRkIfyYvtbs6M5J9VRpmC5/JpdUmwhl+80D2eVfShRqcFs2r2WppH4zU/
I3og5ipc4I++00+VY3iWtsKhiUIJdn5hbJhHfC9lVRv/dG7i1Itm0GiSDXq7EQcf
8moTpbG5wIgTNVtP8Xtri6acGBXySp2YMEZfwgYCTX1lB4V1oVxP1THykpQWwY8h
Au4epqpadcWOyzbTySkCPxrTjYQLwJLfFIaiOpTrDpA5y5DYixs0aq7oJXAdf1Fy
ZwWa595KHO7TXSulaqTDcsCvmKCZD0zds9oCTd4r9dcFhK+uSsttn+h5IAd9S8EH
AYYAK6sa5NwgwwGozafx8V9SDTJ0Ew+Ubd44fkLbRp4hsviPyu3lbGTuoLo588n7
73uHHkJ1CfeNkHrbx9mPXnUFdfVgzNH+hnVcb95j3GSzzydw7Sf5q2R+9I4Q1SyT
VFH0NOvp9h9D2ENtHWiDMydjrd+i7lrgBarnilBZzTeqCFjHS+3yiXL0og1zwLgN
sOQwBddhB4mIIfSFX/ONQhWyoy7PLLdQ/qDfDb/Me0toAEQVZVNKkKdLo+GZQMYt
dX2KNjKh22oflZ6Tzs4frbAhBnwRu8LBXtmSJo1usa2pt/ffhy102a3yL0G//i3p
9oaawOiDDI22MVlypHq+gQMJh1WhBPzjgeIsLmn7pgY2hmka31ifLCUj1ubJzMjS
NFJVC6mqZKRl9Jwswoa6T0e01BKTiIIYVIS74RqdIg6/BO0ew2eSMM6xmRHcI4QE
Gqp5lQkYpWbIq/CplCfzTS4251MJ1pD9ag8wDGrxs/tBSZMk02de0z4mKYH6Jv06
7vuzLfxUarrKvBSrV6XqaCunsKKrA3S10e6tzoamvxZNJIaTnGaYsZRikU4QmiXw
ARf456Gt21+99BMoezdnVZubVt3lYdI6hWJnaLk/NXJ4CUMn4JHM7pH+lW8s2IVn
iY39m8uSeA1mJYwjSFn5s/qQKIsN0p4QjpS4IKn1tx4zpBaBlOiSZ8irqbgH80Vs
HhK/mynEHu/jn40odG7KIbh9HeVyrpNPX0RMEO6JA+J7+2otTkKCGnllBseaEk45
yAYDDKTWC33Q2L5tBlB0KjZQ7+lSUmwD1ZFGFh/0EKL1VhcG325VPQgy3MQJ1VES
Bt59Z9vRT6Mp25hR/xB+zJl9lVciCS5vu8Krx9fNaIVlzj+NrdJyM0xQRt/mtcCz
6WRRRbunr5B2fiBQC1n2dK1gKNQo33U2qbIDAIUcqY1qKe7BiKv7Ob6WnU+DrN9Y
N3SBSkGH1aNsI10cD81VIrj0/TlPFtgZ+uAjXwpU/JbaBP9CP4cyyW+j1Dg1KWR+
QWlncM6pPmdXWM0JZhR2ltg/5oxxHDqKRXO5ujigS/bLOFMvEQzFnmLnYhA+17z5
CHvDo2z5IbjCE02UxwKrODRQPtt5nrfzdvA0RUiIzBq/dnjjj8jNXXmW7NVmFh6e
ijuHs3UCEnGy+p2Jr/oceA6+i1dFdpex2tnF8elYQlUqx4D9mtssyXKT+Auc7a4p
GwtIqoxr3C4mfZ+8c0vjvcKmig8q44FkuxWbG6/XIQ6ZItaifry3yD1SfrgRFV/7
d9AVHKHn5KdZw8XBPtifHiH/ATft4P8ixaQrzyLvkByH88gAb7Ut46rRHMK9E5Db
gpFi28VVMNS5I1c4qsmZz6YTGVUEipcEhgd1KxVToHd68AfbMAWcJExzlsNHwUbV
2alVfZptOzud24mKTKQSDZ+LLrcmXNpyaJLsUUceFEKyf65GRwuxH2Rdrlf5TPp9
0Ft6vSWl00Fke2CCQj0Pjol70dtGZ60fDGk1R7JZOwNwSjsxFsrl0AtIS7C/sD4m
XRZZWLrEnwWlx/sGq0a6IczmqX9xwurBvsYoeby6uAYYDSyJkbN5duSWFeXt/FuD
WE4zNsUIjdDHPS/zdz8IklHRfHpUEszkdYdQSFP07XakHHuguDdf1bwtIzVsxT26
dcs0S+tmh6em6EZ9BECBkOVMt+t1dg3QupKQBCONN2C4g7Oi9tgwsEaeeEY/83Rh
Z3/2QiMz/lQ+RAhYZycE8VeyN0JWKzxuXmsAnscI3EiiTi++PwajmDbA1TNNQf0S
nOfO12+toPpqJHHlmRB1+5aGLsPetd+8OwaJx4k2nVr6QiM2FEvA2HB98cF/snru
yMMQ0/cxcXJXauBEzyev9EiJqBWfRP9BQpnJ1jEGX7ZPGDrDRiHvK+73axZafj0K
q1Za2kt0zabfmcqR8mKggo6qsdrjk6onT74CPe9dUdrSPBLi67FNvDLvOr9bSlhl
8s8RwyS6lSi7koxBB84OlCP5enFvdxxfg05U3ofQMKz7bU/zN4OTpQ86rF0Md8U+
zdx3h0GZzi1ruYiJSCFYWH1AmPOmZOrgmWc8+VDDTj/EKrw51QkVSur6BFicpcUw
AKwgNdpSafQ/6rnRQmmcXx41ZhQyq4cW/lKDIgtykSEJsmuphGajJF+QEqW69+06
aAjampT/CIYC5oku2CZ5YMW6bOswy3oF8iO+loFPhhxfL2BFC2U2eBM7O7JATfjA
jRxDV+mdLfjvDAzcdJ+GKwlp+zPviRIulPFq9y30LOfs4RS6OryUZkhjHP1P8nGM
/PVtcyyQZeyP9EufQvCzusU1n50NeCg7PfbuXY9pI5jsh2hw0iK/C0xPf97uZASc
WI9HBAfoPp8+vEkuwQOS80zW8/VahmPtphZu1Dj0s66NDaqWFJZrFMgV6ZhlU45t
Z+1UEW2O754ONjFt5kV/TdWAYHx7zNYkpleu57OzEEY/Y1JtejaC3ybaJa3wDOH9
8yqZL5vYTvwNKzyCmoI5UBNyutjB6aIuUQcc2DCiF5OEvTa+hTFq8RhxnbqbrW0u
wv3e7EaMdsNbxLFlF6ddB8Ut0b73gNjSMJPLJeHxXO4aoEJFA5HMfSZFnpZ86DN3
v2KvFM4khBJOOaqjlYyE51Am0dObE0/+xaNRnqdxRYIvmTDA1Q5Amraq8QXZdqWv
oqFVWmXtVsQ7dRQv+NtDtbMNgGcXbZOi8N1zJIqQiWY1Tym+jUZFdubVj4ZZ5JNo
JNB7AIB0oZUFZte6scBTbm77YjrPV9zw1P+kSFEDY8nT4+a/hG6noix2usxJm7r6
eYCeNDtPfkPBVEWMDNhh4vCovyjlirracbXlh18cWOR3uohKn4uhtIE9q5mdWY5F
0MPsomR7vlQRHrRjOUvzX33D2wpxzlXLYynDZ/imOqGIINFrxT2BnUWDdt9T/++5
5hABWxvp93ZzaUNMosTpk18fB6Go/TdjhGlPwJZrtcrM1yAnv9D5LqVICWhG+oGV
TO7SDNAOfINNHxReQIBM4GSgF4EDRkYbwiERQRZSRf7gW6OwjOr03TRUF4gPV45s
/RXSx4mh2C7EUOguEFHg+WMUx18EQ9TqUjsvbTNN1nv9/VhpP8PbxV/aZKqRSr9P
cQbQrbZ2ODoTAvdxHYycLSMD07l3lSz4nx3wg6DnRlM9ql7o0V/alGaR/FOfCnwV
GaMr9ZZKvY6WqgTXhu21EzEO13AAHYQPBHfeOooF6BgqC4aHjXYEzFJ9U7f1/r94
dMmNV6yqqngBol0MTuaTSwet0K3L7yf8p+CIhDU/4foEbx19ZeQ9QbpeIZ6Um+cR
wco6nE6Us/K4RgaHqTpcg6B0XWlayN5r8WJOfHl7jbwsl130ZnPqv4Oa5mygvjgg
9cwbqETdX8xCL9r47692USd2MBBCHgaOtIRfeDszu2FpRJOGZerbrpjmSRkShbI6
74BZjUC/ivI0e2j7MB8h988z6nYWZ2fru6wSGPaS6A3gGC6nPUc80wolfrWfVUqO
GswvVly1M89/FHGUNXxHGYFlzrs0ITgnwJZRTjwfv18ZhxVzViEht9lvop2TQ4V3
cP5nky5fGiD447Ibu7VWb6Op4k+oTLJvtkixiv3+OlzK7AlBQtRW8sxBkkwh9tKx
St5tFTDjfe6Lqy3lZA5vqP3Hy7MjQAhRf1uanNniKzds1QbEfUwedGPsBjVEEUuj
w8EBCgCwo+rxtYSaGah1T2eGcxA+rWz+JHiMWB8ORiicsIS0BNA5J2iC/xg+RvJI
We1Dq9p9XIePBQMLGwogUHZoqWNs81saoJ9toJQiq0YJtKz+9tJf7e6ag41/2ckq
t92KOuNbRPuuq5opZACOdYnX9/4g9m7dydHsZQySIWpelMZdqUhL8HFM+fuCV/8C
2HOr2W1CHhOgGnXwA1KXgN/Z0rhn18m9JWYZyNOOI03MDVnnDwWn2UTVkD6NRTNJ
GiT6NXPty5RdN4TyUfRN3+p4UdRlKJNOeTTjX0pIpWdc1AfJXV44vlTnnqskzo64
P2ma7/HhjHAZr6RCF0Dn7m/4nLfob7VKm8LBMmbtyLNCvEg8BcAWVtgmeum3AnhI
qGzwYohwAt/N/2WuMj/P9yOxvijod6U8huk0JqoLJPRHnT1ussggDhoFOO+67KXy
/JJ4pGXLw0+dnHwk3Bs+5l7wyeeOS1rIl+JnqcPgxF/Zv+Begf3b5bg5ESPGGJKD
7f+X1phCkyzVPGmJAMgD0P1pRHMu6f4hGR91y0inuAF4vLf1c83A+CW+Dorg5Y2z
QhrS0X9jO1rtpMlYRoGmG5SoUTLuwat1aXu/6rI7upQTsIKAzFN7GKK8IXGqgKXZ
GOa9Sdm7b9WRipZ5hQ79KeBAeEvC0hF1yqClurSuybMFRUN3f5EljuFX4jhUDauf
cezjSDJyWkMOD7WMIS8SApH3spQTqalJIzdTh8g5ZcbvcC2GT31ZvSG8hkh5G2cY
CiNBFy8WPIbk9qGnVc9tXNNrgAdufE2UhdCY8oQB3W7AxsRiEm1srsIJZx6fnVNn
Kr5EDosoXba4wB8kQwZJ+C1cPiXl3KssjxkxCz+IrSY9kCxjNu0jGwftmvwx6X/J
CmMo4esChTwpWHmDJPGFrOj0cgrJVS7xdJl4jfFF6tbvckMMk+zMJKZ4fX4eYUZB
7nCSiWHnfxtlm46JoX/TfKFKhSe4EKssWlXK/irIiLV9F04nq1nB8qcAgh/0ai4m
s13UJ8WPg3VY/8q13fBS6RFOrZov6DJUhi1WvVQaq4F1OwSKoYTGXkDj/HDwhWlj
B9Lk6+haU/ltikf1fNFRJ8lJue7AnG7Nejtz4eQj4BqtOF7TzA4yNSxYBxiPMQBm
q/+acOWH4z86Gz3TYzan9RAmpOB8OTYXyFfS+ERVeo8CujhIX2Wy9zj149XvAItP
cmpeqHwJQ2r8ohgTaqZcY7xOOfS14AuZAHUwELctPyvVKUc4RnozqL6y1vHi4TJw
GNRVkoVzjMxFHwbYKPV0/JZxlweBe0MyaDwBgQkk0i7MEv22eAFUi9cFKK9CIOkH
r9cqw9ckYBQccSj8nLtAi955nnSAJcLCNaFPGDByjvH5BSKq94CAL+p0Z+Ryatxq
mYoe5eYgCUkORt9z4hANKWr26tWX0tmWpWmj64xxNLRAP0VY7rjsa7SBdDQ78MEh
VE5IarLT/UP+VASZF2SJk4ZmLioTlnHTyFce9t1aeOg2BmANdq/TAQnONfszB2Yy
K6aE7ZvogmM6TBXo/9StFsuchxmwL/eaBXydovDHn/pAZVXQTce2wyHslkFCvqcR
VEP2++KpurxKNnvLh06oj3/kQXsh0oLwwZ4h3DggOFuKaEr0ZL2++yXpIh9EzibV
Mf1KB5mqXVaobPchHnD8+/4fRlWfHWkf05fSbLuZcaMOF4+4VuArR37pgZbthWIJ
BR+CwEpFHbkc5LFfSE/KbKl037Q896IeEFDJnM821sfTRPCPkkTdFzdS5d4xIPXF
QJE0fYz8YgO8djB/8dtwttHetNEUo0/dqUiaEFKC5wcv2GVBXbyKSvOa2u5hI4BU
lKsLLLS7mWBG+RxpSSR+4X/CbGjc9zF72GPmprQ+HNhghCUO//6GNzP+S7DWjAJb
QGbAWWg76tCwWuJLyK61H8u5N9y0G7F5QYToV5+YI+lqIgA2Um4U885AuKKZ+YQw
Bc2Iu1a6T3hH1SxlIUlR/6YE37PK4w0d6xkh7pxMtqa6BsGLH2oJjCQcziQKDZJG
X7/cu8Ff9YRgDL2gKOQ8mPjDNRc6C35bG0WaKnxBXZMe0hVuvQzXoGjaA+DGBbyw
qnfK3PIWMe5PwqEPFa7SqPHmDyh/Jy1gozOCJVtO4i6yyq5dnA/gfeIpoSkzBKD9
inwkGeoluTABgjP9HiJ4GRMw2dYbggLeshbmkxSzHI3q3SmN+uIj8KEFNmYHQ90X
owMONzpA5bMSlyQCBgTjek5Z92A82EG85cYCqvdZHk3C7CqSphvX3OfWn94Qmttz
Yc0KuBD8h/d+RinbSoRS3xZFPCgKMX3Y/Zo5XYKQVfIqW9zZSVqthqQJlqrFq+4r
vMy/rWWOhp5dEThrBMgU5nsKQ4tjcWWIxzYbvR2vp4DXezr1iKsMtVEaCiMko5ZZ
vXcNECeMEy8tLRha3GjnssOWyu1lMCnDx6I68ENRQvynjJ1X0/qN+nk3BQYgNHz0
SNIKb5ipARbOWqC9dJAtXniPtbPYgZR2Hgb9wsD1lX1/66fYtG+gfAeHGY42CRWK
OrZ097KSn3/BHW7RTyddK5g957m7C0fSn2gDnOd0uE86p8PwebtV3Sebvt85Lan8
GRpPKWR3juOkod4/x3VU+PVosP9WtZs1YEGj899nl3RleOHVDAyf7+iyuhRl7CAo
zbkxg/MQRtUcb+xit0YM0p0e42QTC41PGwLcsuCtdM26ICyHKjN8oeovvtBS+3u3
KVkHO3tJ72mciQBpbYda7w9biegOuC+cjzU9zCaDuH55Kx8RqSHEp+fKOxSInKUU
QK9vOnu4ScboVU2X/kxvmsh6mR0tq/T1UfTEimSamo5nlY+niHgI5ZVkc7brvt6p
CXDigYOU1+taJc0uyRUHQo6ZopT0zw4+vSB+xTRQMhW9DoSCufmHAGsJE0clOQMN
ydRNcjaZ0iBVu1QzdevJTHK6qnkCI342jq6kI+CaWG6XrXBESoz0wnBN1Qz5fQVI
8CnfuWAieJikLeHBp3Ed3UshWnDIRiahqgucH1jdorX5gcyyT0iq/jVv/q8N08Mf
7rvYDhIXJiNIM2mH13PIBaBXcXX7QT9em+ORSfJ6t9WMHnOwDLSpvu3PfJv70rLk
Q5qWNS0ri37noNyKwKOiZIx4OLOppinOBQPLVZotmOUPOE9mBzcQAITJUdaEt+zF
xC57X9jNHO3C+EcNNmmzzxQmGsaEHI/yK11qx/OA0lCudbimzfJPxUhtZeYI9BwQ
bp7R7aRBt41oWOCoSkA3J3kSTjZdbWl2mwMPKc1lDIk4svfKcKxc7+dtLyRYHp28
l2JhVUfiIr2/UEVVsoOgVByKSBwYBDchi1bdr0UPH0Qf313yf6kZRXO8MKrYlbu/
xHqnZ8KD6HnLdHGGmKaKTL+kRnOIzzW4hqewIUfM2PxB4H1uVb7/M8K62traG1fc
ObzZo9dSTns1btH7/ayzQ3aZMToVCj9aVkVYw/lDZp7EKYAwIH9jrtD8yzGpG/5m
kBr99LoYU1wiJ/E8ChFyj0POD3e+EYksqkrwjnfMsSJ3+x49B0784uQdSweZrPDB
U4SR5nly+kIovFfVoO97LbVryyQ6p+JFcGUruu1Pt1CWlF7MOXwVAXxaRtd4Qg5F
kXyKCJVMHdlr7ELSoneFCb2409J86Zs0hXIAOaaBFi/wv1LxHPoF8IOQ7QkAN5H5
jFAa2/kSx/B8MjuxBhlXZDhlSrwv7YN0FdpXgCzAiw96KSXPCtXS0HTh+dwvm7de
20ymOxICFMhgvZN1tVIkOmh3HJsC+KY/Y9U8GA6lntxTi7jUYhaYj6R1SV6o6bA8
rOOpHsirh5P8Zft4k/HzAQTzOG2vJ9iCxMYqpAmGBI3FOpMU2c8ZDpk8w3Ul8alh
k0u7kRN6wjqp6NRVp/8oFnNa0eTVAk/WvXl9/dJlcVapZ4kmrhDVjti7YDkpR6v6
QBqHJunejb2o3YL67ZFcGOnqrILJKd8lpWg/yngziLdCNiHB6N/M5QKy+2SdN4Xb
PIx799lh6Mbo7oBf/V2z66zQnQVkSaAido8Xp9aLikgKD0UZDHcv/09tfPOHqoR0
I8CxOxNjEvW+AMbd8s8XJ3UOGUs8XzItR5crCJrGX7sjdErjoUXgBeKTRXVxK6kW
mf3iWNWa+z+G/FlBs8VJ7krwvT8TXEA3dY/kQK6JHdcjgB67eSjS4sNM7/vxHXyQ
uEehd9exH6GNj2qFCECUuiH/UklFWwQJFvtxatio8s5QjDpp/8ckBDUMRKsrOwoa
mtkJFaTsO22XzikRcYso/YNckQ4+lYkwf806jkid6mNkmjZksAKvdSU1R98/YKwH
hm+eqiMo5OAoO5fc/KAUPyeCS4DmNkIyBQeplPmYMI1f2Dsbm+JcwMZCr9KfdA2y
S7HvW2wuUn960IA12o08csfHBjgNaH/VmyRtufE/Bc0Vwg0RxFQGC2dDU3vIqscK
yyMftMGNPpLPiBeGV6SpiPb/Azr8ggvAjmRYGHGdBJvKzCGxG0TxrtQueqwHfrq7
QrHzhDpcupKSxscVHzkbJjbKm8jBtC1oAuoE/WoxjPX+1wLIqsLd3Dhn8RYO8VzI
BSnEhsVUEE+zGsoh711hOrcssy1kLRj5o0sYvE2kvnUh7o7UywAyFOcCNcQ37AQH
2Wn6iU0lyn1+Ybn61PsQqwXBkkdjL8XDNLku3NJ0exCQtFChz2JamvUpweALThNu
yEzwonUFjONqBcUmISVC3hz9yjexS4Q1krjivJ81bwv0j9KXCkorZqqYKxMG9cLF
AzgxtK4r/d//yevnF3TEaIDqlBjjdpPkuFUar9YUg+JGHlhsYejJo2EGBA7L6y4Y
Ypau56YomU3NDn4LBx9JsJi8xdcau2oZ99zaByZBfmQIf3KvfiDWwvzV5+h6rEG5
kJUOpJdpPb7vdiYu4c/6zonU5O5InvMcTNK9JIEyDCRL6yyZYs7HGhFTF2JybDqu
6/zhtLSxzbFLXtSU+8LwriX/H9A+dobS5ekTwZ22XQmEQlGJFL+ovcxOwlCLqjz8
eb5tWmv5It0Y3f4yEC7TYCEX9gJx/ojlHeP7oV7vUQ5Te/yXQo4Q2qaLsHW1ps8n
U7f0w5rTsdNY8UggCgOuwzrJrmuE1As235TzLhFIwEQ5ZpNxAtpos64b5t9RYteN
OBeONZvmucI/f3oOI6s0h1ezoljuaEpIqfzBuOz77fuOYcmhLMPKqo02hcbWmaBQ
/3kfD3Y8YOeL7F5bWr3xx2D95ZXFOy+dwudO3h5U6PuJ/vo7U9Cgy2E9k0lcbus4
6n50+IKRQfFV5Pi0pwTCJXz0lEc47wVmrDsly+bazf1yiXiFUeqH+NOgRh1XKqwL
LEjbiFqzXJGSXrPvnk1+I66t8ZtPSSh3HuE57N3IlQEJNxNC7UCfUxegJWvmzHdA
2E40JO/C6muDs2N3XZhWB8K3n8Eoe8RdPCnaoWNx+RzxvSKdwvcTAfyqAurWANRS
RLxMIoUBpdAiDptLtUVX8rtNExZ38k9Hd1d/eqoikrjh7+4yxxoZ0z0noQl2XMjH
ot0WqybmwROHfTyzvZP4wKBGc6v52MUFC2+QZQXvRIL/JDaT+28XRzfY5YMLlLQO
7FXUr/ECfN2oTw0kM4edoCyii+7PxqXPBlyI9hvAK0zScVSMNdpuGz5cYQLoiAH/
/m9qsv7K3MNhCOulzBlJGWUhbucUUDNnddQeObc46o3JY7MbS5xBWDwS+Uctq8Uu
NyqjMgOKksp+mdr5Z8CDDsKNWMkc+4Ks6Ya0jLZxYt9a3IvOULIXXepyuhvkdeDh
aFFCC+itd4OYSqmH2v8ptvnuOQPyLiEzc5fjKwPatlI9Topbz/5O/bops+eLPLnI
6/QLK44whrqAv8Z8WrvjtkCZZKLzmA/E8RHuTMHuix7sY0k2PuGMiVdOEaewsF34
9G/geOfkA6YHr+fnKaa+NobyGs623q04TcnxOPKx+ihHm4qm13OP3Pp1Alt5wOdB
LL325btpRIydUfbPvJCfQyc2k90zdO7DPmVX60iwDL+Gvowk8zD4xUPuuw7x8C8a
GV4jV416si0lUJ+fgMl2IHCS5FiYKgArUSR2nxM2kPG/9YayWFAIhIOUu9nn72i/
pWrM/saApM7hgcs0ze6zhlK6MLDC5dGaMGH7uKYAYMJ0ru8IstTjrPdCE/E0+l8w
zHG3OtMukCXV0o0OT2fxuwYv21SO4ZA5Dh/t/od9gMNn7nEbYZ6BGRqLzcdfl+QR
I7zXs0/M3FJQHdY650arXJm2+/3LJrji+RFcRjjQvh5E+XQkY9V28dUkiLqpS5S5
413AmDykPAkipYWrGKXkI4QnOOK9tmqXGX7/Otx0VVhrDxU3uvswPR4Nf/aeUKt4
J6AWB9ZNhi77usdt3roYBcky350Q1T/hPiEBIUmsEu7FaoFZ1qWdHfcZhWYMqKvC
NNLvuyXjv8ZB87jCNqQIc/HN92yl0rFKG93sLklvHiGsv+YB7FAN/LFI6zcRi7wa
RuMHhQGgEWk3OFC6K2u6zpWgvmVV5OfvnuTM3efKLlvU46Vpx6cpyGLMlLuVhqq8
cDOPjSXEcHOAB7rpAP1M1K+3gyRfpnCjG7dxFDZyYQAw4DSSdTCgmrrLPQ3xqYxx
0GijDiIezowK9fY1LAZKkZpwOECmiAGvte0U9J+zzgdiYlnI8unZrhFBL/EbeIeB
tTkgEohBclH3bfSz249kNjHOnHCfyZOg1wVDu4nbqZ+xia4Q8hysXCVQC4dTcgDc
ACfmDRvLCcMmMGA3QZTzUONtXE1iDex7lgTKtlJOd0GL3DMylw5+E0dX4M/HUUXc
x672EHUSuQxfLqxgdN/cOjczZqiEtaVzjPXL/KLiuR4e823y0vwexmfAH5pYh1Fk
wMYfUA1N6puZNMLOuz8y5ul8U0uPc1tvyA3ng0CJut8Zu2jsv7gVWxKztsxsrfRy
7NNyVr7MqhTn8L5A/vsGxM2WIvHgiVsX3t/J3MgJHe9jrS8wgP9ggprBas+VQqsr
QV2dm18CXDHTUizJ9vV21Nw6s5xs068F9WNfa+XqPavcErdU2TSiA6RB3rnnBFut
Ql8eoCDQff9A1M6CWLMQdPqIdaOC1hruOmMAKqvoiyB7sDcwTIJ9x/QWUbONgbu8
1H6x7rfsFQQIwbIJZwiZWEznn+oAFUocDJAlTMT9J61x/XdRDqsekuX+VRBx9aiw
khCdbN09paVWF+JFaVg7OAUg7nmTCNOoCA+OyztRxMZk8Yk2tz3w2t7sEfdthy1P
/R7+sRbG4TpypaiPHrxQ5IW8nP5HyHS3HnRm/AnijRe76W2iX3FWJE7nGv/yGNNc
ttjQK0kB8R1o+iNoRgXVhzOpwF7La68y5ox0GQtA9dD6sNO44WA/T08gVxqgAuZx
WO5BhthFRsgUo9zCbZ1DCdqx0Bas5aCgI7x5+nBZhysYh5a26H/3lemcZvgixnUh
Dq83t1RPLjgX7blq2O6fVN/cjJVXLTSUA3yAjbU2/i2J8bNs7U3khQwvFOH9xILI
Dob3Tr3jQKqHwiLzbnf8kMcGfqm0bh29dLd30LlzEg978p1TLkWJob0BjYWfh4c4
ZiblhBdofV2MkCJvY7uhbwx1PaRp6N1AgD4sVxZz/H8FjykUSTN2/Bg1wfeOQ/60
nMGCt7HMg2K26eqMUqCvBiy0SPwkDtbn80VKFbpiYQwfY/giEDDMx25RX0jPrkWI
lhAiSZ8dvWFOADtfDTqkK5vfwTaOQh0Y3O/CM6gMvZp4nnbUJvaGbfEdQs5yZOiv
h1ByFXrPct64xI+jnAAlO0SuJg4/+QGe7fD18vVEfMGQ/L9X2if7fBVVjNl+BFd7
o87OvOauOQwN0cpCsMs4GYiy2qcp1R5Z5XlBgFSzQWcz8v0/MPD81V0CXzsujRbU
I7Dek82PXGmVZIKI2H6jVILxNJ9sYXXUisWf6KZ6YTFCRrcTMICP6/dDyGT5wfB4
hjXT5rz93oEJOcAvRTh1DcEZjoeJWN7nk273ZDw+B0er/xAqoMQdJL522rv3lgDZ
b3sXVrUFTl4Xv7WnZvaTS0GM7GyVqRr1iot+UVH6tLYKOSG3mIF9aKsdsicQRMkR
4jtep3GAY7o/OqBa2br2F3Oh1I/RVEekAjZFtj0OO4Qdu6wWYJqz+VXnioilSxEX
zH+/XXo6YD9AnKw1lerrELBWRFqYvedWCK5kxW9NZQUU+8xHmjSC1vxv7S30d8mc
ysTaLi834NaURC/u2YYymA51enI359ImEWk5bbDAozM7nItJkT7g/Y3S7WQxHXzw
pvIUQ1ikwKGoCcAA/Vc1OK138NDRviibG14JGn3wWzq/lOtnx+jpDQPvjvJNACZH
KgpOwgcxfEXerx22f+cfoT+EgCraLmQDsJwmFymbKvIKXJxBUnswYVkbse5at0Wt
HBZ3xuSQtmtztYOTrLaI1+K9aqO93JV4JtsIYGoA/5vPpPB3Q5fdiHkkieO+D5He
AFIZahopwWDej7DLDTwD5t9RkFnD4kNv41+UcwI7grtiC6gtOYP+6EB6vfPp6suy
H8RYfBl1iBO19pD12ifCNadGeQjx88IZJYx78ml/TQQoTBfntIz93G26yANRm/i+
8BN4OGWJGGZnz2es7poLYvAoPZkkvMu8j05O4UxR+GTbjXuSaSAIuEjS6KKpz1Xe
hDSC6iX6lMMXnRbzGmrZgZQLIYKrNNBhZwlsjrobqN57MzUk3bDdHYQsuCh1U7g9
kNeXY131hYmfyzuP5QW9h2NouK+zISlH23tbk6AQMT5dNR7/c/IoZ2//Q8vAGrGc
ssbjPiXCulNeIGiQcECDLdD4fCGVWBB6GjvPgK8Wn4M7TYYg3/7K9lhcHlE/owIo
zHWV+5VZDK+sPWl/r5zonVGRU63ExL9WKHgDieouI7nze7W87Y+Jv+8QV8f6imqR
cJnkGynjYZUB9x6xb08SO+IVePkhI3WpBai1p0FeJBDk0LI3v33USwTVhsuc5YIq
EF/9XpICe8fy/NDP4AeszF1J/lOp0MyClzSlpXrGTR9Y7eCvMcMaawB5qoQ9Z/Dv
QnRvmFGKGzYepbetLlNyoTh6eRm7YOugAuoJaf55v9XH4MSVC5potxCnvjfN5Cza
/i1MxT2A4bRgI3tDZYFIoOxa7EG0aSv0+4m6rF7NBX+KBqCe8Du9i4EdkeYMPnOJ
MgZ2+kFfL+L76f4Cqc2QwachcbJDYTLlrK5LvFKIAW3X4eps+4xud7kj10MA8JGI
Yi36LpBwc8raZaQEXzPl407ZNNcQSON8lGdxo5lWsauZHnIZi9+SMUp1x79pxE5s
FU00E7i1QaH4S0NeF+5JGkrZP4GNQNrGOrTzgZYhSS7oMH9Dr1yFc9NfJAV5Hv10
W9zzp7abK+j5+CAAH8949bC7U1ei6JTbpUqIqE3yRAs6+qcCL9RCNGCLsBKAbusx
C/YRyuT6iYrmJBKvgMdk3CfHPYJ52C4WyoCMlZHIkWRvjNIkkaJEmQntMIRwm9tx
5hxXuQhAVA8lUC5WsnIuzOQaoZBg/J8T8uJ75tfBIeTzIa+hvFddNPvP8STxVUHU
GjDbU5Jbyl32EuR8y2Xsd3bxxQ9aYrLkNRGV/Qh05jiM4m5pXE7YwrOSgsIOQfG3
Jlmoe45wVQRfAcyatW2zHOe3Zl0N0wNzaRESe8jU/zDnqm3fwJB6Ij9mOsPP0lRn
Ja09zIdUNo2kZt35Ru0gDlo4J4RLsHhBbDMkhUdDfxdzELcL+vK58hD5GWkE/C3g
bBvvqa819lEZqjlGIlrXSSXDadSnq/u3sgkl/I6TtTIwd4dovJZFgg2v8Yxrh1CA
xcDD9yStSFHHv5ladlZF1M//L2ksGX97HB4FReInG+oIVU8F+CL4QgvaTv9mCPlT
5TAOrWvFry1Yl392KoRr6szOZsmeoSoIWGM5+8qZAO/ZVIia8Aml/gVJQppyiBIK
+zV6CauCSlYXc+9S7byhi9yaXFluTZjC2E50Vit2FFVTkLIZzX4CcWKwc+671IiI
V7g2/q1WgDgkrgD8x/Z3aISmjjz6eT8Blc3HnO2zVgzofTWcy2gAuWvQbiGStwL7
zA054BWTbRmzDdWovj5KPWHWD9YHd1ReaLq+qcESn8RnMh/cBgxnI/vmyo3n9AFW
S3fyRbduxSx2TAamJImhTuNF7CdLVvO5bA5dq7kxj2eHB2L1lP8HgmubV1fkstio
H7L+kqVJH8/ciOWOc3pr7A/z6Pis4G033rw7nB2rjulJbjcTZK3c1bv9RVgIgauY
VdcoyzzH8LC40TP9TsSCiKzO6qNxRDI6TQgke15q7D59yg8/b3VFBHqOBDuldOhC
rmMSBcocJ8DnPbID2luUNJ7W8DfJokCY69JoQbsW4Q/nUAwRePwYUKr3fhUbLJ/6
aO//51LrkhDt92xW1CXGoo7WYkT5AvdaLf+KEFZEF1cL8/Mz58Fitq9kLp8G8vZg
cX/kDY0sAyLPDsRD+ghSoa0EBe+7hHlHQf1S9B+GVVm2r2QFQhSjiWyo9aCAG4DZ
dWDxOgVlnewCcn71aBdrDlpgyWlMglAdPK8qsbCRN4N4L3wSh7g3Fq42SVZXh1KV
m4iphjSzqkvr4+EJrINk497BBVNJsqxC+qh/1hc+QXGLTLfSVFi7FGP/8aS3QxRx
jUN+iQ9x4rEuePnEBjpFZHuSuXnLTRuosrW4Xqx7+6ySZuyNaUzm8cJqyHBCfJ4Y
aab/Q7HmYBYgLH2jMDD7nQ9m4ryB+aHw97LaYdtvcoUMSwts3DDdZzatP87ATkEd
v79Me9GGIMwvmCg3iSCl0BmN+ZSanSScCsfvBhuw4vEGLuUvouAc2Z+FSUhiHSH1
G6NcA4kOltjt1fgUNdZF63nVvWabZii5G72Kf+OPighG2thIZCkXBQ0erWPjOmNw
qEo8JfLZIfE4qYZMzWYOjmylIc3KruBYXjgsoc0FOjbERKhFUf7L1A7bYH9zso2N
aoFjbJJljWtnOjAbnuya96Ouk9KDmiJsk4274ShoqSAlRZBGI7sOLKG82Vpvzpm9
nM59+3oJj/p+4o7pGdiTax+bKjelrcgT0vuEfCDnP0P6zHnqs3+Y+TsPrTnCy5eY
eK6JOt9CA1gjLu2nDIQRGDZVKthPALILHOhurYTgvMYtsqbJK6Cy/vxroqHgTiCQ
nx7L5KnfMX/b8KktRDWM7s9/JkINrJURXLiNihyAHwkgVAYfsj9qB1X/YzlbhqBB
mIUejIe2riGdZOlK9zyGFvAywQVQZIqRamt7OlPVn0HOntetwfT+tsZE64RFfO65
UJVDssT3lT5dTXVtEdCP3U4T/T4hpXEbsUIPard9K0FtJvaonUCHCRkEMzqhxW7u
85mELAqWz9Q7rkmH7+AhePiOdmuKM1eLzk9KGzHvvKBKHtv41zA+Bb2cEIGsHpS8
hIXBg52mGvkChmeUl6cK6eaH2l2olGC7I9Lv8ksVH4tisiTXXwcfKIMpKkCplHYq
3d1Mo5LpMXVX04uGSdyqecs7fLedDXNk4mbfc7UjVt6yR5pZ3CqTy2eqWGiVxLmu
1PYk3PvSYqMQaf3Wnh8mlKQFPhdBh3jUN/ZPMjBMfPWdV7gZFJMd+SFLTEVbCYmU
zZfcK1j/MFiYPrmdOWaWW48yud/4oP249uZITAmFZ51lTAtRHQuHMO7hnBVuJLB6
qeIcvfaQ08WwGMxVl1xwJ1ePHpSrpGyJ00k+g7RrwR8rA9ONBz3rf+1Ue12eag/l
ZodU7GhKKV/cBF/6tzYiGFP3DwX4H3rMi0gKyWvNfdHlXfvdb1jopfeJ02Yfw1lW
Y8f7dGlVnJMRZF0/mOTgujGPoW/Vs4OilGsZjQvXeqoPIdUEcGKzyH1bj7qn9ygT
SKSrQd+UsqNYIMNFiHrAz4dVVmtoB12xqnt3xXdGVpuSmqLItLqbPU2MXEr7BnIh
o64wtPf3NEI+tZHFkMfa/w1rXy/U1KE3tZcQILHczTTBBRLhoNwfpVRohxlPpaBo
2ZcKlBWUbD5w3D9uXTMf2941dFV6RIejqSwWQ9Mk480JNfj5WSa5gvTJeLqvZyPO
beJ+XrMxvYVyKCzBvJ3bd/aFdf9znJGMOQtq/zdl3Tc8uQOlE1vRwv2SLWRcMnWp
AyYgP2QYnY7yaIhwk0z2SghBkUmlBLR7pFf7RHCJsfImrkM5y/jkhUidzCk8zcj3
ytii/a+vHt/UfelubP5yBQlWZni7GwWhQVPRDmV0nahFD8yRfAPfPtgk7uTCQsyt
F52yKKzk5JvawRBFYX68DoR1HUijdfg2UEarmolfMSeKk3UoRu2JLhnMjin/S1hS
Pvq93dELCKMtViEWf6kuNOmi/wtI7v2Yi6M9RiwYAq8x77Xifou1vJ5IjNt88512
aJfEMDqas/OHW1dngvoOhSv1Q6z3LSSzpQqIhMkWVhF4H12+morPltPJ6sRwIHNr
fenDYMFrf6pQ3XJUjH7deHfq/egt6N+Tt5/OuNvjeQMKI8JscQt+3PUHbkfxf0fz
VcVxl7Pc6RC8HU9OvrnF7gJLAnGKW/ARrmHnhSL06KvB56+3qd7Vro3+LCwh5eAM
V05DZrks+Vb8T7DhbfcFGtJ8No/k2+GtsZ23SfkKdf1TuM4yj5O+vuS2m4mquGgO
Draa+Pin5h9/AJaOdWZA7PsKUJBVvo8SEWZhdM3A9c+dgyKx4QqX+c87k3g51JZL
3i3+zlxWzSlAVjnPMNaw7hF6S6+kqQMSyqiXiH3r1TyKebG7nTWSqUgIDwq0yDJ4
Qsq6eaP71AlaihzexcVqRE7RceW7LqX7Pf8qk2FlNBFF9QsT9X9dOpHLkZz0n6gp
cgvy5QPoOEEr4dmPnybXOfPQ2crehjYobJHLhKC+QZ9Nn2tRYqzy6FTw8wBtbwTR
zjUd+jFWRI7w4X30WqVMSmBtkV1bfLAmEl7jhxuWcSo+3ZTwXZRKrhdbMOtg4xv0
qxIhL8LCao558TvYZrMJiDHaFAeS0g5czBC/p2XTPzApDSiuxUNPQBPh0yZR8pW/
OXNxwRxNC2T1agiF0wCnQVnPA49OtnWrP5GXD5wyLEtMHflFXvgG+/7Wb8y8LJgg
TC2+QK/zftl2/STiTkbgAjvgUBX1G/s+T22/MhI0jsDaOA+GRMUXA4Pgu6LqruNe
YI2x0adFWbeS+Adm8wPJCBTg+TTKOYqgeuZcLVOyRbzBvybSFWJe2p7UaPCMZ6JS
rVkm4D18TfyI0DtX5E5cWuPrY5/efm9CW7c8oX9DKVSCd2QJCRA5VDMO/jp00bp+
lG/l3hksxtL+HD7I4p0XMeqg7zuJAgz0DlFqH6fkajNDag6gsZOk4QGstyD9wfns
bXJELITbVb6nybr/a4+bB6S/+4fdwBBBxFMuVkLC6OR0lPgFozE2te0oyPKcz0NG
huM7HxuONGflDTVaWTrT/w5iOuYK8c5/0qz+jSVZ8+2kK+dy77w9FtocteHVL4TZ
1qz3z0VIqZ7cFja5OmxK0FnJDWDHBpE5HG3jB9fUfeTz33Rbv9zFY2g97+2xcar/
mAfDXhyQtoDhjYPBGlkf+f7Cf4f1h7aCF5Yo3I8oyJPqai56H7zJ8BySJqUHHrDI
3yvraccrbhdi59UJfVgJeGWQPekG6I1WpH6tXOd9mhCBItz0jqrUQxARS+d1nWFr
qSXrCf/0GM9aTTtzweaY648oRTZqs9VN65kZmx+nguelEDQPjmdPWiAT/cw8a4Ss
Du5Uo03ISE++v7uFizi/h1YbF4eTl7uUSsK0ZrPGoEfvjYwcbHuoDYrl+wfNcsQr
LDdoU1Jh30aFM6/CoFg9Zgs1IL3G5GeWE8UyDvFQe37rTzfNO2DhNG6TsKwuHK5Y
iptrNlIqtzLIZnENjbuNOf4FHiFfZVOO0mv0yRlNgihD6EvsNWQSoPj550DaT3+9
krKKIX2CnthGTyW82x82smuDfJeNLkPkwzCl9uNLNofaU3en5pEP5pP5CRTOH7g3
TztByOKSceFSnwvwTrYAlTK8UUCgYBK0suGk6BcIY75gEOjY5MIJOcIIGl0ppY55
+5+XjAptOGAuwMb0nFmpEIlHY07rMdEvbmg+sRubu/kl6K3gzEOVfugse9buIzOd
L6Qstmb/Jle1ayvbWw6KNbxiHGUI5SQuoOTXD2PhPoqLYc6i5hVzW4kejh2tCxed
AxeUTDNDkN213K1zyPLduvYdQ4J7Ov1PM/ijGFSa0YEw8FiNsx1hDoSCo0gowhZL
pBpsLeruWbXoyG9Gv+D4k9WES6+I8H2IJSUfC+FWXfUs4P+HEl7CqV8mMOL7maNZ
6x5HxAeCn4otPLf1sR/wFLRbAD/ePLPKlFU17W3Tv2W8KD066dZyAXxX1hkYB5xY
eNjqtBHQja84HIOQStlw42/WxN8Kh/5HmuCKUa8hKrotGcbgxrkf4aGyJhUlv/It
4YAhzLImAAuZ2h/LgcCvVbuv5mISAIGUf9gR8Cihnm5hKUCgpxkAmnDALmWQcnWN
bL7uwTw1I+hHgnrCRIXeWsaAblUUEs6md8mJJscqID1JSg48U3etJAzOo8BtSxJb
vbYFb9AbI0/KowR8ubzrWSzr52r6M+fKc3lD5x8Zt6TY68AVS9anZXhHCJE+pqQN
7piSAuM8UwWyYtJgQUyeekkAXLxTcQlFXVof2ymZPXQ8zP+/UG4krbFbYZjqAXA7
WgSTkflTiu55dRljRRr7RY9LCXOdPALRpHhvXY7wwpm+KBtUF6+GY7dr/KRlnRrh
zXoDN90OjkfL9j6lh6V0hDW/1pTz3eMXrwA26o4JxZC893B6qrNlmowzFhSVCpIX
xpFSogwgr4nUks/is/7ftcvHe87MitP4zlzquNIxpIr2vIKh419IvAoZtOLxuHIw
uKElf7FHxrQYuGUR28Tohm4kHTdMPgLj44l249mlP4lKTFDeScXvXlm6/ZpQTuUJ
cIgvDhn/NTgk/kJKtnQIwtFMdaxy3+vNv58uFwAl5jsO6QqlclBvA96sf2uLasrS
njJ0FCS5seg5CbXkSiG+HoulfXnwATPMVDqiN1dxz0nCJQrAZV/NqjSqZsJP74vr
IcOj157xJDh2FLpcJNbppr4ooFrN7qbt/tivNybMGBIU0WKZyBTLUOKz15pYZMir
1T52tjNLiu51Ga++lqBEMenEFTzteFvtMxpkWkMtl1eg5NyC/1IYhef+FRQ8vMFp
gczr8TydDLkhcZ2ZKOu/xCidXhqqP4WPxiJj5ArCKrKBRSuKwy/rFtu7gml4z0BL
tA9HWaqUM1y+w9JoS7mC4hgSSWIuRe1OXelV6BJRJwvdDEuJqkpKpm1yja2DnGRy
M0AytRsXS3FkQUlIh5kZfolG1+05oZMsyFzhiXcSCbV3wFVDRS1Ypb8Bs5ARzgZ7
VG6fu+dSIgYjRInT2EGhRASeSLGW/nURiGgRDyV6bCMSnT8YBzn66up2tIJ1Et7L
JCQvemyLQ9TFIr8d4HAIKO6Wgbu0eillZRU/ge3tSwtH3ReyUYGuYK9pLj+fQuG5
vgijY7KRjDvEORD20/6usKS1y5Txrz4V6GmHb2z8GS2ZR4SgdPzWrmM+0CGozyKr
2+Ofu/ULOtYtPhnlc4RSL62TLX05y3FoBfMktyE8pQgH7cV6DWgBpdebKCu+6hNp
0yTjF29Dv0BSEtalSPsRTEx9olJgFtItPmW5nJQWGK361HecLYBiRmxdAW4uYgLc
4sIOTH+kVZYw3lOxZ6bplrMLti8xzta6V8ne5JSFs0e9pJgHDZoRPe0LdPdkTrGS
iIK/tNvRrQlbFBoznOiBONnc8xpboZHU7obDx0xZ75N3n9rGqe5puQz4zBQqWf/f
L3wd0AaVDrRXbKao0X3c0ZL0D0NZKt5rAGms7H/yNubMyit98fOdghsqfTwqGpeZ
8cdbjQpFNYNi5K0AhV56iCyPkO2s3JAc1kWF7wjyUg6oUmVEqQHt44evBnu4G4t5
s93dxPN6C15JW38GGhX1IQRd/+HbP5COY0Btf64DiihJadxiHBarqZfkgZdKzCYt
THdn2RC90XMDqCuv98l+6YiZqKbi6I9ksr4Ma789pM9q97u6T1ltxLyS8erPriH9
tFgCPHBN1truzlUsVDFhbCoLyHiCx9iwWcWB4skQ7zOfkfV1vZrwwIrE+Leu4iv7
gu7ZV3He49+OfZSGOHOMzZfF3P4gEf3FcYZAltTair8H9CR+ZtQVwVfSIZ86W581
nQJUZ54u7eaJVPJosOeTigKm5Xh0BO89t+hroPEnoQF9ODRS0bLWw8kg8wvw0nTh
U5KiIOvZxtNnHHQUELA+LEuuDm93/QtQwY6CGv8boIr2b7c0HFFftWluJL83cy2K
xTiiGp/42Y3Avw4WL4bsKoJ3k53kIWAVkrnUPFhyAvc+hIT3ddUhnDu3lWCnRat6
umIRwSiAw0j/V6IKsSmiYDafflxQqjMUF6K1BXgAPDoS4gltuPfxU+McWCFAp/Z+
1U0az0UIXlPeS8xWQMEZ7Sapmfvq2BXJ5POe9cm8nsgysRdpvwN9pMJJTD9j4vPQ
JUDo0R772aioRWk7p6WlsI3hjeKEn11XB4UWd/UH2WzA/5ZlTssqV0fQb/6nHi4u
GOjcoHUgfqbtMN9EKRwXWv/TYk+KT8d/8xWHOAuCrssKMSyruumQnY66H+NifItH
DU7p8ZpfqKJyTbMYWQ1tG7n5lIfE+Na/v2XAP8CSc1zsN8WtpLCid4HMbddE9Ojn
O1MhoFiHGSPQ+qpr5s3/DGBOqJkiE7at7p7Lv6PfAZj5FlR/FtQ+YvD7YZUxMDp5
k2LMbqloTwGKgSVLpqf7QRkH70y5MYpxKS1mtAjGCnRFvacANkx6CEvRCQJZLAm2
c2UUKSwu9BJWDRs3ffbsR6kQKxvJU1U/vOU1z+p98vTUGhcqMLlfNasDzK4sGmC0
eCsbyFk5rKQ5HX5Xitwj7UIAhhCjcfIL1se0SwDNLSiDceLzARWDvruABcZyMBeJ
e79g1PblIp8vhCw3DshGC1UAllj4IayJacjMv6KLQrTovX0Ap7w3GqXWCIjsDBdH
wbEuw18lBzWaTxzLwB+7R6m6GUcgV1hM3SppVXJX8BxnzdxfR2vWB8eQSVUaKQvn
pXnjqSvsGdsSxlGI3e7chh/vk/XviNKvrHT47LHBuHmOkGPb/dS/+Dq3N+jGPUCj
77FjIb25bPTV63P2A5LMi99HiGGISlFKh9CE/OsKlVkkpk7siyzzszz/3R8f9bIp
M6DPrthjn0klEgY17xB8YCt+pgZSs1br/KOVqC75AuyyLGrmQFWNIK+WNHxCDyPP
IdT0nK98ayHjq7TpkZB6mwK3sCx+0gBF16ll5YUaJowd0I+vVgKrfurctCvUBa7t
IzhzrZ5/uWzOBeGS9BWgyZzbUo360s8P2j9k8iSnG6c2e8FVM17kTweKKVt+oGc2
9lSfQ68XzBbNuAyPRe3Qj5CS6/vI6yqArg7r560llqdBz7KC1lsNAzATLsvf4+2K
Ia3xIi6iau5QYWTOn6YFI/TzTie0yr9boAlW8ho3MmLstJ5mHJkYDJVUOl1ZcsYp
IZNbUO6tZYdaKZPRXQqFs/FRH0vhKQUs1JmkrVIem5/wbV9TJ6LiR93iREWv5kMa
juw7tuYsaRQnuywonAVCvFkymTEM9EGAeLqogkgJfTYulu04olvMZGIK6jg00k/k
kBp62j/Mqnu6lLD9l0UNUCmFyfjG5v5YllYchhzmOL7miDZsayPNpE2WYUP5L/kw
q2A/lYuYbBUKMMfBxA/5Lvjb9bxLxzArtTx5LAZuAf7aW/AK1lw5W9yrhAey/ye4
h5xc6sMxZdz+TD8r3R+5+Iauj6iB/BrDBBCHJVqkbxBLkVMc0uoxa2bb/DSBewJJ
dcZOrhC0/GzdBq6TFdJRxwvfbPwtYJnJ8x/0Z7seIQt24boq96/uwgHLcFMknMGA
URkhj958h+qRYUan+sCwFr3ZzHm+YeayJxsdHlWpRI/Z6HhbglNpdhjff/SsHnmq
EGNdE9AugGci+olrOzXbk3g4NIFGoJIXECzTlnaffsdj9OUFNIltWkP5c3yF2ovi
R7BsOAUi7wgjRMYQ4ci5y/CbgsMbZrCnUm3jt83Nggd9LLD7TTdk51clEVm/DwgQ
cwGrQRTxYVJIoOzsGRULcTgBDVVmxnl/4hQD45+DGdrt0vtmMynt7I36StSDRtWJ
u27P+wIelHlldoKW/LNFYlZpZi5agEs4nAzkWBc4m6Key1iqe6TNJH+B4IahwAWS
dF/ZB6kXJWUSPh+Wzcjl2El5TveIAi4O2WK8Nm4VyRIFFFk1sgMNcIg9S1RnKuEd
WUAC0svh8tD16Och+b0KDmtRPkduTwPzakEtRXEsZshKXS9H6hPskCGL4MndyYv3
6f4+2DrKbNhnIVcc20fRrjWTwEWcOw40nT8WNOb+eOtUkxFwEM9l2GqaVKgHkMzY
uq9jSYEsWf/+hnBZlYFE0OV2T18Lk8C5XmAaaXycpCTYuh75PgPtXOQLvLkK+sbG
Vlov4Oxe5wUEyon29QUN+EBobjDFoZxQ0NAnxVq7+FfzLPOXa7XgSyb9JlkEQQrb
4G5/DyWtDeAcVQkdbz98ljSRq2u1VNCX2gI4JgsTKFShK6s+PV/UwLKfu+TWCx6m
NfripOlZnVI48+Z208o53+2jimdDugtG4KUAC0GOAyuan2hu0hn2shU1W4TEvChO
UR9RojrVuVCLbx2tuVAGO5YBLFmHQgRC6KdPZYG3B9nPYuZqQKzIMT14a4ubL7LQ
DI40o6fpcOxQWrJ9wmRbQdFtRteMgESGA2QSodD9MwmowDZS5bh2f5NntOnVBQY+
l7FGbYqmYDRZVET3JfQaIqdPpdtvzbCfdEML3X2kU214gAZnpnnEHvp8koXCP+ZV
clFnTz241WZPFmrZEeqk4ja/a+fMGxIoeif0nJv9U1x+4uoJgVlneHS9YgdTG9Aq
DgQ88UML49IpKGq7QJouq32FfAV/lGWAx4flwd9IzLrrXJV5BmNHZ+gOsHm8CwGS
xkSzmAOylnsQUPe8Chp+aOQ2A1l9L/wtKtGnLMwd978TuPobbIk/WME3x2L+1g9w
Lu9wyeBbvruFJyP/U2UuEBRidgwS+QKhrGaut7phLy13e90M6wg1KUDDCkxYmU/q
ku6/tJcpwbTsydBUEBHgAOjm1AhKCZSY8Qowh8iw+6J95ShdazPvGMGxK/bLJs+e
BmtyzqduFrcdgyToNhnAX/xxgu7OPth+UoXpOOoRqrJSnuBYXVaytWEAGo1r/+n8
jBPMrS0YI70EbjB4z6186rm6mUBLqD8ZmGnTN3EukLq/dpgiXJqkSnJDBykHESZj
cVatmM7ZbgFXNQ33z6ConZjCY36stBMFd9VDcP/rMttP8rOiFXjuTTerJoE+EN8S
sxGBKN1d44WR2cifzzlrufMCmWIvUr4lCHRsHE9mNQfbIfKdQJZMm1C1bmXVQ3Pm
Jr2dJ4CVO7IaT9x4KFACl8a/DR8VcIJcGSzNRFNO7duvQmrS9XIuiqstYFBlCrA0
n9YcRL5dltKB2X1LqLNunw0C7lXhejpMIPBDt94k8F2gAHJ+TMHudZ2gw+Y3WmqZ
zTNDq5NYtfwCYlUyvcogfSRBrW8cEpqMvCdvRJFAKJML//2VNRJyfDYnNjdHjeBe
RsIIdx1bhUu3Ahi4lzibH2TKbgVFJPqEn4efTvgQlesv4XOtd2zwTlN6OmSUyuKb
Su9HhmM5g8OFr+LsrcU6njp+lqDPgL9Wjv3EndOQ/LrdnYbbkle6MY4y/SoxLW1c
lNsmojZz9Bv0FSugATACdGtIHhBaOqbZHFLV4kexYUk6AfN68Tic82jqvkPxdhoI
aHSLsAbmRD566CGnf8VCpwnokATG80LBC74WFSbXd6WBzMgfkGekerJ4io7zH7mX
0l3w4kFu83+J3cJB5tDBjDGZOwxrpgrPBBYR8DOpgwdKKM8pNq8oHqFiZwz0+ib5
WJ9Q1w2d2c4jGmTNrfp4Qu3iORMNtcOV6DJm4XPAio+plK8AOujtk9YOlunJJlSd
wNtllZKMjdWjSnQGc9xHDpup3viugz5V+p3CPKQqBgWxWb1fWuLObHgq9R0FLHJ1
dVFwmGEnFY99agNtredaVWJot8XlG+56I46Akbgk9ZuEvF3wPIgsha7kJ+cnhdx0
FEvF8UkXR/2JFabtMnREn86IjCbbDn7ZR2jJWRm+9llmjd0ZtPIlQEi7im+BB+KJ
G/n5O3oLbcMYkedQNiuQlnblY3zi3TxrmDrfjQop31iNgTjeNGdLunaE79bGBNep
fF5Bl5yb3nG4AbExjU2SnMXFkF4Mwub1f6lLs+saFYKow11KpZvel9QuahNnFtpz
QnKNAxyBIGi85iThweEyJAJvaP/yKpyRjPNrPs7yFhWmBlEvcrmQrRDsKq0B/en7
LkuhWr2ngrdgKFmCMG3WCytUJ1+5gG335ZELG3Dkl7ifllm74z+eG3PGkVJG5kZB
01dWMOl/VBvGdGIkFSXItj3vU3aoI8xsmMx7b6IQU3Zd9dxKD64XLAgvShZ7zVA7
TMKNpMzjHQYuRMO/HP55bEiv6wjJ9TkMXr7u8bnN3TFpf3bohU4q1BK+l3a7xu8P
85FyFjYuqbAe7IBhyrI1+K977EoH6Bb3a5NUTQa3HueIZnqQ04FrgJjHKyT+bFRr
VoRmlktl506RzSxHsoWNfySupSxT3LBr1m6nQZWS/RSkHK43+FtKQ79F6zpDrxfx
HFW9KFFBpFbFpx78F/SXIs5h41diRnW4osfGQ0IPrKxDEnHcZwD5u/4JdG97WsxY
36slNWDVkSVDnrQhgesscY14c2FxBY+YxXJ6nYVyXexa4YyW3JqFG5BoPoDUQeOZ
OCTyejKmF7S8fuHudstuU9zyIpNOv50/46qVogynTY+18mkUByiEiOK3qYIc91sS
effPB8WHtQPXbC1CkzQl3TAh70Lu2ebiFZ/iIs5rYEX0jb9MXgeaimUFbqUROShW
PCFqAeGOoXJc1fH2enPnMkwX46Skg/uNkszfaeTTf9Uu9moqSGlrjl0YVr+8GCtc
9ExggXs/3M6qX/oRp38COsmf2zxsNhEA7RXifV2W8L94mC1kqN8cEVmyYzU86Yev
ozZMbl8YF+OJKyDP4nBQZiaUEZsGL4pJMGaPLfYK3RCjRa9796O7csjZJPz0Kw8l
`pragma protect end_protected
