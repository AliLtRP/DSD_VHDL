// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:31:29 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
L8DYZ5TmsCQWMwz4OJ2lotVAZMaoNGa/ULfpDNQjOYmLt2POwTQU8qDJmioN+JJH
1y1+yq8dq9H3/0ojixR1VLFRXRjzX8Tg4Y7Ivw0VcIhFEm3xcEchizbHFBoS3lwb
CRXe6JX4TnR9OEKwqJWeFrlQOJJPJY+pgEQUprU3+Ys=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 62416)
xaklISGuHDLPAnAac+wrPENtKj/MEIQjHJcZGUhioaC562xt5Vui0E8kT8EOlS0T
hVsYsoY/Eji2WgNkmW+Bxr6Rdd2tRadi3//1aqiAekEYCg5zYhpwU7DaKi6u/Tft
lYNHhiGWYJF001f2kHTVWpTfX02kPHmUACWIIwagfDTWA35T9SninDW+IAoqzXJz
gdxaAj4P6W8HEOlbrPvNQUz0xI2p4p0Mt4boZQzMP+Vl1v/mxAIc7hFVIEQ8WkjJ
ARlrnuKa+n25/QljvEsQRNndWmzUvqtKz1tYY1CTU1OjmTK/mdTwMx2wRmtyymXS
2QrmV4MWnr+HCGvOEgg4d4HRR2qTsbIactry9CPumQmBVXfqkGubIAGqGFMaV2D9
pOIBFdtahPWK2a+Hpjyt1MD0i4+22WRLHfHeuR9hWtV8mL0agtvAsp5FxRvysT5I
cOi+LfaTO+yIR2m3yf+KL19m5CxAq6ya9DXp7c7QwWFjYwU4d1YqNMhKFCQymL2y
Z0bz0UqCCQfuZiBdIy00Rc0+Wgifn1szYG/8kkrGXi5Vws1Y4pfW2xVZ93AMSJ3W
I6VRZFzc5ImzRKs0NvY2gfUUjrAf4gipKGj/Ilya4pzNPkouk8VLr74GTVDfTgkS
wmTAi6gg5btpH78Oytaj0vTXbddZ6sZY6VGfjk9eS2oRgVx5Twi3HhUqFkctZXog
zWE6vZxT70aQjSP7zuRKuMgRnnetO13gBkBJRZQeH9qNWDr7ESXUEm5zfIGD4yEd
U/SpBY5+iTawDQVlfMOxVMKfA5sEtcwFGQDO7pRdXhExtbgcZ6qe2dTgs7cJZ6u9
V4yESMFRvD0NMrzD81g9xunCchIwjkxyAsm5CFV8T6XaufehqNtyZVANaFuVpQ1s
lkYpidO7ksifQ3NFrx6YqxZSXCPGI3PYQLYJcOoYtYMebur/Fk3CJuqLngXv/3o6
FFdhMbjjEGsghfjMzbMHHgGEhGSSchJEx49qeQuzTeb1pp2dUwV8lwElnNCuUmx8
pyOYuG1xQEbfeNrotSQHazdKv/ntZbPvM9FtEvGYs0rurB744EImfd8crFrRkncf
KlthcsO/8WdQk1KN3akv1k7Qh9ZgnTPDTPiPEy2ydLeta/X/kHh+YfFl80h2PPXY
20m8WfyrDvrBfrCY7u60iXhBt9BJ5N8xph4mG1AdCTAYaXbmIvrFYh+2vcgnwRJM
kx7SqKWTo3ba8xLuavXQLoL6Ib1PrW3ls/kWZSKihhgfphs/7ZaKoRc1pANuL0hh
pmeKaPn9RB3WkjDvuGktIZpxvZgLSX4JEiuyjLXKNXQJtKsVCyZFh2e4cuD20gP7
GhVX9WALo+v996WJKI5HBtO5UEbdOsc4pXUs5ENn8tScpBkVxreIWGAglvWPyTfW
NRcMSLQfqnYwOkmH/lUbctNodZ5TuDfpk3/aBxrd51n3QStTtl+FM0XRs9gOLsgL
orGRFKcsfQ5QR+XUY4kOU3d0HJDfDODiz2bP6UnocVwNHVnRNp84Jn5TeBTXceJk
b3fgx8BuWJbtVtn4SiwhYW0zWuU73R+SS/pTpMFnhP7D/9hh6f4HGFKWUZsx2PHj
1g6lec7CzTlO+RdVD69xhmXHGKunHqlorQbWfLFpv5AunIE5k+6/MK9KYF0gMnc5
xlFVcj868YspF6ntMtSm7jDr38IxAeJVM2bYMsTTgJ54tYrYkMCR4B/S0VhkwbFb
wRq61r5YSaXT5t7TDaE8yOjTbFCbpPIE+SF9ojJrWaKxQmQjjByeeIcgV8Rm6XIw
3CNxH2TDN579dZTZYL+xWe89FwQ5lbSoZdCtO1z/8SxzSiL7M2F6EzDVlJQAlhbm
VCKLWEOvaw4rZdnjcdnOW7lRGJxJtdjg3//mi/BERq89qBUlgOsPhkx+BTyCFr9i
hAkWoIVxv0CB7cAigwcVnOeo7P3y6RQ52l0WPeM4j/YMYgOU5BqM8GMbVkem+yjs
Im/a0qgP1k6qhT7wfVeAOTuNdtYYMLh9Zc6IM5vJlmES3rUpeHxGOOGwhTCtO6uN
2+2RA5EeilkYqP0sZ+bNeuIedRz/kVMQVj1R4TWy2y7Xo9hKPi3wHyO84rrv/TCf
av34r+ZB9hRD52fzHwPGKAXpbdgW+DUJEenSPQQXbfET6x7aVgUWKYD2CYBkMfgw
ZcvVnhP1g3OhXPuWesVDpoqiYT6XfrxrHl812hXKpf1sJmfFU9GrT6VhaD78SoX9
H/RN2pC4AnzxvFc01mQYukj8SJ8/PPA9hqARq2lQ7yV2IlR/CK60MueYSoL9dNbi
0oXCOoJT1HAaeXr1tzx9Pis4ar5i86/oA40ueSVRuA9s7CE2zDLQnbu2PrZEh+cp
MIeWiXKUvpBHc5adM81VpIE5Lrr6HdVJuPPkANBCWtrQi71z0E74czcOrVq3v8Kb
+zcF58V0OvX20F3oaQeO42aPAMuS75eRWponWHjeUberLTSYp5PT5GMTVkNOcLJc
Q93YTXAUsd8aq9p5hjiHZ7zWzY1Aq47IbrMJoL6UsbdUQyfDPKjxPQl4eHfiAoPS
35E3pNgJNBy5s4wexmINeZE3cdPFVcoxPlldf18UsHrMiFzsSi+gLasfnk06NZaE
rwgkg5OhVpXVrsj4Ql0OUeqR51vRcB74VHagG/ORc4y42OcS3F3epcp8zGfEutQ3
Ja2WvWI5R7+My9IjtDAb3NA0nnvheCLKqAY8fMZXjCUL8Fr/8Yidi0F1GCBqr6YX
61G53rinURA3MonMVleo2zciHGzxSNeaoiCj0T2UdSb2KDEhCTyhEYaPnqvWNcSq
1wj0jACIJKjb+E00EZza8ggkv01/gEPkj/t64H86nSUewcOFgpvFI6Y6SLN+2BhN
ls+tvy2XHPdybCKqG7hVoVfc7qpvEIYShpTKTDmCcf7uKqvWBo0q1wPeZgu0rPBz
kLGghMHgoLL1w9zySbKCSB40gj8Fx33So6S+koMbcpig5IE4nbVRxPaTzzdGyPVq
WKJ/pw/f7/Wl/AyDO2R/oCTljVkLn0fy3HO7qhMUSH9TMSOsMmh68ESmM7U+jC0j
46rEzr8hCnfMhdsFnPWadK2m34zcx+3LI3XzDl+aTdJNxi2OHqrWC+xS6Oh8FsXB
9Fo59kADt76SJg7LRbIlC1lCS4UhR4SS0Mcd9+GSOxcEypSRfPe3TR9Eibh9CISb
J+CLT6XXC1tFGdv4B2NQAc66Bacu1jDXH4yap7wn0jmb9bStmZ0G9e980As1cJUf
k3RGCZGOmVy9mr0twj9BJb9YYeWSJltIUyEe/KJY9SSAg2EhhvbUerZq+WFmN+Sf
RfbQJAUOgnbjysYDJjswKR1aFjIYNkfUmgcRs+MrQO8Kcnz1hPr6lnx2VOB0ZPHX
PeBgejY1G4+qmaUVhSXZy0JmrxZqr1MuyQo2Xm5ny74t3AGe9mQa+btah6TNypYJ
qFLqprbEiFAVm4VRGeJFN75efgV8V0pLABWEAY0/8RH8JoHp13d+mm5+x1NSoh0g
yKOKX2PIKryU+bfvTZS/g6QDVEkkAFtos7mXAMofiACb+zXEmW+6QleW46RH7WVF
Um+91Ta8h04lOX4MCbjIcLENnjDephCKd6YNpY7EhgHLqL5Vcpp19iuT/UX2aDYK
YeY/z/N+dZPOtjlVtBA7quw9YVbkdg7oFDSmHw5ctN13xWJf8yJY4gDvODhti7o6
UgbK/yNwZHqIcWuWyDsAV92p+zArMckXjR+jv3Amr2u5USY27l8oVBoHu3ccfuMg
gKF2qcVRojGg4N3rKtUDkeVDyl3D8h4NvP0BPf3xiHPbrI+hBSCykK2kdUNekk5O
D/kcixqRO7/maGwqT42qiQhnpuepkDpQ0Oyog985FlMB3YrlwERcANIaNb4jNVJ2
AuYPFJehJHQV6g7f+dqsuASoIVvH4DOUdgM1J9+thwl3lX1CZfO3aQpicfKV3DzQ
PV9t8kH0m7FN2br81WhIFfDcW+LdGdnDVjux6hUv3KvDGm87Fmkbz1HAID4ic6Hf
1B7A/bG9QenFLzFgVu1169Fz0lcGxF0jSduAzT5jhxAM88Nax7nE44nnPa/aVo7A
o0NHV1rC1qFdRHLEsFJ4Val1NSfFQB3EmfOBezAfXCBPV1z4DgV4SU65nQcbMJkX
1aH0pLmvp4NDD+pXNneg1QBGe8JRZX0nJ1/PUnymmtGF9hAOjh0igR1ABZOOydky
KCXL0RL8MLhMNUuMbPlAv11gVVNEjzAdaZrZmbGwfiMUMOzeqQ95Rn9TH5H+dQSJ
2A01oeKKUesU5/dH3IUBR2ARiiFNK4daNI22qYY8e0i+VAlMdvLoDfq/91OjwC0i
aeH8vb4liXrb801Ti23yczF3LBA8517h8Hu8vLdv8nxrm689Hnqgyth+SLNC4ycY
HZiwRZ1sUkf6EKPcSeoz0FQEMvYNuc//Kpk135hA5l9u9SZE/4A5c0CmJFz7eeqY
Xrw6AXbHZGk9HHBC92aQIDlbKNYce+Qab/JiDJqoSofoulxTZdsPeSbncwYUWb/3
RJlWmzDFm/vNyYo0WdD1f5wuB45SeigHnMiDu4vg/S/5EhnVf3cLiSbkF2NWAJUT
xzXDoAer+jjrYSppMys3hSKVp1xa12tlhKZ/6mr2hhG9cXZDccriUj5CFjC6PZ6r
7mF8Qw78DgnO04Or/Iam6/32e9FFBy6OBLUZtpaF2n71PsAomQLFWMtu2PCPx5Zv
D/Q3zdhdrGyqJPA7a1/i5FkzZDX8U6PlT44I88xHLBuKTq/g3Lt8vkVcwZ61s4tR
e60c2ctqJxFXPJ9z2/qIn6NtuxDV+yxJEwxmOmkr3lwtNzfRlGHKZ3+NVo17gk4D
PA1XuNZcH/CkRTckWCr6LAa851VuENf6BeJ3SwcPKFaBfhOxHe90q9EqN3N6wGm1
ZusXwsYrOfRr6B/klJM4xiZwmmsK4fx5gaBRgiqzGTFC4VCCWcqOs1YNN1L3xX9K
ATP8IyqlVw5Ng1LqyqMfamTQSdmydU2DTTWAouTXZJEZcBCLhSusQMC27fIHf1e4
1UuCTqrRTx8bn0KjDoAbJl1MLXfEgOr+bmkhlFW0Yq+HWk5czhevWJn3W2QACHcD
nR3rpW7wTKRhsNAAPHYmnhJnyx0M7wQyhgnEdd66OGB4XQl0TYPqtxsI43cZENsO
JUrJGfJqnki8tkW8IAqZbzO8vNpL6LqSHeVd8wVAcSaF3jtKXmIwt5XmLySnNSxC
uO9adrM0qFaLZ4IsLN7Xug7U5k8v9AI1tprOBnIgmj+VtAe//ueqEx96cPwqtnVJ
recQqT/bcvDRWFfkljreqZJLHBD3cGUVefeQOf2lXS4ewYOd5fPfiOXMvo2XrITT
5x7R/6GQXGvdGQjIkCi6oLzQDvRElOAmcwtqW4Am0YudLSYbuHx5WqqiloqV6oqs
TEmthm/3c2yne9+wC4Qb2zQ62cpGFEQeohHhA3CVSn5gxBoOij/Fcd/MzTeKwBal
vBvF7pjk2SYWrj47/8HcMwHGBDTWHhchVLUUVZczg77jEXJHdDps8BnACyT0LfC4
yh+Li/nlOgYS5M5MAdHB7Qs+7WYyhPrRpfFGiZntAe5yHUIB3uE0wfN8c1i60WWq
/khEoEW9qT/JBempJ4PLltn7AtStR/lOZKmBBWi5Z2XmAIhPFWF9HFku7w1k8ADf
ekNw9vOZD+CLW/gYihrcDZI9tPbYyTHaUYCqvnyrGC2AoLerSj/mf0oqUvr5fROf
FcAzuVvhgwRiCMjsYXgCbG2Y1mvmb6IO8ZmGIJ9MVQ1VnMgFKlzkQvs8qY48gS4U
/jApGe2ov9eSMENIXpIwOdp9y+izNAsEs3NGRHoc1T6jaB5vEAa1F1CxhwClhgtQ
9eWwk330udTN3oiqYcNVci6VwdwqmIHfAvDBf/tH8qjhfDvBUrRhqUh7DmrVQDvO
SGQBX35JXBLzllhjnp6R2SmL/x2yH6/C+WxnxClhRYaqbbTv1nrFe3NjcF4ysJuC
iiJezttULKU4PmWRQdR1bbHZELgnfWeTVEujs0id+lH2ildTkG8ezvEmtLPh8Tyd
E5ys5SWmwasL2WDAeLLQDwjERgRIFIu8nN0KXgexP6NmYxIDy2Qqslmt4+xdxYe3
URx7WH+K9MiyLN0Uk46dvdtZg4jsLNOHNjnm205/5MU+OsywUnbAybgvWZiRCaHR
2yHCZojbNqJe5hNL6FSq5d1nj0+pqc6iD0lM38jjpvuLhZ7ZZ1qa9H4aaZ3jqpsm
khycQC0TEnPQ+3M0AEpBgduN4McD0QLh8d+dtQEr9cB/PugePJyfzwQtn9DTK2B9
enI4qW/R08dErl2qvjIpaYRnlt9f8Xh9uMI/1kOm65UIb+s9bxIjaNWVj/TJ0ei3
F/15WCudUeijIjvh+6Ug4LrxtaH3lWowM7XNccT6vvn7CP0IZlhMlTXT9R2mF1qt
tcrbceW79y5XSWMpTpfcbKK6W0GUUmxI5rX8UjY5FDfSdLsZwT2EWKeZvbSTYg8N
ObPCH+A4KWCDsuYL0mQ2dHwN195D7barrEmE57ddUgmtNPFwP4gQmEyihLJ4anBa
O/wvovL5Vyng5bc/fruj0bbOPynRHHTBWU+s4Qwm9lu0tuMZUoELjCloFTmtLcmd
LCpaYexXLAnXz+HSOrVbt/EshJs6jrZm+wkvGtj0mC6JHLPtrP5ixFKtOTQbH5k9
rplMTm1YRw8sq2whefxQN5JQKhGZrjHZjjNdSWphEHOBwOKJ7TBZZ0sWB53jbttf
E5Pf3ttcpg/tJobfcW0IUR0CX4Ep6abp54inIlLjIzk5WmpAZjJbM8fGHyLPJKrE
QIg+psBDKyOE58z7qjq6bGsrRPvAwVqtrSCNoKG55EWodkc3k98EtP9nNgGmTQui
vBdxvESFzfKEoNe+bPqGTuHgtp5o4dZWHplf/FQ0rkmJYidWHbUMwacBfCVAyuHq
gBWkA4TJLwM3XuRt0ZF3gtv/SKZL91bdN43i/dqmSQ0NoZsjqT/TdCtT+wFk6rrX
/5W19RwCksv/OsO57638qPsEUOUsZOhH88wnanxorCIz6JOUqDi94ldSfEsEtzMG
NUObvfAFB43aKwXNyrt1Pf+1pRQJaJB81ha0hw0273/JURV9t60svrUR7OuIZa+Y
5kzOPAaB70ib/wgeYgGLdNUkgEo7cDS2KdQgpnHjAWQgIxXqBXsumBlm8QMYm7Rj
EBFynJ1Vjc0yyrvcERa+23CAL+OLEW5DDBCgsR8gJdKTwHvZ/MUI13Wn9j2CZ7ED
Ujs1iNDkGCrbSAM8cLHawC3xgFLuL8wrU2wM4YUQMAzFPsRxPT/okB22WJ85QdIa
2PL5urG/uNFROm31G8jvpOGYc6UTWoB14r6ACo9kbgE1UjBBYlMMQhsUbGW6ox4U
2xZIj2NTsKnwZ0YVOw2ti4ycXNoliJDzSZIBCm8C3h07iQcam8pacUtvjWZ3txPI
/euxNQdzHaySGkPrhYrq9PUyRSFccrJD0XaympS8qv8NMuOOkLTSacFkK7KVZGWV
sxCWiiNgSGPraCtcvJP8bwzr41b7NStMe+0eDiHwbJDSc8CUgOnB/geMINLFhCpW
sN2TNa8+wKE+v+FNX/fve2u4Ar3b/GgEtztTSIjG7zD1CUDs5wRvQqLXhUEeheEx
uJ+XMXE2QIyLEjJZU0t9P+FCZ8oMPGiQedDw8alBsufU9LS3J3cP/ebrzfASjPIS
VkOahbH92DUPkV4I0ec0Z9xJHaOJJ6lL7bTJ75RCFCCRuKcds+v2yZgs/LnxtmZY
fxY6KcVPd/y3E3x8fIKczsh0Ltc2CxDnOc/kEYtBi6/BetZJCkpYrrs4Jxf85hlT
WYjKcAXHbFRJVMgxTappgh5r40kXvca6ul7pRh4UZIro6k4ER9J5nV3yQk08vdBC
pBH/wtlmXE7J5zvmCR3EFZ9xCG3/XUMShcxlJqnaQf2zOn1nsprzW39FMGw785/u
H7+tWfcTZ0L2jm6i6sxnZ3F1cjCjIPIOHaeM1PiQ8vYVjk+KEfLUo/DdPVv+k8n+
pYfpMmR/s7ltzMFXgGsoSlub3jLWBDmlZ9AKWRiPOdbfrWbCDFmk/sSkCsYCCKY2
s6mhQ3SeO6darTIS+DdOKXQIQxN83K545uuMhBOdVEd/3RZ6bpzLTK8h7VEYmX0d
xKAWOsdFHKrHuUCr/gpooE9DqKdwAFY2xmtujm7zMsonThqNp1LkhHRmhxewzzg7
uLbAofaSZhXXS6K2cwzFJiVp1ddmYhINCxyOF3sNJvIql1b0pl+wqBPu1zXK4O1u
RWuZX5QLquZNWaJ47/QlU0HdPIoxeGLgao2nbPjT7KRRfO2F/pprdrjQyWqUOvEY
ckyR90bPYWneitWwu16/8YPYuinNt8t4nOcxKTBFbQzhDVkjj9Jh4vIKGdmwcfFX
RNJgRy3kJo43EEjbb9mUwCr6xycKHLokKq2UCNlyKddNwcy9q4y+GEC+CcYu8j68
llhAuWX5weLRNo5mWk3LIqsB6l/bE4Rk3RxmT2zsgkMqn7+IIYTMIGQqjCZCn8Pc
4CfSeiQ1dyuORKE26tlcgcud1J9cFp7pOFNb3F9IILlHKoEepNi/fqe85cNxoM9e
GBFsOi0nc7xV6TGbPYrTjC19miFkBuvPzaOSdWEZV2EVY8p2O/spcMlrovpnkoUC
8elfcCFGLsgvw5wwmIfPEpJHNrBOO/jUfsMLpSP0+dZaNk3MszEU92mSVh9+3yX6
MTBskgiQMDgjJwVhpaPBEILr8KF5tuS5P6FEicG94x288btDfiw/uzxVncVxmJWJ
5w3pp0WFfZ8hHVxyC+DOixm5rJmrahpRLWORuxTRfwaDc0piF9FHWX3DCBD4Knhh
wTKGtybdYAe+E5FvBjgGEGSsPktnmVhKm8wrUvVIBldE0e9IPRRgwWLOiZFZZUJq
VWQLP0bI8umM4ucqmjo7d0RanY3B1Zf5hQ6AUa9g2HaKOpu5VyL87YqqS7efH7z5
+tsCLZnLSkdKnzv+zIL4ldygYFTXlVX036mfR8aPgjMaVA+X94Q7gTsZDAS+ovOk
M2sIhY4NkbLsU8WtmhtrIyYZ/E3K0U8lwX6VvxRB5qHRl3hcHqgxG44hktVnN+pp
rjYnLHFt5qWIuEvLQktJZ1sRkuR7kc5rwbLyrqd1fhrgl0NPrkWzv37B9AXNuBpt
b0iaVLiiIHsBUdqmdqXYUE49lknsVXOSFlhCtSwLqXKRDQeh1JvaEj6mSemMJA0Z
XnA6BF5m16uvvQuuH+7yk9BV9JZSGLvKfw4NWje5eY8m8iMHJL2wOMBgrrnCjS+t
zH9OyLV66Z4dGU6UYY/GrCCYYDSBq+uhqdpYYtUfosMS+sS/nUZ5r9DaY/2xXg8r
yRz15vnPklHlS5V1aC1UoXLzpDJ6E3W4RBQIVFsxOuPm4Te+TmCVf/aAEXL66Ddd
/ys2tMicQ3DwU0P/Mm8KMhWyJfSXtO5RIWvbrKliHAoPrLJryUW/1ha0eXzfwTNf
l4P0wa8XBjHGAyMMkN7er29Pfq7yEiSj/xB9qONFXobKRFk9ydichKC2DOEX8EhB
FWrKQp0Ls0SGB76ZshiVEEAodF1TeUwFFKxBWrcod6xW5/V5PA6NoPOFBGlhaAn5
iyHc7zw95yqr4iM7IFxJTWROFebd3EsnZ8WwEo0AC8bcpicQ60TvhR4Ml11nkPWR
t3gAxwxGRtj4l+S5JDOWHg14xQ9nFKpwrarsupOk0kJvI0jKNrtEt289bE4FFhvA
Ro3oF27BFQB+ETq0T7IX+LrcAbqykPYi0iSeZKDP6Ji5GnMO+FU6E7tUKzJssw98
CusSBrZMrNVA2+ckA2mcNtkqoHI3GG71UDIWHcmMc/a1abV3qgf5yLaNbRoYwZxK
Gz6SHhGCC8w053YLJ1JlJUoUgYjVEpi3nyYddnEGV6c8VRPfaXKU5+R9C2XCuzv4
7XdNiMvvbbDj/W7yNs4jAJJu10p9F7Bb3yRILpnalL7V6BfOdkT1lse7sUMIImrR
gqI84diAOs3Io129PF9IteXipd65cer+6ydPsFnXKJ3pTIwiHxysCVBNI3K5/cIz
9ueWafQmDXoH7vAG1KUN+NWC/2kx7btzVRXKD2BFiDJfW8ewMvveoMIQFIlrZGiZ
eFWmfRQVIQh0Z2YmklbGOVk51WyRbakVcckUn6dzRJN6rCX7wjhrU6+/i2igMwfI
IIrsq24p1LUPV4vi+C0d7H6N6DcJFQ5Ty9kLzy9n6FcK/QsrwA6OwdDXGdZ5EmCY
C4RGTBFVoFHuXjHfJAO+j/4GKjk/Y1ZtYFc8VER3l+7k1LDM7GmleygD/G6KAnJS
0wsLMiy+7MaeucxgTDXkt09KesGx8BMnM20FqBtUrcCNMcNTLz8TM7R0Yqklk+MM
Jh5/wIYZfp4+HJrth+I+YSWKkah+p6VMRdY4+w6fQcfg5K4DdP86haKzH+yR/wbt
1wEggwDM0xEBgIjQdTAAg33JquEv+DrulClt6XRUA1tIUoKPXmPdv8HgGf/ZfmIh
AgmsAL3ubacTy+tkQITp7apzFRxyugTsh778YD8yKY6X/sx/hpmmgTP87jxHVLWS
EwPe+Qwgvx0lC2aUxRxhFn8Zsd3L+5i5KW1O5953bGTYD2yvYD+eQ4G4prAcsNNr
8NXvZ8kocUC9GGZwa1vxjANEh5L/JSHo+qxmX+ijQbr7hU+kM+BlnXiWbG5HHzj2
zeG+uM7RQTRRRCGcU/jMlJDmY/vmTAU1zK8oPMZXbyNEeDRuz1m8z8Tp5MlHPbtY
YHQomQNsovv1nldeXCMpOampOuF1reH0CiOm/SDlTLeB4Q/GEbjYeJ8/3Rs6uWYa
iyOtaP265+KJ2jc2VIGe42CWlndF/WGLZy2M55RT+P+8mAbBcP5xT8nS9DONI8Sg
RtnmNQTfBVgy3jUK8WnpCExY/3oFRi+vDqyE12IC23Gd7NbwmQO6Q9rUrxo9bdb6
yPnm1mYRbdrpvH/FKDVdooKvnY1clM3ztCpTzTOwB6p+KiIkWZDesLDhEyepI5ea
e+ILT55DtYxgSOqcm0HRUGncckatkszSz2gIMA/tJwuTT0geviBO03XrbdM5fznZ
BcQtTurGGttwcgp8MYeI9hh26hUH7o7vPpZdvzafFRGy3o3sW++/8M20U6LuwOCA
q3PbJ/GAhus2VMhW9OjwQ0Ie3TTa2ZdFNaONy28BSQZxIJp22zVEAK/GAq39WOBn
xDPEFk3enNe6ChJBQmtBZX/m+JPra7vQmrJMeOacrU31q9T8Dnk/ByLy6M7w4/2Y
uT7cV4hhIe/YtqFe7GHpe7ShgDRvN6o+bRbzRKcza1UFHMZ7AyI8w7zDIwbqhJK2
l6d8MnZJxL5NolNEDjRmCqs/1WNYRJo4wxMIW6PvlntVdhQj/dJreaimPAUIMGB5
IiGjz4NeDXdgZ3UHwro2NxVbc6m+wYkg91jUjfVChmjLmUVveLkTevThY0kmiMG6
oMcKjG2eINIeAUkzJFTOL8eE7h7Kb6oPiPdKuVRN7i3VLBMjDF6TxC46Ut3taeYt
BPH0HOJhInFDJUFnRUWpJkycWLwey7dVUR0QA0mSISDrfOMSiXr/xYpWpa+UPteC
i4kAFz4eWj3kYWstNTeTNVcS45lpeRbRbjk3YGSfUb648K1vW9MjMbjBtT7caVqf
dt7YtRLsQrHTvyoecG/b63JpdUAj6bsA7OaYvYrzyHIxuCUkJ2ZGG2vt89ecCgj7
3eFR1Uo1JfkXSSEqlvdBEi62DtUqV6cmbDf6KSvbUeK2SGIjL9+g7OH08+tFcq8p
Trbtpj0oO7dEQpjcz1R3UsghCt3UJUKQaJ4oNBny4G7bQiVmJXnVODpIlnyfFGcC
Z5yjftSTg34sgbd+9UUtMdT7t4B83V4iN35R3HtPK7+5nYfcTzo9Y6vYYC6xZSaq
Q0uiZd4Tin3hxjFatBEM2V/wp0UqFBEenmduCk/F9kA5xwQQVVoenWR5tPGJI4Oa
1qjfUsbKGxM7mhEuv8WxgFAgHzPxgyvK+rggt/7GDdSf58md0VT0bBJxW6Y4d58m
pyHH8DA8qsGG90aW9jZrMQHNvRbEQbU5sgQwvGTw3OhrU5GEIoO4VGqn5cM8iWGX
e7oJXnxq1SdverRFxEDvRb7KpYatm3OiiiN2whyw600WFyzjKYjISmPHIOypz+gJ
DB08DXZhKpRqTOrvLuoVE/gy2Z4fnHESzSeuTjM9ORsw29diCkO295DKyAe+565h
suluovr0hqmsrdNEwd5rkfbcsZ7xfIb1pJTUq02x2N4eH7U8JIBxB9THgvwGGWvG
1zlSFXRHi5qvg8jFzzPXF7WN3sE6ErxhuQuVVjumrAW2R5x3yXOEfQy9dtT7LXDZ
KV20nCrwTgCm8N7Ehsc4TKJ5u9ZiwxdQA5KDeD7E8AWDrnq6I6i9iBVIZr+pwFFe
duGBb4mEAWST0FF/cKnESz+Y0TBV7MZeKSpRHSLuuehnvCCt0t0T5BAS9vtDDx/i
sWYliCCG9+m84WKJcWEeov++rtrM2x5hD/S0ft9bH7f/W62sqI2k4+QBgWUyJu+J
t4AIduSkNHZTjei+JSjjuchrMYxKa3O8wg+gMHQlXa5lnibs+iXfplZbkAL41roD
5vmsFUum0LOHlTOqo2DI9YPyP2Y1FTtjZQ+jnJ0ByrVcPj7FkDTizo4wN7NcSmLi
6rS3wsaReqmaM3fGG+Z/30KRF0v4WoO5ZO5yDxJaYRc+5aV1gxLxL618KGIjk2Ze
WH0yneqoeRumuITJohT6FQhAapBVi0F8Kj0G4Lcqhj6ExiBOrsuke4Q6BecnjkxN
CDloF497BFhw0WjOm5GuwbtaVbn7qeJo85HPpTPf5ua1qqN4uAVJKVCb6w+bxbn1
0TXoownkUqTo4uuJ+6p2QrNRx0hga2hnuodDiEluaQWP2fjsxFar16TwGw8N6aiZ
VJP8UF611mjJrCvHdY/8SFBTqmxjphEg090zNLbJXqjJzGwm+FyB/yQF/dmCKUVD
oWDEHOtsxUxEACswGifcg/AIC4ys7XHUWJL1LtPFfFYrYKUYOSozjVlftjQBUVQk
F4VWooh+bgyMXf34A6QEnXlrzRWC3HWdgSV6U7BrgbA7/lZSRU2M6xv3y+FNTVXz
LKc8x688x5fZtvKjPTYSryszPw6/oVJd5Q58c2W/iPKCNgaz4nxRgfbEh1fH7lsk
tSrZ88LGgfx+vSJWfadFlCgunCbr3JvAOVgWJrrxYvvwmFqN4ovCuMg5guLQqVxz
T6uEF7bz0OG1vNmtdRuam5rAtMLk0YnGbbVKGlJBmyZThll/N6BlK20Sn7vWt3mv
DSZxpMqSacSmb4o8nmXZesJMJCqi77ftzegjBVajdta1SeqE95JPzOS0b+aX0P/j
DY2OIerH1kJZZV7ZrsRg4tacH0NjddcT7P8QN9lsHH5UprGj1xih+xypz+HHaOSR
Ndbkp9A6632F8mWMnuWnfaaqoqC6ifTvLRG37C2FYDSpik9aZtDLoUXQ4xdIF7kQ
1SKZxeOiSEzBDqb+tFZVLkEMN69HxGUrzyDfxm1JzSriYluqNN2vK2eiC+vGD0CJ
oAEgJqyi3mzqWTCaJoYSlkUZq/hx1DtFvJSdSY2qxADkOym0Ck2H13H85fKP9Odt
Gn8H9jHNZJ4yHSRZJjKQl3nj1072Cx9yRWcj4vT6FpEhy1j7ZGPgYkCJCdv9+05I
ceeuUGnWWs5okGruSCVrUDZbI39VCUZ0j25Mmo9H24hjOUgSdrhNYFqDITjdXklU
qJsp9JKmS7ZoqIKBlP05h1lhhOPgeLCjxhYSpLmF4GmIDJcvLd+wF1MjXVUWRAby
E38ySeCbTMSIhjxLE/NnDABqzMXqa+hzrtvgbqzLNgKkRmVCbZVFGp68TdfG57w+
oWa/bqv3GV2CRdKkEE/l178tYpaZIehJtFhG4sZt9k5Ovbv1ep7zrYmpCyOn97ye
bUYUzm+YQSjt4lS8uA2nK3Zz+4tW9N1jk0iiMC7R1+MgYqRMCXDBlRcTPE4aztoD
bq8GXRSYUjkxNJJubQ6/9nOBpZx+A0LFfP1d1P22m1SFyfQBRRpW9HKjahijFqQ/
6fFikcdPMPVFftRA+MsYI89NRbg9Y8nyu+IQySpG/kjr1QNszQutpjeV3try0bY8
KE6hmNcDYUTcIp/tXbYuB9GRNXY/AOS/0iy6uv/QisNDHdRSuJB+vn3EZnCtrwsW
xnvcEzb9GOookgcOJlqUl1ymGn6XbQv/smQ1tNE7dCkFYD8taMYiMsTwE9LTJovN
P6Qd3/rbKvIYsqwhB75gjaCGfbNbBpG9+qj97TUHfTtzxKsKkI7buLKXJ+EgA0Ir
g2Lndmyowi+Ikx5mj+BvL+7Oo6r4KQLYpAx3N7uSjEbZGEDpT57IQUoEnqmMR22Y
Zvh7I2zvLqi2ItqjgIAH+eIWxT6Dxp22yYmtSZZic9LSDxuAa7Xab1hhWHBjlhgS
qvDNH8h+Y4M3cxuW/nQx84SYhv41wuWwDtTVOwZyZfN+fvk7r/vACFDR7OP/zvhl
nGySwWha2R/nLvmZWf6BWIwygfSLGmUS8f2WvP8cwHSTM2vBM9iT7s1bgAuWEgYe
mIl5JPEsdG3KLdtvuawnZuW5tNp0HlDVWvWjuAEOb8GF/siU4S3Y50M+EDmZ3XFH
kL+xgj/4vtPPZlyr9SeYXgTWKSEva9MIBC0WrC+UndfabrJ02OtqbiujBjvAhTke
NlfS0k5ENxc3pwaV5b4qgb6WxKHsk06mATmrlyTNZUDPpGb8CicQCtdW74i2U5Jg
KWYMPSG2E/yDf8kGmODVOletSSx6HMdQXySG28mRa9W5S7NxTmBAFkbZzGSl0Q0J
KXO1GoGCDE07pZFTI9jT7RAWfmFT0XjCSDeDCaqUqlfjlMC3P5I9bL/zKG9tQQd5
fop4UG0IfDSwOUTEbEDYEr/NZz2W2wipQStjND/EZ2Io4rVRh33aIPX3fWEZi7N9
kJZQCNhQtwG+3XWCwSJDQ78zf1iZo/S5bfmsFiZEV6RAw2vPQ7+hmFVgq1aoE57j
dHop3wrfMtgLcjQHEl1XUtLpvsF+mvHXuigl4WgKUlg31dwEdLnGakhWpP9pqsWa
CfNsMl1bznEoRZFHDzewLDGZdDhvEhMZf5xz5jgZz5dwuI05fmeWCQy2KuvPgDlV
d93BTmJ5EWVf/XBeYXHh6NVCpEJ198wO2Ym1n3bdY5FOmZQ+M/3/xv3t2Zwjx57Z
gDsbOAOSu8b9fQB3QxydIIgb1jYrFvGRPyHYiGBNNSOCNSI1RVW9qr0Pj91FyjBX
dFwks5ENrIFk5olsEx22XlxX2lLl//MQDA1TrgAHLvuAdlbFCuBzvkeVXt4JoQDj
VWCz+GeT3IPd7iT1FUhjxKCa5iJV75NPEbYu1n9PpmMywu8tZTRQSgWtHURxtNxx
xOUofSJ7Q70K3KwhLlcP0Se1i2ezda19UtDduQytGM08qr6WDH0UZQk73Psy2ISy
kDyj43Itg4sRu3kC3UX7/WikbJol1hRkQPiobt6CeuX2RjV1jtYxHpglMf1lg+P9
XpT/hH622VqcadkhTXXZLflrhFLt4QisSx2pANQXGu4R2fXh5DJXZDtXxpDILCsP
AfrsrIBcgKmYiKdN1Aqqkw/tYI8RU2t5fXpmvK+cW6d+s301Zwew+RFdMC1uReNP
bc5MECaGZ+E2zjAuiNphbEgQDnLBZagc7YrzvR8Bb4+NzdV3ge8k7NnoLJwoPpMq
pVMX1L8yE9pA5XpCgIq7LhjYhgxyvi65tEk+P2S9dtyEgyJPraT1sMi63FTfDz7F
n/HDeAfzRYah6KINnYWXiJlbPzjpj+3yRaUcFu8HRc1g9RXe15SMKoh+rLBFKgM9
mrwM9scYYqecgPj1E8NNjmizncc9eWxKhAcid7eun84SVpNBC5BGwz20m11Q7wvM
JnGr/An8ZL0dFF+kHPRdwY9q9PBUTqOpfqbb0TYaxLEvaUAxPuOr4xRzFyJ27k0w
oEkYZA9b29bJbp6Hx043LzqhD5f4LcPpSn8d+92+IuZSQGOIUXflQpQiQc8hkGS5
QuEbWodlJEd5a6DlDEaWB73eeVJCtSlISqg0UDN4rq16ICTU20cZx6AzOdxb4LH9
SfAUwyrbITCx5SA0O7OzC3hYzATVF3V1lTBI4WU0vIo7OHk5bCqzYgjVdzqRoo/G
avDtG92iUIIms4u9fLRP2IN2ejNDyZAZEUcx5xvl869TlbtyuiA61FPi2rywfse0
2aI8se7MAjbzoQ+aSe1LYfbp8qHvv88nafQAV1ij9M5mR5RzdUXs0wYd08hmzeDV
5ohxqBnvh9Y/ggwJW352S/QDmTSDThyK5Y79F2v/qm54Tj/CYgBNPFAyliSpsJVd
00vWyqo0rtV88/jEA2NJwr4V8wgh8kDoJvXF9ZJXQSwFpvwn3qKlfZn+/8oiateM
iC2oi0BvNCwQMRKx/1RfM/Ev3MSo/6LR0/Hc7KgySCTMRGtDZEQyz5OthPOK98h2
aF91NBaTmVpvy+glKcQKC+fsbvGZIXyiH2DVaLpG3KwDHg2YcFTNM1RfNxIhjiTF
ibJIBttcVXPEj/Eve7agI/xvWv1ocO7fBXG3M4GpOtak9mnLNXWmUWMTcfOSKYPa
keWf/gKlZBvxqXwnF1Pwy24pMmkqvFEJFqUC8xXotKcsXBHYDFnnURk/smim+7Jq
f+22J0C8NyJflUbh7zvFyfyCm+BGPogmqrRyeWPOkSLFjR4d7GE0K3QC9z6gBOQj
RhD71TuLlSQVVoa3fww9XSho20wgste5CsxvwTZ6Unw+dDZsCYVQ+BbaOxwZwpoJ
n5MRL3RzJM4W/LN3mqAVkZReis+OgxMAdIVqup4JhXl292iKcpvJTtkb/FV5WbbE
0M6erO6lHvXqzY+4WiI8e8SbHAeS0xtJWkW3hzXh8mTVQ0t6Pt7L7o2EVV0xfVPB
3l+iCQvzycZtCnFRwo67jSLagS1ON6oFC7EJvBv16/1QYvUA7N1dvViboJHo0V+v
Voyp6Zk3pVlvfn5lG7gnxxfcoC3J8bGb02+nG2vJ3DKHUyGt4U5l9LNVf4pBhroC
b4sgjXJwJPKT/nw2a4vMBm0Gaa0X7Q52swHx/3WVYi35xCbemfAQ5h1ER+QSRk59
ZGh0R+VTOQoPRCqSDqVz9LQebgK1AWmjnzDvE90AZ72UQv7J1UJczeG4RXl6Vkin
EjfXg14b1tw+PB/UWpfngt/65TimOde/gbm7fIopL8iRb1QQve8ghmY2X2xjhMFE
InXIDYMDZ/LWCD7txEJhMPLZ2U2Dko3YvZIsle6jLpym7eS/O1Oki+4re+uX+q17
Lcz1tfoiw6CIDdOgpq1stZc0weXJCGaAR+6xZywOMIja0Oa/YNGQoAg/GFrrrfXP
zIyyWfyMHSwbKaMT4HmGBLVSlDWmljGRWW6b1LCR6UED/zeoPm89XL3FEYi6lf+f
mnde0ptDLObEyBNu5pMbyEUq4ons0ndU2sJHgtursvLOhAYdOxWn9CB5UAjgJnsK
VIGr7GhShHzvzcZrSu00nGPYz4QSHbwpOp0QSzfS81dw6Iv3kp+iYloP0NeL0BYq
ueQ2zeKUQqJp5GxU7ZYeHxLVYnmwpAT7GV2l6tw6lgVV61Iw+gMHKOJbe2w0qngr
m6zI6EjgQXxBKdcn4QkJtF6x1Pe3ReNnJbM388pUFaPLmYMCUGBmA7Ax6vi+n4EV
y/4/ak5EmtfVY6UEYK2bqu5gZ90q6uWLbDNMAW/VQSyII0kcJ1sqcFTxVnY5aKwT
IWZiyJg1jB3/A6j4iH8kd/TVWN18tdHqrxRkHJFhwBQrWOnPvQ+XPEc18Ps2Oeki
uCgzQiVz2Xp6iRqqR01M3B5mmFurrUBNQ2+zjGWV6WdNnJADiOGSdfxK4MwZvtpL
pZ/ZB62JlGEZH3wGSlINK/DBzRsm/hIgyoaMwyVPlhBZC8r/HiRd7r8X5QjXjjEh
6Ol7NRIvNbHqFOFNrKTQ/5duA4z0d5UlCw6mSQdcbBrpdODoO4p/zyEobr05Orgo
y6GzxqW4sfp3t/m5zg02rBuDTmXkSmTEUp4IF91g6V2GnrR3wCrixziYKssB5Fbx
NE1/lz4OxJH/9M8Oofd2tT8ZrCiuxCr4o9w1VPc1+je3U5k6+cAsLT8YsNQ0OSVF
E33FnCD5Z5c+EI67x4OcRMoGeQFeV6B+im7virycJghNCzMD4fAtif3k1hhUmBB6
LiFtSaLVz8t/m1GCDQkhlnKJ8xjJXqhf0qDorY5DPg8Tx4UHEWWMj5DRjVOXwc5P
oKhjgyqxrO00sfOYDexsJSt0DJtu4RxJe1EGQC4UY5TelJe0FfFLR8eAYIFMkBs8
obnPmAYd3FcONRZ8o/OwgMMaQNin4gj5VNQqWObNLEA2CpP7s1Bw0kUp7NHt9RKs
9G0AQaOAZp1+O6VfodXDHaom8FPlIzQTcYtrrirv/57K6vvofyj5YA5RxZ8MB6nh
FpnXhRqjrpqVfRD4fXrhXoPfeAzhwncZSY165z34KOT9DVoFFPwRxWMHr5Q227SH
/Z7zdivO0Lb7okSXLNxtPMlTGg2p4ZIz2HygWpxg913GR3wr6DddbCcAbZPkTw0c
nLsmGsJDtzn6ELpN6DC396dE48b1Wy8LnIZkzVyMbXaz8NQT3PqVZItY8X2cGLbb
M1KYM6YndLzXbUOdCKZ5Lh5+UkKwh07ZDMtZL7XV4X+WvhuScUHEyhXwvsyYmwGH
WSSo27DQWff2EdjTmNAhRe1uIEwbd62maIMlxatEzq+fBjyD0OlNfjZo1zDbrNcg
S97pZMrTo2N6TuwHuTdlFq9+ViT/+bFYXDAWnpdMzqyiMPcGVrxCdUQGF88ypyxt
vgUVzDfrJnOSAxAqmV7xnaf637ao+iF/XS9jrJkljyRF3YZl7qjUEz9wEAnD5KP3
DYnxwfrJkQFc9RLxBRRif13pT0Wsa5n75YUsC8krTpypVCpynYcorzQtjJVvzN7K
kIOgMacUL0Cvqm6lklEDWN7KYC0zF1IxhPLBxlCC0UI+JezSVN2hYlO7KCHgETmh
GMm5zJ/VT1Bg+qu1Fxjwyphq6I+XuRs+96HCVtkXwVMoXh8J/Rz7YIUVh3zSjYrx
91sFiGnWl7Eaqkt7walePWaykDyel/vlneIVWDQMrvBnbdbhOHXUyZUKFWW1tjRI
ru45GDKgtCAOs9SmNx5cVuW+ss5Uudf5KDsN+4uem3OqNBTPMniw2r5N0FGK5uqn
B5X/G/U1FhXVTaiC0Gm0tS2H2Hmn44MFr4VNPjS5tJPagwL7ZSYvrbz4d6N4qJwG
ZGLUb+sUUR4KDOC041WOuac8l9/KVoaM7B3zn+X7xkkH6UDHIISO4oFEWskl1joH
lUwyFECjlSUPGQ5lGRId27YJL62r0egZa66eywRER8uDzZh5UslSEQ5W5GFDFbE4
tvIcnTDRR2jxroN9NcO0HlgKtg78Oxdl/dcuauKB9SsNgRwgdcA0m0+6cUDN/Phr
QPE00KisE6Jqr7AKD27vExnG0d+l4hnUmmG4TfgOeKmfmvHqbLluR7YwnUsEWgFe
6q8NyBz0yRAQZlHGyMmxKQj2lTzUYlelBpYI3VvIzt0aauNslV7g3GZqhKwnt1PP
NWEzDwye2FYslxsJyxtSjaNRwNUqq5qrxMaVnsi0Szi0o9SFWWDl4Z2EHotnDP20
5EmYm9P1E/Wg8jmBnKFovo3QFkEetAMmasxZabi9z7TKtEltv+uEGi5aLqoYp51g
N9O+YkCYAETYj6gZFGo/D8YnGkyFz1y+VCq9E+2ZXtwwoENhGukcAtPsJSykI6bw
L8vTkpXOcPdRAxq0Kt8HlD7UX4sbrOmNZuUGqnLyOfYMZFmXRucGd+w3STk8bnV1
TEWsh64NnlFzkItzOQ+NCUzkGZ7ZZVPThn8jWkBEkYAvEnhoC/jj86XNJmj/Q50G
y9WGlYvSH7IwkvqcDes2G1AYQ+ac1YGGCB+vY8sNKhm2ESI+WGXH1zVm4jIFQYTX
NemTMlyixWNb4Kqu97AfK5IWO/U6Vn9VbwcuBILIyF6Fa1cOAetnFjO0bi95BDin
MnodggBGvr/i2tRTIYD9b7WlVC60eMX92IJsRb9YNEdlFfjxtix8JLrzqzoJC0xk
CZmTJcvZ9kc9HzgW5hApy+7S69ge8vhnGqgjesyvY04Nki1KPr1veX63TCI3IpyN
6G0s99ZM9lsZqss2CQ56DeQSx7IoROb9rYqoatokp3mJrYp+M7707zXsbaW7d4DM
oUdSXWfOe4KiO1AuG+uu+0FcDm6axOc8EFPwmnKaJc2Sg6MZf9Pzrc6yOWw1ieNO
qBipPfBCpwPcMjnpJJAfxo3qvSo08wG+VY6u41lUuXxps04KBIwLiRqS6MzI0Vji
HHJ/ctiafGldk1on8Zd9vXZEsS1O9ltQV9IAU8XD5fnSqCbM+gW7pxKO77jYAaPE
dn61/DC0BLyms9wRsi7Vl+zarwpxYYadJMW7df3+WtGvWUn7+xAwfu97HSVFmcYA
BVW8zxABrO99IoQ8Blm9/KcDCqG7oELBoKpTp4Beumfs6ObqA5AjQtfrMebdYW74
JYkdOuxbnDaXRjn1t7P+9GDEQ40XfXqZra6muSh3VwfEuSNnbiTQu6gyjdd+W9xo
skPkTjwvSwtMOzzoaasrqqczBOmxzISLY0rDPRZWGObO0OerfPJ6NbwVd86NUxtb
cbB/ZitLPHaXIVxMrAfMo0ZS0EinsyKNsFRXdZk7PiIesCRJyYBftD4kI9wEd0Zw
2yR0ElbkQpVauQbu8mM7iNpoOJ/mTJPwcQQV3wH1et0XOWni64k858NoDi/Z+F25
USk84Dk59E1We4F1GZfT3nhRxz4zBbQluv5TXCLWk/O4ze37tZuqz4yBf1h8IiXI
61yl4/3g8fNoor/j/ijRD+oUaIt4YGHM+x1cbFOqD3GlAVQeQHKyCbzKs0w3VlzG
5HZ4Mgk66Iyzn9mef3q16BRVkkC61F1JOrhc9/FcO2QYts/8EbIMF/mYJFctgFbE
buRbK5fQJ81TW3e6k7tKa+6rgsG32CNyNlBawqe2ImfwLmNVxl2S2DNzSRyHfO0o
eCPyGSOo9sSV8am7iW/yo832ZKHq2/nEG54oyZRWty9vl6fOQcpHLEk2YGkhvMZc
dgLniu7Olxv46dWxuAcorTcZ4d6tBSx+ehgGfZmS+scwCB8emdPbATJMLppDAaXP
uXaXXs+Fy9CWi+aqPaY0PE86SRBFWCGKrLfU44Tz1wBg1YAGA3B6qWBSzTv9U6vG
YXe+qTTrjhd3g8OyfxAmxex8p/ogBL+bnJQLebz816lkSXp9Bx2/OGcsKBpZvNFP
U4wCNPGkS/7gq/KS+3Mz9lmiavk9Bc/+1fXl8Wdidjz1T9iIem0k0s1YGvjf/KmQ
FxBuaKfAl1UHqBuxL39y7BZ1maDMAs0QtR4rjvDIcqBNwxsp6HWSAs1jNoRtEicN
EQyHPA1ebqqorGT2PnAuZHb0gSOMt4gOMlbntk+aXjC9VArR5soWp6BEuo4KyjA0
tgPKwWjBSVGTAlUpl+uIFsixCtWXF567GxmyEN6oqE7jRBKBEF+jaIv6idJmPaaf
cp5zOC6DauQdSklyk+CumyviD92EpUVMovN7Gz/K0Lldp5arlDyAkQrMl5O2RBX5
PxBlEwQz2pRxrZlpVo2a76RArEsVfCga3qtRr+54wTEJvamiuunRUHGi4zUET/6N
tW3WXb935bykWtXdqfNH6zc6I0ZDxBEI3vOqUfq2Mha0n+Svv59Bz6i2QYEPvITP
E9H7ezUfXd3HYyQf3t2/Qid7yFom//yti3jOMRGGZ2DSNitukZb5uWaLkPU0k8U3
mqb3qWZWeKnErD5S4Dua5L029WBdC71p6sSZcyPnGGCH2EugnYqetS2poiF+q2aI
hJut9xuaSCauJCQvNVWSkCVZqexVmDoAIhLJVZAdpcjnMmD791vHsmb5uxOjHHhZ
IznkoYZnHDqEhMNu/TJH9ERMqbEGwK5SqU6OCnSvh2Bdm/WTlhDyFdnGwHv0yuEv
CTOvwF7wcGr/v0evTpPyUKK19QkxNiqMgNuIezdqYFK/RwAuNGU+LuxDSD6Io4cE
gZt383uUeeLz2hgnb4Cdf56Ph8J7s6bkqJsTWnTShCHwNoKL6T5/QKwrVuGjUOsj
fQpfxrMNH55d8Y82KTGemBs6C/3h1Arv3QcLaCiI6q4WfmCvDTTy78Hkghr0hLKE
xck01xlcUVB6ZgHXoyXgpsP5UWO0N7bnofIo2YLzYFR4+xnKZom846IhTJnFNX86
+AruYgMnLzpCWtNZqf1Q3DXbUyMXWrbncejNwYVUkbhtfQbVWdod9hDUU8EAN6d0
U8mulTFQQDJRMpwXC1ROKjNzo++yC7bD9UqVFZSU67lx48E7oPbGU3lKWIW1xS7i
14L2pWHalDF2s6sCg3QSLfEceY7Ri2+VyQ0Dvlygz2s+XRiXUnWLXQa+oNxu9Pyw
8WCiqZ7MCrLYb/a8ZR04d+AZhXds8mZ00rSi60fO2RhsjGZX/fezfInNFlNn/qrZ
kKNvSqjTju6kDtP14cVellz1Hnk5ivvWCrCb0xWN0FkjBqmYB+KLRstnR5s7/EvC
Sh+BDoL96T0pIJfUfiECyCZIWE1Q4yMvYw4lzhximyYPmeFWXXNWkVyJgyxtVyat
EHY75HN9oCo+83VIYiUtdlthMfhI2iR+4F+j+6j2hMKGmCbpDESDBnUewXQgjKMz
Bjr483B1uvl0bAbE35mTt9BMCV07RVDsDldV6D9GurD9kryKGOJrZmcAOPuWLPOk
XelmzIdx42Xp8UP0d+N7RbIN/UpPz86tl0S9Hc/m3jymBd8i0eN/b58HqJU5MFnS
ERfp9YycLnyAlduK3jKbBC5/2JkAtrBT0uiJBVR3nZD5sctlombF3ifp4W7EdCJq
6Uxg+huWKayBgWx4Q84t21D6qyu39Bjs0FjS4MrQj8BM9Z4yIbNeW5vJP4JJQz2E
Te+czVgy8WNTsKpT4jGrrGYM+0Y2PCn9PgoaAmknSfazaPQwvA86zDm2v0fjLvXb
0A27Zdb7xp33zx5YFSwixxRMjCwMiBZ/C/AAIS270T9OBYpzhOaOFw+ptgavu/NV
/j/2G8cIYxhqSiPB3vUPzMFhhWKC8+IGc8FQGc8Q+Upxf0Gkx103P5NV8Bxlbxmz
PEK05fJXjXcnK9Fyf2p/3LQezNvNYRaWgJGEFB45ndMKow5kvYAZIMDUSEEqXUFf
tFsFkdSiZm0+k4QtviGwaxPOKG8+9Yw0UNJm477t3ud+5CFWeD/iiX9nSIULNZ6r
km1+tWBiVPjxEtwrGNEmi0O+6durciCf1wv1quapkXHWTZf28YyEfS/X9tMqTASS
AEP/D9Z8Xss3Rj+XpWviwm5dyQlkb8HG7+4g7hu/xs6cCW1CvkD3jqIE7mgga0lw
Wr5U55z1NvtLDbZ7d290bmWAOn2gLb1iriLD8aPHnQUtCVHR9mQdMNI3VLv8nd5O
IGwkrHi5uvqsAKeSqYnnq+9zd+UVby5uip6SKYFo2+Fdry7YVsof382Ox+Kq0lNa
TAareQMqEPZjAyNkTPWzkQ292aamH3unqfluX8P6cnsXFl63l43DojRLcBxuNLFH
Qe70PZrMJDW9NUOLSNWl8aqguREXPSQlegWbdLLT+rJjq9RVMqlr8uCHk4rxNC02
D6ZzDm+YgPAROvlMvJnR1RKqnHOR84DinlhdY9moE+d8EwPCVSpgDgqyKPTj72hq
6C6fdvQjLX1+ExS9HQcSPmuKc2YPOooK5RrfjPLNCmPbqxB2yxYa2ira/YVc666T
OBIzRD+6AeXaa34CxGryAVyYXBCWk/DxOCgzsU9WfGeJVie/UPRGk7vwJlftmQpb
rPU3hGj063W3pqg0Ux/cDcHZ4gN1g34C3gSm1/aOpCfRjZuVhWUpUTKA8AZYsaWU
Waq7kooAjFVoaXgKJV1iWjqDe9oNlmzpksxIIu4i18lm4NoJAVveTJjvDkmvd4rX
Ue0k7OwFKKNLeSe9jEEGxt7Kp0x5Oj93bdjnxLbAj1PEtWp+WSugTLXbMgZCJHvW
4uW2WNJRsQAEZPJ2qq7vDYueW2oo+ICof4L9xwZduN4fkvDtmbK04MdpOXI567kG
jRLy7HPr3HRKcPMjmgNPumGT5vYke0gPhiyA9n7pwJUiw+AmKdMEA9onquxjdcQB
KvnRFcwsSyQnGGrA7pa3Dw2f/G+C0AhICTyjESqMMJ6ohiYyk9IGoU0GmpwjZMZO
mbV7jP7GnRRh/088dMt1uWSxLRkPDGCYzqDmm9RaI8KGeLSN3xmSiJ1YJUAAqQ31
fXIsnwLxcN4wuwtqshOoT5MMAcIePpqhOgiGn695BQtmWC9ZpOTq/d1QNxq0NYkn
UzCKdXt8czzGxdsxfbKwRjMusnON0dvQMcbRJCI+J+STIOPX2iOJ/X8+QAbK+lQ9
KZuBibLlJKE+Y46hSKTM7rFO1PRifQv2unLeBvmT5n9NibHrucWRmk0xxwHwcB11
4TFWYQNNBo4YULEX1nKmwqAVYBFHckqtHiEKrApP9qYGudcVz7J5SOgmchre6h2A
GKej5LmSlyZ8bSPO2OT6Bb+UAk4DD3rdk0OvCkPztqgGl9aoS5+/hlL6p2qU/9f9
I477TMc6AknjoANbcVxezRaGGOL0c/shxGgKvlhSJSGn4ZCdcCvY0MgN8BZ4akhR
Yhf6oh8Y/sU8wYrSWcaun80b/hIUUwW0kD0nwLsWgeTga3RN+LCzJ5aBOFqvzyK1
UEoPwpYdeVkxmn02+n8bK70l/yr8FTsJywdqzuP6hG67Yv/GafYP4xUPhoScngrd
Kd5eJ8Xbzq9YWKnv20/8HGCzxo/oIFbdtFYRgwRrmhymhAOy3C0S3VrMtn8cPOtE
xaZ0Nd3xiKrk0+QnagrNhfA8UyLKVFgqbjmzub1w0mvvWYc8Py2A+6LS28oTggM+
rXvQ+oN0/5W8ABiuLQTkJxcwW4O9TzjRM9uXH5hv7j6XgqaAQoH/I9fJxJLZX1Rs
PZMcHKnYFdD8OXpeHkWGJqBvYuJMZPWjvWfhdTWRBFZxbn0VWpF27JZ07VkheTUx
hmaWTMi3iUufKoeI3wuwOTENMU5QxUH20jBYlQYARqETzBfBz9V6vFQCtpF2hQ15
/+AiS75RXCeNXtupApYsN1uB0j9skaJaQRMUYvpUEHVvNZcMxr1SLfeEWfOmslkQ
QG+AuT/RYo6hacTsHK4jD9EHc4dCkuvUYbx9/LmgEtdTmIFNVWWIEs9eaxK8XiCB
sN+2ZvGVTU9NmfIjTq9RQy4yFvJDHaQOxD4eCeadfFGdRmDpTigbnWetL6VTV9zV
whPovW8SsJFHnxGlrOgDzaudWU1wUT9grqLf7+X7pk2Y+IbUdsbmHMfhGrM62uO7
I9EhengURkH+9jI1yshh216VNJK44loAaeIBSDC74XjN6X1n4qkZ8pgCySuSHVKD
8vuk1UbMkIqElrW5k1lSyY2nEJlqhV1yZEh71XIpHf2hxSk0Sawaj9taQFTDp+YI
UV7GeP9BIfwOFOEEjyI3vN1raxLbYeUX8SeBsKbaZIEDr+/C0WJzWheIiR6qGL5P
b7TFpPGdlkDhUCXfAbEiHHihI5Q0KWsSRrf1FYgesOj1kBlQMtz7kISlmfpemU9Y
NauWqys43mQYkLj63vGWbqszc7WMD9C+TaVllQ0RSQNvAF8g8tOf3yIdJRTZS+xg
6vtPxrB3BeBBu3vKnlqSuyJ93g+ASrIprnXJqKLG0OGMlIl/3LkhdxYaP1dYh4AF
SNJ7loAu+/J8cZlaOq817fmt88qSzmUGJy15qBYrucl/YOctkyrry4M9ZzNOFQk2
XVV7ks2ceEtI52YqaCkwFQ9RMgsGZ67yq6H01J/FS/KPcPi38MhEblQSTTon+KxS
w3DGcuIDduxRTmKV6Cemt48IpB2RxxyRT4KFjcmqMifiXQ+A0oWqOVPBQ0glBwCh
DHJZ6ZUPgbPj0uqcRTURXk+ZsGT7N6XfrjDDtL/mFx41UdoK1p0LMMiFBxkpjgtG
8Epn+SRUNxry67lW2lC5IPteaIuj31XP2yrICSMWxm4ptotG1XfJ33GSqtBkRGY+
iat8sMzIiL45Y7UImjXIPt7QWeabsddcguEDcxO5J1OdMB1DSdwKGeDhNK1NDU6I
B0iaAPFmt1kDle0WCTgKYGUWC5lUCam/zWILKXL/qyAHV4LzBylomrfRB6GWgRQg
+ndSu1MVYTkicG4MvXlmHPcv/lgWh//HKQBSvcNKyhgZ7RNupxldgODFUBoxiuOA
knBN/R+sir8FFJNMlhBt1gNJq8N0t5Uy5Kufp1kxvFl7jI3ujJxGbCIG4Drc4vz8
A+Uqusz+CZ7McXTOqM6BDmY94Rw9rNzOcyQmCsrHeWQazlI0BHcE74w8vznUjnBN
WOkFAXY6VowonHMNxYQ7aH2zFZcHFjCGmwY0bAjbKW0AaXpircORPqTbD0kYgq0S
77/u0qWL61h5Cul4Re8T20YjqIRWRvWXxHHfQ+dyuSerGrFgX5B8WcT6qqfMmJq1
/tRPGZfmDYk5TVpi6VNRQFTBnz4rKHT8qDACpG+fnONN9XZ9n/w/uYYX0aWZ9StN
2AlAVDePgjy9JAK7k7I4JRQCfhkYyUE3AyvgR1oL38XPJJB8MQi3tV2CJ8pf9cTO
bxCxPQu5RCsFT8ZG6HBNnknJloeYUPln9Hmw25Tpv/2YBbxb6aCBQmxBwP6jGB+b
9ckxWB+DBa0q7crUjgkr2NUb2OsicsBRVGjRaIVUvb6MqFoNdaR47IvWy/VfRb+h
JbPiuXqzTBR/I/bJuv7CjH0DzWBAcTXXVAmCftkDjj19gqZ0j1fgMO/MJW/9TIYn
zsJDiz7XtLM/2UKu5tQY9eSanPlfc4yQniY9XM3rJveAdCgSi+6Pqg77u1vqSl77
E8HySGx8uyQX0CoEYo5ftKgCVmw3MwpSVqv9CevJ9JKZVPaOMkaybBehErJm2YoQ
Dy+wJbqHRI1KN/VNrsa1MsIuI5Y/Ia8ZmRgRb0wXowKq/XQyT+DHl8f2T7swJRmt
mZMcKwH93vbJyEJJmu9xV5jpRuX3ymwlniCDsiQ/iv11471xIKSaoPuKzp2ZQ13H
bXSfm4gjJ/OACNkLDr9O/0sPkD+wolvdM0QdI7peKDwTP1r/04jx+uW0REZv3ehn
QQ9KIxyuzDiHvtAru+VyccFu5OJUupu28z2DdcVy3yUwDmv1EBIKvs6BG9iD0/b8
DHCclj/x/F39GvAs/ip4AGj8ZIbxYbgggCPJ4XIhnGxZ8rRFX3/gBFia1fzeFngq
k8C5ZnGe5WQyhpwWTgpIMzgcqJD+8lFUILnQwbWKpjnXX6hOsHdjDG7FrNFL3VJS
4raJszPnCx3mcWjEAut0LV8h2sC5N7xA7YrMWMEZr4qAEZGMTe2oFfkxnHFbGCxc
43xbwYpqOk8du8oJWVDY+tSEoMBnrOfBptCfHrEb/liKxl2HJdanoLritt3ey6w0
CBgEsCDbKO6jkRIA5glXBh3wycDZhJD2xgz9wzH/SeuwZrjEUGmbxhdqCbHZik+m
oXa1+jXygvSCIb8BjY6VXxuaN7sbSdyLIuYksNsOjOz7Rp3MECcjiOseckf+RjtW
UPkA9uPufAC3ta/GRz/UrCa19bA2at7/I/5krAIipggk25C+rgTRXdVqiTBPHeOo
htryemt2WWbqdu18o/tEY6ley3pXCFv0lltaLAHM0DZNAwegBrNCYC3PqkLkB4U0
+YqRMeKL05EbXSR+/+bKHe7qPSgmQ1xV2G0913eQNVOgxKlzBn/IO4JyrQIMMpZr
M1OCbN6FnKbVoWNJ9KOk9iO+s62RCr/VAo3MMyJgQvYKDDi7nWBqMplvmgEXum8K
U86wokLlAUCDtOpe+oL4RjZx8qp0SaHBxBZxP6jBKRc0jEhm8+m1ffwlyxzUGqt9
7c7uiXXUT1gt55UU2ZQL45aTOxx+dpxqslglnUZlNJmP3yNJ9IhRbw3ZHqUkcSX3
ZBl/rheScBZRRaiglBXHsev3HcKQ6GctQDUovfJYtDyXOyLc9C8ct/dRsLZazuqQ
nY8fjcSE/lLAC47DgSsFNbeXX8xH3u1F5U3T60046ChKDemN/g2fFqA7UeLPgehl
dLAWLMxneC7I5m1P1kLplz/TWE0k5xDVI9NgsdzPBqGuMqIF9E9gCmM/HLR36bb4
o40ZwWwIyZGtSVnHhF3rx88RfgMynSNsA+3ubuF1ptq9LFdGhzLmjBiYs+gWQDqb
jXgaxafL+EgyrGPWU6BcVKljZ75C72rPhQEWWY9Ih+JK6YfvsDUfrxArMG3bJyyA
nuuWKV4Z3XaJ3s4/uv65VgEEAwMkogZ7Jbjt0MtfeXchKlXBIRNFtM92UnLu6XXe
ecms2M+b6iCM8lj2hl8CtkwdyWzbYk2NkmDMg2yTgvkmbqqormNRkQ+TgKgKoeON
yB18YRozqum7kIAB5i5E7WwxGNB0AnWa4tOQeETfK8Ty0F5JAUlngKcEZQf68v8j
7KYdfqLMnkayIdtDKevk8gfI2XtG/qIwSmWKFsJf8zwiH38dOWUPN+W5pnqhabKG
/fnjKTsol5x3lhGPu4QvUWFAXZX89+t1drudtkOZ59ZbXBPmXbxTt9zBGpjreS1+
6VtcFRelmY+bm4svgGBpigxtbyKHTC7q2l8/YM6Uj2mSGd006PBAgd6BTol6wUAK
H0XE/YlJrFYPckg6Vo5mrxTrQVivUzFw/cQ4c4789vCoJKSTUqwD85OGiHQ1Drh2
7byk2lnB7tVIYAvH1EqympFQ+dvXCcF+g4qDKbw43HRReMqKKNI6+oDAIhxAgjgj
L288RMFBsag9nJXldTBKSUfOgJdMKGtRyVnhFsUupSXa0QkxMEXPOB5q7oBz/px2
EiqGep/slFMuUORHiEhHQ+YdYUcrbryHSDrwLrh5c4E7TwpQJIf6kZQ3rOBbuHGJ
MvANQHmeoD0S1/TmhdF4CSiF47rrrgQhmoFF9M0CK9/0DwahYZgs+VmJa0//jX8M
x65Q/iwnKyJFyEfouI3KaDwj10wlR7xEdimxDz+QJ0EvyYDsM2AzSOIgerFYay2F
3NncMWKOK+rMm7yWVVIAAEOKT399bG3xZSCcPY+8GiHB5PCvAKFE7iv0x6SRTJf5
IMTKINsr3JJMGdJFQKs0HIrskyAHlcdYu2GgC0QicbBi9583/vpiq4hf+OrLb+h+
I8MbcnEJPe8y4PG6Oy/q6l2qqF9MSxM7IVJHE6hrnUr6o/8OueF/Gryy7TU3DY6x
viYqGa+tTFCitbp3LOAoubQSaGYKdGxLlSyBpDSJziJptuxD49+DDIdCWT97DiHE
ZATkD2N7VXhBupNjOMBD+A9qfHOiiFqbQS38Bjq5yJIrI9oLORn82aVw5vnQKuYw
eLgI5z+JXGRx+pFsnDfIuV3oaST5197inDJdVrmeUdLiXIcasj61uL1u9c5HMBAD
C1Wm1HNQzwcd0AWGjSABkyeHhEamDESD+KXznIC35JLnO1E9JwF0IS5Uf9LlB9cr
YO3O6QBHePdWbTGq4kGpKaxK/Ysanf7GO2i0azxKWtKNigRbkR+SWaPz19l7reQM
lDso/wzsEKoq3H/b8RYwj69zOcD3EJ5pJVnxwmx9GC/QJZa5zdlPKN+TZShPsjV9
n+8wV6dyw0Squ6ahGuDHgGbw9tTQZwJN6w3cnXpK/9cDL8ZkpK/vTigYkjw3selL
0TbE96T2uOpKRXWzLp7n+jOUUVM7y0N6yF0TiNFkcEmirHfknpiXNPfEsLHBLQLO
eEFMizgxrbPym3sVta9KrteN0f1vjet877YrXHbE8Tj/EmAqKqGdYI5j+mECx/5n
qbMC+XV6LVKk+G9AOmeTNQAyLUoFxvfwCH9dwFlCHMY24+sXToDrx/E58Uc/Ga2p
7Kg3XxSsbl5F5+T8a93coUyNJsRmu9oZgPOnBW1AczhBfLXyQhX6hr89ym0Jx1aY
03NYw2mB6Xguqg8QlNmoFIWHmWRJy0Xi47f3teTg4d03zQBQ5LjRXR789P+E12n2
nd86VyO4vNk3OX06BIke4j+zVNtK64DtB3zc4217UOMnDDlnZGCvs8FMccR8hXCO
vYmZkgK4LJo7DJg+jS+jbgCKFO8CxLtcey4aaUpH2lcDeHZ2PScYt0hqhHh6tjI4
AXNePUdgnOqql8mID28l9gSaeyFwCZc1CH4UcmLZzCCqXDWHZpANYwgJ5DI2XtV6
c40c0l9O1Bv49wjTvK5i8nLEAraV+x5iBtxZZfYUDc38EYGZgS7wBzrGEX1gECu9
ipxJEG0U8j+tBtbhC07ceORBrTGWOaQUXoog49/E3lk/MmcmKlXzlsiL/7PrfXXo
poa+BALNZfPahRgqfqxADX74Z01OVcVm7PApsuYwSqorNUesbICzPXaQQXoVxlQU
zejiI5w8ZTB0Z4GByV+lRUc5S+hLCN48U1Yo5sEy0RWogwTSOZiulZBJlW2teh8h
z4KGWFk1kk+5q5fEWwQZ4uSVZMzJ3SkuARmy9hJyqqvNLrKcz0Ssf7ZszFtJC2gx
7ufn3MAOaG+KwtFh0WRGBJIm/aYPOwzAu9iSyLYeON/qCL2LbL4HYX+QwPvrt6Vx
SwuHToi+oosvsqOGk09UWXpwIrZxr3MIiy5O3HfGMpyMvLg9s6rTM1XUftj6gmod
t9Bu1q+0lxJ/vjrF8LlC2Tj++X0WMzdHVcNVBl1X4MsL+uOf+c2SzIkI9xrF0qRP
aqDiKwQCN04tX0v8+mpEivKx1/De150eWIWBOJHy0DC3z5ENU/z2dOnk9ot3sUY2
SQkHtiozr0VTfgmvh7kWTeXlcfudC08j+d4qCAbtTHEMS+yY2NhGi8IZKq1KG+UJ
cW7xzXwIKUSxWVky2fwAz2Aw3c0CnM7RklEN5O39PjKh9LOCNdwBdLRsmKB8vo20
HoJlZPSPohVm29XUtWq+6iPeE3s5dqDgKqllPowNMP7wzsSsQj8YEFj0WMi028IW
2EuASwfTJGFUDQCFOSHRc6x9a04H3bEPCcwMEYnIQxdDf8fSDa/vYrEMM9zwEWlH
ckfJIGGrD6GgqybmUw7GfdareMCJpg9YXHoA1aKa7TRxVdjwFC8CRTFkvS0LC727
7UZGrZnFk04PsXujc0geZQzfj/xMpkNVGOy3YlDOu30ZEK19Dqu7kMkyUhh5Z8Ba
ynJdqdwMAA0wj/b/WT5g3p3cmyL2j/CVLbhsAFb7VNjvgKCM9s/7AcFjlJwHFao1
9ibDG6//a3U5t1UmV3yoXxf1OI2P5sX2OW2Lb8eNEUguHPw7pz33pqoOIeDXDPwn
QcjuV0WK0fdKn/IJrbhMxQ+112Vf6XVq+wbleq61s5lRw2cErtnYP2RkGzJ3duEt
VFFWBAUF4PFCeUy38qMOA0kAMfcPhQyggK8ilQkWS45BFUidLlgR/B4+72ZRQyJn
shr5D5ss+zTkDWG6NhvL/vfq756IreR57CY3jragrP8cj4ntw71KMsQ5L2qPA302
78v5bImLYMqmcbvAuojG2UHryk5dv2i5NpRS7CGoHKt0m9PSRtGDN4J6wLDNDqhb
qxiPZJRkj8vsVy7HcZTd36DLdYlIigPxhKtVOAN6KvrpKV4eEgqfEE9TgnKjsmVF
Q169JUuidURQ1GIEHA5PFYWLDdBlDAWxuJss+TsaYLYDVShG2f1JIg4qwXoqqIho
jdu8Wwxz5M8pFwsUpD8SetN5z3BOlw1cI34nDkMwqe1Zltgw+xh2MjIU/cK5MZ5s
wjL6nAEdBNVWpGXtWW+O/ilZ7i/rEz57Uco6vmDIGQ+Lg8/i89H0tz7Rwpe+M4YO
mr/YpMhTlRayKeCax5f9oOO4R+DAeEr8HS5ot4KXa2NMUHiZCCEOKb0qb9tjlzEl
Xa6P8Z8bI826l1JtS3Dn3Y+M5mDDWoTydBQ2zIaucGV4aUb6JZRwBuiR58Ac34f+
jeT5EDIQIiYM1LqQRKnIOs2q1czyoj+KR07SjFWtC1+DsrDK+n4SlVZ1Ff7Vh8nS
It8unMBY2a3tEHWZjzGuvvjurvj1ASqQSjTeCmdDE0O2nGc4KCHAT5dJC4DR2CpA
hFZn/HWTM8Z+X+ho2gig/89tn066+bJaJJyLE1Q7ATXDWovqdt27TjbATcM5iext
qKxWHeY0qVquzNc83+AYF8cwQqPOY26FkRrU+lfk4xb1RfaOUN9lmsqEkWGJ7sAX
D9ZVMt1PKJ7SgTCaftpjEbiZ/DlyP8TNbFOqDbC7sE+tTwjqPgsSeyZcQCAQx0Zd
/krq814hp3mHJbJfnkf/xYwYZJ8k3pj5Jfz8fpEjlTJpQqdopxWmWw/RlF6sGUHm
BYEeUt8FcPKEPJUlG+N8v7Cakhp0g4ihzPOX1QpAYxDnS5RQvMO3+3HmKuhW6P6E
zQ7VmE6s0pnY687ygrK9aJhZ5NtIyH2uHr1IDfBoP1Uu4HgOCH7yWGuJNpaHGU0c
z66jBjNxpW/V/F/M6RyUMDB7oaDwXm5pXwliNMrBJ0v/qYE6/lZqiXt0wSWh+tVK
L/owf8O/pDijUVyo0JCh5xL+ucp8YDyYctKbr1KaALUIfl+qTde7LWDWXQ1gWsLu
dMxKfSFfMq4d+yOaV4BcMj+VNUZ8todFRDYN/fKUAj5i5RcSm4oeBt7f39B94qyL
tFZnr3gO4wMF/6WYFB5iBA59cB4bcQFnbusOrPc4NERpiUjFXV0rLDYFMXUgN2WU
RIZGdCBRU+OTB60n7mdEDFpFmpeRYtKdamrkv5KFPXThk5BHwAgf/uGLhQzbLNKe
dl9RYyO0fJr9T/wqaZL1NbB2vaXdM+E9pkdBBcIs4gLe2Phb/A55YFzoSjrxbtla
Fl0E3rLwF17WejM+xF5R7+DMLpekluIj4sYDJRaLUlb4U0ymaeK3ZORohkpiob83
hvtaBomctdtgn7Z+FrYBzEdk0WRr77WgdmpQYfM+/8Bnq2bQ5lOcMJ+CYnRQUG8D
qOUJjnVMq8ydzmbN1Mgleu83FbFEszmjLX6kAiK8RK94eqWmpRyZ2rTWLIFnYmjT
O+/Ei7zyySnz26TcD5qo5CQbJ+uvxylS+hCJzS27uQJ8vdN2LslNPzwjSpJo0s85
ibPFKWJjdk91UwGSNgUEWiCJ6fyk7Xob5vU5pyOKSFzUHRP2Y1Oscj5snUF/EEC1
GdXAWpN2/JjYOx8fHmUHGtZWxRN1yYB+v51apixL65F78NpXzH2EF0l8NLtFqg1Q
ORTpKqaz6KxMGWnB5vGUc40lH6ICjnP2zsJlmd6ZufVh6RQX5cfjlNSOZJ/P3lEN
CqWNxHxB1jQGcFAag+RK1NF6fzcOS0ybOcLkgz4GEf1yleTLG1A9EJapoRfYnrL5
97uljQSgXz/GEcmtatEXFcDRrdNs2yKg6dD+DM/6eiC2+YrlGMk9kD+J0hF45u5p
NWputQ8eE8w681kZ6BxnTZAh9QSaQuvpk3kfirHsj30PnbPntLtlGWTB2URZWbs7
njhSq4yCWXYUYE7H1ibubyKS0WlPV/CmqVvbcTegdTazOtgafwZvijx3VWUiLIyP
K010qqhLa2U26ZvrPj82h3KukdPRNv2DZyNZwPZBiSa0EcbgKZWmmZKpi9Sw/mmT
Yc1deOfosanEEycwsv94Lx3SkVNua05lo+8WZT98L4ECal7goXkiZFYQKwNcP4ce
hZt81FDK2LTjvTQ4X9N2tWc/OaXlfVI4psvOzhaIZsOZKEqecD30hlNazs2IsoEz
00jUOwsALFGsKs42aODd7JY5WIPuhcPPEsOMXF1lEomD2GOZjnzsk/TVOo0TC8Jd
a4xPWjiT7gnw7JXqUZm9OZ/1DPU3oHbyxU2TEKfUWZeFKm4EmXl/8JPjh+ibdcKy
hDjy0Xsz5seekMSIa7NclGMU90RwIVixI6Yw/GOcIXbe/LF485wX73tstww9ef6u
4wdEjdLwHepFsi+jpa9+JnO0SnrG4B67nbywqCAl07esQzo/r5X8Qw5/KKJOaHBX
Tr5kuJglWiUShI1/nEZhAynXlEPHqF4XxNRNTQ7DfiTBFoa5uLHPNpw63j5aB143
SXzmw1yTydcdw6nKabvLYKf6QgZGT4LHxld3UfriET5W0SJ+ySmlY8BDYBW83bXe
1Wv61zzJQi8I2GNfRXP+MaZ9kyEnHha6vZb4OXWZCRe2lsfyGFsrHFdSho++eGv0
F9u04GXKJOs1QBuQUeprOOsqliMuLP4A2dPu5iY7bxmX7GmeEypZmkbiOF9rQ0er
pwzO1oISTyR+BdaGkEm3sIKXDMypCzeQSByvieLLrxe3hXGaZP9OW5FW0RhjvEuD
VwGL6rg/ynMbwtOX8tXVK2GvCKjA+G4lBlawkgiKj3qtpqw/n5L2kcb+mgiF8qcb
TZV8uI3pAZzaiO+mVPQV3fPVyfsqWKMpAMZrWrlBSMDYmGIV9a9xkcNHkdX7qhqg
muZKx3CrSFH1R2Y0YnwGlmcO8MJe4A4fOQmah3Wn3y39NtiW8AUFqbwLP4eKwMzx
H4x4Wm2zSKW2/7Yjzqf2gVvKw9HnrKN+UDiWtXSXiFPiGCnA/lilyoVaoBjYfYJx
qQixGSya3aRCkR8d7NnMbz8RLHfsH4MXop+omzLOxl2RN2+xxRN3fso9rUyjKfLf
U7kPnygr/9dKYjyOO2IL/GTUbdMb6Y2XexRyLmvbGbmjUZI1wtRCf2jMucCePb4I
B2TxTvbhtXllVSELVMKLA0F+iEyi9gDPkd64mDxC0PjeEc1vek0BKWSom6FCSywi
XveYfAgw/bMLrUnccbZ59ZlpELrf1aTvaIpcBNaWbdoBm4QTjxxxqocGPbStVlx+
vUjRYk+P1OVtEjNYKyV2pdT9g1yaDwqVcpS7m5GBBpyk2Yna9TJ9HcE0PeyryPwo
o1q7HOKwhzY/qEFPzO/8SlTWduMzx0UfSFz+0WU/+MKGUD2hO999kCJ9wTZfy/9m
2D36h+BLmIRSqhxYM7db5L9Cw2Rgy4+aa4ZU7TuVo9dAt074tllyZPooosjMb+b+
8QQ2JudPKli75fbgrrCBY/xEAOBV6/JKGMUjKSORPjuvEvAsCGOkcy0St2m9T1UI
17FWcsc7OM6T0ig/dTftHKSA9Nt0mGfOLGjxnCrsiLdBn7ApdZ702GZt9CJxid3l
pDXYJBWmboRc9IP+pNKAfXx0Ict/Dmy/5S3djBvldiUmLk7x5brqW+WD0aaxZ2Lz
PeC/yEDmBdjkHE8RD/Bt7wWbbiAXhUdEpSHibbam+rzc8kqJNp7JUrAZxlP2igwx
HsWFuvvHXTnW9AreHWjM74IqZFe5RuGDyjZ8UvQiJD77X/5OyLxeuQIU3y97ZabN
kNVVfvRrIxFUtXqn0uaSU1QHcivmaRDnhAo3ntKKuTBg2xnTEF+nYbHV599Rb/Sm
ohhvsGWjuesdBzGUoE8aoS+A9SxFKNzdqsDbqZfQHUWHTyuiZNHkIY/Djcs+1bSm
PjUT5Q9IGF09K/++tokmu4qacFXkIrJIvXC5ZzdkCcrdtX/aSbMHDXGixvB/TgsP
hOr7Zg0GsCVRHolBZ2+YOzr0DD4PJzVH1oldUjWqsSfKPJuXhoOP50rI5ESKLkqi
CBH8V6NYn9hZhO5ijd/kw7X3gGsFHk+H54ROEPsMHYwrWETUUuI+zH0uIhgt+/Ie
Dkr7KtnozV8qLk8sAc6XTjrSNo45J4UNb3QCx3jfE0ghRy+l1zPIYskrC7K02E9V
79F3GqTbCAS2d3OybUeLgD6tzH63kPlIjQ06y7sqEwEmDV1hlrsI75YbgC2RJPUK
Q5tzGS6y08E3sYvtbMUN0dW0ICKBh8Xydqlp+FfaRhOoBQnDIItO9rdBdgZrevTe
3k1iaHrjX6HmVHXUzadsf/E3dtVzxhdW88FnGZAc+gJTYFN7mBMah8BaO0xNXQ6M
QC88QuddiGMvuI6GewZHG2H/1sqtSdaxhIFKvGAkebygian8Gm5DC+Hhq4+X2doH
fvJPT7z6wOGljdn2kkGs3mVqnik1k6W4DFR8rr2YgzUuv/gYPK3VZwNSx/zsduNN
k/em76OkFXuPWi0uFHkei2SLj+WB2F7lweZuNlrv/FUQCsn8xXElC8hC0anBootK
1YsHdQqCSoVIAjo2dqFqJbZ8PkExz7wf0jey8fWv/jNl44lVoWWlkqEGZH2C872N
3CSBXEiGGqhQ501LQIsYPM2WvxTb3wEnKEF4x/bbt5qm6mD74WW6TJOvvpUb06pf
ywxy/AUAZc+6MFLSCkyaX6yvSMauGR8PGlgE9HA6akVGUPll4IMpebXTuTQ6PRjY
InTM8UXITPa3MM/HYo2lUF8cinn5nMVifsddLPTSTcZXk++Zn+9AMAleJmsmGKwr
46n7dg8SxIPAo2vyAjMY2jLRT951SXKeHQPrgn2jkU20DOqhcFFtrWaec7xxAHeA
lrTwEqnV5vBzVQxeJKSTI557kURNGaYH5XeJRS6UeNoYQ4mC7jLXsyWJNwVyuPmV
dNSutZd+xXYP2YEhhPv0OgSH0NHUTgisBxXLAwc3K/vxVO+qNjSfbEkhV4uMr0ys
vEgnD5G50s8mb4YOWRJ2EEqqmYOwwraXEifcmZoUrfWr8SsSB8w9qx+oH252LKDc
3XsghOv8tnxjAF64VdhWpeiQ2wbxFCpn/g0UeZeuUPsOQ6Tuko/uwHylvMDKwfY9
BjUgg3s8ygUwcWMyToZdZPKp6LKI+dwN4vaXgvzRfTpD1Nz/D8kJNcdst4fKSelb
gtENYEygsjtSjHyW2p9r9reUPAzG5FEVWR2NSJQPluSaa3Qd5/GRm86i0XxNeFAH
ulJydVHbPe27T/vGhnb1TivtQH5OzQFSyTQ5F0Cu+BTZ57mlB0imwPynCD4ASMlj
V/LBBrn30wu1YMaJyaoq3qAM9HcHtKOvoVoGUHhrD+RBs4h9KjBAwmkxmQoPl8jl
d/9/ZXEr2avxOKQceJKBJNlt9XCW6KVgzkVclVROnDbgdmGY0W52hMI3ePySylBX
tcQLZ0WlHWBwwvdhPd0niJM6C6INNM2ItoPdd1t4BXU1/VpCJjeZdc/JsdrfLXL5
UZqg02fLFs3Idai0C7dZGFtIJSrmjOIhVVt/sD87+tazi0OVgDQiA88N0bclOMQq
C0h5QGRgLyxLE73rOT7sNmrB10xTiv1JMH4qpytLTeaOapf61ljcRuW27odiRPYU
HXW582cEX7sHw7TGF20Tr0nzzQkmdS9YDwzORVNj0iT8E3QIOCTUiXuOxWuAuSaC
dvA+/wIBfFXUvQfmVCrJVsIyKttzG6x6aKMMxxfRBPQDINaVussTGQ6y8a9aQ5R2
WMbiTY0DHHrd4o7Fo/f3RQa5CEF3GSY0ppHt0YOXgZzUOEt1ur1YGO324rFRTDIl
W+Mr+l4wq3M6Got9wU5UcUPMFNEueRRGKXmHRAhC1n+6gwARhpxBe9To5Iq6YDq+
1HXqHXiDTvBqvW2HOnQxiMR5d0w2vrfyqLG3KHus7t8E6NyRnD9sByNQRlKNbZ/o
K7vioGmeALtVUpg9uuoaAAd2PxVNO6rjxRPR9KViNT87uyJKjarzWnUKXmmeNYAm
kpJ2YUP9jBJI3pFwF+pdYYqM/DjreNLUwiXH/yoItEqvy8iRhsVaXq23cvNlxz8D
l0+icGbJvTLzZutR5eWtdmXVlm/UUyqlYIOCpZzHjBMTxy/FfJIjirz8Rwmuv5kh
rVbSIpNQyVxY0gS5Ai+u82j+PIzwkqAHzjSWQ+0/y18yzBLCPFr2UKzPF1WyDECl
OwBlFsQ/L453nTj+dwX1cFZo4FIlmoANmAtEDoUCYSSNAnxrXj80A2/HU3lZj6Ey
enA8E8Auqsk+rkF5LAOTIRMyga9PltflfQAHeXvTSEGUlRClCFg+g+kX5e2Nw/Uh
lS7fX8WVt46Dos+uhXZouBM7vd0dcS83fkbV1AbYqSklWN5hPhBPB+6yKiEg08pA
8//c1JN0Q4xrJI5EDjv4UHIBKhPXLhNGHTDQHsP/GW1emfGvbPDTMm1zTye/HflJ
Bi/a11NpxbIZkIESC5uBzTNUEwOJZhkSErRG8F9N0UhTX/eabuyjE+IwEsMyxAgB
nWd4+01gFX9JUhu0BZIOQNrGZzfh2s5jJZs9TIRyQJcOIdG8NNf1NeQw5QzlbGZP
3v6ZfzemG7tkh8D4oDkZ2vRkWdXAgxkPLzyAD4d05ZXmC4a9NWLPt8I0bAmLFOn2
x3pEkpBbeq+OhQ6udfSo3IDw/8xUYqDhfc5bCw5XI6BNXT1PbXsrWqQYpPgku+7G
yKF2OMeK6Yrqi/MM9CuLCdLtc31qyzkB2RXeRpIZCwGVvc8Yw95AzLdxhrUH/4cf
G2LxaGQQB1gwjqKS+sYr6fzVilbWDxdDiYcmEYjoAkEuaL3MAmDznld0ncX7lFaN
UjRhaNx/meFBkmuqmf2Rn9xWLvJvyDTa6Oda/NixjwV2cv6juXw2O6YyThI3iLhE
SJYGS+MU0TTMW4z114kwlVp9DaI2KNap9cypJa+JGJyc7X2Bj7bdf2dC5uCWCyRn
903yMs1koeeD8cbr4p75Hnv0PrQb3kxcTpAvOFAHGPfvZ+8/klJ8/rqfomA9DfRB
n9VOHmIwdyin5tYkkRo/caobaFFWj8E1QrQQ7lK7OllxCQKJilAClLeUm9Be1fSv
NUz1Jqa1wxjuWxTyQ5SSPJVZcSo9q80s9Kg2g3x0rbNwnnRDbwfkutc3x9EltLQJ
n3R5jmbGeZ7uDgxxNkFUYiTn8/iNinWYzgxB/XIfqGTo6rNAaliFlu6FieQyZeat
vl8X9y1F8R+uLpIRHCwAmE7GWOuvVqUcpqqqlWNXbydsyQuyj0zi6uVjt/FMjvJf
DP5tBE/h6DLGwi+aUw62gvlHzyVvpp1w6OvER1C0mtzeKmXJSG66FKDP0Q55TWrq
F3nNLXnlc4odDnLTURmD/XRZZ2RKSTvHRuawgpPuBWY4sx0KowUwqoygc38vQuvU
Lc9EtBipWO7DZhGwPIZEhTn52t2i1e5Q4zq/d68iFTpNIMTPy9d45OF04YfWG/rK
XsdPt2HwYs8YI1lP0FD22nhUbiuP+eWE8g6oONCR3rRC/d0kE8dYG0VCbuV4Jk3t
lsrPwayDcA/Pkp11hqPjreh/M5eS1mtKAN+BZG/qaPM//wX/0BZ53m4F/VVsdcgM
N9WsZC8q7GGpTz5Oii94ha+EuTwiMPD442fmDC2EeSy78LTkEGueMJlfTbV8nnpK
ebmkNc5FoPNqA5X7sMMrAtEcv9Wi91WuFXzjSLKGXPCpaG0f6Tq7eMA54BmByNYH
M3Suej7BFRnc8UHaIdAI3ePQMeKmrhXz9iga2iHAI3YfE0RNsWJcviSUr/1qF5kr
L9590t6CK0Rvep28J6HKpYaXBZaswFLGZQzkfA9ULiXgF8Ake85qwjsOZLfmjVA6
XgvUngBuuveSRpxbPt0y6guLdb1k9oKbuR5BGV3mAmx8mOZfRIM1zOIAStRidEWa
0qPDWXTjh+1aDPH6U6jVDPIPg7lXMxn/cl/L7BPAc7eOM0RnIErLOu7ppHDqyVUV
gRU8BgI7zctoNHEEDueVceEllNCWhtIzAX916g/liu5SS4DtntayzGKYx2P0+2g7
Zv4yvYxCGglDzR3wzhYuAwWeLHzQ7MBQUWZ8dUr9XuRGUUI++bCqGQWDS8m+8bf7
sTGnLLLDbNJP34cUYAdjNRYDWiVrfLS8rT6MXSxzcvFph8YG35PI6swhQdjCkkyo
3WczvqYnnPoCN1pAGIXlqp6pc1EWLeo5X/lGDkcqNaFS/QUN1XeY5OCPLfqeBgLE
9MJ78C6/zlLcSzsGKx9aDArdTytVOqfZ0tCcCDJfcp/iwc0NKX0JCOKOZSrwgmvt
855KvyBWVzeqkbX80/NJofdatgJTFR+A54cGN3laW8pAD9m9ZhQsbqk9P85+jIrQ
trRT2i9qTG+sFojNrKLvCl5ad1QDzrtYJEGKw8qrlu6vb0/ipYUWwV6MySMtX10C
jn0pM1ySxV3Wb3/z8WNPSRDxaUkEIRSKMz4VD2TxHYVIpV16nZOKeSslQoQcxrU1
G+4Ti7DFvatuQ8J60c/Uo+KtiPeFZObST7YL6bRGLg+ghbaySqw7f8Jr1gR7UbJD
ICu2fOoVy+crpKkCS66a2FV7QKt3oaa3bTBlQOBKhG/Wg8Wh17TfiDPckdhPJaGf
1t+JOl+IiIL6t7SG8mTvaBvTDjr6mlSwKBj1/hDRffXP66rUVzaNp1U1eav1Kfi/
Q80kqerFSZ0JE1XU81p8y7TnVo9VlFZ58E8yTLV5KVOwAXdPtBWYVnpj/2CZfjS9
fGjmVhASTslYy4HbfGtymME2cz2rvgHslJ3RfodM+Q19vh07j2+JcmLo10b1Q199
4uqFMph09HiBXCXPpQFuOJMGpRI30lgn1OaTXQG12HBJtwb8nJ+gRDm4jMYCqNr5
9m1BUd6FJy5u85KRSb26fDit+oq3o4s4w0PgJwzYQOfLQ5zzWbcgAtoLEDuV7IU+
W9QCnLtTUYOr+48++ffaujHE/VS2ZRPuY1YRwcT1qKz0/uuty5o4jx58U7N/ktna
7rl5AVKVtGr8DSkUojDJfRSaB7UAmV29otaDq2Mwdi3ZeUUs/CCDgQbwk4vzX9Rh
5vS034LF9JWjojDmanjBOu4Xz8VnRfeWb8wWOHcYxMhtLGgadjNARpCDlfqy3xsj
Vt4D5ArWRJlNJNTF1uUHhMhR+FEVZpznaovLjFQgysyR44WBLjYQhP063jNmbAas
3nJ3VvjdU3ah8XSFUl41bP9gSnjoAxzZH09USTJPEUj6nKCzlFmCYFna+T6GevGO
I8yiUsGwVkOPth0AdIVVF4HwzCD6hEZr02I4S0OOxXehkR8JXmwItKgaN5mhj2Wa
za6brEoKkes0lnn3VImWeUkmw+Tfiw0LxVa4siQ4AVceLAEHP//9NvQK9ghVVIwW
bdggFuOKWqpkfYX36eZ5gGB+gw/xzG4Dk7m+TKXhCnh+XBY2A2phzuvVMRCpaGmC
JN4TXZFb70if8mazRhNpNTh5OvxuaZB2ZBrEP9wWHcMF/1z853csWtXfvzOtiyUC
o3ztmlVGR1YM0qD4//liCXbbkTEvbSPcscj4eQo8TQpm7d5lXAc5JoLi8bLvEmk+
iHquqWyuvvnBExPFzNVj1agIXb6mPgcb4DiUfJYx+y3vLnW/6B6XCURtazR5RSoU
7GyGvEQ/TXJ4NROQkKUvnp7TcRf4JLUqTW73fDot8oA4aoMA41WmvA3lTv2nQFKD
/wrcDkY6Fhy3hMJEf5oXrwvwb6p/KxDhodM7djCWIWCz654UtUeR93Png7t/B0tU
AJ/74V95h/llmwQE9Du1cfNG94cFxUjhUI4N3T3ondTL0dn+NhKJb1VGVvzWi5aQ
m3tDqR9b+MUxE19rQSM6QeR/jgZmlrnoCJyFeLvlhFUF9DJame1l9vkJuC78FS9l
OyWKpmqInTD42EqdFOBl3344Hhg/8TmqwEz50t6aIRCEDC4RGWQculXBpw3eyt0f
ueO9oliQ6+iPph68ZI+fQqB1ngfnuC21Dn8gKmtvDZrRmnVoPPBlTWJgR5eVtf9y
e4a8IHPSxgb+fA/gHyhJ1xU+jDmGaZ4ACmoUkHAGZ42O+NQFkuK9RQoIVVumTnIR
sLlNFj5CbH1krHEWjhmg+VXHxLTo7IwjK/Yh5XGsat0sOxTbP9kuW0gWhHUkF3Qi
JDYENMf+paKoA0ypHPcYWzg5c6nO4RDsz95fYEHUmXr3XWP1E+01YoUwCLswOUX+
NVk8sW6n3ZKQfXa40nJh2phTV/qPvBFc0LBVveLd+j0zetP7lO2qzlmdU3zg6xtE
OGcSEgrmIRukzVAND9mCv4b1REdlXmZfe48JdX6pHLuoXjuHJ/HNVEh/FVHNiNCA
KS+g3jbnmbHgPyyQy+rIc1aCei76JubUZiYTbnNhBEJ9vZ0FK7Xam9Mrv62+VXG4
tduXSN5fp0fU6sLJkiNdLu7YdQ8LH8NDCPTaC8f1H5+cRkNPJaiqt+/oK2TlTv3c
0TZdBFOhRVS32EilLIzuU4/9rldzh+NhyJacVpMh5EbaNXiSsHIT1KJLTLHJuM29
Rl2o/raqaavWtT50hU2vXaMEyRk7rb+/PlwRiYPY5Lds89Av1LaKB/g5Voo63usa
jdiyW8iokws+iv95Jl/IAQirBSZxzmc20wxUQPbuxscAmPvdJpQHeAuL33I3SNmZ
6ZJc9a5w9XV0RJIHzUMalGGJcFxmLjl2G2UQIzv8Gx4VrOleqa4bb+fT59vWHHFi
+ywVnO5dR6hsEHZ8TiXDaIuDsRcjmkKXDayN9LfL9DJ7dInnm9lpqpkmLRqfQcRe
asI4ns7GCVcdisGOX1UailAgakzolwBapRvuRg7P4b32IHOAZpTw4DxJCLsVbY7X
7tdvpfPcEkM3cVW7jV326ROaOdsTj4wUUlj69o4e1hli9laDuhwAeR4Al1RhokBj
fvUIouyx905Q7EoeHu2OqTJaoRI9g/dXzD7fhOQ0wvFFVgXTPQN2jeQAiresGbeL
bjLWgyXri0KjZ25pzXITru8KhhKchMLWVztgPrsycapcfZ/gGLENDnBUSEAavQQZ
kwH7RW1iagqaj5cWk0ECJzgyOHIM3UpsZBmyKS726J7hSmi6UsTlhZKFDU9AcdjY
L7LASNo3MGytvL/oeEHK368C/CPujObokdrkwg74dHCgRz4jWbnkoMJBd7GBI9Ig
IwT/QffNqWuKN96e4C3lwqO35ZPzffbhLH5FaSvvLuQXq0fPDQmgp/9CNqmABMDn
TjkHwg4ll22voFCJHvW4s7O+fu7gH3n4TIHxTcBpP6r6pa44a9EvqaaBWEik+B5x
IpuJf+6GbNRoU0RYMQu+kIZHmM9y7GAp7EP1RDYsCDCi1Kx2rJ8mdviMPGxGjSRy
844sO92ImbguzVc+3A9KdbmHM91JBuZy7EVntXgsLRcvmKlQ2VKUHrjrNjIJGi03
7sdHOqXI/ABLd8dgNgiU/k6xaNmiCA4VNshZiXst7/qfkjsGqiWScEyo3S3FHkCg
hqrViFWs8j9PDBp27swthywcgMcY/sIPtLYDPMcKpdzBE54hkIVjIJSwWB6nwWtR
6F345QLRyfqwr8aTo3vtm4HwhcdYMPOHJIGWrHIZHP2mP1OmS2Rd+M5V1tx8n8xp
SwrFR0Jyk1GPfp5vsLodacwT/OflWx1J4HZ8AsFC+eZ6jEgf4lcawzzDmjkYGzYJ
AwKEgxhwLWfZTYC4aDz8b5UQXmNSkvjMyNgWD1GiP/HAU7gFmSGxTeO4Of89RqhE
+bhfZOHautf/bETnsW5q8L0+gejjYP1o21rmbfLY0zg6WyifQIpdFqPrPk5K9zbV
/DTdVYMHyTfhrlhw+DwzZi8I8XFlBZjcxFfPRtZO14XXbjhp33Q83OD1ViZ3qFyy
n5wbILYoNSqpiAjppQ9a1iiAsjGQ2wfTK8KbAIpjAJNoocMhrPkG02+nB4cvq8RA
HkUcI91g7/sNGx+f0JMtnnIybVzVHOerrKJ8ShRwKA2id8s6p4JEJ7ioR7bytFV4
WvF1wKQyDQjPI76+iGbptgU9eDJJIuAFBsjmsNJoIlVOlHFC1JWvSLJ/6YVcuLTt
LoaFfz6dMe9/ehp9P/VjICBb79nYfs9JoslgfrLn9Se7n3y41J1U9d1jaVTLpa+Z
r6RgZUj87z/nZhrG3jinABOPc9Ji/fKzibar5E1SChp2b7adG5+c77MA+VkVArv5
4BlvHRVX38Stw9mRA7nfQwcIheWG+jJjBzijZ3r2Iq2K5kgKB8C3YIvi/us0P+XX
yPwnhxfgLEzzGHYJrG4lM/wCb2KHtLBDwrFoIyY9hR4FSpvY+bEj9nckgcImw3/f
dV67bv0jngqKJLUyKF5Qz2h0wIAZya1JHPo/i4R6NLPzLoIhYF0v2IIF7HBVtrVf
HsuWmZEvNMAQkFrll7l1MGXJ1uzU+eQNm6bNfrWyWUpcmu2IphhgQe/VlZYV1Bw2
oXZ2cV0zgFwt1lGW/2Bc5entTzJBTwBmL/LDfS38lPRCT1Ffe1E+t3vojqYidrBG
6n0XnMi0PsG7gk3C+3i58kVP23UpWvJC6LMt3h3sumFMGgjL6oDcMdNLSYNelpxm
SU65Od+0r+fRDHqeBxJhnTs9Ag/3Z0uVfpMjNe03CKq02Mky0n/gf4/nXQWcbJ6X
9H50lYpkAEAyqQWytlQk8iYWnQO/JWkrfair+aktv9aDUKXIP1E1ZKfpGT6izmHT
vmZMiRCKs/NKHXUICq68yLLUXHFRFo3WlLxiJs6v/Q9yuOIB66iKYD9W73IitTMa
Ynd5vjfRAXDh+3oOIfMEyeYYNdnBiF1dLiStGn/I4yWbHx1aSQWBTZVa0HAIlWot
nNVSKLhdDd8bODPtLaeimLMTFdhJ1NKX3lRvwt4UK/6u7m3uQznWZz3WvZdeBjdu
j618S4ouuQk6emLHAV//VXwe2ZajtUn+LKu7pTWhoWoW12HozO1oTbm7empqQgeW
EudW8Ciy/w94ZAox7jNwC8uQf1E3oJ5ySzO1U/GRNYNscDjuHQWndt1+0b1HqAYb
gat8NvVmQ1eYfbEa35+c3RIdZ63TUmnq+uiHlwS+3En2iEJuwE/oicay8oVmz/Pf
WJywLErUUZYngLS9gUQWj/pw8+tm5OyCgWH7zh6kswp7ldyGAQvU214r0JObvtNS
PTAdmI+GFhyOfupbym5z/r1YVXcqWXVV8EqBrAlOYUbKHR/Lr24gPIfWfYIEwQ5P
MVqGUx6cLOTYS4261vojsARR6oPSDN/XexVuw2YRyTIJYrPjjQEd6YUaXSDb9CW/
M+bjkfsi5zUS1qsv+G98NXht3rGLgXzib/n8G0kJv3/jR+cfW706zaRVIvQSZspA
WJ65Ogrt1GvUwEbPxGDGmT9L5lqrBaVs/gluPZJgy7NbfAj7XMoXg5F7Sz3Av9h6
ZeZE5CwzAHGDu7pkVgstsnRJfyr6MjTxxisV0hGZAuIkqwSj9aGAJKVL/1p4XIpQ
EB08nd8uH4lWpvkiYcLMpMm0rcnwi2anTqdXqDcjtV8hpVNDhynccEbTLFrJHrYL
VJCmCWnncFylL7Ph+xpQv9C8BhV8152StZoZvgyHGi5IU23iz6l96BcC5pYO8wm9
ePjyq+4kzd4U4GMX0YXYEFzfRR77wxJOCyDsW0GK8RqpJ6yLsiDNvoPDSA8Ufqa2
jlBADLf3ICtBtFdsgI20p23JyEm+ZBmHFBlflAggfrQ4UCdG8FKn0lhhfVF8y25c
lc6PNkh2PiRbBbZcnwOChqym5AEYBPC0JZNKj8lSl5EUjBoUw/jqRmf1P9BhYfWS
xSpZkY6rfKjrgdvhOivkydMWlprd2PvQSuwCTcEoh0ggZOgRZ4Dynj0plu8BiE3L
IQFJAmLh6ZGkq9iqrU5hGV547qGgv8sJV5XHtaxVTvLGoXEdXj4QUk7KjLxjWdwO
cPdwgCRJHaqi78QVHrKyQBmxuTFo7zx5RChQWcgHJmKccRSxQNEZnInGjFtcupSZ
Pgj9Cg5fiTAjHEncLYk4gKmdmxxQp01F8tBCcXR1PmUSGWDtK0q9jqAwdP39qaQY
auP1OKXnjJZiGeaDwX/OVuOHE3I3oqJwB5kMc1VUuOkm8LauTrFXq3+jBeK+dV8g
7hFHctmm/ZVZyqDg7iVF8MuLqhzG6rRECsDGqfJ3ecJBzO6VmVumsOJ7nmrAEiBt
s3RHlR//uoI9VXnjcI79FLk7S16bWk9gfWMLIRCLbkDGHi1nrmN96WnhqCXuhDZz
DY7GjRZh3g/wKTZbU6p3XatbbdD8WuJ15nKC89Nlyesxk3aNtLv/TtuVKFjjTcCJ
MrD88ejOyTU8EYM6nx98/RwwvZfqd2nQ58qx0Zi9K9uCO9ih9U1ZqjB6unxWLixC
Y2hPvts/lDlFMaFJ/O2tVxrZdVfRpi9VkbNedV7Qsa0bkryYMq+tzVA48Jx8+5Jo
B3W5CgNHs8c0WRy+qvYXFSXgj0MBDBEKqV7/j9apUTXZV3PosDIaK9gF3i4mfvGF
EazMEAjuAS5pJehVe0XnsEc+AoXQTeOm0abuCxFwjJaH3+SU0VxyFbF47r4w8L70
neHls7UFaxwBQccnsrnRuWL+G8ayC+qvED2rJwv/sdBoc/ZKJo5qIChlCtFsVSeJ
MxqCHr4TvcAsZw+uUrV86n2PTJoZdN1ICWMSTPBzElYf4VYWRaym5OnefBgddPV7
MA9DMg0k1SIN/qLuPcXo+N9hALIAgA6NtREWiTC17p2y1j+mmPVNe0ZLEnD69PjJ
Y8gMZitemAmZLlciTa3IRYMxNYrmlcBoc2GCBDDQ9lR66jfRgjegBzfQq1umyKKM
C5gfWDFhFw7ce2C8bcJd6A61vD4s/lZOfbp7I+WeOJBG6KAABKq1EUArCDNNlqOm
qtk5V9T9+KfUY9FmgrI8dofUKwxMG9aIogPoNttMRyvPE50gkAaE9Zd3k6jM3ZY9
vnaDRiw2Lm6XzQKsApt16hHe5r8WHUNNVBBOXMFwVpu5aMh1Mwqgs9rZG62gyGkV
Go+evyU3aKekpPT7DKzPOcwVmuC/Ucl1Q+1bYx6Wa7nunb1i7sZWrzQReg5nGs6z
q5a+kWc4ah/n0oq/ICZNpKeHVsPABDbvWHDJbgZgbqypskr02l6j/NiaUMPeLwfK
CQQVqHmQFCcmEXEoPHGaq4InhX/ioOgdX50hWGGZnz/VLu6LS4kEOt6hO5PjO7nZ
2y78x1NIOgmq6BFb/cAk9otvk+s5KfxZuZRxRSUypkuNMcxzPPVMe0+s5BcoaeCT
J82hj4J2JGLgZPGPnlrDMmvt8lo0Dq6/NXzBjFXxC+q4FhcIzgJje4YzMclYPskT
jvBFWEcBsi40WEN9carJPXo8Mt6XCBB+Gs777fOyCb/soSct+t2KVNfDNX7WtQpM
i37ZTuL9bFe4Jsh30i5/HhNcaRpovy6jm2ivzTApAFlEtcEAT9fZ7M707ZRYN4XK
pb8rBcEHgx91u8SdWMp+//ldm5yhExNHqd58VC0b4N4BSes4pM073LzBykWrR/t2
8YLNaITjSRtUx1GVf8cV9hguPNfpyh17EHwisRS/fRroQ0ZVkL1txRwOQURYQPMJ
YqXLn0hB8EcJ2JHjxT3/n/1CitRi3S7PsBUx9pT13QywML/P/JAhJn+LasxtsZyP
dA4CouFJieOiM75LvOceUx7uzjPQ+NHPiLhBBFijRNGWOKHntTXFGKzqL4sZw5Y8
yVcj6rOP3hmMwoyeT8H+bEVb0anlDm287GjlKOXw8m5LWKzgt/MEgtF5F3+4mbtr
WLzsZMjyxgBopR5O9WwZrfMFgf1i9m28OB95S0ouJc4SxL16QYQGM0y9e5Uwqr8H
jBw5sme27szJ5uCmijFN2U4V2ogft3jzTKF5fbeaWKc2jzsSGSVZ9++U2ysCbe/T
7rn3DuiMbz0tuTKmr/bb8yop+G52g5nJAoEyjoEOSYDa4Om7nmVRcqhjD6CfSOb5
0F+DP7U9Az/Vy/KLsIAuRDD6HTKHuKA/NDuqKR+LRc92UAEOg41R+P32m1qklpwJ
dfjLMQBw8E9fDmevmmu8eP6rVu6PNI9ga/PrgTuIF8FmIJAOs2YmGqSAJ5NaamxO
cCU+gdCLe20ITNfm6ZP7M7z7ONPJLoxy1UTgBnXZq2HQtCGbi8D+olBeqNsrzDvx
/6ZnHCHwhAtDP7bO6x/EBu/wPi7f0JgCZgUTzsXHgzRNxDk7xQhMCG95mGYxNthG
3oSGVovV7ldNDaj9VTc9UEk9L4jVkAEnpmxW220tEM3dUBfR2fhPqwRU/TlT+Vy2
aXDWGsV574OQxdGVeVN85GvelPFXI++VsSiZ2P1R4cC2IUuGLdePJvFyQUuoUwr7
6i0rxZT59oNVCNS2Bipl1R8OQH/QbnFbdVL3Z4WBa1hNQXPXYeNvqs8Z0DBlck/T
fBt7h9TmfKvtuPChR3K8l1cclmmbZk9CQkxKd1PSC/6111Wo2Of1G/UYaMZ+oITn
UuoTEyIWcjX/yhSsntkLY030nDSBcRi1w0toefb+Ehp1bFv+4+dK0zc4jW4/hp1p
+xOvJpbMhnHl2L1+DrJRmDq2ZrTnW2ryYbqTwPJi3/qL9jma8NEEBBpdYB3pWBgw
jBCL5ggW7BDZUVfhjrYwPhviWtDiiR2Xa0uND73u6hd0Srjhewu1ie5Yt2Vste4Y
QP/PmWd+Jy/flIIdlw/rxOyt49CtEyO3EotzvBTMIaeixh/+UIwWg39Qk1sigfux
2IbZMZxiNv7y/mCKKrQTg+FGajQrMjOK0uRHV0gKGuh9NbCqGEAqyLSYBLJfQAuv
E6i63YgwhwRGxFkOBsDqRqa9r6u/POC550h+hWsczK558JJD44wthpNtsBXISTIF
bL/pyq7GqMNFNDQEk6vFP4gLa4NHqes4Y3otvEmWLr8Voz1CJSsAid1OAaCEZ56l
CyRNG91syOQZJdd9T2WrHdp1CNDch7z0pO0mo/IEh+D1yvJcBpJNq2Ocg57evduV
HNYuttdTKb+O8+gSQVoKsz8mI5NblBquxkzhsyY2EB31w+Eh6+t+a9UDoVnH/17f
c+h0h2C2B9FUT+zlLQkeUKfEEEdMwGZvZH4OKeOpil5vuZlJwPp6Jj+uT10AzKg8
FjCs3fvDobTlsPV4p9n83px6MXG1SU0Gr9EQdl/qDaRdHNOS86yGZpSf1D94Gt/h
tsyC3D8vwCUezf9SrVHZe3d2yze/OuCc3N6jNv3hd6TL6uZeVmTyfJ5hY+0wArcN
0HoyxbKsN5n0/VkKyu2tNe3hz1PWXqhAUAzLrrLd7pqkorWOmFcx8eN5BVh7qENI
Dp4wPYqID0KoJNk500f1mfkh6LoZxExzbXsLCJaP+PJuYHrUuwegmq41Kst6UWYZ
ZtSkulf8vfEZnot8de4qPaUbmcDGeMJWXplzxXsJg5+5XTe2Ugtcd1znNgCl2NsS
cD1UmRCIXb9mYq2qE7V/7naS94sjvlgnebL4uAD/A//fquA6hRSqSsyM1OBN/AwV
q3zxQkTwyh5OYfudlbVLdkRyy1pw+HLrlYMMfYzVKW+dS4ZaXK+T3oAwP97NPmeQ
pR65F0d+t+26APmQcd1mRZG2Iz7Rwnn8Q53xjm/aKFF1YyPYH9G7gv+/v9dlw7Vs
q5nDtKtvS7xj2f+AbtjySbEytlq69jIzKyT4EMrQre0X9q2Fg740RwVjm0cqu6sZ
I4xTXDqVGeTiNbdXrJvjXH7y759MhPwaVv3e73piI1PVTsOFN6gPxve/UdBcZxhn
VKwLP5s5Xy6Px2qUk63aAkSBDHXklpLHut6GeHzFuMqycQm/QYbGCIEDwws7MbGV
ESS3i3WYtOCKsILXCl/GotWGsDdTzoo1idIy1wJLFPRakueHunZ9JTL7WKoezKtI
+348NDiZ2MNg5WWSDsR0subZ/RTzOfACgv+FCyH625I41gvsxWbjXJp/lIAff7oo
zzUibzBkLEbRIgEiyuGK5Q40E2UJoORHzz+nOlG5Uz8wbFtm+ppfWRqh00FI0BBk
PKA0Gj/9O/YVvqYn47j9F05T4983QvtgFiaMQVEfzH0H+06PMjZi1z6GaLgch4d+
SW54X2i7owgUANVwvCe8nC3MpQref4e39DydAtjJ6IQ9sqNPifSiSLL7v3MLOnNA
AMRPOktb+BA2DZsYe+RQHUVPoC5jXA4V97FnMR5M3BrZM4COdjFHqAhnaYit4Dhr
DXwjheEbfVP2Hjd3e0Ov0cmjQgg8H7o7Lsew/7CHSDkszqaUzM4b3tF1v074X84/
0q76Wc91Qvg0lie9kaTu7yA5HWKYSRxJsuQOQoQd8Ht57eZFwCmtfxX+0vA5cani
w6dEmXb2NNT4q0k2KDdpnFw7O3VcdfJHoScbZuKr14KRxds0GWUNDylal59McUfY
0/cFXWNmQwslSlU6woDNk/1i1fwsCmU4tD5+85n8gIMGNIjf/peb8U1QyzW/leGX
+2m6hs4yOODMbBJdctibMAEu/nEuKmmz6BU6Sh4XSVKOPZLT5YBCm3/i4IbI0dBr
y/IMUsunwun6gVZxl3pqvQMFsya4GwuphDcPLCalSZj2s9FfRPBI53w1ddMHiSDj
OJE2Cv09AZ7vqnzSM6WdLn+zuz1vj46GXnyUqYgLpA6UxRZMFOKZadccQTWy9XlY
Zxt6wCFc5+Lt4hrYM38BjmYeOkZ/gYQJdEXHBse9ApwEr7W031Gc2h0Ru1LSI606
qHC7oFKIYp9eSsW7wqnQyOcGhxqI36+4f80N9CNebySzYx+u/NWTzd4f1L9BF2Kc
upqqjGqH6lYi6pogi/is8+qGAQ30GnsVAZfknY66AOE/yE68MrxQqyIerChgxv4k
uhy9llRP7VsZAbPAmlLVV9qRznrMs1WM2wdP3M4h/XPzCgfUcfIjFVkikvLscQ0s
uz74NjcvpmLCrCE2Mp6TjK+zVZAJVgzP/JF3bvH2Sw4qrieVQiw5CliS8poA9fwu
cz57ri+p8UZ5eRpWjaXCkPAIsbnA0erYZ4N7Gyw+PkBpwFK2EDW3Eze41zWJciwq
2/iuUbSNb6RvN0v6kAJYdGntJpvH2CoVloDCt6H7RY3tvb9YewYQ+UE4Iy/WmWUm
JozaKPuF4nlp3uChpgteJTmyILRcmqnDYGxydFat2VvY0QECTAg/ec7XMWt/YO10
5LqDudIIOaMFyVEqwWP+/N71WMwWQ9nAIVP3odQQ+d2soyMG8/hcVezpndsnyMFC
MccMig1Fss+Sqn/+yax5vun102+NfHqSclzBukTEaVdL7PDZUKbKkrVASaNaO0Ye
v/Pqi20S6TjAIjgTdF0+c3qFHTDtO6kerIemGtKKEhVl1TQMJFFUwD4Utvf4SyKZ
YwiARpXszPPXTpZhFUO23SUxHu28yx7N/mpoUR4gW28+rsQl1kWDeJRzoT/rDK2r
gyaITEEWWBv/ENTAgMVLGn4CInB6mXa+q1uV45wWgIUEc2NCW1s1Et7FZ15cvT5b
JFHIkBtn0fRdaQtJR5hMitswzXIUwfqUe6Qlbg3QX9MtVzRqbZZqzVKlfqq2YWw4
T4LcDbD4zDYjiRNuANfX1qmTjYPiTrgYFunjwVkCrA+pPNLuTE2wqatK5i1QE5km
Bw2ngU2UP06N8XddSIB1mu1ZYoyzPDOegt7tnsx3MIhZYcpYwKlb2EkXh3sHIFmS
RX34h4Sov5dssv1zEweGQqBY9IdZiG3+0RZQ5Z6yqV5hyM8EgSfYIgHegtC+gb29
OuxHV62xyW1mGE583vNIAfHDTPyVj58Y+o89K6TkyW6202Zgiix1LQdeCZQ0jBZF
GlT8szTBUoy+oHHk9L8ByR5s6g2wMt3lWU3katYB0um1yqCMCAIFmuFiUjLuIfEy
y4A8aBoJjEnU71z8UdCFVEDQ7DfisLQGoYcBacEtTmkbtNgpaEstfrLr1YU/6w8x
dFzWazlUDgW/UK+cKJ577O4A4LC4fgxh5Lnq1Pm2/WYk6qDEY/TV1W506bXtAo0m
cl0xwcMGau6WHvYLfRJsipYniZjNQD4YrbnJSogZkkCufh9kBlQsptwFijiXxeyz
mvGFtaWm6B6u8UKvb6gTMOEqBn+YWE2IMYt9xI18hqSXecZ4gY2YwI/ZVI9pno67
k9hYNI+wrpqI6I/roZ2yo3DErCoCGU2xipNJaBEy71DZpy39E6WVZTN7wh5mChPe
/4DCwrRoajA34UAg4Yu22CS0bBHQ1mACqMQYHW19mK0hANuS/xIs1uc43G30W6MB
+hWFfvvRvQRFvwxkh3rf7D7bFGNrgmE9sngQKYJTtFjO0l/wOOpwaEBjk2/mK5My
raCDHcd1l0sugN+mM8s6YRiHNA8WaEtApdiP6H3J4CoXVin3ewFs8pQwLNV/80IH
iSDJvrhQnWvP+LJQvQ7Z0HXjGorBjpTLIirWTo33OcE9fslFMunD5vclNdNGSGdp
9d3cFV4mpJWPqqFN73EfQcDhhLJ9mJh86dCIEkGz1NyRyY4zoprewpvhKyPrL3eW
vtrE5r8W2Injz8Edeig2tgboYRGOOk+wQrvBd9TXgSL1J54VhmReqi2xru0JTwbO
fScvA8hqtlQOnGcAzsf2FXyLJG9i5eaO+KpuwbwAGhy/zKhXWr+gcp+R3EVXx5Qy
lrCVypt4gAMqEnBtr3moaraDuDmwcdO0TruDcEzOvB5dqY6QmdxLYiDVd3t0yIaA
1UqLE/L4DswdwzTY92Ibr7Dluj4ttXKlVwu5vUZ53oqfw1DQ0Nk+25sUNelKSvO8
o6u9Pp9NsCdnEPwZCwn3zz/i6xPljaBL3JKPwMbM71vGz+guUndp2Tmy6DXZND5W
8rx+6H6o2B51tN/sNcFUYgrYEncBPgbvxDIp/mauQInpCmOeu+KIIoDyCC4mt3xi
iqYEV3KzNanDl0J0C7he8VUxZhYmqdU1Lm8fAgN0HWF8oQrKl5o8u9/txhD/24z0
mHjFGp3COR5OHpay5yo0xrEE47NB5oF+o4MIDvGod0ERYE+Q9envm9ql7bwXvMou
q28vVy4m9vdWn3BgbV9JPjWiRx7WkAmlCyq7Isfh5QNa0cFdy6/NlW3kuMtPmGQ2
+YBE9a+hudjBQUyRuSSR52l+zGsHcdndBBjahyFPON9OTEy20AFHMDCWSlnl6oHt
zoMZOhbdYmspXD2IRR4vdciUTZDYgWCaTnuKQPYthmh5GJcZBaO23RzcBRTad7Uy
EPTsOi6EvPdPZSELG2DeDhXxk2PrwCerDr1Sybt1rTWCvbFceup5Uqp649GAPMDG
aqNEZ6hpUju6YKJ50BrzqfTVYaIY+uQJPdTql7JxCNuKEXWULIuic3tJB+vShqtQ
gZpPhaYz3tuo6P4qJxZcaO70PQvDblgOr7AAZutymkhvXDLVjSlJrevs+zArbb9z
LwBghbzewTRThYEKblaAMGf60GaU0OUz8f+XUbF+spMcam31KQNxaR2TDpCHASQF
Cg0LYs/M66RDG78cRIHdwGm45zCA7dz5DqKJYCsC7OrMQrFZJph7HE1+WGeai46B
3uyPAT9veUIogijn8dpqs6La/8RKaCaIM8u88cZGQSO0W3pZ5yW2QHWNbAiTfO+u
hPxhCCe4OqJ7D8/Jk48RMfs1ZOFdqMB7OQnAD9I02rE7NOvqN3H8DayEMS0F3vNV
agEfyQ4h/HPVcRAPRx11HSDNfWGiVHwrxfPZmOnTMNLrHxZAGdLkXkSE+AQGUMaC
SR8Y/ZvZyh1xh1WUp3g3qxM/tWSZqm7OTwHeMtkhqjdmlCo4DcSll+9f/E6oOMtI
V/zQ8TwRUiLng/6c08ne771PVFbojxIYCC5eBtUdwB+pw1FaNnBcC1XNDWBulIlm
fWMscfIY3nEkb4WMpW/GA0U/DVKPyVMyzWBRsr9jwy4olq/TSbAQWM8QEPVue0Q4
N5qqLIvUcZi+k8ltJLy3ZFQdRGCNQGGKmpair40ZUY5m8Z+8pQsjTYUzPIuRpiLB
TdcbyyBVkyoB3dLNl3Wsw44tIaQjH2zSPDdK5KH7vIyzI7z4kM0f3EazwwK7bWwB
7s8wd+nIto+XuJ78XK9jrnQyj8hrmrkJMAG8ffUr/lxt1LtWrIa7QuJxzWuJFWdT
6AFljuanyW7gM0CrlTQ0xXsTaG7RFQyHJAOBOFIu2Cf495Zaf9sIQo2yeNWv5uBt
xosIK/ENJh3zlNFmwuDnkLDatQ74VQIuqahUR/zGp5tnWdXLHarMQGtAqJzv67Ne
Qqnb5/bMlA9Qhd8F7hnwGFcIaZJ3Esoav4l/wbGaLnwRutPZp/dYSwr/bJ9VuqOP
1l4DD4FHQwVo/tm/clo3q1B+H1a6B8flkjlCgmBt3ilSZPZ+s3WYQbh7kVUYl2YP
wsrdYJnD/txElNU9cq4D1QtzLuLLMVDv+jGz85s+oP23NmtoCLoOYP/UL5pg5KUy
h67v9SluLDg6kWIsst22WSXvFU2VGUwr6qIVRRQ4tBQsaaQhpaf+kCVuvE39KAiS
bZqbiFkZBs/Fjod/497cKfMxFzD+hmuYbw61dXLAcCVHXOLJdF6Bn25zEyBzr9PW
01VCGB/LzEbTh8SNL6/VklCGKJ/oI9nKcUZSrNoWgnmLNdPWKmyFv7Fqez3HlqoO
qzskh/npqc0mgqcign8d36uVSgsBrGgRGurhFDrs9lHutXSqUiC7wfTlZFQ1y/8l
+1YWufOi5YPetYEzIZRXBGfXDvzSKHLpyJe1jiyyOpiqERpZ9DdDiFVW+v2KCc7M
5j7hYNUp9CP40jmhn5ye/ZAS33ES/lLIIfvRLmLaOpnyY6/EL78liKwxh/A0lol9
7tziuj5qE46b8gzozem8qNlNhXdTWjD5QFnCMRVIRjGoKHYpVvIVSxc20ijjuz4K
GEbeLwqrXMyw5fQeZsc+/TSCTbyRmjGlmpWdMgIH4OHrAfOZWTtP4Vh9IYV5lV/j
maf52txxmPAYDvfnWX1LFovkA/lO5i9iyhP2VpUYcK6gaMqiqUzdAoHmYMHip5eL
wMaPvsYdXRSQjcEAc4p3eQCNuuJkW+PQbIy/7BMPQdGmQdJNB6s9LbPbXzhP9ESL
icpyZUbVFUAaInFU5W78VgnHo8sCFF821BwClmZNnvsLRGbYcUrcB2NqyXXLp2u2
HNHO1tK7Tnq9AwymIEbaWXZXKzub9R60dMlBZ2Wf8uUT1a27ujMnxNB5bpIJe508
oIvL+pSA/uOO9zKQg5aTp3ipecO26qU99/yoif/pp9VwU+WkQuYqY7AmnILF4EFd
hPJkVE6Q4Q5KkBIE6Q7Z6TzW/N1jJOIOR8Z6Nf8wAmxxGFN2dhZkMn1FrdfGNy13
7Qs0TtHFCwvdlUuNffSr9nen6ZSBSewDZlnSk1J1vTYPmErBVkgMVT62NJvXvyc7
w/Z9Qfu8SQVNafbhO/Ckk5h5xKsQPf73+HvV2913sLSIK1nqtjfDdzZXv9huiGvN
Y3EQOEjGj0KIgxabfn65lsxMORBbrjiCz7pDE4yPcXOUcfFSxGR/1g0LAmbpvUfi
yuv3D3XMQJHqngWipNCWTXMJeYubiCD6GFv6ruRwfuvJ+N9o+76tK8jkRduuYQH7
Wau+vEgMlgpC180Sed+PyYkg/S61ChtavgY8BmRHxr4eZb5fnbcurbEf43bgGF0Y
Fr0keQijc4pvE4yULKXsN/E/PWAXP+Wy4Jxx9KUvEvI/Ca0tckAA0H0LpaM1W9jL
Rt/Fi+olz6AIy+RUbKJGQTt0G9Gmvyj2r+dVYxTxcLvdhsKwWgOYV+oRmfIl/rHF
7FiYkH9rfqOP+oWCl7koakSCshl6DJD4j173XbMn0KpBKksp+9BMnxiRqmoJxX/u
dUyhz1wu0Q4xX17GQb/NsfBFKHyWmUtQFzP4ZjETts7qozWAJ6f201synIG9SyEa
hkerQHQTQV0DEHeHIrccNvxLkuf3RL8gw+maZJ/CVsF2LfA9JPdncQYkSZmFVuE2
CBZ1sXegV6AIbS4fQr5Mkc0A/4mE4SxaABGPu/d45IL2WjpinR+RBNmO2Qe3ZIHC
vw9uHXIDtxC7IyKtg0277YaLRkhVLPN7msTFOL1I4KqYQ5IAIEjmBmHPIi0R79vh
F3fBGcLi+ybZuUg2YQKbhW2md9/YNl9CBkcigiI3LxCpc5Bx8ELxRD4J4aqNPhVy
8Nm8s693wmg8LegMKFnIE/k0taW2w8BZ24czFKCX9/Sf6xZ8IReeVLavbNavtg8s
IVyAoGh9NU1XzXQ5S23NhnhWQQwBBG/l3HcmEPMYBbkd8EbN9qv+3O/oT6Nz1svS
VCDCpOJVxJayheiXWPY1+PhfXP7gYec4hNvMj+uhZ9TWS2QhF3d8F4Kj7E5MPfd1
vJoojprIESwf+RiRNdWkxrQlnp1JR6v3o0gHE94IWCBnvs9gqnNaR4g+C+HKSYJM
yW+zraQ5sjZDAZcu9NlltJbessMn7SFtE9VIVBAtYR+G5pugEKBABHT3jB1P7BVM
nLkao8S0liC16BBZezkQ7K49ymIBZ0lyOPATLavnEXz2707db/rBEzcG1RWVPKwE
xpysiJJTvPZUHrWywp/zYrGF9ZWNVtwcAI+RnWUeYesgc7wKWdOp6OyzzN8q5V0j
1QnsscNqMmh8tZI1rZU5CYnPZaNf3mWM0mnFYySSnU0WH8J/LvhHXHX8S8qbJHKO
EqpzrvTJFqdo7pvuyskZyn7laENEzRMTU7BEhLiIM1B3zSYPdvNgUrEKve5x+nQT
QNHq5X0iEjCL4CWzJZHWAPo5bZfWQP+SL2CxWVA5PpLfrOUBAc5M5JnxXGdGNWIA
AWvVyCG4bIzHPoxbFDJMrsYfD8jS8sHjLZ6Bg66J2f0BTtNSI3BrmlUttj0RjgoR
Ipllv5JYlmnX2rFeBubj9mRX7pPVLvHvcw8n15yT+rW1UsU6ABaOPAt0DpLqnELH
ThukNhOKSfNkvNOleHQjwxr7EDxzpzqwQ5pwn1oMfBNT6ahI4k9glIBn32wdNOUI
N5RTdeRbQQVWQv2BJrSO8lN1loV4SIQDa9E2fzmfeFndihxJGNRQfqe6UOFeqA9/
Fv8mEbvpNnkY5AuGslL+6j2yICQHmRBsdB2Z2D+Y0SK35FEtn/KpInb2G+IKXYOf
bO0BxFHy4nhLD1QXQO4rpMfZg63wG3JyHqIGgL79OJhRkJxXhMQkHM7AkNiV0ubE
Lqb2C7l06V0MMCXI6nYfuofzOqK0K1NL4eh949sypJGD83vIQo9zK3jfjyUnxWF1
gFG4app9NDpBmjnRn35d6bnSJWULNS8XCsmYvRwMSnwuVpPbQtUs9QOjsn+UoY2n
OJ7xgUcqvYBw3Guh3R6gEl8l8Hc294fdPlCtXfTcxCSdrSMi3bpTQEIJf49OUQuK
//fWP9Ugvx7qgxhtaewLNpDw5v+rqn4J0thuwf6OH9IfbmMTeq3+P3/kViUQ1Xwc
OrX0wMl6apg7H3ax+Ke8dSEwjHEDYiDEsLKTKNc3lFIP14bfntZN/RI7SbtJSA+u
Nnk0c6jeevEylqu1f9jFgzN/1+aiVwVAPn//mRSHfFmFz+kl07Vaon/Lp31CfYoE
OZvvGfrHmTqngrSZbKvoeRuz8kpjbngxdNt9Tj3C4EJQjI+WZ3eUmmfiRqV+ji2X
4KQ7IwQLqsP0MbFtzKFO7lCcUpHrAvrAIWg6a5hRQBDdaUg4TTlH8CqIwsfV+4Jy
NlQPP3UV7q6rj7/izSLo9Gh8ZHbsojANL48f9oamw4Ba5CRinkgHD61ZJIhFqnTv
Z61dYeOf5bK7gmcNNEgnyeE14ISqhQyy0vGiaRumCtEmvP5TZtJG/Rh1bh1zhK02
tOYzEkj+y1ktuz7A9KWhYFZdzc0Xz1oPzOiZynx6EQKukhqkliIgZgGdEJg/NYS/
llIhvFUjgNs8xyVfGChJSKU2F/Ss9uu5vlwtoQXaY4vUu/HkKz1dzO2ObNxVJ5Xl
GZGwtz0eZZNee7AoA1QH8MkWkk/zAaGVTYUK3vSPbVgVX15DrO7lhldVxyzWXeR4
BPEpMJKnx9T8Eu3EthGALHtYzF+hLnyLW5vY/uCq5wtuaTyhanSBqNDkASbEYEVO
O8UJWHvjHGSsyXy4z7AJKbObhORnm9Sj5KkTDdHtrAQJQW4bOHF+ZSzK1iuPfaU1
u1DqcOzJFMX+pps8JsiLpeqXbXlUUywjL9pw0dASmScZSfY6uztsLSw4iCd9Uhus
B2ywIeIlZaM5O0on70lvnlfRVvdXJky5YZkjLwWhaUXvBRuBILqhw5UjRwjyq1Rl
aQiYErpOz8L7Wr0uvf59TWBeplP2eNw0apXE62pkLr/jiwcM0NGLZRVwsYWrJZlb
FrRh7sRejYb40G7xPavA2SqnrO/g2JsKDHchYKYLIGtvmGYRQNsWHG6naQU25LsA
9zel3jzNLhWd6rnjEmnNniPxMWn79tuxkKCxkcpRZ12544HnJ4J6QLjYsyf+oljK
vActCGwQx47qGu6eNNOyo9XACAdawq3DJVHjyvDc4ERM7WD18KiglcSab7Cr/Kx2
oG/rEZdh7pOADAOeBEfp/c+mXT+7tm9bUCl8OBuu5DeUrm5JmT5rhNKHSnrjY8LR
eDg5iihIx9AD+5/2kVWRmDFeFcSxjwia088QwovHuDeQ93CcSrbi9R5OQBoAKBG7
jGqlHkCGaKhBdt/yOewfDpK+HmPgbovLbS0IICep3WQMbPjqp3H7GuFMjUI6UN8C
bASOyqYiBkfyGaZglya8kYK6CWfrtZZR7RPrJ2yGfOGf3WVD9CpR5EB9NSapRY00
lyKcwErnLrXSpp+Gwhab8rK+H7Sk//uMYx3r3WwE4/086SvsvM0TKKfk0nHBExPv
PHCcUUfFOMR7nw84f+cQCqu0vKFfiyrqmwKtn2vF+wQhjStLZryeMDb2Hao7D8+4
6YDDE78dip00dVQ9yfCorjm6PeOX9AOW2v1C5Q/24v+AQu1ZVXeKb23MWoUUSLJb
v4ZWZjE66DRetwoiX4x5QkSnYPtFY6E6+JyGzv4uZXzZaOwMu3O3oj+HdG84sb5i
2BdO9n0cfc8ANB453edVr8PYDFdJkMn7wGLTu7iT/XtJBV+x9KnXjPhildcQ/VID
V5HL47i9GmsMDDhsB2PFn9ySyQi5mfN/jL7Gi1Yzy4TAP8hsSDcRVxGL17MmYEA1
m7p2yqyN39aRXMQextQ5Ifnft1RHkUBpJvfVkFe+flR+37+JDjvPFq5xlRKoSznw
7rorCrN0ISEueUmDiOoJLg0Sga+zJNz2wCjTMqejiANFBvC+3XgEkREyYjglJIW7
Ki3KNnl4ebB7dJTkoZFBR1Hd7YW4CjiKLE5quFqjHpFrF+X2WFISgLsOPpj4RU7h
g7eYshYVstxeKpYy5f4foYQXcxy8d6gV+g9t0XERzeXn7rtuFdz/ujqRysHftcpr
T1tOwr+GHXPAsmVwtMoPillUV9uhT0D7L+sn7lUTqDNeSmbKO0/Pkhuof+RZa/IO
FTIvOy15PfJL1XrUyCEcWoDTvSydAnVpA43vWOOlWcOiLzzmjpNjV1pcNhk0cFIv
42zozUX6LRJJvdNrKokmnwDfmt6KELYsrYjs3nubYMNYGGA3Lxs0nIKc6J7CcDFz
gqGGo6KY4FTT+xQE30BKJvI2oEbP+DyTIsHHPM+m68HqKp7INGXvVdbtLVvqXKUE
GkQej6ExrVcYBhBA81u4OwBWBTx6js5O6R59xHETykWlJ+BqzilSWAtiQtJvo8A8
mx15XdLa+bgGnNIZRM7SEJpoe9y369J5Pr4H52dpGV0Hj4wvEWNeibpDIwWGZG9h
UetFIIXElQbkE+fo3bqRq8i5+adwD0Nbjq3fjUCckWGqHcEoi3SF7YBH6FGoqFRX
uZ3yxruZBjf/n/hdkJrGoJ3sAr2bJQ+yh1I+L5csjKmPHs0GBaE2MvnkgBVDSBa2
vGjfQcG4g24JRfSB6sHR+2T/eyX6an3jvBM1PBEe6dfzSx8ghkSlnt0b0VxUscWc
CBO2gqCs6wc6PwRTL/mqshbJoA3ctZ+22CoTtO+PKFsSGY+G/MNvBV4fZN6NhUb9
EzcLUnee3qqIb8sFybPAEgPjvW5zkhUuakte62ivGbUThU/l+HfXbQeH/Rn4A3eX
/TFpEER1PFr36cy/Vx3rwbY8epBmAgJkSBHsDfXYYAZkUz1BQHdHFVofMVVCF54b
YNpkeUnJG5RDYkE6SIfFtG9ceLwKP3d+VfNxQw+ZwrzgmGJuRrDeQQEh7GEpduln
5Ebk0EfOTTuK/pQmb9EQq/Spz68TccWkTxAi8ZCwrxEZ3E3uU9vQIa1dw4Fg0Wzi
4l2G5JvmBiInTZQtCgQU8orK+gS5MCROgXE1k1mVdsOkIIO47PZYezT3vioop/fy
vQBxlr85RlfLFDI5RxdNB/sUJJc2UvqmZgknKmyLLbDz0WAg25StLJPeYvJu0Fuy
fmnXusXBQRgj8AFOi8gd7TmTji/JlPQEGzc/qijcg0lzXbxEbpWMgbM8xcie89BT
LZUkk7T01vLAUCv53PqhwMvvwe+yXTsesLHwnzLmHJYXJlsvFYjIh0W/2bHMkoEc
2J9BEMJCrJxGwxoPVidoRjTH+GemYmpYs6KNUM8DDv1WF7yQDVa0h75JVWZB8CZi
kT9zELtpLr2BWF1yzZQAiuBD9vYvJSCsasHNB4SLMT/tdt5mQXTAaxerAIrfJtA/
ESEwprev83lt9OayGQYZZHPhHO4n1XHKSSsv3mvha0KpguUBUmZd2oxQWFC6rKgy
+G/s9l3Nu6MrXk8W+bNbOeVPUAFfUBNTONyWPsJWF9itrQVXyBuRJS7+GqB6UC53
HnpzicZQKQdwDkYvNswWrWqPLSMx7zx+9VNt5X8dt88X+P2lCttcCRZO0aOOnhc2
r8WCsuPJFsE+9HZ1YFnBfqixRPvFHBHfz/ujNsQmmHEhSNeQE6jnsFeuQz9xON6O
G4HVBT3M3LOgv4ulhCVlK4MpOORkHIZsxRfWQyyEPQFV3Ma2ld7rY+LNXJ8I/cQq
dS5/hMKCwPu7axRqWEVK4H4cR7ZX35R7RUGN7h5eBwWPzSgXQmn2xb3AvcJBu+2k
/Efl30EHN5iP85gSn6pUiMPCZaqMwTjtuP+wg2HkEV5JqIjlC2jEntTzmPSscm89
SB1CZrj2wbMCJ2u8kJNBY9+aq0TqQ8wUrsANFQTdUpAoEuUmqKihObKFtrbEJlbV
6e9SBxmIEmvohCbQDzioXD8C6QN5xg6ldr9iJ0q4kv+6f5Y++aViyYin6hCc/71T
8DzCXDG5qi/8GguGRAQwlWxQKMQBAnHZ0r+/IWX9a2HmFMhQUMLb6U24hlb7nfOD
CC28s7+RiYHSPYwMV+fo26fo2duvREM52VR7XRNmBj0EvCrKuAoskNSsVdjcM8ih
+DsNcW/m2Ew+gJvTsvqeg57ITIvgAbY3QjUlOaRnDkwH47O2wGNV9cigDTfD5WbF
WZltZY6hdm+piMNGAMQ5zfAlT9biILOTxk7Qqa/HRH8tDhltVAGCsWWTIOGQAOyo
x9OCpsW0s23WIetU+SeXvUcF4iPySQORCxxfY5kf4X2/YxAc9jDkSuqr3PKL5snP
By4HRVDWoFkO8lWxj0KoNzcBINLc//sgha+171PuDFBMdatwaJDi7WxSQ6cy0fPT
3FKHzns5jg9CqvtJUijKg88y9LxZraX/Cgs3XQt4HoxEG74NKXJODesCNsA/m7zp
pA3ZNWSxffCjUZzzgnrI/Ek+hdEuPyOXKCaln9rNMrpt6WO3pU5YGht8J2PeRPHe
oUxLXVI5jvA96Xm4V3FcDduLfmNh39jU7P3W9ADvQDI8NnIOQtqzIVu6Utg2n3Mu
8HAGT740LumKZxTcv71J2Fp2NqI8q1Jmt/tpAHCn/w22FJAuuFv4M3Y5C3U6UbKp
Z7DN9vEaOB/qT8OymIaF2Bvn4AalTBY2luyqYdMold2hj+nYESWeNj1vY/vpADp7
8J1ds8UVjs8vrD3XCo6vMLbvprGaN/OcNu5DaO4FoIV5xmcyd7yUPHIi+5QRoJ0u
uqCHk1GzF15w6yYYF8O2sLeXOu/XprmacWY08Dx5l9xk68Z+Mj5dHVWVTnfvvPEG
68XiwIvaU1fBrPUZ+8jyeLt6T1oI/qioSi1Us3t4rIC0CqbjgYa68EDFonziP+kX
qwUPD/IdljdjjdHiRKHfbbc7o59cAP0CBJ7MUKEHqgdY7rx1SsGvJMQJfb3xRApk
aL66wX1yFuT6PRPyv+y5bysUJZHzlF0tXEWRUlj1+NhUyGpjWXyRVrt055G+BawQ
gvfEKF905NHar6Yp+hky1wIprPqaBgB0Otzt3sMUiBMh+CG2ttmxOCSJtfeQDw6q
eZlLckhaeo2fDAAlfMe3lzxhZCucIG+QYrO/2pRB6JrLdkmP7NbsUVZvbMPR2TDL
pdoaycJbgkewXSYoelacITCnCQPP9qYROutnkQKufMzVtyybT5dp/Ws7MCWkA8HJ
ljGb5eVlKHuhwnuQOlReriFFzxvagchJXgHzxv6qDUBSQ+bmGB/hNQ4UIs8uiYY8
8KMIz8+WSc6WV08iMNxnatwFhiRhqrHho9hCTNQtNJDdPN0QAE2Gr/YimrqfCSUD
SWy3Kp0Iu/65W/I25Jwlshkjo1MUmMbtznVdzphYBrf5NzoShk/B+JvtSdpNHUDX
HUSs3auQfUaMIv9WYLqbxSGVNEZMo/sFDQ3UHHHdk8nSi9QLwdxMuyoOmX1hESL7
rxZSuYaGwcax1vuH0xcy3xPjtMF1AuCJ1nnBqJ0zlLqU6TU12vpViZDZq62AV+ri
BMhdWd4aCqbt2QLdazIEwLe3j3mNwwDumlF172IuC8V5T0oNvY6ATPkSNFKefQOS
jGsbB14iqYPYcikX8sjG6klz9T5aE9xCKeFCvFZRdGgP89iTE/1SIMCRoE/7l1m/
A9XsUNxUArKy+JPS6Il78EHz+4y90WnYoEzz7hHpw5tB6uSVXLo1hbdzcbSCNijB
nOXimO3gGmQtGyJCwp2TiqeNyJmKoRcDQ7EmNluLGLbe0VVhCYUe9A3LouttHHnM
gKM9rLK/XIkb9u90wUcqY6cxSaMVqR5LDWJYCwGMWO4hFUi8AyAeDnUcFgEu07vd
bA/+g9W4PBLHviDdxOV8ho0o1d7xbtTSlM6bgs+ABpN8lu4UqsnGnjTW2auM9QYn
wBJjtFZ513rwAnpiq+w8RPQoeBr7O36GaaSI+EI+5UcdehDAwQ5P+lsEvpBJw3F1
5GnPjiwjbkCSseqT8QPBc2cUpdxYJdqXeNGOQ9LM4MPllg208Y1PjTR9qqrir6ct
nD4Ldyu3GXGWFeruC7Gqaau3eZr6xWLqLmOEYNhlw1m6mnqg6luOHcf1bxZWIBTJ
pOh1aelr8D9K/p29QyCJI9+wqQfySac84f0nr/f8LXUFehVMlZOQ6ee2IRhgplt3
edL4wgHhw/hbuSvEPuyG0pgklVlx1aNGqD/7H6gvWu8nRB4MfPozlz5IX14xQNSb
TO3LO3bgEZXYeEjkdYH4BCoutxiAxAjbWEYZDtTaULC9DrKObL/KkpaKT2a4BpUC
8CxaV2lZCgV40YuxegLeNILTu0dHWrntYg6EVj5+kQyWBh3CW0HxCx/JrowxKYyt
MeTBL3H58tvYfwtW8JUvez7tuOjmWL4RPFrlg8RwBvNz04VNbYSEykJCyV4bxXNV
EMJXSObUcaQ9PWF+TtpGdqEFfUVRKQjdj0IinEIu/K0OnVD792XF1dEwJeTKvQKC
07i3ed5h14Rb/GahQVjMQg2PB1WtueGYfbnNY3HToTmWzjRYSiOSLjIVX26cPZ+Y
PEjsQPK9piC3SFDMdk583DJGDCOdoj19D24fui10gvtwHrV2+RrkrU3luxhsL02l
JweghxXgzS/Nd/tlhYuyqoCYY3ulqYyEZ5GfpYLx36/JkrYl9wbSpIelBtKykTdk
AubHoXT241MwNHj3b4kcjQ1aojZz/pY+f6PjVmoVfH5FCZgaWhIAoQdJzAwSADcJ
oj1qg7Rd74KLjIGJosPBjvdJQh2FZu4IgyOjW4OEOxf2ZPsxEuskGGNCx9Wq7k41
G5nJsUrm5IwRXlL6AfySxTNPNZNlYrZwxlC+YMufwt8BBmiHanj89TXQwGpLOJqd
yU8xhSNUhcGaVpKdGFoGUUiX1piOi4OKv5miKK5Tco6uESYmwQCArynloNMgHpEV
Yl3a9RQufVPG4jLDx1SI7FRfgLV5pIMwbDFIrQBU9D1dDJNskK85juTBAQ17xacD
6+X75tkmq5iecRcLfb6kwkHvE442ge/lbhCGflWNOt2wmg6rGx5rrfLofIA2UfGW
SZJ3aYh+gHbnkqfH3uXhpLMAmI3XIy363nNjwoEBZzzXk0L2tCUrpxp+HoqhGOX4
kdoedutNRQZMY/v1obm9ZhTh+hFP2zUz7PYYRhNpZ/3P9JYYgfyF5Dx8u4Oxl9YH
8NLD1zPHVka2qVYVoCP0aDspU59VcifJxjX1yqICWyN5vofXaCJGgDkxgOoSJHmk
HfbDemB3hOgtUdbONphyQlcQgO8u3H3HOFQqwz0jHPFhyEIqvDOm/mCitS4TAzQA
0ZzHDVO+FF3AgeHNy6DnbUV0Wr8KpCZdOvc4Txut4Hb2HhXyow00hRDi2FQtphxc
D4v7giJ6RZUzYT0xmaJbZABYkYqScbZ6q61BcZ/cgLa3Ym6E7zk9/4Tdtqoj8qlD
cDm+436aNqGJTTX8bVAnn8u7HmJ6xpkKZazFPX6foed2YtJbm6eZ5J+IS+sVAwWQ
tbUDyyhCcrZtG4dknfBQnKk4BpLUxpLeazhYM7uFtsPDnJAb8dFCyyaTwzhVgX8K
fkdHeQiLbGzn0DwnYDRXjlhBWUSL3iITmz7Y9cRJjUwlIewfrNF/UTBpDZ0h6QFX
8wdep/CPf4sYTy4Fu+19GCSuBPJEJ0lwNPU1U33/P2QOaYZKg2BwzN3I8unLlrhB
VMp+I2Jj6TTqGFL+SOq6JSCrQowrdR/fU9Sr3GnLLYt/sZf+QLj/wX5m4F14VCpT
+XFjjKgdsW1nYowBr+acWZkYfVqJHykqhsDQIwce4r8hZp5q0Dt2jeDqwNuO/3CL
PX/hWu30TonFZ0krpoOlsLP3uJTSDhBYqw1UoGWlAWCR0lv7QY6IpA/drL7lSUNA
bxTmzHhd87RgCN0m3T/yEYtgiBYXVlY66DzC/VAB5m/W5f7w3/wodqxoCbVc9Ryk
7ZkAgorcaSL4QyHaigMKVrpgkWf6PvQ58Gbr6fWSiAaZsu+aVJYUbnPWuDxK6hJX
Gxme3Tn9MqODlhTB7q9vjgBhoSVg7knIbgG7vRnNlS/f9MFVg3gD29AzpLd0EQFX
6gWyKn3qMM5RHxhELyd7mWIpNDlIVb6C0/8YgK/m5bVyloJDO4Mus+FFtCkWD0Mj
6yPQQ4FKBwz1xfTBrAlkgGFfPLNs6W2aaQTLo0Fa1r30sdoDOPKM5P4g8n+0B+MY
NW7OsUj8bBYIVv1SGk6/5q54o6VsbhZfI3Pe4J/khjPCwKoCpYeLkGjgmaH+jU3C
KK/jxv2ei6YRVRlK9K+I9oywVsrth1Nj/P0i389n0niZFFWEng3jSjU366Z6vBCT
mVcjAmad1+xhedZh5ZN0BSwqGb8aJTiKYpb2tYPoOj3Agbio96ro1D5NqcJ0ipBL
7HnP6+QcDTJfPuOGxaw0qjhbclwEfSDZunlquMepE+zn8t1zNQRruPtevzYDFrmo
Fhg3cr6mN+RzH1IHf1jYpafa4oTuaQQp5YbA4oZTtNbjnzAJkBfu1mwNv2xMPXYs
BJ4H9VH0xiuIpuca1iASNhn/hx0CrvI6Kt4VIouwEGXJum8uvVEEEnN3jVbKI/tC
gP1ZfyRFjK535w0liBqWA8bp7YBf1/wiFKv2JfIksCWw3qzO0/6MVlxw9ZOYhqup
ksAqzSqVdD7x/gsZUNkgMIHZlJk6dPT3TH+tQY3C1ahcc9XbRhVxdvaRGpoj0bP+
4K6lGEI3qIN/83k8tM3oUJsVGK8mOBa1DYl8S8mIN1k0mlkUMYfXuWZvexcyEFPU
avBoFvQjFts2kwC1E2VDH4wmTcqwD7uC8hPUiE4BYLcBDlnanLTtUP/8NI6oXC7D
VHbFgVt8VPXeeqr6r/ZBdYJebBkl+Z5qAYQE3wbcn3lY/xIWszY7oQvm4x7tHegO
8zQTp3Zk8wb+0lUVyXRvmQ/qturxWab06X606opRAZ+2AQ3+uW/mCRTZ/HszhKiR
MKP5Xgz/FPwtA4OedHWU8ge6yy5ExvqBTXhD+BHwhOQ2HXKhKHZZm3E5SKGaQakz
elNA4PNg0Mk4sRwAho9sYCcqMPuYt/CLoO2D+EsVpqhXM4EL9wZQWCYbCd5wlAw4
EVcdKmp+AecJD99QrcgesSt7Dcdpkjac9RcHSev0hTOiK+6qsJ/FO4Fr8OOqmZ85
bpnnkjEu6RUyFFgvMXJIVcJ8dPGh18EAbxwTBx6l431NT7wHPihagCyRC7ANYqXM
yUFImxT6hesMgrnL1pCdDUDHfq64VlF53vHPI61x7H7XtF4OzPz8SdaiLAyPgs17
LNEB4Tq0iAsQEx2sHMpa8+SYH5PbnCYv6Vm8qJHG97Xyceohoy4MeGvjL7Rd3G/S
fgnuc0h4nkR55aazcfsOoTTTvFj3d4BG5rW2UhI0PJiAaRCOZeFunOqCM3a9RK5O
mGl9jCvJgkwhMtBInqtJ91sd7hRtQJSELAcGuC7KNjMmn2NNWxkg6394T0nMRhnq
YS5UoCwtQE6A0MibatSRpdmxhKN+fkMlRNUAxXe1xMxmqJRLXOZwLRhgqxVjIP26
MMH7S8ato6wlXPX7E2poLeo6k2A0XCjF25+4DLv/RG5ydvEVwMVLsRal2W2nUgjT
54LT/E0S8LoNABREJaN4s7IJqg0yKbRdSqqksMUXiBmWjq28v2SYOLOxvayvWj6+
7vxuPXlZ1fM6huvXFZPyl0Psz+EuqzxnfmIgh/DGnojD9tNcZBVWYI/ZkUP9AjFs
LlgQeJHP9Z0Dw8xRXj2s3POVRh/BBROs50N+DhX8P5qCs19YEERpkEagGWJ/2xbe
YcG3c0KHxQGxneV035t9skG+CMSIVJ6L9R2RPIKvEyqEEPZW1yF5UR7tbkH2UdQk
LIgRPw17ooLWp5o7a8tS5afJohUY0GZNW+o91Rp/8LbYvrMFDMpcsetblt83DO7b
n6m4/h3m3k8kELfTSJZ6LH1daTh/S7J9u87GtHtx7kdKOhjyayE+YTYPOR9m9ChA
YgYAX5B47KkFwbhymBMXuN5wRXRJo59Ekc0ROzNBHJhJ7wTMhQvKkrE30JtM6caC
SVzn3hJuLWe5rNQnJNJgMKIn0WmA0L2WcgsIb5dO2NyvSwwU7DEVKze71eAjeabM
j7r1C8BPof+PTmWNcMVznyhtIrkDLWmS6LdxuJAdMo44ULAZp/1dK5+TzwRyuNTD
Du4yzlX7iAZVi20PsiR9cQEbiHrX7BMetWCygr9YTx7HhlE2Sh3NZPAXZRpbYI4N
Ql8IxiXlvxkrqhANgP6fabCzl3w2PcmM2oERgjGm6H1ZOs1VCYmIWTZwDA/U/eb1
UvO92ikRYK95P2FhDvyYeNuRy3EaT5KcvrH5X1HrX/MySpAXOS1mq+pdmI4g3HVY
jw4DG1o1bmdJ7mzR1wlD2m6CIfto8akad7FMTH6M+zU3Rp6TAaWkjVJD0GHNvZXp
SbAELQsf7fjVptcnjqnGCa8+nZoVsZRiWkP9Zosbm+v53xWX1Rnwi9QnQpik6SRH
MjTxFHvLMIFbUJy9zaWAfBNIahWmvVriMcPdz0Zy9bWlUeM2cfzNbXHy4zcSRkPn
FhAu/gcSmqnCIxvQlB5tBJ3PQOkJ2xsxrcOakyaaWhmuMfl49YkeNaqRWESZO9gU
hbv9EOIdaF1iIqGUVqf6TFa9jyUMqyFH3GUBItmKTB9RZRcZ4ggSdyH0WXSOd6Ho
yd2wWYmvRxucoxMF1uD9CBIBK3Ch8MRzVy0aGC80ZWqN4/eHtFF3ZzLZ1CSRrSaY
dquhtjc2YzxttlHXD9oZKRSdb33duYQfvBV584MAeTklnwGMYu5yCQw8D7dqOMOc
sSqYNPQKOKvsCvhAjkSlgNVlQZB/+O1WJL/lFLCRg4s4EwRj/V67HV6LGB412Uqd
kz3hBdeMd0mqHZaDHWnV3mOiDUvn7goHCg7EwGPJEftX+xTdAwCLVsoEC9E0fU1m
WOCr5PmEYl/i8kCNxIqLSlvibpOP8pHXQl/sZ4E5BeoPnRRxLH0LhY5kdHimVo9q
kZQ7GjBmvyIBZ7MkOSvHvczw0/XkTjtc6407yvHCZHdym03N7s4K5ktfaj2C1Bz+
QTL0HAB2Rzp116alZ0ylmOnn/nQTStVjmsMckjMkNgJKasLmjwphhZEGFU//6LdL
IDFeoI89SQlIZqTGDdxYkB39h25ZwcNx85pzHhKcTGBjBW/QLaq6Q1klyzSrIvyd
gu/jxNmOggfEmYoevhC7nSwAQ77msZdFjGkt3xuHHAsRU4tummcwEa3KVR7RuJ/w
x5qUFHg48KxlApWguA6RKYz5ffzAZaHCiO7YGTtI42rUq6+RACRX3Qh24CSWBnh+
Itok1awaSlLNHfGfmX8PX1GacnhfuUpkA6IKLEFNZ8+npxhomhWpcsJRJuN4oArw
4vAaq/7F67NNf00ZN44TzhZ0WwblazWEcoJwMmEK82hjfmTZMLM+cXN7vDyydnz/
ZkBW0lYRivp0/0AHm176L9SstHS94cE5CPYJ3FTpIH8GF/SPc1duU8c5X6bsxlIt
Q+R2ppRBOdHdGmkXutKr0cl2fDtaZMipZQn9Hq0RbRGt2WIm8g3cvKCCa+TzL8RT
9GcOUxwQnQHhbRdA2MdLbBBCT8BVNnApXZnTF/55GXCWU2gBkwZzr6A8hkNrRZQR
5Geb2p5bsWk5r6ivSl2P2opaumWaWXC6YNFReQqOh15GwHn+crwOLwpcpW7qBPhZ
Rd2LA8DA/gMcn/DkdjJSMucZxTCoTvDVxe9UiUJWw+iqRb33NXtf+ClkKWiXwcfG
M9AvQKyfeM9j09JV/7xWEfSVoRfPH8P8tzdyeEyEV5CF2x7XrgmXlGCMFQmJ+PM9
mmhmD9hEpq7HqAdKJsEZf5ab9jPu4V7MjtwClm082v4qkQgxl8zY0//kRMpmtp8X
j4IgIiDlRYxsoX/szjkvbMffvPxNtw/BOdJvq1JqKWwiKYFMq2Pv00IM0GfvwJY9
TyFqpqWd9H1jiGLf88RmIaRCTuPm6bGD7jpYb83rM5rWnXnOIJWWHmT1EBOi33vi
aeXGvPG7VIZg7gBJyzgGQzzAXV+8ZwkYl21SnJW/7LLcU19TEbiAxEfdrAlUEMW/
5b8QANx2a6sAgFoiTIVxh66BmtoCRXeFDaLdxhYYsUrBm4+OvQ/7oUAXuUQJT/Ev
2DtHNijfrKkI1fI6LKCnPgAiOyCh50L0hu6IR30zOQNS8ElhnBKQa8eXh6p9Pvzi
9HRAa1Jq/OE4C/8EZ+FuzdM3ChctAM69KhdcrKObNpSA7GYPuVM8q7tNlOEhDZhm
WEqmjP2I8Qa6mydtjv/2mgvSCWVL6+/WjWqx2VsJARqd66n91jxlen2Vn5Xl/C5G
+mNWPNpi1pyg2FkQxmWuLHDxwnVsSWwEWcXFR6l4myBtBK3JTU4tFYNGndWxGJCG
sMBIQRMrMosLr6NMijD7pTQ0buJHT3Pt5TxbFdNMNcayltlyYYK6vYSmmWFZbf/0
vU1ZNezu8M4fztyunpEovQz/8j3mVieSqI7WzcURS6C0SyDwWGwRphN9FyP0u37e
T6Fb/0EYEfhTolrQfqVS9es4rIHDkzyZar49moDN97d3elA05EyKkaPrT8SslzFx
Irk2ofaGVY5v7E6KoRVNC68mhz1bu5+9VbNHoEP6F74uHObtV5wFZkqRV3xsdp9m
rJw6Z/8O4Naiyf6pqke5CJMskmpdxHWezrETBB+LQAtEvjY26GNy5KcNHDVlLuA4
4imtb4DGYBkHKHvj4PjOrzbpXIJXQORrMU/mSeoWPJBIHrYKwiC0gV1PxHxtj2Gz
p6NvwyNNO8x4tvFUbfhF+mD3uK7Mw73tKfKZ0n7zaAN/bD1GcmO7tl3Eys98GA0s
vNUo4y6UfoA8Lj7KJb3I1eLQd33SZ96i6JF/XYkEBC8qZUP6tBu7z1Rx682tuP4d
yckZ/ZsnlUIw7QgRLcW/mRPO6UXIxIWhEIG8EWudnoAktosa7aSZITdGoqZ5mU80
YKbodkPd96435LGW+TNHgPF9Eo1R6ijnAdXJ2E2flsNhaFPzi9yhrkUmbxo0Xaee
T1ycXCr+/90lRhmK1gsElbL+hzUJ2Id1Kdr0BJ0Sb79cx6oET5zZPsxSFcIYWYyW
lKTEhcO3oqvdfedM9DEVcS2myF6DGv4ZWT6Mg+5VaaENTesnDow9plPOoCtLEpdh
1/bLWJ4R2TkFNkhMWMUOLfqyEHRG2dRJM+RfKPp28JPZSUwFQP2FpDubAj2M9cwA
as+ZFpUpsBGUq9kErvDhrZY2sYbrvcWbiR7JBaD8YtloFzyOfMumFRbIVLFUNJaZ
X/qqfrkcQvo+YpzfqqK2VT23re60+KV75oTkMeA24pm5hwi+0v1LUw2ehjrpMZWg
c2LDeKy9f1Stn+B/rE3XOneI2EaSXDDlxMGow0peyLdlD+UN/emIYDTjaWNFB7AL
TazFKQdEcJ7pobSj7TnZvMZU5XNomBrltyN76gfDRnnI/wZXHvN6xC+ywpXzN5ab
Di9muszHY8IOtR3bWceFY7wpGPCzw0geuaoulMxoPpPS494TyrpHsGemvhhSkglh
NCgBJd/UMLMRRW8dOmDuftlFjUOGEb1bTsXogKX4uyq3SrIA+qT+6qELkOE1cUqF
7hoQ+yZ68yl4swfRw1cdjvCJCPKhrQRn3Q4RyU36za4UK+8rPGXim3Xzf0LuGsbg
n3K0JXYCN62ubgpWA+s+NufvaI0Zee5CXK2UEiqBp6aCA9wue+VMgufJWsoGUTTV
h46oZyu4gX2J/qyxsgC+AhU+6GEngT3cIcArJD5Gd0U/OU9DNPEa2+2a9lmm6LGl
mgL29rjEkCCJXuVrL+DycpoYrJ5AeLQbcG8BUCuqEv8AtWUl+xhWmTUg3m5gdm/M
VdavM8OobdVJO8IuVkPyyFpjnk+UYSLa/4rKAVlN+vMqwCxfakz5qhrZydY/7Yno
bMuwQI6yZ8KqIdBAO8mAsl14ipjYddREkv16NUBtJrZgf+EMg9Sjxb5EacWgOO9e
/gu5l4GenQ/7Pa4GFn8RC/6oSD10p9uw50gSMCXQJvMr1WSMlDfcIl2tSbjzcqzV
OWQAyk4On5qQzuuD/6KjUxBnIzXoLSPe/eFCwl1CKtsr1swrOzo9W7sApZZsIlt8
RuZdNy5GtIcyuYQyf6UEdXcA0yw6/Tv46+SArT+fRVFJPNwXWuzX3Ny/IaDUt1Ke
D5hSmA63tnxSva7YhSQKpT5eSkuReIGGj80XmkqKn8B0IHo1hcz6iZ2rgdcULJGK
QYl+qmrdbSTSduO9akTZtgoWDhJXQRGxo4d8Z6il+RcSm0+Z1E8Pc/WlhXpWDm7l
v7V4mw3DUclroAi0TNkYhVSh0uIXc/X4SpHi6wbGyRhgBNcoMZdqvc5oGSZ7ENRT
561s5XcmLGdYfC7Wkx5OPKFlUh2Nf+Pmpb+fALsRqdeJ3oLl55kdhcfk4KMHGfMp
So9ePHSjhImTDyChxsK9XHKHgXv4YtkMp6e2FE4wCcl2+cSmUEhpuBGq4ij1xyfP
kkCMo6vcW1lmH5k0d8dQkL8CpKyjni1eQAs11nlEZkhfYR8N7ez60rrsHd0uHWYa
oGIiNlA8v42D4Ma3bQpyA/uqOH/0T84fQ5T+SmXKLzm8rMd+VV3uuW3Zuz6oe5Hs
IwIkxVvSvzLEjXkVUk4/6CVRIG+Bw2qRnb49yY/lFMw6RPvJTMgBkjgG/34PbwK6
eHulyzZvlBfbZHyCr+FtWcaWszx1bq4VHr6UfggVUo1tlkEMvfRLUgCdBhIoMNCp
T/SYdcBgoR+XJYJAMhkZvtEsJgH1uIwG5aINb1vn/hlsqnBHuACI34g0kr/vboxE
oKKCuXU+RZ/jsjEL9Q+GaaREC5Yy8rk2cGvCkcs7qMXRKoOch94Nhdr58cKGdD53
szM6kxSoo8Ng23fd3DZdJsdOnxnJL22bamxHw7RgEVCFaTVg1m8wAdlpI2CFWo5e
XE/OsJXIVlr9ondazhLs3itdt14PDBz/TT6GxN9WYxi5mJGSNETYbQTe29dxQs3E
ZwcAWjjT1bnQ5dCeXn6JJ4D9QCZdGM90X4KgwXGpyR+kzqiXp9JfLYos2nYZaZbF
D92o/hlAXmWrlM7gBo2Vm/7PJ16GOuyUZ4/ynnI1cBmZbhgC37Xrfwmv39KKgo/0
vw4zoZ9Y96xfogI6S3K4moW4BKegM/KXSHPnlNIAUeFP+9fKS0mVVKzTG5ryf1tW
8x9b5qtqRzyYBcypwywNC63uWRyBXxERYDNppNE5U+ohBn9Vttuw0aHKErIEDC/l
I5qXHIvoKY9wnV9RQaG0vVZwJaGWG9JjWuIsesechTeFO6VAdqUpb2LoBiNhV/IQ
87tX3zxVFnVJk4x09mKP3Dv2MRtOENJR+VQGg61brMEdSHUye/g8wrqpr1QwVCZK
qpnQ2SNHyURo6FuyF0uEp8XRrFvqr7qrOueQDnHuTgG9o3dvy+a+MWCAFrbmlE8c
Oiomb0KGFXWbHeu0TA8dn88/Bv3FZjvgm9edVV9sfGcLPzfVzwRYxKpBRp8daUKx
W7Ofw8td4fX0Hp4mEdqGqa91QZwme0o/DSWOZEoXasHKEv4ebQ1ScMuHaXpnqVDa
9smZxthLRxOmWPruaj69GJlWrE5xMND260t7OEtIixuVHIo7cIvHbcLKwQIN5b77
5+vCGqr09L7pVT+qOFBLlYVrjuIFEZbWSdL62rXJQQjEEhqiggzU/L0ZJV6JkzA7
t0piH2slurXMgj5ZIcgLqj4fwBAtH4PJEFgPG3AgiDwmM+Z435eqcoD/Qgms5aAo
Y817qg1Msl2CnapGukxCfqHsiuTln9CJBMkDttEUlPG8Rin/He+ZkbZARJ0Eqmiv
/3np3K+G3zmUdlGLsEdN+FaKNf0TwYxYcMFWF4jVU7+8zd/QXgd9vTQ5ACFw4797
dYG4hjoXpcpT2z4lQ/KgS/TnqjyW7bMWM3XmYESx1EzBJ/fbJF/8hWgnLLvpIMgj
PKWakgX/MGBgQ7MU++PG4ED+G7wW0LRqYJ8jSfWO3f4mt9Z+ajot/MbCBU0kqqcb
Ie9wNQ/MfR8mIKy8/2EevG01EakSDi57JLbatNB12Sf6KIUJwa8vn2sseO76oOHk
7+4H9djB9VAHtCIejx+OPuIBiZ9OMONDHSdc9lWrfGqawqXApnryWxMjcGzV8NFR
tRaODQ4siUeoHlVCZ2kkWRvBJLBP79Ce9vXhG87UX7A4gzrH3bBUVUvToPvP0GPu
esuO1OyJysPKkHvm9McmibJ342umi7NF1vPKDczDsjeDKYDQrxWW2Vy2JMqLrI9H
MfSvambWKT28moqz39YIzehHlkT7twqFSplZ0Q6vz+DrGY9NUrMofO+url/4n2Eo
moTt7LB9IP3HC/xpAoCgowHLanFiK6R+kjnXRAnOZUzOrHRFOaHv8TTygszmOj2c
DTJTZKnW3fPzI9xME5PsLM4fEYa4+JRENjMXBeKNxQKIxoewAPYXFcBcpGE8wP4B
wW/AgEJzwvYLMf+FcvZBZDXeo7VhuAnWzukSpeuLuPEiKOzq27rOJBcdo02beZTM
YUtKBphDJtXqNLaxWxVnkFQCoiawzB4mDVgg2KjLt5HuIP3S+5+hPPsM2GFItL5z
iyZfTIQklRJx93KQMLHMTW0TxnEFg/oB+UYWa7etMnao2PQe3WifrD/64piHygQO
EW1CQ+01AX6xRpuGa71fasY9Mpmi/q0ej3+IsC0+DQ9lU3bOafz9D4OGCgzasAh3
oNnEbuN9sneMmMOFrtHCE0fQ7ucHWnjD8Al/0lRaI368vEP8iw29iBiNAF/RzAXB
kTX9UkBLOn/OVZG3qHlAE9uASyqV4b4hVr7tqdxP79QeQueH0JZsvfw8JZaNdaEs
IgyvmC+qN+d3S1PGwzaQ+e+1Hf2ri4pdUeSToeY+gaC6851aLAANQ5bj2+dlfSr9
PwNHJBJrmSKTWNc8rvVWt7EwqtXj95sG24y7xPfKVUb76ka2LgLH6G5WMBuQuHNz
JW7uQ20+YoOI1C7I9iv3OCKihqdskl8sZuoZRVdPS4bZjSTH4SKGHpaBsfy9DEde
bJmwj7Lh1M4vQrW2CF0VxPMaA2A2Q96l18XryUoOs5aqGidP1m9fAszSD9ZyfZVa
S5dR9KZhkvi4wcxL7l0i7IsCuOr23UYB05iLaGBO0Y5jIaYP/y6RTrEjR8Cauw0g
D+ORoPqL4Xaw5MBzxIEEErZ/lhqp6uM+fq6mJMIYMzK9gQTxqZdHVH1pRFOwTZUj
rNwNJm//1maRZS3wiXGpEuSJYYYdYnbNC8jez9jRfAeZ1IfD3z8O24JIW06NOCaF
dtpckOKZoAY1uYjiZ7oVSXMM1fB+JJyNbSDLnWjPfC9DV7tzvNjMzXRTnviucXoh
fy9uiiIvqNgF+NLEq1kH+BMEAVpknMS2f5n8IuLVYyZaCCU+XOcZV7B03g8AMRds
kpg8jjQplghX7tBWwgGfCykIStLZ7DyztMxMQEiXyDScwREU9JYQ5VQxOHheoteN
zbhTwQSlmh8g01uLLGOXJWWLzTNLwU5S7tOqSzPBbrfYtpLsUFtdTdYSadzB/6ve
078uEt2w2JjSL3OthOND0JhNaxOeF1Ge+vMEv8dUpnMyJJ8Sbwt1j48l7mLjoWiV
wJ7atOYxKLa/dfYc1gbladUlSMlKZylSfAyTmndNwhxoy/hi+DaDBwdimHWwFzgR
o453ceyCvHZKhWvP2SjhOZhAyD/X5dSYHdw9ydhMcyO3aeLtu1nBbaIwhTZc3CW4
IpRKnWqFPpwSrCR7yRCZ14n6ldOE8sYQ+qTA0d60etpIBB5RFKvROt3RlfT+A79u
MMN7fCN9trBsb/V0H/i0g4rO8csV5zdCsekgWSt1jgriC+BuKt1LT9KVcBwK15GZ
mdsSYkEHrwy3BLYUiKxtpwNpEL4EOudoNxss02b+zWnz9+XH5H5kr3/DvEhEZmpx
j3UdMGoxIZWF3sjlmgFyNSnTGKfhjkh822RTTP2dOVrSP+BrbppvuBiZZ0XJIB5S
d/xcd85dv1jWncDVzLy1aXemqd5PapmAWe442aOYdmGsqrv4URYy+IXf2V+f2NRf
rleM8nc9+cHH5ILE/R2xJ3OZ2Bap+bjryNHGCFh1yXtUnbAbdm81WJoyIpCgsEB4
7ohZ4IYPC8n20d/X2MlV1VCcMtc6y+kTMPvRdyMFreynf58FXMDvlHMy90cA/sfI
TIxAP1OICnGhUBu25ROIOUasmDp+yPdt8bO9WcUjNdSaYKpw7wpaAEw78zXXA+xT
9tou+Ewsf+o+FDkWDmjKK7UK7cI1Np/pYffZs6YAFEFU0M6gGwruEakjHf0VjsDH
a2Eh0JO+hhFDP45VJc78in/fyfdckNxXBYxt+MI/k8FDkl6gb7fGtyXx+WLXWWzs
cno7FVQ0aSnjivxd2luGPWmcoCO9UozPbiw4BZucjrO/+p/PbvuV295h5lh+xd+y
1CoeARiZMkxXNJ+TAerKltgwPDrOYBlE6ts0qqBfO35ngcl2pDRgchRf/n7xdH7m
0KO4zja5Rmb97xGdIebIhIUjkPFzmeOOEKWEzKF07JjU9LQZSU+47PPxeUBMn2/U
me9LZkX8uD//1muAwFH2zGwEd8dGDWQAVvw73ZpNBWGDACWDvkfTOtGmGJbUGwaD
oufPdCKfTcBh5wD+MPA2UZvXLQ8vUSJpn5f20zclbsjYF0CXno6OnUDaGydIFSM7
osrMXyrpvgWBHAFIE/DTiT1g7EXmW3tHCSGdMmZ5/ru2iufRlLFX0HhJibt43IKx
XhwdgMdVE4t1E+IiAcEu/bWQ4BGGuAHCW4v2uAhixebaf9xtwVd2Cf4g9r7/p+Pr
Rk4QP8puzcYBTWSvcTuj9fOsQq4fEJ+AkICUrrumVsRUCtkhiPpXNI1txZnF6a+X
kji+mhpUc/XCH54bfa8EI/0gXOMW9a6w+qKhHtiaB4OOWsOpi5aHYQC2DXWdv0Ri
Gw9D3ysVmKqKsCWDajRSUwTTPjXlYZ16vIU1GyQTjrD8sLDZEPDSigU1lyz4pqIp
2zND4ZD1A9juCZf79b+pViOqtp8o+9VEdGAPzyKOt10fazJ8L8jVFEAQUKDwcjBx
ipYA3UNgKb73+AvLNG2fgxOARX+nyrXY2xbpSOhzlqDWpvE/TcS2vDFNiXa0vSwF
gul42k8DOWHBAwTgkFrB4VNA6nrH//ezgi6kGVWze+I/FK5Rbf/dYPBX5hoc5KNA
1upKzS9hMAgByglTTqInbCLSgUppR9iWyRrrFfwVHHse1DJAb48Kr4bcY9IcoLVD
M0eNZjbvVCXGQLxarm+kY9Z4LJi06aWIqH+6EB4Szw5Ow2WVGHqM/iI165gSsIuu
3WzRQuF7SrRAoFIUbuMr1lN9jOZ1OSJNYzTb6RS/i0sUJiIXVysK/ej8CPR8tN2w
6Mib/CqDXaRI+gpKzABbnsZUk9UwZ5OINqTu11QbJGIqPqY1T4Sv9mjYHgOG48JA
5YhgiPo0t6exG6wFAIRiWHg35HhVPr9OcrqxOrm5/fAafpBAbdphDK0iGVBL3OwU
MM5D2hs1OzKcuZPWVntG7Ck6Ol7g+Z83Gi0TUkL1l8W8SgihVwxz+I1pDj27T1qW
S4VR4FbG1CKL6su/M3mzhGPuWAgpVaRB/8H/H2CoXk6GR17p5/aw9F2u8pLxL1Db
9B3PdCgH/NOFesQaX/qh1hVfJCNHQbXVIWFjtU9yqOf62NZmOOPO2409SKW/Duy4
1bzVDgOKL/J2mG4sU7/CAP/RvYviZS71qv6Iueg6nGPTI80VMdWCiiO9SLU0hrvQ
1UC66F/Rfwotqa64AQNcLPh0RQmupytJFkOjGiyZQI8I4DMQOF+zxPdc5Ni8k/tY
ndi4j2sE7gnyHCiEGO+/TOq5nmrQbnH6/VpyhwXjm41IrBhzTVjqlBWnHnVOWpuq
B20ZtvlHUTa7SGTNal7q3DaP30wbfRQOk27nKUXT4Fjh8e8AWvyQ1C64KW17zqd7
c+BFsduvqH/clqjf8ujg4LEovMDoZvtANJ1ZeINn5OMZ8FKq9nHl4D5cu/uGO4a8
R/Lm3ryNCSCu6z4x3n3ALAcTaJ/3ltr5TtOYJnUsodsBoQ6k8i2zENuTU3OCJk+D
PF0U0QhVTw5a3uc3M3d1gp6DryG2dZyDk37ipsj423tiu2ruG/Pj3uFYs1gFV1fL
2y3GAR80qWp7La7RfCByEzzN5/MVLCjpHnW4ACF3C/cjqPAuQQhSAfcHvdvydLW3
Qv3jJmUWYKIWm38Ks8BMi1Qr+SQfi3Rxiun1nIyuDeW0EIBgjdAF0qxic61ZLmv7
5wLPkj1jOfMxe9588kycQeLIMCD7lU6gxwylxN7ENBhUX6GFGcCzLKEPRX/IL9Ab
CmU9OYBu5QjcZy+Zm88VIXZZP4jNPlzMzVLKH5YNAZtwRiKGFumIfDmsbwdUrQDQ
wR0YYNMBix1HStX6t1UMW30GpLX4PvvWcywZAke4Dlsy9Te66appcSXedM5gqU5t
FZY2Xpl27AjJR7fgJSZ+3DFbICghQyRMFGeWHMzZnYO7rmjvdxDLMgDK7h1SAEeb
kBdwboDBOl9lmHum4HYeeILl/OYWkthw//vYSu416ewW/9ODuJkGhymRCisk1wTS
lyk8rdUza/i0itK5Gj/on4jORxr0d+bFBGMLKNdBu/vdZsoVYfu05PzWBKKz/FMM
/oBtCM2ezf1I1CdiWFZ9aDeWb5d7eSAhdDsWfuBXrgWH/qJXpxI/wTGdu7X1QOxt
oc5VC4RKVgxCPRmzGTC8rHQflZRxRdZGXzfHl/CPCEhPH4oCvj32y03r4yI6lVUR
/hipGzY2Gc63xZoYsJvucz6+B3wcD+fzyZADFD3ghd73+Mxn487CTeAmbyfliPO8
LDDhwjO1pTTZh1LjFn7QEkEoBvfBjuDF58axFs2QUPHOUVUnT79aDsncrkxi3SvX
sUS+holdBemjzwZAETT4lNLwp5BTEtlF1oZog3BImb/Q6j1TFSGXqNHSvMN5HqwR
in2c1JieVTp5eymtjVICuxzL1GjjoKjqZpy9bmEyo4Y2vyy1LvBXq1Wbx4R/J0sH
cjTbT+P9sh9qhwoIvk7AoE2MnwN863BSUkh2otcgddFLIqKl6Gm3BE4ef6tVx4TX
qivocFO1S6Ex4hOrPiA9eXpc8cN34uy8Fb5WgclJuecraO1hUeMX1o27sZgl9WyU
VLVKisSiyyqC/CIaFFxlXeX9c9WBKJMQP74odvYkWJsFYM5Bd1WlQrERKZ2xZl2t
VKuz65qEebwPnMsR4Lpkkq/0UHLMMnDiGmEBZM+bNSgtXB683H5SZMjIw1vbBheO
ZLhxrxDDBdgRzp8cnetuQ4B0OohipW8u3ynTvXnxozVcHsQo6aKeKT4EzU/ezstU
6EkbYP5KoENKPl3xSk+nbWIizp0tCT/3Y9+aYwvQTLj/LzIJRejjy/+nnbtYdOQf
J7oOivkjmOC4Tko/yb0x9QvGHjtVPOg0Gu6dxkuRBerHLkDEeAvAqvnFqZk9MOSK
vZ//UoqSncQsUnI1icSwlxFonACjwM/zTYJ1wngD8LjwB7MgjAjpagzjsqDOGtGE
a4knPrnWAwKRKGafzjTcJ8nC7H7m0PT/nFBn1OJGV3/BMrzuKXgvt+boyNF1peVV
8+vBCCur4PUxNy9quChLAbbagnRDHnfIXaJ21ZDKDhW3yOXj0U59rP61b1qFn2ks
Hkzl12WHEXDYbmGIVIjzNeb1AMB0L+YIfO0LFWAm6APED69NITsr3hbKUcqGOuFs
mmm0vFBSx9m8G3N6z+NLfBKHKWcc1mIoLBgWCti129rA19hKGrm3oS8En9oAS4jJ
LxtgOVFDCvHORVFxbeMe6am0hNV4/i5DC+Q3vuSoBvy55IQ6bNIoRBdTupVX+RIK
boa9kKSedM6t4QhVltAkFw+gXLtNWwQeaknjnYzvX097WysaXPAzu1yST66M1aom
k6lDtsuARyz0mJH6ybG5zqXa15YsokZNtnkEPVrfqSfEDKgzZE3XuM5h3poP0hne
tyh7kGzCr5ppoxAKWF9NaM0SqV3aM29xr5VT23JhomgIUM9rzGppFDaQxfNVKJny
G6LG9Tp1BBXsbsLMSJsK5FOWx4CUGycfTVsyJX8GWfI4JB4J1EUQ3iDunw6Rdt0m
HZLBnWuAcqvHrRm2sCv0tnerMpV1k6c7J+xGAqPDzmcgqW94dCpDVOKEz1yWAYGL
PVhvg4MO7+rF2mPGlHo+orxaM/aA7NUa/6nLva3+4Q9Aspgw3WRBnslPywpNJo2/
sGzZ62Hd9hCHVCNMnRjmAz2Ilv2J38IAdxYkN0R5ejItHgRKDK1nXeQzOZfWgLUQ
mlbEia1b5g+KhplfIuPUut79mNeeZjC+io5/mQyWcOvjf9Rewocwstm02daXpJGi
kSsKBwZUdxi+Z8ZNbhxwrViDmfq/ke+vVvLTcXp8kmGcTxbT2Fg+j7z1JqikSfKw
5tN/XUu6KRUeAF5rhfUrj3F7NlPryi4rj1EaV5TGLBNh3ey6Z8s1bcGxl/lIZtgM
6xYjQl3MUuvdCDzValOOfwM52RhwaVXXq7eVYo08D3SJaj+V4lkKC0+/atiEMC+Z
7XB7K86UnGdFQbWM2dUm8VWajzq7BXQfUNauVOLJN6xFahgrdGuGXLrszFW63UB5
xHoLsuyRwDc8IJv502i18ZjXxFw/oEVEzq7HZadGEmSIu8geoqNiO3yliFDMJjDM
hcizQCFHDoYIqEzO6N96EIw+H9Ha2pHDzwwYKs6awtWJ/wvSa7JtsmADV0a9TW0E
i4ONnP656G0Wk1Q2vi5/eQs9tX91mhlnHSmtvN07CL+k48fuzFjhV613+bQF41Nd
SLWnwPjpgXERQDJPpLPJq+lxzlzBZy3/CocmhJrwIUKy5z6RyRP/mD6KhPP6okPT
xO8Nea7i7inShCDgF9bOFGUH5tKHKoo8/2O/Q+J96y47yYcndFZW4+kPZzfgjJpo
71H6H1a5xcNjeVp0jZhIlsS/cLsTOX412dDQs/7TxCH1K430AcK3qTbHOslL9TxG
C0xASZxsB9UomJcSSVnwXefKk21CXWAJf+9dl52FObSFcaX3/vzj1B3wWbdZ2qNL
khOu0wQFXKJ/hNKtBosRB4BRxVLyxoSze59Ar2BK13IgR5FWdBC4pT+6PPBlMhrO
rpSJ9KEFiRarNUXOsLalJ/tdwfzW0wzFHkdkp4OXqSiGWMFxWz8TcCbW+89yme/4
tnkP9xNQc/A0a7b+JB1/CykpTBoxa6QrPHzf3KUdpEKv2JIOhEbJl8aoxCTp9W9l
qKKArMR/0bemmqtXjMnwuT9eClnNRxsZU0u73VXIy5CGgnMhNa67a/pIahP9Kwwp
zaZhWfY9Ho+TlYjN8vowY1LHmBGSpFU6fEheJFT6ktL/sAU2dCvOap6zC71eWo5l
mfCwNsnuKJRPQAOCXaLVo43tCOpruvign1XUANdHBQ7jPnMVAan9Sq6l98MhFsN5
k6/SzSG59eUfONxJ8pNsWhLWyRsDGr8ZTdC2X1E+pM6T36wPmM1pHRL39ap420Cb
Vg5u2R4N/JIIDL/U4kOEdyEsCF1fILzLGTd2vSyA63u/WYy1M9wygAZ+C9iJzKNQ
d/xSRAXRTSlICQQ3mlhyUUg8DIsTyfkRN27ulabmdRWM44wIdNOS2ZItWjRqd5qc
9PIElf+3+WCNSJ94TvvpFNvsz+AkBr6klRwmNqgSA15VD+boWgfp5XN2cZkNnpjf
HcIOQF1lplotoIyM3VkvJfbNB3CHvhRnUg7gJTST2HjQSPHuAbytKYs6gD6nHN9Y
1QerfDB78yCkgovPDdPtAkr/Dwptu6PKrrwuq0l1ZYN1CniRgazSyW5tQjAQRNaD
66q2jAO5LtJ33KAhtsFY6RTZjjgP3r2phOoPKmQDelg04gd1w6lSRp/KEMAnf4jf
p8iLMS3KOmxY4X8aRuwxTPPhdy/XtmEgfRQO8K2BIT6StNJOsO1IaeOmUqXM9/OJ
twSK3IpMs0SqCl8hLOK1fi5m3fmjNJBnZpj5sHJI9FTIZK/LlIQZwyP3C8IHnoGb
73iLCet+b64rcEr/L/yySzBAt2nNRcmcYwKLK9FSvEy0uusFonqDE1mIC7GqqvHy
W3BhrXrPV6q3XFFwket4iCzNbz/o3lsCq20cuO9LyOc48n/reDmXHwrr1nSjkY3h
5nPO5/UNVzbUiwF97g/O/ryKd5HQy0hUNRRgfT6bXCFqqvL+ityVzMITQkfZ9Lr9
nFhm0cunf7+ILoGHmLfRJnkfJ3Wjo4ISmDyvXWiHRTaqV4PJyr4YyfDrCkp4xd64
rjPitpMuUxM2UaYwtsi8QMwVIy6sZiRRrS7zxOLY+LyWLZCWF3dnZ0sh0IS9jXzc
iVVXkKrsYZoAh2wjW1zwVriAsgBsjWBePnzDGiA9jOlQePcQLI8NAu3jC1L4H1Ac
+cSkLe3JzLS/0YhPUtECeWYPJZYUiJNMu/FhaA0CWSenHtnnH6Y6FVgmKoBnP3Fv
QyhtOFjYgQPV4Mh0PjDGcD6NmvugjaDQvG2rH+UBXhJ6uuEmtCZ3wiICUV1Mvr01
H1IxQLlFr7zxsJ7dvZhRB7/CPh8EmtQMAB9yRz2QTbL+h6DkU6QJBDhY+2+0VFef
AeKnUVi2pi7czbcpwiTBso1j4biQV8XSSgrO1H7hYB1oYXrHrWUHW/ngu/p8aHfs
MnzotPp7y/K1VLIjlI01MWQ1l5yJ05B+WzOu5HfHFT5vM3O8l/IQtg/qsA7VY1rM
Fhy667jwM3KEzoeFzX+N9Sn8waCIXLytojUae/r1svovQBgtmrSbNDMdkiT417X2
kx9eL7czCsQrI+r9op+ac2ub69AQvnG8yWbCdD2Mg3QwOlBhplRoLnyWkuZ/y/vh
S2Q+z1eHhelL2Bh7EbqrniEqKYXkiVQFm4XZ2NYijEG17BXVT7QPN0K4DZWeW6hV
MUMr0SIpDEhWtoOXWuU2CANcZKjzmdpncchq/tBV23gsDZ6Ykx9/Rve45RlSJlAo
kGsRuyY8BgasSDnPKenvdc4XlNOVVfvLtdvox7y1JlzPqa1IXEyruuHS1biHH81I
KBZzABJFVBwWucsPJ05c1lBgnkpYeyr1Eh2TtReYK3Yu3pylkD1JSUOIckU3pOA6
9LDipelQKj2CdxFajGYLYc92FJFOfXBWJMLBr+xpwsZ9iGkadcQC0nDqmD1RU5RO
xyam8cSmo/0evehelYcn7lqtJBVtRnjHisBUE69zL5TCyAdwj+5ib+e3Go80qkVn
ldil1cGKI39jpXYLKEj/plP+YpUhlSiSUuX9KwTCapC8OGaBc39ADVVvLIstvd38
5oS0gLsLNFlVSNfWGeCKuQCw7QVM1YTIYtQmp4siH/PlpfdN7Ke+kG8uncwqn/0e
E24h7qUXF2xdQYblORFiaC+sHHxlVO/BdkNfB/qXChDdPplEh9EIaxR9iMrzrssK
hoI9I4GRKcFAVeH92h6cAwPFjgone6Rzvpx48RTip/DPwhjtqOO1fYL8Xc669fTx
kZM1ye4Cf6UCkfPS63FbcPnVh7NvIz4WkqfuhFySPlofe8PQtNNY3viCGR1Cx9fK
WsHyWAyqJLGbukxntThOldfTHPJdJc75sDt4+afyx1NViUrPlbA87qOQrrd5EJ3e
CbwJYp74rD97ht/sH+GUX7teOxoAbw2D0zX2/BTw1gVHBfuH3MZ0mwbG/kEd6CI5
Ow/w3m9gwZ4VzpeH/5b8qPR5GMzszlsB3pvtadSXs5Chr/aTWd013GsmL8pDeikb
JqWXIfE2R5Z1ufaOPHwxsRqBFRQ+z6OMfS8rhBoM+KskFqfvrpcPT+/1k7gODIZ6
/MSeLNPzzI0tFIRhZg9uzg4ICD5XVNen2jV40ZS4V5qwq7DFUdIYgHoi5TWmv8Zq
0pkd41mPoiXaqHpUPZkWCTvlbMOzmul3SXAzDYXqDVb7HEIgG1GiwmpZdUOKaYaN
Mex+AdPoU0RjxK5ED6X3NPF7sqhE3p25pb57/NBpaEcttGbweiJ6ap0xIG6uucNv
/N3Ek7jOtWabw3jRCs5rAA==
`pragma protect end_protected
