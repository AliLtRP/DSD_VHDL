// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:35:33 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
lgKHWE5+7+PRZ3slZUTjgb8kLr6Ujj4eBWZSE3ukv2U5wNlyX9HMDc678nKQSCCc
7tqrRDcbsGUvoOGJyNqZEmrQ+RfMgYM6YzJo19vKzoR+1DevH0kCHYNYfuAeCypQ
tjzFYSaXrsO9Fhjs23mcQ6tJcXoSxOz4lsP6pN6fmlQ=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5792)
CcpNPGufAgkcEPgZcqDUgXn4Z1/h6ejGI1o4n9VAyBk22HYy5NV66ae9hDPWDYT7
aibPQPv75OMvEAU4QJ3EQAtfT3ycL/g1hp3fMqv8tTBdpwJVglasuMjmqdL1EP19
9Y6Y3Tvyu5sv4AYshUNSrwfO9o6kFjqVl+S3puhd4lUmK1yGUcmJsUZYGbR93Bo0
Jnx7bJeqn9qIfn+fCZjG+dTOGSs2WGTu9srBOainTZLPOpBUcwiIRAgEcGyxxCwB
YuFOA1zLebnDcKgGB7c5RjfY43IDC5OpXLiY2U39B/WmsYJ+EPAspzt3G+w+s/jm
lxVTOxz2F16wCPuGruRfi0UhRKQLK6YyxZU1RSV96IH6NKbVRo3KNZFfMt/9ByUV
OP0GK4kN++ABjMUfcITuBnH60Q3jjbGOxBDj4zPCPcuu3B7lKEcYuezOonHKw7zn
DX9ib7UWVtNmdBS5nDoneTCDRdOBUU1nUg0PPOKA3vVoyBo6AUOOsc/4URkYLYeA
zSr/+1zS8/WfAvsbzT+nhIrEPYEzw1e7FAvzJOord9y0rkUyYVnuz7bJAXYcw10I
cKRqa+r4h1h3Egr5d0BhsLwGtdWLYDwcfBdQmLKdcS7pf1ZKBzH8H9bBOWFECfXr
cZF6+7slW2kgK+u5g6v16/Z66CqJ7YmghpuR0LL+AmpT2/H/Ke57+IRRr3qsTYBi
WoqwcivXBYHptbkOO6P5YszdUpWbenfxSlrpPiPuxCvG2cJNz3dQO792Ldhd54Jf
ubZFd55q5JU9d7WmlhaImgBAHh2AgG5EJbkez68nMZcLnaDCctUx1cHft6KBlx8H
QoYzJGnSCAp2Z0xIVHGOyjIhQ/AAFSKs47x0d9v7w4+ZaE838kh12zEINmc7Ejyu
JsTRttpGlWHZCbMznV0d2HnUJsi+G9IxZJiIrY5WJgkvtCI3UGStP4KrHNR+eQnn
cFtRR9dNd/B5hwdSyE0CNiZefRHHwD3vMeOM7N8nAqPnlk+ZD5hhLxaC+PfScX8H
QRaeN+9wTGo19ybD3TC+Fw1O2IA87vUlHnCwPZut9niF7SKiqD/nBzMC79r4fk1Z
N9CevfjX0aeIfIVMLaVc1hKzLE7Vk1omU6Kpc9BV3B3m70skdQeSl1s4DPXr1yC4
KDNy/2d5juvc//FMKqgQsRjhlegXv/kiF+ICFl3h48fBP/6edkmhTns3G5JeiMNK
bVHdzRl6QWLwyIJuB5ag/viki+U+iqHzvXQZXRa8GHptfJ+Sd/rPUQ4GNyURABaQ
w8zHFUD1NlKMDzg0+GytycmRvPzoQGhk37ELKHW0XAt3EIXnF9gKK60NFy7nnIJ8
JKLgZzsTYfTOvvxgxyUmxKuYzydHj81sgWjnyTrYlLIDAjbZWIhTMfsczYPq8vql
GYxrYNimUFfJJo8PzUkUXmdyOBMVDJW/hH1hDfiMhzZn9tHcKxg0n/whOHkliRL6
lf/z8ulWImWYMn8+ufVh9GfA78JKoADAVdLmfG3RgXXhPyq9EDPjagPWgXJL9DHm
UvJ+3x6+VuU+ta9jXJ9NntaHFGPae2y82ou+hohhni3BSz6XNAcm/bDqLLMD+7k3
/n3o5ywJsWaYBNRFFGT8aGQ+LpA8RfNrTYRSP0Svv3RdjVO/IrWh6Eadk+AIq7Jo
Io1ayiYDj88+OzXpRDW0/gwWJ28HHy7FpXaBGIBgzk7a1EtyOqOESENdM4SC1UJS
Zwj6FcfJfHdfwBuxbPNQdZaIWhNdjOuZg3gy31Mu1wuvT6gZX7PXhAeF5VveM+Oz
VAENWCrEYSvatOZwlCSAf6uPp7J0jjbgsFHtuxzRroYsDq0Lp1c0XXuJfcZbETnk
cozDg9Z4rP6WJacVix19gZGw5+tPU8i2igA1A0S6bQ0gRHgiN3atrzPeoDOIJwLZ
Zhs0AMdFWwa1SvnIQZU7/fxeHe81iKYT5SC+qGuZhbloN902MyAVZcPapPhxGSbh
r0SWIfQtglHxaTwLAVVIwBYf9IhtfTU+4GeeoGxXGjC8lxN6HufPJrJw3Acl9FP4
cIOJ/+W4+w2o7uRxY/IRA2yz9Ra6Uw7pKJZQfp3vJYfQGKg2E/n+Zun5cnQ7fzbS
GwOIbzXbFZRQdPrBjxC4uLECH8zoXcEZu4N1Il2ZgnA5q+9a2V4TjUzovvrFVs02
40a+Op+nfqQOv+vU1MAdUh+XKgfqIsxljxqIZDWxDGBeM0KBO87DkUHtZ+F+rM8f
YNsZPUAwMWy8tqJCSfzZD3d5nsyzcUX7ymO1gqEHR70PTnAOczs6rwKA6hCvsEWe
hyYJoXdFxHCFhihSq6MJdorAsIthhC0Nc9pICWMy1kd6JmCkbtMSQQHs4XlRb/bX
CVPdjWvuTgAsCXfkLiSkP9nYrGpzXDfSrReN7l4OmlutAjxn5nmnEbRDvXWzOx1i
lpc+yiXUC62QdwgWkPn3CR+7xuBzvK9BsBr5LtCnp1ijBfbuOpy13x2q9grGK8qt
Mro9mpIWXH/7EbobG3a09g/ZCx/Hpb5xverjejx+xaLQXPzKHQ30f+Q8JJIN96Ho
GImcC6yLnsitjEiAretsQENumQQeEWgcqtFYSnobjAIVHc5dKkbarjZyWk1DcGlt
lvQlrK8CwfnOjjIk+Z3gI1HGFzDaHOO4tWHXg19xnBX6ntcxD6fN1DvE45ReEyZD
ZfjGswf7tnespogsZAgjcYyKp953YCt/U0tFp8XUpqQX0XSkwaxl41o2tHOCIsNX
Z8QNwffWqgfGURgyuYJu9TZchlR8zQDtPaPdLOPbIG3zUq8lPLo+sn2PCy+TI34+
9mZq/xT6IYD6ZmmCOnqAAG1UfaMqKJ4w7i5kZeWonmNUoxcU70/bK4dPYQpLG8w2
DqZsOPLQOToY73GchZOo4tdHGQjLRpGKtIi9l4b3aDuiJyOC4wuJXNAVqj2clkWT
znqOSXlulijAelFVHNgDhKeXoaLBs2GClUNlCZZ80N1aWrN1LmHnd0zEDXZE0+aG
lkX6XhoFaIXe2LBePX0MGCnZrXkqq1+TRvb9PLOorYsDZtC8bHj+o4ffL7ENoyqM
xDPUy6LC/VmELs8MibSXEBDg0U43F1mWEHahI3UWEzX6xc+sOa59K0/ndks09e7o
tPL895JcdAgy/tS2TQG20Kw2elSBv5GRhbe3Y0Bt2DmTratpewp7dkqdY1EAi7rb
QhEc47qwKQ/XtBRVwefoAclsHXZ9ZhFZtZt7k6pwyAjWNWfwkfLXhqp3KaBpmP98
8Xng9r5wD/IRLY+qPAqkelFc7iHs0dgskD6CyJNSwjsJLCzsojkRmh0BWTTl3Yg3
cVE7epY2c22PTvrh6LaRYkIziqsM/jklANbTYklWzvEw8U36T96myxjo1pNDFPdm
P717sp+1Yn++lOAm0nqx7xG4rxkCQSy2yFsX0ksJ/JKullwYpW9XHGNk6b2UCJYC
gsFxi+ifNXq/fhhwcdTD/mqnRhzHvOeCgP7NMP6QTl+FhbaDWrBZnpjFkZzwMpTx
aReMX4xaa1WdMmTNr/VAsGjpyWxxNQkYzeys0ZpHhqunnYxurr+4ckPaTM9s+YMZ
rO26Lhepvu5Qd5HoJobauSz1NSWZVC08/I8Ui87Q3W20nR44Yohl2OR6czroOhNc
eKtii5rY0xSHcF+gRCK4SHzgh4XXj5gPGkGiatw8ehYU5FJIZYgmA7sIEsJN5iOZ
KZs85tyK8Ni0kgQeDeO5Ie2xdeAfp4raCGQIXb8ZPmvggFZlLD56/KpVOR+SueND
MuslM10oO4nDgCm2dwFmNazraMCwZkLt2VBwGGpQX/kxTV0m0q8Uo6dfSiNz9/aO
7n0Mz8H0KlelSVgv/Tr0HD97ynthoV2F9gw8CerEGnf29TQbCRyoppygYqfn0SY5
Kpl8pmyspkL/NucJGeHSoCNRa2geY9Eyk0V/yQZrM5D306yUbLtUGb1NA4gQpfTC
DEZLKNFottZ/AmfBWc6eqYC12QynbDcWP7fGhgOjkrf79pvjtySs5iAITT49uDNT
0ktIv2QWJP2g7ghtQOrElhB6sW4Ds5DxZHSTPJkPNCyoVI6+y+2+vyQ3ETPSCh0x
SvB7G5r0duDJWHpatkBnBlYuzrnve8w3+iugUk3k+eM1awD7MTMFcnaUn2VRhOSK
TMyfCsWlsT07xzF4Mx6phCPFPEku/1Ar6T7JH36fGyidT2MQGv2OCmfjkjB5YCeL
8XXJPVEZ22HQvd9aUu3vogfcLI9a5btj7qw2eKle3hYUMLLNNGsRcnwIlZ3P9XVy
0mwk8dcGjlcksGrIe/ARK/aJ2T6hZuBWsrp3OnqLcnoIhBveoCwxcAAKRgQ2hboJ
GS4BA8dKDrMvB95QCNgmyvfyK5v1bubShddoMyh+B4GiP3Rp4a2mNfXYimw8rUms
zbrrpkIb/XGZko03Wr+aHVd+1Xu6zzqdDt5hUBzi5Xp5FuXOGyq6RV6Amo+W82fz
4pspYLa3I7GpPOBhml1+NGzFs4ADNsYnlVwYQS9RU8GROZK7+rO6pIcCVo5ivMO6
qA+0DTuViseefrir0ojFfNRiIaeJ9q+iBlSEely3VTmbkv8T2prY6asC7RoHiAK/
+7O+VlwKK3lvrTk2RDWavIQ2tKsePQZZaFzGjv/4HQRcKAL1a2BtLhvloHKb5Z50
scM28sspkU5jT1zpLRLfnbjpdJXRO9ER9A3PPZjOmtMPqZTJ+ZNE8kIFs9SjPAO5
e/X4jvIxYwlfzukKFUpue8mthu5ZBHHUcL8waLs9BEQCLqYExBKe8eQ0Pf+vEOOB
UncNH1aoBpWAjaKjZ+1sqbEedJsY4H9tQSzTLsMLq0lpsf84B+k48lE7l3GgpGx2
wAnZ1mNzWtYd2ZChor8M95PcqsryDHdfCTk0OE/iQF2W5/kk8Q8MYtcMNVJxLB2Q
LJZ4rfv7JihcuBxuzJV2RpBiaIoUSlEsXzURzZkO4MMY8J/1hCfqvdTnkCfinGFJ
Wr/LNRR4BZfTD0OtSJBDXxtJ20u+MyVs4awXbmfRqApOYd4JO4YktDUBhNxkcf9O
7thkGlyYjXavfLLeZ6fdIHDkRy8otWgJCOP60mpU94LZMNB4XhrMQe7vejq5LRFB
p+wKR2WTAHHeI4mFS6ARiJSpe1/2nROJ6zDevSmFY1bm65izb6PI+Jin2q4noI0M
TMzVVMA8fk9ObXENJE2DaL416Rv1/onDlPEZ0rRk9pksDOiOI/O2cyTXRZenmkdU
qJs3V/i6zugyAKs/Ppc1X4P52v0hTjDz5tcpHJHo3MrDnxklf+Js/V0CBxLlNTpq
THbal5T23T15gezF1S+f8r/sbpQzg2EyIATfc6zN+dTKlWDWhoU3PEYxinbfUqvN
RJWrE6vzXJ18suxs9XzTNefZ422byZaa6SvknyOtsITnOl+AV7Oa51D1Ruab6J9w
32oJwSe8tQ69ksqkpCr9M390Qu6emMRhrxdZVUg2kFfyLKKCHC2Dqx408aa9IQ0m
btFDrWS1T36/5D7uc81gXvJoA3ZryaSmi+Pc2XR9W0a60sXizFmph9FgwXKS31u3
zdPTChmueAknnSmCUzFDVxw0N21bel+E50X/9nTmtEm0qne+fSBW3ygF7ZmbQ1zW
gJL4cYdN1kmulqSZd898dHtXBBHJ5Fjo+1eeVQ4zR3rxR+qZFhpdK5RcOSBuQjfV
7dDO9UEcMCSHbW/trVDz5cecXySP3l6hve8IF4KVdmoH0Kw+klEOvjcAW2RCQytF
4BUzQ5Jy9J+ENFNYBAMEllO/2oPkdM7Or3KGCC25bGDGR4pUE/cfIq12ZOzspFvV
ldbPf8BKnaAq3Ki2ZfY0+tVS3x3kclEppv4hxA8VhG1kSvrNm1sVJ8n4R4PBIhNj
pI9miaoMPvbDsHFMp1zVeYr9aFazVhehTOl8oVgAvOyTSEfMYm0LTP2sSqnVYptq
rh0odgZvHj3YdhqQGgwxQbHsyiPAe4s2Bqm4O7RBC8p0//fbv9Tn+OCGhk2nlI5T
fYnwXT6oIVqWW0fmie2ZJjqFRoIgaQTouedonaE5vPMqCoFICQkEs9JdZRzkT7gp
z19XB62jF6L95GfhJiSRalCfptovqRJAtZD3o/BXysijyY1o+3ZBwap6RD8LeeNC
NMAfEbEPBJ8OZc1jt0GNre/Wp2CXGvM2a9tPveLkwDPUO3ON2JUQgw5Pbzh7COHl
+pIAsD7PWK9Y8DoRBXUztZOWgyNueO84GV6VxTwA+OFmLaXbbGXvfu01seaAs3wg
w1cPMAI7WhS67RuR20ke/Zo3wZtu66GRfdBYgKVdrMIL57zrKAgMBT1lzgnXy8Vn
uyyiuPJqCQbGzGTd8/h3c82wd+8kd8EuvT5Lj6XL3N21LtG2/TOWB/3h7W7DfW0c
tgkn2bnljPELIiifMdRfgErHrhp9VegNEPgXeAZrudSOwD09OjyT9iFjd8IPYMF4
6eyrB2YxyozEbowYPi0EZSgWqtQrcm1Hph6eISEotQKWxdH211UxCjAxAlsBdSCA
GRenVApkuaoTqPRoeWKNlEexJzeFU4oAr9zdLu72qFbuZq5mMCVnALIirxTzuoyc
f7+FXJ3B9pY/yS77ndd9Z0IUMBzFnHTexVa/6T9DIx30ha/UfA6BZ8UEY7lWr5n8
8+p2SIopGZIWlRnbUbZDlWgVOVPGTBtVPHxR7Ri+2BSOLV84j4nWPC38mwuTtIju
T0p6L/xhQMez50ulI0514MJkecI0mli+uS0fikJ+zv06Ie2KpqE0QG0DrD08tbic
MuAn1+yhpKTLtFwe+aXHGuvvFbi00oSEs9gcvPQ1YIVtzxQ6gsOv5Ez2WvlE4C+d
wpgdB3zXxkVgI7NvujNDGGy9R6jZWQOXRGuyThY7ePbb7r+XcJNfRhiXEmaoE0G6
YrxIrQDPCeqnPrkV45KyWvfcYOwFxKfm41sOUTCq2O2JDz1mF+U6HFBrXlfCcXaH
DQTkQnH/Iwh4lrvJrD4GxIKIGrFlpWZ//n1UBxOixTwwZmj9au3yPXAvfvjFPa4w
+twBOifh517A2m49r38OD8ZA8hf8l9+bn8l7Fo41OEOGOYRdAGmTqmPYg9YmK+eY
tblpLRuD3WeX5N7iSIUQKhIGgHNRByGSHYh/BiJSGwnkf1q9bFqFVXJkGHV6dugt
A8d/zLnCOiiCMiZ5ELEY0t8BdWmc9KuIG5XRzbZoDk+IH1lAH8phwGfWGi3m0bkw
uHqEY6SirQaTT2nU3cd1bnaCOxufzDJeJo14bjAHHXz5rO+9UI2OrXuergS35Z+2
hLe2ZHYFJweC/rbqjGsMN+bwOfC9jHYa4A4oQkVWehVnRWHgslRIwcUtdmmrqUyo
d2mWVKTelL0VixGSgnVPrb5QmSkHGsT7X5ZLvOizmz0jylcOe5iYSWWyemCz1doS
C3unrcI2epWcOiwqiKkAX/9EakdWJUAabQwCPd/J3AspE2QC1Wsb/AuxpZwaX7IY
lczmufSUYFB/3UW9HXU5Hq/1Op9JW4ucAvTR2nyhYGWZwlfIPa1HcU6EfngiJOEg
OnJKkTNramyRyiGvOKQ84YBAvhV7ZYSSdezhX2kL6LRUfNvVsUogZdb4wfRK4Qay
attwo4WAJ+ysfmwmWhj7ZU159P7kLwGcaH6m4KzIULGhurcHZu1o8OF2+Y5Hk4l4
ItGh77cuYzm6W8pprorezNomZ6CB+npUH+nYvLLXl+s=
`pragma protect end_protected
