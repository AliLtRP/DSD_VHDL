// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
V7XKkHjb0MrjBflucapo+iqcXupqvXcFSJsx78f6vE3OoCO1V062HR4r2qLz7hoziGmDkf+xW2DV
IUU/upBowoWsWQFBlo9pRCCFUyVwTOfAAsi7KWacAAfphFq30q/AxBk0U4/SJyyER47x6v1ooSvN
th644QRNg+KZKz3gIelArCC3Tf8kCtrshnaND8uq62OX6zNkBbpgA9yHwS2g1EtyZCbqVvKolTyW
J5YUDt3vY1czqq68EXNOgckA2RZCwWwt10YdxdLfVHw9tg/p8OD3ae38uLRgDD0nNwUr6bHiM0yl
3oD2afTY85P5A8Nj6Z7Sf6p1cMDZIHlLEFz2bQ==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
LFAx7MuPLzj41CEE22RYSIDPGLuMACtj8oAjvBBIymTQwrOaOOLHRuQKp4DiZ9vddf2RkJaZrits
bI7Y+Uq3QYU3kZsM5q7aOJI12YoyrmW9onLimjh+pKQLgFspZhB/GYbWqcf/p348a5twl2N3nSAL
SQZzw0JVhYH3hAWZ3fGrSaduK14gannth1QEEz/c31dSXcW/zquH6bjfU6vX7NzCA1ciDX0MgoM2
uUirb688GGQsQykD3MwzLJnWFf7zd335Ty6ZoY3DajmiR8VC2oP+c/8x+Eh9S1SlZvCEKsiv08En
FB5HLeASXUQLpZNEClFSe9J8OIRCT9U4ZuQwvtGTzn9N4SBckFypDVWCSnY1SOeK0ORJvl2c4Uwn
JLfoT52x4WDLO7+zEri+PhJRU4vsv6H/TqDdHbtXjmFvFU/XDzz9CHtTpmvfCaOYtECHF/EOePpx
LgjgSireTSrQa/IVKwJaSzNHzY8KDz4IbbULU/UOc6WUQ4HacU+lLm2UmuN4jRU8YrvM/1EZ+jdb
QQAjNEXGf6z25aBJFUawDv4thb2tS7YPF20u0a7JYnHn4rD/Tysidzclzm3ikEJrKUkQ4vxGJV23
VXJNBrSyS5Zh1aTrjvdKWBcdTQokuo+d57TJUqp8MFrBLy+NvEs/DFWqa98a70ipGYOPLW19UW5n
HPIaFAxS5B9krh1sL2qzHHFNLty4RcndY7NAO4wQPb7wnz6a5Qdr+FxZ8g+ILUTOTfiMPqZ8YVKr
cOBnl3un+tlkWVy3+d3b5NOKWI6id4tJiCntDVMgKA0pFHeBjIoqD5NDxI06XjD48hrOp85ihfLm
EGqf+4GhqWdavr3poiP/sHxD6p7FUyIm6Ht1CnJoGfUWkStREi15KU/ZdDCi7txm36hQAF5/fu8e
rjq7Q27Jenv1u9BowTjEo0tmasfqetALMase082mSIQQCtlLSmxfq2uPUdWFKeXcznGGj3It5aed
03Vzpafst1fESjMIYewfXLCjQ8iy0VpuGglxjZyZagyiLyICKUy+AMRggYj1oEq5lln97GycskKp
hoGEPuTQ0oM5lR+BnyJ8Ioo3x878JtA/NQLttZoj6PDsQ3gcTQUWPLFlo1bpYkraIGumXn5EDlG6
kRUUUGit75uTPB6PxRFX+tEHFNj8Bep2Q//bgYK1DvhXZQA6qfSyva8I6WMsd7PR4DBZmTLWWzv2
3fRB5ZwrUbZ4Fxl2tBqbDe3tFw2LB7zrBGprRaWc5eXlQJv2Fs86XhLuobp11Ivi7CN66Ml2wSAZ
llepmNaD6l6yuXTzc1ByJHYXdkfWyQz7bPcy6HqD9smO9oJlfi/voI4cqHkUECss9KXaenFFPyYt
bwVdgzelrK6g+7acqU6SCOjHBNoeJlLaB25oTXcvd/XqNtr7R3qAwa/X/mHbsgfODDzWAfzFm9pN
bu3xEIiuN8exgzUrcYbfdRSjiJBsqJsreyOVETlwZGe53tp2CGkIxxmhL4De2yVq3te1BWkputq+
h6zxwj32djfV5K+YmYuZGc0ZMIbV+M0E9OsGPSLVbJ+fCqyTzFZrof5XdFB0CzpF0PvkbagzgYJH
bTPSHT8K65fIsNmIK4sfgkryj/i9Ax+id/ssz4nn4YQ3u+H2dm/MrfBc00ywfZI7/tTXUlKCUJEK
m3/XaihLCKP8EcCyS17toUGJegFDpFBNki3J4mi5Fuf4OScgLP7L4Hjo0WQZZRDrHzBkgBv49T5s
VHm3vmU82TbT0+ooNyvZn6yWuKfwC3WbJyU+LhmFtJPfCSPgawNkPrKZvXMdVvnYife2XeoTnKQO
Hmpt4QUEk7DK8eBQSYBdd8NqrRShgC87WgoBInKifyYrxDlQcI3/NCRu/du5OSBmEkrwkfKcs1m7
HglAQGJu8ib+ypJUqCx5bOFptOWZ/kb5RKM7OCxIVNNK65R3sM5T001y6+PzbE5X0KWbt/3jRnrC
iQjGJECFwDolpQsJuPRDAKYpe00qXAq1KT4vYE8u/R6YE/kJqUt4OkYboUVrB+q+hUgR7I8cR+VJ
Zzv7rm1lpeyS+fwuIaGK80lwV44nj+eZnAyH+StzX9mGc50MfXx0ysWJ493/v2fRt7DKSsduUEKj
sTCqTyW3NP7sVIREwRTHjRRhji0gSu3gjksqlsNFfN1KfMGVcyjPGxalhy6fDzWhAXFwfRmC/yYN
Z9aFGj9xHgUYplN7bVWeGdBXqOagtkdaxm+NDeTZ5Lxgwa1DXEEnaviKqeoNHwd5Uby/7VUcAsKJ
nkXhFrqHsowqxa/m0tPKsHzpbBA7VQDAjD+OXSP/Z/ewpU7kCP11A9ckZSpYWKQhlB4xproPpGEH
MkgZrKGI4+RJWL9XWt4SXxFsnP4H6c1ke1Y8PAT4YGQZHtve8XGGlK9nvYofv9GjXIgLVIrjRn6F
6ZeeAtkosutWtSgjxyYFlT1nM4iRuXwwsU5LTqx5c09zW4+XgR1vQ6FIheFToEgX4LjR3ax/6KCL
6xSPEpfx1G4M6WjiRDbS16N2+PjS2VD61x0dg4JTl9TFaNYOIsYui4y0/Xn+0FKv2lRMkGPqFm8s
6OlmDrGcx0LBYiJGkJ1Z4pp4Yq81ZSAdkto2jN/5RnA+F0FpLMSbCCqe+ycOi0C8/hZSf3kMGwJ5
5ThofOAflbJVfJGn4sMZvLGO41Cxsv+jeFcMuWFEYCZADjNGu07mx9sxgzCBv7cHdidGAxRNNNlk
jDQ130uHxjSlKGg9DwElsHY+wIxEdCY2Rbf9YedthRwe0O8bxR0gF9bQOS+rGDATY3tRwsfKbnuP
zwwhvfH7/LgZSqu50icOl0syPR9+vviYWgmvdko3l71Rn2VkSgfQhdl211bNYT0hJaZtf+0KGjBc
BiO8qG8RdvNXyRHbxi3De14ANMGeQwBZKC135MKP6loRiZygBi842P8L7WIC+Z2sLxwekx/3WVWq
0HQRGGMkziB82KxynqkJ3qEQez0FGravHDNlFmjuless0Re8fEvpljb6zOuu3N5CiD+xrbkv3V+K
oe3KFw0NOpMyp3EXnaMgwPZ+qRPB+EsGogXpaLRVbZk640SSNPfocLz/7Kdv0XcT4CtoO7Z6yScv
TcX5spLcmv97rrZm1thbBWOcPSTLzw8zwjkxY8byN9z2MVhjm75UrFq6yK/8y0XNnlt8/eq90e0b
6vGplIivXPWjr6MRWkPcVQ/tVaDSJuiejKCd6qTg4VSlFRqFPEfy9TgLBHeLX/q4mPKP8X4QtfGE
NFYnsIIAm/YGQHG15Y0An+LVmHrjVMfKBOskFTJPRgh25iwckHZ/7uHuufXOjeOzFgxcyC/BVQj3
EsDOnnlU2Vk21T0xnLbLa9EdNch4RkHNfLOTMzBxxI8rY7OCur6hdUfA+R9D4xoKAaJ4DGjOTmTZ
kKQlR49F1vqsuEz0xaXbXcSJBfWFjTYhjNpwvVoZH1b97Oy7WNhFTil2vbWe8icM0FHtkamUaG5q
UJWbNFdKHFw8E6VcxRuEylZpafyitNtsaTlE4pEEe2B+t5wm008x1J2X6mYRiR9FYrVNYzKoO98R
YgvwQOfx6jqQU73qwKuWcYdJXUSo7/SGAKSKj0mcaGVeD9hyxLTNTuKOSyQZAQdIhxY1uN0jma62
I9doY8H0uhIWGKrjamHfcBK78Q3sCTiLs4zylshey/AuaiyWq1iS0p1OJcreKTG7yKsmJXYeAOjC
/M/7s3UZEFqKLJsaNdH4oF+OL6jzqzTpxSkNTb9nNrhWf+qZKIUnmTazX072WtO8vGb613WCI9bH
/qRHjiO2amyPe3duh87v7U0hMGlVCPU0cqc5OKnTUkg8G2g5eVx92o7QwR84Lh1lJb16BhzBZuxh
IQP3kMRn1B/bunwGbkDHMRh4z/m11ytNWeukqdHU2nBA4u/unKUdrMf9W+IqCEjUV2uIs+MCkjsO
vvzMOtXdfnqTggnDrd5j9mUYfXWYKbgQLqaEP/FHVEsEOXau0SWcgZzYddSib8JdlI1eve52shQT
UnmjQUZtyA0cU9NtkNES5XQFuzQPj194U9u7c7tEvTznoYqfNX8QX2P7Ves3/bgNO+9sxAus8pki
las3Eaj2mOwOW4iXkA8fypWzXcDNvAcT8G073y+sL7oEvKzVikvMuYKe1ORzI6j5NLdrURegmjlE
yk0QjclW0u8fiah942oNDp7ot7th2kAghPY/4OTNZuU+EZFgQQ7DDna0Adla+DF+7l7N9whgjtKW
ogfK3mprNA4+qTu8PNZU4ZBziiJfM/rIicXunJ1jq3O3nam0ELzNPzaWSUys/gBz36UOZMCcGjT1
7ijFfTl9v2JvqT/xs5Rv1iJWAqU7KZQheO47j2uP/zm+p6UGehUGhE5Yy3gO0EKz2C9j6kSRNykh
Ujz8+cZwPi+E/XLFK/RpPBMZElG8L0dtkM9nV/lZDuCEcyJWLco8YrOnCmbxguc8q0k789QPajq3
mNIHjERLcZ8oQkI6oenPcbkU7ACOmOZOd/HXU1/F2L41AOwzCA9i5qjNlDm30i+MPk8Ti6xYpVDE
zQhZ0NuI+/8f03yeRX2OX2ZDln54ySia92hkT1eajcTRiXC1FRGABn77h20H3qmPy3JrdMgG72aS
N9ek6G2AwMtBYwew2nsYZANwusZ7LqYtC6svqO3pdOs9AJQDIUoetA5/eTE5oSgVU9p4rtmtgFn9
xSAz8vKmxOMUjAttJDahXwpW1ieqSpgbkA5pbo2H9vkWTXkqEdsgh0ayBH8nIU7D3Jvy393GEcm6
8j6tR/3qnUsIat925r+R1cSvlH0JaKCkwjvHvxYW99XNsoFraCR2ihhmnLJMwRkxPjTZjjSGhAyk
4Kq8QyNPiUu9B9I7zuMgldciclhu/G3BYhDfjJ96/e+7MlKnOn0jV0bVi7I2y/v+jQ7r4ubGewbw
OPwR3FyePj2lgaDoXVBJ9ZXLJJXEqpben+AIi8Ah2NqcWaKF1WZkbeVXz3O2LvPbmAyF23SArP3i
cb5h7GhlVYvjU9TsP050EIAkLEPYxDKGT1A0vGWP7yAPgASliE5xu8Ino4Mz4TjTG07B+6kO2LkG
WZZyn8TkMOyjezo053NXHse5Xut3QJmtz4neQN05yktInwKuGtwQZGed7hDKjTnLnB00QQ3IJ8Or
MdtD3HJg8wmsJO2CgjysWAa2Pys221GBSE0AtmVeCV4cClIWUIFOunxBxXs2KKRTvNVit6wpCIrP
zE/0jla6XlxFNt8jjbGXYJ2IkYw6gHS2CsFb2Se4elsPVU7CasM9FnsEP3juA16oW5P3OXqCOSo1
PLWOAKJXfpaobYAatS2x7MzDPKQLbdb08u6PiXBK4wFEhXCkHlLQ0fqUqeOhHl+e6kO23BS8l05k
0LUURH2Ki0oOXhCykpyxetQKZqbYRNfzxdlsT3hcxiJzt8tnZNZSiz7PEh5t46bsr2a1xRWCjb5B
sw0WXlD/o98FxHWZ0Vu+YX32oVaQ8HzUbUUdX04ZfdcPUC2ljq3LMqTjEX/cDJgUrymjqZOTZ74w
tgDKUQaZgJmilsSo4Ax++xYLid2SJC7ygvIzFnG+uCPtkpcCtH9WKBEEprsjbD/ObGrpFX//ihqH
ErB6bcaDSArlSdCWk6VXsKl/mFchMKDrLK4gGYxnQTEeKBlEoO7FZ367+TN1Pd/EKaoylu3YCg9M
msqyncMKs5QfbrfE8mM03IcVaICQsR3W1ToE+OrF/xJSZjGQHFsNvosSD2mARk77/G8quPrCSDUv
bgkZzUYYB7cZLQYVaV4qTJ3snvdxOJrCceEm8PHkZWPABwyQVdO2R+kGwBGvqwOiJpKH603HcqjY
JNG1gab9qUpHWYjkEVAMldyGEY8skQGH5lkRKGXO1x98VVRrd/Gb393RM51hd1tvy3D3H3jM8esy
jU5RfkUwV/fDAbN0OORpsRG0mRMknL+tjDdgik/YefX/Qmf++n74Aevvv2T8lHU5FSgUAFLQ6AFi
LUQVP51tXVNkAZpSukkdDJ4APk4NiGjAP4yVogezLyIDufM6f8iNgPMRgCBgwJ53opqylfWzeUXT
pDAhJRbPDS9w62XDl2RtNCO5ZVxzeTf+Xr5APQjtX4XU+T4B3uJ36DazNBamDLFLjdn9eVN30UDF
KbxSCHh1vi+0DVn7gLI7wmFO3VKbStGQTXhTFSIOkaH/Fmyfq6sYl1pwhP4QmM8JJuPVwN/JCR4d
g7DHBXhd64lJ8XA1E4bLRgciSoclNb2kAJG6NgLEHrU3TseMxjBPX5XhXCdAaZPo+XCwol60PmPn
mMgKpVYV9Cqd5vomtYQnwhMBoJGGw4Sek++OptGeGxyhTjoKoYjoJYIg/d+8OAAP1Kf1eDtV9Okb
GVi9+vGlzbNSFdMHHONyqlWO6rkL5Oe/yjvamQYzf2POzcaO5O00ocN/CAQ8i5hAqHtqzAq/yHF9
ihl0mrbfc631UtQ3MyIJRjG8lCr6inAt93etgMoNUSCtjxwy3u7a68nLWIchu9K39C4HxqoOa07q
jRl8Zem08+K7eOQMXzo7qcmfDXnN/7jSzkzbV+vapDggo7FRdlPHt1VRJV7N/KEfQE837o4uncTr
UpVkdYpFrMIV9lTwWFrdsllon7qwO40Z+vWlzyXZPP1L3kgFEkYSEA+lXHkfEN6NYitYlkF3ulDl
OZOWZu97t6k6G1pEuQPMj8sMYbFiiH6Z7XEmO+xi/1Uv/k9qoYHBRgNj9PHzAe8wXAXw1/bU24im
K5ARjgijL6oFchhWn4L8gu9Lu42IPgQQWYON7/jtQWSazYj/epsbI57Tdlyfcn5rCrwbtBzf3ngd
JMszQL6Qom+uEm++Dy3PaZhNAvMpvnbbuC1+0BjvkGzVyrKqjJi12GQd0sCEIbuRxPz2QGZgbO1N
EwD4Y249mmoFUmpHDhuWmthysDAxCGpP+A10gPWeFO4TrYoVK7Iddp0s3MNzXonReg++WmFIrSKf
Jz4Wr+wb+RAVRUDWly94mTaWmlLTQeUA2Qt/+oDwIyKSkyjhseusGC94vcSBKRERT43Skmf0O7z8
kiUJVvrOumClegdZb2luZ3JGOx8alBJ1PPD4lNMce64xw8574mHmm7krl3HGkPCORUAJVymvKyfk
reLTubBO55DbvS35p9ot3sY8uQLPPPhkAZ8nyl1l8sacPlmT5p3oShpHHOgfbzfwfzH+IK/N/UIm
V8Rwc2PhkgNsw2tw4wCxyE5afRk2e2E3TPU14s/3NCKqWBQ8v11RjDtD1OdXOr78gFwZo/Uth2Ar
UxWzZ4JGIeqONjqEAl2s/vD3lasP4UNBWLB5avzyvKTtqUifuavZbIJoDJ3zeWJkc90YweSz4I1F
77LfYpEz5rLd9zR9tPQ5e9WpsuUBz2ulOlvyxAdMcMbYTKC6nkc5aQq5iZF7W/9ssYaltMSu59ub
viP/CyyH3KAMkxOZ7TX9PSSL8/Ly9mSk3lpFXAIxma0ExBcN2CddHiA4eXn8pIOLXI99PkAJm6eh
fvYoQ8iBeVdQ0U2/oA7l21/w+aVviGLNNFnFsiiUnq80Uw1nnHM+B+f6yKHgxxF8S82hCfHX3bIZ
ElDJ7m+TqUhF1NKlDuy1e5k9p8aqCxCl2KNlQ1cPY1HA9RehoqyA8iUh/uSMBP5SFBvaRFwhuzOE
yknvLkmj3i3Q5kFWBp01RE59xqzpnlemZ4wS/cXLYcfZ7lM57ttIo4jJvVJuuBLoiixh3dKFva5V
V0/5TBlKaqeidj1/7YXucttvZICadz/Pnhqa68/a/u6XBA0Nuvb5i97cizdMh8hALVWu7LduFsI6
NP6ttWfVlPydwb/mE70csYo8oWwZDsI2TWf/5i20WUxsRzcC0lx53CTwwCrFLfgliTYVqimvkNX7
txBV8RTEfnfWyE0TJYcQDTeA7atnuaW9TOSuTon3tAK+eRTag6LxcQm7VPFB03KbX5tnPdsOY1P0
xHo2lMC96WMqyxeJjKlUuZY6kQ9usFsk32xB/kZSe8rz3e9glH/E0T+yiTy07FmG86AohkSsQgSR
ubftFoczxgz9gS2kYISkQa86ClkbGWmI63F3oh5uA+1X77xwxELxxaLH0tE/IlRwIdoXkLssh29g
aOcHlJt47sRI4uViS5sqspte6oITFTY/jzvvi0L0e0pN6iTFCIvTynxPoA6+B3UAHw52EkWbjcLS
jk2r/hHkJtePufiigpzLUBam28QSf/CEfbRzKNChKboBztxgir8XWTXRZi9tWB0AILTZ/33z5+pC
KKhPqQ4LXznvg9WoFo0HdTF2aM7G5aec0iEr9I5pEK2l9qjPk2pAGGYi+EK4hgHVZ2IeQui6JA/g
mOn12ryRzrsX+GMHf6RMOApsLnbaDftKK8o+lVY8RMWEFMutD3wxPkfcdTti3ENjQ4qLNFieRJub
sRsoauoeXMJ1Ra5ZM/gM3mO3jOY/OMSH2+uJ6fgNmhgrz6oE4+quvexntxH9+m7qSznohA7yRwxX
gr+Fvryx3hI5luiXOn79eaPSFyoEItTulbtVFgz8A7N648ruN2+t6oLirWbPgqGZEYL/91D0D9rf
gfiqUUc7Eo+HGMaDtwDDsCsGnSRyEh/qe5QbYfBgVzFyYeqST10JwB/QtmNzHVInI2LB73Kmh1y7
IqV6G4YkzGEz/ioxuEpAvQEbjZynKgii88F8WM0a8FVQU5ji8ZM5M/RG/DFOL4jC+2TjlVy/hBxf
MOpB/XTmzNA/Xee0hIAYVCukMYUZRJbIX3yEXex2uyFJ6L8l1uLqUaeE9RmP06tMDV0tjtCavxyE
autqQSHGXogc/rJid1STMHom37/TVwUJwDTjhpDgCuamg49V98zZqlUW4sEQ24uSqNotjlVu9fo6
kzqSHFgheyHHOD2nhBP9o+m2GJM/doGx85p/sM5yiajOSZQOluJtKux3QJcbyiiJ+NTGPtb/d05G
BBrOIICtQd5ewOCJ5pP7gMc/7JkUl9PJnhSlxYICcPkTOXtyk7jPFScx/0t42iOX3XkvzFwD0hcy
dLmDtx8JMBsHEJn0TvrpLDWeQhy90ezfY/Wqr4akMSjY5UGauEyiL3qFUefVeOTndDtOfgE/DwsB
12lDNifLaJl0V+hzYxum3k0+6RrW2pZltmx+VkQoyyvoz9BwGduOztdu+DqLtDxQnN09Wd6eG456
/422QSayzswi/xk/V2FB8TigdJow3kvY7oXlW3XVupPBfHMzMNy2ns0M55vPBkv618/Qnm2SGuI9
DutW4V0ecwgavOHllNKxze3MCmwZcPYkmPG+XZNDscb9Ehm9m8HBvkGyhdguOEGuRFT/BvAq8cm4
JXA5DEXav/S/HjpmCZhQL7bxpUJDP0Or5ZQhGWNaiKsB172e/TTSiK4NOwgKcJwU16TvW+bSXhOs
0HFgIBOww3LTyC/OTWDDPDtZBHWyH/pY9ezruN/G+OLLf8qSCVLefPVSLLUZ54AIkaAzTcP0AOk3
p958z71Cvo/yFKp9ZnO3hiU9jP6VgrMQZU6S2kmixTJyi1IiwxV1N8+5NIwSpnGKbjg1iambmTbP
bcrG+RgGzBsXOEY6/36dByQgouTL9HkdHDYqOhC6Jh6gKWlCY2NkfiVzBNwxgw22rgDJuYefH0+E
Leb5aTT+vD0ynYM/xkFwdOxUpGHLwtGtgTFp+0Rq4ha3ceadSStxD8ALc130tBR5d5gBcx+Cqsqi
i7lKT/bxOSDuvnTHgBGFSxNMtg9+FX+Fl7YNhUx9YX6Gp6uux2f+JnPs+QVVqC2n5MQcOeSmmGBW
L0Z2drH7lMgJZRztoKT/K4iCmpawLAT4XXOE7CYMb5+clmgvfjN8f+tOM1pMcjt2PDXjxCRr9Q==
`pragma protect end_protected
