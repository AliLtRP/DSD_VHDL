// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:31:33 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
f9lt3yuSD2LJETcV58AecO2U6AQJ+bcxV5CmyH7S4LTmqo4yNQPWOh1mTc/tdfpA
fUsrpXE6//QN550iTfPEbdcDm8bilVjQsVKsxJIlRthtTFoL8/P0/ZIQ7GyirUi6
hqH2vPsdSg3gb8ju8QrcpSqUO4IpyAXUdKPWC6ikgqM=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 3264)
6dR9/bLm9z0G8JyuP/vDNPWoex5NH5Xv5pcMRzrS0oLx44K/R2dV9KmRXCNmLklm
CG4zcAVdasJaMg1Ml9skfn1E6E/bY/flmPWKXXE7Er8WrPog7W1c79qwhFJjhvEX
/OmWrLlTBOwPggAvbSdE66NLnQebpu8zAUzLT/9RC0WBA3evfCuJ29tfkGxRlOln
jemqMFSbay6RuCtEL4ahiHJA2deh7CrcnGIBo0ImySo74ujvXDT3F03dTvzd2aHg
aP9g6PyAXTplTOhTXbXVTSGPuAQ2HzmIg0mAtomAj1woCtZVMuKBY9BYRTKX0EAf
JmfbVTjWenJUi6mn4B6wDaZQV7Nl/viXVaurxnmtaS+5DqFWZg3tq3l8E1H0uxeb
Yb/W7rEgLMh0IlrIP+EZe+F0SzDdy+guGUpoCgtApxcJUxIJLjh2V73ojbqjjsmM
6DeVyYgTVf2crWz/k9GCSnG4uCC5qK0PGGQ2V8l2Uxn+UmD72f+3FVoDkRfm2fpN
fYUj0MdmqVffTos8stG5FSgV3be7cIexp1kbLkO5v+mWdW8FPXT+tydpiwXWtCFl
d8dw2ysKJ410lDlPxiacA8uwXY1J230uttXm5xeuh5gWomsfzR19EtV+HmJgf7kq
89fgQU45rATIzmfruzMAJWynE5NgJHjv5u3jlqf3t1lbH57u9aN9XHszEXiSbjmO
umtdLog42hNNFDd5c32jtihL143T5hZHk/xqAjJlkO7h+P/NSqlVN1NntEYbIDGY
U15JWlarw/76kH+ZKMWpinJvVPCA9gjMNb/ORgntx+x4t9yhL0H56Z/SUc0FyqgO
h3xwx6x5DCnnp2P+Z2z3+9N/D903prJxCGiCCVE7POXRRzCJnrMwf5bM//2pOk8t
IFxxN2sOpMTx2YzMlX7ZO+PZiUszeaR2mFMKiR/DbZgLQ5j+jPTmBcyniXW4p2YD
mzkSWNFlObIEIhWpEuxM7KNpk96SkbnmdJt+KreOAS2W5V5/INu5ZF4kYCteswn2
PZWJ/Kd21BOMeDxo2R6Wqksehbe8krrn3TR+4o6n5bF9VA8oFf1n0Yo+0SfEH5Ot
R/b30NkrcxOPzg8i6oQi/cX6wDIUY1MbJVI45Lw7OcvTJKUVPaQSMJMfa+4fYIbM
XxBiNFJVEVXHZ/2ZKKlY/a/7xyTkhcG10eGQGz3P6dhJckk+qqpdChrTJY1Z8PKO
2UzdIXlk3z/YECTqdfyTafd8YSWDo5izm4Z5PDMwqDujTzJiSFS+V0vr4bYupoFA
bM3KnQhTt556WrL+KbDS3hxVW0w+6dlTldMU3jlo9VmrW+mqK02l+CLwSeG0JxOR
GQxpbGz0o9Cui3g/HPv7skL2ayaQJn5y/lwwO6iuCbQOCTfg1j1EUrNJVKDeANSH
oWrYXZp2WmtUR0FkuAnAyt4gyYBMICZiWd/R9A7bhGM9zerkUOFJgFemm8GLQW7C
IyMVlbKUeqXmtHbZE+ZPTwDWoxnZQ0TtgfzacbO+26hnC/yL0D733dl0mBV4Xo2d
TpfKyCsPA1TCdcLY/3Adbn+zixZ6qVFfQO9pispPbES+Frj9qnGw3iyjMycQg9u/
j8Z8+yCnmBJteFVS/fV7yXwgHnJag65W5XCgaaZjL5VTYGUgx+Z47msNAh+EN2ne
LqYZWy597YgzF/M2eGCC7fw+NkKUOF8RvDBNWhVG8PWwSzfUxUmrTWi97tlBSTv0
Ee7qPW/VJUvGSCW8bSRnxLlS+zIsE2n9CYBYTDpdQqoQ0QLm2cMLMaeuLU0dFuhO
zM20YBxN1HnRtTRroaUJ/4aLRa4SbD2U4kj1ecm67HMKewSPZxOi3c80es/jABQT
Mzb9PlJKy0R8fCL/ZmqLMB5NA/VOEcFkD9wCqC6+cvY/s3WTZhuKNlUoUNAtmXGS
55QnYstGwmL4uz269UQlQWi6g07T3LJ0W2GhbjkiHkHZgi4tqY59oceuJmsw/4s3
HbdanTVrD8MQlZ/vGfTpwCr9cDzWcEuB+fSCcXLm2UheNB+MLPkG88QpPmsJDxx/
asgNKiKDdmm6Xzz4jELSrDy/FZaW5029etGCuuErpv7saxQpgGdZbcGOpcr35jID
1ld4JL5PH4RvS9ssAdKPO8R6/ohxTNwdbbazaYtV1V8b2U6ZznGiDP6mY/b5QOPn
GxbO8BJJr/hUyiyIAM7abyW9wmXQfQuEMOGIX3dD5jmzSG9ttO+UkPXH61Fnt+/Y
5GIMdgGKDC7NKhP3j61h2jnbWiVn2IDsqGG6mO5e1whqRuxsvptnQ9Tn3kdEKkOZ
u+SM0MkwLatKdDGqUoOtklbeVIvJC1lwfgz+qZ4CZcRWBWSR7OGOBOCAhxjRpDjF
wdwuLUNQNFc6FlQSWjTdsFJcvGeaQJUEe2kIpbvFjVKuHbXFXnWayEXSWtJieYAz
CNy2CbYKmbH+u0vmJWBLhh0Iu5ufc//vwD39NaD48yLRxSu69JyEnVChOpt5CiuO
57MG2p/d4tRlbzYENXPNeezFiE4h9jQ4pAQFncC3fLFpVvOsvAmAW2sQfHkJSLN7
K5MYc6WyrDrdjni3+NKBNF5qmAN+jQKg2B0YIon90u/U+gjsYMSzcWYLV4XZtkF7
z1zCk8DKusanH3sMMSKoYcdGV7y7BOG/Fw94zECtjYC7e0JI0UEtQ2p5x9avz5lF
AKZhHhHQFYFhoDbUw7HFQw8+S3k9HQWA04Co7eu/JB/773Bxj2m3rFbb5zXEe7hq
QOfMp4G0vuzY9PKRKUFwxYSAhvPVGN//fIysCPKCtlQr4PI6ezp+HVfeRsKOv01y
9cmtmiOuJBJAqYOMvGjdp4sESM8rybqMUIDUqtVDRByL6xEFI/GDKnknDFhHZ+zT
f9cX4MdPEJMpXl0SIhQSN49HEU2kOwncoSnVH6mLj+S4EcETkBFAVbt+zCW66ttB
2rTDxbXT7z6iQr44b+66YqJa4ArQvnVu7vLgKYUQL2TGmRfh7m0MSHJOfgmf5i2N
TA/mSUY+bGn7KayBNsmwG6Z7/e9IMZ5WXNJaR7x8rJvxGNraIHXLzY4Q8yrbE0B9
unESmYUzLPdJM57cPScAZY1UK5AAj1NHHCApE4M9VZjQR4fqGFDenUd3ZUlHHwm7
2bO0yT2nnK8OJwl0ChGyAS7K7Huv2aJ5UqQ6wV/wT4Qx8oNYYSri7Zi0iD+DDgNr
7jGtR2tAYmvDxJoO4CzsAblNoW2fcESNkArMxdqaeKLI6lejpx3tQpQe1MlwJHYr
VvqiHWFDGUcKyZ6MeQk9L0A1SBMPtaFfr1niS5F0bD3UrAdO6DVzaLjVVVeeUrCo
2nidmZ4b//rvFVkl0kDlLgREURaSygmT/3/++u0HVzsuXKcPxvKH10BhKYPNRaJS
se9/hzJ0cSkbxarK8JYb1cpTzRy2HblYIOmDcB5yPFWKC92Uhnc3TrNvuwACPdO+
24sga/oU/ptBHVqrWEgJIUVcQQINY1GpO/LGEbJi4Ck2QO16aWHVEPrj1M7Ex17T
ZQ/hr0lMNRfywHrxjhmxjmehtAsUGyjWAvaiGDea2ePCON1x5AU9xQTVFyF/dtqa
Jyc3M4j8AjlL7u93/uaqfYlfZEP/f+FERJiG4YUHCYkgMA6K/9Apx+DdB/gKflaV
Ya4xvRtVuSQVb2EGLZ8F9YSW2HHCvYiVfEnhFjVIS051CHIqMbLOEzzREJfjIKNN
8NfHJB5qMqN/B/a0RIcNJfAAI2+mVFDtSguxUaavcSw6kB3lCme+22OaSZdYn47K
TiIL/NJFDbmkC7Wnq4UkFII37SvVdFvyhOrvXRCFYgicXF+AsfaYO/vsVqx60aDk
VZnNjyrakLnBBwIpkhQBbCtfDUnWR+hGx2JrM6YSb67RoLq78u+Qiqsf10b08Eyl
0bw3jVMqtMK4Lb9oN5YX8u5w5nWVqqNDL9tZMO44Linw92qsMEWrcfJk4V5qCj/o
WbYqoPh076Vb6ziEdNh5aCCLBsgsbMvcLMH1cl93lnPmsCIyjv4WW8wwhdRqvv6X
IXM1jgNr6/HRwRDDPdfB+0OgYdXw+s/McvLkUFZKCJgi7LefKVCHnDfAZwIQ4gvZ
Mr3Ut82f82d4TQzitK8s7+QuEni24RqbGQI9wuYl6VDpE4LcfZy28EpawyQ6qbOY
1FZz79tYL/7B10iIlJ8FbJkhWEpOUC0IFAiMrkO61jhZ9eMksmuN05fdnEZ2RNIN
aSx85ToyDIGs15E25KnImEfHzB2x8OD62/3u28Gfz66jmF7jIXNpsNnB54wSBFT8
E4S79ghEXrmonsW8wZbIlZejFO56nGbImE+v7kwv8yF7yFQkITUxsu/FQBtlRr+L
`pragma protect end_protected
