// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:35:34 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
e9wlRRrJ+dxDv87px/q4KhwzyGsq3yco+L7OCfmlL2xs1eOWoHZx/86gxvXbcBNt
QGkdAO1wxbemFpf9l7uqmEsUuh/FRcCaTFvPcGG5toht9dDvpBo5zmivzInaih3j
e+BIsPYtNwclnpCi4hBiYv0RJABHPYiMaknFU3FZGEc=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 11120)
IMDQ5s9hWN+YL+nQQilwQiTHUvZ11D5rnxRumjksKwqO7SSZ7ereUr5f6os8Y/tg
ekX8Jwzu9SDUiWAWB9y3o/UQIsbr429EnFuWoFkP1lD6h5VzLQX4gpv3cGBk9JIo
JqhkhTNVyLKQw7qiRpbObjwjf6l4F+w3IW/XxQO13qucdjQv9tU8rNHtcEHo86Sg
XA/baNZdC9IpbxwCWFFZAy+MO/qJQHpOqrebIBOxUsRxlEXGomc7Hw9zYMwdAOCJ
UJQD9SVQ4Ktz9gVUKalnhmYKMhCqD0YiqfPMZyuthsVL3v9vwFz7cYbzdEaRmTHi
BzfTK2tdxm7qSCJ00O2Z+6GuCttFgoHtwee63vWW14UI+lCY4hwdw5u0XEG9Ely7
fPSVxtbVgXnpnC6PjCVlI1aVXHQ1b5U+90bQ2ITYYfOKw9ULQj4odYrJzTRnzOjI
kIaO6m3Ftsl8/Rb8+8hsMoEAOjWAA6N01suhLBjcfrW4v+OWmfVcgDaVwKdZbrlc
mLQKrMcQujv9XxdIlD2HFW3yF3G6gmN1lhTp+snVpR7pP7XmnEUu5mpspMFt1fxW
UtnealnunxqXtUX1KQPz28mZu+2/0OrG/NZTQT58PxB9KoM+3SPEB+eUXak1xLuR
voz1PhG8b6xTGkMcM6foiMNhjDovhoS+Grmww1DMPeU4R/KwnvsqdRNP/fsDgCO4
szTk/PNDdyw5MjL3hfJQD6285glEH+Vc48XVD0SM9r5WXbg1dIcq1UKGumUeulNj
kYqPPihW3AmDTodqckcgEkkWytpITJLGLFWAMSbz2pSs/ePDQdV5Gn+Svo0PXRSK
06NvWIK5A3mT8aqSZsGjMYlgcSOOMbzvuJqL1A6qp/udlspwpf4CAK3aLwdVV39L
3q0K3LAokfnCHLmog3Wbx3HzDnf0q7TcnGZomImR84ArGT7TZHbKvwwQX0OPW85R
O3nmXlPY8m17GniiKz5n/SHjRsn+W8StdOSY3ULLRLAiQdr9ch3s4BUoh/FiiLX8
3vHFoipcXWeOr189dwSSvrQJmvV7UxYRxVeRWMCRuIk2cWzE+15D+d/m+VQH8gac
juiTVEVwEVK4VkWp1FJix59rOWcDJhAqWZyJ6rgqlW6voTwhCKjlXUExNhl8gYME
/3fzJdSi07boM+6WQyoDekWfxjGY8ArHiUq2HqbYhtmZm+sb54htMbUZyAcnB86H
73rsL47+fy1JlnG5oWDZvueYl+BEeGGnfCCAZ7g7lfHHeVHb+7rXerhWGy7rSv2r
tfTTPSNjUv52VBy/tNFt7UX1sv/UVFYRN5FD9g2wwcyghtKUxte/wTS4k2wZIWHu
YhcC4ImJbTPO6HbG36wtsmloImM5GI4qeVprIw/oPiv4IkqodBzslfYsD4qK+rKj
uaHk2rStcrKUBUmxy32xmWhjQCfdaFVyRkIc5vwMXPBkm3AvXoGjLkKiH9HriAJe
j/I51cJKWmbYrcO6eDjh5Y1t+v3tIR+NjxfEEvwXythCEYRBODYjFMIxBLL6R1xm
7rRBylLY/YterOAO+bNjCSpAYb+GIYKO1oQzusZhl0ien3XF0jKfxnrlsWWK7D2x
DjuNTQQ3BlJgf5Wr3RQkSfcJKumrUj3U2CO6uyF29L/2R3DMnszipCPsZxRZwt8b
zeQiBGe7KsDjIUmZF9DBvi1M6M+uX35kuf/vib9zJhGX02Xh2T8qdwJ864PaftmP
PkBB5MrxtzMtao4cLzONUkS+Vzgg4PBJcJ9paLGKzEnTcNQvrHiz5x/dF8glk2KX
AUo8UnGwvB7QUnGwpdNOkhuy190olZ6RwE3mU4Ni9VMz2+0UgSQrEbdF1KzNaxEU
nq5FjSx+ml2sEM41CZndV1na/RLh+dYzMxLcWRTtLFWlmNMbhf8TEOUzKOLz6DVc
t05eq1EurPKWcb9gfD/HnpxzOE1/ia3xJe6gezV6XOLQEqvK5wrMU5mIjOxfxVWi
mbGrWjQjWDBZJV4aKaoKH4Bhzf6kkVo6r0LHkZCJLPpopwHK8w81xqXZrKj5Is7m
kTjXWDw0gVMSfaKUnZsLX5LynlDTybl03FJ9UR3GOBs6Fu2Nu2xUwCsR7oEvjNI/
83qo9PIAL5ZlXwx3rdeMPqGGARZ+pRb20zQcurQExlT4lBbTJBFLQ8A4MycXLRLe
46H2zXZUCrieLRxiAIi+l2fTO4Pod8tB+ogDm9uTF9dKzvAxs0VGG6Y/SwIeSWSA
p+JIRf7sykPo7lJuAAY+cBXd5jXbyJEw0R8Z4Jr4CF621TznbVo3ctftV3cjUQsn
otyX3QAevS79cCgrd0AS9id6qzR1XSNTaC0XVnaQ3JexxK+Lk8eO17gZv85KKj3e
R5tAYQaWd3r8jUMKWJu3kFuijSGo8LoJ0BCJbfenQPkMJrO/H+TzRLUeTP+srSzm
JTdbImVIy5oWBzq50aoUysCDSvWG9MYPMWVbJzde/HEaZzGzAMcydb/WpcrFhzAE
Ffmj6q6ZmV/YcfePteBVqcc/ikwhL3RfbulTLmSU11bxhypPvrSbPESYREDjlStB
y6n49XG9bPjYb9Sa69YcI3PioZY5ltsdaWxa4hO6Pi2jGFDD5LgNRZSR0LWdloq0
G9uyRkN3X/SaVIUDctLgt8gB/p64cr11wWnlttjIYbOP0rLrc+ni8sMjZxW4Bhf1
V0r05desTUsGv3qeS6tQuP4BwJRbdStkWsHSAYoNELsP1FiPmMkWo6XcFiXVUACl
pL9veBeNO7hUWjBTR9fQqgQ5Nmm9sQ1dpJHkNAiIhYQ0Kf1jo4cfcceaLGyG0+Hd
0yhT+exYmzM1SqKmt3BUYd3jrEmY7YQA8nlRzwpKy1ntpEO3OibsV9z5ACBUapqm
YQpnhQHJVvnk1BxCxVqDQuHKLybpNdjBpFrodVi3PRAa9/as9Jqx3CaxCiXy2QFH
ajuJG2LMASmjcIOAg1qAk7j20Fk+iGNyq/SPkovh3H+mCngeV0y2NCWtSe3Mor34
Ra7XL3c2F/vgoGH80xekYpwDWn4Oz3ndBK7l97kbLwTm0jEdaFe7a0dt/o/tCCox
1DHeNUFeoXOWci3ycm6MOIbqQbCGJUKVJ7JFTzbaiG405rS5A7esdWTQGjefoqvv
DivGA1d9TQ4WD7w4XqLvkwEonLqHYzOFhmB9Mx/ajz5fsGYKXFunpklw8gufr7WQ
JKhC8HINvJ542jVsB0ChkRZNryccqSzc9Y4pq0wcz1vVrBXCU21sVWnmOk+w2YU3
PeFT/4MfEgY4Xnz/khA7SvNfH1TdfOcteiZSt3Yw1+dbKT0AFIGaPIoTMyupwI9P
yEMBRQAoFNnsDRVYQXRZre5fk9kMb9EKjA8xyCUEa+7XJmQJ5+FnRun5ltyS2xMJ
c2bbtKjCXHT8DBD6K6f/wak0Vs0AEKmWbYLfp4w5CddewbWiHmfvFwOj6ch+GNYg
MAUpj1hyauygA9dD2oAA9qG5zA8ZC1caHuW0cyyoiN2PyhQqpWrpRhuDimHDqqwO
zDJKEzYAHLaQED9hXFOlwNC0h/Czl+7mypZN/lB2SmKna1w24oQ4wrGymA7wirON
gLNeKg05Vdzy0UdtnLSN6GP7DsmCQbMBw6e2rQxjJ5sb23TingeRrkxwb4NNtyAu
oQhHSK54H2qCTvRLAu4PD4GAQ5n5SVrji2FvUyGyPdg4uCUa5mJExK9NAaFptqN3
G+QgaluhldCtxaI2ErHzm70DLpA8qhx09/cMcL9B8RI0lK/X5h+kN89JcoTt7b0S
UcNnhMFZ+VisldTaup/Hn0KAMvtx9VqXpHoWH4JVWAgMMCv8/481Msvx01RWJAUm
GBgHRgnoLQb3v3IoOMHH+KcY2aKT1BUEztiGFoE/RJS+qZcnGuqLgwL2VWmTDkvp
K8WqOaFXV1U7ZCRk4iXFyn5RRk4OsSZb06eQi+d8ZySs4whsYUTp0/jIeLS/Fh9Y
mIm4jlL/Q1BRu9SlR+0HqwVPKqTMdpQAPvyT/HYN3uaiNn8b6q2LTmBc/wuDjh2G
grplMvbZfWL5qLqvlJ4soND3mrC6fb1QwB1eKTG794it+xT6ZHX4IyRaeiS1xFnU
wZn9O4gFwVyGpFAyZdWEtVS2WijAIgmy3/zzm0D/F3S5gYwKmthYFrWRZ+fV5A18
OpHvx0PQmbqmi7fEy0iUSCkI5Rt8agHMzpWYQl/z8LnZMtrrv0do9ahCtelYyLYf
pu+eRqiZdsG7rurMhRzFxms2FtMs5/0fWro6sfQzPsA2ZNlAr0nOJ2ynVFbDo4ka
W1BVgBe5EexzdtYULLka8vhYLeK/rP5wkIO+z0EDc6474en2Y+RF740xhS5xrMSN
UY7LxcKjdG2bEt4RxXXn4zJ+T73GyWoGtLhLmbe8emChK/8tD1VVYqzkG52zOrFR
PXQwNhgdfjHaUpLBhAGvbccyHy1cV4yTLEa1YaiAnODvRmxom57UCgR0B65CgNhf
5nc97M4ooJSPMgkAgUHgiKzGUmQ6+5zXY6A1Id0lfkVf3otJDfTb3vLeGmhP+yMy
U3ABJ8mhxB48peEsAyfmlmT/s44yvr/VgmnbXoHncCFe8ukKmWK3IOa6wN2efhn+
2fdP25M1iasknZC6LZ03m8TmSdeA8X5Cv3n1reOxDq7zDI4FdvCxnBeYWxxuqsH0
8yxmLJK7fcvOgP8LQehoEFzw1YV9FykraVCs/1xiqMwEGdTRarzJlIFGazmOmxdc
RRkl924zSXStEcf4oP0XSoq0URI5iMoaD2uQA4yIKM4UBtMSSEArhTl09sQu+E4e
jPoqpAB6+TlCKjjtONBVqwArA1SqeYlH3WCH1jrZ7090sHtr5DzRCEUFN50C6bI/
k/waSNju6i2g48mbT4XrOC08TQ7ELRoJ8dUNxbeRGHId6HWY9Xvie2i/cbgxYNDw
2hC6ZshCyUVLDLGeX+kgQ60KxbtKXvNhnJZAuDxgay/gdzPy+HZ762sGkD/65M2O
yCZG+FKUsbi9qMi0k2TIiWje5Y/7Flt1CHRgswGtawhhgI9QG0qw3h2U5wMwKZ9Z
JwONgew8ANHOslM0CNElPHX5pinlreuihlL5bGVDgxtrQNZIfNM4uA8H5gBj1HaL
gzPyygKUqwFeDyOjPGgB0ydlfJHGw8uBonJosJCzQq5N/VSDw+ZSkHr8P+Cv322f
7gvKuHev3GxoNHa0VTCC9nNxhJch2fGaJzBgH+58CyGVViGEj+ups1pU97t871ET
rLJ+OtV1vosQ5NTpUKgAz0G2GpATUr+6aU9jl6ZtFCxCy9XOfdbBKpb0HpD/FiBX
XQviruhUpLJY4Iz6Qc+WjAoWA7EVG6ftiUFaTz+ZUZ+SI12L/gL030T4FaYJLbbd
mDq1y7CDAzf49yDskngrACURlqUk5GJHw0fWNKNwPZt2zxvIIQNg6eS/EankadO9
tkrlrV4ZLr8LcLMdx5AhqBG92YgBS9cuzUqq+pyab/zDO8L4fe9/+6virnnuQWvD
VRyPpHKFHfSeLqlag+alIQYU9iew/sqL78RJX52p0uqnr1SJ68qxQW12mwvGnPO7
dyiB+f73/OwScjmkhIfZfZ0p8/mOwRhiOtzNQoKdKosOqi9Y0fetdux9MVgRj56U
rk+7WfPNcF6PWwliY71i5wRwgAyB0dqwfV5QK/+W4o20ngc3zLectxLGTf7cZhSA
h556yvJNQBNm/YB9Y8XF5fmrx5zcxoEIxFA2FV/1uIfk93inxRPDxBjxYsrXH8DV
198fcXgKVSoOllU96ZjXlTw9K1cpGnxstdjwTU02joAgECCXBz384qOWPTYPx8Ld
DSyF3POMTHYgv9edh4RPC2oJOnRa+AxopN9YZtdXuwbku34G6dsCSEB1j4uHJBZG
yg4a7qfwbikR/lCjpf1wpUX1jR+8k7ue6M3uTL94vfP9+fRlPu7HQG7uBselXZsI
7YavWlVJqUh+H1/dfvgR1ar8QYwUxeRcsSe8ijsHaNHlfeZqsvuyZg/OXXHMyOkk
UYyaPWMjHajEkg/Z+Uc8HP3wkydY8PizPpLKwtrp8h6a1zV0vgJts8gB/hR4zeET
zK/pjPi0vW1RueHmLUiJ9Z+WnofX9pk9IZCqtcBnQ1Spw1xWHypBJbxj5dC5762J
BlY/hrPyrguyojAGadRb2rwn/ETPQw4oNczq3jYU/di860N8Nv2XsAmnUiuhXXxJ
fd+tw7rMqacRzhcPdges8m+gz0ilqOmvv9PDlsWrEbkRONtzkqWo4ZQ0pkmpyF3U
v13XpYGePXsSgXeaRRT3uC/Mzr7pGcfg+7bFBnYw6C5WDne4nbxCqPd5jiXdjW0H
pXaLYrromlec0P6olr1BcBFC7lJe+2Ju2eh/CLejPYVvkDk07UIWSCJHmTiVxvKN
DY5BQ1Z8KdUMVzIvLE6Be6YnRuX+7pktp+Zoz6717BzVkvPxyYQh+9jaoidQkZed
HiphKuSxIQKob0B7ofQ5jiA0ALq44k9erlMPL7EzqlxXnIfzV9eDebFsEXVksbEM
yAJ9PfvsA6suOlZEh8YXWTO0HUhWVMWgeqMCM8O9ZruiDPxHz+wh9CCN67hpejIT
9p3b8gkCmkqKLnsEZuQWK2Sps9+gz4hkiF19r8sGZ/24AVVT2R0cjUcHfTEmOc8g
f/h4L5lPimt0OLGrk+kanGsuXPWyJhda2JRrIHm7W7dN/1Qa6y0KTMDjZsdr/z7B
IOUQahxrDUycSHg+PPRnBqDrrAZaHrMzVZsyWfJve0ntPpumD9WNrbM6a7XZd5E8
E2hP+IvuGh9lmQirVIlX8tZibADTTfIwwYjcWhtCgeQNHik+aBmxWbxLrNUYPYpN
53MKfYpI5MqdfFFsSqSkarOEV63d5jcak4ll9jhK+eAN0HvrBiXLe7+C38mjiul9
hwWSyzX200Q6ftvSbsrr4pW06dzuH2IXeLFrNTti63DyinRnVEo6VQcUVQlgTkmK
olXV+RmpFaUPFqsfzKjJoPMZygwF6wswM68F5OTWwhy1Bg2suVjlBkOtclUBqYU9
KWhCViQUE0KDxMotbCG14ilkVHCKkX/CCFibLSaj2sCI0+SvuD3tPy0hNhp6vWUO
utHiw/axS/zxnlEGWM4LgerKwmWsKKaY3o7TmfU3kK+opQdmnD7CIPu+AcWUg23v
fnaO2E0FGcoK3WVenfDKTcs2lt4b3eNk1qdI2BWKHpnIx51vD8rgphY/9QOCv6ob
pzUHoAnX+uforRbEkrvE5+zz2bgnSVFbd/j8fTakeextdkbfVWw9qCsbcfhwqQ2b
XIs4qujmgLuGYQkK966sGb6jaVgSsb8WjonCgJM0sxl51K/mhHcd1B80pVvCvlu5
Ez4BOLLVCxCiZnp0CmxnEf/dAYt0xlFuEinl3jM25Vlflp2G/2ruB4lTGyjwOLYi
yUtfMdWKUVtchKYg5Uucs2wA+SoRp4dQYfAL7k8v1HrTRtMwHvBdRpb4SJ1BLcgc
5xk5f9j3n/GRu0MSILHhcPqEho2SwdD5kEhJSR9BIzNkNMika3IUYdEMJoKL/bXp
18xVzCz2XL08mKhP859lT1AhZqd6SY7fcB7ECIvEjZ9HvDL5+MKgpNbGLukDV8gz
W0LIhOuqh9h5/M/gc9OEuq4FmDqp1MnKs6vjLZKDmdjp13n4o64oVuqWTi4Nh3aD
CvHt/lL4/gjyz6dRF7tN3SU0tnBMdCcIj2hwSqDqtABSSqeJmPjpm31T3DFqL3m/
SpMFXOc4vDgrOrS9zWZ+cmroX6e2AnHPebo0pV1cd4kXaHuDL5MnpsTS3C7nv0V+
ypE6z9h65mc4XPXReq31kdv1SfeSPNGg1sRjzj849C4CiZy/mICiy+odPyYWyrIC
ZqY3qreEOgFK/pr3TfO1zw1/KYhZMocqp0vjF8iwH3xG6VzSno3wPbA3j7JT+vrh
cGlT+GCDLxPLEzgxpXbq19RaxCBIcXWSKTrWujMmAdTqakKXqxG7ReUdGtbbLJoD
4Eq55WEMVNjPyfMY4oB8uee5By5S7SF0TbYsu7g2cXq15TeF5aDC6aK2r7nRhJGH
a/Pmw+Wdt//QC1lflQ/30SCDwdxDWeBC1aHYo2pq0lnjtG/6rkey/AiVEkroruN4
dC8PxsuIySyo9nF628UDGIVKGcTO+hymki7KiTWt0W97mZA4YgY8582aZwNsKRiL
WTg10pfYeIPM9ur3QQjjq4pEQ3DcGr/Lw3q1f5dmNG7it8BIyY2CRB7W5mjoubjy
m7L0GUoihU+7HLoJLFTxGOUvhagyDaxEa1ammnQUDl27ab0DkjeCdkq7cTJM1nRl
sx8TdlGcoDTghqZCZBGS+3Jfbbeoyn9gLt6qucopZpxEqd13yuEgx7OWKMXKn7Yf
K8zh/guN5xYOAbxM4kmTcyDsvAe4l9iuaMLJJ+GTobc/6Rx6W1OvnG/B97WniwK6
IdgQ2nb8V0WftZ/oeH785VkFPxvYp27g1pnBqmtEBEyQunudhIYw06I63pkf3zkN
sZ0lheVzGXtfZr2YNGhSt4CNAJwnpXXOjf9KsaZBNUX8QAkIn+WjFHFcsbltk+mK
ordjC8hBXuQf1c2MEzmvPx8KAwrL3vgjz69KrP2Udvc46j8fhbCDCi70UUlm0vMt
OqElCjOlY+TLQiNddZIOmUPBeDZVpfNcN/YWjyUCBZBCNKu3/RddTEo0AUGqqfxe
cuhTJ3wIy0rKCjFVMXZbWD96ZZCQ2j/hD4L0GLE8ZyCwg3xcqqLE1zVk6NPHhUAi
+rFRJ+gl8i0JViLWXMptDblk0/wsDVSkvHevLoxFhc6s6JWvFJQpnMnJGu8TYloE
DDjlpbrvJrzlzf/7ORq4TTUS+ZGnUVVKHw9viB6QTLoHooXCQdeUQx7gNEkXyc5q
1uYwvvT5g1RUco8en01y3WzqqLpoqmNsT5N5r6tm3rhvW5EwjdipX2MLLKBprqKv
JYVjIy+Pueu8PJZEJXyS26rxFWd67/Zu1LSrD2FYVrwgalDnWl6QtrW27tRaXeiJ
Nri+2W6kMAlZziDrIhEsadaEXYgzzmH9eoqjFSNZ5cUNB7dm4bcSJphwBLO3yaqC
yjXzx4ra9ilsQFuIY/DMSlvdLwD92VY/FY6/b/G6235JLDUKNVMzVbJ6CVgWhadB
nyR/Q3AE1W0OKqMLT56jNv9304yB/gJeve1dhfH7X89JS2k2RRgSa5Czv8iOMzpf
K6wZDjn+DJVbZ6iTcY/kqa1OZKIF5xYzEhMiEWFoB3p6gUxH16Ov+M5+vTcgvdxt
KpRJDe6xCt/XlGSPifHpoJC107qfQ9xlrBXgIpK2P6YzxBA0dye8i8fLfqWBiwOp
wUwh0qTR3vxMv2OBu2RsRLiH/cn4AT+gSB+2pScpfskvW/Ug4fOV08Mq+RemtIGk
fFFOlnMNuCRxjiFt6HCRS66Sgtc+IghASFOZ88aMeOx+wNPtVMtOKflRk+Z2l8RX
wthkgcn8U9gn9Yzkxl57bsenvRHAWOvXHEpBpYQTPIwsdo1Dr2nuJKk5phJobzwk
YtFAmRysZov2laUk0a+5op5GpKmZa4uaGtn4AGWI/+Zw68SBWYVg7bTbI3XdnFPn
jSXJ00A7tb212Ml3y6RQ39JI1NvNdQKyyYezkjrbSVBnUMLpFvwJWKs58fTFoKHH
mvpOT8WDc4yhag5ceQ04oueXZBj6rEcHJI3Bpo5e2CGLkLePT4NdVYb7J4fLiofk
+gz9regIOxABGckGRjRm9yabrxVKab8qWSdyeEqQW2bPbKib5AU1yAlka5sx2NLR
MPPauUgPpsVN73/2Gufy0bnZJMJKDk4s8jKjsanEitjkIbIvOhIPd9wYPTAB4/E8
Ocm9QXKVt96MiSH04IE4n7DNHaZLlD1F0abvwo8MBMGBHqwZON25tEOGGgqxw0yG
Wa+1EC6EzZbdV3+HiwZj+2WIE8wh3KVClrBV1HSbtnjMWX90/KxMQ2JA3nW0smM+
9i0sW4GHa18TR9YLJIH+oF6SViBggwMSBTwujjRUWTkIzFO5Eqx7JiF8WI0PORpn
VclmZv9oH1SKgl9is00hjwy95NwZpY1+G0S1zOMmwSFKapMRyRAVP0vQx+yfE8E8
scsVuNZf6vhxyGsdDKAZcGKzTIkoUIcPPI3/+Q/GFGSXZMwPuQrsmoG3Jk3ZcHR5
SiGd4tu8mA/NghmfFcUCvTBuDHPuIPEiZ/n9nEW28gCTePdGMmrh2YaeGA8WAdcA
qYGiyIaqHsLqknZJ7Twbp7/BF4CT65KTBUGXgGYLm96KoYpJNQAhjEUiOyVFtUK7
bBA1WEV3+fUjL398nkwgkds+PypRvwoBI8D4aZDsMMALxgI51Rs+k2aVsJ7r5Pbl
YvgDU5AGo2k+KBpJSfx5A6Rr1sRDlnWpygc3gTql0hq1ts9V+J6mF1xyFVOcvVxc
D71a0zE9yG3NY3oMxHsXW05TYjW5XzX8fBRCWqg8yEA5xLkKzEnN/0yGxptddVPh
8iz13k2uF58dsGVWTdEfH16dZTjLlj9zBxjt5Y3oRXjG9ZfnMhSitzSY+hjUaRgZ
B8R1djvCjPXlpKV176bT37NAoUhouPoTRMT8KW0ep3epLofVOWvyFaqYsNQcD7sq
ZExEIlHeAqAHHvqTe4bLsN1A97OsaiGfbZTKjmWRTg9ALCBE8YUYmwwSNX+UIvJO
sMiiaugMC+OAls1KcJ+5P5zdGDVdBDU06sdKuewX03UtigM03g78/KXq6PGir7OD
dCICwh/RDjxafI8YCkVQWFc3qJOBv+8m4JHDk9y4iW0Y03aZ7e1Hgu/lWaDDxn9y
3UhpWxT3HHeF+YOJxL9/qCV8RQ/H9OHTawZI8EPMx8tE0lGLUMnofBmBCWTIrqef
4Po9szzSYcbFfuJMOQ486EakWsT7Q8xFLCZ+1Zt5N7RgrVvn9478cwVaxHBZYj/H
B2jNo5CeelsddZ+iMwa7L+PfttVSz9yGEZTkcwxdbDs4o9vEZGgs158HtsH9PI2m
IepVMSOGSpN9WPxUX4yHhv5za5kbCHCB80nc2jzRupkoNV7izZZ80jcAsjXhNU6x
w7i9P1y4EFq9pdvsCcRRs18Mqvq5IBBYksXnMyP7rpOOG68UOEpOHTNrUij8TQ8m
bGpYiLd6Ec3cxpjSw8OFIlRyfP6KBYX32AB5pqwwes976rTnsAdcF5FgdZmkN1dh
O5iHfZPDtwGT1Ys1rik3h704Bctui7zAMey4mMMYj+qi3MkYhI3HMtTJr5qTsjGD
4yVIjCkI/6whdfjzcjXLcrBclPn7V5R4Z32fL5idSwHeKEFjAYj7xhnc1+zp9AaE
xUuLG+kS9fIR/AFK2Q5QxRUirP9B4QUfTF4xMas9A8vGamnH/Ptmqk1MRbAZMG/F
6oIEiIRD00Gw/bgPvJrk1SsEcqxtQAFw1Vvgo3XT18XaHhy1VbPleiW4GiLYmTAW
yNaiYI0jc+3Lf1nF4uVukeqpE8HxRKYHst+64nB0bTm6HtWrBuv9Op7YTu7PBShx
+m4CI1reWJCK9Co2PUweEIj4+As89AQl8M4z6kdEhOPnxvxsFXR9CHXSQgAEU6hu
mWr3Q2zr1LJ8vysfB34GkhVZn8BiEdfJ4Nc9PxXp+S4feGoElv6F9rC2y6uNpR7Q
RiwWPi/S/ImvG/zyf4HRWiXSygZnsKi+CXAO2XpBuOF7br6JNjMqqDKKRR1WLXY5
XjJsD8UCeDT9PfAuCV5K2XpTj3o0eTVktrH469yFBQppAZFPknbAFozan9wHkEZu
8OD7VHQNPIwqlUc5Ak5kT6M/I9ZSOwGGMEPkRNOxLPSmGHU5vye9sbDdRMG8Uns7
SdY+bJGcBChCdMG1uiMrmvnz04/Q2p6BHtSYw8Xmxd4VLFJH0KyeQLV4mAy3RyqR
6DEoPcz+J4S/UIU/FBvLGjT3C53DVsQkaceMRIptKYgvtAqyOS/hFYSa5hSisujY
W+sH7QqPVZBzrPbz6+9ECtq1XmgwHHxzWFwqmHMGIwK7BXIuoejRjwEGOkGGd1Vy
+kSnhCtHRvwrOglSOyDpcTiZRiPPrFY0MGlXwYFzmkJ1gW0FP93b39uq9yDfWFF6
0QCtpLz0QYqII3znUcgZPx00SVTILfPcNlpyclordnjL6DKWPOF0w0Gw9Q30uBEK
dVFTZvMKfgD5pzZkTp+R3GWH5mz4uut8CYFfv4fZlFwdhNzxemm7SwWoUvKufJJ0
1Xa0jyPc2q5GLq4y4BnnJEhYjhJ9QZEMGSeKIu5aTdp/vv4abNdRM8XkxkfU7bwP
wN3myHaahD4ZgHbvh6/uf8DBOVh8AqIIMXDu4mp6g3T8VO9Y66uodCwlW7+kpXdM
/El4LMgifxQtqXuxzyHdv+KBVfPz5cP8uNNOLtFKBDQL7KJ292w8k6MzMJXXdtXH
+OFl0UYcNwq9hkDChkX3JoDWfKzYP0IONYh0juj7BGdQTP4ZQ2vUmKQ5BhnIjIb2
KwZIlcHYxcOSWlm0Xy3cK7UB20GmGrjwqa+GS6rYF5a+2OMxK7VB8Afd8a8wSIp1
zCtfAiApU0LvbFIVs6tskroB4nynRIDPtCJ/THy6b9yM/sAQDD6csYAM60VwrF/Z
xppZJykWdsMXmw7mzTgPviQgsCI+7mds7CCCwpk1cMJclSaJt9yG3T+9C5kILoIW
S07HKPfZk644+VAqT4AxLKs8bmY9eSWjrSCKa3GgpjH7Dn6MEgPOh7RhMyc0GeHv
IuOtBMUlDoDU1rynwbW0C3NkkFbkERrLjYXnxg1lvFtCHJQgjslQNGflg4PuqxHv
u+PwNP5au6tj/SdVQVnY2qhlTRDJ/+UWzaT6zT3FH7vcrO0pxJ4bvzNhF0t7nFzS
reYu3wGCUhRHqucOMJ3KKpABiUVe+F78tloCE6jl4Dp+UvUb8eSNRQrfTl/KxrNZ
zE1GhHVI3S+ObWTk2ffN4KqXUUd1BDNCpJhXsYI6NgIGgJ61LYBO9GfUIZCaOkV7
lCDe+TbXyoHfuPpwVRYX83hoR7zMlzmxKrEmjNOLgfA7kTWAt5Xmu0CVWHylBAxq
eQ8YXGY+IxuhyK4Ku+rJBivCcptvFArkwXeWKfzrzqcW9zCp7vO1jNNU9wMbDGA4
M9TveM3bGjplWEHy2HMsfVIt/ZeXD3DfsTdHWNAafzZM2VfkTm/BVixPp3r/lf2K
KztqX5/r+BLlZKhgvKhsDiZ3toMSrjTh1d+7baOD4NbHYb7fOKu/pMXTlrffMzvm
0vvfnEdw6t+94hIGH6q7cZ5/JTPbe+mINVl2RUMoC4Qlh91JF5FWXL/zaZ7craq4
fgRE0ztd2WqEuFn7mS9C1AbR1lkLCAJLViTrQEnCByW9CHI1m9EAp9FJfNxnZJwb
kMSjAvDJ2vTxcAs6S5ndP5kbhh4WoCRuRR2lC+HJdSZ5L7UPOtvFHjiS+f9UuWOA
+NX17zpTnm0H2XYrePQ2HKbaePzGRqHS99d8yvsgYQu1orMV8/8Y2deEN80aaLgD
YopNc9sQ4HxfHfn/n+nY6rwpqV+4gSkIVYFmZRjis/sbqvmFPNHz+KDWce6JJCJd
IhYdEerKQ1ecc9QslEcWgkTG3D/HZnRbQk18o2o2pmSghrHLD/IZsYshsatEbESQ
E7pog5sVZ4uzm6vPTistqLpB/FI5ejkyc1dlwwhrGCXfePeasV92Bp9XcWbdD9eg
vr2430vpZs35azSRr8tSh8G2MMv0bJiZVTPuV+38nSolk8/2CGQutBzvR/lvvF47
g7TQulCPI8x5vkqw9t6gPKOXp5EHE2Lw6L3LiPn67bBjLh9NLw0s82LQBrV1O+Nb
bRojrAXh80c9LTVjfmyRUMSexc2TW3PMaRePApc3QNbHY72AtmCTCpOny6VTRPAv
PXXXfvvfjX/MSI7InbQzzvZ2RMPyMbgmkrX6AmskmF8VI1oB1tWWONEXD+8nuOSC
esqT0ilkGKmxc0VtYKRppVctpX/ZBztbrGPaDsSO9QopqfTB9wIlqKa+bfbGdWeX
zoJjz8tlciJFoLYgcn0i+eYO8SMkEVT+3U/LgdywxLkXqW0bOJjUzg/HZ1koo2AR
R1afScEVF258VcARrm0ng1YQlwhXx+7uNYupsK/SWUQ/zGhRX2kjUmzQZMnNsA+G
ImRXx5doouUzaAtD4tXAgp8DlBEdS4yvRmOmwlKp2fpXZYPCHGjtcF5gwHEmK3lN
GKaXbH5UuHZE1nL3LEhWw3w1kj+XS1pBK1On5SCpspaZUsWBvRFtuXkymJgY+CDm
zJOtovb34Dw+DhIz9LfWJmyux5CopF8S44E1+rvGXwd3TsSSpGOT61IsGB/RbaVJ
91CklndZPBZFGVcwLuOkcbLJLJm774WzQ1yJdllZ+/uhV3zVrKFTcSpFCRPew8A8
rOIjhW0cihmOZYUT74LxfjtMjU5akGaFLPLmr9eio8moZ11nR85zfIm0YVhjTMyA
Uy+79t9GgVcDUucP24AHoxZs6XUqARMuOZnQMMYbdY3+5qYdgM86dj1RWqB3bLFH
6JRXMXdQmbUVhCDjnUkYcESK2olFhDeuVo6LBdkeF1vN0SLI7vRl/cRGEhuvnyy8
BYumHrPVpMVTQIU/Q5DGDykmst6G070OUGLjoer9aEdugevoQM/mtmfGsIP30Wqm
7GPqUMDtEBGL6EqZ/W2VayQkJxNFezjzLe0Aox7nH0M4BHqmZlR1TCM4E23IzTur
6smZ9uVwA/xZ1AZVtHV/CksfJ8mxlGZWUoZR2rnUth41Rk/gyMfKMFlRtkinD79Z
gvhVsyfprL9qsTu/CYWwAMpVjwJ3x+KcihMRylppql0=
`pragma protect end_protected
