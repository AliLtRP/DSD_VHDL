// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:39:17 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Txofz30wYq7DTF/e956HYrK+BkbmL0CVVSgmUAKk+q2t3hJXEMlAq4qLKCF3tHff
2X9T2RLngxwlsz3i63BCLZ1FB0kydoC1CptvNYmLRzGl+JuqRDG0+7u4nnkIIV3E
rBnGU7lvQLgBx0bucHMEOvray5oKJdm+zwzyPzZaNR4=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 8592)
EobCgoKS9bWuD6LhtAzZEdH/S2E0tS9mE/HhED5ESjmlsoPl5s3wjMVsNNBRWeJ5
mOO9gd4TT4WYaVUA4OCTOjV3XPfL1iGhwNdK2N5jIj93uwl7be2FVZG8VBeCUlRV
IneZ0RvdNHFKITkrWozZAXJOHn0f5bX/5ngZzMx2cAlJ3urmvS5KdJL/T1RM3j/0
Np/b/Hcdc0W+htbOFUpXHazuvFIr+bjRSN8YO8ARTKRm3/XPPIlyxbLJLBf3DIxH
uJKV4PBigRGBCr2ZV0OG0mgLkQhWpf4yRwyUXcvnpcl4Qj9gAkKuVm3jQd/bqvph
8jHn7GWHyifImZmMe3bFvTKdYdrPWh6BoGSI93M80/QJYZuRpsILIkT8/HOguMZ2
FrjLr/MpqUascDBtxtbfgZ8TwtOnwlgzcVq++UAlDhFJUMUrcF/8Jp+UqOHqN2hb
b06UhzPpdY56TaBd5cEf0rx4XgtNP2I6xe9UBQM37XsmuY6a2yu2m5LAHRJbGajf
DTEoMEB9GP7SrfLN575amHYDUp3G5yR6fifirs5ve1NOSygPv8nu7CgIHXnYd787
qd2wUNf6NHv2e02dbg/IVSh7hNLFck+I6SVYwGOU8eB1cVd56zUNetorY76ejoDI
EpiPo4nJdth6lmWSQwbR2iiyRCuMRX71U5IOl1/ggGz9J2yQNMiNCgLgVZf0mgJF
b1lwIzvJJfCXCDH3lzsItIhQD6a62PvJnQamjIIpDbUsddHo/TcZuXrJoWFS04Jc
iLJzovYIxbPbIeHl2TRAwNWu6fK1qU6t+ttcDQrBNcEZP80Kq+rYzkbBX6HCrpPa
gF3hwGelBZ1VZojQz/qbgOX9i7Z6LFyiIeyCdoM+Vvo8sprzD6YM3DxRNkS/eWpk
q84RYiu3shylNk5WX6PXCcAzRk9VjAlYfP58sRl70XMgJUeqQCm/q4qc6LYOfErM
a6TJLgto4IRcjrOdAOI8YON9yOpC7bJBG5pOAVOGbnyRWhTq+jBVAvCXKqQEBvga
Gq+j1TyNcBDrDZvLfarWhpAb12eeDP2MQjjzpbpnGkV7JlcOtqfNE8MAoJz2dbjZ
nF5Yn7pQd8tnAu/GGLSIpJFcQpntkKkpKHuGu/ju1Q6eFfMhTwvtZjGx5BFn1pk9
fTm2AH6hHLjHfJeK7zc5psGLDVR5BGAniIBIQz2KYZmg+RxNvj4a1GpS0B/YRGRN
+UYxPu8pbMYBshGrBgTOmCVXpNxklZh/DAlNtsxC6oDxLpWA45v1xj/tp4iM7w0h
8oAuwy2/JV7S2GQYPBebsu6bQd3aOzaxejTvE01q26Yc2xiHsgpXlU7O3T2MXoE3
vRtkRfpfYbpgh+Ld2mizUvQ9L98xNslhRz7+B1kM64YT53RIBDRTswmkcWb/7Y7Y
CFPAKykaEJCdadVr6g6IVr3uehAhT9//GYEqr6wtUn51dF8KAKDajzLNEe/SB/pm
YjHZ3uv6ouhmlWmGIL4QAmTd5UVIGvDR6eFOYlHmSLwd5geLF1Yp97mlMsR6KMbg
0c6i2P+bUagDCzcgouN4ZJ2l6WV2I8pbA5P4ttcu99R9njt3MuZ5wqQLnpnk4JPA
UVzEO21Osqu5Pi22qx+XSOvE6ZLdhLGd3UTFcGixYJ/1Zq4iQ5+QqJLr65n1fEAF
hIsScNfD51ZjOsQcJ5tSOh8MUSJSZL+g2HSz/EqPxxcPhI3GSlvjQGTtHrT+zDTU
4Nglj6ytEH7YNJtQX//iqJD85R3Hrbf3UE85YweQRIibXr2XWwPxbyiUSjTeE/0B
rHO21Wuwo6Tm0ShPH9wq4qpBBj4qH77ERbLgb21HN5JKgcVM2IkkjPw9cmLf3ycq
nDBxINeIPatjJUFX4RixFTBfLc9PgBsOWTaMFLOwZD9P3dGWhTK/1lwahhUGJ951
irFvrUC8mS7FuU99ybjFrmdiefd9tFX3t9DiTqFk+LuxWkYWNPDmKaHxVMOqdcJ8
OrYueYJ/RwP6lChFQ78GiI4o0kNr6lIkmEMliuSqKjSOUjzqWdTK4dn4eqveG8wi
KGyxGW1SfxGcEBtIikiToEaGeiaQqntuDmaAiJKR7m1Ml2JnTh2UvbD/BVjwG/2U
Dx2lnLl7drVKcakTew6irVFMxo/iNR1fA3eH+rVouCtZaR4KuV5NEnYEsUI2Aa1I
vijxOaUNpLA1UEqnc/1zVwoskfcXpJEyYOLfeh7i8BZHqzbGxAOxQxeijZBVXeW1
vZ73mvYsIVTg/++OJXC6vaNCoz5WWM9+wHNxSnsvikSwisjTzIuwz8J9UV9FnN7G
NYC4MJwQtn4Q5NKtBsyBdq0Ux3esoXC4as/Z1WztpQJZbheWSMbaXec3/s6262d1
x7zH8MFQBouPIVzP1gNgcrP+vISIbMtCgZy2XNJFN9eg6kweU4L+G5G0YE43S4w4
EZPCo1rAY77QDwr5WO6vqLOPNQY6EIwQm5YZATZkurhy5qGgLMdVx4ueZuSyBgZk
tYKeWUS5H6JIJQo8kycP6kMTUMumJPFnnn9ywXRE6cJH0EiKbLN1QklUjLaiaViT
8KUWkog4z7APZV66OVaG5oGCi3R2aLUMs+N1bjvVf+NDqR5F/F3tpZPeGmB1kwFo
8O9Gw/LPhlNnoE8gx5hLwJk8jj7p/Ja6+UcHntJk0sEIkOo7q5QMEB9rTm5kQrDu
5IPkzwDevc1J5giuPRJn9wasYtOtZ99LYpJWpCqPWs5q/gWPmihEvH0P2McIGlM+
BzNbB6LBaziJY923lZm3spNeAfB0nIs2Nydsqpp/FDrSfA2h0IW9lo/lrS/JyVz7
qAUHm6reckR086PEXZgFPgFJbIv/pds9RU4/KyvQzG6lZQLTIVW0MMAALT3ybHUq
yiHo5XyzvBxIir01Uz1nCOOEVS++ZvGTqjgw7mIru3pqOSoCB7/EM5ZNOQSi4zJN
u0M/n8wRqQ41tpDIxq1cO8CS6XWO02J0Dap7AsbrjTKqqspIysn/YbCsxzYS44ic
IbCBEkI3hPAkh63RmCDRmMsTbsCWY8xVs+5EQYylfm2ZnaohquQgYThZhdPxThg7
tNB9Cm5bsT3RtBFdubH0yedAGpSVZ785EGs1hmxAtGmpWjGbjAE48aDewlu4arID
cq3wepXxTnWCa727MXt0c+WH6Lr39leVVMxm2Lmdx1ypShJzlt0OZfuUU5TTGosG
tQGZMcDaaD94FgLYAOPy3hI0vcSSKj+y3oRt5BQVF2Rf77u4CLMb7Y7sn0TPPMhI
nAHmTxIYFCvP7iNfd+o42Hz5wB9/fwJsbGHRr+HluTaagAbMwgGGAKUnPm9X/1S+
4h+2JjDKiSAb/yMIZlgaAzSOQFPCOBJ/XfOcvt5DZfWTkvIo+c+j6RlpdhpeiqQc
sXOGyoB2B2B2kyfOeE+Dn/csMeIH5GXh39d/YWTEcHfRC882yT+UuKHVAapQAGNA
3RXa7SRc3iGAmo69hFfIcnSwWnuvNRezegvSHzkzYhzn/DpSN7cic5WQL5TB7U5L
DisoI/gmMj+Nz+ROohrkqWhHo3Enxv4opfBWz9M+vSOV3F5YDMokEiUde0k7ur4L
AoEMnFDNWBhGtqinkPR7j+5dLEHtYBqPdOfbXDjtbaamNUY24/fyo+3FflkcUyi8
7vbEapydT1mA/UGqgoocHQgpAg+D+77uu5YzwARpUjfqgcj9jptN5ivHNaaaSQZI
onc0H5BuqCQ5XMSXvRP0aZJSkpLQ8u3bftgUDZJ6Hwv2d0MvcFTo9JAAayYEav4J
tBAJn5rSfXh9+Yrn/ODtNPiN3enAcTFyM9rq3kqDeWoJu/izdXHNmqt3Aa9ioyZt
XMAgCs52JYafqPlboXtuOHva11aWONLwY7gF3iUoYLT4a/vkt1z7EmpA8uhdtczT
raSgaUeZWqQ59OEI602ybEWa4eATze16iqpD4BAqJxnQzgSGsXwRipDx0loHd4gm
QTiWU55R6K3SnGz8g7BH5f6oFYC4k3EK62v7Zaco6DiRJb6io5to9SEzsWnuLcfL
9JZu6O7lXd7wXl6oLY2xfBH7FX5Bn1Ygsy489gTFhUizfuM1GRKYPMLpczAUwpB7
u1ghUDX0AnJXLrdlIGg37ErAVIxJ4ysQUj1ZZTwf6N1TwVkXsTT05f+NzrN727wC
EtspprLGgSp+q0ZIvIa/CGkUFEpfc676FD7kK8q1uy0ViJnAOzCZhF1TLEGlDIeq
k6lKfu7JzkTZF+3TfmpDvhC7aSQAI+Q1wlc1qp3+npnyBtK15yJnNmUgtaQi8gT+
hUtmOH9MmKEfzirHJuHcBnuk3DV1V0Vuq3mrIeDgJP1eb18W6fwi9Jv5pG9TYmgG
+39suySM3BLYdBf0j8b4kMtslEVSQSSoiPMvO6STRafG1VVY2BcmQR1dziqHPX1b
INww78TAiJBaMkZPGeqyZKU3v6rFyKyBhuslHiyoNcsVHrVhqR2Ijlo0YLzzOF3V
tyFTiP42EbopQBRlVgyiHzk7Rt30kMgcb5nEwec4zOCCFL1QkhHIB6Hg+0ZMOKpW
ZIrXfSxZePPTVQK9wNuvln+qLgVSsPvApW3krInusVZzw8hMhLHCd/WWan+xZzx3
UhnhX7zKtKaPyHpN/nivQ2340geGFnkttFxZhu1BWwW5j3lR7Fan6yJWcTZ1pVwY
1fIdMTyRCRPnRNrLl0VPu4K6dkhNyrwFPpGIRxc9wkdSTlAmejMORujWHd2IxmNF
5X9PA7T/Ihl08Razzs43glNHbwJCOPtMunrLS+5Bcz+6vI4P/i/VAnLhmS5o2V4B
wvGimwjbsMVrjBLLbYcl4bfocxdgJ4yMNXhgqnMRnaUVBtxV54xmyc1K1Y0QFiT+
RIVYnW6crQDobe0v6eYAoA/FYsjpCKo02EcoBOF4dI9nlsEzJ3Zhvl7MoPdboIPv
XAK7eY/IiK17V9IXDSmCSooEhn/YGtqebX5zORXYGYbasX6Tp/dm7isOZXd502NA
hWbnIcmTKz7vA3AeylDgTXqzkzMJRR2qgvB2UD1f9rZKIOiJ4c9cgJqQI0c65r5S
KOFohwM14vIk/sXdyTh5SdxxCCQ5PrGQvbVC3L8EneXWD0IEIouj+4Y/Hp3Yd6cI
WL5oGxxlFbFuhbevrZx8n+Y4cXexm+bbuRH5dDVJYAIv98iSLzNSKsiGz3mtdAUU
QptsT6mavr9oOXKBGSo6izH9z+SHK+MfhLO9Lx/ks80k/poge3KQO2AfatYE3XJC
Xc/sQMq1MUVmPFzX9uc1t18Be7EVLgI1491nmr3kgp1714uhBtgtONlnSQSGj7ci
cwn4VrJrTPG1/Z+UqCLmuny8HaDZcIZkQgTQ2safusXHFjcr+zIQ9M1zPDwkSt2R
m+ZZJ2yXhLfuFIGQ+K5ctonQ3HNczg2F8CpAywKVbin3ZURKO4A3CL35oEDq+lh8
kt20rn6IHbmNj2Ad3+4RhEX5Htgs67rluXM/Z0FvHXmkHshGtl5EBtSgYa0hikV2
5Qp0Vt3PxgYoAqUqo9opOKwK8/r0a7axpQFqlPdyUVdho15MSg9kQLgmy7fAVk2p
MIHJIutHvYAjx7jrAuQTQWMgwdoOSnkq/VUTZKqXw6LpcY1KZzOgo7IRudm12Q7H
4gPKbO8VJIVPCUpBdfmW0LZUp5OmIMrsQ1khyUMjApE2Gh9AquKmmMMsKv+8Tu4O
9LqdvITxUVaeSbFwurv+AeIsFJ4K2JalIdbJW/Z6p7omGAYr5BZXsn4Bsu+7cTeP
Ee7zBb4zc/guaDApb1d2dSeZyavIrNKkA61tTJMRBlchZV4EMq2bApG317C2PKkY
p1nyicTE4jkb3Iy+i3aV/O9plTrSALKnfLrK6H9FelHbuO+06D9Kh+H4jXnB7tIw
2VxXcVoTT84eYeN5P10Xnz1ER5nQPtq9ySAig/ORvCgBoeENeAzygprVN4S6cx9q
auAOu1Ow7ivmuehtjmWKeQsVF5JhA1htaYG5vNKEWlNRahTBm8Bruz+ZO8cM1lt8
uMc+GaqfIhYIpBz1SFaarb521cVBnOIX1QBc+IpZp2X5lGTPes6gdcSdlwlIAEaV
punv6AyB/vGxTe8OrI64xtFjUysUcaA4jTVDMa01WRcqX1I1Vb7MQqEhvxAfHslQ
HtooVSk2zClU1TeOz/bPHOuQgSzgSU8votCEY1Og/q0OclUohk3PNsnW7De1fue/
EYk7NgSGS0aoaDB7vcIrEeuBiTMKh7hWA3dBfDycpRHjpMx3lLjvpjy9fDkZqWfi
E6lbpH6GfixORoG7+qIaFHghT5lVPUxX5SZyXaD2L4uz8x7PxAqK4uapPfXhDYek
ClqitQH8PQkyn7KerFri48kuKCZePgQQZ9nSF9dJYN3ntKOCOv0HUVQYFXnv35I7
nYvrdg+cY08HbOtSTfH2WyRE8D7vHRXgMKSdZZxCM5VIkjDNU1mhnmdr6p811jjR
Bd8scXbFPeogkbat6tcZiCzH8oyZOSUfPHKIP4QRNtM/kmxLsX4tcXW748wGRcQG
MEiVkR43wuu4WLxycVjHQDPwmXXNQJ7PKg+OZeUR/UOw1QkuL2UIGSLWka1mlEMI
y/Fgb3s02cx9ArBjTKSlRQlCJt9UK71XfbaaePBDJf7SmbfG7TuDv8AP/ZZvwKZv
TAQ82qT4ejLc0CzUsNWdx1zc4aYeYcRtWBWO+IiuH7G7WoPWAH90oNtgC4YRsVQp
M9YU0FzsyMJb+Rbj9AZDjDkQPXko9szOPUSoWnnm2064EztvqoNIZ0aBdzg0kfU4
rf7y+rRZzecI6uOZQfET7pEhqi1YIXf1WL8spdQeBAuDwNco6fPhXvmoubmrz9tu
SCblfjhwIt+Y+YimuX1WWY2+i+c5S2oa3xu7e+mPot9ACIkVZGYfsUyY7pyfB9mS
vrsSrGgHOfId18GBf/CKKK3MhqqwAfleS5euW6Bb14kAikr7D1zIYAWfXFPctK32
EXtM93TUs8NSofFNOCCI/1mUajSvKx4TI/aerkKu6ljOndrqcfG4Yc18phMPoWyJ
8+/t4uN/GC91kZVAtcVXn5VqEzudspqA5Cz8z5LPXJmLysXt88wHz9YtG/kpl/5e
F4TvZdZzw8IUnbIAM37XHMgmvCJaYhtqN7EXurOF3oqyhYQL8Z3eYXNgjdLrbnQI
Y2hcBlRzefpjSIoiBHJZRn9k1nNCFXezoSxxB80hzfikMNTwmzfn/y5ax6T1Rq9M
h/STx6hmvu0W+IVUOeQqtQuZbqmcYrxqHdQ6EZFeKieWDTxJNuJax8qVR/eNqf4V
vl4xxKfUTSSiom9vVgDPqPX3gxHQtTer0PpV3mKAMw0K+IHb1I6tsY5qcS0N7W9l
0fqhu0KVrjbI5mPcBYDZ6Xv80n2bThjBkyYGcpLkHrXnJ/H7EHq5MDx8Dur1Uljb
LJFbgSdbjZ1vvehVvcXBiwIepSCkv3o9mmOoAGljX7cW+gwDexEk5Up9GtfzN6eF
6hJO0yYwmvTNwShuAAm6VjH9/u5hQsPNsR8URPOrjCv2kmK6zolrV8kyRheIwoNN
EJC2pkomW+XQTlorHQzzSiFoOjf3KaryGEeRRGcinBqbX9pwNsv+WUxmblTqwuZj
NoCA2AUcBbk54ag88VTMg9xS/0B0DGJqMvWmJUUby4Ni22EyDzmyooMcH39Owfqb
pCrJBLtbkGeM2dR/Rk96HqdUXbuNRVZHalW+HYNCQ+3VZHZoBTpJXAvGt0pmFQoU
YfOzn6TFAEJWkx2KmMZp6MWpmi2+DF0f59y41Yypb5Sf9KTx2TCE3DPJAp7Y+9/n
tr6xpJx75r6FtTMFRtgzdaMIHDCnm7TR+0gHVxaKpHW5gB3D6jr3uqKlp2zGOfVN
uxPJtbxs0BXjcmf/bcaesQaGm8nC22Yc4akWdUjew//llskVyM3QfFlfUzKBmxah
YjHmTUaltE5RP/Qsfkgb36tF4+dhK+/jBWlAXyR4QbConGki1taP47oFc/B+xbRM
Imu3JnAq8tZZdHR4SuqEOLPk3M/rax195fY1SdcV6RzqgGpDPI1/ULhS2uqVHRQl
aeIQEvKZwMwa0o+QJeDHb6KGAqI10+RYLRkbRshqM79yJ92jyzMqZyICM2267USP
IQnlRCqoSPdrh4zK+f6cDp9hfr2xQsJdhgiMJxf0DyzR0GZb7BGn37HmLZUHLZS+
hQP73NrVjnlUlcuyrmmEhZiBlOWODpZNqnZeYIq3ytqXY1+I4mxPRHZl+VhHf0Gd
CERu4Vo9daSVF1CTry0/hLAZF738sii5EVPf1nBl3UuP2WRg/fReBCQGhqFyvbBu
223ZPfh200fzr5OiMbtBbHd4V2KlMx+DSGfcIRZ5FSVCv8/gfEJpGxQqEdMjQTPf
I4LxSuICNxdkquPHfsaAwustgoEVnJdQ3Pya7SnGrkgXZGedZP64kczp/WJbWcrN
Y7SS5kTa1fG8N/ueasBpsbQzKkay86Ib6faIlqdse77jxszWUe24L9l4/laBVgMD
vY7JPMd8iJ3jVrhggMafvxCjQi2Vjf2CB9vewHey+HeV4LgGU+yZ4t3L3SBZ3vRv
Agy9Bqg9bNzE8RCU68kY9p/ThkznK2omEou/cidC//g27QFH5Cm6E/u/HhidooqH
xRtAZkju5bWvHsu4jmkgiE70H5tT/zQRh8sBHL2bFH5PwvKz0VyzkJKWnuYCDj2U
mt0F6X2L1wAJEtnpMg5ae+ImjA56SPUTXPjM8pgm7juRiMBGRJsyhsa/Wh5Mg89+
ce/inyKiKYygUza3giGmkQ1H7uLY0v3zXrSVQoNFCNJVJi/04L2x8VhXIGVZIqC+
cKPkWJ7Ls6uzdGRmr/28UnHDeTOFzqOVEfK+ahhIdon9EPrxLpAtj2LRbw68EG4R
OdosvdcYLTbnJlRKUtCWcIiArPWmSoGxvHni83NMMgwDVoEONLNohBzRgXxr6nT8
TrATl+qfPtZFJFElhipxDDGrgzt68S8DKcrQ/zBDnhTn8Zv0EgRw73tHT7JZwMGP
xOtw/r3Gj4CubnyJQbGnilyEhAjKnjBVIT1ENRsiCU9QScSMF0VAuxpEyttdI0mB
7Suv+VZ8RFqr0cbcWNIAcxIzcEESJt36Qf9XKyZdKwFf2PpRpKcVuJhUilNfRcyH
FYd7LN3rCWobmKj/BWh7Y639sSswZxLUbtnmlKd+hjck4LjZBVxxiThg8WLZag1I
UQmDY7g2v3fVcfwGECFBLAqRCDgweH4+dYroHQdjZ3UUvjurD2MN1uKhK2fCJmrJ
AREX6ELYJrvBfz338KkJmGrNX4rMbWYhKJ9shNo7y5sXdwPvtLQNQLmW887CAVe3
8Sd7GTBlxKmFq/H7VYcIUtr21gRGRIImxwdxYDktCU/CiHx8IUpfj/HtkDytdVDG
h7Puzucs06aIlLpnmn4ZjBqbgXOTtGt5+tuGQNlH91AcxdIncW2moS5auja6w8Kv
FTwyFxcpQdOCk5t1oJp+LgYk8AyCSVsIS8vIsFRcp/pyTuVR5/x+nV6wtfs3tl6o
xEt45aTD4E7IZaxN8inDKus2bOmNOQGTKMALsAIRw1tfcj/ZZe5QlISiD9kNtRGl
WYR+pyx01Nz8vVDNbbHnf1gP9xbSbKF4VfSb3z4dCbTNEnPe+qygAXRY7fq+Wgw7
7yPk85pykmR8Kt3J3u7y1UdTIcMgUXu1ZZSCSWAdtX8JNrLvQ6aGFbiHBBiLeIx+
wH17hGJj02BCAn/viMrEeXCTiZKU4DdH5nwmu31E9F4F0PqeZC4aAb76/xC+rljG
4ae4ivunvS8hkqat/gLGO+UKKwEYchyoqHt078S40PgDxhQXPK2hQx27zsz0E5Lh
kPrdicIaey8RbrLv3Lu3m/jpt4CygSwuIdYRcrzxHuhoqNVjszUntuhJLOc4NoLG
Y+g0ats/4vd54empzaXxmDbHzWw6Oz1UQrLbP8HrQiA5w7/dquO8x1ScEajBStd0
0/RtaavIX+vsRAC5nYxpHU6jdLElFiYc2aqO82RlOS82uwEmR2bfwgH6ID/7Qp6m
cnVMj0hRn5Ks950KpVpOSQ0gUjlhSx7zJWoMtigPdGgMJPpohw1ujQ3I66ZoJkeQ
zCYJoXrDhqAys8LX+s8XK3agy3CLvQ5w8f+0Ey4CNt+7aTwQ9t0kFM4y+SnOpsYk
PBAxGhfpBSLOO6vmquP69xNp7roUH+GniIvPjcQZEaUdcu0/6HmN7ZeMMS+WM44t
3zPmRZ4berdLQVww3MloVgsj0ouoDo8ntF1Xx8vM5+QDoye6Lsp+5NRfx7URuJFr
5iiAePDcAjGBf1m7wf2g1n3IiSPjx8FlzwDlC0BDXhKEycjWgLtxzDm3CF4yMLA6
+LhS8p6j4+/NoU6+uTEF2CRGe7HxJRqOD7xtWq5CGoROGOjuVDm2x6Zy9u0V5dlS
LtVGbuFAjpNjtzFvD5KH8RNI0ayIQU6rVP7crsqIamuB6+594jl5orOvEWXte0AN
A5s5iccG1qyz5/Hfuxtfv5mgdrgX1S0bwdA5eqks5VDihUIAv1J7xWsssQ/Oflid
+x6KdE+nH+mzlta/QZYEU6QkF5+e8BAec0DTK7qDKQi6RL9ozfwVgOz/1MSLn24r
8CbH2jfIJ2jXgAXg0IMXx/e3y2KN0mLWRdi2KATtRXuuttd+rJBu8TKNiDfe1d9L
FLxKq1kXH4/jmx+CcBAAvflYOf3epkJFXc1/KYCMfWvq4jfAp1+ZIIJCJ0gR8o+E
GSa0sN0oEuq6oEU7l3FxzZWUr4+G6nudjG7fjrPIUsUZbt1o9KOcaNWZ05yn3esk
F/JU8j+yV5CZ7sik5DLJ0DpMixPelab/mMFFON2WQv7I1G10dWVaVZs/i0O06Vr3
WcOAt7VH4t+NHghD4s+m38b6MUWVzx7LNanx19PN/lMy2416IpMpB83XmCDyL4dC
iqjqh704tKY1ZKRwbVpBf9vJnYjP6vT4bDHcMAzE1eNYoLm1ENH68YQx09/7EXy8
GlNcQvh1KmVyhoVMf6WzGaZm8qF6zz9+/Ffn7jaYcHOVt4cMzBYac0/OE8KErNcJ
+5gWtI02cJhcUGLbtf5WgE1psR+4a+X0+5msOuk10nCZPuD2LYhS1x3mdjuk0NRJ
FSH33DG59kU91z+ufFh6q5wN7EWGK1En9Q+HWc8xTibgTXzvmp3dexp3VJicuEXe
Zxm9i27mijEEDZagGwUx6ZV7kYuV1jWY2gTVuC09j8tm1e8GzmzYoAVvQmBMh9ge
VvwZY2ErSHrYGkddHZ5mwcAxbzBjhGhDzX8p06j9hRRGZKca2V8JuysnKhm56PuD
JsflPdl4WrfaYbmEZjQM8nQD2CxXneqIFWsWe3tsb2+9bl0aC6fUd92aqSVInX6D
/OkULnVob+4wdYj2ZNJX07tr4wVeTnlRXSGA+NZjCjV1ZsaTbG7aS9j/dgS5KYVi
`pragma protect end_protected
