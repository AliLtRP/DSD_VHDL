// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:35:39 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
QGGxMwS9jNhpHIQJBV0lqiUyDlcnnxONAxcC9AIrmLDZbOxs9xbL9Zr0CbcQaakx
+gx5yQ7kgplQzVVb9U7Bws3Pqx5rJwN8y3M+3SAyxpz6tTkulg/B5NJjbrzYzAgk
C0B7Rhj2Vbs7J1svzkE95Sq9BwCu8fE57i76EfzzzuY=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 10960)
uCkWB+GojRfQXNRWoFG5hlaPJpXz9Kz1ZeILcQfUbUiB6MVirCzccL1bwdw7nJDy
5Jnip7bQTupdbcvXFwxpdO1xbSDPUTNnlz++ZBua9GZ2DWuvHu+xXN96oCvMUNYw
XE/U6b8tEsjgoTzdLMoOH2h8/4xQN/+rZBlizrOsCkmWB0Wo11vuljRSyT4/wEVp
+H9W8PeMQiOFpNjlSWuss3CLJcsm7ygvhEBvwIQPs8R7XWhzwELt2PCLYQDkkQPl
FE8h4daRkTkJJozgdmPx2A9222D0UoIngFDnLN8h0bBpCRGBesCM8H783Nhfh99x
mKaCnkyv5/M8m5gSeE4DNRTh6/G+e63nezlbGTg2l0cl43CkIfppbci6e9vVVf8e
KWIwGJR2aewpzAE0a6LEaomj0hIz3f/+cY57kvPHKO5s0Cr6NXqjkuv2SiDLnYpu
V1sqgVdsLacK72deZGPsqenR7oBdHXRXYD8o0/nMCDBIu+7t4669RxWaK1rmyiU9
MZSM4Elw2BGN19zVra0632f7PSN+hn/y9iXVVJPGM1p5HI8ky/7QvD2QlWo7DzKr
R5zpzS07k6qSF6FZbB17jl2OR972eSPmfPbyy6iwIZfh3EE3X4wNIeMqc3mNZ4bR
xXXQ5ii6viDeVw3r2INW3bp26BjFUT6gw7AOIsoChVoUHk6sPRz4EHWwVRz9kk3P
OHYb4endlI+rz8Au+LbqohIM1jZ52AZeXcTw5Sy/cVa3viIgGGcToDS7b1azIRDE
84XL1U4ZyLs4LLJY8SrqZSmHKWt+7WjkiMm3vNfaMqshkX1QQePifNVHJwkCNYOp
Rr/rAqo1PpdGRboRn7BZRUBzz0OrXD8pS1Yk6rzKiubgOQeu3cv0bhbPqxVYzJrb
TEfFFd87Kd7LPg/z4uCgm3vYXlppJriVK5bXdAyhfaS1lCGRoxNI2TEwqg4EZj0g
P9XdjA0bY7KLPDIv1WnBJ8rr7B8MfosInXcyPKr9IgdBQ5EdPenCWNVLsQ0mQvvK
w+RgcXkBcYc6+Cryn3jYq1h459tIaZH04QLhNCCC1wed76qlg8wp5yFRtaA7Ijf3
XVFTwNowv9HIP8NfeOrQvdE23aZrMugwnADFCoM/riOisgpIfBcS0bKb5XmQY+3L
oDuKEbD16LfvkioBp/89FQGBOPNLaT1yRHg1W6GrEPXaMLwaBzsFVM+zpc7dubry
InJsLNmuuHYNZI+i/GYUyDH2hUjEg+TrWZVqiUdfQH8lVV7u+9vURbi8F2fE27fJ
wclfbFxsLO+kugiyx+1tUEaVtPJ6pFSuy108V07Flk33fVyB0TxKY3jwKMYpQBte
viBEKOLPwQK076s4vEE4ahHUZX7kqBYKv6PtJcN2BJ3cPGsAcELEixpdSb7ncpnJ
gzcGUByh69T9D6PXk3KxTzZ2MQc4YQMpbwzgN63EN/31TAWQBW7i2VZvMJS6VGbu
iHeiiXjMGzLgrCzhymaXknSRxYoJHhx8iuk5wvgY07njSbJ3NlOWV4sexMUJAc96
jQu5R4r4XFSj3E/VxLUfpW6hlTwtXWy1E+K5k3jQee/FcRsQYisA0qx3v6sODaZY
qrvyOHFG1oNDV5VcRGQ1FocALaZdhJMvpzIs8O9gN7zCOO8hFUJFe5j0m8L1HzKQ
6/3UQCOdmUniCPFRhhIXRArFJ5+t4Rm0KVXHE3jXsD34lRHNbK8x+NEqo8Ms/ulp
D947pfmguB1qXW1BPDkqTIF6SEfpBDBJDpyBC1+h9HgVBELAojNw3MDgCmlRymds
PLr2fscvX0sH3pNtD0rrAr/R8qre7YsjyzGY+fP4tZKHavkZ621jCSxjYQQkJuOu
kS5H1t9xdqmtAwuCu5M8If8Jignj81FmHI2mjcnx1KEVWCSVAWtbN9qBafs2FxSb
PePXF+yCYrVTkSb471HufuoWHgcqsDYf0BUyLGR8fRC8rYxYRBMzD0BpLgiHBTzM
rTZsZV+jjxvvrvO9cNqXQMx3bBPCf6S3QLr9x2ATkiOxzyX3SeroXswjN/noPcPF
mJwQ1MqdVlvYsoKNj7J5SCnxRqlcEkwk4T4bj4TXutMqpzmh5PuDqjMgz3Ir6cI3
u27b5mIcXFxuNXwx3JIGPlBnwjh1fNSWChLRChT00eK+oXoHXKXYUmI+WIf/fmYQ
xfaRu2rLOLnsdoyVlpbuJXk1QsY0TO3tXb5Jx3d2AjZHgDgHcwfp693xvZhfibKv
+fk52O6Hbw/8yL+RqtS6eoG9Fnz0xNwWj9EvpgZlFWH5cFObQrMzZRYqLL0FJSy/
1hWXOYi5DlDkw0RsBWmeKQwZJylbJOulp/0Oy1H70q45ZPpvy+E4KCZELalqIn8s
S3QexZaXBr+Okx1J6QnqPvjwE1HL0W8Vo/ajM//tnGyNCH8YYA5bU4xiPU46r2+P
u2Fd1LDzZEq2Q4WuHoMYPx1D2XDg9hz2TV7GPCcJCu66rbpCKR2urO8I+Saef0X6
0VXKEgq4n5XtHZtfTR4gb+FksCvSbvOnbIcEcOW7NcskD89r3jEs2qr5oixFAAxu
UNg8gF04da5LHz3rXwsldaSDRC4bHYHWN2nOhBp5NqtVka4EpmEc5HvwguifDHY+
CkLgOPS4Rm7R30FhgyyHw0xFei+7IV/oSUJJhAQAUI67zmZ1A5NoUu2IUeTpeJhP
cs6g7phG2Qe3OHYgHZ2qkWTC8AjVxso0UfschMBSox/VOuW7UcQuaKlcYS/w2AwY
0ntbY5Ehs0fEtl7SgnInYLvReek4JoLSOwUX40wDEWZcz/P0pANXPDw+UGlgJdDO
I7vvc57LcB090lMHNeTjlTM6di0zdandpxRvbHcon9ULkHwfxHybqpwJFyjaA5Q1
w7+6LSXiQYJeHvKBe3Z92MZdJIyhpUIUXGtU2ZX8R0X7rlmuyHGjXPpTnKAuNJ96
BJc6Z18waYi8MlXzJ2S6MxX6uhyLvg79CsVfGsPKrBLRvrQFS+p8UeoGyHET/Xpn
+qLzxUpShg/6PefhIGeKdY1ePFrYQjkF4G70mN3rhiYjpKc6oPBs6MkRqXSstyTK
zAij7UMvALyKJtwrKAcLNsEFEjEShfLhWqB1haFoOBC0wdmLupSJRpCtGV6FhjXz
21rLVA80SkR73H4v9CTQyqshlgxvvlyFmbFu9WEG400zJBAUf/cqHpI75ucu2Z8i
y51G4CVKJmirus/bbp2Xdh5Kzzh+AACftgoIG/B5mdLSo/cjHKTwpK2m9Xlq3eKY
qo/NmAMZncn/n0sHJGYgUgKsDlygoFglUE1TVYovAo6f0pSEhTUVcr/cZiRyFae2
gwxzjQgLqcg8tJHRcPnyrdtoIxOsEc2Nq2aKrkfZ0AMDAoCRj0nqCfjO+2SnAY31
2/6SCCyEW8t98f+dF2JjtOk+jiSxaMMu3y1ULhpBVSY8Rync+RwyVeeJcoIwBko+
4felOd3o5Ez8Ns5oEbanQz1WLiclFspYgHss/v0hymKDlMmWGQddyOot4dWZflwc
ATwyYG40rtlj11u5h1xxKz+FTz4CPjxJBiHAl4pLPKVM+LWlUbWzJ5ArWCItfZ0h
t5L+0jDD2ygrZHnqiADyUvfGSDdFeBmCpGs7Nwp8eZCa0jGvbcPyRYMlDotUoT1t
seTEdxMAzRCDmuxvpnBtzQFqBwTtumoio8iKwYSjA4qG9nTZVC200MEH7kPLGpZ6
mObuhxpQtBb/By8+LEBcy3S0f0UBxxRtOPH2kCqihz9zmEGF1jsQCysPsqnSsBFR
wLOOWa5Sde6aTleXFYr676wLYhTJ3hK4mzqAtU5P7TeXSQzpZEDMwS5VVxQG8YzH
0xsswsVLCmwRW+gOg8UkvFLsPt3/lNn7eKPkp6ZtKRzLjiqaOT9vFVJ9kPWu/5Xv
nKL1PBvw3saQBc/2qqgI95y54HK/hlBw/0sRRwCKGYu6sHiQNWIJTZTaC1COrJRg
ADd+OlHT7d7gg+CILMCHAqnzoXO6vauGQNAY2qKHTdyNUP5FZK7GLynUFarGwu4A
8t2VXaXY6Ir8Q2iibp+AOwPN5qKULCcRq3H1jwtFFvlflZ86HtR9r7MfYItrJEVO
P/an3RXtpKNm4hBJlrGAXqFR655xlegyrhEVmAPMundCvtEzLUqPkSeuitRlL2Un
BC1ydvF93cn0aQERsDjiKERh4JrOJt38Mj9bzJf+glEBws1zquU1gGUWAfqxjtxe
KTE/XGsApbM2iRDP/kyJNjj/d4AJU9zxzA/ZVeUQUE16s399zlV8tqxt6220pYpJ
SSXnt2P9fP7awsVWwRle5SL8eryx64+SN6nG4SlJ/moe/2/gbeGdS/XrEIPm83Es
LllChdCSav0nkJQGxglX26VD8UCCp3LN+VXR9j23mcpC0mHXEm4ET92ADToKlvKP
Tqn0zXgAo7wGwup0JgHf1j9P1Dbkztwoz8/JkOdqI82lfQKVnDAlvwtmkLCGjiVD
O8qDo0hQApoKR5OWWJlj0i1pe7GP/HtzB4/rBKR8LhfDBU0ER/PxtkoTKbSxSMHq
V2zLqhjYOkP1fAsQE3PxePpYGAp6Xq5fh7IGJT458uf5lxwQDClAxLHUVfLGHU6k
84Ik/advwq36lHzVXBp4A3pmx8uEdr0VMOzmXd+iBg6/PpMQ7vR6BXSuwl8o7fFA
Fsrftqaqy7LMUt9iYVJo5aWPWuN8iH7O24yEjJhIRcXN5JqfTqJFzk+Kcujnqgvv
c2FoaHCFjc41nUXk6Z5Lt211yzdbrEOUNsEZbZmOfX/akwSBXbcZwxRDp2sgHElK
jsRq7SQO7WIul5IsOHee5ixZBYnIZHgRUDC4gtU5Q9wZp3gTOE2/Ib5HhXyewRvt
mnoQ6m9bSQSHQl+CqWTPKKccWpONc7zfgsI41pwe4FQyG14oV/9+gwmXcKIAUjrO
4n0h9JR/NuhESklLbzB+gwWkDg2AUJo90C9ISBO9oyoM31qJsIPVGGJpFqS37fBp
olOeqVpTtBbAWpx/zFg4SofaZGtcLyAGykGtXbqqEgldLF9jU7JRiwiFtnF0ykhh
VVeV9+ucVy3yu2D2dx+me6OtcdLcSqtxK+y4UtNHm7H9yPK8YfE1DwSkhOIQl+PZ
UPCuDyB447cn+QE6Zf2qar+stFANRZeyIdwQ6kMEEpXnquRyc0YDlmaTB6SKwjW1
FFFl9/Y3QqasD1VGU8SWL5Guja4bc272mFBWbj5S6+7HpDVHbPPx05Fk0ehHSiUZ
wnU2zrTpfrg+xft/khde2+ey8fPiXbAEzJ5YORs3SgBYrKlQgSN4uDhvoKhUbDk7
G+gHVgT4jI3NRsZvqOwNufiapE2LJq7TMuWo88wq/7YxeV6UmcpATtxnaQPxU88/
+fRnGLz30J3YUorxOIDrGwX3/+dXTYxlzulaY6Lm7auwnQNiyfP3ZIetBmEEbpo4
lfOxQQORRBQmN/86dxV1uj1cIcAGwhEmRPSByysJ7i51r8ff9/vzdJyZkbt02Ooz
wctxPXx+FAUhQbFIIQtPokZiLxBrVDJbHo4/vRaCjopgucvALNfSLvEWPHEH2cRe
+Cc3mLxTwhTBbi61wBVHqW1PKSmSWTdKVZAvCbYQOZYygY/yOgWN647DLlwzK4gb
w73dqsPUI3pnCGXNbXHowr/A/raAgUSp9g6u7IheKRGPprA0WCmlSNaWjizzedrv
p6kyFoRCNx5deQntjHkGE8Jxb+YNPZ5n+Kq/LVNOFsBykCoUM9vFXWK7j8HSf+M4
ijuCV+Ok0SH1Za2/tNq8E9b0JpX/F+Ai2mgh9LuhKUPAq07nH8w+DUWHCpC47J/O
OTQeAbxp5FPWk0BCLdoJLwph+NWR8qWwaqJlSZIfHp+hrQl1x72l+MzohY8dKhQq
P43mVsLujWS0sGCBSUs0mt9Ugi1DofyIgz3IJzllSs8TXp9OFTwfEwjmMj8tSmHP
pWSpxHeVnYnVMXhdBHG+dL1zc8BjI8UBsAyUJADY2/C0sRoASRHdGXkUi6viqgxF
FMdzbvMkJCJF9EO6R0JzyFpzMHlRIuKbRbgTSk+81UBQbjcUvgOMCLDhgmPEbrKT
r9B5VIh8K5nxc9LRXRJfZopKQsvbdx7+R/duG5wSRt/5+wWJ4xTQSGKE1RdgzQ1D
0C95T5jo37oTvcM5g16lEZueQ0GxOsSkJgp26qOyqyR3jQb0mcyWwQsbYIWpCfE+
pJ3ME0/QcrNoVhjqg5fxOC8LzOvNVSeVYyCmudZdW8mU5620/21kGqPB1ss23VkK
nnO4uL6zgHydM/ZjCD5Q19Ir9sYP0EGobuK4iCMCWwdpT9equ+cLIuhqaboc6xE8
zwRMlroQOjSy7MAknzALc+y9rGImnEXSIFpwYjvOducp1w8jr/haqSsx7ux+YEi4
1HRI+j/q6cGexkzbDbn0nZ7X/be/0xix5MDh2Uj3mj925bVJSFRyVdat7ykOvxC3
unKiTd+UO6PWn6OE6XrKKEg9UF9FELS0ZESdgrackjYwXxV4YBr+Fc9NPu9jMMi0
xCam3LOQ4MAFTYZwmenYh8wvmQmP8gfojLt1E+FantU7KdP5mViK9ONuFdWEEVyP
zhQJwQDh6BoMPXqEbtDCJCNM445ha2TBkh7CCqAvDR/rRfUg0QPQFsi1RvA4Dc+I
4k9sd1Ue413trSB5sRi7bmAi9/a6RVmRebbQdF/uAjEzLpX2qaKb0GW+HEMmCZfY
Cd0t97SQLWMk3r70yYcBKM8GaR5NFtVsEhpjADXHB2CD6eeGggWMBQrMh1V0S1We
9LwwWoD6rsMHiz+V+a09+H7jAW7BmSKCrcxn8Odhy2ghwO862NpUYLQ5qyyOvmtt
+ok40p7AkQM5koFqOuoRI9S7cXwYWBtqg+GIwFjfiN6iOLlI/bVFvnwO38SbJY1I
Az7VJNQdBsab4FA8hfaTyscETmLi65+ztRH/zbM7gTiInlqwSsYR+cZXyyEnn1Lr
wtJuRniVlCvUyw9TZ+vMXWkKYBgqm1mL0MwrDL12Rr2NkL/XhSE1PRtNJxtaFHcY
Ol18eShhod5QwFWgDRBRFKvHTstqju8gmM2l1C8SRALnYsi5ey0k5HxUuCEOQnWi
qb5KLMxMaj7+TI8tDy1M32Nct07bd5YfJyIQhjQ1TnanIZPwsRTfALRhGYjnM3u2
KdpUxBOHCrdqJ3ymJZ/3QEq9wewztTyHy+FBH0lC86fuO+easttzLkg4VbNsvwgk
yy4DSvbfLocpzX55HGlXFumrmqWo1qjMW7oFohGFzJfnN4q0HoIkodIwLwgiPN3F
9Wdse1e714+hVo3hRDfCyQFUzk1jSBQfLxx9M3fRPEQ80nmbTOHCEYPusMVvu6lu
p4SqP7q6MlZR8Gl289H/6Riv/tX7G6cV3WZph9oOrN8F3O+O45H83xI8JHoHWBLk
KFGgy8EREnKwB5xDFp9W+SppO0wcfUxYfg+5Mg9UJwsLcqjAQaFOOfqpOEPWtN0a
JwyFFRM84zRi5XXZiSxDnmlhz/zbKhHLdY2By9JATNsYx7Pq99xlfzEU+ng0gTzl
J4CWQzTVkCUF9XGTYEKTxVeCKQkX6Ec/Dtt8Vz7h6OBLDB1Sm1hH+zw2kQ4F1GUL
wccdDOOxOJ7YthuHctAovRC8IRdJMtRjJADEKBoXXT3f7zV7YEy1Wm+s5w+9fw+H
VN7csu3lDi8AnqoZb8XA5oLue9Ut1CZ1fddt1omo5zeXf2Wm5sXJ86kQ7wsLbg5y
UQkQEzjIxdQfwB/gnBewQt/Fhn8etHpuRXZ5fvQih3iF+40N5mSFfsuqqvGay8a6
96YlFLtN66bch1qWyUzxkN3shfax43TiTDzcMjNh2a+V0/kkNulAK5hNRziVDXPz
TGvzdTe82DpxjSkKwVuX2KDwWVQITdc/rNQajgakaYuhvrmlRRYUGbixFJG+AaqJ
2fWsiHJF6vWOlONV+lPbPPc/C/yZ32+e9UHzYzNoVpyb/f+r2I9pxuy8azeGovuf
awdfQqpTTwlB2sQoLVVoUgxfBfYrR73yjCL3PP971dxX27UAGjqXjgxff56+Tq9D
n5DmJlioA486LUCpVcePQUNLOBHrPoDojSvkyxkHzlVsgxSY3o5gwYQnQ263Ng2J
qZ0gVuY+VtyArxrrTOddocQI5fafXySO50aiy0dYJ69umwdDf0/k3crh7Fr+1u7M
UoOKq9OhvjlPt9qKE4cZg56WNA4GEwIxVNoiFkOap+Hi6Iz6SCgiwFNUfpSmenIh
Gs6zQ2v7Qqw/uT8lJBF/HoreAtQ91uJmpp7TjZ4N+vy9bLj8HZWVM5rTctr9XImN
10GW4skUxFQmsKkOXoOnWNwIW24OOAhS8zdWYy9L0hg26HOduMDJnKL54Mo850kx
UpiLDP5SLLgsTKE95B+5ZwZQtne7pamQKLvIxolouODwa//tKeyIStGcQFx+Nz6B
jeAwI8zTS1CplE0MqqMdNTRVYtYtQcFkgZibZ0dAv3t94a804/gbsMtb/cOztMKy
/tGGEA5PdL1x9bufPUBT9+90dz/TbMzAGE0VgI5f4JkuXn4YPybgXYDrdwiBcb1k
2PZPnf2wZHJS6S32TwD/jQ6sHrDzNXpItL+Qx0UXQYyUlIlv5ytKeEFb5PXmSgDX
ijDADBJj8Dg30fwrO6rwZ/cFMmn9ZBn3H5u2XcLK6tZoqQRgfdGurO2VNEisuV42
QWcBHADKm58CGkvWHsyIQXKGUiYhhTAgCSnmf110ePUQvLm/cGECiJwS52vl8NLj
JcuKbK+ERLjCfkv/T9eH+2elwl52TQXtZveNx+JDC6tQrAjAFRECb7gDdy43x4v3
V1vY2UsWrY8YfhPN/XzMX8kPyLinrVUc5N0M5bKzekIqKjN0oGOuMfOpL+9qbrn4
ak0PsLjQEJOB6AVwmL/F0Y57vE41SKVyzq8/8rq5F9BPYmvkL+khQXGmRlVdH7CN
nVoXGEwIcUh+8JCrd8UKT+ixXUEPu2bd1JwuxbxUQr35Szed7C309monf03rbEl2
NTeyzAw/aGmNKY/uAesA/0/z3EZe39UByf2f42/GhlTbTJg3M2xaGoVdky56IsLT
ZT0+fvSamWZXQPPDZkgyIC/v6FfKjAcDO8igAxttx9p9QQZKfnzBkcFt5fn3+QcH
LtOMcTAH+hXNPUXlPo2emQcsNmco09/6brwNkNNZj8iZ8xcc386/rxhRndnfhGOl
TD0NDOxcsmx5xvNQ0kQqDYXcw/VcfkipD6mzqVae4jYpS7tY2sykZ5rwHmSxso4T
oiE+5LAroQ5hniBVi85XMUMZvbUX/vdIPgkCaDU6QVHVQGnELp+zFDic2O2Tb6LI
H9NnSwRq8HajeTQlnAeYAkXk22AG0jYN3/IF206mHiN9CGaVZzF9UpEI4BadOKMn
YU4+0mlXcDw3MbJSTG+MdzZjHi+L7a08YeJFpCm8TT4J+HitMVAmmWv4itPTft3V
4G+cD/FGlU4WKY8vFTiG1bxSfRkQkrVEXPdOk2x9celTa6XEITeTIqacqcH/tRDM
2ZFMblbHUeDryH+QpNiQz1qjnYSoMd1BmthHRE1IAzANACUtj4bqSLnulkdzMTks
gdurGWFhnYfXc932ZPBhCR2rALarHeOhxMkyx55REB7hxnBLzt27CZ0x0ylDGplL
LqTNegANdZun7SeeBgyiY/UA+BzR9ZvzWeSwiERShUeIGdhuKg/m6Bg5NrcpFZZ4
UAIEEVfXlNty7cujkWHW6MdAGYCPp3cW/q6BF0bEa3+VKtvwmtdaW/W+YjDktYmG
vFPAnr9Nfb5uzQEfibnGV/jxhKBsnc39P2xhAOkF4DPg8SFP3uO4Fu87MemPhQTa
l3+1fPwn0jB7Hb1doTDdc7i+PCIyEDjzI9KNXqTpg6Zr3tiLms/n0PKskTqDJtXj
kzh42yJncHclK9M/gB2VdGbt+73RiF17+AjPeYIMD8UbzN4m1KBmt9IBEIy6XZHE
U5rozFqAcYRfXE+Iwr8ogoh+mq3//+nkOIBJXpLn9sSaDFPOV1va3Jpo2tJum70W
n0Vq8EFIWqtdus8BQS7Xx/LOx56bQFhVCoKqSS7THyeE1d0i4bxPdnxMjdjAYIkx
3ufF/mTAoBLCNwSt7zpZIjcJ0CVFuZd08Fk7xQuCIT1bsDn8vV/eGPdKAkO8NuL+
KoSm3HUwLyemiLBzn6upV8J01AGezb40/luizhICwyMr1K6AE3Bm8CWLIMupQfe0
74+MntZ3/MD55sbMMR69Tfpvg27rmsqEfuxMZ36K+0yCRUXxuIjDti8EioXpfpI6
CpKhrjBvRl5qbbpDlxNccgS+vCmEwJUdceIn+7PgIdozQrjFuR4+xcwqvVIdp54R
jjtDnazKkqa1NqiPtwalBr+In82o4eyTJHox0nnF7zIBtv2HLdIxvws2MVIQC28L
bJ1o36X7RW/VDF3qDWfxp6h6brqiaSTcJCMNa5460BnclJYsCq2WSIKK28ZpXs03
uJK8vZhFGWyAn7fDZRljmVR+R8P4MnX3Ga4IzgpptpTSMebl3uBq0IWtCJ7igawK
3uuVaNMAXVXIVaA1jdfaohArPidzwOTpFHBZOIMiaRapfb5f5kAeqjqSmZJueNqR
7PN29kNYBzUlvxjNYeKqDZULj5X3Aa1M24k9BbE0BTfTZ5nrDLMyGwh21m75p3BZ
LfhIJ0AXFNPLQTDGGTRuRmLSbD0TsZvONqn5blhjs+uiHTMbeYpThRFOzYuZz6aX
p7XY/9Xy3hPT0qXtWkkXzmAZmxB7U+e3vY65ZwJ030PTyL1WucY534CWwvMuPoxc
sizPlSFX4axZYn+NNwjiZiIghPkYvrOH5kRF8hZHETJ99fshWX/FMSa8IKyt8Sve
kEkd0NcuVvfmIPn0KABuez0M+kXLES/ax7UgmBUI8mIqSlz7xnJWKc4ZHtp3rwen
yRw9rzfSJ3phBPuxouAxNOyp4ptEd9lKJtQnvHMmo1jnYKgOKAtOTKK8VODL8mdT
JvzNBdvSo/RmdFSm1dqQXXaYLQNsDXzp1584QeqzvUWWI28NiU+6/++r2MGdRuZk
PjW231zJk2mSJUBWLOzF/wKouLyITT/Ap3Z5TM2RE0POoFAJ4NiiojwiEAeV97+u
ISr+mrAvU3IeqXZr7jqpJ8LeCvcPagblD1M7yVhpVd+kfPVs3amNWrtnSzAV4QyX
xdcz8qXZnNW9lbAv3ve5oAeg8Q2PLIpRIESKos5IzT610gPxQZi5S1WM7xOIS0ZF
138jKV0XPLYSsQJsjjzLmLldZUickA/+F32dwrZYAtDsl2okwK5GAaDIswa52gbo
92iq6pnxD9zbTpEaSya6f4VxIqueSAsp3MntxHtEJC5P9SIi/TfN+hDz+Qftru3q
ib9wGusj0Y2sk7m2zvD0BIG3CeenoOt5BFdKyU5EGAzTu343syB3GixW1VibmBnK
uG58kTGeMI3QlDcWRrqLhRBPiEoHPN02VmiqpN2+TLng/uOqQIXaWql3oph5NDVH
mTo0iNUM3nAD2aZbKAOSKmAO7GXdqFsTFuCxEYgvtEdSBL+oE0YtLjqE0tvghBL9
te2/9dKjZ3p9hbF0iVbxVzPxpFJZxaAxh0BKnARAFJuYXApaD1QFqDHAAsv7Phxs
GRPjCjssa3CJaBRuFTcL2kHxnwAQNicHNffkFbb+wDJXz08T6HwRPk33bW4EI6cJ
++L+L8mi6+mJgqJpEpjqStyr1nU1OF3rHUAKyeVcXKnpd1NrJ5UNKbgZPn0oIYv4
67zufKwne150DFT8YUs7VExBDgO0Q8Mi2SQM1GL/Yrpq8v3t5wd7cFKEAaAevgGP
snTB7B1rfX9LD8spkEt8UMFg96PfwLx0X2WtMaLy8/PSs5vu7eEKbLjFRl6De1Iw
OdATak0qZzs5XZoGb4D6BYvDj/rqqcg3+6tiblarW0IJU4WENhBeMe+6txyoxbp1
4MgogUS81NQUWNI4RvNp0PMua3CTqNVICXY0XcmoyKwJbQ2d4ASjHLLbgz2nh0SQ
p6OJCCHcICX2fPcSi7+TAGZ+Tl0C5bXP8kLDpySKbmZ8lCx0g6rZgNGyEW9Oo7pj
5KLZKU9p8hpriWVh8Bl6PYbvy2+uCh2r6npN04er1tAGfMX99v9jAO3vX/j2crLF
9A2Si9Kr07JaNTcWmAJpSqcg6Gwa5r6CjaTSwuUyb3WmO6JnByHEw7xlK9AFUO2s
wZo2oFeOd99L22DCLHfKH/EUnrbhrsl4JvuRYvipVFR0m9aTx+p0VbZz2rgKrIkS
7D11EtwYIW78GNBmKNjttj2DAPpcPiylfnK7vh/4UgKa3pOzQ335sRGBDIoqPjIP
gubX9dv8cDV/2vo2FQ6kniDft9L47V0tWcjU0F8AP34RAze8fdYTbHgYQslTbDel
i3gTGXwtce1gymxt+zj29ywdwSdDQpDBjy/4XGwFXNdc5ctZl7nM3CMhYZGPxY8V
HzbiqCHct9u1r4omXIUcaaYya78C63bECPdPKSErtBLBFxLVxmtIk5FOiyWSX5Jt
H8N3Ft+g7zzhQ0jpZaClwTg+csC5sSQkLYbdw3SfGqOP/ML57Skr7FzjZPpGgQZE
//siQ54OWF/EkiaZWFFzfwX/j8lzOizh0moIrVEXhg45psOjcjIbPfBnP2nyXWAa
gDf+76YvRcCFwWt+oAt/A5xZtPHsfe3rNr07Y7NEgQMsYdOQONWfyIC3rCfrCTfm
j84CTY5D490FwEAMVdXym9lIqH+fen2rwK+D1mQNkDkSPYUyUOmU+t+1j/LdEofY
nbS86o8wHbWMKMj2WgWfQQwKPb7H7u50HsmAKciAImyZ8K5sjgq+jyvid2BU5M6t
mOV0O8mN6+5f/+YMUveF7YhUkUcgUjrw2Qjp04mRKRzJoMCVYJlNG1kHex81+msX
EXHoerbKjAXzcUGMzOQX5rcFWqvYewVeRNkvEImrZlg0KkSO9D/y2rd14pVd7BFT
PxMTPU25b0iSXqidSyRoRTny5uh6RyqlnJW2egliaBWMDc8hLqnnwfOAupoDO+ZL
pDICTxXbNO+79rpiy/TnXMEz3E5PuYHgA8XHh8iFxw8kzqMdaV76Y3dPLgeo+KtJ
dm3Za8S83XHqWoj20n+ohHV60zcMKr/V8BKgiTEtR0dyqotupmsQo+ZiObZveec7
VCh/Efs9p2auDqw8GFgOM9AsmrrDi8CofCi7TyY4mRcrnBhPR7oGks0C5kqBAjLq
5PRAWm2s0nvWeUN7gQTQ+MRE12OQNFM4K1HDI1vAjAXafzuXFe3AYiuwEdzdjOWw
YVbw2O9UNd0ABA6dOJyqUq1bdbczGYGa5k4avVPNAdFSMtjVQs/WrrnyUiCOzRPA
Y9GGLPQbuuXnQWxyFk+qUwAeEVrv0YNK6rRyxWSVm2XJxnT34kVi6nxE4m5BB4Sk
LjtFYvgnGwxuxuDFEue5jwntlOZMVIczARA29bYdWci4WjupJyevg+lgGdpyPSjq
fhp7N+yX7JVkhHNz4UhrXSa4qMK4AJ2u3CikEciz75pPIrxIlRytPO3XGTb81lCj
phOL72yhO0MTALJEhD7fVVeWfLFfr4tJ9kN6ipBCYTS6iud0FjpSwAyntDHL2QMu
BzqitCdc1Zv6BdQOqAAtV/rzFh+8iAuz5mpCaSkA3GnuUj2erQb0R7mQ8uqAwCIX
gxPmToBzNbiZb0PuvzpmRfgwJEZStv8ZDg76IA76Q4PGuWZUQ6fyk/DLb83+t0L1
6UzYt/NufvYozsAmUYWk+D9ADLuG58moquws5+rx+f5e+awKx2i55otMpJaxMQaR
Rm/Lw37WkVrIMrlxM1N80suEiHAHG+3aws0rnrsmVZWPQkQuMuIUeVuIcMCiOSIB
CXBgKhBHr0IwCMtTGiLM7qCZN2FeHIjUGXiD127KeoRHL/w88YTF0lA9pqnnNu52
g9ZsdKKvb9l9PUJuxttCVCzfzJznKLn5p21M0486uOaEgZ/yl26iKeQKaH4WJzrH
NnoGrn5X5epO0FQ4/6xJup/SAb8xCOEfG9ecL4BFuzPAIqlofBLaZbR1i0IV3Tua
58dkNwK3Exjcv7MNkQ5Y8LT0rl3qiIxtYMcssQTrqW5kZAU0KWQ6RkjTg/lu4dWl
ExYFdKDmvXBleQGE1bJ49nn9gT/+MnrLMTegwsUZ1mJRALaPLIg4rAmCo/sMSHlB
12GQOk2olTGof9T6B+PJOqZ2LIod+Y3V8tzIa9xUVqV9E6FjRVyh5aoCoxuK8pLq
sf7k203eD3FmjBYEYdV4t50JIkfo7Y+iMyrBYsutpcobEIzjjoNnC0hyYWP4hD9K
NKAA/Hmg9q8Iiis4ha/z4XNSrh3drRYDsVNP5Iee8Ls/8jwlsd3wH2r7T3LotrFc
hqdbZV8bxpedwgSGXaoE04rhHOxhM97I9MQxAtfEQz9ZWm91MwQ7SRt27S9onMdz
S+iTCsP9HZhpHi7Gj+07DYL+oKtMJOw1HNU1LJ/sImTKsMJY2rh4R4CyNqHL3Xkg
7SQZIJn3XbhPrc7COMjvMok8gSQG0fDiIabxjvJT/btP2iaJmrPhryigw1cKofdA
Z6pejXkTqK2LsSHTL3uTyg==
`pragma protect end_protected
