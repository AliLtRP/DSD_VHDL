// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
rI/DHdQzOKiU+Ubr+awgblxauZfudgmq7tUppI5IEr4croWP0oA1Hm7AVxJ5m84QhO7dAopNC/ic
OKxc8XsHnwW3XJbIqTiIgargdswgPyOKHWMNyvzBYgY0blSIS8FaI+tvzRHn9ZHHIsw1o5MLwVZv
mpAbw1jc+TCn0VeZXtPnW77DTE6d1HJKn8194pAG+3BDKlIJd34TNoS15x/7meR2tyjaHYcM70EH
jt8oWl4nT7Ut5j+lE5r6J7AQ8CniAcpROGyP5trb0y9mOgKU9c9zIgEPtCpod1WpgZS+Ue0SXbhb
KhT6w8p0lYzsvJc3qZ7k57oaWCnCZ93AFRffOw==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
IDI35tfnxxJ9FaWR6D17Q9TmXS0Sg6SyQscRTpZN/FsR2AYuyfUMOc1/cBRVvUenjTonbnh45/Jq
lGe9xD2/dkyJdnLm6C4IpJTk52Rb1Cyfa6ZsJmu2gjUcZsVHBSvlllodYnxyN5ad2LMc7gIAqA4K
tr95aTO0ECZdFnO/T3vAtCaAN7fBlhnJjQ4SQ0DA99RVm1k6tVWmvgkQYWS3Gu4OkluLtJXqviuT
JZUKTQYN+HrBhE0GkII7aghdF2ttETjyuS9NNX2yoUKdkWH1DjWbP+12yQkw7K/4in1ivq7eeMcn
XdbWlMnbcK9XAm1aOwd/WeREguYrOHA4Y5q6tei0/wes8dZo+/mYgLksksUQp2+jYkqvErZ2eS6s
TEsaVTv57Cx8QgBzNktMZHzwMlcpnS9lk1cC0y2upgWGo8R050p4iqjj80swTQB5UhFzsMNghu0s
9AjM624CVz1sZ3iv7B0MCnT61zmiSItmHdTro3uDaHnuuxzx7xdlNGEFPNOeFgSqmmtAD51546go
Tjus1hKGlQhAzLtNj3/QL/PPhZuAtAuGUXDQKJCsAHO3lw/ED9w2bhPL1CykOaVqZYRc88y/ypVQ
UTtP0474gmutt905uLpCW6LyPw+M+UjRC5DCjX19ZKJoWreCndNd+qj0Vlm17rkvtd4rDIF5SfOB
B3J3dMs9j3+3nwUxzfrSxYghFotICxEb9776h2at0ejGjKafREU/+BP/F+7q8F2WKQrMVjK1w2Aw
U6Q5XBKVM0yfiYtFf+u385CRxTh84gjgwiXJ74fhssbQzNAcJeeS4huXxSAVr2pcJxu6qj4s2uYu
DN/pslFhn4nt2ujwWctabO4tkzn3Su3WYRK0UHK57quR/Em7BzjIciVaNJEc7sR2aLkvhYjEdAA8
zVEnjl/AdzyFSEjUpv72jyJBy07KXcBP1pYZn7oFrKT72M/8gVnq7Xz8EuO0xtOrqROfubnyE1xj
b5RNUB4eAbzR28AXXdOLb/Sj8rssDLrjbG0EwMB6wQOULVLtHuzyPobJP2Fhb/3jQpOnB9Hglghw
jlaHidk/Sy3wGPva42JhSs1I8KZ8v1dz2Jd5XxgkBxI04lgWpBCN8eMlPFK2kxrrf/FlPhxis0Ww
z4H5ZaeP9irUZXQLxb/oh75DhkyhENAGuL2X9vKNu/vSdDRMSD708VzbHRkq2FY9Vp9IxM+l0Ue5
6lfGJecRdEtPeVW5uio+JKBLDDSwX5Vyg51yvpVd6CTi3XgHFgnzyvOWzbYYWQYSrDuyPN8L9Vov
1P39J1K7f0gWvgezUq8rvoIC/nvnIF7t/vX3clj81/DT9Pl3v6h+2bfLhvCuGzL+vtX/iTDWxART
o8wV6nOJjkhwWyLQ05hQg5Zhn7NAk10udNedXsuwb6jrUsMNr60ObX/MRFNvS39YgZkjdYeFI1R4
TNU/izDjTKKysln0gr+yWucbXoVKAsfH5tzvvAdJTOqirlTTxq8/stoipHKWHw8330TwGAwFNm8O
aB+knZoUsVVK5L0VSYGS3oktCSYQgJTfTr23YfoI0bmwrU7bsbf+nBfE5qWbq8S53psjzhTZHQVA
yBW2ZcS8zzxk8lAlTBEkOKT3IsXlhszRhq0Fka+ZMrthzBSoK5guRtVv7+AuBJeIP+1PkbjLcN7A
jTmUko1RpXWH08uFdYloueAZxQkku2L5vBhwiHXR0S/hdjJHKwrGyoKQe6Gyz5VIaL7IEnQ5ex8z
VIMSCfTQBLU0HlDqnDKJsPj9XIyBrZfnIiMsWo/tgOLuag4uYTcMGvgLbnwr/8mNlxir2eaIcuzu
JKY+V6Vx3hOv4Niyy2TByfr7sZoxnC2Fh/cpOTL9GbdrNWaFYMDKAHD0Fu4EcyIqSORkkeQlCz/7
58qZSU+GB42LP0yMz83SfQ5T9MIJuIXhQyKRhNScaPqpjoWzP1fYNwMp2KS6K5INB2/1fRdsel6/
vyx67z/IalhEFcRS+Z05Xb/R+etKpOASD4eDvX5Nyx4mdpjNBxLrIQ3alOBX6J67Nx/Hr7sVqP5Q
vdvPB3bLWxcve78KrwQc0ixphTDtfVzfPVxujr5XTOdnmJKeRLOQVkJAHLUHx+1kNyvqaF+WASDJ
SJ12ddIUB1WTgAuAkRFc2IsG/BDlto6uHyrAuGUDH64dqzp9FLfGLNannRXLD5u05IMWMvjUy+HS
KF1jXZbplAaDIs1zuUZR4zL7VfvjMgHeDawWQedASmxAIkeW0eiNep0PX22X8ENKSMZQRGnl1ZnX
emd7CYWVcuWamDL0WJdHgLXeUamESsg8pTA7kB3eRVaw4tetvLRxGTPF1mwtnV3Kd/f3xG45AOWC
0LYVz/72msiuVIq66RPMKH479NhsJSC+PTJOnPII7dGvLSGZgaphjgJrrzxBwVuC+q8g+I1TD1sN
D517UwC7N7vifNFnYI6gTa0VmxnS0F8qDMqa2lY8LcowaNii7nh6A3E/QJheCZljSg1vM196ztJn
laL8daexg9Llnlr4QPOQd0VF/5+B47KO/wuW+X6nT+q8GOAgfFglfxHla5ILifnvPGA33mfWhVAy
9Zo0x0TOzPBuz6SZpZ6HiePYFlVZsm04RVykgvSfgsty7jjilyoij3U5YvaeB/AJv7oJiSNdqWeX
qisPwyHAFm35jwUe2sK8qfBpZSGhNnAsjR4jqHBitr1tvYREzJb5QTfwr73EaBzmOpphAntteaYq
8Tw91lygztJLk33XoahXCqs4CAjH1iF8IVUZaa7yAyQza9JVQkJFaLD/l5/c35wsvHskgIsZzVVd
QnsSsG7UkIy3I9BLSspK4/VmM8VhtmzoUJXBKOSb0egFriAn9nEyFWgwfHcCeb/zOtgQjtskhUiy
WGsXtr1IX4vA6iiUaJnCINeX2tM0k1i6hRFKeOV/KAFDUUpWu9F/SJ2v4l4knSDEtCHoMfBZ0vD6
N6G9b4bmVlJiu7asAzEsHTdzVkmQI1Wq5O0OYZlI5wHgF0VgHxAabU7N5lK5rJ0NmHDXrhk6SV77
1Kx9bixWVwpCDgnyitP7FOEtOshJKc8RnyNJKaQy9Ma0v+dxfBw+INXAYx1MMyEr0cfL9jNwD0Id
sx2XEpmRQyNV4U6F/vW326TeK8WsqfZ4gM+ZFu0pngjQ83+5x9V2oL8v6jb8+qfv2aYttNntMNd6
tLj9gTnPEmzxXU2KFQwCQ5VU1pAMsGWkPPiZ5FoBMKFNAW5s2ZtKQCrxxqLQUxTtrDSKURZ7amUM
bqaMyznrbHJ/C8/Nn1B+lfoBV2GR6VHVoHwJVnhDoDN5bJo6bKN/sGiBzkvFO8rEyRBRGDSpJGxG
Mu7oPpBh9iZnErxmIuMR0Y0sEx9t48pCrAWI2db8w0m7DrhF1W2Eus1GX5TztLyVzEOoPdNVTPWR
RPtEcfhhO4yc2x2taEpJL8aNFSCt4gZ9DNhfMGjOusEyVk/IqRpiK++3ZTY3Tk9NJjvlvQda1eKT
A21v2CzPqKTC1qISBPfXTwO5spDjEjr06d1CtSYs2HvEtrX5WDrlysAAECvfRNo+TOPgu85wEuEq
QK8gJptzC4CNlnaTVLLrGoXHrEq6ABqcYYTZvh4zKqdoFs9IM4KA/FBr4VFzXyMHXGZ7mEqEyKf3
tQrrUD9KdWTxX9MlY2u4IvQg+XoEA0dztX1+/LA7RFvbcASFjDNM8oOm0s+GDqsXvKE6io2b/+4z
qpOY9vDc1fRqzVQ49AC/KA+N9kPovp+V1K9IyicastMyuOSTe0s/vxZAYb/FqNyWM96how3bLaSZ
oCaWpBMB5XLxqHxLTtrNnl4cl+9sCcNP21Vydx/nu/dtqPT9PK3nzg3cD77u+a/cjM/ZtBzT5w0t
X8lb92x8gxXZKVB0V8z3Q70epmgJ1OYWOp4DqEAeYTk/yPw8OM8PpqVbhFAmPaowks5eHj5sacvZ
mhFH1FgBGxrMV0F3wVB6kIdRHomE6OERVkmlXUlSUkQlexCAgD0J9MJ4rokrm8AeubKGfh8dF4e9
ZwqrqvMPtRnvo12P1pjR8npt4Hkm7hrpMTBemC8GTZSaKL0w9WjlpHm/s1qmoT7EogGlEGCzBAZQ
TQ3hnFODUbnDNF7sQeNo3bf/kJh3nKFgp+CD242sqKxKDARAAjqntZvuHREy7mCtdbLScCCUIbpj
VS1fp2KG8hza2Q1xF8rzgtu2M6CIzkDOR5tYsN9nk6Y7+KVQo7CidBwsMXiu4SAkYaQ3xWfV37Al
dhCSMmL1pjABo2CAOoLRbXmkYw6oYtVAHjYbE+X+dlAQcnZn7Ml5242KzSp/lfOrqZgW6T2ewE44
XXz+YJSdqsVjizWw/LzSZyhgrrjdqfVx79KoAkPuGdMk8Ub/x09B/ZRhPEYHaD/tSGJVkVbagrXs
K58YauJL4HOKoBnYyarif8a60R5foLIKeor40TF+rNW7ns6CXP+i6Yh7Y0NHrk8O4EUws0AyAGEa
CNb0kO++kpCHFzdZb9VjP3BlUnXJwb4bg3Ny8La48MOIPE85MJ797IOrgaz9XheFUvi0Qr0MDg9u
Ehfi1lt5NwJwDFkyScOQEOizJ648NbGAns2w9M+1wj0Uw/BHFzKQZw7ggPCA9gg5i7kRwBSfoDfo
IZq3KFv6mce2uvcJ3KIGglH5s0wApQAsmDRW3e2M1iD52LZr9n4c5lXmWDPFhpYPQKT61DxK/7xN
ND2r/bHryZbZhHVBUOeK1okFVkgzRFUhpOoRdFmvy/KUUoQeK/zV5nqbCa5MvoMck+0Pu6k48gx/
qaV8Qt3qxzQX/SBtzu10S5AquGreb8wZRPR1UNQTj3dxP+BaEHW+FbQGPSc6crl/Dvpnvfw+2AkS
YpUvjatL3ganaL/rQMtIhH7lRQyUtul6SAfnoHDj+YdhcMRbK/cw3WC6cuZ2KXPNer9QV+6xdyXg
0M/dXIn9Ij8fARbt/ivDXuyZMSK9PPkmj2hw8HbMvEwfKTciNswkYypMITLs3fPAcqOAMzsqZXfL
2SNJku9P37ebrImw0R7KnyKtoT3I7pE8yylfvOPPGgzsAhyBHkdpELKHUhLm3nDAf4RFxMjIYBSc
kmb3wV4RB63l+Mrc4RnpSGvS9QMbROAy+b30YTdNrFdQMhoWnoizpRDgIiyW/SQzY5+jwAoXCbnc
6hCt2rplhMW8fBl3pxuOqK/9+yFLEr4JWg1tcnxPAaH2kslTj1sshWgHnf4LD2smP3LPD7bAcx0s
vSGLb++DWsmvHg/Py0p9UIU1Y9gwGfnPsTzqLyIDpF7u+lwud9YXKpU8NwC/nEUrUUfEiJmvaT40
0YPNhMCwPTN2AJ36Rt+rMN9UlHyYrcNpfU9LrsGsNwVUvdwv8Uhw6oQe4M994dB7HjTTtX/KwRUM
Uvs2b3Wl/uEbqomDqAFg+sPpMOHRAnsVFsVRwzOL332BgfVGhmn9BQG4emPX6NjIwrwpboIWsbMa
vNb+WnTOtS2nehIhd+aBnmyu1SDrgrVbVtNcEes5AKxBTT2U8UKqRfbHwUZCHw2kO0ap9WFDFcNt
JxckzRr0czLgv6vlOiDd/1C8frdMK3Devv7Xa9neIJ1PuNt7ahXPvufL5PjqN/wgT1pTWAZHatrP
xIu6rp+tWtwlkLVx7QEmLo9HumwTuPVDfomE4pyZp9UV72azkOL8MR8/14XjiZZ71OuK+kcPSM5C
fv6pZpCArWfQOr93bWIuOPotN/aQA/StpmI4StgriMaKfNZnEWB3XHHYCfp166fio/7xXtTIS+wu
/8/Z32pbXfXRQM9Y7ebbXL1VdaOrg+/ouFIlTOCOD4ZLGTZJypEMEbR3IHoMtf+wqAYCY905RNtW
Gf0qNVRRfNxxMjJGLykMjiTH+ZFmOCx66Q55DW1iRxW98OIMu5ahvkRgFJjfOZW2idYG4/k1MBqo
B4aGX+TcfPOO7jaGxapbjadP09I7zqSLyRsiL+TikuxE7yS0HTZiJwFL5NOcKovgCoG7943RyuSi
FWXShoDMTtk0UsEP2GgCIDScTyEhUPkD4imwIXxAdmbzi1E3NWVI8PUdIwnX4ra7RxKLAEoGqgwM
OsdK5rtdVNV5EyS9CyLg8kcOXcpp4fY97J7aAcpeIOS8l2AxOp77VyOQ9vCV9+KGBB+yAZZmlgmw
2kyB1k/l8WqEtno2wWKj/Ure8aj9MmvGEGv1+4YBvBpGYvKxUVR9iJ6Aa3nAfsEMiECGASKgGkYQ
h9yQYQRgLPruPbZs1CDLSxm7WJ4d1Jly83SuPPfK9IWw9fKyJ31JG8DYWBM4A57ewbwCu6gdKcek
Fe3rHSFqC6pkR/ProDSV3kymgQcWW6j5GgVHD6Dk5b3P1ovygrH9I+80Z+ZFqW2ZmDmEUI3TGUF3
VJSeilwb2k+dyyn7hnOkYeIMdxkMas1tTSWGhcbE0E9+jxq6Sb0wD3+rza+c6yehdZUZBaMtSRdQ
LE9hXlYOfZISjDhIWkPGCdpI9y7JRq7pFznRZogjDacIc37a9c1az9bcKkP2V89q0XZ1J2Y8qeg5
3OKKnhhXcOlaw+PoBxrw+kNjTcBq1QWw4wvY8lPq+YrT5jnrcuxB0YoQiPJzE8+5AgsQSE0DYoff
Mw1F5a3bdeFJexRWDKya0xh2mzc21eODn7KmJ1Sry3w1r9RG13Hq7tBD8vb2sutPixfKoqMpPNmu
y3Fmw6v/EaaBU1+4LV78JJKTuCKyFgePsZWmVGlu7rf/dXTKeAhIkx7AvwGt90TBpyEngEjL4qSk
wvrG49c+gYgOEMrLg9yeqdVA/V+muzJPs4pj0dt3t9fS7N/0QGhZGGXfk4ABvbSyECEY/PIbQwRZ
k/Zgh9umL1TcIDrfwEYvvNURtvsf4juWlEVpnxCuvZwe9myulEIV7pDT92PtPBeeRDEB4n+H6xOd
54aO+8iPOP4wMNawBouggO0C1wp4rG2ZgJkvjd6KN+SUXNCBKOnfL5trQ2ARmmWrJ3BJJmE0efzc
1FcmXwdTSvEyacST5bKbL6B9+roBdqAx+S6QbTbpOfufy4RiQVf6Rro5dv/IVC6E5KnXj+ELqFFF
hsRzS2gL/GcoU8wrG3wrkassX6aL2/+iPI7oy9a/yxB5X6AeVxorMQG5mYFtELzIGewpnzvnoZ6S
dOCTHoIAXAmcOkSOplTGBZHwqKGJZ/KZ3tg2DRaNFj3Fih2CNJkpIoogbo+lkQvgqkk9m/axDt8v
PWY/ccLdR42FSEVQ26KAF3ch4HPSUHb5r9qhfNDU0F6cMkAgOKkX7jo39vrPyqwTINJvm2qUF4bU
PLrY4H+pf5LppPypOaUfVPMGscj4S2D6Qw+pE/pwZ3qTkQl50fC7edTpkYlMVNaxsdlwL8fwe6mf
vrb17X+/n3DqF1klxKJnkiEIRR3QbFqfmj1W4/P3WHYml6t8wg0TKIEuRKiMRHoirA1PQFfrYYBI
LefwJj5FnERl1sgeLNFWx3nNfvmclGtzKGg8t8oONFCqBE5p8qNL3w3IK67Vdgk+HqDCuYIn5s9d
bAFOKbk7ROkw1pOD3/JO01BEeYb6SaVjDmsNm78rtoNjG0eimoUcR0yZN6dpGkW7hoZJYZCPN7hM
T4myMFt4AZi5n3X2vs2XP+R1NRUp38euyN3+aCfF29atLT8qzVjv+LVD3ExH34r9jIC4ecXxS9Eh
A6Qb3K6T/HqVhG74U+Q9L8m0nK6cdlp5ztRgAAndtmiapMGTZ5OKPVm5CaML5Qt64og16sSRnwQR
10ZTmDWu9iAVXBY+d4mFnNEb3913VHVRNWiJYQoFYuQbXbBvXMhdY5Co660nTKnwhbrkOuVAm3We
Uwz0JjMNYw23XR2GygtJ6J284/0Zz+0m+uAFz0EZ2SilZd1TW1zx5x3mnnxkTJ9TiMoIAz2mGMAE
7SiistHkE33TRjZlPRWDRIwYxASC63eAhEncv/ZmnMWpNIsyQCTa0iPY5UHyfSUDKWrEA2Uk/tcE
OccyzlwyI3C9Jr4sfE4pZb3yelHhjlEyZQqYll+i0Z9nxG4mwTOuPffz7it1fvzXFTlx1Q1wBw09
ffxZ5PDZrbRKQkOknTaE2HR49hct1d+OO7d7c+Np3y4z87ErgztL5UaFDzr1cqLyznpua5aKZiDU
yJEfUFYbcBQ4v+a6AH/4okJcpldvgHAYOs6NGrbMeGrwVTap1le11pfYXP7BJDzwOVZDz9I/OwBg
ZAfdUGVXkgQEgThk4VFOnlugqSx42aGTNuUkvgIsrDwnXi/2gznmU/yNhFCP5ol5LnEf9tfwn8Ta
e11IQAocZdJqWHnIEMRDVPDwiVoVyq52pnUnJPh2yDWD9VuVnI7ZXJTJaLeOT2OA12EK+hYTU6te
WcumPEzeJ14cxvv54NgC8brrZx3xacSkulwXtW2vpJvxWBxUysiFLTYJmebaQgnSHufGmtL0ao8G
H5DSMDZ9TvmHRqRAEXwMxE3M/VxxiY/vF+nt4j4gUNg8f6HyayR+BSyrqVAfBkBZqp9mJHZeveCb
55YnYNyPVjsvC0XPo603UWfcg9pO9qmQs+nrVf900arn+LQZbFwIGjte4EFVokaqQaff2tc1mYId
LCYjGxIAgMcbUePl6LgVRDsO1nIPi7ZS2AdI/h/fr60HoIuisY/R/iDHN9OTgiVlAFFOZO/OI+Ln
mHv+16hWLmDT5LhJiNSdYek/ao9aQQegkomzU2KSU6/5YPnDRnCBqVtECXDC1baAYLAoXR4tRMcj
n5I7yv576uGr0l1l+BnYhgLl+Wo2ibIFVB+Iu+xixSRJlpuAHd7XyDK0V195KEo9jRmuQ1TxDukb
ZKhbJZvxknOMNbhBuMY5H9s1xDZV5B+/EdhyouJ88LM517Y+lk2U+LglEjG/XjGn6ELF9eTJGEGD
0z9cFwPcewNvIIqHGxaWJ7GPlOeRhR9U6icRXKd4pqfXyihJEGBXh9KWR+7WqwdOFGYuK6ol4jNM
GSzSj5B8bDNkh4e+WKQqjqTicxw2yzjCX8pxatRsBxxBqJrRMXPTjxQRL7+8+B2vl3LxzuvLjbR/
4/61ZNNvtofwaSJHx7eIqek9Gf7sVKC0oktq2Po/aX8a34TDgVjH19s314mgZBPjzZajhZD3slhf
ep0A3wH7c3HGOsQNEERWeLBTvXnE5iMVm/AudvNUqZIlTdlP9c9u6tOaHppYFCr8pQsvWYbFKgRh
keQnnkJ6ZvAtMQ4LQ+Us5CITuRRVJw0OT88XMHm8peq6eaIjkEEE33F0hHeAQuhaBU7KvNP6mPa8
rX5uqzmiZBeZrgNixDCQjR4f+eXnhyDqM7Ho5EE6IhGb/EIJcHMwpcexsGhDmpEoHybdE1gNbQr6
ku5sboM0TCO1cwBQKdnCRjsMbWgHzKXSreRaSRmJq/ufSsWsdCGniM7B7Tt4Nx6XL0XDKer0kqm7
GLrYvLLrgbOWM4efNFYVgv0mMPpovs1/G8sItkxqBfibVnGF2bRMGNKm1oBIR11Zm/mZtNNPfh1x
qPOG6M5IDwM6vGUD16F5YwkXSWYL+t13UK3f1GV6hQccw7tyXs/0uM3LJibvm65+AGITdIV5H6pQ
Ic3+YA+o0oVxTGxdUp43punzJiuj9lMscKugq0e5F7eHAJRBD8TaBe/FHzgyO5hm2ENdMTLHCR0+
WpLMstydVOJ6wJyc9/An+lTPpinUVVqbkTJO64Sh23ao8rTQgwJ9j9IwezQgqNAQ+2fCPPplgOc4
HVG7vdJDk4RLKcJmSpX8ZJ8Gr/aLnD0FSfvYOI8LiFenOdMBbueIHq9LlkdaPW6rEZpXiPVqD+1Y
7HY9NnS0dL+xwdC8M9w0y+T84WN5M7uSqNndGhmBICkXCpMZCbKexipHNlY0zswg9zuUGS2gvSGD
XOeU1djlbyF03i8Q6zSi6l4/dTSpMn5yv7sLZF4g4bZHroTU5/F/D1fBXgKeMiRflk8BGwW3vYqK
E3KT4EsIv6NRtTu4t+0JGFBDY19J7gofwFJi4N5H22nJHbvV04rmJ/0tdI84wG1Z1PdhLuKJHgqa
gwo752v2FqR/UHTtqGKnxnu3mswPxtUXmpg6iG4cm2DbKJDLxw6LzrFWvN3bH850PO7aF/Jvyi1M
YHEfe/M+m+V3e48NKwgqYlvExYd49FFwkM7uAK0LsgZ4dH/4XFhpowNx3uaX4a5dQWK/GXBqMxbo
N04JgYg9LvIviGrE/YWuAPt+qcz6/o9HMtEfk+c7YAc+0nE6wo+Qb1YjjTf4VEJwSm+B1sZRsemH
mRsJk5sdW73pBPB1ewoXZ7bC2ObnYdXudKqUg6sn5GZwkh/B94HqHSArV/pQOYVcl2mS5xkGrqHc
6c233kfgabudPdjvMhhvHEXYxTBmMd0FdAM5PO9+B6ZeMRc/UTjS1KjNE/68I0UexGA4Fu5zAg8F
lWQvCwEHFuxmAianpPydXetst4uTvHE3HhU0YnT8mU+uQGm9D4jaB/Us+E6/Q/V8KvYlYzWUmhZ+
k/vtBjyVoY9RBaB1sp9IjQDPRN4YazvlDY7Rz4LIxiobJUG9yLjRv15+8xpx3luzvLMpskkkYYy3
/krLkBNXDZKLQNuDnrFjwV0LP2G2LGzHV3kDMKvVVP90UIzW0VtSBIT6dkS9ghfdr3fLxO2zhrzP
l1t8ESgTR4yC87wELRrt285zHDiPgnmr2aE3Ms+cAbxDZS2NZseiPLtUYQOjvjSW7J6xgDl/kIbR
orhDLamtM0ssvazvqXrcojC2B6v4ZbMCIlST+l59I9YYaQiC1+0hCm8Z539v0oIe4kQDFKP5Undj
P9oYruDmKgD2rrCg1ncR1q/abbd+blNAzobNM6nGM7IEwQM8z1UyBiKNJ7lkovW/2k+DJvtSdXgJ
sy17teYOO1d0/1yhB7N/3iyVLNFoOY5wOxo5jPm0UekXb4T/8SF7kLtNfqyMPVI+QftEc2qX6Avi
W1uN3pqlQx7+qar7M262Elil5Z7plOuHWidoymSiPtgj0R1vTo6FghaYDMywT8eoOO/8EeGgDA+M
qpAXuT3DuUuoUDuxYO3NDx9j68OmEm02fhj2f5LLun/tbQkVrvFwaywFvxoF0/S89QfKFcbNR3pe
7cHlXTAwG3rEjcZXBf9FqW/7xr7SU2/Xp0nC+Oc9qih2hA0Lp6HhWWdZimbE6sm6Bg04YvsSKCti
HLpduoWkX9Uk8LMo5mo2j+VMf5CfklA75tNCvIDc7SjRPuiNuapbsxSJjg/HTrTxLlYpez4toIu6
oefg5w5LGYbm5n+DCp2D+1uYEIHx4XbDCPqhdftOkPdEp+oPrnbytoPH520YD3vDjCz+hDgVWNwY
VRdQlij/5KENbC1jmQBO1KSzDNfvkhIZZvld3gA2C1NSv8NHl/Xy5xrRh/htDp2vlxNNYKDdWWoA
aP4i7pUvSfEXerU4dAJGYiDpHY/tGYi3p9L3OqR7vP6+n/s7OqsA40+IFQ+blp8Ja3bnV5aHWl5n
t9tdokK8EDcKDXNF+woPX/x2Zx6pupr2e72flHIrZiGqC+WG+y1ot2E7suo9saKho5zqR4sorio7
LDwvmoNhXh7rCJOU0F7gKw9g2nKJLE9HlttQguEEY1H857nQGgoN3xRpWnf6GaSX3anpQNeboavo
qYCkTonnjjFb5zwOmYYlFGUO+txNXmVuyhWLRfsascFCUa/cf2gk6BIs3HqiYXkaNxAhkCThpAs9
5xxyCYt+X5jsNxdJGECaugcWoeV0WyfelGV+gYfnwhIy0hjgqFsmU405ILred9Cb0WI6moLescaT
l7VpK0vvMDQ3mLyfgZOuZA+OKHIPqmHTtMNhz6ApBLUiCjI38jWC0ZBgWVySn1qyvi6UuArCdinY
sVLGMC/2BbJtp7VaP5i8Ura4KCiYmhMNGjmBq/kwBXPJXbqYox691NI8Hv+y4BCwv784tp9fIKRg
CAdMFniLDQJGg7P8oUinAOGdyUIXh4y3NB7r7hL5z0s6NVqZGIWkMsc5HTQAT5doayCIx/cheyAg
prKuybKtsvke3IKWAB6ZQt9dF2+FiKe8nvIcK4GoFreiKZpOi9YMQedWB7YwALxVCDzN2+otG+Jl
PMLyCcYS3YO0WZ++oTxtHt6yItQ0T/kMhDzD/3mR1+TcnOIbvGHJ2aXUAhv/0fUb6uI2qLTc4KDP
fFLs09BUDVssdKOWCcRaW4TVWQYugMujE7TiwvoznBRv7hjqZG+nWat+P2ON6Qqwhgnt2QOBezdm
q5t8a/mNi5KNa+LJim2uXILZbpuUJZiVXeZ4VdozuiPPVa/4z+g6IoBDtDEcSPEuX+K0bihFleOX
o9ySsNfskUgjG6Ebk/PcxP6JCF6XIcRMaZVorp1rBk16EzBtC6IZ5L5jJjOLMKX37knRAF3MuWAe
2p7Hy5mFKLxebVn5ix+GqZo7tm9fzPNymu0t6QuD3q3IbWCGumWgqHztC/wN7erbKW839iqTg+YE
ZZ+QBvM6tivq119q+OPc9XjJldw1Idx55MKWcg07xut004+/61mFwCbrdqLcJXNJTmj6o7wFGp4Z
Bqsgih3m+FKlfveisnGmOeDv0Ws5BqG9t+RWILBLZ29pB3nfQuLQGWqZ3pQJhfpd1X6woj340kFy
Y2q44/HcuuuRvgKnNTtnY46yQG0d56oMeXSO2vtgLTOhriUKYzAmBhS/OAFgL4T4eD8jVkjn17yW
KNAoYl3EbXlOgBG13nfvoyM2LbbgywklUmOlDgYGX5SCdKUKp2UzYHO4h29FUP4UN60no9SA1J7L
btBObC7mdaH4kYFLLL4NWINzg//CoSwNBtcObbfxSZ2JsoquI2R8/SOarRjWs4k+Co7IPNgtasGR
6fK7FK6+ubpmGJ1VQKyk3WSCFzTc561ZpWUI6u8rIUpMgFsV7zrUQnIZmQDL+z56Xf5sPITUShYD
1VKB0KdbvnauE4bxY+ssgEcSRSbKum8sO12Fl0wfnVbfCERmYbY2eACmACEill1GCd6t2q+mUyGE
yJzFS5daFMzWmN497x/QJf3t1ma8w/BYHZwZ4d/md79xY4CJnEniwzDkS0UIgYx0/Cl4sc7ivrx7
C9wOetEFb19GzF1Q/fSHTTr8S8tlxTpRUqguY9ytlvg9xfDiUN+TmeUBoga4pljcBA4e+E19Yi2n
zn7lDoU2WgdyEBs3O5YYC1wW6V2MXtLBbdddG0E+neYHhAi5+K8zQdOZw8AI9UjHWVYEEA5gtyqY
PFzlJl24mgQWwve5CuZZlFDpKXpPV7LSrDUHVu0NNB4+683aa6j7Q8TXrpJGVTYFi9wR6zc00pbN
8/y6ASc6Y3oI3OGIl9F6fnJOigRBkMpV5Fmxw0LmbYOg6JaJYaBLrJH6bOpcXvt50QQf518u8B8R
OzwmPqY6zo472lpg93XncHmur2f+gMTFmVKG/vepFuRzfHI0rCzUstBZU0nJq597iYhJjRlGxVum
LmgUz8YI3XTt0a/MIv7twuPjqVY+ZR46wDMzRN0IuLcbfy01xbIvEY6A4ddJhrJV3vzesFUePfQP
1gTG59rJm+uHn4szAD2S0kGTqOPaaTMK4ZET7F/59h8vnzQAyghYfFeG/+Hy3ZlAau3nwgUVFIBx
hHVZi+zFOb1b7L9lKn837HEQ0VD8/GNc2SMz3h+ho4c5eVglZWGBKEg+LzRpymoyW5XZOV0WVagi
C3QU1Fbr9epbc//eZv9Iy4CSUi40ew4V18YXsMvodfRqwTiBvoWbMqXyRbru40j5/iFid4vXP++8
Tq003MqBWYNxse5FD2VAezT6cfRT1y7QeRr5wXEVK15/KTWHCgBjuGV6b2m1Cfw6TOynovd1PgqJ
AHXsfJU3FH8CbMpNujuUCOZtOiFOoSq6Dn5ICYxSkeVT1Yw6699OwSkHqdKEbUMPBrT/ek2UlI97
Vp6JsWIZ91itXKb8JcfG7bFompWDzjAdOH0+GoyWMc9nmZfRW8nyHQ5X/ewGUSOIBB1aBmZLC2F5
XvBbydZ4nuN8ua+ur1xSyEThpPKxZKCZzeGkJYSYPtz6mWyAoUiaMp6BveXNi90fBB7yJH3hzLOw
fw1fsqC/LZS2MFzeDhpPx8lQWIQFOtMHF+fXEKNzxE1iPGjetF1HD4bkzQjR61g7Z0+4B/zZ0W/S
i+Z9P4i8l+m0TKIqcrzBLfYmZfjNXKOyNnMHRwvJ3vHAojfSKLbTHX56dBd1JosAhWJsNW1M9zq1
Y88o/NWmIOrf7pmqg7uVN89s95kKO0beKFgPPxExmSJfM3GoleLDQxWwiM3C6eIAAuRma42/Z7OM
XenKtpziXYVvFeuI3JqbwoUKcbZs1SAxI8KWGELYM45u6xZL6zasyEcn4KWus3mmVTdZwINFDmHf
RT54mGVU2Nv9+9Kad3W37PC0mm0HaqwzcjckdjVNmhbO2l25Wp1RHhdizC2JDpAT6xZJXisID1Zy
+ZW3j9kSgFp2RSKr4ogWZ4rUwExqAHV32Cw8+jEciaAIMXMJMZKDwNU3JDEWTs5AoQEANnc1nlZ1
5M3V7+7kg3fTgVOxKwbTMZfBUkETfaspmhUf3XbgNRwb84e4kjAgSP31tptnD8j3bwoWatzcAs6z
+Fbk+BO0RW43npX8jnmmqsUI4a32e1spvdHowEMZLW8hB/5xCts3pTEq1tERpkmob/Skc5oeSws4
lKykpP65pj8rMI6uD4q7NfikTu9YRYVVo1dT+8q3OF+4cHeJ7fnR4xZLoRqwhi4yFZaq/ySY03Gn
qH0VNC14KryfHKmSEIGnQkLnR0csiwWcTPVe6lb3+LdmhWQRjjPtBJMd9iTKazWFJt7YK5B6LMdT
whqtvfwPy2KjM9pwXJp9jvxqFnwMwMjMl6t59HcpJW9j3oqvBzXxGVagMaTSzJJTTmc+yw0E1DFp
SdQ8tDz5cJ+AwbRnURJEEto/vMkq7xZqN16GTB0nB+mwC1bsAZ6ld4NS5Vt3SCAxy7lvG7B+X9tv
Sx1ELlreapaKfueGKiijzYjHyGF8GYIeUyRyksoZe62LmCuK5+AHROjuop2E2Zhk2olpLziS+vnR
z4+Con9ekTI7EpY6Od+NmRDJxZtX305Bumv2GtljsEJ/uohj3hm+Z+ptbRpH2X2pMuk30SjvzlAw
SYKJzRroK57+QEiTqcwnz+HVAFUgiRaG/2Th1KsWvUzHTS6/i5sNBpvPO6zgScKzFIqN02ZFB6aH
N6rflwNHjMWZE9aY++uYoff8Um7rSdsTFG//8oNUnbec9UOLi03B+TYMuPks5KIAVWFek8YbUEQ5
sZpPhzwhxuaM5HkvGjQI7PVEE2X8EN7yo2Y8O93ahjEKxXkqx6xBm5A+gJjwshb9PG1R15kpZAWL
GR8D3j0yaumbvIodSyvN+ZkSbKJx7ZfiYTiI0nIWAE597kgHQbbqb681Uc8KFNfswP127a/G6EH4
CT4mjfpRTKHQzqszjUwMYigwDbQqwi7wp0/bv62LhFW8kquym/2QiJfSlPyfinYYh3Fd571wyerT
KZ5Et4NVYOMozK1jSXZqaa8XA61fQsOwVk2DsbYGkiN0BIiQPPFy7J0xNwbDbqjjEHDTiEDmLrQh
fViBGllkJYe89ISrGLHW3CMLirxxZe1YMOJmujO7ydOzRaYykJ3TmbXUxeAV/3Q+/ZraAWB/v11K
OStaBskW9k9RHbEuQJ+8my7/aTHiGF5Dmjt8XrwaEMa/pNSFTyuA+NE96+yC9Ili7PuvU1UjczOh
cy0iU39UAUzY0+FJzVRlmhjiTG12RwhpORkkvRySpClquf0n+AfEc9VXuG0hUs74Q9GO2aThSwbd
YvZUC+QV3kZzu5vz48f0ElBy6AsoR0lB7rYBjXbzEd60RZeO/Ucoxh0n06xKHVzuhkU77drUvF9u
mBYtPaEnYylRGGURLbkORHQgG+0eTsO22jFZ6Nn/ejKn+77QN6gtgJx8sjuvZqAnDGgT/kJnOMpN
Ky1InRVBBjre2M5J56KlivlZzqqyqWBfs8KhF+Vo5nqkaZcxb5VS/9W014zwUCteUuczU6cm6gGN
1qt3Ffko8bxCt6cJuzlLPZvsC+1Vq+ha6ysh3BZfWJlpwuRuPNvWUXl8YvDgmGipYEoaWMKuetlI
EUhoHzPnhTvURFb7YbP66I0WVhySWKrMYdz841gdpWW6vXRnT98aY3Ee2VxUhx+te62Waq/msbV0
/gEANNPrFbMzjFkez/K3j55iBtUuFTkmpefoS/M7XrUOjOowM/ywyivGF/4LQIVG6HcwbTRDIESg
tu5v/uIJqg39UsWWyn0hatDVs+DEOmj8RRG5L/ueW3pj1IR2Tud3rI3ro87MhE8P31vm4nn4Hd8Q
4gIp8UwULFPrvTlWhlWjX1YZZFMbIjnwovlG+eB9ZflAhW+g2g1lQBTL91EChNC7I6B2Np4ZIjhm
Vm2NVBW/gDXDr7i5CY8Zeue5DbsG9BPvJ2iAag0R3lL16bIfCqSVxFuDj+KDpb16lamf1nbUhFK4
EwXMPVtV4O+IwkuAmBZ6BsDknJMrk/ID7abLAlwhylvTxMA1Cxq1UGsammhwHlXmoUm17GD57T7E
572gyJYlAHwWGh/lLPOYM51yKzJ5VN8NuxhhFHtdlGE+dWdEoh1u/XdT1FzImRPUS+1xQZprQqrU
PhXEDMdB6BKgdXs9xctcxLpFfmTwRe5YBMsQlWdgbh5HRSvV9wjc++dWyhacoO0R9ERmPzHEMWKM
Hoxx1NJ17Ueq+pmmo6hHR0nWcwiqUmEEtPBZGVPva+KQAQE/F8LgtF8K7TGh7IVaBYALGCw4Xg+4
4sm3HOMJTHXC+oWhyEtXMSr3abc/TDMYBQn4uqEvfUBC4MsGu3KZm+5yPK3zLoT9vjkbv0LJDRdX
sL7dtrciuA1RhlG5xv0R75CzN0c5GZMaKK9DKj5YwAcb1kf3G3e94uYgBrd4Tu8fbO2Ft3ArpgGK
9Ukh2Ow15yoU0OBuc+LJqa3dm8wuMBo8VwcEQmEEt+1yNi3K2D9QMi7l1Nc+R5T8ICFpdzx46Vh8
gXnQmtonTRWRz69A8sM7zKIZZDXhqfYRK6QymVseDws3kAt97+5aTOnaq/vgUOGRTOcWlmuldGMt
K4fEISZ8aNw6F3S5vIR4FMw5ENhGYu42LidLMu7yQ4PDmVvD1+1jFoC1aN46UnAn7IhXf6rL++xY
7W9S/rBqRLkGJs4eWQmqC1J+p90RVArw4IrH9gexZOjIAWfW89qd1avFL+ANJ64x1hX0HMHMho7r
mEnytH67HFyNLKrS1gE/0yRdCxjRvQ+K/K29Iq7PbjoEdIisFJ6mQRFnKxK3v0lno8hg325Nn2Rx
OQsgpbM1rK+rD59PP3xhxJtApNqkfcCUYSE32SxbPtaw53/KhM4a40JQPG+r+27fJkjC8hmWcO6I
mikFAMciQvv0BgAWwvmKjrYT6RDHh+0TCbSzw8Md+pQIGTw5+Ia79fTp2p3vYoe67JnASzexrrzJ
s/qFNjxWdo3cpijZYulYTsLtZQu88Z735unMmZTGdIaXFxK/4br/wMEbZeGi1otTiPKruJ5X9+Bu
BQw1Zrv1dR+eQriLmVYq6brlgSDCTyi2TXCdLAEdBKkj8wE6EZByyvgmCUeJhvaASCXs2AQOJ0HD
hqbu2IcR631/S8hCFfHSlZaNd6Kbii8IJ5ifzhuVXtnZW/v55hPHMu0HSgsHZ/gR1+ohVnNIDDf+
qtYStED5G4rWoSxlBNH8TgngzFWYyXesYQk5UG44n7kojcy0xvVaYTIg0WjbJ4uFUr+yrKjPUx+Q
5s77Da8UX/ONj3OS5PfuK7zuxdbT8JNtbHpTveQkvGJvPLz5HRGo4dlj3Hgk4KIWygO6HHSYXXmN
ZhyyMNCPevHt0SdpjqYCly/dLBV4RmEP4nF0W7qVkP5nmkl+9mEJa/40UwjmmNsyKCJ6Wj3OlF9i
nkK5D12PmOuTSQOrFjlhP89CAdVQ1ww13OKcN482DYPDgNJCPghRN613gqi9KwZJTcLMhTqEwScE
FxB7uI8adq0Vju416koyJOHjLw1Ar4sYfwJRQY01y6NTsDD9xYa9uzG6DpJCCmSvu6dTXoTiuykV
O5rhMpNFz7jS6JbLoj5AekDI9A5QCr3Xh33GNbGxQgdX1FwDYcKFHS2NDAE1J9Qoid7uZxxSW77Y
eTRfuKBtyRnVE7ypj39jwiJ3yZmrKi01jeCQ4WZWYOhTxFPYGCjNnh+vrQKe937nPfWnkk7JeteG
tk0As8VXwvnuKXU2skhRM/JvKxcyaUvskhmXIdsRjs/TsAwRlUROw3w9HcH5mLihxt8gJ9lF2xig
APhX94Ix2SBHoa7GCmteN2qM8oGaXZ6+rBr1cfhMyLW5btFrnQiLqpFlIwDo+alhlrvfJhKYTlQ6
JQpSFyBPo7t4+WfVz+0YO3uQtpPaJ7Rf9WvT//Qk0zO7oRLN5NPmWD7oawaNpR/JAC1aMQcjNd+e
MQRRY6R8R+VGtd1p5FinwojUsCq2vY1S1xY2SZaAkM7rbNOiKFuB8RAcDEgDjcZ+hv9QQ3kG7nT3
gXj1ptiesu7ppCPrLzSLcMln9tf6ckLoWGHhuHqy90DhpIUp/CRNhLy2PSlFZt32OW+3mUTT+LQG
tEYlB1tZgXVWkHB2n+CPVK3+tHw5P8BK2ovefCeRZ3nWgZsGSvysNOx3360lkVw5lZ8TsK7xPQ/d
Bv75N9R3HhViNZZnWvXOIjr1Py/ghFyk25hEqmsCRZFG7EyUkHhl5qMG7ZAuMiul4ekdNeGpqIRg
N/LbdbxV9PjXNLvCW7acJ/yjxxgZfpR4ZYZyS5jaEJpHjYHASAAlEe4H3ybEhmOGnZ0kyl/D6SgW
nVdUp0MK87bK/bhbWTn5nmXEK8s/qnVTRtEHJz0iUMFxnSEKH59bCtvRznXKbKkX+Vl+mTQzjuUE
3S3pUGq1ya6yKT0g4yVkPsWVeuUFJ9b6VbwSSov9cQI46rGhNb9YB+RfMRWzhyjIceMkeid4MOxt
FeuJOzYCp1ERl6p0UrfUUHRHzAxc/Kjw6ECMvfBXi6DckV4ZzjYPZsm/s9Y9+JjRE2GAexmbOahI
UI1crBRjwCwaN/uHR5Sh/vxa8SEQvipa8PlStKf/v1iEjp3l4QnuZ2XsIhFMYfctuMJgxdJP0q5o
b2yYgmZxUEKaZAXNangTCkvIovvckjW8tkl3rE9eSi2sbX1amrcx3jbnc/CMkZ6J/2JbDWoiLIDI
jSNAJwmNDc/c4zkNNyuidKaNaPKIf+6IDtMhg1hyi2bIzUf2wG02UEc5aA13hiP7QalzVJBoMZdF
9fvPUHkXYfvEWxy9m3XIac7W+a4EOj/yb8dC6Y+k+IoFZyHpLWmvg8cFTCbjwl9Ad1PJXi6vWek4
OiXdV9umQ6GX2POaC0Opw62pFNoYw7mCZen0r5qcRaC5CXva69YgptQkKKK79px80sPPjqwJEt1g
mpY+oqk3+ZwSJxL+h4jKgx0+spqklAf2v0a+kV60+RN2XvVI52aGAOMPVVD14n5PO6nfLjLLVM/Z
uNl+icayurESRzvAWdB7tfvGxgxYlxToaBcy7keipSLLhLsmrP68T7vlJm6YIC2oYZonSMDSYteG
ADfkYAQ5gIN+xDVHbVtDYBRUJKmQYWbXD5s6Pg4hBrbXVmlJFywgzfnoloyI9fIoM5sLE0zeZyTg
MGTLnZ4mQ860vHhDiezm8KGGd+hcibJHfZ0w0l4oja1b0KA9iWmFhZhVQS/ajjZbgvgBsVfxutE+
TIEnWyVSm3YsqUD8foBxegcZt59DpzeZJRfBpUvIZ7bMDpipcWPU68c/9+xR12EFG9gtZgteh42h
eDb93d7MNUXlhTAmUmiNR8b4SXEC/orM4Oa/Hcp3cUeGOdwMhTckPBhDidcLV1WbaJTd4JeUEXrt
spj05lxoO7e+eKYhoxFNMkBpWfclTSvUS6ltQRbZ3T883FqkK8NBcaw0OchxIq1WjWYkZ2ydAR36
6YauZhDfZDSumelDmP6MCXJmpI7MsyNqf2nojXJZ7aUkzAPdI+ZrP/75aAA2iCNmcvTdyIgg2gVi
DJs1kGD9gE9ssuB6e6OJUnRADxgbLuwg3cylZzX624kIxHmul2aekWVZAB9PWBW9fIi0HBptttsX
tQJyo3GxUk0imRxlFHAEYOMEpS/ImVja339l20uv3W2GTH4tZrkrPlMnGs2nb4DLfVKCPxPXDdlq
o9OaWOlgeeI0/y0CQI/9FCibr3wWWgTsUA1IgWxb0b+CZTmLQ9AqeqOWqdObEUQm1G4yYab1IXay
05LGlKdzYyFNrRA4j6BF1XB/DaEBHrQYKk+cLRcw+Bmt9SK3lEVRUD3HW4uLYfUCMS0Y90q2UPCY
XESROX2UJu12GZ5LEo8jhkwvTZ8FAFn1zUzOZLwlQbthhYC6hwqgMAmvtwWr91oY7kIbL+okmBAi
cdTzg4DiDYSfzX+fdvqSou8+bOXYmDfkCcYnmGb2QnWpZnA6IRUBhgQad/OsB/0FPljovF5HTiVY
1qVz26f9HtUBHFVA6KqeXMHJk//MdY6wHZGo3uh9SkzcZZni+9WQImUKEfl7++4o9XGon98d4X5o
eR/ryMjGVW+paxAd9MiIyVmImU4x5X4dTC7ZkP+RcYfmlsvLN4YazmevzIpsHDt8NKvB6e0wdxaU
CqHo4NzAcPRascXfxVPdMVMLzwvej6Etf0TXvoxg5AMJR9AeUEHICp+S6/2YM+F7LXr5dvrvCTcU
ROrlh/IeraptSbqdU4Jh1xdJeUmuR42auNIoH5d4XxvUVergTQhdXuknF0rKd8Zd7MSzaj48a4aU
SpV72RqyL+rY3vPl5rK75b5V56IZrXEKDEPWrTiib1lfb3Aj0RjOSUTPBeSroBZ9lxTOwNp1aMPq
UO3Z56vYRigGMdbw5Zw/FJIM6oWFJ2CwivTL4xjZ4n/OEo50V9k4lKc1e1K7pJmfOcHaAHquQcFN
3XMY24r2ZeV2jLJNoyFP6hg7yNLDAxoaU8w3cK0wTPLASDQHHyJBkMNGr2RFt8QwIj0umrTjDEML
4PevAgONMTrKBZQidl17pe7uQnpWEPwRplFQvIz2v6HyYrWAGPyeaS7bEVrOrqh73PGoihqU8Mq+
9aK9g5+GZM4Li/6sPaJ6YXJ0L3JiqUc2UTnSARNO2dlFzIObMPobyE81/KoTJserLjUiVWquaUHE
iFpYJQ1+HpIlq/qyNMKBgLrRh/qILibR8aPlUPQ3fCmWMqGeIFHhgBitgcH2vUHRIJJkCX2jNHYl
YBGzmkGMCm6BwUWBgEomnZdv4sFYU6MvE+SIak1TTxfvTB9r2cc3T5SdauLZLA+7OLBYEWRccYNt
C5QClCOQQrf1SZyQ5PQiAOT4cYu4ppIMp5XCXhGZRxCgXJ1M+f/xH+EvzcxPjZlaurKacqE55kvZ
8USqywaObpLkuxQhCB65x70Q8w2rAK7J7VH18wqk+bx7tT1SXOvlesEmp5h8JAPpld+TdeHl9QdC
ojCOVXLTv7hrWR0XXjIDZ8GxZ8PfHQPBxi6poNCz7SpUPXImNYtzGUpvNrEVKkQr6u2ta3KRHesT
Qza4ukVkVdMBZOg9lXKewwv0DjGxS9+ejydDYDSwHen5dn6g/xouKjQQ3OKYDyd1HlSgOztoon/e
/pXwjtRm2Xbhbdmg83/wIo52O3HRvCBgJIDAXcAV/Ks3WkM8zJlyiD+5IFfmImueoRcE8j/Y1YIV
nqdCMaexb+Qgo+x3ne3ns9q9LLVfqzGAr1Aksa8VR/OLbr1ZZDW63vhypfjDxaps3wG/j+Ez7UXu
5bofihvcHSFN/mjk5/cGeq/xvpKC0TjyNXZ3enmo8BSJOKgcZAr15wWI2NAN3cjoXmaHkCL/ddst
nBic9CpsaaFg4gnFNz2ql7fB2ZXZeRn6DOA9h5e03EhSgQqqRX1nF2P10DHFZRkEEFuVZwMmvMg2
fUoGoZvIY+IDSJ34seszWsEzTri75oDkb50QaYI7dPDct8Nh64tmh0ZPBp0fJfsLO4tyqhdSD3Ee
pOax+WbfEFCVcDYn8InowmIRS+pPOQYdi1JX6v0OLEij6GIRV9Gk3Q9j4jmg1m93VIBNWLbzF4+A
bVWuZjNZFfsFsGWaP4NkBGBHMAq0/D9A5w5tbNnFhepahCo5NQIvu0uWbUwihMvgBLmLGcLVW9rL
EzJwC3/9TnN7d0GYCEXHnvvk5au4lcheK3cS3Rlxz8BjFbyh+kAVpxXhNjRp17tQZ7rTpQP1Z7O/
uKZRaWwqwiGvjEAvK85rb1sji208/AbjImuyisq2+nkRusYSrqdks/LSK9myBsjV9HZC12b/e+x/
Ylwyq3Bi1jMGNXlbuQSKthagaOER2rPQyRY42Wiv4ObeHUPQQc4THTME6O+aqbCqaOsLrSFrkmnd
QkSWEsAoTbo2n5g9AUBdR0TcTPalDdMdalA/qImV/0V3Vg88DmYw+35x4TO15Je/+W6uKkKVO+XT
9+1SVVGGufn1+HGumX1Iar7qLW7mjgIDitAn3q9DSUWvcudVNdwPXnnR7VIzY3T5CxjSxcNgyjWA
1T5LDBlaujYAVoRwMcusX8+SDg++k9wN909DP071RQgjT+w2IwEormiMjQncTRwTb1NW75MoSKew
UXQuEi5cjFNzu33pM3ibBhhTe0HmxzVBtHg4ZK1D3FCWC5EOX3yxyLLcm2y4QX4vFVb8YzXrURsQ
/q/dmJ2OgvAV0s9E6lbkYDlIyc7YvOuknovV3nkfccKqcdeGJOqTDVp2R6Do9gKZhsMnLeLlmebh
cQuG6R4ANztiY4P357T37+QaCokTxjWjv/mY//10mBvK2h1soWuoh9ypOZXf8JKePJzlV2E+3FxO
vFdDlcArTSMFeLljCqf7YuFrhr+dT64CkI/YLFksRQUL6mMdMrAXvzAjBbQ3acxQ4u8gTtKCgTvK
LQ0OxXxmGekrVQxVqme6+lZhy8UKTbZjtyOREshOuy/l+mmtRykYVhikAT5jOB+inZqZMeEbupCt
+xETPw3l2L62pBL8X5BkaPEjS8O+ZOziUZP0XwK+2G93pdsvpE73ow+HdMhXNKjYd+PIqGNJ+8ku
TQijIlqlbf3bE1jX6QUVweI/Zk0uSqKO2yv8sSLJSm50r1hGgnMQO5RtuTiHMhPN1TUIYzFNcwN+
k7Snxfyz80iZGJf1gw3O8TsvD10zuVmum7CKyaKGIoc05cnmT00U4VxzZT88UbqOHnO7zcw/8COe
u+qBe1Gbm8u2h0LCScBrakQe4qzu8OFfxmF+GJzYJj5/imIOqXdWHcbFeHL75M4zPRcq64u9A8hC
LGbC00VyE1ey1Ejc5Aau/jP/S4MzcvmZ4CLrnALKYTRDZbRV/vdjMSByFeoiZxvAGU9SKHRHtrTC
6bHKjqjb2iswgA0FPCWv+/D/6wJMcznlR7pYQjIuWFkWgoydnUaSMTLrxPbXlqavig0lngLThnTk
M30mHRptygmc1IS+g6ZFQLz31swO/xgRDUXMeIaqcqpbPHUA6sVhCtTgv3qLjDPZdC1vVrrsIU2M
FFHBpPyr+2xAv/Vv99cu0lyXoZWaBpmXxUnt0NYw2/ZUUYQklsfD0evrRAQqhFJ8JWwI7AzEBERA
WnQ9BoBe/bGlSaowsgeIHcoD9yJyPDntLPSHc3DAZI4wBXOFphP3d11UfXxSPg8DGS/A/lNJY7Yf
J0s9KTeinHxk/svIm+rXwUasv0kRW/TualrILwf7Y5BOhKD+FpXxZl8kzjU20QMStO+SvRVKmBQC
vjm3PDdEeki/7hmlAp+rXevKCnHbQIUR+OQj9Uf+dxSB+gbUPgI6L//yJAjy51jnfxXqLd5l6iq3
Dd+s2MD79BMuxy7qXcBH1J9CQc2tovVMjNsbRWlZqQbzuRyL3DwmMzSVvZNi9xktFQ/7RE0QZqa9
w0r7N7n8JFJDsPYa/W9Lanq3OvvrFpGJwHLlpEwmhrtLdwQW2li2tou1adMKwRr7HMi6VjcUDQsG
PCPhczg/e8xmyKm6MfHs4L1IN3q2TD4p2h1kjTX87dau56jUMolWHdntmKD7w++R1HvDh5zrZCWJ
7uy+55vIgJwVqe0P8X0m2S2L57fmtVxZJ66E25qgzGKdhxGDsAXYFeY1DJYtzTbH7zo+I58zgDZL
nr5MIhd92tERsD+p8cwN8UfeWqXP+1RhiFURZ/pAEIyCtr24W9t9hmbGNYA0VonT860KqGFZGw+n
x0BfV/CHb2tWXF8pN9mMVqSzKG9X2XMEU8kCC7I2gHhcqX5W9qlRX+9JtVhk9fiHNwW2uRpT4wt8
LoKKlNoLGphkJLuuxxJUIgHgTu9gi8IZ8LiK80LsQSGkdl7eDCNZk68zK2yGq7aG13wvbrJhYyso
nZ32M9qT0GUbINrTWI2KwI02qgTEZWZJJrZiWl23oEPV+A3TleTC1OsSn2TQwFNbIhKV2r/HGDo3
ulxY4Uzws3BiUdLt840+z9OHo3P1WGSBP063/nLoS/g7u7cEtLdzinRB6qg859YhFLfDth0XUlML
R1qs88NgOYtIIRUWbj+7IAtvmEAYQO4LmDOyIMJch7bPEd2Vzcbtz5Ch1RZ8iqnq8SuWCf9Ne3AC
n/RRYCt7GgOjexybBYYn/Jz1xq7z6zxUjAjFPVOJ9yJJE61qWyo1iqHhmFwnyhRoDlvtkXaKkDCQ
+ZqTPVtnjtYx0jQfWAccmxScNA8H7YldDVRDkezP3uEkR/lGkiHXqfDFZ9RIcbzZc3nO2qM4OQsW
PFoM6M5zUAI7Cc0MkkVed288sDYE/NM1MYtaYijyxU+mQaTbG4nE+LcIi3jNH0VjI5+o2NqfQYHd
0ZhbJJ9fW1MCbyQA2KG000F3KLr/Dck+0GyWIcvWe2fmKE0Ch+Zb52JlMCtK75EOO4YlTbrA6PCe
eu7CNWh95Dq35LNp+TqHxLvrwghz7DxCOeIjho2x/ytBh9O1WPbIaeg1R4RvLMwmd1IznwEClFLC
/Fi6EEVYfxtyWO1aDHyhqoEDW2pLusJwjgv1ZGMH6k1iqliXcjjqIr5cMzTUOeM9FTeGxo2uGAqW
0GTxSzx+v/1zeYkmZcoaWi3lvW3rHI4Vegs2zlGt3nVSza5oUNvbHtPJfj0i/XbhvEzusDWheQQe
YUo01b3bi0Yby0H1GjRYA9VYw7Kss47+LJGerCrHF8dUc5nxUPLrZe2obbsGOyfmeoi7RqK4PEV/
mztBgBphbJAN9saVY+CDS4JUmZ3sbOr5q6EYXGA+3QIsIybOoSYK+xY7XV0PbuVPnxRcjTJpBAHA
/yt0MhVDq3ync34rmGbHKbCusJFgo/X56KyRXnif9Q1R4d/OicBzaVUYIB7i0oRBfGqdESWWlksi
rqcutN2m2jcjDvlJaKO8sBfWYf43XLANtVHtPDwfbMimXAHIznWOQls1bIoQ5vd3X6J6ETsTg+4d
5/4VcxKGH93pal16Egd8XpFqdvnJ3ZMkscXmdqqk7UGQftPstjpv1Ry5Z8Q+aP8RwNjr9+mxK6R6
23qfg2mt2naEWQ7lkJYtn1vT5NKIW352tMV+FwQtZmaCdsQdrb9TVjMy9jd76B40dt52+6PHvqyV
C7zNPrDIKpDfTIVMVJVY1NWEdzNBdR3wt9R/e4phty58/+ITdp5tl4OEU2h0in1Nj+8Y9c4JEBYZ
8VpdtxtQZJGZXAEN8m91wnvW1p3r0+RPa4kt8n3ypjjuvLEhoL4SywPEYOdQSBL/b2eN6Pk//Hd2
0w50X+0xjjbpB7iR4qVmAX38FDu1IdgsHlLoelq1u5XwBHBYUnISe59N+PtX6d0nx32V1ngqHDU1
/Kd6TwbzuFPpgmfPa00SQuf6Ivzl5xvqnM5nsGiLk+LIvffi+vZ1inOFvPiF2l7ICDTbXg4Cifz8
mSwrtL5TYRxc4wrgVJAYAgLErVQXnhhp5PjJnugEAiK8twA/VtZIuyvECokYuaLx9MLoxRsGy52W
1lzKRpKF8MgCSzlZYEoQoubvDxQJIZU69D+pFqlT2KTpsnqRNU3IForkL3KR7hlz5HRufc+UJ0P5
1Yd2vP2b2fn8pN2A4wCOLhMzXwnmngz93ArCP7Q6mxQLyJYYHuQMvNBrOug9oMXIiKeVS3zcmNVy
uG0St5tZPYlO2RqPHVj0a3y//XHSDFCPFvrrHjAGnnbkIiBo+l8Rw1rwX09P1LQ2qriy46Agg02P
ehKvwW9BatvsVIoAG3jEHj/xcfFuQXykmR/4oTbmCaWuvfbhWTfiYENJkDivEi8sMRc++whccJ9C
B+nQ8ba3vVfBUFB00LYVe1MKRYUSGcfuAArafu18TOzMG6AhTUw8swJTE3vvXtfDxayRHPDiE4il
wvbqAjyEhWnf4b3vFLHLlgoBVPfzQHPSl/7K1EIq4uNs+8CCco3HcvCf81t7EMs3EtOqq0aCvGl6
Pwd6bmYQm293broWEjaGBVlgRUutzzoF5ry+dchBEiF1xBaj3GRN9R78THmGjAG0c5D1OsW1Sxuk
/d5QjNCpIRqa/2guzhYVAxX08bs4tGBm9bM91pUSvp4diEwVXQtA4pN7WZKooTRAjq0yrXJXltaG
xBMrJu36jbVjy3u5CJJYOOGUJtzefI5sZahNEnrw8rebT+5Yv5g3WPHaI9GTm2nnvBssDsHhPULg
btuvcELy9WKW0YKyWvRnhHo7VhI7VsieOmNZdNPxVB+7wBEeHZTsmzQ1UH2HwZNvHsDPxKJYeF7h
cDyx7zT4cmRBVkQQ3yHwCE5OVoq31hFPFl8S5d7nRSTIu+1+LWIpgaoBU2qk0AmjClIhgppsghv3
b2QFFhaSpgBwf1zMNbRUeJ8Doo/tKjB+0rAwL+XcfWmttl9b+h/8cH6nxb21+htLiCYeHFtr4X+/
aFk+nvZi5EyPkCSNSbboPEEmAYoFMxkAv23DgCe5C65/KCfQ5JxZqcaY2Am2DLqmn8LGbd6PezxJ
amK127g1QPRgfEo25dOQsHxgeL5AqAZqHRDsIWsRA+a4tz9xTGa2j+/hcUdp7I/Nc9il/cy9jucH
t8FYSljtJXfI93OF8x9kX0Z5cAU+NK82adv49xcmpP6gNRN8vktDBrIj3AD1rNjbLdsKuwKqZciE
iZJr16vOh8uEFOBYnnsTrVobcGUQyJAZcrauz8trBMl5gziLDqh77VScPFWI7YDjg3hfwomXHCyf
ce4S2uwyywuOwPIIEoj5qlyj0sMe5tga1vzP0YXJTyn47zSMFhmFIXJlf2lm0rmZlvbSQj8ACWx/
De5Cx2XIWZm9Bxfnhy9N6kZ3XlP1dISWrdaBxSGMNOQPSESpaX4I1bEhYg52wkLsLbY06G3Nf5aa
WOv0sezkK60uyCIt9a2ylgzZjV00GYRId0BfEtJQ48w2dimWuz2FoAlvz5PaAoqkQj6hUN3I7iYh
G+wlRUeXHViEcnGB1IDvqpRPcxaOxvyzurP6LgZ3HONjUeUTAHEeVc/njG1tsaDRmZ66BMk0ddid
/I4RnuzEvXzBOaFnd4+EJLR6VVM0fwYXVuf7F3tthW+sVWla8HFFWWe8E7GO0zRrElGD0dJiOlzA
FIwrZUQdRT9tmceAlMEgxubshc9ZWze/tfcv8QoMuOdjGgdWPJtAjIpI/U1n0+2v2KDPbKOjU/ke
J3nrXcPdq34o+QbQqAyrlHG0QQNOPYXXjcy/YE9pq38+w2C5/a+fjsadN5+kkWRgR8wlTQ9zpdWc
Z7WrPfddarvNN6xLsr+U3NwNDvJRTYBvMG27nHhw+esKXDJGcU1oQg6B4e4JblVN4QO7UT/K+jtw
2jNAX+TFTF90kMHwCvtDcjljPJ/S01ONae7FWNzx9l+kM2qMfMAske/FOrBz7Mk4R7nOC4aA8yYc
VzvK2XHqSavukI+Tuj6z9kg51HSyyFYbMl5Oal4UtOTOYuHm0c9dFpAba9E3U7ppt3sPEQbATF5a
vVT8nqCX1MZjJSeTMw67tW9QvbkoUt/3mGR/o629AKaDL2l0dAJIZG5UqZjnzFHT36d3Dqyb3Dgv
JAmHkMIQ7xz1uZX0jA8dDLeBPiXCgBR6VHe5p/mIhmHOXEYM319rIIeq7iZ/2YgIjvW1++FJ8mBX
3C9Yeq3dX76PzQ/skCYnqSwOU2RGGOusRybBqIvp8obu54jKoNgzHyNyJQRFOHGEbQC5ijW3t/0y
fvj2cjf0WiX6FknA+YnIA3HTz3Qo+IOOm7bqG9mrHXkmpJmz5TTfo1zF/VADtq5JtffNketk0fye
YqFt+FL9Wws5FeOcH6/9MZ2iudk1GaGVHcfgCMDe0l01RpUd3rVCnLHzoKwNcdCaJe5EDjz/LvBx
6RqtHc+jRpNPxHA6NewdRdX+E5ZQOV1ZMTshDZv1Bg5SEyodm3aoLQgCwJukaeWilUJoRBMKdaXi
OuZOfqUsO24XkqY/A1xUrLdozrigNTxo41pwyxF5Zbw9EGlPwvEcgUbvBxmy/dlu0yyDJGPP3TVM
sE7THV7BxtboCYTxsfdqtf+l3iIpGaWzyK1xktJ5kAWDIJioYkO3IARniZ10g4fGp7HQcQuBzqar
2z3DM/eI6C9lKE8HdsVLLB2vNCzphM37BGnCZCX8rPwJM3VVVFN2Kt7hMSI7o3eZPxBjxA3icjLO
B8h0dbBLBcXV7FTYMS30+vrtQQr1KxHrJklC2WoJ6JuC0h6/A1ygJGzo5IcQRmWk5dWYK7rYaaJq
ys1u8KU/mdtASVxRIyj4pr7XbAQ+TBAwTvbXK2y16HTXal08ClmZpJEKEWnEck8ktBdAZd0RZsUR
PiTV4jSm1hewZ/FdEHcXGDnjeHdVOr2odrIGH8q8rL74GjeDq6wyYge7iFFxwQLQyMu7jnUvtIbG
Pt9cY3+Hq8ocp4R476hUVmx3DLsZopUBG1Skni7zEBv4RNPoMB/haVb3LWrqiwOxlGwVEFeef2hF
MZbI8IYnz0OtA73hKyg28mQ+ez6nQIAjyo8C8gbH64hIoS0c9aMSES9wzY7yOOY0eLqAYFfoWaB5
rN77azCCHRmW+fwdJ9Cw1M1Zc4gjWby1d10LBdr+lrgnsIqDiKg5dyn8wiBm/8kDiIEoBcqbd0OK
2HbHgAKG84xt21YdfcJZrfOr/XIQ/LkMbAd6LHOlO7/AeZT9qQ2S376/IWwGGxUjqV4J7UHPTBw6
RHJ7yXyXmBYENljquucw4gUh694/1aNdIHE3t79zw6rNnMO+r2ygWA2JboeIQi0bhg/5IzcgiwLB
d6ac8bz1+31pAstESO42UHMj+DNN7j/eEDxJhlrl9CyPXzLt53FNW8SxAe5YXM3FuaRU2Eadn8Hf
+FdnpuuRL+C8xoU7QaowbCBV9ACy6XzHAOndT0Uq0qOsOfwTLNcfZ14exwQIMrnsuWTe+Ve1LzFy
ig4hEiQALZV+yxQqXdoErsliH0RxPb0y6FdxAWoBqcdcvyPVNJOku8rzqArmIXoYaN1WymX6Bm51
5HiJ1cml/qlmfKTJSWyI5WrC9RitD7QroguZKcbU78raLadQNXyR6kaVZf9wUuEiW3NqIt3CthK7
0eGFO2SEPWvUy8r6qEl05egmgS8zeoVyDJoUneqAYmLFwFqJObFadPt1Bf8FATQIR1ht/wH+bAKC
88dhc1jbtzQIERalCs+x1SeZhWm3DfRBOX+gpeX+Or40C1TH5XvRUBVds/U8zvrbk8Jq1tzffR+d
ro8AiC+YzyYR40lDklapX2v/ISHU9WQKP3YrrCKEPOUHTjSxcEHSpQ/GZcYn3zZPKSPZCkOdJkfl
TNLdyLbabTlzUG7tdJEa63062yF94NlQXJ6eN1sYc4zojNIwV5NhhuzVE311DeAMMF21nXLnk0Ab
beIWmiaKAET49j4YWoYWumxqHZFjwnk6u5sgzeEcDij+WSO6Qjt2UHlGFSamigRifhBheFhr0DEN
yBq7gFKPIWHxIHBGsl2woVcpSj84tYW0jXhPOGej7lxeqIXM2ep+WzmNWOx/87Erv1mySHwAB5/o
A945Wl7JUi8aVUkxJsYT6L/usWxxUoFUoKoGEzzdREJ4EZ3BppWjytmnx0/15JBzl129jKub5Xx+
aKhidaM9zoBSngRHnA6uD4MHe2dR9uwZ7KYNgQs59djFkpGJzBtUCyolhxafRqM80ebHiqdpbV9m
uYiHps/kckANA17x7Ti2xnV8eskl789EBxee8VXfKNPMn8byOjC4r5s6qW6WQVpdkyOr2wvCJ6Xp
7lZ0cbvHjIxF2VHQjAnUBV2S
`pragma protect end_protected
