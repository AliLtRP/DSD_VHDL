// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:35:43 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
ZlqhSEn4/pprh/cYPpJsDrLKoa6Msfsiqy1WyozrI62sYIBIp5p+kYYFUpr/jueR
UlcFar/CqZOKarX9G0IDqLjH1H13sBZHrGxANirEATQ51jSQl0ArXD75cmp2JgcM
LcJxfVBLNM6+oSnrOGkh9ijoG5dfMes4P2/Abi2KtMg=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 6416)
hKseRgSY+sC2LsrCoNUwsp9RAu0X/sFb6tgiRyHCJ9Rr8vktggb2G4M5S4JRl6wk
bVjRc76BJ6HUTQBsGPlV8IxuG7vzcCLtMSWG0BZIVH2E1CttlZcuxJXuAvzQc1z/
lSHkX5iDBEHp9WFePJVP1XO/HDKOwpQ9rLv9/54wSdb2sPA5fvTAfpGBB/xwc4ln
pDGHcDWhAsvIBFawuxLqe5kyPaVxIS4MTCDeJKdiGRvq+L8fuAYJd6ntlyG6fibG
+SHuvlm8Rzv4kdCmXFpXJIxtTvwc7V5oSCPQ41l90oPUYUWi+ISqAj5MB+gu93wy
ZwEvDHHL3l14k0BRi0Iwh9+pkQLF4v10461UdsprqCB/Cvu0HotiXBUhDCCL5IUG
xEHxK3VFamwrvNLMh0BNg905NWZltND1Lg9gcvXcsgLAWdh5RHdYieGhdLXiC5Zv
OMOAO3vfRyz+EUXWwFHk+UttgYSjUKzYP16pwq2gN/2FQeYO/pfdFiY0WeTiC5r6
JPyPvoCCLzru/fP41x7A7135b9jYGugNFVVRgAGbt8cQEV10Zaun9HgJbewwnrhq
W/Jj5dIzcwxx9IeuXJUSgWoomS+bf5frsrfU1yRsVr20ZpzXKPVzKexBdomVzNzs
aphjhSb6LZSxQtyCHLLKZ+kwPpPeAx7wxsQ4GPuka6iVMiMVEXhd9jgXWqa3trSD
C4RHpl8Z0tDsYhpkx6c5T2rQPw67u0xTLNJWbryckZOLkxkDjx9KJ0DXy4nUZPiN
RNNMGOwsKIG1byH1WfZBmbvuAT1D5a4rMEZ2RjOpUQvlPjheccOsa/rfau2kZnvH
ItDM4vsvwoGQNMtIlXODtQrNFL5RkuUa4dpcSdLGGDPf9lYKk7ZXU4GptzmJ7YHa
EswdJkE1OIOYEeFl7rTiV9QSqKQa7A30A3PnHch9or4SzJvxoO6kPtOjFvrU2iOe
SMpW7IKD/zTo+IXwwKm6pgt2PYoRSF/6XKbwB4H+6Uh0PTSpBBkNaGbaRYDaEFq0
6OTAANHyEz2xPhAuUQ8ePvNNATjpB0fijd+t44hFmzPRXM6/1zYnknegZP4v/b/J
KnfR+yqCPLjW3GojfVyz3KzHAy+XpmBNGszsfTHHnzW6TYcxylTjWe/6ffsNZ9vU
p4Pl72fA0fZMfKoNR0PP2GXarRl9iXSSoz6Zum8HBVDnfom1aDiSFUHjq7E/zHLq
cGXC3SAYn6a0CDYM6+ic+/yLq1tynn97VlgOElJECTrahwlw5VVlVO70kVV72Xat
u/KsvDsVJ0p9cSHcLKTZE7c86xH9o4Phj8DsMaWKhO7UvTdcBcm6Zwv3BU2vD27n
nwZm9eYfgdnaeRRzOZaVfD076/5hZH6+06x/XhD407xVF7dTLiCPHOxh/7NmPw7V
dGoHqo+ZqSjZPLBiaG+zpCm3SKwyfKa5fjY/N1ygRRi/kVagcGEZ9K/AcQoOJOYA
q2jZaVep97F8qNZacSXuZRSr2w06Hi6Lr6WPfQGjDGB02Q8jiIlw6jmG52QjOns2
phVDma45bv6nBrmMQ1bmU7bZZv9xnAfL9+hhX73KW1epsJuGMXJZj1+UTriGv57Q
cxAX1lKwdLwcvuizn/gKSwJlProPRZ8PR+KDdaxAAonC3aOUtjuvbq04aMIg+5GR
btJXkIh1Re273ra+C/ZLB2KMasfJ6BhaVX+YTUp3YHvlASE9Fw4AX30Qt+c2gRzJ
Ye686m2djjp2CKxpxqLjj2PzmB2EhKaYzTblHJRPJZBFqWDOKkzmVm3flaLQHYKg
XJJlSHDkuI5pEbCPaB8oOdwtiV4UqtlXMOD1dO7z+ELJy2PT2fFdQR7FMhVurbC4
79uD5ricH2DoDk9DTKXEltprPQNWhORtgbTdAA+1Jszy/KdbpA7XSh27BAL5o9Kt
njAZzcS0EJ010wNRx+aMTFj2Vvx3xbX4yosuyAoFO7/GHuMLV1DauBkfvE+4ZBTj
f6u/lIpEx6VnyjDWZM8MZSh3dNry4ranulWlLL7fsHNz5ZH+XUXc/5ga6OAoo5dF
PA7XyEcD1I8D43xjKzMyF1i0QyV4Ty963+mTAliLzAl0INWMtLOEO7B/L3Jhdnlf
LAwWZjQci9/DPsctNNhdVJcv8MA4PRdq4O2Frwo/MdLhhdGC9UjKdOxF62sSRW1F
90UsX86zMm013FnMDqisireHOo6OMr92ZsVJ+2l/pz+LeZzbBB/DwK6+mEjFlC2U
BnId8QXY4k5qbfafkWlOTx6khdFQeC+rSvIephfzVq5CLoLJy1OK9/iUSIUqHBAf
dIVaK6f4s55HVMGBpI7/3m+P67Qd9VV/YZ+u7h/EYwSOY1TltvYoGaThPJrjtDwT
dJRRerUiKxABEjHE7N7v9Dinz2dlE4vAUHHIYkPfOA80HkapUIs93UMSEAfrbvwm
pONfPJZgapupX61BzJpJxsZt+XVShXpTIgoo/QXUE6pedibAINsRHlYpPDL+2QKa
VTC0t3xO8udTjOn7XiYYjX10wXqiJIlCdMuLhdHMtK6MHu8+/Iz2MET0KOqnIcko
KL2y0CqcL/ljCtUI+HhWJJnF2VsPFis1m3dul5r9Ervv3WTZM78Tfhtq3tts2BvH
ScKtMUup4deG4m0Wb2IgpQ20atYN4I3ZOm0JrGkRHi6YNpLOx4ebk1nt7379UooH
AAOJWiH5uf2ApS0J+7BsBxFgK837ATrPXcy/6SxdG+T5V+7Q1prjCekbbAHACG4o
bnSE1hzRCmkDF2HfGwgZo8MF9xPjq5rYMiZXjL9uXvGQXU4Kg9xl0fkuV2aGVZqk
xCl5GGCIz4xSyqIp08r8WzY3hAHMzjOI/INhDNYDYHlKQjqyCSb3lPgYMmPiuXa6
AHpudRXQvgSymhtNZT0jmnXMCpuWfvWioLTe+Wmtb0FNRYafWq3ufxzXZPpOS6qs
tb5CjAAdxaHAElV52f8EZQGd+EF85IfV/wUY6orrQUP1mOU1xrYAYcuL+Sm5XhsQ
5++Qx1nypuDe3j4v50iEMLN5APwhjnoj6t1FGK/a8Cskz7TzRk6huOHuMkWdI4Vs
v8/xAwOU989pdJ3aVNL6MYTQUwGfraJ+bxMCTZzkjW4+N0DQPn2zLjwN/6ol89dN
wB5vEf5V5Dhf09YspQewVQNzlELVhUdqcOVEyWoLn8Y2sOhaEvnl5ivz0Z2j2ldf
U1BHCX6Imy/y1Z2Hvt9vX52RaO+FDZFOf4OYMwvBi9NjjyTVugY/OBBAvkJQYtzE
xFOrMOEqkMJhFvPLYHIUBvjNxYgnhMujT2iQ23E2w/YY80QTaYjgNj7fUgArGU4X
e8jq30o6OSg7jryuGwcLMtQbJ6NUcj9oyZT4XZqwFGS93+5ad/HuonUGz8T6HLIb
VBpaQ3HIJACjHIKgB3ZqDCMQdvQkV0gRq19g80KTyNh03colOy8a41d8ap6Zo70d
SdMGFAwIzVcK653WEIONBHt9lly1vXz2NoNZaxr/XEIi06ZCglmpLvVpBbFHwtXa
VP8CBNBS1vueJUV7NhgTXIFZ/MvsUYyYsbbJbQ4rQdWwwpQe3/CyWmvKM7UiKRP0
341uw4oD6roPOGwLQVfUEBnwAgA4Wwp93dbSJfAO8+gJtLDGbgXPIwa7KiXcilRw
hkojxlgsaHF8qlC0vq8+7i6j27NSyPUrXntPZVnnKuh8tN18q5PLJXMGq0AbJ8aw
MJuKYX+j66OQGsO/NJMx/IARIZW3tavl/4Mm56nH7BR0x4f++YEtlueNhkINj475
uj0hockl/ZI4XXsT8eF8+lA195TNTmGhG6hBiKb3QQE5R5yJh3fa0Tbh30bVEEeX
dVXWRhQhAJ+El3nt15IubNMD3rYOUR+Lu18OkyKuojcMh/UMyQy8dQ97QGM8WoBM
DXG5YGqQO8Ijtp9LJq2fVNQCznhfhn520yWg53tdahCjKRjXwY8YVxLSlCtm0u30
Ay4aA8uWeiQvafC2wr6s9/SGInhWsXua0VNnfXabzRoGBsnpXYQ6pxk7aH24fVxK
pkgZ7tkUkM1E3yot+Gp6GTgaaSGuxOgDr8wtFgdIqJya0Dmwm7ej3UCMtAcPg3tM
1FRawGvo7xBvtZg7PWWHuBRhsE6XMcwYFv8ABIOaTEigzRYOyNOfRM1BQp+/xnLI
QUMgsJoykc2yUHzVZAqHmbR7uoFgnNEdus1hYrMtkJtngdC2XF/1CDj3v86y47G9
XfkvhLl59rFffhcjnQhNhI8AvR+Hy2/hERVUwGX6zmGHvceov+LP4CeS0Jd2BNEh
Bljg4wS8zeegDpfKaMxp9ks66qpEZ4bMMri3qXQ03gJ9iKPcw0/aXNmWOKAeVm63
hoUSJNUuInOXmXEfNar87GnYN0DuPNpg8hDkNVqEj3yn2oD4xgH9RLdF+htxATSE
OVbLZtvnkz+k+tCnJnD0cHz2zhKtl0WADuIdJvWGcY+XtcILSc65xfcx8Oo3SBBh
KJW66x6rjwpC3g/7jxFQDbQoKnmKNRJpmUQgwyZErkH9/FGWOf+GNTmdpUSUArob
KvQOCidh/hXMK+A5yKy8rQALQWfDc8yMzFgEgaz3YP5H9wj/8eqqpNzkDPueHIPE
Mv3RTxcY4UQT+oz1BsFc97ZELobpGgrGwWHjsqqkmr3NyVEI72khk8A/6xXyhvOk
FSvrloWIcUnKuooL6C79XCXEzjQQfCnK8qhvK3RL8nYVzWjkUkemRsbMY+rSsx0T
Q1bVKLaQfqlQxF93k/kbU6dIh6WXmWbeuOtvuZJY2+SgZtDrI4TxN/smYa7Dv9+4
43HF+SRBQYLf0C/0qTk1LH0d/niKf2iP9W+ZGVm4ycNs8cJZIC8Qnr+DeBY9J/sH
ytKc7hsW4CH11iL+aJnvu8qvgBfCvpx4DuUU+4+Sd4ev/kyTD/jJytuAmwrkFyCB
+h34onNmfcd/G/iZ2ERbSVb/hoxZNb4TQA3v2PtFjxkCptgSGG6qq5ocYfzJoVUG
/QzHH+TFsfcPiC+Qg7IwEIcgzNNdmRLUtmVfBDgorgGUPzcg9jLrR2ATGODJFd4R
Puc+8ebVLDXABhhyyRLcPTlHxRRVhWX0EI3HbJV1s0mZMKH7FL/lwG45TwlIiXMi
pCyOO1Oke3U5gtPefsDuBx95f2MTMvQg4Gy9GmajNdYD2FlAeMBEtQ5lzz21Rm93
aeN96PQMjAoUeBJ995/zn6J76rsbrGhgq4itT/descpVfhcoaRmxzn6BRyW6Rtdu
USl64sf5H8oQ7CXWAW+kgTJ45zggzXXuCqpuiz64CBW5/NyFlNp+iA9ZtPbvQro6
s0dWYyEwDu0UkeJQEpI5jYKPelalaX479GHlLozjIPkNqn3BdyoDEIXkhJbkUmu8
KmZnxOCkAsh4ijC0EV13OoCbrM/zrh4hjh8JO+YgOwKPpq5FQiwpzLLRTUVhuQYF
fL9MNuTtLoJcnw03cmO6bnyphss9gD2MUW/4BtnfGdHptqW6oNv5o/eR8/KL0PLP
nRlu/23u4W8oOrzj1Bp4l5sNZFLgwyvInoYvNPhV7dg39i7jjCzj8KTYwcVyiZe4
HbRaa35gPy9Nrd2PWpZaMJqUyEM+X7F61R5CeLHXgnDs+XXS8wDIywZYtC9FGWHQ
IXYMzER0ctiSVs8GdmowkOCysofvc7LRbLz1GhlUe+DRaBMs6xcp/FOuY5K4Kz4b
k7lE4fGz64Fr4MaBy4J9TBnRgRx/ij7J3FMxqkO7G3GoAEjm+n9O3SvCwmLvmOfk
yDqGBgyUQdFWM/bKB1iFQ6U6nMg1VisfWUWMzdAJZLWTG91CcJ1u+AO8Cl6uABEP
Fj6ZDpmEztQr3+12mWBD14MqVpY1LHo1Z61S82RKqviYQmh6cNS/bNSu5EPtcjhT
ulAJsnHrIzKstCt6FD+i58SYSh70++DKYk6TP4auzV4+9AHrsZVrJYNHwj2won1y
/spy1eWfP/oWbiPUdzeBbTXJCtX/fSvgS46RCQiQdXJa64RYhML3+bGdG1ORr4XR
wxKjs5qEWd06lAtYRAqOZqcjsPMLECeSzPNBPG5vokNOz6VGiFmepuWMTC53wkDC
EfSF9bm688tfmWent2Ylb0iL6TT4rR4yM1uUip4if9BV5s/D71wA2g06mD64h+HL
YengyiRrtIAIxTdTd398F6TXfMvFwVuyGIuKa9TN6/ZJqRu+KFopBHrF7GsXGZyt
7GOylhVf80NcVlITZe9PI1wINMqCj24sguBNrGsLW+j1VWdclBivjLELB2KwmB4Y
qBcb53VMdDt+hWXU7DF3gyh8QxZqvXxXb1E8zn1ulN7twKO5DVdfVsbywuLCjUiE
1Sx+74Nvoa53ErXV5sxc69Cni38wD01zKaF7Xu8eaUE731W6/aKpoi9usPemZWpR
03fnA4h986imNcnsoHPv2XA5aXWGmA5EjFMWqrK2dKp30EUoH9emmf1ibBUbsdb2
yhaOAl+OPdDhV4coMvPwatglmXeaJ2ngtjLr9HACbiOGPn5ycdo6u+X7XiB/e8np
bMBf6NdLdSAuf+McE0pC6rbF0Vi+sBwQLcuRfXiEWiZdS5/RgBfJ98EjMO0iUJYX
cdWn3GCZi9Mph6ls5b1B6bTAyoX2dyubcLxBVjzqrkwf1JiBgFPi7mtMTPr46Gl7
d9kqSP61TkrRVY6Xo+kjB4M0JD8KKVdy4ZGaotZrhYYlB/lkwdFp6PcIz20Kfv26
548ggDn6qcexOwx/mlylRJkc61FAPNF6TvX7aCazUCBh2wXWZ94II906aHuYy+rI
vB3Yg8xlK729p5J/UykTABRH0DRD4UDhvKpiPe/usbGVnbeuzr2W6kXwPo//UKMY
MobXsLQVjm3CNITSMsGk6tA8pGT/N9kcF9arBq1391ZIlRWIWxqHR+PHbjLZ6u1S
Sv/DmJQoAN9xVUP4/Y4s+W9sV4yQQQGhAUUWVLYVBXL9fuhp0Te6wDHpL/TM9V0h
dU6duB7g7cRqwqpLEOvJynOs8xDjwmiNpCs6JrP0d76DvhR2ceOaEFYnFOhAHf82
ZW7VBwrAd7EQubpR1GWMohkFSefDjVW53i3r49mVEmPYK+yl/L3hduPJrETM4hlz
ZS8DRBO8cPlIOrCz2xE1qh+pSttBcpYIZL1U57XeqX3C0LE3CtNSOhM2ooYBbW8t
AEhx48aUOT2sk5pFXiJfsv/S279HLmAXV7NWTOO/jN1npGjHl1yzPQaMrSCuqP+F
8wfTmhrephcqpP0vRRGgVrdmzPgzWOCycavlIWWycBC0zyIWI8nopkAgWVrTgrsn
NPDUclUtiSuFLe005tILdicN4iRUoYdYG51PN5cFzvEj+OoFYqeYjZUtV3lUcANB
Mq8WbPSI0zJGGFknv21vi9sTxf/FdKbP0SdnplAdtkjYxPEazu53kHY5Hp68DBsV
Sq+gb1kX3Vn7DwTrGBYDvxdolGglnN80vv3AuJlozojnxASsw/t1XxH4oFUiddrZ
0RNSSV2IltKewjIbxrAJb+4HWS2UsfSmnQlSq1TpQod/6Z40PNcUsYMNs2RG882k
pEENKNZi4iO/rbGKSrfbb+KHyLzAF4VDRZTTMkypTqrVMCv9ck1jlWZajhkE7iZ7
9S/7B5t9PKHy43ZLlPnjd5B9w3V815d91RDO50OMDm6cJqOfRum/3WKIY2AKhiyt
m/Tk13WAF3AfriHFOc7jzsZ7nfridGVPq6FDOBI2soEmpgbyRmwxo4oMflRtircJ
6oHr+QKzxYyHKa7Ck/JcJWnLNZCrJYnwZbqM+yJPzvRp7oMOGzvvD9bb1MF/TRoB
AsOKlWGpAmVvDAamH4nh2kqbEmCZnbT989upSlH+u2P/rKVmD1gOcoymh6YZmYUq
g7FtV/BpfHfzC0u8DmtRJU+XGlMT3YLBQC/6rflIobuD9ZBmXL1YTBIYGYon3YFi
v4zQzZalejU2cBeEcdpr3pxTGUd3kparUzR/V9+ZZZriM5g90QhYU17AtFwFkuCz
9hSfw0IEMI9HCNzg/bX2WfKDG2HRAjUybcjT6Vi723pJyRZCxydmvOqxrlLUFWgC
fEJ+ay5Pjl98fpuV/ha59Jl+NLaTnNla4eXRxt8AhknLWoGesZ8NN+CmpA+PN2N+
nvCcX20YVyvGdWkY3XZyNfA00XeGqI1Azh50OxQ38A9m+B3blzd+MVZwonLuzAJZ
Z+c8oIbX9B0kRFtHUDVNwVsHpC01n2cYoHkdPnfGGQZDdl7Tura851G5/x4Zid7O
iWdHPfA+oU7ydWnc84ST9YTFRFzrKe463ylvp3Qnrt1CjpDNdqZ4cipUDc8OJUql
UYLXXfP4+20sxGGvHVbYW8g9aaRWSNY/p/ytl35bN/l8AaQipbhtoJi1AYSh2Q2F
VbkP7U+3PFAYoOBbcIKr9ENomvI+6nAnq5xJrn9ph3RRKmxE+GN6lrL1JnSovHYB
YJMwmbLBQInCJyoUAGPhT1F3AF8RnzYWzPNeX6kw9BpVVW+QlWYtK4jAGnHotiA9
7F860ZLcgHx4RVAxisYvJjdLaYLAILzUHUBLcd2sYF0=
`pragma protect end_protected
