// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:35:29 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
PP6J6tz491O/CI/aowcqtkeMIfNo+UsNxTfe/nEdSmGI/hdWYu4ETZgzcaq4zX6y
gkz3jfioRqlXnB5+XeahRPou2X/2hWHHz5cI6dfUtKHwoAgCWy6uuNrngRGCti3p
qol3h6PmJ1Mw63uU4ZhEY4LW6+YIW88CDm4Jx7OaaIQ=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 10416)
9g+W6CyHY9qldKJ5MUEKUKA29MRwTph4xBEDadr2CQBXAErk7tnlF3uJktbwfjJb
NZOoKg4rze6xkqBkl/V6eT929GMQjAyaj1cimOivSq7c6f25e4xqJf4TafYvT+8D
vXCoCl9qSuOBEuJ/hbra6v2FLsWn07Xa3slmXmNdLGVz8QOxynfFMRFL7LgVJ9Pf
oJrtzdgDb+srBdsi2xzqnTlyyg8uZc2Xdz/KssmIJSEFMQONPuUtJoU4z5JsbkGq
o+i9KVhRB88G1pUhBVqYaz5OgYfmLcaPFteYOWZHbXV/wArjeAYIlhPGd3DTDXz6
nKSq6CLv/PphxobWY0ieWNoxT/4H6xcmzIDtEzVVSSV5jq1P3osefG9Cqk2WH67I
kFuoRX0jECSOc0GULFn+P92trlvryfEwpj1iM0qzWluyph9iK9HQ2t1F5ZdO2sKD
k26JwZTKCUYtRQVE3CQe/qHQXiLMKuF11Kp8lEZu32VhhNhtNvnNn7raFiSDMCEZ
iDzZ1O1QEzW81QHOk18OzG77YSixweIzQfoZoLDWD4LLA63HNWyEqNK7/AMT7Osa
0et26QXy98fEqOf5RJd73gvBBRvyE8e/kK6eQwEJ86ZMoSr1NILI5CV2jWtaow1R
mpQLJHngoJ4hfc3eGoTPqeet3hbvdZl9hBWb/UOF6EtohtFIjR2aRrpcdQD9DwF1
wYgZbVKVTPoqXQZ1cmWo489A7lWytr3TE+jxvC06+xGZt7UV5wcD6lQDuPvJG1Gf
ilS47Kxr/aIKD9LddVZBR1QMP3elqKa2c+88ZJ8NApJdU9Q8l4lwrwnwu4KbbAa4
lsBf3QUN+G9DGVJRI4Z2cQHSvYg0Ewy+4eCSIq0hoWYeLuBb35aaMymV1lJYhcko
LWjHGjfJE6licpCHLYRe+ggYsEBVJeM3gVj6/41ko+vvN+GFJB+7Pg79j3GtBfad
KIijND3IrmYzyhJEpbDNrmjgnH4wJCFcVjxYZf01EIaokff3Zk/U/LDN0gT2YsfM
pQ4bVY0Z6nSE3EA52mNz3pc6zPte1d4naIaA2B9yGUcp1TJfsgQemDCZupJW+jfZ
+qxw10iJ5saVrlnn5aD4G0JdCPPDM4gnEyZIFqhZ20vE4frdo/AVKSGwGt9x4ls0
rSogxygC1vlI7axUoLiYgwhZHudFn3DDUE7ktwMBIzGOIbt3DWkYgZG0jXCE0IFQ
FdGAvIbyCvjIS+a7JOdL3iZ4xUBh4H/OAPsMJC0CGSFTz+4zK3Z8f8n6zssAZnhh
SLUgxQja3q6FWLqWW15EXtqKt2AQMAR1oHZtcVTJNt83/hULi51Oq8l6NqpLgaoW
xVYyTBi/XZHffjfTEqvqkb5URN7sbh579jPRxL2Cbuw3o8zt+YyKaxpoFExWQ2tn
HmZWeMF6v+cEWbVfowE91YTc8LAjt7Goja3KFj11ABYhCosH0PBTbJ566rIFr0hd
egR5SOg/nBrLV6BnTGYBAX57Tj9F4z09d3JBnigRpF02mG0uzHQh3E5Kza1kgx9d
1F4omA+RrR1tqs9U8VPQaMHDE0Kxkw9nNRTV2NqK2boV3WscNBXFqHOmo6JYayPr
4A95jwvcdRoJGXdhCiVK7lW8H3FP2P+cidFAawhiNOQHpqsamvMzwWE+noLc0r93
sLQq8dxYCEIsCFtUPYtlvJsI/Xhuju3/E8WiINUpF/14lI+Qlha6TVLW1jsKMpd4
suuQnhCOnG8hQAD400lE3xWMsGbbllhLB8hIKtvLX3qruHKfrqz0NVTMGtaggKBl
SPcdY8X0gNa78ei9Ci/ySJTGRtd5rkjTrxoe8XqNoKdxHE+nzeFPOpCt6XAVCniD
KOeRS4OGhncdJqlJO+zmXQGWAbAO1tzMoK+0vwZegcVk6QIYspbyDuHWEaKzGYLl
KPd+qOWLE7u7hVFY83c585Jovb5BH4BZ6G3PudJBTW0OS6CGhuCXkjUpDFdsTHJX
eo+6hnmvfS/yqeLi3RhDWtIalcXDhd/qtu1od22VK5LBKETGFgrsEYjoe66dK5lX
1i7dgvROzwAe1aYf1iUYwl0pkrmwSPGFlpxHcqpTaWiqtcn7faxNyKxoZoBkHR8u
NjnDeFOlLIOWKuQu3nR7EDg5mdl/5AeiN8nuQasADgqATCYn9v0W0Vm2VgtmA9cL
1ZuDOyPeMplEDFmcowAo/s3LN1GLm8qmHtBZcPvzUkzLIBsxY/AGG9WgnenRG1qR
yKQEZKdTMuqoNezVF8NPj+HneuebCD+aDrTIwvww7ZYXwO+kgC1lA3n5Wv97oJdl
Hu7IvGIURXDg8VF2U9ey0uKH1z/Y4lCJD6E5TigbcbQa+En2pYIVPUm5csNn/cRz
RTOiPP9kx3LGhXCWD0dTfEzqDPASgojaQ00RDoTNsyS0uEV+ltIiR+KemhmLFX6q
ugPl39NkRV0p8YXUjz5zKpVfb3LyjnIvDm6a7sXjuF6XKTyGPDkpSjE+Dh18pTR0
+Cz5dkX7rJSi4lS3H6/TLbGIo5Bom0Ropow+Lfmxq7Gz9qC0MvZLvbDC93PFB0Kr
jNgKnjWLRLc3JiOeJDbFn++sIMBWgsLskeYCVT5a+vNDQKj5r/xwxxHRpLvFlVXd
Z/VPEolDSuGW0vnvWgVkE4PmXIPl1N9mlDXmFPV0mvP0oMAgrvdmxSJ3nzh4fbuZ
BlyWiukBYta5tl4Q9m3pUiBboDnVCksPPqF0Z+7mmBcCQX5etqsz+mHmCiyPQCEu
GJHC9GMo6b+VT0RlAV+UqkV8ayAlHD3lnEU51Q/pSUT6Dgh7XPV1D6KFFxH71Fv3
S9EaJNHPpY9ntHhEA0Cf3FGWNpIxhmlKN4wum3KWGusgYwy0Ynimjbf/y3Zvc2Z0
xN88GXSNEJHaM87+HBTXHFH96EG4+BppYC3PFUuTGxuvSp7syU3sOG9Wh5PwsHHk
hJnHnMa/wgpW+9EO8XZRW6j1EU/HBR1Ifve0gOctCz1YjzDR105lS+UL6vJE9KWF
20CRr1bvIMFMu9DGLKN1JGW5B+RtDphkUnxLD3q1Kjh6pQcxPinB5m4BCYUBnucP
00TZ0vQcOLHb1W+oIEgJ/t7HXRzYZSE+CYEs/JZOTBjGugcISraaBErRfanewyEl
LoX/O1i/5szWLetBvhredVBFrD/Y5MIOWvl83q3qKIvyjmFRjpvq0KAyFG1eKL5H
MHNKgw2/O54GKgSc4m90adeWu/0+mHH2y1zL5lYuebTLfg+JGzb1gXsSu40XcoKg
+Nf+dpkGCo9RNkVnquYFhnS9rQ72XCQxM+MsAO+W++shUyc/MuYBc0o576hCwb3y
vIz2a6HLlqMbpOvbZ63NjrNB98aeUA6EhxnjjRviTs410OZyT/YiUQITlwRoJcKV
VbGyxn9HGiLxfSDaTfmSGDTuYZmZIRus672egZoQ26zeLmw2culYNup0bFS4dXC4
2HD78iTEeBy2Kr7u9GlcHx5prqdamarcD9KSShlth6P014GRqSrZfDENjFKTNaVS
CdizQ3xUS99AJKLRj+rXdr03ujANWL2/31TOsNQjOlpr7U4NyuZCOEhKgfx5oz2T
LA4iHjHbR1YgoJqM2/fhid3q4MVVHOvUFYNR2L6/OBRGEAMUbPuKQK9KAFSofTjK
0C7Z1nSy+/cBaoXM8crnsN2tDyP6LszHBZwXBuFXvwD6Am+9/ZAY1GlgYK64UF6t
k4fgRd/ei/L+jd18g9pt7hLcfv2+7uzAMQlM0yVHaXx+SAIxl2W4KFFB8F73qrBl
TDfJy5fQl/091NwYgpkKLjupWk82KWOqtE3Xvi0J19FqOqVXRPqrWVfY5XIf8F0J
pb2iAoLkUmBQzmV3mIoyQGI6Zd9nKrRfpifeVpk0AgMy3fE29VP8eNB11iqywC9a
SkfWoCKHji6PZqlkAMKJbiHC91xgEzG0gtYn550ptRgyIIXqyvbLnyp9P/hBhspf
3kzIyaHrlnDU+q/5/RhGBSlAPe8olKaaIqNu5Bts1Yt5Z4EbyD3wxcR6bLfcKQdb
pHd+uylw6K7WxUY5wQPOyvgkX+CNXe7mFBiqlVCBvW+jg7IMYgz8j7eASIXjFtEb
jaWC7w0STcX1SgEC4akph3f72ccMHz7GrUhqm4Hlgy7hXHfBTmGIw+Tw3JDEaA5A
2wVrH8e/61H/dvTrF7/TiCI5TkAoIJ2ewm0C++CJUnbTOTIKgzketfJHZX/ySkVH
SFJffO9RO6jR5T2q1pzjRodQnhjgsG3tVNiHhVHEg2vsRjokdOiSJ8dnomSWk6u+
73xwBh5UcToCVhDkAo5BrXW7O7nIsECBuRkHfs0jIiCymP1rqMiFvKcn58PK6ufI
IOLqeEN1v0IXvBH+E9ZLske0bNPv+S5VyvXEeO2DDPHQ3A0UdZw44AJsDf1ZDn5l
QBeTDlLetgRW8hy82idQHpd8r/6HBrVgolCzYHgJahFZJxqiFW9DeyQi7bunUhOF
V9tvbdbJYixxgBsDemEA2NLEJUd82qArkhlE83FsT0crZP37P7bb2EqMa2/gwuOq
oJZyJnuOJx5XxBh0q0v34QbE/UXZShazNnSXwyy2vY7eMHTTLHuCaJRV0hXNUG1z
npLHlja2NX3DgBKe+JwAA73l66+5EEo//jO8AOsLw9vlCwaMCy1FcQt7y+n1GcAK
1qNb/4Tkqdiq3wKnPG/gZYNdGCKnkehV5xQFQ4F399YOqRz+3YiMjbocMbBnQDzj
5U3JigM4VxSNAJX/G2L68EYpoO8p+SlxVnS5EXpPx+pvTCuah26Sr0rY4ulUXSOq
bXtVv3fhD/byG51sPdtZRHBsK5jGvlCFxHkGOZhv7ETq0z4iZzic4NosBNBoUnNU
83LE9TG6ooDfrB89wNnTRukufP0zsPIEZeTVfwc/h+SRF0l5wZJLXr5QCgTEqWqj
XRJVNUVkK/q0CGUbGAujrRvxUKRGOLWeYjj1CtEjmo2hJJB81DJjwGP5RI9FGeTC
7L/o8LFJi157D5qqOJPznW3Ao9nfBQmsnvzbD33nn2kd8Or2eg9So56L1rMbMkIc
5m6cFaDIZJ/bYWp2t9OhG1WnBGHSTogYGCIZ11kKMYijEQc8nXNVthFk5IapnAeT
TWDNT3CQq8DFTApTDpMGb/1r2JgpCJHidhX71dgCWfBqc6Q3V2XWzH3Yn2gJtA/y
3OCUnB3MHWdnm00xMIvzMiXOum7iLyOtidtnggf9KyyOowiIAplbHoWdrSyN8+lf
1tsj4E8mhfKHx/o3VDgG7bSU1RXC8mMZAOFsBFA0KNvEFdvjCbga/pNFCs0+bPC4
uaE0R8KCJFV8KoaWlWLsdR7dX3MY9qJStpcazLooVCUWEanP1401vWTHnv8aNdry
m8MMOEDfr+qlEsU+VNq8NEdTU9XRiMLad+a3VyP4Ka/eoooHrnGyNzJEGk8I2vRX
UkYIVRXg0AG8eK2By7ZXR7jLZ7iHnEaxgEhntbDI3teAgmu5ey461z/eFgI/KWDp
kwtuoUFox3ernm9ZRfjGHuQq6J+ypqeXTwtxS5u3TlAm1YWJxuQ7hbPPsZhqrKIU
3tWGrmueOf1O9+RIZhNa0hAqQUwt+0chYL3f6iiWTwdLLcNaEHMnART+HKyeBnZu
aiB0JfxCuTlEbJntu72zOaJBLXi7gbUlJmOQ6iydjAZTKYHBS2znVfEE8jvtSWij
2QVDymLHmN38BJJ0PTPIMcVmxjBBhPT7ETVxVo1kVm5N6ceAMZ1s09csIpkJQMEd
v/35UOGLBROm+7DqRpb0+8Dec8IMqwYg8CSL6Cd6VSA48N5vGYJtMakCkbECsLPL
5g+e2kugSAFkhKafQbvFmFpD3oH7nRdvS5ECVYV807LlEPJZw57mv9WXq+9x9/QK
sA0NByfyUX07KIfwaimludQ9TJbhiED5Mg7yv/O9A4eyZauaBmrGN+eKVSeaWMZQ
L1RxsHjvmiHiQpW7b4fWPHJ5onx1a0Q6gra7Fo92m/hQ8sKGhX+t86Et3MJ1HKjw
CvpnBo1Lxz0B1AdzCWzDmrJJEhhPA0pYrr/TJ7qJvcSTbmvRL9YoukpRiT/B7zH5
MV2M2XsuAe7Xd7Er6RnG9uK7RHZETajYLc5h3Qml5aenc7w28ECdG3E/U3CGaFah
tj0md24AMxiHdy59psnvSfHOME4m61dGR28xtK/gH3rjialuh5jTyFL3UvKkHbF+
jQYnh832orNL3fQphNy5FM8qfPr5FjEnrAkC6nVW5pHZRpum7O0AdjJ0dPKMh7W2
JJZMs0b5ADI0+Tv8/8M93nXYzqXx81pJ0BLKgnoVbkpqDqS/dp2E17Xhw5mhvt74
Qaq5Woz/qStW+q0Yjs+FL5h0aYLckLeDiC3a75BurGDnqvEEzHzFn3x+wlfKtgMS
2/5qnVqL0jCQQnct3wCL+oxUW9j+D5a8+p1gBq/GgDFQAACWHoYZ2QanYHlOhsY3
9ZhQBYQWi/6nspCuFjMH27z14/jneYtoeq7oXZrsPqqtllZu0x32u4U/m9KF0N18
+B9HZU/p/qMHvG1WQm5i6ZT+uAZ8j92kiCJmDto9UPSA3DlAU1JcfvomeMWfPVcb
mfmQ7nSzL+bHOMlI1kgR+nQsPvxhKBi+sj2d185PV/Ke0z7WssMiZSUsqqn1aq76
oQj0zbUWcqWfXCzA3j6tvzkF3kITtOsvxAg/+Y5Vvxl0DBeAlZj2f2zZAKMr7tQm
bUPNEBWPgbA5EvGXvZa+3pOBLZSpNN9DSH1tg80Kqc1mZRCusnXjGfOaNvjb40li
pr3GW5ZjXH+Q3tU7tsWU1VGar0aog96VKPOs41TuAhuO/IAvYL/K3o7Jyk9Xob+9
tYuQ46wf13t6p9EErqqWtA1vdu1AEHpLqbvmQTevNxqtXbNukxT/tpMyj0lP1mBB
s/lucGKWWVNIt9TZmw/RTaPMPd/K59jEeH4YPYjotdBHAI/wWdrxMOeuZj6dhoC5
h4ew+g7AO5keoeeVY+Rqn7jb9WB55C8Ooe6CRmYz7MWvLujNpxpIuGNNG4HXvFOp
Qndl14jLYSmu0E1ow4Zrbswc1cEmRc/9UAI0puoyTRNNb3cdFF4IgUCvY+BwoibY
Rz+bZqdBcYzdxf67W5Brwu2xTVf7x+IDvEYsxChEHeKrlm9VPSSzDoHu69b1JGgy
L5tieMrvYcXH+ieepVkcuYyTEssLDnpOdYL7na9k0wjAw98PZz23E1eAdE3GfboL
LX6Y8ZCeFFW7r9KY5HhSis+mv1+K1k8pDoqmVyHqCHVxCYDn8ajMZJyO4rE7DhLQ
Brf0oL8BUid7LcaLTnTeJ1nRmHnUDk+d205Y6SLoBqftltrtLBcdIxGxyVlL14E6
543zTyWX6TUs+hUMmeroLsTNpy11m/YJaB7lfx6jTBiY6K7K+r1Eh3j1/HGSDtZd
+TCkL7cV+XAxZbjmpSAqBu314zSiobVjHcef8WP4JinaGUsNeHFov3Kw0G5JWqVM
bk+pDsvFXVXauZIgJ/cZuHrV2i3D+txoQug31Ud1nyRtx5wixEBprVlkp6RI30Y2
CjSd96voRasasyJ6Q+kl1am74QFE6io0GzJM6XZHV96cbFX7Lgwx/+bUsyvD90nq
Wq0eqrNNx1vXBHcy68ZvvPEoM5d3Ui3D4ygjrpmoOiY8+oVqcAQI5ZO0MpXKsCzm
v4vh1ytYwxPZzxuQqpzH3doDZxOFseHGqNlrid4IQhZjIMWD6J0d2qF3A6lXFeLL
y2ubBvdWRWrT2QsFvhDnkeK3PMBrYi7VvREch+BUVN9SSNdFuVZx7fekXGYMtzv9
Y9W4lvP5LEmrsygsmIEv9Zvn4XBAZ3CfQrzBFZcI2/XCsX9bqf8aJQtxMylnwCGR
MiEiKkUg8S3+NVntSontcNJtcgWC7AeB1pl/bJgwBiNL5jT6fD3B8TglmYol0Lnz
2aHrUQPJP+XXZpv8h6DU9K0jEOBkny90uxDumHBugkelF5kmxhAGxZZnfMjqa7+E
53tOM9qJRQyMiRuSDtUEoZudx9OA15DyVvM65771BWirKxElwuuBrTHSAuWAPwu9
K+5atsQkGrMXtMJYsKCyiv8JyTjXT4pPWciqMKtFVdkZFziEY+CzPjTvVC6zGfT9
ptcJOpuJnvDByqamfAZtvaDTNZkAlvYPp7Aa5G1gdVn6Tn4UoWIwqC3zeDuqynSp
WAfoPQSy7gFToKD/4av4MHKRJhabjoCPpsJv4WP7WB8o5FAqkOw6FfdYyG4bpPp9
E0AVKzU6l8RZPPGT8qauzznzFconDWDJRHpXkPcLwWWej59piC3OtR6asGKTjp3r
dZ3M3dGZpHG24iBv3/OabIlqpee11r4mbUrdsdkOVH7bSuTBvak52vkO40haefjd
WqGkYLD7I/8oJejK6ROBAJ7/UetvenZM68hue1GaJzqfSnuIV0Ss0MoxMGzZ1whD
XwuwOdrAV+OsPCvwoi0mgncqWGSvQEL488q0+sV8MchRiDivbZrPCIiO5lz6+PYW
RwRkt01X/RwOFgJc9xFeRy32IkoTdO8wlNbbyJ6tSbw+RjDbJXfyS4SCrbyzJCOw
9w1GsqoJUI9TffgK2eYPBGxCpCKW6JBLhjuu+cHJZRbNDa1KxbSgh0QW/mWd7w6T
RHqpJoyzagWOKAF5NBDqUcrjrreHBOeLTuUNzMuKzzFXW4oTo2K7aocBXrFm0LyS
vvn3p5Yqjh49QLMn0u2xR1P5ZVbQAX+KhmcZFPFC0+o5Is8fr6CHSlIim2mTosVp
NJIFPC6QJIsEl9E9XVuSSUDDaOMQlXIZPtsatTC1cV2jprP1wtXbZwIhRSD+HgmF
gfq76Tig7nWkZUGq6x0rpCjmbh+ExXCpBNUJ6rmWTHiFmI+DmQFia/iyuRTuAkmD
ew3vVQSVEq/r3D2VSM3GlbQgxh+Yb5Fg45Blr2DmOqSYSGJqwZ8m0tD/3Fxb3JPh
JStudsHBfYZmnAoxWo+qxuyOYNulwR3OaW9e5SgKQOsZQ/xRlMuUFbN7d3xaRevc
VtkCeSRDNQgysYd/w5zDqEjPfhZpu/FJ9aj8EQYery/IZQ9oPtfvwTEAh6EAJGH4
LFDXgUvwSlxqUpxMQAQew1I1+c47jsi1i7C2jONmN1aQWZqm1Lz8cjr/nt1Nb0iS
nwWuwc/XyKnlryyeKLnTQOHUnVJJOoj3vBGcE6bby1L8HLVpIhlCuSNqKqOz4KaS
fafPZgys2DmoUJZd9exBPOjujm5UoGkFPEIFyB6EJLxU6xN6bh5wonCkTUQl9vh9
2WIjvd2NFFkRh1cH9DuYIP19xSGFyr9CaKlV2V/+8V0QuMS1uDgUFrHZIIi8phg0
CDJ0vmuTdDN/C9lnlitQHXFcxuTtDYnfVtldmtikFMaugv7I4Or2ru2TqzGhd2zH
Cbq79J3uN/vCV7ABWciL14lTNLr3r6Vw7jTj9o4dgsYJQerhnIAFZorryCVhgFOl
8MEtpVn1NqqFsFkZcO9GXVeFRMMTRyuY7hUr0crDBjANQbJJFwxvLn/CG35P6Htd
LkvXwjCUDx/UcsfHJ0ssIdijmeinoS3ThiDMfsGgHRAt9Z0YTKtRj46/XHbOcJPQ
JrNiQ/EXz7Oxv57HjlN9kOs/KDpKeJlSHcxLFf4C4foqsvgkxU7WvMxZvjusF3pj
J3fGeFJ3Qw50m972HjglDWmxL2Ia413+Nz/fjIFyf4zmrs3Fhmfwk6Yt6+aZHoAz
erpMfpypsioJnSFmGOAOJoosbiU6PbNCYr2WnZaaxFzCuUeOCEKNehBwbixnSOxa
2uP6nATgHFpeXwqXPIMGBA20HV7hwDGGkx32deM9eSO8OmjEod3PKfDTStwLk3hN
hXyfFUetLpHjdgJNo5khm9m17N5wCIgT0L+n1GBXLTWrKCq5/g2Tvvvq3BDu004H
U23A/D0xm3hXxVj99q0Zsc8o5hOO5O1ov8PTnGKKLVFSj5G+OCYNeVh7jLTs44v1
8AaTwuMoPRDO7Ic/S46xWo3gzsbpWZLYXKHQ6w7pku3IMpoouWX6lFNIopccMVkW
U1b0YtL9GnfPOI3ud8PL8KHufEmpQzRUwFmbCLMtDNF2vAjm/pRj8h1CQentYpaQ
LEEONfp4Lbdwg3LfzKDJguVfdngyGmToZ6IK7Q3bNluG4n6qXZz+bu+c1IgFoAnP
qYTwAVN7K3AWpR58XGkSs3nsQVBdBVlcoovnYsPmncyLaMdc35cw0QkBAAjyzZ5X
Q6bejxP31M0YGPJU3RDiALq9dCdCkSv92bJbBbtqXu3M1r/LSTeFC9G2rTmmB8jU
KBjjp0yM2eSygGHihtawXijpCQxSHAFsD14m5We6X8XSiV9XOkBuaLgw0uhHtViy
mmIJy7uTSlRU7NuMDXCjBaO4gEwNWqJoPZoxjZ20BuDw/dxCtPh2FDdRlphdn+tb
0wfHq29nhvOq23KlcRFCqmqyjFlikddWYd1g7CzkKTlxuYAJKglrTmYFtiFJ6/pH
VI5hgSWVQ7ZRmTtcMVQj/+EyOV3Mmt3ZlAxgLH1+e7v1yG0pe41m0psXY0gqOdt+
24D+ausY/S1OBt0Su2kfhZ6euSN2ikBm3VzOWYFsjgkWAXiC5avvAL5kxxIaFbMi
KwOVT7Mt6Z8eUWxtLnBPBbvj3X+u7Jz4J1qSEXbS7OR2ICzGtxgYYGqDoNmfnQMb
l9Abgu9T0mSf+3PBJmm3R2jSc3nC37sYS2S6JIe2mx7ZPeAQD/YlAxPqJxVz39MO
3tKL8YCOBQXo9/6vSrnX5kQq0/21DqzNuQMdnDGkFlPhXaHRsapIDF1Sp13hKZVE
aLBaJEIoP4sWu8ALLtXVQpvmgCT41RtRXPzzg18KGWz5x8E1XuPjQeHWxjhbg/Ty
3oF8uB7Le7EdbELIfKTbycKwlloGsV7C1ndB6dgrkFm+Fk01b1xncOcyZSCwowc3
K/51e9eNYG5alIuBmo0lap2i7sV7+2QJ1XTAG5SjIlrv2BC9WJBejBTon7CnaF+s
lmHCZysPOgyPEx/HlaOJYhMh3IFIKS51UETQBJZW4zV7t9WsnLK3zJnPXHYODjE4
po3+JjY7e7UFMLcvlQSTmGBl83qpRUEq0fZmi8kDrtYMqVFtybbY8/bFIXVeCn9y
zuvrZTZOtaPCJmMJX/cqNu57numH8Up9tMAfRIbypr9XPRZG/xuGzi0cZ63m4cP+
iDBHc6mv5e6gFnTQ6i4rxwOvWYiPHhKUucfxoy19idyawb2heTq/YflKStCq0H1q
0lYqEAShZJzMsmyy0250ekUlUG5QWnMvPWl4jJ3gPxAutXN5DOP3mlRkIoSsel1n
LV+7KWJdXJtxP0Tj4dfp8bFJ76WAKBrgUMbYhqX58nTzpmpRCYY50YdNjbR4Lh/8
jrdN8LNNd+m7G8CGx/0xg7YJL/wK34uNlYb9wdxrAUWqUXpDFKwLPYgesNhr5dd0
RTlDp4s7/POn+Rl4iESZ97jhCHXsTtCXqQyfiKCtkNExN4Y1aULi6/rSVCmpZKfW
PWcY0BHz0urHeBJd0hO1RC8PPQruEc6HdnXAG+1bZ+kdvv2ynDKTnYWnqdldKCMY
5fAdpQvAZy4tmwgJmvENEx5AxxaNaDKy4M5NA8OkXrl9u2Fjyu/bxtiEbRgdYYso
SocC2TzR337RY7SAJvyPBEvBDAdXeuz4iLrCVVbKZ+/1Xy9cQ7cmy7gEmnohibBf
Z0ysD87kulB6TO8yjrSNZgF5qFfHdKJ8K30u6eIW7Cm907GEBEpzxQPifT1jUzr8
f94BuWZZG6Vu9b3Vs5kbkJ/D66m+/N7hcuom2NtTMpRy36i/zo4Z2Tv39xSZjNZX
gDGthY1b13Dv5/D81CEkeyKeNyQLq2im/xftJV8FmwfFW+oMb/pmjHt//FaIJFDd
Z1esFxtGP/tmaEEXxbHnWZWuCl1Ce6PXlzU3p46dVPMMC/zlGvcor2tSVSRMJvKr
xfOeFNarinBd2HkJ83pUz7eDz7FDLyERjHyEdSrgR0ICGpJTdwds7gnTgG4c2xT5
MvU5bTG2eum+RanfmFWE/rsOb1UzTOknoSHSGo5X6yf3jvMwu7hA5siueTeNnCB1
BtEnkdagu4mro181NeDsEFqeBCBqVfWCDQFzuWUrfqjmzzVARsD2gv4LkzozavAS
+29nd9Ubp5QijrOR2Ux9S3QbvT1jrz97bi2uu2B+FN99ehuyeXjxVqkzPqZ1TmPp
Mqd/APSW4d5cD2zS+Mbwq6iCBk/Jpl8OJSzsNGeDuT0d76Ld+TnT3V9Q5Lgzxbbx
7FjfLWj5hJS8ClGDq7t+VI8BW8Em+lEE3GyP9M73K+Hqnxa7fbCJ9sx/YH4Ypi8q
3Lku58LDqxSp/SmAwtUgD1I7g6wnv2q0EsS/zvWVfIafgxYdLgDiO0UsdmxgYVtl
rr8nY3ypmkxa5Mh1HsmhCvXOQQByjBQABbI/kn1hTe546yKhCo0rhos4K4pJ358C
OFNpiiSzyy4dR742yI4A04k+4r6P5m9GLYioT+mm0mwi9lpebwq1P+EnBxGMJ/de
yxgEe+gLMn5H5w3/4LrzJFeZtUvNG3IaSXNeDB4UNveAJEYnz6bbTUaPDJ0bNEK/
yogaIDKnNt3O+2jFlCjDhPhBD6lUv4O2juT/DMV8s2vpNhx66YgrWYY0XI17eMrI
ipLbKYQJlDyHsWgnBhvvuC3kUofYkeZ12V4X6x8INfTx5GhYJN2RZaasjuoCNHbc
DlOWNMdvF1T2Y1VHdDD+mQpa0YU+4rEi5B6xr0fBtdB7nPnuIT98NLNTHC/zRM9z
NC1uGKY8+aIyY1ReuZu+AMKKJ6riV21fpcTmvpALkt75m64NYt3k1GhoxrdjFArM
ndS2f76hGvO5ymKnMIH0fxWxprDUPt0+3HD8wt8qZRiFCUG7vDcuhELYAIk3mpz2
o99E616n28VGl3b0ZaEZVCmGXgjRB4BPABCP19LGiO31hRs0vhJWtPcsvFt6Y9Zy
+lrBaMdsefG0ShlW+KZDyh1B+OuwPYhlP4FTsiUNMwfB1oX4xWpmlx4/uQRGGJQD
1pFDHevwvIy9la3Z75dPBkYtA+4QtbTe8EeCRDRAPtrl/0q59Tvs5yTlq0mxv7cz
tlLLDo37o3ExD74/3132+hgFRbYVIBqZpIiR8sxvV8CKOqzg1UDALrMquD7gcxAN
XtGoxC7uBYTFl+0oO8I6nJiSi4Us0DjxE/8CiuKX4qDFZDyZGQoam3EWh/5XRpCS
b53qAAl5VbZQFhY0lfqIlQFjcFb6HY3drxlXZysL03MOMNY9FpSPB4w0E0YATakR
ic2lCXe+cgi7p9sD7+5pMLmUrnQw1I0OqXdGu1noAFo3p1/OmYhLXHWAk+gKOV2a
R882GdelgCufuZgibRf3JThQjnfgQPYGgTTLfdMM7JtvXDSlcTiwMkEtUeEYCY6P
/nBx5mmP/weYjKPIYQqBNl0I+zyWjl+F07LRhQRphc1aqq1gMAA/ikGlIuCNs0W7
+ckZgJDOwVEafLY3T7TRmbuWh4wcEphJLoGbErVoHiV+8k26SGjPhylEfXWLjd+c
MqfDu8giNrbLZsCoTKdrbW6g7hSZ2uq/3w0+0AqB0zoXweeuVpdmS21XGAOOyfWc
8yC4t7eDDS2vSYnJ6Eugi/tReeUxE9LUO/e+Xv7AsjvoYtYRk6EbFbIZnw5mNB6A
vc5RZ4usVqTBvRJ/muTPh0cirSz7JThjYWEtLYPwz5Y0RI1hv1xdZ2cJ7+J0u8sJ
6S7fzI2eVRQNc9kSzWgM5ddon32ObawTq9JM8dDRvmYuqqhOqleSE3a/De6l4zSZ
k/UpkNnvYne1aIOCqlNm4kWc8BSBbwd1PAV/MrEEiRXg4IJ7FVL+YzGq3M5R462U
`pragma protect end_protected
