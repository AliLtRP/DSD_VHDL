// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:35:47 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
GbE4Zl7Yu+jZrk2Dv8+iUgmzPFsLCvBsAgvd63EY9H4qEQDemk+RvcjUliJcG9YB
dQIfSRSDUhlTqeRzRJ+bidgPtdenTrto7uk4RRyvJ1HqL0IxIxRiQkZ9FcEl2b45
aDzXBvJFVg5afVk1BnfWX517lPfBTr+UvCrxSE6YBVo=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 2448)
GUc7EgxuvoJNnO3PAu8RNIW1Xl8Ab3WrhwcYTaT02JtmTBlZRS5NY+qHDeoXGRaJ
gWIvRYgjKgjntFBvha4fDfKQ+o7CoCe3vjr2KwcycQilRIlBb+xEAG82aW49IZVM
FfyvynNPBMhXGvsk0uglN62TF9JDw+ST6b67HEHnmcoDIcyI9O2jy+ICuaHMz6gH
Tw6e+MaJxdTvL3QLzze8m8fqksJIi3/v9/5TVZNgix373Z3cz1dhFX0q0xOMKy83
16IyNtpqMfkKNPRt+xRZjnmQoyzOb9unZfqz/CrnpStBuja9S2at+6IX94beSTmv
GeWRH6DdVOZOs98lDPDgKoJUAcrVgV3rAUdB2kkuRhSslMwB3T9X//Ll8zODq+OZ
y3yS0Zv93ul4OCd8mzYYI+FdR1bPS9AdJszmxW3ITmmlWvq7S1mLajnxyCbDtt2G
1wA46xXpTuvA/y0yoCQd2k/O6hyerChTwNr3tI5vafgOkEHbp1zjPaHJ9bI8OoAF
9kxg/7oHRu8GtISlyrr8Be6KsfiS28UMJ6wYMYyMwCmAp7kuK/BeuJCQDcHSJ0sH
LZlsYqpFBFGBjfBzfa5dYyUngcW1w8isCZ7j1K2lauvNKIX5cclglftEmUj54Lj2
HncRcWM+vBXIdiVk5sWoiBzDw4nGzKJv4C2FOYOwtRPHd2w8Tx4lhBgMk4JRnywV
cdkmTOnQY8ZZeHki+/VgRBoUJFIuwnHGm0XCp2oEtraNYhx5can2zr7TSTaRyFos
W29tVnxPuxNSK51hgB9feTPBNnol7Mx4jwsnKiXYEAl675JFdHF9GHoWNzPDS98G
+7wX1e5qt+3dWLKrBfkJY6ePB3+u7GCMsPYb0qPt64jvGbH5IJCcrHpURRBqujCR
LqvQZMz6lPTdJhCq+kg7uzR1Bk+PkQtTkRE2gIcTl/xNJgicxS/MFkDUeCIe3Edi
eG4m//JcxO1OU7w1PD3C97AlDj+FAbJHIIMLrHubvRD82b3FXcc6treIsHfK0pCz
gv+lIPjtBNsoYxcmPJ5J2n4YS9+4eRBBPzZVr5Ye+jlufSrtb9RC11F8fPNY/yDs
a/f3yoT0d+EDCO4cH6mHQ8WnurpvK4fBivDVrIxxj8GO0YE0AM84TGieCVi2opTp
J0vhx349AuWDs+9yvpBUUSmyyfzi9PPtWlIch4+RyvsxUv2/mAhgKEUV7VvEOzG8
bwH6PVjxWdZRCAjI8j0tbLxgQcqTby3+YX6N04i6XI0GsKhD7B4E8L+PRtWSFZYu
2Q3Sd1aDYk9XMpDu+zdsTKr8kUjeq/VaO4NrcW+Gzz5m2O3RaaLD93rVljVoZACr
l8jfkdfNBUP5iQeYFXvxBLq+cjd8ngCd6feS//i/7uxUAPPUoOIeTBKN2NjdvsAU
v2oKmnLrb+DiL4EBFFckeuFtYVnN18olWHdlAYnIfW9Vgucu0A4CKa35iMuyagCs
vHEvfqMiQJUuU4Aot1U/20hYv7KmXU+tO0uIJcxL88XJwaLQpr1Zsj57eudXIczP
u/GeFVinLkdOQhfCwRqmP5uHxIOjIFBEjja6NgbCBvkfYkzfnyhiNADnDnbGfFYg
avRoCNPT25jkq3nZr3xGsIOScCXx+uObaSG9idiUDEXVrMWfV6wHKH1O2GVnVqPb
LwDbiTFxNJeNFqNi5GcaCF9WRMJc+a75fyS3iqCikbhMZtHnrTWclrV4UrXvlL2D
a/nT3z0bzEM3nYiFy0Cce4wUtsV/RB+GyMIGSar0k2XcgTxXGnMVyrauWc+Vd78b
v/KGhCvwwV66UYqi2p47UfN+W2774AmsCpjQNwC/xnreWQoTKyvGkWEnqnQy3VBk
k6LezWfhfMRJtiYqD2NwWPX+pr6w5RgQ941EAzcVNgvgMnedsSySQq07VlrLMXIQ
nOK7Gpm/0/LgAHWJorNCKyMy3vhVxWtUbS6FYME5+rFmRJO9Zrd1mpziCBX+AEwE
EWCYkeojxGLijYpkzwAJjYqwQqs/98GpOZdVwqMsPs0Vxn1YDUzyU/LhFJsutiix
xrplj4Mt7GNhSGfj1oS61VtGe6YP3c0oxvIr+PbFKSQZNRjwS7n+d2CXuHA2Xos7
YVWmeOwhYxzgTjfQva4rW2WJUdLaP7pPeQBY0rY3H4ocDJs5f0vQhldzIPaNUWdQ
zZm1wqXAKGfamg3NQKnBuiPQvS6jGzC8intCWg668X3Ah8p5+BtBUV1E9nj0dkSV
Sd0qsxt4CkIXyA+DnduEEoIe5bXXeoozUcklcsfm+uzLdc2jxoEstEAh0dUEpC4J
b1ahoEtC7DxX6A/EMFouGpD0FU7/SbuX11R5G6cgI11jGnUOYJBcFiJR/YBIJqsF
VoLasjenULbVnX0IN0oOHWuIfKxf9qR6Ovcd30beX5At7kNZy2kv5VLbUBRFPRDB
cnIwQ5P4jexG7FX3wQ9uviK7d95eCRNCt2clTh0GM806d+BnXtZHOM4b+DOlDuwi
ivWllbYdKoBnMEkproFCB1cPx1tqGLqz/ttnmA9eZO7k98rdQj+i1EExlXmXV74I
tpnpyX/KaQXTHFWDm8+cEI2CTX98MZTvnVmV20TQcz/xcJ1Ro7mNNWYclXe6HiFl
6AH44m/UQ1dSCKc7hPflIm5luYXsd8Ln0MZDktHrTajHqM+VMzpmeHNCnrA6nag7
X8ccwZCLECtqw93C08z5vj29IDKqY1l/bAp7AntxzIsfsBk9lNKG/+VqVaIxrxwR
QZtbnAXQKeUFUehgJejyh0KCVT+jUFh2+Wg0eIHyVoEeXCTsrNULy5wNsvBj0Orw
m8I/M4m9Ult6BQk71H+kHf2YZDon3A3gU5BjPigEFThAp+T9L4WBlcseH6XsPCKP
y7HSTL9hr52BfdXkKkGqxbNvgbtaYybDCeOYrzkjJfOIlL2qSiNRh+hszKKoU8Ht
y3cV53tj9Uj4E+4FRhWLlask2Jlp93t53A+Bwuph/2QWbVXLqR5N7J0GoVvzfMu7
QlmRHGZmZhSlvbliDqFnIXnXAoS7lkwbnB1W6m6s+bL363DzFrxsvdE8TYvif4sD
v4WhE8jz/XB3jElC28a8IBsoqeQp3GHsRJHpn/udVYdFL5TWrrLWasAvdmQFhLzM
6Jln12cnBsNO/Hqy0kjUPPM9HJtTYBRwMUEnTOpQhSOGCQzoG9KP0tS9CsrzjPBL
b8s4vwBu0yorOwR3NBTndfqv0N6Nq/yFMujcj2iRAr2mUGZtcIzur8ib03vyTkbt
`pragma protect end_protected
