// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:30 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
eW1QW/mDDrT+WfVYVpM6lT7/0jMKl49M6sShQEmbNhjbVYvDvGkLsnVISt5vzZI9
eS5ySZ84vZnM1t7aJelu/06HyxdULavjaB0z/Bn1nhyXC0YiHkAHEm/iegUYH4Zv
Z2G2/GCWrqHlEqNamKPPskAkduuUDKSFT8rwjbe7acs=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 2896)
JPr3Z+J35vxsj9CNbwtMYoLUG9xLkh8Yp94JyeXduUPCDngUx9SuZBCPbuZ8CqBv
2WV8XmVCtdtIaW4UoOjWups7L8RlqD18bXoFQ8rdVkJxRlMea8Zi251qqItNiIw3
GEPItaDPloVm1evZ1FXR7zroGG80QXJ6TYQabLiIRMkQLYsu6qUgA61MtBmIDOPc
lhO0/RBzUV4atVpUHUicpqG1DaLM8mZSW6P+xlILCbhE/p62FBso8ES3eQ2G6Z7G
bVA2whsKKVC9aRRRdDVVHhJuCoDhidVXZ6F0uTVWZX6KP7aMu9nZrhkbSwhdHcvx
si133++c46dnmhWS3PhZHNu15Pgrq3EWtvJ+RtOIpKvYkpr/XNpJDvgOrlwP1daL
1r+uxwpSG+Xh5UD0NiYpJEU20Q3aI6etpHaNsUQwncjnKV3sWzHbGFaLv+/vEUx1
UGyDDKv/0UMxbgiOrb/lTepSApp6t0KfIFFiGfCd2mV8zBnJQW5Ha5L9vMetEHcm
7tOl4fpF492Vr8Tfop+yjcv4k8r+0yzP1qUdNY/sxEBHzI5p6c+RKhNv6GFsDdin
VuNkWPA02DH6WFbU1yzp2Y918KTiH3bbQp59C9825b644EN0cJacehu8OAW3JVDW
gF+4+bFgQmIfjk27YWnmalwdorb3mewvxcAsYCrO2TcxDpUDY2Dyxlm2+sAv6t8V
AHQ2j6zxE35Bds3pwO3yRdiciOFOozkA37Rmx8Q834PTDvs7bpx1NBNcop7mE6/b
yXI3gwwlsnviQKiXH4LqAomS1DS3zS6z08nrIBL5YlzzHJ3OZTu3XsTVPJI4+3vM
vjkmn/re41LgZl/7z6cGMRSAIygYioe3gNtNX8gwzDSrlMg3Xip5KcM/BCNTQ0BL
+4vgMZe8U6SyZLFFLDOgKMAREkYYU6MK2I/b4UCN5lvxogCcLjWKsRIy5OOfzR38
GWwxMi3RtPqjd0heBjenZqvjM8vVS8o5+HDDWe8TygFRV2pjbP3kB1XRRQrQOhP7
oOrxk1GSw8xO+OqF7R8DyzgKGzQFHGdAvgEmllR/++ZToI/DjxYGOtIYTreIdgTL
Hahx9u1NAyeklUwHa1sJ1lXIQWPRSM633RiNOBup0Nik5ZnRWfhHcPErkWuNpwA7
5DyHdIjxugJfZAxQ+Ays9AiGBS3ZlXwNyC+tVm12WTTXLTJqP51xN//pI0xkHL3E
lvG0TRFKx2SIo7wktr1pJhFp35zywyhCe/mkDWxjcNlDDGahT2Ph7iD7d9ah1HXM
d+H0Nsw5GgVhDLwun505/gX87+whp1kPi/IllYn82ePSZyQm+8p3sUrxpC/EIbHq
GyQbVcnDE1S9hirXqdt3v+jmPL0Sl+cdd6550Rswt5nOQGQDlWPaYqvT2cg+J0w7
GeLVicjpOtHrg3u5YB6vwi9OtILdzMzZNtlepfoGCljyZ+NVRML98pclANDezkxS
6/pgrx8p4I2Ou7UmD+/MRt4XpDUvC8DbrwCrZ5cj1yL9NuDkWGxZ3/0i7JvvIfE8
vE9vEVoEl4uZVlz9Hu/7EwIMs4a5jokuOGb7G+pxbmCkqPgQArU5Xl+PGyJ6/Vfg
KM8k9/qjapPIhRT56gyjmg4Eww4zvBtdUpQxNFgG/0hwyR8ZZpfrA+sS07SEy6t9
e7UuoWoDYv3BkgEaKyydRLiYKObu/8PisWAMobNXc9Inu2b1RB+NwN1SFZT6bWcP
qBwbGFo96FL55p1i6O9vg4vwbctN0xKmQ/qDkk90ThwyAMaie2QW0qYeObIv/tuj
7Jtal2xeKg56dos60j+3anTTOzI6z970vr2/Vvu/NVENY0iSNiNZeZ3/3MpXyAbw
Bje1hcfjkYuwr2E3UnS6ReFzX9uNNjOqY8gZMXV0X8GsKOVCZUjNlTls7weiqunD
huykw9gEUkySu+A477SCMLqhwW8P3dXnswpypAy8iHREddpzdLr0x2KhBOW/6xwd
LS1hUQMbRLaIfrVzghvixcjNtN6ejc3oBnmaFlSxvdHuBjCdAALXieXezbBUaRA0
NzOsUKNmsRZk05td7BIyBGa4U7JnAiz/e7p9xb639L5+ByvkU69sVEnQE2F6pr81
87yhZMc45N4pb8HCtq/p+nCRLDHDFx8Ni10niKuxkkm+Af3ABPrwb328xi9xKmvl
Li7bLz57YyyCu8jLdT4M1GRCOKjZWbk9FOioQlUI5IzDY5aoCq4676JHqKmdX0wf
lOCa77ZFne1TQIgIWCdVqonQYg2yJiKbNQj4FkOQSCbysLsmUP+TA4kqZBJgBIka
yytr+vAty3nzM7R1NML4YoxyN/wDk7nCC/Qt6eUitucUlKA4N4JQoCG7CbRWF56O
pR22RlcEa5kBY+INbjC6IwpV1LHahfv4ZgFXXgclb6PgKtR6ZZPd4y3kCgzQUDnX
yeg/KSJ1XzHw3LRFLnZl3N2jq9dvnO4MBw/nu39yZGKRQvy9rHw6rxAs9Mwofwve
bea1c3Pt0oxgyXTcrBHpeBnie0xEKyh6C/bcHnUESHTK1FzBMGJnQCogRNujldNU
sEsgaJHFhVh3gRwPyAK2g+1BuQIU2fbJCIHYUALacdXNOYB3pAyeFzUoqR7kajjE
ZhbR4jC+Ji/kNUjKwTAq0uH1sexnK6mwQFvGD3AbiQMphlPmT9KFT42z2OlfSB59
cKSIw0oSxP7DAGqqAtpE2kDVcol7aZO/zkD+ofpOCuY2UujoZHIBO6tRlZIFFs03
ImVtBDfePD1aeAZ5fRCNRL4VLJyqKGSMxH5yxkGCADJ0Xqefp/mikuO54prkYTgA
STHxSgVrB0JLMb3rXIVooBm216D0DfwBzTzXIKZDW0Pp3m+iq3GSBxaXuPYuJrWG
LPaALdwwUwVJvh6RFr3d9VFaZY6zgYSGNv1PRZ2tiRao+iDyoIDqHZ6LhDP/OuMK
BjJdC9URnNbrWPUEM1k85rDe+EFUrFsviYk5V+cgr0IYf681EfDkhUwcx3XZ9Eon
4gq4XFIGN4gddvbmoj4G2eKwnk0wTBTKNEEoukP8TjPHo2pUp+yC39Jnwb0cI+iH
olM2VKGo7S95qvS4mnkJtgsc81tpUCHphvFhggDY2PL38piONKEGq7yg/2L3TL9a
Ps5cn8AIBKP1IrnrO7Av9dKQw3vejfVG6bddGbIJLrtHVKQ4VNRUYyWkm3ySZJSM
FRuonQgI1QqaIZrzWbE+Av1AiCc+gVeqdyhzkVY8PBFskFJEQJfCnxVDsZDsnAFM
e7cDOSZGQqDFeCf2haHYnPHU0J6U24GM2pz4H30HDjOcfUpTDzyhGKpkpctuJeVi
4pVmQHniX5pI7PJcwZ+lU0pdJ+Od9pD/O08BAMuQmxmu0MpJTsJRhlN1bhsHPgxF
PulmzupJXWMq8LA71fSpZMbbDfPvKIg/kmBOoqSmQE+XyXhnjEomyJLFMJQ21jHY
hndsig3OhehWZGg48L0GYTBB8oar/+T1BLQgk5l20pQpccpDOaL/wxwJF3DN+fPV
6E2iXZKxwXiF/uM8P5nPD+2Gy6Ec2vMIJSTC/Kl/NQ1IxSKPSgpcXHxWTnGH3rJ+
tGCEVQGAZbskPbPshMMBtPfRAJfQPxAE5Vbhq9ECw2B7V9U8B0fpDfX97XXRL42U
NMuaoSn2vksCBlBZBjKX0gSPtrM/F1SnsjEKtYV8Vs3U1R91kb/V9ijpO9SpiIU2
+wFdauHV2qXuCaVpkHwYTNpRMkhST8bfmozSfGWuCHdddvi5CQifZs1LOXCh7O6y
vVARWgZP6MQ/2hpzB6umTdWDWSR2M4uZ2wq83dA0ZWgb6KPJUMTmkFhdgXHSaXLB
QnXTAcreH/sNqVcPL8x6fw==
`pragma protect end_protected
