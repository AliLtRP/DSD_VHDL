// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:25 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
rMzsWRcDzanOxcW15bIWjEDovxDJUShKiDCQ8puKvy9D0ijygdJYXEAdo69rFZ4M
Uhuzp5mDivz7RrOcXMFl3G4DLdmJoCMZC3AbU0EyqxtGVNKIbrjuB1AsI/CTc9iq
d5vxyvcEBIQShlPvqDM8OGBnUpg9UkD76aibU4zB6LU=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 25024)
FBreHMSIZh8OeUH6h0pUmDfG0qa549ddSsSoMrPZKUWYIK/4dyOQi34Xa8Wka06A
vBHO8lc6RNYzfj3JiNQ7Y94naoigZSanKgrnDQ0YyZO8lsRcGNzAIMCo0e3DwDJd
w+lIY8FXA+N5+iMinRQ7y1JqU+B8UM93P9sPLsF2ISLCp4NrZ59DKi8J58YCItI6
R1c4YDLPTs70L0DYIM843gYnDiwj6OgBKtKlS0Z7sVNE8/pAOE8wUihQmUGn0kLZ
AsOiUrJFNnak1gYlrK+45YabgzsPLaSkL13eMkHkXhk3eCJabK+Zh4vC0oLw9T3Q
VqzLB1sqQmKjG8PuY2VP+dg46Oof35Efm7sNv468vjOcbMZw7SbB2ejr4fXFYnI8
37X960to8Zw9YqWqKsF8/aK5C/LHEsP9NyOJPy2wfIXYMYCy+ULghee6OqDb/tJ9
V2vX6LXf/lQczkTPXLRWW/csO/O3rS6SRzuLWdtIWkgpBp6OvNEmoqXPzquTed5J
vxbdGSy+15uY93EFvrsxy0P0CViQJHVoHuWgSrrFDZ0wGqUxVq8WIIvfgW1NQVLC
iQM89Lrfb+l8dFVncmaNvdF+snpmkIDCnfoOL4YfcMrlbUCzHrv5miWXKbAmo/Bs
0QUr1ho9dFOlXXqDvEylroOSgNme8zXVKgZHKiLobMDK7xA7ukMe3vdmlmVvHNzS
B+Yd1aiqXZPdMpBEx7vxTfAjZntng2O1SYFKKoJ8+JcefU2eRV6zBbveVq0ulJ69
BcUnlCLVaDzF1elTHQ4qrw+HGA4Dc+W1e+J/uPndMVpOZVEhOORWgvDugygBxaU0
81zq2yjiIpIFc8Ubu/O7q4RgWFpMyXAgKSgomFfZWnqJp2Q2CPVo3espOdegIRAj
ylGx13yS6caH6my/I0SF1ys63NAR8Xtq473B9W7+sPcTDfy89iYBsA3KnY4xUBqO
uUZQRypHaJMD9dCK2qtDp9e9LW4goAqgV2JYl8OZdJY2zq3hFt6TrpV/0Y9Nez6S
6TTMmHJ1Rmv6mKLK33tRZUW3ayDf8SkGF0Aa6IcESCJyeVT/ajIO4jxkqQMIE5Ul
44yZZmRcfaiR4WXvBV017fsIoRaNL/xYjhMvNdVEXN1jABqEDYdVaJ1GYD6fJ+E5
IhRh/6c+R8IaSpERZ3n7blioI+KG9hIpDbvRGhFGFL3bf8xRfHcpTDc9dkP3NFgd
VcqrznpYqYYMBLeLbWKmS52fZnkftumDG4Nelc/y2rKIrFc2is0kqwbD5d1xkfi/
IuQfO658Z68Dk+EmkwVa4YeAH8mmRKG4Trbf0UG9VHcEGBAfkqcbd6Wmjqz0Nf1I
TBkMiy7PqlEr70oODR+o07uhQPRFLOrcTLSkhrhy8UFxO0WUs5pBCiSlWGilAErn
9alp2+XY2rSmUWcItOBiTbck6cBc1BKP5q74SQZiZXREJFJGwFgZCjPvXUz4Op6m
hbetSQIny623ufruQ4hkXI2HffdxZ3O5CljwCI75FsU1977eZ1tJlNsj/eQ4j1A7
PoP0MBJPPakD77p4qWduK3nyNpfLOSpNQqyjoMtlLASiG8jCQhpVxMp901G+48mM
QXw23pVa69AiP220haYJP5TvSGytnUx73dYHmq+H/xeTarDV+VNgTATvU9RbgswI
Rrl2iDDXLnbb6KanAlFcsU2wNvJiXNLA5/zCdQnGpI7dkrz61xz2fu8P3I7wx7H4
Xm3Sm8lk9jOV6YLdHdvTqUg1Xtiuefah4eKBP4upFbJqdxLDPRxTlj//kKxKlAwS
U1b5ZHUDWLffNikxEQHhTPbSqjfeGegQrljamZ2ZJR0F9/iKwBKo52ZmNVX5sTRP
f8xdMz5NR1xUkhba5wZx1Kz4oFiIN8mlEd/e+7GGaEx9opyAAsE/C0xDPfT51l0M
tjnRNrsWhzmLn8chMjrmHVDTdLaeftaYsiOiGWPHbVBrK/d0Nbam7gtIk+4nVYqs
sJ8/h6oLyPhdgDm4mGXVc1QQK7xQjGaWx+70aY+bcE2cwh5BdyEtkYasLdqP/95E
xrUr+5IrEb4jfkRZHEO3ay5+YAJTXiZgQrvPzjQPZilNmY+9NprfVWdNMzgq3jpz
Q9cC3ESQ7ktEmUgHSxx+TOzDeUfGewW/ujv+TONg3z+doCuI+0mEwxKLCToew8P6
tLa+BNFpfU6uCETbBWy/U1J4XQBIBfMJBcYFmEYCdfTkwNKCJ3Ru60QEmoAfMQuH
qVwv+dgEpYhiHtdgNQIiL3Tl92OIvHisxSWxCPRkbz610GFgz85zZtvTscwxCo7d
P+lJ1S971vfwB5nCCCKYSuppOaFUR4hckwq8Tr9gsNaF0GMwYtyP9YdZUFWloDau
qN7bS1TmJlQvJPb+XH4PPovCmt93d2NCt6LdnuC/VId5OnygEMd1CmQXVI7qE14A
irPSBh5G7ZUQn/1yRTzJUUYFZPINyDW2G0oE/AN5+sSqv85uE19Pqg98lB+YyOhx
ay09XsNOpKxRM2+UPn56HnGf+DckV9Q+Fxc/gksFYGDAF7TI3lNDtstMqUgSkrkj
aKzm/hR+pKep0aeF+x6GIp1RihCe35z9SsmQyG1UTv7h0RParX9tX72HC5dWJDQQ
s3D0CjT3Kw8/nYyjvINS+X8kBxHTG0fHib5KusFdFUa6OY3mvhSBKb4o88crKC3Q
Q6zQgGp3Txt/jS//aGKGnzEImONfMKThIhQiKILoLyzaibQTbGJKRQOFEQwTHhKk
cSeDiynkXbbNCjzy9n95g5hNHEytoGEOywy72I8QrhOJfepGU/FolA5juJiatiFZ
BGH7A4D7BS+kPv3u3+xxE6ghkoIHRutV8sRRPbYkgvpzhU/skO3iPPzKvH4RLbsM
8EEuUv+i42lNPkup6V5h9Geqc0ptIANp61AV89ZVVIOck7H6PAYQq5PtglDQ090q
EIrN1aK5KeS5Y8OHl5/fYEifCverVcAJeM5DnIKYR8DW5YQQ6xN24I+CHZxaYwM6
rQoe6/H4bJsOOtvgK1+JYPfoG0ypKqC2KMefH7PvVOrBcmQrcSkVOFrhfV8ejk5+
nSDAIbbDWWUaxyl+QMDiaw229ha2zcCJJe+OXrC81103upfswCFZ8V7m3/bwIVt/
ch8ddYCVxDhiY9JML0Vv2f2uGTuqjYkk4UgAJUOBpObqAa9TK6FPPkPa831jiVGY
iudtduvJ6QnxkuXhIxme/lCBUfSZ11Gg95+JchVaZzoXAVvDrUdBHvWBpS4q4JGh
5CnAoXNGi/r8FjYIwaT0g3M2Pd6966MbxbtxzkSH7MO16oD9nTGr7/PrOtSolh0v
IwLlt9m0letvZa72OzaaAuzGY/cYLexjn6Vp7cqTI1Sz+MN59BRYXA/V+yIROQy3
UYcOMKezLBqGmPBosZmPW3An7yXjjQmHgN6wRxMXM2hAZVifSuWyYGX2jvJnoy6Y
nY13x0Q+A011Oa+wIo3P+HEeeSRelk1XL1EtF4RHRjQCaUOyX6QO25iGVv/q48HM
ocE77wYKGu3mZurrtKT4P+2/Tm6y+QIpgkIBGUOYMV6RU3C2XrOwbVZhq9zXZzDu
x6NqmIEETrqCQ9pT0aanVsTa5o4uhh85uqZlrKE4LU/Z7n4yddRM1JbEl4x3Iosl
CAcGqXrmautVb7IoFfcQOT3/SPXq6UwtzV1DhuiHeUk0eyeLWUkMkKQI2+eOOye9
R6shzucQHLPp+575+OCNKxx0DqN1H92Dpz0YrN9xyeuvKy1EWYvMg+jtUYYyjR2b
abe0Lmv+LhXHaehqykJ/MozHsu64VVE0izfgYB/6KLVCPNambJnHFx+pB9/OzRQm
/49oj8DSdnphVWiAxOp3TwL3oIR63p5d5t+XQH1bmgalJQdKP8+TSQNNA/CCXn01
nt/akgSuCM4M8baACA1YMHK7KtukNkjjDdNBG50VKilcPAjDtSeAKuOeeNPuSjaV
5EKGXDJ6iQIv1jcwqc+40WXc4UqT/gn7jXI6axPnX4EQ2AfEazpzI6ntZKkxYGaZ
V9sf14S+k9lD7irUb1J5vtGz4cJGoY3x6xfxt5ALVLF4jW0wtHYnSLYQ6ZXn4EGM
0D4S+w+ouV+4ztQGdZsJcCAVnajYq1HcxTq3EuQppO1yUDzHKnjUI38sVdDn5/NK
bbbU0KWOntV277qQffEAT+RBtSZO6ggaewKy8kHbyokQZhzrGYrunF6pl/35IxbW
VYM0OA1obZ/aN/jHK4HGMKe8xASj/xJiWy5wWHYpfsJ8Sb8XzuFvbIEycgAAB30p
OUx2q90qPG0lNb1EqprFKXBoee6hCiL8IOSdnQqDmwps9BnOLyUk0/QHavPqJOvQ
oeM4yIab6v0x9kvRXs49Ph58AHJBWTPeR2kcrs9FvI9e2XJQkn13UExjHJX7gpu2
qd0g1pWokT7SEf18zVrEpN+LNjyGCQxpyiVqdpno/PpeHszOScqIagzAhlFI3sLJ
lj0gQZzGqv0G9KcfjHWXMLdH0nBtWbV2V1jkCRLdyaJxPcvbsfSSpDoGmi3Tvg6c
BL1/ktsCjsAssgWufJ7bqOAnV+n9Nl1SHrLvi4n2Z+EKpaD7HaXBR0zjlqUwKp5i
diVEKYKwHiR9EnRNIrQmQr/90cW1zEGCKkMOz7ULr+6sAOHgk7tUQTyKbcNwi1eu
biT0IO/qUH2myvA2kXK7qYlEceWRo50PTfwxcQL5As0KOtjIzkwxpVcBlmzFAX4P
zBmaGrXhuJkr1kFFa1mWojuI88/wgd5GC3YEK8niqW8cGxtryfqsWfO608RTfOxg
bMYdCyGEsUgiSAsImkDGuZ0b8MccWy59sMZJje1MWDEKW33iObzsqzM7YwxGMcq8
cqb/BMQf7/wQrpPArnTgpjYDmCk6z4qdH5THHxzUnRhU8Y5bb5tOaGzSNknRBSgz
4EcyqFTZRBP6GElaiWe9NGIzScuj0QaNNdtO6sXNOpTrgJCdgH66Pgbby9Alg3eY
qGfV69Z4Bln4LM2FxyvrJ4fqGO6XsDAmDqjQ+xCNZ8X8sKiEOryEuul7gkn7/efl
xIGPppLixz797KdTYclmLHjexfPVNN9eHR7sEbqtOuYIFYbof6pn7OdK9FLaZhXV
mMvBuSY8KzkZJZSECXgNE8vh4PNl8fYGp3ScbUVzkOdci51a9/uCLBbhSBG4LZmo
MTFsMfj7PGQPNs5ZegPRTvci0VcmLWFi6O0QTogmxQZ7tJxw5wdbT49OpPrfN2va
tQg7AiHN91uyUPmO6wosVyAjUPd6eynfUAVsNBG0ks+ySWXgC4GzcDAberm13iUa
mErRaWRTIejIFduhpf70tc2FmvWo/B43/WWfs+N4hBoK2elQmMCeJ2LtkqJFyOVB
5IT4rL38L3TgA+NWyXyyRRcJF2IgqrsxEezDkYQgABNjcFz+GvqhWvZfoMiYexRC
OYPtCvXLJGgfcHEAKYujc2CLuyqZw57Gw6bERw6cYRdpH2X2/kyj8uNhQdaGm1Zl
CAG+G3WU0rsQZ8f/VXlRs7kJESDiCmNtgykoFWa95MA0DzmYXOkbtTr5XSqgLjDT
XOYlT7KZl5rtlhIVK891X4I6PJ2u2UIf9HBF8XYRQla9VegLtsOyuWc8jAYoW+cK
jt/zrrBsArB3frP24OjV+8lV6+BZLsjx/jKJ3ccWE3565muBVrxsQjKB+C2AsrYt
zAgeHLbBHH1pbVuAZhAfT4kHc6TM6Y/XkIG3nGxUHUJ3XiQ7t9DM8EUUO/aHio/j
FMkOpONClp2J8zAwaZNMgFel1BBaunaXXhY8VJPd1vh9T27deo8q2ou6cgFTE6Wf
4SJKK9IIPzBp3DA9RSgiy8d3RgaI9LGbH2FGSNyznyEvr0vx3NxvFeoo9LMo57Yy
lvzo+sjopsGsqUtT3kXo+15qytJPMicg9Cp+X6CBtgG4VZQG+14n/xKDS1gINkOI
AasfEZS7YAiNPHJ5JkXD4IolkSr/uDu3h71NOV0Ftg3tloaYOYGO0DkTLRbdHHnV
pcA+awuRsSnShrMSq3yPbjbUS65+Z+rUCDQIr/MmWHzKngTvc2jLO3MKQCatVWur
u3ROVTqbqqndq5B37C6/6mfrN8rOyjUGG8lmjzHtPnNWKVWNbWLS9RdENA9VgJ5i
Gm48LQHLys7GwxgHtejJaMiPimMdojv7v4NkZfiXGiIybmc1rfTv91X0agDU8KHh
4iceXtBDNoZTRXqtCtyOmCk3Q71XweI8P0GShW06UqcsdOTXfOP49A389taexGTr
0ePgsFdmX3Dl+rl+3c95wOa11Gp3YvCGX97oBsIwXepHgJGK49172GejzsWHiX2g
MIZvUrvYJvDHuqFhSu9g/DjkApyxx8nCjQTbHFkJspWMGuKq8/FFndUYZ9SQcImi
jhOITdz1ymjrjZn1NA71t7utbra1/LPpP3RISXKRhKPxZjJZafKszbHiezlTqj+j
YZk8MEOcK44KG6pwdCAaa8j+nXeptRF+VBdWltLfsTGeBa3h8iwx5mAixBmR6H70
W3BT0RUFf4uHcVywkwyrkQZm/F+QnAGSjqJ/NICBa93X0qLT5taEAymin+79sVdn
4cgT3YSCcXXl4GUejJL+Km3y9LsF0DoDaD4jjlmBpnZZEpE8PL5Mfyh9E5huuXiG
bMBAJqpM4dVeTogh1L6TF0ge5Du8J0Y0D9aWYt8nIjnk5ognt1eGFwsPOfT38otg
bgItNmzEu0Obmt58ME4ThEnMydOeu0HGXUkBmD+ucD+slpyeeO7aSNxA2m49P0Qo
prnptc+dInvuliiHg+YheLmYJhrZwCuHncOPHYWZihq7mQG+ikxQ4YDNo6ZXcu8r
LYTwxV8OrCTJA/IfqSzqBy2++00u9o+oy8YM1nQl34ymPjCNbrEpaiHqqvsgX4R4
cobYMjVy0xRg55d4C5+lNKEQ0g/BbqN5YSiq0g3aYWqPuxcuqbqKSGg48xS1jpSV
XFf1MTSMcusH6KuQvC4SlQE34LNTcgwfQlv4rl0F1swnSjOdWBCDVsmq3DGbnXKD
WYcr8SYb59n4/eGzet1Ydvj6LET8njWVSvIoPRk5gxhr4OUy83Y6P3jgmE7oQODL
jYho/1rodl+PVdmX4L3tpVKCV4bMeiDsXr7uBVrTT+lyc6kr/ebLwiOlBFiqYyWs
vQ7PhyIGg728lBXrC+uXy+66oF01gT7aL5niZCLmWPSVVr937eHnRlmfQtFwyt1d
HjMJYZ8k+qVAdfGgBCuk0UAKAZyJCms/5viHUIMXSaAbzO5c7qvzoQOW48+gCRoN
6958QNGlo544XBTSInMEz4FFD2LHU5z1cpXsHsjAMjfxWK+h/CgftO4FgGgpn2rB
RUHzVy0AO9ddPbght7d9zCDaDcM70IknHxq9CIgnEqCb3Fe0svnZpxr8WZR/G/zD
1RjodFaL6zIotWZBWtAdAz2wAeQ4v1ThcotlX6xKBOPjtayjpZJ5yDlw7MfdYDoX
qr8s0bXkN74XgANIEJDusP3zp1MnmHWejyB475zk2tFaONV90VhXXmoi8klPGx/5
uhxVovCY7it06hA/XmxGEn9M15bexrqBW+AjOEW/Qx30DkHa/ZHRutdOzC84xKRF
0/ctYfV5i7mC9e3I/nfAy2EmdKhc1ezQv3TjmEE+XlJozUn3XVXl7qPtqXvAAovH
TIwWGSzYjWCRrLpkTp77AFIOMugbvqvRiIpHKOipL2OgzK5kmi3UOqwn6+I+tkDk
3S/9wFwarqOC2GfTCcWYWGx1zYR1CdB4Pu9oGw5soHuJFkzoVYygQo/qZAOdET76
Tg9s7z1cnDopNtiW8xWTtD9ZGgRZ62N2MrGWk+PQ5ilXSh2OXiyiAtEI9iYZOaZ+
jjWhv9MXqOBjF85c3X005Frg+qDola5r9omHWYFkDzvG/Tnrd4XTJ4zeaJrIoqhv
gulUedgalypq/KPOrFEdpHhJ7wbciEJFvY/b7B4Mdu01h9I5TObV/vH0dgYo5K5q
snysTy/j5DEWHZx9sv7eknIW+pq0HHIvkCZ5MMEr2t/3CAqmLuKduzg/takELHOa
9VVWEcVDsinZYai+vkRFAazKuGCsvwsauUW1hxuBDMacSsQZ8pJakkLc20QAFo01
wlPs0m2/ZgsNwgyfu4ZCteQ5NGNBENcEHfJ9PUimf1x0XbhgRxQRk10IHBv480c4
OD9nMKqbVwYgP4RCdzK6Pn3LSpmU5hv73/B9IwgP/Baa9O4S8oZCSrUCApHR+TUO
owvpKKKx+f0dYT4MKxG4/Nw80ofVSvf37yzEur+r3whiw3OD7I1xFCbD/NzbX4Qa
QGd0UHlE2bmdJhBtlkf6ExbPjJhgC7YLnw5bGCer1729L7MvIabVSzhpzJn4Tuqi
V91juMvJ8qhOh/xw/EXfCVOuVhNYcRTmvWpVH6YMFydjzVvGzNF7jYE07JhcjgaD
jpg3xui8+8Tfen2B+2DpBaLMcQCiTAuq9B/3GY2T0qGXHNFPYsgj+wpwMtBAkg1X
FOiUmSwLbnb/3nhrCIuf1t3L3EK6Qlj/ogBeXVMYdx7PR/DQgE+4T4O2gyfN8vW0
gLB1EB7jLiYV/9vQIp+thN82Skwwpym0IN9WCUO3adODmin5lJV0lXxdcPLuPINp
jVlBjkzjlKUWOaisplWuw9UQu94ObkwAdHwJMDHrMqXHVMz6GMpkgPOUyiHcZzCC
WWUmnryyyfn4Hpl/K58/45KQqbthhNKwuQFtGS2Dsz21esDMQcttz5lY3GcN1YDi
PoUWGe0qc17ThFb4jLebEUSO+AMEtYioVrLiGGhSJ55DTxBgceEg0nk3aeq+GATu
tFGIbKLDsWfxzyww9bDAlSOdww6FIOijrhrlpBPFMiS8/gR7d3VM1xnsfucpkFyr
vYEcSClGLgOGCN6Qk8iSD9yxbTMWHGQ2BSMphn7k0S0qnUGHySHPY/ivG04n2z5G
Q/15qVuIf/Xr/4bAae2Jlu+TqviXRnLT1h+tmjgrDkrKkNj97vkOJ+aUwbTkelX0
sLQPI78kTRRNMcPbKQ51iTkjp82pQv8lAZCKUdvpeWWx/Vg1G5hIvXaSIygce0ud
wf//KV3qthKmzi9mhDQz7HOJZ+Z3QaVd0vDp2NofZQbo2Z2V7wcqpobCQ+L6agoK
21xzYgkIm33jjscF+PWxSK8New9qcsFDmGyGFD7rkN2WUl6jD0ZjrI5RvLyW06wx
axfEOQeVZ0hzsV2equqSFoE9ID2U8J6F4UcxpVbA39TkiTD24P47Q1jqb1+foRz+
2CqeoVm+C4loHrK+9CK/zxi0Sxg+dNQyDNRxkntkii+HR5x4vK2YYRShHXxIe34M
5FnHb5RiDuqrcdZKQ3ar3Xfj4Tuj0WMlfdhJouCLbDWhCH3XjWXKUvs0a1GIfKd2
9w4JakkRpZDpF5QCruyfG6/OB5EORZnkoLuv0Bc61Ormy5v//42sWA6eBN8KvXQI
Hqmer2O2sYi2trwtdwg6B00DAlnmS6HEk/rs+yU08EdZqT7hKWIG7VYCXXSsWOnT
Zc9teJlORPtHPDH9geTSVFfXnvBoER+YmMvTXJ6iqjM39TsAMpMTSugxfR4ojXob
Cuya3Z6GgRYt0q4Q9q9sz+yLf/iGKlKAcgsQ7oPzJ6b8mgUZKHKIrlx11hZr3vrO
TV4bbjRanXD6p1CdMIwDP0iVovR7GMbQR6VGFwKyEhnaXr09L7KEewRYQBK+KQCg
V+Wng2n7x4SZ22htxqNONx2yVmVcFHhcbUlT/U5fMn4F0ztk9rV0bfCs8e8Jjmxu
mOzwF2N7XfgOMjWx3K9wDwgRZXg9NzVe1EnmPccIS+a/omTAx7BgI2f3iP6XvaG2
dwEQV5Ec/X69aNJQTXf47YFW5bUx2eOOWsXza91lJqr0pm0Vpx47GW65opagWy6e
+W/VjLtRFFkSrQrlnU1RVpz8OiuRT+KQBTpVvLhNCEtneRxMQpMk3FTtw/51bAZn
xm/t18gmukDNFGgBHN8oXz76MXshjYZ51QES1Zk+0PhAH9n2MxU9Y75OWBf4UCBr
WVXrLLpJ6dVuZfz/1CYYZEpI0eG8PUq/A62M7DTG07cANmV3C8E8kENZ1nqn6GH7
Nqw2sSU67nUtarrvXFoMKNsHCg+yGTzmCDW2myn+3HSfLwF2xcqnRNGvLITdTlRW
cZBNbLqyE7EaP/DlSqHrhoyzi1RtIldL7bYBxUBg3QHurC7+4KWenNhTyJDf/Fjp
jJAaoJaTFFtgSUjJgAa4C0s2e2fc54K8dM31o1P60FIh+tIx0xbKD/Vqrraqu7c6
GmOXa6V4k/5O6QGvG6MWbJHA276n6Fbi885+7/zMxNeqbQbE4WvqJ2CzvHSm+ueT
qG0iSG1whLypQghaP7YZ+3sKHgcEha+Wag1Dy7FBuMK6Fxk8KeZBDWvmzebXYrh3
fvdAE6ShallcffQoAaQnxx6XILOsXnxtWqn4LWML1mue4fzlR1Ihc9RL2ovCjT9G
qT0uC3SK29fc+elGTKigeXSqK6YZjaYfs7rHbfDF0v6MMuzBfZ0hxoO7LkEjWgDN
0iE6gBxbZ201J0brY5RSe3mRKrbmwYRnjwfbGMoFtIXs+pa4pXa4tQ5Sh+/zLR1X
pfvYr6KonjQ/wktPnZH8i1B4BU2C4ziCX5g34QyMz3zKM0NAJYexxzvTl2T/fu0i
IvE9AN4lFhdwXt6W3uH5npOCAgAYCn0XPjsQtqdxBITHgXSSYC8F3AnYs6U32XuZ
n3qdv9nBnaq0AFsGeLCpqEJT4acBdzd0IpPI/mmnq0GKUBwGUvVxmBrLznQU+pz6
FvtAeXOgJq6wTA5hV4YV3JkAgdr6/Miqw1q5LcrDnq5oshUFbnB1/nKAf1bqaRCd
NxafwcTwG7HoXXiHodcV+MY+UrEzzJcrL2zQ41KAyAdI6Ps7IqPnCzbbrsE4XsLV
0MKlNS63YT6BkMUG7v79qo31x0pmVoLJ7dviyOX/eWnTo2xtHXfhGBmoW/7h4mRM
MaKWmQDQ9cooU8OhmR2A43IqtmirPyZH7V4dULsCwyoJ1O0aTRPojdc/BIqpImsO
tcPqL6pySG6IBZGoKRzfseqCLxrUthR1ZMiTBQNxgqQ9VUrr+nejidvvhjyVst03
mg0uedxGI9X9x5+47EyRHqb0Dfjt+YoOzyJGQ3AADOQfx8EQubU0E8blfwi/GcEQ
BnnWL80QLSptsz800lENceUUwiG27oMApMzSwzEUBiJVHOEAA3u0q3/+MCJkO9S8
AryqErmqZvSOh0SXce7hkw7p8vUhDnvPXGJvYfSoCyI3MUOd3QUubrXCt/TIbEX2
neRILPvf13cPSWA92loKUJNmXypThCcBVIyYx3pFRnBHhubZP3Jc/RHGmeKlUW0R
xn/4jrZ2iycHOB/tSsQkL2bV+bvNjB5rUpD6xf3rgw/X7XC6a05z0JXZPYArj6C7
O7fNiqL/da0/aOIMGjN6VwEmxyby6g0HQLnSQHtHBevSn6MzZisb5bQ9KbAseqW4
RNAq76vW+HIVEk0iWS6NJ4cnCq1YJSVNjRRCqvFp/jYassGzCxxYdXV9O/dRgFtq
kKRt82/2BRFX6BaodbZrhylpAlb97HZwJDTg4Xs8jSSlLYCxfmIGChXe91dPfznt
stsGYCcfWJzbTAjRL6SJFx4kFq/1AxtiU9STtR6WBn3FnX2I2miuf8gTIxIl301n
xR2v6H5moFIGXhbo/apJQ8eYVMKKFgsoU28c1XcwMr7hH1PFpBfJoN4rmeXZrSAK
GOdu3sdmbY/x6wsfxdgrFUbdEC0Zhpi/XYFzWK1MRcO1yIgbAjxYudztEgE/o5fE
NFga4HkVzChK3zAv7wfcv+BfbI58piw2bT7gFxanV8s0Gt/SIQcCVySg13PGQdHm
Af2lbEAD3LalNHPD2sDRG1uZmzAcjnq9zNoEHM9rUYPQJsUfwDUNQVFByIojQjX3
R6eyc3qzAg7sBM+puCLsENlola2AS2KQqtU7xqP7RufMXSLKsIAZN2PrpEhEd3fB
rzZsYRwxX44BQW3LbfzO1mZY2KZj2FWEeRiKT6viqR2/11SGVcJmwYr6ppiNs0Qe
Q2mNVkIpLois2F2El/QkAQwNGIdfjXjFD2vLzGEPgX4yKzoIogCQuQVOnyHJJ0I/
QYtRpc6Q2YG7y2uVkDToodrAUcXlkvMJ6mVMaKVysrmtDHDnI0SeS93OQf4ZZCxZ
K3X1WENi8ijmn5lS8SqwG9CeSrbJzqClZGbR/3P61Pr2vXhcgEM9TlF1FM6vuLTO
o77ziBfyGj6sy9X3xMr00CwFWk/anCpKf8GFmMRQXqSmAi4tSFz1DM7ovxRJBxc0
5zYzB1jOjkG4C5gtHiNUPDPHUa8WswQFxq7MP88worrZNgtOSs3n+8K1xd6ZG0aX
Y1gnsdIzmLRase4F+BPkKhFzw2afFk5mk1v1thMSFnYx37pvvBau4a8I2QRU13Nt
c5SbZrQxMyDDIA5z0yPky9u3sTsAVi4JaIIdZE9SAL9lK+yWGpwyBF5v6BDVcG87
crMgK1OQSikwjR70Y4D9QQ8vjNJaxDFJMMRe5p5Fyt3EZJR+LHHWhDHU6IGuNtlS
o0Dwwdg8HCvi29M6NtV9tlIYimgfgNMfGvpT5w3ZZLgPqjCuB1fCNfIJTcZnpqgI
QnZjvNAi4xb+awXGAiKhVTo6TOhSX5nvfXbtMhNbTjOE/RwImMHUUGYFCupYwj6t
6Gjc7DthgfLCTBcefC/rGlslH2/lnxj2LEN+ixXbAiYLc+nKzSvrFcfBjz9D14O+
nI2JG7B4uQcLrCVcdcNxv/6C9RWnZkOBwpTj/dG98lOrlJ411P3ZtbeWp6PljabA
bQuhLyMW90MNYY12eY1FyRBo8jeMsxRWLbp4ud7CgPT195i1hq/x07b/RDDTwVpi
YigcXaOOFk31LGeffm0Y8NlCK9h6xXwF3FlzjV2/gim3bdI+iHKL5Z0+MQqUYEtf
Nb7L/4uMIsEydBL7532pI/9Fokd/SZ8+9O/BKtAiZp+tnIMBAN+aVerYx5bqjGlQ
yRkQj6faE3iGlXLtjO9zxvNFF9biW2rZNmu20qBe5xyzGsI0xiesWNeLCd1r0hF5
+Sbe5ANVqs/QJoADRplhrxstiWXxQtN4tOv6pAJrBkAaawWuo+qSOpFXb5Fkb1Qi
FFNB4ZefG4P4Z1apwEam17Qp6HUqkhvWisz3468EX2xL1zVkTcGoUQBEqvc7Dxrf
DfF+gxv8rGPv9IIiPYo3PVAfkkVjM7MyQsZvbZfsx/FvC958IJs0E8IAR1Dxgr2J
hhYhYOnf+ipVYE4ktdD3nZX0TsrhFUheCkPKu0n0QmIOfjr/HcXBgkyj6mFJ88QW
U8ZfPzV7x/t9xU7rXAYHJUbiM1gpRRx/ndx3SNP3cDoWSaxmioKOvD9xwWoLlpEf
F8jyIzeotkhMei/R5hZWI5XKfcT9B5fsy/Xch54YGVwyvxzWRmV2Dna6Oc2CJWoR
hX0n8Sj+Y5Xr8IYQUqPP3Ys6Mep3TKzqYM7IlMsTSb1c5BaBVMdq+lORJpk9N2dh
b33Z+n/sUKoyOKOtMCuN8L1le/n1O35JkD5l84rAj6YyA/A4Va6dKQHm8zB1eAvx
9X+sdMyV/vqgOVTHDDMcp8Jo1KzxjIMG8cFri9ylbkE15VjGEqwP04GpbSaTNnCq
efrZm9+lj02Tv8F2CAyTMo1ElEUPy6S57kyNo1JZUaEj+34uyKxXwzGkTJeFw3+r
0Mg1IGtV6kjUXryLuCmCA9xVSI6dBSWCddS6m4gVcoMX4bs1J4JYdpLBpcarUl3u
+9lMkTbkx837PyWegTzCHFyklRvCRFSDuYo79d6GdkNRhgIit6ExMzlt2TkaVh+r
sQZsHGWHtFleVcIf3zaMvPy+K0RVtlZ9cfwfW2Q0t9ip+Iawo3fpwiF3IVPHODLA
oXT8nKNd0ey0Kmis8riw/ly552QotU1GJc6hQWBPlYV0R219Ukeo1ZdXsNqd2Dfe
qxh4Dv4LEeiB4jlH3D0lxSTvSMEPvDFKRQv1GgUrvp8uKgJTgR0RalHmfOxl1iOD
vP7PiixOY0sB+Mid6hswgf9836iO4CpX+cN7Kd0C6TxyByyuJDYqfxMoYxMw67IF
o3FBf5hTUdm2+WECKefVzrC6xjaGNrDXcntSH26GN44LVmfdjoPVuzCvN8gxzebn
UV3FAnH5gauBZvInTpJNeJ4lnUdIwz7FMk3l+vLv2g7nX2WFQC3RvhR7WqHQN3+Z
VbmU8sQJVlodf9wJ97/weUfSOc/yZUr8/6GEig7FJC2+xc1e40ZcYQUhgUBznv0m
uPmgXhNftxk1zdo+G8wo8Y0gDonQ/c+HbSS2H88dEaxdXNUWWJhOZlXU8BmpPgGR
egOYuyEcHNPAg8Gt/WpVV7bqlN7iuJerb/OgikhQGxlC8r/L1nTgmKJ7Gi4267lJ
UJzgY2hbqg7+q1dymLN0QUCS5NK21KmCu2GXr4fgbO+g8zGpFPREcm3guyxcQSos
A57IfDLblYVbiCdl6Q9vLvRRFf/mzAr1f9YdWXCc5+2T1YSN11v6bm9pLZvf3gOK
l2esAMHat5gxLOJ8kx0NEi4ZDC1VrG99XhtA9CX5RF/euo1ggACCUXRNixb1elYS
eKzWRPdbtxtIesaqhBVQ20shm/rZfi59Z9g0Zzr8kh7vJgklRV2T6UwdwT7bCN6p
e3jXVSCLTTI9/d/hDdfKOIqHtXCgXIR16eTuQ5MZHy8zxw2H5QLs21USSXH4PA7b
IwGrhseG+KKeVLW+x+zfiYlVoBoVHXAxjZHo1AYH3qnMLZZ9NN543EzZHVWYqipl
Qu/xCjeKGNjvnmhFR4d8SmAX7WGYO7Xu/nw8m48VEhuQ9rcgSmKwmzwLfMUXWFAj
K8hnmj1L7k4sHov8thWp2JueR4NZpijM0LjAAkVaPUvUBeXZisaUwQZmwsIS7qBR
TxuAy3zrcfw8bQeCe7iSB3nOtML8TX3+V58oVbr0/N8S1GPGCNKhm7YQ1M5c+pvU
Wyw06xHBVxxIwbbAUoVY2c2AboUa+uUKj3tb9yaAsFaCAtWXkUVdUhgS5YOfaDnD
pJhVqAhWTVvpsAzO3oebqIK3dJ7aYFMa7ExPaerLegU5SOsfqG3660Nry8mh4eCk
696O1FARbnFyokQhCVg8PZ8rg/L12MkRrSZrNtr4se8mUw2GPvw0YRM49AJYXod4
5QzVPt9J2fGujXZqwBdMICZdf2FRGpGHPmDbEUO3OMEcazFHcHdDwj0dDG9geSEq
1gfEysVRv8l9DK89MW9HgVRWd+8Uth+/zG/ntpbD1V77LYpvJj4attdXwGMuQ659
7f65hFNuTVpW9kC7HqsnQwecF1T4YLJiqnWbkvhEhPNzktSZbIJ7xfvwxfGB+KML
F26zpS/XFp/n/RVY5Z18xBXm8m+FsSK4KupJ5f7xk5S7x+LYoYA0MguKYXBYQP3n
QKGLGQ0EToDoMXgaUR102JCByOH0oON+waRL+VqzsOm1RwdCKLx11ty11dzWzM7q
951H9ZzS4sWzlyCNp7SWnRt3TTj6vXUhQACYVRa/wN4cR48+HlX++AKgAt5RgVFR
AQZFocqAfcEUopmgVo80QlS5F2G68FG/Kp6PHpyooNt2v9XKFZYczV9I3z3T5BMG
KazV6guJ6xc3qgAHmGQfy8efx5766+fy45mHoDk+m0Xwlngk4mDyF9UUNIoS4a0r
CLThqnUZ3hYa5d7hUIpDP3T/yByq+OHId/y4MvxLHZWEbbZSDh/WbyVKJsPhi1W2
Y0lSWyZXpMgxU+9iPsiHWrlrtp86EKaJRj6UAgKSYeFjvegdu8OkkfmBdwaCyD7E
nwF1XDypUlb35Smkm2+S7YaLxInWVeOGFPi+j39YdK6kWU+EpJwMHbR08d5E/f5u
XcR5tFXGc+8yh6X39KlG7YeS8ED/9UUgA9KWLFvqc5oE8HEiuM9TRDBgkkpHs3rW
UXHsZKnT7epy70DHzrj/wqX1nngdVd1s44UFuT44tRrtdIppu6vSuYMzKT1ovfym
oQtKp6wmUjqF65JmgzuP5Aj0+oweueFKmT3sybTiGGly4pVvQ2OjhSubwXoHVzlE
4yN2mNxOAndxO3omsyePP/Ot8Z90S3gdsEGD10C77sdafrYCyHcKBCj+z+Q9MLCv
tTQRQMzLP+ATGAnBb4ei6j0qTaSlIp8cU1XKbDSH7a42ALPanLuhpkTbHOrHS6p6
mY7nYdzsHt4Tb8gFC9EfyzkMwIkKXDu3YWpGz295M4HmVHajXzA36XqfNCuwGk/2
x9Myea9ViVmsFoTbocvllg7amGkkWdItBx+En+BV+1nLJQlzbJx+gZjpNt8QUKux
zEPFWiJQI8dNWLn6bdkQuR8FH6alldbedchjM/eLlUnch/9ffT057sgNwXKhC+9k
EP3fBif/jugfGoEGEib2KIV0WR3X5+QjUTixVsKjWHV5rBC83dCRucI9ND5EENxM
jMFPFgpDlHQuiGatVLOAoFq/HuoXGd1EXEKGMNdL+Xqtz9CuBr1Swh+CqohYFitE
sj9hkZ1TpkEFhfbSSeMCfuGLj/v4ADrk64X7aLZst9yk0Row9t9vgBi9hh6/silr
p3W4g7QT5P4MfVD+PrARcGL150x8nXn45Y1pfXrhOczNLHtakLAIekZQ7go7ioNt
6QCXB+voA2yhutaqTIPMdaenHLedhLnPGDpRSoCL0lAiimem6iYsFbgu6GEUkwga
vBwb2DCGzN7ZVYxOPcAtNo6BZI3lMxPtnENGkwiv7oWzXT2iYP3gYMFVExhuO9LT
QJpAUFT9QnxlGNWQ19DqGRgi+kjuJLNTgpVvCjd3gyF+B8G8Xyko22/1d+2dhYid
bBnqTQL5dAsEFWt7XsRktvspND0gE+IIv7QOCzCrGdcJapwRj+KMtp2qbsnGtDSe
TbuEQp+NOwZhRGVNVbTji2ifsBq4Bry8C3hfyeonrCKiy3OyBwdN2r47LYhsT0oS
/7hGPpEaZeysZAHzENs+yBWA0EXW57XsFVV/S6820GljLmeO0IC7fSTj5dilOArr
n3/1AYzg7zSdqd0S691Hmwc+G8LEsYq0cOO7mh/jgi6tlPKUYQORK9GBVKWEbBpD
b2A1r+rNwLQsbhuqoEgG2Wd/9xEod+ufW4X8VV6ENFuXmgG5my83NZqSjSxreUbm
r1gmKj1fhmnJm3muPX1Nya99MTElOe7WIoZwM9Z9k/11BfNj/I+lSSVbigpRNIgu
2xwfZVEsbThs2uUT2sIJ19wCsXE1tqmjTT8A1bYiv33QNyUvzTqsEmTELjqGT5zM
fpLZh2S1jQCglAcKTC1OgH5ju19WSJdWyQGcLOhQ9BFUeUM53YiJfkGgTlHccLoO
c7QEUm8h7kX75OKDOFc0tDCljpgE6aa4kfNoSndrd8nSAKhm7efawNUm1rGtf6Zv
R230qA9i9vPEZEfcrO8i/Z6PzbZTdQgfWkA83I0HDSKB4XuAKRod2IJ4UHYqKcFV
P5udCj5iSKRAytI6cgYKI5iCiXE6bnbHENDZ2dxsH34YNzE3PkAmAPo9IDG5Sfxk
Z12YtLJBqi/6e18k8jGvQvEATLz6HDG44CZuMFQfdW4gHF86Shy8oFJJ90wUM048
1Bfb/J4slFktlo+44r0KMUNWSVaBfOgZBgTYF3BkIB3K7MK9nn5WL2B1XkB9rNM3
VQSyIZeYP25xRmT0Pd81S19rpHdQT2bsRrBQY5a8nL/bE4rIWuJhBZgJMIUNeLN5
2v6tgaA0V2fDJ1SnxuHZX+n84qZptifpMPOrkMStn/uh8HG3MSmUzFKntItfJ9J9
fq/W3MkFLGVY4gubMdf9wsRnUe4pAnOPQadLGMWoF8TMJNEvkBQ7y1m4DbWvCGTo
ELBbHa9b/7nqy31CVqbsYGynlf0ANlLTyHixiqHbstyrBlRv3PY1VxMfoaBMEKNX
nuYemqxnIxWVenHRNKnMSSI0l4MYJzbtqQu5UlVpwKCuQmUPGw+YB8xXSe1AERxi
E1uI0cQOJORQ5qTfOcnSaygWsH7qkq2fQ+3Hfh7GBMGE5RmTr1m7bEonNz83kmus
iyUt94G9/GP5cT9e+sdXm0LXzEvcfN9Hb+C0s3ozobT2LtMo8FXsyj8jlKUgrBxK
mKcaeiwI9nBnnAg0UZYz5dDBKLPhqGZiQCE+XxWjcAmQsPN8R8idcDL2y96YQ6Af
LF4p4GZirlH90KljyoKb14B0nL0wDPYDAaxaGYm0fLxF+AyEHhVY7qzxBOo+WJUh
4jfzp2whjTe+sMEVxHCfkLhb7x3/0pcbi5caXOuIdafqMywgsmvHNnxBGsTRGdY+
qExAfKgJOZn2bmLuTfjgb4WVRAGCD6Uy4yQ0OUVSpvo78LR2lqX0COzNDKnNg1kc
sZ/cqAPMKZ4vFkAnGyinLS/8bB3FqTVAtRLPGno+yHcPTIz96jfFWgVBU4MA6iEF
PsxJK42nWP8bNIv0ZoYOS1kY+tWJABGfOnMHHFrHOhgRPQwe6I9bM/1a6MCIXHRd
5KxUCvz0sTi6iNQG/XbghWwUnHWwDx59mA+EHjgnD9cjKXxt2Ux7NkaexBt7NSd7
7/BCEvO+KwgTGV8frqjuC2LJQIg6RrFk2f3sC1kc3gTZZiu4oBVNxabsgd2uaoou
+aYsgt9gvQsmXArGSn2kp5LpnFy48odEXcUOL35mDvPz7VPqRubg2M5ezDu0c4gz
8SrI8q1RiMXO1z8+1qPDf1Vu0rT0ouQJDmR+3fOgw4lBjCAil1UCG00PE12CAuEU
pmC9y0AMvDEQ+cuYVt4PtUzQNPHL16Q+YM9UyHY4hrzuLfMEnNUuegjXtFM5mIWd
OKnIkhQ2FqxX10dwUWLf6ZNGZIzOVbBoxZJc47CJ9CnLm3t8dUe27a5OhqYPLllq
1APICllAmAc7NMSrsVfzaaG1BAs1kt+pUxieviJhB0Vrom/3SGGSI7RnoF0Uy9uO
7hZVQZXZ5IzFIAvBWOsoAOvVCINOMFioGK5jdcAbYgRiQ9+ClRsPfM1T2OCX6u97
BRMdnYBBBtpn0dq33yRc1ZXJRyifp/cRgqtVYfcQSLi2LjzjOr74MOmAkPKQJ2mD
sVAVEi0Et9lE8OWKj1v02qPxxG+ntceAWH5fUQcYcgpYGzgszRg+sFQ0yR77kSdc
D/IyzxQEf7YWG+hQGPqk66XT47ys/AsQC+pv++HCCbUVJTa7BQLCXy6JSfLeakst
gzpgwyAqZViwiDC7xEYzWOF6nNyrBrZNApl0gYjMwCht9mBWkysg420RJmPLEwC0
avCdCq0rGoh1IviJCTs3Qp/UrXs/bdvzVI6ZNZgLRkDJV6GB0eyMuOjus0ezWkR4
mGb6WzSLYgxc9gtHLAJRBiqzj7e20xNaud+MuCGWrjxFBHBa7pIXOvQOBA2Iozk2
rHpDp4p4KKsEd0BYzFt9dmCUTv3ZT2w6PshzVSaM41QvMrp0dIhQxA3dvpvEzjEI
qwhDPh8Xi2WJSrFgZiTYqag6EbXAn/YPHmZL189Cdg3kUNDL5VMbxAHCwiKny5uk
ADos43kbUjlktjBYOsChTtbhVjYePfOdYv1mHWJ7sJmIZTT6sgjlgunj/IbIzLQi
EcgmP9G9GKrN6vzp/fF14dEl/sd12Mj01DVj137ssPHFIj33iRo1CD2ypto3j4cx
ZFhJlosDHcAL3x1vB8L3n2jGV+EksxVNAmtSrRuzAOk8/dmq7FHCar4xHiCnZQES
/u3uLwRUQ7WjOm6FOaOUjOaRRJpOHu7t/06zGI5DdH3Jf6j99whJpZOJAPux8pBe
0GhgjdkmtDnNNv81Mu2Ni6i9gAKk2fQpKhhpXdDeEkvgXQAoFFpNC3IXXp1wm+qV
qE5xeatCwnGhdpS9DME8LC8cNdVITVcoVTSK1QMeX4iQuta7K/f7sfhNiFbnCyJD
Dw0G6ODnygzmudQDIc62NHcEBOetgvTU4U8gv7EhPOQNub/g2ZtMSdVJQL64zdMJ
1kCLzHnry9bNsf8rzufxzBizWotlI+uKRrkASmo3VmwdAL6ufzhBA/8McTq4MZcK
iChjRFTO0eYlWhX+e9cQXRvRqPYQOYa8YAMViUayH7TlYb2bkBOUPIcMwyeqV3i2
2vHX6MJHYIsjtn6Bl9dQUSzclmA5p/h/smR87bzuacsYh0stV2uTV71WeDx0w+j5
Ei2GFocjQsGbF14oaYGC6IIh7YsiZwgaHoNqoQkk7yfNOZCSdWGS+oR1aF7SbHdD
DeFZ3dy2TFsaf0xwT4RhLYMA/1mtoG/ERBTSaRI4kf2gBy92gQVpvWO1SRSeqijU
ATOKQzmDWCrom3Qg79tXPy70ugzzRFcrOz1m7//pOcKthjErtbD19aN9Scad7FLu
LWIoKmf9z8B7NcCHBlOFU1IKb0YAgq9fbQuhtx4tnQanFn1lXcS+JPJppKJrufXC
gqsouhV+qxcuLzaOP9e/hEedN00TFR2VD92UVlfauHdgX/uLwlwaH3QmaJDd6hJq
3STbrlXPz06tYRn8SddC1F79L+UCw0yxEFgDJyn6raur2GsOLxZ0BZTheXL2A4ub
aUU+rZU2PwgO+2Z5kvrVNM+yP6c6GdF6Zgz3eEz10C4GqiapshiQoPAB7QCL0tgw
SGtrouj9t9edp8W/XrUVRvWZe84vjmosNPGbz1WZ2fRMOIltNZixxS/AVphzBpRQ
kSl3Xgo4svFm7EC81iZcwG2bjckBfZ+H8FftThXVxjzWviv/A3itoqlSsTcF6UcG
eYS7r+FrRMEN0zrXLAyJLJpjS1sMzFGUEdRrxacrykTelhCfroYNq6V8Yqa9kIC9
QdRP9y/6CQWCPHzTiRdoWy9EDxbCT5ZC8tHUP5nty3iv5ZenXqPYl5bkWm3mo8FO
U1Y/M1idFHoA/fZJtLY4g277Qr7N1x9z0TwTOMwQLuqj8SOhD4Yoh+623pnoO3a3
40e/eTwZ+/vTSF0ZqhBKFSvl0Vrkr4MK2rOlRVZjihWHBCCh7V3Bafp1LNFuW0jo
jVh1FRolKhCJkeicDZGKoTNgV0775B3JqsGET2pNgxKnTMrDKNKZHWdu1aLbEHld
BzI5I0gX3LUAVnxBj8wvppUfCTxW/6y/eAyzlwsOf/OaX7KK1QLiCa2jIkaXHmH3
KH+M7ynj4lmPnexA/XiL+Xb0s7yvl8OWC6e56JJz9IrGCeR2yrK84FmPTgFcHE0k
/rqz/5RlB3IRi/Xee/HB2HNB1t5uxRausfNK2w/E5m5xS/uwFOPTWAunhlD+0d3W
WgbnueYc2SB01PErQW1QxCwsWV0578sYnIP099Ciu6oZVWMZ3iZaVYvldc6IF50L
sNB5fA6YAOK+1f09DdwCoSMg8hdB50J6euSrtTuj+GmHcXhhYvW+WTVCOLPyiVst
7/JBHK2sSaAQ2v8lLO61ZracElRDZVHa+tBaQiNQ6Mb/DgnfZkJMIF1nOfbgizZZ
YSJcbn3x66+NqnBl+nfhS7VprKPL6RJ0YS+OYwfKLQr0l3vvhpiR3gzLKgalUVde
WwLBZFZEz5MzIB9Nc5uMKCptI0KTecORKVlBcy2Md3F630UtRLqOxOUt5CAxiZo7
4Gi3PUKETjCYAmkQ7dHXPVvSmTcuFVQcqmZzgqkOuaFHsaYxo8YyVOKdmGSGUMNi
6fdAdZMB1h+jJh8jkkeddP68JNDhczga6ZA9NbqN9B+Dn/myg5sKRrIJ1aYyukGn
WbkqeA82f1C2fuwOhDFMFZX1/QF5OkGdx8o7KyHONlxREIvrGFRXjFbQbHCmRQoE
TL+Ev1JLthLiDhLG4rjW+r/xN6nVNtaPyLzipttsIAF2rssDnC4zxM9hwNF8F3vR
byPaJf8TbsDq8oQ9IyYJdEYJW/ZuC0BKFsZN/V+4QoT15IEfRpkgTlU5MtJdod1A
19XW81mYDFbaLh9JoOsNFDGv/lzt1rINKZwQru1UlFe+tY4OqcSTQXzQIu8DvBj9
+/TTe7Lhj4coAk9jin+GWhBZiNYRATa54G+5aSHmpUAwGt3G+a+lBzG9hL+mpH9D
U1NSiM3FCrHacrJVbbucCeoP2eZKzlMzdmbdKTAyWphFBGFn1CxXr99Afagmaqqk
p1FwVvqfWGMJM0yJEy9LGg8geJPYEVdYkNBi995zryDZXBb6j/8JxqpupHT1k4Pf
1asSANotUTJjyW6lyfLsl1OCriRLFT4geAHv8tHL2H6admjrHvoBf6gTlv9e1jtG
VWiB/8L5ZJ6kz13Ck0Cjr3+4oDlE6OYwZittyShI12HTAJHMsQ1ab0OIYlY0+4Md
pmt7sRU7j/crMkZ4q9ccWFfDVVQH2GC2htjR4AoseJY+JXeuwX6jivdDdGe/g0/Q
dZ2L+2NffkkLOCMyX2eW0dsu2oKZy5fF+9Hfa9sXGk7vSgjHoca8aPc53aktMft3
qhrT2/ch609TsqiORMhL9BvFxTKq41yN75tOUCI2pFQ6CDtvO4/pyEqlBf4H/Eft
yPoVaPCJaENYWtVCIqdJUJ8oMQCYD2g+Ch7or6a3e9VuP2ZI6acLYYVzntXZ0uns
JLNJFT7i7OsIeGuYc27e023xQocfZr5CKoYTEVPQngR4apGZuGhmM/nTSAIdZjkM
GqhamOGCuiBqYOkl68uyQTBvYlCjrkBpw2OtX+mybHbQFeK+5K1bXMZ0lWTYeiPv
nzNvbl1zVEg2ihQ1I+Jm1KTfkkjpA554uERVgxALLk4GCenH/sKtCzv6YJHHqvSJ
SdSP743nM6/jrFI7UE1bX0fU9W9z9tVmQJEkxY1PG62gszq0DT11LJDp+Jeas0wd
cfGdPYJB2eJePUIP98pgKOFOkbgONJKCTX1J2jMMRDRYdpSUdOrHhfS4klFXi0UF
WlwOhqezWkpqt6wqx5ZyaF0Kux5eswnM2Wp5vLd+kKuGT5ZRn8VB9Pxh43rQGBcK
jOAbV0l/wWGMooM8gbuYHJTObDco0gmU5ea4LEEv+E0Vu3xXbV1dZcYedw+XkYSD
8WXtjBaGJhriZZI4NMbwy5Y13XW1POvbz1QX5IN6whMM1kq91FX7h1NpTk/lQgb7
WKsoOobK73DW+8/AAZQE8hZynqtbdShnwbaYW1j8ZHtJioln2TnFLYsEGs5nBnPE
o2tCWEtXZTFgFJHMw6VaACOkzg5Q0Cfd+NFC5XsiAQPs0+N2rq4LCKK9Lq1jeD8O
DhZoyyPwRqJ8DhYExTSAGh346X8MJAdARALZqZpzxR0ElBUhAu1rcOv9hIfeOlCM
mzvbpPJucjBs90qLb9jE0ye+cM2btjhdSsVUSSppodsvAQjFE0EKrj7uZ2camrom
MGWsMICilpN/FnVL51iBDTMkHqTw4FFfu1/LJqRfFGfjR9uGSjyo/faaiK+xmrzq
I1+CjOmqeY1NZSpChltj1QJZPRyy6Ndyjc9FcKSDHnrD/hDA/W6z8zcc5z/o6v65
Aj5228aHh9YulkWEYHMIpImrLFZj/8vlFpOMNN3V+dtkYGLdc00K4IVxBXApQcb7
xm8RHKuuViD/7gSV+5/uYYrQweXh8xCaKiwXXTE9+zDg4iInzkYCu8aukTiC9GTJ
zpwOTXasnD/M0ZeC9P24Zcl438FsI52sL6UA3J5EBdbcC+5hANna3ij6QBbcLZ4D
4BsF3z4Cmd+6UA0nCd+y2iogG+r4vps3CWmMzX1Snml4gS19gcw8N9/e4oGD6oyc
RElNtroDdkUO0JgcjC1RLaZPp43UfRF0RVjbvrYeOzm6krVfWg7ZDAZpIVAZdt5c
cj4Tkm9ppXnZ+Y2IF6gP85AGJggm/CVsl0Cz/kUoVxLH4Izzg3twMoq07e/E1T/f
8GvBb7NIInBXh+tEOjBgf0FyJe5UN4oQ0kpAkimFPF6xRP92kIqLGnWri78pSyFM
WMAiR07rrzFVkJLumviwo5q3QS32qupvNOuItAXnV3ySlqN/zZHukgmVQc6Xvieu
UhuiPZDsnwgVVbU62ppGj/NvePWKLI5wu3RJ7L5Q4qr4e5c9LMu1HwD/szliXXne
PUc2iK+HbMR13d6J16BJsdelA4y3qjdFtaoZxMD+4S89SaUtpCpvcuTTF1AODlwq
gYdmxXSdlnMDDmAAZl1bm03yIgitzx9wWUaki0I6a5NVrnWdxGqVlHHwaSc7UyGP
YPFYXMjzLob368gt9UUnMXS2lhnBjo5s3tItHqK/rfuZhCz5tSIXSQGYmZ/V00pZ
pNMskzas8EHgY1KH+z41pAcumBj8kW/XHjD97BbCJOqQ6mdXeyPtHLIwW1joH+0V
Bz1kcz/N/EXjVJ0imJ9fDFZ4g9gMGGQo75oyVaFCI3LzSOUoOTSZBkz4PpJbCjZb
niEWR6/Kwf1smuV0Seoy0GHH1VEx3POB5Uq5pOcU2g5AUoIaFBoEm6GQDSyvDevL
cAz565CuZmcYsFz/xgOpx9GBhKSXhOKZcwkHqN2fJR92uE7rUyIo1EGBw452cZa6
evvU2R/YRjkkzQb7YevO25URPsOg71ubVsPTzEg0UQm5hEB4uZte/oNPiDy/Hd7z
DbbZTo1Exjxfqman2frfMoj8Ff++lBluSO+EaMK9gea1AI+Ug20fPFSo0qAeGs9X
KtSS4SXYwop8Tj5ZBgUnjJQH3YGJ0S8m6H7+dCArll/SgGDcaQlEN7O4xm9B8WcC
RQYM1ZYnv05xJ6HJMA0AAgpzXLsow3UTGNn3MMJiGRAF9eaMpaq5L5EmEMdXpRRS
ShdXvnIe4Dgj9Jo/yS1PblOdABziEijboKWBBpGpjzJdGgbrdk7DpqTvVZVVbWdq
toSLIMVympfpp7hVvstPBIQWwR/UA/ystSbx15TdyIjA0T6edIopHbd6IIkSNOiS
g4YTMiOtzvnMgaV/FAsSHxlH1TijVM0F57EZki88LiQ6u2FHyAsyC1tIHI5LlvQ1
pt8zo/U0dJtErhyOU/1JWFwtthtz0iCrqVHO35Olcor/GPgzeYN+TgXbu7pYINYU
dN8h2WhhnadFOmvS9HQ6KtIz38hV5No/tyfRvOfOAJ8hyGlB/0p/gylVP5Dy8GeK
zpsq7cMo1UtnbIaTeVGTlShJixljPj0Wpi7YnPrhnxi2FEn2zClcgvh5v89Oiy4/
SeaYzcE8aKgdenyI6swbqPthum4f+Phtag5MM1O8eR7HnzBG+i6m3VtZqXPs0DK/
WGaJl5aTXWPZqxksVHFZjnq71T/YQpsSJTvt9QlQ/7Dt+wEmEmtudMY+vNktuxIh
dLD6+rygvYL8o6a6Oj2UeBvL9DmpLR5AoHEirxRj5HjD2J5rzA/pa7IiMsidopQu
f1cZp0PY3dV953SdurINjIkRJrfvtHrKBqxqfO2ksnb7ouBVzPa7IpbcwjzmDNuw
DqWa08IhldMUgYanl5wxbZfu23i2IVJb5GKQeo41tgwPhhDk5ubMLO5m/R0l/8yC
ZJ/aQ2CE+FxUv6TRAkzP/XdKCbYwDdWZuESQaPVkzo64unKEEjJiZXjPsDb4Rh9w
MofSNt+Ym2MGumoHayk183pVj8a1VOlGwcAXF0wN/nfcuHHq6Ue6SUcKIg2xdU8P
Dw7EuyX/y6cR7hgv1zrfvkv/2DaUOaa3YvGAluB3QnyRbVgRmrV+sSCyKTXpH5QH
1WhZXOcwyP7RPhoGJbnNuyzDOV5m/h1X3SX2OebyJmWRvwRrneCdHRrWWWBXpgRl
06ZqGEGUXS4QLG1CshMt8b3r7P2FN+kD8oVxh4yUcVsg18XbVjdI942pgD/N9V3F
TgMI6KEaRCH1ArcAw6IETpnIuTHfzcJoyRuzvujDmbnu8gD7Y1ZApvy2UNmZqA82
Kh2eDpfUWZzQjyjYGPfI5Utdpn5/ReGBSG2/G64EEihZKOmg8mf6rIf1kcjt5YL0
b9XXIBi3wmXBqTgS8BApfBOAR6eJMNV421Ft+n0Mn1OBiAG4uZ8ea8iEtpOOApJo
jCqsJ/8WEgIv5+0u+j6g5ffHE7TCmKCfWaFmvsbFfTNFxYBvsy1Q9vterMeo9q3U
qg9xnTNr4DE6kfSb1a6A4ZmZEGkxR2CaMo3sJ+qSN5e5Zxx/5yVf2CsNfU0qk1ke
axGngnt1+yK/zeYnDAtEG6hO+uBj/NmkmhmbAy6Up/9JkNuCSjfecN4cyRrG8uH/
izzVpbVzbDnQaXcjAjceAgW49LfpoijOIs54JC7zJUjOMDrwA/Ss1iwByjnbUrSJ
JhSgYs7BfE9hiYyb+Tzt1iL1/nd+hg5mvx2Q19KD1IOIBUe9tY2/31E/tUiyz9O2
IUAKdAtCI5ApniHiBSJtupsUh/xIg0JScHiiatI3Gov6Vybfa/hXLfqbkFSe7B0/
iGE45tR4x2z4HpOGWFqEl4kEht7eAEfAfGwDZBFpUbE+BZsJgSnU905geTz2bfXH
aAb5JS+675UuTBDsAGhCzZAAeAItregfgKvMtrzNJ6IlVl6tObTZ30ph7IknjvK2
y4Ef7qXDEGJleC8oC0wJ7ve8HVX6BelC6IFXDQlXEQgjV6kefGhWqFvztpsTKAwW
7CD7C6MVgG6GJxbp1il8r8k+Ze4lKNuKRwynuZTpXdoCraiXnMkqoMdWAcQdQUUO
/ocE0bnZSviDBTRCeoKD9F7vJ8h4N6QJcTkFDTpgedKE1HwZqgzx6BYWZ++RLMbB
MxxIOA/dOvn9rkCPYUJARXjRxccalp8nXfAtSZD2v8PMnTas1Gz21eAAw35ujyZ7
wPo6yIXU9KhRqIz+C2ed3b93CgHHL8HWrv/OK01QfAql/TZUSlIG/jC/9bBjHITq
y14pMeYVUk4/nKVlPHRLCHxvLfmxY6StxbN2doXOaKtnpHE4h8zt7m3oC4MMOh0J
XmjXgQfrs+pkDHSdgMb8h5uA48pQmZe/L2ji/Ln12MB1VNT+k3eHnBHBzCqWwlLR
B1nmNRt8Jb1SzaC8IR6Jl8BQpgjI4VctN1TSeDPTn4Zcvi23k43qWSPMaHsLE74R
8mCqYBNXmXWkAMg/aNhgXK71j1WEBRLo5FV33b6Ao/twNOVOd3fLRNWa5qonAN7I
qf5eHOb6GDWcla0gonU34Zi1SUZemP1sFihCfqnf3oBXo0NZLiQcFXGUyyTP75Wn
mC4WjyjhpXmn0QAQkSr9CX16PiYAq2q1PzOnYl79BQeangtM2NFnk+vZCw6/4Kug
SY0b5lveqgc4KJY9CnLkFmDgAOX2J41wYxEGftoD9ChVhiKxzw6UZXw5lYwo2mIV
0qtZlEKmSRLFyEfI+4owSXWZj3WBJ0crJv0g4J1p7wkkwBSebxVywuCsj+J+evud
HIqO8xUKFecZae/feXPVh2pf4xH18TFiluptD7maX8LLEXd6jzJgdIN7HYYT1+3F
hZLuH/44106kT9P5laQCSpOF2XlAgpf6i3AEt7ZTVdamGhXpSOrb/mD/Psemtpd0
rGUWYm/Mn4PL1VRwlGbwfKECSZLhkuHxT0rjL922j1m0Kbj1FX6Xm4VcMex5tP+1
scJo9xxIur54C5AuX1QujjEXZYPx8syHF5JfExo47o/qbcfeG5kRCAvt6xutoLcH
M/FLah4BOHzISkxb9jfN8uiN/HRFrWj+PgQ31stUBcic9IO9i7dgbE92UZG83l1D
Xrf1B6KCMn7caXhIiOZo6VqMalE8RycKTeY4/kzser8EiEMdxYf5YJjf/agdOksa
WJgl3he6xS64sif5vOj25wd4Ml8QYN8vhAyw9FbMJCuAzvP1gAfldEu9rNFZxuoo
JrmarbqfRPH8LN6CAnWmARDsz1OQWb2Cy8nULPZDpgHOyv2JgeALgZduHb11kwf+
oKXaBllFG/v9Cm5709awBk1VdolVNrRfQEZxOn9LkOC2CBGufJqCxGWpgjViWnCy
BRAtFPNaAKseQwX7lDsDX0RnFypG3b6K0rBsFtKZcHmVFBsvqVi3jH7/epmkhtZh
W4tTXSRQ3vZ1vWJQITKZFGJ5WC05+eYSlLoZs3lfWDP60mAoQhOQtA2KdAfGLG0k
xlG9FXJRym0I5+Rx4Oil9sNNVt+8FDe6BkqT5+8WHn3szMKj2QE6jG2To2OsgC8l
LSb+lwsLG55E28fe1Zux4uH45MRxune5FSNARcVOOlEk+/mfSwfUM5zdo7eIBErV
HxQKusBqz2JD49UdwH245yxJ5oRlQghAqsVScSSaRugDD+5NenU/A2DG8YkJZ8wy
cBXj2DOm8ZFd/PTdZL/valeJznAVLlC8m37+hKxXzUTa2BOY/HADorjNYr9tZD8l
SKHSLuCSEInttnz0aL1AYWMvJoWgaLJuPpLve9RfVK2M2HQl7LzzJqz1I7JrQsBs
sQbZ6jray9rDGyPgBWNkbMywwmFfk9cMsJsAH1aRKOu9UcIcxqBB8kX8gY8JJuaS
1n/YFso5RI75xpNj6mVxbhVsmiF0HAfPmPYdzE4O82H6sD3vM1EvFHDLtbLAgDRs
K5qPJTFkoInxCXee+y3aIX/GR2Nyy1W/K47TxIs5BK7VvkArsIVboRjX65fCmIH/
Qo3h/BFE4HqxRaKqj0I095FE8VR7weAtvnHD3ftju6j3W7UvuBGf130hJ5vvhpxp
xyrDEVovEDn340SGOJGS57Lm97tgKCVq+yMuXCQkDtpx9GYY0yYz3TM89od069CY
eGccE5HiYBFneZKg8I+z0rGKEM1X9XThjupoD2pHQx6cj/S2QbAeEccnUni9Y6Y1
lY6ritQyq9ekjSpskBoYmCySMJt6tJDSa2n9D7zRJCfrCCsIqKwI6TB/efJQPRAu
hD+ec75ib+FgLesgvXbtZCqllxbeDzi0mDtXFOnGbW9Cv9DBGZDxvcB6eC3YXRuf
2P1yIiebOUTfdgf7GtaKjG6w/eA5mMiY1WTeQ37VSnk3k8IjnOlb7pHmSA77Rjwz
VZjwNLPNAA/0rkXd2T96vZLcmxpVUoPU8AIkqzirNjI2zk9muno2Kl2f1c+DcaUF
LhU9zvvTijkFcA++2ncq460OO3j0tuGrdeNAm6e3wzbnJEI/G+t2mrenxyqPVa8f
AvMQ4gFqSe9QTXfscHwGS5D/bvLQivQHpsOAf6duHvdkoGXOZ/tyftfEEm3w9jNw
oO/cmE/bWS/YylRWYnMqrd/vhVR+PB6OCQNjrl5+I5EfhkMcq7Nh9eT50i4ShNZH
sVP1kZunnkONjcJtGhHQcdkfKZ7pXN6mn8zzI6fW+nIBNCTlyBJFx3aJ9TzPvtsn
2aLwnQj/MjXO1Yvqpeu1uv1MgQr6BZ7nvIc+Yuvi8kDjr9XokDLr0bUdXG4mHv42
YYkr9h+zfjMBL64r/HfNpXIOFa8tZHyu2+5DLPT9Bs1sf20CeaDur34457+I+KTY
SffrC4wj+WRdmiTKXSa8EG1RAVRQ/MAxlqiodknOoX7t0pDBQ8KdyrgjuR4ES6QP
HqQxaz0sXmGr5N/VK+KqBf1odzqSyw2uTlEa7joFBkx84jsEPI3rSvo5yaOZKVd5
2UjnhOtdNVpm1DXSydjxS+OE2EGe74RD7LZzabAMrBophAMIJADmxlf0INoHTMxE
MEsXakLiGk8rvTpKspTlZf8nw8akFxvicKiLsed/LDe9gqBK4wB6EjSxi/lTZLt8
32n2LVhYugwSKIhlaYnpgn28Y9OtkLpVb3pt94RYZXbZdcspYhfgiur4cLr0CMkS
4a/WeF7AKH9+q+AcLPHcoxckLY8MJvFZ1Eh5slaCfBscXb33IgKGUCx23l42r+gs
I3Q7jYDxd44DBhBNglj+HMb2qgTyHAyIRs3HOt0AHaHaNo3/OpvtcUc3TirBgdeA
oefHsDW9Ou/YvulxTFVIp1R2PhrwYqg0yvb+nT/0B75cNSjZbARTQX1mjav/W3eI
CUtXZj54Dazz+6iVyy1mCWOKV1Cfyx38MIBv9RDIlfCxSmaBthAkwxWEDwTFAO9c
6u9w8y6e9/T2B0NfUzH27veRa58sUdS1fdTWtRMGej+cR537PXY8m+hrSBxbLZqc
4l2ApUxY3nzn9QlEMR4Ucw4uY8DteL1CG7jt15HH7wrHjxh92nLQKzXjOx/D+sv5
kFKPznP6sEEFPHnCHGhdTzYxRGKTQAyNdncAvIoTh1DgiLheRVPUKQA6IUmikgeb
apWqIuO9iH/l8DS2UjHSQeFGrudPZm+wUUNpEJecwOoCOU13Vl4VlRjzWHLMqSCM
nYShosmddULThgpFKy4DAMhMYiC/Ql9RKgga6+GmN+8QXoN7fOHJu/GK6R57pUx2
uGtFMp3k+I6PjValfrEXCaT8zBqMg9Jmw0Fr3K0k2QSZ8NxIOO/pB4V8a8IogI45
cfRKnCQhML1GP4QFJwqzxCpYr5LlJFWgfoTEQx/tqiXe0ESkUTUZ1VVaJdJx9YoL
2ewAmTk68O696aiucOn9T/xjRhZhltvbqw5c6DK1zouzuhdt3Jg8AGTVHhGI4CVy
SzMzo9DMuhSxXBcLfV5HacM6kpI1VgUsSr4fVGHpntZY3QXvUEURoNAFmEEe+zJ4
GFVvOvO7if5H6TyS1FpwN4QUWTRbrBKiHiz6/8x8oi7xAdYfRKAnlGFYOFh98igu
3D0OAADBb3YfaRJSXLBerXa6cu7zMJId2zWpqtO2rfviG9LBngaOI4mZDfil34le
mHilOqKgAdoConh+PdKqXzzhvy8DNHzLFCXprX6TS5TaB+SItB5Uz3C5uFua28ZK
z9GkypUKMDPH2u2jv198O47KOekPpcl4tPaO4isxySEPcute18TwmXDO7AVAhZFI
K9b8aMEsWuVk5CueJHcqtz265icIBNJSlatQzsoI1zzSfRnGNCrd+8QOWOzCeds7
NvzmguOMEeZ6b30mfk9hj7Qm+g4XRu3LjQEdiQ/1zbedfkLLJZNXNO5FITx+ZGsG
YLIi1NBIcDuzpcyojoXWSGyNX4wFzsCCDjp9eVhDSgqdp9qFVCVQnB/mujSl6mi2
upbH4upGybl7pazggbb6WLvGBBKhe8dyfGTO7Ck2gIOxtZhmRGH10bYP9/5CdCLC
xdiwYl5xroDFwzYzoJaR7q8qjTygzZFBdRGfzUP3dCJQkB5E/dsAGKLVlqgzXthB
7aPRWtD49VeJv2zB1PNXrJ0tjU1yCs06v7UpeO68c8A7NkOH628RPe7ZNvALRDoE
bLMy5ZPyz4QYwlItHYJP+xtTGscKKvrk+wMDlJiCO+W2hPbzdXU8w9R6ewDrVmGU
FAfpIKvF61ESRC2ETDd9TokpLl/FJ6YG0/gEXo+w/450K0V0PVl7EM6nc5/aDHu6
ToNbsqVyxAjyqEafrajAuB4uACkt6WENI062mhoGu0/loJ4zMwu4js8bJyqjS0dp
ZO/jc+XoIisBfksSL6i15KwjOUqzpv8ljxyzQPqO+AsJ6e3MMOTrty5FBQVusB3v
FFVPUr+OoVORiHD3aVrYn8k3mHJ2pN+PEymNkD8SUwpt2D93tNCgT9OMkQUrPn07
s2yql5llAUZeIr6s0RtkeP6Xs3baGP5MRju6qpeVQanmsdg0h+prKLb/LCpyX1BR
wKHzZvVMjOuo5pu3IDtuCiJDiRIvfhBXblKnM8Km5JzpztQqWLTrclG/UQKTItEU
Ch29QzzgyApY73tHcq7yHqaNz0I5ZiyJ1AKhuCpV9nxwVUS14pSSPJtCd1Bz6W4A
lVqa+d5VrbWhu+yBVOKZ29+J9kmHy1VGQfbfG4Om0fwljGX7om6lOLheJi/Frro8
txznrYPUWVa7cRd+rxJaehkTVfsC5U0c7WEjqMqurVetym1OLUIZiVHmKDTrLKO+
NtzNvS0iJkYzVv4L9C1Jwmwisos6qXOz+HKS5Jg0PM+f+PFQLu/xCTROxfb+vi7H
Bd4fXg1GaJHI3o9zyiqopuKU3r8BZbtNasp1dccU/ZrK55NKpvp31C/8ERUwQ718
JHd//rOiiQgA6C9R2//LDbIdJo17cNFy9w7MMUFVrlVqF+2yVa219pHvOwKdndAt
NATP3qKRjrfAij0xxjcPBgeFI7DGrxNUuCYNEZY8CzesZFOlzY/6jXEHg1za86MS
pok5ANiTN37o/gRFZZqnF2Fz084bsUz135QUbwtjTRIuBH4BEpdVA/xndTDEAoeu
v1klJCJp52D26beb6M/E3YwfBz4qzU1el25EgslIY0Di8BH9daI1G5Iu+bmm2E13
UCE64i9CSsQaKiBjyj69q/KPGY9VquBglF83ejYNpV7Mnh1hRM9R2otwj3yOBczw
Df2nT/FDFP4HgLt2t7qvbrs20II4ggL6lQlHVi+LYNzTXMHjsBXALxmXzV4bPeQI
53Ih0owDNw8heR4XpBLDKl1RM8KenK+9n1LVtzlmP6MwAdO1WEEZc0v5nI8PIcco
dyUatVsp/FYOyLqrv/KHuvnZ/96+f+ujNJp8H0vjzM6nUs2ii8u/Vgd68tsFDrsL
S1yQXaQ8CCGF5K34DEjZGfvP7BYe3KpAHCI+4RaiECQJ8WqNyWKD8w0UCkcmPeZr
vncBCjQHQsZckq6ZcTRiSYOxbOX7UfF/eLtG6GULxc6zxwJj/RWyoLDEdYCmVp7d
3cq15AWsTnU5E5yFgdMS6dXQp1d0MrgPox8JZTANXnh9bQHPO5jwfxDBHF0oIj3O
nNhCEV3HoLby/YYdyrls8m4vQhAldGTFXJW8B4yScbKlPsLci+0AkuXQ9J+SXrra
ustvc+FNgsKNS1CGYjPrhI6Xo1dWnvkO/QDikbO8OUNuLq2ISlSKDVicZ/4m7ssO
wJefjuN/v5FkZawwKJFRSAOL2gjywicaJjsa33LlKfzrzJu12FmCdytkYH1luHVj
/23i/S7186K8RonAgS/AP8KXAioWJxUbvKoeXoz5UQB8VMiRkcI1CL8N5nsinsLH
apsr/o5AmkACYit1J6sl3tja36hz1dbTp1kUs6K46kI6mvCWrhbk1fx1moHvId7j
iwchf/AHY1uhvyZ1ZPTbWXJWyJDAqIsSBBTlHSvlYbJ/yfv0YskVD3hXSArDO3lD
FlaEGsyEJGI+IWA1G2rTPR4M60FNJJRwMg+nqTL+pnHPNybwIiaefy0+Q91VFT9Z
2/Uymh1uveTwC5GLUqGQ/gVJz0fKuyi/U66XgTvfYak8ciYRRISEgL35Ffw15+Cj
p8d7U20zNCGgYpNJKiHjW1YTXOMDh8/z2eGRJF61RKqFL3xcoQ4ScfZK6QkxRmNj
xiBN5MM/lt0aDH3T/lQThdtZC7/5pr3GyHiojrgOyzKBvGyvPNX91Nmo+++VvvGW
Xhi10A20Hm2DNDn8QliTiEHxnYMOju+KwAtabV7D27cNfvESHZ9PAe5n2qP4fOfo
ypNxYbQc2uYJUWQg5w52zQ==
`pragma protect end_protected
