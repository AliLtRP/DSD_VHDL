// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:33:34 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
jaxRqTUvzTUgLfbpPplzGJ/MYmmG8IWXu6rJXzqsGRCggs5AYROPHNdld6dH0oxc
yULG4M0qRXqH8uSLclmX6IXcuf7E3ZbgFidw34J402q6As+mRNCQ10wd4s/CzwDK
J4y93NihRE2obPU0wg2P2X8Wy1GIDzLs0nVITPMljfE=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 22384)
0YitSUNBX+E/wkcJHnv2beLSCBvv/56x8YDH8bxjitf5eTEigD6PIjbJs7OGTK/O
ozkvthu/vzEyHw2Zkr7X3lde5rJkmZEM1yABNTywGPVkNMS50mvcRmADiZ3ASsEb
5OjPSX/9TNrE3oATETmzWS9uZkm3ZIzxz6IFtaWEH0uoQnLlqVv8PwsecqEjub/8
+s9BfwIxKscvEyL8wWHBvD6tq+R0w9AHN6MxlO0n0m1ZUj45SvNlBvmmd75NZCK4
9R9Qnqzm6f7BQWoxAA9/A448SOxKQIuQch8Qk1Jwo9y8d2S/nNpO5lms914yN/4f
14udkLmGtlmM1UufV+7g95IXNQ0qRk0Gan1w67YxDTRYl3nbrzjISA2b8LWCL8Fu
i42V5shukbr+TmyTg9aTye2EKutel77lOthsnDDU1RLkVHvci1a0rPYT9xgQxeuJ
GThhElN2Iamxa3p0+B8AGut2TZVdWWQXZuf84iKFO1cxWjfHb8cbm8nYt7qWEZVr
aJBX8lqCnFtUvvZvSMPJiJpklt/f6vIaX0aHOs8wht/Eoowuc99jeW2oAKS3L4k7
Ine0kMziMOGEGUqFZHee8xwHfIpP4KCQgvghhD3kg/Vvm9fVc7zJtRU9u7I1/zv8
kCyVB4aDlgUZL+c8YX08VDDYwLxXBxIE+floQ+SfMKYECgKtPn+7aZPwFeazBz9O
wfRtpfvUP2FHdKssxcsG58yYUi+B3IajznYolKZHgMhVemMtVXTNM+YyLdnNRsJB
Wh2DruZsK5OPMG/LmRxgQgaKkVs3TiPEYyuia7c/Jm80lpootAGttZHY1Sr+anrX
esGqYVc96FGfFQPcAoF5flEkiKaeky7CPCe/NYOR+XErZiqh4IOKxjEYTtaw5UFy
4vp14OFv2GHr4o+vwjLHGFqPxMzHYUK/UKsBbrDgxjSnr7zMz8YajIeETIeWFIUx
9qaRU/5IfhPPyym2layLo5GQJm97eUYb5GdT98KoJsjPHQchUasT20KLvWdXOyXy
RYqhzqtEH1rzCHB4DZGXhgD2R8Zv9FtI77GknTrxuGJMrlIkpiPa9BtsCgxM8XPi
G9q772MESXxingxa3qSoby6ZK47Hape13EDQR/572GpHP9JhkSpWdRnoLwqdpuWN
AypLcrY8/L4SGstsH+cCZyStAcEuMPCI0oowXPE1GBqvRayuw5InpUUKgwvClPvN
e67mg7+Isa5jRgyfwQFakpthQRyFU+M24OOpOx8g+va8ot1NG8aGA6bDrhiJWsDh
IPgwea1x9j8+53XL/D278/F4a13C/O+/+987CQPxunekdim+Q/uJW8eMCMKNHcI2
qIqW9vOBjXOBCtsg+H0Bse5xGYUtahxJLFyO/mTZZU5/KsLx+qkuxcdR03d6Vu21
2Dx/jmX4QpM9i8Mm0tTRqrbJHhjRN6pyncDcO5ojo8Jg2Uay1+yoI4l2xehPFYHj
6I2bl83QqBAc/9Z8kUhhbq2M/vY+vOHKt7vX4KY7BZhS5MOuzdG1NTnVG8RGmHma
oecAohWUBmyoeaXeWKU/n/4GaukgEViinUewVXQCAxeRKkN+jcAlfge+e5+AnUC4
3hNQCaGxj1Ddb2P3OllP9G7p2Lv/UxjjtZE4hLBR/RoZD0dpwAnQchyfiBhkSGBf
9lLHTBk3XEc59AnTPKSt46LBxBjvAiZ7bsncCpCGGxztD6bIDq2Hws/FSt4bgZQI
T+RGvrp9cjHUhrq8jsxAz+fB+dNfW4fcWHikegWEo4ObqHa/oy5iVIPa7+7+WeCu
WKFZvmXc2UThr+I8+S7FBf0uHJCI5Qcn8E8c0zVS2BziYNcSAwrILyIIBs9Bsr4r
WGqMqQpuVK7YK5EA4UcIHylzBdCMhCluS1y8l6cWyhOYYRPvTI1Ry8rPQJmJpK1q
7w3JYY956MgDsSNY98JJEpBuAl2R5UXb/SmH2BVynq30vIXUt37uexDfSSaCSVUl
40ZR47OFONjeve+B6XXc+pjndjQ/4QKmcF1Cmtg/7cvWNnrcwXpLVgFjfAbibh2Q
t2p7XrHO50cQcOwrHXVgMNlTo8s4bl5dU6O8vbO7RIuaaIaMTCv1c6t/Dwb3xuOv
F/acnSVThPqbhOxH+k9SMQbXv0+GdECu/E5YdqtlXiyby+F6AKJVeeBTsX/a28h3
If8xpPecu1g0mbjs4fFoqgyVJZvJmX5+O3bCFkmAlJcv+gQEe/E38Uzh+Utf1/aR
qspDv/x5ApAgKpacDjwUkdpKGxdT7z9j0DRzxkzr5nV1D/ykWOAONLqAE//Io2F5
wio+aIGmCMe9Vk9u9jZExNiO35RzxJrKabv6kA47YHTNVwHPKcjFb0jA1ECHlmc7
rLVSdW17zCY7RG9dqJ9HFLUoLQwuV/HHp6qXGy1/lxEbAEly2Y+1tj7r/um7mBwB
u8lvU2Mo0ungyVYDurllFifTCEsMMOeKXuRkVLyHOOLgBFnL5jNrbKaUdVTp7G4Y
zoepW2RLslF0DssBK0YBzOqkAu79qTE7AhV53wV17cI9VXMUihlCNpb1QJyTVlKQ
zYkOY9v1koQNeAjrdkFg095If7vodm1/eD4rQQEIERdeD/ozxdEhd5cdS3dMlKTQ
TY517A7QUT6ZX4+ZgI6VzFWy/OLWktOHl2a6hL04qEit+d/e6flMPDa2BWnn7t/D
+Cc6GCA4AnJbMe8Kgf14NhIBrpXna1l4Wvq8Dzv2Ko9TfuF+TXyBortmZ8OpQYTP
78VBDz+TLUx/APl57ZrPgEHZhGUcP1KykBtWVhWekEI4Iv2NWnLm/o/2HVS8IWFN
9Rb3+kxGqS01IsIEa6wV/mHX2zdn5iNO0P7Jw4FHNf+diTuptH1uNQ+9EggpxtZO
3Yq3Pl19mgZ+YYDXPU7ENCpALAHJwMnYGwFpUANh9MqMC5HzUXySUvVe9skd8cUj
J1sx42A9R/1kbnGRT9DKKOL1iRW6fvnBZkwVNHpeDp5J70D8GiVwbBXTFOO9GbxS
yLLHEU4gl0+e4SC9N1aUEpMHvxOVljG/STHqeDjtDdHwheJVWzM+OjMg0oW/i7Kp
GkCKBXZznmnlMkXyTCfl12JWG32/FBoDk07q1KAOdYX9yeGA0P5ykXCH6gj8wvrP
oH/sWuqZGIWXtjcbt+51t1W/ODrYSh/yTpYBRZlkJcctlTNsZ7FfBo2IApke5Cb6
zBlrr6YLmcKuIvo6DIdIgBeHdf2p3yx/ejOfcMhT8oW1dxtyNsmncfS+StZVJz2N
D2/EmbLx+7rlXdPZxL5xGTDwiYvkxRtKYHuV4JpkoNsUjEhGrkan7Mv4kRN7wCYB
4bqbQjKZu210k5lv8gBsaakik0Md6hZcS9NzXiwMlqATyeIcmH5a6Rbl8ZAWnQT+
JA4NCcdNbh7Y/Ad9fCA5XNPZ0lIOfu3757qRjTIRHiIft0yuVLPHx9x3FFFeUv3u
XTAJJuSQix2dPxaEFJzkX/m7VBHw6vdCCWIK6hyZcYC+6VFg6dn0w0ECh1C74Q9V
cSFsKfp8NfCyHTR/e26BgADU9s69iHKQft+8h/WpIPSUDpJbmu0J1/C9uUUjgTLV
0B0UeFgbPh7aOp/6CLwzni5ktXGTXlYANcEclEY3w+ap6dqAKFmhPXiCpHArbYdb
lVCyuXaCYbXYnXOrJovdoeSuxFU88NavLRDkCq5geEA+hX3VOI6k3dMwy76WuidL
4ejMOLyuXVnUcyCr8alkoNt990dGCE8id1xyg97E6uecEG1imKM71st7XA7SXkI8
pAHAwfEzEN3Hfw2y0ho/U5Xsmm72YDEQOoyupdxsytx5E/QCQ9k+sfigwBRQ/A3i
iu9gHXNwahE5KOj2M/G3odIv1v19DD6dmzoNE35G3dna46OOm97eXsUxB+hVyiDs
zMVJYEDeslK4QytMskKk71+Hy4iA+F2gny54BKPX1uQ/jND0jFvQ6YgLpqu7kE/z
qDHtwR0RPB4wnaaAPpi7B2Hdq1xKcspHh7Q7HyLCrGqtx60eQgoPeM4X34tFHKM6
oIycwMatyeqNyVCZCECzwRnyZ7XcV0VDLWk1+/PQB+UgDU6w4Nh594z6gwPtACPa
FJN5pMTrXkuMahylZm+GSABwuYSH8SUDajLGg4HZc5Ps5NQYrsrdetWJ8Jp8Mrph
TyFIPQef9846aPIOj2THqRYoSJakLdvFeWhnygmmnSK2pW3Pc91ULSvPMRQq7OGx
MJb6OOZtWH4uUp6sMinRqPe0Ib6sj7QtzTmd47RPzrogWlgH4YZbkjAvEb96kYHB
rvtrqrWlYSoSdRRTrfvi1x9+MAP/7ejCHdSz44PEgH12moOnWMaF9CvGM3CyTRto
fA/0thvlamTcoVRr1iliBTTixkc+PFoT+CEpNodzrZASufF2HWvh3zAMSb+YxUCP
RngBS12GFOh2k5seDV//gJVidJTqCUJNs+w87iqSvojETyValSuj/B7KYl9bAv6u
uY872SNrce4gEkfImrKBeeMFEoPhssy/sDjrURovUPsXHlHGa/4YQFjoFCHYNkBQ
DOv2NHDmRT6J4kc4Pef2PIevv9NfD4lYromXPbMcHxP+hXyLtj1xjK56hom4ZMhW
pNFaR5IbETl1dvEzV7B0tNpxkCpqP4YN8864LaackC6KBM3LU5VgKzhXOi+gGLat
QPxjibvNCjKPWWmOZvAXxzU2CSARVuUjqutySmnZEjra/ZfCRVKrg1/ppO145JSc
NGswl3B8Q3piXYcW7xKIDj/1gXpQS7HDDKpKMgTwZqHZ7uq7WN/xHvWHYwp5kAul
nINiC/zxU4kwJe0ofjrpKlKbRzgDwA953LIccmNupY72D1XkdkRcnOndmQ/rRDWC
RFp+hPW9uPHQRIwfVMnZ6odk/IXRwzs3Hr40J4TJkdi9APCV8La8B9oq7EXjjEHw
ZrNkCWJP5hUXAtPBmgYzM+lqsLl4/+e6VbmXHIrE42C7bZVnsNnGjRAjsfW9ADDe
OqKqy86sp7ur32mISov7FeBmvt7ISLYgaDQhup7Li1RiRp7cHPD5VV2ydy3UNU7U
5tYLS4b1KmMoPvyvHrhOCmzG11hRbt+fKYBvqqn6KYXXR63rTCQkBaAdGw3iHfBa
jAYCX03hKUUXQ1s3Z4+gzW9BPsWTMpKNeIxK0/RdtfQMkutXDBWz0GjNKMufVUJz
peki3KD19RBmcTu1JNoJcIv0uvSQtU7M0Ny3I3N/zRgpwlEPW3cp3BVMOex0uKk3
Lrfiz7qiKTji8D07f7bluiHM2DjtQMC929oJHDoTy05tN3tGuvHgPKvEKvPVeF3m
Nm0siBbUMvYHvhdq9gpFbsCepFmCbVa7wtcUWXDeE2FRp3rav9XliIkgmRqCzdf2
eAG14tzKga5jj0p57nUYNmjX2V9FbLmJNgYzUbX0Pr8e8NMVIR6rckf7C4yOy8dT
UGSZSkBRxQu7Jc2KbHwCcMACSfmzxlfR0kiKEmM5rcJzPVpy4okbMRcIvrKtSYMQ
5rPV+43xuvBUMVRudnmqSIm/T4dOk068BejSmWKZlxcAQHUGArm02BosNLRBlF1V
+MpTLyE/lh7uEJmNhR1Q2cOpYVPzwhCvsCiImojyWnGtdrq6E6GV3HRrnL9FSpEL
SikZKnc71rfiIHNuMiWWeq2IEijjbNOg+oTj1jEa5PVurKYoNkdrL/LZYrmZF2mj
ArxM6Bu2pu6NCD9VMfJ7biOd5Bh6kma48BO/BSB/0iQszNfaV8O5a89vOnqSMf/7
7N4Z4INQAaaszbnMe5zbyJE+CUVtu0XhX3oRhSExR6p2eNothUiVM90a5NJKZz5z
jQs6QnIPcsFQ/Cmky1dEAvUsGGKC3v2b3gAa9tY2hB2ERiQ9lKqQP6oo7nfrC7iS
5lEZNuVYD/Gh80RB1O7dPEcnMKecWDVvjhhiThXIlWrdFqXSjTdGP3FIltMBScO1
N/jCpV7fLd7ZdN6CrmMDb60L3JS4oK7aguFdmjfr9fEodGcUVEEKQzIp9hELH7DP
Y+AwiX7y6gkT2QcS9HC9CKIB+TRfs0KawFOuQew06VCRvOojQ3yCbgzvxkm0ik+t
HzBxJuXchtHCJ5kOdnWgVp1aakKAfHW2S/dY9TMY+uKdA2ybh6/IIJKe3wTIKx1R
leu0f1eHGKsyx4pPxKOPufP6W62wfcADyayjDk03SkFSzNw15AwFtOI91LMB3UNP
HuvME6rvFb0AzJ+jXCnF953QBX8VS05T5O1SlNbNJZZA40iesA1Y0YxzovAQxjzv
jw9iu4/hLR3vLERQlsOy2NLlr4z/nL3MoKTVcT7iCDtmUmJqXseLHjKAI32ZQUDv
z6pKaEO3GHbT0laNPzaQAhMCLZZ9pk/GMuK8916rd7K+qD/ZlAmPnenSdXrQWs81
i/fh/fIKLhBJJyg0qZHN/othTezIWmOORxEE8SmzoMLX1FYS+OrXGdoj20yZWfQX
NKCxTzYv/BEtIqc1tzlct/Sxfaw6cX5Jo7pFTH/AbAhM/wmn0sfJ/sjC1fqawCYq
8s+ItHs4cUxiUb7dLpSNDIiMnvBe7vbwRuZYkSirKuzdPSyyJyhT9nAuGzuukzE0
M8Nx5KIjFkQmaq0AOOFc1BdIs6HKDbqtGcwK05SZKN4y+9PrdWutuy7XWnt/MeQx
dpwWXv1BXeNN5gV2dLcEAqkbDhcNyalTN1n4PUbbcTHmEZDkFoxrmT6N4/yHiS2A
aPHPwGGxDuHVELbl42ullwA3ZY5Emz9TTKncmyjjFCvhujrhdCSTwbNIAB89j7qI
xu9xwxTxz4GFFF+zRKWRu/9izCCVtLIJfLfW8xLM1y9nLmZu+5eUYGo3pgd8Qs4z
SVlTtn45vDQ+VW+dkP9AIakoqLjBH82Lk+A6YvpIIQcYRz0vRmdbPYQqVtNWJQGl
kdOKACZvUzbCY6+SSa10KhniVmAWCXT1PLumHrQ4bceqjxMLM5GCHnnEzIGmpHtT
fsW93xotWimofbRWNMkSlbGjcr8+pjLzrpgWOvQDokysc1hH3Xv3naogg4fRnoIf
tOnEL3ZMDfXfC9Ox4aNomNfqG0oaGlNXN9exeQfquED6jzz0PXEWwUido4bEuwVA
+tSBBaBMmkyfmoRDt2U07p2LqQHTNaM63Y8Uz474G95I6pfYO7i6yLF2yLYa73xy
Bb/uy1mFyrhJuoC91ME7oblCNnXfYIdCuSmovsB3Z83Al+R/xgqyQBsLJNdKgfMi
NhBXjOSEjYJKLD60fW/Uanp7HH8B0abrBSHtLIgXVAf5Drxacmjsf3+Ab6Inuoay
R9tifp9C0QcDhzlkBWMvsqP1zXgCC4ygYbRh2WORoSl2AroFPz6r96qpjeW0bz3x
sAYqtRaaTQM/cq/+qxk2XtNkXEfQBIpRZDHea8bAvhOU5+mfpdUNGNRdgGcfdc4v
p4cQy6kzh7OCu6cFfxCABkR+ICzr4a1kWqr0G0ZTEM8nPjZtbHKTNtn24vSVihoi
FpIJYp2vZKFhGl6mIFMTvrTzWlo6m8YDx+t+QwyELaY5/N6c46hmK/mDhG0AYJ6w
zFfIM1jsLNPr0yIkqSBUX1VI3vDqEu3cCynRGokBmMixXmsf7r6X/8xSLDnZ+V/g
2ksEZ/UilDCSPfNvCn93CwmLL7T30d4Q1xRMMzgd7u7Q8YGT6nss3M9UJs3ad0l8
yqUohIX9r6jKw7bqgn7zLwtbhMyM76LvqIHb9P44pysEKH/Nbq6wL7/HnKdmLaZV
F2BRcmIgNfGHYN/ghzotYcZAlFDgTJwqAGkYKN5QOlzJR9Sh7/kQAEAl5rJlf0Nt
BX/U4+8WasNWSmEYe2KRSTc0tZU1FEmIdGbIU7Mf0dzqTvXlmEz+13r0s69qhhaR
M4fRS86+h2r5U8if0fmcro/crNqWS5PxjjpztQ2ZZ3iz8Wa0ExHGMvy/4f+9fZ6O
Wz7PunwkosaBOX5EuNa8AnStnzn6eOm5fQXqr2vadrVBZZKVBMbNh9r61D9RLaQg
vCztcdN46pyjfRQhQyjtGSLskvn9Fl5qhdTUmOmugBhj9O2je/W2+5mN5Fk209Jh
zQojzBtzOnBIw4wKAPeYvue0LeTnJrpPXPAuoeuOXy2gseZcUxl97WckcJgkFE+5
4AmaJLzrs9cFkUmCLOonXoc1yGLivpeUnTr+3Np45NxEf/hZb+cX5JAoQkMh5Tgn
MKFB5c2+ayrdbAFoAgywodeYRuyOcMVQuTIsjc+1wI42JveQ/RdpUyctXOqBgVCV
xJSQv5ouCGrH7Fv0ohS6kQ2d6M6YftTinJcZLqTe9eMTFmHrCstU2+Sz6yzfux/w
5VX7NRWeainfv5BdXeKJD+0/OPscO4WjHik8OfGma1onuCEUVw+MNRVP4viOxNJC
Iykj5BTPmT1xtBkXkIg5lHjufsdJN3OmxKINqrfnAatMLpQVWeXS/jgrP0ZdGYDA
eWugO3sHHZ/SL45VQvRxDLnfKPl/k7c7ZPRfiKWd9QLbaEGSawKsHMJsv8ngSQRO
cPqRmgkR7TY37gq+ujPZHHtXyZEQ/wVl/f7K/5E7W0h+cUGIfK2EJNcrtgPt7zQA
VLs+YSEX40dYIKTw0hhx5D/MM2z/WkkS8a3xtr2eQO2DZVHyf+xUYg151dZqRle5
xzZdx8gRoSsnlv6Y1Y4YBMkQSp396uRJam6HA+DNyF/tmQzdS912aW40Ni52LLqo
LOd/WR/SJ0VJ0v5Czmtac7LR1iCQPidMJwuPAZHYua8bG5HSiKSSYM7YzrRylXT6
2g8+AJeQvxtySwLkWM+YNndIS2TRScnh2sQXGgSxwyEskFY4qsrhE/XwZo9tPC9a
C9/ZNlKIJxgLFDvyjOrznJRY6k3HBD/wEi5UElzLRA2kC97ObNXA2qN7L/pHcXNV
at4Gcz3rkNR9LNbVVKAO9MM9R9LC1Cgfyksg6FJDlcArnHWm877RzIHgeoBQFPvV
2MA5NWDOeOTJNZnx2oR1Jnd+QuBG9SQMOswhb7TkR+ciyy8ctNaJlBs4eiUWTT2S
pRZx8Sivj4ppTMk3/aULV0pm/hdBlH3WX1fm8lZ//zNONM1xUI+gzlPJjDXQnMiK
B1bGVZOwpHck+Giqfrz/yO46KgsFg1Ez4uKsa/AX3SsnMGIvzZiQk2Yke9S5Fs0I
QZDBjMUzgLimxX4AEBvJwNRtufEfGEZ/QunqtD/MQP6g36wrm9yQvCif8cDJa3kL
BbaQvi+ivEoVliF9buadi89MUwmRBolupKDudwSkMujKKQ+lURB1/n0EiWUgKTWV
sxTEC3ds44h9ef3QAaKcg8W3qkQ5rYY+1Tc9ZurUY3uQKqndKceioN9LIMTFh9iL
5U7bQp9gm/wVLMwrK/g9OhVSrZCXZQa4fxnlDsRi92Oqo6Zvxz8Uu9lhffUTQPwf
mmjGbqaDtPtz7S+VSPjU80soEjmqEZ2PZa7mVpzrYdZ+rrDxy98eusbB/dkAA/Me
DHPDPOM1eoF46mGQCL+kDG08AVH37wda0KJXooJHjz9dSjEvgUdrilYErN58dLvW
Zadz5FrkpPPhxnLZJYHMpfZWzcWiEBFjEHdACX/V0CSqjsno3JPozjCalOj43RIG
2eaNu+fKu6H9c99rV357cZN/T2Vb5K8T/hX2rj1yPU9gCzcJKNu27FLnpan6yVjS
2biSqoWagAYTBw5PC3sROw9vm6VZ3eXVljnlI0KC58fg3acSUwisaAamMEhFpwDX
BS/xH1+nN99DEuKL+hDQAE5urqBtE2y5pNQo1L+1f0HlUS69clyyp83GQ53+Kk3R
rH04NjmS8DDM6vTssLMnzhAwvMrQomGshBvQgIj5sOFMlCpYfLpG3i6QkzVNP0qE
mAF0TYaonpPyeOE/FVky8MkPe5VSmmeiVMU+AxXz0c6uW8vYJwqHgjqh5trbehpC
61YooT9m2GvBiLjK3thJDXdG4YhZZGjYqBtU8XI4OR7sWMwPkJ2sQj4VJCC7BEoI
iyTJ0EPTT/Q2cayGrK9mDztRTS30kuCBe61zNiknyI/HKjztiyEZ3h+Pk0BkSBpy
G29DdsVHveva9AWY1Caj5I4ghBecwDunpeg/E8ApXApdm0C5rc9jqenTDnUHE9rm
m7uZjKzGzq91MG7Hwpztv2kFY1jInebxGdMZ3Gk4TJQ9NecRtEyKHhnRqAAmcm2p
gSCiWdmzfPdEVQEg6jTcGpdl7n7O8HNoJMwNrfo0+FwjmAK5jn5VcEivyLJki10/
OZxaSRnh2rDSEK6il3qO7tk3oUtlWbAHhMkeu1yf+Xpcggi6HdPzCWUwGOOGkish
iv/C5gnkYzjKXvA8gJEpl5dMyzeTTmArqKevm/5hv0An03lI/F/nTojIcnQqUIb5
Fqs1S2Ca7m5FN6Xg2Klk6zHmxseEuE6lCUQ6JG5xPjmaSbRXQPICPZa7azV2vBQS
moLwBQVEbcbqlum4PszqeZVQGqdRMC7ZAIQy083tasnsP8s0Jf7cGPen9iM9seI8
fjaH2SK2t/5rw+zdP5Caw8eRALzXieoq2BaFDSnYvtzxKXNnd7I4FtS2PKwyfxEK
b20atERfT/Ea56uSJaPpE+ejWO6XwOQR6okRDcM2pktu2whWkzbo72hysKOXSvQq
qQLS9BBwehlVv5AkBJiQIit0gfIvWlBTk2jtRYB4niysuFQgFKSlE5odYE5a3VFO
vUQ2ugphV1edPDQiUA5xKDJRxMbRvgNU1D1vBQ7uCaPWEqRAlzZPr1Wd6H0mVST4
XEZS7Ck4aV349cZhWdSU8AtrBPEM+If70vH8dEoqqoATANk5WmMs1JRm/VNLFnww
jzLbP1jwoE/m6QUqxx91EByI/rsmy8nLizOoWH8aOnQGqNnr6A7muXbLnk0ZCAzK
AT5U1sBC4NKbrxjAKwqvxsc4pni3DIdwJGWxZ65p1iQbklBYEc5OAhp3zucfof8X
ucJtIkzUJDzHvNeKr1uIGJPvjhgC4ljvKnvWvQQVtZF2RiVi/0JM+Y7SQfv3dUAD
RCWMbt/kEGlh4a54Xspj5eFSJz0YldMDOUbsJK/GW6C5Sj8T9lkGvX7nLczwFwlR
fHwCvFh89tzTBfE8Kawff+Zi1Bw++zLFtG3bQYQzYAl/HMLirGzsrsvL1nPFWdla
opwNHCbIH22OqYlzIncCoS/p1rqp/zsSSLHwuIHsTZtVSO2TYoWWIpZktG+sXwKY
hUW9J2CQLkgmrlwzUEIxFGqw9wEMZnVdy+548e9tM7ykSOzwoG6Fne04WpiBCPib
SEW1GacYit/O58QcjfYYtQIlcx+bA97fURGrYhL/wBQszO9PXVj7mFXXQ81ccdP/
pKlB2s4KjGR/biwEpSOKPrMHjRfyJK8zn7l7z23ILuQhjW6pzKpsgT19t2T9aAZ/
1W6MkoQh3+aaqBH/9MFU6WduPuwLk3JoZq+vjm68rXabyPGjJ8dm+Ur0B7T2uuv2
KMUwM3QNcO5WPV9r1iN76m45FUF1nz08P1Y+LyJu/b4vBVLTzxKOp9GlXK3QLIu8
rKdDrzfGc2qiKymE0DyRm6MVdMfRYsw4QjF//DUMRUE9MzVI4X6oU2feR9eZu8Tf
qQKaaNLKh/DGufbv19P+yXoU1elG5T/N2RVU1ZcP+Q1PRHjbiiOXiOhQZL+fBHIY
scweXyua1GNLlRZML9x6TPA/P1lUAK0lYDCUV9UbqOHUDPCEBBypLz729fXveY+w
znBXKXMaY/J1WsoYjq4fXoad70CCZaM2o78/+NXDooU6t4EMI24Or2II+HcT/6Ky
0bC5+uzmW3qgFpy5mdus0HPwl1b3MEvd3UYy1jvc0M0cIt/7VqbCmddE/u1vjsY+
gb74uwW3gEuRGl+iXrrocpsvmzFePq41VX12syDAX7/HzanzofcM4HpgZIoC0VaK
kDJJYUQf5hA+ALnt/n60U4KXceH/UjIVjEZvS6mcEvI6AG4D7ixh92AgqL6mqAA6
8FMXpvxE6bwfa4ZHuMlCY5adSTfN5wTi53Ccn+P4GGz3KudgcDsq63vHGuCfAC4y
URx3wH1GoirDuyrOG0Vx2r/B7VvqbR6MDHF6gAPyyX/f1u2uohsxsERmfecm+1nO
jkHYDe7S4MmCabLJKCDl4yr5OUgFzkNaPS13mHppBLbnEKKAbxvgsMJL5NouEU6Q
MmalERZ6om16WaIH1kDCIkUYDTVdeeA8T62R1NM+Hcf+yAsYjSV6DxcbWO36JjWd
aKJHDseCy7k+aOCVJ7dhXJIhtg0+7t9TiKZ2eiqEpEDtU4RKQLPAzfxu5qyTSurt
tN6W7AgHINCmkijMqhEsw2GUL0kmBuJtn2KP0QSyQkOUMR6CEmxNyxwYVZHOMa2m
v4y71sKSVo5pDp3KDp9ENc423RG1YTpHyXeb3Dq0VvOfIFBFLjMfebqjum0da7c9
7Kgrpy5z5pX3ZVu+U1p53Je2CDdzVHAI9lidf4UY/dculEIJl5iegO76Jb7v7v1L
dRz+JSb7InQav2k1WI5ghs3OBv7Q11nIteUSGWDSkybnY2cfmy43YnimeyEiKuBG
LHvaai33Bflk1fcRVXUaaTL1/uInyFApHwX8xi1L20/BwzYncX9uPuJu0KaTp2/M
U8l5/1E2/AWbsMRK0GtRhcolWZP6a283J9mCXiu9IjujugN83K1out8t6GFJBde1
gP8HP2PhsKwhObZg0+oADGlFjmxxrAZc8QPGvNtwfM7jr9SOfFjOaM4ntGSU448m
yhZ7J6KYYJKOVDpQbWBttcxP561x0f6xOOvdJtvFs2t6XUrrJNHg5B/qJ9FYl9Jk
99d4pWFI9rfTNWfOaUaOrni+UwknJ5tVMlepAUJCDvZYK1SpOf2MdgXEMkuUcFXW
Nzvu0KSMF1JRgEeStSsT6t31cTZXlYzRA780G/4elywS1ow26JYW9z8PWsep5gaJ
svZezsC8Kw1bDUM+7vmv7mNhKeTZaPePxwOwbb48tZmauNap3z/QSP11YELbKpe4
QNyayyi6NfkFdB9o4sY/ZjmG/TGTtZXmRmsaPFiqtBz9C1waZmix4jeQaVuReMtz
PsTjbba1NKJ3ALN5EgConXA633wUJ644ygBDXlxAlzPRPQwGbczx3RwEoTgolu2j
TbNWuSMYR897XmD4TuLov8fIID25P5tHtMk/94Q0RDK1L6Prekmq2RDljOQSyz0a
GVMu7FQ98nuxpFyuKpDqsvvZq0tgwfTDq6EieRC9AkGgrxSElWXGWb0dvbI4ygbS
kdeqRYsHBcJUnY6tupWyKXVx5yHafhEbQFw1hP7uMUK4i9/q+Sqi/kq90/oXesNZ
XweZoWbTahverQ1wrwkbp8EBebKhrttI87KsZnP7KP6nsR5BoGM5auGVPqiduLvh
y08GHVP3/1NsvJgedBCmzRK4mhL/JvqBKG7IvnoZG0268JSu4K4QAqDM/n82kNiK
PZ5+6sWl/7/pIAgIMGHKlwNwvB+RosZ1Ug3FEWKo8lLxAFuJj8K0xNiZwyVR2fqC
xsVeiBxps1mKd0arNqjPmrm7g3g1X3QuvzR7lOzIcpVXoyRMpgBMG2YPgtNgMP64
+EsTwHCnI9Y8wE28KdYsXk4bqbtEk0enVULlNRE5AgCFeNn2hZfTyMxqRR/LLQUX
NvATE8cRi3wYo0rn8YtYjjovlNyl29lt2OQ3Q7hKRGCo6hyLJRaFcq0wz5L08Udp
ZUb0/SE3VyJylfIkuEIG3C21BOZKqNNivwNdH763iipXy5q47D/BNqhcjH8Li0X7
xBgN3jK2yRqQSjW/hki0xXwueQSTjONiqTZWx3oDcnoVEIcEciSxImmzekGb/hfn
j79CNSOduwFR5OmlSabu9gfps4V+6dB7I5ByICCu7UaSui0aKEu6FQLRXyEj8deK
BiEzmlaDgzYsXeNvB3gMkf0qMJLCFT37NZ2PF4331sMU0jhzl8564ToEGLJw4HZJ
mOPXhOlqwJ+JvdCB/TIYkm5snxXwHfr7I/9lHtvxekv9JkxeMi9FTIbZ4CBD5+tE
0HeQWhkepF3orHsUYm6NPIRQfGzEzmdKH1I/XYQzdaXeouBZ6bdicPwL2ztxselW
9HVMq35KSIKFTCFxHBoisO8pJRmSiQv+jySpa41vao9t8atTnwVWzdncWZZZ+GOe
GbzTXmG177rH80+5UWIDfA9U7QKsTdXXIjRzXyjtZ4+l/01cjzvBM5qu99t1+w9I
ES57Mpe+4OmzjijUrcE1jkYpXoaVotsh1X9SmoVzanqvVhd5Oekl3/KhCyoRQqLt
QiNKx12fHU2ZytYJkhwcB3HFmEAbVtrXE2/3j5jPeRzkzQ6d4ucZsnDv3I1cH84M
onQ3hlNdDcvuGHr+HaAp8v0NAGIAvc1SiNlgyF3UjavS4q4+3N3j2GKVFJrBD7es
idBS1ewkUN2UJwj7J0qQHdbZLqdezA8k8HBkwSoYXV/TBRUFk0CUIUA/aZa1mrQU
pk4nJw5dP23064eToaxLQX5uzcz8rxdLs61YHSFyI4AniFrhyanS2vOXRgxlpP6r
bSRJ6K+6VNOS8uagv8WvLZC1DnC+uIKDdu5hQ9E1X5R3TUrbWQ4AhgfD7ylBsUdR
swvae8THm6xEX84jA1LOktM7IZdVURlf9XEbBTBCk090LtF8MQ4ZVppk7nkC8l8Q
Di9+UspGANSZBNAo1I2I22rlj0bs6dm3iwO3FMuU7UhHEKLPGEETJFg7Y5VkKSj1
vqfuG/A3VyEtAoF+ZX3tP/Na2klIOg+CKNsh1Y9h4BdVJTifX1YprCWIte4lhguT
Un8epW+ivTSm4msU6YfPWYF4cDBXxVNT87J2uwHiO2OcxtWj47QrHAukhGdMSsEq
cKmOjX5p1EJ2mpIGDSCNgkxTCe+KFBexfD/JnSfbVQDufM653iQ+8gN9EGZzG88q
wY6yFQunLaA7U72Ctm/HoTXrZQiwvJSQzRI7gnqsDjFT9XtyrLtrJBt6K0zjd/vo
4L7A8zuJ7gnc+smVyvOXZaGlTiCPPpYDpBbygBO0Hkugy4H4y/BN1A/ZzDs2Empg
Ubss2chEoAAzFgz/+iir557Er+VVpTB4bJrw5JjJmT/wdhq5Y09czfuDXrEPqG7o
kKmO0gqyuJPxZQ/io0PUmYg5AaQbfH+Yfr9O85GWekAE9T5viplHHGhKxbGe41/r
Q2DPrzde2Y+WYhfFw9RHPs+J8nhaXw7CO4o4dCvOOpWKT8rMDFs9VaYoAa/I9j6/
ilXT56xvc5Dwe+6zojdAS0SYIMGXyhdEr2JyBZe7blX4JW18ZTXDgsI8KPHQYpiU
lX+JgqcS0RYpO2vfLY9IBdS28ZCwZGaee53cwldRXWZp0B7ZYjk2L21osrl3nxJX
Qq+dTPRqe73MjYG8DsUxHGH02k9HnwqzdF9J65TgbCd44KqOK1WSdIEwvDkzSGu1
UCh8Nrt3A+OQJVB+CKxOTJg3qWKff//Va6xr2CHT7rrYyPKNk3sneZKlMO5GUanQ
mgqECieI8NoWviGDdjWIZoo9B4JDMMMCdHnw05Gf1JEk2QnEsshnA6AO08Hcw6fg
bL6FdO0zwiBmy3phi/ZP/QhJ/4WhfhOV1m+q1pJ1cksMEglDWzSSYJSqnMry570+
ZYaK62jP62PPAf+thoZ1Al9Zp4Zw+wa4WPeTDb7FXZFeF0QtoRRv/xw1W0zU/tGg
NfLXtNSm7nwrry/eS+UpB+GUM9pt3WDDfe8QgZKEuN5AT+9w2ssx3Dq4QUMu1TNC
wI7j+NDx/khe57lCiJ7rYzCrprwtqj5KuR2JGR+sIvClvj98ftyfKW1keaSweAOT
8zo/q8wm5JQQzV3nqscEgc8DS3wrpbmL46hZ1pdrZkcXwFQjxMd0G2TTXaipIgXd
fFgOwrrLVdgxnXygTBFj9THY9k+NYkyK3QvVQat83WIsFJA7qQQE6GuIhwwcZVYp
Wgk0BBDrPGXllP+RFpLmxcnoFJBIm05CfhQCY+M/BxtnzLY+93+Gex5mJoCHc57H
x66j4Wg01Ga22m8pW102YQT3tc+WO/gWGoTkIUdKgHZMp/tdwjBBHmTjIs/nNDMz
3tKSCwOsOhJ+FEdmJss7Wo+MFZuDGTcLmYMEUq9/EFrpCnI18M1gHd7FrgoAdQIf
kNiRAGs76eLt8QVB0PGuA9bs5wUSBMqQvGFeUOwJZLAAtGl69V6Z1LE88dAD0RAh
PBMwKH4GxZitaDq0MPr6E20AKDkywWCnRtaaFilbLItmFI+bEXCnYPOj6JrsoPYk
nZ5Pr2ADDpXr7pk3O/bQvc5GWnUN6cTnCrLL68v6w7iJb2+ur27GxDzJzrA0E1Ra
zichNXrpMx9QMzR2rt1ziWsQx5sF1Hpzvy0sY+t6p1dTDkjuuMZI5TmTmLiV31Ql
Cuxc18ATglR9YgKyE7Qc4zx7QEDNsxLaN6aILEFuoo4Da6+RZflJj+Vw7jrW3NWr
XCWFGErk5RSInCtwp4mbEji9kF7W6kiMZNP10HP3IJi7ua/nGRSd3wUUXBq8O3jF
clVm9ZW+EeVBqR0qAkLIJLgNAtKBEi7u4FMO26Urk8YpGWAn5nv2wZMropu/i47V
xU27BAB4T3Qew9uREvZKbrHOZcGNshyzePg4kEKLXLV08uaLU4VS8yqY7feg7Fz8
SRLZn1rq7hd73TPxFlLGbpaDb81HNEzpdY4qeCjjZcbJZz+nJin6j/42p5cliRI0
HeqRJjtaVX+b99aXA6/9ex7ylOlCa6p1UfE/fNxAa7TZZ9WLVRe4lDnZwvQm5yce
q5PiLLrC2Qyh1XjuaknQpJrgFH2Fkzgwtqm0oBhkSAIFFixeUQWlT5ghF0aigBrW
Mje0X2i0Ha6V4G3fU0/TholkqSFLgGplhZhRd4/tcuhu0lo9lNZjnYKaUggDDNG3
O/j7NKDMbClrRpYSe/kaSw9d9bOUjuf8nQm/tq641jCGGrJn4Ctxu7G/iUpMfI0s
4BkbDq4DcaxkpeqI/wfxfH+LqxVaX4eVoKhjTGsxCimwZBOzqEB5SrR761cxSlq8
Ph/vlLW4XcTJWu6quNLoZ5meAFsDFShvIEDpOWfbQy9Il7QgfG4MqWp9uuAVH10w
ym5WmAKgAVaPj6Qxx6dlZbJleiJz366+L31qsHqLXBp6IKN7e7YiJeiVjvcxhFkC
8KDvElJzN6ndULVCgr1DWnjcHfEuTM1xF9Pa02zB1zArLQO5tUSNCNTEk5DIok4c
e3xrnVVzKvQ9OvUc/Bl2T4Xr4DV3cmLmWqoxT2qFUATKi02Dgk1x5+viMVjROUP9
Y2cyFPnDiunRvFP6fxUYJd/FpxiLQ//b8H+uxX1QYWgcLZTupeuLcDAF1klo8sM7
e2Ye/rblV1MH+YZJXPyZy/3y23swb5UV8Q35rKLJlrfCpkTfbaY8M6sF+K/eOPHk
cJLXOFq8002b7I48lEbmIoybMiML4RUC3BQ9t/QiNRHpaDckToOFJLCvrmK47JAn
TRVGGQS6JnaC8ZfNxKZ1iTshKpDhjzcYl4owrqYaYMx9jPQWGkhbkMQOKm/Cesbg
yT8RENezsiOxjTCddr5ME1vXUoj9y610AgZ7/hFdrxo5UUW5LkPfEjtu7FB20FJk
jeNBypCUKVz9RdYeAfVqs9kCDcGxDvPQFUqUTC25+972na/cXtTBSUZdmcGgKp++
MLGgZXZ9XHmDX9yMhWT0VF9zpufppPXABKc8xWuOwYtFFSB4xgtVB/aXvLJbN6Nj
DUpX4efuoTlIPhjDBi5+fx6soLhnG+T3YjPyC659d0q8YyHZ8ZotpEE7pHjbNra7
fSRMDks7udj5YWGxxmaJXIS0pME0ER9b+LXDN4CotiSx+2IfJ7OgXGIL3WwEODkR
4Rubxp/cFQa8gBP9KPdOSH4/R6bOs0DUsaAth9vBQBeq8OtLqxGvqrnhO3OVzwgU
0lHN1Q/eJXc6hYSov/aFpNaiP6QieMCEg4H102YPY+Apczr0nyeAxA2Alhd6zChK
/Yt2whVibTSlKr3F6UrK0vXwQSuRSZCLFnk2zb7QvWHdYSyULaPBM5bUaKRlmkvh
Rmbxc8AeyzYd8Z96/Ffpq/khtv0whMhdMUt9hOPWDhVxTZdZBjzfjCj9oP9e8fBI
6JVVHjPGINkXx2WA+ueretmgBU1R4gE/PbQiRAjlk4C7GCB2Ca1op1wYCNwWWx1u
ZorX4A5qu/U6jpBv9gyVP+tolLd4BLDcSierXTHlRjSz1/n3zBo0/wEKx6tqWlt9
a0FR6MH7tVJEjJqDxb4WyllDINeXO+ugTYUTJWn3zngmDQAPNkRRHvry5736dpPX
T9YI8IYw9fhE5i5GuTIWO3FIpOsVey/dm3p9C93K0cwV8j9DHKjNHH4bih4oW2ad
fg33wI7myPdosNmAb8CllTuDAIyNctCu9CA0LtjZaylYm4UfuIRIfUJd8WRRPAez
pyVNE/JywJ+21JtAAgKsZXMOIDQEpA7+bYTdLWx6A3W69FW9DjbiR9RVREIOqiv1
NyKjzYp+ZGkjQ6MkaLMMBZkMPIX10Dx309GWLOUQFbtSnBesS0+akW1JSUj0lKDe
L1vmAbLzVn0M3N0L3Rf4OPEu+9dr0tGPhlbPYQb6TGDGRP8+wLmnuJHHu7PhFOFv
3+fkXInqGpHqwMOI/4zW3m0C8L8eE+qcJ19zopSmrGT2LmOoB6O+pRePgIuxK1v3
1bb8+Z3YP+457MHCrPCbnazMu1dQYFq6JEd1KQyg0YAbVUPuNevO5I9CVRDS7Pri
Yx+h1XhIVo3FyYrtRew9c0LxWFFeIiM2q9YBytPBeEsxmAX5vHifAaJ6WemHjEB/
5EwaUOJCQy1xYFeAmgjEA8Yf+s+RXLPUi6kYnWBRpMvgbFJHnoxzq3H8TBtDei5Z
qQnDkXInxOfFVgPKeOsS4240GflP5YHLiowvJS6DsB5NL7tF7KaeVfhYnTEbCET2
vLk/GZlPcrT+4TLvYqrGiFwt37zznZbyeHyiIX2Q5u8bSZvMnr2oSWhVc8Rg9yuP
LjmbBcGyKwvhhAxG1uyc8K5JAcIdRWEtjMJamxuWef7AjsXE7VTyt+pTToLc+QSf
cUnDPeaqaTrXlZfw2VjzgnaEPjA7JXOVHy7Qtfwt6o1KkkTMxXICXjdESJgOna1E
4E5Hlb83cmMu0SUj+U/Tx7BOCrZ65FAvaP7/sKk1iiV/Xk6umOrUbXPAjPtbgJxt
CVv66svqP4wpRnlOaZmcvcXFRMBQtSJKh6PlWKMuTUNtx9egzkePCDjzaaOtkqpr
UpajxVesYS2+i7ZaLTSISAsu/+PSAZLftx4U2PElLCPmx4rMPVkybNRDy0OIVC9T
9BPkshRz02BgiGIOjAasja//Sf+q8gf0ufH3nn+8nS6Baxo85PbhbydOI4qDd6DM
HreF4TUk79VwxrYhBVcwKqSf/N1Zmf6+nhTMtm7w4PAi/wwbIMJDLoouzSBbT3EP
jAWGHM56RfICvUtA11dkwdy7MIYrcM5aYgM3BCD3vZ1kzQIgz57Txp/J1RMaA+Lp
ZyMgcGq1k+v0jAvSSDzB6aVFCBTu1C6NiRauN6+CBu6zIxnQOoILejBhnRe2fx44
KgcwpT5tiApePG3wIZohPzSa9mvJSNBSf8Lt4UkcXUuZMPPZb03E3/h2NJvYsIh8
SVRU7XRBGmmSEVfCuch35cEeyd6CY8hgt1ovBKr1jdV7OysKfTqFpiI4scVrFMth
pERw63uGUn/clHeYMo1Dt7ZgiUTwyzQFoB/LlEfhgE7b3j/PjiKz+dkNeRG4UDNY
dStOP3BRWi9eGASaCPvPjrRMnGIxIvdjAv8OrzzxR1zbv7SC0rH+2qSzAWoSwJRI
AwdytJ/CxQf1iqq7WDGB2DskSi5J90D7BNSSdNRByjjoOI7UcRnZurKYtxehpQaA
86piUjk1ykC6gpPwDaDhoZxh9R0MXtJ3GaQT+yUy53Jj9JFsDoOTq3uLkARCHqOR
4rbBiXN2Bmpa/q+qcLa0JcbcFcsb8OgKBBm0CPB3FFdqZ2sxDotQyzuyLGBXkdbL
QkY5KNhWVYuca1kmZ/BxXPUeK2epJC7x73rZVWeM22ninGi0FMIViQQkTJQx5Znq
wWxslZbJ5ys/RMnLqVLvUv1aH2AQmb6heT6wnl37Igi1xFcSxK578I3EMu+JgqrO
YPIwzuE81G3nVZxL9nekbRisyczTZBOmWVHeHlHIoPA4PTXL4CQybsaBpRz8VGJa
icIBN9kbtxebUcQ6dDRhkeen4rmHZ+FDGMD6qXYoHMJz7i1s78KhzDEknozwKJav
ssx4R1B5JzHMM5rJWEHTVDfT6iXkrVknug4mJqM7t1qR852z8mgBSadMbQSPEU8h
d3tKhmDrRhA6LxqCjDoMvGqYxyErCm+Uf7hYQHeHNIClq5rH/Sc8yizUsdiv8s1J
Uve+oVjwzC3032XwVJzRuKA8Vo68BhxZO7dWNeeHNgz184K+H40wclH2vxawA7uW
og6kRS/mD4cDGoq2Ir3zgNScn35UJ5jl1/zUpqXLkDX58+/G9v2j+47rVd235mxZ
tvOEgsLoy1CJXR1NUOiJQPjOuCotFhM3z1trkGeUz/bhZTTveiHuQSPHlYqoKZSZ
tGzzTtiR243lnZdiMkz+MVCujll/9C4KbYbVzjgreEoh0qMPHntnVxsGjR6Uet0g
8lCStNXcQ1w7EDVzO4blyY4F1Ry24JCnu7tjqmCDIY684f7nJqq5nog2UlRlZu40
qsZ/36XrBPOoRD1f2CaHyjgv4QzNlhAYmO4zeCBPaEA1T8XobClxj4K0aw6Vly/D
r0Q6Ba0BMUiIkqoPMS4fzsMyufzzOy7tXA9he2en8++LFas4dfSQK0tC8yRliecE
gF1KPw+6AO9frNGUFWNWdApkL5K7zebL765KUnB75TtMi2/KnjMhD2IPbyxYw9q0
E9cNoivEBOq0Q387nUGZrSPpv7dMI+9yC92KBhhbmKs/KZ+XPTG4KS3sWvb4sCCL
vkHrfmsonAEH0zvJJrq3scnTnCQzxhWwaup2wXv+6dJIpKFSxFB78ESX1uK2lid9
njej9+78WN4uAFtQZPJ1nQbTXCyxjtWFInBxM7w6Gc+gKHaVa0UI+KgEP/QOFnVt
HKdshkygjSd5CyEg28zDYlhbpDGqNFojVzqD9bH6auUgEPMEpMrGpxJtmiEwgu9I
BJSiHAuEGnXN0mOC5uejv5TLcfDxfy1XclUpyAren3ZvwkKDNs/eESV7Lw/VRKa5
rw3BNRIforJh7Xpr0I5l6Xe14byXYuzPG9iQjaQ/9TbrclAUh3Q7Kj5CJIHKGjpr
wK3TWpncm3nlwILAXj3QqQ4PqKomOB2sGHEpK5Ep63dclrrkp5vM9VM4Er4eDhqk
lxUgsLLllBYGhDVngexqty8FMYqcI2Hjg4hXZWQvLrKgvyDm5U3kZPFap9YvPEdj
ozndw9CbFxUDuDxg4nA3dgm9GDFo/4HcaTRop2rP+J42vueKMP45hLzljlVpJIrF
15NpJFy9pFGI/+O9bn+qC1/99ryLDxGq7/mvfTPR+ZmLE2i9w7Tbhz4QCvze8pAy
h94VHarnZSUPeIB6jVoOYqb0PX+O4nQ2X8e3qFZajESaA2zPkWWVUC/dmuxWixkO
AGl1qdbFfNsJmy2JEBN5XPm3bCsBeJ7NmrIjN0SGE6bvuBA08R+0BT5JWyrWlMnL
wvMdBPp0FuzpKvDR2y7xrFCyqDkK9+8/THXLbo/VjRJF9zP8im7BCEtYRXzMOrXK
+8TN0Qg1GEfJSUb0sQjk0O5mftQBqIFyplpZaA4KW0lKh098fy6DoxGetcH/pUQM
0YvpFAVbTDtxxxsg3IJ8Hs0ixElF2iZg8Sos0eV77aEFVHz6MGMIDjhRJlrR0/sB
NVllLmnuKydGmLnh0qwqlPJmdFbAdwWkww17wdbSHTzeJRtXaMbE3hZdCkxEy0mf
LbZbGVPiIfr8nv+4Go9h4fXemNX9egNCtl7LYhuPWe2iWyfi52hRrG8+X053QSsY
reW+vzDcmE0/AW7f0ojg8EsL4+aAQJpcazbuQnlFDrAhznez3SdFU+Cl5/MW6YpR
uqbVEe/njhbPtxNvQTjLaQ8SzlkxTjwg+34sJIkfbn6r2Ld/1gVavCWGVYTInS+X
tT1tWKTKck7I7er/WLu5NPQ8XVMYqNU4NY3pmphAhfjYLtHkVcYdPAiWRIMAWnqA
SQbgRbcpy2oY8zZX3ewGjswpdczXbI+5acfiBNM7Kft0MDJh2rR7Ae90eOAfQBG3
LdrDCsLWfjpvzQSAapfXSuukIaHCAkYq3xVM1hW7+3VozraXDTN6FNulQs14sVoo
97miXraICIoC1u+tDYYHZaH2YW0wo4rvJlwW+84Trt8Lqth720BefuHLASdHt9Kn
G6BwW9veqZ4fT7hQ3KxCyAH57ZPusATS63h0sAt1mogtayI0jeDISGGyGTt6Gi9E
15kcxNc8+ALDX1mGkvnBRtDryECal+xUzewpt09hW/nE5Idvw0RYHL+H3vHT7i6U
c6QWO3juIdS7NNc9TSF9jnQeyfpg5Ty0nbxKM3uhjUdCUCJZenT4dduh5Y1fFwgf
r1Y/NgzHByEkEZAP3YCx9WtVHdftagiKCQWLtHmL5yBz7w73Rnxb0aO5MFk+K92M
EMkDTKZHgRfgmXJH1XbRBTsqRG4yDZO7AaDGNOmAYOHWb95ir/WZy984kCAXcWbi
hCYe9kGySHfJESStxPguKlJ+WmjQGMXIDOSUBX2twbIE8MPtwjysgdw50YnGD18h
SKWHiHHvfIGOEsPSWn+OQQffPYQ9grGaXZK3nLX/KICJPaY16Gxb2rRXtmOd0Wtp
xRXepzuAm0ZAD+hsfhE/1ZZ/z+LLn0xDudTHlVfEEybvqN+XtWGlTqu6LXTjvN4Z
XrF0B3QY+OJFordGpEC5kOHObj7FJIf+dRaTnaFxLyskgCek1v6vhLgabA5WoGZS
sJHs4RYy5hDcMYpPun4O6O/fnMIYLP/Qsd8NM4EXeBbqhyqkKABvJQDVUPW6gH33
48eXeQtDuUjkXt624ty9RBD3pohbZ9hFxE80bJuC7oLOhznD3VlauMhFaMbNJtTX
1IkCuYKXw1qOgEBwiOf8aABK0SHOlGC88/6TEgshF/wEG8eJm/cjLeLg19ioobkb
6v8JTmgLVUfPqDnUtsjX7wcPV53h5W+YKnpEyRfs/W/XrAMq6uwQ48aJaqx2jjjH
ICiLfJyGTK/ooX0qzIHsbPhmWok6mfsSevucm0+ALvIicPAPEdIjqrtoheeCkNMT
0BjnyeNPacX1gNKslDIUcVKUDNHEbX/QtNcShzDbYiUcAZE4AfktbabpNkI+EmWJ
Xyxs4qbbzlkgy/dva//mrAlC0TGG8glPkEehF1o4cTq6I+DUh4DtzQKlziwrqqVL
i41VlYnbmvs+JgnE/ImXB6KcNYathV+EAjmXL+f1fanfn5fzJwTin/EOkND9eRDR
tGTW2jHjJG9oHj584cs/a+SssAi2p0Jsguj9e4WI/zlSUDNVU01fYmKuPnxHvhGF
Ez/rHH1rz9z4aPHpY2wrQc3s9z9P1WzN/CnVGhmYIGIQa646gZIQd+E4EbJUU1ut
GbYpvNcQTGXM5Wu//4VZRY1kxHDmM0ujhj061sfcDoHEFujqP3uz9A5GHDBcBMSk
bgRoPrWz3NrveX4JJFiR7g/fbrqK2uk7loGH/ml4pdWzo0+XNTDar4GFhWXYGnIz
+V8CJQBG4RA94JKsK5LhJC46b5sjLqd6N8Z9C38O68oYUHECvx1t6mVBKtGmOpHO
JGkAUpKA3PvgWcBm6u24jtHjVwJ2RdfmB3/mQ6ibk0QjWWfdM7mtbviD45yuPa1z
n8x5WCjNS9hnlOESt3Jh2FnqlPbqsL9xBAyhDQOEgcOQCtFll1QM9Sx3AYLhiB0g
p/wwFXcVAJ8wuREPbib6cFRNvndbXzUSaDw2LiTasI+gSKhv5FyNXDYRb2ADU90T
HSyhNoeN5Rjys2KywCTn4K6MQzwBAGm6gCErJu2q48VktoGvFRVHxprQlDnfwBOF
EfkHjiROeIJgPJ4R1j6IgVK6TSLrCiotOf/LQpzZlhHW5iGavPQeUw4NUEwrAzzi
zOZ+VX7fd3iw9uBgyoOd72omqf0XRp1fCsPizvI/lUv4wz51Ut9g5GnOEI2zKaio
v6X8Y1AOr1PS8i/5ZhDisKhT9KZ9b48PYqE2nuwdai4ByxzcrHQDzo8LNY+X4QaN
wK5hnZtKnWsXFS0q4/0hPi+fA5SBXhjBipb2400MiNTagqczWEEmWKTU0Utjodej
Rxw0HRBhxcC9bDmNQLgZPMe9EeA/yRO0/nUN35BXqRiaD5Iwn/WATW5Pl5xIjDPH
lXofwfCuP1dBpt23Dufy1d/95p6jbpg6iJIaj12HE1rZ6LUyJ6RSeplxJl5RuxpE
eUB8A/gtdKxihS++4XbcFM0xSVg25GTjv1VJAF6fMnRgrbnJNogmdWx+6scrZng8
s9a3HpyOWWsxyo1NR95P2Yxs6FI1vELpb/F/wjMgorfzEvKOeXTA+IuD786LgYFL
tZCR6l3MywoQMHjgR/BllOdVtLMbLFQUWzPt6NRQrRqVpxgHPr0HoWzjmFx2vYiC
nte/t4SxDpMiKJoAZ3tUHhfYTHMx+013Q9Q1DCA602soDCx5mLWq8oIDFx2HxIdl
50ETp8okPTNWgEwC6kKcm/i9cRP1/mlpR6w5zuCISnofTbmO7MllEFVmHVCTJnud
VV4wW57g1YHb4K9l14OL2oE3je1EA85+reWq4ddMFXpv/HjU/+TauKEPjWCcyH2C
2biK2hXpiws7WKit+lEyywC/b9IUCaGyf03eMdhqG2xv/ZEdNA+GECBGJa9UE+Eg
u4ffbN3CVnAFI/22C9sg0UB5XYv3+YQs+AWp45wnknkX+vmHHHuUyYVnvfRdwd73
Z4unUt9DjsbD2LpjMwc4po0xgI1WzYedxmbMIYqfPWqjN/YkJhHJpmCLRXvwyHRl
OezosdDv6q5U758J7I9b6FcMjo/9+exxfAnFmSSzhX9W/t9VJ3Ua6d3SqnBZMZb9
zIBYHwvEjQWbGgfj0UMKhOIhGHUTV3f/b3YPD4mUSISe0Fz97mDr2Ap/dppG0V+Y
akUkrEgQNy6dNl/JZ9yakb+njmxbvOjjj9JDW2/C+5SOF+q+YCGJQ3pPGkwb8DFP
W/sXKDIqeho2+r/+HsmBTZZNbXFzVbJpv1tZvCTxe9GtlJNro/PLW9gKYutxhv5G
d3PIz229ouD4AasCrMUI2p1MQJDuB/lbFAsOD3xwrc2g++JiDcTnld82+lpfldRj
9W3fOYZYw58uXK9ddEgwFpdlMDP3YhY4Jzjn9aL9wW0ggEUU8iZ0vBOKfTbCKRBP
HrCrJtAzwrHqF/av//8CAdI39GRSBJjLJqPeaGGqkHrb0Ok+dCcSUD38i+UXkTx4
g0FHhsXR2q7eeexHP54RqwHuOHHr+kErC1k5gR9zabGDB5nvGuZLKrMIBRTbflNv
K9SZPY5OsrP+ai/XHK4NGhQboRiz7r81nFsRpZYUuPCe1bsmo3/8KNwG1RXpuBr3
jQaY9g/eOnPXGTqOCL4l8F0wdZsQtWsVTGnp0MMAX3MKpDLfqEBuVKBZ2qKFQYTU
haXkHy2ygNU80SId+yevWQUWgYoLlRE/N5NNOjanNcRJGLItoiUFI8cLkYqmr4Mh
4J6JYplmoK5J2kJim3F7Ez/TCE0pMsIRmYuPEJutUbO9Xj84XQMxvPHTCUTfmhEN
OPwss8v4ZGgKZrM4uI9ayWBoPS3Yh06f8QRl9H94ZEQkkh9upCh6P9jmt5kpvg0t
dDtEYKR/KS6lPcEwZj+7OMC/trxnPzX33FLLX15NYesV84cMpWfvgXYcyZLF+0qk
uUxYQS6tBUL9ZQmwQLtwepneeHoBIbLiqF7wCNzrbJ6PFXYFSm1hPP829wBNS8ep
oyD31nqR1kDw9Sz/6dSU3IwGaLacuMB+66Fz/DwpXn9W3U46AKggueFg5X9dW1iJ
WjOXhmR87emjgs5KjV/aTyWGc5mBh2K2iefldb13zb37EGXaDeZoig/0tiW+CEiA
Yb5PAoJd9UbgzvGSefgwgoY+GNKborXiQWTYNjBYNBonqSVqXAg8gdKuv/hBqqAs
HL7fh5vsrLKstuz5LVQCr2NMcyR/Dc0hrUBW7FJZdsAKzDUuR/Bfftvy93BiaIko
ZogMJUWs2jPCuDV5dwNqnBtfMpCN/TmplFS9+DIuFg+VcsnLHQY07BTACR8jvmFT
6R52ViR4hL6sGmVL5uClwdSDivtNLurTTiebpPPohmM1rReKvQAj1LiBYY43YCaS
sqSLOnx6zyVYKiv3fRkEYET/JiUfW8zQ+OxfdWEIidR4ugXyoDiUmnIfzs7nuUF8
hWEAMGAu38TRH+Za4Rd54OgSt1W7kkaLAgAEUAQdGn1thAsMaA06jc33xj1wodKY
5cAIrNxwfWNQfHRAsLmuKXyfSNqihVCmSdr9RJjeI1/g3ZDLm2RubONXC1X1kmVj
Tuqb07wl+xXw8oTlv4WHhNyVy/TQGQ8bG8oH41hIiSIeg5qZLkVfd6jeXb41qIVK
ndz1UmUPwAVBjlFQF7FMncqVPvI1Q1bD+hyL9OfR6gUVOXJk1pMUri2EfvRKGi9E
7S6plnkGm2nLUnRxUl/BeVdAPOMjmSh8/Iul+c7QWjKGxAI4V2rYom6WiUcrXv6l
oZmNC4ZpVsfjc56U3ffG4D5F0f4YmrP+91qpbnCp3HZbRw5vu5blLh/hK3HWFWg1
JFFWKQpiu1/nfacmCBsKq955cPIFQo41LIhu4UmCwx1xte14EjeChvdQalJ3ob0o
OBk5L8NxKSzQ2vSgkyKT3VcfVXB0R4758JjWAqe120e128gBMqMGVwI6IyNztkDx
sh9UYV3ljbgUPOudbSTrYzR4BNOY5LzYkcNqmvC8t1SODguz96mtrGLhPCFcU0tc
PXJzNmgEnFT4hVoxl2z38qS+k7ZOtzEPP1eUCrhmwhQ8al0L6WZkLOW5qEbQiEYM
nJrGE7sAOncuS/F73tCVPe0rSrLqSrYfb4B9eyloLHuh4r5/XwyC1t5QGSnVjYvA
MwYWO/iBIatSCPulE5seJEB6pziAMcIj3o6uplyGasGbzYRT6vz+FWDG3cT+s1ad
4jtxT63fYONZ1dWyrQzShB1va4Dg6S25isvuieu+mQhLevm7YlprG1MLLaAwoaha
Ql4kY4wd1QBypQqLXHO466ktJQ5VMu8je9MCcJZXtvS6uPIWUcn5YJMfVzs5LqaK
xLkB1R4oehpSEoTtEzIDJx+nDyUyVSQm+FDoq6dOPa/lx77x3mWfPhk36KWUqadw
YO3h0vhtWhbHG+eXWKhtw4YGU9iTOtPymp670HLHepkUeeDeMWZuVsK8e6A2wrM7
rooj5d9TV0dELWouBatIaozTZRqrWo6ioPCOvayKeOe1I1kXetPE+BH60JdOtY16
/aclKFchq5goZz0cfBuqbL9UW2LDsfpa9TjdnQbBeBexSmQM8wiEhZCBAeqH5cHp
6zH96i3GdhyN4IBH2tZ7i1bqCI+8srTnkKsd0EtB6Z2ZMph5KCf7gwJ0riKDK3zd
bORrtm2olaMjNpxu5oCpEnttmcrXmdxmS6nnjjmyzUJVH2mPcSlpIUOhWI4WXpNI
qNRgvTl7BtirFK0c00DTFR2tJs00t2rIeLISHa0ChfaRQs9Ri8BKGtBnMch3p+4+
h/+PjGnIsDF2k0u356fhQ9EiR9zYsFFXlYkjIkEGjAvU46VQYzwq2a1cwqFytRuh
LSWD6SFUO28nmDH4ja+zlUj5MVvHtA09ZbXpde7y7LossX7oo3xuf1y+Dsaqqg74
wyBz6UHwL0lQ5JJvMwY8GHCb5sNGpPCsHUiIigbn8fADjO2F4ue+7ZQOMKqqvNqm
oawNGtDQv9sWw0JvUD1MpriyD+Fk+ZcevY5u8GofLxuhRCzvveKMqsFN6K+7eMc4
y6LOhlRB2h/DqlHfkj165gwliwzL2nguo6CC7jElhVKZLd5PMig1bjvGFizpoQ5J
2OFarxpxilmURiJXKtrE25LiX9NklC75unNiu2R/DHAkHbBTDe+azRHnlblyxQqb
SYm+pmMRbKpFzJpkN/yixSIMBnEu4AxKnnjwIY2kVbB6b69ncaGwqj3y9201yj+M
x+AdarIODDvoYX4BZpwb8pmRbhPbeiXdUEHsEvNOQXeYOgXVQVu93oZri9f4/9iL
LsKFsjkbz16Dj8/6w9iXvDs4ydcCK+x94UYk3OG0PGwHGD0UhcyKRv3Toz2cdRTY
7Q0ikXE3P319/bEWhW48f8D15HrKlX0IxAfd6BuMlzKjG0SkpgBmKwG5bgwFa2QZ
Qn2YLktDThmohTxDcyNvxIpzWBcJq1F0qwEuuuICgP7MNN5v6ww96lMGZXA+ZbnV
1eq9913of8TuKTPIq7Mn+7QdkH3NefYxitIg2lVt0D84340wGPmeI59uCr11K6F2
9bnTh8W8IxpVjXXSAIwancnoMdNDHYeYRznt5L4IWWot7ZdLJz1MaqEle05EEa3n
tiDhcCljBb9+HO7g0A0rvxRMn9Hp/1g39TXI/76zb/OGvNPR9K66YoQsT3xe0ERV
/g59zSbvz2ynbUoNX89FmrvyHeCiFM8lwTMcytnMzoWGrxr/Rw5CXlwnxYgs2Cp1
SIiOiRHbsorsuK3pYgg4JFncwn9TtwMm5d6a9QtCAYVy7WeKGQI4uNjcgxG8eRSl
6eTReaBCesBDv/bc9p1NhCdOpMG2v2+2tVljb4G4kDPbyZcdxUrvOZBZlfzZBIhD
/tUk03EUPGPXMQBOZIqkLs4YW2FdRoqNs8mhiNrdufX5asS5pZyIP2iPovXBPEu3
B2c6WdyZaJbQ2JID50AQOs/nYc9K10jYQ7QrI7QXjaZwXDDHPlHKRC9sZxpGDpdg
smT/h253BcegwFZgMoB7ZQ6LWCkJQM2pBsOUFm0wHUrAP44LjUCLpsMOyv8tPh3j
NSx+6FruXnW5mk04uLabJCxb763ytOqY8TxytCUInsSfrcPHSKzwp2aGmq0Aav3M
VMfipOsKzCV8vdt5PIlx/agFTsqya+EBSevX9Ug0OXUX6A5+04F/Ca9m9nT2sN8l
oGpPL07geVuRihdcwHlaUvLNEZcnUI4wVwbQuxRccjUlKi/c3o60G6V7FZJpJSX4
h4r7h1AL/zYHDtz7yuri5mAE3T1dxjPS4Yd1NZid0bHxWlePQcznOItfkJlO+4jN
ksS2IniuEXah7A7E49AR7ja0tzWRVlIaY88CFluYeSkKbIu4tgkZGGZ1TBmiBI7o
wPZtTE02HAWkVPmgcun3JcEsrfzegpeQx0V0TL0sm17hXjLOCpBYNlCRMmWqCFCM
aNqQwnNLY5mAazEFfmZM5u4t7zNQSBcoiU6xLjR/khXtqy0oxZmcGD6oRo83U/ug
qcPC5PTqw14jDO4CMdkaRn8/1ohcxqHq6+XNXh8em1cvxUIuJMNu3xWJbGhIGlZs
3j6ZvTLBMdG6JTG9B0T/rBT4XMgPCOb8gi39VDroBtgSsjkPVnAMAHLi+wfNiS1c
oiKBgT5Wnu2E6wnuqbWkEgVb8nXClLZ2AJT6PmbEvtJrStuqyOgNoDW8pLnLMV8U
4SxBFs7kUqht5rVzKf9FC+tPYT/calKCfNouulyIerYD0X2qgOR9ePGAf0YuKT2M
Gyo5ptq6CztOBtGoSW0b1fjEdsKo/uokun7hVu/clw4ltCGv9x4V3ZyIlVSa93Wn
wb5TSrkdROssRsGlZe2hPw==
`pragma protect end_protected
