// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
hA+2tj42iNALXa8G31yEhS3OZfsMRbg06epFLCjRsSyHDZ6Iu5G5F0iAfd0KTgtmyMDhaxNAVkKN
+6I+HblDUz2DfuzbvSXy9f/V+PE0N4LdUyWwWRK19Q/waZAZpsGzzgByLDPV1BQ65GMpT6xs6MFV
zJxTMQLtooDbXEMk15qBGlC2HLAvZunflTqpjoY89KrNVXkjQ4PlV9zH8IO3olxkygA6fxrJnD44
exfQIrEaTf+ZTxSjmrwAu2KnrSqxdSBliMGTkz3LsO9kVA61FYXexc/IGv4lhAsvb1flEz7LyzGD
OkJxfKO+TuOwHFaeh+QHSdyiem2p1WPtVByPNw==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
Q79arXTSKrHYBgQPWzE49KRb/XSGlX8DocJnYOF7YZk5j91m2zYIGbYY5K69mf15miNnOrYXQV/A
ghitGm5qbY7velpjW6IVD8MSy70yKZenk3afY/bHcghkW/5avNSXtfr3D1I67L5xt49rIlf3v8AZ
MaaGd0IQnLsiKvces/sym9NzgxZ3sHJOgWx6F7uHQJl/dWlksc2saofZKHiPor6t1RcqJ0Y5T8fe
9kG2M0sktxWhe3ad3OlpwVXEXi1FCuj1JPxaav3Tc0nkCOTYjIcRXG7Vs3+1Vtol4p3AUowsbBa1
juYegEFcmYu+zBVZVo5LGeHRIKNoG7NTeKVDIXUNb1IeYK3JyqPX14PAic317oMktZx+351/VWTN
DLJmoQt2xdLuh5kv2c36KBMOJSSWEoTHSmUZ+1H0w1A04Bu4JIZsnlHsF1CMCMfoBNCillro2MKe
P2SN1LTQHonSKnvKVZsKtv1I1SQeKhbXB4EVKtvQNx3jiwln7L4fKirgJOoHgT/XAmsr7uXD5XKy
NhucRqD4iuFv46Vl/0TlV9vuAlhBxWqBFfZmTRB63butQLu4/LPun9ojPxXk4IVSlMwjkdgIeOZI
IK7BKbFNEtIUEh/Ks+vdnmUnPeCbjk/zY2DqGorfSE9MbX6NNTSodKBpSPHIQuExj2BcymBGyznM
9I8Yx3SeBdqfx+eM8TKdhQfrhCSjHLBkVLT/vzAzq79DOxgOksmvIT3yGxPE+lJdwC8YKtPrp1fI
r7a2oN+ooDqp9nRSEMeFMfbPsnXFk9MGOMawVHmoISLVZcrwz0+gaImR1KblMKVa8QPvATBPYAA+
sg3bE3sHPDmMmKd59DRSoriq/kYTxsxX+4Zt3V5X+sIiw8XJkXl/UsC1/REGwA3B90Kjnvwki90w
G8meJkZrkMz1zBSzMRTEH91s4ogWqWAjjw7VrtMgju20xGuZNrbJ2AMGZKHppBcznnFuVH+tRnE2
4iDQTjAcm9hKrLVUWoIiew3pHlUYpKjvUwkHovQX5/FgMV4Gf573vsYpT7BmPPll1WVK9sNRvwM5
fassLne7JQbiOyr47aCaMCa0Gjwt2ZHvrQONmvCbZaI4kdB4QIKjc784o6E1yneobZLeS7RzSuYB
FQ+Q+144UX/IzePZOXW9e1fIdQ2heOUGzeI4IapDiSBIZl8bdKsMa77zmA0n6LB41TejHtOjlY92
Ah/4C79K5JlJsp+a8h6oXo7Hx2OSuocXMsOY+LHellEEqOdqdkYSBtVBYv8359wQCKz9IkTydKwK
lUTBbs3EHhH9neifmLkrRRaHYxv69vb744tV1BEUK4d+rvGSunih20DUku+ug9HTLLg1DNR/TB9l
32nWO4jAeVuQnnrMo/mmMYeHEvxlsZEBdF1Y4527qWSQeGZCCEGEyaVPdF3T4xnC7Wt7rE1qV9Yz
KDH3nGj6KbezUFuatp5HjgnEpaw/Q9rH6N4EwGF7JdRUIsd96ZhX08mQ0i3gsR+ze5uCL0pzCojK
cCYLZFQM5KD12hsCnX43rNky3KaLUj8IHfKMAUkiFxqtG6UZ2MGxGwI8a+PsYDPczl01om+39Xe2
xtIOFY3NsZuZf/KYwoyzsmJnQdspWsyLfke+ANp3fTP0uPduo8ifi9OUKh5sxE0HqDUGDUrQAfpW
qLE8o3nzt/Oy8GEbmWCIoGZB7jnALHiW3i4CSjBR5hAWlxGs0upOOxHJb2bcmTKKvErc8r9f3L9B
9FatPCHCqRF9L4Gzt0ees+jIjT5zIMGH6ikPqBwUx/HRo2ovEd+gjCsbw87dwX3A3MAc+8xCepJT
OAuEm+uzm9SyNz365BR1ODQJVSQ27bqE7rhzJd02hejVuxTn/AGMBmVB/8AIvH+otZNHFmK5Tvxe
eOO1BFx+XQedF5Q4pB1HMfsB/4+Qjbpy0gXvwT093kP6Pi3bBikU3cDA0J/GT/QFzjIY5QmHVLb0
JEaXG3ytc4a+727kJff6Izoi3zGNJnHjboGqGyO/7n2qXp2fx1lThLrVFPScP0+DqeBGWJzk1B/1
OCHaNM2pE2cj1rWe8EgVt5sFmMHmD+LhM+DTJJvTHEHF9VAvggR/hsOTXAkttRexlzklGq6fARCt
6yiWXigVbQVjGDxVpaQZBs8dvCtx/UrInYYwNkDyhI4Zf7X3I9jYSO4/3SVIi91X8oKzgTS/njJT
2T3++sgALKiiHQ7wpMzucVyziSmQVKjvn5wrBpeM4/Y4TAmR1be4F0pyzeYWghr5pOW2JF7601Ha
6MJCNpH8mCxJ3pVRpEyKHvsigeXmjbJWLdj/LGwAOgR0M4ht1jjL/UiUFEcxmp1CHxh+8iqhJG/i
R7mH2/YAZq2OWoRFKA0oNUtESO5O08VIjM9eFG1rmOduui114Zb4NkLd2CNnF6Hh8bpFSup+ElLq
fZ72V51Kdbj1zbaXKVQweW0hI7qA4VCiyUYkIi7JiA+sPv+qgs6i1Te1MMlo2H36eLohzcE/u2yQ
jjraA2HfNv3AGqjRZQv4w0cQZUtJno95a1/cYkx0nstzhiCc/XdXeBsA92Tk7nuCxa0Sy5HZx6ab
hB3G8EtFSMlDLhndNua6qzjJ0iUOEDvbPzOBmSGfjAyXBIqnfMpFWnlvqasq3dxtMIlmEmi6aasE
8WjKVNpOdGK2MQMS8Gzfk31zOn6jl0D+bfFXYJu0OLLMn8LJxoEohRddC0cKfKGwav+jL8s+yxKp
59cALlZsmCNqpxVwA+lv1PRJH07pBlTuXEOg/DM8thi+1Lst6a5WSBrb/YPSDHgiv/cnOUFfRYXY
C8wCUHUoJJfFwv341ABL8ZSuMw==
`pragma protect end_protected
