// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:23 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
QnydObjbz0LUKuuDoThI7Bk2FMqnMeRwST5vej6jI/SZjWMf2TJ5KIIwuY0su/sM
+CxJm7GwgoYKs+ro5vXmeLlzj3ApbdjmTBowywJ1DLSWPZL/RHHfleuvjzEKgr8c
SIJ/xbyZ8YoU4f2bjTytBkWzF9J3fRJ7bNa0KVqtz4Q=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 6832)
08mNewBMl6+gXSX/RP8Jaum2/ugU7P7In9pjLFaLdKfxv6umOB5LtcIIqvd+/Rqw
foq+Z7Huy9GfOC7B+iBT4nC+blWfY+yMHyttv9z+4K5ibpg9RJ+lk2UxZ9sL2FGm
v7hs/wliDidWOv0XUc3hiPSLjO/tM6xSNHp7PnX3HC+2UQucJ7Xh1Kv5RrqCwZFI
wUxYAcxtO+WhLUbGa64RaNGgRpyGmKnibeJoPBydYbLh4WG6aohVLm8J3bcijXZn
L4dV8Fkg//gjkPiZrFcFtvtuBxq4zD35RvHvW6nyiJSQlqdKA9Tm27OVSgpC/IJn
5xCR/GfSQAW5Y6vZUcTLI+np0Yg0BrTsG/l1Ea4+68wK2ItZG8DOC8M6beJ2G3i3
smvvaPCShf6YuBEKGzh26F4jmRLruDRWeMNxvgQK4TCBT1/v8VKcAkrTqMeidP7n
6dpSu2HzHS/FTB0BXbxVpSIj8NJ6QCMY6o2pPLQYsjOE9PnXkeI194Ije/Exwm4v
H18d9fCgAaI9s0B/hSTMAQCHlLcAY1w1gfq8KfptvEiPuR873ZmcnDAQTQzNSg5e
b/qMn7mvXYwVEbvDg/nOusYzqOJu9vTYpkcjoh0v3YcJ157e/qIsyuToExd4x5F1
g00u0hcbaC41EPp+wmZcF8X0CW7JFr+HCAam1rcSzD6BgCoftndoxj5A0dE30T0r
vvI2xdfXgcup2Qcmh0UAEjBmltO0eUrOf5RwUPqn0+jHI5JI3D2O3lODsSksmxhm
OqKx+X+FDt1+G9jCfuXlDw7rpwaQ1t4I59VRUhRa/SokIBhIGi7YjiUeEOiSXz9f
iwEvt7r75eHgV3exPj7+XI/3U2caLkZqxIUiDqJnfZerNujwRUtUKoPEIuGTALQH
vVBL1pisqojo4AMJenBJvnC8+7TwsEWV4NZYqu1WKh6KQQYnz5VdiHmuWjH8UZay
7+xK9QpHU0Js0OWTV4YLqgevNkiX2MU7sq2yLGJBMa3gAc6vO9pd3uDCodVmbhNB
UfaorHkPFRcxwtBALdZHqiSu6NUfHX5IECPc4b2ZjSvsfcv3YK1kOWOAYiG0wZCT
P+jrHdWjuXwYZ8uxIiSSrpZsUANrUgiA/IfqPZnUA3vgZV+cJD2ew93dCaMv+j3H
7sBEUiwVp9YrVW5it5kKXcIkOS87IfSGCtGXsCLqAr/B0XRLQ2oYPRERsetiJK2z
/AifZXQaz2fJl2KBYvWq/ll2adCB7zzHu79zzIk+eCbmiXoP7FSFXSszMitjSA7u
gzkYTwifE7AwcrtN+lPQhNkhOztB20Bp6cq3HJStkZttvy7GC9qRzL/noFIhxv/I
lZgQapn4Z5EFDNqM3smzw2wfHg/P9GQ+AH1C+JpfumayViPgFo9HutTAUCEEHzS7
iKwB2RnYLGq0xDQnLB+C4D31WUU0YExcnO9C3Y/VEihu8SCXB2tCgqob8xbjMS2V
9T2v43W5IRKywTk9Ykn5JN0HoDEeBGGaDvP3R6KATFHz/mDipsKzqxYH51Md6SNj
3FJTkgS/9PPYgM5x6iLPPd6UuUdfHuyvgbMHCf41PAs6NyQtzM1TG5dGJVrX+DfD
+wkHKBPg9lL7Ff+bePQOjJjHOkGpAqxOS3ekFPQp0TV8Gm3xY7SatKgbzMKrwQO+
QlFMHeP4Wdbc5E0AvapBxJD1Y31Blg9gQSn46k9yaqZX13/sz+UQToQkt5GZSKCX
Gzh8GPk0OGm8KA+Z7cq1T1Fkc4/i3K/47xurc71pPY9PaNxRR4ivBhRmlTDr2Imj
NFJaMgjvGahxZcRF73GiL6AJaf4HLhe1jUN/OgFPhw6v4GschwIcLBU6HW8rC1Qn
EEjnTtAp5IkWQA9tK6AjSrmwagkgXiPiwtjiKX6AaE/QCwETPxglpDk9dmm78ggI
g8nvv3WV9yEZv0M4tJdPKQKtfCvS5dy2Sp8/rvm4RrXwvA+QNt4IheBHX7VhqhVq
SJznDelneHmPy+sERthzk+Er3VOpk8gPgA5i+j17clKeoiDVkZfAfMRaEJiApsup
s70glqktShklhMQTaCToGldoKYOqLz7yQHy9iaMdRCvdDXFO1cAx1ACBf4WRiK1r
RPyUkhGzS+1yHTcOOCJE5OShkmcU8tCjUoQmB/3rM9et4iA/CFaq2ycNHYfClq8I
eMbBkmC+SuGPsVLl2H2kExBs3xbuU+dtTSfPbWNL/uAA5lGWhBdNeNQ+cZxaz393
zg6bj6p/dGMFxMou6xiWVV02fQIjjzWOJWtbwSrkavQfWkmdGQQcC+mw1em7i1o3
l1uFu58WP2oPXSFGpUXlG15RHBpaRZcCe2zCHDoL3tpPyfDM+pIAKFecU5+u0Pwq
niA6tfzl8abeR12J8yf0qb52rII/vy1c73vRKjpooVme7wR60zhJom9d1rNclfp9
4bLGjcBLXzThGFYRw7nZ1CHFnMS1EHpQx2lKapCNGeJN1/sVw1wTGOYSouM044KL
TZ0ZW+FDivnIcj61vIIOdEJuPHjSKkVMzBu/Bp0So4jx3k92h3l+yw8Z3Olfj/7Q
SEexFwBm44ffDq9UUSXdQfVSHHrEpMmd5Qq/LZlD4eJTWQhKyixL61a5qsUo5EtK
Hws+0jG9If5/vcsk8THGtftfgCsvNXxNPiEGKA/XmGzEC8LP2aAnwYK+aV89XdTh
JRgS5S/TUDhfAUxpBJlllgWG/d1FnjPVz6C445LbzRlZG9qJjFHGU2dwuB59s0eU
aOt5dIysEtBH/WaTdEbKFBpsx74tGGyZ310G1FdvndbwaSRYze8McKJfryxKcaj6
EJW0eH+9j76XpbBT2zUc/yldJKQ7Xh12p/l/hgMley760xL5jdGotsx8OJ1FimU2
J8vPyAWi0oGLWjz6/OygE6NFlR3jwFYWSdT7fkRqtHo0oEjVPkpA1qx2rvHB1CHU
1EzkSoRpeZQ7/p1n/4Zr+ObxMCMLz7tx8tuguIa6sw4ILzO2WqaHw3UM4wYW7sQX
K2WAV4BUnuaJWeo96/OhiPZm3BJk2Acgvf89XXYns1E6sha850hMgNZIWE0dVbm+
9hzVLJRzR1d6gjFmmFqTlpudrvGcwKVBWIOBuAz4QqVOWrh7U6eEmqhllwm+p+Pu
c8Lx8dFA0iLs15XKc1kwSqjA3lZK0BvSKOcfhGZBG39vRowrp2s06NF6LfnxRRHC
TP83KevOLvwjmrlLlVpuzhiSv5PUxyIFnISCXoP5Ut4UlhfooDDH4u72Jp4LL6K7
X9ZWj2++FV6D/Q4Oe42+3gbhCFS4t4NzqcG2ETNHDYGxr8SrJmIdSzCtBbgvHjc8
ClgMCTFi32ghGo1nITb8qIgowU8U2ejZQsOVotnnj21lFIThdjl7kDSAWFS/SDGl
kFar77looJlivOOmAuoOzCYeEXTedGvWN2CkwP3fU13rdvTQn7PUmBEAqcAdbKul
KfZiAbddcp8X6RWEiuZu4aoy/OMI4SJTEYAawO8nS6Bbq3TuRH7vOTUdOVfn9TBJ
4oPYq9rHwYfn9VfFwf5qHJxMaUX0Je0wycjW806kubPgdjqebl4MKABERUqr7qE7
alsGBZToiDscfY7QSIH1vJW/B0wgUeNX4bgcwwT9PejYBVc/OcniJyyIjjWysHbu
sHTlGRjEz5vSGPg7141vRy8mGBLamP43+hJJ1Xqndrs7kF/ENFjfFeIPqgbD6Yfv
1iOlD5b7BPnnAJpRlUHPf/6Ls0VX9MplWCytc05HjwaYv8YgK44mNqQ+K4Nj1pzS
v9j4qseR3nbolnAIf+jc+RtOAY2ZIieuzlvxnOAikK9USeHSBUT6Wv5rAL6izvla
LnmZI4Zf8YQW1lRc+lGwMU83Xb04xqJxOCrQbbe4brXTV92al9JADNK/2/K7to49
3ZgVDeOldiql0RhLMI74XixGUTiJFR1a7auHoue6oO9lXa3kt0TnBn+4urM7J5tu
3A65HlL3x5+K/k4YZo10NnV5/IXuSGxlLGX5TlDPLIq2dIWNOAfgnQ42r6pMGTb4
EA30hy/zH0SFF6tB2SO3Upx5HmJw9392uJbCQ7L3MhoQodUE/XT8IvDRZODaGRg/
/H55B4Q66PSRWo23LIwN+NYn9EPAGul5ilk3NSh0ajo1xjHUWxEdKLdE6NaPoapr
WuLYCat4zD/J7Kg7a51ZWUpJwSw3owPR6gng50yLRSuXiiAyu/ZS6h9chYTaWR5d
98KTOq56L7ry9bDFTb+IaKn6rL8kgZfW/s5bPJibyWhx/iiiAQcaomKILZhsdKpr
NSxBU69ayUPbw4wzvIbAOg2R6EWmvmwobW9KBfedfOJpuv2RubOMQLwZUn3plk4a
hIOWXeY6pALDo1jHMtWFMV8zolsWz/y/kzA+K0RpkFOwDn/K81p5fkZwF48iatwV
c+ftqiIoi2FWHVxJBzX9OqhpgtXpdkcuL++0ZLVPyhVbIgfaa6zfNM2t7xg1nDQ5
z7dC5Zib7A9F1nHrgr2gL+tFL+VVXKdm79scL4BnbEqza+e8ohiySBruGgDh+RID
O98367Fq5ZprnRlVRGV2RVzALfCegz1Rt/tUu6nJqfwSogdQQJt0cSsdoHEsYxjf
JitlbNUBjvZQ/6teSZoADqdlzpgSs7OhrCBh2kPr3aX9Yywo6JCTknfWTF0xRIkw
rPWLdNLEw0bfkRCKNd4XGfzR5gRTTdc2NUrx+z7Nj2btTkjaQYuTTO2h7pgRVshS
Z0jAdSp9112gtiswU+no7xlnXgbk6VdDQ/7LjDeHcF3oBE+I9EqaCkjaWq6SfqTP
CtBjiqWCWvdPWocAExgvzcfX/6TZGhNQZbfu6xQ9Posp33crBmfH3lg+OKMpOI2X
EvBX6IZdrafsvLbhf7Z0rmIokddzlVV4p1E8T/HUtZhdYYxkXtMulnMk6xlrJyvk
430lk9jm2LYmEe7I+RQsAjcjZGi5GrCAVoxI666qlapex0QfCsPZqRou+XFjUd0V
EcyM6AvIt6BD+S5I8Lzdut029TIoElddG9vvvXM4y2Ry/HHTlODct9yqBC2rceTM
b/O+LKKIQ8GJfbRTUrk0oEZ5cbLibA5cENSdK4XsdrnNMcMUXdb20dqAQJIhZfQ8
kA29E+P6FeUPrYr3wpjVfG9FBKbjaSy7J40tRgZAc1pWEonbXKZzNFMVMFVceLKs
jH6lwyA6ejXc14pvdHj8lwLiUww6g+WeSgXdhDy94AnYoyXgsE0LPE8eEOAKOTrx
qQEy53eCQ1BffWw99531cczQ0J3NpTr9C8NeoqryzDiOWchvziyqF7EPCAYq9CqB
3m+qzRZjw0IqgKZWnCcMzQ8dCYJJENUaYlOHAq24K1w2rAlUKcsS4eEBBKBGQVsj
E/bWxz/8ETSH14ibTw4wauEsFNuktQkIDdOhOMyZxyApLtH6eMnnd/0gAO7g580B
tColXCk4hgr+y1W1lKmaiWNbHQOf0Hk80YC2bUBA0ZYsC4GhlLr2AUhUhF0FevCL
ir5b++YEMYuxdlIWQLZUBzPlsYwT8PyEZgGXQDxcXZp0ueXYPqGpLGN70qHSC5m7
w6uW0/oIsp1v5N4pRNhu2kfs8Vn9Gj1s1S3yUSFTuBD3qE9FOjGCl4mwGtIEsEvl
4zrJKAoasee+WurYuID7Za3KSq0H/V8571StdkZ9rET3+KGdRwQI189kRmbWVQa9
PVaNvaZGRufs+ICHGv9L6cIXrOw8TOCG2F0YUY4XPC5sN9O6Lm5XZLqJgRFhWJTT
DS7gbevUSZElP6Edv4DkAea3UVxB+JP1ZZ8ZT8bc/rDs2aq7UB1873fxsdc4UH5T
hpNSnH//TuQO3lwTpe1RhebpPz1Me9/AVTkRe9blW6Yw4G3+InlQGpYcQFwOXKFk
F+jaB5ai08YTq8c+akWFcfaQk7VK/Y1so0t/yGF2JkvZx8P17qJgjafZdy6TO8pn
IGn4u8po3jTQmhDWoNVf6hwvSKuaCCzlbtgTpAe0+hf3STGhUo9fQrqhNTgkTb7S
ATD2wvJsghApwAixwjo0Msq7GEJeReXBT04kZ02JHBrngiAuz8CCv3Y3xUPdSR8I
Y27BQ/93gOwXA9TwPkeeN25l+PaqGMCmYjpPdeHuRQa3loP9XoQCdnCTIpdmKDnj
GXaCPO3yB7YiVfQVXAkSGMJ9bVTxGL6qKdVy87X00/4bgc9usQ9QvHvP5BX58X8w
vCkmCe57qS1hOdz9er+98A7T8z5uXsYi4zhSUU8hFnD5lWr4pS//rRleqy4vaKtf
6k+rwLSx6vApy9YERh2+qy3sAyI1K+7Bo4ZkYQDsfDVTF5hGyBJzvUjb/hnO9aCK
t6iRpNlNsB5nVsEhOoPUL2rLKqVPo3UHzz7pmj/xYKSdp728O0c6aCEeYdKUkwqa
RZJK8J0GqJLP5sK8tFqAaiDu/VBzpMisoup62W138IHHJvMrZZwEB0I2bdgq9tXZ
5xdFjoKanEOefPiywtLNJFmarQ5arbhy43giww4TNQXcH2MBJ+mmnNnCuhnjPnD/
sChFHVJY1At3n3Zoex78bqTmkx+vhow8TG4NsF8xYpo/d0DJRiQaeoe8gxIKKeJf
G23OLOm23eHBLfZ9+z/faYPEMED/+kBPUDJ3bZccLp1PU/RWl+vzzAd2KVOG106P
zV5WSVrHKXr+PSQ59Kq5SfcQA/IlzOFcjkRRL1Yx3EyotDUBQUPXgN3CkfJlhjf+
+N2NOohCstraj+m/mhUdozduvMqZhXYFKpzzgqOgq824cwimXz3hQlhloT+pix0a
VDQIvmtcIf1ibSvkiycfYyAGy69NwyqsexKX1hWhBDxsgtirVCa3NOBNehpNuoxv
M6SMUpK4K2bYYeNxk9RJWVyXxBTvEtiNQegW72d4uiOkw2qYoQaQM5NStwkRCh5K
sx4UQFKzN/xGwDXBVyaZvH6qQXDres/QWidjC4n/nSr26t1zowoFV18bddC+gtRC
e1l7nocXXZk/yuJEVReSrfCVeE+qXJsNhLIEXHLWnlZMj4t4MOZ2J6eVkIFDcHxU
zw1912/lGC80PjxkZCLuu+mw7+hlmTgga7FUJLFkw0y0irnp3KZV9U2uMFprwXGG
xvIHPUEoK152FEQ2DkBqwr8qrXGSlU93Jx7pVvGAlg4bClQdoi/rFCphfhNr6Lcy
2lcadnazSJz9ljWyiArxYMQtT1tFOMx+Yfr0hQI+5INxjnwtHoKWohUxTfn8Q8uz
G8fHPQnb9f6I/Qk7NLueOiGMn2Ih+hhp1t6UvFQUojy8b5ZH9LxE+I2lRARnHvLQ
MUE/zWaHzKzKlGxQHWPMWFXscl8//kfdjOjWspKNpz9VYHFRfoBN7LSmxSwPReAD
TKlZwjwe+qoAWX3c3/tLN6IGtbBSE65pTYBeOuyLL2RefXB48IdoqhvHQrT1zimL
Hu3nFoiRxVlq/KkAGbzNlbwtMGvdZ3yOv7IfJrzNJukPRSpctIbrIFZxbBzXG71S
xNbN6CMVEf9GpRpHsNEZLTx/BsYa+nV5J7exdJLQFH0xwaLdVcfKzzA3hSZAsJra
g8HREKzABJ4MzJqATBE+Pc+Ka1vn3AcPFrkQ5veHfntB5RTJ8IaNuRUzyiSckcx+
JvPBKYqgf9pXGGdw3qsWajldHF5qoTthfGEwrw2Op0PPQLUxuOyzSpwV9opsbVdu
A1cWezWOzMr4aQb+WsSVYvDDDDhNva14nenn9+2vWKWCZpagqZ0o0/qJuRLO6aca
yvVFIwYGHHqyNCh/vWF1rBmaNL/5BAcgHY9u4M0BuMs2UP++3FUzVS4cUh2/r3OF
GpV41Tc8p5URAPk0wfO8omRtNb/4wLbjP90Chq39vTz9S83L3hhpbCIc+3kmb+g2
hR1jl/JqdtawaRQNCdVYhI7ZsDbVmMnKje66JmbY4QJid7XartXxp3hqabKdDCkS
5z7wJ7nLKGUgg10SS6yxFyacjzm4yzPRM6lgz2cs4eBu67buW5MNFeAGZicuHqPE
u0vEEJBvcrb5mm+lh1bfa5F/M3UrTWmBfTuI8naHcevFfamGPmM0VSuKF4bDGBm1
Uvw940Jmh2OfCw/CDYk5eGOyNsKz76q8snnz/TNb2Z5cQK403nQUeCd7rEMw2Ua7
sf8mbSb/X8OI2Y7DhAEZIVCKXfhWt1ixq/ygkMApTXPMYjrpU59jf7Gymg+j2zX3
qC2ysERdaBYhvgVFiBzHcNftWxnC2ZjI2vd1r0mmiQAN/N3k0KY+tOTeLoBrZyr6
fWwG7lxAvZAUlHLUQtmPtHaZXaJkUgZMXMGKKY+42d038a+SyB69psEsWcmcC5+b
Veh8Dd+3pZ8vCBNP4TOLVazcFLihA4YpXFVTemAzTiVA20cjqUQ6ZbiJlHT+CLiv
BjsE/JFlM8A++ZCCb3ycMWVG8B++xoG9wo+9ckrCyWuMH+bStkbSEs5BITAmgCI3
4NdiXj+CrwKdtECLyMpSK8gTmEiLNmsQ6pl3lQdAQLfb98pp48Toleca/664GE/S
e4V8dnHXzpBRy5Iq5v2QFNhFXZrTcv/T1Neb0Cr1pLqp2w6GMRS2F/nFiLbXUVfj
Ve9P9Rs0qiZ/fwTKwGHtAi3VMxrz2kKTj8oGxhZ4lD4EjY7pLKML4tO0wkL9rWVf
Pcj5+7imeipkJaZCpclCFp1eiXIKT2BDWOuv/hx04SZBKtQyFZekbaVZdDOjQ1uL
q4E0RxXpTcMScO35b1lAXDVfcniQco+cZ6wz56oeYzO39U1y4oteW/hLhiylVnrW
crGY4yWLEfx6xIaTINmzCOaEyCMAPugnFiPR+Pd5DQdIeDfJN2sBgmxM8jTpTKZW
MwoKd1WbKh/lb4ylL/m3kJ1T9+0XGJNKpUe9DORX4thbH9y2gvIf67vjNNhnIMxu
VMjvnLmVH08e6OsUAcd8MfLACpOzP4XJ3RFgTwY0O4I8FT824+9+KwDE8Ux7Txf0
SxpzeeRtUoGd/5pt01TSPeoCFhhf06Rgv/agp48roiyw3YB8xFqdPZ6YO41KCPlp
d1fVgR+L79TG7Q3lrIp7lnad3bDih4SBuUJI6VFNKWEldIGZpA5ACVvK5pWYRGre
DULjPKw/nsgrVD/obgXoPw==
`pragma protect end_protected
