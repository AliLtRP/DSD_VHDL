// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:30 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
VLVA3O1P5E7M/YFr6/ZGNC54ZjR3PPnW/EgbdaL6LxeunnjfvrR39LAmZPX0/q9B
lldNgGyWCjWHgHqS51zLsU2QJldjEHinUa45xWrZMAVDf91Q8MOZW8qxMUYJg+uW
uUVkY1ktu7Nrjz2tEW44CkLSgRl9X8WEQ40Rfg1Nkrs=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5600)
02BDYFjn32hOIbGwhjlitJrvak+JuuzbpTr8EIDkgMw/R9IdwCQY0uu9yFRLY/y0
1TgzhqP46aXUieQTjlltXPho+GSloj0RWjDYFzJ5wNJdJvajUumqjdvyLh26khae
grAkwVBVf2afBIk52Ki4PekS2Q8aoH0dZzVIfU+HnU4VWuYGyvFcS1S51XqDMJBP
QumX+9bXkYGKAUfY4BoPVErfwMVi1petVEvg+wch9K0nvwBMXBIezOfvdCfoOUUq
DA90C3PbwWTF554PGl0yo/jur1f517i8CvIcYl0cdSfwpOr5YttNi56rYCdIPGaP
S3v06aGESQtSSFNgSgN4ysqU5KqGHU3Klux+VblfnFttdEDOI94x69jprn1j7s7L
OEh+tOr6wh/m158XFUr9aKdghIAtEHBDb1dji0clvpa1k/LGImhEtNyMnKEaD5yL
338sWZZqDCtu6pJWtO60H7Wwqpg/kgi6EB7CjBqj9A5Far9Of4564z70zPetD92L
d5YYowk8wTM/ojhpT8bT/v49tDXDImJXdUUF37PCZ/CPGrXYnsfFWlmtj1X4s/TF
KilGxh9bM5D4U0i2fNxOx/FMKEwyKT4lqez15pu/5+ImIGYWT8xUNnlFHCvYrIZS
gbBWAqaN+5ymtwYLg/2wg8U+Sew+lfiNOwJr8mona8GtRjRmFT8ol1VMAMRdytRn
6mdgero/zBTI0W9EjQ9OZVHzl3o2Ig5Bd7n3Ui+OjBL3IlIMJwdwtold81+8a8FR
y7N3SlMszOOeZ2yWRIzwh+W5v6vLzHo5HxdUV64JTSCwcI6hbKBVQwHHML4ohcWC
Lb4glLjxDmajRzNH9dMnXe44pKwRmcuDtZOkqKdsDTfbDN7syKqY+sbz3i3y7plP
+4CJcU4TYbmSyw96yF7/XLmKEYDgdBdbIbfeH3W5Nv0QizVh54bBi4+w7iU9lFed
r4hurIai2WnW0bQ0s0j6Dqtj5u/HLmrRnveBRv3VJc0v3Cwr45bg4Lw+BAJgrsJb
E1t1WNx5bJi4I6fR67U7BfoBvzCMJ+uq0l5Pb3CFSWVCXZm5TGz+CdFh0hLbPSWx
cMxoGSuChbY2CrU26ilvViWhYKI87tSBpPx0rqu7QY+nCCy7GohRu2bzZg7jAaD8
b48O/OwsGzRu5AOkXyGyv/2htUu/BD/ZR9f8oGGxDuhB4uGEh4WjnRHsFGCa4VDj
HDDLr5ChT6duPtUEVQYDIa3MwTgelOMyXjPw5RL0t5C30m7riRnPuRO74fsrjcao
RGKicIZNl3peoU1dt4JzNQpMI6UbIwre0+n0QEEDPwKw4FS04eGZlQXyGXd3f/yz
ZQs9GTM6dNvA/F/MmHFKpeOFMg3YJxuO+M7kVXaYYl+Xa8eXKXSFVMXYObi6qS4e
PZjf6mU+VojxQSMAfJzSHD8b4xIMYkCXFO2YKb8kIsG0GEiF/xQYVlIBwtkrf8cd
J3XySByWD9EaLr5+O6mkt8ZH16z+atyvpIO8kCzJGzwbkuGhdv9VhBDurSiF4Bj+
2Qqkl3VgzF1aAlp728UV2sGvqdm2d9fnXivnRNuDCWSRFyiu61vmq7DmptKN2x7M
t02OcWFzo5JmkKvMS0AQjLaEA8Fuy2lAos0uaslb4c8BI5MS9znOME5VOd4KRZZw
5F8e7cyDbrNCsOOqVqF+rSIGS03YXhMav9wHX79tQJz4gHaxArV082/Jgi05Z1qe
bq70NZ7nJ2RxDnCbHl+3z+7o4yRdmjoMv8eZf7rn35scwiDVrClReeNW33IAi1Ri
bwEboKyjfTJx3uzgCxWrOFzCNN9wJDlKG37LXSiFOL6SW4Vtx7ldqUsgPyTNGZzh
Mkrp8kzSEucLz2sQ96+x3kHafWBOlX/YJhmsd9x1epO5E/9DtxvbdBOG+0iw95Bt
4nDXkv6cK+c/f1+txo5hS5Elw/MfC3j6hhZ932h0aJDNVtBhedLFpv0I0OGH8dMv
tSOX/7F+xT5JUersbGPvI0RvVnIWhZ5yhqyOEeoVmjMty+zUuRa1y+VUv6Z6nN/d
GzzBM9CP42qed8WaG4j6C8csappprviw5IZ9mJE1elR0jG1P2JC1LejrIjIiPg95
DmDXkSARxL9DV57/pY4VjrscC1QGViVpOIlEWBQc58yk5h9iOCGG7B4ALrdmnwsY
5U8fTznqbBrW1NI6KL7iA/zAXDT9IENXyC1gwaLPCiCX8UY2lMhrTObut0rdyjtd
X7y7rZMZ+n9JNFcT9qQr5itev7hKeMCF7Q4o1eaLQCAWARev152PwJz5TdAzXe47
trg4DDrH0gwKmDOLOMCWvVrDem5j36BP4eOTsSmzE/kvXB/lmJnjRFu8XszIxOzz
lSflO1Jtzs6lHyyu7LmIZBbhC/7fwY6/Et5ysBXiyiF0PynKdOlu326ksV1L6nUC
2/uU5Gn6rXXmX/kxuT0F3Wu05phW9gujJ3oTGxudjV7BfoWi83S7xKmjlnEIDK9R
wTydwQclA0JuQTMDz5W/FtOObeGOrtR9SIYUBwjMTuO+RBH/CTE0CeHpPYWApXO9
HPMVK7rzYh351xfXMfi0S7F2mo7bKUEWaVOGiQ88zRG1kMjPinQJKhIYwE62V0xh
lv7b7IUa5xS01BVFa9LX5/TlQ36IiRWD7jGdzwbeCturl535PKKvY/f4qCa1bAyw
zNAbSiNiPcAoVF99W8fWmiU1XaZVkb7Lgz6X8Rt4zjkEQCwC3t6/DFz7ukuWMXw9
N7PZD6fhKrtnWx1spzSAMtRq0zkzHuoaZtsMfhQMGmeBCli2zFtdRSr8rLjBWbLv
UkG87xmuH1SxYj9L5sYsVVkHsYYHxINBQScV0njS+BtfmyeyFIVtXXnfCPNxzf7k
MxoWewPztrwa2AOS5C4D+S/hWAzR9NAW2YTFtg20H5gbBfMVjr54Zyec9qA+XMKm
abzgxR8H/NpLNsEYAF/30VwAKeiESFc3F+ewgrO9ImAbGIqEYGbn3oTK0I5Ki+eR
FQARxYntHaie42g5L5kE5cVGo7P9atwmsaNtO2iNroMsCYhYGbrFocgp6Fm864L3
vcj/CpSXZuXdRqUEk8Cz5hsuVcH5NG3LXbTul1JXVRTBMalBAAryhyKrZjUg7gaf
iHdMkW2+hLLT62YiYrz1nbVJ2SOyZCPP0eAa0X+enKLpr03c/vkLsHABzMY/Dx4c
X9qtU6NW7iRrBzpHgokkwPZI0LjZhOciraVnbxSoDXsYhBPFb10J6/PS8snnuAAG
/43pH5WK7PODNXZ9feSdBXk6Rv2hgr5dWZgrWSFF7zrVScOUd8M6ghk0YWOj2fHr
RH7U0a4799YbTQ/cZxKdYYvpNOlhzSjM3jD1qHoG9YcTFJ7ndS3jM6PQhRugZ3En
r+8bFIrNY7PvTND9y0GG+FCQdGIjW4wfQ1xSk+TbsIj8EznzEcEqw2IojwMupIm7
gz5IgLxzCPCUsEW1PVEit4L8V5w3wL+H5R1CD2aCwtstz0EG418jtIJrUkMyHTxU
juq+NZPcuTS4tITqWjlLJbXkHPpzR5MskJJ2/LCYL82YeX//l079Q+qGKuOZazVp
X0nmnB8SD/lq5vFnkFdbN4BfCklp85+UqBwVvqsOo9cMtKIeTO9ZvrAbtecRiFy5
wJD9x9Murv7D3bCkHX1xHJvomT6LPTohJ48S0Z0uf3VEceQBpsadVNs3fh9Wj9My
dyht0lK8vhf1dqGxTT/gbpx99MiSwA6T7ZXZZAxsrVKg6X3wo6pF0ZJ3WZ4mzNB2
L+XtXOJYKUKVPWjk5in8sA88qpLul0L5QIfUYVu/FjJgl9tqJQPy283QYnEu5Rsu
tQ968WLzlItTeyM3vkLrEj9yutewx+hH7ajFpP/QWvd5LAVsUaQjifjJR+xtw0pQ
lB38RuI0/EN5qzrw6ZHJyTEPYTLj6SoCOQTVkPpUCM12A6fdKvNaASMLH+yBr7YZ
inCC7Aa2f+sJ3P5V+n++naDRTnX3FTW+m4F1RHSpHxsSeQbBBF5N1zen4rMA/Ytd
jt7fqCRWSNdaRei15nRCDetS28GOkX99Whpf3Cq0dP3bso9nPHdvBPy+wctAmDSl
RO+fMiXPC8NM0fx/qki3fYNjGLj7jYmpgrxoGNB8bgMGFrD1TCTh3jJVzWzOOgZb
+x4hayooW//HFUIKdkXry1BkRBikydg0Ixobp+BojGTaQydg2wf9Vvb529tYhDUO
zusLdLIi2K5dXUui6rSFy9vJYh7FqmjURkcuD7YdL05GPw1euiX79gpIzLasRi2F
Fl+Lu7rhgtQflGoPVM4rxlqyLQrYPQglLn0Z03cwQVr4CU9VKPDE7/KOGh2W1gWD
p2RqTbiVGX3pgsh/0vLHVZXoB5uCmz7h5dKJxu8Sueal79DwkO4SngFvfq30z36V
i7R/f0O6jgB8pUm2T4VeHIFPYw6AFxFIRBWDcC/xZCoycbIjuVMEXYI9vuR1aFA2
AYhnAbsBrvQAQs5lzj6owqY+OOUQbJ9JPSKcvkKTOII6fx4BVL+VazRNzRkOoys+
zPEhtl586amOsp/pMgpvxwUGi2dT4+caYyih/Cjo6Eu6fXPtciphrgp+n/oI3MO4
egD7sfeNZI6YmnEqmG6cAaEOIPW4aHIvC3chWg3dCc4XLEvc74Pr+vpndnBnge94
gLxvZLqw/MrhycdKqv1WYXeaJvb0no8SYEuVqA9DFcm0l6WN9uaEcOdjmTSZ73jz
Nj2RC599dS+iEZq4XLwp8n0rheLYIBUIt9UaekXBiASVE5ltVCjBWEhSDLihqwCK
8hkL2xcQAlytNjMTX4yl9LX6DPzw7/+G4rqaTYrhHddOuU2cIgxSIr/zS3hwV2O0
y+hOHxdxHhXs22QCCCQr0lc2PycQzO1MHfxrFTeoV7QfGLhRiS5Q/sNgOL5BDNIR
+yhD/Bf/B4Xldu6GO130Yb3XzNtBjUOXrXjoX6LSmQWjUAX6vjjpdPSLQpVNPXqI
nQnki5jq2QKN7LI3py4pknsTOYJv0Br2w2reWy+gy4fYAjTqqcvzHIdBFrI0YLPL
6MSAgEZLL7jU1gvBPoiS4Fr3vHl8lZ8x01VLAXZnAO+z+0bLm2HsyywL7ehJjSRn
ju9fTJv0StpwmsAb93xTXrXavl+XzLuDR/adCb5F5JFQNk+V0O+nWi9sCk7ecT/5
T5BHmQ3aWUiCXx1hiiwbrT99S0XafNbWIfMNMzKHkCn19rgTg1H8fGqGk/u0y5JT
0mR6GJMbijD6MhBontvhKMB6LsIaGvBlBN/QGNyb2UgDh7JoH6AeltL9R+EvcGDb
0NGlcb/LZ/iM5ygVceexm7Zxi8oKzJHvHDN8Qk177XZlDltmojw5wE8+W5f85JeU
1NqR/J/uGTltPjSK34AlWmgYJMa76q0GQ9SqAyqQeJLKsNb3Mw9n2XMo78f7me7L
IiNrWyqHkbtmmrXs2C+ZaeSS6XW0kIQ8hlJ5d3XvZ5SRydZsLzFppWaiBGEW4i0W
nL3YpQ3Q8Fz6zD3bUkFxOB3JAK1/tLOoFOkSpej5aP+cadJf70Xpr/y6cKys3bRP
aK8xZgW9VtePw8AzPiF3VYCjw2EdZuMSE96BU4KD84v9HppaCosxqUDd4lJ5wLV8
x2WgiiiqQrHkX4b1RoHi4jgBjtvk8/lb4pWKDrxnLJ5hCWp89hFGyWVJI/toSRy8
+Los+JbvAYcT6qRVrGap9JPFjtDR/88BD6YEZSIY+O/ImH7KvD6rfNy3XILm7pau
NNqqKSHPg8/bxYkiNRQK+0o06UX3tNJFdc4zy7Uqxyw3UHpF7y8AkYHWwvtHQKN5
dX7ns3dAEkpGzsCrbTyKd9Y3WTtK212HDIq46tpgprrna3DKIm3Ah952bKJ9lm/e
gYUU09ViPgWvCulmFpcqPbzzcRadNoy38Zci36O/1Q72XJcepQWgqcD0ct+0dNms
UShI9z6QY3JB8p/e22/qFz+HUIJCOErz3tbg03NqX23Q6RR1/gEo27Syp9qXqlPk
PrbfETMgO1EmbvRDpwXIQ+1N4Nm4WzpLqVPiATQx1HlVSAJYQ5lkAvo84wKRKzVI
7hREL0yPkydMzrDDXx+aet3SaiS5kFOJgRxd0pG3Ikk84QIaBasD0RbdEOSCqclQ
7ArDaToi4XLlT5qg0TFXJz9JeDK1kwospTtzIdEzc3VOt8pjMzyoFXSbmLt21GN6
XVNEBVCkY6AwF+MzUI+9Ukyfgx7wC3Z/sUBqrg88nyl3yuGQ2MkJX01HtRWWa+le
2bKe1585wvtNH3RWGNPNc1Vp1GWTc55hgUEvskzdaFNEZyihRggwaSXZVw4jFBbt
LHE6UvS/00xUhGCwj7o38VfaQfwhSUkN6gwUDGZjvvAJAlROGe2kCXkHgIfyJQWi
wrfyHGLR1A42F/vQooAW8DesPXNpAvPlr7tXZ6o8w9ZuUDLEUr1N0FPGLd0MproZ
HDrvs55UDyZDVSdld6tmRBtqDaiqp9ztjBM8aZeuBrHSejsPPWdGMzrFrP4fOjYV
7qrGnzkUMrznkKFGBfl6M1/Jzd5pbsrW/5w1qGD/rMuRt2MrfBkk+XL2EHbQDygb
k9Y+ajZu8+I6kHSDTq3q4Gkp3Z+415cvgPHQmH0pjyKcXfLu+a/xnElgo/iGF/wd
4vxZYlvY2W7CTCr8w26HPbpokdVun31L5vx++KysmPuau5xVDaFXCE9mq18WSAcL
6cfcaDRMfV7mdfiRf4KUSpjLO/MK4P7fMBa7xbzMpgIaTxovrPtCG0gwUOKVHl6L
yv50UlbDFHQnQOe9VJwXIdYurQktrRg9rmlYZvJkEz0r4N5ILxnnO81r85F1ZPpp
mlRVXRbnq4zaPsswPJXlKVFHCzPiPxTpm01655WIdlguPKzE3RvhhECOLcewMKD3
hdDNF6DpMt1W7JvddHXq/yjjvH9dugDldaMBonA6LlwvJtbndhOrJGOizN7jjgL0
TtjDwoeSvJdSiqbeBKNXwUYPq77NBXckUyXZUqz8zgolkLuYB55vGC9uxXhgaK7i
UrjS03sICxLNcMdFEZx4Vkp6VJ0a7RfZBi4q6ePFneNyQxa1GWlkya72o1Fpqn76
+cffX/HpmFRnT1XzRt5kkA6SCT8/XrxyKlvDeWvqT0Kxil6UtmJnAmhd/PT7GlaH
PN/TGLgzKu0Bsx1xvnY8VcNMSYcpfW/6UAWbO/+50bo+Rp9oIIvngSfeU80TkGAW
GZuxXNm2g49Z+wwG2N7+YWiNkUjYunUtGNM8vr5w/293eIe0/4s8c3UWygecRgsL
kRUUf9mskddO/2xFiz49qE4PwK8cgiw5lxXA+el08TN1X0LfQvA5oitpp8FwJePx
bS2imfOk6r448vwqc2RW/nqNLhNgr4Sz6uHa76Vi8OHtBm8WhKuipo/y58CxyaDx
UpHMS1FZ3t8ZhpSdviepVuo5GOjuTFahVia75eTphgI=
`pragma protect end_protected
