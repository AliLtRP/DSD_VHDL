// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:42 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Szbk5OgSoW3UBsO2lt0V0iLmWfZSiaq1uNeNZWpAufLG33YEBmfHalOC8e1di/qq
VsP8Nmv1RS3YaQGb7K97UxNC9JxpFCYHjRD0wIxETiK9H4YFmNSBzUNaUXJu+qVc
XIn6K1xBcuwNjy1aIXTIvrWqBMOv39yVwUbU1Q1UDO4=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5088)
oe+aSKYrRtTE2SLkic6qXuJVvvPZ2/VMQUt26zXi2r9wvrOZeJL3PHQu5eVDYPU5
nRfRPJZKSaNWy7pUNYgVeVcbZfO0obZnITKeK/zJU/CymWwz8lpjjCbkpFcTX6FE
Z7TF3yqFQWvRpAxm+aEQ08J4Ac7lsUCAGQfvemY+yv7ATelvMLlHoVvF7+o69cm9
yUXA75Kcxp9/2dNbwNJK/7lECcu6V6cE+y9kbo7+5+ZE/V3RLo0Lg/aKdIHtQMQ3
o4FUT1CfZyPfgEFdCTXP24nhFyfEYQTJz24u72NIeY3jQfbUjrEE9IW67Psw3P3J
MS7A11AzyXnxX8sTzKLS/hnxEfUhWyKGAg4StVNTpiuPVXA2Kc621BXxzwSWUFfL
UfrAi+USJ6Ak9vz5JpWsmlB40YB2UzVffs6iPRDTt4EnR/FXdzBcwU+j45zP5cVT
elXUMOOnuLzx86WyaUxe8djhKLiAJ5V6KNQ5S/8J+6Vv1ImbikBMDdVFuUOdeIPq
eJtiZxUtywdkR7ngws9i0/Rsi9orv9xyFrUkSnxqmBnmMNWr3XhLj+SOXOl/Iouz
DDz6biqn+USM/TgtIL0n6wMAkZO3rNKMlzw+OofmmLammTQrQiN1ij2AgNCfWFJ9
D3Xe/HQc0tgGMjpgS4T9Yt0mMaXtG1FD9a0Zh5fFqK1UWZ8YSjYY0bnBiCjMPDup
AlqrPikbRf8hZrxiJa4oWckk10wIQD7JrLwSx8kd5cWdt+igmEJUlza3JIpKF/6P
FLA8UCzGQ9Zq1yWR6hwSguiw+uqaB7EWJFQ2SlDGCP++k5B/nmdegEPjgHoYkEfd
w+U9yWCoa26wObjqKIis9jtOo76tsINvYanaytY994FP3PLck1eyvwjO35r6Hpuq
pcw+GWDRYU9G8Zm/rg7XN2EEPL80tryeSQRuUJKDSkDrrq2r1en15gxVb/kGHy6z
UonEJpz1Y1fE0FWwt1T0XT8YQWbeftq8ifCpB2wgr3QzK+QHd+g7/FVL8G1Dw1ad
enmwJLOf8ksOPeUdUYKMwT44YhgFSGL5myWgrJsr/DGb+rk1XIrbkCyynlbaQz6/
d4GxCpHjPClhWfh1xbB/XOTCuTsulxsn1vttue17HheZfbTOlRQmRqSjTr2WDQyL
yPeNIP4bgL1P6DSW3wUrjQVOq4tjUE/o/LflGZcy0DQ2IKqKJNF48feOKTFee4bd
dH60jbw+i403P5gKgLe3h7sSuexB4LKVQFrmLyaxsRnm3XaQEZmSkoGmkYJoahph
z/leGXUEGlpMyv1Vh55Il6n90tAiBuBkEO1xGKqogt9eRpn8ec0Ktt+j6CLm9hsk
PK6h3Z9KYhFMAMcypiGtO0RzLZRdG8n4tOZVeBGcVJEmgxqWR2DpiOBHPIxGnS03
52ZG/xYUTjOlfuNPylBAlGShnlzzXdt1RLjJx0BXXIL0yzbOuFuux8L7s7NTFC97
uTQwNyNS9s0Qa/JXetO6GTe7UBbjTWz+HP76hqsdUl3XSKTSUIuUHBa2c1ORNOLL
k1tlz5PjRH8qoTmzABufmTS6mRPRJHfY7J9nNXRobyVxWcRinwt0ft5mE8OZKqm/
C7tx2HNQ5vMmz0BMRODvBdHmMb355JW6nqnHIGBrJZNQc2rCCuDZWuAPimq1pxZN
pIJdjH7549Ph7fCF9CdIaBA1+sFoJG2+g8lyCVOzCMg81SYTHVmzg9HzRYgsBD7j
B+znl7+Fee0jQL/3NS0Wd09/rrSX/qO6jKXHqNWfj9U2JoF79Yn7fTLsdk5HdTBa
Wy0PyG3Dn3gBZCy1oUzQUwzTZ+h6u28XfIVeE7gatQqZ2ynNZW/ds8FmY6yvB2YW
T8CRVmGg2yoEW2nxFUWwruaWIHX2ADLcuv3G5VyfnVyELQnJeZ/ZHxmIYWvl4LPT
dCMb2fAR+pXSvbUEgLeQf5R7Q2YAeHhD3NI22lhH7w1cMVd14HTPJsHDxo8T5VUm
9MD1PX9g58lO+0ud7l13qo5vJuXrw6WdHcl/d5Tvmn0qsYJLRo+5eAvIPdYPDjD3
vhYbV0JUgpsdoibH4MTf9nSAQi+B0aWbaEvwOKiPLYOk6PqMP9wvLQtKk35lT4zR
ps+Nl8HhYQL/Ut40zUtUl+vRg6PDVOsnCf34f1/FyueRww2ZM5NJG0yiNpLjxOel
UeRCTjwsMsj66f0/Dx+EL4Xoc4/GiDryQKplCgUAt4D6HAwkJFMbKJt2X7Dyd60s
RpUiUuJVXYYq0l6gqlTi94UyPSFvi3cEMgFU4ms5mSnNhrlDqzit+EE5L6fRWAI3
nTXWKIaoqQGFK3JRtse9jQnDZzE9gSHy2pm5mnSe/e7ghvflYQuF4j7oqSf1kvRm
k+3BylFjRSUM1E+YxKBz5oDICNB+iNk+rtxu7Cr4PO3/X9rxjepuuNV4gCWb/HvX
ezbkc4EfrcLFsjRDOkJTBrhvJbRKZTv8OomkTNBgxeK7B7QayMcm378m6YD+/AiL
36d7nvRKQ2kHA74yBiviZqWl5Sfc5V1OJBrEwPT+H21pYMDgxWcr7ty7RxL7s3b/
zrejOGfm+V6q5V6Z1XNGhhQGWL+GQvwGjKflKLMNCCEInojpsR8jUXy+IwRSgbfg
7Hzoq9BmFHp8toE6CXRwpMSm5G6CQitCEb88BazLBq06bVWmhfmqadJL/Z5ESgoj
xc+PhAuCBCqTIwiKsuTA1kiHNvYnux1Q9oJJu9AgRv3fBaxIuG3mCnLjJue/ASZM
C+tUOJDX3RFDREA8BCU4b+McuRrODAFSz/l2Kbx30puA5QX/WSRH5ygtsIaLLG70
9ITWqOuashM/WGXj6IDqOmXD7WF7r5Rf3U1aSpIs7asN+c2niRixsI64JEqFHmE7
OgtSPwcbAweHikzEtVIkIyYfrStQeNyFniU66hnkGfH41zuRV2Aj7fbx4N6p3BUe
mHa2jxDoo52xtBmBybxsuA2p3+IlR/Ns4oZcVw7yZOxiW2xxEpC5F1ejJPriyGlJ
Syz7Ra4CviRgcR+jiOwxLs+zpfOVbJ6NQvUu7OYvD1i0gtN/V5NuFqXZGeiL2rFL
1NTfuZKAKW/kp6YM7tPKAKeOqHnzodXV1Su/w+TuJEYoJd7Rv72/UTQJ8RrdKvH4
lXUXYHbatXB1+MdTTrT3tY+nthDqA4pEssD/x3UnrjsQYWxbWi38TIafNJZPHjgW
5es5T4z48/ByKZW9OlxDbm9XvozT7LN+bitlXFEzcRimTBYkez6F4rstvNPeLkYG
mMIjNFIzhuvESAd+UOlLYEoEr8XFNOLevKHFFCs/h+bVhiu3L4vNNA7abRHXLDjt
kb0hcDLnPyD8ZvzB4WvFqEKDZmB9PLPdlT9E4rqSWwGGEngb3MUQ7kQAuORY52wK
RGJ+nJJoy0BE1HDlTBwPN3RqOtS/RHMo5EXEvfvYMZOiMAR9Q64qlc0c+uzoSZxf
Ss0O7sXJ40WV9W6y5qOo43qQz70eJuqaI0/bjjxcGPs87QeWlxjMPGqSPKvoIsI2
FKyyAWZziPoFg5txSomHL43x+cIlDD0M8H6QhRjHbyJMg/72Dir0NvYue+HnfAfw
DwhpQBhOi8hLZ63CrOYHHHQUXUZ0kydxw4RhuBZga9JStQ6B3zpetWiB1Tagp5fF
FwowZ9r3rGz5ADypMPYIVEvkNbAhfch9AywelDAUGDOQ+/R804b3/HfJ6gRWo/qm
uzLISZxnSuGaJCWFxfAcAo9oq9WWShgSIwiMj4KH69fr/hwKJGvKaiUpsursri9F
F4PPhnJ9ywgMNBaUG6YwGJRUmp8FWmy0KtWAHBWHOZSdOck4TmcicQV27mVppPRA
pxEsFx10xW13nuh2Dr5kBRYhMlXBVmlZQW9BKyFx4w8GTHqaxPjwSXpTTym5Ekho
+0B6AeruFg6nZfk0polHxf3nOs6OAvTRXw6rAFuE0UOkchkGvmhYSveUJJ24kfJu
upExVMh1q/1z+Vo8xBBPg+W06uCNZNtj5+pgQTaYe3is0Jf5ll9LhUvWAFgPZJjK
9KCcKEPv0KH/sxaxOePl8mWygNJnZ01zNpRk+owCOwqPqcn6axO6lPUZ+my3cYL2
eH8FqEKBJUwJWiu0khqzFKERuIsp3HqX4dBzTulqzX8b09BdgRx3xsRLBNVIcdvg
/aKD8Yd/NI0W3tYDQVDEYo+XOeXkjG7N0ph+D8SLTMp33rfuceUey1dkgCWIHNWE
yjnZ9FMi4NJzh5ZM3KOo0qfy1hF/zERTvanjazGHjC+lPzOMu5VzJ6YlxFQpwE/Y
uGi7nc3VPmklmUb/2yJjtVAUUbayCHXb/n0sXIPkykHZCKVLHl+k7ZkHixRvlKCe
ZrVXdRI6TxXWD50iE3SLJDfp73/XD3IkT6mopne+XmjQsOi/pseO+SXO1adu0LNc
GyScLqqG3Z4ZYAD4T73nK78msHLJW6Pkf+VZXEteB1/NwE18FlAk3p1lCAF/TIWT
JKCsDWjtTyUAYei2D3ZYLIrzZAuJ4brmm149TfQyggQ2uSeBXOuy1wEzXk7+AbNs
62oF5UGqAXRkBeKbAn6Ucyiv3j11ZgrVR+ypCSH97JdWdCXTsfrDtaXFMFI3ZHCT
kwH/a3Wue9Yh58YjqHkeRfaU5aUBJyPnyYzAaru2CHA+pCyWKwW73MrhpfBaX/jk
8elzpMP2msIVUQG7UhtPnlIQPelDiJr5GpSwcHSik/IWBcHMK2hwLJR+Mv9T99fK
/IhoXue/DvCNBqoS6idJHUPr8XkUxKp8jGUFeJvPE9o+M5BWzHrsLj4oYw9cIm1v
oGai/h8jl5hYiITmbxnWuuhviQRhxboDuXOb5KF5xTmTVbsXFeFtrs43p1hQ9c7G
zeBQSupErYklQW01DWY8UiR2azeu/fTB6TsdxACjpyZqIq88TsBvyhegct7FhjVL
zAaRFApq6c8IRJ1EOBVbql9gTm0LwVQgNPfHvLlYV+Mwv4EeOZvNhvUFURchIZQO
8dyJEYzA7FRDOmrQdd7Yig5deKTtqjFv1p7J7PHuL2hOeWUtaPkWpSi2x/OVDCwM
uDuOITFByLV0JyFa56KrdH7FEQ79YC9IkouaRoQExqulwINdUOeht16luMCKEHhg
6EmlaCzcWuaHGQ1xxbivfvh8O4BwXKkSzfqMZKCDS/e7fRIeDa848hMcIDelLnc9
RBAj3E3fspfyDxZXprRuFvT1LFoMmXOzAW2WSGHe76xzX5Zhx0zEOlGU+qF3Kuqg
hzdgQBbYzSTK6vTDAJr6Kzk2+C1zvZAswiwJ5Hkj+QJHODmMJq+nlmgldL2GzZy5
HOe6d+tU9nOjsfKr5X4Gn/GzQoXmpCL45DpY4QOE7Z5O/axOeXfkvad+QuBT/vGw
s7NIAeiE8AXrWyzclc428GBJxgAtmfkMwSUteggs39fPJu+pqQMZadtrvht1picb
RyvUrQ4FK2dmBL5bhNZ4Ol2jDwmGTh5QHprjxugpePZZl1dEx/ABjg0mzGah0bGc
94q1+qb7P2Em3locrJ8Q9aJvwNF6NgaFqzz5NXVRVE1/uByTU7wqqEvHgLPeuWYp
zrczjtsWicYkjpFTZBcVgc99eI3jCMSdMEXAS3KrDVRTtfCfYsuqKQzYh+uztS/s
RJksT6iwRMN1/UsD6Nd2+e06HOZA9As5rXGHKKLpv4eRvHhKMfy8S3UTTuCNJwRr
+6Kkj9B8aAM58YiU4vDr+foXDXSxklw93no9IuzHzlK4jrjYHcB/NoaJGWZifvop
GZVx/im7ZBuhBhjdkK5HB1EpE2lzF5Rp6HSbt7xkIQeuR+SiEYx8hXSxFMDvtgz+
uKQOYGipoNcRgqVrC5Hi50Maj/ZY042axEYTPPMx54AYUdfWT0ulnRGI/sEwsoSL
aXIYUG78Y2B4Mh2abedagxEDTatpwyFhzZ3Zt7MmZfx2C2/D/x/8cAK2HXbEwlsX
ZfS/91KolPAimpM9/2MgI9J6Ecuu/Qb/HF+rZm6064fLuw4zSo3mCWhwj5Ffyajh
T7AjCPTEzWT6t7iQMzhoFRSPB+D9J2QtzwN3hb/onaxcIsb5zpuvyLD4gM7P+AAh
UJwXUuvi2dy8nFyvKe3ZQ2aMdq26dOdC4OjkSPdfKlNepect6hF9+MLOdjQcZzn8
Y+IbUKGzhpCiirPEN95ScuAa/W8b8+AG/w2k1IUwIqXDhdBFa8V8Bl3syNBpJMz/
rUOG0WeU5UHXyExsXoF0Xkiy6YRUi8RMJHUAKx7dRPUZ5MOoAhVkufUDhfavke2Y
PdeOlFJtAY3JMc8h5cOTGiyC0Bzy4aj73bGvbOUru4JfK23ZmBgtUk/xnY29JtVu
IgEku6vLncK02wvZDeAMe9f4CYUFQavf7y+VBslSm4nCrIsqD6ZFFHuj9bj96V2L
epv4depgG61Xk04xFaCNUtA0XcRubHbATkrr6ASrNAGbTbJnr/ju5rk2Aj4P1aE5
Xh0brvgKY35tnLy0xuTwBZmDnA/8UGvwfjunQglNFw6MrkYeVwDcHSBSQ36z8KQa
s8aM9FUKYhs/6SnKCvwTZTGeb5PueIIfHHvfTZ8ElIn4M37fQ7yviwbHwAbO8jVw
853rpHQbgdnWj7vfBLpDbBowWcfYpPgjinlkVLVOM3tvhLOIYhXjZlJcEhpctuAK
BeL+/f5aw/sBzqn3uWpyoUPRHmR2+xAoNloZC1XEbuQSFR4O4lGFjFLgwG4Cu43T
24rbQf/gwAW/IkVxpu78lTPd+b7PipjbEWwTa7MGFVgQxENQX8obqExtlaGbsITj
`pragma protect end_protected
