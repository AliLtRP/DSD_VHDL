// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
L9Yuq9LVj74B1hd7rrGmhq23qEeMRY1ub/lwQGZ1ncI/gC2Kx7q9AiO7PfbCX3dCDSttN/iPAldT
1rSDEyFL3ooeCPSywNRUaDbnyFpGgiZl5SWskinTT3oxgdMBEPLpnHWE6+OsddWmZDfhJVqJVSRk
4QqjkBYtbLd651paDmkvHE5t6Ncd0A0Fl8I/jPOyAU5wWJkTN2/sYlKbzVr0q4+xEe5apmZaJRVd
5VzUnxzkd7Aq7espSAXz7YryUi9Kc37XiyPGo3xYdI8f9sk7YCs5AxvsvGnAoLYvRHUxIZO6qRS6
8jqgHSDBQy1KJgzfa3fMj+WWK+jCSvY5vyw11g==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
JKkG03O/rzvjgb59zUkSekAmITf7WvBaqBdBK1OFgLQspcQwxvZPXFty3G76gY8RtGsJ+JnLoQY3
0qiOyBr2tD/2B+6/eaDzhY/AveJYORYgIEZ39zuLHkdd9AlxS8S1E8SbhkqBrPKPwfmwlN3U2b3c
mf+1RoY8v6nYWc9fUfFq+sZWb4Ycggx+VvZw4pc4TpYi4CPR5L1k9CdZyVPQDVq7oX9umAkk0See
TbVvnsWefhPvhwZ/97BAb8pA0u4P1EJSMAXgQhazmI/RtZd6dE5yu4VbqeeXYFfw+wKqDB5Ls4pr
zoD8/zvfponQ+IT/weCkgGL/hLSSg9+AWypn2E1o4x/LHRtRVu4gt1G2Ofi18y2NVjFCuqV8cjb1
M98VCntuWUm6awNTcur2nOHj31yNylbXXgmD1hSyAKugOh2ZgJBJ3YsS5C8tpPZvDb9RlVgSKpx/
rpKPsVH8MIghgmySM9cjLoQS4YZZFPMGXJxE4qllgYqYtVXa+wQYCIWVTEa7cVAjlfWzvlLxu12D
PvloNrz2ruxAhAPUkp++mSOeXgyfRYeQokuWX7vP7ozTtomVDDFwnreubt9Gmxs2k11YpXJokXPl
2ozgbVbpU8rkLNNAG3q3EoZPvRs2lJq/BAjoUeyjXiQydknQDvBrE53llQQUvSu0GBsIanKvVWe2
frX+A3wyi4/W95qsVR+I6KRfv5ABjOjsBfE8hATEBzgSycstDNwHu6ROhh1QSDN3SX1NHfjlOZcS
jUFMmdbUlNKLgPB9ZPKWB3vELoPhfZidrOLBo8zphMZSmRGMIyFy6LeQcMKXePim/YEFA5ggkROd
6jOUUebE2h5NeMzVNs5IccG30sFwRPro6foZIfOC6Om9lzIVbLKafaYD6w0pc8Ifkb15UBSy8toX
XzC6EpgKjeddL3xrZjZMVL0Qc1TZyNiTXAgRem5NUOpa5fbg8LniL1pcMEz4aoDFizajYxwDDY6t
cgTP+GTWD1/z+XiaRdeVVVOXSXhjT5Xgi5WYvaWZzs6uCpH5J4lR9EpQCx1QBTeQOsdUw/CQHj8I
dwGwomUj9eUV5JlJlzaE8be3Uw0CR59vPqkoPE26Ol5SEfks1GBKtcLRKvmchl02oYtyDQ+/rsh0
RkDvZV0W3063g34cKxHOZ+3vWpm50pTOOXVxS5ZoBusjsGL7UzHFwK+uwMXwhabkj/wgz2GAP2eW
q5mTPczy4U7dWfaP2m7lJpHFCYcUp6Na1ca9VHeU2y60FYNuf+IgrDo8vCSe8dcZ0neuJ4f8X94x
kdTtNQfEITpAOTzrGl8pTem4vWQs38Olrpc9IIJo6hD3CH7pJQPrUTctyAuYjECas7kquwVQP0PQ
jsYKrHH9GwWuZyFcvNv0wxmayRIEh3fKjXC+H8/HgHeKdL7wxZbxECSI5gadXy5SDJcfyjg6r4v+
R1hZy1+NEuNtgqLFhPzCRfmgdgSzNvH2JJpjBsEm84XdV6tpzBoCGnOTHBvQv3RWVJv5Cb9hC8qr
jV7de/AB4WdvgwKksbrMmu0a9DtcQhyeXEOYZcpdxF9X55n9KS1Cbhs8oZvXWI0YBqkWCr/e0AGY
H96jIPZT+QkKzSCOzkwAskAiGQBlNbJ6E4wLXfODcrdeHuEQWs0ON44+upIx7d+iblAyHHBqx/gG
QCdUrmdll3OplKzlYezslEmquzr+zsnaA6BSI23wEh3NBh9PtITShh/cCekIEbCncLJR6Ue/Hvmv
/jqdu7mgcsbpF+VZL/oXJdP1vQGwr0wDAoUHfyv58evs6W0UMSNywUHj0ZHRLZZuChu00oToqIs6
6lhRNwkihhPMxnu53QyzpYw1ZUOw94QerDrRkZXQOxNoZINNG3ovhrJ1GCncv3aAHmUROonMY9CG
7F/Sefy+gvz5c4d2Fp5mel9iYzeFuuQV4TwEWuhnzTKq7tYOtDg0JmQx6Tr5elsG+jNpfvc8J90u
BlHJdLY/Gb8VDfhCcmzRc+Xcn86jGUj6jHqhxHEi0J8PWnRF6U9CIFryzmczgSkHqN6Yru00ugH/
VeF5m0BXIF6z4es1IP+Ryjerv6GhDUhrd6mqHfjQ3qmjUcseU89WraIsJasOrPs1VNQ/rshNDlRh
uC9+qQjomoDj9rIEObY+GzwOTy5qMfPmAL3mxe4A3cGx6KFXucJqnoP+It6wZgGDHWqKNk6nqLRV
plQGlV3QPVpFFubOAPIfNf217TyReiBl0/vNSEKTErL0a2kAE00EVymWZvCi1qLNqnD5204+mj+1
51r5LHSf1nNqANmVVdtmOF7EgLxAZtqCQIpENTOXq4FUDi3NG0JjsBK5LaCiuzbereJo7SzxLOAq
bdstFF16DHlz/iLu5D1uNEcILsCMlQ5ndf0/e+ho3ZUoSJ8FtkbU9BXBSUw1ZFBW/aGNnvvPCvYG
TECrdUElTa9JcU7Ejy46ihTTM7cbxWK4ZytDAnd0f5ky0IjrMsaJCFbsGJ8ldsZmxYx3E8nAsvj+
TE0rb72PrIiTmOVbd8/aEPrYSrlSMGP8N7Bb04/jXIZnGJdxm/omhflNpjOyG3GKEoiS2YNnw43r
XEISSoDvyWaS+hC1Qo8HG3b8X3sM926QVGBozNFlzLWmkITpAmwqWQVJSuyt8+XPOS/77oBWoQhd
fotiYTlG29PYYNNPQhO2L5ZmmqwfHOpaqeNMkNLtYixyGncDURyRUZ++yBL2s2YW2SJepvFeWXzn
Cbt56OOew00GMvqYmIS40uhstFU8q5LNLTXPWxDnEj+1MmgeudHtOBabe0j2u104GB3sZblqL/oM
/VUoF7/Oy+q8vMsnYYEFaO7oXhSVrJyZCJotUaOv3+pnTHdYoYeW6XyLri4gmYc7tlSFZitX1QJ8
9RaEObRcoVyjSmruuWin6uuH17rn2jUYC85+vO6LBav/tshTc6CvzMvFIlq5t0LJFWY8DYvy6TwX
Bn6+SAIfyR25lMu3uZWW8ozucNLvoHUJhmEZ63HqjxeGfHuYeHwDEjFboxoK1q2PKh6pQ6j/S+ma
pnCJDW47WenTp8jK19hlkJmV1j9LI4a/PkFQCxsSyqFt/YFSStHCwarTmGL1WdhCegudf2a3P2CU
C88l+betCycVC7EkK1qsNHBvnE+xY9yvq5jN3oYDo415KgGrcLY2iRi7/nYSAC7xK+UFzBWwjLN/
EXYtoDNu9bGLWSgKGQqgGQLALCA7iHcht+D/jU6t5Y7Igp0ut77g4tZtOuMnBGFFbhcpHugK9FT0
tSfFch1ot/bGh0xdkIYicybuyf4Z9HQzn8J5ludR0AG8u70R3/lvu6FxinyjiAUMVVlBk5DMCK3N
/5ded3eWoaNRUDL57k1biNiGRPdgGdQhCvcVepP14U+lNj7XwdzgWystu8R46rMIRGYP/ZEjFlfC
ekZrVvpAVze1RA8sce3fzclqaQSO+ddW2PNqcBWZLE3ao7X33datD7sCKUuq/vm/irYCPhB+k5P8
zwz0F6f52/9EkOv0XeiDP8Z+3X50qK2Yg++2ui5Qk7shex7zUbm08XwVanfqrpXgZFFuxlNdZ0EY
ga47R3gm15c6faYjpnfDe4V7YO5ZWPmVC/0UBfsL2PzraCqL5z5gCl36+NtCFn6wYEsLz4v006+M
PT1mFNjU2+qB2q/w51kViZeJvkAVNBgR1ac8wOqH/9Tk1nn8hOykr5Gqv4MYX7Q9kvaAjE6BQoBF
ZAgM1komDbNlKUYFJG58uUHQN4YSpIUCjmameCe6Kc01MEgET8zalcLDY49+4tSMfaVH8HSqV1LP
gGcIMblPUJNHD14JULBOb9Pbb2VpAEcqMr3EzkM1l7jZm0mDFER34Ni5l6ofvomNJEPm5cGOncXG
P4XdXgawVXEP1uqtjLZ/nkVpBioFWb+NAqLSZhV4VOP1eCSLL301ocJ+tVQXvmDneNhCGILjz5bt
MfZ9Argt0ZQVeUiyfJDnTT9q6wCY36b9q9kgnk5HfZIToNTSKBD/AgT68e2XWiaSSiZocfd3vv+a
kM24D3QRMhoeMc0h3du3TMQaxhUBsu7DCzfmU7HRUg5PxcFhwBagn4Q1iRfVFv9/hKHYgm/aCStl
CF/fDoMWsVtgD685uBUoLT87ACnIB0Eehs8O9No1vOsSHnwV9mkcAVfzFiK4lPPcIjsN9wrTPCPP
G/+cAHAA7K9SUNJKTypgn74a3G3PatyWxNa0GiouZ2S7rdIxlaF1cBNUNTYDlWBmQxhS/51JdOZv
nAVjD+U5xkmN7lD+At6HKb7T4RIkbVUFKhFTyUdJKU7LyMwCMtIxyvQ+0bJnhjHMuaL5RMZQ8fEE
l1CtuJPpTji8gAGo3mcY8yGC5OEpUPAUrw6maK9eF9fOxGO9RYmL1RMBTQtbO9JfEKJCHHgoGMaQ
49NZkW2SGcdMNab23TeyY/ZBdFoH0wYhyz7WIHUb0Rp8LONhIzk2FRqymJ/vcxdv+4b6eWiKBhnO
bipkg49ilKFAQHqLiERVwgr4H6v77+vmYmZ6vGVS/iO+KqGr4nyEbmwwUH1V88FuiT35w0r7/UPV
SYnb0Y4UHIqQpUgxq0fE4P9kmTAgMMnL4Py5znooatUj2s97egY94LRLY0DbFmd1n4nJc9Nql91x
zdDeefIfNT1ZOCBVsp3WH/pk39QCLaDlS/EAkHY8CIcYdeqeb4oMQlOIfbznhjxiShVe/zafjnNg
ArtFZwOhHWfgI5T+BfSuAvIJ7rIpBdn0D/5jNMaAg/nHVUlGsu/sAOCsxQIf7DA/aH2pBLyUPVSE
K7CVBOyyFozSewzhPiv4mzzU3iSBFYfYOslC5VZqHOWrf+2VIlBjOr2Hethu7uKed48X193OyypG
UeBwp0tHnGAnanri60XUfT/eeNxdTP4/HNtVPrg4oTnZsmE20tXdf9gDwOXqqOArjzeJkQ7aYpXd
oL/2uQ+sDW3hqKHNRsz+j9NguYbPiTJP2Cdiwv2xSahcHZIBTU6hw7DMNUCmKfMjXSKYNdoact9h
5zq5TaWSut0ee0ScuOOua/ZoRhVEk7LTj1QoQ57ZVWlhm/TJ2WqB+AUGg3LZuN3X0Ko1s066sV9I
sjergJPxsJasdA7uj6mjiYjPbINFw72xMk8pcX34WOaozLEGZYSsTxx3KYGDuoYohpn/GPbn+5wy
jpp1ikiC44QSs5zrxKxdDa7y46FhtKASgVPTu8QHbvvdeSCTCJXfEEAl07JxX8xzagtz4RRbIInq
68tChlrCNc2bIo4svMpryZNnvUBbio6BowKHyPfnSNihJS+KD111ds7+6qu1cnxeuDX/1cCA1t1U
6WTjs20bSish/AzI/N0uRYmKcYNVfj+t1ywpo6i+LC0iok8AiSfi8oSotYuYx2ft4NVJViQDfiXF
bAMwffcDQStJ+R3toQ7WhFQbOwAyDJxTdiWqFH5JhTIxX3s3R0x7Kg7rznQJnRzsK5c1WNqVQ98S
mkWIHPpN/e21dcSyoaQaWW02kDovgneMjEoHXWCq5ldi5SB3HziYeJfSG34HeHOuiaRq730Bicsm
kA/9PGD6GsvhxkfWmpXXiXk0UbNnkGb1b0fNkW0itVsm0PTXXpGhNbprld/DeGVI1xYNpxTP0L/N
OfH81dLMXZFytZ++eQTr736R8nfKRQ4j7WogBEBnxmrlz+7eSgCb94lPpTDdRYcfghE19pP7jLxA
a3lNObQqR+VgWIOPSoxaqC1kb/64KQXrUSJyQLqSXBkIq1/lNOz2rFU5K528ngGav+KYE+HkFYEk
Q4ijwoQK95GPjzJ0WWQYn6dxjHTT8AKf12ej0fOJzmJXKvBznOrCnc5cHPXhlXAXzEHZsDwLBTQP
XXp5EUUUSlgQGYN23P2O1+q5LheZKFyo7ppUgHk/dvBNLNS3lcbqGDeXjspFTjHQj0uMW2/3uiKr
+bTTYBVkOM1wLaurKnSzekqYBsTjXMGfMzpnorzfOLtGC6vtfqIF0GA3atKiQL+/a6o3tpDXyFaC
HymuunMzvcepHkZ9otxPe82uvl7qmzpslEiw83IEsJ+FnEfrofjzDm2BnfXFCEOfHOX/YO/ngHMQ
TQiCClXPXNppildouQdzVZj5hfi7QwIzzxRpfWXnzittd4g3B3hl/1KySBdPZz9XLTyGNHn0Y/f0
kIgDEN9Gj6wsxT6VHbTHXQ1XphYPq48hv8VjJzveIGueL3RJ8/7tGsrrAgAglA5waxZuyUAiqnwS
QUwdYeDE4lj5IH9jX02vG9sofMWCug/eNvVH4gG59/ci1udxKEeUu/8l/TaNafYukVLL5EPBsHge
1GavVgpM8eWMAqsYfFj8Qi5mNg5b9K4NnQnVEfH8rez9g4zbFW4G36xvXY6DOIc3ucq5Xb9WvLBp
ew5qGDwqt+wFvXznzifoKBFktF11xt1CbZVWJs2P2zxRAnYrIC/0NyKWzMHzWf5XsIJAwSot54oG
KfxOpagcS9xZzY8noDmcCv4vPTcC1CaEbp8uolHHnEVw/N6w7NJHE66ubNGTy7etZvw/PTo+MrsB
pKUyQ2x90th43T7c5QmDeeK0PcYUVxlZMj1+xAjrOo9vpVx+m9gWso1d8njeAleJ6hWWdUaWwqWN
49mq2Y9brdPA+DCjdbYIthnB7aF3CtO+dWQLWr5bwc6a6gz+ND1HlnNdcbohQksbnkVpGmHcb1uL
UqumxuWwNcdn3AjREUjGIjMQBwoOJVn6g14kX51eWfYAzg7XCf3AQeDDwRqyG/yK8I83I/FRMGJP
qhYNUIX/K86Kl/1wIQty9KLCtTzjyCEY8P+GYjJXblQx8Luk/uwEDTbzgkRW7NmpnZxqUG4eWapO
BdQiHWp02pyJPT5DdJSS9kGbOWkSaQ2skonL55Q5CwhjCiRzdDebXpgSuMPm2uOycr7iNS023HfW
2TSdjiit3OKYXJruxTgjR6LC7PjXpPOLT+m8nucqmEfJb4f2Dep9pMqVbYugoBm97Bv53I2002T+
UMKrVsqJVpHlNijYSggYS/jHyk+0v9Mj4L4YDqma6ICZvujbPf5ZKcEwDkb/34PrJENivdQA6Uyh
LNfN1APA33I1Y2G56wUyy3vhfmfI27pT0QST9by+0A/azJpTxF46/z/wxdcIwuUZK4H10jEW7R5g
uRxKshPbmVOUi0cd+R390lJr+3boXxnoqqasY7Bx6TEoI4/ey/SvzlWo19Vdk/UW1elHoEMjmbxF
Q7X1cwFG6qUcOk8zgYznF9vPuipTjEqvODBEXfIq73Z0a4cAsRFbrZmWa4bb8lZOBPYFuox26fIN
3nWCVc8/EZvTWCRdrUEbMabZMu9DdowNCOk4U42TReH69bQBXRtY20tCeRa6p0K6SjZFh7FtIJe7
l/9sypJg1h57dc25es8o91dB8sHS0mazCoXmdsB5BZuu4aB+PocG89OHoDwhIrnHHV3rBVnUHXYE
SdJ14bTJ3VSqSS2AJLviSsbMnovuWXiPrBluzdC9MCi7xq0NhaAhN3RssZNwoDSn8t19tQH2aLTI
dtsWrgpTR/dfPOtPhG2e67cpFZ9UiWMKgG7PLjj8SnfNBaFdavZlaHRjq0GLL40D8Ly8Zx41W7m0
qXdqQA311BY0qy8AeQ1Qa8adW+X/fMkSvJdV5cvnwlAk0Z7LTOkeiiCBseEeQ/J1pifterCXlV9A
+dJVJ5iOuCZrdFgZGJDlhxWxzqtEipmQaTlga1t9vRM8reh48pYbiipccRZ1d/9B9uD4T4x0JmGj
EO/WH2kCxeCvLpzVU/jueLnaNefhpjlBu8lDHGj4RD04W1FS8mpN6bxG5mP/OhmGY7c7Iy+5E77v
lq91j5zNF7FdwyQej/23WDgjcl1I6Hg5X+KypUzxu72RwGFlWJSt+JZn+iAuVRQzYqXgFnW1qOa+
T98y+5+T7S11nNebFT56RkKUe9qi2D682RR0IGQ+3ZFjW08A4l6fRC4v/zzcIH5u9J8lljThIXLn
OwrG4kHQHGGC4R9AHDti+t/RW3B4cek0fxDYs0TCniNi0/PguKL4wr7UcKnoY/7/EPvMBRlXABDX
zSDmqiwcp8Ks6j41O89C8ufWMsmKyzCdzcj63Cues5sDpcP+XhWSbUq0IA19N9AnMefYU80958Qw
uCGm4YNUI+J0hga26+2wUdSlYWi9HGbmHoz1AuKWpIHkyP/x23QggEMEVA2IOVTcjmv/aYio9ghL
mMadS6+5A2ZrHoX91miGhHXdNGLNBzaq4D8KnT60Oe/ExVBXSxSGO/LR1I189lmgXXhsdugmsDb7
HQXsjk/kZ8eJgl07HS6Mj+69wC/Et8r32molJ9Ch6g+TQ7TfHZhZMr54V7DDILIpgVKAPIxMbEyf
Nhr6orDNhWgCXqSnbuCxTEHV3UekQJ4nor7lidEYj1nvlfNHR2BoGwjNuWRZhZqq8s/vASP0lm8f
/KBe5qGOeDa4CIXJ9GdTmph1rv/U74KNA1GTkE9bQ8iWI1H+qVUXy4RI2h9Csbu3h9uchL7c7J0X
0hpmkHDF/+3jK51c9rI7XSQNnFrCo/t9f5i+enUbPpDgTrH3j7AHpldF857qpVE4rcbWbeNKYqr3
774UYlotLa83WXuUSEo3gGZG2wVP2fOnasQJZVzbm5lIcBJieg+j7OrXQ9XDBldwpvdnMD5GRUk6
zTZL5DjQCKAW13+nAMjsAXxpN8F0upqf8DDvWGv5o5dPpChGJm6lSO2bvjHb42w01PdT+LFckZl1
1UJ2tEtFxtrK+zq7u9JOcWgph29Lapp0TFy18hAnMN9XvcH3e8NKx0w2Ktx+IksVUPWvGGutqHV+
0FjrWNbNzIumm9fpRByKWuNo/BqJpuiswm1N843O/jOib/bjastJ1ANVdzAG2bKT3HXkHYlPwoKi
RWo7TLOHKYViUwhieyhUpaFNGYVmidKHLmaw0yGZe6HfiZMM7ANwQ9wGn3hsLvUF3bu7gBXGyq4y
MJ22LQPhluMX6vw61j+TBNMzq+bmPo62CiQa+hYsmXIRwNUkD5szRGH43wQkNI3x06l9YgY2cEMD
tTfQsRqCJG7vrH03N7wFywXbnC6wGxEi6z9SBVPyRPFdfjr+aWpWJIeSAwatJJpNn4RDuQIn+tCx
PBH9Zd2SWYTBg0SCT8XV+iWe8nqgmY9BMLZu+4UNr22izTl6BGIH38avk2oKd4hWQWdtKHE5Pdel
gpVZcSLzCmLNwuOtpqHMwAE0kjOHz3YE4dp7aq0h4fYv0rXuqpDAkxSe9jsoeWImECeWLYpeul1e
GOhI/++s83N9dYbIGkVgeWBedhsLCsaRpnPbse5ia9Tnzi6EyMhh+1DDooqI/qhktTRS+cWb2s1y
HLLjeZwoaxefclQ1SxHKmbt5qTJvohzndWFSrz7RYobcm7dB+3Rh6KS5ACZZ7dEzcgCHZADr9fnH
s1YZlpOpQOeFTrVB57mXT2VijlCClBrz6DtL0ncv670mypaMAOA0BHwM8jMGWlXkjGnAGy8hafts
tPGuTS7xCJ95kt/rg9sYhYcZl4wJoqgBBJHEA0YRYXOO0DSC1NdkantjDhB3uLkgdTvcP5d1aieb
xO9EoB/cGhXNV8Rwrrd74oLe53QVEa5nQSoJ3/k3OZ/WelvBoPjH7DFRvaIz+qJTSywZPIud41fQ
Egn6F4xKDGaGeyC25kWV9CLfjZWr/zWIKllKGPIC4I/xhr09QdYYgX6sDWCkrDwOtP0Dvbbq3aKz
HRLIOFP+A+zuNHBgL49QUetijldt9TTYUEU4MvFzVl1YJ6WoDFxuAnTcj7mttThGBykse+SQ3iqt
7iZy5U16SAEOJv7FYmJ6MXReLw6kqxDz9PebhORDVdJChhrxmBzv626tjd5hUe7wP6uEoE1fm2vL
H0Gp2xybmyY8CWsQYzQyCwAWG1FmIPk/UaCVZoOhGYd4OeecxZOOWozUmGdzBmy7Ggn5Hereq+us
kTxMtW9T1HPzWz+DN+YHHwWN0Be7a9V1qelfJoNGRQIow2pnGYSmY7xbzF2fP2EpcDXEcUl2G8K2
Hf4CRLu+Ap1fjbPL78H+u7jFFN0aXxnPG8WA4R7hrtCnRugan6+xTo9SRkKwCahKPlWqHZc2oOpj
2+vrujZqa2pFUWOq+EREZR2r8ecaRjL1zWZ3ozR45L3RGYIc0Q2x1QXgbsJaT8YmRls9PnzXNo0z
xL2BPZleC2K0X8gwNaai9I7I1fQ/KjpKNoVBOx/Sgu2w2pVPWPyH0u3Cw45kk48jlzdQ1LXgCYt4
ODTQxodqJXFcPp49dKW6wWRh5c4SkImX19NS7Ji0uo/GUfjCnauSJfvQqPQop7MxcxougndoxUX0
HsP+DQynE5WZBIO+a28ELDYUpCLis1TIzJLjNN80+ybFcBK7bUmtN5rvcuCZK6ZCD3sE6t0/SDhN
8IWQEfa9/5RhXzuYi1Htx6YIqS5Ciekxp1IAHkPtfB8lBBoDLdqoGZLK0aZtW/9QzjdC5H6ael8L
6QN8FpIBr+2hJcmF38Kq8txl8J8NDb3D3UN1hteywUHRx7UiaFI2JEbES+y0KRlbf6pxiZkAQzkS
RqyrKQfaJ0Kis3BM1KaP4SF/EHHJ1LXMRhkfB5HfTH3LVNLrpT+S2rfB0tSzM5XZM722XpURbTJq
ab2++tpnNBdOuG/ffMd5nX8mk9KenSRyck4Qj4sej64dVAXp7SyODgJkZyDs0T7qxP/MApFvB7lA
Kp7YweRMk7WyvxUG2uf7UHBrwml4q5tvZhjImPdi1mNNyJdDtHLvVCo+I7XLiAwZc+r39n4s/SQV
tc+dlHdMPZvLhCaxGIIPch8sz3CKbFOkqBnvg8N5iK0QTSOUG6iW+UrD+fnj6nrfDMvgHiqkg+x9
zo4r803WZnQnJTy0Po7q8i3XhrtME7H3zeVtgW8aZ9P+ZtjMbsow6kyfcnWuRqdFcinuOLbaJ588
H6VF0X7+RiGB+DW+qoUHdHBGOnzFOTRYmhYJJnV/XVWtM4QI0+D8HRiup9ONPTgMAXlqsseD3iD5
5JEod3VgpZufRYpN5sId7nNlGnwffLIlkjN6U/Cr67Zl4RPtw2ye8EncJ1Lx93pqIyoyG+9NZqyf
qL9rjSwzMvHBdf1spbQK1/hQ/WekRRu4aad9Pe1SjkLdg+corDH/42cW4yNUJb4iqyvricqtziuu
q6rZ+TfiyMgKhN8ugmxCf0TDX52IS+OUM+PVzKM/t9l4KU38BH+WvHiVFlkCoab0uYHe0KJNUZMl
GvmjJ0soLtkHWs4AKXql7yVBV4cSW1P7u5K2jIMSacIiAAZ/PuhYDoBRFhjK1m69+ggZFR7TAP94
1msG1o01krtqyJNXD20gqZ4CjMYH1hV4gu0wUZ+p2RxxDgwbCff6fbuwGRQ5BWo40dah1yZ6pAlR
cCelv7SNDjqxvNg8lVuCgG2VkMnkqFEkY8c4AUkm3YzElrba63nAKA3m46tcK2JLC/KYrN3lo0fX
xMovXx9I24gtR0dx4ov9cyIQ7vbSeWWYGmjmR5vug31k+YjwkD56b65+gJkDX1QeK2+u4utZbKDr
IWjZQibvxcsutOWrVlkkaT8Ij07A0KAZujQdGaYJm43BWin5u6Y2AhFAuLzHejBM1zi/oFX3zZyO
GRrpHn4ORfZjbaUqvNPdRHx73TP0wqzSndugxeruqm1Q2k+I+Q6MlTUO3ut4YLknc6um4FhwX2IZ
etYksZ6Bq8y23zFNXhHJNyIfVGdnwDi3kcyV3gH3bpdzQihD0N4xXcwvQ0U8cJQGomofQsEwosO/
n04q9aoOrOWfjgyg1q2td16oVXOI4Y1CvSN0V/7p39SQqpzs4FqNQGvX4Cvi6CGkB7JeqhIDXF4l
Y/4oMZTuYjYItJzeM3cxbjOZiM+xXJGzTtTIg9Q3yz5VK9TPI1HT9J1dLdZ4TlleNqwIF00r9E4F
fjYZ79YMzg+qQy+XT1PYxIem7Otl/edFRkvj+zsqzdSd54Mdd5BMdOKcpbOvJnNk7DpQpoVxi7at
+9dRCTwDxGAov/HhmLMIlm2QO5Rg2I4U+8DqUKPsAlhUAfAEMS4yGrZ3y2E7MQUptuxtnYG60Xy8
952/jXW+guIoQ6cu1FBNpdSwHb9IJa5GBibABZZSO6HsqhfAUE2CB8RupPOchuRtMYo9HOFp7d12
ICF5BPEVZjTV6seyOpfV2vq5kJR8P4bgYJedvuBtM35MCuxEpF44ntJIC1lYXFhpjfGh2y06Xzka
w4+fSfiGxoWTABw3bI7DSz1ZgitTJHXZpQ3v3JTvUxwiJ3s8QvbS1Cf8bLUamvUy5GI0w0dLuups
BN3KiqExXA8Zxdxn5G4ZdfP5GOFbJCzOTrK9JgFI5puFRBjD+WFL5OCMOPKhWKbRrYI+cuJAp1yd
ygZ5tqIZ6UQfahDCJCB4TDeLfhF5HhJHQ1xrE1/3RH9m9PHHIYt2wYrnczrF6aE/GJWCL3PPYu5U
wvwNyRHSZAjJxo5Jbz3FySTQ0A1dlFIZBaEKaIz6d9wxLfFvxxVxP/NWYVXLJ2NAvsXvHnBza7st
eaaoaecwZHyyeIrMECJQLdQXYb+FkYzjyDZzjDHNihIrrx3ZUxQ7tMREOliqeH24wVUEzvL5AZ4H
qwPZHGLLEzkFKn23UYXsZN+pO84NdHN+MdPIBCPo3RedoCosfGeTJ+Vn+hX0ZVO0Neg58DXfRuIt
i84BD4GxuOHgfqUEEeCvOudWss/1OETcEfrqD9dxzPrM3CY5CN4n/99Y8WDxBBlYyBXjOhXDZCH2
jtl1QJkYpwVRG9Dt40WDzAu1qoZU+Z+js32KcMfTEQeIsJunmLkVeHpgv2mQLrO7WaFbjKTblWYS
ffyAoY4vIApKu8FJVdDT2Q6C7MPTvCClmaP7Vp9tmP6Xb0iU3QY0FTeCnFPyS4fUGM6CpW0GLGgD
mVaWiCDvrVTWpYddZWZnzyCdfdU6kWJqCq8p9D5FYbZ0cQFwIDh6y1F+Aq3vopd0nUaCXs47WV7Y
W5ZfRMjIb5JBIE3Mhh3gQK9E3XMe+Vvb64QbOfwmZDv4LqARkhhgpchMsv0cPIQiMiMjcJS7CXEh
IvP95wCOIIWmups0OGUTy0k3kLjiK19VqtQ+H8td1yn3bctyQ6rwqMJfvzkMyC7Sr34Eb0h9aXaR
ylv+Ytw0/heYLMNUGp49zW3DJZKTz/TWRnRYxOIZGq6j2rMU3iXOj3mn+nMeKlT+vYQjlu+FDpel
QxH2hnLUggB9l2YLP8BmGryx4y3yp8zTk+EGmSxHbs8i0e9BX9tXkyHcggZRZsbhjFEeodqDOKI1
Y8wSfzd2gW8vFWf8boEQxlfKbYz8VfVdguh4dQrzaPwaYB9/fqNarA7lBJNdtWSe6QSGt8ZTO4Sx
u6CUFB7zDJl4j+nDjxTM9JXzUtBPlB8+KNwDAr6en+3UB0XzW7dOIrCgFuzmQpZsANrHF3dYEP6N
UNdEfHl1NjwMKqSUBoU58cB4fCVuOv2nXCwLc/SxIJtOEwuw9gOq0Fm095C0/mXJ04NdX1K9NkTT
+naO7pu3NmWlGY8FvLDPG67eN/a8H/JjAtydVf9Fs/+2YWEcS53FWo+lc9cPQI81nLrQ5V+kmFeD
DWKsOZ+zNzGoVyNnhLaQTDmxfTj5diwakBoTawOYjEDj+/5Tosu4/OHgNC7rbXofHSucrV/MuFn+
ySQdBwKvMLnFo5f5K2atc18MhC/zPeSDtwuMxtSCTlZtY9Ftds3WcZBkbjIkeRU8Xw6fY6KRH/Cv
8ZIqzrgO3pNWL7NTsyVafXY+llKBVA7XwrX9laKT3y1MmHKmBnrGujGto2ra9/YckCVkSlAt3zxk
dhXdiqOi76FTBoXCic9vlJCXYfD8ZY+L0ScQhnJTLI5qsBcvRCO+RJDNs0ypVO0nzi3wu8OXwa82
2ZDd9m9NDGtpwrJOVoacS7VIsbq5LPahOC51F6VyTdOQobYa9DqYi/X205PN0fm5misTyLsjap08
uzHiJ5vz0v/3p2c25hKxRvSSIDrbHHTOhTN8jTZdf8jaiVAMLFy3H8RF7dIpXJAxCqfwlVvC8ug3
tKMi5ioL7FeJH0vR900mnazEGJ8rLy/XA+Vk92Xxe6ChjqdwAZcTITUBzNl1VVw1UEFTYTLcS8Lj
3aaIG8N2vTw1W/H2QRMgxZ7l8BSn88TY5GV394lHqdr7zGH7sZTFCHa7CV6/O3+h0BI2FUgvhDfs
fym27aUt1tGXAJIESLAU88el3bj9cRUFjjUBWsOrHj+4aOtGWzheJWoTf3/k9GctsuwCKsWMad7K
SC+y+d8oVKZtqESEEfO2Whs1CA4DDAVmmApGwk3aMwyUwL32C4XfYC2ajYF/E6jlq+HkA2mZz0jT
ZKPFkFnqf10GSpz66HSD3Pn98sF8xYc7G6bIza0GAHR8+m+KrVJb7qjvleP7hklZPEiuYr05fViY
7fO3T6eqSho8pKQseq9X7K8QJ4RjeCXdkEIu1dr5OGYQNWqZop55/e00RsPiRCZjJ1tUfGI9/uLv
Nz44k8jql+PSUaZjKZT4S7lYHR7AoH5JR8auBSH9yNvRxcwrmDR0iFYm2MzcSob61EHEAtjC2g8F
hZDDodB2HRSI6esgQRF4BuvDqL0fNA08HoDNItcYd32myrkvHqgr18Q5OK5SNCM9Omh73KuXaIRV
B6o6MwecwtTicVrbeUZHzOWh3N7jTHLW19EfaJfReJxHrDP6osJrq2Cl4NBEs4URnGrfsCybvbiq
EY7mVRUzHn4udNPXTodpjnRcdKYhOXOo7of+a0S8GBkMiLx7q5Nth7PUZC7VvT8wSMvZa2pvT99N
kbpbBrwQUdJ1wN0ubGwiB7De1mLrDffn7eFnv6GWmox9SwQpolknLwjD0j46ta1z6NAH4oR10FHU
+OoH8F0UNpm732nw9R+axijHF8LgDTuHhZv+2udg1f0nfCg80av2TUHBatlbFODLz3BUU10j3kVB
79+kp5NO0FpqFe4yxVFX5Qv04Xo9XPhNk5V11n5YzhXRl7NjsPdtCr0oWAFT2oqK36yj4tZOaat6
X6tsye2rhbWEwaMOadocXomhl04Jilw00C9KPRTvos/jO7FhueNYdZZuPEepZEGGW0KLiKaEUl+W
eCfg79ywq3WFxp34KoIO+T7rD1nFHAAHT+clfvrC6ACUyhK7C/v7rZy94PQAmf99j0KeRLUpEAMk
tWfSR8KGYKuU/v4cAwXIbw3bt2XHJoMn7OSHfTdAXX7cVlElvJqqG6TPaqt83VDhoFguaGoNNixs
9dMfLSVQV7dY7bT9q20x/on+Qw8MKz6+UwfLLbe4lj61jMg43eqNHN23fUR7wXS6QnsZoGeu90EJ
PouCqYrZlcaqOxoEdSENOZ9nz1EWF8R864ebiHLdV069fk9prog6kWKf2jd5GHLBmWgh7+6XS+CM
x1fduSId7HV5h9AmXh34VUEL/SD5tk9vMXzhIFRvforDwxrB9IOX1Y9yVSKXXappp0UFMI302ACZ
J6mBvKzCfI8mczQ9sRLJZr9puYdx5RSorN+/OFbVVXTU0LDwJTjbbSe2OZHmcNSj+yvzDyHoC/Km
mahtUzPI7POMkS2Z68P3fWdqkFUO1wZOI1//kh66SbvcVUvgNvEcXYJBQMxWzOmNGvp5EuSSnC/S
0PeLSUBA9vsyz4y6Q+si0l2LSmjAc4wzrXB3+mwmlpGiK/2pVXUf7lH13ICO2yo0kWYmGirl/juj
G1f+/quQW7b+S/TQxi7GOdn9bH0UG18vnH1T5OkBeMrmxraT7925DpfxfKZFqgu8iQwDZ78bX8so
eQ7FVedJojqLHULxkLn+oHY/JQ0FpkecO4587fWvZda+FnSH8bLYrZA5NVjj4lolWjrXqOANuukH
r22er1HL4ql1Np3BynwmrC5UH5x0kd8HlvA+9mp0rUY7T5nXN5hEQRxKhLxTcYQScBkbRtDKz2sG
WZagSnhm+s4OXRJAmuQIuCpY9dEZ8VH6qEcnTIzvKlZ5bWzJx+Hz7VwFg0ho4c6ASgzDwEgVlRdM
Km7bDArqaIEZ5TM31nIYaON2vgAW7NZaQ84I7g21Zzl+oDX/DVDaKkofCR/5seMIwGkoC/NrR2Zg
bsW0CJpwWpnkPdiyoicd1psFM4avSfn/efj9IQaT7iQZi8rPYUi1DYDOA2UMiYAiiy3BEzzagKDx
Dk730q6jQ4auFjkHtVDEalRvIGdXpnrKkxYmQPiHwj+HvLHdGjjYHub0GNBGq4IU8HLfIpSDWeu8
SwcQqsYHyp+ArAtcQdPZDMqIJMMEggoBc2F/er9v5P8SO3Ie6UUxzXD2L8argIdsWk3wcjOtVjqW
9uhulC+SlMzsOvCNiiWVQxU8T4ksKEBhu2Hj/PUXBZ3rDoe67GXBX1aFMMlY73uSVKwBQZTMhP0W
AirGJ1sZcEcH7Uu9lZHqeo6XIPVhp8AvlaIJyKrtMfDVM9Yrrfo5aEtZdtN5VXDXjV/xSQz3zurR
MyqTcy/OLSSH60kFM1OnKdDOxWckxKS4QpqF/kUupSS4P4Ia6pbVzZE9+j5NHRVlWEIgIFEXYzts
GTm1i/YG0bdUIwPjCk0ZVV1AEFpIT+5Kul8kQPw59FP4bnzcbGz+JVJE4+emF1EnHTWB8G8odE0S
JBeS691pQHAAkA0YLA026Y9vxyJGHLR4Pl8UVDAOTtlWU+JMYUEql4uUdF11vTCL3SLOV5B1s3wO
RBaWlQzt0prTN4DNa+xdkU54fcNYzMP4CW6Yh/NZUUFyZcBwMI1a0uKAXcwPu2qg1LQq8DmFzeCA
XkqP5aq9HbaydoCjcE8vNmKnYuan55vdER4U0ojyA9WGsTJCSwdU698zVU88OM8ZR/f7h69RL55+
sXw0CvN6nd66mDfvEoPqTWDOc9pXoq305dicFnhD2mFW+VFURwj4XYV0z2qwoU/xy9dSJnK7wioD
S5UHMa2ltb9vlHyTCXLbvmE1TkETBAJeNdEX7jBmtDKXUfqxWZnKGG8zHxmyqBWvS7G+aefQGeiG
ejAke6PZO1+I+TbTMGIiYwFwZKStkfc1Hi5R01vS7gDomP4rs9NfMC6KtzYJaQ1W5h/HV8fCaxtC
m2JkItozXaZJYfSZhqGMduNkx7//71N09dgK/Alnc5jePNspidLo4BLFNawPU58JAfTnKkYPybDK
e/7T2RiLLpsTrPepvwwoIYIBjnonzA2h4UDN1ZOa5fqOl4NXyaQBkEVzxjHdjGEgOTLjbeLjbBpd
ERPKm//OUXkN8m2hScohPd/upRKX0s3nap8uwyQCIbg85QdRKKazRWkKGoA+rg3XelTZGeJCcW2s
kwvL2x55hhGZ8L6nQNhOeqnKHPtRtH7g2yUjlJYJsLl99CZgGMMeFe6MKW844cn10aRoYDl5I/K4
xwCucLDpUuyBaYSIHhdzAelPSSOspr5ThB76z9hOvP+OUq6KOyeZOmhQCInfUBCFFI1hb1L6kpLX
0fv05DieKbZ4IY8FVMJdydVyxrTXtWkm+eOzgoMmAKGylKqrhEsEwucj+2QXn0aKIKU33XJ9bB1F
Po5R7XeqJxoYwBV+va9Jcs41NE6vW8ygq6Yyya5tkQ8vY0yIF8YJxymhqxxvsAg3MgOmspIYpsAS
ER5Fd8wULxDax0LTZFzaZ5E6NqTEzSPgzW6axzOH2IDl2ozTblPgZCsyYIvd42Gz2z27jAaSt5sI
ZjnNnpIfz0PNMFq5VUzYDCpk2nUyxoQS7kcxdFkfTqY9I0htAgqbFhVwYEoVxjCn97Z70h8zYyef
VtiqMvjSlITytUodtpHj+jNaaPPbycX9sylsvmfSA0VWfXVtiguaLdY7kSL0cZdSUud3IXT32uJK
q2R8jiIbtJWd9ZQsQrLGxiWGT2yUg11Cm2G3aRtOHnLKjed4YEMes5mWW/IQ7znwXzFDtkkDLI5c
wbcamcWa6O8Csx9WAlw+5mgw53xqPWYwUvZEie0ElCQs/EgwednJb6amOKuD1yIryNtX1VAtawe7
8VqydXnZkakPaYi95N6Xxvs8wuLKIdykdoxrEfQqYuUYgxIm5uzM5qKKWBOUUknfU9pYoK+/xRn8
+eXWveEAvvGu+/h5g6zI76xAnXRflSv8D+jA1bIbZM3nmFI7XAAOAIz9Wt9GvFRPHQzyM5m0cfqz
vdqV3MzIkFATehFMZ70TvPfhWZH9b1KoORCrgf6ECo3Ae1Hs/lSZe7lH/fgU19HpST36ayjRBxXk
Q01emf6PmLEDrS6a7noqA3dnZuGKjlAXMbk3pprxG5+FQw9W+VW+9Pl+WgqfNA6OVEPMEFDjCOGI
EErylAzPdnAArvjq1uA++ZqN3j14rrAPBM7gMtrVBT3ETrlZFaECswmyWogAQNDcr1YfMHT3XBxP
KJubUyTFKbB0v4UYAqluuPtv36bFCPeFEYrlyXz9l8Y0jvPkT95NLUCext5yP9DTcuqdJZYhPFIg
m3VDsxgVHZUTj7t/An3u/wA2hw1E5GOV648fvwKoSLf7e5+oWL7EKSDBrEnb4Nkl963cDEbGIoZQ
PbCCzKb5xoq0l1ZGzOjctysTgaVauXaEDRNVNU5Ki/iNbF8njOeudENU2+/kpVD1KHvz91wMH3qq
A2fXx6mPKdK8noQawtyzqmouAGrmlMq5WBdlnmFYaXcFCvDfbP51b8O0cnkJYGpwVzoNWk8WsuFF
94ymy+ClMMQl6V1JwIvck43Oty+HpPClx8UvFz6NyvAcL6wizootvSweLhfAncQNaxQ2NJuQLWl7
xXwiPu3yyl5FWZdrgfuaf8CzIVZ/6CM2y3d0XIaXL5AM/rkCT3Jv6I+3x4hn/EiVIKUYkmO+Vhpw
jEiT1FFxJUETBmLNhHnia8VJEbnuvHWoMoBra7r/HVkd7IEG+GPeLE4nsaGhjITZ8+u1vVjWyq8O
ncaf13QRnSGaRw2nuaVZfYS8yNqbw1pyEW8MH/ErlbiID6MID1MUy3DAuHZYQDM9/HHVN4DyMTQL
FvGeFZfaqcP7Z09dfVtzV/sOYuKZRk7C/afYZY8DBSRcKhi00oKimDVeDRLB4HEnHbKZak+LuNa3
uRujimyg+FamPmkTicuO3nMQ7uH79JI1wJrmIFLgJrLzORN62OOK1OUpGANfyvFEgLdHFC08cYw2
7vabbQEvpuYjZfWjN2/aGwBAbLQ5ZCCHlw4IyUrdfbf0TMgsF/2mVf0C2lp5zAAI6PfFGQ5MYVsj
sd5eqIMIETdIQMJ/7DhBuXR1cin4Gap5RZsJPAMZ2P3Lu2gURYUFZWBnu2ap+4Qrtnq1xWf7d9kb
k4l14wJlKsMPk2PFUHaS2hLqGFEii6yc8MOPwhjf9EIgj6I07/2C3YXzdTSybytrt3PeXn9aDKPi
j7xjAq6iB0sTsxop0QExVVmWTwmZ6PSBoF6RCXi80RN9/vtH/BXvipdeCENqR7gMGTRnA0jI+Idg
BNw1w0bEggjxRXFBRXMxuHqgwLfvQ7KdbuGGiOqQxxAKnSQqiBekyqblEdPOyGCAoynkK3oOwCcC
gEumf+Jdw8GYorjigjHrX02wzETXI8L71h5m6aR11DrEj0Ux0Sgu3XdybtOlePpta6qnLMNqpoBv
OqieHSlMasjIPaGyA+7goRds0LraTku9K1+WjYbB5LmNtjv0I1w/ybk1YxIU0fcrjW2vFXxXoRdc
81Korge3I8lA94Sy4z2OBGcShuaWlaBrfz0GIOMUboqD2yr9TULSSFIPQB9YOXqB9f4SsfSQuXaj
zbAtsQWj+3eGUqfN+47KNBpCoaAiAYFNBgvujG9EgKbnJ7gzpEtopGXa3o97RGkkq0bPDeLHSmwI
vDttc4bGsgcfAyKjMLFJy/vqwWzvo5267T41dzlqqGHbe6exxTVM+yS1Qgxup4hzIbJWhmb/avHJ
w+er31N0wLeNGNX1KVnsmx1tPM1bPOeHAGLR0L5sxkelpta9DtjGvj5HvEF4oKp8CWXsHPV6Xbba
9tTAMhVmHvptxM2wKI0Os3eYVJG7N+QG0vjp4jPQ7MnOT2K4Q/9sQ2F01jVrWk1cjCeZlvhJjW1K
VLEFQ7rNU5SgExqqSYMPwWM5dpPKlOIV5LB7zQ8H6zE1KsEWiJbWF3PlhxCJUvpb5r4fF84wQRYj
d+Ek6jx5X4yBpWt5h57msSt74N4J0hev93TwwVfqdhSrDfi7FjjrlVC3+wETvMQgAOPC1/6BNEMB
OHhki8yFwON4M74dnqLFweaTTmSQEiac0XWglrZJN3fvQFSLkdlHFEWsIbFhuyPkhaUxFl9db3v6
P5fGjMc5tzM7Y8z8AVE7JOjqaQ+tYI8g5Noyro+duOvXzWidiYYHQIPjRq8q8bmHBbXzFFZhZZUV
I62fs7R1Q6n3Wx76KoAbcbWDLvcv9ISwHLMGBiy04afgu9TFSq3YFng7VOnWnpGnUbYFy1Q8ajUP
oJMIp73xrkFfJURy5sViIRs8bzlz9HcwMqFZx/UwKOpRdvAwDT+b7gu7aXGIro5kEkfciUzXo4v+
RVddw3tD7tGoZ0vY++qBx7fS7LREdPQmpGFjmKDsiQ16z5oTHh4ukcP5VtHthYKkfD4s52gs1Vws
fUZBiKi8GSy7nGpwbDZbfrx/ONzewcpVdg3GKihDmmSxGX4FD8oiIDvzzdbACG4RKQIQPQD1wK52
yh/UfqlbPxrnheA7DSvGlFjBmSWcyxJziPt+YJV8OSGHlw5Pg8RTsMYAcgmn2ZX6aM5JGHkSrc9/
l9fXTxcDjdTueVL9VMeDHi8EhgHo9Hwx6GNSyAFnYZzLgKucP9MsiD7+Qzp5LSYtpuKZbg9s9Zz2
3OUQ4nHaSNyo/sriNmrt8YloduNLJwtA17qsT+Xz4vKhE+k/c8WVIqz2eudZZLxiqk8woZ3vgpmo
9u66wdfvGYlDV0RtEgHLZUfpyWCGIIWWUUNvxSZR/LXiC+a0jGxudTaupBKcrsiQYJyP2nijbj+9
KdmMS9dDybr0zIN/6bSC8nPJlVzozU1g0hjutZiLvHvzG/IgJflti/44Mcc1b6A93LrnDFUfjpAn
zp/aCayYumIW1rexhrNNa49i807rXdilsEzSBjxIdNjuTDEhf2nGCWsg91BgiOi4nRgwHGZbHHuJ
Fu9Xu5R9JclPYgL1mEkIme2GbM+76pBPbzjxgpJjFJwiJCEl2YPwjgUIqqgiL+AjPzyNBqUwR/QI
RJAqBMr7Ux1TWqhIZr0xId3pkK85vIVl9fn2HabQrT0SCHXJbjVPoUK1dVTVd2igxmiaj7B3okdJ
aa8EW5DZajLxJa8rSTvB41yltL35VTe0TRl7Q5WnZt8mSduoo0tQddh+5Kd2I6HiNkUZALoED+Ek
lp4MoKgO0Ttzi3wYSycZN4QFk30EWCIWeyp2ncqjDydY92FDA4sIu7oNb/opr+kPAQA4azMSqEmv
yJdz5/a5z9JuQLlSP/4jO1o3gk2V4StZNNRR4UyqqkgEUAZaUCMV70EzwL2AoUTueGjznh65Q0mH
EAHLagHlbVOrjtygUrPkg5+UZUPIOrg1UuWe3jEminsSnbA3h9R5lyUkMUQ5fOioTY/wI+qz0Iv3
3/AqxiNlumaOboji2yM7J8+XPziD383b8v668hW26j6WRGi3uSYJY5XDqhfEyOiW1UWIhfnXAGqY
UvyYIlUaxeMY1q5iMKQME5ReRl0U52IhLY9ncMbfyIZ0EC7yKDkteHKTTBA8uFWbAHrxOo0r/49U
qkbfsnCr5Sdo1qWfB55wyW2vQZPiPDXbi5Q/jN1KbXsFv5q8rFxnYYeLwhLxakwWLOe/lqcuPFk6
RgzvsBRdEmnCxs7KhdJeARxCSbFpmwXUwbBxW14yLSJv3fssmGdcl64Q2fIrKb+HxAHx6R6TxKb7
6CQmLEn20ANFR2qSp/nL5pUExzJwvydAVpXzeNqkPjuvYs9K7ddmdC8jOL1aGCC/otuobfZlaZTw
tpt1JhIdBw5m3OQoCrEa5CEjPcKGsICMkWdsH1Mk8uBActHDFic4hHDXddtWpWPpqPWZW3GEp3mL
FKIbM6pYEHjA0yQaHwZDh8IXM2XMtp69O6ahrW3Ut0yfF8YqejVckQgfDq7QuNJ6RqI8zMPiKTCk
to+22ECDPb0gcjR7JsXNMKL2JELNOkMliuI6+R6Rhjf0vBNw3CkFpqvbag5ON6TaS/ldIdHRLBAQ
ElAeJwh5toP0FqnjnWumzQI7Sfm08or6IWb05ULiLa8Qhxy8hrToJW1UIlcz+NT3ur50jX+WCrcU
R5q8mSiOZqKEsbAPyYlVmNa4Q6SsvsTZ+CrWiSEhQ65G0a293Loo3WzM9D5oJxnHeYpU+tKDp3lI
u7oMhv//ZX8UCEvEL90aRSWpziCjLj5Ccrb0PaO9ePe2icIMys5sLdZmq15XYgtBg7PSPzpYVRrV
Z1Fg7Cu3HV7Q47mPY3qb4htnOvFdx2sJAlVQ8I6/+birqMUWCyLigPhS4F04NJmX8v0HpNXwK6Kg
xdVyCCrOQAkxn7/zwKoPfLR1KjJIdwQyQ5tlMIQoWNur5m1P1Ul9FD9aR5ixgaQ8bLutypagltCD
5wb3cTVykIkplLCLp59JdMtEIhLSijbd5PJatQJBXGLnss9DI1mf4C2UjtYjD04a4zrtGAMiovjL
66JHBzYKy1RANP1QPaNm5DJLFr6u398Nr+lbCT+R7VOeVaV/rVCVkK/V5Jw+fYQvWpF/pR9BqfKA
+oDOEDwvMGCP80KBoq5GT8icQqnxobDdnypul5ZTsj65IUrQJcd8n4SIWiYXWTs+6xfRQ0Rcf15D
wkFI+idvdZmMc8K3CAXDrZDdalwP7dVb6tyISDOo8uq7/jO6ZNgpEAv9IuGwqDXnh/i9dcKbWRJl
slqe1lFJkJe1mfEOTC/fsb8m3dbP9+eWm/mSbOW/0gqYTXTkQxTAlSh8GrXJ3qAKQfrxQPKWZ/Wx
fbL1FXFSt+Z16ZibvUpizGc58DErzCfku4vXsmVQW4nI04r+U/nhuImYvjuyGazQ1zpfLWGURjRo
KTcvDMsEPuS6ioBiiiT/O9J0hUu0QD2SGDhUPHPh6E/U+IcBPxxLN6mVmDLF+sU4p1ARdUcwTn28
Zeo5vcevmDDimolbYX2MWnnSKKsWKiWnt4WvVuJkggtHOBpONxKYvgxrw0aQlh7N8uXZCDAU079q
OE+YfKcOtVqmCnYH+vLm2pj4VRkCnDCk3ij7XtncZTO2XOL9hNz8iZOGMZuu6RuAqpvvm0/kLnSM
gT736nvWOs6hq8r/UGZWYYPauLvqNl/gt0AGbk8xZi4NDVAELlxkufZNLosBYaMS5kDM06cxUGez
UNIweJvLtrYSBNwsCGeAJ7YYGElQRsYAJzjxEv/7ZWmKYHgd3RORYTNCC/V8qYK2T37dlSQlFe0X
kM7sjWLoAJhD2zjCRV7ulnjXZ6pCqpX2QnrOExdS3VcyV+BFT6BgdpqudnL9iC7gJf2i54e5aHIE
n3/68yJ9lsvAfL5AMB/ZF9vYKSMCdgolj7ci82KIK6yNvzb0oLq/ZfIpc0oulM3JvTTXCuGJI6Zj
W+Jm6P5XbJcJmMbDMU9yEasyUp/12JIdldvSkyt8EkjNsXhVBYauvAYFcZ2Y7lXDqIIqTSv7Y5ws
7BOSzRm1Rw+iCA7tvQ6UIkSurGZZIASRacJ5JyqnEBsqbALVj4eq0PCxG4uWTLb2cIKYm5QWnUv1
U4kUIHPkh4R3VTWBLVgijO3izWtUPE+4BlcD3/uiBZWYS44YfXZF4RLXQfDaHhPHUR5YUjtrKCvB
Ya2EElZDTe+JY1AazU7UUXdu5L/wE0r38JuCCj0mUw9TlPHq15jmoegRzgAqfmbdisg6Qyyv0FSc
M1USlAv1VYHy2n6kMdrDR11eg+990f6LMyiFUMCm6mg+P3GsVZKiKu33r+vVuxQ989tmWt964bxN
XhCIyVgH3aJrsPdLGC3JUtM12mzzn5dXMlmQi3PrNJP7tkAdXUT4lqD0Q54miM+NrDThWfADMT29
r1YOEF1UbM3uWjCib/PaC6CnRvVE0G+F+qFGRmULTIRBSay61MPm4B2DKM/nzYmr55+e4ajNFXY3
1Wb8RLMqZKYernEn8DEq7qN/M8b0t0vqX9daj2k0pOdu+QhUSy2Ks0TzLfpMOVombFuHc04BWAwC
Yqsq+2bLrli8q/bto2NGKEcasuf2FKaPQ+C1DmbludDSonOicFZmS/1IwHHr+2reRrDBrEAImH5u
GApCua5GoYobX1gRzBcXzPz1AMja9XjvhUiMkVEHRJ4Oo6y+RpRBjujl5XI1sfVFWz3m44EGTdhB
5M6Ycll5moNO0h/GkYX0UhLxZuG3qyjA1OGeBeiti3csSUoARZIKzEdGnQb7wJlRdnWJcfXRJ6CZ
KLeCPVM24ANoqLFafbk6nWn6FrpHJwNwZwulNDKC/GEcNChi97OMOf09aQhB3mbsh47uZzKnOcbT
gM2SFhNqWQtvQADKBsZ05BHISyVFDKxmopgSCur74AasGo8Agfd5xQX7T3Xep2bjouQymIXoafKV
Y/2TCZ9qCskfiRcpHMQ/Y++MqPQvGi1Va89U2u0OU74j31hUHm21rYXsZIHSQQE0+lXbR4tSSp9C
jN6GleXArA7w9UAh6Pza1pnWaVSMru7GFn0xuI06fLO6RjZ3NV1OxvMzS8VBB0U7QcqIhompZsXt
OQvHVSA0j0jf3005SyT+QGfxAwj51XAhhPJjxbUw9zbi7fDGHfjosrHdG5V1tfJneFemZuJ3Is45
C16CEqTGFZwj8c8rJZYJc+i8ZItQbiKoQG7JK/4+ERAhSLoKCL6LcqVi58dmNPKv7QLEUt4ln9Ic
yl7QiEZc2H/Qs9LVpvzg+83qewD+BtlMZlFpLJyPc9USNbqsskXOOSIhX1HRJY4eTfQl521rsqE7
/OcW3IKzt2ijNML7A0ZpxxnMy0v0fJqZkMdSCehbkFJQHwE6LcnX03m/feCafx3FL5sR2NyrM179
IJEVTOylZEQKcP1ERG7As1pk4A3NKXsLMRxVTvJQJI41U6+YQc2EDIOARl3nK9wG7qZh4OeFjHbA
gsR8yTiDe3uQqIHuzzMCBNCTX5HnU3Md/8TjnG6CWvRS4mYF8y0VdfZ78PZ5KGPdLnPV32ZljPmr
nyBI6foFtbUDZYl+Ac0VADxUD1B4zlA5TTKzv9ADYirFUPWvydqYnd4xVn3oF/Y5Bsda0zKIDiI8
owU7IGNDvxQMt3DmNUPfZU2QsLROFg4HX0xED2TBkQjQ4o+S53sJDn3ojnB7ipHBA+S3qV2Fa+zV
ISVIgwdP/nV4L9TqZazP2oSma419txlnfhbnxfqyOEhsQBJnbGC4SubwPXbgbfvYuAbR0LO2OPoC
P/J/nNdM2mnlIUVZYK4qgS1P+4gpeEnkzxVOP6cWK4x1qY37dxKNS1J11pfvhPH3g1+zUeHJS4/C
mwZc447M8UkP3d6M7bKrNx85BF7B0Up4vuYK3QiTmp7zLfA7V1MgL6w4YFrbHQXqrO70PeyRVakX
E9jcgpvXtpLDgtTRUOYqefI4z1ulzxn+Lp4vzw0ICBxx1csHVMIO+Y0L7P4eYalvATrQC8qMDl9A
OLv55EMkLkIWUTLbuHZrmFL67XnWXPn3Tw8EA7Ok+TcX+TLm467prupktBBrsI34YkrI6+QSXuND
otlm2ejg8PoZcsIWhuHnYtEiIMJ6hkwYN54TGJlD/4kXwiTrzyCCRluUheX0d+yQK6gaqC1/+SLH
h22e50Cmd8M8NEZHxkfxX+7YJv7mbRnUS1ZxwjLLlLUKLop6SFHDGAKvaLeaB13SFtqGQknE49BT
/E4hK4YeqKQz6+oaMFKCmOgTcPMePtkZYh02VRMb26AOy8PvrNLi7iZ6cA4CJ82ADB0c0YqwhFC8
PbezUh7WCFlfDrFlrx2o1pYUQ1Pccq1jHNpBrU1jnbgpf4yeaMvTAg5UJbtFpRElRLAshbTYumdE
FcyA0iW2hYLNMrVwWMkRPRIR4yRij2L1dB9QGSb6RGdVoCBJfz44JkJlM/M5fwMe1/1Rge6/W0gT
VwuFdGcJo+1ieur/SuPk9QXo0xYlbR49+jYwthjOrP5xxZxLYjz0Ldsgr8COCIN3AcEQ2l7QN7XL
B0qQDRF4KJJeQDQfvg3R9kuFlktqjuWKXWRDKNnZleBaZGY84mlqykIPfyNam9Js+SHvkjEKHn3x
hrWUj8DtpHbamSRBauNmwbEkPxBiA1TZ4muwGHyGUq1XqFKiIQjS4Wp8LapXO3AQmheZZZ5sKzdE
H+Oby3V/piKiRTKd34qjt0Zpn/R/cdy6rXPVQ/ogvOnngtv2sUzQM2e6ez6hXFMdeJREQpQSYaPb
qdZEERANhQE5pmJj8QRkcTBp0F6XhW+fIBxS6pwfOUIFld+GWUTiSznUgcPAiFDNBpQFXl1/Jvve
0iwx4bgLsnKWlmC5TASu8/Kl70nYFZVbppwj0JR9gHUO2XkTMh0d0eqMPmZxVvOezY8nlGK5NAsq
mwkvJt4ZwLTV40I4yHvhBqTWRAdKaK8+iTA4pCLaHYzPrIA4RR0vmA38tdxliFniFa8MBMXDjs4W
1JR103EKdm7q/0d/8GpgPVtlmvnqkPc74RMK9o4kma7Pf/qFmE/+BxfPq4OmjelXxnHXhUM4LJZF
agLYpxVvmO3EK73Tuqa19MHk8s+KJN5hN4K56y3FpBnQZU2LOhy96uguxdI4sSHy0lcmMrNXGNaA
S9w/x1l07VdSkzInxK/a44LEEwOZmRlrtuDO52WGvLW0eO4rd+sTTnZBkKaaIkkSCmIr2MR0bdsA
3p/1wMHVnGxYEH5YRxRvxPSc/KPZRo5/RS/P4Tcv15/otSmwt83YdM0GvO5KB+cday713zX2/y5t
Mt02A622ibidpqJaKwzMkptjNoTC+XoHAeCYfsXYdpqNY8jLj4t6hy9KDi9UBDqmSErDxRqXhjA+
s3GUlxdP2R/pPPcS61yiCKc7/6HSJ9tDO9UhjCSBKf05kdYW8ts+y3eEO6baLKBaoqk8DDa8EsxS
i/geb4+kbdh61oNhHHOFhPZdLzpeFcsmlJekGBVa5ITiQInkSTf3pJf+3QGxf+1kUCWQlaLIeW03
2NUtbTA9ZyGFXGi6mGfwDUnNnWUUH0NRRnyT+Vdr5pmQyReM2vn2sGBOdSGnW30pmIffaRVc4BCz
jb+JFlzgnmilq/ubuMRSWoTzLrzuPjCCUXS0E0TZWFUi+ca+nFL+5eDpQ8Utn6Y/fHDVZoBABDel
JrVCIu/p4bR7LpL9WHt43b+EYy82qZHHsWsbpxVHhaAW/a+h1edxWf+SU3vKSq/iPiYhYhar3KNV
17713FYgRUsHY6h0+5XAc97TSKyJOJTw/qoL/HodGDQq9Rhr/c3MeSPwWiH8XG3AA4rDTWxn49dM
gVWmErFpLLFPn8Yv71JK/U6x/kb/ShTIUqzgCbAnkBXXIyU5XGJqVuewFqeQ9LZUG1Yoi/VETH5N
vA4kK6Phe9UDAMnxZOyBaQviMb/QIVC79W6FaXI8u1QRRu/kbGCNjEqGVSz83PaNfmhz1li55dE8
6OLRIVD5rIyLbwKitdLEYDQXPPuA8PQjQhfHmxZENOx3RrhwU9WodDnR+UpEpq+x8c19xLaC8c+C
F6CYNp7J9PMblPJlLImbBsPYzmBwGcWbbF6V61KFbXU8MVtXGqF8lnFFfAR8N/WpLtflO2NioBn8
Q032HzcxCsGRiSCc42EfFw9nhNYqEDzH+sNPjhgItv979OpOZBzt0ano3u88Si2WptcoThB4XbO7
Pvix8Ys6DMTYBh5vKWvtGpQBe0rZ5tY8LlCp0tyFxa2mEcBVeDWQOW+f7C5Dyrl1VBS4ZO3JMiPB
aYir/eBDsJU1OhhRYLdYYBMpv2UQKw8jspnIHNq7/Nm1Apsh5MfAX7BkRD6s2OCc7WMWPBmmMEfb
XfjP652WGGp3icf/1y2cTZCYaQ0uPntzi3Y70+2ZIxTquU3SF9Ad4cmnAFZrEbmH17fVioZaopGI
0R42yKl/M8fEmWZrcPHJ61vURQdNEXVkdckBiNDlsu/vUbO7WISUVyVqwbRdIOhdVtROpGszCNGd
vX6UIozA0CXmZMn5WW7ncapsOAf/aHWiBOLBVD1xWQ1Cs7g6Cc30d9lYI8kqoblOcWZiaWXc50Iy
bFm1wSVgwvmFxSJ1D9esuussHzDirVGbRzXWfbInTt3XCPcyxX9VsKY3yB2p7YyhPx/CgGg+AUp4
qn0o2FHdscQ725figAn8IJtAF05YoxMFsatwRAbBEmMffYiwYcSV4UBojlo28yKqcQtFxgNoIVjd
y9V/Hub+tkiouTyWCuOUS2URyoSGh73BUQpvk33QuEfA5P0EkebyravMi6Bb9LEoyMQC5sKeapsb
DCizWz8UEFM2PQSZf1G+oIzfaMXrLopVg2uqGjLqAYnMJpGVmFkTowO1LkiXYlkIA8sMALyQeuY4
pjF6d0EedKbOLb1xwsyGab8CVoL+Hf6peZO+PsyCbrgGuUOqBOBm961uFNs0O7MvrQ0LSk9mXXd2
a56SgjfD6I2h/g5lHBGgvmbq4nFRiofWfXkK13ggJuFqOntmVwfg5vZ1Ycny9H1p6zB8b/hQAW9z
M8Myhfu9Wl81FoSfB7X3q6Qc+0JapCermYptnkF1BBWlrbD3iUqBLvFwq1EJpB9bVaq06/xhlLsR
vNb8U+WFp8HmCxQPHa0psC5b2qnpgsmH/oj8fiCVJAGZMe9R0bsJwxWv+MwxJpUIUbzBa8iPyeeK
bWicrTC+Sc1FA+Xjkf1GxCV3YZu7k35Vnu82RAykCUBFjtw8A4b8/C8N4mJVWbvqXGYSTa7WVYNS
Agft6EwraIi3Pm/N4lbSyWXd51xYockh3MG45LLtOMIXA/H0bDoWBRo0I336x87ccUy9ogsvxKOu
wH3Qn5VbsclHy2b9oPR9EyBFQZFlsoFV4YPkkNj0WyhhbZDQWct4tMqX4nVpw2S3fx+HNtvNlqIJ
Kp9zvd05p74S7CHhGEWGnWROCDEVPvNReEVOFR5utZg5NFGFwSHr+uNYe9SsY126h0LSKJR5oCOD
0wcD03u/wTQpHhgTw7b/TsxpFxzSsv7dWR111poiP9DKS2msRRnFj5TM4luypl7vriDegRXcb/GZ
J8VzX01U+YRRXAd8ZW0Qy7fGYFZHg2ZLuITX7BSoF8zvEEC4pxTrW7d6ZTJYPCAzunYBLh76l+xO
vNTcwEVuHro78F1lsId9w2jfYEaL390BkyrpDHlIJMXak9ZrIgzfGWeRR6Et+z0HSJnljDqQ9MmW
Du9TZ2A0+us9v1ehxjoRRxPvJkHr+ioulur5zfZS3kQHZE+cQwkZ8VzgN+HBI1XQXK8Agb/CqX/D
JDUg7e5FMm911C0FqUKYXfq43HEjjdMx6g2vW58/3BNc2twNu0gqp7b3IlXMa0+Rn71ZV7uC6fI6
u3iH7PALdk4mHkSxkGPGHxNL6FKXK1BBq6i6BWjXZFhARmAscvNGZEzdAlHEY/IhmLecCFPhJUsw
9Mp2wUNiClASvwvhbEAFHQFhXIw94xRyMz+hsEwAt7DKrRj7ADT9LC6lRuHeEHWq3FxgMp2DWayI
ftlG7FNgfeDCpTfZMbsB1B4O0TnCFv3eIMhHECgVDleu1VJl2Pn0Ev+WAkIy/z5p4Z5lXR75HeRn
MyxCpCcf3hOpEQihb8+PFUZh4NuH4bbnYWbDbMUMAbqlmBgtImpfCDsfu1zSMUCAQRsEFpgeYu+9
3mc6jNTfHwgnhrUE+l0SN0crzW5Unc/Hxezs1v2KOP8KjU+7llKC/NSJdOgIv+YotVvCmLt1sFVZ
zbsfWOOA5xqFII5Z5/NFPMdGBFjBpD+PsqzhW3+7+UC95fgWZz2HvLk5yCadXivVwhNVtN3pPLOp
PWZWtzpPCjK/Fr9Xiki2c4o/vU23yOZMzSJbLXMlPJrOAhJGOjzJoJnQchtu9PiUlXYa76/XigIk
7w4NkXCqTWLfoZdqJKSgI9ZGLGbp2WyIzZ1soDmSz+uGaYtD+ThuqRuI6X7FUVg9JDOjQ7fcPb1Q
x1BF8WXWv4g8QG3n01NTaHOiu+XwoEE2Ij8/6pc60ig9QYSdyARzYl03QTm4XcfsvvAbUAuvRSDd
Ieq70dPcjKhhhhUIXV+gIYrfK1aZuAy3gQUXshC47KwlpNlzyY6Z42gDiVIPJAYbS4EQcUidh8Uj
Y370YRx7pvBy/7u2SJGDp6aktNRBMOZpDtv/cbJ4/ukzMPmYq48tFVOfJTfsr60weTFKwXRiT/cv
93Y6C5QMv/vbGJ4khiGgHGqWyQj43ZwzJnR58D1AHgiMx4fsA5iaWbOTQ3iL+43Cl8UJb5GkCM//
/BmXJltoW/Q62QcxXub+JcFSKOpOAjj1Q+azC4QpPHK7CGNxVR4HGRYCYuZo0G6i72d48+5XhtLr
U9PwoPFNWqJB5jNAjAyRfWoj38Fu8wEvH/1xqiuamg9LSaO3JgsiGLKMbxgxrL4CEdgYQYgfWUMt
imX/VVrAVBxbvaYRiqs/jn3q3/PN8o/FtwXOCct+BuZaYRdv1rqvxpgQoSU3bAnlumIq9bM4lC7s
W2mzpxYR5GD1eEsqrEo4V12jmVcNZ8z/rIrDqIL6mduP6FcdbwoaqAltc28/rAMSVTcQXSf6Yf6t
5BktmG099sZs2Kbv4PBqAoKCcft8S3sm5VfmU4AuajfdAfAx9KNrM72C9bfcieC+YAKBrDHSeKCh
vgeaXuSdi9oYW6KHVeWWWqEQSJRpMIjB9vxVlhyolsv0J8JJJHc6T7ihG9HmMgtkbJhj4YNPfXx1
TU5CUyjViUbD8KVStIt83YbMlRgK5DKzWYcPFoAys0aw04AitBQaTh8zRnX4W7jfDFtExvmq3ego
ObCDLAugIX9P+C6JEM+f2UblIFHTVOwaCy8MyhCQvkciEe6hCYcNQ2yEDoNRp2LwMJaH8l32xrt3
icAtOnUL/81BGuGrrddgxs4rMqoyUc6BoXii9FrcQydKK6h94NuHF9otukfSurs3Pjb/jtQU29uc
0THB0BmcWC0rmO6pSQ903zC+Lsur5MzFuRaMqQHQrnmPEIxr/14nFRaB+4ftOdxtrScy018n28ir
/wL2viZLKSaZ6JgyILzgTsvMuG+HaOKl+Gnj5fhvH6GDe1rEITtaqp+FERUsQNdl9mH4rEBrWL+g
UV1dPlA1YW8IZSX3AQ4QKBhTWTubBhr3Nxwajf7ZWB4T1iL0/kKGCTLJvgREX7sSnG2uCwtcRy42
2+3jOpoFzvdnTUPFHv8ZtcJhei8vsoFiI9JsyzHKFaGFVPbBjzcX9xGvgFF+hKvUiCl+ellmLz5n
nbJJfjASqDcQSwAZMlE/E/h6JAq66Zyepv4RAhdeXz2xdxYOBJM0iMpBmTmbJTQTGkm3goY2+9JX
FKAUttpuGzNSRJDqGNig0/4kJM/pvdPtSYTl8SA/kgN3WK/teJMCaLSkTCzCt3h5tIwrxajPHLH8
PJgIXk5sojW/K0JN7WWidjCGgrNuPL58MB5QDxKsRiqCeML9QzdsIAdOpLr4QBpAp59b2K3Xc140
Yk/mObD41EcOjb3u2uREqanMNYe4E5z1YU9y3n4yOWubNsRMvCxi9hp+jN1fpyonAnaO2LgvkyR+
97UDyoMxzKANU2uO7Bp5T/XhK9DUG2dxMW/N3eAFiemllE2R6dUZIJraCKwePM3d7IANYDiBGPR7
XEzy5CF9WAor1omywmdUfy8O8jo+JqtoX0IQczGJHMQxyXPbnW1T/6tKAM6fIH7/3esi3rvxauW9
0RVTyRZTiO2LZoHNAbIA5dsVe05E2oBUsi9KKeGdC7q5hQR3Xsos/QuwxQF5ZhrqjeVFbcugJjLA
oyCu4uMhw6cF3tgONhfnbVX6CdcFiwKY6khbDBfnPLLVDTZCEdx4ZZgaRNVDHUQDugiCFNYpu3c/
TgdkPZ8JLqefbGCh0+cSut1+FBDmGlbA0niGnys78pFudtj3JlEes7RJSReNeH6kE4EsExlGk+Kv
3BonjMR+6MdNfjM3vv2N35opBvPpVkeYCcYSJYzxP0F5Vx83MDQpiiJsvny62H94KwnWksjUPQgH
90hmaMlizKRKhYj4zRsNWpnmpLwFedwPUetD20SsYs4BRbs4hE2sK0SeGCnRSsteRPqqRG2W9PB0
oUEGrtWdAbWMa3II6p6SYY34ypZuMa9U2wccWzUhNyvpCyV5PQHHjJg2dn4hV+1s7pi7rIjCVAN0
YvWkdHldZ2rWjAfD48dlYZtU09F7TKAYfDl1vsZUQ9KbYcppNWP8z2O104eYBo9qN6Cje/MxtSbj
tt2XhcSCTXoLhi5Lw5270c53j1t4UxLAxeZZEOXnkK4xBx2zpWFL5cTF8/4H4Pmo4qI0sudjuurY
IY/y4Cm72TUaDcyDOYc8BbUG2odT3D3nNoa/mjHhSIhs/YAPn0CZIdPopLTDInbvYZbKPNd5Z0Xl
u9k88tQV2DJ9j2E01MZjSb5uKFJfhMZxuniQfXGzfTfB+gmOTwNNNdYwJSBaG6zfwgrhIvHZRuuR
BN+01wQYLyJ1CNJeBEqHF4FMQbzGvkyNHiFRf6fO3KScZU/Y2dailVjghsFBpjmpUYxQ4BspnuoO
L2g6Z4VhqzxY6dI+VKiD5diF0yPfBq/J9xtJW6SY5T2s7cc9dACsPOnbY2UHYdgFmPO79Txg2hFs
jEY9P3IAtZQbmwlivjiLGAhn3JyXkNyiIHOlR4A0uCgrUDhkcOQZ2PZnqzSPT/o7u0w2/RG9Rt6E
zUOuMEC8ns2TvtwJJB1wjmfQy6HYKRkLTt1RAwEGt2fnrYoPPhLGAbE2v4SIkJTiCe6tQOFrxPTK
7idMEVXU1KTW6QHKY7VO25IxijyFd5e3zcQif8IronCtH/+HrXaD+LAv9HiyqKrHHc288cnWvAdv
LLi95xy8QVkiPHTn39Oi07TwcEsHSUN9sYq7TLWoZTwbLQHa1+uV59kGyBpR5TP2RF3XSTcTZSR7
1Zss7z+o/gj9QV/nONRaRcQLXGJSlW9N5iFYvws58MGUiEyzhAcca8zBGE0aIK+un+b+JTwdsGv7
0LkHaD9BH9vg0eECYEOo+rhLpqBnmmBRZ+sTCYhL3Xn+e9rorIUUQxfBNrykWA62X0AiYyhBKgb+
hYSsq/PTgA79zvCAyEoVSc4wdvquriHlNfnJFti6Xin5LNp8dyibNI2kJL7jauFwlEQJhikej190
r12jSbw32XASAEQ54dO2UMQI90V73SAWsE/h9LlcZFNSilPvIypHvd8uQevD7UkpQvr6Yy0Q/v3I
1MNmrF7MaMt4Ie4ICkCq2iHViKg/uAIx8L5gV+xulICB8vRZF7m3YouidteIAzaMWlSZzFRrkVSv
Usi7cDznEwVZCemeQiQDAHBy2IQZ2We+bFTaIMckT3SQiZBRglOdiLT6vEyCMYvPpZ8T9gGUaa8G
S4UwOlV7KelgYN+P6KqTTKuj9ZS13zzlCAhgdEhGuxDXCE17JDF2bPnueT7X0O1Q9UoTMVAwUJuu
IA7hMKVMXh/SlSqWvASoikj20+MDvP/j8Kt+XC79bzY+SHRJaj3D04pz1YFkVhiN/q1VIFRUxhAk
JzA/Y/8TIF84reeyuMgcOFSST5Tzmd0J4unhPq64Z1q5CWaNPlW6LcMT0CZMEg84w9Jtpycd0Dbb
QQ0YUd9aT4elRz0tLgCFZgyv3bUdeuB+DFPYO2hwxLinE2CgJbZnWCbd5xaxJE1tPW/bAd2ndY5z
rV686CO65l3MgAIoUfiNgqhYLSgqePSpyqOQjZNu0LnS/ZHgQk1k+NqanssdCGNO1DfMrHkMGpw2
10WXTduZCvRNoBQkSMXWNUPO9U509daidL8wlAQ3Ef4Kk4qAfm8KBiuOQ6Jc0jhtWlBSGwVkE+ej
W7R2YU0i6f+T60KpUItWGplY45hUrXn1iDOYIzreCml96hkEm3cTKD20ABnPbFA83Dx0LWnBNRs6
0EubuHSZXwpyx5CHKojIuraSnMHUDdvzN9qZ6m2Pul2SUbxp3kNy9QbBZfqTP3+/09XpRu2FhL56
UWOXhAHDezifo80boCEFbrqvI2eC21/joYegpgSbOFdSbmFMMfHcyvUwyZKJ0Ajw7ZR/XNI5FdOC
qa61iif6He/2j7eccpx3o6W6bbOXQ15ZwaTtjrY+F2t3pRU/r1k4lkwW1rUDk4PcKMwZSETudW1d
58UskJnodmzAauVUNSLd322AE7fcfBNDlo5Mpj44uqwfvC2T4FaHW4O9KW7otum3L0QNW6J7aCoX
14zQEU96HiZSDMqGsAC6Cfs6onBielObbNPkcwV+yKXdL1410TKWLGfp/mdxeYpogzKS84MVppBu
i7UcPZJgq1WNpBdx8Nj9fFAmCwLI+EYhmw4S2fQDhLaIgzq7Aj2TseRUDytH7pMvj9KUQthX7hp3
6XOD+Oc3QEYuWBOmNNiJ0F4prLP0JyNFfkbnW56JnOoehZykbY+xYeVpfLZL810T+wCgCoCCGFSq
gJJAgWdzadG1//0k+efnhv9sa0PZk04kO/Xk7iE4Ruzk1fmD6cWkmltS3HUlV8bnBQGo1Q+FuBFw
/EZWBxhoDPlAOxbk9UwnV0rHGoiTdobIYNk71gIx3vXB7rhHoCCmzOHW4srqSksOFSBPh3Ix2adf
yeUP7aSlV86FjqFes5enGNYqKKxdlQzRvQsewEJkRiKMu9ee22vxRoXkimMhoxEb5FPDXJwJf+4Z
SAX1BLt2RxvvEnt7LMcjJ5LWICk0yJuy7GeZB8icOZe58S0ML9kUs1y1dnAzAacptzCyfNalmdmd
ddweSn8z/mfBgFJ7WOrHb8Z1qqAyV8QqpuYleYOCYSPrjOlaCYrCIawTOAJujq654JzYKHCd9Zhj
BPp6NVEeuKEEw0hg5kjF4m4vLqHt0gtgxw6B13MIgfxB+aPd2+1N4T4tXPy0OxyU/qL7DaU0cx4k
0acwbFnxYt9+0wDedNMMUsX6b3b8RVJsEp0Gm15C0pG8qDrvSHpG6eYnK8LOc6djHqdCLsEkWUy4
eaEdKotdDRoNjc8fd51viAcehmWElBSc1t9nzOwUMq+RupKJR+Hp6JBjWIk5iO8kuuco5fbflY5Q
hoqVcF7gKlUYKBB2ojAwo/9AV/SY2Ta6vgFT5WZBH9U7/KoDo4ev9Et/eg+u4mn3so7x0+PAKVqK
UM26INy3/RwehZP4jTqZRpB0JzWUkkZrm4yTFbOecDNyGobuGtvm43MLiQoHRL6GYI8ZrK283acl
oqeOmb8mOICBreCF0KaohezT6p23N2KVA7Fz0PFUL6PF0ClvqVzm1fzGvkrK6G5GpbG1VLqX/cXP
8sUA9DCZOg9R3btJ633jHWb+45QijX2UG2lNSXN0cGufW0btsMW5glmx6/mUusqUzwPvr/DEmkYm
LciNUKP7LHiNeQbrOvB5dFLDV1jz1+fctXJuKCUMfHMZrsd8PLpiIhllCtXE88BUw4MHZltXnnov
TehPzSwEvMb6d0CT1shVtWLIPEGhh9uVoBbz9Y77hA8Nh+pnMfMYyZGAo1MswvF0IAvlHiJUOnkv
HK+ctN6F72AhgzBpYs18ww6V/mxwSqy3kPndJGW/LUrepYtRaPLneARlh+AQ+Iw70DtVdDbENyPH
bxL6R+vPwMZLV3RE7tAJ46auc2IB2RFrrO8FdejHK8b6WfhOs+YYZG5rgYYa3ObrGVMlORlQC8Sj
BCmzYYCp41eQKUBf2CmVOHS19z2EK1X/WIqUUDsSgt2Y+BZCB6p+iVlb9GRkrpT5Ean7gI97d8Z6
EDCxMNJpXb13ORal0N4jVLqWAdiviXpTL+cyN/SxzJGQrIsa0GwvjQIjP1uS/iMDCxAXF8Ocw8mj
ghgM93yl4bBStR5J9mMH3ZCxIlb9Vvggei94mU3cBUL6K8TR5XaQbldwLguTkgsiDhmkb4bo2Jn0
9h5BqUjHA94YJUIeuI3X5+emxmyONJtGj9jUZXtQidbnju7zQdaFCbakJzoVXpIUrDCiActnAKcW
kRPgg6YVNV5QNByTZbePG+XAsgelvvO7cjd6OJJAPNlO2GQLapF7LB2dBF4uMWcHphftrEzuCt7h
Tk0DA+m2MUOg2r8/4uAKsnoC5BHR3YzX7XqjUy8K8bKbqMp/fG8CmicE+WEJid55m3PLeRPnjeGo
ULJFrdTQYhum3rqenE4/KGWe2oiV5yHb6vVLpWjEfrTKc2SXDKbck7HY/1vXrNnDuucfGC4IqrIl
SxOMxz8aWu7QWOLJzETs5S+KYOyhWOsynno9wkih12/y03zlk8e62m6Qhiu1vQNgH+k84lfQqt8D
+c5KMWxHQJRd3yJKb1RES9NIPSk/LKM53r62aTSUPvid9CBi7eUa9ys6iQlSPioX5Iml8ohdOTvY
Bnx48jILNBHbXSXqJMTwZBJLoubWjo8KU8NpdTB3lUzxsF+pUxcAhRN1GbYRV040LVF100+P98EI
DEI32A5k00bNrV0XjBElpgWrMdjqWzNZSAmigP6cvBMUelXiRhtIr6egw6X2uNpAqmB3tw7+cF1Z
RBw7JZoN4sBvecoaQSS/3BU6h86MEnV4mqun7GjxW8+lKyd9t2sJCxzke4Nr74lBYGlQyiFvirMc
7AuJn9245vBrJsyRZpVhCulof/weAc8f2Ah4C/RYm3rCD4WSSf0QAldN6nmh/FW/yvQmLg5I9rFc
/vbiV8DI/W2u5IkqTFGrUrRnLMvRABuSHbqkCXDThj7fz0Oy+p5rUMgEhtUcdeiKrHFz07nNyRG2
dLqUmsL+sC3XnvdxWEqDrSbeoQMhrtQJegRA05COYCA31tPRskJqH0O/2ZYBwPFBT9t3uIW1jGvg
am6bexf12P2JhVvN53cl2bFTEXAV0WOFTfthdZafD1qcncd196hAcgqDMJKd8ZzqQ6Cs8NC5v1WF
QbsdLzR7iqkOzfuMWKDypntMJvb94c6SNOBEW2kzxqpTx6+kAWU9yNLLplizi3TS4jLgSlpVL7hc
m0HwRqQ7bzNnSnrXO/IULfv/1MY9CLAc/XGlCtmIoEmqES4XiZq+Xn7wpK8dlNhwabUGCiWGZdWM
2QUTXYgjWVZGAg4s0S9B9nKeo5PPu2YM4C9ZLLfbMpPBeI/+ymGpimAjFlmHDUd4A/sQhuemslKx
vg4yKd1QDi6fTw/h6Mh1J/MttJF0olTNg6ae/HsiUcW078toQJj8BTQle7G0/8nfSfJRs+elDeRm
5yVvnoVsx5jgv54N08GXv8UZleashnLJnn0Uc1n8/MzXvikh/QZxpZyjucYVKf6451qq2rsMqi1M
c6vvyCB5hcmrTb6EGNWACcZVXg6jMY2DZlgo1fCiKq3g3LCvTrJMw+RJpdezVYoLPHoXPKGkos8G
W8K/cKVnxzrX+cjnmkr4KzKADcCWHVUDO2LIdN1vKxjgozCcx2X7JtZejCd0AAYW4694vx3ItZ4T
zKSL1DBHITitQb3wBBn2FG+G/C2E3S17lVdaUjkMOVtfvzZ+hCRWqndn2Es/ogzve+Ql0T/p19jC
tY4glMc6TCkzdviRbHWkN/IJYABtHYoYoU6fGm8gEg9sAKe1emEZLJX4nbWqqPrLXyJ4qUVevf76
gZnDa5WpHQfMVh/7VlKeyShNeYr0UoTvYIGVQeC/B+r1qymfTxj5apBMWxHLBHsJdGxR7CkZAKoB
YPUXe2w9V291Cz9RioLJvLZyyx3qMZTR7tIKe2xxXxmZ9hT7R9SKLLGvupaIY+ntFG6Ox1XyhKzR
u81aPvC0HibBAQIix6Alvttfm9OOR/F4MDuwOm0d1/cr9EqHDC3a53+lMXJ0u5rIsVzFoziS/jJx
YMCUaL3w0jF9xnKOIAXXCd8q5zyFbKZ192OYcB3IkWM3rAAY7EtxTS3PzLYgJ+1rtRasPxM5IYcX
Xj+koO8z/xUHmrPGTqbUeJEZxjkHvRmt3LswuZUKohhxRvdNsk5mgUUoakDBzC+b7zoPaDYgjDpj
jqa2dwofQzHc/nwnSwSy+1SGCfYSlZLT9FUVKfq115u6fyeXjSyzfp8hmWoq089WRpVCd1ErQuV/
OJ7g5ajLkdPpsw3bR+SBsCMpDCBSL+0k4/JE+7HXS//88cKLgN/b2hVJDVJHOEE1yq8spmBzFCn2
zIRDVQ4vakVhniGQWZgVubK2A8eL8lGFpMgu+//YSgE6M5ha/juq1caWXqaNrz24ee3IZHFCfZzA
EGqaIsda1ytL1rxSr9liIyFpL0veBgZMQwrefIYMl5qdVD0+BvomXV83ER/7GvDJUemJydavKYdU
4bmNATazxaddzLlIJ88lFT5nS6n8Ta7jOIE2jiGlBQHWmkUchfAiieynJZBD9r3p+87o6kZvA4Wn
fzsJFW1AQVOB1VEEg4/9gvJgK5CfG8JVR3IiN8w8ajP+tINRzbMgu/bVYsrqk9FGvHjqvpoiq+C0
WG1pK58bLVhGEb/pBMcywXG7RD+JPIbYpUELLH3hqGHFSXj0mazXjKPapjhOvOS+94Q/Yt0zN9w1
8iyUjbiy4VKMJvY/8tOFSoPnrwhrsiGC6mho5zkTLkot229JH2MpeM6ya31Vbd7Jq7s9ajPtppCR
IGxv1yHqQDTmF5elZ2Tdv6pO1IxyFPyT+9RhppIp2stbo+L/j6uFMFvDF9VaCmESIlbj4rCn++jL
/ZBkGuC86N48ZK1QlE0MM2fpFyfiB0A8N/nYg4y3t9sXwCvEOCdECvkUIvIk0I4/h9DHT1caXlsY
tWkh9kn/r1aRmYIf/Rv0oox5raz7Yv3zknj6DXF/ZHb/XVbmYW+1d0rhiHP2Lx+PRBsU3Ka5MZ/F
iYPafVQEFLMH+sgh22JMoqpreOpWim/+XWFwvUViw5JKd2EhnxKCpk/WDB5Wt1xA4vCJ0E5VwQV5
S1VMIopKYMUeNyRqI4P+o7/rrVK15p6wiLYYqBPar1prj1xBy+BGRXMfTJXPYPaXkuNpFLtuogei
QR62gFHZ1BAyaU4EG8bfSSwfHkHeFKAaGqgtP8GxiG94gHQVi/k73cXYCjqN4WWAT4Vr4PUmZrPv
boKOvlVy+YtgfKIfjPWY9vziUyywFjhNj93GzB2RWat3TqRoWbTBzPImjUaw4fEBuLxm/4jAhu94
r4WR7F3dRn3L0BD2MGaRjugFN3+1bPn1GGayNx4ASysL+hoO2dnX00aCES3DcEepNUIDdKsr5Dl8
fBq0n20inZDBCllRGe2oBEzlsH+xRyGrdajb3b2QECkBitfEYLYbEI6OeK7mta2lo9ywJJGptJ/+
nUHoSWTIymzfTOQ48HNb5o+MfL6WLkM9RsV+bu4cdSlb2fqZGoyMNdszLbBdNam5PiH4d84O666G
RX/bAq8L+Xv/etn5N1TP2FM9Sts9P9OZBvj+1HXCFW4nVCnE2IvNCR+lnlaf15yrYu/9R9Iar8vw
w3BfaMDcloyoBaKk+ku0tLJQ9z6elzShO2pEcQOk/hdHbUg1KX1es23PYfkdL6EWHtNMHrbH5YSz
+jc4mQbzcKW86eISJLVkn1rvlZ+azJwB9Aw1Bq/Rby2pBmVQFECq+ODVVicPtxNsTfJmdVTGMj4B
n0AZX7wF43znaZ0h+OvLJDahiKpoPUnEITE/8nXRvKxtu7G8WeZOiwV7DShjRWQt2FmHpslqgE0o
vdyTdfLPGYofMRLL5EPe0UjcKYHKVzyZSdx6dAT/1RXaTQwDtNJS6JoQqCDazsjs4/kp2AU0rOvL
Egy1yve2VPNOyENbC4eA/4k/On3pSVNuPR0HQO3IHOdDUkejeSTSc0Iv+zwFSEiFxKzWh+hj4oRF
0ntu6szhsV7+Y4DluYEDSbH2KqQWPEHz0iF3vgPtXtySnMZYROl3sQ0GZ3LbPM3FWvDn0W5YAQpM
jlanfuevxC6jFu9wor3hgWJX7rTYUOMD+zIi3LbscXfMiLQ2dj/l5tOyuwJ2q8bo/aLlfGprIDOh
tkmW83xQecHiOfsBs5Yj7aY08yEBDDpaPZpWwHJPLd5GZ0zGSM1ABzF6zFDccnJ8oRrXgmdl2Q3v
TswgJGn/1NS+1gouhwSmahA6EqTAX6qvUVLGL/nETKxxJbWvSoiJaRupq6L7fjQxI2wQmC98DQU6
yOksBdcc4csBuXP9Yptl5tGI9WhpFitpNmlQfdhId9b2otlQuzkJN0QKVCxeOjXUp5xWJxuA4uwO
bXY/w3jg4vr8z9FYHVbAwBRSfxub9OyTBdPda819M1lJQAOAWBx0fJM14ecQ+7qecdWh9SualrIh
Ow1Dd10IVFGP8CoheVVW5fZ5Ys1tenitWOSS9/mWc+dc9jzZKKIRuW3qv1gRKB4nk+T1/5c9Lq+w
J8Jm8gNOgLSJPn8RHKUzjpshgmDxJbYdt7hDNmR34lQs9IgX5HrOuvBzMBSM3G1QGl8Eo220cJhK
MqTa2t2i2qtj973I2jGHNlNHEnMfroa6YUuhXY4kGxuZBCgwoElOG7UHz/XRjEjlWuRQe0iaRo0I
g6cb/Vqf81cWS6mPla97zxC6jnA36F9pYy5hpUH/NKemHRxxKa2zeHT1w2EltFEXZpiQL4PPI/XA
DbjjT3l/JqJt1PNEClb+NIqypVtQb2CTbIEPfBGTlJnIwzo6lkZY3/AQvW5i0w3H2s5o+0P/73Hj
mhewE1hTpSbgOv+0z5WEoTmiXIL1mY2wDWtJrgXNL1r83I6zkZcHhZHm/SGmcygiCkDSNd64Ujw0
Vf2EE0AQkeFCErmkQQincvCtlJXyQerG/sKmMgTeUTxFzB7uCV6NtsUJR/3pP70golF7nFN5Raxu
AXRMmmpHUIjQvsH1XGWBgMtvcA0mvpnBS1yArwR3HRfSLptl5hkzd4oWJ3GVGD6V18A6wfpLSeG/
MoJ+E+hWJRQjQSvEx9R4TXgUONAxAM/QRaTIB0daBBUs9Rt1kbuvArnqphD6KMOgzMDQH+tIiers
Cm4SWejXLnHJNJbTyFc14vndZoLQvM6MhPRkbvGZmsCTBix7mJjJnP+BBdARBfNHStgdW3AIFm+n
QlwdgsCdupozxfTXLakamM283XcwPN3eKV2ocyJlaCQ/Njvxn2jPIvNhGOX8q8VJ3VoFCJrwFYnf
2Ujq8uWbG95xWHazXApJ3p1hWXOq/gDqkhYZ/Kpiq3N2snXLVhk3zGeMsdsNhSA96bIPOHmdEMAM
BF9DnP8OUMNt2aMDCkgS00cwiN85azMsNM3m7dUJUgKVSVzxmAvboKzfPay2hOiFngVjg1Ll84hO
zaMBTD81rBdGca5lm+vXgOWqi1JRUIH7qamDk9VOitN/w4sgyjM6Q+CrmwxHro+CUH6yaQEVyLxS
IopcwXbVTXPzuIHJzvOdIO87b1P9kaQ06ojjDNmFwCY9T1U5wEkAvNPxbmxnixwJRuyW9o9Pwrqq
cKVyJhdTbrFIRlRKrmRhg4ty/EmZX11Z8s9T/CaNB82Yb8hFAA0881HeTqpltDp9slzaE392iOs0
pu47ElgzPAgp4IBbQVAkN36k9oTy5eTjb7AbuBSkGVB/+gCB9FMR8nYW4W1dVpAjKcZya0AFuUKf
Sg0rx05oi7OHKHLVJCauOX9o7cysfZLt/HOZ3GxkB5Ug3tDgrZ+Nym+XrpBqTgEmmG/nSujcK6WG
jSnqGPYICKmkWn0xdYHyfh08vbCLDQ4o6c+PbiJaLgeJ7EKZs6dVTe9cisAQAXL26yAljKO1JuHu
qvC6reBiLOew8ythZ803w84kxn6cOUq7T2nGeMqDez+W2ZCSheUiVtBFYRru6LpiIxbOM/5Sg3CB
RdaYygniI5OIbQfC8YLm3C/e8KZdoDYysFxLsKEjB8ggxiMNs7wTPom7n7F80Ad6uCpMgyN1w7u+
DUZpT5IPOMRBk8AWOEzDNIPgW5obnqSbs49CLPWsiGnGF4eVPouthYDZwna+tMQ/rEtPPog/4sKB
xvS9kywBnloQ6+k+ds6WYccRBTpZVaNoHQ7eOM+zG0ZVDvmmEOfCE2V3C3yubtE517cvtTX6LaJw
JZ+cFyom2+Oxka7ng2YyxDusa4XCXMapxrkSoA5AcnaOE6Becuvf7ufUBDReXscEX8W/Jjm9IXOt
fw6rayc5mP+8hz3UQDbwIZewr8aqPhgSbExgDb2XKzmusMOnf2kLlHqOskHeQwhNsX2Ob7TNc4sc
kGagKPNuMlsNOrSls5pXsVrKERutWmVHJY8qROz+YSOJlkNQ/i+zKc2+HOxO40OPp6YO8j7SPNxk
BebQh6PZiuQe52P+DBuiqdL1IHOUw11sB8Vgx/TIDJb4FPdM/59KqGBbKgJ6VMOvEf4u1AIY+nFs
PVksJTJ19e4SO1m4jvIzLml7SNYvB66vRL4a8qCIPnGqPyuEVPbMdiqEPt4bFuEQu2fGI/mY1rHC
KGObAypfI2dRO21qUcXBjmnMIkmRWHyOpEdwb0CmoLQgbZpfH4ejYgIIzPvTLa+GZ3mtBTO8dIM8
ct9/b8/jJssTV3jCOz6oaiHKtBQrkuUWvICJRqXRJA4Bo5fZfqLPihqANFcUvkxSOCJ+YI315ray
VGmNLB527/+btBY3rqPjM4ko+b9roSx3UwtlxIVGR3pkRyS/Syv+c7VmP2Qu/4cX33xOaoehVBBV
jWH2selEvdA1OqNfgcpQNotHgjtKYEScJJGD6+qHc91izl4NOJsr6csWfMNLBpeS2T86WNQLPsZl
abuYM+kkHT0PRzAbRtKajULy5KzXStE8xd+w1V3oEhfpYXNdK9ACsFohA6OZ8dLsZEwBSGLajQuU
DGFyOeQ2/TT1LkqqlTm5RoAC/CpwiJnb44vLOtL2DqfkN9oVE9jm17D/jBZEC8S6KmrMqd92S5o8
e516s7uFbU3296mHZpHR74zZ7qsM1xqo6r4Hw5JFHUzFaFxbfwo2Cde+qLNH9L7jK7fQkqgO6XBu
6Ml1vGHAIqcbTS8JdoInQ4ZyxvNtUI4RhmDlmKwsIhpmZicHN2Q1znR8QieRHtIlhTWNymJPJb7+
ufQL2ii5xb5AnOsGeNgbrJgYBmFkYeRAwld9hWU5/nKlg89jd9lkD89NIrRAlVhtTWSmFfbJRX+S
hNJ1BcE87qdjw/c2chhpuiJs9Vhfs5NxEEqReM8gfxjb13TAimWKvdv5i3ruuk9Ms4xWfYxkdGKO
36W92c1wVD/ovka1AHahlmd31pgyTydtW/Tg3BHj31PQs5FsyQ2IPiZ0lRtakI588A69iE3MC2GY
nI22zNBqB9k3bF0367m25vj+D4sxek6IM7IeWQYTaIxJ553qt5MmLvfDqCCR4SJYn0Y5heIDWAyP
urnnvD3G/IQd6SoTe07qn/ilRjLEEHFgWf2PD0yheUgLCCAiGYP9JuEiekJRlE3zPo1S38P63zJc
utPbwS883EwYrTX6utu62zGjHfnv88x8ZZAoy8e7ur1aPyOBy0HmjV1igo42LXKcfvX5CCjI4MSq
UDixdvhQzpmSFQZ0LU/ZxsGeTR9OIGLE6HUDTboJFQewjG8mMKUuR3g84C1Touf+7M0O73MmzDx9
9ih5RLWST0QK94Swq5E8TKxzEZihyx6Tl7YdGQAQ3dQMJ8dCOzggr4DBvh4mkRBeztsGwvO8APYS
iukXMsOq6FB3KGrGUD02pLWeEcXxBInBI7AGFx8eftfPCjzspBDnrVsPmymTy+Vp9eZinkoiITK2
ek4xcdllGm8pI6uuGQcvKm1X5/NZqhBIRcRBIoxyE5JFqsyunIgVCg/plF2p8OE44rTLBca3tC9U
RJM4VVAb713qS6xtxmhL9MKGeYP13UvA6oGX9iBCOpaInTOEcrLZWWf/0S3ivOOj4wzuAD3iP0yL
4muZnwVbdHFHB5bf23cj85K1VP0LnYncZ/jYBB7QX5WGwohvJWwwLG2M6NWHBGti5EFoEMvpwghx
M+1MscrlVOvunf18w/wj189HdgPWOfxDNBYnMBa2sFZrE/mWecCFhFNGUDyFi/gA/MFm+Hnr+ch7
sYvgZ54Wv+unGMDbuXWL/7wrhzlwPspZgG4JTfIlxFsWum5NwcXP9Q+dYBJW86lxLwaV8nh051O8
uTFsmfBdd9aDkUeDjbISOAFuTG5quDdNMzOpB1jTpWHs+9ui2KlSe2PtLwhbMsyKt4V1yD4qplTN
0NkZvNcx9qGqtNCdBOVSkGSvIyzG01+b0Om1nV28vvWNnuFQ8mE8DGORwleclnb8Z0bECtu8g1J+
cJJmB/n2w/5gIXNWt0BVZDoZZlGs8Y8GcaRvyviLtSCksTcKsQGZUNNT9JzWc6FLP3hUvQDo6AoG
U5CwiZLRjW8acFO0dedPvFDpGpKsnk2gJKrnBw6DUYDhEETecYfCPzfFg6WUVqVozCXONsnRzeEb
pl/mWD7HYgDIb2Alm7hT9PIodIDsuFu81zQkYob3gdDDbb7Q1bYD3D7B1JsABxxCI1QpwmssSuYt
efDvDiwwAd7qAyaSw4y5XR0US7FSw2xqg2TAEKKUI5KIkmthGHJE+8eTv6ax0R0eC45W1FjlDPtV
+Qj0/+8Qh7EfS2wIPn5KK6oAwYQp/pfJALeHAl6tLu4bUNcebxbQVHKLnJnjsZ5yz8pNLJadLacI
PakU8UPjVohdlZ57Dx75muUpqVNSxz05Sk9iYw9+qKUNi02sYJk9f4Bv8RbZ0nyZkZ+ILhiRBjDJ
76t2hdnMJY6y4gv6Hws+gqG69ZOT5orcqQ6yzu/T5s582MsO1jgG6I1ZYU5Ue+T4A57bQXeN2Wx2
84g9LjONmXBAkR8Ve0SeNBKC7DuQkfuL+WLtCaYyXePa0fsnixzlHRkawZI6qYKok9zF5kqhU7Al
hA6N7LfAzGkv3D0MSKtaQ/V2avTb8ecqIDO5KQOjoQ5GollArhdzSsHyfOLayY3vnD2kYSfBmRE2
XFea0kQuAiGCGLevvakX52jWZSgBI9rUlAQEwK/FQwnPGhwD2oOpPQMoqmxA++DmUxYQdSNMd5ea
xNlYEaLKMsTIpA0raKl5FwCXOD88KlC4KtmBdQx+e4V80bSxEeMj4FU3VqQt1LW5znrpBMmdhDqT
tFndZSdiz3TpURKAbykiYMu9vSJ1xhiqqPUsJqiT1m7ez+hUvP6q310KmHuAyaKcYIKKQB+WRNCR
Hfs/YV2fhUPICBrPtiZqEFhDyW6QeznDXbJL4eupvUPNnDemvVlxlakVaqBefr2eD84grI7P85DT
0vwfM/JoW1/6bz2w3Or9iR5cQ+9p3t+jd12TJzkLZg82kBDLYYFIQgYgcMPORm0lKsGnqQjVsJqv
ec3EGNQjaShinN+2xwwwah4D0jvpgWqP54r8EwV3c7pY+7oHeB3aV6mbjUJUYZ+K07oI+SO6/lys
nqpdMh5BK01mjxS6pTLlXfy/y91ChYsRHkX53xkO1DXcCD9yJPDs/GJDW1rGaxsupeSY+K6XsM28
77xFysZjP4pt3k9tfqYN/L9t+a4qG1ChUvi7NcOe6VHcxlaS9l60+XsaZc0aqo1DcezYWP+aEiLw
xY0efub15c5eE5c9XwMa5Hb568Tmv5iyaj6WmzADRU9mTu5jrK/Yt6NM2dL+t3UxWsUcLnzD5vMJ
60X53n9KkHgNkbFWyryODejPXT7TPhOzXqQPWp6alFG43zM6oJCW0qu+BdZTjJe+h9I/GMuaabNq
0tTC3zoCpwsNtdYBUpo8AnP4MLEdVhT6N21N3gxoiGL8PprtB5b8kY5Xk7ODRkkqJ4qlmnv2Yr/A
1xKv+CkHdv4vN2ijzLpJaEejAM+ChADXcnsjXlrc22UcJERC2qimaOTPBr0PHKjGGHq0up9SqdvZ
ZcElPE5VxeHPZt0Gw/rKhPYXFLAkvNBFJO/OrEA+jYgunN646uTeAIw42ymcA1NQ/pPAS1sDHJCi
erubRG2i4c6W5hkM4zCqZ/Y1w2ukazZB8u7CNs++gK/iAZoEeVMCEgWYauegpW0hoMNequ2PXHpb
HzD18WbMOf+zsJvEgNOtEo2g407yWHGkCPV/wjK0qDD9SW1nIOlC/kIOAy6IxlAgi3u+u5oLusZF
EqBCuxYCqiivLSIzOWnN8DxP92c2H5DYVXYmapJSqQMAmzbu7yDtwOJyohkq4uWNrkUVzXP2XRi+
RHqoQQz38sLMDntGHHlV14SfhJMRyOWDq9uNWtOf7gucnO04YK8nBFz1Ab5lIqUUu4iUVOEWF53q
gSV/Rs4Py3mK75oVw93luaJiPvQv+G9xntTdheldB6W0lHS/1icOrLlceqSihVY1nFiLbrx4wLUn
O/Mqxgr/eS2VINCMR1V1qtwQyiBY6zLlueNk0ITvqBosRo6ornluZQo0i6ctd7gl5uu67nP8zKJp
PQPp6oooQqcdH/Vsxe5Aqt4TC4n/v03kNi7dLdsGtpSCf506Ds7/w3Xo3BAbZFjpoNPIeTnbGdIF
XXbj5IZAdL3M97dINxoHX0Am0RMUjZP57bwbrNN6KacxUuGYU056UId5zBSQHYRP0RDjdHfOUe1P
Ah8g+xKdv7tr24bRYV9Ei4Nc5dl/FGR9YJWRof8LQzGjkc1qu2f8SYf8vVGb1s3tY+AcbUaCFyA2
ZPqeEmBJc98oQEPizhcZnPwtK2kbCvqRU2LMtSJC2IULpf3Tnbmg/+MSnAlwl7WX8OR68pepydmC
+1w/Tt8+N1xPsovOcLOcjgEVuSDYb4O9X0ZJo6tdcHH0MlyI8AXqTLKv83h0DNbhqBewDlPmh1ca
FMelYbLsW+KBVzroL5x0X1ivU2P2CPLPrn3bFCfnpJ6qmcer9OwJg4bNT/m4Hq7WLalszytR0UlK
qHqOfYkBE9KdkZ30O5WojDpnuQnMOVWGPK+mMBA+6CpJh+HEzlQDu4GJkL/sT55L76T4G3qPnBaC
bJbZYEBR9dpmjCvlt74/hnYx2ZaHMaT7njMqeHqcYnVpQYySker2PmaZp1vjmUershL8LM3+bQeb
9m/m+tP4IT2K2axtpgl11k6ficO7ZnkIOVVYd25m5qlhKeKsThR6u3d3KpIcduHnfBi1j24DBKBT
A7BUhGlf2fOxkRpWHEicvS4QT0tKQVzGaJZOUwsU2+cXLUqDeuR5eGZgv2/+cSTJUcYfpA30kAsD
82Y2s/1WBtLc1ZMtVbtvZdWwTjlM5XZmL11HFK4sKjqnOkCIzRSidZNhutEJMF+QmiNGq1reItm+
b0oSO+jhLsHLvj8WeoJAy1nSqtBw3I3yh/3ZVSNdxlvPXER/jzAqvDwXrNXRmHUlU6ACy2j7Pcl8
d3X9+1rkzZKq/SZQVcu0anLOSu+vVdSxpw1uWiO904G1XRBAwmNxzfV+twplLhEqZlskJMGlm1yu
S8Z0woeC24xbq2SvbKJwNx3+9h/6GPOjSfiHFdQ6v1OyXeFeZTM1cZr9g8Ua6kR1FHPxhzJhTYfT
rMQTjZrYdGuN1fEfPif8iM1yqcmnG1PfKNCr/aB2wOYj9ICEa/xnNoU3+MNrwx18CX1Gi9oNlBtr
Gj2eZhfqhQiJUUsLAf/s3eMrbwpbzaZ5zaXn3yBSfVZbLQNFWPwtXoBJAGxKv6V/LrwuzO8aDSht
hH+QMwg1rvm7z5jnN2HShB5P11Ue/6dhoHoIHzt5msKUdukjOhgb+TwiZM76ZTjXRzP/fclYgXFB
5WlsY5jo4KQg7UhxN43lBgaG1xmYBVLLjO/vutGIZZ//hvO8U0K6y7JBxtQw7mjBzS4YmLK2qjjZ
zsVEEp7oG9CSH1FXxcw/vo2v+1kroE1g/+oTlNDULoQ+38N8O0oaF+84Hv64C3YBNxmjN7J2Nf3Z
45QJwbtDVSvtnX8x9KBKfghyLNlFdlESZId6afYnvzC9nkca82pYYFiWo8WGBbhnRIDzXvEqIAAg
ZjSpQe67VHBPMDq4wQAuLT4ZoMfnLiEPQwknL4Ik3XXGiiCqBsa5g4O+ZkaE5q6qSWQuljLuCJAR
XyXN+R+8ZNHuZmMSYArBgxFmk3JyySfFKiLAmGR5Lh4jJ0h4MIyEyjpbDf8h+bYO5emRH/OyG8N2
IPzBgPJVvtzn/EzTJ5XWLBGD4nfjZfyIpu3Q7pSydEsPVnHqeVhhYzxIOd6VqNrNTxTYlkQANGxm
ov+UyXfQivWf1P108iHYbwyDZ1mYc7/9r4r8wk8nKnr/QQDzyXsfeqf2YLz0nLv45c1ZK8wVJ/5G
rXoystGNTxLUvf264ftBTMH/M+r/7PgMRZiEuMJ6FhKFJn1G0WJytYcmmX/76X7bVjCipsht7TK0
UxxUpnJUGoPl7RXTPwIRSrh13KgHb2qxpGeoJPt7SUHjOFnzfKwu/D59oxobpzHPu0leTuO5B4jl
RLLV2YPEvk7/u0a6aCQg/dBJizCgK/RrvXEljKN9LaZvZEuE2Eo5brzI2KrFvM/7hTa2C3tXQ88y
U7e6uH8Wk9U5gOpnqNw1Ov9AbH54HkV+vsc4R974Ho2ImZtTZE5azwNZJd4VxrSp8Y2PzPFryuSn
kfUWhXbA6thdThacibfE/JzblXh1q5Zn+aziVi4nfxZlLgCICpPIMO/JFGZn3KxC96HYuFIyZ6i3
UAYC9LTmE2BXMIBCtShGE6lKrA1/Y+qC66aWyWLMc8YMlvAhEbNNkSf+CnG8td6fOn9qaKiimdsw
TRA+8ogTgqSzKibIhyixLOwAIdfkMHTEOYUKVhzpsEK3AoYTeFZuvjcyQme4ENWk4OSh0f4Quhuj
lx63BwqPp1e+0M2qz7+cN0Pl6Za0eyjGdW5tNdI2K8aGxv6tt+YLNEWzShypxnuEefle0EqjdCIa
YIDH04IkufC3DTeoAwlTDTNEY1Kl+3cgRXLH5s/CXvRRYLvbOaTFbC5JGvrGOUh9W7enJrAe8a2G
tMY1ALiRHypOGAEQ/UCmk2AmgATEhRDqX0Zk/qK2nlC7iNvW2uKWZZWJrbrI3PFw5Psw0KXxpyMw
iVgIEgGW7ZtL1ZnC2V5oxyxmDE4LkBPW/oLgXauldwFfzWfEyIVjiaUH1KZjOdC5K18DTgWvBbtU
t0JOfVWYG1pcCPVZ/gqKOazm9GwxL/AtA7DMWjq/2mWJDr5HqCouKlAZDgSSySMLzrwUGy7j3/SN
kQqTSo3+kVTE1YjkGv9/1XEdioqXLp+oN86M8Sl3Y6BXSnV9IICmVF0rw6hhKL3E2d+drbg+OcqV
2vdG1ETjn16tTus44JfakkAsDrF5E8N0dwyREDPUq9W1nATmJpNykhlU1tZ/KCUrw+uKNMya4vP7
E+5i7ZW286aHPyqOD50HXroi7U+T58GihaO/20ovVQI3ycI8GzhhWQOjbEPGoqoIboZshi0BwRL8
bhqsG9vgSL/aNy0v3SCGrpJlabXv0ZBN/us7auCEHKKdGJTEctgHbfUplWRbe8G5ao3Olbs9eq2p
GDJwKU0ioj7m3/prK7HCgvKw30VO2Cm7ESQ41trm+DBlsgCYnpnmRpPUGM3e74aPWnGTP41E4y79
dqhcrbqzSWBzYzUhLNq6lYF4z1xQLa3toqKSbN9HwiQI6dnqCtpPk3sMV0BvrBBRzI2FNkwYy7jf
fqCxwS/N2c4FZlJWAIlsO3pHAPJuBr6fsM5AeOZ3uGkeffi4IWRKIkdcNdRZMFUIyOJVeePFlgbi
JujsziPDNbJdzQjJagInDM9PPxubq+R6VA1LB7DTHyQiFt5a+xW6+0P9DRPVtkdXojisrXQyvo/f
kQ+vWF/d1zKOLZNV7hWjm5IBRZg+weHwPZKtzXpnWJCoxDvErnMd/p2kYYZYo3W5Z0c7keY9J1zS
6boLNb9bH4x5VklIEVesX5BDz97seMOcfB2EteZ5qZbqXwSahUCWOczUjtpuLIK1ht3fJ/X+CvVE
PmwWe0aLoRlQ8fvTZlfiLk6IKEgky0om42xlxsurQNdr0KHKcHvvFiqD6itAsWkNPFfECYOLjLyg
EGlJaXTzDn9ZgJu5ylnRjS/Rynds6dLrTJtjv6frheUrDxTtsoVZ7toer9CYFXuwHFaDTALAhV6E
9tvNHnb8nLOnxUIa8qak5fO25yguStlkKk7X8Orhp8yRyZLc9zYFRZBRZ/ixFXpQnEl1tWtxnivW
bA8lUE3Epin70a/vNHNaULrRuDSRhpPA3lnwVjlU4CktjOH2sSwkjWAgYNMcNsnmgTYu0au1dxfv
p2+EoQ2UoLi552fHaQx+5/6OVGX5xADaexYPXkEc0fXZpEpzwCdaOf/Cz/6JC0Ug60qTpPObtB4w
dMFP/+YrYKdYVQKcdappan2x61YbCu9MwfqtH5YZUo7AeQtDrHscW6akE0CMSXZmbzmuW/bQBPPq
xk7yHKFFzNSro6UNPqZpWtCWtZDqhankVnQL/koLumqtYF8x51hn0qXca0iU6Vkspi7ktIbUf5FK
AC05OaOTf28zf++4VUuvqNsr9wbYQIUVXAwSjZpd135yVzZ7BPiaT+9NNlLeskuxiBhK7IF7VHLM
t1UFT4JXpfMM6bR8bK/Gdj5QQaBzJx1/N73AjUxnZOQRJzDj2Dce5vdr/fnSQou47XOMSqdbUEzp
8wRJabVMP8VA1//Twy8K3ywSolLtZV50HFlAo7pqoLO2vP1Z4rDlPBqTungTgbzWIN0CFEsDaOhE
K8GwTgSsYZNfcuGjtgvLwi75tOj/4FffUNqSoPAlOIjMZ0Uxj/4xCfjIkj3XBqp+clpqNQm/Jm0U
VIcWVkVuT/6CZnjM5XDKfef1E/yobkSP4UBJyvF/ycbcWQZ3AbDVqtLS0OI+z8M6r641XwzfqDD3
AMrMtQmkwGNR4G8tuZ6udqE/zhlBpb7OExULmzwiVnDB0hWUZT7smj/8Z8cMH1hvcK7/YpU+O/M0
mE37E+6HPiwGvbqOcmV6b8K+lRNQRPIuhuF6wt7eKFwNsR9RWqdR87vhZpPPeoo9yxGKvHBIPIjV
Vm+u9pUuFU2t8K+jP3ZPwuxGiYRcE0D/HvPuP0iYGuTVwGCtl9qJQTt7G+wdpdPmi8YW09Q+0w84
oegF7Xe804y9HFzrA3Z5NOc434pzrRCjHg2Sa6d7AEJKYWxkbqII81g+m3Wca857oypNr0aP+agT
AC4u0lgmoTPqlEKUMsEt4boDR+7+ip3NaJFaoeakd558UBr2ZjjT7WhfGyqZFeTcrx5QKxSVlYOW
HV8PEBjfH1z/5pOWaYnWcwawaAIrZf8LklH7APJRRs5gfexrwa8hftYIyD8pJ8faFvO7amxyYBPA
u3eNT61Af52inXcbUkJW4U2ziDXLCakW63HFC3w4kq5GChrbpvac3l8GG8AEgMFW6YFBTUyUDpTe
ryjUYyCFb5X6BGGTpdb240JBu4mJGeHG5UP1Ruo6a8VNXsat7r5bPRi3u0I6x3W6iVQkVk0Jpm81
+c0kDYnaAgE33zNleqplZ8OxmMPrm06p/kKKgr8IiJIVgjAtywklP6MiqYK6xZu+SSOiyLLJtOYA
nIL46HrT3VCF8QdSHTizi0lwdY9L+xEyF3tGNo2rJWB7N8AEDXKSuL9KWVIXpXCdblb3Pe58FUeS
aLaihuWVckvInm7fPZzjd09+BrmgxkxhvqBcRlfIBgTQTKwveWI8QIfw4kc03rt6SFTwq2kkn3hW
gyhXAJahfspd7eG8ZQsDOQnrptfcU2KxWj/UAcvDJl6Nc0e4Q+FKNjtcnpjmKWz3oa60RHtTRPOm
wx7rH/Ea9eliVZzBfKfzOg2+90BpR+OF7R6AghHCu2QWZ4JTv46ZinziAaRGFTCvJ5yONxDvhASa
8I2A45WcVVvaWM6pNsHe6K/QVB6zTvR/k79aG6Ua3WOWYPPBXZ8ileh//wTKh7vEEB+g2Torlkch
Pn2+YRuy5AE9T44w7nIiboE61rca2VU9bfRR7h9H8nYq4ox96/ZoLHAaTzYFPQkekSZ5Jfhy3L+f
b/8KqsgJx3DAcMVkA+1pYXH5zAVWKbU7KaZ4YM6jtRIPb1aaq4VFkdzdXiJkuRlZupd7vEgASpUz
J3+LywOWF6BruXPQa0xHMV2fSR6pEdBRRS/btt5z1LiM4jeAgjxuvSXhygiVonZnyNqDuTlRKde5
Ceftcpxhq4xSuKgh0ffjuAoZdE4dc1+g7S0mJARIcwUEEJxMi7kOK3zuIYBlH5OCoGUnRkIrDXr/
JxD/sF5IO0HNOtE1XD3afDSN7uvuJtg5rto8L4dX5o6xs/LLBeu9iFZbwc+uq/VgGI+6b/XCl0dj
N1WOMMrXYIIbqYHQwIQRYudnp3bBTAdnnNypqsqEKtKQd1sH5VB4jh8wqRWncQa0HcCvHgOyNZjo
SKdHj8AlqQ4auLp3tQ2qaiZY19j75uYNOhxBlcvQ4S1Q5yLESunBl+m/6JDqtYDWpbz3m7g29DxV
aKtgzl1082kw2z2KLefMaAji212yQ7l8d5spEriTlzj/m6ObCNkOY4Yr6PM66/cn8U6HJm/jgwhu
c5g82caEBSbL8CXfKOH2QsVU1pYsmc8LrJ3IZO8ES6r+LTSHkyMUDcYFGBT3FdOFd2gLaSz84QVL
1LF1X6Uwt0mKYTVFCoS32YqgRe5HXNY4wS4YRqJyrtKlW9CD4CkXuakiTmIOgvzzn3axz4J2jkQd
na7b3N2cQSwJ2Y2ngeM+1mBdNcjFhmGX+2xbzLHiDxiNfmgLEDSh69zqxGLJUU1S3lTX/moz0j3x
CQq8nMMBKDSg352Qfb1ZygUxVXYiR70Sil3wVrGL1YKpMRL9PcINOjvHfEnC4X4JmlY/MaXNaRfk
uatB24HKx3a/gYYowGbzfT2psvyQKNBpf1bwIaNTdUQW6FYWtXuPKJhV8H0BFGVfZAk67utbc+J7
+YEywJBM50Uwat5xM9gkubOI93EqU9r1O34q6nSkWSGlFy7irMnkdLAxPOwHsofwl7VEiYUjmzJg
w05H4gt6fo4bYISyHV+QB1TKCQc6gIBUhPtSv8V13++06m80iJC4Af0riNnpEKldSR29BrrGTNzI
w/0pJ89vGonNxtF5uknDEJK4Aobbv7TlirgBP/vXu702JEr4/Y2chcDrSt90tT1zpbLomtr6v7Av
7/o/JiJD1DFSu7FQMBb+ngtAdqr/0EJJHTs4nmFZ9KfZqA/nxuxhF/noe7SbeD8Cs784i0s3ZsoQ
ZqtRQK1CMhE1C4VZOcI1TWMwFLZvxdoV1C/bbu1rsRStZZmA9nvrTRii3LbFAPBNzKrorqBEPR5S
qsLix473MGKtHIa8kHZIjF7FWi18FNVEgm8BGE7D/oJZJNk9g+g6MXPVLDHLt9guL/Q7psiA6BI+
YTolreJxrN3nsCXm8ncQWiuOQPWt802OS15LGgjCzUE0xyNr7bTkFF2zyUxwN2Y+fnp4oo/178WO
8N0EP0tiVb7GWoYT2aDapYHHAuLMWQO+DVHbFo5RzL/E0GMuV2yMzA3iNKC/++fKtlyBbciLxx0W
dSU0xHgbOHCdw3Vcl/qnAVcrdLY0Twti9eHIrVQC2Tks2iQZzycMtsEbYK7Q7sCDdi8w7iuhtZHG
TpvwDfm/qcYs58YoZnct2PKziAoYyHTsfvtFeOPgxe9UHSHRCyvzqOjG8yNA3DSWb84jFBDj6C53
GP0v1E86bhCIBJnrW6g15gfs8q/Y+wod8aiqha4ARukWA54m6wJp9MSkOAhwsA5uw2dEBvfp1nYs
dEyzofgrEHh+lUTJD27mxa7AVZxd1Wt1IkO+DcWYTIVgLzaNQc5GvCBxaMSmoNaLpSpOY0EXf3Nl
5egURfm8USEoHw7YC7Fw6mdAKvE31ugdyQBIqZLQDkYLGDPb2i2g4CVPq6uM15k0pgHsEpHN2FVB
hPjm2KcOtyDUo9RTb+8NeUywPv+Yj0i6CheaT5UCrBRXF1YKXMGR8tz8622eo9V8Nkbvs7ypMHSK
OUYYpuzxyEVvtFwXlYu4MUzMSXcis7HmvGg86Ryu/y4PfsmAqlY8FYPjd6Dn3ACYv5rkwacbOCKB
RP4hvxwcVs6PxhaSyvj9RZKyGXr3XRhhX2g2omUBtkyl5aeE/LAExXJB0+wKvehfyU5NFQbJuLc8
csJI5w6fQ/R1K6usk85Wmrjx5wHQaEE67F9PIfiGSsp/HQmQCJd0yr0Q0aOjDI8JmgjtBXQlrZBz
Sv70y0ADaHYBRd6e9ZOBVXZbSQCUl+u83bEeb99Wv5s2UxxhDbIqig6GKdPXNwaQCdktoiCOZm1e
+hBbn9ePWux//TcJdpQ4UmY2xMYWHqIeTx1X4biTMW0By6/1zMAN1sBMvo65AaHHkluK4NjadvmF
bHLTK/Qbx4EVa8Wo11HY448gE2VJS6t2jLL25hVko4r/rD6ArmwxgdOZe5YX09a4Le6hCXkGIOow
7QfM7whG5ivlCt6cHwBO/JQKL2PYIm769IvBjbRUv+Y64mZEbcM5tw1EteM+9L9QHWGdFMZgd8TX
k6KOdHOhRsAgCAwdHH9SuCB1dpht23kKYdB5pklmIOmBdrWLal94QMz+Ovi/EMdu8Jj2NCLpFDdR
MdY1lwI8B+yLur51OFUYN+6VHAywWCD0QwvWUsYjrwP0dN62k6DAaNH/xvR1lqSXcDJ40mKidlQj
2+6LZkaAxOnjBMQam6jV3ao3nelxHB91lSnm6zqNRydn2Bv0ifxKc6++0wX6C/26iSznO5gISYX3
lHThmsHYUNq05dW0owkzEbhHoBlBIZyjqfNTPoiHCGOYbbmWSVwhJRYklVj4ytfbiVmG2f5v4EAu
w8di8/wJ+T9v+S/YGOEHi4PdaTgN7j481MR5IIkBf2xqqqDSLq4yv5mFeHXNeS0xBMOr1RmPd19u
bzte/WaTGlC+quvvmQ9Fj2F4QmdYzdZDXXHDzamMBQREeoUSORVNf/D6qjbW0Ru1K9hJA83i7vL+
gPftZZhJE9Xa5GqNsV4sXM2IO3DpGXK+Coyyxo3LRRhKMp1xnm/UzC7w/0gZCKqoAQq6Q0qbWoOD
O12z3XWoAnxjWvHRSSupH0RLBrBkn8dqZBMUc1jjFt3DD1joeQfIj7MCecpRCHOXf0tFsxuuR6+W
CxW4Uo+SnCtidEFSZNShDNwNXA8h81WcHUvtv/6ks6bVuHWH70Ach9/53tR5dyvidZ1f4//rU5PS
3KLpLhFalrxSOySZTl3D0+k9Ici/1hIjLQARNX53Ne2oZZqPZ9rggCp4AaUTSgJEixFV6CONg/PK
/bBG77hwuNwcMn9RBu72hZUMuHaHKv9CSG1wpM0pRWxafshSE+yvA3Ia/Eobu0zHT0iR9g6WjqH/
a5lAGhviaUNydvyuGFwIR90mAuC2wgE+8rLSIcPSnX+WvAy4/wP4SCyZZlK1Y3nI+3sFzukJblWB
A4ENd2s9wEb5yYTrXmZ9PGsAz3KBOEJfIuoMQJRyQEvgPe61kN5Clg+C5RLcRPDjtBQUYDdVB2SB
GsqqMzm1EJtJ3b/MrEHBprRa52fkgAxRdUDHoNzVjnH06H5wNQtQ4Kiu/xJ8H++Oi6RRgtheeDWz
gQR6zblw77zGbbzVYnSYupD+MWXXX9Rm+Ke3MyV4KW1EV4JpZN3fYl2HmETyG8k4a9jQyzv5T15j
gnG+d+kE5Vho3/iLtDC+lAnIMfKEDEvq7g8YzDMMeSvtJu8Ru2hqSf5ku8m4TDH30ghH12WrjniR
l2xIH1L4UVa/DWsJHFPcW0ZiT8ShQRzMwyZe6x3RsX23RwGBXT5elR1EpkQ6A4ijRfIkzELCEPc1
5I0r0esd4x5kXdhHigE1rjhmSgIvMfw0KvXrI7qdSXnSB6TKeOfRkdAgAdvA4lKAboP6Qul4//Ni
IqGssFz7Cx3CIg3akc1uE4g/ict3nqBXO65X+eAP8bi1BH3USqm3e7Fm2fC3LjgthNu7eEGPmRDF
Ry9KchTPBc5SDdHakOYb9BHP2+TDiA/VjaOVQDGlNrQupHuPR+V7v15GxIayFUCE5U0wqERGXwM6
3nE7h1lZJpwJgT5IRuYOErSo1X4fNQO+quAkO3IBa4lhrxGkfYEL5XJp20XxnWksMDL+3nRxc6Zt
P91avsF97K9WQ+HUQdlgEnit0DLaK/5uXj3Q/Kg/HtVZj4U9rnLP9UWynTpk6cuK/yS12W1gRJ4h
c6aBAHMn9iqIyXxDSiDEplJFLvdVHfofk/6enxjJGuQFDEAfbUa9HV2TpCVqtFc19e3pX96V3WNJ
FdFnSt5ae/vTGqc1oWvVmheNlbVZev0R6UXXguPMDCGQ4cpWFuaaWG7f9kzKLEop9D6ijnCwmmv5
XqMHFH0oFZMnkEwoEhx+r3L3o/THQOMUS92Q4FfqEMGnWHDG8LkLyaakVMEdIwZip68mzZM7Dwu7
EXgRRO++hkFgfNSku2qofGnIfCiho2VOWkS2IffmFVjKS76h+ZrS67mbJ6SkY0VvyczLb9lFlanL
mQBIA2LlYvVjZjejwocLgrWeR5tcdca1sMjx9LD3MhFHFYu2quvjC75GY7wG1G1SAJPx9N4LK/zC
kMYAdB8aK1iw2HQfwKDQL0g3A9OxnvaeCedcm/qM+YQXD+3Y9UoddIyDr5w8ZVGLOGWoyp/jXoTG
uycxvDWJiXWXfwW6ahoBNY5XG1kEgDmWhiWy7z/ZfwRsAAh1Ph7e8yBo6b1kxEacff2ghXG8YyDN
59NZMFJsji90Mq4m/xnscrfC2OYfqdFFHFzMUlmJiKiodvfW/jmGp3pM6iTV4+8e5JYfWyu5OyCv
Y+FBPrTnSK0z1UpyFvawgYeu+Er/t2tQe8nGWhZM+mUhtLrywpQmWHyJAMPiNTaI0iDafTW7Vht+
2Kqoie+Em8dnUZV0mYpis9fYpBdg4fEqqSpeAUSQMsaVjkU15n3ubpf1pk1cMlUGb2E+M4TKPEGF
Bag7j6pD2ARH+EhokP2fNZgwpp1JjG7DMMrmAi850c1E0CqMcgvVAvkds5rFjytEYbxbwIVMHJgb
twG8DOmFGRFcdz7rUeNCg5+Ck0Jr1gOYc4sEM2Wazo/8alHQCYaU4utyUSMxanCdbkfUAMvlugMs
wUCT2bFSep0wLMo2byOzwE7tF5hozI20Y0c/ec+aqq2yphHkh/RPrBAjRWxYAuuEsBEw3ZZiuC2/
GbO16fC/NfvtheAgCbdjIESaGHtI5ZV4WUuAklI351xvsQcAuW3xCFuLR7Ju5hh1cdsIWkDlAq+Y
rUzTMuybtPrNY+SHx3uusCc7owY8Jxc1XhRg9jukW8/8YR1xNqSqD7AzGDJ0CN9eyESTww2Q+oPA
tkN4B3CW8cVyAIvh6+d5cT0YGV4iaslFeeKjl3VTzsUCceRGzKm3RKqOruS0PyUCqWCq892SI2ov
BOFj5cVvl8iSbUCTCjw1HgprLTt1cocuoq9oOfGNttyukqNyg4376hlJSOdWXFp23z7/TN9tNeHH
bSX12MDr6HzYsC/TRMWSCeAzmBnXxDrhT0RoR6FJfob8KQfydm/PWl+gssOJa8sJYAtedR8rrzYF
NpkyNIX9FZn7LKOJCq2wnMfIG0mGEpPf3uWAcAUbGo2GitYlDleEKiT3AanglpSzn+a0lpQe5uzi
JdQ+GjpN0xkAWiHGj4XmSDjIph3JE+6joMkP9LDjAd4ScKQGtiH46jcH++hy/AAI/q+SHTf3wu2d
InOLv6O+Lm0Gjtia9zWO5HPuWWQY5UDG2k5UM6LK9fdXRUec+D9pptCi3FHGuUvnPmZ0pDvZsBbF
7fDDbHPzK2GMXH3a8fAnlZWzR08sA+9J9k/c/H2eGbhs+SDgrCVgTDQefFEJxJOyWAAJJwkFLyhd
yLLzH5o92UYssFzUILSXvDFD5lVWQ6h6JllilpyLQoSF3oAsh9ONxqc42ZbcL4A3XEqfFxcTJ51I
wxk0ZuqKQyGr8zkCAvWgxC/+PKAuMldz6cIBpTTRjrQqkeORuIua3nBfQ2r+OQqNQJOvUx+9PpuD
ACt27KF/eAyMBJtwymaYKDBo00FZuWC2td/ouUkGX70qjvQPfYt27Siwh7Hk82c74+tbL6LqkzJS
dTCVSpRh4YZdkJOrQ+IDuY5ETcoH8BvzimX+79cWj4f5oGov6K4RJQTyMvyD1Pu9jQutOIZkXR9i
d2WRTPI4gnGRqhydoGfA3sbyVqxzYdrRCa8gVRimkBZQVmj6iqFm9xDv8eR56P5cWHWzqjrfhN7Q
5rxiYEC/s/XPWmK6YCadaGoyyHiIpp/EUujo6xDpy/sAM0Rs8j42DwaCnJeKw1V3lZQHmWfi+Ms8
Cez8n8m7fozTojQ1/qDObhLX5+Rv4mMr0P9fjUUCePVHVg8oyhBKZmUHzy+000IojGVScJirqKGI
+3a4ZGWH4rEaC4nYBegYVDUeSQ8ZQA8w/Lco3EawoGsvRF/E7Mwoxi31AD1z5qcdFNumILnhVTjr
VOw0Cw5S73cBAXQg9MSt925/+ny0wu4RpwyAChcb/Mr/5sBwTpvyuWq8oQA169V9KImwY0CZFKyh
DgF49JU/aXUy4fiKrEI0G1T2QNN61qK188b7U3d59aQfcrUWutgdQ69AXBzP0VAqK1BlacI3uFI8
eVBvMoHZQB6pq5O4k9uo4g4aTMJf8gjn099JulxvfsijiaFqO5Y08VWrWmtOXhdSND140uUhemjQ
xZmeiUAxosaxNP1O/hXr+UyszmR6230dNL/4ZIdNt5Eud1KK8mevUrtLHdhDhTqMZopCScUICUcB
m7UqwVM+ATvws3pxgGsYS+KAyhRVIV+fzjQf/XkfRNpuSGJGjBmj3LP0rtxHaDNm0Eezxqmx/2uT
9Ab8STpdfj4y38HpATRcBpj272ypll0oY8QjXVcaGSp/c7hsP5nIRYwOytnJF+mBvAUXLdI6pn59
ayjKGZTPGig3TkCbp2rUA3fW//BRXq9XjxBWleFfOGKJm2++byKOdLV3o3oKaQfYdwe3UZ3XkxmM
j2r1JcX/PuZy+emPWaqbD6Nfr4q3YJD7ktZJ8rfeOdwA8F5Ih+Nv2J8451x2C/y1RmPBfEWCUq0U
8VtduaysD3a7K7j3YwMWxnQT/RmVh3tyge9pp0hBLMwVYM6kn6XSBDowua2PzyhVEhPYeP9+IW4Z
IKjcEVNI0NEPQG6yctTFe/CpeeXTGAvK++TcsUfTEXCyyjEzWu3uZsC+AlxnXFKGIzg3GWHOVGY0
yGoUJsbZyQpoKaidHF13tpnlofRBJ5uEBqTFXRqmP5G+gEW22//dfSLZo6rL/Ho1ATx/WRTz81si
YJWFSlf6GgwY0tMbKh7bmGtOuPXUq/KJSOWUAkHKw+budbXcaQpR55YrYSZdov44BsCfas6bcl9j
71cDmqzb7K9uQISKmZRV4O5Gwm2r6funS9B1yaRihwxJtNTwtoLSzSVi6wKaAt28sKB+vxxRgRdx
NXZ6h3QKzsbu6wwsQcQumSCTb/y1cnAfYcj3OqcNXacA3hWP9NLt9FcsVnMuO9BpJ7pF0L3QlSUX
D1tkp9HXzHoy1lbGZxVrrvK/t4W0DqxVPg==
`pragma protect end_protected
