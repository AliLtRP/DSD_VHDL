// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:21 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
QvWbhhruYcvg/8ZJ7tqcY8adylqOaytswJpSuCga6pUuBlj/jJguaIGt8nLBZ7fe
lvZW0/OFLJg7+EiLEWX7e9eyR2AkHkPxFAXLvmLyVRFPSvsdMljkMC4K2v6obrne
JhgbQbtK6gSCKABotw+ZH9MUwaV7ZA1kJKDTOXn+HLU=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 29664)
Y2NdHyVzWAd4g0rFMx1+4lDOXvnedI1sfYUZ/LEclfNJHdr6tsNuazeqVtvkg+Vb
7CjE4qrPljXB9u8H1D2iSPm9w/7PoyW9oDnvOxXobcbsh20c7Nrw/6fEp31QmJD4
zD2TOajeORnAr3JtoP39TnGgYBhOGj4tUAFzK2leyBmNnbnXgmE3U1IElw9CCPOD
y9LBWCEWG8iLQ9lqhaUBs8V1BdRZDG7JzLVlHyBoQlqIBLJBf4RMrp6thWyI/ywn
eBigL6aziRqN6FfgJnhZ9Oq/VsrYmXyzsGuecuW7OVv6jLYab4cZQsDyy0A6nlFT
0tFiMDmcnb/yWrXtweLfZjtIgYX+kk8UQyMvNepaxh8EUohyK2tlMeqBadU5xdUH
WctqobsOHvaGQt7lFHLrC83sFjdzZLMpMtcgBKCDaHxGMI5s5VerjiDy4Rxr5UDJ
6MaLTadvOtPyVLfnvL6NErAnv1O7Tupfn/KzzPDPnPVmclfy3WMUpJ2xg2d58Mk2
dfBI50M//XfCKAhBCURZ9x6wsA2sM5WaEgmpc1vL4bul+oMorjI9hkeKd5anesTd
yfcJu1I5fVrchwUu8xPfP+A1lMAf6r+kkKYcTqv/P9jyhaUCElNpv2KIjkBpKlhL
ePj29qSU+o+5E8aJq6u2Zvi2FDyX7UXq4m/zatri4FkU6aP4eWmHCYImSutUKrdI
0QUrAmcgKmzTtUJaKzCW4KyPjDtwMjyFa47GqjCecnuRjt4xrUXy6DeJMMIpjLPH
SHVA4NswX8VKDttqGc7FM60LdhVlJXRgn6CFZrDk9ufKigIivqU/709jHgYTV8S1
yGwiv8QBIAQ8+JPciqVDDRhOHNWSWmc4d/KuwMnnydbs+AzUNtt007dO8sCYv453
Va1KF0QF2Yk657/ZVFhWmhlACkKB3SqnJRDrGxYtBU08Yd2whyj0dy9+ydrQHlSu
PP+5H/VUIGCCKMZUa2PaI6JeWyu7US243tHUA7XJqubdEDjuM5/12jpFTPcAeqUC
VjIH0sc76r/cidQbrtcMkcGF5g2w3CZx2bys5wWKo1Teb3yZLxe5Y56tW6GjcF6U
ycUsr5kPDdYmMZMm2MkbZsrV4KF1TdAdKR5I27SP8SmmHuXGKPkic+xwZotnZr5V
bYS8t9pJmVsrIkNcMn6UMqMcnIEj8xqmZVLv8drD9TiX8eVv+nrc4JbnyqbJgHcR
ocgEk2n/0YPwxeNeLLXgCheK9cozqDH9AgMlvekzr+JfC+FpfVUkJSnKggn6/vzM
VCFD12gCDuZSmnqmiRtjy0U2FLr142BpLaqReCsDWgzTq6You0kJ4iVpCEFPQX+J
fZMh393bqiIpJm6E5lOPKJCS+iUuI6y9MiekmuePj2FZeh7YnPvTxTXl3T01weJW
Vtc5o7FDyCawiB+kyYw4EFLFm/+6Hw/bU6OsQjUoI42SESsbDtEkXXS/yAXijyLz
Osqusbpjc/fk/xdZWyBsjxHYB0+AEXjaXcCDtcsx0snShrJAS4brMuG2muhPMqqF
l03mBFdocUrWgOYfPgdjiQfmpRGDAqVOFHvq8Gq6HDIHSfwbBgRbn6w0366JDHDT
wz3jr+VuKAgDXJRXT+O9a6hK+Qp1RI8DEyzfZPLCMtgkdDvzS1ngOIRT7Om+0gDX
8cuMKMuoJ5gSSLNsphhyTKAZbMlr0I5WGDwX0RP8p6Pi1rpxjmZJk64wbVjdJqZo
VpQ5Bv5dkZpl/KhL8BkdwKcrLkGcRH5uM3EOdETb+FYAPCleIBfNg52hkBUsdBX3
z9DeJkV6gZ82otZ872RkWLGxJe9ts/rWtIiTcGVvcCmWCJYhchve0Eme2BS1bck5
kMf/gP7+0wolfk/k0lEzQD0XNSYE41KPF5wpt7mpT2rW7CRVFGcygdfwDenaSgn4
IGpGbJFQIJeFnt8710F40Yu009yre5FSxMZWb6GqY0FTgWicxQcza7d8Qxu5dKub
NAABOOfT7YOHU4sRhrmWJQxKbjdbTmmLZzTwnY+9Esn2evIgq6rWSt1EQVazqOyM
xSLCfJ3NYSTtygoA3TPx2dYxHAw33dd/q//2UX3b0H3DU+rbPVYpY8uQ/CNmxBGe
AHGbsG8DZ4W5DS/AR294Pe8hfneA2Y79X/c8p63JjKf20wYZFgd3BNfn3JmjLbZq
A3xcUJmw8eOChsOic/Fl7swdORGNclGWL1uIZHvBGYdMCcCFJBLeHR3d3iYX+dfx
xVpKTKc8yLNlVKJsiPLL9HSrlsh4NYPRpZfW7And/Ojpc53D+O4l7zVFQ7CqkJf+
maDXbPqeZQuzrXKgMDy0MHR4huhoWvnUyHc8tcCgkrYNfNJpJtgMFYf7s12r8356
bL3ONiXjJ8f1clWm1HLyrpeRIIKyk2ZRJxlpX/PQBEI3AmjszCLuI+agOIPrhsg+
Jp/tj2x8nlsBOcw7JaBIe9FyLr6gRCD9+LrM4g2koWaGRHEUcWGJoY2ANR6skZew
18FtNTvKQ+MSmLJGImowbLwnvosm5qaWkOwjeGFYxoVQMzqh3OfOi0qy058sa2hF
h4rtnIooUmHfrrLZDMCrrPp+awI8G6BpjwaO4Yi3HBTLgxKVEMdoEzBq52C1+dZQ
0HCEcv7NM/qMpMhXw6BnEswBronQqcp2dD/VJAYmBO8gUGQZPjmVUv0dPrs+zONr
pHCrOSi8DZX0O5jJXTdHcpFRuqNjS0lX3iBWUio85xek5TsZH/IZfXi3pOqp5lND
Y7Vmgn1aFDy2LKd+Gu/NxtUITktVxyjmJ4pG4VpmH7cs9b9Q6uq8fI4sMTAXcTs0
/cfkPCgW/mnKJGFhEYjNCfHNDDEiVsKEPMx1VOir5ADtQO7D1FuzfZmonixlHoFH
OU+aj0thygE/jirheUw7XKgzWTtuMSHQyyusifSD5uSY/ULVsGWkIRuZXPYY2iiM
BjXXozsRBS21MdcpEb8CJXR6+ZvlY++rkq18nvqrF8fmT3qj3nzcSOlLfRmkzXO+
prCHL0NOpfXk6GH0sveiHuFbIfbjFHUU2mk04UpVOaqFGlhThfYr7k8ybQe441nu
A0+xrGm9X8hFA4stNNHR7L6BzhX/kWuh5XOJGISuIsPXjxlYmGTWtuBVyUR9FzWj
/iyYRbRLY8Y9vKqA6H0gKXZo3JuArhPhgoNbghaYydMCojxN6IhqbItnrowKL67K
eS4+e+4QqnUpjahvte29wjPaesmFTy9nYYTozPsWRHlC6ITv7lYhL0+iCpP01MO8
k1vHqH7TDKG5v7zxGswpi13dfto/e0677AkamSkDyX1VsBWeqerLazmbsPx3npWt
AxB3+kPTHnhogcrEcSlbrDxkLxvDxmBCLU/6wqaxw+XfplLSdYrzPNFVS2M4KFOq
PxHfQ1ZZCEVwdKfberjm4yZOp1n8sCtZ/a7hbThdKy6ulkTU7qXRJPgu68jBIqfQ
cGWEolUkTVzaX1aqMVzhi3ygnuOv6U7Cw3l00LbJbGErtKBrxG5lUGACJa4gLfbD
yslaxHRccExf2BV60TOwaFm6p8GI8Wv3VsTRVB12GwPoyeY0ujyHOeyXRXNJU7J1
6+FdlO10Y0iHcx319ct9a2FOdRb+UjdEDD3w2Ij00qZS7nR1oGcYPg+UkfKRvZ4h
3IYTrAAjYSS78kr+PkdNcv72pnBC1Ywr+z1beYCY7DJyjR1Zysk4j4KbFykLdUV1
XDEV9JUcCX/ggy7IB6zZGFmmYfMAhWVb8rBplYk15/yWur9oraT1IAbNDEzvSD9L
EwdVRnUMs5oed7GDWbaOZmDqGVtO7RuZDTv7hqv5LkXhSaTGMgfOWPSrC0c7/PU6
5e9vB+ohEptnItvvga9sl5ERVe7D7/2HkZyk1y+PerDfr4tXRZ54GMMzKHvjAuSr
pFZlzN+g/ZUiI6en3Us02hOhtex3bMrjFBTA9EC80IfG+LUQutm0yZ9x6rsRNB8x
d4uaieuG07R3QwoVxO4xwsdZnyNurFmh+0QO5Xm4/5dMagohaQ5GhicqM5vZqlCA
QMuxQSp9bqqg/SqYZW/kZ/8rmkIrwNGItZ8piMdDXhxI0MMEXwg6EiKzfuP28Sos
Fstpw+UBXIoyGgdkoUqzIZat+Sb/UVxqNQIUiul/OOMUFOFvnuxv5DWRUEeWrU/f
0Oo56GCQx5MJtYKYkDGRmfX0i1tK9LMzegx2/RTf+frklwKH26unJyohJkHQhz32
6VPMPgtftsejK3h1mMXLBplhzSEBuaAKRbassiQ2TaS8onrEqZ8i0/TIkqjCDXGf
q5DSbDk44HMZjHoaOIkWeCCDdZJOeOa58b/ep+71X8PzVDEyPtszKikpbhhBt7vj
hseJWTRiPdJKYOZzz87ev/lHELERWzwip3BTLu3Dj0S+AAFZEAN86J66x2g/wd9x
LEmWdF5/MTl3gBQ6RfP7o0Rfog6vQxC9RFfe7VhJNNA5cSbs7kRWEoSeYsZXNUqu
sDuoP6u5G9r2YJD2M86Djr+P9njxWK/TlwB5bOZCkq/lU3e5GFvQTXK8mypa3DpC
nKHYkAnE27qpSI7ACtV69/oEh/LK06VDsvzpnBK94tIuKiqUa1kJ+01cjSsPFXwS
p0Gch3yy1nrp6k9pOyBA/jxM5jDgtoBYWDqob/CkL5RFJPgAJhB7L8Pc4/+gV1or
xbRMjC/wJLEeZy/B64Jd3FQtFmSynosK41sIyfVeNpMbce8fZdYrj/hWefGErg0u
YCfdIUi0b9tKshSULMzcHmDGifyOPHK+lavBvGOU1WmhvgQTwLcFoC1Nrhit1Ayo
cXuZFD4brj2z36W4JgWyF39ApFC/kZJPL7PuWgg1hO8qitxUcyPeI1V8hTOB2yej
HYpNrUkwSqC3CPdinT5dj1HrO8U/OeUzzoPJucp3N+Syn/qWLGsI1QJ+qY0R+yUX
rjq2/mNazioRztXnQp8r7KXKbTECxRKENSF1cReANm2PS2CoE6BYoMR9AFxU2aZx
PZHHrZvA7ZHm8lJaQaqVxjYu88B0RJPrNrYjA66Yu5GUdsq4tJpHES3Ia8tsM737
oqE8w6KydX/Zk/X0mhe7otYvaw5M6kSckqJ/nOFvtvbvXIzLqO39EJX1nwZEoKX2
UDXILYWiCk4rUBJZkVH+DBTr3Q6lF0rTCz54UBMWQjqFAY2OLkNnab4SvKbK2xfm
lJ6+ssHB8btc5yzcBxyW7r6Evrc9ztEX8ccTz4ecLEMAjgGRFYXx8B1xmMyIzwTl
EtM/OezvFkibUBvZzab4Zh+v/yu2gXoUo+yqP/ExwLfmG/3ot9LIiRiv2TZsiPYA
9PH3zUz/z46EZk+lI38Nn+eUNGGj6CtFuLH3b+5ST5Mu2LwH5iN72N8SjdBgCtbB
xBfb8aSWXI1JxYBxdhdbn1yMzqDceCC9T5blvuxl7vyhik6GSQE/0c0e62z+iMET
6g5ln3qQtNdc8UNyM+CYZG72TYnzOguzdqMeMYw7lCTIe7Ia/1GHJmOriubutmAv
Li3e1qgwMjZnHhQT0enItzyzJ6f4h/OELsS6CehjamLnKQneGAbVI7ju14AI9Ylj
pN0gM3rJ3DNsYeLHf9UDoT9y1C0VuoWxlGw9Xec3gUfNrmayWqfRaytCVH6hQKr1
5xXRDdST2cu6gfDF0AwlOIKfFkrIY0lXRITWdXAPiaePTZAtLsN2Ix7An1ojLtLQ
KgS4vWRKmkzc3lmCCGjhHJ2bEdMOybPfokTtdAyeGU3Slrmxp0t/7v9E1yu0jAfY
x+uC9TrhDSN2WxIhPYFUiF3vMFOj7w+0ujYx7DBuosgKyUsp3o4wAWDSPg1fmjL0
v+yUgbsOai1jcoEuC3RrWgIgj6AltXmkKmBtrVg9taHYkMSTMP7SKeM2BPXx+OxF
TabHAfvZm42oYgZACOeA74dviUisoC3ZXFvzMlsreDqe3zzRQB/MMzuH1F710Rg4
6wRtMBNz+OJZO035CfRMs2scsMI6vzlKK0Mms3OaHpTdLkp+meP7wZlPIzYG0QC4
LE/OcjuyPpxShPnCQsiWlePzGyW9O9zY1yXQCAYERW/6ma77d6g/5E6ed3hpGpo7
v8oqPurjCqovN2sAIxx0SXzVYtv8ouWkX4LwUwASZcMj4JIEPrG6rPy/8hIkXppR
KUd0heqmd+xAZ3qALqSqqLP6mLjQMhkyyAU5RNI/jTEVGd8krw6fXRVt6aBtmozF
C+p3bcF9BygoEtzP5NmYIaHRV0lHyXUH95qzMgBxj5IAaiU7TgrQyEjRIUqHAwb1
QteebfLmeP3aIsoOYj+JemwQjEc/rKO1Kr7gvYClX9Rs8anBE9oKVFzFZ3sKqhOn
LB1Z3bVm7FWMZuS8mdDpw9zmRxI+rjjAUiLLIL7ss3PDkZe7aRYuApi/aXr83WKw
f+UjcZWSS1Zw84rUOrHDjQHt6F4ivRqD0y0/wj3C3rv4aldKQ0HbQOpvZ3bEm0qk
1oKFe8ep9UprlUdxvQXqRz3VTO55FvfSUrGq0HZguCAGyHotb70OIyvrWlTGpuKC
G3tmTQk0IwENDg16Cqy+uMslJjDH4yR0lhbywVwXSdnE1/YhzyR/P6vw16f3GGlv
YkRlOt0mdmkH6a0kAsfub9GPH5RUfaMVsJSNXxJKIqqyjQwk/8ZrbdaEClpn/PNV
kfuzc5TCklgvCNzjezpWuC1tmVR6pTSVCOBC77/yb57lQUdj/LR+dFP1RVS/DBAa
TzQi79A7LnbbNBAG0VoBnIIAXx1Gy3VnzDktjhgP69oIj4res5+SMNhsHmtmLvTt
mwk56zXKgAWjJDkK6eWvrnRCkuLvX+9IL+FnI2YcZPPJFK79g/0aYaR5GosIoE17
6I0u74zTjbez/+kyGmKlv+l7yBzvBrQt/xyuINQQPez+zPEZOTfQ5W0pT3t/uXvd
yBEOTKHhsnU1COhIQHXXxXj5B/g7sOUhziXE8cvewGMvMrPRpASY6PNvx1OLK2zw
sNFMWB3Q0P4Kr+EzWzI6LzvBqLgRlHbVFT/LKgAdTv7CoVqMjgZP228MC0tdQcxN
HWSuiskyL7/euQE9dxhJyTttkQBYAz5VapKaYggwC/iIILg8RFsv93ERRIVRa/Wk
RYQABeEbIvMJGFFRf2/8jiA7123NgXoNX7cDVjRIDyY0SZqItVnYXYw5BvcUUDCc
Jb6OX5f5dX6WnA0rJSVIrWscJ9ZC9juy6MvCS9J9w4q/nQR0Fm5+7Gr8mlzY2PMf
UR6Mpf97tI51nxJnAdQLWQZ+5yeJV9QVLzgmliGSpiAmuMOu5CdZtHZixAJ1Dovi
vKszXAgm+xgeZ+xAO5ODHbVv1KPfdChrzvnvvJ0/dcKhlqf1SYWCK6oVEy/oY7Jp
DAg/ZrMmwP/fFYEjE6IBo6SBklwt3i5lF7LY0j5ocIZeqnHY1jnDz+EyQ7UIy+i3
47POO36PyVEaOANNlnvLppzyVSFXFlL4xJj0v+Lspotua6JqIrqg5eD0iQbCUQWg
38Az6cTnqgDJTlp78blCEiVVf142G9KGjmndnYmLZc3rqcrnb36IasBRQoaAEMxG
1wvikCCIZTJsibZMoUMJ1DJQunIJEycQuDXwVq2NsYGCg+DDcY2SD4Qt90xxZtUh
3hXuVUHS2qHodrF3h7llxjGA/HkgHnDp4Ns/AxnIevsuI5d0DC4zL7ofEesmTAco
7xhBt+LjbukmUmp2Fs2ffQxrTEKMrEb99Hc2wV9CkICiZwamvEVwh6KV7+rRXfNG
+dXJIw06v1rZ6w6D/97C/93Dbpmn9cwjCOJVpYOO6ylz+YKk9pFrE6qcezDBCs3F
U+fDzQrCrv0k4G5G6VftTG107b8SokqQWbN8JKViv2erp9Tkhnv4Clnvl745aT+B
RtO52VpJr0dgTcnExErK13qkBA583wlR/DJ0Jrk9XoxQu3Ivli+DEcaVwrxOjiCK
FagcPSkg3UbMNoMzun1QXzH8i5HAxOVCmzkLtF11pUvw8rU6tQMiyOOiblqskS9M
7PUzr2S9deAzck+0c7YnDriVJKmq8hWkeY8GVoZNaI0xOqJG7jaHvJsenXAUS2OZ
2I4O60Y3WI8qYD6vw9VZKUvkNoALxZnD0l+EVskWYr0f514Y2CApPd0vMtldtTsb
qPfYD6/5D9CkwFwfuq6FbYu+/zJzIfJbRaS3qCqBVmgJ/m8xApYtumBe2ymGJW6T
3UbrZbuknJmdfTGNzWM1scwlO3VLsJ5RJb7FNQiHveWpNb0T0iMFkLKiAzzIyr7s
4z3JIvVWuDygEyNeQ+aJGOx71TnAetqWsHX0sMm+V4ChJG88CtORmGRo1cUpe7UQ
Zaxw8hhhdU9zfDX32UoFraZbnK+ARp1aJxeYF0iyFLA1yOaUNDsB33+cI+Lflkym
3xyYqyXf/m/VkIUIQzQ2PJw6/tORBRc8ofZkJZbFcyUYF921TNxE/Z9jelrVCMl9
CHRSPd9OkkkJTlFAAn8rM5GEIRPTiEeqqOUqZ6HyRy30eQb05z997rbUth2gj/3W
4dwuzyV4X5LycXJTCDzSsppHBYhpiwJ5pneYs56GqjKZrBJN1R7buBsDF6mVxXeA
d7B0qcA5gq48yKoclRrx51lkyM/qlyX9HD+vgaj8ni4rG67cu6244PoMqyI305Qb
IDVbR2DJj8N4VckdTotcsqgVxnovrEYajFia9VL5i36ZU3TZGFVnV5YBaMqQyylx
GVQ70WOtaI5ySOMdSm8hr2WbrCJpX+yPydl5Sgbg2fSr7xbf+PY8neA14nn/k437
0LJbpJuabqidWEThnrfwRIqMEdU0NbwNe5ZUevAiu3IfO012cWu8qlvN+EMncEfG
MQGd9YBNUgK9Oex8bFrbxkZhDUBS0uIAPwYuW/UkB8i6ic2vgWUaBRtqdjkSTIKJ
lPrwsQHS1f4dz4aBD8g0gOv1DF8fxTsQFD2VVFv98n7pCLNBqA1wMij23qYtnnt0
VhpJ+Uh/jL2KytIKVZiCHsoD/MbqIe8gqvnPnl1O+t0V2gCQrrOfXWitSnmxBlqV
HBvk4kSQX70ARjkac7Mq8DXzQERKAFkXdJ7Lt95DCcjsSHzBJW6kHEEIYCr9WT7a
rz5HSFlznA+MAN4v47v3NkU8mnnTM+7Qaey1lLZOJR4UI+/cIPWAkc+uoGdr9SBJ
VyShqic4ZYE339rGQRiJ93xdAJu0SGjRvBuwUG5oGoJHG0IcoxcM/qDGztXA0MK2
tTXY2EGGgbNuNymOIkcU6+r4nxKkt1COhXmIVilCCVEJ8N2pVV4tN3zox1mL404B
sFviZvc3vhUIQKCY286QmVGqpsBVc+IB56u2tKgXiMXctV1F1bpInZKtqttPYfhi
jKIsHyGpeWVkr9lKtzW//Q2T/oskfZaj2+SsEuw06CNLuA0bNCZbTnkssnKmjJAr
OZv0ypxQyDRt3WV5H6AJA6tGRewEDUi6XJP8Yh4Ih5sq29H9rCc7xtt40D8Aw0TV
3bgWAmFycc1QwX8qhoXPhx2g6mXNEk/y+LtqV/Do8FDxz7zFZWQEHLRUIkX3RO1b
4wyHKMhlgTYdbYIyeeeNM9FSB+KIUTg4M+dRP6HbsTa59iIbups0HGqYZkwrBavL
1Ob1484f7L33VizQ6bJPG/8nyeM++FIY5MlC9ozwcsXYTCWAe+F5/pCUvHBuSVRJ
gFU64o4gPgOLn63CA/9LF1+Nsc947BR/MHiV/mxRZqejAYnxSIuHYiWSaneuRh0x
qGCHUa9fjnHPgPL4zUcG+YVBqegBeswKarfIH2ruG5ZMLCSk7KeyacD9m1Wb+gds
UgNstiSIuqqRP9tf8tg0Zi73Hw+bgQVGu/4ge8/rRndKjhdOHLzq+k0H/XRWDrvg
Y2sKtOVR3Q8zohicg8WrmhZvslcWS2d5eY4MG0qnswV5oHr80I0LKJouhUCfCNy0
kded3mDnuaIhZYWgvS2WTkGAwTr7dPQl3wmFIU2FnlprTd7ygnolBpyCV1TTyPWt
qHn5i5kS4u4ePyE1Rzglht5Kv99aAdxqws1gLupIE9VO1UUmHIgOQLhtFNMmm/U4
wv2JTO6GDo4cB9kbsZPOzXCFv2K0h5lg+qcvMn1XC5FOshM9+Xvg7eSalV+gTT3L
QX/y8gYLU9YSLu+ki0EffdrIVJmmFmQAPZ62gXy3rq9TwFxys2dt5T5wOqWyysHr
EmKjPYYrvdMM+/DdTK/5J1zgrjDvHIuzv84lb1d2peelwPBhnwQw9d8vf2XJyj17
5ttDgieRBMeQUGnD25Xqdk8l1Xsa+XOU8aT/BRuVw1ZQzQQjpS64hLYgcfimyfIV
2uVruLeYI8oV6ss7EjnzOch8p31GH7Ki6yOK0UJYV3BLZ3UzSjAbansf65jB2txR
BI8V731zHudxKOIXqxoANmG5CIIMnV0Y4HHEuQnD8f2KtHoli2JRNmYf96aMfPV3
DlznqAtIkFaDDSa+f14PtjJWseWDRQSs6pupp8ifFL7LKbRPIev5arz1JKyBtYid
kY/Bm9RlzsNpw0jw3RTOppDvMWiJWD+Y5sb4pa5rf46aRoJhW+bFZvWKh7S/RrJ1
HbkrHicMRBg1UWlQV4Zf72xkI+fySmzr2SwkswbTb9qXI1JmT43qAYvmjRLRJA9j
pW57dQD0Ik/3gb2Y8NjCZZbkBNqENN11vTAgdp2up22Z7AHX87QubQiH8m4YLxUt
uR4/Ha4QBcWLqraPje0Xp4bsVMoAYQQKx2imx8gXfcTewoMdfDsG+r4RYH2+dIQC
7ldetLztyowsB1fmE2xBkHOitIgTIF5HJfMbfHJnuTj2YhpPwVDlaQN04x0lfREz
1UqToAiSHWG+vmmmcWj6G+BXYqm1KrRVrzLh31/xWZJ45iYzKwhrA2t/OeKK+sw0
VC9jqwRPluLXRtuRXYbYmjh4UFtxRhmy+2KioBUzJm2TwEIK2HRdcy/pS67gFxII
eHNyQP6lThakHyKoUfIIwUgdq5SUB7fYKXoEkOEwugQwGpWv3Yn1a+K8KC+K7mka
vu/u10vPgCzF35UELDkEaVHQbwM6YJyyOJB+tv7hPzS9H508yEK5ZKhHu9301XE2
4LTQhddRB1I2sJbzXA44JunCV80BaIdzanCHkTRLAXbDhCcnOPbz3bMRayhgud9Q
mtoLI6To18Ft22WVl5MmORu+P1StIGX45lMA2QN1U6mF7j3Q7On6p2uGBpFTmGBf
D7dEVhhG/mOHYYeRhpjens9zwVB+O9XV4wRjFVzqePNHnnBVx/3T/zxbucGyeNKn
Mf2wkdZNs2sQ308WMCANmIXgir4Jh45A5k9bU90rHURpfhkYD6+hDzZuAU0WOp49
dUvuVi1Y+1zPGGRRgMuD+PBiyKyeYrXovnNAL11Zl29D4H0vo5GA0M7u0sLwsruN
o2mbxDdQOHBq0OU7oo1zqWbPRnSHV03Fzz8MKrIF1ujeoHZXcBTLkerri28EHXxZ
k7+z/JKoNbGKU/T2Ln8opAIu7U6rsAAn5cWFpEFDkwIb6gk6j3EH2/MRUj4ynVYc
4mDhwetl2gsO/DN6oA/eRMMl88xc/R1jnYttOm+BH1jSlIbYkfbLNL61JNRLlfpV
hJECt1za+wmJWubMq4o2VB2WPe09f7lSCcF2hcfPVMS3MDXiSZjpQlBBN1AGZ6Hw
MQapXWfCTBefOztHJkVn2kVJ1sxINt/DnhbWIKwpBbS65JTCZnc9uC/FtVZ0qbcV
XVDrzABHzVCWKTv86WcerHmIgDovcpsGbQxFisHvXfD9L5SpZbGsWhVm2K0/rge2
e5LF4+jM+9i3mVd2tJbQb93T0rQUwBGtMkgf2PebcS8TCoVWFj/4h5wzptpQxLS8
sTN51CZPql/24jiEZWTGoI3YiAO5s5LRW2AZHdr/F5QRRG2IZ6XEDSRAI1hxs1Gc
U5QCqtyEmqGhMiEWbsJLxL3iujbgXPtQ3b9oet6F9hdFyrwJl/V6moZ/CQdKUycp
XuSyju2KbmrR8bbnf9vNXnW177bDCkW0dp/Eortz1TxAbooRxSmJr/m9c8aFP7wh
ZglJ2NHXu7YxERI9b1zAbp3gnpFz73OjVS2WMw1NwA1W2ymBZ/tz1fQRAXTKE1cy
vJcfemmMTlNMzCgdMcN346YA7pH3wxV/aw4cRK/KhqR2TKxXZJ8Qmy9KfUHEVpzD
EYsjN/S/IzGoqQCz7vTKRQklxpCEodXSfmPBxe6etKby6RgCYrC3UIAkFo0DhnDh
NqKmIztygEfEtmXcKRRX4Wr3ElxTIva7xJpdA/s8rQyXv7wURs4IeTEjIJETnQoj
eeq0Bj0bHH4Hiop32CG+WjqphyTiI9JXhVclVJVHdSceRh39EPXto7UZn4+e45g5
kkwUGSDVRkLPw5oU1kLrlsGAXeSnt/pusz4jXg0oPyoDExbsBSuBcyTCNRHZ/RC+
bNMr4Y3EkmZcmy2y61stvKvOwP3xJA2RsOXpjjvoP4KtbOSpfOAwdO6TQP8tPiSb
MmUqLOxB703l2ny/9mVI93sT1CWpucUOUNhegEKNrWaDVnUQazZ2lCPPczsuvBI2
YQfzgiTo9IuwvnMKNN8Vzn2+n78csXj0GtYHhapUruIOXtcmBeRJzM6T0g6ZPeZI
71RXNuWkKjdruU18UFo3AH8KPxv9Pck6Tm6OApZ8S7K89TAARHyYXTAbrgr3eLOW
hMjhuT4tGrXuyB4nFRy3pBK0dl2PgppwrS40D+XOpND2FBTtV0+2ZTZF2NlRPX8g
xV3umNtrCjX4yihUwX1yoayLILelfMTZH5qddCuJHA/A3b8syVfGSKeIRfqyh9/5
5+8Ycv01vbB+IEXHVhYT/5xAZa6TuGJ02KPsUs/9WN4kL/6Ra/HFWCydpkuGH+LT
fyK/CArgbQNDtWDZLppIYT+fiURGmSYNkNmUyS1f6CJs1WoHGs9OSyBe5Z/kj0Zl
H+9zI+V8ilANE2FnMgERl12dUnSifOCFdu+7T+pymVzRzmR6JUN8r6K2GDEHskBy
f1kCTxKIhR0GIRAVO4LKritosFhx+mStPQz+9OxyXXHii4ilqqMSC66fOwVm1NPN
80PpJRau1yCb8X4nHMZyUwKPh9T/29hveUN3aJ9X07UO5nuDuj+jqIF1SUl9xdZI
5O+n1ts+oKIjGH5GHMEAoqW5XaDKut7CrY+Ejh8yVDhVcyD/ZQ9CtJpPs3lGtmX9
5dglxyQLDNYMbNhABK8X3CQT+8SBce5lVqJ9nT7GHYlJSGgqU74JOi/Ph/BJt45S
17PgGwdPIkFIn4/UaRh+AEK++Uks4WXKgaWxMnLSFccZoAn6cwL9k6HN7iO9Svdi
2Q8MQm2sf6CXAXn+gJRfbHJKFUi4LWhBotVmCeszhG7zUEbFmam2Fi17EeGTmRBL
tIDirzq3lZ9N36NpLonWpJVnNFcz539TI37HktbujZYDzVRdavU46iVM4prSdqi3
yt2m1mWYd61bG+As4D0D5ThO7BktfdhtRH9BmpFJe3ttTrm+qHCokvxvi0sSUZh5
MWc4uM0CiLXInHQGI3R8xolxQlghSJyrzbw66FghqPE31b0LPu+cyWg25d3nmDAO
ecc5JlsKQYkwnNEeiP2XCYupxCZWwrjy27Nc74/GwxikNGEbHLhzBiXKAKZLI8xs
HIg44DpLEKh0c62NFtBbFis4aaELkyNnljxyftefjrkhfOnpHWfpuATAF9rtZxur
NJcQop5hYG2jaNKzWJHVqPXM8t3/LatRiws5UkdI+fyLqR9JxYeGQpoXP3x7yxiL
CNiYzBU01phvd4MHSM2BoaC6Jw6NiISYsqpk873qYS4/ech828HVo2sdgrFsWG/R
roV+Yn+KwIwBckkfsPU0h3fSIsRbUiLcONqzVNJ48+bV+VCEUoPjtPHnPGAwGMex
454yVQWVIvvTkpHQXjpt9p51s46nJMIS9brj5KMmt4CFZs65M3IWgciexgmUKvJ0
ymmbiFqrr/9ROpIi6+cVvQsP0cMJOdk237va8TBb1uYK8R4kYdHLGq+ZTM0sIYDe
Z9cWEQybau5+dIrAL711kO+uZwA6DwvJKjD98eI0baLp2tvMs+PmEUHYKoirgyak
1ZF2G6pUbjIRgMgWxmqZNHQJ5uWLomTUMD4IQo+hNPzHp7Pu6ujY5RgrewVML6BR
nrr3sr2Wc4yr/2xzVzIux2K1L2QFozEb4MuPgfTllJn5DUIJh/sffDHlGA3H9W0p
kSNVrUr30vQsrQMKCwV8MSnQqYICBD/AJbK4Vv7r3YNCoRrES+PfTYweRrnzyYPZ
xXrz5p/AnLlONCAAQf/seAyj6o1udIn+iJZe7cqeQaC//bLAvj3FD+CIG7olDREq
djYZuHim2D5Fr/mSYkbTIdGUisNgfWFBzLXeOsKb3BO9I40C2bx7KDcpCTNfAWJU
oPCtU8lV5vTJpyd7Naqofhz9eG+aGDQOZwi/UmIwNXqcySUSAdYvm8luzJsZmb0g
6OxPmK9D93cAz/nf9ZtGQXH/Gyyg/lTblsCY8CI8m4D0X4iSaXeJ41LKmOqw6KD3
JYHhi9xPbH9BOPua5c+3sKccBnxLrFiMZOSrrECX4XhTPm1HxGomrkS2UfCCE8pO
8gQ9fa0owMIYCFQVAvO+ij2vskqCWS6xiRJ6s1JQk3VCKvd1nLeMHXzFAyT9jwBY
Pw0a2uWx+3h503D3U0N8dc3OWkaQYbZ8kaXuylN/DRxol3jtlRoQ53eGRX2iMoyE
ZQXuuQZcH47rzxUVv+kkHlXucAOBVsV/jmkO3xyjCvS2RTy7MR7+lHeruSaMdxy/
j+zqjZRbPTAH7LKbsieD3rsvrn1BjeQRlwOwJvL4Et7tp49YW6NPEEWLCBQVDD84
gEDuqG6PWK2/sS00fWfauGKfCAEtnxJtXEOpMcVvosVkOjgLj6tPnWouXtRb/3bD
jkwzVsHfm5jvuViK4XoOTnMmzJZV06P8DAsyYSn4bpQ2lutX2a/imxPkEsksGZxu
/NQkP8XhDFtFRMahnl2Jb57KV5FsZFpYBMSei3MffpJf5G9ftNKXtf9ns6ewKcVt
aMEriwNFkhbVao6/jmg5PXtTa6y3i6pNxFblKqi4XAMOEQgSSRsFrPwJQtLJCFDq
5ZDrYrIIdM1Cz/cIbmSg2HHTXo/UI9J/65oQ0CpEoS3PmiC/kGOUg3Yymgcx0kI5
yDfNqbclzGPnFmvxaO8wnS6Xewvmqyr1bCDlCXY9EwJl3Pxkd9EqAzSBVIwIJ6o3
ViJwegz16jqP0i78R6l3kGwpLWRLoQBXWPVkBZvENQVBgd6mlSjEEvz2Xv6SckBl
JX+ZsjHoZtHqnkeqtfLI/jd8x9CTy9N3ggbhdRV+9CpwbG1J5ZiN43BIPvZEjvPn
LkDKeTTbWy9Bi1abSe5aK2474NfaDG+z5Be8KCus0ipWWJd6A1hExjph1gQPd/4q
MSY6jmHxr4pkKZRbX1kll2Ykj3ku8yxtVAYh9/uDaIQq9XkXypUA38r0fO0iPUnF
fJ+0nOAy21wu/nX2NPwfNlw4mvd1LFzw8YZIYqwXzfxtkwmTFAvrMaAY4V29hNoP
jAwtywsBmA6NiZ70wtCyeWvDQw+G1vipOiF94TL3YAAgvwYrECTubh5wk65GUfpa
lzDriyywpJed8LNNYE6AHrX7vY4fyeCsWRoxiqiyVydjijcFhkoRhCclCcN1q6o2
q2o3AAoTHhWx/78WKeDptBz3y/D3aQhJzGeW9LRrR7ZWHmAQKvuYgXrBgyWlDz0E
p7HdIWQl8ajsCZlJ2oFTcR2p7k1zcvWfaL0yKwy+ocBeuOhL0dI8ed9av7ZYxvq0
VH7QZA7VJDBFgFY4YUpbjSHi4v14WN1FKRKoizakgYS3sN9ydDiee7Hk6/yspLrt
2MEBvR999+MU+2zqR1BDjCU3YlIXSDAHPhdwIKU7rMpmqun+ttGBjJv7VBYlCT+D
txqdcCX6jA7l9fPe1DXPUhBFPkTyrEHkZpNoYK6M1xcuDlk670hQ1aq0WBpeOdu3
rOuUHMge1mEuz3rO0TULtqkuNWQnlJdt+s2aroKJdL38U+b5EzPmrOMcqo5CRRLg
bZPKZThQFtcH4quOTo9Aa9DaMce3imT4n/5bQlg9VgO4vw24CV6EcwiRiifOYG4a
RNpr+GZmEURWbepYvRSQBvUcRF3MZ9ouucaZWyMLL4XEf4oiBIDG3j3mTEMnAM9M
iC4vqvPtmDQ8xmwKQQhJmn1fzOTqnjs+6mmHZ/NvZBXyzniV3FDh02N9/m1pOQWN
1Fe3s44yVeBEoQDIth07OAiWzHG4KFLcKgR4uRo2ZWXHq1VnL61iuI59QvY5x20p
4Z+KoeAA9mWVNGhVeGsJAlbxFBm6nid+BfF33cIzMWIB9lYOPCWdMePYXxd2l37B
RAT1LliM8yaWyUtoNqsG+wgFxUsyf++x/2qxu47gyloKhgPbRXYYVfq6ZjaKG52G
/auT7kBsYZQzEg4WBcUmYK88lL8vSY5HLe5XK/scGA6JZDRRrghY1/f7Ku6dzoBk
o9UKDBKkkq6pgQUMhryJrYDzkfanguVZf9R0ic3jXojnSXTWFZetWg+Kh8ysFb5k
6O5iJuvkmfTUfPeNHaTXfDFq6k/nsyiO/yFrob2XLb4/ob9rb2CkCGuGzF0WTLAL
KDXz9x7kQzSai/aVrnOtkoYT99hdDEXkFiD8YSffCbW7XVEMrmyo4cKOvFb2I3Xs
ApeJEZNsgp3QW9x5/CfSQxRFqMMcWtdoAxAKP6GIQX57OVx6Vm6FUTsJdb5v7qva
hvlbPUMKsmY0CM7iguFMzR8AlyQOid3VeZde5QHVceorGMmcBaEdFwqaZTz0SWD9
g6P9PEyULmFqGnGxK0A9nscLaMx+fwOi7iAKrTpqbe8pst0TpZAoxarFwtzXSLUZ
uUm7yLNrvy86TAZxMxMqzXy7Fl7/fpMZCKpPdKLZPQ08XO3OSbwIO84tjj3vITzB
Pm/2K6dT/FZd2TbKZhQjN4fVO1Y1bWd+KjqENSCMi093cSYthYiP+I/hFFBbg2Hg
khHVE4/lkP1agsH+Xu4tnL+aZQS8ycD5flEN5t0sGA2C0a9Jl1gxvzSZO6EudwEW
GVSMA1CqJteykP+IUrl9Xq7QshSrMEF8pdbHtdjmyF6YyYPmYmlgvcZElE49zU51
Z+FyYYgUWWCUJGrt6vWuRHqatI7C3yN8BEJDzX4pOKihrFvztxIURDexJFmuKEqa
of6piDIpiFaJoKze1/AMxnXdm+gZ19i68uyxVvG7Mdtd5mvFxt18w/cF8qiKMOv8
bnYKknY4aYOtXsui1GYkvq53FexjDniSUTkqOqP9rR0wRtO/Dpfuxo8ZzuqE2SdZ
AdR6KXpxDOHMHuN0mBeKpMNG72MqOa/txoiyUQyLe8QGZ11pE9XAbptL8O3D5mJQ
fBACWOFsIcKNVVo7fxofLdL/MgZbtnP1auyRMm35WqftnU1kmC1YLOqQ/cNk5g4Q
3flAG1Uks1oa1+gle6zHsnm2gV72sLLNpci1pTiQ5p0OWFKRbrRM/cZPiqXxrKx/
Ia5UsJyIWxo9RBpzOHwLBdn1VPDcx7M9AtkcoNO9rOwZSt6RCk/0YfIceuE/6F2g
X88ui7ogWOdjTMD2SXmRvQkRd85HVKeXfyzjFeEnOJdqrz9Ib0miUGijRzR1Fz9P
FcLNWu5p5oagklMUy8jMnN83csUv//2C4//LOhyjB8fDe3bY7eJNz0+jys1CXqwO
gEd1uGcKp9jrfLqv59dV+3jLDlBorsFBkvFy8yjQbd2pduRULP/Vq9+h/lMEnGi2
9g1gy7OC9qqKGtS6jt5o/TP0L1y0Q8wqalzcjQAY9O8VMm1rwPPmpWwirCNhUTKZ
Nk9vSXkrtWSvPOsIDcMdotFnhokf5dz63hL5/ZZFqAWBg/m5GoV1GpAwGS7r37Re
T2EeuYdppGE5zeSfnhm6+mce55V8prV942iBy7KhrmwmxgkAF2dMq7ZnvAjZzBDm
N5LiekOdCXiuIj8Xx8pimy19wFYW+72FPcmbU70fsWRofIAkH5ypGaOqMf+sfB5I
fKBkopilUIlqmwJ3yZ1wokwPue1Hkk6Dy7MKwNqFkhLfNChWxHxNiDfXi7SzPxcu
BoykZuCzWbHwi6FC4pZsuN6sDXbvBQAUf/SzfAcF37v6Ux8wRLgJrQqtDqKpYcy4
iNWcAkz3oqF6pZLIxt8K0HPSq0rsedX4ktTwV3sAU3MWn9Zxcz/nEkBtdf9llk1q
hBW2b/I7oPNg/QqjaM9ChQqoM+onmlBcD7T49qdJDzJJ9BkaY2zdCxmE6Ic+fRwp
3H0CO83R2qsWaZ8zAOkJAAVy+IL0EiQL4sAPvyn4yYjGr7BYfKYGLJ6MqpKLp6Xf
kXNY3Am2p5qOdVrSsHvE/5JAQs3SIYLedeTVMrsKZ2swih8GIlfAeb5jC6T0O4Ls
JChmhNDK7NJUbft4ADSE4JB6E/WXkIu/sIPaNBOcArWJzWW0vFMHCTcQb9WZ3h4t
qryd5WnViCzVbR406W2YPf0AY7X+NeM9cSGHLnE1Lluo7TtN7SEt6n1+VgjS5T4r
q1fd9MxNmJXPK9c3BbBz7HmpQ7qYFs78j3DCrTSDzM1x/ZLSVD+cbznHmYE8goIY
w8HJIr7cchy9KI11Hd+UtJySRqhn8bh64ekifw4+k4xQWf9N0N8KMnQow/lWO+Z9
1oErOrO9vMd1nrihBIENmMhhG+SYzJzFDbs56kBm0VvfXjaaI+H/UKEF3jtk8nUw
L/jDvXCCJ7j8NfIBPNd6FrlctuL1cVJqi4UDXmkthRlmr1xCUbh5Z+Q3/ReSp0l8
lk/djWTouC0GRZ317Cm6VYjtzBZYUBsE20Xd0NH/G0d7SVdcO9ILUcBEBsepNK/e
9FFkC4x1I38aypRlsTyhrKbnEB3kA7dI3xuaYFEKhcb8mUg7sqotQ1jsoOsTpWcb
DwTvduMlYopIzpgz1NNREbaAtGrGr5vWhp3PJZuWDiTaWInTL12yp0/PJfzWxuBW
eszUrlbweIcRYtGhQ9HFrbLoU+EeuUJMxmoE4HioEDB62LQF/blzvRFcSBl8wxOc
7Fh9OE2fqaWV4kDc/Pj2z6rquiYNvdFM5DzfbamW58h6xaaaNCzULGYiTiEhIsQO
8GkhC9+QsdjVPRM5i12WL18vpsosvCuIv/4WptNH/m6/H7TklhRnaRoMbpL/+JTM
DoT13X8d1XzCVj56IrEcoJHMgYLypvKAIaYJI1bf+iaoZT+5mnEWW0GwTbHMEFMW
XfOFPCaSJsUuieqccjlrBwKDgpGrQI2CovF4/b7IkzRnZ1R+Y00L9ukPkDGgirgx
O8TpDGVVcP/+idhniMD55ujn/VCgjZE1DbqW8CSKrilpbRQZQ0EPu/pP7v44cOIf
o+2JttqbL/1omRhtZQS08FZjgfSNLHptcSVy+Q6zm/zwHDS6prHNGBfnI/xK9upA
QG7LGi4qJalxRyqNNDHg+GKJAK/+69CGj1y/BvdNFa4Ct0BaRlaA+aMjlj1Vn2/y
GRDTmHRFkLUDd4m+ENxXG46MM8vZQGZ+MBB/P3sOzJ7ARRoFPPteA2g6rdEH4jbI
b25tCO/t7XpstdwCCijprtuLkaVXLbQogTkpQFukeB+4d/XD4PDaFVLuuX3hLDtP
AcxF6R6NFSaO99MWKtdbKIEXkPIt/yLGA4VfaXKVuu1fCvfkbPODdcL0fm9p8zRr
ywYr6RrYRJCvRxXGYSu5qBq+LnPgyumOTOh3NSEF0CwfvlTR2CC/XOhq0nA58V8A
5uoxDfn3toxxOBNMuaUxFVL00LsXrLl21iyC1WBwD21Z5jAWOeVvas/A8xv69vjD
yizv3rYt/T8S0xxwEyfhOSnfJCAMGg1lUUPJ6Noa5Dm19w8VMBtoFptwK382XR3u
R4HyRZNLzAPNrw8SNLAYy46jVzQWTcphJn5uBzk1Bub6qExZ1ijDr5tROzoD8nAT
c1nCANcCw/IznsZKipQAK+egj4jG5enaYim9qz2H3oVtCAJr4Pr1729si3mcyHwj
mmcQeqhmx5bYBy6CA9BDUHZjN8ETKhsxYANf5y4tJqCKQioSSrv8Fk4cPA2WHp1T
iPb0GT6n1S+3JULCDaHj1qDX5lUcLBfUrs9/DzigRCc7SQrD8icLDJr7L+VuKXPM
0SepERfbuxkj1vfnhUSAbMj/wfMZ/2h9U4pEvnLedYuoXQj90687NyPg7behuZoz
aC6rIqFPVkARFQJUJ+YcpZYbnGlslnXm/YMlnq7SG5sHd40vtQo9jEVTkhFDyYHH
acJh0w/Ff6wL5SMKH3Ctnsyw9vblgmrjeR6xgr/mf9VsrkfLx6MpiemBfXnv2CoD
18Z5/LDrBED+QNO53pWJ0IQvHfUq56XjQNujWxDc+U4EosNxpGkqOmjeecNKnbk3
ZO/FnJxFthH3+4UHmZpsRxwUypDsFYBYRB5ViSpHfxsCUO+/Am6EKmEyK8BcmqTa
Znd0hJfgTTq7TetrJ8hjnjepjP0WZ/8KXs/YN8vXOfROca39+3aIhl8Lt0Kdpjch
huQVtlpD7bN0uL6eJ12jG0J1ExFT7gD4Hi3Ja2VCu4aO1gpHAqEdfSBG37w3OPcP
jgvdZVV+nrFDAc48NX37Zexjl43O+raG5Bih6OhOEuq6Lr/Go07BRjj2TQIeUaXK
uEmob2CBbqeOkeTtajpBP4E+vAdT+eV2Kzy0RBbCrdqzcL4+3zVvzFpTZSvp3mvs
XzOWq1Tmp01vT7QF7YgwR+2WlNkCk12bAeUqajmas39TaMdwkN9VjKU4vJaoH/8l
kzDrzuuYV87SeLcffphlpSkHgI5Ya14JGMbdT9Mj0IpU8iQ9RWZ5VydouPNX7AIO
CJmssk+/yPPBXfUrgchvrtGiYLxmprohVBpTlGZzR68pczWQf9TGr3WRXRf45OT9
byWWcoFF4S9twE1vxQGqqW5DdyIW9OsMhXf02SWgWaG1nZsOqJYd6hw9O97vIeFl
TUiRqdmEQqT2TxN6XtfOwfjKaAqUvcXE3pBGP5I5KkoAmp2wCpfiFXdkV1csAdvq
aVjm6REKXYiDArtqvcZ329V8BzUVNGQanlWrsI4BH1QVvWYWlaS2t00/+PdFf46K
nn60RLNb5x768afb0uj2T9NZam62A9c4FwXu1L+XyaTD6eoad2jSJ/k8cL8qfpAj
QgIK1hdAlWXECl3FYyUkg+ATTsZ85Hp04DBkMvfVF1zRwIoQ1wB0dBXbSHeE1ZfY
K9Pph69JOMl/jHwM1q8QNyt2ckbtl48dpKhLmmt9SUXBSO4KLlHjhrNxh/CkR4m1
78FaL163w4eaLbDuOVRAGZLugy5OPiDsHjyt+kzKtXoG+p5PlIWOLwJbzteGbK/E
A3D1sy2QVHeyYOl8URi5O2X+sav3G1uu7RYXh0QlloQ2PXjmsu9HwJrPgT1jAKML
tWLbYWxBHMA+eO96eRQHCfPpAW3MkFzRYCUBLBVw/V4toAu3kNzMicU5wssp2P1v
SJTtBCvN3OVt4mxNveYW8b0MPEandc0SMyHzXf7vzGbyEwARG12TIBqxBTt3HtQZ
Iy5bVLwL3sxGu/BsnWlkNI+NZPw7c/h1YmnrOrmTgJlle+TGRxphwX2hjBmR0Y5f
fkq6P2FyT10uYQr3Kbru6Q1EqdQfQa4ocBoR/0wZfXcsxuw6mFrnVuVFCyj1ApSj
CDm1hVwYSQDGyAD4VqIGgqsU1guzkS9/uTb73azgcK2wyueQ/jBzkkN5RaZF8cG1
iYdhFXdKI9XnSymG2qwYLJ/vJEWcXbxAhpmDm7aLNkMo9p/LDsdTCcDep9vS08tP
UAHIs84dmgpSAQiZpDRHvEyxZWzEmBWIyNsMlX/Y5ZS1WRYtA+xP8KpNScL1Zklk
NK+EWuLw0JokYCid9eHj2wJsX86+a/84cA48BcZcTdL9TjYc+HzbA9a2+Pnwag6C
aosQiB7pNHYjBheRO5dwoo7hxjHmum+/PRnxtWlyoxMZGLTbwgDdoS3ewHMR/gJF
FVsXRbJEgn5fDoXf+xazoLmQgkTv782v3OnVUl839sYveyMAod2Vr25duWfoLG8J
7lOh1E2MCK2BJpxnnlAIWKeHcEFJlfpQYq4CaHYZ6Oxy+hu+K+gFdEtBLOzqNBBR
6VmS9AeWyRAtpd/Sz7Dbwv44bP2FH/+MnDhnh5rIWL0na+tXnDBHPSmdkj01U9cN
pAIPKjwhAKu1ybZ0wjJl5mMQnpYbQtyZNJuRdDcrGczYPKhPl1mOun4w78Qp/sML
wr5aNZUfWe5ZfRf+BrTHAHS3HJClEUGH2GMbTj+rSZmBPa6xOaGClRG9i2afRYgQ
QLefmn/BVMMBCKASrq6C3GbPyDSe9L5aJMgaKvOFxVH/GO34jDyCC4aBNKg0Y6IX
PBMYCJlQkuH2VvHL3+OZALMMwWWnxQocP7zJSMocXYhrI3plu7iBapLjpoAHjI6O
G6oUM5SgylBf5t0iEaOdg4Pr2bPexorc+A/2ewDuR8VEiEFF7+zceT05JdvV2X3S
yRcZgWmOv2nlEn8TTpzVY/hEgFB7brmelyBpgBll6lG7YsBsl3PBRI366vlvQDHF
lGAYx8YmO2938bnPha/PL3PFdA+voji2etK2TW0CjFnajt24Je6+eFR2MWbONwar
N/K+V73cplW5xso/WP0M4QSrc+nJ7Mtj12IzgpVuDFAuL6vTtwppRzcCUWOq9VNQ
y1Cel/1L5QX4WNN4mpSW9hLykU/OYHRoKmvHYZz0Yy3/K1fN7haq8MAmHBpbdpT6
UOJOkVEdiSFWT7rFBkmATT7tdKqeY5lqcLaBzDhD4O+ZA1rblSxBh1K51BHt20G9
4VV6il+WtzkMo7F8MssbpX0qL9NNCzd6kl1dqlFgPJcTHLah5HAh0KRdKmb3fadb
40VSouRuh00aFRqbLanxxo5IwzXd0ZE6QbtIrez3XGSdTIskFH+j9kOhwc8bhlJa
fTcceE18KJSXWI3pmHh4cFPSFv6anEnncqb+Mb9ca8MFWiz9n+Jkga14HT35QeqC
NRW3BhoU1PPV6JnBHX9V4qjN9GNWa9QxccyHQhJOeYKhMFTyrWgzuzZFk0oxGzPe
qFd+kZFN02ajLlTa8t7aRmc8QY29c+8PvQM7mkfBO1zzn0ntYMjgmel/R33CsnBs
VNBUjOYSBSfaQQqCYlN/F0CFVUdi/F/id1Ls2v27noCJMdVH6hlSG2/NP6ANM6Z5
28a4M+dKRkfQzb1cqfBS0YYrS610xLh18PY/UeowGFMcjQWGcMRncWh/iR3n835R
0LjAm3szTuWXIlAjZ371gtRIEAzh2INuZwRhjowOuUVEl5dPfjuvTM4AwuLXlNrY
1gMcAAtjLJdKIfcoK4HHAJraUuxSZgmmswrsf6PLUBZk5vLg1mqQDNS2WtgszZFv
KDf+9CzXaJExSalgkGyJG9Y9lsm5kC/9KpC01Z7oBxTgvr6amV/VQrUYLJpZnySy
v/TdOqssemAopDJBt/te2VyOrBlc/1phHSmCdm7G+jDilGf6QbKlKujzjZg2lPAz
xxvvpO1dBhx1x1OpJWedpap5dQgEDIa4VrgN/Hp9eE0Rh+3o4VP9t1X+8OinpyEY
01eDrz9kxOiJZFt13Qe52tEecN7sBVxzlKL92Y1NJpedn1AXq0sExnCmZ+HUykAM
ZIZ2BuIrpM4y/cyE5MFKl2UzQDkS/BrFrfpal4wj2bXAllorUlY7hl+969fLbn7a
P12veZ7qjUcNgCnWTd36yFGKodHJKkiMd+VbprHsNVYNk/pmF+LKEsW299O1cQSp
Un4ZlN9czTGgH7PkAv4rWSDcqNWMVu2LCnsb523mnvrCbHMVomZHIKRFJQUVLjjY
TZRgM2g94pBB4ZoZ1ggrnDZdK0F8bQhb2vfN6OuB4bygeluzH/SrRwMlDVkxM0o3
oJCE/iM4c1DtCDU281ejN/Mkmu4o+Xt5teXH7npZqjw1hrVNddqa1Psh63c2zggY
sNBRE9S8SskAy4pW8DZVd/gMEt2L0FKWyxjAhFZ2t9HFQJrriZ3yHtMn1LuinHjT
AQMIvXVVNranbZ3v8Xwoff10AX+3cUCld7AFq5iJyP+WinOt5tJsnRjZ/OR+bLD8
sX/fySRDG3p2TXLyPvUSGTegko5C7+NEr8Ix1JyjDKanHBp72ui14vnHw9qfdyzV
2D0z4nNXDt4LlOkCvc3lO8KwJs3ygo0pzgppEsrwufdtwluL86ehsOiEfcTYQPeP
hX+2a7m9rqMlDSOV6Qq4y2n0TNyhFlIbHk0wbhOVedoMePsLpFOjyjc7bYMUPYpZ
lIBVI3UDd6Jnfh7F2P5115W99myetUapShp9Pdr7Z1xMJWPF0fFSz9dZXyTD216A
F8PNcim0fdISFuI8J3zmfre/LBPalWKIQ2S8s8aO8h7wAzpI3Z9jNa66BoGuAAC9
llAbFzdZa70N7q7s79+OtnbMNaVV8Rc18JfDuf+TPsTPZgxy15cPYsQSO4HOr2MR
yKXBDRh8vInWORDsx0X1nqcxRYtF7vMUU3WsFXT/VunlFzj5PcbdU1FcYrgIZMup
txG9AzTPzhb3huhToICHIsk+q1jNALsJMtjU6Yr3RY9KsIuhbWkC9tWGkE1XRvkd
kLaW+ngEI2502TEXcMw8vF3iNElKeixovqgMH8Vpl9rWt5GuPr67ymuR8Wndug4K
NTFai+0fDr74L7bppZyz1s/zyK5OJUQfgnSFiXAbC+jR0aE1NECNzpyZ0chqtr47
vMysP6r0PPy6h3dBsBjCHVEooVL88jha9fL6aRpB1btl7Ddj5zGvrDLTnSSHPhc8
9n1PvAYLcE4clxsUU8trjgC7e1NEPrVqG4ZhGNuhxGUgwFlGuQTqTi8SRDaeMLvT
ydlbDQydB0IWpRegBXrAjK3zPYIBEBnzKnrjqn87tByThQAZ2bRPLuL5e8qEs+ca
MFYXZVGQpDX0+8a03Ml1pEK+/S2dB8UNGtddg1eYzI+C+0QsXBBuauvh70Fo8d1d
70uidaJClDoyI7pMdtSLsDcPnD9ySRnuffKn7kzUZDUVe1I/Nw3pJA9c892BLLku
9MPwmm9dMR9jnJdC4/z2Zfrz+l6ssolAw9ubbVKkCGrv3ESsU6yx8DyH217Gfdmr
iEqN5Qv585ckhZ9/EAuABBn8MOPWSzXZR3mstPHRyXMtW6k5QgHSfGKd239oPHwr
QqIUapjM0EgfD2iO2X7EFbMpqFcg6atx4omyKGRRMyZr0ELKHroZ0cwQ/kqHVZ9A
G5y5yAvmVw6STiDoPuy+LNceoHq9MpyEovlO2yJiOU8r8Ka03m9q3XvLkgWGg5Tq
6Z1leVdG9veIeLoOfSkzbj7oeWSb2InUMuM0Z/hHGU4w+/fGFRp8brgxwKeW1ajv
mJ99oOJMBkJF3ZX1Ut/LsiLbVOc410Ru6xgAd1zf6BYi56xLKHFF15TWFbn6kFpu
Nc79eyKJaI8jJ1EquWiIaY4zWMU2nfUkxnP0IVNPc2Og/ygFSiqG6eodqM5ICrjK
Q89wbTSe1yIX0s2YuuByL9T8iuzSHk01fvNJIuxd6ACqo9IFbu4MgThnQbcbCQ86
fNp4mr/cZjMDLlKkuNpa/vs1ldK/7CrurJZv4iX7HlULjs+JutxbqW4xUnOP9uWr
unhm1YfqQz5dIRklui4i2N2vBrrtWj5HNBV6lCi35fEyrUub2byHz43bQ5YqFS/B
6xhZ/VdyZEQkGSHiwy7JSJB2WNaFNkWL+Pk6qYzjJpAPHpOgrp0ukLH8BoT274nA
S4CvtLfp3n5tzt/OiB3Md6avQArIsqwVqkMcafStkYw6CV/EMGHP7DhvKREHntHR
CFPysS1vZsLx01uSMGHgzWkPooMyu2YsHhnJqDdnHC6n3CYEBxV7lwODRkrD4ktR
naMsjpslhUxGOoj01lPyIyzPWYOEqLwyyGR9MTjv52kK36eVt8p4EteCjObFJ6P/
jLm6Kf+ZYKvySAb31Mz+pTis7EgaoTgHUSoAKVjnQ0uWUDMU8PyOL0U0fdYJO0lI
qc7fexsKZLaGRbZ8GBiNjYZ0K3myq0ZzTGjfdKuyWtyomyDMYAzW2ntrq2Qw/e1M
MyGFO1YpBKcrSYgOES5s0mHBeJjD0AJMvH7iACDT9jupP1oz4e8Ni4SzXMapKb5D
88S+80s2xb9zF9RZqPvQoJ+himgbmCWoAQEm3ZIkA0gmZbIKmx2FxhX8IHH+lwBc
GjBD7RXeibnTg1SWkkKtQ+WP+Wb09NbMM0249vtEiZcIkxw/wXD4AD16SKBM0+QL
Z/bshoWIXZrtr/ggPpY8saYJdlsLxiS2d4E8iwcxSeOtx/ZnOFuoe/j6rqcLvFNX
34vrF+EZWoUgVIVKVy/Su3do6bSXoLPQcSF3VyHL3rhLnNpNj1Y0CSvJTf6diN8c
tEqNgB0+BCPnDSGMrtlJ39JKlr4DZSvPri6809M4HaHlgIL61LFNo2/YyI6UCRnW
UwkAdUmg9y8kFxuOLXZ55VxaKxkxG40S9hvwLhuG4pRuoUmRM14ohv7lGC1f/MrV
yixX5n3OsP+EzKJCSnk+FKG8V+EGf6TDkGNGibXXAgqG+b2UUn/P1kjMOetGoLzo
vnfgcADOtGJNEWs9DkM+pE/TCWQnaTjJBHAVeVfzL4H+ruDw9jgqluWvLhXM2w+0
1Wbe2Pp2LhA7lQSAUsA9PJUh9H2L1K1CP8i2quhrZ9gQ6FhHGG9mONVtxq5Ofv3i
TjaQEZOWqPldpzCToH7FzeXb+RtZpq1GOLusRXMESn1LYEPbyZMDJC4tIWbXRpZO
BjRjJ4Od3Qgy94MeCdjVq9Nrw9KWxQ+dcORNtFlDxVJRziGSKpOcZP9otAshxoPa
KyYvUysa7ZJm3q4aBKj+zFbOkrKtE8OhlEf6Al9bPEqhDioLCPIiu6oXssgBV/Cm
oUkKL0zShFy9gi76u94Bb9P7MGwOTX3eU8lCGl8zvjSeji6I/idD1eWq9gCat6/U
lQUAlBeKrXwMn2Dnj6teMM8SMpNHZBd+vBh30D8DHPqqC/BfMDDWQg4o7ddbjg6+
rYwP+RI+Rad4pebhcPxbBIrxAjNU1yHw/a9UA0HK4pf86FKbZ3vBr0xWAqLwJB++
RQVQwEZ9iWwtQlRg7NhegGAWawj2Rzis1ZUOYcud9angSvniS7E6W90Rv8033ADD
BZyp9d3iSHGhZeQ0JLI82t+64usiVDL2esc5m5KWgjbRdxi7D1AcFEs/2bZPN78u
UPzHz1hCTObX/4X0CjNGGMKxOyQS4dVv2BP8m+gJ+xFPmz3RR77rTvcmM7jzpcfA
Rc279ft8YTvpLs0r9b7NPPm5fr1D4hv3olqoYhGF1VdjNvI9uHwUoAyMmIFvTPsx
KC4/UMSGwgeRZqV2arN+zDBMo0VD1R3JH6lFZ2n4GmVgPcfmYEFsfORV5x/Brtai
dIzrdh7xxNxOfSxe8VDFJ6aSkp9HC00orVQRbFjvZBgYu0mFZfrLEq4Mov1r+ULs
ngkzsqZnIjRaRPm15UrQYmGWFqaSdCtE5y2+U0Wc12gwGP30iyKJ1REj2mQOKPor
Ele3ScgY0KbpOqoLSWnMUXqcQnctRbitVoOPkgfHCow7Wge6qxzeKXYNgmL+mU3+
eZt8UwRxn0aNoFRcxXuakqguShsqtm2fUKOZFKDWpmxF9cMoD9doGnTH/0C7R8Fs
Pyc0eRv3B63glXwv8s7DJucGNGMTzINIK/39eobt8FuDRmMA02+XfAg7/9xweaiy
sjk4M8EwVqqsJC1+lBK3Ebexybj55I3wRUaRvs8nba0Zct5HPwWwOJeAz3v+8zS6
hN0mZ/RQzTzq3fPuWC2kLK1524LNwFlfgY5IJGOUeCXOWtJZfKWXGq2MiDBWw0yO
M3Owab3oYx5urqmJXuiXCUylaLD28kipjRUnIi6Es3qUaWvbyHlyl+VoL/hMF8aS
WXB6JFJRuvgjCg8o6QtfG9XQ/EVhMEjVAnoAYZ77n85m4p1IXxjHqle0oZRQO37M
kI1nutIJph5sTSdaq65AqWkZxRlSSpT86LsFAIwb9piHPijvg3iN8J2sl3AiSY0+
ga9kpnSCzAR74RA/8Nk6CzrFMAiz8TFBVOk41u/Jvz2LEGYOsnWnzx0x7rrVLNq7
uRQ5X8ajCgdDcWnTV02LiLiigsC//YNKqEajuuvPBYYF/GliwsFncJGAsvnW14/T
WzPHdCA6Z0LQVtEpaqAVtHUmUoRim1mVMp2VUYdswZfk7K10LtRjDAtX4+yVODH0
IilVEJbIgjxZaVrKX0Xupquw1QosV8zqNAgff9HxBzRSODWzjw2dZurys9423Hif
y7iQtLbSte2nq7TJjmPbOE+UFFxNafQEUaGhWziiHiynzCOg+Cpd+GO3P7mO1Qtc
rwiI2PuT43V52zXhX1RorUtHiGw1tItzT5PqhGYO2KZ21PJHPQEuJ+1Zdh59y3d8
NL6unHT82qeyy26k0PiBT2pk9vtFN0Jlw5FMA3ML1Z6yBvSeJc9g9/S39b0m2SXb
8OA9dcM3BeOj0eG2b94xfLr0Y4r+sKx/XKckTAyPYxAh7dD47UTtv4djOzwxSHuN
pnYbMheNs/MzESi95SY78gYGuyoIjsqLr+rUhJeF5Gc5TFgMlXrVrx6bE+BuDpHm
LO6DwpwA0OY1chYpKY/6iD4/OlLO6nUT7tvc1q0xjDWtzd1DWIs4mzZbIRccuBpg
Ikj/jAAZeM8Ss77QM4ZW/hEuNGMAJ3HJLnKIANAwBJ18fFRDNtONg7E3iLVna6ph
0i2XCdFeNHZHedN/uPoaTNuMStlfiqlCjyWPs+T+usfIBMnWyvRzmBV/zC2THehf
JBOZcwhe64q4sK21cxnXL+ENZ6RN7G8mf6vf7f2TD3uoOjplf0uwpJDlsMTm2w2p
8hPHpA445FgaHnY5zlCRo+1Qy7NAhFubw3F+1yR2Yn4uIoGdOakbOzpejppm9Hsg
xUjyQiVg/MijxWAQG12+mhYy2Aef9BCywsy1wlbNHFtT3LtaFtjwQWwxTATC4xas
tRQGKKrXDrgGESx3qzc+X0hngbkj/0K5skoR3VYzps+MHNkbkKQR2poSAAqqHdX+
BoNCLLTTfw5NN49XiYhx6AFtJqFLax0VBIqGD2YVFmb1o67P3xzHBGhrLI25Y5na
UHsapTf2JfCZvB/3+NABsrj89pWo9878+r4Zjt9DbFUSeQEYcOzsLIjnclcbUSCT
IhwbFwO7Yk8CBjib2q8Ml+BbpM63NHDMH9pull7SzbCpzuqp/rQB3yagaLCSi2N7
imeuylsZKmCfAb9FaGjMtyyolWalLeQXcRvuQdoIvAkVmoczdSio+3dUl55ZkK6C
SIrjwV4tttZnYLXRVEeBU8BP4Z8dwAcsrtSwT2KPW90v83OvmjKdqRN1G8sG+YV8
m8uLEMWClrrcqJsuIQbMAb79EcLhMkgSCvjS7QtDFuK1drPKmx8tLCjajdactebA
DmZUCoq/6hBPJB4pza6LrGvm5baQkKor7xVY3v5A/diarb7YUvNdVIRIAqgVQ1it
F0eIuQ2/B1v3QKQOf79q8eHtndcpAHcBNeaeCsOZJtAF4zqXh8zNsDRK33o0dKsI
+JHEU9XzY0AM+VgB0Icy1OMwErxNo+ZZj0fAGZwveUPh0JjhuZwZxo3mmWVdnz0g
lCY0uWaEMa1UiY5g15ELTTypPPjUqlNqOHEImwTNAbyQimY56xauI+44MCpNPjiV
9QlKoVIPRlXOpN50rNtWUA+CqccSEqRSurTbFAarZRC9vA+9QqXcId9n/4qUA6hd
+303SUyYe218GFEhxxSV0xr/AyTlhzv8P7UYQUM1SVihMZERp3Klfp8vqqYf0vey
MKxWLVBDh75B6SJDAJKoFX2PCBO87TcDIMISZHDU9ukIT7zRszqxVH+6OrejmjJZ
iVIh9prnzoF7v19/fixmEHB8UuKd2WpNtKjWq+yLwsB1VJCKeTZR4fvJhdFGjq0T
WR4U9vN0gEoeb5gdVio5jyqI65Fc6UI81qyrvTfgLx6tLbQRBvZnaEBJvuRpZSRz
y1SpNLvg3sAMRuQl3xAodlDB6GML4XdWdY07zBLSjOtC5sF2w+Bnir2AjsiKJG1B
J79+Qccs8O9rcGsFNqJFTzg/47M7GJcw0xSvwgiP9bG/n+d7K9b2u5iUBDJ4MNFK
UA7zBjNYAMzfQa979n+/NNe60rV4P/v0A8mc5PrzT0HHM684RsZKEugmaFssDI58
Yya9QGpxz0qLekc6C9WOcDZtPhhroEiCM1KcqLFERjmxv5VCa/L8mobIICBoX75C
iTeZb5uc0teuKfst1U16Jum5mZYGM1DGmeQeZvT7YSEqn/oCseUcOn28wujkLCH6
1eW5Z3JvtLjzurlcQQbnGjKXKx5fvzAvkcD9uiNKFIrYeGeAZdS4uttGpt1fPAgz
E0kL4K6NRkRy/OGlp1xsplBBF+slx3HcvNeW6JGrroLRRV/SKU4NC4gf7dXLZ+Gd
qYD1bvoMfFGlJDiwHpz9rZCreroO1Mqaw+3IPjKqqpVIaeUefzZhCO0g2Gwsa9hs
0F0ZvymiuXo9OotIcvvVE6XY4ub0/dCU3lWf/fUFn7cpgqWPkm78JN3HH8TOKpJn
kktb1MiiwtrdltoRsbbYE6fNRlLph1X1TlEwPXEAuaOiODo7GB36hMgvOdM0O4ja
0J7zOdyyhVRi0I20nCIHWTRSSELJd/gMUUVAiXSs2nPVOca1P/VBHLkCRS2HqK1n
sIfkxfvIumfvZsrMH90OO2ksdpeMcwjuomo7VMq8fe48/uaBqPu99pWsZVh8H7/m
bMaC12rl+gyqG/HrxjlM+cKoh0vo6wgoWGYuSSUowcell8HwsknuhKW/mkRhfFUK
6PDnvuFNDHcd0Id75KYD06mr/tTCh8H/GoAz+uyMFwvZbTjYOPsp4pxnL5tByPa6
QCVc0UxqUf1R/eehULdVYoE1Mmls4qNcbZHvoUfaaTbr4FwvU4uiTZe/HyPld3nZ
2IjT8RAJrOXNWqM0mCs7nNqpekJ8l/DskzOSNl0x+VYgaL1HmMB6FfSJDfg4VfFC
WbJMr+5t0HQdzILrpQ2L6je7SQn7rzCP1mhc9Jd3X9AcVKLKskWt6UJCDkVtub2C
0a9weM1R00uDpAYfdO+5c60N3rasrp4QfGcnKHWL1+3D0fttBC2sN+q32RvnEVvN
W1XV8uXcnFl5PSRqHg6GkXk+ZaVGGHi4l0WLY+H7/ra7+B33gwoFSmLz2GNDEiGg
N+RU92hD4nCmwqEYOpqwRLTWtyinSSLmYvS/aUiJ/JSxHKU2EdPDFamS2QzcVfYI
5HVcx1OEK3WjYqizsDKHZmvm5StD2FgElCXjwemp70Fe4vusOLlyF07GSAkFp61G
I3HabTusiofY8iTxHhsiR7wbEvJjekgJUVj3+fnM7YufyBKGowpbvw7mdzaxoiIV
AKimuDBVNpbKKYiN+fqgC36jOZax9YcLDaCB1TT4eT/W4kxJmhGRRD2oabG32K0F
ZAk6wuE8glWwiTMLjAPoagP++AQ+6gNh35mlTFcfsNH3q12A2LUoeFHt43UUe2Um
HzhVL6z4cqTqJyKXtgYlBIDqLR2HKVAA1tDGmOvq+vCMN0u0h9ZZdM3W+pke6wG5
RtXieZeC0spMM9olGkQV4JEwEmKAwI4S5S2MEGpGIAMCT/J2lTKl+r/ynh/IbNTu
wbDDFYVIu/s1UYPm1mioEd0H+U2ihv+Ai7QKJfWiADmVDA8VF05GSZ6okgQT/xXM
sKBdbpiDQOdS6Ue7+Mb4g46e/aEATj1+rzpMKpLc0or6mIQwbKvGNLBYN9PfBGP1
pMVG5EsMlIN81ajPEnIPHi8xZOidneKf7sXJOnloe6XFINH4RnD6Ui9azkXBbHkA
nq1ZfTcyIKqJ56FsqqAZuln8NVWTpIkR0JSvBRTz07+8sglswBn8lKy0qwTqwpnZ
CnzsqxCbeErYaLrOhmdO09L+u1AT6rXY2qrPtunDwF2BVsm4FfPXo3QcpI7+pFzU
XLk9xhKTnrVoRd1QsOuqh/nHpBoDneDKk1JDlS2PNtoImXIHC/uXyuMC7xWbxuda
YErE5fRfpQL7g59+eBbGmtuWa2lMgB2KCxxthb63IrMcSUo6am/q+hr+Fvho6cHm
nvpbM2QoTcPn2TfYaocnT0MjKo8sfkZ1CUjRUOOuqni4gsxW/GsKmNUSpLklkiO6
jwXJoAMdHq1sIxDnFv8ubv5uQuEzibXr9FsCpUKzx2WpU6mtJ4wiWcxpUCSp23gu
sY42EfdiRdNkYOM+lUlxH8kBj+Zd1954OyQCZPKJY1ufJx08/XaUG8J4+2n5dcOl
aRmx6tHkZKmGBFOZ2aO3e5Whpu/Ix3DnGTXf3QdXk6hisj0RC4GSMFmOvhsv/5dh
iyhKJvXUcYohTKmAtcF7chL9NNWeI6SaU0MQWcWnnjPTHov8v2+HBkOFgDWLvuXY
dtWDlbjjpQ1S1rBLdrFRzL5LZFwn8H9+wsRg9lzaWrYsgzZiTFVseo82+TPoXSBn
mdAJwU+aML1GWo4O9CbNHg+q4IUSOX1CLZZ4gLsOFb6f6aSd8MfmID+rkfi2+Fxl
epz+BlnWabWgQSmbv3AT/oWsCj8NMy5i/lTYNTphHO/zuDuJbIW50FUuh1rlk7bH
Ndc3+5FByYuKqqifFcsfmzeaKg+2q1WkHf2EePOg1cvRptvIbZzZx9Y7B4cnvdHA
skJMAaZRpIBGeO+BRh/ZquOMrWp5PuUlWdd9LNVKPz8H/WYRCNufFNIEVG/4EvNC
4BRkQYeMehB+NRkSjYdUHAmgNCTDaHKXKuKk6KrmpnsngY77pgttx3q72IPooMLs
db89gD/vV/Fjt/4QZ2xujiDzlFHuWYhgQz98P3NFvAT9bQlQvC/uVSk2C1bMBry1
V7nyfdkM2v5C3bQlpWATyAFj2HpACeuNw1Qlc/+zmp4AtlXeOCeEjcOqouzeWZ7i
B+CS8wMDikIxrSjRkQQeCEeFxv2/95SX1KJzVPzOnCFMgBpPnRtblrS6WztaMXWg
j7SQDpEGBjjcNUGVgr1WIQrbWbS38O/8Kw/PswT4DopAXWfrUAORbfURCmxnGOr5
+2FGq+KZhe8V3VZw4+M6oNbLuNopRmWxApQ2/wcgp7kQ4pgfT917gCdKPTKVCOm5
3v4xIXQ7Xp40Xh6MX4457gf3l2JiDqhVrvGi8AGr5i/LYlQoHYCAQsvloDVIetvm
qP3WRNQ4AczI3wGt1kJyX3PqY4DJTW+f05vHdHrgd5MBsVOoSbxOZgMxC75BGkxw
0nFb3LufraFoIrsGGxwQpwb6ictyTBZiy7+EI6Xnx1bbRv3ePRS3452M/ADa0LNr
Fh56MGPj5ACT21fUEoHGrN2eGHTkCBbvg/VLh8a/tuRnjtRa4FRwRySI54A+a7Q+
OG1BQCAclvaGstVmcmpgPHdrSPw5q0arPLEtT7Oq1ZD4VMXxyNShuStV7tYAFQ7i
egC3wwKk4TELRIIAFpjjwKyG9h3kjHRU2asnvsHwji+uP5Z0uIgm12Crr0Za7LcX
YBIoQefx/brJNwSUAjIPmyxtI0RIobTPpU4t7ISAsX3eexSsvJx7WexmXuiZ0DZb
mcTlVbMjEeXLUBlN2BX2feSkSESFaA4RK97pDHdVS9dvEBckv2Zlvcvj34NzITlF
oJb5ZwYhz8GYbNfabkKiP7lnEdxdmH5PyNYXzmw9xsi9+gBt6RViERjALyORwbUw
shv3ulZeHmjFuNs9Ua/YzonBy+kCgrtkHeq+v3N3m5DkGNDhuCZR1ZmhSQHtP5DI
lm/Lwaju7b+UGv6SuNNQ0f+6VLkG3d/adMW8PYQ/BxS5iY6dn8I/8QxcZ+irbKow
X+bFMdcMPqdS+/z8SgzQmkbZiKfmYLxVoqP4jtHJP+PaW+Igv+HFKkaGwIwlQFqI
jAdlmhnLKzJtRh1aoT6Goxgxewpa2Fm04WEE2/6yY9zy6OQwCW5lxTL0bsO4bDF7
Y4IvF2HjaGdRq0qE5B4brMhRZGh6DVtumK0B2z3W0z+BJyRtuCkTizDRzJzOzUC/
CurlF/bsjsJYd6Uj1cvEf2eXrZENgjrn3qBipYSgCrkL1RLuVKF/D9NEyivhAxwM
PYyoPA5YUCHlEdXfEHZy4NKG6Di0eKmSqMdkubzgXZLqwapS3KnSUquyDUO4WQuA
GqLZ5QyEMTp8U+i7js4C1PA3ZCdmAqEir7BjnQ8pqCH6O0wQNvY6bXLRv2JI/erg
r4X2MntV9SbCXGyYO46/3OvFrj/Wp5jBWv218gkM0KkDRO+d+lqTuaJLYZphhSpe
gTO7Jr+6rTCzmFzLMf+Ly0Lk9rMJsuFrFiC8djygR+w12sfCsgSCU/ZzKWWoRhjq
HnPMzIU0XmxYD6fU8D0ZY2uw1rF9Ooe+pYVccHYZMpMlqSS1009HKNcM01cZDl7E
4UNODSpEPTJmE8axwL1EhNjQmD2B12lcl26AbUV9Jp3YwzYTmHBU4NoxKFbqOfFG
Tnw7GoE5qNtHw9yGO7C2Fjv8/vjQUIcgdkGuflgww//AbqaXttBFewtmi+GuC0gj
qvx4YS01wfzECICLfSz7LdCQMdjSudnWKew5yV0yfHUNbZw/3XsIWabcBVfY5Xbg
IgdOeFSrlEBd84uCJkg6g43Wb4ognK6yQd4lvINpxHcXsY8SBWmNzGGqvEeCTrXf
IDFSJQ4Tk9CMgo5xItbCLlBKUlVZbCKEk7dCMUjXLCx9E9LkjEkoez7VB3zMsFB+
WCErksP6ATnIKpdBt3Y3+Su91ROJtXkMfRAjhSrWxMuZ+ym3JYtICKH5+ZIsDdeq
XoMqcfA7D4VJk1Zt5LMDC6UpZdzQyaqzsjjheejTFPLzlCd7kGurQyPBDbeU+kxF
wxgneIZKzcNv+yH4r54O69Qox34VJvCT6mAZG9KJK6llK+u6vbRyCP84TQcY/I8w
6Hc6Ta7V2OG+YOBhZrdR1BDX8umHEGlsLftlmgvCm5M+PJOeEadNCza9gZVzzROv
V6LJiYLiHKu0KfTKgc2bI3SCdWyDRdkSD/fncGWtXH5kW7owczzTVcnZeI6ply7j
2zuzhPbMQk41xfPMpEYjZxQJQEvF9Hn2QY2+5CGcAJL+DdULI8CJoQK4DdWH8/1b
UhK1F82phFOykiH+whSNUccl3T0Ig/vC0k2BvAJFPLkK0hpHtkDEzMSeB4xrcYee
JxBfcKGWVtSDRyEITxB03wfwSIxddh4xhtu8590V9to8PAUwkfWZtRjCkskldEET
c/5qj/H/NWtbffpCBvWTvOZu+RIk4fdkrnELZ07Qv9Y+F/POnmDKIgvikhQ5ev8F
tVEbySPYfbyl6HTtQoK7fkiUyhIo3CzUnAJO5nIqpRV9NLnswmEM3pqenZg5hqTu
MkXRzt2gzgb6FZEKc6sorOnk0g24EZdXnMZxC8lIwthwUlWvGERlHDuO7wbIV2ER
Ze+PP7hdekFrgFq31gWeQxJASpaeVT/wRS5cQRok9FIa+MdObvVyA4PLIWuBu58D
ASWuwmPsPHHAEbBHN0oaP9vdY4oqDqBCQ54O2U9DgojPIhPIEvA9lBTLbs0yBUai
NIhJ33U3mQ+b1Ij+UrS8AFXBiMWyzKlNYRUtDmZ6BJN0fqGPpWz0ba6GcKe9GHvT
BCKk/XEEAIpf1YSNkUnwJfPUwLhngQbtOveCZlWMsfcdK3QP8Th3dx1x4XIkK9Pi
bggceYS4DA4a/NP5GXLVcmgqHWkKJ18tswv6GacjJ3SqjzhteXj+sdQAfXwQ/nsH
Y9xGnHlpsMQnEiYKkcIyTR13jNHTtWBavK49Q9cZ+Dsh+tp8zP2T7OUQ+23SU12a
uD1T8POJWA2OTr5QUx7FmEb+nmUuPAlYjvGnnjwS+2gHpKJ9+JHaxXk6S7qFlNnY
pH9FyDMoPpSoAUxY8q9yr3JtQUk6LUDoRY87mVTrxXuxhHWGekXZaKD+qxtuCiJz
Q++PlMtG/pbgCs9DZy8i8WbyM8/n55oeEAsmYYnDFvxVTR6aEXYNnQ3XFte150pw
2lQG8BFzl4/VKCFilgOaxQ8gqIYnMupHY1XOYV/xFI5zOT+y/eUsHUnJROMmc/Ts
CmBKrLmAI8BZDy7MwwfWRMV0sKP8SprpQi0MNE039odnfZx4Oyf/trRqdSmLPnew
g38genc0jAHf2GOi0UKynCu2VOHXXdHP+9liRO830M9vJn5nnPUXZ03W7UxA17yV
2rvCK1Hx2Ynfe/2b/Zba2S1fxc0iZcTyfXP1ZtpUeMlUNThJacIS9jYIAC+sXy/7
2ZGtQpn3ZOyYxhWUo/mXL8OKHJ/i2uQN9joi+JRDVyOi0cNLL5uEDyt99O9Z8Wvr
CzjsWIMTg4pgEk8gWsdDRA7sTAa/OkKrEPidK3cMFD9JrhyJoa0AkB4ydnZavJUM
lQQi+JWzp9bCA4d1/aFgRRf6iEwxe8kjUDh5ZdX7JD1HxcnwsCljvscZjUC4n/g8
arF9IJGo+pQBTIeK4+aJ6l6ipmbeBlCZq3PYLejqEvpybLErVt2ikEjCyatVSOQi
ESV8C2NmuTo7Mw+leWU4PFRGk1EAeoUITt05GvLazyeBhRNZu2KLZ0UmJ9dvUm8C
Ku0Th4ap1QPbwa97ZCLTHilwORSaetzOTEuo3KQ2rRnBQGggqFBYb3xwkFDWSoVq
+HOku0Vxslzf+2HNwJMYKcfEW6vx1TPa5/iJg4yZDVI4Cl9E8EID4Qjqt8UH+9mc
EiDg26QvAf2fMmpq2SnTtHA6VQ8Q58vtUwszyUEONGLT9L7HtDf1igmbjuHiu/6r
5TePvkDQCHSokGFedT+bxeAuAK3CP+IV90H1IWrbt/kmhUIKAH2OMArO15IALQNP
SCoEe4Pwqm29CgKgVU+EMtjkrFWtHli548/maxU04Xj0m+H3OF0sqeKPDTrfCffu
latEFmqfoKQ5uzSRDWWOC8Kxu3VdQGqvmB6hihOQEV5OKBdmXjYyI7f8jSJc88y9
fW3YbQ54K1r3fg7X9pZv+VRZjz2S88IC8XDaZgcMp5BCk+z/ltmKqfpdRlTx0bo1
+7h36Mh3hA7Hsij1fjz7Kx6o/pHFLaHFXr0zFyFZ5zK8/0H6z6o9Rquum1XC83nU
1Wm6VJlQjgCVHG1zzzSqvaK1eDrPm5mM4XhLx1TgMpOH1qwCTibS2/sHdM/vOsXX
pvw5AmJNJ8Cou2fmKvrAdyZg1+XydeUrEOXgfgIdWr/KkgJRgQFTfNthgH5Q+pOD
3G+rhySJ6MAaMfqGMdM5Pq5piJaJxo++R+HtC7SIN10kdNE8ib9aehArZthyncgP
mVQsL4oj3WuLSYnYKOgvDI02QK89g6g/8b6Oqt3VswINoiF/+R+ALqSLrQR5m7P2
KFS+PvAAaemmNkCWOK5ihEZXGK5628CY5VZ5M07HQuAAQmYOzjfe1EvBIIyRgji5
9ghmeX8jU8acTncYEOtt+cvdFiuom5hOwOMwhawZKZ9IL72fFwEakSRO7sEoAYPd
9WTW9DMj4vToYeDGrmYMIc6FUiK+PV8Y7wU/fZ5VKsgGWwuNjvAGdqaelFd4G7dQ
09NbhfydrwyHSTznay+W7PxD2XX0fmL/2ZYSMWUhDfqvv7V6qH60cjvtqVEbGeaC
bbpQUJ8gPuNUbj+NxmFwa7c8QfcAsgvcJj4/gOGYBBufDKFFEHyGp3ba3kUb3pn4
i4c2OVX52Aq+zOv5VRLPe6ApOI4lsRfYda7oJ43DUNN8Y2H06kyia27GZ84/Dljy
YNof2rc0JqQzOmBl3QOM4JO5xjy+uCeWxA9vfPwezYqtjsmr47WAfYdVmr2+ojA/
tpbAZUheHaSR8LytI1Rh6CFgbgQI9oFzL060gxi3HdLJHBfDd2ru41kH1vkYMBXP
yxIW1DrG8rZTbkuFkfbcajD8W3qVVl6EmTGQ5XymVHSulTACeWR7FEuyAXnuvaNg
HrbiTZPbUtqS98ZDMTQ2V26WaiFAO1F8n5Fey9YVj3e3GBSVRZTY8/AHWD6Z9HWw
iGNm+dsL+o8ldyLh4Al6eomlp7mER2RDB7P9sEIK+FK925iHwZ8ve82BTxDGlX+H
ZPb3z1iV/F+vEL8VUipZ4cAjYs10wN1aTacAbakF0uMmeif0C3iuQHATPKFgxdLL
181AgJ6ppM2MM/H/qTBS8HfmYp8rz8OZzbH088arav319geI49K8fgQhkL3G1Nsm
12Ogh9l0u7Rno0yat02xJQjqhA8LwxNlor7kkmjTSh4oE6dSNtW72JPrNakOIy8u
T43lXQ3io6BPp0eN85YtFZRqekOMFv+yhepuca/IYBY5kRgG/4ajN/cZyYiLOqUy
ftPLcSuh/hWrKeFaRpQI4ie98xFppe+iSJifkjW23GzW7MaJE1Glw7GOLFbqnIaW
AIa8+sddvY2v7/E/1Z1eGEZWVpraq6J6J+QPa7i9rHO1jzxzRrwZa2rcOVbydpWQ
Dwy/IZeWbz2DseXKg6nJdNNUA5Zuo8sX1OeFzZcyIIYrETkPaEPbrFbqsXT5TK3z
phNyADxaTwaJNCPhrQD0SaGyUmJOB0FsMyXef/mBNRuUw0sA3itb8aTaapmRaG5C
MOuNsVsHrbDWLRp2WL/gPYLPsebG9Skkqr7/4qIlZTCAtU/MZtIf34l/Mo9RHMJE
dWw5isBOsgBYwEV0tGOks7Kj63CvWPuLDQP4Qk38oV0gNMEWE8RSU9YV2+wY/IH5
3d3gaDoFTgJI/9E4VTahxqa2fTbJdixrjZ2j4QwuIJBkOqxfqMDh9XcsKHfSYotV
4hd3GjYY4vYGQ/hRLlLKiwhNhHEhWoZ7ySV1/sPX5jJf5+oFv1SeP27GNPDHUOUw
UvGw8zrw5wnAcn0vF+yuwmssL+2WqCibl1Hd0QTCv5aI8Lk51ANUs/euozKq6m2v
tJlKS5ZlhD9nGgReJKQTDADNg1UURvlw9yvfZG/XhIJhYPB/DX4QU7Y+takVocEt
xKo+Yw/c7P3Ucr7dQhI7P2WkLOvpjrPaMP63O2E1/JXcM5RPpuY8AYthtPqySHAS
dTpcj200BbGTbed6OKYC74gGzofkhjs2CBjHrcZLhedscf5kynBsvtnJO3cu5RCU
EUAIUxnoL1px5hGcMG86EtuJjASQfo8SaQR4wj6pjKzvEzIumTmDhoLzi0Ou5SW+
6PwFWjuACVrEjt48bdD9174PdmMx9Uacg3jStKFBrMejsldbiYQejy9JqigBp4N0
LIcV5VekQ5nzsXtQex3XN/T93pj343sPyhBEDEvHiaH7nfbaKMpBIZP+yc/b294e
2aNGl4QhxrMLeYuh7ZDOuWBybBbdDROkxq9/J1GEyD5yuAvQh/oAayjjYhNS+XbE
5Lxty7EpTCIUgvsPGejZPOypaF7Wi313KiXaSpuDVItkGJIdWddgrMNPhWnnVi/q
vZPrzOJy3ws1ArrET1BCtN0eY5PjkyaHKvEYjYw6RlD7kHkBrJynxceHzwxlOFwe
`pragma protect end_protected
