// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:37:12 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
AACWDcspkfiuhcnNq+rKgLpwO5rQZE5YtJKFPwEgTeeuwr2/0o+mucKNCRz0Z05R
eSRYVITdzbd0uBIGJXwqyAc7qjtk3qnjGOJfAy0KQ3N/YTbGJZ2TydxKxPnhiCo8
0a6GAzgl9g0nOjG1Q2vPHSbhKFwok+uY4Q6x0RyO5gI=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 13632)
hUNk5LsRmXFz0+mVcD61KDZOJvlSsb4BtFPjo8TcHJxVMWcifY73FEdB9Yhcp+1r
bv/0FxvyZbZuPteX68qKOD+iC1eUnug2TBwst+acFHFf0WPeco3uv/SpdZPi69FF
ctH9mYZH6z0lkKMoL/vY0A4S4aYrH7OBZhyjx4TMlgnaNss3wB54kUxR0t8MejTy
sqTxQZUsQpkw5m25b14C+hTAsYpNK8cbdDL+eeJ/l5iSNPgPPJ8iiHF/d54Hb0iL
tWx8RQGOR+tXr/Rau7uV/0/wKOtUbav56CZiDWDnYhBr6ZAakrmICCua3k+nU1V2
W44iQem9+A7Yd7vBqiqi3ONyHe/bVDt+RIlLc4rX1cX+6qkN3y+M+EwV4O33e8P1
QazrcPxYsyDrv/6Gn/dleZtG3H55nY1WlIliks1OLF02dIEdmsGspe6j8mTF0efd
Lr1HCKFYM+8tnBDTKrP3p0HwIG+VFis8iNtOul2BJZWdP240tOGtlIIPt2SCIO0j
LwKm4yNrx5i1rwt/rVrjj9fS/bTF+PEmfwk3gKyKia3KHob0/a/SHKASbuhX6ePX
k15KMBOjbpw0l2/RdyKjusTlZVeVUM6R6rZNGhDW6Z3TRmEy7+nUlMZGl4kgK4sg
C/TsdKNBQ8g+SanTfvTk3V+yiHE3jWLumzUNpOk1Nc8dEbGxoMl3K6lDygIDyJse
74IyBh1yI9KPbT/4jGMugX8EuUdQnQZ9NqgRxirdFfY0g8BU2tpolelA6vJx32D3
BeKhywrjUn1eeX8m9lOVm1xmitksaDUZP8pjNStZHZSKo9DI4g1WVdjgNVPY6FDp
3NFMTTAvqRhpgFG6Tt92GlUzTu59aS0y0UppGv6kPJEWGdS2lTSfgfad+lnVRkPs
xGJ5Wnz2Y9mSyW5gSrNuNo9QIOh2A1Tg5hSdqs5T9+MI3DSg4xZYKzo8uqB8yGfV
05nKRgHvd9zz14R8Wk/qQ+gju5+j4L+eMEm/14FUMqUMEa/e1wPAuCWhCC/FL7oG
ppawo2igz3ArtgiUqgJXvAaWoORBJAlqBiLYvHWQm40rUhgbXqKWFfNIUPMV8DQB
EpO33S5qd4LY6OmbLSDijmZg2sWeKcg5jO8N0SHhWX+6j/7Z0SD9gXEPwxeEg08Q
DPaDWxkT6H5Yw+LIvyaxsVll9nMd+M6VALaeSucbjrnnn0oorE67Z1XpdLoA/goh
eFxGZ9EQweMDevsbnSurSUx/zNvs7qBxE9r3HOEQa5IzsG2t388CsZ4v+FPeckxJ
fXno2LG0uz4peoJwPz45SS1b5swGFngYj+TDz16Z9hd73RtjXPbmS+YxWWDI6jI/
nLRUA4nTZukiKxvB50psu6IzaqB1+cttv7XXNNQnySHRlli5LVPdu6ObKqbuWb3r
IFsV2ArvVT0lT/as72GhL1A6mP8EwI/8mA/qbjdjwgEJseOOVP2I2CIJib1m3RHU
HchgY9hfYmsdYltcUI1Dp8hbrUUSgN3ieOCofFXwEQ2AmYnY5ftM5o/vn6EG5nJF
EGojqY2p/ZYv73sSrO1JYcRQkMdN2IjYDptWbK8vufzlkgvN/yNXTnhDrzuygiLJ
qTSeZ2jCktlX2AmvgmO3KMRnlp0mSFzdYqb2vKDdiiKP5SUu9WAvxRK1Den91Jch
0qDHSVEsCRgKDcpPtiHUavLIad7hNeE3JTAirNCtgR5gFCxMcqJCeGJ6ikcP+ktl
G4SnUJKMVPktUybZSDMpnke2h80Y7G+PTKXMfyX+55pBNtiQ61KoaCLTQqnwSuRf
S8cQsk/hEMttIC/HDicJW7qoaOM5HbPgy9P7wGuXs+zohYD87SMzSJMFo7gkQnCY
JPMXPtNq/+jez3Utsb2ddQJZmLIB+hKetyKJ572kVPiyLbfx7LKxCBejGw4iM7JR
Fw2Ct7+ZDMZtPPKxConL6olaJfBAv5bA6l2a7jP97TaY772H2fxklemvpAtmjMcN
vI7oGCbraujwjg2XK1JDfvnKi9P5IC6F3fjKhqcFwKzCc0kE5F5dXcl6D18eMEOn
AmpvUO23FqNhgq7UMP38gSGGTBIBSVKE8qK6l8WPQLEmpMgGIL1joaXbc0sHLtzT
biAAwX4rT+Ty7xs3VXcs3IaSaJLhmveS84RhmzHC7Ju7qcWYOOinzmZ6A5g75CZw
xbRDoHgrxJ6jeEh+okWVb08se7k0bV9CSk8Bv7coSRt91DKXR/mattxtH2evdNXJ
lOdFQOF4KW+JbPxMxZezzh4t23yOpFvINhsjG5FmRpw8pB4Vo8iDAl7tZzZUPVqI
NZsbN1NodTzadt3XitfX8uK6qQ4gHoPnoOW/GgZBD9yef49eHIWe/ZZCIlk3/U8r
888oen8QYAV2M4gnE+Y/E7+bvEM3MmWV2tUgEJ/G9l/IhHZchpvwVHYALpjCwMZ1
vczwSRo895acGXqmRfxk1DaXWXO6q2BK1tK+IK3Gcz4PAhxUudrZtRJ7EJmdcoUb
5Tf+MCadk5kABUeQ4RWHAFAFlO4Mzt+I7mkOsbnLnx+CC4nwDU/Rdez3vOQQO7Kc
PEdY4lHU+09lLPPIYtTsDMBkUUD94uIre3A4hIL19y74h7Kv7PpZF50w4Lun0yS5
IsMeeyijeBFY2bcaiw1i9VS0Dk1S4Cpi+FXtZSII+O0CcVv5TXXe70hFZNGS23hp
OsuFECmoTNRwr6yNrYIc1wraHJ9uKxh/3/ByaU1oeDyihREtM0G3rviPomnHhMtb
6IAHcbYoENpprl5l7rs9DYHSq2+rJj/1uVPsBHrygVMSzsHSh49yP5wgyD7suQux
ABJN2Dtdfpuget+fp2rm2dk6DmHc4GQ9DXSrg4g5o242zNhJmAcMLTI1XnZVy1B1
u6UBEQX5uWcgqi0n5xPudGhQRpd7nWFdhhoUVqa69QoTMn3JMmWSr1CDvggcRqWW
3Hzyr2y5vdsui0vSzdeROSNavbUNL5yr5zvplRhsmXDOaUW6sbhNdsDkksYD2AMY
sxh43SbWAOMEOmr66gbFvF72SiSt5wlGYSMDF+Tqsib2ZZ0cmnqXGE2mqiZ35ZW6
9aA6l9wzRYEUmSGLKH+oF+FT07/mjrvIBAky2taEbi/l4kIIAEfLS3gVjSJyxk8U
I8eED231gJ5EMs3Of7R0XOqWuUebA2V6XE5/W4R+2enKu62/413eG9uT7y3pguat
5kXwsvxPFgk7D1WT6/M5pdzBWpFRqiY6Rn1COBV9/46ftMcNssecrC566R9T/bKa
ToPacOrk76imJLcnAVkARFCt2R/QpB4zlAU3CGfnwGaDg9CWDRgo10uJkt1mIbpx
Hf1owDnelBkx76fEaqZuLA2C9vji2eWP/D0YYvmWUFhjH4v+Dxv48SVQzkUZhxK2
t/bodOhLMnKuS6qNPDUXBuE9gsdzBVjjVc3/NZsZFdM6rLPNhEcdAAEBXZYTcWDz
4AyPA/vRLlzNHmDMa+J7F6p1Kwz9Zh4xSZCuXNrT4Kxj+guxvxWbpxZobZSsFY4b
salunUbOuSUV/zCB2p6hqUkX6ivApWjaWVFNJzvH12IwXkuvJYRDigthVm+BJetX
qhieLmMB9Nljp2PWp/P3Mt4MXWSGSdwIYNl+cjirNCZZWvTqts+cGUBML8UQf+/Z
17+ebpt8hFFKhB7kkHnVn2TZWHrl0a0kow8oFQRSlnUa3m77H9aikc/FL7ck1PUi
kClsIw0EjlvAN6MNTDSUZINRCE6bc1rTtMYLTSQosl7zIR2Bg5RuuSNkJjuPuGsi
ke5G2pIp8KLHPsylw6SwueJwRjGf14g8VZqTdPEbcR3KNQKkQetlc7bSDJZ/49sJ
eKRFpv8aiLoPNLAKeFnu8m7UXei9ZopGni7oLqs/1CAVwznviOfIQS61ZT7SK+Nr
zc/TV2x6JAkuI6D6CUmVvrVUTDCNHiSsyG2nNqnXwt1L7nv/21sX4KZN3BAnxDJM
D4WAfJq9RgvUpwX+9NGLJJNpNZXFl6LWVsFL3qCpZXTDijJLg7sh7jZZjFI73a6C
jmi6/Z0sfH09za8vByiIfAmnxJSylhH7GAhBTcPgK50upx3Yq1ZH/pr0pFEvMFuC
rE29Hc3EeHwvzG+P/emk1JPLdccYqO+/WCgFFC0/PV1jyXzuJ2/ijddKJwXCmUPR
W7E30DN0ajeWubStRA40ZwwktuK/krLeNhJZnEW2g2qegUVUepjDEUyDro+eqOPQ
u/AVrhCDWG6NsqT1gEZ1OEmN+zgtnpLPkhnULl9hgn8Pgfp21OtoHbRTg6yJOPUA
E1Kb6gY3Pi8tUe9w+L9GOAwRFgcr5LNp7CYMNqCV1KTT5b8LjNE6eu+UDvQGeGxF
e1MzcUjakdziJD5YWZ5T51OfyRLO9rzDIw9m4rJVHlDsCAUMniev/G6LM02Ge2PA
PJ4zdS4w/Dir/HSLj34+Ye1YfMOfaRC8rjTPdlurTy44dkXq/hhgsH3U0gvmg8wY
1gTBW+M8j25V+mT29pVV+v5SUobHJh5qNyg1FudZWzQvnQn31v8DHUpFAXcSixPP
JmN7/7+5FcRBVtdxnFF8cFk0lbZM5TiKRgJ4PnRmCdtOjSGPVMvaH/d8U4PPwG3j
dSlLX+TVq+TwuhxI5X8Es71FezkDqwnj12EkeHoLBLWiMGhS+tTSUbQyumXEWU+n
szlcaNX3Uu0GlLwc+MN25tHFQ5ypthqkXv8u9q+cZVlAvaz2EPQ5pvog/klZbHla
elxih8H0sy8T4C5zw0lW3uBbIp89HkH1Wmcz83EL9ar6xiKE05wT5K28cAdrBMe0
HiTI7SC51gWanyubzy4rWEYorrdgjsuWpkJ24CrDV1j49mkiNx1KY2O8KK/EaBZj
zrcaXFktDJVXW4nOG3ieL5M5Jbc0dOaSM5M8fhlWFfnQJ6VHWfH++O7rHYpx2ua0
3YpKszUadjHn1reQQjFZtnhKD5x5PG5qBphoAJ5Q/f9jaDENtnbhT/fOIlsT04g5
ucvrLmo+WCVWvz85PlE+N9bMeUy4G3uxH4KD5zO0RG2xopoWjORaqnBVco9w6Oz8
DzDRyFKLCNzHiIFt1rmKbthFhGe9JvOIN3jhuRbEgRia2SWpuTJ+fYyqsVTAwIIX
tWJHGn2dRwMQPBBfqFZ/lVOoaar68ZfJjtdaFpl1RbgYu359TP4paIxhbmoHHUMP
TakYxLpqoeSfqrZznqQB+5+Q+34OxusTmzZpHWYWAi7r7CHA3QP2TnHHhyDoPD3s
xCLl8Qcdi5zVc6EXQlePh1byxRCDtJiL0Y70IZ0nhZi5fdLjJ1KlfQ+lMbG4S03w
ZpQdD//aD68fjIc42AgnC5gnjrZp0BLfOPe3NulThEJ2sVjof/7OsrLw6ga7gz6P
dgWWqqWEiJ8Mq0nXpF7zruxC1kydAu+v2CnAjaLYORsGQt1JvzuL6kpS/PUlYhqc
uFWy3qwnDNFaOgmzVwan16kuST+K6kYeX1X/fCtc5O4pypGn3C15qkDzn02DU5od
WCpG99el1HxShKp5MWxhrbIC2jkdIM7Ek50YlnMdg0b+WZgox0M1Ma4l76WgqGaQ
DgSJibqfUEdhHMFrb+7N9mLD9tBYE1nOT6fKRfevaJEFq4+IFEKBTE60E/24r+EC
GYKK/PIjRL6VCTGar+Zt1zJsyyMvCMvhunEXlK5mMcmoOXd5B5eGOqMy7Krl3PQn
NQV5HC+m/tLXjbNbkIQUe2bUTmm4k5mVF3UH8H0+CZg7YORhci9owfHzWTt+plbQ
tFW/8FRuvSsgyftdhMFlesXQoy9C3xxPiF149abpt6kvpJzUW8tLLc443U82/Za/
rg/LPK5JeKqiVEx8ZPjR26dAY6ia/VHgG7aL8EnMiSgQdcpwL2LzYY175SEP7N+Z
Dgb2Xm4QXkCn/IwMuVwHEhFbc0MivKihgXyb2MdceyQovCB2kLP+uuRaf5RIj6oF
bFYlxQWRW/BCYFxN9E2IqeXbnIyfM0c1I+t46/vGhm9UDH7OVNh1q3/a66PyujF6
AF/sa3c/chPa3Xgz8JdhCSnbUEzPO2zgZMD8GEST12OkND9SV6jfOtqHix/qYbzQ
Z6wigroVp73oZq0JAPPaO2KO1z7ysnAEgswaFs76ulclSZGtvhnQZgknzMPtXjYv
ZsSK7rTDz8w7kTpo0flzKJzY+q4WXzEPZXZqG1KtfbODDZ2IjsMT4eHrm+3ZFpZ+
5mdKFw6r277AGMiHd0N7HKDWFL7X4evq11xlmBwSkRX67Uv8CznedBpxK1sApyoD
9o02sF8VoMq7uSBCcMNUdj8sOvqvONVvlarfdbP4cLNc7Rj2AbWQcMLsONcb69ok
f0DV5okf4yvzFThrWKJq2j60escI8+FPp7KZ6+jwnqTNd5RsPDB3i283tIF9eYVA
IwjvPZBuf+dEi35bh38Am+fL06hkTrIqVttujZEDpa6QsuERbHN+a4YZwMCAbcOK
fi6cEbH2M7D93uqTUiEWwyMWpvpNwhpllIXBcevEAzwL15a33rTuLuKNRtjn3+TQ
rrHxOH+OX+buOypIuHtGDDnCq7QpAGHigIE76XeKybinq1zPmQUhLt1IqToHvgLv
n4AJaBwErtFKUkRwPhfJganVRJ99gUQ1/Eb3YQJ14dW/G4aEweoYKd89bYLJiGQY
1HX42IEdxJdvQiocGqLw1u+M+Jz+pAQbL/4T/l6UsZLmteB8GjchfOZ2a+RE7pvz
DE3KwUcBy/mmBtea6zZHNICXvmOXWRiDKQYCUOoMHlmQLKBDaPcm/J6Ah4eyyFH+
APqs7EmGUzO2M1P8E1nnIv3re8z7ec5SMoIXE5r4sBpA6y9ef9DlUGc7rAMWbb/7
YjvYI6yL6W7iExd4cb5nDS6S2XDbV291eSLPQgMQEeU+sUBD4olRMFynDvnanrrc
5QB88o94lvviN7YdqiOokNyX/VWAwYnGHMP47dQ0a/j5TXdOIGWlcySWx+OUkRu8
rRbtfQxII5pp1njxcLzReV5a7LAaqDUPqZZG2cEeMG4muZZCnPfDdDYqxMMB08pO
bqgf3VjzqTYt7Zr6P38D2VaiWQKkc/XvMJhecPk9Ia2JU0of6U9ErA63xtbxbMnV
Swr/w+tFIeDiWKb5Dwzla3kyOFvUvpG0oT+vXI1RwWJli4lYmO0pqn4W+H3C3AKd
FA+NopWDgbBzv3YDavFG7PX/5LifOB+H5sT4PwL2ysRP3q/q3sTX5JfGkzzagOmB
PJfqAmCGWcM0pEhGQFnwNiKw+/Kf1Tyu0NIwODXn0vt1pIUhkuin5ZAvKQKPiIJ7
/3RyUmvprLamX0cJiC63DaAJOCt3VCuLeyi/5j3AgExOgqmPXMfJXcWNlBWDn9cT
+GU44t0ABlLrwiG2Vf8ThnN7jOALjUMpz9yzBa/lrmqdSoC096mMCc3uER8cuHHF
Nj7YKGPfqMGUzS7oUr8vJiQPJk8BexOSIML4V/kluvTWLiGRBV3mGfhLM0OH/wt6
0t1BoLEkKLtKlyZqee4clrz+iWFjjwOZcqzJ/9TUS3SEUK4dNGel2iC6Jfaco5kH
Fu6JKpjvOpZlXW8z7e3x5PW0tfA1L4o2K9B7ffPY1MoqJTRJxYYNoYTjurEftDAR
39f6ppBYTAKnElsfac/A0+HpNQqxjXAFokhydsr8q0u+9SdlZPIVtybWF7ekcskF
4cAkercxuZ3UgnS38/wspPJ+BfjpzeXBGArPuUu8FFz0Er6cBUnqKzUvvBhrDJY+
fpUBKQeDcrliV7QALCLDeope6O5OFhu0LIaPSNeTj6t+9ezwHImudUhp7uM4qN3W
hKkcpx2aYnYTzyouQG1naTdq9P1IIcYRmzQNX/+amrrCbmkkpXluywWm6kgFTpIt
BpS8tXr+gM2Dghc52Vr+1Qi2jk6FU0v0tn0c+Smnv+FtQRYSVZiZ3BGahFFxlBtS
74o8SI8vwXh+X6DeNYSiH9y6HHMdfaMsdVRSgfxP/fobSEvLOFhC+Tm5ztZbYmsV
BLi1fYF5jnrtx6eR/WdY3RIjgWHTMs+oT4ZjKgMwX31eGnGjpXTn3vCKzTwshL2Y
FKzM836na332gP2ciWWieRpzf4fOvSCAR0E3r5fKqvzdh4XzQaS2Yl5EOQotFTSO
LRaNhq1Z9edevRxzmArmMAQnOe8k88wb40c7kZ5ABCyP1ImHf8FuEHsrZIzPtrDR
qFnVXx2PGTQ1OyZxjGvJY1flqr1Jn2cXJkumfhmVqQ4MocF3Zc3r6dwz8Ha29wqH
XyZrctgJ3dDp9yEsgkQX7IuRAWmBl5/0ZLemALcMkYie6n30ay3Zku08IjejTpvx
+2Dh0h5tItkRCa0PCoaxOBXxu0vOvCerzhevR0QqJ6C1w5Ig60p3VIt9FHwC6i0p
IoDjVGHufycDp5TSbdyByLewdyuF4E8EV/vK4xVNONu2r6Pspiitl+CPdwYiG/J1
rr5GJgXSRUzocA8JSiiObd3OI4U84Pcp1vdaOlrQrxQXPyoWqwOg1YYV9rBriOs8
jjcBe7dtm4VSff79naApl+QWqrwg4sdiS1uStPzlT6eky5W490F4wYWtTRRWteWw
p2ZnxlsXE4uSGCTEMQnO5I96LbY1Tjqvty3a8CqwM4TSiCDncD9b7JhDED3RAuv2
/ngTJVaNlMsUxaF4fMkUPwQaiHQ8oC2G92blwmOmfC82kPCEvRHN2bernjSS3o7E
Kh8Q3FGWmMVNst7Fl6x9uXn8cJ5wdekY0JkX+rzIPvamoDJeZe0EI9+azeL5NcEE
ZjaUzCD2HsAIVxARTEHHpbKTCQH7qYa9kSzYoQsVXAv7N+4R0PiGDj3/ZtRAWT6L
JborskZ156sZt4JB+448VYtG+fCEBF89355PpGDUj5F9rdNWnPu1GnButE2DFPux
pbDOwHM4+hJbe4Ep0U9D4neYaFmSvJXEg1UO7uMwxbGJApV8ALyzB/A1NKO9bhfi
YP1x9bb4m+FJ4f4sBu7MNB2j2YMvgo3qF6qrnblHUowf32yU3YkreCJ3AeHOftVA
ERSdfFxEEIn2EulqvAYYiKzXNbQ72XEHIU5oQXSa6IpKstaV1q33CBdbQjw2cjuS
Be4O4Nw2MjH3NrtBRrlUCcbJMIR24Mg2uy5EXTruYAB0Q4wlhXijZkoVeM/zFE70
LrgXyIImVONJ9sFa+Whq/qrM1dZxyscBH5VfQPBcJibXzULRFUYG8/52KTVquuzh
hcnWMj51+z5C5uZOrQzB4yk7BYgzLKZTXhyxCtCY3fQDc245GcSwGzR7f7ooWM7O
4oYQEDZsCiEMi6ShwKopqVBIpJEIjpgB2QfQZGoj2oN5LXrdUAr0UxGkJb7sVVsy
wT4REx3P1VGBaL/lpYZdDiZYjQkKDy5szQgDM0qdB/s95KqbeqpXad7Qb4BCeL3x
9sBI2/SFxS3to9fxiteJOaDLsv18ggeGgTTgxZH4K1b840BCy4KQBmf/97CNwNBa
7PzWYHH688vg1l/E5iJXDDNFUUEky21p5o/PMdXkrvPLNQIXmYdo4AnFlqiFX2vU
Org7GS1X2ghqZrhVOXFu8P7PnHvNeHtjfkjUO6NmDYvbzgnP1rR7JbMlHQHg0iE0
AtYtQ4KXF7YayzF1u440niMR2XEVrMv5IpOaodLRJmz1T34kcTYNW7mBKgcZblbg
i9TCj+3CMGqpHcy1cqBMzHfJ17VVq0L18S3Yv7xOJSuN3dGfO/b6Df+8MORmdND4
QO2PMPCAaYKrws+Hih3Mr7Jk2QWQFqOrXHugHgHQ8eQXpPQuGfeDqqubZEsp/LjU
nBAAqvk3RZwrZvr/wnXyB6xYChZC9+SYBnVe2rYoCM0bvj+VxfCihsHBWqI3Q945
gHZKReUpCMKMWUJu+xI0vS/duBbGJuLz+MBFQ77f7XOX25qvZ4Wiu5Ss8lY8UtuU
CR0L3/hOXz9XJnt0ADp6SjCaRx8TFtpxCLHTpCtrNUuxf1y6TRszfG34Jlfe+rJ8
AdV6ewCyRLCB/0T9MXm/tEeBmmcX20aErmGi2hXz75DJ9hRScI285LP3BfUH/sXp
glKo3c3iNYAm/Qdw0+0+Gh///o9Ba4eFxuY/UZVs8KbFVKqLup8dG6MPoNTlUFGa
FkoidxAfzm0KN2us+2bDmm8IhatvjYmnu3q5dyoIvrEO3bv9gjav94qA8/frjY7n
vI1SxLPsQU0wQYUYD7t7lAn807BGMQfNOmzeW36pzf79Fzui5fvtH7Wsw+wIFXMQ
BMx0+TwQPw/WtkpJVFQhmRSuKZmr/22tCIEFSOdaWdaEvxzwSxvGd79ADutSiJHb
2DJ8C2SlCdVUJCZDXU6ajjaurEMV6CBPZIfYYuZ33eXjyviq8KC8IEQ8nVs4Ecvc
ayRz0mEu0gf3vwWasKMtR8uLTmL8nYlSfaGwl561eT+CCaK28p1J9zWqvPPldzSE
O9CwrkxI/Lw/fBO1tQKWC7GGXZIM8wJMu+5O96dnX8UxaQCO2+64Htz9YkqOX2KY
BCTcXFv/Ol3dILOLn7B4pv/FXGBiARm5Y2MW/H49sN5po79fJMXcolQSnvUClIvV
oJJrSEqvueaxpf3DDU7hQI+zvIq+2Klud1+3YVHMCel/GVjh966Ccx8LBPlIRe1a
jNuYhIiDjM5TvOpNTZKRw/GCfDfQPS4n/oxu1DLKsY77mXoTguEtuA5ANOCloz4h
HXMJ7xV4wWwNvsITDRptb+0bkofgydVOnQhYSffgmjPKlDFFK+WRrSTfhl/tDzI8
fzj1K972I/t/t0v9JUDaZgPWy++xR6nRsQHzGXtuEBwh0LLZ8muvGU8rxxHCRxHH
U3koentmYRnoohhF3/H5fx4bBvnda4ZTN2ZbGFLAY4BpWnZhocGwykvxy3eDLn7r
clxEHIWo227dRp958+reZXn6+yrHNjoNWoozaF9uuxEUFzMFvV+k+R9q+OQDUHQW
3WR9gpQxN2cQNXMv8+WWju6ZaL1HJVIIcwpAAXQT2E2LiKBB82CAgW6ekYIdFZJi
Ws1hzIq9UumHLhC/XsG8ox+kzJcq4cytwHScqukh5ru51AIQI1TGIvuJk5+I7hoA
ZmM+xT8sDXPW5NNpvIf+Tu6CXikuBod9iboLo/XCHxESbQeqm2q6U3TShkZIcNa9
6mYrq7dyzijBDSX6R8OwfpNQf4c15CgKd/YYEq0NcODNQIbKHETHVygRjlEzsgZS
YaA//v4qwH85kYMLIqIkZNWpp6yEaecy2thVFP7Tzc1ciZt8axd7dO0V1OGpllA9
AJ5p8dES5nlirigXPrnrWXqj+p3K/E4hCEEX3+wnRN9F11Cwein02ExE2pAJJrOx
t7/T18wLRf2kNyE6e2tD3YddmLzy30Daxki9hBySQRHZsr/eY8uJEEM3SRUXkvx1
87hrwlcKyyw9827fwnvlwNyxDkKx2g8U8uqtO+abcC7tqNUn2JdMj+CWJHjzzUFN
LKaIP+mh4jgk5JRdbyLQbzJacCv+SPAZu7anYaKnAGd4ysfAIVD+Rng39EYdnWRW
dHNYYiaEPRZnJjjPgTbZFlUA59rFQbpDbnaPp481UPshdVpvKlPSg87oYmRuUEuK
1vwJ8N2AwRiuEjesvb3GXWpAbpV5lCjgCMizptqR2xuV8aNaBGWmWvJRYFTU1NJd
F9vqehrxe0H5Tx4CKwc7JmlGrV/f674Rc8+llSrWJfe/T4uohTtwiggzLPplqX/U
yTJgs/i6jNlRxUZy/3cqhnIS83ZOMxQgMS9gm/pibKtdMpo/EsnsMOZUBhbcZzgN
nG3iceSPdC4zl9dZiV4SFhIDNjumuAGczFo09E1AM0Ne0VgVLrmzpX+P7fX4DnIJ
CkPc25dtPvMhE9mOIRfKWjCxGbdSf8HW/xhwoodPvPyEleOe5H2rtVHiyf/rwvNs
xeoeTO11LSl/mPZblGXOOJZUc7b3mduqikWPIpDxGQkv8XUA+MiGd2EimxRmqBzW
j3Hdp45BvJ9lP7zzL/C3VEq8OumP+EMY9ATMS8NicifgnJOEtLt2uDsofjlmJpEh
/zTiq8xcxYWEmynZk9Zot5wIrWNrN8J3NC/YVhbo5xIVcgZXSr6kIbX4UI236vTo
vyf7DLaa5yRRQvIdTClnc5iAX2m0s3ld6FXa/Ct8scHARkt7oYBS9UPhcCsk5AbK
V/Ekr0gHbyXf3MopqH4diA3FoO4/1TvdATP8IbgKHvXPpc/yYN/WGuaqFIqyFn1+
VQ3abotVVaglr1w4c+Tz8oa7KDJ4WXhCXey+bo15S6r6/QKPHMlBZrYdfUlG6jog
UM5dNEwMUAAfvprkqLWhUM2XT3pZWlLd4d+VVDC+myeVANmRKkN04n+05dun+SZN
oCsOZoI52reVoIzTYpiwxS+KTp7tkFG+i7AZwgnZgf2WgQb6OXWwfdtXl8jJwEKy
zwN12ppA5dLJ2yOAP3MfgnBg+yAq4+bCRB9BkaQPZA5AmHPvi3xuWbBu9QyAfqaN
3a5Pa2grQXU61MMytVur7ai3UpqzFC4qBdnCtm27pInhs1Q6hawJLC88teTmjlYt
JVLaQND2ulsExZjQih1XWNFbOyhNmWwD9bRPfYnPJZIamrMR2m4p6oeY5700c5lF
1p5Jcu2be3zqIpb4D7V3iXWGGJoudbfwv7k9toC2lGKwPeHXwOOYC6oTb6nXnmaO
3RVRvS1FLppDyVDXUA9xDnK5k11FcYWi7MKH1b0ASmxLhn4I43Qd+Y6XkFxQa+dT
HPETX27jVhiOlUvCJtK5Iqppt1MRTkPIqtfkQ8c71CfnledPzALVhFTNIt2IEstH
D9gyKrAqIJO3GUGiMGZDstKRJkfGp2nktL75UIJMVlbyt+UZFejKYfQKokfiX6b7
twhR2/PvRYurxiscJEGRMWEF/rcf15abs26OotfTijfBjfH9hsWAvaROcYQupMXU
fjmhWHZsPsQLwLss7zK0UBORDrupQ4GVcHal3cHXaAgZkiyugXuHyzDfafA5OslN
MCG8AOB7ZpcEp6YYMCIAAj7f+fwcmwnfRSUzORjgWK+DDBI/Ny+zwoE96Tx6ccBW
vUmqMMrx1Olzj+8pkoHlJDaJrr/h6mBxt2y8B4Go6C37Gdwb1R/xA/FobkUePUS2
DOBzXtR5s213yfINLupMPChfLt4PNPsqoAWbd2SAcTw3SlZYX4itStFtEFKz3roA
tHr6ijm8H0+ontUuFYEn/2aiv3yXMcBVyP44gGXaAgLeSllYaqVAsQ2yjV5rS/Mr
5NHn5BbnmRqG6CNdeQ0bjhHPFaIlhw9wf70OSLZCAY+8uMZhDOoogz2l3/NRN/N6
91RFVtfkgMmUZI9ZSGlFBqynxJ+/rUCpiH2Y/kGJEtKHroXFvHK3M2nqxaKa0VKg
3q7SMZlOJYcn63i4N3P2BTbeM+nzgIDmLdlZ/u5X+r6hWv2xuM7MxIrFOoOy8tqz
4TCKsh7lC4JnJlo1bvl4uFlkMDrtjHZfTPcPlhbol+ZL+34LRzPLd7IUsgIdPcyG
h3CrRgvO9djT30TGG4Dl26gbxhaVOdHnUbXtsU0lfw6KgciqoCsDPgwbuClvjPvB
3gGdv3GpC2JnbxZwrVJ7RCB2ZRapCMeenkQruLJBkZv529va7EQJPH/ruN5YQHJP
82U8Ur49NQeAyA9jRynpatwXgjX2OOGiD9uPYVh+8T/6zlcRsS+JvUlpbSgQibua
EAWcqSEnbwoHwOkDwww0hYJxNUEVYc3ztZ1cE7Q03hEs2a9WwOQBZXag8fA335E5
3/FRN/05xsGUiiXklN07gPGfFzhmQfpqsviZPbqAXWZs+w/K2MzJkV4D3b3ZlqUR
3ma0sgULM4cuuf9PWy1urv/Iec+L2nl/TrTiPtWxFu20FsGA8cSVmG2MEAiX0J+K
buOQrntK15rZtKARncWG4lTbFyrqS8bhNrmiNfWPWmJfTewtWBUkqr87URcc8mXi
dDRyVOZOv7KCZ/DWxt/xskNZaa3yeXCLv2ramy1IiP+hBuCxOLz4u2kGSMtQ9NXD
m0cxlngxWAJ/+GpIziGlJ+ljjtYo+6vqQleKfARSgAIM4ZgL0TMTPrKOhH4Gu8O3
9GjY/beaxABkfGxS07oBRdQm/fI1Y+t1zB5LGIv4W3At07tOZuJGsYSd/xKuuZYr
U+tXv2/vfFM82m9Wqt4oMWKu+BmffuGSPOrSfOltHly/wuR+jO0alyBZbpiRE+hu
T2EBNBnSlVvHKEW8wieHL3Ls8xMuyjsCT5+JvGLZNsUebO7jNJ48vDhNJJcM9Oex
nkYHK15M4WOj7rXVFFqV+ogH/6uVrGIPMTTtVQgbL4QiiLoQjv2vLjUFelBM+EaT
/mLGEMeolQorZx7c/Tf6itzfCFcs7sRKsusZHI9uIVLpINnfkmi1ozv2FmdxmQn3
OVunkGdkaPuoXk0eBmNiJtNMPiegEWErpkSlINx0WuqGlj2TJc2YoEYkpYdbfTsJ
6qWd6PztiVS1AfTPUuFmCVUsRM8knyLvsLweulqM2cie2Ovm/dWsEyFXTtDEqvwx
qgmU0V5EA4eW8w/zldbKabzmuYYo+pVPhdrxCsL6tmthNl3U9hDOPrfzezm6aqmt
Zd+uBJQhuQDwdses6W5NVV2Ze7hsMBgGxwwvPSLdv3Iakm1K6GCkCcaInAMP7Brq
CrSMBTmdayFTvThS1HFPxg23IotHeV1/WHk1wnUoHqHH32IPaWGeuO+Tx3PUkagz
vFPvee4JnTs5P8MzUkCp43WkKbnhtv4ud1w2+smoJiSV8LLmUYm9kSAVtMsGTSV/
bFezq2UyfjlmSHVu7CSu+6YcfkqPuoX8o0s5AZhPXQ9Ge3OVo/FGenXl/tOQ8zK8
ancFEshQhnsTGnte/Q0caTbDrhk1Mxyl14EvNjaAawxUACymmEc37zC/BDA53a9U
XKdtMvxdYzBibhqrh3vxDGm4R3BmDF5CIQgrT1nSHiGSHN4SXR3lmMhtDIWgG4nc
Ywu6s2zmzo0mvzT68VjFX6UTJUGsgJuH2DNVDN4HYkk8XX0wgIl7S2ALC6h7lFzc
pkVq9QkJIg5T+L9h/ETl7U5V/JPcJonDljSqj+ualnAO5YBew46YJ2s0Ym5Kv9lN
yHuDtOHdNBfDWsiFyws62htI3C93MQc+0BLulpYJud5tJ4QuphdOoKV8ATPsXYUg
Mr6mw7NLbr+eQD4PM1LkZoitEm3pv/SeVSBUHax6iKhB+3sAtfzMSxQyInByauTX
YL7iyCUlf+GFM8B8Vu0UleUgUT2Rdf0eY6ITeUiMXSI6TytoiQzksx6vvTVMg34t
kIheCwhjwh0ie0OfetguRxcGHCTMXJo6M0myxwK7e9MZoIQrCygdGsiXW6oFmd6h
U1plqW1LBmC/qnQ0Ky2i63n9kuta+WP4oG2sFQAxE8U9CJBrBNv+o5v5geEMje9y
1GHiSqiiZ1nB09gkKI81OzMzUFyytqbyytE6MFBnSxY6dCojUiz2+5eBgQ7tPrwf
kuTxwP4Uy3lsXO+b432unxtK5YwWbKwRPgtw7Fq8miqU/euXBgsmd4qgfmSmxP1V
I9qAJkZzuY+S+ZxEMK/BRbdVMmMpOWr8/a5BFRP3Ve5ssceKMVpF4WSL85pvQsCq
gGan4qQVM9zycOTJ4oXMwIc5hC150lm+PpKTwd1EjmtOwbKn3xgh9eVLpfhql+bs
/MzB85igzeOlr3anLUAcu4UUPKVcH7PLtwEriK7gq2RY9X50M8Jw/1hVEO5Drz4G
Ty3/Y2RXADoz7K5r7rcu1iO7tBFEqEjgGxc9YUIKob/1i9H3jQnqx7tkO7EwDCw9
da5u12NlsDIs73mudQBcWwqLGHJk5OlyDhyEpHJtzk3mt4m8dy81zt0dVTfAnLlb
tN/UYxX4NMzXH6aHZVFpiOCsyAIdQub5A4NmhREARH7PnFM4z1WQQ9Uup0NTdJqY
K95JNXkO5KvuC6ZlYMfSiaKGi+a6ro05yDCvpIxn7cmnoCe7on/a5SkfFsUrmyZK
APg9N8mEX3Ak+GK3eVU3zJrbJhsJhUnXmrtUiCLgzDaaKlcIU8uFNuVvSo1EdcoU
axcFx4uNh8XSGQVIs6hZ7TX3aGkZ3XVoz+xfuZhKzXE0Z27IyAXbvRo5uoM8GOA0
jplCMrKN4rT9nhJGFrYPsyzWN28C14pogiPo6qvZQcViz08uzewoUX1HyfQMtHir
V9qn5yr3ih2cIEwLxnzSZZBnYbizn+TSg2+ibVldv4Emi5Hgd2EluwDOhb/Io1XD
/4wQ//xHgpV5AgA2v2etr7W8KAwkSzX5/yHRZN28jXmWHxDPoPn7CiZ0lMeWw61c
1KrEY+rS4JfspVIQy/BHrV+vvpLns7ZB8UGmmPxTNqf6D+g3MOKzQIhZD/z0xMKv
ToOOIEGPZCGersoS3YiwbCfUS6OhpC6v0ZDM9OmLRur2hR9LbtTQVqG6nLZ+Opg6
7JKjefx2mztMxsL1/RSS1OrimxWBHy8GbISgHP9Q1qYfw5co4HjXZbvH0nqk6E8X
MCesbMX5qa1pxMuaUoH3NAGfvribe8ebWE0QFJKq4UlzMbjySo5LvO7zzir1sJpq
9hdHp61UBX0/5/TY+dqPbvKL6XtKyX91a9cpuVP5qNYO4/7yUKyE164ywfNeHOd4
a5ZxT6cih+O7XXnAP0ZnISIMX5UKCCnEBlGVjDBcD3HyjdG/YnBozt92MyptgUG2
Mmpmd8Mc8unRxSzfnHzUUh8bOY0nzt2R/WdJb8Z/yTdi9201q+DG/7s8B7hlK/bn
5KvYEuha7L24XVwiAP/SuRtBi2GBYwfCu9oIb54YOW1ABWyq6aXKnOQYUbREjs/D
7aOxVF8o9Hyn5XiQmvPRqXcHB3GFBBXOxR1DsbtlnPXlAHG/UxthLjS41YV9ChDr
tl7kwp4vytpqb757hzwJ0mNEU3YxXWG2xJbtGwLRmoatLjSaSftrLQSq2ql7o0eq
NOeHiKPM7HVzV9BNZE/jkU4eSzE2H7jYvBJ48F4WkZwmhrYyY0mYD4coxND1z6u7
jGMZxsO63j2Ea401315bOWCH/qWZ//Ee5e9UHaw8kjPvMcS9apTP7O4Ju9zTA8JB
M/p6+9Q7scsK9KZBnbaDrCGNBu/3dDgYrAzlyT08QX5Gov5mqb/pwyjC4ZgKj09r
f5zQnROTMI1NnCssAFmvdzDtn33vZgvsWqbr7YJjyQVDYEQXwYPXwWu++tUnZ1/Z
cRgPXtoSv7V2zi6NxHOfy6/8mY9mIxlyDtxUKqUMLEA9Ceh3MJoznmn4ATQuY0ah
m9Ps57nX8celft2X4SfVL4bYz18yjVEqEUNrBO4DKeWB6emlfUbq5/Gjq9wlrdwp
j1k8HzYzan/E0D9R/XQqgoNiMEgLPi8IM3MQC5iMqUBQxy8CsawnJ1RceXK3eeJj
ZfJUxShb62rScNtGvCtOz3JJK0EkRPQp/IRqLLR50vLPrjj6H3pg5LKBOEPdmPn2
KTpfWd8z/StwvlzMHOHKdOxaZlS6X+WtfoaoS7cL6QJtY6vfX/JDqKCG27ssyaSE
8Q3o8/gNQlWEjV7h1U9lp3AuGd91I0KvVl5BbBK6HwAHkAOX8qi9POvCqolCD8vm
MRvsF1OJkFsQZQkclRC7AhBQ9/CUiY38ezwNK63J9eRTJgg5F50ViGpPcPH/TQtU
fyNXPLciw+dZ8BCzVeaCuMOSMSDMtHEidmokGLbgARJHo9cP/BEJvuoe9d1SqqsK
vcEgH/StQU8Rjz8bmXHGu9NXLh0UVgFTdRN0MxH+HyQ3NXhg7l3UtgkluVS2y+zn
UZkCz3+/Ypu42/z/ynV4LEEQxaYHKYsRK+0xcNEpp8Xw426kaW1j/H628rGqrPjF
+jzElP7kEiYEN7rT5czs6uuSKfVM2Jkynazm32DnQA6rIQFiP9HwmV4jjL4OwK1M
QTRA6S7US1dmEPGc/A5ghiREVU9vt/Z8W2WH5FhgEidnu+9Pvw6/qE1+vBCOkHu0
jnbe0q3rbFpNQ6V1IVU1Dzy9vpvPQp7M6ucGIdlYNA+mE2VrcOIK8t6JCjAzIa8P
C1ucmuHoG2sYpxTmAxtZIbYGxsjMy8QGNqQrPmawe1eXqZsYu2oeHj6lcZE5OIlQ
pgiDj5HQBCANnHLevC7OGBr/7zZSStr4EzoE3F92RYUOJZJ99H0wHgdeJ32Ol80q
`pragma protect end_protected
