// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:37:39 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
AxbtHvw4F98595KoXiqLN7hcVJNNLh/lQzHIsxzAyU0BgbMhYtzRTzuBr1lUtg/5
TG1iL7JU2KErMl7xnQk3eetkQX+bZEm2FHQ8OYgLBVXefCl14ImzZyNyUnEHDnTz
rokZyJ0mc4aWUf48ztMQLEQ107BENk2xZLKZgqnE8wg=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 8288)
3gLSCBCRCUBqd6f/BqMduHBWQV9H8jaji7NMzp79uunMyblios88vUkgTUwLourk
PDHnCc/duhnqjAVc52m5ukn1Vu4CnA3BtHeGbnaJHreisoXWEXO2fOB1DMqJt4au
I3DsYgJUEqFI0n5OvdCynF7BhgU8HGu7uKYiORbwct3z7HnGQJrrnYJDI1z2Q/ZN
rq+eKh4A4t0xdYgOmknvuKJfvzkj5NYo6WQcAPJcV217E2xs63FUdEiscyYDfr6/
p2TfK+zzmZtai40DBrt0HeALz5+WaWuCJGje5yvNqfrBDgJA7AiLNWSmKtGEBW4X
LXjLR2tHn84D/lb3DftM4SZmQJSVI3T+9jrGQirhudXcPvIFzW4Im1ebNgIRBa/v
VWhqAWxq8RuFZy6PIYB8zRO8uSlmgifaUjHenF3WzaDrxD4BVudPH2csK3FN4SuX
QHC565nD0AnODY434Jf7kD5UInGlXoohUcBip9VK9hlAuPC92xtdLLrpuhfHTcts
jWPh+Y/oF+sXV3K7QK20s+0cCyAHPdSiqNbtOaqYxTZm+DW7b3fl7i52ntknE54+
pJZtPx3nnMA3XWEuLOU5qtnf69dGV6zOOVjAf6dW/Mc0F+XEZenHosU4wNpyLsm5
v0kkuvjhqX6l8HdfflxwmTxXnuhCjeSYdPUWfKbAzIHK3Q0qsfUzy4dDiCN5IlsX
m2tV7KXx6jJLHc9K4J41rEdgmb5xgD8/P2L0JPsaLQDsw9BziaH7Iv8TxUPXtaL9
B/yOqW+HnJZhqF+wcGyav2LKOBgGNECb5JPBhp+n/7V467VcFPWgHQoMab1Ip5SP
Y9xCQZPfj/+MSYoGhS4A/Ub54aS6kzeyYPECoqEqK/HcVJwNAkJVmW/8OR20YPG/
zL41yP7JijTIFMt+kGsNM6dt/We3wlNP/gq2VPnWTp55Tr46N194LBUll2cwBiu1
BJXqtgWRbofMH3a4KFu1Fn+nX1YnhdhRfEN+sv7CKruFGgHEqEx4xOR4Nha1yOqX
eMNyRr+g2qldR5t/g8WMTywY7lIRSNfJavQmslvXRynsjcV8f+ONRv9JGiOd8HtV
xP9ugsPgu9uHPUbb8qBBljO7rujDGe0cmP5yYhQJBRtJ86JhOoz/qJvpMclhfk/s
N27tY9xvGF1LSP2Kn3y5xyUqLsQfWXny4nEzX0M4BkwYLg9OXqfsvWJN4/XamNKi
GK2Et2tAAmcDU82sA/gs6UB0p7HhsCTHa+TJOwd/Ptlvg029rKXIBtAwClM+q6DA
pV+oJH28GQETIdSNg1rnIP3Zd+GqnLbuLN+EoSin4epr3crjxhMAzRfaz9JCLz45
Jr1i4EoN3XTMGjg2CpY/l/5jSdOiTXCXH26sFryXTao718TLg7mCoZm4pMDCVb4o
ARHpJU4Ke4inuKR+/62XevASXS26f7RrcAuCva/vq1DAzXcKZ85BMwtObqWCTBJb
0Hb+RNUrlyKrtaLhFcJZ3o7tTFiG0ATrjCberPfHkaehwoJbwQsIrC5M+PjqD3Ba
Rw7yshANqX27LPP7cYVjYwKHoKsPHf7B4SJhg563dGPnl+WaqgPxX1LH8u1MYljW
ga0rgZpXjdZ0ozKv4F86rlg57U76stCJBCkfzuvcxSsYcbMLh/ixu6Dr/8N988xs
nB1sS/YkTn4CSxl2BHrevZsix0Xs2nZXnKl9sbMrl6fBedy2019Dncd3+LBXHRqQ
xcShvURVq3QThK/vAT7dNDUtOgtw9ZXvM6a1M6N4zVpT4quAK0e1RvMomPIoXeOE
wf107fWJ/xNl/Wl5ib6WoDW6Ki5xFDx7Csd50Ktna8QRIMlFM4XY5BJMsrsKyWBB
u5zdJHnaZjs6ckQdtIn44i5eVvHx/tN4TG3QqT3eZtBQLGqQn9/wnzF86zg44c7f
P7jwasOGv9wibL1N79akVyNtWgWXsz2vZ74Q1gm6DXpbZTrDp1tpwSAPrRbchV5G
XqZwukD3iFqMQeoIujPmnIbmEPHHhRwRqKdnDZVDmC0PD/UFgyIp21L8uDalu9JW
wIvpbQ8A1UZPRJ7gWX0rDnOR1qfDAInQ07fYGMIYJp/MJ0Ks8O0nZzJoXYbq6cMA
Sd0Yl0DXQndjJLCA0/k3A/fcUYqPREbwT8rwBc07ICce02ygh3I/ufmUbhQZuOA7
b9c453jpKylJNVGP3tlutcRWUuuibTvcABzdJAUYp00ax8SIxOkl0EepyaUxwRE1
txYSAifR88i27ziUfuX3Azq74wATPkmEyZI6++3ZJaUdSiJ5yUznvCmrG4CzjcW7
vohW9vJM8h8GmxCWGvxjCNxPV2Pg2AoIXBzNfkFugOnKoCGndQUzHKKFdqvbI17q
Xx+HQcWhWM7KF8fwEL889umDuqcbAQkLu8Pf5Jkkhspvc5m66pMyOag+ZJC9y/tK
cgUuTzRBnD++hjzi8rpNc3afYQPGqCSNLj8Qe6W8H0bDlAtEExeLm3hx8CaKRHTO
PhVH+w7n3vv52LfZe/QeZiDZ3LliNzpqsZl97uS/ykQBpYFWijHfvh4sqsF5URNd
25Su8Te1hS6eCIlCpHcQdlQRbw0F4qhG94K1Bu3Bgi/sx1cHiWKQEvF6k+9diQSg
P1H7aIadcudymeEj7H4HUwWFwuTnSZq3K/rpZ1E2Q4MPByIG7ys59h0aTyGlMdoW
G6otphFNcmvRvXDz3/Z7uiLeYIcgYXnz4w0iPxMrkWlVT8CGD9YqjleeZHEr5Kf2
FawCRnbh1cDG/3z2mBFs5rEWBkVQ3vKbnWjYnpWoNfPDjwgkaqqWeefdQNOiAeGS
tpMFwn6hWcULKQqyFGPPNIQYNjkCO0bpyvXc9nU4sbPUhm30zSJTaUKXBlBqEIUS
LDLoazVw0Jf5pXS0FHg//qyQxhcxi9KT0huNHUpDLfsCbJ4Qi8EuZ4n5YDcO7Z3g
Wm8b/7fxZS/lTjMuSwHm2fP4u2hhNXt7WaESpbFJXbCL2KQBewhViHs9Z+ymaqiT
AKm5EowzItXlMbnLxfucAHmlOmLCl7lCgIudD+CsbnCJ4HF0sXTMix/diOQmm0fN
ecxqo1K1pThgVAF+CQrEpWWsJtos1D1vAURKjRlX1CsfTfjd13PnUKQcRFeZ+88S
3hHFGQUDXPR2aI0pCUeNO0bB59XyWhNoBvssaf8N1r4c8zhY+aa8RkeHDCJp1sSn
BC1PEuIsG8VioCNRx71zp6Crzq9D60OKvuTaqyI/eBPKPgSDBiPRi/VSTPBoF0Sz
b00N7KLl8DeaHACCqcL7qiJNw+xaQmyjvHGiWK+4T7ABVl1A82CZhs/2CIWNxIU3
d/OGNgXH1kukWweuJXFJema0BYykeUgV6nwHoKD94dKlBTZWK1sHSniRCwT7Gq2C
D+cTfBOtzS7cDC5Zc+zK2GMz5Egcu/vjA9tKRbVpEDR5ixsvhajWA9eBtE1kuhD9
t+4aHMLWkSm9PwYNAABStvLE9MU+kCayyyxOJU32UNx7bcNanZ54YCBvhNfE1wNz
6MuHh2uL+iE1dpeU0cxeREJJH7+MaJhFeDtl6xqJR7e6p8B8jRnA54fkvyg5FwQc
ufGHd3yl087IFCteKmnRQjXkDQ7E1SENbjhGXTZZqJEjPxd7nd9++LVkeAmW8BZE
1tHa2gQ5oZYGhLtupeQt/fCmPjnbLErNwuOnEHK9/Mq9QdS1QTlf2dqNFMijZsiY
An/kBgiarn71ROzZrsY+BS+8gCe0GK9WXrSRIrYfMasrwahbLm94vuNqiVrMKb0W
2/teRU1uCPZY/qrJx3S66N5K/RWpTfyENzQL4kfH5FKp8ln7K9XXUB9Ms6N1JjnO
j0Zbz6HoYWzH3PECYLJ1ZwA2Q0n0+vr2RvHbD2r7+vCGBg3fIM6Rh/Sl5c6OVkG1
Dlx8n2DeFNXiLT1Rvfpo717eWWpI6iXHJeujXljzCGTWhjeI66IgsPayo1EV8cPh
B1eXRY8aKUiqx8eJrh71MpRVS83V1VzphdJbyLs08GUPnfobZkmiVqXtkhiiYQNl
ozniKmp4GrpwSTSxonx+ooM4jJY4nCpS+Y31ZmUojJ/aK/akeqn1kPQdYtgLsOWE
JalXkf4RhiFWWnG/k04xmA8op46qYSgN8bfnx3f3s6cP4IkhVXtt5LXiys8hu4qg
sAI0Nw4meZftAz6wN459Bf2VA7wLFKQgbNfEXQQpp1GT1X6rrMKe3mcLltfAKcDz
Oe85/7094+lgoVrAOmzsW3IxHx1+J/iIgFe/4ibiKxohpmJCwXS0gyuTGS66G7sq
na7sJr3EUYbOzyLXZFFLgtj7HZVuGNunXNcJwmwTPVmltacGKYHoTePNQC9bdTj+
ejBN7dRcqLdlOw1hBq72QAWCGuUEjdgzFP9I3BZP7+/BXXjuamPUBKl+BMkXS78V
ofuA6m16yOqPXoYEYm6va5HFrYH+tc1dBCOAJ9dg988Qt9f2wgRStvLCYjGblyU8
pvNGyKjbDCwekA3AetGwe7yZeZzxZmhje+nTvUzjF23EHiEwFkNmUWrBMj9AxMry
jzsS3qAwaPjNqmgChgFKv1/ur1HffJPH/Zt0efWilXTZ3XcNNkwOzZgrRttleebe
GJwf/qQwWL5BSJIGstjNCHcVm2jtTSL+BLRUpN0S0auZxniGoz0Fx6yRDxRpv4Yu
3aeEXviwnaxRAR1J1CspwCwhM5ZAPBtKa9hELO4EmDN7HeFY4mKBMHUWZk7JfLzs
Q0w5qnfZV0fWy+W0+B0I1ZnQLQIqPIQCA+8CdzP1eyKpyyefOQgT8N5IDWOEAVgN
M7BO3s3IPja32mO0umwwq+2/dwkcMiz+oJ2G1LJbGFgX2fCJglIO0IxXPqPffLGd
D37Q6Cbv7eMBrFLgvOa7FAIgarSWkutT8DS2XJyG9XkAaky6Dl3bVKWEu8Upeke/
w7zkWC/4EWz9HBr/qdJRBIOtm/Q9iBMCYxIWzg0QNQZILgyMlXChzMpgHxB80xmb
YTWgqE3pfRlHkfKNYZAw55DQDMs7P/mAyzD7fECTNu4r4PyUDEBhiNwYv+wjzycm
pplWp0QSbtyyzYNJvWoKg1ty8fORSuRNNFGMUnqcpLw9s0e3qxRpT+K1iPufZelO
hWVRQkBhZeRoG8pTDUkObbdqUNQap4+q2esVqoGkq6iAEsAUd3cjDWPhPeBbOubJ
LK9C2BZPHDDasMvoe2OUi6H2Xme6SZ1y3foCwFbzJtSHfqwT9fDfvfPM23w5hTHS
/Gmz8X/wOrrAdLd3KdM5AXWHvGyRHMR8UTwaILsz98lN/klnh9xtg2a5ShiSySbl
qU6XQ7F4wuHFqmLvEb0dB7eOMm3HcOS8babjfytBhL+CtmVz8ovQtF0C6isN9Gv6
ozVi9ic9MZGiUSCJop72gsYqEgo5C3R0fq/4xPyHeAPRJ97ZWUcC4j4wOoIXPzXO
dNSvQ+dsOZ8JvOFfa/uuBLpQ7K9S7TBrHar2xuxoj7Pt14FKauCQIyzSOhvxs+wf
9LB6Hv3CncWVvBZqZjGHr4AETODMPL1zR49piHOTj3+XFhgqbvew9JiYRNase0+U
uSFt51GID3ENsHxW7fq1ExF9RP6Vlk3IODy4/kfSverhla1B0Mh7CZ9kL+PxQG/s
G9wm1PxUYJrrmMfUbmJGcxU8PdM6gCA7WIYmIP9XgQl3sPolqIzXlZ6cjLrrg7TE
tWeGRqRPtWoQMosjmIH2y3rmhUBoY1MQdzkwnqJ/ENnwieh/VcA2ZOsbNBXzcpuo
fLC4Ayzk/pgqQZhUbwdttJQVH/UiXeij+4nIiFSLBf4VEL1LLe+Ekq17WLKHZHsp
/i+pJbQCYkDzTo+YvuPXuqU8Lr7ZgReCrX3PitteTWIxuLhRLusB0rZmgUI2FWCi
8l1bwpO+oxp0aeajfJqVifcbXGEeDL0SKgvAXoLJEFmZ5FGKWIN2xBYbMmtb4N7J
jyziHHdDh3EarWe4BNtBCBc9ZZAG16or4GCqRiJiGGNTSVmqQR7Zw+zJVPQK+B4v
kalzlfaum4KGvLXPYjH9QsDcNscYopxFJo8zKuDiHphU+R7HaMftDrxNt2d1Henw
ch+UiMbn7BaucnzzMbCWucvjCkaol3ShPGxgz2ojrWVRXjdVdpQuYdloS8DMSi8s
aW2U74oggKO9Ba9toSJm4OJdIT96FsuW4jPy4h2kMz9IQsBykLQvtb3E+vXDLsrx
Qb+zb7pgFrRdYSfMlROnHVYVCVqx3nerZ4ZvsjIdiR6Njx8jaCgoiL91iMvIG+vv
wttQxwPmseXRMweMebSm2d+M4L3eHqkhSn4W7xz3IthHxUDx2W7D3+Hr5PuEFq1w
gFcBJK3TR0pVju2/1IbpFw2lnrH7MROHBUXc1fEYaSKjJkayvl20lOHF9hO1VFae
o3q6cARspbUL+A0hY2jWW9qPSWvhP2yrfnPRrVWiMwA8v2QVAH//Tt9yVvhaVJgm
ETw9hLMynEkcWdKFRUOJHA7IhMKyAOVVaMkt0BIECikX7HCw8gKjR6srRHbGMg0Y
c6Flk/OR/Z4+vA1T6VxPPWAqXi5bOj/h1BqRWU+n1+uaDvR7Ulvvdp/LZrJZxoQj
Q39RG8jT2WhSY7gSPKXdN2yl5SZ04pqSES0Qg2+epiN8XGPzs35jOVw5W/F5GPcn
bUY/3hVxejMOQYhttMw930XNglyKEQ7g1yi+TJvf+xWcWVZlMfAe0dbgar+MSdtv
t3aLRCbzkMWKy334Mn4OoiK+cRZB+zejiZrBxy+MK27n4VfxI9um0poiqEkL3mIE
XhCSvpQK3lsm4kZgNe3h9r9lokPzSJZPoVS7o6IHsW/THF58XOVhdkFUBBaq1auL
nnEHSKolmLw/hFrRtUC0KvWVoe1aGC+0Trd8Q9U0VzEpKdBStfomsf/Q8oLGLEkv
2v0r883wNUbC8zml3N9qdq6Br7yXr8nixlfEDq0dI9ZsniGgvGb0RlpGh62xQIuI
ozp47tD/TYCuzhjVI78ZF1WYo+J6pK6Q/UNpeE60pFmjRp5qKEsTQNjIZPCoL96E
43TxNB8IvGWl0PKQTbhGhDjkSXTZKHUqAZPBu1WjoVUWw9bR+jQINuf2CRc3Gm2e
VjH/8IvjSNO01F7dpDhFaS8tOa55mZDn99F3ombMgmm3Gs2WBGH8rUknAkjIuP7Q
5XHowggyYEib7/+3wcJVJPYEEyCulwGsownrnedlLTUfk0sxsBmOfsbyQVnekSpU
R4rQm4QS+r2bJURaURrGx+FmqdtqdWLaV7T46DW02HjX/6z/mH5ZuoJdZGH9myzK
Sw4TXynJjnoxUsZ9tJE2ymXjaexyOmIRIo/4UOL7xe+YB9OSjoQ8FS01WvAVsSRv
tVcyVIoOUWUD26JKkSJICvDcozg4bG/xeuveS8ELU91r0doNYhOSHeUanfKt7Dxr
TDL8xyXSbYXQsdvupDhPZ203eJC8Rm98Gt7pztLpDZbFuTRBVjHg79fNjn7g/sX5
KGfGFSzlh7ZwlT2NMtiGNOw/yr+uVH83wjtFOemaBqKAqiEKf23XGv+pVvOaH2hJ
NlN6pK48xgpUi8VyAa9enRPCBhTyF5IP+85LFaGeAYZ1FJg2dHJW1u8DPUIl8mVa
46NKMMlRgwAXpA9RjQhjxq1vrevn1MyrAM80cLNRxbLysFzmYw1CUYaYDIXLk2E8
UGg3rWdfskHzlIh5ByTd3jzXJOnWT+2N49K4H17g5sAfg3ZrVPmjFyK8eJ4NauGe
8ryP/ntDHs6wjr6Gh/OePoiIZtC+L34+zKk6ddHELW7CYOcLiTqpAdelgVtCx+Xf
pbDqqfZIuVn52mMMPJ1kNnkE0boCGyJg+sYdPEkke6iqLt3qlnMCdqB9C+GZXX2S
cChtxV/j9KtTUgoJJ3yz0s6YlEQjkg9nJjscMPZrJs6ysdqAr0QVR5h1LVr+gP9h
YLXQLcc1x/B4vEZ/vPANZUt9otpkuSltNXIbOgQFN8XVbvWFojYOCrNbirkowal2
3eN27ITJFlMZU/EcK4QwTholO2/oGRcZ3tDQRe/rfiyHD+eKXZOICfXKltetC8mB
KcXhohMjBir732YR+22sQAf0TV4Vae/RkAHX12n+vnhQAq9nH3PN+kDd8McGPMpC
IJM3NkWLRFOUdOJK1B46PqBDV4h7YguN35Unh77fI7tVeIjGQHcEeu6lXixnaXfB
IEtd+woE/zyFPY8YCCI1cX/xTS1PvlypKSvkE/QnJ6xhqz9uuLC8H8uLrQrwAUsg
U9mu3XDhcr1CKfRw01Y2IBTPY03FO0G+/7ShwDobfjWdBlzFNXEx4+JxBNeP2i2B
8MkCX+ePBC+2EGn8Wkk7uFpXnpgKlqEEBzlOA3vgmcWxkfOOa9gRyJWnvg7fmitZ
H+d9OmjlvwXQi6d7+tjIveo690YWIRPymD+2rDX2MKGoykN8mFPPZIxo4ULRSoeH
4RacEEGivODlvVUaWBOlaBnZ49WjH6PA1J/XcC/qVPRoebHsXR3CEXieQEUumAs8
2rrYywZEJGmqxRO+ngmWV0QqmMN29q8+oggJA+SfMYhbjWOPjbRx2bwBKbj3uPvT
pvtFabEAHH6oSL4Wnz+4e7XETkDc+oHz6omuM/EeE0UoslzG66IDsoSzJHyvMtnR
dHQDahWpUU3wIzYNsZo90rZH9AuTUfo4dNFdxDJEncAGsD1uo8s6e4yM79EJfUVs
J4Rty14tivCysu1uBe51C4NWeC/OkRpEb2KgDin7QpeEucvy2wB/+3RkJMukp7gh
sXcodz/UmH3Q8zvPpvV3bbCxvR+te8VhDtAWzneA/xcujUu+tXG0aluiSpqKyUru
mu6UYfAQFZcrN7DevM8d+JfM6vbOfi9zGGytxrOo15hkdCOYyHJhVn7YtdJ+bn5S
HGV0P+7IQn1usDHx0hMclYIvKFHSeVP5cLGYFgcDMw1P9otQOk/ac/wJxoG6vVOU
7MAaFl7KYsj9fPiH4+DS9jKpaORnMF8VkuaeeApDCWbBbAwz6myp/E7l4XdPjM4G
lK7ygEktG0jp+1H9pRQABdD/h62jqpB49P+elA4LWlbD5k5gPqJYF0xbWce2WAUM
qWcck7iCc66MoauL5oe+hvDr0HL7vS+9Bd4PrUaNAeh31MbLYK1/MbSbl3ljvQuj
F369CuLlGUkB44/zX2D+Ivj6zb5wANEvy/oNTfMquhx+6NOQCkmv7fk/+IjAbOs1
Mfs9GEKrEW61lSykCtqqSnosN4vu1sXCbJtBfftXxg7ZYhKp/za8RVo5GJWHxxvk
P03NyBLJSDmkd265/emruSyy3e9q/uV7UjCO2RdjoSQ9AHM4aM/uY2my+kAlLQ3M
l1SLMq07tcjMgSgcFGvzDYA6Aj6FIORccXbO8vp/KxZOjQ9l/h+yx0So16w/Yz01
vv3XZvBKjp2/XIuqq1CmqES1B2OSt6JjNzUYCErBzkvcnIqQkvPoGyohArhUSb5Q
JeK5LcH04Eg8Bx29Tzb3ZhmN/gwaYud09NDybpGQT1i60i0tqSVEjrj+qJGr+lS0
5DXAPSFah7DiGzLRKmtgDeXx1NIfSg4Cg2VYagdfl2FSsbTLsJy9uLup7pvk+kU2
bO1uQaF3ORhyjBbempv5Crs1sRwkz1P6J7EldA05dk3FmzWQxZCkzCXlkFAyRWWh
9U4lP7Q+9a+IEd8QmCl7eSBL2e8WzJGO/GiUfmnnQ6S7R3mz9pFqLdxXYNc7EKDF
AP/vBdJ/vZgLuK+HOM2xSFzb+ZzJp3/a5kxjka37Gje6EAwq0LrQhaYH9skWQpG4
Akezym1uAsAZ9wyfiKEDJULA0ogNv+M/fXvlKXLDO9bzFk5VEAyEV+kNhnuBe0pc
MuLH6V7inyiKLrYp748SzunvauL+Mb0PV6FIhzUwjq+LN3UhUdcDxiEw/LVfGfq8
A/eOd3UAw1SeX4LfbLc9v7edykM/iXFb+D6gKXgL37Pv5dJLEh2Jhut1ue+10RQM
v3miqpEq7VALkVmaiFEdIPeX1/0Mk/XjCXSSgWtGSfOs0uD8g2DcQQl+4LY5jqfF
b30l9xdDxRGw7rNtH1jZTjpcmBkKuDpfsF9h8+lWCWlYMajeNonB7h/idGSlcDGi
jD28kLUL1AqPgO9JN6IeO+Y6DkCASuAYp4NOz0GETjAIztK8K3CbQTUrjbVK5BTB
6vg8Joos5/1xGJGSNxeUzypW99B2pd47Fge3fjfy0fUGbmMys197p6v35VhNXuXe
jRIL1owBa5M8h3TDPMEKqWvW/xKU1pdxP7X3Scg7Xh0sZ2FW9rQLFJLH2/HbtQw3
524u6lBoM/qJvy7Z+R0GagJaPCrIrkmxMfxdZ6CuCKWbIgzjdW+gbZ+hcGHyRQDJ
DekydJ3cKW72VaxCA5paRtRr9UvQoI+37MV3Fecq9AaKk2vEfR/iznF63zLunkcw
ycwuhjs9D0vJV+pbbtbhbiCdBNvC3ceC356wdQ3QrAZzy7G7IDXS3f1CFJgc2zYD
jW+9fsAFdnHt+yz7X+JcEdATuhA69HhjJjdz1Gka/XhNps6aPxc8OKAk1NjdIVVq
MA6vm3BTA3sm6OKs4CuaH/CCXO7z1bBCCy4MPfigVVVI4riPhT/XHRTDnEeew9/h
r+k1n/3/U3elQS8+MbSta2Bm2oEMce89sF7DQASz8G3av9ST4EslhvM2X+tJTxz1
tVt5ZMu3PJAWKpCgj7zZb3oMEztItqjbSM5bpjerWFZpP5vvgrRMFi0jEc+1PxJx
9YDD4843wmDtUQlfiYO72nm0UqNMyDhKRUvxYH1QgQthQI/eH1zY5sETVfhIP35W
p3/y4xZa4GN5ELO+gSKhHLpG5YKoW/ppiMPKbAsNVhXIjN1mH/X6VR4JGB9cQktG
3pJqj8Al5Ttlke4SqGaFVAmlwbMuWzmnky2L/x+SU3CreIiPDz7tqlrbEW4Kfhud
KMY5EoWHBn6VpwHHibn8FCxLcqrz9UdSaM7ghuMaTmJEljnnHIYQMLxrwIIsRxq8
l53ZdJWsnA1b1+X0T9SuwYHG5cEleDUoITelMvHpxKo=
`pragma protect end_protected
