// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
Mew+Z1G2Nb96ncqqL/My2OaEYLeSbwhqgwLqvQAXx3/gEf2Mhv5Mj1TW7ag6+CdQrr2O6Yixk2dp
SB5WQW6f/DHEheb7Ory8jlhkg4A6nfLl7lCpRfg5VipZ2teYiuWY7kqG1tFU/jY4dQ2vMHB0BNms
cUp4AVg0u0xIzDErXitlFotJTgjaj8fcBqdnQw3UOjc59GzQeJnBHGFpkXpAJqG2pI9ZSrKNsk5h
KHMInrKwxC6ENhm9y4Gn2m7uqicgd5IuVSHg1E36raQGHwzPJcdGkEZUKmezfxIAd1fRMvNwMr90
9zuR13l26g8PWX55epT/MsdQHEx4X41FWkdZ8w==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
1ohFLH+lmQL3km03pny8QmoukpdNZe/wzw1Sv3nnSg9ExROpPDx01oIzkzWjdVCTKiMY28Rv3VdW
yRxVyH3mJ0+WgAUFe7S5/OXHW8JeLHGJzp65NQANa5Oi1TdzusvZqv8LEgIjBKq07MNq2x2b+cKh
bl1oYypviWGEM9KGQ9I2SuN1GoK0cmwsuWFXW+Y7RysnOeR1eDTFdEgHQEW+jX0O5+eZg31ZP3+z
I2S5E+L1qYtKJlwyTpr1pgpImkFMh086oJJFdDdVBQixeG0v11LJA/r11J2G55XRj7l+Rk6r308t
i3tCMtpgAgBJjoXqie/L/IQIu5jbcffyxy1jIy/+qzTiD6McXitutZRiCkuoTZYLc/Ba5XtpcdWQ
fpa3BL6ZZUgMHbbXu2+jYZZxOn67AJ1OFJ9hG7A/ljNXwat/8w57ySeHtggINPmOZqyAkY7uB/x2
2yPWP183xBg6sRDTz9y4Flez25Ib4LNjlHHVrrGin2jhM5zl5Z2wF+PF/3vpeUPZGIgizhAyp8iR
PSkLP2aG8BC0ITz8jtBNIfwRLhvHz40Dj7K4Mqduia7lZ3YEPQY+XEWfP27n6rQlkQYGdd3wwls7
TtxO2ZyF+2ziV2EXq6yINwSOss5IGEx1E5qlgoQOD1bATldeZjGvi+ueqj/k7jZSq/1Rlm4bWH4g
uwIpp703sL68qDfamCo+WKeiNxj7HbpVxJU/LtScUAakXgSmr++oMUmuEQhZu8lh6xvjX8R0PqWG
K8Xidit9rVGUknO+UBY7H9hwTzm+39dIkvjo/Q55ZUPZB6navCC00ciO3VelyNf8upgskohpiitc
0VC9MqBh/vMC2oPUM+et/lVnhBiN9RM6NxUErvaCckbevOJ/L65gMsfacmzg41i30AqJxvYZkT1B
VfsfrU278eTFuZH8UelKTCyy4hBfGan2vOSu57qR+owPho1hdNVA0CRTT7/TISdjklNRCPWDvi46
v3bUCu1oQvGuTQPIu6qz1BqIxg7fWpxSr+zEHuTsqRR8kKEGPIULvTvaWs0YHaVyfyI4LO82vLmt
1ATDBtd4rTX216ytzVs3un+7q7C5qksdsr0g0ob2l16TKkNJ3/P12rwgH+lKuV3evf+yP1eTj1rR
ZL4sjpBOYhaH7oayj5egHOE1UmTF9DrbZr9s123uQGbctyzXnlq9jJet4n/8KGLAvjOrHkyx5sKc
FYij/JY9hYyqy5csMp49YY0pHHCXivOfIL1F2Qt6nwadO5SlqCc6E3vfTKez1I+LIIop5be+JGri
tHnqMgRcdA2IGs+ymumwMWjGRHn3e16xDVcw5NqYTo4qo6GoaYOTpprqMwFMBAzia+sKCaG+BzxO
OrURWnOw9cEV+CALWT/LHfFYNSHFNlmnJKt4iaaBA3B/q24I4EQyCcf4WmuPNDXZ7K3QrxWAyPfu
CYQjBYWN66HXSj9SQmFtND8vdwb3z2dBkR2BclX8C58/Hw9EIygUuWnyw7SN6nslkE6ldsyG+m1+
GgdNvtQbI3h9oOCjkIiPaBCQe47K3EagV76tvNIRshey6pY+103bfjxDl1qHIH5w/B4TJs9YJRaT
bfKVZX8q8kKfxbOgadFNuUVLeOmwhizk9HYwiXz7XJGYvCVuRUcUDhl7BSJGepaMJHRcIuEZBk7J
hNNrv/pudlfvIpnAj3P/vE92LwU2fk5WTB7g6iCsKKs6a6ruP7CllpZ9BwQ69ZiO0k1QWCW6N2w9
xntZFEgLZkEoZaRKP/TRfJTrUZbtyGD/1amrB3qLJ2sXKm5O9PLdv2bqs1GbV1cJKoBmXGAZ5+2i
LTzwvNveJAim19LSpHFqv5D0Swg/U0vIdWK0HwWfkN30WWUr7VXVOjty4zcO7rq2Tn8UlsHgD094
XnjZBoMlF9N3B0VuhCx4sfpw2IAg197XHBlmhz000sns7kHzUVZo6dxDRyqu08D7UDi3b05DJa7S
RFG9KobKQzGkqG56Ksu2/3kzuEZpoW61FHjm5A2vzv0fnXR2W6t04opU0yZERuCWqdu2GWnAr4ER
kpa7fYwqcluMmIdb+VTUzdDb7+6p+pNUr91GZtvsuAJHrsegxj4aqB7E0xNonOlRhiat1ye8Tr5q
FVM9iLptATTF5lq18vV5XqxhcCpg7yEyD8Pf91p6mmt46SQKkAGR+ISy4sndv39i6IwSYAv/NIoB
lKVxHZ76YlZX6ko1COz4yRf/7a9KEIEFtbJpFCytt/FpPSn1FzrjDN1z9BYjh5oDI6SSuDNeOhSq
4AgPjywMiEwXgJrG7JCIRyzQnKPQ7/8rLs9sWaKnCNkDUm0mS6N284X9gTv47KxYrs7j3XmFwyLj
0WdxpDFeMgIPuOiGO6Th2t1sfJiFtLU3xqFqG7sCPhOoCROfkccdvKBSp/D3hgCXMQ4l4Pu07ExO
U9o1t6JlbuFB3jbfciAXtJ85bcPZjtl8/1PxOAGp0o7Z/onX76M9/87YMf85QS/NypTfV4jx67d1
DWfL/mwq53I8phVEoUKOTvXdq3CurxxuxDb09avG2T+QIv95DGUrgs9moAGR6sMgyXvk6ruWOpMy
OVo3XexfZSQ9l8J9SO5qGU8q1FBG63ChWCBCfRSxderiN/cPplKJFuLrjKGlDNo8goMbB1dSWmRu
uIaS0r2eXEpXnng4LieBsMbKyaOBQ7ycE926gdR85lXVlF2iojDHaRM+npnay8eOXs5rEKwR6nw7
JQll11LDYsKcFmLhabkWiOIZc6CHD5JBsZ0z4yBEgdad0HY6vv34gT6oshYa+Dl+pFhOEFVdQXnt
XeKQB+DKLJSBHobSFQ9PA4SdWnOjiTQxvw/OJpZ5i8aPLxldXLtRAheKLBi4qJeRYcVGWkZOgc3T
ar4sIQK/Ibyhei7p41EX/jZjzGz6zm8CVgy7QB9p8Dy9Hy88eEBeQPDi0dqbchnj07bDFSvYUvZJ
rqqnpiE5Ja2HnxCEuue+8SqZuY+m3zM7k9Ns0tYoL43E0ONjGpDjl2+q2n+afvQBta9lue+5ZKgC
9zy+WP0nhRRDFRi/RLlhpCNzNtz/8Si8gWS6365iqh3Jy60+Yqrw75ye5BR16hD1ZBKyLcSwkjwU
Rh4zpB6oq6NrMpTrwrwR6g3JDjjTp7MpVfQlBAYOjVh9+XGIIWq4/Q6d7hexyyEaGFZ7F6MgHZRR
mRuDzOqLsVh8U/SMt3SVD+z0D3xE2mjQOYzTBny95gfTL227EkR0QHrE3Tfcl36b5A1zQuIjDKzj
IdwhCFsV73cA2jMUj11O09wGgDITRKvqUbRD2g/42d0GgqG6on/8D7z7UPqT6YFfZT0J5o0NG8YV
antfcY3LgMf22BwHz+KAgILuliGfYizx0zeL+jaGKcVkXOExccC/NIQg9SKxJwkCUUyOBel1OmtZ
txyWIIwEFM9rhf5sRz/AtiPlUAHtYB83PYcIdQqZopsqnpHzUFDaWONaQVoZfKHK7QHj0cmJn4UN
xiY5I7JasIUGz8al65zuhzrCwSsFJRp0d67pvUeGjMkg05Rever/Js6l5tGGQDE8dp6tb4ELdM3e
5zTrhZ92/6AjM//4i2L6By9pEIvCaoCbocOoZ6x2C+LZD00oFNeFXoMks3GWIY2THBPap56fYem/
/ITjPA9Ic6AEB8WXfc3Q3oHVhuFTHpIV8m9Fjlmu87zGKJ8/qa1Nf1n643cUZKqc5Jpn1X5h1uHj
nirD/dPrJzDMLLrJb1TMRMaiATMGlZgVxoiysv/ir9rk8eQ/wn67j+irpvFHSWA5AEvow2tXsuS6
HryN3Xk6Y5uB0kgit+l3gH73SOn/AzCTOYDwdqQGFPbeJxmBpqs35OP89bwVGL5cJ2fEi5HKBbvm
xdiey+rMdDPEk9jytmm9cSzbWknW6MA2W+DB9/zGRS/rqyPWNLwW1TftkgWU9wVA9wYOPceoca6t
PhWy3nIGzr/JXAH/Vhs7ke/wXEMu+GP7IayYVfAH8SwDpTNUP6yuOSA6riF/ugfQbhlkoInwPfuR
GuDaRsGRj/hJmhr9OM6jreLifThWy+aZsDLVpVCF2r25tanBiEVf/cZiM2O0oy5M1XTbcp1x8ofl
jpnwFsDHPhePQJ4KSNY2o53731bqrwhrNxG+ZtwrVBwcYocVmzYD/FbzcXsN8Hc52EnKpBWXN0u3
hsBtx+b+sht9Y3noeSZSFynsyvljpMiip/PcEJGiC9Os0XlLuQlVbnX3UQCfD9oHCLtCK0z+NCKZ
6doNmJTkBlTWCrV7kGZ90fmUYXzegbMuSp1YhW4YtSBuW+sFP7Z4RFG2QVUQ1lcaWTkNuImsulMG
ey3rOaH7FGtlSuqKuy4Aoj5Rri8KpVeS3TuP5VdOvpjDfKp1Nrh+UPn42PcOkFvGvnh/AkRZR8BJ
qHPpwSH5cl8c0hiPHygXDoNLzwx2t5YaYd2QsThBnEnmJSx0qklyDNvL2C1o+tGaoN5g4OMPFBg2
RH/avJlvoWtW1Ke5XsOpGyy44aGhfDwinISYcpmGNMV+Gj3dUfkTkYafAQQFTUZ+23yhz+9q2ZbY
MTpVK2unqg2xjURhg/wiY1DCApYXD8P1K9RtswdMHfXNtBbjyfVyU/hsCiMGzQ7KFxPsFPLk73TX
gjtrHVNdd0gggpqsentn/jQQAWwN/LxTYYYYZlHNVuNvjy+SpFgEyTSqORVgLfQ4OsARxKucZnPg
aHF0AMcDN9ekef4IxibUuncaONpJWG1DgAJ3UPIzkeO0HH8SGnOww9CGiFToCb/7K4sk/rtztSZg
ROS6BXMNf5uOFH2kygmpK6gYYZYQQJqjO3I+RcYdJ3QIQopx+mpOS7CBgx1YPytiNhkubF/c8hh9
oXmTyIqZ1JK/P0n7kEBWQgrI5RVVAH9i6E9FL4kDiEaj0xsYFdboDl5ByktuNoLMOO69vOx3HV1j
mPIT7jCexERc8zBC8XSrOyDF2VJdJQBxLMpIdyc1aQ0GLl4zjWjLTKX8tVwFeyE4/zVO8P95ePiN
auUeQdGa7TQn6C78FR2DHa8B3OIOnYH02sRT/sIlurLppLzgJVT4XH5SAZkr6j2PD3nPFcZPfw+M
ozm2kQNjM3N7kyY0CHiR6xCFkJlsL9xt39Y2VsCasjPvtJCqfM4e6pmB9+DZVb3Nwxw58gKTq6f4
C2/nihZWQboy3AOEjGwY+ErLMVTTk+N4pxlof7YEIsskqGar/iOUlncgiDVO93RqqJTgA3x88PWV
I/IyNrm6EISD2qFF/oZweqCWoL6WTjzWS2h1EjXrZWTMns+4OvHwIbv0x1p/paBZZUZw8qKsK561
pv1sNeYabA801/Xvsqb86jJWjzrkzejMFfo9cmjdwdn4G9uUKBfzfVJc0gHXvW+J1ChA/Tkq9VrO
7QuDBKJ5YumjEZ10I1RnpknEB6GiOkDjH/oUpibVsK5Bma0ipps3FM8ak0FSQ6QFY9zspDT0Aejb
nti79uV+cLp2Zm3aqIOj0rUFeo8qooeGq66rlwfan5tZXScRg8kGQox6GdKRUATYA5Po6+5F5+OH
gICqKOaMJyqGEGM6rJW9tyI2ig6mwzi9Ptro946bsZDTDTZZL11lc3XjAAKZvRrv1Y1UQdDaYK14
mXGAfcu8oyE0dNy6NWK4ByJ8o3gRz/rUITYM7ItOES/Ia6XHIKlmaOeBEiamPYg3faKUf46BA/vT
om0ccD13d0t1b6E6uJ3b3iqxWIs6/HylhIHKjfhGhHAk+W3JhqDBEQd4Ug48vYX5XZXouWBhh9Ne
wgXsKEbaBV4B2ukkPFloWPPy1fxUA6PnhgsMVCnVdn8KuubYyZ2SGp/W6vZTDBBd49MJJX0kmVO2
uV9PaYEiXdZ94znMeZ1Cwk3KDWqcXtkBt+LwUJ/eF/6GyOLALNbaQZjJTujbz6+LtvMQAYGR5uw6
gjo0ZS9jMbEmu1ZqHmnc2edu5Fy1CcFNVPSw8DixPoj3720fzXA/+VRfMQaiQpuhrsLsEhiAteCh
8UT4t2cmhL1cHN9iP4DXCPlAS4dYoTb/z4ENm6HICu7L4e4nF0pSPWDN3OEU8NdjqSq8YNouHaCu
CFyepTCb9V4wj8ztmA4nqCrhUvoJnrX41y3ufBlP4FPdU3zgxFXdrTlMin/0J2c7+6fblUIXrV06
qv3ZzL5UqmQ+6dL09IiyrTyycjMotE4Ci//+vF8diOw38e/BYzSHgxES4Ng+ThpZqN61WDTe/TRE
C+M4vRauTdfaS8Dn2QFjtjt/SctpfCTEcnx1Mh7qiY6XCDkmqvN2Z49Zi4LOtNXlMl+m1BhJB/as
1yw2sSIieZ6RZD5ENLQQuDmoCfx0UVtciRQpOR+L7Iz5YBL44wYOq6yitt5dLWuqzm9l49l2IlKR
iVJ2Jitq4IiOlgnpUCYvHJdwaaV58AWCThm/YhSxgaSdpb4J3VWEXiZZQZmHpbLI3nzwb8tkUFVW
yiqfmdOqMtv77B3WQ8Mf3DYapfYX/PZD4KsdtlmQ1d/OatSTzMLnKUrqvaFUlOk2pxamZnQN9bq/
Q/ONj4zG5m3qV623Jxjd9kPKbLALgA2PkWhBkJLW0dfJGiNuNWC0DkNAicHJCwSDtLNhqmrGsgW9
GGo4QtvfBdO5yssvxLJqNn9+LKHkoVzc5C7FMpcDXuwjJ2GuEZffbVqKIfaTHpzjBnA94dA8D8OG
vLYsWaIit2U4gqu1UXQPgPT0BbYVBhcJeVOdZyZMj3A65YrgXGpq0pwv7tDJOrouWZO38UTQYBZX
43jNSVkUzFfmRlMGAdYPUT9a4+8dkou2UynIOEpTfd73vUKcES6/HG+H8Vsbuy8pQnxP/loqOlTW
8Lx0wFQDFoudz7pgrOe3I4LQA4+geNB/hBFF2eXDxs/j9P6BWfOVWtCpo79eMKhf/hB6tAhFwfan
CMhQNIVgqUQ7yfia/V+d5IKsmBYTMPvfDYkSJ//kgFXsXO8Mngp3rHGsEPUvf4zRXZrFJ+QoLWP6
Q3tGLgFglrbgMmeDBL1hhtUkWunpJN2t4JkGbun7TX61AxpHvhUp8oFzy8A7GS27TiIfhmxMWcIi
CCryqQ/wFQm666TcrtL3/IoPd/GGIbANgp/QmaVmZDdl3qlzdoJb4Sd6mGnlacHTBc8ErepIgSN2
RrzHCT6cA0KhYpx0XXIJf2mfeupv2ERT5+zQ99A2sCBmYXinfS6Yxazon5WBPD9xGFEhqGhyluJp
h3E3efeUxULt2w+QicM0C3BTpzyNwbCDQ/LUxbt3i57Tb1X40LpFdVQ6ifQ/rwuQbsEFPjYxMsSc
8od3bqanleJ45Ox11OICo/7jC+gO6Q7CJjVU7sGd/r2ZZ42FU23vZq7dZIaWr6B1Q2dHoS70tVQU
4yr/dH32sGgwuK/9KtkxnC3wajrgaHb742/ARgYaUvXrdHgZE+2RbHZVFO4PAiFnPtTQYAYD9NMi
dNlJdQRj6PjVPiuMZev2ss7VdDpNr+iaRo6vFdm0W8jM7wpHkKqEYua69Kke35BJBiOetJIMF97H
rJhpxZ6UCsTqOeV5RsNoHcC6Rbxm+u0F3Ax3f3ETrJ7DczNnJlzz+2yoITZg0fs8ylbpNr5nhBRD
7P7nBW9n2BCN/4QbtEzoh0VLBj9PuFqC5zUlMt3m1BRvA1wThHqCz1U2KAdpmfSUhUnc/udJS28X
HA1CfuVQtWK/OrPnu2aH8/ZOpMcivo6y/NVLlcEBUP832CwRLOIq2qNUVcmNDaQziSRzMM4nDdmc
eVtSFFXLCGsav7APwNOyWrJ6WJZuuHgVosQZiEjKZVaDEWQ3IyoR6AVQOmV1bwPXBq/NdrN7Gr2+
AC7ehkxualya3uUCdq81Jxo0XgeaFS5ATz5vRGLb6jtBpeKFIw7zr6Wk4pJuZObB6owkLuvVw5ZW
8BZ007Rp/jcrIrzQzJZpXzQwLJcejTkTJqLnm2X6ylbsJDpMov7+fKjnFsp6pnEzljD2mEpri/EB
HoiwJMRK3bMhZB2LSXYKqOxqufF25vFVhhNnn/SsEjgFXkjaJI6VPCUwbehWKVNfOlH86Rxwz3Fn
u25f/eJt8OTTOIw/cUO/WopRSUwMRRIvGxmpDI8KRiZ27U84NSngQemY4EZ8lrfKTFjuFmSoANtJ
DyFL1eE2wAE9/zENEy/MPOqhASS7LZsD/JxIjiCi26YpPwLNlvQPGwXQFJ3oqfy2Co/2yuPBvq7q
5k64FyuNVeZgsz+pBZEM85wcA+xdRLcjWB2HFFmXHfK7V/F5shrYsRgojiEBaPeMsLHiMdF/TGxj
Tjr0QIR1keWXDBUMpPpaemOVRBGEnphMcsIUxGY1jKLAlveJ/C554awQFY86v2KlzC2arXKZojcj
1IKo+mvWtW4/tKiV0fMgksqaRGbNlZ09xTyLzua3E98mva+/Sh0pub9/KvEXBjqSLBFVQxUzvLKS
BvMbUxM55NhoGarPAXFM26b4x1TmDDuxgC+3jGPbW7vDe+equRODumtddazYKWqQ3leIWv4K/C0t
eIeudRw6W03EKCXQVnfWQeAa7Xll7wf0McRkv1x085WJqwGc93dzpryF7OQG1d9jfSOihofByueo
rf3yFCayvDG67zbibVihHwSbVHHs3HJec+i9uBa42mu0fGJY7+AF1gJujTY7WszLzqOIJUm5ozEt
3d0vXAqZGrSaycBpfyn4DCW5coNnfkxY+99Q9zbtJacIghxdpkr/iLF+9SG1JWNlNiKY0/JOkbM4
2p4MpcUv5ZiCL+1kDhLHy8WWCr3U9PXLCNM1NPFg7rzJ5wUeu+667NP8ypdRm83xkx0HYyuk4O5/
Lo6jU6lQxhAaOoaK6il0WLi9iiAG2mYVe1neYw3YUhVbEERd0Kem2qNrmpWLwEM5Sgje+dc47F86
+XpjoSm/LjOk7WytcBZtQaBgPF9oukRRlnAuE+KyzDmxUUWNu5SFpyANyyTNcws6h7W14clETOaV
X5Trs5Cpg49A29lJ7/s+Ra57Y1WxivckNC6XHowXTdnhHHCM+yD0V81tGTDNu1VJTuofN1RpkxgJ
7avxRF5SML87zqNiIaKMPsVfoXdxv95NlaINb/rHLLLNaBUykc62uU4HtcGh/7pFtqMy+EMc8as9
h1MXGtXmvLMLigqU5ZWl0ANKAOfR3Y9KYdAt72Qm6QUTcZtXiAtxtWVwrECR4kY8OQ0w255u5Q0g
2KfAiwD64eSpkGBFs5P33RxaMSMjU5zVXke4CutA75P64NhsuFKfrRgjN+AtR7K7IAyRbDS6VxrA
7h4mLnqmR/iMAqrD5CN+5jdwVjrNYVUOCVE/Eq6QPHv7L5LR2zzcecKKdysnogrJ91E0I/PTiic0
yjnx4++IMTHURHHqAhjg8zTHWf9kuJN2l+uZwFDx5DszmlxCHfDaWSgubKCjdGuBNIVFSK9Mn+Mj
M6nc31QLQ5XdRRrPOdRGbI9e1LB8a4kT+s8c2Pb2RW2e0neI68rX6ZrdpK3IPysq7awzlYltmaBs
TBXqlS7zDmD4ULRzNBNXhSm/lhET6mz8A5GDxC1AxrCYkKZiX+/nw3/Ia2M7n747ayZLxpnoB4cB
7dVAyVvPzzWiBbemtjqVLCSXmlX1HG6KfW+6YQGDW0fX384xgcf2todxhgOauFW4lQJeJ6/9uTXO
lOQXiFNboPmmXFPkWd/MgTQpJ6VM+Mgn8vwcwAawwaX8sgZZqDth0l/laHOQOgpn1wl6Np57DCc4
+qUYXEnF2R1HHmRVP49tBIP3uciEEE+Nmy126nX2+ezRbEmp9n6Tbo5wpzoHJ9NIyJqPnhYnSnsw
qmJNPVOUZcYbwvdNFzK39wCbIIj2a6v4XxtnG2Ga51sTV5nAD1TQ4PC38HYHrQtUi2ifP2J42qep
0nTeKZZO4DHIthYa9pMpoMgkMcOGloJSRJCXIf8HuJJnPK16BEyM3s+ujJqZlVI2bRItN/4cprf2
hCAS/3S02Qux2dPqlSbAT46ffomV3J3O2z8mcIBdbIDw4eU1Pl9C74pz5naEWQRj+jeDQiB0EC/Z
4XWW7mwFKXxPDziN2p/zBktqNtDrPeUO7ihrX2P3atvu/d4SuR1F7mg3DUuRIikiyrjnR4BRXjPp
EQra47ylT2Td9OQd09ruzGTRgpjEatNRIDl6DoVquPr1AM6lLmufusC2DZ358gt4IEThx7d1c4au
JKtr8iq1snMisOtg+pgKvZAr9A9ysM3EcecXCXIThfES73gTpC8UO5PsERQA8653X3CvGm/VFSJN
R2s/VU1LK2l7mwMWo+BU4JZa/tP0ESCoPl+ECw0QpZjewR8c5JFWdmGHKJnvmWXJZTCSdRtGm46q
kUAlyvJ/XrfvGzAmUekyxGerlitBBBT4ZPa/nYA3svSEgJnfP/s2COGGig5O/2OT55lcz3YopUB2
3aEydUF4E+KZrtaKTAPrdIptEcUEtZqWG3/xbtswSAWM4qqUTZf1CYBZRYKW8J2yHMl/EvSjLsmm
jC6qAufPLBPNRcGqRg7F+mQ57VAGxl5IBsd36bkURSo02Jc8t+wHiheU2PPinISVG9qESsdR3qAM
gPXZwF52yIjVNe6rti5OU7rciT9io/XhV2YWRF0ilviPTAbdU8LBzTWapZ4HLeSkYp0pNr7y0G1c
tfiayIABt4msu+aVgdqKGxSNUArNzv6aS7ZSTCpBlblDBuVViK2MqSxHg7tT8S6MLWBBPZnNEX9S
2G9ojFiskrg3oArucG2o46Zq0C6LgviiovF/y8WZV2msrJzpl2RybYDe5Y4HGcOuCyIodpsbJJTo
5qaRt9345QswpTDgUr/t/xzeX2iXZnUiENXzYJJCRE277Awoff9WiWSO/L/H+4dn/4LYObV2o9eV
j850sDx3d8Kgz+s+JyeunCD6fZQJgNIuXY/bdxFIHTC5tYLRSQ0eRiw0n/gygN1fS/yTctN+ZV59
9rT/OOQOze7CBtmdQdaSGFdtWlsV9l44d6ue380KPApzY04swaWq4iEsWnVJ0jARFQwmmd1f4Ab1
0SjZ2rxGApq+pngZOaITs7thYocY6wLL9TQ5Exjnac0CnB7msPqIwH2jjP7o5K7QP8HLsfK2QXNQ
9vGIS6r8aWgic8AAXiN4VjcLpV8wkJP8LdGjlR8nryXPrae5/qfzufQ7pBJ/hsqW5kN2YlRpaVpe
XvW3+PWtYsMTQBVeNP4fvZ9C0GZrHpa8CbtqqGBJZhIyIzb6HMnhoJcHr7XUh1Uubg4kfK46TeHD
esXF+vkGqr9LU0JF86Uvx78DmcnduuZYvfPJQZeT/Uy78eiICP+G9EYErqrtVLjBULc9OMr5iONo
cbmFiG7bJ70JYSlwb/U0sWxIN/0yObxaGktPC1Aj+2MbF/3eB13sR07T3iWAR7NbHlzVWkgsgU3Y
wjumgar/NjfZNFqp9ssKAowN+iwFnhViYLg54t2EzEZ1kQdLzhVye9z99LgvKKErDQPPfFQnmwSt
vdv4ev9SyGsX0aXKyVau5lGa/nbEsXhGvcYEgH8Bl+4gULkwthIQ78ShBqJSxxqgCHMmmnmTRwVv
ou0lHR9M4re0dr2WZ4cBeJ9TPHk+ccpDR1FeasVDywNUlTZp2w4NhpuD6QNTe/ROpHl1SOTH7PxC
JmFfy6sptNzLXVqr1nrHUJwVIBqJFWgQ2Zdgehw6f73YPi+Agz8c/nq9nrJTnXXxjuciPnq+dJ75
N6KhzeG/Pho/4lIR/E8aDw582po1o2WFalkGK46SZeyTIho6l6BfC8yyqTuin2W0+F8wj9GGRKok
cwPpMGuZXMoIfljJLWiS2mtNb9Z6eZfr3LVqOVSoHeRhY0wTSgOFT4PDytElftckzFGwOb7MDbJh
wgzPf6BT95JYCm1SVzxxfZXb41LQ6456ZLGiOr2g0PxGGYJ6Y0ryT6y3mmjiI7PCYqYRsZUf9LUN
WsgRFuzhdY8b8ccO9a1VTtIqoURRVUwqv5Xy3ZUjkfq0fVsORu0AxnNiWWWsQmqx9iSheJ4+L/yi
D3hiJ6Uh60k25scV+awGOctZZXVR7QoYc7vXDTJ1/imXoomMJ+zVnyC8gGyU+7eP319QJEPM6uYF
B23SbUH5odOFyK8E/b69d0Lu9FFvsxGN8pWrDEp/lo8NcbYT+fRDqmgHoaj04gs/psIdE1c6tyUk
IQWsgWN+dFMCFwo6c+Die5vFUdGeqIyT2WiGblUomvbpOc4cVApKBbfHWqeGAPQBTszTDKTBbWeG
47APcitrnlcTwUU02JPofs8MR4R74bd2iwideU1TAXcW//WZSjUxU8d61u3Pegu5Wp2lC/KNsqb4
JqMRoPxvx5jFjDgP0r1ZRmMlm5Lfhxa9JqcJ040A7rjnxjw3wG7ObQmdx6rohjBYlEyM4h6sAs8I
IGoo72vpFo6EiVc6UOqyFpTwSs6PmcO3kgKXGWs3LWxAeNBrQZ9N05yK1iQgDEvDdkrqqylGEDRh
nguURxiJzbIRK59y8ryP0242B3CgKlW3x6bfXMi8AxHNw60IiLXSVkHwJVBsiOT9kZvXJfX5/2/1
SjBfeOPTrt3BElGCtCvge8Z1oz7vTtKtapCYTPF8C/OHYMRXQR09Bk79SRVer42nNX7VsIBe83yi
0Y7PHTd9HwGpx40mrouDaszW5eXthvbCR8xUXo5MCvBVmJPFAsYwZHa5DYdBt9bvu2/Sc8mquJy4
umqUYtuB9c/pxU8h+KknjLlv1luzLaINyxEfTo5v1nKBv3MGdYv653xHvSB+zxrUGTk6KcUBGKPT
vz2hI2pZIyEDtXx2CRuABTVWq0UZQcQZWiKzp+34y8Av5KCKqVprzNlIIrZ0SSj/X9QIPKc5Bzxd
2FgnxMy9cbL0GniMNmN5ikPXjsgdxaN+/97AOoHdTHVizFmMG/aiQqqEM0aZlaosCVPy3qnEOGc6
SCjtoi94tU22r5PVBwziVDq6EiIEva+kLQlW7ZoUwcH6tG2M16zyMd4wHrhXvAsmRahgprTJGNhj
ScWtZkDZhAMldAKOQK6CmdG0lJICv/Vc/s+wgW6cu1AqwPtUGt5wWHfAhLSlBj853m3ilQxirF0w
NCcUaQT1xWB33i+yzLzmBw/T5hAUhtYhZzrqsksAkXEkqRc8WHQYksbqiv1dQALqj4Y4pFq5rLId
k3jYpkIOpyDeNCAa9PDSzyppRfSoxKJW120VyAIQVB9r3joVVMR5JGEh3NcGJZN7udlvBMhzSYm6
IHUo8Ttd6MNtOE3FSUG9uMZcQmXvU7fhnw9e3K8n9x2G40NqO4mhIO500fvKYTPVLzddd9X+zxFt
qd1TRu98Gq0Nj3qr22hT0bhansLNfBMoVPPfkBSaSNo9pzNW3Luu3tU/xg6fvjKMh8Nlxo1Ho42d
9cptCYNbFfoV+28+WnrK5OV/IPducY1Aqu/vtLF3XfSJ6Ikpu8qTDlW4OQTQVvehILgr7WNTOSsN
JsJfXOZXBqiAcgaOnyx6+eusXEbPdhLL7J4pqFoRv8IfHhZR7hQPfOmcWToq3wHZ1Wz7TSpIfVpU
J1/aGP8krKUBTtn6byURbv8epdB5aEG4Ua0CiU3YyVnyFjyH46+71ZmbeAWWkxM9gv1ZK58QVGKa
XzGOj2yGQJlO8vQayyMZSagHFgkaS7zW1SeYQRL+YvKV6u2I3esII45F+YgSzcea6CzIejVdhCHX
Nfw9xWSN3+tNeSV9ZHX3dBtyZcr7eCuf7NtQiM/xb3Qv1ZeBC41Buam9SMuI8xjHj2ZspQ+xNxp5
mZkpgC3IQE87l0KjOmPXn3VfX/A8slUwFN222LvEuh8RTkSesT5olMONa7ERakJhXTeiORkfffIc
asJY7KnwhN4e0chRaexGeh+nRaBl4g0DciumikzRuoEQsdTlu7iurZsK/X8B4GFTmpaFE3fdMYPl
a+/ySdQ7Vble/hh/+tw/iCYVzTM+57BEF/90v7VW5XdjDp6rne0ohzfTKNCCtXoNpRcPB5ZQs8KZ
hDb0lRea8MVGXO14if3iSdQKvqHKnvYLhe85ntgJGC5UWYH0lcN2yBGWoqukPwSx7wh4Y5mEPrAo
pHLlp00oM5PS3uDLY9EM4WWSzRQ6tZDQjkKba+dpSYrh/Y688jBHZGdr0ttiQMB+Sb62hNf29gNz
aZITYBXTc5EJsGWpMyrMNMK9GQFNsbtvaNHet4VRC513p9cU6klO7aJnSoHrUMIFNP0grl3S9AFO
vRha4iVD9n98mI4KMVoNWUb/E624H1/PTspISzM/VIxQnCb5tZ4GmYlAf6IqMfiQzc7ZsZqwOJ3O
8GlJsmFBDSec2NaNlOjDW25Jd3c=
`pragma protect end_protected
