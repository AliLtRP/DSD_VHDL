// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:37:18 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
f3GbVF8OM48KU85Wsw1IJ3daVMJcANj+nzOTC1BQoCJgHsfGmylTnDjpxCBKgjeq
4Ds1OCVBEVA4XSrV+4NoXQRZuSS+OckjOg91hKPCDjXrsvqnKDrhfimQhg6wuJFf
MRxqk3LhW252NrJEopB1fBfZQCL5KuvEwN/KMyiSAA0=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 3424)
ehBESw9hB4UHSftvXdQZiMal+Ck5rh6hBmq8pk7Z8DQI6PhiSU58LilKgPP8dUrh
uAHaBx5gyBPbb3r7SGaGT/vnV1NcAIftHpEMK5LPdd/o3ipIUlRusmKQ9sTtp0sM
DpOCcPepJm9mdd9IwusTSfQ6dd7EPMU2+pc/sl6PUzTBpgD9iklKU5wB2UPjBKsT
ZJGK0jZmEsJNqpVD2PX1BAqMkf+MXNQxgmvuipRdNDW6iQ26x+zctKpYl0CGUcCp
NS7nh7TlrJKqEee4cJkTxxBnRT559g2MJDx1y2BbUbROOCu0SWsjszcitb1IeUM9
etN9wFieLDInO/OmMdnId0FPEHCptOFoiY7n06sMmsk76gP3XBdr/Ly8Bp9DpUB2
BVknUNNf3sJtW6v8pqxkp/ZvfLkdO8msOj7Tk7YmkXy1j5rdm2yrISD6gfiJDyb4
f9JJkoBrZDbUVbi++ytm4KTVye0ma+FepVI6o/1haRYVPMmBU9k3uKcelcXL/HWX
HQcXfBZtzKVeMEWjmiN79PNXCX/DzDAOyZPZ0IXbytGHVmwTy7QU3SLmqJAEtrj6
lLCG++AnaPPV/wzKKcZm3MY1CA0nlhMw2nQL969eSudKCmX48xjx+uafXfW8rLsv
pWZ++S8pp1KngsLY1cHtiMD8gM9Kbuh/VBrh1CvusbrhRoekxh9LyMmjysQj7Ifn
Wz1YYZ7PVpAtDqcPoME6P2DosdFcE2kueAIDXmCSkwN6ORZf1uaCQ/fZmcqHefbs
z8uspgmz05aQVe18ELD3jV2bMv9juufBGfk2I1Xzqm7DuFfgh1s6pvcHzAyQzzoV
RqSkvG7rLnAYMGA/JBHGxhhzNaBRZ0ollZEIDSAbFJDiiIeDWSy0TxO+vfJbtvXJ
oiv+zd/RsaUUYWzWvX1dlVkyx8Npc79dzs8JxVh5+9P2ANQf7pB2eZJCsz5tHoH9
ePtfUyJiFPJMl+eHvjQB11K2FXo9rJWl8Ctc4EZziGrYfOZp1ytFU/w17CZba3vo
XPAW3SQFRCohy0lozr/cYPjYMH4OmhOyvvWvd/29Kwc97cPf4wha/JNbqJuDOiC6
8W8vZjEOeqRMBQ2ypH7VU9J23H24hdhY307mxcau5h+ekhMBxAwyfs0L7MzeWFle
jsVwh8Cf17zv+eexlS9BmljcqTUk4zUOe+Y2RzPqMoJXFmgWmPj+e8TDKavCRPr3
+hbJFmd4QE9obDEfC7nuWTWKTcW1vFZJ4DttLzH/oficpuB9Tx6KILQb+i0IJ1ZG
EIy3jqT0akSCEtv91igdGctCJbigcIm5mWpSD4ug1YlrQni92bIrq1xJqTdpIrj5
SP5lJByu0fnYlO2hdH2VZY7i+Vl/SdkYeNwa76xdtpQ+YlIDkqqtCNJLKeryCoY3
j1Il8N91Cchj9ncN3fKm9JKVd3Z5gC1ig8V2zyqdoRnWFepQxnHk3BA6wi8og4za
lUEDqjIyg/f6idkPofGgCq1Tj3Icr7b2qxjPbtgn0mml3VFFb8bnaPFBTcPbCwZ6
0WNlqfHOXvsmGkJIkibtVScRY0d29EXOZw2xgkU6brSYMYS52zkWXuG1h+QYzkhd
1WXveuPGXjq+mibTKYQk4lkoQL+oA6xvrQW6TSmYXvJA9GsoeJCoUOB4vYyvZnRT
/pp+XpnDtDfW0R43+KTxcLzQAyGo3vXd7PZ9of80KRp9XMeS0ot0apEtlBfd42UY
dU5tgy48NmO9/qfnAbgt06YBxB9GQa9d/tUJQDyJegc8XeGD/AGQiRJ2/6s3E8MG
3u9TSwa3rfsxRH+MIvGMNb7ha0mhqDaaiZneBnm/wLbsJKwsg4HxrzZ+QitchfCs
KPS7gwUflkA12ryfmIX9lnPRmDbt+JO2W8FykqGLmtSOtmmAMDixynVwR2k2YUkZ
pncFgMcPgfWy7ZxDjitDg9PoPSlitjUrhP+f46o8ktapPbDbx24taMWBC8qT1Xjt
22h7eOg/rNxlVajaVYmpo1wC3o0S8pLB2T5viMR/2b8uFFuTegDBr0x3D/MgMWCL
1MMc+9cN9ZVZ15XjKPtakxtoD0JWNJ0lFnfZ1LZ1TcQhdLOZPSYA50wfsAhvjIPg
fTvTxd7SrCoZAxkull0qVC7dT7vcOhd2wiLOy83OQR3KXtyIBiguMBHM16K90bAa
VhwzOfG1TSVN80FnIisdwGYydrlsFAbp/Tmb+Lvg5tzn0ZK0V2je3AA0y8slkaqs
97oXhDdBIma/EmM7zFMfD5WQF2fFMpR+c684aM4iAz3l7ZbcZdL+TX19u5f0R5KD
Xby+3kLLMrnNzehrA7UqsH+6iu46H+eVio4QhryQTerZyx/NZB4vgLMhtk5yUbYy
iLDn9eLTFgxl0zaIgzszz0R7IW6lgFftVAvGZq7ByRNa/ncXYoWThiqRqLPE1srU
0rxIcaJBqqFcA+uTK4rXujaTMMdP2sQrWzszRMlLmDjhRj7527dEoXp0vLBQI/or
abK6/nrvdA6YBRpJW43L59UFxdt9UvTg/Gmuj7+SXBi8wCgNlb+NTpQE0rZwuAy8
RoIMhLU9xOhOV1r5UO6TpblJoEOsKeV/HJo8NzPGbd0WUeHIhgkHWmxQM0ZNGU0t
4t90t6MUA2ovFpTIk2fIxNpb4aRHjbqWcry1eTVcS7WnBXgGKNQeYa2lI2rtGvge
QpPPT4D1IvHmiLqRAB9zps1HEKGdrZRPU2l3Rja9kfECYsOng3Vc9ssL7GWQsz4u
00awj0Ziu3fkHN5l0JZSiTD+LapmXUr1u8ZXXM9mXNk9MTmK6AdCwJyxeFUzXO2k
C1uCJwO/NyvrbZvjyZdnUzqy61K5RtDGzxYoZecLBntYRFBylA4SfuUI+AFRYKCr
5QX2VatAADYUtb4TDhZfkV1a/FNgOhShRhAARNomrhZOn98j3t1LFCQXbZnMV+oy
NRMCL6LeJdUvc1EE5Klq6QBN/3/EgTd3fhh0t/gMbPEieTwyMiTyQVXxhXCctxgm
m8YqksBCYM8k+tBg7u/Owo83OdnjlAx3BFwqC/MdkVQTOIHiSSTJUr0mmDSNeEk/
NxNabz27iz/VjpT+zagXEzFIQowOf16HVD3YwzOlFS8YOWqU23NSbfotiboCxWSB
bT7dTn1TmS2kb1wxBG+ODAzV2yfKe9Gj80mEdBclQEWyeFyJ+IafHxYFJN9dlS1v
EKXkU2WtBisN63EhjpsCXFGh9HZ7eZtnR9G4nh9AESwhQgxndCrLoUKWzDwAx9ym
RhBcuVzUYqDHOnJSKk93N24EwbVQVkbRtuz7ryLvyoXePIwmup9GX4vXBgUPwG8Y
Ly4H00jzbqQhJ4kADhuVU5J5TLclUnCQ/APsohx7j2DFGi/t4OO4E48uJBXeOiwa
oz59KX/NnsEmsHEsir0oSjfEOjyyFKR/LUxzDq1Wyk2cTTYEmd7oid/yJRZgkdNd
N28tVhpMIo1duwcLTquhpOSCSbiF3/JkNI5YE/zGpXm23SI8jeGEkVfOJO6wM17a
vywKXEAqfb4Oz1LQNKQHyVhd72yvEYzVtRC8WRr1NDyp6hakeK6sRg3ytN2ZnRWc
Gf/tOpBLX1Y+X82AUgFniOfW/5kGWHIRXR+hX3o338Rosx3ENvC8r2VhRvONkvsX
cO9wf47twg72MyXPaLGS+cUUdyIv51WASV4ZFyfYR6s+orHTDZXc/xHuA1AlBvy5
MLI1gtfDduAtJb4zhv9S5Sq/tKhS9m0Q0qkG7rMrzWWlLi/4+MunbZ9YJ2vWU+E2
07xw7P+scfzIrFr70myvFIgKqM3eBXnuAAivZXKOywvcw4dZ8P6jtz8/k73++NmS
++9LC5sc8ha/lcYpyzzSlJ+Md4Dg4/R4/z43jHtsAl2GN4ZxEoqxwPbezEe7Qv4d
O1z8IqjVZUukPrzoZpAmWF3kWWceB1+6Ul082/tRHo/BSRfrBBhDxxmA8mNVRUUI
uzsBRQBN6sD+gYHa8WFHZmUyFYrfufLAd2VTYY0skp2kNoIzzaivQ5jkTqT97x7u
DOHkyTz8gTphJGyc+wRLYXw5r0KSNyTvoOOr6JGDmwTOcVoD/7pUuxy2yjQNzn/8
plqWLuNyR8goJj6acj26MQeeDYrWb0M2sfZ7tbzluHEJbWSx5QujwQcjtyyt5xKB
JArxOYLfEEryOtCMDZaGGKfvZex6jbaQ66GMkrnKWTmS0g1hNtIviqv+U8q5o3Cy
ojEGHn1RE971PpnMtJOjVLkYERRyplBQuQLPrEhxdg0fCY1BjUysDmiFSJFKZVbo
oHZRSYaUJmBn+KnneAJ7H/JeNhrjO4tOH8PrrxoT3LjC1kHm/swGiVX0cn8J99VQ
olJk+3v6U+xl6DBN+pkcWiMSdei3Dl/mW7EF/F97Yb4KnT2DrvzV+6bix9db3enC
oQJA7rIptxpJHPZjY4Uu1bVEBwx9atb3YfV9PVztZneMC5L18z6vMx8IEbSpB1dZ
p+pebI+Ncg6dY4UIZecmjoEWABu4JGKrF1HO3bGdxUlcAbTFdcpQgIdYLrsbuCbL
oLKfHVG2ETxFc4KK1raIow==
`pragma protect end_protected
