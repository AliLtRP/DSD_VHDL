// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:35:31 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
d5ZBOUkRdZCNMevh7gCNHA3zep19yjld+jfTeARyFZlyhDhNyrJ9kEMYolxqnzOi
pWqdYy5yu6iYZE5vZiHEkh4oXU2WnNFuibiTMdSn/OmL/KJiNHDOzalNQdPQKKkJ
MLXKz4iPgoNbDPV94rhU5koEhcV6hzy11Mj9SFH/Nqk=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 7152)
0o59Z5UnsP5cfk1w4RIdmUKWETfdRACXZP287L6XoRzBpql9Fr0Fgy5exMWPF8XY
AZ51GIWTdLecGi/wwaJxV+Bb21dylq5XTnxGh7rmOJNS+dUQBDWbijtPquk+1VME
1+Z2KRp0FyXwjZIJKBKfclOPAF99wGK8iPEvopFz96U+l2HuKMm7OMlOnNmwM7YD
Q3LrTE69Q+tZNMJmrCqR1iNs8AGIiINoBH2LWTNrZ/pP4TuY/iqs7csWOSbDhwuZ
FnpiLdf69XEF2g5KZ0ZeSK8GFbzp3YR7Of/fs90wkQ+nH9LSqCA2tKuPOgnZSPwU
bYc2Br6GrSReytBmdPUdg4XDbq+sCtpblLfpXqBhIYEoCxgRQmxSzG2YaRSWXd+s
X8wKKsm1nXcmRhbmj3mcTZoXFgkcXjbASU/yZN7+rWBY9/CL0uYK08blQmUkkgHB
7SkE+pinXPGzwD2GUTpJEFB4VuQKSeLw9jThGtrw4AzCmoh+d8aQTvxZcj7lQl0y
KpZMYyKoZbCzYp7qZTFHhNPkUL9AsjtDXigCSAijGaNglG8xVWkauWqQJBLu1fH2
ZXWyGN5PaWVxPvKrRnLc5Jw/uecOfkiZ0z8syh9neG2i4iFRPUQsseOhF93pv5sl
iJj+6e1MI34ou+JLlsiwJjBtsY4Jm29E4wVYUq5Fh/CceE3jI5pda7p5AytgYZor
HykdDKy2wLpzIfLFGrG6Djt4y/8Z5HdYEvyE0BZQFJJRoqyrlkiTv9joytdFd1Oq
2UoW50B1YC5DO3Fia0Dcex1lGE2vuBjiVnqFfplkAZX5WTPS98jQYxAvX51dq4PI
54y5vbot/GmiQ2CPwR5+37CA426rZlr/M8y8lkQy+xrNiWSJ+A59B+ohZXeF521M
TNnsNcmXM/7K/fFjyQjNvDNEtNp/yzJnxiML14Y6mVEDowlMpbjzw1ZTRTh6Oeh2
Y2x/yHmgSV8kCYExikf2FtXyclMrsNAPjGdLec62W1Z7jCTLZvk8qLuNLmW3IqAD
E7NpWZ0fnEr3RBLB7DKS/zGKA1y28g80JiJK9KXsCk26Xk1cEKsVJtpXQwqlXzuM
jlFaIq0oIuhTSZoqxBUzeXqqC/eOz4IUzHvbn+zgI1uSBOVYbZ4cnavn9DxDuAyF
dGNg+zDwAItvfIClQAX6Maa5+AB10RXmOyul3tcTpezBeclIJhsgapyOk8uwfwuX
tzCFnRv6MCXoUMEGK01+B7+3y0WIMQ28PpZswl2K8B0UyFhQbYm5F56i0xCqFNIe
8usP2e0I1CPjn48XouUF2lyunmyv5WLJtYeY5SBy7U5zZlFtx+LEui10zPi2IO7G
KFV6QqBX4c9+Onj2fmv5EFJ8UU+F4IFHxd5K5gq6vpykV7o7YVAK0HvnPgH9nM2Z
juEw2ZnT9lSRpEWR3imDlB4GHYMXGrOLaN7jB/udwF9baoFBnIMQ/aT9IcEMwVHS
+c9HjCexACYTn8omJOd6UvUVLno3pKQnaheB472kG1bGp0EpeKx/E7zzXV13A9DX
VwqOD8MaY+eKgHURu5FWgH8iFFLnFVUzFYFJdSQRys3JYk1aBrEYlLi6nkRVN+cj
xfmu0JH4Icb//MoSMNEewneIZuUF+seLfAobhG3NZvRcJnbMRQ5c38InPCxLkQou
6JHVcgFqOv1dGf2A5sD5iDbFJo9bJgPAXr80rOjpxyd8Tz+blT3r2q5q4VedWVkC
evbiai68zve4aCHqIGPguCdekUfyc+ftkxnVhiWs/sR9RFabTVLN7aM79/Gv4eo5
JQVOOOKFcC9PV2jV4DGDOv1Y6+sIAWEreuVGpBOWNy87h8mzkWoRDsZiNj+DoxWG
yFdSZqBHWC6LYlvUgaetDAssHSUejAte0bmpwXckr6LyRbQEdm7Je1+GC5B3pu+d
mP02+Apcjhmgdb/ze8BpCQRW7ZJQu1N9MWjy0l1h5Q1QYGflAuEO4RxPJ65pnEDB
eUKZ0uAk23pPub7jZwH+XMP4O4TkWV3BZVuaa7Fey1P/80ujTWMV0MNHwsEjWsDI
RS9zWyRLwqY1KORiG0zx1HGSnt1/sDhhIzNs8RdfpjX4vz9Az+KJfe5RqVxR91s6
RSu2Y31y7JG1oEmwHYmY7hX5erhqtnamYeFxc4dQaadiGkqVjHx+Oq0JtZ84y4pB
XhBJrB6s6B684AeFiXApfJz+KN8GFymIQOPeEd6IW3dcg2ycTuQH0GmD8wGlaz7S
SIerW1FWwTE5vq2vIPpklo2rnqw36pRvnSIx4GoTRU0iEf4eWhJpZTTVby+p5FX/
0JQruxqoNY0cW/zCOD0uW8ymG5Pv3izgSAsyC7Jxka5wSM2Kh2bsQpcxHwx9Riur
mqNaFwLGwofGsesneLMngwso1UuluJiP2R5xOpsy3YzXztG4LKdIIW7J50kVUj4O
+OUO/qL7hdk0z7MBvbvJ5gxJCFY8YocygW5GxLfEGrTCkl8ALCpYEsuaqdOHscg2
bX47CG5cHYWk3PLgHxOy4LVHBmyrjrE37Mv8wvsRl5+BgSVxAIJU4oouTheyCWER
3ffpSpAUx1fT9f1GxMktFg0eG3SmHRymx87+ubqp1PvMFkznHQWgqX4AvKggHma7
aR8vWJbSQerKanX2hobb+hXC7K7Z8TKclx/9W1k94Zf7XllEY3mtgdI7x5hxjIyo
2AyXlqCrWxxJCtZDK8qdp8a7gJb0U9okgqjj6bUZLWgYJmi6iCUyMTB0Jm2tg70O
oE0NnpbnqMiGKvQ/ecjje3cIHLrseoF5mAZXNT3evol88cScsQ4u/vI5qOunDJHh
tDSlKnZzs+yfW9anPb+mppHpxdYLlPbCujIDDKuutVkXRhmz1IzVpqgH7fN01fKU
+maH7Y3JOLjuyIieQ/aljGSjHkf4Z8PwyrrPnVyeEoUpkM7vJnjwNa4Wu0oiI7Qg
KRkz8IvE5GXORQWdSTd2PdoLySzX2yNsITXrFEnIWMz/7hAJk/XMfRKNwG4m+DEp
bLQw9ljodobTJw5/TjT5zpXe6J5o+Nz8+L0hUDedZcKtJ7NrvodomUdq7sEVYHOY
tbtgpanIYILU5wnaaRuh5DBDZFZF8ZfVw7YEme+tX+FOnDxNDklsZ5SGvF8zoFN7
b85WPy4cPLj6cMYVWlXyZahfiqmFsFgZZrcM2kUVh2Xo5MSqta/O5P/hJY7Qu2RH
iXAtpvb+18IUEWw1mDnUOWe1kU4hdEtlgFCXeaj2aIf67Wy+UoH8uT5oKFH9yuOn
L8Tn+q0CGA7XtlnCeBCaNcs4rMuMzRk+E4FS31zcdY5oAtLKIJlXDyyC9hlwNNX8
k/BGE7dcCGdlW/OzD6o4gGxnlu0TbaZEcowzSerib8PlSWA0QuyabuZ+YD+9nkMd
587NI0GFpc0WbBR6v0oJpCwjBUMtSjZPQDA3rTy9ESXvdBvtQMaMHj+kuiLztbTV
TuzJb1vE7BI7VKVgycpLiRqbVx2Fbe2jBk62VoVo81PeJP3ZvzTCBFo5Ef/XaNql
0y3KMWw4wVTbAwpXIfKLO4ii7IMabJNGhg+dxSPh2IFEfhR4OjbSjfOWRL46HdFk
nWp/BDwOAt1cDwaFLZr8h5Z8nh47vuxnJr8HSgA0nteHF74Nm3SOdXov7nF0fgKW
PapHH1rf889F41WqvvR1uwBAvtzmhd4rhp2xqqU5CwLL4VTQzbmExThlRA4M9Acc
Ti9Tuk0xp8JU4OFkMbYoh0oy76+GykhBaJIH2CRuvtcNnMNv8bGahkYJ4hw0tavt
y9jzkqqkW2KAKST41Nk0CzF3mT2OQRJ/m+zf7dO/FPoo/4WxwMTAbhTKqOejC8eW
Iw9ffI6U/so90BtEJyuK2gnMeWzVV8ciBIZEDBzm2q+pto1LY9aHU6yawT/Tz2Ta
Niw+qGfIeQMscPSrLMCY+tJzAZPIbJJ9nShyKm4Z1W+e3h/UVzhis3/ljKjpJ3c0
4+BZ7xA6LiNmDHnAl7BQx6hyxx+WkreyO38Hjwt9f45TESG9ceXeaLQEx04HHqIZ
QipiPDFA3eB1i1ukWpXp+NC2pK6WF7QufZR47ODMmgZRN9fICdJv6RwRQDYB/6zq
8YqDWe466mS80ZLVxlxmI4g9ns9SVtm1bO9SkxVgHwWbgl2QsOAi62rQ4g3QwdJV
18MvuP1h3GZMdFp0+Dk+z+djLutTwop1/QZhLnbXuFYicij4mG4kRZcPqJbtEJTB
R0Kwt76+/qzadgQjyADXSj1P7yyaSpvKxMx80UG82vGIcLOw49z4/tkJ94FByUmh
C1U53Y3HPGHQGPVP2n948BuUAN8FSs5Q0Bg0OFOdnIcwJ3wITH90avazuPXkDeFU
notBIUePNxPTZd6Dmg8ojQtiQjzI9uh85JpW+O4YP6D1GIAEQ8meoyc96TIyGVcW
tLsbbDkLjVY1xPboYRD4ihe8B7XmsxcpzGNy+CKHRYMkvDhOTsFC3ZkRcMjDK5Pa
B5oMcsV3xIxaj9yY2VXZMF9QZAS1V9Jl0Aq/Sao0d+Yts6swdNFq2vESHhL862Ca
d6ksDcnUx6JKo49BHtLiWaJPwSvN2sTWGcIOhjOhzhWZazjKsgGWAcBLCRbSFLWF
Srjt0D8RFSwVuMOExjpFgJ//y/pwqkteKs8hM7Z5/JmxLnV2leHW69n0dC2Guyoz
1Jx1MyuhbHkKx7tm0h4wWUHq3rknwKD2lLSgERrxfCVwQY2rt4gJlSkHEST7QxRv
/orq5k3Bvjgzy9G3wspl6pbTPjQlgs2rNcPTHRcoqIHjqnqRWpSbc52F6bJkIeoO
377tL1lP79fLM6v/JsmGiIfUXr1Snecs+SUGHUMzmYNdvuqQbixX0zSnEGUUCwz4
btHDZj9JwDHGdhyUkz+pFpP8RobnZt/TkcxG/WNiy0qSq4e1osVqZ7xXkKvxzHY5
P+02eH8m4StkzDl2hUBms6YCe06MhGY08ic7p+mg5gQy4pFb9qxMGDQ4PKKKOdjd
7mCpo3DZQiMkdeaEJTFjatmwVLfn62GmMQY1GKD3fhQ+x1/arQVfCXsADvTLPTtW
awJ/GOk2sINL5Wc3qFE2vMDUQt+lU33vx9+sWzRTVSJVfcM0aWhdraU9K9DYjY8o
Xbu/lU1hBt5SEYG2BBA33Uib2gtMNuxTZo0L0nsGennbWutvEH6jMkO5lvofafL7
v2acyN4vogLGdnDQpnuFNLz6L/EWOcb37zVWhNkDfJbDatnkQME7mOerhUTjFwD3
BkRFEvNbr6bN5pQKONCL/kp+DqHbG9hwSw4BLf1gGboXY4iB+72EkWKA1ENqSurb
4aFrmLI1h+1tipi1S5GqOcbA0xEpAMkqfFIWbqaHMN5SteG+sDGbveuYIFudtI8P
TrLDq3uP9fTAhxYoe72+P+M5wpcPKd45OCYyTRzOHjBwX+oJ/+irWWoJw1AMUC/2
ckIKLxszXB3GFkjtMokbxxx1LguLAXCJ7XezvjWCpvuPKWwjKqJZ0YJtOCpg5EJs
+JNanDV9BjioACT/uDKfqKw7/rjwt/A7P6lcIiTk+Hk2UYlPtaehyS6xbaO2Ca8F
pVh/ZbSc2NeMivyebczBwTHf3EBFA7yAnjnLpZGLgXgwCab1UlHkxHuslTKD7GHi
jZy/Nq6BCuaHrcPpUxCysCAGbhvJppotsJjvn29QYSSQbKX9lEsWRFzYlkF66YXy
5FZwnFnWvobVbTPNqPKDWWilfIzclYUPvN8hXASuGC3dSVru4dBK+lNMSap6XEWy
5Q/zyMhFKZfDxVA9C7EUM8JgXr3UahY8b1HCN4jMNadbXy+3OUouYi/JuULS78I9
J4LzwGUkkPuGvFBknV79PyUJoKEZNWmYW1LTdDgV9LnTe08/m5yq9AcxgviPves7
EVz161y1lWGH2+aoKe/k7HBr56R4gZgsiq1F5e8VXkOiFMbh0ZR6IXSslGzfs6ib
QYVwrza7WQn7nxhKgJvsMkuDr3SqGNW+qeIi4dNV5oyvb/U2AgjbWNXmwESmeOkh
nCHMViQfr1cMgpCwBNDCyPgntDxQajJuioZ7c8Cr+lemuv+0q7i7o4icdfjbnKiK
3WeTwO3F7TsEG2S9NJ6AxYhdvMviUwwwhmu1hNAT3XDejFrcSEHQNjM1b8pohUnG
YZVkuqBzcBV3NJja95qyLZiuQZn1HbsySIp/v8duvbLQ5FkNyaqgTEfPWNwc+mDQ
13e9aHhQDLAD2M+f0yBxR+2sJ/Zko2GIxgV4Mmar6DN6gOI7SMn2oD5IOGCZFUSK
xUVyn3oYTFTIDofzFMU2D5eEL40Ms1I0GsU0SAQ6Xhnm2oFdmuD8Ttqq7ODkZOuQ
z6wcls9+3y+UpcW8DPu6gPcsn3VcOXjTkhqN7YY1HUg8fUo17l7Hx6p0iRnaET3m
zzdd4nM9D7r2kcgro+Q5MJFB7eFruWj0P376UmQxc7X5d95yeraaxlyxku8/AGid
Ipe+MpsLvWR63nbfwdSgth+EmgQpXc1z1KGt76uAJ/8Z84nr46rb8AtjbUUG0ytG
lpqvxMKj0bfn5wFVnja5nnDdNj5No/BwM/6YeMRF5WDH0MZcTmhhzfP9/o4kK3QN
DJON8+dY/XOaY83pUs1FQPzWhCr9VdIOxtT2yd52oAYI9PSmeaFg/GrLqNuGiFCw
cJCTRc2NHcjl88whbKTAt29W2tF5dhj+eAohumHT+de++Rskj1og2AXFV2Q9qTvk
ftbSSm4H9XxdiCkKRK28ZHINPFg9713kOEIB/pdyiZ+j4y8qpA2aBOIe7D3LiSa5
7IRKoDk4g+6n0+unuSWcpOMOqnu9mgG6zkroVZUfkEZcjGctLm8Tc5n7/H3rQIYG
IyZj/KevLSA1HFBu/HwYAhcRV9Pl1dA4S9uqyV6VFHrFnosobUwRfp2rb+kgzh0t
3faMmyEbciPTo7V7BeVc4XdZPIMJAMC1IA9jDfBC29dvWhKLEFA3I+KEdkfxvo8P
4F4WBiS2OWGMnWxGmk7Ksr++J9pFPtCROXwkRkN08Wxne+XaTBQXJMeBF7EWwQtu
2u8grfURvSu+nuj7YUVadZDsLTUYZ150v3kexAzxMJBUyZbSK0tl5o3FFLDJlOfa
AtsUKg3eB4JpIpre/IWgpjoOBvHZT73ExuVEB5eXkfKuPGZpr06g8ts3qSzgJicr
RREJphAslT2glsY+Rnto01GRFFO4cWL4JBO2sAgbt+N9quLxajzPiKGZZMebS7jt
7BCaABOtOZG36AGjcB8niU8Ls7Ck5XliUr+KUGJV82XTWE/nqEj3I6hCLe5DZqdc
Vrgm7MKTSx8qvzPvW+3e/NX2FmOjbUhgZMj3nw40w2YXTiZDQb9iDk7IEB6CIAaA
qIKl1L31RbNVEqR7UMEZlwW7ct3gxFfdbqkT/EUoVNTRZDhrzkOfAIbDWW4gAPJq
GzZ5ZEVKpIGKZPfnzyX7nYyeQlStOrdyIQaVQ44LPGG+Igcb070ZXXZ64B046jKk
SmYp6FKD5VkKIdFVy3xLwik2VL38wQk3v5YjcfmJaHsgvLocslAInXMNdP9ieAuV
ZXwGamIpAqjtqNQShYt8TpY/ItIL+D0/Y5mQ/k69JgwODg08Q0A0RbbFka91VPyC
bNV/eZPZ8YcA4QTRHST01A4W0lYiwUtl0oBZUUAA8v4575bnFaTVSzAASSwcUfg4
zhY5Yup/mN1cCDIuDiw3izrdkDxMNTaOcLqiLNNbcPbmiTgSkPpDGVSiGqntEdzS
Kr+ZDOdqEzECRFyTG3b0zQu1TZesdI1KcWMqjTZry/SX/JAysxvJR5TLF7l2qheL
SOSZZKe7H8xo84kjzeMHGueBZAmg9wGZKImAaHKQCy6IqTDrWR6GLyXjfg/A28T/
LCc/bKSywY36UJPW5cfZ7mL/C1e4qLrlQF70ijyRWFXMXStnsOW3yavaejZ3jHsi
/AmBA7Tnlvi3JlJJLOb4fe43ZTAx4Itkz1cGue26/Ski0oR8/iPOAT3rre3Cyqw7
k8mtco538OJD98v4NfsenRgM4EZOVjdNK9/Lkblu3bOicr9ebC2feoEbTBZwBfm4
e/LISu0FYcdOw4WE8fPpZTWhIrCQnoFx1KWjurcijjoB8avziwKt3hBinn07RtI+
T+hUrD0ykR5dZCixz5gM4T2QK5lf3N34IxwruCEJfkA7qDq0uFLit8VHNqkQahhc
5GjvQLU9111qYf4ZCO/t/C3UnwB95ryRkE0exu7FJIs4UuJsKHBO8fxlXbsCNBlj
YJvdSe/pFs+Nv5wrr6y7Zz1g0p2ln1dzCF3KqPMsT7xrcdvmhAhnzl75nw9Zhgq0
V1ZwMSdtmQJ5xyAlALk/9z6w6GPYfSVi7/vGvdKm6ofh9PApFGCKqFcVGUx/MguM
t3wFepAh2gwbGbUQnwMtXvlVfTfzxj5n3m3c/wjghpOiV8jPvqPfbdSDdNAtU/ku
ejJAJK0TNJAiyn5RLhYAhOB2p2/Y/BD+G7jXu1p4o0y6E4+i/qTPBfwwldBUEG25
3nm0ZXiFfQ1iRuAgD5BgvqlBxuoSgbnG6fZZSGjE4qvIdcLgfsVIgg8ToIsYcQrk
dQ2xXnlsBoBQNcgTFwxCBDIjxMxoBt0Hg9kXxQZFksskovSmWaB1qApdk2UItkux
GGNXjPmqs46ydaLMaK1KI4YPGZdeQXfxlQhj888E4BrhDJQiFRTXG8B1Hymjzw7Y
4jRZnHOBCSYT+1EyVZgR8X6Efg7yhkr9sMVWbHYqcTvkk2i5rDHwsSgwOMTnScOh
8UwUH26kuWdjeJy/Ml7k76MSlfo6dEdKjwKgOkoQLe7+INYHGfSMpxj6EmwqfH9L
l6OBqF5WDR82IZzmtN4vOr/PzpMW4cJSRySahWzz4BGKVmkf5NH+SS54TR9oC3ry
+2LIVpgYYm2AILPxnZL08O4MKku5KlpADD1X2WwzCEia9KsOaJzOiJzVI3x74fqN
/iO5dR0c8c/iMfOYbgBFVpwJabQIrcaceb97MDr87hgxYgIIl4ON2FNCNAjEnlU/
6fn8twrWGNuGNy2mvJUPIlAvO7XTDxcoMn2+DK+rPVm88+bXdGObk2gppguyGtT6
q4pgomwdbSP6THCr/ykUY6nueJCeIftYb1KCcQtwVgeJ3LvwEChL+SAOeYegDw6/
By1tuepne/erkk0NC5VJwOi5bHOfbnCYcpEepTyJaaWLWdHLQ+/J3VjHkHow20cT
uNlOnkkt8jDdsi+fwgdPaGze1MkZJa6S5NI7mRkQJSWTexZ8T7fjx4lUZQrLC0sn
GtQ2BS7hQWNYEwV9bGooqzq/zi9vsHZ0UUt3A5TBumCraVQkWj7oKHhOVn/+5ili
62A7bhA/KF5KikG+41i1Cg+vnaP7jzXflBCEMVkf0NfPS9ZA2UZdT5EU9gjC6c7B
zfj/yP7zHdKg0FVVsQ8t5hKs89/0RLN2MvIvk9vPgZMOWjkfIrHmmw4MgcchnNPn
vs3vm83ebhL9aq+Rx/T44et2RTHXEw3vk81idhaxkk3gEVXFrUboIjojB7c7FVTf
`pragma protect end_protected
