// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:48 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
bCGTYJAW0mUIOHaLe5mx/DDRQvajdRV0qpfWj+zwguhyol6OfKzs6ExsOrtTVn3D
pSaeaxNrQbt0Z1U3OcvvNwTW6qNbASkmmvcdWTD+IVOsVtyRaORlHMHO2THLHOdm
IWf4U3uORBDy0eI8UPhwr9pbU9fJSJjr3tL/ZK+HD/0=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 42592)
nxDgsC0oH5xmPMlfSwxa+qYrPUDt1dNHgAfUzMOhbG6RAVpucJUCXyIidvTuzwC1
QUVDwMRBvM9tAsbl+XxnrqhsXwDjVoKa8to7KN7Uwe6a0VaBNmT2J5WAF13K4kD8
Q85odkYqBDjkBOsVKQDEPAKN/aZDsBbtDNjv4G8Sg1kkDd0eZAN8C+bOjDUc42XO
fA4VzdZNXfd9WIfswemqEmM8XqtV85+nTmkaW7oiC/4ghu0IdO3pVQYs5rnYQ/Oy
tMCszXqNohDSiG0UzKifecjYsY6nVBhwJrZQebdTNVLmM/CdxKzqrxEeeyV4liNm
eoq5t+qadmxaHhWn0CkxMTnP+TDZMHBkSWHWadzrnBKaIU3xtx+Adku2qM3WNUXF
AMkk7xcknJl/GSEHaCZDEQk54UEeEWCofh2K/v9pw9BYuCuyTOgbssoVBObrYSzU
8+vJ3XwSOz52NjW2dkLeUiVhJ0etAXzfctgeC0A1+/Reu+rrold7chg84p1KtVVi
9c9B1qxKZGt1WygN9ZmxBE2uuWAtQUxm8BP8pDFmb7MC4FdJ75RuuyV0svDPEoxk
9CsQkIkSYXKg4Tck2PWZQTM/H8QbfY1lsHJCcfo0xkmn8ul/hhXMat2+g/bm9PlB
0S4IGkZCTgaTelqgqjCLhgHuw8NKPgmH3DVMaTty7gntD/QKPuQm3rmahhWngu7S
SLP/pAhFvURSWhl5fMy2AI+NEJr1iFf7KhaggSvo/8tccR/3qV7/E6yL4IGV16jB
yqPy7o5VLZPEwVZRiRaDdPedmcDyONnE6cOWm4vI3S4XKDnZTOgG5WJKT/lZ75Cg
F3gD25MJpVL5fVQmzR0HlNcdeR40NcuXve5tOtTVOoeWhhj2svLPWaLlJOOLskzu
q2iPelMwpjCHh5JFUhT3d73u5/hZp3UpJHdR0Qm6KMS6VWRTboa3YGWp3M2g7a65
sG2LXGT1NbihKh5dpUZE+Tq0u4CraxpiPWa/HYTTJU/dIqsJ7SS0ITtusuLWS6GX
Io/cePq4wfEo39JzeaWojixGgOj5gD3yJkGWJ5LislsuDqCxltUo/5HxkJJPKyn2
TXSaPUH005Vh7MqKRs4hNaPO4rQyvcuVhmUO/scVEXGKedR9/2+5hsZMwdYoF5oK
qrVQEECGQfrBkqKXFhkVEIVQvah9n/OYTDKfWqnuFoZGNrXEgySDseJPApT72FBm
A7vfJ746aD3ez6zBpsV8w773G/sU/6+EnDRkiLQw+fOV11TwkGlvGkPbTnFpLPEp
VJwo62ZfTmsUVBwxtm3tC8Qe5iPRABYINSKRvoDqGzK9FIP4BesxIRITviZXUItf
HrXv1Ae2IEm9lVQw3kM1RDyy2la/WN9RuEt9FriIl38SNov7Z0/mDu0HTxXsIXLK
/kqf+rPhJt1bBHshrhosCVihrCo3eWXFIfjJaTKcMRD3f2YA/GS+uDz+H+sYlHsy
339z6KrSiU/1lNXQeNivwFlFxEoFfvppc5Wz5WzuPdJ1S/g5rYvBbSQxzm43PKyH
TrVEpLS9C0Js4qR+8Z8ADW7eWeyEyMwlQYqCC54e+K8avJ0R+vHr4LSDIvRSQXi9
bo34IzS33eGTs3xVVHleKyEBWj8tJFgSVoQEiPv7IbSdTDRD4a0+NBMQ3nhaVoC0
LuhfnDk8NBs7bFofPm8S+oxBbpTLVfXvyyUd6JzGKWIrjym7uzMWVdFLvzAkbo7e
wKf1Ca++LKVOLKww/jIV/93BMOXFFpu3qmQgkCZeStb2WNhN4vED//QYTUAbofAx
EGgJk6LOXsaNRn4E10Z0X3yR46/gX3dQOhhe926UCPSqHH40J9HYXAPA63rsOAc9
vdrStXsFCaZyN1YuCKWmWtfol5PcJI+8WBJsHfb1KUlMPRI9vMkfCOEENXIpqwf0
s9o0185iCOnPCju1mGJVagZF9R1W5ZOGSGubKrLCYOPQ5kS2Z92pFCn4z+1VuTjY
Lqz5Z0HNyKOTRJfRZXBh91bjHQy9oiZnhggrmOJtzFseUGQHpuzOUWiI3eo7Cxp+
9SAFCJGOZai63Xi+iKD16YMnbsdVpaWDjpypH3qEj8GmhwSmjwuik497na/Iq0GV
1XADAha6vM3u+2W1jcvOw0dpCx+dy0N2OMa+wjxrDHLwy2D4unRSPWv5z4xbPKG2
A9RrgvACAAMPwCJw1MPfhGGhlmv9o9kWtHfBuPjXAlBWDQ2V8VIOlOLuIGMZjO73
KkofJsvKXVz+d+77vDtskvj/dawO1B7CZJCKNF4a+K5G6LmX/po5tJdS+gc2rGcs
0O+QvUExlOsHRWSjdwya0r/cmOuV0nwhjdSuKxxPZmPxsvviV33qvPKh5ygbkKdE
n4BOKVAk7xExRPjdb0g11uCmEctc/lUGh8iKPqzV4T5Ev0k6mJTSe7UkZAgdauTW
3RvENW9VPCXbefE0hkySE99WE48ZqDJDpHc4/CqQb/ldz2FNgKw8ZD9M3zeKhW3k
l6REkEQqgwNR3baWShM5iBk/SzZ9FEt3dm1jXKCyAkkVRtM7hSxHlp/T1E/Wmwf5
1M8WQ/qCZLJgC8kmwOprU7gn1AgGreyAHWbPCqMnIGcbuSLzs5HUiP38IqTVXP2k
96iDYWwDKXW0JwPKFkiBnciMgeCvNvFBA8Xf9Twa3YczXTruV6JuH1EE5fDJymTM
fDRJNFEqhzdPSqLk7RBhvnYo2+Bf0D0fltCng74HdOqcrz0AyPruiKJWgk94dGv/
fWvRMlfXdHEIEhh0tFCzRiBb+8Vhb/ul6wI5IcAJ+nmj2qFCgiZy5JKKudsG3gOl
kTUdx8rmKlqgNct4aaRluchZZHDgbAtlnXd7ndCSxevnAMrcX3o2cDgghB4hH5FK
5NDJ2bjeQLmsSPokJXCoHX2RwINGKL2jZs/Oom3fTzDesElie6MimaEKDwMmH7o/
4sTnCBIH4oi2PHLNhKoyTVd2iul3NZ/JJGPn5G4r446vyayh12LmRwJnI1eBvXUy
gzP6492JoqBGI1N9o2jzdem9CTjPcIH3K76t1J2t4XR26clMwN+HBpk3Gaez60HD
7qVvAvfUu51yvxz/CmCwAenFMzv/Xd8M8470c03de3BVEz+b8NtGITh8V9YocFIq
Ais98RjEqGk8nxElPnfklH3T06NtfilZL83f3UbWI8Jq7wn7Td8ZZ9ltgsz4b/E+
uiJGY3a6LLsdAviUwlU2RpjPALP5pYPvg7Hugfcx3A5eWjwqWoQzdFJXxHumH/qa
6EhNTkyg8qZbrjEK5KmbcLQMAv31Dlg92mp8zERcW4y2Ssk1rFc1ZjpJsZYSKr6c
7GOUp/5XeXeEAnS1xONhxThJozdfKI2QqbnK9QGF9isxXQufnlDgEIPSszfG9Fky
5JIEgdtRSfJ9v0QnhrOQ6U4caPSJk6oKlqLYaacZeUA8U5mwY1/nqy3iQU4SXXmU
R9wMGY3dg352aCTr2kfkT9akfplEmePtujnnbwiHWtMUMMtbXJfrLL2q9HLTKq1q
fGshPmuRRdIXslqILK2TZ+Ohf3Na3+6hvc0+Yyj/dsxJ/AWMdFWLfRX0npyj9QS+
2M+nIgFDQZ530UFvzER/8eSuk6pTguBvf3PJezCXRQVy2/KteKvMkbeBtefA0mj3
3I86fNbsetG/l/ZpFXOKIfs4BNO9em6+o2iUEpteTUzNoJz5ybpkLGS/5FMnkA+7
wrB3MqgKmonrSVRiAN1uB3WOdIIVCEq8wFCOKawHIenPq0RrNCAR1ardFmhE+uKs
QUb7Fg2+YQSP6pmcT/CgMwq8ZO79P+ZRCPs7gTEuzU7A1Z3zM4Re2UUqTNKac+wo
KE2hPr7DGPk7I2GXPAUACEoQHSnEFE2kbPW/3HY+EeO78anPHGxcf2WZ/U9/RAjn
Wi11G6pT98lXxoTqaN3ifBZHppOtD4ka/jaaGPBizB3Ije79F1DlBoHxPR2K1hcF
ibM7HBCUGc1k58nCvZQ3JK/2AtPhB4dHHr8WldEAZCYgg+pLIJMErz0DtO1TNYfj
ISqOWv+8JyxCj1iIvlXK9Q5dq4wANqDUsBxC0No1AxuC7VDHLoh8xeGABQvM5qpx
uXKdTVgbbiGCyE3Oxx9tJ/n+HoGpuzucPUEo2VkRUTwDGying185wOlCGsLdf715
R0a2aD6D9iQoLeMo00wkYr9as9CkcZZ3uMGfjudPrHUqNYhF5a883CrT1+WOlvJf
JHq/rjTI7hHJgEQUKNkkJnxJiewiVahX4w1/6111IeQHlY+dI9AXkm2kMB4GC7wt
6yj3TE1qlY/mzgPsMQ62bcqhDLjxwPaQiS+oc9RYvLLW5TexpGjiEBSZ5x7ctLvu
nfzQ0wO9eMQdgcRl8p29MsNOiPhmTiNK2zAn9hY1V06+lioWYi/XbRJHihpAy+4W
1rPQAla242cXkkZlNVPrFy3fM6ru+69nqoXZNrZE6K2YpTcQnX9LZawuMlSZrhLI
YfttzpeKyBpSV600XCpkPkfWZ5wUxCsJHmG8pHaOSYdLShpYLM5eGXTKfx+pgEpH
N91JBB7HEDSEuGynTZvWBVMfeeG/0mX4tMyY+aBG97/BrLhptth0lU+8Eb0hbWFn
1d8QUSir9EPACkRKTFlmfl4wpyQzoS/Z/synNyPvmnO2AxyqDdqjCyPcxBFxRjyh
a4g/C89c71QDC6Lym/jkki2MytStJ2EejQ8QxWNkIF456BKm/4r0dB2wtpc/nWJa
KAkU98vbiRrHH2ytGtEs+lYYJ30u0VsZDht11WvLG6A0A0+RxvYuTT81L3c4C1WA
eOaB/MBN7kUj4m3CBHhkwxqOyoWRR58QRPU9iamrQ1iuONMj+Ll3ZnF0zQfSIVR2
ydgIt8+Yskcmm4w3UNCJk/WiaVRrue9jG/njkMHntuEQOMf5axacph7VFt9oRxLf
OCQeownJFWAkL/NxE0KUKRyzdSmnEq8lcRfVSBpwxA9THW59gLvusiUVMOAA1ID3
u/e2/q6BLkmcllNqcM0FYX6Y/SyN2F5eAkHpSsFnsaHoTgqocxDFWeiKuLUyF/R6
6BhltVWbTZ/S3kviJ6SXHtHUTbZXjRH6JgGzhES3YZbsyBv0X6K82b/KJ3XsA6/I
riUtF9T6Iw4rJvvmtmemDxzppFL0OEPZr1ZrsdTT6hRLWhaZq/ZEl0rzzU10Mvbf
zhkB62818pwB0tQzYQqSUat72afPeM7mc4y/9JNYxz/SBQaidRxXrv/uvzZkPlY1
HGl+/VGe71l4+s+xws22h6c02soa1QcFCNffqGjizaZXqqvU3pTOZcOzNfho8p/A
HVX66c36sCxNrwnvYEfn+n8YtISEoVO7JTlQBzmS+N6QiggQSjWxJkY0P/oZRuMb
XSlDPotgcQUpddJir0j25TGFXOT/qjXydoIWvb/ap5OL0ihBqgNpCCTH4bGwncxb
QCYmjjqJXgZE1WNX4bpTI7fenw/3Wt5EaFHeTNZcF1EOzCVpjXkdygiNqTdA+19U
hOmPDRPNYNxLa8NReULhhc/l5yYJePwSc5YM5OUyMMz4UQrrgIQ8mn53NNsHknm7
8giv6ce0QVpy042yVCHMmkmCmX+JhC4y6+/+bC4ueHgbGiDU27GOkCIuqhcpHOVq
8qSIBXEHoO6SgSYbDrWG8q2EjFmO/6opTRfVn3O474PFj+c3m9cR/l2V9SJhKRxx
bZcgHxRQ7jx4UgoWPVpowjfyJyljRsrQMY7P/HqKK1T/v58AL5ExVe8yK0JcUkhE
dmUjMA3FnF0fhkgIIRgpN1izXKAOg1RIYj1oNd56GQ7Lv6q94VlcJJaUB0IAC/JQ
qN82SHDW6SmZqvyYhbqa/gcAGQPcko11kUsf96/EN3AOMIuzZ/DzfDzTtbcJCdsr
TEqEp2Nng+1U6XwR358YO+/wHW/agQHy8I3xENJqx9SEBE+5bsY1wzn+w4wgN8Rf
sAoqi6LerLGpMa6voaPds+xHzgwXWADG0e2zaZ8fBbsHeiUtgIlkWleBdxAbXaav
bRA8Td9JBN0gy7pVgWTrFB/P17suPBGl+bZ68Wq8utgVaARVz+l4Z2QJM2nyHUL9
/G2tT3XBu1fziwrpVyZ9tN9bwqx2me/pJ/4CL/s7Y2bHESZtaBc5qtLJoR6DOxW3
eST2fFvnYy5sP3NFrpQ00XK9ymE8GmZlY8CYGrMrQZyKYfeLtkwelFyabxtCf9QN
oZUVn5tMpwyQef3HACITxjm251PD3U3V9jAGWIwUaiRV1MlAPsFf6Ae92ATJpCjX
ONFp0Rcbd+a1Qm2WZXzwIUyv9ClchknEXLzzyIOSxQmyKVLcSU8M6uDnbgiAF5Jz
4UdmI03zjsWpNXu3Oky9mp1H7z4Go3Pf5IGYTP2SbuojpXeQym/DokLj4L3lb60c
Mu8D5WzBBw6Zie95/rvFn1mam6n+zS9wbmeVf6WqPfcFwxx1xdH8svj4IvT03TP/
SALDg42PiYGMAyeaOtpH9lU+k5nQqHuv6jCrFfaoZlpdp9GNC573zx/jTFYWN998
UHwQZE1qQlbjjfmdIWJ7V7zLwTsI/Y3NTVtoCT56gIBA3Z9duBGgG2NDyR8ayEDJ
oU7aZ0yCPfg9kZh/NVP12Rj25hajXePhnCWiBeln8rNGruUu4KGfuDoL3UD87Lgt
vcJErgXGH1QDdAou/VLgZO+F1C0G5Hyviw35YBwDdLzR+iPOowQcN7XMqMvVvuCx
TQDCanJEu5I20QTDvjon6YQNRi1VPObUSPF8K06Aq0fAv3vOg/cW2k2VkfpjpV9r
AP8WAgTitCzzs1yurlr0CBrDFG9RKHkPeVVu28QYyawgrB36ndUKR0yb+6tVH6U6
HLoJmyr/68+7xw0wnw3Yperguqb9iYTKBHRfpVaCSY6C5D6jRT7RlhGbFwSMIilC
iAvQKCp8xvrvlMllYC7e8O2vAe1qiL/ePQTHmU1/LpJqc1VlbrQYpMmswECoeHmE
ac+Sz9hpkaYn6KA92rWPWlDzdaTScoGV/WviE/ZTABefoCeQMc6kgwzPOj0wNqsV
NCwzQKnwPaAB8+GjGnKdSHP/TelxQXwAKyxD7NNWvuF8BDfk6teSolSXJ6+0Wj8I
GlktfWJf5WmqxpENxSxUBiqJ/Qa2+8GoyK9hUjBlILxm8gomp0ntsdo2mu7I5ep9
Af6V24cQGhuvCK+Akeh+87Js2iwKAf6EQpQWf8r3/lCVL8Wo/vJdvXbXPMtCtD63
RMeaX9XoWGU7wmCY1QJQY3i8htEb7bBXhAmMdR5/H6XOY577FMmDitDEp/eXzFeI
HdvD7Iux49B7Esd2RCMwLcS5FPZGD86IlI3fxASOJ2eWrrm3gluKgE87PelJ8b7D
S25/l5Xj25ZqTFe3t3fQKRLAkTyOq6QAF0aicICboszevQEkkImZfe8duu7F9YUE
GRJLvPksddXwchVMH9P45x6mrNALhcMX+IRo9yWF/leTRyasBWa1uwg1NilbZ4da
CJbl7EJihFX6pxhJP/4hGcu88az1V1+mC9XJiWR8HwOjsk/6sCBIl3+TeYXCzfZT
y04SyfBIw3XpnYdjM3QXj9GnjnpTeQK78JcHwm/Oj2obCRfrQQdMTRFERz9FHhJ7
ZuhYKUPGsDh4ZkwNto5vLmWtxnXLStCp17Za9nMsyVVKxataVJDg7vCPnD/5kKn7
ckOIla+O3dy+Z+0Fs0pTB4mE5p+CW4IxURQ6hzgvQS6mfoOe7Yxt/eM1SueSD6XS
k5iPsGvhxX0uq7PHjwYRLLV8jL4HpUQoyMh/H8EEvewNL+U/Og25OL0Y6CcNJWnP
Fi7/PUqISLHwWKaQqv5P8ipMIwllSr+yuX+OH05WBTl8+svjAyPB8BBM2uPdW2TV
PRrWF/Qg0NcRfpDxiB0fyAZYMkESjedUuPTpbTanqFBHfUXgniBboXNJmsneGy8P
/06dmfNhkvkT3Mkfl+UQ1Hp7LZDeTVT+VoNZ1VIpd+BiDU081QRPx91LfqeEe+rm
9o/kV29lKSfxxEMOYiJ45ayHb/8iE7A+fhq1TEjZFsyKLnH3dFcQAFF0nSFqkZhw
iSiku8xF7yxCzLnmiPHf3skXS5dJzAL2qFi71s6GFycr4AbwH6hBwJrOyrHZHt3K
7q4yH8zf9kyM8F6klR/O62Ja8MoXksrEtuib3q8ouUPIpdXjQ2AJdjtGUhFgX5+T
e0Kiv5+1XaoBZ2qtFD/l8LMLCSFyOwZ9gaD1U9Ng2DQj59u47CE0mbng+wQUbdSR
phaa8iT6ypoa1PBnHfWnLZYzaItMmxIv1i9RYrN1Pgw7M+reXEpnFZK/TMZrcjpc
F7yNWyr1cJANrr0yPSKYSZnBF5iK/0GXH9D/vqocfKrBehmJZGygM+v2+waZ42UW
E5QT7JFs/ksdWfMBXkPbxtzL51pMJ5RMZaDC9sIoDmhbFrgUi8Vfb8koit3gKoHz
csTttsf+TtjVqHcFzIshN//rLAlfQucKS6MjWkzOPBxC5TdVpN8fV8gem/DIMnYy
aDQYgDtlFfx47EKbCzbNctjwnqylvCu9/chA1S3Xx9KxTcf/ANo6Wud8fQxwZ0xs
+K/rF4MpEcGziqAZaT1u30Yg0zlJdLXWAnaFq4oHDnMt8AhE1EZlLcGhjNMU33mt
5fqaFGw7TPIjgKUSltidHaInmCLSWhbk2i6MypO8Q+KLy2EPB9uVCEap0YbbHT5M
KZP4NAg1Qyt0LOoLckTaBeYP3OKWGlFySPyms0aLEtUoLW4KttXKRnplE3x8UqKE
Z+PJc5klEjmZRhjW0WgYEJgjIjNUUMBxINfC4bBwwPSruT/2PONjjw4Y1rAERB5d
6OsODJzzILh1aC8JVhGVHGfz1WZBJd6THJbvn9I9AhM9pPjrBUYiacGMO3ZpzLmU
tNOT+5w+8HxEjnC2Mor8cr4IpPUUWHCsYUM3qyhr96b/D6qmdPhq+Hog4hEVu84b
AvWckhNxaW2o5q0ZI9Ahf2bzGqTfVZS2HMeq2JyXYfFm5V+VslaZ2YgEds2bd8bk
CvJHku7GMbF/xb8D4+jFF39S3qDTkkYPkC3QqauvrLGRsJr5u8XM/yLgIhgqbvVY
OTCAv2vXheugQFkZuOKfP0ACQkV/9TuKSeIH40bcQG7DC+KenKZxn7j0EOEe2bQb
djMiy53D5Orbs9WZowHYMUF0AbfsnX4nnURZHI9qRUxNxVJXOcn0v0B2RiI3Cajl
w2zhWcwKWhbRjwSmNPx8BcLZhZkt3U6ocxbPKftRW5FjwSO5vBHjrcVUjphnWXFT
gx39qzzAJOonOx7FHfYGDSTyVGzRJ03fAA7ifCrodOrapCRP8xCWfN2YElOTSN9D
ZAEUvkontufgYMvlSjxj4tf1Py0LHSkdZjSsiZXk71lzdMTKkRQSxDkDUg7GCehg
K+ZB+jXEpDzSAO9bxgQgS9jGKKv2r6BbDUvcVtI7eoIDx5F4xWGsaEnMrhdhjjfX
5ZlzUQ79pDiqNYO4rvtj14AToOMdA361ym6OPllsYQzMdQS0BALzf9ZeBDGTg253
hVtxMR7TFddbw9BGuJ6s9disXTgwspmDB1uBPr9tkf6dxMz1iWo9LFXMkvfFPhQg
JoettTRJVa06ezhboK/wrLvoOvuVhjEuTLoYr0ehFMaSceP0GDn8HeRa8vlFPvgx
yLKxr5nqvEX3J/GkPCkjo3XPa6b4aLw1e7JIyqEEYP5UI0iFZsTspVuXXvCc68iW
+VySWzP9GVcY5S0Y8CLJx8FMoMn9FgTOO+JotuH/fh/SankUCjc62B+DJv9nVWFY
IlRz2h3tuyJmGjocxiLnilj+FsQSv+uZzlcKQxO1ByHkuLZ4A88S1ZVrhiH3SJE2
N/xbPqUuAadaJjrTndNaGwaO2NKLaY8OsleBaZ/c4tRV+Nq8HAiqKaUO/Z7MIQCi
8FhjejA/aJuFSbOWTxeHntfqG4oDC/BHx8aGOS4ozP220aG+YJtucbqnKWY+TR+N
yV9P8ie8lVkvI0RkIiL4/khKAI+gtF+DVx8fcx+3jgKfzW//VPndtV1/+i9uiy+m
w5Z9u3BghUojb+pW5OSEkXVmrwdC7A1gcG8jHg1L68/hb0gn/1YZ2b+i4PS57dh1
ahEZwaIP0wOR5XgNZ05iFGWHb7EWs/nzLUE9daWF5t/Vqsh7xkrKOXC0rzPOmEM3
BqvKBG8NEM+JrbUC5iJ7B23TVa2DjP4xuOH7L4qctraHN1wR1rlS4bAbLxdhhm94
iZ4zfkD0EAyFvNjj7i38hNNgtUEEq49XpK4ausp5u3hoODIR8LZTJgfElWdcneJS
MuLTVG+s9/ptgPRq3YRwmOkmR4h/bazzkFHx3LpAyegFZ+6z3Ec1KI4oIWV8Qrxk
cp+ubI4bSPQWyW+2X40ztmEL23yQ9ddPcC7IVyvVGdQ/2P1AkRFF8u+SPZQo9QNG
bltfkqXeeJspbgQRXgyzkOiBTRG4xFsh5H3+3V70RK28Rp9V4DBeFCxUuQvkwym6
yMu7igq1MDiY6ObqnGlqvQO8KBFDo53GDtC8yrlqXvXLmK6e2odMPDSys2oZ44sS
3E8CJcKiPZuWz6/CSB6av1MtOOX8ST/ioz5jFFva0uGBGkcte6Wl0hZY44i8q1CK
PJ+tOS/NANU8rhqWQ6SgoCp1U7NY5rKv5tPhMzRfMsN5DuMgi2kco5N79Svvwdio
o3PPho5agH01YoMjvij67zZWeY+NmMoxU17ilEqSOhUrMUjsC4EvYW5VQFij1aIT
Tbnggg9pzQJwMcyr/cTdpgtS7HbToia+iCkRavn+8Y3lwLPn+FyOhR76E08yfrbT
YmCUGgG2rfCSop3j+DjyqJAqZCz8oiqv/4o7yPd90FzPyUeOgMkQwFJsfcADxrZ6
XrQmMeCwk78nQLa1iXecFktNjHE0r2EQ+35qRmXsMDn7WWhAQvFxoo1sy2c8eFtF
GaWtq06pO8UCHYwlWipQVusSCtkIs8QyoC+Dl1yUqwCiGCOaAqjyJZwaRLLNhVbu
QOtBP3Pbx7BhMu7v9Kmi1klIo5ofJVI04Ug4MxVP/pARWrCxkfIeOH7CDCKiy9+8
Vh9Zgp7eljtYydp7xU6USTfd/8g3/Rv6Lx2tArNxsKTNGf5trnH3StFF/WBVBRx7
KETB0h01Y8qDG/ks8euCNO4gaRBLmofhV6wfffPPLHlmAI1H0x7vhFyDP22Ljwo4
BkwIab6wMiUHa9ZkwRzpcjE5MvQ8jIcx2ZGsCj5B58qkl5QWib1XlAdqYgjtL5P3
C2e2R9aFKk4cBQPgZAooJ1sJoWkcqUeZY2cwBPAttFHBBb45JpgtQm9wB64EW1hB
ufjzYP526DfA0cAzq3cGDnktQzTMfpZfSSg+qAjKpF+uWCkiCj6bpFxEnildJb90
0cE7O2XXQSNYVIqPxpPvn6noTI4LyJBqJ9Xp72sLpTxd3GvejSc75MkyM1iG+v+Q
qNLsFeSBsE/HrgX1GjqVgTD+JUdLN3CdwNrS4Ssjb5oqE+7qpBEL3ptZ2KkNVa1B
UCK7J1JjfOkalyTAuBRl+5KX58xV0wwflfDqrB6FIKHmkk7ghnQX0K9a+4zJBnma
xmhq2DawukdMp9CnYxkH7txNcIr3P2WqKhr/7fXp/65MMAwTMqmV9jVb3P9FHBH+
pX1BOZB72s41sxWUSK11vg50+H3O6rfrRaB8EXTB/aCjWPuDf6VwRr0ihK70gIy4
UCVRmB7JrHsg54VQrQDbVX4W/JxTPZROi2OYgfcvFbiQzp6AMCqtdKURGVHUR8O6
OzUQbhwKcHl6IdmWiyWtlSV0fi4Leo3s4t6L6XxB7hSlzZ1aFIJLTyxsdf9a8/Mr
3noMNwww4x7Y15vQj/jXMi8vDYgKEf4G45g5truFg1wqdT6zw1W80LJCi8WZ4WDs
k40pYOgbZpX/Ef/Pxbmx5iWhVVLPijG8w+pU70JujR6F9okAbYzhrV6gD3NekaGA
/Q72r+gsyI9RMCfJKlREPi9urcuYHHvuhEWeTy+TNfU06r2CBSdA8qb1t1Rc9B6h
U+KrV2wPqP5jVEfSbwQRQVB2e/vbbgKzTazVJJW3HL0gHoNqLLxMXiQltUbzUrvz
yzUji4h9zUUckrKkisG1vIUZcm7irAaieqdPEZS8ve4KpHN+ocrxySlWd/Lkpn6T
TsAI5pDUA+DHwt1i/qWm2dakrdHwwRkotC3+E01j1g8yC4hH1sKxmXvv6tlVMHCT
U4EV61rCyfeV1TC/SxawouP75HM1TRaKCioGWW5oXcdsTSeKafJt7GZtGsheIO3X
qxJHuFdmA8QDJpprbT4WvsjGVgw9kCRBbNuc8lUVF6B5O5/sIy4p+O/+pu8pz/xm
xL7jWLJdRPePQ6nYH6fF45x1Xu+JHpqaIn4pXmmYqIEzx6W+gtXDxlSKEa+cVipz
CrYqg4Wj/qH4UezrZoV2S9fRls2yIwIhcsYaL2urVuN7GYy6Z51qMLC7zL6gwcgs
wNDC9fKwMjEPDykcBD4/eL8aDS5EezPJTo6MV8GfWf8njVUob9zWzBsWTaSPNc1t
Zr1SE/WsT4xtgJcbTehuSB4r8qXDqjs0Usq2ziaNpCnzfZHKPxXMdktW3FbpW3ph
CdE4LyyFNWyyYKnWxKDdcsJ36nPI8beEGWM/1wwGhrDnvrahYMAjD0znphw+bIqL
x74mbzUAzAiBtKKpNfoKIxNUVGmLRZ1ZKfLe8EY6HsH71AzlX6kK7t9aUhXXsnRL
tXwpach/10AuCgK6P/f6tb8aiKJRat0Bbyvl8Q7dNPPYA5toPYd7Nd9XYCeIfWkg
usAGUrLXJj6yKHqci4HcNbTtf4JMKBcYz8w+UYGM6Mw8oQg9gP4nV6g9g5jzyoIs
yAldD8aEk2xZeVYef3GXMZK3U7K0VVE61SDhvOSCsnaqkoIBfh+/PQ9CNq/cAX1A
YIG8ZffKWhYTynnEYwoD9ztSAW3AZax2l4iwTyHFJcKP5u7DDEJV/JS+EPuXKtaG
HVucKDlNsQTkebC3tkiBanI3I9tvb74va/QtgfUAQMtmdNfcgmSa6VyQlKIC5i/s
gqMOd7aH1vL1NLKL95VQItBCYs6U/pHyXUuWq6bjQQx7y+EFPy1Em4kOP2+O4VaW
w8fyOCYHBbn1cfM03HeZ6ZDHRa73EKUz0O1BQm2q/NtAuPvHIEaP3hOg4AUpPOfa
xz1VTARA0miSfRngwl0gEldeEFW50ZOlTNqK3UtkHaog0DzZiq/ETup2GP6dFyqt
12yu7uvgDGhCPkppMDq8BP+HaGssX1vWdLo3p2mLovmLr4oQVzimAE5HyYTT/Hcb
03+ZR5r4qUJ9f86RQwNsJGglfhOO448emZ3EqbIzMpkl2LYBU57Y7268PXKeyE+i
/YV2eEUaWawy+Tmpxt6kFS+3Eybd49EfcTFKAOpL7XDmRYRsCIJARb1PHdDpozze
eFq0wUrDNsNzQJpHavHkaYqJH1b0EE8/bjTPEjiXF6ViC7wSyn8w8w/oCBowtOoa
5ifvCSG0jTVqobgvpjs2q+U9be6F8jmChNUg0Dfn24+3Lx41tFidATkXwkWrc/HK
VGMqGfP/i/MjkI2YXJ6+2bs/AAnYFeiWEfngNWBBZrhUdHNUT5ZOYd0h5fLN5LGn
rjAB/morFATpGwbhwXtG2gL+U6xfsgsnpMUjcPjfMcJ7rHhpKsh6iozJpSyFekk4
AEUwbHcMDgl5y87BHB6l0lT4s4EPkaSdcuR54IVZA1dXfx98d15CdaUKXNdl3kF5
W0iZ0UTzNCstw+Qi4yMFhoQU43m3lAbYoRyMcDuaReHMC0iL/YN7OxI9nbRpReFL
mF5cbr2aJk/2tOPkONcTwWswk4TGTknuFSMIdZ/Es8Pj7Im5tEF37nniIXfYKC+z
4d72YMLkxiMjmq4YARwzt1Qm3taz/PGePqRylCirs/wykX5OPLu2ClQfAZHk6nap
awqIngiBjDGKE0mdp4mDndaJ5VUERJsHRLrvELiw24TtMUMytTUbSTXsxDYD1GsE
MLR+CH19Av6Ua/QH1DQWmn2zwv/AEaIKqOSwotjvrLi6ypWyCVu012pzpgrRj+Wk
xNWGTuWWNk4ymOwpxDZGlmXgkeAAN//oEOKfQFMrJDHGM4iohnUf/+n4ohogTLqC
kdFIH7kep7djVHMsLWZul1tnrd8DEd8aUOXPwKWUow05OUNggce7XUiXUWz99270
AUcDfjPKAX5/6XPs5a3BaMt9q/WUjnGbFhvHUi/bpjIlu0VST9xipgWhS0vvIVTf
yca6Dwi/ep1tvccA8Q21WSBPtPXR3Abpt9W7wJi7JK5QAJG+UBvqLTJY3K3XnFxI
/URVNfA7BrNx7MoX55mjiPlmZUEC1z623PlPcdAC5ONkLtdaf4s4e3n+oKt9BL4V
rMT+lXYZl5CNqGgOAcjhQs1cFeN2zbINYw6EK7uLL6qjGrnq99Hu5z38P3tfe5WJ
TM0DmJ/hX83LrYgCbGFi7i91uZrN63M4DmS51igMJLezXfFW7LQvegYaZ/ah0XGo
3raXSshoaOmDh5+nx4jL9gPgdQsdP9YWfBqfJrB9vQmrhaS918CiEXIvtFZwjVGC
FgA+G9VZnrWT9eut2VLj1PsAToq/szFZWjX5tL1wbtddBoJqdq86icpKTL8+QEpd
cyfGrWqsA3qwsz471gk65yqniQXLtaUjrPwbO76rAD3HMoP6+N0GbbFYAE+TFWKw
1O9DapUgCE6eayZG1sUc/sit5wa1RSN+jcVezkL2/QixtlerdjQ9DJrhJ//4qqfh
8z7HyE8z2shdy1WZBq588N3XoPf6mOybKfdeAcRlbvT2OuQ7VADczpCvNk+dtZHq
uJcJvmdshYOGU9xbqhkVAYGthUR/A/nwb96V2g3611Gbrv7TCA9l31KTCzg9cHlc
ajeCRPTZ8FP2YSHa4B+Dtrp9SJWzknHh2fJKw0kzrxn5OglHREiPOdTGugII94+5
xsS4po/T7yGFugu30bowppt6cp0aFUTUh8OTKnfRgS29vdMQbiSRTkFQEMeDmad2
wotBK0f1QcBNqEJL46EgMmOoYvhXDYHc7AgmQLxWVRXRYiBerCPSuNZC/wrmn4r7
I9IMigD7yLuzdpr7OIOLGf+XUq/Rcv9Hhq4zIUsxl1ykZXh8dUw+o3dfs8JFvAmY
4SjUKToyaqWfZV0C6j8VwhTcXZfaMT4hW7NrlAl2Ms4G4nr/8QBJb+RXp9fxQSej
bL52nnyje8Y+FDwCW9RnYKkzACYltP/VvHCdKbpdZaNfljLQXBhRs8dGeQaeEs0r
7KrzdL2n7f+RfRtqQQIckjIMdEF5uMtdu4uEulf+44dCQpbIyv/pWsWWoqTsrArc
Sjn3pd/4r6i9EJAOxcuiJz4c+neGQA1KyYskDmJ/IZFXzdUDz9Jr8WwYOmHvUj7E
tlC8B9lm/PX8wNRggItiEN0iXac4JCTAlTd+HwXo+0Rsb8RaZgjS2yANSQ+zApxI
nbDIooePUU3yBR5VKS3ylpG9qOskNH5hh60mGHvsqKw8kGsxAOrlgjnMWcbJT8AI
UK5Bj3N2Whrieu82ynrKmgQrt6zp9q/7I4S1Gq8tTE88vzNgP2vi5bxjm005LPZE
SQ/79Y5c3Zy4tYRO6I7RQ6tWGSEYFsk0AGAu3m1xmcC9vYvatk6fnSIMmz6eGHDp
dlxm/+UL2SDFKXEt+63ERufZL5gx0kb9S0M8tmW/s+QpK0ozewc6s5KsW5r2UlWE
k3gZasJtEnX2+1m93+e42ZlWVgwgGjqQ2acs2ZXLVpXOsDZEZNrncnsTzu43efBb
1YTc40CbmfM/bF5UNnYbJkKvkHeJItBVPf/RqRPXFl5hKDJ/elz4kYd+WhmOPXuo
83bnFqzWdAXJvKnUVK8AeQas+pqHvBduDR7EhkjH6sZxuKYCzv/FbKhZ5rf9OU3O
ALv5AT2CZEe0ExuqUseVCknCejBVCdAT4SEm0IM+48fO2mU91tO6gNdFTWe9ROVv
IQ6k0vXzB5Y7rcWZYZls6IQcPoCtkiRSN51fOh+SkHm45xatRP/mWA9u/u/tR39t
RshvCK1lIQNmPu8pUJieqkFchqdijEXppuvR8tzw2ZWaSXaStvM2HBOqx678hhI2
ePeirIs3GiD638XS8IpruaYfVUZJRAeMJgeLXB9pTFAEAE4wbNnffzZtea+moEHd
dmCw7QIKlDH8kmPQHQeJ+lWVlpyUkkfITl22TEA+hZoyUoru+8S1Lpo7++rIh/Vb
zyqBUVFKirmYP4woe2kp2y5aYuNuRA7xkmcWJXqQgt3rtTXE/8jglzDr/zDf/qRu
A0YBLMeN6TX/h8J0WmFkoCrQ0yA0yJ8B20dek+VHrgElrxTsZ9dhHFPTRIo5Q1fV
MkA2ZpXVcLRxGCmwebGv2y3a6JS0My0MtCb5Gb8QNbWYC4p+koOH5q0yLLVd+7Mq
IzChvDoyby/BKEzupRmWd8P03gjeKgc2i8Ub6QxlhKlpdsUIaSeMTWfdQu05dYj7
Y1uqlayC3rHPM3BksanXcAU82tofl2Her/RD4wkwHk3HaV4dajLC8HRzfrLuuXfz
NV0vATt0X6BDbz2GkkU3z7/Ovxn0UCKCadVOk8JWm7Fmci3V7oRI38TAJXNCFlj8
1rUsP252liArMsFsl+usYZe/eXaAk40d2SYS/XHxcWPGFF3+ewFkuqJiylMu1LjO
2EQ+f2oPhlGlTzQ45WwBi05lvtdEeBBg1U2tPIYXNP8VQ/rW359N3CfH28uKvWnO
hZyLU1RlJUAu6bflSziEtIcPxTxmdeuNJsOC6n3uK6+Tti+59LOQZhTpQKO8XJD4
2nTBjZtfPX06Fk4ND5Ml94ipvbSDFe6vVqfoAr6tYCggJMYFvVxa/UqyqX6lYjC2
k3bRj+UhijckIExpASjdsyVa8eFkd09jbeeA9BqA1u8d7/soNX5Uh2Sp/WYX+s/A
quQuEt+wIal4Ks1nMi3SrfUF9+0RwCQz7n1t1oV8/af0tSdJOyYf4Vq8ILPDKbGq
+1U2qBY3ET3ERJJTvJAAm31KAJ6l9NFn9OswEOREa4RH0fv8co4Mztgko63vgqcT
5xEfUzlUh8CN8UEgeSM4rvkgTLN2znLDlCfM/BpCtlvUxdQeykpkZD5PwyGvki/l
wzPF4xmheisUeHTAoc6m9+mir0azfxSDpNCi94jljQlvTnd7B3uJnQuzo+wQbze/
pHTnY5Pka8otR5WKhfQk26qkqA59cJ67KCfq8AZxYRlasVehORxbU6lZmZeEjdRQ
gqpKhOmtwKbPAqM1ik82UPPJmMmql/Z6hlfBVX7hhcMPaXks+/8KW9VtABHi723S
SZjbwlPkNN38KFkCfvjMQoGg33Cepw//GrbYCjpJIuLa5Nn92MOtyMLjQYJw38ui
iw9A/0BBQRLUeL/7TcPyb1YRW7GNQ9/aZOxSXL9jqoUP/9Z/wYNHe9ikMKudBX0D
wDc2f1Cxl9Z6zcborFltZYGWsw+ihEOh7Z3lGxY6JHKJeRZXQnmekEL3yrd20o+Q
KtgOBxLUkfQ2Bu0TA6Nlp2Bky4y7Ix4J8YLR0cBC/nHxzikp0CKJt5OL5csopA10
NGZGluP87b9BR5zg75aUrBLddmp0sZQ4CBTek116tnOL9eZvO/BfXVBGNyEZb7Zo
OphOV5ovE2xKW1iTRKAIZdRmLWLTi/jO7sagNkgMyXqrQrBZui7r9UEgCbWG0O0v
Dw6KmfED/Yc8T2tLeUUvR7ffz8EvPGrb+mhkO5XGBw1UCptzbEO09JHleiS59lKP
XQk2k3zRPNz1JOBvPsZLGQ2TU6ixCuqF2n0LpPwFvkNExZzNVqJAdCfyMs8AYOXP
tAloJSIyEsF/gLT5ahjFTBfVnXK1exk3RGq4NM2kgcvDzbSsibO+zG8yxTsCBuvb
1db0c7v6y2tE/vaJmZ/F9toWPLk32nMVj0cg3+8WBUis5ezb6q6voOsGrYQmgaWI
P9nT6K6HVVhYRLPCSx68E3aLuTep8aSJzjIHOzxXjhUbbp/KNqZIQ1pdggtEaxeh
3GTI82AwVJapZ6HyRIqq6ftEEout2GJ1u8YnSs0ASB9NfsrH4kHQhVEeBqLhGLFs
AEHR1sSIc0V7512WEO7TxJqfN1DVtqxnVwszc3aUDcXVZKOzBVRePiwFagwCe4JC
cbBC8oqSFlneq65LqgOPl2fJr/LmM/0GzdDvPiK9BeZe9X729q3WjCCFYDITioGw
7e67J7XoTkXdy6Ot08aTezyUv0XmUXuhSFzoUtVEDphbqXG932FrQsEzi7VoNooY
T1zJ+vv/lATIt2T15benBMZEWWwTchy+Te9UYlyQja74AuXNlwtkbV7fBlcneSJw
Hvvjz3/83HKCJ4dkE8ES+bYrSsRmVDGik28s2yvTVXTaS7spGymdZbqp6lc9hbVO
Xf7Pdqovl8TaKLs+oFAfsoGHIACw7Lw8uRgGb4hOm5PPEVCCuMsMpSXY1qbb/rHm
JsT05R9q1JxVviB8dAmndgMNgMhAn82itezs7NBgZ7hkoQkHoHSzEq80McoVxJl+
dnFWoxVaeZsodh2FfszEnIhUW725quRXsN/OuMvJIMPwvUlol0MmXoc/WQiLhsYr
6rme2i1rKXAuosMsWXIa+a+KByKYz5ZM+hpgE8JRJx3ukwuE/2BmzvbX1gUZCd2b
hlxFbu6D30/UwSGs2wbPx8VPq7sfMoX/Tf0QSBgJK4g12Oigts3Z067G0GlF18og
9nBW2TEvUtGoYP/s+RGa+srUz+kly5PmImQ37YBheMmnBIdFOVc+N85QQSy06Jmc
UX3/3He3tbczQjdjS9d2nMwk3gYbGadZVV2UtupXCj6LQ5I+0+sD2NXSG0+RcqMG
qFH5sdKjLlAGFiD0yABRK8glXP2xb1+Hvonsx3vP/vPQoZ8oUjsLyc/yrlbKymZl
mut3QD09Si5twv+NYK948eKfs5iWT/hnyBa+55x8ugI0gF3n1ElwiyC2sQ2ZBAvD
Q7mHzYNbP+wN5sHkNivLve9m8Sil+N20nqWFksNdhHUkfcG9zzv0zvYpyCDQtp24
pUPxmce6O0XFV+CbPT3+/NXwHtSF+djszB5mc74Ey1sVf7g+QmWttygDjGmwAMGi
LJTDq/8sd0zYskAYcTvcyH0lUAipXkG3io7BoiDuurBVnUxqkQ9t5EufRc1jzOwd
p0P4Waefm3ktNZGW/zXwAh9sT7vkHtHlUB3sJh8fiqMEcWe+vG5B2odzczOqYxdW
DxedBLaDjkwdUG5WkuYwDkHzUJyuwHv0iSoH+ZgqMIhr0e68JpGK2/L5vby36jEP
FUAx8LKNSN6vsOrt7GHK6CcOxEZutNiFQxuNH93EaxSSNYqU4zH2hG0xbMQzyeDO
2FrcVEIBwhDhGQ/qqKxl+rp/TCERtGeZP++foUqZwPLmz0m6dm3ipkDmLHe2D9HQ
RKY6ATFLOEgytTI25RHPLqlC/fP+NW4g2acOZD9z+U/73Yks7R1jhlFu9mNqx4+3
iKN9gN54XlPVizjLiLquZJkGmZP0UdGT9bHvbsYqSIYi1khifIDGdQ0kxLRPrtDE
Irza6mtO1i1mH7N79D/MQ9ZmmqENS1F0mfgtZrdlQQ4C68Sj3LOcNJrxr7Z7yAP2
zG+Xn8mB0vEPLbFxnYQmdUO4jHfSsf9GnOfYi6zJk0wMFbCLHT64Yg5MFonyoWan
AlZx/3ZgRItk+L0wPI3Th9SqB9H0jXJ2XUSPZdDnqdiKD+lbeDXzk+IC1uL3u2Pq
ur+jjzkUBFjxM3wT1/nLO1DoRUlg94ODG6SAYW9tcFDcbfh15TZPS1xAlKGnpOJ5
olhMpD2EJxDGCQ3S8X9yV3t0gN1JqhoZdGHy6HWJw+UYxB8YKNgimO9+1se+PCoq
6+hI25oee9JRcDp3+fiu1rjqZTn/aBiYaj3CcnifWjHplZEO7N/c7tdz+tl4PjKy
6mgYdEsTjQEOca0JZiVULjT637SvtSMoT5fhRf0jPcLdsOHuek9jWlU5VIrFwVR7
rMeLsh7RdYG6b1K0RdbZ1ozKveqzKiCiMmh6my6jnBtQhkryR/Z/wc38D2ZR2NoA
Q25bYJRWU4w+fwLkNCAM+iKsoGaDFJBkVzY/DIQEkang3LQ51RD5CCBfx/gmPZLi
AZniPLmBEXos6vqTGdhhPqOcnWu1EmAq9inLGdsUgK0YJktXFFO5cEqrpeOE02s/
N8Oow+TYtSepigF9pbLRbsMaEPQynFJz/tRP6TJE9KQ5k5BEVdPGcnKnOngemx5z
+9eK6dZUSMf4D1QqrtZt7vJQxLQRqpfGidQaDZxAu9KFsrOXrjP033RDMU6SyOiN
FuvqT80UyJFFWRSAh/KV0DUTjse8YGJ3HNF5JyzDTQYcmxyY8qM91FQ59vP9esyH
KwHyOcwtkDGMPDj4HEiXrVK177rEqZrPtKTCZ2/ovKNaRubSG4IAczocWOihBJ9J
OZRBi43fYeBRZWshTmIKBjbOiwxLlZgL+uyvLtQBJbDChG2c0Vs01RTs1GqpkpSl
LhC77v69pBlDt/uGe7Dncn8MDOagZtr/uK5OOLIwErbTsw2O+VSIXxCKt7BwuRCi
sXIOS8ERvqa4FXRbw5Q3r7zeqTRido/1cdmPztJVe6i4f8Q1q3FEXzWXaowa8Sbl
W4sLRtj+PDNy5PoxlOxK7RzrgbOpeW1tXVpaAh7/OfEsx8Kc+jzDN4Wb9IJrYkdp
HHs0FTqgH5gkRuHp695E5gYiYKvkEr38lD1r9J7l3VqHvrOhX/WcyYSp/Gg9HnR6
NDQruK8SJdjR7tMK1ooOKrpQomOyOaGajybYIh5AgS9hW4YheMDGmTUFAcMfE7gz
iBFxGj9sY2bC58Q5TEhbwhI9vGjwlnztcIWw8ZNsX2XxLeiH+UDarVdNK/JwHctu
ebYdedI5pFRFcyP0OAazXfDzGAbGCSyEXrM9Va+z4spLxhGwWWNRXXj/FquCsYby
by5nS8/d5q4IAByka/CV9W/7OebgDYDzcsiY09ApHqg04Pbxih+IfScreKAfd9yk
6Zk7tikQG3zq9Gb9OiTUa3KKs4Aq3e27/ylF0YWvbqfqR0RqQImgx/eXiyJ9gpY5
8p1OH0iKRBHQ8wJzoQVKgL916e3nOFnfcz/QC/ZIPzHG7Os9HTzVXgteyT1SSaMt
Yeu2AbjRIylW7Vdo2EBiKpSJXfySlmjU+QVS7US/B2meKGIsRtS2IsKap1ARwoRm
iceATG9fbUewGurA9uA0W4TmuShf/GjAiuNb9np0Q5oM6IgMyKt7N7mOF9v77HNV
FmGqelD71u9UM6v7Cqk5Foz1sq76bVpKctB5Hi9sE12AT4qBJZ2rZy2PNGsIaOf3
SnAlpRkMfeVsaYzYWIHZ16DOelqfSRnmpqGajSb7FVvdF2G1z1VP3HqTTciD1uX1
srKrlXtJy++R7rvYJk7iVqOdSiQD9Px5we6fzK+IzTOHBU7PUkKsmBd1fmq86Uxo
3NT62X0gweRY0pc/FFZ51lQYDIwetaxQqBZ/JdqwmSiiHOzP9Ic1zKmbDLQloXdf
bZIHVevVNMEC9xZLt66/IXkV1L+eaugGUrJxU+1f3M4bOPTEQcjtW26UnD12MIN0
DZGdccptI89n76UkjLBL3z6MpRx3blFF3p0Wut3bdY3CigO/wv6ctLv/fxrTpEJo
eExHw+zM0VWxqcaARXB/0kfAZPK0v8d3+AKQnEMepW1sPBFu8n6FD+kvmtMaQjNM
RY5OCdkD1x1zFnb+O5kDydeL8wmsNEkNoFiqDwhiXuRk9z+jKxr2fD6O//2N6Tr0
Qe1/IkNX2FySl9bDggwMJuQy/m6sfpTN8s2u3lsqGtqh92g7PRZF1YVvYxgF/VlG
Z5Lt8x4MOvikBuZ9J4P59JF7byw9YWnsngilNFzBQ6EzyzmmDfIzBi82a/6tooXA
Av+93n2q5d0fIXi3w//7D/4GxfYfbn2vn6RCsHuvIwlZfbRahIRYLsnkb6mbzTCh
XNjREq6/KFqvrfNGZinw1llyxNz526HHQZnT01M2e75/N2D2xjkhiug3o9pUd2XA
FquhN9Ej9jB+i7u8wp8RaEAVm647YT/npruPq6BDelCiCwaA0YQxGzU0d1oEOgUv
9cVRacIN7n9lvXtkUCC8WpFX3I0Izvot5CmTbOBQlhHVKKa0sSY6VKrTg2FodBNn
xtX+hTLmdgfOR8uxs28ApJYdO03VTB+l9iF+hUlQP1EF484FhaXy2+BthRRJB3jA
hsFlfj6WdrksDpuwGB88/K65qJo3v7nDXO9WQ+JWpNftH8Sl6HxSW7+ylxxDxyeE
/mMLxyvB1fhzwJ2VINotNJ0qkRSYLYXvRJKjSPf/iCJ9MGgUn3BZSq1gGEsW++Jv
W51uNbmbUpUYDYK+cHUFzLr1VFnUzmALqFMNG/bE0uMDpvYyEHUXYfxCbW8IGjJ3
58rRlhJGjmZk6Euiq/S3NEy1heur/3+QgDgCFboeySFKOZpudxx5QpB2XzHUFiLZ
RHT6/EWH2EtbfwfxEdomf6zZl2lEGp1Jlc+0aNOFS330j50hA/2JdnlczJGGAHPv
vhGzvLbCx2iXrVivfDOcN88fk0E1ApYSk0DmMW7V7FGQ7/gLXCKgVE/KftTvOkBX
9NUvT2Sa+DBTmP/gnT285XHtad8VgdzHHMfb2GqZysUnElBG4EZ9rTrjoOiHaA1W
aIS2hLwE9ydZePN4ynX5bDKxK1vIvrIS7onN69L7Nmn4XmRAQhiYEFDlo+LGVBS8
xuaaHVLGobjr0viuTVhED1y5lq7eh47X+GVinLl2Olu5KO9Ds+DVuTvGJaCl7RdQ
uFXQzWcFG27kIXkw3kGWAd1BMs0osev8X93MrVXN4KnZQ11mIdTNQFjJQvqWjUL3
ilt+hBpSW3mCMO4YQJeQZABxcKNahdNu7bvZ+PDiXwixZ5KvI9+4r1FLSAs5dr5M
EBQohslBkMDIMKvE+Vbv7WmsUdqJc5NWS89ROjFHtcQ9xLZPT2Jyev8DYBTJjgK2
sxIP8JSqmEuPY8RNuwARsS+OaITJ35shBumvRsCWH8/kPFad9H6z6hSXUrh5/vWt
5xVgGhucUD3/w/5TcZlvxGyhQZm2WxU8WWqKXj8MtEmskbu80ulEk9H3+CEg5coL
1d+qQKVBX4Cw4nwwgpE3NcumBT8B39Wt7GJ9lRPqZX4zRvGxpdockSmKwYeEhRyU
V2sZhaH5bWrhhvHrVlcc+yIBgFatReyi+/UgHSAZbZswloDQA+JxvDolNDvndDB0
tP/dTA7FAxd6E0fu9R9K7Q3RAFMi4LeTqlRcBMVjhtOJl1jafClUEmx56eZVvXUa
71MkHLDdBmgBHGnp2o8ejDKQvp2TP/yotN7nVitOnA2NAWbQrG/+bZ0YDga02WJk
W13u4inZKpYwRf95YTd/VxkpYsf7kyHBnYpvpd7Fo8YNcUe4A2N8q/zCijmvZDNM
mVsWhMMDB/IpDh6JC3hLPJeCwPdDwr6Q2HgdKvTTEkacN+mEmiFOGuN+QMUXCG3i
WehIOmbbHSc2un8Ua0JaFjLkgrGWOCMINen5GZWqPWf6vwc3FyaCj18Vb7ebZf1m
cCBqkwzS2U12j2tFtg95shi8rCrTFJLRXXQoxWawtt2Qn7+UomaCvVMDGTBDzxVC
qbbxUfVunrrfPJ7VJq45hOo+3WVM+SH9fLwIWv/lxoEWJHqLMVzCra9kDgwhtd2N
0HtVhQtFVt7uwYV+1miPVZCR9F2RoQlNR1mv24pyYJBDzlWU63pWgjtZivJgqSQT
fCXuMKmiN4oykQWqbYPkvL8oulTHSQs1BPiSq2yod2lqA16jUwL914j+pEKsqir0
TokldqV19ZNGkgCJj7c/aq8uHFCa15N6O2HANAr2GV/iGY0tmLP2wBSoGc4KLkj9
6MoiezWxcvJeBkY6KDvnatPawAJJQVn/aREXwj5nkemKm+2F1nrv2DKchFCIIKp9
m01RtwqFHQUfbUXHcvaD3OuIKqCoU7S+BV5VIBdDunc4s2P1VIl0IYEFJNIS+7nH
3aMhfnf3ZZYY2zsWgkcULGg8XtHsUt2+wICuGEV3AWOX8EssM+nR9HNxnwwFUAzC
KFPLaAWBw9/gG6xVo0yFNoNP9WonN6bjb9AEIn2IzJ868qTed9j+hOvfeS8Hi72V
Ec/92dUdEPuU0sL+OV5fSdkT4Gqbk+ypfGW+PiO5QkbWyFUs0XWmWbQQLJcPewOo
MrXXFDU1nKkXYBYlWdNxFPPor+v33tw3PJ3njMGVTuovYIj1E5oarc+vzodBPj1g
hY+qqi7v5VhR7xBlohNfbLDHQqtoX7Qz+7i0deN4k+q+UUU4r7EWRNjpS33wRtNp
DToT0T2/pNmkhEeOeobA3zCbGs3tVVvOUK5iKJ8nppuUQOxDz8eMt0HXiLJf4IJR
l93oX0GJIa0GJnYWAodXet/h6acOmLfHaBSjxRj62TKX3ln9yjKIMlgJqBf4pvvJ
TEhOEkpJAvhD6T6+rxC9nidDfXgDrwZAFBtyBoiSVySe+uO/FtdGanQAZ+HWpjsu
wTldzwbgALYCh2f4shCdOZKM7NALFtEjGsWLc8PlZ9dpbcJetYG+IQ1kNo4j3/wo
pVk+lAlVAShy3zW8zXnTZWihkpBFfjsWANZ38xB6MBQHm1NU1r5Kt1MVgxBT3Uu8
OTwIHrly2FnAKqgCvxS/gpTpdHyRkwq/2nNuGqLeX3gSRu8jDA2Cc07GaHdpUUjb
LSIaSyZ05DuI4l0lXGN4rQMC6PFREeNPkBl0XwK0ScDuW/a7+Aq0dIpP9oAus72V
MzcVX8p0eI5a386BKKElyEFhfGF+JwMQ65ZOvZOSp0J+8EiOfYaRLEv7718VUnd3
7R8+ESvLMN2puA8+ksL04k4uy4JIhDp5jVID0ukmfsma/GR4WixyFEmhOZx2qlK0
o1C5PNiBP/ZRp5HqdCLiCaQhTF+XR25MTIwdIerZHOkemq+jDDV8hQfREsX9cstA
Dl4SEEzB/c4w59KB5bIa0rjQrsEQEgyrygBs4EvbXzzn0K8N3fvCk/Xydnf04f81
HJhTmyVN60Hqc+hLlrsdRrQ14AhRgrcyON2RZjfIUcOzDTCMh9x5FUxai1GFwRw5
7jYo6OdIF8UU6nNW72Kq6T4nHeDQ7lCkXu8yQq09xIJOJOzBTjfL9l2VxQCnXWGK
byXPKdrU+HHwQR+luk1w93c5s/RBQxb2xx8KrcFPEl8oM29cdbEOxnOm5KhL0ESH
bgawSwyDeHS5DUhVtljHtlkbdbNjzNKQjeSVD0IsHG/Vd7BBcGJdt9MPoIgt1lZ0
3ECpb9h/UMtgsDHrM11B+flVfUYD7ElPCMISO8Vacuy1NXKz4hbrQ9O6/dTayuNp
Ijyp09vWxwLr2YRIA/6Uq0BNkA9gs3WUF2o0fP1LdT4yh3SxEB3JdDYE7Tf8Adc0
jPaEYveFps4+NXkt8Ae1QxVWGwOnXnYV5/EyA/bjaDXWIEOmSJhd7maF59/pdf87
sR+L9r2U6115O29yxQZaIenfNZj4W/p7IzsbCxgiorzuvJHaOVUGsQ+L17M+ANga
EovJps732ueqlfde5OdphfszMz/4xcuSOHh04cqwqdGmXwTmZH5eo08JfvCqqo7g
3ziJV7yfvA+F2JU7fN2nUX+L/XSX1rufihD92vwrnWITcvd+kuKb6ptusVxccfJH
XBtewGFK8bkdJT2NVI53ZzAPRg7y60EEXO/tVe2I9FQZqqiHzt0LfemGzUvSJbzV
gR3z841zgfLq763OXRcnF5LZw3Cm2HXjUeaKMmfdzM/8nXxOTwYXt/WB846Jn85w
3PvKOlxJ9kIwXk7kUw69xin9cV4RD4nN4QevkAKKQlN/hZunOTh9YVVdi2R3IULN
xYbqdH67whxRd0BypxLnXliNI60gDpl5idlAmz2tGs3O2BuMBhSGkrVn7xm6Y6py
KCT3EBa1WYWQqd6v4qaA2kpXz2PvR3NUueJRbskz9sN5yW+y/Qb/8UJQ9oCjv/tB
nLyptH6skZs8ccng7btSBdZpVsgUaqOeqjqwwrT9G09Jcbo+Yp1VvYOLE3fgKC/U
JZmDyb9mwFN+ZJMT2Hs1YLCJldBhB7OPch1Zi45ikz76JOFy06tE6cKsjJeOZtiV
HbnWmarQBe4ehzwIrtynAP5N5C5Blb2WCZkdgUwhuAm+c9QPLPk9XtKYPAM6phtq
nBHoWwJy/A1XEwKMZ74stoABF5cQTK304IaveSzzwZIhV8kmNaJ9Z4XXXA+AQOxA
BUhf8d0d4diCvearf5yA0f16K3zgRry4yS/78XtkCVop+Pi9+6U2WU5wGIwVZSXH
5y+KJtCaNOTSN6NoUrP1Fod1Ini0di+hvgeKDH/6Awe89UKfaW+30CXUip/seLbv
JmK7gNo1OZC28hDp9+iolmqv7QPC/jmEBK74R4zZaTQr9oW5QFlfsRq5T37TaoPy
1cLkSl8RTyftPq+hFy3RqQ/Tj28KWgQSCslAOq4HnXLBVlxGH0b6ZKoDBkxcQUzx
XzESn+yGMDXSBX3sCb5bBotovldLZreL8kf6i/zCDaQiIST0L+FHCc1GxN2HQW2H
ccT15IZz995iVI3d+vgiEJsjH6HinT1RfyPcEC/N8CvQDvZREK0VCLIZPpkzeON1
ZHwClRkMkxhJERIPSdNasFYTIvcafe+Niq7mXSJn8GzTO7cG3bYB00HnVUXGwn1Y
JIg9e01OCDnfe1FrEIk4qkJzIeHm2IYdpNWjWy6nkn6LlJgaTQtXut8kYsswwXh9
8O7Goxh2L36as+2hfM+zLBUMMKEG6yzztFVVLfPr+CF6YcbM2Z4nbUUmzorFZYQ6
YIxBVWmA8cElacGLIAHpwg+ZQmuq/b2fJ7TmCfz+1/w6aFCN9z82ZLjiGwzYS5iS
Qx+MIWULjYDFMscZmVwcJsBLrvCcMo5mCP8UZANI5ogQ4O46TiVvsMD+prCXZFnQ
YQI+7UgOLMlm055+db806/axjWtzlKU3+Shd4qu/DjwMEgPhVKkhEqAlFnPBDYvu
7RwvTQj05hqbkEIKv+afLGA/FxirS8TGAXaUDcAq4F92o6DQdaLFI2lVIJwctXUf
bN/d2PtRkLnywoBD3sZ9gOETyoKxWJ4c+vbQ7CBctYYwo2sDOTMCXP4rGTWIRcNU
DNpWnhReuqd0JWCSKCXWQWVPSBJiV1s3w3MYOo3EkQVJVmlqzAIIOYgMEpa71588
+b3mwmCXhwA95m5ejRKM0dV7uq7lVOeVvRjnfTae0fd3P4wOy+epUqfrFH4Js140
jGgGF1JTYfUxhESsMpLi+swcIR4cjOQskXuSuhzQN6pLkPtJVR64yJMDkB875OU6
oyi19Vp/2QpVENwEwN6TYRyJgp+GhmWq4CCitdDCvloBs8E1H1QrM+EUzn2i66de
nXjOtnCufwFvL6JjY/nn1ZxdlDe3q0vuRF0fGvCNxuY+rsnDtd+/VnYkwBajECYr
auMCOTW5V2ynR9opL1RKFEJgNibeuUeXQI6YBDVz3c84qV50Ix4EuXErIyE1r1RN
hPgc5YOwK2oYNToIbkDm21TCrWjtQXTjucyjRrwnaJ2jH1ViSIdtXph5LKK87qjV
NpEzFBXUYA82SGCo00hBW50Qzzi5Oar7ULrJwvqgMR/m/G9R+4X6yvkfmpOW6rqz
nmeO8iOQx8RfrNMquuww3Og1sv/CTxoT/Wt5ISJnjt/pj1V3wkpDmyaLjlQTJoXT
PtqegL9hUAnEH8K6twvH1cT4jxckv/gAUaM1Tcsoa2l/zu+dHmQ11ZU+TZKlXcns
yCeuI5Sqb8+yu5AuuXbZJsGMaimngghYMxATnJ1UM2P6DGguRIPfAVkj8t7kjVGK
vK2m817J9nvLzJjEDhwaJSlpaFOviJf6lScoLjn6Dwu01wbqyc7qls9iH6wajMTO
o2umyJOt59tZN0eyQnhKvAESo9kL33O65nC1LWNsk6NlaHzy0anF2OknrFg7QIs7
x8ZeYdlwCYBnyEAdf9x0mWmOnDN7qdCXAjxBEveM8fT7zHLh8YgnAo3k2pZ8syDb
ulLE94L0qx+Vg+rxGzE1nNMRC9R4cAZgY3UXwHsLjeQh/iN6P1jXfila9Vs7HCWc
DgEjSOzCkf6ZthXnLM97IPsgF4+k0s/DBhdOOVpX+G5nh4bLdk/IL7mGg/NaQqK9
ugeqvPEkKATmqQ+4anWNhY9yQ4hkXsrNdQQLx+wB03FlLeEMCwwF4Bde6U/9rwyv
nuTwQqm2P7wNdnhlT+eWV+mi0ZvBOd311OTDu6RR5X51tf5LhhDp9wjKJH1iYNEa
80sUDR52RMLbvezXIKrI2TrwLukks1RxlsDKo3NRhogm3IGE4zwACOwswkW79e7o
Bb5YTpGRfIYJVLZq7SEIr0OPKrP+1PIYpmBa73uPLBeHxAgmac6ay+4nArOXABNA
BlC9FZ4E9A8FUArKfwR2xt00ukwvOWW+3uphoce1rhmDPIvy0K3hEHqaGEhAoS4K
2ZuNds7UCeGU8oZVemxzgdvLVgP8Nk/OK8SZBEfEk08LxMAkUlOcfesS+9sHiKWQ
oxoHoM8lAnvWvpgV28RTaZFrG/iKrS+vvq1eqMYka1hDyUmgxnyaWbFzhYk7pONg
rXitOqcJ0vjb3QHziwRp1R3VRsPr799ldCMt9dRkEYnaT0oKm4imcZVVRqjdkskJ
Cq+jYPOZrgvLMm+hW2ytYSrPPmOtrIhdtOInFawEu0uw3WSm53xusqzF/ath3Emh
Zqcl69hVsK7qxWE8y78LQwxB7vVg17/Pmk7xxJoqaEYQX9zib57TgxZZAihGpWLU
kuY4dFN1uc9IBIrqdsA3UbzmO+1rk0joTzWZqJ4ezFet98hYSdVN/xVGxKL4MRi+
wfspKihtG05kRfN/cdBS3+z+UMjX8cHECFRmX8atuWYK1L942poDmJPSWcf+H+EX
t78RP7HDpA92DYRyBL4WUxrPGsBMyv75o8erQlBtNj+qRXtQl22pFL9El2HUGJ0f
n9rPB2rWHNa/mMoXoRGo58JMBXPmDExhSe9Wa2R3om2fnSseG2cNOqitPamKpABP
IVlKgozUdFfhYqeg7LckkIfwZ9rqSXm2h+JGRrymgcI1J0TXCnRhLmG120ajNjsq
TYCP8W8yRo+hj9RZ7TV9nP35eCdWKbdowBVMlbEtcXhVEJZQ3pme16QF3pwJorze
GkUV/5OmBjSsJBMMFuW/fLn8thnkSdQ3PLZ9udZ7XhTl9xAWeztU9/32ffphd62c
MzMyP/khp1W4bD5ivmLrnOS0TPUPkqiVRDvoiLtIbpqSYwKXEoMuRHdYChnise6g
/4KYUVo+sAdlWs0HtlFAEAL4b1zKo1i1Z9GlqOENiUpWgzvPx6lQwUb/QW89mHIB
hHzibbx17VaVT1KIM5eny9qMU5lW1jRL6tXZLeY12+tJq/XGdK0cTfQnOOnVCyWF
ApUNlboWkI3kMZn4yIly4ksabU3ol45BVBUtTFDB3vAT9g71ADslHlrx5V4hWLlE
MErwA2CmMR8iUhOIk738wUWMDuRXDPvI3/p1wvLwa2nXpqIYo5S1vvc6PPUEC6dQ
NZsjNGJbVHOwf8EVATpYzr7AR+jJnUyRolGQ9fWnAvy+cDW+QIbBZ0fAPWztlxkh
uHAuWdzEV0BwtB1b6xBI9TMD6JKYwO+ZLVmYq84WeoICfehkJkso7OipNCTMY4wb
y5a5gwDg/X6PQvCJDe+EXih5VF9osy7gbSNZPIfCVSXkLwU8vsQQjtAO/0Q3PgUf
yTl8xbIFRzG/E2m0VF9CoS/atehUQeYuyLX4kzClocU//lKYdw3A7PVS/67wKkNS
HHcZGw5Z6qbpPI1YwCtRgBM0ShUJH7lRcYBKwBObbvCb3OOPbrbT/ZxuqMnqHntx
lAK/cUZWmikCqa98k/JhwBDrrtzMU8cIA9k2KlT7u17I3EnCT0/3QzRUn3ZKmKDv
GdD5uBiYZzXGL+nYCjawBvAuQssvktowLC7lDy/KS/qE15bzupB/NyzGIpv3rHTs
Gu7AXoRcIFQnWqFBz+29F7y4XEzubJZV+s5mVtQua+yrMP/kxJwJIYVPQ5ZvbDNW
eiNlm1RG7h/FJAjgoyEk42BguTqaAEyxAMxjVax7Xc+wjPn3m5e2t2yBqUniKcaY
pkXO8k8CBvfKvP7KEjQz+R2K1w0pMARAiHtXmU0xQYqlyjRBEV8Xoh2sUiBeOjnr
7bvOJnSMu7bnGk+Ar9Zz++IY6OF79lLgIfpU97rIhd1hl9dsTuYnOKUSeJ7cxomx
mgGTGOyoLm+Ov3T/zJSbPxqECaGHr1Wvv2leTvXpKrh3La1IyKtLjgDu3JLQvDhY
0IC+QZ1XkT5OErGhkdh0A/QPZmxZ0soVbfalrUw4ns40shLpMRiYI0jWann8iQ8q
Eyg9vbvOWPq+91CwV3xwLG1uM9jE+0hwEMH0tj6226w1sxIE6XOjUNSRnKQQo8LH
MJU+QBEL5Vif+Fq/VOs92ijw/TL/lpEOsr2TptQfdJMZZpSDjRoZRFxLiCBbRMf/
6+rU/n6nGX6+1tfwZIcPZC3hFaEehN+D7s3U/ZOaFfWxX+AP8PEK3D76ttx8f6YE
p1SyXC0DtKTGumAlpyqv9X/UiGhlmMPj9IxzqAfo98XCUSt+kOzuIYxeUgvw3GGY
oTHbRhj12ILKV+SV4HsZJcd4edl+VtsOR0PCSFiUO2V21k1BnQxo9zf4JI+ttIXI
SPK1+p/G/k44FUNvyiTYViOjaVooF27/15aHaXuIzNnP23oeDBwfM5f+/0PMXc7g
W9az+7z89iXn8YX8l6y7kbOSKMeqyDvgi6ppIqeq9gAvNK9esgxR4fnNM4pwL/6Q
VFYBNs/V+2OkQsnLU5JqKnrGl7/j9W0hfE55RG6L5QgqK+WS75SSBD3EgtPF1FLw
sU6jb8Y62YlwrYu8gMBUj8v7b8VY3tBIK4vbbuBgD4AvCDDE9FRz4gu0DTwYPCUa
Gv7gkESMH0NmL+w2rb28QIBgZukrBgl+6+7WhMdNgjrUeRkX+P0keq/4EAYn5XTK
OhEErHwLdAfLs/WALtxULXo4O4NscuYI+Eucyyhhy7JS4nFUxajWSjMGXlqYfCOI
420au7PYbqbNtcq2dyomhBawZJ528kjuj5NhjT6tHxrtpVZsP5XGcyZ7Z4No8Cz8
ZAGHKldOM0QRiTxxymSJmbNuR5dzAB05hkJVQ9h9hxm7a1BQF6assV8t1riFwAhO
PJ9Utm5eJvokdWkZZFe8UBVOY970XX2lvLmJM2HEFauW4QYzcz0V955AgOZHLA89
4J6hOvzhjKgMj+VECxkh3AbRhIsq00+yBC3Z7C7g6LCYgWWFFyWgj35xRrQSLQ5n
gMhEKB8q69qdvmyOeSntmpKhmE6t6olgCbsnOdoKAYaRMEQo0KRI0aqyGHe/NBkg
Sn5Fx5wVPtSt/v5maSfUGSqPzkUGoVlgEqk5fNrF5qFaEGbg1DQH/Dqp98KcKxXn
pMUY8Aju7NkarNM3RtHfioC91Kirt0smjEUvY6D4rWmD7JXTJrfPlniI7ltvOmQ+
0BiIp16taw9lBNjqdGEhnkxTcfFYY5ActaVJzz+/Pv9m1gKHikMm57Btc98pqr9h
PV7DcdWY9HCnZMADM68OqDKxjm+hIQkgCRW3hgUVR7NrgYCW6+gY4P0PUn2g8sFq
sV4RivM0EQuqoFa8A9TZFdod41eNbmR9yzxtMFICNDpkAVGonmm1Tv7nxnHNmbjL
EMWnGfFCp6vENME8R5B94QCKzkVS4+GqxAwukla631F3TyrPZkgauFZx3UZDik2I
JR99EIwUFCCpgxwND5/9N6mTWEgTL9XJoBBCminzIZzqB75pihluXt3BXxQ92bvn
FvIiqASpviSTiv/ZA4QgEKQoFG4vqakNQ6nAK84Wnn7eB2nUfBUG7HTM+l3SkvfO
lcMQ8zCoVH3Zi1I93VLtFa/w0pTbV3+2zOYCiZxLV4ETCS0nwG2g/bm8OHqZH3Sl
W3EEDt9tXaldPPyWganl3T9x+fuxtT+uBJxQmKb7fXHRbNFEk7HZlvMZ5AWDwhLO
ODc3utKrEtp/HMncYc7xNEphpbrUIe+qaFHJxmn2CBr1Nwo7kvNGOrrAI2JmJOKD
yqrVeMrfTTckQ+O4wrI2SnaS6pbZXIO6g+DgmGrfk6Kl1krL5O802G1cYmVpmpBs
jrQjBiUfOf6qOE922NDgijRTWedUb06PrL/tIcNXCH36PmfR2EamGHBRM1q+t1Lc
boyjooiEDfneB0/69cVL+XZNik8PXyQAi3SpUi1SVaQoCF6nxGfqnjiI2HO92auO
zDDGPy/TVQ0744G2kIXQN1eIag99rtPSlmIEbb9FPMLp+Yhk5RyqffzQrfUsh5Rj
6sxOUjmJoEiB8S4v1SAldvGxQjlDgyzeQ0VhhtlvLSnH6b+5gH5qIhanS9Sl1il7
D3B+xAAogt9u21URuBfoE8cLdDgTjeGb/p1NcWHkJqH7flnddLlPXivmjuXEQpkn
XQzubA2P4+7AMp9WU0AN4AeZ0khTfoNz4W1h2iXikrGZ+TyODOlPo+6s3cxl9kym
hP/CVByo6yFUSLAvE5JY1Y389KARb9n7JCgl8Lf8SQQ67B3mBgYIk8vjqhFpm+VG
nMufqCAb/a5WLTGqaMAE0wief5UMpTeaLH4cRlX4MtVNDZiOz0uyIktIL7IburXD
LeV5XhJr8QZBFeWkq98bcLeLAQVaVB2Rod4cAKASPIR2/tZTJtOPJ6JkxQtuRiFM
Vxqhlgm0eryqEgNegmJmfq3n40aM6R2WE4fZwMDIvAMQvvmjRZazpxWKMNsSeeJg
+FzgLI7uPmb+Sr13TvzYnb3zOHmHhz97gjt0Tud5GyPVrAwhizE7zYWqSXW5ISb9
iauEm76z3LSpJmJTdWR3b08zWc83D7SxTpsxHleAVEEnb5rVO0G6HrlLFMuAaS10
L/wbaSLEV2vjsp4rtwYfeyJLrSKnfzGHrZJ5Hz8tLzvN3D8V40z7kG3JuqbYh4hf
rOjAkETycZmhb29nu3U3ccZbQJ4sfiF4dbxEt41lUKzyLKt0Ah32ER+k/vofbgej
PD4uHDeI2whfPnLJST7L02pIWdrJoBKxP/zQIr4gYXNMBcywxB06Jdm0wPo9Gbxw
FR39MqIuvp+wM+s85R82jDoiHUhKGZ2Yv6hggeOBCS543ryPlUL2W1kShjb4ZxZI
CG46YFDuEQjsNBt5b9uT9D9k/A2Ae4gLXyvRbtFoYvMT5a/mlM2P0emCI6Nt8n6P
oRNJx6j++gOxc30QFE2C177jWZb16QVQZlOS2HmMtk3GUqqlncxEI4g6xxWlJ0mw
HcK5gn/yqxoMHShs+5ZgxxMGVj+/3Z7NURB/5euYHwPvbDJ4j8zv+bhoZ3ahqIQ9
MjSrFhJdZ0rzO+xVcN1QBJ9Hq9oM9Uok4iof5fToF6r0ybj18NXewGmkMsbggj2G
9X9twrXWGprEL7ATGOq6J+T+XAaBdvKXTQE/enZ3WvQnj0eq1A1CPtZIFhPsJtas
rjTY+c83W6JyHQYsgEbKmE27p6PPq2u1BhQ4xOCYoGv86hNeMqqccEslBbyUzoVR
ujayQmdBBnS4iOLAUArUDl7JTLO7gscbvg0Csv1ENUWz7mDRkjcwoLpI+flXwxjN
m+ATilHQ9pHekddCcWs73OGV1TnrGDRXIDgFDHOM8xSjgn7KQSHeZCj5ZNUKaJz/
/84SASdqoYtAbAas29RYRsjn/8p6IrSxUnDzm3afCCZuzRV1aVd2T1MsteyA1ff+
qv8VU/4mcU87jeNqmw8OiYJVy1EdLPy/ECuAaM4QrbH50Sm/n5i5JGC4en2Mkpav
/nsLUVPGRN2eJiizmv0fblyr6gLlwJklJH73govd/Hb2ZJy4/IXA3RGHkU+tdPyu
ee44vIR6Al0p/0UhVl5VU+wN7KejMHc7sl9FWZgGFmS/3/8rNutOh6aJo5CqGpbj
RUEuWvx7maxNsXFbqRmKvJIuZhRtwJAfwCn7dP1wsqO2zuQWKnpI37HhJ2I4/fFQ
121KHcSBn+eMCtj2iZxRfUPr7zzMrKMAu7rMRSGasu2fTMTvZxK6/howowVdlDFc
Dl2Ey/B6X3BxcFbeTMCM6pr28V7lGKHr8HLu/eI7/iUXx9/Eei6pOSqeS15/KBQ4
SAWE1yIFtlgtnPzRpP5266iCsGhUDoUilbrckb9S1pnyiKWgm+zengEEuw14WdU+
/PpyVqGu4b6LZrS/P7V5ODcIDbNvLyTcphjepBcONBKnd6XJl0druZeNRnEVAr9j
5qUNamG+eSVEQm5I+X2ulAGJtU9Bl+MuHNVaosQ2qEw7TAOCUE4XcIxCk1mjNCmc
6cb9LkP1QWWgEEdH8KbvVx6O7EwOvYPwNhemil71NI5xB69OzqBSJLyRJ/5z4vwm
nzZZzI+iChReiCXBZO0Nm6xF4u4/RlOsOEkMf9kvRYPa5SrpD9kGWGQpyT9UtLAV
pumY87iPck/NTF1nEaArWg1cxYoRLScBFeFsSQZ/5c4HxZsA0U47eQr+ZfbaU0wA
AdF/3vDGCYszESQ97pbnUuQ3FQfg0xIC+tPVq51WxrrPjYvRZbBEEkykinVatxOx
88HvbL0t2tEz5mR9XcRATkg76+orfwFtquBv7WoBSF/wHHEbXPk1Z+D5dKVzfgH8
pBGQPy7u2NpH+pczcVVrxnql2nj3n0GA4ZVXDFTtmRe+FzeRZ2Iyz7ahtrfpc7iY
Jq38IJoPCbeXGZhqpbQ704JM3gtaMya5fGlHeZcDcbCtz1U835DyiYHgHQAev+pE
Ge+BJPqivQkY0PHUiy9dgj9Jp83kfDe9oMupUbJvkCUjXJm7ZtzV5BbeP3vWqC1S
yZHMqDfFMnh7hh2YTyB16qEeZRsTKESv10ZkPMNXbf4ZNs7Ly3tzFa7pa1MTI7yM
zhC1LiMnaA3er9ErhXZECY4KwVQ1XO8nw14xIs1nR18AVYuDpw+WyOF4l4imwUCf
kBf91uNUafaYNgBzrtMBGz4mTMsYrHGnmNa15WmFEpJkp6+/A5IflAYOIz9nZvk9
dvNSQU7TDDyJ99rUHcgrQpapWGvz2r9/nTuUM8iGOnWUXlnu7gRsRjJ4pcyK7jo5
FM3El37aJoOD220kxNGQajtIGPZeTJzSPrw8PxnKmCeGTHIpa0nXcNaO/L+oU014
cpfYmcAOioP2wEj+Vbf8XbQlIoJ77zJH8q0+Nxrz30EdzdhtxK6niXORlkfVKjel
ElNvTzgsmrBIGxuLmikJK/3xN3cXH3QB0BnraZtQ/tFIJ/6YOskHwl9OOnWqIfCC
jZKGHmT6Wu3j2oq3UNhbRMwnVFvkDsrLgpxAzqSZYpSfHdRbAhJVdy0KJ2lEbOQ6
VWCl6LZMvJWZ4yXQ66mIlq96/npqsFCviBjaFnEcLS4eh2kt16JhSu+384BnKJ4Z
fofPgdG8z7L+9wi7HKmF5pAbXZ1v+urvOTyrlcD0kcgsOF9UtORuzaWIXvvga3Sh
/CqOK28Zw7r/ASoFxWed9X1rr3XQfJl+7ZtSIWTbZpgZcmQfLu+zw4WI+9yyW/Np
Zxs9G/C299MvTIGuz4aKDvb5m5eH0CFsm8KEJjNTGT33LfiyyWKap/dosUbIsA/Z
Lt/M8mOPDUlJ381JTDhuADxAY14Zx6QfuIUdYYJyCR+24NFbYLtaB18JmiRuP7qe
FQd62yjD7RC46KZRvRdVFGOLu/TetDo06lbiv05ar0MVvuISd4UNa4JvYFu2DJaa
jOh2dZQyDC7WFT4S86oYUfoK3wwTSHQGVR4W5ywaUO7sQ7raJ2n2fou8Clx/+jJr
zxRMadg4KdMgljHHq/2hTO7R6YX43Gcq+CLk+AhHCKvgSnrAZ4L3zkJJ7LgumiZ+
rTIES02D8gqbM4TtmKgGs10OGqUJtvJWholpTfrDWpvS+Ji6spDHKcr9nTUQKY7K
L9lLyaX4Vv7YVeuWqcDZkSihkfa19bRpgo8EByGaHg2Jf7KUDO2LrbvS2eNQ45BO
DtWd5Pq+Z9V9Dd98JJspN2z7mBSYY3C3tquxST70XHAFixAcheSD08Ok+PDMS/ZM
+NWIuFvebUagqPq/Cp8orvH/28DcUagNjHC4MAlL6EkWNC1E8Jkmy3Hl9Lm5vEqv
0m0OjbDmYElIVERzsDuSfyuztckS17dQUxZjxD5TFXdCoY0Aompy/ADDmuFw04SC
PAkVhvzI/p7NkAx4NBl6WYbIIHwa6WB5p/hIEbxnEPd0foreNw96C1HJIKrOS5T8
BYoPA66GOdoTAPApszjP8mSnqcQJ1AUMf55gvMCplJM9WKEAiFREhkmT3lcGvTq6
nhlqKiwY2ty1MNW0BG7xvhabyD/RoHW4GvpydQon/q6gU2hPb1i5IADLlRuGM8tC
A08JHjlI2LtVEaDW1ZXG3qeyw4IO0LJQq5KqmbpGlOpuMmSTFvy3GNT0VYKXDyQn
RJocZuKZTEa4+rLsiGPWd2t6SNl6hemfS6c1Z01HV3l6UZr35n3v0ZmNKxKQP6vK
o2Nl8npSGN/gh1B/nCD4Al41nFiYIx3x2b2PukQV6w8AooyCwysnc7aai1K5XOfS
2Otpea7XbsxtsJMJLxdBJvsuvmQePwkD46c3KeUbh8yhlBdHkUHEPpzEAG9fUbqE
W6idPEJ/CbFE64i+mXiQhpNe7FRezXx8S7GUur5AsLgfqT4n4ik0ev9fgZ8oYRGB
ZEVJtARKGjysAJ9ulIFGhWqkyBd5DF0iuSi9xDI4vkG3N6rnagsZoKO48A0O/zUm
sKoozVZ+zpkReS6OP2fYvK/l+D57p53VtSjAoVdssFZENjxDzDFhITGwZS2qrXk+
ceQaLT6E8MJWNOpJSnfiAaHnCPbLHRkNoNt8dkjK6RCJVgf7okJNDC/YyjbUrM8/
zdXIhA1uxDAFsAHtljLBWLoSWAAzeq/vnxQgpTdUg0I3SdAO1m6eRRwbpmnYECVV
h7O0owD3uwfmnsZz2hz8VN0t7aju89z+Iwg81SERGOdrp6VPjEVOi6KUsd1bn/O9
2/nCfs8lIQnerJqnhy5ACza9QxfAOLAtNnnC0arERugPTbpaO6g4FdBLiFRXv0yb
eU6aUKRvvNwJgsbFykMN/+Ntg2Dp3uMLRlTU4eBDOPwbwibUXKwuJAqNomZqH/26
3Pqr8W8Q1UNCC333VtpnpjRIUn3/IooJAEO2MwjWw1z011d9hlG1rfWrq5GAOumE
ud0cXDLz03+d/dhiDWoV+98yLRC5aI0bBrolJdM0SENgaBFXQmz3Cpg560npIwBt
xL2K44qqdfDiNDV8aHhwVEM7FqZNn7eOgh/R7YuOhnwKBwgc+BzL2N25JSLzFaDF
mdg2YZ2ukwAGFrJauB7VOtzqA39wRJTawgaDPZ34hUCG2CsUt0aVMXjV2E4dy/q9
WMjs9qFlkfvxTZuOcZwwv7wPXlT6+CBXNeL24oXWQo39LF6ZHboVjKgcrqYx8ys+
iWE2Gi3UV31XV+ritUYoDAUoRuYVXG/VQd6hDGS4JKnI5Krhbuz30lDBAXRM83hU
lQtWlmIByzlNDr6Wz/pX8sEEFPgJFrZ34eMpBwy08MOMiueUKEsAKyLGbJWGfh/O
YfuHWsV2098yEJqw2nI9TJ0QA3ZkeF51jmDIi0LU4zygeh68u5QahEF2WcjIqUFL
KinHSUzH+IAa7OmBBhwoBv01uAeI9YPS9A8ANX4H7CBqEBVj9ZU8QkcyLey4YUJW
3zAbGmj2h1lnEtEsZIDtoYYJhI2PiBD9nGTWYGOKwxIa/zYpkmdUmp/MTBuDcrUN
6fKRpsCzf2K/WNs54SW947QJwp8JGNuasG3YN3z4tffXVvf0F46E4sDD4GtRNVgV
V0CSswTjyPNMD+tB+6NyH+g3rH67ak4QwoYaSOQ09O/w5E/CPsf0Clj8Pb0wAx0a
7WHw2Fv0KcmhdF6OKTS/FJpDfVPBbUQIbOCzt1j8TwUfO7wFwQZkwMwwYw7STVmD
9C7Q5m2Q+FWf/yPKBWmiq5rtrhPESQ5R6Cy0goouJjWiVqyo4bkbc6vRCOnhTEYi
fGhTFHTlbTnqEr1zqJBCdxMdB3+Aw0v/61YZfk4xBKs6e50IEA3eR2b7+TczGQMn
KTUyyYWNq+LP+lQcrmOe8ora63m+TnbXn3xmrEzuQXHazUw8MgMwkbAuEGDwCHMl
gtnHXn8pTziRkUTGz0Iv3wJ6Y8V9nIuvgm1psgKFeP52z8g+SU1GEYpvYlDq3Vgs
3rUV9tEsbLqIICU0RkTpdG24zIIBJLJgbMEOTJa4bAbEOG0poZZ6Ociw/mZnzkNK
jfbFyYWVnOnXfJ+uzv5atdVxatu6pRn1gzfeLU/Z4541rhTiJd/pnbEz4inBYjkk
JkGodZOSjEbeOKcKqTHtzcv8EF0qIKnEGSfEcRXBE9qS4Zs7p7lQAuTZAmlDDqP1
k+xFdHjojYGgCeMFhnaMMuLq4yYu4UJvousOeBcfx5wRHLkwdP88MThJgaTVmzo8
aozo/OrouD0DyaMHMUYWxlLAVWgA+wxaSO3Yelr/zX0ES5w5XzDLTZvzk60LfsCE
Yu7y+vFeW8vSj1C6kfHh1vh/Z2Skpoid8lVzB+SGiynxLPXBVr413L0CUU9Phrg1
7UvL9i4L/6VcoXvbMNtAuyJB3tecBtpVRcJCLPwCla/tK/Q2TEftOCbdU7nilWgM
0KtMndDDJifZ/gSr3s929rrD3Oeo+UejVMwRbtStnr4BHFb7m29CouCxuk3CUOKE
mwZi+74g9XDfs6lYiHMnRpdaXwV9x9OwmY1jI2BZDdYsjCBEo8m/eGVOyWOCNZbX
AEXUz5+5RpdFhef1wtTj4prOHd2KroOxQE9xN8Y8wHiFr+ozhQmD9WU+WC3mo3uP
97gGgkQXSKPqdDqF9qkwiV1Zt/pC+zTNTb96J8ZoeZhKqL1C/zvwPWUu0yWXpADk
Is8KYQDcWEH1ZIf4Ls2jGMj+TZtYzw2fExJahQb5wAJFhR12cOy7U+IrqgJQuClC
0Nc6v8Vo66j0IlSJy6I3S84HjKGQbyNqH6UVMo2+WStwVBMH9PcZjKTUxPOTOwQl
mlttqm8Lm60DKmlfaPLaIJTCGO89clfJEUjO4JrbA+bipGCTQ8p/WvEdQ1D+h7QC
FJLT/Ikof1uiD4PocfulCgGPPG8T2aZL4Qmept17WkqRtkc7mxoJTP6ISlNJP5PD
ON8g2Xqx80/85jkDDclhYMqExVWUCYCW8T49SG+gqgWrQI+kRGUFuByL2KOVhexp
yUPC9NAy7lkQCcW23JaiFDqgA418PXS82/KRvCRQ2hWnVp+9O8rPOAGDrzsEHI3G
mFu9Z0UQrdJ0yjIqCQFf4r6n3Lrjcu441CyaJBS/ILLojBl6dpzsrc7O552fxstr
028uICsbejeozF35ocTjS69fUWeabhZK9zE4PqWqba1TLnYUjuyGWwSqQliEVuGs
D4qeRvZ88WLAkp1wMsggmY533yPTKr7bbBc7kank3b1ViRNVFi39Zf6QhN2apeEo
kul9SnHjhaIMjNcWAnTVnTGvAPGwOVJdf2tlDzSH2LjIp5L7XrHrYs2Ckl3lPFYZ
7LOaT2n9YUECl6lTrBehv5h8wyQrJdfE5PeYCtkXIvJgv1ZNF5q976gko33AcJey
I6nyqzeGS7um7Bs+8n9WzfTtCDNnDAaKYXb2gWQE/iPqkFbOJlNCTdnGjzRBVY08
z4ITKjpbp/xqgLNp7r1nzmF2BPT1SF4vaNoSdNUiBw96s2QzgDQK+cF0dJwjD3kX
EGGahS7LP+02xyxzgiuaBr3hJFi5amdTUZOdU9j5s2i9Y1fnS+sa3Hb6rdF6tD0U
JkMbJeMbkpbX6egkQIFi61EYvnQe8Ck1712SuILlGhfdK2k5QkXnpj85hKE0IZx4
PJIZiTA2FGN6+phkPtVw6zSkEHk912Yf+NavwEO5Vfhq5Me6m1tUX3ub0dQOEHNF
w51ga2/ub6t/JEFm1ULx2hZZuJLGVrEszabzGkiVaXPX5OAmURheIiWR5KXFA4nZ
Yi39/4RNpQy7GywBBPGR5OtvgAuLpOMLq/lLdhYFUVynlx6olQCk3rqYMcOnFuPq
gkHcgmsWmM/BLPzz6ZNucOuEQD2/kSEy4DfwMrv/qRgpim1cK2ibiBUbU/Um4nJX
qEOpJnfC8mcRJM6XrX7nPaw5J+5Lm7ZSm2Kwb3O14R/Gghiwmud2jxmiiUfIMScJ
goRIow2t6TqmpPgVKyW1Fom1HCOD2/oMYIs1ir6uECczV65nyxQswqlGW7DMfXZt
ej8qKSALCterf/DuVOfnSRVtAOonqCETOvSpodJZUeuPbLtyRObfkPcitfcmxK/k
5Qj0d2i5a2NxG3A3M279IglurxOgJraoTCgwW0w+lMj7fb5lnS70QuGr2nhUDn+Q
mYKPuAEKGWNahssV5y7AGtWhk1xDuNKoEO8qM9YYgJ6PO/E8/JgqQGUeaxdeu9gH
MHhqVLw6oUp6JjBS5K4W+ki0Ln9vbvGhN6HklYHIZ6msHT8Fiatv39S7WQHVTnKN
yc3Ypk3mvBEHpl4Y29UJoOv3VLE/EWYrLiJ7ut7IYBlnzJogRnbozf+h8hRyate/
d005jstoMdttk/Qz+EHFfTzd3+zB+xIeSi9V08+e5uhfjaMo07fiva/SwFf7k0Po
IyDVkvvyL4hK4tjbDiSwmBJYLM44hAc3YFGXelKPitki2rz8M7yNTWMArNgCOR9/
IEoi0YKJmRtdnSnFRrdPtWEFj4AViSjyjIrjFJiu8+0OAqI1pIGS1pcGappF69AB
7q+RF3YQ1lLkujTNRs6L8R3CUM1Ik5uBBHZLq5ZkVp1WzjRrfjUN94vDxinynIqP
nNsUBFOxU3jG0vOAkWt6E4Aq/c6YiQ5bChOtrFFDBbWiZNtqSwhTUk6PBymCggNm
NuJEuhTcEx1zNHn4NJBnE2KsQsACiR7ofNMTezyblCvHEg5SBc1xFau2DshHrVPA
+ECqUmYTwfrqabxBRFFtQ6V0/yL1QwV5LPNHCNLNYz3feuxm3huPqn8vVz6Q/cPF
mNSYMLiTLss//BiXJQ/EP8Z2cEaA6CizobkE/7d3bhznl7fXCXdZYdMG62yUaBO/
HtXvRibCLJgNMHU7wYTOK6alfr4g9VShvg+Ib0V0+/dl42+2xBNbgb0S4igWQIQL
ywRHJ+lgg4zeNaCbXAEwjHSxPg50RlQ+f0RKwTN67ww/GbbXm8oP3Lv9sEqsgU9w
ydR2WmtNGgodHBrkY6B/LtRwdy1ZanEjL3qMKuHR118Rrpks+WaJKlOTmuEVB7NA
a1Qhjd3O/203vvSG8iXVTsSiYvvjY0moyc9Hj3lM/B3oudM1HqBZe1+RDDjgOrI+
rKDoh6SbTQyUkQoN+u7XulcFhXAur1igxqGzTmWMdiYUmJEZUaNYGpl//MrCQtTm
blHi9smv6AeNVCU6O1iILZiv07Yq2GwaW7q+clydjs42i73orN1yCKx95TZw5RFP
Rz6MjOA9r7H+4qjYGxpB7lgYzLuSmd73vvj/A1Hg6UgC/2S1ZxXs7MCU2Ijaqxq2
h/A+ELnJB52G6FY3mA8YuVU5BDGEiXpEzLjYtawyeobXaOWiGVPDnFdaw69PuSCW
G5/5a25GL6CX+yHPw3s7QfcjO4XkqKaoDl/CmHHPxkUhO13bS4tGAhX0U3NlrtE3
xD1m0fDxFPVYAdbFszi4mwgshPHzIQnQEM57qrEnG+VgusgroyoSq7vzLUbVM52J
EcjvdAX+PlXACWBDiCA63thyvfwmbSSLtLcUt3QXwjRdQ+r7v+FRWG3L/nmqISTG
qqC5urL43caPVuDLnIoB6/Ru54gXVeRCj7aTcPaexKt5AYd/dFr19kNDcnpcTs5O
cfz8C8biWQadyARHqqweezEcOUhdrya2JUENRcRnCzGz5JQFd5/UBr4f+nqeq2VI
VV+PVh/mmFhcR7IDpJOhFXRNQwVGuQTMDilnpWlJfqKvpwsCvQ5mLc1JWqM7QUZY
k5MzfBYJli5uAae3EOn6G6UICzTscV/c8Q+xnWZHhHYav46e1FNyJcCNltkCNF/e
kONWmC/+80mBwGAEuh6hEvCAUQednWAb4D9AxEMLJSF1OUzqxIfEefDU9AOxg6vk
gRjrzh40HWh1yOsUOXQGn5GHGzUAbZPoUcPg+NtGNmk7KlOUgZ780fdulTHyMz5p
vusvJVL6zjGL0dkTqtI8AkP2KUv9yyZ/cKDjMPu/XAxajNMRQEwwe4VpSdzeGZLF
yMF2yjZmHlIlr433EDuWXt4Bw42Ts9AOjrrAn02BLGdV7hPIf8tC75EPDQUIYYh7
A0SO5iDM5UogqD1Gw/YLUyT8yiIVM9DfM+6m/1KxOhEDSWbt3VypCivsC2RHOPP/
v9AkRbN0T2CIJLu6MEFSEOcvAJgOx3ZWqD1R/4pjB4PsxilDxO3fDfUs5s13rKHJ
2+1tntmvFDx50T4vTZVwIcEt0xpth8ZTWLVrLtEbim4O+xJfRXtPagvvn+LTJqbD
tWy6DG1PM1EkePjMS49tlXa7aEVQQupbWJGzIzIldr/OJocG82y7oKXkqfBZXT9V
/7MKVYB1zayp2Dz4HPUsUD16BnOm4kZjZm+Lvl+7v+w0Aw2pMnu/jv+Dd7Yaltlx
6VPHLKD+Ik/jvDtMF2NGdix91+iEbZvG1QZJ0qj8gI64mttZupdTFb59QKOQs/J8
bj375xYRDCdrtHSa1gi2J1JBBYWfzq6fKhPDrK9N9zf9FdG3SOXEcLHZ7/8YEc9H
LFcKbUzaGDbxs8TCF7P0g45+elchi/oUTUHp/i3QIMPd1nme+nlUaAmkM0xPWCc+
GhArS+qHp5HNKfILLO5f/ntw535rhJatC0vY4IRw7j6hB66Okb0wD4zR6Loszgez
dXYhoHsdqm3hIYNK8Ve2trD8pZLJ0gg7HXNCBDHpyjnmLhueR6Qnyx9oUHKtOcaM
f4XnbFu8kozHeB9LLqCzrGV7nnWmE7jeAegXheU0kC2ZgNlwTVcXgTgQXv7WRm3J
Y+8OiRHDXph0BlYN0/tbjbGxQ9kkyGcaPa8OODKma+WYmWtSyUwYEeXz67kOatiD
RqKhYQoSo/w/Ju+TWNrxRurlZFS/lGKCelEUVSs5cwDweL/TdJN173546GFCvyNz
ypWsqLtq2f6AfoJ/QY3WEkYeY2o/FugmjTtn1+p+98i8hTRFbcjFqaoPm2dIwKaP
+mHT823H7ii+KQ7C09/dN9tXcksk2rR36ya0Q9W51cOScWxTwgK4hvvGuqMsWSfw
XvoBWe5Y+DTw72Rpfu70TCC16yRCpgo/X72fX8sJOOkhzYcFnHUtMdhJDVtdqFRq
4riDHboo9jZXXEZx3qSWd9pxWqpFw2nzgRkKEieshCHVHdk51pHzY/uv7BeM8zR1
7O3kcgDluHwNGxqwQ52v/yWlVgq74+Tv7o4cpxicW2+gUmwPsRjxksL6LIbtlr6B
D20nZcsdcYnMvi22N0ururZYha+QH/GsvnRyFN48b5J9HUfMuDcl0bm1P58ctO6Q
D8eeorMKO31JQKs888UwBJyybrodrE/B20Ev2Ip7AeVCcCyjoXXyEN61Ee8CMlDI
Z6lV3iwM/85Xyz3QjQFOpDVdt4wuFjyCAD9/v4uVy32SM30Od309pYkxNkZfUB5u
gDPkeAM+/T77CG9vH1GCzEqdTFjiPpQoul2fZyZk7ZTlhFkNorZ/bYN6tIRM5sgD
WC3FuVyehKG26aNUSbNGD40OB1h/AJqgpODjGjpp+bpUNLoKfcdvFpfB3+FNaHm1
c5Cs0Kkjfb9dF+DQovgAI+fJdHS50vUz+jlTLetvXw85EUsMm2QErMPuLO1wZnNS
oGbQ6xKAqkga0en/U7h0xtoa6/VN57mY2DtP5trYA03ViAPMfY0p7oR8oTaeNyZs
PD514MzNwBgoCH/sUh5pytxs/VEo2ZCQ+8MDOSuFPCAmEEKBOicbvKqlSgOCEOJB
GVPDuitSnO1pE27uDBK+jJPK6/u5EnLSoeYpMoya+gqznJC2e4vuyAJJPaQXJBIz
KZF4Sgksh16edQjLaxZWlxy9FzIXBz7kiMZ1Eb9S6bf1wD+qTf8cQ7wB7l9Usy/I
1iqINvnnttBfr+Sux0ye/ph2H0nOEvr9uPpvq7NI2drxUAlDSANuhebpWSG2G7uV
EHbHLlG9G/1mn4JRSYf47vD0ADGJDg48+Tp7bXjOApuV1ISQLQcOZJiKodlYCKK1
E1cKLHPBG+0AlvE/LDtP7c8BmQ33/JCT69+Uvukrp8mk77U8R7p4up3RNixHLT+A
QnpYZl43Lb4wtkv9+Cl4IX5A7ku2PyLntorUJ3HKPth8V0CZieHdIw1Z8Il+ArP/
+QQseXUnHDE3Kyl+wsKVLybLihAb3rCZtDMiRPB8QF8iocADqnyV1QoMy/kgM/Gp
sMPGwVsg6rgydmN5FSaSImpAuZSVVEFEXs0skqekdFnEXBkF2zxiUXSzW7Zo5qYs
fpCfpkDLuCsjVv+7AxKHZRxoeRylZpN27qkNCr3LKAUbBEzYRIOXNtZpnaxmesMV
k8sRrsA0VzT1WRuZNwvaZKmCM8WdI7CI1jzE8QM9gAQYD56ZJSYfSB4q45VrjVZo
1t/NMT3V11FEJwORPD4ZgOJ55UzU/Wag1EHfLrkYA26RuG0EpJQXX5GNDMXEqa9c
pvAxi3IhN3p/qApphz4RAxF1X4E6zUmyRv8vM+1GvmiUJc9g9HIdTYpUf7lTte1z
IBmx6XpAwBkdGRv/mPaYXYFbHZRDMlHJmoX69FYCQV9Z6L5I2+wp+IhmZgNaU1Th
3IBaTA1y55NYiWbDdEnZ0/aHNAfs4lpODwKbLtA0rjcL27TSegqiwLdFxDKlAkg5
DWl7bMobxPbxZSvxC4wp3joEuCxXEWEUSHLKzOwgGFMj2ZhT+vjsV7xwlWldgEos
5+sUDdzh24I5qx4ge/p+6HJfiH9jkYnAr3M57cz8cJZ1jArAdP8YAgjSZ7sDAvcb
aAUihQsIjuTpDFuuujI99LE2AuvcewEiV+i0YW5oqjIOiH6QwB/3KEMCdRj3G8Tz
A6tyUimZxW1m/4QQt1oXhSRM0EuuZfPK8RfLKxJf2MpXiDuLH5rj076+n936xls5
mohfQ5f2QKcRUGBs5O7g1VeefI/YeKE/KDxNiOEEATGLDna9KgqQysOF43oK2dHp
UqojXiPKGrmGKTUbJqugbmd77Op2fmeDG8uBfSXMkQ4GWL9ObJB8fFqDkKH8/+bG
/eAafyLBO3SFmySoE9oODr0OTHPPq4SuqnhH7MC7quthAcS08HJVuVYQOOGjvjSu
ww2ByBZg7eaAp8NmNR0CSgfsTsTeCNVTYXTpF2dy/1s3g7i0WDWn9lZY9qUpHLJe
rkNgXc23YqbN5QpkAAhiuI6fFI2J0QtGCBRPGKKaUk8JSmllbPqJ4t6Y459i2EHJ
imKYLscPjsW0vpykuL+xrk9ehL0Jbfw53Wtmw4IrLbJMjomMjhttcetvCERuwKRn
6gT/GPN/kko3Q7VlQ+vTr6s9JuOjBSNc8JWHyr8J5KejzG4scGTPLT4D3zbyUjL9
jrnAdpeZBvVZrwAT5sJNZXzqGEKWCiuZ+e+qIpgEG6/NvAs4WeQLQc392GYcK2vo
BH3agUh0Nc7H/n/j7Dx1JK+4mjZaB/WFG4y/nSVX7sm8/6WpdMTIkOsmnMtXjwuq
DCBIWZsMVg5brQV33EfR0SvugpnY2ccXysH5gmbeLcCz1R2KaFoUFMahfim4hAoN
uzVQ8IwwhPhYzJpcUeoPR704r4BraOF1xABs9UNE0l8atOa9fLrs3UN7qhqFfL5h
gZ6IXgzrqTa7q3boODZ4p0w03XwsYSUsr/nz1bhoaECMLWx6eXEDeXw/9Te/mh2Y
si5DPxS1MFj0GItkXvghhqg2KzCpPSrQUuweqh/VOtewgo+Q0C+AhlbZqOXoQ9UW
KmC+beYYrlCqXDCLGSLw9vwalNzKSV4P5NdfglgB7d+c3U+sjJlGTrPKiY88ZhNO
J0Ba3FIxnQvV058gtHlVw0CBRAh2lFvlT83WXhbl7fvLjt9JVV0LVU4rDKYiEY73
lsEffyaU18dc9jXTQwknYp0C4jcpHxHrUIEal8quJ6HxY1La1++MpD6VtE7sz/Hy
0Kgo/VE1PfTHrXNkDZ0qiei0rEgwfIVn2zuSvSA/HuXQDQ9gmghA64Fi/lD55sDK
x3SVeQqDXX/ynXESPHr48oeKEvy9QJ+YgxnV4MdIuhjIsg+IsHqxgoGsS6Khf9j8
MTdSYQeAqqToMljzucraswYdMOeRe22OQvil6fisKfu0HlPH392JHnhWw2Jmbvga
0FStgtrlIytEG0QePYkn92PDyMtmmxaPc3/jfjU5IULqY0DZF8gIGwBpPoI0+m/S
G4oKrbyVCb48tPvEsifSbkEJGqNM2SRfCVaWT0Evtmq2EYRT1Lms0CJVB11AzxDR
55lgekRO/CcaqxBrq3HB5rd9s4GVaJd3f1kTvQpLEES2oxujhoxKFnTJHYiWldg0
RFKNVAxdU3ZbeK5/tAAxSDxCN2cX+vldZnYAHZOGQB1tpt0LGhqgdQyWv4pPsFO3
MvFen6MDRWvqkFikfvyLaQg6UZyWzchFXZ9CkpxgYHn5CuWYZt5qp+ER4aFWwT3o
qqWAC+/HREG2d81SorlG8vnvMvnLSKxAWCHaqV5vkUr5JhkLpRtXaE89+F//p8lU
29GpMXRRV1hUcyD6asmJnjxh1hrlxYY0SXu+QDaYeR/2qBoC6Uv2Lr/m0l8iQonD
855QZsErlOekm0tHplvATOKSGY2PWqT9voKTL+Gi4Nwtjb+zYLkhmR+LiZ8XLNfH
ShCjgz0KUCle0QM8sFqPg9x0nfnmpHooO9Ddyyl1M+hViMaiwmBPNFi4VKtg6m/8
eK/jTf59V6QR4v3VYGIFVjH7wJc2z2XLr7IoJPdyzjnboa1wEeCtgyGmj7GVlF3o
XDZZFmyw8EBVfYzDllaRe8HXa6ZQTVMJroXC8k6MCBS/iHw3s2cL7EPfC23SxgT9
41AWrbYrFXbGLyn5/A2GMcnQgRpeZib0RTnBr21a4c/77YdRDhBxNrchJmn5pge7
xsgkyAIwRrOSoydC7P31md0+TuYI3W3k7QsgpH5ZMOwdsrO1yMfxlPEveyTjfvAE
FAD0HYlwztAqnx9JukRah8WN2TfaZ8NHkL1In9snTXdD6lzJinoKQsGhSiLxy3q2
cAvULJSOUz3QhChjMiqDR3QbySi6KEc+fhbhciiLxdjMwBL/RZqmMt10sWthpuC4
k+IrNIwqtYIx7G0RE+EhUH+J+bTkTpH71HpMEgwZWHLtB/6ACN4OFIQm+U+9q7Zx
s2GIZJdtAVJaih1nRj+gBrnR5DNpKM9C9loWDM1F6UwqIfUTjeiEqDOpQgNqgDls
QGuimGiAoQ9ACHvzsqtkGnEbyaklpITcI1lUhcD6IGFyCHiFlUYwyr6ms5bLwebs
VSOTVXdXjd7dG32JRIiaHtkskb2R9veInkBtj7Ke3t63T8clpY6wQ9q4yhdX88HK
vrPAW8lu+duT90yAr9jDLdCTT4wxBiikEpLDquHkzY5bwI/h+DwCDg3FtiUbdxQW
nt84ieCgs0TGMOyHK/unvZexU3dI7x9qBi2XFlfyvyUTbwpp13U7MptHk2+R7OPU
TDfnNU/9Lt2+laTcVvtbRgZN+0b30f0hVfa4HSwy2MRiQTaSt7hbnuJrc/dHQ4cB
1SbCHrLAKoWiqIRdgTW4/eTrnOYkfP9BOjW5pT6tvLbj3ou9nyq5O9QdbCzqII4a
bkxKDBkckVyV8i5JXPMkrw7InUpUZlyaK6h8whh+N68gywXleXLgZnWrATZ/o+Jr
FW4VFabPNVDp46mM4Qxw0rdx3wMxqOQjG0CAe++5DJ2nRj3eXr25SQR81WffEJzk
zpYydU9cGSIesdfW1P1LqPzicHyMArtGmP1ZPhqiSEygrXsC2dymPNrHTerTHQBB
loHZL8Z6JBhSvz/hCehjdZizQDpHXdd9/BzXxTinOFe9MsHDpAYmGai5G4BRWGft
+oG1d5vNqjNq5P2iiTieYcfAzb9Vfi0mHKp4Ywvodi6ZE8ikx4rDosX5xSn4ScY9
eV93tuQTeVYhQk2V160XZOVhlBsZN4lznnSw0TTU94CnMRkFezk0eevAS1LfeCSW
sx7wJ6F8D5fO37dqKDMLkuT07H0CUC1+bKMumSEbm0SC4e8/v+bKLDKku2wiGKgb
3YNpp4UfhEYCvanx80CsJpDDR5sXuNshk6z33AyyonU8gZS+my19l6RxVsBOkfhz
ejg4bZZS1kuFhqf5wAbikr302v2KCZfTGFUuGShKAj919CMA3Zuk5P9e5pccZhRy
gB5CdWhytvs2ama3lg8BT78ZskCqlBYHepQ3hKy5bMCIqHUhpHpxsIgFx2qbw/FF
cDrb1Idxcsjp4rduv0U9iDvlSTCvGib3S/jOE5HgG4qQnqIen2f64hYFR1BRQEAP
KYcToh0n/sxYhEaIaGvqLcNzUUmUY0y6kDbYXMrsqjRR97g+I5mkwjpqGUBEwv8h
DVhaJWbN4Qpz2MTmikSwA++NRbiib329n7/1PdNpeHqSGsHZGC8+KCTM7ug2BYSS
MuAETQK+qKdY1Gh/Kivjg0j1auR77aDstWZCWOMeclSupzXh/ytQz38mySGIfL1m
z+GlK/6P0+FrOuhNfmMIrXCItxsW/r1EAbW9hrrAtZ2hAKksjfuB6DW0bLYLK1HP
uzpjXh7pGmYA2H0iA5eXIGwuqADUPIShBF7/xsesmEkTytxcre18KvNSpv2f7q01
Ko3Aub85RzjGFdqUpQbwWUf+EO7qtvmBAsdGSp/zTIAY6EsBU9on+bRnpplaJgC+
Qp6vfos2T9SJwkDjM09czqA3079CEv+GRl/t2/9XQyxXXwzi8xbubugq5c0XVtTa
dHoH4sgjG4lXl2yHcg+lrRRW+A0F3ExhBCComqJgGaka/v9gG8IURpTGSM2oROe+
7kQ8jbNncCu/isJ5N7lSpwuEXN6vhCaFg5i7Ja2Fp/uBTzadX3g6VYiDMA2p9v/d
uys6wKR+dHi7G1kWCPJQnSGBdboRvTi6HXPqEaW0yTKkKO62z+ixA60bQWso1NRr
IlupICDpBPYKnf+2ag8RYhNQWDMDQ42ndGcaiE3AER5wNqZCNxfclewasIvWcrFX
ul2NBbVKNyx+RxQwMg4XbR9uqkxc/XdS/4GE5d2OpCaKTyZ5GjTa8AheNe6OQk5H
33SusZhgWCqFzNHTSh8VH9w7KgK7zcYmGA6CMF8Cg0PyNrRDkERdCb4p00FVZew2
EHDiKPb68ocawGTJNEB59RdtcIAsTGcRbLOFy1ARgyj0tXq+TGpJ9OIRjoxokdHA
RzJORo71kcaZ7s4OEBTHwHwgNl5xbANCjk1/f8XUXDnEIu6YUqhxycX0ucQ8wELP
ArYPIXZ1bovEntJQpdtudxeny/dumAKD+5xrTReW++nJXqEoHmZMtsiy5xyA5Pck
+z2CzQ7qyFhoCTR4YKdwLR7csuo8/jSOIhnCvwFnOHg+chpxzOM9TAc4tcWfNRML
buodE7H27vEljd5QiTipzlCs+6KcYVko6viybtqpzlbWSxi03bNnjNVel+6ZXqCo
iJ9KnOrbP9INUo5rnnTGCqdlrZj6ueDESNot4+TQSsaXGYwivu0arLi3xTI6gcQ1
a8RK/INEYa36dBQo6c5F4uhFgHbM5yRY6jW8cb01yUUBUwrvMMm0Vjd1F/vH7efo
2zBeXjzjBPYW2dKoJ5Y6g/+47v5EE70xDPNSkO0Gm2fXPZon4zz1Tw76nc+Lu0mo
5f4UU5hQPonzWgAk/pfjivRwQL2Da4lftWH+NcX8fwgF9nsayL8boxGA9zRSlHA+
NtkjQ2s29u2TeQvftSlthyj7cW8quILI1i+mSR1UJVyfVTU0n6K6GTg2GxMsiP+Y
lMC8uVzFpL0CBOCLA7aDJn+vXaIjdvjLaAYJgyzkyuIw3dxA9iPIh3gQjs4UAThL
Tu4t3gBb5EB+o3ohNOBwXJOxh0l+ADF0qsMR6C8ffCQAOrZxHbWobOdVuDeUenfV
DD7fvkzNIPQ2qtQcQZvxa3NlFIXwpZj0sOneZY+SSxUozBSJk/LJ1g3LeAkKuX5v
IQina5X6RPFWE0hKdBZyDwzWqbi9N215e5gbrqcg2ZUCKYyyys6p0R7K7W8nz/vx
znPV9DNiJxilVmOdTPQIFTFEZrcuTYzeKChzHE9ZWsCdKkGuBqK4Q0G9O3gcpNFm
A5tER/bGgwm5Q5M6a8fZ0HEYDmCNhksJI+/EdLZ1rRBPX6CBi6QBgCwaCLSzOchk
2OtVpG7OhrnvVUr9gvyD3zsxEpyCVrX4vQhNataldIpDdqOpZS8hGhu1hiWqV1wv
/fswrhL/Fdn0h9zv0rqgebjN1CbH3wZRnNmgFcYMBcH8spGpit1I4/oFnodyLMbw
NY1WDhxvAH4iMaqpaz/OpuB/2YShz8RSt5KU/5jVO6V17T4HmmlUudQeY0UsPpwV
eVhDf+Hp9dL1M6noGbYbZCd+jh22zW3wlvYAcXYsEjbqPgQVdh6o/8NzV7Qsmy4x
FSVijHd0SOtW7idNr1oJjvcBRf1prlFjiJfLjJ7SZcx9GFyllv5xr2GHeScZENI9
gBWfqpFHjOo1RWS1D3XHrrEd844/ceETzVle7GRrn5Xn0Aj1DNGy8O9KtnhMrS68
c7MvHCuAuUaCWFR3TwPvYRZhYF16lLDPweKiVY4F2xCfTz/tZkI4o9ZWy3mKCP9D
cCfBjHnRcDfrlfcA6zs56CoHg3RVtMrItzdXRZbTRJEdG/OeGFPDF+Fy/9srvmKU
60rSCkQdQnQDxTn4d6ANFNBq5eUV/+QhKWueKq3OhzGB6HRPbsE/oKRijdCxhELo
mNSbc++s8XaYYSYI3LXr6vpYAOnfqEulGFzm68INPGY2C87krmyseDfsAApFEjAN
tHtENJV8iL75DUWLbRYOVNiR0dr3DyHIIDoCZ3ITfj/IgAaxywSzdW701SQXKeIR
e5FCcqVyOVem8VgZUrA94A7d4+kDUg0qprH9lUcxMaHDZdArIREkl+b21miRHaLD
L33OL6zIyVjNKNIXRSxvou7fimagPBS0d7UerM9aY8xT1nGhdW5O3yoL96tM2kOv
1Ls1p/BDhtilN8LzgofSr9iPbaQ/FYc+JHiwchgADiE7FQt+09YBtLoLsQh1jONB
jHRVScnKDVlBfw/8toZ6gLgDFEpY5QWQiHgT2jbMay+5SctrW6T3gKPZfKVzB/hr
Yiyt4ozi6IJELS3CYb+oASWqTCFEY5LXxhDLbL3yiYqQUaezLjDqKDH8V8E3IBTh
hXRjIhQAc1WS8tOkyzfWOuF/z/8HuF84nK4/6D6Ag8c/t9nOZRuSxBZ6GOFgEpqi
Wt9Zu+p0vKkZm1Wb4ZldzD/o8HygMyCNLjUzCcjBaGrjb+8fFB+1sSUPHBN0rbck
h+STzBRaUwAVnU1woGuJsMzvpoYXFcokPjjLPBUZPPID7HgacleCfq9tDaC6nFzi
YsCEPUvIvC3UoDMvm6PgSNgg9cwxWSuhwNMpd4rVHyvWQjCE1FrWsfRVi57JZKT3
hQyjjM1pcMofRtEnS++zXaBldpv74jmepHR9PK0PiojyaZFZ1hR6E/XEY/dPnzUZ
5YMzgcpmgiSoou7xj6JtQJ0nPZfd8hIbzXObREZpSf7DYc13S4Xuz3NVww1eIRto
AzjY/sbkx4lPP364XW9sseWn33lHwKYEcqLJHu+IEnEvz2Ydc4uzq/S/MlSBl/wZ
ixlrvcODVnZIOaMpYBTQ4YPr3s1pWyfnAvbVZRhMfcF+7cCvnvGpvQMtWR/NIJZC
gCwX6HrPAGjOMkse22fOnbtWYupNVOvOjt3NsdrCBpTHZPXy9hmrumqe95qymAsC
diQ80gae8k+OY4DgoO1SLG1OFZ2P9aP56yVZDMQ9PQfUkZfcXm+XsrMia0QM9ZwA
7kBMW+2AH6hDLgu2m4svrxFpCnVR4nF6HpR3SwNVLxA4jaCpBba1y+C2beb3hGS7
xePtEpomvwUBOD+fr+xy/abcXd4EqNiJMI4DYRVt4OHeb8DpN/OdsYFiN8hWidu6
hztD3sedOt6kcB71pzowHIkdMOtSyDkdTDMUvFFOjf/WpAhogoMlZA93WCi8TRRV
ky9kFMBnzKQ3nRvzof8fCqWKuUR+wnHLkNNVSjzmJN8Ym/iko6jysZ2Mv0AoYve/
L0wXAdT/cSe33GuhKeGf3FpnRJQ99R3rgpHphpiaiwFYXjYPmqz2EueJeCFoZYzZ
qlG5mBAg7bWW4YCFlCOapZ49jqdWrWgvctMS/QJskPmXqCvKqFbEaMCKjI6aKf56
BBptSaxZXHNcaOWpDNZujgDouSo5CBBBVn5LtM14D3aNXwvzD6SOCLD+9Ug0+m7R
9ZHUmw1KL9LNk0/8IZ6P0NpGx0TdryULJIKkWLO2L7hiey5O6pVorVpdB5la6GcH
ZS+Mj42DQrl4ALERJqx75R/MVTyF6cZZMYZdVgfWeB9LV/DCR4ZneoLSpteOmGnK
nYqLCGX/x4UipCP3/no5YGJhZhMVqgK/vm9i9IMwNF71TcY7Ja+JDzJVgyTvL6LN
sw2Xpw9uRJkKxDZYuRDrxwqacdqHbObmlNm9K2Ox8yrXaHrffZyS1/pULBaO3zyW
PN/xfP2aTp3copYfsUy1WNJUAVTfNF9FA+I0km6Xows9u5Ql/sBQCDsyiwagBShg
iW5l1jwsCYAXGqSeYOREEYWBqoAXJBzGwVkweHT3j9p4GKGAUBQpz5fpGETdpMY7
1ksMbaTD/xYdDAybNNREfVSZFGc1+lAJg/xlywI7PWB14VuW4g7VtzAPFzDmoY2s
v8SXeRJoQlegjZWaa1PtuNpdpnKl6DtEi+FgA8pQXBs6tTV2ckMFCT1RvkvMeWoZ
G9jnt3AZSVypPHft4Cqh+UFRvpczKyy0L4+TrPvqbuo+nS0nKrv4ZgcmDfxd7GMI
pm3QT0EYKRGRnWwzA4uV8VDD9kPx4QL2qYRI+i7pwQDSxdZUEojbJpXlaxU4GceJ
0OBm4zkb4Ak+Y0Z12XOVtxlegl3tJmaByoZejH7phhHIfDBHHlax440yn3uqXiaz
0YwHJEz90a+h4EMRuSPH/AtBsyc80srg2BkM8xShfnjUxosw/hF9sL1Cs4BiH1rw
YJnCou/r5FUSog7sQpBMEH1H9ABtsslDVrItGnSgg8iAXp2sOnP506yqd/YE8GzS
WzaNTt38nIO9seDNV/ymePRiEV0LSnWhPsw8zZ+dwlP1aBmDd2vF4etL6famI115
iM2XaGgnt+NeQQSWamLZ0Fv/503tNn3yLpHf5xpJ5rDplLfSiLx0qn5eIoxO/0E1
tsuR4gJmCRJhH9pOU5GJn+BTwiVaYQVKTC7PjjSkkc89B7oadODGSfj1QMi4nw5C
uXItJtkMNhSXyWQWKT53sMhHtTsTL9j6DmKSw5Om6I+HJkorLn3rZu3+89hXn6+B
kSwRviSoq2vqrYr2j1m8EqxxzeJJ1ochrhURu9t4wVxfbDGn5k4f4Fc/fHJEFhcd
4+M48tj4MtRx4m7PJlSn359Q+r9CUmzZpnpJyxujob4aEnN4Pqe/Dw2qDd1snRm3
m9NdhRXyLCqzwDixpQYrMDSt7C1aTmyuJxmwhB15jMAJDhZLzG/i+Li6WPncKrnY
GyQxcZTZ81S1tcDc6ODDvthBfWuSoZS35Kw/y4ez6ororwOJgL7PUn4RfIAuuG5A
N5+5VhAc5MeL4I/ajdG3Ob0L6Eh2SZI8iHKuJ4y8BIW4ko/gGECuCrkdqdSLLAN9
gqoSJXlTT3Mc4E98J7PZU5idu8RqpTp5ALIe7JBf5XaQXuxLlxyvQ8NbD8Tlzu7b
ZzK/9OUUF7s5yXRMgmDt5VRBwEXLgWApqtwnxjHVxJRzx124cec8qpjpXcOWx1g+
GoN+25kC2Uiec4q9fM49MuzxHgoe65f37LJFVUsvb5wAoDx3Fj2qdV0rbsYAYrFm
aKO2HSZ6ES79RqG2yHqIz7k3dVQrwXB68eheqOkLpkVmtyH8ssoHI0xYUoAlwW/O
YrrKy1oI12Y5lMAZ/Wrcfv6u7Kzu3my0nl9QdFZSSmy6Yw5IfwMoUE8WeLg3tauk
k62Uy9T0vn/8Zwdlv9acHXaz/ftFsymswLHup2Vq85muezojDOUyYqaZnesUYE6M
/AcQDruVB7IDwx+wumjs42KP35Wpto+pig4oFKeFDqeukzr4yN4k0nuV2ua4Hbvg
bvwkxXtIl0aFK6XXoc3n3wkhC2ZRoDW88e/VGBFVVDdLleqO44dj0Pdy8o9f/nDV
gQ99DHhX4RTUcZywAQO8mSXtkIMJmk21LomX34btyPldhgGkLBpI0bTPun/eSw1n
Y7BcrYk2NwW7Z94KQa604lQG7DWfzR2IXha9wCU0h9gSoT3uE4txZXnj3gn8yN6U
JoOdmWPT16wh+m99AfEzMUw3HzOUtn9rH8X2EJwUh5NssepgvrWcMGz9Ggp7QI3v
lplxaVIUYr6lQxUadNwrIG3sN2VOr1OO7SX8zDY7wOGWlhmuRqgXfy+pf2rYLG00
7v0Uk7R88os30mnTYVHbUV359RPwftoGkdcufc6ayn01a+yX4MDDs7nzpCJthsgV
jjpSupI5ILtLKb7aIuSewT3dXkeNOCSZzMSbI7Q9KcMORV64Nx5XKTgr9Z2o9hT/
QxSpqQnO41UsXgeUUE6Oh/D7uzesO0lICjvwMh6csaMm5tW/Mp1NB99zJ67ihqbw
Irvbte9kj5Y6GpNlXOmNNuMqc+nGOwxo14cMVoltXB0RrhzUju/kc/6r8dwVX8I5
l60Cy03R8dPAz0ScAYyDdlQ7ExXhYkRiOmCxwmjwQqpS3JoHA4C3dzsm3XpUC4+y
nqH84lykYbQxRKno7b78RVFfVlOTLQaX/WRIqWGaHNmTB0Ac616xQn/H274F2i3U
UOLh9RGOA0hpYf+e0wzKItxCMrf73f85CeDKpwCxr2AeyIKFll0oAiOJ2/qaY1tQ
xTiI2qNpl/iuLRdYdCFocqSARzjPPdTULiuu2v/eaaNVaGovZma2dwTLYaJxBrqH
OFvcmosHxp3wqdv0NsouxxWWhkD+jIsqMII3hG0NgC6dl3iBl5Yhz86gN+LvKEt3
+TCP+FgL0AtnSjG4wso9SVnvWrR4Wt5MUNNUCjane9+5X7TYh2WnFICFYhg6dLvZ
jVBBO8Ov0rKa9k4YrfxMDF7iPD1kWglcDtQs0RCtyJWu8HlbXFFk+N97WqVhX+Rj
+btcriHB1+xkhJunYeO1DOtGcWThzpnmyq4c1U7frr6W5BFOpzIKX4tYC/QRPbfS
MFHUBcZrU9znxQDfhJ9fQFtxQbmFHGmCL//P6OS8TNCW6Vz7GTk+SY2wCnc5vLmU
SEbbHbPFTRspQapfEn9z/pMwZxL0i9uVzYNlyEu9sdGcY/Ue9K/lZbvXZbOHmjLp
v4fh+q1Fx19PbWkJJmP+9nt4H+ZfVVVFURwIOyysRba9pQmUc4WupusmMy1OO9q/
rdEDA5HdmBF2CqM/9veLvteNgrog1ASlClPrOo13iXeDzlnZ4Vm3KXR1UDfvbHm2
SXTmDUmE/iOOIBCBKK5DsLBYvDwvRhZJL8oLfyKSqDvY7FRE13uI0h5cjAgWOqGs
vFcJ7PkcCDtbJCcKhge/uu4rqth8WhoOOGWUFGuh6+GnTZ3XO+Dvc2y9RGuliLXb
dHUymTBHavTTxtGnc39ptLLe4O5Otg1DWBGrkm3KQRSkh/wp2KXK4GVAbVc1iT12
3FnvzGZEwMRWUtj42ZsEox7c4GWNNnqmT8GG3YmTbsbqbop3zittI+OF4A7+Bf0p
f7GW/UjYTyoVUsBHGvj7wXx8zoxizs3FzDUtlvzSU/rvPkwKDyy+9Ut02OVy3RzJ
9yxNdZtVyFc5e2MBujZnht2pYYcES37DyV6QEhzEAKHdy3Hj/Vbxmw4uFuv6dJpy
fUH/7qNLs15BqpJgCa9qWZtHXRW1JMlTeiZ5xZ7H7tdC2l8MaoGIJJj7j9pOlqtE
+OgE2VjYant6F90Tg3R0gpgUaw0wkeT9+63ltvbhskAR52dQnrphKgUaQHIvQIwq
49I3/9N7BHE/bfeN3XiBOT8J3SOgEfvN2IsUPSlL9eXDq4/ZMeOnE5FQjQU3NTcd
OM4KWlyICbcH/OHsr4hMJ7OmWVILYkV7Par3Rm9fGuiSBQeHN6VQqXLQ7d37uF3Y
i3a/sueVrCUhblwOlAED9eRXYBof9QJi4W4DiUEr5CZy2f1Arw360uJYdZ4G/I58
Qz7nbbroSg1cQDVKc7XnyaIiqtYrJltGyLq9GI9hVLHy3yyi7IYGAkUugcc96Hkn
+sAd7zI6K9eg72s3ZRs+VkcYy0aFi7pGSf0ySQZ0aQkgXqYzZlO74ojqDGqsnKXt
mPdc7/6PTmQljfeiqvrEqYUJMU4daQZTezRc3aj9gu59DN7XqNpCSFym96iq83go
3fX54sQkJrU0Cl81idXZ7CEfwjnkx1vSN+EQ0yAYU72oVHSdwO5jmdP8NLl9uKNa
58ITh/LxPZhttI4XnqaGlA==
`pragma protect end_protected
