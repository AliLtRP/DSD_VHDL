// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
nOX5kUEkLYSqQKACNeOeBKxTB5iH3+8pKVSRBi+jSSltzPEx/nszg2WGQ+xx9Vf2IISQiuv6/RgC
Svkgkjr0jb0KP5/d9h8fFDJyp1tvn4oTNYBialBEOwLwPx1cAKUU7bnttWAAQnNFvqzN+Ax2OD2X
AaEI0cjC+VMw8qoY+z6Ls94WyHeLJK2do68C34NpOBk8GFg1spsuxXvIYCagkVVaM1RirM52lzwX
c1ekdd0oK7ITfP4Irjv7eoeTUZnjaK7k6zzGPjtBAQA1VTLFMcIP/0jYgp9scM3Vwzv7t6Qn00ll
YXz9Wo6bG8O2KyX8FO4TEdPV9H9mD0aDQlTkFQ==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
4mbOqMHVpJk2EwidoZLsDXgdTiGz0TIwB7fn1Or3RErkCKBggmRNVOf/vxw3WtuTsCUptuZOTvem
SwNVk2qeM2wO9wQk8sRG1HQeOl2czpxcyiFkO/P/xL1dJ/vAYurA5zMNA3jgfmMruP1+tEMshHlB
z+r8ivII8JBBJKf5+rdAfqepWlca8YSIljAJNvbnK3Xe0tTM6L33BHppcOyRg7H2OWeezqjgdhBx
ABbWkd2amFy6VpCM4OS1zYFW2r7A4mobjcqQXlRpQq3UdR5HbkLKkcyvt0w3p+rTJP7TwMTA0Dsj
LKoP3neYStkc8GkMcLmZA+gbJ2dT37+4pZwWF8unU/J64PRt+4x8jaPwwn2DFYdciCoq7NvieuF6
9OlBzh25UQr8Mt1iguf1RSVbC0bED8qRAuDOd9BhByC2mKEuxlvrQKaHtPBIvEpJeKLG60hz6e8y
exLZTHWr06AGhMzLw+zYCxa5k+FcErA5+b0HPib7OWuPZt6u9/IYVCRk8CAkvT3LtIoJJm2BpgnJ
6m+DG5UC4tDiW8YroizdOxtgDRi3+h8NadvFKqoKfpSowfgDMnpV41n3qqp7wA/mVA2jczsMaFYF
FUbrWDQJGfTNRKfom2PwLVWLtzZ896EunS8fV4Gzmq0+gsN0zFuoFVffyznBQYqCgJPKixACQdin
oODr4AmUekzsSDops3zIPPz3mkPN29RRb9r9OcjQM1qYzZLodjw6W7B5ZwaxybvTg7pP1xRIwO5P
2K3UN5YFicFuljwn9iOQsEbV4GYteoumilKd8SqqbnaNfONZwljV8PnQcyBc9mG5SbIyI7HvI0Q7
T4oAqVJVl6nkqUshUL/5SLKf+0H/EOrKNrRHpz5cSvLD/9yqBsPclv9RTBD1jxaM5tvM/a5HoVbE
1UQTtzbpBONa1p0eoWv+mrUud5J716b5a6flh3eoZR2VKwimIL2d3oH86bpmMs5bJL8DYTiTmfB0
tiJ1wNJeW7XV1Nnq78Q65rUVIjke3W4bYapgAeTVJjrMdQhRWYf7hxNxhtvluJZHjsg5YIN8UQhd
8v2MdcazkgwOOLkBOdilzf2e9WJLKWaBR0vD4BLELMooLTp8QJwG5xmYDBadGEL502iQsnoGp34z
SwksOrAGKy15tLTQd8s/a9HmBQHEZsYNcnNrGyIlgUXUZZfF1uW+S+lJkQNdY/plO48vsRQVOazC
YQQB8hyEobjxRNxy84Iq6fMp6iA2Q2FWHjftmRUIWydDn/dIQckGm0QWdWnlHINOb+rh/l2ryxAi
9SXIqjLUFedVwM1g7o8hskVlZaD9qq48iIa9/a+ZLjfxNbD0TcZWstt85J63CIHm4iMbOIC19evH
GjZ8gcx0/8u7LGms2eu78F1D6MlwhGLt6UaU5fgx5TcgsfAu7G+yUOO8twRQyaj+E+QuqTAXefA4
yOHKA9WsLUpQ1nLpUTUnxCr9v0g53q/0hLcEx7Mg0lnTYm46C7oJFJEDoZOuFRwBi05F+uRI3CEv
50GLv6MiAAz67EUs5lL3dMqZ87EZrprRXMz7B/vA6eTfpVG/kW3JL1GUd/e+3X3xQJch/jiqiodt
biKz3AhHMJuwGXEql7ic+Lv3/9Ax2hsDAOYH2AFg9TkXejcXqr7c2q3V4ucILihlQ7yuR6K+L1tY
O5jy6DquXg1g1OhbS0HS9lcAQed3riamxFddhjml1WTbNdUD+4pG5+KJbjHVYKSSOimilELt3lJ/
IPfpc8qL7/7upvO/aYJbrJPxk5CLWxYFhRItpZ8Fs2X4uvb14mWeHw79GQZlyKUNy+u1HuS26ixC
zUUN6R6VMzcjjIwo09+XzADQX4/IoIvLhFOJ2myXBr+6NoT9zCrFjfmFNNgkzyvvrXww/ZV8VG6M
gk/gMeuBSotaqP6CDCkvYlm4fEnN7UPvt7u6fRtlN32Oa+FVGIIP5BAcT0zWFSyTM9jZS2r33HAW
zGKz61s5MmM9eEdLUwEJms1ezGutY1hJdnO7JJfEtg44e/kFi0yMLq6vg6zwU9KU1qNv76F5vnJ9
swOf2pS2c/Vk75G8d5lTZcKHYZBQ+/AjtKLcOi+vdaKKs0PAIpOQ5ZBE4QtQD6shyAbpNyljJ2NH
cjkNaQa+w7LjDy/uwcIQTGZBH/tcEt7v/AP3c9wSampN3csO5Wsy9c3bPGbpEDqq+4ETJZsugQoN
5UutqkGyu57968Wsdtc5wiOfHMpsYYB16LM1/LBWLTjINwTcxrEjip36dpT9dzZi8PqETehDNJFT
I8WeS/zEhlHTnurq8aWgnBXdcGRSZy5QqXN54cZjTKvY/accaZIU5vTBV+qJ49Rnx6rOiE58OiPt
vC3Vz8lEIC45kT7R/gcxImKTC2Oz9XLfDJshWp4SYxpr/8aJGCJmVF2h/LN7y1oc5T6Dum2PbPYg
KEblHyeo/hoSNNEug7SD2T1ZRUJG1wc+NPYejL++/vKpnHE2xaX0oYWhsubDX0MQMl4/78mCJa0H
J4IbAXlBD3LpoCDj2Qachmi/BHBCt3ZE4Bo8Q4RxMdZ9p46a9AyWrKNa3zswyKJ5XQgsjRNSMAMV
IBWjMuVYLO0xOfKXnltqUGRGwlhbZZ4EXdtRd7DcMANvVFKX4JPPuX/ZiqDNLqXrzizV9YzEGMWt
FSW8f7tAhiZuo0HCc9belwDcUoLUtZDa8HOckDGwy7+OO8sFC7tsekalHSm6ZosLkdYMvnBK/0As
yB2w0IFZpkI1kVIH5Tf6igxANk54mTSGRMFqdeYF41yE4Ztwa+rDAmcFRDdSy47JHh/5JDbb7217
2gWkFDPKaqUyFYYzGYPgpPwtFMzpzEGDiGva9sPg16IcG5jZDnmI5bGN1WIxOzJ+KTJGb9siDMDd
b8iCT6pKF9+CAteevhJnm4SjxPkvQENKd7ECTucbAk02upIv7bo/N3NZu6vk1op5oU9NorTaCfAf
TIpYgc3Yk29ZI1dQvb61tWYry40p5Lh/uB1qeT/jNreiItY8GUdwsYUxqNZcyJltbzqqH1U4noYO
MGWONvTtDNPzXSzbOrB8DybrzdxSPxFSG/8dCN4bPorgjFuff17nX8q6N8Iy3ih25/WH+x5XB1jb
8se2gH1uyXKfgrxiuU7j4yimXzrMEVjbYtqo3pEohrxQDqSTc4IlWdpZ6TsYsUhIZ7SfA/v78qkI
ws3m3sNW3iRdYOE2wIjKS2SS1st9/sjuaNM6QoDF/f4PGN3ZJU4HYgbw3oVfJ6eQrOWIrEL9Zd7b
xCxS5CsVb6C0Rpul4LIVJOLLhJMTLti+WljPpX8BlknS2qBIq92KBzrRCVQ8ujeNSyjqi7IhpPG9
0wFSoctbMuII+TtzuhcUMSCwK+TmqazX3uzH5nzsBdxbEnU86AD7lIheS4i8u9QL76kS5FG3WXs5
ls1HGrsw2XRami88meJ/BjybKkLwW4wh7zpNMZoqpSUQ0nmik/ULgrUdZM+L0mRJEdVafmfHc9CD
uKfS7wFkpXgUBMOP3JvF3/dJvmA8jMb+hmZhHZoKI1VbjnHFWGn34uICa5DQpsXopK6VqyPaV/Yz
WrzvSQEdq6MdFQvApidA5dXTDjUHJW9Tib2AiLpjUl0KUAixR50a5VZBhR+Efq8FdiB2eyTtAJa3
SKWVq3ygfh8UyP9qaP6+lIE1J+eJbwvfIWf/f7Vd6lmzfoOOqBQyXes6yrK6LEZJmrpPqU7EB9US
WWv4GOGWkzGiIAPsjp4w0AvD3hHYbMLO2EF2wpkud4tRzfYXjDqBuQ84e5ejjPmbZ9bw5N15apBf
V8C+5t/U1JEvyBjB1eXS1F8EcGnE1ckdDF/2PQiV7Dg5jUoQn7fwqy1qzVgcYEA/0N059sm/Vbwp
Bzktn7Q1WbvT3yXUdGh34CyWAMiE325mAacQHcgswHO+/kuEdGgqUp2HKWyhpn21+6RkRgPZ7ins
Au79KCgdXRnpPE40+zcBfOZwxP7JbkrTOZvlunqonC2uCnr249GjQ0gXIlRBgcq6sBxl809f2jOZ
c5Q9wWd0DOYbvBSg19Y9eqxGsnP2Xh5ag+YGPEm6AjMw19250Ncr/ClUDTmH+Xu3TaczFVeEAE0+
osddfwuK1vIbylfpiKd1s78aXtXaLdTM5ICn4pFQbeaHrYOI0wCiAzQYgs6iL5JIQ2QtgGsvlxab
mS51uBRjT47V24DRNjn6OnUgs6HHn17M81viQcC42BvKPdnJmlNIKphm+EwSl/k6p/PAhspi0ezr
lLz9R/Y3fZh53+POC8W6jkbwf4monQCGA6XGY3J2PvkADSmUB2/E9dURrD8ONOgMHiZGhF3DVeR0
OzL4+F3yOgkB3iKh8qG2KBZQ5ZbHraw/GC+NyM+meqtv8YapMqGC32ab48y7NUTr1BXwvJbwpuls
AG2Rf7TCUEXJy+Ps8r48+pLfhG50wfGu3a1Gy680nfd4RiPkxp9TLHOoSeWwJWpxOz0ciuK8gu5k
LlIqxLfsNUpp3hPKQ1DRPeSv4+N8UgcobK//ZuG/L008IZlTlVPXEZG2o1y0MxWWVj6LKgSNPq3+
KmjpvqSKkG9u7ZsnPMTZ/mg7Gn35fDPHRW1eSWXTNyX2kuRZ+qSv977XBjLNpuhInPQMDLkcLKz7
47ZYn8GJsO6xzSRA5XQg25n62lqM5kVYKjyW5c5gDQYJrBvmGcPhLwayLglkteLS8doahkIsQ1r2
cAVImLvulICf2Uctj9krNRXYBr6sVn3HULKsP5SKUV+vixSBF8kf61AEj+jCDaTgXMvmtCQz9EQH
del/5V1ShFoefb/jfouoxg37DjYbqappen4TVozLMFjHThwIhhWzMGWNPg48kv646JLT6hh7X73D
JuFPInA7DUKqcrtKbZu9JZbMM+7DJYukIcgjQBDH0qU5BfDpqvASD7L4QZRLd66YffrM0Yq1ghFp
r2jcRQxOYgiTeMdKIwWiZvA6VmO9trx3lChzUWn7Mz9Z9Dml8I140Zm0VVGeG6lhxzXQYntE6oIe
3JYfQDLW94uZw7D+qD822GEgGwzqstVSgPHkqAUYuk+vIvGUOewpQ5g+wnCfi1DFsxcwRrzyzahI
1CDQL+9C2YX9MMqOO6vGa5JAuE6lYLI+v2r/lbAXHcV8DvG9vhRIAoNzWmk+IvRhztl8M26yXvw0
Gam8yqFP8+do4TLQkT4Cwrb1LN7kwwLxPcvra/PLFwbKm52GuXm0SccFMLS9DQ9YTzokznZYflrC
hNFVHqV9Oyd5Y8F8+4kAAlRWLZnMW7CdGeiXkdVMtzpxL8uxa4tEaynBYyb2e+3u0O5Fud9exEAn
WVlFXIDzLmMNKho0fbNNBWVTAOcsTcewcsQ4ahUg2N9YC4sJSwXXRP0mlPLbUMiXA2CtM4oSt0vy
5M69LQdbmPFgRzaXhnyjF/c+AV/2YllbgdcMJxemsGEqATHkQNF5Gbf3KEbyK3fSwS4u0G1mj8OK
hqdwBfvAbMcVpYKQK6bM74OWVghvTBAtKGFYSav/CQK1mj7G+bhg4nib0DAqm7XbuDfKSqp0ob74
jWXdByNGy2scJ9I27VMws6vKAbUD2GSfntxGg4o5cAbsLf+Nr2BdKkdOS5KPffkES70Ag8TqQrpt
Xrah2CEMKfEq39HLXuvl/1OOIqds12LUGglUHKxHzISNkR1pg3mS8gnihB6AfdXtUOrTIZUe9xNZ
UTWNd3iUH5ch08oJ/xIpQ6iavLVaoB1/hReto7ByVXN4GibIl0/kj6atgNaGptCINwr1MUp45/WE
FUmC775j0eeNd4RVTRKgdV8rJmwUFOckhsZXLcrXT8fBi4s+GtpwypSLHjBlY6oejcimiB1/LHFh
rKs9a2f6c9o5LSEgEx22kTrN/BrXi8+cu+kWNdL5hhsidM84Yy23eRL0j+lxF/OEcNKmjb9bMb3T
FKA1F3j+W6MLOfVNicu2JjLNH1n65hc8iY1N87IX3QXky6L+Kn51eAPkI48dlboFI3MnKKN5p6lb
qYK3bBoiJFlISbsAg+mift6bOyJu73WV1T3ToxNlMS2N48QaGR2jXDo+XkqcLiWDCiQT7iqCWrgc
05FZjSFfG3DRfVEyoQqgF25ebNMpkRUeB2HE5BPcHXp1M+UYZrKGcGxkoV6OKNwQUZvCpoKpobyA
CqD6ZDIKdiNeTg2YXtF8qmmmN7FpXL6P3T3t7ye/h8zdKnt/FpByC+t6fwVHmA/MbkiIl+6Iriu9
X/2/d0wYIaDG29aRP+xRkIKZ+yYZeo+RbWksmAUrvQAlNT06JAd4tGYxmDkz9nicusIaisFJ1619
H9K2Xr5gU6jC8DP6hTt49VtweOqbmGdBJFyD9goXVwmxKg1PGfqX85plzgr5XWmuIETsM5E7UuTV
fq/njTBkCplR6px/GDzGY/KvJYR9SkUdq4t8gkiUR+T2lKhi9hwECM1AyidZrWAkVRskybYI35Zf
yMIlvv15Bb++buY2Jv/5nA4YGagrb5e5wwbJJw9aOdoFY7MNvuU0kYDAysbv3vAxjbZ5GZXE6l9i
9cgVzIEUcEwWWiE2b600TaqZZAfjhNxy6XQE4xfPIMJVCUOQmHaWb5Kazmvd7eTmgYfaWKZgI9yj
ae8JA/fqba5wXBgrd7Ki1qKakUuR5zkHdGAxTAqfKECVQdDWmHkgtpmS312t7nnbFUL5JDvOmyA1
15KHbOet2xEe3+HL9rKmle9mbo2HndmcJKjQUz7sDVVvVh8L4YSMo+28LTBJ7MzxyswkKYJKMNNL
1GZsIzEwmSVzNF5qWJnZU1LNLpQvSuyB2slGpDtIk+/8Vj1YfNfhvkw3msHKFzPnKAKhiyPLGyT9
i/rG8+v+JhyJVtiDj/DRlY7XtxFLAzrqbo0RH+putLLvxogBQbnIJ0vsOuHi0rLxzztAZ/nj8NbJ
s3gvK5vNOspIc1jmcT4PmtQHrfyZGlfeAG9uDQdNAHR4q9GgkhPosX5y/CDj98sfB9PpucEByRsx
04jLasMyqC7iBdrNOVEU45tDyohslnfjn9o0/IB498qYjIhsL9GAvVJUp8bpVzbmJGR4qlNdb0uJ
q2uQHnol2mApUvGvjdqfmf+le/jH9KCFV/q+W1bmeLSYdey1cjBDRe00ogxqBwRcwZQT4Y0kVGMN
iw5q0+1kEws/6qMMzU7F5M0rGVGay3qIZ3tggnizoFcu9DfN4VcGGrAutCnk55aDClhLPYEwXvyo
ZBHB7jdslXFrvllNIF0dt+KLbiuY1GLS0UKUioBSoWs8Ty8wEeUsTcz8qWHN2orIBFyn9TDakQaw
9kLK0EvnoON2+yJJvW+8mdZK2gchuRWfvomccMXQ+JeOEv4c5rOlfbsjB1oqTifbfrTpagWqZBJe
/gx/IowGJkVbbK7VdVSVY1c28KzogJNzau8fk0G3Lu4m1BL172BnS8ihJLjMBaf7hskEIXK7u0So
uqL0rcE0zhDJK0j97dUsw7nX7C2A0bFzp0fB33S6nPw3qW3lRrDaUHTP1fGCtU13s1l5dBIaN4WD
dLWxDuk6Jm43uUdfXrC3CrWi7gfHM7C1xpzYl3bEiKjlNqV989GyusgDK3upbcqk/+344qCYsgN3
Rn1B3Al6PcRmL2B/wVW+nO+/Vis0Fr8cfak4+fYPN1oy/EADUU8i9m30NwbLbwbi7bqWWlUIbyR9
9aHztw1VYd7F7JZLf6PLihwPHUHOBn46oTFaKy2MIhu2qgoTozE1e8G8hEoF2SftQL++CsthNgP7
8/Wg7ZVu4TUcsz4t0E9xm1RXGZBhG+fhfXqWyRFJiF0VCDOfxdvs59eyHsy+R7lzMirqARECjjMe
GUQgSaOYRrFOZAyoV3Rj0eRFn4OKzDnsrvoOYadGg5saUlEnSHwJEy+jqlU12wHobcxWVez49NSD
wOHqQbN9wtghG3BtiScA12EUUDmxdvynlQVfNbdeAPsj2PElKlT5+bS4hlpsOwjGWyRipq7SBVE2
z9t8OcYDPKEFZoG3Xtr0ezMocDYWFUrlF2alHQtnneHhLuEQ0yn10XJmrnKFZziuJO3cKUy3pBEj
0tekSfwGA5CKLHEZE6Ii8xRFevzdm4/k/TtV4GBVXxgbR4t22B4kWFNcvB5EMEVwr03VWB5m+oID
66D9H2EPV13wBECyUaq8sqUn9qWm8TOdYGGLEDgAlJljhfXQp9cKfFR3mB8BG0NeAwEyZgq0LXZU
pQx2QAgcrs7JZ1VUCKJYdjmRK3st7+za/hV9Qa8bkT7Xwop19xj1Nebh+8Esuv0nI7C2wPkXz31S
pbIf8lW0NobLXR/W1FlCs8jaOrM6NA280ErVem+Czuqt2F8tpOiN+/80PRlGJRVMlA9IyQhMpxYu
D7d9uiQf8ppgrdXwdcKnEu7kVgdMFVZvglG7Yk6wSQ5HGUsg2WBgZCIA0IJoicniPgpDY/4iLK7S
zi7rBMua8IKdVUrVwk47AllMByv1UhNvnaIeclTayuW1TGBb7x8I3D0i1Z8oxx3CRu0MoayTs8Nf
60+q8I7pXLnM9BHn65bUmpeQDIZ/+jydYOXhIVPOLtEL3pXgh3J9c25WaIY7sAvZqbH6cN5RygYm
RUtcWHT7zfGAEg6Zrn5Q8pfvKYqULLnq/PC5BuVlVgiX3ed92siQ+LXAzv0duwjyRFonh7ZwNSpG
Wi+CHDqg942fKV5zNhrE8agAxrpubUKSOPVdt8eMIa+uvH3whUPenRw2s1QVv4DfMqD2ALUJ5/CX
fcDrZAQvU52c6zUNzqZGrj0TH5HTkmQ/Jh8oX4m8Hza75Wpq5FdQpUJyCD2Hb/zs5WaA/traaOgN
sXh7rzf2vuUVLFWpih/1ODO5Lqkyv9ky4+0Ck5GxZDu+vrnBPbCqWJLfNnTGFS46/+j00sLpFgJO
X5JB1wfD1FWwcXhtkkkfou/MBZkFk7XNVIsxfk/YaSQNHgBLcSbhZpQNrCDYP96SlDiY6C52x/mV
bCIFmbx/DxSYxt6z7ab9Pw5/aKEwmSDrDxwtDm3i06SwC98f4KU+K0iNshI8QeZJ6mdWi6s8sPnV
k4JDE5XPD4TzVKlheTluG+kFQqIG0soulc7m8+4bOfR3zF3bq2ktiInb+m4JJ6c5NJUJVF8CQ5u/
f6epZU0eUgO7If5jSm03IvJd2XSrBLwhPRcU6w7dit6ZRHAPYxZQDV7KeFs/0dweigi6tHECwU3H
yvdpQ/Kht1yObSLWf7SuM/XywNe1dIntoIZc56fYDz0ocFyb1E+7xgcrrDlz2qcFLhDkLth781Dq
LmYOkamtq5OZudxheYuwwdlB6XNJDP07TRaKh86S4oFxpEDUq7ZWihjveymH1xy8RKMns0ioU0Q3
935jot6dFgyRWKJBba8YZ3vm6pQkoHm/Kedrt4vGWz0cMoA+mKAzaPubMHH7dDLwwfmQF3GFHE5K
trhUUNLqgkVUn8cAaGFvKiuTslts39nq/nIYpSiqNnZ3PUM4JKS9o27KjKfQum+/XJQslCRKwC6P
mtQIiuWwy3ADo/6EHF7kEVeY+5z09KREfCiUvFniyjJUnExnClL3Zzd/L6h6L3sEfLou/cggZtNG
Vn2IJthK2obSGsUSuFtQaVT/xYLy8tKxSp2drFt5kJ+OqPwyIYQCZOg81wjSPo6T46/R4oYLUd6k
uIwTPUiMHcweCi0esbb9Jp/S3xtvi78/mlokWW4xqx4OZaRoO08m5eHmXltGuL7aCpKyP9FHH2dk
4T2XHI8hdt5x2ylzkxwsYC8llHYpMq50G3QFAedi5CHd7IIHbyPlzJS2wEo/rjt6X09RoRzW7AKc
oO+cWJh4CJ7MyQ8VZLzQQZJClXAOKktFWaaWQyaIV76x/EEioqcKdr8ci7q9R2KH4B26QokJ+aaW
WhS2Zo9Q7yCri7k6YHI4tLnveOhkJmzQEjh7+LG2ruZryOsQ0dbTVVS27Tzm8SeDpECmeMuv+CJi
hb4DQiBuZyP9qTZbMSvdfin0QjHm8kNuzLC0yEi8Q+HWBg0nrdJEJOk9m2M0oqGXko79wQzDjaXk
fTBJr6rlBg/zc6pk0MseHd40cexikveOgUxROLJK+WfXZJzs3IgHShryl4u+t2Ls8r4gh640XpzL
uUHEVephH1K8Bt5BgZrbFb2i9czy+Cz4IjdV3JSV/J0O6QXt+g8xhiXod80kQvKshgF5ms/dejDv
wwpKwQEWzjbmE9zBqj5QZ5fhu0LvE7ry2p7t7K2/PB2OwVxWfR8s8lc6EqYbAXELzJVwPtbvsB/A
xK+zk+vX//TOidSG+SLXzaa5ICWbyXL2hvAETaW/HIteJ4UAay8SQLqnua2lJOsEO7SFdyZ5CJ1D
XORtZHUnhe8CE4OY5gLD5JdgO2H6mKxEbo7sW7sPjZVSC5rizvLrzNmmC+/6ok3jIDPo6zXs8jA2
Ao53CqNmawYLv4GcOW7fhM7S38XVvdJYHyfkzn6dR2pVrRRyRoH+IGVj3DNzEwQIZV5HwqaR7IsN
MN4i0a5VkSRwNU7g3p7OgWZKY9geZsvI51+0Q0SYwSgEapzKp2ZHHLNuBvQeDU/8DdRQAJtu686z
DzuBSR35R/fa8H7Kx3kAYS5v7jFPtHy7NDtuEe1FpovG1B4RjiVj7z3+dAxTMZeJPg1okmrOHDZF
+2hFfBNVTAufNuD3W1JIhepaK6dwGi/iNvDXlInAP5UQ665e3v5RNyekTvvGZ0HSkYJuFzibpl5T
tUOCmCK3gZHXHLm7VHu8Sle8Rx2FbtP0cqFejxPKXQ3w1fnXfp7eybB2sdgCEuuK7zlb3OOK65oJ
mzSMVBMC6e0c1WgCrCAJ0r9MBWqJbl2hMjHqdpKBOtdecCcgi06humJBCf040oV6G8NaBI8/x88O
aDdlUGYUN7s0MhBS3R+4RofSez69Hb1XS8yoXe4XcgF/nQcvTmj4jXs020JCOk2eZ2EqXO3WLL+8
YENT952DMN/UdDZpKAiTfTm9cNnrP0SYdUBVMqky9PIEtP6byY3fMj7mpRN4ObZhuOuUQy/6lAfT
Ys7chyaPmLL2yjEsGSzjoeEk504Jg6T8lKs4U0Q2+RrdQojULBGwb0DFKEC5xLPuC+DzGF4Yw8AO
P4QO/32ly3M9QXDSELdRt+r/h1ePtmJYrP71uFaP6XYcALMf7/nzl+fhsVWqwUutcQd5VWTMCKaq
ieeeVVsWjPmWXxUOrwT5T7B02+i8MadMOaux/CWaKM4Borpy+nmAfu2NpQWbfOyC6x1C8FULpy86
XRiWwwBB3MmbT3UuXYH6zOop2xZ1JkhWhf5sApF1SLICd6RHhs6mDbBX0f6iXwCMUx0tNqM8hXjf
xYRN64AjsAPNy+4GzEPNcvumL5XHgzb534F815fTusqxK8Dg0stvku2GzjNTGIRoGn8xztDAMgvS
Z+42BwTnw7whe2SRLBj07F2lCy64z9zKsiZA/hEq3ozl3R530UYMQsvndhZO9giG2OUZwwKcTATo
RhIvJLx+cQa4RtxH5R20eTvkOUtVIG10JkzK9C271fkQphwPCJwTVGkVwSFWySov5KYYwgw+yRx3
eXl6mPmr41h79Smc6qHj9jtAnUxCMe5mAZkXP9ynF6FcwpE+fQ9p6knivLyXtqyhyxLpvSPawmQa
KaKRyKADaep3hfWcn8wJPjny75ubj+xnviNlj54Ty0G2cyppprBviVzYp7FsF7psw3X9Jte52QxH
VFi7Xnl1nU74xy+e052ZEcvJxPfS4VuJwGBdaUkGgLbgDFXDTVY4JrDAW5oo8HI7xUIR7mF724wp
cvc4KLikqycxTHyReiJ0gBmaDfD7fQ1Y+1nxsTmhbkYHh2ZbL0UqFsv0QhQ35Npak8wXFoaui2zN
9KhDK8VBKscj/hpWVxH/RYf9vPq0LLSTOaHzz5Nx+27i2TR0uDldCY++LRqspgijy48Tpt12xFnk
Zbm4UVYpNAnvFzbD3afuL0y92P534nAgeTJqZ9YGOOY8FNw7TpUb/Al9WibAdcMpolYwUWdPikFE
exGBzYXEqXg/p1c4SX1ensi6YtXOu9UVs2xDmqZmUu+NwZqBHQsyZc4txevI+YuIo7CcMUvvHVem
wiEoMXdh1jluZzGxZIFHHEkmukgnqUFVioBdiHIIOdbv8W2bYloNmb6n11qx4yJwO+gcjELOfxTA
pma+MXDWgmqJ2Wn/KJK1Fou9ipxi3KH4ohpitK9qgLbT+CfSn7oppxuNDlFTauntxOWQ6ywSWwWX
Lf+HNs6inXcY0/Kx2Bq1+YAaFiV3qMK+G1gvTUDu+gJlS/3Q/U9vzxEcGZB9WzmuijyI0rCXaExr
5EAj3IaCOF3lSoCADfjEBxl9BS9lJC0xGxQDy7WQtRJ/Qy9VFxnd5t2Hn4XO+iIDT6a9Bb+VmRtA
eq/oMs3s3LSaRo4cGEjHtWwGIowwO+tPzfPN3urzPaqBa0OhJaGcj9Q3Xml+PgPQp6L4lvjrYjw2
7irV199EsQDU9CpRbRf87LmHBo38mkAFGJa4wScYQnFfcb0wFMgE6YNOVEQ8Lh0sy+AlViYmLNgK
w3fjxi7scClt2TT/W1TsyzgRGXcJWGHJVinr3xYcTkTkzacId5lXdyjXllCvy284Wxt1vKUa0F9f
DBhdzOzsLYNnKdXWq8dcjEfdwO7B/9gEJB9ShCNiMi99N+q1iGgorQhOUfx3iEIC9oOnzgBhCkD/
lq3IOZDzqTmVY8tvWZ0QabRR/N3NTnfcX44tgmfXdNTrxtLDykh8LdX5r2ifRZD5DPYxuSgfj6mS
Skat1ob9mWUe7KHQZmgBWMngFIfmatLSoROwAqFIdqgyppPY3cfT4+E1zPas7v8NYOSox8ovyo33
iYJR7I7oOgyl95V44OqfWiLk7djuVSJFhzUKIGeksc9dE9l+En8bTRlKlSKeZ3bqs8LWHx3NAnlX
1xaJbpxSI74ADVqVkEBNfAjQXK+RqVnMYv2Spu5GHmY0qnlqeP++aGHHtsfh+flwkhMFy+X3DIiN
nyb9FG+yZoL7EdxcF0H9ifsTCIjL5Gz0HO80g8k7gR86u3Ks/NUTXPmbkz9TCc6+UbDmV3pKqVoj
V83lvg8fW93CIuy0QDhDPCiWDw/2eYufV24Zt5K7LttBmUQX0v1CA7OjsDW28/OTKL8SUcsS7yS4
nqAN6luGXo/NDwJYWnml2AS69Mcl/NDOT45qsY7OwX9kBDHqYGUPsAuLg/839/CoBxIGvMw9SEEq
TKfRAfTovStsSJC7aY+6SDjUr/m5mFu80wjYzwRZqNIfpWnIr6/KNwYRWQHIGpHRwnRPpYCm4C1U
7EiyaxMDDbc8BHMgwX+hArx/veAhtfW/U8Bd0R5YWlPM+3fhNSCKZlMDybA69p3OKWhf6ejemIPe
iv7rGLsQOAoVGXY8f9QdM3O+TaogxhPg9RJIWfoUVtaF5tL4Gpw+62dwcD6syq7xVHpuEOm3Usiy
nuss9yWmssrhLnXF9VUiOL4IS0ZDcN8nMi6YwdB38dcdxwNIHp90Kern8W4eMLJqfGcFlAAfpuxJ
3i80R9eFhmoh+F4ecV4D1J63ouzj+PYII3yjPfsHrOUIsKxDQzVTHoZ56fXzb07NDDXWARZ63gmw
Hzi54mZAFTi3DKDgYp7MWXRu1Rzn3pltNqqYlCk/jWch9gs3XoAV/vhL7/MmjhWPltAQyIv8buWy
Do+JTuhbiCd/T3HM2052lnOsOTXDh0d3YZGYTx7l0Lw5EuwGwlBeXNZML01KB4016RD4yj9JUg0A
lqypuNy201mpaQiS/MYRd10Y/JxsASuq+mcg1KfW8hxlOQB8RtL4gaKPlyNFLUFWDdp2flt6BDNd
nvwR9meZVn8zRbcvRRw9Ty7BhrD/niqwcLpQH49FDvqs335+LvttbG6yd9SUUHHOdn1mGa4TfWE7
NXMpkbktSfUvWXS6tTW8O09nfaX3ifGoPU7POhcu8FkQ1x1DPZ8+YF8mrsPTuMphvz3L/gRfFec0
ie0Q8U+PC8gPW3igwMOgenm7r/6SIw08oWr+rC/OX/HBrlKNSj1oIPcTsMK6PM7laRgS5oP5U8aI
7+W7RaTIzAYe+cMnpf+ekYl3Et3idWAQLyU7NByWO4eSCm/1MocMMFY0/A30l0AMS8Bxj4dVsb5I
QS+Ta5bXBQN7oGrZq75kThAFgsAnRBMg1fFk2SIIIBXVmy7sRYbmc8sh5qHb/i2pvNHTAPNO5T99
y+VNCVy7qRN80gOkmjKyBXd3YgcIt9IO8AXlavcbxA7dECgCwhORlVuPwrcDK79tyH8bXS0d1K4r
DW57bqu9o/g13h1Enw2+JEtcawpkPnHI1aDfX/oqWCW8zzlstVVhgiJYqUVB62WSQcSOgUQQQunM
8WcYZRjdQNmvce6QS6qHLh0H+v037eoFFMd/MSWpSwCkOpdCaEyI+06oOsHK0aB7ZB0o3Zl4w1on
zxXrS67FQlPpIWTZ0O+0bbLC12fi+e++lUX2hjrnUDMKD5GYs3uoIAzZnY3JFhuMR51FaFXdk4Dx
/BCbG9pqMynHsAiIwBJhJ50m5zWgbrVB1lgFKc7T3Vd2WzxAJkLZvRsodip0qGYmo0Fxz+kVy8u0
IJIZMYsTofp+nGf1Kb8aPt//ZEIp2/4+SCeUfxA5B3sPPvOpG0Y1Bmhc4UIMX2LEeE2LpmYLrlgp
rlti7eXzB+yf5FbdRNKROEeWOCs9aCCBLgiMDVUHCS49Y48QXV8Bl8yc1nP/6JDhquohxTj9i4Bu
YNiIitXqoT33o7HhYFAUCaggjUP1wBV9QDpdHklurcfku5HVVi/RbRKh1C6LKOHa/FqK4kjDAJl4
YBU4M2z7C/ykJatOmMzQWbZwRnjFrpjz93PIW0GuvNAlU5wb9Qes8ORUku5Rla6Ubfhp6k+Lob3X
1IxfLOGczaz1jITTXHcxou8hOP64UBkOsKfSAqDXMC15bqHMJ8UMIxQYe1Ng1zV8hzvNmxhRQ9sV
FGI3/1Zs3kEgq7Y4qi9QhAoKkHXh93hL+eu/EsJEk+hf76+Vdk+A1xvmRSKioruHlE46NszIxVuA
TDAGA9OJnvminfgij2wmkGiRHORWZoIlUJrTbbkuVPVfRp/QHbOOI2AGpfbxYiWV8AeMHvdMggzw
nvEuG3dkOC8uMztdFrhPxbhcA9SVB0BfjjeQOwrc7S6TMQVJi5HsA8o9HrI6ryoZ5C6YvRySozwx
+CSL42iKSqhhX2tYhz9SC2w6r78cgODmH6jJ8VWoO1AJxdf5aoV6JIFYJh5ZW4m1K7LZSfYv/YLN
65zzc3OIKFjT7uC4vlSBwdyHs+TUYrvNldj7TnUfS5lt5rFquoZGCzBpR7TRAt7p3NANCbrI9Dbp
P4s9+Os5FYJ66NVua0eOTeAL1DvsSinMbU9MoOaRdceG4MnEISKBGUd0yoPpG4vKizulEMzbqRLo
XW9WW6YhvkeKq26NkvZ46RTER07IXMPbfUNrtUZLUZTST0kED4XQ+V19xHAX8RYZIBoWMvL1+Zjy
UU9MCDRjfPrYAkKOWRxQrMu5Vc3kUmUVMctbtgeV1X20SURXXSX4GJQWxtEfEGp31kMqSJH6BRPh
jwbsKzN54zyNNbDzmqCIek9swzn/zXNhye1gp5lbxvtlOY1llN/Fhml2RVjBt1V5X4HpGJT8jlAs
mIeAMO3UtGScgsNoZWfdpPRRFD0ZWfmjIK1/+ZNlnaelAZAyKxOrzERcG2JX3kbzK6+ip186o1Tu
D3jELZ/ZVdRGcKtrvkqiztbPDi440I0KStnbzTAoSkdT3648wUkFUTmv1dUSHO25SD7EgchO71l4
t2iCAAS01qcEtTmkyLuANqaLy30jyViCk/MoCtv2yv8Gbz22TiuiEUhd1vV9un+KieIdLJfqPFfe
bW6jntz9Yf6F0HiIJ5a5/g/Z/8JC7I8CB3XkmIqXGPN+vppSFgQ+TsipfFofkVjWyJGw/gLBSC3m
pFKiQYvT3E2W3M4WZWk0+UnYOanYQB4kpR8bj7E7dvJcmmpSxahtm9G2t90JIr4NIcEZ1p/Xuo9I
+0RCKZGF4/ZtorVm2v33BGE5ryNmCWYgXV4XmlqqNvUkSJuxORxcW0yJNw+z9lVorj3+xJw+N1V4
aJVQNwqsYr/ObUnsth7cbUe1RP8CBHHsI+MimlhkYxl0qjZ/n+2OtAjD1Op41pzzacyPNM4QJoGa
MidFmDtkK4I/kxufnpoukqfowpo7JiWIyH7f+HrVTO3unpGMkXIWpdRhHCUfUWQmPRxx1hdXD20x
xOWKuw0Rtd94k4bb+aZ4tZoQlC2wc7IVgS7JDpXyLhjbwS/sqCICRFTMNGxyhzge6MpL2TF4yUZX
tXFWlpXOjF2Vmoe3kfJQyhv3fj9lMhs4l2RhNfvmApsnNMCbLe8gk1p0KRPhZkJcJ+ZxqqHVF1+W
IyK2GlIFYfy80r9rGOc2bagky2jgNCI6Tv7OsnHWV+RZqEc5DzNMdTCY0gLsv0HvCwkZAoSvNpdq
4HUyhTIfDzsnnVOivDT4BBUcj9C+NPX88QWD+BDgloZkyzHtb6Hhy2YFeTjatzKjOg1pghCrZPox
82yagTTaJ3jZ08oSL+8VLoHATy7LLwa7uw4BodiixL6/VObJHl333XBbFuYGvt4Ixd1A/tjfTe1K
wwkTc+TXIMLbN5uu8gksQjWgN4Vw0uFRXv6HitGAwbPniNh1+OpW6ONtFvu1cCadT92aCdOsgvgw
VpFDF9Sf29zptFqvGhpwGXpdyuP/qInkP3YPbvWPAGRuvFr8CdwM/0Nic2G7wsRqQvLMRqzQ+jvV
LFkBRfFzeUIAOxI9pFbFCYB7iLXFCpx/Pv6/ad9CMzAKJ1NPKxg2m0+iEj67+p0jVBACv2UKqeIg
9Gy6T7YtxKWfIBIERNp/rtjc4pkD3Be0VUMOp98sMgpFC2N2/iUIhSr9P3fT0IB2kizPVCW/NyBD
DbkYgqyWMUwqaRycv00HjM8AoT2M/PNDuiQorSsG3jT1lamvabSkZeEgI/JZkZdJrHI9u3CyA7Lo
aXwNbbZlHp5qBYS/VQ0P6nwdIYrMh7dnokZztkSpkLRRL87OejyLS2+owum8RUcfgrt41++7dPWP
7AuXUUfOlhEuvwsgwZuTOFpTyleHpaZswaH+rLl5iT76yF21FiWJk0sx0x8McG1UmNMBpwm3qOBk
/WKpnNu4VlkSsNPy5iEyGf/wSYdqniTIYk1V5DGEHO6vDMKrN/ze/yL7eYM/Bg0GrC3WhqT0+wFy
aizTkSHwwjUrgnl3KgLhxWo20H8AmBnBTOz1lSeeqn9U7f63nR+tLdzLWp0qwRZWSeqxu0az0MYu
2Gctq0Hw6B0U2jSqDFs+T+9SEcdZohGHADnYJpAxceN6jVdcC55xdgg9Qug6zqdKigaOxEBFbWzz
2eFS0hL4Dd1L9I3L1AlhkKtpKBh3xR7izI7dQYP4SAtmHhU/djS6UM96V6+iTAdwsnGXSdgOV8HF
LqYrg2sd41bPROz571Ln4IjWAGAR5XlEbNZUhsX2Ms5kQHgqc64KsxmoXv8d8TE3jLP5YA+/McdR
vE21ntdtU9bvTse5bkGP12biwJg7vGojXkXFrtb7ggp1wSs046lRbcVuSfVaDf55UfJ1eeTiSegQ
I+aOpqRQhGad4/3fTUO5IVQgnMHAPrnNTX8gdTlVmPRVbt+5I6bS6pA32RGqj1X1tTFbEzqlFPNr
y6pVvn6Vs1XDi4BkLpDqQEAIPI0R9PDKqgsz1Lzd0YfMPLVYBSqVNRCqLwVXl3o8RdiebDpHAv7T
Dgq/f1RQww+tlu3zw/mORv1Zqghi1hOjHlXgUrJcTDGUmCZnHbdef2I7AA0e+K+eBD+lyrpFmTX3
FemKJRdVvVPdgvzBamA+3vnylU6WeaIeURsm9ABYg2VTV3kMWWtHwvjNoU8eg/au3c/2xxRYScb+
wTj7d+qzeCuSfotJmZSrV/XWNchWRTaHGL7Gt/EX2r48ZQNOW8alBaafTPXN7+hkb+xeh/5ato/c
c7ZqQNIIqUODnFtWuteRvpYqTbmzik4qg6f44ddy0CdXSk0nSnIsv9w3c9xtkBQjm316WU1C+Uen
NNokW9Oz6iL4xC3hgF7wW38LFaajsqFX8dt12+k4Rr9Yf/NpdRvCSRyP0/nPRcl29EgbOpX7JS7C
7B1qAXgcTUeWu9hSu61xCuY6N/JcHPDc/0LM2gGFt3uaVsqgtpZuXcTV7rsfB1voL7GfKpq4USlA
N8qzrhvjijQMQm0HIjiV0r81eTVm99AOCG14VT6PrcbzLYTb4XPE1Vuu1CBRPRSflnr0EpAvOH6y
SxvugiAussCCpp0Nhp6JGs17edn6PdpQ5l8L1zjUdEik5foiCLOWiWPzPEYfILFk7yjuVF0nhRjO
/fTGRhujuZITLAvCE6NLe6oKoW2rJ7ARBNqZYzRFkhDP6W0JUlHoHlOmDUvjjwzqb12PBstqOQzI
tdo2RWG1oSTaFjNeeearvsaomSHRFYit9CpSU3GJoLbA5AOW/TMrx99+zPtOgfXZfIgri9QGHypg
9cXhUcw8jUTq/Bp+BvbKgg5og8+JRjLNPMe1CRJiO553RCz7CpuyEch/tRd8VALXfaxa7txrQZ0/
0S6dLfU0uBjv01mrSq+8AyHsfDKXHf003Qnsg7NtAz48s8q0o3hQZ5QSMWshWUCwaphtsEkk4dE8
6H86E5PnE6Oy3+L/QkYWhatWPzNXD+a1LeTxh+ezHnAXg4ros60/xQkjZAnNXNGVvqHkI0xSSwWJ
8jcNKxSkGXeW6sR83vl5KAk3zDs/4mHevEnpPH34md7VQzbt0WWJ496J54aXOYDdQM2CC5lGawly
oCXUQOQoC0l+75v0sCauHrq21mvkTo2HmbMkUaKyeVUEsdkuWYA73Dl9gcxmoHBTzPuKEVIBSAEu
ThrdDld8Buq2rBVsnAx4QLoM6xHo32CQmcw4f/t2zEEO5Vv+3O97GIJATGRu0aMJFHlC2YB0CNMu
/i8sbbNBgcRvvrpfvnjAeTHFkqUMk90peH7s6cvVWqBg7S2AUqmoWWsdZDe3fhX2VHcDdw22BOfN
+DH872cXipv9Vok8upv3rBHbrqL9nLeZZuDRoSmAeYIWQN9Vx8cOduV5RqBBfpLl5QsBaSMPx+gL
VK5vFT+WssLID+F/ZfblbK1JwgKzaCIwNutt4LHIGkGMUYWrwBk/8IFNrwU5K8pP5I0pl9oCXZcI
wN+6vi+qFTsEf/YOyJQiL2VIMAoP/McfzUYc5a/RY7mlz5wJUKB6YoDH9BhlOyW6VqcCVenunXBk
RpeTzyZzWBOiXdbmOM68maMxOcM7P2FMu5/00pCm4FhIalkA7QzUjNCCF1Ig7rfcuwfAQGsyGWOW
TVojlIOeU5Yjt2nHroOJ9DsNMtsKqWAbJgSMvNlK8897OFVMWgAKsa+As1fLzEOYWO6qQ6nVJj0m
l7NIdEfkoqB7wywHOSFojKbSM2/WmF3feyyDc3CBO5z2zoOUHqcnAOp9RdOnFERl3qLZGxRYRtUW
2OzNzu9Lg5jYfEVfrkonOAdyc7iCYlqM4cm2w6bfDjdOFVXWta/hbwbcYUUEvMLKXPU6jRQqxZgB
mVN3p5WNipFG+6WHXgHdYugVoci41uhDccWmaroGeK60JRD2sqL/FhvNXi25Kw0uN8n5r3Vttj48
Y41mvwNuPElyo3vJ4ATEusDjdclzdd+JPfKgXeE3PESE5I4kyVPh6/4t3DLgoLisTL7M9zAV4M2v
JspHOwQPMXAODqRWCwRqh0HhcfvnXsYiE1/0KORINjCT2ErGQ4/qUugM8EPBaKVLP2NqiRGFAhYs
4KJU1ZgZdLHd3ElBYE+fB4f6AeyuvIxUSZPzpaTNm6tFhAK3/6yiyaG6dx/fCJ3LAEhZHMvVlXfd
Ud7nyUoOLPRxIrgZbJVvCjx4zOHsKvMSg8JpDUPan6Ksx1R6StTsboC0SPLdQv3MScmlLJ53dDOg
J4vSN494SXMwp0Q2oLVTs8uLMZgfWRGmz9/fa3U+CvnrCWdq4iaGfPhhc7naWEZFCruPFeLcQi6A
yHz9SJbtNIKW4V32KbyFrf6jLuuNzfrWYO6TXqcc7f+qKL0f+GLRV8dnnoSGzfSqH69cefuddpJL
he212ScB66GQ0PvykzGHlLC3stqSfDdWzDfOjEHuMdTamXGSJdTyAcApbqPKgPxLA1IbguFNmFyn
OKWTxnSLHNSetgtHv1uIPtA7tb60IP+11tin/6wE9IVgAZ7dZyjFPJcFE8jrHkN8jutWCpZl/Apv
MNgOkthZft8nT8NhDrGMP3KeR6TBpp5gg7qIUdSK0ThUCUWyUfsq8YKiTxXE+sdjGs8hzeQY8sho
zcsihCN+C9ejYHCwUUqNDH51YAe1qMNPzX0cZwhSTGnGpeNqLQGV1pxfuxNjRMISkBr6EFm4sC+0
eLejWDsT44v4Ze7ys97EBnYC3YDCmjtZt1CEryi0H4rJTG/Ge6yxSWDqPrwP3sp6S2h89BFk7zsD
AUSqbyyF4sVE5T3U7+eMQ9jxqH/SGEhFvMcmzBwlmEhoUA9L+SNCGsvlAAV2aHhuF886MfuZZgHr
jNj/e+95LlqTrlhUOOrJfg2clHKC+rLwrvDb8KxuBSEJ4CwABjlQVjzxCWqbTfO4/TNQWgNeh+rV
gZL8SqzWQZ3Ti3mbiT7+YjSe77FbpBVO10kqEG8TRC+Z76RI1VGK4wSwl9uKKs0BZ+noTyQKcg8v
1LSAgsid+D7pNyz/DHRhJCQTlQ5dMlJNwxyWv2g17PPWr2KBbNdaWzcVJ7TEHtT+AJpvcwCIUvdK
FlNWJXCS1oGPCygwVUW2F8KqU0nJZxiOKjOk2QiuLvBn1gu4DpJX8rncRcgoBCJ2Ym/goNVM44XT
fSrpsJRfRZTjmT9xWi8Ntbi5tl+1EoVP09BfGO9I/zWsLANzZLaRE6zu3kthNcUnRqoJivK/Wngh
tYQRg4g2URPWHpl+2s/q6e4I5tj5cvHH5UbUVnScDBc+cWR90R/L1DbZog2iwtU0e0BwX4ZuFr8k
PCwPq2evSxe++3r4Q/e2wGNA/M+jzC/OsWjhEMVho267ISjQalPmUZpnO2l4vdSh44kY+6QPR1EH
XN++aFYLD3E5BLbE3V4eAHeEB+9pjEAPd0Eua/kUFopjrAanNJaYR/abpiEJuAEQtzu7kSWifwZa
OE/1PaiG24t8NWKJIVYqvHMfWi5FzVhIC/UmNomccMGMrpF8g/VYqEU9DURHVdzWVY26ZieOgRab
nF29AaY0cwsbScXO3VdgEesehzV/fJe6An+16NidG3GIlyTB/hGCDcFB5b0aLdE1vHwbIsn0jWyp
M95YM6kf6/A1d0M3spB0JoHuo/oJ4AxwWxZOZ04V2qqqcA0QAtx1C+TA2gB1852b72kALubx9Yy1
bIqSFA/q77bLzgvTchtpeXaGs5v5IG82RL9pbH8tIRMc7o73eIX4VHwot6w/pC74BuB3x9GDgyv/
u916Q+tX1oDKf6CKMXtY0ZIoUkvpmKVmrcpXQPqHXp0kaUDCNL3AxioroAW3ympsyQbSox+ki7wx
hrCpW3gVxQ9+r+ucdaZvqRkd1mOHHUjymDtjX1WOxLCga4dR8IV6KOHoJ0o22enFHk2oT0AnFtw5
zubZUoq3S78AfPcTj5sLmGempc+12G1UaX2Hm617BsoR/LOqKMR3/GaDkuaodkEtZ/RvBy2WSzor
Syk6PQ/aW1Bo87jsPiAYNuSW4ofp8RVlOJtSiAh08eWGYXbBmMjAONazOqgZQWpQFLiJ4JjGnkRE
0JsbALy/e3jSHI5kLWaAOM4A1RaP0k0Y3fW7BWqZvVaMKEHyMqmUT5zTgSCRdBzggYfjv2vX4VD2
4P6QpILxcpqITkrhgvnG0VaTeox4D+0+ofj172xYOYYqxC4f3TWRwiqaXmC+1P0UH+WABKSkLJXr
YOIVPM1LUshT/onzq2AgvKx1zhTE6v7vBU3bBoVq60KWADwVbHLQddtLPHDIAU/LADp8tsFx2Eb+
EFQ1tkPAuDZC1FiyRoCd7VwUloEkLXepl4zPj/1xhLuzUi20VJnc6GcwwOGxsWxNjyuoVE7ryrmT
CkUWNsYgC5Q5o+TaYrMrtd1Bznm9kMf98wb5PEQJbcwUdnC10U54x4yJDoTuenL3fcgXzd/m2VMM
ovDiuumIg7AihTNbFbpA+7T9aEnvt5h3XUlAVKS0EOodLgJQh9nG1URpGbz9a8zBnumgnDrpsa5B
/6IDRuEXVZ7t2Gx8XMIzgI4vFtlpW1fxzWGpfGchahr1fbShfR9/yN5kUrSVNaci8PEYSgAVm3yj
uOopYn9BgsI0yYK9XKL0DZ4+wBDkzhaYbx3DkQtlahNvQu6eetgPuF4jgvt2W7PHlVGfmzGslNTz
qWERo0Y/Q1SKfcLRn6LrMDa4KVkY0C9tEoSrJN+KV/xINc4kW/+QH4Af5cEOs1CEgiJ13KOb1Yul
Be5yVC17ITD3Uzu8jeC8kwarpDgq5wzRH+TIxaKXEamtcPkOuFFfdMMRPJrXMz2ilUYG5rGVVv23
d5NXTiDBkwVCihTk+nMuu+xuNOE7he4fVjpo9wiXTUTjVvVApcZOEVFgKPhGCuC7z1PrkiSWPj+T
olU9ybolVoMDwESb5dMLX8WgMLST3vrNaH/5kuORGJM4fqTZOYiBm5CkzLzVRc+1KDh98izNOTgu
OJkAMdx4SdI3M+5vs3wHnBPAB0n3XMC3SJCo4LN4HsFyjrQnNLvma/80bqoOhAGSP1ZznLgXBgxH
VvAKFPw2aBPFQJ6r6JYi0eSaUkDnueRXtqZcMBkkdc4b0CgLN7jrZ40THxWXXEJP7XgYLf3rVmks
nlKR29KMDgCNX+lJnhKy7t2/rmo2cnkwT8j8Uz2VR90vHYVfOevD+p06aQWRNdyCY4DFTtvLEBYi
tVS70odCqWzyeoc7TMdBgABKftmqNseYaOKEf0t+y/wpU/e6M7srXc1QRb170NXOsd4CAuu/dmFK
3uX1jyqNnYdp9XfIfz/O5uVa2qofI9NjJfiYV+nnbP3w2iHz2g9sHtirilaALZtxIAjuexW+JE4h
kkHOY1JcyxX3WS1giuXaA5vcFKv36p1wbune8lr/J9oB+BP1Rd+QxhnaYQ/9jlV/3UZc+5vW0utc
t9EcatDeZ1yiPhLXhRetApvxvNUNgU6ILKS3uF0PBXPC4d+P85xP/GFb8ctjgUPDQ9toHt2AJaA+
biMzLg6dg5hPSJa7DZ5yGt0O+GzXMs6VNnAnIaUOQ120bHC16LqDJR1Z0wQtOUwSdw3owYFEol81
AF5h1+WKvWiXcbnHrgxGcT1QqAX9VkKJUKLptUFAQWTVVP1s+VyDqowYQCv41buDIxdmi04F1Mfn
LJpxYjogbUA+TU5jAyEQwiGbRX9le/xlT91JmdmViimVMXMwaq5D8SPzd2v2/Mko4OTeoUoesgX0
Gj6HnQ23Vs78BkExCZfUg4lYEK0+a0h2RAp+wzvwbG2XeJwOXHK4AH/F24OL8ac7QIkeFbxEVph9
SsvDFNrqD6+u+F2a49w29ZS2i33Bl0jDgB5rrq5HWdZRYwn6zKA+/xy+iuPK8GRsNmEnXER13Fek
EKNT2juduIfo8y6Bb4mQdZUjMnL5GL37yKoYw0lqlCeuvP8Yzar8V/7fey/sAnB2+aIFy31gg7H5
gJnN4aqjuQEV3iyide2VBr0EbPspkqCHroYvJdahWV9fv00ztmPkGa8CDDnLTq+b9X6sb8l+vbow
jLl5IOZGvxDYSEnbwGzp+0S9xEL1zIGfqiL2htAPmQCUcuIxBzdocFdCLb1tF4VnzKnlpkPTcBLT
xDCDmuN6x/PVnabdR/0aJbk595DUUr8xcsownEdxZMil0YlSZwTX8NNs9Zz/klHxULgoF9Iv5VM9
xxx76XCUfgBP5W6lyqjsvkCErP7Q2J0koXyNEMHWe0A7Mi8hgNyOaKisu4yeb9K7MGTMzJO136xG
QyF2Oipnees0dwzdCRTj942MT81e+c5L9Yz5G3Z6UbS8CJg5AIrDDkc86a6T73USbt/LA/5RlQdF
GKBmxAMMF6f35R166r1JuxiEXfRBRnvDqDx9yeYqeqeYBOSyej4sL/VVXA==
`pragma protect end_protected
