// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:45 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
nB0+SJnJ8ZDc5Z7ikcM/y7WkXL5Kg86flfu03Vgj2VwrxLtG/kW4loJBZQ/AWhOg
aGvEwJ+s7r1UPB6eYXPvEWnj5mYq+MCht4LJfZGdVSPGr/7AUIzaz8flu9inb1RC
ynFIlDciKF2qB3A2ozIGKfkF6+1y3iLsy/ofX1IKWFw=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 4224)
yasajoizGCRekEHRZSNdXEm8/Y8cHiYT8qF8ujVQxwWvFl0cPIkuGZ4joH8no5vq
bYpTblBKISf+W2x41yPROje+kvnoLEmXbiqAztVZN1x3IRm6EUL/IAALMKxcIDL+
r1+DZoISy9kKzDVDvbh5sElcIu9fhNbOoYJiAgRL8xFvS/wtsCNRqCMBWpIBzN+C
jReWx9VyYYbC7t3drx0xKU8r1ZhpIJ/uNhaNrRIg/TqltcY3xnM4ywUPC0HW90ab
8DjU2sJDxg3BIrvgy4zNIGVa4FVmY+Gzw+dDBbBmcjRXrMDPZ+FB+BDm1dvhJppj
0M2ec2NIQEMVhKXgSKs2PyinJ0QFxCTLIX28k16NBEAkw3R4aqvofoK4oFiNrHQt
Yk+AWu6+ye9S1AEzWcXP2gR/nMwnzqimVfmfBZmvLC1tHumvFqjoUQLTjM/obwQt
DplXT/OfdXKFUA5wChL306fjYZl+ws6oWGBs3hky3nG5zarjvKxw5fqqlNMRfYIx
9fc/GBpgWfl2HsshPZswDe83aRzCRvbYHuTx6LM9+7eVrgt3sxtEK1n/MrM7iCJC
Wki6F19u8+uO9AOgrutfS5r8eYhGD1eLM7lXn1XEMm2rYsMndpy2h1B69nam0JT+
Suq6I+cu/7i+JPdWK7plsP70LqBETttAYy4GVlXM0xt++d4H4cI0DjmGapWsrffn
Dr4esZll955pPX/Z0obIRFe23msYfQkpMbe4phLdfP0kL/llPjSQ16Ckbtl2VFZa
igSG3BDoUM2ac7gCunWv1UwWEZmb7fScC+FlohQqbymxh/qOQmDePywYY2sD0hNo
OG20FEzmHPNKq934HfXfbQgqoOrtHLRs2sEIqFRwd5PHiT2wTDlNnjTomR4EHm7y
D/KJbKTGqoEl0wpuxFkSAP+RPh/OTgUj1ucZw1PDCvhfqTrsTb7GqvMZdnzzJYfH
fgjs8prVGfJoV2iZ3KcW064ozN6C57SIpQsc21gieGI9UcH0sVeKW3tUtCTB5pNF
L5IJkjrQ+VlkCTMIPMLfG1sdvbW5iX7Yr0HC+aoHzd1Odx2UaNSiUGdxnvN0Js60
OEH8d3T6RBwXOkv4t4uGn/72qwTs6PiVWYFnFPazqi025DWEQSWhrciJ4y9KFjQq
HmCoTPoHdl6XXeG0LAuSRbSxXhT6sGaTiLxWuyaqutW7pcCoeVSacIWJVeUkfeLY
PqNH9Epne5k3NrsWQt8nKZZAlEj60uvs40Zmpd4w/EgFw1Ak8fM5nhOgNgeb3tQd
ynOCahZhUBgb7FfWD5j64UO5RLZGFFlErdLDk9w/LrwMiQV/AoIw3iW4uAWYFiAJ
2M78ydfsnOeTtpkJt0Ar0uBoTCF1sjRSyXbc94fmzwvbuhG1k7O5LzbG8I8ymMS7
dQCkZ0r+F0tqIGFA/wfdnDcHJ8x0IfDs1//cF+ddBoYDmrVroJQq6RKQCzGmwalZ
1eAncHE1sXsn1SkLwhxancs7QM6J5Gixj3PpqtTanGmNI9SD8MTz/uHuxlVfp802
A2nQjY/OF4ADDoETfaSg64HsKX9Wd/hrh72RkhLcW5+YL4vaklHiWfADN6PoqSWC
/z5WAV9LLGPqAzgOuw8Hzvo/pSagaE4HZatiz2p00X6SV1n/Oh7+DX4Er0B52/a/
iskQWu4GLQm07sp0+lJw7Lo0wLRPjuSYd7bl97QxNq2tVe+JktZdv/ebAQPRzUU0
7GZURn8UwGIPBZq/dp65P+gOVGtKz2KuJMS1JV1gW/csyYRg2HwqrGFKfP6CThqr
h1krqTev/iG6lR7faJi/4zY3S1aJek0v5DTjd7EbWMFI+MnNsXMa2sbrxUZZ3rX+
RmWKV0KJWpmVjZOGBQ/bTNxbTFqZWFpxChvU4F8Dcvi/0eIqD+nHAyCLg4dUmNwG
Mb4PmhrMuIg+D9HzFBKUcMy5RbTiz/SJ8LNnSFZ7fbe2aBJkUIIpOp3AlX5f3oNt
21T/s9xGkEOM695LRNKoJaHmvOyi8vGrw0kPovbnYRPZdIKMxCOMBODfJu8iuetj
kxonChE4vylZ3bJVbxRzJKmwwUsBid6jxOyYjkgTlbUQl1+yVQTEUtE8wyyMxh+h
afIXCqnVEBXd/pyt0fLnTl5i2LGKZom0D8q/ECH1kJPcKExMoa/UMUkYTu1wbD+x
kc4lW0nVJndoqxF0lnKuaMniYNFKQp4IH3cK4rg347RQd3Yljtkdm8rOXtzE+DeE
nO2Hn/OMx1xfh89eTLnyXYdg89BnawCzPZ2eA5wwLPXXIbdEu1fix8LOShkMhVbC
EXqZCC5egjDEOaml7ncMblQfzxdBD8YBPz7i9ORlencjPcbLUs9HhrY+1gKzzkPy
Qb15yNgR+Gk7ZAvuYCq8OQ/cqX2MmiFb6roM1rr57IIVuSzG4v6UjogGxvFBLij5
UQ5cg8Ui3Y+vKNgg7mdH5VUlmBvLuBl2sE/RZY924XiJ4wGJoWRyq/w2WRvQbnAi
niiSx2wW/HBvB1QLpWEafEaAagjIR9KL/VFRXSDdJrm6gJ+zmcRIFw1Ht4akslHN
nJCnCqgXn9BgmZsHqx6Vx7425MYHLSNRxI2mDMMm2P8Nkxpiega2pzzCjrfIe1iZ
dt9tm0LlSwYr3ETUSk4j9iKjI1pwRjizcAhLFK/g98tH77BGUvU3SL7MjX5RarpB
oLzxX+Nwgim1Svy2Nl/bj7vYmMcCgQz5plzqjd0GMfIuycLawTykul1Zl8+LDfq6
mTG7ZgO89B9NsIFWJhV3Vn9O7VTR8bGn5S1DH1AcNflVb+txQDbXbqMWiQLGHkX+
U3AH37PNDNlxVHkaxgRs8wKDzjqSTrCpk3jaawz9gJpV4HmSInviz/OP/UdT+fLc
uQ7ANo/VUo/W3GG5bdc9fiAN3VOfaFioTynV2DPRsTJNUBfoUkKX54e08V+82Eu6
W5icrqvHLuVs/NMmJdMfFvRixjy0UJ30YhrRLsEvNwl5LLjJPMydy2ChK/45ZXRA
IHrjINVciAECfrPuwcd3WiBZzU5PoOP4ytJ3W4huGLlMXNm/u6Rb2P1dIwdZ86P3
R1Uzku4tDQGknyIyPi7YepjaztJfRSwPRqTV/90zo/O39sUIKXUOUaPh/t9mGEVQ
1pRCrlC3l57uVtPcN+v/MrQ9bOyWTlpPf/n2VaM1Si1Jehma1fh3JqS/VdjsAg2V
7kJLrFaL9lWb1dgWG2SNHZ1kXElZCy47XjDthp+2/UNaPmetJTTICdQv0Xdzrch4
4vmELANleXGRdQZevtsLZYUhEPiKPT8NbT5OXD9H8XgqsBnxK1dJ/eAkwqIxmMH5
5VfKctqp36aCmMUwlhQylAaRmUfbl4RdmkKwt5sSxPvaRzowaf7kbeO9PPl1PeFg
VLK+6e0/I+n7x7MRzKAdIqUjbOaVi56qVi5rrDP4DGOuZB+zqCKux/GTzq1zvipo
Ab5yo3OtK4IszH4xbBx1HGGFBex0FGUGW5+k7D5CEpStmNR6EZfWhGQLTLgn/kem
6nEX23MmtivrX4tFVs5meDAw5P8sZKIaHDAl7odTdYOk+eSHcyu/VYC2ENtA96jN
TjXLHKg14XouGS5okELHKTJeMUjnwGa61CgvfvmggCuJ3uy2TMYeWdgOIdclkkMP
KWP5KRN+gmXvtw2bVFqACKl4oZhefsTT6KdjH8li1wUB7R5iorzMiPXMbX1OQ5lL
9n50Ica+QZTx4VnuKuwFv3bqs1FPo7MuVOEg+Z5/cKb3fRv8WWy1Xm91FNzlzQ4Z
LQC/GRPFlLGXOo2u1b5Xs1woW5DxMg7nFrnJETLO52CC3L97953F8aSXZrg+EylC
X6mgYPkqNVUuKVMd0c10VdY3S+5St0vvljehdUDwCJJ+5tNN/SDGHwL1jSNw/APc
w16s0IZNXnl9RsRLvi7eWt/LIpRLBwfRyNPO+d7A9liPVfn143GC6kBv8Pd7Q7/1
TOZI4h0jH3WRMxEuVhJG50hpdEimHC4yMt89KeH89CUwzDGj76GN7FmeSd/WhIio
LuIganMySQvZRXKNNHelbycOh8mZQX9hZ2kIJoxAoiyx65OfdTUUsiMJpivOAyIq
ppKtEKMK4mm9yLY+wyLmk41gTq+y8F21BF8z3zFFZIspqjfQauU72drHLtxX7dnm
TLF7Mkq24+jZRKjnUXWY3pseZCHu776xEQrrNVo4qybN5Zq/LVNvdOx359qE0nS7
aecN7aLGRx9JW0+/8PQzGG3d+OrDTGW+BgWydY4TtJxM7kWs4BAQNEGF/LHNd3Fb
IeWNGXFrvhB2DuJKA5zoDCtktWyJpxrMjhChlhHXy4vZ6MyQrH3p0nNyTWrJ+jfS
9WpzkamH0iVhW7KwDW9H4eqHVuXYvvLVygdspLZsUKX92v8vTVH+RndqwDC2Yn8o
yHWIxvOInPHfmbkZ7iSPMeSQM+v07Ahj4xZVG4492DBMrkBCliYmnJY+bCU17pMv
Dw6Cl2/P7qKrecf37wAYKsCMUgF5GvGoXZlXlsLEx5FqfMIIojJAxDQ6/iW2w80J
e2nOp0vwpxUeRwEmQrheM2nv1fOCeBrt94sKS+R1XJCsmYJ295qNjgtqRgXS0STr
tYrqdaQk9TEqmh3ieJWyEGGuPEIDXkFjPHCW112TC3k81hZVeRCmzysSfWHyV50O
PkyatvDG9pIo792QRLGlRhUcvd36O9iTTuZqqDUkm2wXSyu5QjaIB8b8iy+cVtH/
quwr73J3zHS/9FVjtMBm358HKODk0CuUNBGZ2UfYxuqs6vs9vdTlcYyEq8/A/Z6T
W0O8XDsrSe7cj4i49D9I7nvTV4/w9XnjKVGt+KB3tnFARrBWbzo5EduNlEvck8MZ
4zFTiEIsOTwT0t128wfSn1HqnYMdSJ9EFvDmtrS9ktf+LN+yLxNvsokU6cwFobi8
jejgZMMyK5j93elU9sRnjFrDti++r+ZUUVJMF7NN4fV2OKM+i59PJgc5Hj7yRZ1a
da78MBBkQ1WSuDxKsBBhLHp6Af2zs4tXw0NE+Y3Xxju6hTQMQ1lqkTezPHt3WQKd
A8kHyqhCshCYBzyb4GDqmcI57xAs/eg1gcBi9ws5wdgq2EqlC5LA2BuY+OJS7X5q
SI0O4jSekQoueqlVWMYP9fBiKvurdlE/roFFFEeclH/DCvFiPBzCA4OW5E0DRseS
1WXtpHfDrcod4VmkBDtDE6J/j7KjlavxB3bYLHDQiNfZDa8bwDSqaJMwKxWW9Ifq
64ujxQ5ksgDwlmzd/zoTPjYmh8EtUIXy4Rv7TiB/L3Rq1OjglJl4pOzWDrveIcUJ
f5rrzg8Je4iMwdaxYCajUJhGBRjlzE3wZHwGCyUj1iccYMe+RNRedvqzJUYQVu2f
4/hc4jWIV2sQbs0yYX8IA4Bap1uKDk6KF+w41SafzP0XjA3ZL9UcMztn1hHuQ3Km
QLgoFsqbsxKsF/kEk5x62hKHFdaenvDd1w20tkjx6k+QRlMPe3GwgL1yVs/OmiaK
VylJg+seFomNRO/wybXMr6u0XivdR56JYGfwZ2eizH2gYJ97Njbr1WoRGrD2YoqX
/9o3Yifi2zGil8JzouKcygSwNFKYjSUdAm7xvstqUI2b+FnEds44LVuXq/E325g9
`pragma protect end_protected
