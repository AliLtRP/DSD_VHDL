// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:35:48 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
jAK1tdpG23AD9/xjyDOxga9BerlWPD3zJBM5HzfgI0aK3BxJOurljL2BTTJSyLAW
M03AfY74xNLEoF7bKRg/YXYoJSols7ilZrXn9hw3nWmPUA9qFgmW5u1rK/xZiiHT
lX5yVhH1HqwFMdpy01ZAtj2HFxG3dpiFawfVly1W2CA=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 2448)
jwudgEPzMB9Xu3pfTETQRbGcr6SfR0Le5Qkv6z2o0QZhJeIfJ7GNmbedW+FjI9U1
6TLqAkyf6owBgRJnbODL2yA2eDyVw0rnFF9moMwDhTFZjdOMwjAg5d7FRNYury4X
ylkpDqo8n9XHC7Lrxr/6IeAxKqjcisGGWhFY71++1KMYwnqRTUhilaq+yNUW6w60
hxZiNlZejc3KnuzYdP/rY5/IVjv0ZdpuL/M4yUQuQ6y32thg6Pn1k/Hlso5wr5lM
DCMsjyYKzIoe46k7p5gSYXcE1R3I0W8sYRTIn/lGi0YIvP6ZpT5LFNwUXSOYqtQL
9B7Pma8jtzss+0mAtvM13MOGVsMeUDRgRjGfwuknh70JNbZoBIYFx9OfIaNwVp4A
3lggn5KfGCOUgPmEWB0TOvSSdfbDLR71D2MYUh84giYiH2Y52gc+0zOx3HTlStE+
RElNSSphwoRlSkM50kXI8++yQSPFS/hY3ARIsXrd00S7EMD9qcd6UTr3zdn7dYj1
oVm4/q1Pvu5vxu1TtsF5gSxZ73of+5jIyoiF/YeBFmqKSfbmmn6sZHn/HD8+6hd/
B5U/Y/QxmY9NBllp8Rb0oLCaBtRtOOUnbdyhaURsbgsm9lHaWf08ZO4zXrB4k5Hj
1XbNxCr9N60JyVxrrcaPqQ4jvV+pmqjEIR4Jq1yFNDc5NLG7pxb3y4ctw4jeCC35
gbD4M6mVx+zNvQiG0qVwftVhoXPBaxzT8wa6ji9o8VKmzOS/kZ7h1ejOJwdbvr8N
Onrj3BxWpQLrHCWDyV1uORLidFpOpWwCLp3eZC1lhKIKdyTebqYn9fGA3ZynlYUB
7pikU6hy9236WJj0nTrsIJzMxBSGvlQlqxSQuly/b1MJYK4bCu4u3zYF2pEMGHwN
fh2ZiMJSFflE89aa4f0JKhQggVJO16w0nMqPfJlkYyNyLJ9AHOMqT0f37BUF3UDI
viGW7C6vShK9i7Wuz7MyvkWhNxROaD9dfAXxuD7jiwxmZ2dihDRhCZRw2C700AgC
hkuGdqdfLZbBwQyCoJE/H2WKBQ2eL5dRzKxLYKrtu85s9h0SmQjOr9L/+tON9MRw
a2gYa/2eS65Bt9mjmMaiYiW4ndDm+yhgaEmAK5NTzHcTIuMVjXN2nCW3S/XzuF87
k7Sx6mPDREF8ZU3awvFwLlWgu6TGiuYUSW0q0ARbDOjIfAUAcd6GQ286uMiCbHe3
qT15gXHT3WVYNlD6OBFTSsGqVfNdhbBdVsm0/QlshA9HD1yp4pQxom9KW9jG9FHZ
2lYBc23zRu1/FCXcNChVsDuP/0Oejtww91NJJh0wpclimtI97Zt2o69An5q2PRxL
Bhp6dcajjOoMnFeey7Wn5UJmVvZwUBmgoJGUW0mojh5QGkn0KBqR6gVKRN0Iatap
mOD3z9FWCueAFKTiVVBJK9a/Bedbz0HW7ZpAFvLkUdXsflgV+fsDksgGV+jzKh4v
8vJFsiKChfi6znObmWch5/EuJ7+kdq71xEj4l66iKbUpn8wIgGQn/eOZt0PjZV+F
UsieyiAA2NpJM3XLHAuZ3zPk9M8mF6JI/iVNTmD0BOzHpwa0SKoHpZ6s3HWKYrku
qYALq4t4M02q3qOf++48JPw1gm3tj2mWmDPPn9rWmRK42yXgvYkBSuw5+yQw+Jtc
MLCOWPxxY3es0QK3K9NN6IE0UHXGU2UNylZYuHfTpQvmgtcdWffbM+7FUQM6tl/n
vShNbAN1oeRrT8eb3DR6h3FTfgVHy3wcjWdgqWONVh2UliXFnC4nwAoI7Tl4bhI4
/URiBe+4evMbdTMzrl0plk6VKI8B1D+yWQsqTcwMuHqeWkaY3lMpqNmKx9/0h2Dv
WZfQomSCr5sGitOkxU9sG2SsF/o7gPlUPNYD7xE2A3s01OeA194FNNNC3mC8vmbU
z8lRedRNsJZnA3+zU6kSp4/qwgwDERuXztja3zySebwx6opM4XpvQ4Ce2PvtdNlE
0BIe7UGgw1bkvJdWUSftxX9BY+MKKfLqKX6U0UB5pRDsZypKyN36aBt8bHuJ7Oub
sK/ainluFmMQklII+Jl9pblchIzCJdDV8dYdQFmEvFIbiyAF3GTTJdMUaKfwS2KA
hwx3kCcfjNgOQSs9KhDykVLS+g4VenF3fxvhbjycRSdPAN6IFwuaW3C494Dnq/ci
Ixb7/vnGPv5LOcFKzS7Xb1Cu1uyVK8l3TbH8bYGJUrCkr2PIFshaWhb734Y+Cmt5
J2+V0sNNEhwoQFozFS3IwVIjO5fNRnG2rw15ZaToF8s6ZxOswbX+ZJ+jEmriubWf
ArDbcgpgDetrGk1tAd8PpMGzwwowgNTqlpIgvUszLMUh9SldOGwcAzaH4gFXnraw
jJ63u8kAQTBIrWnRoYl/++G3UTX6zAhmb9BhDkQlgXl2e1gFvuTBRAF0rssGP8Av
8DHcj8gfr4xRVaFCXaPZUrRqpFbE65fU1mhlBFv5Cpbzk1I37mcSn2/mcHD97jLb
LLyMvqnImCxxxyhDIOzz834DWjaaEisrAcQGrv4kbQ3gBsmjfZ95pEij3VvU+uvH
saQb3XQ+vaNuYvLS8rxR9mgA13Gckmi+5sN5gPJf+w06+bVRypueO7JziSzRO5yC
EP6IR2p5SAgYb8AyxVjaQwTXu0TzJZKDA8myaAba+Sw877gLef7l597yUyoCO9pD
2XghQ4eU3coIsh/+MFhiKDVGjLuM2WmNzuwKQ5IMwRVrRvxs7lODZzJie+CwcgAH
G7RExi0Hj/nHjYVBt+jC06iCuHs/sLZ6fDwr1MOmc7DU+J1LcMRkMpzIfkhCl0AN
3KWIPLYwFiwxh/O6xKjHterX8/EQ6YTtwNfuIKVooFLpLH3n8Ggq98G2LQBmMwUk
w2ZToluDOFss5Qo7rikI+LSmeoQeitec6B6AJA0KwWHcYm5kCxALfEAmbqkYH0+E
YLxexRDdPA/uf5NIC59rEAkaSIWyDDgj5tIRqZtYFYQnijtlDJegWUGBt7w7Afuk
TwzW9ysHM52X5BNjrsXjlHi/LtFMdSWuVG4Zi979/xPVHKovMMi0kw80zxeK3YnQ
xs9o9NBsbiNWhK+8SUtE6TP4mI6y1SpvGgufPQHWQtA4Hm181BZQb2HJsEHt3fa/
Ui9Kb4VuhjlzGcEx7Adu26Xk90LtRZCX/gPLllEo+rZNtKJPT+vkKlFRLlCIUAam
cfGQjpYkdknLw3V4d5nxtBaGu6DauFk7FuYv2t3cHzJEH9zVG+4kYPL1wePOv5m+
`pragma protect end_protected
