// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:24 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
LmVZqghjckIR16t1vQueUznRO+JbvHUjZFnMpFX9jP/euPIRPBjMBBPtEpCBaA43
ePDg5OOHZUB6/yZTQEbAeRJUBLCv8UqGo213xQqg1XDsrdoxRLbvl+4eCUKEd6wU
GZ/8MNvnSdpXdGp2qj4Pdg5p9YaKw7PSg1VGJJ862ao=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 8240)
wQclwaiMjSSZMMPN1OYDK1KaGK4R3XuVQhHZXqXSlmJgYSE01Oy2sGZRpCzvI2c5
wMtxPlZeNs5A44mm20UNji4jMFQmObLM/TgbZGNOnfyARTaRzsTRNp7dune8UIAF
b5uNY7b29oOeqbFpw01VF2Bn5532bOFAYGGJwR2w0pL40Dy3bqm/A5nW1fwDhY8x
m9RgTyJv/h2uylZvDPoXJ2Vtku+vt3CWk8Q93wE/Joi37eS14YEFvciwFpPlkzQI
CpiCoojSn9mDDnCtz1vvwgq3kOYlXM5I9Z33RUr0H9+6NDKQDTAnWms+VCnujvn/
F1jYEmPWmO5e1vZjyAAnLG5ogW2ELo/xnlmFrxCOb6ohyZSi2Ixbz4O5WXJmatCG
d2mMWkO2tGc6qO2pityRvVWE/ND67Msj53LBpwHToe0jMujUiKqfeOfS+RuXgJJR
7T8BRKFFtO5S61/a35gF2+bI6JrnZuSQX54FocBd0WnbrKYHTJfKmWdc+qjOxL8m
dsYBvtcXRYWDMc3VWOATLItv2ZpSWbqkQ2HeW49bdWlYeepgXf7qiiV1mpvHIkvO
FyTuM9P15Q4lDlD3PsnTF/x946z47vUV1czOY3jaL4BgRp6c2T7bxqiWJz1oqNEE
brNLE7kwGe3jH4jTwWMeDPruovZZVsS1mtOh9sxFOlmFMIPT+Pnf33znR+SzBt6/
yU1oFlgh97N9WCl8Iwgq7P4e3d+A1TJ1zduyblnfhlwzyELJljxlRfUvBrI0esNS
mjhLa361Wztin7UFxppKl1l1DBsitOO5rtDI3Wwr4rk1PolK+l0qSqZel3To1LqE
lL+UFhk2oPQCzHidDwBBXWXFblFedrjqq38hC+XnP/tmLeXqKw2wV8jZ6DFIn9H0
F8aKMepAemUPq3d1QNrK9KYbB9pHN8zBWrLzyoF7cHXkcqWtkSVW+aVgUoIbZ9Ag
4XepK+5CdHEH5STFm+aQq+Jox4NBwsyv4eWl5KtqZg/YKVSJ94q+XfIA7Sv4n742
2ikyhtyppgaEuJMEcePoWnpHsh1iWgEqtK5pV4QTdaKsvyvG9KVJSFs56HS9iWY2
FeLR9vHuwqKPBegPjsXrdmSgXKOJZzC6MsZgomRRwe7//zTNg6FI3M6SPcVf7u6v
mvetP0I87Lc0gsxCXa2VZOU6TsecS1kL898j0lOBIqj3P0ZlU/GL/QQQUrGZ9msg
j8L4DWbHMrji4XgIa3FZj5R0qZAsGh2vET3Gu/CHxQVL0e8bz0MScnkgxkbheJqW
OW4HttF1qVc5q2NWsfPSiWMVoZd7N+F2VgQox3E6+uGsuPyz453TMRlxFKHDnbEi
0aKQq5JtJ3P8434aA6O2wPJyw9eeOlHkzvUVdqUxxaDZEYNHRhknZHPRxcfvBKJO
jbXXc+cPeC9k17g6c8X1R6p3fAfjh4nGoUXdeLaaf4NTVORj30pMqtakX2l1pvKv
UyIhIGcWSdsoqDg6+uz5q4frVDJ+u9h2KxC9RHauVeef+EFi/GK4FjhpHQz5suu+
4yuRjlmYMMS20mcjlcMNQuyA8PwinpqoxZWxXuOyzNjMpS0g8/S93fufL8eIzrzY
fvKQ/Ai+x888c7eYyF5eipEjZZ8vwJGifUy6lmndUN/AnAUJGR10RncG6fcjLh9Z
EUem72f4OQ387D3+O6lLXa6+Md9k+aV8qXPXQ9QKfpk5/sL9DjYKuhn04JFgiIG3
zukupae5KQmSn2dVKh6nUABxcTjeLPyfdDqwWXpGSMSFbEJBr1EIS7P8560IRGxX
E2gMpSB6UJoSW7QHojBKBw1YDtcB23v0lU1BgSI6H2F2BnB7rul/sDyrRbqX7/sp
Mph8Wl2ppaenuNl3DNCzQejcGmfbUzH1h+LySkST6lvqhiwKQDZkjg2S2A5mhqf8
vaIaQD48cQbkStW24ASo0tH8SllWJEAxcRzmyPm5mIQscYOCHHXEbApGs6wyUjj+
1oE/vJPyzKGZlAUcPYxbJz7RuskdlyfdRjosjrgV7SE1rIArJdT1pkwm1wZ0/baM
ITXG99TAOfYvoVzZEBac5Ld10MVJQH0sleJngvRGpR9kR1xHp4EQCzeLWfrtrbAd
PhzmeQPWbqi2QH02bmo+Gv7S1I71A1vS9xqv9xmvDD/269HMK79bJuJXlFO39tSX
OELL1J+ajSg3Q1vMDBd4ECez8JdafbOIyRfeq3fZx4+4EQWbIwux+DxtKFn+bgJe
EcgJx2Afp+IjPgkuQiIJMlAntXZfCWXiEvn0+QrEdlPmqCKibWErbOHo05h/9Lvw
Pto5+bka+oGZ8F7gMdS6zVBwIK+VGwoqQv+8TefCmhDRlkL7u68JpptFJL6Zwi8U
dVgq9z2BR1sDcUs0XgMKDpVsI4+Wp3SrJgSOcaIIfm1+pPuDPM+6q6gkCFucI0Mp
leXdjr+crNe7NTKT4SxtU3GXNY0NkgUGbDwHkd7/ZcPubLjMRcYAKLL93hOauCFQ
5mtJ6dsc6AqqLRvWr3J98Aenb3WyjshA517qEqOrPHSV+YB9OAI6KsIdBprps4rT
s1XOmI2saM8zAdHfpqBYgAAJuj0GG0zPhvjMQDuE+KuyGQiO1cvO44jmoo3V3YyQ
lrPUrVOovhA1cS2SmJP1xH4iVftAV7fruCXGkyIPne1PpBv6WbOCAr1jYBYHMYjb
YCqUPIucZ74aOvh6K5WWvdXOydt+QEi1g7ipYG70F6eQMwDbP7nSBXmrAEYLvrJK
csFP/E0B9gI7qdlONcdDMblEzsD3RjXDyiqV702Uj3075Huv8Rnn6TznDnpTgp2x
kww04J/CMY6KHroUOXTrhg41k0RZGTjQcmdd8CTURt5JS2YV4s+F0opIjh7rAILa
TiusLeblrLy3ibpNbBoeB6zAtUV7bA8yYQTEHbIj8lhxKcy1TjuDXUPpcTI5F2AJ
pf3rKNYv0DXbbhdH2+c6JtblTrSyZTiSyr3BbFM4a5UTJIqy19OeezIWjKig5BVg
YCgMoHumVHxX9kRTHpolRXEZmZdFE0L2NPfVO5bNzREzUWVDpaHsIVLX+Jnvu3fi
+q0b48KvGmIelgNPVoJw4wAjcMGMk2BY+/SbZuvUsAu7OkzQjEIQTF9UXZ6dFwXv
t0j3MBZ4npSVlYd/tNGxm9ecO1+XfExXknTA4f10EK0mp7evv7+ID4Xcjphyu1sR
mdG5QRtPgFVPqvI6VxqMj5G6Vgz6FptSwQ5DN0idTKQE4uiFGHToQeXOeM2bPpAo
vYC836uyexJW8TNI/iX6Sdp5Xh8G8VCI8odCNjMpzv9RFaz7lqu1tO+Qej3VaTzK
KkQhqKp002MlCF2vGxv+Q4r/WKlovqQ8NoVjAFLwzrPI4VndJOget+nly3PBgNSX
DcsLNi4Ufk7hW3mq2Fja97mFdnu1/RDqHZOj8KyuoJ7iaQ9ePn+9AaaG0HlQV6HZ
c+fBYG5O4OgUcP2cJKv2esvTBYKcLeJf+1U5CyItv+/rfltkEPg6nrQWvKrzKtGn
DASn5nqdiZcrUg2U4OT3mxeoqVnLeiMlZRwBwQhkvApMEYPKqk9TNmjsqv01zBe8
iR44FG9nogmOYg6LFthFiCGWLkz8KvJyWCrAcWkAuQby3kENjjj7veMujr7LwBwd
ldSDv4guz9W5lVtB90i5QpuDjI3biBu4xVHR9NvUhYgVVzfVF7H2R0ExUaCVnaTL
kkDf5AIIw1HH/vIrFWoAikXB82UfGRImdsyyxHadq7HriO1SANUVwOwK6PWCqfr6
qEAHOM+23XNqEZ1XiZ6QcaE4N5y3EsY19jemdCCyLumTAvGVcM8q1VfNtGj+zPdG
FXy+DfjzT9okjC3LOaFCGrlL59aqriblxvW+Wy8xM0IMbpvg6ALS/cmn2IsCi2ol
+Xnl87mb6XQtwc23ghQHTT61VxCS0Y6oJen1H6m/wAd81Z0ll1BOLTyAL4PvbHsj
+HByKJfzsDgbkzswXHTQxo162y8Nds6E8P4f1d1C+tEn+2A2+5geyho1KzQ123yf
qlh1Kpkiaviw7VMlHjiJLa2js4aAJjBqayCDg0uYEuBMcvrnSXXgDijMW0UFMLkH
7vRkPWXBYD569eiT3QW78Oh6y+HBBKlKRX4y+hllpk4+2xCnYAqKnXN36SGs5Hv3
AmiMkZ3F/G687VHntSJzuZMu2lMQ/S0jYVYTEshpwKNN9xO3UCWNyEFNshkEGu1/
zfeKUMaS1dlhLaABKG3VctP3j70TG+lSJiwJwwCuqrnHz3EhWUcm0upGE0HGz24U
VJzHkhWu8PBz84710L0v4+zOAhRfvrLPNKTkV/G59/JgVJYepb2p4yUcoOIKaayK
MqOCtSexV2A4bHnZs14LHUlVVI6ZZr88v3TyWVDGMzUfgnp8BguycqYQupbpGZM1
fDR3l0vGldr6P6qkIodwQ0Hr8CtRowgqluuZAtcNNdhZP+SuiZNwruqILSAfjvyD
T5xoOlA3lQv7lN4+OFALDWgikqzUGipncxcvcqaoLoJQc/0zR7dlkCyAsq4+0y//
X7NZQhle0SlgFp8FmG5Oi5b88GqPvLIeOvAEbHA/MdKbD8AtHv8RUp+o6Smh3K/0
Xa1IICgFdnsXNG0ywLKhra9Oc6CmKR7gz8WOSAptxute/5dOBhmVOJ9E3Hjn7awY
cN+/Zmy3UBQICHzpoYnI8pdQfQXcqwhpFOoo4Zg9npxgiBMGVhsIYGWgkYgLBMhJ
rxkJnIeprr5m0RQCNoK6ri1TGmCEUfhXsmy9GdiwhmWdOZX+0dicD7vfj6/5GfM5
J49lNp7xSCFI5xU61sjV7l6FAVUsmc0hWfKVM/g0zI9TA4sGd0F7HtcIOuC9tvzK
Cp/ct046g73BQrczkZOOH2VCnjTE7RNKXIoNddF3j0JG+2NWXEvKFQnaKsbDNHjL
d8lThHh6Q4h+iJGrvcTGvV9AJjioEHpLn7wAtVmb+GktvPNGuTKgUIOPVrm1plsy
ltaE5O/elElqYiyV0uSFYxFoZCAnDkIjzVA1c1Kr5MXYkNjKJy71SZXJjhUScd9+
UZBgCVmQuQ54JeLEehztnj/3V9+v9ghw+fmG0rhr6IVsS6BaPWwO2rdPukJF6CnE
+KnYrzgliRHvUdG/mAUQO1wVnZ6C37Fj9Bo8rbHti6CdcmPdRAGQblBzhwCiFC79
rw4GE57grkGM4JBPtDgvm5Qh1/VpPBynYSDS4d91Nxw/Z4JnlJZu39XV1fUVuaD8
ciraHwyOAg1s3HlCUQVABWpMEiJqj+XDPZ1zAG77GrAGsySNbKqBPwvOgbYdOqqC
xuwLE+lt5D8sLJs+sP5Hi1+5tPHaZHvD/5RNvV2jnzwm8rYvadkFrVLsH0zaZEd+
NxJEIhFZf4M8fCka/20y1aLkUmowmnKbfnHcsdVdEPEPHTURXsvR215XtK38qNIV
jdDDiOw6bKkL+t4CEzv0h/+9g2YyKqk9m//2ovxdBHwMlcbdo66UNNtX5yOF83aw
adOBG3kjsTsDYqyPpF9rwzQhXpIbtkonQ4FW+qah109fEDWs9YZcfCAvbY5sZAwI
bdjeAR9XSG5HuTLxYrPl1qjSzJlLlTq4IhlV798jpPAwnXTSNFbwsYQhJfrBniZL
x3kvmC6d1Uq9gt0OyRh0DRCPq90cZcLjF/N6F2OqYG6mEsIEQZDmVDZ/w8sxy6Rb
gDQt0/onX6xaJlmrlvAuNrbuW754OQLLfhI67ZBve9v7WJZJHCCu4YkI6jyXNx59
WlpAQyPV5v0lDnvBoj5Z6+2AMgM3R2Zh6lkhEm1zMa901exs5V+In7SlJ6nFlLBC
Yav1aIolG/TBBf0CQuoMKQDoPYs+VDa3g4KLaD01SdXmfpoTjLpsDQ+993DHtgtb
46ZE9EVEtp4admFsWxW2IFu+JflUq76A9Q9fzglSoUbAI/sQMXn6G1ThMEN9zTri
BzXvcmRNJWzQygG17pCiZQSuBzYRaLhApYMGeA9WrYMsuZQWDxvbfuEfNCOrOPE0
Zhyw0Vyurqo3rTR+wJBY4sMSc5aG0IY3KZUdgEugmeozRMfUtriKR6q66JTKfzRP
gutyW+et8G7gp4Z3ZRlEqIaoJaHj554x6fvWV6w4lsq6rzE871XQXht1nbBdt6yM
blT2l2T3Mu1U+cd4uW3jhnCxIvQKfydua3ijDqphLMI1zKaVuHoLzIr9S9BS9uxT
OcHNAKiqtF16wELPdHAVBc67TlYWedppwFzjLfVFwpWyIaAtTSOl/Gf4LnZf3R5c
yzDBrH3T5h7hdyL07gA/gPUvCX51mB4ai2yNKYd9GXTiJrjXSnFX7tpxmAOhu+9p
Es42sKz8HFpeXErKIG4VwCAnfV6TvWj/VthbGby2y9XO6uLXsY1ifN16/OKDZel5
sZBZtt0N1iIOy8hGwT+EfZiiXmCbp0ZdX6W4BgZERq45Q+u4aiRb/oRIrlvQUij7
UeBFveMSnookyQT0MeT+MkqJ5MhF5eXTgOz9GZvGiZpXDrSufU7P/hmDQg+1rBvH
yy+3ICbEeTcweZmGRXINsd6uDxvKCmEDQfmevaueLIaAKaiPOJXGDdR4nO0JDXtO
d8vM2WJrUQIp3Ic2mYSeNhZVHvfKQ4qtJBnypKioRDgODf3SFMNvbap6pHu3P+cj
luwCsmVnRpE8On0OduKdGRuUMmz+DszJQU8hbuHf+FwRGUryQrecvlhvp8ToHjlM
YnDPiZBLj1Mrk+yJwdHrzkUjScN8WK4eJ4Qd9EfEimqzQlZOgojBqPy7N01Ito+3
81fiXRnyZtLlonjiDyM6BtEGNF3VnvKTQX8VjyJGMyJA3QG9RHOTN6KbR1rxOTnG
srqFYHzxpDktoMOrZRUZaAIdm0kD926SKJ0TKiMz2U27RUZR1IQtbL13iiF67O95
EDjSm0hrJdZ+rxMhTmOivVXi+PZMtONUiakLvjK364xT9CiDoLOGxTxzsX0UHpGQ
04tSKkYnJIaANTueU41QB+i9GV9WrqGQs/GGHgLHM0se6T9B4IpdDgzv/M7cqawq
u7Kf3ihaF+al3EK0wpBco6mc6tx7nv9Xs22zf1eAEb4tCUE/OPQ+2XQ9lsHqXTwc
Lh3+hiCGvG6sDuPtj1Es2qC1Ev1jcWxODmM32kFN7KsH/LdG3ixKzNJfKnd91wfH
TQzAlS0C0P/Q0Fff+kMN7WQwHj//TSJeKvR8XEabVHEaW9xE1TetRib9knkNeoq8
V5VJsU0ffeYg2ulysTFtUaxW+fYPjF8AUeobEz6txE/0HgFX2bQax143iH27o7wR
eGFcAx+L1DmHX9+cvtlVubeLMb2Z6SrceNGke7LISnE36FXCkDuUFvRb0rubsd/D
JrFgR6e19YEYL5JsaL0oZxV5Kl+FjNAwKU5AtHrGNsJ2+xP1dqvoAwkgRctGUzE6
hUTUPRvdSdu1QMGQziG3TRRldCeDHbpk6N9XKI9TczCFXZYDSCrIdbjOcAfw6/d7
XmXFe8zN9mvlU/6NI0hO6xMZjMVCkmY8hJZACe/tCqjS70QtO0VSkxyns1A5rZFK
vu6tl1547O4fKytwvERnN7IdN0UmGIs1tZ1lhWBcLKipwIhGjo0nsU9zks9NdgYp
QcoIeoNkiRLvcWS31JjyWzMy5DzAOG/7HoGVSfcWRsN7kd2v7oLGrSAdYwl8kmQh
2d64wyYeydvXVaqyUKsMVtVsiZZ9KYUeH/5HbLmg06wFKApq9zlqSV5YrXpRYkDr
TBeenlFVOSF3RTyH4xk1mQj3UUQej9KPP6+cbZyhcjns+XmTiukqoHhNCSXqrQX4
e0XbAK7E3N4io0eVKpGYrpZrvSWyg1MjG0Xz01q2miyIBatQWBh0k7FaiB1OCPEh
/dJ2u1koicdaaM4tbtGkruHpRNA2dZ9xPTjBdkUx/9kPl7Dkt2atiihBkoniURjz
mjcAe1ocQAWpzosIskTfag0LG2xFhxVRj48iJuSORxzUSZmdaie04OUy+qWsQE8I
WjfVG2qaIQKY7P3q4qnQ8kPoxnvf09LLH5bI7ltzx7PC5JKjk8eiEo+nheNEm7UK
fgm5amKQv2o0v4b6r72/LZv7k+WjdpO3627SBAImy40iJhk2/X4xGHggDTWKTcOC
1S3ADh5+USh+3s+m4/HzyYzu2OPQHyN8IRn4OF6TLY2BysAB2emhgYgcnWBfR+J8
yDhnC3t0gVHXFzvEn3oiJcs8YCNgtY0wPznAzb+bwTFVhA5kasQJ/ax45U8tra89
wOTmnOYUBPAM8tbzsNdNlDUMYYSraz2PwpAMIi1Vy0i/Uq4rbUKh+z4Mz58CDRvp
4EHBRi411CVqjtZ2rdxL7HuZln5/Z+B6/RCh6l8FhS9Y7Cqsj/ynWSWKEHPWLJ6n
+GADGbXCzCJRH5juqGBIkxLAESASzlefN2waJS5zgwN8GcyILvU3eBXitwIBLMFd
LE41GBRQcG+zKR1D6DcT9POAWZJ/CEkMdAhOt5+FSJLfXt7l8Nxh/UOxDEy0Fgzv
hb+Z2lw6fbpq4kjyN0anikV0+9gvkNFi674PsudI+4Cbwk66lcSB/R6azpaA50l8
DDAazAtlLqfdx1lVln3WpoLu0OjmHsmjC5MQtT8v0XH8PTgbdK071Yqgh1/+PY3c
kkO4Q6gHnw+D5rFlnzplPw48gpgh9KCSwLcWb+xH5QNehixlD0OQdpwMzGdIgNZc
sLv5kyrNphTtBuk62fSapR6yhqzT4ZPbcXpzOhjvCGSixVV/kibWqyaxhq1ewW+R
fsoSsp6oRE+TPkdUuYIt0blvWIk8/bEBAmGvwGT7IsRwbjvIlID/gRZuC2VBqkqA
3EgrmH9mCwKJXjU7rKlwNRlA/Ni/3ocBJkKSFugBFaS48SCWaFzFF6XRqcc1Iynf
9pF/aN6I/ugIdlypllsXIFTl6sZnyxp7VLYpW1nqstQ88uGkzWcjMWgxOE8ahLEl
jkSw1sA9ViNldc6MoWpVu4aIiLAfJp3uXd5+q8KWVnchwSNQA0UfQiIpS6Xc3AuW
IKdOVwvz8m3QMurh9DTPqjBs1gdkt5kSsicbfYs5eEHrtj/CtJGOniIX1rHOjP2E
n7JnN4vpfFVctzp57A93yR0gkiIBsLsp/I6GhloFRpNpBMneWnQDPiqYrLlM/gBk
AKtk6TrNsdcNCINZJy3LH1y1mNcknydFAX7QtXGQsFcAAbfsJ+JtIFEuJibOUYCv
0JinZ927SarA6NHbH1Xul8RoMKK3t8oOUk9ckEgKEZmR4tYi4gRF68WDEE24h+Co
06zsTwaGlKNFXdjIgaPHGhfSJ1Ymuwp3u6VTYN/mK3pVlSvgkcb60UbtWtlnbnx+
bLMsQsZJ0z4Qu7of7q13x86Okj5qyzDb0UwIGOYG5aKlvVp9gZKqb17g2WAinmhg
ypM4OQN1SIxAkoGS9t6W25k1JtTZqir2DpE5r1X8+ImGYBlL5XLUZPYjrWMpuSh1
mWJHQ1akgdIZWY7WH5sNqfAQLO8Q7oQQd5T2cBoIWNvcoT8sQnZ6qGovfNIWRKMO
QPunfBNIvvArQ31DoixcSM3GpiY7Bzzn9YZLaM9uTJyYggdyjU2sWD2zVuHY6/3P
Tt45/WqHP8F83lIp/UORRihi6G6q7pkv+bTd+ncNhV04kUtXhLpVtY/GS8UK+wYJ
+XuJeCjiKKIoV6c9KU7oQHryhAsZu2qYcmoBT3Vbd5jpeywIDh8JlBEM05HBADiq
kVIC+FEelQnVcPSC7e4i6jeNRzXzQKVZzKuzqwXsV2QMeSjxq4aUViE5xTGqtUdm
3xZg9PH5k2w+rgVzYADUOCPnHkAlVbc0/ykUEfCGKCKprvn6ni3ZD19CQy/K8uda
aseOqJzyU1z6oi50i/PLw8FFJiFRrqU7Ufn4wBef/+KSt1Og9yRSziTT8mCSt7Pk
JSqM4SN584wCITVa64Fj4iwMbpv3+5Ovua3OkgFn2+H5/JkzerK3ZuFnDhyF7zs8
wd1rlRzrmebY4C6RcpnojgsGTUsfPSegx39Cz5rDZh3O9ffos1e6qJoBy7GMKE14
c/RevaFnT9BhUiHLgTFCnhsMHCnF+6qZhlLGTVFQoxE05xthOhFaCWoVoJxoHuiR
vkTeuVmVaWhnQlQ2tKnfPaX8lvUAIK3BVxywWDwR2tLzP21PEx4cS1Yb42NfZPM/
LUka0N+SB4Ro/TPdWUPMpLJ1J7+BDluy08Q60Fau/VDYYW3on+ZSDFLxcO5OtXm2
Q2v+xOpNNAKzplITVhF5Bj1hAFmjPzEzwcWTS7zcocQPrwqhbgQywr13fzTahYCK
sF0EZWL6kSJJFNeyWpF3BehMIeAYtPNpZ+AW7aftzm3RjYpD9lfF0KUNAABSpfCT
IZlRfH95sO81alNqaV2ci2m9kBKHyC0/uEvBeNAoNyKH2YvsGsFOW51E+12lA3dH
U27WOe96mll/GV7Pogqa0Mo/1RRYz+7Ujio374X51Bb0Q1geooW2v8x9uWRlqUM5
9SnFDpB9WDSCndtLLJAgql4Vs0mgPrV9otQYWr8SHTRFocL6cv0NxCw501q2N1Im
WNktpB/Rpx/br2iNTW8IY+EncoFm/hxV3SGQXfZT7bxZzQ0dTleN94yxtIGCluh2
OyI1LC5FkRluLh/aFfymahFUXgsofkx4ywuj9EyLDeJwiu4AYP3t6s+zVOs1j2lS
Res/3xE3tbsSAm9EAd9B78K7P7q1KVdwcnrVO7z5sE0O+q1COV0WBXjn+YnlcQVB
wz7a4JjMC4btG0HdaziK5ok0+0YbLvVDyYsQ/Z4JIJytDdV3pl8WVQNr3NUAbJUp
HddXV/3ECvVNDfkOPOdrL5ERZMJiZMc0LwjVhFTjkQZfPkut+ZYYfN9LkoRH0qDp
wP/Vh45bE8gAb2Q0eBnuWDWvEL95KQSvbsZ9zxsl+F/oYU/MZROiKAayzsBrm4bQ
EQt0wtIOoiARuxMW2I+cIELxmfPEwphCPjCBkqMiprs=
`pragma protect end_protected
