// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
GfodCVaeBNMxYvs5rgkmphKT7h0e+b7tgK3nzewrI5iK+idVPwJ1OH1UKzf2c8GMXlKSPelfTajH
oDK2Rf6wzjjJIaediIbiCVXPJMaRSzC3h3Zx0Y9kvG/sPcypE0ARV26cyPCRoJhkBFVzVX/3D60t
21Mkf/6W0a5FD6ZM9ofnq0BOXO7Bj7ZpkC39CLJk3BH/l+68ip3668b+kYABeqF4RVEnYEzqSkcL
0D+6knNGBBtuHmUTZEPLJB3YStnIw5fRSWL3PXZLsdGI4u00qcDrtYg/qigrrmn7jCRFyXvrTxtA
z8frvz5dK98GGsYK7UCxmcrgyJ/GJATv2OStsw==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
6fxpd4ztxa8HlewEjMBqaaFufRY1aLTxxil3A3Fbj2gj1eDW+vZI3uWvrdhOG2dfWUm4v2G4C+wk
AuNdBR1R76/n7hHvlI7e0sJN9L/d50UBLmwrXfHuXeMTUS2l9vovbJucUKspMM7Q7gImKsXJWZfJ
eIlZOUSJiHX8AUEoCd8x9IYC7o5iR7VT4G4Y5/2h1Hb6Wt00nC5drIFladefjGPWmxpKhyWQR3nj
eX6moS/J5ePwu8lA1WTFmc13njn9caj/ExnPUejYQ0rWv28ucHGQyvvC5AdHR05a7QEOZtYyYg3O
b+44T2vOzDcqEam9CR4WHOCuSrVKWQoikixJ4zbHrTfIxNPlY72tKc7HbCrC3GqTbLTV7UBlTBqu
dEgvfTBQ8DNK6vCI6bgMPYD5yywsvLbMqcs2KeLdKkkPdKyOkGRdY0L4BuaZTUH5cylPBCUxSKgm
kiVODRMmKtb74BVDymAZojAeO7sZJEHSDaJ/7bGoj8SZaF3tVyO5aAuieS6FnHbgjzN9BVlVKtfF
DuLlQmSO8+wEM4fzQKnrKe3PBf4oDIL0KtJqxtzdDIOqHw4peW/mqHmG9pW46wGKFkZxsN8/9+tI
W8xdZnPu5V3dUgIIMoVFDk39IffflkYGLqAnqBSW313FRRxaVAN42Prv60TriUW4BAv93QuTSWRn
ejoP8rOCkoRStKmGYH5UCctihevzTtnjfMGyF/dbdo2anoNPWfSU7wil2cndwLIsBYs0GMA7I74k
w448Hi2l6t4eWkjJG1avakklOeNpFEDJAlZWf8gMeb2cjJRoQipL0hGiNRu2fs1+vXmIQRQOzQyB
rioQ73njTlEBE+JnqM/r/0opfhXaLnLPwZ4q+Kq8Q8pXEsyQVngsXwWaX77eJISrWNNgUgBsXKq0
j/zVV0Vpf3ACvGQ2SgC5BGmIpOkLiEApTalLwyEqBZd/CWIQ7KyY8CmRXh3wVLiLq1IItQbyIwlr
jrdsvZxuz/Jd8BHVHwEMRtaIB4kcF/H8pAa/JZvg7gIVSFcq6HZAjIAG0cKbiJxP1ihGOqvNYdPy
W2tTgI8eHcyTaiqce/PAri1HvYAAEblhZfZdqQjL6psdRiOMOcwKSvfM+WByghp9uksA5GOYAui2
z3Oc4WJEcvIiA7ijHTLKz0UJSijQV4GP3rmW/dRY4MReX1DsHdr0HQXqnZh89rknwI+8Uzq9zcoC
ULQMjdPtPRuZI2CCbD2ZNZAFA99RHZt+Hq8wKuxzP5D1bQ8TXLu5LzO+/l0LD4pla6NosYmqykNT
8L0iu0jjbPK5Pirp6juLtOBG/+Vnu0QUqBgG7KTKNFKtrhmdB69uakaPLOSUkmvxUlwPj9j8epnB
EIg5s+43/v6NfaAJ+jTrqhGDmRKCYnObDWKeM6h4ZACTRMkWKTOv5IQdxbbtIySEI/lRTbVeu1rq
gcJc9BWBGyMa6xmW3H5h9MIzjlO/7+ijwiQCgpdbme8sHnUQGJ/at8F3u0xRIpAn9FS6B7YFtgjy
eRVDWs7TnLkRf9XAfBiPXKtL12To+eDHnx8fGFUOSkOT8yWNl9thw3iFwP+d15Nwj7ClC+DKSJ73
A8eiV6yHiF2nKzDe5X1p9y6NR4qdzRf61X6AlwaX63fZZ99djxIqoz4Jop4tCOuHSpI9GTbfpMQX
fnFOdtF/BtrwwxwEYZ95fKPIaD0SlHDDktmqA5jxfe0PtIsa2OCmsI9YTciKUGKzuDfTD0dxE5jI
L/TEbr3L49h2hTYl29RItsTk9+eqIpYJQ48iadb086IxUvG+//gFx94Zsw4ieRlyvz/xixoHeD5H
f2AHmgEBxCTXLDBttsQpPignAUCAnayfNj9Q3mOuvXz8GvvzE9m6DS1WnsS0vImQAqiZsDoYd0os
4vYG7PMQ5Icopg6+8GgmXtylPJiODDNmWd2GIgIESDgHrMfjMaPscqw9mLegRsoB3DJu6+z8LxJX
AJZtkDTBPinvZ68NBNbzURLN8e61djyAL8J8NQlezbYzqg7LR/Szp6ZbzZ+pXLpORCozEFqpYmRS
kgasgZ7O0hGK4W5P3gj+kZdhKUKbIlitwwTs0SNJY1lxNmCJaDTn+rlMZn9VmAfz/x47oVQGnhFS
HIXaNK4FxFTlPeAYH9+1RQOYQgox1HmsO0peekJ3OqK0s8YKDlqHqzeklbgDlACsuQRa6ORHbilK
AiYY0ecs3Wo6pAg/B4xeoyEZEMO0ebGeoisKBP+7RNxWKmbzLlZhTHWfA3N2DuQv7NPlPw1MQkhE
dzvQIdJMSCQhfB7CNEjHho5W9ySYhl8fU2XXRdrmZnU60wvCjEGcJndAt70chd2m+1KCL3J7Q9Bl
qfcaSY+nki0gRqf8YwCjJA2h1pyMome8ARI+DgBnhnrWs+E7vjYFoKQ04Zc3lEkzaee6AVLPTx5g
VBdAbaQ3KPbDqF4ITcDZEtmYdJba2rfIVvdmC0oe4PLA5NUSBhlsOsBskF+5va9gTZDGFw3H9e7/
NMGDtmrFXSs7eTqejMCQB8VYo9L0v4ZdeQsoNxkAGYJ37m5+TV9vAYX093A+3dYClpuHhk2uO/aW
38ADLleA8DXB9Gr2TNAoPBo5BCwzMBDR957Fs4WoCHVTO13ulRrBldtw/vfCgw8lDDut3cATfOKX
Wj4smVrgKyQe6qzT0NIT0Xo8TxtGVh0GP/xn5Tmky98O2l+/VYRyxzovHmSmtP0hiYvsDGbIYhla
HoNM4POPsTZmWd4de1wjn/Pc7Ojy/MEfg1zMgXUiN/1BW/CZfvcv2K8vQcsk0WpT6MBnpfjGl+0O
cWZPcT48CWlCcaSTwziqDEAzI7u8wkD9MF2EiFeL+qxKhhFT5ae5juynLxFbdLspPX2MtoOpAORt
kuI2KH/aTrTrW38Io5hl7tXeiQBc/X/VpFDnky7LT3eKLZSto0M7Q7ZyRvI5iKPJiIdHwwm1eYWe
V9Fa4SYU/uL9bhKmqLS1UU3mDSpTlGj5nSyBVuvstw3/rx4aMih32/1josqVnJ0illOaMMFsJvhT
MrXvWLuyuRk7+6OD07GJdc+nscF7Wh4mrTBTGJYt2tlSrv8fxmPWWexuIIeuIw4BL+q4SqJ9ysWn
rR90bvXhaZSAHKAxwDVrUGTe+HUlQwxsyExsb/P8TZcSbVjbRe7B+Sxk/thTcBw8tSaDvAh+sBJ5
5nV6V1jbnQamcpsc0JLQ+pmSn6tqSWpzBIz3ryrQq43upISuZprzAn/xq2z2aMq5TH41QdTvkZAN
4zVIrs0EUdCSKZIlMJJ+n34KVTQxx9Jc0ymF7builmFaqKwelwQUNyR9w6T2WnXl4p4Cthy95Wi1
qCtWmCj4y4WV08QhOoL43pKM+ZYSne56hTWVjQxiX7rq81fJxR9CqGshOAWuX4xf/iiyV+pkeiOS
XSavhFFVM6PF/iB28a/Oov6aGue3tGsMFwRivBePHUCwsdpzfIlcsr69Q5cDrlmxmLjLV5m39Gwp
vTYA1qPAl+fc6ESqGltWMmbhQdBKaPh4uYfkhw/6f97DHUZ4pZfW5k17sqzW2fEsCD/ndUoVwuB6
sUVplXyrpDcimfMetlvfUcGFbPmOTkCvemYRdPvhZlry7SgiOjykMV25BMgy92REz7CYINUVFmuv
QbdP7TUR5IVtCNoTXy90b+zD6QVh/D1GRCRv1DtYQj8MvTv8cjrp1gb0r6wH/z6r6e42FtQQqFUH
b9TkkyyXCbcLdEbplBklbiT3FUfy16bp4D+JaR2SUlvR5hBQGaUyTky47BKDvgUTScc7LZ8HIxUb
Gxi2Gben4VFSdwxvhZmGlcrT8KyuGZS6gsuYg2YytKnLr3jdlengCvduGJidzMdRMsVraIqwjJk1
qqrF3XxPRPSorD6CqW3caI8g9Hn1nWyJSK9EZaiyP3KjbKp8W16Z6X2C3lqqjKXluPtLzi7+pqs3
YqlsgZfaAN4ATAVFGDH65zxAeT+Co8po8tuVcUCaqlKXIpC+ZsrOZ+gp2tLjAhKB8HnaaTMCGwwP
Sn5SKXqyrET1WLHthT2UAciGBL+JdQ5yDUX0CLtn48Vxu/YDlaxSeEjguCFUkxoH0N+8T+TPoc6H
Snf0TA9YDvYfpflhe5WWtcZUJWxwsF2XmxpDUInsSH/YC56JpZGuoEsAdd+OkXoiRx6nEfUuuylE
cxicW50FN8DYfB0PsAkxYLtNL+g45FTNH7LNiCo4tJfXKLw636pRU89TEyDXLHAt4LoWSTX0Ct4w
8vNy3vwkpogoRG7mnhj2oZe6UpNZzzDfQPA2O8twjXqmX71Wpwr55I+iEKadzYwNP7eU+abjzr9/
SvDiWuREro83FQypyxDoRiUAHsi6UFoZMHILVX1FObl7Gmwxmz/a1d5J9JEL2Xuck3GlwELKH5If
ioNpJoJe1aVkCEt2YDAFrUVJU3bFQ5ajq+Q9S7wa1Zn4WFIXfK0iWQ4kM2k3Yoo6U+B/L+kPlfa+
BiF7CA8QbENP72N8eaXYLNnCzAGh2Fnwlb/XwdJ/kaMq4HOkqnqTVR9+NhcP2GBp/Rsg2XiJclIk
9NS2VbO07g3E007r6S1NwIYvW91a6Qmy0fmn6mHYnbzR/JTeLfbDtrVpsln7TXrpKhyAPbP+X+i7
Vzx+zrdpkxwjfYGeZNLGUk28xudxpMGufwClIj6JaavASOs8OMv4tPKa0WjzuSs2+St4t8daPwz4
PwGflrk2DnBpejRHjwJiPEbxqMkKK80rxEETrbmieKXzyPwixjSEtf+3lz/0iCrxyxCR9DMq8ioU
rNHRuPN2GH/l0HXdtNIY6n/vrZuxpR0sb8RHSymwWpzVJfRfkC8zKBu2XvIUk5fjmWJIwiVzfqGq
RC4CqMVV0LPm3eS/mr8bhkQh+xIh033XaXEbE0Cs3n7SfzhJkuvQk5pOUyA6FyOSr5XtW1VjGY5d
mA1s67JwJGwQqurSyW+zTUJWeCyboTnzkHiLsw4hXbryPd4aHBD04GzDLs76kc0PDBJCKoztprAy
q6Xta79M4lua3m28YkcMqc+f5sWQZ98KaL2XgvByeBVKMBwm8Iyz6zrawppUho7qKwZnPnIflS1F
vQStj+yLpVZ3cghPxhILVehrBMSr3Gy6ZpFX0UW+hi8whUE2sVPo8hftS+IRR041nKgfeMN8wG8C
2/f5p7pzunJ9oVkeHEc4kyw3XXO6U/PrszkwkcFJAccgd496U36sbCqIgT3IDSa8DJVe5IBTWCV/
yZ7XPH972WEHwaFmyTGyOn3j/JAHQ7NP9vZxT5rzS6G+GRuxE3ztT0hcfGD0E/eEQmhBhdzJGuWN
2lm/KUuBL8cCxGyog/KnJO1B+6/HqizHs45LChSexdPhut+J5xtQ1hG3uDUTUL2keyGO4LuolOxe
8QrR+w/lR2GOPmnfFfyQDzOGPdqCf3G4GR8jNfshtovAmcuy++h8OhvfZo0Bnzf/HvwWlO7WkyzQ
wKH0nLFoZhjHPoCyX6RcptmEr9JWja1ccFkEvbWOmTH0hONwoiVZTPd+Q5K4jgwxyDlZSrCccA/u
WFmfbIaIl7BRV7q5EUs9lKvVN7ZZA7aUwT5V6gJmiJGmfoZnFKxYnREeeS2nQ6RUQ6R2JuQP47wd
msJEb5i9vjVpFaXWrguVYQ881EVOIBCAdvWRH2rRKAtmu9w49G9RHFeZ7Cg9ZpfMH+LmHKRo/ITK
R+k83vASXg17wNC4vEsnTekD4GT5N1c0etC3C9LVU8EMU86cxchPuNv5dmmnb9zMUrWB3bU5ig/f
I7M6iy4yYdCy58eucB+ltFnGl0TA4ppSzyHcCxE3QbmErzMFiYinsVQf8jcjUI6feqsGw569Td44
WgDbfHXJpKUmduERwsgd8hZi+rfc5wg/BnRmwKVs6/HqZfKXr7Rt8QDO7boYqGVZXF1+1iG7kuXD
VJz5gCxo+VbIPREKf1c1UjwciLfGax463jola9cU6Y6xBiMgLj3sGwWAQe99fGSYaszkdQTun2ZK
2uUHMfn22qeo/gOpJXx2EB8GkOto57C2Z7uP5d7FZc56MvBPW8CAV4wV1RND+Nov8XzA1cz6WoC0
fdKDV2c0kww/bRodc5NhU8K2v/wD6Gc6gK5KDh6HfC/ftsxaRvN9q0ZCA1zESNw5LdNDYpSGh2TY
WdSLIV4XrmnuXLXyTOB0s69mEqhoBhcyeQzlvVdTHpPjvKESwVNl5iZ3FpkJagvO5JrWpwur3pu5
lVzI1IBIiSxIWJBzr7axeAbddOYURUEpcH4/P6cmzLxAGTzDWkj6EDsewmH67OLuLbjFWLqACNso
QgC/ZCY7KQ6z+1/ko5/NaOfygNOSUrMiUk61mZpvuHg5SLT3wCg41gmE0dRe+5yhMC8xl1YpMLFp
yGr1W7iLXL4PTPihjxMyxRnl7t2fF+dUuZqgimkAbIyXqV8KAR/K5fmP0CbF3k1u7WL9F1/ns5wb
+fHAy9O++RyXhVlI7xXc5PFQsomjr6ZVWtOZ3Zvgh7sgxtPyR6VvXwGdGsHYePUE7htObw/MoqH9
iXRDPX1bb8G8fBow+TVa/TdF/VrHpEBOhQT1S9Qx/4LTVAZQMa1Hgz2sUKTl4meAa8TAGx2WwtsF
CZElc6txtl6J2fwdr1py7rVU+hMRIQ7G2ezd31JqdpJW9XKbrnl3yOHi+aTCROXxh5lV89Udb1xy
ubNuK59nPBKiN0JYJWwF+RqXrFUKqUaEF6PJNnFeEkoAX0M1NzV4u0p46Z494TQPWuTRJ68JkZ7q
pT9RIZph8X4Nw2bdsY43ndCvM8sKMNvoN45jAS8GdD/s2ewGhyQ5aiBHnIXkDr8rQxAf5mrL5SFe
e3uS9QKl8cYahSWX9rMtQKWkKfNjyoNz76xmMRA87YCfimlcEpeZb9zZgpR8RygsacHDk6Z7CET5
AK2fABzqVyOJs2cF+B/QDrnxkPddQ1miV5mOw8mFvIGu4Ahin8nLDf+++xnGhpeDy20FLYWeMA1O
BSM2H601nm7pjeZUJcb+RS0MosMmJhYV9QZ79hcs/r8QCQZBRKvb4GXjRNz6WBccZQ1/V9YHvIu8
IICaQgaaxavVzfo1E0llEd77+/kVuZh9X5dFNosAOfg0c58lbEY2WzUui4GhOOOgk4YBPRl6J/B/
1mzVhJD4tMe7pW3jDDSGWk3dDHRxXSr7nU8YW0TpmIFYbGKf3z2qHIgYyH0aneo3fNhR50QtvPyK
cpnHK+Lccc87UjfQAqvtc2lKE6sN9XNMGtoTfMiaVi+OVRKuEtCWoU1DVNqS6UTLlY3xASJhdoD8
sVeBDcIUcxUSuF5J+beQAok1niBQFFKxQnfWhAxKaKFICztf+YH243WtvRq/Po+ky0CjKNZKZPXl
AIUsf+hwc5x8RlHa5Y0xQmbfTKpeZhWAcQJRUkpMW89UQFcMBnxBpno3apeFmzYyiPURnnUdgkvC
C05pQ8r1d+40L1wN4Z0KMiT/4IEkGAMctySQ+5PnG++lTFuxY6arNOEb2t6BKXssxKsUg/Fj7yGn
/BGHhShvhtDo8ik5xPqqrlD1TG/Ma4bphGYjwQF8OELpa7e9R5L52Zwg/aBI2h334iU8TxoevDCj
qqM7saYO4hukMudDhoXTHQXgdUX7UWR8DoMmEQn6DkegHoX5zGzTt0wF+YAqgEfUVOgrK8IsD5tX
YGN/4nXf48vV8NQ9dMA3TuspuHk415v4JH+JIyC3JBstpXqctsf4AIZx90pZixCroJmGIaZ93DhT
rnHIhRwuWVJSwlp7vYRv7yl478X6jFrEHTewnNKue+igVlVjWXUMV7XUZn2BRSo+OYms+8hvsqkG
5FvtUqSaC1tKhlTj2Tfwk6l2DMXJpBQCmZKOfNxv8G1q6jX4JHfD3OWfoic/W9COFvLVLN+49BeA
JjpeLcbzTt51M2hdJEbxUOcpniiOAryWxs5yLo5fjwM/GjY5tNIS5+1XY/QlgmaB1Ef60oiUgXrd
1BaBsSeYkcKfSInWID8C4GZBoAWYZOYOuEWyun1h3jKcbXkgEBJaGJD1MrOXkY9PEcvWN+wqfYUy
cQJS96cfu9CHqw1UdhD9DkkPOmxFkNwfI7BTfI+HkpXY/O2lQ4F/ZQb+1kT+HiBBcosy5eenjNL4
r8i8FqZVrHGtNlW8isZVkloajZZy4lDoZxg+kzZGOlSwSEDOph+ev6zEMe4QdOQG5gFgrwWkSpZ8
LqSXeFi/XFiGKaUfyXKuRocjmIuzCXVYjVKu9NvzKUk1PPghnfbyV1xzFMe9jQG9b28gXg99uk5t
nqKCJEY6cwBGpwcdJdiU7/7BpJtueU7DrIGuoaHxf0REgz5LxXpXJCi2QoUgB3/j0ixK3qcqIBAu
GvX9TCE21dIL18p/SCfRRVaVAeWcJRCYIsCsmXd71G+dophSaRKENzD+M4bsQvONKqujRNjq4n0L
yfrT6o6X6btcZ+N+PEPHoRo4D5SXWfh7vBeJl7Js1+Ke0E1bdMaJI6adui/Npr0qp5LhYJtrvEWI
BGTcYXFPB+mXgg4Un/1vCmGS6Qulvqv/hriZei2wo+X9BGZbdDBZErGeZbtORkoOJLPabinjAuzX
Rcb78J7uh2KMqZ/gp/2RoG3hXGP0cP2eBdTUasSY/gj2epPUDuRAT52pno6ElWQOL1eHJsSzNBzZ
rWj/w0PiSGP2ZwypYxV0BpdysnRpVZI3iYS2iFFWs5HBkXvbdY2ZKigj49NfXFUEQqxFXz+z6nvX
G1O3duP3yx+rq0/sXSggwxGMZspNEvTNoASEMqCaEKkkAXDXoukiWuTxVlK/pWT9iFDaZYGP45lZ
VZGoQuvPIWnEcBhp6ZrpM1S+npW6+SLnGFU26n6Wtvig2jLGtn/1ffxoqLDOe/caYoVjqWFJsvXP
/xpYkE0jbxh0zAZ9qsrEyF3pQkENTeZy7i2etKWjPtKV2RE+rzEUyf0CYrIZ/yXY7XtPAqJ6yhce
lFMhGA/LWIDWyn6ltpas64xVK9GqT8vQfRQBLIwnUwZJidQxupFW7oI/GasBiJAt1JKzA41NE8GQ
oa4UCyBMsKDL4Sp/bHOc6MZ3MPNBeSg09ExRjo9p36I3+GSgMlEWWN0kDa2ohDgHS1aicTzDc1JC
hWyTZcsEaEhDGezmGNaGBMQwt1EuL/KguXxmxYDnXnMGgSiDIHm9UGJt3ae7el1r6QYejsQAd7yo
Orz2Z9tGrAqoxjb17Oqy5wssEBjKkfVQqkznGVCP3BB4koyjiP+FMcyxoMDAMg42sEzw5dbqrRow
bShb/1KbMEwmefDTiKOXo3E4goI8dcJRNWHHEPHA7707aiTSqP4IKZCzahQ7BXlmMlVirr7AbOs3
pbh2InJadYCOFksEDRpvFlHqSZJCUfPC2QHEKRN/Bmx1n2mCylZsxgqTK5CqFa3CJhtLrSf14Kdl
JJIPaVSNjgDcyFA+Cz1Ftg/FOlCYCahlo6ww+9NYxkJ6OaEKXc1Fu3LD2qObOajc3vrcTwLPdeVS
9MmWQFimgDGT917ghCpCH75jroQ4SJ0G5wZq3CB/ckfDgt4a+51pmcIpmb4nt8o7/BRLtURAMt00
ufG2gV1oK1eBwynA0yE0bYdn1OH/QEA0ijCsIy13tEuKFx1RXhA6ya9v1nmpmu6ylTZhfloXC5Yb
WC/NbsDYa298qWd8vzXpuLSMFAt9bt2jjzcjV5s7xMPQIfWIQP2wI6oMSqwXIdwJ20womLRljifS
CueD8x0+tC5bbakK4kesxgp3IMHjJQreyR7nBu6lNQx+d1H7KT7VVMrnbMljN2Is0rmxHSFDTYAm
VuU7/bRaY8fqyv+LLqirwPosEPWqzpBCDEj+GZhrSY41vRgZPotYf/hhgfOioBzAYlV17fygTsZa
+Qre/vhUItWrm6Q5f6pjXpGRITVlebchq2smJzcEnfOTi/vUOfdFeBpF8FHvJ2LDxvKzZOunRcyA
LLjPC+g=
`pragma protect end_protected
