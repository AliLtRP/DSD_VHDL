// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:37:12 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
eg0MPUNKH1j/smM+PT1vp1qB9ZDRLJJwjOW3qKVnA3kmd0P0gzGM/S/ZUXJYeh97
yMfCF+jqSU4XCjKRyJoMKn+d8GxuLXXwVfl68hGKlEs2I9W/JyVGT2vilr5+b/RY
y5FmR5WgLE1iaCD4c9bHNOGfTNRLoFbtz3Lzv6M8ilY=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 13856)
jJ9xq4jmPNMXkZsYrj/rtP0ZKfqXvNs1P2yu1Yv77WPXqENOVB9y9iYmLY3He6qD
Pvrfzj9fLChXblnWhHcf7rHJnKtqjPIFwPMEDqPgDlHCEohNXKGRhKCGgZwXpMyH
5+P9bRv5vcoqWmSTUYC0vCTzxiMgKeImtkWwrlDbOg6odMV3N+xyWelWA2hvD5fm
A399jEjfJ0CDBOZF7fadmFYJvjGTuM5eFrCCgTsApC63qezreWTGyNKlQ/7yyLDd
jQEUtT9ruYipkQwt0jWUq7Ir9Vq7yZrXhbR1+V121ELyoq4/+NBmax4j9keypm/F
Hl86Yb9K4xHwteGldab6QKCiRzqkvbHiVABVsX6mkMHk5jreQpRt8sSrvdzgkxVL
F1bKbcHMla+BFVzo068H14NBX0ngpQvlD8JGU673DD5MCymnYqouuyXM+7Wx7gPh
k0pBMPWr3u7p71DbEsC9TvVuHLATn8Mf9KfCjlxHaQRi2I9SDEjPUIu4LY3a0bXw
tFqEE/ey0PXrpCcIElG2zB0epP4z5PyEqgM03me5OaU4EZLImlNyOPMR6MNU5cxW
inJxmDcg/Yyo7wjN1buBbtEmVvT6fjAQCBmw4UYGNWmDCKpq5G9K6a2LVIJfmNw2
9SLPvU81gJBCS8nZrUncZKJWjfjkUFcvBLYIBtCdLXKJp1nsr8wwK+RvCnyFT+2+
atcQX2zoDf16fyvdqvwZ9tJRRukJi/mC+RuicOJQ3NJ4Iy+/L7fdUaz6LNyqYToP
owFK+nCVlzGfmOti3rg+hWlyJsvSDkM/jgdLoeQud57m6hcuBFkkDkTDhTXlZXE2
ploYnv7FGmjMTI6Yl0ZoqOwzP3w0jzoTpAw3yVPhNTBLkwfnGdey5KEj1INvIZCz
K+I45hF/TdOqPlnbakqXrTWz7S5M8Fn9iycUJmGfrVf3zbmWjA4n9ZdZ3yOCgCE4
W0tS7rFtZBAvMJXL9HSImHOlR+p5NAAJSrA52STdceQGEvBdckLc1VhmPu5OgHs/
CLaso2TRhWAyzM+D5QndqoUSALW9VTaLrmO9/ZN9BoYDp+umeynDBr68Cy4ImSI5
iSwcj+Lm2++CJjGG0g4K6wt8fwKI2NOlT04/hJeWnJUOfCJtLZv9COwR9RVXk6R8
S61mK/FrB+zFoJzhRizPF+KlsJ1l7Xa48BGkQsSE5gVU6RHNwHD2IIB0mssQMWvD
lRiih8ijGKMmvYmxNPPJJlukBVpIz0ZRwE+KGyxss4wawodKDmQhBkIz7zf4G0i2
GLCJtngslyTV5dk/8VVmg1pmmeDWQ/swqlwiZ8ybkAcmtvDpAEEjGfEext0YjZSz
cEbRiRG/hBTktCBMM0suxzXRv9/d8QpY4jDcuZg977CbOG7rHvkZnzzjlPM7ugp1
0akHqk+ACHchJlrLOrrg3qad01CNLXavJNN6wgVgzDbLgUDzW6yPuEhE1WAENMSo
EJtlINgSj9AMtjovAe8TvftmyZ3I3dkp4W0phatJp+rHXyBIXJS+5cNwCsORdrgZ
B6UFm7pa1dtYF/gS2VoiP3SCf1yWkN1y4ZueCIHrhH7+KUsPoJbL1DpHjQShlldl
01KkYifAFIif1Lw0Te1oVYM7zGT43WGZuakn7QvP/umEDgSLWt4LPskcCC8uadba
wly0w2A6zVAZxDxZWlzEIdCM1fel24Xm7ixFD1Jt3kCoHhU9cfzDOShmRIETfzat
w9Yb0DJgjo+va0AQH7Sd83EBP4j3Y2Xn/W4sdbjbOSpudPFLkmy2/zMt7XhiICV2
Pnyn71oxWPsr8fE8EvdtMJdRDTut0HH7oVVJI63uUT3S40ItgM9sbeL6OavEOFRD
HGvlX3/cGhlBXX8fCXLyJroi2WyMQtcWNEcDUZki7gdjsMbNTRpDuji1NPCRa4ty
WHPkeTfqD/g5x3ZJLXlXOS79sTUpFzRJvavwo+sU9mRhuaT8wC2p/F5eATRvHufR
zYRkhmnecJpzSav43/9pxI6+pe1h8w38bb+HP54WvjoOqxfoHDlEdmsACvVSr89T
hsdDyDFKRqihCH27/dGReRc9X7wVpmkAhujxFijMUfRjarUngJJ8at4YtSDzTO3f
YxgG1NxsjA2g2grPotgrWSfgp59PpydXJA1SmWy60ekBOHTyfW6LMBnsvfLsbivL
QxK0owlxR/W0wO74Go8+quJ4VVzf6iRB+ocdT3Eug3uCMnYV6yjiBulVf/2yKhJY
tVnCOnGNqpVSZc1LxWqC1B1YimOtgGrzqbPlOnEuk+97awG8Wbqk8a/HrB2o7apS
7HNmPEHOMkpLAoT9J8HufeFgJnJYx1Fl5zpdXqDQG4gW1FA7eT/VYxScFQY00BVf
fl2aqxlTZD6d68z0SvqZCT1W9Kp84aihudut8U6zmB3cXNO/4f9KH4cqxbhXw/Py
/ex6OHqdl3BxT4tKeVH4QdwVHyszE5mU34cSOPkPtqUXJ+V7s1SC2EmdELPG6iYO
fV+MzNRBTaSMrIcjcsD5fcYqPn9oUA4ab0sp7tXmnQR1W59asqa7b/M5yakW+VIO
eofNGD4xs+vTzN4CiZpPG33buHTXHOlHpkztTEEa4CDndPGvHbNax9BIbbX2VipS
+7cK8nsi3mdTg32nNAQr5KbAIQTOJ0FxvkP5jmujiQCKzb7d/xe5Mm5PQMha8F2B
iYeDRPoQu9xZTSi2YxTY84tBtaMDXBdYg3yO5Xqn/YBJVww0CJ0QHDreKXs8czlS
3OrW8SkVq422KJCBXjyeiNxdttzirgVfTmiIZFXWJgJeZULkI2OPKVEV5lBGfrf4
oh8e1JRRDPV0icUoxGyRc5mqrtKFWP7mVU3CuAiT2APwI/H4FwrEhWP6diwl8m4h
yzX9tlh/L3rGVrOr3/R8fjRs6KOIrgfjArp/wVR/83skSK6SWWr7RFxYbIlQ+iiJ
oYEllHM9IUEKGdSAdtFhT+gkKZfRklLZyyK9rnbJLf+IXUJryPNjASC4trGiEI13
GXBAvE4RJoYH4ZaApSokXrYe66X6qvEaesFd/XFWAxAZWdCFzji31xTKINp2YiEv
tN6Gh4QJ6vKjRR5u7S8SA+osJbvmlmBCVISx6v3iQGOroqrT8qqKTm8QAseIbn80
+V/bDjK94S7iwmA/FvwIC0zvH/P9O7YfQ5ldlacVkw05SBkZsvaNgr4FaR7n0Y3o
4jEXuVj80mg5xLBIKAmjgQAWeiaNsPcEVdAbE/ZZyHEnqdPDLkaBmMTLYVOTxrSp
sKQNwe7HQOhwxaLdlXxi+eJxVRUZD7onJHAenIY2ikZyw4FiuXAXurcXLCBj8Wzx
twYNUTDkjUt3xl3GVM7o16mE0ZN3+b4WEHw1ji46WbKMlARJ4/Rhrg+Lwg6qRghh
iiEOIICezG8wWKytQxHI+mdCFTeoOycctxW9KeRZQbtDtE+k0TmxBtiQtDuHifcN
g4q80Tl6qsQWckfa2U5HqVTkyg3WlNWVeBML6qERYQwr/gbRAa+uiSdKuTim1qi/
ODHURUlVIHCYaiPYLVIp8B6bL7a4L9SZluzirmLmyU2A4VPxAsvdp4DIrE4IlBhd
qCItYQsrB7gihq/5PtBEvp6wr3ZkDM1Ed2olQK3zMRfM0GLnRc4SKSc/53Uhwi//
fT+ezSWEk5nF1cZj0MxApDZ6bOe8PC8Nu9KLmJ+GaNhjp8OHUHAHGWOfgGlmTUmP
9HIzD4bugdr7a5Ywc8VphrzUcRp4ZyfjpwIY1GNDO/BZqQf14Y/JmluQBNC8432Z
ZfiJR7/g7aiUTPuEwxcYbh93laaZOSnxcouWkXaTp8qTDdUfVAVQB0tGios1aEfB
RTthoxHLNeFynaYQcDre0S+p5d5ZnfXY6iysrr5+SffwNBmSpwouNlslknfWZzqa
mGDNX4ZEEWfkikGKZEm8LEv3hFjS7T89RAhNJoTtWqAfRJYLQEKxJpPGWWjMswsv
mAYZWCCCMFvwEcQ1cqIc/6v0whmHI40dEw6NhfKfZCc+I4EQC4DbLKb5MV9KtJfw
Hse932kQ8bWMqOq6j5VjA2E2gsUkybxpK3xmIVheImsBaa6qWlMYO7bB7JAz4/qd
1/Eq+pHIcjknpZKmb9HKQBSu924jtpTIF+vWPEC6vp6fNR+PZMZljR0r42N92csI
lCGYyFgyNI/uu1+5nYtr8NrTLfF2ANR38gLqwdCXDr7opaFv1mcrD15+Oz0h+ld2
/HRUyLjdt+AMH5KfUPP89b+8CJUZI5ykCAeQfyom68Cm3mB0jxEJdpdBxRxpo9xr
9N3k0zTxesPD0t0IxXwjttaC5G2Oh5CgWqHqKZ3cRlA13bDCzG3XNO3RWtxZjQgu
aU6RXynEiCqD0pOJrlOttqyZktW4LGlnUlOQs0Wk3TeZvNYTMggURKQcK0vXm4u6
6iN27U7FmfdxHoLT7prGiMlRZeupGL/kLbRnu1M1wriLyQ2KKPo5dlGdukUoI3Is
WSMpu3a8zoArl6BnxQe5exBiyIIctDRLgyuMDH5Sc5wZlljoMtLUozifUFXJiVnI
01828uwHSfwnsTt3e7Mz0gkt6l+ZC+dNJnuL+ibxhMx05tSEI/trBopnVm8xiune
fV46s/u+BFYp73oMaTrdx6fm1qM3D/7esIgud1Gsz+xp3bpcHXidi7oOKPaIWDf7
ElnBNAmlrRUx9ehfBOaGxDFEei1HTTJpjqFXzw3Sk2Wce+0jtno+mxns+wwzkC3K
hUJLh9YzOdFOpvcCdekA4X5isrGVV2FLz7JRdQ1qByx4WdwsFOT03dDCvAmzn0RM
eC35oAUyQxDJhbb0tL2lEKPaRGzltLk1yPdm1pWjjIn9MtizuKNouP40vfPIGS7u
XkpumQmYa6wd5Sy+z7R5fPL9xzlb/YsAbXXUBazDmlZSCKVQUd9CQGBJhoufJT6M
HRZ8ALRRj2XrduPM9ukVxj2Xa8TOqqmodvzGzZWpD4ZEKr4xD7uNCmwepVaAYhgx
D2QUQjFoaHVgMkTp6+8PF20OIYwCOitSh7PCOn0THY/01zn8TaScmZKbDXz7Jvgm
TS/ATClh1wcAaBRVKi0YqdmqGsHMMwUWYybeWdIP26w34c4uGyOIrDgQcdnq05HC
oCMtkIftL6ULPjLvE3oh4bjDxCTnMeh8Wwzo4t/8LA0+BkEwhL064Qvy10sr5orv
RTBE9EpqsO4KbsD6mPbkYAcf7poMwaSaWRCyyryHBzBGsugUVl8cRgv1yklt+77Z
wwmtTkNmjJR5w+9q/Tl3tqRCyKL0X/a4PD6yOMNveXn+q0TqRgi+PCOcRfI6+6M2
xm+tdYul6TndmSc7mSBl075LXmM8a2Nb14yNTggjZ5/4y8VlD64qcjvgNDEZyX8S
/FJw/qJByOgvaF94vUqKN8AVtyJ/uhBiwtQvfb/beNAZIgDNKcxlwxcDrasyMeQA
3i64IdI4MpsQAuUAn558hEcjEYrnJM2VorxRPOpJXbhBir9lSq7GGxiWyRqQS9bF
jdXaTZRDFtm1+l19vMmu79PeHH/4kevOOwiviMBGhNNUtaZZIhztor+TEwD8ZDTr
usRH52r7SoaBTz8X0hz2iYHL++8ga2D8h1fGwsVS6JQq36zvTJDARwxu7RjNVuba
zppZYMW8iZXaNejfa/eMhP+GUrsFdD4bnujzUS8R1P/Rt6sHzb+0NIgnyKUTTtnP
ZFMpsmLsiq4N2yZFV7vWFq3pY/be+HGysTT6xFuVwLM/phr+1CRqZn2YDRvVOv7Q
hbB9BshCdAdbme1aWKdy/RYnIlem2oO4tuaTCV1RyNnzSoE8WaWsT8875k/W5qZP
jXgzKKH52iloKZVYsXS2rcvV++CR87FlyXo/0PMCYt0jGoyPdf348DH01WkPYUc/
B39ujXE0MnQpzw2QClXtBSVlzqGyA0VRrWQFDjAPE9J3HjPIqLRudBINhEkxnsoz
X6KNwftev8yj008kfSHNOUxv/NbqKoT6ZdnULLU7YX0YH71lKRdr/RCLeytsJGsE
yBjLcFlNOneipowsklC5+kkHAbF6sf6QJwa/mEym14eTmH55wtEMUbs2Hrx0odvC
3/QSrQzRRxMPPVNU60S5v/kqgE1WRDF1Ns6TuH5V3Z3NWnpjv/26LgVtvgYlZToN
FI7+7aClfMcxf3CLHYEyFh0FnKGpewvijY7/1YEUVAKnrUjp3NdiNXQejpa8bzn4
ns7AhukmZZXnmYESggn6MswEj83i0ieYGQhBBve3zBuh4uC1MniPiEpPgP4y2cKf
mG9aHrBzxFGYHfrPSLUbJUXXjQTSI5vP5j9yZ/Qf+ZUKCotzJ5TVQOgprmBxCFRS
kIIKMqBbzsjM0VKkvFGw/+8uW/zQALaDzT3RvAavl5q1On9AZAyo7dUm7AAADqQ3
L37jBlvQ6vRHdm7MmZ+u6bcvoj+Y2Fg0+0njcFuew9F9AykDtFL9nkW+8sK0pvcp
AJmm3ozEEZeiQaRB6T8VyqPXiGRB9/NRk6xyiqcLJXfOsdtVcnSxVc8FujSLUGKm
9zHCsjlS5UupJ137C4p2/+OTHYpWCZuVkhulhPSuonqtrqIcxfZj8Ssowpfm0uDw
RTcD5IftQiS2qRehmUGxp0kbt30ebNoG7m4NIAlgaqOAtgNwSNSMbpXzEtsz/87X
uNtO6+WqX1Vi6Yqq+cUufrNmbxGq0Kp21K9ZITBvjKf0OFHCGXDM6yiKSDNKu4Zu
mTppNFrQt/3d7foD1nYPgX2ztWMnjRQCarGz4RFcFRrOgPKzYv4JG3+KolGh0m0f
ZPxfpqE3wYQt21Bx4JyRs7gsN5YZJFtbpkxwaD9SeTthmpQYDmNyt6pL6+v94mFs
XkrJheDu5BNxxoybzKj3XOJakNO3OU1EF+5mwUPgzpS183E0ykIfxYn+scStClJC
pPu16iyHKN27tDZNSJsJpr0pWrjqsycxa6uUHdbm7tDihdUxsIO2Wr1IORkDG7xz
d//+EMmd1ngVkiWbCvxGvXK55ZRvBBdrfBxLDacse9RfaS/yi2A9SDVqsBrIvDft
6uqfsjHF2ximxKMq8K5HJ9LmlFf3YEkmidO+5hbR/stokDCQA+1mnyy6CDxVIFdk
EUtD7FRH7rqduIF0+eD4rmRvida+Vxy30w0HR3X2XT3Z+1JBfnrGpDkKRfakoC5O
blDkPbMdJ+xkRsqvlrW8kMfQeGNKZbrmHlh8CDpN/ORIemNKTd6pFASVl4sCxHWb
hIjOs1MWlCZZliwr5g6/ulT11VUPWcC3pJbMA1jiHSvIIZc0vQESCwaQHsTTghHT
Lh5hTkDm6SD4rxyU/pJsojRQN/OTVCIlRi6XJieSS5qtLqQILlwsj/Ovr69To8Bl
LYoXEL2IjWuP4/C07b+LOBwGI3CSRe2kTEiG792w1T13wHTeXAUeEk8N5NwfT55r
VAMG0kTRC6ngneBJki6RnjF3dg2PFrTECSs8P7TrOVpDHAqRfZpRiVotnjIT65TK
rE+iTK8QcnZYxO10cuqd6k0spbQ75kgviZtIqO3keuhRUEyMdS/S+RBC3iTJsqzC
SwoinaR3eZOfwKk32d7M/wP40ss9IyxTH3SMu8iz9pRdhTL4KG0d0PWFc8H+zamX
ckFily9MAMmSN2R1wUadgvkG+x//L/Gqf0PWPAbyQ0G6TMh/wWobVSgT+nuFfSLj
2paOjaB4z4/jX/L4XbLsCd6wDS6zU1P6a+xE5Hbfo034ltqcNwYUXYvOtKfaM668
/gKor7LIHEdyeHhq4k9lTZ6PGClE3/OhPqRRPxxdzQK22CwTmA1+uWLpt5llvEuz
gTSAO0VlfuxpmtQkaYuMiRei97BhirPw2xpfaRwdZp6kNNTvezQjRFnBZZoW13OL
3ihD6MaocHtqfZCpQdg/IcuI/ssHw8LfoYwarvnI4XXYVUed6KpmEawe2vCIGVpW
YgCNpdD/bX6P6ZBNQv8rKrrFT+GrPbSMI8B3I7kRu0ptEkdrnwLEftp1Gf5VDaoZ
l1C1mf5K0KiqI8Yuqduthxy9ZweKMA0F56s5OBps6Pql2pU/ch1ymAEATXJG6ao5
CQbCQaJ5dqKTFYCw6Xs+lrVpNWwmveIiQcafQKfIziqH1h0pFerETdn0uvQ8Nfum
NYck0Qol0qVUdhm0+uc+VpxXe/0z+auYTkYpivyVAWYr7ZZOY2LAmUQfdKvEvXkW
ATDFTNopbpTxn7OuIqdfqaY7stjDlX7AI4VMcJBUdlW12WzWGXRZtGEMIJHSI0Q5
/9dVH7qskCtgS+vUMoeCuswlW5YzXY64WEoh8MDE1QZ9zRog4vHQ7rYcDFT33l5S
5/UgTLBjyRSNZc277q5xiITuYRbtlc8yUs/L5yMHGEI+eQDIhup0UVEDlYWFmPas
TlLDELds5qXMwTUYrnzFq7Fw1Zq/rnSzu87jqu0PV14hHxc2BSVFWj7/TUoRFVKq
ZFXck3CtyOcD3cggIeob+gbVuSYtDKW6u1/qshaN1PqTOyVSngVvETDuPeBvlRmQ
bCKb6WCO1dgazNrI52E0rw5JVGSdk0jkk1ED9FNQqYX2wAETOx53ocq92DdwJ+ko
a3oJiyV4yY+u2mbllEmGYr3apsr3FOqvVAh2FAiVKdcYSo2Z9AnifKJgxpZ9Mlll
pjcMEJjL/PBvMkbUOS7mx8b2qZ/o478F0Hvv32kfiGe40hlIJOyZspitVUKbOK3D
9ZAEnfh4rhWxjXIBgDi7iBRwJW7P9B8jilO52XXRF1gIoXtORESfkNK1eK3sm3o3
9WUhMpm14HSRkaI3Rli23Y3kD7xH5MCjNGmsDDna+JE+ZAdwjXxoMB0EOb+Yq136
1ibp78qLgprj67wWGtwgJ2H+vqlTMAJ3KZwY3g9iJztwnXk/CB/Z/+L+WseiXPMJ
v0FBxGmtXs/Wd4f5lzBBfLdTLu2y4IBoQHwJfCjCqCiRyVrxeozviJeT/4T6kMXy
BliAlO9gUcsanaT0ZiIFpa/FZ/w9datza7qLXbOzgerW3zeaDAoDtUyUVzwVm5kA
hEhfFJiYE7AuJgLQ1af3n5sz0K65ICWu/XC5jxaemgexlrAVegsTBPZ5LUQq7CMp
jj9Hoy7MH77Vdippg6Fm/Tt4DSJ9punol180txawVsrAn79+ugDI6crsgsxlM6xM
ziT3rwQsaud5y8E4TmWEgGfUrX9RMFq4Ck4CHsV+Bnc9unyClKGUzB2DIp+D78cE
zoxMwO1iNQbbjO47Wg8jyV/qGeBeH2Ct+I60DhSyDV5a8IVZyYanaxcJMXrxFtVc
RhgBdvgsufqpuS6kpAhQxNo+4wx7QJj/DD4eyaceDIPK0RK/jk383Ibr+CkLE/ux
pWbNJO2MiPvkx9r2J5vvZgThCv0gc3dEeArYBGkqhcYaLyKszFPHFCmWtvMMQxzY
RSFXXz1ujM/gcsFmzyoAOkK+E7cpPQXsNVHOTwcjOsRbczQg0A0xNQAt+iLlasYl
/lRc3ihLNci6F/dA6FmHfdca9o0v7q1a2XdZbtScac02QsUjoMXnNUojWdUuZ+cN
OZA0H0dMc5nZxgiKkgMzg0cxFDOjJ+9Jyc2Jh/54JR4bemui1ywr/iMFb7XYUewD
mCyvAXTOVxrcvVsL2wiUB1Elhxte4d130GWpx8b84U9FfzC/kf1Z3e43HAk7h0Be
6fGlHTkEQCncZ4yEuLfkov3mZYj5CSsWQCjpXUhRRRxbkWXzbvOEWK3226CpO2Wk
YOxwEHEAALTOiVlgys6K4k90oGH5XlzKTK0zsYg98Qbr0z4eDQ7ZcDdHXSMB/5xS
d2VoE6JyJn2iIENoCplEyf8NLQtw+pTGzq4zPVT4/7YCUK5NNyNvx4buoeJa+f3F
He22Zdru09PLLhDLaN/wjJMbQiiopfl2P6T7MP1lP2G5/szY34b0c38YFCAz2LVM
yREU0vaBcFKqhSu3tTBEoUtVcDvT2GZItNONTbpxHR+KnkErVgihA7E3c+f3muv4
vBk+QFHA2ub171YMtAoRCm1YMtOnoSKno90EKjBsnBQvQ1zvX4WG5Savvtqp+FMo
JS9JJfRJ+Pfux3mPdMk39lew1UPccrU7FcFeO1/XmyVlZPBflBTkeJ/lctMY7aNz
7OaQ5WLXtlf8UdKywDDpj8xZ8iDKTfIZN4PLv8GcIITNEsdvCl+mriulX2W5Wl/r
vm+MPORgEhp6XgoLXynz8bGogrYiOqnMWdzlU6SRGGG/yyb8kUY87OAReDvE+kMe
BTqwF7+Wupcgkqfvn05GduKq1kPmQAbRGCvZKr3WKpcqPQmttWuv/dM7Kc8/bKwX
3LnmBQ87Fx4QvANyZY7+/xC2DZb+XagbOMBmLRlkqUs2FTh0IuQNFyZ9GasD9jBv
t7+L5k101U9NjvGCPQ9Hs+XgYhbd8v7eRbnRSH4d42fP1aFqmDq5bmzlL4sdVhUd
t8Qci6UMrnr7VfIPpr+VTMmpDToOamn6waud3D4wNuW5Bra2F1uonsXidQk4PsnV
Ip6XxOM9BYEGmQ0qqWrxeeIs52BdxHidAbnXL94FUjJAVbBW51U5L/c53hXUs8DC
JkNeF0kgpbPA+38N1SRJw/p4U3ARb2prWYu7AWpwcFBir2sQDhkCPmk6yS+LK6MP
shkcMMqwUur+6cmszX5W4oKN3ih2FLDuKlIkxzRN0Isj+b8mhak88CgVBLcNEI1v
8Z3V9FkhhI2/8zBy0rzh82k7U9DvFc6JynOyttr05PElZMo3Gc0vv8IEmEH5idpe
1jF1DDHSdEA40mTanyVGiNJ7nuBRHlccY1fgnEfjbWcBFWUCc2854v//R8VT/CVv
FMgm05a4iK8tW0YYgIcQUuQMmV90ZtTkQ7Ugd1q/CXv6FHL3x0H/GdvTpw7nUYe1
W5HU3/NzUVgqIVzP0OpUGlV4nqlmYcCHnvbD71NZVZhgDWAsFg73omxTttvsoTbB
/+6CoAx0qJE9atD7xdcyJb4XsYjF5GjMCa2fy2MSi8bMaxIDH0TEG3K81nKMSVga
vMYRj52H6Z75g/qGZP7gOAnvbNIhPzrkPvflZfk6BkMKSCR+Uh5ox2zNpgLD3c7g
PxRJ/5dzSFhaBLOlt8obK2MPzj6pkMN0L6KI9LitwO/oPR/YT4732qsRSubzjITm
OEPOmfPw3W4zIe4a3ZUA79xnDnm/BWUjC9k2/im7JqtYEGX+3zy3SO6CpfoCDVEH
ibw6qzNtCk/2bHfALfBCdcik5Ele3MrKLyVlZ86Wonl3MCGveM0dtePk4UFPwJCA
cYHxJKOeFAoTVrjoHAEsFUxcxXhFi22j2iarGv/uW2La0PlTPQbSZz/MR3CWKUWV
rEediwFZzF9tVwH4TKs5e1u3kCJ2II/ja7CjmXIZU9Cw8UrAxlwOjFg9AWVG8mMq
BRPairIFWzJh5jkgb+fEIDZKitcYnvxiMc8+/Uy4xcPJ3noNAAPRd+AgLA683Ev/
qNGja2TVI+STej5TufEcArQBJR42li/ypcuYVGzVSjmImam3S7tT56Sg2aTabH0Z
WAuE7D/waMX+J8/cSohH5QZrQ6QZmAlCfSau1hoT0r3gu6lkpkfHPlM0uLkmd6GU
RCcRUyCyv8fsbunkwiV1S8EXsWEqEwRrcHz2s4HRWv5/VN5g9VvlR6lHxeHWkH+E
tjxx1rUttNn4WGTaWBFymsMIa9Y3kD3a+DnASxJW3hxZ5QNfO2vsNY9oWzu8r7Ne
feuSo/xeDSm5AgweWXcFYlyaYs2UEjQySHnlAH4Qb0rzYEKLUBQd0e0iLtFd50hI
hKiPBcQsTSOBkBVMXzBZtgLBLoXJF5s3/ir1B3h2OasGA9JRxZQ+pG+rML7n70xe
SgQWHSMygUq/iHv1PsCgmIR3RuyBTyyyy04mg+7GF95jMo2KcVWOlbH4PAaKurKa
b1Hq776TzUPFXCYa7EgFMwDUrl0JZeGoAUfQhW74ATJIFRchkzAMZNvWOISznKg4
CYnMXb8yN3w/4GKmxe6kq8b0tesD8NeLiKquWqH34ESGdFiQtnEMYoxvVHtSMO6g
w5YcBGHCGXwbkMRF+TYNMglIfmUnWjOsIm9kvPt7gHml/8AeKGvRKPtRD+C4BDwN
gtgdNYjJEQyIYBdSrKwkvKWMUflMoyflsBfu0y8g9DxzedGs649BSvkGiroNwmFj
jBC0CdcjlAYgbFdeMinp24Ab0HGwIDaVyU9IG0/iDWquv96lH90JoKbOcpO1ESKo
KCKTQxKisnUaUDuDD6XDF6S82cImYxdTxKmboECHnEnBEhwA+qqXQmIkCTbGuNNP
KbIRI81sdAvvLZN9Pzc3dP776qDI6pROyX5uwaMkyG9hC5sOFKuqGbh+Ily+ymSK
j1dkWCG+qqmJY0Q8mhRp7MaS67EnGW3azsR3tSljm2tZkmYO4Zbg7OvVJREFaXu/
SvpmaQ4GXG1UAfwBcMTUBphE1RUX0kxgB3xSMCClTVJqX6X0f5EKb1vkywpJBvBU
7EPd0Q7UAPeXmTes5pHwFDMw6ac6NzWCV6QrC8ob1L7VP5Isb9zrNRVC8mPjfZUT
5CBemu8yVy4wfC12aHNMOvpQZLsusvizSHsoyoTbuWhzOQzWUjyIHLZ6viwxWU/M
JyH1g6+5KmraLVpCNSbyDgMKNUOFsE0EauyWXTMqHQhr3POwfqxhoCRgMK83trt5
efF59fF+FNmMMZh2YmQCpcSgN5zxSBDGlJFfEejWVjIZFLL9BL30YbyC4f+5Gdz1
0byyIzDIiYUSKu4wRXe+Cg/Ey0UlyAWXMSyNmsAUoC18mc4RQLv0iYtixKNXI8Ld
n3+TKeklLb9D72kKIY9M3l4H7RptE4EUhizogkN0ZzGPh281jj3avPvblzL4/P1U
3QbOUGscSIiH2j8imCGxZJ6Ky4pN8w0hroma7oOYhnVScYGQtaAfW5DP1hQVCdy8
a8UjFpg2d4BIO0hejfc4CX0c5jMFMpOKv+LetF/XcIKqzobk0AKwXur2LPYwgCGC
5oQexVJEQlvr3CHg5l0f02eo+yxt4iQDs7cME4vUadsjfsYvAY0XXtYPZinxzntg
hRKt1XBxp+O2+665166zy781etG3pte5J/c9mNYR3x6NZaGVHrEm7e7o9M+CO91X
IXVfihTSViEmKEsnb2Fc7cJQ2pEL4cZ7TZWUQ9QgFve7DTsyut5clFr7KlXKapGd
QFzSMU3/P8O1RoUIUwRoX3e61j9Q9cdZDZwqxaNTzWAwdOOVB0O2VyRhp7ekpxK+
QXcPx/wSbFjEdQo61im3HHfYqwGIzJ2AbkiuflmdxC7iCPbZd9V36ENVpUIn/tfn
PRKc01Dyt0hAmNJgsqhNNuXvcE7HRjs16IZCN8GrqCCdRYadGIYnsyCWDl/2OO8S
HzxxlaMl5MXnCOiG45nbCOR48DW1oMAhEsCtbfX2v1DQ18xt1jHTN9WYB9m6wsNE
/bNJLE0JdoQk0uRHx8x6eNNhie/ukx2VH5ZJkXEcScVh/GInC+ziF4aDEpRT4OJX
fK9Wszj5hXNa05xEXqmNiZovqIsil6GiHYCf1T9RyYbYmpo2hnAkkjyo6inHv7F5
KTi/pJjZ98vGHDhP1OrnERDVQiCa+DX9Zml5krR+0Rv4XnJog6aIMhhIwGF/EpkN
ApvZC6OTp9o4ORcc8xCWWrNDDsOTWXfN3u5pTKTwxlkKMFMgEp/zjvf7qfzic42V
Gx1cOevnWd7IMbu4aSZ73jp7SSre6wvyBfHX2X6AIBTMD/2lcBGezJ1+RCsmV7tA
+bfrN7JppdY+6sII7GeWRZ0Q5HBQuZzl/IaTfVGud7y9xBoHsd0JdK9Pac+xVJWl
gioGDpiz/YuyUwDAPgcyoVgDnQD7CkDAJ/uAiS457cZ2WJTdmUac9s8uPVkOvKK7
fg4w90AfkXWW4VbXEkeeUWENjDkibYvGHSH8GEA4T6SGPOh3l/Is/mrrhW3qw4FO
O/+Dfbx4gUXkxfVI+UzqK/VNdywSq1WFGL5cHbtIXez4AhsmJJyRBI1rwOd2E13f
AHt87lLime8pNvdTlfUatsrHLxXt6yRjmfDDQiLSC8cSsB6E3BWM9nfNTA5+KT8b
yMw28mXMcA310WehLsGH9r6E2px7mNFWMLRIL5+Ceczrdcg0A5oW8Z4mK+EgoaKf
fD8JcCA9dK6C5ypBSJ8O9BKXCQNsMfEZY2yHKcLpk+HkLI0fT2pz1pYOmdZS5lQf
upkxJwj04YatGylGF+adj9dVT5WxkGw8YFKH0/sLZeIdCGyZ83lDv3O6+slaOuxY
ErvK83jhAY9uQkxaURdYnFGUuIKWueb5BY3LmeuwvrRDL6Y/3/i8+ZODnqvYmeuJ
oKHjhV50TGs0zoY/HTJ/wpxmHzjAw/083fq5yKTvMYeWQ2MDQqMtACvFum6G38Am
Edsz7uKTx2eBpYid1sBt2rj29zokDRNvh7B1OQwSVv8VNlhwWntgYzk9N7Otkg6d
OQpc/SMKhRSp7uaZP7eSObLXp04sM0WzhrpYh2ASN5eThYoCKCBZzGHykF50szeZ
/mTNL17rDoO2PoNa8GJ7LJgmxEa6+jrz8P+6VwZTjo4fg1IAXvqSSBEzvjOxAOFD
vs5X94g2NJGahlZhrpN3lAusZIy0eDsTkSKoC7pok9ipP6HVL4h/UIi5lElzm6ws
0hS5/V2dwfrcmMozTSmg+PtzYYACze5xIDz10POmCblnOeta1SKzpqcc99nxlgzZ
lp+/zAcQOA9nOG5SZl9sMhMwyN8txqEDHRfSVffP3RsKms+fNFlvXU4P5SRN2Hyf
yAI+7+WCGQyNPD3PFB3AfPKNyQIirdmjBavxmJxHzfCXpil9EMjO/SjeEB16A7s+
akQ7M/4RzgReS4nnVx9Qy70R2moRkY0nn5h2xwbcgfx54MTRLYhzGxe4ZEL8KNCn
aBUim7npXdFD7T6Xa1JcYU2Lvjt35jmF6ejP9r5wTZQq1v+WXHQWaUTeuG+/bFad
VOhkVJwb33MTm9kXOuUZ+tuRDwWw5Ajn0mb6lsa4JnRVcuqKRcIn30JHDa/4hsbW
spaS//W/wEDGm2ZQ8DJk2ouoghT3bvEvzaAoFJnKxOiki8eyO/BPTp80rKsS6jvm
XBvCYUY6SkBY3qPmMzeSehI1r7iuPqFFeXqNVq31yk+j9wFTWcIKrVm35qFwnFhB
xsnX9wRXvTD+oyyr7cCT82mrFKm6chrGs/c+8EhXKCkKw8N60jbnHunCGneLDQ6l
O6i+HImxeB80p+x/Q8c3S0eScWjbqvvXTRCZ5N81HLULFcf55TxGQBnMMlQS72+E
CQfi0B4aU19+0stwG5YKICRxjSyCrzB77TaG5+pjS0w/AYmGHOsCcvAsWmPwnq1t
wgL9qywTkgVhfh+UaCJv7afR3q7slCogHDSwME39mBbu+FkjNv6og232qSXKnvDp
4z8Ga56MMuS9kljO4c0ywG4SUY74Utnr7xxtlk+IkMqBGt4diCFoGQ8irRoHQXtA
Ge18XQIry8UKe0s6ebkC/YZxCMf/chcRCRyMUUQCfNMrozBPwLTXsJ7VRvpsABfF
/8T1FD6k3riy7SQykBAflRWf0jwh27Rufgwx7IKopS+KdJTxogJVXzF3xkydOdMt
YUuSgOQCQcMPoWLDbA66MYjx+gG4p8E7nzMrhcUvYAeM0OH0hSS7VMJlsoYRwh5r
lcDDsFhOzav6nbhh/8/pFzIkWYf0Gox+Ewsd4kuLO7XVgRuZaxu7WaLhWfJr9Kxj
nsH7P8DOR1ZcuIm34G13uP5a2O4GdKvg8zOL8JyhZLXK0fIRXEV7n7rhrgJ6KaYU
ir/do9AGiLY4uugbk+eKLLnugZlAhtPUzUopl0j1InJacD+XSCoxOzyFZUzbodkN
755br06P8iF5iYN3IAF31LAT/N1gkoAsTZou+gs9qAka7/TiPtugaE/yY2uaEAlJ
hpDI3vgRMepsuAcyoreYokgqdWNUe7nSCkY27YZyChuUFanrkWY9Sc9kMwq+6x64
WVz7mcq35tWvKS5wQ5SqMm/DJ6wEov8ZrTVfsjzRykXHK0okM5m0J5jtD/yt4ko9
UWHUg51kdZDxXyK/qkcXOXelE20Ni9zRbbgOecyxmGE183KNZlPVBpRJ2fi0r8xg
AHwwMLTi/OkqvRaiY5c/6Wre3A58PPJAFkn6Mw0pOgrqfdxRevR1R8D9kpRYomSx
dgSPoN6BmxXHhxhGe3hLuQ13c9RWm94chGxWHxUolGm4u8OhXXaT+K4I8JqR3O2J
yYBjDPTNsdx2ExC/vQmeJr7I83QTHrPPmIN9N/zYv43e6H9UN2b2ph0OMXQVPYvD
SGmCMwb96t82oL51MAPajJeCSXYSBKImxkBZwVMXIEXyHtqMGZ816/xuy/nOZyKO
aEwblqdCKnbOIGupFYLUukYfUW1/9jEJEuIPzEQE6TjeHW605c2UHWD4SV5MYVFA
HCATzHCKxJwz23FcDjb/z1Q5J827KdlgRISXc9Wwt+94I9EXGzLEOJSUepLAf2lr
fhkakAe2sV8qVTrJDJNdx7GtCuYIVZoI4sc9T1htAGk8fctkr/hkbfxe3Gq3xa5R
EOyJohNhNm9oSKoGxGg+SuyjuWEST1zXm/hAJPgCgITdAl7vvJnkOLyim53AKAA7
7cOnkBkjSelGcZdhRQzO+/G+DvV9NhoroAkGZFC2V9EPu/o1Y/u4hPVH2KLIYyvM
paO/HtNma0Xe8u4JE8XUWqnXKgOTBKfnw5Oztqve2Ac8wvzqh+CTtsbXCUHCQByF
btWQbUawwJfWTSUHlC4OXDBSHVKTFF1mKKLPIUgOWsrQzFQznpfLtQxbFX5ReIER
b4D48y/8A+J0pU7tM3XF9elzERtiSHBVhhgndItiGpYnHWOSmr+5H1a+fhqUCVf5
XvXBL1zMnBngt1ul1lGJKrj8tNZRu+IWWcsZrjpXqPpfg91R7I4PNg8DA0F3VOce
Vgy+TadTr52qW6CQhMU3FKY0Hx4z58cGgM2C46upoMFp2vWT0Xf+Oj6yNoJUBQmC
MLMplDzfmYiwpMhMO8cyudR+r+pwruc1CbM8BHY8T82NP81fqZCoeleQNMemWnzS
5uWl7bhDg4w2q50alBIUjVPs4gt+5M8b12VU2joA46tCeUpbi3fzUglIL9y98veC
CyYhmyTgzjnNYpHT865+1u3WZbnJ/2ZlVQJ+/SKG4E4wjEI3r2y51/wT9da8jtpp
GhPTJhsPIuL5uVKIdFP4WNwFx6owrjsHKce//dNx9YSg2M4gc5vK9162EGBh0Ffg
RaCZb43d79PqQsdZEAsRW00jY7/waycFf0nefmL2Dcl+6FpCwj6zY93MmXeOqIJy
V/R0pWvAnSjmPADM6c4pJ9IPQuE/fvV5kitdkr+wFF5C1Ay0RAyTpuikCMFEJiuo
N/FOQmwDLSnmHA3+ULISkaY8iMvGg4c/zwmBRVPf7630O5gLSNunlAdvDFPGxJpk
OIo1Lq9i5rldQi1vGaN6gbX8f8YxhGNwPHQujehFz05cZdPdlpZJzy2lBBZwX2bd
rdlJabJcAc42DqEjPDkTbKFX+eA3N71Ri7olo4CEb8ldI7Ulgh4jR3rz/DP712jN
2a3TXLGWyaHbQKVQMI88F5GbDWdGgMGH9++MKFwOUr+BREhYlboFltJbhE0vhSwx
XSz/cilU801QOOXPQXN2K8wndas2OANA8hqqd5/Gd7V0Hd/wQb+5RVLq22YMrq1m
8ova+F+MxAKej9wQ3Y3uzEypHha/uc7tAXbBg6DxpknEun5DvxyeU4BeDoUl88S5
h7tX83pNqW+PjEvuUttzTcxlfkZEhNGOD/tAhZE2i5h8FGmeeAVg88JXM5lJzd6M
Fm5BrPlvVo8VfcWyTGqL2Hv8aN/k9XjD4lxLXxxD8YhbdgaMkEP5RLJef9imyybw
upY0+CQLPIvcVrO8/71w4xKlKQkvL2rYQaa0DXVBDqqtzuVoBDJOF+GuxcPNnJNT
Qfig/NOCR5YoQ++okTKfyDDD6YgEvmesgAQ8lfLj9Re8XnxVorygmEvDelQhxbCt
OoR9qrNcW+d48KTLWXLL8gLDPn0t25dhr1xMtd8uGWWxZcvNzlaTIILD8xwrtUJO
cwb7k+SP/PwiNctDjEbbBofqtYWHXnwgrcDn6s9uf/HDnap9N89WbP0nBlSuN4XT
/fXPsK4fL77mxvholD9aU/rH1wkameJ89cd79NQcbHDmmavmEbMXPIwkhi/g+lfv
X+rAgpyusudYI+qzrGsidWCelJdgp0xDuztfawA7d/P2TYbuqK0gdB5Bw1h280ja
hSymycpVgeUHbXYzUIhrm+1xGlNex8YUv9QgNzXFrfQv6gx4bomA7ibbxt0WOEb9
Dt6Ci3vXiuj9Khb6QUFaqEbLpw0BglMP7+qvfVjmv4eqqlqQ28SFPB9ZFVqkKOIR
AhdGO/y5h7I07PEsY6cldBqfPeGwblrQaxVttPWXm4k=
`pragma protect end_protected
