// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:33:35 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
QP0hJ7vTU7Slv8cW2Cd6/a7hNqdsJsoZnnYqRGXwtt1nv/mUXO20N1ESPlv7Fh0Z
cG5li7JDi4CrcCXNKcDnuQcnhHxhISlK7R5vGi7y02BwoRXi+JvACWLmsplGidMT
Z1B0dZhCbyexI1F1k77aU3pAgq3Lvka6w9WAt8kqI7U=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 6464)
ZP7eKnITdggw0rEDUeF8HByKxT39fBo30JcVBSRXflI2BitvDrkRVzI/RLQyFecy
hrAr3SRYhz1KWaYfEgYfhsLsnfDGniGpZewY7j+YAjOVOhqq154WLkJx+j8A2Yr4
zLJFBU+ejgAhVOu2sfOWnCZzpuAmHkjtIcvoAf2Pn0KtvrEUmemtUiyWS0KAIm2P
Oi0Xw1/MAiYGXf4P9J9PS3uvGP/xUuPYZoZSMJdE77G0JlqsIBW+o04ZaG3VUg+S
JAtBPUKqZIv5BZv3iVnOss8X4Sz4U/U4K1G60r2kxF4XIia3Cb/5UQhnWz8wa4cE
TVNMj6PRlkhdpqEassyQOEnqCSxt4c5EHK4M+J5S27yjfbFtgGuolAQF4vz5L6rt
s/LoVxdsq0sDAGd4quV/ZMnrZlVPB9SgcrfYsN5QAbb3qgjDh8JMI7XzpHdwS0d3
3ssd00WWoCZ7ZDHfwibCtR2SA+m0j/eA844pmUWV4mJJW6jLcY+mA9nurzA1spBu
PmnYPwWia5oSN23bgkByqPRG6M/qkjrggXYDXMbjx7BD/vF8YYxQ8aiNJ7KU74zH
BMSL/9Y13MoYu93iF+FqorchN/4Xo8bZdeqm7UoeOCyJf7dmhLIjuUkNFi1CYVzp
5BojtsEaRimJeLSkuNlp5fOFFnYbOwbM5rdLUPaScrXMNk84YMXS1PMbkPKZ9sG1
sFKczw2Fu4JxBGGJ6zw2Uh8tMWDAaDFNEFYb7dIQeqsbf98APHPVpzAy2JcsYAFL
4+C1cNpVkumb8DBzyH7ZwWjyBBWfFhOYULfMzM7uOjz5q4gihWqzSkLoWqwWhykX
e/hxK7Ak9SHKsa9lPdiAierJv4cjj5rpG8WTQABWog0KdoY57OJF8JdViHFKDdAG
qoF9cUVX/AgA6zF3aJRyHe2AextRocVJkUP8iLSnCAXFRsUFNYL1h6NPDn1xRXFc
0+e18wlu0RVerIpirHYBAySKXsWNPhnQrsG+KvZRCVpIECB9HSfGmbtT371HJfFB
7cE8oJEFfZptjBZYFRc3wOQM+OZ8ib2jmli3pO8DCUvpHEUQ0q85es6O3ZkDT8M6
E8SSdTM+4b9tSiSQxnQcDoFtRcut4nm5DAAKOCcdizP4sEblEeLrjDdKJq302mWr
i3XgLGasjvx+0qxMsS7ybPnzJMAnDNcT55EaFPRnDwEbgABS3Bcbdj/Sw/yETOsC
PbbGoyXMc4C7XpSna5FSFydH9mn//RUvGN1oIZ3OgycP+28sFOtsxSN4u9+fmuNp
9u3UxIpRb88mkeUQ/QweGgFoekDgjwMuo68ZdvZQ7zInTG+khz/WgcagLPb1UoJ3
XDcTTCH6F8+XUlm4TYG2k9Ww1KbOwbcB1rvIZESIkmsUB9D2aEuCQ5cZsAjeyQ6x
sa2ijzq4EIBtrDO1jeTKiCWB6DFOF+MZ53KQfyuij/3HfSyoxQ+MvKxsjNPi5xIH
BBCHeOPiw5liRjgHLPavTLiQ3hgfMgaAeB/zpmwvpvkijU8vzkAaLy9yJ1tZ8RCz
pJkK1Bi0vNyJFosgxD0cct01WfQGtbWob1jDIM4waXMlG0cIbEAHdYGdBJi9y1Wy
uCrRuHTkrESEchUQ3UUhN8JA153Qa/nPpjgSIwjtcLXkZ2oHxaopJBh8ySMkoOAX
YClhb9TGQIgxQhT4SrPZvdv/AR5lr2wfC5xpIrxlbj0yp9edOQlnB03ZimGx7VEc
JGSbziJcCWDB++XP4e0KSVOHMCQfJZuN1sfEQEhbV6wKAsaFE6hqFTjsSI2axOT+
y7LzN0mvvgh3JkVueTMhsCS24aJZ31BTmfD7CqIYnqv5c4He60R96ATqkRykmaVn
O/bUca6VyrfQE7yN5xvJrXGeoayjh/vINHBEaVYM8hHuwdZCThMb4LAhXqC9vJBW
qEnqPt88wmUj5v70KeByr5Zi9ltbp/KYX5B0s/R77fekx3IJUxhhiQdHSo0H5sVU
m9HH79enn4iuhYhBlP8QQ+oY3jwEcW5B+WwaFS9mmbLzfJ7UoHKIot85zzoI3RAb
9XF6jMVWfBAfhNpps/aJ9XAhIdUZhn6KtvvRtqrPRqWpR+MNDHzxU7IsKH3nSgvX
Cq1WPJZaX1IzxkkV/DIUirb3z+retgNR+pQUu6+TOB8c9Rb9+kHAkwf9Ak/qLYfh
6BF8bU7yRuOyA1cBxHcyEO0DMn6HiwKuM8dT79/Aqg736kDOvuZBxS0Fl66T5lyR
DZaxnTNT4Zg3b3oSMooNsQzt6h4d9DcXcgGP1UWlffVywl/tX1HI292qqBVT99wc
XollOyodxar+X2uvAAq0uzrm8fMu3CMjjp9dpZiXGJCHh0bWz9jjZX+EPrvXheKd
fSpE+0TnzSqBrdDQl0UV0g8u3AMuogclHg2nHdjsFN0AbQd7TlAy2eoSDIk+yGCA
Lx06eVc+B93nLQ7N9J4ObyUTcdDrW9Gm00oRZUUNaxJrTyzUbNWBOftp0ERInE/x
RKuATtngzyrep8aF8lWXAJcjN4KvtHTnnobTAyCg1zhK7qYlQPssz3v+QopVAKUg
ZKOxv3Ygu2Wl9i+TUKrmRhtAqYEXgMmA5KGvRH74rD+gLhR7ubnqvyG+t2Lex3wB
ByQ7EuZ6p0SgHnGpC66uBlkxzMwEZzMfFg7N7a8KvKg5tBjKnBeuWCTjPtP1dOBs
EqG/u3nlPViLRn/xVW3pMB4ojOJoOpyFgrwTfIUejy+wktGQLC3HQ8ZacIStZ498
2QdDGXo7WPE+AXeRObOPH3zr3GoINKsYsGeNc5AoA49RF8/RTZwwJc6h+HGHZ6aB
4SLKQLYtI6nKvZf4FBQrS8J04YBxO7daaTuilnL4jV6zqI3AU2DYJ/2/TSTEm0SC
VWAbgLSXMFg7yuUqmfgJNqyktmxpmCd/47aMVc5bYEWFGWGMwfpxkKJqJXGo31RN
8GuLwn4oNfSK/XYnF+KryRKujPjYL9f26MbCjJ6yau9vYktADhfZYFWNhbOqcjy0
0LHbIzE3+U97AUxtnow6kGHm6DKWjT2TVjRRCWu+SmyO9EtrIMXfwAYO5W0JjigG
o0iOoPVAuFmZX46XDXYVh2N3sWeeU5KIHG3vLsQ7+aw3y0uiRQDoXQEwYPcur51/
EYnGOkgOPf9aZHOaej+kZwN2IQTh7hgMsz+Y0BRjtjBADoUirK1RzJpMOkJKfesR
L/QuZjb5wJ5Us5YS8XnsLrqL+zObPfFdmAKzP6Iz6tGestRA8Ww+WQAZyfxgzGdj
XAG7nSGLpCxtIkhkQsL6npevyIA3tXxvlYL1vOjr56rJBy5nB16a7iWwSoXTvofP
uQEcTBip1PMpCp9djz/HmC0PNiWEywwBrrnO64IJKe6Cxt9LY/O9p0LuSuMUjmRa
rgvPM2WikLdtHf1M4nXmqApqUazTFIKGOS+ZsF+t1x1WzvL4YPMCQT2pyGfMnfE8
XiSPOXVfCzrpzq6VyLUk/GX9AjTitoJhSerZyQFdgs18iJ1LavRjUTcl2XM666sS
yqelaPY2n34110BsHKu/onOXxbuEQISWGkYyXF1cyUqgyrTGSHxdZXxYFEVFnBow
op3zdj3H6R59a/kL2iOCXnkbVYqP5vuig1qJ3+S3qusPjB46+WNS5u8HTErzOyQ0
v1jAVRBTFBX9gpZ8/y3dPTR7igqhjTCQb6kn22NJ0ZQ/v7dULP0AY7GfNV79AVKg
WxMmhx+tsD8yoG18wBeqMZbDcgR2/jt2Z2aeixKjc7lkkSmAv6iT1lFGkfmCohll
q4xstXMfqmfxz66SX79BEmJcb3Pi7moIAibJEKVl1RQS/3MP7inYkXD2YA3/1ZGf
YT4EMTniiT1lSu5W5/OXPj1hm6c9PkEdBktuGEoArGQUbrSr9BHymYjz/i6ed+FH
DZDqj+b2wq9sCMQ45ybGkfMNB2XowczQjAO7WH5omJlNlbLonUCrl+ssMBJwMo/v
q0qsWWcZIdLZ1olt/tnSzAgTMQ+8RzqWoYMLxhut+2AHwWWDejgRsPFo7f/Lvn/C
9S4T/smjyG4h2jThNncABwnaQk4dFnIf7gYtgrkO9pnvytgwUGRtvjyuziXOpTzo
FIVcoWb7JC/V0z9BzWx9w3241AWFonBKFPdBkBcnQ/DX0fw3W/MvygKONIPXTGqg
6OfFPWyBKs8tlSxqF6YPr+Eu6GUdaamaxIx+BYK3sn8AogNz6bQxvSl98k45WMDs
Fm8AhMReWoFAuqCuL9uqmowaSurM2pZjyl6Y7vcp8OrsSZwQ/PGAwCiLXdJo/hAP
CAwpmk+CXlPFfVH/Dc3tJ9aavMkNuWpDXhnWv2WY5V0RVWlDnsZ+8lVo5f/hb5AU
MhxBrQwVQgHZOQyOD5n1C9rDiHPfz0usFjv5Qdd+ZPcP5MOsVQDg84dgRVr4A1fJ
hDG49TOCjv+shzwM3g528YTmYrBMU2dKrtUrBDCLySdkGNk1DiRg4AQrQgmIZugU
U2zxRQjXVrKkFTCPMTyl2rUAyKp8Qh+Kh8OzCeBhDc49wSY6NCk7DqQek4l3a6q3
sUsOqPoiRS4SvEnfijgrXRoJ5QzTGBX/4WynfUoztFTL6sezwTe39PAzpgj6UEU1
xvLs/H7ydXN/vbaVp4cILNcletMsurwhLQ8Gk1RWwbB3zneyK2sLQ9uLWKMRrVhg
eXhFTxLt4ittEpBuqnUgu3I6j+V6fPk3XTze+ivGvjdjRWnCEZmoGloFQsYhEriH
vBncHJikgk4DqTP/UZZC4SqRkL4ZjiHLSgo/C+KraJKkjtxMoN2Hhj1oO//A22wo
l/IN5qJLoktdow/li32gKw3HbDn2d0MDfSeTrZ7uktgaSqBH9vdr1KUwfednxBnv
i+vybBSCubuka+rJY2Q5Plq4FoCW6so6WGv0/zlq3IHdZewyMA3GL7x7XQ4lPn+I
F/EUfaKlB26unooeDrKiVquj3bQYuMnZ5FZ8nwWeAtM3NCh+wCfv/QvmW98MYarf
pE9Tb8r+mzwRAZFKQwdnexPrKtneUT/nokRMxrV+zbqQxSQ8wXobVltCLx4wq965
qlyOzWs/6iaSv6E5Pj6MRNHhLxfDRQjZA4LOM6zWxmjq05IOiX+K8XsGUTSi+xuq
lqhnBc5fIXLUYBFiWt9PX2RGLjT9SjlCq2hjP0dmfSuWdHtR6izrgAyz9ErNPsg/
CikprvRlmNGSytqO8tatfzhpD0Ilixhe/uDYZRJPCIDdyQ4k59zleMAc1a91dQD9
iuXKxqtNX3NNtsX1ps5CnxKAtdkV1pB+56LA27GY4R+BlltVaCv0R/LooGZfxwba
Zp/H9DSsGEOayYe/Lan2Luu0rjIrKDfFWirJWh70Bm/65oYxCL+Nxz9RkKxjMS4G
DbAA2qzLQCMP9mKqhfffXl2pHBPXf2dgOdVH+gUFpq2LNnZ7/0BgiVIucPh4LPgo
LVktRjnMv+Egifc8gwpm3UEXHFTiX1UZr4nnDWCGvPnW/z8nM2fvHFpxKNOH6XsG
+VwdMoQ5BSp5PPyJW0fQz38a7+BMGWz1BazFpYNp7UIFzB6fzgoxMVlRChpu0Ejj
UG9J98gloiXpS0WVpvCpstAM4xf2BRkRiEKatReqP1jIoPvDaSZ4VEjI4GJl0kcy
j+oYagfz6SR/EVSDn3TXXAQaaceUiN9lYethDuwbtbWVfUkXuEgtlOi6So3xejvy
PkkrVpMX3rKbnx1JuIHeq9+dnCtA+hOz8FCyZ8DgzP2znFRZPchGszHXYmXiWghl
ps74oMn04kUgk8cEC2X70vdVsejSBjH7ucC2lyvLq2Kx9kQn1dfdlhfiTR0L/gzO
qw+oQ5E/LCz1GICszjpWMCwbCUUft3BhNZaBSAt+bekQPXW7lewpl29EVoN+vUjJ
Rrq9Posi2p/oTIZG49EnjEzImHVy+hblyXq8S/CGqKIaEaRrLdUMnY3WSdSpT1XO
XUgpUjxChyb/5XfiExDwbRagKLkE/D+pBOX48DePDHrzR/70nBBNYHne2fC7Ra0g
3TiZNiZPIDgaoRyGFJ0GGNLVQdYenT2IsbkNdzCOWpDYxLeTjut8G/kJ+YZKdGnv
49dEyj9xl5ewp/zTWSvTYJ9m5+nFDL8XKi3LU+ubaHCWo45PDvFvUsTNvCQkTjbW
/hk6s/t7evCMf327c3noZFYa1QvFrqSWhaWb5eV02jMxi9sCmquDrT7igl9A6eiN
fzxWDCWboyB6EdFJMlqjOXSPpEB4XpkyrJmhC9sOYVgqvt7TVUx2bPLKzPvRqsc2
InMkpuKlSjmhXfIb0UkbRoxjUTj/FU2sL/5WhCeNhHRr2a0VOgsTpoXSzBRUchjc
YCY+ermSm3SlBCVHJQJJO7lO5wLJa0F24B/S88A1yduXFx37QXBHxBfkwzWwYhe3
SoGd+eAcp0U3j+22DDfT7Exy+2fcS1rOht7uyyd+rEsZuWCXu9p0Y/VGi5R1fsrT
grQbQ9uH4RqP22JDWvOQam5YLgYoREfo+kp+9Uox3pAtwsUzVNOApU1Bfdn/5DAc
e4a2CWk/3cjhkyLQU+Spa5WqPgZiF6+pgQNPKmqgRn9pPR7K79SBdFGeV0v8M7EN
QDKXRaPp98gHvpqqbWwwwcMS0jwn2BGxf4Zp+c/PBdL20psE7UnE5Mp0/26GHW6A
Ln317lNKx29v3Vu8jzINgmg30jxpgoqmMMrmCuQvELnBzKHbajuwqO6pEIAiXjJW
V16rYE22IMzD6NpV0xGaKRps4+tyNk9e3nAWznsY2PiQFBeEP3K0IKymBUN/sBM8
6I0zZh9bAG8uIu+qGnv3bosSwbFKigq4pILJ1FBz/eiAuV5ukcaj4wC2KR1W5CC0
Ae5PkLeWMGLhYcKznED5BXOFn94zXTd31ReGy2GDWMaKgBws2VH0QpQIZj+GIbVH
F3EWWZBkRD1slMIypdj2wjh1nc7xpPx89QKCloDowpi2I7ufmaJA7krbUUV1xBAL
73RDXk8ebg9Cd2ywofOuodx1qPstbnZ8t2XJ/Z/MZoZ2vROHRp9zePpOinyEQday
Jvac45/wKJ1PNxFOfWcAKX8Gp5mLDD0aAlAcW+nG20ms+H5RyT691wDcwTDcT+GV
tF1UiU3MceSf6ui6//yeiIrBnVKOLdnb5JmDSdgmD2hHXPRbge/Q+EMFjMB9XmzO
kNcuIk0sSBsNu826QA/D9PsTDMSkXl/kYmNuLesSvHISG7eYZ0VIj8lcPpwLkNsY
kUz075vLhIEn3xnM5VreAXmnOzpgJ7qjhvhBLkz2RB7mde0F4rboGIqqJND8PPG/
12yQ2is2ec+zjTUfS9X+bKGJUNUN7jYMtNXnyD0A/V4gXPZRrD3+FkROK37ewloP
3SPgzhYjfvsP2RlfOgjsMoURU+4tSg7wQFqmv3rVQm9ZFcILQzJvtPyUg9Co97T9
WNaqS6FLgsElOMbJQUnervG8A4QNWtZ4k3wAifiicWaGhfoQT8OTfrsQwgt/JWbO
ah/5a44hMzyIqiiZPqR32mIHWa8R3wVfT0U4UnO6Nu7kPfkR9PQ6/gfigg657Ax8
ph4JKLAUJ3acJBh5KT+E/cDBqFMpW3Q3SLiUqeEpCEB/tPXwW67hw/VpamGNz0Fl
ztpl9U6uc7spV8ucim4btelionZXnpjbLus1PMezqLe5fFvvOFkKbaEhFMFdTJ3X
nCtD6nSGNlhPeiOAlj5x5dhAHN6Q/cHarbX+JrZKNzY/MQQfoyDXvKBV0EzIvYh/
kPr7i7Agm/UTxJBUIJHp85w5j1z8cL+YaNZXWcsY4Q5DTPL+NIj2jrRmuKMes/Yo
9L1tPje14uEzv4qvt4fiSYhfLdoccAifyF40SSQrqccIygIAg0H7tUjLv70qQQ1H
cQCkF1t+P3sYgEaN3r0rydkH9AjGlmQRNa+sesG0WBq8az6xu92Bgez1dKffM2Ef
l28DrUAKonwOcWA3rV3mqn3JRoH49TtsLF+T6XZucn8lhXftzpDL7iVPTjBsDnQN
PAe+uuab8hg0NHVv0Oy2eRL2rXuzphqWMQt45/ZwfFXN+MfzMGNnYLsTsOSXc+R4
e1mHvymygFG0W5MslfDRnYLCLRnWhJIJMTLHuMicZlYskGP+kJ7cVmqVpiwo05Qu
1mWxXqNT5M86W2PWTLOmoVkLZ1QpkMmvT0leGLhIpG+K9D26i7QjjOMMdJsbCMbU
DoLbJkMnG6SrkFqPnZq7IbpZJeAYcoVXwy9YUmdnYyuTq4SCKDhNycSh9QUSh8tR
9CURSvJFZYu12iK3EitYAZIJD/Iql5z1b0Kr1oQZZjliQDbl/cLl7dwoZaWJ0Giz
jCeWW5d5QcW+MZEsyr4Kq6pY4L0iGmsWpZK6K/x3u9SZDyn+wGoWOw0qm2bogpG1
mkfpU7gsMVUkcNM/mL1U3QCYLY3G6r0WVflN6Ye/vSW0Yg3RJ65/CrYq4xTH0AjU
LnaPActdYKlntYnr0KuTO3myPW07FxBqzyissFNiZVO3W0X0mpVlcB4fZ443a1aW
xSxgx9X+9Yl9RSgqnefTUxGbRe3C+qprv/p83QgMIEg7oaNjA3CCtq0yn3OStQ8e
C/3zzQeKi8RMdbMwqse3CQJ5dsrg/TNMknuF8CWjT+Y=
`pragma protect end_protected
