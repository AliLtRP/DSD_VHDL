// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:30 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
fz7FgnRMxhzO0qz3at5BaS48b6RKf4GPh7WqRTn1/8ewSHS0uFG96ZP39UR/OyGg
Qpe4oA53CqxgPGE/O4A0xcFOmpdkIG0uYR7s1rRxdWUqdMIOR5hKXQYh+F6V1fIk
t7HUYJrJo+sl+5KZi+QKrILQrXENCMwRZ4qBn3WGRMs=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 3104)
we8vRA5LK296mLPL9JO4uyEuq/qiZyIyU9KOgdPzE0IwnxgJai65ec9EF9m0JGJl
hU3GVqCiaDiBDZqnFsiTwIlKk/Sws0PKIkZ5Ssh1h768pD6pNQOJURD04yG7u/TI
LV3y3wESZxJv02sgKjtn88wwKi8616Ai7SwuItpSv/yuOaP5WQGVZbA5wPI1M3mT
aIKkbTxF0TzPnL0E7EpFSkFFFqB7Z6kzdbmMfcMIto9oyHlBm+eNe4j/wg4rOX2t
o2r4EtrhFLGQurRGb4eOuvPmgjJIodCjvIu5FQiAdPakMotM6PH5N8p8lpiDPjsk
1kygaOvwHsr219gru3wYyTsm2buSNvffknUAJX9qLVfUan+pxHDm6Z/qKO6qdhnY
n8ftBjXC5HOH214NFAcpkrCKfPbCo9jGOeGrbUHQkZlsqXnhV8OlremFJwHBI9h5
aYBh4flagjjfN9S2YwAxeKfmqKPMy0BLPuk5rZ445Ti7bpYKbI73zyZM85VNFLXi
PCLPpxse+0xT+iW7W4kntAAVW67RSZhp+fWfE7iwmDXWh9llNu+n0NX6Tp4BL+aG
FAuSdG6Jy6ngcwIFiJI5XupWRO8DCL7DSUZGiRNNBVzgrm/Oyu+NP7hWjnXS2/um
yx1G4VXih2JpV3tHhKFYbUiDC8Yi7ApSLBUuR+7ZgccuoYH+G8zKsiy7OYILGaol
2q0J2BkukCL6g6fiG5VXSm2kMpIChoWlwDpxgeqt1EbloqMtPJJhBeS1Uf7HDg6k
NxHP3vgbNoK5hvqj7OZBX6izPdrJXUarnlkuujS/n1PnqK84OsC47FtmTSJPQFmP
q492TGTC81HwxYE2TMMpQDZBMNiQ5X9Ae8oUfpY/8AXZntsm3o1bDS2cGzEOAPT5
Gq/kETlfA+faffqZ1nXrUClFJFs9+GR4vYhvg2PM2xWrveQ8Ss/pFSAJBcN1EAG7
aCCxfgTXioDlUs+NQcb5P0KpVvGV0HWKlOizjRfa30HyiHDiO8ODn6QBZBcXcmMc
glTDrfjkcOv8/fkx1PHBtoHFQne2l8Eb/pbgpPWu8E4OWXs3YYwmByHnZqzuLPsx
omGkqd5ODsFsUw7KuoZFJIQHHz5Dii1kusQxE/tqrYqxpkop2eLrj2ft5b5GwXWU
cBv8rvt0g5hGNyLkGCXwFtnXMl8mEt5GxdPuTfQnUWA4N61bXzEVcjGFxBnjO9yu
HqwsnxmPU3obxzpyxMDB+2lwNQlCGeV2EAL30epLQNQII5+0vIvpoRgYfxs5AQCn
r+HX2qoVGuHD/QCKIj2t6W5POTDqr0aM8scMCYYPjqHXxNJBID0Dz4cjPjdecQaM
FXjf7gof7jX14qydUjF5jmbVoxb6bNsbiYQQVuaPP3QE7drB0GJ3rQBM/rrrZDZC
G8NYSOhPDDobvK0GDz4I3K5VBJStYPNbb4Gk8bVf9KEqucff6g0HF4qKhbzW/wiW
neHenyDMKUjeAaG9Cx3xOMsHCo0TVMC6E3Aq/ejrV9PtL8xeYAq/vauN9wnc3QUq
jCRapyAFh9nTtGg2B3xlJ5kiAcGoe+Hdl02c0TatBLPc0TFr+HfKTtBlIOyzDFDa
3Ujkp70qbggrPWLRqyhui05y84UIGrxBrL0JnHRlCZofPn8NvRpEIQfPiWpCqklF
/wWkd5Iw2+REZ63KH+4cNgkitnsfhbjABUqKbatCYsSk6jTKEOUin02Gs0PdMH1n
1zB7n7MJ1WYvetmVE31oeSGxk+ZSaiZtIoAGkrV1eyg89afcaHivjWOU/OwAYqy6
zI6gVqtqhOAoQoltazPaHJc8wSrcNL2CyN5YEPS/GES3VEKpxVYpB0rgdIJ2/kfu
s5USPxZDdj3ZT7uHFTKHliGBru7bCKt/wsZcKl27neBfOh4cdCbBFW9CHyxYFz07
R4a1qPpOkBMZjfbmBADrwBMPCyEhk6r7t60wOW+h5c3ftQTQMuKZeY86BeMhf4Oi
LVAEPRAgZuNXZi/owh5cJ1Hjg9F9WuEIlvv6rsS9u92q61r69+BEtrPRuK+KbpeS
WVYz0NNhKAGygVAiJuRAqHqxKCpZniuxqPnNoRFm6216CN87yaAw9Dz9U2iVMVPQ
0GW/AhJwdw1ZgLkk5584TuANPps6XEhmuEeJfj/fmKyI+CJguR+Z4cuoZ9KLo30Z
0pvl0AKKfgk7gkkx7aaOgEfHvq8u/BQ+kOtMn8ml33ZcKQQwrIC5d6HSt6g/TLQF
T26saES6jA+6mcoZi9iSGWDLk1yEaHieQAxG6G1+K9TmThyyRVoKe6BrpEQrXGbt
7KuhsYKn8rjG6FrYXpnK2Ad+AF9y0FY/TR6FkHxq6BFJhekds2cJx/RrOVg95Gp5
aBAmqGHzqcfJU5FLSViA3haA5Mtzsgzw4WunaZOux/zNEGU0KCAyQ0+pmyBak/7/
807TUME8+GryYpiKH281BFekg0WlvU6hg1v/4TCQPFB3DLR1iBrLBn7BsQPJbuq2
b0pnCTYcguL7YauuInxulSUnnZIENd1cP6NhzbBJaTCM7foslT1hUpMxCSOf4lBC
5Gf4osyd7GmQRK4LEl26e0xs7R/CLA61qC4Fc/UtPok//mCjiu/A1HyLRKzMbr8G
4WfDD0Vc88291PwS3xhw86hZPp26lsjG3/cV+PecTnYPrhx1VGS1ewmG9kWUkXnG
7okum0nRcebWFHL3FTSs0tAy2c+e3/XzrmzWZEAPCnJm9dnbOHqL+EMfdC4Xs0bi
Ivor3avP3z9PaA5+BgA4yq5j3U6SyTdMeTcQiADmpv02NgE2+uXymkThpow5ZZOb
Il4AwnTEipI0omlNeeQObVLAe1vr+zQYWrg/5/cvdV4DEdqgCXkHbqd/QZJ/elHu
6BzVh+DdP+4OmDyuBAm9NfNv9hEq5UV1F8u37xnIcbItsGHwmoxsHY0lky0kTFsv
mXTuHnjSjRMpJQ/CN9ybwWtu0cshheJSIiMAs+Pdhct8rB02+di2GDXmHmQNig7S
MRvPeRDwyj+llMq3iNLtk6D5bY0MeTlmAcPPVkyopffNwoawDGFvvxMlWD7czl/s
6k532poSf/F4FlDc+TAGMD/W1UbSNsN/JZ/AgATedR/SMAwM1rPYc9htIpYScqI7
r4/2aG44800ltoBg2KnNUNoBb3+ApJu3wVFO+0qZluVoBEI3WslABWxchtuRrZ+c
6XfFJ8L+bAhajDZXS9whw4CtEYYY8GWRpW/ExUZiLuF4GCv3Q7FlYToHIQwAOIkC
lrojFwv7uaYg6kMuYsIMFdHP0qCEKTKBmsOeeKMCXagFRIZ/5dDqBAEob2ElkAzT
6LXEw0zD3AZjWfYviqtjyGGfTbkXcpaSVFl+EMbNAd9+7+Otv6+zVYtlejosLexA
DeC5kCEIdSl/H+AzJW3Z3Il+aqGmQ3JgJMx5jw48uEifjzCsyEyHai2bLJ/Zs7gq
Jk5PggOvg/MbQe4wCInoSxq/Q56g0BgDhl+JdBDXr4gMLZDEQN+weKg1rS+mxgVK
TzbxhZUqYsh8N8z7DBHu4n8/bOBtgmMXJwe0dtAe2r58+HrylZTUIXZ5c+aoAcoV
PNxvnrhD1Hh6plD7/LGV07WkHgrUsAAgi8j7CTv0xyZhtI7QLTrSpHb1JETmJ4z4
U3u+CwOeTIsWqJdgc1lzfQxGQdN63cngGJ7TaKVTHqq/cLYkEdBZNxMaQBmB0S3r
9xj1ZscW/5Y7qPZtYMqinzlKdlGPiDqoOKUVicyks0z8r9/Ge5wJ1uze4bYEPRka
WX5hgW48SGbQxPQrmzyLAENKfsb/w/cuCkcGeF8uGL0GxIOb63npg94fcoEr0ETZ
WuJkInVyKU9R5lq4gPY4YH88wqcXHDEPnmAVtkSwghyXwdZlDXxSYSULO4Wudqro
HHvYFBnUR8PfIovC96URFsZtz/KyZEATnAVKVYwf3q/uG5ct9xQ/z5d7eZnziofm
DPJO6lmBUlpiYjJ6aksJnniYGjs6D4pnnm9yDEzcOemMw7pwAUS1ilKKd7bSWpA0
Aa6RjHctenmtZ7zwlUgyQgTVfaMP72KU6R6nIxkkC8L+GQklDAiIr/bWr2Xb4gRc
Rc4fWcFfysfvvHbmOx9lJjifm/VuTNTz4d8AzWwgKb8=
`pragma protect end_protected
