// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:35:47 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
GDbzdpdjpPSwnvhTazqjN/FX7rHVh+HRF1qtI6XEOyGNm3Tb+5pSbQHw2kgSlopa
gKlCEWx8WlNoflFeqeXztE4aYuj9fCQh20D//550baigeuJpTxn1pMWOEu9vEDBU
2b0pcjIcrzw50qTSG/j3rV7sbv9s2bb9UBbmgSkZtXQ=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 2448)
ykSCVGggQiogCfZLmfF5hSUbmZS87ZqMzdfZts3NEbOEp0oV8S32TvpdY0V7llGX
t7lQdDOPuA4o1F/mCHREft5Vcpl0YKm7O06L7st7njTMNxll+P78LCQnCjuQ+eWB
3c7UM4KckoRqNF2VKRbv0iBGlS48MQPHSJNT+bXLWRJccQoeWxJZx8S4EAVEA075
sNoj+dxuMbrEEpr8DwZX59T+H62g/PHI9HGhyZJ3gm3uzqBOYlVuQaKRx5KhO9L4
tdgO2xDyR2vh08DCFqRZUBUJPzp81dai2c0XGh3SydSEeBaOYbHOyvEsvVVS1Zcg
6Ba1bIoaukY08mRbbCvV1GMyAWZ5jDu2OOFzMRWmw+OvPBxnHW9pIEjWS/qWBVgq
U9vJBgyGbtuFj2gNDi+0xtI9xzc9HC+ljT6VE5o4hCGtZREbRZfaYdynICdwZPEo
asv3ltU3ElVVz9+xo6uZOJZsUWpv+NBoUPzOJvopAkloucOPdg1hc2PJn1tNmSAw
Z2uFRm1SZQ0blU3GapG159dLB8s0JZ2h75t0qQQOBOdpR2RCT7pXFXfBIIkGaAkG
ru242E3cO64YFc+xKMSlUwLVjZOwHuZJdT2/y5OonVa+e++gJLXk1q+h89v7QZzJ
xyT2Or2DSdEsCbAPe6obar5IxtVaYEv/zQYxUTQSyzXqFbYrJI6hdvn3O+g6eglH
QEQD3BCkP2trgy2uhs74AmIt8gQ0EGDt7qZfSr/1GKZ6ps5uv9e7Fn6oMGPf6bH2
ZqkTOpPBD1U73qznQ9ctHPVQ2ZLbRP7AvQ7A3b1Hn2s5FlkibCYM8I08H+aysHgY
tdGGtju4yqXtOZkgxahW0KBEM2UhzlPo2zeyW8BPCSZgbjX+LLbdlv4urISrtMaE
hJX5wHVysewKaKjayvcDn03VB0WWSz/EGt5AoFSjmCMYNFp5xE9smuWcdB+VIfwj
qOb61XW6wysI0UdEy9RhGJYd3DU2a8TvHGzDwvknv27O8AXPV/j35FtOHd3073T1
eN7n4SPnAIeus7ImUwoE62VtalHiCym4saf9Zzhfx5Q1udHTrYNKiLvvC2l8L0Yq
kmabG6V8AWqGFl2WBo20ULAfjZHg2MKOfxEoVRccyDac6qid/GklrZQVr7lqqljc
BnrtdwzRaw6jURs2yUEWgXu3g3/7OVd92xDVnznDVD287uOmmj/WK3rj2cL93aSZ
82E/dfXVG1sw/BBQzHnOKkUuVis8wT47U149YRYAY1oz5znMHadsHKRvcLiXoSru
6Gso885HGXlsMzUy8kI9BNjfM9h7vySEr16N6IniolhunJIo4AhQJDYacqvkSmpc
6fk8KXcqIVxMvk02A56w9l7/Ahs8tRaYD3emWsy8Q5vax3i7aRG717IIh+L8s9kf
LI8UYudtmknXNNd3VlBkrhxB4MtBj4+ud5g3JOS5kThhUw72L+o0XREv71ZbmM5S
pcjBYZ2C5aanSSSLQjsxEAS33U0iq2PRJD6YsGYHURbDa30CAl/SmWUbg6/Fg2aw
H8L5S8X2niIsq3N1+ni/RjbU4LZIskk5Dyqb2N/COJnbMrljF84Wz8YIshNj4wMD
Q+s8qPYNcfUbJHvcrP2rlGSqqQqGtXaZChMb7+A2zsZD5TLCq2z+jK09myZ02/5h
OB//yCPLPV2icy0Zmv2pX8uPtZLFYXR7AcW66ElUINHKb1WrvBDO9E4x5xpGc0XH
kRFalSKwEpGjalGv/N9gAwFWSxGMX+mRUpimhLoY6P6KHtnIWvrwvawSUBpI0tur
eKIqKa/NenNB+3NUMdy2aiKqW7fTlCbCwNm11QQl8OJRKPdVr/Xu4gUXIW+zF9oa
x/se6eLal9FOg9yW5qPhnC8x72UKYVU2yjf38MeOpGcT92GH7zelRBSV/QRTxbTb
GDGAtuNfLoatCGaf0iDxpyBxJ5sPk8AlZlek4GU7tnc8bMFoM57p6yIK2s4sQSpp
uxZXa7sLnTZBxDLGRCR3pn/sglCmCUT2h6cH1HkETFq9VtHdezBWkxw6rZQwN4yt
wNCT9qJ7KuQurbqDf/7ipRNL8ypuAlkQAtBSzBmAuRWaULsFN8isihZq1K/27wEb
6t5q6YY43gc/sTaUwezpnwZfSpQtn1biImAC12pof8afHMvgOVnz0ZBX3JfVi9tD
4plBVtmV6doHbXbN2Cf0OTsXBcx8JJosXZm4QsCLZuS4IYvU0l5neT/8ltbv1oXJ
02O4YtXbi31W2yvDMkdr+EJkQ/0AYcCTCrdMnnrcqfCZ4TrOO/7hTCl4IzmO0orl
lwCX3rMgInvB/DPSY2+l2zvHnf/ty4O7v6ufiSmimBX7o/ceIrmIiE0Ig/Mm2tiu
MXn6Tyk3vItT4TaBg7SI0J0ZgWnQfKc/9uxuc+cME+C6XJoZWDdPsnVR6OHRd3CB
KY4RyUOCul7wXN7n/t9Ez0Dl5X3MYTJ2Wk1ZMMZJSJY/3X9+lBMxb8rjbfMvxHoL
cdk4DFe9f1wGn69yj+xvHKb+eqkryWTE6QjwhdYiqcWWq1YuxRiZYIBHZDgUCYq4
4NzVb5vaY/EH7mhGUxiIzVIvE8A/wxzR4nNoCaj+mp+yv+Yo7KNJmvhRWxfoWsXy
1ZnvR+yn8Gckop4tG2RDArYCCCLAvac5yb5FV1lbDj5cVGKORTPlCh4yyDiTXrzB
Q9uk+lGbwKDe3sXexKF+7mug2Ij+Z0H9BTQjYEMRsqGPkN8swJvXF4hFXz7wrMCE
2kI0toWWUF3xDJGTrDdTjMUy2bzMbr8y8/FDr4JS59NH9J4R6dWfLxfD+ZP+NSN1
U/r30Oh/CmvzUQHZgoh7buLB0McwiOyi1LY6b6pCPaJs0CxXgsW6G5NgiErEB01s
P2uvTD3N/AaMdGlDehB+OB7+gweoL4aSznKh9l48M7bhYMJ3Ktwlkj9XopaZXJDV
AP+AUCxZFrBp7SMAwiXWYkVNRZ8vZ3q4GGHpXprzl4jpZ6amybhOAoaLLhttoIkX
NGWh+3NhUh+7xV7tCQ6ZbwbmRzaMqMX4o5okP0fT2b+N/lUNW2xkiyVMz9zLh55m
b8+rlPEaGpVEDnfO7sD0V/oT7ptWxqghtqYwtJ9qZA4zN0P61xUCjYsiTAryk3Xq
dT8MbS9z4blpmz+3bg79o4Y84vVWmXWd9duVjHg3QPpQwqZHH8hr9UebFdP+7yaP
43fbZ+gyYAjoYAn5o+hqXfR1e3F66kJLR9Uvvi8Va6VrBO3nYqCm29bjP+eNUh0r
`pragma protect end_protected
