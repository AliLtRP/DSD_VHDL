// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:17 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
r40uXUnUAIAltpgcOI0lyORCn99uMs2lXY0CEN87WcDxzbzN5+X6DqIn33C2FhNh
bo5XGvN6ukwylGNrtBHQF1ODeza5F634slkR3or1uInClewnKy6vfN/w/4NdjONm
lW6iMqYUBdhD1kBb5lLKtMATkQ9RgklSCSNWSL3yCrk=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 18912)
its1BE081JgpdArLj6DzgAPYFyKPvUxvSsnCSkxTNaSVj9Ztox+4mOZ08Q705EUa
8Z6mDDqKg0u4ib3EoZmkcjYZUxpe7gkqeNV0tBEIR0rYqgFyrunffRpaLAOT8eaH
TSvN+ip7+osHqtZ3zdFlgtgG1Yb5gTbDjz1cb78z6Uw7UlhzOvnd/PUogLiQpuoN
LLJu7ibQNoMil/9tOEZ6/Et/xZSEzIkfPNWG2/HfhbDjXzMp5lLp2ZYFZ8diUqYp
zo+khkwhx1Fq9nfeAup1Mnwh8/i9BRGj023sgCQCQ5TVrvHodIqFCBEenUMqPKkx
gnPgks/TP9bYA6WUfnjhth4tJTRkIVEtzvJqNXCKylFxGPr1/ca3zW/WJX8woAMm
PwDrKxdANm7hPaMLF+lRVo23qyarZm6Rcdr9O8Fhc5XN+zWO7ukITzruN3VwXFTc
ELcjHkfh+5RWd4WAK9uMoWhWHaCswYJyaEHqP6IErp18UXQqqFo1YEVHA6YdZxkw
5JF1S9gCSCAVuIVqgRd0SMgsz4Y7x8cbHxX3li28DY/PnaToRLA1GgAhSE53pcX1
MJAAaxaPXcMmfFO8ik3nbFFErcg4HHVIOgb/fXA5l8XDU3v2uE9+JsQmBtowmxYV
frHVEXJDMhotr+34XsA+EzfcRFLK29sNASsOy9wHEBBUYSOrzboIY8ahvnDtyylt
9Zu3aSTOs9OQSd6cz4Sd290tok4uQUjD38DhvogkI8a9niC2BMIzXTePoZyTLvFn
q/5cJyTWOZepyXBbKiJ2K92xyG0sr6u5kPSuYRViLmM2YXH+UMwxzaMTxZ2BkPuS
88vMQiDnK8YlysmquvjEWPb/3irJnlK4Q1Ej9+3MYmPYJ0I46afvbsHy2DvBLtAK
wnIqu+BJLOQVvHMjhsdnnXJooDycZUrqyD//U7ZmON9/vAXLQg9sFgIpfLwuNQvV
Q4KLSx+EqrsSC63mvm03WeTfrHoOLXdVoYxdryR4UirZ2/DJ654i0yR5dgt1byhH
xxD9agrmlAPDXw6L02pt34IcSj5HRKj9b5Hwu8i+77jgHQ94Vc3ztHPBMYmpDf+C
hXvu0ZWwYBlGLmg62V46Mmtd1OzwTZo8yhleb+AHhgOjBLG/8u7RlpKXLTP9+fwv
S+FF8Z50ym65SRJSq/Gpy7HKWJxOQ3CdHstTSbnAxb2mguzlql+s1eNsCf/UmZyV
wlUIr8FSm6QutrwgDPhQ+B2EVcDD7oEgCO2k200rmJGA0faDOm6YRypO7HxaMX2r
9p89guRS2lRde23ndy+T/Hrcf+UikwAaxu1u/fdA87GOOT8nxDCXpAOj/cC6MZlI
2uU7DSt18RfpVuotiRytRWgWAOjkYiWpIHDk4RQkjKIZxtiMHC4aQ38pHOv2D424
oPuYWNc8JsOLaVPYSEF/VxlgqBunN6JkfRSxBUbfbFrtPCGkwG9B/Kyby9mk9CN7
4htxcjmfDM/Ch31Lsb4orYwEpAT5bMEOpbm4zrM+Um9eskB6GGfl4AZGo+LIkFOr
f8XW/01MzmSKcS6wJET16tc5nEawv3WIwD6JYNUZQYrNUbTvO4Aj6hRNYCEUDAgN
tY/XN99OfEqvTCW9PW/JkY/B/O74Cnxl7ZagecisfN9YOVXoZGwlZCOyLwS8vnFY
zM9EFrHm17K/vYl/537deT/EKHUmixjcjXyzd/T9banvrzkkq0YBwAtju9ntzduZ
ZEXWdSqYUpVc1efIEC3teJ7WXdTykFxPVhCJrsRSErO0eaF0aeuPCZkpqf1UVUhO
X8fqZdH9yO4MSICvTwu4l8j2t6qLQXRw7HEPzSLz/hfburVZjCKmldgT1Ot4jpXg
kW02L898VPkscthRoRtALKMmazwbh7wj1bwusTQNdxeflXcbNjWe2+q4ZAFh0gaG
kJUfKGQGF/cO+AFT/yWRPThmj49jFIGf/0p55tZdNe9jDRzmifHFs89jVW1DOgcm
GR2l6kYqn5XYwGkHa5S9kn+A4EV7Pf3XO+gqYrSxipK7iehcVA0sVGZPXtPBMfkT
96ntQ/MNFuasRdew1wjlse3XVSlQKVDw/pSxRlYDzoMr1NMRCKZdxwsWTeGJKCTd
FJgWUA/oqLQglKlGe3dqcFVUHnVgLMOyjUa4h3rbryt9iPk4faMmiEOYWxTvUV6d
55OdQADEAZsoVwOa7TmA4i13EF1o3GxYoPdJfcTj+8L7JgdexwGhiYYRuBnBZejw
5QdXgxX7vdTHmZ7FUIvotZIT0hxICnMKGIXw2jB1xoa7AfwDLXKFY6nQjr/JrmcH
azfQEC5oB4DlmvqPJfipQmszINBb+hK5o/LqN1eEZhjXwmGOk4nso2RTxSLhUirr
N2PTKaAUB98RdMH2ZPhSJnkei05NnJClRePr3h7pAobBQvec48baVdA8+QJHIOa5
kpif6ZMJzDNo0ekzLAZeC2AdV6ehLFlxdfN8RyReuIt6vXM+rHQ9vf9z5ZztFLyg
WURs02YuVZFy3Y+OH2k0VxVxQ2ACy8qE4n65+e2nMt80NILetT84VrWjw04Wye1R
FYUeOBFHC7qYwhneFx6RpbhflW7vO6OoZxtmXAz2Uww1xu9aSlcfAQHOE70KBWWz
a7CK//wtJ93zDq1yiqv9u/UWKh5pUJID87KSfUFpBr3FazypiBKDO6oVUYtiFk1a
zTykTAMb5dfehZzeZ7UDe/b0lJRPF/70012rcvZqA76YekvdQiGC3+V3M/cjKr8I
DfnMkyhr2FCqFOdk/JTqPVJz6U40kqnLxwH4uDNNgF0FeHDMGuoMChWVFWsiwJs1
VUxPSkGmxZhaYYFZtSMYLQ9IW7hqVmxGOxmeKBF0Q0aif9qrGWVXNtWkUdswUrTo
hEjBtTd1tzynLwdnTO5KGYKshsf7HWM7RzJ7nwzjAOhMLBp+5XnWljM8C/sZ5DeS
01LD9CugF2OX+ZtaYQkN5KT+umD1I4o9E4LjkR3rNQ5RKcqN+7qajidAC6mGHqlF
HT1ytrhNeJ98w9u9mfil0hLL7eGBViLbWJg6RgyHw79/noNVy1ixXjFXFsdoifo1
fMXeL28L/YoiL5Gv5lAENJKKj8q2aUx1xWhP5/WdFzXWTHICLTN0eeGRGb1P/HDZ
VrdeH9LRgosHExZAxP+LNhc0byFcY5u0dpT9Mu62zszRc6A/ZnbQLcYPCBI/esGh
i5vmbwLSjS1QX8U/KswCz38MhwvakXkX9x3AjoMsotJN4eXBSwljJ7Q0mJ8QBNga
BHomEUoNPQ4eP3tCc1Ralmr35py9NbCe8HzAi2ugXvlaRvVBQc+ANP1z0BxPTq3z
SpJQqbruH+CJYwoK7cJLpXU6j1OI3FqF94/mExBryG8KyDEtwVLqzwRBkIWJANkJ
nysmUs5C8B3vUvcaVlnyEpBQgplccnfl4UYsoJwIiW6R1jHbbd57k8MV/XrfdJGR
xgUkbJk/E/hDIbS0U/zjybwKYUmRitwR/TRKQ8OH0vhXQoyx3l7+x6KiSIximvPr
clPj47BgaswQzcDISuSsRtTY2L/tBDBZliCu2ICdBbGUBfCLvLTYkg+uXra2JlmH
+6uOWc6vQRgiUFLbkojhMWBmTJv4c6Fk0VKD+aPO1VSGPpIk+f+AmwqOUw/5tS/q
jbt/8GQjhrPEGqIb1LmIPX3d1wAxDQr2hh2192ep7YnbOB6z8rLHnJepWE+bxEnz
BKFlfzJCNc18sptd1lUCXkYI1QwcdDccbhgFS9yqUsr9hF4oXDSy0H6crenSIkPv
jkaWbkwDY7hiZF6UPFhRirwhFbSTDTRdFhUZJoP5cXkYwSJ1fl1Ykr9TkSvoUAhQ
MmF1RLoeR0SM6SOLuoi3g1XOPTRWXZDKXKDiQn7tRd0ggLXdQXGTvc/RzwdpN7iY
dyASIVYk71TTbnezv6eXHj6BdzweXCJ3HanICLHEJB0q9/drwCCCjTL+QesnLnEN
5rv0D5hRbfQDlHJt/0OIoz7GHZLM8xVDeYtCflLSro8FpMOaF4ulg//xoLjUJaOG
T5vEwu9mN3boAAPUnFk+SnxAxMg+mv9+ejsakOz6VjO2AT28IsK1xkfLFhwBwils
3wV80oDQGWLQcalqcBouNpgHxqLBQecqeiRsbDAW+/4uz6iaQltzaJ7MK9AYzPuP
6T4XnderF5hjrOMcWBRWxSW1Q4MUShulup6nabNU74csGXVSm/D7yeBi7iPTv29O
U+sf8nAilhVvu8BdTXoO/DTLY8txsYaAXw+QRBUsclF5CYOSIKMmL/Js8wMlGnUx
4crif+xOnpDk9l4pOpXznHehCkX/lC9iSECBDuRDDShJdEAiTFcd6yWTcaCJL/m1
9p2zE5I9bnBXLho+zvFeZ+Tsawd32+79xt10AHx8Ixq9oinE7nHtLh0WFVHPY16N
rcucBOv1WXQW+od/KqBXzCv3SQxwBOS9zyujHK/cIHnyWgEhqqgx34pITbF6QiJp
scCt7ixe1doa/Avd5y48mmDpfZKgMDVzVZOZE3bPY08iDLc12Ma3PzLrW6J2RnMs
ElGigCMrnrebcHKWduFVmCxe7ti5LKdHRyACbA22hFsvbPMnKvdgICU1sRsgFSNL
JxDX+UIc77BDKNe6a+y1W3YCkUasW2OaoHJWBKHheqrhhHT4bBS/7h1cOTviCr8c
tuIzEXKrm6tRzj+XXMDEJq7LDgNFFbQ99Z++lml6eHesI5WFo3S+jUIsy2BFsbnE
SjjMj3+7j/rFFfFtl3K+JHYOXzXimtMi8z82atBKM6zgrfDQjkNIZcDYi51r+nV5
LpZ4zvTE4bFXXTkhpwj+sU7gbuuQ1BWmcgqvfCev2zC7DHaWru425vHIEx9ucRFr
c4PkA/cg+ePntjo5UKy+wJRnYTeXV4XtVz+cKSX79XqWFO1b2QsQa5yWM/XCZAfB
LBDD6OOq+O9ZTEfPyZI75Oc5flrEGsu3Q+dHmzggt/3ciSHYhJJEKIFTYAp5XFQ4
KwCnlrEkrU6uIS9V7vEUrur9HsPrUU0uvbp81XRsPquN085sk/aGb89qvR422D7F
JWg8hzbGttVOXYsPNzsKKjIBvCqByUMsrQVa3W6ziFjRV/j6fJsA6EICm6x2EHgK
hN6/l3OZDBxpwiLhgCxs5DhU5nmuckhzX2DpfPK7rtRYjTiZ/K1xn61pl1sXLA3m
cBU1pwctbQ5eaRpiPcJDZu/KraJWiYLkmu0ilGn6Z6aMrLzsFFMQrHtz+rN3gBzX
8D0tluJ+Z+w7k21csaVRQJ6QDWem6F3okr2hgk7uIj+qUWI6ziDu18IX96nvk0Wm
/iPOvMsh7x4ktzwQOQ1fgUK4SLR1KFkisxkkS2uLX/O7mFZ9VTvPTE9geaHLz24s
vwYsiQE6itiOUXk72MXTZAO7HCelV7MKG1XPxDIgcNty+W15KlgIPFUaVZn0CLnb
kImImT3HAAl2ctohI2WM9pdvTGdWWkxDPMTARFBESq1EL4TkPipSRZGbC0reemjQ
IJuk2obLTmlPUE0jbTItay3Buk5dyToyAcfJk63NjCO+WdW1XWcui8SwljpEyB3g
FRa4IkDCHIpdPdnD2dlgjbh6WpAgcrRH4LoqrAVA9Ux0ds+exvG4IknQQ/gztmJe
ZXX+DaisAzPSBYqift3s5eDh4+6CG5xxzhV8Q5wyOzLu92GaXPP6iXFptK8Kpi5R
xXYAyUqCaRuehZ39fIbFwWMt0AcouslpPAR3Hy9cTqYQ1LiKBq3uGFBTFVDpfHL7
WApjp/woB2lE5LqFO69FS0mXqlivDl3vnNBihUwYVfPyEry/Fxi+s2n4Y8lNo9w1
lxx5OkhnyvSFi/H3/kljAEyb5ImzjEhVx9A0LTRIA2Yq4sAuHk9wTJg1cN5IHwex
R/JU5F7KvUhx7q9CFoqf6RzZccSwmzmVarCaGitIdC8n23hw8ZbfAZvw0eD6dAt6
9m5pXoXTBaLDt2KKc2mTQfPG+kVHruPeMIYsRG0IYzoKiLsKEPk4zLvbK0lnonDE
44gh/EhESZLO81GbsYva9GyqKRdnTbDHxZZxe6q7gXqHtqCwuzRFI0FQ1YXcS4rU
HDfklmgMNJLRzj2jN6gzsYgR8Y7G0B5bmbWUOzqbrnA7a3sBXRdGg178ZquZbpwN
EDBX+GcHUCjCXD+8KfJHUDkxB/9VhQYc5NTyDjatNesIC9Oaz6wZozP4QM4OpBAQ
QZAkHpI6aZ+xJUUE0i1YsGtoJGYTZPL8RJ9EP4p2lIQE/wdTRZFWyl6JOYPQXDXw
dudMu5iFt75taMvT8cQdyLIWwt+5GeeK2JpX+Ezd+5257Wxa6NeqW2/TXUJMQYHd
tdM8ERH8uDBZA0MeXH8S9jiLdTJMLNfzD2lnPYcMkTs0GjQ/oLVolqMBB9B8syYn
+8/T6j/iRdvaUKn3Twl31azT0t4dQPbfYvW/ziFnVxZVEN0/H5H6+gf6tOb5hCnc
5DAV8Pi3Ah6y74pMezfaYSpk0F3nerWqqh9uBIdtqmx/J7FA2RsW2q4Oc0knsCM/
9lLgbhXvK5qnvtK2SFiG0uu5O/STH68qtiGwIut618lc++FrHIhEODq14GiJ3qEx
qP/94UJmoN/vwaBHbd+EKz5Pul3uHi7gi5Chct3IsXjG8oBV+m429U1pUJLdxaBH
DLmEaL+r8WPHqylv+DoCMN0Xr6xLmt7mHWEC6kNHNbt2ItfuZMRqZtaannWOuIOv
I2xdaPuNBJjiubts4znoTri7k9iM1g2mFqNNhjBLmZ1UnnnIiuNpmdvgj07g9/CK
Mig15gtOEHfU2CKglLmj5RpQrg3Yn0lYoSYhjQ7Pa1QBtKQJ3xt0xG3clsoLmR0T
3TsmelAOWAQEuLkakCLCdf+zzi4yF4iwXaOw0nAu5rJETdCkRcsaH7TLzo59ZEdv
m91scdmvecLrbNSVPm7NSzu5ZfKHpF44ZlyWPK3+VXduq0bILtEG76R6hy3y85fx
ntivtbTzMQeOdWnj2l+fYiwLswL43YITU2Y0DlRmm8xn9acoryk2liEqShqof+xw
0W9BXvxSBZrG12BBXknJSds6kIwK0TxK89cCLKWqpOE4sct1nWLkbHVTPLEMBtjw
UYVxrGIWZdVLtPQ4HOZoqJFaP4/qiRXGaPzPPKfpoVaXNJNudxX/sWyIQ/0LIaXU
3OwBBFBJKDabu490TvdGQXS7oSa0AnyjUFYKkS3CznbHalPDSNbhAQa6LBysYH0g
vUbuvLxr3f+JSz61GRZWsJqS079r4wp1u2XTfXeLc9ywMgnExotQBSnyoHIbwkZd
gipkeTypw5b5iHACBTD0R1NBaB0thsv01wp24Cng3csBO4BNxpRcGhlI3Fx1kY51
ofIQ5kl8ZKiRXUtghmRxucX96LBA3b4eo4ItCJoFFafLsv8hoKi40d66rxBxNOHI
njdyqR2nCkOSOY63OGaKbVVZytMFcSrGPh1upG5E3KQpQW6tfmgjBPpft/RWK89+
IWphjAxCu+GKetdwvhZc4mP7LJ2a8OUB9Ca+H8m3DGlagr4bZ/QxGB3K+cErbJUN
L6OPkamzOv79emrQGrXB+oLcpwKFupA05/oAh/N6Z6ez6zqwLdLwk8xrlE/v06w0
nTNU0AXzo8dh4f5GhVhEGAMk71xMeDK7RdLOVl4Zc6eV5LkqAZ8wt0zF7KdLiRFB
yTERcZKiR9NrJmAuYDuDW8H44X4PWGuw+C6my8Y8EqZz2p5Wt0FNdrz4t/cAcV1T
k0c3fOucjTzOeRxOb8oKjxL0HYNLm+UC5UFIV7cUVrl+ttkQkczvG/WjZA84CxWw
BNdIlg/LnbC9xLqRjBKZK1Tfe8uwgJ2cw4J6PmSWoqKprQmh6HS64LlK4k9m2jPO
mfv4+xYMngrlc8WQb19fSWCJS3aMA7cnpdHlt0vtoKiUG3I7lEZe3OCiGj+DMhhs
0pD4dg3mp1A7e8V7YfLWOlb8r/u82dfJ4ysoL33GiJGoM91Oda3HLrq6dK8m49Sa
/nWU38gCCJT6pdpw9Dt079sk49KJH2ZV6S2a3PtqfAfsErShMAOBO4BkSuWrOItx
SagrQO0Ndj05RD/8wtOcZb5xzB2XMJZNWaM7TaH7qtQJeDE0vlYBIwLx8MJdqSVa
g94tv6oEwCjTkkKxW6mpjc7LEZvKh4CxpDlqNyUa/bKUOPKxJIfmgMrW2StnvemQ
dEbA/pUXctTTPmcsntjhAbhHi3NNQs79f00H1qWZn1OTklSEn6mpZXvSXZhUInCb
oPNm1CvJiBfWBtILhgMMxg7GyNadLV3AGDIN1zt1dTDOCI3klxbCPC2nBsxpO3np
y8nphpq3pqFDtegOe69HleS1cHykUqlgl/QMM7GAlEh2TYXjtGjYh1ri6zI4O1NY
CaJlhAKaSkbmBMDSQqQr/mRH98if8VnruNK93ZlFUHg5bjCF+cTBLtd7CAE0GvNI
CClPhfpVXVsOPPmauyQkowVzoBo9hBxTomoCXtLJsxJRcIGb+EIoT5U54AaxtEkW
KU22+hMHhZ8TDOI9cgnAib+eE5+BUkJ4gU3uyYICh28AGUMDdD6CM+DemCC9CV5n
YtXkFmbMC4MpvzX+POk47tLcph89ij0aOXuBzOpxwP8lD3RpDvm/GfgWLRF1InRf
9uMhqVY+uOH/bodtibfHWzylej73fFJ2zYgA0DnQbewL5YORhAlX/9f3N0Efo5pl
9BmCwZWRb9XuoQLYdX+HTDPKlhEnyxMWNlrQqaWv+YfhQmHTJtFJWl9ZyXWYiK8h
Zif86GL2LQ17ei0qPM1BBbURbBAu3gQK9ZUMQV3Sv93Mi5b/AzY9wPYrxOCor0vz
JRB502NVawco4Svpxlk6ro1zCN068N0tRy8m72ut9K8EG8wflqKKGyx4TuhUO5qt
X+7hvmmeXue7T8bZT7UlSyzMRw6dsqTTpT1tawj4BvyxWSyhEe0WXiLp3R05r8SJ
5VyvWuEaGZNcM6nUKpVqyvHCGp4uD3sreCbSt5O53Du4b8GEx2UUS04bV416soPN
FY72GuGeVq0kwZ2jdvbl5/z4cJh9n2HnvUc/PTxOFdDsZIF63/ZN6Oeb0YBfDFpZ
BmPOtqP5I1sD8OgCIgSQT6lI4I+lF2uo+UIRBp9VnGLQC3ep1BVO8/bGYimgsEzC
WwYRrkeN3SlAt9sUUcMQpbi8hqgBMkPQPQGuJqparS4I5ucsBtaOomwsgh4J9eQy
E8+dip+Hw6t8b4coxVaa/Y5SVtmuNfJgQCs6dOrqWlLW7aJT2aSrg7mHt4uUcUWB
0tMp4LCLxHuWGMZJ8CRkEzR+0KrMuqU22nTypuumx/E1tmB8XRL8x52ga1tQXgBx
F0S0i+ti1BSQ81KSRNh+DNBjg5K10sFZCaCss5P+rGnj515r5XTLyLLoP4jfM7Kl
baiRWlvbTwek+oZQ6uA04JDd+LZUpzdXrty33iiBQaPF+F79fRKSTF7mlpFD83FU
DJDLkBjperseUbcJvdrJUMl1S/HQDZaBboM/eD4VjhItwcmdyBwRo3CfnvTV4BES
izFwdZ2WwJYap9cM8f65aHrFDKVUlTUq0ojRtmuMSoXaIluBqiUf2zW15wljYIBH
5ROULSkPdOGCBMD9wObKL9Z1Fv2ZKeZ090YXhSfKoShwRklL12lLw9pYwe0WlbyF
IMMOngyR15/87p+CCq2COPXZ6RN8H9tv5kPbhTfxKqyk57y4ntYr2kK+9eBVLYIQ
1ti0et9GSoficxp3MoX04fQINFwA2GaI7zXvNHHU812TN/1OBV74W4vT45YCdY4x
c6nmpKuiT8IYb4HobPbfkP604qBNAkwXg1NiQGNoMNW36F2bn1d/VplKTjEG+9un
z6lhaTKc1b/ePWpOfQ8vCy5PZCc+v+NsBmE4xhjilSYGYiy9R7yH3RQgmgbPz0Zk
jVrLHZxarwFwhxHFAIhN8YxUZbcFgtjwGnMmiF1Mt/l5rgjdPqoMX5qKUd9BIJpD
bMOlfSrS94fl/4rL3RYr9sqoUD+AWdvKkN3B+whgkxPWRciyrbHeEq4s13AvXpEB
09EguUYy+ux1YnhCoWWpGofiD9l7TkyKoEbth1RKO2WIjkpaJGJYaBY5I2LT07xj
kxvVKCI/DNiC0Cu5XfYGFWY+5O9jiQEkJ+lZDO7O/R6duzL7hu5IFFb1ss/60ymr
/VuR7bJUQDmwMS6/5N65o5YUH29BlLqsmgSixdllQh/bU7QXIL8UTOECQNE4B1Rm
ziP6MzdRWONNxgt41jUwwhXp7a7wAwNxQA/8M42Dl0E//0MupMSkjwJYLJX4zylT
1rLyGQ86GygVfdGY9XFQGBJCZlilPTElsEgi8dcQoIjGDl+UcV2sYxAL9ZplPYb4
oilvwt8bZNMsQxOsuZtqQP4V3fhjuguqkbyvWdWSY8BdDhlnvyvtee0gDMDuHkze
rufBMYt0q21yD9vX7RD8ImOAheO1oqHZkLDF4prHUe3YaOz5Z4uzbMmcXukxlOcu
2i4GayholYNKJuThh+/TanGMdYFxVODaab4hYYe9rdxRzRAylXl4bSL/SZya44ox
9fxxGdF6Q+Y5+LVpsovTmOM7gFcpvaMO+XKPFOXQfWIPeicF9zrv5eTR6SH/K2z8
9ktwLDWEbl20lCeaUL00Z+DC2ylbvOiSHj4u0DmduCMYXBHPPt0eipu4DFiR4j5Y
zGwFnrHq/Klnh+xKTePUZjkzitzS3pRMloTSQYQt0mkRAP1a67GOY41NiRTfpaEF
lzAQgBZ+BzLM9oxc7rz25Ga7m3KxHygo86lLtMbcMPBJd5QnwR+VYoOxsjgEOen/
ETKmpqn9m3HB5uAc6FNvPNYOrGGfd6vU+n6xC8ApluEo1LGMpxJrnmoKEA/Tn2DQ
voj5dRPWmRXGkX/eEb+6qhXG6SDa6linc2+UTygsz6Hq93T5Yqsi3Z9ak6HXu3YS
89TgeIC6BlZqS3yWKj8Iscf5a3PlFsTfThuoApCF5pRZCjnEuzNvOZfaLrlOrvQy
9uGYrUn9dCuJVBwlLrqJLu0Gfe7uOV9OQyyJJyl00UVHSX0zgp4H0xLQgSP3f9rM
faq4eGLQKIKiXjkXCXC+ygW8wJQzaghQMwFdWpBbVnJRTmXT3IqmegBTYaWTbXRr
ToN+WfCBwdjDExpH1wHVTeJfFKLhfbrmxHRG7/xLO96Ly5OBpiW+FCUNTOuKydjy
F98OwmClcfE5cfHgsdTGz2wq4ub/PWU1ZnvMNnyvBCNN+PusA4QCWumoE8wVuLBT
n6VwK3pWXw5lPkVzHrX96CxVB+B0tfsBqiJfAjBpUgMGb/XOEVX/FcOdA5t3CRKk
1RAeBu60hMmI7Z1ZWB3lr2SDefmM66hS1AYSSnfZNU+U1gBam5Pf9ToMSpddCbiS
P4gr7LlWCcEvKmZh1aMm6mTPdoSSqvKFgU4pR8Msw+ObV0BOusvkf+mPEhmfk8HS
54CMERO82hZj+DXjC9iPZn8T14Y4HLC583WYrBG0k/3OiXBrEM2IVTcInkxkDmiQ
ABCNq6HLaWdWZWIuyc1tSWsM+eBHe6M7l/GA7jbwNvt1MkZrvd3KT5pYo+DyOk/n
VV+xxuEGM7EjaFI1aKK7Kx2CFkLiVkDYqH/DVCFVz2ZQevCDmxC6a5flOMn9Iups
NPWEoS0NZzMSfYUIqxrE0wyS2Nep1UJ48Z2LHlMFZqMp+8jk397GSt8POjthTC7f
4u9ikVIhKjmmJA5eN2pnfiQXNVH7kUo2AHapwUxS8jlkCDBfhRV143xl3JvWj7FQ
ugjkCXCNeRH1VU2YUApKm1LsOQsg1mL9wCEl67K3gyb9/d8NlaqASC0Bjc74VyRD
OPDmhklcUWj0LmGGZNRQe9uyDSAhG4rmqjk0U0LSOOG/ZgGD+MjjSoUFZ9e4Unu8
TUx4sRzI6mMMrnNq9Urc+lXJhvzIOs+X+pL65jCoA90YaJGoTzvrEULpxaVOPGVn
THQR+9LlqMncv+jepdeDMBG6u+z01IyKMUw8A/yEt2rAAVJ8eNe47szUsAa98POg
cX2vxHhoVNxTy8QBOErJa9zJDrdodW+ElA74yKYxb+qdY04jLOsP45u1BT8xP1xN
zhmE91Cu9cAR4GHBmx9amiL6uC+hNWNIex8sLkueqzt2zicsqGP4IpF+AYOawFPy
jb0Qs5joManQZgno8CgGqsO7uPkTiJPfXfoKjcMDPDIB6KnoM65lqOOGZgSAYUtI
ocJjKUNodbTwgucEIEBJ6DrdGUNReaXhDj6VEDfcT//M/wrg/o8l53S7ZU0/vhaH
DXsBvc7K3GM2cutiugR3yowE5rBu8Ww/ClVYu6K1LIF4682DATqv/K1iduS4QMkb
nytHXKI62GVh/WFpfzG3KCkbx8babO/NYGri3CkfVjUnvfU3MbdLp+9vhxK6XN4z
EbtV+rwdctUaEa6AaGjqamJRjt0Fq1LgTtmUeIvkYHFukxWdrUUWHIsJXkWVrrTK
ol623WQmh6xzyr02/csPwuTepsXBTS+jJAnqr5V6l1xFUlS55mgq3GxIxyGowIh8
yd54fUvuQcrUA9RFWleEgrPPhF6k8S6ch8s7U0EcBW3Tee+GBDdTwHdB+e2n9QrV
CGgDCCLE7iTgd7QdfX1ajDMddVkVlwIf72W2NmK2g/jEwwCp/VJvGVQa3AKzSfjL
F9l0WdoEngD/SfKUtlkW6GN8o9eJNki2qVkvwNkRK0p73tksWxeA9Iy4KiqYPBD+
YGYj5/4VKgkXUkbEVPTdKih8nwfqM/1HCmpyTszavmtp5VNvFVisOdvqIlh4scJ9
+OoWDNud++yv6sL9G/tgynhU7pgdWL7LzNpWSspD5rKk/VtWeKg1bsPRjIZNrysc
hnhvi7+G41vEO3CNHC8JiC2yLnwurIT8NDbyomc7nPeZKzOuj4p78zE+H4dM+eaJ
UFT/ExergSeXDETwMSv+ifDY1OiBy5K4jWKNxC6ogw12pbm8vjR4BQFx0LW+vzZb
OpGvA47PXyTE2RXzkLp2GQ9TKkSaZq8W+cTTt683IUqTfVoJeYrIU3lJiezrBlPy
6Xwc2Wa4FJRSh6fh0yOPBAJ1bP2JgSaaDDxdo7muUhDbwh1i0z639FiVuZAjzCWY
NPW0c4quePVluzow/avGB70U2X+m8X0/nM2UswKdERaOkEOSERW94sNmtPe6RpI5
0bmg0nMo6KUdFsdp7cie+f4RQc2atn3Cv9bEMwukPYMsI0BoEa1edPzOBwpk016r
Ypp8bJha+F/uYxk0lgOm03AlXRv175yT1yy6daWjjo143R/RlljQXR6gbO9Pbj3g
7CNP+XDPSOV2CcH7XVfcaJnmOYFKGCX2HCkS/7ICXXHz74pQv9xqmxDmLX96AxRj
LRU5hYYRlwXHlyCVOi0PflCFfLWQytw6aNqm3V/jL9i4khZr50SVoCidn1BDiEhV
WdOURx+R6RfNoBqDMafgHvbvdJnaB0xQ00eHEOe/XjmpDdb0JpHhDohX6fUuOi3v
7Q3iKICrJAVw/MEQ8liUtjh7aOrIlEx126/T0r5DkuvzWT196k3mWtOlE9+4O8lO
3OrCRxq4cozL9pLyBY62QMN5F8FRM9zUjIazzlnJQMZWYJ74QXXGWxxqfIFFTyqj
UoEied0WB+pIPwauKfvEJbQ6yVtDUxGtohJvZ+RBB3tg9ftTNuQrFsBU/r2QZVEj
A0Mtf+zJ6Kwnw5MJYvh7/8sWVxjzLT8Az9QmlgvFpoRsmFQFU/TpBf84vH79oAry
Ed2sDexPyNCxcrNjWgBLuw80b7XRvEjbnYHbikzxOKO8FRCfDS0RFUAivWfaImuY
czgSrrlcbEVH6SP5YAV9X0TfowuZW1+Tqw/fVb8YJHwiP2nw822trv8Hm0zhdgil
SMmiJthb7+ANFEnLfsgJMszLDYTdUMReJWCHQ2pqCTMkir4m+hW5WDo2lWic6KO7
xdkYsN1hnaYQVbEn5tGlPtcLCBmOfMZpqdFSgRIP9DwFFIM/asT4NJTthcOieau3
3sWNdIAaj1EgoEYd4t+ZGF7akHVVSH35quwxH+ntzqEKjdHiq/qQngQj0O9Jc2Ik
ip4s0y3i5ltmHnRIR4+cOqVO9N03znx8dx7/CzTKLbWxzo8jBF1pUND2vfCeOVkM
/zd87aI0Qg1X9uu06TW6Vg0dmYLOiJENZERE0N1vJpdf+/lNhrHkK88Uee/JxCAl
c3PrD6nyVntQ5FH9h3yzCT453ETe5o07cu0k4G3dj9hH5HDYnbG58kjULEkmLq0b
FzclPAi0CzEjIFqOtbIcNryq69zG8yGIstPFTjvnAKnZKaMi9IWAKUmPN4qUrGt0
iR88Hg+kU4soyXMNmgPgyC2d9ZEkmWGWEGpjjaAZyKITZ2z6N33XIDoNQ7MuWK6/
lLvo54EToCi6piH6RH5vc+GCC3phfMQd9u91yBGuBroXQgXgEwRr9ZPdaAyY4KnU
vVcSqFQ3PYHI8JOg47Cm2AfacmDP45qA5ZWdhvw0Uk3+5EhMWi/Xbcihl/AgT1rx
wkInrb62O1OwFLlmiGXBpb9sWI3riNo4yasCkg5VJL9Hh4czIFM5TL9nEwfLCU0I
28IVaXp7L/Pjer5RH40jbeQclZWijNWNOV83+K0Z7HL0SPNDnqcZ1ZCJN3yV3wS7
ccmzMxr5BzoR0ucRE5F6H61MVd8PQ7azdNgaxA4bHT3zQ2lw0KFKj09SFpM781WR
aUp3xozBH5B6nwFs2ASo5l4t2da+QeIGdY1ZiQYE8mhfOFELlvadR7X9XtyqSLMH
v7r3MrvtFR0ko+4aTksQxci9z+QaOVgPvgy1Df+/xl1jrhKYg+dlmIe13kx+OGGd
6obuRsi1OiwdGTr9oFWBZrYggab0i5KcLOhVvcwExWR/czX8vbS440WGy9bZq/lN
Fr5JwZwECH1G9v06X99/9rCXfD2sQmJL4BuBEqA8MmhCeX//EXrHFuZHv34Zf/ES
mCyJ6yS1BWzOPlQ9aYeD9ziXP+WYrVNXIfIIeTQj1lqPb5oGqLFePPnowQ/T8hTy
KeijMM3UcUvvcpUhuD29joEtVqbtOIUDSSagi+1Cm+BjwpxFuoDSW1mRZxAid0SL
Wn9g+rg7WYxgTdsn0K812WqpsSt697WsnEjFRpyiKJf1lGPBTFMGn/401BjSv2zi
GB+hp+P3PtLAgUERLg7pyB6e6eK4KkMLjVC561SRIZw5tbrNyz959LsCuH0ZTrLF
2hrpRdxYjUXkDiWTElctYuQTafBZdTvE5G39l8IuRtSkhCkUKd1htPC5+0ofK9e7
mighoKn9yGzkRxgjyPz8NjpvjYoy0ntiSS+OZDJ8FI+NOmsL6fJURobcpMnt+3kB
HNS66vTVLpN9BK3SjN0gRxLGByxIMTZLIE839yK2aLM2U/LU3Dq1gGLHWE9iCtit
PP6de7J7MhwZA0iLBjm55+eEci3wPTh/eE9l5+Kqd0dbHA00CejzmPZx33hkVsuA
lxdOpA3d4Yc8U2vwhSRVQaeVNooH9Gak+LbfPV/Wk8sWJjLS1kaXvgWxL3GQnHO1
uJRBHJ0G26ysIVPz4chXibKv8Y61Js5ogLWJAsY/FkMbi+6903ypXtcxNtFwovxl
s2LVWpeRer2a1miWkWfRobP80P94qJCRQuN57zMHLw0Ca1RrjU7GDvcrjrnPH+zz
FAKhzEpKjVRrwa2h0hY4ZYa7GujeUufqBohaPBtvZDbxS8imUSN/DigVSAgECFYQ
yYMO/rRX5f1cXkk+RnEtPnfJrN9jJfJg8RZ59zh7Rqs7jcjcp1vJBJWxM2J9Ov35
6Pn9U46L/YenhcJZmVCLAvatRR0dbxrMfdWe64KjMBiwR9cU6pSiubxC3w0nCcVN
gtWR38k6kc1atMOpFanHMg7gLXgvTj8RUCezA47Y+xFM26q6NkyJhcunyE2UqumW
9SMFzrGxuw08cvR+HkzXmxgXwbAWJftM2s1i7LQbId4VaMQpvMbXRk0CCPY8yeRH
b+wLMCy8FL0s7dQaVlqlTYjrNmHj9Z36oXfQkEA/yteYXg5pQf2/nimPz1osz7dH
et9zrZo1HPK5cZ72/qs26T9Kyk8edDdi7qnBKc5ZZn2P3Wv2FgPEl66fvoxl6sX7
XN4WQGv+nGsM0f2mJcUi66TfLRVjvpWngpyqMEhmhz37CUYj41PN8VOnyPxz2f6N
aFm46r2yDdAzj4ZXqTj3aa+H04ZqN8dDpzP9rtK+BFk2QoCwLy3Yec1qzujPI3Ni
OeeTyhTuSg6SF0QAphDFJo9YUl0yqoCR3H+WbhWsMoJHkk6a6/6IJv/FoVgl4QC3
TmaFNJrTNzCIrFhEbgvZwKhm0CGAKmlnUt4D/sz+k7bk47vlCvchPEbBXNnlc74K
ud2AsCg5G87AzhVIq9SiV3Jj1VHQBZ7QhoFDQmyS63zXxGA9pdCqsqAefRl/A1u3
NmsoXhlDImcwQ+ZgMUk4VMBGtQMd8QND14Nitqb+zj0uLbDSMlWRjn5QnvzygYZM
fNV2VarOY/9V06LvA2fQ1B1Rf0PEoEzDUCTTetSuAFhGmOa1QNPTWbng+iu1Uh7M
KHZmA468M13kBnOF81unSZbX+CJVZHfQmSFCRVa4hCLjNsgUxVnh0k08TVyiwnJN
UcxHmK9DWIINxBiZTmE+SDoi0oa+kz5AGNaoWwxDaHftDuOqJ9sATNEypa/ZFCw8
JNilpJX9jicrRBMqxyV9JJ7XJESyul1kzi64UmU9RQ6acJ4ijHr7au0w4R4Yh9e7
zO3WXHc/PvyUIKn/iDdZWbrGdkP+Mp7W5T/4kUyexDm6TSEm04nsJwKr6LAY45Pe
GW6SUYhPOfvrLX5uODzrs3cxpDlqWf7dRTwrEhPxUg8K3By//J7HNhpsqToqUAho
6nA+qDwXyby6w6RftK7KEb6n7M/it4kiyL5tnvBxS470KehoVM2YgiM6AdQBMzDM
DBb1THDYWajj4LOU16VcjbfoRIJ6JcICH5dijz7HXsRmjttcyioC3OehHsyOh5ZD
nhGdQc1IgCe083E1vl1vC5I2ETVEklXdhWSaRiyyS5jr9uKbPNKiA7wpiJ+/PT5v
TsjhiPFf4EpHlTzk3W4nlPj2SFt0AJnW0ZeBNoda+xFTpy8MyQdeWAak2w5gaDlc
w9F2JPH57QUFIytU5UeDQiKm43qyBHCRKerUa5O+7HmsAjddSkJExKZMXsnGDFHj
IH4+NP5TZhb7Q+UQkXB3T5ho94ac6yIr9dc0L3/SHoP8oxJ4Lmm8X2J23mo4GX8W
FL6MtRQvoqztUjeogUgAtJJZaEL00cTg3DUTZqTQDGx6Veazz2DgSPb3PZ2CshTv
M5NPGqk6aNj+Ok9E2heYDEeIs7B5TJjzsTPf3TpMp4nMP/w8Wm3QpssQh2LBgHpS
d/zh2uoiUy5veGEcQEL6U0eowazkmks1FQdLxQIkSaM2E2W/WLup/EtlYCcFbHjs
AVsJcCtIWOMo1XjVwvsmIZbbUeSVtqrtbkp7KTD6WGaByqhxTeQ7cjeQ5Qr3Kvi1
ffd0N+z9CGe8Z6Z+p59epCh4/BTKDRoKi0YFvsKilCaGwpUUYu3B2lxJl+knrNAA
kQIZ+nMZdLBom8CkdKP98X37SmvkmbwYCXXlt9adfmZ0snOxGT5T13/L5pyAwJFe
ne/pgDdt6DN0O/io5n0Y4Q8PfpAHaov9g96Izr6DYTWEbc6np+aPdjcWrvu+FI03
EWPYXwtu1SD2Xw77rmdQDUw5T0CZDBauFUu8y9ZyHeGW/3LUzKcWA28vfFWUsBN8
WGmPzzPgnu2Tbm06aFUy4uylfG75Sb7Ql609C7iWfmv8M4AxKW19PFEhneCsFy2J
6O2jv6Vabr9HuPrEMXH4XsXwbe7eECj/pxE3bDegHsx3gHmvAc/1HNYDeqjOLgDl
birsg++7L8IL67kgaNRzek+yUKm0NIEZFXuNDQQRkaCP2ko3ztvQoACn+AY28PDZ
IrYN9rKMkc479s58gxk0HY7ha5NpQErL2FHc4uYwxfygcekx//hIvnHYMQyS3ui1
YniVXpeXv/J8GJxq3/75VwFfR/YhPwsopftYkC34vdLwOXLVK0Uv88WlgU9TStJN
3ealnJAJquYcgBvo1tA8bpO+1Xzk452yWaSj4qXruUpZqPjCNT6NYRoloFuCuAqu
gElZgf/Z7U3rHfP6qhNHo4dzuZ4Gx8wYGWW0RwXyaOwJS0IB6CJSHo5LyEZL7x5R
7ozpRjeART5a58N50rdVfz8UY2WhmbAD0G+EkmK64NtYxXDf3x9y7rO5l9ZehnKG
UeLLqJhX5zAS3AbAABY7GY8MzMjO3gkjAVX+uJdWa4bRsBidVMgHH5vH0LKHd+6r
lwBtuOEWYGvf90XGKYZGbU5ogszMiWJrMRMfiwJBBtxwuJEuVLRFLuXCPaZk5Bs3
DNokY1+5Y9DBvvVqY83MBGgNhKS7Wyru9KZel7954ezAmqfxFVnOPX4EkixDGvXB
m7GBMziE/vjSPv9Tit+6XOlsDF3Fl6tQXu07ZDs+eKX03KchsvtE4eCb8DQKQBXp
ttFAwcXJecK86GzrMLDA+isz8B1yvkMkYZ4TgM4gwG+lvJ1h2rzdvvqGCa8ETdzx
MD6xFGEP9ae/smmkNT2GxxcGOeGuW+8ZsoKliO43ZbRpSHvY0ld9/TAgT24PgAXY
ob6S/t0RystqCPbLt28ff397whGXe/yqP7A9dZq6etqE8hEMj6kpBuOMw5ePaSuM
9X67s0U8puUhgvFS57w7Fh+Ts3XdziFyG9MgjOTo2lrBjkqa2qCo0zOzOScgNPgz
AsmqqmelExwchADfrDqR6gUdTxZS1BAc6QWo3Kn6PSElqwCzbFJ26ipg4SqB1em2
QgN+96fZNz28yQeJ2KuocggAlSEQDheWotWuVpOfvZHYyIWnRj0AQYK0G8dzphZQ
Vir3JFHiC43jSes/opMcV1rmsa4B1HnsA8zyBBJYcpNC3emJCCpaNxkIM8JFHwDs
uA5CYlk0dcGkXimFVjVn2JD63u2bbo4WKBlqaH8ybv2+LuVXlJ9/NL90r4LKVGbN
U4cF2o3nMmlPIroaIsY02EOIgMT/8jN2HPGe6oboJISHNJIeAgQ2+S7bWSvgWTbD
4IF3w7DVcy7BiWAdbBKyRwkg/LZl3sb8V05egRgWwHTpWs9M9N0ot++9ObdHn1FA
NVP2u6xPTd1mP2aHCUZLjCXCZi0SQ3DDOiduABNlKZwfFc0hPkxA0gItaiQ0rz4L
Z6Lt+AYW5CBesII5vIZ80bcGCjMya+oaZjsVZJuNU56QZCYqO2dXFXKJZtlvOobU
ZDPZhwuxZiHkq1Qfm6ybiXbC81i6s6TgttkXFAaJLH5ZuMqX9yd9ILWcsyvoqzko
SV+P8RPIPD+WqvLIN05dgfeqGgPpwdiY7Hi2bycyJ99A6QY+V3GMbKUDi0i5foD/
PfsUK+x9PFuthdD5pLn0CRSdv23NQQhamViJo1hHnR2n5Ji1tDSUm5+dcKX7b3wo
0bBX7ayOSxdYkZs5cVZGukN5ms7Xt02+9+Z9mvO6mvBoqVGRFyAI3a4IHxFY1v31
Fl2qBjqAk4sFD6AmKXY4CKr8j3OgrPJVyq4HEH9r/hdRWB3osh09fce1IRkCmcxV
1bJftqOAK3wGnUsxLb0fOsB2Jm0wGhKNkwxPoBq1J7Sf6ikFbsqrUOQVE9TlbyZD
SK0r3ICn0lmd6+0iaqxulvqNIIBoF/RkypMQmQhrHi4wf1masSaMeIpD9aX0Gq7G
U/ZsI8psbFCZD6TfuFt1NJG1MsYdA1Y2bjAwC/9kooXJMgzRhAwSw1hGOiDhmsmQ
+AOsWpDT9Gt68tgahIW52ur+fYUkqFIVgnBdnYI03I2Ll16/9cvFEORd6VZWL/8H
I5M4cyAazT54x+My/BcGdS/cDyFCpQwlJ3mHc/QBF++3S43BZvztwdI/MQNvJu3N
oQgxv0L+Sd3S1Y+QGLRXiS1ks2W1SorLM3lo0Y0PAcp1mBBiT+n5yMEVpwFGHHc6
Zar+5dmWzv1y9Y8tCzbqXud54pr7lDdi8ZpR1BjSPlJHJPqgx0T8W8Ik6vVRBmKp
qI6IYBCNufo2ETsUq9QDEWNhVYBCRERqKTwzhVSEbjaTBkIEi28AXqW5Ty/z2kv6
hjk/LlPFU7aKrdvnGN/xoqzUEGVXBf/ilASFrJXazOwfhEHOQ3tuBrBIo07juBRz
SBw+GzYQv4B04DsAE+VdoJKRL4r0FrcOuSb5uHJekJKYNsmMP5U8hy7fKnfkcCG+
Ihgxu10JBpZt2jl1wsLeG4yoyQSlZQURLsnp+wmrflmF3+zwadqSK14Zxk3mdbCg
GBeysEoy2aMNL6NcdemdHj9pjGx19unOfU/ep2kMoWSZvR5yd0g4lh44TsPrrOrw
sHjVQd7A2Wv7baGE2BPdc/3IeGxYC1Ys/1+4HQtJTK97a+pxxPcWOukmqLJD9jlk
PheNtTZCgHa6h7UoKKBDvizKOtNaSklxFbExxHz5x8wGfs4XDz89Wf6PTn6HTI6c
7lqClsAEH6IZv+efMCckb79W7t1zdej7f4krzrcZ0cQSNjDET3ChYj1mRKcPEPsX
flGHyjA8dwZ9iW4hH+P2q0YQSlXyRJerm60ycTQRQGlTJwk+V7JgIoxF96ZZOwwy
uOpQuXnA3xBQi25UnTYqf90GRH7Lji2x6foPELw3YyNR8p99uhkmbx33jr208bvo
yjU8/qzPpwWnHBYzuvmPgvJZdRjrxKVTN/1o2YeLaPFX4mO4H8CaGNMTAUhEQtSU
yJGakXmdX+QySEpTWMNgA0GAP1/f18wO60Id7kiloZBWIloprEQ9u6lX4pmLJnvM
XPwRMu0zUe9UFQyuHp5VJjTd+sEcJ7mebCVhsr/WjnOGCa3FcG5bFElNtid83FFA
9P5+5pMqjd0qqtUMqoPKey7qaJ3U24Nf15sr70foThyYKsRBjCgAb6p/tzJ7taPz
syEU0uZm9Dm6xws3RheKG/FvBjo/2ogFSpCwjWffEuRzqq04ZmCQmECP4McJW03n
544PAKIvEFXSgNTVEqd4vJuWBD6ToKSAW0aGKyuUG8zgzHZXSggJHdwE+OGueDKc
CyBnuicZ8Fv+ySK9RqMwcJ9J5Gncb/XtSUchm+whewVRqCSzdI9rrknyqXAwSIGC
vkKaxg4wKWcCOhes+CH1wwNEYE4/lt1W92tqf/k+pgduqZy/M5ta+MawGQUhJCBZ
pc6LG39paoflv8riAolPLb6Cjh1aq5tCpHdHqIkmxtH5eKEhlco/goIHkC/SO+gT
h5xWkxB2+8lyBX8ho7LtH9HPGXJ3ROOdVfgpDCrPszwLKgCYUcJ3ofAaU466WxnD
Srojj4bA6ZB9A0l2vDJ7xcKje12nNXt/+IFSEY/++YQv7+qP/0H6y44NHPldVAiJ
brJ6SpQJRZgJMYUh9jaT/sIqaK4Wk4jmsWA5J0ph/DdSFXOMfYRZNL1hmDrlofkn
eU4a+pLUWbpj7QF0dXvDS2SLxbZuBBXBGrJt0rbSDWYNtSrJXCpG/L6/6g4qAYTv
+18EPkyUj8J39zNPH8ZOSMsKQXHvXzIqpOx40J3LFJh9WiXfS01wt2gg36AlaQLT
J1kTOAkCFgaj2gaTG5Z78o6MyKCtWNiMAyEeNKmfsOzb/zZX4oA/2H4iTfTy2ZQV
FtEeCGww8oE79T7NDhmVtlvnJH9Wnq7fDA5sO1SDOmvXM2cLoGU1cznpQxD8MYRN
XxeCwv6m/Xc1nhSoE5oTaylEtARc8c+yFAtCwbNbJzbAvcK0cWmDZNMvJlPsP5KM
t5xj5js2p3Btz4Y4A1AesBI/Ab+7MEcRj0psit98O+UIqesKA2poWa1ZmnOCi8BV
EDLrkmdkUW1h0cTL3AqSHSImJq01tXTGfyXeZS6uH341wYbuZsaF74c2KQEuVjgZ
LCHaeQQ3yCSxRuagwOFwCzfdR7UP6MdRTwm3b1C/8jKu2hb6aSZ7LhvBh065Z/eg
GXPRHpCvprFr+qCMh+i1iRnuXRPmaHJR78Fy6nqCbY0i9MYMvWdm8AJquYSwDmU2
cM9Yp9Mi/c1BGGmSVEtwmnsFKkP8b6Ih9cjFN/rK46MrvoOnglrvAKB0xk/MYHlZ
aOQ9jbsJnbZHPabZUijf9EIpHINLJ3QFtmrLjJ5iu4BIgrs5bhTK08p+JsPAWzFt
LyYm2VhU6WU4YtAkXiiJvxMgAGuaq8HwcKklA5wPIljPhsj8YZz9JbxnJAvYzQx9
sDoqNOIjDuEbhfmRvLcZSBcIF3aeOUB1BakOBuqKZZmNvBcdsVgZmN889VcnxRI1
JJ8nJeqNpPpa8bExGwoOR5iCV4+/LeklPhSpw6D5ceamuSVcl9NcoNKjqWrGL9kC
NsxCzER7vkw5DjIUrw93yWTopWLKZ7s1ksPxYqspnoPuxjiMHgYWuBSvHhrhBwy6
QwU4toMwM+Y1DVcMLjvNop7gtXskVhtK0bi5NQGebC3O6rdWUHlmvRzwDDg7zwEG
I5pXmEmR9q5ANhhPRZsjLpsHEyOCaJk9Oe7Y9fYWhPnHP55hW6iY9vN0014NRFEV
1ulclZQmzh70Dds9VTxIwN36Ph8Yiq7qDmywoqTpzhxLniPDmSGK/YSh0RV3FiI/
EIjkomRM5vyERAx19fPwqE+dcA4OSniz5rNKlyw2zxmwjBCQvdlJz2xBmSnIR6PV
Lo1SPb0RnTIG8NA9E3N0dQ21Y9nxm+8mdbJSMQB5khx1uJjQ4/nq8cVVVNbZ/COq
nd+IzB8rVnDsIdXrxaXeff+b/+I0pCu+YO+25ep0no3AgawAJRPSuaNge/fMsTX/
t6WRLrlDNXKQyHZ5M+QUNlCE+ieq4qW38vs572sv2m+GQoiasgAYzmduAaRvAPBx
DeQA/eIo5bKfl+kkH+y2tjWbQmRSFu7uL2GJhBam5k6ygzTOG90jwR9TWOC4IVaG
P5dRdr8qCO5/ylxkxu8HW/5Es+pgCT1Js3sj60y/0p+HFagY/jzOfhBkaL04zc91
/FwG533xcqBvDfdnfTGTj5Wv8dYJJipaZ1euyYKkdhd0Uw+BrKseWpfRisHynAL5
5lXwsvmtxUQ/2lEldIn1uB6RQ/cLISDsBY9JyYk0rOD5GgWtAA4HKVdiljNVKOKr
Vc24US9Tky52ILpCY5bMMcGV38FvHZuzZkSiMHxQk4JfX37U2sKm/VfSHf8Quk0O
rtpyblovQmSx8RYYXqqA+zkFIroGoV1OhgoV1yXhy4AHMaqzZuea2Dy6J+Oq3hB9
yAfvz1xuMkchZ6CoFdH0UnY8Bbvj82mqaUpeaM+2Ip+evadAapBgFFpHYp0sH+En
+4og4D2sFsRIaN4QfA5JSUS7MyFZG0h+WO34LL7tHkEyKuPEmjdHNx3X5H5vi1rN
mvNDLRsaxSukXOEN2x7k12fC87HDZY+bBG3CCOS5HB2+LO5mwqU7WdJqdszwMh47
xC7kE0pebChMv7YU0shVYM3eDLDi0oUQ0+QHSsZa4+rkIPjleRpIgQROGxpkwTKw
qwXv2znB0dyZ31pSF3fHimk/2umx6YWBq6CsfH2aacf3xIELFjQ6Y2Ycj4zHX9hk
G7IC9mOt4BUbnsIq28mYVwJMq3m70uHadZ1aJfwJxVlmoz+VJHnptsd/CtLtchau
M3qg3sAzXqDyKe+8VMfnpODDfcchdHSUWuFOMLBcZoccojho4e5W5SfhpInRwpsv
ZR3dODiUN6kG/lFBCRRRvjLuRec+/WwM42f3JvmiDVoPCgSrzTdGJXYTZ8xZqqVa
xXSneyuTsyvBdmCirgIFSNikWbjfBg7SNlHE9oTXy+755F1whsVWsngKpZITmKNF
FYX4pHJ3SR4XNyDOw5rXMVFEyeDjQ87cpgnjeUzkOkZNQ/IlRJJHNUJ1BOvfWRwA
I/XuSZpUcFYs+G3D0pLXi91zOPXmgsT1NRna9aOTfimIxFAYnyM8HEaoCke40L5T
3kDJo3COvAI7Leo2lorVlumBTLpaiXIPQS8GDL2A0qbFeuMpMIc0D6IeyFcHXBeU
mUUGDqdDUmQJWQtSNd9HbX0eW1fs26CqOHn0OUJRi9XtM4wmw9CXJyhN3/MN2d5D
r+OQzM8MDzRf8CAK3RviQxn5xifmWj7zKjHUu/SMk9RO2DPjSPiqdLNlvI2j0ivO
C7B0gwvqKK2I017eXtvyTq+RfcSMz5dO+AwiOKO03J/sdLGR7PFuvG5LYKaMlxol
9dp+6/5gX62YjX0aXUkiKRzyXqId/cCNyiSbBxjJT6lg1ElcEUSEGduFdz6x2yLY
gwpS7gPN40CVuGOhC+EB7yg9JPN0qb2Z/wxa5vqLwBb9RG9sB7EXZsuwqp8NwVAk
Q0NQkVfKWz2oUicayncGxlILYO+14TBFL79iE8LRm9WbMQZFPJGohPfBtk0734Xz
MX6UozVgwt+oU04Tz0ZX3EX9emoiIQaub/N5+MpiXI1sojlMQpW18NZGgq48W2yh
cwRdYAFuTO7HEw0iGm3ea9j4E/as6ZDc3WU1B4y1fUQr+r3688Tk7TQ6eH8qUk4v
HycaYZ5s5D33QAJSrFlQe7Zld74oJUZP5FXsPJcULmBZHo/WFBKuaHni1CgSTAFU
twfGZRCd7H5gCkzh+6GetCWp4yVDYrgiDHQ6oOvqf3aB6S8fQwDAWFHDGexxocBi
Gw1V+TIMGRpllR2s1crnyNoS/k4FIbvrQOPG9S3Oq87BqyUwbPOsFvhJHGaKU7BH
7bFIL7/ig7E0G18tbcaCf1aGYAqSRfx25HWMoF2//JOTUgGf+WSAnfLWl96dK2lD
CCT5qANHzQxaA34ezd6hAjyauqRzmkxFEMvs6P0SZQMG+Jstz2AszW332+CJcC8s
YkCYhpxmLUK2gyesOb/Pe4brwrtM2NxIY5vq/A5k1lh75thW/raRWFAOGfxBXiFV
QSjORmHDY/z7h9zZa6P867Y95eiIJCU+R1M7FBl4PW8G1GJ/s/W4ZBj9OPfH+n2V
Z8FPxHRlf9IFjqD0xUkOBB842UBPz5gzO++r/lKKqG6Yi2gKXBRgXzNBE3EA25Ck
TI3I0WPuywVMhrWqbNcWoBZas9rrmTQV9AJbek0X1AK9Ue08SdGgam+2ez/JVJYd
gIaDUZvOMGK04UMgCD8cy67Nnt6NauMUhT1TCdSrU1AE96Y/cfrU75+ICifNiGqH
`pragma protect end_protected
