// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:31:30 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
i3Prw7dylPCWsYJOaZHg2iaQyi+BXUOHCGF2naHYUvHffVjv1EzfM4WFQfxbzMoT
/j8rSujxt6pAP7pAcex7MQ6jlY9NTT1LEL8nAv2N6N2mHluuPxl0nWl07poLbDMD
2qaJUMEI0sjVRuDEkz8rAN7rLjrR+AnXfHNEARhxiuw=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 61824)
ztDcDgR1EhPJqgc4wo5zCulA1n/QuCcd1LVqWiq0vW+cW9+lCWfHJj7jnhS64N3s
4CyL1lr57eHk5kUHkznHe+rdsr3UWkLxt2pvGQJBq1M0uKi21KB7hqGJJr9WP8ww
N57uNgE+3GCBKWEuJlXQoVHwi5EXE7mYGch58X2MgNjzIN7rwhZvrvUmO0MsjYVy
+Z/fikxMET83eHJqiiPI5uzsZ1nX3WwH6Wy+8PPl/Ug31kY5JxpKCNUqkR/+JaRF
+SLa52e6jrdPrxM+Ot0fpcd95mlW75El6KK1nJOydUWgloL2YjhQ5EN5fbWczPbl
BBvndl4eotek35jLLVG42o5I32ImsApsdRT2dMuQsAmTy7KKWf3VmFMDaUskZ5e1
hUN9f70LpW4kEGqPrdLAC/Uriw8Z5mrWnTPp2sJvJiVuDJ22q+odRbargYoBuqaC
MglOVAegzPXtW2lDF2et4S3K/7J43Qrpl/e/Yhv/gD+owXLHfhFypJnP+eNv9oU9
nZbwmlMfRo4BKGlVkAf+xwhemJQme4awCBUImHT67Rb3XCkH43QhsfxOVNGeuDbk
RAGcBaE0iMG0CDj8elvVU7BXywYSUscKbIDlQvaJm1STT9CIs3rnikxK7Wd1YA3K
bVfvdEqjk4sNo0S4lk7Mrk25JGSg+RH9GKSloklpGdqb9+oFogrB6RJSq9AaVSUN
uTWn9oQxhqxMc56tJHW10EArAoR8Z9t5+gfuqjaUR7VeakgZwDov9MoPjHgLT088
cey39+UtYkziKlgLzRhufoDJN0IYIYQGMxO5L5ZjkUm6o04ZK7qEeRQVInuP2AZq
zpQn/Y9MyIqnlsX4l+mBDs2ZMRu1ZVlqf2w722OfSvpziDsXLc2gWPY6QuR3B1hK
LIT3dUf0WpTGjZdd+/MkMAmYOZTCOEP9nwyUTjLMalHXDtYpR7uGCMSYvsUmRpgq
6/Uv7u/vRzvpUqIpXRYP7xXykau9++w/jrje4/HHkAWR2NG2uDfPERt+VwftduYk
cmKu/jp+VGwiENFBWmt8AZloVIbk4ue4HJ1GFKaNcuxuEEuqpXFZ4KDdFYrLX9gr
OFcDThQsyLnwjG7Ut9+HL5LGG3NsW1yOPlcDzVzVhtlBqF7ffTjJO6PPcpD00g3k
GZAtXjaD9x8Y2zsDgfVb43y6LBOfChS3z2GKJKyET5r7PNRyH07rZEOjD7X06Ps9
CQlcVl7/LUMVUiYbXBjSDIoyVJ7Guh9vzL7hPKuQFVeKqcS5L2FuyasJ/dr603sQ
iDvfj7HvQdkimPLVJQLLAM48KqHFJ3QGev/YdszkyqzVDQicsFXMPqlywU6cIOrA
MN9PQLB93agvb5CIh5+NeRtZ1Zd1J/nXmHt2yRLgzgVKyVIg8dwV0cL+E8qJcl76
DvX3RaHaoQiwfzbpko5NDwkwFmR8H40S/gGAxDSfq91UEX8csSxednb811LskR61
QgP/cX+SvPLqNAFy5+MJr2Q8ww5ARBdPEDEOT4tCJ+BeQ8IP5cIwon9RGPRgGOiX
BDB/i/mBulluZGEMwvrlyvJcod0GFIBPbx2r0STGMv0dUdsB5chS9L7pbWn3pQZM
iEmj0JzLhbZEzVrk8fFtMN8HhDimHHuDzG2L+7suxq6yU1KnoF/54aO6CfD4D1WJ
kR+q+CKIUbEotT0EHWT9OOSYgcHh14jJkDbzywdeeWYizRz1cP69G6UsxGR67xFd
PsuLf8Dnk9VaKxZcPNqL5+obSihpMm//QDgF3Uyq16dX+uWOSpXRmymLl+b2uQas
qlUrWba1f/gCKE36lVMbwqawHRoZWkC4Ip0XubIUC8jeY5Ku1mYgCEV6s1wFnHkv
hcLfIfsbtB/D4tgjSEknK4lFJZTnqbwiKLfqE03LKB02ipc9+qmP5nGA75WK7tCn
f5bm9pEsEgeq+NfYQY1/ONSKrHi1rIl3iM4Bq8DBQuEK9+SJW3QQsUx5W3YxZL5w
WpJQJEe4DUxgPwa/rS51aWc8nCTnEONFi5CRCGm1GpFUqFTiRQQK4rY4fmEnYZ+L
lwmlkD9l5BP7HrxGB6/72zoPBMDE6x8nsmfzso/PS2mUxvBId+nfsSEp3oPc13wh
clzxyryuOWDJ3c01LP7f+4umTKdHGI0fSrBK0XcnXuXUUFoYMZWmJMg1QalgE3gO
ss4FFFQw87IbsNCp5uQOaOuMzQg6MnAm/wfllOM2GJVGa+nLzz/tBX2sQ3KDGAzM
ZDdgFWLt6VHcqp7LdIdIkMasQa4CTybXheZIXcSkKe+dDRXjI9a8szt7aKo7IY+k
OECQJAPMCaBksVQC4Eb5Xa0dIkXhZ4/9fPQNWMjn3J8uI9hyAuKVk6fqoR6lvTEx
cbaqhtPe3g/dUBv/FBdFl7xCIkdB/31urv999pNfxi5WlfhPw+4jw/uW1ysCGacN
A04Y/V9fkRT6PiC0BIP1Bi4JSLAbH4j1p1GDScVYRbquk9IUWz2UoR17R+NR2jsE
1SdfM8TLVdbBmC0rl557DyXOT+O7fY9SjPeufefJ9c+dLkXRNJlZRjGY04cMdsF2
Pu3lrq1cYS3WXAdRWxIZCjdrGq8MtihKuwshROsfI1KGz+HuH/zixrSqvErpA+Dl
vlRzHmiZ8UzJBSvOU3nh4zS2o/yX5wxgISb3Tha0o1ucV+nW3C3TITFA/2nHRy1o
H0LyePExDGQa3a06heMQkCKX5CffJoxbEo+5U3/5yDXeQcfqK9EbTUI4aboeFilt
DN2O/B4t3rtwxUvqO8uhGCngXBnz3xLsMCjYrvt/EYz3c4ahKzVkRrTVI3o0jFhw
02nR9rsQ18eH9CPW+voX94XV0Oe/3GAgHm2U/mI7WZ1DWd5wEjhAHEG5zrjAaRf6
61sQRpHxCttcXJGyjzLNLMLNz8ORaJHHInSypw2B+96PZiRWBDexVM/eeVpnxMys
XTqD4GWBdp6QquLRKzMyu94ec98BEfK7KiI6ABMmLmwLWc4xPrrTKjn0FLaGaoPj
mQdLuwYQPemk93OtWcBud0ul7hKaI1V5VN+sxNKp/VvmRGfe1g8nPLQ6tWCd1WSy
cJ2x1ryFI6jmSC/gM1h9IsHEwLjbnPEbNxR5TzilOjS/aMSxY/eAIDKjaRpoerjs
ZSesu9bq+sat6XyEcoDfzhCdQYYonm7lU89AaD980pIAkaV/bOxY/MO3j6UpzzhK
KObVov42U4xRTcMNwrQRBy/ePfwljVLp16WI7GwDA3Ux6nrMcQxEHmXrui3Hrcq7
yZfKrm53TFyWGCowX++tKuzXI4nh5Ethy+c4K29Q2DfJu+X/WseIULpvtH1utBzk
5nwQ3rHsypHKFZ9hR4p3nzVaRpQw/eGEq2c/KeFUTiuRamNB23OAK4NXx7SOgRId
2HJ4MfbMC7jxi7hBxTgjsArbhhI5qU8ir7y2Vcj50PDfyyDfsk3WtOEThv4ZPCJ6
PErq9XHDhSzd7Ta+VgOL2ogk6B293Z2lORTrZCYo4tn3kKvNPxIjqvfFO/RyrSER
Rw1lStDlC4fj6uv0qTIOWxVtXgunNQB/0Thbeni0OFAm9NK19GTxEidkbDsDqyoV
Sadyh4icdM7Sy5Hvy9lGdMPnlvFxU16BtbM53In5F2rfRvwQRfzdCxqUGlVSwoap
QZVJ5QuKzauQe7S8aenxBzds6D3571ZHvjBpZ9UA9q6wpfxFPI4kV4pWKvJwFvuB
0v6ao39/dM2zhBxCfIytcX8UhHC84NWIfSHKGCKVwA15Mctvm0ExJ8SGvCn5PgF8
o7B5Cqg4sJ6bhKTMKrpfBGjMZR2bAKOm45iaUeVD1dknmsx7jOI1fPfGIe6SQkeM
+0ZJeoDRGhyGWvExFVMFudA3ry5Pj1o2hN5HMTD6v/tMYTB8jH4UrN5r9Mt8Bf51
UWXJzZmesBC5xSf2bQO2sQLbJYfnTasgIms+OaipsqKnaI7wRfT2PwsgWfyYzWuo
GKGfJWzubZxv/aZH3WMDGD0lA72f5YBKKDHC97IqVLrSSOYYFVIAKZ/dQDnpMCRI
JptThPFOQKp9tB2btSZN0OKH2nqx2A4trxHFlplSvSanZXZMB03/Rxk3xGNLSvMI
w13tN2FqnoHulAfJxhWHFqqy0rPp0/0L32hXwIKw/fes6IvhTd98se3vkz5XxX+w
o4cv2vCLuZpFXshU/EylPXTYd5BMxtLlpig01l98x5jUFkh7Z5tYxB/N2g87Ng6b
0EkPw10NM3XHAHLdNOM8fOukX+4fnyeYBCCYSRt8qWHrPOODbOfxhXBXLPXdQnuG
fdq9694WHKgFnmJC58XpYnZvCxrmZlzNwMMOLEilx32P+x6ZnXypf1KYj/KX6F9A
QRTr5JTA/Jf4OntCjvSwmlB1WlK1e6YO45I0savxlh2u8fa+AuNpYU2cuzz0c9ez
z9Gkz0Bkh3ayX+fkf0SDKfadwQRFpPN73Ou/X1SWDAkk5nMQ2wXF/cATk916z+LN
zFcCBuAKKc6osTHxzYyUBytSYgo9s6EpN6OfeDiJEnGNPSkcfmWkqgdhkRjSu28x
dZnGAxP9QcjolKIgc9N9HWmHed39FjubbTq12s0AEDccXh+y7beWqiEFgchiDfXc
9RsdmoxeY6LbhgqJ2N+GWsEP0OBbAyR+JpWMyqcyayuk3QTKH5N+qfKlHNAhqO8p
r1p1+wvJMBgEFe77565TK0h4BVK76an8JXNGRtY4UWyBBKUrf6S0dUZONUwgICJA
pOiHblpK1MVcJI4o+bkiFHqAcIhUS1FVx6hOZ8hxTP2t5Y85kjTBHoM7XhvVGkLv
K7gJzi6gYuoNPGqHgqPrAa7H4so7dq28oZHwEkLkcJoKVtZxX/Lue8bqF27WXAU5
eX/gVWXjbIEDyUX5H+VK9HhUfi3ZrAZu0MFhvnNfmKlJRzVhIQdO5Z76Z0jyQiKe
sLGgdgLRuosU8hv1G+JUGF30Zot0TM+fdH5eveAJjj/e6dwWKE6zgoWWsbNRT2pD
FGfDPhgkUXFCxuBgfO3pO4TV0nslh1LevDueZgb4XgeG6ZOjgzAm6lLjIMtorjtB
NFW5QWk+qncoZ054bwTFV9G9Iv06AhEdu0NlpO4fZFWKzYWVeOXPWAniY1wO702M
w5siJhNVGjCx9FXFJOSRtk7OoLpn6v49/MzM/NsyEXoZ1qJHe+rPIhRUEb9tYXsO
0L+Fy8Mxtwqq0dAA5NvE9j+lj5X/Bk2L1klrjbZp3oxgFtiUysyAMTTyeDnX8RKU
gmYceS1ipx8m3U6Vy39KX1dDGzy7ysxZZuVXVEzMQJiW+AtaqfBt3xzMHRpUUg+3
XLdnnAqn6gZhsTQsRnmEopzpmE6XMCxlz4FqPAS17VP2nBsRh0fmWrAMG01xSRyI
EgsOOZigI/S6kRsOmP69PzeBOF5TsW50AexXz4N3f49/3BHkQkpdDWSnC6vxzgvL
cRYhOsou9tzQaUAAFkAKeqlrYcB4Ib+ow2tu4BwDLRDiVgfXp7W48667zfgnxPJv
2tMvZ024AF+3rI5No3BRHyrH9C53oGWm2FuDSbhQw+ZS3iVnFQL29zyj/+MjAdze
sWG/Mu6pIsM48tm5n/fMNI8AWrGJddAUedjyFkCo+QXUJy3QkEi4rKR26z/eioqY
JYCogOIlBmEjBer3QwPJFzX2qtqaUVnfLwZu/IcCjAbSkG/SAw3kljn/EqvfpBGA
wBc1+/V3BMly/yRhmIuw2+R/E8bXnDTOXRMmWYpYiygzrL//Iu5QxI9meU3E5yzH
0yUMILfpOhXAwwLK0KYE6hEQ6XQV0r4+6RjyTaCKHxYdiZSOzyP6Z1UI+BEFGXRc
ErpLxc5MUi4lQXLi6MUuJjJ/QxhuLtm3HD72KG22oC+EYYIcVZ5TAznvxkYwD6fS
4JbjNkQ1DRj+jumIdeLhm3y24wQNqWitrsLgQJ+3NvdmAsfd8sBI/53+38Q9vDHC
gCES1qcn8JmuFH3uBSnqHNBCDENb5vG2XeVgTD5mZAl9IlaUnf3PVhccjGScM5vf
zCl2/LOF9XjrkP1nyKge9eyvp6hQSnflfXciJWdpe0r9Dbdtchc5U3ZGvxMBmMpa
nFha3hkUqzfbjsepc+1TMXE7gMcECXZpjdcZdASiKR3mJg67TKu6/po283qTuzNW
YRSFofnA1ZAB0/Jxw/qmU6BAA2EXscB5hk27BCOD/3vEf4UV6IfE8gFU58grFbLN
8Tx1A6o7+PUHKcXgE9XUlmgOvNhs3CjzP/yd2B2s1tw9193KkwSKWogyN8+1iHd9
NzLhwLquuu4oZ/pP3cVtoHNETt0wzQMB8fRqtpEfUDWoAg76peaPLCi7DMn5QVcb
/SGID3o5CAbxDPvjCgnJ8NFtfndYb4DXwC2KTI98wWuAI2PVAH7CLeVISTo55URK
Gcno2n/JWgBjAFsMGT8FxlYU7ty5yogLSQvSWabQGD6k123IjIcOtwJQmgbpmR5f
3omiERMZSE8toi00LQslKdSQUjlmlQt041i8Y4CfeAwCeghbFo037Q6vOtZ3tA2K
qalJNxZnj5EnM7dd2JpjxsPiCcUwYsHy/sb/liq1UsrEq6beLTdBLWFlT/4za9db
fSIz554qt4vwtygESILdxIPnDeq1QZd9nassMTSFy1bJ8ErwDBC7IKgsN0pFeyzM
rlyrhEmDAFEXCSCC4OCdfS2vQah9LCqhv6zDYWHcxG4MDtUeQzaSIW5PaXwa/pa4
g1j66nPK+SjTy4RDv5EySNLe57Jj/zY88YWkcuo4ILPqA6/P48Gx7uxvBDf7i0nj
wHDPksDeHqHGrJVRIw1SiPz0dSsDGJXWh7GF/jIr02S0whmyIIBEdAKW6/6g17BD
qTCGWha0lzgtzwowMK8nPkISyT48HBavIf/W/1F+04ow5iC3vOFUPBoH/ZM/Cbjf
7YLY07LydIWYyVm6tRx1CdqE9LIsF2g4s03zKufrWv0EcovZS7bCOdkzrVHyvTyx
AafdMIDFlPJZKQYeF46WQonrRf4scXy3q/3hHTNEM5+dGQoLtjStIFHA7plbeQXB
b/lEanWZlNIxTH7LDVLE7/YQr8YL70FRQoaUwm6gspVfbVo51ujnQzts6r9MJ7S0
JMios+m9Y3T0EaXAydCATCjQFDzwkfB4D386+hKZJoJF92JUGUeAUY8fd/84Pf1s
XtIhs7H1Xw+kKbDKZeUkHhYPEmM0cmuneULsp5wSD6ZrLV0G3lMeFbOSv7iJiPhb
1VR69TMxDsJTeaRsnVHD0qQQtMaT9DlVNmwiwSRbOSulxbl3blZuuHsA4jsn2H3Y
1hzlcbrVUnQFD/iiuFBH5lFxD8FhOsLcTFolpua0ylgj6mXv3/e1jiWUCkTougVE
V4cRCYjQuEHkM8mrTpkvSmKcRQKgBA1Ecl1ZcZg+AKZh+oe5+MGQECm0AvcrFjRA
Rwt0bLtof61pBK5GcvwBTnlmLLteuDxpcrDp0HNlQuYkDzyPGobn3eLz9sFxsDT0
2k24PaOIRbUGAmaMZB16VEZkitujSnwCK53PygJfxpFQrviutVh6I/EQ9tBiURUM
L/0fXK9eBplb5moZssHJY3e4WOP/hyJLgFwvyZlmBTIIG3vAqe7MoSX7noZ/e4G2
fhWxKMqFrk83bLlUwW07MPDIUAaJUABj+3M9VICfeRdObjCMkU97hATXNib6Chdn
Ax95ZTcbmdpdkPT6T0/Yrj3MTaQPjlWJL/8fZRLQzu3thRWd8uvfFu5qYZl34RGp
wvs1C9bsLluLJ8jBBmLqb2jihcUBw8ZX8y6rpCsqowe3T00d9Y/7xIi+wYAPrRzs
ow7JOv59k2ctDZwDBYHYSMkWnnXZdLZoverbaKAl4zb2iOnh1FE4EzSPQPmn6mag
L3zi/D5fE7YcbzcXB/G/5zL/vcCvZBFkcKlJ2svTgehmajbfDQ0P/mRGvauRYoug
Qpms+tqiVURKbvOvxh3+WlmTXiTQdz3v0WCIAR2w74Eo8o0kyun23pHEv7djmADa
n74A3uNS/4dEqaFgIJMvIABLABvgIODp1MrvQyHtvN4C1m1NP9TAHcdPohMwAkeR
NCFX1ppaaKUbo3CID3g0Bjkf1Phfo1EIkIQpS2EVVS9a3C2oLkJwCYWh3VQWPN1y
rm4Xtxsi9EC8ociRWtwzS3TwBuZu0n43b9E1dzZAf4+AGNDEAm8J6LS4ohDwr4Ue
ZmXDHWXVBb4vtfus0rul6TKrQRv2TnaZjahbbsW5DunsPe5TsnJoZohGZ2CdS+E/
wjyZHmsNx87utg+z/i+QcBwJCalFWc22mw+GN6jnpZ9iCtdRrSJEFWtG+6l4gWUy
g5fuFGguiFpHMfgNvBEVfAel9epol7/HQqOb7WVTl7yVFi8B1eL017pttQ/bW66W
xpnnlBs+G5mY6/UeRo+xvAvi+Gtk9rKNudNZLrhqeIx8CDDws7hWTYG1lM3R0F5j
rVwTNZzaiOG6vzsKrVRrxzOIvKwrcwuO9htPhyjGYAJ3m1uK4YIjB+Hcw/v/9lrn
AOC1AfSuTL3G2h8zWejXejqdtPYEM6zvM07d8x2+03PJx1t/18CGS5czFenPFK5x
kmldvTQKUdb1hafjt9kcxY0CAFMHF/prLfoO+FhwO2Wko68IAIrdMYKG0uqfynxf
O/CB4szZ+whlCEOdBFo9wVg+83sD97Wf/28QcfDWTbZCXZSKN8MMn0d0RNZwx0jA
agupwpbUBEIL/cJCqdqeKi3RlmcW+kYraYq8XTZSP44lwoPdhZZXoagC2Q6+6JqN
jezuRLQpZUFkQaKEfQ/DJG9jMMCGWgsV100hqkp+Eb13DK0hsBI7dVgOGNJffvX9
LxySM9/lIgDEJ4TjcIu+mdbjjvx1iSW50lg1GxjjniSS3eVJNkDLdPnsfvlvOYd2
ncRJl/dpYlCltYPr+5Unb6lxgXIzp+4uyEwGtTUvo89o45ssnBzE0kyBDfqOtR9I
HesnVA3MzesLsgDk3zKwa7aor6YQCjFKfbzADMArYkJzl9UIJpiM/Z7ugdkFinF/
WY6KAcgFcOFrBOpI9qoBrlYTuO8Ei8RIuuH7t51xt6keFDEHvUmNtgnE9LFcsJgt
KsH3hx/agNOn5UV/gdfmMo2WyKTHZdTV/OAvfK9VqliCkxBau77UDVKwNBtvP6hP
c1akeAvk2ix93CUqIJmmSX7s8Z+P7TKXmdXJAdRfUJzs0sZWPpsFm/63jsLMnrR7
tX9SvBuXYsF5PqNBz1U5wBNn992Gz66fYj4Bmn6pukcWp9jKijq6ER55h4H54Db2
fqZyQPrB5E+xwXN8RJgtms54UTpgrEVLY6UbxJlcYJhIHD4dXTe494UWQdfEefje
yFizzP3RRsFSnIbTJIxFpIE8U2dxDxMscOtr7znlfLI8FQLu8SiFqvBPvXUSkrGr
ChD6yzp/AXsgfwy3DHxt1wnAj+z1PB1Nm3y1yG+og7kG/VjkLIwBnlRO6qo18tuN
1l1hsPXkOfnXgcKmKc5nkn7AgDPF6myhayzIO1JPtIeyZ8f7X+n/3Q8jBd14L4JK
A7AG1EwzWYtmyxx58FPiWC+H/KRoBShCSInBpZlYDgOz5sDbUsFagjQ7sdxPQM/4
pgtlM6QdYA5V/gYA4u2j8m8fW8WqsJCasJZ3IOqa8u59qA4I30SafLB9+LsyQyiQ
ZS69KGs2fBNGiGE1ND51TB9lRmKw0usXGRS+O+w5CD3lnkZWwbh4ca1XnyX7SxQY
bIPQ4cH1O1ini2PI/RB8DHCKwNbFedy/Lib0oz8sI/CSKL1wU0/kYS433wrHAanE
xwq3GFv4DKFauYzU/iN5B62NZxToEUg3i+6sEV7lzOC/4Vk1RJG/qRRwE5hVNap9
cjFnCMYhvlEfsppUk81Ri9t3G5Kq9+LjzfSjm04SFnkFH/XrlsH95RYG1JtBdpUL
vliGLp6tuq/axYHzstFjPGjLSRt1XY7FVUKr5SMQzn0JrjiB3VCJy/1JH5CdHhZH
+r+qYwKUQLPd2LlrY1CVeYRdy9TVfHuqerg9ADuwLu9A0jeyRcjSMU1Z8RX+hiGa
mEiNunqTdWqsISeD4iTAsp5amkVm82kfx2XART4Qu/xe4/SzANOEZ1U2+3NpfGFE
txauDH1W6XEO2qizjMLmfJATJ5yt6fWnbKXQT22qDWO3XP4nUBwYVoWiS9OU9HU8
fdFSfSpMtl7TYE+v0Q57p+qo4RdIyTopE0DXcG370mhls3FBpt17FlpSa3ahdlgq
tfX0cFyYj5fu6xst9wNli7TMkPtoLkYGX6jmKGRChxd94A0nulgzR47q8a+1Me0V
i+Pxl0Io2t7lE2vXQp/K2GdY1ac2fRrSQh8uYLQFfgEnteCn0SDOYci9mbFk3o6J
CABfAvk62dsgrsI8OPbFCEXjmpqhZC0rVw6ZTbbCkV3GJgGPtSDDMrMwcTOQAWEI
ziQ1Bf+fb8HgCMh1ehd0d6kri21j70s6GRAqqfOQws+3ZRZ2BCR1ua4BiY2dLxYR
C5Fh/LEU1bJ+3KsTyAzn34op27kHh40tYpOtwspDkOuzg0YLkTEnoiEo27rVZboM
ZLhG+oGTylElEQgAGOgmIJEWBeG4D9i6ZF+9k4AUaBVJEEcjm7xg8fkgVxO6nFhZ
e+rYDC/jmwxS8hop+7WtR2o/uvWfRATo/JHe7R+8D6e/Tw0MfNKsrsRwprryOR27
i6HTN/v6fQheIqquJUAxAuP0iwqz8Wi/KuxGzuyZM6nzoaTJCrA0jx/G4vgenQNS
/XY+Ca13c1OB8+y+CwoIxjTPbWy2BogY1B2v6hl56mNaY+2P4lB6tWOBwBV54VQp
BexhgyMf43yVwFxlMlZtVS9MXAlZX2K+rIktmkSiDlID5a2fEqyLHb3KOlw3gpD7
0ygfziKkRuOUbQzoeJVtgZxWm5lsbpWuJHsW46sItIcl5t7teOWwy6nzPOYocyC5
nsl6Z/bkwuuoqejyPjEd7GwGl8i9tqHvXCXRZz9WBxavrLB/S/YPoJhXBoVm8E+O
JROTQrVQnlEtq37pnxyfTYooF2tnQ3lACqu2E49FltdNSNevr9c3MHkcKguLYTeL
+orbUvbqZmk2LBumcMhf42EKuhpPlLQsbZgHrsAuiOefdOpJmMW8c3ejjYCjlO7T
yggbJsNVI3ar0Kesb8aHLDgW0Ae1cSP3MePW7pJAVfQttlLGzQHtsCjRdTHe/B+s
FgErmi3NxdZpDbmOCeq2Km3icgo3r5KYjasC2xZIoQ28SzfdOT9m3QRk2Fp7yx2g
Vd5NmKnOkBiienJR4deh3e/XOMPaQZtf6PR7H8fac+gytwJCN/vl7uVouoD7bR4o
+5bLVMVJKZkg/aPx2Uawp8kBrXVCbIn5pNeE/VY87VeLkzQ8FaQSdtXIh+XbtgzW
FcZ7qSD/nWCSqRRQ463KKKPhzgCvJi8y5m8UnwVTyEro9H3/7Z0yK7q4stZSiPzh
sGqny0JJg8b8pI+Xmsf4daZCKon7xUNHXr7OEQFXGZAi8ZGg6oQMy1eP6dti6ME9
gT+kdKKPhEHdh6KuH6JlyqCWYhm2HbUPRC0fkxW3XMnUYgBSCaoQoG0uUQssqPH0
9ojtL91uTqWtkjJP9id+nxiD0SaAcnMvsCXkM+szs+dvnlBcnfq4L81zBLbGdv4q
ZVe6T9z1ETkPhBVcNDfv2omepo1JBeE6brvciD++kh/+mX7NFcBK/ykzgg2nMKwS
NfDkiddHv29Tsqb1r4rvblaqZkBsB2ypW3VZupGn0f4f/cT4pu87wKH1rhOfRSa4
rPKQzPTRvySC84WaU+KQpqYwdgKo1LGa0VixS8uYUbeE9HeB8gQw3lnz+41S+l9J
kOvOQFhWEYQ8UMrCwQijBRthnV95EMHu/kXlfGSoMmuT4Q5jtKHt+CPdRXLmHMy+
UK8lwZKq7Aag7BXlkaVVW4WILtnERS/NFb7aLlXDN0o9ORZw4vPwzyEXkSd+fyo1
cS14lSsNOF+Rx34n8R+waFYnVIws3Pe63fE3S7umTSyne61Tm7LlTp3jodTznclh
Ewn0m5RW7Qn79jck7V1Ch7elDX61gP/sxdCkvr4PIvadaeGHyBH3AVj6KxYJo3aY
BKmbBld4/oQmEXCnDoHWmUyq1sm/RJBWI/jsjl3wJdJBpB8ExONR+0JSmDGkcxs8
gYGjuYqWbYoDSj8ae+A2HF1IPikwOnvylIiXJphMFO1PIY1YIkLbUo5aGpfooGfE
6XGZm9WblkVaOqZk/bXylTtKcUwZ1x3kimazCperr8Lwb75kpVl8v5LzxuiVq38B
s3FaK1BbQwSYwOg5iTAhBDfQ1XJSprzMVBu5o1hQOhNy2eiiOTnznhGMlfdgKk0q
JHsbUglwi7KQcfHLmaYUGBg6LtT1Rh972nRz3IpMJ5C9LCM/GaV6A+ZNjDEx88OC
hSXpdaFMnzLbz52EhH6IyyffTPEafb0lp8A7EboCmpEPGfJZVEw72eKor8du5Uj1
bjbOZjH49JVGjIv+SJsfSPx61V4nBmebsYjIqBjrx8kIhAh2opOHYhKLH6osz3AR
UkYRL0sxUishDyzxJ2NLqDP8joy01maev0Wto3QZqj+sI0vOC5HvLLKecqOk36DQ
2Is8Aq8LDPJxizxqyL/IFJkyQiRi1LQ1EaMVDDOeBrNgxktFtd9vB6KPN2pPnAWr
Isfvp5LouYnldZh3v0/j5UCqIJwNfcFVMLPsLEUbFpDWstQn8aOZLdyNfIMDzHml
P+1XVt7uUg59WwUrtnQ6P0RJqEvhYXYu5d4Ll/HNzK0OD5qZJ4rqbhF5wEHURktI
RDkn6giTWoQTb633NzOar9s8BA08EzA4tCCmBDo7yILN7jH7zONkfTwiL2Ideuhn
vxdfwSoxVeyHBDy2AlhCvffgm1LAqHPZEuavbJzvVPEmiHBBLNoPOU3hkxM6MMyR
WEyph6eOmCYimiTWe8YD4MXXO69o8WV8Et9rb8hO8HB51IMuFQfv70nSTMJLi6sM
0LrFF98lQaKXiZNnvfzVGKZOJXBxDhare78jpTQY2CbPCbBepJspQ89Q/iB2Opw7
JW4G/N5hEMntEbhETcBU36UuVXA5iaey/qpcbMxEM2AW9bH9GX9Pt8EkJYn6nuzj
XWJPpAcicqe1L6wJJYixljnPwSPj46E0R7B52JoSxdJrnWwgEq696LOHNmdIekZf
NIzgW6KILm8tu8vd+J1opc660oM32NA9rE2vRO/BJwB/rhJqzVSgQbzN77ZV7wxr
DnXNV7OOelQGjOxsCTpriEwMsnAvG12v8ddX/Rk6Twe9wgcwriRaGehgBFfAsCgQ
/t6sx5BKjfZS2n4N3oJ8N0D00nVMjoV14cDs89RUvCB2S1p5aMxrYAeq+zZttZGP
rIKo+GvAi0EZGjWHwwiPZ0Vf8shE24u8qs64cAAlUy5Axw7kWt0yIlJ0zdE56D6i
JYFEQRicepDZikLHNqwruoDXaAVq9uSR/ogLKqxL2yrpc6++CqQAuI+BHk35MNXm
/YBbTMFxmber1KuOdAaQXcThgj/zghYK3W8iRfKQ/oxr+HZ/9kg4vJg/nPm5oX0Z
6NSrNp/4iFB9cO1pa0GGOVCuv1QJOR3RC20yLQKmaUpP9srry4uJ3kXyoVwLCTAm
5Z9+lH/iWbmnX96wUM+a1Li+Qa5ebK7O1VDhHuvUl4gHmj7kkaWUeuQxU0u8IS8Q
59dKZbfU7smnAKam2+Yn5huXZLfapIDTgAdaZPM6oJACv4wpcDd9P2z8aqIqGYt7
oo1r+byoFOuWLlmTDcEeNQMFGF1rOvURmkp6UOfsqGKnZWRO4uQFJquzj4Nt2Fwq
30SC7CulwBArdpxxUdmUYwtWJSaBke4ELe5upa2eCXhoBH6ygCRNu/KRFMUbtfPe
0An1u01KFAmrEZcTs5/qWsQoeNWeB+ktjE30UxBatt2PyDhTC4FbNLflB/3GQTsC
pD8eNWOgLq7QfvRQPzfn+h7DRGhlGDW0rgi1NkQhMn7HQsaLOPyV0ADuOOkc6GJ/
9Xs3MjML8HmANJrmyBpKP/xBYJMLgzsfo6+KRo2fJ6/DFJiNwmHS1OGjz33CRGvA
/6S03n6x+bztTNMKYMvRLigZL8CuofWsLeHVgzhL+NHM2IpQ2vF/taMNRBNPkw6U
P1qYyeoyEDVQMe4Kyw/E43jNINiKc1x/qq1VinW4s2K9l/o3nx2KlWAcY+OnpicD
m5x4y4a0pjXg8WWot40hQfxwSyjOCN6phW5WE/0hll8DFY+mHcXu4YprCdWlNdBU
wyQNCrgaIVdZ3C/03nRD1Du8+QbXi022fQQgFWGMrklkEImQRrJzuIQ233E4mJ4s
EXstg48KxjR8qLm9jIYR181kPDbgil0DinfoulQE9KbhOeYJqohcLLa30xlFqe7o
ziOyBX+ZvdPeVSaznPJO1VcP0KIbwRpeqAk3yHSC+9OkSGYk7qd7enAK2uUemW47
KoaAosn9dm3BTNhe9eZ6cg8iyZvU+UA4kIe3XZyzF5IXnsHKaZlNbxq7btcA/KN1
4RBMZApUpe4G/rVNZ4GuoKjyh/qbwgFMpK4CKWOUsJhsxupgCwaLMK9MRfcE3AQC
3m3AFGmf8ft41121CXNSJMTpqvM2d1yj7Qd+gWiH6A4Jn3kZpqKoPW+iwsY36B8v
QxnLZZeeA7y+OiK6wcD7H5iqcKLLn1H+fI4eonskmSss5sjfntQYtmN+fkcUyYDP
7zo43mw5sQTP90zTQmcFvQztnCCRYyagHnszW4vcTxEDz1jO10BkyVWXtIMWH3c5
PgCFNFBflaTJbBtTqFmnH9uNkTyhd+U9VyWsTbu3+X1AWeDE/U0VQMRe1PwkuR6N
tSaCPxQ7NSO/2swRlqD36vBpcctkLvNr/h/6CSjVrOCHn3hBMJ1EXYCan8y62IFW
ZNRhEeaaUVIcXA3xGN71mB37tBFsvbP2cucV7Aemetj076QHLYtGmg36LMQHUNBV
uxh0xUHJ99Ed+yZQ5G6HKEoNdBm8pbeVM1ZHrMSyUJTPmdDKsHKnXDTFBm5I1XBv
tIEtO0B54wAsp5iA91XbQsYDXJxE3dmdYzKnR1Ua15A7UfjUYRu6m++CFAxd8wYE
gOYUGESodSFH1e0trMooHQb8mRjkGv2HgiAH+U3YGECjmp4b243+HGVV6kwwpXSP
kPBN9mQJSX7YVFOhUC/2UkahUcz3sxyNIHbDxnVZ+ZgaDTkYDuu/dQlVCqS3GzNl
hkGCcmWq9IMLfn+jDafgJHGW3TblXl7U6qGyJS/5q6rBB/EagUhTDxxFcST/gDd4
cCRXoDQtclGNgOr9uL6OcS/FyrbzbZjmUzJew1HLfa/NdcxEYhyg5mJ5DcqFO4K+
G2W95KAJ+MX8M8uX1D/7damzbiN70QHAQQCDC/yo4vxA17QgqvN3YvxqyBqo5RUL
hgNG8xqBIk7YBkwvtWsB3s1hmodtxlzXXtyeZ6lZ1qiVAIQ1H2gv1iTgkueMa9qC
CXSF6TsuOjWjoocb4gfdwU+FtvPZFBsJmxsPTiSxJSuiPDwNJ7WeP9sGm1YnJ0ub
FeQ6K2HmgWudK0z/OrqdXgsPnn50wi4o3ErmGWwKGKO2TeM9topRgFY70y8UgZjb
/dIIyvHYph8Z1X4E5hxLbRvcmuD1yzWoRM4HB//nnvuZ/ftmAo7/sflZwG7JgrNo
KvFTR5Ux04aLI8SJLaaBWVSfYp/DW4NLYhZ6SRCWe0Llr77sd+e8Cs2g7spfm2ak
0stuM9xdAakrgIuMVSEsKaK7uOZZwIAQdDYf41bv1Zf5qzisg2AZCe3PsaoPZBNz
12ZhH9jLsFMbJkAvzimEo7XAYskKw924df6GSEy6yYVnAgSASOFqCZXXoiRIDMxD
vP5hc1ySXn2MYFsm3P1Bk3hHEGRwYxTB6zF5VU9ptK/FidhK+X+g7yI/MWO/wAti
b6bp3rPuljTVWu6dk842i8l9+q7wSSWiqyKm3SSF0nC9OP92X9y///oADoPki1Hh
HoZs3hWgUwt5l1JyiGblt2OXpkUmQo8TU1Iak93FZosyYfnhAat3U/FiPNW6mukH
RRnX55XZKhfih+pHUCnG8JaaGE5HL1ptVrm2Fi9G8GD/iET/c2EJMZXxOpevGMlg
oWKmHAfhsWsihhUDucNrBK/41zp+wVdZQlcMeL8HQZ13Qsrmpn94dk0pM0+kLFj1
VDMsOaEcj4A10OMx4dlYtIEW3NtIncuMnTcHOZwneUSeRWVlDkEG3m7QVrCGYTUo
ZDh1g2T7Py7lStTtSjwVAkRS1jxMc9fFFb+2OP5PU/7+n+vnYBukeme17uWrHeG5
ipoqV5V2+cKa8/NwVh8UUeXOInaedj75vxuMs2Lk/8eElTQScEHPXPPZjOd55KK5
Zd1AhcuvO+ibp2MPticGDENWv4AKL9q9h8mjBA3tQqRQGDWcSl2s2reDYlXcngwY
Lw6ccg3PDybFlyuulDuC3lFVfFdzHzJWi/+tpGf1P6bjbych7DOmaYp5LsGF2/lJ
Hww/H+K9HDOYcdmZrAg6k6ULxsJWAYYmANikOcmd+CQK5vEhbTHrfVOw90MqPI6F
wYiOuZMvcaPzh8dhw0gUsP1AzD4cnXOyw7mD4Ec2GSThiVsDvHVgyEdLK3DUA32A
2HSAtkd1UughAYNwueWwZPH3VYHjM+I/rEjLVKaOWkIIXNQFX2DGWiATwnwrpaOj
vj1IVV3+WV7HU037zzwJResOQtWAPKFfccp5zXRE+b29rKayp5UFe9q6XLFNkZaC
V4H+NT+JQzq95Mh2nZAAEm+HkQ6z5aKzJcFlpkVYtypi9FA6sPNO0Uh6T7gllNcL
V3QqVITwf4X0UTp/GNR32m6rlrX9Cl60iGzvfg/u8lu12Qc3VkaHdtfs4km/Zcj7
9b3qe8LkTY4hWF6kCEuN3pTaVRCWeMYCMrWAwKAVhQEGk4ZwqWK2RZdBoqrmsoZt
vUufC6Z2quhJPuq1135LqdCC2hfW/wC7e2arJHpon2ejiTo9ymvibcsckxgy67X0
9YqPPvRUf0mBnceJF315XXIEhMmZu0z2cmSCL3UcaU2mmOaC/K3BAcpJtI5U5D6c
kzwkK+SY8REGhm0D3VBS8nJUpy5YmCfE1YQmu4g/CgzQ0tc2CijJHe6wJPrXfQXe
mXl4YaU5mt78lG6m3pew7lxMIMZ0RTe/SuYzl5IkclsBvHpVgHdxJvW2kJWmdm9Y
5ZlBHrfEGsVPc3deL7+tRALbSaHYpgHwxnaGU0/UJxvQo/qEGQ5PXrU/MMR7Q7Sr
7vbpxdg6izSkxIgLLi4DMvGK56UVc4dtQqlXAV9VfFpRnpQ8vkbtQjJxgu9Lvccc
rKeklz/VRSE0d0FwITj/ECGIcmAFYSbsT3JVppYmQ5OFPzLPXdv2wRBiFujwyHtH
srtc2i/2wnKU/1ixWWMJXmYYwkLXXNz/Hi+Fucu+b/IgjGYe1NDv/P/mxQe2iuJj
lIlPCaYWuFij6hUDXFROE+VPXJvsWO8UuNf9RnhRyTt1AlBdlJrYkuMODDU+sIDf
eSH+22f+Itme8CfuF/C48rGk6HNmkd0gng/a7DRD/iTBO7PxloFEjeTSzVeT6Lke
9835lxxl1ZpWdIpOxKW9PVgPxh0XiAZW0hpRsg+2MuVp2PuQK4WZYrJboz9Tcsk9
+ZqSBbkbCKoGrpqZyUrS2fF+DTuCxFAvJWJ4ZFRHV3ZYXWeWOdqgK7A+j0A8Ub4Q
xia6gu0j8xeoTygdYoqH7AjjcG/abRxbeg4KRwFrHMI0IEMjCcjDj+PU4T9YlFaZ
QLmfxv1WwKNtMRZUhpgpoSwbBXDVUWe0s6fQt3brPpuhsb5gfnBd89KZnY2GMMyo
mjnxJ7PUYjmgAO5WPF8FUFrEYn8v81Qz0qodJQnbeSHkm32dN0Q3RacHSfQJ0IRy
rHltsYu7ohf9+6ikARpLe/cj/skR4KKH5Gh6KTx930FSaV8Ko+H/2xnx+b/QMonJ
w8SQU+kg6hP2C+YUa3aTo2PI8iTlI8ZpfGRadBKrCWOWOqAy17C3XVsYsMYP//0R
Rc2qNJBh2aeWCEqrstPSIKKYPol8dx+/ROewQUD7ykYYFdmu5L3tfiC3rY3ZApCg
OJDyC6/S0MMPpWLFymkofEBXl/znqnQPSGY8C/2LzFf6QEFMmrggK7QJFcXYRo29
hwoZ0scKDyiA1os2zFRMDG/aANWrZe4SKVtZJFFL3GRDldGOKpAMrJbK8+KPC7Eq
RO++5P/o3XEoI5bnj1KNa8yGEpMH8dOwU6cdIaysxkjtmjwE0QaM7XZDDyn7ZgX7
32WKuRyWI1GufIddZttqtI+jpFAVg7F1kE/PkAE2FHvZc0dclFjNK3VsqppWLsaq
pxPOF6EVcp3WPTQWl4RS0s8E3t6mgfEV2b20Tu3GzzLzwRCDQNHT9a8QMj3LvzO8
7xb6dSHLfjlm1O1bkp6BANiZ/hoCaIDq40xTxflb4gLR9vKqx4IgVYlCUlHPUy3I
T6XB4eshlTpN9u0j+4xy5JoUZZ3n0B+fbTGUeWNze9XxDCYejzGCVSMYbBSUNxN4
fqmZQ3xc3fVAhMfzfVLcTx9q8yOVD/ewerCxUYiTvxTTaGcUOEJldZ/zdck7Prj9
0zoOZLsihSqg61H344hg0tnMgd6jDnXG+wb0kVpR7PDyIfWDr5nt2RMmM3pg4xtG
Nt7mBfkbiXU8nMlai87KPUwdZR0UWWAIVV5BpxbK7l8tDT6RvRzfggUKQsgG5mn3
J+Ab+3cY2fSQwymYa8mUaEg75qLFryaG5QsLxKX64khEhni9us3XDMg3F9odgYyA
PGJeoRS2gbGNpLdVSnb2ioabiwEICJLdn2Cm+wtp+rF4SDHaCttRjVtDoX0CSHzL
6t9rfId62zJDIDoiJnIRHkeDph/XTZWzh7j7YfaaeGVejJXs3BHAwYM3fF/MRDrM
bqL3zfcYzbL7nBUATZA2Uu8aeE6JOKrcTaWe+gmMzCvff+OKIYmQSuLNwHGXcQDM
Bzf5jG2PN0t2skcY59PDLOCHEaR3E2UapEowA/Ad9Ja5v2+8BQBJ2GBBzo5LW0sj
GiQTFmWCfJLcpCkNgwdQWTx2mi6zxSEGpEMlyCKV6YHzgpMhjrU+MTTWJAGHl72P
GMIiea1cXZ2Qsd1BGq4jzv7XWovO+1264wVU2+ZMMpHCEPRFpf94fKyB3mc3vqB5
5Ope04dzFynOk31Lp55d0a1niMV6WvBVJmckw2KKardIOD3EX6kaR3pyIoXkkIg2
6cBK94a+t6+N00vyNR+FokHzCi7HRoA5E9isZlDByOU0u9nBCE3zKISF5WzOfG2g
dQzKlE+5y/wfRCbuqQjn3G6LWOFLFG4YEyXMSdgqpZ76pZAbcfVaQafsvQX4vOvl
HNpBI8vw1xfyPM/K4Nh739guwQ6CgVi1+v8qDnvYVDuiYuHsXVyTzGqNMvB1kSKL
2Co7uTRyY1kATA82o3DCZ0cntGsfFgQI0Ejdf3UTrPR1LQBo2bXycrWm+KrOzrhh
AVp4lqlDLwIryAf9RFyGAhjLaor6fZYKBUYq95wKQJ/g16rPSEXaElXsEi6j5ArI
wXDqMH4fMjawLo+DoeeFYLaF1H+Uxx4tgc4tkzb9jKAZc49TwLTyFYMdn4axT4Yz
hXtbCLdqc/ETBB7VgboqjPDgvKWGaymeAwhXmPJIc96+rytdIlAJ0cfJo1HkpuMh
qc5hBJlLwuCcuIWJH+5x4wpY8fsHu7fMYZl3KDuPrQKp8G3DXSoX+7bJ2j65RPpM
Qoa6qCju+X8e22QYe1Lg/VLkZ9EBo54vExU1z7bQD3SKkyYbx9GZkz9jLRqPHBHD
hgQlszcSpZT1YEfsBIbyekR8i+YPTpx30IhSEj8lhNTmdYsR01K9HvmyHOCLlaMr
2voqy5miPaEG/uZ3E6/PNlwQKV6jjIGDczvOk9rB5J3O+0TLx0hVppOabqRkb+Za
Ak4JVFoKAZgZUc62KOhL7cEN+GFG7a1orQMm+R9iyeXoiKmbioYv/BInqsR2NL3X
Px+1QfH4pbK6pVsLF7RjDWmRdxy6pk9LgHo9FdI9tj290MXV/ICWVvP+dDzutoJz
lbgP1l6cgrAoCmNvEh89izcxG6XRflVdYiXKcPPiMNjn9Z/RalJXGYD1wr8s0br+
9OpTeNB5HQgRQs2qBstQ6hcY48kfOY/FcmkBaLiMmQFMGpum0hkD+DNyTQBWr3Bp
NChWwYBKNZ5oCnnQRz2av6ZHjvcjy6zI7LX1tqgJWgjkRI6T7iku/kuY/JoL1A7b
5HOWQ+BMFCcDSQ6DnR3UT+IyRc7Qkx5zVv+e7mKV5yAlDzK7W20gPfj93l6Ylgi6
lvsXnY6vpP6ExwEDztnAaV12r+1rIP7/YBr6Hx/qGh4BW0PPjYlXkv8DGh8He8RA
oOpjNUBF5nK2YelPa0iYJLXTGlj1r0ggSwRSA2UdeD4LScGG1ClJNv7Nr3sWvCUK
RB0cW0sAJbdckWD5AkG8k5HIt+7ET3OMzLweSI9GO8+yNFHzeeK+cJbMWxTYvirA
xa7uc+oqv2rUCVw+Awd++gZxFbE9snE1xtKapMWskgzl1H33KsBu3UCQEgudIvrd
Eh2PqMpd3XJCPR/AfXy543NpruQSFrvuk+LHgaMg8aYFxvd567pw9WA7o3mmv1KK
7LDcnNTtIdqedRVnGP6O9/VFr7hpDXzqjCIR3Sxa1ng4xMypeoM35ldyUp+wk5VF
zu45r+0qC63fiR9id5M+47KN2FB/VEr3MfVL31QWShMGDxxgnk8Uk+wvyKwAl2T7
rOtlaPfk5WWuHNpANM8gIQXxz3qJWJM7Fb5Be/8PHpE3fgAC8hyPYAl/Hc2JbndB
10OBCqrdU8bAWdLx+40Kk2FqtpYFZa7QTlJ1P0NBOYkJqm8nG6arsZsp4fPM3HC6
bICr/aYJHuBE+GFBx8UiwiBy3tgbw/vkahsjLrgtpqhMxnVFaF2y3n2h7332EF12
n5HOkcfyCV5YF2KqRRmTO7QEx5ViMAmn0nig1VVq1hNALI1sD9l2hKA5q4FuMvAY
TZB7HPAuXRjpjgAekdgZKMRaGT3Cxe9zJ+PHStkWQbXonYl/gHJjOyeXxPMXt2mu
wQnl8zmdvLnIyRzWup5kZzyHtWxOO4ycJJhrfE5lG7V+nbXviDyq2MeTX+dSM15Y
cGrUdiTGhoe/2J55S33Yr6afDG7KwuFTtNxBs9CjhR5BGFUcQhwItlZTtHriV+Ol
pC0HP/6Tesca9WyDcbC7VTWr01giK2YVuEZgU96UShgVdAUFGtnLjGQw4HgaIKid
GLBElwsmPKiwVJWAf/NN8l6Tl3yYelEUvPzO3sx6SEcOu27rrurIlInLi4JIsLlM
bRIYYxtYqr2y0JiHeZyxdd5ECBxY0BPMdulqhVurz/15GsfmfMPmdDKRNginxfZA
PPQTVfYfOlyqZfeJAa9vBEORMu/LHLiXYyjirTMNRaeUVVMzbt5vyqVGOxdKSj+/
06v4doYwrWfkxSwF3bzO1YHgwrpuyftm4KQyPuX7YzNSxflQM8dodH7NvftO4fRP
VtE9WYjh35mr7Qw6kh1EQFSFoEUGD3mANc2eVkZayoJOSMa2Qa7il+0nKsRSnSl6
wPoDC8yslgMgahRpijIRH13me2l4YaPgS2drTdlfAcloXGH0bmfR2CaO3sfaWfgl
B5VlEEPRRFfE4Xd/rRLS9OhV3moixzsy/CC4bM05UtwlZeFRtG12a32zMDxB6GhC
QaDgpHFPjey5kMoCZR3h0JgS9qQlypKcuIKUiBQUGmidHrbFZZ+639t38tT7gw7N
BbJA8jzfihQEX0A8NJPCTFyrCAyAcO0ZV/u0lZDslXiLNtWOOcmm1D2m9BmsrE4I
Uy/F0HrxorVgn1pmydm3rC8UAUyTW6Aijg/MKfrVaEOzKzIhwZosRs8li2fr2Dyw
1G/KJ/EXT1h3OCn78WYvsnmvIUbVEVlm5RHajrcSfiHbAkp4g9Zum2A45bElG6Ky
4g4mN08Dp5KsGnBGpXd9prWwf+12PoJVIeEomeAwu/Ycj51xI2LYk6aBXaQVOWrZ
ppjwmxAy58+Fw2GqVURO11cU/bbS3fRo4633jF98Jc9t5pF0AiGGw+up/bcyg0nw
eTOZqqfdXnDM4BogmxuknJvZVDjgTXcQpp8HKtvm6BSfL5pj/Ksmnr1pazRFlPwW
AI0mZaciUbR9ruvimMYWFQwxkX8ylLq4RQxyBTdJZAjxEEfHxqxsMDrYCoXdru8A
6ji5megW7GRd8fTUjs59jeS2b6GUMDKhWKxyGL4kZblGRVNyPL6rrfrRiDyaI4L4
E6dmbn6CuIBDYJ9QL9JKsPTLGDpV1Okw0KCpys1XJ5mWTLQjns+wd8txZT8NooXi
cn+thVyR6BGstMrpz3M4CwqzKHrNtgynof3wRWSRPf/w0VuNgOYeWIcyhZz3bfMO
yCavf970y+WXoikh+eefHm7q2Nc6IpdUj5+z5FdNRw5cXMoiUI9Rv7xuKI3R0s1F
r04i7+3CS03rN82VXJV7hjr1JOM4iScXFOtlXyUfNeNkN3E5eBc0hzMtB8r0H74R
VmlWRzOGd5PSvm4aMu5rsWCjrFsHcIquD0Bhutq9c6Xncenr6eRsU/1oIKdepA2j
GYPZWxqph/nTIQu6+IW5W38R0slRI/cBrC0C0eJH7/VUSkDdO5TeEBBtsHgsqgKn
ua2weFdDpTJxaNWI+uf5/g5OH8DV8Ftah6/7mSH8WYKzMwBdzewCQYyt3hOTR5ZD
JpjqmnUd8s5LqfMEtYASZ33kbp4BBoctXeNsZzmoenMrjQ6UJlAgqJscaoJcIO5S
k2AaJZsUaRJjMRnheaty6gtvqnbjZCV6WhWrpqUGyKPz3iJcci0/dX4Wks94OLkk
jhNf/cvKqzQY6B1lx/cjOAyUdhO4llP2SNLdXE4ueHuEJUX/qX7seT5/vMC4la2Q
FqFe2JUywJyi8v6iSo3Qfa92bAsNOD7B1Z1vx3cEERtboeKxIY3Cn5yDzLAHyZUL
NMCV4Wd/XJUXKqbMLbsldZR09U6uVQVMGD7bKMN/JbivXsawkTVNiSiQaN6EDu7+
HlRbJUR8fREU8zZuugoYaKO/fngtkXo5Vzq1Ox78j9BdMluuUu66Re0hH4S7G/Xg
saROLLY7krhxaOnLWpWgoyjjkEoG3WIGwHqtuiPcdAIyNXIr2tIiB4lggnxf0lc+
TMBAA5GgxhoR3xJq+D39YplaxopksqyFwoP0tnmmHHj9rnxXICCkr6hoYwdlHsgw
LZWHwb3u42BU6SEE0zBoQl+QX8hBhaGzP74theDH/kcN5o4Pi7q5jIVEJpEfUkOE
VHmxlFL71YSS+ia+7GghNZKjmBKFW/bPGkkSBY+sl7jYDGCyQJeaUTG4RMV3FNa0
WFYKNuhg+/IxjUJjbEZA056PB3eRDWPi7sKnyLTxLCOijq9Ek/Pa0uivEJA/XPom
d+C6tk9arwdH5nfkk8X/r4mWOHYodvdqLdL47kQfZR11iGaj4HzI+f4g+LHAmc12
EdbBpNutkVdmgxf5SP+Y0Klngbsf58uSnofB1M/XMlclM53QdnLyACEpDmC6zyJp
g8f+NC68CoXmPY1qUFZSv3vCfDwMGj6rm0yRy2B5VdSL33O0gXo56Yqf7/tr2x9o
a1Hdbx6hurCO1Kcm6y93dP9R+QAIcEQ9b000LQETnVxDyhRF9K7aujxQzeoaphMo
MjSArOpi5yynXlY2hpZesCX7hAG1jD9dq8pRp3bmgqNi5KzLKX6jRnA1m6UyadA3
bf63UB/DOniZPa/0CIIG2jmVYR+yYEtFumw7HQAmD8zLYOcgEuXNk+XgqFECRegv
wv5yRauiCPja2E1TG52NHsNzJKiWc1wHnuO8A9L7bnMs2KGcWyN2Whroz/XnVWFj
/vrp1lDHe9IfXkyh3XmbdSm8RGpFTNg0W0GXJhkGCzra8kPoY6m/HEszHqaqp4W1
2nOqNvsqUCAbei923WzCkcDf4QR59BjTM6rQdHPx8+961xauT6brmjsBHPOTIXH0
KByCMIsZDWXFg9a3PFEXizSIh39pnNA2PvGdkL5ffiu4TNVUYGX2pjo3lzBFFptm
FnQZ72L++WjgqS1HUEjPufVx09q3EdtMKUfsanG+CRLb7QfW/sjM8lspuZglLbdZ
KY8RdMZmx4tCXHj1uxNZn79LC5zKIbZdGPZoSLgDhl1RagKyhTnBmKZI5nYiFpbk
kDNiVrv0KRn/4SS13rZPSpSyTnDPyeS7bgEHiyhjNYnNICJ/Cn1XDndTO27qPBXG
NtCJND/+veOP988jk0rqODBcEOzrIjNVcvezkEqNnovS2lVFocC/vt+CRVSYVUSb
pbKoI5H3k1IzwMugCCcLkBLAmXLMLnAQTITKzfx4QbdOI/UuKqq5IstJMQckPHVw
N2QlEcPrh+3kjBD6CaNeerLE/Nd7fgwBmKaC86AnajW7cJDf7vFkyhDGoemZZxS2
3hRn2zPlHGzZ2LEQLShDiiVQnQQLBgD9zZDzsIXberwigsUJRRqzs3Gc5bThN7/V
hdy9tdy8sU4XQhZT0lAey3OlM3JneefLQ4yCf92tCD3FCzdMq2WBFKjAvYZtHluz
fsExYT0cjsu30Pfvls9WrDUjmjFoMUEeEe+bLLX4S0mYpaPJUwkuJ3pvaj3XWwK0
kDQIm/zwaFBn0Uu2YOMLSCZJbkZ/CPK/JOp6Ilzrg9895nvVn+6rHNfqnu5p2EKm
CeUaoPzDR84+SQlUSdIp1ZV3VUcIanTNB0fN5uTJWl0lAfH8aRLi4AbN9mhvy0HN
T74VW/pfUTV2rxqSx1ZMqw+nbvXRw/SyjgwtHiRlNp79SmePC+c/M4sPXVv59Ya5
MQFWJ6qOBb6rVAfrBla+QIiAV9QEPq/y8taMLw2ZTpj44aRAUOAjiVBN1StdeSbm
7QCzgE/0fdue585x6fGqbsnBBbhPs9g9U9xzk2w0Nwx+NJgougfTLXzvMnbpXsww
tUx4BNQ6tmROSCq9TNZZ4GMhXvMah6O2p2va8B8hf6mKAy6ZTeEDfBg/iS5EnPoo
BNFrGjOm6k1Jtj4s3STOiX8yO8KYati+8+/XUeNGnwewm5jJxPocSkvLyAmuLrZg
seZBMD/N67rXgHMuoHqUrxxgkgxZ8FubxGuffrMjVkl4XOFpLHAKObqNuUKvet/L
rFecRtfufsbyNoANzQXQf+/V4AN9Q21p7pz1fn8JNVsWO756Os9M1v1WKy/7mfA6
OodVmflVqXRNm1BaWcpk7mZB5KEaxN1tGwQDBQMejlJD0xKKbZRxQht14nyyrUuS
NWz3rfJF65l2hyTRgI+U5c+cwXuj9QFITGMEdDISM64XL4mq+qGDwvBVZdOB5EgX
UHuGnLEahbJCDpAFFx/OSbiWkaTN5gHYjT8AAb++maipUsWo+lnpbIwImr2qYSVK
kKCQEZITNLkLMkaRfWqZ3wa7tSy8o6DCWP0SesMWCibndF4RwlMWLcEBKtspLVKq
Z8jqmXiaXYEECQ/UULIqcLZuZY8lB60raZrNkEmqFSeFbfDzpSZLyJSaKiDdeoOj
/IgPg/BjUe7TWf2rBWyCHzx6j6VM9yPVaNNrPm/Coc3Mum/8Amj1vDBIp9GknGl6
UjHKTkx9JkthkjxwIsqLgEmv6N5TqVZpH1whCDzj9CZBzIcHiDv9Ec8ha51y5+Zn
Kx4O+lS/veIyvckBhXI1azFL97y79bSXiRLseXhFK25BBOURbMy8Efm6v5wNPy3h
06kskZtpvBQKtI7EPkmvSbR5Col59VWe0cbmuW6bMiMnwnxZWdpFKuE0eX2ex8C9
PW8qYJLSkxrdwAqFfrXAtnqTuyHSM0DQIQtf7mEuu3+CD3jEj2s2yb4zdtKNWDd7
TdjcmGbB6VfRIII+rMmSRBXyKRI+wkqM/rEgLBCsbElEgg4ol5BqhocT/d7aF6co
wHvNXbiWL9IqS/y9uLBD1WvRoG1BJjA9fxdsClrtMr+N7wWIsyDPNHcQDyKmE33V
7XrCER7XlNxZzvxZex7XEBf62DMrMBnK+uwuzzmoVLDwgA2YNBqc2zI8VAiI/bA1
32wna/QSAbnzXA3nH8iOvnnFkHoLrXuPOD0cPrpviynVlAF89ovsuSlNttsygy5l
kAnKqxXDU2cT8oXbdU+OgCOXcOqwYsIa+BibLBVOCcJBnT5n+ROwRcspOTL9exYm
zcKICp2mNSFE03o0JyZC1iDCjV79liRymYtxb+T54ls28fi3bhPEtn+G21OZw4IQ
UZg2vmhPSW3v3m0+gT2xrYftMs78U26tfqhdsyUVPWTYO49Xq9owJrnaDskEN/Fs
R8aZhuhk/+RnsQrnTOMBE/3mlV/6Vr4ExvC3to4fMc4CVPis49k/NCcryEDtUeia
kw8zev2mtODBXsR9SII50CLpLWzF/K8kXhlJcfOcRj6F4WsgQiWH9MHlGWzgFq0A
G4gFq/uIlXnPptWQv3TriYNC1+dMpYK+EXp8oERcfX4Fp4ZhO1ucKckhbMLTcOoB
YynVSLDhWrOo54IrkCRxugsK0JprJwhmVhYALTa1k8mbYUEvPbMYVvP3ckYhoLEz
bEmwLuPpVPKOdSC81IPkPDxahrjD1U1rkpaQv3P5tlj+CFFPzriiHLS9YrjIZmnx
myQFh/SbtcLyCgrUdr7EOZZ2qRcY/lu4kUHL113mnEuzf7g+BM7vj1tXMseLttJe
P7Z2IO+OUeCwI0qlYZgnwvV5RgK9SJaQzFihXwA3gxpqPAMVqSSb3bdwCr2GYA6K
l0A1cr/IDRB3yq0dHWmpHsKdgae60rC08azLo8WsaPPZwRfYgZQA7p5W2ucMwQY6
hQ2ldqFcmg2rB4QmWGVE173ZfoLnrwf9yTsEvyBAKgHQimFbMvuvDGZhtK9JWMiZ
G1L8PVvuoZ+WuM5FQigs0BCWexu22fZO0ugrwo4YBO/SL8yw2DiC5tVq2jCIDYFe
TKXdLSmQh5cgdR+8OB/hUXJbZI/TLRR8d6NTpcC18Z4JudbDloE+2p4k91pKng0t
+/O9ZZq59+BqwDOjNqFh+gu4GUfhh66LiSKD3jp2S6qCJyrmLdDPnj/UNijL3NAE
kcdzZ7bnn5IQ6ZaGjlTAIMp/WgxHzdpK+ABAKz+PVm4wFV71PWf3oiSyhvcXAjZm
AD2OHTu8cKt8z+EXWKfXG8nOuS90n9hhe/ljzuDsH0RgtU1PBlvY6EfsC7X24Wsz
Gb9+NwhMs0K9oxZxfxRZ+3jx1EjQfE4pvm6DnJ/S6A8guuJAtarfu0shCokPmJwb
AGKImhVzhL+4YKOQ/wCqUV06UM2Uqf+/u25ynaB3FRDqNK54Dt8MtTeMaw4DlFiO
SQDHWl8r7K3XoAvrnOxPHMtgPcZ97JYmw7hC59HWZ/SzmXuJNid11tuzL3ZGql69
TNtJ8ZpjEwWvivIYkHq3gQYxFlOlQCIIdUVlKhUP/7PxVtKbGgow4HNF0a7FB5mK
pVEZvu8qK5U4+FjhJyU4B/lF6U00/ulvZNBfl8aqKef8aor8Dm5ZeKfQjSFBUiuu
hL710ekgAprzrH7WhDTOryYfiwr4QvLbGCtE1Ur2sGniZCk5A8Ek1tD4pYYXRBl5
UADURlR2jjRytQcfmlbEUFu6G1y2RylOD/Dt9+jlsnTkm7fEXBCYOZTEfqBi0LHm
CtTDKLdUVMKkPNHas0QIJg2AEqmUgq/HhG90KVhoqSo9eNICfkQJ1qfLz4eAzRZi
G1Q+sCy2EIUFZFoLjx1EQN9AV3w/WtSZH85NktRk9pBDve5y2KnnTywpirffuJif
HOgNX1vD954azXQkvFOhoBpjnQnnPCl8S6+8ZrIGhJ0iwKa1WaTY/L93U7QPXuyx
E4SdFr51oWaNeDW6sXbflt7bxwpcn9WrKKhHeOqP6R5EqgWH1NyeA39FJb9hJ042
RS3Qx0y3soLS26wcGfLUUZd5ckkkQ3gfM1IWn8mXNiAWE/A9+FubrL+aBmYg6QpW
AUr1kzJczbjnEaIt+l1RnmUSmx70y+nIp0f1kUh4dPZX7v9t2cq37N8EL2DLQbHL
Bv6JtYSWRa/7L8+8iuoS2raeHTlwt8Y44Uj8LotrpYxfoSQN+eqShivoAIGvybBL
szF8iYRxdrwWX5sZNDGp6fvLY7HI0fwHQclHSJCnZkEhILdsIyyF2wexbfAI27mA
gdFLikxHNQz4UUi045xTM9MV0UdenlL4ylqIDeWLasMbU9oB6Dp0plv8AnSTPUyC
vYBVwf1qVGU6dnWcpd1CIi2EiG+NQi7OMcwcduZK7xL/CInIiyv4lOiRbzPaMB7V
vxpB9as2B1LOvs47oJedjkFj2xSJRJ96y0lhKhPzsuC1+m9TYuDUrL+p6zrZMH6D
LK6XhDnzFoxMoYERoYhq9SsnXPAIg4k0pvwj+hi2Y1ci417w+TsqG9yZX9lywU1k
QtSBSgNUoVvu2M/9Gm8e06gEAh/g9d+eismNA2p82WdRmf/JFqh9QtHxceSRqTxt
Mrf9ppsJt9wlRyQNRm/4faZwv3EBS/ApVNv3lPWEiFU+jOmF8vPU7OA600AJ3rFL
7LwlRmbxb+Zpbb1udxY5M+sRNJKcyllKMK/BfVBrfERi4PBDMrC2WDbY9iNiwY9o
nJ7Vzj6YsU1GvA4lYm2TSJU4AMRcteQ0bJsOnoQIPRuIQF8ijoSq8pqArGuio2Su
YwNZf28Pm9Zn+ikescic+HKhviZ6OhEsb/OUuCO6uNj/2OQCyxlHlKKZGOUwlyXx
5NRBxkuRa4VUaRZ6RUClfJdfZtGRF9pYABFZ3UgchLCcnsN296pJacxEkv+KvUg3
FMb03QVtZ8X8S7NkvZAtK/3RhgztT+hAH3svQIQn+C11kP2cB3Xy+CTZeAjMs24i
LZuMOnJEg0s/1z6R0tXo2rAIIpq8A8XVLAks9ybRONbu/vezQ4PwEHI5oNol2YBE
GyXyr0TxYbQ6Kl9WdzVf876KOcsUqjfieZXNbPzrSK1yH1EO0f6ruo0MKU30NEbM
ycPcI2uoo+vPSIGse9v+WPG+oIS/uEmAnVkNsZghij3V0XhQ7Sc9YNsSkT9+/B+e
AfKlr+BmL8wKgx4EpweHgixJHznQLnw3wMp/PHErqpCNUmkKuRWKFzp68IYc8/Jn
+PzvMKGCZi9qC2ERFzP8xr5bzkIS9C/AnG7Eh4+PbhCDt4q3t0f3xqq/ZU6D+2V/
cPMLIUE04hYRcUMnZAFsH1YxisCQKyTIQFb8a+5vRS7UGt6R8JnkUu0xUEVt5mN6
b4Juni+6QWQdUDvhIHotWyG5Pg3tlIbEE1XORo1Fd3GrXWeMWkW0ZJTJpwi9ikXK
HZUZc+ddB1O3iouqrzx5MYaRhp8hDjZVOrqYug9N81ZR0CR2f4qrcmiJwHXKqbxb
d/7BRB/SuCLoNah4AwFKQsKUu+jtk9Xh+ii9fPX7b/kTdJBF8mDLg6M+yKF7LcYH
5KGrTEligXTuTjcToZ2LP3O+r8rQkllWDK+5GmaXf963Z3YRPunQfQnRmhWkqz32
LjbK7puHUkSUcypDknZ+Rr/lHTz6Kc4AeJFYywRIhDDCMNlK/q99G7yBndcEIMx4
Y/q+Rtk67yxG0HyL6Gcq0yrgMJa7wuWh/pCGhK33lvZaDQFhahqh71fYy0Nify6U
xg42M1os9lLMEkycCyj1Ga8ZOhYHv8eq2iVJNjej3iDJDm/5bcFEFAmMn1uvcZNL
X3cEyYHs3SEtZ21VHkyZc6sZFcTAtpX9mYfZRd44R8OoO5ASqRm0W2gxyh/NqTzx
y+QPtR0JP5bvDS+inSQ2khgSU6xyOSCJzXkrIsuusFuM3JcKGfW8LfSkrHtMbRrT
ni45laErQGzp1kA2h1RDaZIEsuej86e+0/ueT/gk43wQNoi1PWhlK3pM2oOOK9uJ
o6fKYC5iZ5ni1hUGVBKZXpl02OKl1KZxmkCIy4Rm/bNXPKqpkqUrTgPMMx68kdw2
fagY7q1xqzq4On3Hi73GV1W7YV9Tg4gkaq41soj/KcJBFyBjXeq6xvtclcBB1mga
2NVqvbGtKGXAZOtYgPRcl1uv5IZuzmlXtMu9mdl4DsEv9PRodCOjwGg+fQ6iaCzs
V+c/K8oEmcy7Uzdk65uG/2+RSg7tJSzgthyY6+L/Abkm6dMQAbvqm2VxKerl30re
cI05yKP7VHTHZrSHFvC1MlaSayToqa+Yb6wSBmVix4OnmBPCztGZFLqqscYrcAof
0Gz8DO/3W+Ft3qJIYXiHDSsgOIxygdkQuyhG1IqLalBiEORUCcIFV6tnvNpoRju7
TYAlCNOKBzjT/obdLL1JbFmzXv11n+j+8NKhqCEwgzgRVuI3MIJ9AAYQtr1tuGt9
xBon0DidCySCXvRUhZozdq5YhFXg3SqyjmD9X2MSBOJG9waH1OY4HKeZxFq6kQ47
KDsVaOWOjV5yWH7wl7hvut09RqshdA3qJYAfILeh9AmzRUEITtddWD+hFp/foEKG
PMqmzE+IGfkeKxUVaQqZ95TuJG+EWpw6g7VVk9SNLHdZk0MpXQmoIw52THmF0hWG
VDsZ9r6i4A36wXYKgEqDXX/K1jBWdYZGOmQA75PecEmYWn+2ZpOTkioM3wjiOqLW
iHLxviJDziOCsz9hGum1w/phht5N3EQCDHbu1jL8M+G3wuuyUZuOxWA9a9G3+fUG
lsW0C2Q8dXlx7fwqz7UnF3R/dYHT2LxBBemoxUxrTRlVHnZpWdUf631NZFn3IbVT
yS5XIasvwotHWUKCL6nnAmhoY78sQowHcgshTwNO9W/MPiVKupufkX57XocTPgwb
v0rRhkBT8Oa/K/+dpRvJLGnb1TMHkIMdd5emmbbOrnkgszmQDHGK6ei3NOzefcpd
J+2ZdXEydO8tXEllmCVETMSU038SWQlkAX4dodM4A1O1dpdG0/MIxjtAdNQe9/q/
/RhUAi+6HdKXKFEIBRkeS1fSTxDnXYAlQoYu+iHkEMdRQxM/jSKf3dRPGtJSIAUr
F9OBFe7siTrj70TfKw2pHZVxkq+apfe1zNauAqPF0Ker0FDYcJZOkX0i8508m6i5
cWLhoU6AM5M72MwHaqc70wvxFFBToIs4+ya2bqr1i737nabV0V+rLtpunBxs0URS
jWckAXz0UErP6pRzb+jT8JaoWyHXb3G3angYD0UJVXVeXboCxT0AtdqPdZBsgXn7
bafLSIVZP7FZsM+jjjLPsmYOpE7DpLsnFzXPoRDgojimn3ylKiffMUcysqV7Dac7
DtKD7Od4FiBh35X7DAn0yiW4e9JqKp9Vu8zgALmpPbj7nLCNJSrHoGE3FX1JOGS9
2AyOd7LwRA6DNoyAps08s2HE4F/E54zo4M1HS6qFNOpLyo0GTvMVx/NlPvshUkyY
YR79nfq13k6GnM4KuVhNhVdJA3Q8Movk31pYtoNaczJcCSdi9sAOas3uMIBCjYJd
UYJzQPk1re2XWpKByl5uSVszNBQpAx1aFHcNmjbYeaMU2glce9LydR6+5sOrw1CY
VBk6SYDVS0/mFRYkT/gkH2dFS5dCH8OCeOuNG2mtTAKCgdx0ik7/Y3OsaRuhjELL
GygJ1Q+bD+nkCN34HAmj3WNSpkdW30ef0/GPsgDli5rqh8zTdIvhj+AG2Ux4FcvS
AJKPBTS8bQIh2u4tTLKsdBQlEs1W4drDzOoBwiMn9KZTYfDJxiZqmZYAkFOkKe/4
+xZG7X0wLjwBwYRzn+m7vmqEWlcjfiR4DKK2eCPh4PeIR9XJM7zmCeGcZ/7PIjt7
zkppia3EuytH69tyGRF1TUAHfC/M2KYPMk1/TA/NuTZLQ8D+VsqP80zDs04n/jJ1
rlXyb0HPTUIX0qNvSzONYOosBmTxWt9/el6Vd2E6Yv4zZic7iYDaNRrJLOAK0qj2
0RMJtD2bfaEIx8otkc7jSW1x4rnksG4k6Mk22w9shXX0B62LmZegO8vP1PO2txfO
6pd5iWNTR64Mc+VC8H4Rk1rt/m6FVdDp6SWBPW6l0mAM2eIS36PeQjapV4pI6Bqe
HNoqsLMnFJ9xlTRDu8TrLSBVDyO3UdhSCo1m8IIA9HQMTjTPkuOz42SRwX0jl9+A
Xsl7XBAGT8VKc6KTHIGOu9zpIN45xcf+aAB+TO7NL3zJ2B93Gw+xC2CBdQ3yeU1H
/A1yWIaIJvLrhDvE2ZFYr/7L6US1C0RM7OrgN9s+E9tin8hS8yHyGPSPLy9hqYFy
P4x1QRM7SHkGJ/jQQ5+C2ZlKH+g3QNQbXDySKOfzdlSBgo6YoSmFUrbgDQQFkjB6
MtqvH+f67fIo9F2InsUKNp0844uI7HdShx0nZMzlb9nkzDnm07QbT7qioaRPwF/w
zRwJ+YvW10SRgl5oGH/sEECk9CqhyXAhb1p1fHo4mNQcIiQrLnZqtcqXMlZf6/tn
4CHvzAW8OqSnVGE1XDXVWLNDRcMG6YvPZMFleQQbqvNCTej16RvcM4+ChohPN11T
DDLQ824OCOoVR5OhLas+1zORYqjR+lmGa8TRJN6na1AyI1xeHo6oV57+kmgUFZ1/
R9ulwlFgXMiYi3Ff0FJHSeMkozlT8g+RorMXNT686el0YjUegWQClFXbBBZmivY5
05TzjNhC7GCYFQlmArU9ugPq/L6tMWtp1z9PDkNln4IaaDW/yu2FPxzBaA54cVdG
CTekQZj8PC+0rA/ItWYbfflMkf23+Kq6Ks3N5fGbdDbVHexWMUMyh8WdRBFoahyf
ta0vwv2DWSEvtDHJh2bqng4MEuBrPUe5mWPcgirGPuttDkahOrF9LMSDnfnZVa24
WXy8eTvQ8UJCitdeng3Nknv2zivBzupl1DUAxbzHjPY5VTmlgDPLfYDqDwJU7CBQ
xUPBIIksKf7/EDNYL/4876QqFYaOTvv5nGHJYtCAnwuRiT6VAw6Fk3iPznL4Px/s
wXOhHF9/zJdbZtfXcAS1QYEOpTgrHuOBS6OnKy4T9SqNq4jWT85PH3Lve5UwfJBl
MyMSce+lO7O1md/1I6r5YduQoDCK2IkcC6dSJiQGTaT+RxGwXLbooVW9OZjS1UT+
fKhIjAwo2lCsDpqROPeNxsnpEIijfVASdwJ9blsZni/faoPU3XTvDc8mPj+2p7SK
ZJC0M2izzTM69TXT4WAhh9zOTOKc++VX1++DpSCSqoeP2c4UWHdOgaXzdSNAXw9m
ENfnfjvXzadehVSeWsUacpDE8ihmdMpNYL2S7rKGRI+eMa4hQd8k/3XRzYR3Ec5S
qozWOWEp+hz3CLCjyR9zL/jg4dHSpVy8mjZ3W/LiyX1CCzCZTQyIAiQXeKGv+MTR
4wy8WlREfmm+MAb7c2SaNHUhWZ68iE+iVjWQPQ1U+98Y/07O6oh9FE3njbATGXj1
BaFWCyFUbYuy2lloNn8aLkoS54LjvFV2h+SqZwjJTwwuhAhmvMinQLu1wXv6D2K9
PNuPlU5rs0LDFYBu1djbw8pswVKVenCFh1kB0QnFxA2ErbeTVvDHWO89gOk+s/Tj
+kEOeilky6C0RXqltjfqt4CuTwCzAizU+rRh9+PBMCXAjVBlzRaPg93jpMvkAb/2
iQjR2fnErRlYvy1w4j0VYlNFzBSkqyDfysJS3USYOujR/yDMZ/syd96etaOK7mb5
PkHSlqJD78KjYGKN43Kvgs8iZCznCJYWZPvAEMwME2PUxvE0Tfitq+I8F5ycSB/Y
RV4ayMli/ZtWayAZSqh+/RzF5BW9Td5fT0KfVeun3T1tmsGPFPzSePQrurCEYX7Q
He0g2BMfDMhvI0ZOF1F+bVLtSr8XoUdhH4kr28BcZgVvkkjf2bmYB5gD1agK7342
n2Yhv+UQhJWyc+fEmEJ179n4VnBTneVKXyKj8dJIvHQADJXF7ggAL2Sj5NMGZw3c
iU9dpWaSjiHtRUStVZ9oa6S/oBO4FETOau1cSDNMruwj8S0qvXnBE9XADxdqRdgG
nC5e/an3i+ZNK9P1f8sxy6XZ51NAw1kU8rr7r0kg40DTpPJ0dtdFfHf3Me+rJaG4
limcZ1tdW1lLFBkwIoWTd59bs3vORK1DEJ6YxjogrdGiiVY8Ffsby3c3g9s1plmI
RE8mXY7vO7k0TrsmC8tc8tE2YBjX5PSiOiU26T5fPpEdLQrDo3BeoT4Q/REq93Wg
jtni8JtyRzlqhuOfo/4pmdn/CWXOynTqMDhRGkhY+JVm9eFJnznU80+lqNXZkVlk
8aMpn7TIxSdul+Sy7rI4Rai1jl1aeOVKei0mPZ87G3gVr3Jh/0TLT6IjLe8RLWrh
+HrSsl8+LkfihtN1M6tu/jmF0QFhGqM6FVKttyqrD+qE45pt7uHSptvqzG+G9jJb
g+7kS+SjO4vYDwQh8pEHq1RGtsovT94NvGfoDLf3SXV1u5KfBvcDlfj0uhmY1ooV
RjrPpq/VKPBA4U78AMB0q05IGKBrvUjyz/LgTUJT+SgNAjoXHdxpF23vZdBtFrMS
xBGWfwj16pSQUCbgaXyrg4T0vZ9mYd+Ac8B3WQq80GsrDFBprSWLeROMgpk25cCG
72m32Jb62GG875L7PIUYjcbQPv9cVBl+oJ3QrBzk5LU5ecU3NQMfkREMKKTCFYB8
dfQopxAFkJATBDXtDyMsOuvqNexYbN0qstkK7yDmjGpGZmM5uQ+g8JQ1o1Yql9wt
Wub9heTyapzPydFEGkMhfJ9i3rnEKVOECiutajW7z+POrKrxPetaBURS6/gQKzco
5GO5B7QcdNjFF9osv3eeTMR2/athYAD3q3PW0ZnfP76X6GGNlwakx64lHVobZkJC
ISaalPAXh4Oi3vcce2sXwHkhTArbRSky4Qx7tsRWxjrxdGW4HQHh5SIwbD/9KRjZ
aIYsPcU4lZueijqtJSZ1E6r8RDrtKLYP4Cp0KgsX7O9U8Sv2MqggOlz09ZTVOuYP
i/5xpg6+/1ZmnnrQnA6T6ysUZWwea3bkXAVhWVggwM3h0Izv56F7quIE3p7/0wFV
/pQBKT/FAAkYNHEE3rbkhiaLhQogXAMc/RP5GowuJIQ0eV8V91+lV2joazUAHyXn
sxchuUcl64awsf/aSb+K2ufL7IL9ecN5m1BZWCv7qHptS7O4i70rCIfr7HcOu2Si
PAU91zsJAm8y8AELSQUTAS64tFhAHBRLsvxcTeXB852TMdmBwwwia4mrHoQwVt4A
GfqtI/e3xuF7If1cUx/kwDblrOLmL1gE6TVPxb0EDNsvD0ovBtH8OBYa9kDSzBzr
opa4Wzwf9UFN7CT9TY+eVkNbbe/cktDLKXwsoMMPaaPUdjtKOEylu3+J+0sqMCkY
RmVaV/RhI/5KoTCGe9+D3ivS24t29rMY7kTEY9W+2hmTnXQl+RNnIvl2lHujg4Xc
P/iawa9Gqys8Htm2NnziNhqmguNHUnst+aMUseHYW9fwDiOkLH91Jrf5xFshf4cZ
Qq9CwDkh7I4qiaeshjaNEODeEzD7NNuPk3gfu+SqZ7R5DnQfPFoNLAuivMxiGY9P
fdfMbskbTXRGSjJeuHc1SUIr8JeTsJysHBqHQc9Mc51T4q0GoQckKFanr7xjkAok
Bq6+iCDqIg5bPBZCGbSdZUQ/LlxLdJ3g9FC7+WxGXIingLQ/oN9T4N+vD81I+Ksy
9QqqeZtzOIe18PRiqLhBOVLiTVVBS32kPOpQ2qbWop3TZN6nzDdmtIJmuttknqHr
+LuXbT3unoRgDu6uV63RAzVcQJ+LSpChBltYlQ72oMbyuvHNQpFBLQUoWgn1jf11
CXl2sf+mwPZ3TAu3ZD2gjZ0u13A+dyX0tPV31oGN+Y2t0Tj9SpZmORKOBjsxiRHz
Gcz/mpIL8hDPisoXHG8Z5Tu0f09i2unpkr1ZzbqOPLC3mVfYYwJCZxiyfoV1iYjU
5ter1jTjU4Yf3EJF/hfC2po79GAUbxekuVW2i0wS6WN+eVHAHsPSnl937DmoXi5E
v1SxZR9nADSupekTVGcv+/IQRDvCL6lrKilpzobVvsI7DLiZBQtuZnYYJmkWgjCO
+SoKnIeIwSDAZzt+oBaf5KzNj9zd2bpRqaiIiyzSzHZRheFUWlhiWcP5QjlBW8OX
B2f9pRFiXGOUqvoXufNZTRihPjj0Hq7J8huAScrXviYw8qK6vnv9D0PWn4P7NGyk
mrydVzQ9M/qpmwj7dEGb+tBINK5txNv+9a8ggmOUURt6+H7lRyaxWNEYnW7yZSoF
dOyNxfF+gEY3LCxgihg0XJi1n8yGovErL28X96UAHrCvDM73jf/36g4uVPHXHnPx
jJrvH+TDlb8fw2+VSYqqHsp4p0UJ4GbyDz14X38LcImS3cljHgGmT4/3YpU6KCDM
AU/LZbze6YH064L67V2j4Zt8UuTvmwl2Pkq4v31jG6F4761kgUAaab3PORPs26Je
sQN67UTnfbnrAKZB/dXMmteWfWsrBgiiiJl5MErU1McQEYqIWryvnPOrNxzK/3rw
o5gDbqKSD2RZ3tIhuZWEmnXXklzhV90dNpLsudvXmv96nLXBL3/3FGyb5tUqEzta
Y7ulRpFs4nQxvbC+/4uXnszvdC7diBmQfs0qwyoMx3lIKX9XSykGc9IfDWV8SOqJ
Bie9DDAOkw0FC/Yq9ypx9AkUzSSHJNi9YHuoLzBwgXVqnT63lZvAdATcdx/uQsHD
vel1cYEMVvKskuda6a66/D8g7pu145DdN2I5Vy/e2XrA5uaX9L7zT3wFYB7X8CtS
85poRsnhYaMKe8NdEi1y7JHjPfTwkR8G36qClZhoW8w7qvlY56LrUdnZgoMcEdkL
M0EM2ePaiID71TAMj5O57toZIC0j0kCZP4R7BG7UWxsdxuFpyMICBy6HoDch/cDU
jyty8pgJyLxQJU9PWB2V+z4qMgy/zR0dp6u+GHp9zAydCKQOGLohU1Cp5fJzsQtN
fwj9T46DiUP4QcjFeljsi8bY6XlYauezvXUKtttYrqfJHkYcdM2UF47PToVQWd9m
Ith/hYE9Z55q1jgQiLkpIXPwFqOdqD28KTXcmFz3HG9skH3rZl81+FgN36Pfme6Z
1uvxVLi1KYxmCmLjb1zwXbanK+H2KL9FuwvkvtL4wvGVXs12odV+CKPZsYMSyYfQ
C50mjf8S/JvmGfQBfKNup8Zwbh0jYjzfWrIyXFit6We4mKF8xalTjLNykAJDeug7
K/WFfp8dfmoDFR70JflQ/0M21lM+BFoXriDVEciFDJMs/IOkvKzyKNVCwpGPpmHZ
tvP9Ky1zhvWIS3ATGFEdYDKGrd+D+77NPWIBu/NEuhisQ0Zm/FWsSdGK1ciStBLT
7KfZbtEQph5eCUS/W4TaFRtpX1dG82vZ4/C1R1weEEvn/GEpACdM+LTmNkSWOcmc
mXStdDp0a5tI4InBesub3wiJbsdg6+V5E7yzAa75oZz2kU8+4RsjstBKr7P/aO5A
rd2+EcLkD882Lx6R2f11Q65TzxbXObUWPRBPo/a5wlBKrF4Kw8itYuLcuGuCCLQu
RHyelfNUf2RLsMhDVHhGp7f/r6pP+snbUmEXqeZTfc75wQLpjpbLZbml5r7yBQKJ
1BUMNFT7MGWFdR07F4Hc7rCpqSWzoQYcIItw/yGFyJ8ec77OcFL7oJHUG/WZKic7
PU0puWNsNoIEgSmKz7Uu8zz+H6gLIPWgJyrkn04wNhlQJZSorGMmoFAb6dwiG2I9
Vlq9IhjmfM7+YpzT52VuCG4y5pmNe43tihCDdvZb4q52ebsI1Exf7s5ZTRCltrJE
SIFhzBRXZ9V/Xovj+c5yQIyw6QNu3UbH2CX/zQqcGlZJreAb/vABeMOdV7i+hGy8
uLPWQwFMOOmx4w+4D/uflmjqWW2X6iHgRBEhYPC6BCLcpFK8x3sIH7y3N7UAlxFr
nOPY8pItx3WtFZdf4dCcEMhjUtpVVAmZ8C8XDZBeYWSQ60nbe3zLBvxtC0nPV66r
QB74fWOeZDODfE4vGyq9Y8XPy2j9XSdz5B6E59I+iUg/50LZyZVYCOu03z9hN0Jw
df3nCV76pG88ZlW2W/tv5l6Z/mHXvJVLro/ARd61KeTAYHnQLNyKwazqs1jCO57c
LCxlCXCoRwnsjqwLOXhu88JRcbBJ66/xZyjCRfHuXpmdsi1kTD15HVuMktDKBTFJ
vh9x2sjIoEAkc2tO052DwMUw4pQDEKYeNe8nYMBiQVMDOn+IwHeBgiJJTxPKxWLv
k08fQ837V+SKXsdQLbY23pz+5FQLtCUIGlpesLdHfJkvr3Q5FD7kb7MS8IINOGnk
pxMKqq2GZuF9r6QySy8QQkvBsoCp8pqLz0lce/OxopwRftC1yzsCnF/823bemUms
vheFRHSgSw4mREhZIH4PIJuXzJvyyA2Ly1IxMTY+PNokYieM2Cq4IULeqTHFSVBb
LsYKLY0W7V+IUHTJYlM1SXk5XyRpumoi6wf/IGtO4N/KrZTnLRNDhmxYXJhv3uWv
rYSk41JRGFe5l+urvjeuqZ4ZNxtJxjB3zcFEQXrioq7834MQF0+pupDIozr0EJw6
Ql6dPKbnVBikPfm6URKxmrCYuMRUdSn2Y00ZYaRSVlg1QiaFl+70TNT4ATIUmxO6
0WBrpqPSK1m+3bIJ6c17YLqEYCT2HIi1Pdy+PtOPo/cEHKL+U2nCyrIZMcGt68ea
D7Bo/gNUOX6pmM2P7a6jDOKqfukpQBLXuxkDOjxXqfgw59mk/Q4gQAraf6+sO0qY
Iz6N41wNwZsK0MD5oe1xJMP33pjQS/OeSouGKw/WY1iI+cGC5I0Px9rJlHQSQhIC
GuqtdI4bMYpACD4uHF7ut2AZYmgGoRIlV5zMUfcFIaZJv3Samg1Dc17EFHUIeK3V
N2aRyWOeJZ/gW2ikXnQj+vpi9Nx40XKy0t4SRL66BqOVZ2IKZaZnk7W23Df50Zvp
ljAyt0SXLYWlClXQvcl34ahMmA9qLsu+nNyVAl4lpGWmbwPwLStCPFXiCcFkrEiF
WO4PUT/ZvJmB9qcCS+RHKIGz4WQnzWmC0roL1FXlJ5bwE1JjNMAZuBFu7oiuSOTa
kZpDs5lGzyI7aZnt+ni5pouJsdPuFSS+C/WUK7X5nnDqLEzFC3lUh8D0QKd1sbVE
PhELFi9TmTwuT1UVpSoOBJPO6wpwCxSXGj4TzLxrXQfv4pMQ35MMS24ilIRzuuZ4
GhdgvcQbB0dhhgzR+V83BnF6F9kZDTqKY70O6oUOke/dSvoofQDcAHRpp/vKWem2
fhwGzPuFhDXE2Tu/J+D6Ef7F7b1gG7C2dQVQAL3ocquWdmk7iCHKzX5fR2Q4pXol
W60HM36Fpbnz89AEk7GIeDZC7Japo+M9HVOBJKxNnlOFEV1d6AWveMIN1MKIeL8T
E6WGbh7lKAKH3ohlQY0VeM/YVtFUgUsivOW+OtnrIWKaM+tbZv+TowZUsKpIOXTC
b2n+tVi6rHiX+us0UZbvGw/y9s3puQLYrQGnJJhudvGQTZMxNEaWOofU+isrG3f/
ERwvqASs0Fd8UQjn2Lb3iUS2O7iYo0hRbzoQ1Q4v21tRqrwXQbFsRgpiyLsbBRXV
tI8pDbT8BpN3ll1HmfScQWvUBFofQsrwJrT6Fd82fgGiiXzjIXQv7h7fAi1YVprP
Np4rBzZMcTNn3Xz9IYtm1/HuD6BIGHSYORaGFhg34ewcIxrIfmRtgBKu7jm/+Dl5
UtpNAghLMiXltt/MvHAbMGA5eLWKy0ByHTkxSucjv/oVCyAVPbKorrv/VONG5Z9q
z+6UuTBsl4G9aFxS01Ek+nQsNf2JuMLbF9ZhgUZ+2JABkrT5exOhgwTsqx73jzUl
4pEL2/UW+zBHmAt2gW9z7gH8VMAFGiqL+4ybgJpYaCQrqbPmtjE6LE1cibmM6te9
zaiO/rvYrfFMge+pw99V2E91VClFaVyfkMocHqbn1AFA36Y5JN3SirtXmW7X0RHP
1uXdCpB1LDDJKat/YMJwe7nVsh2iQ9Bg2ROcO6476wuew4Lx3cEztbILbRN6KU3f
mwdlObERl4ILev0v3YmiNA3Tg8Qr1gjL6ZeBB4ab7VKUHfzCCpdJa0sKoARuf83Q
9tWuraURMBDagOg+4RmWaEQNf185+yw0BVS3vwchPQEbo8TkZlm0/eELeuTBTTCW
L8+FskEzMH7tZM1/tN4FkUh09uV9/fOkDOv666NCaJ1RUdbg3sneClDCJWQUPvsv
gsg+XVx9AvHEpeEBPH0g8t0EtVd/bl/03oWy8l4c0kwjReJY8Aj36V/GJobsk0Ey
jXTjmrlZslrdcGhuCngi0ncri8iLldYv6PsH4mXktcgNWsKdGXnVu9YB5pB/U4r6
xlWM42CWWs+cbhRw1raCQfpE/bPaF3dLOS3KlSkOrhP5D/pRcUsLTnHGzINnibPJ
8v71+1pyjFix/grKRkwRrTXz0orKgJSUOSlOnY8hVsgWJ0ZQhm0g6T/mK3UNPm/I
jhsK0Ou432deqvi0SzfWa3GlNdvTPmUceBEQ36kwouUC+RQP0YLDLRcvWLXVo/8A
RcyeWAeyuATmrEes6u7m1RbifWeptBrAwPdD0Fht9Wo7dq6zAAfTU2I/nc8tmF9c
S5bctQUTqPmfWsSGzUsB+0ArWw2Uhn3B98CpiGz6mHOYe/lSEjCD5F1Z93EDDimk
62ZMgwsuISjknZKmADR3qlMTjvvXyfWhdm2giBNa6rnR8Elb+7Yk2/5+l9oWMWXK
qm0NK4l2RoX5d4VXXexg7tT4iLKhRfBjeorplWl9/duNb/N93FB+9CxrwJyAiHRG
WfOxOdlM+B4KhOQorfJ4IP3gSdheKB6jf1bJqv4efgEn9RGqbnUaSP5gyWJWk1m3
zKrjBoy/an/pzjoeYF4pis/anobXtGZqADXaKkp/4qA+Ng0dpcIZkohOQFShcyGx
B8u4z6Bz6/m9A3oliTP4JaEdiSSoya3FBrsZt4zI75HM5BqHJb414D0KPoklCDVo
vEsUgFlftIw/MDsx1h0LTgiF29iZ3z7fnlfhKKUH+Mq3EVXZRJTgnZl2xZiCtPzh
w4d3/gEEEDTn/BpUveAT2c4ZhTRPyw+BOE5vF9ou1plzSXjPAzOFCLwLg0LK7LkX
2D/nYID/piZtXreHYnLXssPEKf0osVDzmdgscZr6+MxS47fe2zGa+tB9q3aiNvNq
qOcdI1hgkcQ+g18/p4ClTaQ48HaNZV7CQrVrvkwus9eiUYhIxsyZesgHYJ9Vwc/E
UEj3QtR6wQIfZ4LJWSo6IMHJBLbtXmsHzGkbH2b32lQC3hXEfI9fKpZwQsz7lxZD
elc/b8VCVb0oW2BwOb88AaVQHLw82dmDB6fpuePZbTpqOLQpDnMKhxkolIDmIGdg
9IdSBddWlnHv5pT4eb/qOSWx9+m//NEnqbZIQKO6iEOIemoopcuucm4lGdQ+oIHi
q/FkQ1lKfDbe58IiymgoMstgpZ2leWqAVTvTzh5JFCXkEBedQIHozWb5xWMusN/Z
hKCWj7VdpCTw8FiJZZtO3okJTmOn6wf+u+9/j2psOnUPJDX84Y9IK2TrYojP/F0n
XeDEMFBgxkZ6DFSKyppvc36v2W0+hrR2YgP6lu2kxxn5z0HQGVHMC9+D5VbqyOkC
9J/L2kWTYcaaowx0AV5bh/6bu4qKkZcxJe4Iaw54mBGCXIlIUU4VEBMiS2fWTdnL
sJYn0idkW8/bzz5QirRut8S6qAOZ7QRrY+ksqMDt0mrzfc9NW27jrHWrfkiuTZ0o
yX8UDkvHzjwv/ATYEGxUtRXEv3CO46SjhV/HnTnvmN0Zf3DqI4M5HGEBE8ClTk1r
bAGp916jkzrHyV9mdH1AQ4GERaYVAFLCL2S0FSsDU3F8ve0oX4zcMfaDxraikV5a
ZgE70nC64thSbOttt3poMPEnQwtAZuGydcOp389M8VB1um4Xuv0AUzDXEOm4+525
h88HNvfodICzuO+Hde1+J4/nyhjh9oqrr5+pkoRb+PQr8/g1QPZPjMa+yGW9CyrM
bLL7XjHla+46bgr06YYNKEylOTJUkZfSrT3j2yojixJFXPSaNE/qNZ5Ep9o0kG9d
6ZYRtL6VSIFzq3Hztb0sB6zyQqpROjZFgrVTw8nUV+8uBkRad66eNM/tdEnYPjMG
8p/4HDC9NsPAnVb/FX4g8Q+LAcryhUd00RfTS+cxYoCZMoaHFSE+djPjK5TaVKF0
9XQOku/kgGYFEoDUv+N1dWcAr+sbvjzJTvztJoPLFfVXHwBRixmSk0l+VDtnlEY2
7d8lk8pjtqE5Ym/0TjCaQXy52qqVrxXxwJ98g65aM/Dk9XMYQgl0vPVxB1nxQt6Z
V+0PtaboBdQXnQcm89piAa453XvwbAMKoOmKF9GPlx4Ad/2Z17syMX1oeTKi+nrB
KG3i3T6cW26/GyESsR9Kd9wSAGn4gxCc79lcO0+AbglbF07DVnddurKGu9golpck
kDMCDjHPXQn8g0nRo3b3/8hgCKX9G/r/fmp525UWqBAraeePalaKdfcUySmuVpxC
HSRyHD18uM3kxYZEaeWPMlgGD9J2qHi1lNw5y2+jNU/GrWBriyQCtLTzvCToNcth
NzEIWQ87mkr9E2AXnUg40CivYWSsGN7C3Uj/a2U8CYTDLsZdtIhk6XAxq7Jdq8i/
SpVrlFl17z7W87N0Sp8FdeZ5M9JeMhzarK5sFeM/Y2SE4SHvtmPXTtPagwmmV9Js
D/bwjmJ8LeCacJtqNZetYi9gjRcoE2sabyS05BhwQph6vS2DFelbr4Uxjpm6Jywi
eP260+MIcW+L2VZo9FE4ANYvDTcw53Nx8jbeEI5L1FCdSwacrjUERt9QUd/FvDkF
uWPhL5f4L+1P1wlgF3m8FzPKenUD5MG09Un7xZT77F2MX72VTvKIyepJfAF3FYD3
wcisJdmxo3smbFGqGvNM4Bfzek+kWU4jyScKyUrWFUmMIXExXbgjdBjdsknUT0/O
ATfPrIjCBFZq/hvjj6SBNDt2yzXovZ7912MKgBa81L29wGRhp1/mfYmmhqkFYmKx
0xqWNJB7rLgMOAfAa2Ofw3m7+i/22GiTQPKUpBxqU5VnZRVam5ACdnCUPkSeY/5+
JR7YnJlDV01NIOdPMk4VdJKEP1QSjkCEZpTEGvMUXVz2j62UwX5fVXSKCrVS9olt
T2QNG3ahhg4e6nGMTyZTbxUmNR0KVhvBIxbkmuTmF81RU6xnref7NESXW3TLSvB5
4rJf3ivWMoh84mG+/wpdznrXTzwrZXt5eVLi1wxZ58L+9WrIA9RZ4I2uqpYy0lar
lKdjnQFJjgsbDOkjjpbPae4Y2h3PSnVrJmAvPGoAFhu3ecHEZI9IPgXFaBuowX3S
oGYDKlLnYm/zC36B72qLF0ABNk/XwiB3FjmNuJ9gTle0Ls0rAIQ34PHOc/K9exBU
r2Txs6kMuedP9xin+wPCoguhJXosJgUpyC02pwzbrlaehB3f9HTULc0cwNYoFp+W
wIQH+mhoWPP382hoQa/+280LcHozGmiSqGTa5y6RHGfxDWnCEKIWHFnl46DNwkPl
U4BbRcMU5i2oxO6fIuQxhE5xJIzKATNWZ8AvPWSvw0mEBlksj5o+kXuMuDlnskfw
wYgOpMMtvMth2VNBp7FYfHPcwhAwnpdZBQ7wLLifDvOOlDoPZnxGRuOii4PkSqHl
te05BhFZqkncrRwFylRkAf3OfUspPy7PqpMmYskAmzZL7WZTNZVKzlX1/Ys+WKZR
EW1b7fdvoXAPQZVVtrSfwBG/c5KEdx+zsoLe7+FxJVBQ94XMMR4M0ncx+tZ/Ei6C
LY7XuKcdAe9Rs+LDkqe0Fg+RfO06GTBNv++uYBgA3was7j/bXAlmpamG3DGz8CEx
D/N6XQ/wFAeEGqrKNAUWGSyZPmZ4L/u+dYxgLbke/xF715eo25/G5A6IC/K7Z5oB
/p47CRGkO/5sf1m7uWTdZZ97kRUwp/eTy//qc3pMXuoFHvatULyIIsCAHCVmPoTu
lOaa/qaXBHYn4y8SLWG0+GN9PcuVabNp0saKiFYzUtzDcBAZw7qgkfQ95bFwZSpZ
JbGbTwq/Q7txq6ffOI4Ee/nZWneZDEQuDKqTQkF1CuKrUsoNd5b6hQGq12MHjRDS
rN3cPMAIkaXOnMuyJHC4WSiZhx2k0DxXtwvQuk9ry016i0u4/vvYJYcumVZq3mxY
GpihY5GX1ZKpUwHiBtGx4sq84NfxqORhCUkLCWixE1CNda8qniyLQqFXHkYkDVgM
Q4i+tG3acAO7+s0mZt+ICm64ZDEvIqegbumBOkBspCrE7WxfKT1cUjcoaqksFIOH
H6xwGL2n0D004NJ4nv0O3tLmkUzCpUzX3+MZjzvE1l7WZTFiWn8uiLUJ7zcM1yn0
GjTWVmzEpdJRRFgXGNwIfY6AINxEWlJtCVrJsKpgdFf0OInXsCD1FTHt1pJ+/xxt
jEwOjDedruUzVaBOFzPFyyFPegrkBjnAB3FNpKXMH7YfjKzVjVAibfvCbyNN+RSG
DG6TcUqcBZGZlIDaN4jL+l6HyNlgc75Qv+Ud3f8QKqkLC7PWCxLdxy7eR/ZW/ukG
36Dm03D4woTHfrJ1lCj7BvuPqfzaEUTRt8wTpIQMaS4GVPOOuoptGvF/izGQ/LpF
y8ZJtYx8Mxk+uzPjNVy1oXnXchyC2TaxCNalN3nH3J1V7VhVJItw6lcsVzOqLr3C
k7nkwH5tdOjjJHBOsYCaOLIHo9HexiVw0Solydc1lnX5351O+aNFJzlAle3QVbmu
A346Wf/axcX+0W5FTw75cPKLQGVTv0n9xuD3AvTmRto519h/85swTH5I+JYPJibR
b0jA8xVUjaJkirqIwqBf9/9PVZmg1CFydO+6suLE4Q9HovueR+782NT++xFjjQWv
Kso9L/Dng/MZMERX3uu/XOKKJHkSwSorSTPTeaj5HRMUtKS3aOuhDYeALORHb28K
F8BJK0X+2JHDEttgDoVO+Sl9yMzXMnc5eHeUHkdA2NPcxX3McGdYw5Nq7lTiGujI
OIMr0AUVdQ3piE77lMAKZzWmp5Z/c1kLNKBGB3ALGOT0jzTwxAjYq8D7xfjRY6MC
kacHq8nNypcbqiJSZGVG8dOVNhdA72NlSbzJ65sIGgTwCbIzhEuBK81bcLS/SN+v
ftYQDyu+ygLzUUE38nqYhDYDWkExjhZMFT5zJJRfKzKf7u9YDIn3YZZcw4Fef23a
hvSbCOTsU2/tqe4E+Ssm6CD7UUrCQ1SnHkEP50uF1ffsJ2HCkbf1vYfIK8jspD5x
cjmPwFUAowc/hkH5uiu4WKnFt6S7z6iuiGUaVmBEBtoTk+pkZcsYdZzgDsl96nEq
bXWoo0QZAZr/4QDNk9xH27ybGYlYNjgQZWT8IxooIg9bNzZdeMn25F2VErqOli1P
UucRRmDfl2P+bZovQ7Pfn7aYr1RrvpwwdcFDpq4lw0cpyjlhsaYXWvronuNCZ5UC
nP4RaeYZdxP5n7fc+fBWxDu2+DycxrN/L8INFtvIi4JjladmbGGH4KXXKtxLQnKz
MUJKGMtdg9wFpm27pMi6QI88OaJaE/sog63EIVGYHru1lKCPAvPh1nnhs0sOW4ys
klLuTH9lF0fdzhPsNaPklhfT5bXk7fbkkZpdF3/bZwqr1v8DOgCsnPGtie4XAdbr
RhzkeL7eGq0WzgJuDqIWcN9rLKunNyNJhymetwsKP0uFWk/44OKyX12HhymJ7cIz
jl3zlW+3PjBTrX0wd4LEHY11vyGr0OXknOSKsyZ8Cktkm1LFcPmiXTS0OH8mfWMo
WxfJRaM8fFCh2XZ5tlrF9VZUlfhXp3DG0TiNip5N6V06TmwEjdfjK56EnaLGvYu3
e0dfs4qHNjAwI7zJa8lpCNmB6jw+J+y2y6ml1qG+irg2SgYBj82tMkg1oAHBPZEK
lkBZUqsJ7xqdFX0kKzCLd3HZE0dc7ZSKIgN3olis3Tw2eMNu7oEJ+yP3NunEFXVv
p5nXxqWyq3SLAQ3qLBAlVU9RwnFWBf9AcSfuMLOyQhiDJFk6EzrIWyVv/wIPhpjK
C1vQBsr+huKpqlKmYOYiry72GRvXiUult/ifNlPs/dU4ppIBrQ6mOZOZ/hfyeCGK
f4nsJ6zEkbTI2J2JR4GCFZivVKYFV9d2707wG3V4+8f+C/fyXh2CbTdNyJFGJ4Jw
VT+gbschQVjkMbgCfV14eLC1XIyWI5MLmxiLsGDMWmgvZcG/cRT/W3F66Jt1xuQ2
am0SOewXLA4imf87OAFPERD51XHNue3R4AeuBsJBgUhTxfLGRd8GL8THS5Qoa5y9
dwOKx2aTT55Ri7TSUViUEhxIVhmB5s6LRLJ1Av2R3aF+htciQk8/o0vaE7H4xaBI
+2zZ2BrQrc4RdPa50day8Bx11IyprrKcwhFjqcUITUrYAgd3tGfvNX7uJXaob4MW
Drvye+hTIHmYxaJHenYTe0lPumE46eLxkfhIksMJYYwo+rgQjeiX2ikUomTqEq+d
iupcSwyvvMJ45t3MD+fw3jAlTDKDGe0KjTfMYfOi2kMwIrRZ1HLPfuaIiSI1ba9U
raqUV3UyZlnfbK6mrv9Hq7YS/zdPkA/8NWDJWD6tUv7As0hHvColJ9Y4SwZGOJCu
s0fxEiN1VTk7GyCVqUFmEAIyc58sQConeL3tmyDKE+ff/8gm7GKJkpEBjj5Y7/VG
HBYNFaBdLf044W9K2PfXivN3gH8zoVdBsRM6gwcrPI47/GFUjkZFkP/tyVtT3FGW
RR/1kbXH5qMnOUtso0Am6uo8x2EfMemeogD/rnZxi+37KTWfm1j6ACDi393qtn2i
TgJrCLyF7MG/0CTnokd2IXWd8LRhxF8KDakamfuNRKATGt5HDm+hpnDRfHkeruY1
AInzEUWbiPXmk5FJoTtwBvW8PT0IsEfI/OW+ab8wSGk2Hw5FQfupD2TtbafrH02z
fclSg3Od6g1gv+A2c0YUcIw+x8sUEoevlcCneJsxfbMszPaq106SNLzHlSjjYflq
RbZAgAK7rUmEkn6CdsYYpmF9JJIwTgFMBo+AvKBHH5kqUjtNTwJttjgtxnTsBUVt
Qm7u9tg9Ws1vpvZFAiXSM9MD8XVA7u1Cf9PacnH+1NSvsuBf6psbw//CrTRCYxr8
ieGxgb0cZiwpDHNm8KbFU4QD6S948jPd861eesrthPSO2h9raI5tPbC4brzpjf7o
gY8eFgiB4D4ikd2HfqaSz/uOglF5dSOS/uf1CfF3V0onRRypQ9TWYY72BznvyOx4
Rio50xVBz1/5oP0pDKDBvl78ygzh8M/j9y220iqHdxDIz4DMGaID9D2bAJ2EPG4I
Ggzjym/mGuj0is+ujTWZHf6mkBrtDyK1Ayrj0DV4LNLJNY2sZn7qvVfb5QgGarCO
Qvg5H1Vb4eL7bKE/OdAN3eOTRnTL1O1n3oyp2EG15Sy0ICjfR7MsOndSWPUXpRU8
cVSpSK2vUutqDR1v7KdxU/utUtK8wOZkyNI8nCsxeeXm9mTnzUNOeSiw1xnL8of2
/PvDkCibATSJN1QDZRxvbKanPPQhH/4htRfVGesty3kV88CkgKnu7N9jenLB4Q/m
h4+sUXJIdbSuidlZkL5Ir8heJ1L1US0fICNkVMvOZ9Kb1ClZ/GAi9MjTkh8qjKzX
qbzvPAGWs77fAgJ2Wu1pn/nznGSvVn6p5SWQhClGiErcyfsr/3Ejsz2auL/WdomF
gzHuVhfTMrqSF0jgxQW1q7r5+/btgkKDcnieOLMbajHooI8uJIfIDPa/SDL+Q2sd
y8ia0q71PohKxvk+MBaaJFu1JRZizRcGns8HW9nISRqH8Jg0Y4b9Pjx1PNqNsPqI
tgreoVh0oK2OzUSZpdpXD5sgM+YHFSy41qSE12kAPaQ7a8hLpO5LhRc+jtVC02iu
9dHbErAlAmVQOAS1q9xWA5clZ/BcUSKMroVmTypyMps8gKnl8k1v4IqCY07i6vDE
m0SZuj3V5CVXtTUSUfLIwJODhwWzazfIC9nwUmt7N+eNA17+OzI96/ipZLxA2ZZ3
a8jCDeWi3SETN0wolSxfb3SH5j7E6nukc93cG9AApZcNnD+GLigZ2G3oxark2ka7
OK6HgFp9t0r0SNrF72VHEAyn29vGEwB1kmiN/2eBN7VRdudxtcB2Z+ESff2w2d34
L7ygUpEq/Ov+4HCxdTRHVWL9khwVt9Fip0JvzwAIvVvLM9UzflDrrTMY9eu5kl1s
ZHsGynyqZZrY2vlvbJ3IO/hnH78qUQ4rHsSXZzVS2E8ZgjzHhAtmgq7zAAVV5pV6
uqtT5jlbCFSiqjYVUqdKFORzK3hVIut2pM+2U39ZDh7Rl19QmO5RxydH2GEKcDpb
GzJaTwLGn6kcCb3uy0tUz1r++UBQpHXi6ZhHqwBudKVeXIbJ6iSgwsuWV7rly2z7
3WfituoiiUhzp8xBjVadj6wwhoQafYyBZj+PzCGr+g8xL8oCeF+dv26EVMxycfN5
pwt2NqVQW0HYvc70jEWE6gLIhuVqeptb+lY9zEN+uO8yC2cJIt6burGHR9kH1+jP
/2lRfPTy/5IGchxkxRGkf95ZlXviSRuwxjWlhhuM5i9zKMG/gdQGr7cqyme74+NO
i2yrjGdq6AkSXnxZfN6yDlkfNjqxhfp7CyyRHGeGq8WbNKRSvjirqkNI/od6P1nd
UAVYxtfbXehXP3zejvzvJ6qAsV+cN5bt8vQb6nt9neIG2BFBAWpW4Mf/zTCmID6j
TWcyMZdgD/i/V4mL58/22Wd79fKVZWObU4dYGTsR6fTyt3KLGkz3FxBj8JzcwZi2
XznvvTC6qamsnFinnv4bYY1f/ayo306Do01eY891e8rPEIM87sV5oXLqfuAXMHZH
KSJOoIjsNjEU7yhOD6HilCoV1EGZq0+qFZGYm8aSsZdlaTKpVG7PdtMyMAlpfM9B
JzvXnITBoX7LE69NzOxwuxXkWXwluDzT8JsiZJ6zNtw8Sh3uVwMJfCCElZa60Z+5
79QMXiwarLjF4iEzc+lbn6UZmeFR/NVp0SevLpJ+jDmGv5LBceoKfOettuCo17sm
AjpGHNWjd6jpYohSsOg7VAoV+QTCJczNiMEpDIBQECL97CsHq+VBURjgmVPQtOna
6cqqxayMS2X/ZR7Go5NzCWWga7BkQG8lqvlVO7EmKQrXRN/beiCy5/K/0ZMgzX4c
YOboeDkMbLPTHK1iakL82BhHJAt/JkNCbKxvG9NTGK+KTOp05EcPcX3L2lujEz3B
PQVldDrza+kOKelHgiCY8Fbi5P7RxQJi1Q5O0nuJSH3wMXjectAvNakLMUhtfeb0
J9o4XD01Mn0qEE1nrqkgRqWSC/M2FyMVRpQixzC9bgSLVMRE2k2aUO6aZwedv+yJ
UHsW8+Ecwk8LJCJQfWfmIzE9TTFGHZlWN8SsX5C6aAGb9DV749mVTpk9UKaxD8+v
R0fCZoXmhPQcxkdNPrFKcEkpZA0LZ3barR/CqbQ5b030nlmaPxDvv+3G6IprQw7c
96nL67r2SdrurphHCfKJ2AqqF+ayC7kBE6papjPcXZxFk6JanuvHARAsX9ncnYiO
bahmENL1tjn9ekjNQJr0qeJn8srybT+vxdv0W/S8qmQzUyrC+zMvshHvWJZXxbk0
EBk0+AkYZdmu++bI4X2oeqz7J0OU5pXdceltrv60f+du/0GcHZIOobTaXyN9l9jT
fHDm015kan9ZbZUMQ73b2PrrXjKwMj3Xd3GEx4S8X61lQC2ZujlnRS9tH/t0p+I3
h+f+nbyFriTd+IPv/8vgd3AzbkX3N/AXzHh7FObyL+HWjyS5l42n3Cet4rSObr4g
U4ddHrr1HRVG/mothI6r+ZlviRt2HwjkyXwLLSDazncihBLmjAdRAs879H5BYkGl
oEqR2C7iYsA8t6CEW/fo030QR2b6oy9SQySvrBD5+FdSH1Mewm8ezxBm5tTSj69r
scSyZKXxJlS7tsR0+t3YFT50D7SqHyQqH4YmZz68PVEubX3mLnUiiRQRyUBLTFAk
X74py6QLmWWb5QD7VjfpB3AlJhNZFoxdlLe3e6pGfmPICGCnpCqjstTZ5k5ghODm
cuRYXKXoU7J2omvmjPnovHhzD1SxTcehI1Dn7CopDTaZEzrxOdAdHpEN35QgORYW
38jo2HLANiYjKQuhCGedBe13QADew61LoUWqOBkVCUUGzmp+/feLzdJYu3rODLCX
L4jVC6CPJT7OjccY7uIdl9BRlDt0uX4PjOyL+wvDQaj/EU43+JsWPmP1xhSp1JCq
lpqnX2laFMF8rKjkemqbr6qiMnJLFKAd6j7dM5gHwPmaYeZeo5pqsjbVbRfU4oYZ
lNT8j9HW2aWr0kH75KJHhyKEeNBpzWgIlxGaJASQOiMQ+TMu4effUfcvvaKnOi6o
Er9iKSEIJA7g954oEXQm8oXeVJblagvzaJGvpdfnmwK/RpEr6m3oyEP/IESFnrsA
I1BNxmn6Luc11NSDsTkSKbnVMondkJ+W0vuO1AbsDrAEpUXEefJKbVJH5cEjarEV
SNyk9luVCqHRGlV6roSc1kwFe4ZGKNr9WoxO8G6xlpEAzhXTck4raFZWImT5TtM8
o8e+LwFdT8/IkgTkeuSbG645HVljnCCpbG6+vKtXoulVIrdJZPbOVPneRE2GMlB7
eQAZrRKVy701mtJsK2otR7i+L0FbMOcywtbKZ+2xF9LBrVqFJFqKHP2pCBEusgdr
FwD+pZX0jxrGp0d4IHNXIfpNzhKbJRW2vfcxwdIObD1GKriTp2D2ASkO+yYj1qSs
v6RQc0cnH3OHDaCAD7N35qqsB0cbq2iOismEeUAYMLQSdjyJUBlvmpYR+mjtlT76
gm34OfgHgAIyZyWOhieS5Sk1vVSCIQliV6xwmivxRONwug593KCzmmMUMX+uv/ND
RxK0Rach3iYVZhH4aBBLEriJG5KECpy5ffSaQIXlIOlW8UJpT2yFZZQzrVa0m+oS
stiWVYmte1lK94vIfVQGblWJwyp9HDKSGTY5pWoSpJJM3c+HY7lSXLtJoqlaHdgH
hZ6MYdrxFNSrPN1giV9fQrV32sgF0NS8lXzh0ePtZEjsd1pXb6h9e2up7a5lrcDc
4QcIdoopXkcJJa80X44G3Pm/7oCt2qq7hA9o7JA25Pqahmgr7LjlvADlBcFTNbYa
uMc0HhefRCsNkwyPiDKuFPEqPgZQSUrWckJm8s+WxsHdKB8vL4lpL1YEbp2Hhb9f
bsHUzsTNJOV9vkIG+viUOwL9WdNoHloAr5DXFtkXr14BWi2kOaD00es/h+sDAr6Y
ikQtxjRy/h1DwFZu4XdzGCnNslRp3BVVQJfpf8m9Z98zJ2c4GjJgPxl/p8oGhuau
zt06k38yaM+wh30szaU1XtNYn/kF5OWwsQpw41EfgWFHtk074YMCcpqzZWQIf/gt
Cc5c8Y118g5zKtbKfqbIY6Xcg4+R4AOSbw3n2u6nDLqgbVZ2+VnhMppzXuGc62+9
J0ITl/JwXWfo+/a0cypZFIY2xI1VKOG8knfOyQudqQBgapNB51i5j0GC3Zj5ech+
I6I2f45RrUBOe3QO5CuzPTKDI5flFevlnKy3HVOk78HmTDgHVP+k5Dz0BAIsJfX/
3fT+gQ5Bj2tb5Nc+sUScgIC5TyE0EudYr1pE2nCTJdq6/toiaAqvRUIFdPeGBUYn
OrvExgvPmTLOo2qrdhYW/SErawEf0WrSEN3iEYM52ek5xwpv9N+Lm96hnpWpGQvk
XCssNhEHe+AWlLa+Tty1tFgZ0rTVDqjsj9Q7T6do5u69CDYWiM4oEai2ZuLV1DS0
pPZQM2E0Y5P0PWrgsZUTw7fNkQ3C0EI+NfEj2x2MR1TuoMAC6NsXsMJL6/tNxopM
waH0H764zBZOs8b49rk86Hy1F0TtNv+erTsV52FzYHBmWSK7X6ekUpqspYLhPSrH
WbnDe4XZWI0bKhmQIKCco8CKSJlRB8/M8daHwWDhM8KzJc3AEzS6u/OP27a/m4+I
MCp9NKQ0CrzUYKsciE6aDFNNCoTb1Docmg2F44RAq2x5PhNEaZte64V1fcY1HcY0
E12XvTr8AvYFLk9iqJFh7R/nfU1b25tt/Cw1Sn2cidSHCLcJpXWKCizVDdDIU8kT
WYqTXw8f8dvbNg7Sy7wuh9AiRLUW7HN3oMP6WuP8MNWIVNuJtiht4nwEyfMWZxx4
Kqjusrsulf2I6jyiOkHZQeupglkrhALpShvwmR3IBpLup2SJmgFi9MaOiCbCbOWU
eT9ZvjoJYhWhXpNVpy4boZK53TD3MebM3KAFLEWfZRVyKElZCKFiox9GphYHCXlH
7GeCnin1POpotqKkv+n0bfESh85DY2SbQU+K7/LmtggUiC6h+aLDKsferb8SYwFs
ptZ1NlKFyildnXzJR9e2eqFmM8kmZleHaRFqAWNaBKFSdHWrMXfsHGO463tnIBd6
UKI22hsx+NHGiJgvLlQ3sausur2I/Knf8LSCS0IgLMMdAg1F4MZarFNR6icr7vdb
gyEYZHnEeZtAD/Bb9eWFt9Sy4ukdEQ3YbPPkZKrvdNqW3s25uDU/cO1vmIvay9vv
l57WxW6ZbH+cATZEpMKcZh3KWFXAMfr2YHvGQLR7dmxbW0KSnoDwc9enOMYNvsMZ
F6ATJM7wqjdMUvWC8pt/0NNu7XNsYrfwMkakzFuwdPuQPpQxn3ndsNLXpEsG7kFj
BfzKZIpSnA+6AP1mi4CDMn7Uj1oYrgmIOtKW16YIiLR2tQJ7VxmHAif0Z/UZEfq0
5ntf8jeX+MmFaeNCwWb+AxEdktSEGzhZjhKeUzYLRrtxyhpgqJewzaJBAwJ0jDs0
zuu63JM32PAaTxScoSbhVNu7P6LJHPJzB9p86LUCg6bD2NrPk8AlXXuRP4pWhkxs
2AN99sou5dTRWp7dkQT9QfaqPseaohYYi0J59FWrtlbySccZZc2yHenUBFYTh15g
e7QmVotijO104/ljC55t5iRFGAYjbhGQHK8Hcy66+YNuuhaBpYHTNQwaX1TySuOF
qo4r4TYiL7TmyZx730lEhpEwjXm30mLa6lgaqhydGZLVbQx2xTjEDypr29WnCthx
mRTvWJ5V5chLl3YkDWW1Ftnqrfpk7PJYRqxG0+L75Ob5WkDVgY0LMsndGKZA1oEj
3WS6VKJslwT1IdX6g55vnKuF8wKgtS5st58DUnFHr8fiPSVmO2SLip6ssR4WL1zN
9r6Foy6wcaBbQUEnwvxPSc6TvjmVe+9rck5BqnpmlCO5buvtDXA9mkBfD3vCll6/
FetjN/EqMBEo+ShMJNy0E/YcXOxQnLOPklRtkiHrUu/+dowmV5vuscLh4u0hGy2a
lf32p/BFVkNu8XTjX/goz3TeE5K5Vz2htaIqVY909J85Gae9GFjW5kGKQQ3NM5St
sMZfmWyiKipBnJuOyV8g5DbfhPTHDaZowSUeLw1rzdYogTVQfVX5dGhPNAmB6kXg
/d4Z0Du1uEjYoLGs+1MIC95MPncZJ5RCEDD6vSJ42YXK0JZHy4n50KQODSPeNLpe
pfaPiaC9b0AjRVQnUNTHFjaOx705D/8orG4+H540HO1f4GGIiFIzwJuxSf3VKru2
zj/xvsiCATKH1g6UvnWHqD6DO91RUCnneENc4ufr5ih9uhbro1GjJ40UDiKozTvk
54xfvSOPsFCEvY3dMWGV2Qp4AQvQkdD1mtJTFlFHBH7iZgzwxMn08ouUOOo9dLeB
8Y0I4wRiCuVfVjDP3/O91o2P+QpmpfV1V2fb8AliijDapPt/0y7BHP/TVmGyrysK
ecIDt/U4L96v1Pdg6QDb0bGxmqh4h3S1Q+q8wn4eeUWgbYIIqqsJh8s+JFf38aUw
d/diz3pr3phI2s6219bOt96zaljGQFmgqYlRzKqr2z0c9PpNuV5GkVxzJ52imQ0Z
rdy8TGbWx4AdXR0L71NYzF5aBGoEzo5qIBbGe9l0QZ3FlzIfhYbnt76hkJl9Fw7n
WKA53vQV/nlmIYrA4Za1g1MAeVXJz9yjy0FVObSLsHPYahKYuiv2TNItla9tkYxe
qibl8CjSrYfCJ+yPCt707PTpJJMl6108kkC2sYPIWCgQx6i4AqNVLj69QAysJ+Ws
E71pRiatMX1j6D/wzWGG9N6hEp9YDsamFH/9H5BVt2cR0UoCDS6PLqPRnO+4m/Wa
QSlxYWfZ0BZFSdqXD11A+mRmRi+tqBmwXy9//bXibf/L6vq6mNwvYqxWjqm7UIrf
rTmq1dQ2VxWVXkBQghKWSOUOiD0px2g4Yhd9ZEsg548ssjr+LTLckIQTIfTvqIEc
KUMjUJFR5w9hvtaQUW3JBF8P61fJoAr4tFX7Q2CIzeNhnCxkR1KCL7g3ilqx/Eca
ctjrEoAH8NWTaydW+muPcUOFbmZfjXCjpELL8K9XU+WYRax2ET5dCWvO7ZgDZO4K
+xqsKzJoDaC6ruAwQKqcwxAn8nKX5tnvQKGQfcs27ykvXf+x0LIj+z/wu60BlDWa
tPRT11YbhOGA0fM0rq0OOweyG0bENInoOl4QcrFP1e6xn7j1zxXSnsMV/9+QcHQK
vdccID0KcXF7PEwDpBlONwjhVQx0zPxcPQ0Ii0CqmqdMzElA3eJC6L5WMgrZJkrW
jP8TJPxLivy+l2XjDoH75Ig7/tyGvNkwrcm+ftre9zC9StKA/Xvw8G653v1TJr4e
QiZfosHyigfebeaIbp1Al1r60lsTneLTrkwVKEPAi38k0DNNIhMPo3CXOjPDHxd+
nja/VvNacI2IaX2Mr4lxoYBb2nCosTxG45OH4V51i1kuh4k1ZPZI8o07JOYIa9cK
rIkoAmld1wKuqt+KSGZmMi3UTEkcOz1bG6Oje9n7+3W8gVCNsJpX8x9JPY+4zvIo
b35h3enaVIxoW6NrZZSyF3KTAovMPWjZmMCdC9G09czD0oQQ9drQ48oEjjOMMUVh
Lf2e7196iKVFuN00Ew4xrKiKMSg2To0G3Bxv7VSKoXeWRdZADP11JLkuGeYrNC6I
9TpsiRZQcFrgQt4G7CaHKVjCZJriv/TBEpalMi8EOIcUogyG5Pzz1+UDsF2bYWXg
vwLYKED3Vc41//fBKmGH0L+YpVXsRA0ReoIjA/3C/h54lc+WO5PRHS9bHYwuQVBa
l+80LfC4zep8p06J5txXzozhoeNWfJpOlqZnJyKgL/7kvXGxMnD2stVEM5klXY0z
LVIgoue+iKQvWUjdkKgtReTbUlcJBqg2pRJAu/ZzM1F/v21TcRVgsCdMlbBYTY3L
ClhVjfBeGfMb+evTw1QS2ugMtIzIaYmuvMd6xjUrQHQlSZLfcwb7fZO443+3vRQD
1jDYNu3rs2dj5TyD8LcscL/Oh943HC93cz4RSEc5dUW3m9ucvFuynKhJRPiqeTDS
7IFf6ROZFTc8rK8S50GSybpl3RNnLchn/ku/ioJ+VevTrQj3L1Z2U3l8p/yQyEVG
JCw6NQ19peQK8161uGErhL/PI9jrj9JpLEk9Z91gC+oM9/NdnjKyGIm1/Qh56Eoc
Ul3WDt3k0eqz5080M3jKS7x0WeW9KuliZWYLR2W3RN8usRS0cdlIg9tqEmaOGUVL
MCj68qKbc00SdetEVp57oJWdpf+6OAyiZo+wzXEyoeHhYoVFt5qyApJntQbPGQxf
l7tssVAR9qampcV489tw03iwwWrMLy96WcpHYIxqefSxCSCrYcZfxEHNbhbHmwzI
z3I4EPUI0aOE4ANG7pxVhjHMkVSdYlDj1LGOmmB98yifPiKGkNEcZCmKbqhE9stE
xiV6R15/ITantqgxdqMm5rw9tAN60SzFxKo/kDB7+moJSbfOfeSPUF4GYymU0lc0
vsQ0LyQENt5/ZOYjFge4tdyhvwdhbmjoBdK5FWeNuDIu+cG8P8xIVWYWuMfhiLr+
JAocbi2PzMtFUNiXEm2Uvqg1IZ+PE8V8ZdDa/E7gF6r+K2ioTELPxPwhoTgM9BXw
7GM7M9/DtlR7ZjBx/rU/lb4owVAykA2HfTfNlpdKCTLgy+529Rx2J/sum0J5bcdw
f5HwT/LH5EI0obkSOZ3L9yN5tiS8dt+zlre4SguXNFMd7fBjbGp/zL8nZH0Cv9Ll
WCECFfDE0Dwf3jfnY+YKUs4Pog7DpeFuJ6zMjr54QX3DIe9rcIpcVCNSZtxTpwpr
L1MK8R+JvcofQYzQZJ4sZyLxa3/5q6aBHRvxyjrxanEZI/UpIbWYmw74w/hZ0b+t
1ldSmoJrczJrh5ENZl7tAZlCk5Oy5KPpyB1xcx9G7uSRQTGZ1CQ82FxKAw6G6T7k
a+jDxQGHKcZ8/GFxQr0P10uqLWusKNryH5IDGMGp9+mqG5OEUysF8JiyPA+QhSmT
Pl64Dq3Y80CANThSX63118ZUkMAcUJ6ytQ4f8s0nx1KEFczP9Asg/h3kjWn9CMmV
ucDMkVu9G6JNcJImpNHSFEiZn/rgdvKqF8jwK5JRypxNhxol5BEv7FF7ar+tN9zz
lJCBq6MjpviNGykfgbxhNdsZA3jUMp5Zjkh7urvW4Nm00HVOiKbzNJy7jWCQMeSh
KfMWcY+fGOxLtfIYYyqv0aq4Ci0idtBkNr5LTzwc225AEKuprYHrqcSA8A0xT/DC
4cIVYUVd+u0UgH/vfzlMEpoQ0l5mE4J+QkiQZYo5PfYlp1NyEOxmPGF30/VDcPli
aQgPPfeesJDMX1lo2E774X2cmHPUd4SadLNqf64bavUDoNJYFJK3b34k/wA4ZJTm
UhqXrKhfXS2ddrSRA7FC0C9rqe/MzH5EgFNLbjDUCorbm7CIeBeDruSopUFmYphL
1F18haqINFgNZyxHtH85aZKdTvpKyOz0mdV85WG1whl0MljF9ekak6acTfx2PDbg
XReVk2n/e4hEPzsZtw/uTV2mrLcKyvyxz1brmf83pOp28PU+xJJTB84S6OzRBClv
PBuJp7O0ODJRWsqf2syW5JGiIafYCPnan2x1Wnx7mov3uxlT5+3rQ9bCmalEjG2Z
nuP8TxLZ3O0m85MwFffKz336xxzpUw+JWNGX0D/CpbpZLfWb465RVcijX6rV+2Pa
7VQS9bMJQgNJMM9qG4PbtTe9f94xU/eaOosAi48iluVZzEmdNZc5rqnXSNsSM4Fr
GC38itEIJ1KMbnc6/eF7hkZqZjmfACCEpfxiulbzpmEo+IVKRFuw3gpWUEyaGVwO
METDllwk7Ioydtx0+ztSnFfgoZdU2697vcK29NiDF1nYzX5u8B+VYQgeEv/7X3w/
d4pANhJWth1uhjGCahWtheGK8C2+OMwghD/6Pvzyqm8dWqRqwvhNjNMsrXBOtFY0
5XUVUBskdf0u8SmeYoxyPqGHtkze+bDaR9CkNPgQvlOICvXvFAWO0cKr3Z/mfGhu
whawK/pOBOgD3vFaxYviYk5xKk/QhHVKHBoLUdPkw/CFnB9voGSx46RIHCpR1h/N
ke6XmDcU8Z/KCRzDgXbhgw/ZAJZPsEKVWLD/CGEcZHDrntOgJ9PUj61oOdmQoDPL
AGvHOec0lSiN804ggQ/+XPzA7/d3o/mHK4d6RrpFZLvo4Va+8muRBnwL95Zb4aTy
gArs6gsiALLSPyOGFCq8YdVTPJMFdQD3i/+0XeD4kuHgaBDPwWaMx1UVisKnOyoo
7eiJkf0CX/nnXHiyxr40BeyFlZV0E4sh4G19i3FGPExB6x0gbCmj/YarcoBNyuMy
rfQtuaNV3qavedSmTJjU9OU6epbnwbqQHMGrQ5C41/MTM4Cf4lsx05cUHU6IWxpf
pTjTjCyfOctJ5avvfcYvv2rzMBg3PO4DQY1oYSEylWh+Ndu3uWSmvmQHKCmrRxLH
hq0pf2iOUdiiFexBg5ThtZUZwBaqrrXlDnquXq8Kq/u6biAdxetZsChIakbRX4r9
rhggwsMRCc0nPqbWKQsoC0GdegYaKabLY32kTzlHG0Hqh8EN6k8zBHTPPfEfog05
s6xJ26WE7xS2s3S06acJJsda0Na/vmeedHSNbhNpo/GofJD2fW39ehG2DRu4nnkQ
14ZWhIAHg2DaSMuntjoG3y/3nnSBZu7BClZsmRe9KSUvxtmOW894ud4b6Ir1ii6N
TksfT+39YGwMtnVJO5PO8OrRwxYuhBpIrvliza6Xp6F5YmLApe6NWRyhnx19BnJd
0S/I+U891Hbi0BfQHP65DaF+ggpfLQOuUP6oxAX+5FhrpLqhzoxqZlJ0qWRuuPBD
NK1klyCmQAQ0qqkfrl5B2pRHTVjKdyCy09qbWlEQwBgE5I/PGXiMUcmDp3gA4VdN
p81riqeP+fRI2RFsyHT8I+5aU3KaX4L76boEcFLTSAK3tr0+eZu+vZUv2elJhbzl
0xa1fQdieK42hJebES6ESaU0+KO9kOwc0qzStYx41M0ldmCAmouBLpCYqN9ify2C
KkxHKv+lrFEZ9LWJMScfgYmiLitCAUAHTrj6g5d6+YH1SiYChlvOuAvamHjpcTeJ
ogHRFspZxYKSF+PzLOe7XWtOgF4XF43mo6lJaBCMlOXzFgG2EF4b+M/lrriP3Uj1
HpliFygoeIyuZdB0lVGFGZJEidi5rfd3ls1UGzfPNux8EMZ0i7UQPEJ4vIVTbEeR
rFXtfbATVskWNnCdhldim+qr1wTjVYakVFUIRmVNAr9GZm6B/Sk5wjchKOfbWW/G
UzF8nHxJKykKNev0sv6vgRsCY/aTnozoHsur1zNC63IvXsl099GkuC9A4TQAGwYa
csxITn/w7ib56c8f6BBFbOlRL5X1xJp6qbSCPjv3KuITY7o+ScKGpW9IfcSnuxm5
z6KoBNYYbba6Ax1ru/EyJ00vRsFxFBGKaNFlrTi62ClkHtS7TORsiRAnxj7ec99W
d7gaFgf9kTam7ikvIG4qGoXRBoKZXuGnyQ21Qg+pPDRIxdxDaoMIFWVHLj4I0ogr
roAr8mVPzJZiO70ExiuxY1i6NL4jjYtSysQuyJo9mCjj5mauymkwq80+zD0hxf/8
EnY+R/b6zzpCNMMjx8P+0N/9cJmBCBkhtllSP2Zof1PIxc1nWwDSQhTjONLuCXE7
q1hR45ZrwkMj30hxqwaxVCzjz/dOayFJtskwJoeA+wMSH9PCTgYPZQNOG8e4H1KI
Gpx5r0jWzSAFb2RaJAbBmcPNrkMnYPeTsks+iaY9talpWgxB8S/WPeS/T0i3nKUu
2VfnO4M91x/H5khnpGesdI9Gus8+QvENKn0n4cRwREug7U020lN3EbpAie+cijE5
EbvFmkQReKNTKBDJ56Iu6K5d/jPPSBt1X6B3Lk/tkjEpOBnYy9yGNplMR7+4C9Nj
f+BWPVc5DoCK9o8BCSb1wXTx0QzjMJ/BBuxbn/PdAhCNKZQU4bFae2O9FumWgj9Y
jACtppJdJzd5Ay5RD+rPkcj137cLg+c3P0D+IlWYVbic7JBZ5BypyqQgCEaFO3D8
9yKtl1NmFZ58nydRDbsperG5EfmIsD35eFldkJKEdmdPKKv1HxoYvHMiWWwn44/v
uapRGIqcRJyMIADCZrH6O4uaCnEj7wkFZqGmKSFrjUuWyyWnCW4qY/6B/oJhK6p8
KrxJhrk0lRFamAFDOiA2ibfw4SLGch4jx3GEbYmhmqiQ0ooe1TU0SI7vhtb0QWmS
9McH5GNuhG6i2hrJufCXJWjeVScMDSm7s5BMRQVf4PbgfmfTyIQhS+4oTskZLeSU
UEG6gSnOjL0Qfg0KBFLRXo6l6e61P8EuVvanPsDtzUo+ntQ054rNBPbJBYgCeiMH
2PSCrxE0suNrLuiIOcdvjhECHYVYGS3Reh3/ec5xJvsFZSzA9wYdrxQawqqlcO1B
5UZWnZf+ECZPv4KQUTtiCN47kKibzv9RcsI/5fF38pLNuFnBTVg6V98JmY3SSXrF
hqv9HYtyscvd9l/iprmt1owFyOoJNbnHviK08tsMnbiyzztIZ3WpHBpUtLaE9kVD
kLwSpMiZjVxKg6Y8aInGQeJhwn13cP+dEQKTsI3vnSmiCQi1qN8u7LSdz26uhFDF
B295VnskAaHyNuXJ9JtmkJuv53uDMJ7P7ECOPw+HgpqtV2+zKKCvT4r9nFrIpX+X
nz636p9Iupn7hNWjCOn1Kbv5rscbVdfcPjqLffe4tMtmO5zcVNrYV0MeSyO3WtSS
dv3qyQYX++cr4Q6UWPIxBQ4g2542WLv0E45uZCq0f10NEiglan9FSa/zGkkRUAtb
l/ZQxYLac1W3Y7raLhOUe1ZXYzUdYCfPxYm46qEifodPdzcObuCJhrdD4kkry8Dd
HCLLrKA2Xq69pI4MrXfo+1enFYQmmuxeSyBNm47R8ys1Y66DFR/34GRKcs5Cd56C
VLSLS+ZY88YlxKXXRaRPQjZD6NERlCc31gHsoBea1kv4LqLGU7RJbMsEKRsXV2Sl
nbiVwXQOi7/hldL+c0sLDA94Sb1f7hqWWHW5Zc32qxccH8uj6kiZ0DO3YXj3SzdE
jSJstoRasR27qlUWCSwSoJTSwTDEb9duLe+MGeW/5n6JRo+VYbw2vZnmoxxvWFLe
1TfXLdSfvjOK01YPho7M/CkQpHTW8KkV/Wu/+LLPncv4lYHMnq/YEQsg/1NmUuZj
SS+nc+snGFwX73XjZD857L6UZ1Bis1hXB9Uxm2TJBqTBTZhfEj74x5t4GCErckTs
CW+ZZ0NBVvIadpV++pPJYg1fQ7Hg5i/vUWc3g/Ogv4wL/NmQ5JJzPLea8Hdq0V2Y
IE0gQLZRTaT/WTnPsJQ6qhR128JhdLvfCKhbi3RsFVTNMP4vwklXBXHAXno3Hf1A
AV2mEU4epoo9FT+V0UetL2o89v/NRtKluI3Yo6jCG42pchvA6LpMezRymglAIpvg
PJKJh7Rkjf5ds+iHA4rMzuEXCKyrFY9A7cQWSXCIgmV7g5/68owHkJacLg8jzr8O
uB1opymaqx9cNFk8LgUmmISZ5FahKZqPwi/E9KwkWcBv4E0sjTBre0yU1nQBSH92
zhiWvTI3Ly/qvkIgdvqxPFF6gCQ8q8bVcOcO5IJv3wKC4nzzZMF6Fj7bYmO0L2wK
bfQe/YZCTQaneL5+uoKdc3pJzY7LJzKYZpfW4tC7RRivytpYkTYT6h6cErVWRHhz
RGd4mTeIgfZ2IDE7V/453HRaT3OLVHkjcoC7em6T0+AKdHJbcw7qXzY2sXKm0A4C
MjcCaJJbNLT3a/972xlT572XKUzKyGtbzSif0c4F4ieCccbOouL65dwD/19tvSMt
dOqcKycSpDMDXJvOqvY8RctSujW+pQwEZzJ4x9RB89a1MVWPmBfNJyb+vPPuUUUK
b08RLKUkeHl3c3Lv5h9KrQ/nX1NLfqa6MqaYgVbxNnvbhETXinktz6y7yyXpmvaS
FX+Ik+1sg/tF9XZNt8ikBbVdGB0UG9r3fcztdFFOpy/bx/a0uhzZhUflFhqiuthp
lMPeUxMTmR+wPIMwDn87vFaynwGs5eCKlgpFJtK1wTWUZtUX/ApPZH1xHP+Eq5Sn
nyj1xKKCxa21vwkfXjILoSHdLhZp27dPCH/57U1DYATZjWlSPBf/QGqZZ6HZb4XN
/B+SKzn5ttrFK/yC5I8Cg0hJgJhojbV49jmHZJdUixGs9DtyjbahlZz5FQlN50UH
uzmt0pu1nFgVEFI/itLrNqLfPwhgMSyAFiAFmmsxpcyTTtK6Z6L7KPX6Uye35XDt
R9gtpPs71TM9YcNOtQ6Vh6tsCRuIx3ojbjwIV+798MsY0RRbmelkrKLabSqsHohy
JTieftUhE1P5chfduzIskT0+vd4Y69I1vMIdKtegRCczVLaIzX7/qg0lLcdHw0Df
/mOrybOys3O7yDUAcRHqeTj4NF4EKvVERZLjIsf3YhZBsfvdp6TWsJC6p4IRj8KA
orKCd07PYrzail6mu4+33GRfcokqeSnGmcesAIPKz8x0Wh10QxNaWBE6GHzZKqsL
wOl7xfEpisUsoYiyqVqd4FBVnT4zaTSDNm8Jm5CCLBfiPcC7wNx2iOLTdijUPcaZ
dTK/ptEXuW5yHEjNP9ZSFJSwl9GdZ0dX+gfuyJBCJk5Jla9imnRQqazGlJOqXvV+
Xood5t5XdFsUomh398jk8/74cS844ceq1c1rc/BrBT7EKMQKnmE/I9vFGtmWBkCP
x9uLtOxnuqVVHn7LxNsPzguAHy4w1yAxyJ+NNeON94vDHUWAMn0JqA0L5W8WB5+g
hfFpmL8uh4sJcIXeQsrdB1RW2AbcejdyjYMYBrp9KGeFt70eJqMGdUG8XVk1kR+n
xlpGd71VTW4v0JyNYtFaxP5Jc7AGEGiIxaQtf1PGPFSqLPY6C7YPrphXNFDe1cUj
N1gFUsgJJ6XoGaYZxyLWoGm9rAGKLcYt7eamVpZ6KJUxqqO0zItodxfw1ithxGGu
Quj8gT0D+PPimApW9VZjK3+jF2cP0KbTpw0G/7uiqybD2rEJtYCcGuJnw3i4eQWV
m9pRhQ5zKhIRzQPkCIQ4HsW9L8kv+B19s49zoDCwIlnt+8G7yCIL5qIMdSaw5i1e
SAoq35ypM+T5/5hX/iskEr84FBpa/hP0Pj30dd/sYJGpGwjTpd9yjSXlgNEG/kfM
FWU4pPYGcly0rBtzEkAtCLU75gMZaXeq+6QSsA7E1GBYunJE2fYBvIcVefJ5/Q1V
oFqcdb4dtB9WY7mYBfAQcPS8W0rXs22PMpYk48ESdF6k095LJVf+1iKy1mpa+y2O
JYIMiAqlv87BDViDlyjzdBwdiTYoS93qFBz0MPt2lWdBbin4zweno9xFlstfF/Ui
sfRMdYnZTcBtR50O9VC2NvUcyMBsSxi6oaVorbvWG17ugyKhBkN3fkSu8uwGE7E+
LXgeZXCg2rOtcsU5QqXMcZAbXFrM6fuT/wMctf4eKmycGjYuNCCPr6yde0l7bL1J
VJWL4Ty/7b82/JVZTGCSfsPZkGDItnhnHTJKsmodttFAEing49iSbMvgkoYg/TOn
+Elq8kU5ZJ+A+G1I6Tsfirt3YM5D4l/ikW00BpJVxycra+oKwgsHxl9rdBZxeJZL
dk/l190wGQDEj5ngq0Zo/AjMH47lI4FBex6J5XIVJlOR6kaLUrKKJXd7ruUulead
5qAPU54f1d/sdY+nmZ1t8WzyBi1/zs9CQkMpQvVE2+mcyhSaTJ12FRNA1rAFd6qB
BG4gJcc58CLGdM7Y7O4qhVIj1FpEtH+CWSrHvzzd3VZEf/FtpZeazN1QadEPFkM3
BFhGSqlUrkTZ7/w62XN9vMStvM8eC6+Brdzbkd8Z9bdi9EVj+JXZ/VbWQwYUEhpA
p0R6VutIX/At/GzKR6VDkMrDRdY8owSqIrQbKorFWWZFKZZCPqq9/P8RmVaqKp7s
7lOkqar91eIaS7rgvIEZzVwhinlM85QCm0Vl8jjGegIjH3lSI4AtXLZ6ZQEixZ8x
X+TWyMfbsG/GCdXzEuUO7dVriIDaYKJjgwKnf6cEjsRmx0/jIbKF2d1/BNqVSjVQ
r6Z7cnqZc+Hg1kcdsBegfcASU15z2/cYMjblCaReiJwfS7Sv9YGVFWazL9VzgW9W
gJ4NtCT5wSlg1gN6WxP8Mht9scURFEixszwelSBQLlw3gi6Bp5cg/BnmshZU6mZo
wXcRo1ulzBy7BxjAU4wmYNUAfwxE9PeMj+kfNk3l8zfjt9tlrLFpztPAu26l1P2T
kp22O6uzLV7LT/yIiYAmxdskIEfH8hwWlp7io8G7hqPrZJb4PKbqByLMfgiyRyVs
KjKTrruWr8UrQW1dTPtUyRKHEt/r6k1HXUIi8mNbNlXIJLuEuajEAAuFNV/J5qps
C7gwpFt2bw+VC4qiqDoJ2pV+KHEYUHxUo7Gs3iBkSMVON8rwlPBPur6Rq6/EJDzE
85P3q++Ohrd4dccYLH9phtinjoTONw5zSBPDuwDMQpAEuzjR+cql+fGfmI/gcghk
NJBZPlspZGZECAJHTSPlvXsBPsrk1JI9VVQwiBZG1S8y/YOUHXZej1fnolL8bh4R
gq9RZEXFOmQ/vDTF/wqhG89Mz/4XvCS3ot2LcgFIxs3DZtsiw+bx+q3NpiYEzo6e
uKsLrMLIERZouDZWyMlJa0bbAlm4Kz0hcwEZuUs4UqIyuqYOnUEipgRcrZce0v38
8sh4SYTmzDRK+TtqfYQg9dskXxvAQAm80zGDNiCSJeLd+SjAaaHd0F2dUEWfjtnM
riSIpl6djNYzwuMGwONLkgTKZQ1ce8E8SHTF3ZR8a3jhQ59iIvbHaA0Ng1yThfAh
avZdD00hW3wpzowccNxpC23XmhltQrAIMOP1xycIJ0lnny7lWf/8np+A7iKxw+T4
OI2wFNLF0AkL9iNkfFgqOX4YxsQyZy9Cv14gllNJ8bEht7GXnxVt5hdMFQgjynwl
bxAH8ORstwaCQYHq00Qqh5Rzb7HFgVkzuvfd4sPRtxm9Xxeq+6KEqf9pEWu0IQx/
z+3rMxnmtMVefmTNTwuaQ6Krz0YaYh0V9sKbu//K+Pb4H5ewxEAS540fJQrejmLM
5rOwVJu212oqoP67iHBHBD79g6NDkqUhOj2Ley8FXvRpCKarPvHshkEgcB5MJpOW
XeE6X8zzYGzF3HnuHI3qHXjsvC7+3iqy6J60tCpgNgezjwO0tt0JC9CMGB2YbCQS
XRT9YxMYAev6Jp7WK0/9eNuVmYZNrmdHyPAkQJomlhJC7u/1C+y7KCfAYTdnFfBu
Mc1+tJr3lxYBRunIRTvQAGJX4Z0HcqArrvUNLmQMGUGbxRtnAcw40GIu2JChJPLL
VCnCcvSNLkwbFfPiuyPTJx+WZQ0xfZpS8v9t3qNG/xbrYM/mhLUW7lsBl851mYon
mAzymLrk2IFevccwNBqkGGqWKRDR22iRt832tC5a21wq3b7IwWtkZ7qf3XBAwqnu
Okvk5+MYnbP36MkljXF+eaxfZtx0YqnupjY+YaqtW5ftWoMth5XSgD+hmbaX+9us
Kr+r1nEyql4d9w+dmjoMbB6e2NcgqaOliLQqywfEps4VNnxLbVH+VZ9yWq5S2pXI
PkfrOGK0YgQSrpxHfu6OzHsG36y8p/Vib1B9QiFAqetSE1i1brgZPMSsLKva8arL
TTxNaR+KmlviHgCJX329M2paq2FOP0QHgulxEXfSTmZfWqyAKC+PwRf8jYA76NRW
r9Ivbs4afbM0W15W59CXLun5tbfWq9RyrCPH5dNCA6B5uz2URb3Ba8vuYdi4KVdh
fDxchk4jvau3RPa9M/mxrkTghOYAlJJdRDcceeqSxtJC7MvHsylHLDSKU3PHXnh3
xB93n7mgbIgf87ivEBNJByqvsprPDfxk1sYyUd/U6JiawZwbPVh5luTYknWCp0DZ
dFHKKLDX9PSxcujzTy5cXU+j1rJVmsJ+TCnQn3wWF+Iwrr+hn7jNqy9QNtCWw07d
TAtijpyWSN+Qfx1aNve4sU1TghnGIFn6NBeMRfKaqt0MY9HDhbUerIwBuDUYDMTo
5XLmUk45U3GFG6VWfwmJAXexDAhABxX+hsL+xURY/7H2ZvmaqQE9Y6+Hp1zjaTfZ
eZtArOpNy3XoiYyXedRijcICKUIEPa0ecvLdyGG180gYcw8cqaf/mFSnsLpuW/PX
cqN+lZCOcvKPpqN27IN1J3CtqkQ7zmv46+8dHUF2qbORHQ5doMqdz7W3whwe2HaW
+e6W+uoXDc248KJx/H/hcwCpnEI1hkXhCTfbtS2fu8Wl1oZR1nHQFMRmS4Vge4lG
7lx5A7ulmXwZToN7tGaiYe6kFmba3cLve3/xYI6BdzCAqO7y87aYcQSH9RsELoNJ
wU+a45c+lQLKAa9i+ascSjJitn5SqQvEF6Q64RITlLBzu3wfeWZd/jsRBD61h83z
sbqu5uQK9XqAOOpm/eihJALra4iIDA1zFCGNfUpSMcWP7KS446T5iTru0aMwvtPL
iRg1eyMw2tGhUqcgIikoP/UgadmV60Q2BAQLbWvxox8z5e1ty6SHAU1MyVCFUKsN
lruYLPFYhltkrYYctWEDmZCOt8/rNVXg+V2ok3y4xsQX41cSVlTA/caz+78s6i9V
KkganmW5yWMZnSJXlopzYo+XjsFdbZI3I7k/itIWw229EHFf+NozNz/zHu0IdAPY
aefOUlwTKiABQnCM/u+yqXzZkBu0xy7EXPkInYoYQNHw7rlzlJlWhXu+WZJ9zWNA
6IW3iX+4zsFW2325Hp3R8HPC5+O2u4eOMaRFkpy67ZnsUi+tmO+ZUcrmu5PDiZ67
w9swITVxgTO4UE4D3fpSv/z5+hzk+SZKj9HU+tqRM260g8nI7l2beYRzG38sb/4m
eOl06S8GUGZwpID9XiDiGcIz3g6KT+2Bg3hpTUresEfTKORZ12ecf3EauOBVqaKk
XZJD/IpkrAVrkJzRoq98Zsr8v4ixby3o+Ci4vf+H/eyRsRULF8ATDqPRnNXGLuO5
DAxBMeMNHYRPB6Y9NxxSRmPQKhrrxNO6D5X5Z9aC3mUC2CdVxWMMH3bGeV1+bjp5
zJhtF2jt8yJYsbQfKkoiLMaDVO3K8NYRRr7vE/5IIxR64kVHqpFA330gGHb6rXf5
WNbkodFZePj7HI/bnpfjgndIQ1dZ42tS8iAm4lgRqqXskcTq9PXZTc7E2v5u4f8X
IBCxD4UHjPwwOyOd+oTYjikWP+WyNQ+82hcLIaX6vvhgcR53bNZv57npD8Yyvs7K
Kxm+GnyLG0+HgJJsOLj6cZWVkHyyLwmP46QKIEvVYxyyNx0/loaN+czwH1mAx/2r
A+5xCym8kWu2mflR+2Lod/T5nQO571RKG6hALJQ64d0Y/ANJfrHjBXGZ/JJTVwxt
Vwra8IpZb7ICbysKg2TTnwXFJiNcIAdoQcUFzf+WjuSenDGSS0GGIVT0jsSasSdN
K1irBWGsZdcoD+Odu8DBsuJ9tlIo3IwZdce7fMeuRC09+Jg5ahud5/COqmEhGOwo
sE1T7Wx9PRNjcxhpdICQX1fKuobLfPmFBPh32pQHSwwd2XPY2yUvwY3u7zFwx+fw
wr2NbIl/VxWbUrItLvHSj0BCORP+loXjVsitHJY1Kh6rURkQC5uWi6RoGxuwCI0p
RBRfEwejtraD5o/ubVTdAM5l3q3KS0x/uMJbTl4Hrw2VR8tJ0HVZVzJRO0MYHIL0
owKRDbhROOombPDSns/yHcvVyuNeT06zdbJcf+0TB9wFIcHIXi2/qRsCqh6JTY9k
JJWCfYOZ2WprmrFarJ0AmWDI6i2wKqidX69q9rpGBd75KuYMD4maJo/UmYYu72J9
XKARCeeVkxiYbumzg5NSqo4g73FPF9cNnzDbUaHDZoh+GwKM/j9LkhpbeVc525kn
9YTCD2omZl6w04RvvIFVCPdPqCHHusqlL9LkEQ74UJkQPO0h8DqgDuCcW/j3ALHC
MautZVV2kqaojAWgUEdcl0E3l4yaWJFoPPAoaKoq+GugjUy1gBFF/OjBCgLxkiMt
DskP9FWdOg+VlvCCZ5CvpHACJUL6EshDg9yYfpkYUmQxfe1miAE6GbbuJFo8GOSz
SKPe8Y4Kppzsue/PLadSORFWT7Tg7/RhH6/ehtySV5bFc4G/rp4YuMS3BZ+bpyYr
M68ZXj9Mx5noXm266p7Ii6VPturS1ZiNGJlPDVhDsuIHzrDdLkPFiqpcUpdMLYU4
Zugow18jXKPE9hSsyJgHLJbYacGa+SKCHxmWwYVkKpd4MUygpYK2Eib6iLePeTxS
QY8HtcBTV3iFNMyCtvzCmMZAb6CHTtTB54PId30itOOXt54XDxJPfMl5oZu/sowU
qkvJ1aUa/rG8GK7ag5cWfdXX09y1Rbu16K2tYzRcxU5/oFAv03ASiBodD2grT+Hc
sSDsoD81UhhixTSJsuHM2hPuPJDHUTvHIfys7sS4YqtBl4j3pUEabwt8SMlvxOCn
sz9+ETrP7Ebo8rP2t8CbtWDJslP7lHmi0WkAGzV3j3P2Uup+amDbLlDeVrMfSvF2
bhb0KpgMzEwljRcRvCw6zsI441+JP2pZRquoqr4XqCkjzzf28SEjiD4BIkEWk/Mq
s2LZq53lmObU3ZnPkPc8QChWLaPLz4hc5c6LGDXsgqjPQ4XwCm7IrVVw46sZrQEN
gGmDtui/vK2dyWRJ1/X1FGHIrvTQdF07RQEQq+xzwZ7gEhgk0jRuoIyzpggWPYoN
BWPSqZo28YiHyFTMGHa3X3Fkb54NqSDW5eovLICu3dfrNjrU5/e2Hp06Y68JEgDS
sC3zSCXUk4t+AkqnGAXvr3uEVWbUR7cgxR39rwzAecVKw5M/GBR8Sa1S1KQroUe6
nyteFqW8Upkf3Chve2ysnroixF138v8M3wkYQvFpdty7qMaEQZVO1GbLeqKHiL+9
xCy9OJlxeY0pavd8BXxbZQuHOfwCJJtn7J7yu/FjMOxdpXhYJKHDU0IebG1wgd3F
h6p3LTTZ6zF/RBgDJXLe2Sy4B1GffRkDAwPlnWyI297Rfhpz4wU5n/1D8pm7IGgK
0Il69lxLpgnCNoan34Urwcrp7XngfA2NUeMbvXN2FTAmWmo7XYWXkW7yh2RWgxis
d/XQYG9IdF/vDlbdM9IA0LULtMtkkknh+avtmy90lH4ElaazEEl4gShOC4z0FAnU
4vqKjJGwH203aDxd5WqUM2HHhs5MhCnWoxSAW3etjezTQj1njHyZbxP69a0FabSi
jgR89WAlKfmMazf7Gp72dbY8bBjBvfBQytQkdruY1B10WZ1/L0LdONzA+q3TpVEI
nQVrBaVKZgIBgRrZNIZZWy2gjrheyLlsia/x6kIdcW6OUOzRparn4Ct0PO+foM1d
xqE/oMUDOiAmSV9X60bu9FVdxSmeg+83Zq6uTEnOqcvk00Ndz299XQGg3ne7H9+d
d523fQT4th9fVZx/NlHwBVK39hqDVQXj8+VvUKZ4mKquL0Ja/7WiHnCB4DvskWj8
e4HXJ6I9IwcThszFu+OzMkOv98nn5CQ1sazqWXFv4Tmaw3FHMRDzCxU75a0RsvHh
oP632US+B5cx4KqRRLTOKAUr35fu/y7vb5c9rWcolBN4lUwxVmbGrXJvpXt2BuKR
5WdTsgEAp0/zHBLhk1jT0QN7RQc/7xSxNJYFfv0LpOY6uG7voUKgfEovp8V0C4lX
gV8kWyHY9EGhLxCBoVCfhag7FBOP2rtHxx7yw07g+aHhrjjNkdCvj+qWoG+7/F4L
d+RduNMRo1Di7d35C74l2zuOw821BIfcMpiNQZgY6aj8/QkXb2QSTua70AW9nsbL
fjH8LUydstwEQh2TdaA4eMyJXDKQjpmBPdi3Ta2BT3wcMBJzzjhRfvmS9umYgtbl
TSKuJhcD9eWvZjhB0IP0p7AAotvvqrMAlrMu2hTlfx6J0vvgRi66nh9c7aJcK6v0
phmqKPqTkiasmnmkiuvZng4dU4N+i2Wwg0JllnDxk5821vEWtR3oaofHwxGwjHqx
odzHB956b5gN5HdBNjNe72XtkMh36MRhYpaJSIQQwM1+11GGj0+g77NWpaec5g7F
9QvMwRqhp4JDMVrlpRQF4Jka4e8sJMeGlTGnYUeXt3MULQhNCV3rUScI0xYEDS/J
aPj2QXRSQ3k1S8edvRtXD5PoyrnUfWF+eUKU/HnstEp74oFMbsbHyKiiopCxScPY
mTTI8Yp/w4kjq5GxFQ3eALtPGKQsJQPYLv9H/FUq3XDyImSnCjwQzkFU7tdrT/N8
NiafPMb4Cpo0yDEMcRczgk26GRSO+BUka2HeI9U4lcAFoBlkKbfWWZghSWhI1+LL
xbiAFBxVfmlJ5fLY2lp6fP9C5xOZGWKP89API5IuiMg+EybLSdwjwWmRKSdOlvef
lkMuUXatZO32j7GUW3z6YzWBfzKs/CcIWepIdQamowU9nOGnZee5sV7jJLXGFWgC
LHRfek2ZBn1yWkKXOVRGB/oD7YKxKBElvhTd+cdAQYGn3VD2rwQtZ2ZxqzbsAAm1
EVTZD92A1468yAQ78K/GmuHVUM36NIOP2PDAvfLiljTfW1n/g8jMMU7j1zRQCSdq
50yr1PhRNBt0isiTFWY6gTfmfwbIJgDXhMXB8btWaBoHb6sUCoQrO21ZDt7/46e7
93YLqVNQuuaX2lzGztGvsBlrQ5ATMv6TVyVtyLBiZNpmRYtKz8DVwkEo994h6vO4
ng+GVANd+AdcGXR+VCwkc5f1wXzmdI4uaXU6EFhcBup+ahLt/E8dfEGpNaTFVEVx
XxAdycPRep4/VVLt4EVgKCdRgGW60G2xBKe/402orLpTaW9ETXteZ5vrX48MHmut
/p08a0ZUOwskUXANSFNOE7jag/pbTrrZxOxb29ymsiFUQC/tX1aoLWpqYNT5rqBT
AmsBq6Sxv1D2z5oy53fAdzxzkCBUKZkvNRMnHzB67lNsPdTfMYaREi528TNITwhZ
fAuhbZgj/RrNseYKEX/aAwUqs0gQF+VKJfp5/QD83UXjLeSlhUmL5KOolckU2pBH
V/8RQkEwdHu5bQchCRSRd306zcnU8pYIo41X672k9haouvn0hCiQ5abWaaYGiqAn
Pg1dibsHX+Wvaosz07y4PX91gi7dOQYV3DW5y1JHcJJU/9x66hqBjS5X/WIDcAY2
HrR/yMJacMgbQJiyKaoXmiyqaCPBysX0dLwiffA6b74k9yExB5Ngz5idYRTASjV0
XSk/xTzePsgYHdMnP8XsA9/H2hCfC4OKH2psChRCs3J7N65WZRQM1VH8UGcXuvfo
JSDyuA7irsaUNrLIQeBtlVbkgOMt0QOb3WMwoCov79GCvM4WDM6OedqvMfyMVsmn
nxE8um0u7efBS1h238n7tb0f7IvukCWDHPd/Wvja05ejifydnFidvouHRF/sI9DO
jOJNud1qFytii8WxsA/maYC97dJ8xya+RXx8mWLSD2wK/UMlbf6e36/PVrVrYQ/8
iIaaesHniKKeSmCvpavx8kPU2MKHqrBP4VtfY2ntl4G5YwxweOPHYouO1CZKIygd
3I++6Nhh4SOjaO/+fvS20YfQreffSlUc0xiqo/UPS63W7OeAjiWq+ncS7Ub5h5if
y2Jt0b2sb63MZQLZQgN6NUa3Lg6gCpsxg7ofoaE2YWshitFHuQCk2ogTAA2wMfgg
JxTV8iqp2TaNWZa+IE+z6KlfEiG4wO7MvAD+czVjCJXbE1tCTQb7bJdxbYqz1YWo
1jg0V1sQbXKUjX8cA2sb7eeePebr6ort9baxGQo4RUdTXK0FEtogM5p8qVDXu7wm
JcXWsk/m69hwx77f6Up/d5pq7RAJGnjjbPYPuFq/xDZcocyxpLh8Bq68j+C97Fce
ytTM5soPcfslME/HPUyE/ZClY2aOjwYQw5DkUXl894D+HpE1kFm25hkpHXu4Le2V
RQWYwlwmJocQWSCuLthXCMa78iwqRTP7QCyS/Tdp4iB1vh0pmKcFx2oWIeIzK8jO
cosS93ocAD+pRLlxhBu39BSeFq3rh0uJWNl98JT9T7EzEo/PmXts2R9Mp1jcfwQg
8Wrmh1OwS10ZhFGnq4SGIDfGS+8o/JBoFwbOSBofIjQvSJE4xckkiPhIqzqqQM3f
zTxnyO7TqyMW9wEwGfDVgRal+UCQHXTooGqO9fLgZ50EBseXJzinKsWPj2gKDT8l
kgN/s549w/FTF3Dpku/PUUzfzNEdhIT1tMXZj8cq9KsEb9/sRuyslVF1/CH1MICD
ao4I2og/pVeQtjA8lVx5pViU3hh6aqV046RURNCCYNBEPKgNTEK0S5/VjnmSerCK
73P+NeqkjXeoP2ZClmGCmgGvcY8H9nf0tiV2J9U9show/i9nWTeGTurr2x6yHJbd
U7nqM5aa2ZWTmdWDZuRniAebDdgjcULt9nBCaITwn2vaO5PSgeJ5DcElYmPlHOc4
vD2IiQRTrIQMh6Skq9jf+HVAgztTR0zhu0iPC8XPDIg3B3AmhdmbGYXghaIDraFN
Hu51mwRVIUvBPrwXlTSrBhqWeaspOhohWDIjGI7FQL1lC92Cq9VcCfH/WhM5oN9j
ZQlFwK7t7jEIAlKAYVtOzPVxtNOjdX0s6BTBfXZMLRPYMGbscRBPgV6RGPfP4fjf
Cq64ixnpUM7lYSPzgLdGmFRs165AOygh4yz7wCqWLd7vVzf0L4z6v6m7yqDbeMU3
rV+9A2L8Zu9uXjvP2p1eUbFK2criYcgUKwArPXHRLhSEfauO45smbg3lVhnE1SwS
gZkt8BuUny6BEDql3MHHK+/A+P4htHmh3VZEq4zfdRyMO8c0Dp88+ABZ+NoGLFm+
UMDJET7demsig5VQpcSD5RCFEGkCWH5KfO4EI2oabnI0tYxH3ZnADqeexnCsIhP4
SiGOa4LhFnx3EnY63CmdXZF32Lwwz3+IVI1ZCkdCIZPOiAkVLSlRC8GJlyPZpaep
lROu8wkRi8J1cS7hR1bdmCEyPW1HtadBEvfihG9aqtM0Ufmb70RmOvG1FyofkMlI
cjqR1QsOXTi43w4psKTKPHs4W6cUmWh4zAn1wQl7n73rfTz9rEoIfgPK4CIussCe
lsGjM8ooJZ4uQ9sOHyyrIfb5mu5KlnR7/afsIrWlWmEfeEfBr9J3tNsZhwFgt7Ma
4p9+cb7H4urqftmgnpYyspOBp0bboq19yVV1Sh7qNdQLcxpn73JT9mTrEGLe0iGJ
FWNUWg/owY8bmOhpfdgQVtgaKEtrSayHz0xpnqn0iwEc1P3WrGyvkQI+0fZ1gPJ7
+MlqDJedKOU7lV7Ot9h2bnQF8To58z5DlGpK+dfMQy8GhuQ84+v49n2+F7ucgjz3
4ORd9Bp3s7U3Z+/taK7kJjloA2lXeHc4ulK+LHVUGtiYAzz1twtdMkVSE9jmffMI
IiqX+DBJS5DlzP8tOWSLiUATqwYxXDOuaOAMnjtJDLTksnxWvE+mbz9xZYCg2MkG
am2SkwZQEzRr8P7dv0up2YfW4VXynTEECl+wJXab7Fo5s3VDUldUO8J50Sph0QMn
Ag0y9/PxS0YPPkk99EvepmA0zVq/ZjMyTH1SEtTWafdoN+tjCl3G/Pc4ShLgtPRY
yr9Eoyqh4bb5leNuY6/wWmmdrDr843wl9VhJOGVH0UAuGu5NM14STqvZ1D0xEusC
mpyPrQnPkR2yqFuMF01QgJpzTOJHH5mbO9CdrSvQRm7FgLhPC3bwhtYbDfAPnn8f
NwiiRV1p1rsOaZJjhk6Gu6WD2cbFKuCNq2usZgWXwm93Qr5rQeuRqjfdYshDU5bn
jhdGRarjtaw6dWJ8imxQyz1E5simsIvocnA6hImGuvGeCI+gGtQMbeRLEkkA2foq
8O7CdEw40OKKXfqzwZqJ/1KNEin5+faPIEmsDwW4AaUXOd0jeSRYbUhtbW4yg5tL
0TcwnAOsk8RDSGU2KtoCei9fxq7NxifJoIoBKmp2SttGYvaH6QQpAsTxsNHefpuw
99Ln0jFd1xDl/rS1QNQsBFW6KCZJwbfbJMdh7b7LHrBpPIVs7+egztyugcs9xD6l
DUyrQozRlI/7SKNbZbFKvYW1gpfppBpoFcXcW6X+E1IEZ5xwJcIYvn8NCXuQdMDM
vRr3S7qP/9M2sR1KBBeEwfwnkWJxkOzYzdGJHKds9QulBba75bkHc/gYwpYMvkYY
Bcv+0roBIhizecgO8CIv6Rm3ttJ8mmRLPczg90ANqVWN5JciJUYCiuQDmlqJZ/Ei
mNkEbKQBqOU4xWsKkGwFMhhg4sKDk4UqUaL5jK0Uu7r5mUgVKIIGMDQTJ3XPUXW9
t1xeLiRMrilxznpVQYinBWmiKd3msY3tLzDolq9CMUuHqAqYpdHzn2XjOdNRHHdP
7SOR7Rf4VPzpg3mnmsyR7Zr3ckC2VFq/6pv1DtQMVs82wCaSw4w5p9R2KPpqXvTD
zUwjyzv/fXdWGSbOZN4yczpnGUzXTgJTxvllN6g5ItmHeeDSb2TecZDbbgNAy/R1
7bziC6f8JlacrAgvhqlrxAXS775uAOETtBvJCRsVULI1REDKAMybnWaI6fIO4qiY
ciT4ZopcKKc2w33K7NIV1uftxsCQkKS5ZgZq1y8210xgC++Da45WQXP6yalgqQ0g
16bPW4E3kKq9GJ8+tKQiU32H8JxYof9O8gOZo7M543Wc+/ag1KRHLe6wIBNNSs6l
CyijdcYMoWNQSyle0Ao3SwAmaCj9BiL0GAnYzML0K2W7CN5Ju5tLORGcUZcymN6U
J9lsTJT3FIlTqP1O89d939sNjtfBPfnXCzdsgonVUgc/6zrRFvpdndGxjNohLM/X
Pes9S6neSwPPiS4F/wJVKy2H1g3y7ZewRmbs/mXH38rZ3fkmCsnl7KTGQZcnf8au
SfjsUhkUOaKy1s0zxFJqSMqt/BP2Jedv1vMd8//bdhmFJx+5SABPnL5oXAr1LP5m
jy8zbiAd42T9oqO5ZZrz62k+KiAtrQGQB2+qD651YEI1bsoSIf5AIgfmM2Oi4IcA
RVZWcRZ0AeiaUc0htnJ8gsoJLDW+v/c81ycjo7YuF8wP1As8Z94ZsFI3MFxYI27V
vRlPMB1Lh6652ZfpNWnjkc5/yc+ZvWBTNQQJJcxchUeoN9xIqCZr7XCL1jI+XHG4
06HeW0h/KPn+R/MwSX6b27wDsJW/PrOWCY9xCQ3tpMs3ochMloZqQ1WYoQn37Hzt
TOr6DRnRR9h1Jk6Nh1FjadRWyggMUiSZ56Z49Cz43GC5bJyNutMm/wvDslOg2Scl
oC3r2leR9Atm24keImyAAse/t0bumovuaSISZnZyRdRqravdHT1r18bJMxXI7bB6
552XUNPeZA+FG9SUB7SVjwUKKuLkXEGYsf/rWO7m3Bjqw4XApBini/bMfMVoFI7W
ThnfNQP5HWOIksXoG01OkNovcOhUfSjIEJsbQoRvNCzWDhs+ccTL4xDpPxzfiUWs
+u+qrhyizKWpmDmgAQlozlKCiD2jrEyrnYjqIjvoTfCsav1Z8uPhD1g6dSY3fewD
z6ziCWUfehd3i3sjoEUVG8hWv2EE/INbi3MkHBeAy5h3r5qxCjMVNBgt4BOlkgXv
z1RZ3KW2eoJgelHYoqJPApHHRSLMjgn22Q8Q+XzpHn2ccbikfJdVNkK18hMCYcQt
aIW9CjbifAcRaNyPFLN/yKgkGKYOHxX2gbFIhPhJpi9oOjKwf5yTJ+YpMBdlCnDa
V4lVLoWTD/6eLH/FbdEFhKgGpr4R+SDBNOj4YjNcoMCOjIwNsZC2Gc0U1ApO//8g
pSvIX16nHLv96XRnZn3Wz5wiDVdvNhYEnhJKhYc1CpxORQKmZfnY+yLyRPeUJrep
UJzsoBl8kXCv3KegY2apAnIt4HP8/ALapGMWH9QSVdtaMv42pybJ/jzAdXJ9oPR8
bvMNwZKTcaZoBAjHUDuSJ17k9oZuc1+8UtwoYLSiZKnFy4PIYbXwsbhRC/2spJFu
3oqWzyzZs7kQio8ZvKg7keCms5suHP2uHRlh684+HHJ6joZn9iKlwZJ2DI8zabVu
j9vK0UiaJFywKiNl5iNgvUY3bD+Da36t4e3rfRqJQijNJPEzqz0BNfWfeh6zBWbd
ONKMNfaXYbiZyxODI4G9o/noi5yZoYwePaQ4VkPHgG9aqWhF2+5z/uAhDsR0CZmT
zoijn9nyJcGEkKF7vWy7tXgjSNZaaZ8LRgGxlsxbjSkVgu9ypSi7ziqL6Ss8G6J+
TAFR7huQFayUI4vydyeMRsqg2PmJTSn74Y06pZr7ZjOnTbNJj9ilnA7cIai7I+Gv
tywbctrYyuLmHkTbp2goCr3Xr/GGvkyDd+zWBj8/dS+eqz3wX+M6RQSWSSOQcOI7
NxIv76KZvKwziAaaEBSNJFfSRgKktKv0pCjNAqTQnsgwX2WAj6Ob4WLXf2F2LRvE
ti/x6q8h69tn7FFLC2v2Cw7MkfEjtV9W9/3UQO82b0IFWWvG6ET1owqQgVEez8Dz
R9Nv+awONrYwhDzFV5R7YV6Uqbv8CB/Ye4QGMIv9Ro1rKC1AjQKNiJ0nC89w4rxS
y/OZCSS5Zo6mvUUaIZBI4at9cDe3Hnw2s4K0V1DToHsISCTv34Fy73rdPAB4YnsL
T006u38ZR+Nhv4P0XiMcqbwouYstkFOcAshFyN3Diu3F+OK1XoZe89C/g2/qRnEP
zt1ltB2rz62xwcCGua9S67FCatkV24Us2WTmvdUxKIefT/eUldWmDRnNbXDu3Eb+
YkLauy0cwj1ZNjjLo6yHNIReWMlSE5BpRN/gyirc9nwJFkCc/QFQJuQ4gZBwESmT
sQwrodCtUEqlprnjYiryZ1y025r7zPkDywHaPJw8dMOu7dWSQ/ICmo7x4bJYsMgR
dNanGlLTiuIwrC8uExaro9ONDUSkJAplfvheQVw1WIGOhxbbczw76+iXtc11hnlM
iu4A7hdHfPaZMR7U9LyneefcG8pDg6JNC38U0keZpqeB6vpjaSHjzxzRhO4arb1b
dmqycBU5oSpNDKeUIDzeDczBnb2QzjE+t8rJT5fAJBrhaJeWazEgbMOHcxZusWYo
4Zq79Qghl6VKQwYPxS81hFhL/PsXTjpNiOuYtENSOja7TLpcFHuCymfDViIOHPpc
69fqr0axah2nICXvtjam+G0/bc4UNd0u0sG7Af1Xh+hOXQt3HbqvQdxmrSt99c5l
FXW+9C0mpX45R6Vs4W4m8QIwabGGoy08nXSBB3TLifMFiDJML6Zl/sStIz6MxTi3
6u0n7YybXJLDFIDGCxUVwPaqmpChkysmm6j8Trbfz3n8LIUIusWx/6X1UzyXNn2d
LQx0altY3CLGFYsd/Qanrt06TXiDyIclNJ/fID5DG6y7uMekw4nDYipw7iiWBpkw
M9AEiF8LCeQ/1ZdxWrdspBaniz//j+5pyj16QvIf+70F15yxlOaAi15PlblQViED
JquE8QSv1HOiSX45eRKskAubBKaDcgfHqjkZqXCpsksJgrJgUb1v6Pq183IL2ncG
N9rQmWX8oKamEYJzCrIP2TyvMW3LsA5DBw8F3tsnXz+rp1WC4iNayk+l5DEJqemk
s5StcWjIKizrXxpnNE519fxYy7rH3/Kct+FsDAyebOnw6Xf0uZFs0I+YmfZul/3A
AryrBtBSfYemez/y+aG6OvxcfB2cPSxuN+9xaVBe8vh+guLPaLnbm0zD7c/r/goI
7kYSyQt37TdKZRg+iIRYAi3kn8QY0TCmnv1utSQ9eZaNUaVaRRphbPoexK+Adw1t
GLP81A6757wDu5hORBeFmemg3dVK9tF/slsIue3ceKtg0SoyojhWWGKxAmdMvdZ/
AZR31B046XgH0v9u7HFXlM7LWSvaPm0uOdz751/L+ko+9OPfkT/uPAAGaQNm4+7x
9+MUDjUxFl44ffqRsROHST0kmhDSiSYn2aUfA9sGpB6afFJsmxU2Aaj2YrgO8xay
FoNKwOArIE77DhUassijp3qI2a+C40KPLQUbBzJnGc356nM+nBaZzStQr3Lsl4Vo
zNa0Ihmxfb5SwtPXA6S0etaeb5RO6RfY5kYyZYcL2hCFeHt5AyRh0JUoja8YSzhs
Z2AJd3znjag6ob33oHtCs1lD4GtWbY7vFtNeKH3Z//4yA2GfvkThqNPoL2lbpy3q
WoEtHUacG/IpPunFSW8T9QmA8MjL+1jkSzgMGed7Ogz14q37am+yVAcQFIMWL6uo
7p8BHwHVwxybb0wLzp31qndZc3BpAMMOQrxzRZnUNNagOtv9T2smH1XsFG13hBDO
OYUchU57YXJ5P3pib/OskGgjLoD8FUue4MCHXStB2diO6KIicVaBvbLWS9jIJ0ow
tgHgu26smAMpL6XEpNJCxF1U3tJ+i6/kB64yV1cLFTNedAJxEkFR6HzIC8Fu7JYY
f3CTcGQQPnkhbXI8x+OFByyvMc8wGqOnaiC1AY1tLiOe2KpI2v8YQv6LICnYrZ4E
ilA32HaLI1WFVy1HJN7jebD6gluiSfv1+RfnAIKUw3lavHjTSdm90YYy+YbePU1m
nKE6U2Lxq6vDyq1yCDamceKJ6r1YLIsiAfNTAdunwq6X/ZJueGyDM2WFqeXX5XZz
ArEapYI9WqE0o8l0NFpOBFQXemxSJjQFxrrIx7AR4C6awgexHIADpIR/yJmmQxNQ
LRIdxfZG5gmQoxTwi7w+uD1jVM+Lpc6SjFHCwy04wg6m/KRWUtKJjuYkUzOgorCE
wc1WCumagGO+Ppjf6q9dyB73DMkUscKLY4l6JFp8FmChwGzfQIdIfz+z6mc15EqT
gzjsr2kKb1iLCgdXNslpW6J67YG/UN6TSBlDdZM5fENXwxiuWzCAGfID3mYZMqeX
3DgLa97GIzG2DtkDioXleAokG9sz3hbgcK/awXD6wCO6VckWuCgISR3WMbvMgzpM
5/PdDNO7g3TVuxj20JrIsiS6WhZ5O2VmBo7KumhI4KREoP7zH2fZ4W06zEpDQJQ1
BBPMVnLeFNFXHQiMxusjraxIYH7fIJoiP5nDmQ+7ItjViiyat0XNv0WXq4hUuxA7
GZw0RB8cJ31J3KqFrFaKoI+zo+eGmvHS79bb7CH4nuu0+tZERszVzuM2cuvSBsw3
VO+8g7cN4iSHi0TupQh/qrf37PeU3SlJGtNtrd/tqHoIT7SJsO1GfpxlWkXn+/HX
+6vFs5dNlXGBIkwF4gMhOZiwS1qzfRoYvG9fjtCAAGzVmQL4uBsi05ogr/GihpE+
7HvPMYyKDi1d4KDAVyrphClBbBPXEAOpOg7w51dfF+00HW5esiX+PfuCTHBtNrJx
dFFmg2L3NjhN0btl0KxIAJ2aViYz4o37tXIBJ2o149xSOa4NtkmSjxY03xmWctna
zAZZL/gVFFk4mIVBrQcFjM/Ix5aYy9l1NHWqbt2P18/JmHFSdoEmCQQ0FwgH/wqA
xhc79p0cUIvJsbIh4Yn1iDbjSR8QqVrZ5I1WgE+AeEdauZc4aQmf1rbZl91i+JO+
SOzAX1SxzcYw5AavHincz51QpcRLTL0wz2s3KLPf5rZlDVHk3H4jvgfG4npzESwL
eEXH6eFgX4JP6j7v4I0i3PcDy5Ni4BpGlZ6TrqAaxNubNIATlx+7pkHRRlH8/pMQ
/6ZhIMhgTaUoKNWPWgGyIYyzl/Vz5+l7Aaqp3WDljB/cpOT4EzJrwTSZsRo+EitJ
LgmNWBS3sPIXIteIylp5O5t13GvH0JDNZWPKTsQ/tDuhBkfEzBhIJsNx+ZFrtreU
rEFI8JcMTNRWSdL3g1s6KAC1EyFOMUo0dCgB9rnSt5LUijIYeJU4OILbsWW2hX9u
nUutuu0EDnTw0rUL7lWJXl4TV4DJdmP4wZL5L4BQtUAyJ01v+noqnHRaCbGOMwO7
5+HHImNTuHkryMlyGAa8KcUxsIO9SGC8LLQp7stbV5cxk1cFn2Apc2uYWC7SA6Mw
TbueDhAvWiLckHx9esZSrgd41iNJtrIMbPSz8nsC+AA1lOz5oHkxR/3QqgWWFPYb
1Ve1Qm9rKX/oofBjMqXkC/0JcHGR2h9HelnDDdZiylyqX4tl33AVzYe+G9J5UykR
2QZVL7Ph1ESwpz+4DqFzfboEinRcYxXSgNRbkz/PDyMInvaZMAo/QDH81ELzHAA4
XTlnsoQsbVjuuxGRu/EMgi0AQj4chNMrbc3NpePOVmtsAcRMrvnMBmjk+PeSWt13
7dR/XoYivqVwAfZDVz6C8dM2yr0cVza+GxW0JCmJ/K8jiZ/ovXb2aP/HryFqAC9b
yCCGQ07QOR73PVOfQB5E7lKxVhTvejW02O6KWC2CxO+DBm5qAybnNMxRPrSy0TSf
L6hFD8Qjdv4vM2+uFVl1ZeE4oDU/f+thUWMtLtFffCaxKbABwoGwfQPh2oSV/vVE
xxXfpD7CLakv+EiTdFnJuhY6YO3YXa5w0RU3nE6hr+i3SV0frLzIkrWRVc7gSCUd
d5IPZ2asg6Pmbm1RWuPSFIrJ52qOJxlBmdFNb7luX3iML0PNHM46QqORoIObzlJj
MH7kqLgsrZR6PcU1E54K6GGuzDCbEC1AswZRApWTdQ8ibXCGvYzGQOHhJMv/1fPM
8DMISrtH7AP3swm4NOtSnsSrRrK+NR4P2H31ZlEpJ0HadrPS/Ppw9L5i+diGtwFE
0V0ZLcSMUnkqnf3y9HcxzCD63GB+7LeQSZsCr8WnPl0yX5tEEvzUH7z/DB1Pr6HV
/exqhqa/mEJAk57Nr3kfWSegIDff/p51scz47CKFKK19P6tPTK+R9FvS8isQGDV8
hRQ6RFh2VPVCnH6X0j24azX0TVFGPoud074AkKTc4os4omFQQFRgH0m/nvIH2LaM
qZWH25VKKV/0IPfQgLc9kYE7qg+fjGAr2MObs0u6wC5lrPYaCMqFRgdEEsbPpfeZ
mO1M9UqcdMv5nRn7wW2GFmdmfASoWMEZHR/8x7GTEIpyUkHizfOw6rQokA7eGaIz
3TfPh1JP2ARnkfivWGArftZetX9uoL5Q4WtHz1GC8DRyetLPdSw74D18bDgh9HLc
Rsmk3uahw+/AgAgAxq3FvimKTQ4brFaBP7Am1e8i/YDZyu5ofY94UcyVkJyS/hyK
OCu+YRqHzco/LtDCbzbZOVYVQ4QlrVnzyj3ForZs8v/Bf69MVBBXtyuvq+3OUvmx
qAoi1TFwiFk4nVG6veJ+8hsY1cdBbFVlWAizodwmSWkTAenpAB5d4ptRG5ogpYRU
oijdJ6hCCt740TmYaGqPoUBngZiS2nUVv9SOEVf7IV08TyeKItexVY9NRbMJbAW/
umtIo64wUD5hNl5VOYXPUItREDZURXqE/LtRDrW+PkENZj2x3wuWDClzr2k9bM73
/U57THvH2RIVkQPbQs+OukEEvdPaNYdztYTNK+0f5ML5Ha37SgyG0JS1xaTwwLUa
fmnvGq4WeVN9YdekjnhwBRa+54efwLF3Td0IrrMXwNxxGh/KRJWmR/riBZdJ8i7+
bLEanh4w8nrbdrHVY35ylQM5Jp1fZPLhBnfPYKb+dp7v0x+5CR9gQurpWzRYrB94
W8jH5r5N9wBxFD81M54dbn039sgYtLBEFUtX9Q5j4+DdDO87Xlytnflc1vCPZ1c6
ra66hQNr8A7M4kCDa2nIJE3kdjo/FUQ/S/2BZQ+G/fy3gip/OoF/MGb5SBqCV3A/
25TxEQyumBnzE68GJjkca+pJ33uVB8oRB7dlRAObvCW3fmvNEDzzExx4BwdY1XA+
9oorkNowBC2R9JFbMUVDD7K3ahr8wS8XHdSgrn/apm2fVw9qaXje71POP6uvbYb3
7UmdDvCWa+hwTPfJfJY94cUN5HxUWGf1/7ESj6p78AzA2lDWpqqDd6hwQQXn8VzM
If7KFbtbIUvDkrgGBkxMsjINonxrdS/wY5xmQ7VwvVQvxYGAbxdPd6QivTiyViZT
i+fJaEu1QB4zr5CCYvq3dwZgajeiXVUHM/ly3yAkaPDSSO6De6UFZXj/NAXuI4xh
NrqF5JjJs0UfcNdsVk7SOTEQoziDQsmKjf64CQJ528pEcKqH5LnUkqO+r8rtrWdN
VkVPCpQ+lhOqnGB5q+pzCj1Y0nxVe+L75HgYapYSDmAFJimCeAEeqiLIGZYSp2Ue
/yUlYGXiyo5/vDBC7+QjNO6lmdBa9RvsFVfptgXIugIWgWNtpozTLK75zDCFCF/K
uLpywhhoK8shoFFbMWk1p2osF49/QIw/XKN6k63PCZRkSvwqiSJA+gWSZ436t2L2
eqt9jbShgclwLxHWXN7t4JdoumH2FfVmtH42pq1pFu3fRAwjbilV+HG2tNfz94I5
5eqFfgDr+E2lXxrh6mdEZHnu6EKccBdFlmjEiVfBlct4J6pusYaX0n19vhzZQ8x3
M8ER/a5GXSC1bsUjwiG3vpsDRdzcp401lvLZ+0BrGx0vS2IGb5nyNXibTNzlsNz/
uzN1L5WMtvFGTcoQDVASF9vC/6IhvHMIGw1li6yz7+0weRXrpqCl9jWTCZCXVqzG
XDAxeXFh6+01XrT8W8TLZAYJX2S4wTg0TfaWf3t4r0k/bCKSHZp3+nItIfxj1LvI
JVlTjgko60IQvsy+WU6lEtYoTZwng05zwotdfbU0hMEXfws9iNQON7Pzg7w9qbbO
JR5FXL9JqPup++TGOIBHe5J1YQqTHVWahEx5i0pdLYbZYmeIvL+n3jefyfmGI3Up
rX+g3N8szDJMuhVCHz2P5eTv1xRiADymLA/1/K1uCjJD6zi5X4wCbZXxHIDcGCJV
jWXSKmcgYiGZf6kk3j9cno6DenkbwvSGgorPXYnOywmgp7BuKwYH6vm1GKCT3LHm
Dyc+ht7KJeCLz/XJMYL5YuZgkhz+0gbna9J+frnG3D7tXNcmPllLOOL478eMtjuO
dDvinpvj91+dtAm1S2LlWBtO+UIEyoH/kMMOnqZymqhrxR3Do7g+Cr052Gi15Y52
kfmBfMxciorQeQsMuJFxPWwsdpQGtQNW0fyuoQHV5k682/iViks2zYuVMSxBuuPg
tvM8dv99vJlXsIRBpIDVeAnCevfRr6uyUnwt5dH83725jywYCf2Lg955gAXJWliX
`pragma protect end_protected
