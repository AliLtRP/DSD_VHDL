// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:33:06 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
nSA/zAaCFfRFp5lx6a4jKtgThC0mQVy41DB3maoSfHXKWqKeMKp6bCdNToX/3x8L
53mHXzTJQ+LPZnx8BX4Jwizr5V1JImmLAdI7wXVgS9zhBq22Z++k74IIvKKiltrx
27yhrmoUGu0hXFtGFsknKTLDNRJMmGarb3f9QHAFysI=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 12176)
HskkO+lnosZha42twtJN7M1sQ2JchKUUjGW6wxI7HbkK/mKouIOqJQITvyoP1xII
k+HCd2HtUIb5Hs8vTVOG6cHM24jii5VGRiUTf8bQnxwNCivpTeCC9ak4TJemEgZS
Oy6KguyN2436rxkb0PdlM64HIMGBF+uEAwmvB6MXPFwQKE2nbMEUzed8C2uKEfmp
HOKQB4wEFdGGwIPLdrZGtYGoJMnkfoawu4cHNGJGo5MkKdTJeM6uU6J5X95fH9gP
TytLXD6H3kgnp+nkVZvqE5tjBt61onULpGXJuHsu1iE/2VtFIbRBLAJZLvzfT0ge
MHgy9LXd549FxLQnS42xinhWUSBHjyoDvLgeQCqB9IVufgxvmy2AneIQa5Ch5pOp
bl4W6CImjV3OBqTAjT4e3C8ej0ZBeDOBCfMfKXIEakoOFb+qMWUUz6CkttwRu1af
vhyJZUYIg6HmvEtPI7PVIZSd4SOABI8KDZSK1zVrKJGLviiLlroaa+VroulnfDZ0
J40LOi3wgyFmcGYc7B1VeOh0J32+SisSeqkg9uE13oPldIOA7pklxTQhRQ/MSYv8
msxdUNuLHQm/RXYair1Tw3MVddRRfBCQ7/ZPH17PW/7uEk/EHACySBIk/LUuyCwl
3N0Av+ozRy99rjLsezpjMIhtfbtPr33ppwGxOCY0u8Y+CR94ggHFV3qV9amk1J2p
+A9uPD9EgDhJaG0KgKeibJaDk45/B9KFHtTaDSBX9cC6R+Ssoaza0+6R0xjRf/sZ
k7WAuzMYGdJ2+nBizAf27TO5baeNSsTW/kORAZ2imVlBkF90FjyJWuV5PzN5GTEz
lozENqpbICQYMMkZinbhBfdLqyMcqIursBNogHpMyiFUsFO0JpHgdZCeLcCLexY4
DcnA5QvCPZ/93GCYW8gJmqaxKtzgL14MWw5B4Di2WVAiLlSmmy6FbBudlPNSrDqd
COw1ajp9nUAb1D1XuRqflYh898Tt7gt8V+ltWdHUWJttGBJaRzLW0tk4p0uKJenS
8T8F52DarX6Mzrd3FRubzHkkK9gQqjVkj7Jhn0uFGLZe/meZn7Bv+IXxnlOZEpZ/
bwmfCm1vaaqEyctBrMN+TXtYeJ5Sa3XVUx/GUXPTIx9R1PIbQuq8lt7OorkGvula
y/F3COT/inha1wMpCDZ1cYNWyJCaXpddUoeQgPc/Xqjanb0RCLxJRWdbvuLqVh6o
gAAobwYFiE/mHBPTIjiPMV96xphBdJzgmS2B6SrwParB0T9OWWuZ5nWP1NezBe7u
s4GcT3E7mtaNaD6eW9XjPMpWQd7l73wzgtZHPOhN0y2mPNR0o2JU5t0w48Azucaj
X/KE87wnsj4J+llG/kQ7GknvD1DEaygaFnhzbzxFmsAJNoIYXTWcq6rLiquUTMB2
8jyRLHhfJ2YG2uO0APGYUpVekTUW2pm/yz45jPx0aIYNzh5sFXyZkkymjwrS5zkH
3wTPKQ4ixdr3dxOlXS4Q/QyG+r8qN/dx92dmK8sA1eB2X7WViyabTYs5iQqhAdUs
Zp7qwIad0g94ZjfadxwyWPS2Tz4l3zZ3NViqsdDfGD3vY8fIgk5/omGbdb9xglkL
KRn+lDUE46j5iG3vsoCVQLP7KWdZR1L7IC4oz5RLYkKr1Bk90qRUMPe0lttMY9u+
ENdTouMgNanv+hqpjdnUAXKtIdWuH0ZJPCxm0RYSsJyrHkMI9U5HVCf1zXmAMzal
hQNAUnf48+/xUO65eLGzwQhy56qTv33QEn/spUkSMBrA6/zZCBQ/F0+ZhfboYkjG
w3SkwnLMoRToqSDtLW4HA/njtLDZq1zxCVfN3FU3q9hsQW+wm3X5ZsjqoK6NMFDk
PV/CTt3ql5Mw6Esx5eCxz3fQ21rKvNocR8IRY46a1JANspONgKBow6cDD6fBVlxu
G/CrJLXWOTUDkXaLnp0gnPdGs0btQp0ICieP2lXsYmXRLu8NMNrlq8IIPP7znKFD
TVaNbvP7dBhf7+bzWdc6ompTiDAFsziPhFuwQOFkolVdc85YXQX9OGBesCEcwDMb
Xs281QTsjrpVOSHOaNzN7i9r3oCsEkb75xpOFMxkw0i3IqDHyLVT88HJYvYU/AWP
Hi/lK9haLqZ6lqqA4r/MFkGZDjCoOVH2HoAU2xMVig+QB0u9YL44KRxgaDug7z4q
vsv5DqHgnao8+1ZQRAcR8Lr7X5gV8p0oZ04TDHUoZHSVXGYf3VWymuJbLs+KVPnr
HIEuFXQUtmGjTuOGzXnV3FvpCcCpPhoAK+CEFRNhgxYrmFZhr5bzYPe0pYmE3bjV
f1TBvtQtDMKxrt8/adYI97dB3qaPxQQ29xQO29DG6dzTJCKkJG0WlTEBfhsTDmDO
n74/Ddv5/EpX5L+FExMLzChTrpPLadNKYKgPMpteUYQ3zor2m0KysXd8yFP+jhTu
8mIReDx+3DMDTjVhA5NRQXXERuIXbvvDV45jrRyKA9tXMaJg/a1q3Dh3pNK8MRWO
OdyqMnJhb/0ai/r0MAxKO4ex10kge9M/Q/+13wyZiaVtF7caCuiBDEJIjBKgIuDV
Vpm4VHGQFaGv7Lr9xJo5Eh/eF9IKRGykEIOBG9KB9zFYiB30YUg7REGo4Gtr4Wog
YjjQUikOIATMf1q3NMrdIG//DY3bdd5iMEPoSlq3csbK3QpLHezsWn5v1DNWxaCS
HoalhRiLXn5upsNV7O2iahF1aVqwt+4UDg/LWahvsMxm3bXIcgXXLFrkA5t68p6R
f6ClYqhMb3vLB8GLZ33KhZAv3TpHc6mFoCYxZmk4vn9dIFeDgt8eBvxz+U+ievtZ
ByGTp4ur9haMWXQpQgAQo9xCpx1uxlTVdZvm2dkENuvrdMn2hVI0XXRSTCm+/KMf
UXt+GWpgcbSMg7Kt9XBl4frlJkXBiH8vCl9eU4ei++w4ZVQUzE8P83uBIvUWjUf9
6b8a+I6mYzE6OCX53hoqZ1IQkqGaDYay9n5VLHvYUcTbWdXCU/5R6mzy3eBw8kCS
wfwfJDybvrtsF91VXrrHilvDqnr+RWZZz9J/eGt2NUOotkZEy6wc0wkWB8kITBQB
lZYg7+W5NJeg/tzngVqLssfCBy0CTOo19kigWRCc9zWPdt0ooW06istFcEdbmRLs
mdUc2cx/5jGLuEElsWuppzEJVMKO2UXHyJbuQqlw+3asB9/ilWsg8GIUd5kT1Hlq
G9/VkkWWODZSNSrbV7fXt0/v9pfOzuHGc3tdg4z680JEVUt1XM8LSixx+L8ks8AZ
0cV7IYa4ZeETZrduB/TVslIZwuCoiNA5+EdTIfCVIaKcIlTQoNPZwl98v8fm9dsn
GJhRY6JQ8mYM6u5KX7yoVApaDwIJT6DVYBGDAtCRbUA/IK+BeS8QZx6CK7fNvss8
oGIZ5E9LPejmB26HnESgnk24bp2emwbEjTFUfEDQMHgWglPFEP93fgc6D75KC42a
rVAAy2uvKtN4OqbCrDNfMhSco14S5rnjkF5vvibdLM2hVNBSfTlbi8ZG9o0G8X9/
nFFGTeWSuhBlpltlc7K2Wyed8EmaVBozGp9DikfX24zl1eZm4x2WteM/hBYF2NZJ
lm7edfLC8Cjorh3UeUr9elHjUYN1UozK4r7INLtq/dZaqJ/EJ82eHvny0DUTHVBx
3fRJrUSvSrw9MNyhpUl4RW7KeAuTfvb7PDaFnIxgbz87MIUyfOsmCnuBsnM+xyPi
36Oj4Vt37jWwG0nu5VknZp+DCPploT1sejYl/pr4IbGi6bsGWRYhplkqSN1uFiTy
AC3XF8T1vVbxW1n+5gC8+M/A9BDvtlyfGFmlmvPUOthqeUgn1kVl3L0w/WXgPHR0
ZttGwEXnQWLcW6TSRUSk3Th1P3E6mOBAParZbtMOtubQ67Jl5RuG96GwbfjD9ZVy
2koYyL1qk1rbsXF7dgoH79p98eotkZj6h3pAX0Ik2fBWwP4zgFMrAUxXv5cJIhSc
prRhMzOaEgpDQ8eLDII3w2nTE43umrgxamAEs4JRiGA1yadu8jS76iQzcI0O3LRR
X1IcYnAjBxDyo3wZTUZcG+smhk0ATX/koHwkeVgQDKujzFBWE23mDRg1dvJ9oJHK
5omk0AWGke53jRsq3m3eNK+PGmsPXVRaX1OHFjsuURJD69rUTCV9Uxq3r+n7F7s6
ojSGtlekam5jjeotgUYtp+KqGGNUvVhkNA4eMmJv7BYLhg14ObwX/gT3rfadrS2L
1AicOlAWTgLW2GWLtmvg0lSKKB9+RKwWyirs4AHDVfRBrjqZHQsbi8yJHD6KMRxk
sXj+a1PvvNaBFmKyWaFDjnb6C7OsS2P5hHU1ySiVSU8I6NcUr2HEheAaRsjzy2cW
wy10rnF6UfCp2HgjRnXWmj7OdJ8XxVElUHgRPDhbCUsuxWHDhhyNzQotQrtr26Ne
YIsTgEw1Nqm7TIC5RGTHRE7srJPnSdR352BIgEJNBTXupsFuLy/8iU4npA+QlLFw
HaSOYrqVJhThT2fJZ8ayyzGmW4AE5TpROwqoyK6kTHIi/Pi3xuRPOBY+bvYYAEQl
L/wiuBI6PSrNZ9iGZuCwxlkToqmB8BOf53tD1uJI5yLuvQX6h12x+dqYlawFtJGM
QvIrX6nZskLTxtFRPgcrOrxal4/2tr6W31fJ05olCYotfXD5ftDLndvVO1idzz5Q
y2HU5K8QTYUFGGCP0qVm5bL27NQN0e0gp2WjeiZWk/Y6NPMwjH2XxPKHb8RCi/MY
5mAwnc1B2GfN8Oa/RFV/NzBBh0cBrquitrRYxvKkFs8WQN+AT+57RwDYCiu1L597
/kCspJj10kZOnfbt2Mu/8w3McFgu4BEXZ4k+iZY+eb7oim9Cdl1sMOxtN6Mt7YyN
IzZK8PK912HNoKAh09H5WgbkqArEAbNJtc2f98OWfjFg/1oPSeKLNWnB/Ri6aXyb
nml/sEhrFB5iCg0NL1+APwxyj3JhIvyrvjI8avi3NdqughT3zx74roHHVDIgSa8+
coKbFP0Xx25NuaKQeZ3bs38QKpp3g1VXK0hODV3twQ3Auc3QQTPlxQVumTwOlAhZ
yxZbTEAblCISDRbNSFwBwhWTyXVro3WCFMDS/4eRgbDF71HZX6HSnkojAbJMSeu/
z5Mq/9exuiY1g0vS9ZxcZx3jlem556SxGia6XTBVJGUdRdSvALtSSHd6HFIE7Yt+
OZFX4zHHTiDI1UJ+CZNHpuvwtWe5iMNvnEfZQA0ljwiw4uW01n/8i1ttkkUCQR5A
J8+xUnSVfj/70qMQwQdGq7tydXtGXqBdD4rBsUiA+FlAgPwTYCJS7FromJAqq4vH
KfuvWlL8aCIl8x/DhQlAwwCmq0vja/BdWz9Jm5M20uJAvWShAXpgUh3+ur6BPStr
SE+6wqH6QLt61dDz8GfT9tZwDuunfQ2t4sHV/fs8aKzdg91tOgcQlNJZtP7jvsSW
MOZwirTOo9eHhTdgE0c3L+2UOcxTn9nG0J5B18jtjZVJHxeM+dDxoSdkmssCBn53
zHI/xaSibKYI+R4q8LY+2Lde6iYvM+qhmFZkAR6vU+y5UGtu3gPR1ueM4WXUs2Bt
4H2eK0AhEbqSIhOpb1d+9sqlGHrWT51annk5JEEOONq7ipcXW/df6sQW+2uXyIpo
ugdhtuiAolXTUjt/WnOztuJ5UY0hD3x6NASoeF90CGbpG2jd7V25FhxmWThjhHLA
fc8A9SvMBGW27dtEWSEzeK1MbFoVFZKPPaxUZGe4LNIum5uvOzruKG0kOBNE6rU8
3lbEJ9474y+gkUq83IqXuMsFOgbBTLbQyNC7uqXz7B3ArAfH9LtI1QORyxufYmOE
L2PpSL2Pq3qcasMpAa2oeNXuBHzRCzOmAtqDjZtSTNTAdMbs0oDju2dPg0+SHjr3
sZWXPWUX6gU/hIo9Eh/OD8eJCXoM1ECj9tU9P5GgLDK03T/mipUGqJjIEV4ei57k
VFcervMREtBwHUJz+eS8A3j9bfcHznmkMyhhs/KbG4q3AaoCWRsBUd7J99ODxmU3
rc8h19BkKGxzxGrRI1R6goqle4Hhy4F8gE+FX8EP5NlyOQyMFgGgFPphNPf3sMSR
s5Y5s0vr4k23Bom0eC6iNfdowOQ1XG0Lvjb3Tn4zN68scpJ2lpp5Uu61F58wENHV
7FlPJGzZgxNnZfUqqXZT9Zy0LnV2eTIrXKy07n8eoqQ2hWQrnMAh6nxDeXy5a3SN
9w+qVmQ7jUG8PcKL6NUpifXzxjJSnekm8XsYr0VZB9vMlkUY3URIxPgt7TkPfjzJ
XpKkfVhEnUP5q1oofu8x7XGdNxXcJj8XSQvF27TwRNDFygFVjci5oVRTV00OVS+m
R45PE39JuDHY/8UHRTaL7FYr4GfLljVekFGiObzdl9OQcxVSdc+tHdWaRqzpDPZU
N9KJFO/d+ejLI9ByIhpQ6leIh5DWZSBWd6YDj8YiV+db5EfibEv2/Mvd1VdeXfok
oiQZBgo+kvYztjvEWCevsAM2VjqsdtE3+7E9fkL+VBKezNXOxOX+R8Kpb+3sgkaq
AICAjIj3WujYZO/awJWcZsPjsI3463VU0L/BjIqj+JWyVjwjGj9uie8ma/6Xh7cE
3eM3/yXrgfcuVqZD8y18wTxUIvWVbUGUizVqEDHyuyWSQH3Hi0Q9uUd9iLuzuEhl
JkYZ2hj3JOrUECDO1FS98As6VrdDvJfXxOLh1LMdLZOGGNxkpo6FSGSftCCMWS0x
opKBKw858EG4k+NFvcEfroQBCl1KRGC4vbZJ4JHzwOsH7pLjvMdjr880hz9u3zlt
x5tqc8RAL+BTxGYMxEbWwv3BzEhhk8vvJYm3d6YzS5vvwjSI2S/HdOfQ8byvK3H9
bEAdPM/8hiA27aeD1dDwN9B4cERIAECZOa0gRtdQr0+lfc3Kw+oojH5YmDhYCehX
TgZhisIbyS4Oe9+rlWL2Z/sI3njg108pI0nAbLLL1Zw2Mq0UBsAw77hjK2gP14F6
ufd7PI4oFDYQKTN3V9Y3xZf1cnAdie/e+BTGlxb/mt4Q92zRkDIqTqKMxyW2GMc3
oqlCbOSdeEjLX+l76LMacbRg8T/YSTcRQ2eV9vaKlZyFTshCOFoRJPjiD/Hv53sH
gtRSj8JjCEWIV3/uuz6EXQ0WfuD0Ne6rOUgU6WBhDxcSeens002xNy8EWlshmtVD
9sVlDDV6mtaz3WIgQu5UFPg/RnggcVVWwL7uJ1Bd9TmDhyFO+N4bw8KlcROxaBwJ
qPpocnuQb8gAo0yUJLUyg60pcsgTcRqoZmsdOZ3VLJtNtAaXuAMbeAlKqa7qkUDt
hoyYmq2d2Z2JD9imIav3yFzhFb/fPGZoYdn8l+8pcdcGnzciL7bk/Cp0iNzr6KTb
sdJX0LViiBveAbEwyMGWSi644yXAuZqgYda6RIYVhYhe7RUtKH3AA57hbFqOyvGl
O8+H3aa3DlIFK1vReW+iTSPrwRNSloVsD0GEdySQQ9QV56iNByL0/Q5X/FNMsjLh
Z0vUnEhJxhKRYX29jehcMBpUi4TU3e0nUz78ukb0sSV1/Eq7NeL7/eqnxLe1F9uV
HskB1AGq/1FDI2isxaUSugB+KOYSTFPdixUwfLoNE8iFkPNGWFd5ZRXHL2jYLBcY
2+MPZNT0pxAACNOxmidn0xPT/W9CNVVTOCEYH9GaR2BgJtPIaci2P+EgrYsS9Xn1
byi19qSSuhZYHlE8D2YVqH7Gs/R/rQqHgDRoa8Tdtdu9Zy6jyEUgXOJtz7D2CVwo
CKoZG7+4M9PQpMsGBbCbNcW0/UNTPyAksxZGRDYK7mD+sf0tece8+4fr2M591AgF
0IxBh38N6ip6QahFiyCBCdH2pWMbF69xiYPiM9YQg5A6mvhF9L50JyiQtWiW4yw+
a+4XKAzZxR5w5O2AI52gw9i02pprNkiJfuaUsqaVPmIhL3pslCghfBUs6OA+LNAW
Dff/9RY7qHwyN9+tBZ3zw259r3R47xpVQx7NtAQUBptN42GHU3bDLFqwKW+A/A9I
5m+8ny6C3TBmT19G0Nn2G1Pgwoh/cUx8iGEZwnmFjTQ++YiLZ9I9eYo7zC7f5Gt8
xqXYNfnx3MvNH6THiCplQE49S1ZRL7pa53awamp886D6lbYS802Li4gjLmrrljVX
/H8VUgR7nTWhHpgIhfvA6fbmlK4pRRsHjmY9TDHqSwUtA9aIC90Du3C47rDxYH+x
RzAUluFsIRLYpLSCjDIwJK4C4MXBWf6Lu7Jrz5O7EPd8tZrUUGnBrYWV1ztalPKf
DY4LFBmAy4p+/SIzcxwZJRpSuRWaf74zXo5xFZRo/159tXU1M+kIpcEhglWmvErf
1VT62F3jfmNadDONPj358sPxiVqM6sz1ehrHimrzvN3pC3xDQpo98FXGn46VMIIq
KmVsAPqtBwN/zwLIPaSwzz3HB85JDCWF7AkeCrlInEM3gfu0NjzRvcmFpAsHsbRN
mhhdNOW7YOOtC0J72MKi2CHgMeDaG4j569cMx9BzwXMy5yTPSFz72pW/+rOyyUNh
ntVkwnmtD54YNH9hpP8q6CdYVBfPRLBl11w6LONUTltFqUWMHwLmIiukTtBLxnp/
ME0p/PVqgV9iZuWr/PnXL/VRljBXUuQHmENYINfRn8MEemvODhNlHoFdGQPRM0dV
YfDEAQTaew0afL8khsS/cEtOC7AI6gt+XOlK7oZyKp77P46zmjM445rHmbUXM3yw
0kP9MMpGaXCSRhrFvU8yx3tnQYz9RYntza4/Xydg/meslFTQ3HpG3GZLk+1gzMgN
PPKtoSGo7viKDx2qXM+wFgYBXOSCOqwpMMVsejPNyaPmG5yLFlltj1Xa01HnNe9h
xovuyzTPxnk2e5/dHYJOvWLRdyTIIS6iTYdtaBRKuY3YTtcik/xMI0E9Z15tnrw3
cNbIX3Q0lHWIlYzdXkG+zTyaztoXThqgvORt3BEAUxQdrNP30nBFH1Zw9EM0ztzR
MZKW9aGdGfza+cb7KdxvuIVooCEhfrF3ozHJTWwzNWOoepNCfyK+dYz6CSFAHvUT
HTcqVtX4xDUZFeIHpQoVh6/4DCYklQBsis9/y3/HwSd+7HZBqZC8EVOlROjX57IQ
aZ6ucRrLLv8blRSFYTYRRlBFX9y+HXC5ba2dJQ1IIVkMkGawGV28FQVrdob6gM8i
8iu6pt9jDYeiLJf5ISJANFSGAhI7LsgBUbyoS15rx+mYSJZQlRQ6XcLGdo/o8t1S
Rs71ma+X358NXKxohA2smymAIuZvFcbdUO02yJkG+kpf/5rAMH8mHwBv9Ger4Ocv
6varYTTkvh5t/Em6Jm6h6ud5zXbGjbQepbTzAoTM/qLn+ZoJzwrwLbJiUOVWzy64
i4p9fN63OWQ1qTQpZapYX8UK0zDkdDnvOTX0FksTdhX8Szs1lZScix0roSBeiSLE
oHdaXNCElfEjTu2241xodScesiWedKj+ly1qWu5nM7qVvh6iYBnbsRo+MComPgsM
GkZQIa5qgK/XF2vWxLF51kkEFMmLuM2kqOyYrGbC7ScmkYegVpi/SmiEcFvzDpmb
xzKjf38EYGJjFGRM51yJRASnH5axkWQ3Id+8K3J9wUoDx5wX6171QNJlLRj7th2m
0U2jM0Z8UbPeXOtN7ogIY6JxRK0SG+RKfIGg10kHjceq9Mck8HdIZbPKh6mOIgD4
XfdkJOkfOzgSCS+vlzShaV4EDtlEw+XSxgAgc89ix+ru+/aHCLrxwTCNG88MU4cF
fjK2EU9lvqipOQWJE7yG7pK1dLESwy/e5Sen99nrdsjxjwDQ1hUSFpmQJi0XvT/j
jQORKbWukuO/mO2LYOlEQ1SYdROG+nocosgRwxeZl8KjqgD9JWcXq39QTBigeT7X
NjDix5zrS8y93Kty1JAaGEXSF36HNXcRKT2zFFex5j7yR7vbYGKuMZKSD4lahK6l
yN9yfH6uf4+qq7R8gKd9uT+vErwmFFQ+Pyh841tzLHvrOEbZAm03d5k8lJE6jAkw
kchXAN7CB7GUrbC4Tyub0vqDLdTJJTlPlKRvMHm1AQo/KRtO8JIo5fKwhAoLiFyW
Sg7fOqJb1dczVnfslD+ANNyT/xmB/2SL7b8ms66caoqatA9Q99lTyHsbUTNgyBGK
gIdrPb5KE2lbJG/Z7hrJs0SuW8RkDE3neYDFbJISGd02Inq5j6exQXt+XU6K6RUp
IAIKh2IgN5+KrlsXJSffgMkWB5tHj0WrPUNpdjC6mlr2jhULIVqlHmbwXDceLSL5
n2bV/MJGvSCHCO+5XsXmKnisSxi5TPFQBpu+NVp2WAbX3YuG8fku35j5mIhIEGtg
2cHhZKtHk3lK2HT/rhFNQ2/Y7/5mWL32VhQoNJTKSFYVep23y1/XnDkY5YFDP8Gi
wI4QSQ4ygkn3pSdAbU+yjgVAVLwg9kv7vfjQ/3j1UXbOjl339cU1KrK5eslu3NbC
z7sW/fhd+rXNiwgZZVKutQPD/iqpwOotRBFlB7mMO/mp0xv/VjXPOr+9R52yijQB
uHnKvmkmnVSrYrs1Ao+WGk4QSmKDu8MquniyIibrzRjxlWnS0G0NVn9CIfSanhps
f+uhBK11ainoYI0SG6gTAI4ttJ20K1Zifz+E82VTAIZ9cCOmTFGEmYkTbxoLvkLp
2gnGjaL04+NizBZzS2ufGfkFsJfBtFAfmk/w7Mwp1Dx1encxOnRnXyyVq18J5pAo
f1FmZCohPNPpNa9sXlIFUw9I3aAL/BFCSrzHPe7DXOK81qP2Wa5kE58MklIgyLEe
GJjcDJhxfFsXKabzugAOX86tx+fkQxN1CFRB6+xLJB69pTaDDsPFA9A1epMyXrP2
BT6WJ29RMtWooltXBUtVHyr1K0yfwSVIVQlCtomalWeQn91Fjg1ZFSqNc/LiWeUp
pMUXZxLeJ1wC3xMkcuq0lkVXmHr++pynTWxFi+GnixlZ0Dn+WxxXkvEC3+SGUvVr
jVAM1//PKoUHXB37WpjI03XmsErsWY/9paoioTjwJjjfe7O8r2W4gWUNjp0tp5Uj
1GYbfzqUjGFm1TS+pAv8qnoSWOjpag/7P75FS63AGohbk1UhkrGzO0R79u6BwvJW
sUNVnqDB+3rep9/CtM77+wFtDpVmUMLwk/8cpeGLFqIS42gp2XuYTBqQy5fIYJ1g
QEj8IYlHD1IIqApyvl19+AakWNkDuRjRR+Zw9SUAbaaUOO9+PwtVjaCpO7OBWjzE
3wTUFZqE8QawUvSQrKwzOelI5ZirRMm8nQooHpzjpUIncPlfqqIfNxR13dJw+SDB
DAUjQbQSibM7WW3f19j0nEJEHn5AYdrMm6HOLbVWOpgvZUKswEp20PirOQAjrl0Z
48n+GBYljx2I3xhIpmhVPuwYSeTGS6G2nqTAckHj5aWwGOAw+ifQ4elEByLG6+rq
EovWWqWkeC4766M7iekiUc/m6qR0keyRhnnc0O7RImqYPB16ts42KM+G7kVvBj8E
zPbRrCb4gQJjGSPwLGqiBGqTMoRc66S1X8LcNQEAd9y4BlfQYOQc9qO7pY48j592
t8eNcflXf89tAzwh8jZSXpFqv1+DfZ9MIGzts4Cgw3c5w/V+riXYooXQKt3ggs3Y
cjshqVcsL29o1u6z7/JLn0vaikE4sQCXt43bUpUvIpXTMRz5z+bxVTAtXCTh3ek+
WJfiFzIHSU9u9a+zrdvLi+F42R0ZALz/0jNkBtGQeY3Mr4+Xts4N2nlRDTEuOG7o
sbnutvM1lHlUhgWhTxlYjd5/rlXKm9lyld/oDCG1P3FksEP536HWjOw2JU/Q1F8P
cPidYOtmmmX+mdzDWwKTeeT8p0jcqGVxcAlzkhM0wQm5dSPtbYvp7esBHifHpIRk
wyjm6JUc6QDAbkDhNV5DBsLhffTlVcwVGCVK1Fti1kkLwRPXLCnyoCz9On2QyaPg
Ph5OsE+qDDLhdbXpGC18TVDoysgmWATyPheBTQASL+o+3BtzvLlh5/iAZ0Kl+3MW
pXEGFfKk5nO/fH21mhSkiDFcb5P1s5rei1Wg74Q3ZNbtnXPyrtu5EMExDpFv8MhA
qE654yhymBNDahm+AmvzncoAhxt2bQD9TveDB4oNjVp/ZgY4nYS8hwWLBzVJgxPG
a6kIQ/sCd7KQmTEkKmTrEef6YoRWgjHr90NQcUYHNozid199tLTui9otY/xSMWge
GQL9sGQ3zm1zC+pEW8FwSvv1VFc6korWqYmHa3lSGc5srIVTKrly9xJssUJeAcTv
4/70UpU2nalr2CxASCAH7mbpmOrTITjOrr6+ZlMeVJ1qWzbhNgSRHOPjUOzqhET1
lZoFrhvGw9WmHkE3T72QZqnyxfv3qIcO9dS2h/LIkNc33Nz1GAsoE/Sx8TZaI6TB
p2qCOLxcGxxWPe/OjRECE37YJGXjA2YQdnZWv/Kjkp4KLbsQpRx+Y4XY/EV5QheJ
bYwYHEthHxgJvWIj9bAtvyPQjxr5p9M4dvM0TdsLAgisNGe4+aN4p1LRy4iNYGIc
aTcvcEIgAUPsrc8fGpZ24RiZQx3C8C6EGtTj/Jh1V4wS4znoKNmKbhbYjM4HTt7h
KFbgdCtEXiyb+1+sSV9/Yhy+nWJT4GIaermcgUduDNqWHbpYqDgjqwFGkjfdCY8S
Mky+0Ldkbjy9CkxehZfxR2lWfrr55++VDyH+mw+YmqKd3Yzlsf6uaFQ6sgezrov2
i9bclVxsheFQOox6Ofj4B21X1TmJke+EGfaly0hFO0QT35VzfjUF2uH79BeFCGkk
0/tHE0jYOklWrkqGl1KS7Dh/e5NOplusdUo3Cm41zTZaEGJvBi2a9NkZNOP5QfYr
CfZkck8eG+2ghP7Qxa8Mz38Pxy8wUW4mz5KRlMPxv1+5m/k8mtX7ecvGeE4HmRif
wQZGDd1yPdb4tlQogq9GrshxB+BxOtfkLk7uuMMDju/qsOq2kkiqiIusg+Be5N2c
wAteu7Hi222o7lK9bnKwtlGKooW8dDbUGxUPs+013Z3VbnxORadGp18w1m2iJuGd
2WSnpf/5cBxHjZ4wWeYGSJdPtvB9PAdXD50eEnrxchyRvS1nVSBUKFsDejV/3YQR
q+w/9qFeMvHQAysmCnzTxD272oPbaZOPXQrJcjRYT1s8u23iEtOT09IArK3VNRng
l5dtWd7I+agGV/yC8D5sOxdhT5GuvUfJY55bq3aIhjgCQ7Q01EFcjiUTLS0nza8v
k9wPnum0GjsaJUHmPjwHDc5hcC3kKT8rdkKLnLmreKEqbcYUte0+dQRs2+4F54M1
Rx41eSZR1xYdJLxUnJlhzQ63mU9OXpUOFGZXG493fzArMfJ5mcX4fxAWv6E/oEkk
arEhtZb4Xwr9sRrTaPzqGB+9rQJmc0uGucV903Nsqic4uTVDd4vDmyOYM5DMNeFS
FnxkfHcXGmfyWOxc3Vd/xLvhub+BC8Zo1BhiYXfVHgGnhYe7JX461hnb+wxUCcg/
fyukpuiNyo2Suaifg10cMYeCR6AnzyCinbvmBMNmFPb32VcwcZTtDhYscvpBwrNX
91Uch4Qj+2x076pqY7+OaRe781mpJ69AjKKIF3YSw8+3ulyoROhPWZrzHHteP+vr
U6jicWSVm1a5m124CMQ+xax0yJzQZiJ+Ns1XFkdBLuVyestJDYQfGs8Q0QdQSTko
dkiZ3p2yzs6WVsjWIN0uZJADoKLbHK0KMGL05xh6sZgvbvgK5nNuwZsnthiFLCi0
xL8QYkZF2Y6gVLLrUWRzzsbu8XE61thvy8rTBBIVCWi/oM5IAdCIXP9CYPTy6rux
lcLishiQuzg71t3IguJTqu8axZdFiWW0aS1D6zEt02iUO1etvl0ZASX+NN0VKMni
s4Wlifka6VMtL5J+yKepsT7Qn88pBxr6L0vQk1i9l1d6uTomFe9zIc0KA1qlS21G
EsjdC23qZ3e9Lp0nNvTkTfhoOv6n/7coyuw2mGlMRKqcNwL+PXsM1FaANZ0wxalx
mjwyvdZg80mhfXMkhEytrWk10sReVKk4muCbmkc6aGwgBPwkLnO/ls5oabraa5FJ
Z+iFs5UT4zU5alBrqqkL6/rxkbPtb9oYkArw4RoLIHx9PB0oeIcZaEl4l7/ohbfM
UvV82zXOYZ2L4XcFfihqSWtUDXSDO5aW7ryEZoCpWCcxjHffEbUnvgwA2R4qDt0u
Wt+FtvJHT4qa6qs5OC7jZSqpjlgyQcwH4a3xuaQL4MDpDA3Gs/7AoSf2HjrPE9Ip
hENSrvqVFKqE4awYTvJn45kFuP5iHAa2GCVY5C7gKYgTpMmvmrBNM0l/JmwOVSSU
DO8PBQrMZ5Jwnthp/I4BlMswbftIwea8ejT8oVhI27SgI9ajUU2fymt6ET7U2r3g
6uxFiXrVXWS5xSo68DT5Jqnf/89fHCETX1TNBjLOJA3Phl2S9UiUWNPGfd1lG7qE
7aTc7onmCDth1vV/4QGAQ/p2M3GaN4oUevD3zsw7Bjg+mE6Pj4pnS+AO2BElpTkr
nP1K3uq/jmGJYyV/51e5aptAkMukfpSBSZ2Y3OYDvLn1uTTEt+siOlmlHQ7vMzho
PqcanlD5YpvmQVG9yD1q3ET1lUEPTQGC5akgSNgudqHL1SzpSb9dwMUZpkGa/Nkt
eVT9ilko3hGmYQnAQVW52ALf6jC70Af14BOgJ+dCUZ1Oa2q3/fX7r5FuN6r5A4us
a7EMNofB3C090K6TkRgMVR63tVQhNrCs3hbjpG8kGdqkjwIyaL52IhrR6VD2AKfU
t+HtXPkwzRfV0t7/tmBbXSyqzlZZBVCZZYtbcnPWdl9EvGfWB+AMWzD1KeJRUeTd
mhpL9jHYjYu4IUo6+72KjQEvpH5CCEVipPld67S6m8DCXC/L0OZoAlLa550UXLDx
mNgMKxLEyLc0eAJRuuXN6rvHFNW8fbEI2siOxYlKY109aRy8ph5iTdCo2QevQVqf
eOZf2VfpDgWgqTA79GEhVQEkxX+bPCeTmns/XSkntOWaxrmnXGsdPRVKpZ2GQzp6
D+QGBPFdcIOfi9vlkfFDVa1ioMqr6Xbp3KtkzGmoUNl5YsSZL0R24Pkto3ZdWYXY
AScKxXgpyNYHxDMRmhL1tdectFpfYmOqHRhGKmdqIcyOSKamYaoXPgPI75Mtt8S4
rqjRCFRXPHllvuDg63E4Duv+TBhQutDkeI8YOaqm47kLlki98P1C6hu0XcBcqU2l
S3bNgAXru39dbSmRS2JARwKoUDMWzfwF4Wja2rGlnGdKIhYmuBX/9gJiNWOdR3nz
E0ki3Y3sIlugHQFv2ePgTsgbaqqSEbzOCgKSQAZrML4dc1ukGZ+6MwLNlJ5CFlaQ
dkiq/K8yagLwpj9h4+sadeM/02bBzjk5ofnI5m+ep2fFjVIc1tAom7rsZtKfM30V
s99wFbE7Q8C3gOuuCIzsgqk4hChV0Cko9vAwGjJ2NJbh0XVXZCGugOZioXVXe35q
MHtiNL+iTI0TqAwEytxnnuSwdi3r/nmN6QOzqpXJTrILOJKqPlD5VZv33N8pvxbZ
zduMuWAncnj6TndClUehlcaPsXwcGKF5IXoZniLRm1Fos44GrlwPguKHMSJC53xL
Av0lyjLEsVS3nB/uDnncG6u3Ht6qRogHwHsyDH6Zey7bKrJGBgiNOoIZwl/PuoJq
VFWDfwBoig70mElLw8ub0BEIWpPT8sWMZqOl40dsyTqMMLaJwUEubp2kRb9yvCXf
eplxeti0klqNLKyrYHohuo6CGVqz6TRCfThC2JH5bbncLYpc/9X2OCgX3S+bjGQU
vvKJtLV0URMSpKSBvib6Km8eH1Z6ezatXZKlxB6tPzdS6l+JtXOjRYoAITEMLRPc
79+QZaV3EcW61k6bJ2aGd2yHzIWNVypihA8ttVVRvPJfv9K+iiYoAkh7NukqsRLn
GJn1ZXt/R+5nRJXFza9gkl8pR2MGlzRAeY/dj/VY0LkG62QWgoCy+wyJD0ojCXx6
PJZP/ENsObbZEsFvxgxIgIwuU0Nvy90LgKsF1a9iD6jvzgQeovOd9Tkp5iGdoCrP
Gg4Fw6K9vxzWggMZjqoDP/sJfYpAhxjDftmbdKew3EmOzUaMdlBk0HXEy5a0pGTx
xS5K8gZ4c6m+3T22B34H+XvOqFZICuWgyAQiyU/2sdW+SSy14GfbV4FvdJIjDn1d
fDeODzDUZgVhT2wWhM8gAh7nOM/pWqWZifS1uHYzn98aBIgQNuqjv3oqYJ5VPXpN
dslREX04063P12m0YvllPJPHX/0jcTeNLe4gNXaixik=
`pragma protect end_protected
