// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
J4yNlQu7AOZSy3BHt+DQNQGUPk7wDrOn2OAgGBzeZWtGsNDq4AHv9r76RdHX3OHw5xgAxKoJFNjA
ofn5I6TYEBvLedwc6dceeiNqZpIBGXY0Q8gMdbDwQs5hwp6q6+1AoovUOE2JH030ODLsE/Q6j/6R
2XUXsSRJte7ydhz6GP8kdjiGAVTeRM17R8/PqnrHKacpt4ts8P9GpHjQ08mN3Nf0QLAT5UASfEmA
qgv6DUNI3dhj8xlORNuMxeJfm8K0F2G3ItroANs2leyXrfcYAkp3q+h0kzrkp+S5uIbN3B0068FP
02XFHmTCC1GcLCSNi2h2qNEOJY7ygWx6YbTKzg==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
fkP0erk4ccHpMIc681/hqAheqIEkKB1KLiYQ1X9QPu3hhmObZ+0x2EEKDCCeUM7+WLP2o/i9zDuV
vgVYnDENUn/52VCGpkZZCoN5oGvi+VQON8cnHToLuppK1a+LjhmUPrdosC1o2diwTe1iqEnIVqpa
V1q0XoKp3qcorNV4vzQobJEW/RC7OSVsHP0WXhD3S8EUDFxjr2Bcoab/JxvHGebJvKHJQW3+3MUb
GTyb2OCDvLS7o8VY5jkxIJ6iywGzw4QuyMO5Za+GjbhDSf5CVTIu8Hkawym8eE6kBVp/5j6dRMwc
vBn2JplTAxsaNDgrzeuQPw0nCt48Ie7rdfnrWheQGn+OXZpGsCAjVJPy/U0Va2AgYwMir8SNB57v
yYbPT60QkB9U0z5IjghkLzi1VPdViIqlSpSYn7B3A5vkwLy5aoA+O81AAwRc64Wuvy7n8FyFFT9G
8mGhgibNeNuyoN3H8P1bPmKfKJDDjMcTkYLrR8JN0D5j9vvaaAet1W2Px8rDrQdm0qcPf+bywSem
jR/Bs4pbtqKneY/GrcwzBEPxr+EBEZvbaDZeJ2oPBlTNophLtb4vOVe32SQWcLugfx7hDUiyLXkl
PO+Xo2wgWSbKBG8Jo935xCYBT2o+JUaVZQIALcwDEXg2YhRx75pCzqRkHEI0vXFXYnWkRXqheduy
vAMoDp/wvnA5c2BTOf6I4UWvd+sN2fv96Gl8tK1fCY75ubyPywMeCxTSeF+BDX4wVnaVSlbnYdx7
Rlg2af5YieGi/Y0eHExIz3zCfK8vvEuIGOj48V4FJOspT4S6fFuglXTx/ikTzQzbA5JbSU3YFPLf
3YJLmh2NoUQhFuQkbAreYtkylG+fAC14ot67wENcwXxqH/d+53orqvRNuENeEbgEGmt3xjxyY82G
NO3mm3kAaHOM1FjYsm31H8OcY1/ZOLcr3708Dqg2wI/i6Y4MDN0m+k9jcZYh2iWfFw4Alr/UfOHQ
yTVmnCvd+4F4JfBR0UrSz2AJRidpnG6xO7ORUUd+Rxgh03a9aXiLhlA+ZcQmIMksgGCHgbjoiCcy
heaxuiZkIb/mz+YDXjqm12RHLk53pbR1miFS23D4xR7Ct5Ct0I5STrZpoCf4nnSCL+ZmczJMWER8
y8msiooIwOHzumx63ZjzR+J3we7bFhBR8/Y711mRrxJ/FYbnAqm5rLIjLVBNVyyk5geJK6MtMDZO
MWot1udzMlOSmIfy4K60V45o+7kvVFDgKhH1Re/fpMCqeRCzF0x2+pYZ+FOZPZJMR3UHq3iNsTwf
6QbjwEy+xOc5aWz44KmoYAmDTGw78oWC9RRDWjFYklQBZCWx51HqCiV9jeqQZNC8OJuwmoVCccpt
+W0yCrWILFBFnMz3tqfVh4DIlPJxdH5orqwZoFdMP1GqL+YKxWUyrhRGTNdQ31SCHOYP5pX/uKVf
jDISyFDzWrRuIWNooKv5r3FM2GcNd2XLAKI9E476/Pp3fsclvaSdH/g9k4UVWT4OgQyWOgKGADlq
z1pnzmAmzLlDSqBezKD8jCnS3ii67YyFlrBzc4YhFZ4wzfqVCWBwbkRkDyuH+2vDvNmJgnUD8E/4
Rl3kAqlNxdXMhETaetxwxbbPB/8VZfPEhGFbRjVi9u7IseNZgLoiXI56aU0K9W1jLEnmELBmgTYi
vs1q7ZkN02JYUpLCfRhgVezMapCiGzM3kz6hS51dumBTgmwdzsCErBBs5cF4ly9Qbb2DmPhFOG8Z
+8cbIq9doi48+GOZexqAtVaOzhgCKLr2gdDT91lUlv6Fz3jK23RI05QKV0LIs1d/aA/cTTWi9kgA
FmnZVwCSH4JIFoXx0tvWpk92nKv5G3ZppjG5r5RQ6/Ht7qTetzKcJjp8yJil78ljUlO/iR0cTT7k
GcRjP6wx/mK9tQ0n7ZyXTQfgX8Re7jLhXDEU5a4sjKBv+WUsBKNzDPDVaC/yhWdQ/+naqjLbizn5
qdS/hjUBXE78aoErvevlx6yOIcTd7fetfwwMK5lHB1OLq14nyy7Ucx+0jAgiCuMJdQY8W8pAtm3M
zOxfql3BU7GaencYGYzRFzRrxbEtvJQomdl/MvLFtrbQsg9xM9Da0PhPkKy4EEDT1yxaRqWQQoy8
lSTz1rfVovhuuYopnpMar+xsA/dvj2edxAts82TCJhTNGd2OBhC7aAqz0UUwAW2a+KcYisyBFzRe
ptrhTyBCPQb9prVGAaCg4zi0faF8zDLNcIiHSCdmtH86N155JnpTS4VjJzJbhVCPGD6UtW3m5aR6
axFgzsZE3UNFCbmoaRb77vG7bSEtoLGVxSczXjn0uK+Nel+q7yfNM2LUYRGQ8PeT8I3QJ3LlY9Kr
09STiPFDOm+spZL8BBJKrRs12gmNRAWbmyxiQdh3cYt+0SyjoWuYoCEJRSenou0VfXVLQx1volr9
UhNDuNT9vvy87i02FdE/DE5vkPeACzFo2J0z5RTooQ3WrCEodx7/0zibOmCIeVD1UkDR9L3rW0H8
DtIAAbqpGkjJrJb8mEkwM6HwdpA0Ol4j7gyRW9SiaxCN9SRc9ZeKlansHFv/u3yHeaWo/tETxOxj
idBEcgevfioXDvabcmcNiNvsgEzgFfrGQcE7RgSroo29xpOBifRm3UjKfExigjkHJptQUgYgUTQZ
pu+kNoN40owNZlL7WFuqgC+JdjZykqrDa59oAVd9eBT+vvKYJek6jP2DdxF0bALmbAXXyRZOPwl1
Nd15cKR8T4Kq2mtV/ge/F3EdHQVSb36/5RUvoCqN/s1PbKjevyDA8GT0aK1UVL+KrMQZQJiT04P3
cRtY52kRd8B4qZiTU0P0mVyZE4orRU09OjCGNOqx/tH/fr4a0vnI76uSRAZZGQRcYO6M0IoRX/mP
mfydN2Q39EPLarzFwN86Hoe6yKtFlvyjQ+5iWmf1cxoPBlc3q5i6ai9HfqmJN8oSHywU6tM51Oqv
cmzg21/Mv6dm0B2TPCBm1y2K0LjOyITKBynh7L9wuMGhZaRuVU0+n5MLmeLRUULXR8kKLCOgXY2l
vygGnfstNiVjVfRUyFNC2tpi8lir3DCa0wbuK+X+SJzG//u/GAPr7W7tj0DX8A2IDWJMzqegThwn
gNkotz9kGG2HsXD7dzjHpNYhm+pFqCq22T5k1mRElHshX3MmEyzxQoU+cCbG96Pzu6GjfY8y4sUx
Rc7DkZXGaiBD3+dxymRECI068lSK2qiLcf3hPvsahRr6LY1XEZnR1azCbQlPUf9iCY6mOjcLucf4
A/4+Vs48KpuX0Qv+YtwYaPqyom8pVhvvjUEUkFpL1T8MZ8ucU4rICePc7DQupKAaKVPSTsSt1lxU
PEqnCniJlMfRb51b4VQ+MEdMUhMbpMWp21KIqYO8miY5L9Z0PK86yn2s9p+74w8wmu9DvqLukdTt
7rcvZgTlv84S5k1+dfo78p0FE/lu3oD2AiDruu5JsNB0/s/sx6qlAFb5SkST1Xt61xymJer3KwvI
zb02alX9Zx8YVNX499Q2quAQihsKZxb7Ci7IeKg7viF2Eu+n/9/Nr1A9AkvpQayqDltlL2x7M4Go
EvGPo9lyb3w6dFohe/RpFKQTp1ZjLoGEOO/Hg4v4bOZZS5ftBeC01iA9K78xJTd1NKZqXVuHmUil
DEognNOZLmM6+L6Td8h554u1uQwu0qmwjWRNY/sdoSX6k7XP9rAuQgdNtUmAtltf+ENFfyHuCAXU
6KRHXJ5EC463kDMK36OYeX/BfE1tHAUs/2lkBBIbw2yIzxwWAtjJII3SMjm80N2ID1qHNuEb2MB6
sNZswEkNTo9qVK5Zsxh27YO+UJ4xDo4lD4u0J2veBqIHDYOD0NC8n+20q0lZLTR8eX8zKcL33TcT
7hex+cbxli4o1D+IVebm5IX0EXIDBPYEhcr9+PmGlATKFPb9fWOiXlF+1v+nhH4DVPup5Qbx3LcB
MII1L5KJacgrp6AYCv+whcY8Bm8P2R10U0iGbvKHMOhWgvUDlZiAUuQyVkzzgEi1Dul7OIlasYGs
zVT2AKE417pYDVhPbCjcsjSemuwMyi2tGakpnptmN1wyn8S/g3jBkEq46kZ1Ns1/wOrPl53K6Q6z
MUUAKjHRZ+fSOBNd8/R7YBS8tEZAeVMylBHyJ4ie82iFcP52ZgmsY/nwoo09GkEj2ag6nm1UrOFu
A0jBF+VSSMNmy2jm1j2t2pt7hSXNhXbymO7O5RY6mMfCsugi1jfC/yG862yE6K93bKoH7CQ7yj35
rxwVnYdxLsTTH2LL+hcr/F+li0wa6/6h2ws1QhEOZkx9a6n0k5YR6uR7GV9TfJRL5w6iEmC2VLKv
bcmcXyF3u3qyak0Gq45E/2UNCLNRo0Qs6e37f5OMNevmTGJU2SLRan4sJYbhTbltXtdTRQOiG2VE
A1tU4Zbgm5qhpKD4h0zBdNySbZ91a6ZysfV/HD8Dzjx01vZSOuoOd1kE0pguzScWIu9qe2XRN2n2
UEScS6iEvniunU6/5SX2BLp99b6YZ3fSPnYu0vZxJw9G4nIStrKh2LQ3oBiZVcsVpCbz5m79XlhG
2Y80DJTdRqiBdmyM21oF6PCZFkYeGKyuciwq0knXR+KS3H9Vh5YsdmZVx/xEBkNhit0oobu9ro2L
TWZh1Ag1Szr4aTUDqLPc1WcPXu9DFbAa9rTGjY+kjUOkMKHskrt7cbxJ5zUiUGhGgyOLpQ/ou+bX
LU7iU4AIXYrUkCgejkjGLpQENQ5xgogiimxm03txLJ8xDDk/jKXspXsJMHGHrk5RBA2LT/6RivbR
wguEZOaJ5RxXGc3UyrO/2Fv3xnJCjxM3M0YJ0Xusr9mS6w5iPAzyzXF72ydGsjysdduhgj3J9pv8
BnjiuoXmBYJd4jUZqZ5phRY9BHlzXJxCByNITuo7yi/fPIzUofy6LqKMkAqKPdlukNpzia4NKA3q
hsAREv4VBOcOZa0Ztyo0FW2sfoyAwo1Ch5oHmIskEkzfrqG46kRttzOJn2tpI+ImkAMwo5EHCurA
126F30M7FLNY5aDkkDi7W8/UAuKx5KKMrwDiAWQdg6edK1QVBLtEcvHMC8pubn52tLgnjDI2JrKK
R2VzIx8u/CB/3uvaaR/FFMK3hI44BjBKCWna04gm0G3IBG9W6LMZiU5CfQxDAnE+ML34XhoH6m/g
iQ8PiFWIvGA7qwwO/3hyghZ9u1IRT5MyjEhBJ/UxWLT1Zjy70PpIPajxw2F/GpTeBvuAZ8SVBJI4
QIO4EGOvZU5iDcqH6xnbcPw6HzfpSbVBl8RMEOE3sZH8TH3GQyC7sTTrHNkEDgrD103c3zn/ap/+
MCcLt7fPgIAh8fc97KcRJd0a6eyeQO8rLlgFiKXVMioTnoQazZvaoszAlQbHTFi/r26Z0eTDWkdm
L+1EvRVzwyKRWet1vL2I7VQx6EqdluT5y5hEBdxhRR8lbbEwSGEANaTMwC2fW/fCh62PRnssHQkT
RB8fw5uXKFThGf88ZKgkrWQ6mGAUxod+s4EuwamApxAYWlN1jz/eTl6Se3zmrN3XVYUfdne7yOIU
MtPx5OpplfEsMe0fIiKzBo0YA8cQYVMEQP7ZZC0p+mVcwhMdsnWmKl+taFIl13i2khDifTke8Sga
75tzR2cZNLqv21f1lQvzUw2Yu0WiMeg3UE607RFsBW4X2j9l0dLUjNDOnN49cAA6On4uBaqt9G70
y7H7B31aNZgg2G8JioQgitNNSsLgtx1S2W9GBLoHbnyiHlvZoqxhsYY2Pq0ukVLXN3k4s6xmQucG
3Gmitb7I7QWGwc0UGuX0yoMb0KSdZXDTJDgo/cGxNtpcNCMoH2zeF3Bat+VueK59zHPt/3vUw2wB
Xc5UNpM2W2CmvoFrLmTPrIA+k+7CbPmKAyV00ij4XUTKwHNB3jdtuXt+qFzgE6ksRPeuz74xPinQ
y+RA+WFyGlJGrBdOKCalG6nZSvDX3diqLSI4m9bqpBwfNDwBSF6YXn3oVZ3yfPwrvKi3TP3AmBGD
ZteeTHmKl87RhLpP21kaf1olhPt/i9h+qqpv+3YcXSZUk9LjwKdq1HidlXoY31JF98yVUAMq0UsE
u0bPIFxtB8Wx9V1ktNDEmbn3uqmTaC8b987RNQfkQXid1wvPI4hbK4g4T/TS0/3JHVamMl3TaKp1
6XcjdQgKnE3KJQsUktErDvti6eguEPoGcPiUgOt7qOoKSMBqGEC8IQHV7rogr8bC/s+WtuB8Bb77
TWOyuFkg/oixBNZHGv/Wl+bNQ3vRVUikw/mZRIT4F26VMzFXdMIn4/5duuh6AcxmiZ6DFE9T71uf
f+xFw+WjD3os3o02lofSb6pFMyBmYxjLWzlkJGLs38Ug+eV3EiOOricLj4S4a5/CZThk3JWCS8bY
L8f6noAMvDxFD/R/oSdeEjWFfsjZWtt4o/JmR7W3Sq8fXmnAcNruH8eVU+28hKiwLgl3p2rkYWHD
ALemO2Sh8ItUtcCXvOdm1RVFfXuh8GXWf6Vvmg1eEintGCXmmbcnk8VSp9eIZT5gNQDGE14C0fPI
ZxlUgw7rV/UiLl4BsyRYfSgx+APsDLV7oMB3fG/cd75X7b7KRnirbEjoAr0DsvymCyOq5TF5j/RF
sl7YgOOZDFVNA9H2ha9UWwc3C/KigYx2wILt2DDICYttedIIHB2Suq80d5Ss/q+jCGtvcFn8laYx
4PQIAGTFRZeenye2xbuGbwe+P31CtK6HqpxRFYeZauOW25AeG0s+T97/4IpFcMJVc27Sj6vBAoXg
4iNEkT4QJbdjNEiOI6F7vSGF66gn9O1oHC9vrhFsUHExa5YnB4/4hqyPVAhFluuJYVHyokPo5yig
Y5OICuPZGU3wE8vCCKc+ziZyQHPuK1BFt6z0oMWS7pR3Oqc/w6Gj9VvSi6ErvVnMzDAs0qH6WBlp
cL8w/+pViboTmr9KC8xRxrxvUikEmfxjESmhqzObII3RVz01aE7geafOn3F8uFgKOLlYf+ScYNPY
tpU+vNpdz3mwkh1Jq9kvnZKt/X2bXzfrJgvez05ffNCVDA/eIQVJTe45V3rH1nN1+jUP5r2CnaAZ
gHo7OL8uCcSQDWEc4kN+Cz5fu/3Cw7E9R25h0s+MvBpskWdGqeB0BWn/vi9QD1IVk/YCjGd1kB6+
gpm8quPm2iku7r2JblzkFAj8i2YamwnCK68XKlMMtL0pFSOm97oPlKAfTd859VJxxnlqVvBwEy4U
MZ1qAjLOJRwRrXUo/nkzCXJQv5sXV+o7nvFsbIEIrza9IKxxQ5NlG75Wv0qVFKep3ppZBX+LV2Jr
oiVjTVZh1Lsl3HtFLfkU+rGX725fEm3JCrD2aZIDV3d13JuVdGaG8eLPIWmCPLaFyrol2EBa8yux
nPMuJJtPr41GCqvVpb+C1hlYKzllQ9UlEvXY96Gk51yRpn5bvXFuqen/vOIlCXVdUBPw7W63zPJc
/WKzgVZwMg5+uo6OnnI/VkY49IXEA4Cibr1oAeStEBSkq1FXmZFV6Zgmn5XUvFizPiiUBrB6wJLo
KdeMlDWiru/vEPBSOYko0ltGOtYGzKt+6KMtaQUwU4VzMIvn7fdUURvgg4WdRIxiVSxTZ2SCSGX8
bFRTx26lEBu3GGDggDxM/WHw9iCCYd3sOx3PvQKE45D5c5Vl8NWvINmLvAJn4lLkxQ207ayMmS9s
+CXSWbm2bgr/2E8mTddkzBhB8C3iRZUJhUhys4/0CDG7EKI894IevOz7ErUdwQqZFgK0ljz5kHZA
eOh7a6qVRG/kJn8HO10kM9r8/cdwCUoUTqNhGja3vhGhZQnq36+FoAE9OCvw2KF+F15TRHv4lmMb
Rnz5dZ3olqoqXk/biaXKH4NvB+HrC21XhBamDpAueEMh50Zzm9bNoQkjP4QOggxGLGogB1BrGfhg
dIKU7jj3MRX2X0IH2b0RoVbNB11pRYQQeDn+6JnE/L55VGnoAzzmi7kDngS0RaJD/8n7EtbIsQWs
Hm8ux+/1/qnQqO7svRuJffcqRrsYr2xYKLzNCTVpgp2QSdDVmC2lPLje3o6AJdN8rF9sPEi/kgEg
HGbvxciUQ+c95kYx0sgrs/o3s4nq9XqDhyeVwRykGvXKcUjmS4E4YEeRuE4bNHqbF4zeI/L7kZ+U
TuFet/qfwSUOV1CuK/dKyXXB+Q1rDgJAENO0qOg3QUjCHAgK1nZiObLWkZe3E6ILTIi3GLR863OS
ABTu3zyHiW6IW/hiJXeqnt6Km36N5TWSutzuFRAYiiPoz16yp1PUnvExqsgZX/qJvj+ph64KWaGg
tNWZ0ByIiTRdp47adSdIePR8fy7DIODpAgbWF5otCafJujzyGi5cHdruOC/tSw2ePCpYU25yw7mC
fc6Mx/13modAQX7UFIQ0cBkGQAVZSZVIfWUFzF0+DGYHssxGZOZ/qQ6qNC7saUSHHW8Y+sWpYuRp
iR2muB99n66kjcdnzyE56V3xLR/8a5iXxpA33es6fffCdk9dhQ4V7scIjqrTXkPqLAAHsA68YC/d
0ayzan172ymsSyNAAiDWYXjGMCj44y3/miEvepNchvfPn7Mfbcp+HXFouVJk7vbEZh5eO6t+wDAu
2tzWOgvIiUQr84+MWS/vSfi1mczbiKxhiUXMJTkXLPV5GkHzuCbZD2payy1RhRmNQsM2lJT1E3g3
+N/KDCHmwXoE25PgH/Jrti/h/sKA7GGqInaJG/c/g6umubF0/Uvx7NNlKY0MNO18PXZ7YSF4ZzzT
RlctnfZlwalBNuaEeTJNknCCDCvSYGUNF8AtmJ+mjxx4R5X/iETLH2NcOu4733joCGhWi5C5AzkG
JSWRsgjlUG3Tu70OTv5M9cGJtz3uSAK+T3a4kiSMMVXPSdeB81kPm8qZ5CzOQ+UGNxCwS5fjQXpg
HvZ1YXIJLrBGYoFRoF/tELPnC4W7Z+sBDkcI/y9HFzPeXfsuOG07lB7oNh7sNxul7CB0VpapyIUM
+cLV++16u509WBcIII9d7gZBjsfbIubephQzBM9uo+0bCq+n9EzKN+pD7/I/TJPDkDSWs47FuKyv
yEj+1beQ4p7VJr/Wzlg1igrrFIVgZoVaDpf6zwTRcTl5dW9vKrqGwjjS/cjIHns9g5InBIZFeiTG
xcuOI3zGc80L4NgCzCrk7uIL76/F7E6HyXVbG96gAokchOxOqPZQM9E95wAcXudGlXeLo12Hz/qf
KId0+Ve9VLWrxiY+7qpnA56dAzhKS0D7ksW4IF3F2iXMjwdqRB9d/QoM3IXNvj24xYHEdmGp7gFt
PjzIswqg3IQT0hKB2LeD0i0wg2gF4jL97ZsE4bb6XRubESsPv2jWqXw9oW2d+jp9M+ocE1vB6BaO
l5qrqn+GZoDl5R9vWpnxN2dfOr8Ln7iXa4QX6IZzw8nvnuBjZwzhq0yWUThi3oIE5Ni1WSjAQdpx
LuzsNPfImMD7pIcUZZKz3A5NM68/FDLwkiz59GsonHW+qP7cD65Q8LPiNCpQDgNUJJ33E7Df97NR
ZabE3CsCDarjnbMwhsktHBdarofx5vSHT/PCO0+vCXBuZ6Rgo6XoQoE9yKZISw7Imt52DPSyXyxO
9iuqgODcGVuZWL6uHwfNByxy31ufwgHXm9CPl3TyhzqaBK3SvNRZF7amjg5YRuxgojN/ygUnHq6S
gOVHZaN1MKZQPyuConE7M5ouy1c0ePDjc08GWL5Wf4nA1NnmFvVkTmjmzuNziOt449acaHEV/7RU
3j+zKL62g8B3MFZ2AhbaFmtsRK95OTAs4WcT7qr8a+vBo+s+5qymb2ZDXEdxFjv57RY8wKMYwcim
jSfOS1QVQ5l0f1t5jJC7sQBgxqDoclk/flrflj31k62kbfBpCOX7BWbUduai2Nud+Je6udx/BnSZ
VlxTSxuS3bhHB/57ZENoFyqtY1wXWOZZ+4Sq+jHya6BX6TqZ3ejJJvOhjFOR+gXORErhyFbVTS1H
QNOdmZVx2leBhZpohU2Bw6hIIfNdLen2nIAdWvE8fnS/T/jEnQzMO8DzYWgbkrr/cZ5zSQyjDnlz
aTffzNIvcKrJiy+9y01Hlw2JpuLhY8YPVPfyOWuGfqoqnz32JXA9XPDLKOUQzQKvWarLTm5LJTXi
sOaUJk18ZzzW6p5T0JUFLfkkigZUkAVLEKSdU4fonpyLGnQeRzjBwgbM03rVJxSJn2Qs6N49XrC2
+5SSKPtXbI3dZxjPXp8j2aFMNAZH2RqoSzt5+I8yAEaf81NhwUEt3NEu4SQ8CcXa1SZSZYbLb9SW
fqBSHiqJW9hp99mSrkBQ4WCjsgSf+9HCaNAOd4n9GhBfqYzY3LRuVS7ogrBidiv+favdpN1g8CRK
JYRQEXsethLYoHQ1kbc1vzlfXWadgzpKdmFWk8UzGcgq/e3hLood4yzRpA/r/dMd7fyMml5KA/Dp
m400NjYdOD3eYPy46cNit3raQnDAeyvXHp6iDi0ke+YEtZ0kiW/GvzZ+yNuELQBR5piOgJCyJIOC
kqXMjXciIoiG4Bt1yKQge0pGiLUJNdjqj0aDWTsODfGfYGnE3LxyEUsExYVrN0n44z/RzjZtP6Ps
vU2AzDsfr3zaJM+Yx3pxyZR4P3yML2MmaJ1+mQ/q0j08ekf8xNcvuIMDqDB1MwxCXUjpc9nMEEnV
Lcd5K63sNNVeuxK9GP/joNeQNFEEGjlINS9V4xUkrDpp6wkd6rfl9bwbu3yG6LJZIc8KxWYxabwh
wPUr6F63PAZCB2jlsJRrrYPhe16goLffL6qrp6xgM8zye6iEXCFkq6aiwYp97GCATZY8TNSU4Sb9
Aao4zzkQZNHcH9K3G120lHWOtupR2UZdCHLbP783TgcSvN5YBfllL/PxdQU3G/Qkh7ys9HCyx+1e
e/60Y4bU0jgKE//g/X04PJijKtSkBer4SEugM8M3lkpwHjmHICVs2KrJ6lgyeT4hN7NzRCrfKn4i
JNArbIQdTmogZluBFzszroQlV2asmEQ7z8pzEhaQO5np94ODkBqw57lDlWoFmpQq7yFu5YSPqJiu
1EdxjDuLhXKD4SZisvqTxsIAIAqzf+Ze215f3DIpkbyTZ2xRpZttmtiJ0xjdnxPDwSaPsR7QKUUa
HD/orT2K2XbBkVyLd3//KdUCuVZrAV6SwLru9ccr7ekoiLitq5GjWxtwDzW8QdlL6O4WyxZnLowf
McsaL8BUPRWfBgN2IgBWR58qN/gEk5Mg3r2dDDKlZVu64+knDdG11EQjHQLT7rUvnGFnUbepqgXD
s4ImUkIKOTCPf5Dm/e9rnGpxqUYe1c0iFJSue1GrpWsSZ2D08ClqCTbG4XPdBZj6+fr4vdGbZyK+
rf6dFjhb8+WSqo7T3kN6K7jhuwHYPqzXVCZ4teQLy+LC2Wrcmjet+WeDy+ssNqMpvOocdk2eovcv
/hYybPO17QaCoTNsgfdA+aCB5pVAMBog/unFAWIreXrXfIIxPVP5LvqjceUH9iEU/ZJJ4tc3O2uF
zSO8yvgk4ltr5piG//K6f3S17awUyYaGf66eeQ/2Zx4XGnrFr8zqGs3mmJCQ4fYZnoYgM9b0IRuY
hLKJ8f62TeExMo0Fev+zE37DSzA5P5LoivCZLrw7EuNOS5hCZG79l0wBi7venZuREqx57W/iFVrA
qIfxHGQ5GvwhT7Ar3QNAY1ufXIUsytF/1YA8GdLSY5rdVh27WUALUK+NP+OoXMBSbdKr4ZBGpVnN
vhkpxAA4CmgVInqVmik7mxtcgjls4VsjeIaBPR91ErbtFHPwJW3+DiEkyOmVQHuMdfo47sKUf36E
yZSQRoae9BGUdwd2QEFDdSH539wNLZSNH33r1FfihyfTH5tuE9VTNSdayAVgkCaEE8jN7gIsvZlS
4Xz67BIVZMdtaYuU87wNq5IL4icZ5nKdOqqsPbbs+5BLgLsIeMwhd4ejqXt0NYnSZ5JHv3F83Zkk
HrElgVDDgy1RwyN5dxFzrSJIeVF8QuX0as1MH41dCcMjB19L65/noamz/Ac/5lOGfwmc8gTkzb/8
dyn8IJq/SS1d1BEHpvAsiPSGd+A9VT+XCNvrAMiFdPyC0p2z9WdSUMuaFK8nGONMhGVm2ZybZ41e
aAw/virIeVB3DccQfuL6YOvOxWnKEniAuK7ehKFy/EEiaK4DUhDSVekbdW8bsZrjo8OIb9jPeLQ0
HhP26xVLmZMK8f7Ry5+QWriOIt8nDEpDzlqtSDsXEzQrf+VaoPhXIbeKtSFXZdR6JTv7Ad/Mqh9b
l//eNeG52jIWTBkz6ixulorRSsN9uZSzT1p883qlz2NjEESssHLL4Th7TN24OMVuZQfZEPWMOdNd
klQ5keyDY3vU2MWOc8AKBBF3fUNtSXqoQO2eDqqUJ+0uZJYQPSmDfSkfMQPddIqpKJ5X1rGtdsd4
ti6LsP7B5kl1yE5dBj1b/7n2udoQU2S4j1naN7SEphfPCcm1aUB+a7Sd1jwBMLZdm2Zdos0unjD1
k6tTHbghlfrJ2KRvGsceDQDryuT9NQEYL6XHxWHjX/cS1A2DHLiW17Wp90dUeij5hmkzcGh9BZgA
NOuTQvw4rZ/VYymgJwcItYbdLNdsFDG2D8sYXu2/vE4eSFpeCCo3eUt/IMjbK8wPlqzIqB2fYiG7
YdkbXIHOLrpP60Ta/tAzvn4IU1IYTE5U0mbco58hAzjp+dZe0zubt91HMTFGO4HMKgstZmlhSZ1F
EeS5V4CuICV38h3AcKpoX9NFwZI12Xiogbyfe8fiW4NqfWmcFJTJQJAXm/w2sJuZ9LA8kIbfD2j9
BqsBYUwuGf9DQB9bHo5zNaGEAyV1oEQuLucZi6/Ggv4emN/9o7X12Z5+lEPaRPo0R3oy7jMm82nP
/QwA4LvxRK3G4OWyssxka/jndM1VOPIYXM8qcdO2yNI40nSY4XBuSUlOPZxsfbsNJMxUz9uzOrZx
REvgohp60omO72jvILE33yUcGFOBdDtfsno3g+nPvW5UjC9VZa9TN6Gbx/z0Sy73iIJN+uLbK40B
EGR9RLA5lfm9s4ezYe31WPRcklGZB6ymKSUJITBFOjmek/k7rtgmAoi6D5Td+Ct7D9xNhHyV2z4z
gaogWvEQnFIUrzxXQsIMudv75vKV++5Y+j5I1Prp7bJfnc/SEegLj+G1NZOOb4pLx+jpBLRvoTQy
zIqWX4hps1uriYppbz/TAaOon/gTOpHmndhDXlv1N0atliAyAivlLxSnKDhIYnnNL9A/9v8W6g8O
GLfLnNSV6U4TNcrLyx47c5QBTXjyuLl/4DnYs1UxOUUVw+F11PMdmKusCuMlROYu/iz8guKqVKKK
XBI5bZ4leOtdEjlFKTTsFOZk5r7Rov6lxdJBLcyfFkPAxjlB3hqMiOolxbtL6HvXcBxciXqxZbPR
OIRDc1VKx0Ue4KIRvPKYpzoHMqo8hWIITMw1SRq2DE9ybgI1zscRiEhuKERwc0VVZMgpVmA8OtDG
N2uN0MCtn+PDOeckvREcW/2SQrpC6sIAaBmKEc4WsxWboO8fqi3pTNxsB6VsGqO1wcUGpe0U1lxn
DwCfHXQdC85j1IBCD5aSCv8K0+3lEAYAnYnTDUPseFbXpiaARUWYE3eDAQd6q2ngthsVYvDFvjKq
7uop74NTlLCbbBr8YJwzN31UzXa8kNod/KWeLnDHBl6VP9tW439t+F1cqhFiNUTzZShgyBt2YNGs
C+g+mzV7j752jopcwdCuAnH47FWR4JWYoVXvBSHTV25oyhJ4E9kkTIlF6vi23HUdTQ8MTPSkksU+
MAT9f1IAMQr7bWAcPnqAC5QngGvqM/5hlKQ5f4NTgbea/F81ICOzledRt3FVSJLHh+G7Jo0mw9es
0OsfAgc1aVweWgXbc3t1qKHcTL2XiEc+kuXZGKSwxrLFGgmuTFFv1R3VEQv6/OAzdcpoE9iC3WfX
rdspE2nXAG7qe3wltyb0K7ld/QKMwiTKZmDTxXJAVyGiyS+w8Em+Tw8E1wZ4SCYjsYgAXo5jAbGG
A743Dr9G00dU8U9kKFWsZT6XfpfZAndqCybC39gDTOdItmHJXR3a8wdW3a0XbzOx35CH+/Ot/a78
Zv3nnD0QinzML7mmV2xki20EYXkmytIT2J2lHhUk8U33WE0ZxUF3Xd1o8qGxyoLGNEPwzbyLlvO/
Cbdj+hioa3wQyVo6EwKLTnbIj+14aowfFuVupq1/ybcO3JMXynh1RlvvQt7IL6XnsfIB4Yeqzw99
LXT3VINtV/cVwDL/X/hFuGjoGf7W/FmiQeHPnMap0h0pzCbF00QYtlrjFlpLdHxA/Mvj7KxIimqR
6hvHcfETPJ6RObyEB+80WOlywmBf/CA+2dyX2gOFGS38ulSYDqBeWsvgwogZvhaAENgZu/4L07Ww
2gUBRPTNHG61huC+fL0b2L+x5/kfVnPr3ktfXneNag3smm8Dh8NZzMbBRfMaWFDspGXHsel1smb8
saIAh1EPWXZkHdAoENyXtmqTJhUg6rJxYN/UjNg9d/rXksNKFC+rUNpJqV3JQ9mvcjaCVet4EVTG
QqGooo7iG60rB29hgRbzw0pCJFExFZNcL83WqKQbQyhT1ej2gwUO7cjmLJB1eqj8dsxWBMNCUMlX
PzzjXkrOHev6iZfzQxCtXv5eFJfVk4vvHf2A0pJJEfnd30uf1UCiqiS2WmQWmy6lWGJN+3TdD9Kw
ep9FHeGG3nQqWXZQ/s02w6RLwB/HE1BqOg8dmvH8f2pVR1T1yc4UpWrZEHi5sMgAaG/xwJBt/z9a
ND6sCd5ciFQK5WKcOeVQsYlgY9Bt1Pe7hnl9ox0ka3dGTj0CplfR1z9GNzlQUV3aUIIHVgAOJPw1
MvC6gBg4J/vCx/+53TNiLNxXJao4SSm69IXQIVdxweW6Zf6h0WLKzw1VTKMiKjTmd9q8Ihoy1kNx
erhnc5oYEdq/voZ/m6kDt3HgwjmZShs3T8nx85hBZyO55tRG709ymmE4vDakFzymwn5PTn7qcw3j
5jwRQD54ATVFZbXvaa2OXu9RRx2T6jcqN30+8tKXvSuZfneHk+pUj09oTnGdV0c/qGwePVUMTh/Z
thqayc58uWnjaCdoUAxiv3VzUOzcTohnR5zNLkveYU0jyj3U/IxOtHQpg6BegAAXmMxvaPC36SSx
5Kf8Xg8GXmZnqdd7a+h+e4F531xehZ/nvqSMFle0jKEVHrq8hY0Jg7gFG1Ziz+8OK0B4NmMJZjH+
GHns5R0gP80eAOI2ZwiKSeodpSX+F2SV5qhYOYZHXr2hmB5O99TyGPgmB5HbWeGsmxTNprP9aGDa
8RSWrwZPTFSfwJjmowdgc/0jMYB4etZ19OFL5DhjrFot3ofCPg2tSD50ZHThrp/vZnB15fevsxM9
VxZxPK1OYlt5GJn6wsUCzngpCsmImHrxyn8sKqkpje36VDBEwR+o3H+e7BHtylpVgwO/pMd/oFUC
e7KVPdkfvFPXiOpfsvF49PwykR5EgEtgMOtn+3IhSfigy0XJ43CaRiLh9ylbcKT+xxJ4byr/vewP
b6ihgH4oN/dw3o//WyhHxnYFMWNlp/nnsoLItFx5X7xKP0S7VQ0Id7QD+gYyGpWRt6z395fExlxo
dpT4c2sx2DErz5YdMD5kENE3TR9TDZcOb5e0lxIZXWMc+QNEegeNGKctGyw3Sx//WCbZEdspWZly
R6wfALOWyFqKno0GE6fsD3nO9SeqMVeUCjApEhHSmarLBkOk9J+yjuI/PESjaxMq6vIJOJfTwF21
Eb+gDW6EF3l7cWxaetRhDVD6h1DR2hnlKqlr1EStbwjoY9cbkP0o7GgTtFHRZsMGYlitB6yD4Pl0
ReFwhKpix5gQvv56o10iWuXjnsPOIxvBCeThEZk69eO4SkkBWHn60pmZGaVxIVWhWnML6wp0tDz0
AfCZ4lAxidJDNt4myZuV22/7ukAVyKyyH7PAg/TYXF9CsOzpU4eyOFi2Ie14Q76jPEqwkcBEMr56
phFYyTJ2mInX3dltyX8HDprHEelyl/1B2oSCyWlwsKviH0QfQkhXL5VadCHuHnmtGizCe1LORZS1
vTINZWnCtaL4qJViAl4TAenPqbYgxh0HXiVzaagbj/qeABVua97RbeK+EPsRvVZO7vEQp5zGNiQ4
ZXuhuRgKDgFh3+8nKnbxAupwqzofmQWA5owVF7YSAd5c97eKezXgC7Oh8Itwkv4op5fUEZv9hYsh
0Dptf+Gvnw3dtiH9tZ2ItoSkV24HFoGtjjrwjc32k4O70jMusJu9DgZaGPEXCj/ysMWFj8RlG9dX
RNDCVUnbqNtzMT4SmSfpKL5O+LrU26dyB5cEPylzuVcmTXu2GKr3A/SQ9KXRnEQr2nSfFrKhkuac
d6jKKIUgQlPcqvVuCoJscpzsIqSWPJBAvb3dFG0TXn5AEM2E4ay6XrmaPWD/n0ktH7aORyW5GnGK
OYVDAsnsofVXFW9NaBP0KXcMHMS9XdcLPfLTJgNRDaIz/2AkF/Sdv9lKIcu+MVfzwTT8J0Fu8TAZ
FgTPFWqwm9jlsTSZdC9Zg5q4N6JORKHO1ud4iPXZ5XoMLHiybq00Z6XwiYYJIcf5GMCCU8BPqtTP
suKIjHkciB3zOuCOykNo5QKC9JHIbA/D232l1gsf5YRKXm4NZgtE6j3pF4b4v0AJzqSM9gJX2NVI
F5p+rxvI58rLCkxODifYXCdCKMXAzgb6W+1i7D9HDaaYcBqlUkELeg71D6cO5fYRC5gvPsUQOHBw
ljGH2C4SaS1g+2m8k6clvd44vcI+ThUm1COmY8fCv+O8s/iDga3iK5w4WBPcAbPVAF/V3eRU3dYo
IhGZw849AKJ/ljmr3ZkyUU+4hhzuGV/1Gl3wEylnEmOTRv0+op80/jmM602p/wQ5lJ3B48b54dcX
Bxx4Qf0apLT4FKyRzKFkixGfWLqldKngMrcC+wBZwE1I7sibHkKA6U53JqO6W562d1xutHoVMp3w
6uOHVT1D9F1jaPju8IO7RbpRBYwhq5c+f0uSn4Z4wnq8hSw2T86Fe9hNQLfFrQ4RC/79OJ19KxkX
rU+QNrDR2eMQHgkpj6pV34DmrIVPuiH0NId39tnK0zN2o0M0ApLH6df2FTA34v4MbDdJrfmAXEIu
KNKV67U21BzMwCMgt2Ddt6zyXV8+y/908mEjMbzwQVq804dEEJRXBGZnegcUNdPhizwQ6tXC/du0
QlH3R/5/vGgxVnlIKyBorc71KkP+KJl7aSEqq3Eb54JwdILUFpyTyKyfdeWTx6UTyaGXOC9FvBcR
Sl43hk+1IggOsQxT5aBQ8laSkgHI2hdFGUQOav7fkrXRXfJIRjCUQHm3OJe7WoeTIrgAbhFwc9f+
KZVb2Ew6TF0eZddZOPpq4eOIKhwvSVwD5bcVlV1b9BzkneEpwATcfloM0tNjXRU/dJlQaP+eVCiq
kKedMjhyXWYeHGmFqqJlLrhkxGKOWR8AnPf++NuSnImteshf9FGOfs5hZVIr2KDfgwx+t6Q6KICp
YJhbMIOrZnxvXV45+bP2a/ORU5CG4zA+oj55oNGPxjBksmg4UndxtJ0MVN9qSuoLpE5z1+R2V1FA
M0igOXnGDy9lP+HG0g1IqQSNXWivOyk+J5Uah9kBRmoKd6vVCMTbEn1f7fWHF9IKCwCAcvRLvSQ5
tobrnv3SdsQvSxfv6cZppD1cYIlXvYgT4+3B1iXIzECWee9XwXiUKIudWC1PH25lGE6ev6Or+TbN
Ci7ES+jchY1kDtQ7OhhN46tfCLH6BHUwdx7IjCxpDPEGQ78YphaHvgESw0TLAxMx2O6uuyMTZSrk
ae+L6+4DYkfNQh2jE+4MVVwyG+nrtcvYfRLRbRI6VpQpjLGoUg6nEpcg86xsVivcdzu5cUpKWs+J
NQh+AgyQbnsKqJIRL04FckCmWA3tOQ7ZoOGzyd0kBVO+l5oCJidotPoXJj0CZA5NPblXB6xWWj1U
B4//ionC6GaCdjWK3B3krUxx3uwfmdaQIZQJr5ut9+KEBPyuuioQYJY3n2WKaEx5g23p6wRS9bbq
cQySDGNxzSeiCwYcSq/n5hAAm038MssNuLgPqlvT0uMVoWk38/LIzrTKA5iPpa63tkFqn5+GE7p+
oClXnSx+2aJemn93oCIcykRRW0aTJchJwgtBwTGinBQ7hPzwtPjmi0tERndk16K+Qzkod609Vh3D
bj6vmO1zh5dlqUSxmjVruEafot368VGgpdY1wt1jtTFtJVdpbhISnl+A2WPrxRkFgoFKbijTCxae
mnrsBcSUvIRVWrpaVlAYXqwJKgIlBly/E65uaQMLswMhE7GctFSSdephvAUWv/wvcgvlSS22NaUP
m48NNd49UfHWzQUuVJVtMXYKsb5TFQcodWEoid7mQCYlNxlDi+66JpvFUcwZXAP12oFRwRtemdLQ
JTuM/tRRUFWcssP/SbIRjs7aAsxGw2gjRGNvEcype5u1FAa3UCEbtZayqDjPveHX1P6Cb7r0aSrS
0T+/fjaI/Bt0fXyZvOHlJQSnbhQj9mEteN7wtKH5yql1PS/uaICfa75xQzGoknV76WurEJFLNOUG
Y7bucdFmyq+DInzDtXC5U9YuEjEDRKBxz3qDIBJtFAS9p5VVcr0YVj4hTXiq6jLzBvZ/57Z1r0ym
FFyqQhJwDTQIq13l6lflUWRg9J2r/2FNMaxTXN9QYS9afX4mRMXYVr+J6z0QxIivAbP670CKSKzM
RmPm9X+Be/ArZWLtGN7fz5iAEdLaiETXkn1ENWFYcL2b+F6aR5w4r/4lFdj4H2xFFmpQAS4FLl5G
A9j762J4jbm53Y+/h3XAvQK3fB9FVDclzoej+jc23Wgmiv3OHtH44I09rSPr6T/FguEgwjtunn0s
iQK5H2ec7ezZhQLJLSn3Jr3Owk01gNBkZhEim8LcKPhL9Q1er/mXl9VHtLhMqxoyoz1gbsSoVhaA
hzK5L/3lgL+QmhNdyE2YnBDg5Jj8DnbGQ5Y+firxeauGe5TMOfJ0wO5eBSdtjsPMDs04yYEmL2Jk
YsVTdg3Okz26FVhXPNnN9TgEZtOk2rsafnifO/rmHj40G0t8xM8GaPtwEs8JW+xOp1WgKR2bCABp
E6ICfM0d/K6QktYeulRqj9GsTV6p7oroUfC35Ze/vDWPVbo2DxQkBzapML8zmzKlMYCoArOhfWOS
gW5txpHHxIQxVqH07nrQcV/jZShNiShT7E/G+SrytQgZWaqd31ReQbYdZooyMiLeaeZec7457vK3
ljVp8DjTrxNWmrlJowrxvoaRJ+GWEQvRx/PwsFOlZ1Y8UYuE8bML6mwIU1/yINcBzdmv1xgeuqzn
FuRSkkWNprbV/NIhhF63WUuqw1Vf4Tl4fA8WwejBcmYL7yO9IfhVrjq5VAI0eHyE3ZjW02k30qmp
vr0BzgQWzHeKLcuSH4bDXoMe0U01sooWnKc90S2QDqRxtn9jgwh/cbRl4o7S7c7D+sKifYoe2n7P
fUfqU7OvEBjV2D7zGBBEWIeCLyKUMGkx2ikr9tNi0Azv39fYgCl1Chd8K7YYM8Zm7R45dJphf1tj
TTsaxbnogk0sCKDK4rFnP73hmp4p/6xNt2xm/yj3pyCYOl96hh49flHoneWrYDAHlLLVBqpBEiM0
95LoITnz+ID+SFYsqcHU3AgI94N0ZUBI8Ke08palfIFmLXwmCAuedCSWx/5lDPZaCHfbu69Z9UGt
tywy1zzfY/CprDv4xn2FfIzxpXHtZkA2XZliXF/mV7NS75ZVcgRlTreK2nOs3iANnaEYXY6l89Fh
jaDdGExRznSqt4RDfSRGrf3bb0Tws77x4nHsWLtjzgSpHKau+VdxwxTqV7GlI6cEXaF0DubUKbqu
3cO2BMN5MwcRBCph4N4fxZGCDXn6xc7IPnorbEG5gI0yPX2hJzjL+qGIHCuuJMqFW3N9jisMvJZC
Tsri5ZSOr2mJFuwh0GbrliqtpayfNLentsuxCZrdcVTHsIi/okZczHwduAfvssqAxa2NcVY5wYyy
EZo+dERulaEcVKJkES4FbFMJRRYtqP4BRJHDtlFLJnb/uvNWZ+lvDp4nG5wiCcG9ObsaV4GSjafl
zF/sAeE4U7IK6nNfae4SquSWjoXRs1z5AndsS9wlYv+RHaoMP5Yn3jW1zSaLkfwfERbIfoSkDwku
d3VIbUFXEqsXPnE21ZixO8iMoazmqLpm6e2L7QSAGR0RsDi0eqhIGH3VgnzjiUhVl52B2010NQ1X
uY9ZN4p0IIUjAai0+8hl2tDTuHrvUcBghJnrMcGs9sKpQMTIe7ikTLWbjo1UQRWLPgdXQL4McEB3
RjRgNb9XA8IotkGOsCShFPEzRoqHFPas6sOJ514qoPG8QmdECcw5YfmzL7BPOfxt31CiVy0XHsg6
0rm+tVWnY747ZQlEovAgaamR24zUGyFYanZo0W2MXrWagIm+Cg2deNDQ0PYdXfO7tyGLSYwKU8dL
LIvnx/1qxtzjKV+xN9b+Sjbyps7ntcCidFx7+OzUrhduQcmefRcFyISfNitnvY5CAv6thsqLwlhP
KknDjtirJesOKuTOshJqjdSD/1GwN+rBYGM9ZuSRUtrQqBC0OmuIRHIHhFawA8OWHNqSF1zxXpJm
dH8Gn77YnpFJnq4JcO8hjDrltzHQSMqGw4NoCR5uLXbfkWqzE5flSbn2U4wzyxOPPLKhikE83SM5
JU5xqtEjMPNlswN7QnoxRVUKNJDBRrjVX0lbcuBrTz0gDSbIbQC4wnP9gY2s/XYha3VH8ryCbspA
Zh6x8krZ5txgedSr6y7q4deGMX+XZuKseVeb2Lyn9CH70nqcsDwSF6f1udUL1lBps9nXYXkhoSG1
2ZTY/3/Z5/eY42qtbJQz6TH7emi/449Wo8dODfYY5+OLFmCAUA2TQFKJLSQN/NxSNZ6uunkTMN/r
LCQT3QGOIN9LuwsqO61IATk+EgfGcjb2XNn/MNZZHj37CdJv/h3dctOYbAJlJj+gbKvs2BPzBU1+
AQq7yk0IdcMIE2L8dfZLub6A7T8BqrClzayGkmAUYWE0DtszfpVrprFUg/jKmvgtytBeDlTQER2p
DeLZwIAhnyX6jyMXWQAxPD16Q3tqJ/DNaVN9rnfHhWjeiYlLsHBvB5nCsiVKpFUk2BMfSxRwjV/Q
FkmG03EMjQDe1HB8Y/DiQ+Jd4C78ah7dDTHtn3p8bTLnNoe+IqAOIGQaLo2toq4T4SiZJCrJLMS4
vy6ZRASvRiefQr0e9gBCo14a2spCdjEY6yzP3Q5rcMfxQLx3xWt2sUo2RRERUOqgtzHM0LAPhRVl
FXQivqbMF46hWCak8DFHzQYbDZKRYm7c+rzvX64LVCQyA4b8NlRrHsx6eGlvuXdYlnHOvvcYZ3UU
PkWymDNB2vtJX6hBIX6xrpb+oQgafBlMzfEonCoQlsE1rOFU+T2bho/ZMuVwWWSPAyRhHP7fPPYL
O1WUe7mfM5fxvbOpO6N6OSc/vcgEqnUQAij81A1eC68NmE9JXAqS4qJTsJCSAq7m2dsVUxqJakGh
GfUjpQtDcH1pOQtPy0vhpbgfJUpH2ERRIZwCk8zHDS63+k5ayiPvvM8/EiswETqB9HpaAsaBbgt8
uhqABhJ3Dm6xhABgfk9w0NpIJPTBBc4Tjmw1qHQ5zUtYhP6BNiag/Xv0yRlE8L/XlWJBag1KL8G+
vBgVK6m+RtaXx4g9sQEjDv3cV0iAWyl8V7HPTZrFfDRNP8zVdyptABeWkEfjACyCBL2C6NXbCy6m
xyYxud+VmH6K8xCVjf7TqaQb9qOjxctSfGhlaIu/zmjrL4FCcK/fZaZNEDRt3Mb5AspIyUF0dRyY
Hk/wWJMPvfJEKpmT24BYjMuFHpSsB3OXopq6/lrUS9K/JGMBl2ups3WO2YzWh4DPJ2quWgGMyvGG
jleOOsgd9u3RIR3TFW8vtvUREQRkDLl9AVkePTtsBOElam4nl5+dNEAOO5JpzI4m+kaT7l+8y8dm
s9KEJP/6csQJJY92+zQWJkqO6L2w64sstCO4+EFWLbDsTsf2rCegaQQS631vzVYwWN4IsKApxicT
DBZCmU5dsBroLO1+23kTJhHVXJ1Jqafe27jMo4A0ZGF72+C17J9zILsmJLrmky+bwta8gJnc8Ru2
n4w6J2xz5J1/kqA5MdWSEKI4dNjVTvtwms5XvuqsNETR1D2tHoJMxNDG35jTrHi4YA1r2K4ibhZ9
cfbDQj2QtAcwe4VvKvv9BqJcmLi0ViM+7wa/QiHpdzMbsNw4SLfkwcnEfISXz7VxpfeIGh6CUhV9
QTNzamo1e03RxfFVM2yr7Bjjd0mK6ZEC6lTgRYXx3d/+0gvSpAI1f50lPRgmREo5x82p4j+AWcYM
O2qZLsROKIFHBmS/NC5oD4bAASAD+qZoNSzDTJNyaLlOs5nEsl54hKADt39018yT8w4NMvOOBqPa
fPWEjmVqWgctZMqiWrV1NIVknJdhRRVqehWijVW+hWKbrWhGB3rm+xbQ6MMVvHqVnsOuNOGiLzFK
UAClzcX3RoYl62sDFzF3t4d/JGlClbr+54Iovo5kfEAh40g5GPpEXF2Ev8G7qW/N/qE0JLVz10xs
SEHrlCAmVj9S3aMkDdZF0DPSsOH8wde03BnA0szqsc8g7vsA9oUXa5Bd1exbtpLOYt6VWkZGgIqG
qaUeVAtELSwQAJLJ6da+9ta8Z1w1vvGO535A8jeuNhMMLukEwMgUydAgR16hmMWpDuzge97745FD
jB7Q5t1OVYh75u1wfBEKJGfst+QmshqQd6e89VFH6AWYy2WnwO3a6GITSQr9Omt54BcbpWsWQnmL
F+3axSLalSv7rW0RL442LrfJHNnM1VX/InLOUgwtbRJob00GWwoD6NRU487at4hI8C9480fqOi2N
UMa2PkhrN8Il4fjkOcb0Z2g6cM8wXTHczQsEQkPVaR2rLJl9AOPGkjEfdQfqXQbs+K04djcpsfiy
rLsLUiWdvPOeO4Ac3VqrX52KhLMt8Cnoj15b4peM5YodEcITcckMb6iElekmJnud1VTbun2eQw/h
zjlGxsDWr1S8lUkhWlirYpC6JMFUGHZAwZZIXOp/Ti+ARAjv40JikV8XOa3qz4hwSAVAisglPUPZ
9ShJU/W7NJ9/BY9nHrD36vxvu0UmQgDxNgmHRSuH0fPDgR9YwRcf0xyu8g8mnkvfNRmjtu7kKrIt
SS13/20iHUYl9QvqOeeAQ/RWoeAKRy8JCMG2suyAvWvFVZNVvJPVobujCjgRVCj29U6oSqnYkHOP
Xrjn8547uaU6vW4jQJFoooH/lZIbbXC6xHrRpT0jjN92nBvFg11S6rPPyOqJBjXhhxAdRBLjLyl4
gBR4S3FOiCXDNlaXWdNzWPlSLoWMUvXH4iC0rYrPMc4Lf21YUp1Jx+gY1uDsVO+a0il4GDQQRaOD
KYMA2d74fdyabKTFACjddAB+7P0nUvMguJ4zP9gDml4yxstv/bCcJF+FeDCi4KYneIzMDe1B9ywV
Z2flUxhefFj12MKf7UOTKYgfnapRALCWdzfFiIaoLCbTDjiqc98kys2x6Tut4deb4/MhO1A8RbpM
oXEcFXlo3UURk8q1TKvkW5ksesUwEBinB/kdgmweTPJrRqUBQI9+9LBul5Csmkd/v2jVeI3qL3DQ
qfVZS9GUzbA2ioCDp90D4Et+NPoHUpTh952tNz6GJHQUKS9aUQQTpTplQVYZSVJbaedNoxeSAYaT
maBINsp5FwGuU5ZA42P22QeUUwnzyucQnqVndJ47soOR0RAfTpvTIlw7cw9caK4ND3nBoiXOSHK3
saqfLMYbDAUjhwDVGBBSZqozZ/d1BgJ1q1UtnU9f94x0O50H8ImfA1U77XxHBt4vTlS6N+96riJg
/8eDUonIi0k0+R+ffrE8D3wM6y3oiHK5Z2YGDN6Ytu1qllq4iFGL4kH+Gkogw3mJNjFTzhZQIRjM
ZEyH0yobsvi3Bgc5VgbFv/BnXDAzA8Dr3guM8vF0JJ6TvHw+6v/m9MO39KHojbubbWig8U/GTRYj
dfAjJzD7o+6sXbfgWsyGs+Pl05NvUmEH6+G6zD2a9KJnJqHkWtO/TSc7W/Y/t+h23uWpe+uT/2c+
L3T8p6Vg+lJLqMit7jdOBq/Gs8r79QZztaIHSMkjDNv1+UZodJ2shXFg6y0rmKMrWYyqmyfLoJbh
8CRnN3BCu5buNfGi1bU+dcE6CUiumP4e3SA/mfBYPKg0ROOmBs34EVCpSROj2uYcW4z9/KVv+TE9
mEygyy1L3qveTWd+Ax5J/HymWdd53SfT+fg5A+/biqFBgsWSMKd1PvC3YoQGuF4zuelh7X41XpkE
TAgH+m5GavmQg1mZbLgIuuTygkcU2MZSYlMJQ6JtL+x2wljKyBtt9ScIGCew3AHIJ2IyvsZ9pRPW
POL1VpdqqPqwQ0pwj8PlCYoz8cXWn1j/IP20lab/PD5yt9yLrjbCSkPP5/O748xOsncjN4N9W47U
6ws1RNdVNaEtcCh/knWFSYutmA0hIUXA4givbhuFHsJPeQpLeBmbeyslQ2TNhcbaialAlZyH8UzG
c+KJmM5Eynd5dztsvqr8k1n69dtkFHXHsW2nG0HrvdfKU2RgfqkJ51MIVw6SjISRRsJKS6Ak+Vcw
qMpmmN2C05v4XJTc/Creo6JFZbC5UusHqC5x8prtHi77Dt9Rz5rovj7e/hoRuvGnxdLzN9AF30v/
HnrgwnP2CKXnoTa/ZTJDi7dyjy4qG5AOIyFDkzZX+Poi2wFXJjs0aQinpKN/v9ULTOF6p6ey998j
h8CdLghfaBykoBjhfgTSEEKPQeSPc1uhApmPaSW/39deN6cH9QOVhYLRMOEpptpwmznA4NqmXEoA
AwLtLtqSOhZQJ5a6UemU1S9tyfI3xTaAdEdb1hZhq+Pk5eG0DKUJtCcZweVVdrP1sLF9N9D/0Mw9
vXgwm6Nw/w9Z8fFrxECu+THZYDStAPImE/ltQEZZWIKKdECn9iaLeSDenGorc+6TLDcWEkflzRU6
Zv1oR7ahhNmuVbWGxf2ieUdGQDFY/xa9mfUDfFRu7CLConwLm6t6iLfokTtmfUAr+ZnQINPLjjM9
reNhJhvsjQWUs54+WJGTN2KaA32Y6GRq1cWdSxTJzsh+sE9txCVpdha/w9EdWrGxfN7d3KuuGW8e
LZsBfKDeCuQ3whOkbzzDP4+yTKtPPO+rd6zQStjM2kEyjWR3NrTSET1JT5ohb7hAV4gNRJzxA51g
tuR/75U+DFAd+Ib0Wl+WCsEladJ2XXp5PRVZ39QAufgJHPO5SGZ5/w1hx5ioSJmTy7SnNYo7h7Tn
J0i29gBmlQmuK8PaP+GptvDeE6NUt/sYQPqwx1rn5L6tyae2uDtoPNGwt5J0TxeJKzoX8hQ/Mksl
zyVPZytlr2QbrSJ208lrMOgbQ3qf1YIkpfdGUsuPzEaixxFAcRNiUiX9P1oPk0g8CjUqa3yVJEFQ
aEj3x6j0k+4gYxFEeob2PatduZpv5+UDQHBolcLlIqLgKlljWdYTKZhtMevUONYeSznryRkr7s7y
M2tDge/y/m8kvZW8KGx0osVm5uSZdvWozR5fN4YuNvhrFYTcdjVxEpw9sBaRlSnRmaGgRca606vC
ob2ZWPpqLJmQuyMj0qSg6UWI4LBW1NhIMprw0U5qrQu0p2FH5uYDB/weLINgt03PML3rRcMe1BUh
7z6vwvec++fTEiZXawe6tgXipKPFXvZoJmFvMS38S5ravkO9DD3/RjfJu1pJEKvm36ZofhsG1Cqb
+VZR8LGYWm4j0GA6i/97+xrNMCCycs3z27lRnYUSa4z3n13h0kVQJu2HF4PnxUrO+CUFIp51HLVR
98lqN1oslDXxIOpjZhfirNjZAjiXS7ESp+mqah1XyMsDdIPgTi9/Rin4CgAPD3Wu6NWy2LCuqa7J
ZWyieBdp4Kf2MpIrLEm24Y3D7FBhLJYd4F1bJmo/DJOv6AI/jadPLvmivNkDxWmwwiPM9Tf0DvyW
0VfjYg4osrXJwPoqCCFLMnM4UrYEpYd8VAsckDvX036TjSSKKFUS7Eac62cPfiY2wZ1u6UC8QOpw
y6MTNt5AyAHcx1sixh78idwFNq+J0NBhQezRtpwO9CUPbHSToHNt7Ej17n7yHADPbpEma+sbjAZI
dsYp2Efl5vSJE5wS/RnIkOYeU5x+wdHKnzdIzE9qpCOU4JwTp8EuHT8ksTkMZ+h6b27NPOex3kBm
olhxNMf6ofHdk7Qu4YDh92s9FBr3KUn7UjErgzyOQl7VmiE8GxKD4pQASotdSHXh3uKnf1tmdxqu
XguFxQuZ3AhRwz7xnHXqsIMH0BBjFtj/Svs8qn58wM9yenEIlHMC2f+igDYosk8ayWw/n7bRYXfu
1yqdpWH7IlijKVJ4oRMUG6u5n9mF80l6nimcM4nnZEba0YCkhOSOfI2VhJDb+FBPllBRmhJncdeB
51WqZhVh5i2d7SxLlMcArQ4NRUkuxWzjIYYu1vZW2GjeUAI7HBT1GBOOmCOzAOKG6hRGC3i2Jy0c
8AOkvfCG/Rv4tgYI5rIL+b2uK665bPXVmRbMgcF7YeV2U+Y3KM45tm02A45Qpx11oX5iyLyBS+hj
WutlZQR/IE45awWStHmDxf27dkodqbvZSzDCEBf8FqsBWzm0cLefcycNkx5Goq5spK2QBhU9Vbkl
zfkbHKgSXbD/ciSw4EpNfpNNKY1uq84YW1UjTbOgVY+g8JVy9Uk1K+z4BB8nqp57fZhBB/HUcWia
OACSQ0V5v1pz/sGASbMAheYFfyXKAnOcWHJikQIaZc6RM1pGSw3YXcn8hqLX9I2EUwlRA22ZJDSB
WgUqvp0ZJwYhZEtgCAlrDfTIaSXBIArIUCbs9tajV0+BmMyQ8XnjzvYsTownovOg/fmXDmqmBNjK
5OYrreLzKECDC9giUFpnTBd6GVPUDS5JSXOWEkuJycon6PE5GRPqizlY9rKEG+5qytbfdKHu4wwM
H195upFgTMlaN6m71eJG9lu/dLoix0G6mcDt6lf0Z7tPhD0L73Yt6QJdTD1J2HEeL7vqeIf7qEGM
3wy4OzHG4IGSvdXj2/T3lc6toz8+gOqa2EwuubxhjrnK5ZTKNFK3M+R06b0D4ZXsrZUbGraQJbwn
hRRx8Y7iWrOvsNU9ARKwV3+Kqe2rBsJHoyeycmuBD0TP1ZuSkpJitgmkCIdixwSS8Yyq37WTknP5
0YKdQLJjGqE2ETHhXSUJ0NUJUH5afTn/j+fzUgDv+hofcsaeWul0tJyadkVAFmL4AFf0ELapGi06
+vqH61A51xrLrut+DscA+dgtMBUBZrpg0V0Aj+HpglvzqN9RbwnO+BOPbNV8t0cK0XH74Oq2wrjO
YQJNSWsduATOZUpI7tRPq+1d1OLOGjPGCbs7J/047bJzAl9sQFVron1UPhNy9p6e18iWNxyyuzy+
dBS4dku3ABNa3AhbMAJuPjLNZGT4qlerjKqX3uBlit5WP6ZJWJsoaI39OcAocW+S/t0ufvhkDvff
y5r1RaG3ZpggTOLLAikwYZxHka8iSYGsLH84BY7zKpco8M/yb5p2lvNXkUfsrjlkqK8YwkTkzIKv
EVh8K8wCYP6sUJMPpaS/pPl6gkl5R3NJW3wA+i+fMeDZWlKVdXbhfteYm4BZb3hMKlt+vEFZ1vdU
5NRRf3Gw38M+H8Amna944sKMD1TGAsSn59h0sawiLnRq0zDXqpkR7+hx5MxvdYgMUQDEdFdU1xTG
R1V2NXLQFbstXb+GvqxeS2c+eov6yT9wkmBMbcYjioo4jz9ICGaGO0ZDfGSemsq1hfcRgKZtSkHk
vmd1TZLPLMYvR1FgUlLlZ9BghAVOLItW1p9FG2aLyRey59v+VXRA44biIJeqy8uO4N4J93UZm8ro
oQh3Z5gDDwfJkIxuyGQtd2tNlIH5XkQrKneiCBHCgMsD33QD+2TL9IfxM9rfauZVqO1a05T9y8CG
NQGPeTaAVj/ArmpfpK6flYOzRPAZ2KOVNJyvR9KTlcVBkjxTG6vz74UpI/0xyf2kxVdFWxgABwkr
2Ccj0o6hirlx55RwoqCHC3ybDmc2r5j2aUgFYfDx0yiFeL8eR7R6aqzr4sr/4OdWbH45UfePWlXT
HqKPFmFkwQyHxn9uDv0JZVrju9NDP/rjJuQvhlVnetLe8LmX5JwqA6TO2U3m5gqnqcZ7keHj+rvR
HUMAF5JrZP4os9miAb3lkQJ59QZ6orXh58bJAtO0etjSS2wSmJv7eqe1CaQh/f9cY4KgaiSWRWaC
pjXHtoy9zFTr1751gK03wYJg0jVkdcnsQ4D/fU3sYOrEh4c9Jedf7brk2W1V1sH1NgXuopBMxf+r
DAy/YPakSXRy9+Md1uU9t63u0j9T9Hx2xVqMNxzxCi2SU7LsXaqqp36/+8XQhVYTI37DxjlFnpG6
btbgLW2YzVEPaNGoc04qRahhSHK//A2dz3zVLaGXthDbPYoMfDZrBUTb5gAYBVmzYKLR1X7C0BKs
Wvg9IBJ0P7gfofCfhM1Jolc1Al6s4P0PTg7n+2au5mOiNMyC7zi9FwlpsitZKl1chzh/KCK9MXxv
e8lbOlAFzIig85etZeeZ/mM1JTnMm3E1snFpHrSz0/3xJq0VwGyo4S/DdVxUM1fDvLQq11HyYfT7
vWz9a+iuyHUI91I6soapTVmRtwxnKdbNK/uCOZ682hxx3Hw5tLE5ljfQ8wbfe4j+fR7/Omxk1+y3
gaFDSczSa8W3wp7dP5pkn82qPQPHllO9O6qxYCuIRHDuKtUmbKlLCFs/LoMmROoDghtQXJALyzL4
DzGOdcfnk/x5QAFxZeDucpfvIPPLOSHHGb/iJWPDvT9bu8MslrEFdzqFe/+LOQGOow4XpBfzDwhy
bw1HTwg59iruJ0scF3/mIQn6Gczc6S8MeMXXr7U4KKtt34lB0M6ZIK/C0gaOKa5TeHUYmzdItaz+
2AWEheD1rNJqp3EI+GRHwQtZhdQz9nKAgi9EnojhLD2ABqujk5XzBy7e42DVQV3ZqTIOHhWlGp4n
NiZkipYNr93P8mi1qTiHbPcjjqSI67MzcX5OKhAKJzLnOIfEMWj9YXsEpDonx0Zzv5rWUvedY0nw
MqYlNfp7yW4JYTTP2Jg+epJsVu5o22RKfRZXUrsQyPZmqlF/1rMBNCNoKHtxpk4YyBVOdanDNvWe
GcacdvT/l3yYHA3FOSjqSOU0ApUUYE4ycdz4Ft2eWE5gilQ9kadB2v/KhXAhgGy2qrssmbvsMGmH
yzgQZ9keig4smYk6X7cBMid8I7kBX8dCksv0YKmOx+nHzAnaCmfFtH+RkidfmJ/XsZMgNOC/O083
lh5jnGcD0MIVxIT8jgifQCEQwGs58ww2L6ZnCIytfTYka7VxJoqMl4WxpS9yvAjdIdyfflRZWfTh
CuMi9zPFU/dv1c3A+xaRpCkf4nx3W10FfGBPugz9LKvYa+6lFoutCFCRVNeN83bvt0QOGCDdpZEA
6kn5NCbl7I4SDvEKRiL0PMA+qkQwGc85e5JL0AeEnNhbbHL2/l4hU/+4dx50r8six4lv3aVarsnN
0yA3Li9FptwdNJIxrTAjJn0aEgwW2pIR3rzKDnPbcblEYsVdPlZ5DeXOGVcatmjsChy2YZw6in26
jeU9h7Mm2kJSj3F9UxSqHJl5DFEDpcXZ3MIoa/XhS3IL1nHhGobNHskOJVqaLuM2x2hhLxOVWErL
iwvURKQd9nev1GZXzwaGE42+2CG3YUvp2QNusixe0jAeVlRlEAma+XJ2DUofJa/p5ic/jP/dSjb+
iT6Ss6pCIu1p5eh93oMZ1kPektIRxV6Vq4b3qmivRx1sTFx1JAc7XFYymrn6W58LEmXPVNMI5+b9
d+NU8B6738/SzZ2lisWy9lt0f++7XuHD9KkmGLwqklxL5Nx/zS9fRb8dVXp3fe5SesD24iUu44Tp
6T3k1D32ixxHlt7YBMbQ4I0x08He2JlC1yv1MJq680Du/rxW3veEtbjoo0yHu3ZZ98EmfeXqdRfH
La+JUrfkUlr8W1+uN/+JzK0LEco/SaXJWXpK7G/1dHaNnvU1blEHZei9J2Ym4EIoZgQKyqJ6wWhf
kWovzNZwSINX/tm+set4RptQR4DEIGALNvaUxK3Im37wEKYRnubmXBVQ351k2GMA+Ze+On5S+XI5
7nhRZYG6Vc8kiMR69gNzum5EhjbRVzstXNEuMvwYmvbEKB8azmW6FgwkaAdtTMtGiNVPkEwaK8eU
qkPesQ5Fosmxph/c6ju0ElsMeDIEYipy62BhCnTh7exIZmDV41UcclUh74EByVEvjSMJGeGaCrRH
diif+MdOhyHgNhP/tdXCGG3mkTD4QnXo2+YeCb0QBOckeXBHhH/6KGtGG2+QfLwunOknTq54XPXL
ZtZe/6dqYAmT0dmnAIjvzNgmFskuF8QD6DuIcePUyICgdrgwNgjWwERa4sHfB3ExTypqWVrn/Qn5
ObsFjAcRJ+ATUK27DrKCfS/rQ1ZGhrmmDsNAYYletXNmqJDHbbrvQklIUPqwikSGq/wXrJKptyNx
tXqSxRYMZWHR+VksCgKF2m3cJX+t4tE7mwyslcdOlsPebVM5H72H7glKXkCxjTkGVWiQ5ixVgz17
AqPGZuKdKAWocXAWaCKIOMjmJkHAR8GMffAu1U/fv6SPOdPsdXFMvICaZkJ3yTJvzHmFHwiF6+Y/
Igc24+/m1Nn7iKHGvqlELaC+jZAARjaSL9YdvOYQXrinHi1oGNfzkjEeHfPnwBuoB48hm3dy7Cxr
n3ZyIjLarKc0GhGpt5F0lAAttoTUuHFq6XtnAC6oTYIHIUYpp9rauoTEGlVV4eFiOJZV4CPMZ0/y
oOFBEb10/hJ9L6tCd5B2513O7s4vymRQG2OypBdNUrafKUeZs+AdLAnCi0hiNKQSS5U2yOyHrTxl
NFcrnHQC7sMAilZi2/UQWJL/P2I2ESZ7DsxkLK9MF2SAMtMLZnLgOpommr1JDFh7e1WKxN5DU55Z
kCR0r+5Wb8rXtKOJiOrnlLGq8+brxsXZn+reODnGTqkb2uwKx0jc4nn3srMK0fxLXZYwyGpbC0Dc
t4L8VACI1ekUV8+lUamL0yGepkI8R4qnWjfXUSIUXf5TSKFrNE7+FgHYNQ3yOv0tz1Znpbbg1b8T
XNEzkptF4SwGS1TtyDg2vZC9TUMvUKrL3S5m+F1xux3oQPK6bgpgsYfFpVF8jeaZIYDdlnWjs1Sx
2xWUY9ji/KDp7sV5z6RX9bnCSQVwHGINtTxM0dT5zYiiCJscw+9qgfAi6xSvjc50AbetQ6rWpI6r
6dTC46rP6sSF9vGM/xBTg4eEuJ/OIuFaAeUwATLIC0d34pB2eJNBaWc8A5dXg6d7+/kr4wRtrSuT
p4Mb9YUaRl1XqXtIm1t2+5yJdbuwlZja1vFAKOY7siQpApd5TNC9sBd35KLBvHitJ6+WVzGHHYmy
4fjvJubbEvus0otj/kUJXzwMvW7kX1sbgS5CsI2930lrGTj8EGgMhMityCjNVebLT1ut/PoGRWfG
a3/dBxxKRtwP8NDI5QgbOvce/VT/j5KlOsGanQMHrLT4Xb1kg/RbST5Z7Obz2yytp7Rkd7xsA0ER
kIWz6sMj8LFuDzhqppIgVIb1ptqEyrrSJzpIcWG2CPmuxwe6eFuTR+IT2xIvo5dzxKsaxy3tDzhf
fpOXCdhn5OHFUYW2gCx+LlkfyJqqQDNhjOfWfXEaEAsSusmt7ekL1TqNXADbsv/2ahjKvU3tLhlC
0MJZkMPuExVaYxSHtWztIKJdKiDTrAfCqr9N/h06qgs6xDy/sLWO9lWYaOEr2djZEorxOWi99Ztu
iXoc0/+s99p3prDQYhXf4UphdYHH5UOroOlxdKqKohctXBM1RH8hFIJ3MmagXfdgcsQqOXZELdzw
hzwnNyGwKar70gLWPADq9OJd+3d8934XglASwuWrxEyfiTFMa0SqZYWS5+8baxMxZjXtPyF2TNWb
eT4p3Le+iO2sv2m/hPfMehpTjEG6JMirsOru24baKLTrbnZhnPM4j1zz57nAUny8p1q3mPuUjtjS
IJyRi1hP0aYgWW1Kk8TlKQpbgnCeVCR6hgw1JRvll7ljkdI2hMqm4BxCpifOpQm6UOOBhuqLb0j8
VjObOc1Z4wziK2cnPvIicJBT5a+DGSIzdUDDDFnVkOzmGGekf770oDncOwRCTAeS+Uyx54ZfxiEI
IMuZ+CCt2eYcyylsPV+ftNW7hq1X06ZtacTc8ygTLaqeTxoqOZSlyHnHRQXLTUoX7lk9Muf0//Xp
GP1EAlEQZX8jYK5H1Wem111kmpMLO/o8pUG7xqpG05Kmrs1SwrLpUmobPNARJoQd9Hlc7IuymlVv
Afbr9HfFzYnCUO2mhThNTgiMgYP717mF2Mcpc67WtKIGiW0I6SU+sHDqF6Qux5sTt3cA3ymZNqqc
h6e9JKVlY/1DHlYbXVo5aiFU0Q9peTsJy+Xu0HucRmGfaF1ENwEYsrIFUx0SfbZcFKWpfeza7kLr
tjbTLlTbhd2k4phtZ1G0z2rNb/KMXpk1kXtG/eIipD1GtiLvlCVcpy58QXw8+MiPqGlI5XPXZlLR
bcf35Zz/Y1SYGHwxkEMfRY9v++KpSms7E2CG1+aknK9LdQdpIqK6WpkKSzPsn75jUFzMID1Pznxb
DepHJI1xVwuD0Ap3BCWpAkris30By48MYFJAuH1SBX7cUhrIAms4ferxPdZcCtQDtUyCpIiI7CVN
oyZajIbMb38aHOPMlszwYO/ebvnf+7Me9iB1RUosaSp+gY1F0hIKTTckWTis2ewWK/494KTRM2L6
b7RhZJjJd/l+x6xBJlfdGL51Fi/3hgzNZuX1IhdkztD+3SE4sBAbqEFhuWR0saE3dpJoRcWSm9uv
nRYfcknA1bw2aAQ4UR1FUjn4J8R8uYuNLx9GpZC2scTQ9fyhcJnaISZk3ym18RSt2c/ixuUGJKYs
Zt0Gk8/GEaQxRLFKMv1v0tSPT2LW/yMFYfMcu1hpaOvyrMGd9DTLlt1Hr+2udEO1NGJwyGI6nn2M
AZPn4p4ShAoZt8k3EcNRPpz0jInNHekcVey0Hb1gZGOYoKEsmMea2c+/TUbZrBF3+/QmTeYa7tV2
TwL7KBk9RWQ6gviGohjFMhNwA6xSPlrRWuRiRCHhcnL4GiR5QdNSf0ABoneTZ5075D5uD9UuAdLC
EQhsfl5r+VnksiwlARGEcbfmso3MFEOiKXOoLjH1DaKJuHl7mrGN9h35+nCcbAqcns2wGUF3qO6V
iefCDe9TmvRFUVLoJdvwiQ34hL2soykxeTDlhhiKgkRiBw8Z7YAxmSlOtArOfFrgpFbcEHJ0pF8I
hZ1Kwmz9/OmurWFIJn7f3u0AFGbh1PNmq+N253Kk/wNZ6zdIP7DZqgx2XskHtOJ3J6umlOCojkmx
/utGDv5vwLEB270vZgiR8m8VSJN4oJRaPBGW1OyaIYUA4QFlYZ6shKljr1cRrSOe1NKgnfiQzdX1
SCmMGvOZh7cruZzNUHGD2OYRaoG6fF6xS6LOIMxM+wqzdge6x5P1aXWcVEr4B9Ccf1HEfC/8KhYo
GgmLpX56D0pf1WwgUKlF5OeD4zVXqkfyFxyogjD5JsevVME5epq3gqQ8u7BEDcQFc7vL7pqHLGyc
RfMPBINgZyjnmt5Jw5puaanhVkqN18yhMCJF9t5A+zfVN1WtrJh9pDHNyeifyELs0s0en7w8OiZ4
2yRzu3UHJNOUl5GCcNm7ok8MvGWubxNj/IKHGAqPmPNvvm7Xi63dfxqyttqGzpuFJKRTV1bPSbJD
y2oVGIhqtx6ORsCW3QzvK+ZVYMo5GTofJmIlSJsFf4PlS5sASRYiyNjO44NXEaD72a3OR3qvkvAB
4ay2CjNIN1G0RzF68D02CYa6hIQ4qZMZCC9JB5dYZQEqTjZUYJbZWYp/JXxTyVY2fnHWNiKZRq63
5D24TdifdRExyqnHdrcGNxhnLrkU3Tz4AluBHtUVQcQHBE6ZPDl6c3Wyjrhjxk0R4S1yI5vORB1a
tPzUw5wqciv4w89GCJNv4G/abZxXoim3IEjx3ac4CuK3vOSWu8eigApSkle17wFyZhIWlIdoOOrs
r+VIotD7xz8jntBWlJx21cmm2JgMYYAfesaa9rFPqyogbk4EW6C/XYpidnvdOcFUUKGb+zli1zWK
c3EKeFV+uENjK7v3o0OdIhREKBhDWBNZpWn7n9+tuDzYvYc9dIRmRYox5KhJXYoMbtBdUhF0ES4H
eQHphAdNkboPOjmq5/1IADmY1WZ5VrDu4+cGuN7fejQ+2VoTwAa1LWk6KiOkcpTwXGB47xXmunhG
qy3/q0KXDNb1fdcK5djorXYIYxZXCv/X3bOfwkMzZ1P9Nwq8MTSz4BM04QYEHND/sYdwN3MVHEwp
mSqzPCkPRq3eEYiVEwQqfOSQqoQEuegpBxP0BKL4hPdq1c9aSLzlBu8LkmyHshJEBAcuysyuN8+X
06HkAJg+GXdDd+fnQmWRply0l5Fe2MCcmMB4C0ZtuskyhO0q4C5uXXim7SUvfY+j0vDJUTbCPjiu
UTMM0xYc+YBNI9iPHzCxgH7BvfuzUvdFL3Le7d36J0DtqTFycD0FKpiB8Kz2wck/1IHLiX99MWHO
K0mIKRLIsjiWC8zbi09WYbxedYhd1Sr65gDUIlEpUdZpMn7ku/rRhHwf0ivyUqWbo5E8TgGF3s+z
3IJcCURcAlpg+yRJ/wtwvl0NSw8lTJoqYSp5hsnBWxQwqxTJZZZJ1pLb4uGUio2+1dUmJQ3jRuEv
PUTKLLQVmwR3wLTd4E46FvuscM5aUjAO6fH+c47Yz8eDwioL7ARRwt6q+QXWMDpIDHt2PPIHkaYx
0AOg3HHgw12zM6bEJimlib1PSNXiQXHnpm0MBzI/jfVJvG1DbTxlfwOlujkf1T/TWp4FrHEHN7UI
BIw7+7tqPri+z+riSu+eqZqFOPmDE1+ViMAg8MA/6MigUsjyJ7mtepSfXGrWZqeksxROgYXAeJm8
FQRka919JwhvmOp0t/Nhynhm+GzZrNYYXRBuf9T+0fAJrJRZ6HqF0ntfOMCWsmFNVep/FSIos5C+
kBGYp1h/ENVtyPLP5yYsxXLdWxGIxpKDCD1N1j3SdsRLrE0HPm43z7S6IxqxsAqaiT/bsZ/4oXuM
26dY2wCt7WveyKE8iXVWPz9IuIC1R/xidj9CoP4trNYehFQIJ+PlXl2D7DHumdvUm+IWWmoaWYO6
UThgXpe7UYWrMJq7xS0YGh6GSm4xBC+p5fAGEPg2OoYNPyUYqmK/YSMa3jpyAN8IkLIKsXhHRj8x
nc0OiKuEmweF+9YGiiRmjTJNxqUBlpYNo5bBYdr1CJ++WVs4cGkFXOuVj8RhFbj6Gu1HfNoTw3iR
fLsLdTwn8eG0LsLnW1anjVjNVLqdsUXie4wEtBSQg9PHfpbI6rtvuqureDY294rzdjj6dbhkL9SQ
mqoSJYps0L3iYy0LISVvYDQPrRMQzg3nIxNVG/DS86MuycoGkGZd3vyPc6M9Yt4x6PvTyaUMRo/C
L2TNzP0qSqQnI2lczXmZ48/OSL328isiQoVCbWRkqUZmDjwp4VepwhuwNP0RIW4GSmyrA3vpAR1G
ZKsQyrczpbA10gDfjN9rfU/duWiVIQSk6dJGkbVnk3e0xWSAIccxR94OqfiDaqOWeH8ybrXkNXxs
GkMN5l9gZ0s5TJqTDd1KnLW++w7drXP+bjZs1hmjmUKCyE6YCzlnOw0lvSgkIMcMaout4jMt9E/R
k2+2qBE9Mz+IC4GYR0gbSWGTu+mQ9M9yCv9W2nI5mtjcRW8/4tu+OBkB4jNy34kPnqyiZt1Q/DaR
hUEWus29GUcm+M8O+VzBpZXmuPc2XvxobRIfTKr/al70TZZ8GITviqofiMrnn9pb+RBWxfZeHSme
83cTiVVMjLxOPr7XFFZsFBL/vtMpK09i1F+PgbLaS/T+FPlrn8Jf8HNq9NuVrwvQpmQPPj6ACWMG
xjPB/cbrqLxl/xrLmWDiRB3ztOwlNarum2h6hlogsDPNTPDfpQzCua4Cfd1R0oEQEAyBnMhw6m7v
3hO1MIlvvqy3nt6PE39zUTCK6DBkepYCfg+yqRHVDNbWeiBX1LMfGs2wsJEi8OkWtKXTt+vDKw6r
4YAjWe74pya6NLmbsnEmdfLKXjlDUaKpOYczz6IITnXbsgnmjbdyeNbiBBjcH52YlIhrovyfD7Ao
kGGn7mHyKzJLula1+Ou6q+lFSlDcbLf6mneRtH/PO72Jd4BN1CbaUo/eopw89TLHZ+4eJ1h/nAIH
MDAu1mTFvrIpfOR4noh09m716hhvGM9uO+xKUmeyM5TJBMQl0EkoYidetlBxHpifHgTlsnTltpkH
4S+GXufR15Zc5oINkR61CMEpuyz4VZ5Y9vCjWFkdy06XHk+a0nHwtyPYkNZ36s/Va3E/TNbJy9JL
zghaed+3/6zHITnqN2RjnFfAPEvv0DJy89cD1ik+IPUgg8agbnnaTLb6wTXeZ9OTyhv6gTt1WCUa
Lh9zQZ/A5E8KkWG2bFzyEXCfBJvh9JT5ma/TBxodzkBZ8+bLO49ns0yUqyq+AyctwA9Qd7T+rEVJ
E0OaEJ5C2xw6MNaf22gooviGFRFhuunwVkAL7qfrtEoC4B26fCb9BkkHiYRBpesgsJ1VMktIfxeU
UuSd12s9alpbYwGcaIK9cRiMNSGFBlPhzmyKLBzZ0YI/X1EDUFHXJPxc4bMla80nIRzSPsELgGod
U1emDjFFUrpuWsAzw0IQ7JobEyjMwZWiA2cmByeiJfOViLNEZfA+aSIOszBSQx53j5yQjgpGfbrA
x3XjEzTV2w3OpQTXFeet4hGRiUU4ID/jXUXB89++p6QuYXGOsZMT4rEogqOn+ZZMdB8hTFkmUhOq
JsMiMX8gNGq2LfDgyvRf93NClijxUYMNe1N1/If8HmXbO9w140J/1jBys7tRBgW4B2Pk7HGPv695
2J9yK4qwRTeXuZP8EYWk2BqYVioxNS9guf+MN5s5eJtIUFhQkHbedWUi2BTe14DbK+lxe1zdzolK
kTBX1Jykp+S3VSf+gyG06wMZP/iXgUgV7hm5RWOLMqPcl+oIiozEcIv2moOuCLGGh3E9DjHx7hOm
JlaycqYmLTNUBgUb7W1NdelYXXip3s1HFCr2iecb+Qiur5aAX99bkk1yEBjgRUzn7LTzCsgIxs1P
xSVSRZJgpXgRsFn1TJ2nToMQeWUTF2gZ4dsWVJUmmjaE3FMEVcIuFjRF4bVoDWBAj4XP+oaxRVi8
FSn03/paz84pw5LsKzphr7CR3uGy5jOeF9cRWOjOBsADKanG/cdhLRHMqBALo+LNWfo+K67Y+EqS
atfS3Br4auo9wZ2mdTyqkKNvyUEavUVueg9AkfagkI5yk9xHo/zgKXscGT09z/kzhlIykZTqXxei
i2/nrW84UJ58oIrFUzc0PBkAn0pD8PI1KExKL4elHsPkwlPTjGt6iaPzXIR0dKGf/AH4g7+++e/G
Omek0Le4S6/1J/viKYWlVD6D3VTvI/z85cXnka7Ab+m0EdxmfeZrDsnSsZDmqQTHwhakmzEAMZdq
Me8jqPDOtgOgI5v60Zd5dJc83vEwp71WVnZKMaCXJgFQ3JKeG+tsGmEEw15M5VOKWezk5V3tYE1q
rBudGfH1u0w8ZmmjlCSbUB5SmW0ndIUZ8AkX5UGFmUmtYBTFQx1aftKUPheEgIh078gP1jUUPLrO
4iAcAXKTMHky4FaF7GBsgeYJTavh+kqgRG15uhTIwqokK6LIqQ+qJJA52O6mPuA094l8Gl1AuIXY
yucHih9iM5mbcha92BUAykj5l9lFPkILm0lYfmrD4ynkq5G4na2MNoKAfzajmUDtYe6dF+Y22DRI
ZvA11nIM8AGF6fhb0jJ2hO4tLuDKkFMUY9qJlWqUUoJM1jLuznTSYvPzpGMog3X3NTI3J9M6DRRT
3+A/lR7SrTfWD9K+jbXfFiPDdEQopvBdHhdXdjgb/il/Qc1nFX9N0hi1EnKs4IN35ujYVt4oA0hv
eXWpDeWBdTwHHs2nB1DIsJS0WcCP006b5z7FEEhYTxyszVgBvEQAh5pZsuIgvY/3+F6m5UOiWTUf
OU7ujXjmLsGZvlpj5LyFPNljTW+sqR0ATsN3XgqubqROdx7tfQvMakPt7PqyWeQzWGsCulnWsAwx
ymQD7xHopD8wNyrOQOcEv2PUHRdIy1FlESiJb9jCOxXWOXFBPRwBR1eh2rf+dGB00Xl1OQ0ti+LK
zYWzfehpILTCHHLJ2A84cej7xs/WLudkRuNMryC9nyFAivnMdXcQdQpTPgLlXDuEG0Iyjy7N7DRx
JzbXv/mtyRbLb3wAGHjqgLMhmVtT7WAft6o1gu7CCV7JheEbquz/HyXSAyJ1aPKiwysl37iQz2yr
dhX6FLTEyo8eNysYWLW5WsqkX9Gcpw+ivxTg4ujnMFB+DM8MmVcDIRq1zeG7v+M45m2qHePVxFL0
tud6B982ls3kGcARyy3nnkMN7yMqnHN3qtsOD3CluXYbaIXpWrsjjEg3kj2c15N4nU22main1iP+
7B6TW3VQ+azoA2z4cjrbog2KFQ9MHbOaBae78TtUMpKABaWVL2FZqTB/FM003gbiSpF945jsD25Z
8nUu0Oqkc9JNlThiC7kNPqAst7jHBO5No1oC+eCZcAUkpHCYK2NMefbuAW5px3cbyUZUpfdWXtGm
xkOEgYtaG34xV7yMhcFsEKJSsuMcylKazlZoNfPF3+9SS6bIfC0IEU7EQNzMaAPt6fAJvBNug9sA
/FlFbFbtUzJY2CS0D4ua2iIYGChNKhilaAALkvXm6iiHgsGg6NbbOBb2QIlJYFb/P2i2cdPeAZpM
ac6sz3j36al3Pd3MyT7sFRbFIMENhhzA4r7rYoNzSlnp4O4pkC8yMACZyJhrl9wQhqMdhpIHDiI6
p7LvdBH3hpTiV2PBw0SZ62RRWY+nNHIuAR7BjAIEvf0+hJxPRUI1YyszvwKUJccEGX7jaIqLXMe8
bCGrGP5dHw6O/2zOxHZO62OW1ueMd5tIvQ6J8MnzP9rYS2fbz2v0f3hSG4FPcSv8yepnqFgIdneS
Z4K0PBhG6N4MwYo7Hb1uzPU0XvswhUhpAoXCRz1rTF8r+TmRkWGewFXTbkZeVt3Ynsj+JYBiVflm
BIzw6/HEgxgnyf/AoT8+2f36CkWbLhCoJanxf2bnxTKvcMkmPZp8bkhuaAMblllxZNebmGY1Oq/G
Y7VW2numThQotDJCRCgG3zTy3gtFuzrtiWN7VTYZ7zITGnpALXnC6lJAQZw13wsKRRD9LEgxUY0o
dkgWkfben1pgm6OzfMsvTb50aJPNVu/KX7fgaJokz3DrsPsIDOgZKbJsITG1jlyz6uTfaltcmcMT
0ccr8p8KChkh1SNFOfBHdAh4VsaN2mUPWbpEvl5yhoeppp6j8wDhVXuCKXWhD1TvTQkE45KifMMy
CLWjYV0AHhJT4iySUD7u7JE+nl5oRogMyxPZx0a/fZgFJzv881LbjXmgB+ZRCrUG+whcDqwTXYiP
DFP8P8iPvvBQWgxW2sjVlxdEU6abczJcW8FtGJ4ns4Gc7kwyFR/euY2CbbjUAIFmfbcAgO6vVnj3
yTXZPYrpld1zDKWvuSRhqHp5YtNov8gLheLw5K0VlAvze/mndKiNQdleejkL6HfQyTJdvb3hHE1/
COSq0NZWAAOOTkf+seY11EztxNErFXYLJnpROmR3o/d9v0kccow3e1hAzkwEN2i6UvTtbYJtQiQ9
lAabPlStVY1Rzjp7ZQF8Y6rlyvRa1EA8eYkX9KFBrGHgDpOtvehrw3tqysFYtwMSE5p2discR/Rk
V/cMUo5v8qtG1CONNi2vn8/O64pMpQXiARkPuTBp31UUcTENA+LHGFzS+v2HPZEodz+cK6f58B/a
wRoutgIFxgCh5FYOKlAGGhSsMmGj1Urw4bhg4Jjq8iBSmAqKDhTmbn/KrhKDWBHfLMcFROvnTgS3
Tsh5SeAWn1SUOhLiHzXyVl5GvMo+UKJeSIy/P6DRZ5P3Wg2nrQPtQbEnoYB67gLh7IHvSc3qMsi5
O7XrmRz8mangCIp7SP5wffyT3S+Bz4Yy+YXnA1FaxtQYa8t5yOVfZHxwJCws1BiGVQWsKIVkxBEf
rc72IVxtK7rQWnmtdO6gHYCHNy0VYmdpkxS/clW6Ai8n+2MOwyfsjDHBs/RXAm7I7aVNXcKLtcmh
CjqS1dkHH1B5npHk7jwBMzGPe2Lr6CWs2mj5PIbQUUMPao8pyX82S2j9Wt1uerN7yHs7yj/LPJB0
jcB5imXRoeFzLW9u7Bx/9bscpINXs2S3SdVM9nKFKnggXL6PXgdoPaDNg8RzMvbJEQPrXvkASywj
/rNgf/V/uWCq1wgnUWhi0wkZ8Fs8e+bzv4XWeKx4s46pMK4wnkTMZaumN+EZEw8F4mgzC6pg4jac
Kcu1w20r3ZrbOztaaXEgOteRWqzFA1OtBLoy47j5+fvtRLgNQiIYaZBcNc6bXeE/qgR2ahmjl0pD
eIAiR0yEesIJWXgi0Fn2zG8ho156m8BVgxmIxbAwATaE1QwGNd3++iM1NjkaoHmT8/xK3pckUveV
1Vd0IR2J1N0WUbbRJovm59t0XQIqqaC4/bfQo6G3ymnD8n+5xvRTt5Z58TawAjwpy20vBXkXWaYT
hnb9IouB82yuiw4r7mFSmFxl2SKOHLNWNtTuHmUYoJHE4j06wov0EQC7jczWRNxpLDVbrha8g7MC
ZFiKqzlSSzXiSIq2msImkhJTjvOokGj4Pe2NkrYWaEmFBFhNUVuIPD52CNXMaInZSFN7PUSZhDXj
WyYsuufiPhY7ccpB5AZBAYpLmWZZ+91v+6AvOjCFQ0EvE8jSr+RotE2lv0Fpt9tdRefrgYhs+MrJ
+jZOjGFQ/BZ+65qbFNc710/Yb1Vlifpn5V0TlEvy3vrr/5y5QbfQ3gga/yDoVEO1QCsUWMVh25Vf
zL0m/gv7y0UgmqGNMT3AnF27/ZNRSMc5W12Ko1mb4HueBstE7Ve/asSA7poDGTsZ0ew5miqwVItf
9nOuw09jtbaQ1Z2lXfsHMZgAUtFbf6PQFpRL0KIt1t4Kg0QvurakYyUr6K7XeioO5WjG/aaFHuMg
WbsSpVwgs0CxskQdw/n2TI9yV8xyPuHuINKYqgH1ka3+eVTtXECyduKrhSQuX2RVOppdPx7O6Qu1
D592jwg/2Z8NlRngAVCSOfHsuuSz1xc7ZbqJH8X0RtDm65/wL2dRFSq6CG6K0qQZcPvpF55jZG22
gab5wER7whivAjbMtTTKWmUJzRRYaASeWItx3LTvVb7U7UsOO5x0F7Md2DwjU0CBFz6df4g3B0MU
zd9GzzaXLv/40YPPb7IF3crzQU8NCBnJk3+xQYRrB2LdlEZRGiHwTlxYHCbRhne0ZfBYpNUxlBFm
KGGVxTnM7fij9y36v774y1hcc4vCWVsIy+prYCp17ToxfRCQNQ6kQqVj1LCAVW2XwiX7BjRzCuag
5iPdJzLjY0jGA2mt1JDIwqZ3HjKPBypKUPO9Je2jRrMtBLdZVsnnhMonxQdZ2Xz+9P7jJLoWik2V
Dv1Ci8+VZcj2Xr+cPIYHVFMhXu4u/fZ73Y+8igBSMIghxv/xj1hymv+tVUONYcR40KyIuRBCnWCg
cg4EjtNSTtnjq1DMZXgHEwr3/BFcIwFd9KtDgPbmkX7Lebv+ZBBuF6GD/9cEDF4C6oYt1qgtIPzE
z2Gk2twZxoEnFmdkwJyfqH6F/+HXmvWRJlGLjgzRrHKBIMSrI4pTd4zMeTVU03NkUjTgk56PdUyB
SqWGNHlD0rbVezr7BbCRy7w7NxQWTjVbr4ZW//BSbXAcjiWTKIekR9A1/NwseK08EIJeNFTb6uM5
5LZYM6SAoOTVEtIYwn5kBtYMkmhRbzDBNRhbLytQqkfAcFPeWNBRSgk6qn9RF+fDn4try7eIE/xF
QIaRYuXy+a6wGdaYlIEGRQ65psSlHHITgh+5rTBL8mnw1Hc1cQ2GAXIivMDi5noEzZ4y5dW3M+i/
vIPuYxlKJKFJ0xPG6Q1RXEtMU0tANVY0M+rFcmoA2CnXEEUnoKhUXm1J4JzqFoa6ZerzwtmAgvTE
GH0cCpbW/BVIaKJnsac704USLHrCIFQPfVGa2ANV9J3mKz9+m7jcp1PGXnUIY+AnVxVRYornejnH
5hr5DP5uMFTeiEfCoxM9+1AbqW2SNW4kdo73cocl+TJujAFQt8JvOg5YvLazG7Mm//UbW+h5EYyw
ddfVwftTcrAbWfi5E700OwDd1W1n3M4kILwUFeJEiSKnmzyoD1G/PeHSTzQTIFwrPaYO5NJzmhEg
nO1Dhu4udP1ja6E15t3dgwetOQVeGYGkHtzh0QiN8MTsZC6vyqtqlzP9jB+mVgoMUdDw5WCGv8iI
gFO5TTI5RX1K+8M8s5EujDyG5YHUvzFQoK79trlSvgPU3Qpj2Z2ClpmpvVhBr8ytUcWtEeI3rHLh
1frVsvbmSqeaqjJfY0xioMDCNIHUHhYMm/G5qLTdXX/xeDHRVVpL+3GbOVmOVqH6ObwlYRl/bH0x
78xyyvFjsVX4rmPXAYnseGtjYD7jQSdFk+Yrit6kCG4x6VcV1rUkFWk2GHnb7cluvgFuleqiRat0
JAyxqLAw5ft4B4kURdtiTpw/IhFr07SBHB1sFzpzc9cqtZUaemNVQHpphvm+SYcdTw3haplVh1Tj
5Dm7ex6vQn6DMg8KsnsA8ZjusMSoTso+av/hgMoPZDUmu7Hq0NVOBpLFk12/vXcWPhYbK0KQUzeI
TiAkufxFMAkcuxzouB9Mtg7fF8L3KcRsWxSsDwWkqa4b/u5EeTAdR02c2RvVe/yBG5qlk+BsD0Cu
iKSD3QKjZWvBFXmRip5EuWSNtI4Fix32D/MOXMJbm8YhFwosHL+2ditDYBtDEr0QPB8Ojsc1BGRH
wYHMdljO6rHw6UtAW6oc3LmFiPEE5lM5LbnpszNwiGs51wMoQwnLlye2qI/p9MmfgOASYnNW8uzi
AkU3XtlzTQ6ag6hoxrzot+z5sHcGlg0YydIGxW5Ou5WpwWp7hGYPctl6q+C2VUVOW7XBGhS6Ctfw
vbQJZcmFIBp49lqdCVeWFC7DYbNQYrp8ptDPH/+H34Bf3mCPpU25KSZ70UU0qzzvS8iL/gLQYNLr
jU05wyNw6nNCngn5fWHeapLOYOtfrN+J6QgUFpoWb7h6oLT8lPPP6Vt5Z+SoSrlgjP+Jd4uP+ppv
P+y1yQnWEXumn7UQ4Ik5fwoJFXTK03WYuJAElO16mxywi9yfg1vSaAEFgrqS9ViNKhqY4Sk82U0W
gNhEfH1/xYxvF16CXzN9Kn9RApRDy3rBUwmUwYqqXzFOMa4rvYye+ukrLjMOdgGsSJojfMavudSl
oGh55CkdsO8cD4FV/tW6sV73jP6CIkIqG1a4lBnCmE3taNxa7pXZscg0noXkphOkHCqI2wQA5GIK
ojNITKawckpo9yuyTM2zLvg8k4d7GKde6phTG5UzLuxgdI80qBssMi3JUIekYlN3UryPQKl/mgli
V+bT8Tp5/2OatGncYyTGtSim+esW7HZwHoARPIssKBc4KkF/WAX73cvuqqaf+ztJ/3BjLC/wFeDc
gRIiWn1gQTijOk0yjnFfQF+eAWiYuXf0A6+J+iF0cvW4wk2plfOu68/ckmr9hm2AQnWFPLcz5ydU
llw1G2W/5MXQ1vehlIdG8HJXjVMgymy4no3UhB3HAcwF1mzCsTBrqQYLT7noPB3DXrOPiRl25x3A
4uisE4wQkOgPajiN56F7fcXrc4qOH42GsrIV+oaCQMibBA+Ln6+NbdHVjjANyYvMxj8OtbZ/epwM
8ttEjfCmj7PaKv+8hNWZ7NAtsdVYS6CwwurWtiFWc8QXe/CwenSnprJnKEhYbFOpTJjORAtYARzu
yAs7A2olv1SrQCLiJdeyBQiBmKPbHusOxxg6XgJdDkot9BUj5uOIQ+GuOWglyBzdLX16UN4rMyV/
tv3i7gmG0t3CZ5G/cqHi/DGcVeAPcuW2A8N8SNiRBeyPmoAFuIcDQB5KUBTFAAixwtfsdOZ8J3Z4
+vxufh+zDn/VzoarF2E/EvfcFUdl6xTiWJ4paJydFGiQQ6PalTvioBrUGONAlKOthW4+yQUF72cq
QlIwyGT7NBXLdRv+Bl/cS8YxuBRghvU4X8joLTiJCtXFzUlXegX9QeZvI6Wq8TWYVB/0Ps9o1eJm
wRqlhp5t9T/lAhw76Uji/QENn+Rp9snNRZEfps/pbF7Q/m6lqRImcqxZrXxuh26Oi6R6GUQJozb9
Nh7rZtK1xvVPchfpBs0+jBYaq5/L1rcDczRNqzNXHx+FGmM9ObTTED0QuEFQpfBjRRTLzJCW/r+3
8YzWjdwfCTUtYXrbblIk8F51ruXps08+Y6ycsVsyjHU7xfQ78IZ3DihSMPETKXGsxsrjl+a8Psfj
XR7MgH0KNNHrDaqyZ963xEJNUkr2Dr+QidmeZ3mXNsKhJyilJgO68mUqqSYIpbPgSdAUf9H1/Qzc
pLHR6gWa3Q/jHjE3FeM4OHJ0xQq5AUdc46AAvJBQlEWWZhdZ13BK0NXqusvWcam0tWzB8kKqgWrR
doAizhnv0YuxKzcoKS2hSjdQ2H2+wfuarL9yv4WtqZTgoQQ2AnR+rQnpqDaQXob6eY7CKvCh9B7c
b6lJl0NClFx7WvHyixNad7znb2W4puRyT/hsUNAk6aEe8ep2jCcdQCGA9kNPST+Cf3angoy4ZJZt
B5QZAHHZUEvyVF129ek8eFR9T4tWvbWGSkSiSexORkx2+ryJONXt9FwAVEj7+ICmmB+gIR01BaFa
hTzTI29kbPpse59Vw+wMvkTNQYuaOv9rL79kaBT7GIrNUDYreBQFgbozk24oJ0mTIxhGvjnNB9A+
n1ez5YXNH1rEYOX3bpiaJpzoKRk328xKA4uM9vyUSftuDGKlSThxPT8W5WMu1eLN2CbBLo3vEK5H
1GFiEiNqyuzIJiJKTbNPB+j4pCTr9mucOS8AgefxPDPDQNXNaLTBBISgn3KzxlNYJ2woEAt1reca
Z+5NXzQQ1HWv8kcJfPiCz+OgncUsXNFBsXw5/hy7VNqSlm/xPCoaBLw2aYKKczHQBqCmo29gMmZT
FfKiHq0Od+FTprIPaOtR4jaianpV1A+Ygd7e9myjTiv50HZiGiJ9ik9VhZro3IUH3f31e9PWt9r1
gi6ECG95Kvr31hQ6zpxp+x8tz7FiMm9EEk/AOvOnOaHIkf0zoOLolnkZxUFCMUIaSBCYtBmduNRR
llS/7y7SIgwKg4+9Nbt0ABJ7v8oPUL2aXMhrXfKWq9iCMmaKcEF4dlxp3kmGYJW2MigS5gpL8DLs
uguDn28Vo43lNzx39aW94MCuBa8h1YZCNPivQxI/TryyKyJi+p4LRJjfZzAt267dWIRB0FXkmiKp
eewxx/fRdoYG6ciLP5HVHeS74htyaysS4vYJ6j4uaTQdMYm1w1ElE1CZsC/D/XYFE6y1ViNu4uCM
U3RtlZZhru/QQWR1+9t8eBM7XoouaRKe0je0JYH1vQ7WqTGMh59PKCTw8+TH3x/eddM7HChfZzMz
C9TZeJARipG+XN/xSGA/8AyeVBiY+RmG9gCBTXskRLMNhWfNbj1GnD5Xyp3Wx8+NPRrbvZrmRoXu
ubBzZEEZ5YWmgkY3S7DGv612ww0FLudsUC46cfKFNg7sGxi8VUOBT/TvV1ZQbSYWcU6L8kj6HxBa
tyxWgiDpJjtEHBIuj+cgv32Mpy7ULc2ZnEj0/P5YiEJv8lql2cvtYqD41lnW657nWMzAFxB5B0Ma
0NRDHG9eY18JWuzeJSqn6+z6Li3lofsOYAOaf7GHJXSi4a9HxrV+gvIVpBw4mJ6Y49m5siTAIhSh
uNqXdR3f1rtEl1KzhHFzGvXbaFdZG97zt6qaG9JmkdPef9bejqf1XVMfhXbDBoGU/vnlcMqcZPsz
9GxvgETH4O+p0MaVFXEyKUy2Q+wh4v89LidQMIpy5b8TDGsUa88QVpeKAiwBCW8nTyTx7WXEiw4h
X4xH7an3sHJoyppqB5QrP5UXFMXv5wgu4RkRsx5/kngkRETuC3XB7SbCYEWNNjcAFhO8aLMOXtNb
WnCg97G8406E77sdcnfNHGYmXdEvkfr7+zWH3upL7uV5ZdksFmPJk3Bg2QNnQTuQvE72XNioxc6A
Zo8zs0f+MK49rSlqp+F2PCOjkYZdo47heJ1kSvi840bmLyH0j3CMFLuQWPCwjSsVRhTvNnz/xJtb
eLYCqQwCxryu2zrNoPIz/p1cQU2Sn3A0dLhf+l2+Ad9izSlk/27IomcVfAYw4osuc2+RAt0gajS/
L0dvht+Du5546bwthAtClm4uA/XKgRXbcgpCeXv1yvCC13mcIjobsiq6teGUJPUo/QqtdJN1x4+0
ZyJE47wLYTyR8BpXaNfqHi6XLGHtx0D/6cNb/9ZOw0uKsf54cmkVTGqk4fM7NjgShodMabkMFudG
j59XXoVM5vqmSBGl86eKl9RvLrCC2NYBHhJ/mpxpyPdRC4F9KfMmCRK5KzNF/jaR0y0KQK7tpIk4
3vhTWy18We/jA0HQH/Sr7ESL/zXBexrIzCkO5xflwjprz0MAlimAltZzCBlHULQh+E0hy9g3W1nX
A4JaksSHh3LUGqVWu/xVg0xponYXu8IUWmhjx3+yNEfR+ndSZzCPyvkoB/z6D4YmZlZLF/3GMFuU
9nu/D/MJRgWHMN5XLUvymU4r+F0XDkLHM3trY8mRdC3Qz2HV1T8STxrDYlDAEVnsLlVstS4INa2s
E2Fi2p7pxW/bKHYBzdpNj1A6NlSxja/h1fMNNsb2G72gGHp9Hkd/npHLvEotUyEz9c9HUe4hFYOw
deLQObrkjT2M0Nd/kQbYyHrwOTEwWRwx8MIPVvE3oVwYUq3xFoaEbgTO2CnXvpZ4MkrbeWfPzTYx
bzePvNprHGOFA5Vt7pk5Tpue5qvxm/zR1lIXYQOjaors1NyxGL6aP4KbC25bKmdlfAgYZFRuHsL4
5CRqgIF1g11NiZ+5sQD2FgkzTioVNwYZo25jI+SEhjtSOmnHNJHM3MuAuFz2Pfytsy7K3hcV92ri
1xLlGdQnnF8M1WJAR8Ni35c+H00OQHeb4PRTXjYh8T+vnb/uDwx/kEKS6u/V/CSFqQWizs+/xfgH
djnDyKt29gPisTjvgWZXvh3a+cfCuht4ZV8OkqSfDGyTVSTwSEw8LUiYkxKWD5WyG7wfIbwoINoy
ART12Z0F1kfWElb1UvdgICY1Dl3Ja8cjTu27AuMydE4uLHuUJdNLqtkKrQNpyjFQdMvbGICZP+x4
tQXlaXzPEQ2sd5L80vTc72dVrNXKq0HKrIkOzO0zZAfrWKIkXlbqRerZGGKgzB6x/+Zqjo3P3OQV
duzdjHdiOeQ2XeW9Kfuqr0Hpbj681AE3Oo3RlTA37evc/tdPIrbgI8T3zpKE9p9KuVMNly3AKiAp
Rzq572nxtnzN9mv5PY5nwCxH7gxMKtmzMWcUdpQ9ZW37FjoOGYp/d8y6ag2v7YEdhm9y6FL1Efjz
MO2/rtG3THOfYOLklkMVmAk9STuo4ATWL3AbCH561j64elMZon3u6i6FzHb91pw7p9vbphgENRP3
jI5G67sTMWaVOTJKqtJB2qS3eSbqBD5YyeNYgb5jbZL27fAiC0dP5s4qM8HLFy9NIlMgty8FoTHb
g5bnVUYoiGR9cJlYLKh4nzX/zoQRx3QDvNb5z1loQR9R+xNofcVgVXl1O2ghp0/WbEuHm6gfbczM
vjF4rpYJeb/O65LX7Q+Q1wF9ix3nuDpSe3uPiZubzvIIULwCdHSPsxSYlWiMVDG3n2np6jD5pngT
zx/rejsmu9qYIa0R6XxSOifsEV+0eqar5o+eVcmw8Ec2a4Z5JY44wE2r+qiMcks5cMA7qbMPvekg
53KSKrl2fEPpH5MRf32qhbyaDA8N6MMmRwf1uTVHtSgIXcMaJTirIznqd7pQnrOvS32nABpV05tY
TX6gp5f8dinxaRf+Woky/Ejl/HqNEwt3Q+c+4KQDh+YXo/KQstYNPJPur7BI3wVjQ4l4uWamMZQu
akxnJRxbLT91k7vy6GBlEk4ZObQv+YUEDCDF+xwER9t20d4LqPK0VwqMPQDBRYJsZIZtuiUORjen
oI/jqm4qC9JUPTuU3rGpEGeI1vE77hF8LEkypVc89p7N0xyQQCcHC/e5QK3EA1SPjsILBuSQaCEu
08tkqZOaZK6YM+3zAai0nvjx5Urh2rBCrqrSjrjEuR3e2Yr0SvBi7J//lsl8iVy7y9jlcvX/arlt
s7kJAiyWi9aZ52nUuZ3wkKqwX2TNwBqbrON6po2FiMFRvSl7TdAp1MZHDpKnL0FBOwiJ034Ux5KF
alu9FbbVb/pnyqDMjRyKWCT/O3W13iaCO+/WaJwHLcWntx+tClSp++CiEAnaLy7LG3L7A4ux2eJp
f2aexh9vxoNjBL7zoUyfdNB4Tkg0DiRxF1pb8/8HHZOdzaq56gR/yxcLkHC00urQwe1KmeMx7gx/
4PR7My+TGiFPYNWN4O191hKer+Xwjv1/rpjDaPSA8qeVcYdLPie9VR2KH1TN7OFPSqPiUO9S7P8r
BkngUvrQSQ+Sy5yQEua5YF34g+yB8fWlUpCV9pxtLDMvxY61z/dkX33FFOSEmvVXgrn+s1nitDCr
vrNgH76YCIRYFr1CBJJBF2uLxGKuPPzkMCnjXyyyw90VrBKxJMRt2jOjsIe8WIGu4tLyMZO7x3FQ
wAMuw1YAK3Ztzz4u5Ci2f5EzVtuGPjwoXwYLhOSbNjSn1dr6VcGfpzcXgZtNpq4d3AqIl30aMWYB
O8TRBJI+Qdi/favinU4rJMTvO3PumY8x0tMFl+kAHxRdF5uF2vJvW7UX+uKYgmDpHIFHV6/VS1e+
JTWk//t0u5xv2t0A2nVgmxGhU4TYMB8D3eDYzUwMWo+bUxdJKXVYkCmi6F8SjaCKWkHx9hc/zqGG
kP4O/yeCEBBovBw1CVdKFJgClqM3QDZstl6voRWv70IBoU7PkEV4QZwcV9zRe/6bj3bkRr1sxh3H
18A3RuGi1WyZ/wsHVaBUjOHvrxs9vrfpf8N2AZHAC8fKaVkKJqqjHqC0dbtKxhdiAbY0szD1NuId
McTvV5nVdq6BmSkc27bw2ns31sTCbEAPet9c6K+lRPXHbSyjE8zaH2Jf4ecXk51KXY7YfW0zZofl
qPdOarGvGtvhzWcutBsb2WoDSXBL0IoNfS+mvxg77u4j8dvyLW4c3BZGEqN+O89Tog2tYKlIiQKz
BvE8tm0LCrA3jzHOLNILVhLbcpYMl5ZgjEJlkYgcbgwGMVP9zYO6JsKDZZNAzXBnK62EgkEkz/p7
wRab31yT4WEIFjAi1U6nPVB/Ye1gqPVg0LdMy8M1RxLRFWfQ/6B99Haoa1aDK6gV1Z8rZdOBIf6Q
aInU6JG4HyA0jL02cZ6Z1JJ4mT/PAgRdqiHWPNPc50G1+F3BeHWr9MTlbIgassJnRX5oN5sM4PSJ
B2qw5MNtozajSQD9nqVpde7TcIbLxHVr/tolpdBVQKHid1MCqyMREvX0DX0FYO0heWOO7MjT15fJ
1mtCXPFgigmRFAATMWDJxMGdlpUbtaLG1zk9UVNrrFx0I1/vBXAf9Fc3fT5nO/1DpJHehKxTvLIv
CU0hXiLBbwa9LRzlkc91NJXMFs1NzvQVfPVEz7Jqhtlima8Gz7AT75+rCfvNtVj/+WfZi8sCdF+L
/pwuztqgyYU6+X6m40dnpltOCMvuEU0dQHEHgKAp7SEyrtWj2BK3hRZZmwRqU8so245WNvtCixU7
AuRah2kXqOzd1tXQX8UQL3z5x3x9wy0ci49MFjvwXXmhmx4ox4wRzy0LgCnIRLOKZCnsh1YzVBt0
asS1QPn0H0ckgnb9GuGJBZeETyM2D5oSACwnIIi0XPA9b2NzWdC0RD941f8S1G+3OB1GL3+CyUuK
K7v+8xPB++Ms+0RQG1sCdudCaGCvoUMafjp2ziNBK8TjertzQZnPIN+QlMX7DNijBrmN5ZbKKQHQ
3AP/WDZznk6W3gGVXtA4Gg8BWG0rzpxDNZgo+1MeiNWJMbJIsCxGycxK01n6MmFtKY/STLZOpxqd
DKX+Z9h63mziSZ+UzqJ9vd4GnIv6SZ7tzfpQ60yZLvdW47Yj2g+YewaVTY9NC77oSLonvTpn0q4O
nkjfuie1tfLGp3G3lJdwb8IK7jPP43V4cjM4ljXqVebS2qkEfa17LN8U+naswsuB7ddpNA7uo6h2
uMTNpHf2Qyr3hs6nk4y+4FEQ5tTGLf+fZHxBCcCUVOHcBVAwG3gJd0a8P2hsLpEta1n6LF/WlWrw
JYep+5iFhn4kLeKvwBFBnpCjM3N8C0irLSdHYzlF3U64oBirlw41IQEx4q0k58q41zXuG4IhXdw2
YSTI+LpaLB6lSEibR55uIVhCoQT8DRYhEo2RAm08RF8S3nE+KE4KaOgVKf/BZA8bMPljuwtuIV/4
rKPYY5LCuYJ9+HlW/CeWNCUtg/Knome4FnDX7G6S7KxACbebEeUgX9pF0BHrf1PD7934QZjAAL0o
pORIv+aG/mQo7nfmVIpO7FGIXQZ610oe4HqHy6kopzyMJNtd7FbiBKCzJkDWH77WWr6zzPSA0GVb
1h78qYqG1F1QP6aDVRFVz3dzOK499DPMZaE3yXG24cU1e/fg12P6hDdeLjJJuCUNwhxTKER/0J/+
2Pb8RhGj6DNkfXHviBTlsRFxmbMSbitpat7KRndY8tGfZZ96n2XlpumNyHdnfLTUN6PDvFlZ3trT
dXp0PQVT/r05Lo+XhCM3VlJiCNhXUnZiB4jUOxdb8DMpEsrPrGW9FzZ4/3KDaX7f0yLh60eEucoh
BuzNIuJsy3TXem3DOVFZnC5oTxnk7NQHPQyoxFl1fa5tyRB2f6ezIAsuToyryLA0+QzH1qzirl/i
PWYkHKV/j8XrIocwjDu/qrZneYilcPcn1E584HEyBdmQXNQUavAlGUhmVzpYodiFsq/tz3sTDmdU
1JU17j3LwfrJvGhpEM5z4Pq78nqwdzzHrhs8p4btCbH5oBNskuPQk1cHe23U7hmdikdk1WfaWfgq
kAzdsoTI+OjfpNzJ1OB39Bdp8Xcva71dAyvOllfHDgLZhQ2wGJ4+Q5szl/jWIUaHOZMOB871ZJ3F
RFBVyiNevdgskMaXKJXQo9uzdw5If9TkqtQvX05O+S0uxIz4llMYXlRl7Oon6/4ed5f3zSDzHNRk
i19fcW+joWDZqwsGQwxqpz7d/6g+JK8/9UKmQssTCesjZWDk9XnZopof0jeQkAixhJ9K9C+z3w7P
7I5Y4WU36mULg9zlhbZvDCRUP8v8CJqvvTYEV4H18UHi99AWwlnaGfAKJnNwuzI+9BKCUHKBRVBa
7s+vtYF+uFtno11qr6zcyvgUxEBqifoRQgO9YEyk/GxfvkeEEOiQLlVIopPdueLRdvkx2v6OPxTB
X89zRyvngXuXKoAfyTiMMROvms86iXfISFi4JaYBGrguZ8Q3ULNYDPvidsfttwkpe4gnjtWqFu7+
PsNxN0HYkMg25I4mhJuPkbkuDl2lD7jEMXH+qClLGMPR+c2yG21p4oNwkj6v49urIGGOwEmyuvKy
L4NDdY2sRXBN51Nf46aHATkV0GUcARx575+9u6/nOtzDcS4T9QPq43W23g1ccfDWw2hPGtnRbOGb
fcTy38a3U3ZtLjl29t9SXFcrCswD5gpF/cIFTkNoa4d8asZJOcNU32wGcFDf4owUR6DU6da9tANL
D8M6ne2cBx4l8aCJAv4lghOvY3k0OyxhXNvVlz6S9l0TQ15cpDcOt5DWMDDhe5Wuan+vM154Mx1Q
GOTm1VRa2BsdK0UNixQp79qFFc7Xd03y2rglf+FzS5s1FgVrDUEPYybq0V9HM+iaMYE0qF+vNYEn
QB0BeFDu9Vy97F5R/VaTEJQVeEtM2U12LIq7H3ks7V6HVCQf/pJZTyfJOcs8P5nrdUJBfQoPNpeM
LcFgre1UA+qHgVeJtDiwdbiWqIzCztQ+Ll9kJ2bZw8SU8saJmhv2ov0ED1lTCrR/8YDUrEC6jth2
5XeQ3uDhUh9wpm+ZpAbIkJlrWKaev9KYY7BVGztXnK4/tNZvOivm8kKIZ2vurThvcI4Vj66MwC8i
gvm1XzqA/L3aDZiz/hjdjNbecJatrM1gDJQ3Gud+7TP9afYG8FwKxbF71n2N6Toh+sQWHq6QEvZD
kVVZ0hWpFnjRc7z1Hs+a+Bhk3jvXknuzKjgUCILj0ES6WPSwQGPncMylOEB8o3vTaJrNrNKa3us4
nbYZb5u0DqX4eLZp0/NEMN6AqpNX0bcAtWOvkvJVvS2DUtKpvhtOhdUQHGIxx+p/Nw96ObAoEy2e
/HkG9+m50tvEvWjLkHYO3uielr1P2S70IiM2gL/o60WhtNgBnERlPtATa16jJElv1Rb6W0/yg4uJ
u5jux7nT8yMYvQJhEnQthf1Revg6AuqQUhKm7AeyrkzJSHIZBDXUGAM1QWLKiRbJwAixaqBg8x0r
1OsmHqsJgTXk1HUwBVgiYOslyCQ38D98GQnDm4aeDjCtT1LAuGi4X38RDxKLh4Yj/kwAIJ1FpbMG
yMGNor1aLLPZbJMY3ErfGbYoMtRe7QP3zfnNvVOjwVL2hTmgLdj8/Res9bHysbbyZC2rPxdi523q
TmV+V38gaFYLJ4HVlzzkPKGZkn+gyI+oWMKqGIpHX//bYfrTIn4J7RmMDydH7S8tWR5c4vI3Ljxf
3i/4Pfii24ij2qZ8E4tI50j0YvE527/SDGb/EshSo6da+8PHUUr4FO436NusdHEm6qbRyGnTsPNf
AAK1xf3Al7NbB5Lzn8XfB1KzsCKlJWY6JtVihFrCcSmSEL76N3f3mmuu5vDbKp1fg2rwbXuuE1lo
D1k0aaEXwWBMYG9Qsv5lwC4hQR5yRrVOu59gA0OFnX9j03nyuN1P7VMNngFmb8WcXrv92gvTIa8K
3GqZFNl84WXeNnJY6b12xFGNVJ68geGDNxMo8HpgSWq47+mekV8b22gGF7+Uhvghq08WS1dcYuPQ
4yH+YIlHK4Isc2o0TH3NdrWwds5TXXPLn0+KiiASnbzYbNXLaKUhoc9M0MAWvTB4R6nEwABzFi6I
fGlZ7XI0S+3ADnxo5qXY3X6HZF4opx6N9VC66F5iKnXK02CjEobLc3AErX5cuNNflcsy3QVUIsoz
cm2ql3QJcd46zBoB/bMMI5U3rAmcNO5weXd5YA7ocnCXf+flfbK5/VhTY6mF9vyH9rhIS6oqIcDa
K8A05Z9/6lluFPBZGHlQeicezJ/LpAUSKTGSGA+l7ZZcoY3epv+aeS94pzPGuKdzy4lkd4yMvj3E
kqsrKpHBbzO4BpA67VLy+nHUwXWBcdjSvxLyaUcztOly0RRdRMWLWExV+uSBNu/l59Mh2HvmcSv+
Pm4gpJT6OAw8ceFiuGXPMO603q8Ofenrm0ogkUhTixzkn63ht0Wz4EQW4OZf3fluXwvkMfPv/MJs
IroDivUlQMrZjU1upRyPiJ1bqM55tAq2irhODyQqwFuxrQjJN493yUoc5BIAHoRsy11wcErxiTrg
5rqDpf2bGXeXhwe6lHHa64vgMbHi7iqihWuL9ln/Ra9wsOXdnWVMAfdWRyzhLm/m+s7/yndqpOH8
Zw3h/7KX8SWlLhJpJsIoyUch6yj2B4FdpB82WTQeYGyA9s0Q6/3AAyLkMWe+Rtv/UiUJy/WiaePV
HuBBetG/RSDFPEXf+PONF5hPbPs1YN7kQZgKI9MnJIhz3TvEereLQeThuP0ENFGxHO64Qmz8vBDc
3z2m62Nn9fJ3yiJOtIrawllFH6701bhb/EwFb2PIybiUmbuZGYakCBfKy519YRtb37jAKPV8rEgq
4AL65U9Sf/nhXkYcYxljQHvzALVe2xoftfshvcvtPzMy/Oor/9SMJJmXjeXgiBZz/1A4adbyURvR
E7wGl+BsBwfXLgmAmoeZD3cE46xfu3GXVUqsWbWlMnaBadmtgEUKsxypXrllWildu3+7VDR1/PGo
V45ULCIz69CZgTxQmrHbXKQJ0q1ugAjU1Qfvl0D8hjQJhf3TTmPEVjkyyhxuU5foJpFDT91LFtds
ZG2EhKjpwWvWL/gReoNOBT5rwGQyFQCLIMGZTMi76VxFk/piUMrVaKY+VBTXQcAy0F3fqfV2QEOd
yhNyBc/cU/CWMBBqcPYrT4Mjr62rcWegD02EI+wtJM0K3yoX5/QYq2bPnT08b3AGe8CSQOIMA5tT
tu5QaRX5vvd8mWcZhN886WlkTzIQRIG+bKYO9BB2rp+p/4KPTJxUUgCIrBRdIAHqmOCW4zpTFQ4q
WbNHkCaXJWFZKaN/pFFabivLDATB8jE7myWvvhUJv+hzQuV6OitnGl0gyF0Hc+SPD+9S3CgpnLIy
1LnB1yZVIAvaIyFfGukLuU3BGqwJJ9CMASqoAJkRjjmeKTmLLp9NtGrplXJF8gLs2gj+vv/KD19B
F3eEe307EmZ3CZaWkkKfKIoTGVt/jcA0TdiBTJcpv88hPOdeQCihi0F5VTU2y4wPJlRLQUe5fjHe
TNJHsBWjiOgP1vFoUJpkuVWfm9yr5cJJ1ss5EF0HEHzVOpfPEKVvZ4b+6+Pp1rLQhPZUHySEoz29
GYEFEYrlNLCXjr4EpYbYIYY4cbjQw7WhFj2BE9JfZTSEdsyV7rio1uaXlo+OaN4lV6+IzV6ayd1i
yMHBH6WnIaZYLzfqltKQQFTkcpfOUwQ7AGLKDQoquEQZWwduKNlFJ+Eo7RNG+UDs5oufHJNGu8j7
F9gCw0zeuXRnbqkS+EuBgKt8JUHXWtBjZa0DAwoDuCETu/GzQJsJHMawffXCB3wOn38ESw6Su+r7
LcZ2rBRwy0K8hP0+fLSBgmFIlsmDpSAR3MlAZjiC+OtN3waIynidJw2l/3sEBPFUCVqi/ysqVoDV
TGPqaj2lr6MUfigJlT6GSs0UZssbEy1HUstlvBLPwLW8LCKaD7V+/D+qBXZ5LT211eXeW0OYdPex
LjzErAZ2l4RH3eKRdL1RFoKu8R3VJMRoFIWqtkjANW/a2o+QKIiHSBU0MyU7S8drnrlTXcf82BFO
PtTJchd59flVMc5423Hjkfhg21hUqpmo2QLLUyoEz9xDHuz+PeJ//y9IPLoVQOrZeVBLNI+n2uqE
YB9VRyVyvvRHe48PSgNeUEFRaQUCm8CN6PsnsWkRfJQfuoxx3q0d7KvhAYf9qkw/zcLOIqQqCW/O
7+RhetN4vf4w9t8CtFV974LOT5lQRZrNrZeROuqs/pTgC0FTyqptz+mGyN5nDHABnfBVJcPu0Oh7
0p3s/iDyzKExaM8r5OFY3EXJr9Z32tY6LRDy298tNM7dsBdpYwmfmpP0JOhalgorymVYHiRHUQfx
uw9i0M8fOhJCV0A9zSqbngcdTk31lykyj1cZ35ggLZiwKioEiW+ZBRlV4JAExE56ghy2FrtvLid1
iyZ1ilBOjLPqnvCbBry3WVks1ldfCmre/yyvnY6gPBHBemZcmgq8kJJmE3u38fH0USnLZM00HCvN
AwqKk+zkjk6KGojbR4FZfRkaIJVk34w/aYaqXZpp27syI5vA2jx60BSf7fP5V4mfrnUsKPIcRGaM
g/bM477Ru0UusPOVGezPR1W2GiR7PMEUT5UQbxInRcOEpjceIGCak3fuKvUYrzTnzF5Cs/t1GGnI
WIC/dBhvjsQgWXJZw8YwaicyeQFC5pDgemGKDsfQWz5AepwSrDw8QEZpeSj351hld+n+PDBxDXY+
gMzbI0BLGUvRSuk2aESCJXDZAX1VOr/ZDLM1zb1hkAcmrWhB67o/FCSb5VyfDL7RReKnxejrZJTk
ELxraA4r2r/p9Q358qZOazsLA//m84Co+WSfXpibFFYvJeijTly+zfrmCFSF7C0eSGE6tBnUQuJJ
BZAfFvb7cg28aYNQ5YBlaZ7PdiqII6wLC2C0v0iorx88+BmawOc+y0Eedxoh/zNvuo2ZeovV9x4z
zPW1NKzbt0cx5d68vctHyAX/RYJGGoWbnPsV2VhFU3aFbiF5Z3uPxPq7Yp+GYDKdwYMtLMWs7zbv
UAet+ggH01AFBljvxF4DDKOjrjWNSRM/YFMYpDMr+qJg0aoGV8RDkJJ2VXucv+bcIHyC4D3S/XSQ
ycWG6uC1Bfq9JOWQD/9aWcCiSPXEZWMiiJ3mmsqUlc8dpmjH7Wb+3Ti8PAKm8+4tNAqd7m+OKbUE
orXfeR6CrnxO7DUR9ZGFBtkmdZRgGjpQwc2/9fl2/WwZevp3zBfibsuyA8QCWTdx8NgKzPVdXjiE
NyTVqBbgTypoKIAHwyHq0JnwvwsF/hphqRZcCxNUW70L9g3QiRLf5EYwjHrLjSJCa20jWaBXF1+7
IaNG0EkU3V/dFES9vRhkjJguZHe3GkSCy4TN5ty5e9mosn5DqtD/6SFcz9aJ6LJn3AHe3Esa1HNT
L02QDZOKNHhY9opTjspNGbq8RMxEbSmFUohpM+FIyri7dBTh2dp66Rn9cOwTg7XWRsgpEzDcfA/6
QRvwBwnGb21jpvYhXWzjJzyP8/7ehjM9DZ2gO+ZxuOMftEVsRa86oSf3VyKnerGIJU8g8acmDNK6
q5RJ7CPNxtUf54zqQ65wsmEPMTyC4oxaLBTYI5FG770dEP+8hrpBZ7jY56DqLaZT5ltFDJCRjJ26
ja0x9IkvigLQ7116O6ABMaxL5IpF/zbwYWB1CKlQQPSrMR7uWDR4eKq2ShU4lDOzs3Mri0I6uFqR
ebrefjhgyShlPUmgFGAa95HjtXeEi0LXTRG5CzWrMxAs8/rFvJVqhXvk4yGqZfXMr9ASe8+mVOiZ
4vZu58MrBSXhtjwE6LREsyzqsETeI9By+mfvlh1ijbbBFQxNSL8+9B2K34bqHa5W0JnSq7lcMAp5
3y1ziuWVTw21Bqmr6oEfCgoH0vjBs9gWwkHQV90yCX2rWAV1jbXGfGPxjCZKHRL+JRsGUjazI1AL
KVSvGXNQzKVc6Q/zdYCR3NTTPodtTwlXxyttHdrIZjmk85PFaMEZbaf7ylHrKRGrG+z7zzjhEmwD
sP33veJ9jyCmEfXOQZDEfKExYBg6q8wXXOBKjImtpwfdS0le/hIKaqJjIDXFdSRok70HI9XpPuTz
a0oeg6z3q/uBK/8l6n4CwS7aStqauI/Td0tkvhbFnpQlQ1omJkKzguKEO0YEgQYxhoLv7o+qn9TV
UPZyX8Y2vs+ruI8/K2Mcyb1TFTkmKnr94ACu6xJgxvhmjhS5puSZjeFcedabqMw+6Oz7k2oAtxdZ
TX7sg0Xi+S9q+EOL01yR/IneI3ioMK7fKoyTYDtHxvLfig2lqnC3+J4GZjJ5i3E/CfaHoIu4g599
cSYLg1uvS3Odo3VQW9eBseCweSa3TekARSySzcumaliFDIM9/mZtE2M7DpwlgmrEC7m5DsX0/PkF
8QtC9VhAbzJio8bL941VjKXuScpqy9arVHPGMQiDyjLegHOBdNvqmRCMhnNU4RSTuckiCFy57U5y
rVOrTZ+btTRS6zur34DILhKPTYvecfBMKTEjQ3BIzw4oI5mJ96fWRwPbdOUjR1R9cXfiQQEnywNg
shEriWAYDN7ssRG6sn+pWK3gtTxjavK0MGGdHAqG+DgmiXzEjGQuinA+ndCX0MN7mAMf8biVVufa
OBD2AY2WDPo9bhO4aokkMXMXlATpFSikPd/efaUJBNHo7fsAabDEJwpqMSJN/v4kDwqIazU1g3WC
aAudw4VH3GBm2yq2XWD9uMn6atXsiet0OTT72oFq0p+lma5fxxqvnICs9o1dsMS+yIz1Bg7LhsB+
d+KzaW2xwQ5zyaAYxpxxRe8b9ghjXqwlMKE7fAB7ER4VDh4e85+QAJhQpPjP13ZuTOCMx3G0qLox
0ZmeKyi0huj5LlKrnw6L1QhkdeO4/jGljtu4F0vPTMlHKOF9HMUlCubCCHsUVIKZEae5thiSJgAx
8a23Obxyy6GPlHwC6XPDCzAdBwoesVFczG4N6zO/Wyc15JlwEh60jKti1lr7f+Op7rtE1mPtJZf+
pDToLxz6yrvMv1wuJjNmqgO1hSyZLwMKl11c05ncXKI6kUmwK13dHGVVAlq5gOqavlVb8Ujlc3Oz
Jkoo1Z9G2Mg9UT+jlLPqXa+cxzGDL+MLdhwcY767onkXg7UCuOA8yIfici8iTiOnz15GKsCvt08h
GrE8v7GvEA2n0Neink/pN6XT/G6Ad6rqr5Gi7LMKIVMLqbhFC4WuP6LQuY4nvv+o1LUh4fRIQKWn
V/stXQchA567sA1F4G+Vfvhy4RvuGg3SmAwdHxaGMisHpQ5004YEpTp9mcSWk6CBMTEQ1o4hVfGG
nlDEgzzDa08YSlZyJwjQ2U0Xz+7u5Cv8qQ6NO0Ev4KTp+ICL3JJyqVG57dikEhmVIakdWObaMlBf
p+JiMpCVDNJAtAVBSUZFR8/buVUebgGUSmm/jTxBlraIclzVM5HZFGgumz1GIzxpBSjOTbxqmkhA
dG4ArcbKpBa/fIVUr1qZJFLtOGQEXez060aef3mGRzq1Z0lK+FRZPKbiapaMlmdQIRS6fCmCqaJq
HDXtSDEccsPTxIOg1Cos9jGokoBmcmfLYPzRvoO992Ky/48b2dz9K+t4/GVHg4hUBvHQ4DhjeLXd
LrBI8DgdN0YJ2lE848DcF4JoWoQaznEFKZhY89RDP212JtlETdV4imsJZMq6UeF5ZoSwSSXHh+JE
Ee+hK5qGYczJQ2YOoW1Kypj4bMVDm2FnOMrYETmTX3PBmac9bmIzGLXXlr6DLwZ+EtIORUSBDnpZ
ctNN/aA0oXR6AubAo8pIgMPlulYyD+KYZtxF2Al698zGs2Wjv9yypeP69BVXE88RTt5eD431ClDE
WouQD3BUuJWSQ4Xm/H0iajdxvEjEWNBalNW8Z193olQxb6zAPAJatOTKzf9xK/vlKVZeKRKJiLdx
5qWk7dHGhTBDJT29Tkt3xBaCzAnpd4WAd7eAZE0yEnSvW1FSskIR4j3MOgxHaGY7f0hwSMgMHCft
ompFATKkJdkinEa7hJ8sWRLTdoDkkdZAyJCttKGGXKCtkJcYHuQM28kpTVxHDkqALZh3Tawrznxr
6UTKGSo+gQMlrj+NCr5wQn5mqKMOheddjF2paIhwoByTqIWn8x1zdsA0WnJQ3BdGSOLWGTMtTuSw
X+646ur5HRoULk6DGECEhCd2JMG7UBYA1Q/nMPz4wCqgH3Uqf4qzQfevV/2hZtam2vRUqZ7gcJ1t
jgo4sQpuul/cUgmBlm6bFz/glryYPuIFyiTC40BOl/fSXJMR7Nw7IhkWcylejRob91yjJqtYyQmA
MJM7ht5ghrgKl2qp6O+E1Or8ydd5oVCJyZ4V3UT6fpwwNxgC1xDYHEYsXt5JEgGBr1gQrWdm9dcQ
NYXdP77h+Ob8341x9p4jBB25mXq9F0i7jIEVUnEK/o63RGUqFZEvLjf0Ej55ooOKhaZJIgkZyFub
f0LTiLGOqqobOjnfrtOCMir6W9HkgUlQi90EbRM8UNIVUjODVfsTt8hsEnj9mck1xz8k5/HexL9+
BOj0EBeIpC1rwHJQJZnNta2i2whg9Gou3dvXGZBdsQQoYi6vVsgbuheJceFPJEDTFB5FtUh4f8PM
q5IraOGJzg+fDwxIdbK1Innv2ZUk07jbDkL9jDHTF+rxqvB9+ktb9lPtuRNXg8LMyBZjxV6nT0EZ
OP9yACOysRlQOgbNHALRDXmbwwdPpwVP4rfUaAmOI2tnDHzqemiYxowTxUQW47OoSEj29vjdk9wz
kvhMqCwcQWtUcDAMI8qKoXcPWo5+8KL1Um9KJQrcMgrQbOLtrZpEl5Dvef2te0LjB9AXQ2OGw9Uz
CD4RKKNiU4waGoX+YPYhvRoSsqTigT7ClnCp0drUCcwhPYxKFGt0m8iQtJWqeu2+KrEmHxBtVJ+M
hjnETDS3TCZVaxJqX5SIgtbSHxYU1DE6BRTERvMSosvkg0aLlXtsznNEqcMu7Iyltbu6SE458mRb
vjJxZhoacUgI/uflwxYcw0UsCHaejOyJ9UPb1DOkrbpjMRLc8sJyjsMmupwtOwwUWixHlH6QLXWp
hyRNyIsGnZNyOv3BmUyQn4KUgfFmAIICuASpcZkBRvrQtYs1Ph/aVNVKe4F0uyp2pdujkYwuaFiP
b88vuXbeIRCe7S2+M1iO06Sg5+HWJ+FJA672ogt/3HQsedJEk36uZHWsRq8RpSiLv5Feiwy7tTe1
sdu9+Yl7PyGj1PEVjtjjspavJpz+eU9St48lzZuDWEyWsBihYwj/jvuKGWZraJoqEtCLDrWhIFMR
easricbcOTMmV+7QlJsVTJQotEm1t7SHRZ6BOg0rrmRb09E/7dGH/iiprQtQmYtlHsBxuk01PTRy
fQPQgN8gtW7rOjdd9ZPcNCXeMpcZcGkEegNr288ue0iUqStKX983m5msqwI7mRavmR8QLy+oUmNG
97D4x7NOAMsF2ueeJFsHLvzZcBtuNiMYGgOJWT/brzpHMof82KYJb7tHGWxKY3lN43rLNTFLIN25
BX89LWFHOqttRZ6T7AhFCIWtKPpb8XGstXH53BZL0WOTJiW0nzcUzcqLCqyontENeyHHCTYWUyt/
yqqRz1NhoDTSKIPhXed41PTTOrmbGMa7SsEPIJCO0vhuSTslTYV+l6XB51NQeXOJMYJsbDibYmJk
/XSxXXYQiaaayr9kOWzv3XpVQY6n8Usg6lBOm0Q+mASFrM1DPkXrHODi7uB8DR0YOnrp81y5BqUH
HlG3AK80smn5xyTwTtglCyt6g7WAjHOOiZAN8LE+kmaYAzUrtwR7LYOG2vUXnH6H/jtX1GiTe+zZ
nR6qH24HPphzkab6Tpe74tYDT44wvJnqrQNkr2DbNJfkpzPZNlfGo7yuK6PqfiGDIsaO5ZXoJNNa
R9xPqzr8eG6oiWNuTNJPpJnvBDn9mpNt+1jLnL6o8narH3I5ZkcEQGJce1aP8gkRgKF7EIUMaH53
sGNVma7LGAStcF+yoPAK3QorkfjdwHN4eTTH21gAMSoW83lCfjM0TkJaLAUNr1RnmCxYEAmUmuzL
U1tDCqIU3qDASkJ9d9vgL7gBkdC1U7RB5yJ82RXnBxQTUiFfsu/5h/n+x4wUNola/Sx5+o20lhqp
a3btRHom2LKhR5ic5GxW1WMXeUF5Sg/ATgx1iRecmuu64u+ExqYpXZWlc9ziWrdHCTNEb0jvth1k
ju8DXTxl8c6dHvVu9FzpFyAndlbiICmpBBHIHdy2cYtsoeGlssGkCEnAvw2YtoI+oBf0SaDXRWvB
d2b9hufDT18kLhbUOyFjEYY343mrBka41DM4ZPEwGW19saEYQM0i4ZbItrJsWtrMxVv3zX09NDNb
FUac5dFYxA3TtfzWsRAjsMWDvfGu4VPFKD+E3wvxwb5owAwB+nB8hd0ADLO1SAdPCTRkB6oRTR25
rMZ6qRI2ZYymfDAcKEmY+ZGk6LQWer/MiOyLDYxZgULuppcS13phNy+GgZIgR0pNQNttbaQl6xFP
wv15kZkq7vW5HDa+DknIT1QhztN7FFAf6ojNEqygzlNJGsjZrZcsQk2HOhOL6v+CDbbBE4mIVyZ5
nqB+j9oMDGgm8nKKQPIJ+OEVtleT5vt5cY4Bc+wPY4jCykYBISv/HxPQgFzvOuHCN+hz/XN+JR32
uBFjajwwxpCX4OaDm6MgQKQQFNF+GWczBZuUx6hcUtNk4iSIchr3l9MddMb1WRVyjoRlqdWC/8Bc
9okrAWQUd0MZOAi8NGxv7YhB1Bt7N730ugm2aPZQqeXoXVJyLx9/XPzNUYSQHJ3Jv3Jf/2kugtdS
B2EW94PiYTUeaG4vHFmnfsWfzsnp592lEhAOK/Hqn+oKuQgcgwS4WtuERkfn1He5a8p3pRPxuCPM
6bh+rTpj4P0Qf9+VReXj0d+KzB7Kp0Yr3prROpIj1wEX6tRrQ3JwBaESWuFam/040ITQ0PsoJs7j
9U6iwfHfDbpx0wwSYfY3LnNPQE/PSrLZJMsavHwk/kDi9rmf0/vMAavXwLr3t5tdvK1bElUqzYC8
DKvH9iFsr/dtqAQD6KPRyUFhmvUko23Q/Q8zQqPRFI0qsnoCBGtoZ74AACGJFPtfaKwTohiCQx/A
yw4/omP+T/8rsZ6RiKZU/2fF2InnyrpbgS07srZmOCaEj9Cp3AdE7dxiOEEGp4cTgtga1n4hJIuG
6k4GuD1CPlXI36KnJXFJVfZzYjsGufY013YA2a+soiLArIFGpNjGtCVIHWeQQ7Hq/y8h4WlphFVm
4h/0L8DFSJN/SgxWTvxKHYRFSlxF+yekSsWC1SwXMCNY2IR7fXOib2OTI0EEqEYEfqpHrrY3atD3
e9zdzb5DYgi2G1uNJEnYTqce3BP6TzmwXa5lyQhzP0ICXZZRpObOgm48eQiCedd0c5vzR8ELE72L
Q0P48JepKHO6wYkDiA+cTEn5Lry/+S9XbGIFjrS/fK9XQ0hhIMS3VlQlzt+Sq4OAjLwq+I+dWJba
h02ibd8b+hyi5lmp0TQlWdOn18ESdRuWtzVInIOqN5yrZTe7FBo/Jid3H32FPoAwQf+cqhv8MhJW
inep4dnux+6+h8owu3Fzp524iLboDJCnppYOO/QpxBA07Ij5OYarYDTGuqYcuTTQD2jQI/BjeENr
586B94uEapWYDxJOTheatssIHBaTcjcHojibV3mLGI+uG5eP5du5eOcJIA+T5fMXVtRO/Itfio0F
MRKV74jgNxrxbub1fBK29BjDurAJt/xK8EpAYfbp7AI2sPZKERTJ1MVRMdFi/30B2sQRg0LT5PWM
vRYrw3o+q73y8cfoWendai6To0ralWGOZOHOf8wUnDBBFBgUKqts7moNWkhF//vSkFoPuNL6d26P
Z2eVjArbeWOitKvIk/4lLvZLSlhvm/i4jYc8InXfouteIsCEDHk0PykNUmBAr6e0hvVaAHZ95MoW
HVTPSua581bkifMFeSI10/STQpxKzt3U6ZjMCaeaLCx00qOyqi7DZqwxNTaTYnXUejwKkZO1XR4I
cPPgvtvYWsGkCw6NDuGe36emq7qpmqlZQRW85pLZfIBEfJSGdOewo4paU3zvDDIPafG9u5CA2idW
7Fdjn/hQagYJIVmjDfHVhCeaVsj5Gh4zM/XVLaJl8dp0I0LJKx6GFU/zs1HQFnd9KadMJ28G3MN1
VyKuPSyExyAuRigEAmBI9DamiGIbAYTbXE7CQMIkhs85fULwC7UJvNMGv8+kdna71+ROlHvsb91g
hbS8Sq4Wap3SLmxiWhxwCkt0Kp2+PtQzAruxdclej+I0USnrt5y1ShIsvGshJHseMY5DIKvMzVcj
8daPBzDsbGsBHvew9aGM5h9jhgiDj78z306WGwT6s8+LAzvVI2+MEBHse/Jg+lp2MrW+wC/nh4vp
F5s4KaRtDeO2fK6u2Lj/A0n4CUpGVBJmvXyROTKRJJFbZGYrHnf6GV3eA+YxQhUCqcoAJ18JpQHu
aSB7DMN4a26vpARi0Sa9y8MWtT5A0u4yIwDCgqMpHBEEB7++tLWOAnqdE4oMpmIC+owKILrScTSl
MTby9sjClKM2je1lwXfq0MWax59B46IGaKLZi6AA5VOFWbKjsJT9JDmhReKQ8mtbUwCz0uHpOpqK
7yGNa3vg/FLekz4V41CK3tOt0XTGm3Q8gI21cUiv6sjHbaLWNZP8uUBAxAq4dpEOcdaVntx/E1bM
HX0gD1oeO2Y7W2ry1eEqq0dhSRzVRe7QCNZ9kAZV5PpyK2rhGTRTYwr+hF0AL3zhs2U9Sk08uHYE
9KINa/UfGGllHuhjpRC8VsGCpChycsvXc4BIwWaZdM5id2ETLBi13vyJF0AI76I1I8yYEezCm/QY
mdrcFrXz5a370D+ZcNzQ07/JO2iMIAdwOdjWuXWGUHE6nz8p1A4jr4oQjvjykalqLgv1L44VYCxw
EObrqSQBs91zKDy1Vo7tkTq7mckcRmRqtJkRs3pIY/oi7vXko70L5YZ4pXX+GqfZ4SM0zZb2sfXV
GgPTIQSRrzJSh1P7UrMOmUESYpio51YljlH2UAoVsIkoe7QRZOQ9jINn6FMY6sPGEACNPHHcRmeN
eGv3DagkxjeHFC+Kkn5X2O7FBY2+UkTV0HsyneAgg+GZWLNbbbyxisUCAUYeJklU2vvpqzyxifG+
bH68hFJ9oDqktKs5tw7D67XEAMK1o2JTdUj9Wo/zVVphVyjAn0wn+T3Y/kQLX5Gjw8IO0zrdN6np
/3RlMpe361ogfAEmYXAzv4QJXNHKgQmr13/Y5OVVZZ5+AwgOKPsOm1nA43hdYxj1oRNOjYUl+wYe
SQGfIykF/l88hw3fBQT1uVI8rMheEA2tGxoeSw4thuliETd64TtsawsnCKUd7rYx84TksnTbDceT
4UgyIUAOqmXshgY8KRURbYWdj5umGTatgyAdh2INmsqoD1ikZdY4K1lizIHNZdRBzUjx2w9BfeQm
RpxsxxNcIN0GGxxHms2OwWIJDgT3BCzU8e4ypQH+1f+8qrdVf5XIAXK97NgNE5xTxXRxkTAd2b6+
TlccZXiCm1DwA0ggQSi0gKO4wuBBRJVz3js7PDBsdJBJ9czZx5tukrzUWMFCoe24yORfMjCq2m2p
8ogtv3RIZGtK3RObKTvg+RFMerV6NKytl9/r9N5eZg7qIoc3AvdViFrzU1kkpvyG12XYgkbWS8+k
n0cOhEb9u5ONDP7pi3fftsF+5EA++oA8FXBwKjNiDCjdEgGXIle5zEIVdS7xgPpw8yQIEFFvCe+S
bpbY03wt9BRf1uBhC5VKEDUIN2FaKfLfqCcvAmSAvLsGneGqoihPGwgCvNP3N3r77Q8wKzo15O/2
IWNcbOSuL8iVpfPCQaXrbWcY1vUso1IFjAM4/4zVAp8DPl94tTAqRPf/j5Xr2VicQRm9+zm9zMLm
iNLdRja32hTAviI/IlgJhEA8IWTaAsddEo7E/AZWgY8QAfY82hZ3Jc+epRXfy9rl9NwENU4/El3L
DRU0QRSwIF+AvLx+MtJWZql26/Wp1/pBK/urJqNhwtJvejVRqBYXRIJaDzwpwBeU49NHhO9JO3DN
GuLnSAG2Pv9H2voDlPIHo6B1k6CzKWJKyt9uIU62efciIB/PWQmcjkXwq8FT7zsdLMWYDzydXX6u
aPcwSQCCE/Oti/GmtL6eq1VlW6o2JLlfyQDDVddRfTzc9HQe01zzvqULtdWROBbAomSj6CyC+SRk
JrbPYGQ2HZ9k4Fah7aT+sHoDYXOcRnfg6Bet5oTaFhfxOKdByJhwcwhYOGzU4VFNAN8G8FVqmxF8
fXLiugOFiRXKka8xzLOlsTOyPryWiBsOQsEiUS9WlEldjhxgEZ91P+B/1lXGs3NcmvfLm1Hq31gJ
O828akjCHtKKXhI7GtdgUvJWPDGP641J5CPtRV3qMlakxbniFHRUfnAAdboXTNgr4h3CuKms8nqN
4hTyaNHQpd9csXhFToEcVJ+lrRo9TapBz7FkfhcrKrLEH0a2av1y5QNVAqTBg02HiE7t8SCVv7Uh
oIAnsBN5y/d+W7GgxWUNwPBm2jrue42Z1Pgr2kkyJvLSnU8eJhh2er6edqTZmRgVxr79o4vWh+dl
rTdrx2GGkPxScHd/1AUbgVXU/9K6rm++ESWSZM/FPRv5Fr08cWY2pSHyy+O9lLIiYqy9ofznz3cA
ilpSrHrDrCnwMZVWKkYUSp7v252etK6956AkJ3B5RDPYsU2EWFJcWrYTWl/yyB1U4xBWQLfZfQj4
zTeJH4965QsqaVpXrlOMl09yz5TlaUz83J9/JO0k2FpjcyJy5iFv/lK58ezSGVpbob6kZF5WJFco
iSwKcYtsQl3wqm0nGQQUlfZSn/9F5R+E/vDu9sJldfl06JnL67X7g0cYk3RdNe+sDwJ2iGkpJxeX
VDd8BO3U4JhID5ZFMfLBWqm4qoLTBRtUyTaTJ+KgpoLmuUgjcOZPWSeZYx0aj36LH/a+0dYOQ9Kr
xnQ9xaODYn/LSk77z7JV3MBCUmSKqL8+8SEr7LpcTArtJf/9jYpLQ5fZsMLFr2HhHhtZCH2LwX6t
8pRwTcnbYOcISJfNzPGJuPSaKyfWVx/evbOe7TzwxVN92IcTNTEbZBtBenqaVYExMWyq5ivDdA4N
ZVXLzVRe4lY588bNWZm1f9UPV/bjkl5RlkGjixcnpa6TfqJ7OH/iRD/cgVlxysXtPcug0hoATRqB
xufCIzVO0f6kWqDoluTzj/guMjZ1cG0W97lWEer8wYc32HHM8IBisXmf1wwnImA10GJbfD/aOXHl
I54lPK1NahhxChBU/W5ITWxSX/rXKew4rdGfh4rmGN68m2/VRxiRYZpk9RwXNdTA0ZEDIyy4T7t2
IWk1tf+RyozZo/8vQOXIJyFSAasvf7vNYSsOx/2RZS0KT1SgClTUpOZHWkBdEg9ahfYCa4eRgJUU
8Ubfyy4UoW4h2JOFPuVHumxRqYpxyS9EqIhp9QWvukmHl5RD5xf6j+Aqdjqc2JbqNojNEk+/pj46
WypxDSW1X5gfB9OhCWqVYPejIbAUZ+9qMkXkgq1TdbajXXAzUxCWugbf46yqcE7J9hQNqKqQIBT1
h1P3ZiE8z/XOl7HWq/rdoACYEqhcW3LNBS06jlEYkyzY1qxxGdNXH8ejdAMaVodKgHC3qv1EZeeW
ACSALucp90KAPkA/bC4ibvM5xRG/1NMnOZF/eAoZMNc4tJikTcmGGlnXd0eZbGpp3XmWFN5k2wxr
0De/AM9VpqAvEY3kiwp8+c3uz9Z1Wgf1PL4vb8fPXA5v7O3wZZ4SEglzg8Dn5jT3uYMZoIGhPRa8
j3FAmZ3sqGwgzbJgOfl87XrYsbbCWm3eJdcBp9qyn9AiRRPC7UuJssi4oyvcg105cU8LBvjXvnZl
yjz4KDytHCOYiontfN8dwb6w/704mYGF8hJPu2e1H+7TreGOuLmXa5tEvmmFXn0KUH2nb9g3pk7d
T9hImr1Wio0cCeOO/blzhRqp8A6GIwO/6ZGS5G0Fn67H3IiASgfk5nfR31PEL41UcA+BbfQorYz0
O+oN11+S7qNSYOlZTsjqlWOXWkdIhLwMPs9Oel8ooGoZUnY2IzU4yssYfzcQ73PC2W573XDgzgk5
npJdmjZIrTOmUo3eguhK+202H/PTV59g6BCihAvQIihnFTbeWcncblRx3C5yhxjwWsWCdAPN270F
JyqdBxJo/oCvVAPqtuiwbI4Leq9j8mO23x3EjUXzhxpPmWcfRrh58xOTctki9Riw5eNMsgrjWvkh
dKJcv3cuCx5+oJ3FL339+UElL0GFheCMKX2oX2NOhMikb/Jv1NDnLY7BWwKZewpHcfNSod1HLn/z
i1glQiDe9yM5VDaeMfTzS53xOP+3Yll57vIZMOHUn01uFKhX2obxX2iI86s5HPpX6hL1aTnm8/El
/sYu+wHtzGqWFhDrHWrdgGZ8f3VCezbF6/QsFiucs6PulKbBImv2XYJe+ummDJLnOOfLIuJipwHN
tXFwBrPskD3dbubfJU0Nw0zeMUmidmcexq1/c5x74kCeJ2tmMV0D7JXGcsiGW8fP4ZdgDTH7466b
lK9IFyDpdt3aWEU77HOSmbR5JUhIiKrnxQsTRzFJT9Xna7fdXvO6I3+/Jc3E3GYRgxamMQYkHd9K
kCSC71zGi1/qV/JguLSeVuYNAWJv5pyAU5t0Z1rGO8/5hYGonmeXzUp+Ak8CNw0kREMQmANibzDs
l4iwVWXO1wC9RnUzJTIHqiyyU7S+aI/DVl2+a0FCwpJRbwYNLTc2JUjdKsTNSwcYQf7irocOrJH4
6bs+AzCqzOyYY4sRzaBMCZVOlnkxLJFVaoMFf3qLyKluP+Lm8H5honbxdJbUXZFQA28QvzfkEDan
55JNxgBzQrWoxo7S5RkUSdGfTSo0fQZMXTE5K8skfn2BCtrXcJ+iqfalpcrguIaqi6c7g6BLCnHu
BVDrQbK1dCMV5kv4qb0YkouBxrgHkAb7hU9gvoZj6VYDF7SVB2aY7zpYfazcnnLMZPx1M3FlTe3A
BIoIHmHmIYMTstWBuqqf62XsGyOIAJCC0n3zuyZZzbUbUqMESvjTFqUWwxwpQXX8vPOPP7Ilc2xY
WwF57ll35DLgK9lihW6TZoKbLq8BlAJlNm8Oz8C//cN3aru7XTm8Y18UTYJhO2fJnK0k1wJjIPay
Oh7QUUmSeBUvj9tAfnL5M4CwFeufbTVG3XktnT6kx/Y1m3z3ao9lTGD8cLYQh7Z/71xikNgqbnrr
HMOdmFfNzF/AguguqwxzSI18ql2pxmczKOjb5F5+0x1Kr/kAYOWR8yoSKmv5L9E9BCtqljYYEbv+
okLBPI3k3c/IR/7ahwW+Qf2e/j4kjxJMhZ1cIG9JlMWUon1H6jZfAxtnKn+RtvA5yzln6ouwKMfQ
TKBDC7XdHCn5yR8OrVbUY5c874e3CHGEmS+NcN1RvGV3aE5pYKh/AJHAOc2kQXlvGup7iSmX0u2q
3O2lc8TvAq/jA/k1lpsIbuFS3bWehtaL9zk95OKvIqqg9ZxSloWYO29A3IsS4bnL2XILehpml7cd
cO6kjrQpDK1dtZ+QeeKXaAAZqUMdxRdJIhR7Wkr0+qqsLoexwOWGe4TI9RjHyHvHMdwWyX7pIhvN
PlYu6cHcdJdYLasR+yBHo4pzWZVPatx9xXC3L3/ujOiCrpg/m2qOf2hkA6ZXZsXJ68drLAs+T1li
63qMljZ7QPKJh2MLObq3qkrEL5HU8IcyNtwhvrUqiw1BCuO4qkh5BPJLBCE5r/le4Zof/esSZoPr
TubSr/AFWMaEqnvsMyCOGyUmiHSOv961U8ObiNA8K92dTCMWPjU8k2KSwrImvCV3wtdzihwfimN1
jIiRxyUjKKg4Kara8zayY8sE8pxaI8zQhRSyPjiV9XCDwK9SRn4C7YnxuLdG8xiwPUJYibavTxJ4
OlSwCyl0SBfDHrwF2ojXNQf+tPnlrODTa/p1EVq2OqoZKJ1xB5A2R/ROawCiegaCjqv1fhz0I337
cze6TIRd6sg36NXXtxZaA2Es/L1mMR5n1up1LCVa3ACxopILwoJAPKP8cJc48vnkdNqUIU6Bajf/
sN0UzV9r2n8tBYTIspB5Nf0WzT1V9nr4cRDl289ObjzOAUko3G9gqumYYIDVXh0aT3tXgrqA9gT1
4z9RQcvfBKuRq50jic3IhrX6RfQfHiau/BVB9Ut1XkUpSHgFhT54jzHVV6phY+rnQUgFd4CY7Y/w
w8MIRoAy3oR4a8ACMuyZqVVoHoKGABiedoEtMu/zzCFxKIXBA+kf8xkG5mTgJRyKt2iL4wIaTPBQ
BiE3dk1lvEFiQOBpzE4dAjEJtyjh2/3nZcIKiq63sPxSq1ZWnimHKler0g2AUVNgQLwhPHQWc94N
2Wgoo0F8VAZjAa6OJ7jdy+6r1PQYRbcma9JKFryxqP7wFWiDP9BmlLlp/2rthlqK+MJOXah5oXTX
2JLmu0c2pFMs23z/atpl0o6s6CqNxl60ORaLqftBud7oum+dk2MEatYHZUTciHSJhb8J6HzgzmeQ
djNruwiUCAU3lblkfOohQgktwb3VRpcbcNJIj848ph+n82iCpz5LW7PGrlsfivxj/NkLDHVA7g3D
3FTvxs0RlrkFOTxELLgrbS4SZoVKB9kIUEvWgSg9tVWXA/MT8egTIWqhml/l5szQHKwcecrCxlL2
nlaO1ZYGCCE4fLfMDudTChv8idQC8q6FyQHpsFiH6Y2OVYLPqJ4qnA636AsVUPV+jFWxbAeIUsOy
UTOpN14AIcpVBhgqrRscvOcr45RBjqtqMVXW7lRzYAZFWTpUTAEMiJ+epHTyVOeRX3ERdzIQN+PH
dL2j+2EG2G9447HlcxKASsY/JEABmiPRCkpmxFwb8QcS+4HR52lIiy36N/IUJM6D/rfh0rzhUV3L
42EgTjolwPpPlPDQJ/MNVdpV9sWPS8PbxQVfc1tsHWVuqjt7CIQGmFCNY7GlvOosBHG1UmwlHrAU
xlzMBUjj9jBrxZsTagQ5hfsj6I9mjifPaXOifGe0nNe/Pt3Dg5Im331xLp5zzwRLfQBRemKPLkht
09hg5EOzD0/sXndqN6IMx5iMZn73/bVALf4p+6Z8VZtrjcxubc2hXOPWcZzUD13SutN4AotJCdYF
gJrbP2jEUaiNSfJinmP+kM0ieYpY9a72VWpiD0YvLZhuAdGJyTY1Hil4RNf8pKPEPXzsQfhb1N+U
P/ZUme1x3ZHbAUK7Iu7OQ0zTXVF+slt6mQUWhrL3CfjQiE+ObgYwoJI7zREJqcxRU9ZWyLXCH7sK
9bRuTCIaW5mdv6wdEZeAtNduHE6vtdN9ceSMa34l66Y1rQ/KZHsNvk0f6t6DMCwx2HfRvviTUUOI
Po+XOib+y3T6RK+h2/iqSa2FQIQLInRdRAKiwAxjMjOLiKP4kXnr9/XwEbr6r4IaKic2UB3irQRk
dSn4Y0fqbTPo+OMC59XoG6u1Kyue9h0WRRkukyMQq+c1bs0XgkOGY9Ct722e45g7rguX1DO7FdYs
qqld1y7WC2YOjMBfEd45jt2aqMONl4sXTbrHcflS2S98ljk0Q63V97bM+75dVpbLWlRJGqb8IhAv
U/EM9iMPIF51e03TZzJgXgSLp0jlFz3g+bsTHHlpSfk07J32lCUfDE4a8r3my4eyACQF2WXSJCkZ
RVcgZ3c+pDJqhIHCDXGxyPZyvnTYBfa0qolEaXSUKe/Zzou4RJHMXYW4mHUoaOwFtXPAtG25LuHY
TlrJ5PRxZOAlkSmHolaMG1qI+9y3neyTJuFOdOmZQAXWCYEE2qp7R22nImVUqz5aFmQEtXnZBcrT
uM6I+QFXUMRm6mJXJPdcXC2FX1ZXJwxzbCoAXii687BIb7bqA4w4cmVhuLHRxlye8h/Vbr2DUie1
7sNOyyinBeOFqGVPbhndFVXlyya8/68z8J7VIKay27h3WnRxfdTu9DW683zM+smsooyzufdVDaB1
QqCDQt3F6pkqiM1sDO+OEZNJr8k9RXwohmWkq6dqpmMC0Dm1vg5cLdf7cXXCeavVjqV5TKyzxaj+
CW7OyPFzM02iKBnC95TbC0fSxKtb0hUtSAfVamiG5ekojb1vqWTOQD5qvwo6yfipueG5hrUuv7QN
Ae6AAoShYMFz6vmc3aBxtmiUtYq7IUkipiEDUMwj/kuPKIUTXC7J/N7+PlwlISDVI7sHEuq5nuL3
PW2MmGb+wjZtGkLtILXoAn2ceNBvX4As2Puysq7BkEwhQQ0nDOnskf5flZ7PRo303Rrpgug7OC+c
x84Wsne8FuCV0pgQHMzQtlL9lBLsaQPm7zg8foHp1L1b8hsBTd5kYDhUrPQGs9+pScSZEYUvQifQ
GG2hrpG1zGGsMJQpc8u/B/x9xyeaHnEA/7vQtF6ksHSOcFAKq/MkEtLRVHo2ruKq9OqPiydEiupN
0Z1onM1PqO4cD5st3m8dR2C6HtgYvqxqbWC1rDotNokl67N5Q6uzjGgheAoFb1R4CJ1Ioy1EMp5j
o9E0or/RxGOKbJj1BwG+j2h05IwNLS6BchNarnF9mK3ClkJtP3CvBltHB+wwQ8Yrma2eytlbFYPG
9z+q9zbJUM56RnNoDhFTWFGqWprAF2fC1V8R1ffN7Nniuw0HrjW1Chi5QUvgejFL5PQntZqFRLlg
oBDIG0VVNgACtImJxun22PNNFANJ7TATsqsRVjxOSv/lXzxCAQIw6iAA8Cle7Njm+KgtUCMwmWbD
BvVKER23AQGwhTLPBx4XCz5Lk4calOSrvIkEF+fgM7n2JGDXKy0sjkQ1Wmx1I+m89PFJ5pB10aWT
LiS6Xp0r6iyUPXAsuJqVVx8jIO5acB5xb1bglElMWlFnKDL1ujg6jVqqLS2XHYMWE9/U0Ni8oY3b
FnJLRZTLuqdkmiWUF/HfTwBfWPIG3DYjjiE/KwH6RTPtL6AVRj7HVjq6MAQefFuNWkRrZXCN9dpK
nEUCAcSThqdybXOY692M3mJlu6CWnG/yEVnwSBbRHtyn2xTQd9GM+cy8mRMH5AhnCumLz6psExlg
I3HGDSd8pw2c6teNix+y8sSXAjUKHOSDaKwyQuSqrHmnjav9oXtupcnUDo055tsUZFtMsIk6PlKL
u4S8zFOLNRaWqq7rJEW/wt8d4iiQn7eHw1EDDttRqI8nh/khQ52FJzPA5jUOyNtjUTxYPLogkwRp
IpmC3ZWZmKKYixb6szU1vyW/A2BHgcws6ckJT2UrKUv+ABMzf79dSSgsxyOKpuutdoRgxwzG+J52
S64rh7FJl21PvSTRk/rSJENFhpx62n5FQ1gE/1gdwfAjb4uBYBf+vMpunfhFj6eLotgzkxQ2MeB4
3gon/F3Ym7PuEN4umJm5m5vP6VI4utBAwouo3/Pmoo0n9YKmLvylBHgfU3doUX//i53DXuOQnZOs
dgQ1lXwpnUBzmjjByr2V6YSQWJABhrRvNwf58OFO+O879UVW8pL46AvxwITAaMVfr0bsyD+wqgOH
fasd1TeLR2fG+2HhTHgTQoVfnMPzrhHtqp+bjVkn7EahwpSeA2RJhGNx0y5kf+A/4ufwy1TGiNcV
ogdlJnqHncKZT8H4FY2zDce0KioI+RoPXhA5l7FcuFCr3T8St87iKzN9oPKXqm9MWcUFCMD0IUIF
TW8guC2MzjWTYYGWGREiOs5N0hRII64ITPh6+KefKGYnzpa7PvmCKmW5qBVFCoUOYkVp1/dIDjxe
YicF9FyIYbJKZOuT5F2ihQSzIIp2Fg54B4QfO+6wpKbWiMsC1QxtvZ9B/iDV7kWnrIIEta1AzWwD
FQuodMI/Re36vuol+4bNMiajjPDAhZGXKPg8nkb8ygPxegdqMslcZQVpPw5ivUvDO4eUQ6pn7rks
aDUKVLp3x2wm11QKKMU+rsMKktlQekr8kxhMBwIw3x30ZBhyWrnDAVcdY5ipkCX0/Wc69BbQ76fG
WAlN6s6OqaVwwrY5onAb0XDLz3HvniP8XQRBq1K8awbQHZaSNxea7LYESbHFJxAD+aCFyp7xitPD
u5QkDpOiylFYp4kcEF9rrBjryHgeq+1efhPMQOiund04kD6TAf+HROz2Gppf4vQZHzs03Z+i+yIF
8nQZhLjkLvN0lMkYMp0n+6I/tYIYXIoW8mwgDOW8/yg5QthE+4fjOVkRRlc1HUKrXqytkcXt0+1P
umzASSK0G+kTK8eph5wNRhXpXHMbGQ8mN0SU4pMgHUlhtgVFKXIkheBBJk+49OzX+E0SjMiRdMrt
armDZUkRL6FkhM+BbGkTIEpD6lzF+TxAQUx9eTHzeyywhaO8IzIi66EVUzY7zPz7OcZ2E/GdCleb
biEFWjys0FMAos59bzt1CNXqNZoB5LVfh4BWczalzx0nBjpFHJwPJzhJClCclfuwthKDDC+yISiy
j+J4kP5AQjhOYEY3dBCtMtI5hkb9pf0PyYCS0UzZqz4elpANPDC2js0IaAp/cwhYakP3Po9ypnr1
K0LaLaYrNeM0Dr6GpulXtlDzkFrwHxk8ZEcSQ2eror8Ct9s2vGop4QjYWlfSZY8Kly7y17lj8zoj
qd0l66RSItyJgsE+kkNn42hFuUC6+gdKGi0rpWJHe11BSBc/UAih3ZeSq/kZjGNzOsqyU6xNjXSr
H0wtAOrApuhlyrbs3hOPC+4NVkY6Kyl7Yu6YMuy8P5c9qumKmoBHLvej/P8atPFZdJAgCBM5ysJc
HuvvizVUVZ7pnVMsaVO5wB41MCFL43kzb51JizM0FT6ZHOnpWTiDBnwKJtqu+xaiSwTJtln11gVY
auYPHaP8xR3WzFI1cDAVgIJv/wy8IDiGRs2EOGRILUOjW4Q3IBwAKlo3EGHjMUhcte0+YzxiqaPL
Py7vhBBVk7uTLbOxE/UFxV6SNGLLikANfv6G0VFI1TjTa5KSslK90flv4IOPqVcNo2pItef0A//4
guqaebDfhDAtGfbkf/X0v5lQtkT9D8Ep1B+RMaeRd0JW0Ys+IsDk0j01nyg2F4oh1FRlGLs+MQTo
B5KJHNKXhmrkh4CFenv0jFCnvCcVyj+TeoPVuHvjw7BX0tp3KHV9VnnHd61ZHIixJDSXczP4EIDK
90imdlvXl+n/PRuSceFNnD3nj9oQOP2Cjn/1ins4sbtRq15PwoWaW5qgvthBkQe9JD4lxLbZJRfO
Aml15uNBekYTKFZeiZRQOhnYYbqyilgs47ZF9GQGMZYuRKkN5tjqGN5FMbHY39Fm4D5M9Zck3fh2
ks+woPoQ7tDuF+kMpjkxMhNbZIkRvkUNVx9P44+gDoQk3D/T7ln2nI38GL7Hge+0skZ743sdndWH
rG0Rjs5nAo9TEarYB6ktsihEumoByI3BoCkxovMLyclA+Af3kvhBLPcSCqhPOmNgrbkDPvf15jk/
F6kmBCYmxlMe1G65L1E6JIU9V6Pm6JmuPcO+sY5jkpsnr+NypE1Rx9ycQZBAu6610re5oXqCVrrQ
I9oCCObCKIrzh/7jhCTXa+GXGITVw1g4Zkq0daWjsYpk7trYAnjafcujOjZgFcazrJjF8l3judoq
YifgA59cpgTfjPq4FrH+PEig4OfEQMYCq7T6nPP8XSw32lmEd7lKy4jxtaxbheK7pcQue/2Kle1K
Zn5QtqbsKAkIhp5NAteQ8HGcOmYnnMa+TOtNg/CoUWOv6mp8e60mUfzN2dkN8uWkg89LnZiV7VDI
WNfrUcb5M0hUS+saCrLXQFgvjx3McGKpK82thjOcKJY/npVGtGvERFlMIn+nwGijiM85iYbjXjnT
jhGrFZ8RUKMydPuwJq5t7+VEb60GE/jgieI3/2XM89kirshsTtEUt28E5StbBJa8xaufXPfopQVb
peHZWRacAFYIKj6k1vUPQGgsCeTYfo0lsIALleozuzMrTTjVvly4MyEGbCtH5G0WqynT84WDP3yI
P2VB9E9bgPziSb4OzQJkWIt+uLNnFK2+t1MhAZhprRGL5GAhn2HpndNlWEHHhUzx/nvmGQtM996f
HCk0gAObTj0INoTK2nHouS+fSFic8bEGBhEsx+ldJmA/Ks0h/w6HOgE/YNZQyh4BMY7hKAZ1waAP
Q2cOWZDJBdXJmsMNDKmE11t6j1zM+4xvas9DRjMoi4kdS2VIMfxTFpHnUycq9U1c7K7Sp81+kPsm
4qiwejeq085scCUVyMl/QiDPuqOBMcrAl3D9hVBZO9JFNekqbsPwMQHxaq1eUGF0stKm43RmluCk
4nJSDxz+FWp2hl48QnaN1jAuevGFnyNcmudnyrW3r0JiEIOq81QoZn1+IDeoxdoSshO0DDAFSzAU
u0eklTJrUluJcpYqTgKU9aYnKMEmNZGjBgWmPQ4sKDEpZyLWhrNXbpqimBZJhggyTSIG+frL3xkw
O8HwKvyKoM66yUNvUST0KFJKUxwzpJ0Rdx/jlRmCId/1gmTs8OFItRt6C1vdYRDE7U7CTOP3ueiJ
rY2rJmrB8ieqhrJfz3avmr+TEJvczw6p/kn3lLj+UhZEWqGtygItmxXiflABZU50SrhmhTWlACwZ
JsLShan9BQ0zVIk2SBwSKs6jwj/3VNbNvQ1U4PLH1BR6hflqHOzKONqFDYPuta2vv1VS1xPB7uIa
0jwmOXr+GPcN4vGfFZk4389Yeb04Rrkc8vAIr6RE6NZVdePfrbz31rTBB1JzzxOr8fV7JiOUjkF/
pT1MQ6qjLE0E/mH89MMunsW3uI+QpkQ1cpKkmyk7/QJsI28G49xfGFs/oaZaKPSZ/Om+kr32c6u+
h+PAdpahspnjj+cXm740Sz32fJ5onzZnE1cCZve3OQ9izM2318goUOIKQsPq1gZExWEqSVlpzHlW
onTvgtDvlatQ4t1wbki6bLBdgbzWThKkn+j5kHZQTV9UIJ2Tn+prZoDjhN2v+otPbbqBfYeY4SaX
8r0o91jX+gIwMSOaz3CTRXnQB51X9yIPsoLn06I/5/y2ig7VGNa6qK1rR+u6NSrlRZsQRb/yabIU
93muv0X5hNSp5LXUnyOfeDmBu5vv/younqoGd6rDOQDrGvZqUlzA+EwKZtYvAYg9JB9vy5MnZiUf
1IMXT80YKBqKoeFnG2Y/2Ij+laKgMF5z+eTwF4PliSlIyHvq/6uxV+zrBA50CdxmZx0/iZ+cSgtz
8uT/PwlHKYvXQc80l4dTk2lAwoChot8YKb67J/VVkWhOgjM9KsoMUzuKYWDKRT1l58m5B/XOkdMu
RYsGVlWkranWXgjqMojeC57sIIEEjfNQW061eKzy4zc9wrzCee3RtsuYHrNgSbTf9lZ2OJXo5yzQ
kMkI1xI7ZLhl3NKjd8Q+QNzzHzwiLZdNyOO7uQ1ByqhH9tvNURDvsgDgoi5msvzs+vGfQ1xvRJcp
QlSjXuoQ6YK2a88b+lnUT7/FjuoYITKkicE3Gosy1+gvs6yXsqseQqtdFieoyrD8xCBXoEf/h+DL
FTcP3e1vJ9wxcVhuFuXdGcCvypnkl8lIv0N2NEaq8zbIKrosC1EWInxm3ICkmKxxUujp4Y7OiCR5
gULenjGg9cFpNRud1R4k4m0uDhaZvHmZL4SiUHZpPbNZBlw4hly4SLp8B61d+wiNmFWJ/Z2q7bBa
sNgGFfO2IIWCrUmulQ5kRxnvB/hWBBN9G55r22PV5+gfSyljeDjkDmAqCiG5hoHL73ZsxxBcAyID
PBlGmto2itHumPGgo7qu9s4T42/A6pE8QxlkFgSfGA1pmkADP7dSvPiAm/pBTTKPHLNL6QQhjS+I
ZYLxTRGWexWiA81iygev4o8mYtNvIqsUt7OsB0BftWu5C9fGVlqvACmwLP3zuOxhEAXxfsqzqIuR
GKgFhsoFFTXFsyWBAi6vtLBnsdjtP0au0A7jEfDjVGktYkDXdwe3vJFd1Nah71bd7mhUqk5IVn4T
4z0UPNf2m8J+t+DrnpcaRD3dpOaZcpGOarRzYcwKch3nZuKKJeDqYf/82GKSWadDO0DMAwho65Mf
w/ssv1LCtIOj7g7INXKaWCtCL2oVR4KVkzSeL9/XX9062/lhF0/9GxReD8OBApXhkwm7Kjmxxhma
+cQg42qiDgbmLXa9L9de2RQ7/dXjPjn841ZNSZM68hpphKNC94BJ0jaOKyGEDOeMg5CI/gtGnRW6
OurRzaax4Tbw8E49VJzDIhoRuJtn6yw12YiNrHxV7KJD7lVyD/Wjhuipl3LpCN1v1Lo7sSLhfh9t
rNzulS560EVfNgK3uaFwSXB+JKuFxLPbio6/0QK8cwrzJCrV8On98qmg3fmHcCtMprK/yqLnDXFS
MxnL5x3NqfJgNgyC0Q28I8OBdZUOliZykWihWuUWCTe6kD4FmdZIGvlLEETfvKNAe4qZqA0pgqPL
Pyv4Gpp1GuSIOiB3/4EvozOhnQYODB5w+2/C2AMipAplvSDITsuzrtl8TrlIL4cuGRMrDk83jsP7
T8/64ULNUGtUNbZnwIZ7zAYZjPDf8HvjXFPoF/GYn9VqvzH2G91e/3jcahvSv8sWc7d08ToId47f
gA6/rvrKybhtA9YW5O3c/VMmV8E9i18kge3kangZyqhDaMvGxiaCGg+RHSpL1K8RJ9ti8CgWg7bB
+wAlgYCbJBtVP/gbdqEjzazr/QcVJZ1NEIOfn2TK9xZ+kF9WHfvOwUSd3+QZ/2H48PCFaxu69D3A
yezLQ7nJrbEao6vBtN2FDGPIkyGCDKzvvUxVw3TjCy/mHbYDtdWlZFgtbZRn5W5ukh+iNYgdIq5m
ib5I3yXM+Z2JiXAYAiGP3amlJ95AP1djm7x2WYV6t2X087El04YDUwCRpJ7v+pBmHmZhEySzcS50
9sdv+ojsUaSKQhiFkGm6RBTQ7ldxqM/qFq1iLBFsLg0melO6jvwRIdJVNgSaBoNR8njOqvlkea2c
HXC/TrtxzYlL7SJaRQ7l0XPjTDK2zaj5Sd4eLspq2sFviOS6w9wfewqi47DczicTBnJgp5JDOE39
5TuYTbwZC6AxTDzzYha8bhTuHEwEGE99SjzgpUNB3be8Z4zdEl3h4Gau56YCoxFHJ+b7nd7P6Hp+
AuVM0WduXBNCG+TDStb7Fqo8rAknDgRMVfiGAenDfuZTzdfTWuUrEaGOnzvmY5oBjTXyHn3AWDxy
otSrZUZWhVC6u3SYyp2qcoLeTws3eDsQQ4w2sZFqmTgmynapXNQL1n72bLuBwL60Pb0mtvUIxnDu
sdwR8QgtuZLK1OrvLvbe/xwPh587FnQ0LkD6bNG9k+L4ZF/MFDDpatHu0OVfuI+3d1WO8FhKJcBd
R2Tba1YoGGheh4LRjZ74zJsDAxS2W6JRS4p76X03fZQcRMaoekAMF0fZEcwSauFBSwsnYV3hVyV6
YXGG6ybRUhJnhKvxsSp8IJvW40asecVQw3pFiTEwQzbs7GJgIUe3qKZ01IsIwhgym/713Bna00F5
0ZUPfZOKBQ+ah/IysWkktmLcawiGCxQIAOUcv6LC5Z/xMOuYG396ndDyXhm12ujGptTCC5D2EhtT
hX1MngzK1GeY0Qreos7a1r8/ljOWDBjwnC0aJBLbNe9bSsQY5lqXo4hTQ20bIG1ltTljvcIeyUOf
BuF4lNoM3TxxW7YeZ9KG9cOoydIPzC3UZQjjIHVsNz9o++NytkK2PQJuoIW6kGyf/w6NCwzk7EgA
dsIIFiyi9VYOUqHK8+eYpJKgl2Xw/Yh7gfqxKOD1ALiqWJk0q5dLG7nbjdgGN/R6ZdL0clm1Ojbj
WuELLcvhUG4HltYwD5bWuImWCN9/gwshHvCfWRlxovT6Cy4N+D9qd78mL4dlWZfv6YkDJSekJUAa
ZiUuRkH5MF5cLsxSOuF5+LJA3nz2XWqZiweYFRAfED7Fi+ugIsYwt+mQ+tz1EAn5WCDSuufbduCC
ilvqbIs054gyhaopWlcNRMMWXAtGcm7mKgLjw0jvs9MJbeXVwd9ZzqyPYaIVxNJSUKi7wgmOT+or
v7INgyomLUHHMK+QwnNdp4iQdT/I/xd/4x7Vg0SJ2xtrOwGKxuglf31p7i1WlQ7sFqflbeffmlfD
h0wATnJsNHcLnre6DeZqOSblK8GeGC7gcuuwxnxielqvK9d63lVXb+qjAfDCM+2WgP9yG8Mmhwpq
lVEmgImHjiv8MKqTztAc1PU8TOCL2RIgI5eOVr47vnj2oSL3pyO6kgOOANvVs3IykdfQWJ1YsvD2
2evdGZaMUTa65eHehI+WBf0k7pSOUc7LZhwjiiDnyeSMUVuRNsTnvUIXbDbv7blwNnwW3qpWpanO
vaRt/fHFEeV9P8I4iZO/lICXB8symuq2YJdAK5LOL4A8PMFb/MDxzOR4lZG6G4Dl7ZsNYOjyqJse
Yng/4XocAZxtFE4FFDR+Nq5lbl0GlBNDs7CIFJLA/ucexnSnD99u0eYF76V4o3g+JKvTnbkySgMp
4pVZsrI94eoDe/bWLdVjtREPJDYHf2gGTr3ILrv0QU51Q0aC2fkTapID0OhLnXl32YHtaZBtm5EZ
Bsa77qJROUIqDH6ZS9warCWyOU4laJk0uG6fV1pPoQumm34Zxg/uv54hbZpicMUt7/3/ZhW10F15
ZO+Q4Hvlm3/4CqJFXpjaRFdjTqxjdMb2ZJiwo2HmdRcnjDZKzX8elfvRj0ysUbGMwPPqfgNnNFLA
M04mgLGArDAanzEEAgxA1KpGUOVwQwcHKwHGSWu918Q5nw9DW01c4ikwL+/e1IV1ZYqqkf2jWZrr
Jrs8wesBYvd4ixi/MVa49Px3cXWEIFfTMbxYHFda9rdX+GWLyATcnQxWxILfPNv/Jes0oW/Kmhtb
+G5ulzEc9MgXBRIHCaUn+8MViBehb/+4A0PslCTeyiGwqhnQA3WbUsc++rYbq/VVdvEH8U3ByWfp
xZB5amttzOPE2z3yFpv5X9/sj9dL2cKR+Z2BgKVlS0C3HWlzsZobWXJf/rAdV2seuc5oPvwyzgB+
pRvwa4kpabQ0YCiRo2L07H6pWE72BaxzG9tMGst8fW/GF5zzZSlgm7H33yfiEPqTy4x6ATag5Xwa
c7GTfX4UTda/awE9A07k3rAb2LDPhFkhvJlt/8BMJ3hKOoh7kT5nF775YToeEfr3/vpc+eD/vO8k
GlAeU5XvnIgAj3JC78E9e6lAonGgcyHpsEdDiUkwft0qrzASFiRCTsgLnRzqFJZubMao7JI3MAdr
7lArgYTdHB5pmygQx+fh44JEJSWr9mrNqsyRkgzvMj4K+xX+SmQQELEsuWtKyJUxQrJYNobqLCFr
8A0Bk/W15x3FVrcyidxIjXLCC3VMzAUu4TVPdZpevXHrh2ZNYwj+Ks+n4SOppZihgaHHHpEZg5gS
gKQNJA5JrJI17gdu7dIUZ/Ei8HbDdNRZ/okHGS0FUbTPfX/beMrv/wICA8QLj8xisqS4Rs22Of/o
guAu0tP9I98eKOHh0WOA7iNuOKcNAa4KU2vLO4hCy4koGPe9uXhK5jFW9Gznnzx7medHLkVFJN9E
vsWP/9yQ5W+AbkCI1KEJ0wmi7JYZw0hbASOdAMyHVHLTFs0N/9w+bKYxvD3n1Tx3GTj1KQi/+yiT
74EJ0FGvOnpZLhxsbrbU9r7fXyH7lcgsReVxbOsad+h14/H1r76cI5xMFyT3kXgWscw9ay+nxE0b
RYIFmcfWzYPg9YwNu2ws5xyOrF1JpHNWJaJhYHICAszlooz5E0FhXWTFoIukN24pFFQLL1NP1IjA
rYx4aDpP5yT69bT0BvQBDvN2xlTk37bL6LXdIIMbM9DdqgjfYB3Fd9j4+M2nXfycrdeLwhCPUFyy
o6k4+iSD0Jne+SXOC+KkNNFsf2xTkwJlB26F9vkVNzRJoU9m9EhVcgRkmc6uan2FC/K1HmttheIw
CuFGDnHVXU3S4uJvp8BZI6LKwrncCiFzpzYIG3et/OT2oLrjipM8oaXKmlE0J2e4BKgrossINOzd
MlR4geSCGP9ETMfGzNVZ3AYhx1DLVrgOR9OwpweB48yf5f5I2C8tukuivVkZWZZIsN4dHLKYQnHG
CDaHHM4ygaImQlX20h+y0faHi/9yC1XL9L1FKF3B3BgfJbHcpCar2hSEv/CrUWFX6wmMVjOb1xtQ
kyATmdGPk8tuMiAlSqlXV1SAXYLLHvBR58vHBSkuct3Mr5Td0mJPbs4V0BDaiUdodo84bjCSguoK
0MzOtHeskI8QVbvdVWCp6xx20LbHJAqK373gFBUGvathBf40mHUo/xdQzB87hTK5BEjo1ztQdcd8
Xa0on3Btj7jfAPHnCRslKs23H8/rfWOv/DAyHSXpUEUg6pUMKeCfxpyEfUL+/RkjJ2BFnbAWyEAd
H9EMAs9FkX0mnkmxQ5FpoYV+rbVfIvRc9x/gfp1hefqqT9IJz1sYVsljNhS2eOnrkCyhVeY0TpyG
f9IPc/+Sl9jHapZ7vpS8wcqjtsBPorgiSHt7QGbvG4K04GFoDrUIGKf0E2nvun/urUUSfX16FNn6
BcaUhpeD74KsKGGr+pc9+6JfbUaFYDfUyAqDDO8h7IVO7Gw/rljIA3ob+AB1sQTJuYJWVjuDoQpC
ZfMTizHGo+jvbvZVvgVPupKtrbQxLvudt18H+HYoucdCXJUXX8nQN3Iv/64CKg5agqTvN7OqlHrp
DFvWOL1tdG/LfO3yoCTKRi9O/Ml9cnjgCao1jA62Q+Ot+7jsmmmK9Zcbt5oCPi9rybfesGm+jt9H
O28hbJOtxo03I5Zx3679GMykf72w6QuoLjPX0vdcoZ5uyxnATPgFNDVQ+N3G4rq9v3f+I3LAO9VC
XvmKdI6iaBowo4dXF5IWWorhNoTHbuxCA5y4wXig81mPZvR3tgxs4QnbBTtdtpNvin/nKCo6Y1vF
L8A71R1YXqZ4InKYqJUX/cBkBjOc8+5u2dqPF7THHxRhMRs2f+CxOkMJdW3RF16XieulTcuUk3Lr
zJT01VKbuWW17kjmG89yv7r8LsacmW23z7S8Cp/RfG/TX3N1xltbtvcnKFapcjrLMf18+G9IHqqe
kNkqu9eoZ0+WJU+HCZ2+Ltp5nXPNVKY6X6arcDA5kkSySPr/xdwYdasSzBfAgCGtNoP5ja4iMPxh
XlXY4xMThIpkVlS4mA5heSrTTfJQYdE0FA2lFslDbeTjVe3bkCVQ9P8oD16vTrmcg6QahQI5F0N7
HU/QL4kvkXyB1mnj8+OCB4QTjrtqPehPHSWnvP6WDCQk76P0MnvdVtxbHxO7myIK3k/5k6b5g+sz
g9r7YeRVTbJZS4rjhAhREULKwcNUsTv5t+2l8ru9b1XlmMXnzDxFp3ooIgKPoPNL1mfXlYsb+1V/
WOlbzuQvMJ6yC0Y89dzIYHEf/mK3r/IPiBghCCtXvQF0pRV4V4sSXdjD9Gf1iB7F8V1QP16xmFIg
OrVdavfzpcCt/WL+k00KTPlbl9XMkqko6zx01M3stHE76IrGSYGFD/MObzHmHaKQ5rC3kJyJyg/B
fL24W2EzwNOV/Aj+7mj6ANlAYp2hnf2t+Q1ZTB1ROKOYIDo/TzqnMW/OdEZ17eF+CThncUh9rtzA
mmMHoPsexBdcjLqReZ1YnIHe2fw092+e6CW7XylswkIfRJ8R6nRASr7sO8LGdaWarBTYOlGOT+E+
ihoDChQgGOAq3UZRFckMl2PjUgi0tvTOtiLdw0yFPo2OO/lXdszQZ7aKZ5ZB5vZy0Wf8wsb3xE7c
rd7kL9E5ryAKhvY5jHBr2mIJFM1kZXv6oe0koysNwpLWkv+TGo4F3v+TzkekRT1Pf4s9qWCRDiEN
RCRgyC4PAMiSMkubNWhdM8P3N8RVHGZV8au0IO0Tn+fY7dMMiXspcpehjOKAxEWqjhoigw4PZRuM
hEzbSbqxf7x70DqzvSdpo43LAQ/ucWpeP6+E9ajtxfSDV2bJ/3qHdHQr9UD1xc0SiygLLs0XQ0DM
oofs6xn0ijs5Tbl7F0xuAyji5jGusOk2uRgeZcLfOs1Cg4Z29rsG2YU7HlbOE5xGYT2RBoPTPkPr
xCdEMsmh2BK31o+uO3O7xSJNiSwOiew0Rf6IYQVks0883B694RN8ZRbwJxBFXHgpOwp18rUE6T/H
Y7euogJsQIQ4RBkhB2gUSkN6B++LLtefTc8vPVCCrGQgqzA5vvTx+9HhRD8KiiAzEHxLJX5qmOP0
A6/7yYhlfEtr+6poJjYqGcTg8+0/696tv7GwAmsBJXZuoQod3WnMfFaKSs7u+QO0E7yNqxTdrwNq
m+FpsirBkmigGBYeh14yyPUeNiEJAv6xVXO14VFTI9sStEVjGBg8iUssMM8kg+/1g3ff3AMvxDic
riXZEenunTA//1On4Xbx+F6nFIjLC7EkzkkCLSGis+3rl1bE3/5rnxUbDigFZFE1o9Oww2EEVLhb
776xVhLXend/YKpd/1gsDDZA+Z0R9LsdKjxihanPOSfUe5WIjTb4EhboXLtSQ9bTRb1opnT1PYPL
eU6MHAH732OCYXFhkgLBOk1UJyXNN02ivO28F4+Q0EAcoDwfZGQAIb4qqYFiIIrkA8W5NNS5Bi8U
bvtVzAWTCA5dAg5nLdELZBthrVJYWWrSAwFPlqdJFPCankQIChofQlKlPciQDHV0/qnpvsn54HiD
YiD8VdJi7v3b6lcKPcMuRAa2/aJLr3JtU7ERgNKO45wPU2je//suVyh36lxxjVF4lojqzgnlDBVd
vQgm/Jl7QcS39DpV/ZSlh5QRWxfKWGpeEnvKCsOalLYB1sJdFdqRAKIedDCcge/uYwV5gBf5js6J
xzbQHYl6w1jjC7RSHxtU1QTEFbKQHeHAyg2u9hwha5lUPPwT6DlZdy09Kpt/9MSiWzp8xNOiE1Wf
OgfIVln1XQl2c3trJ9wA7Wx1QzqDo6zSIvABrXGuhfAG+2NFjYBpsDCk5RUo8dP4acHPKEZLujPH
F/MOtcaPwOYvIUNXw8pAL4lNoetqiJP/GOPqdomSnd6s0/7IYXSz/vK3Y3jPk4+P+RE4zrHv8QRj
ClKx1y30iyyJlp3Mp0WsPvVLOyp/PG4U3YsqJJ00AO4k0PwQ3A3TWBBJS9lNhgPik5GY0B8+b3zX
SeSJylzeE6yU9pSO1C0m8X30CD/z0RdyFYe918VmyFVetfBYZGAt9zIcrbwdpGmlWCrsNOnphC8m
cOeyYX7axea/JUYb2lQmQjSmmiuDKTFzEBZDVo2/B1c0O4A1JF7gbKr0aaciTyignizd3KFl5rDQ
k3owPRld1ktNZcSw+hT0UwSBOfQV95lIJNJ/7FaAS8QSS+NNb04ZMU4cqI4RPl1ry0AiU5O+iEqF
pxLHwyjJl8eLZqjySK5Km0bTm+MeVfa3TpGpsMQdYg5qqpbUc9Eu10/tsBbZm6/cqIlsldJQ+YNm
mLEr2osoPJsGwZc8JIzdT1DsK8sq+DbQb2x13X5wr5K5Mgp5dudDLSQIzQERxiT5QOGzm7pGgl+G
SOdYNi+z9BtIyXNco9VO4HahpjKV5z13j4WbLy95Uj6A5JzJU146ngbpDTTHsKsMVvhqAUCvVeQH
GZWdeZbNV6ZISF2gWZIUj+S0MFIz6jkVy7ZLcVCWBFY6UVqRqfOol9TkPy3NBABKDUHg5GaF8pcg
6htqhi1KZ/Uha5BQxxGOZ5DFip/ECp9Nwtzh/09psyET9CZwxsHwKV//1CJ6aUelRUpzRBT3e33y
TLhz9Ecgnwus+yjt1WCxqh8b9e9jGTSiFJPvHBfyk2G7znRaj9qVRlvsBeWydx+b0ghxm3BCea4C
rJnrG01coiAJXcqSpjhoYDKOSGN2osF8YFmo7y75XrQNjqDWTi5I1eZUQsLpXx8TOtibKkhPAkCS
xnDOII3RRF3bwJqhcRg8fPVlzKFhqwt93mP08Pj4lUUyvenHf6Onxrh6Zx9FDCVtUsrW/38t5BFB
tQewmmbpiAUQm4HqyNs5dOzNUedWdQ4UFWRn5lBm2UglMxXQFjJkP28a5uoqCbsqFCzQT/PPnwsy
Z4k0rED6V/GRpUXEbx16pdSs75npOixPZ377WfQpl4eY9/DgDJ0V0NErniFt2l8ekZHCgKZU86Px
9ilOi1ow/lcSwcyoVyvIb/hGX3Eg/XX/TbNs8D8VGT2LaWZahFF88hUjmfe8nqHhkI+XV7xYp2nz
9Yqz31NGMaoCHzte27gNpCB4wZW7qRxKoYeOeiY5QoxIweIEuwmVWeFGWJ8nZ+GK4eoBWS39L+mI
RZA25KO4ims/84pEnTcF3AxoCVJMMrCIycjVJwGds4M67/5mxq1tZ33yLLQ2UUR3KBDJDat15tbl
BNx22ec9lAB0yxLjLM3bfybEXM5KEEoQfCwpjokwERemKsea3cg0BC5w6Eh1sn7zAXm3xcsAZO6S
kCtshYBokeETo4xqpeUXv/KT0nyK5Zum6i/PKw25QG68mUOfX6gHjvavmnXfYBI4s5K7KUw9ZGGF
6oZ0D8U24mDiC/dq496sXjDj9V/0tjYIxrcPiUnsuFAxq8O7LE6JbN3sAVOTFpq1ZFxNBFmLJ/0Z
aPaBjdYOJXzpZ1odietLhEp6woyxQnVxLLQp8785kNw7i1jGHz9grNVv6rKZH4KMujDHmhJ5Uv9o
BjKhxsuKmJwr9sRsf6YLxnIIhSch2HpPW23a8+xXMihPjXqvprimVbzhMzf9UGSf/D3Am7ZDsv56
NMvo3YeAim8OU0iid4gaWDAN/WEpuIDMq+YlIC7kT8zlhSxqatGKlwKysOs7bXrBDOTf7SsokbM5
nUN3tb+jtpInwF59vTetSERT8uXOsQK4s9uGfouCkuLnWBb+QNGFJMK5WiSqEQwYcilgOr8+Yt4V
Bp/eAscxNxjsu0bcqcWWEk8QzEmPJctLlzqFKX3uz1mVvX8ElO7VkqhnUmcU7tQy2j42tWZVZ2Z4
fmGw+PyM+SraTyeoPV5mdXTy9VKYFhplDOaq9ZTxLFLOjOEvhY5j2u3Z4ZUHRvuMdBEa8Uydccua
X0Ofe9QvdnLfQrJcmMb5QV35Ed7jqEmZRXC8wj0q1V5un7Bf8mRd7j3LktmPIlVg1isfNb8FL6NB
4wwsi1+nTRltyPo/ZTdQ89hW38ynF3MCxi9gE7PB5Kq7fGUt8ZP737ABPgyDnKzFFRAXu5V3ArX+
lIyHXEdBAhozzNp/WbliyVkw4o9HeDyoi14tO8W+DQ65qFSw2jCaQCQEV4cyyDU+u8YSkoXAtVIS
+AFEU1rg38qzrhCPSidEt2pgMCFGpxckgsYR+fxs4rTSPgacUePrjPQPJXGAlm7Y8ID1aCam7GON
wP0Y8K+5oqKpq1b+Gse2BCx2pVFB/WJl2hPw37/bR/gfPKcpjvxdA9l1E/enlvIeaQmv4ZIaPK+j
lGuwMiDVGNSrAOqv9jsjdhDgumb2/SFASWxhSkqzlbIvwwEW1t6RCR/vQMQzLkuQbqHajVoHgsu/
ETQudZHQG0tgNBEAIFv90UuxIQQRmqahZCnnQF6AtFAkbhAtawE/y72YV5pO/5Hkv67RGF8etYlq
73Hac0dgT/Pz2V9XFWVgwzLslHKeSpJ3BExB8dYqJ2LGyW5sAIriP+1pUzISo142WgzDcbGiebcD
HzSfvfwOYqgDkmYQEj2+KI6vU8LWeh8HgEOg0Ro/QBKx4g3BY2+frPZqnaWlL7UWn4FrHKbh/vZe
zhTrO1XP8hBApB+gTrLTrMZfhHiHgEWq6OarFidUiitaOI36NlDskTP5VRN9HtzTCgOHKUrJnhWm
XtPWIDYSArivTOQgoaylPyU5P1qTkCqiU0w9x4hYlfXCNGz+zuG0rdG215tmGH/Hvs8ICzTMvjGV
nMTRPavbQNT5Vo2mYiQS1wT3j1Qd6Oewy3kF1A+o1qkb93DZFP7uJHSyajHFG/5RTGeeaCORmEGb
ElP79PLwmBdxijzQy1qGmKysCB2yyXlQY254DXH+qukNVs6zrjMbosBj9/Itm7eDdBAxdFD/pzTY
NgRwWysNgpQbdMTNYfgHi7Kr682mbtwkc2iGNnI+hvn8Ct/B0+jbxuvJ4qDRsvJ0p98X8hRfGbHf
Z/AwHre3c3ThTvwnB52tES8/bt7tkQ68rVY3RBOkD11D6xnwYrphthmEvSNU4zDAslhFaQnhhpDf
PRTnaVAsy/MJvrQ9BohVQAgb68YoEVPcWTejVt2d7Uv1JDvrYk5eptyXWOW0nmuHxoiSO8Kxorvg
nRghrVgwucAgsohKBy0x7dngRCM2BrpKagEpUGnwHgYjnwfTxwv9gBdhqW1oIPL8DYyCddjUP2gb
ZP/MRgVKUYddtVK3JFYWwP7Q1/Vkwe1Y0n9WfyCNjfnYC315oiUybB96e93apf9AQCugeMZbcq+y
2/JNBxjXrxC9yXjMwq3prROzTXT8AUO4wMWWtjRpS8tu1/MLwOc9zIWfM0sQSWFq5er/deHaTs4W
mQN/56IXGjDI7iXu9YNZSqa8m/aPBK6iWn3bB8SrjVqVRv2JNKkDLfSH6p1X3y/5bN57FYWtk6xC
kJZGlnjZ2jirGk0f/irO4v6E9hywSjFt8y2C1wSBbjchXW6yKmRFYL5JMeQtkD/yDPiv6Gy9t/aG
2EDs6L4Pr4YgsdKskCxhRfiGcOwfFyYtoQBotBPVhDZBN7SfXgpaEQG7LJbo0qWhb7WqOFvo04ax
EN0xfAn+e4W9p49xQ4bmeBy3WsGJbbO9XmHQOsfdDjU9sttrvBEu0HRgJdPn8xxToqKhmsyoUQRB
bTt/Bpr4ycNCZVemNLtZD9/Tp1+4+71c0Ue/GtiaHRMH0r1KlszlN7GBx2/euK3OkR1fW91hEzxD
VY3UZCEtARtBDUFzZOl81fbCiz1CvkZIBR7mIp8RF897blIMyWPN52TQxOCrjai7ZmbnlpZWBPCL
cSKkucrg/xftExTng0enhxFMhAWIzdxYwpVuaAGaNDJx2Qdd1m7IrE8okRdm8zDIbex523RuOQv+
c7+Uj8qPhCeCEtrDx+8o5FInHe97Ixsf2oFwuCCn7qrVrGRmOr9SgZpueQnjZI+Bj/ISZntcWgMX
mTSv2m+vzbJ6Jim1Vf8troaCVp9xteLZfGawq5C2IpK3fTygT/fh2uCighMj2fj/ch83DkAsYC5S
/xWenUqXQX3O26XH+U/oCe1gt2Z4GFcNE8LlP6gM0Cr5Ic6lfQw8h5+WgLV5i+HSCkD5iuqVxcc8
VtUeEi/qbClS+jS+kWd+1YeiiDG7PcoY+S0CqiY7KN4fHU5GgRmAhllX1Pm2xrZIy4FPCKqwj9eO
sv2kJFtPaXEKcwpxy+c8p1yIKb0rjdZn+eKj78B8//N6WgUhRohJwvj7Sswltd4B/qgmIOnJ/AT5
MC7oPi4kCPbyITdy/Vgu6DXHjSXV97afyvQ5PqnYS4yVW5YQwN3bhU5Q2qmEqEzMSYihzYDQgYyF
6SYMQGs4pQF+XOe4srLWYCRtcSKSCjlNkgVBl7cpwj/Scl3egUQI04S/bxZCc28AsyPbvJepxBuA
F0rPN/+nY/NffYlSgUIWzPlqY2tseXM4IxjvxbGog3PwB7QbAdZW5c8pFbh2n1Eeq1rzlIfb139R
6hSU6mxPj68XPr8zq8mJwN6syIch6unHuphh11SMVuBURAsAgkeWE8+tfEbHHjUzEVIVP/9mU/y1
YqbSopC1demQ5RaXd7DTIhKSZh5PB5NEDookyOlh5tMZ3mzQHnetk7qH0UZ8ZjSVAxFTcFROuxAP
b3iP3bLxxdvRJhv197wD5hiDaXl/CBlUu9nZQPZHJKQoV0No2xHWMoFNqN7ZY7WvH3v/XCl0Cr72
kIf5Se8c44fYAKBHJadsspWcUUCsR21saRmzRQmV+tBs2R3BK7rrwJg5ROVCmFCdD5JXYunVz1Sz
VZCqaa75Qvzkza5QrkFcyYdsAArBNiJ9EyzVBzIHtDl5nDVSj733x4kuUetB4N6NJvKjjTbc+y9H
aUX2KN9ev5Bx6m9nBW4w8bFUVUwOn1ljp6Mnff5Y+N7AYbkR3dPGhCeVcMd3V1IEDfqR4lmbYxvH
c+xZShy2H01TrnSe61CT42q45mwlDE4NkWUOtVgpr/IhD82XeG0Cbbcwm7sn4e5LGuKYaQp08Ba/
zWam2guVdgONJ5ta9726ULZaIk5l3pfRh2S5xNzpVKvDftRoaqztUHyP24UX664C7oFAMR+14svx
zsyWUHjlBIMDEhJsPauqWrhrbn5dAKq49kOXXNrEliy+esnb8mwDas0Ym2xJXybDNy6f8gMbM2T2
OcV11lbWRxP9r1TWpFrwJbTWRPqFgcOj1uQNaKShqNZP41tU8dK4WtwCdlgcB8hVcqLpOxADYZoS
42RyEnO+AdWZMZA9vQN/tXK8mqcoX49kaM6BzafhK1eG8flvYZjyQ7QLrKsHWcmgMh8MUfss+8pi
PdE+Tc1Z66DPdH9vGB5v7EdKm9YmrzpPocx3OFcDyWhwgp8FqOv0WNfn+s031wMshoFraqZjC+ZP
84TDf6YdSOEQQjhoAJjbzbQB11YBphd47qJEdx1jG4tlbY8+8xfaa/7SGNh5JmDCnVALDlXS+83s
QUBsEbW93iwiXzERjuCqDR+RuC4+PczfeekWiOAhFmjZCo1/xhrnvRSj004PPr3tFps4AWvfYY0u
gDA6Kap/Gk6nRTxm76cs2qMNy3pAxUgfnt/z0edFVJJtNLir+/QC4pTUFLCijmbeC/MxBXnMv8St
a8c0qpISWFpe8AhnEgnb1ZaZ5Hql0ohZgRLQHoxBBPzTJSQ++FE8l/S6LUKLNJ6xo4wXtAPvVXGy
SaDBqpEIDCyv23L+7dfbXFe/44WYjAXOywnIyNUWM1qDtqljTXl+w1SB6hS6AMDgDU/pw6Aycady
BNu0Zaepu2jr+Lkkz4hVCz/oxmfNZ9niZNms74oAApNIs21zQQkR1saOs/J2GqoLPz920vW1Nz67
hrl4BAKSF/geVxJ2EIg9GV81auN/8wit61QAqVSISa3HHhBM2f3sMYBdWav2v9EzgaIA6XiI+V2Z
wB8ehp/Ybs3YrByZXMmGuFRN/hZBJbggxCx21SMdA90l6GtoJ+XBmG+suINrAOS7S6mbDWqy8McP
N1eWsT3ZQyiUXZ+aFVx4KFu3idRCtgeOEIxzqmQCSzdao0L0qIPVzcqj85KYDyxRY4wO8kE8lr1l
dtQ/aM0jWcfmF8ZpXOW5B9+BNgiUhuDA+zSqWWeQ5IRaf5oKA50jx/PENpKcnpDA3ejWXg2abHzW
7rg+FAU8u0QsbktnYKqxQasYfQtBUDSIxgEtOnf7TdGej0AKbdA7RRaqfML13H0JiqE2Dpsz8FTz
rsvsW7Hht3yYDomf1oh7QIkZ6pZONwsgHtyf9pEcCG/ALzHsCzljF5gQdan1UdskBHzFdlDjt32u
jCKjG2v4RM2Tf6hoDprS8xWhEYB3Xv+fcoNOgM32vX1JWWL2qFptqc1DmqFC/NR0afFhrQoxoWLp
Xk/L8J79cYJNia5/GUOJtWO52QFihCXgZ+jiVlq8k5YmAZYKb3vm1BggBrSQ3MnQmxY/aGpPjDuq
h7akrf4PKF2VsordBHle6DlbgYoqlPatws6UW9jd32JZ8XxC2raUdEb/m3MiedT0IiZHpGPNlpHI
zJyBDw0Ksh0lHGUelOmn9q3jMkoDFWD2tmAadIcYAv0ltQ2NH/PQRuYAy8omDn1ELuxVE6KfRcs3
CPlMAqAuc/YCdx7kcsVfeawlj6xcwbyph88hnKrjOBP7pCfn3hD4k/EuAuAqV+K9qIDEeXXP2luk
xW5sru9TgB0LdZE5mxozcYhinthgfAN2MYa6ag4oDUhoCrEHQLhp8YOuDrlDbybEannpyRJQZdkZ
CEuLo2oOrqd4OLO/LerOQllbMrgQ4Fj2fMzYoxxqfJxjSPEtak78qNzILhVswPTRgbtocsK/X8+K
55EVuXJ7byorLZXUM/clV+rMTOG6j1Sm9w86meXyaSIz8WSVNOG7c1YVpOxNDtmk3HuseLyeFdX3
pkgrc9ZxfLMlfHpWFZv/BrJsuw6Ad5XzwqZTz/xlgGp53Ipu7V1Tx4IgAqczb4Q9KFjY772LFOUw
waXc0LfJ9XVd7GFJo9vtGyUjZKOdZv6Xhn77ounEKUvHzv8qkxGIAM7YRS5eNZoAzNG31qKJBfUi
QOD//On3dLl+UICnI2iSOB3P33GFZtVZbum9O6baPlkdHSuwVRsBSMFn0wrJ6Sj/+qfHKseTdaEs
BNcQav+hRhxmAmYg2r5PlqNuRkBi1h58+ieycDISEdXNzfYtOyIuJnc3eIl2a3RhFiA/olVuxP0Z
akVEH0Aqqc15aF+oOhiUZBdifzyeTkBYeXZnfUcDIP8zp8Vq8vU1HHe1xdCRcVW2PHt28Y82TBHl
UHXCTye81IUBbeNA83R5MrneTWqVzCtNafn/CfRS/fY97VJSYmSuX9yoCzgow02z5TOLXGWFnGCR
MQry7+cHCZt0keSktUU4nyhWS3e0aJQAsVLa6vRUc3xBlheHRdRh7eSZ/daGKeKUFLK2ffd0SfrV
KQ9KEqvtEFcoskyJ3oZg5Ak3BEMqclcjfCdXClDqIi/8Q96UXzYHgmj7jcaPDp4C+DobI99eQ2QP
qKDEYqRJdILwRYDKP3J8VXYMgdxgiav8vPoeDhQa03gCaH7+ZhrESWenH+POq3asRFTIke0pDyBV
TlAPzVr1tmY7FEtoz+i43RqJTtDmmHqL/BguC31PmkiEyC2qbiBbQcvNZlSAnFjYW3qn0QaIK+9t
ynVXSAvq5XO7utFSH+Sv5Mtp7txsijobYfyLsMzk5Nb4bzfZD3rykewSFCbpBc8OeGj0VWVBrqk8
6Q5IGyKUs6cnM1J8hoeGC7dYoDtmMQ2NRWW8hybYL5IiNCnTjE0b/IuIswF1JtT88bKYbvGnU4X2
ubaOeTrBPPB97b/JkrKpLYCgKJUWkF/CrnQRje4GrykriXFwWaMdzkL0Fn5haWW3ePIDF766/s0U
FYx7qxAyj+mEZF88u9mt8LZxWRWTftcXvSKd9nWwP9uj+95uVsQGM4c1ZbZH8cEb/joPpS6Nb8Tg
N+enVxHtBLrpau8niAfByyusbEZpHhCObgiuiPOSGq8KFB/+jB96kXnWkacE50Mr9ObtaMjKrsE+
E6QyFfrWf2x5EKMWEok3NrDoi0xsFoREou5Crz2GuWwYmQfbXVIPeHG5tY4risx39TV2rZwzyiqf
v49SI7th0Jk7GI1UwZAsExi4FIaAU4fAKxnyoXkT4ZvwolIqNtP028D4NXEG6EsUCAZT2QeCINaW
bwQzK2Qv7AEUV/BgkYpkq4GZZsjKirYlidPG7K+uCTn8bg7yE/JTaznOZIVa+vn6QmjGWbVfh0Do
6EQ9qAHoQbbiHKX5M/X2yCnoWay/hKcNjj+LqbxKQRsxT/mh64Zv0jrZhKDwtQgg+tfnnaEMyERJ
FgFipthHs/KCb7fhi6ri7plGOkvc+r4uhz/HAYqnZfHAU6tAmEKe68656P5YK8vfIIIG2n1LCzkv
KJf1s+x9zWlfqwFoXxkTcMbriSIVxKQsJ8tj35PhKb3jrlxBVfwC3dbKs+wp+DUxl3mVc5GvkeU1
vSp7Eebwou7Z7BYILu32Q/tfY+wzLhoG8aW8xoiOCbNuUOV49Ulc/RtfdZSNSuYD5vAvJEKdBi/i
dlE4KqS6P4xSMHaq0Ip0sPmsjGLMFiWq0Lo5rWLHVkf9Th715Fkij3KLUx/qnW3+3uD0B3e2GGGh
Q9Z/bTVX667xc3K6ERAZjYqtHah/55NNLTIo/ezDYUBjaZF+0Gloxtf7Ep+F1iWW9wy8eCHFX9RZ
6Rtht39P2VL2++1ziOre+DrplT+6Jl4/BnhlaHFhc0L+qBPzl+qsmFsUA2fo7V4dPiI/q7b5Kt3V
+ZF4Bf6aI8Vzin9KqruiljTGieR6b6f7czBU/rz4QZGDk7S5uqKFaEjR7cs3ORa3rxKS4AUR3Wd+
CojmONqM7APPcq69G22knJ46PV5UKC9P+wcmp1Q2TuRU5Rz8vymHBLBdlutNaDQiitFClv8BThRF
zuRwsISU+mEyAJ6K9QmD+Y+jUt1P8udNo/kZpXZFGkH+DPXWYEAFzeRf4FPSQcz1Q/i19h2u83Sn
GkHOWHK+rqk7fZUOq1fiCK+5K/kEkMYeS7IAIfpTLJ9POzbdVRbjvIW+jK85kCfs9bavsP7dBNym
Qy5dwRqZhSHX0imALWbd2sGzFbghvhYe00blD12HwvgE3j8ZinumgCTyxTwM20DmsPB2xLwEbFRc
No2QiMu/rT8l7hCw/sekgPjh9LpgPx5DG41SIpSMQBM+Nid+WV5vUZfKLhZmRHeWsq2vqNFjtE5e
No/0NvkASdoJAhs/bz3/L+9KjLZya5ggAqOWRh+ONGwGBczyzQ+/Vaq7+p1XIcIQiSVQTAjlUJfq
Iy8eJZN7+UdMuBxmPOpBzUuHTdwN6r+LG685EdRMe5kxGwtCMLfB9y+4ZkSB0ohn8NZt/cNU9B6g
G0a9Aed03R0DaX4Pc3qTpQe83jMFubn9LH0U9LLsWCzae5PAdLCWW5KDBGN7H/+r924o9v+Z2qok
8UZcRAEHPqUp6AoR4O6mwT6AC+ShIy9WY24yCWsMxBatSnQ8fm331wbmzv11Z25X3eJJ2LYvppC3
6AglQHil3DjnAKp+zC+9a6otaPrXmLWP/0gA8dKYEj5E0xXuQ8mCZq+/BAJ5XTnIX/xVlS/jtMQp
oTiZI6f17KZJaDRWrm/OStSV7Tp2rBBwZZooyqjv1fqdkb9oHVL5Ob5CWaonCYjrg5QDxFFSRAhN
nHa/+C5btrcnF1B/+VBFqQ6KTJuw/M9kQitbZ8hvBds+Rql1d0CzV5zg4B2w9b3ZI4W0HBE6oIbn
vxlFik0TV2+eLR5FJ4rzp0cJM+esWjoGRDrllx8jUaZfo6mxGik1aftInAUfgInoYIdfNNxDZPgc
e/eRn8FWw7r25NSTJruEWTk027xweOOLHVQuvSFPlR5ug4KlTIuczY/NTvzrerM7OIjVegEao1Nx
3FbAoQp18WLXLBTHQ1hrUlaoRaZFLoG9TNgj4mREJGQgFCKeoFGVIwIIUeT06lkrQHoLkYtUoZxF
jO+hYf0bRmzOpq2jzg/qjtAbJwFpDuUUqVVB3VRGxV8tFQh6LEwxTMVfsaTT47jEN7sS2pZVWwq0
t3ZgA9Hdl8JR+PDRF3IS17RQp7rnzYQCMhcZBuqwevoYFz5NhL4ELT5TdGFGzSFkJ4kLA54duU50
fg8FJKWPuJXZa7DjmR+mkKkKAWa9QQc07oB5tx1cSRQ4/OZ/SZZ5AqR7SNt6zqOAETe4tnUloZij
UoPF8pjO5oY11CNOFuKag0j1gozBm+lv0ajCaAohLM+WgL7QzkJIfpqchtYDTEb82KXSR5iLqx7Y
EsN9IY0NtsumuikHVOtc5ffecWQcXZYHovFhqhdd7K6f/y5lmrT3KOgVACIKZbfJo06gT7PdOyR/
0Z4lmpj3YoYgGYtY+ERCoIBwJ9saVuXBFsHKbXcxpIKmWALUExRO5QyCRJdbkeaeWDRRexyOHLqc
2RlDaTURf4mNA0I0UJatV9UWUcLMoBVaGa0y/GMWxTwiCmc5RYr5o1lqge9YHjxFgVAoAIH+4kmb
8K05n4kCAumnMY2j+2mNYiavqw8UYa245YKRpq2JJbWu1/TCTMCCF83CrDD+yQpZS4NbigcklXsu
MVWp3m/f3cXcMVzwnuhVDv5oz7V3G5IoHFXeE/BCTSmOvNnsOq4VSW2oWxUzb/KNyuRZ3wbZqqaa
wmOUHSIXEgMCJRBe372n3KbnWfcrYxM33Kl8YdPSSUhSa9EtYSi/pLKYBI3r2+OUB9UgZoEiVcVY
gW2vCWJaF/D3HXBfy5wVQivW/yxttslLQhk3lptLdUZustmojAWb19Egazoi8spNGwY8fugX3INh
t0QGNrYH9xXry6D47sfLkV0pZq2aQA0BQoTNoGsVb3f2BMpqqYiclJre2yMA8/csjyzoJJF1OLUh
6FRnnpfr0Am1XtYvj6eRsjCW0ma6lz1PoGgl33/Zo3PYwQP9xiMmb44cvVCG4DYNMa44vDAw9Pwx
VNz2qhtgbKsRJxXAPQhjdrXix8fyxJ1JA0hpuQ1IhEbC73aSizlXUDJsYb5N8cVsJnSe3YwLt3Pu
0WJXODxc37QL/5Nvyl+5aWq+9Mg52D3pLZ1YQFMIF0yacUzzZ2FNB4pKRn156DpEX6lKP4YlS0L/
sR0h6GW288BSHyUzm40tZXIV91XXumyQr59xeM/pd2KUzBos+zzWbxo8NlSOk1/xLrs147U7mn3V
V9KSVMPbOMJbx+7pkk/oTKg+G0VXxheqgOkVLKMJdhgfwwzdApJ/VtvLKF9zNuI0OdhEOL0Mz4/h
PHdYRKDPFCXEvdC3bmfK+W5/lCZNtTNAAx5sj2uHmFs0LQNAC/BeAJ9EfzHoDM2sLGroV/kVpEmt
T+eTvmWqx6wNJ35DvOl4U9CBeAH+04hCPkk2FTCmznyYArUsAEa9Jqcx2C2TCOOlRKmJ/yUTyXoP
QsaDc+vuKtBvKvweelueTCVLBn+Jhi7MaY5/Tu6NrCd0xU80IUw47ID5VozvtDyp8rldxYVyZpGW
8dMa8a7PXDWU5jW+VaYJuhLtt0Dno/vrhPXyfpy6cqXgnsqwRHBrFQ3JHlrzsblXIB+lOVAslMNR
D/c/t0gIhUt3o2TcidltxRm5qNU8qfJ2BaGnJJnWyTG1295I8zY4n5fMn/Sy0JGELS56ofVir4wJ
5RiJwKztdNncVNp9NkPoL/DlnqOYC6cZjQBYsuJgCTi/ywaGikPjDuEz1N/fL2CRavWcTxPutMRm
m0bukkO3sTO+emZNLHUSfenE+CMtwYj8D6yHsh/EVQz9wOeyR8QAaG4ORicXajMjlb9++iiDpEyD
D9pj1/EkG2SmM0gxJPOTU24cTh079bDxZLwmiCMGZuNwCe7E0FkvsPJ4O741tzUgQoKWXREqstYh
BOcvDurL2YfRnRZy4FH2bFq91z5Xelgd9wHC20HVmIv9gLtwEb4xTixbwRuOyrcT0Cr1MclTH+Se
2CBfThktZc2t5WaNEO0huDxypFjaieOQ9m7qs+iztLKR2qsBKa3zj95SMk8QUiwccEoVpq0WQHRM
JFJzkCfEFDDuwPprfEhkox6mP+J+q7RTW8ch/FkMfH+YshXf48hV91WnvhY9KI6udV+vbAIEUIMb
1X3IKHiJ0KbXnfHKmXwmExNSnn+BrTMXVvLGPq1r6fY30714FGtDr5dytV78biidLysokxLmw9ew
TXJv201pKogkQu9LGxu11Q/TR/DokQNlCMjjmEaYiNz8SuqCs83D1il9/xu1idC/oL5IbRvtP9vF
/b0zsfe5C4Oe4slkgsMpVBBgJd4YIogDxKEH0IKBz0vf8aqp7oxlVSL2w+yy2Xvf0TX5ovqo5oRF
52HNiUKvy8PoooOvIdvy3/yyZnFGhFiJasFhBG8+iUsgitNeUdb15wCBuyIEnMs10OnUei8hc8+k
G+Y+Ww6uvXbsHJZqIjSEP8JhDwoqEVMeRgAUM0LbAo+11kbIAZIL5fJTkGP8vBNAniUUpScIRrGk
E5JbOiZRAYNVLw6zLZwcWfiwwyodotFr8rBarD7FyQGz5csCvvYGNkW/TXPYtu2Oia4GP4hC5GDs
H4VCSsdbCQms7KprbfASpiZgg5GITOLUHNEXGi5X3BOva7W4rYhqmZ40loZ959GOwc2fh6gwtV9r
gFiwSsMK3n0GeN7svLRzED1c5VfJZSANmcwctH6M6soTjnjKijJDWeAjqzW+36nH60Fo20MCdNkp
UDhxONBhxg/NNU944+I/PPSZqYZwHV1ss68ojKRysFaVA0CtZhLDZwIFo/0Gl9zy2ADWtf3RkST1
R2deROYmIwrgThQi+ooGcfFESIoMqz9s0lYE5yhoSC3x0JhsI33jAuMskf1S1qluZBlJo3bJcGm0
TKTfDz1OhkfLWL4Mxk4udMWx0EuSNy0V3Mx48thgLmcC/F43r1cMdFJjxzk6tb/lYsbnZRuAIWSW
nLQq/fxQ6gr+gffUVKyPWG/5XldzpJ/cxpgKOIhJGN4r1ScI2oYzpF4Boz3QNeQozfiY6iixw96J
QLUHp+6jIDBJP4SzjLPTn/07ivSOZheuJWtK9jZvgUaD5RokUe6OUw2J9/26Gu6Zp/Vnsb+Iz2dI
M8oMUR6tNn4qi5WKM5lnePkbaC0ey/0l+7r7Lv40Gipa0vAmyAgvbzG5Dgki69BT0Iqq7DC3MkcK
0/DO9MlgXkzXbKH+a0dLIaxltiqDSJphRy+2GTwYOtSHBbdnsD+0Q1RyCwxymVDCjmpC7vizys6T
PJlWyUaVMGZXbe8lbn0tP+IaX6zvxC2DI/cUMfIgW7czPjuCMypd2tylY3fidJDc4m6n9LfyVsbU
wUv7JAgCDQ1+xRqN8K20IlK8Vl/TURXpCjE+SFE9tKakALsBqW103dYmFfi2CRBe1pYOHDuOgbWS
qascczkpPHjhhkM6GDm1EhqR6BRMLNzkKzAulmf2zKTtCLg4v9FworF/0FwFoQWTLIGH+our/mK8
CZ68WXAcoikRohspLR2wuzj50G0/GLOx45cwha0/ir8j3T9aeuUizxRP4lhmkttTNtHKGwQiHKTG
xcgs2aiWL+XgE4cX9e7/zQdquylnVAOYIBNi+zeOG1GaKlTyB5bx8qWkFSC/I0GO6JyPONEZhkdt
2mSeXhfBXqaTLUQBWuOCZqefEU/W92fwKHeiSlR9jI2Y6zUzgw+Yik10z5ypHc3ZzQTMQgHXJgCF
T7bc1xG78DLr5aJgW/YQPEoITNgetHzsgUVyK3E6PIxE76VesQCyMZGOr+kulU4ElmoT65pE0bCT
hags1p4zSp+ShsSEA//LRWf4fIgfJthpYOdnA8vKicCWzOZ3Tqo4jTKml6JtynJ2d2Omf2659m2I
vaeAFWyGINAVduWWXGN33pVPID2VeTwVxYd1HJZO9EtCpR3t8TopFj2+Q86byz0R+Vo9Kh/v1Q7m
d2TZ8vRuQi8ExgL60Z36hvWEMsbyvwi2gyr1r6sCvCX+c8gol7aYDAcuX+KqrH5FQOfMvX5cT99z
zc2vCNFNAsCGZcclqgYCbeX4H3/lmZ0yy7+mrc3q+93zkrj64M3uIuIDXa20NOAR52W5MP91dF9L
9b4TBjTzsrq6q1tosYkTxGIJaSEA6x/60mahu0vAdECFySMo09DsCysvz4+ngKKqP7w1WqJyAEQ9
R7gWbNnRpgaoFonZgEavMIBD0LWoj+4d6j3B3psojAhpoWjicR3h3M942hwBHrTtjraTbN6HACPO
9gkzXaCZMAjCRSijMUK1SUtMw3BPWRwo8HdOkb1236N4Qkj4IuvzYJz3njzCWrSKimpZpJBLvp4i
oLZ2t3A7JEOpNyvZOptcjBNYHrLDt59RcMa9yfH0MqcIcHYUjM2tr9En6wpQDLVd1nxhcYCO5BYe
eal5XwdHpWQc6KJUjlqKU67033HZ1eJ1QEv7OYo9BMEvgBrygoFzTJhZ/8fsJ2B3LUK2cI/DE1Xl
ppjPHixlGOhBm7NKk0hdRzaZibnIqHUHM8vXn08ibYSlVAp1iMZLkyOf5QsQbgXZ5kVC3JZ3HVZs
8tZlJOM/g39arRG+gvc0CIPb/rcuxI44xKGHGCNoXDgR8drwfaes+pNZPncPSKnVHzEW/88i2kgF
V9h/6/TcFLc3I04Hky5HlQHK2o+6/iDQ6F/hJDCuyUtpi0XD54TJSqnoJPrmKsaMM6aLMMJbsK7a
uko9XaT4wPNwsFpcJTJFFFJ4SWICmFxyG0qQ+I2pk0FnPEEzNiYeuj7nY2sAoVFO1JBnpgjruyfU
U0+wpmY75AkCFRSwNSRST8gVlVZnFgdLXCKOYMRsJ4hx/GjJJoqtfHyXFKV88ETz0t7/QVVUgTiu
Gum6eVfI3HRc/5OVePS8dkb0BvPYK732kGsnpj+P/CSpBItjUVtBkqgZJ1Ou2HtR4f4OE0Ks5kE7
Y7ii9EVsRah93aMlJ2+k7IpaFcYxMX5pwocfCA7cCD85XpKpgQo/y36vRrYAlREpSgz1A2BfThoo
mo5HYouF19WW7p06B0uykaSTUA8VqGbXfbN+yDwgE6jILtoWBxupUe9nUPpHfvBAzrdrlKwIJ7/o
9FU1jHZdvcSFreXGju/Vfl5Ryj196Yo+ftH3KKHuRqxJFyiQeA9mW+oEq648y6sFBdohbT4hkoi1
rSTKK1DHOw175cWo3FAEOrjYz4bjpWJUZXurfp+g3tRDaJdbEn/JSZe+VjCgJuIDTgJl78JgUdre
wIQpkufvTsEWtHR4vGift0K3vbcoWuMz2IiN4K9QqIIu6M3IBHlC4bimqWAzl703MJ77jAblEgel
Lw69zOXTxU6cJ+9SwoNkv6nGslRYYId9/mpV/8Ksr4AplKZwosOr/8+/XFM1PqzYJRdZb99SMECu
yggunHvjoUd/9xqBouqgQzlleyM/x7M1Qe8tGC/W7i7c9MvSf8PWxv+8BwyySVlAlCMFyndzPElH
YoOIOAuG8sXXlW2QfFt3raP8F/zkoMILnq6oHOCXKv/hoiqhKbsefqU7cAo/Sx4Valuun9kkbd94
mXBHnup54oBzq0V323QhuQCsILkpmmAazAZAKybfzaFnQoWAb0KyMxhQ66T2G3Zsy6kYuOGD6qKj
Fb4DPHuksYjDCjLYO9nyadWLD0z3RBp3GGQ3kMDflalItAlz9NKh5ioHlWM5SZyZgI6dg1UeatUE
sT9AtFmwi+hTFnJcSljLdPH4z+wXVb4wOHIuK+3ZxdMvKwK5jeEEGs4V5XLqZ7K+A1+99CgyC1mx
OZx49uvdXK0RPJgSLCqLEtQn7DbY9dQQkAIKAHVmM5NeIQLbGwV4LefKXwEsLQkReV0unaB8CWyP
LBOrrvMWmYGW12l9SyrljT8fd4u+I7CSs0Hv5JZ2YhgYudlPmgmU2rxTShbyfF1AgxCP4Lo1yxpU
315Yvq2xx4DsBlh9g0dicJs+BxYF7YkZsUiZ6UJh13cir40EZGhTGbmaWzs5p1FfCURrzj4YCoeS
VgUQIBXIORS8mNPxAw5r3RDTRDuVy84U/SZh2zEc0M7GgokBonwbfAXc4T/+1yPECjlQXspXhmky
v7RGwnHgXpjkp6hKUg5ElwK+DYIer62efGhm6b7JvRiaJ2W+TNjixnykmssNCcmd3GjIF4/R6s35
YVYHV4naf8m6WPmm+cTjne3b4UeuRhSyDqZupb6koavqX2rRaBlbHy4guWBCWIp7EoRtjZjSpqtM
i4rigHOwhvMZB2HBBFfqY7HipD/eVKOrlP7j2KKkOWcDEE7DjDvxJ8KPnjHw4eCFyr37SL6s0Swp
Xl5VQc4KgaI0Sdc0VS7x8Nu981aSYEQX2JWq6KEe1mvdywMzZp0e9mW9F3IiyxHHOvGaY5Fey7qW
Fns9/GYV/O8Q5JbGdm0jSxaD18YBsexiy6tL5gIPYtXiLyhAEV2nM4MGJeEGRh9hQuvcXNVuqP3n
VGBnVtsuRfs9wPfAlpJeSdUMqJTPzfPkwZY0s9AirvNicbDN7xfqp8IMCe30f4M/hZXFelaNa/DB
YJFS7P/yI0dtbf99nQHhMPCgiENaobEIoCeYq4tkVbXNNv8TC5hJTAPlqZohS9Ao6U7zgFPv/eDD
LXdl3T2sy+LtoqkkYLh1oQkk5Ps8xsuIIUxHUBd3G1xQO8uURMsRdbedrgYVDqwx2L+eZhOO/zMF
20s1Yt0uJn9Q/V3Bkwj6oFeDk01qVbbEAT5p7r1/nwHiYK/yr1LlsrIhXhk2RNFQkOcjnO0g9KVm
esxokB3yTUEKiO1q8xtRlYu2IjwenrJ5v1/87stjlYMIq4hWL7PJgFC4BcRTuBDFG5XXQPZSyeBh
y8TTZ7uzIuOCdDmmt6/K6qN1FOSqs4sT3Eozsx6mctxeuxpouVRY7MpmXzwsKemarRHPEmbNd/XG
46hGDyNNjdSE6oWPxLbUvTIw9rIUQTSV/RFVOdOfr3cFC1XyBrhGHIHtjq363nH+JCKwnNm0/f28
tCQ6gqo9vCCovmH0sLeU2Q3DhPDNL55mOxr/PkIRllIolfWj11CzhcUGgVWJJuzzYgOz1ZPicXgR
9bHArEgikgXIK4xWBCZMHYfFawSYL9A+Qp+t37JQ8Q+ThqndnXg+biCPbQRIRqn94aGRkLgUG1P9
W8V7pk4s9eKgtaZkKJ4oYDmGjD1kgR8DthAnC/V6r5ZSXNN4xDWpM+MkWmeVS1PxDf7elKrhO7bV
lrfuKtSeG3GKmUKEdugOO3dZgM5X6qdGOVakV39D8o/eC5uxDH4kkVepB2sZHRQosSvrreJJM8Tz
U8iqUqAfi+xuYHMd9A7sD5b2U5aBx9x5q7u6es0C3giTWdBUafldc3SV/21fadYY0oQzGVAahet0
adfTNEGTSOGPtxYTYftxYQ9sD+0oPGNGc/vkRfPHdwpy5kDjHuNDM1BIoqiSFeSzqF5c0oqwjKcH
PPsDushEc6oQON95qfHV9S5DWV3HBlVZOmRzQ9UJ31RJT+ZKW9yhDpkpx7NYTo1JVqdQh7HNTi+A
lpLcEx8sftOZM2VhF8Zehto3GXZw3Qkk6glzOPB4nqkXS0nLRdbC9G7kfWsK4ISwgrmGn/7GDdHM
aznltLS/xx2nFJbzTXr3B9fPaJUle7d1mPxdyII+n8gqi0HTO24tWdT8euI/9lBx7DhW/erkySD0
dmDl+3TcCREKf55pjaheO0434WxjlfgPpCtgIElbEojM4kNKP+F/FYQ7hUVOEgveyAytS7Vc1jFc
8k40sSILtwbH1ekr9ShYajpHdx7GknbxxTO0dvDlYIAZa3ANSJsAh2I3pmdl9D9rWvCJgQCxMepb
Uh5WmXJeZI2Qj0nugUB5wQVr+qS42ZGHW/ajoRynsSqLOEGL7AMNi08gbxdD1SB6+5V9pFIZ4Eze
VohENE6kyyC2RV0MFj2oPZPQcR6dpExx9AMVCrxFeYvf6DjF2MDWh19HCipRfk/PpfFHlt+7RwLd
Ya8zjUb6P2Ac3qZjyGlVJwM9+9hBfrNiR/zIeX3ZdrbWPVtNbzmkN03OX2xNtWXb/RhQ+gPc7CD6
kemxKXG+p7hnehj6IY+2SK3dCNIQ78h42PxtXRWFJefsUpShVtH8URCY4tSh5DFE77nVI5wWSjz2
vJGFfcaPjZ46wCZ70DQU4iSzPeQxaw7OP3IsxqqYJmM3uVRTGIO6MX/+eUt674jOUpGy8EYQVW6g
KsHvi6KIOv0OjN14CrJLghgfH7Rj8b4v4SMP1wvg6Vpk4zTMBsNH6BG6D6KECucVlJx6jpG2+SjZ
dOOW8zwP9NwjFOzy5tjSrcufv+bzh3VtXTQ0CHK2h4OeDcvCXNkMSuCEBv40NTdxkqotWtZuDJkj
d3sfAHd89sCMdfm8vXQfIv2JIP8CLKKphkpWC6hVFaxVzQCLmcbSN85O+RhdEAmyY8FFKNoarZ56
OQksEHSwWcdub4IG1PvJy6oUJRTH3l/tVu1po1R0fdbiH5jWiotIoCjIDsgRkOe4p9kU45mpKveM
XXq7XSNsylR+3b417/FG5P7wC+Niv8KiudDHiIQvj3lk9dpAw7eXKFSTVQBHR6GFthy8giE7WqP7
8sR0xl8n36rYpUtid0oFyK0D/UGy5/kgnrdXRPqU+79pLN+zbn+HqkGO/Z2N+34Obv5HVIezUHgC
NwWH4wtoUDJCfPXeEJjpfkoiyGoXgaQmdvRVuhNnGRAz4FmtU9HP4Q2Yv0JGoYDk53M58vRMWm1+
JBiMIIXPw70K8MU95mgacYzGbeevc9J7B2JPdU92Tfc5RNuqCUASUu6o63VaB1mOy2EzX0oUzMvf
tCxyRLcrkn8LI4SJ+MQi7W6QntzVtDORi97pkawUf6JPBb2jz6/j+wAOaduxXJ/LqzW4vfJPyxjq
GAQoXau8aphKUAhadRMWNdX2WQBVinoNcQzbJFcQHOVZ/+GV7pgqZ0NvsFXyPuq7dVmTPKfE0s+a
Ui1E/7Slw5qyf08hnKmq+iHoGwNvAb7VKL7i/kCOi90klWfrc+I6LBsVtS5xMZJcWMJ6Hy9bwGvx
kwuOO1NG9+GvU+r3FXmkUodM4XEwR/uyymMUaGSQrns2bFOzvHi038duSp/C2dbHGPrT6YeXIiSq
L1fGV8LlGov8A7pn9uiISPT6mRpvW7tmShLwLV2Bt3GlBu0C7GpgfAGEAD93U8Ovhq3m+C71sUR6
Q8a3vZPI/DLMiJgrRdjsSs5hcxSsKjsZwruHkUeCu3paJxVkKKn8tb4Dqf1qucB0cwKNwl7PWGiQ
V4qUVqcwjT2Fs+lj+vjkBogLTepqRijNqgLs4UPCLhrQ1twxPa9l7XqUOjqEg8ZqHPv8MNaV0HVo
xYU5CLKfzc1pP/Gl3MkBKk+cSPeBJW0TsyKG1nBHs16dD8yfZ8RusQ9nU0bm+9wbLiFvxzqCBT7v
ApoCBdSBhepK+hLWoQ/ealotgPv0QuYLyxFS8Y6IB1vJLirdFGv3sokyv4fu45zzV/nx3UiwPaAs
ZLiWdQ84zB3aDG5t84NpBxewYMZiUJkNklBvx6flDIz15OmqFlEvLMzQ5UDhVsfaZB6X5gbQfXZe
0PCgIeyCzlGl9zuph5O5MRarI8MH++j7ihnO71ivhakLA9cEocMec4zxLvZJwldZBrmL7K4MClKV
Be29Go6TX1/EQdRaeJt+8tgCIwe6aeue4LL+E5NR/f6f0c0EaZMtMb2RmGdEz3RVxY6llQDXN95L
JxwMB1BWY76V/mtOWmk4wWPTZ46jkbYb5IG2mxmIkPmhQsd7SZCTRvh2i2vaNNJhjUejl9cM4Xbc
bdVRf332IvI2q+88VvJNNsDvGcQjfTnASsPB7qkWXn6H3wKvoRuy0fj+7dACumVWpRq+ohqGAytf
pnl3ynItn7L38xVXqciJxqbWWJCCy8G48J4LRUYDtoEuWeqUu6mL174275aPDCPa2p43UplZLkjI
ytuTjLLmfoAha4t6GhsSgHXhxcCfmDGPvdVH/oFY1fk+F9Xfg+KooWYZ5eSbx78bDorLaTPmOP1c
DwMeQArJcIlxKiIXf2tJ1hWuPB3ItMxIayhUNx8tacbStfIB6uFpccVTyY7n4ymO9j69CAZYF0ff
VPplEvTqrmgEi0VF851KuGt7pH7ZwcJoRZGd/1OrZISdGyMjkN04/bii7s5Vd5i7XvtZG1Effipf
J6BFx1RqyTqqwLttcDydFwEvtLUGC6zry6i2Uh8Ut9D/TKGRdhg6Dt98FgH/npaiqdi3ni2fLklX
xDGQg20nvQ6GVLHWuNw6sOY+gFdsCAZS/5FiVRdxNMK9uKp6z91vjK2oUqIfhoKVz4DmrQF1iRYb
wsVg7RCHNRY2Wzl/73AAUg9lryyl+PsftWQ99r9/9VtYz7Cm7PflpoBd8/KvqLs2DtRIN3MYGeou
bG7MpHAsKSHlEWFaIdTApi8VmsjNR1L1SP7KamH8RnsC2HfHS1+tHYy6fYvMY6X9TKdsU7vt+n9e
4qYP3dJU6MD8Wlr6WI906V5vfL2yK/MtcbQUjhsUQMsA3H6HlNGib53yW1S26cMlCy3Im36esU2t
LhWEKqf8ccBZfEGbMfDDIwkfO3mIyKbG6AqTTutzXurL/nWcGhsac0esv+0OIVzgl6Vp3+EHCqm4
Tm1aD+hXu+QNHXUPiBTAU43Z451tUgs8L70/tlwwsR+hWeY4CaYQCJtLZl/309eXmEhFh1q3Da6L
Xzp5Dn1Nqcmw8ER6yPXo2kwAXCAi+f+4gruAbB+YWoEcCh3b/GIHH4kKEXr9zMnQn/BDdeQ+a+Wd
sO2lWPnSf9zf2Y4+5p6ZllsRPw9SjeYJHhswFEXUgBCrGUgQ/IvHhrvcWLe8dmmTIUP9zX3B5mQf
kMyLZBMNHJZudftIliIbnT2+550XTi0C/KpiSw4il+9lmND3hO96b8+XxlZvKwjBd7nsLmeqCQfY
dxCiN/tFhGuguyuBJQ+VFKknTLUTroMYfw4h1tQMeWqcmPdV5lIPMnndYV+qFoUS6yiyJehAStj1
tm30A4uQ4dcHDxX1oKgHkr/pLeRLDXd5bhW37T2J/0FR9B969y8ILET9PqO/XeOzdzjZ2yyoRnx6
cctyWr96j9wRSygz817p8Tku5gtRe0Lq1Pz1dizO9wK9XgZNi4kf+zNzyKN+FPV6i178OvG2VF8t
rjLKUncljv9ZWhX31pfUCndnZY/fu7kfqdVb9HUZJXQZ4zcuWaqWcQ6v/bD4aI+MpHh+iyRExm2I
CnkYSw1WkDZBhyoJZFLjZDUdyuljUR/1mSww6MU8iEKoULaA98Tqkebtfh5zSaprHEQ+T7kM00xJ
wpeQxk49DDGJHKnyV5QT64QrMRYa8x53zidYfugOdj4nCrLb+8WO7hTFNf7Z2/xMZc8nD1jZX4Xv
cg++JMyXX/vhoMylMOoOd7K8Pg2Co1QMK8vxVsTgMAgNu9t9XTQpRfb9OgDr9wb3aIu/WUeuEpEH
sJHi16enRLLQxPGek8wVZUCPF68uPv9CyC5ljnhylKPjaijiZ1ENcbgyLKwtKSOgazdLlqYa3eAs
JfQa9KBj7RucgO7gzMe1ZytOHtsog3vZXOhHScJLDBR3AIy4Us7wsQP/w0C+IZWef3hHDpzQVrac
Zl3Dl6ePP5jYRCkqnTgz+DiKEbFiFZtQQOd4X5d9cONi0QUMi0FHr5rOdXPHXC4HteHmAfnddp7D
gWLBH7M+jWd710lcghAfM105NopKrlZK/6lq+aIXcdZJNP9WJCfxoIgy3V16Hp9iso3ELcjVEYtp
vVOIxZoGiHeXa3lj176aqtp4d/UiYj/CCDG+UuLDhlvCsYmb9dKepmL/d3wZKvv4YwHAbO2+AahR
XTqm6i4zXm7x73fq8lBghMUKV1pACH05ZpOZTShU1lwoaXK6DfK8wJi8XHxLbVW/bvzhhVVgfaAV
hrQokA223enNy3cDeAhTkARnT+2omKXNgtRuJA8A/C139D9uf0qVYNitcmB45jdxPLZ9asQFfRLd
y9kI8sFzblMpd2f+rwf1zxvjB9+rhsI6SXyq0tHaaRE25GmcuTY/WKzvSQ5wqV16jbcsV7pniix3
tOuCKwKxmQYGwzNABRrKT/M5UvZuDa2PpeVFuB8bsIoKLbOw5uFHO+o7zXP5i87n9eyUCeZefAao
iHW3pmxdGU4Ke7FxkgzzFoi3Kw09JjA/Ugm6LmG+JsrtSLoAo98165GbHV8DjVdvyCIZJfiI/4ea
5ZWPe1tNBbQhrDlvAfPT/ZFudGM+AWyd39oBIBVPQB6CDjd/TWp5UftgDNNffJ8l9wFiMSBIDnOa
4fm6p9tH4gxuFUVnh+aO34G3GsZsRSgtNJWSibydyzUSUW58HVL4RHoaHusHCBJyAlNUwvlmVKVd
hQWy8vJ3+2UyiY/ruDDIUUJUyZHWQQ/5KLz+txtDx4b0/zq53/IUDtxn0JRijhZZoBFI8CoyWz8W
F63WOU4SQRgMMbJpxKQqgIoWL4Dpdh26DKA5fcBVvDTDF2vxCxkS4XFLGkl7ED3p2Bi7wpO65kJk
By+bUKfZUbdJTxoejmjtHp683CmS616PR+Rnl2ZzZzyI0ZQlrSYRUZIUGJxMu4PgmTovCO1P3FLW
tScFxP23j05bFmj+XXU1Mor3YZJFUoe0WRlDCrg4epd7wDqjH4bNTg4J4VSdzgNKHgWgPae0q0Ck
hbG2FDpWqfppE6W0E2wZk4SP19fVTN+nLLIlEph36+xw2/NNgwypQ5c1jrCxCfXJIWbtHD3grr8T
64CXwjZu8e4sBrY1y7qYoBrPppnxMwuif7TVOZjDVczKUh7e/6WeSDWphX48xZacc7jXNW16r946
vVoHP/HwhXrfIYDO6cH9seanWEm4wHZ2CyCcX2WH2Vb79R1RFORxMdxfqxEWT5ZfPeaQht09zP8a
9SnLM2E4UBqx+zEgIpFF5dOaRgqmx5h0zzIqM7QJKRtgn45GrZnYHi22uVnT/gQnDTVg3qXB1I5y
iKQhmFoHhLVrAh9Qvgyhxeo52rsCw7UpmH4jjTPGKZgXQGx00SmuHucK1pYLIo52XjKy2f6e+m8B
P1f2bzQQpaPcVE1I7N+4hxaKzMovspW4T0PnC0X4FI5YoTkAF2rKauxU+DMAS6iPDbuSbWQhdTDO
T0QEtn1/lFF2/oI/urVJfWkOw8hUGukVg27kW0cWZOk4feiKEOKMZKl8nERdkNE3UrvOjlCLDuVW
haBij3lx6af/80gdqIiw0V+wHM54TLqbMMIVz6sLOYl9JGA70D32bO6EpkcATfK/3IiZlnSgXUBz
pEiyw1gsOnAIcCNAVHv3whPtxcx0KQnRJftcYE+s0ayWHg7NvgXJOywB6iWBI9/WVqZ9ckVVulXZ
PlnIK00CrbuvK+JL4ox1JfOUaD+Tr98qTsiVf1e9LkQPBGD+1wSIDgop8H9Qt0SSEtQQYpZtZSjE
3YfBChbnieBy0WZYArpApRKPCCYohByC6f4F2750lUiXWDnC1vNt+urcmm/swGBlKBbbQrXaDP76
TVkkl/hQuvl0X0evnI2ZLsp3tUX7Y+Ikdri0wRX4e/gNtVh+4hy0KPqeAAWeWHN8IqVjZpHYuqAz
kTA3VcBw+3v8cR7RNViBb3ig/6/aXUu46XePfImAbfYnEtLCC+74DmevK3cZZhdFOWFp999l/mgA
DGxWDO6iMUGtcXZmp93S6pa/f3mAiFHdEC8Qj4bA42KFoDA1IEsfh+WGCuI7aI+o01Iwu0/7crbG
BPJCndhOp9PcRRfP/WbvqyTyBf67d9tid63xMxQv33RziI7ksxYhJamKRyIx6CAdLzYv9EiIL/jp
vB74xdGjUqHNcouj698lUO55iIKEwmoeA4w77Zo4I3hQF6GoHUtPQafUldMk2bvrFeOyfFqc+LLA
LoUzVlNsclA4l05xWn9bdics9u880JdHNdGxRdH79UgaKFolJ8bbuJ1VcgsQFPTBC/zw69WEGZww
kHCnBqcHBKQR6++x9VCn6KfNoK+uOCY4iddU/yyexWXZgj0R1Sh2CSE8DUbWzEkL6JrDmA7MzqfZ
Hgmn8FXLjRl0erzigIsNB5gH5KW6MrTdxsDE6l2Qw0mzinNul2CVGrc3YllTfSpttHUnjd7dLvOU
5Do2paVFOuJdjv9egERTrum0Kgvm/Nhkh54u7cMEfSQBv3ze2tNE0M3MEu6aXC8JTuhySmGnn++n
tOAB6WhO0DRF8esNx7e7nirdMVIO+uaDDWxWEwUoqvyEOa0EGg5y7cHV1Br7vuBm2hLgpc9whqoi
YoFfEzleR8JYsOdJ8/sLsUqtSgtNUZWlpP4YHIaP3dlxhv/V92cJWI6Xm/KPLVHZXPEQ2dNqpI1Z
xJGcVuBp23RZIkWhGJSjIVaDRQ/rQ4NoirDEsrt3jW4nfVinY0pwHqJdrgYTNksMamIj6B6PB3Fm
y56x77cW4gXY+xVukg12coBkf+hCL6ZlSfU2b7eku4jtKJ931TUHHSmZeq5ftChOyuxwBtT+y51q
lhAnNUf28mZzXFXFylp1DV8FGnap2zJJ7U5m5xQxkH8I8ifnSP1YEYIJZzqAQyO3NdxKifvHwSjc
Vez2YxzfP92YRzft/r1B/n9yknEpyAstTjxkRDf4qMJc6JtPADHPlSzDM1EvJWiz+xkenEdp+bGK
+Pw4HNdAEA+XJWcrKlJpM+Tefs+tmzMxdtbrMIeVUqCkotu49pgnZvDTMPvu0C96wiRyQaumkmgg
w5BF3WSZHPmT/62qYRzeyaoXl+wKX0e/h908QHjHbcmUZDpzGkz4Q0NRlFLe54/zAadtUP2ikH+z
QsWVKEeJFV/ndGghBscaHJWG8KIuA2JrVUmFZdxJP/VWyFo+YLCn+0dPAwx1oOXxa2uMudpLhvo+
SF+Y9s9Sdm3Hw5WQsFNWPtnhHj8Tfp0ltYxaVHOR1SjFxK3LzzEoGpMYVyMKRS+eYhoqDYLAxSyv
2b7kcx1Wc1WD9om3hoDrpf+QlfmGqctKy2A1Qdc1NqRercKuzmUYWRaqGRIRLWB7V3aIKPD0AM9i
tL/crphn3+WTQLKvLYdGSK/d4rBfdHSMRn2PvlKnQqgjx8Dw0SJlhXYveqxGYFL2o8ejhlivp83W
txIk7JO2T9H+/osw5lLRYq/xja6a7Pgc0mAZybnlpE/z/FEJ/mnRDOitLYs5goQ6alQNQ0vJV7hy
XSRi9aQ/JBGr40XxC1xMNmU5eWBvd4MH5KpLdO+bU6VoDZNFj21RNhaNj9Sti+wqv5/eanbTBjAE
fHodoZlkIvy/ATyhfMiq08H4LF/3zDGCGqOxOEZlIngWI8ln7fsU5NRY8p7VPoO5N8U2zhfuvTvL
5wyUCnr6QLyV3KA4/f6Addeht/jQ2r9I9uLR44DWYjbRtxXsRMAYML5gOLTRZpJHseXcOobE3e/J
YG3hx6c/J3+MX0d8CDxTXUKVvuvCmqZFbV23nbX+0l5qmE5F4ZgcGZHON+3xZnBNQUyAmMZHy6aH
Ma8y6bWD/+BWgzUP02VJIQc0NkuKOXZ2iXn5j7PyNWuy/UP7R+ff3A0tNeyXMve0P+Mr17NWZmw/
Zm6cEgoHohiwtu/hdkSKG/lRdCU8bgjl3iCvKvb07Q9il1tr+C8R5Omwb2zLTYwLuC/0rnePgr5w
6vQx0qdc5LW23calSdNHue5BCoH7q16NaGd/yuniSbMIDYthHkcRLpHvTx9rdqy4fV9ar8ciTyik
eFxPTtMPFi7fIwKL/JZYOounhBHipCa2WpC9+uj7M0poPnQdWNptVJ/ynGHwmx/My1HK2jLApeKo
A4qTlpqlr918irz0tgC1DkFEo618Xp6qniXJEl9o3FleCtor8p3TfUsZmfcZuDe6LltgkKtLfBGq
sGgJoGO2V/lhDutJxKzgYkBlTY2HSLafQua4cGc/O55ru/sxn5lLJgihO8j2GjPG8lk6kDImKix2
JBtvxvX7kNrlOBEwKC3gGp3k5x9wFR2MzceZyJJqf5gmr4F8wW8Vj0xR9B6ckibV7N5S11TTJEeG
dwswIC1e7fSirYIv+3swaPWA10WpYGq8zh10GeBatnkk9llFs5ZOQOBmYG5UY/dSmtakJcUZNjCH
hhGhKv465ZUid6ZbLA4rJgkVxFLSrX0pL9HxfU8iZeqG5PqaUpV4W9ukztTj8BP3Y/T2Ngw9EcIQ
/6YDcoxBqED8NJy2bqOjksc9z0Mpkobv68/5FYwJzfCDSZFDrb9StMB2DUooviE9fsWx2eHn5CVu
H8BRMtAO5u6bof1X3Iocb6iEI/tF6OiZXoKZv/Nuh8G/TQFrAiAuO3Bk0tvbtMnJHLYittBmJC4E
T4CUlbMBgaN79fc0PQISyt4XVNYblRJUmzGQ+xYVtoleG7WlWwy+LEpv0Dtbf2vAqRzWEb93rEG/
goTDAubzbPzhL27/raDM2BUHlChPE7XXHabOkxy+swswH/+xJacug5EbiBwLkqzbEvw9U9GyAnyM
Qktjxklq/P155ooqfpmelXkYJ95LESxh8OcUEOiFZ8mXT+yX9W7+iXPUC8e8pcfckwavlMEnAfUi
6ULRbqCosotc5eAr/vxjZC2QptUi/yyFMjl2NeK1djafYf2KzKbwkVkQlFXjEND2IeEWFxIUGSEg
27IOTwzX7vnSWP6bF126/fPdzTP1NiC9m5nrAbzBSFqXXeAvna1jeYzsRBu3Np77N6q9ylqIcA2y
CZi4Sw2U8FfJRd9a0JKWyNnrkyIF0ZQ/w/ALDKI23o9FJYK7ZIcLMtnTiFRhp329G1lisfVkbxBc
kxg456S2J/uociE4jvg02t6SZfmYu0/6IP+YjLNrJQvT1VUwLsVhghuU8BH9arn6o7VvOKRPVYyD
gWSbJj/NmL4ysuYqUbuFx9JcAdiBymD/pwffGqQeLpans2LHBimSMiMq/R25kXbLDB1g+RHguLSj
4ioioELh8crlWodNLfJgfrad7QqPlFdPpBmBluFtVUfY9dDg279d8GOH1MXCMXT4YZVxR+O+4Qv7
6O0LGCx2SkJ+rQBDF++oZ4wUz4ofutnojrJKKVFLe19NJQyWRtcKjYBs3Ua1moDo15V1t7XZzmS7
5xLMf1lnYC8vtGTfHsciSk/GfWSKu+UsmWvOZmtUnSFY7rc4GCXOfKDQyr7/bwBEVNEPpMzugEuk
WRhsaNckZRX8LXYAl0n7WFdsSLdGbsT8TToSjohYhnhA4Cti/7O8j4Y1KrLx9w55f4oFgtpDEqXQ
0XKskoabgyp5Awh041kyb4VvddFTFHr4VHkxNw20mHHtpj6EsZHAJM9Y5n4h00DrZnJKIpZWQJxS
BLjPl0drJmn6tEUvikyBxznfFzMzSTO+OA74+zquxymAwWewtmJr/qoa8/E0LUnGTzK0eEgJh3ka
7vOagL1sni6sdyDet3v5aQLuO1YPYM2M3g2E8gx84EHCsdaT3nOJmWBphJbylsuzfhSnMB5LiEt5
wFdGUCve+ekFZH96jGi/+EmkWIXKphLu/mKcBXjYYHbtkN6fcOZoReDJfgBRtskA/ZjMrXSESGws
eShUy1I2AjjKcgiM4oX87Wv3iHexa/czQYRZ8mjrvvjuy/pGRVEscqZVdNPGdQa5UTa6JmextMFf
61kQ8ZXA7YigsqdSS5T/LYOSKRZvJcET3G/nXEZZ6OgppHrhzrsptcdM2ThrRuv4tFQ4rLninWUu
5nD78JoxwYdMDRFrro+179LLN8P53o8QmLzJIgEZ7vqfKXLNyaX93rsCXdSLsQKD8OhDMrJQ6SOz
TSPcb/ursQh1y9gl9MrxSvpWtJg6e3d7jf+wJMiR97xZ4gIZSVwIvzikCN7dLfgMY3nSjqG20Km+
HFAw6Zw4wq0GpCJHSz+mqyeEdan4eZ/yQgz0D9KfMyjjfi5qM8FsAaZjk0KKex2kIk1lBqXKV5Cw
Na1a4oZiecPXBAnwBGxCP/DJAtd/dstrxE5gZH7u0qg6bW5xRRFOjRN3HjEOZZTXjNlET1GqwLFq
5I7YX8KZvdu5eHP1um6SXQLIeeoF7DXP6+08tsHBSBGtgai8xxsR+pej0pbE+NL+ER8gUwGLh2I3
QWDwE36v7dgvODX1JzVoMAo7d7x8w47bOKBQYsURWmHigW5YW8Lno/2LQ3BiDKLU2KtjYo5KbPSS
LJ4VTmmJbjIqwYWgcAKfT6Nahxq7vkLtA34VFZdpzZ7NGvy3xIzebViRJ/wUlacMGtuLopUXB0ST
Kdkg+ezmX1wG4C4gAmGQeNpWOmJWEtY45OSMuolzSQYTpyLqr1/7LPUTzexn4kyonVpoq/D0QWC2
IDdTmebmDkZ5qwNezxI2FxK6ZG/ArO2RLrRpHVkGwN4mdLgY8/IywTOy96WztkhLeNNbj+EVTSt/
GqaypUGJSg4bM6LSaaY3yHhfDiYZV5HZhwGOTiRYkO/gluqOlwXqVca6khgdXhGMIHL2bQjBWjqa
hioALjlpT/Fc0oWCVkBEPF/1oasDh1R8bPPdBY2DDO/1LQQTL0qUZgKeFFRVIwawwyYTToLb2ca0
ei1ByqId+uSiU8F0xKpAiH2WKbAcZNh7osbcBY9xlfQJps279qkwPyH4DaBtT1dVOwQiV3QZJbCT
3ttefDzk1Uf6A6eb7PEpm5wqJE6PSXs9jQFRujSfEgUlZP+VdHTRhsk8yK0lATSFXmtxNJxeePa3
fUQgHr1WyYqYu6Dlka+waw0RPeCOuGk2HIZSbqUAyvoDXnxT7YTmKYrHAb5+x0onRPfWagXA2mOr
O3FOigO8lztZSYGKSGFC5uIpBIHEz7Q8lv7krNE7KwfEBGcDT0q4qTfcS3UDb13nigK7Eqva9LV1
j7PEz/p5ERimJ1R3PtKcg0oi7Etilz+rK8jHVmvcpWAJRBQOAnpnVudboq/NK2+Ys4xbTcVtJJK0
YMSNt2qfeZcQdQ4PIcX+K3UXpX6ZYBvvY3O19hsyzycEMguy5ttXhJBnDjtv390WkJmXyXNc8xPb
SyJ+SRTfHlAhQYehH428dQHal7CEPis3lhFHIw1/cBjq9cwRmiVILJW4/5ulNVK3Pku1+caN/7Fb
nGx++11Tw8IV0RqA6g2DhBWCUwtBVUFz/nJcaBjGlPlaJdYzAHUjIvW4N0M4+VYNpUmx//V3YepI
59chSbyfBibQl3kA5X1l3bws8qlS3oRZSVaFEkBva6tEyTHwzgn1mPrc4uImUzdoVEbJMwQQUNK+
QKpMo/OjIIuRInq67l6F0aEJ7jpc4K3QrDYt4AVl+tEfp4O0sdNp0x3QnL9qvnOhDI1jRPinBv9J
gc7D2LHcOB0tElDL8f6nNvx4HObgXv5+d191vWVgMKcCnhWLpUuoRO3mfevPMwurrMoj0+qLyrto
yCU2zNM3Uw2cR/5HrsRMc77fq3MD7BKdBfRTrGZGhHG8znWDK4AVmlYl5zI2CGVcQnyJNyKh7BKz
lWo+SpejUXBkcrXBkgDqGZbxmU8tfednsrUDdsd48MdBQjPjlBh0/Z8fRbsTHRwmDd69ABeh4qdK
LkLK0J4psrKinILwlxA5Ml82Myfsz9lKBynBrUrfniAr6NC9ICVqj2VAErm/w7yLd1lSScKwo20Z
2acmteFJYsDUuwxqPAdpxawbGSWePfpCQWQT06+uKa9lFcUDOHmqYbElbmcwULSk+DEKpB6jNiYk
xcQGNM222ynqkXOicalOpTDkGt1yA87cVxJQoVGo5F4304KGeF5CuYceb2vq02w2wuDvXdC/iU4s
/dMYjndLPcm3lc2kx8OeW6gMvQPXgE+ASBQ13mMBegUI4ekenwA4gbIJhlJrlacOOPiyfLslcUep
zKQkv0Ow+0NVMAlrMsb14WbwZfjiMOcZcIUwN12Arz7jM+BZVPSihz9eLcNmejw9y90sRAjqE6od
BwE1rI74x6lR73bR3vtIjXq6eF/L2wnjgLPKgr7VcLirKhheuIZurkXyuFj0e3Do4iauHcmUFV9b
vWUz8kuwsJ67UrH2Jg81b+b8lDfMWRL3RDAuKP/vbNarKa6zK1BHiXa/zR5yWN7ef5YNiWH91ITK
vo7ZXTHKyJ4ic0WIQJz6JfQ5UNkoriZB958DuUSheV7aH6PYZg3u2OZ4K159MZFj51Bg9u5Mmv8X
GPxQSvhUf6KQ2kiKaSG5zIugRxwZFG9jlwyTbfRAw1AIeacgsqqgVNjeai8k26Odywdlw8rDd7u7
fdFhTWbJ+dgd+MfL5GFJiWcx7ihBJQRFq3elDZJpQ+duz0rp7zCrbwwdUZ22zPHjxCfqyNFNZ/s9
9EtBbyosa64DZJykrQJOunmYQEHlC/WN3R2rImKnxVCOolEqWyWygxCeK37J37kxxkPlPJ1aRcWC
AdHdhG5/tx9JLZPEEXGslfrXA9LStetHnj1ArlGTX7vcos5QcIEQYSKkoApmpXfbddbBXjziDXiS
qqzX34U+v3NmFFHDslSD1b4nIk4hcoaQtxlWI6IaQcDfCyg1YZbWhN/hYGXV/6tXWj8YA1wGb9rX
aQVZyfNlGJspRq8Ar7kV2FBxStCjUiGaSHvxVc2WTyEmsZg6KUXhhEpFqFAn9Y5AcwCVOkEIz5U1
n0LsWF/bBMp9zGkkUts+3GcKIjUuT3u8ZAkmsCdPKia7nYGZDu5Exj7Y78dGgyiO+YvV6/v7KFsw
hTsMFn6SYcAkPvEask2Yj9fJAl4Axrde7JL/s7NrcikEHkXPR16PLnH8h4VJ41zsyOMtymhQooge
OA0KQ6kkJ63QDmGG4d1obTU1kXMl+HgHnjkHH0zuXsth1yytFPu/S6gwHvCJzJsIf1/eqk2qsZQT
/p3JEl9EUYu+NwMS7oDo8wRrEk8MIAwaU7XW6eoGln9k+TwKbet4//g1K4mo6kVp2eku74g+AHrL
jTpXcVPuKbwN35oL+bMqMjob2nCoX0zyGGn7WKu5DvWJjeHBVbaK1NFdTnCy8bYrOTXFYVHzRclT
x4zjelPq2OYzyfup2UvQZDM4+loEiK3563Vsb+sz7v33QpcNob8Jd98ksmqkJbb5WiGe7W7Ej8Dp
Nj9Ugbjxq8PGwJhmlig3t36589g4t/YFKm0E3MO3OlPWe1byJUiPa3yDDQAK1FsthI9mWrJVi6qk
E/kh/fRVlxb7auG0PmkzHm22reBA3YcyPjerIjfXSvbgQUVGUMaMjjrxJuOGQykkQ3UV2NkeTdtj
IMUY5nQCohFmWL4KJnSCmkEctKwIMxXhNqVWytdeUPC4SOYrashSb8tbuAlJS3If2ufAqB3hUfBM
vxQ68wgegM9GyGWT8G1Hi0EjNczwljKjhptv7ajpj8SIug+I2vY8yFccipq6spWfOmriEfcxOWOq
2sYBDn3yQvmxYPRffLl8iPTGzYXoiAwIn1hfjyzCPbrAj1XB3SCj5aBSiwQjElyXhpSjNs4yD78r
IhC7Fs3cMCJPg04YGb0b+e/IwPAuvdMw8aEbQZDgINhTxwJyI6Sz+RxlvKj0d3BuxukjPdfKhGdC
HJYKyoarf3Dem9EhWVUim99XUwu2+JH12k/Wu1qJuEseSjjivkTlFHZBsad0tnKfJ5+Bze6P1vtc
N6oRr/AyTo6DKynCU/gES0HwwevR76IQrrB3D7JeVozwlEcQRCcy2yhSYc92kjFvJ5stqZaZtm9z
SFVNhsQbPU5hMSi7e9nAzCq76QQoxZBsl9GuPpJ8PdKLBIcZm2Hu7SJhVv938rqIy+jJodcqu3jX
xo0bMY35aSaq99GZqRyqIKcoydVS5I8ogK0MKVRdWvhPJvYRiGxm6lmPahqbmleyTxSkQ5sQb9b8
TaIXdougYLdoRbXBqZqe3670ajnivDls4Te6nCbdn5qeNihS2J+Ez11Tna+uSKQmfUzJSMoPXC/0
HMK3qXL8Su6d6pSSiYdpaCXbfSOvidD2AjKzEg2MI/FG8KZhjEJSAfcqJAb9ElIrHk8utd+C2fYW
aVFlukv4vaVnRxSchGGWuGfNizulhJK8MmP7VJqCz0iu/wKd5nn6yMy2LsQHrHiTo5wIVOjLRruI
55oJ61A/fa24va4+ZCNEYvnlcAlYmi6cq7KDtbJuEV7LAxbyUv2Z3ItsqM9AO86g7/e95c/KUEkw
h6kjFCwFnT5zqvevlnIvi0AgT8appn+DCIFvF68iloaOTYss8GFoRcFqoJiH11GT+KjefjRym18/
Cdsrc/xCKrlru/m9sWG6njfM4UzY+4mXAEGX294cusg0oomBjSjF1NC1sTN6L70KuZ0PfLkGVd67
fRKXi/Gz2RkInNmpCzCt/b7yfkmh+V7b/MNDtvPqETMSS54Z+Ho2EH8JC81PJMukHdjMT24HXwau
T/4iORjptyPvgaRah8O+IyEFTPUaPgGJK3VhQiJtIwlht6X2QocdAmMNvE/Nftz+o+bIdKtuWV7X
kow7A4dX6mlDf6UqAUh0m0HHutiT5vxlDFOJETiUhchosfFg4vhJbSeqEJ5eHha20HE4eHI5L4tt
idLGV+pqk87Ag82sU+rSBjEuG5xMMCG+m0yl9iFIxGuj8eeTEAE9e0wbGA+oHoWoV+p0bAFY/l2h
yJ0gPpCYLQVDrtklEo4+mYtNx7HINlpR5cLDQOv5fxuNMF6vBv0eF2HHwoXFEMH582j6CDaWBfRQ
cbT0lNrL4OF0/HEmmPyK5qgq1UVcvbC8ABQPcyYHzJSPtm1twYo+X/5uGosPaTwZA7qaehOlaNwZ
VCP8+ED1Xr3HupIi2+3HQNu4Qrra9Pbr+CGjxi8nVEhrl5t/Q6ABnbVE2YpYo8IUYWnGD5+Xt5DH
dZ8sDhDWna7vRYAAfkkCk6etbKAPSvOEc60Q7VVrDfFCxd+dcCbQ7EryipvUq4v/K0c8Xg55Zls+
BRQqIqQ10Ix7GKYGMPCfFxA6P3Y42KhM05JDr8KRi0F8+U1ImX8G1emlMPzS2tc/5hPVE6o+a+ex
erQfP6va0pU7d4gCOmjZ/afo4Ghb4IhBc1YwCMFQ51xgegM3Utx49oq0AdL8RBl1TD3j5DiXrSV0
MJrPXi4niHo6bi9p/CCKbq5QV7B86uuC7+LN/KBKWYbgwr1COX2nHszjVvZvDfC6w41qIi+gGCxK
8rrEXDTjZXv1l6MJ5qOllQHjPqVOfV13k2SsGfwzUnpXD1BByhKTb7UWcQDM/ZxJhCU7FL9BZ44Z
M5dPmCBP8B8k0NqitbzKY6CFQK88ISyCAylQS7ZRgjgD4y1vbARyzzv26fcyUu1vrhC2pj5HYu1K
c7bj0qWH1lyJhNpE8PB9NVOUwbRdlqAD15eLuenlhyfrJrxklry5//4m6Wu2lMjpl0s0QPjkVEQK
UH5pjnCEKhekHsVmVKFjBg+tp+6GEOeWTpYxt52dvx5zr4V7PF4iblnWT82lJ/sjc5/vN6/knA3E
wfqzLXsZsUMInrefDNn2LxTMur1GIF4e5vURfeyWqMrAgxv5PVBTz3VHOFj6MI/1x71TgPx2GuBk
ETQGLQMo2ATrHuq3tp9iGmyBeZJQDarfwRgvB6dIWGw0Os3jYlS6b/Gj+Xuw4zJHc4Uq3GxKecjG
v0O2WFbjRR06CXMU4T1jv9aisKKK0JONFzdHg+PjaITEFSxpIsOfBsyXaGZcc2cjAIkxPPzOnBru
5/s7sus2o72VKYxCdwzWUZ58kfrKH8/0qYQDyFxn5fsE7vbjqyiX4gbllkELOeWDSgG32qBCl6MP
ZYdXnuK0zSzwBhbmMRncUuhjNXjmRYeSafxiD27f5EOxg9CdEUfyA4rhrtK1YFGJFQqzvwZuDzao
Az2n0AJVsCoxFTCLLnqSDqDUHCQANRK/bPDvBhBH3gbW3Aa2XYVRlE++X7TavYKCv4b2cUJxO+Rv
Mi3lAc4Rrgc8oYV0rGRcQlAxDqcHp0TPPSepsdjSKZ0edlZ3YFITQ3BqwSS0PB/EQKPzCXkcmvZT
7Wn5BKH7nMrv7/TWnaCRil5bxEfRR7JX0XZG4g9tLv1WTBwAmPGhcAiywU4ENKcDp8iYGIsGVbNh
qAREe6fNm5v7THYwxR9wM835AhnSE88VqyhexuPakFf5BBH6cCcETU1bSjiKKTrY52aYnuYl2DHD
KqjymKY4q8u3hSNQoXJeKQ09MjkrqR3HkkC7t2AQBv220vecicRDAjPelTGqVJSwq+7chFOT/OW5
aLAfjAekytcCZsySoLeT2Dgxuu/wrBJEnfs/URc9/LXxa+E/NIH26fPhv1Zm8zd1J5SLqXLmPG6B
4DFOHRLUHM9eHwNv9IkeAnx6y3WmwnFHo2KrMKRija4LoyGGPkrO8MdWNrywYKcQtGMX3ZohvocY
ZT2sZvH+G5zK7f+K4KLQYIAiYwSnnTyS7o3ZfhoMa00CSfYcLBYl2O4oKb3U1M5F+Y2bdlLjV9Hb
Lxfag3GHNgn7ThOKLmWaZqnnsALekf/NTAuJ42T0VGa/bFLvsoykhT/j7erRrqlfPB5pDIo3twRv
5cYBPdZBYAEBsPDdWcOYDBJpGAEOj2Tdt2plyXrziuZGlU6eFn9KZdz5X29DpWnsotkb+O5mOn0Y
Jg30cTDpFw2I41iHf5ilGz3JT9HysN4jnbU2vapOP64onqnNcpAIhInj/FCWq1VmXQ4KnPlTnvJG
a8IQuJDCSWHpNDNIk/b4f6LohgPqmwaVt2VAijChQCbHieFwszP+hw5y6qe17t9zWNZGyK4q/zLz
7JKlb6CwfF7CYbAtDqGe965YuL+XpH0yohOhAHz8xsXR+7InBZhSCToBoN6qQPFb/8eI4tjyUpio
7LI2/GeMDzx8+wf1k/6v3aULg/5+0XXQTXhu4PsKDoRmz8nByuCp2o8FOvYrvSgvYSSBKj9MPKi4
aFFSMoa2Dq+raXFADC5G9gbWpj705U4C+Zpj4EL46S85NnCmiLY58ie15EL9BWbwIrymqPdziEHd
N2ETrhirwv0oBUSbytwYZBSxjw0R/8Gak/ORk/anlsReB4LDBDRbjC1yqZ/K2mfsMOkf6sAfrZJF
KcZ2YdU+oAkbviePV575Ah5jvEQGJXDqpWER4vyxYdlHWIYdR7tHW9Bk2kffccjXbbrxgqDc6d7d
z3UCRA4nlFor2tuEv6WIDTtpCWVj/zLCZj+Y9ww1lYBMOasdq/+4PTT9s3Zk9fFjndbDl1OJsbQ1
qtedU6jdarmnpUaNmOq6vabMusKBqeDMyyHAywovsAzu+kwiCwvjcbA/nzyTFxwPRpspwgIzibrV
w2Q+bz57HLW3xE5loRJ2MJYMUoRRtNaOWcCLaErWLFhI7BU5n49rYc3hJRiKoL2ficTktLOMXMXy
VvHb+8OdqfzPJA==
`pragma protect end_protected
