// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:39:11 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
EoTGoQxQsMu0iJn1059ZuN8UTZrHbm4YLgqJyEz4hKJcgdv8YAukyD6VO/TaMdC4
utkZhve+Bv/gwYz8RJ8FiRnBB3+K3TM5lr6ljyEnndJeqhO5n/ZmY92pOlYiL1Z2
7hTrisCg1GI2hqA66Oc0wHXygqwW9/y8a6YmeE16vFg=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5936)
ofInR75qgJeQFoo7KBbNV8ME+kIplBSEVC4nHYqVtYX6AkU7cFGZzMf1jSy4Vhb0
NK6efPVKm2OyojFHmA1mxZoPsQr4V0gzRNhhrDmcxbCeAYeN0ZNz4CxCsHP237yz
xPkbRkh94GOl/DlGp+mSOb4yy8ttbpGeus4aSY8woZJrdMXSTpO0N7Pu3P7rDXt4
Pvr2KRNY0Oblsu21L4f7rylHevXhspU6NvL6sNAkzGwF+1/ocDpQI4riyWhSuSl2
OmfRR+B5pqQHq6rUGUFT6wzHnTbT0PWYtyV4qUYl/MwGpiQ6Xj6KFnZiD6En4aRO
jl8bgVyYrYF2N/kwkViOuN3cYLtJUcgZTh/5EODlKwzrFeTiJBfDKHaCkUZtkgJ+
+j4Qgb4SKwvVbGnqqRl8CEQHYTWeoeL+M4e8xXGVqBlixHGbEv32FpsUym0TUKBo
EMqbpuQE0LHphs0Voux+fCnNyUfHnydtmlq2hU+ZY9gECLg1G8PU2ioLeIj4Fn4F
bQE/RTNEBDCG8IjZhhIup4MHVLDNJlTsZkcl8wtXplx+2UX/zFClG0RhtjnI21fG
E9XIij2tkl1szqdGFx+q1VcDrd4Z6PMA+GejjSjZR2cUFtsEtW+TY3iplfWP3e3+
kBKJoKBKH8jp4hjBzC5l134/K2wJfsOZOP6KmZN4MZu550FsuHXlEucIhkQ/NEaD
PScGOsUtKHHlLLy40Irqr/EBJTbbMR9ymf9UoD7bZOOv2LwGDE19cOZnWib5P+uW
ZTzsFbwUAT6WZMxdfRKMlgXpUJPjD697cVyHc4V/QiTNc5+x3IepeV9kenojtDwJ
uYRwlgojL+AOn8tWNdBwEynSrVsOkpweFMAVMfuZ/tl51BhhHq61D5oSabRT26eY
4dvrKzCEEcZ2Rs1+Ta2erac6y7qWetY8IE0MXdgxtwWFY4X67ng2JRCXGFkZF5z0
9SL+26yFR385LOHeIa3YKaOJ3HnUjwwrzsnLyZSYLKIa6tMFwr8X5/Brffitc0Kc
QJOyOMiU5ldcQPh5wstO49NdU5ZPQYnE7dE9UQqnAxkByQJIdOUiT+ERyC/5zXhO
TC6YVACCx25j7wXo7aa5rljxSG+TftE1u5/ErMpV3u99u36w4izvqRCEnMPK0QlA
uas5oVQ4FLpvDCAoNvlKeahVOZr2AcTI7P4b5pokzPthbNYl/vpg4/pgqt6Lh9It
L9oi7w7Mugm6YAYF9rhoK+biqXokhtQ/M3WGRoI9GZxr7b65vavhauohe5WbamtU
MGzLHPZyOi6too34+mH4dBi2Jr4OkZIp8fK6HTvcihXIVlve9Kr3savjmlwEnqBa
Yxts1F+IdrhNAdzXWjFz2K/iyB38xCsx+iGulsHNdUcev1ZiAHC5sOwcorygDDoV
6H6hw2VxyggHT7H55SoXEUj8qbcKGaW6bmNp1u0uDVo/noVvzjD9isHT2JA5pvJK
XDua7hcCjOPSAF6DgHY/WiiaycHsi/c0C0l92CzWqHKue/fUYy/NPZ6VxE9h255V
NdfiqKgfvly0zTfm/heMqH3syibiSWkQFJNwcYNIXyZH97IJjmuURfgiqKtBTkP8
ID0sUgbH5o42na3efs+hwDKp19ke6fQuerYk0UX+8ghjy6BZcFiIqzZFr+OUKm2C
RvRvuaIWKE4PhXZmMNjJFGapnbhF89ln0DjGvrXJPxXUkHlNdZRqkVoddbwnZDsI
IQ81Y1kidxd5Ylf7yyQkEKkIcPHGIOlHPVbRlBPCiSKgI5LX4tdPpGCQwKt2D8Cb
mRXvEpRCQ8a1ar7RDiID6JGsTutGga6jJZajstKNUja6MB3GevrKvx7Yap57Vk+w
QWu347/7qJUnTFX5LPwZsWkLRqxgQIKpCwEjk5oXwruo4PqFWBXnzduscCp02qiY
3R66Vbmum271TIBI4M2LohauyKI4wzvxorM8hOOVmNoVcO//hS6EybTzZGjSrGg7
3p+YLcAgmnX6mR7MXKyYkI+KS2te0VRwkXfbh24XJwQVIKYIYT4dGZXh4RETBh4h
wVJxxhNYiZ6H29Wpcgcoil3p5jJfuDFN8SSm4IA/cBOUZF/BKg5q1hyKa7qre5KB
Nyc8dAGmzbJDBFBoUSrjH4h8SlYS1ETulTOELYlcIyPXqex3NnYVpgkSo71A6/2X
Ig2ZJVn9HfHyPtkL4uBfuN65U2GnuOi/zcDezmnDx5qBaDR0GMaVYg6dFRVjAj+p
kn0rv/DvPbsSs5yhSw0k6EJXhRTfTJd46IITRkD9vhdB9SivT3oYCuTpZZqQYAt6
6uJNnyITRJFFSlx8PoW7Y7KAj3CaR9X/baaA8BHeDrnYk1prLipnf2pXwue1msJi
TzfZ09aLVFAd4ePl51+SgWSo4Vk1bTG7yO6az/NJ8FhZaevDQUphxlG5SDItfm/o
HMGR0ezZNbkK5ipxCGGTF55uEsJc5b6uKZlpTur46PHyNp7rWBrNlbXgS93JZXNV
jAD1LtzRo23YzQd9E8V2kPlPNvQV4FbVaTwDH+WbqYHvn/OdJMLy8AiEUEX2Mi8I
npFEMZ701S39azsmtNbw84N5SIU8n74iNj6ok0Gu5Rv9+bNZu/Z7exNJ+lIPgszM
YjIuyyDfrICAZjs/DXXvov/tTtGW/qO1CQs1C1Yy23YmtncW3CRFDndbUDb0rh4B
P8jrWPE3c1R5NXfzdwRqN9xoKUCDk9j47LcXslpBnJ4xe2Q95E49JiB5w3iFAF6Y
geqwzgC8iNSj2zJOpqs95rAwW+ysoxH7h5oEUbdmoD7LLQCKwiEAzothQ/gZaj5f
w5ckTnNBxLJAq8/1iC2O61TUgUhQcFooyazHdUd0NPcjIGKTcnp891Ns8rsa4TFm
xQz1Y8poA2O92aeX5Ugb7KpEQ61EDTPPs8qvH0Z9/Hvwr8E7IPhBV36V9qh2aMcI
k243xd9JQg1LrvL5XkJzGfdu06N9vcqNB0QkNDXTGC9AsUwYyubpDe+CxNZG8U7z
YXiMg7DO/VR5+yXZalCZ3xoukY6Z7re8uBaPPJ13fo/wE6TNP6ohAQ80ixcbCQmM
3Q2skNxdhMHulWjynC4At0GUqkaVBtEYpN5ssPru+WktkVwR+T6zx62wTYFvJQH+
WKOPSyBz8OD+fqi3TIJOUCflvazBz0miqBcybCtlcNll6Zj46dpvUsBSlDHxTkMb
4hZtK6v8ogUDMD4/0syRTxT/VPwfZAXdL17e6ZkmPLNteXN7HLIS8lcs2sz0cvvn
sflD34oBGBLSajjRkXzZgU+EQOBCIHGcWjh2t8xqXohOsRGUdOah0yZPov75sy9e
Oyw4P6Juy2OKmZdGLFlDG0UCxdghgIeH90zn9HOxkx5LjPvjBJCAOMeyPLCrNdFm
H3L/wO1VgQSZDW6XApODZmjxeysBuEkmAzmLmxjprWXPqJ0kyWkvh3oXDlN4FI70
7o1Mu+uckKQhrhdARNoLTuxIqAFYxUKdHLqnCO98FOOLpAogYAg55M/uoYa7BRmP
YyvJmdcCx+oNHPePAOMOfZjc+CwEKqBh2vRtJ2qobH3iTi/XgzzKSOfh5uy3qtHY
AYWPh6iX8UWu2JJ6Q1Pqe39ysy+NGx13gSBwzufu1nqJYoLKD0syDcdQMDaFU1d7
JJ9BciTX3U/Dw23HIxMcfeoCww8YPbZ3kVGUMHMUDP2aO5kT+t1kLufssTAFEY0+
lcW1w5la40Prux3QrH1t+uPGvRUBGaHXYJbrG46VYbvWsLlyZ9nMaKY+MH8QSiUS
a5KTjtVG+7HTusgBptJ1SCDqs4S9uJFl/CjPHFLAQIHuZcCvaLzZBDOH5HzgypZS
O4/1kg9WjMnDsr0jaoLMnBN6gVAFHJ9Aqo3sBXHrqekpeCVvHFEaNDiyh9guXJm5
InVGw9pTGJPOkJtwHY0k64L6m0cy37dag37goMF6oJxEwxcdFOOKiiyO3tDUUwqq
QjL6SkF1CI6xpPLRGY8B8a+bKT+J2Rq3hAiGyYzD9X1W3hgJcxFXWvK6oASdgiuZ
zn3bYisGzTR8PB9IXB1QZzWIRzUmGjd9KgroEAImVxhPxlaDZYq3208jmw44xy4C
+XhEVVUim6xX5NWtt3IXpY6gnMKn/k7yLEqclTnwZmwaPbMnYBIMizyBVCMt/8f9
ZrelzKt/4HxiMiZgCa4216TaJ57CB5A4UGwdIr//ixXvcmJwAOQd/G3aowE11kWa
Dv674ykyZx2c0PsRErH0drDtqweeTAX+kBQK06NB82au8PemxCHP2SLcBejQRBr7
3iMfhZaDF308DyOYxXd4wKaStEcVpbKZVVXy+cJjeCf/ETa3iKZotx7JOh5S/qFf
PztFoUvVPswZ5W5TT32w+0H+d5ycxnG7/SljTwx5TUqsIQw5Il/7tFS9pTGZg6GA
Q0tBxUOmGxpKEyj6gyn+Y7bayhVfFZZjQq7alMR3o4B1LkJJGT9RxRERGvTvFWhm
ixvf1G7JYX+TabbwEj3FZlsJc9DPUublTZBs/k5AcTcdeyRkrtfovvz/e0oVxXVb
Tf8hl1LmA0lfw714I7FHgbVYtWniS4ireMdYY5BtJZ9p8h8lIcFq2itkp3cPPc43
g3FRkPjzbq2fQTsLcoc0rqjYxByTw8GtHMXXbhZhi9aIBCX7i0CwxBZLQ+qacJS7
bqw2SXzuS2ErTdSuUFqpc74MgsPIAQr3rWmT8TY6imiw7a6nKNfLSiUpByIkeJ4i
HYh7CS7GMF36fx0dsEqEBCQWqEW33KttSa2pw+PzxjRDbobWj6Ml0RlqZ2R6knO1
zUVCn1SGd7aEThjgb9XC6f5oEg3TIkvDs49AS9ADYVOFYS8tR6TeYw4NY7rJIKBU
q1nVkRdLOFkbAXkW2wZMYPCAxQ1oZTuBC7ImKFNHH5onfTZa11mewjHbLS/GlECZ
Cjk1uzvWbF9IT1QnSFJwSY6/lbi9tfWEGVAPCJfyNECqU8jtGky30iJnBXBocf2E
LePzAVIsQGCMGK0f/H4e/v+j7C9H3dk3OggcwepPNcNZqQt0SLYsK5uakx25V4Vl
2lQkYoIEwp4W/r/Zd9OgwQ5a7hLpw13j8Bbb5AJpicnlcxu0oPEVIXRAIXsMzRAN
U9Gt61YS5ZNoN9UTJQVxrcY2XQoCs3uKkDmZ3Y7WQdzChEQSo/SH4TPHdHi4pevn
RFBOwd5/Haz20MCbpBUqp1CQ4oD2MelARMB2yKEnoemwRU10JLLF0KFi0OE8bhSf
yITzmgvL7OfPTN076MSzNa8x17AAtYGqKPA+95RjOW62cnL7sJuPX/srI00BchK5
Nm0o7iU4wahGCjxvJHjrRov17J4sz1UzSi8UqU2ATVeh8GTrCXPCW03LzxKedEiH
T0hJC9twKf3tJJS3oEMFqUbJ+NjRT9i/zBWEXgbpmRKSxH4OtuaT/GsmNGWx6szP
x1OQX9Ou6E3ci8tRqXU0992ri1YE9lhahqbJaIhr2CACkItEjdnQRDA7hrXN6LZf
tKZL0rg/FxPWRK8NjCOEpuqkUWhe7uG873sPQhDTkGfdmWHilfN9zK1r5DgRKZNE
9SyPeV7gxAFfdMtXpr2z2EH5Dmf6IJdtrG0K+iDE5QVkm0BKyazPQJz1D37yJfxu
NqT0a4OxvFb7fQ4piRNnnzKGS1O6vciZ86QxWZKPPb26M9w1vVOH/Xlj11aSYNPO
IvBw8/0KOijxGAxBrpJPBzfdVlMN4tElQN2ml+mLLf2BDDPsPr+9hPuynau/gAcY
slegcml95SEEHPjFz/qCnSBbwv2U3I9v40/ofZ/b1xx3knJdGVHZh8P0L5IISILw
X2eSdNmkxTVI92pdKHIIcGwnQvEMDW/KHIgWkQW/5lh3MD58reMBpbVQ4bJE8wb2
cepAZBx2boNjhnQHo371qTHqnCTtw12HIkK1nI0g2bL9sJsrK7pYCKuJwf45Bvvo
5cqDXwb++Cnla8059YyUD5jFpsftSi1lqMyP8S50tAvBIprLHfkZ9ifhTKCDP7wx
lnpjF6krL1/L7ndghI0pC+qpMr3jSDPqZpW0YWxDfyIeYHlWggFaNQsVbLIFOY3k
+0T8Db6yzygSZM1WOa9Kjy6zl3vVEgPtU9h4BL1HVjGF0XPV4eeWwiA2HosGACIC
HFo+qob25srzf8CXnfzem9cshwvkREeIOJKpqPSgzi6GSOfy7XfqbJfY0ahgeMFY
5EaKDCorG8qHR1xm3pArkv36IwFF6+pis30mE15EoflqtyOcP7rVeCgZMpTNyc78
X8TAgY4w/7xdRDeQ8hDJgOHoVKudHetLr26aHPhJJ4K+VgJ6FIzQSIYj+I/3OtAP
D5IUNoxsgaLU6jymlIxCceAEgYJt/Wsk+HjUCpMUoK/9AICu56f+bj72bWWBkmZK
uA/tOnN9nq6nCMiXfgsn2/z5/0tk6CKalogKm0GK8GQlNw3XrE0oXflpbJsqypiQ
Ds/a+w48+2IAwLUUR0IOv4eCw1NjFwPWKhaz6HvI31tsREEBhFj5zuq7zs2fRfnu
oGADzzQKbjMdiDAS29xSYfbFiPezAe+iR+zXNcVJsW0v/zPXPwjFGTefxt11gPq1
4Q2/4tIqH+KGBifgwAHAqDA8Wk69onqxWzB3BcgfBOH+scdogChIpzJ6mV7uzmuo
x8c7e4WA/3hFXhZVelrWcJb2PoQTsrsapLYyQLGqevy38qeckdX8LFxd25hB6Xyj
5vssoKDKwZQ1HldZtT2aAV3gjK+lfmu8Ox/faQn68b5Brw/DU8PJI9XjzsNZVAqA
pFJii4tu+Vvm91COTfKbaX5WQ/mf18sJtFjb+XyBEcseTUghMhQtVff6+E3KXjXB
t176CyGU1Z5YRDZh9I4UOX7Vr2X7e87MreGtTngr082Tck4IWz0L5m0/rTWoEg+z
ARchxFsAkKa8dYP1LFR9OMVmvn9WJVAk4rpv/gk/nAo5LRNqniXQJE4LgaC5zV0e
2doui84/qHsgbTI1nL+f78jRZgo1SIykpB2XxPm+1Fya8xK8IpP9zrzdmLFx28s8
wSaz2X0ty1lw3m39No0hUpzJQISZL47PVhzYFFhzLSC1JUYzsYSz2Ux9HmA/6iZc
mtkWx1eCNz16hnVscyl2JsJihJCRQLjP9La+cOq/wvZN/OeUhXKg+2EhZ6gE0aH9
3cvtTNQca++Rm3EF1QA+80ot4CbabQ4kEqXdFeeJmwSTqmWg0mrjLgaHSJRZR2XG
zbKK7/7s5oFH+Nl0D/ByOoWVtjPoe4lHfUUWYiJbrpOSFByyNAeVx49Gn75HFxIc
ZQEjxQCvGtG/Ra6j9ROXfdJkBHyV0YzCbGbPXVpy9OcEaluuq4L/xjut26sa59Wz
bg1V+0M+sPzCogOkjrdb7UOm3BfayAt7Jm45XZaVLHdeJSxa43EgM4QjgSJP0MIk
D2tIXvkb0yaEcWyUakZJFgWRm5oHruGBKY2ltZ/W/a/v+8L0clHPR+L3wRvqQbqw
HtEAnPqwVnPBh6rXjTRtu+bW/SCLSTRCEiNkhw04wId0OOUdKB55CwhEtDFdJfdi
w6Fun+Q0pm94cUy6dJHlLOEkZOdOFVlGC4mHd2cCn6Gr29y+RDyE2X/+Uowrkwlq
eKGurlMLdPm+ooY/krn3WWOqADpX0f1tLs8OKWh09BlRWDaR5g0QCQep/ZNUeP23
HMOMa3UAcpoT4nNE9c3umTHKxgeamUnD0Gr1uulY0bBcv303DU6tCjKoyChZSZko
U0kEvVWYlg33VvO+75dvQpJI67Z84gkaBKYAcgcVn4I2lrPVSok6gAe64lBralLO
xW7o2fRK0myJI7GT3fmkQUDkaRfsliBIbhrt4u5H3vnrGoJ7dSXgDY1zoDDI23WC
eO4c0UNyao/pKbcahpXmPX+AYScashCDDN2OwtSrfcM=
`pragma protect end_protected
