// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:35:26 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
hO+N3Q5nc/q3arH9kJI9G8mshOpIeROZB//6avf+HdAGrKNJhnDpgYbtUxDa+1jx
BBn0RMOWPkoPif61vYblqpIVpO7LQ+oTtiv+KVwZwyeIk8W7ehBbuYOv2Y0lTtTw
sMEu4jU2OQTsDLVb9KAKb2ZNBGRZZmveH3+94WKvVms=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 6720)
O8d8WqSQpdgkYBatzNuXYQKhj+M977vthTEZS8Xut2vSSNNzSceAzPgeDnSrtEjr
xgL1WK1HaQayzhDmehgVSL+DqtXP3g607lgufFsbltkVqupw14QjtFxkIoOThfll
5ZtBONMJTgr4YdWZJstOmIp69Kkr0GLtgt/tGsFxXrNIHmLd1HGnE0lalGOEkay9
0EoEKwZDWdPRNkWZqhEaUaxBqTRTl4M5/nLXIYDWpMDQB6DkAE7Css5oZfPBDY4Y
o52zbovYjYv2FSG57RZSOM03v56k3+35IHVDiJIF8931WdD+Y6oidOgWbI/x9883
jOIy4Rrnq9os+4vXrOKAEcBYpSDvqqRQqgNqsdGfdXD7KLphi8WVEHmSFWZG6PKm
L+jzNCv0op1LEHOz1jJseWHj+ahVHKIDZN/soI7+CB2G5f60jnun1sxM+xVdg1K+
9YdhsVs807jZOp3B/z2AS8aeITh6aEymPaJ5gteGXSyp1F2jwPJUhRVRHxk/Hzaf
f/yEMBiTNv89fdWxDu3W8UODvi0vANu9M5xxCOdDT0wjXAuM2nCgpofjfYPWasSL
qMGYNGwedJWZwCW46WHrVROuE5/ItcfEF5Vj3ct6hazug0SuFgXtkQ1qh7k9Op8Z
HG7QETFMaixVWANHfsC6jYw1rtth+3AThuBORcDeL4QSdcKghiFRkOWTY6Qha5Bq
qVXehMp/5gOzJ0tiY7zWE9vyK3hh2zU85WbAmA2f7I31ju/efNOOul2l1f4LT0RS
au5DksT7pNeQSirvg6oM3vx070oLA9h1NOP2GL2fc6XnmLsVb6KJHvU51Xk8ssuY
E+eGfPIG4jmIfDz3UXMMuxtmOycVnXR+0wUe27bqyh+kBYxOPaotfxdQuPTUtktQ
7BhH2miOmzlNEvO5EyDcf9Ktjl9jgNM6AXnZBttDRioG1PVem9Cb4VB5ID9vNvHv
5EJjP3GhKlTP7p2FSvQWV1gI/LXtCLk1vA5kW0Kiqi97o8X1kXpFJo0pZGg5deRv
nZ9g9jf92e+SgEz7a4QJ1sHojTw2cWMx2pF5nOFd7oMEi7/pLxP/g48qrAKcigHk
FAHdUpwVViag4SJANwm5cNggNy4D6cP7pCflsjvI0xEEO2/oHrH/FtQwbx6ABSXH
NeaSKBlqZWAoX2KHzvywt8pKV6S5evp+zt8zU1KTLMKEaPiZnFrfTQJWmysqmO3Z
JhYLOkIMtQMHOnWs3FOqM4FGPOkmHdJQE5gdmvGlupEv3DujQCRo0TAY0bXopXz6
Ft/ce/qGHCS6UO8/Cud61W0t+B7cJ8Wkz+Rv8IEuAq2vv6ZGDetnD5mH/y294aF0
GgNolFdUHzGnXB5Db41jknPDKJhXZFbuODnLudQD1ak7tR8OyKqfPeB4z3DOUMdh
/dcijOx/7FF1+tHTCZGgAuOLqoRPC0CP9KWY0FubVbeHdeI/RdUmyFgKTnfBR9zq
oyCexs2u9KhGVCnE5pzRsPkbn0moc3zjgAjYowBrawZWAUAk0Qi4YInWj0oTTkt5
Unbt9/IB0/2c7eJv4WfOqN/OZN9DSG6g/X07EO8ES0HSDSk3BCWUQlFU3z9wwwLh
STD7s6sl3Tc4PbvdZZF8JdwndTJKQWIhAGYPtQ6LNsNR/bojbm7aHRzrwwPHNThi
fph/7GAe12PtmaUgwjW9awMLpAuUycjJHA8lm87w3t/jpTXCo61RWieXlAa73iFl
LT8SmDm1y1kc+wIg9wHwev/uTh1l5ebjlEUZI37045tyugLmA0seUgyve1H2g7rQ
r8DGeM/UPnbfYV71btpx8fbBfcz9/j8W8vdAcccGh9wEKRqeV83WmKXgMl7fB7yu
Bq0J3br8+1Up4/vYY4j6fDIGAW8VNvXNx29NoUfDttu8tHVf1QGucvNGAqZ3CFdm
icbUldNPTDS96E6I0mBL/NdyepzIT0zOOkLqf3BXQO83oWCzAzfnx5Xt9bu/adMd
9RQLi9xP3qsiB2zNU41+aNta37lt/EDrMJ+pejd0Be63SXJOwaimZCm36DiXAn4h
5TlzRi5bKhX7LQpva3uS4jienp2W+IoTpUv/PdUBqgFuD2f/WqCKm3+PEK5qqK2C
E/+1s4asWQUj2Rfwpn1NZVyTKXVLGrhuZz/ctjAlssIUaLbYVm1ggz4FKiwAUj+e
WceAwo4LtMdbp0XqRouW1LfEVc7JZFfpr/XchwOr+tFYto17gHY/nwXN67DOcIFg
gmtI6RsVSdBQnLwxCvhPCXhAgKCI4vJlmlb+jZWQgjznGivylOPAGZwcSFA0c5N6
aQsXHmK4HMqv1Y/9qea07xOH7Dj96fpqlXIzeuDJ6mAUzMqLP6ZvGXS3WiHu4pXv
B/f5DQsEF54eXq/pBA1/PIcghTkQxFtZn9TzKjThfU29XnRfY2RNSXk/BAi7flZX
m8aHgFhB2ZjLXFDhqs2HxBhtOQAP4f5UgaIJfW8VZngOf2FnPIlWnRpAq9tWdIzO
nI1xcq4GeFVF960VL694hyykf/D/Jt3cw6CfmLit9K62l6L68O2dxeaFrGVmouUE
4/M/AfjJWDRAIuGQruJB1qwUZuNlwHQfkC7XQGve494wN3YVukrvrLHzFge3vqg+
g4WmgSFE0BocC6owKz9MaC5nHsfuhMtCzqXB43M8vGGMFsi7/7S6uVhVLKAgoeZj
IYPX4ML1iEnmalmz9zydzeYabEVV27f/mACY8KujBRvEEmrTLYhkWh/CfB1IhuxD
IB33JdwpJ/C3z1h2BFlmf8HWwC22dGVoOtcB6tGRgz3/qjQqFiywYJ8jDj4JqQa/
mn6iHXFLwFs4aQDu/guo/Kg5821V25HKpMqgZaqAeWcseK/7fsKtE3iVwDQOPggr
MWnxsmTq1GKJyDSNORwbH0KIlM0Kag3eLIYXG3uWP/Li7PrHCJaGmknrB952RjLB
Ub+G2U9xM+sozZU+jgXJEIUAzw+TMl3+aM6xFSxpHl6yi/a89Xsfg6itHt7HJLck
t2xbFXOpbpZFBxnPumv2M3o28/ZHOZaMyWI3bNyZ4LlyhZBtD5Qh49KU3OnRyq/B
yr3PDQpBuSG/uyY86n2qssKuQ+5tD9PtW1pf2kHxZkGwyXL1l5FgLnqqsb1k+xUl
mtZru31NdTX8G0JLum8wJsxd96/28L8yecuvhSgRQphk74/cY9fMv8V0+yk1Q5Ds
S+yZzS9BDTtyjRpoSEeu1M/MDyuQhSxERY6D/ab8MhxuWlhu3Bj17UwSAnySIH3n
PussnEVt2sLpyueaGno5SYVuW8Bu7ir8Jk5qI2f3DXVvbLwIMrIHP2HaefZxpJ+a
I+I51mksnJInGQp5BT0xrtZ8x7F2D8FkRgQJGqeFnoUzkq7d/pyE89LOhtXJV5Er
eKll6xEtVNya+tqNWnqsJUE7Mbs/X1G11ELxA9klCvUOge4bAjW/0lVIugwZ/gCn
h3aiME49egtqrXiNxsjLDOeMQQxSwhmjC+S00W/Zll8ud+QrHFY9v0xhdhRKhLkB
7gxwPuDME8NLGBhVARgn62o4Smycy+N+29vrjBG6smI5fPjOnfDCyPtdGwrQaGYU
eyjRt0yxUDH9E4xlUoYB9AQbmOHsjlcEWASRiUK1m+48y1q6xvAzG9/PHeTntkgC
ceqNNepUyARW+TGzLRZTj/U5eJd1iPibb/pf2atPiCnF9FFolvR6B4gkS2+8r2Dg
YXQCHaI3FK+VocXeT0uDHMoLkL7fpY6sJtL9cawFJ0OZb4aromvqujYkI5RXUDsO
MW36Yaec+hDeZvmkC+Z2l/Lzd6dMNt5Lo09xo/6vO0zVNhnrTr1RSrWR6WmpTJ8X
qLpXRKyrXVWqQxEhAgWTI1HliKh1twcE+2PfUQ9Ofw5yDwKp7m5g1H/hR7xUNaPk
kwS8oTJKBfnyhwZ7tPIDy8xnFTpN+3Ex5vfL0yNxJjKtuKBHjUopcA0pvmPjV+nP
J8CRgeIVmds8OaDRsngyekbB7FRaaqOci0W9W0G6hPrb6qU4YJ7awPbT8kEm5kYN
lEBe6DljXK8lq8iKNbvqdz8gZP7Yox5gOEHsFG5yoz4uY0MthSwm5EqWGbkmahrU
0N8PWsH13luCvyBLACAo6rgqffmBhFs3USUp3t/3D5yksYhxEEk58t5Fr5xIMi8p
Oh9+PlxGCt1tHxXHatNlv9vIqsJ3yvoqXXvzSyjKS4mF2087baRzyvqAicG7xdMN
eEFLZUEjlRBsanC3aBL0/DysYRqVElLNazc+92cSiL5uWf9icU/1kb5oWdjStws1
6mPB4c9V3K//JxmIJzAp42wFe8RHGaLHr+iVyOs7Y8OxU6LiRAiSk9khjE1cT277
LXj4vwEo7qMEW9+Z9Y86zQclGC+5x+RvjL4nx8cLKYM8839vdqFmm15e7QLzrtEb
SHGdmUVgPZit3QR6+wPSoI/C5IF9tRtyqBMG8gulK7bnurR9jt83x06pw51T+qQG
tycZAfjnZp2NE+mJxE/UpJ1TT1PyGjlXVFuGrrmuJuc8k2bP110yRPjy6y6bwwS2
8fmyLJkrMs+96V32VHShLzTfhtuUUmxq6OdIajVWE8IsdwSDXQsX1T84w3NVq4HW
YnJDGEZtcEQ3R8+GZ3Kqwj3qLKhMdYSt/vyvuE269/47u0VfSkLItyEB+TqEI1Li
JhRrDTkwKTMVy2HcbaLA6outpaoORcuSuBTdAAoP2J8NF6NrudrdtH1p9uDc/Ilo
CDc2bn7vVqhnazWNKwLykLxr3RhTiKi0noEn+wTMWdI4Vb1tVozIiOjTL7GzHD7p
wGzo8NDwfTFY1m+BT9tmoe1NUgoAXab4j0LzEmpMk+ZGNHq86YtE7+ihiRUEM8QA
+HcIAt77IZcaQWisq8M8/bDjKRsHzI2epl0wXQfKg4xeLYxM6waNy24JuPUhGCaQ
WudS40BGuSQ3M3K4hLKXagOHRS2iBLJdy2OA2DZJyksNSa9Ch134sSIF7B6J3M7K
6Xyo6e1a3b0EFXLTz+NSW6GAub78H7MpWUsuMtA218K3rBhr8lki0mGFbR2GhuCi
1HodPoXbC3ZZ9qBSb/1vW+l4T2RWhZhNmTq8An3izAM+suTSPgjjfp31YewlLf4q
olljP34FNgjZIUh9zElF0ELXMkIj02Mc32DuHFRuXZ8cL7l5LHDxeYFs2BSy6FQw
68OGoPFL7ifMSh61ZLz0VutMVIeVOiK5twKoHmZtl4kQVRBVhoGK/dNEDcH/0aLX
N1PuTC/PPOKGAGWJAf7i1NHar56eNF3qhbagOPlTnQcDJ6oSQatIgX5NK5I94WOQ
BofGCMkWl+13TR/kT2p08xSQnuWGgZA2IQAmeEiCLiuyks1n4RP+7+ZBK+XaYMfv
wkUpGObaF9c+c5kFkIgR6x8JoxvV+wuFXfSOFNSd/jUARHCHXEJyGwJmFK6SZpWg
vFdSCnuDPkV/R40HvpbEMTsRPuJW84E7ejdgLOmZSgmScLzessEmo1cGiHO9Idtf
oxopuSSgjIBdsd84O4t/PV+UJoP2vk3LdcypVClGIsN6CB6J8jirpRxGWsqFIrnm
PepkWRwDvJS8u5NDooV15CPmEz3V9CocrJWQv75eCi6DY9ia54kG6gbv66Szm3O2
hyqIdvjlCYSr13f43nWjUzhWnqTHIEcgAsBsB9sskYR1cY5yN7TaEScMxbdmHExu
UwPugt2TBEpyIOlbE54OXPkvUUzQm7bMMaeIrKhrM8xCQvUdKsVBKjMHaU+azpGE
EgMjhJEplIcEYxfXFQo8nnq1yyFaj2m8UPvYqKHWJo6QSFXs8MfMolRAYbkuWz0c
aF0K8LMHM3KyV2mJoKuoX/4NIfrHuD5UB9JZy8+fxOxQCwfoeprwwkX8IBe/HaEI
8qSxzZKN3K6dV8r5O4Oj14YEKzi1LJztd+ANRqSWeYoIqzSsCpB9Jd1X+VRewn2+
3bQRVcCG82bij9hTyDTQdssNcNOb45CATgMkw04qfa9jboDFaoQntejFxtM96tig
c2SQ+GnWnhZSYCp6qsHcreLrkXJ2RULH/N/SO5jtP6byMweoiCCbUPKqGsfuIAZf
KhB0SaXA46ATiaOSz+d3d5X0taJ1d0u/DwdxYIKkIW6bZoBdOlIjd9Kl038+c2Lh
bT7pu0TNx0rR/BZ4Y6C3lP/iH5W6j5Y6RcBD6t5JP2dL1Y4Qjgrhh/ZNAhXxtX3k
lf8Eo7Z1Xab8UJ7MWXZ3K6o02s6cu1eGBSRPSZe5qK6JBKwajMjHpEFqI6VbhnY8
11s/5NjL9oeQ0mzQ7fmxasdUB9/bVNZVT0X4PcDYayflAPL/HlRq4pfNuOpPm9Pa
1YMcc7YwJa0BrBMm66fqwch21j14948ZYSAFUZgtS9eI/C/31UgM30uL+kpcyAJE
6b3xQs1Joz+wHg+buiRJYYdgb5iBV3/IOOM1n6PyPO85hyilMC+9K7tBVCPUjS9Q
8+5ylvkvQ+yIHISUj98OtAWZ5woV7casgXsXjZb99496mC6BUpT0dem0X0VEPG0/
8cuxVheKcwKRzCkpHIlrAhGQ/udIsF/GowjSRyUUvR2b0JFZf20nOQ59zPCYDJ3J
YzPiUHdROAUnSH38VRzUrxw5cEXMRpX2BQ+jBfK/WKCm6rv7js/4KHvmBM+S+6EC
97kvJ3u9Omw8XoUbqydtLRoC2sKySyDVSd7TYhYc4EXvD+tLuCh840QLs82LL3lI
irSzNJ+FbfYUwfKyddjyIXnRRQKU20I5UeEuUlEf66hQfmpXDYhKHqC4yWkhInVg
xdenhb6k0KBc8SFE1ALO9QMum4FoXuZPzJWZPQb1IDELumOyMxI493CzG6ZHOROs
Uruui2AO1QNKdfhV7eXPKjNwaLsP1bQ1TzMbl8k0zyz6TtDIfv52WoGDOgwwiFCl
cOxTbYYdSrtBAUYsdU3vvkMGT6C0XTuda6oQVc8MUkj03ko19oQbeoiBizeO5rxm
RC+H/ObiXpAValDC/N5uHSMHV/hUX6DjJAB3TS+8uviNF+Q/6DhnN4hXpzwE4mvR
EENcLu6lkyjIm40oV/UpCOep8Zm+tP7aX3c/LiPnMDrHfynTJn05r05rUbsXltjD
Xai3MKKFSw85gUcyEyVKPIgXzCwf9fGNoh/+9smFQsJI76Rj0ml8+5j26cmzjg3r
7YpXjULbrbx/hbVigUs0pHpAdbXfJjKIxRlFAutG06J6sIBQDs5IRAibEam9bN07
NUjgb3Zkvtz9YSj+b93Tj9Dps7dopMs55PBJYTsO54ZGM66fMluenpJ++wJPWpy7
+ojRL1lmSgdlYMWsa5W2fCdL5rtZ9A4pvE7gLzc6wtWxcj3G8SUNcfa65XPfyYIU
Bwbg+Z2JI25Cd9Na+zbfjV/j4uTmTyTKKzGi3ZY7vAZuFzoknHv2t0KMvR4f44XC
YKzkzPk5ium24znzSDZlMilqBjUIBAMqpd1HF4OqnpoxwwfkAvrZxeA+tBL080Zq
48Mi8ot6WYAnhsEG9uzeMAgsQqhkC2hcrmc4/hq2mllZf5lroR12L2b8AfqGhPJF
hxTPUUW9Le3ZwfFRr89w9WlbJyaXU/AsOVhDQ6k6+nzbDJnrjjOS+f6l5S7o8V0M
bvYKX3/oXxWB8mfzH8q4oL/Aqm724o2U/f6Y/boiOhovNL1Jy6Eg2fK35bHTo5ZV
IE2c1EgTQfF3rx2kgZSYp2CTacsSYviN+84vj7zXAvvuIR4aHE/lCnmDyApeRygM
cBeXh9qfMX2yLm1TVhCCFva8sap/+9SqcYVmanmPn+szYcZuP3bj8/TU1y7pgyMR
MmevPJUGUYoM5w087krpL3M6Ub3DeDQcd8/Y0euirldTOGGuNmdyImQP2GaUUoe9
yzflrRCKfoe/J6BULg5XHIsNLQxXV1Bp1kmOxEbYPAmpsCUmdYPcGV7BwdLUWscD
VMrsEM7kiw57aWKbj+eiC9E6/1rjmk83mG/mE8KbdN6BkInTVs1e5f/+T7PGrbVX
fJRSXy9AsOtRGr9wQcJo2zMe6UmlTnFROwzslkgZ55aPCuyIoXUaT9PLYl7R+RoG
/mqgRh4rVRUb3iCqd3e2sKhEjrMETioxXlmHHI22CEzo/L7Vv2mfDf/RTPZAx26E
zjju+gZ6uI8R89Tr4j7z+cVLiUDK7bK6g5MXp/DxXCDcenYnjb/d+7HgrQMP2cLw
1LeY5fTgNJQbH9fBKh2XUNgMoXXWh8dfTw3o0iWpen9+DmzU/xBVBFlJtEA1KK+K
fiqnhiudJO5nrywW6yI/I/e6fkMjNHEJtqodAK/cF3VGk84N9DCTM/M4MGnxNZ5k
UzLJN38Yf3FyYqCEkzI2iQMKyBhLjidgY0KcaW5c1VuoMQRJAIqO+UJRS7IQPiXe
iUsWSOO8tlX3Wwqr3SFYVQfYkPCxF28Jdz6Hsh/8A9KGgoOBdYOgp5bhgHCcYtFJ
lDgBd4Yrj2bkcFQcpGHJAiHVgr6bsc9fzsVW1Yxol/lNA+4PFn55B4UhAdjTnW4Z
FHH07rTw5ggTYmuJXauHFyv3AL5yGyEyn/ouL8XR0WwBlZnlpi7+9PrdSgX0tKOL
vISUHhDoUmxFcVIWRf53aub3YM6X4HkZJea8rBhQQibUe0CjuzwrFeKpxnI2AoNQ
HYyouvd31D6sClTpcQ+djnL60zMR3pO2g2of5ABp2o92gRQtfwkCs0RSWGhwM92S
ABYgwlQ7mFj6nMbqgMOC0Z04LiBSitGteUAAyDfCtTGqx1D3GxODyS16WffGZKXn
2ccOvr0wbfKwYD2nf/ESm6kvPiv6vLCLCrb77g3Ama2653S4xUTDkv+4FK7EViEO
n4wlafcYsKU8YAzQ3X/0dPWfMe4DW062gsyfjublAOp914CM3YILJOcoh8ryO3kS
s9o7mQwD1QRtYGfGknTwjXanT60+EDm8R5WKzIAMvZHStiUUswKjT9KTrCmGx7F3
`pragma protect end_protected
