// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:34 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
GpAV3BCnYR0iM5lddf+dpfIvlsBIjctoNPqTvcANlGaJ0LYOI+LpsuSOMH8zJl6S
v5nnEnJIuWizTy4FPPrBlW2AIJsxRGAucto3uB5ODV+yRcm1dEos6QAG77GRsRTc
CtkHGkQykWt+y5JJk5tUOJtolNrhSKIQX8lKXPYlxik=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 8624)
I1RBqKesfwtbD2BmWMYMc7I9m0zrWn/w1vtBXinv7uzV5RzGXosYevspn/LL+UO5
TEejpJZKq1IQQMVG/iPM9X+ZPVVuRYfFX8z+pv86pMen3decH5pT8mO5qceM+SRn
e3GShZ5zZfDMH6Gwdy0TMgLFA2TwmyUs1aAcO5VXOvHWCjFsI5THShSAh3ujYj9L
odYTIlaAPYYLql5dAmjuSX9tfH9ffxNiLKOif6QFZg7snmZsdry+Q0fIYhk7EOk2
Gqs1LdimGwJAdQQwGLeUF5+0YyjT0uWfL3OdR+DP6BpYsWusZApcLb6tnEL3cKs/
8Vwp70UbdIAJArTEWSl2P+XxrkDrr0o6Ghhtn1NxnNZz5XdjiO1z4KIu1+Q69nIc
Bz8yzS9Wlg9PBQNUs04sEfykh2J+h3fHKCRiEIToWgtfu0DKFUQhM9hhwjxif9Bz
SXx/kkgKtsymud8uqXY2uzzvdSFtjBLSQSiREINpGokVVQ/OsUU0TcnhARr/IJEl
O1WEvrwkiHjU5osEET+u0pDEmAFNHMefwzyQzOwBqe04yJZNH4HxI1KixZTWV4Pv
x2s9GRoLXrfy7kLLEhihllHEya7TcMUgaMZG9dxw57Zhi4NmNwRFy9oUHiSnLuky
Ex1jkUYBZ1PiZjwAlpFyzjqQWoRqgLYexbrBcgS61LFEvKHHxvdpZuIAto2N8u+l
KKUKnhkznneYQQRzSH4LTXBKlCBCsLEqb39aY6PGymEC5vv/LPwmyUziTcc66cJC
gftcuFXepNTqVjXC2th8pf5S/ZtAOZm7+R7SWZ+8HWsznhVIeNX+fnRAhv3TRLeb
p199rGyK8t6BC72txgPzpl6WRVN1peXjvT395b3Rlq3vqcNMNSHgEb5jVD9f2K8y
8Kj57Pude5JyPPzdzMXyoSVtSSty85APuUAqIbOdJXVoJfyfH+bO2/HbrL8WnAYn
VdJH5iGy4d5vYZaVFn/Eja9+noLB6vsvbBJ6WA1hZomp1FR8EcANuAO1KPd2fGVP
L/6ATvHi9hvlQ9l6hezxmvcukb6TofmzEiRoH7jjPumFIUfAZ+b1pXyZVaByqlYm
gQVN9UFgoer+lvAJkUv9kWOUjV6cGsp4Dx/hoWLFBb7WsQ593Z797kmbT3b5fpYv
Tnmw1dqIoyCmByoVG1WzY3CeXGAn47Fms1ZtpqEZlk4SVWuw8UxH8hQkUI3d74g4
jRYEOQz4sYc302jodW4fz6Ss0OexOS0m4pAi1+XQeb99C7xOilDBqAI/QPCtAzLv
W22tIohi2sX/G46m0NxpPo5d171o6aWrT8nkRukYCBak+7Q7LPXTpXLMFvXz7afT
HElkSk/JcQeQJEThnfQMSqPnzANQ7cWpYoYpmcxYm0UZBPPEawofr2BQ3ilJz2fk
pjxNPoFpHexWQ+Myu61hFiOqFogCjAw9ilt/UiumUgWoyYNdpaCz6j8S2VXHQz0V
lVCAb7l4jOHP/H7lECKNCavUtrLkMGGyBIA+a0OTrGKRbh/cgD8Ok7ZoA9jRFkre
T7rE/DtYKuhqUexPnwCrJLMuDj2IS+ckIISMTlrXIv8d5AkrnJnNp6Hyq6cVvqmo
62iXasASt81REusPp3GmtweQ9psP7TzlbMpTvmDlhvt2R9F1t0UfDY8y9s57WnVV
pxE8ol4C/TXIUJ+QSnHpVGnGNxI/q/WE8Dc0/FjGC3gg2vKPmGzc3kNxwr4NXgPG
BoVaYp9cXlrCAiuOcUNixE+gjD/gn96eg7rcb7uzgU/MnPt1prQ6uS7E16VFHvqC
cI2IEOXQW7+ZyqyRy8O8K4mYG2IG7+LlAlDcTfIxrAOS/BlqGWQFLPTtYElHXiTz
GlZZoBUUS2exGaq6dBMiwDgEMafwBbdJKdT7fG4qKzhH48UShgEdrxEy4sqzIjv5
F03CxyaOKl6SzwLPR3zRVo37SFG4LUwInt9yAsEHHVB+37OcL/I9aTXa4PhWuICf
SZ1D67wi2Kp/7OMWcBOdErCF9LBmDXoyn0MJBWPrC2T9yFaBu7sCh5J1ytjMj/O9
ntjhqfYWHI84nb1CpQzTWHLYhi3VVVA3GRKKXHTh7nROwukBw4fD4OEAt1i3ORIN
kCwqXKCj2y1/Oc/luat8Dgp0VhfSk6qYvssDHQp4ZHbq0sNaJCvWkrC3tozj//mo
XXJ0gKzf2JWFOB0XBXw3Y5ph+VsavGqFRKJnmVoBOh6eX7yO+ro7iFrq2e5vTjJ1
gbe4osH22cy9kTKl7lmz83GFKexOJmnwzm8SLgFCFbAFIColgx1h+IVbdVsW3iQ6
6+eAPsmn0zUlZsBmtBcMwz0buZitFggvpkhI96ufZMBjNtFpawdH0afTZYhZl/Hm
Z5u7MzNmrb9Az/UtGeULmwry4nSsqXknpBr61hPM5/WzVg9KED+c/ZfUyWH8agET
NVfgHzZlYrP0ynL2R9OoplomtctN3mGjGO6bhw1+DC3jQDo/FWqa5winEa9U3et3
PKAYIXy9GZHxfAsm4Ix3MFVT66FNH4/Vcqe/4gsAjwUzsg7qAY4LrY0DJ4xr9XaY
FAPQlrSwr3mx0bY9EN92PSQ7Xr31TSWWzTHxLpLAJUYGb2+YTSYvxZQi1cx9uM42
QtSYJ/+FcoxjIioMdVkxcp2yb+Kk+74X7XdY3I6j0+kQ28uw8zq9qdfoQH0orEnh
LdLkxtQfXQW3CDSXXEGIMJhGt2ou5FXdRbYanU5b4TK6BZLCZU6YlFofmp/7Ocnp
F2QgV5UFibPS7pGD9B0+C5AYwLqC/Ig6cZK5AV8w989LTRN/opQtZp+JOF/63WqJ
X3s9HyQgLsVszpU1YVF5CpXBczg5IWyHL5UMQRJhUQ40EKa3GT3Eqg6C8AmeHX2e
+pWHrM+xY1476qBAXS4wan30B3e2NyseI7O2PVCNdWhbCDosrri7diUo2Z2qcMr0
Dv6/D/QffJzc9FJW+FVCXOt6vBR/TBAy37Zer/YOdPwa2xmbQjC2QCEywV1zXV4j
Ckc0yxiYXF48pYR9z8tYcqJ/NXqbjgXxH5nIg/rZojqqOapTYmKHzrXTHw1QwBzc
+F+Bf/m3s+aIeDoQ6I5paCfeM7C7DiLpzBiMoZEDu9oIvogAxR3plcRxQBOvgyEH
pCyyd0y9mBJZ0mdbI2RyYGTOynsPEUApRjjWu+4SgaBOCCZmb73ENFuQy57Xx4zb
tq1d2wv1iD/cuOaZJzSyZRUxdFk/0UgXJIVVNnOSZCM+qK0gBneO3DUFKKJiXBrM
nTti+ZjAZMkydU1MCRejq0AaFi+NQm8j1akWOZ7i/tWneThABRGmlP6ewYNEEvfZ
Q7oo1lG/odjDpAyN033emuTqgzZh7VIwPwJ9BxEOh3FAe/Wqxo2czaeecAiPQQH9
g+nmSR9asvfA5BptXUGonuxv8yH3omlLRi/w5+gpi9C7+ZJZuHcoirtS0ce+FMY5
FS37I8X/aXB7NLte33kZZt9YCknVNil9t33RdIbN0kARzUgVmWAoWU7SpahiRTDu
TTOAsZbjrKbwxjsZxdTiOE3xXRGoRgRhPCiRqw4K8wyjpxQPzOzcn1Xp9tpmLCCD
gD7Fs+oqvmHBtk1FLrgbWo2TB9fFmm+HrYW06pFttubwnQNvH1H32A7sRTLkw69r
GNgAmJ0K59lB4ezarzUXfp2A4zwCo4gqaGJ8fXpPkFv5YDyoWXi5NYj8hq0irkjW
XCQPmuCIbIBl6/+MJZKxbg/x4AlP41uzbR/tY/LMm6Y4IAvBAKMu3sqswt++aE4I
CnNJL5j6Ict0FKpnk09TYdq41oWatusUk85MIwEFlguyFzGCtNGOTEsnyEMGS7xE
lss0q1Y0y4M89d44VliGkjNPH1RszNz98vX0MDL/ufXEH0z+3LNb390AS1j6IDAp
XzX2E0FFmulVY7JQlLqU184nF1HCb5pvipMXJo9naqt64aiyfxVRduBkRqjE6jzY
3zTHiy/0+Amdh82lszVem01ULgCddPAZ8SErH7oqPqmILYbfPh8TISq3EAN3kh0J
t8wWW/oWeSmqtbL8kQ1a8SzKtF96vR7hCXTWHNdflXdVnHKNtrpAxiud12bbhs6z
J5E+3UR0lBlYqYrisQzAxK62quD8GE63ju3jXSKksRlDbbfZh3XJFCDYfHkxcwLr
433QVZgLR0QZFh4u7E4A9+mysX+Ot3ot8G04SDCsyJc0/T8pkJ179o/q7vsbj9u3
IYfdFangQtMLgS1qs59/VdyZ81Z3XCEcwWpigUFu+MXNH4rKNn+GnC6hYoxx0BGV
BMI/AKyd47xF/W2uqcieuySxPK4kNnuy91i7lCRCH4OKuerJmMVYsaO1x+A/YvSm
eHr1MH6PyRbd+vSL+aJOF1KQZA3Yi6l4OdGbps+r1iyZ3DWEGYLIjjfpABvFL1c4
8M5s8t/gYr28JWaWQ0DzsKptMSiHWKxng/2Hcfnt0lxV5Z4GldbFlC5RsGBqtoPk
P6PJe0zav5J07WbrbetQKm+6+EA8O4in29QmLsva8WRx1WAk40P1fH/OUxWv2VdF
RINh1E5TRXOSbrInZfIKcKQqRXSsD+3gSyuNrS0pnf8p7jOHpWRBeG8LWryenVj7
cyI9Wk/JN0Ij+EJjL8ufoNrVIy3uRSXYC+w4Oud/v5/LdVpNk+DKwrWGuQcdAVIG
Ya0vhmpEatlNTFgH2Z6w5FYI6beslC/71/aliANAZt5/ZgxDzR3/NgDt9t88Gqv7
g+YMNityGK7l7qke8nu0qZd9PMBT8PiInJAw7zaTG3dpKVnNbK9q1M66lcBzy0rU
T9d+l9Izn1b2naCeZGEe0Dm7eN4s5Ng0bLO1bfY887QF7oNbLQWeNnm4BovMMAFZ
iOYnWpZC+3nQKvNkMdarrvyaHioqTNnVOYkrkkYHgRGla5aTC9OEUqgbqC3ywbvE
8gxX4vKTL8b/LU7FFZtkFn54ybeIGIGrILwTRXFbVjKZXSLPvWPFFWeLKU0mmLLD
kQIOfwYnKtyJT9zRXEKKIkzutQPbBgqv7v1WIEZNknvNAK9uYo0L3SErIdfaNMCG
Chs03CRtHFfrTi5h3BVzEhr5Ivru8QejR0+wguX3MtxFyY2+dSnEHrGa2f7PMuTD
y18hOMAEK9sLXcNC6zoZTrBaezVVKpJEqE42p+1vAHKecda4uiVTVbQ9v8uxZFaj
nojakvSdI0hpDOkApqtK0KPSgeox9QXfCJ4ybLQblb0tLaqshkFTYaiK03lZ3Nvq
HGVZYDYsanqgo54tT+EZf0qHGtUi0nZgZ8nLczbfWp2B3O9GmBXUR6Z0lGnFEwiq
yi3CvHtRn5VIJ5bGRNX4u4IXRDgzbA+3/p5wZA4bKtDr+Up2qvFW7zZLcaal/5gb
2dUNBIgCWf50hj2VZeTml3I+l/HlXXvEmSGPkAYPb5u+fTTZ55xCZlBxiIbq9iOQ
vNn/k6Jmi7gsK7y2mXTcmVDfgyo/XeXJz4HjVxGony2iUvbvRqWQZz3MWPfvrjcm
vt3rcIBHUPjkGx+Sscw8X4alPgeb5dLiIYdpbdG931dRWIUSx39xEEXDk7xmHJS8
+A/RvLWtuU1lin9OoiNnsr73S74DkhswscsFZ0dOuHzFDaxKKYmEMvGQx56qKMON
d4QiF1lwPKdVT4Q9d1rhtWpTmx1bJi6T0kfpPMclQpbmrIvK0mIyNOEyluCHm2/T
Ithu6c2jyzM492eldb1ElEXya0FkeM8K6kLbvtsZf1OsgkamfF1ExyZ7Yv9B4Mq7
Jfh1Iy3MVqkyz5/jweLEB3OpgmnQC6zlkcBBJUIDKN382xXPcH3BPSRAHz9+daUU
kIPz7GpGTz1qLFD1OZdxvG516kiUrU2VTPgV9s5JxlsHpicidPJ/PUOd2kzK+vfv
72028oHnd0qGK+LbVJostD2GDeUIpGMAYxKmDThkUGwPiFiJNs9NcC6HTWo2Ik8g
p4k0rU4Th7sTBGrfyPnGaKZFpAtluNbZ583aPdTjzdjXYNhUkSL9GUEshrr+Ufo8
o/LKVwj/Bu34YgsiUaSoFUikDSa+HrmQtc5ijlvCMOlgqcb7zrxsWVgIhQpnsOUl
bE4gW7DgluXDQvtROzT/dIStaTJy3kutMhBHyJYFlNeXQFs8LqgOlG5vWC8kK2Se
3A9aryi+OVNm05bDvJml63VDIWtjwye10MemGN8OaURvHgB89Qu5MKlCZEIVzQSd
wc4NYzBhv6qbbh6HmWJEo75dJm/LnBrjd9lAC3GGY+qZGlTAOOyJZFHLj0wf3fwZ
/avLWRS+ahdOnIv52aLEaoDsZIkFKS5Lbsqfurw0s2t800LkARwiNW+7k4CiWXWj
mjlLZ2vHz+B9ExCx5kM+AAALylwY0kgbzn+MHeOixvJcJOeOhVHzLCQuxeXsZGQ5
X/5yLG6jGxhWAmYvFSCszz+ajNjS1Hq7I9lESFbDkTQDdt5phFJBu+TxkTCzM9nC
jvGhsuZRtk4HjsRgD/g7ZgLUMDaiyOGqsgRXZD+41oUIbjt2hMxj5NaDoCava+mn
wILXPCtEJzPB1cn01qiedGufdT69PkqAsMVyFTbL33Q3bmz4aOyusuMTfSI2D9Xm
DwIbUWQ7cUZ7BeaHuTCd6OYr/0avQexdEtFnEkYb6jBkzAbycImOhmjJ6pIPmDs+
VuGX3p8OTRMKQ1fa65K+J/Bycr/uInfptS97tqYyHjwCs/m+/N0HuZy/6zNbPo/e
kkMKnyJbFj1NRna6PuAZUAIA9HtWnKnApzD9tzL1zH9oYpAUdFcfr76M62vz6SvS
7lFjjAIFqurW4j/h+5xe+LdxMgMAsB9Lsh1Na1AI1tRGrBxvBbw4n9baV/lKSHIX
L223p8nco/oY/7Niigae4/IUi8oYN72SlNIdkfbuYTOcDNBgzKvCYcep4aEnoSlh
xl+ygpz6CGUbUZI+8YFg32x3F4ks36e5r2C7/DlXnTegLhzy+C+GIn6JF5F0dToa
x5PuQgWoTU6CVgYm6mYwYuVGWjBBGC9nJ4xj7Df7+B7N0KqLtgih/pQ8kpk45GLy
cy3gly8v8c6Gx7ESHgm7R0PbZRnPYyDKibPlbgyHSFd5nJtosLMZjLwJhqEKk8hC
BmUHOmv9K6tugWDw4VLT/yNBXoQ2f9+4MNXfgN+yLvkbuMEb86UKY25GjEV4RDYq
xe4Em/Os5uqig0UIq0UW286sWBDwfAZI7DexDzSS19bc+/Sr5guB/kQx5NQBB7gs
X0g9usV3Lp99mo5G38DrXQAEkeNLKZFBBmntWlkhGu+8I/KVeEMZkOm17cHXHepu
m0JLO/obd8u35nmhopIcaG4ehp3lPsUDIF4Zs9OaP9ZCPFNWRpzIWHIIT6AWui2Z
JlADqMp6y7c8+OF1jkHgTddSWo3klNw8a1D7x/o7V6rHeALJB1ux7G3x44OJn290
3MeCIByeQW0BcnNk5m26Q1uLtZloZAhLb9yD9HXX4nCw77NmO6PJQZcHgtX+MGIR
slWleHKPpPMxRN4XtT/tsrn0vEY4nh3B0RtsDOnExgNtriGE7h/lJeKp6WlkWLmv
zMaeW5qkUTIcBTVhXma9UZ3KBoXD8QHMnBzCIcLr0dbI9BG0FR9zrjTGllK7CEiK
8YI5sbzf6wyaMUcJgDI802MK0+eYErok7FXaO8OrFn5BK275baF7ogS3G3NqH38N
iT/xu1Sek3qTv2BPYrS5xa57ngyqR4j8LqiXXVeIoS3HXmtH6QkYU1HGF+IzZARn
AluHMr1BUqUyvxCaMPbTYg6sTTMW9394LDr47gLtOxxJy9/GmG4RdVewZ15+Gd3V
ARbxSCS1ZpGuHs6gZuiDOFry8iHcV43cBMnuscfj/wPct/l2aOUSQyiwBSqi3iEN
V3pchFgtAoAblgKlKPRqWP95QmIZVO9B17FTnjMkGzbyHzhRFYspHvkYMs5+SHYo
InFmc0I1k532luIp08XIKxmvzIVKlYWeXlTDfgN565B0e6RU9FPh01Vqd9JtVXIR
gpiZGYJVQwDo5piEqBA2Umvix/UmmJqGK+wZ/xEvvLs5fxTYU9ghrbRtoJTo6d5h
FtQjtsUxN3F6zIu1Tw9e8ljwqxHTt6pS1W4ZjiCIULJuD0ddCxxZnw2d+HZ61knq
gGeqSmsSiwO+BDP0tqLw1/AyOPxi+jk+FF9zEAc1CU7PN+Nck144RMle+6lylmIk
1OmQYn7lnb7NdDDxuD522PCPbf1zAJcMFgdhlPoMB0JJpnjlkbOlQq+unn89ayTK
a5Q6YB6nVUtgtF2RbHoOt26yd+4yhs/SFYH7qP/PP1kPJsIhAiOKiYpkMRi3/msb
7J4C3hOZnihaL57CQYyVyYu1RnCmpV2MSjhCUf3RFNAT4eSY72fuacoINrC1g0gB
QZusva9RjsQJQoqM+3iNvjYh/5zUIEkbjACFO+yzp0NmXlnCVKaULegW3fLJHzh9
ybDQxj9Y9BytCaL4DVo6Km035C2ZVS267SwFrvhq/ZsMidDx124bXPB8iK19uZtr
JrUlnLtlmoB4TAYit47sFgAhYBY6u/aEULWIxxziNQFCZCRJIluS27uX1njHWQfL
yaWT40+NxUVF6G1V4PunhWG9KKZRa8M9MMS8vQ4ZAn79ByIK02evnXdQT07rFnDP
G/7VKE3aVll+uwRwTt5D66Mpjsxg71V3JxAemNM0KZxyCJLgIadkLF8B17Bu+XhB
I7f06ugY581ICztumjmsnDLJIZwPCfkXpaK/ctKCH20bdwI4nSwMRXLaMQu4wHqY
hykb7irTT3upRKAVMHL7teLxpFJZLa9kIf3c215gEdXJsBNLxXsEhu/QoC6kpEmk
waVl3CrQiN+kWQeYMy3Go3BfJJoR1z4G4N6flgfcYetgA2LYamDW8YYpNFRH7LlW
zIpP2pXXxgMzDtr5ZXWvuIAH3iYxrT+bbO/BRMjS1upzzy/CskZ4GetSbuc2MoCP
2FdMJA0y/Cv8M/xGkem4a3hEX2kvR1PapTsm1xWl54rYHJeKZmbjthVY6Vzf/0A/
G7Qfyvmd9Aus8OTHFlrho3MSoZbW2BUvxzpwdNTrByq2noLaPMO3Y2PrSxul93/V
8RFk4PnLiGrhngZd2vL25yrJdt20hiEM5mAkIifr9+14XvpVCLkHTLr1nmCca98x
1LDNH7EpT3UoftpAy4TYBX3wmrScrb5SI/tK3mPRJ3emGLRmADP2y2+tAE4KwlzG
zKA81GJrj3/YkyK/ODPgFJDRQ9sf1L6B1BrbsgrLFooYrw5JrPB1ylp7NWR3Pm3E
GcabWIyiLfHOFmf3yOEP7E4fDf91bb8nVw09eTmUYHvTKN3pWDdi0C3VnyRhNowt
3sa5mVrGuIn/4RFqzS29chUQBAV/h1VqoGqdMogOCv4EcUgyTow7XqP0Ozx/yqi6
wmQZA9Jmf7SbAkn2d+W7Z+ziwi/6vJXz7pQ6qZRk+RVkDBiO6dt2VnmIOx6s1tF7
DI8UiRk6p0SRp/H8kqq63JNJS0J77qm3o/puw1egMtx5cWlilBMuBWMgvQf7L1p5
F3QbFZDXVNxrIvQqGm+vOiUCzRkdgIdbbhk/n93r3NmNGrXn/+YXusEP56MW/Zn/
G+gl0XnDXTREyTwYL+/eil/ax72uCwcig4HLzJcVfWxVbOQimARPIVwi8X5U6B6P
7WXmzzXzzPC2le9uHKCYfeLnwWEehT4RKxas0jm/DGHgNzfoNtrDdJh1hZsdCwJT
kHCu8El2TJJfBRotvvJViJdDa2VYkBnyFd85bB50/7KOAoJ6QAcUDJ6hVS0YMWoa
kiEhqeJP+/hnfZKk+jlJB0yZZfkYpLO9o3Lua4WVReV+ln0xNojSA9/1yzicCCIr
ts8ubnjt3ik/bg4+LCjfmyd8rLomr5mJM7+ZegWL3X0Tv+OE5ajnzLgEGOq/Z4C5
wSCyNIFS8EKW8ZoeE4jU3+k7IxKLZ1f5ab9O4uyAiyLYqOyb4ykfH5D4YJKYGEZr
F7PNO6qT21F1ZDO84L6YmoPe8rji0DqsPLgzf5hmvMbdwSTcBo4GxOEPK4knU+X7
+Xjx1l0y6sqdbjux9cmvaakwixp0R7LHmF/7GwrGvXICDYSHKAr+SjfqRjnGHXgh
nzRFB6qNL3e2zN2JXRMsvLS1QcvjLUgITHnCNZ/Gk7azAiJPspgNHt6IuAVZ9ujL
Kvdpgc5WTallS/rkEi6IQi9OZuBsr4BTfFo3LJxDr17Ji2+kHHRUU3QEtZT1sUar
LknI7DyQN/5SYK+DuXD08MyS/TWLjBCRXDyfKIW3HHItyk8X+nRyEtG1sEFQ0/l6
MQ7DY910UsZ1YVuRee8D9BXVcjye8kkqpv3RPWQbCX/Izl2uQlTCi+3Hpeetfj10
tVxNVHwJIsPHuoHLexGn8cFLXdpmuSEeUChW+3mWx9+JdgmZ2w7oGlxC/VPZCLzo
x/ccqWObsdcg4lOoPDUEoxlz9UoLaO8shCI8IteS3g2IsrMbC8An9VMcC4LBLjPw
SLz9v9PcfC10Xg2LtNZAX4nddTf4XU6YusTzX6qg9TjDqcXet+2kp0cQfatC+UU5
XQ1YENqmwt2mLQdAHd+Zbhm0Rmx/ApXLeGjbKdxNq8koj/Jc0nTV+p+Ul2y9NAZ8
PlijQpRhb4GoefviFM0LzouStSdNq7wvKbWwvodo+Kfh6Bv1POt14s3N3G0U8DBx
hAKJGcznSlHRLZAPptK2BGzg5Gf/O+ldcv5LtNCCaWPTvRRSUs1OMFI/kmagMOOv
uWMZwh5mPfce+XpN+gQf5Sam8Uu5lECimLBiMtq4Abbspa4HIRxd5+FC5Zb++ImX
ahtwmO0C5+S1esdBXkv7FdDTs9c521u7sKZFyrFPSSkzhLKnGEwxbLtWm3iq2t8z
Uq3LGNMzsAsgNIU2bhNxL84h63pZ9cHr6zWbQfas8df2FnZPyr+9QXGOVDa7jMld
vWUfNK2eUPYOWzjy7k/m02QbTaoGiv+L8yo4a0mkvaK5TOtG7OSI1KfQBkFqItnl
PqZOieH+BzshrAT94UpDBL6E121Qo82vWpFNOx1drWOcYk2xJc9GtC3xpXUEfy7r
a2oXnqt1t3QBh8U2Sgc3zx3qBixDHx8b/lPbfzRq3DnUVO4HHblfZRoINm/pfaKF
HWXpJ7EqTJPzxYmlcBEaXp8C+7cDyalV9Iq3DkN+b4DhD+jRbEprBjMj5HJADRVX
ELqigAO7qE7TXtlaOKM7BqRIT4XykwjjVOsWywRvFkn2d1SrhwXvcCghJvDECL5k
rgi70zmQuaWzK1Db5ZajfUGZ4yuzpOryYZe32eRTkpTa+neugdKNPelBBdFLTr/d
XvVdAz5S0qRsoLDYpcHE2qg5glNebYNWS07gi7tDnyChhIq7B0a9PNpYmWphf4aq
64fu3U8KnjuVgpYXEMsO9x0paKYFX8EFUlvR8xbO8y8yARA7w3L/ilRIh2enil4j
WI5XhsKyXAyIt1CT5DbduDV2+2A9URe5W9WTQCJyIRw=
`pragma protect end_protected
