// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
WJwwDvCdCFOdmWLpq6dRL91GC7nbDSOk/0E81NpnddAuOlp2aRmL83FaOIsNpeTHFQsN8bV0Zgg/
3Zm7AVRgfsC0ynB7CqHyKlrfM2xx6ubPnd2/b9ha95P+a07+PdXnh2stkyhQdsBYVWc/GiVoV57M
vLOk2FnxMYORJfXCdeQaIDb8TJB6736h1+7Z6hOhzprF2zFLsW/oJaS9fZI+JCn19oaTTktREXep
7O9gec3S3Mn0jFy7+c36IkT58EpwAGfZGhejJruvoiLcS/NtkMvhX6qagqg1GfAGSeFoqfJMKip3
Tc0f8lrzovclRL7k4+LyTYncXQZHrUHZWNhSbg==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
i/JHRuKP1HJXeSuFcqkf2pO1vFu1bC15tvTgzEF8Uq1XiV587jW+r/c76WyGvsHSUPGE5rdmxUrI
+S7Il0n/xzRkcfUuMkPmL890Nc+ig7Hh44o5bubTLjJBfTPdIfOUpr2e9O1VY8J3JNtyKoFmvtA8
0wckX7ap34cpqwbkwfvzuhwHP2zypU02V/phiYDVGg0OBTv27LUFZIEhGfslz8mF6kawVjOMNK8w
q7Pbpvkg4kZ0pwjI+RC2N0Zjf5YCdRAimOcsAbrhOnFokXGPdKoTAsvgGNENHDw8d0J+EkYOf6Kd
w2uK27jqYdy8A+QLPKNsTTs0brS7x6JROKwtVXVAY2nQ/eKwgNR7AQ3o+8PQmin8p0/U5Os7EaIk
fcz2nX73cwuCfLTF3F4pihIgAmKi7KKWQkupAJHEPfDe9pXL06a44KyyC5is4xUydfh5xihWtjle
F06nXocB1eo4zdjAnXhKZJCZZbAjNub9FUja+a8p3HehUosbC4sewbxi1U1UnINjpdAysz5DEDr6
VP59xT2i0PPIveELJP6wDU08QkrKO5cEoNoCWWetE1IFdBOVUfNPDZ9VWJCRzQ3fdHCDqyIDAjeZ
9quzx+V4dksC+ffMK5USxZiMqk+e03Co0JJiZpQDLAf8HJ7lKzBlPNDJyqju6uXHUZAZ17RXLM+l
RkG0CEAVrluJ4u0HmtyHxC68CVoT6G111iN9KuJkQd4ufDMqyngA+N0jxoY0mE2yg2YY3CRQ9AQm
4yuXTDXuM34Gcx6aSeT3uJdF/sb7GKrf1Mk8E6dc7GbuSW8F1LE2QTH/mFHJd1wuCdPZA5LCKjLq
ei1H//ZLH8+zFtZttGEwfmwcAal6gFmZygPWeg5q3ccHtMqcqfhfIp6okYglDD0ZxPdcZKoobn2N
52+hY7WLmdflWFLA1TvCNzCNPraLESCcWEQPq0OEoyV1ImAnbaP0zwYfN6MU0f/kcCEPiRbF4Hqq
gl2SvvixxUTMQXgobzFzdU2BjBfAFaRUY/USRVqE1iLEmr0VhIFkfJ9kfwcmrX47MkRZWr63v7mq
7jz1yciX5Gpl/k507apFSl7P8jY8Mgiou9aOvuCdKwdicpmMf1qKbVGK3oprhXdtZxybstkOX9rx
QmLJFM9v0iAD+sCCmogAgSrBNbeesQM1kKSE8Dda40+RgcMSCAKA8yt/CATAhZY13fejel2SdKVL
eUX+ngHDeHf1uV+lwaxpxIHY9lqeJo/CUcTMt6iFo6GCnLiA9IiJZMEK0mPMOobSSuyuT04tHLEB
QDqUb0UK7HH0oUTDw0RwkK1HcW9YZ/DutlPjUbyYjjmsKA7ANqLa61vYFwlVn+TsbO/eULKG8Kru
wZeheYk5cJptnMcYYv/JwIIxsdPnjRc/DbCzwCOwATgtc4VmbES+KTV0cAiMZLfAaVKDnxFBTlTM
5W8+WEuMTGV1S/rSC22AQtpmTx3B3VkSM4c0AXlZV3+YuaRFOChNSdc2lFvAgaato/2EQ36EeMTO
jAXbKtEu77B1PQzk3AELc9T4Xbyv5IUs7gGo/uipOcdZcPJ8th0sODEsAoCOgVX4TiXkYAEciCIQ
0UFueb9/wMBKbCPNgF+dl/hvIj6F09LU07GON0voHVSmkC82UdapU+JTzuusonAtXOqqwbOUMOB2
OS2LJlPaKWiWoWmvmT25WC64SbxUlEj31RYwDzKh03feNSAAkZcuE5sRH5tuzs48WBaKZzvfyZyu
Tmf7C+vo1HhTr9aj1wgvMRO6VApJLeaEhwLO10S63OtIaQRgnIyoxiRnR0wai2Q0t6XGGSWD834N
wZmYKbn9ClxNXGx8gMEQLAOI8DUVWNW82ScsYxjS3BP3eObp/SdNfjdtn+8b4fJ9+7kFaut3RWdp
ra//RdUhc1PN59T9Hx8Xk1MrnYnkWD6UfGzuAza9HmhiZY5t2OYFysLEkUy5B6KLEY6wuZIouGjU
wmJpBGxsT3XZaEF92XRDu8P8enYvNXPBPu7H4QjVfTt2xIhBqId3/c3n962g25sWViw05Ksc6KbV
bprGR6Tbqw3WMGLxKOKe+4On4gyMfDY5UtXnZAJ32kYQfdaSX2VXn6V8r+wPvUfVHfKuTLSlJ6vC
xOT7RwxH9DbtQQjlXMtmWpooGnq2TUV3zk4TymRqqv5c1PEVHvv1DzwIv4vlYDJDgLd5U2JavL06
A5/wjUB1h0g4uwJbNoIVIyu5TqJAfoWfyWs9Aqxo5vgK39LevzO1SURhIm7VhR5VZDqLk6TttViy
OpVjThwr+yEyOekwBJjbpEX4MRRwjf6ChiA2d7G0MQ8WDKu/m1MNCAiPo1aHZQZjkMcLYxk/TgDY
sqdD9exHq0ARoC2MRL0ixlbb/mOPVw+pz9uzQGcPlcBAJGEc1YPlOMGxvNr57SRGlbnA+lEeVE27
IypDGwGwhmivgnIPITSWHaeYevHwMYVAp10X/chfDgrzPtNZYDesIvJgvEllRP3FWEcTR0XL0+IH
8l2tVb0DTtKHzJEG+5xCl9YdXEqScSs/uFCJ4S5AFFkEWVqJLIprkf1vNpbju/EXogMl+UF4kZH/
fCCHmuIr2B84rL8itR570Q8Ne561KHspLVSxgkelGITIKbB6mpqB96HAH2UfO6engvreQrShNd2B
MJhIuPA6n1MF0txuU7duFHi6h7LTU5g8+VLZuSBX+0rRgJbw0IQ3QupSWs3QhI53dBcWdZc2BVa5
GqmTIRF1B7QtMPPOfCyaPg0+FZNkCb8SFPzARmmzGqwXxBMTCSVMCbrRpZQ8HRFYf9YJBKWpgtSH
+wCNbyQJ39HboyrMRVlJWJfzV/LwdmOWQMFnjIe+y0ylAExFkrKE1VwvGw+kfqathXTW7z609YAM
1SH4uzSyBEEmN25r8UpnIezYynoWcGAyqCbijt8/d5zrWwfzRKHHDC8xn0WztQw71UBTFz9+oTL+
SXxPDKrECIsFc+zG+zmD850WRHdZ8jY4GWL960Vl0T/+S9x88Gk9lkNhJ7BtOoAREKPN9VZBM/Mg
vpNtkiBdW4QDeFa0PcsTTcKMM1JbN0NYc0vZZ73w/4ABHyywzRsE5WzywDzOtDLDbrItpP6qQ+NZ
qfyvzQ5PPyjuW17p1e46wOCpqGHEA4792mz5i5s23mGdu8/85zccZoBQ8hvX6wYQkz3lbGokNwFH
cp8HVd8wVZL7Se3aoely3Yr9LkSccvqDo/BTmnpi9BNWEv7t9WxMg67czrdVRBC9AD1sRMKuLbp1
NW2jtkzaTYUckej7isH7uDLLoRIZeYOE+arZnuD8hEuNk1NIbudd0Bf+RUqfP2ESAXX7kZMT5VY9
tMAC4drMrVk40PEzsnTNzGmXtgNQPRSU/zR6pSDWUBgNnOlcpxukTTdR12UkZ2N5EjlyFHVC9qrd
L+a/gMG/JkOrUuJSA/5mcwJKdEUYG8KHM/3I63EIwlA32LQpFm518wkuqSkMY4AYH6+cPmjCmmhi
okqAAg9IxT1iVYuKviYUUw6OHe1rTH22C/srRxuT0y1sjMS35ZW7a1tbBUMCTilHfbYIjW3d7IK0
d/xuo4H5rgkwLMLjmQTNZYdGTm4DwTrFH4mxGIgaLdPW2q/vObuL9D3iaj40+WiT/Zod0+c+OqBv
dwc9UU5eUl60t7liJH2Qaf9i1snHRiS3wouy1+dhHmIb4nM/Bnmskc+Hm7gXsLnvJYWjlBSB63L3
/vhzcN8LZAZYWyqFitKZF9E8pyXTD4Bg8GmGzz4pBzhIVWPgOuCIBKVfA6KYeI3IYWD9sKJoCyhN
x08Wu3V63CuIrRFG8iobYQkZsWqZd/DQFbxrn/dH5KAvXfLIFigEPxdqVZrqlL4t+GkTTFqF23LA
NB59S7tNICP5Q+qgz7/D9ReaU86VloWK9JMuojFDjnfxCjeWUBrrR5VqJb/i62ZwAn8ax6lp7Ylb
7vwYd6XfcWPtCj+q6egWGcTcSgjBTtBubziWSF+FKJSdfva1/IZABKAHf1X6sjJEtfWn83ztqWV/
fBQu85ORulI6ouV4YTBRlKKQ5IwD6LSey6ZyJQdH+uZo2XAHZYYjOUq640DMMp0Ur53KVC+sfNf6
TT0MlQwSppL/0k+R4dnIFTDfH2FgDzsFGsdwMA3Ecz0zPDEzEbIgDvFm+EFhIvZC5KgOGyyLRIof
CvN+ClLSlB9RXkdvmiC6B1AbcYJW3I5SWRWO8ccStuyaUcJJt5Yv1w6zzh9D5KmKRg5VjOfhRbXv
ne610SK0aMBefKyMtmLblHPlET+EFYmmPJQYCm1svmMOrxPxmXMEhHYEjTk0s9locPsznQsazYYz
FxpBvCaWfNd+AYqKWUk6WUOvXJmlQ10tQM/DO75ijbZjDvCmBzedpJPMcyZvbFCDOik14+KQ6nZ0
+L8srlw5PDSLFf06dkZfMGlAh8TjY38kFbeL9X2LYOUo8x6eYxIf/WzCobYy3cZxSrdM1JfAtjcp
hvExfviBgB+Wqu52yXXlcXxZV3fG8Trd+jioMUSbzDSDJ5cpUUfGy06fovmuy7f8m/FW1wOr+qwu
kw7tftifPbSkxNy14bFvxDSu/PToG+i7hXihMmdbWOLrM/95D4xXsWi/n+A94GNNwanh0xGEYhe1
M6qWB8r2gdwQ4sqQV1ebVTZThvAEDy4rfg7950bqBnecfMwHrsJfcrbINTYpoASii/rRWBKXhZUQ
ILDJOA3a23P2oaPEeYGW4obmgxP//RcEMak5bCCtV5WKb8cML9efb5l32kWmwtC2TV2thqVg/BxP
onSMYxYUrNmP/HzPeAWHq3NxnbEMi7CAI7x1BdSOw5H/NIzjAgcG7Pp4OM43X5XWvTbTykXDtnoI
jS3TyTNcqsXxV5ACzyop2+UfAJKtL806zRzps4oIPivsn212CRJoFu6UjZH5Zw8Jfsw7zZvu7nib
nsNvqwTOQ9upwLd+QoWlBwvOgxJEfpRk3f4zK4A+oyeZWHYZQvjGEMCQMbNZ7x5flovgwUcwv7Ya
KIRWZoLBZOvlThbc+vctLk/fM5bCUsMfcI0zO5J6Z2/HxaiztRYQXHNnrRwKGCoZLFMB4ySgWrfG
4klr7jn09c/7OWpijDqeZEbHeNv1dsFoBFisqO/UzthB19P2QK3ziUlf5KaQY8YDRFboQbqt9bOy
6KeB//w0gVxS+N83jf8Gndetv+r2iAksjZ/+7BYA3qnRL8MrwOx57H6zzdx5WL4nIUmYH7BuiZI9
g8LBlizn61nEWZnDiDnmfF53VvX9VmxaKBMIQ7N9N1Wq3QGrfw0wMC8rdkFQREfkGBTjObOS2Jw8
ZuAm/flcMy2mGuv72cjkTcrx0rpok2F6zHOYCIQaTNhfE0UVo3dv+Ag2cg0aNb5S9zHeKY3Z0tz9
Yg1XYR7IMFQmJ6Cza3ojkp9ZTmwjdAsQiwZxULhh/NEsv/B6N3iwo9FF4Q5CH9u8CQ0q/FwwocN3
/qbhMguK3wWzlxhU4rwCad5xGNAvoxCI+Dq0x33f7Tat3rQrGUUHl1tr3fePRjznsg613h4TcxXL
Plpev7u57PpHiIGPbQW5XvPdjx8hncUChD5vRyBQt5TJh7gga5ju2jBL8YCePUS7KMJCFSyj0vQ4
My9XYu7xIwOrfxx0bL5hqQ8THUaft0gC6mmEa4ewZcqbIH4vTl1wCKkgKFS+Wf2+Jn7u2lhz9l7j
xj2S7tKZ3YShuk7GsBqXboYvN5p1nNKgbefv9P/Y9wtwmk/mhpv7cjnQuqk3HPqFlUndMBOOORdH
UmdmpusziOykFc/ZPIuA0nUtRHujJQh8u4rCcVHQ2vyDWyaOMdj6h7X2D1vrr8bVZWk5H+Wys+tT
4Q02urh2nx1oLv6xaJG/pCyULwIBHKjtdibK8drJW+EXE0epGISU8i1oPmExjlftJIP6xo4Bl4Se
qdZzGfnmW6piZqGFUmkZnrK4sZdBcwapy7MJw5kByseRSJnvZfVvxfTP8TSWqwsYCmre/TN85wrE
EHdimzNFr3VgO1kvoRYnGuG4kA7tV+owj6EHbXq4Y+tfW8FKdwtejdVFfAqBU3BKU5KmLB77UBfn
MNHFzeH2dxBXZ0t9tYX9eFN8vqAKS3/TcxXKBYtZHxqHhTjpeSyqU3vlHRpOTfMvWlle07m03PFP
IfkVczS3amIKcKS8g73WhiaF/TDBBmjitxwjG4tMXfkfZ9BYdoMFb8a7l4MqMMoVKixUWqmQ5fU0
23xK08bAWnfG8ZSf4kKGPR1ZTcTiTmK/0Ze86dnJGVhjvf9XMVm8hxksvFlnbkBUc8UiL1D4GLht
PP0gq/dEGLzPVaKY14thJKjAYt8WyagzQjXAviMj1dV33Mxie1uMkL8lXcjSzbzhNXYabEn/IKD8
7GcsL1tp/UtVPqKSJRVAVMszK4e8sNXuykgRbgtxHz3qrjTT/ouQORp0mZBf/d8Qe/8BGv8EOLSz
718GMG1xk5iwlxiqgxE6Xc3gzbT6m+niiPD85nN9myDefnp2jXMesPAYVT1RillPBGKH+ZP6MFxO
ccTATXGGxSpg9OLVMQbwJjcLHVn8JJXy17P6T+v9OuBLnwsymkwXjB3l5rLswNAMhWJo/7EgWgXu
ZyYZHsh7QYLXCO3Xq+9UKN+3Qzzb46wNshF4F+pbhHzGxyOE1Ysbe53bOoHTq5tG6esx8Ux2Alih
lOiRuGCZYf5p8hheyBQA2UMHFEKMIKj3wKXpbXj3cj0swjSIRs/BE2qkxm/0cTRWoDFEYX8llPPD
20p5gWmejMalhXhaOuZ4gTXZXA+SdO6AcvL7M9jh5mfq4t73kIsNmbh021rDOe4zckwrFPsxkw9p
2wCOxX2Y0UfNoFPwXBZIc3sxMFweAFZ5Bkmz4xH2RLjQ4xh8fw+/F/ejcb/+cKlCDkIK4tuNbhLi
RPp0gRApN99MppqO2nwtxSyHyCkOEwmxeS1eJoFYyioUuWmO7ZDkEf/8dedr1ebb74QqUpe6wCr2
PBLk0FB/dW5CrfBHErDI1tg1Hp/s9q8DLNHAv80dgoAJxef1cFFwOwRSygSJEOtdfjRYZsPmi3/Z
HgdgVTGmncPOtH82ibtDjs/vMoYCyX4dFMAeZfCnZ9VhTjDGk6yC905aAlOsIlz2k/HHqlF7R8eM
YbGIQbxzAXl2GIuWq7dWTO5b53RTgT2KiGAN1X/OQYyVca0nqtE1naAk2Csf7MG8DYWY7ghrQZyu
U14Ctg3XgLhoOtgT9cWcwfuL8QV3GbhBT46CNlND54vmSreSTVjHcAFoOTQOW2MPq4ybiJ295Xf6
dffKCHRhPt3PlpRZw24GIr1ZRsSZdJzHGEbbSIJdv0ZzIMqn1Wv/EbSRHjU1VzDkHdlJ44sEDGEc
ypZNxzQKyzWldC+bKUEvlKR+6CrWaR39lJMlhMIERN08mnliS+tK057KAcPA3a6ydGWeUUvkdm8k
5x5w+3VGh/j/sooQezXlNYhpZtNYyGrDPoy9aTFJG7Q8w7fESAEYwrVqa9284q+O0eodnhMLxPrh
U4BBTuh4VrciBb9/cRKgaOGADF3kqZJWdSSHM66tHqN+qLp5e4Qynr2FZVyvqk03ZcwQYn5bK9cN
j7dCLsyheTf9YUjwKdW0NgVNDoXWHrMJsB28/lgCpYgnf5RRRDtIXNlRLqDAeduC5h+kZhOUewto
O9x3fpGdxqepCaMhgpsbpXAVwS9ttondve71Mw9yplFXCmyanAhcC0qRKDMud9qcXxo2FLRjukLw
dxxzHLPgy7xufe/MlFKb5ldSFu9A3x6hbDZZiNLU5bP4Coj6RXVCUi/+nyRdYdaUX2sG9rJurq0E
F4hr7y5bYHinRGMcLBZ6OLLBW/n4VKDPfsostgTkEG/rhp+zpV3ae/7887lI6AzspHsfs1i4k+NR
OAQk5wNwk2IREV4zwjPS69U6/GSMZ/1zNpJono11jB4KV/oN8SXAjWnoqnJccKPhgZ42L4VsaFKF
qXWEtTCthDupm/EGCAK3PWoHMCWCABhXEIL07CIa2o1DRjnO30EA/HcpJoGFWEEmQbAHVchJNXKm
mcwLuSIWxnXj3eNKQRTH4OXok4Xhg1b5fo1Ass5vmL1DvRr7+v8myCDfF4C9PgX1j5pCjmlZ6F03
pj0YgvXjdT3yiidzxafrxobCVdMMzaaIQgXTxpDlo+LdxYQBfILGOpoVb5qBx+xTLhWNf6Nx8Tm9
hj9AYF6Q/CBma91bwdqE6vfWyYePzx4x0JxSzG1e2/I9ab0NXi8IXOvyH8vK8Z7V0uFX4L6hGhdp
QWlRVD9T4CuebhJEidjemk3a3kVfN9e+OM32Hzf+XF1nULdjnVAyFm3872EthPtJDx9k0bjjm11s
J+CxAwdChVZR9iLi8akL89Hf7iKF4yIOZ3lLB7bNGdZ9a6w3ykJHhc55f/XeIIaKco1QUzvtIfV5
fIfBNHGcHQLRjrxXSG6ovTFCpa6kJA68a4BpJFNk2Vc2F2x9igUGv1WalLOON329lgT5FK4FBxUf
wRozGFH4ea25sirtB6+uHUA6PCgGLOOIwTdAuterbLqWIb5r/FZ8dj4mYqdw+cuVFaXxuQqvSbJG
EKpHkzymu/86ZlmIO0NPIRXh+kkSIJ+c/hy8H6p+nLZvyKONKAxfjxKRiXoNTEopE+AtOj7hoV8S
BCUSWFRHcNOt+78BKdBceb08NW+TJ3wG6hanzuEwciaMsGw6KY7Ks3ZZqh81uS/IO8dTyHQypGbb
6RD1vr2ClXOYGzfLYScWgpF+Niu/xhumU9ugIpvMeJSGaM5PXIKFxMyBNB/t1wXa727qd9p15sqq
RixFI5uYk2qSHRpTO9QwAJGcMxNz5C/kbe+wMZpXN6HviJ9Y2CLWg/vYt5soN+IHLoXGgx2uNk8A
XLWXvda3mnsyb7Ea05FSAtozi8eGULlrevtxOo1YOeHPZf2GA4Pdtu7zb6z22bTcRwr6qDlkw4Ef
tJcvSKuFjm+ULiGGrkwhqLTBqncFkrQe7Todg64DetMUYs+QAtA+s8Oezw2cs4pzKxX8hAvpWl+W
KQjwhLIVBPMlRAUNmQztP3b0bWgLu4FE9pSWMfrJ5YaICTDz2WN3KkiCdonQ2hxGDqEh0cw5lUOB
0OpgJ1/OUWVlK39RWhErZ18PElK4z6C40XHDyiZhLfJSn7IUP+o4aA58WVgXyXBycNc6yx8n/o9/
VTjTnqA+riRuAXxSLRTRPRKKcxIZxrgc6NI7oe64O/PwvpRhs1NI9WK4B6Vfmpl050ExOS3l9S8q
MOXGHqhufEg1MaMf/azFeDq1TpQyExHpveg80FRy+zXW9eeoPxUhuTPfVxKdvjPaxDijpoGQDYyy
RdJXtC/FDoXK2I9FQ6ojgjvYqUIKY5RcTR77h7vxuAz5DDbHsAA7OsV0HdKVRYZxjVAOlTMv5gK6
wtvQmmXVVeu5uxTfE1/o4c8GIER8HQCcPUrqag2/VxMYFwvPhBDBnnonqVv/WXOMZiEZHxJD1igs
NOcdBv6ttUhMVTMy/PFA520k+bQR2rb4qJjlnLrqN0Ds2/ZiMOuPDBGartTtsv8BnB73r1qIy0QE
Dqj48JMBVaOLKk+cFAenAdGSPIYVi7GHw9Y80G5Vwhm6mIUQHm43T1+u9pK/CWjyDetSZAFPFHjf
aGXhsNNkPGj+H5YupbCcTcePma1uULbPYYdlvPUnbNup8gCIopsAIfZd89T/HFHFrWbx1vIi0uPN
Lz4yVUDZAhRQxNvmyLMOuTf5GDGp59yy5RaUYcTtHR9XkUXGOjKtw5HYbOCbJbibnt2MIZ5Tt7/d
5G5RxAf9Xlhjpe7CRYRUFzMieOp50oyOmC+MkMXbJF0U08ZaBY+B/bXeJfQha77mmFZIomj0k8P1
Y5Afud/FA4bX4JOeS3TQ5EX/P3QIQxJx564X8SwiWHBBT1GCBJkxVgRPFRlkYQFt8pA4tJG2RBzE
1fg17xzbNdcZ3W7RCEUV48HGdZXeCoeP/e0gYd1pNz90JjReFOfWmD+g1v2jXTRV0FFMY6XmaYVu
xSLK6Te/iQpocKeKVWRyEkgY53A6EyFKWOT7fmzE1ASYIKO1Oxypxut5sPVaPJ0H5vwEMYGyuYxQ
L4ao9NdBT8FevOkjcK/qwcANUXPO8EWh3t+GisPEWvFpfBkhKbR/nwIKp8ycfSsb8xRomkySc6Xh
Rt3nk3etQr69fioksLk4WW8kyD7PeVPGq2LnVmCBVPIJxMsLFKctwspf+TniVYsJfbYw4LWV2plb
tAgYhqLIdktCnEnagAoKyVsJccHX4wHwDif6a3uFrT1+awqoKfcVsdQcZuO4NwivhVSt5GcpD3zw
lEQi2rnSqgopp1MrkhffyecWLNEZPL2lY+1fUqgrQQJVyQlmrfR3zhgkuYcvzBDdloL08B1HvGQV
L7PBwkyEx5TSG5NOJfTm0w9ldnIJDNScXJKyZkCIHHUCeiBCjYKNVt6qxrUQVRsf1WPGOTqtCiTx
LmazZOfxQveLNwee4xYM4aie14U5TnjycXXPoPgm+nw/vpNaIlwZXMEXDS3sQ0ToYSdD4m+JZp26
jfv+iDoRU9muLA4y09/X7Y9G/bNS+2gaeys4wxEUw0xrPPYIw9omLtZr1g9Ca0gFEmF/xtWPWJLT
C5RYs3bW1Hcz3+pLOQF1sy+AHcJH35R4T8Kp8OAIZdJ6PWFRzMFkXUBTMQEklWH5jFP3W+OBdZfW
3Ky7vtpQu3yshEihuRJOfW5luTgKdAjDBR1+Vw6+FY6WjuDzoYKDRJWGL0TI6q87WNJh/7UxJTqF
wlxSEWQSHg1/vtta0B1BZ//OsZSzqrmNKiPXhxTxQOE31DSCVGp19ucRqWdn46/OMDHwb1PqsBbD
YBQ3EvsGU+SY36etJIM6dA42GiPgDTaZC7taygE1Ey/Hs6xwCTJJdiM+Z+XBO+kXaXorf2t0li50
M280/75vLyxP90wImqxKqqKK7fkDhN4LhvEZV8Rs2iN5vVEdp41Ru7E0HT3Hh7Yp1xJ9eDJPuDoq
Cf4BRfs2H8aPTNRhvnIo6q+F1+7p9VNAH7WRn4vzhsB8FdRkoYhy4uS39AaYXP2R97TckH3eH7+v
rg0Rq+PfIGMDxwRIHOlkFi+WXGVuXmYV+aODZ+hTfo04cQPSHaVEnTahEJqtvXzcpMI93NbJ2tba
nILCpE8ZVuHYkA6slJKEvlO4Oae977Iq6+Ne+Uij7yKQEpr/VCnmAp6G1S0ybIXyrIUdxAKc4lxT
OLX7KgBk/rO+4W9dDFBHVFhDpBdz0DObypr73nDew1RcxppP1nQVVEaZWQSiKTCovyE4lFOSocN7
0fKTpEiSl8xySgEUPXBBkhexgILnZJVOcO+fzex9HmBUxWETmIUfZseNJFtiqZt0+fetpS6iB28q
3EbKEVV0nw12YBDMoErlc+Da0d/sYo4xZiPI3IXV9UiV4XdAGXG6yGp70ehwgWh0VAgQC6tbj0xO
YRR7Oyo+ZcmSJ6XTXX1Hkw7z5ivPdEMN/Rd5lXHVOjDdJPEdF2xbyvEF0aoqkhPmOtB8zWl2XuVY
kZ3+PrB2WPxfWcIdqTtnhbeVGRFR9vzkczJfptgz37k2FtnsUh07Hlhu/ljl3v7SvtsLYAxCCynX
jyQS62xzwNtza6AKViQ9NuG2GHfQs8NCejIgTZ8OUaPZNgR1KVaOlpXt+6QZ2QNsToEf8O49yszl
HoeGEA2ywrHJPS+xWJOTNkFalIRCnt+CQyYorA0n9Zvcs/wj1qKNhrsgl2MqeB+jKEjavsCOuR3k
z/wE0i6UxfVZunSIA5XQjV338ydo1mreOtH6TRf8ScpTLBitbjQLAwwe3ngVXo+6coXtgMmQ3g1+
Rosd7O3Y74vHjt9Uf2VnfU6jdCC9Hm0ahwOm8bcrPCPeQw4QJI+2JwHa6Z9K+iDmRZjAt4dRWEWj
2Z1D+pC/kOpbvn+DvOjUWB8+TgqajjRUVjNvFgF/1cggFLl7NGVYBhVvM1LkIBkHrf3yIXoviYcv
Lc4CTdF1p3Bs+KHmM/onzKdiS4zlsAJdUl2P/Y+hxA2S5omtLEsoY7t5+lbZEizRldFUr+53Bm7s
7NoYyukf4Ww4ZLbXzVyAa+eQjLVWNkgLTcjCBCHLY+uE4lUCgErLKr7c6k52uk7/d0/m+5Z6CZTF
gyPn8L016hpElgVQcT88bhAN9gSI+72BXpPY7bDDngmZx7RJzQNn2pZ4tVHVRQ/mBJ4LiIEghcHU
4LLLsVZEliqDKacNoFQEu5YBth6a72RKTele02Vj97AG2hKfzxv9TKqkGjPypQ6s32hyP0aDFKkN
r/1Nd/Q+VTSiXuVOuihFZlWH7sApv0CiVF8HUA05QGPZSj1SMedtYKWL2AbxqvWu+r72BmoGdp2B
vP6a/I54moVELulDTDfXVkl8/wbEdwYBywGQfXx+TVnBwmX41K+77bmPGKI7O59IPOPwnZTvzLO2
/DsWyreP1+wcL6waer2Sncvt4TLgkr/1xVkNFa0erEGhuoFYDjndmX1ri/GT0uEO/v+c5e1NL4ek
BajZf8M1zr+heLBOo8Sz6S0uyQA4at5DDiGQ4UH7+unRI/EKLfWtOolnkuR/A0BZgJxMMar2QjqQ
3s49WBF76mts0yjgZGxl/pE3muJgg4JqU+RgqZL7KHHoFVEW3fweZQdLzqpA/T20wW3n7wuO29ui
X0J6HaqXbYcgUFVl7iKdiGPythZjnfcX1Hbf8LKc9MkMeafEISQMpM7iH2iaCeMCdJpSSKXm14e4
pprGvMSRZn2ut1IybMzEKTBzR/3OSxJxR0BVkJQvy84UmG15SQ+J2NNLrjxYVB8P09nS3BaC0gxU
bc8TYUvhENVfmYWX7VacbhCr2+17ibZqXIXUk+v5BfnQmGjRu8WJ6d1LUUtomP78/ckW+86IbYH6
XrdHJuu3KYO1QGoLoPMjd2HulKvnFLCDN0rOCy/Kn3DzNX1DPF6Rz5XWR4u+L0JcRDNBaRB5goiZ
70Sb4hG73GxB2fsG/20rZjY58+8Z5V5HC0z4K9foKwQsbwgjSsnn/1yT/0O9hZaUBtGQJJ1zNr+h
omo8UIKO7EGtHDnwc7ADTLv0cCFmWHUIGFcvLakjCyR7OdO2QvLbmZ1CCXvr9+oILAHLcsL456Yv
5yLPKjVD82MkYzZ7GBTSopOTYVhEn8s9T32kLziCkDcP5qUV5iNkKVnbs3B/ayB0fS/+7mHhJ0IF
A5KYD7FbAI60RZfDddDU5PZpHmJ8+KiKmQt7qOI9r/0oL0j6VwftZ8SQ89Gerf3g+4kLxTRbG4uP
bI7L5PgXF178W6Ov/GkszoD/fpI0ofPGtHnWZ1XE8qv2BxaYM7DzUE75y/O2jJiRUiHD7CN/8bkX
AlarnRHDbqYU86MZ7OhXuh+ymOZTSK4kCNbeVqaM836lX9P/ULSaxtAwwIgQQ2pnh2SUEIYdlGd6
e4ddi5ctJxno/eZszaIfdPopjKxqt+f6eho7GJa8L58YdTYoe1bxo/n2hXpPc4DMX0VpFCz9KzG5
r1krVr9aXNpQEsWB7gvxItAjdRCyQGKEC8a/j9Y7zUYfb2UnJoVaeGkf8qPOr03jR5MOhDLH5npO
M4D/zefNm2rit2O4euP2+LT6AsF4QLJQVnlXMh38YLH1vh0j88yIkc5fE3xwbl48pKxv7BJbiowW
7jwWNrvL9WKUaz7gGnliBVmP4hixYp2TCwmrBvsPCxBUmJO2e7/HhHjlitKOQf/ScY1Wu2pWnl3O
+5/8J7KJGtMC/Gq+3qn2N77/3joQ8MRk1Fef+OE5Fd1r/Up7ng0w7jBpGDQvKQdmHiKJc/heALtY
gFNGaShOX/YFLTlq5kfCuVhuu90AnR/as6tBrEmkkBSEemqkJkibO3DRYU3CaeMaPdgAJ+7rLQP2
WtMv0NMZyuXmigl66UrdMV3iEdcrdsr1OrKZoxtPA0BHyRG901EsOUiWF0vwWiKMSZHbjMRnYm2t
Z2m9RddCCWI0lvKf36Zzr1rhr+ymt9xfouhGQiAYB9rOnKmFuXFDkYi3+Jhr/PsWkvbtGdBCJYK4
n6CTah9MG4BU0bkU2/pBlQ4HUBFjMPbJaNCLsdI+ExSvvuh+qQeWRe2tg4HChZI5s53Gu1eIM6Xf
5zVJsW6rmLs7PvEoA246gTfNDeUspk21zgY3ATvpa+D5K4aLFy4Es2Y8gddsUcbUwgF2LwZInV8Y
vtMUU+1yQVKRfFdOcoBUcqvDMuVhjpdTbzkOVe8NhFGRyU1XL+8fkLh/I+j3SMSwjzXTcxTfg/7w
G5UsJv3Plwfx4+2QuWvodC/b616Sojy1Oqk05rF0pwaKWIfETp0N/+qI8NFdvD3VtwwX6cgCvxUh
NuY//HrCxUcHkvt7cHlPMrAb2DhvR81k3oJkoRiU8ZDQPUVNyeC69dimPHMrZu5Hxa7JbhZKnIW+
NIvUIWt47EY/aXKC+6BKCBBQpgnC0jQgLZz2Tl79pv7KfrCbbMncuRD+liNsDzHL2WivtUbRetJ/
eXOlVwqpuXk8z7XSWv4QDS7gbAjjpihiXqhPs6k0kP96LaA1sv5o1jrOMpbHOpaUcwVUbo8LWCAZ
KtfEs8U5BDqIupoLA1JaTvZrEnQqY9/ctlEik5O65gaolmnZvZh6VKWeQktxskZPd+wECRINggbn
axee5VXJF0/R3ms01jp1244gdnY14fkQm49DV+gUJk4L2BfSIki1Pv77Ot1MvNdwtgkhLo+WlO+J
b7Owdc0Px8oXOXkykJchiPI5EpnPBHdg92eAb7gEpFlWREjnnVfbI6qUZB/+LnEg1ntK0zN8cacP
Ja508PmuyYDDjJz8tT+fZAl1F6SEIm5LETG6I8nqaMDsdETWNc0c3yuvfW2cfsglBV53ZoGJitM2
8XeUkWUUKN9uqtKoxrHdgL/eFgdbrY/SHdxUJTVZlP0xthQEo0r0H/PhY1ann/epkIi/DdzqCo1c
h+ihvjTqcHKc57MHV+FDPYxQvjJm0p+RbCa34nGjL4OhmmE5ICBl6cb2XElaFggqog7Tt7sg72Pc
otr65RoVpr65yrLlRZmrmLuDXkFCEti8YhCzLw7RttyjUcdq7iudpO9OQKSHMyJU8bkZMt2Zychz
fH3IFg1jN4IVJg3Dn3hKEAMe9hbEP1cnz7Cz23vuV5hNCaJLBpKG8TmTGL+CbGR/R7IIeOPULs9d
2gmtqWGWdfoDnw0UK0s3eUEOEKmE5/GZDFkc29NFU6FMrbr9sDhUVUZ4ZIBmTKoLqY0fVf8tosxm
WkWTsrHNlzuLzn77So99gsmPS0K32gfAja5jum+vtZvZtQCpoY7Ol9S4OKa5UCRpkShxCpHVlqlU
Hpiq+SpxDqgH4TWsHFcW1srx90oOxlxq0xZtMDpnP/iOrRJ1zjK3qYxV3kgxmVz9o5V8FR07RoAh
HVpqHlPL8zqAEGUe/n+VwbuVU/5kxI9EzXkYEcqiV01iEi3yPACZ9/z4eWUket46p50jTe3k015d
5JMdyTCttZYmKUNpGpy0iusmlR0tJipJhAYndsKu4hApWePhjSj8P7vHSMgBk4NOQuCDL34BfOym
S+92hrzHV5GIeS+fSl/lH0UxgHacuc5UKXP9ThZ15wskXlg33YCf3D3Zh1eGU228EtgfQRT1qz5/
Sw27emskHCdaSTOoeXsq+MOrpp6CO0z/cHEM5Gudqt02OPcBlB36KTSDBkN6fkVlWHuWrHZKVjZs
LVNXMPcGmNPpkBIocWRyh1ym9uaSX+7Bd4GdiO1mZ0zY4j6GSTmHndFZKslvljQJzgqigLuqFVWO
zlBxBxHLHSPikOHVGNMnq20WqfUYyBGiiOoIRovFMz9weDbZFcETgVAOdF3t6dklKw3/tJD6RI9X
tZswrS6Tear9ed4Du7tWAJWQBDVYdyG7QCmbGr+URVoP5K8EOKHCj8U7qQsjlBXRWBbWomvMwaCa
GwsZ1ugIvU5mjz5sxRzqi5/5ede7YOlFRFNEioK2U+JlZfoRBh9wk4Oc7DpTpuYnSpdZAFGrAL0Q
Bc2lrGhh/B8hcm0k3+S0lAllcIjhmrAOw0ntjOt8bTDOdTORZBaoj6qThfuz5DwkqnptTOPNdreg
72jHenalSyGr8uJM0ARGvG9BIId4v0nMVnzwtgPagseXbZGJmrYY5EkMTlsG1m4WzslWmZoemgaF
qHJhl6RkO4uW/xGkQZOGu933TL8306qsVS62MkgwqKi666wJ31atjKssrdtaPMrQep4PyJTB/OnQ
nW1Vvw2LbZOcRz3NulbOEQRs/Ayd/mnl4JqNE7SXC3weVYPiv8iCLuO/qfB3Xiy/Hn9ORuMixdAT
tRbhQ5AFYXcy1yae/lYqsJblJrez6KUo7bW7UPG9e9t2o7xkdc6cQFwMw6/xRhRQyhZH26Zz2Ps5
+qZmfp9v5/doZi1gbb59l0TwJa3VFz7ls3VlsnM/AFDAcutovMkucqCHCOCVljrXJCJg3Yh+YM2e
UTVLCzRNbT/VyS0yxHbqxD1eYKLBZFclUs0Vkbuwya6TqrscPGoYflAuFDZ1hGUeCLR3Wba6N/GF
cOYctPB8LgSo+R5gZ6U1AkCmEZqIbYOS6my1wDaimzmkgf1nJ0L/eWmuyI9RztbiysrZopzwKCNM
q4eoTbSaGHtEPDm7LAZBj1FWWhqayRIH8gOHmXoHbvWjC6nqjlEi1Fxy920jhiyh99S3JiWrBLE6
HbFl+fQA6d6RHh3/u7gkLdVgDqqfCYdxD7WqMZoM3VsCPlm0wyDL4/3XieYwqzWWi+va+OgWlJ+R
G4yCBftmRRo6T5YKIqHo8wIogHhCSegKfOn1dXhlv+TEezczlg6QPv3FFyoviJV5uYA7EC/ZI7py
xVfSQoppqElT2iwf+A2C3NLlIpZ19pvXVarAsJoBY0Bui8YeKfp/6eVZlIFLwFD4ljSdmEULEuFy
KUDQhkrowiOblj+429EAWxsRsrw8kKlynkgKio8D7mbCU5QkSQ5VhHriD38DUfEjga+SZFLSGvVD
Li0i3Iv4+DO49uQBXdqk8mZhA62p/pf8m/Nl6mq/sIKsIl6mLaR31Qzwge+NgAr03O5hqunaAIjT
UVglxH0eFf1lkeJNXQFalLlWoGdke6KDTT8hMopeBDYvpU/lh1wCF+Fwy30tk2xfWn6tlwdJAx4g
Aml5LitT4jn0UuZvgq+CoeO8EY65AFTMfY0WxSUPJu/0+BfTGPBLRAgHkUgZjn+NRG/Om3kVcmhZ
qGMXr/7bOKknFNvyDeQidY9HWaPIM+SVzrFXSV65tdt4P8ryyinmzQ1sr98SkUBePZQbuAwBeGtx
wr/8jwuYxVYhCwSQoIRnN1/r4V48h2kn7mF18hS5LJe60RcFolSpyq67JRMbnJI7fZNQQKykF+lY
/f7EdplJeWvrmTXO9CgPsVfHLLhhvI8WawTNQoziBI3S/sztCmKJwxh/CqUoH3cIkdolvh51Fyk6
6g5H+ojOBxH0qqlqCDH22C4v9X07VSFyWTUNEujrkmFkrXTBSirkBxmGNFhlJlc/wxS3WbNuyRDJ
Cw+RSCtg46CY0C4iAk1hd/iJAm7oB+mClrz7kdME9QnsDFf+XoCYqJ9EESYENX5C4uzYI1jJTY95
gObzjpY/gYoVjy3QBmu4pT2EyGDwhn7Y2jCmEAkcoBFDk64IKuDS/9Zr5v6TQMZx+Nc1dsLwFo2I
+sN4P15zCjsjKgCTo/yPdoZWV0dZfCql6teh4RcJIGuRveE7qb51NnYK+L+3rC6fh22IkoNaioV8
wSXym5kIIiGvPW7vD+umdvCW9lcPvCd4wA9G30Ozut8i+BemJLKSdikORULd21DvBj4M89Wc7o7c
byBgw1/QfnJRYuZjtBYS6dLJzU8556Cu0tSOX8SHRDIqfDTFo3ZVDgfXV69gRuNFeqAF4WJNlQNL
Jtb8vwhD2jJnIOyQJzzMULyL0EuCs30HkPNWx/v3dfEM+St8RlmRIzNAIwUt0kuZsXcsPDir5lvG
50SkKFE7+I5X7k4jmwxx+y4fx28C4M7MJeG7U1Q5WlY5ERZqPPTxOC7TmC6qhTjiFCtwJOU3W6J9
gj7OY3ET+4mTLhQMV+44f5CdEHTd0qRlGDzgceVM2wp2c8VQJ35Orw8806gJvIh1axhAqYwnqPwo
2RnnJl0jp61rdcGkRrx7U1zC5LxnnjzZ8d65wl+sAbsAUtEIIbjLBy5KAb7NXQ3pKrgIJWA9bZcf
JuTMGhR4HCcWX3M5xVJViDOOgUvTBInBQaJ52G1/g0ROsoln+Uxb0yKdPjUYy9bp8AugjPUGbR0d
AqcK9XaNFtuZKJDAEzswfYs7izA4BbWRORenzS4aUBktewe/cBkikoxlhoB1fzvrHlQUjZQIZgBm
7dF10OZ5GF/BzSOqQeiiitDFybcu0JVk00f6yz08hieW1TfK+M2q3gkkjgFdtncGel+Z8jxKFanD
gsW/CB8WAhNmRjlCL4c+Qnqr/54X+wrcdfyKjHxdU6u/aBxqttn13e2NoE2puezudJIHHRF4xKPn
bg8SmRmaazse2UKY8u2rKiXmd1RC9zL+Yjjt08da4TtMYe+TJ/VhwXsgK8Ux01lGB/tABbt6q4J7
J3ONI0F73xBklGkAqef9sgpUua4aPLQXfYn1qIMmKrji8HKEAugbVHQ4+YJtw8Wu2HDpXKyIunWp
I33MsT9L0hO05Y4nkB+zKH5/rzc/hgmlLS4esoVQPL7WdgeKteDifbYsyMWUWBTLp3u9PbfUPOE9
b9Q3AeRRPhpKuLCBBI9kIrxy/t+fWMHmU4JzMh+bBYENvGCZFokDPhPbU4uNTSgwtQT7X6J+n0tk
slQfo9VtUxpNMUhy3T/G+Mb4Lh8rQHbgf/4f+9o5GSLHClS+UnlAmWqCWEDADSEQ6hHsYBNfro4C
dtaEB1w2b6de11OEA7PmzvNv6h4KcRVZnq9VxTuDl9m3oEWnRFkmwH+SZVKM6nCR1/dea095RfbU
tj9bxeNfV4Z2UNozQVisbP+fSmtf54dAJW0pn7QPTWJwbRvG7b4h+BL+ObWnlxdlviBmJE5IrsCQ
T26Uyyhq5nl5XV2wYo6J4iDxsWvWBK5TuyidgyXBpuphT+r6BFCK9KwvMqeNDSCAf1CnTnw+2HH8
ujP3uNyF62ZO0lBqndKbqag/QcMcHgUU7hT5rAyrnazYmKwLNpqsjlFu8b1Aj3LqDhqQsyCdQjVF
T01P8aJ7ry4BGiIRDSMWYd+xQZT7E9YsnGwXWewTcGZLrMljvgvDbN3kOx4WZanLJSniWmyGZuLh
T0UOkbZyU+FRaugNzCzwwwGf+I2I2u9ui/3G0HjhEwaQq0m/t6IZpRkytmk7KhxDG/Zm01689/79
7sw5kqjPmyma+bvVPCNPVxpWOPZXzp1WzxRpxlAcnGgTKSLuBybjbFfGVUs70IOr3LqqYVXU2P4h
4+e9hljuYE/0xNICtoCvAsjz7kuD2ooG2JXBIbhkxiiCZSKpBtXp8nKY41crYREA12MYE3oa0iMZ
EdvtXQ9EePR5tNemjG53YspXSnieFGRcQQmVp9J1SBiF/Wt/FUUeatWOSRxD5AFip83VI0ANkaPS
0Vep4cHTZWNY4p1y5kVw/bYrPS+aodGeSAKXzbJAahS/ZK1yJBVIVBHKhZtELFdQiRSoIyODVRCQ
zfbIg1pMnMy+SF9BdLzFz4Bz2tze5I2ekw4K+Xt/UQjFDnn0ssf6EgeZCFgOL2REeqj87O6VYn7v
6r/NTUezYY1s8fwvOQlNRRtBsSgmk3g8sXC9txrr8OqQ74EanwcCr4oIWLaBlJSLgqBnaT18aDM4
8ZrY3rvvks5ek96bE50i8YETEdSLW/COQOTeW/+8XuV87493E3dXrHbY8l9AMUTdw+NEnZZ/mybw
8tHWdBEtZnXtC2VKdv/IFbLMV+yKLdyVOQu3P6HRAW4NMVvrOxexlSCSeN1/COGJFu+fybHhVcgN
M11bQ+94QadI/FzktB7W6EdTAKPXLlSaEOVNOINV4c8YbE2zpiRKXWM7BUvzy2zudrokXhjbm1bH
HSdfk5/P2HaWQvVx/rtrfOJJbHY0G0cw2kiY4ZG63QsL08cSaHbM/Nw5bqLVlB0OTlqZZ51WtyT8
BzLVSLLojL6ZqnWzQu7SNxxnJn6rQjuEZuhZxlix8pXzPTbNuyKIKRsjdp0YZiwpIOfOfChALSn9
QERmUMNozczbmbOBJHd4K7pJXFcrqVBQ+f42erhySFfkC7X+X0l9QipdP1fZBlniUIrGL1tuJAvA
kl2TK3j6kX2fOpp91IzJs+3x27owozLuYuJfbj03Z83dmAzUG38QrN0GiW8B99YE7yr7itcy5t9q
P7/uscdlgec14zBvLQ54qJ5P3EehghEla9D6Y1D5irgqj6m9VrnPAqMcEk57Nbzjj0UBbcQMoCUo
1sPR8Cc2uxw0rNrolE7Ly0Tb8Ow7KBHEtXrgQrk/GNFW0TtFM1JI5KmGLiCQD8RqKd8/yIEVYeCl
DeoqZ4zm8Nm9sPkjOjV95Dffp++AlZFvaI9fm6PLhuBVger2A/0ljWXo8DtqxCu/783Qnc9ufsS8
/S1SdfHUphugh2spd9QO4nlGhW1sSIEYQ8su2CqwDVg37abKko8ekyg02FNcDx2h98xqOBnY1htY
SsjVJcKSvAO04+462A21nFaSXrueSQLMzl0d/5LtuJ2Ul3q7cgGI40KQXVhvaMRUDA1IF/qfesK5
4hyCKdRnqDH7a7wwRK1AfV3DZwEdhiBiVGlFY7K9IMsGMZ5zW2kjoVkLJ42jddQSTjIY5p3qO+ix
NyXw7D2pXjSbD8oE4FAN7yZWv5mD7bOQVM+mIp62nyxFNQtFy/r3t7UVi6HHkqE5IeGbK5YXjb7C
f/h4UEObxpNm5Z6P3kxLugjyDlWCwlg6T446H2ig2xlm3sFglXpvvlhbvgFcFgEqp2TgKl2Zfm2X
iUtgFDkM5AmxjCBqpB72PnZ52CHFcbWWz7GL5lZMcndVZcySXaY77J0rHwvsSsv97xFKcqrcS1qT
vC2DLfb9J3lY2P6h1P5GS4rQogZB5WhlSzKapCwImZCQacPYqhmazI+olzFaUpmU65qyedqOH7B8
sEpgmFMaIlnEyZ1OPS7zRxWZ1AgidvQKS3g44yPHojPx7lLwUjkRozKUQye5h1TEc41nz/MNSzvC
XjGfo6z7Nw4EzMK5b5xW6gYR58ClvBwKeXnXvFRQoM17Vjw4haKiQ0A0R1vvw6WTz2nW5Qxew6/D
EOVpe/bc/X1Bp65k5+aqmlMUGzLLiRCbyd41dcXQ1rhNQgdaQ1psS/JtEK/kxTxXO6oL90z8s5ys
0tHE2qL3Ljs6Zin+zLdggpMIn1W90pm/Z/FisHTpVMmtk64Iiv+IWdRHdWpPEce/ebBXnI5kJF0q
JAvr8nNF9oRmAJK35UUzvoP9ozbD49VhDlyRBH18cEL2TWFmNLZF0cVWtaDmrxO4ySxMs3xWCjWR
DwS9R9HHwOEn3+4DKBvEfGZgmnnXwA4HzvjVdDROoKe9l1bntZcdrEzeuOowCr3sIBwsDLLpyRNg
e8aN8VSBBDKH/7gNdOvHaa8bMdUeA0A7cMlC/oWU/15JrOYPLFjceY/b5smX4klOYxSQ14o7+Lru
GNEH2j7sdRXiCklY27gOwN0wJJNYO+S6RowfoX3O4JdsRZA5/6LBR4+nBHxC12rJJNJuSLWi8H0W
fJzC9bsP87K3dSNKV4NfLdgsC29ciZGeswkfYGSJUlxfP/lWCMOVApCYI8497rMk4keUjdrJge3M
ok0mEaE7HTXiWxdFdOvjoEvZveTH/0Xe1PtFizfBUQ2+OMyn+a9FYSKcvyLfzrGR79/cHdslX1xe
E6/W21urvrQIrwhmEt4Y7T6PZ/DK4UqhUqFn4FbmNoUnDt0AbfCG9mt4HMGE+XxTzbm2yuaKxQuk
fulsoEe2yE2Y4iieWgizDjnlQlxaueQ41YmGyvSflO2PDeB0iNAvuKJZJcvV1Tjm3TWPyIsrCWW+
m0iw4EGO3EJKUfsiWbrDvsLf71AUBa6dhDamSqI6DpkXlu+jUERwyDEGWioIezC4NMkP/9IkVHdh
y3Ml+tcnV1hY/4JvuSIcUFqbI7lWgjN5wyE8hTUT1APewbORrWptqJ6faLA1Ev+COPcNhrea6y5L
voJ/pnm/pd9J1B0oORUoOATr0XpTCNpmzK3KCJdFez5tYOGIP7oSgmZIT142GMJ0pnRizE66hDom
IkkMVI2RWE7nSSZTKuMgUPUvK+YAncFJZSaGgohbZijPxgJfeftoezTglvM71MPrgUF7VQ03CUbZ
XzD16Yl3f47Aq37jeHHnCQBCVO/i38v3HHRMXCegmWtsywa3D253lerVJ/QQrJnHccxj3B9poLqo
PToCqTwGwgdOAnNJlEKHl5EKiOpEeZXU2D3ftPkTqGKi/L9awHnjStlHeo+sxQQKq8OOaZ7SG6zx
GzLPfwYS10+Y9iXZcIZysSkyBNNCKD4VjLj/yLHUXvQuA327bWGWLgDeUtZYcS35hGDbcuhg9QsX
Gd39adJOc1kPmvmZXnOkog7xnOZhJV3bAsHU5PgXaNDPecoKwzpUyYhk8QDpFpUgJzSsV9AD0Pxg
EeKU/lcsxkKwyGbne37ysIDFyITLQG8dw3byGt/RPNmmrna4oD9OwGidYoCaTl7E/E7+atiLYeK3
1RFw4kvNSRoN7IWJdK8QjgGW06iwHxCWlzpaL7BOSKlF8JLcQyFdrDUm2bDdyWLCyWkEH3m6Mzu4
hIPsol8D0IL9JdcdJsDdcAR33Zq0LhbCQVxa13ZP8C0sSRHn6/X+Qs23JLXPcVtNmIR2HoP00ZVe
YnzTe1KgQIrNQ8IpZx0Wa5InpacMyQJPvlZ2p1/wMn/EFcce728D33NI+/ZK4n7b0fXFYGrVY4St
aQEk55Kn48GsF3XPkqaXit1Tw/69/YkAxstahYbmPNLR2mallljh7ykKuQmnRseHjOnXKGiS8JNq
VQm7wCbbCCU5JDcYmV/+23YUpkzTF/8sJfpCquupjSe0CcWl9BTr6o1jd2Z1n7gSO6bNKqdj/WW3
wiKhb3hGXYwqgUKyPIm790qlukdQ+QoR6UxIdyPAlS21bBdISukS8ilbzUUebSvBXfIn4Pkl1ZKl
6pIu6RtA9dv7AOIX7/pIQuVRWJMdhmhEPdnlxaDWTArcyk/UkXN+v6Vtd4cZFDtE29zcZ3X1B+Ql
yJ5CqdFzY90gjOeMl/KB/aXZegIuxZAGSC8Ez39BeCYXdNOJRvaCd40mEpT9fU+Zi/BjSnk64IWF
kPdV2jPp4uuPB0clNjaD72cIU99x0dmm0J+yIxqTWvIIsVN0gD0A5TXb1kVg1PJls0UfrkVDEZt7
UwIHu/V16p2fpirhmDqje3XcTEa5obdAVJ/e1jz1cAfTikLT3KAdXqMwIRIo4Iz+0pSuNnWOxIQR
Nc39a26y5GZldsrseGMzZOUtEpLbVr63gTClRUAcMP9499a8Pi2AaleKUyK/TTkglR5VqIGs8N7b
rzz7kD6iVNAFMQn+hHHANhDGwTQI77bmYx0nZOVDZQARvmFAMFE++mWdxi5LPZHke/tgFAtmC+pb
K6mDFrz4nl+CchaqRguEY/pwlw1uuPETHfiuXSGVoq3KLGD0bHExqCYrTstIL5R2CFIO9pUl4Uw7
DQrSpKjR4j9AsW2wI/BwX5jh94KsW/zU++ZIKzVFpTkqLmn7Q2PH9mWKchV8kaHz9S2v/s7AHVqY
3x6z+YkJSUXRlt/z1sGYaxhAuoj451gMXnOGL5spDDCR9Woy7xpRBBunaYvRiQ/xccdU0Hi4HiVN
KucFF46desyuO/P1y/uIT5A7vqMWqaJ1tNRSg/cViio+BDiHavOTkJSjonv+qJOeY99ZYJpqPpuL
ragnaIpT8qDE+cipcvWWzXlYRNQ1x27NQSK4gshECy/2QYpyn5e08d8WHW+1PLRPBX/CDP7Q4PR5
57rx0I8XwkScYrs2M/CK6fYYAxP6K8fFVArx+4CB3xIWiEVnCXgDcKLX562mh1KuQuazO9xfopRS
AccGEDLCuLvy8tz9zySd64f5fYjaOTf5o/5CZv52NtKejaLWuG+8F/A1tc8JNqr1XH/M+esNdu1F
A2go2Xti9QPUA5Q0lDQ98kEXF9udjKXddH6OCHI4vsVzHHlotbz2BHE8KSTD+BeHSW0GTjjzIOBf
vzyeo1sW9ZNbGMOKFqi+/AzTElRx+7Vx4NYiMuPwrsbLPUJS5MSeU+3NZuhallJ3Z/qOVReM4wy2
yLbaZDH8uv7LTBxU3EG0Etdpw4OBt2+61qPFFfufH6q+QF8+RrD/MvVoeq7QB7ZLmd7LlN2cBwXY
H+g3ZyC9e7izk0iZarMUgDV7lTF5yzuuxRORerWIMmfM9XFj2pR03tBS05Wu7IZftOAno531ktnJ
HPcPCCwmS5xeiExElxzeLlgEx+83u8qvK1V15yVezIDyBrMixr+S+OCT0kxGNT6cP+rnFBGoCIkR
tZd615F8gUfb0dijYCdSHoEt48nXZfAgqUrgj8q2ssyag9Et8u7guw66SvL631i9qpXYRac9ck+i
UomW1dVAF6qmtIa0XOGzXDZKyNVFVslCV9qvvQtplzZwdCMu/e3MfBn85Xovji8Oe/JdmjTJvJvz
29/I0FFdkfo51zqLfTuy8ZEp1yQB7tn4VvlmdrMKhXIsRBxmJ83qVfvs3b9sd6+rJLuD0eKE/GRd
NrTPIkS/tANfThm/5y2PeULl4zMDxPFkAUZIKYSNtzh7bKijDEIAs53Qy++y0midjyRFwB8TYwhj
mNm6tjT0y+sP3MPYkXbac4E6ovD3+SSkmldJZ0cEyjiPnrzJt2wgZwetbBveTTl1PmAXKu3tf2Oo
79poDiF4Ybr7KP9HR8vMg2/0rGt8X5AsbzyKbwrW9ZR6iZb4imj1pP2/HtpWLQu0wx1JwthOei6T
C6g60cLtF6i75RbaW4hdjJLpoOGzJEmirj0kTt9oqRBaBiaCocc0pmF6UP4LLSqSi9SaKaunX48S
RvrrY8INCXjnI5RtQhjqCj2CmzcLsdK+KAl99rOfDtc9Nd8CBsC/OOyZ4EQ8DEH2cNKPKjbpLjTK
gNHEWy4lYVstIhJVrn6TeVUwaanshVscLdxUeUUy/o0/5enhmUoNE7plPeyZF2QxLQSAZXVZB4bo
FeU1CHqJbaips1ccF2x9SbezfB6NPg7gldyFfcoBA4nCfFZ7I8PYWhdCk3y3TsDwvxo4EZKn6bXO
fjDhOn26DP+j7RvVUviTEW9S4Oa2iiICcQYyA44/myasVgpbegKXUrQQ6Vl3fE6kYcefBcjlFq4N
MnhxBJBsvok2tjx8gAuOPtjv7NX0MT6shWdLkhmTkOSa4KI/u959DtGkWeNXig/3RvQqKZ3I0Wbd
mhPadnjNO7/53r9Z6gzwSZGDfdus3QNZNZnhxUcWhLWmTs11Odae5k+dUQN5YCU7Go19OgKs+pQW
toCfrBBWl3F2Akt/g8GkMVwajqd3sA/9BA0ujMt0f1saFFl7Ey3IXjhRInMNJTDWhtukYhwmRM+k
ZB6EGC60lL/LsSlaBhHBenVOPkSDyRVZuaQserJvN92xrhNqxE6wpC92vsVMhdsKCsZDHWEczitG
yjYpv59SWd1bCF+F436bIUgoEnqkdVfy/8zu1nJstaiePzyDHcL1M/E8tmrxiIt8UBeC6TfJVvJ7
ZEsCxOJXOFd/EpRsuBZazLQ1YiN8HYIZYInwXj5DZEicc9MsaDcFaVkcAn9bZ6wjKQlkHHMvHRoW
0tMCKg/UtYjdgwxpVkrMRRe6UAyVrx/7ORHUgLd3yUmSP4EAKu+B/q7CAvm81k5a8ivilcrwj6/T
WEJ4TeHPKTtqcFKgih3ghkl3NYI0ZngVzQwIYaafEFQ6K0okmwAyxgOq2fBbTu4/d0O5TdDcPzgk
xzR1KVBAyRMIB3uNdCmUDKARz2FEVbTvFfXBEDSR86WLyDt/rNKBr7DU4O77+HZipcXvnbz1TdAK
eTjgwZIt3vkGupSRjDa3fOicfK4IDqVrhXRO1wWNKx4kpqn9OATl8euKOcwAKseQ/rWk6PpoJUPL
eAGfUTh5E+Zope3tmNQpfnBnD/15XAZd7QS2IMmcexmBruMIWrVpu9zH1/WqKxdAPQA4OoxG04LU
LbfYoLmycsjq6/8rM6HfCdEfXJf62bCtxxtdoW7CEBtTakNU+r19yi1jUpkALbbkx+RvfUT3pTZn
gern72mpC/Jh9Raj/wopPNW2VQ0mGWZV1Vx7H1vtLlEZ7GeSStNbGz1Cthd5sAM1zB01xfg3nDRx
UlwWoKNCKoyJDrjryETTJX8FBR7VDpZCkRYsskhU7PPTX1q/zZSL9tCGZkWPVgBVpBRXxDyHXsp9
jtwau9IlLquqajtwaiIh/zZ9G8KKKDRyl2sePd9Q3GfDeKeBbTctTSnRioPP1XaI1eXmtRbrqCpV
oivebosAGrnirVP7seXmknp8ovkYjYjpNemxkPOqquaxbN070nly3BmrGrh784T0mQldsG1xa2A5
artr/+YAfmICgUISV6wmUwReSrcTxl5pKw7jZqPtDolUEAdz8SnxAAMag5CpY+hxpMNdateRwJz7
tnToxdEFLz6Ro9PG3zuYmh+XNjeTXFAPEQTiAJVh7Sq78V7h652L8OvYC1tbr4IdMtJaFl3XyjN5
VVTzx/X0k/PM98RcQfZ0CvCZCQbCukF/pa4penbagUzP560JM7FT7TcOJpUpyDvDFJfiXaKK0/U4
y7whtJjwNhEK20GHcaSvmctKBe/fcxAITUQJzul7wTVG6YrwwBmPn3AhWeKV+cPjQZHFO8CYBrdB
y+bxAPPJbRT5pI3I4yHeFqflIfNIpAx1HG1pUyiWDEOC43K/T5MjOjpT0wftuIQhPLS4fc1c8V1p
ML58YINDssAo3AMnG3duqIydSAmyjuOtT3N02d9KzAtIZFNrCn7Iu4Tx+I/6R1trKQMb6iLlG/Hk
VW6u+5vityFD1sZMjd4AmUmRy7Eq6UIwAtiomV+xUjjtLbNH9tyENKbOTmX8e9N4jWMQxmXxbuTz
vCMKHH5+Z8kcvGSS+pvNEOtAPj0mB2F3f9RZgtE5zDavalUpAaOu7Bpho1ygfW+WaoQPrHi++5zg
ReGw0eF04MPScba7/r8plcVB+q2DBk4SHu4l60a6Dk7oW2asxCqv6wLm7UTIdNe1tBdtAOk9z9dz
ieDEEP1v76tb5WZwMG3zL6gTjs4v3x7r8AD1Mj5P/Fqgm8KxCXCXmAGZOmbJAXJjjv1uXhHXtT6q
w3FG+cS8ucCOEXuMtMKWj+JXAcqXkjpoK0DFo5R9MkDxT8iPgaQsR60MDYRAq7AKWMVvzVtWJBxh
tmTLXVuc3Bsf4ZYzIpR7K0D8fnl+QyWItLWRkAgIkSN5xA2kropD7ocxSVCg66Hx8kbyb8gm4EKA
yemhaAzLWaX49Q86LpGbhbHAN2u33bMGwM/s0LRTLdBIWCBwQlLcLKOQtlbqmLQKrcSr5Wwd6Vq1
ZQOd2uLbCQEEJtRSiXdmjdhEWX3c1xRBprbb2af4SM1oS9KZDlC8V/CyvUqUVRsEdeXTUsCI+BAC
nBi9YEHEBLCkcPW5s5P6Gz3m63xa8E7H+1Llx6yl32NgUuiHpfCmT9sACyN+RlG5/ObaxTykLoOd
yhC7Tha5nZ6zORoorthlNn7aHW2uq8XfWf1AWX1cQ0jbv9kkk6U0mKO/NK1CecMRHLr1djKX1pcj
Xbu1d2iHOqTCoHcgOQBd5C6n/RuFZFer91A2L29nrldEBtaPSsXOUYJ54yZK+AJIEgj9WX4g+A8X
NbjNlR7psmfeRZChFPPJBNJto0+5uwwymtEhfKRoM6PwUxu41D8iT2h5EcyGJ0LR3xrpRhy+33jg
y9Y4D4k27vcPkYwkk8+JrQqcaHTO46KjKoYLhFG4nj0a7/weQRHilAqBxyKdtkTugAcjuzmwxe6o
G9D4yVm+nhs3qmryGmjHlxv9Ezz8xR8+AEr3QE4geyiVzp6tjbG4kn26UxW+BMw2f3k5wvDt0N6c
iiJ60S8LGpWdV+3vYClKxBZ2opnwPZRXKjZhnY90f+HuW1YEfqIDdJsx7NcPHQZPfx/29v85YY2t
4T/ch/KIXd/l1PXmh6dtgg6RuSThdjJ5YQ/1xwcaMZsmGjmuVYnhHunsUvreO6sHhQdFqS6awMFD
a0AWpauL7kEwRcvheebuNwk57KzHitQOpzasRLKOe+ZArLKU+/QtJd+sb8Sg/iwDAVAvkWXksaeT
xYYjON3uOfDXr1kkOH5evr6yPE3XmsIhkAoNbGUtAlR4spJbdUgiBaqL3sjfgD2/dyzJKlsWdLlf
YiUSR7qo3To8oSG2RGlJBtXQYv6NwEIUeBkKsJwt1FtQ9wiErE5Jrhm+oE+a7sSda/0zeL+2OERP
ttEEZck26XdnHvBMW4dG2CVmulunMfeg2Am0nSY+0p7M6uslpU70pE711/cXexMl7Lsct9NAd5J7
BPG/xgEHVBqsCCG0ON+gPptPbhJQ4VJDa/kYuYp7EJVTfunQLyjYa2eGt0EjT7NetGzNTNOVgwnE
s7VXr99K+OCeBaxIePuSRIW1g+Piiu+15PJ83i7atLe6cbcUTi0N2TP6OHyXWydYjw1QsE0rO0A1
bcqeFGVWUukVkI32dfrsQcG13XL79NX2PwT5l3F29X7zDyeQ4A++XSrY9YxhtpA5BbZSjqNFSsmB
mJcTel3L4os2oy6BKMKIWUo86Vg+57XQG64HVJCzPE3h2wAC+xZMxLA9N9lu8ez7W7D5TIesK9M7
2r/s5iKykHMdaTQuOemWj3URElIi5oIs9RH3JTSUqWHZtpZTZH7o1RTzS2uRk+yumsOYIQpwKjIb
o4RRj6Iycl24sbnD1GLC+kBZKg7LeQ6r2uv6SaF/GUlaINBwpPMXplExGE7tzjuI6NnI+SlJxKzt
+pg98QYIxwlap567m+IHkTeQ0aWZR7PYmolORhpUkoPZMIIoLd/2kAwyDwOkrmwQ3WW/jiD9Nh4x
oEghpujvGMga8GCVn8qvIUzzWCRG/SHxJqu6Qd6QVzTGToCHCgcE//reDp2K+lI0M2SPQSTgYmG8
ubbfvjqKbOhPPZHC5ZobppI6uxXTDWLQlYy1/zknbTJl/ZwuYBzv1Ux9N1Lp2eed9WXEAzaRCeUO
Y0dT/T/S8ggTTErJaM2ST8wv1UDeh2kg6c3PMFtonkdOfgA37xZV3z1fNCI8AKCKekH6GUP+7IRc
Z3UoaY9n3ffzmkBT7CCySaOVR/kFsb7VIqNH8a5CXu6RBf6puiqwTPhEoSpadgB9yfPEfSlLEdPU
cmij1h8/YBD+XQOFSZ+KJmMsRiSn9M0uYYs0w4ffmFuFs7mK9S0ur9h6DVA7JpMNjs9WxGxwOpik
06fX2g7YMnVN/pwbMoQ3ktbiNT+IGDNSp7gZa2cRs5Jv777f7kEp5Lg0FS5fV7sbjNFJLNxne4Vs
Zw9OeKfbo33UykrASCg2ZlCXZu0lPkcVu5eW96otnqG2WSHaGuzgtVKSkKUQGfomAvrT3EkkjfRv
38FQ/+MvsncbLnqM7Ybg9HgoUNquY563+7PIKeDXaiJRAfarO9ClFvbxhTXr3GqF1PTNunWUSRQ+
Nv5inCQDW7FkmWlLO0y0eFDJ5fxlHx6t8kDcFQLv2dLIzYTLYUPLHeRc/e238pKjonfO9msSEup0
B5t4bcd2vtQsO0LtzNammy/Ev6DgL8pvwRKQoAla8SvNbXEFAQRzvy5aBrR4TirjK1q0wHs/tx1z
EcOGsJ+aEP7Cxk+IIoHTySeUBm/PKkiQ+ir0+bFzP/W1niivrukp188S6an4ywSg5RFzkxpWR+rI
fipYiOVSy+YBQHAO8kAc8aX8MsePvxlPEsOuSC2h7OSLwTZIVJCO5Fee+c/ggR75uD8UateXJAOQ
GKjjeR7OuzzlX+eMAxS4FJUPcTGWYrDA8yzrFAGznTLDXx2Y9s8aqL50WrKWD0ZIdpzlxeXh0ze8
ATrNa1q2ny+p2PtsNTaIZuuqMfmqnqa5SNJh+62mTrBqML3orpqFJFnGPZWJ60VA+/9i1Sni4Q/q
vWmt+8JftXPxBk/Ej6QPq+R6Vr3o+gvEqIci34gWfjfsrzNbm/5ekByl0WiV2hCxBluhban1H+Om
6jBR9cljWtU2+ASpHDHfufG9+UbP9hm9UEFx3lhiS6tLjEagAGEqpEe0Y5BOk6gsA8ex95Vs9K8t
9GYsW3E0vHKGYYos8VTrv6qT0QStE8R5P9gm9IQvb7w9IQCQqdVMGVzhgJIwma2927dR3CXyWpvq
24k8nrpYTqHFc/7m3FSx2b2xrZOrMhKZmDRp51koK5h6V9S9D8NY3LcnC3BIdVKNw4lJmBdme82k
okBvOBVwo6hGxW8nGD8GOaQV87Z1DPQVbYEtYEG53mL5AlP+f4lCIJUpdWNFDBpA9CynYJKJPIk3
fMv9WVFzcCzw2vLq+3wlP5O26/x+GbdjjV1N7b09RF/mhvYCLj7IqGC1k813a7bbAZH0PfDNqI01
qUpw/bts0+fVlvtZm23uEMGFCfCJYqMQhmbcm9Hj4V9z7SQ1v1SEm0Juuefyy/ZFFfkHKF/dJfrp
h7gEN1XW7LAd22Bm+hXtpynM19nrCcHSOousE5zu3JXJ91I7FeRraKCeO0vOPDa7wSxO4sOFzACd
QAxj1NJQvLsBt77lPb7zbDSs3ag5T4+Rwclkg0jIBcUbqb0w4fJGvCxbspfFabyfjBVJ/e7bijFj
i2gRIiog6SvD7XhmFKBy5PRXxB89lH4YaNRyHqfMtmnjFMV57eV0Qg7YXT66ODVowY5tccscTfHv
TSKbiaHGpBtSx6hOmRzqD2dCzvCtzr6gQNBqWPI4f+cvgZzTLoWW6hd7uZMb8tdwd7GOD6Vht1pK
YpqE3OcAUlCcnA+f7G4z9d/Tm5C478UTjhkW9C3GIZ308DBMp5L59URrQPxHLP419VpYEE2+Q6Ej
nXIdqfGp5nXPxLEI1cZA3/9QAII1OuylOc4sxsulcAkw9vIp7u07R0NY34qvmBcejs5gOqxjs/Y7
szeGUinUfSjp18BXWLHzTq7/W7VJgRILih9oImXHt3XgUZjha5TpXLVYTDpNmg6RNJN95vlLQ0Jp
VMVEZ2hMenXr0PG+70GMeEfAu+TgbvWbMdhnTtvXsL7YUNBsXiVIpCkffz7FzGqFp7jC52s+rWke
iMveA1gPMw+ng2HQReEOfpA5R4cgLJg19RsWHvsAQMB8B6hbSjlRy7n9s1pLwS6M3ipUeTb6+eTi
grAm5xa8WDIOm3GH44MiqzQppFRqmB+Yw/tpxgza+7DmFrMBszZmxCkVhuqlsK1IHipU5t4SctP/
2qXJOh/Xb6LPsjORB+4srK1Pbw9jV052541Jcn/mF+YObz9aqsv/7jFouILYI4pqrhE/fqrvN7yk
ewA7IYXpUceJBckNqkcZ0S+GAbcvKrsRxdA1t4ALjglmjiEdbal83Ewn/kL7G4LZOLRexacbjKR5
XMNzP9qOHUgE4Ayg9A/hSkVRux6fD32HVCvtZmbprdFAUngR36z/S1KlARWRoX2ymRjcbX+FuqgX
ONbMJFKlFrkwZBVeYat5ElRVFv1/M+yor26TaC6UZMBCQKXMwyGBP2eqmtgSc/yArtl8enmFV5v4
i2MFlo4B0pejcLjsB4FdpeX1w4aN1jYOi7y5nlU8DkkqsLeb8a9XgPNzCFmjuk2vlimVTTrjiQy/
ZJUA8LApdxZ5bdazuLevKC5GuZeskIIFCku/8vXKNdPRfim2+xYTzQB82IKdkgajgK0il1JV3Umf
hkr6Sl8SDCbb4puRgDu7yBet4nyTrlI9Z+Hwha8yBXS2D2q95fKSQl4DhBuzpzgH6/jwhn8QDpth
MDgHa5GaDTNzLAHQKlPHVX/2Oix18cDLZ09iuxocviFPY8VHbzFzUfhcpKeVBD+c6Bs460psiUKd
qe2wQ5bL/l98dWqyJAzua8LVsN5gl7GGccYoZAi/QP24XXIB0dlkQkM2XNOrMKTAg4cUF8dzo56g
J+ARsRByRz7K7woFpap6xPdPboOly5TpiiHQDThbIl4MAW74NlV4C4iYLuo9+d3UUoalvr/DeIf5
+22qZHQdhynt44vdQNpLQvxxkjuj7wkwAB6dUMKv7IRGFHjSUC7zia+7UKlBeGMOGLeFZg3/bA5Z
qzNdp2eiDO8XQ836CZbBjOvM6Z+eDKTUd6cuWFPDAhSA1CojfrbpT7jfeXatbQjLWEBlG4IDc+qs
bThC/RoxaY46QNfs+r3ssxnhK0nrLXy0OxBGiqIdMv2FUWJHaHHxOy54Iw5lRGLl3GGo5XToLupv
iPr8WhlS7ksGYk7DlAS1aylB3IJjKbp9HkImmxKXcoYW1OLvhD4MF/3KD1VuQzgd5c8pPo2ENdxp
KrKCK4nDZY9HXLeMYLEQjzzM5EJizlOpRijT8yOQWrDcxfQoQ/yNg1UbQJgIAJ6+C5Jdt2PZ1Uka
PjlV3jkfWbvuRJOs9zw6q+fcCK/TM73Hs90NotjecGFynGcfgapuUOOEV+O/xJDPvAULfhFGbD+u
/9I0uwoQ3QkCrJNsvLhALLY8zCJFeKBu/5wKmm6pnxuAv4cXCujhK4ku+TIYNn5Gk0MPJ8RLZknc
vO0Z5euzS7BART4C1C7YZ+m5rxnp7Ci0KJsuSx0AYtBGIh4f2O8nGD/kjWheIHQ1i2+35IQKb+Bo
`pragma protect end_protected
