// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:36 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
ey9SHXPa+uFgtdgQv//27gy1rmp7ZyaY5w1wDJdCbwTOqSFRqzQCRiydmH058Qjl
o5Nx7fcbB2ZPPPdy93G2ra/xgHyzNaAgVqJhmJHtMJZiNoX6PX5VMbdK6G7HAXPH
A+x1ttbyde+qC99enf/oMmhjdTDpK+5evKqD3o6eSGE=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 7280)
DjNjI6xXVrgmhCGpp9OuS48LmY9M+l+Jlzz8Yx6WpU2OHl80XLWG4QxALncWj7l+
IQcuabMba0yeSsfqlzmq7QLrVK6HRjk+TdZc7OBLgteW4v3rl+s//2ujiozDkHNv
GAG6dIU7vQlr4ZV3wOTsj4lnbLAPHM0p3U0flKLZ4NJfEhksLq4caT2WEZVP2r7U
+fYHKYbcPF/B2S/hXjOBGwI6iQNTfztX8pvljJqDYKUv3jowFAnbC4RsC4xndfOD
m7VLL+K6LzL0fcuMYPI2jpfH5vZ/JTNBvh6L+Lp3boOKTwH/mCSfi3n013KSwT7V
qot9cwDJxBLrIEpvxOqQbsXHIk393bwmXEjNDgLZWMdLUY8xfwz/SOagMDgCwehc
Ppb1XYFpyWKnP7fxbno+f/YqV+Km4QlQd9jhA64i/O09yWQF+CeuBfJwFpL8Orjj
+rB8FS+PJWCVrcT/FI7mU1qNPmWD1pGPxJYSAB17H+gle/XFWMKVxeNgFfp5JoMP
i0neeP43e1XP0pmzsDuxiUDJGcz6AL7ZU3DqQJPFyvcZTTwPSagpkyrZ2Mh/yZCz
pAm6lqEYpHKQLz1H1SjtjR0B3+PLP/dQ8EEBRqim3nOGmZACcOQ0t7VNogUaI1Vv
ToQEZDoXcv0M7jmkOVsVXvhH8d4WKuB+bn+oBmKxFE+syq6BCaMsQIAjmdCMKayn
D5ZBLU48XGzoXOjsHi9t5vAHf4FjeINtmu/hTyJ8OymSOHvGW99suG3IW2eun+WH
UIn83WTXhLFxdSS8Zd+Z7ape1uMnbp1v+DKwBfnIOSdeIE3fEkQIInictFr7c1rS
zstr6r3S3dSPv0ZdAxyHksWGPiZKDGlX3OKHty+uZW+tfLXJty2hv85W2El7X027
/xF0MN6fO6/NEHFuT71Sf/bJag+Du2DNODPZYd3J2RurUM5ajIPaIrYjZMn0WmXm
uF/PZW0fQ3UY39J2bPEY8i8PkylPfCCq5Hzb+69gao7mY4zCOFZOQQ5Rg1DyakqR
RS37sejP3HcrGFdi2Wos3ErC+f7W05OdGy8djhcHYGxwWu6dAtJ4lqKD2mdR7jOB
EcxWmBX0vnzghLGfZBj8GuQwTqzd20CHM4soCL/ZUHsAj76ii19aR3658SkTvffP
TAn7YnW9ZyivBbipiVoTrG7lmwogG9AbvvDtYq/3jSOpiuacdS6xgiTJiJyMPNez
2Eaq3u/lcMF61iHGFfMUVHMiENEGLCGngrDB5HO7a3fq74y4PJU+IoUrdGYsB9JK
ZreCwypkXl5RAjZGC82t1Tm5dbtF7BpbR9/NVttDDGKdt2DXqjzQgNlSUJq+/jGc
ewyXUGp+AXKjXejooZYqnTiYYplmzWwCgOPmw9I+QAbu7UW/jn0yn4Vb4a074uqJ
cuGTG27oYBpIdi+mFYN6zFN7IrreeI2QvaBwpjVuwfZTMnahkuTyhoxe8+Ktunlf
pVhBdu0TuokxfjRbdfge5yptgrQq7nscB069IxqqbKHaboqmk35O1x6ccXJZ6ceP
IwTyntJqKnB4eO2O5E17zypmussZK5AJlrKqSqwEZKZ6ge5gUp9gPsB58YL79JC5
cohIm78oY/QW9hGmkImcXWTz0WcP82z65vD6VKDBeZsF0U9MUM4C0V1rzusrwNqC
es+7aGKiLpxuFgF/X9JYnnUokOEqM5TcFOrakaYa6japuXjO+52KItJMEPKR4Jgs
T0qQStS/dTlNNfuthVWoTxD5sWROoPbkn6zjoj+uDSl4jJyeaiyVPSHT5r25Qtz8
LOiowGeWbHVQlprhEkVCsU6Fv9EtDUdAy45ItqZmc946dARhjIViPs8PTfvZ3oEp
Av0nej53nW2Eji3m3yrxdBsh8PQEP2200jGJfFYvDHBAhZFW4dqEsHpwm7czmmkQ
rKQ+nmM99GoZCmGCCQIZYjjMUalcW5taMDpvuCXhE5lIZQ2gFbttqSUYQ0h5GDWZ
0s5qnJtBBBxXzrXCRr/tKmXCPWLG3JVtrQAz9pTHBFF+xrvscXTa2n1klMwVpbe6
23j8c6l3xh24J7beCMG7f7HMFRmkzQTWbPGRfaA+u65VEQeNcuNy1hPCX/8NUM4F
ZAxs5RJVRsFRkFjmWJmN/Qh0TQ+aotHHkGZAsLwJW6nGEQNXNvQI+5hCS3P2E0LO
Bm3i8goQzyPKm8j5mudZdRGnkdioJV+NqCLd2QIfD8LwBcMKo6zPB8fwrABnr9g6
7OGrndSrdBZ7W6xYYfK0iQUenY4YM7vB5n0NQNBrEs4kf7w/RMLCgpVSPdolpoQF
dlFYcqJ3lqdg1qA/dr+P2v//TFIgvP0a90Ul7vPCeMJgu7z6/bekbvj3qq34M19R
WC2JHDGXaTFdzovhziumQmJ9zxG8O5Hyo9HlysK7A/Y+FOG+/EiQuJjBs+kpc42s
qjnRsGsS7+9bDF/f7cbwvVYJvYr7BMhXMQt+Xf92Zml3uLXlrGpow5VMQY9EMWRm
MutrGqKJ/iVIu5/NqN/7Wbt+FIPycozeTL5YxY+2bqSIbY14Z3AA4AypcGN8eaWs
vNVHaSzw2GFqEWAqL/Be0TvH75SJ2lV3Hpm31knipv3WZyzJUcKNE7VQyZOE63tP
UB+c9n5n+KJehw16LWYHAlHJEcwprfVit/jfB7CrXa8aBgYg9EOgXBEKXZJvuY9x
1AG9PddZ9mm4qvNXOxHe58VYraWKeT0h+YrTpzRn1pYww2F3TZFpWhoqHL0g5ylU
V7gTwaUHDtz0xvj8Jr4O3XuCzcgnOXjOtC6f1yMpuwH4AhflohxsjDj+yiZLRWBK
3PqfD0H6p3pyggBx5UqijIxRtqM88FsrgDO3uHBhdYk+1rzwos3Suv3AGeMvVeMy
H+oH65oSWKdmCeretQFvVMIXMl7D960PdWJM6qYUE57S3VbBrMM+eZcmzPtPJKJA
z83D/A3t6aXWKQDfAzX43SENZppaa2FJcZXKzPNJas8gWn0IA8JCivj/C5YqCAgH
FrSxrTKA8wYRF+gp5uv+JZErdWzj56cFf6bTi++92ne/FOOYBxlQmIM6B2o8Y651
LrGzJnqlLETB0d1RZ2oerPTYu+ZudKY5C+FpsfLE0APh2uOhvsY6TulfH0L1nvq9
uMyFAmnx92RMWQb/KubAzIa+l0dVqrVJ5yu/o1C3EBfcU5aAngoaAJCSS3PDGtg7
sft2DJtq+Z8fncdPiWkL5vfaJcGq+FK/TxpSukuPQNFwwwGDe/Ulieo5ubNkrzJo
5oNIjcrHg4q7rLewj2QcjCAzcmUfBOyqDK0DtQy5pwuZMfgkYlj8NPCJjajAWs3E
QjUeviXATFrEfreKXput1Y+9D+gjDq8Yl2bE8YAaeAGfAPjQI+yODLB3IikDunA4
UrJDvDazFqdKdK64+mdrLFMQFYhjpoXV9Wt6/2e6cvil3+PeuACSHXgGV+umJBIi
TREypzaTR/82ldVMF6Hk/dCu+8WMba8/2rT0BgjF6HoIXOFwhZzTvxTDbGN2Li+E
VvR2RgwTnXUwctW/1tTgGZyVzZyb7jRPD1AYrv0xntph1V7QpNjopozQxnXToyo3
YqLVq5sPp2ap8VObI9niYTarnCHOXfZ9z5WCXGbm/TopYfqm73kpSERGyhEHy3IF
2tuBeS1tay6ztu6aGANz23ctMndWOxyn2EATw2PO/wm9DanALP2vpYTcQCMzgxXC
G6zCjHmBjKk2MdfPdTUbc7MNmsxOji0i7wuE5tuJpkcgMtZYlk7NdMkPJ+WOGkDP
vxJhLi3VgnhPUxVf0BI8GGi2P01B7yUqjZZ/qcqcHEC2AOu+l+hdqk5mZ8XZAdGQ
nOjwb7/UuFHH2F5PLwDA5KB2W3YvNJrH17iLzYoIx3XUAAlvjnPE4nphBBoEP1U/
/EDE6mCZoGl80zfdqO4ljugoOZWcJbnh/vyiLSe8TaiUzYwWfM2y0H5iYDWmy7bM
W+xIxi9JPXydiyEhboBNZOZWEUvwZts5dl6H+rKNFDXp+u+mXyfydqz6HCKyRqet
quPFZf9nxWinorFbjKifh01alY9DtrnbPcQB5yaDrk+2efxy9G+hXaJxw3V0aIY/
kf+crGjoHEWFApvTPKk6PEAKKRpPvDPv86hhGV5xbf/LndPFPlu8KdzZ3uapIorA
d7nAt/BAfRMCjFaAiwtbfNyiBSy0AyZBRWZ8od/3pEmzXu41Ecu41MqxwlgGGUwa
H4ZLVG8m6bKAeXgM/qCQ6oykSvmbwxc+ch46HlG4vDMQXGLoYSRdRNzAhGMr0kXH
Ua4yucTHwk6n+o6TcLNrwVtV9dBKARsaFJGtMJGxbfXKypPsScKu6x+jKXt0IdjD
clUXAA5KUOgPY83P3ZpC42ryr7EpCpRAwcoiI3aDzABgt2vPZtJRcIs6C/3WiHyY
xo16SMZOQHXbSHvzQQoS6bO7TrEtRR4pv//vEeyAnPX+/T7ucgVMi/xkBuNUCuNG
0LbfdM7Yjng9+Xli0Mp7gnOgW2ntCdoX94JdrXdK4akcGtlkZVAONZtY/pEFcYOu
fbkdcj24jR3+pwsikQahEkeAz8qis87ijH8DG9uWuR7OU3o07OMhAwJzobYS9SYF
OV+ZABlGR6mwMe7Fr+0UBZu4IGmmVVYnYFIJ6nmRl/nkkGKSGYmGs/WDRa+EyQJS
eUTMNW8WNIGge8SKeJI7vF6tnlkT6JRQkAOStc7HgAOI6up8FDmzepbzR8gcu3m3
RVnGjq8C3fCI/d+5afiA2tyQM559lKM4uTMD44o3OSNYs1rBq3xgIBRE1WpFmT/e
MN+mk1zupT2xu2i1zZ40MxrhPBMuzSk8jBJyqibGTb3MNqFKLHC94vSVK78HjmAX
PvxPUfx9hvl/HY2V4a/FxqmSCc3erXCa2nxKgKvl78Tp4/u8USHErRf/X1l8omA0
xhWlIiFExsdnm38y7b8mJSg+FcxBHEMtr7SRi2qq9kv/56fonOik5qkIKJvVbr2P
f3HXUJC9Kc5XeyTCgrK44OOWIVo8I5CxtQ5tR+O1MCV4Ni4AIcmNf42hIlNMDqPk
lMWf12wPhbXilSGWQ+LyX3AR/pQ44sxenXIGvselz10URE1dBPZfzINedPzt9BYX
zzvpbxaRhUjaRHIpSBLJMUv+bo/IdNjpdO0VYdNST5+FQ/eCcA2c6wuOEFCQIp2g
xUg2nGi/HM6XrkeOpIj7QA7ukDbkPduVM2OgzJXNU8ieKy+fV9QJHZUTe3ZvbWIe
7h2H7hMLo7Cmhm7xJ4gz80KhrAF9AW5YkG09X9SOQ/f1gvyi679uq928AxWs9Dv+
8jynTfFME9WIstUxakVeo2VPS75mlqgyR9aG0cBrbjwKlVEVmEOmXnmT4j9A7atZ
xbY6vBWNk0I8KLxWTPuJq/mLCHrL+YvclP5zJMHtHzTQl7pf81NGdiiZLAbhabco
9alBWe/vxwzfynifNEbC0C+ztnVhC9MDkFAagN88fPJc9VTm46+Lcfsw4YFffB9r
x+CKfK2SVEIErxXzQ7pbAKAg5TyaerfBCMKOSceICCXUPEZbyZu7mXweh4NURvGd
O7KbPhdHODH81VTN/UshvqelVpGXbwCVYTB+8dVomBM0m5iAPcWaP09WADbpnlLW
qzB2Sc3URYlpcdVFUzVheDj3123YJohLDbsbXl3XCoeegfKjrzJHhnJHkHfKzFoE
Hw9D2FiL+s0zyDbXlWBryjcFPasKDbkfWG2r6ltvvU2ekYebxSnneqCikfXOZEfM
nleb/FlXNrucBYBP5MG2IXOgHxDNF3TEsTknqYHS2cr1k4zkA1a4Q0KRwVSdMQGy
xefinhBiG/s9FjeVMbuikLZSyrcOblXu7wXSEOuiw38yiW/4n3zPYdI0+KWcCks7
YCA+zwvYWRq1kKPV2v0ELnk1bRlL0QkS99X0MuR0yz2pUu1lfsz4/bOEPZRp93+f
8d045hfN9muvTyOrece2rVuJmSftrwQAYGFcG7YDjSjUXv93vyICptLZFdth4Gka
n7IsIEd6dtG2ezf+sEakNmZI1RS5g4aLGscDVDYrmbXFkrcVtnWIqCqpkhxbAHZj
mOMPiVUrpw1wt2o0W+Fkb2Xn5QDgQc1fv9ChCjrln448Hn6eCQzhSqHPOg5BXPFc
CDHYFbgOCTgTHy5wPwu+r/iStnsoNAvL0Bjs4OJh1LDHPUiid23lp6IRwas+9g7S
T5diKthYx7+YLBWBBRcoLFDEc0tEnT/vM9xrTVERB23Bpo3Ia0kGxiBm017sFaqJ
EHoUcp6L8KuU4gdAT7NIWdw5lc/OX1HcIcldzX38BD4UkUv45QvigjJVvzV/4ib5
+554KNUq1o+FbwllEjMviwc8FlDW3uTjsWVPKhyBXAA5JTBOBpz7VcHXl+kYFmiG
LUYDyKk4VYJbRg80J64sAxWlEW2YxNt4zHjIZ6FUlw2h6wz1So9IEtqilXSDVLsw
Z4y3HnkBj2HY/cpScJCRmSB++8epPmE1U8J5o/TiboMSX3ktrqRTZVTeou0JvqjE
i+KBNKELD35MqN8oYIdL0wY+4VPJRVNsPbKkRbnR7p1SGMTxhZlk6lCdpTumHkyv
qZA+gz/sUFXAnQa2bZsweYGj6A6q0Q+1nkoFg3FOZbrjhGJmK6Hd2KjwQ0W5jcJY
qZ575E1eb8onTd8ZQEkv3EfI4rbKtKHQ0Sp2WYkWsPij7/uHIlqmJvV9icf2ilWS
UetWwYoRAdWEyeMyi3xkJWYymhqXqqdGadHWIWg7gG5yukUMp9pajoa7jb3hX44f
mld3p+oeJeV8tUDCO1aQrqoe62kwg2dpeAm5d0vkUz4eyrLbbjmN3SHDbYnyLE7o
ZEX9msxT6DmrGKrnNLRAlZThmx+VY0fvyCcpe0GlweqHrd2inU79FGk5dslSYC7x
SZ+WCHGs3myTlE3iY/iTCs/mx50+TN5ifgnZ2I1NWDri0UK6O1I6ryEk/PsznFVq
j4S2+BsQmPg8faXN7U/NPCzhF77VjUDPHGUq2hJat8E+KXMGRTvxiwrffNm5H2CS
V+nc8VAfIR8daJOT6kd17Vg+kkSN9dPEtek6zPE/7n3qxwy0484hn/31EhpQw4WU
Jkm/CUT10dniH338n0zOJn9soY7f7EeHv3KB9EOXXDZMW3sYPavyIcCZ/pGHi2mt
fb8J+v4N1H42/Pp+sGFi41ZnGMbp4QxkTy9mLOlIMf5fSwuXLiB/TLdRfOX6h6es
ndRvGrgLdW7Kpfb39PJTS5AJKc7HMImF3Vewtp3xszj2SuSM//hfkWaj58+fJLS4
30azZ/XcU+FIQDTg3m7p/i6LNV1xaaRdcWZfKVGyoX+EfpXaS3BRz0HEPJ8KP+i3
/QJbSdbg9iaZX+p1gqnfLuNq4CZysQxZkr/FUPxDwllEkmtu9EUzfxYMuTjhdUAn
9kenArF5atWZUpvzajsE5+Yo+lREsfHULceAel685x/6MSMvHs19X7erJ3IuQ17c
SxNvTmyIKCqcPMTLxBR9/uKnJYLdE0dO2Cyrbwd4UyVkRwMly+XGBiBMjhSkr/ZI
dYJbSyCivF/UQ/zR6GDzEp4HnxuOgBa+z9V69Zz4coekTAIZRbyD9Ywz8IHPj28j
k97VPG5OiJjZh5En5a+e/5xSDlQzeK4857SO5z3X3W5j5ue0p+qeftM0KBYyqot1
9238qI/GrRs4tyEqObeCoWbcrPG4FVIuIPZB3MUVoYk4/Ga4dgMxkF/YFE+usYVN
sJK03z9vWF1kVdYz/eZsqMsu4mdogyoqeMehHIWpEWqvfjgW/NosgshWDcmqL361
GXtbhtXNKOFJxGF8UquwSWj6g5yhX2ExVSiWvk7p6Y8Y6VeClz8h6xPBNhfiogek
GgEITNdONrEr9Lvhx80P+HhLzPwAYtVlzmFpw8FZex9ErsQG8Esl1SN6uHqujOob
vFg/jN+8TfYQ8XcVO9boPjgyAuPGss7Grx63COFu8lvRrrBYJyCMM8G0tAMFBj8g
X4+q4vp92AHFXjGfRJEjNx1c80BtXhjRsbLERSwFTc+ifhw7I7uYsCu3gMpf8FPV
Ubb4GeSARyzRVMD+ecUTpKafTvx3S7/IvtyBHQXNtAW8wzP8mwyKWnmRSSzA+iiD
ok3x3Ctmyh5VVxbeo0cV62WvwQzpnYimMCHkiGL0i1hkVx5fAdseHDupcXdSq/us
sKvs8nkYLMRuCHa1I35/zd8eJXFCFWTTIBjjuvDurd8xyd6e3K53lIcov5573yG2
c9QRsAWP0khpYeUrESwohr5PpH5fxsc1TUXjvmoy1ydct9woNtEn+R4ccwqtTLpG
7bLKTuJadxK8MxtUqsMb6prxbSvFOqxBsTLANoEYQnK85L55hebIiaOu16lwTH9o
dDgVkl5Qjrr0wcJLtiZJ/HbyiS65legcnpmnsHFcKjYep1pb8TbnsywIOLgdZbnR
8DBnRZ9gaP8Ll7cBeUjBIfNXtJJ4EtnhdI8VDzo6LRkGgyt50z5jmd3RX1rQNIzh
eMiUdUM+uHNL/qjnfJlb8R96iGQWTOFEfnhBKiR1c72vv6DbErSFlvv7eQBEI9/k
7NiUpwblKobQXHIliW7CqvR+NEKSHGsz0ulu/Wpi7+Zd6gm8im7kkES8xAkEcNRF
1msqvsKO2QLHuxH8pHVe1dcuFnmtof9uSBMfWbPTXvAX4EqAcFwvioLaRVlHVSCJ
KhEEJjQKwhkH7rbbDS3xWkHvJ/KyMMQbvXF0x1UXS70COEvlYzRB6lCAByl5UwjU
Cf6QqwhJQ04nVlJWY6KU5dI7B2APyJDwSsj9hiqeBNkfLL5Z+fwGdBoKb5f4CfJW
AlnvOmXFSaM4IzMw7W964X7vV+4LDUDunZGSlaCdWL/DNDJ+VfKcHHWdAUkBdPly
4/TWZIceUPnAzJXaU/vOz8g/uOQvOTM/8X0dYy1YSTD4SgD6ppn4TH7m7d4VO415
h2q+IhYx5Kw81dqcwrGExnTkFTgo41YYkLgg3uJPoaj8IXzO2vasIWjBjN10TDlX
Vl6BMNENLroSiB6kV7TjCDvaIUnsuu3IMrQA8N4A6kkjvuTHwQAHx8ozCql43Q1c
CKy4Yv6pKENJjH9a3Rxc+uXJxyCIJzEU3P/pL3gBpH1Cs4jDDiXf92J2voQ8YSIb
F/WbBE5U1xPAtaVDFCw3qvDu1kwBRyHcPSXZgahmp/XdLexwvyCsww3vUy4kXfBo
w6ST3m985FcF2g/8o4joUcVcKADSUdVE5CIgFQaVGnvHKH6r0sqg+XY4F9kH3o4o
RdZ388Lg42FmI9c8lJPm5SmDWjEgAtjEMw3S+wLw7y7bftPITfDPHoo0qW3LDE24
1Zd7Li4FbfrtpOjlKyBaKCzFfBTSE5BC9rZ69OBl2wIPMNy5c0+ZJsInRXjUkTIN
Pw8KJz2gw6gvpbrHRBUF3LPzKEfgTKwvooSVXUlcnABc9wfme5U7dNbbM73cbQME
QyZSisQArmmW6ZcCMsi4at02bj1PFCcARHYoLfgySTo8eY+zqICgzLeeJ7YgCh3b
NEynGCDeQhYClLPCa9rHwweFJ2hYAKQg8DHO1WJBSCrcKxVSnFBThqJvsSrlol/a
mWpALikBdXEGk7lqNIJkkr2SxkfSM0lr/zyGfzEBfMD9QsdXN5NvU0bFzgMs7zjp
ASILs6kKFw1pKBqll14ruXleDJz2/KxVVorItb4OHBk=
`pragma protect end_protected
