// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:44 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
nV0BKNO/auaottHY8BoY8iucJr1kwMPFi4jnjbunATiiAZmUMvpKNn7AmAakSgqt
EsxTKzOmJMXbxOwL7WaXicvfyTc882zTSIl5kGKTUTIujc7RfMpkO30KaaWpW3ab
x/dEYEdNbHlP0j2E0JKBLNkhzowmQ3nevY70jXP60Ac=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 28000)
MlCwLfi3y0Nuarx892KI3MUlmKpNfy0keJRp5fU5WQHzWRC1pOWoIBjif8I2D5ts
OqxEr5/jkbeMb9MP6ORC12kskW+qonJIlRKim9V0RuyvIHrQdOzK5xPHibUxatHc
y4RHEt24JTgDMhxRJSCHJDnQYACLFB51eK9h7J/XNFM5ypCGZrKYvU7G5E1iiyRb
XJuRskCVs7IQ7leGvVcnjXkpup+tbFdPzk+LOahBAeOv0/DBJpK+J9TD4i/uoe3f
9kHle7kGpbH1yt985xfrD5F9p3EYrVxWJHsJNf+8agaMdifq8REV5fWjlNIhlBz0
Vy66oNxyu1wapTiDLHqx2rC4NoKIrTyD07MXPY4FyzkUOxH50MMSVAbKld0i5KWJ
E2om6/3wKpj5YVZDzI+Pw164Hi6FEkb+6WL3HBATywx00HL0JPzNtl3H059bBue1
9vF1rVRAsLqEdjAEcw0PrD49OHgUIU2mLwqHR5ds/4xRjWGZD2dMUsYWseXezHdd
FwAm+mn3UvVUwGpM3Jk++s/HgTuOzNEh7Bnt/JmuToLgo//4Y6fybzEy4xJ4iGQn
0gYdCV9woVJYKSRFgdmHcpRb3s2v1k3t6kFej+MDDpxO3o11wCx2HZDiK/Vdpl8w
CCCkxj5yRHS5KG+E1Q87MIzBSnw0pkuqebXl/9aSS1k2Nifuyqibj5jIy9romcW2
f676eOQ9u3660zgei5O3FkmmZpSuLJEWFt/wgMLK9VB1VrjMTL80ozOcJrX1fsV6
RUywotUIxe/26HFtLPNMMQnGgCiULMRrruPU2DGlP9dQt8qFIEAJnyMWYNZFskfY
MJSQIkR1iIew6q0+jVqapsGv9UF9p7deGoaaDgjBAc0lQVRVQLJsOpRxcRetki9d
9sRPeM9nD2pD+kwVDRDD5EP8nQeilcRl9GuhuIObgoo7KZ26/4lxOycPGhEYt+JW
F5W9M9OxuehQhJcS6LVU7n7pm7lkYEhtbMpMayBzSig4ASdGMAQw7cXR3Vb520yb
prg/Bo60iSb7Cri7E6GXNypAMIwx9oOxKA7EqttlEusuZCcP2F1PxT5e7F00j3km
G90uUiK4IO+1St00gsBqj2MJ/SLoAZe+fKzZ6Mh+aaC2HRmaPZ7meAS6vuInWJP9
DUfo5ZDop9FWjLpKVnOcG7ePiO+gtFufLcYXNDrA33NnwBKGYrbRTSc4rJx8GBAp
Mnhp1Vl/d7arR41A9rLJJvk1cIlOt+IxMi2us/aaXLtA+oLBpZKGiBJnlzwDcQc5
G6CLR6EApG9C/fOTqabpEFGs4/ucXGyl6L9SCUcqSjGHl3E/Ri1adp1jCNvR28gC
8huN1Lo1YEX/H3ixkZ0d0r9goZ7yQnaYJZjYQ0hK61gj0gjbykvTPp2g+ShGsDh1
WwlsO57SY/PTwvs95OE6VQgWXVaA5Aqbht8fM6PR+8U5DEq7GZIqBozHiErodVTQ
3bLVrPMF5MK3wa2Z78HadMBFxDibFotAQ83diRa8JM0QEfgq51p3C6Z2q+XoH2Ix
FIMBNmpYJifDCF/0XgKAX8Ezc8HpEmdkmC0UTDqXbXA4Rx66omSSQsZ3cu+WNNnK
UlJRs7MOX/qPRHsatXPFMbGCtPlR9IiBCnqLsjqoS3qMTCPNLtlxpOJLCGZasITj
cjGSo4E+WlWlKbZ3C0gm+FGvPqeVbCXxGIFSobrA8U7RwC0SESBAQuCguwkbwhBN
t4V3Fw+byS+ER2M8MUQa/o6dq/lpxO9WGhhnykSFMFRiRAbHufO1DHm7LhPyc9X5
E4PrB7ONvjx08+IC55F+92jUDppIjKDI20AfvYiPMLbRjAdb1TZR0K45TwOTwmbK
9+N/SM/SJZlR7oHegllnV2Zgjqe/3Vflldjh42IVPkzUsujJR5XQsxQF73wzADrw
PAcPTBNpf+d//kW6quidDWun/CI1gabELEZVq4ahKmXXsb9c606CO9l9NlTYhEX7
LY5Q7heXwy1OKg61aXwxwAlK3gPy/BLkpjLlmg6tpjCCi3/DBC5b8QEutASzZp0V
i87VWq0U7UXFWV7HPjhajThG4WekgD+PFeps7RA/63TUhwjg2GuhvtmJ9/ce6P/r
etvZ3PVYbkeWUe9opRmHBiiZQJr8t8kbmLeZQUcCellErmfAsTthNNoVNdPCoG6v
xLUX6oqYnCciXjdX2SI66FaQr/9wPsPNvyQ4+huiT5FTohJqEeS4uMpzecAAbRxf
Eli7kDbUqdCWJTbC42bZF/J9zCYUFiF3B+i8Ml+fVAs3d2mCkvfFxTFvYuxbKRWB
AqVK6S7Fs+lyqdKUNuWDbyBbSVoo+eFhE0W3d7wi/N9IM52gjahPPccEJNBQJIgL
Mr0H14LYtNoxxatsB+7uj6AY/xGn5uz2CFzjLCTZv3TnmmgRQvNvq9t+ISnkNpyV
WuT9KjTYSiY96IfIQhhDaKcXDfr0NMayFUzcoHfGAWjI6TsstOxTsPMh1/FeyXy5
vjvd4ASuHA3W5asZFoBz1wYJCtiLdq93t1vExYjRMlx0LLchM0/Pa6me/vWaHeiG
6+N6YR3srL3/TYneTXG4udYuZX0FuEysubJ2b5oS0D0JNB33h01yc92rXm5GErzP
mBPmFy3tX5H5Cj8Q/RYBtjMa+T7s+Qwpte3gJupPhTbWI2SZDO1mGmIplL72WxkB
ztoTWhkWVuz8yyDi4O9mz5Y3MfKGEl558WhyYomzFazTZSboIJv3KBXAduNujC1A
uhboRM1248se/dEbSDroYvPTHPqrsqOacIcO3P8aF/RzrtmT2oFzmTgzxWIq/4K1
GmfGiGifKwvBbrEg+PUxVlEJt5FjF/ptu6Bx7calc2dG1ULY3R8fGxP7Qhg33/57
w4mR4xdh7/I5Qh0/4rlYPswItVkw5/QzS632djDriMmZt6WWHJ6Yofce/7dtt/Is
Hp3dwCTehV1er1eFh1pfnG3V+VJgDfNtCB/2ispzdy3AD5gpHZTVco2Z38pGGUL6
pisauxAhULl4gkFH9pLIGFURyoCCxUSyPk1IX21D46BzJM8WRaEfAgQNNvnOn93v
F4bCXNJt87dj83ZIz2Af2K0yrWRDA4n0qe20qXF8BtJQ+SxpvN97D5shfoGqw7x/
KUtwevzZoWWT4RpyVkvGdOtUEAl1rL/ZMcT8jEwwk3sTIJ3qi/LB5Qq5cfjDgxXd
thbz6h8QI5RCsFogZMwmoC3B7veHs4/9udsZDYuT8choKpRkVAe1kw0oPD05Chvz
tjQLMxL2Ca+4XV/DdcppLR99bJ7stLAJB+qtmggpbYZgQx58eLktZE39CoEW9aJi
juV9JrnS9vt4PcdphuUAwXZLFOjcbikKl3eHHppeioDbbIRfankhPJ540QpkSg1c
s5wriOFWH9dPtLqOzIc9GrjbRVXy87m/gtAQ5Wq6CyXBw8+cHIEJH8y+kdkTOwHQ
Cw+ya5osQX0bYHWp3FzNuCMw2GVwv1RbVEavWhR9dJKdaplwtV/SpxCKA7SRQ0Uj
SFW7RcsIICaTt61Hc4aZ3hxxWWn8UBH7QMAa+g5nLi0n18DLhMCee5L7LAVDDJ+U
o2/Ht+GQ58B1g6p1PlYNCfSrZbfU3CN2lebpy0k6lz3tBs71vaDRotXBhRShCd9j
KQ5xXmdduYN3qCPeRxk4YnOwJak4q5r5SpxMckjfwDuhhe0sp9R4uplhKQTwTlc1
r+5qoV33xmigR3tA1wGdtb+3Wz9E8SLZfD6Rhr7HZI9UegBxUwjwUTXKHiHoJAJu
rMVU3i8/Sfr5e+RWrMMlzGgkZyWHTiOuBZpxu7IR3cFe5CqY+D+zI5K0Kff7elhh
PHCio4nwrucIu3h/hlPfByt6MJSV0chwdZ1y2YeHwWGIj1tlEi9ykt4O/t8hyLAw
bjKkkINBtWEWnoB9nXIjyWAdulk31UpcYO8vpKh5ldzIrQclFvw7aDAs5KY3SL/f
98l0/acE+0SbcxOoQMM+wu0B5Y1iIkqH5SKHmClVH1yORcV1dpdYYpVzi1Ig9NG+
BPANWK0dOv4eylG9WL2iG+cgMZd5UYcv4JFst7OeyZaQMS4kDSipVBlo0zGrxDXN
gO6IY9S4AkPOcg5HNFva9mljPAKzLawI8GVWFCwhGzGTCtIEsPP/mCP3tIKOnljw
kBUXeaDzr6bEmoumPbphWbAnaHz9+2DffijfPaTYCsBOIy+zsw1I3e7C6Ev93RpC
BvNzjGEBoUJa4X3aIojc5afkGFPXzP+iCagBh+/QCFQS6IoXeGMOlKWKzifxIkHk
j4hC2o1MYIsaAygKXf73jfM5MmsTa7jMtQetYQ1PFyVAD6ULKkAOKcWr8P1GMyzb
LsqlrcnvP5+XixhdIBt9srGpuIlQu6R9BeFwODPFtYGd1CwqL9IvqcbLxdUo+1yV
2Jf0daNiP8lHMjZg2lC42SSWBGApzejvmAnzuCtsTd+IX6Nz8LlClFQR6zohSe+8
0QsoYaOsbgMvpbDorjucFBC3FGuwBMlaQTSp+l9zp2TAkytE3hMp3PklwVz4aSjn
iiiUm8PD72dAiC0hQQvFvWkm0QytLe+vqXYHMs7JN/ZLGx1o0DTGcJc7yYomytZg
zoXhIf7V9tguMtifZIjdjLKnomPe12hVa9jNCG6cJojKP7ck8f6H1/C1n5TzTKlJ
gs9jGHbRoGejFbUy0Hc5Dng90yLWHjXm4DN50LC1Vz7Q3dXDhNe/95+ifXzKx+kR
YTqXumpfXLsvII/2ts86lrf1PRgplzkPSiggUucgFfntR/y9/iaPFGYXmRCWh7DP
d4aD1ZoEceWe5Iad9hbCSAAJ8qU77hzEM8v6FfCTn301Rdfcm3sYKqIw/dnVoGMj
3ZfuQDFdHhbKPNiQqw7/gjz2SabmU/mKZURHF/7hzHsB2gooG9llU6uyv7N98c4e
L4oeOQYK9SVwc386DEQL28Ohm9B9Qc6JT7si/ecw0vN7h6RMjfug4go5LaqIPiE/
ieyybu/O1pmwpC/vjrTwkWC0deTuBqhd+NeiACh2ntJnaamob+pT/VaAjQ55CzKh
DX2oR/kauwb02IHg6OOn4ENqH1wAshFF89KUzvVwNxlMb5LZ6bvFjXFDyb4xS2s3
hxXp2mrfFrb12rhC+7T0S8pZCVoCQT1biEkPhUIjfMHo0mvcnyP+UXBPk07XHHdY
i/y86lvAhuY/7HaVGP6woHuIsQ51jN3FqrkYn8CttnsRCI0x4755qMxcnEcb+OWG
u7aJ3sZfXQKyafVev6BJ7FPHVuVmjLYMphM5QdJwrOkkwzR+KGErWFcvrZ32C81W
5pIGjHbHqWxEpxhEI4aVu4jebB8TOmSE68k+rB1zoHRXGAU3Nn7kHUVQlvBEGQmc
DdzYC9W/KDpyx8tTkzdXLSa8oUfO9DIRyWthwH26A0uo77wuKu8PCgvovu34jowJ
/JF7aUw5zf/kGWNVypLjBRGaAbs+VmjnjZENrp3/N1BlTy4ktcGd94DggPcbj8Nb
TdZYuuFUnGBXRipsVVcWDyA/PhoKGvkncAidPqi2JeGDSqzj95eRznp4dmFAK6QV
qEj3yrk6EjZeM50dTH7SBKyqY2Z7bd/Vmz8FvauXASi4oTaTPUQJgNMVvgv2ksn+
/e0W2xi5BLhb9bqzjh8z0+aAtunh9R2snJh6SyFvsaN+DFfJisGTKyhU6jPAomOX
3ygo+igQXkpOblhYM0Hh+44+48zvBRJzsLpWYtqr1a/d6Th48DafGLHZk25UZXGk
TCsl9LwtbyLmm/0wYmVOv+nEeow+X7RsmRNH3bFZ9M1cSls/Su+aqEe4S62uSQQY
1+kzbvWsfXWFBOTo1KCOwq5V6YbswvUG3toYABoB/fIGyZM/fPwuO25KNf5t3LrU
JtsQxRXnR0llUApaWkLs1wxJ+oXKCReTG0Ug2dzI83NrhGllrIdqALKHBaSidXbD
wW1MAS60tUa0DhOhnjC7QMmvgzsGp7bYC7a2C2oU1dvLwYL9GXm9jEHacl0F9E0k
fagxuIMBUyUhdx2VCrprxbYo0n2LD4+7G5eyCWpv2TEjgjLJu6DAzoM5Up1zml6i
fEg5uR7HlnOo/UAwNRYk0hllMznhYXLsfMEbpwyjpDHHeF/ATVz5SXwKrxBUnts8
TtGU3ymimLgJ7AmVTYte3BYvAKWsMKR+nXWqS/j0SPhl1VpxqinvkN2W7Jb2DjEg
CxdtHenF/K6nwsFFii/fs3YxQQuQ31jjQdpWVw2ZPzH4x+o6wNVnu7aDGMlhR+0U
+ajgbZubMDFhVyCNhwFjnDUnSjX/K0uLROrm4VqaYwjfHXMNRntfq9f83dOCeOgE
yj39ctrgp4AvHwDDxGZIpF03Fshb1JG273KWmBDOjRFEWZIeco84m6aTUqSB99ng
xOaPS/K21OkxFNtDlm5Q8gZjJjpa8dJVWNpHMrFOTIZepZBvxBdoompnlqJZEqzD
YPQeTNv69ltGccPcqMVaNHjhzukUJhk9Ti9/jWyiB09nfCvks2jJQSG/8iQjShV6
33BUbs0Iy7km4D+rZYX5vWfwSVdMwFk8Xad29NipRG63urWMtxHasy2T9AldbyVh
HBClHbHMAST6aeDqon8YF0roW0JpkZZl4hMlBCFzbjbjFs7y7cg74QdaPV1BGhk8
Etqmr8VADr/B1faWcKqMvvyyPVMSu0D1DHe7bpbS0oXK+DvUa8szgy+0r2AFKL0R
MyZvEF9n0i0tyZ5FbfUys/vYb4JATiz2mVrpk9fJU9xD/EMTOledXXEDIkW3BhGE
HajImxIYwQFOyPNp0isMlv1uVbeI8pn+RPthiPtCIepPH3KhJz96aXljDK5vW0q0
uqQkBxFqNPogeddoO/U0Vqd6+0tzgwjQJZrfgFeYL6V0Tugh02O2b9xeJNTB0oLY
t3GqP62IJqQfFPhW98vWa8AwyAbhbEQEjAnQkw0LTTFskYj0r9D0wFqZukzjw2RA
JMAUTye62IEXMGWSZDeogXd86t37IJo0k3z0XV66xNYrT+TiN00JDASmpYF/pW7f
hPc6UTcE1Dn/hEFmPk+5VRoJjm34RInjOGwumiZfvc3kNPFiDVTltmNS3bx2nvTs
/9Dj8ajquFWGVuWVCxIQP1oRkrAPrX8CD/pM7e+49GjAMXwz8O/0TWsykso02M5C
1/I8ikaSb6YChBgjqGdWq+hWsNQqVGX9+qcKP5XuEO6FmU6NMGTvNcaic5/vZC+u
Jry3uJbOzbOgbZ3iH4CGhDhHDG7IvWYwndaW5MiZ9suYNTeXkWHxWVi56seOOV0G
snZSqboO+6TUEe8tO87Ts4BOXSFAZ/qP5PhASfLWgrZxCjj9YqF/QduKmMWlm2Fj
IL1uxKdxCsQ4US5qOt5k61GRf8+hq24baz7sh6IYPXNu7USr7gW1T0s+gdhMjkQL
wbWLlEKQ1HHeALxWYjSTMthfUeA++QnJh7ibXB9payNzrkSlIWvb67u43gpi1B5q
un88WpubvJejlAYEO490QZU0JtpzuMZhu1BkOPEywmeGZj4CzCYadiumO5gf6Td3
g3Cl7B45N4tK3JqzILeT77PJ9o9n2vNQjnTPFnTErwG+lTUCHJjc40HvfSx0vn0Z
WDMLyiYRe00pga/ndoA3nk7OF8jfnLURkXEIKj0vrFjRGsFgpvqowMSwVR4bKTHg
ive49csJy9Ajq4vEbdvWTFSuvR3FJ8Wb6gcb/EaDwOPOZGWNwrrXd+gsZ64gVGUx
Gq+NVQ5pHUArV1axPN33oY5U28IHsWt/3vRD0Y4MaCDLV6GsPVhRKTFY9/+96ats
xYJxBbLf7pHgK/Lc/4Mz7Zs3cqopAV1MFUoFIMiLXngqTQEhc9zmgZe2GP/vANT3
Qq8rnzHnT6LnmnHgliIMk38aeNWhl/gxF7cZcI+Rvaug9z2cmnnDNXBW0GzjyJ78
6rGLUAd0Fa5YxYNbOIxW4PxXVmUfdRGkbsiCKy/1hHozaLRzta9Qgsmi+8usqu/K
eSD3WIp6OyCVll6dnQhTrXPZetHmxGgyb0/vUqq5sEv5rW6IHqYcIBvEqajoPtvH
MnuC9kmPUfl6dkwyGnEpr9ulmHSEJLp1OIDKBejhSo9hLwK3IMah2LEcoh++BM1r
rg7TMuQ3ZwhZrEHvM3Iu4qEsSSJkWlOG/BZ3x1KdmcJ4NgotFtf3zzbiOY0W3E1C
jKTC5I5uRgCPcx2BrtwV7jzI3btd2z1DGXh50kspaKOCOr1p2jP84rHCAlag2leJ
1VDgsUWayFE8ftKyoR80hZriizYYLC48Q2UMdGgzRtE0Spst9Oampt5FPL/C1d9M
+Y6WmnGGJVG+wsTGHvAHzhbW8IHBjF9FEBJAPwlVt4K2Trw4VxJt7lX42SvSRUHl
qDWruBhuIXNPreoIDGMETkHrqIN8P9yetRkEk5SwRwTy+q0aS9yo0hVEr5Sq4FXB
nWgE8CwKzhIOw4MVvY11TpfM9+48RKfxmxuhEx/NHJZywgryiwibIjdG409WGvN7
77zxdLs5+VHFIEskScmpdYktTpO+XdZ/qziMlaVwJW6AzJLX+nVYwS5qpi0t47ce
QxRbGqUx8BebpcMG3R8KkgdEVyMR/9yoitwhuAtjjNJ5/GJYUeVaYHqMfcBeTLtO
lERmuh712BBJNAi13114tD2CfZHPPT1TaooSYrKaXK9MDRBN8GiCAFUXNKA66eZA
ewrPXss6ws+e00AP98rKVt6+XzOqGOjgAnkM42YBtGrAFCFGw6kgNldtP7BJEv6y
sINH7+gZ2kfnsVVuh0QVlQwZNTy6D6H2XUlTsxo/cVzT3Dflco8DIJjov1UG0LGj
408ya7nSfD4y4Prq0AP52gPrdnXzlR989nOWBMrk7nXBwXCXFD/71D9vRiDIuGBj
qh5c+GpJMZs1Q/Du8P2k6Z8ZohU/9BC1jSh/bFdE/R/+6mcQ19NkZ2WFXmrDColl
UBZC3FuWU2Pteopl3FoBTn0NCYtdxy3ATc4klHbxw3oSBbpU8RBrRU364idTIAy4
CqI3Gn8RNX7jneB5B5+d7wkfC5UK2Go3OaPVOJHd+p3xfJQv1X2K8e0PQoffIxtV
lMWrSSFh3iYkwkT/JZGAfRQTrQi9XUkJwpE8khYt4BpXBo5FSbETVM95l+IqPCqY
ngZ2YZrofc5iCN+ayKiCsK/stutBNgQqUqlCBpbo83iWqzPwOwdYuR0aTc9HAt9K
hC3B6ok66fWN6eOPvQrMv3YYHr7oySa1k1mB+BCKC1bPsRi9wZzEVD3g4XSBEpuH
cDZBg3cJ58dEWqbuX1TXauYN0+eCVY+nvn1jg1LR7TRZzn9xfnSd3Pe3dMe9TiCw
T+UbWRYh5And4QS/owv7poI/C8GNFSXvp7eLNhFCaHYBWFuR2o9aLa8SEUF/qNct
V635oze11AeSZRq4i67Hieo/PXELmJBJQpozjc4bkAqPiQ6xL1/iwf+eR7OPc4X+
BXgmQHB5S7ZL1auSjIdHmyZIiP8hmr1qPG/nL9TE4oKas2mSeC3d+/HR13+8HYvO
nwNWdsDGv0uQbwmiKXMkTOKOcK4Q+FySuezLBkTk/FibVOsYZoef34NWTROU03Z7
q2fiRHHjue29BtBaDk+a5/Jnpr1O0mwahcBWJEh3tcFEYN2s3a7lotdfITBjt+OM
iU4fvOQiLIiOeidQywYxdfKDxqT1hv9LkHBxQL5rjRx8LBTG//vg3pIeACK8TSaZ
ekfyrjaUSfqz5Yo7wfVRqjn+xNLfk9JQwhPy4UEfbpvVUPo5oOiOBd8itVzFm/OB
4bU6YX0C2qb6WeqcN/OiTUGu7BM0GBBm5GXlT3F7EKhG+0EbT76hHBoZ8r3wAoWL
EWITTrIk4oS5Qad8BqkzOk4GH7U8kuBb+ezoaVJ/L1i2/rUgpOS5yi4ihVfiP6ob
TD6aGx1wDf4Qv58QCMsVYUOrBq9ES4WYtNYcsoUgvTIZo33nUy6WvmldB+aYkubz
IKcyavZjJh70feUDluz9h0bOIuaydTuLnEB23Yw0KdSG5+N8cm58rL8V7qeJOkRJ
93ELQtdkiFNfCBOXS2IBszcVeK0h897CqNp0Rs9MzkHfOfA0SfrG1af+quUwwbgz
zlWqwr0LXfdAWYKgVMh2eCDYkL+43Tb6/7/31YMP8kgGumrILIwur1uHoJNreUTp
rjOeotXH1Qg8PDP0nvoq2nkat/DHidCPUgK4sI5EIydv/8ESkZV1YsZja804hbp6
SolKBCzpS/Z8EAnImwlHS4ly4TdRbPqn9e0GUl56p00nfs0ko+gIah7grG2oh8+Y
hm4bMd23XBMjrxAghgm3Jdot9Y/vu2CKQliu6u7qWV53W43DuooVToDJS5FFhj6O
68aqTPkXi/GCdEGQ4FMXAMNHWr1tL7Ou6Re4FjWz7ZnELa/RUhpeMjXdrTzZ/WpI
aX73n9sQGnMqQV+5srf8d9nzYByUzsK8zItO6DHm13PwesmcdRmBLb3pGcmpC9Ib
lwYNoRaz1qtxgfw4cuGnoNzDdRes7q4EIY66AOhj8TNjzcTQBKh4DXQw/n8qatpL
/YGRbK8P4TrM1bGe/3YuOdkO3yRrJW0atMusqR0LmPplQeeHfgusibH17bXK9ZXa
gdBtNSeVzUDFK8M9IF+G4BhVRXtLXoNuY5FCDbhXi/U/ewwIsthB8qyp44kNX69W
7/0+89S7G7Y/kZ6BXake5xLiSGlUTdkVC1gNFvuc6AJw1/PWVf44EzI7LTUwlXY2
/6pPxaGRftmxnppcuOtqC/zDA80Zku91MAH4RJj+SKJSFRKddlFhZS+OJ1odC1yK
rGLROlkk6awpt0F+4RtV9PlaPLIU+hNGpbaq01D7bCp+izOyh6kBJrWpJLtVE2+d
xchmf28//pAypaY+WaKk/kJFFBy92IxEZ3Ju/azAE8DIWr59EH/Fs6ZblgFGS6iB
L3og9XsN/5hUOVsziz7hysaURT2PE2Rf8pRrBLFKHcre6oaSEsa3E66WY+8KrEhJ
O7dH/5tNn44QqBp/YXcG9MDZ8MIOeZTQsWllabNK3ND0U1al8JvAaKCUAzUvj2sf
oX46PGNRBIxz87goOIPnEWaHI4u0KjI346dUMBH1QFWhQSLcu+rlGufcHnQp9Lx3
5VrFogl3brOUv+4JhnLl5M/EkUhVX4jH+GCi7fBxT/x8q9zNDJ0X75yIt9pIe791
9fRN/kNo6+oE8Xh4jwQhNIMZZQqRB6L4DzC6btQNgVUGZzYNAghmCjaDUVwZsmvW
Qt6cXv/1z9Q3lkiQTG939doYNo1DU7Evv3SzORB5cfG7IS111Tv+kDdM6XmDv0sz
hpIfeP3hxvb693LoIW0Y8KNZtcW9KPVzT7QUf/t3aEKBqsSQaZZFvUDmNqEVibZ8
Bm/kHJmFGSzDh4yhMmno3C1YEgPMlOiM0S7J0dawM2omXEu0AdlBZfBT518fY987
r8+ha89kEdOcg0nN5e1BqfRb3cNw6UN19o1Z+COrFVBKpiOCU0SuybmCk2OM4vNY
R/xNqcm0u/gOP8+sHeyPPAsiI5npVLLGEGQV6niw4JBu60WWtO6FH7btPL2ongNX
r7mp6E85voJBmWSqcZQcVKy6sQ99wOS2rBHCq45kPs6pqvq1UGTkROAJSDdQTwac
nWAZmKXNUHpAXpXcikktyJ/c/sX156HOEAc6Pxd42twZfKF3X6qpeUdAcw8TzJxN
4lPjP7DHY1cHJnqDgHJn5Li74MbkGxq1xzb9eS40AdBhqEv8jKFdHOE2tOR1c56u
sh4VjTUI74c0RM8YptI9kUVkroRL/gIdTtEIZgQiTAcqy1NjIua8TlJlgRtcH6Lb
OY4Cm7fEsbmxmNU9DBfcQj1coMptc9z+vfjMnuQXexOo4sMcoFxUNvGmt/pI21ko
DdPsLQOxihlcCM3epCefaCaiM7TgbibKJbpbLiGbXXeezu6LJK4w5UXbLKrto1cw
L6SMWoxedabaz+n7+JnHq0jqooQTpZ0eg4IxqgT30/KrZnoeIxRUI8P3pUAhVhZL
i+gTUj18nZ7jCmp24Xge/pMJ7XExMHRKGdZur6d9DJD9MQ5jRipN7dt8XlwFuziT
F9c8SQnNkMUbKapZqq83O7FmrrM3Min7PzInd3Kkr1rZtOnuNbhPPLzNN+VNRGTj
fOGaF40rBLMfMCUY//mMjoaj98+zoIEK+uEMrWBok1AeyyN1V8wiD6N7dlC1yWRe
LKDT8tFTWXpMrIsk7xGe9owqBm6HJK0VtHEkTcD/clDB/E1aPIUriaxjMlEXAu0B
sZHs4+KguxC1El9dgJP4xI3XjsWOugfJ5PQXgh9KJI+63HFRS6FdDMnwMTlGj0bH
klZa95CZ92hp/1/LyL/rsdqE89aSwmuAKS26haSG7nCL3yl+iPQ66NfR/tMCHYMd
dDIW7i3A0xYV/6+8vW28lRlfFB81UxHgq33qcIwVGYSQKj3jSZTnnZtCkE8XWO8z
i+xgiLZVTwW26QC/UfcaDVWqiKE8ycRBozhQINOWaVCUOi0OsDjm8/b4cdBN6TPz
Hs8WXjo9NnphROmft91ogEyPfxMl0XFEGxxUC3pjvRPRIHM/51uFyykeXVogSwDe
RiLQC1RL7x5tDCwxFAmNxkFea+5CqZBSv3ooRWf0kLM67kvuLV53y+rogzmHUAxX
2MaLiBimbuSEBZVC4f8aq8f5eJlvoCzzksQ6mLwJORRAIQthXK4sd3CYAyNCejAg
cgqlsv+NV3bJubfRMlaIvUBNUDiVrrcYb56myjSgCI+UQY7a3/2gt466MxBZCEn+
JvoPfbAYC+/OlvPYiAfqPlhcLnge71xAjro7ng9rjSrSAGKgNxMnYKmlVZ1kN50M
hP3arMWxYgUEmftRIutxyPUmooSjpqB7kXrjQGJmMMVNuj5nx6TSWqS5JitHziA2
WCGfZFU+ZWRIBgmi3u8aZEY+5gpKO7fh1j1sfQQzJMiDkJSzzr0ALDoV7k5re9Jr
V14b7svhmQTgkBZnZraUT6c1HAyNbtsW/Tai6xtBU9zPOwdRWqAVMRw9kE2r4ZY2
xU54kwidnqe4Eapr20MvnPnkvE7Hdceb5QCFO51CuvQ06FzwhJvmvaSbfcsoFcFb
Tp2D0IVIoJW5Rsfgp0YsgkmDoDnon4vmq4ZpsLSFIxxOF557SpaguGhXyadRedX0
+quFk7MGZg8U5/mUrIi9rWTbUbS6k2G9nPT74SwvRj/cHihJjej/gFRbj16YhcUG
/7fDoNEXyMIJ2KUTR4ePgLlJkmK2Y9ixFVVF6nl9b5bdZjFWsCQjkXwjTQSxR9EU
dyNsZNfKGEXTYt3UYNpBu3IUFCLaDBCzEEOiOS24xr4bEuWybmv/tf3an9nARp51
WIX5b/JuiOUSDprBiZE0d0gJdZnlKza+KR3W3mM7QWSaH9wQbPLQYMZ4O1SqUKG7
SuCMRi8Ug3lXj+MAC6PYBLhcrJzqodTa7Py5BstZrZ/f7MsK9SaBT9t9Rv91cEe/
FKLVVT21RyJJX4AaJEWqtf/9ianhFR1KT3e/ITXArKrctbCFv86z3ZfUlrDPQv3x
2XfSMq8K2A8FiZv2vWv8mvBPpy9nl1bkrUzBTgsCo9sO+LmFaXht2nJt2Qrh9MF4
AmqWD1ohyoStu7Jvr5EFbQ1xPiKcF67vzLJ380dzHhNctZG6N1JKv8CEYLD/NtGP
QvrB49NnzRWlWdFEa7nXhlTDsXiqXMU487wWuk0ccnosZvy3kDzHTcG4vO2olicD
Of/9eTXXcG+rIL8LVO+MW0U1haFQyLqnfnM/jo9uG+BFpgUE+CK4kMxZGf4txYCa
6ONq+wEfyMsnVBBCu6AnY4dnxrpi9UXp2xwVECrhGNRmlbKRbIXCdB+wH/ZWNsYi
qAnp5jTGcU++lor0wlZhoghTiAQUdMzEHWFMCDuv9vhYTrAbiJ3ZFvPyTp2yV3qS
7cdgNu6SMQf7BrqX/73NsIqoaPXXwJaZZnRRt2C9UT+TRaUfUau5pYgDN/2ct7BX
2zDfhDOOD+bKgUJqTGfIs9uyJkBPG75m7+h9JLNLi82XmA43f/lrg8qhg7VOTPbT
TqAHPJQTxcQEBGBG8madVRDdd9J5CEpwES1Gt+CfDmVyi0jERZOFASaGSMArGmlT
NZLUqglTrkCDei4Re5PtsVx+zoefwtea+JcTScQkmvA2pBm1t/efONO56P3U9Wv8
Cwygbl2vFuTiDdsurnEUVF3+Av2b8Bfw3XdG53soOArKMdM5mbYVcOIV0kbFG8/N
OWYj7qQjJkruIquekbHDvEUDaTblfmf6Nkd+Lqzn1o3r1SksxKyqPlTiuJb1gE7K
6vLvVxJEjyCZyHFzsSax9FvxORUx4GHtI6ody3dEgNZM2ajWxB1h3r9A98qxVp4A
McNXk2RAvbMOyjwTriBRE7dtrlb7uuF/x5a2PV4yB6/d9cpfcjkzA0cQIWTccjCC
pk75xMQK1pf3/azE1r0IjDkWpSmNxbwIi4mDzAEKp0zsZ7nNbzI6NmG3z+6gaKGu
xROhxI9LKEb4YbfJt+XsGV2WpACnqUr2RqwcN0D1CCCT+f7yxPlqQRlzuGar711M
k5afZ6RfA2BE9C8+6RNtRViwnx1kjTJ3A8EuW0Rc0ASZOPcyeAGu9ZmR15jr0EWB
emx57kBanvna0EoVHyDZ9hqLhHFNNEui+IeCLtQh76o7zACCJLlPuNSeXvVN0JuI
2yAKDNWCt6bcTk4wMWJwgciPD20v43joyV6t6gW05o6zL9PVv00lSWowz0InwXy1
MQJAaVgG+CpktbX/RY2AdsJ0q4CPfF4zsX9YYjnQkJeWuT6Sl5h9KZuoYEK2rRnT
ncUotLbXrvUCTSl9/qaWqT61k42Bu440g2VnUDkvd+nIpkQtNzeme95HAjzt4cpf
dMz85aarXYUzfI4CATJqixUT9xg2LS3BfhpJsd0RqgUezRP/W3ajczch2NcRphBL
8fN72/2oPzxc/Cu835l8rYpRhDZ7sjlBKqNVwjjDlt5K0Y8RioJRyxoPmmMOoK8Q
8czEpFgBi2Q/4dVz9MbhgqWhfymvRi2REqVdLktWidDHit/8deOZrBrfOh4BfJ/Y
oZoJnZUk0UVRkbEyw8sCH0ZbI3VBNFemcj/aq0pgfegt8Z3oqQGPDJ4qda83MPMO
K19yMGXCD7isd3KL8wSeOBvDm7geMJC7BvJrDJvgaODzF6YkZaOHOz9d2zgc+N3U
rzTPbWIkjbL/ep29N9/4MeizaMeLMbcGzGCSnBF11XZJlwKexHnLckmVpzI2TRqN
zQB9A2Av5IB7hPx9Rr8YjqL9MSGTD9OFug50CUpzghcEabsmHAJvCkrPanKlR5FK
Vi2+kP2lGW02a0+agg7GMzmm9mFBzEEiCMgutM47znJAA+MKoe8jADyp4T/nRQ3o
X8dBmVCiam9pl3kdhh4Igj2joWKbb04SCbCvWjdQdAJwdeF6lD5M1/akio/YplgN
8t/mG1612ALzXypbDjMATElfc756b2rYxmPVhECpjbz9Qxdez0HHTdCp/KwN4AlY
l9FtohaVWhNM40bNV6252MRITUNCfQ91EV6eQ/QaOOjxb+qQpkGmLH2RW3rpGadP
GhrBhvweGnJN8lA+x5DmlRf6xQdC58pvDmLKwi90jAvOyqHpD6v+lgtaqZ/aBCas
wstDgKO7X97tycwNss+Ap4g2tWXwj/rwkS2QLoBvKDUk882p/gbs67JJxfmUxVVe
fE/1F6uqj+DfYX4bNSb6uw8ALs7zpt/i0xRcnCNWGDW9Zn9nnfm79+K6aHyCDAg1
4EXyUVnRxCbphUzmB0jMPnZa4qdUiRZR68Z07BDFm6rhOs9Xo8qMjld17l2IWR6l
ASHs0Od+q/8V+r1jOYErS6WUE+wV6RrxOPhM9ongLKrN/Ms8ftbLXu5S+sXCeRFC
VezCrfrAM4Lwv8AL+eFQE/4iPCU0WBZ4admNuHdUCdZMEglDRmunR4sqCHqQkV8T
JpN2VZKHtI8oWpTSdEcTvBvZHlsctuIjyrwPbweyNkctNzbKpOf4RYIzNrJ88uyV
zkZ9502E4J8sGNacj1N/PPouSGiHBP/EX+qN6S9yn12RENFBGsTi/LsY3O+7Khgx
ChcpfrCrfIFxvbP9SmVkSOy4bKSr3Y2N+YFlH2+0d7K0iayD+HzQKr8GAAnT6nfb
W0oxqTB5wl0xrtY05z/ZmR819JoBVBatB7JT0uuZTj3GX9DbQwUXkc1NIchoM0xZ
Vn7EUad876uGE/Hu/hRmTHYdTrrH7UBpGtejZVH4xkZmoMwlbdmhO/Jz7RLJNrNC
Lk6Ka39ZsvZsRLF43l6OUQLeddh4W5R7kLkq56h8K3EoXwivmUmRtlgXTDvcATjw
+AiAeypoztZFC0QeS4qZ3EPAJubh2XqtucJG/N0oOanUUhywCUj77YluqGR6ILEo
yx8aqmGy+C2zH3zb6rt+vXUQEWgm2mxF96XX5SHm3W183VoP+/UWIr3qXRwpXvZ9
gjJrp5TdafT38NtOoY4nJYyR2xFJZyrLbAhff2EnePobAMEBcD/tlcv5KHRYHidJ
7XHQTHc6r5LET1knjgj7rHm1Pxp0++f+OtYOpiwAbKan6ZdeMmAJgYXTBeLdAkdY
I3n8n8x99G8j5pNAS3OQ321xoDU8YjihsnVjgyE6fnSy0By0/nLEgSaTpgWg0kGB
ZsAQwDtHK6Y6jijFgZSFnN5dq/iDdh22Frgql71pYNA62uXoetcyWji/zlcrpljc
jflMaJtDtwZKibscl5e5jxAh+25sZcfY8xS/QXNXiNcBt7uUreMRGjZqNbxC+NQM
I8BAIyWIuQy1ps9noz2IPjghs742dYl3uzU93ZnloSGhBfmHwsRmwq5xGczLdALc
FV2J1vnDG/MOL6hXVgN8GFI/B4bDBj116OFdGxLla1RTkQhJcoy+uWNLt5YOVmE8
7PxYIa7qyPoWAqb5sha1sfiawINuzT/TR01znfoSJjzDztekp+pcO63Kod7YNeIq
VNbW8aerQR2zZwFrpKB6US8KElBYWX3z4frsUgjQ7Tek9B2sbbXeoYmGRPDW/+0e
hTL2sW2CoX3KRMRXb805vROqNTXd3XB1uDpccfQ9N/bIU49Z929ap11RkxSL8qWp
OUU9ArWB1Dx2HnzigEcIkXm6auKl+zXNS3YdaOBbyDXkOTQhmZMNi3uOYVsUt3Ql
aPu80t/b7pP3MSWqcq7oG2/58TOu883PTixTYPcNfPl8Y1jh5Q8nnX6obrwZxZet
63xZXLprgPx/P1kpL+uYJtP3ILlxbil0bwSPPzvXTnmi+Pbb95OkX8JkHCG4PfIZ
0bJuf4cjgsomZkc06b1i8tslb+KtekD1ErFh5YBRKdiEBum3ARpKVBDMURGto6RU
F8I2ln95EMUzFx9L2PShX/Kcc7DWH1yxr2Wk7Cdiw4Y1jqNdqso8wo6BVtmyUZya
eHV5FPbu43ezVjWYKveuyMbMYovWGCwnTSXn2QCy2G47hKaEOgL1JxkqlittR49a
BTLaIVZzgVKoDgwaonu6L4ZDXoysNR4xCqBQS+57W9WSnQz6IOZ4g1K6JSLX2TZW
asTuWERCIMfozhWOzv4f0xwLmWUWHxl3rP42vJ69H0xc2SfzQ2m9QZpNpATD5srD
u+RIEG9E9gaxlkmcyBBS0eT63dLLAZg2I/XPAopCiXAbqxE30CSlF+woyAVYuVWo
EGw+4aWB5ouFHHxpJIxjsxQCcYYw5uhq1AHuh1N/vN440RMHZ4e3boO1V6yG5NWE
KxXfTzgIqVmjCF8YehM5R0ebcdVGhPcywCyBX6fU1XS1vq9zmbih9/eE7WMHyyt+
YKl7vxUMesj52q1zVvxZP2zWuey1uvFAN0kWBgPMGOVa3uKEEpISFMA7lWabLG5S
ury2bSfAvbmVScuSyWI5nSd7KVNyCwvgTK89YFYRKouNgYDkgx4w+1MTglPp44/l
DuMX5PK4PTWsORRzmDpXWvOHHWyvxMXUq6gYw1ZHxsft3otamyurv4stijehWMcM
wUpfaTY/Wb+lKy2N+8nXAlL1X+WjbS5F1McR9y/sI1YuN4q25AtFdaOhKjHoeis/
Cl/jKkNXsw4tav1LRwp4XIirpFiFdFVwMpFt0GTC+Un8t1elnZ5IjLuyhSS9SG06
LKykjWAQW7P3tXid7l8MtPPFlqKgVwL2ZsN8wEDYKiVXX+jI2ysrU8MIbJ3f6LxE
UNN59FhHHc+2qMe5gc033O/jQ+RK6iOQKBzKFCQEc5yD3RoQw2L4DJnZfWq8lLIb
bX9wlrygUR5EjevB6psnyCkcjQzXOTYkkc3Ir/3h7DTOdCLvtcDrCBLFXrHXMj0L
J0oY2ENb2nQ18zWxsf2pbalYxGN3ZLgAKNP8ZNt3MiXAaqHao8UlSMJDtw/40WsF
+0lPhSxqvIW8yk6Zb2axBlEn/fT4wOvpZeTvQNLDymksCcYGgPH48qMipo2YmuaW
YhGYIRPIXzo2nShKa/R5F8hjM0VNBYaE0aSTftRiaRABmwgOLX6NNCf+uFIIxxwK
iLoLZJGi0voZlnsxVLhsWSzCSaa0kcyV30XODHDdzdKcCHtLGb0Hdgaz4zCq6aZm
FpsyBpKWKLOhTZFlSWtpZS3hq8FIjcyDfpjblcS6dKgJj5Br+Qty5B0e8FpumL2K
MronXVhbTEfA46tiLE0IrD5rNzE3D9c+W1s+DBl77GmWnca4KJkndBGRO45LZdw9
Om1FW67O6HS6yd7Fnrz75jkWULMWjCeI4fbt2YqeHU/H38Q71M4qehpWvgqRg4Si
t6mCKSNemb7q+XXA+o38CixW/zSZf/E3BBWAw2dsxtgSeeZJUdjt0P+NZvQOppI5
x1nqUIsUmlXiuNhkh7vhpIaDfCZj/B77X3vJCSPzQXcQHj8JNY2Wn/d9krsR7hUp
6/nG9oCJDdIhFuRw/5yhw3Ao+mTI9qrZg4kMGAKJvTQMZVu3ZAh0nKGKknfgiw+B
hE5GrjAClZNaZx/jSFmK3GQv7oHnZ4Kb1DhtQtkLYRWv7vrllq9ZBdbBTwa6/MUY
71RzYlcu6M9tIT8/or/PoX11GPhdkb7RrGobcvvjXzqBMpABkB2NkXVuqNfLz6Yc
laT6UACGvMlKLj/HZqb2EExdnb8GEBFZvs8cYAf+OFVMv4flubzvItalRelcMVKU
PBdHF4PnohIN8ZVcCxJp8t8RFMWHZbNo+k9CoKYLYDXKh3Yc90DEbfFTl7AwBQ2p
Mu+4Y+4hhTQJI50JuDfA/L2wQT1enOrlufSpqrjg6NzqZg1mqjCJ5CBAS6Ah+PHg
sAQgPGP5Yzd9/rMJ/QUlc+7xfx7bdGDdz/OhVGbplqabxIL+ns9g5uwOzJgrHpzj
XIGkCBwyNZzzr2/r3hHSA48sMh48G15FfAyiGAIN7TPwY1pQtSRJ8z5Y/n+rI11r
NTLH/zwCJTLQmtn7IjdOroy67Q5M5sljE45vjwHo2O7D21x+vzeqmFpYS0Uej0Nk
2hex0p0igTX22JoRXlr1FcmxPDei619+AneqSNxH6JGpjhb7jG6qbN0DJXq/jHGV
y2aVbq1NkbslU/6BXjchYz9NVm26vsYKD9bTIh3L2JagDlgwA5i+wsI0aP0cJR8/
v7hOLwM2k0wosJZV7ejEapjHd3Hj5S5ddhNPPq8rfOFvfQs5WVG6m2sRpM71QGgg
mFUqenabVRZSjW3CSuLNFLQz5Dxl/ojI51i8n46gC1WTX7wpe63o2mT74kHowbLq
vLtduRLlJYxKvGAIlKu7feb+eOQTe1F1KcQAmCsVpu0gV9xaaGS+jNL8gLOq3UwL
oacD8Gs4ufjxyM5i4h6F/GLVQh7pmipvu/mFN79HJ7C9S3tacxCDpZjDON4bXLTH
TZlpzdOfX9nCRJj/RMnNyM5PhNJ6mlY2G90VEwCbxJEyGLrSn3RHilXQ/rNXV8/F
c0mNv8bEmkLPrUl7vsiTaw4hICAjhdVh1dPXRNgOxF3dUDZ4qAhAvqzzN6EYoyc3
ri6AFwyj3JHsl/WVGZxSU9eTHIqfU3A+GbDRTYw0czlxG8m6QaAITkduuXQFLR9i
yg5C75lar6eIM/urave7wemL/VqUEcLpc3Pqo3WAh05nMU58mPDfHIm55LdFMm3B
xZdRPzJllsjLV95lZN4oLbDYD8uVXE4cmzkoyfi6s15wK4p/rXsULkt5ZcXr/YtU
golBk9LvstgIjpoJKFSGQUCyVBCMaJo/iD0xhnSSTDpu5SoHbEL6DIDyWeBP4Xs+
JtzaJaIYuvQo4mTwbrlXabFB/5xbuksHNu8D58+cAFIPrntu7a/tu00lqkKc4vm4
/C4UsHyWwmOB5deJJjubRKMoSzfYsUmxw2FSPa9muCNNJ6Yd6i2jwTze5lhWRhBG
Yh1el09swnj2qmtkcT3hjvMBRxICXQ3YYCFO+D2EAkhWvKeu/sDq3bmSR+6LG4vX
1chYNhnwQrxhPxmt55SmLfl0QuFC5b6T84htbQTr32xa6bo5LyS8FpAjldajpCfW
nNnOrnEEXLNmJECEeRDmf8hQFtpkttnBdhgB3xwpQNb2MZHByhbf36QD6YZM36S8
EGK1rl33t3J4+0zr+EZY8omwT23xgiG/MdONdR4cH5kVfZ6+SJrwgL4ERZQn2Enk
2hBVu2PRNyh1SOc+sQypfLFMpk2DR/nya38v3R83fc3d0Vm61dGBhJkNZvNMG6OB
xk9ZL1Up333Z1dPizx3Tg4lD48ao+TKq2X7oknaayVtAgfKHJOphvss1pej3C+rG
CQoxruEBV5xqbq0y3JOlYK4PEe7KnSVbzBvA5x7Ujj8/YXB2pVhNDrAN/FFHUjbz
QhzP38LdCqiMPWaSlEtEccxiv1JkPBBj/k9pTBrDKzkV7mH6QLxDlpNYTS/jRyyH
g+Y4VSlYyUWM0HSk/ZB7wiMWAC1rEBwgxbgwv8HYlQbr2H+DHt6emXux9vhdUJIE
3ryliLS+tGGE+DwyjJeoCRbUSR9pjXGsi1G5la1lYbmbQBKOENuVHY5eC8b4mk01
Y1nEjsT00FG27gkMwohIgNy2kFWemkMSfp7vlIo63PTitghV6jkkaohv7WDnsG8j
hnZuBZ1IgmOdTpdoOJtfshnOn+log/AdMftyXU6evRZiE4aeDTWDnRFiE2hMrNfg
k5kSOlFkgdx3BRs63Zvrdkm1tdOiJylzrxIdPJ4Qnu/ih5v+HqdJv/VCnCEGOVOo
Wm2DqYDXe9geanlcYHYxeSAwurV6+/8KioJZncYihTTPkbYfFF8JbYQ93Cars1VD
MuQk1GAxWtuEHueH/1C8y6cl20maPv51DN/yuOy134X2NEGPt/h43H/7GXAlg2h7
8rnkEbyERChqBFnPjxhxvIlRm7/+Yo+tuoEZUH68p/VbNio1emWe/HlRCnxWDKuP
fk3Ex4vGztL1eH7Z5sOGiPkEHJaH5AjBMyoZjLKqkUUwwtI7w9dhd3rb8rSAk4tu
7LxxFSqBHBpM8pg8obea9qiH2L3didzoBREIIeGxj/Cs5RfANo0r8+J7ANNkxHlh
2FxGYXrunhZz3vzZEwaDcQaUEkC+MqcLF8Ya2kXBXbm5fi07XcTpfyUNgs1u7GMF
dRvZtmDWUIIQQi2vDSKBKSTJZ7gsAh2De7VJZV3XH2MGO4H7UwPe9zox5owYI+8W
GoNabs7Zau2UD/OsRCSDxShQoKy4YdaqO7p4NXlk8DJahkcxdlm1jIYl3EuqJiHv
9CPF5oz0CR6xfsLC2jAfjlkYbSyn/He08AywLNh9Gu1e/b/bD/Zme53ji0xmfS/p
xdbgOP1B5PeKV0rOT0x1GRymNnlODF4scvcoqs1aj/VxGHYLC8VQleeXoUMbsxKq
C6wFcMT7rcpPs3vKFiyKhISvFY9xocHvwF2Id1hHmI1twrhRr2xKkiIKbMM42Zwb
nBC/HCCwYd7Dm5i/S0X5j6y9hc3KaWFZiNJ7naKBnXx5Kr/q4klVWmhDZI8NOhr3
4mzxbG8E/w+iIXz8YBSsvoqbIsR/70wVR2HwAPQtmFbXBDL8O7Ghz7K0LGrQAo0h
wmp6nrmFPSnojR6YeLZnCivVLQ0q3Euv80Er+VV/70WOIVWo601lvurwSKUDkEqT
RSgK8YJoe08To39R3i8Ok6LCcSoHyvtgYRL2CzWXTVeJspLZoUwMsO38Er9lkM89
8QKZYmPZPuI6eWjtnXOcGvDoM1bHrWaNuIAaq8+7EIUAAlaoyRtKKlwmgZDAs7Wk
bcf6p+J3t2ChiHHMOzI7/6pjyQ9WYOkxJTsIT/66ZH+hB0UBwJrdleA8BQF62ygb
aqXZAsISdTxJ80+ykALA4zCb3JiVk4VTt7PMLrD4IRfPZpKXObhY1eYZOgCPCnS8
N1o7FG1Hd47n+IntcuUsfAleYeF8rh9o8Qr+1WVoeZOkk1YbZmhtClIcLyhZk3C1
Z2IylK11nCFhBBvMi36Tg9cuU5mnmSIobFgMsW+J0nCt1PaoYUC8dBOm7ONHYJyx
uzOT4VBEZcykov6OYrz5tTMedQAJsdLa6jGOpaTAZsebHdJPcGoTLJPNROis3QZj
df7lhdgBYO+ncqzU63cG493FC7eHo82mTpCg/dSLgAu5SS/LjMJaZw21lXNRPxyY
nCPeaKZh0QXm2/gHJL6to2Y32WUShleF5HZqecGO3emikOwur+te8wVOvL6LELeU
YZKeo0JZltNVbgoGV1z9MsgZfBegXQDbw/rlAOS6H0tFvbZrrG8T/zJkwU2FANOt
sSJYE1F9Rx8mkCHnCJbQEEQhJuL5Y/CZ46Y6OOBzvV6xn+soDaaySS7P2yhXxrtn
1+H4IwdYm2i4zbCMNNRZjWfQzRGemZ2S2Qp4QWUA8y+ygwy552ltSUy/jNfHGrGi
n3KWwq3POiNwmaRcB/LaDqed/2w/u1FZrSZK1qLLovJiH2rmzP86PLzADMO5yNwk
mBSgr9E8Jn3EJmRbJOxrIfhJ5/YmdCIqwLCcbXDSyqw60/yDcBvgeoqe7ILOkNEK
2Qyr2CR4QIUYW935oC/+Q2gwyvQQZ4R1yctTGs2qonI4QYC1GczkK4ZZKjsfFalj
crADGtHRRnhPtsiaqvAnr9d2ICXIRsfqTpkUDdurEeu9RhiU2tsJUJ+86QZiiKie
tvcWaOte1frgOl3Jd5bBx5XVRTEJ3uXxj3nIeAHruhs6Odl3LeWCbx161CieS8nZ
0JEzYoLTwebUWTWWvRBo+nUqHdYbrFLD1Xmsaon/FuZXPCX4vmtdzRV3OfR2Cu7q
Gj8hCmPojTDkuPitq83QLFM/oPJAyyN+hzGRBZRBCYGkpsqYJAYyzVHvKHt+CWDw
s4g5J3v57UU6LbBSQXVflrTod6IxKAZcNbJbSC88TANeRZVIKf1W4st5SwUXhHwQ
95eHP45uALlcmwVMMyo5DOmjLnwVJfZfeGWYHnGeEAEnsCCi1IkxIunV+vuZSyWO
N+PUGgDyK/lauF/dA7NvQ/C3NhZt95rAViFeYV5/FItQgfnH6Xbwvjtl1cjzPrJi
pU/GfQ8JAhtnQKls7qZP5AINFgD04OXyKw/mTmoBWW2SaPEtGGuNGH8Y0BL8zaEC
XUSKhr5sGYcu86Jt45V2+9oAMOLIOMkn+F4s8w3LeSn72CwhfQ4hXmw/Dx0mQjhC
L3jawASBaXmz0Bba2CorxWdFAe51jGFtUJul+6noiYBA3fXvRZR5ml/SbDHH2mEC
d81okjAk/nQ1xpvTKZUBT5s5ux+2gllhcSIrYLMv+j0DCp8LphEKGp4xSxhS9j7n
pKr/Hg8LBCrQWM8e6fnNC9+3StmV8NLiJBKeAS6+vZhJwI/8G9mxpSutIVxXVjZS
982ydvvBNsdLSMRYDJeoA4X188FC9W8Fa0HSC5fUW/XKP2JF6t/L/Jxgjj+PiPvF
oRFg97ou/r565R1k4DQVuNlMBSdnEZdMx8IUKXQep8emwOeWFEbFopbc89vqH+++
Wxcmi8WGcBhCqWhGkXf4ocWjCXGfcCexxbDumNEDinGIRiOTR9s1darooAPF74Qf
ER2E3S5b5bxpJYqtEgl0I3SWs+StVZ2zb42MGDjm7kRJwvAyhfJtLD2hpqDS5eXA
xXaxZp7+i7PJQCOu28cOX+EAzVoFz6OqZR/5DwHfFNTS/q9T4OUG77/rdmYPMsZU
XC55D5CViB2HseRTn647ZkQW6cF62pEolGhDVI9QI80QE05igB6HjAppVVELpv5u
+2OUnDFyXe5xWL87meln7QT3d9V79jG/4FUCfmFMCW3vHzslpr9xYyJJGYWcvCys
raeWwyVPjjV6L9a8m4amYMqzn0pkFpMhH8BddZrvf1fG3q3d1ADJBHD79h/8rHYg
qjUq/ysYvsvjh4od28Gim83eCNhnI7PsS/S1K1r0VeMFIrc9LLMmtAXTpo0CbRCn
nmSwUSnoum3rYjlOrhzk/kFBnmakUJazMUFCrxTqv+vuAJ/3QiWpHwp0QBg1YaGZ
6l58AmDtrhYHUXtoQLcP2Sxsi3zRTITWBOy4gHjdDShJo4EHHwIninc9a3b5JW63
lBZAtDVdk4dZ1pM2xWHTHbiRhF2O/5s/8CpZmx8BzOh988ummwI+Li8WYd/0gvvU
w6gxErFqvHmZM9eIByfJkZS6BBP9hL3n3LrbfGmvrrYFYLAGv0f5YIq2CJV3naaE
vEV3L8gFc7zfGPr8c6okN60zN0h1JVka+jwpLBqu/A+vE6C2CvTBj8lqZ2V6l+t5
skeszqro+ukELtsp44ri529T8x7sPEd1ptmlcE/0HMt8558+DlJpkz+LNZzBOH40
YyabLt6NSPEKKcsnKd51xZkSYpSor3sU/aW1XfZpyjmkjRMqh8KQBmtX8wuRsCzS
MS2GwckhkMNEgUFpNSBHfdJ4Z/MnEY7hPmocX4xNsl4IoHLgD9qXDpdh8Ax8DaMF
BDiqPIK1fR07TJ2HiFGJ5qGbRXT8sw6KyHr9n7n9/tJAdxWn1ZPQ60uckY1Oimlx
FUgP/y7GkfUEYnokckIuedvX/FkrlrpjvX5E71+NPg2baZBjUoYXvTlfWLvypkLF
3xJelpFxiGiDlPyHchc2Gk59I3fb/NloP+SNQdOrBmLANOdFRdQFlakqdJpJRwBG
e6lV9c/95kg2hkwjK7ah2Wl9+RYCHnQeDvk8U2xXQaz3ewRsv41hWQgf7K+fgsiB
cF7rmVoDvlsp1uEQB19Yyz2y3FuayMeMfs2qt5GyWDpyZ/MvLI5To1LV0SL1polf
GviUOKIPI0m/VTJ1fESapiOwFQDw3TmFpgK4v687I3iVzNyny0SWryC2d+oxO+12
2IzBq69qqXWsPeO/BXX2S2JFx3H174UCzjri+/qi2hVwcjPndwDL+oWkms1/U5Vs
HV/PYvuI4hHghrAC/tNZ24LDVN0gli5z0F0toF0vThxuXyqU1PSz4Wac2MExpJtE
VewGo/W4PNUt6dEkZyph5L2A7A29xpgWiIO79JIWrQ8VHax+FBNEc4cdp6AIaQVS
HLV43/K/629aXW1Io7G0dBpAe8W5sTGTtE8lzDdK+RERr++/NvI82qrpQk0wAUkS
9Yoj7VAWCRx9hNGGxa/OKgp56japa8TS6cOL44vjGOmH7AOLpmxJPCTpQzp8Lpmh
PhKHuuBt14qT5/6ulrkoWWHjvitJd1YtXDCl4Rwi4hyNQtE/w7OsSiEOHx3zpXNn
vYWYfU9aIdPiIe/oUMFS8Qii4oywpgdL8QveIWSv6aKr969m8ZKSrgS0HTe/IOSj
Q1VO2krpmBAg80tkysF7NTZaTbGcfDp9l0garrBP/2MwIqZxYM9roQVCXvbMg2CK
6s8h/zV7TNp4GV+aLmTFUv9/WW3SvKz0zeVaVv5cxS/wyagzxgR6jKTz/56xIu9K
DVex7svjpYiu3FMk/XImRvza+yxDu75eyza3qyWMia+Ko/LxqcXX0V01ONthcrqN
TCznKXD+SdKpy9IUl52fV4AtIati1VdTUvnAiVLaKTHPzZWxr09i/arWeIECkfFQ
JvEk6odewOz4hNhtE7hzSLeK9W72bsGNZwCvIk/vTy4eNdOydrZgbtnrP7r0QZsF
MewL7q5FCzT1CNz7ZkxZoiFbh+0BygM1BiJItQFwRPIf8LcuR1tfPu95Ib2vTvcj
1rp09f52cxcjwlA1pD0JuXpHFWA0jVzWwl2gioh+4rLuhZop0FgKYQuH7dsoEkCb
oWBic/YbfantsNc/NL68h8D5WkoJqvMtUSMFlmkfDnuaaWs5u7G2ogkwfMgNafoR
AsUEH6SH+QNB13mspxuRPduUBuboPtP1umGDM0anQZcPgG6EShhniX8cTB7vI797
iqba010f6HpOtDyle3KlY3D83MiixDKSyLloUaAdjiOVvpXy4Cw0VA+1shXaKK2X
PBpULUSaYZpGU8IwjQ7S3ZtxDq7nciCHENd+QJkt0fRtpvTHE5KiK7I5jsHNffn8
u00zbWlWGVDjoKV5GXgt0/JdiDtzWHrH+302Q16dNEblaGqxnYvIh8mz/L3jA78r
4fxJDV4SYZrXfLk4P5dfMZfO5BWHbJ6M+QDddUB0hZxqnE7YGSXPrXwHr+BzC2Cc
HykcWkLCZC9b8JEl7tzbCQDV4BDoLOuaFgFe7TGPWVf4bNYCG/2fJDROPHLp6EXk
lKJPTzDNpE0ZCe5aV2aXq+vf5MfKbgSPMRp8H/VNRK3xLq5fwbNEvHvchc44q4rM
hu/K7OeuwnOsnWSpj1gwBQ07DLxcdJQ+gvK++BJzjQ+jDulm31Aviu0RKmlz/Vlp
PyvJirYZgcBDfCQeAGlRbafgIOyIlOlcZ7Zy5Zv9xuuh5lAC/KekD5LqTD3Yjjam
mhYoA5onLziN01kFaH8v380NqAbolN+06AR5tuTyKe2+NmgvhuUP1b6O0VQOBIdj
j1zm87mv8A6UiOLhG3eGtT+dYscvXPZqwFe7eLD+83QNyucYc1iaw3FnpHBrVj9A
OmAcUQ27xKlfBtHdusR4og1sXnr/UcyzUfZPnLHhQtBNeC+fUWqhotGmbZs3c+60
UtA0wW8ArjvELOt68UNwBZPjWIAboI3Zy5YrUiJrLbOjlNyGaBQZuDfQMLVR0/q3
zj5rBqDPC8DkVeIs3yme2cy0P0I7S+DpKamsWwAWsX+f+NxGerfyv4audGa9g3+u
xnDPW6xdKSRnnS+gP2h9IjQR7lXTCr5hhpqTpzjsEK16BnOidOvaA1drIO7RJ66e
z0TOThcyC0vgX2I10NctkL29XOIIoL0viY4Np32J4vQjU8V+KCqeHIIgVZiEyudv
5SeSgQyEf/QkCA9M3ZgKlSsgavZ8FqC8NSPX74jsNwSDaXRzvFSvqxHRG3Sg+obt
TOgVfUMgNUC2C9YAwoAnEF+eSqq3UA9wBwaL2JlVznBBCGjSIiG5GVgC8LKxLzEv
WeVn88E/NdiNFRQ7RvCPmmouYCxrOuW+2wM85UJxFiY1oHnzGxcQsbmQqQdfoKH8
/BP84BOAxlscsjBTAXSzj41DtZKDwJLGOV6uT2wfczLCNcVzLh09j63WDNQDhrDI
i1vu4BlXCBlYN5vHifXFfijEnVrEmLJVyAbkAjprzzayR8stp6Bz7Ggf+GZYkJui
i+EkOJHdNHVhIVGDfYwkwKMG/SCYD65vE7VrnaULwDcX94pXvueb9quhR9TWlZb5
mEYoW5SesX6BYIjCeAsj6CVn0wxbPJ9IJaJEg+ySd1jTXSPzbtG1VqY4EE5a7kxj
vIrCGNs7htXKVR47/k8dKaImoa/t5K/aSiIDFcmImKj64fqrRuJd5DjV+U8mpjgo
O3stKwc5S2CSqBVYSYXXGiGcDwTGUvpOis5Ede6A1UOdyFJr+PkN4XwuY6Rt8MY6
hM3/hbICFwG/mIg7e0+M5uWyM/BzsNbxmwmKGX6JNazoMxb5iLSSUrEySW9ArK4j
FapcKpfYZitDw4vrDrdFdI8krqJNQ8hGthFqWMotPwv9vvwD4Oa1BJkuKcjTtN6b
QsDgKkohCJpzRtPC9heE5yJ705aSssJTWRgNUt/461Nbgu3N4L87Q16Qn+nYZHax
Vz82Y3pNjj92N1wx0TXlJWsjsa662N9O2SKbivqOzuUMv7iRP3GUoRAokkxphqJQ
+WIAl1yyJjhto/uv9wuMZJq4H8MHDtDw5B327k9FcPpB3BK7S32/WAeO5zFST+kD
ZXEa9C3K9w1cSAMeJ4O6ly9wwvRs5pBUaSy7/sljOlhD2PKgdo7rXUqdHZWOzzBL
4XPHndlXxI6n2lcKiisvg70LIgbjow91j8hNfwrtxbCgNu1/Y7z8RheyEIxMEEeo
KAjR4mlHMLtUOHYcdYd9pefXY1Mr0MzBNKYSKPowgktdy3/tC3vSJ+P88Uv4aT0w
r+JvruD7qmJ+zZmqdcEujoo8dMueV3S1YD9oUWFrg7JF+3RvYiRBRIdZmseR8pSZ
FBOG0fUu+H+F5DiXjh4/WGNQkAR3NdJ85vp4czYwasJLInzlnTNS41CcrV04BOf+
f3QyjZenO4ZcgEJYAByxS8Z04YwaUB5PORkwmP8g5UZsse6yoEzX4wwKMxjYM637
6VbQfUjpNm9ScGNUBLYWOqu1UU9nfg0bufmxLtIJXlRICi/Cquoc5YMt0DlzyBaV
IL9Vac+/ZIulyFadGNtGzANqw2enMj6cMfiZTVYvCNXDOsuppzEMcU5H0yttseqP
SyiAioR6vV5uq9iecePH4k8R3hUp9/tsmQYD+f856+a4msL0GDnTps4n/g+CA4+b
+bwZH/ltQ5e/jLSMC3FOwO1RBhf8B6KFQudpF6ofFRa8Fp2ieOWyyYu7iETFcXyz
NjMPjg3jXkPta/fosg07eJVUPjWthW0KVL60pX/fXeV+YHvWNjySzaXy2FiC5+uv
Y5srhnjf+ZEpUMTrN4fT2gCV7ZGEvmgoJt1gpTCbwd+jigjfUELlfbTM9q1Ad0sJ
cdV9Ib651PfIp55F6wHKtwnfeu39MPNb4iVzK6mws7vA86OYe1pE/nhlHkUfOxVr
T+e5SkFHARsz6AnhwlGYl+eU4fIxVDDbmVPq3UcY3r7gamEYMhtKzxcW4s7MAZZ/
PjFl5TkKaO6LYV09rtOBJD5FX42WYBPXvJXcHrI7uso8EdkLGL3bBPBRuAss31Bq
eeG2DyWe6j98jRTNHVxfrFVwoKAedBIUHHlI+yfU08Zg49XwKI7xA79w7AfgcDFK
+hNc6RXgdbAvZ9MZk000QDE8E+6hmsx2dQ7zXLI/aCKi+/fgR+xLONQ+YkdcS0MM
DCLQMx/Dezl67TNZsvY+JX6zGc25krNijvm5owVdFT//kIyAq1lKAtSmHPk11Url
o435cuzgxNxYMgUjNVZkduJXwmxQySsbWuVsEZF8A/d43DWC9UDxSXtNghQWthE8
/ZUoaeo5iqNcEqWAqyAkiEHC6Q+Tn6UyPYdFD45BrYnHu8xw7z8M7RzjSjrUWV0K
6YRvPUWyP3KiL6hkqZTUGgKGRFL+Sm78eSoA1D22OL7WwqJQ1TIaJPGXOthpAemz
YsDhlpeH2UmoASA1Y+ubK6jy9Ql9kAPzUk8ZuvMWvkWq6FYn8r7u4hMVIwPNTUVk
gQ+ucBuuEPwPohqLSV+lb8/bnQmyazA2lRlbDSf32+N/xdxQ0XYJ9jaDQ+g+ToBe
3vnsGmRgtno72ifuqV9YS6I+VxgB/H4Ni3UhE2YyMwQnqp4HWSv99VSAIJG6lus0
LWiOCQxXbMlWTVNg1tcXs1UZNICcRfQkPKyhsos+I6oo/zkfAdWROz2yc3u2PZTj
jUz//EvPcRk3ApLX/WgPgxWV0qVw+LA1cdFmaZSMLiQbXIkYPDvM1b7zHlYkG8cJ
ZFB3y4F0DnlHbWdXAFl2B2Ftf8jfwjGE961dUtHy0mvXw8CckkvK2JBTGlAsjBYR
vFIYazHlFChXWhWdH2Ai6fv0wViEPo3UoldYPLqyVLnYzm/84yeytmu67kmxUtrF
7vBLprebqF9cUhdwJLjVLMdCrxm4SaacgeTrG59wKO6ZQGg47iCzv1Y1pelh3mkF
aEA0Bqv/E71BD3royYxs5bVuvI2LW8W3Dnx2BK+i3c/lQxqDME1MpLTw8qFYQVtW
pS6cDvTTT7m403engqjvR/IPdKE/ZXuuihDiKM2l9ySPG5yXL1gRz5MEfFbSYYDr
/jc0PaXi1dd9vq1cF7cc0Rjsk7eAknr8tg86a3L1xu6wzJHG3HSL7UV0Xy1YqpXL
6q0fJKdQwzrF8Jm4P56ikOifxsyNsxczpxigY6u+xH6y00Irbjbez1MteQN7rQFN
/XuNX6M40cd3sT7tNHML8eGChedYv5IHqJZWCsR16Gen83AwTl5jwGsVTX6tFDgX
LJoY9+zwG4il77DsbVzibGoJNvPhp5fDL0yweB+n1CZxw3hKa5X/YGCcludb95CP
6FCakgIiVAM1e1p75AxZlEJBR5z8tl4cFesl/ckr80LZaKkDRQBOx7nqxtVpT4ki
fo1aaxVz81imCyHDq9dWhC3zL7/9s5qHl3GZTr9H3s3vk5+Gcx+FtTo7nrwXHv0E
dre1mpIeOGs6wNV9WSkvpZtnEkBy/FhbKKf95r3wjPZvz8WXlxsR6rWAt/lBeUKA
uuDYs4PFgfezXONfweNwr15SjgeHhk7flKChX1BhXsmZ0T70PRwjb5sRNDPmXI+e
cHxASpWCVlXqQLQm4BMw+aHT6Iwgo9dFcb/xwNBCk0l8RmdsXl4twRMSpZvXIaWs
pUugVj6kQ7b4FIC+FkGQByDzfQOUYtTp3u1mqX0RJ11Sm1ZNVYTTZVzFr/1YkzIy
wxlfGpMAk6Z08U/ZPRXQTEmlKMlFdqFIf5aGXYRTj/uAxHl/iLf6M9NjnS3WB4zL
zuqZnNJxhDdlHJ99ZQQ2kU0P7IlfLakqlEsmmDS1dNfedqH2bmh0/nc4yOnti6K/
NkKxJ1s2DJFQWnWA8hK2Zt05JdthipzSF++70VwrwaD5b16gm/rd3d75ViX4QnrD
O99YNnzbYNsWxyA70oRQwyb1ANX8OadWXc1ZGxKct2sSZupPpO4Z2z2r7D0VEUgL
U8Fp9WOPvb1F3i9hWFv+Wclt0zICtp5rAxyhfOE8bVunkmAX2uqedfJvqHlQLa9m
Wdv+TRPXqkOFbJHyj1HWGFAC4oBPbiby/3M4KnBP6eBFbhaampQARYRUTkM3gKOu
JKgxZsMSEPu4EhcgPDky6D9gk1j8xUG6XmkCj2Xsmz2XisA+kcCUqxi8tS7zxCMl
TeLHHYBiQ/PAWidCjTJEBH3rXYmnHzGuGcIrHC32M41WIYZBOSZ1/i7Zl98XqIRb
gJgb39HzAXzB5X0KU/Tr8gK5GApkP/IxV63TB8lhf++FLulNc2iIfRUKkebVOFki
Myg2TPlgJyLV2O+R8hY/+3c86b/BskS0ZaVrcVRdamavZiqz6aXNdujTqokwACxC
vdCZR5WcKGVZMWBoPSxImu0G4tV7s9WTUMgNlevaIeIh34apbsbi0PIJmaWiANyx
w2Gbsn8uIEBYX52WiORV+C7uS/ZnDkVXFPY6rmG6SDI3h2QfdY0RcpOSDFb9GTx/
3KIBOiHmQTOk8O7bfHc0Z3qfbIDriuRMnMWpFdTtSASLQyU+t3G91uFLlxoIdyEJ
xNnZvR1HJI8YO/PjjorUxM5Nq/k2osySEbHDMOnWWGj9NTVoz3uMqKKAOJAagCLH
D9vvs/sf9rwGDWMFjYvg0v8DEBZYVB0HR85amAGwctjdpljfEuNu5rdFO7uTOmBN
OFXSby2yXJeZEiIMxEZIDDWSLPg09WMnbUKL7tYNpBMUpvTjf0i7ww6NMOeR0BFh
Q0DW1+aaIDKiPR7TLsIZC73+kmrvLe42V2vbpQkRwW2Lk8A8esGvyBHyzBG8S1Vc
J8opqNqL+09zJ+j/+uV5H6maMl4k5faGtE7wOBYnq9OqZRNTRhVAkmVZnSP4PbU6
g7i2TbB5eAdYJGeTPNNKFUCMHbDJpROgH7BN5w3aDaXULRknp+0hkcmcrzfUomCX
pTElLyU16/uxH6UtqneM3xtRy8PKr9r1xVdTu5BhgEAy2S29k8Kcv2kpRqThKemy
gbb1Pk3M3shqQrW8v2I62UzZXR7rDjD2D078zTi2NMORK5EDaZhXB8VP7KEsmKxU
UlCzFTuRQCxOuGia0p843DwgW9KRW27aomooH0kSAA5aiL5zUqafQnVh2u/DwFKT
4ClLUcqZokzIO+cKU9S6tTz5RE4bIU04i8jdPwXf2wZTqjJ3904xoIbRxlGdUFfD
j0tviU+9TtWVmMJ39X+XZhurDiBokSWuZQVFX1tYAWeevIsGYkeCgYc1thq+cjN4
a+aqBiNfyCfHGlF07iM3uni5yMG/ClFPTa77/kJ52OqntYuGZV13sJFogRKabZ8m
WHAXrOzInQ5JxPpNZPweRB9FiLVu3u9/RLs9KKvcy0hGdxmqzew1qJqZbKG2Rnfc
qrZ6y1EY8OWj4g4B0oFHQVkroZIaCAtgu8A06jScLEvoAasN5myRD5wD+/INx77q
GUZ4jxDNrCWIKHYwq9A+PfOSOJbFcfvBuyrPhhi6SdIe/Zn+iouT9zDTquvXWkT8
xm+p2jkgJJozdu2/6Q7AbyukwK0yJsySi9fD95nf/NMim463suAwAzKe6Jm8J/Rd
KIwjofpq0o+pIyQ4g/3GtyuX9XMAcVf+/kT1Ek4ZPMEhhNX/s1iY/UhBZhbBzAi5
bvSHfi/5zzCl6MeD49x+EfIS6jQwQaxf9J2RM+cVdmfztLppUNyK0DRbE85ISMaL
x6uc0U+2upbxFvLWCukFtiS21mRhzoTGFOzJYZumaal3NdwAh4pYPXQzQfiygbBK
A3Bs+nPV83qHCxOUgE8MRfs29fduogWmjBOWaXzxt9BxeOcftZ0RKxrpRBj2l0v4
YtOu+XLnC6X7ncytIUbcfTwKCv+Y7TzPDAMgtPtKnjpi1c5HHX+//rpVordPgiKE
b7iYboGOvGcxUM1z0xP36nrSJSDri6DX4Y08S5rnElNpkxM0lJE4mOkyl+pjqpPJ
K/DVeUPBeCkRLUXkcm18p8dp55G2wwSkAJ3fvH1p9MCsk5fHR5tKs9p3BHZ65eec
AQycy/ef4AC0EWz+lUF37efcrUemZ0KH8/8wDLQRtV2ruO3u472NfKh4zLQ/sLH+
n1ayA4X+Rr7WPmn57Q5A1xV/KKo92RmptWp6Jkv5ITO6bk9lhmUvqc2oeAN+FjhL
ZaepLIbQssXfEVQuoGXW19NRvGYV9qNll4WaJI/HMTvPwQWgTzG70oACRwMijJ2Y
TVVsUrd5ppaUZnfYUSsnWMZ+qgCaZsOw6ioYZ4QDf7DQ8n4+3/QwskXureFNAy0q
kVVk6nahLAsevZsfodquJFhYtmr3WqPonoqC+GSTPje32K6eMew+nZnzuVWANko3
u3NiwKqZdfb+Q63zg9dq+kFC7sZrd10pK17p+R2vmZxmqkf5Stq8J0rTmIwQacxM
CRM8hn17g74H2+oCLwb/llZddYFVP9faTkrnbEn7kc+cuYsKkA11qU7z8rAmY5Q0
Eaze9YNSSdwPrw2SZVNUADRKs1Lr94Gdcn1j1RSHvqfSW6LZVS3Xp20omiNGpaEH
PssCsovLUFNJC5joBESfIHukYzfKLwOBA+ehMhe8pTz/c6ldYZOWpsdsAQASTXQ3
6AYJfDIZMYhUMqA1CKWik3igHP7a7pk1M2jJjwZJz4lpTTIIXzVU3OMHxKScUMiq
2ejSPl4LHuXOjtDiXt9gx7ZgaIoTqU15YvREBc31kr/GuiubFHBI6nwqO8bO/tYq
uN2LTOQmEXOveyZ5z4xFXXEdWENVvDzm60JYzAnmgi5mEoOc7DhPrqGN65lW7AY+
zGYH9qkCPOn0UMH0JmclAwTeppAz3Rjadg+6VXCmlULiWyvgL3ou1O0GBlq9y1bi
YL4Z4aERMYlGynrGdMJ7LZN5/RmHAPeZ076vkC3AvjqMV1wWTWkxXm0buHRHT9oB
//zb/yuSNpGZClA58QY8LsAue+ejQ1wKrs1YWIhbOMSeVOPgNOiVaF7QvXSwF8R2
blu541PZkE/str34Ao8FrqeTXtzU12iiF1ShoyqiJ0ZQ2nHb2VAxZCrDPdHFI4es
3/9+8MwfIKlzbKV155FaIySwrs4z3g3QH0O+huNUUVvIwvaGkAq2UBdu1cF18rA7
2Ez8yhKmrN+Fs0A4j0DzYVcArg0s4DETadCqbKFZPyTG4z/aQFnoCcWAKRvMvc2b
eyGtsdwF0h+yiQIfCI+CkOOPqQi5ZyIQOju4LPe3Yuvd+bhWtueaqgr83mpUbh/5
bJDlmtwNdcjU4m74rnS7TPP1Zk3gf6J1NJJi7AUvf33BvL8y4JgPJ25L0Oe07EVs
qPRrGCcMwnUjNL8yqSJh98erUf9dBYwO3aYy7sDnfnxIDGLNuodIEgU5HrDfV2bQ
FFMs2w7LEiB25wfzzg/wTm874O5P10goJ1Tg4HVBP59AHKXOe9I4Hc3Ra8xkGyf4
lW68eXXRpPHX5jAlVBwhSIViOjWeE98YjdFSsSiD/8vNlOH+oFHkNut6D5AGWM2Z
ihYjJtnKMiy7PQGD0MZR1cd9O9zAP4eAMb7E0k1qDqqvy0uqNdn1b4rZzeftcboN
VXsJLS6MdsDARBuA2QnIe3aYkb4TJ2grNhZrqkPt6KhU3iJN7GZvvocSgDzpCLjZ
ZpcfMrv71JCzLzTb6MqE8VHwiS0/gDhMFweop0jiMNAkFzgW9WtOHuPkskUmaGaI
Q+zuQFEsn7AgVJc2LduXrloH7vAZmuCEiagrQH5rWSUsMvFR5drS4Mo9mey5HdHY
R5IXlgW7lj67h/l+o2/VYU3ww9UQyULtXtY+buu3oHjRF95AXQxh8I8rJkrKPBs+
W360Ckf125MhzyQdvcaKaP8hRQjLFK5nYwk7TkT2b79A9UYeCLbYN+GZH5rrtKnA
wTRE8rsGRIYVFKjBHuP+yMz8m+dj/EEaCVpzlC4o7/Yrk4hcHwBxKuOylmkuTG3w
TYGWuvsi3h5xmRThGY/BmDgxhm/gP9rFKBkR7sCBv8Dil6dIY8Dkp/8q3M748pIc
IkPSbp+NUy2AHZvkxcEClcDd7VCbEESNudygp20GqOjQKC+u6q0ZR1H9JYdGG6rc
AbuAe+5nbxysa70RfMJ+2/OGalRTpLd4T3xm305R85fnxkhPnSKWJUKCCbPoFLFn
ua8xJqC15HNbv/RicO+b80Wkivo5DtF3RFRutmTNarsTG+rYmTO+i7GPqf9BRAUF
DD9fO3OUC31ZDvavtTmR0H34cH9em9XGa0SxJDLUxhF175ODdi7zzhf/u7GJz8PS
AUyGIkgY/Ly/78wkOOGQJKLoB0Y5H/0K+YvgWhUmxenYSN2/LfXvfocgQyEs1Lqw
VsxGhmREyYJFduKw2LVxtvqqIfkTr7BxljvUEo+ejznPD2UE06+7zx1U8UXw1Bgm
ZS2986eqY10MYe6DZj3FBRtZfw8FgSyywVOXGxbsLRhONZS89QAya3kgPlnUdtou
RcjAgEAtmLd/4tXWQHOtUAkwgR9qjMXzRroS6pes7o0hevibnyyR528L/5LgxNO1
1lLlCKT488shMpEs1zpJyhFM+fNiKpHIBpN9E2Ed+ttjNlt6i844b3Vy2FZAq+FK
6YhwLHxcZP5Wr8YWN0zZjcsLveST1+mQgFT1nmzQrlZ++MHxdpZqTcRIVFdQIv9k
hWFtZsvgFV+jhl3pldJJli5hk0KqeMUPoyUNYIi0PxU5HGGmzq1mkz6ksL2gjMQZ
TgcXHh2zYo+QgkpJ7MC7aSQOu+f0sHuHcQBgvb9hTEEnBkp6GZggftZJbUoby14e
kl1HFutHviEnZ53gJcSGbDK4zp8HpHyBkxyi7OJht/VLx914c5XHzzMvDFMsy5YL
ynPdZM1GH7bSGIOB2LVIDgu+JiI/vyfzQypuTBVECYmLRHlcqhXsU4vIVT/x2KIo
MBMNUk44NzQMiGv3bIv86ZagT79sWMEZ8dYAxjOM9X4VPykTrRVsY05iVdxeo5u7
WE5ZBfkNltJM0y+EUDX3qoym57zpAupz3nDdmLi7gCXmpHRg3/UnhBQEosk5CtTU
R5+7b4+KWU8ntG+ZC9Hk9XYgyeCt4dA0UIghfnSi0O5BH9yKsFOySHrffUjqs9ke
pQ/nF7BrTPBhkEUGhcEEWiNJ5PJrMkb7xIkxiQoX9CdcuktSkdHB2EpdqzGeA8P3
+AOF2HEOSVgWveRPUPKSqUVD+tJdNnLzODfZub5zx38PtyzS1vB4JPlyft+vUvYX
hIc672A4vefbuYAKY4m3eS8h4uZBB570u2DTwpwFvUiowcaMgfiamRzEJ3KrzoTH
l17EV/NU0Imvm0R984XXbyDNOt6LBg9c8xgw/MBmSLMCR32unnVCjFiUJleyO5SH
e8EY6bhJuH+djEEGYaYRc2FEfE/YcwkTKR1HnH4u3BPcfqvGG14oSJ2TcMMob0Ea
i3XKJWEOnwgLizIycfVdRY+R/FHjIlmK3/912ySdthXsxAzy01w7An9p4dlq17tL
L9wGQ5lkb3rghu+f8cOWEhy0p3BJ7RV1pUYaCWyh5CGxRxh5InqMfwnCrU6DqPjD
Nif+yILbCSU96XclhOpvqiDuHu0omsI4xirl9Y/JW0M+LGBm2uew5yc/nYx0ypbi
98719dzANd582Mej8mVltNQUtpB2U5uhG5gDNYjzORtig7KiEyBSTP7ZFrIN4n2w
oxXuSE4T8nCZDYtDH7W38OccA0brSLQ/JSh9WSfbICmBqvUNY/RZEK5+6hkAUxrt
cMCSgG/2fD98z0cRPWp1RpP7tROWxLAJrGVFFvEKy9xc2LSx13H8a4kXSlzP8iA5
EFYzw7qMCVrDLfIDdx1GKDCgNqGhvx14DgG5UbfR1OkfS0O5uqgtYT86dnA1ve1S
O4buW4UDvh+0iWch4Dbphqv6o6sw7oipIVCwC6MQfkWqZx97a7XXSrEFocRaEmbE
8R8hQFH0891wvmHpx3PimJe7ilhEbjfXmG5ZFd0+y8BQdMG25+gLvwBEdE1UWeQ/
1loYyh4uHYZOiO0ICBwiEja87+0hNRFKe7nxxwd/7kbzZE3bbhVHcSFmsl8djHZN
Rik5WLgJRA26j8+XJox/q1mvrztOqg1DHfxO3vWXPMa7Kzym8Gcg4z7tnJq0ZA+U
8yL8jIO+G2oGUZvynfwdr/Bm6c9B/zdE/iJa0sMNEpWg2c5NDK+f5noIUYFcqRmN
d2QEU8GWpXKDPNP4I8txFw==
`pragma protect end_protected
