// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:31:45 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
lfsZyWKA+PXbPQhy13TS/pjJeD1o1/5NgO7K7qYIALMYj4gI00a/x9zc/K1kdh7z
48+moI83+l1uH8xL6WmZJxWmq2xXbm0pU3ww5zDlBZxBXIhPRFZmTcYklZdSDgNF
5sC5Y7bmVFsRqseNIXbb1CNPFIg1tECC6SIkl4zxcs8=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 4720)
j35BAAuovqGtnrlzfs/3/F3Ee1KY+tryZvwz1ORFjUrT7AbrYwIs6D13RCQdXDzo
3/UPapaRRF6m7FWUY1ksdPDfl0Wb0vPrKN6n3Jf8Es9g6fX3M9EsY8QS8152W4Cg
YlGVXofytt6N9oGQ5zo5ZilRrFxpr02u/0Ij1zKhTukjF7aOzqmn12uQTGsoTLlB
Hf9RJ9fGWyyH/rEMNtYSZ3Qsct4KLTRIpAAe/r1b5QNmhWHGmqjnImGMciT4l0Ry
nFVappUAziHvZgS2oNutDId8F3rG8Qvcaa1zxJWKTrxmj/bNm4FVqe9QJ4wTrk0b
JK5DRILsDdry33V3M8py6UWfWsM/9rvO2UqTbQTdRFkd8hAUgNbyAgJhG0eVbzBg
IoT4qOQ6MfCoQ+Cf5W0F2p8Nzv3l12WZw+MZIiAuiKRhXhbyyaHBZbGYutJMAWXp
aCEd+MXDZ+GwwpImlYzHs3qZIwXFe8Jf7lhY2jOvRQlAhe6yDI38qwc9fYdyKgxR
uBsj6B0+C4Gwusyvaj0d4BmJuoYLD6tNuGrWDJnTZARMrs+NuntugH56hgh0OFPD
Kv7NqEXWET/Wjf3LY+lqB0xULTf8aZPgdMev/VvWWvSsFD5ALZXMT7e0haKlf/2u
7IYnTKnugpOosEbLody3zwLJuNp3OByqj8jQu5pX+lT9R5DZFgStPYy2AKo9vxmY
637TDGe1ngXyKQYl375obsqNpJrCotQdHtQWiiRl60sluzjO9C07/oIYK4KUTAqP
GYBrnUntiysRGiNE3G/+HxM6JWH20v3aoRG+YUC4WMn3RIFTJGGcawTd6Twwe0k8
qLD3mS1NcMyFS1WU7rKysklM4sZh4eQ0uXvcUn/NRMIJNHYKTgaYozq9HeT/G8Zw
JeC/c486rWdRD+SuuFLFDfapZK86mNt91Gf9Vm7YNO9Y/US2m1yqsk+YhAOTOziy
YciSsvPOSXdBUU0B2NzhDqJdbGKipyUItq3BAfs/nFr3JHhbMh3fg48O8Mg068v8
wL2Y9BssgFcxBAKOB6RfyRTBBqFavCsjPxttG6OBO18FW1CigbqZmRptQaEpBC/9
nyCaKnO2iud+VbW+6VY6FKys7QGmjq4riz4gUOpTsS17GPWxb38C/jbdeEE9KCEw
MQi0SAzu1HcEXov55vEv7GeDhMT1nEWVJ00tMdVAEB7OhzuTOYGy0+tcKvzEza5H
1+kX0vc+cBppaWbP0ZORbibLo6xUDV5D7gzfB/H/uMU5XXgazdhePYptXIy8OQGt
yfpHLiRxtk1AUQUu4zatAEsmh37dGxxLZIlZw3LCxzkumhaxJ15J3N7KeRVmZsZq
txKs66BW742fEbywxzzkahIXHkTw23/Dn/i0/81hh97a8l3DEun12+o7mNkh7cix
JRy4nAW552N4/yDZWetpD1bacy+n72E/vNLXG2YsM0t3K+SmM1jAoAqSkEjH0616
81W+iptagQtgmfUD2+kl2L3V/SUAivid1/uPv+n/iKMM6u/LUJlXI888qJr+c5nE
mrCZFXrSi0THWdCDTP9GUGyVFS4+PdC8vX2+jbbG9minhBfIYdaSaNDwGlIto4yj
bnRS/9cJ+TYKqWhcmhb7aPZwtDH5vGDZKz/L6bDJCt3QUjaP1wmM2hQMVRXRFhew
52VFDY3Doc+ak1UNcfE6nBmUEAnyLbQA8Rs1uBwfARixXcKQ4+i7HhTM63qbBut6
jzE9ZE1NXcnKURFLzLJKH0RkLBW8FDdX9o7qijmPgkyH5WOFAF+2dxAP0wuLTPVO
zq48bI3GUrwo0SASU4ZB3s27OlptgV8EfSBlOLCNmOPEie5orwrHiONChm+xoJzO
Eb+e6gWX27PHVl78ua48ylRYD2z0gyhMlKiHLRHiFkSP/apaC07LNjymmVc3Fzus
Okvy7mz5dGucaX3iezCP0XjGfNj8BEZrGYbYcziEH1IYR2s0BHKjSI1TsGssSmKO
OX8DpOL0yEULj16Ma23SpAliCkWip0FbotjCgv5Llnl5qyd2DG+u8bTofkcalFd3
+v2fGBXetw8OfwtLWv1QQYi48NOKWCMIfuMCFOUPKAl9wfaDHzWDN6/c3bxLwaIP
jkafiUXPyRQl3+ga3VpU4OPN6yMvOg/x8mgxJeQ8GckXpDkSYCap88ziQmzGGHfF
FMxtStvana7ZYN0nmoFhdesbkj3rJoAZViDWx33dtARV9ihl1fhvpXnTalWGsAVw
PNyd6omThlWIxwpFkJvqd+UJXBdMuhvXhclY2ZGUqn7PcqY7HMGayl3TUQFXkgfp
k4Qi7+Re6IHFJprJIYWduZkYM8QL0DDKR7aFR0zS1rmrJt7n7gxpG7GH9EjIUc7E
D7rlQa72ldvoQ4hyisjSkTBPz9yErvs9+YEVyx+HQP7v81Il3ymqBheOQr0LXfD7
owwHcNB97pVsKbZ8r3bbXbxF5Uyt6hAKMb17OR5pO/jQNaSdIS33j0Wns6cqHQpG
ABLzT3jH80EvLwpe8a496Hu4bP+ZsUbRzThg03ZMW/wGLMw1bZEnJKA6BVgpdN18
nXdU8sSG9r2/DObDSyopqUU+4+e7V+9ffDDacoLbddXveWp0BCi9doLdg2WWoazJ
1RoF7tzdRbH5wuYGAWeWmfHNv9QE9BPGa6c4WoeA0nEu4SpzBTBjg4AZ0GX9Fgfl
bOcQLs8LiHS6BGIQiTXh25jKxBhlO6J6RzUUdrStqTkcfNW1ZlkQpsCYtcAy7LTu
eCH3Sh4pn2grztcUPVjhfALHpyG2BkgWYx3nRkHImlT2O2UKypMJlSQvhvzctpG7
azOOo+hxO/MGLGg666g6Ttjtqlk19MkCLChaWxpy3mpvsnJOozCnYd+LWh0aSkvx
JEEFrr6gVRJ8hSqS+RdahAmyNMNLAp1aLiOx5kwTu1f/GN7+Yp5+StsaOXC6TMCs
5SCLBiz9O+6bCfm5KPmZPrYgMVP/cxhf6ZXk2A0Pu6LSaLDFhKOo1/+BFmWwDQKM
fHcrZ4y1cJDJYFOnjadAbWxAe3KfTsZZfLrVgiPxjzpI87Ph98TQCDUImv4/XDwB
wSjzOHk/qv1XZWyeSaUzW6gUZHbveCOv2+IhWGf+RSpr6rZOsUpY/bPP932c8gyQ
u+THDyTydqLLYijEcPKpssv3Y8UAxCoQcp4hYq0WbtbBOzL0jmlp8KG4Ju7IXubU
o5xyUdUR9XE0F4ySReAsqpFu2EFpgW34bfbQrXvlu3I73oY06wleUhaa0Bh3iC8N
MIYk5HQr6xXagD8W2OondPs4QyWd9dtBJgZYu1cseIqswjCOexYJH0235gTg8O3m
cqp90MD2StxGhWEpxL851pWLE1Llum/lxUHY40PMg+4t/QVd6+WxolLKpKdTRUOe
UobNY/VwQ+wxf/84pkU3vZik4gg7lpxkQcZdtj6/CnvaY+79s1akHuxYZDKLkkX0
4ZmK292C9tLtprMR2nTxk7535PLYxTHGnLAWdE+H2GZgpEdAoqVBtlGmErbOeHYH
VL9Gxi1IOejlg3BhCJfqn0NRxUSgaXKGmINVSEz0giW8M5U9HmrNkT0L2i1rrIfu
pa7IOdeKStOk37OskfqAz8nU+Qn554a1njcpZws7hjjuqaRfu7l7m9cV/CDlbeUU
3r2XJhUdWMCiQjifYW8iTbtTl7k+yD85FpqzvgKGbunGO59mE8vIUjy0zxE2H60G
G7xheUVyO54Z1aexbA+y7H3fxm8sA5wUmFiCsEkDFXn9dQG5YnXXXo5gOnYZVR1B
x2ANR9a6fXVdMefMKSevAoIX+Kyeu1jXJaimf6drgxxs9xMmI4YiEuW3pAc0IKYj
gFqk4bBfZNOPei/xw0QJV5N7ojmT3lJ91cKHVRALOvd83nWIMhz8RwQnm/I6SWI3
GpXfnsIyBVeDAzpQET7277FV2F+aCU/CG/kdebp3osBzlgFqS2r+DfwsctZ7Rlul
J9SRxb/ngyGAjedr7SW8Y1Cj+119rP+d2MT2pZYK1ndb/zXrH/KUmy6eGpnQ3Qer
N3xm+c6s6D+TnvNeIMfw6RQ4YaIrWw2w7cPF+SEdPqJDPRdnKkWu+fkCjLqOpqoU
cfD113Tn52P+ryjOQD0qvpF/8IGBIj+fOSE2wXik01mJBlx0qJhiAl0LktDfQflt
ePodyX8yIIHSDaKPv+JqBAR0gh0EEuQpcOG8JuTr6+DHz02r1hQP7RCOKYYnsr39
Wn69fjybYsN2FGBk9d5FukWwL1OOKjowYRg1/BD9K70bC7NLK3hhKvfotyc6fJtF
VW8mRehAmjvy1qfxCGGLi0+4SxLCtisFaWHVi8uQE/1DBr3JLh01j6ogx4mzOjg1
A9S8H9MKdP6mLKRm6ONhS77OUrYD+MbU5mbVAbVhXGvdP6y/Ep1lpJbqCJ+gmKUT
Eic8q3Yr4JmJDXcKnvuP5IhGdtkWpNhF4q7ze05qTcHMBnahZbBWGryNXXIe16d7
H/axCUPmAXe1YgIpCvLBLkVDp5DeveBaDeqc61SiXfgQHFdvrMynYNbNey4OTDVg
XCT8BmovkQRj86tf3Sz/rd2AyTIHLC4L1a9sMy3SzCthL7Ql6YoKYKD091nrmChQ
4wdIYNqsw6ITYUpF4li9x9cvKi3NGtmZ5AGJCpMB+H8Lw3eNqYXzaCuIwgv5maUk
GDBFNfa+grkxg5Iv8Z1X5IR2BJ7WmwUeAR++fcX7bJuZc+j5ossxG8vFaRSDJjMS
GxaH2QJGFg/tMB67bv6SyT07yA+oAk+amfEY2Owa7Qar1tEEDn6UKSfoxHBJRNfL
6Gcz5WReJgLV/Et/h50HKNWtCE3l2NGvHp0iwAr4qlo8aJg1M3fyLy1R6Wcd0xUB
VEaTXHq3l+bH5R1pSdbUAY5ycjjgny0qpKJaGXbXBU9WqGGpBmMnMAXbh5ed9Tpo
xy0hyq+Wns7MpqY0I3/WLnfidBBz6RFFSbONlBNbae2x2gIFRsGnhQmD3zX396KG
OA94sr6Y44+xUNgJuTidwJWJYEYzI1yIay5eJkJhacy+FPe7kogGzuLvkfsB7gkP
NUgj5qMwCOrz6XmxhIcA8W1tYQg40pCxKf0mdHgMBG2Zz+TyhJYo1B5ViRu0aF7C
AvDJJpSVRbmvgH2hw/rnoIEcXMbQfegSEFFAqgWOrkTzEKwCn5mU/ICGOs+poGVp
YkA86MibC2adA4J5LpoJvN6WSOox8/WUFZPeu7LC2LUmoDTjq+TTmcatcvzjoJ0A
ek3LG98uy6sBXnH9IdkpuocPF/ZKJKDLm5JaV3UDOv3VUwFHWlBEBs7D2ztdwCEx
ob30G92w5H7lJoTZz1BwV+ZlFzWoewYmbHWKJVqutf0l4FaW14s2AueQFrbxRZkC
irVFnOPP5lxvLitQloknPsO5bhDuAdvnJGLIQrdpjzXdE3aDka2xQTGJjjsc1i9k
OUw+hSA1bkS82JAJF/hecMDw2eOpUeRAQXYeRAFeOV+KcGnsiqUllXy4EeUAm0ii
VtIps2QQKyWaR/O/ixgWKHZilG4pfPXFZ2TiURcLPrL2RYtk1PeGNEVh37FKLTFx
CRXsUjdBX4mHMJ/zs7uEE/tUP4EqauuN+b1Mhx9PQwfaPsXiUIlq5L6xIvmCGDb2
voMJTwd/cLBmmHYSTRjGmDS4qvt/ubnjgwroorSabIr/3jzhvZePf29l9xD0cHBZ
bMwE0W2gC3zgYZYEVUNHTFSgheoThOAe2cNr+alOU7zjJdWdGTgqZ/kNbiMRbK18
Cinh4AYFZDBDBg9lp+vazVaK7cWzTLvhuqNXR+WU2FieGgpCTDV0+1I43ihvMEWx
ukwvSNqfbF5wS0swOLS5ZDxFO2P9wg+C3p/RLsmKlaNMHlYdGjzr5j+jNOTo/LJM
Aeso83Ru9ZBky1AWThJB4UbYH4y/2CI2GWFPi+P+PdcGJzwzELke50B9SXBZno31
9xyX7HapEI4cyPDIenbde4kwgmEdlE4JoIbuFnOwruE+aW5fLyd23xQgIcaVH61W
HrPWLDU+GxkMo0DRwFq2x5lN9OgKnTEJuCujk89w6Vo9Tw7DZvY7SuV2+9QX1v27
ZvLLMH6VV9L815HXy0MV9tT+TIabc+R1+GNyuHrIC/t0qdQqocuie687jaBl+Dv1
P96+br0+YZ5Hhp8KcBhjotoCG7c8h/SJqwA6QaAYQpR9GUXwiiA96dR3VggmFA11
L9kHJ5gCg+NKmMbGX2Zlabxv/d+3db4dhO46O9rfJ/LjK5JoS5S9Wz6fziNEcgCc
xuD9vzMUDscEEuHFijlPPQ==
`pragma protect end_protected
