// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
OlESwwY0o378XrCbyIADnCD25PdzJaxEp95o9uPmmYid+yCxtEJmF1JiTNQEQvS/v6lNDjPbKAbv
HU4Xiz6ZEdFRIM/81W2YFcjAE8HkNER8GD1hw0079TolII9XHZ3Of/gKxWDMOI0WyoJFHdtf/yKD
dPp4rNu3S4wEUYj8IJHjsfXLH9COeoJSUBh/YeYkKD+xuJz2aEpyExrKF/nG4q7Tvoh/5FEZYJd9
F+/CSvfsALelPFXHWeYSiIqcU71l2jpUhmk8ayVXKDXe/qr+Mo/7mwsttzaFGPL+4OKH9xjbzySR
gG7U3qirCyJbZtslleVwY1va6tKpRWH9e72H/Q==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
WxiXz/Xp0FUuC2RR/8lexQMIga09liKM7aH8P6lP51Tt/WVWlOriybUT+c46yCjeLTamrf89TPaS
zM3sOq7afAEjIocixzt9IzKSrrpmNeAu/gzx3TnZAx2+2KIaSg2m0RYFUw11w4ZXhapmjM8FAByW
11Q9bm9pzUsVbvL8YGCgh5T6Jm7CqfOsYwt2BpOrtOEQXQjh+h4GH8v7uxtDsc3OBLHwcboHkLZk
+dyCN4gts4tZCW6DQFKDUAk2OfneqYycX+656oQJAuTBUgjx9Ea0EfbKVQqP5Tfnutxog6G1L8Im
KWPbnGo/mzGWf+DayGZX+poc0SySr0r27OK3iNBB7zN2BYGBb+LK5yQwi8jbnFJGMYDlobFXecbB
Ve+yftoR0SHA8CKloJeFFY/f+q7mNOIVyidZQnmHka0y8dXbMqFgKMwIDnW308COZz3D0G9Q47/G
lRpC6O08hj2/ugW+skxJr9PizXbpUPJZaO1LW/jvV/oslHr4b9sVC2vV0NDCEWe7nieJ1wVQh1aY
LmUObPkDB2+HgZzz4mlI7Yt55eCpg3jhQ0Oh9iJ91yYgnL8hxTZ1TfRVxbj7dmKNlIoSvn5+dQqi
Ojszzx9OFwQfbOf4to/qlLpj+8UwcFDFTOaGHYZ6/i183JE1Sv9l4+67FX5IC2a/sSGmS2Mnf59p
x4FY9j1rKdz9mZWCzlc+bdT8y56CqmjegJEMaGM+Sq37JdY4c9MC/1zUHUApbZ1ONVbGs3SedhnA
PFoIjK0ncL0bxn6e+ZAMOWX9MOms7RPUz7j0TvQ9fb9m3aDo7Z+rODvfSnGw9hkA+2IyLTRYhjDi
/g0BlBjNTCF+Le+ROXeFKN/d96NF1ByQ2XYDsem/+hYx/zsK63TCCK4seQTcSV2iFxDjw5n0iP88
IUdZ0IVlvgPnFigbDA8UoBMK6e2N7InflbycCLJb0Z06SdgiALbp3b1F/KbcocxReMCMDNQukb1o
W4jLpNv1zcMlu8q14sEqUYv3AT8uLdhMLaB9b8AiYr78xVXWL8aARnVxVah1+n5IUY4FOQYBzmq1
rc5kPATa69lkaV7tEC27V8dTycNVJs54fVbjJgL6vmE+/jYxsVOPv2GhhgP/ouoxiG2rLM5ZSmin
gW+TysEGVLw8bRT82aED+vkCkYRqx3JyYRXq2c3Lfi9cvwJkbAadH7XeTHUK7E+kdxZ8N72k8zuM
OKmSTmZZSfBWXN8gLT5Uy6G1J7IbNN1BpIiWolkrEXlF8nKF/jIfIesddmykJtB0InGXEFqfm6M+
0Zd8cQq7qQxGDW8GVKTx1XeaI/ddsVCAzldNWmKfBjKZ6A0B+Cx+ovbSSJCRlnVRALofo3qj+p3V
mbCFmiO3lJ1xFstb+vs8Em+7Q5S0/Y+PDMq5EBZiFzRahFCQJ++FC2gD+z/vVq1mzVFNKi8GD7bv
heqnvr+qLgQFSNxqi4SAlkLjJPFzkt4CQwOPRFqRgjsL0hkMBslqp6kLlP6TvKXhxiIfbt7jOF+I
uye6OPvX6AY8qXpofWpURaThZBBfz/agrkeYLE26GinJUaqX+D4JSYmnGGjdKpx6DBMce3Hfrfoh
T/BymtQrEXKx4VzkSXkbi0XJU+anaryIKNZwHWbeE7GZah9+ri7JyZWlWzn2QybcUu4cxbb53nXw
II0Yi/jCZCJU/NKqV2q5Q+af1JXoHLPGtZovPSw/AwHxsjh2h318ZcO9u8MIVqkHaiMYraAtxbq4
sUOtzkuzs+NIybhw69PlwC6hWmn5yHl5Lw9rZXqu5j8TaFKMFLdN6XfWWz2xqIj58mWJ597zxwOx
rtkKQxyqmPpoIGDoZ/VAs1ZXhJeZGys/QhUx29J0TocDmLOucemecqg4YDrg3u4jK6h01PQOZZcI
EdiZAYyUCMsJGJIOFqgGjL7oTD5zr1hmUhS22mPh0xyXojTbDimfjNdvtrTUMwpCoQjCMjawRl+n
NbBi0N6SEVsxqjguZRcgCuIiOfQPcccDfmZiNACggKhHz0BvJBGKZnRzAcoobGLCfCR4QJnYkLq7
C7e+XzN5qYTz4E9MACCPpWyVmLvbNWm+dzW82u4o9wDegMZa6cCzZbmZuvZXauS3+Ari4XXFOrXa
ij6cYMr1JuJRtyr625aYS3KMhVggsyqvUcO257Z/3ue+rkWxScBXPfHpLIktfOJqqxY2WWEPbKw6
bmLaFYK3Ap1ipikEX0sltFmk4eTW5o/uKoiLVTasVIRfnQemRa3El5yQyjb8IxAX3eNPUPmM3vWz
0AHkupl2eqLsqcKZOp+a5I8CIsAMMvE3CEinq8hxvVePN/wd2iA/Z9eL83A6j9ZWOzTG/Izhmmg/
hCcP54OdQsV2rLsJlRMPPuEAMaYl5vihXQM08e7IS8i1KXwv+Thc6JmC964C8aAKXGPDYy2bdsOC
6GqVQBT52YwXU/b6n2nVfVjeBcAxl3r581wfbzIMaz3al7VQldsGqbZVHGIBlvcvaq+XojeJnD/S
xd3wTGHWFDfVzowlS0n3VHrfB8HRQCt6s8bngP81meVX41CW+2qj1hjVoal7z4zZsyiWPczGIMr1
YNhWxTW/sH3lWopO8gqmkne16PT8pAqfXhwrvkr8BtJ2ush7ou9iRYjJJ/H5VLjeQe4qIFN2cT/6
zxsm25qnbPUV0sYwkh3lN1sB4JfljyvIvV3dc1U/Wct83OUN8fz1dktVeI3wn+1jRxS+8ZTb25S0
JU08F7Qd4d4D5zCqaHfQ3zRq+mqkMWrvWmI3etLwk7PDYe/xI+Q0UwKoz6uOcj63ACAABGVb3xQW
r5uDH2TNh/8T1ZuT8bTu5klQyrWXHadX2+qJBQAL4u7ZSQ74Uedk/XfkpF4e7/RWqNzo2zk5CrDD
jgH1u2Rg2n3Y+falQ07s3vdwUPq2fOy+KMC2vs5xc/6tMJstqedEIz0Wjj0+qq4TduIfaEAUAiVH
F0nVEgdw5CDxncmqsTx8FhQfQra5KMVy739MqTZKyo0x8F+iR24rztCNBULy32q3XtGx7Wl8vNnq
1Wl1DM8TwXCQ1LJuBplpMrmH/hAws2CY6nW7HD7gx7O05SZ80uM+HVSkwieIoEs9JB8W8O7zVdgd
hYP8qgdWnzGlV0JuPtVqYa+QBJQjWLFgQSvEstyb0zwsuA2zCaPnAcMqQLy+uaEtfkzldbE51JNn
hDYTMnLktSiaHMD/nPbi7s6+veKb/lq39MJCBTnZ2lr88WLvCyWUeVSrA2P8yov6qcbDBXtpMVEL
sgTIR/YIQd4TtSONGKM9mYoA5TjHdKAAUBOuK9W+wsTLEUCf6cgswvQvLZy9tidv/v5baLKcalbj
sk6IArQog33QzeR28TcJAq7RJpdOSOpREjyloQJU6Lh2+k61QLst6a8ZHTSDAzduKkVQoNth2ehd
a9LRK2+5vM1puOEsYk6xl6zBw7NIyTHuzJ55hZDNs0QGuWEPGlOr1Re6eN7Kno0UpGf2SX7+Lk9F
HWxx4cafKx1DreZMC8P43ttWGd9MNspvP9S3mOJBLFdGHtTkOXVK2+IWBxyl+TUmsvocqP9oVoVZ
0/jKcOiHk3QDNBl17twfG/0daGmhASPtcidDzhiPMftJIdgIp8jxBtogwO/E5hHWuiu8ixih7vSK
DJebNUigsGRcc9l/5944s7pNCAznRhfnOPXQ4rIeHi7Rh7Z7w5JR/IswCfxUenKhVCgESCEmwUMJ
QCnM3r9RqOjvVINITq2+AmwNU7w6QllR09cErx4lyaPxahNZKUZzapcmDBl68ZC2lVIF1pDBiO1N
RFcfQ+ifj7SQnkqeKYu1fY7FhITLlw7XYGkzORYuigo8fIyy/lo2UHFSsg5eZXbTvO8wYdFg6rmk
3nXdgfqs1qpDMEIi8oLip+Zo9QeDe0tPpcnl6vkLLBEgtd3I9vzo0BVDDF+fDXOi1oGkkkAjemka
H1THjNcKPDtizCT05LZ3nejnmyXYFvC1VJcq12+bJFLbzuC7L/Wlze4mct3lkbqd+y3DyxSxRFHy
/IYXkwa3x/nn1SNwA/6jUd9St/qU66xDSpynOvokCVOLXuUICkYcxxZS8ahIv5VGglL/LJROX+ck
+abkkIXCYJGFNWp/bK3+6m6Go9M/INRqmByApX2ouUZSCClafabF+xOzDDp0A0paQYZVKe0iDsh4
DmwTF6RFSCY9isKdODklSdvGpTRz2OpkS1nhbIKjEx+X1HwhPSz0yiSdRt/r42dnxxqVZ/vHN62u
5Cg82Oj1eTq9zCbJhGWL2tgTfLavByRp1h7cxzYvVOGPCh389DyKPXBiUCarmZtpRxRHbCXXsAe6
KZ3tTU9qLeNjV2XUJMAP+LqEAjbPJG6yZr4t3RCu9llE062hXc8LfCjEQ8NcCCLHT3JUEhiPI4Jm
Tv4maldDoJSIrx6cAZCs92tHyPO6FK2fNRvCIm9W/i3nB8Zc1yF/O/nNagj7/xRb+/+RVxyco971
aubQYPz0QwQccm5Z0pyjQmQZcQUeMjPNNHqpEGeLP+DT5ib6Ta4VX8/KZRcg53i1o1tv/xr2cBp2
jDxyPxbGFU2rkYIzeC9bBXo1UbwRQr2x24Rj2u5ID+7EuQjnPFqji2OvClz7VfJ6tetcHrtYGO1E
PeHelqAGzEa4E95ad4dk67s6OLF9MR9pMm03DY0RDJEbpNYCGWl4xZevgKurhQDb2Aaz/eS1ETys
WRVpQLB/V3MpVThn2mlIunNY3xRnvdz6ZY3kn0ATc6LHHf0ELOq4pCG+vM3MfiE0of4qAfheqT1h
5kwwwcMVyidtWGiEa9JsRFWcx7V9W4SCmYPaZZxi4rpbiKhnOvGwqc5AI1rriXLMttuDNdtqTKOc
atKkiEx6WbXOzstr+X5FQb8mKJNvHFh9M/9mGCsd2DLIqSMX+uSzzVabpnQGuaquOVPJtYvoURib
diDOB8sO7HUbn+rRC9zqrQAmdx27xHdPzZe6E6HnCPK4U24z4wRo5IJpsEiLjzOWr1ryREJC5pdp
4wNr7fyIHTp4Z1Oh5U6CrCK2nPyy47e1liwEw2Mo9w7XBeUwgN8yPWmy3bmx5XV0MmlOUPBU0kPf
2yrMQ0f9AKENeKYqX8d0/Sf4veCtLdlCu1PQUhlJ7aFr3vD9pZ6TO5SMZu0vBPc364Z9e8zWIf/J
bcd/LdSQ5IUlEDG+1KBjP0g70pyKa5UJEwokW+kXg4NwDKy7kbCbQmbD5+k6rYJeQ0WPM+d3yPvz
rEY0pEXYQ2SiEw0n7Tng5BsS+le9jUHSn/wbM5n139Lrnn+yHGtERqqyzHmO5RGZZL1oc3RtTR60
LORzZ+TKoJZuZYv94W6OI0xmjvkF8kr4464ZsY/Q0DR043utBXTonedsAwIaTJBkwUvuEF42t5DF
PmUu4y/sw1H4gdf85yub0IGtSZW7gP0+MJXjnDJ0h7bKGLsh8bOA/2GjBLORlWUtN4t9VxDWSJHF
BUaIEhWFnSL8fRw6OXLtaPScR2r3R5C4/gt58oaXfNqpC1yVdyJ8zjFWOG6hk2FAyiWvAvdWHKje
b7ZEIBl5+DSUW4D5yvKFiFTj25CpHM+8UuZ5VX2aYCClnOYS4L426+le9lysbCu2MdSyrQb6IhkM
N6eaxyr9+4TJ4MkWRExCdoo0I4d2EEhELkeQ4GRwZoowVhLFOxbpNfKVLtwpGqffvXtTk4LYdBEQ
EhnwiKjet049xkcw0xQ5gXvIBZb+T+oPO3+ZImzk+YXDQUHCX7Q4mHHcBqwzTAnNiRocvlVHA/C9
FaJoOECTFEoXSnCRG9ZfaufJ7qVWaImbme+1RevKAJ0xqjhqSt0kvr/eyxd/IPOGpGpCXByo2CL9
J0UW12CTOyQxP1RDnUxyfRxK70rT7kKF4kdH1X5fI9ixjTqxi2QeTrPKQNy9NWVqCnSgeG1xb9jy
xYsNIYQNPG+sZqfPnLXQZR8Dkw9QgKamZHAZEIajGkD3xIu6w5xnPcj5CWy1OroZXZFvyArS5eor
NDRAumoOSy99rwlk6hWt42GksY7+Ks8Nhh5ufxX7AFpL6rnEhPqDL7FzhVWHT1EAlep9AuL/bAY5
bUsaHh3xURx5mSjP+pe72hKi1aEObxXM38ypzjwj6QzeCRAu36wL+oE0w24W2zdF/0ZWrwCJCk7l
XBp4WeOvpg==
`pragma protect end_protected
