// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:56 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
fVmbDcGNn//Ydcyzsl+grWqgwVZiIk/bLopD8/cnYTyZZ6v2FLhg/ufRMWMeQvSh
Be4Iqi5Lf4alXdRXQoFEnL4QAB9lzKq3s2xpe05zc06Dbu7Uk0v+EUtBjqEWpp5b
R7+hCJND/T9xdFzdJp0OAQTjgaTjPQFIiBaPNFhHn04=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5248)
cSm2YZhiZ2DLy0DkxAcQm0y3wpKdfovU/HIH5NAMZVyiyz6EaZscdQ5RmhSMJMJc
e2az2wVPtGgWXCaJ8g4ZhQsCCGhRT6nwgiHxuRi7IgKQ0Wskh+NK7HKRnmXobgyK
li0ac3wONLHrZcqJ/5kyFIuG4agxFLUUvCkB3rFE69y4BRZlAzaLeHmN0ZHxHMYj
ssOjc54t1A+qyG2lmS8Fhkp2fNE4Dn6rzUMoFVI9Y3Jys5DnuqqDBH4RXxRiFyWs
3GvpUvGVrwhw9I1leOSw65UJDF2vP5xDqO9YsHPvUvDHuU0LvWzPKYOKBLLTgu3S
RnAtJKRWVldEt3hOxTvLECSyUyKw3sseTcUOsHm5HFED8c+4dni5rWdV22QmUfZq
KIWpX8cLBCfJ4HraUdePw83yEMaucL9kEun/tY6V097C0X/AcJsNFvDmgnGFJGn8
DErsmukdrSCAt7KoYDhx2ZXoQdM8GeSUbYy39mGNo02JQ6YUvRCH79CNQ/XOLtvV
sbfOKWVNvgHBAF0Xrz6ZXp6Ae/W2IOi+teGg2890KvIA/iOezZKs3SjEdr/N2AbK
gL4u1dNKVkIx2mFqGZMhyrfB6CesWz4VP9VEU0INti+dDPukVrF7G0i8/DjstVXv
o2NW5Qad2TZuvTg31bxolUDg4k0KV8VbnAT+gURkp0ttX4DFp2pQcS2NiH1PdlpE
+TJaLPOuFyxzcG3VfkdrVwGJ0Hj9ksBVLZSMtOOa/5KxnydrQYTQQ6HESRQ4VzmP
JiiienKfBLihvV0v7TZQAGUBhQkeFh0wTwA0UN9mbtyr2uXf1qiydDH94X1QXHy8
Y2nbboTPiua9xWPM+sfpHgj1cHuX6BQliK7eip7TZ+hXkM5N8W5bXkmZE/91cebn
ld4h2saMPNTIUUBTOj72rwgRdaOKSE49qZjS2F2VuHs2Hn/wGhA2mRV1wgIyvOpy
33dD3tzzxZb+M1FEuLMeoGenyV7tx07muNvyZOLLqK0CxjwVNvcoT4O/k30mKo8W
Up6goSQGwfekny14U7MF58lHb4tMk8M4bOkFimP7mqvHNTOVETNk6X03ykVlD4UG
SwmQh0eevGBws8f3+OH2GYMj8iamDSANisUN3PfWvugdBfi5+b2gDqIm75iCdeGJ
5GXItJzUsU0qrNMhARLTatRbWr6wqR+cc6I3q34RF3N8gfyH9RDR4/+iMo2xRhNP
DXpFnmAbfkqmeapF4oEH7krbXhczqAg8fnY61/qi8cYrwBDVgbiXWulhR9FebVkv
nlFijpEF2nJ4TwS2PgvcdQal8KFVYo/MBi66yM34M+i822t2OnLD4wJXACSMY+IX
I6n6xrygAloitkqenK7mm1UCyVNhvNcYcpqGMHYPJjuJfZS/+YyfOnOyPa4cTAW8
GH2eQUA6WpcxNH5hLVsdumMI8wkfLHUT1hxB/i9YNwv1l4VD5oVBhjB80WonfxUe
KDW4z4QP8TGrwaC9Qh01Qp7eUevVPFyru6j4zvKhiz0sgVHVi32djxdSOltVFHLU
x3ngZMCurf7Ie82OVltCJxf8rfkuUePnRi64DAymp8dOZH+ND79u9zpB++4PyRLD
wWOfPIE7w14WKbhoRLY8osxcz8/naQFBRE1KC19tx9bNHcVXWXqwx2mAsmnEiOtA
XqfD7/8/VkAVwnVRzDSykxUocRf+AI0Uu+0J04I+zc8J3tFzjjT5k5K7In9EKKcg
lCl4HyiUPAYNbxScJCGdeR8m8Lt5oAfYx7nu13CMrgPUxTrEECKGF2YutXfkr166
10gBUQrLY0rfDZs/d31fKvoh6uuR43/tMYrHmU4jdTfEA5D3slQj9NrHZP42SjA4
fmuaIdab6L4ZMrGrlDUIpSHiACA110hjA99jiO+q7HYG01MiN9NfBMExvq6/+BsV
Jr8GWRZkI6qkWaRLwQQKuL1W5EVQdGAyUQxj1Wbx7ILiVw4eIo9/JkCsoAxmBku4
jjRBvHwVJ86dnyc1GXj7Fstivdv49slik8Iisu7lX+4Tt2X7+0TCoSaMSXjuxgw7
vHSuHbkMvrBBVuL600xuxDpzJd67QdnZeKDUhwvPwspKlyx3DY/9VdebZPjxVsQ7
U1FBH1SC2noF3JDJPFFqUG+1KP1VWzkjL526StV62NJgu4RdmMNjp6NdposkDwIN
5IeHXkdamTLI5IHMnwl95riTsVu4AprfVe+rLn8w1d1P0VAqOWy/zVXTxVJChtW9
zhmNYpn/Bz9rZcKNCo4HjL1Hp+QeWQnW3MorblIbHnItbagMddFVTlNj7oWJMIM/
dDlRX50Monw+nRtVAzMlrMpt6r5oRS8P6T/MwuA8rAqI5tYPJiXzTtnHL2nTIvl+
VkJB8J9727g54Lo9VDOkif+4aPnWX+KAgPXR+Mi9SC0wKBh8oHD0UPUem6fdSSBM
Oi3Y1d+d6nhSjXVuASt9V0mM9Bu6LY6LYsLmaDtSEcem9p2mbWFysj7CbNJoRIeb
Av1Tm/wugqUAG147CswnHL289/sZs85lc/XHVcsb7v5cXAuqY0bOPex1eZ6NNO7k
eqL4A4Cv0AF7O3yYzV6Bsyd3L/IwschTClOcYhKTV5dJK9Q/+dkdlPe386T9UHWb
tsDsXWaBLQayWGt1qj5dZIZ2SrxG6fD+eeN/Bynvx6ubKFbwvVRWObugJEx+sFe6
aU+XQZe8YY/99EOtRG5iA7cxk5qhpf31XvJbEXpSAXH1QYcBkb77SZB3KUUsJC9J
kcR3Fnn31TooQgUlThYcOLFdSzkYq1+BkouCr1IhbFqUeKqNKrGp8sfE5q/wAAbY
herDmiuuiDYF9LB+G5u2ezlybkA5W6ctq4ysO8lVE/upD9F6MO1LmEGI8B5RkmIK
KnWRO5OqZuihwJPcl80kaCDQJMpFh2r9bbUe+dQEE1jMIiHgWmLrQEShoYw/Tctp
sNqw+XBz/M7b7K+OBun//awRtR0VNmIS1wU/pMlCzrf4QHKKSC6z50DRfshDBLZZ
5G44Ut0+Xe52lees2mRGtjaN30cM5UNDTVcUjrH/xWdv3G+ncU1AuvS2/iyz8l3K
mle02H+8JFeNW8oNCSwqn9sNJsPKKgb7PlycFS6jn7y6UioM7BJURSHu+Hgw0Xy1
V9NTIRRz9QJ94gmnv1Y2zt4LmY68g1BXO+0Ky9xrdXAREP8RqlxYg8Tc82093GnR
aElKF1iRNfCSipX9vL4vObjmiMPti5zcjh8VjRuI2bTtOa/t3vZu99dzcvrkWlQs
d8F3+akSM12dCd8Ek6ChPSLtSeq8f3nhCHlMxuw0Kj3Xie7nXjtlxWQOEjq2klaS
p8PSM28AW6GG7UQADn06zAg79znnmTu9414vxeM3tJNKsAzwt1NaqXJ2kgAgEipW
z06EBO6kE/ro4HEKgmnz5mZwYmEy7CbCD60G4kle65DRvOecsokc+v2UcEfiXGtY
m9XnICoVmoufremxp8KwuHL+MZWQ+vsggF9EqyrVD0FqjS9udP80WW9W+ULqtoCn
QdH9wzqnGhRwQDQxaUibj2XB19artB1lvROtyhE8a6L5nuTngG6hWksC5neSfBtq
F7lqTCgOPj5paBEUBEnMfWRbzbvq4f4GnBux2VPKPYrjchP3mBk8tuDvc+xhidSB
WyyhQ8wo4WJ0Xc+7vUdndZgHVc/wBKueAKSAnlVjAO4KfBBQl/5kqkYG1ILyksiw
d+lJ+7LDRyO5CSbbdANr5K3uezXcjz+J/r7m0wXUFRIA4wr8YZnU9Ui/LvUjs42D
RurvzzaBENBsXUH5sUsU+Win7JHYfF0Y/WGtyEHAGwRqoyhPw3HhGs41XNnAmTAG
JgibDRq/3mGvKw8UqAYD2Wg1PFvg+A0nkJy80LAM4r9Qx3jNk2VNJ4JW0pQFuNtC
EWqIEx0kt8c6RxyhqFW7LZV1mXvOEzPShPiPgh82mghAttxKP35T03Wtt8ebuxez
JvI7FG7FAeiHjDJm5fF0+DsLbZXYn3tuxqP8E6Em8HshsKk5XMOm9xBmDP5rXYr8
Bdnm0bmgAdxebazCbfviuyKmNQpcm3/D1kVV5UHJukl6VWfEVMNSxiCEO8mYmj+k
96N6BKsSYyndLw52RY0OXxkGyDVUz8+GVf5R9Y72hVh0h9Uu7ihxNzjlJZaQh4pa
dFOc/4/2WzD3eOEQhpkDeZwE56eNpjL2Q2qFL86gDOOWQ31ACGlSRDZMEJRdzZ+q
oUcimbXLfm1uDN8QsoQdGEa77cIAhURJzyflxo0cP5Hx4P7xbVu5JDhQ/WLtSHkg
zIg+ky1mT9TvSPd0CZ+TUp3eHkWDZKcKmAa/Os9JUUg3NY7NbPei21akBj6u7Exw
M4qjyqSEOtL2L3aosGFesZtXyaAqUnCw9wy9CM0oOWQXO38wf3HGOvypt+Tr8Pc9
EGvxNNOnFlsxNsitWC/2kht3QRz3+Wc6ov2786hEYE3p0VY1fpys4QMVJsc6bx9s
VDCM/mo5Nhq6QLkWLjf6pwXfN87b0/cD3KZlFDQHMBEObMMdAH14sbE4pp9M85W2
rhs7Ax3QC6INicsHVVXRS6C7P5teY9IrmGclm7YBJvbm4q8Bazndp5VMIs6e3nR9
QWNJglSGuYAW+Ol7QM2gnw641NtgTXPxPFM+mqjXXa9OXMgAClXH3yb8HFE0WfeK
eYnFT7L/vL1+EIkkXqA17ROxQfHDGIme7QKirAhGwoj5aj7OVBMQAu8FxuXp8cBa
xN4OUCg/o66+lvodx9k050pCSoLsZZ3KuA/bg7ow30CR33v6Goza/CwmdhZXkd7D
Ic6ugNTEHIIG2nK39eBfFU/j72htVM6mkC/cwZn8UVJhqvX6usAaVqTKvrzPq6qR
mtyNyuztlZGB9Ph4vZoK4MTn79LsHvJQrNtB+3UL52/n9MxF/ZUqeNQC37YMXJJs
3mKawOXvv/LqFtLM/wR5XI+mHF7dFNQO3Q/hCoZab9Rz2iLmSw9HBRKNFlDDJXN1
pNi6NlEgNZs7cz5kTc3XC6AOZrVJQgrNCPhqmdTooqCnw7nrZe2grw8wJipujqz/
UAsHKz1+bECk0WxJhCELiNiN8z26El1v7bwIKkOT0yA/zplLYhU5ljOGr4aB78Vq
ZLNY6bCeuLamGYHuU3FF+O4/qLboAY4tOjmOatlTbF4H/dMNv1wAjb1Y6fCrvTyV
b2Ndwk6UHNQUhHLSPiRHO0sxt9dBZYvSLPp/jIcbOaYMu2Pw3MkJgcRk6sYGGeGu
1bIcyqAyN0KQ3cX7ftfk6sQRWPonfR9roaM3RMUVtxnO2AjNrGpHPlBmsJO/goQ2
PwJlNEae1MlDm5D4kt3z1pmRtMCVv9PEMckYICusqofGIpeHjF4vdnwbUDUK6tOH
vJzZ4OZBThtTElEea9pg2m0AV6irGKFI6pBSSy4fCkwQZvrt+wRdsvb0+1ML9tEA
hTdy1NLJvTAEas2lIDQ9CW550vHPP6sMH4ieItdFydTXMOyF3OCjpt2AZcIsfYMb
IajLSa3EK5eGbaW0y7BuIAS1Rp3DiDRd+iXMMGOPjKD21fVsmwxUFnGXPk9NqOzA
zBvRt3pdqWBhMrWFluUjKDTubj2ecfg+T/YX1gLyKl/hxDpvkPwuY0K4sgQojhPr
eItnEG3HhG0z0cXscRS4Gb4eWBrMD4uYPC25BI8TZMITp9hO4TKG4vy4TiEEIXIj
lt9cWI6ZbdZ8da5GW9DeFE1Fy/Lbsq//5GfCNbUE7hc1Ua+ESjyxxifhaGQ8VyP/
JsYXprvulo+9tVwkDQO0etxtvR9VcVO9ZDCsFYHb0eshwR63hNMs570/iJQbHlG0
83t7ECjHuXj87Hw7WeJs4kORSgBnEvj3BcabrTAorwNEgw1ZpuzZg0PWUdLKi/4V
z2nEq1+5rCGOFjJ07audB2bCHc0KFahLwWdkWMhnZSU3mgF0zfCG0TBqcbW+YFVj
nJUuhW+Gy/4OOxLbvgcENLacuapiGTJCcz3m4JT3TyaKdK/3vlecer3MlYN/iWeZ
UzbKEDNszlZkrDude/elLmty+0sSkb1Jys4vTPS3JqDG2DInJx0i4EfLcOnCTlru
0Jg2SZ4Sz2jo0XrlxAYgJ/yPsLroHFcip0fz1xjiBVKku4lhflIV5naeDUvQy8B2
apdVDPgQaEwNBfUk0tnFkTXCjEjE1XTPwY79ojdupNQFGcdkLG5engQQpOJ+pL7y
T6s4lM914Ap9BLANi7Mn7kmq1tJtQrgO4nvA/hjXp1bUwAApLv8Q2VXxnVnhsryY
0v0HsEqCUWDmkxvFqGuA+iSnHWJSrxiwkIVJD3+SxTvz1CPmeICS0wksNV43oDii
uNgF6/i7urLYALhc/1zG2dIAGknFd5fK91qtRvAzCPibgcN6JA7VyGS51eWYtSTS
9uyKlMPqQy/cUk7pthZujgf+R0qjo/v7aCbGoBluB827NGYNQX+1b2iwNRr4NPhB
a2NuYU9QW3R4uQNBZ9dDJ3ZANBXW3AdoqltTui3PPvJPPDyBtBUlod9/aRggnnMh
r3kLk6FNAkoqMIeOzm9+IwSE9XLomhdRe5c8f+vF5XXMtq4FWzOTmPN8zvNzzFZr
ZbjCGBCMSA9xnxNB+UXjByFE27WR/nOR1z2jq/TNMIC5tv6lV/8nA7gOVFtY/SOj
hcpcwQhm144lfC7n2FunuFwLGHLQsaQNGb7Mjh+Chg8F5QPwePiaLOMOQ0a9HMMk
vTM3MSXIgc9NKF0Iuz1fvQ9fH/KYrA9ZmB5E9UdSHUVrBt+HEoII+5truqQv7Y6N
UAJaXy92FuqioNVcRepZrLzL+XJcT+p7cW3PyPn2CtCPFRpn4eGtx5Vwl1gO9Clx
WXNnDI+jjVyOaFpdAgBe4/IIRfw+SlEsZ++dGweJEhJMKDhdeea1yWIIzSO7z3Mu
39wb1mCuONr9MkBP6Xf1BciI0eDTx90PYmOXyj42zAChrouFDe/q3DwTZlcA2Krz
KKicfAxWpHgrWs1NyHthkw==
`pragma protect end_protected
