// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:37 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
IsHl/1FLhoRi8ipLaPsYak1hFMA9jwdLDUAKWHRkjy9dYAr2vDvHb6DK2LFPgIKm
6/qSPLufCrhg83bQnRUlz78QF2GREPRO5m0YC3ebevV090CDpkImwWi1qh816li5
+7zFQffPIoK+FVg/ph63a4f+ofdEdQdyWCqH/Vd08mU=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 10400)
p2y7EzuwDNBu6E0OcjV+5kJM2dh3JWz1AnSPJBgIwgBWzPDAfpq8A7ESMIRJb7jw
+FFxiylIfbUDGucKJfKy/5Gpux5BK/v95JQuHPXMxDun+qRBfa3QFBZM8319urrC
KF1k1yS3D/T5p/NrOIlEvWHxgAmvCeBs/HQL1zSIkjreQMZt8G6xPiItDOdmFy5g
SBKD8R3min0dlZqXiE1sJnHlxAALEYL3z5MusJf7MGDiKRk0rYgKe3GafLt+pTPi
4GYdEwjqEbzrrt6W0Va5z96qeiqEPH4b8vxiDEliNN80uRJEUiykdkKHGb7NKcy1
NBKGDa9h4a/9niIVAVVkFsJZCv/WiP2MDVAZ8uf2ZG7jXmnvyrarUX5n6M/YMhEt
WBTE7ZaYOqpi1Jz9aanF2bnRsVORVKdg7NqG/xDeGCCcMRVTXK6rNqgxvktKp/tS
0hrAV+Tnnt2JViETZNjqaR4BLObcT6g0CmDlaHs+TOeK2ULDu75583qK7HYnlj0i
rEcCiIpotXuRIoFoPs4MRqCWmlftp8j+7vZHsTgKUgF7ZDrePicaweOCzRimevm0
+PXe2Zx+zUuOnEsLb5yxS0Gfcp5kRKpZ8VKXNgGt7OOMGroACHRvYGq5ju/0Uc++
7bWzYibzzmLwOoeicIwsfKi/Fd3U+wtFpBvEwo0tkmLeKXfFOz6c3wGmNekqDCQG
qNGnMGn5reUOCj/LMUdf5dyUs6XKRyJoUOiKfmcErdwWVBX/S7FWT4szsQIqGFv5
FL+Ffs7o2NjUadggmQvYSleV3TmLH8ky9L1pY/CIwU/B+tiyLqRgEdr4kvsDBRLz
p3sIH8zOHd50v/nX4Jb/DQaetZYN/QMpMk2gmYUgyEdQAqrypTKPyqFQgxRdh5W/
05EKmOg7+gRufi1VIB7MskCy8pajfVSDCxQmOG+OlpJ6wif5ySbMNUVm2Uw4CsNG
iITmV7jOOBwPWtRTIQkkWARLhIF5j5M8O5BZ4lxYO6L/9LGJeM73nSjV/MfIkfyQ
xkG+VbnGFws5A5ide7VsBOqetLoqpP2G1XfKDovH2hGadkJNrKm2qPfWjyfON9wq
GIXg7K+z8aQr73NlVYrsnnRLPbVquZD/bbIPI44zDszUfe8zhpPEHeZxC7iSjqOp
1Xh4yDbGn5e+UbjM81M1GAlnjatTPqIPxX4c9e4buU8WJMg/7KHvSgPnrJezGGtG
wy1OwbMFQFqZSqR8iBTTlRtX/lBMvuAOhcN4oVjTjVcugXONyVy3HiKVRCdZDUPn
3pyFit4NxtO2k2jXVTAsBq2HLM2jtgZ8rJtX2vfe4VH9ukMrl+1tdsfhYeycKIaj
euWcIUK2NGJsi6ITUgA9NxSWnTqHcVQxw+Uu30EX6ENipCnD+0yC3gfOBlXY31oj
XJMspgXUKBepmeQQzHqHqNkI0jDO7I+MFed1KDxFeo53YXTtwS6WJWmKE4T4S70Y
imaE97NORbNDh+3mlnD2uhCOppfLo5Ak2fpQrKdkow/z+FbTw36E3oJiMjf7CidP
4vcTZyT14WigHyOLSgFCzFDke6/lKbMnAYk+ROegl4fxOwpdqkvWMYkyIq1K0XQh
kYEWS4iLk9AiF5+0UlPeEvKuJrhe5bDmGDtqtbQLmc2jWBe77lsDRC1r1c+qmVsa
Kq+Y0wE+6po62cZdRMJaiYb4HWKiV9cb6XKScsu7vi3t8Fi9JVHtuVl+Sn7d4Irr
GOzirb7CqIVUf9C+dk2DzvzpLzlVscbKUzczVpI4Qkie9XUmsKxHexAAW8QRMCjh
nYMDCieSG8fqSg+Lf62pJ/NSkZ0xa6YDPLpdyJqj4RIOKYRTmIskR+ZjoeqqFgLb
xqVMD3GgWn4M0vegC0f0tEQp6afRs2eEL9BDZr7brp3zE1NSpwoifIWGPt++fKhG
lZXMaxtgqBtSQ6n+l0lQmRr+WJtt9fDJvnwJ2W6j7b5LBGBElIjlkFhzC+XMdgGn
1ow3yqPBYUqD8R582sHqtUDiwQCOqjQcSbO3DN8LiQwaBPX3Y21i7f1dtYo+ZUel
FQtkogGpdZYS43JByf/yYMb52Rhk4f24vR3969Dcg961XizSSMKhfVkaziZYPCkm
HUMhma0r4yFImLhlIzokRKA838VXV3sKE1ZypSFP7kWh8TsLvgNjypbdMAMQlVEk
3SY+iK/pyLztic3VnMnSjVDSGNJeZtMQdi/P0BpIa086l5Vh9aRF07xlc5nsfhkJ
sQ3WSpQT0Z3eAOYXVzMxLfDWv+Hy3lUdW/HP/k8fNpiF1H3FWGNFcHLxUWXibxJc
LPgq6/yA4Ll8X06LrZcgdXv1DU0u/dd4QahjT3+53rgm950tN7Y8LITHqsy0Wolv
GsQ9vfviZhoPP0YWmTDCgLpOjDl2zdZGYtZq7hycwQ5q0P7SNtEKTAHDmYSLuyiv
mPFKbj4H/GdrTyLNopy2Zi4AUhEbQPdMK2gTe0UtlkPwOB0QcOyiIp0g4V4FzI0c
SOSpbDYFxTqGBET83aKenlC0it7dEE7OJnJY5/zHG2wldfV6RjPc4KwCz3L4GOCn
tFivZCAFXgGhGP/4uvGpTwPzd26lwhtiHTjXaWm0jzz4/PG8xSZSLuf34dfRGdge
2lSL+oKbZM3cEJ+Dt+BaXpZchT99P8lNdn9bYobSal+V2NfMU0lPL9tGg6Ig+yp3
NK1YlEJAbir0kJN3W5qXszbL6fAfC0qqvgpcHDdTOMrC1cTg8nppO1qyafC9ycWt
+0N9iWVGsHWlJj+HbQl1aZ7+YdKA9b1+PDwsNtBOGS6Ty4/UKCrslck5194KHFVv
nvF07GtsX7zplPirRjW/w3d5fHYyl8q593W1qzUeUg+EE8wDuyOhBDjDeIJ3XkBO
723ConRPTEzgjAuET4m7pMox2XNqO9ENn8eEYd3b1ed5+hwzQKZ4UJSh6pYEaw0P
i9i9f0CYzapCG8teviDThZFCgRwlPB65jYPCfdldWfUa7gFD1l1CkqJKmD+wBeKY
/fOe19f7aAWdW5ynCM4eEZEdtzLRP84hLv3Rhnk6KZouvtrRYp2bBfOmx0vBGzjH
KiLyiEnPbiwJ2jxoT+/96nv3UYLu0oRzXj0jz2YOOr5k7nG156gkFVfMY72bHw2f
FFgTnZFQSQ+kFapyPwnacLeJtLRnfnqdcokw5KIcvJNOZpIRLiLNDkSNIPPHGH0+
HpgL6cS7lOfKFOcx2KiNJhbJ6OSCRaneW3DTQKyllwvNIBdLozUGq7vlcmWf7LYA
GZniOCC3ljVAnYj7PI5/jKuXwL1jDa8AKjBRiMIr1orzDcceS0TSJi9axYHSvZID
C82QEBn4U+jFVmVmuoezuInVNwyvmv/6KVcL4ggiu4n05pmbHVwP4bmrDtp0Fcl4
11HxOVsQIyJa9M+VV+rBje9/RJD7sz8Nt9aHICaV3ICWTjaZ+Wz0gIDAdL2jxxN4
m4OVFCXixWrmgGxHb4gxgBjohaKc8vjsdML9q8+UOWvwARisP7XtL9wgjDbTWgd1
HJmV6iDl+IYVrsJI2iTHHWkQXwezFmHE23l2divS6t0YGzYy6jKgKaxIKA604xix
yOtt8EqLDJRIvJZ3eWeG+iqQQSX5sPAtsqpjgA596+OWgKVvlyLnHuRmYTph4e9u
lhsrBVy6PakedZKiEXOv7u2qRIbbNk8vyLenW+0NQiYGiFkrQ0BT1J/oycHyH+Ir
7oOEuyjQ9bH6jkX2GgVpgTaApGnT0DqjYuyx26IQGp88dvmC36NVCv6osaFpF43d
qdRNLk0wSRwa4gjNDj7gtXq/YlzvsHvUXq0P0+XYMNqst2xpdZc4VzKQRK2wyJ1r
ptdtkD+ZWeotwPCS3PUtwauexG0UB0MaKbo3zeajPN77+zczofhYDIt5UuxUc0JO
dqvhgaYWqxy3ZmC3fIZqEAkbE0YtojqQ2NEjFbsk/8cxqIsn/kGYi4RYSNL2gZ87
fudpo9WCHQSVmgFOzSANAZxKRmpG+1/F53dDTozeTBTrsyQHFZ5lM9zc5jVH6hHU
1lTrSP74o88lPns0uWvmbPk3kaMIeSB4QKsCFIWJLiAGXDat0SMAgBEnJetpDdqZ
MU4bppGy8W0/E2ksQ0l4hSgetSdLmsq7EWSqRQyW038QwAOpGdMhYRuMFBLFjYX2
cDbwPgm8HoFQMIIo4U2AaDrsnLYHc1CbBfAbLdvBfGGMYPVBIy+GcdV5f+7KNRf0
v89oS/m06PlkcYsVqDhTrfbPe7bQtzC5chWGxcGR4V+tTAtGN6z+a/cs18cahl8D
waG/wmuGWsjRHwv+Gb9S9kOXa4GSTA9ofa0MHsNSa+TibZnykY3mt1H6zLiU6kTj
GBhwW1ANntB2Z2sVSrEnk0bsY/UHvikPEjnzdsq8lDFGM84XB3UpYRe51VIZksoW
+0WUw3Lo+aBJhoRoKK2ak5pwwDGil+oVwwMSiqVctQ0+QJnuzX46r/IZwMLrytMh
NKj7E/x8xcTMPnHcPNNrlpaX8GfLcmIewgbNgNOuCodqeXwH+3oAE+gsPDmbt4hJ
0n1mpe+BfIT4vkfUfniEnZ8ltC7SNaSOFvcFJf5FmcoOUZe7OFU4gAcTiNia+mXc
GbHn8VU7MqqNL6fbv2aZXNBJdQCz4kD6UYkt1cGyiPRWabHSv1T56QlzPXle3nCO
trs2y8fw2YxcQhBMYYDqJQooRQTULUTfCXdZUhLoJRZJRUJbHSReswFKBIgTkccn
FhEkQpXUu4CyS69zTgfn1eUQkrPl82gnPa8j/81A0wc9/Z5SV4o7IIvNTnXsczPW
3qsE9opUAISYtKlYk9Pk5NgAHs4diI2juBbrZk2NE4wXcdHL0IDlZmBFQBk4M1l5
iqp2C9XwXj0ZKIZ8zL+/u3bZBqR/l6e2zU5lowtgl9L2o1izjOqwnwUi5MB1ssyM
vDN8gbBHPr+qo1gMgXMfK/2Gbf+HJpPWvb5YgUoHE+2GdaCltL6HOlRy4Zoy0dGw
vwmnvCt4qredxjUPxTviYKN9UcjCUGANmGO+hYxltjOF549SkJ3kwvcMfJfOaDpQ
FnldGLniQBjzdqj8BnAzMsa7Fl8zke0LSgQROkcDhlmA6y08iybXOaZOpa8l1IN7
oFOJuTc9McWv2Gdb3Q3ZGOWMiOsB0DLDAQC6z+kQ5S5soADhxH0fpn1PplYcKJm0
y9OD2H1HIH8wEJN/WceLW9aQOUuaAaymsleIXtVgC3orJBekqLfJge8VObxU8yj5
lmj4CC/BYBrgRGSbga+rvP9XIsWgbiPU09GJ6lRvfqQuSJsY5vkAtLZEEf9tBJYg
0s1tFqC34FWlc23TqKEBbseewhDPfN9+zSvhlwNG0JYzm9BwAYK4NA09P3gS/Xt9
pNk1fDQ3J2g/sRvU+PzgEhrvBj0aDIShvimbSzvv7pELZFsDt1yUOBtkoFxJIn1s
iYKIvIV14w1V5zvgUX+AVJQCq6R/4ooeyrKB/SIySn3wCZS5bWKFl6E5myaWoQIo
/wkt+ZcIWrBVMRYcABEA5LK6gCdY8bxGg+bgjnfwoEw7wE579SWARza3JqXf4n2Q
fZKd2eDRG7rO4xHxWwoR1xMYZEqL7e52YX/Y0HsV8eu0/pc2ZW3qEp0GR+HIOeCG
foVvJTEm33pU0aiYbz2m0CTvcQFVuj/BpdOfzg/D06ZKSkb622COqT9iKugnWE5V
PH1w/RwHOubCm8SiVM1v307oyZ2ZXQLWXFerJ/HOuKN3Y8BQYK1+xUJS2MhGa4dO
gVBnbABfK5wPdUlSMHNekkgrz2qN4JXUNnL1WEM2F+2R+Pej6gpraygRypX7OmZV
Vw/dziWY441O8ruaRwnoi93CuDstoyBdHNWYRHSvucGJ+KYGVpz5ff9NRtd6F0Ab
jgkwbuuzP2spBNi2o9KDwzEPZH03UYxplnh/9wEDbBlF6Ipd592p7Q8CRIa11C5d
X5HjqamlaDtIxmCsNmXltMp6AmZk59wYthJHyH8aFZVeCneEdhMM6CbghSaXD1sT
TQrjLKkmgb8EpdV7lY55kTZvzpHOsi+d7Vw9lHrevYo9ofF9SSdqLMQ9C3rf9o4+
S2tiBnPd314++Xg6kic+1aTZd6JagDu9CW0yWGXiuymocwLmoehNBII6Tn2G0g+M
5susUFlWrCP+d0ypmZmJur1ywGXdJ7KYD4v9g1y5mrRFTEVvmtbrFXeJC4g6hoe1
uXw6dKShiBXJZhgSO0egrhKiMOz7I0GwB8Po+9CKQvou+xNuVrDy0VWmzZABvnl3
P3b65TWwxghiiz2aZQQ6eYk0N8RYdbYylcPYjQTdKHuyBAdnfTgEYU11kwVWQJ5s
JrlAhIDSLbGQKktnJi6/uKLF/DWWEbiPGwbVj4IcNBgS5tqxSuRIj0w7wkyQpVuC
UduPPKOTxgG+RPGWbgNI0f0lBBpNt9qQLjF7m5VYpEycVu7ijwyweQHK6q5+tF24
gO2wtHTa5ay1v40S4LwlwPBx/0/jKF9KNY51EdoLEkjitZDWWkN45DC9A+9e0RR7
02TZ7IB1w1//YcOc9nXLMKlyGSoQOxkvxXNI4iRwQgD/t/sn5nXbJacoQZJgmMqS
uLM3FVg947DmeklmEbkF6aX0DwZxVF+74L41mc2grxsk5eM93wsuqCVaz2NyXx4m
ENj6DhFC1vFD2FPr4aOZ/45jul7vtVUAXGELHQV2FfZVTWAljqMAMuIuL1EXHIYy
3mrgdD2buBA+o+WNPLho8BE1JJlO09TlHI0Qj3qAbOoAT9ov5rxrZuPIqkZugUpg
ta2bMh4uqtBdGLn2pNaeH7jl04QI0rTknS+d2L/bDC2Uw+bm1/Ry8SezsPdRTQQi
AUCdm3nYy6NUnM08oyJQ9bk/HNuM7TRYU6W5xpp2zytwAotVfAQTTFdurrb0Fd/7
Wtd0ls/TVRoneCEEB49cso71NqJhMKfYFhfCgR/qc3Fv9lBn9lyfwEPc/Y/bNWkq
u1sILyuyQr3FwASxunUpHkmoDeIUn6gnhZeQd+1GbkVQbVKKnjZ2D7SZrFtyd3CD
OcZXL7L3CPWSW8Gu5qOXKKsr76lMv03Kom40fgq9qqQ3T6a4mbdykF/J7N6tW0w8
9t1oAhzeF/IzjopDxhM+bxnrZCnW6js4g3YerbxgOIv6nT5rOiPESjFv4Zu+NMjn
DjR2l9vRzXamE6fYNNBm8IpBLN3667agTYQi/oB/ITbnfZU/+tT/X0d2V4FVKuQ4
iEPCHXpaAHrbcD2NlHTfGrWxWDNdHl3MUvLdHjohOmRwyU4R+SMRGGrh9QkAMQf0
f57Js4yWQnrHj0we0dHoH5IcAadpvkMU37AkR6wf9KxkOVXvq2/kz5m5o/2n1VMi
WaqFnnmka20tSBdN5mJJOZU9K6ijXLItCZ+m3I6iSsXKwMt+Ix9uV/v56SN9dR0J
lzTWhDLghxFU+NNfA9+yUyN2eEaVjrvKVxm5Nj+4YEKjPXndOj3GogunGhhScx1g
BEvjcHWoF19CreFzbmmBa+B9VgSb5yRav6/Nhu9pDbUVjd8lspvDBjZ0oA0E67zK
f89oP8EQUBYvLGyIVLkwdnCvHAvO7u4BYyzirrgdSNO4Hmj1kxzk9M+f/8rlYart
pIF748vzQbmeRjgyVW4meU89NnVLHYp7MoMGtbVj/6tl4EHiZYKF23PH60DVk430
bVKSWEytRpluiqW+6lMNtb1PU2inOPqE3un2XnhH/GxTqyi6EU5y3whNQIW3WuYp
rz+UzU7S2grdMR1V7Z8GQwlcjQ98C1myD8mb6CILMe2btobSz4B2nSAJ/pqCssbW
izXtupAoHWCJAXNLFk82x3mVv4VL1GACR3s9kAAbX7RMg5we2MsKUHs2qyID5MyD
y0y03c4HXdrEwfXurt+FEGJJPPjT4hVNmatNa4IWOM0O70KvGba3Uit/tV1W4GN7
qy9Q8Q2pEPXwVmCaA0wEagLXdcbFXVnST2tN0vrswFnGsdlee7hBPO84tMo2FCsO
wxun/+GGIJmej6sn6aST4l/f7q7TQ/j1dw4L/Srx0zDiO6F3vo/5CpkViV4OgnTZ
vc8a1yov5r4+GvoAGSwaC3S01Z+HMtjx1pJcHL27CoVma1jK7P28ZnV4bULOAa9I
lTibZ3NJB4JyrhFQub4c2dDvO+zEsctYDhyXGCF5SRklfH4bBTONkubip6sx694v
qFmcaMQ9TimvFH8iquLPP8OF7vo7LKcfhnF2O1UC2klHf3QAdqhd8QtWM3HQiC1N
YBpxdbtm3lehuk1R9g16zR6aYOzReVRcoPimEcsD9tp05U2j+oRG0WG2S9iO3U69
izXLIWaLJ+hWfRceyg+ChS59jvXKkhdD+JeUROBKA1BzKUhgVOhpGB0SxuhIMydI
blDIORfFH6O68KwPeQuBxdy7oYwIzvlmSEX3Zjj+bwbf3ZnmSQcbQ9PQrMbSjXX3
70cMK8XU1VK1hhlSn1uEFKsYpideyZqu1/lDYUfiAJG/KJ2lK9Rr7J2ISuEnbUvu
NkisCFQxqXlwX8RbNjPtrlOdqUQVrMIHSjbTVLYhRWh7++3AYX4UmxTpajaPvoje
e208SMSCMHO31Cki9QlWSGawUe/zn5P1nzO1lngnh7QAl1lOROtKUcEOt0cD36HZ
nvepDRiUdWGolwr4t3j5iHL6kRLyaBLvX+4fa8NBzZ7QzI6JEfsg9iFGRZ/It8AQ
P0TN/Mn22qzLEsoHsxwHnq5JYmj63aVTKhr7A2z/Vte6uQj+iL3F7S3na7RPCLZm
76TWjiAk1qGnrMg+W5dWAlQTmewKTurh4gLi6ggpe4dTY26Ek7vH6S7DJvF+AP2k
YQ8FZXgBVYWo/mxqCjL0HrKUaNO3qZ7Vnlc+Lxz72OkIVJSk6WKe1jzKPrpgmP5R
lEPvP1tziK26gAv+MTaZpSrW9lcHui26My41jArbvSQMZaNBY/0HOqKA45uw5god
VgA5Cv5fxwHpHiGSSk5PELGET3cM6HAfQvqFOWXdFq+nPo3M52p1IOeTl7dkx9rB
RtX3vdcMA1ARtvqAXp5g5gNvZU53UXigoU0+mBjPYwyF3tmRzQZb59KVhHSFA1Yc
HafiC20X60mFxTxczRC0Pa7ycNgm4HNQ8qjNE+MGktMZ+W3A6PyAFkPjboFrIAPy
7g8sbJF5zZt10C/lb7Q3DbCONkU8ypQMwuDNp1x8ldogJkwfCoychdf6b6Rh1Mh4
PU26ybk7iX8HhakVfOvHY6X3juXDtColsvXhHH3Z+rqSaKYRUKzUS2XTwxWeDEHI
3oPCU+TSk9jHo8dw4b8JsNusifWyuKhF5+Y5MkQyKtNoRSU4392DrXx3+38AWIOo
8dYmZFOPg8zb5k1uYPaTLuwAYWTgpBLK71W/f5wGEnrRDOocRYUoDbP4rKWl3Pso
rgUSLQAJPjNFAB8ZCcFtoQhoD4+4Ba8z8bCTW6VnjvFZ8Pd1gpa0ClOzAj/DDT7C
ju5mBSNzwGY2mNZligrA3DHVCd6D24xeopFu4+t9Put9lpoKiPSr2v90XeFnhCm+
upkNkzaDvxGmWpmhtq/xPUbwzN0CMdynl+7WWMSqjLGD1ggGxQpjYQ4piGyYoI2C
L31lZQ6ySazNvfKLq/IfLbbJuXj0xKrtPwMEqrH+4Z3sI1NFy9ePIFvT+A3QbU8W
4jagIxc1EXieuE+CfxzSHvZKzSjBRvtbp2tRw+14H9dhLXnzlkls6F3qkIfch2uG
7YptL1T8Z19DxMoC7LA5HJ3eaKQbwTbJ9/QDx0m3JaefZX30ObQcQcvUU/V/sHb0
40QY2as6Bz7/5ITSdTinvDJHiMvSqMAzJZMDO9+9WkvjBy2pTRWvSAdy8F0o0PSJ
NjUa6wntN39A5oXZ1RksKvQgxtde+c3fwHFyILJNorBFT4I1VbfGmCoQ7Cfcp1C3
i8sj9dd4BLr0l1GsvS/kW7Pn893N/Z77xLb0BfYe/SHA9e8D0/Tjo++7MvgVVZDJ
4KX95szQ43qSaydr/R7Vb1KWRs8FgyPhwTtZ4YDqmwlFgwi4x9CBEK58+kL0gK+i
lBO2v2auCjPJdDiTiX4h7ON9RghWCbQHa8QFiupSiL3PKsqYIUXUm8HqoY8NWSzK
Qk9UxT0fNIEIQbMzU8r37hHZJnpeNEQIX1P1av6LXy/BmG9RK1LwxzOd5WB1sciF
I5zUFU4OGi4VUSvdxCLw4YnFLbBZ/D0OEDKxOIFBM1eC6nYuwCbhORggl/+BaH8q
tEQU6+6q/GEG/g7b/PNo5KUJCKR3sUarTVb/KoL1wsvJgSKJ5svY66qt5Ajo3WKH
Jfa5DFcSck+z8yYQa+pO7SDSsWbwFpv8DaSO4bJP8lD179fA80wA3FoodRL0heqC
BCf3hj3iryQ7+M9wDykM+qCn55/It57plCv2IpOvyD/GAPsRooOVpUwvNRNCP7c6
zOp3mOLYXFpMDZmt6WTftCWZkaEY/dpNoRbufxcLrl6jw90p5jH2RBzrLo/8Rwsw
iSeYZzTS+YFoZTwCFE8LaYNm8FW1SJjR2HNmZEZaS1gAA1MTl4sya4bNx4nnWDZQ
h8CfwDb2FPO9Y4tPwzBYik5P5sapGEkKeINHTAPi1QRXBt32PfuGWMD4pYtS/N1r
JTWmWDdS22o68P5DA8Ig8wx9Hcx1inx23vuQ5FIBi69eDUcg1Ja9ftpU6DB1nZyW
DHzUsS0NfiLPp5eldyWa8WLt+9GcmeXONPsogV2gyj/lZswkkbP+WNGluc4hoxTk
04EIAJ2Nr1He3zFxV/r+eCXPbeXuKYubX9h5teQ8ChgOghcJFd/C9+IvLc+mxWWv
o20DGV0YKcNtPsNvlMgc/ES7EIIbh7Bd0ZTTVHLL+KPLNtSnoT7EQVm/Oqe/wryI
OQd9fzf+jKqPHWuK2UXp+biSIaeqstvPYKRyjUaPoLCQG6QRei1xKjxq4aJ+e04D
zYNjr0mz5WllfUHPyzUos+5SkKa8c8cr3CzfAP+wvcy9ieHfKzT0ZB8xaxfKzW0t
HBdzswvdrMxf7Py3N+fOQJRnp0rZTBN5oi+WXfAwYFtKs8L2kZDhzakRmIbKV5o2
8DyqyDApbWCK6iu2xjd1d5FQzfK5KPGu5RQLHOI1OeAJJd77X7d37+PaiVYN0T5l
YpefCXPTvcddteaN+Pms22Swks7hnk9CH6bMVwzWeKClvC1g7YCaFIlIV8+wMfpw
F6N+bIWgA1K6q2jFRHgVM9StE3qswNExW/Uc9k/gwBz+zEZ+dYtpFfmvaFL1/GJi
AGgCMRPLriji89f9jJNi0AkO7oKgj2SmHDU51siLjvcqk/8qck5i/tBMVIFOnXRv
Kh1fRipCn8F8jj1+nXWhVB6+FF2m7pUpfgKjxJfEBnq0F+C6rTMuw5b3L2uHRi3D
otkNS3+NZAF9w3JMSDBB8cy/b+NnPQOQef+r1FDKCnpf1fhQOqXqPlyfA2rUfFJO
zm1hAWIu6waEZIXYBbqWiMp/waO9JYOII5+rPm8T3CUIHSM/axoM5pm+BNHfrE7z
5w/MQFfQEW9ptI/EwIWJPtZsf0Qvk48Bowm47HzqvZ4M1KlqbY/mUydImcORYuvp
ZjZs/V6wXLJvnzE0t99/kiN2xcAN+4TNWmXbLY8F00iHQSfd+mr7aJZ7F3R3DGrz
yIljKuaR7XZBe/wbMAS2wWsGBp8C/dEduTCO0Mx+R4tIsDfWnCIqaHDcOiE9gP2A
vK/50U/mJt/et0uJz2QcXIK+rTz2LA1c7Z+HJlO2x89uFSnV9A6r3LZ1PpjJvrgR
U6PPUlgSxU/uztS+Sf6Usq44/ocLXCasM7zh371UyNOwq9k82S0pm7Vmb1zVG3qP
qu2Vi6MqIa0riRBEHsuOZL9x2UCMswLBrGp5FbjEQAIgyq9M4nXriOUDhkOAhgLc
jQmXpwDODug0XwZAkmNDiXfY4g/8J/jwdF5RJQ/aS55G5MRsn1R7BbP0CQzbTR6e
R3dpomxPDvld3X3x5xX3onvHjlj5d9yizg+bCwsR2NwXcB/hHFqO4xBtXSSke8sr
VZqo5hC/T4CxfYeZAMvYv+0o2EJskPesSgaOsShNsbGCVJeZjJ1674q5vozR7sqq
/DYvbUKeSzCXrjnro+ZqmBXC/mieuC09Yall6BHOL4WvKqqfz4pwYB+INfROnCtA
/txpN237cXLnvPypQR4bwVMFtnJdoEdtsBrMy7g6wgjypnvfSYSwirl+bQYN8d1v
ICYef2ZUnKR3k+/BTws3G83SwsQIevWeyVBOH1Jkq2sGr0q7qtcNz+IpD6cE7vbo
JnJlOajCdlAcHTn7wx1b7cJVsi3cwsjclbpmMP7IlYK4nYzRD7KZXVrZkhRzZwET
48mQPXGr+kEyDeAm8Ggn7EYxUlKmAKio82zWOpNNuezFwFgRFk5SdTDB7/CmedLx
/iHN8/WBvjUm5m3SXp887GAsHrZOBwR2kWV7+jrMeA1g6BZWgfEZ3SAaewUb/MKV
8GyEpbn7Cjt9vKpzyJpgc7Y7TyOlzjgY4LvUcefvcQhXNEcRWNrMgHOOSIPF4jkV
NaJua86a3jEptmxwXS7Q7dnbZKm+qBjpH5UzKZ2JGOYMeoiHtaE/kK16a/8RU1yZ
suhI+NxwkHcl2RB+7OWPiZAzhEmDE8PMXaOypoW3B1i6hee9o1GhqtNW1feTtmqV
7XQ0pcUxkJPfwW4stWOKczJFoOapoqwoudn+kJPPOcUE1K5L4uPPDI9ZXfKnPmC5
/lcr4bNBvulXCScm/2/LDKQxTr69on+ZQV1vFIfgx6I9IS0Bp3zttwR2ZipteTlF
DOK6aA6LqEpI22Uz9+E7VGNFyV5tt2ieze0Mf4Qr4hAvUwD1aQyVFspwln91B0Gp
I71mAFwqF4A16eMdDJzzggY592/UTImzaPcEbVnIKh+MY3HCKspNH7Sqyp6dvPYC
AgkpI0zX4Ran8iriDe5viJ7zydlkQ9QQ8Mv0KSRa5okQhKlvoEIKYs26617up4mn
cUTolfXFylHmuYw6kMk5fxEYqCrRS4y37I/ZzXAjRV8h9UlutrL/TX7C9NfONb/d
w04Bfdmkyc+hc49w0XqtAmIIwDhYPfGggayp6ukBUuG4obpRCH3fvOpEfHaG0N13
/v5LagZ7sWppc/tc8YrILSylyUagbNDfr6F+VNzYSWRT+XiFf+wzD4UElu+LXRPh
i+Gbv9Te75Qj1+VnxCoiQqFiOQFBI7N7XbesvrJrN4cjC4OrUDHjapcKMCk9gJjH
w//6ayzFo+0LUbFF1zb6IFXxhBaRx1c00DEQV7/V9/Q5adzAeqHChGdN51MvysmM
mhllqt/eLg4GG9YN0etELt5IZG9atTBZ/RFOEtXy/GAHH6g0IG7py7fsVYDJS2MN
sK/9GeUazJiSQcwmmjZY4nv/58/vd4eSDHXWUTRJzFTUHEiV6F55FW/3hksqVupH
RySS6+9vs5kXapYFmrmoOVdwCgVyU5gKbFIQmgeIyHcq9O0FiNKDbRhYC1MbCGo1
0TpET6Lz0qWm/TKA8RurSJ4uq/P/dfycLkSTsc8SP5UpahAtznmZkNmhMbdizQZn
ejRB5cD29uA4bd9gnQtSwVF7K4RRwehxUO6i5VVkfdEnqr4C4ezRLGAZRSEvV3fN
nAfO6F0EGaGxGXHb74F9yRHq6oinubbJlHKKsZVlApAL8RNJGzFUKyke4n0/qkR2
4djnhfq00glqJtJvkAa8I6v0uaJmce7ieV6jyWYmRh6AB0ABrijMV8X5rDpt+ViB
lrVsJ9atDUIM8p/fyuKnfMvtR8wcf4LMoZPVFOvDcD/SD1+z7xcJ5tHqXmad6yXx
ia6Gj3XNuTHhRpOZ38geg0Pcw7nDXRFDhlGr/L1j4QM=
`pragma protect end_protected
