library verilog;
use verilog.vl_types.all;
entity mux_2_vlg_vec_tst is
end mux_2_vlg_vec_tst;
