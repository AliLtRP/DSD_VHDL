// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:43 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
svA5EVWFbKQRqu/t19q6SnaeNhJiu3Pz4B8RSfsNimxPQUoOPSpOnG9U37GCptQz
/Hts75lwoBBmjGTZyaPI1KcxrzfWmoG2QEoEJqORBprK4nvrPzjQ/KXECy4niDp6
I2KAA9N0COD/4Tdtk1O/WLJdOsRG7ceCPgyTGySSsTE=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 46288)
FhqIko3hHhGzm2LQIhYzNmjLevrSOguyT27H6I10vRPmNuP8zjwU3zCo89Iz7+LY
L+o246C/lCyZpJlsf5RMPFPhHOjMd6OS+AHmiNMy9eMYcUUSfWIoth2Ss/cgutAU
+HtH14tLvUgueb8WXqqkbkhM2rQF92XKBeiAiFL1vOX3CRgkw1w4bWsG2+DlZsyk
N9jxDBnEu5h2G4ychex+DBGfGqr8O+EBmO+ucQplGCR3gAwtyB277iORbGVdZ8eb
ONP/BUJOJ0dVckwu0GDqcFWU/TCWQBSUroNN52CM4zt27nUp2skOre2tYq3MqM5a
hgVpqaloiu2w6Ic/1tTJhBSWQ3KjHeXWEyK3YropjFklW76C8ief9Dp3lCS+OSM2
o8Q/wIwY3qAtUFZTBv/Z56oUuZgPzShRSZPhMF4F63QVGThQu8LTAgMERBN4Mzj4
vzmTHWzT0J/Ys/rjDsl4mTRqYfJwA7BR0cnmnD8qQrWyWOx0aYqAyQPlvE1DjNCL
Ml5SEy5ZYK9wpWoj7xR6hdRb842PX92FdtXitUSD6ROEwc4zYM+Zkyg/Xz94Rj/j
k+McnCdLyKfxhFdxOlVIK/AhwIhpw7MMqkYegJhtjb8uX+n/1gLqa1j4SFxXYmsb
yXj0mblBKSCYJoPudZP+OazCFJxZfFGCBQsLJpsgvrS142vwT1G49AmlveYEAYpZ
8ZX/hxRP8J5jgNWe+3RNcxbvjBwquerWQ8E8st1KyXNErHxIq+VAHp6UeizPP7Vc
HuBxmC/BFvVizI8d7Da8wavLshwyMmSTGQbjqOANalz+e4XO1390OSIKt4oqgB7x
lbqZI2ZqGHTXCodhjBPydsnsKpotxVFP922LKXqscrp4VQJiPVQfH3oEzxrFLoiS
4L9KuSoJNk6QLPfW/pbiWA0Z/ek+iSFKoziSbZle4aSGoIoB49aycy+TUKdtIdgL
R9xdGtDjnYGtYBDTDPOKRMuO0gxGN5CW4rifUcH9gavCWn1Z3kJ5aWUQs5jd4P5u
McpH1+r+El0uyd72iwhu7h6H9my+BKPPJRHhwZNpf+ejYX5r8jpg9x29fPyvFkiw
+kq76HtBGpFtYvmy+vKHEPbqJ+/8c8B8I+QblwIqex5Dmh2/kz0aN9DFz/I7MGv4
Vy6p7GjUaBSJ8JnnkJzFIDnYbHOYa2g5CEMuah0cJVBBRng4UIJ7xamVE/qgMAbJ
oFMSm/MkBPey5SA8GMp6sdBNeU6hMDMeL7QrvnPIqGJRTmhVrXa9ZNi4V5/ZovaW
Qh+hOrj1jboVsvRxlciMUlDB3HRl0aFV7CW/z8ooyOlBQourYD2WZrt0Xl1g+Gjh
gWDH6nM26NIfl2bC74qHwMsW6ap2kydWWwo62/gsAukE9WIshqKEAgtuiI+hmtad
x77BpF8S4cjWRzJGUT66RPiEXX4E/djSd/1MCIJpf8m1OaAFWKx4qdEMen+TRave
zDf44cqrf3azu+aU+xk9Id2mM4wFQkhTQlonxNKxqc4NfBgKa0nEOlAWY/Vq7Cwn
CKZRWws3/IUAsjgFR+nbf9VKxHpCtmL9CLRt4ZGOx5GDRZy6ov2itVMl4htc2mJf
Ze1IvHtwb2iyqRU7LSgGTqyjF35RztK8TdyzGO0M8HC1SEiuxRoRjlOvNtfortib
cyLnFuiMjdm/17bX6Jwe1L2ZfqsRGTIeBqgcKdM2J/+LZ9IHp8amrHTqkCNyitcW
qHV11zblBLCzEItcCIgs5YUBcrKjd4IfufFJNCCNuz0CRp3M80GiUHJO+3DQBu0B
p+QT4+PiyFtAkIGbzz91hzgxuWYx2nGrbboP1VM2hzq3Y9NXngv3d2TY2vUEabDf
plvxokkniWz/a7rCMMXQ5BxWNdlYD4RIVrkTzikdGdoCdvxKlBmw7Rz4gkE7qAQZ
wH4eUwohRqV9tjmkRfhrf2Gg+NB2Z7LbnbwjCsFsk1UVeuBYo2ot+yLpyjCirgWY
c8VYEenhoFvm9omw5I+0n5aJoLU7/5V0d2iJVtbnJIE36ohfjEC2BLEeCfgQC8/c
VwNK2Im4PqQ3v1lVAhnw0UOkPnOjJxqyWNla4MB26oysWhKsvuZscBmr49J3Y+7c
3gaWaoabocMs4uRzIO6lovJPdSgA2sNrqMnEay7aL27BTa6c+ynDiDfCVYqcOwqZ
SpWDBiold6849bP7f04AUsU6/vsVo1cxyw977tHEdEv+wySeKyDbCpufSb7wrs8h
pQDfVd6Q+8UmT+wAebzXO0/5Wu8smIBu7ibDyokOvi64lDGSJ2m0aPpjJPGWXCdR
9GqfXayn7LkcTqrCU6b11D0klaM0zz2BrnCUjQGygANi7IAv77O09nHDExibxrt/
8xw69CN/EwFH7MiIhsjc/sDGADl0nbfSiC6qVVS10uBkPYQLuTCx76dX8eUxmaC3
eMbjG3CGHes292Mh/3feWphqSuhKZe7hjYEdVEKf+jAQHB5T6kICaPCmuamb6Im9
2iFOstVsKAk2GWey07OyiOaJHA8oNzqIdeymjOjqnKtd4DXUmzmH2tvAXEZEKp4o
/wvo4N5ck2KDpRsfyuroFATI/suAe/CwEIBE+Kj27NvyoTzTHtu42Y/bPmleSDAq
GkBfzpnx29JF/39Rdf6MwNC5aQPwn/cn34Mp1AAFfxVySrKb1/k/QN9qZBjXo7s+
2VEzZ7Tfz1/oagRTkwPCxAz7mpGSWPGr4NrS1DxqiD7iPu6NXVQc4fzod65MHRNM
RaNHsYZd5xpEZ/QswgtOYMr+szvqbZVipxgnjhbh56h+hAqt5vlfmSDcgwepH9yn
H8gjPdr9ztIoHBM5Hb9PpPRpjso24yyGdoYUXK/fjRz5mzyiop3mw/DVe7CHTAMI
p6mYGTxXqi0Ln5zYVPe8UrPTmF1T6EBRMKihj3P43NWLN2DpK5aQziyTlC2WXP5z
6jSqs9JsIPkj3O7OB645xE5AekAIS9w4+i3natqu/y+PwjUt8n8crEKAAlOGuWl7
RqsKCsj/wZ1ksSfM5jrouAFZoGK5B3BqIYqZqu9UVPEVTyuKhVeVqBE28aAh+sj9
/P5daZNTwGrb0n53D3Kv9EbeYMi+o8mt7l4FPy8s535/1t5bSn6BQu6szvo2AaK1
lQOFVoaCQaCz+mqI+21AwZ983A9HxGr6ZzaMaOuQO/ZdpWnTVGEvXaETaTre85Rz
JM74+PiurXkpdPmsXlv7ORDhGrBwXnWLlt/sK1GyOeC14HyvcaOycDMiACzPdEtP
7xguWJAVfjYfijbDOvcU0ni0h5FSg7tgky1oZpkikEYPbJACXi5HsMr6O0S5BFW8
10hvGBVcGi04/eF/MLKwXn1QeWvKS9OvDo4LAUXcPEAIFUw3COg4S9sZYIiO5yh+
fZKvleBacpDcXff93VPsaSsBdLpZ6KmOYvInM2cuXUGXLK7cyBMXEVJwk10YwFFs
wlbe96bwNzfEURAHnxc4o9t9dXSfUvxY1FqPFWI9yNsWsrpiYF+sjItoNyZ2WHOn
6CZ8unBnLaD82AsxfW9BdTAqO05Smv/JlhrItm9IRJ+UtuexJMhu6OiU4gCkc34o
1WdXcQ3xtqZqVgfCxC2IlyBjYF196KLn8IRTvAr4koJBrI5WS5khI3ShM+yNSjFr
PYQb+a4cmz+Zgiio9wqMsl/sdturAgJhoIwPjS0IkQdhwhtEyvdYijSTe/dPSFda
WVGuKf93cqwk2M1Il6gei0bAFjzR98wd49O9aIjrs7xnjxatF2cNRnwGH2Tf1hdk
fvH8HITk0eoTdeEb1CCpTvbD49Vqq1Brg6tiiwvyn9x+vy9M6CQxg+wbqvY75BU+
SbpeSjrkXRQOTvf/9OreLzGAhF4MET2jSaGnq7n9neJD4G3V9CvjYC5Omqhcuf3f
CUrQC3nt8v0G1mBKENK5zlrjQ8fU+0KK++PFvg3xw8MyyyQ/oW4JiZq8uzwzN4lF
scrffJ6fxDeMom2QxL+CmAJckY/5d9aeU1Gp+D1pwh+Y4G9RjZu5dNj3A2Lxodw2
NgrQpddOOPF0DE0KQeQCrFA6gLw3zuskELaAhGTQQ0/ar9dwpASvSR9hAB6rCoT7
8vFZFYzq21qgID2klypm2cB5IldMEULPjSbwoE7CK5Vylr0PnpjIYR4ymM5wV7yX
S8iawAgQy4GZKKFlhD5o5EEuYme5GPdST8/2RGgc37xROxbzVjAVw5gyrQopbpLd
5fhmFbcwxTk9N0DXAML1mT8LvzHVKJWp+LyJQXg4aTpjDRsVfamVyEPSDdFvG8c5
Tuin7NsQSAlkhxg+MbfYqkxUavr8rIv14bIMocMRaeGiVeEgggE7I57QiWW/f7JB
z2T5LnVCLEDW2aoI7syRyXAGIkWhFzUd0+Q9B1XzEvsCZFP6v75Ub5F8O5l1PBBy
sk8kyFNd9oRWKpc7bJ01pWmFfHgbZHIGpAjKe34z7hAYIemwHcRJIi36yTSGdGY5
scKRlguJjBrSwjspWqRZVLwDhdfP8v89sx/xGjf5FfiKWChxwpyyvyhx1vBy9U5o
eroQh9Qd0sUCG2PBOvkalGxB9XJYXO9UDgnattOkRoj1Ep6qWw2bzKOsq90Ita5U
sFjts2jiKzXJM4Vm453tHevAqxTvdkJaOL5Qe3p/y1oy8kNdMp+MMhsInK7eSe+E
morBhiYYjD2x9YWGce2lTIwn9isJdosgW+3v7JB8EO/CdK472KCpWyskFMLJGFvy
gUwIbBuGpNdPL6mNn8F7NkKbSsMVhNPSok5Hi7DHGTOHMV63fKQrOKWpSPqef12Y
0D9s2hJfoG2N9ZY5O0Wv5nAmQt8MK1v+I5jgWExCEpYmdkXpuC63o8G92YV5R2Ns
L1WnRI6XKm+kQoGPwjPCScBFZ9fWnuhFSfzleHQ8fElwx8r+RQqplw9QwaEMIYq2
2z+ms3Lwp+zcY9nlJp9PxzYPUHlU/rA94f8jb7lPCNcrhSoREk7sTVeOKUOsDztU
NLDpg7OtaiwLAn6upVvrRRV5rMEOIOLQT2tbdRxDw/p1oRb7J+vZHJwFmTcTtOeb
uiVItyhRCS8SWmsUJDYx8e1WCw9yA2tZGQABlWi+rqsf3t7lMN4Np4qXnYxA7k/Q
wB6u0XkTThzZPyrOcYg5iDwbp9af4/ix3muI3ddJqFmQgN0OvXF74kUjC0yPJYUT
1lVYOdZLDPUMSQ6Tm/HoXCabyaow/k5V3CIF4jCZ08PrQtnZJRFNYgizbhixJE6Y
1j72gZqaems5hgotV03Gg9O1lj33e6xkWpDJLWX9Tm3XeWs0O7EPSx6ypghzl70F
tT+zvcOvFLwLmqRJ+PVaKHLhYOn1S/sH+6Vap5uQ2iYLLtDeuNuD4aXqCRfyDzLY
Vd6xIdHTVFJLfpOOEB/nYre3nAsffFV2Oh+6r3Tt46sXjyFP10bLie+YtaIZku5Y
dtlgp2ktTfRJfWnAJOnrB67xvWlGqry2L1eYJ0Xhuk5r4m7muNhaNU/5M7uU7E6n
50ziL55Y97mSNgPR8ABS6pEZyZePS3r/9vFlioMa0FmRXL91YjU/UcvV/WJUZzrU
+iMWB+aT339OhtVRj7Nn3FAb4V8Jvq04t6NILkBx0Ksxov7nJkMkMxwCZmbkvS0Y
pdIrmKivXBBRzM0QBkGYGaZ3vZ725ZOPO0tIT+Y0UqQSbWzRCfZwr5OMHY01pmCx
o6hS0OWxQm6H8dax5XXjZUNqESpoaTFERSfk0Sl8shGa681i3eZDr3P8DirnMugp
S4Tf4P4po9sBe2hw8tVj1pM5bB5k2sQ9dD4olHBuf9tbQGZHxjevVLoUMRDS/KkN
jSK9EHB9xlf66SAUwiL0gpWza/y5JLyztH/HC7O6zLc1lCUOHutp8GTMK67jbTcS
sE8WzIAMxBKMM249fne73KcrRIVVSR8HuALQV6W6O+W3i9mN5UOpQVr3Kk7isE3A
bg7gHuwkm8X7ZzDW6deqzbXzWORwrYDm/2D7zKQC0h+maqijcZqmmZM17nzDbS/1
nOT2bojI0sPAg6nSqQvbMEl3SSsFD8WIackxXZf0maBq0YEFVahSasY0xx+ZCfRh
HjJVujYwcbx8P9TWtSr8vGQzsc/6o5wFBhfElKBf5GLwNkXQFefRrBKC9YiLhzFV
TTA/K1eGtAPWY/dh/5fkOEEUG3ZEZz8vZXwF7Q+y2C0TBj49YhADWTUNC41KxP2D
6z1tIbyB4cHbjMC8xwLq1EvQtrMspR8WrHO2rCNb6sIAYoWi8ZpZ9Ilksbw5LDs+
Vf1GJFocVqVcoZ1lWtYMQV1WMAiCGkBX6q0SByct+8aJTvJAy2FBEq0Xw197GCWM
0bpscr7d8qN3Xt4hRoo/dZxm/+EGMLjtP2PrvYoWV42C8eNbKpBJmAvRkmR2khHy
Wk3WYyAwFv+GlTwCHBj6GM8l8AbPt/CSI9AjkihekGUTST8adOqtEhEPfUlxfiXc
XBRld/WyiEm1B2gPfZwl9i0ULBhqSAG3rTTdDa1rZ031U65b6I6Ip48lxZxFfwNK
oQ4C0gnpIkMY4li53rV+bdJ5naL0+O07qRVyioov/I/18Sx7NdCp3rlfEc3ZCF3C
xQeszBjyyYnUbprjxtdQcEoEAH5DvCb25Ddq3gqdm2Tc6sgEdqNaYg99v9++4FCe
lmEepFqH9qU9TdM6EKuZJ1ymNvjp12RqrP+KfOznMLtdAm5OdMymYYaC+AIgT7Ek
Vd/RhuQvPpJ3khUjGaQm57dt1Oba9kOnW/WsbglPS8IPljhG2lzGqbwqsPHuj8Ck
zsjsEnh9+VZPsl8NVosHRIYKTCI0mlIfSe+DmaAikYOO6OooE/3PJQj4p58UIAWk
QxwPOp8Z+97LlV+6WS/ulTRhTSNgcHWa/uGWSti+IVQ0NTZSKMXi69ILopgYp/8e
v6H7u5711T9aazNg/wpeWXlHc9vJOSWCIlPlJ7msW6T7Ampup3TRS20B/2So8mLG
o9wxh8DQXP7vC+x9VZp/vt/zgSwPzVCqlRWX539d2DzMae9ACwCLIanTNQ306tBk
RVC3EXblssG+c/D3m/lTcrI6dmcq5SUHwPD+1nRaSM+DknaPCTDR8cO3iBTLV16Q
8aqtp2n7y1TUm0xCa8W09azrmMf1i0s2gKsLNSROiy2498PF4qXEeDRnaNrciNlj
7OCzuA590llqWEPn2oVIDiPNk8H71SYrbGU1rsndGZ7ePOfpcvolNmNEqbD3K1gY
7qX1GERpZjgN8PcDO6tup55nX4Lz8BUdQg78u8BKswDmfkx0Ax5Y+jcUi8QEFxYd
Z922IvcMWKU/U7bx1IKr1TLsKZG3MES7Q61xFvU2tpYvBiUFzL1hjukZ7qHQY8W+
C62XF62TJtGo0Q9ay096+4K3OsmN7rZIJVh1BlbvWBleR1JPOVeYbNZe57bY1fVB
d8R/28dxYEjit893ClzzWQc4mtBsxhK4/S/kXa8Z2ldOjeS99qQnNWE0md9ieKv+
+e1FMDLKHc/BqYmcQSh634M/YcY/ekKmcmkfQavMWqtEPHjj5xWT/J8EYusoB9X7
4elRrPWJhDevlixG3ZUOptabRNsnmH3rh3PllaitDJYaF5ZmsS23Wu0v7Iu6Kt0v
NBqiWLGGQdkaaGT3xYhulWr3141aaaYNAnYx5MKujY4yF2CLfIo57W5w4DgLbV3b
aNeAtuaiwvsAE++qTc1E4nXD1H2JMwgi6EeXxH9Lbl9ol1ClxabyHAwG9f1gMNRI
5LPjEbu4kIsEB3z1hoC85Q3p61HB7RNmW5HxE/OtuSQVY57jIhazw9751vaf6rTf
vtes8QCf/GAg2E9yJg1H9yljhEPPjdGTBS1RrpJruCILDd2c6VWg/gzvFaivwqfl
e1XdOcSp72suRqVQK173dmza62rQD6Vl8mBO70TWCCO7zTIQkP90aX+JBZo/mbJB
VhS0vlpW2/7B2lC9sypWUzQGtTvyaKX/J2ilb8Ohk9oF9GGfnOZR14sQS6HfrfSe
9hGU5gS5hSDd9nDhqUGBoMXEu8Sw3GTNzruQB+MbRgrOCTq6MJhtP6N0ZI+DzFoG
e6ZPSPcVD99L0nGc1OCswG1d4g3kRj9iy5/tW4Tpbud7hHIJrum5ioeCyK6A0DqK
mA91KJ+EowxOWjmZ2wSunYtmS/M4yROAbE4kfDaFFY5Yi9OfdsI4vUtOePYgI0Rg
bRximjvi3Scs27sKT5x6oJ+hXjKgOKdedmmSd6SQkz8lVsBi+rNcdwg8xgRapBUU
XR/qEepJOyd/UZeJzYsKJI3rBtCCxkkl8gyzksj3xxADMsGwPbovjzegaVnbqaZb
5oB40GOYav+e//hlQMT6ELAEfHa29++Wc9h31eNdgd4XvS6PWmvislcQvH251eVN
36E8szHmFYGqCuxFGjNCw7KJ+a7+PlwUT+oFf1eypKU52Y1G6NlaZ792ccOY79AS
f9gnK/4JHMH/G2583SdOKhIuD4uMvoz2I7593jh0bZ6yW3mkRyr9SJRAz2ya8fLs
FjikPr4YkJ5jVu6FJEj7WyyoxXGCvt0I53+liU09r4Al/RA5vlZJlkzI3Gy0SV+F
AVUyePouhs8xH5tFCHKqTtkqhGazxOMrVPJJTG4wY/vMUxXyAQ2jHBRfbn95RQs/
bldLdHc5QsJCrW3tmD4RQgLwx8FsH/LugYFn0BkL7Lb+oLa59UBnsPJ3kWd0qrXc
QFW1V1NBMy4uXZUXfaJwnq12QoC9BqM6UINNc/T+f7plyVnfKfsEdW5IOX/gI5r6
PZpUWyG+FywoZjW4EgqUeTJMG7jWvtuXOmgmbHCjvKN5TAgzUTkk2QULMivH6K74
3H8FjCz5xpyAxj6RuAoz2mZwlFQ73DjEkLEq1Oem7sIwuzZs07L+7A6RfGb3n4xg
RUWqb4wqVywRnjX0q8JYHNz7+rqpvSHU/ARzIOf2W9CcDX3UHvTW3y9KiTgFnMjo
UlA24YplQhazZ973PKs8fXQs+eC9nkzZDlyDuBRm7XvNqnorVER2RC5etnB9AtzC
LPRZ0y3dk1pjc8oAptpCzPLUkJLnjUK39/YdX7Yeneo3zaxCWeVPjNenYBVZSFtj
JsvORxBK1uNbJLcu6W2bDECvHckPma9s/jzxyrJr71oUpZi/ds6msf8/4p7BTeBd
DncEExHieOLwsWycWQlhJsBczYZotCRKx2ooiSMtE/Pj35DSi8hr1+L4gfd+zSEe
dduLjtvINro5bdCYyLTg+6FFEJTMu7TArZNdNA5yQWSsNpEkKnvoMKUIdQ2T4BKw
BAcblvQUDqWiuftELUkr7hfLwYE/Y6JDkXIihtAvh/wlJymh8NumfQb388Mi7ZJf
HAhTs9wPlZbzVvjL7NNS8LAeQHhsJeLbJ16AyuSReGuCoOszwzUgGIg1UFdSg+//
O9/sgfSXjuLZrp82MuXU79lkCWNhTf41HvmVRce5QQGOc+dEEbZ0/UogTPg8Ng7Q
0EZgmZeMBJSaU92bFaBlINhUZ/IcXkAwIConGnwUaf/jTGtPA1vG/MJSziFJSYCq
Jdo5UMGeye/KuVQFr9X9Q1f6+yM8gmo2daHoe7NuT4AHukfQvaQMB7+LI+4IXDni
u2VhsoTuXQRm5d65q0wmnNiXiX1+JRLdXO1pd/BUBtv1daG9iPTLfOYbzTeq6a0Z
bsXD8XW8umqabKP9ToNA3/iKBA3JSoKKlMFTd8xrmZtFZMGhkCHRIEswicInD81T
Ui0bfzSGKXJ3lPd7fFAzIIJmZqsqLObOTYKkfh7xFGvarUps1Ox9MVk5qRW8J8HP
2N00NT/j1NtHNYVx+rQ179eVWvu9GyyvuYUDVaeFfA3Cs490Z2lkVPQK34tejXCK
p0NyRj2AArLwjHKOPZ21rc0LsJ8R7FyqI3luDGzrLNSDkGpwmQ1AH2mci4Q/8QE2
wSlaUsRjloe0C1RX/1XyxWc/Ybc9iAm37OnzK1/eRkELLksW9YPNu+uehjJvBGZh
tBMn7zu9frKSIa77VUvOo7uwu61JnhUPG698zqf3/puSmak+94AklTieZ60Wg6In
I3BuwoMQaQKZL6Ngwc9XW5Qpo+HfpmkKZ7yELHa9LJvo9UhI7oiNLJ/pqUNvhjAw
3ZFTIZGuIJ5g9++liLNNcHh/Op0TQDkVb8cV7q6Vm0/6iApLykZZmI2QDZf1WDUt
6vJlHNfhxSFZ8AGkViRhTi/6n3nwHicZpBKHwkdy+VKs8utSaEath/+G1vTkeUOB
2P3bI/Ia120GlmyDFvuyvDacwhNuS1TfgyiTS9HeeTgQIQQSQkcfUqnbzCR34aGB
jy3ceMU8Xf+0y2Z9x5F9jl3hyEEmseM49mklc6ETok3hoF7pM5MUGDajECR9UZa+
zFMFthbPOB5BWZvTbWVcRJjnoFJR6jJI91aLad5bf0PnOw8ulXkCjLSJFlB1SwJp
r/QMa8ri7FqGbEl1/GLC8kqq9I9MyRAQOlaK7Du4DzpxAhduT5jA/AOuWhcdcyaX
lBbh2t5PH0h1vVDPIfBl3F7zPuVu/rCF98gt2iu68YlU2LSYRwIy6imZaKN29W7X
grHeuHG8brAOUXKR4nV8H0Qk+oQAY60/5EIEMMBHa8eUT4GoTpVP6H7CGyq73r1S
NZ6yU1jyjPeTAefkJvgpMbsdE2MEiK80HX+ZMyZZ6B12Xw/mLS+POyd3QfM+15qm
GbRC/+jUX6OAvnAL2JR54+kwTA/vWleTq7HjGA2hKzMJ15NRH30lwbyM8XLJQ6C9
cM8PPF/3lVCwcx67PXBydZuEwXeFuhcmixEE+dbGQXxtjRqnsJG1J8yiENCrVGXl
0tK0DOeDnReRvkNxN+vg4lOrZk3d32HNW89MTcWXFKsZyk7YlCUDIedjet8eDPhm
YQ2AV4KJ2yeVHBedJnv66GOH3IUtChZFk4SOipXtCo0239q/crwk++j3Gq1V43V2
ogekxj9yi+Y/k+X1Z4OwO5A8UmNUbpoKDiPVyoPr3VWnl6+ckx60N1Xph1AEuFu4
OqnWdrauBQuzxTABwIS18fbPWL+UVYNqNLJGeE+2E1pX8rt+9LNVJ6u+S9CjCUR2
HMD7AtdANUWz3wT/2jQ6A7TYW3YpLI9Ry8NP4e0vTE1mdwWBTsVf5+NwSfxd6Ey6
MR5lMbmbsp7H1UVgwbUYVQ9AEzG8o9A2/GUKiBc7sGuWrsp3su0AjogmnQh0T4Mr
kQrT47g2EJcG8rPsPtMmhGM4Z7ztKbjX1LTsSg80jtqB/qvmknIJIFb99OCx7uQw
QPsL2SgHywRIuehILwoE5uegMS0THuyc2FfLNkM0aKG7kyVnuriVUA4ZdhYrOG5y
U0ShJ+uwFVvYJ1G4EX53eNehtWxbhfgv3pv6oCJcqIr2ccIAOlFzVN71MlG9o9JX
RX9mHIXL4IRnVEE2iSWopzZxPHN8qqLXfN82SNZCc1kC92j/FKBpiUi4M/+k9MAK
DFnNFl9uU61Ml4ziCr+3xxuQWTiRgisBmh3/LxDCm/Cp5ntVU3Jb3eCZ5kOUamSn
ccqVIvz5umn8SK2knvES/+Xdl8JlYyIqdAPj4uKSMHJbidWgeo83wIL9EoJd0d2c
geoZGZ5rT8ruJPfH+k2WgLCRwOgd5w5ys2BLkCj+yqEj9wWyHO0fd2PZt9iqi+Iw
tLK1lgDOZL7aFLYuzzApGYf9kLokRX1uxtXTLYmO9paSnQt9yN4FqJrnyx7/LtHF
OJUpxBuEnIE6GQS3pe79hI+A4ok/CnM6madhfobRklzBD9/3HdA8Nvjx64YEsCMz
LuN6ThfDakdM+8ZFPNv8BgBSokN+6KH8TZ86nGCBdR6xvwq1oGoM2e/JldtAZZ2I
4NTqBfwjcp9kqddyy3JEBWOk7K2XvP/TjIsYJFsJoZvS9BzBsb469v0bPhv8uiPa
lUQ4/AuWnZbS4yHF+4kli6fWbo7zjMIqK2krabPuwzpFdDPQDRQXA3PjoX9plfAV
KX0vx/gIkMB6klzDIuaLFqsJdd3oEPY3+b160y51YvfCItSBDRXSYCxI0N1Wuy/g
kBsGp0TBpFHBI/i6G9ybvnm8FNwwyH7HwXsv1zcqAJiM/BiebBK8YjPGA1U4B0WN
hk2Az3c5VmZaaeEhX9sHuN/4QEoghq18qtdqfs+rAztSqZotcZQervjr4g+N7WuS
MogamuE92uQSnlkIr2dpLqzhPDfwrr3rs5tA4iTTZT2O8Z1fSXnu2iQLViIS9O2f
FTBCf6YY1X1V4aaaa4xDsRrCPp8E0usXLG+h90FI2itkw11KsLTdhVzkvWB4mm6t
A099kBGQyt6mkeoPYf2lj7TQVS+8TdG1IAyam6fKlb0sQnA9HKGhFORUD3Qmw9p0
csDHLjqA5t5cH+Yjbo0q2aW4/JlY2HUTOpKT/xPBO05Xw0/eAd1AWBx9VM0s3Di4
THcrwOQz8NLXjh2DYwAJ/0O0YyaGdmL4/GkspRxsrfnrVTs3DWrxqLBLSGXy0X0h
0rhMHVd6CDc3TtAP4ncTxjrqzJFHQ8duiVZpPNnamMKrGxRvVHA3PuX/aiLwKVxj
DNZ4id9bHCLv8Gx0pmOWoCn3mnIOEqGom/+RBug667MBX+bghlvW9G11u7aSTKVR
LIy4hUO8+b+fj68d7IsxfcbCs6pCTnjl3ZajO+Kfb6wRrtsTYEfC6/ddMl4bMp23
84NIuugN26Rp6RXN2x300ypE7qe9i7g61l/msVAmc6ZkFACSV/61tuu/KvPVaczV
zLwslCKVZ+FPKGkFDsrxIpBffXOc9IYLC7aj9WZDyZYGzeoVYU52SWzV/uE1HC0J
mclpgewl7CBw1wTr6X5jnlUNk68wHrb26P08OeEL6iHvMHQeTvUZP+NQXifl+TWn
t/6tcZGHjXVewf9ddbsQMWLenzc7vqFqDc059OTlmo1u2ecvl0LdNhn16wwYY6sM
HKBkUsetXpOtobFVz8N4B3p1rWDFXYN0iRy6jxPdpqF19mc0hRpqa9HFvhtcIn/T
6doMjAgig99amwecLT3KYhUbBj+ojJBRe1D3Qq4A0Lwh2WCXIP7wWzvoBmfY4Dd+
RoB2jdtyUoH+A5AFs5WO51LYico4T/ce//TZbJd0qwnVK4qs7CZxHwNPZ5zdkZCY
L1X1n5aEESBQwag8SojC9HkK40873ayNwByq9poUyMwQCrhafCkwvJCDazWXL4Dr
SSulDpbhqwmoibyEKCVQlGaNtUaqHvoxIRy1CshP4jiG7GBKUd+GmYtCWSYmzUA2
dEUMmngKAhIX6cbs3Fg2dWEF3/+8ncpQQPvQ4GUecIbTfbEEUv4Pu8jzsN2vh7zg
9fFmEZ97hgQF3LETw+p/1mA66OublF11nTgWozJFnRBEMWi2GP1gDdWKp2Acq3rt
s4srVtIySbj84i1319QAOk+v3Q118wlaSBsugrcZ41jC7JI+TEN95ASFRfgLOAD3
tLpIzOjzk1IvudDqet/2Ii6B7FYF8e5eeVl/QzlZ4uuWeciIox+Cg+mgx+9nZiS1
CWwcMv0lSbrQMq7ddgwKh1ruGTC8XzUDGl68UCe0lGF0VJqkvQesrsOvGKK0BwEY
ANdvlT7GWzPwwgBvFUUMtO0ypbJPlcOGJCu2tUUV1KOICYFH/LNVDLryxsS3D8TO
1zxOKgH9eG8ehZPiNW0ymWxFThnTkThdPtF95bRF53q05RYZs6wTEjkTqNH5sbLn
JO5A/FEEqQjCKaEfNEYf7jB2yOWIvLbAQJLh5hO2aUGLcALwr9hfL0lNxS+328N5
iEk2Rv4oMHi77GJtpNpDP/hJAaIz+hyauSw4Sq1c7M88SXtPhE4T9Yy8kXlGFX2E
nUjHGCUr9/AIu+V7f9T1K0c3pGtQqPaGlQB1UcJork2qj2+pSDBjs8ldLrVVEhOm
l3hveh4Z3FhLdRF7MI7Sp+ztLACzvNdNrXvNzBJ+geLcIwgEGeXJrnVz/KkWVnXR
Ff4A5xCe72Lw3wWKfDyhIg+7w4bsOjc3U/H5Sx0TVnX1m50Gep0JHUxP0XM8hnf1
3dvIj7uuwDJQXPZeItaVeZnuMwKrDFzr9H4UePOowBJJJgnrq04sC0HBbsW/P0xO
TP8jnd+wBo9QphCD3Agw0i+Kju0a5rrXOWLmwHQn7XO2aslxgyPxsrK/ZlUUsqcg
sfdFQ900OAG4PC7Hz+lU0+VdwhLj4kH7yPPVbeTCoRIyUkpRrpXODvCkEDfua1pr
fso8g+6ZI1876GJKW1P6YmUxckJhB6Azl3lREt9LNGJ4IhOhvmYiQxatxR3iCHMk
181IFY/t0GeQoIChJ8fdLXeSx8bsrDi2Wbydp0CND6bAEj0TJNAck5EDX/lIX0Ab
5/4z1vQlHj9SDWVbBMu8K32zyClVM/Of550L1QqMsiuHwhJ5TtuWZNb6GoPG8r/h
lUzN+Sk2cmDWSqzmjm4M+hxbkSGzhBoxYX4tDYmVSY/UK393t/HVvX1+5GBPPSMl
vjuWTflTxDgIBDWsZYldxlLe4ynQaKnqzmpiErLsgBzHjwedh6Ou2/+e5ko4vnC/
l725fDKzRsuk+nekdVb2F2Gvnl5pfYIHk3fY0NjZ2Cuw2TBOAldUv6ZCB3ApKKCp
feOJ43SSegh9CbOse9BYJ3mP2S4bJDhCmMYplLYi3itUR1OjVBSOGgPPWzkuapaL
N15AQ8dkK0iMjrqmjSvQjJpk0oWnWG6vRfmxedoLlgr4uG1LzsHnDBOcpAZShHjL
keLo1Q9HOc2cO8NmAfhanmHqAHt5dGI4iEQ8n04K54NBIU3dGE2lppsQzLdNQjYV
p5NbccUIPhXdmhNIYUgjCJ4NTT0+qnrCr/i4HH8IuqXcciSIYrei3e3c5tS7YRkn
oTztKj+vBoN/lqPWuMpknaxTfPi1WxUMpe6bPeRbKbkuRpgzOKEpP+LLHsPzSYh2
qXnDBjdBS8n6KNh0bMWjRtHi0sNns+s/5IiadNKUQaDRyJFdQD2JHs8kbHgkGOcG
EvZoEBHxLnzuzlhqqiAz8UYXnX+W6JTtI6lzISmAAfFA4W9O9+Pk15NMhOyaT+cp
5EAReFzhchEEM7MJsF9HqV+p2fvR9/OsVGa25j4xCz8LcF5enzQekMmx8zmmfon+
s2yLu/QyGQP8OyxhDAvhdnZgEH/PX+SgyjUQFZOSTiizU5k7KNAeq/OgM04TZdlU
Z5vkyqrdRFEtnolV7IhBqs++UxQBagyumb5aLrGvc2mZiCVCE+8Xme1mXggjtY01
Rv3Qsc8OYoFlC6FMEUrpOFxYn1FuXJX88/qntIsFl79FXyTXyCbAVBegeAMvuxhq
aVivKPkNPbM2v1UsqS06uJ2SZbH4Wex0iLXo30g198clErefsHnDJBgVqobot6JV
xMzLkQcZCkwp6oM5TjHPKnN8IZgodP9x9iFRD/KnFV+HbcgaJXmNSiI1J0qYmCTr
LjAr40dTueV1aJfT9osmmEUmiTXKNYgaPaFM5OE7W1HbZTWOcaY40uTGtZbKc4CE
A87O38miVgwFkqkRqeRdPhFffR631LuppGikTXLKtT41Nn5q+YFT+S0+xrnUiIhJ
sxepiONgNY3Qc/02+mQanV5vm46Up5+7xxvLdlt/rm2GNjShgdk6NYTd2sUVDYkv
2dKWIjNSYtBQU4Vz28sfGBgETClFDbK9ltj1lC+GlhkBgsYH2KHQJ2RP8+yutgfm
KM/E0D5+u87fodIW4CtEkY7YMBDrffclGODdTnWDF2R5mPvOobCLE1JvuI6gfb6N
WfzHg03i91oile0PQaqyemXb24Gv7pVrhwfHpLZieljHKMexZ15W7Yz6ktgmNF2z
+Hc18Gx7UBL/nw7HoMhXpPtantaRM5JnYSlDOG9sG9e8UbEJuYs7xX20COIotOmH
piOWZAl4TBp4sk+RZlyQaDg7qOxCeXlEpzmm35U9ZxL/Xz7E2VAEnxKq77ZwM7HT
TN0MWsEm3O+GzHL/pHE6wkAa9d0qUiOQnGhu6IyVCFn5evrGRkXYbMinhCWpjv61
fP59wVdEQc++OYxdcu1VjfL+ruJF24nR0Hjjj2lhRZfTYXYIrMCS41gCIJgi8kkY
3IRP1GxmVvLXeUxeyTJiR4Kttc4uAQ/SsoiRDuaPkF3dkkqbj0DCmOP8tQYkbMhV
SmiWJktkZ76bhDMKr+6OhIsiHncbPw1rePlys85Zk8nET2ALaQNJ7fr3s1HswolV
Hq5XxTV7PhNo+4tOoyzV7YzC9a3EiiK2WMdxCmMMvB4pq34x47FeO6v4zltVDOOj
xDyD80wsg8ceastQ9LnSK3bEZD5gvzAHKiUfqvh0B6tbD9JsgoiclYruwlH+30Va
pmFb9uU7JXVXpLXmkAvlZg5DiSb/ywcXlLRibJuZQlSIGsGM0aBpfjPmGgXEWTiz
ym7DCXcMF/JSYY3pAMp9vQeDr4rKh1sybdXt2D6aDJ7XysXZXlz/WSxCR5CrS4Hf
kJaOOOEPm/Qp/pWGgeNdV9uZhOpV93JJZ4eDnGIUruFmFfHDMhUZhtimWUDQfSb8
lQzvvIT/EJKsjkhJzBG+7NbWJDiKTKsv+N8I4FjCkRF4+pnuw692LS25DYygUbTQ
q6TaPkRQnXWatpSDAEpdrj57g90qvVlNIYr0m1egQzRO6BVgxu8uSndYugQyTp9g
1K7LMYBGBX+Vy5t73s/tSSbYEb2Mjbz8SfMihIXRPuDkA8FVw0mmsIPtyb6ETl1L
JKeOZS2+WBB76tHlLtJBfR9A7Gv21UnoH9zLH0pxI5tP8geEOoZriLf4XwVmKiYE
gnAwMJr3kyKxOOWMxIJqCjh9cjoHm1VHFETi2INe1f3tSBg1aZvDkTe+U8nbC+dv
i0i0ATgxmu6Aa6P++H9RRYMZVZVq+MFGISQjNaI4vgPDlMVjUJ98wAT8tTDrk1Me
9jy2BfFbY3r2V1Re7JtCIUiC5d4e22a/T8yOxzsghRxijFk4x3hLHq1qAzXtBC05
rGqHCXFsbkzf51aR4rjWhC3jdm/tK7RCHf+cLpj2vJMmnK3yPxuIpIMazGukgtcH
2whhCp/qAL/CibkCzG/h84U8DV4quMjU8X/D4D1FRyUIHPMzPBvxzJ/+acnES4Cr
0Jf8wI+ddbF7dCRDSJIbumVe3yKoOnv3vH5Dw6COkVHiuEE410xH7dSp0C6Yx7iV
r1EnTUVRvSF7Iqh9JvfTyBUvlSDyluY/JAZ2L2Y3Nbi6ep9WblUXobBItoOC44Gz
5TocERHbCQrjYokIMF832kHx/BdVOaBp2aDMDkQ3w8QxliqDOtF3fH9E1xbGAp0b
/arY1zLPP54yhg60jNbp7cYMeyAMEVEDGL+YDT6+vOTEcERXXTCy5JNjZ2TSRKp9
X9x9KXVUzdK3a5TuHaMVBWix9qkpmPhy1LHYiovasqTnWSwR0xGWU8t5KCogkjWm
tT6UJQfNmtdXwNNetM4FrlBZkOU4rdEc/RzllPTy0FAGP63GQ3S+d0dSN6h4jmBu
YPuF2bpBR4l0Nr8cjGEFY7hrzWNFYNFNVxiihGM2f7x3jYt9pqOapy7I7svtbSO4
ITcMf4+JvwWx0oOsIXRQbKP4usAqcR6CkOhwDXIa8k63iteFwUxr0avDs7+FpwPZ
P6pAu1G43YitL5qaCgDBE0z5lig9AThn4AxMO9trDcYzGHx8QziLjkOsUlV1sUQL
4IgUBfN5a3e0OLUAlJovEvlBV/j5epNmNIEHQi6RP8KfCjRrtXP5r9KShXsKnZNp
LJODFHaS3R58+l35gCGjK5yW4VqVt76iwjj9PeHgQa1dBWyRCHDzKA6t//xcMGg3
o1XTWBJsmgP5/aA57Oya+VaNZwE4FYCC5P0gQ3EUabxaXFPu2qjyquUsV7LgJ4DE
xDmYa9cGoOI9p+rWsmmUAZsnH3m09q8cKU2fsu2WRjpFDFbCtfZWD+IYjOTdNC85
AYk3ifxTZRdEB8tsBmW+lk8VtKJ2I/Ga2Q7gfqocZiW1dTo5dc+q2umlr1jW9nCT
pXE4t2YCpvdSnNHb4f6tx5NXOZSvfbH4bC9FY3nxMtix61zwm5EI/xqnCC1O1ABt
sejmk9xUbU2SQ8xgkZwWpHlRdC1DuXAS9b6toSwI8ZIPtJDvCgoSy6lgAD7lrLgo
/Khm/+cVjtM8A+ricK52j3ocxONDfErJD4IJYgYfH9qp00Jk/b+0p04+JqWU5KS6
7Q45kNTU/I96jUh5UciK1/FTLQWQAMNJRyWgacf8dLYdHDTQIBEL4UoV4xeJx0u5
l0ATAz1eEE9HlvdN1y9ae19VnzHOdJBbgcFJt16aacQrCxrquO8phLn76YqEBXvP
gIaSDVtPSQxoXQm3K/hVtLmJnISMGAnkDI6pA8LgL7kdnPmVUYZVr4kMzgzQqNuM
t6aKPrR0MRVWCNUzOrFp7YcTBR3qFzfPUkBhjf8RWXe/vVGSIHNxnPoDMkgkJl2y
LhKMh4v7SHNpGE17HHw7xqZ5qgk3S1feWyEknnF+b2FVs3N/VWJsdGMIkurBJVk1
RMQ1WpaRjztYUTr/i2kC7jPR4gaTz3MkbW0sUHcrOJV+PcsI++VMoLCUIjrEtqAL
FUbCX1BDksHgZkxsV03b663k7jgpHYl469sl3ZG58Tm8YL8CdiDEDle9MyCtmo8u
I85P2I+gEUh0pgUuA/hnZ26awI0pPsn8pw6VKoUdUILGFIe4CgnlvCRf9boi6WIl
LmAychYe2Gep4WqSWaKE2jRgu5y6zbywgFS9RK7ZRTVR87PSMW2huYD2We8UEokO
jxbBUgvwDlq8Tf1soQCozMZ8M2G+1neWKvQHQyFPRdCBekj/SESSWAVC9abHZMUg
19J+wVF38dDb8hevhSHxXav5xa5dbpgYPip8OYv002epF0h7WA7WUY7vdpgCBMln
pNr6O3oVPjf7DrHZkjWTtivK0zs+4B5lSXlOeYO5sEele7hOr1xP20aJ4zbg/0of
ZrOQy8U8bC6HauCrO/2gABcZrfo1JpwZRPqmVLy+/w/NuiNt3cbYKE2MPpV1guEe
miWxPCDcAL2fPRdPAvXRzCsPvGmVjxtZf/IEYw1CpIFq1PX7zC9duOX0NxixNF3C
8YWGxUf6NuptP8yL3w3pkoDGCp8l72gSQRVVUH2eXbBKYNFwM/k7e3ZCDG+yqejE
A8ADLYV9sUwioFN9kc2Iqj1ZhWSuBXq9NC6GR9wEeci1ctj8K/STqeFLs/4aQ5Mn
bfeemKOeUZwQy/lEj6r0sxA6FamecGCVe5ebEJYFqNvPm1cy/AZzXmSswzyoGeS0
aPEucAwr2XQnXFVvXwez0pLpEEO8z847mRrdNPxZlHb70MiAf8f5J0/ISPbLX8Lr
/I8zsIzPVa+JKfeQP6mBd5lpD4MuOHlDm3j2cVzeUjdU6LoS6ZGgTXlcCFVU/rzh
B2KFFSvouIEAEy/QshWqk393P1QaWtXAetJF5ehclopmLotlz+kfdQ75FnmOmu5Z
dr3P3wrUwOjhHKHNT7uAmVVhOxDYGqUhe47jiKMKiacJ2Ttmpxznony0fhK5nkaB
MqpZ0nCA45wynAGJieK3b+17m2eWcsW1jq0lA7PIqDJaoXC4tak9zoWD7ZzwLCkU
mpJUkpTC9k/BF/XkPtVb2AOQ84IWaX+c0f+a/9F9Hy9R0kr440XLD2eMrAV72mw4
keOJct1fqUg0+aQZpCABoxV4lKImQo0VeO3VkCCxHVorZmclObvD2kTO+y9QJSx/
lamUZcxgtXxv9RJUzXGumOtVj28FANLwMziALQ9l3Om+SVeQEyOBCXQGISXXCjAj
7aNqcIcZqobIPvSrWe5KFeu3lC4STyqkyXfU47OcQppNLfY9QuZGHonrlVNBwDWJ
d/AOuGA2kGDdAZeb5jzasNhMvPOSBRAUD0EJyrv3YlltyZs5Q8tG/kEEtR2x7Ybo
OvDkjvFC/EcvmoubpolLbjjEXfM6amGlP1bMVOQLc7kfDQWxfWhzFV0JfwLOi1bG
dPb0Xp+gPKIVZf/twVbZgMf/PwCU6m0weBrXC9xuGUXuNuUT8rr+Q5quqbyr7xsT
PPCP8q/+zcvX90iNmhJmbQzszWK0XRdNGP5EM7wZsuHTflU2w5QLCJYfRigMIQPe
pju9aPMegeGQHvahtq++pCIRu64eHrO5/+BwU3VWTwId/ABbKYr2MqMlZIM0VHDF
9TYCQ6vfuCF/naaOwPIO0ev9rbZiXyi1YkyJLa9IzIXAWIyRHdI7IX1SnlOV9fUy
m3oRhFHid4ydKAS1VQeDu4rqYR49YJyoZ1Vbb/xU1/DS/2fWfWp8X7dwxWWXvyWl
IbJm8qfI2lOdpHgiVFLQscr5iX1yjHTkDi/0XShccNFeiSJ4W/4K/443erimc9Ui
Wja4jfyOkYAS/xRTSJ0K6HtB4ZA0n4jhr62H4dvGZpouNNYygwgXtk5zscX4N8+K
xnYyi1v7vpFmL4bSLw8u9I9hej8oVYEtFx/Cei8/aXDrspe+WQt6PmaZrq6hQVyN
eIMULem+lGAD9zV6lExER2Lvl/nAZ/W9RRudyVnTT7spcY1RFlLeMkoiP6b8KGg7
mwefo0Ma1RZBfjYHa6C/pOCoVuMwi1geC2uK2IqhkXvamdz80dy0GHWuy6agvAee
Ttf9Yin47QwcWE5y8Ay9ryp12UAo+D4Okw20ijwQ4OcVb99hPMabuLHGJr+08ds2
rcsUJw1fmHIyMjPXZqlpBe9meu6W0CmNx/eCHfJbZNyT+7RcXw6qHuiVM2j9qcfh
x02zlnijMDqFQz7jtXP/z5PKMDSm1CKniIvs+YE2m75ChTN5WetrP2WV0Th70n+0
dR1c6r3fsxF730ntUFVqls/dN/0EYem9m0Cl76+dJnxWUPSf61WLXpzi2LFl5bbQ
Ynf20xuGPMHCEQ4kIiyZYeh7/2anWrkzVfY14TyNL7Mjao9xU6IcZXbkqpRJSEPp
kUNAQLMEwz8+rkXDsWS909SKiEzV5auxBmX0JWP1RWLT53qrSpiP6rh+Uu1M82n6
nXGJufl6w5/ITj6DIoEhrbPXlxgcnLB6FtnpayvmeuFX4NsIgcYmwQK2TKn/nGVh
11S/v7NlcEHiNXJQL0zJkBVJE0CoKWnEK0+Ys3ep8/JRHpF6ZxAQgtcTaBIwswJO
oMgGX/QrSolyDWFUG6VDUsi9C+dHTomanLMDrdcUHg6Aj5D/scGOGmJR+dHoKEok
vRSO0p8MMRYWIlsOKIMjE2Ah5o0d5d5VbJmzyk+Cm3RhllQp8kMp7NJ76l2yPOkC
G6h8NWUAIZq4ETarOvLY3gzK/hSA4DKy84r4j49w+je9ozX/tfsyVBHZmA2pMsv2
/J9h1mI78inNhh5DOgQdpaVvUxkgMTfZiP+xCGoOSAixIbWwgFF1Hkkgl64Xu1HH
UbG3+hVlMKtnPFZOF/1ZbpsskEEl7Mkp7IQF4HieQojB87wXpoeVDsQsCfo4f4ei
4HVlw++XE+5DhdSBBYOwPZMuwy7/bjlhPbB+1IrYdL7SZ0JP3H+LEazs5/TUaNJu
u8lV3ch+yf7B87m38xohwIYuzy+YTeCrLAldoccYujoEqhz0gHyqFnsjievfW5Ue
bZxt+6LVZ6ibL6cWbXJ2bj7GVFbjpqnUdRHi/liUUhEUk1oRGn0TGXW1/gMl1zPK
LEP/SJF0duFZ5ka1tf4yiULXd760BtWRT0/8gPjFOnvRcf+PkLP7XLvgE16vOi5C
liXw+H0s25BqT2MxqYc32+kaQmXsqxdn3yyuAtbquQ0w6Nb3M7V0CBwuKhn3mjGZ
gYCfY205BbhPmJx/ir8gma5C2DPRyJmkDdaz8SV3hIwv7oYZn40JisY89FT4siIv
821Rjtf821G0aHsejezEKWCcmf/GCIiXxBwJLzF1PUFGEaH6B8Uy8Nh+HoIuRgue
azW53DJfK/N5KFaQAVZocWqDh4zGmT4/cFOsGz+zCGDwkLu2CUaUdPH7H9E5ghFr
4ENnIEvwncWVLarRd06yXAWgUp4vPRS3H2Tgpg0ZSLe/V+9mKT1yaEowqB/2shBc
UXxgr3IWQiHlHxvol3X7mdHIZ7eQ1qhJIhR2uZYjUNyRgMybYnEHJTPA6RwpVyUT
7ydd8/b2KuGgFvitS+M93GLPqfR0gF82xLLmkxQCJUxRD+22B9wCQw5H1iRkBFXv
RxRXN3dZgiUiWCA+KvxT7tI594XMk8WrJzjDM66fNVUbbzn8SZZWPy4zqxgntbNC
0pF+RLpp4UzshvQdolA9MK5TMPrIhnqH7UBXMprz6fc7I7GPeRZCXv6Pp0dUcuBE
t8wNQalJzD8qF61UU53uqFmEZYZWlDdkvwbOADwBeYDvyULXoQU1xAt7U3l4p1IT
BooG+utT0/0crara19mNtBy2A7mxxiAo8IXC7WBKxontOOdn4z6j+T+2EsWvSDIL
pmxJb258GxXSeQtUdJ1/ekfRrpv8PC+GfbdiTaWT1sS37oGhBwSGpwwsEw+FhtiP
fMe69sClcC5g1VDdEY75Cr32awNsj4XPaabuEh7SWl32DYfa//qltiGSQn8z2qks
QhmegZSOLs7cgdSovPk7g0meVxMrAVFySheb/f7+x+qjmc3YXaZbMbAP9K4oblC3
xChv14dI3eXG6nu1AkCTu0liw31zaq6U2Mh5Nshdf+BEqhanOjimu5XzIsgvR05S
uKK3Smq2ioVGE3PFO6u1VU1a2igU2MfXAHIWMz/0Iv9+Gn1TSFVV3EpWISMehoZM
NZ7Xs+XXDSSa3NAkFRKDKQo20HrpN7H+yArbPYEjQ2hJuhyteIWFdGGZNyLc9uzf
oxb2JNudZUSnqnSvcUaqfdptGvGzbQzBLHfVk7oj4ec7A543zlbUxRFRmDH3fjsn
W7vOEIxuCl4rS7FtF9v+dQIT6/Kkd1g84UPsqi5aEmLLr093Zjoz9ArDyUOqIZPd
xUMmdZfR75hLXNTGCKEDoqquRqTSIzaeewefMEqi20hR7+0tFgD+4J3yNRJ6gha8
ruHtFZBe5qlytStrjWBRbLxIwQHZelFHocNg6S2v66STVGkqpvsXl2/t7Y/tFkpI
UxWbYdAPciGW2DEuP1lo/MwXtI0NB70y2o/1oZmKqS8AC33J6ti87k1c5HQkd17W
G0WabjDSIEFePHoxguab9fV6++wTH2UbibvNalWca9oKscSxy9wjKi98jZk8GKX3
D8EpZkV+t5cqlrIVB1jbquhYSkSn0igKkkPjNpaz3gULNWrQOCqYaNJpt/IdF/W3
F/V6C+dvi/QMd9uYTWO/pw2wVblvSLQvmJXlUyuapaxvz2zJpRQTH61G/RoaSEUF
GKuddzfcm6TWSA5D0ZqjZPaOBA/CpTWeIPbqRgLFOfOoXDdtsiVdlHPlX5/PvNJ2
O1zxxw3kmOqWwEfl09Jule7k2ORRs8eZ58NkatduhtsFHnaz2tMe/PjVd5OxEjYS
nxeT+f626DbRXB9yme4KCeCa9PR6/FD/cU+9YJul3O/15Kxdm6zvTpdjOS0mLIxp
vMhRMOkCTxYnqWEBxO5ULuj+avb9INteQOpKWtQldYiXVhSF2jvLS73BHtaPi+YQ
mZz/azgZU9rsm+vpDozgW6GKeyH5uh18PoHqeQqrvYjnjAA100KQRug/i65WmPNA
3F6xnb8fEEu+L57rvQOb50IBdvsIsw+ZJChod25CrbTvTCmdO058TOq2DbpDeokk
ku/8CnVmxzKosNROooM2XFkb4iWFxJ9iNZXfJUTuUdoQgVUxmq71mloE07PfHzbU
xm7Gprl3VLTe0pw56tGsdm4XsPBLVfIHf9v50lWT7W7jW5/mbb5X5HBvGK6Csryk
pddhvY/p29qI4YfH/xxP2KGXfA/0vaswcPJrajEOAPPkXHKlHm/juXGg9COk5Amb
ZOmGHqTJO2MkzjNnuMoUPq7JaxUZfwWqx+0bT7vbdSTDjpgLIAqPfO6glbO4jCjm
ntXshGPdlYtjA44WLROakDOFGhGft81C6glQm2FRh0EFxtv9Cna/57A+lyoiQTFt
nilbNg6demYVUvsc7hmuCSrx1c5/gij9Fd6tRtMH8Y+3cYjPFTV7LXp99cYTR9pS
485hQguYWqNoJDwAN9FecwcjkeKs+8cnid1IYuYwXykhFrA4HN3IIF431k3NyPnK
VcfmXM7jtH7+xSRmz2wy2QtHd33U8hwhsc5+Ply/mJ7LAtrWLi6iLcpxspl0bKW9
AdFnOfFyvW56MtI10TP3OH4Coh1JHBpcGeFTTHR159+ke5XcCXVP3nOvNaSy/wF+
SF0mLe7Cq8IxyeM13Hv1xVCaBcFgk8dsq5QWL7NF7zRAhFe2gCavNjpfue1Ug4Sn
Cw6529MheROAkxaNqz2v8AOqC8exufUpW4GcFq2IrxWRJ73JXDG8ezTrflFnnIRU
zICyGhVBHWAPKxO3TC1OSz8TuUFF/zPLI5e4TpjH0CURMt5lMxUwx8MIbllhmjed
TyQZLxOVIbV7UVbu1Up2gBvlGF9voJtGGjtGncdOGP34TZCO+kD+hHwoxSv3e1RW
j/oES48I0bXBgO8g6MKL4WauPhqq1rW5czP4HSj62pSxMUGzH+Ip+pA5s3QCE3ag
m9pcAmP0h+hnAAyph18Xqm1Yg2xx8xqJSpScZJigMGYAVrgckQ/L4iZ9BohPHxw+
aUp8KgkwHiapy17tYiotM1+ItPg31iR/AiLBTfydBn+sy0wv70SThsZ8b/V13f72
8H6g+R+cieKVF0Oiz17AedYRw8wMKJJciAH7RT50cb4ud4jA47+EsejZIrhOTlSC
oJAqO/UmAeE+OLn6fvHAcz22w3ocuv58vJVeJg2uRcekug5x4rUGkj2Hv/EmZ6lp
yIBpsSYsBz9W6bwbfNTZ9zlL8kMFwFsqlZp0amUzPh/VqlJ9OEs42RkQWKYOOZKH
gz8qi4n5Ze10DalJP+UT0DICmvrA8d3O5hMcRuC+ZUXFYlXI8eYL5/692TBki5xp
MB/8QsaogVpNI+mmw5e7C1y0xl+ab4BgOhjosYAeO6Rew8Frm/wdksceBdeySORK
pRcP3kFPiRd1P5Ey1Ym/VLVUgBBnY5BAqCQWa0gr1/4aqHgxuhaN4nor8bSFeZ++
qbFCqxwuS3M3WwSIJ6RMDMkMZDNIgmW/cKsMjj1c1gDtseNuW21NNZIofWFaJhKa
zwvuzZkszbXVZc1RwX7c+WxIVsldd4/YQmJMaNcIu9C5jg5/+3X5GeqyiJEtxxrt
eh+GLtWJZ2LD/Oq1mhoS3jg6vH6R3DVxtbVmxns8aOoWo9I2rS64pYvLvQeJKMpd
/ytbj+PeIk/pYZy3/4CsXh2vJecYLLlWgiR22fHemZCif8j+GXoSaIks2nLa9oMF
/RfxOGnftgC+NFGsWby09HQC1rDlZ37kIfIQ4Cg4OqfKyTRstVcjv02KGjgazt7y
xa3x+1Y+zMiEjLGPZazCN/5hnWEbRiYbE2fk/Jzcn5rLJdGbyS287fJgg7/0ICCa
S2pwMxK/TRsZYgngmOmQJfarh0/RLTmH287TDylt3+rwWqoaw8X1PTTCHjzAxGDq
Bc3yPvC2ipwLudIqjfI1CYPf+tkvOi8+Z/+9furOc6s5/hS35T2OnvhxDTvL+5OC
ywl1FegB3wYnuAxLH+GCVLuoZlsoh18VcfdUC0lpu9WC3IgW2dSGHhzyGTgDApgg
61SqGNqahN/5FULRsc5qqAwL4uus4plZe7tMznuVvnYzVEhkg/uvIKPeJTNV5CVA
KAVUYbkW6oe7OzPXlrPmrBQ70TrkMf0RBT2JgA81yiFydqnje0fn1cuIaUYa2ehH
tDKgoV/LsqA9R0iowB/RglPhR4L3J+FWcXc/80K3vL4VdQzB5yn3UorKXhADo8xX
E4DF+COGIFgDA/+SlvPzWi7KPUesFHT9f83R3FLdb8Euz7TVvJg7/j3+k1bt+PPp
T/FXKaCNH4S8MjAviGGC33cpSI0SN5ZseSwK0q9uagwruEGHcX4QzLrGAdEg7GNa
j4ZFUqNCGkNHXcJRbYevbavj+MjsPAKJi4bpZZbTkArjgNeI/o4kdQFp72vXmspL
xEU1CIOEWC9xhSILGrdCBx8zm9ifL/epB+j2I28E1tGHKXxOMwU+3C9S5B38QG7R
ZMWB8y7yE+3wRiaiVt4brHT1iUpdZSzeo+vXA9RNFX0W+Id/j+AyxsABp/vGcd2m
6jF7DTfiih4OB7I6930zLdL459PfAhvo72+jUDuF//ZMMqHuBCkac7csQtW17pVL
zrSLfkgz9fTxbUzeGw3Zb26IvE/WhOuCbFNEao5YB36LSz7foC9+BCbrH9DaxUBn
empJ6udD0vPNqfdyggsvP48FLUMzLT81bVSAjFNnBSkVMuj/KmrootsHeePqlHIb
/g3ASGoYs/ti9XflUxmyiFvmlAmVtmdi9hr4NTugJUoLeYIORkRptoQgQXS60lAI
2zM5/DN59R8oS6ybTgoNymXRTxctbj3p43mSzEyze2JEV4iXL9yWkNeL/p8TRLlB
hY5elFt94BO3gIarWV3FByTEhj9KmZX4QbJXsFLBLpz1JosfCuTcbwyQDegG2hTZ
iX1UzCT5d/5nZ3gbs8FS36qO44JBtYze+N2tuWQKl70dVEHahS0ruoGKUpNT2elV
0NALHtYp/oPCajI2WQQbw/7Dst01VJSILISJkwBtilS/Vi6lSQasHn+bjjT+nyy1
9anbQUjRJXTVNyJdNd3rWvIhsS2g+19G6M5COpO+DKsXW182S3Q1l7/fz4fO6q9x
lm1XxvfP41l2tnaXg7hj2r6OGjADD/Js3T+zeSdSy+g8vuNQC64Jkmo6XT7xbe3v
C8S72sPfRz5S4POW9fiMECT6pg+DTA1eTq/FaoXWgPbLyuxP72Gp/nCDIhG87yuj
ZMaPR4BKaEfuNIlxYayfgwsKWfKv5gmJNypLga+3d8IAFgjwoLG1/iKEFxpykIRw
0XG6MMPYd2XUfzGWJESQ6fDRNYaMJ5oY5T+T8U7dJgtKk1ew5VzJZzOylxv/eQRA
kvIdYVqrtjFDGiNwgW/QsyeAeLpeTKwiBuIN5L3JxL84gMlJTRjsLAbqpsKwhod5
MJQqtS7LSkIQ0vu4NB90rOXDwR3nQ0B690tGdgBu0BhJMs3kQlt2W26wdQhngFrL
DqlX/tIp2CnrThNKuMd4DvF6TJzxVI4aeI/9CqHphjQkyR/VnqgpBipeBchASnQ2
6pbe7ursR16gCOb6TIWwAqSeA2I/IMx72BTSzrOUBwjERH1ZSFpQO4T8o+LTv7q1
atMH+Tyd7/huA915EEkobhSNdMHL1pX/HrYx5xusRYPxtJ8ZwJFEDNi73EaFnviW
lK72N1hvf/2Ge2cAQVJEE+hHI5gjw+qlA27OTMDt0MDH/O/HtlReHx+rHsxanU+B
w0QGScuwUbNNniuwcswk+o9NWNDH6kPGWd028fSAurhlbgxUELB+mNp36lr7G9SB
yzPgWTvVLuJKqzQrTxOx7CkeHoz3KWG90sB1pDLMvfs3e8jIfHfniBFHnuwafymM
IQWzxONwL2zga3aQ88H5TJ/7jJ63O9PZYzD30+uSW24DfkVulRgv3ujf1T31YeXx
yVBqamctlX+mvfY2ZUblV375ar0w4sdbKi/QPG0/mgAJCUG7N/K4liVhvpxSz6Eh
wn51x9AeqSV/V1UqqpdvaXIf1ZYOT1vf4JZ8wnkizFGR/ddflhCuUjeVYsw4hK9A
nz8M3fwxFkMLTjhuOwov1rKC6DzeD77S6YIZW3yJ+TsI0z4s2pP55bmzBd/yTKzr
r8blNr4EpA8X/hBO3bxsdZMSXA6brWCfRWNwfayfCUaFMEbZzEjZpKdNt9YYE4xg
XdrGiPq3EAkrac013fEM4q4XxUGd8N/2NhiUePQkA3+PjmrrfPYHBBOLLxaq49al
xUOnng6N30ObKq5MGX2GpxMQhH0zV80c5+ImBm2bUg874ygY/wl7bGU7wKaoPgAm
dbZYwzu7JmCmULEXBUUGBMYwU5iQs3j/xirEeT77AcguiGW+trks+w+dcSRzEMMO
Ou4UsyWGHps7yAVUnl0f4tCVEUSlaDzeBDcl6e+usrQpEMvzQgh4IR+Cfnd9kyJw
LrmC2FFrh43GkFosZC5d0zDjQWatML52lfZ8AzLrusjOWCqrKrRVsOonCe7BwWNq
opVkFABXBAyheLc1xKiN9ru+IPOKo4mkZwwfOv2qVG4tDQo4kHPPuXvs0ngQLCy9
Pdi0lBDDNSCCzjEquq5NXUQu/s6VT3Y6tw0wHBH8fe0DIHcBXp4aGI5UHrZU7v2w
2bdfHv3jOWLYxDO9yZxKDLIUogIvdrNIbN2aZA5wIzTOP724ERB1SHD/VqOP/L5r
bPtG4/lhL+AzMqAzxgASDmNb/YKyrY474CVC9j4j1cxOFlE/K2UO9xDHofL7Iz/C
SXb7deTn5Pmqi7npgyQB1rcEunslw8dM7VCmxtJW3bMtC7Hb9xuousim1qFNYFmC
75UA7ZrCAHj4G1xgLley2mLIidIeexsiN2pT77/f34E/QlE+0q9QLUf8ahIqAAAN
a+ox17Pqz5PfhGpuY40wUc1hqBD2vjyvQYsC7xQvKPr9sQeWeLvDi0TqFAnEG0ZW
FNzKH7dsYRJyGndwCvGIjFf2KNKZEN6V/82/2PG1Y6V/xoSkr9aiK0mhTCYChTK2
Xfg/nUA8kScv3+jFQyQjW1+PTZm63vsWhF9nTN4PXmTGuoHfJuF17MTTu0gdrUIr
1Nhu8xB5/apuq8s/T5QBiJ5L2FZOEg4DcBx/5YcuMGIRxiqaaPfnwpa6ryO5fcFv
qSLotFf27TEo0xSCXzou8rBu1gh+xLNnRaCCbZx6orZA6BFZ91IP+t4uZqpLlGlc
sJ6/R2DFvg8jEu1o4TrvvEzahD7/HCg3UeuAJKwn+WyszrKQOp2UZOUJJQ9kzGdG
5G6sBJVyP3F6yYfSBUCVxHS7L+1SY9W9FqNQJ/fwkLHdk4gqRbYONCsf+szFuLqs
LB5ABQ1kUeMh+XASVBWBv9d4hPOaiDgwkq1p3Z9Wha5J+cP8AznqyHh4/tPIk55e
am3C44AQCakgFGuBdVP9r5csFoLO7Ef08r3hI1+KwSsURf6P9PEMFQgzp2WZigDb
4vWSPuLngoMnx04TaHT4UHco6oiTiVO+ZTyG+2SM2ZZJkNS0XKADuQBV8P3AOvLm
p59RoXFqDNyThfRHNHC3lZdEnxxwTuNVDgpZmDnoe/8zy/yUwuFnAGDv0m1Xu1jR
t3RGhEQIBtOX+jMysEpdWoIoeDK84TScmE/4IZfvHLCWx6ribRQ8nIkIF4XVbKyd
77iuwV1z3wX0KVzs8LqVc4R83wZXjLjY9wAo+0Gwj3Os9BVx4rcOEFE3cUmEm/Mo
q4f3d/BZyzc/nQUMsF9HYfRygcZHuvaUq2HPnIsP/QFcAwX2+usi9MsJzQOOyxtp
SDhPET7BmF0TfGKB2STL2cFnwr1YmrtehxWz64y3g1dsPNh634OzCfZGg++bOlRd
ZU/+fbxNuooPeDYQ/iVw2TuCENe+rWG7K2yn2Qqfn6xyDVeqjN1SDul04s3W8Ev+
xYRKYnnIKwyTBi/mOX4kUGAcyzJe/VZdsc7I2Ms/D2TnQd8sGaNCLxeZ9i1Z6KEs
1TYptA6fReuyPZwlNQNl6Xr0ymTZNvz5HmpYU3FuId0nutDbC6FnCDVF/TCekbue
5osFGfeTwliBM4Y6EZitH/qGC8OhB7Z7P/exc3Nq6Rsi9Te3cyXHh8sDQ97Nh0kt
JMGlrWm9J+86JEcMgt3fem/8Udg1H8FUtEV85yTABYJuj2+vryH/kJYiUb+dspR/
w/GacilkhRiRmdj4GS9Ijy6oAl5RQYCBDpXUuYxvwW2TjLH/rT3qXy8luey14hk7
ZwQbbWm0FCoX1TxKmmgujUsG842Bn6+40KCEvC/8OydiTwoVeA4lLYcWL1NJwcil
d+NZJk7CebUgtwpN9mxVHl9QBlWDc8ocath6cdOjThIxR0sR9B+2aYgWH4edk93V
JTfZ/LSvpYqV8InVVaJijWiKcgtXuwEcQ+W5qGWAFwgTSlGrFwFAdpUsO5A96jvn
cQrOKCRTJvZZYbQgXkgQ/l3NU/t/PBHJfaB/Bh2TbAHos7MEmY1bHD8xNSkF7IfA
eD27r71edmUdxmo6GxctXGfOOjOvdcaRBgsv++7a9fOe31ZDxWpQbLnUCnpL8Eq2
hfjBskB+dettsdvC+GxkzP8fKtHY8ePMGucAw0JlDYBX0/4fKz8saattySgijDDo
ymC7VCyerlSLfEH++nzhDr1W0HyWNkVLdiMhxE/tSb1bLCbjqjRAE4j+j5mpm4ss
2Ks+VgtYIjXpkYk8kEsGONbQTL+ZlQoM4eCSRVGPSo4I2dFlIIiYRIVOqimVJG8O
K0eCFkyXOVeWAt66BpYD2E0hYzXStW/8LkWp1SFrZiThYxXjs0iK3KHwZjEr0M6H
5kWQX3/Pnpk3Go8yjCFWFcSRLz6NdNjRCy5XidmZnFjCvkKbcos9CCmvoCRWXJsC
AHLsXzAIeWQb0YSCfWIttVd9FTjZqGRyUz2moKDLzHg7ssY9plOKX+aT5tlpoOz4
QmPjbwWSVCGd2UrY0Wp21MBb3xLC10NQa+rO5/xMpKAjXmENqNOi/aJxf8BCg6KW
LQgnYkdpb78cuc9NrSauc8eaDfq6q8Q45YQpjPmJUVyHZb1hYsre0FFSOBFdBXSz
hemZHSx6VtQttq+fE2UEM7jDkceN64+KGQoAVWZfDKJPejow7Dg3cGptBsBkMgMY
KNdsFME6drXSWC1/MbkALqT83ov8YKRwQwQzW6jg/KrdLGnx1DZQ5kp9pgp+9Q6n
WntJaqMWypp9ZTquAGysBBhAgZEnNBmnSF75zJ4VRETsiU9j7iNacRLhNAt0gE/p
WBUCC4TJnTI5zqS3zIbdg1kD8wdAFIWun/UlmHBoxLR1Z23L74Yf0MtjtpYgYBdR
gjVvrl5Ujwgtff73opkQkXIepJoBTCEny+v8XF5N1BLgNbVbSJGBXamCt1nSUKGw
omvTs/YB8BYfQjV6Naz6tfVmovDwXht5uJUjWY8DE4C0iMd6E6uKZLcs7ksBmc/O
SrwNaWPbEwlo/h38SDwRogReJDPfgcLkwRg9zZOpvUPGbdQddbG6+0wAilbsIdjd
SmspjFzit5vvGKZJ1z9wn0VbETE7Sf7wqcI7g9t2A2JXkEnp48+mQU2J+Y1E5YFK
OmuoNzxwz44kbHY02WwbVqN8PIyKk8LpFa8+ISP5tTP54a3irgYLts15JdnKcYnt
4wIQzyW8CvQvYshsG5msACJJESzuylpFUIgox17rdu4VgzN6oB3zZhy8ALCBojK2
Wqo6407dTO2S8Fc7F4lb6Vutv0Rz5/+HE6qBT9237sqpkzLaqfDemQ3q4NMEYmAi
ZHqdAUACPSZrtH1+TK3NPCmVJbrSpL5iqqxitq+bmGXCzBs3UvyBtNyvvJAo0DqY
UJb6Z+K/pEd7pDVIuK9Vn9+NY7aNw4CnUeFiEWqzyAZbgUul02Jo5w4kdG0FkS59
zw8aLSWrtK2R5gZBT2WUpfIwHk9wWEGDnABvWr+yQEAIefnpZ5rDCxoBxc2zsUJm
TfeHyvsEQS9OGMQIzEHYt2Q9mK87i7NM7ZW4LR01dXq5rTn4ov5pGXaRSFNQG1tu
ZlynZyR5XexxmZV/hbOFYDJ6DaJIqeRh8QjOzc2U+pNuvGyVsC9y/fdk2czUZVr8
ycdR/qrSNYpYDswZI+kK/0tYZkbxWMa9wCTfpUSlMcmOQAAMKYUDb4Ctn+2ltG7f
UrHAd4P1kJ5VFmC+e2YZ3Norpno2q3S5RmnoAb9ZDtJTSwlWSwTpIFdbbwfxhnhl
kU8tXU1WcvGdMsr93J9wWK/DP5TfL8psgAjpMr6oUGVt7Bu5qzhEA9PwNu5xYHpV
1jqt0kQ2yZ392FxzrvWEoUwfrClje7NSkIl5wXJMX6CMaXjoyhekdLupSAYj1pO0
Mwz+5x7R9bXsIdw7bZIAlUIlms1TGdjcgs2hX4KHCudRi5Y+M3WSPh0+2PfYnAwx
RwmWXpfgRtOF3NtnXufw1Y/FuWSXTwkcHtVtgoTpRlkNxl3M2rKY/uASeX6huKBG
L0PvYJbaE5inOlwZ808QLBBY0qGOPcKylO81TXt3gM0gwQ9ickDqZSpFH2IPU5lV
pKchE+w3qITcXg2WJ2hqRhgfGYJRVkwfrzWnqU2qcLSeYsllnBf/AqpReflC6SuD
rtuaUaaks7A6I1r1UM0jZkt7LGrVod7D98Oy79jhtRgXpizwBApend2dRzdHjFGN
Q0KrDx6l6yvnmUCVO5u1jJlTbIZZYhxaw1HJ7gQ1HeKPe0XCWdRzU01Ck5hhd+P3
4o9RTFK5CI9m6MoFh2rjzh+Eu7IyqB6AesHq1l5LOpvLTtC1Ls45P6MfHMyqmqda
xE9bVDX3CD1WxtjVnoMwOKT07c5g9fz1Rm+tCvun6lxi1ZSIr1MY5xx631YUjwEa
4je5CSuJqLGVpIeYwoNdfCf/Uzlj5Nwj68qiSNs/aVz4sJd9msjtAU1zSRHrPi+q
zzhmjj68Ujy4zeTfxI1UX53Cg2ujnakiKmeZFhNd883IL4WbvlTbhaQlrocUnAKm
vBtmOvKroUlli/fR3vkIv52D+SWqIZyVEvwBZz6amluP1j3TWmC+dm3fgB+fK/CW
eza2nejb3u/hLL3D2Go4HAgR0vbxqXUrvZWeQlisk41PrFFagriLSt74g5poSeH3
36dWuxjmOdyF2gDui1WJHs+Pxtu+CsFmAH30p4POviY5wFD3613VlmhTssTt5f3F
7iCurnhZ8nSBoppD9gYCx9T/pp0HKpq3eAJ2wLnTv9WamBUva6CubkxJgRP6xtP2
tJRkLLScz+MSPLCXYsfcOQjXHT9O4UxdU3NEKUpJEVIWEDL0T7f4jFgRhosnDl6y
QZsjigca+1Me900IS933b7aYqwNqgETnNH0sNdgLpm4vR1HLyN2wII4LRMXMJ23L
uQCV69ifWhSQebndEHU9Kf57y9jxXPIcTX/zb+cgf64jXbyqNVMSD+VRUx+DYxr0
TctqcujM5/ZwS0OsW5EZ0deHi0K/BgT6mLNeAigB7YSDYgbLueBq8E4NNN+RC2kE
rIWu66uUuSmFqS6xWI/8cfqVRAbE8mr+mEBdBXdgIu0oKrT3v4CfIi+KlvSmRNl/
nKDeyAuSshQGWTpPEOJyLdYa3iOMNk/LcCWXaCZTvum61hOj7RDBSDe0YmrFYLSA
x+chabZ28LaglfolaFszCAIx6w42i7TTzSY0LvbcBFm9D6WlaNGtIgaZ9OQy4uw+
ptDjP6eX9Wmwfx7Z/sQDWXiUcQW7PV59kcXoHpzC7IfB7aRpIPd/mUCpGQmB9BRp
ESiM/sLg8g/tVR9d1mJQIrWdFI4R0Ff/uwrtGsdvMhK6Z6xMYP2HBgH40WTgpBOq
Jmll98ow6FyQfe+7MmnXXF0umPvHS63bUP6ezmC3wStNlRfzLKWjwGKSMqd2L+k1
voTVo9MFvRKjf4huYTs8tUNEIYOSL9UboMM6e1n7ES5C+6edNPx6xPqsVUMVUK06
g1bPfKELWkxktiyMM5Sr+xd964HA3XtYRoMTN8YRr5vqh3SZC9K834+fyv6qYdPx
DQcTEBlarb0zQO2jpXgZltqGyBm3VD/c2twAz9h8Q+91cz/VsI8MznViDsiV4Kr0
Z7cSDAXGZtd9Wr59JBWfu7p5jahSNoxBsLpEeOkPA+7KeJL+y8yqevG7af55MYfN
jCYIelDDMLuOEi1dNaTrFSYLt4nZLCRBDwQwpUgJw2y7RZNSQmiiSp8TKtzFgShs
wc/H09miUpowVn17NB7o4J5COGhQbO+Qf8lAFjkqN7Eq30LbguW2Qf74gwaQHydz
+XJn/mdAqd9v9VJoZ9Irr1znE9jPElUhQfRJIBVE2hFyBmlw9XjPE8rLgjUbH3Hg
V4x5xCs53aR+i2gWoK6stFD9QSl6ETu5BnjfRoZgr21sKHyF/9zUBE+cr1cKKCNk
tmlk/Mtt/UI+wH46xFJbnc2K/vbrqa4fp9SBu+o5l8FZMHgghZv7EpVLEGXOvMvO
M3/gZRfRvQNR+zmKlky0Tt/3bufiBwimNgBQknqPqx4pPhl84cihCJW2RbzaRbfZ
Da6Xo+5B6CxrJkPPIudIyko8OLmzlkTsyyEhPNZFrv37Rm71vrkXme3/Hhcu0a/T
LJZcOPQx22+nq8wenq1cV83mKgn9Fpi21VdpTAKoYHguvDJfQA/854ZpDA+6+uyU
4VGARgIIcoiwrGDKwlIRsBcM9xm01o6ZAuwMrNUqGrhN9cef1Q4N5LmhgCnRxIIZ
xJwcr23TQg6yS0bhIrMPTHWw6vru6qcNbwbe38mdlwn0Mw6MgQHSE7fLNXsJ25fs
CNuW8w/BTg7L6B+T7XGhDiVdIYHoMB8GagDe09B4F/64Ai0sXAZCF4Nvz7ronO4z
2+J6VBSKjdvX0KRGoz6qpcaAS9/OgBM+/KUnmP7SRaw6c1OMDOF+2yI9ztl2RyaB
yhjPDzpUBExPz5NSsPjcaxST7BXi2gQWQkNvWYpJ6i2XALU4zwqLaJUEvkZ+bqO8
cvUYpCD282+/ENc3PubbI9QKztuFeNnTuqHl1JwLrYODfBAYu2qV+mjbeO3s01Kc
YA8E2BCWT+xuuVRMrZeuQ3n4BH8gmmSMtW/5KOf99akngU3v62cIKiOBKWVt61ki
AQF/JSTNgV6LArVKza3DIsKayeOJOWt4rR1euUgpSqoyI6wYqd9L1TJUncyFD86G
hHKzgQSU4LCoj0XLISM2SborKiadYSCiL9bN1qnlcTCoPqumzw5p26g3SuqV9UzB
Jklx3rBAY5SIQF5jBeEOFLSclTi/H2Psa/ZJLyHolhY5/H+PxkD/MgJpfcXr4EuP
AgrDK86d+uvNCll+Dxrua1RPE5GF3omriWIFFu0MXMSosJeblC7fq+brlxZoiRxy
DwjxF0a6MzYi6MKCeW8/z3ZT1jAWHSZWKYbZk7SoRg9Ltyjq2VdLiHkDAp2X7u3y
Kzy6jc3TyV95wBklGmLdfzCxm6lRGzEwcjWojXmjGZ0WePEccA8MiwXqfw3b6FlN
kNPBcFgWOHiJij4sKK/EwnQMPh8P60Ov6TXMZELozrFG+6dgmHlOnJ2wKl7120+Z
h8/mIitTpML3ta3df+tZ4+Z4gapwSzmCgNYZWA6PMIu2tU3OVBQK+MGcAHGKqR/K
zXOtFjn7316WTCJI3HonIKN8ScsaswSZfq3tPVLGb6g1KcktkhTWt3vTTGSO73As
ceCtite69nXmlM2YySKHUW5/AIIJ8hIGV6+wQPO0Ke64KjANYdY0DNV1+40NYPA8
aSutWeqtZhT1s86rAFKnFWib3YbgmMvVGvI3THVpZVGlmK/XRVkxDmFxFKOUdjFM
/pZa+cmtWLxtBMntKkYo+Q6pOFjY7EHiuWlSPLw8qmVGRb0N2jq6s9fIQUBfbXNO
abjjkKNjj9XUu6lsc/o5SNVG5qLHrP7R5WsBGDvSb/i+p1DLq6Zo2GLrlU1mQlvZ
3MxUh/253eE7EL2CTRaMrg6NI0P1NTIRoOfMtF2/0zhEqdJ/obFznzWqW48jz5OX
FQPoVYwCMbM8KOZkSPQKRaf3h0rSkBtu7Zyz5Lk3HybAx9dOWDXD+dc8ufAj73J0
K7JBVd7HuWnpiS6nq22MlDeuyn9HmVtUTXSncyopuKwj7bWJ5NgrN9ydA513jGnH
rlF5UqWqyziGgdKFOFXhX6pYM8LU10UUhpARKhZcyxedtUxDp3h1VejALOLFOIgx
nQrn6++qD/oI5hVAUW3nvcZZUKF+xKsQeOPeHBPIX4RUdGKXf9jMZyCVPmXKuRIx
05E0S61Tsvi404Y+2jJM4OFJaipdavPAG/E4xniyEbMdlDWYvmzOokLfaiAVCiCE
NC6Z0h8YmiJJ34MwlzhWWsjmspVoJJMNXaE/6feuocsqOZmUsyBrg3prJGY+c0JB
9AzepnmS9R15Q2PZxcfvNV9MYETJbEoRv35W+AgEnPp7FRv9rjSkxmHKSWIBy2Ij
xSIBKUNoOvc2SbSJu+wdifz2MgOttOADXNGW60IzhG8M7d2XaJejmkEsRNWILAC3
ipoekTD/v5uhjpt+KZl/kGixPKp5BUyIOX0nyGiC2dYFM2qqDClBI9/hCYupBOh4
aZsPhVrrme5ACveFv4KZ0zsZ0vpvBqkMPjXS09kJFVJyUDAQ7AORAI4Tu3IIv59d
ZD5w/06Uly2XaNM1DF68PB4anpNjfP12fZa0JzwkI8a3Ot4thHUTdG7Auf9oEpka
5hdhkptst3NOPQ7TGm2dlOaPlMIrwNVth63Ret+dfjcEfjH32gq6fy+1l/coVgiD
yZpph4uAAsdXELKSSEMSpviaZMAFeb8/z7COjQUyU0kNpsItxdxx0+ABKafBansD
+ytmWji5rG4MMRjQOjBOtGfaSMkD1FlXNBHZhDqpZZTixlNzt+dG3If/GTEConpd
VQbJosXzWMS3t74F1Z3LL39gtT2/7pQ1zWnglc8Ed+saA1JEvnEi++ec8yF2Gvi4
S79fdnyeP7ge/iV3hsYfKudH7N5QhIZYYmq1pxQsuGDZ/rYFvUYUd31wS4DLnDuQ
liif1l0JdsOz2m0eMWiGkN7NsIPCjMM2FzpRKuciQI8m0aswSoQ7DKxX01DrF3cc
1QpLMuCRWXM+m0YC6CILYKbOqiJD1m/CwGqz2C2eP2PbT5ewAM3GbEINQAtTGf1r
atSPrajnrOnzVQFKsQlu9+i5THTHOjbhGLY6EENENYJmTEXYqn4YTaL+yHy+NjVv
8GMW7sl/9ZdBCuIcVFCjfTXRwwOEk0zpYmNAqNzgGmphZ4LmauJjBE9Ny0xTJFt/
j0WolqHgdcm+EWOqOgqNrTrqNybBFyPGL1EiiXNeTS6LagSfjpkDoSIvBPKFQooM
5ntgJi+nkkzLxoj+0FQL335D87XOzEjryWBXcEwVhYWEM5EqiYHC3P0oiyLsifsx
uQ2pVp9WGMN4c4SdzuJPY40ZMJzg3uuCSLF+8utwxHkqk5WRMSzep5Fm8ZCvKO6p
UCh+caxAjZgwMpIYPvWZdPXQ4laUYvdlkLOEXzpS4Uxz3qCYYjPsqMEJBU+vQpKR
4sdP6k4XYPGJO3lX7W5KQBDnZqt29jhiHLKDzV0OaMm4JT4tsMsXuVfKgjrzwXT8
E0AdY/bbgsgAym2Veod3/Y657EuQLUnPxhh5qb/pnHmUwrZ3wUy86mud29sejrBC
1CRfft8rRZwRkvXQy2s/27HGhoEFelLaTORvf1zo1djx0E+VdvWKkjjHjxRLXGvH
ilrFjE6kHwoTYFy/i4FNQmyb0UsCyszdb0Z5VGWKSk4NiCBt5Igzxt513FBwglpT
eO41dCbOxj24tzmnsGqoUg4fKVAqnZseZuapGG6hKsRu/OhQk/hmY5aGdSI/5EuD
6ArRSE4hln2Zsxf1O2si7H0rYZvoW2N86IAxIY6NMOKkmSq0vMm/HKcuzUob2t9Y
3zZa+rhKNJPBQUAZXXmztRtPOzck0jG2asBedmdTNQrReWHKqlsE9Gq1vLctyRZz
Cr9+HxCFpcsMedQY4haY1cVI0u6annpo0EZpIyDCx7Bh8bj3WYpyi1PYG0tu+pd8
Hi6cfpPqEVVPI8TzkziczS64vg0Z/ts/PSpWkg/3JHOHl3dhLboaoFJFgXVb9K3U
HOvMhmmaAontnn1a4Lvdyc/TTjWnSYX9d+Sww3RRlGhh/a8+a4dyz2mthYPCpbBm
iMf2vRVCPWRfKMQDMhozfRwycTGLQbvw2PijO9w9gk7/hc6GIeJ85C+pLPPQ9lV+
Xzy2G933E8zFQbV2LqbFgdgGhu1xO0HGWFmYG91V4/8LW94TRydV/T4xmYqjVuRw
M3TwZod2nqiJtdeP/LkODD85YW+lMfGriI3sESL9x4F3LSlzCu4XH5JzvCaqNt9D
dzvAoSLKMM43ajYo5TYYGfLK+0R1FGYvZ7jx14rQoBJ2EYbPtvEhqqsM21HV1Xxx
lG4a5Us3mSANGgUAqiY1una2Y/L30KgJyduCcy43YwXcDG4Tf128J5sA62eY/0i7
sCBxnT3ogwGHNkftiKyZSdhetSjypfZzGatVJsLK3tVnkA6bf4QCF/lWGcp6jcg1
B+Ee6+AqeF6XOKfKcZDZR0lBxZtqldXC8umciLO5hq7y6k0XPh4euJoo5vBF4GEM
Ji/koD8unHU9hdpiS3b67rn0EhBfilndnGW3hJH4czWemFUYmaywRLRh4OVqRC7T
CwOXQgUK5HH4p9yNJfjIN9H2nVGEnkx67bvGTiR7jK9Dmp+cmbmCmG3t5/boftVE
30U6b6K5sgQgii4K4xQb/8nAUCr1IjVJxYeFFTlZlTq2aO/MFOVzAOgogY1R1yAZ
3gvzgx1Uoz4d3bSdIBs7nZFLb+KrELo+54ohzR9caCv9Xmr2intpYhOFuxE3BT/1
vXiyuIO3Ppdu3CHw/08x1nuJtRo8TSketqjQADULojK5JrL5F5A3z5kKu/PSshKt
dedobxluGoJRkVwo95lLu5rb8YKZCLSH1MFtKyBq6A0BkEA2O3gX+AopkaK9Z2oj
27DMmGkl223rWluNce2GOpI1spLp8El3wFT+3ReSdigKy8YoLkMcKiAlR8zBmbFt
+mfV2qrp6DaiwyX3KVs96uodIAXvwRFJr61Ho7dquaByjrOmjCEgxF4RzAFr4/no
v6JZKIBOqzd8SuK0QarwNvlc0Ooj/OFJ/D6frCnrl3CSkhw+Sk5gSMg5rtr44uSm
bj6QN7ObprETnXLTj6EtEX3V7vI+0vD7QxG5PEKuOcj81lx7ZmaDSlwhbwBHMKMU
0wTD0VqLc7oF53hVqRl6XeVOVEjMZ55XOkjpgaKr62ps3jvBXyET/yWl+GpTTvyf
zpBDlW38HT5lAxBtK5QyOZWFXLySL24rfW9z70nkr+uBuFelejCoWRW3IKnOKcnv
ayH4b2FYDz0gJkPlVVvVvBaRwpQM0BCyzisfBGmWSZ/FJlO7NXZ1OZj4lr3mZf3C
QTCL0RLh2q/D+fY26XF1Lyvk2UytvMOAX4YH/3tCUgTBabExPhOpmv9qEJEmSBOv
52P/JHnrqEICYuE7bzxRCGjHwFKbM87qzmRtF0B2ekqY5GN3rUzwIUDmLW0lTCmZ
S6QYuaMfxHOueVQeBWDcFeaKJT2ajrorDhqffNqD4x3wHeZk1hwc1v55FHCu5h1l
mLWsCaCIb1A9rDJm1kCc3G7+GMquz5ODK4FBQpalUHp1qC46DzbEaFxa+xR6bv3O
/QoW9V0V4/ZzdAuEYZL5tIJiaUD9SGQFdNblERvM0PDcRoVOEttSlo0JfCP4M9tK
17UI3VOckfwvoQ0pjCnY+cW7y9dVb6Zh61W3nme3g6nmjGdd3UTnWdo6TjdrfmqJ
DqhhNBk5cj28z636J6/WxAxvch5DJXygEUp892mcNwAnBFo33pfovqnEXFilmBpm
UbMpXweEI1jiV+HbWv6xiTnj4AP2AQkDKvwrFzmHmfUAfEhoQZ0CqWbeB1cZTeAq
5WeNM2Y4szHexxQH6xLuxBcf84oOAifVB19cKph+7bMWJIfRcdlemPEg9S+7R6/Z
ruuKb+3pKJVsQr4DO/utfxYLhMD65mp0pIxuK00ylI7DnF0rTfcnGiSmDXCS7n+Q
GVRTY3JGjOCq1TH3enWP/kB6Jf22q66nG0eki1+/7UsYe420B4aqDNsUnHr9KZsL
FCLvvC7Qm4lMHT39ajq7CbWtsLBpS1G15MepIwfN8DDh3fY1vsfgX5xtPxLNk+6g
lSPmyeY1UNtfFC5FqfQrXw8gcmapJ7/x7i+xsbWm345CO2zpZTX4MhUsIsHdLPcC
MhwksZmT9jRFfZ/4y0+kgyUmtjiWxNKdTHRCCmi2wIQhUk3vyvNOXR17O4f8evl5
SxcVf37b8LGWjjASGb/h7EdeNA8AkAVUJlqolbnouw5K6aspxZlcBkz+NQz6oR/A
j5H2COGlD2jaIjyLPlp0WWUka1YaJWS79dbUYhxry9zum5S5Yil9MONgYYBPP9/t
vLCmYsMVndSZsHwQ8igNg78JTaO2QiwhpmoCNc0GKmDNSzVi2xajgV0VfnuzvsFC
BzA5Q50U+me2w4CNW2hpmnQMMIsoFdiQi40NoFQtZron165dCa06OXxE/Kl+XXq+
T5/eZbzSDWQcYaDEjUYr9w6AUTZnMjpBpkQNGYRGthjXRhSD5ju/4UfVX9forwf2
soFlVvpLEm+8hQU9xQx8FnmooSlc/4IGogStApI0KAaioNH5Aj3lm8epTZOh4TpS
Q1fs/qGNx2nhp4M1wgda6Z3Dyqyt0ZjgVUkyQ7ehWikOFMVSaIpXlMqmPlT3u2Du
WnpMJhGKbYNk6N3uVR13wSMj42qN0kMrNitL8PkYcYQv9eH4U28Uf1dnN6qk0bEv
mBWsi1C/SJr6p0iGNu5onPkhC9O+j7zsJM20yPYu9HcDUw+T66pNjQlWiWjkV8YG
aBUfk5wcV1M67WdTtPmO1io3FUo80zQmu3Bwr5mUsRzZhiWAj//D4fj4/E59Qmxz
UqsW/8RFaJkNuzXvvftFMQneT6sMgW2Miz09SjvygbYbO/ENzB6ohfrTk/soZ/04
rm4gil/4P+xDm2sqp3rVrVO7bp8b6MOXOBcwLYY6JA9+HmDrmUr1k7dVlMWNuvR3
APxzk2CmedI0VlG/x9mh7awbM/vpMbnxy4sjl3UN8d+l2znHo0+t2018h49qqplG
6qMJqLtPRy/IPvwHD1ZucykfsN6Gsl6EtEs4+glkvyZxhyhLaLv++DFO1ftoNt2i
WIoXGoM1M2XG775kbPh/RslVYt1np4Y7nDtyVdEISklxxHf7jeEsYbytSpouzerw
p8LKJ29mxeXN+Xe3iKgWlRAR3nKbrr5jdVyzCeflTpFm0AhvHAPVeMAC4J8EKrnk
DDtRG780yMI4IfH4qJhsrhQUlqV0BivzfklL0XSMMLvx0y6Ppug1a4U7Mixueah3
6neOuQecOjDMyY/BoPDeOP/ukpSNloc4oLzfNykTh+uqsDrE+Z8F1qIRa88YmsUw
1x2aXdcBnhDQVhP1eL2VNAT3R+y7rfVwsiDDqDP4YVxon/5X+izfs7eiRLY8n5MA
k28JLcEczrGmmEfoG0nXrAyRROevpO9egCbJIUr3/93te1E0K9RHadD26HMkfPdP
EFbliLehTxai14EArthl1mTAyFfWACaL3ScxBSb1HNg0jkORDRFgX6w7Ylq3tr4l
KWK2+tA2ylIZolkudRoz92cUZnJJ1UBWn3q/E0EA5RdTZXITWyogbB2rWKfRB4zF
WpyUFhuuMf8/grRYzmRaDrM+cuppDM4XtwZ65RCdiVZCoSbr+vl2H9q0G11/n2TH
GGP/lTd2FGXuLi5tYyB4iQkFmj5S4SkCqt3GERew/FIuOmGhFt8IXyuHd0O1lylH
HUe5WplJF8ujbasIIpNpyadOmG/SCs96HHm6t1gxtYFBfNTxfR/Z9KBHntmusKvL
Yhnc9iXKlD0qoTVrqqAZloA8iJuYU8yZoiXzJxlCUgxWpXAkq75wnF1kUtHYawJE
xv6roAuiXE42sn+aJr4Wy0ZDnGjZP2jnaA8FpDOaAgMUbJ9dJfb64Op8McnNUuLW
A+urXq48fz6q7CXLuHuVre8h2AtECdWdChxbVcseTH18EDvAuqAqsyrbXpBuO8/d
Lu2Kx9WMxPQ4eQ5imNMVL14uAm8iNRnE5dBPhnBBGcQzOr64r+CuJqC3dVUUjqB2
B3scPTrRIRc8Xu2mtVspRVjL6OWITn0oEGVOe2GbjU2+nMhBMNMrH1lXlhvS4aKs
9PNektr3wFAm3hPbzqLs6byHav9G9uWQ810fbVok3UsOTRx1Nzq8Bi0U0bbZmuA0
o3/ozQqXGUX+s5EcAAkpqTarwIH4CjRpZZSkS+VP1YMvDIQPhXQNXbpwgpp5kF6x
sMAQl+U3eigqbQuZ9yfV0ibG2xvnjSgBqaOmm6iDRg/55ZejB+LTUg4X+SPs3ynh
o2U5wa1OyIEZcE4FcSXqh3EEh8KfCWNHfVDhElSEYtdMarx5sCuQNdREP6yU5gWi
zLvbkmQEngVER+0LyVZxhdou3N9hxGE56eNUQiKf2/yocIOx2L8wJw6sRyFmpwxu
CugYw0EHKIvufH4PtWuMm/80RdXqaSA6Y3gRzIy3k/u5kyC1VR2cCK+enoq2q4Wa
o26A0K03zdVkh7+05Of6byWs1+cZl2znqZeVcjMKf030rglowI5QQwlEK9pi1zhs
6e3/F2PH9bBMwbd6UAGq2NtgEVNKL1Tby9aorXZydUoujttIajQu8W50QafPizJB
dhfUoQmVB2Y4mdKX+xDIdjDNKM9lbYO+2rz+fWlgi5ReS2qZao/cXgFmacVXyg+p
hBiIyR83HD8Mrc1AmNSMEzYzZ58VaIvtOxX4N3U+eM/yEvlejXIb/ab66k2+JOaM
zhPJUnNDL81FRDopG5/QAXQCwLYNj2rVDGDPOBtu3J65nfW2C7YHvC4rvWkoq0oA
gGqt5DlZvxG6tl5QjrnwFGPlNrjfeJ6iKXaNdl5lI61g6hLbuA97oSlpFWZ+zpH3
YZBgj8jUkZD1zk54Ul80VKgJUf4UvnzP9zZm5Gp7k7PqyHFkT1dtDEiRdHfxlJeH
KKLhyBiBBDHWqoX3/bF3LSjfdSuxYvtUkeajw5wh/zOrnRqIVH52QSeVWMOhM0aD
VSMSlEBnM2QbBQKX1QqVK+b+J2as+XFlU0Rz3+Vd6w4CPzLuY2U71Bn7s8VXoJcl
psQbn4dFv5tW3VFNyOh43l5/HNkC11Yo1Ls6P29436rwIiU6xNi3tWZcbZKl64al
8oubcKMNaiH1xF68ARvQEiMZdeI2r1FnabaHxmAOvqtowNLTTekIQdLTH2I2+K57
v1LCVSrP6MrD5dbIsTUGQhgy5PQS3nH1fL5OD7fz6S5lbWsZ6CAAKEWbKxEYJ3qW
d9Qw8lCdlODALFAJSxOeJtxv11qxmRpMjC/dxcLd4IaiPNJr2PZIJQgY297qBZXy
0IyZ2GD/1bx1g1jCwUMC2rEKMoXkxVp9JOnB/vSPVG2BUOu+XNR1dCRbL1TzUREc
MOCWKe45eUYMIHdQH/YEXlgc9W3Fuw8Tthxzsg6auaVxNNwJdNB0qNxp/Hf9G5Pc
nGWeJxFdwYmvenIt3IqwITLw5DZly1t/ql/SINcgocAO8c2rtMpbR1XJB3LwM+pB
Fxs/Cp4GceiT9rSJExJRD35FmNvt7QiWPibI+Mv0jIBSAZ2/EpkNES/LvF3A6XuQ
8cMEJ212qPB8Y9LCzuirU2A9fhs2FusdhMcJnGPXjFFNPaUsSngg0c2SeSkCVZC3
A5taqUSAPH0IXASjkJeXHGtCxsuAvSxuVAzPO6SNPaSUa1Eamde9lDleeqkhBH+y
1ZoeQVp6nl5Farkqdgwi1AOA6RDuQbcIlCCqE5b9Ms8yu/KbXxby4pRyAfQNo2Qc
vqwCQwlNQUT7gq9e8U8MrSnFL2uSjY4032AnQKibT87VOyWqUNuaEhCIiD4L+du4
c5plWciM4+Lmvm1j41o9pGBMb/94yw+xP1gtzNUDZhzYpcxLsC9troeGg5IvgslO
MRA9PIZO5L9WdiJRE1IBNQ7tYGe9HHu3+KSfyouWRZJdXHJORH+ZDqgVLLEd5MbG
mE4ZgoCCUnEQzJrgKG2dQWxvDSrUImQokbmiNGOkRNuDT8YrSDx+39dC3lt2dO5O
6G05Z1plJyhyIHKjblB8pwJ+cel6+3+NZQBsOt2D7DkleGamLA2dZRwul1/nOpDk
gvRiguxJHYv+3nEPURWD+ZIO9aR9BsgUB+3v403H+fc2CLm9DAo5U4hQNBZzSYiR
xKcGiRaoiwZat0Vx3NbCrdkwu7VcDtnGgWpZrl+r6MhBBm1KodOh+aEPnsCYrEq/
xMKDlL5sVP+ZKzHck1C7UehRtKZ+Eu6hWZEgCnUV6uuzTrFd7FlRRoKEemdLL8Z2
WpGu2ah7h/AxeBV0osRCtbwGX5U2k60vdAorXvEDufJsabhnu0MelmqWDywg1HtR
AbJX2Bv922FHMswDuT3zcRvlSk8/R3xqMsRoA4n1L4htznxMnrpGcICoP1Qta1K+
EQQy6h8UBHtpbFMmK8rbOgHzcenVFzpdc4KWdJTuFRqKn0aoYFuj2CXjnA2bla65
dOrGhXtqEjIy06X2x4TnSBMlC4lmJHepmIcDrxIhgfFVHReJ6XX4AYgbN8ti5STb
YwjlAgjULH82kRBD8bpW9fGBY9zvyABlBfvolFMM5F2rfUBy4LEGL7avv5R94C1h
s38fMBH5BFr1VDb86s36oWokzTEf/8J6/zL0xs5v4/67rKviKsqbxOrDq5MVHANm
X6kifawt0RNpLEstyQ0GsyaV3DtyRSScnZLONDwKIiZR8R/ASY/ZJsL2N2vjiU3q
BE7pUVDKxh+mLMA6SNSG50k8n+pl4ohGd9hT+fArGHzWKtlRLCx1LbeFCIVIb+pz
67aT/C/Qp4gJICluHNeOE1HH2fpKEJXdItWs1Z0u9pdt7S+fcRYVYbPl4jdpeXZs
hnZLlgp+IsBR3lTd2KTe9nA2OOHGySUKWUOb/V7i/D/EWfVBjOQwjRMxVx6EQY1v
noeRoB1hXteisMrY0JlARLoQXR7QVlFlyjRsNnrZZqvWzuAIE8rUV2ba9c9ry6ko
1OknA5TnQMUUXaP7KdpeVSBdpiPQYDL2ojDM/YBbMbW8EiMFuoggQP9FhIlq80gQ
f4Ifksh+iRzCtZ0LS2ML/ZJ4FkAd4bNEMJyPs/8ClYbdm1KuZV8lz/pixixbX1uX
jt3kvCyTXQ2mnxt+9nipQM9QgYTSL2Uu8aq3CjRBJTR/6zgLfdhDR360Mf378kPr
NgrxlDE2kEzWcWvx90hfKtLuWIBvsftLScbEPSVRuAxjAy3c5tdpDjQQT8BXa+FH
sUV+yBg48oKT9fp6t1kfxvb/uvgjBkfRq2KmeJhPylJXj2Rh7laSaOGWOpMhjsgq
fyTkf613F0xBfc0xw/CYYg+Ieo0+syzfbPBuRFKx0di54M1IFULHAjar9DTniPu+
kNo8QrpBteJ4qk7CJgZs99YpXA2mQpYajbgcQE/WPl9wjmG0j38IEyPv8P6cPFJR
5uSN4hyorGirDc0Bu6UKHDFC4JVhjrhHi2Ri9u8sYYcWJAYuFGpsJuVN5alXgDk5
IxvjAEG7yZ0lfgkkyQqdbJny0RvmuMle95BnOUv5YHtfx+btuyVUqPKGsq475Nz6
n4v+3EouYCURRG2511G+MyZrBntzZKNiDdKGi0+wlXyOY/ZhD1M90mVID6jb+Llo
HeLCCxCk4Z7jUZoObn9hV1ttNrXkC8PbQ/xF5qH8ortwyAvM91LtsJCy6N42F6xJ
JCxE5eWHsTLscs4nQgmymJwTZRO4DYtv/tcOY01DVFlr/5xfUAZtIExqriMW8Z0o
6kYE+6Z3KOSKLU+5hXbRLXaNfpLASuFHCuyi3A5eKzuTiL7cllsZ3WJ6V4bq06YV
CSqFyuUskZ2/loEiBBT12bGMGhb773dNYOegeg/ZSCqPpd4cwjfERHQdM0JEP/c9
hqXQXXhP4vw80SzQUefEEqkIVrLZsRLFLl/lyvcTjQBSsBHzZUoUqoalrm7LYLt9
bWDWkWm9vFwLCMTcgKoYndAbY3U+F98EZ+ZfFHrPvkI6LCeb1uIQiT34AgsF5bL0
jom5FsPJ1K2W9M3hNtoLpaqRiG7rFltgmpFlm0DpVY29eTpkVZ45eCKboeOtxhIy
zO9LzqHQ7LFnZPFVCSdF0kFK+mCWewNEebNCwEJEK7Jm/uenrZctVTL+QR4Fq8hq
xQ8eRk1EEWF8Rvza6T9AHCHpEaNWoIxDauUMZGIdSEeDun7POgXjfGBbx0xPNbgd
ugvrqgw81xH0hqnZAMZdmvieOKC84U4mtCiww3kBH41ZUjoEcotRaZ7t3c1JQ6la
/IbFaHY7unsIQXNOTwaMfZXG880FlayMu8Eph+bFbF6WEwqM68CsrdgslDAATCij
jqE4q7QYjoqhIGZEt/szyJlbB8hvVMgodYCwlSWRJM5W5wzYdYdRL59Kv6qTGUHw
nisvdYjyGq7bsgkrghK5vR9qd4MKbfFW5uSoJTFWMJVfAGGpgnzf/c3VYk2m+5FD
mT0S6BSayw78kyt2ZlwyYdZmJiT5D4JUk83Re/kun36RZlvfKRfwNs23PqmDF2wT
5YdlBZdgW/0EpWhCN+fs3pof2Kj6Z2jROLQQv94xGYDrOWmwCXRbsejTLLdh38Xr
DyaOhkqk8LXHBycDdJlKnUqwJ9qNuVPX7d2WsLOwr8LxMzmRG25fHGTNTLzDeqjp
rcoqZx3w5b0pM4BVSXgEJKO1A4JXBUCBUIAUikfLr5+moR1WfMpLRsKpX6FzgUMp
JL9L8PcHgTCoAeclcLT0s4jclJQJVAJYA+HlGXdeE5W3yOKzrdpW6kQtbNKvAVrR
PxhST/aPKfwSj3w1kafAVVWQdQUTU4nG8102K3npIjXLM3F2k8tqMW04swxOUEH/
pAKK/gWgkGfVGRORTp+PeKS8kn04ywymgsXa5sptaQFVsEivJ7OUxpB/ZoeYqHAn
qLSRgNRrmMQNxKz9ljGADndJK4jJLmNgfIsWpA5xMLzH5b89r0vceEkWeTnVvfXG
Kv+8GKvMGDXptWzW5+qq7o7eQxoTl6Qq1jg8dnpKdbxudReYn1+1o4SEn6xhxy5O
DMlrggdQKgQ/SZRAEtMmIcUbBz2o9iaxDiUSzPdRU6ph+gV2tr/Z/HjYA2ZfuVe5
n8ntMHfVIwTFn3TlOJoUuBUBAhowvHVXpaUjruOwGfyt0Eh7yz+l6IdBPRuSWbEg
PFn6OvLoIXDAaAj3iJsbY8pmFec1sjd0XRhl0HXGdxQYb/1pc7ffFdSeotyNNn3o
dpzqHE6/MyMARGTeTpOQR71ZumlGkL5Kv1nb0/tl80b0Huhql0c7meRpvpM3bYS2
puvF2Dc/Uq3G+OhrvFQG/sOAqbjjDdmgaCMgYk6ug4mDFxv0DF60ymRefZvdhnfR
95ufov+vbHnV+rsE975BW+ovQ716o6rZvzuZhb/EdoIKE25V+NEB61SPKbqTcVvm
go4pjxAMng8Liyx21ijeQel1/v8TiwxRsbQE7xGvO+nUNEWXKurTEc5Mbvlj0xGD
X47eHmnxJmaISdGwfHe2RXxr9vBNMvMwEanLQSJ6FcBpv7SJaiy3dr4et7NdI4MJ
inlyhVmhzs8QggnglwPoA2VyeGajBUQFLt2MNEHG3Veso8EuX7faAPwgctC0q6z2
Zbaq4LgrEDFxoPTF941FnreXuLP7bZXEVa6lnruDWn0pvG3V/hBlrSQ5vZNQiqkC
m1ZDSGcHUNcBZ1gYjBqeQfVGBx0VxV6GID5Wbf9aPzxkqeIpcQrFi37/iQJP7hcF
9KP/StvbRcjaXmb3dKIMCGCzA960DmTzMeAN/gkXo+b5v0rE/gOfhpNcfX601MpE
5VN/yGc0VHFOT6d90pFq1+XkWZztcMCjHzCU8yC4r/cs46U0pP40Xr7A4cCs80bh
Pe1DO576W/UtUacI1gOTQqIt/QW2L3OLp4gl6POu+gb67vVFZfaLu+AT/5Awc09c
FRP8X75tGAoriwFEtAxVESk4g5DmyR4q9JCtLE2zGfZh826O+6TpTBRdBLPGb4cm
1Y7y1b9i8TRdWEPnZEgLEIs2VPVmKI2jl2hJA9Ca5Leil+nflVEiyBL9dKKcdFzQ
xhlmEdqJBliWv2iXWN+gxYF0Z76BQ7jCMbCKWT5uYlaozSBKB0JBwm16/3l54Hjk
enXdAsnq9PDblMpX83DcDW9ElqPTFgSnUxGKglAAEWBIaJ+gWe0k0QZpEYQ0y8C/
jJIioVKsa4a4x92cqEI1hYVNB9iTmgd2ZN/1ycRlIyQ9cP5FxjFKtcoNAopuA2aM
3kjwDDNpFN1xxMvRvc3CJlgRj+XSxVMzBL1fT6MOs5aorJqb3/qtVLB+KZkLP1nD
uHAiEtnSpfQhpbct0+g5LH8XPeuJSTZgcNuPAx1Vf2xq+9/YRDyuOec6z2EGq6pn
HNEatXhqDtqcbYobW2B5jrbYSl2dr8ugGlxCprVAkbCZEQM9lE1/E5O1wJoh3b9Q
wwgX3OzwNLjQMrVe9aAjhk5tlgmKfYiIeQCBi1wWSQCjRE4o/fV7dRJTAho7Bjui
NxThwzX/c07LCIt28ZvVZd5ErIflBNZz5EW+ZbvXV96DkGjJoc3U7oaB5TCu1LDY
iK8Xs76hyVZpSb7uKBBnchtngEgcFbsoS0HFIgPVJi8vu2+zNKHtoXH1cJYVkKZN
4lgfZ9PC97JZrO53kvn0UXjegnOMalpPpQQS5oA0NJDIF5okg/nkozqrrOYXHkuu
TSthSjJ8bci8OwUYclbuO5QNShFI0VsOBM+9d946Xzkoghvhztg8LPEfHRihxVnT
qnieRO245t2Bq5skKiClnR0o3Q+Y/TY3j7Hjb9kLTjBy1mkvLilvFBtdxA7biHUN
Ax4Xja7WVYX0PKbmnqapld8JmqrKGtxZyhqib+fkP+8lQBq2tTSGk0COyq1XRk5D
tdpsapOEvJJP6shp4fXbSAOibtGzTIW3vD/LUh6jedVuQY6FJ5qknZUpqJmbWEAt
Gae8An1ldTDB/FMD/zh53ay7dbPiVy8b2ULXMe6Z63E/VvK6uKbfuKzcHiuTqLOl
MPmoI/jLahbNpDNRVMW8FAm+X4WlK56BCeDU4dWm2drBJcXVMAS0V5B75ocKDzRf
n+2tZI32irvKmobJcf97fdxvbHBnkKSICYXDfPjisUClEbwRPgp39kEn+KhdYYFH
SbzOGrXzxfTj7xCY3pjr7yRxzV2jLAJaZuxNXElPxknOg3qz2dXyGThQY2pJwkwJ
1RBspOPsCt5u18AcSeBbptPjmLnlZvZ6r0C8d/rnPwiJlLhvR2kxycyfMt1K3YRd
gIhN9C0YnbmlrLJkDuBPm+v82AjnBZixRdtTh+WP+JXvUL+6sGNHgnAV8YBqTF5p
6sLaeqvu5A4JCaCnOqAJM/XsNthkf/iBbxaXLgqu4EwHw9idNlLOY6VLhHSKRJlQ
e1mSzFCpQsL1sKuGKf00hpvdyYqS16qOILJysdrnuGjXwG4qtTHKXa728+8NFFGM
JB6911aVYQCjjlqLJN/TWMiPB6DZByGqxjsM1R0r5Jx9Q1KUqrBfPTHgBpRoZsdk
4rgN8pVB4o+ksryH6GgocqpTG6p5jTYoV8fOjbn7LiEQcDX8PL+MP3mrzikSQUvz
5hINLzFfSjzY6x88jH8ZfhmObQywkapGDF+R1274ELECezWDSChmxNXh8QSXEbDQ
1QohVBcUTG2uEbb7AgOTxz/iNWD5GEyC5aGglYPdVGPxAFilZ4SjySrSR1jzUhFk
dtKIemZn5qFs2IZRr7RNmUVpE9h0ixzrofI8oiQPr4dDM9q7McoDDoIR0D1rBUZa
XA5/l5kv4JO8c/bGYe0TSsQ4zD3aZVKrDT3JgwLiYF8KRXSMYsKsvdnUR2TrrYjp
oyl2i7DcxVvzo9zUJSE/WV3x9gO73hfM9vBPDmukL2xt0lmqtN2lGM1/rbKz4/vX
03ibCU+eI0nO3RQZIN4V/BcjcOYZBoc4aDW7uEtzrubXpr9jdG71V/UTd7eN7IAN
y0rFh03CdSTkcwcMuZc3PWRM3Zv36/7rDWF3/1lwDYB4tPJV7XPPforCGmF2W+1G
YM/3PxclZC3TKP/vgQ1BwDQ3ggPs/vnTiZsxA57s/IFR53ZJRaW7YIor66RYJAMG
fw1L6MNOjxSxgHezgZOFXBNRspVBMQVxp23qeUC/3HSfumv0KQ/JYQuFL1LPpomu
FHJT06TnLlr1J4coMldiGB6cdKu020343qemIPH7b6mFzisZLgdkf8t/44HtQ+be
u+yBJnP1hEEXvZF+asvrqW07MLAFELeDTFEKBqnd1YsmuyD3dDTymCzb1CNO8jJU
RFYP2bQxpib0fhYbCW2iAbopPJXYCcbyMCHLqogZoDdnksZ52+oA8ajWVeATMiq5
fGYWTxGRA8dwlVbxkzj0CMJPDdjZWc+SB8krD1CfgSgAu8teN7HDEXVQbMebI/Kx
IXHuzBnFyyFBk2lpTAE/hyTZpameov1W5CLLgyyVBmNsAXxbMwW//+Aov+zWXH1M
G2SQYcT7+WBsJipQEIdvZh1YPJnopLYZoicwkq/HL4n0wSJzJPOCsHbm/8nj6e9E
SYx39tT2iGwIcP6kuEF2w7h0C7pOcUu6V5oP/6DSrK2aH8DamambRGgi7vr7va4T
Ci1JimnjB3o3n+tAkN6VNREwr4+4Avmh3jSBaGupTTp4hY5dRl6QRsObzqjo35VQ
EDkJNOXLg+73BBd3I3wpHIYP1CpgOmdj8M6CGaZU70K04Sbwxeo4Wcxk3JTrcPcC
8z76j/ugfVvGkop0SITLaYs9Kw7tErWVAvKy4YX8oS+7ymn1N/UBllKEDDson6ii
x9ZTq86HfDyaptqhh/DsukH1ManjNdxZIPw+8G2IDfneZ70Fs8kZ7717lrLqAcRb
i8WFVlr1J6SEPBXwTGd82UTbn3hYEMSuuEUrAVdFEdo7yg054pxrQCKfWUjCqNrr
FNNfWMy4G10IuaEGFtBacboW7GIIOlKSbK+nbfNSC07CC2hWoqj1XfxwPrz865Fj
HDiAWILMXtE3/BuQiJ0k1Azk5TdR3+BQboPMdrT4/vf6zWYU+NNLW4dbqckKkska
XB8Fu8Xxg+8WYHjHNofJcXGXsDl2c3QiINUFGprmhwjkzuKLl7ldyAGhzVg6DHIy
hdBWiKtkDVG48Vx+ivCWrKmpOJyWAFZfh1oag5uyghySeT76sC6p337iN3coE9iN
7Be4OEftaf7qBT1oMrh5XqeKeNwFJ6DM5QBeZV4j/ze6pyobOL9KSNxWihbuS4in
r2jhew1/9RI10ruIGV6G7pYOS/lP20EcTeZ5BUFP/H0EbACnUQw5Vs5skJtRvnUb
I9YDk5GgK4KiiiP/J9XnyxflBv2dphxgVuu4qTvi+xH4f0CwJWy34nkLzLtISiuv
Xhgudjj2/fnXCC67s68+aYpkY01Neg/vC/xgF84Rp45Nd0ZVfC0/brLq0aE1wjXr
Qkg4OiR0yzviabViCRi+YbbwLeGah9O0tNp/KruIvyJZpg8ZYTUfCQtjXMuImg0j
Dud26DcPcba2g3mCs/P2tA4UShyhUtMyig+gQRnzkCmivRS1+kp9iHJVT7x2oZtC
jD7FlSIzlqLP+xMhV7Z919h/6M5pz+n0mFrDPc2sauiAYuiint1KnSlnthrDF66W
sflTSm4EM10OPLzY+zR35VublJLgQ1QAWxLrT0kf7DNz8bQw1OpG4MF+oHXQDcQ8
Kzqv9cJ/ntjz68npjQD5NLi/A36bKtbu1/eELs+R/8iSxo6Gfkaco0I7oA2DVXhZ
NZs04GPboBG56YGQJvRtwjri7lGhD/eoKZwtmaxZJLb0rrxpSoD/1ngDEF2t4B1Y
9zO+KozGI763rpio8CsFLF968LTy6F/TorklnlJeqVQQ4WAfNZxWGf0BHiNTP7iv
bg0Co8hBoAxlaE6KZaGaSFhRSBPCBtC0wDfbvGu4VqQEXcclYAvetH4a+NT9kdJ+
zt8Nm6gR5upsaFIj/4JeixrqGjcKu3xM+NWUrcMUbgFzDbuG51LFs+TWISQxgypK
tbJz4d9f6vqhKy1xtB+xKtEqXjzuonZjvD/uXcYMrG/VMTUeYAfvUY4Hbdvf8VKy
ELk9ng2lqQuijAiFL/rOX9CEN3kX7njoIODymCi3EgW5DpuZzNhE/xHhpDF6GKzi
U1fFJeISbPg1InjzWMyPWfiP/KNPo8NeCwX3tY1cOUJDW370sm7C243lJFI3x9Yl
jPT5LNwb8GvG62iFAAQ/dG7ov2tfJyIXmY9+6EdwCd69N0JI7FmRT1Tf/ZBqg1l7
pVlYBumhd9ZWdExx7VK87Jx19ZNOWMO5D7BljJRT8BDRQ/HEaZgqnjO2z/RJf5Cx
CpuM8LNMce+9eoShaajETEVkF4fZCEH0vamvZTDsLBjuCsEQN//EiSGKTZUr8P5S
P0afIBson2X/6UJd3xRG50V8/As1l/Wc5U5brVjtwV90MecjcLhMvKn9MP4HRSXx
qA7beb5wiEXgefRwW/A/whGltUAcjhc0RWy5V8iWqU6WkBV9ZAOqbj2fTnuFTPNA
O6xcXPpWBLg+OMpRRl2u1CEt9FJcQfW+V06jzFESGD9rGRFqmhBN+JiMUDwFexRR
tRjOvoi7LPAmQ4pJp3hHJmpcaDMbJugNXSwHSu4F7cDUzT8F7t/ryfFZU8i91Gji
uSwl657LeQO55S0ZRlywBC+ChE4cGeHVflsjFzcp3ECqCCUEdTsBiu6ii8wY78vy
eADU0ljifeQYyz5R5WEajOBf51O+stuy/i17ekqrAMQMy3j5LeeekBTN2FMrcc0x
yxVBvME/0JeR4vCWRH/fQLXkFAz3Hm+cIva2E+CrUaJCKKwRgJn66WDijwRUaX2c
pD2FLtsdafv2xt97o3N2Fy5FS/Wbo4oNzpGLMefwzf0RoHb0KDSFADxaQRRP7Qza
3SVPSpVItBbD8BlfHJ15ofbHl/lj6Ge70QelrtWxrj1psW3hjCX/Q2OqzqzeZML9
9RAX9fjPpBbHRZw8KCsCS+cFUBhuyyCAbBf9YNATt5D/y5kzXVqtMtRJLR71DYYE
hH0pGqHbnpuKokfNOAZUb/z28ySP8FUjc5hLsVYTV6b5B5rpggBJ8uEvghq4qDXV
9PqA7uaSlBwy8PuBKsw4oAbt3gNnNnYoGPtOwF0RyVZZ7rq9wHS1c777pSXjbwM1
Q+cZvFQ53Psz73YCbSloQsxrzSWvWhI7PZqy+2iO8G/LmIsCr0av7KEG8aR7LiN6
RGpLh6oJjOvVcxoPFxkc2TwgIAkUZeHp/Y1h67peDZvmJHfYWwcynsj8r5P5Zhmx
SY0oU63XVE8+2MFFzQmREU/bp3ZTG1MgsurbsphxM4Q1ybJtnkg+PBGGVkNhpVpF
IshGXjjsJDwlW+VdaHw/ww6DmE/6gHjCBIaqcVKTD1PcEOYAsIUCWtUPfmXlA0nt
NVkKCPKt4IelrGyw+bBWWMPkn8kQaWRFbSg6k02q/T0oJJbUVhSD5e4NLS3k1Ycg
3h1IcJMVB7x5yDuhH69ONBqIp8aZ+VD1iLxUDNraTbk8U665kYoig3/EFFDmdCvh
0HXLlbqcyKxj8zOnAc2vfRrXhEq8qylVTxVzQjlg496mGEySyHLZj7FSLvmKgYxV
hLIbpk2n2LZ3WVi/irVes7PFA183Je9MKj4DqN86hLL1KvUEZ04ZgzlGQuDJdcc1
jY4ZFNGxKBITMRiz1yVK20q+yiqQRDGAzbnCFY4QL602rGgfYFw/bY6qU838TeLn
oIVTJF+4bBMzLzbUR/8gfE2dOBjH9krWIh2QwOA0iAqGP6LvfNY26w9r6/Jui3uS
0Rk36wWLvyXqxjNYAra5fvViRjF4qQOnbi492ZRnhM83IRiKwxnSIF4wlq0ndzhy
NHVx4XOAK8V6b8hhZ8sF+thKEE7NOjRabJZLG7GoFMTEezNNiW0j1O3qXf5Of9HZ
iRPAnY+OC/ubiLRrJcfbT38oN7gmCzf6XzenGTJ6BiQEutIFXXLOzQgiAvr25P3c
CdEEONO55wLTeLFP2tkPVgyxCxuy8wUs9r1KoM/1H/CtPFQJBcnt49uViYWQCDNA
kMsIohlcvPXyWcfhj9okqtlqOPO/n0Ft6J58QThhPfvySPtEu/nmQ234X5mBAuKu
YIx2+Y3OdlRBVBuBMF79k0hivPr3rsnyfnMEv7jiaoy695c1K3aa2WUqkX+p/0iQ
nIaF2KfUXaiUgYlHQKRiiXZ2dxEfIDRTk1c25RD1i4TfIWeDmdmehg/ePa020Ey3
FJum7PefqHyz9EOby4i9xPXSosKpgc0ebda6RBfN+cIriOxoDZDjyvFUCScztPRJ
XuECC6l/pm04Z/9VBhe6S39GaQmbw31ntTxwBAWbbc5ZH3V2CHq397TDY0/AmD/G
dwoZleL+OlvV+h5AAkHHTh4/xEog3YCx6Muwp8aO7ocDUaQQJLa+PkA9Zh8xjmzy
FNmKMk0dW6YseKOL8fjAx6axiy6oaGIJeBciHBaZwu9/S0Obf7PTW0Bt1bL6VCW0
SrC1EtVJ73qM+jf1uBnxfvnh/fHvK+2QU0y4qdWRKpSLSjD0s3voMotp0izFWFA6
OUzx2CrXFzXACeNVAVbJrAEKI2Q9IGzZy2SLMjp6u/4x+6TAs78nZ6Hc7hvcEKWZ
JgaoOU/fSxLd9UsXsaJMdGFdovZ4YmCkRXwYUrEa+xQsaLkdZfCIFq2gSia3cE1Q
lpZ+S/jPCAVGsqSIOuBVAEy0CaLRwb0FncBIDJ1WyZ4Wzs4ZR6olSYVbQCn9L6QF
3uvTQMAUHQuEWViLe6rjpU8kFQVXsC/RQ4n25HQ0WFSejQ4IqoHvVahm2Q0hxl4k
AzIS6Z512cXibfx7aDmqbTGdK8dftETiwXqub5A8Qcjs13ITZZvkCAg06W5ZPRys
SBhQaKomvl7pT7pN2851jt31I0LvQH2I3KwFAJLS6079N7OUXVCy34ugFUXU/NxK
jg3VXSHgo/RIcfh4fIA7O4EkL2nJXtYVR/hnZ/EXWJsY5VCCczK0XQ+7RbznFWV+
d1Rnx5uvnTFcwIRagpdKtMiy/70nPam5bS+vwdOZfXsVRzq0ATXfIVkXpZAxfJB/
ErKXmWFSY3UnNdKFUM3XTs6CuSn0NXQsnuXDiAJxZ/4dsfVp/4KG5oqio7nlr0yr
kkSFSPFryDrMwiu1u9DTokR2LzK5VA8GPdl/6uc/tvPH7TOzA0+x3Zx2d6GGZuFu
ZJVuOwk3ERm498ytOeIc4PuS8H47NR8kfEneV+yoX4WL8OMhMwa4pr2mo2i1BqOH
/O2796abYOX57VXAbTp8pdEX8NMgpT2WEBHLWsoG4ZNZ2POM096R6fvNDB9KX3jn
6UAqgFA4N7nqS03UG22WDQVqbveI/8obsr49cmNdUquJWalVhJUFig60P3YJY9zA
H5Q2kYw73OC0isqW/Mpuyls4z2O7Wg4CylJfIegHcHKZ1dJPskKbFNTxOjMYpZ23
K3bQYqvc+l7MTH7LsqwcmtL5XEBUMzrdSXvpmd22/NoxQ/hKFqbwU1nCKPmf92pu
YzQYI43Q8OqPdmhMVHO9LGgzyYcvOrmUc0rP48SqEPXdnhcYkPB5yg4PdwMbH1on
x/GMZ5L9YW0uwx9ycBh4OZWf2uMC7hOVa7fS22pjO4mkRYunck4uv/Kuqo5Mbwbo
mJyFuvVNednqtO9aC1nGuuMFIGLq8HBMYvg2giQJuvq01f5XPx7gbVyMF2ebmQd/
e+REsLkgfTWsPZFKJgUZITErQ0LmdLt1PWvnziywZ6ZRsPBLRe3+sxGD//R4Yj+m
TthCD+20A6QgOvL8/u6qmz/3EsU6MmYYmo5FOW6MimmRIhNSy3lqDuYVGUjq2TZ+
nkyJfP5QJAeh9tuv/zay9/lHFuSRYL3/D+eCBHr432kG4pAYESkmFyM0895u8s+O
d9oQkH2qacyAxhJJnDGpoJiYzqClbzAXl6s01RsWc1SZyQUtDDX86WfPjkCIlYZ+
evX2Gec5PYxqRlrX6CtDe/XpxMJ+MjLtFDHGmF2/czx+vWkGMrKMf4FQGlBefjsn
CohWdI9+qwangC77EuIz7cZL3HUE1IC6Ex6q8xkDzkhcplxaGnZhzfySwQj87aK0
5b7AlVfvuMR93Av5wX/PJKEvI+Q2Te9T4yU9BLTJ7LYt/VV3Skfj0ylX8yOmQ/YD
IuR/hj786ZBL1vlvEclYAanAaDkwSW/yAumltNd/QlUQwR9jkYoBwAe1W4aGXRDZ
Jbe8DxUrXndz1faP0wdxKhzLaONHHJyc70xWVOSqwzt5EFLlNTvC9EGWH34gv8le
LLTkajBueeYzVQdG/XgLLcbyOjZuJWulr00PH1FrQ78nWS/BV/bc9UX3r+PCFGHt
B2im9ctOwQm0TTxKSgZ4ozZaga0YbSNtEb0oRNB2JGPO7ZJwYJYDNb4f0AqMSZU2
qgbLEGhvUXy37+0VTnJOcx0IM9rlQH78nFOap2wGfq6UEOaqq+lBZzcSSrY+sdiK
iI/O0OyYKfO+J8NJKo5WoPOX38hFfKTLpObaYl8j5H0ohcGFcN6oxCTq7eABoHAi
YNMY5w4cxJJgwPdyUuE+ow6NgAkvhMhrVwtcK6Ad+Wl3SbOswx/ZtcTeZisQs0jP
QUeFwcuKTSbxrG0MoiU1qULJ8YGLf/p0Wo7wUDBxRSMsm8EpcTc/3cvdjW/+ZOhd
uPEIn4JKRTra7BxG3UqkHL2Lcsw/vNnIP6cNyKcfhKLb5a0cV+9CbwmUvE3Q4SFD
f216TyAZxq596tDO0kCG5tToyT/9ouH9MQ8Ji/fwaqU2VoFEYCqZArrBTcW6Cwhv
/obKO5VE+QhAMXti7ZFrc68wJe9gtAHanSWL7uQCc3Mo/rZrYTM0Bwx+VlIbz21E
J9zWuMc7/WbXVNoyDQCQRJl3c5G/bLnq9tisgTxL/WEY0wrLdeO0U0x7xpNCkqED
h7sUB4nNZdmFHmelgwRePQgCjWsWaOa3NF1Wqd5jFrVMQpUkDCydDPhKMkzbXlAR
59wOz+YTnc9XN3Zh+kQwm8v6XLmyNrpr4AGFBXdD+U1nGr/SEMj+kKxyNMSakX8S
z0OQoLqB1VKGr5lGydmy5yCQyExCaPLoyUzfdCj+7a40lxfhZfPWapDKHsEI+Fd/
omuuRI3zvYF07gmuxz3h/N5+VjB/gYuI4yo2Py5XH62IddyOZOr/NSevJC+/ckGY
UcBrWKAWk4wm5pT2ZqSwBQ+v4M/C6AKIPVX58hvqz7enFuz3vWznxWbGmjzBj+LQ
abvlz8eAlw9ugy/vghG3lgyD1DcbKAFHia8nNYk51ZgHDMMCKGxVQv73GMVawS2w
t10DhI4WLyX2/7Q2neRSdQgPuMZhQC5COqHXNKY3MwqGscbvuiCRll5a1fVHAYnb
3Cb6NH3kY9DtoyVSb9cggzRq63UQLZq6kuX2yS06GsiNRmmydMXpfoGqMNft1F00
Xu94aFttMvc/+/NVuO9xYBZi6Gu+fynwO22LWr4trOfiJ6b398+5ggui5SguvJhr
GSLygMBci6RJTlqUcINYOE8dNXSI+s/mR5dS+GTmFiHvIsK2bV1HmjUwlejJUEX+
wkD27mpPdW79o/rLHcigZHY6TpDfWiFM/Ade6Lv+rv4sUJh6CfXfal4u7K1SmMJL
3pqx/dDpAUGy/ZST4RfU5BJn1BZcIQRNfus1xIuJdH9z2RyYJNFtmZ61pk5QCfUm
Bx3iX3M0okS0spwBwHFUs+ZX2mbdEHWd0JW2MXhOl+wAGWN39AhYzIr38jlUIveP
OXP15HcIS96tZN/O4wqe+Sb1po4Fd+DfNOD7UyzmUESqmOiPxXLFSsMMyEzDn1tb
sVcB4NzRKMpsB5ERWIt47KGP0QjQkVHYYWA3DghSZDU3Hg27o5APT9SmhpSPlFsq
xXHkmG/IJBXNxd3LIbsQAMfm1UfjMc4LFrDUk6N9u1DXR6N0RFwtEb/1J38j3/3I
IRBp/W1DZquiF8QcQZumR/RWvHFqEqWqGxe47rdJ6MF2cyfeGqxdK6RUoF/ktTUs
ZcyfpiEuQS2GgKfEc9EpYAzpW1IStZX6vis4gyKEP5kAKQ3ccWtlICSXluO3kbNF
nphm5eY6tR5GwIhNo7tD+Gs+0xSY5GKxw6LGvyy8i/hWIVMHMc84oHHWCIXZHgYJ
1qnPdbu6Fvu4a4Cai5UPfumZUnPDyyp2CgFBljAqUTC4H+qjXQrXzG9DpgNyypzO
JX3L8Nl3abOJCEjchwmFd2NSCY6GQE7tmkFHygXGFb+x+XsDLWtR9/F4mBbafsJF
zUKeaA/iaNhIzk/Sff1/HgjwBRbrWZjWa/KabI4SjoAhHwwmE/Cy9U3wrk0JuDgM
8Llb0GG2fa39bJlAFtZxk+xs+WxjoP2xRl//Hu4kFxkIAqqaKEf644C7vrCVoSfQ
y0xwsVsrtKJOPop4wI+6kfcPbr3Utp8digGmu/34Ih2HNhuVvr/T+3ogJ30kQ5CS
FwyJDovzmRog8x83jr1DtJpOeMmUGm3qaBU0Mv3S5ZYVO5WOgM0jcSkwOlYD/MR3
cKzDQYckFIlpDHUA8is7u1c9FY+l0aeqWk+k4orLs2lvZDBo1W+W+QOESeZWPgxp
kAPApKjRpnyegPP6Z3KFNze5ynVRtRxZJyaQmrpv4L6HQMHLlStwcrpt3zOrQZ/Q
z5mFydDzRkox5KxQnL3skK87rGhvFg2AfrhZTAZ4k9/ySfAhPYVq644YpoY2ECWX
iYuyzGD2K+kZ6GF4RySGyn8SN4H12wYZ7aQbulVmQwFV+QIfXpZYGxBP07v6AIV7
jsHZfkHWSKd58EXJnglOiSJ2ixD2QK7Hpn4CEr06gAF9JKNy9W4YF2THFoaouW6C
FcMpHKjqALGzxcGlgbiC49eZPh7dKDLuwH7u4Jyf/A0Hp8ZkDpZN54rz31Da1fPi
HGC31vpA5BfCiYnwoZdncJWof4yvU5LTJw7u0whOgVCu+e4qpo/gPADFdjLJR1eL
2WgmxOETDVr6zprHooMWaad46siMAJBKU2CPLvn4BCp7b09JrUwtvNo9vUmFH9m2
525qbraddhnngWoVC3Ztz6DzghCszj6MbgOEW4Hhb8qYDSnVHCLz4g4z1oav87RX
dzvYJel0Le/qhw+FGQ7prAG8zSluffE/ZGtgoUzanGy+MTGRPG99WR424NnyehR7
s12CGjwVrD9W0Msi9uVRJ89QCOhtJ9aFLhBkiLgXQBU8m/vSBtmJAyAlr3p36esq
ZaosE7fANlmnuxJgi4suCWZIij2lzeBBNGP6gNLu1Scmlp7H4khpOXR1wSU7MOuB
mYg8AWxyyHfy/3o+0APna0TMrOhuOlzEr0iDqcuj7+Ew3Bhk23YgeJ297HRu6kRW
DqSkLv5UQJdj8NGu4GYHGimikHtvdf6agUsf7jdWShKFZe4UInVNSAzOiFGy3ts3
veOJUST+NKYzqbuymJ58CttLao6OWXko5lmW0lE1cLTGUYLVq0c5ZrYr/pSTjKoP
SZg4LW5iYJKvRXM+Ec8fZEsDG1SGzULzf/W7bOSPlGU+OFNVIyBDA06/Q1/eFVyX
3pKWG/YGu4qtxP6Yujb4GP+0scyfGeA7fh2gAngSE/r5Gy9B+/+B7/pKfFa4HUHs
s1+0VuWLIR1A+18XQsFqQ3i3WiIPeUaJTlyE/AqP1/aLr01D28sJf4YInud/CvGJ
l2n74w7PD2LLIgopkoKsV+w1PSC1t48b16i8HnjZHtrTheKwZuladuIuHftutW89
fDQLva+HeYFzwcSbZUslMFNa6//7TOZ9gM0tCBvKym7PRt2f7OcUUDyBw1w453u9
OV0yG01sGA1/6sW+InSsgHYuv4Pj3H8Ql1Jnh1lmQXRcVpLah7ZwJ9PSCsrFNxm5
l+Oc0n2QYxDoX4+RdwFFhBn8nTnTV6Z72SY+92BO9zCfIfQJ4Z60XIFoIlQ9ye6U
JPb2Ve0kqsJoo6Tue3Z5z0v6+NIqoT4WoFvBJ/dvtL+eqxT3pwnsJxM2v30VVBnf
f5V0wkse2yGLdxYtjs8yLr+lZ/IaWOr5plaiQCZPoccF9QrK3Ob8girLafM3OOCh
TyE50QRc+VYRrTcwnA1+3wpbepk84xKVD7BjXYyslipEV8Iz7tixTNhC9iRKmQcj
AhT9jG089gzKPZZGU013G0aPK0nNoOfCbUTVCA1SrufNSDlOv2s8P/7O5g0l/kr0
MxWm8JNonbgqXNKi4SHXpdMcWvTjrqJ4yAxqKBEucyZBML+2O1Wq8IWjGZGl/UCY
aRtcm1sXCY98vbCPLZVLcDHiM8HpXvbwc9NgwoYFfokMivaUTepPCIxFbrYS02Rv
Mkd5lE4BXX6B6VSisaJ8S6IFchgrTpC+Hn6vaYYlsFxPXHF13XHTLQ1vVuZ74vLM
hlc6kqBWHuqT3pPJb94YMudakBcftJLRm6+QXBhQxUPI2mSLwUPXHS5NduVxN90H
Gx6rW1gool4QrzloAzVa3Mlh+fKOVdCGKI4BZisS/OLhJmU4fkapBsyNMOLd7nGh
zXO+XUMI0IL3C+nc3p27+Zdcnq0XWLo8YKzAY1w0vV7Lt0Rlu525U/bA0iOhRAE3
IzX2MUZstgEPhh38B98RfKJReQ+XoQNyc0DoiVEg5sjGmc7ImPzl8rUVogPVaMrC
IIAFI73DGcWSErF2ZLGCVs1Y+NbhCQICKiY7J23ppk/1AeiQiYgzDjNRx6dQx/+v
C606kcSzahxw7IumXcW3GPwkNPV2ALWFJvKohw741jahOIX782VD7HRmJy1Ra/vj
3QkMQeVZ8K61BSrXUZwH6LVuRyf2zEJmHFPg5c59RNBemMmlEC4LDe6BWWxzVrgg
v5SZWXb6374mhv6bGNuctdVPyNmU+gsGPJZH+XhayKo9r5OF29nfi3RoJ6AiUOY3
gRktIc0kEsfrFHnDj/2S/M+GTjGMgRlgOEWB/jPN3Eq+FOJvSbW9VtrnH1lI82hK
0lVbvZsUt/2e5/F4nW+qWAL3vTfZxVmFXM+MDJqjzPEg3ehhZRe2aZfQ4xLvehGr
c9icjeMuq4Ml2t5ODKhQb3UDOkynXH0Q8wCKUShGrlSmfx9eOz9AUsmbx7SF25fZ
oouWhHpcyZ451jPATeBeJxmb1gmWyMfpf1gk2A4gjOIdSjFSP1dMqsOVUgzymqK+
BSmIUsKfd7IaYdE+d17Q345hbIS/TNG0tQeQlliMu2P1rjn+Ql0I+HAu4nKN61j4
ntkk5OBUeRYZD+yHbiRtSHvv+SfSX/9GPB3yDW82wlNkgn3YMU4tKXVZsrhclSl3
HqUHesOFXITxaS9uuORes2k967Ac8LZ7HC8kmjHTKWTOyYiDb88hRxAzLd5RQ1Zj
9iXRukWnOVj3mWe3UVKSMuXC4C/mUJ9Xkz3nz/TAvOAlfqTOw/dih3FWUrkGz5ZP
KJa1d1k7wQfBCgCS/XU/J6YuADfju0FMD3vGms1p3E9GbgGUWLRjLREJukxnCd0p
YSxBmR2szjMZmlPcU/ULgmmlPrzVtfzRlOzKC3ehJxg6fYDCyCDkCkdv9+qloeGd
Ro0M4WkvxUOFrXSCv7l6zx1fgUaqt8HjHffeldmxNhu+72PqJcl7/F3QFy3DFOvm
XQl3cs8DFVUw+szfJeTwG4mYofGIV+TB+LoQ/ZECBZX7dZ3aKdpI5tSoXkntaCie
MX9f0lp1jaNq/Fyiea2iYPFziH4qHntucJ1seA6X/WICoZ91OkhjazyxpaI5dwQ2
gWGCeTnABWHpCVz3+ldu1sPtqmMw3Z+LA7jqJH1K2u0wlTNtDYulFWpXYttNSzEX
smPKNb3DzQnA4ZqgPhsY4vaNpuR4d80dxmYoqoAU6Xkhua5AvOPzBKZFNHg5AvGR
U44I4n+JKOOfAXZ5O/BwHg==
`pragma protect end_protected
