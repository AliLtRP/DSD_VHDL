// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:33 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
hvAj+bUjahXOZzK8Abq48Gc/uoQie/tZCEnrpd3t1r7HYp2DwsO/0UFjHo40G++I
TQFbORkU39ms/SVjX4rWoRdrDVTdQQbD1osTn/06RkHKk3KpficnT7C/BLnb3rE6
K+nqzDkFgKERsCv9DotmlEq4+1X5ZrUatOR+6yU5Rfc=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 19248)
oKnE4oCQDh4cS58y53FM2hS5B4a+KcUP8qyVnysbbnQ3h1BVKrDC83XGyl2UtgTK
cSKYruN5Uhuq0JfjhRCgm6xxEJbBE02qjZ5hhFHiaQ6yUwBJ2XD3ToEszQ/CDidn
JTR2jVim/M3E/+ZonD5uSGqBQFedYgu5JHpLPiGVenozlf6ICGlGlInLwQv8E3Zd
q9PjQe+TKHk3febq0VRjuygO6fFLGdgDMY6SLZ523JhlYl/XQ4soYDAqqd0r8Ekh
ktTjKXFMgmsTLLaMXBcfsI0DcRrDWtE5f+gZDj2ecZh2kRUtd5x5AprO8mDQEom+
R4eWBPPOPnPSGJ+TMyKjMheddyNNkQbfQCDxFTOTvgN5TIaFW9DVUG9gHm4hTd7c
cer7Grm+oPUy9lzksxYXXsKNVIWXwjQal3XOP69ws8OMdS4GSC8GObbnkK2ltQyQ
/Y5nANbDhkBox9QfawVxbLJPv+xcqfaIbCNduUk2+e3ZfddZHF7x3t6bB55KaUVf
Ry6lUDkxGrS8UjSZi9bD4suYAtepwzAOYwpkKjLp4MYsLMZquwjPPLzSly8m8d00
6ZBrT5EpAnl3oZ2Y0UmymBr6kobD2lXtVH58FJEdA/VhPaLQooxjDjWXMr8ZH4bj
/FAAeDwGv39iDPZyao8IgE9GHX9ahZxmI+cX2gkrL+Nvcys7dJ5ghr/Og+sXS+Rr
erXT4/Y0cOWV1lP74wiOTCvAS5PCov8qbR9Fz5I19Qj31fvGEp7Zk9ea28BmQBu+
kfyBpzlCCFyMVgJVx1ocMvsTM5HwaDChHENeAdJy5fYAIC6ESomOQMOUlGnbya6S
7rjXuIJHe1MLM5oASDHF5BUIuIpOz/MsMge+Fycge+Yx2NT+H7d4ttvGgVv/bLQe
hC3NtXS8fXMWw2siMyO/T7kMn+lL11wRb8cMl9Wb5GWgX//RU05ubNGQFaoothjC
L5dciVersONsZSyDgVaD3NfnVIuXvER/PzxdNfxGtViMHEAMygGbyhbLv8orZ35Y
mb17Eka906TKP7RZm1+eBI+QdkyQBo+8QpVyJ5r1aKfMX092L1srq5LiWc2gykGG
1vd5lvIliHzc588PbnATfudCA8D3OQHqTYI2Cj8+5mSCPTqNeM9ZdehDkUNWu02b
h9vuPc/ySJijeMBF8oEyzz180EfV5QtjhJkOdxl+gN6GSpSGcYgVqBcYVGhRJZc9
mhLOaTmCUSueKa8AeTzt2CV1TH1HvD4Ay2zr9mWYXSLllXgHsk0cNlls1CWpT1cr
IKfg3niZ3kLKLWqgMDJfMrDGKJHr/fSIvhhqVr8MfpGosc2AaxZhZ/vFrAH4fj5R
/3+tQiA8XHO9u2p2ONowxqfrNTsAjvvtETQiQIzFWwfn/0QeFYRdZeoQYmExvAkQ
re5zarTmnv/ef+J0aXR00Ze8K8qbjjZZ/oCNueBma8TmLTartVuSWBWga1t/jisW
NGSOV+aQpmQhbTKmZvgfUHawEfYicB9yRRRtiJMZ+oqEecZIWIXv9e3cjl1qGsSR
0/0qA4RpHhV/Wko4q90h4iH1pfb19odWRG54/zwCcA6uBVEU+w+aqSCY2/HuYWmR
++NZgPdy9yLj9Cq+eRW+LElZu6qGUbNgA/8rkf3MfFp9gwS72jO/WieyCKdKKKCa
XKRRz3JasUPIA4st//orVRQuj0Prv++m/yq5lXTr7cpI1qjpD3IjCQFWyUopzvVl
65xFH1V+bFPZ7WETqKCX86R9Wikyowas7BCQaWd8FI+oZfoApbVK529JHTw7Wz3/
mzwUwr+Ig/NS3wfCekr8CMXc35H4SwNMjiRtdAqnX9DseqeQYkGuS+3TIlVwY2xx
9oFjZeqy2orVJSPH2skKYbUgedk2dyqbl2eHafQBcxgv3R1GQ16kM+ifPmZbDGAd
Vl57dKMff7at/PBG2ZfoF/4yEL6DUM1iT82nQEMSkhnxPF/cWGplppPkut/RSUka
XCmS5WtZ1RbXGcBLKe14TxtDsQAPsq53vXxkbczGeuv2nmBXLNvAnF6DVi6v9+H2
08Pg3vQnHaVYJjUOx7dwsfdD2TAyZDktotx3mpwWCDftoIAIfghk43MAcniG+iN2
GyYoSUG0P3/rP1CsqM7kPzfj2CKHAVFRiCTOOs9p4NsjLxaT65lspiMmAHRo8AxV
Y+tCARDa10JEG1cBSN9BgQSE4LVGiSYYF6a1woE0DiIQWRZrYzDktZqngZoKaaV3
PJ4reOk0mi5q14iBNymk36igF8swVavLVoDzZ9e0ZZcgHKLONslmqoHtfhGGll71
RBKn0/tC0ES4kW2SmAz690phtfXc1oQ+FxA+x1dCmexfZ0DcUmGYut7GOldZcLXK
PZhCvu3zJRqbJ3zt2uGHD2kD4fQBVRhQht//HC1rz1C7+r5ZqI1bpzmD2RF59hbN
KzjLHZmhPkuYRnSLBa014lzfAOruGU1WhUnuQP0pq+NJchtum/BYi4K8liiyiuM/
F+UTNJJJWuC4p+TepCWrNJzXusXaLxnKxp71AS1twIwTbynehze6YUm4G2mI/XgQ
9L8KS/6/kLeXkYa0TsapYwcVtRcZwtGv/cS5OeAghU5dEBhreoNfjm9omcOU81Yd
95c1/tQ3LPpHR/ERjROdk3T3Zj6OdO4TSqRnLwRY6UnM9CitoUirnKfV7yVOK3ru
VA8kO0HHIAm6/pJUCb5gW6cGUMn6jinvXwxtIgFTeJCTxJNEEc9/cllgkNx0Da7f
iwXmtFXyZp2xBIdVKxXvmUufnri1z0ypnmwrR8Zdin6ntGH3+Kgz60ZwOcuwooAF
S9dznQjOJW4ullCkNkb+HvVx2Ilrw+WSDwWELUjxZ2pPs5JYB+CiSBd9Lb6IZ5xF
ZwgN/I8VW9i5Kmtil1c1gwFDJA7D2gq7AjiBaA/EFNukxl8CywMRDAxlWzPm8mzB
2PYuk97hNGxxGU0+whNlRLbkedVA+sGJ1d7BHq250cPKXbFo5nlsyLcchkSi/ang
3k4ngMdvy8PO2QHTqohPWrYaVmK1PPULhi16vJyOZaAqVLtdKkp+iBFCjpHPzFz4
6KoKZfL14hTEU2/6E9SieYanKev5PupHF7f//pRU876QPdUC1CIDuwWYCIPo3/26
vt9+AqLliJoNrqxq1jDRgZmglDe3MPjyZRpD7htbJMZM1NXCqE+z7N+BJ7i87s3s
55NS5mmtG/I7lQgL8iYgkgH4gEzYtJIPLE9XUhk7KumrGH04oMz40la29sWtX3sx
RDgfpUzbg1K0hYixYAljvc2/QAuCaFGiDbreJzvgkX0delp2JIRzQMOgss/tZdPg
PgIoNSwsNgGNQQpnGtwfIInhIdfGDueWzLaOAT2TonUCV8UwzXut/MBD+RMGDiuq
gglqp0H7V8qwzTqHWekNgH1/R/udlY21PCGybnoryRCHVPu6nmEt3fnDhqM8KbBd
v0V4ziE6TSMj/z9HhlZ6Alua699A0zAX0z0ZE4uUsC1d7cOVgP4PZAkqYqNH8G4A
YogTyXNDOW7TBvHv9Fpn0dLMdnnpciGAwyfE5ZDSBlQwMHpz5gTgZEf7XuJASTLL
BvIEinfaX+QRWyKf+LmzmcdU4TjDcYzVoG4PuUVFVnm5MSsXQ8Kq6Dz9dH8oiPzj
6pPsIVIKuCnHy0BVaLGKWA8kVPQcj/X5OktxKi3kEWcODGxjuuhUfK1JO/HPSIgz
45tIRgLuVex/SlNoBYMRiQd0F0eqcNdNNWpeTeLXRjz8I55MKyBRQpCaD/JMguGo
LtV+uru3COxWPIXbVyPLKMtTv0vghh2vO7DkIK9zfHMQJpLweuOfq1Hn+gYg9/UU
sjJLHTOANIH8SisxjQH2oP/mU4thBIWADsOB0fk/v/0wfVkns81aaONLgiaIioAn
4hRdApj0O0tUDHehMTvhO1we+KQ3ovXptfp1K/QtNCVEb5eIXtM7mM9DsGRjJYv/
sDydi5QUJmGa89+1yIPwBB+kjFrEWHp8navs9NGWIyZ94ECvrkaucUnbXtIEgSfn
/x2Ycg9/qsePv5FbU5FDhiIH6I7rZFG80Gyj+GGhAo5qAsWFcYS9b61MiM5pGNMy
fEnmJiC9NpA1evDEervRjTlfKjXnUjQtVCrT7eHut7WsXDOvDrvs+LTESlJtqt37
YpTwAPMhQtJjyr5AsjOaFaNRKHvVccnexnFlwKFTJydLsXuxH/oXYajnHlpC0+sF
6jt8//ZGRPAI1Za3nYulqnzfdxj/36/tuforwpQtVVPIuKCuqZN1Ke5FuQQwh/Oi
8/gRutQg+JzRYcSqXlDbQwh4e1UtWISt0sOLinOSZZojJPWdW4xaaJnvAV92JeIv
1mARhAbAZ/hohTR8L917DUSC/tf13BDkakNoLHAEI8jgJX7qDIBQqDGSjfIDI7lX
2b0mjyr47PuZRt7CKA5lCvi5cb0Cy8GUJhS0xBUC5A16k59yxjgSxwpGxYfVbG1Y
w8zuCbtkpMYxqS4k4iyMDhHMNzGnePCxQgrrNJta11sOVefLHKzXTirJpt09Ar7Z
G/vQ/3chmnhkxoRLC1go9dgBYJUumkHQS4hEQbwG3bW2IvaJ54EWRcpIsgv2+eej
7AwG0fbzK05XuqielO67HrXFkAhEoegIa+AHZVoeZLH+KCOMf0uW7c6w7Zc31Okp
Ha2V3sZeB3XRT7MhHAnLKN5+gHKBlfJjjIcEY3Odjm9+UqdV5BjPmyCTifkFqC/B
2yi1ZDt/DgjkRij/mLKwhI6ucXoPSHqToAmt34xBJF1uXB1hmj/VDFyR32T0yRqD
Yw54Nmrw2pIygne+5TcyB533F5AajflAcT95kzzhqER6RhUVFBNqabbhxLAG1MmE
gkkAdY2OCY/ZY6Yt/I41yuLknuYATMfyYaLZib3C5I7LaRTIr1gT6yM+VIexalxq
qlS4EeNQ+FoO5pDX5q1bwlo5QO/N2IVJ9XAJMfW0vmFzhxPt0n4p9hI4vNu6J7f3
x6ZDpEzIakOXrz+Jo7+6r4FV5oKaFvZ+UlHVCMP0NjYlyhye+nPcjGrL8fk0veUs
mD4O59ScUhOd8E6AmZ7dIEmFcNVS+zZPVozprrkUDmnHqBsjkYAHstSIa7Gdscri
dHBOATfJfWXuUqll6hPo7HjBLN2GwxUkNGg6UrSrfB+nBUPeGMsGuZ3/dh9tDNqT
JhEGEKw9FQQuACe1gNpA9eQccUTDxZRCQS/ULaea/rTaX2WGTpg2pmi6cHIpvPwC
Vsyp/OKNiMtcS/0qwTodm7Yhv+H5D6kW/23wGBQDgNmQAPvPH1l4Fx9gPfnZL643
aYEJdCAxdUVKKMZdNks2BHncI1y28pJAzuFgWAwqTcpdp0MWSA+xCb8nGETp23Jw
DKCgw9EumwQ75LIiZXevZNpE+xFHLWhMxEfL3BFtQzdEGOjO1IJSZSrWemE+mgqj
w03DIU4azVbK+EGNsrrm/ru+7ePYUmm4yNl3pJeyuhMWbnKoJTMacn8UyxgmXUkr
PsAARQy/keSEyAZTGLBOkDDwwyEA5MJCIHZzp92K4Du7eGm2hcMbBAkF48tFTjf1
5HyLVDG5mLVauE8oGFw1U7zLRcKVjCtcp2SzsYfjzQZaAqP5KJHvbVyyfWTlb/Qj
jHkVToRzxFDhyGfmu8hSJoQ14gApDM3Nxut4ukR3EZtSB43sg7x0ZTDzFPqZEe3c
XH6FNrK2GIHWdyH+QOf5bhSM6s2Ul73Ui9PdHsaanNN1RpXXMk09vjwmobhcyOnI
AG0radPOilX8O0qVXaGGxd5jXo2gAbXPm8CDvOFWnnAhRSn7wFrBfIg/QCrEBhL2
u9hjlOmgxamyXVLLyUlWt9flO0mUn0LB8uyqDBlo2tTYoX4K12tfxHLzJdzApwPM
VTogUkzQTBJfddiyfHhaBpvgv3hM6eDsjyJl/U5UXP7t7Wx5Mrd+FWndWFOc429w
rJpvdbQF41FQEsGdQPeGz26P//9Bl+5GxvDfxkKM8jkpPt/T8bgG/WKZsYDnVJsT
zWuhhFwSIkDd2dqY/ZKAJulU/W1ucBLZ3VKcPT+XLIlYznLg7aYxQYNJqdYAkJWu
lEuF/AgnTpk+L8ruLIva2Sju7BhucUaX8EnJk2tmC/+/0YAazP3+uCIeK9dtvzeg
BShgp94ZwfVXZt/TGQWwHQXuJb63XeTzQ3O99lYAPNEYfEcS+bOZsfNyTyLCK0zH
ismq5N064mGAQ2ATinb1my5/bBiINGAIXFIFcCwfnh3zBaU80K4IaXFV0/wubNt2
5gyyqX0+vbqgsHcZq9nmbNU880yXGx9xqGjn/chWpFKV9vuQ96wkGT2JOZNei66S
65SuEtuw75kuY3fbCqlJxdSvkl0BNCsf2jpM9U4MUUhx+yj1yMbzyqq6CQ3ACEAk
Uo2B9uA6vXMWfSsHFBuVY9xqcfFYMroA1YotdpkyEvgY5VspmOKu/oyG4DUCCKue
BvEXatcCG9zz473jXhIROpeMqUvX9hBwq3kPLAcA7QusYP1mhKcBmy1AKWq9jXNN
QJny4AHKwcbjXZD2YDSGwOT8aPQgN/CAt8xukNC2CgvVushxVHKMu815QO/jH9Or
djEWedtRQys9mHgZB7W/Q6FDAKbp4hBjwlxdorE+4Nhrm1C7fQeGSkV/EqTPW3Cf
EFk02xxqBeIXHZj2Ne7EzVwVE2fW+fHuvLhMigTCOXUxWn7hhjyzo2+lVKrSlhGg
PQo0aIxU5zJzTu1iOVQ6H7q05nTWhdrF6ggIapCOfFTiTFQLn9rS4ATUI/Y/56qM
2Zld7+gScGk+gOfN1y+hhNTBHgalcAylypj7DZG2J2+vfUWbtF9BG3Ig73Ls6SD2
9w7dlbt5lyFWvpjXM2O2kJwIRjEwy1uAn679t1/ynl/grOIyvjVnHlYFOvwE+2Uh
IWM2l/kbqseopwqiGVt4oNqDX/tc5zwHOcFvYx2pCSHyjTSU3cHJ+YYH7EgTNfYu
PDx20QlCOOFzcb1K/Zr7IHHDfbwgqYGzM9vzHHdldlgxNwn1bJf6Sl60Gnd06p2o
cDBkAMqjKq1GmGIU3QmtozHmeqO2fiUB4mZ00n4sZmhQUy4osFiM73ULfk1sn83k
ogaza9SCx95/uHijQiBKIFljPt708GCY2OQWio8b5YqGmtXP7/C7X3hfvKga/iJD
WQaFdFJ0GMrAQHEwOn8gCyK9EY2aQLo62vE5520n7Tjb0eJOK2esBy8Z/GYjlaVN
pRkqDsOB2lH7DDDxBXCxIrEnohPjgqIV9yRX7CwPCiBD3Yoxkgc9LYlptK6mPCba
T+V6xVH+PLIhqoQaM+LGCTzM2LFHdp8QzyHrIH6gOkvjCi3P1Jn+Ci7kPY2q2It2
wlg1x/g6tHqdOcZtbO9oQX1RPyu59UIMrvrpFw8ZGVZmI/dtgTbGjEaCEC0di9Ad
UGVzd+8PL22vI7Lx75toZ/7veES4W+0ABPfU4Q3vG99RAT44DyDty6syv2MuSKrt
LBHusVMfdm+MCdcZ7OqSelv+TMS5G3SbnR4RxSED6W7Bnuv5vjm3aYp7H/u1ghIU
6uJUmvLqaA+XUGB8N7AyYN/QdQvLaEq6lnNN9PrripNlnfqLVYZdEjH65ty1X850
8d2pSNU9joe2sQzRAATo60XfWWSzVJcr+6rpscqjz1bVD7VAtc7vP1Xrwfy0CC0b
URzo+wZOr6fo0NqqQlkCKNCvEFYNr8vTQaS80Kk53LJE4slTOFBZtzd+Wmgu0xD8
Adp1NnA7vIxAoOWG7hoLAzZkVwHIj2dQC6wvGXSK5S59MWoVKilL+QO4BvEyQVj9
IHKOZNXZEmz5Aet95+0GubLxV7wfHr1Ghi4FyIpquL18ZQmy5PN09b7gUM4pxsGP
QZepkzRHAWqyH7zk+XvW4eRPPDm2SPsxmhkBJHnBxQBdf8TsOW9hLe/YiwrLbgnm
9PfRoP7TOFL52SyPFfiWBBCzbYRu0UtRZpWljOKnQ7Fc9B6MCXpKZLVch4b6q8Mp
GfEYaxCGOLjBDLlKn86dmVuj5poTwal5E8MuqR3L3142d40/NprlFV1MEFt99dTL
TOSpVU4MXQBTmyp7OJQJxoCgmNSYufA5nkZtV5vcXIboShyzOAxklPz45r21wv0k
ZmjRNrBSpBxYO3LkS1JayNxwEs9flpaOyfzSV98OceEUqwkQYlZOL44yKPn+iiUi
9pgTwqBnTV4isdf0/dldTYkOQ0jVRiaqKyrMjrEYrQ3aAWqu4Hv5ZtfpSl7Q+1fA
vNPvnRgBwxZY137+op80ELtlYKuc201CokLAKj4UHC6Jv5wPw2CylLINVO9X6X8X
0Wb2oS3BGcmOUNWZE01WZkNCbE8/bF3r4fyNQpcQzhR55ZShO6jRGstL0WdI2Fy+
7cvywpMgc1CivHggnqBr3MDWJNhH0JC+eAmWPrWVKsIPnblNFHr6EB8UCB26oecg
voxsFO+dhK+pbp1M/jXinHObxkbw/EUpeQrYUri/dDhBGh+m2UuolqXKp/c2QjaA
MK++g1R9wGMIGzj2AhB5JTyZ6CNZURt62NdjtjmqKcRUCflkZa7t8rA2Iie9jDg/
HEImc9fl8yBLbXKJqLZ7oH7PUNXoE+eEmu4eOQcRDdsQSJzUfkn0J4z7uwVhJzsf
Ydm6heGhZS5pxM2sQGbCd2KqQWZELxLZ5Lf1YdPRYVHDxxCKRx0EJpLRrWVaceVU
JGFrNey3zuBsqQykzpRmG6Ku9ug6R3V3a1sAnA448QQnCYMia5dYDuK5AX3S1ZuA
UC1leigrPn+mzYMx+aFf/pGkvqeiw1B0u1FnxTBuFgcOg+WLQKAhq8r3OB///YOk
ayHq5h/edH/Dzf53TwJqlGQIrNbY6q3HhksbuEXZBfCsFjocNkNxwMhltyBtxucd
zmeC0K2xEp6sLH4fbwo/9jxJSnndgpyJPH6t3HmXwdXUiG2qp6/p2PSLP+6ZHi0B
oT2vMhAGF6CoJy2MYuLkUMeTq1ROgboGv+Xd/hbgT240z7KzhifTMYFBLYKXEg3h
TduvwiqIkuYIFNTQAX/8WNkWVAq5zQidyQMlBmsNTreE8Lrw2/4SB4gtTor8TZH6
b2SsQsGBX/D5VhD+kf7TXslXAGJg0Rjw0bBzkToV2QLWvgrCq9KUIznhwlctbXUT
onVu4reiK/WO3zkiHSd1oQ63oiYZOZ2yjZqWe5BwVrJ8PpUuP3NgvwPmn29y0kwB
DA56C2jNicgXdEsyiKamArvkwbmafu5h1AXSO+XlsepTRLshu+lwGRRinSaodx+F
UDNZmraL9HOSO41D38Mtq04SyKDGgUeB77pxxAPA+aUa28FGR1q74fdbMPgs4d2o
PQi3+9YoLR6RjKFAr3U+RsnTjPrIKyX/kwzGSE/0nLXUSErrtimAxXgaejRSVVZP
CPkm2JwtFhZ+FYQTjxv2FfSOL1B4Mh8dF3SYu9ziWfbbYeDVLI+2rHeSQ59uyFy5
2T9VtYZbTjbBMxGt3DIW4KQtjs0zsQQPFK+ZAIDrw1DHNom+osLUSsnwo22R+LCm
zPME4DcYjcYqaw/8vO7Db5RlOcFXuD97hmJEhAcrHAccWZJiTq58OaTuTjQ7HCWw
bqrGAuYzBR53LjhWOZf/PnjCmisa2/l0nzhZd9IbrHpsRqv4ejkRMsfH7Vy7i+a5
5Bkg7wRAlCTUjjlyNPVC9sMqTPwycY9+9UGIrAnGPv1nxmAWM6iBOGNipwZAXBhX
+RIqsoYq7TPiKDEQoPia+zRh1CsQ5XF0iCrM1cWr/nJSyqq64Z23dM/Z41i2v3iR
f2SBSTKxyFQq/naf98gv5OVhtjhu7D8i3TMUe3u1VLOmw7pDWMAVXEuBYA81ZJvE
U5EKA22TVIBfjP7F26R4c1+Q8RzPyIdcPuk1jL+IOTxpbh41nyogvFRC/2UjfBJw
FaxhuZGNocb9i2HcHEdYMti0d5L/wr9il60dDo+6fBYdW8WFUE8BW9nF3LiOyCbu
M+D5/HmahaXHEr+cBX+vclrNOLYaZSTUdd8/I1U4Co1+gSPfDWsZUOU5FCrsZNJ/
xoCSsE6QAXitiWJL6rnGzsRZCPUBup/A2OSauF+93TBE4SNwXuU9AOjctzSdpuSd
k8QootPMmQgk0I8rsdlB21tLdphN/6Otv/hiLLKoJSmy1Ur1U7ZR1yetrlR0xbtU
npBtEQDlCN6S5hmEK6/O1MK30gaf1P7z7T/7WetP28AlNqX9sPrNq+LwPeh+7dsJ
pASPw3EnxizjjOlGDFGndK+/RzDJbxSkeuBuR6w9UWwngu8dVInRT+++2EK6kAi0
28DoL7dh2yUtktuu4wTJLnhAOQEKqxy3KLmIH8btdoWrmXIPaXHvBCn2RAhCJ0R6
pB7m5iHfGFPxoRVMKPR3cAP08fK8fGX+llrUi1JC9xhKZM6Lt6gUfFQPBFdhdWIH
t4rKJaxUiny1EmSwcTEiNhBo7wBheZwqciiu1bRnJiz4+QBI7jd2MYVwEZSd9LPS
N2rHZNfSagVhD5RhTWEALT74zd6qro/OMBiE8LL1pIHNhbx4j+LpdGUhNzhyOzL4
rRb1jyLaHzEWo+vAhO7H4S/vJ6S1Sqp6RpdjfdWmhCyMSrfR02sqzEr8YSHRp0jb
fFi7c8d9qWP9nilCWcwmbJzywtG1zrFJUzKeRurFez8Eigk7spwBfdRb+HaTpUbQ
OZ+UYS5lqNzkXi0GwTiDJC+rXvBpoMup9paUIgK4FMFZytQqnmnt890cR/IACbGY
3gVAL075VrXyspKoXNelag1dO3qLOC8GJVHHvUFnmIQ0zNljv7YbGlzt1Q/nDSvZ
1xGPbN7+Wy+dtxhStOYrkoHJ/45vt465mlfEponIlSbftJOpL6nrGqld9K2brjMa
QMyP/KmAl6Xx2/kLAhEff+PfjNaTasneWPGmES2qKxgBBPDtiegF/sT1X8GKJuVA
E8MIR5BUl8HeRli1MvV8s97Om4Zb8wZxaAA/eJEWfVwkNR76x+xvLPdiCMhoyGNX
rSqfIBuqucupeBI0eRn+TilTVfPZ+zdT2nwD4L/fIHaEJl144a/oAs0A2trj22TN
tIH8BSXgbyCMYwwhxbPp2HjwWxk3/gOoPnMRPLblBI7lpYFQ8BcTTrOCmpr5pW2z
r7cjppL8uxUmXbrkHQ33d/WV1O1CXSbWOzQMucYhQHUzYhKJ+p3l/5Kmcqxz+7RU
T8pfjZPJ7q+cXLOZlA8BCBizJkzb1OsE2D1b8jSn+E8dHS9RUCm3fxGsPJgZgQZH
+3vZkli2dVBTdxtGal9ZE8XConwPRd0bCBU6H652qpCOcKirhUq7lBa25QMj/aba
W+E/PlpmJf7KXBWMyam2jVqC5gXq+WwNBumt1Y9HU2t8s0dD7ii7XBITTqXxRp1C
XgV5o6vNeEaNhhxOXRFDJQScf5FI9rsKcBLIIswWMQClfKHoby84QC7WReHjI+Ip
IbgfG05pJxmi685HZvrIpMZlIrxsHIGHtdRcF5kYTYFpedktRWd40ihyDVEJICpS
AzxiJER9XuKMYl3lqptVb2wMALGN0Wc673sECuHxmUXPyuIbexIM3RnxDWuRZo5V
bwvRfIibSL8nw9TM4RNcXulxBJCQdABzaw/YhPpYZWvh19a8c3ER6YYFNZLqUFp2
ZraHowGuXbde71hMP7iNDvr47zOTxNECdWoTWqnD5vC/ZwzmpOEKPWAT1eczsFaC
JyVEZKWsAHyRtFsDLh4SdfM2CPLwvIQKA1ptdw6sDfbRPqw21cwjwJVGRWCNCpWp
frfNxWCz+iZRfxWABG5Fd7cUafZoHfR0PC+/oaMtT5JkE4WLAC6IRLeWaT/+qpVJ
9bMDlD47gZy45fOioRpkbaT3XizrVwFDIEVO/d2YWcDiFGT65zrn/9efl4tf7BuF
MHOC15f2MoFj+tmuScCZy9K7gjpJyynYOO6bsOEd6OG9gV8gjwbBjp7tTQmDwrtg
x4WkdNt2lp9TrqlZ5G+KXo1w6pnEGgzQcrMFrz7dKR2e+mSAEKs1s7IZEPYhwIWH
h2WNyUCMHfn1zz9Gv8j10baMCSkSTvuLu9z4kJ5WOsNHRWDC3VA/BNHm/Oxghx+l
+3v5n2rEI6LQRiy8VaYlKKNyzcJZdSQPq87yzp6piLTfqfVL0+7wrMkelJBSgWqc
655wYH0nwI2ZZZCJ4+0F3DCn3t5dnxDUrLV8xBPqRlyb+sq0sKuYvuqRVJKXRLiI
nZ7mriQMNxAQDVhfLp5YvnKhwfCm8RQiQhzPCje8KSKqzqMMFQE27D+unuOa+pOm
SNqqjKsJoKSWqC5D8Lft382swvzMbiUPf602kf9kWXzClnh9HR3d6Y/G62ceJLPR
MmQSNERPfxLb2R71O3DfCA5hT0qjFdl1kkWzdePSMvdLXwkkEeItgMlnoex85Fe6
Mye2WkwQribg/Z3p8LGBKPbT3bBrLBATZQzwft1buK7xXhoJ82akS8kb8EL4ykPE
FYOS2eACrJQ+VqNsKV5kMfFMu7NwfH3UA2as2ikhyvNEeIRN5gZy2WGbSOG5hqTg
a9lD5rE3M3Zo37Mu11WnRjhKOeCzgwgeFaOq4yW+p3tf3cve98fZFiAXizdlZHMj
3oSVkXT761dlxMNVxoS09WQvZ6phPjW75t0W0BNel7UDTUQuZU4TRdx4DhwLBOkn
6aUkaftcZg/few2kbmxqdQrNk2LyipqsqA+Co14BCG+qJwWzpeTMTYnOCpte1tcU
wgNrJBH+Hbkx13d2qSY3Sgdhp28w5ZxJTe+7bAg1XG+jQ0LNzMbvuvdse5Rd/BXf
6fRJznmWqx8gdu8xWVvapqQs3mLXP1rrvl5/AmlQUGcDhIlEpAMT8EnSl6XoGnMc
+j05LHfpBnaleruWuxhHPSqz8wB0aQmNjjrce/Jz/Vp96GaVXISOawfS0C5Sh8hO
z+/NHH4OLEW3SfCQAQhM9Ix18dQ/YaXAGoxoPYpGAD7QTbz0ieXVB7sBZBWevHAA
m8KoHct55Uhl3WAARYKSyrNf64XKnJyLj2to2pABRXKXgZ4+pjbIL97vIp22HMH7
pFN9unXXcKKsz36SuWd6RYzK38fY2YyeTB/j95fbHZgKyYGOVqufkzNV2e6Ipncp
f40aWuAbGPQwKozRGbGPZRLe9SM7cuaRQ9ROuu7n+/7O/BvN/6czgU686SneH+hM
hG+QIJuqFsLfHqJpGjFQCV2rrKi7o1eM3rC9SfNQ41GWNa5cfG38mal0ZQorZ70R
8LLA8iWcQHxuSCWdvnqULWCbtvrvOP9aUiVMphTA3JFZDCY6SSHv2f0Y0u6RD/k3
Dr1H903KlMmfzITrlPtTud7sdlQpRnvbfLK/a7mcwdyJKp2uM7ZJj1BvKuNbshoA
6maQAKdTTFSUbLDHHHuciPlAOWiGvxvCs2DkY0eEH/xHIUtW4eKCBy+ryhxjsNub
JK07KO5ECcpyu3XKT9bkbMrK1X+s6kbfQZcTxpn7K6VgMbKKqAOltUuFgZ3NLZrx
hzH3gjgJEMjaPqMHCDyp8GCll/AKO0RvENgGoksbRfMmtKjI2vdzZLvGfrWg9Uy/
PPIjNZM1+kYJmmpszsWSMnGcWMsExlTRtyU06pA8A9YmBJ751Ch2EZ9HVzFnX0tK
b80IHVNBjVuw75n5A1462IGwCUJYzGxmP5dcvQs+2W3+pAETniNuQIViHqSt/fGt
Dro+8knPvMi7NUR4RW//yaxkqmBICaNk/uspkunrKf22irnAdvjtbwCahDfH2xEq
gCoAVN4OXo1+3aNGg8gHGgvBW5LTO68x7EeJaycxbxUAHVR7XEfi35ivnaTbUmwY
FuubOCsxBAQq+3UYk4IOgaxKe13+hVcb6w6F3nt0oAB/cjTPi4PyxJ4K7SZ/VMIQ
dTPGBZx0K8DFtnDOd7xqEPSIAy6hFmNUBsFn1MLCfw8pNh/lrc4lOwaBjIxWhLnJ
PxLtARtm3c5Fk46SULRxvR9ApQ+v7aFRPRnYOVXojztkTTb1ZB5D3+9hJgZTIzUF
AmD+CSI6D4smBnOGWuAH8s3bEtcIS27sIvo0tNaexkcRIZW7pEIE5o0fRk0A+8bW
169BWV2SJp9wzGJ0C4oyfjNs6O84gL97yPJvNCTYk7+7K/oI6WmlYiTQsmc8L0cj
hppLP73i08I57U0E+E7lCvhigr0LUn7Fsq8bB5JAkZU3KlMsGtS6qdnD/OIcZwWS
OSdUx4QMaoHckcVM4UWOYoKppjmTr6GmNa/auuKV2e5fb5DO0yW1Vs/uJHHgDCAg
L5kPzRkeGwnbKKkZ1rfuS4znRzC17y3+IiDvA2ureMTr7CCO5MbNFTTap8RNttZq
QgSW7wrcS4svT/KBSnAYlJO/wyNwP5LsZeOy0hOH1erDTCAvZWUIglerwQSGR9vF
iv33Mk6sTVQK+JkGARJ10rRQD3N09GwFcWuDzuDwNwL/4pun/W64k6Yonfzd3PQw
NrX3t9mc7TypG/jbKHC/X9p4rAMjsyb4i+P0aS97Jg3p7DxTYHOIeMBhnJS2adGN
VYZGNm54op26DJlsJe7KwuRV5C4dEvUNR6HwsAY1FCrR1SskjuRCtpc2cHyhzTF3
Ao0AhtZ5Z7GmvicgBbVm9HGFu8h86tEhC/Pwessa+1wvuqCWfHNW6JMDYNs+ZKpk
RJuV72pjPdBPebZXF9Ult/hkSHrPDVQHGm3n2TWSxFwR4IuV6IcFMXx6XZFFSCJe
K3OtBL09KBEQRMfostqg324ztoiZyIH8b0HfsT7tQDh4VYXI2MdS9AignTNHWCfA
HnlyzhXPzsuMihvfDqw1wWocs00otUCBMODV7GE+lyf5mW1aN2S90QdfiDwUfuxa
EyJ5mJSiHgfyRfVK3uDCA+j23FoRHxdigZLPUU7ag1CTTFNMkPSxNyVys4dSh+cN
6Duq3jX7RFgoRU6n1cJAW2M1oDUg31tZ1CnYFWNhR4JiZ9mME4ZV7QpeJQQUMGNt
1iz2bGfxddGpsKq/O4DGTJxSnOclH9iS3vFkOZrr6MSoduoXSYLGKa8P5wWiO9wc
eOu09OpTrAIAIGlkf2Kw8ngSI/kZARol4X7ChLpyW+0IV1VJgqFGTYaM6Jc8KTUg
QGR5UxGBJ61pEPSy3khNDplXPs2exhzsn2b4iOUmEgjeGyYiE5fcwROb/Xvyix75
Bkd8NcD8QPoC0hFP1/H0xTKJLJoBS2E85C2xtrn+KY2bxJGDGNaEK5hlPZs/JEOZ
p6jHgTmy4IyXZURTbliaPkq2oBebcsbp8daiPAyVpl0V4Xd3xqCUYyr/htZ6d8J5
g3UoEXn2oq3aWkWN7xBd7gjNzrtf6FGiEfXbem8XMs4xNvtFCyVJl5koXNlJK8Il
EXrTmlFaHbyzmx+d+pqLuiBHfTZB9zW360BhEJEchFKAf/hGaPl7N12G8DV3pOu6
4vPFRKQQYqraxH+bm7BfcOp9j0ja1y5gxSwQsFMLvQUbH4Wnn1fs0R7vqZdABjeX
2MGVopr7JHxn+0W4gstk55DEDSla8cSJU7ghaXTGB9cGOb762gCHhgbMzIxpSa/6
b4E9xqV89GD+pQXztttSkat9dG4yHwAfZW45YPRUEphow2X7ld1bQFFalFbcgB/A
6nEzbQuVr8hvh8FpbUz8T4DXsqgASYYlLJr14aJqWHquHKb884Pv7iNT5qU7Ve9M
dPhzIJsIUXuws/MFIzN0IACCgapNsdYVptxCgpGuy8nMfskym7PkCJP8Wy56UCnk
yu7Y5cZ0IdBe6nYVeLP0fCx0Bz5004qHdEu0pOsU/JJzY0EBEvGGVkswTzLj5mKl
ivbZh+EwO/YxYXnt3QpPVqR/7K6Nnvz5A9fCJtaGLFY10gbVb4MQ+Ika1nJRxU1x
Cgx57XACpge6RA00cjqwVt/1nx3GgNhtdmUQQp5SGmR3kA8t+LoT8Y+LfUV/8rAn
GCBLtOVFC2fL4PYlDoRsg9jjUfaeFish7sAASPCNYEqi8olhU67KtFaRgtDsnLGM
ONhaREEsXmImq0Bfrq/m06VfVuArstEWQKTBZrUHjbdY/UR2/REn+Ijffm14WIq6
bbTV8fwbhGdk/+LPW4glntjw+myvg5FfWDxXjhHI7PkpvnkNY7SqzapghJaroE7E
bx7DXrKmb7F2bWDBVwFv10PYLiyiMckRlDZNwQpx0NxhMaR2wixiCUXCDIHv/KDH
nwvun/UZ9NuBjdxlFkzgHuu9wwXnG+K4cGhwRwBS+1EM5o1sqkwyoHvp2E93efHQ
cwg5r79TFXuODUmu65Romq/yFGXMwZAyKO0lGKdfjaaljTaquU0OnKsKx8GSjOH2
R20ifG5lS916E9Glz6fanc7xIRfr1M3crPGj5TsexXKe921hX1admEXXp3mHnDpf
WMtwW2ty2/Ar9GEZgyS2OUTkm/aUjX3C0OVTCii3M8ZdwLAXCwLAYBo7EQIir8q0
XBSxsrHKGjbNhQo3Dv/sYDyFgDcIF0PAZSzTBbTZ1viSxSp58khf7gTZkMREZFJ9
MZMJgYfvrWdft/OFktNMwsRX3SNds9WkUKAUBRaLsD93wwPM+D5E6isZn2Y9Sx9q
Rh+3S9/nlBEHvyY5dI6ulR3RHQckEgX3e8d1SC0hOkrapRX/ZN+saB04p9/yf8U9
nxAn9ERwZlufDzsv5qa0bqFAXFl18+ktWF1IPV29G16KCG1g6yidK954VM7L0jdc
/ebxMsONPAqWRTU3rUYU1t/BQEF8k5UJK5vEiA8/ek9Qp3MkrZ0RzTjhJGQ+OmvI
xS6Z3dGI/8f2F/Vlp8Da363l5TueubVYI3pa09h3+OhD05VFzB0UQ3c0UU60C/+m
DyqLE4qiixgAX9OKTY1fhjeJiMKa2BXw+wTtAykAqrUtu6uGKw1OYMdrTpFrzAwO
7iWgV14PmhzxzKjYYRahW8eE9kBsabFwy3ox1fNIcBcXpah7Zk2RaiDYA8V31W1D
vNCgMheihW8JhG5ohBepEEnOkZsrYNyGvVTbsqgoBc/SOdSXQGGRqyq/Qqd0+jCs
UX+hliUCA1IcgPxJueIxj4ers+gm+Om2MSQRae9Pr4ZWaFVSZ5vfaeQyWgmO3ARs
dSOb0SDD6GPAyyirvYYT1QdW74ZAKBSw7XfALPgHmgzpCAIQAkMyljm8G9iBb+HS
TIY3MfZionSeKb3iWrAG3Lh3D0peED2w2n3fmqWWwm7uMBW8vt7zTa9KkBRLeVV3
P0TJpotgyT8ezFoYtFe+yEOSORUTLJDUAeVcew49EEpovL1lAr1+kNAHPahqbOno
hrEBUsMlEkvSal1p7ou1fRI31Nqb5keWHHOyZfed7h9TRd0/07JYQlGlDg3Evw97
ADZmH6e6Sn6kvKwYyrNExhOt5R6/w79Kq43T6M7LO1crB+x7simo+8eEVwHUP8n3
EFLQ5eSmil2Nzc3grHV+7CS++b7PtJkfDM7FkIim19jqpsJ2sKv8KTOHso4GBiwi
x9V+hQNcjY+LH46YKECr44HptAXNoRmgSjm9yJ/9fEr+ksyXVYUbq03t4x4IkuGQ
aDf7cT2rjDC+8cSRPCqF0xyKVJNAfwcshjk9UsUCtALC29//QzGQGBB6vCfBItH8
cQIIafKUztb2ekrX1jkpmlSnANGZ5keVmCz4IMtjJY/68cw+A6seCCU4rE59Cxtw
8/XU7xyknaZp3wMJo/FKyCEiplJiZ4d/KAQ395VnRnDxTRW/pAXCn/mXyW0fw2fo
tlWpQzsyha8RP6/HcIEOGr0WbA19f2dg2kgyxBbwInaajK+N/x5cn2PPIvd8aWLh
ohtnowx45XsqWRZ9nXX5eK+nfzcSP/bG/f66VOR0MFqle2I6P5eYnNz1mhzkZ1a7
V1mVEmDlwrDnqaPpiz845e7gidNGeDVC7ZH2wPujPhWojkkg3TOetlFm7I3dJVg2
0p2zCr5D1GPK3Z97h+pTMh+zu73kAjq1DEnnJeGqLPvDWpAnARbmTtE/88GmuCT0
elglqTNOVZYyZkPsIt3HhvNoTLM+dugXA75vz71kJqGqmZz/DvAMu/jX/oAD43pu
sUCjCKSQfcR989ovazrG4bU5+/TAcH5+2RdWdb9Iv1zkiuuzEMUmswcFv1EVQgFJ
CZHFz/qJ30ediwf7lEd4ha9uQdBBzqmCcXFW+jBZ15bawlBkObtM6npU0GRg68Bj
sZdEkPU6iqdOhlzSLtPCByY/qNlThF2CNs8Nt/uwotQGGvpX8zIRgCNSvlS0XVxV
LH1nmSRjHr6YqPHk4zy6Bknf1WDJQw+TM1cnRnsbEllutVEpRKD5dlyJqklPdIhH
feIuT3p4Gb1+U15sWQ+jJnG8skFOVVJDk25Id+In6oNhI3kx/u0KGZGISg27JoWa
FsNRa2guXp/gGsRNtBPh8CGH3cUX+/gqqZZMnB7lbp83HZD5o4gAdt5gLwto3M6d
dXsG1tCpXHIpOV0JUknjwWeih2ja4a7IUYmP1na4lQsz/xwKP/pvPhQx43yOZzDm
XfRWiGmC9FvJFo0FHXwjEQrZS/XduT0BpMZuGhUEL9vZUtilEektY+SCLzJff5uU
DBopIYvif6VZAYfCQsVvfp4eEIQpzBwvgSaR6asz6T3vUvqq31e6cGhWUTb4gJdQ
FeS34LXLs9OeHSN1hTg3y49BDpobQYKf0FZohoKZM+eLUJbu11K8MaXwZWJikLm3
VK2+wfUTH/S6au9Rw4gT/iMbr16TgO6XnCBklzNK88yZdJdSUcLYfXKnFzdckAxe
G62sd71Kcx+LsCodfz6h8Jt3h71lqLPf7m58LUrHyjMAqIxZJDZ/ruMxGdXbJ5oK
8oDoc2SY3e8myTBukxqolDTIYnkC2bssXvisPCr5c5EtwYXChr47yCz2gLe7Zmcw
E3x70foSfn3gfbAI2Ig4PE3dBtEGWIjkfwDoruN0MyBrfB+aQxUXi/IzVAAVx940
3R8A8Ha5jYv9HPW74giO1ihWx00HghkxSRWUIcN6gfpvChJAw+LsWxsdJ41Rjdsv
1NC9gGdYJoWobXGWsmi6h0T0NJ9tRUNJFtpDDge7Lnbw2Nhs3MGuHb5x6d2fiIF4
ya62eEzpJB0f1zPj60FPtWx9Y48Z+H9dyHohJ2LqkTxsmRtlOho3vj9MQXfnpsZw
6zOUaelFpn5Db6eqj9Xqa7Cip9NjDlJUxBUprKxRDElh2XWVJiSGx54j0+f5c3L5
Y598q4zaey1Yam/HEBEMvvwjaBtgAbX8Eu5CHl5KxVhUgvQ0o8p6Ls/whAFN72UH
2uuH90cYc7DQNfz//Ce26Uvm2wszLuR6ZFkiQ9w82PkR2q4bIikxB0Xq4dB2ZbRC
j2T9uaVEDYVn3W/3QSo3yMwKtispvUwJJVD/ykkxpSzBn9MZlnv8aIfXzSrSSTHl
KrNhJwVuSD4cq8uNkX9JeLG2G80rcBg2JAPpnBcuTv9Xi2dWM6JG9omfntzcnMjg
BNZKId7Dm1N7aB9FFTrjhmz52Da/pVwDj8Yj0JE9Jptni8r3eWsutOwZdLviLX1R
QHognXPVGxzQiRZOfQ3v+cKpkCzCLgZR8ebZ+ALuWkgEDyleQM+TRuUvTr/3zO7S
QmVhGkofDPAY5Rhwmj3MwRpy9sNteEmEwEnsRrKioHcZfRSuQsFVCQvWLeftEYhN
OkD7idMNrzoCX19pfL02FccwnMdlohdrv7PSiXpj4VARnaudJMdfpq/lSSNtKZGY
wuZ++oGDHDybibgqtZqZTgh7Pxn3+bDu5JELCFVQpF7NC5ZgIuv5cNucVqoIUTra
sUhnBg82SCjIClBFBU2LBR/vhiq7Oot2LWCRZ1T7ODzOiBtLMlkJhWsEpBtjTdWl
KtGiNefNcW6tt0TuANtaj0AAvTTvab1yHxfIwiUAqkseMT3RaUz7/3PkeJENeWxv
eeEpx+lBESiflCHVtwdDtMbsaKcJNQGexHpQYpIJsR328ozjk9sxkefFcRBlw/69
n7NHx5B2iqtJCd9Jg7LEjefaLiPnn+VogHDqhrZit2eVzhOLzdwS1kLXd9bvPNuy
gGxBkjb2vWU9HqqMkeA97XP/QH18gbw/S25O5PKbIVDnbqocOEQTMX7UK+Xemz/J
Psk7tt3sQcarAuvSfdtCjSmZ69wLaUKEB6wgYXNleJq+1p7+pnGE1gbAcpPBkM3Q
EGhCNN4LuWemdB4GwHi/6acINahopLbN7l7Lnvd6ReO/ND7967oCPedz3iENGxBF
MqUlopbhZc45dIGYVQaAD3dsDf1TNZZCHeliFFsIUeA+QUAwKpy53B9UcQ1dA8tK
vr1D1q6FNhzW8urj9QOpmoLLQ+IilA+unwrL/jIY2F85trV5B5xshceAjO8ILXFH
vFiIAKMnrspQCvb/Ew7P60BTWouw2hPJYLYmyzkKdMSEPimWVX0U01sXwA0G2vOd
C3tiJZ3L4Dt6CjsZHvGOngcK9OwbtWDt6tdMF+FRqozLEwIwvMVzsCE4kT/Vl4dK
EpIsYNtzDfaoAerXM2rJYkgsVvQFS/qAvkKs4cZqodMcK3a6UkdYc+FPrOVHsd45
afbZhyxEktMjiTOb9GJkizw5nfqr0TmkpGm5d2wmv7uJbiKwty8Lx9SnKgK2a9FP
2QsiJnxskxwRgteBl9wm5nGaggIlkhD+5Kdyno6KndR4lXDeziqvVu7Ir0HERagd
7od8MmVAXcw0oJYNaa6/S+XKJpST1eslyBfcuHzy+BWvSATNDzwxsJhcXsgicmll
e/0EAy828wZxQhwKsr3wkm/njXqXjcKH+D+IUdfe/RPhbvdBEx4QbNyfsCcSvHU4
VwU0YMpC471S0jdPhr4/G2gWi3mKlA6ZXSrrQr9gfw2bOH2AatVOOShJqXN65fZ/
a95YfbWTPxR1l+Y89xV+Cpfeqk81bpR0EtQe4I5MK9wyqc4/5qo83OVu26fBYMMH
y3mMBJR9pQgxEYqRctKPtf4W0Bho01QdYdPR7a9aAnfLMV3yz6H7DNE9g03YTWHG
M3zPEvQkjIdFUt/zJ6+YbI2gqUz0/CxM09Xsv6MWV4FtYVvo8UoCCbXoJ2DbVHpz
lss0u9XdzzCcpdAsfTOps4GJMzKtlIGzI6irmcrqz1Ty+o+9gUx/upRGbfq3qdDj
XLyjY9d45t8BIobUKCHoArPhiIppz3RB+sxccPejh8avqU0o3maOTbO7gL0m0Jn0
u0SHDvx9B1MKXOpPyCIYgd+83PJ74gp/WeSElWKWmZoanZLA3F9ORiSAhZ+q7Zw/
ozhG2s08Bs3ryjyNm9qDviFGIqtWWJLV5tdC8hRwC05dWN0sE47Xpcn+cpjFj34r
1nahwfaYcY5HZPGf3MgMpvO+erqHTLsHZCCV9rlNPwby4Saa41dH3eNjJVIGaYqX
FbnY4EH9RSHU9K6WBmabqky5wCS0PzSHYeoDA0PE4SEzDYiQhammVIaXPeB2Czjq
hToMLxWjTfw46JL/0BjMpjUGhVY1oOc8ZVwLaVU3j1G2jWBdFS0qvaYYO/F1TJQX
85dK6QPDD8XJ8bHYvb3s6oUx5m6eOr1WHl06acyUCrxX47QmaCn0xPUIwpPYsZcL
EIIvazV/KOZZuOFTptq7XJYh3GMGQzaWYPgSG5CN6efXUYkY27fozTv5EqhloVbT
csuLw29VRrB7qkjOSlgR+qPULuGieYKPgEfMe+NU0e3AT0AiFyGokiPjzWoESuLP
BctiTxu4gPs1LRqVVetnu0FM8qo1UIN5IcOx4xjFjixni6tbuJNzqw4rZA99oLDQ
l5nMnVTHhviAID4Kqb0B9tgfOEpH4561SGMhZc1oVLVeUqypNW9jStVK03f61AWB
LyJU8q/0ge9rdLKU2yGZD8xJQTKPssjA1Qm0v0rIygjOPNjtAKjWRVunPTlGvCAr
KjLtLx1GXT7DXHswxdFfzO9wwO4uvBBkcpPi3U3E5XLGcEP2YE8tO1AKXoKnrX5R
ffyN+77DxVTsHM3yguIItHMw0dPvt2ImcQPAQcE93qNxnrDLrp2OgjmdkMjOLWMw
Had1fSY1fqQQfo1RLT3FdrwIvqDpF162rba6rAq9HSxdCkgJjn5lR1SQ5kYYnC9D
rlArWKHw7konLYQVeHwLzuLXlnXKDM4IKLmRBNywQ5qYu/oQsc2goaE6bRKPpHWl
rnxRQwn4h7hsQpcvtVKCfo5W1qMDI/eLzadMmpLqEACp8giyTIB+twvfI1OxAr67
Ld7mvyWZc1QXtH9KbS/07ZiSMavfmwQL8RePTkbV3HrAHu2fYb2NugYWTPq9Io8F
8gC8+F9cPzFlWM+LTX7G1hQMu2W3/CYm2qWyxrAg6udsQFmT51z+hQsAtLK6a36z
nQoB/A2w9l70/IIrYI17QysQFfaTWWP6YSYp5AaL/4p2rD+m7voCWz+923s2RXfh
JyAuzj8z3ubEwZQolz3NA/RslJYuV65QITcRWWcyh6PYt84beD7EGAHe2PWsN+Ty
TsA4r3/l1sPcK4RnxWeFeWxA+sGtftIdpVlBnMJPKOS98J9Q3AZb+vpa/H8/5awA
OGK5BMEj65VJumjftLJkXTtfycXuE/+LtZSUGYQg4JALikhIWH5pw5mvNnlqQoz0
Mwgn7QytgNH1EleLDLKC2beAiQ/ukosuMXAdS3y3+NGdso1fuuAXiLiwHLT15y1f
qsv0OqQLl90EyU2TQm3SbvKxfhwKyWATq5QgY21n4m6T3tjcA/qIaYT+NMTSvKqZ
NYnc7s4W4lH3RojS5sdLYII5Bfs0fyL2x0PjwQrvaFPBUN1sEhsKt9DZIwPqtTCD
qsrbqfgjUWqNu7HpnjMfccJt2hhSl8FugcbtVPRW8iefuBzjdjM/e6YHEPpL9byB
gwwyb2W4OI+nRXlZ+F8WvUZ5tmEySx/evi7yTt/dlCXpjXtcru+AnCynuuUsKZBB
VxZkCpaZ/sYHedLX49prRWqasjkG5hUhWrBG6Ay6ipyi7USznV0aNTL2twttIkNA
JvNoRjq+RXqiuJuM/LA6mwZdLGnM15mq3TCmxmoMKSr7zjfEbVBBcxoBDHtzIj1Y
O2G7hVvNmDz/KCanblC2BvXcrGf5rdSfXy9H7BzKqQ4TZ52OUhjzh82h1RqsB+tc
19to1h2urpXJaJKUBk1k0TAyoBr96XvSXzQljXlvM76uVcfBSd0UZmltCJujckCk
4iCTzoOwKwzAWLigZuzMY6Q8qSoi7OvKFr9MM9LF2FLB1S4MpGUpFPG8JAkm3SUG
mwtmprybIXXLVFlKeKW5o7mrid6D5Dy2fTZSnkid82LNAdsDk4hIiKBo3FJzHnzo
dIiEQFU/n5Rbt8DcNWHkQFuMjKqt8tK2M+p6gsfPI8myHP3lb8ACiwhor2IJiXKX
/tfEUGR03QQX+Ct112bZ1tdF98P4iM9eXV4hpwrYlv6K1rcPUy8LLaDP92lcwwvf
4QTOM+FnCcb9IrOjEAVU16RTKvXj3rqIsidgGOCGT5tpqQLKYrwC71eekuZGshOb
Mau28pm1XMXKNPJcKJvayCKgAAYxRrJ8W+S0CfSvUW361gjt7ERHijeJDco5V0w4
YvdqUcuXDxpoVKnSbsDjsyZ7rmKe0aG7XmiC2dtsr+YwJRHXhiVN2jchLON4nm6N
eSJzg6oCc8CvULRpEJ2muuROnBAVC3Y+yD4ld5sZV3fAJqFLyUEN/2uf/IVcd+0+
rekp4ydR+Ozod3en+p0vKYvuFQdlOoOX4iiZv7FizO4i/OTLMf/LDfXBBXAHrzeH
ES3sxoOfvP6wHVmOolBYFrAV+Rb84yZxGaeHQVHGs83TRNdL0s2mvawq6wUdW7M7
MGZFhj8jiCBoHWkg5/kCaf3EEH8FtKIwJSp5CTOYzAosXJC8/2zPymPXCb/nCs9P
tA9x2IrL/jebo03GmPEbKqJd9kvOuVwjgEA54MbBUIM39LdGhMPK29UCcSYmZeGg
bNyXrSo1tx2PHgoiMwqj+Bao9ywnlBjuetWuMa3FBAwQBqbWxMODJ0ut2cy+dN1Z
sjzeZtj0jSJl+aIgp8bqCrymA9edelViZ5e1odbgnsNIq3MhmpAMB6o3Lv2+zKEY
r8iwDxgS9B8E4GVR2vykdh1gclMR+YQbY20Kse17IJUKkaXTeq8jlaJTaCzB21LY
QC1Y29cg/Zotm0sMWNVBiPxFQOLDhnVhKbtmWIVB/hshRLn9KfJrBzvw0mQEPL9i
oOqcuIv/Y+wX7gR0+7MoIDyBW5MfhAggBpwrw9dXD36xI7nrf6VX1fXJqNPbZpGv
9kEYSElNyL7PD3VjomPyKjtQW0vvNTzexo5Y+7OWR0ZYFDsWMhyOHfet7FyKygKi
lnjAne4J/67dGeRrX0VFgnY6d0RTLZoA+dc4L4DNdIyXwKZHEKmTfze5v/DIsQ4v
g+LrAfBpqvssnsslM98TV/rGNHZ/WbdcT1LOhK6r013zbWmKP5KHlsNG63s0sfqZ
xM/l2m5dbW0fFeRBI8xqqp6Nr1jSryrWAtPrLLsvAuZdqjGgbArJXETkX7kL1KzK
womYmMzjnw3Nkf1rz1HUdIyxuBOKt++wK6Xi4n5LGxIV76HbTenRTI3ljCCvQ2Pd
7wzk2tDm9Lf/Suh/vihrid3ElbUzt82oBB5FlYKdKRD5c7LgZaMO6DVb5mfcYhHd
Kx5d0jbfg8K2B46WcMqCfe55NsKjVXPFBsNnklfiM3mgvaQCtEUPgFLGKP77BXgA
BaGC8EtbFvNkFqb2t1oGQk7YXfo6dSHMytTXzqiTmNR24FjJz2eoFcFNjsk4Xhi/
9WBwrZvV3nSzJ4XARcWGtBajEOS+XX+5ejrCdNgPPlzWwCx64kODkm7ZiQDp4T5h
Yjzm4UAJxaTGA01Gbust2Jt3Opq01qnD6DeWU9jnWShdKkjegW1gqzgMSL/3v6UW
VwdBp5BtjSs/iQyW5Cy1WSMlYmBf/YYXrf+0NFXWWU0WJBcTvW4qOLaONJMmVKai
R+2UfK8dQaF6N8nMf5p9bYzFPSGNfx/m/9k67TWTsXY5MBnUO6GJjAvf8XhHk328
htmKErA81a2TFe1XVLJ06IbyqEfjW0SErRKGg3HvGYPIFbyEVmOlOfVAld/I87Vh
iR4f/FOfbcxxLszaxXsakHVakxs/OhYgYhU12yaGd/2MbBwyLK7loIc3yi4MdmcO
ZjkER7tu/B2HQaaGd3E7l87FHXazrECs1WKNRJJ50laVvkS1hCdnp+DzaUhvUdJV
5z80MEjHnLna8iPxu+MD1RXqz8RNXZUNPDLNueFGqe57or3hOxR+712hjiozsoSs
0aP9EVmTG/MECB8hP+dWSDfDxzfoUoPKzzRwFCtIjh/yO93aqGgoYSSn9qacRmcx
BWqVfySso1NH7iq+MXEmtlvirHDwEReDhN5pHd/8rS+K9kFYzYF9Y3i+XNFxb5cH
29pNH0UIxl3t5bFW7AqyFCw/dubxbJ4Nd6WIP1feJOD9PidTub2bgRlpnSxluauo
fkHY9AK0iYUrK7R2ugHnAYgwF7U3/u5IXd4J/RMBVGWcU2OoaXCJxT6I2lhMZ3Ib
L9ealwSfUfLK2xewCScn5inImcQs4HlhJNxbfcAG7f9idpahem+Lp8hrQM3OHUw9
vXzC900f4yuuqziQ6I8qj6Aaudv/w+auKiRlAvJrc+STHhJ7YJjigKz3x1nLVOHn
`pragma protect end_protected
