// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:33:36 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
dRelzmCccKXU9l0+S5Fgqs0eURfQdloKxPjy2pP84bD9H1hrClaPUZbGLqdKDfWg
51UjCPbpiusg63D+SjGS1J19fTnMFv6DuZpPsAzDmUCkDkayzJ1rZj71UEcMubJ1
6KIHRNamdQlfRvf9X1FMGhRD2vnF/MOhUz4xQ24kCOI=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 7648)
d6HhiCuiWFHM2NO1LH4MJWilHK/UImHiCDOQW4hYIWuBoVVwJXzjmb559/9+TUlH
5UyB8RtMGzkBKx0bjFaYmQ4c1GNimuy4xBfhbTLYuT6HOKQqJA9z6nIEpARl5Dku
k/iEDhquvTpuac/e4Q6qvoKHu5tPW6Z6f8vlUXbeWrf7xyRMBVk+j+Pr4owJZbEM
WRXgjl0UM1SzMkz+gDUd0fL88YNcOpjDmWONJqx6QdinfGep5m8itAGBnNAYJe3C
uiukBAVQXYQfzlv19OCp1spBDkgUS2UcLnpMdzOIzznd0RHQ0ZussqkLdt1O/bfS
kw/LupCGZuYa7e3ICdcEu7LzXsCiDrv42xGsQY3ifLGV6ZsdQ8zzfuB/4EGHY0RV
jU6FF7kxdEhQPr75g5l/ZYEAk0DPxJtRAFkbik7I+7P7UaTSOjiNjeLPGTro9IlP
5Po+zvtemWlgsS15oVYNC8dmQAeji48kF36+Aj5+VhmZWmrGfvPHqDatRIEg/APB
jpLd/zi9Hr1KzmbjU0LED5FGER4jdtpIBNVVaoxprJPsgu+O2+WCmkD4/odN2FBC
nen37z3ULpg9oEpqIKViWxhAOqcgVFnwk/w+QG3GmaQsX2qMdbnf6v6CDMpJ1QGh
I600aGOznGScjvpVJuuUIrNwgNZtTySLwf43WsMvRSJPKHKR/xUykkjaawzJCFkT
SVNOtts/aUZs67HeIujeS+3f16CXLZESOUp+WGI/2DchHaz4z9J4Gfnu22b//x+s
kdPXV6UJcXkvwnrtQyOeareHPm7p1+7+kpwXkV30ZswOJJZQsuTndPFqNsn+uXpJ
4SxMln9cx3BSF/31lS665JbD0n+J1nFUQ+sycR+Bdr6iwND2Vdvah1qBPn3h+70G
PWoZL8nOnchNchx1QYIKnvjvTVWpXEI8xyPdPM2CLYMjkpAlUTO8PBjGfPfyE62g
j4o7UgjYFgdQWVqL7TIu1manIzIr5oAbmuhRG+G8O2pfcIZ1SQ9EORlDzuuG4L3H
jKUpZHDixJktfCQL+oPFxkI6wQ0BesYlcLOCRE3ozZJ5+6S0OBUU5rZGbfaYdDq6
JI0EPGRb8XZvm+l0TdxgQm5Pyyuzzm/qpBsDwpogq+YviE1EQ3Pq/IDDiS7ZbZzc
0SEUb7c8KAk9sI/hPc6FZ9E5cyATk70Jq3BMvR6Mn1rV3s+0B5VprEkGP7vr8Svu
9oTOMDJIkVNdCh4wuBci00HM96e/xVMCihcg0fIupX9mcq26eCFkHH2xXErQFxAk
hvfd5xSobOraTVsFvrHq2QnEvoT/a1+aqowxp2wUbKxGP9Eleqgj3wQ8cgXNRQxa
NyELaClFBnBmcP4Q7N09VpHZB9cUeMfLxvEALaZZWkSGonInuC1k1Mc5Wk0pS1Fd
fkyeGS/bljnZCz2NhkFQpIRMp8IN+kF+fSuhYNM0sjXQKq3pb2+5LItfo6qp1bUt
gp3g/2o63Jq7fiur1XjZ6ztZEDxQYwiR7L1P6N8kq+WjgJxPmnk0J51W8/axtvy+
xmCNJT6LRFFMyblZuaQpN+dTPBD/19gHEhH4MvXrQSKuaEHnO+t4XErWs6ByVe12
GY1FWDgfG0rwhh6rshp9okWLnlbZB+pkHmIX0m48e6U1YW1hNA/XnkD8q4LIZ3xK
bCC/9UlgNnsIqlC86WJ71ivstj4OK9Kc5ddAjrApYrscIKS201Sop1QJkUzZDYsj
aUBa+vfW5WpEpnOb5XXPOlNXJlf5qvb5VzgdY+QNYk6y/Koc6YNu+zub0UpBjB2b
0jRRqh6QLuhPPRZVHVYh/zBPRR3ARCPUkBPwAYhhO653GNPHnH29IxCTkTz9RdV7
lEqx0tAO30QurXEmrT/fckGw3wsSLsA7G/JVKFgZDOy1dirqBXh1BeWwFDn5bvLA
MLMi8yuT7gt50EETepkAv3P0KbUTwil1sG69TonZ1gDyLO7BhoHSpHjRhoG9PYiM
c43OetWoFX3WI9TS37ryfW7hmE6sVKxBdJZ2e8Nf8axOmbVXycOknMdQ4DigQTh3
DBz8U0bEFZtU1pdcvmzjw76q3ioUAXUgJSaYQSfkosJCo5VG+U/Mc6bSfm3X/x5m
U3WDhVkvM6GMGORy29z1xLaORCxTw7dTXhcj7VxWKL/jRb2wr1oE3AxsUnwOeZuh
wVebq4imVpgD3yYyAAhvdcY+HMHytn0cJkqbLcnnK91Kt1EKuo74HlGe8gzElEor
Hx+llwh+CtyrUGAj9yNPdA0JHvNKIh6ZKmeJQe/+S4m8FW1zkWQP9nXGW0ZIVbyb
UgxyX5wjfzEkMLC5ctNL5ck+e7VyUNbNVGV5ar0XmkifyMBJvtmhV2ROOTZOO410
AQON3UURGAXy+RHfjS6l8N5DWsjEwbQhmvUbe37YjhuSzUBKGLqN1yqGPMviIgro
P5y/8bqQpi99iQdbbmVNQvT3FwrFuw/BDnWfJL/mXhOlBVll812Our41dHUSt6Dr
+VtN7NfZs1hpFr+A4kNNX8MD0LqzF8zwljc3mu5s2mspvGX7MDsUcGtlttf3LebJ
ne+ROWhLmalgzy404AkQSE20P2eUmKL0L0fcPwO4+N92IrNTBLpnYnQ1uh+hIsm4
c/l1DykQCo43NOS4ayXYTuuJ+DOha2b4b/EET8hcaYn0+0XkhFRVX+u1VcuHj87p
hWSh0vizCrCDMDsOQYd7TfgQBGJqqwr4lXQZbtCCclW08MjoMkBP695QkBhkLBEd
kS511cVrUXfoh9dcplMeULNqhLYHYy54MLqStR7HmIMiQJor7TEvlk0nh0t9OLDg
evK8dd3buwbL9JaChuAj8l8kKfc4zoLgDTY75BDMzG7eGNCa+JBuCsLXs1+aGeMR
L9QLrfv7yyS7XT6Oh8FCAwzHVVUe5CdenrqzosyVLhNZRIf5D2hMWmdF/RZiDQ5A
N1BnMLmEWE1TScimxIe84l5LAjWGo/U0PzeeLXgSTadNi53DeTj4FIPxSJ2L79qV
xNg08q1j52MXHqS7jqv6HWwnaIFCy1m7N/EwXWxfCPx1hPz+Yksgk7JdDsS16p+N
Yfhm2O6X5KoZImY+w6ToWO+2dbsZ5XQ8NYcrCCGtpq/scA0GK4H+14nidrAoTRpL
FTpidfjPc/SP9jESVzwkYvWS5iHM5qW8/A93t3eTHt9YXgLKSWVHy/rpVLpoqiHp
LbAxXNN15Uph6z0Z3NYP83mqcE7ksmNq80Oi7KwtW/SSQMg6Ep7gK2LU/6gKdp+V
1Reko/MAkgxK/D6+I+pgQT8eoTXPFS4pYn5SmbLHgOoxN4UldCJvdgoP7BqvpUIQ
q0wAwM7mFEBYttiu3LM6UyUkn029sucb5HQ2b/PN6r1X6LiEvW3Au4pKZ+u9v8ji
El+xxlll1qtjtrJa/SXT4Yik8aWwHcrbG8AwzgfaKdH/sfb0MY4HuXWjvtmKqetD
BgOWrOO+oscjK4VF04Sw4727J0P7VGCen9wtYrk6x9Y/T96X5SdA3SONEnMJSSNr
fOYQPWS+TjCJo4cSVSoRNTzKPiG4fX1gylTHg20i3Lh3ckY/cNJ/Mz7q5KKCm2zQ
1NuuKoKgcAlPp4Hd+X7b2IWV4KzzbXvsklyK6ekdnKtBlkS2pWLPYNidRgOvzDDK
bArbK6xo3heNcLSXQLZaRAF2HM+0WwKASTCUI4iGjmCq2rdNsxTR+y9aeE5Dfvun
oKeilzWeHrjNxD/XK31gNp5OESCf2jgDVFgiV4PlghHl80JhLML509shuVOwuS4j
SCz35l1p+pW56j6W0b56c8gbaVJs7UCvzvgRUK83Zalji5Qn1p93FA3796ngq7l1
tnJ4Th1IFmptK42pTszXD5hucVmIebNHpbkgvi92fOsbJZjuNZVfIZjYm3WeWgPG
AKAaLEQNUgdwrmp0cJoxgmAUEPtg5IhmQyq5/kR6FCZlQzOYb5hds+Yrdh5+sr9x
MXQbPHdgN5LjzLri6eNdHCm7WoqvM6bWjP9DYkT+ulfjaOdNMm02wvYXvCi7gQR0
sG9935P56l9chZ9ULT39sIu/zu8NpTi8l8RoyfLyn1GZ2Zue3uei0GTaHxw5Xyzj
hhimyATk0TT2AEUiTpuznTRdY3RKXiDaEYOcSbnl/uejXkeP3IbxvTk1tP+JjbTm
6sKpl5i8OICqvHf0v4UtB1p+0ePCWTAn04TKcoLq1vhhpKunNFAhDN0hiilvHj2C
GKbWNW9Ska8j/HNrDjNIabbpUba0A3WWIt1tR1RKuu8U4HGbrGXCV8Ko3oe2B3Gj
jll9Z5oEosJtVsiMOVkeFO7DYWNA3E94NmLlaCRGo/e5BRb593KudryMq5MspFcl
YDznwnczG02m83Cbqvdv+Z7l7ZbeJuUq69keFN1I8S9N4qBO7c+badLWjKbi683V
TDoCc2WlKIv1MxZVEY/6ucHWy7EoZhnTu52uCs7Xe+8zZUpCHHbGct4SRjp6tiOK
DsObc01USPQqY/0RqTG50XrRh690sjoIFK0NvOMJcF66L3CkEzl1aW8bfdK+ixGi
bFWPqYJcTcHSBHgmmcZzfySQxIXIyRzqL247KMQh7reA6wdXXwjL2D+3f9jZG+hq
pEgi2noYc0DWUBdHpxiWO1Mqwej0B5YfrP0x5a4ZZWzAPHSb9o4mvGPyWVm19w9e
p/WaguWCmZin6nlbU18P1us4hAi8YXH2ZbeIsfTPsl1HNiQ+EiZVqqlOhhgArvu3
0di4WArs/TICTN0kaeuSEeNQ4YolUICvf5wbglw2e1/hjDlZjbFWte1clcRNPPvq
BI0ENOUquatd0MI0UieNKWn2ZVaSh3JFbspXvPVBlRduhWx4JGb/1NELJWL9zSjY
igPbV/9rHblUe3iBojZ+KZZQJjz6mkKiiA/vbyXHD0qupaXW9zUVtaka0YxSTItt
6XCeLmuBn5ttNN/G7g/0xzCkgtuXxk5aewC6KtUdMvpXbC+Sh9cZxrrDYOsl/AN8
W4s8K+6iXtoIosFVJ/qZX82VwdOrD5PJ1HwlAo1wEBV9j6l7e+6a8MH1BIWi/wU1
t3JRCtlGfK/VHnDZ1hbh9bJyO3BEke/YtcmYt9r+zezYZudF6VvdY1odSrE4zEJ6
W2i4gdVGGJbqo15YsPTWXRU0VCqO7pOXVbJF6aXsTOeMu5EfscMIwccmwe9nY5AB
L9uX0f6sJsWmqfyeDPN58NMS3iUU9BZvZtBLFJEw57ZyuxYNRNyHMIgb5yImRQjp
I3w9NQ28+LvmllTKy0hjh8LB374fIhzdMy4zi30jNObhhq1v0tX67CxzYre9Qi6U
PMe44BusH9QLjEsYpwDM7Oau71yy2ohKOBijxUy17p66WyDFwLBnXM5LImjdwxa4
fmQbubcoWxQAQJZuRWm99OAorhcEHuCjNkyT7x+c77iyHsKbf2a12UfRnetIwU+W
f4WDdI1oGvHL4ekGcqW3OcrqSNRtLv9vXFqIPSgy5A3GE//7lecJRs8dPOUO9jJX
taatR+nKbIcIa61iWF6rMMLF82b0WsqG5O8QWwrUUu++60NfQyTUBnDZ1F4IL10s
Wk3LdpJiwmpAUvkvzniTQM4i2GiPDQGvnopaz3+5en9y2ZoAy2/n14cVk1UQLDF/
MZCvM730sQS7Bzv+dhbsAsjDXuhCo0cDpzndme9jL+y0OToIDSnx+r6CGhpNkZzj
XDFDapdcsUChdoASwCjosoU0/5PPmX2kk9/eHsCEutjwF7ZZoKWMFQd7BlubYImd
kRlz7LfgrWl6OQVFy1AvXIiSIh/9EFkVyYiEF8ml13DaCVGBmvkYx9Gd3QI5G0h+
QzQKJL+Jn+0jpzVv7j3Qe8uyMPytWPHIdg5Xs0IMlbvNmLfrPp7NRBXjAe+JLiCN
Y2G3k/Un6xXH686LFPR4mGuWkeeWA1TnbBmJRudE+tYGxA0NAH3ABP5BrVJr/EPh
4DRX/VjcvleGZpDhQaaTTlqquVHADTxkxoXJ1OAkjs5dMMaObyQttqWcBgdJf5d2
+wRAqh0VzCZr5HnL8AWTWTCTfSNQYP1UdCxSullf0PrJJNmqjesb/CF+uNaMJBp6
kGsaeIdfWFXhpooQYWmcJeaH5DwDBS+nup/+HXYQtdDHIdcQevNTpevB5XmE6VK4
ipqD2WZDrP1AUnj8yqlZAS9YJE3c1qnOwzFt07GUQZuxMoEVp+S3LHOhfMGPVREq
UD7EqqZV+YNnfGH5POaepHO5dhEr/tSEnI5xkJW5QL20202S1ipivTlFIlIHw2g5
LHszRFICrYeidhoLHyQGKqIdJKjDh4e0RZfzByjuRJNbi80SN3B6R49HBDIDku/3
Hpgw1mt3GXs1BI8J9V9LF5T2TQAaQbvKciB6jCxdNHY5F5TJDxHAHE09bfZyOPly
o2ubW6GHXrqL8WXT1FYu9LF+B1Mvf2rRkUwQuGokzzqaUGwTqd1BierxqurwPZpf
Y6E69sZZaKVGRU6Yhh1xBivXUdKRVtlQ3SfPM2FOA0wdemBouO3YyolMyhGYdQHO
2MLuG82mEp4AXCFBGULEM733jtxZWc3mHxmyEGlTdcNzvA4J8MwE60NBgtejjTKE
c30v5Iir81avSXjv0K7T/mZyIxb1iqlsq7ZlgRr4SNFoJglLW2SVHLNfLpuiyahq
+s3s3mz+mkbKzu5cwUFVNgKzmpoK4p3XzJjSl3l5L0VE+9luTWeJmBTl7g48qnq5
fdtI5pbt5NU521tM3E4XOGb/bHZycBk9X+6C5RVKn6ok5q7lYpqi3J/dKlAQdbzS
ZSXukrpayFWXeML8lc0su//21iKVblVoltR9pyytrWSX6Vad9IJ/4HupNd5lKlaC
S5GltXwzqUovphFyiPFOeRcFl+bfhLSKiTfejiNVf2o0ozt2R6CfFTuk7xTIOyIM
v4aNWb1LBJxfvF8rkkn4veKyS0yei6tDEjCAoGsVRzw6STqJ2A2mz7L2qCSkueco
Fu2pcgczQAE4POMls7eE3s6J2dAzFJlJ/Mqv4hG1Xna3cq8cQaVCgavu+Dvg7K9S
+BZyVCPyc59MzTQxkudjxo/q//N0d+mfO9RNeXSg94hKzLwVTnJZaze70GYfAS57
lukvz6/OyRpJ/mnWl+2Ow6V71Rea22RJkkvbs+5TVRbDTkVMeV4c551Ho8uhWYeH
eQRSB27OJWuwSWPuF8mRVPJ4qwUJzqOuKIptOHQZdCDecRjfujbWt9UNXOL3Yk33
pVfjXfEYwFwbRPkEnt7xndGUaVKIXsbhgQYPdGfbZzGrkfVThiuMeQkh2NOas6Hx
zn9/4wEeSSZ1LjUrjytZHUcjNsmn/7eXuNLco9Ccrhz77wCSkBhJ/zWSshfYGA6A
bTJmX9oHfg1YjQJF32WBG7l4I2s2S95AdXOvCYqyWWkLimgOl+ovFy3E8wheayFr
iT4b3LnLr40t+uL1RIdBLi1b80Z5FocxjGZSh0Sb63fVlXJRW6KsZYuFFPgOeypa
Y0kny2gyjiJGfdTgXlVlZ6GK+WMuta6VaohqDEQDRWgj8yIrnqoogAyCu8ZdH+sl
wZTtcU1rdGt3FYBGWMnDs0hzDbDOOOXXwntVRbeGlG3uPBREGjj7qYePpPzWu/6B
p097T5m5/aHrLbQz3ZJJs+oa8fBLk0uMSxZoQLocm9bkprA1ow7FA9ujNkLZ5oFJ
PJe7/gl4E+fgHyqOVXGubowJEO2xAFpTDg2t2xFdnxURtMIW1lDrG+++4M2jGXqA
0nuvNwduDEc0tMzctpcDUO6FdW6v1hCBl31FjntP9XaNC9ETseixp+8S9tlo7wUx
evpfsQNSO5LzLqz4VYnxuTKjQnVl98cXx51cTEWdGzjzdpGu6/XElGmdQeAsdurL
bnnoNTAMUwZzqe+Kz+CH+AbJzPSVofgYAeSMtKC0Ahg977UAGpTAJ+8rkHnlD8Dd
ktH0vX8AzZ+F/3JcpQlAczBvmJPmIkzLJj3azdF3bL/P+wA3/qwpyb3Wno0q2Blj
IppQ4EN6z83E5rYj/j72+PWQGhkcH6tLvL9mgXl495EuQOr49b1Derx248cRhbtd
4LBJkdEbZ5ZqAUqR6imXa1opvruiZwhq69Pg20ZAZZ3BU79SADJRIQwddoDPTZ8H
WWS2W9O1h/6pxDgPfVofw0sLWUUZHcmd27GZgFdKsMogY5cDPDLdyBbbrfuUtHtK
xwpbNY5uvcOIiM0Q9wMzH0Qu+c4rjPSNutyftlDkz7yjlU/PRVhyyY0SSYHKXYR3
aBLaLqlmO9Eu2AidSDRTFWdUOI9nWL/SkzZi5WAUXjxs8yBqsNtKJi1AGLUczhj5
817s9VaeeF107/hCyulb5Eh2xkzV+T8F/YX38+y4ts5G96myTxJ+hYRDrOzjIlPK
bqYdaSrU+KUe8PyjdwiUOv2wVohy5mQ6PszSFM5lm38zb3n9ulZQ5c9t5sPZQjhO
9x+1vuQywhFljvdjL3etz6c6qjIObEBQQRewHroOuoPF57DJ7qRDtzE4HF67Y4hh
mtAgeA9631Fvv6XrhyORRrZVjAlrVusPHqWuUIyCZdOr3asZsmlrrsZ40wCbN+Fn
vYbBhZUxMajPu88JftT3qLwK258wlkwPVg86dQ7zC89czcu6SaqVIdgG26C9+TtL
S68EMaM3i7kNuqRB0m9teUHkQcHcD/KKtrTUHpTrKg1JBhh2rGZ9+PubcmrEz6wl
8ksIAyeLCb27b3DSsyshthE+glR6WleFGV7HAyrVoS8o/cwsUMhB2t53QIYgRyf3
8ZK0TZdPkXcxNHLoZuiFv0WuLyZFQxrOhcV04IfKkpv3wPjCq12JpGePmW9xjcen
/ynAAYcXzfrRHeTWwKxZalakpg/tSoWl+YOQssbtR/jFkg/YdJCXeQ6KMYSYRnY9
+lQqzWeN8pcQdRw+KZd1b2WaqrnJA0NvTQ3sFN7HxYY0v4FnzNNQ0w/7Ttnmj9BC
E5XTkG1HjouGWAxo9qdGnFGQmRyKFe9yQuBnSzdxgGRC2r7OfhZyI1jGho+e38kU
vWeQXq7NvPR22WOC9T7aVbmMRBc+Fy5HuzxSHFSyYF2kbkJamFSNKnBDsYH+36BR
OVvr4EmYUqZ5gni/o9+YaOJFwDim5yOOd1gys6k59bKX71MUN40PYMD7iSj/myDI
ePA22G9AbqoBD0BgQI31BZHL1xv6h5DYUbGOgKLriO1H7Pn3ic9OZ8Zj78ACjoq3
rh6S8LZfE3rLnkj6bqDQNJw0m6vFvF0DxXWkGj1kDAwFdjW+vlsaiZUG2UNxswke
0IugyHzb3FVThzfuJ0t0H2HFVw84hKpplxjy77W4yi8Znmg8DPyNlAZwygrZ5+oH
hDk21BgPsqO+N15ksMxrb4Mdzfsm/2nSBJC3K12/2RXALzq1GsiO3PMQFKa+7VQr
eZTn0xFzzbKUIhauEfzgdQSBmb7a5xh3t4JZezs/5WAbk0+vyIB7X6OHcMbFpsau
GwSaRPLFlsom17CqMZjr8zCMNQArMcuMN4kYJcnx5EPWQVZXEsYI/fYvq+dgRo42
srBz1tEbB9Obm6rZpxgaJ2KKiFVXqeF3YBvCWVTYSxOLRb6YaB/jbWNf+lvtl4d4
CB65Rwe62Yry45FHKMJ0hoRb5ZksEowORajSdpP4xqUiIIz7Vm/JQa6Moe715ZF9
ifgiWEg+Io6OYlCsjw+omVVYnSo95aZsEa/cFDPTsqlU0qvUI3zVI+g4NajcyoVT
0TehocrH4yz6Ldurus3BsstkaSw0psMuIyRowgq8mLiYCECOGRkJO9wf6L7ZGYgo
X26ZILzdPPSOSYb196GkCj9/XXqiKUuweIbmTjX4glArJnu3chJtpkLRZEouO8sx
UuK3cK/KkZkTkxWCNj0S5R+4zWY6yH3+rngXIr7qpZXnVO7QpF9RwfEsK0tP3qCL
0UARzEtuWzYNAn6kc6EVXQv/YZMjP2jZB+JHCBp0464d9hiF9dkPOFkuHJetsaic
mMZEi4L00bK5sakFFFDJUtismohqnWU8dRVIHTwhOCI1aIwIr2E9BIJ9p1Xz2HUo
w8nVMeXtNCYowQWwD0snrq1u/LWUu9AgOCNJ+5Dazqdj8c7yRLlSeJkJwARScMiD
sYM7isv2bfxtIEzHKUb+U4aD85bTMwchLvKYGyfVczfbSx4jS/VAerITE75Omtxi
C2kdVCcpkAtipNWFuqLkrQ==
`pragma protect end_protected
