// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:37:16 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
KpGw8cUx5iijLUtATDfNz4BIgxlFG36Hs7Y8Zv8marsddsnDQJHpNIWY/dGOAe/E
j98YbXVD6U7742wZDuf2sh5pEfu15UMMIM2pgOdF/do32pt1gmFhZk6cU7lsDN4d
g3kCFPcG5aTc/UHm8wxV5sLMuw0q0TKpexyLLJ/QcC4=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 6432)
yAJjZV7W4h+La5naCHrp/JXgqhO6GHMCNYwdCC3Oa5U6cnLzia8oyT1NqngnQY4U
BNp9/COI9qKjmV+hRdyeEyg/5v0AfaEADNJXU9dn0JeOjSZD/UDH6/M5yjm6ECe3
bgRbzJL+CscsVmb5k4IXLUvi+p2+vIxs3nAEkR/QljX/0AorB52MMvFCQsEBoarh
MWajCSasOaM7J/v3webrF0J0+/R3LOPrNt+p0RgDacKhqOr0/iNJ/DcVUJBas2gw
L0tueA/aqYvN0WHkkOvZGqhrcwcXsATqz4TtS9D9boLGSvM4o6YxDphnccfZwiAd
o371EvVzuVCl7XpmGDtq9FqlunOgW6hunpwpZZQeP33aa0XszvpBY9jfmT4hxPxr
EdsrT6q5ytO+FjUd1XL9s7eAq2VKX7vBqQIrwwJ4BcWlFU8v7x6Mh/H4sC2dzqFe
KCEnKWaCBoMvT/M6HjsJynDUPX8N+zYLZ0ZAKVifRQPXxFVSe1o7CIR8qsUxcFrH
LbVGM1F3jD8KzOMmtwl1gMaqETz+QLoW2ore3i+VH+gPs536bgW8Qas3098gAu03
bqD+g4pd6AXAiRYQmsXgvMWHlxNfdCnX16eMELRtv83+12rxQAVZf8pRaAfMpn7F
8KSBbjJXdt1c54QOsHqr8d3jqlkpMO4bXsLxK5cK2PUqPGLPMERRDH76vZJbWTe1
Z004V1IT0dBQKD9DXTzA4XVOMDqffdAsjc6TimPp4h18bSayfwjqgH6cw3dMBYYl
4m2AaBbE99I9Ozsstos5Yq2mGqgV8oirNYtIHoTt9ifWvRlwxGt6+6s2E7SUuB7d
5/o1+1qS3H8Z2s35ARzQ/6KnKsUjDR5hrpfk/2GIJctQenVipA+jW9fVgovWFgfh
y9cxv9E2ZlioFjSKU2pl2+SaDtH/uwFvzGfKifPft2Tdf245LKr3enJ2J5rNYdoY
p9BqWAR35c1qQ+I/qvNfu7o35d2f8ZGizIjFNwdquP9CcXkQyyqdXb0ApBV31M2J
c8/qhekZjxXF0mGkGh/Yh+n+V0mPnlexd4wqiSJ/g27znKh4c+YFb85nyWzfvCeC
PL+b5XM9qnv7Epv2R8sYbIx4HwOQ8UZbQrary7D8q4j+PDIhhJXFMY8xSJZ1sUCM
8tpYiK4mDg4QAv2DLjI9S+2Ygz6wOzUjdh9RWyGj8CH5TWu5affbZpctjpU1MwxT
a9zsAs17HhPvByVBa+z2NtRfZPoIqMx9m35Q4QD+8biAVDGapfyQGq4r3LWSMIzp
5qmmyA7HTw4OXjsuZhSIOXS0Dg7u4GAVWx10jGXQvz22nNFl9eowzO0k55UVJ8DT
7sywmDpd0EXVXgafK900m59miJ1NBTc6QzzjzgPe03ip32AKTcy4OExPCfMNK/MD
ueXAR0U31MvYW+a6LtR3sSk48BXwsK3+b/4CcwhDxcY5x8uxO90Yi9R1I6ek+3Qj
NnFxVu++we3g92Wb3zdH1GZYetPuZ91WRMWq5uk+mdJxKs2mYBWIB07GioDWXvHe
1F8h4PmRD+9wZH4ahATE998l1f7lbgaZtOwrGdM8lTdmbYO1Fx+PkhEG+n3mSWu2
f786FPMt2zhw4cIW1umaACfJxO+am/EZGW2D8HhRrmRDBiz+IIyB2dlZNF531NZm
482vCwSm67qkJ3kuRMYzFCKeIswDEfBaBa8fen1Yn/kQYQHQJswi6AYN96JJwWOE
MfI8BmhLWjWdGj6TQ98KkCwUPxLK7V1MxXGCuyXvJMcBKRQxo81XJ8KSe1JpKsKI
VvhkQLY4OBRwsOojWgzK/AjQuoYuyqgvYj5B9pDluuRAoQSAubyLbSPBrPPBDE4S
PDmAjd5eVEwgWVglzhNy1MTshHVP1M3r6XJlWF0q2VbcHa8vLspRlmIHZLJt8s3P
a2F8NB1HXegBBnTgRWQ7P0HbXOYfHVCNVh53Hw6FzPzDk1Ab5qari2KFtKKwErfV
MKFvqxSYjtAEz8xun/WDY8vc+aq6FzvwnAZRbZTMuCM37cIP2codNb8kNOWR8U8u
njrHrgq5Ge1X5qbcE4znrZqsIbTYTMQFbfYjoRekTK77DqGh3zmaLhTSnr4W7aKF
jmFJAIRHu4R+2LmEuI9ZFZSgrZ6I9VBi8teYpctqqp1agCNipMgMBs2NLmZVnEEw
0wOlG8FTsjVdBJPr5WSUnsixYAIK0R3gsOPyLZ0FxffQ0n+8D6oSfo838I09JPwm
lQbUaVckr7oOrJ2CP9Zv3f/x6zCNnS8anJwCtPjNoQUlBfsM4C51GoWYYV48ElVc
llUqMr+vFDEo9pr+OI+faPGVRatYaUL/Cwru9wodk8VarNKwWl336RJe6SXRLfPy
suucnJDfSDLi5cj3vRSVhdxYJYIeLC2y4wWkBDSBkDaO4RuorpJYudHPxBl04uyh
r7UOTE8X30AguhwH6DS2xQ4gCaXyk4yXiij6+6zlUuqmwaTf7WRpzg/W1jtMNCIS
jfjjw7baoq+djazda34YFkukk50iSjumAfarArfmn9O/wiUBoT9r05pYRU30bHuL
axu1kwgVieoOPOTDPn2V39NK7afbYo+xNbUUgVdIa43Muu62+A6r/LQkba/Uwd0Y
kH60+VbXPyk7Ww9AmrXtiY7XWIBqQxH4ZP+sFoiEcPxyfVYcxCmbxdUj7c3Y9Fi2
EgwTpoyKobvIpqMVe0VblxXzjh7d8fRzvyP4dFs88+WnPgSpDQ8RD8XycvJ7J/DL
p+zZIsUilw3trHk+T5aarmthzuUz/KtOsrBxGiVODLkUi/28N8jT1e32gDfUOjGY
9DWhQ6hTbr7JLTvwiT3l5g7Z3PDpDwXXoA0f98MtZqR8UO3HzgEVMDn/HWTZ3eO+
Wl8ZaIbBx3pCDZMAfA5Hzd8IUwNm1/7NB3Mo1fJix5YO+IrplP3Gq2lCOddku4yz
LIvir7meVHQxoDxzDk9Q03OH2SZMrdGB8rC4nVnYsppudoY/dHGXs3VBOr//96+n
Ds+YOFZq+95Gr/rt6WC/KvyPagi88cCM8HmdNdOUmAsSVVkpCJegVaQopyDyAowu
FE9pB1SKCOWq0qJCBnRZRwHAb+BokBJLbx7cP7RTo90NWaKkNk5r3tPQRosDul9k
sg9w+C1kuDS+TH8MJf7sYZ78RRw9mXQ6GefFcNT8Ywrl3dGuXIBnXcFVYyqrI84i
0kd094LhWg/bc2U0T55OPKVliiibXl+z48CjTK2cq7U3/aeLlq+MMur+p5HOs/Gb
OKCH295On/z54w30tX+3SivDi+MwVSYHhUmZS9DwjcB6LHbP2wU/2X3DSLWe82Fd
nwP719d8eG7vPYjR+SP+1eVx8HmPkQVcDQj+EycUv3JoSn6KXkRu/FuXXm2uUxkJ
YhGmFsRp/pykx/D1mr7CcWvEQ5YnYYy6x63macbniQmHNSj0eJGbUTYbteAI3Yog
FNq+4039z6QXaKI3VHuQGvmZL2n3IBdL1SDN/shGII4huOXiVY1bjyFZvKbR754d
Se16G/f3ltYYtHxw4RNQPJNGEqpDYxcGRYQjTu03jMVe8agk88kpWbi91i5oq3R/
qy4rkxJPRXf6yKgO6BKaMZjcxOVmwoUNs//z9R2noBXA51RZvglQVxR4GmZlj+GV
pvcB0jjRaPw+Fp21qpY+Jm5HfpDB57+v943MDTBVtGlWdA2bFzoBbz1YhJwhvTP/
+aIhC/Alwnkz6vUnHiBemz5kbIRrQxqWVPZARPWeoCIFS5nSEKxeAZeieKJuZTc+
3DKXzp+RjYCRQYg3ne/ChJv8+yMyPcSzw1Jlo6VzMqsZt+Q4U7nDyMB7uL//XOSY
PQ+yV6GrWzmDoSQdOtzmGUB+UuOjWJxCjXLvjiBFpG1X5oUpXz98U2vwOWobDLj4
MwsInXYGi47DKDrjNiBIHYQTlK3HLZHOQXulLaA6epoNzkmLh3Pdf1FQVb7qbEaH
QuIBRhEOkSfx/nUJwf2gxO1mmP2ucQI1rRbg9YMlrzkHtsdgo22CwwnoYEcVxhPN
KoaL6D6UW0bJ85D8g0BVwzc7rBnzyGm+1Rz7grN7nEEQB4Dp+JSlUQdavpIhP6sN
soPrrTYVhRS0UYD5fD3pt6sl9NMSmfndZ4kC88QaoVloVOEENiw2zykzTEjUFBzk
59v3WUcvwturvpweAB6hVZUclsXQu8LGltKAjZWZmlGrYX0Fcx7VK32EvkdgmMVb
wpd8XU5lHWxvFwmOcd3iec7WWlOFJLU3+H21CkUjkGpFwCBww/5Mb+AmEEH84IXt
eWSvEZ3Wm1S5SfxnhgxOGVosQsznbLOwgK/q9oz9Y54HIMhasO0wfk/q+lYbO2zm
yGkO9lHfoZO5ZRXDX8zvqJl1ye43lmsWrIOqDuB3oXjWA+G3kqjikMAs3aOoJBHv
E+Dm985jvHFEE9ayRSyfFJkod1eR3BQqavJQsElHUn58fyN3p8IWAiwACHJgMckJ
Zze4EENl3F1Qfko1o99EdkShN3QJlkF6Cuo9E4ukeQBXW/RligwHKg1hqZkgOZ8R
gjctbyNUxJImvJrxTjcU2NV+uBVYv5uV0sCABUfCHqMp6hTrb6jGeta8WB7/I86G
UuR/kSUJkVlLlUb7s856UWjm42PeLiT5iNiixIGjx6PwG35Gd+D2jv+e+8zLiUA+
OK/qKbyzk8zmsqRR7tOczO1pYBKAmI5whdFd5lQ3qCfRr2NslM5TTgnyrP40SttU
7ZPnwn51ry+yj1okVQHN52HVTdB+z+YkTP/ohpiYZScZetrpoayUh5T+nQ7Y1W0p
Y7DF/8VlGlEA6xeZ7FqmyAI93eMD8uXH6GZn8r2pEkoN354ECK5XsUnaTLcrIS53
dZBxBbYTAIIs0qdCeI/GGwEMME1WGntBtssAoyXOWICa4Sn7OEbInQHyERNoj0cY
l/w/ulFgSem6snNTQmLWAkKtbkXks9cF6eM1A6c5xA4oGhMBsUF5+w2pwbYImKu2
nqGt8WrmbJ2c6RYFBgYKNonu3VyKS/4xNXXIiHZdGdQjjy2ps4MSh0vMFmhyzSAx
igNaZmqUjnEx6yfmpfRTwMtdG2a9VvRbgBF+f2n5cjdRYxHG7v+sbuq5mZtihaV5
SkA/CQXh5CBFQh3dXLba48pxbUuS2pbZgyq8ENC5fkAEYeTKyrSI258tVy/iA9dk
sd9QnEHaKTvjdmquTjjQxgL2K3ntpFbaADDmmP8E1j5AnfJvWCaXOzeXKCIGZoI4
Kwza951kbjo8VvGqUuUssw2MmQNItQ6Cc9eP/AGIulFLzCRS9eikduCgnSjUUjOr
uZwBAZocUSM5boY9GymvyU+787YQ5NILF6CCOypRSHlAhovbeCZdcMQHVfFH6tFe
ZbpXVzua9ytBcn/A9w9kVxgaOUMli0lv/uKQ9Q9oKk/U802oGmmQR2dtIC951qoi
a31Ni/K7SLQEozWtvJkH4cF+rXEnzv1KRyLp9umNVwdX5CgoxzhyjBTM+jyl+s63
5XB7gBAoasx4/Y673/sDl8tjQGI7Cn7rVmai8z/K+7yiQ7OabwDF/gFgq7k08CnS
azQfdVtwyDXVZTy1m2ZfQKLYnjKdZUnCKzvmyCahYgADDct1JDw8NNiSKvtcfs2M
85DuPQaP6+l1QuuGj4DmAp+CztohGTdGmubBI6sQOM4zAZPtr41FrSvUBkaT+Onr
jxcRATNm6U/ER6jIQNuNN+60W1UKhktbdeYcE3kTxqyrprJK5RRaWlqvX/qneSsc
ckj26b9rF3VnWu0qEObOWQ7eIJe3CMsvnDMhOEevNcHg+o2yA02Rq+pVs3ZXspMu
nP4wa/cAVQw1B14zsZ7v6Gy9Q5/VM/zYqxG2lK56f10y9awnRA6VVl796bdQI4Du
je2IFDXmmoSQg03mPq4rDPqhmjjldxCJnhGoNyGhqziH2m4ETMpc4wSK04/Rkvt9
G4T6Y45slWmcmhUlHTJ2F0K/TS4jtQv/NckI+hcI4h0UzQZcoX1lvxfSihqYsi7F
/TQkfVxCyafbXYb5znczy85E/r/CFTwYamUb0hUuknE+1kOAfrhEM6Vpcx7oU51u
oEF5ZTihurbVzT3l883lx6TpH9BM248Ea3Zgg+269WTcf7BUKRMXZMyz3eX9kYq1
Dddtcth4AAT/lyyF6xYLC03oBUCmLY3uGYBVhtgb47gQTqehZiYbQKEQFjgrcqFQ
+oHMjYzH/qXpw/E5q/kUSfn0uHs5ugHyKj3s3GlV7rEvftSl6ZU0RWIJAprALu2y
gRJYTggizO0Gvz6hM34vcdUsMPolx0b6MCmPKCX914muK3hdkfeJ0c7jjuXbjLvx
5qePoRRr5F8FjXHzTt6D7QYPVFWFZoSUC8dG1i/IFHzmH9s0ksCBIAup2GBPrgdM
kh0lCJ0AsmvyzaSwsVvrIC41XiHkXl+Z1xiGGUDAzB8UFkcCa51rPkQ+RMrwZryE
Mhg+qNttsYB3VC/CeRscTRRlBU5NurUa1dn3pJ2PTA859a7RiroixgZ6mWgPXXW6
xVQcJh2F6d2oDKyCFgwMyfQ6blkP4/z4jKW9kr2LJN2DveeUwUXLedDWhUg4IR3q
hLU0yfRj3suXmU0P+t1hTW76ZkT2xV7marhNeR9X66OBk1rkHRp1xgnCvz/v1jcT
TlXodl1dbfpvW9o7ZZko5D1sVBtEyTSOKJf7wklW5CUtwjv2CVu7GN/wJi4BhE8r
SJ1sCaYyVXF3EJKeXUrI6lY12bgdQVSQgFVl1cWLgR2TA0d4AB9xIys0pQcSv7ny
JZOGRL5T4wZhkJG6c8it80yIQQs+lje/8gxvvhu78lGwFp+wJk3siq+PgUpF0fqD
2DpYznZRUztkHc46IsRmbLZaDTf86yNCYlihr3n4VniL6pfhyVR+eoCKgirzMb8R
BwRCCG2U/m1Xqpv/AYD4WUZ61kiCt8fiu3uqcJ7VoQPoFUUk0n8NqMSQ9rY7r8t1
4/6eI0MHLGxa1zMeq76AZwv5ne3cPqdg/aTm8DeUB5EmhvXGSwosoMusUHNcGJj0
Zr2NL1uzlfOscs8Bc8W8vDPzu9tG1RZPW2XyQJ+IpWYIhpX9R4hse8VOp54DgguH
ADq7dKu9Ec+W8uE4ImnuIA/xq+ersLgMQm9wa1+Jbqjw5Q1Tas5KmRl1pPZE/1tJ
pPd26CwWG7eI7nwjyoBLkilmlqWYs6TFN6N9neyeYdEoUZpt3/14yw/rk7ZWFHen
pcJtJXfD+1KDpWzDHR3JexGoRY4TJA/4vUitOFTtqKGYA/dTJr4mBK9vscs1fe++
/v38qLoR+SJkrcR0CBifa0Tyh1xgsV0DX2qedfoH6Y6dvGlM93VtTceQcwNdjOk4
H/ffN4vqqqmZqj+97ySaWZdSjsEXCgJ3G0uXBiCxcgs/gsCOD7iNZo5Ea85vBVRT
b8SqwU0WFgsk2aOwTa+JAaqEAwYiGT6WItKsXaJNVbgReXtpFxSPqT40aAkG50vF
OgwLuUsjVPx99r6bNQh1HteJVbqVDyr+1iRAYmRnHpcLF67u/8F3gXz4vCZhPLCd
258b4F7z2uSYRFoOniWhYAK+HD9FZzBoKvjkhvW5wbyHmVn3MTEbO0br664yw3DK
ku6+I8JZijtwnosucWv2S8vz/5Qmif4VIxV6NAP8JjJ2Qo4Ttu37ANRk2WVWN9Jz
UEZWEd8q3dvu2dd2hdfFUTrwr4ViulTuMiU+ntV6gBUB90EbSyS4DM+pADnpREX1
mY4SyCMW0JlTxTaUvQEuxaoz8kepp7aEhMDV/lOm+2KaLpaQawDimBINuh5KPtgF
2lIi2dT/hBGrvR/FmG4biFDIN5J56MVzWoEZizjfjuxMxqFtQetS0ZCvoULh+4eJ
U/yLDmcbfsSrHYah7ugDpGfV9AAWateQ7wX1gOL8TTETbshYoVpgfXmzhvpHQVAV
alVT+MclqBav3356deZ6vGkdLZtqbgBYPKBhz9f7FRlCXA2caLmPMyoAlHTM+zdd
zcrDTsaCnGQs0ywwOgD4AxNJo1ie72x1hDb2U/X6NkO+d+kTKl00KX2mGktb6Ji7
No9F8zA+ZtirUMkMTz/YwkCpMBJWCRlaUt/8GY9XPjUAaTIHxOCnVjnhoYQRBHQZ
gLzN6EW0C+vCJClYlBhzJBOXyQyo/w8hiSsjYmrnZEU0im4aECIE3GUaF8Iij/Km
3GyFH8Du+fmo7BJvyJb3GsQXvJpS+LwwHNoObNSebG71bwbvr/FAswPmW94NZh5S
a6q+rvOAMyXF751mYudjT1/7ccOnsmGB6ZMN6TwfKEd6x9YxjHQavHPqoxOErE/y
9KXIMaETfJqYHZyac/ksPHymxYYMoxFHYpM/R+5QY21ds7JPLnaxa1ihshXLSb/P
6unRQd8Bzh+WfIYGAHup7CVTH8eE9vfm4Y6y6twAU4D8Ohl82QuS+5l5MvKuw7zc
lBT6eCAlCHP63L4PB7faYHsPmjqQdjJEngh5oTmqHKOBETQvU77d7EwGOJzdcaWr
XYPvQpgGqV38vxzW5/GCSlSXea4coP0+DUm3Kxw712JLFo/NYoKJdtLS5X2cvOwL
`pragma protect end_protected
