// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:34 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
cQTGX3mWstgZC+ENvRtWbXksRogBa2LXRuS4vHCWfWjZD9sHaJCPQ7FeaFfSfrcy
RhDVAMu/FpdkBx2ju2FUkANfdyoIHLcHMMNN4GBli9Q4bRtuBgtZiYjk8QTeiVTD
d/lcxUi6oybo0JlXjR8QyXfnC/0jVxL9UjnJRj3zACY=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 34064)
qmqHgxOJNHfvaj/aladU4+u4pFBDtd6CK2zX3pTr18ozBtHMe08vMI2dmGN3L1la
gURyRaiBsBuW/LcyNbb8ZaVSlJn1j9u7b8EMcaV2cSGSXfE0DexH3Gi0ovDWc+vC
TkjTp/xvAWJyUiBAslLKkypFG8L4hlx8fK6oJQH9Ara/6f+R7dGQy8PiVqFWDeF0
1F9HdlU7sHAO7x/VK1/6kqtoTH1eyq/cBKDCWDDjfOhlhALdL0vzZb9z8k3jxsR1
fVtGQ+LXu4WABptMhja9C9a93abez4Oky0ffbJUenIrS+MvvjdGmXgR00hHd8tKd
RmFuMv6VgXwFdoBiRhPKYMTapS1I1tXwyU1C4pnievyn+dPAkjwDnsYK+fbEq7bj
CWOsLx+9mfqoWWkAGfaxBrYxZyeY49k0fzYHu8f/H4M3VGg6lJ+1vmD0Akeaw9MR
gqbGYQgw6mbn1BAGV+g7PC5dgkS/oUKgZPz8wVEEvpw39FK3+At5iXyKGc2fHl1b
woe8PVNKUyHw6CiqbYs3NYH1FJQ1KcXY7RQCN8TVto4Oil2cAUUb3fYwGm3LniIk
jHfsMvamyCF584HaAzLCQeGut/2rRFjNtNc/VcmhjdhpqsUHSb9x5/VBE0ZujamH
4e5KcfqtPd2BUQz/B313tHmWyeRFRlvCrknUAoI/LSXE0KHWvbwLaYuqhiDugIWP
BvuGJaO05oBM9tLaLY5o5s7xI4rNaMQlz6qOcDKX+mize0DhcIma9bS9ogUonB+Z
kZPISMiITW+GZwh94AFFXAteE7fjMK4dez0eFKlqK6oG1hKcF3wnQJbHjjuGt0et
Fd9MXES9FQhrBdo+/+A8XHsqF6fpVWW/C+NYy0X4uTY8NZOuWv+BxKL/BUVYE643
kgsPJQ1vl8nfC+kfC1iacGukNU2ZjU0oGmBY2Acp605eo9Wvv+AZa5z8rYmUObpi
rlBHtTq+ZoyBkq7nkGtn/pnHCZX3ZwI44ERzUyn4UOTXbI0nAzJTNFezFrW6YgZZ
q2kE30lg5vQooutf55lOaEuGFcHfl2pFC8IyLZiYIEK7WaJlbamlz+fbVFveagCj
9AFViegY1QANrL1FzbR4FuDr3aPIV0pJNehxbxkwbXUaJfjC64KeK5TSBbiPV+G3
wxVoM0JaUSSI6tMS5uX8b/hdkirTpoIJ1pVZUuOXzs3dDPy+Lbs+jPUyxaTaZFK4
tK4ukxvTFt/xyEfFbvEzJyl7DIB5p5V7Mkgn1xWDrOtUgIVJA+oljBHr07MxQLld
KpoSY+nDfmZC1AnfUpRX3d4FvhPcGRvlCOOJ/c3QkublG0gBiL5knirgD3zo53bV
qr1Yl3TyrZCC6Sgbgyun8/aYjy8LP4LR1zAT5vyVChzUn5s+oH4XS9jyzE4tDuKy
Ddg2eVXdgJ8kmam16B99WtBhDYQHYslGKIvjNn6i9R6LwnuZOyKMaq0b2v0Ooqjn
miOX981RX2HrY/KqJG++OA8aG03C+rvU1rzfYaQx34slZBviXOxt883sfLKj3lsP
yjdWp7fyLumrgLLxOA8mJkxa2iOqYuaO1CWotk9619r5OQheAdfQTGoRPGCLEQ7m
5X6El3Q8ACgF/qdnvZQ21NxbeuEu+uRgPPogmOjElJdT+YJ0228ktwfT8sp/5wB/
aaMJiYI2s3Xkwwtk9A/yN5vrSZqKDVyLPPkJ13v/o2NFPtAYs+FmFOlHq0xcchgh
nxBFi91FV56MEOe/yxgonz3Dt4bZADI28ltbTQYsjRinIQekLRMLyNrtRs77OZb7
N44upi341ZyQf/CYegkIuTYZ2/EHE9TMOy+5s2DW6zoFJIgV05wI+e0Vd5IpJUnF
4jA3JPSdXbapYCls+rMb9hCFujxLa2cs54syGPUoPF8hz1jfZNIA0oNZAvCSzsb3
dBWWFs/8Epn0oobU4YYqM2O5Se3oOJ+fxTDFjDF8uJ3i25LihLQe5IiDCxTaqsqK
OotmNtywDQvNCLJkEUZW1yl4dbOp/fiBicguTNj2TeHbwn8cy2WUeH9ipZwJGFzB
izikdjeOWlEvFZFXMZOXUX8ec/2sWpg74vYO26ND2G5ghKEmpoPp0ItgI75Bz0Ik
DMS69BJRrNadXm9AySvBj4T7xkxkwMgV74zWuoXMEC57OjGdwvJqKKIH8UEz93Ul
DRJpV6Cs/LQ51Cw7pRzEGyf8iXKUuX50ctAropxohQwGrhsxlwvFFZsvjqenY59z
iC9JloB2BF4h48PRynce1mnRFfm/N5R3g1ySAakRGp9dBRh7hKaD+Z6szb5YsMGD
x6uDxAqRJf1C5GsTHF024L/2cdr83yvSUn9BCQ/jl7/8ExBplw7SVZilaWPyjVYf
m9+de6AqPoT2iiU5ffqknUNERMwjmpmEriqyq0NxYUA0HJCpuat9o2wBeh5exank
p8pZa5xQZvYaG7pXN7KWk+Z/nvL2jOTknpunTSUNqUYK9gu4b6ujhs1z0IqsMgtY
985FiZYmJy9D+FdqEUCXssDCYzwUyzf1iZp2NXbhpFAM5mU9CcSeZKWwpqiUKxmS
6KSqv+2Hqt9z8pRRVdOaumRY9XYeu57H9njyXW0h24Y9/WcpeVxkFjTo2GW9vvdw
UBVBHReu0nniXSi9JnXvlzrVyrWCoIDg22ge5Rfzdc9/73fp2V24CkVNmwnP5jsD
5/HD+lf8D3Z78hIlPEbsWeDWtFFefVXXEDOYxrH0RLsTYzRZXlNnsNYEBd2Z6CNU
Xex6fadQJJavdffh0nEoO8i2PctbIk/HkKi4qWn1pSWTFxprpzNQxeKFMmCTl/9R
smjmp7SJQc410uDruVNQhKLWRTvuR49gLKqS3rvQBGxI/8S4xSrYuTOQ6YCRJjSq
h7xjgUHPUY6h8zuWJMtsdvV9UGuEcz/yQSSYmE+NjltEuyOTAiYNBGFc+81ZTxJj
WzsXoViKAypISfj7BT9Z3sp8tpDr1cjF98VGhZll3O2CUCeqt835BC0JThNRdJ7N
tJo5ggBLOOy51X6XlUsxHTl1H2ueiZAiEGljz2/WCSmP+Sfeu7ZTLgcUiTDAYnQC
+w61UIspBo9fTCoApgjGJuoBUW59VXP/Aii6VYSGGHWbwPl79wbBp2EzskdfXUKZ
mMBYYgpVZM8KXmBz2GNE6zXrU8ksR9Mzje159lrrRslBMrrswmjb6nMuqmyYz+e1
b1VHuUi7hITtsag3Dugb8XV0CxUbCivQGQqaCWzYBx19hItzEeskY2SmZ6ermCkM
OudLPUMqoRay6gLqqAKZupGVDyZ/BtR4GkBMKNg4Dlza3XoclQOnoi2dMzwzqq1H
v6jvr0Tt/pyzdIzGIBUaTkR6Sz2nrnht55whSMLSgo4y2Y2Q8Ip5bFHdL7fbLS1u
xOT/B2cRzhkJa1H5YxcWA7ng7jeltsZXVtos7ImN1blImWvgK9J7Aih8uRSurXZJ
iHSc6/iZ9sFIqXTsWDdrWt6U2qDvBnZv1oV0F6U9OW0+uy1XLM8BwusEcYZy39QN
8Y0qnzYrzOR28gSBLzSHMi7sz+J7TAbe7zROupI7voBMuQxyMUjTpVHiMj4pd63f
qXyyySRlrK4NNssQJ11jL/KHymFbL3S3vN27SwXMeUcImZ76AbsneugG1A6Gk5kA
wH6nA9eMSxQUw46oYEWk1RIPtHGsjHh7mnUB77fSU4sOj3s0lHZnszc63pdrLuab
LdtNNZ3vEY2X5o7cP1fNjZkBDetcgFJgImPSdgmZpBCR13nG6+yX00jvWxueql0b
1OUsTQO4WDGsvW71TpZGqBgl6Satw5cTeKmZtTVFrKfupHc1qRrpS8CgvHTyH9Yc
E014iHZfbnsUl0H8kpwoBhbTXTnVb8oqB0aerP4KZaINHF2ILnbUqTIbKSghWi5u
QztE/T4aIYwzU3ntsVsXFgzxW1cMlRohPPwEcP+O3HmEyPAr2XkoH36pFVbNOxAI
0cIbfvEIP7sJLYgZmRdCAk4/BCaGbjnX+r/4QQPk6odDNR7U1RtrOJDIQ3Z/Y3H2
UV3xtutpyg8QELt5VARFOso2beTEccVnveHy3ZLD7gg1O8AQifMSHI6Bx58dCFIP
k1rIEsQPCopMqofmI2v8W5KI1m4LrJoN4B4Nvf5IY4zWTwjZ55Ks/6lDVyoN2QNu
l4Pzw16Dse2x9SsvPsQCf8xCYOHfbbjIWBc9wHgOK1M3kop7w588RCoglWsB1uri
6ytM0u/mObhB/td/ekWodJmQIbEXLB8mlc/4xgpV198bq95wULU+olHrKIc+gs1a
PHwjDaxdpjv5R8ukHtKit7rZRASjY34aOIy1UYXawqUJSrlGIUHy0SGcT7I/S6JX
XHyfw4QgP6SydjRMF/P6nybks0BinT9gNht3j66izCokZZDhQhgYtZo4OLLFl54j
o/2E2CJHw7VhmVHninpENUdenPL3ZLPo99gEBb+8fm2k+NUuwAbbWLnRe58U48Se
twpab1O8FGpCamwoRVQiOvBy4diQik/8//C3ufIKUxA8Qn44pdXrOBK78PXJjsB8
xKOFgqTIKTpGjmC1shPc3d2AtxTXzAaE/bB8MsYFMqIgXeRyweQpIT1ydfnFrH7F
wRTtDZcExGK0cmlH3UG2I93GROqueZXKPc4p6p8a27I0jXRaiRo8FPnqpS1Z2I1n
p0lw7xj+uFLpxnjB4HW4SOf9bR3twr10QJTnkecU/1CrZUQHF74/lhyMppjMFVab
Xoxfu2bI3SJp78S8bQolTPlBKqsmSmikS96sczcQpbqQYo/aJvLgeM3elcyXBedI
/aqdOMDLVPXrUuyyJNw+zEAeABtvBmT0J32/94IqylIBiEEvDCDxev0HFQIE6lAf
BeJsL3bvdsx+dZrPn8m2VP8LHWeMk8DNYLWe83nIXUFLVpa7qoL6N96zp8NCx/at
l81Bw/sbGrt4ST1ij+FxBWbk5EG42Z+2zceS0UsWDKNkRtP7zpkQdrj5zu27U9Ud
m2tJ5fixz8T+GN3ksdpTABAjIZ5qWPLxJ7ZFlRJUqVKpUVCckvN7N3eEBKgdeAnt
e3mvvWjXDFHiuLtWonWEZXPnnl9QqtAITam02cmBsD+DA2xElMJe67IIW9m82CMu
uWmusnR7xzcrVVyC2+op4o1FMCf2l2OHsSbGTGVsM8GXrchKaDh69ZZGiqcmEwqw
WpV7rmJgqft+BsRln4MmEgvCnagySp3OhqsrjOmCGfq921mk+R0TvojITOcKruTd
dpx5+AbA+OFf/uvkwlJJZ1KXjtUnUqO4Vurk1enr0/yi2dcJo/uhQIzd+wmRCOUg
29bU/wcPVJIGWcoyCj1fuJDd1//re4O0R7b7yBb43ofG6IK61rVz4YEXD3uaVtPu
ze/Xq4gPMui70bi0J3e45ESXXQ8QfWVm594v2BreYqP7zpI6+r5xKP5YPEk86rCp
1ve8whKm6Ole5dNn1/GmiWpwfgw//401dNVKSnMToiH5y9MTHph52IzSmX5PLcPu
6DWXLB+ntmBBTGhjut9IGAzVz+OHmOuvFQ3MsaFQojR1gxTcKU6VekM64pQarHEk
OnjbKoElB8hN/BLSGATd6FHWFmEftRF3RdtV/MPLAE6nWlqyRjlxnOzSFN6vz0k8
LnhSYIfW4X0btZeCIonq5XXBE7fFSMPr35Ii3i0dGEBA3v9ebl9AyzTK/0yJJOfq
eEDHyXxymMjOWzGKLRIcnh9cDoinrcwDgdiObQllTnC1UG99skPf8bTL/1sP0mJF
m491Bxm6+lVD7tUCIFY3hCKi8yQGSq6wbVRXNxZW+2TvfSz2yUqjwKJ+SaTgk5ue
HZO5fb1NFuVn536qeVai2MrrLWzWE7ZqeLIeXsBfp2iP4iWgcPq2CsHy9Ur+JCF9
MnJAdOd4I4I6JrpFn9cEVHaNOUnqqqAgG/eh7hvQME1WJEnAINnvJRdbKk+kVCe0
3UR476X8gjiG35GDLmUeHqOcfhrFnwwyzLiHx5Q8CvwKdJHusn8/+UtYNjGf6ugS
Y0tcaRD/8Rgo+VOm1n/oXSAy6JUmniJGRkFSG+vuRTV7ON/cmJRl103FR34uoPdC
lfPQ2Rb7qYQPmxv5GHSYlsxWHu4AEpRDTcK6d183QsqsO8DkynDIAL/1wMzQrauO
pEBQ6nRfny/S1UL+h9O53Pt2GgN36Hxvl1h6+kdhhiozPv87khfOI85bmJJLYSGM
3udXZsFH7Drxkk+h8LkJREh1nB9ejwn87ItbqLiKxwIkPM1lGbJEOsktnhgxB+gU
gYr6r5jUZOa0fFLtCTBAwEUvME5pipj/PRNZq1FzXHREZR7uyG/E/IIc5cOAWPhe
rrDc6Iip4q5JPbU1dnDPCQlItYB2R41DNYZi7Xa6E28OlV+AZAxBZNpw6djtTp2M
s5kuaTiin6mOzPovinwrjia5e2Z9jEsYcyHE//fln+jvgQzLPnsQ1jmZDJMA4p4d
V2lq+BglRrjtFlgZtumIEnb/li+OBZV0+zB3cl76qbPPz78gCOhkYQWGoKijVfmF
3RLwcM9EJmv2Cu+Zfq8aTT2xf+xOej0OmnpnelZlZGUcZGSNXl3QhC0R7e0R/9Mb
TvkiB9HjKpXN8CiNl3b1nQayr0WfpE6ZXANdnywsSCen9kNy46irtKK5Au52j83e
RtGvQd7Km9TYkUJg4D9rz2Pa2e/SXmkEsJiRa3/fmLONJQ+mf3IE8WacjgiXjZxK
6MPHe3ywacLaUhzj98KLMeJoWp8Q94iMG7xV/wQqLpdsfYxSKqEu6UsS0hW2PCGV
FECbvq7PB57WubCxMwD8zmaoDWiCblJFS0fUlKzLR3HlMjxpBF32SAgHF4aIXZjG
pGtqRlnhUppqVXLOm1QRAJFzPeUniTNSKuSJIjRUBVz7CQjjlXOOAPiWV/VTEtHt
sn3cf+4LdRLjHF5qrmFo7VOznqB2swIJ+9pGV9cBApHG/KAtBDz0L1BpMKzbBQ57
pz7MaVni40ouMYiH/q6C/fLKa3O6cl6Dl0+ZyLWK3xZ1qfqBhcZCH42KB4w1SErE
uGk7KtFw7k0xAUP8g4fJwJeRRqJPQ015eoFnhsoMxgN6c5nosVsM2gEeE8McYUhD
JjG06NNtmh4p/HuI36hm3s78GLEslxi5DSIz3KdkcFyBnD5297xAB2LA2iK8lllh
8vM7G153WcZWTds13MXdtQFOHguioBdN+pDcbIDNSmlSBj6GV7wizX3jbhE+SDDg
1UUzC/UXuDdpM90TbUsccfYLNHDryS4dDBsAruTY02/op4S4p5IeTukh+0GagXxF
FWUdTUt4qZUhj1cVCB7RTirKiw/kGyCFgk+TBK13LO9XhlK2IJCcZtCrmUq/rOji
t6UxIjsfrb0ZL/3X5/pPr3Ftlv8rsmu2X79xOP++S39+qo8/6QT5ge4obY5AFNIb
dxfSUrClbm8WiAoiJqH/aSqqWK8prA299dZuZoEcpn48cP7Z9L5BEvnp0rXuHWij
o6kX7evpSMpkujIecK2RHaqW0mdNeLwzmgxkL12XN5jIgvNQ7qnc0wV9U0HhH81r
tNiTtACldGAI/VtHFQQ9xKZLrxT+tfyJRW/QjJjKACWRoA0wrD53MQ7zhnyDQQR0
IxOJfh30AwNadoCkstM7+3oUj04aK++IPxY49aUp93h3YUzzY5ZNXGdtPGlOnla0
7fZ+4xJDmhgF62sx6yKj84HxFgh7vKV+bFvaBeolnmki2LvRvq9zgx3Lyh5TIq3J
Vi+A/wXmk8HtBWREtKq51j+QfIkQSzd6CaPHHd9c+K06R7Wfzr+HE3nu8A71F4Aw
h8yYH9t9J361ifpYMzKGLqDRRXbtKIejqN3ewQi2dInRp1TlneUlAlD2XB1n/xKW
KqtWysI1zQrskmgBKoOE4M+ZzTJgtbeS5NZxseD40h6IIsQEgdQo8JoOSJcBX8lH
AEKOdJk5sBB+ueamlPzRgLFuxzgvw8n7hkO7m9b+prrOAvtGtOSXW0gk9EarXJ7A
6IoYgwJjt2j+rkvpJkFDacdPuP7yfv15vKh7ZU2BQsAl9ILVplNTwdu1JoL0GXXB
zMmYQftHtGAtMIAq4zU45qqg17U+BfuoVXlfxM4wNu3n+lFpN5AfYREbgR5Emx12
JIiLYgGnTrlxnhbvCMWfK3ZE9XxVcBiwheNFekudJik71/K8pTr+U6O451MOWZ+Q
ra74YTbH3o6J2h1X9bHqYYeUK02YMrf81PCnmfItVYocopeH+ygYEEeafEAdaBcF
l5z6Lh7+pRW4FGL2vMUOcKZCC/uBs/SfIRVmFMaAsw6Mv8k3Dy3pow8XT7KOnElv
EWrfvnzfqse0ZvqQr8pYLyY+858FIgP1zZ+4jhvtvon9La4mWKolggZI5grFZ92S
73A9ZoJ21vodC4eNzsSOSvuKP53xoQWOIwgyHXYZJnNxRvJ5GbvrJuE+LRKMN91T
t+gjYfWHCeZOQ7Q4OZ6QklU/ZKpuZbEQpJX/WkxCERgnmLjSF907WGSdSCuWcazt
Ke2D79SjjXJoJGA5bPUKSAH33IcIH1pGwoHWaakG5tjYuMl94gfkVvdz4hc9Mr2G
jokFHUidPH8qi41IFkCk3nRYr9yP72jnMrHLXbuWdDb9btdWRagTAC1sFWERyIf/
v/zb2y3P60YWFA7DuVtT30V7ouoCiZz0JceLFo0Nj9neFQueDvEkQD24dV1XzzaD
AnSC5xFaVtdpGq8meA+tygxEykr1fCSZ5exTJB8AnsYy6DXSuFm0Q/JUEkNkSwp3
hOMhyLQl7sH7zfthH3nNXdalAxmEUOaffy14S33rcowzDjLn/AaJxN/zy/CFxdx+
K6914g1qFtAknZjjEgdUSQEo9ymDiXToExvUNFw41A+grwXrNmxdmSl0b73a1+Ok
IamwA6rAUllSaENIP6Ndc41rZ9nkqYKxAkNECPMbDmaFOk1GZN0PV1pB1jisi2GX
JPyFl5y2T0NMvdjtqAU7+RE6pGMMtOwaYBS1oIiurjsUAD/MqY2G2fHagamuNGTj
tMX7fYVqRerRWnCHEjmFntgn3K2+ZvZoHb0OtLUNQFoz81jpVNaD75QwoyaC1qvp
5PJIX8FIu9kJO5tvIHWz7d8Sfylesa+TOpiSPuJG9XyxvwDka0KuNUoTE6fO4DSJ
rJiNGhpwLPMC3Xldqoc70s+cnp8ULxm1otk4Ot8ZM+jo9sk8tXrehHTUOtGJVH2i
U5txifJNzzarbL2xZEENNnineJfBMCnTUNKK7/NIi236rkdDujOAUZjSY/2f3zGP
NKYJUlcTW65CpnbzXtvb15/ruEKUMZ5KGLTHA0AIjHbhSIMGPmtwNliHJBu4QziK
o1z9Si/YjYBLRIl5KNZY+6wAghWpgJCWy305cjAQP2C6Qh6KGwjFrpyUzBFmpOZy
H0410Kto9czMwMnXkqT5l5yHIX1tuX7as9GzMEb8N4K0Z9nA5qC05rNQiuGgV0Zn
HFGKzCVPXtuauyB7lJQkjy09AREY9m5j4BmCSdz1jnUVjUSnYoyPpOlHlSzzL4D2
XaIr/1yfJq53VtehI7WoQKk5BDefU8xyy/pDbvoAISlm1jXgjoWUWikvu9/P9Fj5
cQJRIgxYAfkESn2WNGPTCIEnddk+zqAAEn7NhmMaAIw51xs6CMkjH16Rp/c1S23q
Dsyf9b+H+X76nZIwpbKYoqAGE1X3Q4rvdjqkSV10G2QP452Z234JfH0sjjPpyQRs
8Z6vpKo6EjDKK/xJJWXs8sm0HRubKvAFCaohI1elz7INvqVzHR0LoCoy+/eM/JOH
eFDITb5qDOnn1SfokJnlMQQ8g7eGAnlm/8W3+/15vnsln4h5tvgXsJpMek3KuZ3v
LkyeNCqT2TC/6EsK3kK4esGo3AmhWVV7boJnt3qKXh24krtzPM/Z6h7aPIR4jRcL
97xAb4pDghjtNvkjdxj8UP5OgGaC/r4bhQzVLmM275QW37jyVS8RImwOt6yaa+f7
vPcOK7p5s04vlOxRkDFaS/bO5fdUx0E0N3KHUldP73v//s9cSCIC1lGsezhYorjx
xMflGDqzy4flvdNMI1tnlMr4m64PXN3c/+yYJ7PVvVt20RMTzKwqrg2/YRplbk1b
PaBrVOSTGMgaeT642LN+jAxBhrZd8VTwJpMJuP9T743oQbHGQ008wBjN2pxzAcU4
iBJT5SdFxe4e3Ns9FBMGYN1iR0Noi0QvJQYSthB5090BBdmXSeP7chOJ9bToQaJ/
eNKIhdAswxLTTL7DXf7tOOaitZZo8+7EKjfAywI3z2uI1iZV7EwFkkxibI0cn3qk
kZYxDGvFl2iMCY6EOg9vlcCqXJMZJ+Tpbgwp3sL1mJisiA+jycYoUP3tuS7N+l5L
d2/tq0OENzA8GUUV6DLh7ORrDbuYRWu0ACgn93F/r+7vStl+OYOkmz2Km5FY6t5W
ZMmwLnCtH4UtXdCoueu0m8RCiqX5WB5qPoYJ+3RVvLQBkByNEpP/hhhPOng1uQeE
Ou6sVn4gEcqQCLsG5L3ME9sSHfqw1UIpcQQQ+Hn+bp+KMVqFumfyTTyR4wzhUK1R
A00Q2/Em+0kso6q5qSvOVNkJ3As7p3xU9QkMqfvvAPtBGwwRbZeSrnmuDkKhymc8
KQ2fkmVuDUx5NVJwnujQPt1Q0pwygxBMLjUAlSSCkvZ7wtLrwrJrZtksr3OQfXGy
fSqHvY9W1x7qRXKLfec3fLgm9AQBLznsOOZVBzsBHVCTcE1QG2IOizGXkU+Dzoyk
fK7PqeM6KCDoLIx2y1XH8JPi0D22uK1NsXlUvhILPBX1NaZzgY1l1TujeVvvOsSL
0iLFQgl907vbxn7YIz3ic/+fj/NB1FJ+oRMuhg54ONRUbELlmUbvIAmYjGfrEV0D
dyO+PrR5i/CRkv8CWscfMa153Eg/JAOEtuOZ6/kMQEo8fCITdXPxOZxSX/yD2LKF
zjs5nHt3Vp3+QrdW46vPDTjnYNw9PNk1b8kX7MiQnnEuYbiLb6tELKtjBOhxoceZ
hWdKr7ElnZZeqfHoOIgIolE+L7hXcLMOwi1mpuXbqu48hS0P2VnPXDvpxfL7szKS
9Lg3CmNe6dMRPEz1ikZ7gBsSvLvFOCXkoRvBPShENorMk/76Za/ufEdqF7Pdc9eU
9oSedqpz2hUXGYTGcWqgS46Oks+qNn8LZ4seRymAvHfMvBmF9237euxIWe8HFIzk
28WNnwmE+YQosAPok1pRBwgQhWTReaoOrqiwwijX+vmvdryfIWm8zOpYMywdMvK7
RTtW6GGEHVHMS8cnyZ2QGltTF457HeJporwto60aYYk9fNh1FLYOid6I0jz+yoQK
dwVWHNdpbMmuqQfLyzNNh7Xs7UBnKSRtUqJ2SVtNt82/mMqn/HFuESVvugNgCvx7
fhNGYeLETQyFG2SXxOqSISjeOLX4JieT8P2vtBmlRNjpELcTCuyGDZn9Vtt35BjX
9Hz0GyLf7HLqXkTLOc8Xn5frW+fDaK4tDsMo4sRjS6tTKBggrSRlTSz6CnGXTePz
y//LLeIFu6B3Lr6UaMpwQIFz2o2eAPxKxy3ycDKjGFptF/wY9ZG/QKE3xsS32VVU
iDVnRtuP3OmGKF0G2P80El+qGXaHRNUBc9fSC+2FY0+s4rkYCrSYh1DWTln9Kl59
aGrLE+vbhXTEkrRaZxFs8ywj46tZzSbAW+rDQTBUa6aVeBG25kUYZl1x23uSwLZe
WnXo1ecCuEPtTexUEepnW6HlsPyGCmUx12PqGV+wPlolhqYMpC28facNENQJ7I3/
rLpVzyS17pKM7WDH4EB15yLdufJl1PMCZ8RWlCYLKf9HH7pL9AChm+MzwkJQoAUx
ZjgWAQ4rNuUKyowbnQ3XPYMDQJUD09XQFgrkSsyIGBt9vQqXGv67BLqvRvYTJQ0h
FbHaOGl7264UOcJRZvOMmy7PQTh2nKlSN8wyp2IOW14oca6vJD3j5IGBz4NZR4il
kBPjG8mJv8RWF9/C+y9RQ+Q4bmZCsct65B0c99uXtGfUbwB9iT4ao+fPsBcC77EE
D+CosiyGem+Q0JswpHubqojPsphkbxZqMq8xoO1K7hjrWUmbrWLmNRHpURYMXmPX
/iOoLVx5D34vqPCI+zDdv5NjEfhAh7+87vFXT6MDN9fgdMle5Ts6VgEJAMEFT8Y5
JxO4YDmim39AY10Y7GHe7fomH67BxmSiwP/oRLdZDFubHLkNvPyGG/4EWjpa9S3F
wCqQL0FvT+vBhdlph1i1prC5S/Yj3QIUQIG7tscLjWElJtOsfNhHAedZkcIrNuub
nvRBNGbXqtJVV51jo/F2iOEcRvAoJ6pwjfuIFia10AgBXt2HSr8xWECiJZYtR7Lb
xx4nO7pP3WNTRx7iY26omt+p9F8+1PkpnZMWaAW+t67bMbJLkk3HXwqVJre3elVE
GqgtlgSPUK1B6LT443NIhUKPoPooWILZTYfmmoUijWMzpeyKwObByUzqnv/l3ucW
BL862ZXYKmMUkCkiqm66JQ7kcIVnePM3YoPchhKnNhvre08/NQCJozhUb763xzAp
8AC0J1qSLRJvwjFcT0GHU5sqMHMhboCTZGa7G4aU7u89drW07NRZDyQNFQfoTpkN
L5KwWnRm1p/sEKR0FkPo5tzBQ50IWjYWtoiPQLZxYwWXKyUrWoUr5Pr/OzYHsLY+
n40KEtZ9unrmuybXDWjfAhBwy2N2lLo1bl3Jx7fesDUUTILRD2ROHFbdJwq6YpB7
4jIEtddS1rg7kPKEbbOJyNEN6jmf9cpAeTrtuIxq/LcXGzLD09wZRFopG8jbqwoO
2/4+iabtXUOitxUuby2oYC51+I95cCmtVn3AueIjIbhpnWUo8ZvsmslmiwPrKjgH
larYn57Nayu2DUQrBk6ubVILPcOkEKgyKOYcI6thNuW/BD5oDrUNuudGaRJbG+tN
BfpGivqTfXqy3Ghl0hVNL6KcCPMD5WevpG1qvx0qXCmTiiQCpKhMb2jgM9Whldt1
hILOuuAJ4JAKVu+J1Sv6024zWcG+XOkw3QvKaPLOxOfwmG+imEn9Cy1x1hM37zO/
v6z8Ne3zn0tpHE7MtKxIacWs44595t08vxBgUTcyCVi8xQFsVF+v9YbPJKgN1Tif
OZN4fSxnc4Ej+7OStA2DDNNGy4wracxDiCAUVnuyHrryQFvnCT5AYutJsBDhQScI
EoVEj4O5zXyNg6sUn593gMfPwYcBLQCFKgT3QFQ+oKciPTB7mlLg1jvOyduzOPou
I0RwLbRapf/YPRhTT5NHITmzl9N7xPNQTbTpP5DdvohPZh/tf+8qhVxPqKwig1/F
0MAD4k0k/rEMZqVqdLykk0g1tlKQ39Yt0KdZic49sBBrHKzUx4kjLrQLBW9LRxZy
wPeUKB18CY1aRQGqC2wD+EFt3wgzU9BduqZbPqZxBPCPo4as2goJ2NvRllWMjXwB
BXB0CGHBMig4kS8FBc5nVnk8qDkoVJLv9J/SKDHVMSukGfZ1Ax7XOR8/8GxmhysQ
ueKEtAm+2eiUrdVTxHYzKP6/YLT+X5SX54BL1iJhXdBc40uGLiHCflVInQklpK0O
RFfS+wre+vw322M2QZqrDaPIi7BPMmbIdMf0EJsBdCCJSk9SHETSqOsQ85fi40uw
P6ovg9fKGaWShXevMKIoaY8/98WioeGgnua1oWRh/gdDfoIrLNm7FGGvaTJW3mVj
y1PX8yennRr3hiOMSut3WaB+7hCrOFoXq3GIl0J/9PBaXVTmXoe1PFOqW+amWF7C
R2MAW+mvgMdhPrQq54LvuY2mMzYPwfunwhGjkfUFb9yjEVWDpM2NAzEUA2TKkCRd
mzOhttDTfKVadKc1GvmV0OtiIgr2VxwlLbFH98nxq6ZrU/SyBq37K+gRgzMqxUM5
9XJpoP7QvYq7sNMExM3gSRu2IM9YjNu1D7E1+OLYN2Wi6epfKrhLiJJK++lwm1dh
V04WNtBlCOOwSYsLGZnORZbB9SxmAfuPsRnmFcOdiKwKWO6VjARTXNIZs0P55kPy
/70hHiQPRbyTj1VQF48CyVldrkPMcDMYdxOdRZoNnlEbQpTeD/OLJ6Iia/qbIFHG
bOz6kPJuS4BfeWhu3lvhlNV4nAohFNYWr8q7iwm9EtrTGR9rgKa/OSDpxl+cD95y
HtsWjWDgWmQs3RRKcl2NnUFI8KnE6td8ca0lDsxVtQzIXCEb0k+6BYwhE9DbOy9k
rD3tewbd0I0cDAioT0RwpIxLVJy8YlQna9DaHgxfZzI1OGW0azfd1n8sYFURABPE
O98wUdvdcHKlSR70NiEyAZkFb+hz0jrYP9W3fvbs6EFMGmdpm5f8xRU9CM5mlpo/
1yKJtHp89cmn+nF53xx7m3OTozm9KdpHqPlkPJpCdr0VVljH+3dNLySut0NvsdSV
/vWIJ4Jv9uB8+TgXE+ZD0wVp0kkPuvKO0gxnGmXqqumn/ew7SRLk1AusQfxE0xaH
iwQtrUG9S56idkh86jeALUEi1Q1WTEO8n77O5aoDq4Oqtudhbur8GgiuJSbHoKnb
f09+kG70rEvbCFD9/M6D62l5z/Jc3Jo/hJReMc93G6/yIGn9EkCBPYsLpHb0KdBy
uSUMpC0t2+Snmd8NSQVsCORCCAX6JCeDXuu8GZ480psBA5IBUD/LLsrzS8TcDOIw
lSjeyaBgVs95OhUTagjmU44JcpvTqVO6DmMK/cTurNPE8/68VIIZV0wcntbbp7eJ
XqJHDmQbZ7r6tqc+FTsiTYrhNxPThwhtJDUZgZVdY8lucIDi2zgIHnAV4iCZ+fz3
eQuMrd1mNvmbYB2YhJ7cElXoCKOa3FFsLYF7qQRzmitXJvQP6QveetFGT/kwAVyZ
HUz/4rTeMjbJRCCI73/CESmWmPX6LeuKeMBo8gt+yLrkzmxs3AWJ4k7ZivA+gjzl
4pUxl1IttG2CQPdV+tSjo7LQQ3oisoTJlDFlr2XN8rmOwki9BtWDKH26qAO9lbUf
vE7MXwOccVP5I22P+6OpdNa5pO65mznbbapULxkEs7OMsUwWPizL1+DUcdssZLsa
PPXOLPsXQK8LSPBcqdbpWxf8pSAz98xKBBZG7VHTXySrl+otxka2B3UkJW09iH0E
TgTQ4LsW0lhnsBdwi9WCcbpqBuMZF4pbbPJ+ZjoXxGigiBmlx/eMkzAt3+F0YMDz
CxXP2YFGp+RShAhvUHp60MJH04eN+8A84qkxqn8sIwL29kzXLfCbi/y+HxL8DDm0
Bvymlxu06faFOr7PXdYSKT+nDjXkTscci3HDFENPZxoJciQu8lSwhEk3Tyjl/xLZ
u1yIAtUX89FoEcl92XJT7zqsoesWrQlnNnFXboNkv1jALyy88XBKtwdrhaiPwLUh
E2Z5Plsxq6g8KGOz5o/EFqyQN32FOZZuIJWxOLHvpOPZ19s4p0BdjDf15OJeBXZN
yV0LyQ/eoEJJkJo694enqpT/apxWC7waUqC2qA8NZPP+yVecCN/1gnviYohCEWFR
9huzy5OKvaAzLg7q9yK6VgtDzF3TuGF6xR7LPMIrlvK4bJtn0t+SMvkfUUsfRpna
9+frFX8bz2pOqqJyh0d/9qv35bdi8DaPVUVK1vNpG1lRbfsvc+yupMMseXqqNioo
9yE0BzZiDGT7C218BTod5L68QlLQX9G8Xb28zoROtgsu0ZK8yxSi7BNnBC/NUDoP
XVZGr3mDIcw/lncmddFKZ7amYISnJRjSTOCMjIK5V2nQzq+BdwDevxRR3RUyPE5t
khr/g/YSnvpz76yRX+gT2pgoIW+bltUzPWtYRvglDixTs3iBr3tqojYgky7OZxoi
cxOqbfxZ72WuVwUya2xHr5JTpksMc8XV1LDNEclC2gyl4zdFRpcU29a94NeR+bIE
v9v8qBct8xsI4vzGTeI5A4Ie7v8GgI1IAcsI2IaTfih7mN60+33gGiXoTurDwpck
K3HPp58sXjzIdrGwXqVwZtsqjRs0YIxIUwwyTM4pD5r14Vvk6BXF4hIW+pwANXXC
bTFek4Lnr3tepn3dMy9x3v49Kzyvy99xhDKbMnrqw6RWEVf4y42hgtoJX0uJLk5M
6clzp5siEpg+sZcex7ia+uI63+xMxAN92bvINN+VNtc6r5NSw4K+rm92p3GN8BhW
J05c+SJU7N+RYA3xQ+bF9fXpQRMBLQbppDmdTRzdR1G2n2+Jp9RwxGA+70Mv+ITF
ASSDEY19tFCnx2F8XYAfuXmjLuiseHGC9Hw7iHkPFYqqiNsqR01q7I7TOhDt39cR
LYvnHqBIFawMVREoll1NGNxqTfFgwrW343YCuXr5mfklFUYQj0ixXGAnlc/PuljT
7mqhT/ujYTCFdUc4HHvKY2oCrw/DqWA3BoalMneCBthy+G4GmzDuucxtE8YBBBPr
C6avVdCmsjnosamRexrLKtibrWM4WzoYHz6cu4GcGnD1VGtL93jjd9G/tMzmQtjq
IAr/ymTZS1bfuNmXoNz1VzF/1HoIiQxZ7ILdVlzCq4cNdKOyI5+ea7oo+Lsiw2jB
YELOJdpg57dUGB3FBPLuA3BIAbcdljn4QgkXY35/tar3igXEpFCZ3GoJiD6E1Zli
EDcAzgPJfnOx34/nLcl336CYkOhb9jqirvqMavEBivC+iNaqIUVJrtWhYnYcO6so
gMuK9/SzYJjtRcpSIIM/4ySmNYwwjfEW5qidJcFWE1xukdgeravU8MYBzEtN7orQ
/6Mt8t3rJPuLOMZNPmIQqS3A2ehUj3VqTVTyWC3U6h3evDA2Hp8oldOSeGif0SFe
TvSvPnUpWq1jNAFm/hf2W2oUnwAxn9KYOpeL+UYiaw2RyQtFaRJIoSQT6hsat5Cb
jLJSQFfaofEny7dYHIs1I0lRvdN9/DI3YcP6JujKbh5D8cjhx+13d1mGMPKjTBNx
VDTxlpFqd/5R4AGN0UZ2PtzsL3Q1VwU/pviLKKX1R7HClemhdSvNAJmObUs0qUrf
9buFGsMMEhy3KLCuObdemIqlOYOWlksqY2cfKCMtiXc0ud16db6bj2RASTkhoTey
QFCZ4wi6hQ7kAUPYviOfiBVP5g1/89JquIALXvNNkdircB2a07hCsOREBwYDhco1
8rVgCd4lViX2LgDLtLSHvv07i2odyYdiA6uvXZmIihSDblDmZPJdXYdwKdCcTwZh
CSPsKn/LK+YFIbm9Gu/XkbqgRrrxqlquxvAEN6iBG8x2qTYI8kDVs8lm2MIt7aoa
ECQrisldU/LRkgjF14d7YAB6I6BR7C/HCeVKwqKL1IVLupfTI73+w7oiuh2dPReV
5pFJolquWu0lmesBv7wHWlYHOJ9h8mjYS2kyItRCFslXnLHmW92DlSOz+lTcS8bt
a4krFDOlnzKz3bfjEcEnWpaEM50tiljYf1X9NRQUdRD2fooeqyX7J+q9KBFjP6E8
ej/1Zq57saopFqkxseIJSdqiTkSmfdweOhhmY1IZyk0W2UZDBBe3xppeyvkQBKDH
sdS3KEBFVY/RVYu1f1BOH0xcAYKvJG8sgwGWw4avk0+XurFPzvY3e53eVY6lyb3p
iYCQW7Ba36AXSQ722lt9lKN94Zb55PBzlpEyulsOriMyZry+8Q8pvcI3iUBgH84p
Oh1tZRmkHG9I1U7l0J8HgVXhRYPDLr1KzyNEGeK9qYj9s0i0FrbMeB7J1Z9WPw2Y
85mTP7IeYhyvxTdOg04WL1cn3keu/vh7zCkwc/j2Arlm5jDoxFcaOWaNojVOpEis
Hj+YzjT/gyChM/q2deTgzY4FTFX7uK2McUv/Tf2RIFlTuqEEO8Jp+h1FYRsQu+WM
POh8Qrp9yVAO+joLzDl8uv+DCcEmWL8GE4f6dFK+5b2fVdUZVSwd5UdHA8A7oY2r
vvhv80Pd/bt/fLkPcvM2D1V9QtJnBfCqg4bAaNFINCm5Ygc/bC1CqzCasdyb3AJv
Fw8QfEm9nyjHnuraQw2XjhrdlMhIAuytsFqMeIFiozAO+Gp3bFAegy37WyKEZ/4s
gdE1q67nOIbCJqQtx3r0s5ppDqrwWhHlzr9/Kj/jNeamT3T/QaNIzjfEgguazau4
ErbEuMtkTDB+pFftMcu07KNfl6RDgxTM8yVTJ7g5c0XmqnXFcJm5RF1FJg1gZot4
xY/foiwqtgvax+GJNpTGK4Ak4z8QGqAMhQbonGzRki/U4swRXFYlBGvQTx/kRAyP
8LFhskwq+QLfe27cv5L9C0OLbkaj4vQVy/PqFXWcVZWYAcTAoJraG6nd2WLVxqaX
UZPTXbNZEIXUMBCn28Xm3I81ny18ylmfcE13a3NJYn1dlX8MK9nO0+bW4z3WLeR9
MyTssn0n1IwEHi11Tpmci8TIIAaeg+6azryYR/JSTYvi+D5PkT4s9yD/PwHxERAV
Evvj3aIN9SXEt0B9UY8ttgw7C9psUFQf21upOf83hUTovrrGlXkW4QyyJUdbzhuL
Hzl5v37OhvyWWnm7BQZDnyim2Bscm4gsFN++jWmDwFKOnVpKlNnfNCgqUs7/lK4Q
svLh6meT8QbHDJk08NGw3npDfXFVZpFBw54PdHsgs19d1pj6ZScPXZvVIORA6Wkw
K9lL9P+/hMSoF4SFyBUv/8t2ylLh1soK2dKHJPGSzv/rRxEp66A1LTtQr+DxSJ9c
n/s0GN7TjP+oFa1uMfCe3Ev05aK4WOhIjgbZU3AS7muK9kwqrVTHSUnXaOrnmwJ/
/tsYU/VJyPXVro6Iyp2p5FVIbKgdKwUDwbvzJ2xlW23dRxursE1sAqgf7cIoEwVT
AJo6qnOCHJw/TpcmByg78FRdXCKJgSZthgig69fgmT7Z7+Vx2QPwDSIq/VSwx3eA
mEc/qPQyKa/ev9lOosMh/2rfdolfbRB6XcswnoWMhW0O1yz/JqrfhtKwVrR9P5Xx
E6j58mkapCJrMIjc76adNXc+Yms3pNW69LssXdTnZm7vQKjbopNWPoZOEtBJkpG9
V7JJfpTXKkxllCgKcWJpstfGN9Rw78IsN4MMO7a+N/Uuy+VmGJvArpyY+/Qzls0B
EAngqwnfDNgsXtvm2uZMXFy4/EojpSnXwBRI/PxIswnNbad3yhqDh/xdS56qMuIw
GmYUPU6xn4eJIpO4oI3HmTWklvhkEkR0Tj8bUIExkoSWqN0+K8Auf4bjv+3gH3PQ
r2AKstlyN7ViwMF1kLpam1hj0uulKP/Q1sFqapnnmwNXFyoJlm+8dTTJ8A4TJkk1
oAuOJt1zFQzH/pkX42iDYd1VKVjCMaImy4OpRM5OcPCgkaYaLj6mQ8tpoYw38TVG
310R4EyEzo7H0tOcDl9X2uyt0MHTU86krrKlNkmUQIkl0VNMTVrnvwV8WMOquwlk
jLJhIfk+7CoO4HXlrWvWs3nbLA0KSe9ErxdcJg7gDeTLag8SggL8ZYbTBNIZyub+
botB6MDcEW5vytHw72a+No4BJGC+XAd4FCoSS3dX3cInkiP7S5icD6RN0qLZgoP2
mBXlWDXhlRVfdUrNKzTZnXlYoQgphb4DgGlFTWvUzFpM8U+sjqQw5p3oZKTXexjX
se1A85WlDtv1YrVNmwsRwjZLzvQuYBRcD7FCt/UrJ39mvM4af5uixO+CVuaRoiED
Y1hTIwNrGM38zpgYuE7ulZJaKtRd8fR3WKEg+ugsB27skZW1hHjTeNHXdciQgRMs
YRH5DE2LjSsoA/CkSxBRK9nZtRcxpo54FMZxFUT2EssORRjeHs28ouog6qlHPLi/
Yneu/mqMwPBIBscNKUgFj0gPnS9c6lI4Aavir+wgACGT3yjVtH4tWg2iJesmm0dw
TYUCybcvbyxYG+c6deUKtb5+uRAvZGUS1OnEs5C0WW4aUt8IYg0f6Q62uNgePyYn
L4O4jYCOcspJKEykVlWvsH4RUEh2AgK1PUEGg45hTqoOGahp4mX/lLmkxOcrpXt0
gyJss/YGrHzU9RvVfqL+74U9J/3XWBwS0PyyhNTOknocj/GqUgNAlZl/2/C2hp89
10lqmvtJHpun9GVkqxRkNz6Gm8eXIol6+Q5zCaiucAOfee9FuybDiCDyzDRGna/7
pekwU/A+sgY9NLHj4qBd8s5mf4IdOS4F45OcRogX+bl1ItrbAruKHgdjHj6Op7K0
x/3kTyTguA40YB2MYJ/Al4hNx2vrir0+OVPhsD3LovTQJ5ZgTELBVfBIla/17kGE
GFQfqBCV3tMUJuioLzD7mVTYQlNWF7KRmhOHK3n1u5S5//I8EMwFdrXSrHJyQofq
9Wg0Mmyvw04vgmA6k4AFPNu/fJGEjUHAGDV0l7Pom8+/WAbupIZehWe2NUnZsZEC
Qcnun5JvFij292dMQpZN+ZSal5/vgvw6+JFm+KIsdCvB7gySkL1B1ShnCXOindni
8vBBmvFfLz+fZ6RAhOMurvD7RxyfL81hOCAc/8zYnRKjUGqbC1PcXeBHwZVbM78I
6wL10RSjKSYrXY54GSGNU6s/zItRtQqgbymKvIFv6kNmSlHSbnIL3QTC9uGYVz1A
ShZu/tIEhShMaDwXfReHidNC+8j473JS/qeI75o8kFEfs418BtYktitKjvhHyBSD
afYCtE+mk4fIdaXm+tBbBHUlqLIUIp5MUS7tX+IbmgtCquiRIMJsPpOLyufiX9AT
yoV+Cj9rEDBKzHc60Mng5GrvnT09PwO7vCerT988FPAEB75aDWVWwTeFCoWfsQcA
2la/oKfuwIuxJlca/q0SgJBScaFGxQEgj4NOZMLwmUQ6FB+oR/dDL5rqS9qi6QJe
cbcdX6YonoDCLtT8rObVP8g0xmg2Sg2JQSinF/cyq38IsmadQeINorE2WS4jZlHk
gEwjV+HlOCheYlWX970SmrjgypiVf8S4b4yEqlv9TSKd1aEekUTK0p+yt4uOqDUd
ceIygrOJCTI4ULAkUgAS585UkLgmpkG8+t0Ij0pPjP3D7YSKECLH2opzohz/HOXe
Ep0ovTodyk7GTS792l2gpikwwF5QMf6qxC6K+grJPJXCJvgcdNQ1tY6ZG5R2BSsl
+SyHPTl7H7hlboO3DsJpyyiNYALIKfWQw3iBX4tVAEbkkQAa0Hs0cT/qPxjdKIqf
c4dYYGUueMV/ASPhtuUEgsL6LkJfXkdwb682RkvQJecA4H/9xIOrEzns/ngfshmX
5SueOnjkdcsGQvZTyEo0ukZaD+JqF2GTDXqUJeTx0FJCR7f26SGPOkISZl+iN4Cn
FeIXZlzkTqix7aKQxpmE2MOZvMUEsU4e2IR8hpsZfqeQe26bbxhpw+Hw5OkIYvRr
OpnBzyyvYlT30Yneeb7V19UG7nokarV836efQkgQCfhJz9ZrixcMglirj+0zwkwV
l0rXeT642KDOV2u2Gp9k3BiOE7gvDebiWI5tftbIrJDNz781YvK0d2jDjLz9lH7a
/1K3p0jXM5llFKYXEC2Xg3SgWp5N/80xSirvcu5Jsqz9XH/aYVrdq+ErqgAN0Vju
qHRE3EIBxG01CUc6rq/UIOWyUtzPHuOE1QSmUhkn5oZn8YxL8HQwS83d16Mulodh
VA1IrWhuKxTw0I1B9c/tkMC2CO33iyHOQRqwu3XhVwA3S6aHa7CbZF9AFwrFBMXj
v2WtCFuihDBnZgwaaQj+uLxZ5oKVyemNIvy5TOEDE2AYmekXpzp0Z5EmHJJBSFuJ
E1W1VHYkd8rmITC6zGLJMu4zRUu1ancO8B0Y2HouYjYaPvz1KQ7rYGB+P0+g433v
aTzOnv2lD11nbmoEToosr5e57oFR+xDhRF5+wj0Xj8dAS0cv64+bthjvtcVBoc8b
x0jAZJVL0K6xY8Z4Vu7OVh6oHhNP6rVVL31o7CvXvClaFJFgJELrySUJL3+5werF
UKN/Fco7o7A7k0QOPUpWI/K/iY9qGHl66ggRvzK4lyOUj6HR85PbpORekZN/tbzb
9dLBRy+th6Felmv8axir7ata7Qep3yulVprtYvQT0i7OON5q8mxHsims7zhNSQ4H
qgpnz5HTNaVGZXmYdg4V7K2cMXFLf1kDLkj3KyBzkCZEiquDAuPVHpVqTHQSn/PT
nv4/i7PPidhft0dQSMV8OttuPquC2LT77Maf1VRRjs287pN8sZicoSx4riJGnXLE
WGkoy7WtKdju3AQrRgD66qct/c/ZTG/kfEzfm2s1J5ClTspiYMg6l3La9BHGEYqb
inUo3ZrI79JECk3/y4DOQeTMCZc1Ce/GK7RQh5bRxMxf7psfVlvATaORe/2W2Ec3
K18FtY36nbUaQY8x+Q15SFzvLjfFxoJV1rg9ZCZGbTOnDb9V+K87WFoo5GSSNkG1
cwxZv2IGjSZ8wlEv+ty4BjMcq9fZ+rwiCmQOEF+H4ewTVJYIThYpJr9Rk4/09yuU
RdCJphq+29TlI7GlYt4u/j9zkHhcEy3wOHn5yOuMT1L4d5TKeVIAJuMWEw0BivRh
c/A1pfJMeNbwhHQq9CXScgqpMRXlCx7VbxobCaSbZETiqqKXJAZJvh9t4gYsqmBq
LFKjn0ABRwSPuPUncnUmPKmVz/E4+kNBmYTA6u86mT5Y8nMSOGAiZzPMpZA7n9pC
Icm+LcNXmNmHf0rcgKUPlQfMenRD/XjSbBxOQKXa3AOrVeOJ7kCVkHfg/YfG8kDm
x/ubyLL9GvtIdoALDcZefKLH2GdrfYwSWHpBsKgLzM7cuPQXCE32XdJa7gnY+lSb
Ilq1L9vHRghV+hFYrUX/rWj1wyXTNIKS+aRPoGPRqjmcXIc+WfH2hkQrbrw6WSZR
tbq7kh68tduAwWCADMrW2e2Hc9Ynxs5jAjFK/ZxhZOOE0+Zl9CeEKx01h2RuA2cX
l8j2roa/ml2dXyNTAXP3qefxKExdSsQM5W/y22vwrnnm4f2hMbIKA7Hls3na+M+d
8mpqFpGPBYMxpRcp/nsABusI+HCMC5GWpGSo88vaBuopBhSgVditwuVn4qRJ32Ps
WzqLzkCKU1DCjhIdnnFfRiIyNVmMuhDKfmA64IVxfdCfLHCoWwlTrx7CKfyHiduS
at3OuIyGD/n9gMsBKthstey8kYKgqsngk24fKUnQbP2cZRgU852OpTiKrO8K0nIo
p1EF6DXlXDrxA3IQEN36W5QvbIrQK5CDTUab4Odqyoe1J3JBczvsoqGxADqOpnZu
YGpZl+OsaZcFT/T1TmRLq7X/KPZZl2m/zTrmInR6WlJfnQeSNSWENWqAKTKfxe9q
+8vetecJNAlAKu0LnP5LfTA99sno3usMVz7FF5nT3ROIHEGj8JMgmUBDLRSGwTLv
KIGA5lYXROUZqQNLQaWc+rCKsTessYXb4ZmGMUGxj6Elh0SKwNt6TMz3n6PsWbNP
jttbggun3PTi61zPBMkbXRbD1zsNwmhdSaDnURIp6b0lBP1yMl92FEqL49wZ96Wq
n9tla0TvVcXPnndETJpiDT2IuuDEbtuz1tfnShPaS23KPtdtp/pQK6N0UYY++5lZ
DAVlIni5vYHa7Ktv0UhV72f3X44Hb+9U6HozZcNFO7UCvdsITCQJzyR1Q1OhoUaq
xRauEZa/ghw6frdAFTXXedLI7wFsed0dwFW4bYfH0Bnfu4NfWxG2Gn9UpNWvxSF6
jX2MpU7VRSfFP6v7sU3jpBSOP5YKmkKkpKyh99FBbAEfiw/MQu0e/+oYNCItPTgt
lzqUmq9KTHwXYBjHtDv1JNNeuRBVA+rV95AnDuYjkQboLZncVgHdJRtIGKL5WwbT
GBxK9lmTbOZ06KTIZJMDgVaQQr6pCeDKgORuYWzcBN/hHltAoL6Syg8Syit60w/O
KHGOtZx6PXzBowctzZqjfZ5PBugCBmbXHr8IaCyVr11UMo1paFwg21zfbLiSitK7
M9AHxyte5/4xIdGRWLqyBW4yTfqMfn7qsFrUtuV2IjfhK2Bs7y7kzQkgX0euA852
G5ppn6x1LH237rwSHdveGqLmoQAGdmMYGkx5Z284xnTy9Zooxvv9vrM94UV7mVAE
hGpQCDa+mUWakVdxIE3ah1YVWlN8hC4MFcu6N0pyPvFtl1vD79RXc3qgwubBEZI6
UaitxkrouUyE63FG07FH/hx6vUaKq4d9aNmY5SLWl0OVBrkKb+nSIFB0ACce057P
ppZ8QUOqgS3Pt3kfbTsLnNhz3/gos9aQaHCL2BEULGaGtoUtuWpBn3DEurE9m74u
BF62lgjutibPE3xR+rPBo0UCPVFfSA7jLJjE3RA3zZcbng9f/YqEo7RnDxkyeHqm
1NZODgfo3rw1IegfAHSlJpAED3PfoFIxB5WfhzlDXlqbjC8BJeiIpAOkTjwRsi2j
Z9aHy0Ukvs8artZ+Q/B81Fo1CMevUpo+EGrGhOn1fYYKeUMdcbXHE7Y8Kn0qUPFL
s0j6i72Pqazj4wEW0EZv3eb8uIvEKChkTCHp81VHs/4+3FmrwcfVsdOwSY1WIFs8
oDdrLq0L4uVWoz4YBY/ayK3HPOmBjjVqmzbEEaeP5OTdw86h5/IW3F6ukKovLdGL
o3zKv47FTe0Ld5F+t55rJ65syHC7HICLY3MhoJMIGAbcx+je/n118IBdMQOPRTwW
+p7JpPfyvpFkMZroNzvBUWccVUOE1224Nw05q5xNgwxV/m1VC+I57WGp6KBRXYkM
HpXOJML8U+BQsIxkuEDUrd9e9gSiGI296AAtAr5AUzxkVea+bLkQnQLh//hCw+Ts
edKzcCGFCOUA7RXGHy+5G5iZJGCSLnWNxpumJxHZAaAokTq/uFVGR7ZNd2HBshqb
2W/Xowcpi4KmrsN/Aedlkbrvv8XeynrTMvl5dDnzZq0DYJliPEVchE1EsX+3v2M5
5/gaYeVF+USrooOgRPx3u4uQ2PFF7RKRledAXMrFYsPQGcPkdAfQhR1jPhTwEiof
NRwIiMcJEXvmEvTtFpnfDcPRdgHA3RRpnHu7VEEEzHdL1Ja0pf/9RBB3wJP92+YE
Y2xL6ZKfDTDfUtfsh5AG4+huqbcvz565xqPuMv4uIHdpCAA9EkbMApWwA5gUTlIq
EKx8oz534MxX2AsL1ileYfeHidH2ccwwjDREyXgIf5/GOR7uY/554gIcus9Ufyf2
Tc+375Odd3pq+I4aNRm6/5am1z9besnhJOd4LHPvsF8CF5VIuzzIg7RmcIfpr8t2
UePW5o3gyAupEU1+BahgRB8Y4EtkgoTBxwEKa6WhkI75Vq4Gerkd9Lf7Dq0zPgE1
vXAX6YpGPai6AFQ0qxeEk86+MpWA/YWY26H+Db6ZzzqwWtKEWlS+AMtQQo+osfQO
timXXHbv+smZ1rXB3/xzPdxyMCwHqSFxNyMKotdvkCnAx9SpD9vXQ++1hOexRSxS
nL+A6UzSuGNekINo+O48NNfzTA05q+r1UpaqhFAHve9Bh1NXKR3NKQl72efqt0wH
RjkKe4961SFg1qjlAi2sUcYtDlYr1DyLo+LYSRxUaeHN7zcxXUn68xMTiCk+1MjM
IMgqe7i1PqNdQ8dZdSWUqcddWziF4pu+0Z6dsNvJQQ2NfIZoRjqrIaw58GeyLEnW
IC3MEncxt0CjkwpvcFw9cBBku1jdYY3hqF45dpDP64FT6DGTSq5t6AZ0Pfg8712e
5RQD1gbi+fo5uRwTGdqO0mO5TNIPJVk/NzlfPY7WMnqZmuZLlenAkqpwU3YZvGTg
TcA9RR2OdG1AscCnbCIgk2QK3ySBrBov+ktjMfhr+l9u693j16fEYvG+LXVZM4st
hb3oTvdugaiSsKKAF5wgcNJ18ymQCVrLMDCotIRsK2exWNfHqF9f5qULbK3/937C
Xld8DCQdWAyL49RNpD6nKllDdsQZ8Q7/bfptcu1HQ+a9E/Pj/5XCA8p/mswrvYxc
wLlCbrBZfr9yC1YSYZQT6rfVZxD81763e6RyFm/PTn5fdf5fxH+l5EXOLTxTEsAF
O/pYI+nt03+p9uyTnXpalZN0E1EGagHZgwFds7VZFKhHMPJUKVc7jEQzHigT93Uc
DYguKAiheocHnw1i1171M3axkCCEeDjiCU7/UJytkkdZU7YYHvghwHLtlIZbXISs
N9Vc3tpJ0Nt2qbqCEc2c08R+Wd4Ga6Q89Z0X/ZAKrPIvYQ4b++aqEfQuqTj2TaoG
sUeQpdzJR5sGTJlya8ZrfpeVXuRw4mIIfCV6SopNhFgi/Tn2ADXGYFOxZjVcfJpQ
eDOW8PAo6U/1uu7d6LJoJSM/VqWSrCUarFqi4scsFquKMN95tepXa65bhWLeCMMi
snQWGfPUgz6zeQz/V6kG3SpMFksdsgS7w5KWiArYgtRZ+/nw7meJbz88JPcTARVA
WLdT9+81vhmBDpKQJ7MvCQ5cVYcXAknSwZT/QOPyVkqopi6dYxIK7SLb2HS1McQD
NEhY8U3EoyxnrWetSUBSw+6gDX0q5mf+aL3UY4qYYb0g+U4NC/KP4zt0HAapDMPg
lIfFl42pYe64foGpdkF5f2ZYUiw//yeBf91mT0GG2vUlVUjdUsJo7gIOB+pRhgsd
TBnewZnAjnXiHT2/dsDtimUL8DuRaFE6Ecz7SjVGCB9v+jKql0EcE/gPneFZGRCc
RkKCtynL+JY/eZ1hHM/u9mRjYOoECg3AiAm/ifWbN2CvEG69LH3gYPIg1/mw6QWO
IlywkklNu0KFIOEuSYxVHOha2iQ0iEn6BFR09sHPLNTjD2ywc0HfnSsJLd756JS6
IDDxqE2gctkBqYt4qVVXsiB48Xidju6ZO1+FCF0OEYWNN/x7fzWEinhO/4spkWCM
Uoy9xVO2d/xFqiGhr7OQ3qsmsfAocD9rY88s7PXIpW23liUTmu/5v+gJIqlHa6t4
Z+WAqmTKXwodC+wtnw8hWXyp64bQvIJR1GkbYiThDu30t8N2YB0b07OqBOy+vLgT
Xy7MwDmOAOSRKde8h6ceP3q14//mgN+/13JQR/4lGbHyYyuJ8auhaChkEbf3ltHn
UON5w1l7nH7xhNdKbd7qKvddh6rLxycJCUqmDOJXUuGfoSmTx/d3BkuVkUlfL26X
/OCC4PeAOmlatwVzbPeGfGT9DvK1gAzk8Llvn4BxEpx5BpI9QSX0+ykyAIvCwsd7
KCkMvCebd//0ghs/YHSZVP3fEU4HCeHHQwi302sb8O0XPVZ1dpZ8MoYln2SSxxt1
qG3qhS1gCi1S5HQ8T4OItTSQzzVuPlqaeuh8xhQWzL68YnrL8Zv+vKrHwja7Q98A
IJ+K7SCAI4nveaLKVjQRNGWS2/I9OMMe4Sp7u6xsPwscD1jHVRdEhnuy6jJFADbt
HY/OmFQYDrhPcLiAuqJdjcrds6WylGCuX1EYA6BeILhmzagieOeUuf3zP+R0d0iF
WF6P3sTlmjmCuWkT4cs+HQhn095+ZKUG0gwcOX2C/4/Ocq/1WKz3A6uJKteJasLC
YjrFzP9gyH6yF9q3ORW22w338vuhcFdjMqGLldJBfORrEKw10HyTsS1CKgpv0qz8
m2cxcY0OGhDdSXTizvygMia/ioP/KGba8P20uMovwS1Psp8c9Bj5NZ4mdLdK5Onq
NtXajbaqIxYt6rzD+XZKFM8oNI9YP8fWeI5gv1eYibyi/M3WNhV22EzOCJ5BSj3c
Z1gBZkJ0JR3LFaDbLOCIfCxR17XgnFZL3ZzAymjFOCjru8DMPWo+R4y2eKeZRigv
PfMddcQjBdQgiQISxUK4ZFalYj3z37sX1UQq/yzvU5fXNnGFudXYjtitG1qGoN9M
nIWMyx66/N4gr3Kxidns7f7qQMzMhkRfak2Ss2MlKYG30uq4BC+d0HnkWXrc7Hco
qmqrFYzJSUOhbUVLwv7+42ZUAB1+P1JTsfGbEdxy/yZC09ZPg0/jb3z0xUxS7B9u
SSBZboZqhoZUk4WPPPXLqWlg6cjk5aKuIx02yNH69bPf/zQdAD0rg8TdCyjWpLuX
8spiplrmeS+FP6bDGuh0OhXpHZJJQ0jWJNBGDpPqcwsjRQkPthDCEM+AWWE5mRK3
riAUdY06yfcxemqzI65ETm9qumUCwysVMcfNKP0YwS9CtQPBcNF+LxoeUr5xIsRV
7PUHgGf3Op3jMORLBFRnBAYKwO6VxLD6pyA29kg1F1TGYGhpKqkDpZF/hU3DtxAS
VymIeN63Thv6wZzXC3Jea19XFsWInVSoenYPSAODAdONPex+AKkXUf1MV1N3CQXW
xJVfq68VfD/9j7h99ocJRaswu6WL2LfM+FDBObjlxp8dAZFNUGP3aL6ZV0pXHBsI
orqCtr3TDXDSqoAZyMCRm19gq53HKbooXHxhspcZV9P+3qvBc74bIU080MJkcaeU
VWSFmOOXBWbQyX/VCWa94zY54torjVE6za5mkCsHHEMzEVJRFhB0xdoUTF1Sp8uC
ZkasxTKvT1CG9RgMoFNyIQe+x7w7a3VKpFYOHoeyPi0+wZfJb8Hhe4ffszb9f1AO
zMrF0KbJIr1n6KVB/8h//ztYrtkx3w2/Cd0aRayEHZNBRTC539U4dhnFG5TwVlxW
zNPCjuexzj0YbLqAyaisrG+vvFEkQh5eI8AtfCvteOyl8XDIoQ2A6wdhSh6e1Xak
5xN4+E49wIIC/DqiA/qoTdhevLQ3qVn3Fg6MI0TxvQ11D9lGTau3ezX4Hu/JGBow
BJ6GxE+AYk1MP0B4OiFZgqe5BmrQl2L+GF69IDonQBPEwjOf/lEduf00BRXwByg+
tyADDZVK597dg2olY8W+NhMWd4OavYwc6YWEIoRagSlyHSl0C2BCLX95lULJkalp
jE0ZRevPnQlE/Ro1CCmrkUtVC0gYDfCDybK0gC/vOuuxO/pN1SiLyjA3VOuU97Cj
uRSscvy2WaikWlFalW7NmPDHiavlC59559iHGelNcHnTE1xt0MLTKra/w+o0DO9v
qwL5wdcVbbRN55J4m1CfL0vc3yzonAE5PIuf+BLAhGEzpOAPVJ/XMy3mkN1H4Z6M
ow0VqtdsZ59sHFl7px2+yqfIaCDUNiFT0Z9bs58ce76LGvf8iF78+Utg+YSOlX/q
vA4dRhyOj313ETBUYhb9jlkzAgsTDMrUwoCzLXWxNVra9uQ9n+JG4HKigyskH6/t
VeSHBK5iHtHv5qXzem7Oj0JHYDsEU1pwYoFExZ/ocW67SQXso21v+6AL2NLP384W
elLqX9FaMX30gevuVFLID3HSRhAZ6ZDi8ZQoIHvmUxNoVz2OWJ26qhJ2Q74+pSiM
Bfh3gIhQqp70Rt3dasjEZc4TLv8PZYF2Ch9qniOBsoc1K9YkVEYmuRvkzjnENA07
XQkEimAJ/phMg+A/IDTN7lHJFHvZPGe2tudTzObQhff/hEWCpwYhUHtMQnS9/xA3
JbtaMgEC+a5QomKDQ53wjmeiVD1ntXsEbSi66DiYcdUuB6VyELrAJzTrNiElseiW
F0+uSLQc/+CI7/0WoO53idhi0gdM+ofjdOX0JSIPGEWLTaHTnx5ddVTx2BAe1o0u
yN5mfcSPmNHvLMRweel8BYA2rLGJasfqFDYflcFo52boGLFc3T0FpgJZRAo8Jm4s
2uuIfrR57IhbOcyrv2EjaQ8BnnAhAnxxyyLT3m/aC05OtOJNVr48S1jESDpWpOtk
tKPcB//TYRbIz6laCBjPtkthe7cYcs5Xy+H+vT/8xwTLstdt0iODzlJmZhi+1Rc6
JZQdhEOdFZr2MS4DmPhSxIDtR81cYi6oUJjoO4PC+ajnM58Jxz6RwryqIdkkxgnJ
5frAJbAjxu5HLXkPOPwNU41YvjWDMONxsDSUYE3Rg11bTGJC+0DPgyezIHElgTEa
umgMmVkaDTFTiC61cwUrV6VOvsf09lflZz5/+xy2/BoI44XOxWr43h2bxOqL6xvG
844Odp7OXjFU21xWaHNDkRX4/VU5uLygBB7H2znMcovMoxQ6r9vmIPwKl0AH8s72
TF04RviV/jzM7Hi8k58VrnQlIZ/b8RtjegGMWbXYGMRm5R3CPHR0fjLXMG2oOomL
hNkN1hmuCIH3srHozBYHAHyv31G24i5l4Pra1opoWfyHrZFWRDt9ennlVsfEUnJJ
iTmvYcKb4tbeoA6Ja9oxaV9v+YFrbn9mnd3WILfJH0O0RQ00KkKdUo9I7zBWjJmr
Vu5zPHrfqnIfBvnxges8p5rBd5/jTYl9nGPoh2a46zkLqsL4DqGB4rPBdJ3v7fJk
wTUjzCWor3Izgypq4bMNrwPqtGsihruIZlbQkMlJnTy9KCfR907qc4A/gHeRptd4
GXZLMe1x4HC/ndIHG1QrS0JQh89xvf/EcjjmmyuwQTCwBGga1wgZRX8O0EE5EHAO
SbR4TF1s/y/3iQisMxDa8hlHf/AAo43SgGxGCEjgnDu7Z2oloeCr/WIDN/Zf8Din
qVlptP6qwXpMBfaE63U8D+r/kV1prgXjGtYnrmOGXp5JDMlJsbXGIk56f+a2L14v
ORYExsWz8mwR55ZS8opNQnTLgx3sNVg//GlQJB87QZo5+/5mYuTF9mPbrAGP3Uxd
rB4epNjwN5hVUG7V4WtTmB9goolE7nrnbz3oRwsX8Ep5xBnGRLQ9e5eZ77VXa86M
P8HLzZFJV/wOQs38IU97HpofRPnkCK589FObR8Uy0TQBCWGu0GzwDCUZt+Bjv76N
FaRSRu27rIKQpEknc9UA9PxmrfwmSmeS3ZGLgmKiw4H4j7h1c8laQ6fytcICrjhc
JYXaNnZkJkvxh4+1maTMx2hAgDColHlSknDJujoPFs9rA2DPDT4r2h5gBoUdxe+e
dkBXcHKfuhUglbE0yq/9nyreBBsbAmzOaO8cA3V+6K0BM+Ws4gI4Cvcv9uBuWy6I
F+XM3Ua7Jwq4pW9bW9QlCwxuXHsCiO+Rk3Owo6RNMJUkedTjx6KjiNLU9V9rZt1A
omOYms3OAi41RF2KCUFU4oqUtltWmqXrp05mMrahsfxrTYDKgoEZiNbKhIei37Bp
UklYTnYodSs5BYlH9K1S1X5cKxVppmVYQpFae5WUFQMfeLlxCnPRfz0+gz1DVf45
yhxXuOKp7bj+gVafsuZkd40mAPKywmLJiY3uckGi7ShlwVmvn3OcYxhnTimtGrRA
gOImuzCw0RI7QfqqzNsybHz8nWEzt12+QQ23w9knbOW/A1eCzErhiftXixxh6gMR
/x3Ak9NYdzNG8/tLUddjueLgq7RB7pabyqsH+9dHJ6EPq+N3a6GVay+rOFsUhRqh
Ux/gB9xIZLFFbOBd5MExCGChHIF+1y8GlVIYjhs0jE1fQeVeavjdEUSNLi/BBoJM
XkjKHppFF8pVUGDtygt1jRLw5RVOkJHLiiUkFxeMUWxOErO9irIZJBtoCk8+hVRt
3kYPwu4xdHi3R4yYIm6jhO3yUL3Ll1+6xGlvnEfsMVKYdbPHyTBAnLtdIKj8js0J
RVFY1Wp/Q9GBYSXr39g64IUi7pkVg/Jr5KJveMiTP2Ng2zZiW0G+8mnLG/Jyp7Um
mddbuSm2ypUF5yWQfVlw2BqDJ76636Go6hMh2TGk/E7zUOlW3YWDwdvS8onM8y6g
kKrIqUDL1wJStHyLilaoukr0l7uyq8pF5+toMTNJtIivHIyMdK7Fe9aFT5aaaOQO
+asu/vGgqMw/8wv0KW5Fa1zs13QpjrG908CA1/m60wUvlM3iq6NKlnHGLg1vkhKZ
pPgNwv+LjEk9NjOOBFJzIHTNqNAnNrg+25lj5kpVUVWk6iF+42OtDIW+N3jtNvqT
/LUtPyZbnDI4BiwsGs0AcNE/2ShtjT7vsJew9GzZrjCUc+dMN45KEP9nPqK1s3mA
FWQwJr7Zm53T6vGt2JSYd/Xjo/OkPfyPF4FfxfJgkiNd1h6tnpfbqp4OPGqaAq4m
I0kiKlqFzbP28yTAN0iX1HCMB70dxAkES1Rhke52TamzXDJJJ7yUlFxyyJ+9K6ec
/L0A7UH6+u/HT0GUJ69o/NWANrtYWDtn1VAOQQr/iLiHD+cellbhTwQcLqphBTFX
yRiriYdDIGcFTp4H6HmRoiIgMoOykq5QvspL642/kVjFXBeu6dIGN/9tXKCYSsys
iJoIwXjeCdkcvrPZfg7NfAlYl0bK+TUEEGpzuOUNm5I69Nki6avIN8xkzCSyy22J
MMdwb4jUQ0Vhpb36TXdvGb/GlhGfKIHsXHjN0laneb0Ft6kumjsR5T9KCtCP8nv8
8bZqeJ2HXcWDsGmrqK7E21owBxj+G+CpChW7gcPCZUWdFYKE8N956xpHemFX3bSk
o4oRMIia/6VUIhAX/wMCkOXr1sfZiDWGqX0c1GLgNvhTQsL73A1gOPQTtXDHwUjn
Z9NTJbBlLA7sqMG3VBGRPFa7gTQC24S+ttzoG6lXYSSu1xubrnvnjGKPL/kPHGsY
5k43uFv3VRcUmTidlen4W3sLPbR4Iu/0yWwRfOh7lI5l/90Z2yCSdeQDP4FFhwHf
M08Bx/UI9uSjIfLfSlVKZQ9/8QU9ekKwzmIO4JirJxbtwQu25Z04DBEvRwgLUNu5
yi1yAQs1S2+qQvh+62Xe+7jl9Xdk/EATboaRo+VnfrhjnsJn3kQIfKmiArkMbjxO
zEyT3TAg4eIdpiLLoZTl2+bP2Jdo/VvprWTfygo9QqQGk9dieDxGszZMeSwlm6Ow
JHxleqf8u6aUXdN/wX0a1ET3uY4rampBP40J7sUXXt4VERWuN5o9+4J9Qz1mJc7J
qqsPI7xivHOsxsF4lQhWjsPdTK+qv0HzrE9ICFNqkuFfGWgToLvFD0x4Psn9Q9QR
yNF3eShpAFGZRpUSgn0zfW8h8fEWf5dHyWBzsB5ptQqtvioqn9rI136+FmD9176h
x9xqppcXF73uED6bM9AmL/8zTWS6f0fbiqI3f8Ht5w991G6jT0WbCYFU25aXLsra
u5Eg4OjJNKjT4eFm9rEnq0bay08NUTPw0HA+4Thx575KY06Wkclbk+VWZ0J+cZe5
U8b8cKi3gwnnsD0eW/BTQqpydrQeptQ0ykhUZP3wNH3ABIJjJHdfPbDMX2wmjIR1
iNOFyVeP33zhODVtZaE2jvwfocymtRJk18H1UGjaHoSW/amBedHYpy3p4go/P3km
NsGUvtc5HhaGvF0xIdamK1SM/YfwrXUvnXz6245IqAy7IFuS4serTjsqDSqM/lk2
EAzZxKkDgPB90/YZ37cQp/MRLsrDCfe90Z2HJqLn9fGQYQWdvWo9jykxSHSofupM
5Tgy+uZig+F8El/eJWU+S3dHVbKvKXY0ALaanqBhaFsMGsWRwRtOR6uNP60+59yg
5S2xMDhC5YHoRIErpNO9HuXel6s/gP37WpkLxfvQCbCH1L+s1BBoARm2a+qyhQMW
EsRSWmFHJcH8CHpexowjg/P1CgDt1yr3vQthNOewWqVguJndx3plYBmpqbG54/rd
lgyi3EHeQiAPn40sDrg2B6WNH/zDXiKPhI9D9HcUXM4GBCWS76QHsRQM0oR6lTFf
qHGoHlTBtO2DPcHzbFd65+qQEK2gQF3RnOZ917ZMzLnAsRHFNekOCj2dS9KfeToR
512Izm864atOLFgcZZEyMxzy7y61q4gRCzJzj5UO/adpS5pXBPhMYenXUucC4WnR
YzbqugzTpSJODHN7bhoQLbycRh72LFnibxrgT5UJsJz1Vk774D0OeWRwLbkL4jnV
lEpCEfJxQombZMd3TCNaswehl3kxoX5W3mvUzCNC/0HZdcXrRWNaxLtJH04n6sN/
ANZPgNQ+cdJZzsD6AjjEdHJ6XCEag9C/oW8D37cdrisJmXIjrIyZjqF+7uZsHQbs
TFFQxO5QxLSAFAzj+5MF+Iy+1MCBd96zGQOsvkZ2/PrlCBqDDliBGMzJnJluuXP9
W9f01mMaeC4OFrpz2PFVx8YycAUxneFygs4fTK0ZrHIVZ1k27OZqoG5Gcg+qAhkX
HW5TTxUImD20Kr5oAnNgv1eFlVB0bMDleZ3hiwJuxSpLEd+LL4LRN6jS06w9/cFH
C5XK3ygDm7YPNv20sh4hhP4ayty4Tici5ngeuxlPbie/Vssl1H0RndLPduPXAcsa
OJdfOIr6ihGAdYsdVYwUtotsomoWezcvM4IXvfme6mXbN2jsZgtgu/HC8QauazYQ
ulkGjceiCBV2FAj8kb3PXmagH3+gQrqDDeCunt1/pUSVzSOL3QBTzWuOvL9Mxz+u
XK6qvWpqtK0JsxGhMNzXfOxp/DGM9b41xt3drfaLlq0CUqK4bK0X+J6DuRaISWTz
e4d43i5QNCOMu5csA0GnP+9IMahVWHlbWb9FtZrhfFqb1sWeA5JVIbk91DycfgsB
iZL9WCKRANdRhWTsVXUX44S4ka/azI3W1jDHydTpKKtkGkc/VkTMU8qd8JP7fiKw
YU66pagtd4a3dDBI1N9v2VZO7bbqo9VoJYiNmw6oEKaKm10DYsQLuUvSNkLb0FIZ
TmPx3rQ9dkKNN0LgQoIs78w2dRFn52ZxJl0mnWErTiE++i0qGzXihgCRWGpygXir
vIS5MgNrCCnyUmCYCfhj0NGlipUEXNY/IFL5Qs33bIFDuxjfrkgXmlrbpMHOoSf5
WYfm/3fGNBtuDb6mDHnCG/tj1EhFtpz3jL9d/O/I5gLK5PPM2iV2og4uhM07awTX
zyrpDsQ/6AGbP9Qqro73mpkAnepsHfS1MnsyoGuQ7XyNflunWqhgsteIHrXWTbhy
1mw3CNEYc8xmJQGCyulthOhnOpabVdYKFqSWoyqs/nWPm5WOHuGzM5COCV65O4nf
IUHyDd6dZuFeZs2IyPMGSCWeRHh0t0Bg6gvaYAmNXHco/2l1bVkIKrSF99LqT2Q3
a/WKrGU1DYc0jj/rCyRg4CRVaYF6grofpUIIRyfiXMd1PgNiVl/FxQeMpKhaY0/c
EttMwI6eO3BLr6fnXLPEULAvo5bLMlY7Tf9Fz2Gf1yikZOZSlBYkT+EfvB0vTSzF
BdWfqdq7ZsaVcDwmQOcwlvzXDKjujswsy4ayvRblytGcrxQKKWuhQkZ1/bnY/Alv
HWjqvfYsLfJj8ajPx+PAcgZvhdDuR08+o3Ql8S7sdz2BooTMsAa8v9iFHBoLIZu/
kjQkDFvUK7EzZV247NKwv+WlXKpU0bryD1U9szBnR9nwDjmE03OLUPczG/iffy9R
oG6GyT0ubcaHvveYiy6QqtnI8BHQB4uhzGiKkbyJKWKYZYeBgrwKeVUUwAqQR3en
Fdj56ENFAxAeejHWMOhoeEzbeEkRI46YJGJzkpnO0ET0FhUrEzNnGqRgwcmwEoxD
XwtcoS1qAIJcjZPuowxdBshKsnOO4A0BwfRe5Gi1glBarncyZheR1rn4x93iH2h8
9TUN3yeCa2T+PjPPh7YRjcjaFMDI/S83ApIOJk1qzXRjeqikNS9dAA9kXPr6CmTW
DfcfqDJyRUk50pQIt7BxVaU3a7qYyDrMCuw+YakKWw4+XQ/KyLrovlLqe1RsOSpw
2B0qTV35Cy7CyFKx1KuSPR+lR3JY+fbuUuxx5+63b+sYiblm8SK4w5vI9jq8T06u
KHwwcln9QgHKo9kqH859UPOqpWGDX6/GNVWqKt/0VIcyIwAGsc1qOqDWu5pKNwcM
lIMELMPWWUB/X6IfFqqUdnQPlKkaU5j6dJjjSHqNMpn/VfXzqvvu6Rcyr+xap1Ni
zKxGyzLslZlrhkGTywWV+ekTPlAmp7SHveppe4h/JMhXYAFeDfWBTFGjoRZOuZCT
pfxTfg4LJvjDJi57AHnki6hpEAnSh77mEcbl+5bH4W1nuCI33O4vcabRKe1jSBkY
+ccTztFMOTMV7T2cc7FqCCc2n3OcZAEBrKiVTCtx/Gt/O0Fh87iIJBvDwh/uozek
d2DL8ZZh1y5zCsFMIyko2y384gg1m4NoIrttCYduP++jri7PNHG0LK8MEmRDAdr2
GGM331WIMvKJ4crfG4rijD2TVWdBUzgwlqufeIFPgAcNHkRCXS7FvsAq8Tz5kTtj
UkfBlBkjo/lIn5uOt2h3k9gdg5/pNxJznXYXGAT6JaXrwowM/Zm3HgFKmAQpB+79
ePojAbJwNQ3dPWmlkfpXBYcdDjzQRjm+RjCRsol+cRcGuOmdSOga1eNhvOVHAwy6
1o1za8SFjxmpLSxl0IPX0hv6c6n3KiAekZCwlHL5rGuaXp4uPln7IS/Tb2T4ciHr
/uUWQiigx4T5MNujljRRvCDz8o3M/qT+R/955rsWREPRuxa6HnhYUkNfK6j51DTo
YeHmeDr1jNB21RtM8Mxm/rj8TARATf22SwMCNAEM2WpXEFUgGBTBDsez+vxwIKTc
LJwqYjeUnTe5mQPxSimpCtS7ozE8t6VtgmV/zgDlQm8x/1IgRvo23Yn9P3xauyui
5ayRMzNXWT8V3TmM6qCjnHsCypG5U/V4/lQKrLM8Dq+xkxiS5s7W2Ak/K2SGaHz9
4L6AWatyUHcoYBnA2wQIcKCL4BfPA8MJIkPQIHs08bZ5JWLeEfUukCf1DG/w1qA4
pxLxf/LjmNnQ2lEHPTmBAeEoFCXPkODMJNuT+fdVJdtg908u0+s3f7RWMe+CIK7Z
Pnd4nBopVUEZPUoNlnZIfVbyFROlhDvTVvhkEd1GEAZjLKYHYwQkmd24EYzo1JJ3
g0dfA58VYV2VkcdzChwCrPlGf+9T1h4Tw4iS9UsQcNeIjBvdNxBIKMnT58HramYJ
+MXdivD0Lvreh9PpGJUJL/vvkK8nyqJR93j6vTUDz6eMPg9kP8Vv617kLdRySFaX
QnS/EO7e3/8QGt+sA2ojPe+SpFf7ufywE1MNqKSGpGMHJBb0usSeKTuB4e3BTqzm
wEbuiqitlmhzT66aYu/oa8U8bG9oj8phBAB6EGcEfgjZK7Ts2C7Vjj2DNtQJ/L/Z
LyslqjDB4eVQB1d/rZzjaoSYN8fZugqrjTJjBmb3ePDKQLaoibhBmdivczNN1YgG
vrunjajNRqyMpDmzwjKxB88SLsrxUT3KpYtBTkO/EW6yaOBUh4dAcskydd6g030y
oV7gd0OtrCDWke14FEegcsGPGVzyy6bCxypcoa5a2LmMWYMEHab0O5I6sEh56ivc
yCQtF5sZKkyuDblz0nZvnvxiRy+vSxnGdvo/OSZl529d307uo20Rygatp9r/6yzr
atz4adNC4vQCn2OMUzRiVb8N7bs+pT98Qzj33tgDdBT1swPz0wlW9O719iVgNAA/
55W7MAHt70N0D0wq8nzIDlhLCUv01tAn/AKLiWF9Kv1f2GM0s2ifimeGCRzpuins
vCsIzIeI51nS7DPwXdx+El8kZKYcAlNNprrUZGFyBkSQbjdnE6xnA9PLxxn+JXFM
SEG71YbMIKC/uMUm+NeaE3B+hoqKMrMvKTjLxxeZuB4knAWUtUe6WaTU7TAYjMEQ
P6/+V9zAlI4OcfEtB+MGl+4tvWsuUbtW9nhHEFAv5O8a5fMS25r8DoIHXnQ787Xr
raGcHXwdqcXjRnTXA1zPgJ8zJ4gFYiA3YtETueVlf1bQs5aFk84Qz3pBiOPvcPj3
HlN+29MduwjqlumAnCBYndvU1WiLVmqcg9PIphxv3rC1ttHTVW2stXtg/334qI3m
IGXRqFtDq/gr01aisXY+B62RkSPAoMmYjV9H1nuAb1nFKZprgxbOSn4rsN/OEBUr
hlKjcE21SCillvL1MJVU4K7J4uHh3NAytngjU39qPmHBhQ6P4ElYPbFDFvZQC2q5
YoE+XrMMEKNu8glwmKIMbJvzWmIwQuyUN2G1GipKoMtBvxX1hU6U26TTt4QJ9589
DgWN59M1UlLnS4p3xFAxbcdds+RtQdgQrT/sYZmoX6Bi2fEsDK6UiPl01hrq6Rcz
iLVvBMvnPG5n6HCtCyNJ7dJqJLQBPGrxMsSkmi1KdfNIYQ7hjRXUlFu4mPQZljnN
Y446gxVK4VeHu+Zq/KIOaoPDOsyqwVgx5a6V+KUManKGgwRuRj5NJDW/nvIFDijP
xRbs9NWXnXaSF51pjrdsNSJ4VX73JNx1L6Ts/BRbcSGZ1zjTGfas0hw4mbHNt/dL
/Y2+y5jq/53J2QfH7pMYDykQ+T/AzysWzItkGjkCIJO7Sv3DO/PdGODOp9xOrgQq
8Fne924i6aj7QHnTacf1elht31lzyR+ujZcUiBb3fA9GTMRIxI91dnHNsU9rsfYY
x7ErtpK66CMAvZ208S1LyvHCheDvZ+RJUdUl3RY5B437RUiD23CJu6oCwUrDH4fX
L0zcd2ijtmdAmITTUffcklbtVjU+Hk27vN3AnfyNFNSDhtQiZMNhcVWT5uMhTltM
r3f/k4ZFbadOYu7kuoHSXY76/GSpAMD8Ww7PDUwl7bGwh2eUPNBj8rO2fRvXsvJG
fVnwWk6UIpe/CsKHUDxNDzRmZC5kgV2duPMMz7gfloKyFkgpWfBMIAstml66IEkL
4Q7UH17rxRiYIj08MA1i1v8ymoUaUXcSKOhjRPU4L6G9zarN0JJY746l6870t/FV
eZitO6hTn22szoMq3LSHKE6hb2jCYbgSzpe4rHzDYGV6Mtdg9JLG+DTPV5JePWIf
PTZG7ZvgQKb1bFUMPz4Zt5ySHEy1W2IVJ8ZMZdVy3QCrxE3fYV7AIQjqlyj4wYia
rlzh89Klx02IdEOHoPVfrFe4F42DplNsGoHxgGDdzRMfqwSnHw81QIBB92VBe2ps
+ccSF5nB6FkyFJoZ2g+/FHHt3c225dNVQBcVS+cIRXSmGzTm9vEv1bBIiEbxe2gn
Jj5jIq1CG1P1LK7VkSYZfK4qObKBxSCSWIrFQ2Tnll8n+qgQ1aq9Ld+jAbhgM9cq
YRuJ4r150G/wzyD+UAbh0rBAuXSqG2O5FElRCFIHZIL3+h/0KwLVnWkfHibB6UZA
MnEkpM/HOpfcDwxpH5E0YUfbDAxXdrf8C2hLJt7LjjZnCYM0f3CEAVRFe6wKw+7s
Tuy6hAnn2KZ44wHJvs/ewfZrzEnSBIRU7+cWn3clTHo7nlcgRud+mkuM/VxDXA8v
qxNps1KWfyoXAtWMIBXzdYx7jOKI+nuow7Ma7s1zAPXs1hXJ6EZ4IJOOD4M3S+5p
zebJ9Sd0hF4pT5eLO/JBcYbhCvFa3nCrICfcR8EzQ/6bOElBqPMe4Stpdv5YvQKK
iOjBsooe2f/rsvvRMCJ+kHr7IVYovSFmILlDHjuZ21vdGF3PbscZ0eRjpFj0yGyW
VFeR5dBZojWrkOJh4ipzQnLKBv6G0kikjkhNVxKrFTE04QtWvLxizcKS+HZeIkg5
PmK62A1JYuNIMrzCEI8pT2CNhHxpF/dnWcofh1PrtaVFHBIJshIeUq2Ytkn5KdjZ
tHlXuKL+skHwChcHXKfiYi6scV188NezyjgDOwKA5xvW3WA/gbVAF7DUsLGeyq5j
lAUukaTdAsWwZJngYHpL+ExDc11+iTZ7AtZ0lUAn4r9PpjMJjb/N07Hv/2l7kg9U
tBTCz/JMy2KfwHyLN7UwtqJzZ3hR9ev5kpZvyl4C9BEBQJeE9d3Qc0CHYFnUjlIb
nr/5E8yqDLuV52LE6adWy2OVHYEYLZC2igdeW5l6uV4R01Q3oq0lAD1Jto+ue6mm
+vAXbzQ3Uj40JDmYRx+xNSQrOnnV8EnvzJVKU4ewkbhinZfTvhi0Izy5MJzn6kO9
lCG6sIpNUSnIvOz86/n5Ze2IVqcnuOwyxGdq2sgJxpko7ZMM2G9/U3225jQTmPEV
i8NVEieFj2EgEGLfcT3DDllhW1Qt/PqSdRmCPjjmO5zCFA1CrOm6WTb5mFIdopG+
K6YgrC6WuaDBHIvsT8ivJz+/lKCWREs+P1IFBHhkk2x2oyXWHNhuU0/Jy1bD1fZv
9g1StN2vE6ePH9cB3XQEYwjsV85ZUS1QvNHbRpxP4NE4+z+Z4LSQ4j25YQigAYqh
LtAKEaVBiWsxJg7FPNwPm4c52By3uz+D91o3eF1qdDqVM79pwEK8o84CSqHbk7Kg
3IwWERNQpUgvbKAO6VD99R72re8siT+GXmTJ8NoqsQb4PAyUd+5COt2v5GsW6tnx
NzbTgZMxQyoKYEpnZ6WdQrCrpX/HuZ59LvgIMZYOTMLAveFyAiwU5F5GJ6Q4H1pO
kC6UIaW1SOQvFdE/OLG/I5nMd5f3PKN+hu2jAECxLC9aMQ0zTyINcTlfzqd3k/J4
aXQ7sj5qZBnGe+3fJu26nA9+kdG9Jn6JdPLRO/m5g98yOqBKH8W4bOMAsR8qQSk4
7O5rB89SS0G8I7wGhTIrfLzTbg8jtCAIrTYioZSgpvaq74S0DwIL9eNjDIaHxEG1
MkJxGzmrmK95SEtBwsW8ZQjIjiolcFlhNm+LTTGOB3dJHdCgTbzBqrmV3zsy3LD4
eI1xqoVzSumBI5VloBuqHPH+WUvDo4BTLS5yA551ifpsMjgBi3CfCrAfv+vXLGP1
Vg0QqOBcIMbztA8KsXrUvOc16gxP+SMc0k2OxrYzFgsrSbPXouTUru2AOMDjO7/b
cfXzJfKlo7mOHT7HAZvAlux2Q1spJOclYU0K/I7pcsoS70pqb88YNbJ8wJa+XZEX
91jzy/N4ovbBpQRmdRcMCfda2YmmN48OvGVuAYykFvrGAEoSkoCr2wwhvmT1hYrC
dyARjxSkUtkqZoCzjVDQVfb0LNlz6SlV1YQTp6EFT9Mcvbwegfpi97DNaA5x8f9o
XULm4gYLzJOgzHQRG2spPtc4P3fFt9eYksoHctIi35y1AL5bYTQjwGC4AE57yc/X
w3SrezrV3JG4aRinsqWkhlTRP0yNzMigB8DWzFhohBgzzTPiuKOS4FdRkMVsrOkb
ARckcAuFUU2LsAPT64K3CMrJ0T5CQmduP3ybpn/CSA5m9G7OlwQaPoNSlRRgE1Dp
HhmZoPiyMiaLuY18bnDBWG6lkn1BoMmTnuSZNFRblDXrvcIDmZBu/4wUclJGtfR/
YlwaxRw5zV9AYbEZPy7axYX6p8j1TZJeOkqG1HaU0ohKeLRbb9So1HWjIhtjSuVd
A/bx5HrkoCXXokvgO8RPxBgeoEck5/FG+1zvLWKVRxsJJUARoITBeuUxAbxmKvmI
L8AiKr42s//loNQYtXZ1KdvXFK5I7becYE+UYgf/8+Y/K4qLaq73t3aIB2hUO0lZ
d2P3cLU00ySOguTlWdClhqmg++G/WqJbc+Ee+cOdx4L6w32768lsOWMBeMwJZ3VQ
ipV/PVoDCaLBnvp3PHYTSg3/NI3K2iIMuJstE1DcunnEhaL5qM1lPlOT6k3vTDVP
1PADqlrC41NJqZwAP3KvmQ8o0Ba9ZAlTnMorKz95rj/mGN4GEYGQqCVuhiRUGm85
G8hPK8AMqLmTl+paAAvgotZSogqm/Y2g0hnEk0sZq/X22cX5M2zk6TCXJrkHIJtO
VuqR5mJAJK5AURmuJq1UpEscD2aQ4ZM9aSG7AKzeM9K/R3WgZEPj37d68b/joX8M
TwYEmAWaubxdRKqY/ONiqYD0V+cQMbA2njdaroTgV8RywaIN1r91aHcp7G+7LL0r
qYl5ufniL3hG5AMy9pcSWMaRK9yFfYa1m8XZcEBuD5fR87+90Z+04sodiEna82XU
fgZkA/o7o31MtShwWjK1B0nf3hzPC4uCXRBx9HNemLL+lY7cZyZdQwmWCbj2H1zb
nOi95VzkIkUZVCn5ltPuA3lcgMTrtN3ErcTYkqvAGqPDqJUstz/97g3A9XcVS4Cc
5zTWlhUP+PXywNudU4WUBfnk+jwGN3iA2uQ0MhLJZPcMkSv0q2IpIYRbMT9fiHrJ
xgeZmoXPNW5Ns4AGB7N54M0uadagoLDp4rKcOgzMb7O3JoT6mUTfJn2hMdKDzLr5
BG2DhzB2hlhXkZV4nr12THFv41bLcL8Cjb+jXN5fHpt/O8XtP4PPp26n9iAhf+qp
l+6GJYlbTu7SOvZqkn6HfwvCGDyR7FX1t8cPj7+hPKWVacjjphRfeim+9YkFlsWz
+hLWX/t1hd+/EAVY86zgfmM51RAi3hJHAwcv+pLES71GV6tWhRfMvvhfBvO98ylK
RZFYA16sCsJhSjhjMqY3MvOPPLTDj68uywsf4AZRIKfwOUsgfA/n9Xq7wwgTy832
M60j0dFcjpUsQHeT6MrKxQEtXjrxyx8Rz9h1yBc8YFuSdU10BZ/RTFLcwlRTdMxX
t3TFMfEaC6FigzxkameKXA3BmiFrNY9WJeXXjmFoelRiDrGSZPy6TBDCJ/w+GnyI
Q8o8xbZOxefifcjkOt+zD7Mf8zrcAhxIaGbW0CyI2kq2Y/7ZUOxn/4endHWnbwz5
fTYm8Izlo91Z29wcmt2+dcM5wE5HNyldm94aPgMT1et36x4dxNE0FcFTmjkLGdcz
llkY9oH1dFqMpUkNbslK3pok060UMxSvFDZI06bnNsetPshkyG/sk5zGnxYcpF6C
OqqQqq0IWoG0RuAtG6ptpH49NsUgTYRLbFw5CG2iGt5cvtjpIBGJBAii7aSTelA6
yagw9LPKba6X7sFg3vCvAH5SSJqNUTM0n7dMlL48XcymFLn12FVirzuHhKQLMibN
0ct3j1wwPtPijvlBnHQaDPlMeEexUl64X2RdMxJ9fW1QB5BxaZg+L15On4TtDpIY
vLBCG8iau1KzOtu84LNVEY5ST+GjIL310P5GqJhm54xGsa+loPB686LKAYeQHXtY
IuMf2rZqKmDpq3Vh0z+rM73WfmKYcCJyGjsEr6RDS/Cfk0Cm5CY43V9u0kRgXKl1
xrMt9YQwdsXvx5jiUgEbKJ2lxZy1sLsCJzQ5bNEPciRTsf6SBA07L4cBY2BrAuV2
wTL963bnrGwi0zrKQLaUJ222YXIbcaG04p71jNpexlh1eg7cylK845Pk/aOodXer
pidhFCOZCARqGIDtr11vKQvz0NPeSHpUAGdpjmRkv4r1i0udJSqZ326Yi4ZxRyHg
O2Dtcn/RszKmAvVpFcK8oAFpLKzTd9cHYUwW2+RJTmQ9tjc4NDlo3IUqiFARfYO9
312CaEvobWlcpqyntqPeB2GAOmnXsQ0j+nmMHtrm+6NkPJrt3vhzUO0D2R4kmDYU
oCF79zy8jfdgmuf2rilx1ibFcj44ubDpQ8D7w6mLt2DaTa2GSsRwrQ3SFtyJo8CS
ItnZFOrRstqeRHw4DLrAoR/b7vWWm7Cw3Kox0e1JkI3IoZHszkvQA7+Uw1pQlDEw
fRGFXi2CyNnLAPTUxQt7SHrJNPJjexU7/r35036t/4XR0x8ToS213fhbpzlVALmg
zkjeuV/AhlyvEjQnHbi7rvlVMRoY9y8m2LvBOcAJ9fxRU9daPnSWM2rBa+zLvEfX
PwuiPv7jb/aXlV6EBaPoaj93OB9N5k4YwkvvNpJTMLjcafaDT6igjxYEKk8WoOCI
ieIgIjcoZ7qDUg6WrhbShJTtWgqW7J9MTYg81CJcQaai7feDr1I0RVOXpxnhYrQ9
D0xAi6Gf2iJ04sWnwbRBM7abLCts1VU66WNXvyoY6Xh2ZKkuLA8KCoyN5dO6MI3u
RewiI7E/vUu3gDV45DFcZeOyIhA4dE80x4c8bST1nUE+2JbQLJdvJtYBqOPoVyL2
9o8n1+o0wkxU2mWNrO7HymWhiWC/L6a96oNNYN2O2ED95Hd3F5xL6N+SYTV4O+6I
VSOIlduNtrnWO/N5uoJmI7Idy4wtL0nkSdzZF6HE6oGhp/ez7KhOk2asSRHmmO8x
HQS0IozgVA/hnLlN/VY0EKwTxW0y5xx61VCL1iMiYWuz3EQRb0Vhv5O+h6NhASvu
XYkO5yvE8PrEu/TKe/sDyyZHMlHkTseOrICc7ykDMjgDbW+1acccCA4e6oIgIZ0X
H5IqWxX+jphPtG+HD7oY/r+MsruvK8cJkZNarLXFNyiwzq3gwgWjFBLYs5yiqFrC
yeVL1U+alhPDlB5Mewujrhe+lVvdIF8cjIwvirvPWUk07rtqZQJM4UvoQn8gy38r
fXuTYDEY7jFOD1h2w+S4leYUperfxIubGkdL20IG7nk5/puVHCPqla0KJjsqjiWX
oYCCuzcaAaLxId7PfylgqYPsyCXZ26vZYHhzt3hm8Hi19gUEZYWEuV6XtXjHLEuu
wcGWl6iqbe8XgiCnAnpw436eE4JMoJP9DHgsE9vSiSo5HDMxK5ne1Bih4VmbtPhq
nbFyQX4uOpHMQoIiqq3seb9PfevjNDdF6THu43ED7RIUKQsHyNOCwFPn6AB2G3Sw
HUXbSvLBqinzDsYjr2vo19RLxg+lRI0M2IDVwPCHWVGPeFSJTKpY3jUerXKCto1O
MhbauUWPYLxdm0gDZV5ixv3/ygdyrUdMh+RToi+bBIIhA5oRv+vAQLRs2RsC4Qnf
A/N6ec3wp2K8DoOY2momSAtMVvE94hE7ml9RiGkTR0DFZ78X/tB3aQCCxlB7gWWw
3SIO6vYpevul0ujOCnW5fycyPeiFVp0SRBnOWT15o7ER4TNaHRGOhAvf4clhguCr
56oenleKb4vgX9K2LQypijBHMLQ1UrSyxVrnnQN3Txjn9rrn5kpw3n/QY1/e4sFr
BhSqCtFRomBzS69QEp+rpaE0jxHHW7v7hZf8TsieGSh3liBmqNNkoZk/TBH5y6ou
qNpvANLtwp0XBP/Ck1EeK5Z3z6F/i/jSjHmGAXxxJD/5ejtMyQNG9kCKH5Pc6tzz
VqjH5tn/OJmcJYlcfawZ54xyMVYvdUcstZzvT6zH7x8RTt5qwS7LlWkA6CJKx/JI
jwf9i7GuP6PSoHWCqDmXFmwpwgjST1TQqdqEKyZxklLP4OS/PiSVmIgOmv2mNamc
iKog8VTp6pG2G6CKtbcrj+eEA+p14iTpoZNNUNM7vT6HHEDCMnIJ/0oLMWkUAkr8
lmDQPpyRaziCuJ/Dc0AjjLJBGIyOUnr+YBbhJMSm/4C0uyjztqjyom6xLDzs4YI9
HLetM3QQf2C8olS8FJ7wy8CK6ycTdlo0/pLZgKmAGk0wCXSj5Ni18mQOPZD2dHCe
9QumIkTS6ZQTie2bm2P/SK6W8rumr/yUGlCqe8nAUkQeIWXlWWwXFDBH1AfA98QF
qobeowwQLd0yvLYJ6oEmqzuleYiR7SubPHEe2okvd+bactYkUQzwy7PvjDBWrrGb
eEh8VUVbjJUSbf3AtrnnoRFbf4gSzL+uVkE4OUfxW+COqBjP8+ZAhQs8kKh6RFYf
HB3AMsoUeDdjZ3iqlU5DG6QMsyIPqszGT+dGi+aN9cq8g2YD3To8AHJO9dX+UB6N
2EXjNtjhNausWUtJ1MhF/3xSMmen56bGHveHaCp+Ai+zYUHZI2zodh6jv6EmTeZt
AwhcXrwYbDsFN4yRvBbrXD3Oe87n3lCFY9cgPvHV/1sxbQMJsAjHk+EafkxEyNhE
nB513EFYPU011ZmVDBYZ0t+P0mCgD61CyYP4jjGftzOX47naH6u1Au+erHx+uLyj
5uFzWpwZ1gfiwRdCDMueB4vl9Q92baoTuODW7SLF2YR5eEjW/Hd070iTz9uim7RZ
TFD++dnniAZtKoMMQeGBAzyjCdHyEAS3Koh3lYj/hjkCrHWg356cTSrJ5pH0HGte
O2kJTRVwgadprLAmNWBaWSlzfhafREDtYulW+7DBWzw=
`pragma protect end_protected
