// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:37:33 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
W1gVL9i2cxEW98SAYEoGXmtP1V5ZjdXhdA4Iq2epxgedK53vXXUAAJNsKE2zeNAK
mxupsCSzUhUOKjNLnRHp82JMo6jLUTLHQzLhxUwEuEVoIB81eHF5jzjW/wDVdfuF
mg8Xel1PDm9w0+wTNTIE98/jkcEOPjsooDNwEjJFMWk=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 18576)
EclHQUPfBQbvEPql8N7M7HbDbxyWGuxGFOWPMKU1IpDxz2iUU+S09m4mMK0bwcKU
ub7zgZHz6FUAkmva60ahsUdHUnN2McPZHLgMl/HK9jgn6COFyzyHKaeQzECqJShw
KOAD0c52Y3YrJCesRc+I24khjynZilmL3FCbdC2icsSpOWR/et1x34360LDjeruj
SDBGkgN60KsvGr+GBKJCik0xYG75YPulkjFBGURMTUv3irRHApb2+l4U/MbmthUC
KOk7wHBUMbMWtY5FYSbnrJaVFw7FDNUhEnRwK3mml3Yz8cmeP46u2A5sJ1diYgPk
rCTvWmL7pLz56Jv/Zbbvvb4CaLBX/mGLBGhga21WeydkuXIHZyMA9ptlEviuNKbX
2bObh8Yy1dmxxjxKa9JnChoJnebCv/Is2S4YbI9ie2SwO+ZT1/3+aa9HD0ldwpIJ
kFhrZNV7YvytrtlBr4ZWM3uBsahV/Vn0Kys2dU6izTQksA10r5vV5nPJphZmrZeq
BYPn2DtXL1zczrJMrNIIa8RFD/JwjxIkjPezZErYuZJcCTghimSp5DpqU+5f0qx+
0bqH1DNoKShPwrPeQfdGwCDVT3Eq1Kx/cuj87mXaWkEavvtklMVSDEP6d2gYCd1R
T4CSv2BT+MYh/8OkdVIbAtptp5QAuBz2VPpynKm4P7atQtpFB8cCD1IVquDrrTgN
S1p/g2IrhStSRnKY3XvcfNiWqWOusaHs69PKJkUkxqwtSqa/0hlE8RgfIqXGZPQm
CRWoiWsAQqhvm2AUrMgHSDcFavA3DCOpdsz2vByiIA+N9vslFrFuNG1oZ0D37Zhb
r1m6IKz9sR/eggZBrXubCs7UKFiP4GlfVTiq6sxDOvefzKdbAynthz+hyqEL29N4
coLsYYxaGB2IZ3lIrlDcCMK6scnbiWZSDJPy1oYDBIfkzVbPAQ+6lUOPkKD+dIrh
H1Sa9A98R7NuqkIQ1mww5S6xUTqzrXx60vhvGSDOKUu9pr2Y9boCLkg+QUmwQ0Dq
KFgGEPNhYxhtGZ956RrmJmhDpbleoXf9jAGgBpsufxLuoDmLfzxXMpgb2WtXVtrt
msZEzc6yxniVHGSMNYeYPjGIegjH8A+v1OnUdl8XDNYlrx7DKoJBMWRWHa3beZfn
giVTT2pB9eEbmUPGoR9FfV29Ht80r+GI4i1yyEfV3/NHeKSPb0I1rXb0RWfN3etF
y9OF9sdlFFAiYOXXRulyCdFlDm9srydvT4RTF9/ChQKtmyEiRbaXG8cNOxNFZu5+
vHv7D/n/vJJKcTQNMyPnPIaQ0OnSHf3w5w7Z62R50kDKAPxEooNxJW5Sabtl6Fxn
6pMYZNhR//4yT1JD06l66vgzXDOyTdCI/J1vZG4w0M4TQiJLd6mM7NTpAvw6tRmw
4rPuTO+fN/KQuK4KgIMFvGbacmNyCejb/uyzzg72esJlA7+3qrI1F3L14rmKSqyZ
B6YIzCmjp2TL0pgsdz0AY1xfJGURwBoJaEAyqTs9R9JE0uESsbuQGaMJXwPS/nUT
U5cmjN6jmDbo5ROLa3sfieH1pJnXkAwhTevyVMnnsfIqY4q9GIeitsFB7jsmemqT
8BnYCtuGzwnBo+SreivpWhgfKbv4u/+H+n+pkmoTRg37k8+1K2YiGTasEWbxTfpj
0hmDF7yXxgHWHeYPkWQo28+LgvdHy8JVdZa8s7pqYstI7QrASC7FOlK6KCvnlJrt
hG5/4i7LoXqJkxuTVdsnrYBeMLj1O8PL8ERJ1bmfs7eXlYtgsbCxcv4qyruuPvEC
uXjCfK/stznTIuL5KWjNQ3LT71eEGzGIEL9Zo2RGY87Jfsdw4ZkjoYIFKpMH9Aai
vtbaDSsx9yM/vmiRGLzfg6kt27OxoQJCJf5DjBRKwTIUQSO38MQHj3Gxb8ia6YLH
LcxZHB6Nj4Kk0lATc92iyn7jIuFhgzzIKGBV0wx+OW0DYN4jq3WgV5jfAO0C4Rjq
YWS9kdlTBEk6oWuZGA1y4mhjxbIYaPgokdiZZ39D2fR4CjBu2UYwTa/yqonqbMBa
/SFg8YiYtpKg+pAT/hMwrmvTRuZux08jUXhwVeW8lSYL6LpuWqp78cUXKmuuHx34
Q6k5G12xvYPOzi0NdHCiZMqc7zbcIu5PkMhczfeg8JLkNyLM7PQ1UMDdgtvBdxI1
x/WsqO4Fzqf/IXGH4szV0JSndhJZaOWlk6xtPvTAl2cosdElywiBYeYAzZMFXNtM
/BcOlD7HazdH/4YcanHvA907lER6hn+cIM268SaE/6vLbvvcHG2DXV/qPuDLVkWy
2SlZIDX54guHXea8euGEkUsOtgucj9EX/81A7uB88ORgKFsgYP0xmksRQtg+bMtt
d6JJKlg8Y0VlNFZBvPE/DexhC+rBj012OVXW5J2XUwlIGeCD1KquOvddlhu6Qt/4
NPeZM8O2khmm56chtZMPvbpM9R1PlTFh27NIfhU65XEeSof1nORKXppS2CYNdT+p
Wui8x+UADowQOjXVldSyrCfnwv4l7CZyJ5t9dnYE2NemSbu7F5Fg+j9s/HO8edGk
HcgGT31xJ7M8xICxZpKMK3pix12cK7LjtgE2BnSC6hGxI3dkQYSe7thyUPExgGt1
MZl7vXLK3axS0wHh0s4IMTikdAKsPoZ6l1jBiXiB9GZD0zWT1uSpgHD0kgIPcmdE
t78mLZHPg1A2vFb/yvNf7O3YdgSvSnbCAqSnHzcaUE+mPutnCmsg4XnCqsZLgWwq
DUigDMJRcwzHkxS/l5gplzQZbL8yMNMT8rJgGa1Hih0rNijc+TqA3bqxODDW26WV
ruByNSQpvBxglOXL6lxzeJfVdG0QauxrRgvm55y5hPilQr1MywfiRLHwg34/qPf4
CKwqAAk2Q3UqGXM4r4wpJQIapZCPydPLLoWACF1uFbGTKJVHrlEgbRJe5TnaztV/
/g8RH5Rky7BQks/Y3oyOq7zvzdfTZ5oCFrZ6aMpG0XOkwRa4JFPVYeD4ew10+rd+
FzHR0xzeYG8g21uR5OaMJ+1gpbEp3jFxbIJKGf8NhkuG5mS+MAFnodXOoJolVz8n
X5LxGPgfYtSk5WnUMY7P2WS3FM6P0OqjB3FU2/NpbKPuTBZey9SgM45bMgmq+u/8
AyLOiu+NCAslnRa9GScnKhi0XZH4tGrv/Y2eExAgwPXDG5DqNAPMnOhPQHblfLrM
FR+7z0+oe6Qcb3FhMuh7HJBceQY/s9aKabuJILOPNgvJJ91IZ8enVWzrtDlfh8HR
dkZ2zXPLLQTZ4/qQ3NkkqjUmTAEOQ08+c2cZLiq/l08I2OTisyWesPDo+SuykL9O
kGwmqW+EdltXwyabwsnLzkSUUfpAf0qCQYimEvsDiOq1oJaLLgNqshdQemgWqSsK
Yl0hvp99a91COHWHOlGHpH+gs7/tG2jpCS5igYu+os5ySy0fAtxqGkclJD2O/z6u
M4yo+j9kMC5OgsuyDHtLMKfEdSLacb5PjSQE5tqroUu8CnUtXEtD0Z+KaoGBtEq6
jLFJzWlAW9lGynYsIXYZGr4mY8r7Cy04VqbbS2yiJsWannUzBst+npt4jwdusHuV
RHTIoPLeHzLr68HTCB7jOmbtXxOhcpYEA3q/ZucT39JPIId50eKlcsRlLVfWL4tv
dGvlJgq93r5aEmQuZ7SwDv8iSqx0evomrdXb/vXCTPGaCNWkVOslt89ztROk9n06
HOTxt4M8SIJFrHx1um/Lqnp2xLfRy+7FfkswO0K9Hx/t/ESCcujn83GEHzxpiU12
jhy+zDYJ7jBW8ny1QaVr2jKnU93rAUeGGweOGvPPiM6hK4SDo0TQfNlshdqkNEPi
iVPt4dEqIfreMzJZpCIIfwwTAkuQsUDUBYmq4J4Lfh9oexUdNI2w3UlOiGRPFKFx
KfiCPlna62xSQa5HGMWQF8T7T/C/lqJ0lcQQbcAPiF6Gc/DztLmQQxaDPALypv7h
Nf5lHfNp7qDKwMU3PomRO2UWvt3tIVgf+bvXbrsLq52VZOsV6nq+NcdpOukFEvD6
a0qa/skmn3IXsWk821ZgDKU6pRr9dS4dMh9/FY9xBbjGhOLO76fEg1l2JYBu5Xb3
8ql9ydqif0tlb55/IQ8QQL/snz4qbCkbKisYHsB6wUJAcNLz/zIn4XkzpgYSOtoV
Yxda05ap2sSLTJ5zIypxb0kfHqgoin+WKDbm7SI8FmE8vcCvDNABqOTGUsJiu377
VJhKwE9fLAuvYchZ5go/TJlI5quV9qrCFZ9tsj7qe3FQO2svSnO9xAOTHv7ChQAL
v8xnB8uzKu6GOxF9DLdTHCnmv5BloDZtUYe6Hsk8t+BAc0LoNMweRr4mCg7QQIzW
W/4bVaj6mdHSrYDIcFmECBDthVhm19GHTJvG5mEpERr+cvCmKZm4eixdBAnv/Ow6
PYqiHX/sInr9CX43kjzYsFPLgcRHFOxQCoksuQhRbwbdefKExQQ4xFib2lgVScIB
kMfufzxrLl7fKOsEGJ9sJAZAGsaOk1+KEZRX80zop0xsKewM8FUdxiECNd3pNoii
Bampy+qmKnVEkKEY2VKdhnURJx2Js6jKYlniBbRzCFwxJjRtND/3eqmo2/NwgJfh
xUYdn6CYl0rERCrV+IAfDrIYElakU9R9tgWRGs9Cau+PpurByIDfg+McH92l1B6a
wmPDPD2+llhB+emTRDA1P1BZN3w6EK8DtRZtpgecwbVt11KSLWsHhMhaf11yqPiq
4nRKv6F3EiRo1OvtbVEFChxUcVJdi9/sM8r3NWg2aN+fOnOxBbSBCYRaqp7QcM57
e4quh0Trj8/TPOyqsqSX82AWZ0BefmomBKvaNqb1wb33EwjY9kOMF5NGVrZ1Wzs6
9OVk/V3xSBqLYlE5iSGB7kcitDvunzYsfAKCv+Uc43T+hHuoTNOTYNJialu6DUIZ
z2k38WnwXPyA09icNuggBPZTHw1YnrDoPAndGMrs7cx6hwHogbovvXukuQ80aCaz
CK/o4LZEdJ+MVuzaiCv3dbBHu+KcZxUD/HYUKd5/DjZXUOdrKYhDE7gtFH2njDJZ
BlykutztHB0bEiIb2JqQfS7e01a+U9ay/2Q3SUZx8bxDjgkYq1u7ghLyIJSVaOT3
f4svw68HRFFPHgYrO9/1mf8HXg3Yz9ev5V/1a1J+eiss+JEhd1U4Cgc6hSuTeQtR
uK8LuivQrFgnYmjjBp40n0oI/wpY8oPWfCdBdt/oOmGDmiXjXZ3ucS3UkHGpyi7Z
xO0bbbvXrH6QfCGEGzxBdJzPjT1bG/12LC6U9UuvnCnHbUs6ZRT6FS2Nk/tCBApu
XKGgGuBP6c/9VWLPE+2FWbVlQAFjjLRStJdRJbfEws/SXE+9Yiyudgrdl612BFQ3
w9ozM5bpSW28vxCDmL6BTUt0BgcpRsRtkRw8QRWKoJRjxT8IOnGEYNBMxbK26idv
+gWjA6nKN8xhBorI5rqyIK74thYSiPhGes3dqqmL4PeSncCdcXvZ4Vl7GzPvGraL
teN6LfqZ/g3/+vvAUSbLI6gxYNEfsLCyjr1oyvB+OE8NTnehd2Id7/4CV5eLbqg3
VljWU59TKqKYq3l0eb6TP8F1O2n/Phb7xVoJPGKP7oK44on/QJZBIDPp3D2Y/NF9
qHLmwYYaVdrue2S7VfInD3QUh7hiqinvxQoROmcXBfm7GCX9T+DEF8swCgRKbtKG
XG2nwxxfMzI18aNI3n+5BGAv+16mgTSIRJmq4Hfp63IcyRzj9gXGSYwPAO4t3aaY
dzPK94miKwYhnQlwaZQCDJZ2ffx4axQ2mBU62AQ1mb9tATy0U1M6/Tt3CW1jkKFA
MPi7gaX8qOJQAneK5QBZQbA8yYlweOoKOZoruOu1Ly0VI2AcbxsleMtthjdRsaQo
vT9/RqDQg+rZrBodW2eE/ebTx2tjmGazZrzHtRyzu9YffPpDWpOAhM9Zswg75rw2
bPEG1slwc+s1pkBcPP8LnkIzC6F65XAOscs94GNiJNXif71POAw3c0YnuowWOZ5f
BCpbz3C6SxQBTEnTlxRv+ZJ00O42OsvTUEDIcmlflgf13aVI5+ufzG9doSpH6r7G
u9Orj02G0bw8MFbvlyljNn0mYOuVPtX+HYmB8Dg5/hap+snhPPnyrS8LXLKf6x51
DkCDSP+KFZTt/r6WXn9wT2lpF8F1OcpwNaoGP6LYc5nH7CvX2u46jYyifkND9wvS
yb3vS2kESzt+Dn4bXevOyEBS0KDlBJV2vk0/iPZQYCRdu3IRRWMPU6RWMeYwhgjy
Qo+DM16agBGxai9uS0qktWUnCJEFOgB/iCaTcnN119CXmhUZN6YxhIcqDa3FI5/i
QFlOffRXGq8bZIhY2wX5VbnZVmGQI5WXUitzCy+9P39Z45WPhwBzTpVTqAmhu+W3
knrKMUyUZRJ6zbkW7lmtvTnz2E2JBeSYXrY28WlF0dc1gdzprM9lGIe0tl9J3MaM
6oqe+3tDRmMDbanoPhE+GvajgvrgRFBJjdjlNDvoqA8LjZxdpkLe9G1hzMVwuRRN
ZrjTJANgBpDnmKeOcikCE3WwRnvEAAiIQG9TkuAHDc8AuGOMDQ/SjmjTZFRJVyjg
/Atj9YbSVGo40R5kiSzgwc+A8UlZy8UiSdCTjP1oCTv15rUs9GhKJydwDgLhyYHK
x9QJ1Njtoww+THEY58SyPPK0xpicocQzYYA4Y5jqwMz/2LGgEZVP+wh17LQ4oq4c
JepiUIDdZYxO1G9ALtEXOlkFguUnRrvhLzcCOuZ+yG6r0+HmqAxp8PcPSq0iOrOD
n9fbTwxvThbaVttb9jOcbNoYAD93MEFL3gohOjMfv4xYiLpYWLlLxVNNpqQb1tSy
Pyc5e8fdfeoOC1vA24tFyrdsKR1VUrv5uO6O10UlQ3DP+e1KOnn7gMWz1YHSnDBV
3KV+MVfGVPjQViXT0suLezZRBt4V6Z7wxZ5yZM6lWPPhbQNHGSIdnDCmT7owGGWJ
+WGtFYEJM5k7lAr7+6yi5ndO9yKcQCIS/0+9KIrqxTfNWvoeC5WqpJz+PXnlWEEb
jSh7A/yjZvSik+C1NtYAuzpPSwTrRmjkjD9B6XciPEIhiIQMFoN+Hip++A111T4R
q+7f+cxVs43tGkfXHTfNJ2Tf9FyxqqFjcPlfiGBLDv7Zvp+69MVbCWWYLAtgbdHK
jQR8FL+G74jp5q5oA2tiJtUIUkfrhLXUY2xmHf/1QMEPAq2eW6cWcUGO5+a4Qpob
msXNMlXdUuQ1AVikUdkv5ChLj1lBeF/eRIPvDBOmqOt4bhZBT2v+tftLut6nsnXc
sFe5yaUSwm7Dj9W2qfPUPfAawE3rRWq3iECZbvWglNHSayDOUihd3v6UYAOdAOF3
g76yABgtUY1lF9NglryQWlvveRmnq82swcHYdHtX3NO93b0tMYSOcwTao3rEpA6w
wvEiiesTWCh2zv++iT7Y9l3lYZdCgxJB7F9pPL+YrKIuTECX4bwu6Pm/AYJDY4nH
ShANFPT5kf8bTvVbBv/yZC3h8ZiSEm40JUOpQbd8VX8CkyLM+NPsoXnK6n0cBl6j
e2QKwDyVw0BPkgsWl+vWA36aTw70r3I8uPEhYNfaWXF9YvHwstjG+/F8zJ2fe9LG
F3TMpJrdqvdYKCrkRuyOr5zHJZqGGPI07P14uAnKZOuxHGMstVGe0OSGE+RIvj5T
Bu7fW6z50JDMrlCU/+xEyxi6hqPT2macIT5xYZnD9DHlphuVEFgOrZCjs9+3v7DZ
is100M9ALJJILaQNhpYZMPCJCgHDGcDiJFPlbuoUy/u3QsVE7kLMI+uN2sPAUbLj
8HjhhIhJq2tI+yz41Yv9X2LfbMjq2wxY/57MhlCrYoVoPFnDNYm9KVgN0hrpmMGg
9+3B6UevIJggQCnNObsCDDnxL1nFfE6CwADvT5t2PIrSGSsE255VQWX5VY7g+4Np
ebL3nIrcuP9/Qw1dUUU8P5CCiq45sanZKNICO/j4N9fljHEi39ivtJaLtSFX7vuA
VEHW0HZ7buFdYWcDVDyjyjN6PrsFZfpvokByOMWZaiosGRF222feFqbBtK/x1Ha3
Wh7isdCtIGH4/SJCmodDbBYZI8bp+3uuIvtedGQUZXpeDcQWw8FBjHHlUw9MuF3w
ZhyawOTrhbGkp1x8F6b0QfU+jGo0Px3TL253Ayrjxi0OqnI9CdBprZscHdIg0KhW
mjXnmqpuuT2dpaS6CnF7dyOe4WAirWbPflPYBuFkCDetrOyI1rI2j8OEKmFV2sqL
IREg7ypD/6xKKc+RqHfKPZLP5iB0zj0GWapqkSNpk9I/+HGGi/3oEtUPvsM3l4q2
eY1FN7lWbRcXP6vvq04T1Y+owh6TGbjdCPXxpZZlWrAg1zo1EvvRBp5Ktu9zGPUo
8jFVY5mAPDJmcDdtixChWPC+VJKnqneTu6T4Dd8EjjfuoObAqAIFOwvnY+iuqCqy
geg+pZhKZLjhkT7nj/QbluxOWm+vtXwIVn1PHOSIPLkA0ukSrtDqlI8MNEFpfGL3
ezDVBYuuM3JlvpSn3503S9GX39IAmzaFz4UGVMBcTX8egakyXh5lpgYhg6harH4r
LU66NgomIFPrBf6z9mD3lrzR/1PHOq6nIjMLkdpApV8eJeKrIuDg5aDsN83Ukhne
tMoOqy8fbE5sEm7YdcIJXye63pGDpTkbHa5felihT9l1R9J5vUZPUY8lZtjMDMVh
lzv5NwEbMqvPKaltBCQCd8qjRMJtuMTSUoIBI1oUHobxopcK2+CHBJvuhbwMvUA/
ShtdzNswJrZy1052pBdG0kLTl/hrdT6iXGOcCC3Yf/PZkvqw2eeEwg+wRS/Cno41
SqDYQr+M4VylbDr6ZBQ45STjkBhQnlMl3p1ovHU45Bco6Lz9Sgvypp/yTRwOvARo
3JC+HnjMlLyUAdltww1U68UKADrhiTh40PIjCPXga1M5uoAoqQsmPfKVFVppRNJx
7+n9LFse+e55W3DtfnlPHvbA6IWalhpowqH7fEotHpoSl0qQ0HueKNoZyA3ZjV66
n23wx9YIc2yv9HiGGLyl35FRryJ3nAz8mTm4tt5CRPgAbOSO+rBmyd6PFsL9Ry5w
Jyl/GTzYt852GTtmfZUzAq+qa3bh/Wo75st9NosSPZzhfjIGnjlskmyBOyT+a0/a
phYGjvdv7hpDukoniaANLnVKPaN1PXqId5S23mpxN0TbNXCIcBw1ifrb3Gb8M50b
LCtdoDP3Cln5q3TnO7vH8YCS/emRfEAtBULyAFaKwCM4jzB47H1xOhpASw815SbY
msm3cwaoBfc5kxEX6Hvp5542gjbeQgbJ8U05iIjkQs0oy5PzjINa4Ah+E1CFFS4V
9ZoOe0T21c/1Su8kosZ7W9T/Ed5uv2o7fNyKfagEtd+13IVnFJNa7l/Hrl+hByNR
MkCc6I4K6Wg1bIwW4Ijyu7MX3cRnNczQ7lzUqI2CDOLxKIDr84Y8b+XDAkau8mZl
iKJoRa051luwXgYvETut9NYXdnb7GYIumOOYw2MctOChP2gHvm6j+JuXbV9jodST
ubwZEefbvihwPwWKhTmoWcM8LUKMWH6WI33QoXhnAq4518mKB55Su0iPwUA6f2id
SXJM3qRQbHgh9wjZSbyT2ixwioOaGw1f3vlklNsmiTooEIgs9DYgYdWoPY0AcUoJ
odyJWbUoxFkivIZ/LxfP0ULal8DFDMO8gbxl5ZLehfuh4tsDyP/1T26RDIP4n4q6
lOiZEL+BxdkGSV/+utkPFCbvCDUP0sey2sl2NC+yTSb34bXqQ15/UB6F/RdlNxAy
Wrh37mlE+GzcXAvmX1b4GzhM6a+nyYF4oU8DPOz/GfOHwG4e8UhWbUhDj0VgKGNb
g/MNhjkwwtAQEbjuRstVs6u0ZIJQ0MRNfdqU6m4yPmwGs+lYzb7Bywu/VgCjixzA
bUCZJ8BkxwhTeJH9I5TJ8rdhSzAFuY9JjXX/+DARpRU4p5plh7D+h5qTxtf7BuIb
Ii4wUQ2OdCIGdMEDCcY+lqPuXZkqJuH/2uy6ezKv/r/jeem9XvE2Bns9JdLLm5W1
spetzY708f6gWPFR4Q6K1EDhvMRKKRpoJGw70GAuhOInOYSZkuNxQAPNuBeiJEYn
ZJmXM+SQgvTSDgIE28cl0KPL/MCnvLtvbQJN3aTG69JUz33Wi78/O4IEikaaWH2K
OluDSdMwSdD09JpZgjKCPSCWz/aNTbhqB13OEvhw4CgmwRqKRFVe2lLfJ/nX48po
mPeiMImRwcElbl7zEhhhANhQ51UX1oQ1cAweK4nkV6JLHY6x7zgJqFnGq/DhE6RS
E5tVE8SVvFeyODs6RhsUcZYVALUuYrXQlMso5o7kR99RALz8wBzUhAjY9wGqfYA7
y5mr4dopxUx/MBv16Ld8pUNILaoEF+E101CqvbvmAccadmZ6UEK/mtpkj69JV0g/
C+QiHu4AqxHQzP4rctsFjhiKa/DbgTVata7VQgEe2+UtjixJSdKGlTLBjXijBx45
5P0gndsbewATK+7CM0K0qCzKkvEaPCmKMisJv3YZa/HI/3WcyiTF9lrXHL3hgx0J
eVvefzyp034JhDlKFG7zU2zY4IHoogM/wOhY//8ZDF3pbvd4BuXm4QioEzccVM7d
KFo1ivjhoePFJKLL4THMn2pGDBWBPqlqeMpy7h72bapOEJ4K/HGYGOxKZKdv+LTT
x+Fdqd9nnuYV2FDXJ5Q9o5oIsX75G+zZWiuXKCiG3Ie9Kbx4lQrzd09fx1RXfYc1
khUI9tgmNB73xJfa5Rjg01ixZukhlF4ulptKfL8ZFrw6Mxs/qSVbkRshIOF6KdsG
shACmtA1hlL4AcXWLAturJ3miXqzNm03rkTR5EA1ixJlT1w4bGIRg6SLbJpOB7+C
VTIzoWEQVO7QHundx/Nb+iuBhnjJwv4VlZfeACxnx0yu73oS2G876CFy04a2ru+i
OwqeeaDlJMGN1CE6nTE2V++qOE6t+62APX03nuX6ZhcGDKsWjZeYjthCjNILgZgQ
FJTaq8g9NaMvxp3Exc1UQgsH2z0Rz5b21h/Xcl6JTzrln+USDZdO0BPgLUe4w0FD
nozj5hEOyj91G7AeHWVj2YM0xkkcML0zcwN10b+0nEznLFf0iLjceuUGJFhLz44L
97WidWd9xA8WBEXMskA+S/glpkI5Rx0BQLugZqsexOLDy3Mq4qw+ypg4v8PC6YWL
7i6Zry/8m4+BvG8PARs0oirXaPlpCJw0WtfWP6eT7ZTjwx5pcbfIon9CfEbUjkYC
hVcypUMLMxRKW/xQwb48EEV4iRmuNvt+MOb+On2xfxszX7eOzNlRrAS/WxyNcJ06
1+BsfhYcyMjkM03f/hbjOk6N0YQTeOsDyyEg1E7tBZSBOSvwWp6JicES4u2JiBjY
EIkKg91oAbVFHHFZAczt3L+4gs7CEQjWeEZbLUFwyb3WsHXyq3ZyHhjd+kQQvUjV
SaXgKPXKCCWDncq0BN7rZwIhMp1FJHCaVyO7eUjHdjh/Bl5E70/7XgkHHEI0fbEK
c7RSsKjReb5LpDcXqg00rIPPSw5dts3/eua8elzZhMR5KbCgkGqzymeR5qgHNAKk
6QMIyq68asI2ON/zFhXQ1I4GHAb2i3M8TeSMDQjJUu41M9YiZoXervYCyHDHkMDT
sTLNDw9Z7+b1nr0EqeHbPUmi6W0L5MG+TWk0+1uJG9Au/Z5Pf5YTQd3Nx49PbH/R
OKY3pkKw6G1x6HoP7bJbXlqUGcl33jBJDhkZJ6MnqRrXuk+Um8KVfwbdGys5uqfD
KsooejkRTQhhO7AwVWtygjegPndRPZ83h6CS6Ok5RFF9+5MJqkN1g4Y3riOIukFo
E4IBu8pBStfvJajuWJq3dSfZyLqRuYM7e4AZ1w08HEWHJQ4C73WMvNp8ASE4I32D
h8EqIsKkXjQaQqN/wm9fcG3sN1o8UP35ZwD95c6KffB800Lx0PKUnYKeM6EOQbEf
DMRQrpiF+CbMEJC/cr3zwuHiu4A7AOo0370CYDnbdxomvDwP1VBWGyaDUvPRvwFc
PustFZ8HRA3KxGTGdgff8QC50teBWceRNLOmHgasNJ/Wk7MT/LVGJx7ayVXfMNRu
ueETJp0l67L3dJefs7QgVyDg3fhrufF+uUB6Pa4HNpnhXJv2U3D8wpcNoIMEmGeF
GXOz4pB7wMQfoXEfGM6RllsIlf35YYoB34yQiWMaK1bIBU0snL+EJk9aV2JaWjpG
JfuASzDFXS4TQA7B2FgP89IEUvn5Bf8i94ETBO4t7khuiS28qYalywBu3MVhCfCq
BFxjprJxaL0SZopa1l6xdh1Uwv0DtTkoUhACxgLYcM8kMoathGNqLyt/YqSpQWCg
It4n+/xzPKJshf5ypvOANp0ul3tTm8Jinw2E3GlQIGpEESKRCQwNxDRCX8KDTuFG
7z4PZD1qAgJyOTAnn8vc+MMG3vZMMT9iIHX+KAp5SG7+DlBwxt6/dCcbeyXp/s61
hObdCSPJFf4+XgbNAmL1dGWfOU6tiQ4kgwHHJcdqy7LQPxb/8EFs5iwEl1sKryDJ
D3YDKrEX8lP696HyvfhSLDFbMdFsGmhqVDPzzvTzOugEipIqx8Rr0NM7yQPqvn5+
M1oi4cS0mWdvxEOGwaIFy9fVTS9qM+6/CeAZiC4Ex7ZfTj0yK+WSqGLd2e0uNFBH
Y53A7gv6dc0MnURjm8X/iY6a78KR2bzeN4RuYQXIKqOTFQBo8ahsfkzCGRwAzQYo
y7DpFiPnuKFyetH2d4effWS7RzZCImoNc9B2Ub28/3GKBSPiaOg7UHRDAxLy+MEI
1c3drb1O7+gSCOPBP52bvWhHn2FZUmked/BCHaD02xxQzWLCGl6UMGzfvCpWfU3j
IsRN8UkiXIdQxRw66CbXp24DKNPO8N92G0A/xZvLdcHCy6zZELY4vhTdGZ6mjQsy
N+Axe8DdshMHtETKH3gMLKpOUrUerLm6Wt5PZo+0thHHD9fqMdLsOxOuobGOz4bj
3UfyyQOM0aBsBiiGAaSDyglbdgFxk936hh3ff7lo/S6O2ob/MnUiiL2XY10Z/8lC
u9iWpswKhc8XkEuJicbSFU/HoPud3jBvdpqKWKEHigun0BS22m8mJZU4YEF/ESrI
9zfnN0xbBDlrlqlItk3Jglx6H2qyVxqqae3kceJ4EjpFukV5OIIg4HdYZC5LVMZL
gKKNfHD7dYHpEoTNFfco9wxCFEzg4X+SEozsHU5auazRj5ma+i1/Bmx8SbMvKrmU
SHRQpjN1WaCLHubVSORduniKpvgiuUl3l423PqxoBrwcA2REDB2uKiC+BTPtmzmC
ogCpzym4wY14WDfQkkkHvNPF74zGqpnoue7mf4rU//i6U6tySsSQUmuTieKk8GDx
efoN9LKcqmxvGdlL+xuc1soCs8GrNtyRRtv7j9qYJMUN9APjkirPj/a9IdqPo0eb
VQ0QFKlQfzJASRUb0xsfmJ5flc6/JlE3IdudVPv4jZIByx1P2TaBBvNjBQoXEUmM
zltPW+KC+XWk5j8YNEzi2hXolqPgH9ILqZ7TugT4BlqozHms0AVeOheHoM0u4huF
FMiC6Uyn642K7uOvnGmsFWWNOA1EAQBMNnSqJ+Et1QJUybL9nymeeMChtNjqyWWa
Wq2aFz6FHRhXDKunopK7W7mbcUxZwLMZK6857J1cuN4rmdT+YBGg63UyMWbuCcZS
ToJpmrI9xxV3dO/54IkCBI6Ooqa1te3VKUx1ltI3LvG2c8KGeXigW2UYRXKPOq6v
6qiw2y65YhtZvuscWo2838Cg6UXN1qazgPt/o8UlCuPpSfknxmlig1+lHQ+bqt+N
tBNhgoiKvv38E0GqSGwQKE6TTea2JoKWX3yFKjswu6gnaxCvuO2gKbHecW9lgwhq
nfHrm75QKdTWvlJDWBV454Km29kpwWkP9wdaADTB+JvmPPS2eSPcOD6HLvSY5zlR
zJ/1q7E+BbwXGUS+o14ubyAxuMZD7a0zWxPwdCId04CzC86ckQI3gbs6Y3CEuFrl
NFsLMyIZU0+YrIifZrUat2j19fAotXzkO/bE6zjHSDctTEEfYIZyiA2PqbJ9XGMW
mgo5KKRHPiuNx7F/URb4l/ayP2oIc9/dR6xCu0Bn9W/TGACPHItmVpq3Zqo1Xf2L
fRVDnZBV7LiFGl8RDXFXbt0gUATVsqVAGpUmpSW0b6YwtxbESAiXwHoL6DWCUG1V
xqaS571Ynd3KEbYt8z/BVOs1wRuMXxTNQxI8HDTFNdlIhOi7nDGdghFxPPpNWWGE
Ja5cJhqV5Ow1Px4b1RxUMSAiADNTK+mAtiCD2VkWS5Wqy71LegSkPeOEPUReFDrq
wgTAqFUnHzWexDEe5xZmCRkp2OW7gwbcs60wENzVFzOfdKvPDnYk4GQmyyw1hzuc
Zjm7+aomeOe54Q897rnBkWWpHVojzF0u6ltweqwJk5sGaDnyjfHT0zc81o96EoA9
ZB61ibNvDnaYdO4LNMKEyOlu+6gRusc4658xAJe4dKXy5hAK9xu1QI/5/OP3xLFn
5sL3mDkgJiQKnyHOrp6S7TA0m5E4/gCKDYsISjpjYSQwBhhA4v2g3UzZODS0uX+v
rPNM1jbeQ2O4bSDtDHcFotwkC/CYL2/i8TLlg6N3g978aOSAeqaQ1/KfYrmMc3e9
XndTdiyGwhNYOnUn6riauHUONsGYTXkPRo590pqaYvvZ8N5TsjdogCs0qGn+pI47
53jju/d7WMm2rQFuSALYEhJPyjpZf2eJz+RYxNwcJeImI+Xl/S0pSwnWJzK2D0mm
QOPe01ULjW3IpCt7OfE30qaCPPpxgJ3/rnWug3CS9OdxDWMIjBIs44QOmCC0gHKZ
3yykz4DzeBgR8Q7njJceCYOXARAq66UGMAiK0DTvocZPmyFMhcVHc5AuILzyQkiK
dIjg/rJZ6npQmlloRgknsvyFpQahQYJnrKobSollLHd6a7JR+VQRvv/i6f3u/6nd
tnNoNgms9ECjI0EwK996EdEWQUKaMGpmRA/qj+g25CsoovCAdP+1TW+X7wTu0KxL
8BeJdOoxEcTnuBoY4sbUDhepuyUwHnSsfIx+pj9PdYqCz6Mg6cKZUptEYoewEgQO
FCnOu4tEdy2YjiW2VTk7hK++XzrR8CRdDEzQubgLmqCVXhTc6/bfYVo3bMYsr6l9
AvFxYJth4VjUqIFo8Jzg/utvDJxgFTcDNCJX+Yv5Il+m5M1DnMuMqJ1YLQBqM1E+
4RKbjNACw9Okj6zXAiPoZsOYk6HpL1bIfk4VWZmwO1adI60yshYVxqfkWzxs8Dyx
jVprSnyQTAiAawEGLuzO4glQFmrBXGi8m2T+WQw5wjEzwikbCOKJYuAVzk3L/fFq
YDy8GhsKfPYVM+EJKATJBa2suY0nSR4VUy0ZgXBX8uY0Eu0rc5F9cUP+ZE86+Wy6
wZVRkjw94qQagfInYtv/4WR5/n8l5/f8gCkc8cc3Q4gUUzN1oiPNn9hguU2uEOJv
BL1sA0vzjHFmQZ1x6pTFYn8+DHrkakdln+TtgVVmV7uubS9QUwp2fU/S4KjnOY2t
gTqcPgUJn6+sZ82xH/+FMp6V1heVphOg7/YZWnTrP+McsEqLFeDVdba60sRWB1Pr
aZSiidf1FbQTZIn4qCINLBSE3YifZHLi5ZAjSA/o0ACA8cGJyGupPa0RUoGMSC6N
1ANgVFSej/6hWlP2PITaLtIl166i9goeqf5M93vwrUkEmjZpUr03lSALwI4Gxhnf
hiyPRGxbq10PQq/CsQmeFreZTdtveccdd1Ln9EwWpNoKNjjne0gUkHyl8rrd1Y6f
p7DY5ZsBnAsusCUGW/jwqb2p1QQSMd1QGcOTN+B3rr38zghPinjHtI2ipKO7edKj
i1ODKOKkWNKFgqzyyBTwR1T5v/6l8fupMF31DZiKNyTg/AAX6/wDIsaERys8rdt2
81nhrToihLuRELERfHEMCVxdemkCfdf1Ke+VxG50nNwRlTK0eI1sjadU2Bs2ftie
s8eCPPW4fDwaOU40hpUGEFrC4/kQsRDN3vmwqmQ+1EyWLEBW8F7K7K5D81DD7HfS
cijCU0HSj69pv/bjU9Lp+YeqGc7s1ORhfQUIxxn8kS46+T3rPTs61JSWW2KDNgKA
qIp4CoPF8RP2+aAg+5IZMTlXwILQraDmrCETpg1U7J7LiRB0JGKsxmAEVkJqHpJv
A9RboqmN6AiW5BtVqrUWNRCgcQxF71S+oHbsQfxkrHisE2fZW9TZrZMNNbe3eNLM
PQf4u0+/bX2yrGnHjuHSO6PqcPoiFwvtjjJlZERBxdU6OrazN1JSb1YpZwm1o1Pi
Mk2ZbZJFbJH9kujjzUuhEFPHbqrreYdJ6MAilPaO98sqbPvlBDfdIhqzV+Acn+v/
hfB5RqAvIwsqYDjcXNTizqJ2/0YYg69cE77pMEu6S0H/LQER6MaePUERtQm50xku
fRpeqXrgWiLU0ycQJqqrDRFITz2gHbmvM6BDxHFkvvW0XWxMt5j0K0TssIjK8MEe
ftc9WhP4NM3khzjTAqnOb8wcx7HfbafYSDu/OXD7F+N80Zr7QO8CYyFFAEdLdOa1
kX7nZ9JIfOSObbVFZ7r19i/aOEgVZ0GO6kvL6LMkdBIFAi1Kyq9J6AwNghqsSqM3
mJinpp0DL5RwDL4dlLXPrLgqY5Oq5Da+JMOk9+vSaZxTC0bwhevFygYl4DzrrVY/
6dXMGpmmtttIuWUQWj1RP/isTRtuI+VuZgLZcFOBDIIBU5CHNu9SAAX1JVqbwyLU
4Mt8t55+S4IC0pR6Qktx5yLoxyJNzKfFGcVN9PsCjXX+SdQC5LxHjT+O/XNT65uR
4xPxJdp3A0CEsm/g0sj1KfHfhhr7w80lF7e45BEY5fl38vYdgtvV6PXWF9HGDDIP
pi0qSQf6Bj6UOrrRe5zOspv9UvhLMbWGLq2Eci7ui2KhOsoKlOW44L+kjy7eHY7o
7eyn3y8x98kC6JkxcLztCpRRisANWBwqMdus7DV0euoLM30l8ibcwoZY6JItPvZV
ZHf9bMhVUbzXSsrmMZvwf+BOkono79iMQ1wuEsY7DQHRglGWP6/U+OHFpyrmEffv
2lr5JzU76hrrqFqNYrxjJw6pxNlOeaKex7VI5A9TBzGG/iir50prZFPW29/ynwtE
qLy/ckT3knNacIjXaJwsAbzPK+uPryDmoevVbsjhKay4bMgVdWR72YtgX+nYrgfm
6dA1bMJiIzrJg0N9lY0Q7M4cDJLLfCl+Bf43h5gEiAcEWLmeJR745298gkZeIrGt
784OvWaSimoi1ZH3KVVzXn9jIBhiH2O+BmfOB6OKn0mMew8dNGxKPBN7wC6hFsbK
wsnBIp2oEXch+ZB7Rkayr9OFCRNmH1wx5LqzI/93xs1sfpV2iuyFLY+K6EInVZ3W
lx8SmMOft18bDDKZmvhS22lkQEo/OjmtKF0RaW6ydb5j6OiElgVsRh/sPrrCETyT
gMl5eG42bCTAeM+O5t610P15kBFNaZJrv/ckZ5iKFP/VLGSitx24Gpm2Nd4te1Ci
BFXbdlGjJNV7Mf5FyLORMdWH9LxEDYfFzkkTU3wylLnWCTCaldaVyu3vlrGnWd9r
/0erjHNqSwH5VjmkEF15zBQO8FkAW/xG9FoNwMA81r3q7m1CSzObsD3rzaGBQa08
SRzUpe8qSdfgL1yU2v9E1ZV1u2AWONkD9flh5R+Jd0tLg2wByZVAfUo2IgHrv3tg
kuLGtslg9dptkIk3nLYJkcfauYKO+lLIsZt4iSpZYI01lnqlnA43C78k6T3NVgw8
T+j+/2LsdGLTS+zGjXrE6hexwTGGlk0Ql3oZ0q7597HPWTNmhGBLIpQFkL0YVUUC
W/Q21dx2WBY4uOhfjQf3k4Go1jwm1ir8mWq/Dmkr5OyJToIXNrAp2MRKUJZSC35z
g9RLxg6T3I8VFmjoeW1HCpaFOn+Sn67RD6hRcdW7V1YeSUshg0BItOZLe+1ynMwq
SdU1ZNVP405OTDDHbsM7CeTEpeuK8QukRFRUBKIYmqOCp1PI/qwrPrPotbmKN3Hk
QmUW4hSVXt5bAX1wRRqhbnxIjChR4uVO9O6rJISFLA1F/DGmoBQq/OEHTfIrleCR
XY6dLsUp+SYQ7DVJ6Mfh7AXivqJ72MXzj9UpiBbA0VQkNSqYe3d7AEuc3+ATSMNA
mpWQuCWbkDryZXY9trEup06YYe6Cywzv92ECwgAEvsqYSisWz1crkylOqGfMNLmQ
1wq1n1IkGnZ9dZxOiAlB/fxX0OteF6yKtsSIDgvSJt4/UMs1uG1GLdNdrCZXEbvO
2wRyXwyBwHrb8KKKbnjtg2R37J0N04YxSF/jdxJ41+skH4QdaOBYk92T+oo3dl7D
kLefoQzmbVHnPmFPJcDN8IlLfnv6H5kyfSGcYokFL1df9CCKWpFXfb00eANSGFBQ
Pse5NVXiVkHGC4I2CsFuvcQoGuhtWNIc2SYQ6A4+KZa4H/17DkbmV4IRmx/cxoYE
brbaQS+E7sdYe0FDuwIZBszWkOBPenqp6nSDqRDWhZyV6hBgfqiSlOpCFAhDTEyW
cEqX/eMg/GwZKrG3XZrhrZ8BhEupWlt02f0Yvvg83QFCgAYwx0YeRZY8OmpWoVgb
PGJezd6vU1SOx+taJKyKj8/Cx80uoNvbNf6dC4LkGUu7ioq09LZbsOkJTTP+yJnR
vcp/GN186C6QbXKHV7wOcY/E3C9HCuL1ToXj8j9CkzJOg16D98rMwvEG9gi7g7YE
u9MTwXD12C/JfUSvKZ0Rpwq3hATkJrTqw4y5BppesQ26YUhUiufeEPMD3scSWzJF
48UBB0NqgIgR9yqen7PRn9/XJlLJwnafnp7z+M26lDd76ZcaPnTSiEik0LVGtAju
IUiScfKYZVoPD6XcBVOsCaJ0NPyeilvU/eiQ76BUqgUaCTgc7/g1tP5IxNJIAdVG
4CEwl/XxV0z2N8KmrN9X8CnzHz4kO2TofDgc2Gciy4X2nEsrWXrdux6nBr1kP9nJ
+L5BERiemESh3PZDNW8QViyTPkgqp42TRTyNHEkgSu7St+8amoBFxQ9xvMlYoyK7
00y8tC+DbEIhaZpNQ1tCX2Tlz9/n5+YKzbAx5sRTaW1c5N2qF7C2IlzptEhQY4z0
6WHbGk4TJQgNJn8qhCBC+ff0hkEaEzzJbiZigGQ9bWto7dQJECbbtAF6fNAeBjPK
TxmaJK0oKKh1oyj476xjeOnu2Hl9aitPHTRplNvJAMHE5AYqUxDp8mrINOjDyDH4
h6jS6VlrJplM5A6mxGBnf/wWdMMn/EPxg/a6yBXzEAI+q8yLff5TZY/AwUT6CrsC
tmdCPXQLNj4Q8s3mVICsSHD0vmC+pWHTz3m1KRRiuOCLNGu5/s2G+P9FaHiZQawq
9FVhhgi6HFuJSPktByny4nbhRWzcvQj5CVbmlNBE77VRYUXXShsz5ebjQFkgKpoF
UDFOMY+KkQ9vVaLVQYEP2wfEXK17Dlu6li9xt0bFMfL1EDccdx+clcuEulo9JiG3
mS8L5z3Y5pgnWGB3vui1PB89jSgdu/PoQkrG58UJmZJBPQXzxpC0rpTjGi0NeK65
9v2uCGW6GFw24LHxyYosqKGCL/YLTyHZ1mNtTojYPN6W1tEtdzdkFkjeljmt9aJs
R9whoFuD5qbuPasmnNRGVH5oiFHfjk2vrv4aMXtvks6wQLay36zzef8wwcbbRx1q
YvwOR4XJ80AQc4iScOcev2kiAbkcU/TAaPQCB76kQvOC96c+UMAJdRvYYnVuj0cA
JA619opFygpFSUTgqYtm0b9DKNVvvnjvcq9WLzM2jqQilIC3tAk3MbidcAEJeCR0
weytBf4QzD9eG1aDN34e9DAtm6oJYnXnfTkmf08juxCVDogHUs14/suVednWGdqD
lM7xBcbQXlGLPrxCKBSDNSKFhuLycA18yRaARkJCCnpvep0DJahcEG5rUhR/cQ7T
sH0SDcGdpXvyQklBuMYMm8wQy/g4J0pfb3EKOths0PJ7G1TdtsI+mzpgtBYulgaZ
GfRq92AFs81J71VV+WvgxKWdc7bH2eFxSFVtjhN+7D1f/iNQ+18XAuappogAnAk6
a6YxdIdWejn8VVU8i/VLN7FZzK8042jGMKXndIqPSmpDQ5vuZCkWzfYXDi4LZ5Z+
v+2lUmwTOGT0RE31UOy0PhxRp8dUlEAVt6AD4sI99MRbcSHT8e476i6Pv9Bsf3/F
yLuL/AIDN/LUwqQn40D6eOaJTTPnMx7mk9dmrcdK24XBpPDnyS+sWI2QF0KDm6rG
Kr2N1ITLJZ5CUytcEwJeEQ/HTfDocAHOh5PFSYOGIRzcLiNnO/89XDgFcF1wASTa
zTHSJ5n3CIq5RUHLbTbMfJ5cXgyYYtG4Ntt9smY+sGimPm/CXhIh6yfZWOcWn/Ys
RKD52HTDeDyjcoXAizlKJLdnXUjZABYnK2EGhV42JLq4NnKaoCeRRR9TWJaFYJIu
Kf+oM3AiAw+WRWgvrYos0l/7/ViCDShci9YF3lzFzfASWxdPEuwD998R0cHVGs2e
/6tp02eqDM7aE5J6aVx0dwRmi4RyETCcoYkUUbBh+gaf6s3PpqegMliwX6WwIRjK
Po/Phe+ZoVxEK0X0IwPXKfnVMnqzX74Sk05gFZWQiI4LaX3RChFk+TXjhFFyLqcJ
JqvzgxQXJBCbO29ibfvtnwxV72s6bYDB+69Zjxpc5ch4NpBzZzwxRF+MLz9vK+S6
BhdobsyeSPP2WvJgU377m6XJDIeOxZjNHJGBBQ3tVn9SmG9LlbdxyQ7ZgjWQ++Iw
cHOs2n+obBkuLrpFNzNi8WRRE6wKvvuQN3Orwj59YuEec5nc6ytjjNp8iWElAixT
c74bYvfRYCXzGJe0yWZsGTIWhkDWpJTE4UvPD5lkIHleDay57KV9nsw0uZcaohu8
Yq/5eVCBGZ8mtleYfezrblZ5pgP/VLUsG2yrJCdwYMwh/CO3TkR0CjDU6mYejZUR
bwjc1Zot34juJy84EZRBYG8BZFO3CtqWZ3rGRDRfTxUtZS2yRIEqMaqHI7g8aL69
JlR4gfYMrV3zeFld1vAUkP489dqQK1Vfe9oaOEscVovAQeieTfYK7Cxn7wdm0uk2
LYumh08Pybz+xEuU14qJHcW6HzmQGsSKVyhXaQ33DSj4upmVIYv0+0e9V3ynl0K/
qrtzb3o5Kn30/xB79l/7cOdz/Dl08wjbwdzyS1z6hdj0NWS9tBhmUTh0hEtpP7sx
eKVc90lx1rnBRJWXO+fqGm3YPUiLwlvVU9dTFq3ibNjoh6DA7zLcmxS6GfJEmBsJ
MNSixmC4ItNDMGqcNXCRmIZZGHy7AYvtU+3vLJvQZKa6jce8gLok289VV+U15G4V
V8VsItmq2d4nxfdfgkCNWAETpU8YKAAdgRRmksb+VrUtVOxonKsLFg6bJgwVLxo9
FOyuR413jZC85D9LLZtmirK+M3pQt4wwh/3pyPHUlMXGcVyJf+ZWmd4ea9USj5ly
l2p0nZcnGnnUZu5fWikRr1COcJUTGKmWCrNFoEZOpB8wE/2ZpYIgmzt42cmXkRnW
Uv7LopBl6YB1oGGa0R18ak3UN4waEjK+EnfIZU8mdwQpxy2L9AS1OGN40rIB9ZbT
jbYtE6/86xaaC2CIGN2Yvt1n1hVQWFxjt1ssyONiRgRgz6gAu63ZGX9yVIVbtGJp
OIQh2spX27h0v1INbi8gLc43+19ikxxuzmP+EhDaSK8VFyyxQNF6zvSRReqtKuBb
jWieGAInT3rFroNbJZ9IUEeWjIWtAO+pzvS56Th6z/KjwY19kzqEIizqQSGieSpG
2Ygng8Nd7pWRdOco9yvX8zHcdwMNdI3DJ/XFdiq8LdkDE4tmFsJCG1M4aRawogna
aCYaqk7229fQFwcYyN3RO4A+QaVz/HjWStYLzx046h5Opi0Y7epTBdPwd8bTKD8+
iEtXOsSRQO0wSaQJxkPy7AofPpW7PeazgAcfhc834YxWq6bR3BtWlwoM/NAmUrCk
twt4QM5kMt/zVRuhwxzKg2KYDRnzuC11pCOCtbzn6MHNCEuysBFRrOCjkv/z6SkX
RYnNOdwlQ/2UOowB+fAMbxZDGiXNzTc65ooH0TDNyum7CT6IyYpeuJYvjys+/OPf
r5EUTOJlk4c7mjQaUUR5zLcj9yi/vD6KYhX61d6tg87xbgpmsAnPjY8N2hglRIG9
fbhzjzTrqyTiPOIWYpTumMUA14VzyEaVtteOQKj+oJ55gxQO+GZtCj/exRKW2+xm
++jCBaHzF96gNJPrCpPZfdnYYDZCRDBrmhb79WKm7P1A7iwjjtnK12q+BdJAPrH0
reol14GNK1hCTUjuMWeZ2tnASIOnX5NoXOwjIQw4Mpo4Vfh3DaGkzL97yF7XEOBn
m3bWlhzZ7gjCRCUzFXnlFonKnzL81HKRj0Wxj1sTUmM0yJwVVS/y5IR9Ak71f+LY
byUxhmILvmeGGfWHAZ6f7c5pPEz1GHKusyYFY+NyqhJLMwqLEdAqAo7yjMgW6Enl
KDMO1FybID02Y0J8ikNvOqJuiag5/iFS5ypPb8dVFfGTX2ckOuvmzFFhWBpCK2j+
YlEkfbR8+tX0peaexusA26s/6pnCbSqMPzan8zAH1Ucbk7qZ22HVK8IP9Y6T9BD3
AkYAXpzfY9dHQ/L2J/+wNBHLptSUGxgGv5j3lpi2Dt5lMmlr5caSdRFZNP1EsV2S
WDDy0BEbLKhAPbio5sgxMLiC0Q9mBwxJrhy3zVbBRncYGj5lG82UVJ3VoZgx+lSb
Jx7s6ZKcvJDOoaqMCGSxdNlAvvHtgLcA8QZ9YY97y/WrG/9gcQyEIPSp8VjE+Fwi
Pd0gu8TrxMZL172pJN2Jta+AenxOXUtA1teW0nCr4B+XeGm491lAClqw9Jhi1F4R
IdUSh+uFM+Iq+DNVb8qDPfNER9gnYEDYZ2CaRbpZoEbcQ3RWVwlJoyZUGyUBHGt+
ND/eqpsDcoYpIVvgVP29biIhQ2G398EVrP3TJy9EMm+fs1ev1kRJrrGLdoBxJ4Uy
oL2yEc8h3G3pHrCzKTFYXt/nYKuAUg2Du6voFCwIUlm16jIcL9FCQgjryqILbEED
R7BybnY0LkbjRxCZDgHENUpwuQyHKOQZZDcvWQqk5HyVDcyYcRbgSP6oJ9Myt3Kw
+983TDse5vGPDlxCvtpi7KvctZHMU62DbC82OtQpThHA1zRgeqRfov2MywhnaIzL
lVqUKLxh3iOFAZ77JuRnsC7BFr5cbVI2hxOPmeWBkwpfwpxmqENc07rN/dFrzbil
zY6QqTKbSsyi+FlTpz2kLSlTbkOSSF3+lOYPuzXghr9H6jO2ZwRhidBGoq6d8X7J
8u1uT/0+ivtl10CqYDJZC04P/bYfFu9tZXdU+TGUkIo6zfuG0nE7iqfVPXaDUhzE
aA5ob5skqZAyiDvqry8FrDBdFcfGnI00sHLgRX/RuYSYF6+1zIo8fI1lsYjbeEDE
9cQcX/5ctDIl12Jwttqptw7+GP1Afe2iECZicAsqtP/FUKfh7M1C9NPklgLmLtSH
J5hL4wsDkvv5sS2jrmlxn9oaIgkPY9/eBSl5d4eJOXjvIAK9V2bWpDH6En+4SNuG
qMk5ZODRGQCc1xO/OxThPLzDAlVBkFDLpShwU6Td3XONBRDMvzYVIjsxi5LW421E
3S5mahjMqEwvbYT29OOJ1UJ8gO04ZIX1DAkkgJZ5jHYj2g90df9zcuJBK/cFs0sB
I74AiaTccjENHYPnVZt+49UPFgf+1DUGJ58VEmiyeqnyqbxVjX469yhAoCCr51W/
iqUoIkrkPz0pHNByaIje2fpL6An0H6dAWN9NhPjHxpJscj4lfpZmx7FfMUEXGTNu
fP8UY3npzcqCqhHrnzi6YstPnMUNpL1NHbYFGPDN6lYMf8r70tqGQKm0Iv0ANF6Q
jb4yVPamI2DB4l68kiW4RESVU9/YnSQbE8Y+IhxorF82Qk9U0DTKy5ioEpggnH00
fwb87m7chl8TgqD9+XB6yWZon2WU88U9LZrd+E3RbB4GS9JUCDmovsp9/8uRB/gv
g7+oOPnveksmMTNQlOSaaE7jr3icciIxD05s7KjjpGjYwO3/us0nSKiNSgBilKAV
BvuiR2pHAz10qCSg170rvhiKEvWK9y3DZX3hSoKt18u9SkOXzG/noeusa7J/+/Jn
IHwLxMVeFT/4VI6Sk072JT0sudxjiqtnf0ZS5KhN5VVsvxlI4ed7c4anwV/AULnh
xzPkH5/cZkVZv4PVwo8V6r6d8zjS8wv3bDzvfeZXQ49USHmir/a4QSlzmVCC//k8
s/nApwz8puHq5chh4o829fpTPTe0mIbi1GnstUhiXLGiQS8MTKg4hmgGvEtzFy5q
BUoFiyeXz6avzeu3dSDlgr0m0xV/5lxw4gq41iVR6SO/eDyUjmeYlJcHKjvydLDs
6TtFNkHJUBc9rBnY2gl0nNnh/soo1rDWAKeT4Qd3cTpQ/d6axeq6w5ymzL6mXQ61
P2h1pt9Euobbfmr4jomR+bP0YBRmkPl2pVq2D3ZtPqrUYwGsYxGgZdVlVtjZsB8v
0z0Zf9gADImoryINVBSp69HtnTzpjGQubMmJ9elMHlE4YzC671EWw5d0IWrcLtNR
+7oTPHYUvqXpuALDmG9eFiFpzb/mam7jyeGYF/OUrwA3JV6rzOEYgXNQmbaWqPMw
Ze3zAuejaXmpiv7ZOHjOFJBhLasUQMWvoQiDlPum+bE+e/rebSDgxEDUYFmpXEeU
`pragma protect end_protected
