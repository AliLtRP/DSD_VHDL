// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
ESLT6IdX99AsMGRDII4deMxcutRRbyE8aAbza2bLyz+F8fv7mDXqi/SDddQTX85/DGPUO920sFNm
hCKq/iv/NpPoaGEp9DWZXDVY4Vz6XYu4/UQEtLMbzrdBhkyM87Usst0F7zCeY9pobgT7GCMPLNHA
+hcLLXixLeNbqdReJ9iW21JxkqDAsOMQo1M8hovXOy1btavFupn4VT/dZ81rV94/DAf4wGumAe/m
ux0oI4rUvBmlKkb26qvlUaRQlVurug448R2LyrP0jYRWtLCaAoonChr564nidB8CRwMVhRH+XthW
TnFP+417q9LDq1dTSaGQJrtd5241YSNRbBKsVw==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
WO43CyB946mx+HixbFUuqGdFDnSBtyB1YhAB6Y60KCa70cSskSUM62BNkCiIIvx4EeafyVcnh8Ie
KnXXvfp5TGe6nWmSk8Y3iV3tnqN04nGp3CvchY0aQbjTgyOmo3KZ5CEz2JgUQAkw/YlqrqmOO+yz
+q88HftDL2T6AFlzeP1ozmc/jPOfS+eug/YCFHvgHShTd6yBRjZi+Zio8hWxszB1NuRN0fwpB4vt
FP7xWjx7oTYY0IcEaolLiwgWsZct8V0hz7od7rGsLmLe7umBdvtjD31FS/ywiGt1cMPjwEP0jklx
+6lkKWvc/uT1Hj+/uwNA0ni6InfkgITITavw5vzbfMbVJCdBFNNnulqGzBqNM43Ri0z3zoWDUtEH
7s0zWw9xG2g7ZORd4ZabmMxyaJ1329an/dVGqNYF81V5swz/dHwNHnpYzaKDsvjJb4cNyqJawFRh
FsUj3zsm/kn18KzKX8RwKwlb3PQ33l1iuG0VxtMcsar/bw43KmIcBTynx3cbsNDo8WonVA7UduiI
W8LH5haICvFisnx+MxnqV3EjBC/G/qk4IJfouAzVsu7r/Ok+tyvLppVECLYVu9BTYwcuUGfXqv/Z
JOXky/OEJ2eVHS5X37E/q09BFhN+SSR+YBe9knTOL8lR4XfM9mUPZaNtjSJpwpD3QbLRn/v3ukZV
1NqyJyp5odRuHL/jGV50mnb4UZzC+OHslR1y+bXiap0I0v9dmKZI0dxUi3TFpsZRGi9TLUan7NED
E+wiA6iyfEOIQN8TR/XO0upuWfJcjOCKshnknuPxzhlOBlX9scYntSq9ixuRcRENtY9CvwmCqGiC
B0WlnGXJRDG4/icwxd+Iawp4pQ4bvjBptDTiKZGYnijj59eLFlH2YVACPpnwjIg0+zPWnUvjgohU
H5suLeyeRC4hNUcqQWFR0XOkouNTs69R2cHPhbBC5jBLYliv1scuNFqecLjPYvpbb6OsPMNZZfyq
vZJeWb3xamFkTlBqt3rjGdZNONmUqQ9Nk8DCGpJdwQdYEtmZrMhmiazq48mvcXHW2l4LncgbRGDd
ItaOvJptB4EdmNv5+uLVephm+DFiHUcYOduSnWuBHV01Us0vpBbIRkHWBp1UM02lmD9jh7Gg3Gcd
fQBgblj6Jq7pQfk1pzBFCX+Iuxj4L6H8iMq6e6PXhT7qJEQOYazUhM+3g538AAmT0/YCHWw89Epl
xHH+bJldP+Ui+EY8U3QUYwFaCiqJSlIWxKK6sbvmZA6S5O2rAVw0dT4zjALLjDTgsFsiUg0AlkXf
su7dxfccN+M4p5ERESLvakM9ZcLmOkPkqbmPA5ciNXdJueVPPyFZ3je66IO2a/wsJPHfGphPD8XS
+XpgDHK0/2Z70LuQBox8F5DXYdspWnzd3hjxYt/lswzNUI3VWWOYPjAtiKNg/HeVxxICct90jzhz
Y8JJLFN55KL7Wg+ymYAVnQwFIT72Ll+WBS4Km/ZKzjuMYA0YzuwIfSZclXqT7gaY1ijF8CBy9rEa
RyEup0TpUSp6b3HQeLLm5+1yPNQbENWqD2kNCC18RDrzJ9ryMQ4F0wVooKh6PyvU/8l76IRPihLm
cqkti5wNXYHQPTZ92LrkFBJchaGTj4P/WF9SB0iU7oUXwGsKiTx8EHr4MrQGBwb91lO9fAaS35kz
859FKBVdqkaTDjnoPEZiyAYEOcvY5s/Pwe1VzHz+r5rH5QXpE0WtvQhrPX8lM8Dv14WmaGbcZHEa
J7l/3skmrKUjIxZlOxa62G/LxjModWC+856X3J4yci3FtXsTnTUgujIL26OeUjqJRzTmM+BtEcLN
JAZoumuSeJtLkineCtijZS3qui/3VCRasCCHBB+vtjdSCKFGnnHHkwumTLECYWTpwxAolZm5YpwD
J0/OWJGkcuwXQv2wsQfpYpXMaJ9PmJ2eMVGvi1EzRAv931eaEKQQM2yjKreblefYIpGB+aIzE4wn
cFkzA8wKEWQOH65kX0C3B1ruN6Y7UsTTYiNzuaFVptoSBdvY6Ba2Pe6YjkJ/uFZZ7/ssEcjMfcN9
VanF+NnQOSsmtuKCisnAxIh1n5J/8RukdH0i0xGo9VmtGcGXDJiCi6z0s9EkwZ7N41X30umqYq03
lee2CMZpqZT/JECKHoBEpAGZS4DZP3MhmYwD/UlUu+TIzfP3Ln7EKQGKJECQobWrVs6MUtGrBmLu
8hzHAENuy1fGc2LYCYYpEMq8rLQT4JHUhbKjErdDOhdJFaY99KMfPnnt484E9M7fGxzifIqHL58n
2+YAc42Q8KU9qd1eNKhm2ACPB0kJrmSLp0iCafQfe1L9IgErPIPKMvxNLe53qmaazPMjpcu5UwdN
+ziZ+/W5uYFM9xkp0vT08W1AlMpWuYqCHclNPZsdgGcscKuvfINy9AIxizeEPYYVorkJMJTCxabJ
ewzXNmcls1MBe0m1wPjKypKBmVfprjlO2f2lDWBAWpSSxJuoG0QcFLSnI5cb0lib38hu3yIVeQFW
Zf/K4yR75vTpk4uw/5QLoMYYspmW7RMRYBrVnKWDTROQdMU+BOiM8KFj+KXfgHFMW/FFJoF2wIya
6kqABmm76vJLED4HguZUCDg3R9hdXCVQpm3O43WitjpKRF517s6IrJQQRiA3jSkWxVKcrravbM46
ookh4QcvmiHLHV8MS5RWumrSH+97r51xHPe5eUjm9sBWlL+6AU64SZlZoeZ9w4tcQnm9qlPTf2O1
k9zk3e30O/eUdJxAgo9xc6aouIapFt57aF3KsvQAz0cl+RDkuH3c0JW8SkbMalQwItsoEbj2PWoZ
b9COj/f8BjACyGw54bZhQJT9K8AQnFq3vp1KJPyg315jRPkx7mxsQVcnc9lV1a9cGRQslWL4keUG
UUry+7cmNASI96Hr63a0lfofHjrMpx6Ppjna2O3YRytdfs/zGP81eUTFQ8nwB2B7iKjSmIiOoK0/
s4meA4zxJawkeZLaSAij/Vx7gcZIbtCcj3wYEf046E5JvEFUWGmF7YymNysqF1fn1LDRo6QqGcYM
W7ZcGpFxSdzCL03buE11Kbm1VfvHiObeaTA/YpVzqssxAxTDLMTowcobFvbVo6RuZCUOCqZJcmmM
qdvorHENO86yKVg4eKKvZ/Q63jjdFOfJYpetqUEsytffK+yFUnyoKlYinduANkVYVJXFV6dDjPbF
WwZAyovabvR1SOs2yE8oQTpEnRqtk72Mwm5d5jhMNa1HbzJwpe4Gd4AdM865zU7UeL970VeeowMF
8GmKlOr88INk8V7EgDboKDEBc62ZMWRHhnv6c7ABz0iWyNHdF65bFBOdKaYgcXXmC5eiao1QNoNj
Qsq/rtOONw8bZ1X2tnE10OmzHEKFuSGuD9NTcXdm5hU4u2hGIzl49FK5+umv7Cz54UyYhSDcRV47
zuqGz51kJDJMtFg3Z+9S/B76Snrx/a/P8Mmq5hN4i6e6cfsSgZfmhskoQHAPV2ZJov5ZRVTgvWoc
J9lAvbYbyiuOtBswbCBC4rih2KJ3dp+WbVmwElETTMS8j5GNuasJ6Q1qwDPQdRsYlEBLVKjIaeJT
NgGKoICshMPfDQzJlyl8tDS+WDVG3+exrcirbXID7ScE52qakJk3y+Sz5D0N/2LuA08LtfwHiOwg
KKv9a7L5q0UfZuyR2S1f5+0Yb6iAMtoS64A2MUfcGcbnjczZnHy3Q/JQ2Zf/YWJDu7JHhQSL6NLQ
GvykHCQWpxR/Rax+WjMewjUcJLxbN61458Dt5rED1PH8GxO1O6kHxzLOB/njMWNdkm9SqcBaSwlN
mVr1/gTOtOGwQoqMr8yYtSdzIQPiOzmYs3ILjYSAc2uOd8jcacOjDZ+CXZui2r/4sFmer28FFwyG
8N0a3Z6TMvTjgREeauoWZwbautsAJLiiqcQbhITn2eftWNMtRlJosUI/Qg1UtrV655glYq+BU3PE
wF6rJAYNvAANW4GyW0dv31ca2l4tlAJ76vl9D+rDF9hW9sxC41ZitMiBaGEBJeKRjeiL5s0UVRcj
Oal8sgvkDYkB/9lcWMNOmfeVa1i3yv3hcYLUv4jMFIkqRlgi7h4K8Qh8gFoJ0jQ5fQel6v9hA7uX
EJZDVj1ZojKSs1hBMU7EBx26DwVBb5uS9N3UVEqvWlsLOKzZ+DyZV0vvw5O0q2NliB7nD0zArnDo
lZ8Y5cAImbh3GTibQraqDTb21y+ibIrVBiH7yS1KT8qkpOmE0DsHJlTgbhJ2d3lzvAT3N+Rghode
J4TYXVX9r5p5n8q/PKomesoQ1sNjbb6bUBZ9qQhsGqv4UxeLgTCcZ+aOgkPZ/Xz4GP6QmH9d+QR+
zW8Q+OhmkP6KIKiot9jDnVOSxrPdTV6kQosyWZE+wiESwyYennxzbeFpTxG1ZdFlIRRY0HjM5xqx
SVo2qSJQdCgbT1QekSl3IQyfdtgk0kRCqea7LtzSsuI2wqbu9m5y0Q4NMf88oFBFc3L02cF9KqrR
b3Egy+XU8G580JZKkF6NFE3YfzdVhCT626ZR3ld+HTC/RHg7FUiqQ/RIps/muOUIa3OTTUmubY4X
nwYxOlsoziClVmj3tdmLiuYToN3wqlgZiTC5MSdCTusLdYb6Mz/BtB5kJs+pEMd3xLkAtaQi8Hj9
+dv/dbKQ5Qw0bshW5ThLTfKsgfHulZETG32R5Lt2VXvF05lrYpXHOlV2SdT+sza+Q6G4eysy5RVk
bbwmdlP3SKQRQrdfXm5HgLS/W9PAM9wwk6tIOpTXEcciPPYo6E9WvQPBIyzw0Nee266+KoV5HzLZ
h27MVrRZBaLw89mAKJ0eMs4V+ynYwB70EZjI8itkXlJpE/MBgm2Lp1PX8LJrYDrgdWmpnwy8umOM
9ifUwPdowHTjCvvFoMsq8NS63zb/Orr3D22TCNvB2wyp6Yn2OA8txQGoNiMR+DEEBP/w1g7+oXhL
GSm+Vlvb3hRm6hkoohotk22lDMaXUCjCx6UESxr0eycSvpv8ZHgVfU93DfhPhXrsFiPde3DjnCnM
P2nks4z6rY4ZT51bPLPaeabcS/V5CxRjiuzfZ5qeOcqM8/clkUr3ickLXzMitcKTRUcCs5lc1E+F
446IzBzNOJQeozNW9zTQpjy+QXjzPTPv4Pk2yKBNeqGjXUK0SKjlWdO1P4TPG7Lk10zpjr+AtcMt
DWmnPOMhqr5HflG+84RJ34iRGCs2YeCq/P6DgQ==
`pragma protect end_protected
