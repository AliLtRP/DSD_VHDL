// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:49 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
pAJ+d3v+/QYbsXof1weXLNIwfT7qxIbgs5f9f0jOpewgLc2oVrrcJmqDicmXU43u
ZnHHnjbW/lxzcXvUybhC/uk8pDQE8Q/eNPefbcraxCZJca3lbWUyy3WdUJiNCeTb
mNqmsVbeTe94/tQ5zl6Qy7TfZP6iThH5dmEs7cx8QAM=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 29024)
heHzhr9kUtSgOMnB6WehX8srTEA96zZEOnO4TiXBf6WI1C/3fJkOgl6gdojBfVdT
1xNJbb/vJsPKM864eDEsEzKoJ1ALoelemvgHM5UnHNNFCijxw4PrVS5vMFyF2R/h
m9+VCeiDfqAau+M+YgtpD2EQTMZryxvMQcp1PL0Ruw2UTyvUMKxI9XuduIk5Exmj
UmOpZSrkfNx217a3ajYvTlfCCRX287fWXqUeLfBanVwGy/WajqkhYfbDmSP6ufoP
Jno3V5BGgswQDRAM+SWy5LrQ5AVloBFa/pim6bdd4YN8Vte5BCPla5Nj4ZadwG7m
FK5IcdfO3a8NMxxCPpa9NCu22RbLvueWYqjj3Br4fbPt7ibIIUl3gCjNUguZ2Dnv
ZO5+gZrYNjDjyfAPnEcxNTYO4J9V4ZXeQlAHkFJYcf4kVAYILOoVecNsHwuPFKyx
awQsoU2gwNFtgR4UYZ0VmljroR9f/k7aXnL/1B6Tl09D36AGHHa6U1A2L63EHfxM
aWEa+swU2b73wQ/JxWAJ2gxXjT90vFLnoY7/nyB5djmI4DygP0dL0tYGU/b8zcX8
U7Oes5stdJdLiyWxSxtICIdeM3mMnuSZ0z+WVKsNNq4dliE6HlrOjZLPcGxdL2n0
LjjmQqp9HK+UmddWLdB//DtfpOVn144zVz8Ij4y0SFy7vQwYPya1+9+5+ZY3MUEh
VpttWoKIz5ij0fSQeQQ+HY5j2YEEQf2hlPbxoRlpxwM3Ng9vSnKfEQjJJ6jU6iYE
5SerYoSrp40/QKVlp9fJp4ErkI+rb7mwGQTSYU88/7qBj1Bb2nYWGXu0uwt8D+cu
n+n+dmvxE8j6xmOXPxyfKhMuf9/CgGVrjdXh8s/8EoJTdl2tEi/dt/Y0tKYjD0we
Rbg5DPemh9opSDna6J2IoID4Ixc0ebg4EIntwsESKVVhDQyjBPuUb8M+nYI1l9Ji
KROtwXNDCrVp4NNGITI6eg+z4MrB5ZsrwcVbjOfpnjVuQ9Xt4sLDRPt/6NcvE6Va
Sk0Ejdxz+iKsfDHqzfCTm+M7vlB/06jDqW/FWCvjKM0sEdm+sdo6XqdrO3RFGNuZ
dNoy/irBhGBefJEefjE3gZjgGENsMDoFNkgJ6cgd6fyICLyT/rFy1WR5y0HVthO9
HVwhPfVbNogi9VlVN8HiWUFIBEaGMWFstJfDj0HaAezbskfkuYCR7LS/pJXDOH+o
8w/pqP0P2Sy/kdv+DgSnhquU0NSyJNB7ekodO+bmB7bXDqExOGbU9O+lpVmW6/W1
lsV39dXl4c21lIr8GV4W2u7L1q/lsnWNhdeXOZUF9DSgDf7eh2pzR1FKXRnic6jR
xzEgfkRayPG7BEbeke8gnmpbeikfygjd+nmvqS8B07JfDIFtRmpwRyrMpI0isMew
dgJperBsuavYRKtLEjRSQLxAAdSeXTzdaAy7fpo4ePYuw6UKI4suJwtSA19d2WLn
YhjQrJsuUC+i8UDA/UpD77FO+NsfqG/MWGq7YLBRx+kpWevU8u4UDS2S5G2gRser
huOGMvyekYmHCGcjOW9DP+u/vh2FpIsP0KrrpSVxnyNulrna9Ni7Orivzsp+aM7m
zK9OGhvCsv1sgboTRcqMYcKjCzv1g6xxGv+q+pr3tTpk5tEom5Jl5mMEhfbM2LZY
E+pOjyD9KCZSIZ/PWtEBtvKQjQ73NZGa7k414tH1yl40Kgi/i/6Z6umUymovzFug
LSRSJ+66Vjt0LA6tXILCBF0t6SG9asPkYC3mweq+pQ8r6rSwKE0as6gmM4fr3DI1
TUHIn37b29+hJjd1X64I9H1Bz5dDnHFByOFvMEXvUS27i11x7BavpYrD68IvPr6Y
bh3eAX+/hmX3qBbszhPpRdb71xT1IiClXxGdaV+1ajiyROTjOJWUsFHL1nTWLmpP
s+sn4IyFlMCjHfHigTXfreKhZREiy+7yN6lDwDQSkhoMuFH+p8oLV7eoUSfz4V5N
sGmYkj+waFGfUeR9pE8jK0tZFe9N6y2sybCiu2S3baoWg94NEZvtAX91YuKqvX/t
+pJecOXKTgol6uuOHhqM6TGOQVNLJBmIhzZ0o5shav+iFnt1NiY5Kt1H6mMCVn/U
KCLWB3okCJMjpulhC5RwxIUBYS6/Qz+bERZvezWWsk5fcPv2mq3wpb70XgrZPnZ/
Ww8t/uVEHB5lKC9nJNwtClfFGM4FCamEFljhq74JV3kzDGQR9dO+GPb74i4Hy39N
MsqBqEHGROXyG2P11+qE+4SEo07hgNN1Gci9l8cSA3usSmFRjaxZyP/GK9fVyLnF
Ss176Ohpks8HYB6isEOJMtCq3ofoR0yTygv+SfDF9GAj3CMvufMNu727pyIBZmjy
pWFQ0IBwwOEsIVYTdbmYWmNFJOGcbeuwoi2IXK0gseVfoqiPek6rZPXv/cX05QXM
KQnoXxoRdRASe7i/KgW29DzAWTBA+jvhCfEuLDHEBQbBNI4BgdVcYFMaBTp7T8Jd
209WEiSE4vE7YZncNwJm7jsHxmylTQrSUMUD7wqZBNVBhriabrhlpp2DOA0W7y9j
MQjcX/ak+7xMPtmskSUPZeGgVDaU5WoKSHpHYqsMPm/rjxGwDkbShMxDiHguasp0
LKVuxzqJQVBPjvcgdzg5g1NbC1RLO45wJDMe2Vp5KBaiVEliDwRCIr/7MBLjY/mM
FrnfplJl0oRpR2IvUzw67GYUCwJt2nuryRS7vUN3iu6c/7xPCVC5RbKMOeNdz1YC
UagucB+R5UujGw4lcW6a4h7VXfV5X46VKdJC5BG8hO7py9PbFoagOXSn+oZtbDaS
P0opnYFIFvhK8g6XzK0m5/WWNQZyCxK3Wrknyirs7iaTw3WUx69f1BvBLlXITkJc
GcN+jNUSnz/rhewqsrR8CPkH8K9+tIJd6Ls8d4I8u9JSA7bPjt0yGrjiNGQeaDBK
1ffB4qC8Klh0RUnwPdosoE6Ac+N0h/P8fFCvJ0sofaD8qhZkeRcSvh0nPp3UIs4l
fwjswMYtId9fV7PSn/CLhmLVDDt538u+pt61sGHvE2qdOQXLZ7wH+xNh2otbYdbc
ujT6T67KyQGHBz2a0sp8z1QOEr0TOeU6SWDA+z0XymcwIMxT+wxu+bWetHeYEJDs
NUdIWGsG+d3hOuuFu9zt2w9tiFgtQUw+G0FNtkZjGlEF7onRc2jJuZVsNPtlCKx8
8Jv1B25WN17DvLzddIJXd+OUxfa5ja2lltNwukxqRaiXksYY6ANFsyVB3nTctrcP
nn/Aj5OjMANYfj51bjB/SB+Gyt+zjFGRiihUOQHrIJJ+ewM1cI/1T3bCu7N59ags
7P8cQlTUthegZHc6OYsVDAyIPDvL7+Zedb1wa+8FjJgYIpY/nCMvN9XJmloQjYoV
iYS+9ghZqSs4qzm3qmJvFuY5b23xIXhsO6qX4DvTopeYiWvcfwRw83XJloe0RYuE
sSAbp4vE78rj/4Iin9IAIVIulNTSuPf7jBYFRnW7h7yJl2N6XgQYajQNtsHw2WO1
2ONL+OMrm5eIakoMqTXxYTWmyWDnUQc/8oFKmysy3ujzkNp6lhFsG+W3X8xdMTrd
LvhDuCQYWlD4cWIgtOqRV2MyV/kCwyvjfB3IzNSBzReUXrpyiXLonEv+O3vYi5bV
Z4Sf0PLzgFWRodFgEb4cZERwHF2j8yDEi3QCOJRyRtuFDtlrC1W5ZatY8swAOD0V
AiSJZa3Cw15EGouN/3niQ5bRjsruy3XNJ7bn2/945tR2ZFE4YYMXj4CwDLVwK0t3
bQPHcAuTWCtuv3bLUe31rj8pnywp+EGSkDjY54sJNYBGyzTadnofxH3eK6EjjHDc
0TW2pgciyGJxgiezVi8bGGPYA65EawC5/9kiI0LIRteuxDN3lzPTEIuL+/kMpjZk
n4Vqhq3OJsAUOOcJ4t1pjcgjUsxatvOqeiqtbFDuP/6MBnf98Co4VFjvpgrwu0mu
OB4GFYgh7gHbYZMRzhyTH0fcrTJt8H48G6vcSBcZSVw5WON0EYaHvqHYC7BVrXPI
cIBbs9vl8eSVk5mryXbFyUVx4gXZjRLjvq2K9maQED85fgTipFMwdbuBCCoS0Zkt
4JUDiNuerLABRthEGTTdPf9upyEltIw2YtG+uSf66BKQ4HsrFulMU1wnVoUnY8Cf
yqXYh2E22VdNM6GbtNxaJTrV8E7aLQD/WHZlujaLJL9RVDqtSQ36yKvM0wIJapXo
jL5sWj+PetIdhj1r5qz50fCMydtRxph5cAC8IDKKifgW26i69i92Y9H3WzfA8GYo
REN2YN70qHju1hfzY37TvNPAS+pM104Y/powvCCODeXC0INKop7GsW04dMQ45Ua0
fYnmhEFKkOLPYj1Lts/IrphYNcIRB+1O9bv2dm+0zB6VvwIA6IeY++cPVu/rXZfq
MJgntUBJghWXjzK5vmnSXggZZJVeSGnmT/yh6h/+ydLMDFV1k6KBFNCT0vg2T8Nl
BwGfWEVeV4E0V+WvZtrFiitXMRHqIGshChZ1I1Mx4CTn9B3vXvPlSloWNvtEY/xC
QRnI8paBS7pmdGoMwd0ES2VMxxgo94ac7DPwzWgqVxXDyMioXFazrndxIld4CJ/m
0m/kpNeZ//hlkyKre3eqZc5eNkbeR3oVKeE2EwqCd/y02UzTj8Zer8OeNA8Iz5dh
LuaUVaALuZKBEPbeqh84Tr95xUifZY/GfLZ9HNmwEbXtB4ZRg9Wy2W30QE+ZYngu
L3MqT6o/b3DgUHkxmYlqqwQ6APULQUqgo3oUK86UvFBWf8/zTQlUR8dyErg7iE93
SyRC+d1U0NO2liDAzQun3+fFazo+1AwoDYzEQEmaiO1x3nuyTvtAP6DZ3S8t4tPX
HH9wlzz7wvnNuJu5lXfZyZZEs6p96yc7ld07O6guliF79dL8fSKlUfmAX9YfTVTG
0i5WqrNE+jNdlXlTgNLDjSrIOsp6/THOJTPjZDKgM5nEBIijhZB/RZzXY90yDjRY
5cTgnlxo5CxXxMudmU4dqAQbeRX8BPcjiO1/sSP7f8Dtx7g7VMo6AP5dsxG/Xl7N
A7+HY8RSCa29urbGbvByh3ptsWJvX1fGeFOS3brwL3nav3SlS/ztxNDNm1sSCuN3
zxS+xoY+Ed5I9ci35GbTROt/tdBiX0XJn8qdDOjqfBEDSKzu0D5LKl/b7lj3B7D0
mm8S3wEvbb7OwKWyd99nVR7LfcNuGU3G1N/RRfQLYyT1dfSr7ObAjdQ36TQeMN6n
n3DBS3iJwNt71bsEWRUa56HX98Df5428g6po998U2Jbbv3wK9EfTY5aNFoVIS+5E
yUHV1RxNtrKRDLFHPr6ciwkjS3+cc7hTnI6FjGZIlPPEYjY8lMKlVBzrekJncB6J
XjLO813hU4uw6R5lIDhwcFs5HUrUKmEXgEeW7PnU8UGQ9Zzidufu2Tdo0/YNS33l
GjRXa8PMxZGqHOc8eCcGWqG0P+4ONYz1V3xF/tT3HBj3IX+LoOGEN3eXApCEU+bU
TJLeWNUJHfMpJV21x4Lx1eTtc3e+DltiDZN2xRfPbb3Hcxl4+acEKArJk42BNhcc
w1QjHzLN5/KmNyE4ksP1gVowU5/qHg2C53/nYfhmiQGsZZ9Nmf+1ccgq0mLZzii9
HRyq9V/amjoGrVzlWgQH/GulTycq+/eul72ugyLfD8itLebzWsWqEk6R1tOls+Ep
EwW3ZyI9baLvG+ES/47LD1sFzSieNb2SXox7Hwll06Hc+ggyo5ZencPu3nTGMY1E
ME0/VUpvnM2ezHPnkYPZ3BzphSSO/rqYVwYyvw73vZIWyebq8b8GTnAR6IxEequT
uYf/JFaTT+dOfUhjzpLh646Iw7qJFwG0JHGODNU3UuVUaXq746C6j4JiStUgx4nV
ddZQOsvqxB4snDFRFn4dhXluVCSulRZzORD3+eLiD3JmZS/C/O7XB6/rnf7pyJKX
BnxBfQ1dKAz4aIwlvWIZRWSgBvXIqVZzlKRW0krRowrDIl1CzR8YJt/yS8zIvtHY
P05YykUee8Ud6Z1eAwo5y3hJ2+eZr8hE9RMPehMnxDFyNqWwc5n+76m3L0rz4XgT
Fxj+1E28I87e8PqsbC6kho3cuaTkyI1hYczZ0XvnLyIPVQEmbYORdAhHes7vgl7v
uW5hRUL7g/859bZNYp1yV8pTHpP/+zPQoUWTE9BlyWWSAPk75gJxJoBRVFf+ejSk
BpvvNP20luejN4jH3hfJCb9iDH/IN417BdxuYO6wv8XAhXNDZmaJgUxaZC+iafi7
U3dTmrN1nDIITgoLYXxNjvXjwNGF8ya/lL1DEls8yIhpFGICmsrOuXqZB1fU2WLN
7LI/v75loWxXLZYZP0KUL2mHw3o0KMVP9EuWYgG0quCm/p3AFIUt3OxDNycBj1m7
1a0qj7MWcpnMt3jTyNd106HE4pm/4IbLu21G5t2/PX49HZIEaF1YL6NWpp+QrrBt
mgy5KziR8TmO9TyyQ7SCKxMtVdltd+XmqreWXRMm674FZxPcldutyYjLVxW1K+FK
gTWro//RfkYt0cbhyDVMup6+D9kKDvaZGuJcLIUJ4c5rH5uyoz+5L/V0fVUzmxRv
nfmQPdd6Cm+a/F4lTQDpN8TR3pfbqjTBev6PG6y6Tieik4PUKRUPfm1avn4gjtV8
yey+zSZFSelecsTzWTaRsrbDgPKNUVQvubmQQl0pZhE8HFSqIQdEcMY8jfbYaQ8y
cso78n/VEr0bzIKFdmySL2pmEV+KfCEps7Tkwnyc7G50CdrQVcdOe5y5S/n4hRyr
BKxLT7QymvXShOmwH5Rnh7JmQ7d8ehboKHQjy1lNTj/9WnbUFxN53uhBQACTQIIt
2Gum38MsKyTMcan/SNHQDMMJ2E0CKYNgYy+LuE9LA0w76OL64JRqtGlNywTt6fto
+rCrFiXVAlmb5uvXB2oj2MsKqS9pFkqfxG1hepPAHCa5Yt7Xdo9pybccCpVXZEYy
SN8fhEBOCXu5mHZIKCQcXxadffUXSFe6p36Br5zn6RBbl8cYzF8w2tLdRJ56htKf
eK8l+cEhnTuXs1UNZiw5smURuEJDr+XQt2XhYsE1CrY9CHM2DzszB3ghRjHp7xZQ
2DExvoRPYXubakBU+4jHlkCOtXEUjx95wZuW/ke3e7AgT6QiNbNWFQo1PPsiEe78
yfdNXfH8XTp4HHYYa6IMPE+8/NuNHl7LTtADG6im9QjPrS34h2T8xyVwW+UDSJFd
sv/8/U9Ag/Hqoe7fDQ5jqiCVfMaLl5cY6sqlwCo70rQUZGqtJBBDzj93Uqy2IAk0
rNb6YYVyPDMVi6pEfCnacqTRvbVkIVNAxeul4EXE4zVuO1Ru1vkCs0sRkRMYMhCc
SyW+pypHK33A8I3uOBAjJHbxtrOHFZy1SIeaFcv0DevImD6PprF75V1QeViVTLxG
1U/6yMRlLvJuOvrr6LOUtg7Kbcvu5HEmUNeAufXZXK1gSsEOYwfzrg2NVLHFHGY+
vebTjURKC8tZiaBquXQWnoiuVkI6q5ByaZfRzomY65MnWBnlrAvVaHMpUu6wcXV1
we72GeFpBgPNDlG7ytSEbyEW4l/Zu8I9Al0dtqZGGKJxQ5h8gCJbbMuFlgSIl4n2
GEqwwkEcADtp7oWuabDa6FfCYJWoz2vhsg7739GZLim63/8ooWdN2fZccgtJr3UB
AOCFP6e1yG7300ttlrIPD7D43mefLuragxH95/JwxCOou8PUmz+ZJJ48yyAWfu6d
g8A2tKCPeg8SUPa3CjhZ5hHaIumMZ2Mg04lzv0J//ssO7wZVZtSyLFkfCaxTdB/W
Y5U+rzwKMgYA6VSKhlP50ld00VLSiEFfWloAl8Mre4riRIoSnEY7h/0tBWpru/WL
oFX0KXxLgE6NC67A7rIPyN8XUdGHL2CwHBLYq1LPcW0ZTemDfvoXNjJQcQ+terDZ
TOQ30kbsg/61z/7B5qeW9hj+AOSfcA+e/eEsso3oiXcQzGFxgQHD+J7QV4L54zuh
Vu+jmbl67C4k65nG+s84zZBCXfbfQXfTXMNahA4hznOpHieAJcL2k1La5iHIpNbJ
UWBDGe5o8AKnaqPsVwnJORDnegJ+R+1lzCgwjNy9fFE8zPFqpur0BIVWpRUW+euX
xB5NITydhvwiLfwtdMRDecHKq24b4M4Nm+cy36aO/dEeuhlemukZN6H9gjHT+qje
lTiNGScGSxWe2/BXO39NfmmWezVwa0yea6rKgu9jgFAo2D5d3hhq3Rgab0PWAbKj
f63GL6uaKfexd2SPCdnrr2Msm8kMUr7AYf9XdiW/dU1FRc/CBGIU0WnvkmAMAyWs
OVADJKkpNNhBXwCJFsHln4pVBIKLVLBEvqU37t/5Ua3oL7tdqp2qV3z3i/ZP4U2a
hrPGYmCb5iQR6QsYc21OQtN643U3dyaRfRd47DtNgR8GORx/00CdcINBzN0xwXI0
FF682nasKGWPBNmaklnMxuaDKxkScsmRQlO53QfDiQBvAhbUKbfzPkB4frk84GE0
LgUfz1zC1q1kP1ezoWgqwL87Iu4AGww06r59+mT4p2n2Bv8fefHuWpLJvP3eUsn4
KWYbzxrtMotT8d/s0Zl9w5a2YuqdNzTRgoY3adzFbbmSxudKXj1U4T1tQewKvbQm
yAz1RW2QMICsdN2NyCuZVzZQyKU0tZ1/kHYB+NtAQ64vfhaQRzhB8XFK/nZhsbD2
wkszSPVT75t9Lve1axmtGpXEafpxaWLlM+8z+GxhCbGwzpZ9snVEGedlhpE1DQaP
aazY/XEM7UJNdoVPIiJ8olKpOvDkNcigtUn/3bJdKyS66Ccx4xYC8gGV05hX+HDE
QNjWGZrMKS9/Iz+cNggOfoTQYKoSSfyqf33OcqwRzhharx1BM0E8KyGmQoeMfk/m
/7DcNut3HHcvz+yHxMYhD+IH4O5OZGzwG441MDL8ZvEV/18/hYxu3LDuf1k2G9r1
pScK9Tz2WGSVmmjByvHZ/xLczZ/H4bkQlr/1NVGGOXEyQi1uubud6+2G0hssg/Tq
6JwHXNb2XjpsXvn873Rh+uv3DhDNNxmLAAY4xqJfvqaajahUfsfm621FR28fMuRb
eMm8vBNRGCfqiZt0/nDIWgkPLCCrZW/376MlHP56eGGGIqEY2Vxb2RAoVGg9Expa
6+hnutigFueO1/DV+qVSiON299UDpmTvaQe8n+4OSv1O4aNilyg1dX1KPwiRsG1O
0ct/76HL3j5X4mfUVzrP4v0ZXeZWV6ZaK5zkx0uW313Dk+3AmMU9kRJbFx++AWiE
+NGaM3OrBT1J6+dvwAi83tc7Ks1eaM28QhS5ZZTOdRvFGHIRr93GJIyL/bwvvDWF
3iIX7tazkRups1JDP4pRiBxQCv4ZghGcX8MY0cNhZov67BKjogdurOiZC0aLkWW1
DG/6sM1ZQAx+NfmBeHfX0veybRGxB4G5Gj2AnZzKl0OWR4XkQT5/48d7vOIlisPi
ddECJHqP5WAUGTGNgKoHxDT3YvPx0OEtqvDb3TCVKqItEWIPGdoxRTmPE3yolFqV
JOUz5BPXMri9XhvKl0pJNbDNw5q7CiEJP3C+hM59brWTc8xaEPwphA/VthO085IG
ViuyvJ5wmAhImkUSLpA7xmQKdmGQduDZ6n2Ey/d93BnM/iH/cyBkcYIOPd86nHw3
QhYoN5HO7tBgJcC9H6BMfdybxknqyr0yySKWQPqYE63k6a1H86suIP6F749BtrXG
e40BAKtqFMxzmrx5DcMq28AKLuNWM9RUlbPYWmLApu8oLTn+CjeDPFN/RQaqcUqz
SGFLBUmBUZtXpLtW8tI3ZRUhH7fL06pWjw6niaR0hBn53x+iPtunuuX2ZhHXXz3f
DHLWGsI/vdH90j9hyi1Uq6R4V78i0DKWvtxHfDVmlWmg1O7GA1iXS0+XimsiB0Rw
0LFb36W+iK1PDY5UCpnUhrMYC1HmCGuxbcDWD/VnV37kZtXb+x8f/hCn+4qCn+/m
68sq7VK2yrg7984+zgupMPcezZ19bL3Zgvg28msuUcgJrC4VwyBPCsQmrwNJD7uh
XWZIXP8PLKBR8zGmnP4zYIW4aDduW4weg8aG8EbCBl+iZw6HAAh6vEZeg5Fitt6b
pAAL4jrKSL/BD/DDINtmYzyqXqvnTuPD3ZD0jIpKSYuB2k4XH8McXSWXBSK86E5K
SMAE59/3RiFcHhHF70PpWpriSjGCndmkBbjcN9vBYhO2MkwgId0A+7fl9JOW4/Tw
FBy/X3Krms6+utBqyFr++W/EEqsKYabOOHTtnnHGH4fT6TcWg2WivMYjYvmivQmb
ZwpQXZGI6jeD+gIsgil930NKbuz3wuO0S3gO2iEFk3x83h9GdnRppcumbJmWHBzC
VIXtoM1bPTBAVa74Kwr7V958vab0izJoRxuk3FlImbejs+90sPbmpe9AMVBSH7A7
Si9vMpPhAIUvbZfP/4xOnwVXC7/3qH4qO4x4UAHtz5rjTMLsC79Z9GCJXL3muYxR
88ntsQVSSlRy/ks+uz1L2HU0iqgoFULrVtW4OmDJoCpkYVuB2jEmPp7gxyrpJw/H
RzYfXP4ndjUg8vcFozpbxIYykLoo48i/1f2Ob4fSbNF7uyiN/NJetg1t2wkINAIO
OlVgje1CXLWF4E2HSsWunt5RdXCJyULu9NliHYm5Yj9+3sY1xBikAOA8in9eG04l
hBU/K8+tHhwWbWyv0AufemnBp68HtT7TDN9Mz6k69MdvZaioHt61YBIYm6KYQPnE
lDN/6PspMiyNxUfepqjKNIopgFCrlmlWKQZO8zh7PfnRnnobg0jVr3cT6bRdescv
4G97vaaa3lriEoQA/yzybiFxIJFSmEZ3F0z1y21wSw+aB/sOJ3hu4p8yK7vbLf/o
V0jl+MxWg5/pLhP+1ul8E3MpTJqvN488MfeavddWvmTzF+Rx/XhVm16/LD9Tvfnv
dB/iIzD468qyXc63fQcDzkjdfcQtDqVcvP5ciz9iA3FQSbxxn/LKmXocY+HtpWF5
t5QQO+Vn+jlpKeRjo2zghZbJ1xg1JKi1LZdbyPcnK7T3d28bRNMRPSe9yVfNV0jh
FtGbP+/KnRMB1YU7hdxnVEPRZJu76d0lIUjRqfVfBEJgRXr0zAlRcHJB4wRf1qJC
p2YkqbwjyYMGvqrP0xyWD2hrKUOT05ptqDUD3c7TKGW1sQYwzPWTKq6kaUdH0Mx9
sXXr+Fm4G+nKKHijqlR7QYBw4z4lPyGGvOlmUN4HosY/dk55eySKb2AnyfDyvP9t
tE4ZV6IC9P3v2BuecpmyqduVYrfwfXrEJFjOzbYi9wK2s7pHOradEj0YwpCGnr/3
Nc1LiT7ysUQxxGFLjeVZKeiJpM/Idx336IU0W46EUwOcPUTw2Iz/PLYA38x+wpFy
fTDFaVGGV1J9XSRdWJMgecongLISQs9CHDRpixn45HUUxPaUlqrHpO06xlHxFUX5
PdY6inqb5D75cigXEp4g9Yab75yltjZD5YcXOO7RjEeDwSDcyg3fmSPalrdfYFFF
cal/tuArku/3DyQPWK8jgpkaXZdMJe9kg6zFis6HNK1QlbEd3Ej7aQ/eXQyzqyPI
c+thtX2dPxEq4mg/LuJTR23mi8pgxTO6P53JySr0LNpBYF8tQGOuZFKHfOBzVB57
rPqG/WqcrWXGa5qOAlt3z5NA34aFeL4tZs2xxTl+WV04bPd1aUts+GBdcvxhmSA+
RZSpL+zGPPTgYcPUTZzl4KElUO6aCAmthBgrQfOQgGKvOBHNFXKPSQGW8j41/YAd
gEJ7LW4+E5UqXcKPXAUAjnLxj0Nshnj5t2qjfeJyRpOYaFVGOqc7pQqjxk8GjGqH
9cRyeBST9tHbeqtnZkqBeo8H6iNJAMyHtLYf18k2059Vww1S676lp5a6QHMzU6EN
rPhFsazOQOSMW0NiiXrslSazuEj8ZnqYon8c/EbR5VxmNIruyzerCzRaWuU2unth
ohKvXhFrxGr0ODOfR6MebBY/SG41q38pN5mMPkuJEbIQEdnkEQSa+j4ZfIzjyy+e
77XwfZpQkYi+YHEekMQ6ATrf4IP6DpvlF/di2R2qJYSpZq2E6t9CokLTw6slQ4vu
Jzp3TD79m9/xi3N153OF4T+Sl1m2jaoEIOjifPDkL9Mf2GlQBZpCkn6DjM5V/rmW
oquyuP2w3NSUUJlSli3p3RSuCVLWs6OUDZGCfE3JRAhztQwg4MyuA4+wj2olEcyT
m1V8dvf+/auJoox1E2AzzBQMz6K9nkjr/pmx3zgQTQH4cd3IcyMMfjgI132NkyR9
POBkgCHTgpry1BkdLGvmNL4xhDKD2cy25jVz+gkszsw1XKs89w/799fn4TizhkH5
HxGZ6qjbBnKB6yaTlqmHQOhFeX1v2/t6vT8ACce9kxjS9WgebuTDF/zRQX9Q4wwN
qbx55c4/xiNRm4P373067h+8g2C/km0HF14lSboZP2jzknQVoIGwHvdHKH2dN+ah
I0yAno5MdbRVuUf8IQxOVpzcDsBt+ETp8YKk7lpguNHgBJqaeJeJ3Im1mUKhxyt7
h/cIlebi8FTNAu/vFYBut63CriYVL6mgVHytHeIPWYxEngLqqTVXmyKDJs6e8y+O
Imu7dBQ0roPYtKvgvFGTpZBt7pWc+V6UQVZAqQpymzjRAUwtsdCi7nDO+c8cHxwI
7Btjhh/a28KKJuWat0QbqHa7R37wp74/A7GECKwOI9RqQer4iUIYxtqXbqXTQT0R
gXBeQo5p0Vus3lXKhu+ci3Voist3389dPHyICKcku+HokzxhxwH60flc5XwKXDYH
9vInkPfE1jvfHQLFpOsYEgKtV0kIwDXJIvc0yYL0XVRihlNZnJQSdZwX5Wr/lRFB
QwDdRGsvKzFkTqmy6EEmEzwc4/oxDbtswxKcjXMuLkDu4GECLAfvSm1M3FrgN58l
pz0FWdoKxZyXTGA4/SAvrIaIcsNuli64saxU6x7S9kRi+sLrz1EsSOMATBi57/ly
jHwnSnE9VUunZjgvFEbYgCivvnAJueOn+Xg3ATMZpYXzaKil7sFkiI9degPpo/ch
ZIbPe95dn5UClL6QiXs6ogKCpPQN2/LTJeQncIAkx8/Fyi/KrH18PWlkRbijNzeL
mr4vfzPaGDmPvKRymDUTj9TnpN90A2cdH5qBiMNGVTon05sZc+3c8cc7yVdEbrRH
gTPGnSMD0EKmjDFCWmr/VJxM0wAaAl06+/fRIbnjTZjdPnO9U0wqKAv6S4oW6ioG
YlZlf0TnToh3OnfqGRLBiNZq1Ko6o9cGodLoQwuLRpbu/EU0hzIMh4V4KpXVXYuj
393psI25CE5L0eG7ys0syT2XpAK2sDxR5fprO4yzhiZHRdQELSv0Dt9/9ckdRJKh
4syoMJ3497eiZns4wFUUFcwh11MQY/X4LCfQ3bvJme4qWrfxyj5ZyN3ZmxziQLkD
pmjspjf0RuSidsFWdhzfLsu393Qb+uDIkqke6wbSAgB/f92XW09+6CnyfdJDPozM
iPGalNhxKQkcF8YCjT7zWKfG082mYZRtmnW7s4CXzGSt9SXy9bKauKjBwvZPYfoW
+osmOxK/8TXsQ/MSS8PsJOV5WeQNRnJBByHW2TGMDYlAsQA9VD/uZ0D9kxQze/ho
krptynZgBwRZKTePVOvZcQthNTfHdqLzeT+puuMsY9dWrTfAMOobibtuFWBescn1
AvzNi1xEzGmdMiJHYQkFg/BUmFur+gs/ZeBk3QLDpfanDhiN4sOI6JoZx3KnK7VP
HoXts769HSMVItOUOMXuVCOlEF+Ihw/54suiSFko6na5shJRr0ax8l8UOVk6fBUN
oKjoPgeKERhM/rtkeZYGOvSSRJVf4/P9Q6B7u32jTM6HTTsaeLwrxi9cJ8w9z6QF
5Zri+YEw/ZNDbw/pdVeKwigOXszClyZ6Po2MHcfrqPM0Q107TlQkaT0CTdV0ctwY
7V93NxE0dch2UV2RsYYVMG6zSKcHZt+MxRNIEAL3uxj1y2BTie1lRXl40L1MDSEZ
rGf7gtH2Us7g+nVKhwWcVOjQ4DrFayFN/NuZd+wAlD5kZxIrhpMq1QrOaX6MKgBf
ZIZhXUSbyV7mh5cGSYX1IKZhdBhc36hrwSon5MX3grwmyEcIisnABNJaib2qFXeT
BqnZI5Jt92PDMo7VYrJal9ehe6uk7bGbzKP93lHY6Bf/8lCwAiBWZFE6dDBMDrcN
SjVb/pTBFWd2pgZAAWjpkzdT3WeL3tMkViLZK5WzMTllbxNzIAmhlWZzOZNqV99i
rU/UMf04pQ8MLnyKHXVE5Tvuz5RyAKxpuscsdbgqtSInwfF9FqDptlyzdlM6kM+i
Uil+XtgPi2sA6PXNYvXiFt+y7hlZ5L+G22MI2pb1POXTfmMoWZSARjuyYfuWH4yy
Ayyh+AFYq92/qQsNeRDeC568WjP4kRICCpLtp9JlAlGGq09a6V8AL2ZbIUgVJJBy
qMn39QJsQQrgvyNNLER5EbV2q/73z+ufOqAGz8iZCJ+kv9xEezhnvqyXyk4yOhgs
4RXP9FBdmh9n+KNsaxdGwzHV54sU3QpWBV9975cgwWK9Ey+ghdRaKkU9bksksG7O
3ccfNxZIEDlbPousjOCFFsXQfAMklDAQUwUxvF2fKyMqsuMGbSL7CNicxWJb2U43
qPbmRhzi2FGPXqcudfrm0amEo/kX7uqgDH0xCaIYQXBEG7+k+KAE2RF7vyH5U8IR
SPpnUEim5R0HQea683gVpVQqyVRktY7mHe/HvUOYhh6nQl3NMD8pZRwD0b9obnKC
UN5Ma/7sh4MJ+J7BUoSm8oWBNr2ioqTxIdxwSwmSWkbr+683EFK1g8xPfIToS/Wg
n9aroL7BWAf07O2Ct0z5zIHxhVi0lOs3kfxJv5NHGSAbGIt1DMGnPeaHpR3ppTir
qz8XkLnvGqTQy2Mg6jmvv2dHhAYPCGbAee+DvV0MXwH+YIIRB11oKB7jWck73mtd
kmTGkQdHv4cHNOZ6tIQaTCqwxCffdnFmhVOQA6Tg40KzWQhZR7IygPS4mtVwdDgu
3Y2CJYzkCJqvJi8e+rdVuyLutSo6NGRnaIP6LYT+aRqXN20qeE8Y+ft3mQ33t8rO
8Ft+jdWH0eGGPO3gO7jCq6QAHxdJj+pPDFyRCZsDm6kmTHAa0RGz8l+Rq3F5Ybp5
OI4hK6lf/+RVDR69P2NlBE8BnETJmQkZv84MsCzvFZ58t9+OnTrhYi7xUBDs/600
7XrT6ASNa22yXh7iSX4URCgA0M5x6ByG3tTodzEWp93hGK5Loi1ve8Jp/NM5N6t2
UwfUbEKu+MIoy0RbRIva3R3unmjxZaPsXg0kNQx0tO5eupuWNDIP+u+XqqUg57zO
n6AqMy4NSHMlZjAlvqONTClv/YFvLqq1W18OR5MCRszBDdIhqBf5v1Pfmkx9bjT9
94BDlddUJdUYZrJoMUpvhcv1P14xWTZ2uyDBCyDkGU4mSlD+Y4mauK5v3upKVJf8
wfCv1JXx9/k0A0PDueb/4ZT21LdZy7r58ofu+ACvMBVPLcZEQhsxr+4t/B16siZQ
DAWFTwOqP7yK2XqASkI4SdYyUnonaimC+M80dx1YT3XCWTUed6+V4/A1XTVeDLj2
d21kkO4GhPJl4htpeYKexcNYIsU6XW1IRtm6zsDA204gvRkMTPZLX6BItd+t3UzT
iQ2v/mRQu80i0k30Ad1VGwShqyTUpsw8VM8c0c0OutgRPh9WPbpMsPSMy8WZ7ZSj
PCCANZMQhyp5H0i8S8gtanQYr0JwTYQHpqVD7gTHc3oxCLEW9Tth8EtcHSconrQL
kGbl9wsTDUJ72Z3/c9NA4IfwnXJX1S4ukNowusfnmEdPqehwyGttzoL10eIXmC6a
utQvHYz8PWA8/jsek+O5/bYMIdSVTfFvPs894O1o3MCZ1iPiGtMyXyAJAQsuHKN+
xz7COqgeCz3NJUeM5DqlZ3pW+GuKi/oA+QO3i6NpgMghkMSa+mxR9T8ki9SrXknk
c0J5ig92Xmg2dTBgz4O2LXcc/PQiOvmIRmrA9HlUMWWhp4qju8M7s5vYWWHwmSAW
59ebva6I/UKzCQzapnNSoQW/0xb1WVmSBd38Yu3Q5Wh18rlBPet0PRdJMAIJ4ZTs
2cjND6zR2zLaMSG4BKQGOxcq6E64pxmGF3QFnovVxzVgcHg6GE8soDVc0BwsHcNi
9ACrmi0QbEfpFVKTL8GrGTEn/HiPA+ezOwhb5xs0YF6qUyVs+U0kPaNsVW91g8bf
OZGgUZ8H2WqscCGv36hURMadkONCS10dZR/gDhsc8UONBnKQxUsOYh7YX6xlV0C2
FqslCo6g3PXf5iudt4kZBX5hRce/W6N0PzgcKwMBCx4unZHhuiSzrCAstenT9Gxc
9MVOzfyRQ2Qbze2D/cSIyAc3lN/UPNKL+HHkEoX4i3KVvruAGEwZ2g8+n1YnXtrF
4arOpw446h3R/ldW7Y0hEv7Bp45K/aQ16EqnkaRYXzzvHLMp4nBMBAZF6VLdYdp6
9pYdbwbBa26v+haWkTcolErUkNmFm0lg+g+LzFMhHmevSOLl5QfE7q+cN101YbfV
a3l/KRr/21FkqsvtTl3wNcrltQhTwk+QRdh0Irt2woDP0KKtv6vYZqSLG620z6Sp
wQ9RnzgoOk2paqF5/hnewRAQ1AL+u3OzOOpmhM2hcQHrQQNbdOLimk8Pk5nx22eL
livi06Hq90C48mIfGvwTtAxN5KpQYV+nfTN3GxsU6Ew//1k+rL1SvbWItBdyBEGU
G1Nqghq0cCDfmpm6FRTk0Ne4ybYdcbfKptuiWnU994yL2yf/TPvw5RfxmJd6M7JG
uaaypmLH6RD4E9MudFNMKtpTs55MJwdZMM26RDz6qGiOhM5B6wyoK6DIegBZt6fx
RAp04HERisUiBpek9o2H9prd53tjDLgeCdJmCgduxscyvkgp2+igNdz5FwdL0J7f
RpQNa3ycvvvqOLDCgHsY9cCU2rWyYBHJ2O8SvdsMskjcMd1ZqQ9owHTQVLka5FJf
nAYCet37bilN81TDcTStQRVh/MyxWXyYh7e7u96KOW083ec1F0N5I8JwMKIEmuPU
SFobCJF7BYCqTLiTQc8NVShupkC4L3FCXoebK6ozajH0Cks3u/gNAnmI+XRzuilo
NqqUgU9GMOMzQ7HFor6i2Ik8FqBNfBVSrV3Tqo1DtH9y4G7Cja9m0knJP0yCFBQ6
Vlw6aUGDCmVGv7vZC+ARi0pUu9ETxt7Kr7FGLSI+gbVJDlMzyhoxvBAHj+CPuHsr
q9sYCwOj6krgmiqDMu6fn6KDHYDBviyEH1jZhL/2HK6hSkHEpIzaZpJNwg+57eUx
LC2gzJjECmIAi/GGOlaf7qJ6KBjQUO36SJNpCmAXKscHQ9qBnQRlGXt2vfP0wogi
Swn5cGRYHHW7/Xm+t3KOHhr5/Hc8em8t8X2bKpFEfV7NeJL3iKwdCwDjJEivjXmv
o+NFBnObsnyJB2hMQTbKzDG/kUcFHYJAUStobR5TrZXC03br1PXVrlgOxvG8WtmN
rQT3YoN9WZgEGhGg+QXs/7ymPsSQZcoVVv4lZvxppyVjTjiVacdvESJz8jxQDVXV
7e1u3y0lXXCy/85tvk7Y/IpQvWp0Lv4oOCFDmhlAvQMwO5AmmjnaZ4moZYPDRhbv
kA2CZ367dHLiWiWPln2hpuwjetZQl6ful8VWNl9e6ELklIb/H3UC0eZ2FUFzr9X9
zOTRX0J/mVHOJzqt3JlttCdpw8pNzWfxbe4net/XW8QvomYyS9aLj/8qfw6UzsBJ
EbrR97UguM7UkqYhhvqjk2sl17bx6bnmfu8P8gmmz6rg0hXoHjjVUcVZv3z5HgND
Y67FsH/aF4kNmDB+kVlhYyCvxFpaM5HIFjoB8G7OEjbV07eqs8pR4Pfmv62T3vWb
tWUyT/buQgammKcjQjGPqenS59QVpznK8puQ6ZEmOI9VEN+OLl60qvowXkB/n9Ws
qqhbzAIFzurqq/2uqXS3f2+ahy/pQvuyMMVQaWQgT2jTt/LquHMHlux9S89lZTpk
z5/kphmvg5OTUr6rBe0Z8fNu0SXPBQ/SBx/QW7cfSKSyR455VssuSqFaNRA7Gpbq
d4lc4OKICeJYVfo4e45qysWZC7myE/ljnO5zJmA09BVCJHfCQFSP/zNQV+qSnDA7
l52GHYO45UZV5umNmrVLyY8VO+iPXy2yzJQ2AYQ+49AtjBytzb6uYSA/j2eDZsZh
aXeODM8s6wUK6esDOzlLc2L5Z6gQORBXGlItTdg71nh5xNw/uOyuky9JCM2tPI8p
GijekLYVZiKkXqqZz+Fyg/SzJoLD+uvLMYAaWedrAzHgLbK5y6tV1Dz/f7gmiEUd
GhurQBCmwV+rnzYMZld3i2O+RHrzmq1vAv0dJAbixE1L51MtemSIm/lS6pkToiBd
+e+dk9r2QOsfFINpgG3J/K5iQyZDIosyy4CPDW7H27GRzPzkw0zUjzKS8tJUcAXz
T3dRAGMUk+Ut1DXU9zXwngkqkO1X8sWLXmAx7qNLSkdcyy5JHIfiQPBXQCl+HfRX
ijrNzScEd6cowqQmXTveknb6KIGr95nYFXHLSxdOCTNt4l4wf2h5CtNFti1oBSHt
LOj7W6qNjJpf7GELKpqY57j9soTeeWIM80D9n1xgdRm8VLL2ikgh5W+bQLfNv8wf
yVzPye9KbpZwlfN0C3XniTUGIlPUAxeW/wcz40GM1l2MVA8k+4lFlGorOSxQ+lJ1
CIsKpmCH3tWhKTYyiHwVV9jmEFmN8vGZQw/cs19ZZBpag/rwhR0Pgn1/jVh7aOhU
E670oEYdGxgkRSjvjP9yrpXcTjyZhpWh81Rot0sdeRGrr7pNaFuJG4pB/ZH0/jtB
2DSenbf7ZzaMHcuDf2qKQOQ19Ng9xOtCAPEww1HAiea0JwlYoEqtXYzoVh3YvN+p
4z2kYNvwXHzWk7/6vpoGHMP+FcZ6jXRJdMN857/K2wrqinH67BWWwxoO7RsqhKYG
wK8yALGNEvY4Y5+WU5SQXwf7eGykytgLq6t3Y5GljZOwm/QdMH7ftNH5XxqnjPZp
l9swdjGTYcC9MjZ277APBKmJa3DPFMCi9g41MwJKfLUD0/si8PqcNETN8Zx9fiZ5
pudk8o86Jy6iWFEkPAHbNgs5rwjwHfVxiVxK1fz6w3pcUPvr5ROR4jEwTgCsVHIE
ct/Fboc0m/d2QI6+Qtee4ZJ7GS7PZTrGSqpHUKj8HWbJ9crAkZnwE9wK3bKx/xAS
Z804H2ZZ4o01KKpT+miWozUdNI1SHc60PwPgxXoju5udnH+HE0ACo5HIx3Ua37N+
XoTvPIOOAM+uPdOfcGaNUGC7wkeBO0kmqtQZT/uAoaB8dJYmcu8i9Zg027F08wDZ
I4EYHAR99iZVdnf+COMgohNpM9BDyN5S6+P+AqpRAjeSAjuVdRQNjyjqCoRsLJNX
1E8wymZSViCXeY9Mq6WWVtQT7t3GJVIAgRCrpcfg3BD0FC16kbD7aKpYVFIbzCil
653uwe8M0LGWxdiq9mJvU7FDlVemNbWUy1/KnzO6z5zyYGcS3mZ1FRq4d3A1Ofb9
nyt/q65pVYOGt6/7zVKGp/MGXo3Py37BfH2BjMIsDMr9hoCXRhP1HkNTuKAbALZ+
yaB+Zri4s1iJZjM1pTo4HFGxvmiPS9yxoLeMhQuVlkLID90wFsXIa9UUBR49nAdg
wuAyfL2OEfSxbXk3fSh/l683pzJjvC6z29uDHBwdabB6VbjxKvtV139rZaYMoJiU
ASwmanAxh5Oy9QTGg3gp6IrpI9KxW28WYWHn/YhIp6xmBSmrd/78j9f/mRuaAW5o
C9LAXz5mTj0bff7Pgw/e4mVWH8Sp6i2t5iHY8cAvmxYDfgLZdKujW6MacUFI/dqd
DAdhorLmJMerHCTU0j1wIbi8RB56uEqIf9fGsI7x9mOwKXIXbvnmEOAHfGCWniDG
y8a9j9bX0i6I+/Vhx+2SLLDQ133xLEnBOBLU8P1X3emqDTRvzb/VmiUMQxhuY8Vg
ItbDHPIS8/2Jyi+0QyLaRMazz3NtJQi5qJMurfJogEdaKmAzrNFRRgM55btI+ZhG
tjMEp/OvUYAdA8zUmapSDC4Fc0EfkThmPTW+PtFCShcwZqcv0dbe/cyd+3LDv1uq
vI5GRcKCRMlM0tUL+KdQWWsOsDsHIstkliItVEsM5MvR87N1/MYdnep8D0jcwE4r
xhzzU1hKB/cAcdnqoNSAjTg4SGAET6X5CjqMsEAvjla2MjJN8wKrv3ZjX+B9FtNO
+MfV7S8pWdVqAbz2HU6F8UFibwoDTLRdTPrCw8ILy5IhttJRCeK/VA/g2SfprgT1
rNP3hEusa86pdHd2m4+KK5ep8XR4MAUOkQoTHs0WVyP3yf4GuwbqdP+7T7jN56PX
4ijw7PIl9jC+YeDOrmnapcDFvPC4cNWnBR2Mqu8jyrGcQPO9QzZXl4IPG021kO3c
SWV9gX5pC+87vdPamb6JiikRhSkG6nh77gc68xBtYhdP+5XXYm4luCIfDWQjm4KW
s0ePPKmYzfid1pE6UpmrFAOHTthCNyxX3xP/ydX33aFOmEk8c9/Ob/Jfwwu659uF
PRIO2me+C8/I2dYxj07AJh1pgdpagzGVD8hdGoy8NiN8L+Ew1KLUa/wSKian7YSM
EhGyYVzpuP0E2RU5qKVrKs+NDfrWB+SAL2eJYDMBLUCHaBDDVkeoJOXmS4YvGd0O
Cq8+xyHBVbEQLO4k2IRB2KpHuxvbHBa4osHG/Djb/k75mSNQejWoCrGAlRpTz2s1
z2EMNpGZ+H/kqeP42gTO5dJ+RbAn5ytaZTRXr5JztqtGP8KEJsSo1/6XVgOBvuz4
jYR3tAPfpRIivF8seTizCrx1bHHp5oWvIyH/4RHEgQDa6mwEdCnjQgdMGqpovj2l
R/0gv7TX0dxiePAgzJZGIoTTNnUVNJ1XCZcp6qJQAQSJjgBWPEli91uRE6N2+Hzn
O7jr+CneRMDxuiKdGfTr9seed99zSTo1Qa41/iU+HSGFoJz0U7aYbixE9LdcGzNE
FtZTE6+YHMLgtb00mTpyZ9UWXM2JPp584blFCtBJhkonZD/8qNNysLbLcHOvdp4D
HfrQo3rOretkcItm9Uh61c3g4OOAqBUfmGuXBjtkjxlIs5AI1fvaWdbcRbMY0tdm
MTIKt4QiDC5i0dnS39Dh4kqbeL4HfiYioXwNjmVoG22ZFNcEG9IJ1LshVBrLj9p1
DI8i1VeJDiy7jp+ll1l/YEZrgF6w0Y9fp9p16JY9H3FXn3cIlmCjR/6eqYhECdXx
6vFuKtrzQHl4MoMeONn+FaonmynQh0eC4VjA58XhpS8PN1/VGd/8hn0q9qKAVxn8
T9wwluSh6YsrEUhjPU47ufl/BySdOKE2CTg/+/6791eEjKrQYOBiCCAQPAtBSOPq
WwkW4deeuKIYcRCSnxIbtTjRt04MU7YUsJ5jc6Dgucw+8+orKWbkqQiC84nXUbps
9c+n2R57XbzL7rLv2AXZxrhLIUahsqjPChcTqhG1kNwMqH8Twbld4uyvJA2MFV/6
kJkAPm+WgCjwY++y/kRkGo2uag38nDmAIPsXnkRkHqk/21KmvRh1oFg3pXfnk8xg
EcpgVkQQ3S1rAv5EOgbE2IlMXv3mvzmyAPSrl8N9XL4M0cmNHe7ffeqgxHmEtJ8H
lII/s7oBFTpjrGojOw/zDgXGHEnktuwsuYpWcLTszOW0zBPiXidEGmXPz/O+FCcc
1OW5FZjqpAaI84zcvN6CnU5xPWR676mMT4Rb3AMwoFQ6VbHlq/wNqs6NdqXIuXzN
33a33k4AuINJJwp52+eLHl9Lxj9OnVQCx6grKKM1RsHRxD/rrH6KRhtdToGGRFai
UIKNt59y+7RgxsusbjksCd34p38xOu+xQ4Tcuxp8hRQhq1PZ0R9n9kSnJ812iPeO
tWKkQIIegqBtoydA6Enu1NjBTa5xz2EmMOjZUqkjVJD8iu6LZ6Os9StSjDj8Gyg/
6+uySYUlwuMfXy7pDvNzfmWzge1Pa42K2w3F8yJ57iMUUCggtqKx5avCl5hrivjQ
7aRcsUSbW/jrbOVP7YBPdtEKDGzfIhPShR2aRSn+7qLApaUlVgtdF6BEPeCsHBLx
k+T5FmNlsKSRNvvBYBcgfrtPiX09V3qO/1v+e1hsbWcq8dMLOOuA+ksbpdDGYSRL
WDv0dIFgo2K5Mg3tCbM+ftghxYJnUdRmKO/IWweH07A+Gt3iCWpM+7JTrag/4qRD
zvPbMyziR2RiPt0wdQozxSnKL4KoaScfJOj2FY2GqSz5qzQvy2hHulbyIBcJ67Il
7oq7Ca+tjX+7Dc8qWuFskePFby5b1zt2QLuhX5oVEQtcB+vn4Um/UtaNRLDCqYba
1eVGtkMJywpCnCQDX7Wt+pwUjdE76f+chxKfxfDW6KLJ0IGlv7XvxlADvqab1OFd
uUrJTbbAA367NVMImz6WK+RB/nZiqTvJ1qC4fAeoF2+4IdF3IXmk1ladUVMzZMGs
bxM504n++tAe5Qaw9EbTMjEP9/2F+f/zz6egiz9TCQP8xHIdbGnWPqcru1VJs8to
mvuBXwkAIseecknDLFul1msiO2u+ynUxo9Hya/r+s0DWuUOUAmV50hvKrwGqyhiN
GnYArotkZNod/YsDf8MHVzWXe9j5f1Eaa85k02Rp5Yhf/9J8LAh0PHdK61hB95px
5mUADnGFn1SwBZl0FJ3z92uh27ZwY1HmvKWytuuYlJ6FsaKa+ITaspFWDlUCwOjR
5MOL+HVSXKBTcm/nDeBTAf2E8h32EcZd6aimLtOeXJD6lLq1gKM5i3cuQfkdFX5R
tYfZlfUVUZrd0C7IHWmRoo6/tlZfcSe9RObhnwbiyOpLD1aTXWiS06I7wvx4fpQi
XTwj5kvfsIqncH1NGcIozvlAS33Hhsy8+Y0pcuw4OTqK6Zk3KNZbuDxJv0d7VEbu
z2+/+UpvJHho1Mbm8dyeO004XgqJ9E6Pooq82esCVQwvz9mWtagyqDCMrEo6refK
42pDys97edbdkyDMADxGSTIpqd3hLDY49JjD1j3acVGCZnnnbHtbPtgYj9Z/STDJ
/HUlF/tFSID50bHmlLaHeKVWalivrjY66MmtktBt/3GZGaNZ/C+/cRNUulKB7hBX
25V/sFPybRbzwOi0iXgcsy1IelDTaZaBwJZnx2mrIBcfPwJIMrLmcU6dX1fQinGP
AocKtNi3QbXrvGBtzp7Tedfkg/CXK+bwTJz6k4XUHfja0ikdO5Tlq5Tt4RCV0PTg
OTZLOcFjTdIykW9+jIW2mhrWy30Xjsn0eSC6HzicrXGDTK7yFhGxOOcA+AVfa6Fm
NcszciSexbqFr+8QJs6xwnht6l02KjDuo0GZxjtTNY1K0KuTNo+I+G81iI6oYxn7
50ufIt9W5Hd1xzxeaYFG2MUm7hA+NcMxzeht54k3OTPIqCqWV0PydWAtIRk0yKse
LgitlpVbXJIvIpnVhKUaPgLooyyNaVgLydBBfPqBmoXPXZJlGYkROLZM/yKlt+E8
IlE2fbuHJtpMDH7tk869ucimvsm3wqgz8Oxb9Dr0bJ+t4Xp+MByHAx52mLbipEpu
ruT/71WeB9XuFJNqGombf65HSqHF7n4eOwMZjcymQJiNyniJ9VS3hqwa+RC9asUU
wt2xENqsNKP0kCALbcQxy9xRxHHq2tF3RGfZ8iKJugApb8uA4hZI/E9pPerLqqO1
sz2TI10tJZ6xISMRLBj+gXCkLhcEg2OVXti0iSpFwb0SzRJBOsCk5Dr0px0RVKyH
2YtBJ1iX+KD2gHScmd12x9hbe19pM0GGHAHIRxkH5iKGYonT+e+UkftZ0xOmIwcS
kw+Lalf1eR3q8Wq1NNgxWwP1LRtloeJn+PkPwikWo4ybQJEki/2lGKXY8qxXJ6gB
+ZQNIKqOWrIOBUuQFxw6wlae+CYQLL4v8S+whG0heQ5KB7WeRYnIuwEBInTWkAh+
qeVLMKdNYmALGc8PNbzKeoGuyiZB9e9XXUEnz8OVIwbWiKPAkFvPc5FfvSinfGZj
skv0+hYLJI6CCyKlqPzlfDX9PbJAV+w1le8CBQcjWqS1asq0HqD7LJ0XBhzTLWWK
MfE4ds5zdRdp/E3RmNhL+59a7v3SbuP4jTqyB7/TlUXak090YbM8VrE4+WzerLTF
ApfrOoId72+kjdyhl2lAgx7t5bSZFo4kH9qopLgI/Ev81Q7LVK64cM9SapIHsmoJ
ZSOFI6ozSURP+LhhPlJgtPV1K/sGK7nv3w4+4rcfnS2six9RNatj+nTikVcot79N
w6rLw5G1VV5Jvlr4D3qxVUdKHSaKbBWIUADjHNgfaMabErc2JL4Eg3RGG1X/EDDB
llpKNxXtRa8tx6PH+hkHXfsBKxDq5wjkbEQKT2LwHjRuWCSFNFreIYcB8C/VJe+4
Wu+hpjmhGtnZ6s5WaHnZ8mfTQ1tmeAvHJGbqQ1LuTwtxTLoLENw1tyl7soKNIl+S
h3izTeRGoHn6WmiCk4Veqygv+pXfOC3eZRFuo7uCt89b8S9jBhmaGoVkiimwbF07
/4M3StNiaJb4tkUJ3sqjbSzcNx6kd47OpO7vQ9BX9OSjvgX3Ov/bIBLX62juH2nT
qBrmJhwfg0cCmL7wxq6asuHg2rahe81SxNl/bl6xvLoKWCXL1OqZnUvGkLee3Zoh
ZvrwoP+1+CI7pyc2MEeq5jXfUsSmeIFYq3VFFmn9Rm+VfRFfud+sIYKJgvfhLisR
uJgNeFGqz5g/ZRi3TCabCeyYwn+Lir9RwS0Q8zH52M8yMhIykU28ThU79FB0FpzM
RkMkP5icDAQrqsTP556KvK+Q2rLvrCuPdCWirJ3/4RKExlfJjAQafGOxC01AH9bb
zOMsvVf8e5mEf3aATWOJLLUD9WK8rKnaze9jygoCA5u5L7FkEBzgUJh6pBlB4bR5
DY4sJDsBz/4Dn34HGViNfTBVAIYdN50MKeTRrG7glWgClRIyvB2IGrzi2VlSrAmv
dD4P0ufWXs4npORnzhFMX6YCPLPHg7iqN4KV5bHb16h5Wzb4PyfdddCxhobLO7x/
IJyu/QeNT3lgsP8br1XbIdagh5gk4KIHj/0JPGpYOAzM+aaxxfXKOhS701nrgtAk
1SRCkH3wTE2hVC/ZBExMffu7kSqp48n5tpx1DazlZoj+hTXUeV+c6wkOr6ULO0Tv
jG5Nnivle+M8SX7fAougR5dMn/8oDLpX5rvi1cX7lt0R+aZex2fA+HX01m1UzYbq
j5+Q6Yfc6jsXX1TsvCWtTqJSweKlEUmwHOPgb6nxE39DGwRsLaagGJ3MQFKTYnDQ
8J/snyvXb3A9EXAzkSE1okJreBKUxV6erzw1Q3KhTmd2/QXnnAZGAX2L6qEQ4Qhl
EMDHII4Drnd19yjX1OodOImXuCiZCF4TveAPJu520jwIwNUiW/HVqaZ3eWFi049c
wIws47qq4GZt9u/TtM0CKWePb/+W+fOWAzjpjIqP8wEGIV4QtvTzWYolaqmH6MYy
v2CuGodYU9RWzbiyODF7xEhdKMXevfbCc6RxQkIW3aCQN0lRsngepxl7yJEhTR+Z
Zkkd9/4Yc4mhK9yMnYtgl2vuP/q7wG8e/T5TrBalb7YXOJ+xwTtzjwFtDFaLmUZE
dNBrpWjoQ4pYBqXEc5Sod9KVhIG3fl1dRM/B2z8laEzpskKxTdAnzZtwApHJTc42
q+lJvCUZt/GE509ZKRIDPWsUghFjbZ0hCOqzxqN6AgCd+ccruHZPSGgPnxMRqBVk
bxZjyKNNwk5iRGLoBTGBo9q/s7SIpDfn2aLDvXNoPwt4D6gGjoXbT4bY6a1ORpLK
DCbMWkVZ3ollnClrmMSf22jhxkQggdzKTKkJEzkCWOhm+umeW/1WqudQ6Zw5zl4O
g1d+ltsMF69fA6WHOtxqDgq3202CVBaasS2asQ5MGA2DH2U3wAyIvnqpcWrRpITP
EtruVYb0eMNAiNtenTjT7t0NdQxI4GW1BYcg7PZCklfN6OtfmwAjSHh9xAjoiIWX
zJXaQyolf1kI5DqmQH7cHZOJKCwDhvYUBM5D6gZr48VnjP/to0r7OmRIUJOQe24h
7nqknCXgZFzDh3yH+RIhRkd2U5U2aRe5WLIOVeo8dPKQ1kTY8q4JY+yKu4ML/9og
NkVXvvpHYCGbBPBDgfScoPHwFNIhG8ClerzjQJ3OlXvEkjp18MN9LuQtbOQvKi0M
czvhJHuQINHc2ib9Z1HweJpFWHoi8hqKR5+HgvfgzlOtIxS7rCzzPyey2WpE5QAC
F0TGU9SudDFQNCOxZS2Hxy1ZocO6Fgu/Q4On1zFd7+ybTfnHpcw3atamZy0vD2Vg
FZNLG/5fnnh6QxzKTN0eKGI/08Syu3JPJ6FKm2RKDd/9bN5BjIrvfCxGhYrdPcTZ
7JQnlongnX/XQzE6Ns1Z6hveEl2YKxmpi4cKJ/jIRhyWkLXLxIu0zm1hVerzOQaW
XP5CjTxVx5uL1k244RWqZfBGL1Ffb5FVAqo8EE7hA7ojSL7iYoZHCJvHgpqeiVnt
TjHTMRKw/RbyyAhIWzQRgnK0g+Rh5w+2xUh8wF2iVTphTAGwXNfF05sb+zQzKgds
JAJUmqY8qB+WcadLtu7jyaR/PhXGLHb+ZxPHmhpX+SiRjtWl0G4QEjGI10oGYN+0
+aFX/R7wj2S6shkKFAp/CPUjA44CxG5jIUrvM1b44d143qx6504YGro4JnBQwgGx
un+67QNTFbIO4jM43rKkvvGjMimOeg92o079LlmnKmKI0ypLETn0y0fK0SyQCmZD
AYmwMvNsyJfEzyFCx07g+MLXBDqHvrXcDp/vBkMk+D56KzBR9u90B+yugoeSzNuL
oHJCJP+aj7RC5FdiTl/22YklltYkXxttrvHmHiq9DSNtb03uCtdgZiC3ktbn/Hlp
eCQoek3Qn1N9kcLtexi2Mj/7BqN//yXaUHTyrNoiqgMsWbwB8F/inxRr7LJZkViD
bXhzGakw4OdAtfeEiqE7ta8fFN9tU3KTElSRyq24Y1fD/usZzZEWaALEmc7U41WT
FK+IK366wQK6cN1uLWGt5f2oztxYubheLgeWhLecBWzMUjQa8N4/5DW1G+wWB5Dw
Via46NObalk6cxT2ybIGAaeym+GnaZpYMWhqnfuwI2pZ766Q3wnbOuTFFARy27Tm
vJpMoPChzM3Behh+EOdY0N2v5yGZandUbexjVmuRq8caU9G++mJGjPhMS1R59+4c
kNSdRsRGe026L/LzMURgf9UFBIWJOcn6wg4WemUSF+OPzLGy1jUD4LF6H2KeP+RY
+cfYZa3R6EkH3IzdDlIIkdk9F/PFeZjxoFfMsuVjXHE5+aQjXn2I0J0ss9xio+xo
H18fg4JjVaz3kOX/fWwRE4WRnyk2Q+4deCye7QQqipcp2bYfzfaTjjvGNVKL/4Tu
8QCHtohqT/QtbWBm1mrncYbV52CSbgNYTqJqeyJd7Fop3xyjWC6k6UdQCBU+SWOQ
cPJt+rjp+n3Y1h85tBZKGEn//O1ASWlwARq16YiJGzpgpP+/2Xb6MHwy9KJEJDJ2
p38HQwxiSir1TAnk8nzU4vmTX6reb5fPQ+ObYT0VOn4FRH/tQCRasFeg4CWxg6EJ
ybylHwwLICBpYkUOaChneON26qSITfN7LKogVuiQJAH/WAsp7EmnSjdFQAojpUP5
XMgJxRdXVTuIbaYncjX4vbODjdNtWr9jtfd/Bgosn2AVXk9M8r7tJ9TrxCRDDG08
WrYjix/aMSfKJBDdX3gtbDFQH6BAVKLwUGBJ9bfNma5AGhBL/+3X4YKgyX8PpDCl
iR9aeZNqfHAj8R9LRT3yoRKb4c6NAmf7nL4wNT2x9pdKH8SpSYhIU56ZLCHmuDT6
xzk9swyyIvzB4Xd0ZmOoeWKj5mDzGRcpUPlvVV6kycky1EhOGB9Vk0do7p7fbutV
2BflleZUm4OKBtfQpUFtBu8rUyZFJLBmKopCvsEok8/ZWnwsQkWH7c671wvVSZTB
Q76vnrXpX6BqHUjiQvQEjn1yKq1QiLsALC9DE31UE4lDx0GDe4m4X8mTpNeb+zVR
9yW+i1se26hE5XTuajcZ4MQRETtlwbwWrQRYcRXhudgsysTNp3DGnZ+sTjSMjMCX
9lmMl2sZ3grDS9n6A0X1zCtHF0kM4VUAFauzsDPUy2nwu9pzHwsTXDnHWJMhEyXC
OqNiZ1EddCnHRQAp+zk3XxT0vklWohwWn4nD6GAz5MudNH4r5eRRXyZgKMAH5ZTH
yZihJS7Y2k77VvM9p0DNvvFxS3t1uyrzoTN6FsHJ9iNGs5wkpqfwJRpogp/iADDK
XuufEa2xJ70VHiFWzr0BR4RaypBeFgFU7SJNmhQhIHTzunhjMvPEl1JF98rBLZM0
1P25S1imj6nl0ELJbEm9ucdgvHHkUwKa/nZZnkXhgZw0RpQUmzZ59Vk+z6dzBMEI
NNx+G2xuo/chDD/7yYJKiJ/VwCQnT/WxkGWcaBQ/kadurj67YWCEWhuYF+p2JHwx
yIvLvy39pqnPnywhCRBn89Qfx08vLZJTVK6LHdu0g95wAraX5xZntz8WEwDrHkJn
J8f4eJiSq2M0MJ7K26BfC9lpiQgFjfA+VKbjfnT6stZkxG5yG95L1Eqs/XrV+p4a
/ERYEBCN4+DXNN2iHkiuDUfKE2buKqka76svZrspd0LZOcGhnLowT/yggC4ni6EF
iIU1p8fooIPjc9TC0U9bwXJB5GnB+Bk1UwJHZ15lgxCVuVrB0lynLuQbXRkEvXIx
0heuip+xtMrimRC9Oj9m4YdfLwTL7E7biVx36cqsD5M+J866yGPR82nEki9PCMRy
pA0fOaioRE8nOPte7NmgH88Tjis2OVT3eTDny7J5uXY0RSJ/D0FEVs9KVM6Jiqke
aAQSXSyFtJ3gWfqP0eASYOoB7IR3x3bCF1stdHxV74blEm+p1UekyrYWTIEASOXa
Lz6E9akZ80ZzIHLwuh0MF2JPSSoIigInASKzM/44H/j6kMK1qSRRqzqAbIDq8ow6
v4cAc1N8Di3/WrZtiMap3ciCDX3ujdMLpa2iqv4v1uYYwLiEk7jrF0W/TpEWPL8z
DZI9ZV/dKI5ErmpZX/76KRL8YLtVQRVXHw1gqmuBfNFME0tcpKY9iZtix6Vi7SMo
FDGR8zfcz6i3qRnZXSQZn0YHsZpUnd5ouE1nMy6OIc4UqhYeSwvRwncjv7r1MEoR
iHsr5E30THw+1iNnB3g3CBwMD+fg05DMF6ucg8fIYhu+PzqDJpQ7HzNBA5H2NxIi
/wYRWrLw9n4CEKrNfOdZV222lf/9ZZDxf3LY0TKfjBNcQNlMjvcK1SsBPWokqeGi
sfB2UUYDGp89Ae/uvDioK01x1mmx2VyTDPwyTkIgIbISANOp9f5s5WNvcCaZ3UbC
4KkPNIuZD3TGL54SM3qtxoxEc9t8NEIKhoiaZcIJs9S+P27HsBCCQxcEXqsGaUWm
ijUA8zxupao5SlbRbrqH88IreEG/hODrfCtTgiUfiYmlXwJE86gB/VcWFubDWIyc
QANdbDDT4RGQPsCxIgqth/7H1gohMCXq1/VVcOzJNoA1vhP5CKjBC7MqbDS7BnV6
RtrqHPFUOm3eo2viW3juhJ/eu3DIHoKwEelfUk/5oLOsbfFyHoqB9QCyNx2Y9RlS
lAjH9pK1MGbYazYfz/CaoBy+SCz1ncY9ckikNPq2SilQ2D4WIcz9IeyHbcHyHx0w
ugTPqEsvXj5EeN8udNPYPUBjtoP/WDfKfzX69+dAeHyyO5Z+jNPOgIXe7uNn87dy
t0HWDK0OD5Q8JoGiZFWKnL7ZWBukWz2d5ln4C9w+rlGaUo24Hs8vGxOQn3rqksjY
jSUebpe2WwNh8L+nmuQR5tnUR7H/3yon7c0wN9Dso2nPb+BS7EPtms6IjKvj9NnO
42Hs6H27ADJCe9lj7CmBN3EBtHNAuePoR14jpYFwXJhr/8nzKFT+B0veN7gQ83Sb
D9RyJbGJTzpgcmhAKtoBP3fzBkRlKri6FMXE4MYVggpOOHmMCuJfhUVivKdetb1F
FBuWJ5LuGeGpTUJdWT+v4xaQaMwvDUswNFX66ICiqeahfVAtmKlGPzOnHoZLiSdz
Xcpz6RK8OEbgAiWT22QGtCc/ldGZADjEZCF7yoSJ9xs6l0/xFxIKqJHqTtn4FPlK
F2PP7nAwnKP05mnhBX6aWeLXc5Bs3hRvqQjzd7eIOsopBcowjtE5NbEsCsbHs/kh
6b0Bz+HBQNAnAirOCFgMBOW4QOCoCxg37uxcVQlmIOTaMB01Jmzre7PHdjmnp/+E
02LJSC80+MJxN91Kpg9176IS+OqJm9/K+JI1t3MVehHHgNlS7xpgRbzHyVJSUQH2
/rzk4YOnDBVOEBLzhbjrmg6Ov6iQSGTxYGIvtYCI81F0TqvMFTA76amcvY5++LH4
cVzlw7n9ualjYsQDhyxZATh8iEPcbgE3bLQYv8TmS3anGNzN4bj5onsevIkobvY8
R5q9We4V+rTy4LeOm+taaJkz0cLmX35OojkJb5UPP76uQzzt3LJN0zb2SaWX6lrU
L4BLWeZQ8qV2AJJ1Gf11WxBcuAOE6TGFmhNeifQTJiVsnwILhKfTA5XZygh93bUB
8zwAmHI8fWmLlUJfgNDC4Hk+IGmvO0UWIvQJUEbMYlrqT9AKZS7mRdu948/gEdux
GjCBjNg+YYsXDYby5LthaquXtkdF6IQx0x6yOcQ4m/lg9WxYNRm4jf6CEDltbfhZ
WKZhR3wTWtWGFPj4XXzKj/1blWq55Pzlt6Rxgg5zZYjdn1iLvodV+hT2XsLEn1MZ
gOlFTo8CWdoXHa9dblwBgA5lCyFKyMp/iSr/Nt3dbiq5k+fpRKV9yIxzh2vfa2rA
9VWTV2MlqwLYic76shTBN73qan1f+Fil3RNeykYSIbtHaTXT3E1mkUKladybj3S2
kyiioyqWXQ4KPssHsTxsNcuqTkeAPKPlAU/HRfM2ujs6ir8StlL6y0AfTDxas7XR
ZZac4zeVlZAcN/WwVowlvwWCQ8KWMiCvBtq1YL5lvx38KoPkjgeuiYSsKLUYqWwl
R8oQhXx/Lu0bfhn1i4X/5pDNl6ymiLoUnRMfR3DNyHZm5urIjLEW6nb+LpUUod0F
d2vzClnPC1mMhTR1FImmErZH4rM2HQEuCNz+XCckT6dcYnbrbOYnposazeL2i1Lx
NDTQH5yTNol9PJnGvbs6ZsjXtfpZfq8T8tph/lRLyaY/T3v3WL8lxkGoMub2gAzT
uF1RT0ExCgDPrMgiMcZx5/hkIYXEIXbMta6II/0fa/C/nr249heHQGzur7aYl3wu
ziBkB8cDjZooCyH/nC6uaDhA/wDY45fWGqIzD1jxTEaNrwKJt2hsmUwzt0W3kAzX
/L3Zx7FwQ5gJgidr5jbHaEEybrZFxet+7CbvGh5CV12/2v3g1pJ+wf6wCUID9bE9
j4LsE2DyzvmU3/WWOaJ6ptGyO9xxcYCspQYU3TxUCU2eOcJAXLDQcKSani2vmat4
Z21rmE1u5Bps/B9FWo0Up0ZN0M3sXpIJMRbQTVQziVlwtlCeZegLVQ6geHcIQxgq
PhWMsNqY3/QJMuxvM1DWrvKvKVCY39X8inSWqgWBcYnXAclifXsBQUZNxjar4x1l
Qdon3OyDPnKa+GKs67Yqhj/7xjWsPC12hrB3/Dowmq6nGPFGEC1zdtf8XK4ij9v0
58PTTqZDp5E5GO7nmv8MmIAD+e1reZIjHigzi8QUl83eyW0Y5TAjA5SMZZvTUEh5
NklzumepWYXglm+q4sPIbgZDoAUyGVqeSOTgRPrlBWcxEWanIPRw2SbDFq2yavrG
axg/7sLM3mypeP7JAAQnMhtdGEl0Sep4cm49+hISf4x0RG4a4YWUQr5nruT1443+
upCy24EWkmOWPwXDVrDKOUPYjk7iqvxYwGE8Mkp1k7yKS1p/sfc7ms3tR9VT5/to
AmfissywpFkVx1iDuUtE1lzgIalm1s++fzEeKjf0P98rrMeNyU75QaRPilO6iyeS
qRbUJAk3aVF1aw3rio+ZkiyQZk3YYaYIIMey3YSyZjutfNQolTRH21eCx+WrpBQ0
iZvSs7W7MuIq8HkqL1jqgCiet4MTPis/piLy7exKf4mnito0wuxIqOJ40+N5b46t
r1mYaXtnTQNrPhblAmBkXXU6SWlprlAMfN4zCrx/MlnjqpnpieIKtau71KBfBKkv
pfg2U4hAp4f2aYDhi6VAAXYWiAq6E4WdwPvESKJUAzVjRcuWkWDtl3aDFgsCNKxL
vjsjtXTGsr1NJvI26Urt2SiWLrNHIuZHURvWusKVCnvthm1jwKy/Q8UAQzTfUOCn
ZUMIcKZs6pGOVARIiHotW+oJY1Hr091JLGvcUwLrLu/c+YWjdYV4CarWR0EwJigy
9IQ9MdTmeiFaDlLCH36ehjTfc3Mw1JZ6wmyYbQuWIaVf4bGJfOQBY4O4OFVMRTAZ
TJouYCJRPtyL8go/VbWjU1kyO0FPQ6FfdSLf652x/yTbyf6PNPG7uT/SftF8919S
ngQVxARHIZt9L8NsKzAOurMMavmagIWDLenwVRDSUseedCKmJBeUpFNeWt2LoGbU
hgaMxcECXJo0ZzVRi5eqmBk5qM6/fzgsmoAVWRrH3Pc6nS1ueIH5Z+O7AmfHjJAe
WOCBnDPTvzifsnck+/9f1tZJBCCPlMnPbtIV1Y3e8HSKX87qKteGXryLaoZl8sC7
YLYWMsxa7RqitP6KRMjyWs6zj+Btrq1VvFzaQTlPUKIpq2DpMEVN+S9tbTLR3TcH
RjXRAa43lWThAmlWYhV0XRxV9sfMNWkqVtPN6uvl69HoQVxY1GM/xjqF0GRtUA7a
dM132RupwYI3sT0C2iGVInVSmVTnGYmJVj2xZ1cGR2RyR0yDvN6JyrINzAAG41JK
gXdRWXYPINmTTPGrobW2UyDiUeRBva1QCNF16SuuVjGWggXVZ8ve1B6VPXcrQrd9
uce6I7g11b2gkA/IlyPbYyz2toPsnb0A5jpbOGUVN23cDXfvi47B/e0xHpkgXyZ6
RC6oGhKaV/kir/dpadSYWi89aNDUDjoUY74EhXWSS4Ej+yMT+0hsd5DFIOCIhplz
qONF8Fv2cn4QZgFtUewyofi/uDST5wkWTCgfRnPSs6j600apkgF/YGsobThgr4UT
Sxklnbq901CdlkCYTwwDAgGaEpyCsuiUo8aU+YQ9P3sGV3WOT/xK15zySa7Ftubz
/IKxYGtxKGPa/HNdwls33R3DatxgGco9V0ydtt+4qbmfQao95ItOL4UAha/JF9Vu
hCwknZPP8lrYwGisfIx43IB/6O8+7rl5R/WmPg9AUe62ZSK7V+MWAd51f4UKlj5z
0sI++6LNGj9LirXlq0e8WIXBXb30Sx544F0/IC6/Fp3vA703DctEep2xQKMJf/R0
JASxGFiiG0B/PFM+/6o50556gPbJtZdHQMqRm5SOSyS9Ox1+zqgU70uIAlco60/I
UQ+Ouu96PiJ6MWsXFO/H8xo77tXASb79EplFcWovPrbWDF/xDZLyzpsy2rpfnBuf
BByXjm7ZphPSj4Ml18EyaW4rOUgeRbuSHVclEbb0GYun0bX+0GbBzW/i0g28Z2US
LISgdJ8c16pGyUeTH1GvqDpDSPplECEW5YJJWI8VuPWDvsMPxA9Jylnx4kahJ0+L
Ieo7/9d9l4jrhOfXqGH2VbIgoJNgVDQpRrIeTWiR2iIsXvJ3GE0KWAqFd6qCn6p4
keOEZEAbgQKq251bVrZ+V8QEDcuvjLOKGPW3JNbfMsOfAgj4k3f8w261iUZ/Kskp
kgrVBiA/50GYN1qTN3R+y17BFmLzH8cpQiCaV5+1r8UE2zHwyrcqNLg1CTe/0Fhm
sBl4BiV6AkCKM+FoRw7rvoDbWLRMxJZb5dBr3yWmQAOK+OPcTmE0POUHD6yfZPX4
pJJqzV1VI4dZin/PsurLRUZfTcRRxY9HakxJ0SCJ9RWPukwBvy4D+5BZiDEuTSk1
MgQ7aB2BR9q2KIX04bO7kZKUXkM3nu5Y+J/jdZa678cT06V2dXyr+b/zHLVZpE+1
qEXxq5H5W/do4WgZjrBdfVBJ7R1hNBIviTTGFFp090ypQUcbyBAY56c7sGjih9SN
dp/POmDLaIcG6hLiAzWNF69PjCTkHMEH8uyvJ140B1558yDV46J9gkcccP4E1BUd
DKCZH0ysxUiamZayau9xeYnas20dKXRzta6Tr0D03LrGUMYUQySmUDQxqBpC+b7z
CzVcJ6e5FNpLWM2TTWD2IHhJMyqcEe+RtCC3IEvdVI6Z+sqRCEoxY8rPAZVHGNlR
8EHMKgAOGyDViUNn2XLOlc9QHvmgs1wCeej3K6zHrJ49V2OROCqj6VhB77MDJsY0
xbR+6PX/QCvBnFlUYM96a7nq/jP5kUob1r3FEQ6LoNZdJ5ENLS1qrEWoKo3WcWl2
dn+2iHyYf7S8Ss9WwOMcR3/ybA3uZo25xAfwQPk2br1mLq8QY2QcWdspjchaJ7kR
Vp69bma4VENUwoPXN+TP+3sKkSqOvZmVzzA0llGXnGpmnk+js1wYWV1KEJ4Hm/1b
Kgdc81/ER/E4WYgbj4I7B0gtQ2nOnsgPVwH+M6qMPXsH4QknOIG6jPwx0WNeVpSX
KO1igYKBdGrPwKQEPep56DurN3lhvvDr4IgPbaUi/tNvd/aOI33gGeqe/UshYW1C
5rWnfs3qwoaVTPSkYwI/ZViyghVBmN5eWMmxT8WsVL+1LzOwKZrzyoGRWv1QO1aM
WElh/vSJJEqprKjWzR1OunAtPBZBheV7949hvZE/GGPkkvdVhoxvzOVBHJ/pIc7a
MEGxtdFA0Hft3gVe1YG4rN2vFbHyrp+G+mFV1VPT6/U7PyW0ZoWCLRUyZoBijfLB
X28SH947+IzDNMod5MnMdvA1LgGEqWNKUsgpjZKdfvQDkdnMO8z4Mp/EdM9bs2Bd
WT/7RLl7bzKiJ6V40HoHTy+JGg8KrmA6zCIWTc0kF5NMXxR8X6cOoP6vFYltOJX0
KUG1o6Tgq95WWVGYBrS4H+yM8E1XkkXoyQ8izJG3vlyZ8TbfM/lUU5ofV+aCjUhd
9hSIz8ezu9TZKUEwVAgyDvTM2LNNSpq4UquQ2wfZCh1r/b0VDaVxO1EqN0SzcmpI
fnQlRzUB54kOHJ/l47QKN267mA29s4TZLwm7X8iaZvGAimT5rcwZ6ZCvq6iijIih
Czp+zXBqB4QXeN9gfRT4v7mDAZcFp/awWNB52CEnHrd79Wt0BBpCkprsotOiBE+4
vDyAMGHjHNpXnxaC6TdMsoay6e1+GJCJQHY/5PxFDJx2YcQhHaBONRdsabJcqdXZ
HHgakwzPz4OgCaqio/lQt0Xyh9NUQuBNr2oKFWMR0TduokLpvzx1YNUUmR6f8Kpz
HTQvp4qBI8OHHEl2MqJufhpYXLWmD2r+QpU9yCDHBLRUZLBOoFsyIWplMD4RYQhU
US6yFbxGouyp5tsjebwXAOS6s++w6ReSmM64EuMlZF2jcIoctvh7Q7m14Xca/anr
RxIS3RL08kOU7PlW8hlqUsAWzplmAmalms5Jo+cVzL4B0wG9aGuqgLEhtZZlZRRX
kjzCeBqle2pHNS/EXL9aneFHGwuKUTZGxti7OA1on/59V2nsAb/T1fYFIxLgGHMx
vMYFOPkS9eLf2diD7FqR6d8AxQDjcMwYiMsETXDXERTMYaYATQvvhNgetV2kYbox
5OzMxizpFsHQgfOmJ9G9AOS489DFV2RC2OCndTsIZvplpCDjx6AexHI0VkrKLV0f
F0wDQNzQ/ucj3BgA49KcptEw5H2E1kPuzv5KBrIrrIv76qwyRE6lkjQjPkjngeuU
xrzSUolCYy5xBERJW0GHm/OnfDoiEa1gLXxEbFQRezRm+vdSyL3Tu4Yew3WZbcfZ
fsebqYrwaYvkFhuAB5oi5z9vx5o6HEMyXQ6cdeTVGoSkJqBaPynXyn44EjspPMiV
BKt/uKuz8w8aYXisoeb1FiPXe7xs8klcG5zdmNQcFWAEB/QcMjaBQSHz8vEASpxJ
8Zq86kI0Eu5HrE36lJaSJVJNGOyqMYMzAAk3PXr3sjgWOofpL0ZsZigFfPqNkJdi
rjA6hD+xCS7qgsOc88X5mC15KCjEWfA8NKXEKmzBxjYkek6QDtDCXOSQutKifMP5
N06//1a4b2iRdU3aQLxXzWaHsnJ14cJMFuTb0Qkr/Xb0Ii6s0RkLqdGibxhRNlqA
oyYfVMqegi7cMH02jHhVQqpmS14iym8lXICHYtMai3MLzpgPkxyppPAleVEvOl3o
I4aYMelsMsT4zhEN/RluQiq3BzDhQ54+aYoScs8mrhMw0yNw30/nKs0d5H1Tsd6i
AXOjm4/bsOmGrGHv/0zNzZj0w5Ghn4LHdeOUmHf9gx20AHBScJ+TbRkCxt7T+ofs
H7qlbGktnjYV5W71U6rIhX94dHHkvlzY72nh+yhv1kDHBUBP8Msi8KUZmX5uAQAM
4ttHKx60A9AjWKhgrub14oBZPVCUzMmMPwED/aIdiJocqvCpuKVMWlhZ2hwkG9cJ
9Z/IKpvIN/iuDe9SO69JUBIkFcwm1crPUqavldtvX73gmO5xrMdWiQSwras6GB4R
JK9CdTla8uhIVb0asZ9Tn9/LuUjT0tG7vCzgjMI15NXt8xg7+/6Ngd3df+BhoxVI
NN9RRF7bQr4o0phEfeShlIAwVOCEhcYrcWaVHTEvCsY6SPCShB6G5QKmoquZyEFH
y/0Lr+j406PkpU4LGii2gYZpbl+YfvWBOTwuK0Xr+jyY5p3ABhuuXArWClfXjcWT
JYSzT4q12ETaM6kB+83N3rpzuJJ8xX/9ADFXeI7HZnkEo0cUescx0yTEtzm6sA3c
rfvwVFv8KerC162qt7snC5DSLqGyf/HZo9Vr3ftzBc4IrBoUqnnlpOGRMOEAppvn
3JUhBw7JcZleoiOGHjMcPyQNYNgyh0K3RLsGBNRzFSDvPmFyST2OgAsHFD2aHocY
PuZ+8Yr1PC6wW5KyvvaGkkpLwZiV92O8tf4JrY2GFHUQLvF906gY9FVDQHv8EWiG
PrVrzwF/k2vvrYhSBed2CiozIrljORRVP+l3cII7/oPZRW+yIYLubEZJNw6peUDa
85c6h3vTY3lIDik3ZBs4Yhe3cezX3gYJUK5IUpoSItEyd8iDE8gKNn4jcOk8gmj2
meA/KBW0cyJBykwFFQxus19OxkMGYgVCKM5tAu0OUgmcD1o5iv/L89moc0Tqvyhu
0fLqsF2W37FPsy2uyST99TGVCQWGqwUuoWBumge+ZSzBQf9p9mR8z6Y6J8O2rnPl
45yD53dR8HnJ93yheHRfuAKO1rLxYGXkX81HGmzhf4JQifgTKVrCU8U8XDc0nMRO
5PYtH/OF7uT7ty7NEeYbFHifs/G0Cis1T1FLXOmywRUU0Ov++PonREEPTwndyApz
UayPXGflz5ixr30r9emU/WKwcSj5HM9LTvkfQ9/zRIvgoOGYsLc8CO0PREHDP7Jd
ViJAsOymyt36VHLoU4ixThSDGcdVAYnmkdNmGzOPW7Wp/Gf68NbcpZVKvgBl78g5
W+UooixvJkdF8tSX/b32/naUAT8h1rXV6c1hM0/kjWeqcGB1wt6vzeu7fShgKfeS
nBUmgUusRYQtVvmzKJzXTnEySqREGl6RqtLN2/FMsY3F84VPQa9hdhs1Ec8V+Mxd
DkP7DwyCxMVapUfGFY0tz1OOi/RAQZQ5W0qby0YGrOw9ZDPK6ZTws5C5glJj1w2K
ccK5XXrjLhsccEqLDQ3pmhLtnaCTOi+qGojA3JcbqLZjZEyA+x/zDyvL65T9SVBK
ezRA1paZzu+oVg/YfGvWNrhZILiE67EV40Z8ojip9Nj+bDhK+pt4OrEg+ynIccZB
dIjnTNzD9hby2uaNNbEBL6AU6u2JktVqpwjmz1icA1FNE0MvlQqmTdhY3gLqPuOy
Ijk2VoUvWjBnJBRlFhU0hAM1yj1m7Zl9YbQL302jy0qNC48IOoa+HESG2ifsmyxq
caBWMY5u3odQlQ20yMWhiGj4vYFmMWm7JxsNc7OClnYZqAtopIb6d7L0puSrlJQl
nFjhYOkxw+LXpgAnTUPiAN3GWpQ+M3hIufNAOUsC+Xsq7nac5Rcx0arR6MZKj2uj
0AC+PrIiiKEGm0HqwuZ67PesKfclLbIe6+Ji63qe/8dflBx9hCDa9V/Er9Ocpbkp
IgcIkQxjP8SNBrZqHywPR2Db8sa+xNG+17YJqQr/hHyHmcZ6v6Xc9+Lcju8dxZSh
JLLK1pDXX9ii7wTjYzGubzXvboQCv9t6VDENFFen7GKP7Dnpdx/tl6VLzBuGcJdC
QcMIEQKdO+JOGJN1seNHget+6KAxcIMK9AIlJYwKo5XNQrl4elEGhVimONvCIkCq
ER5ZUFXBTnxhJqkkPJvVCSKTpFyHiVbnLx4G4hRGeQlzGzDPGQr7GMvOARiYQzCt
ubVRZw7hOqCVQLH0IpT0PC7cfny/2xI+iKrpiYF2o/s7CImHCmgT6CtoHe4Lt7JG
kIjI87GoTuzqq3vhXN1AXOhnZ4ZH53ip467A6iViSqF/oJ4j/2P3YQdg/NcDwHZW
/cp9CJfAnwSwlVjlmw6iXcfbudoJ/DNHpBV9vk6OF9Q=
`pragma protect end_protected
