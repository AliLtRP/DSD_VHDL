// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:50 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
rMDjPDBoKp79MRv+y92AKSKx+l9ZTUbjMq/DjHm1yy+TBIVABT5/oMWDXH2glFxB
atripY0VAcYeQWlpokH5rhovdqYJcjlAypuVRadXBh4eqtuXTDosFmQcgbrJ/2z2
cFz+Rjatk16QJwStiyPJGzs4zuNsfXu5RSsyJwqKH18=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 29040)
l+6NpQ3pYI2SzBXKcjCK5I1Kx9LDcDLfQCCri4tMsAXVjV0YxenHfpGC7cVliTy+
AE78eekWFD4M4kh7PfcxDfrEB63KVWrFuOzWnUHr/9QMWxlKjlDnjkbrvzomSCeO
5+DVYwP5WpL4OKuLFA86E/Y3l3NW91HADsERPeElU0nfL8N/erOOQqVz6i6saHbg
nuA/2bQE2QyCnCzN6QvdcvQZK3CU/Qk0FTppO6tehOw4z8Si95IToVPqAy5dhNnE
L0VmSmcW26bzRv8iB1b2w4BVuYcI/d/pOsAlxs2DpnNoGcEahclgtXjxzxpMlPR0
iGk2lS+Q5S3yakTtuDgNlacehAORf0ocQ8Zk9AicAC2CTJYvQ7SwQX6DT6MFfO5k
0JNa+1QRHmIFqK4Xxv/bQXzW4ehx212IphF6lIq2HoGi0Qt4xLjIVWlfGaUAJqWr
Zz5k9bGbCEKDi1vSrlSC6HyRX4R7agQ1dyxOhERzDtAogza5UtjYn4LQ34lQLAmp
+XpbACVXIvfGM+7m0H1b45IJDhjvBgpaqZbICLnYyiC8fIoYJnh20QMUfQXyTpoZ
fF3zLiJG5r/OOlAkpgIj2NJCyM+aFlSfvH0J0sllC7q/z9m9YQte27oYk6es33UA
hKnu/KA9+u/geYQJOANAv/HkJUaOzPEvnZf25Xjb6EEqf5XTjShHwy4phfXkLp4H
3oUNvOORGsl0uTGnHOm0fMKOpkVQhPiDErFOf6apsJxBlN2JwtnuUJM85ZYuOT9m
qDobswjhQ7aRkJ+027xJgzYMHrNBLHMg5PbJqKfhl03oED8Hp1bnQjSdRKSfElQG
YUC2NVoG3SDw3ish7LbNPFQo4Q94T1b67/frN1lBlGPMX81aDmv/jwXL3hhqgRTR
t/0S3O4Pb5yn6BkgZycB7gf484v/o3hTTkCmV/B0AHKEPMfwnVsXItqkp2EG9M+9
TQ6CovwG01O18dXLmaoWjqD2OuOfpH1hUuBBeW1SgAK0qHQPqLyg4F2T9MQk3B9z
cGW8iDTte7KpVOK8GugkOUoP1WESHUYAGFywhp3kEbyWXOQAXFJOJGzdKAkbsshS
KFSk1rU3UhaUsLWpIC+WHziwLaNkOg7D+wJtPEwraCyIWFvvK1D4HSLrgVIaqcxe
k4fFBaHfQx1O7ZwSP1XRKCA7XVGEsqVEh2dLYQ7hIHeIAdMZ8JquMoq7lydynwIF
g+ZMFRyEYl69fK6ojg1hA2Kibnk3gshPnBc6qCDSeM9rEzMUw13J+JJsVXXYjXhN
Sjv58uik4lzj0vNDy8F/cIysvqdgxALZmTsMiAp22OpmxGLfAqbsyY8+WpC7wZYr
TOm9VsFw+MIXRml/jPIDvsR+l7hNJTCpV6nhSniiUQd5z4tCNNSNvhmq0neFs/n7
BaZ7d+DMllM9C+lU1TjP1bOkzNgfnbpv2r8bwOtXWG92lH5oY8xAzf19277Cx+N1
WJNar1AEuPNIH/tkVux/ZbtFRQR5TPoAll1TZCxooe9B0tAx0rU+icWOFzZiVlaA
XsVBjex36GHBs1Pkw3W7qeQmggBxOdWdEdlfp8ON/k8KIHcEMkN7eV1xxcfxj4nK
Djf8BXNvw3xH10q8YMhyhUlyKGU9bI4A6oGIf4RttXT0fWVdWBqp9xRD0SbEa8NU
Nowic/1xQoqZlh03d6EwvEDdNDvncfEiboOIbwnix0RanYqXw4y6B4xPXt+4dEtw
XaNAyH2gNulwe56xPawNfp++kvAuhLjAUOJPniaINMQPAp1n6RhPwbtf7b117Ld0
Rtwef3Q358twOZhFTtAUxAD0dnrCDuc55p6nfGR0Qb0ZTueHVsFV47ZRJV/mdDfg
LjURyevvHUTC6etFjos7r+rH5gqIlXyqdIlp/wk8SEuXgGxECmiO4paVO9c0kd3R
fn/lhtWZoKmUSlM7KHql53rKOCEnd9N9boBz/I40mxBsJmy7s0CtHPtwf60jKvjN
qZEudw6gbIJKkJ8ooxyC8lcQ+ynx9aRZYxdHV5vdLBfu5RXPSH/hT6sOZ+/b9M9I
keYH8iLo+/oLOrSCJfqYnXwVmocaFTTooW/P0dbHHIwKqq+U5Ihc3pBgmj21R0JX
/si5RjheiqnqsjofQI9m3XU3ecYAuW9uiivWyH7S/y1LYp5ujzsBwq43yfZINBhX
0t5W/ilrmg5NKDN/GsS50HlMQwzfiebBgXsWN6N2eMDsJmBHLwX3Oq+voZM6PzGa
SJ2LCvn+AXh4jwCjYmb86bWT7SwGamZ6BIggGgLxHXHh0+KgnWqzFJ+V+b4RnAxh
Ju/3NVmff6w6NF+BhjQ7wQC9qpy2T00BHuoXjVP2AXvkiSMEXFNscWkcjW/THkA6
OguveV4MoayLlo8WDnVy/m1B+LuP77bcyHL+f30ejyx70o3fQpQbaq3vLePY6FV7
GYsQ2e5138l7NOwszwHQiKF1DHfJa4blL2lnwto9Ygti5SnhSuTBrmVgvPmIf70u
hHcHj+iSpnk1uVIgSCRjJwW46T55yMafxr6Q0YkXGKDahLb8m+aMOMJ1r0UfpAiq
/a+kBfeuqNziqmXAG3m53p3XbXNF8hqi0TbVRiWygMdFSpudFlSRdYHNn3gTGEQz
44FIBr8/MP1zaM4MvSyeX7jajRV+svGAF/wGKtSL0zmUfhPpl9jZpvjbkSKOTvx1
Fxe5Kf9639VOLZzj1WV4wM+82e6nJQVDbdjpctoCo61PB0gUz4Egv2nFKme7zq1F
oTixA8jpLkxuzsZTEHWqrtndO9Bn4nEY74zjP1ujW9c1GZDjGYko/jhqC61IkJdn
VNiu1tIULMJfeFueuWJSBNAH+u9kJ5PD3+a9DkseOje9v9x3f40DxGYJASmNccMY
ds/kmUYbvC0DSYZ9ld4b8pKEtaz6XuBUduzPWPdbhiLE3HPMtBXcY/kR39Dw+Viq
IT8JyMyUPVAocHc17zH4ydEuZXCJsH9hDojoZQ3taZXc696pdRql2HEEUOHPNBnh
edd6vS7K0tGk00ofgyo2zBwXbat/dOHhY8PKO+GUnuJKAgGT1WmLlTBrYDnAzDRR
Ck2HKnmevEZ1Ox2r8+YU0YYuIpBHwmuk8bJ/e32MD2ErlmKsOnvXNorlRl7aN+Zc
pFmAn/OsamTY2WdAcAnvqregmyKoHyF5id87EJpnlcacgYaRFVVKK1yGmTalNjIA
IL3Y+UVo/VXasxQaWAvY4OGTMdJPB/YYHvM4xANUjohQ5qcA/E5AY9saYc/72Iub
5cecVu9juU/jjbxzcSQHThZL2+JISnwe3E32wp93YWObHl8aBeFNXCYOe0GqN1zs
PsUHAG9ycoipjirBsmpfaNL+kXWENXCA75LDa811Ou1ae6zTmvuRWqMbUABxQgsI
s3zAtjKL/MGKYGP0XzdPxUxMeE8NAuuq+PEeqV3+HVYhPgMtR0PEXxXr+bRZaiu9
hUrXKXDhBcJP3OaNa87KT9oJe8ceI3PChNREA2Z9ITIBDD2ZIBitKXELKRgQbemF
4cMh/vvcFs3N9rEOZNvPWOMU91s59b6ZBmqwf48nI5GnR1ig7tPtEHvWsEQ217AZ
B6/Q5k3spgE3IESNUvJIM8mlT76WqrtYvXc3SbiCMNNWbiUyOT57K3qxJViRLhPO
W4l7OIKP8xqtc7BbWOzvs3EuSUXdEZCYaUu2zL9zV+aHLJGFyo4G4D8c/Ftwocs5
myUXMt2VoFvDfL3EN+Xt+R+nmGaH3JClhg4KxdJZK/hnGQYZeKdoEXPh1yjxGoC9
3Bwg+c4QrvbhQMXp6c26d/x57vrPOGoSbm5Ia3Uv22vnFjg3/6NgEzxb8/VjJXZp
g4hbFWiNav7A9prW3hLoBq9kG2KPtp+8jaQKYaCvtTYozm1SY0fUfRgV7oLFD4vM
occI+Rt2NmUZWSQ3FVtiQIKlDi+7fBNbVAVNWMkqG/N1hbcxhrvIWGYUlMEJbTXe
jghRRAfFujlMvBPoIA59Wu25H0qw/mLIr+seNK6tE1WCGP4Pqwh7MmxXtYpLYPSA
695aIHP7Qy9SgzoPlf4s7npWEz4cx6i7GbhqcALqt/ZP0lA2AbNrpGKYajtrPBlA
sexevd2ORtmDOvLaNpuCl+MjQwbnCFSDleJUAA5r6GsJZQpakFgPcEBdoW9PTra1
8TYndXXx2vN+9T3+AkUllKXhJi4TFnM2zkUz7i96HkNxrJL0LmtBXqge+APyq/cY
NCmRLHwuiqs9vwDupDDn1Id50bh/t8KWm5OPoWaDtaEj9Erp1eLJXfI7DYPAUVn0
Px5TII9XTR7vbdFt+wyESbq27cIcCw+OPezk4QIozhKgv3Iz2MSr8ruYZN9kYtq7
yJqzVVa+nrBmoAVaxM5ojo6LjleXDbi+7S3F4rrz0cud0a1TgSQPFNTmQvtblo/B
FoSrHwl+zL3xfh7ctrBaRcNiROpaCJ/OB8UuCA/S22LZgDNeEyP9c9u5Dc2HBchr
0C3rdbkew3OVwC8wXXy15glySQZ90/GYQHHZAyELpKDEHMODz149JJSPECPXmdxc
DTaSIO7HssDgyBDI2FLc+OArqiFICC4tUFdHGkgLJIkvtra1p2pH0rfR+t2MHIPq
PjHLnorFBOp8gG8I6RA4wxc0zHLEKX5+NR7XI4TzEjgD+qO/cheHc9a4QRM1qDNo
QSDpIXIcr/C9A9vNEEfPYcXDqT8saut1i3/+SoF/C2EPXp32o3c/VzXIJiKLOVDo
/u25LK+6vNGydPhFdaO9i0/0q0hzTltbQ/V7n+y2ys3w2DorBuW9aTgfmhBe0vO4
VjllLAf3WW87lgsmO889wyrzkGGMeHj17GWqNBoeEPii1af5QU6cq9G3ufJ+tZNZ
orvajkROj2d/6IlbdtjzTmvi2uHcriBSS24wTOlYocLLRuhqJVjS6RfSlIkb+YZN
1lsxyiX5cNAfaC/4CUjl8BuqjkFrPdDxAIwXEjSdPHOz5lieVvFJt4+ybidnRJNf
A2b4EBCS3O6ZdxPDNy41zSUtatk//xSDJvtp688F3lf5WsCoz79YJupAEDUmSttP
4eq/DJCWe3asAGT52axgtuEQZTrdLecs/EMn/RyPBHxZw5Uh1q8KQj0jJSx0lJuP
l8MnQDCJ9OetHQpuVS0lkiWVoCZOWijijo2NzVxLRSaqGulyywmqPFHywYmsFY4Q
dhHeJvZUuMZWS5ewz1cwkAag0Uvd8GNeNDrq20RKiX9uODMsXxhV0f9guEmrcdgK
PJMTDBGxZMIX50yJVtncG1aXBsrhEOPlR4apMIdFaEHO99zYOsT/3w1crCZfIP0M
mZfX9Odgx0Chs4mHeDvf5L01kZn+LUr+UYFPTckyb/c2GWzqSkfWSLwz3YHKLEAg
f4YOrFhY4Px6nxkrAVRYZD4uELE0fEuIUWPI7KzQZyFpcOXUQLQcsu7Iu4izsn+y
y2Gw/qFZKNSE33lVZuyD6gFND47L4VK6qLSv35QRxavQ89CnN+dciCfzpK/QmAgh
CPQYPoOkT3hw+JJlfR0zv8Li5GOpYTdVcjf6dc9x4xX0EsLXvVUcVsNgHY8pQENs
CKHOhWS8zOAgfVf7s8f/xfa6//OlD1o+eM+KGWDskxhQZV1jJZJgb369XewWur6f
/Q0Hx/vtaMmXs9mr1sIuz3B6zVGgkCdmq005w6PGL5i32xgMoq4spS8IZjcfMYKm
CTgVRXae6up/ddJiweI4Mba8i+E0+snk87yx6SrRIrZqrXArEdLhnaXvHx3pTags
/av+SBT/uzexp0sfozIHMCFFpfuuprJN7IbqFXfA2D27v6BmmcNQyW8MLdLG5vaN
N+KxFt2oHZxIQqJDTiI0CW1ahGlBJO4VCQdjpENQXZ+pT3MWwj6AKTl2AHZ8XpVy
8z02tVM5duhw9H0dnUObra/vMg/wcVC+90ucovY6M9NtDMJ321ml7nleSd+5n74Y
0mnqWVcuRyuFQjJVlRWSxxDn7owIaH6A+HiZrhahoQBwiuRspcKvizYuD8MW30ec
WgUBBNGqtdyAq9RRD1mf094lAfUyk3PRirKMQshIx32WLYog1d3ayXTRXsZD7fkO
UDODVgTHCwDJDL227ZwP8VQ55aKhBaiqh9Ue1eW+8LyYQxmP4khPOnAFl8FhAUQS
GrCftUQY6e+vEFJwHtlurH0u/n+OTqIS9W4WyYFJsLUDJh0kt2PpvDmPXEqZ7RJ3
wWbmrLNA4ymv5omJdiX0It8Q6nyDWRx1FoSLRPMAlEG7Z/chOv6Xu/ZillAYjTIL
hMSTOseZJnRHKiqrylkj3zb6mWusGfgdOE2M+j/g6BFtx8o1yPU6z5w26tc+gLCl
2EUbPPG1Bufzo7OTYySK+uEWpTfcU+j8CudohJGq2/PQ1PdBgyd1q8vURbK8XBAT
T90SaC5C6znuwgt54Z5dpdkrLlZmyL0nU4uz8J2+QqwXmyrpL4HE9JyySCiTneYx
5HcAahES8/AJUDdudI6XSMCuGzXOgXu+LWsyfCjrWLo2GREKAX9hLAMoNKDzMMGS
bG1HKSj4eKuF3dA9wGpexJVULcmWSdu3C1jimSFqRLuZch5Bt9WYjTXcll1OuuHx
GDGFCyHOhgbagNQnulgJ+TVle7F3Uop+dHVbfNuJQq4HkOX+J4luAJ/4aQfZPdBv
i7tqSstMLCxpU4gN6g6sOc+ROBQqQ/iqqXz7G/k6c05OUuEGwrmTsIS5h6qvGige
1Ep0PpuQsbCN1w6tGRpNhpmypf8eSZsE/jolpktPVL3sc8l3r4jQ+IO/soCat76H
kxvj1LRVjziBvdEHMvWsUGUGjxhnUnMHie5i1I1WLrAeU+9RoecmucKnyXgxHsXC
Sx4H27zBqhldRDo/qUaYiUUicC/E0XcF0vIAhpljTCsU6i32NgW5C8IDJfHP9dAS
ncCNATdgEUNdByUifCz77o3Bak8cI84koWqSCnqecoV74V2kGTfZ+HMraOi3zFFA
B4AZol9o/2VNli0aiExRIMCzrwvQqpBlUFxXXzT0WMPQY7siKs78VzmBse6SfzjF
ETHwlz25Uez2XwhjsIyeQ+dNi+zNGk1UjqNQNeiMGbu1ylSydqJkI/4orcn9tupn
pbdSaQTuZIdZ/a2OpemCoaG3KgXTqxeikwAPCnwVY0bf/pU86RgzMSwv8Wft5xjR
ZzQoOyWmW44gFgOdoOkv0bc0azEPCYA3TMaNmTKSIO732l0BGdHmJNwnEePk/qKH
bFl9JWKTAewY4Ygem/obe72bMshZsrY9Oo/mrGuEGO6Re332Zh3UtDGIipmwzX/j
wlTPh6qEATf0TNQ7nHIroxakSCD+NncuuNa/AttAtiXeXhwRAq3lkbeb1MCcttDa
sLHj7YlDHKPHMzL1kTGss/c4FO/tAkxaZIqWqK29U4q0mWbND2n50d4865wu6eY0
xXuuEdt4kM7mPhsIPq6Gv+AWjXb/LbhkT/X4kQfCfw2paQmWQlxFsDjkC4x6Ah6I
qZsN4pb1FBxe6C2YWkQqnhl9PVRUvmmmx8OBGr2LEf2/boLKvL5p7Sa+h9buKOQt
OXqHO01k8VXOZOSVsnXSJ9qthlUScBbHNQkYxTI8y2syQd6Z8SxAXgB5t1+/ZO5n
Ncu2lN0KA7WEyog401Gf34RBlBNI53l7pz2oDpXHStVn81Kr3gSJTkWhTCOUVJy/
v4XVvg6PUNfHHd+1D8u9CSuzvpl7NQpmUrfdcAkMFx59iyT9gROWha00IMGOH1U+
SYCzfvm32211jI157mpB9WebYRA0fzKmv3h/Pq+EKAAPJKoX5fwz0ZZITqsQmtRW
HsnF3wfRi5mbBfdbMVt31sGIEl/zcFgOMe3cfXApgC2MPJtU7hh3W350+lRbtpuX
24W6lZI60/vNkOO0CePgXFdWsyeLeQY+8xBb5nMxo0Z3JSMwKcf6ImJ3EAWkyM+Q
HxBlHmGHl9/fipt9QuahwfIqg02rYsZzZhTjKjKSQbrdHTd1vkmdrWWxeunGPrD0
bAm62wbhbb2Vs/9P9a57YTj5q096YKrGnqgeR9ZxaIKHnuBhgWfX828hk4xvhY/D
xVKjOFvnDFfgKZsFARD0Br8EVm7aVdreCTT23IpWKqW60+egdlEL8WzUBALZZwue
ZOy+kYoH554ptt0mRHnHfIz3+uLiftfs+Aq30wbShP5zBSeqSuKMkQD1ss1MFc5X
DifiXwfY6VJqle6KYYxX4GfyInGICyzGq7ukBVRagNxAdbDCwHw+WM0guzhCg4Kx
SDqP5G3z23Fd20XnWh1ycP50ZJGgRvIdGAGUYgXDoFs/cAEca9nw1sULhPLz9yZH
HqtOGBEYdv4Sd62SPdtQpkC0imlgoofR7GnY6cMyLgkbeC2waBPPfJdFdPQ1f7fr
pXmUjvCxyWOkpGOIATpnC9KLQPlNwJPTVRbDxFauPSRGp6OQO+GX+ZOoot3vp/e+
TSSZcnYVvDJAiXTqWnm6jS5M49bXrFXF5SUpGPcKNEa9bQGEcGrt3y3425PaP59h
SfTAztHndxFd72tcV08trqjW7yqrpRTa0JaQ7mB+NqgrZ0VpwBZFr/bkuU+SOyZ7
i4XJPyOatS5dy/DPQ1aKGgP4/AFZNePbyFyNZHiYa/3706ye1T1YaOvNOVOioBZq
fdo14mm7TDgQf0yhR9HHy7y4PhpedLYtuxExOm42oWobDrMHRXt2SFsM1ew/7TaY
MkL9Uszh+QEnDxRllXlefObEzH5cI67FTJiXgg07HuCrgrZcraxIx4uJVIhAHLwN
ziyDmN9OkW2lvE7M0GRxMoWirB/sLbJA9A/4tE+Il9gZX189YDIAUtQ5nmkG7M8O
CYHxGJW54t2WAtZK2m1iSLzEIbymDnYab/ysib3YI0fn6QsAdZRJOCIRvaA67g6J
wWV1lMF3ZOaNR0udGBCguOIxTlA2c7DXwAqT4EH1JyemdQ4w87S/TvhVrkm594oZ
HzUgapNycZ9whNYT4dL5XBVkZc3uFffGKbjxaZCd0jxa1PbKUYg9ekodQnh+RFIq
ZRr4WlCjhG/pNPCKVqqjFa6zsci8VZe/EMHLq2FvJRCt5GTd63xZcT82BtMP6oiM
/Va2cGPAobYW3HxzgDOvh9XVbxX/bqlV8oZprnC8mh6kJhF+LUcF+nqbPgpU10Xl
rZAHT7rsE52TLeKe3VaqxRBDOz9MAV7hOFdrTLk1RkLxMLxdBW56SjxIo2EWicf9
3BUJQmPOkjHRCsDZ2URdtNWQQyzDQNRCAqqudrUHQ5meNuv1h8kMyKRUHaFpmmHo
eVlvT87Omdc3iS/XINKaSo2B4eDXUIrt8HXgb7hx9oN6oaJqxxqB+wVQUf0TqOx4
KI90NK7lvyU8cz7iBcjjwDRIgk6kMx3qhWJurCFsPOY7Cj9PPKYHFgD1rjl53HhQ
b8SuvS+JJqp0hvYoqL18OXhgtm72aP7f8XUvDhIDlrJpZsBz7sQ3uWK4twQ56DUO
a39ZnrEJ9ZVyrDhtNJfRpjlKQ319VWyNMjDd5jD6f3F5GhjP67lGqNEtOQOevHVx
uIkaFrZiOZ5Q05LIagZoANBEylCg14K8UDeHBlouLumXJbVyUGDjzFSLNahCNCV3
VSNNoily6JiSDeijmFreOTGQZoaynWSX0xsDgIeq4VzYJZCJ83nG2N2RXE2S3mDc
WnzKN68NAx1nhBJx/6OGSLn6MTpVONSBJsQII0hNCSD0v1ApN75RdcpcHUVYukrN
loWG2CFj5jlbOcT8CAMkEPzwvN24FM4netirQdXTLg877c8KRjpluYeRiH1Y30tU
wizDQhlzZ9CeINwMwVqnkf8qZcZIShVrhlGzzgOtxfViZiWYX8Yq1+nFgoXFfaZe
qk5nC1aMO8ZeJmBDGeB9S2K9VEcmSOqTj6oXKGNGSK7IGT7B+5ZHMlH+77rDmejr
XMCl6v44WBlBX1NHFy5n7EVH6FPdWtic9zK2WmIEzx7bWRw78AaDVeYZHg5zObt7
j3nZC1Eu9CNc/gIzHLhGtcu2F6ZLKXd7zNFSLylqFs6BEdzXEErU9amxuGrI0yp8
eevN/F8PxbR45mc9iS3ixlAus4rVm6EF8aRxaOjBV7raqwEexCx8udh9/qIPqQn9
7OwFnxvY4qPWvCLpJ9H0zhBbrvf4qj3PIzB3Tuez5+BEG5Q7ND0ee03pjQXrFWLF
/D3NMabPh5k9Sh5614WBb11HyKvTEbucazer9WpHByMHYb65Zn3US1HM+N0BjE0c
o/JF1rkZLmdFqTkmnP3+7mBv8ql6PDmvCCYRrROjyUmEacnY0zL5AKREENdebmJ/
UzpwTEhEePiiywtyerotCuoTeGC6KRJbUoZgAj8PXF9TLwBHit9GMr4etmJj0kG0
fUcXCrHxynczWCGClp6fM7mRFeZqCs0OwL0h9UdOY+4+mBs6hdVbIcf2C/NPwwMj
gbhlj/jhqY1AgWJfQSFutGRG+5HwfT2SFVU2dZEoQq0yfQyTZU3cu0eCTr6Wu7Rn
wNBR4KzbWBzQq1uSslEJIJr+2pSXjiDrlgJWBFEPRbLyjfugkmrkw+Co2hblrv8E
83i0OtJhmh+hazeIhtyXBdzXa8CqNv3AjwUJu/0xJDI1VfS2D0uWXRjsYbAxG0Be
E1wIsIVdRX/aH/gPqjkPUTVIL/8qCAp8AJokIqtWg1QIihfV1JQrnv2plPc3hCld
3uN/RiJBlJmqXyhlWC2o3fZ9obvPJG+zujDW632K1HAC0qgCqJ9XUEhWeAf8zCtx
v4A9x9da7nNye6g8H64ox/CTrMDl9h1o9K3XxIpU3/jgu0KeRG6Gcpmw6967+CjL
lP0WX4bBsuUikdmDGTKqYIYRWtwVbN9gQgl+Zpw8zrA8LazhqOJYzof2H7Y65JwR
uk4ilBUbJzPKZlTAdCWMNt94btkiVWQJSmPTYkxtnlLBxMfmDgJ2c51XxQTxeMKe
fFAxCV8ThCVnQuUXDXikIleLvdSBl3QONN4g7SakyPojsstxi//KKgVGHhpOWfsf
Jo1G7EsvV6ExDn+Nv7uAw0EkwXsv9qxUce3LO/1FZeUru2Wy9GAOIIA7BYs/retY
/MirlBQrAWzWthdYM9SBtSLgSzj5/Dwd9LX9zOPscMdp1J8v5GCo/z8dNSNeV0Zl
TRnV/VzjK9iXNEYxjULSkU2w9D72k5CBs8xOUbEMKRzDTyL0U5XqgZZpVgA/J9cH
ie1SXZ7tkUlRc790z6y94YlT5jGxz6TnYgBTwdnim9dC5sxFjQ1swdQffSeMzcOB
fIhnnczPpBY8tez1cmr4xpAgUas1VQtD1iFGdhRIuzi/gnqsTVd1lx1kei7O3SNr
2jgMAV+28Qmu+dXsmbaTudH98qnyciwvj6MhLsw/TcnFkwS6Mamc9JQD65Ur8W42
bg7hRRMJjAPc8hiDJcK+8x1iwt690v8f7pAe/q+SzAYdVCXoE+Dhllc+8+3DrSQp
2p6lhdpn8rSmJ2J6W7ADkSsnKBQn9b61gg5f81boo8VmjHErvVQzcEQc/6X82wmS
1hu/SW+UZHsZMqslBSAnRLBh+ZeYlxbh7PjYRUiFfO5gKth9aI0xhI0peW18ovIg
+TrT3qOz9VgDmvaTnjt32oBuKqOuB6cv4NuP/aVNqMJWudkEN9nh6SI8IbWEFUXX
AnLIB4zaVvTW4L6PSWNr5QiIeUKcEWZOdoz/RDBLkR6s0upO9Z7jCiBxBnNxz3JE
d8ro+10cCO/MFKxIKA6g1reiwxmXuC2BVQAaGw/jQ/uxS3tPq3bXoYRawZoQOCLx
v+CR/m+vkgnvuJBS50DGx2FLkO49YSjARL4kZ+dHdCuuv+RIyL8JRw3I9RfVxAsJ
15f21TJhV+lcnJ+GBIQJTv2Ktn54OixSOU3RQLiDzKgnsVI+IRgiqUFXEES/Db8J
D4w2YXefC2iBq00wAuSppbn6sfGjCZmENrztWVGa/S7U4kQJYsl/NeowuSuaBGL5
mFW7Ly4eFMLtBFP+bJd7a/1J1VC7yS24sBynYWsRGuvJGR70djZ/WRbd1DasLEho
1HjvscaXf3zj8JG+ZFiMd0Usv/IuyZKjdzVqMFqHT69QJ+SkoV9RK0AjbG2xYxnv
EqM5+KtStozt8Po7jNh0egFVXGlMVrTK+CRMTCxwP1B5N0ikBd25gCm7mPz59dBf
UBl6luKpVKHIW075+a6nDePUEuFPFXISw4rang4RmiY+WhLr4rCwL/7Kh1FbuqKx
7N72QpUVfHDzQPcbPGoSC46PpngN672/j4nOyZdsC19Hb+tpzGs14KFZj84Jc19y
RKJITGPYkZ6yCIJP/nQPqYwvXV9XYZnJIo1faru5Qpw1hjNAGMblFLUeNvEOeWAJ
JNopNulnWQauvfz/Y4Wo1eHfaBqA42BEuy8utdIBbcWlqu5iHTMf6E5KJ2JMEUyp
y7JEjUzN2hzSCQ3mrChonXDQipDhnDV5TGF7QQ4ogKnd/w/kiOa/T6DgKbaMH+XT
jmvJn0vPDd38pnlQlFoE/eFbI+CT/0W3eCpRHWg6tEuxo8f35Sk2lz7uirnZMqSW
fyAnxOE0S130PqHu/dy9tASsoH/ynhw93w8Z2Ufpwt5XFLVog9uxpURqFsGjvY9Q
jU6uOrk1FmUucpfHCgbU6xLcxxfMikiYvEXF9PVGtD4iGtUl1f+Jxyx+K1gRfw5M
OKTpq6Com8h+iWF/rVY5eN2o5M82t+bxkXjv9LhRXtHdMPnpA5urSTbZihL492iy
pyGVhBpydXk6E7MV6GhOBAD6yyOUCEgIlgyalCA18afFnYM/cZsuIfPFOp5jBlhx
tvd6gS6/dOQ+WCsOII8zQAEfwTGBC8bh+blhNcpYvpY9mKm2F4UVavlpAGVOOAD5
7HTueLmUx5gpeOnTXpkPjGx0jaEBvzJi3v9gAhNDBYcxiU7Yw7u6zipgxvMsJ/Y1
pXbAuJMpsyfwDvliIT6Gr8bjNwHNZo2xRfHlvvs/PhfCf7nI52UtbjkE9gqt4dZP
CcTGPZBBjw6oqBmPG1BOaJcX2QezODyphzLJZvjg8kaU0fYWTT+T5tAkwkP1TpdS
w3l4Dt8wAEWVZSCbkZIAAi/QO9i6QRe+hGExzswpB5p/FNH06EzHHqv9gFxOUK1x
ODRr0yhQ3QJow5zW2tzS5REHumg6mKmERgHF1SJXPOLMzpAFAP6wkZMtm3iTOg6g
hcrit6ToJIYrzqH0oojysWsT6UDxpAhaTB66JYwhW1Os4WgIhCT/bEZGy91HK1Da
FTd2bWFggqgYYlTOv6hSchLMY1Hf4E5aHL1NCgkvaoIhWzvTpPMXH66JNF/SvYqa
xfkGmn+aADHM3v25sH737Ar2xcSpT1NTws29jLmfkcHwGwVjdJARuUMd9eqsWO7Z
LEXAx4p0LgTR7JUjyW8BBUBLldLPprIy02c7embdiwgOZWfao704FbLS9MyS9t93
+pdcK9pyFnSN1tpkuM6x8p7l9KkTmIWvGEOYklu6sfDxq1zvfsFjKj7GFMT57MHT
iHSf4JRQrqCCu49YnU/5n09wFK8/JtXkVP4BtYFqvCWQTu2/jB15cFAA5sPZTALm
u3ns1X+66tI4fVGqyYCeAzowEc45obXCZ3gP9EQkAIUCvFXAAginbrhS9bsMf2Mq
JEXuHjEBAGxNQbrKUPS+gj4RP2O307Za9Gqs4aDojmaTgPSBFuptW/tJtnEGjXcL
DNPTQQXIZVhUF+PGtd456queGQi/owMG7cDQQwjsOArZJwLCNnNDAA8rM0AbDCGv
od7YnqsoMy3A3ggIkc3Jp783WHX5/17MjoQl7QHtb3bce93mD7aHklSVaAZZsmBN
wAzN3ip02YUh2h8+e5Ik8nZQ9sy/zGRPxOdCMuW3f0oDRfRK9qsGBMIlxpPc/mh3
GGC2vwoxV6bUZSMOrmDdEpfxm33ABGIuvSJDSKy85Cn7KdXbNuhL0E2BdAS8h9ip
D7gDQPaB87V5l8jYX3uazF8NNjArVyajp8ATbVVcSA1JyX5fS0+3D0ZWh0nrnL2Q
+Ny/ZLko7wrxZ082Fklz+hE8Ou5QuydUhOLp2GVC95gmmxAl5mSlpG0YkVtl92tg
YvP0PzabUmp9z1/IOeV0aLoERxlEs0sKq9KQNQmrmRqEW9grDf6erIA+Omr4nouM
jr5k2X53I5f0YGkg5NBkxLV9PUatoK821mrtM7V35dL1+A1j4Gq37yGudrdKPAwt
kRMRg3T+c+vugtoEGeHPnZGNfBB8JSUjZdCoRwbJsmBp2rJKKbxRDbiT+hH8lHGD
Pq7xGPVQJ0VQTzbw/nvZ+Q1lbRzw/0pqCA0PJ4slO7fvLaVzczAk6uZYarpFiAt0
gtXCd0DsAlSMTCjS3K6hon1VMw5jIDBsVXRJoCtvUPVC8aBFl5cEBJLXUJFnGQGt
3By00FW/VIZjzrJhdAhu7tlvwMlCbtFTG9xWKigqZG1xciC2twutrGt4ufYFuKDH
gD0R2+2uhFnoNeCfvaDXSxoKORBstaahfWoGgrMQB/6gMN3+/v7EhOgyexCX9ffA
wLw2K9o5GE1hq51VWkNaohxjUIg3zykV9iobdxctk3IZRF5Wp7mFjIm+YiPLOImf
aEOCuKoDnrZB1yVl/k10rMRzoa7T145dY0gOr7GidXKTnYN1MUzLur37qN9TdZUE
fJMPj+4hPAw2jFe3waxDv4eaFKc78So55q+eElq+LS/7mv4p/XEr2Urn3HnVsuUp
P1/UeewAoewJPL+ZoQ5cwewN2gzaOxOz+S/utkVeK/TMoiw/6FPPumq9/yTs8nTU
q8Elp+44YaL3I0rutwGSoMNfUTwJ5U3eBc1b78TJwC6DXFlm5t+rt0JL7+x2p/aG
qMt1/G2Th++P2DtOcSInkVjDTLShriOpkRwemEOis55lL6CFOyf9sxzPz9iCGPcA
kPiu0abukDmjFW0igs+WTV4Vsapqx+49GIKaOMPDcyxPA/ZjMAqImiMtoOS6K2Vp
nAihtAxEZK5xB5gvci6SeFan4B1yMKOLK9T6qyq5GnVjNiEBVjlBMSpleCV26tkZ
PsKQAlBmeYjJBvOI9MhOjs0+5QCMp89M1HjpsIWabZovveN613r3gWmP4oFZMaQJ
8ZzX4tRtlEXQ/HpJ/qKdGYkr5A99eYTIJ17Uf+M+2dQ+ZithFKMDVxdRYwl4hBsQ
qnT8RqHy8vqSvuc/4gnEj2G83wmA1JmWpxyFk6pZ2BM4eJByMhCvoCnaKfmURnR/
lO6zxK/exO9bZWi1Xs4pAn4Luo/t99us/Gri4bYflsxwChAmQbx2k+nof4swDU78
Nm4Lj290ZxKUoggq8kWV0jXRLRccUbXqBZPPRxUvdS3LrstBcsCDukgBje+1FsL/
eFwagHiWzlGNto8gyQjK08um+TIuglX9moavjd0P/OgJ66sHehrAVBBEj6umP0kf
vteURUISIM6o2DXWA2aBfDInFBTelpiVnJB/Sk/g63HLOXw+pQFiLXpJ3CHxJLpa
9ZbQ98y0CZkq4YPCGzt0pMt8vyQjJ+rZ2gYsyEB02LpQ6/MX6L2ddtrYg1jhLmvK
cWx7hmNGW6o+/f2Xz5VU3rjLjeSUu55ClXeqBSLEKJqpSti22zraGft54qZGYzLc
XsP4t73L3VUA7Z2bwLcMdbLdimEL6Bqrkj0WXqINdwzF2Ia9hhCPZL3k9Do8DapL
KCgMbAh9j2wBcf0RiSA4g/JDv2EQF/99XkbirOhG/pBZSjdZeU+hageB9Pndhvgj
/xYn1W9LpkJqbWG/x80b6q1rOlpiKczRKzebbwA4TqxatxxB9HP5pgc8Q6FCdNn2
dBhGkqj17DaSDFM3DovcImvtxE3fmsHglOM0rww5JRbQ0vNqphlCdP4oSyyVuRky
WGai0mcA+zcmdS2ZXeNYmvPDWpTWjUSzspcBhJi6P7ST04JuH8PHqVuAWz31iZxg
v5EHLcb/UYu3Sw7CMKtbdtoAlvVa6nhvJIAuY4yz6QkWgx7SCAERhwlR1xDF6Hrs
2umZujdd71/3WxAFjz9xNI1Z1qVPKnuTlKK9VLXTa0tchb91RnXAG32vSlShwahq
+GUkDK/uBndfU2rFwL472NT7u1Te9UlBhWu0e/NlO+ABI+JhFZYV1pQkqsxtegQs
0vga89X/Mcp0VlUFZ8ZFOci7bXZITFGOplzaEh4B5t0Ew2jW/xslKUMNVjapDktC
ApwYExeFAzWnx12L2OyKYheYBKUuPva6M5Dgfd18+oKx9jL8NgLhkkTdVqRSsffq
U78D0a2PDBtQbgKwcc101cVUXZDjmBnj/hXwqTtPBhIT/9mGW9FbM7QoDz+Kigyb
Gxnze23iRYBSVZCOs4RKHdMO5Iel0BUUxYByWVfAUehwwur85O97/FzXEfnlUme1
MmH1F8uU4nF0tnU575wHZGCaKlX2aQvfi8VepN2XYW836hACFhV4BEAIfWi/X3Wx
vVpT2fxJtLrnfR5wfd0MhPRRb/U5oSPRVPDyiGTW9TDeWM74gYjCBbsaHMzstfXv
E1rym0jlRS94h5R2FhwQ9lyCMqA801sn/jXGZ4+C0SiJeCXdotlhnCMKEh/5vdjM
NcKbabRE47xQvqsVoqImvAYyvIMEP82akOZUFVf0siFGwchuNlDN6g5ZQaCxaZlk
3VzEIhU50ajfk04MYtEHBPBhP/x/105W6YoR6QCdZ3onEnwJrVJqU5kt0u/k/nVn
aBG/yLAOonfNmWbcP0Wwj2VwyQncSdA/ZpntTHDuDMGG2akVpPQB+uEUa1RYKjjC
ouEBZZ8OrDjMfQCyb6mghKxB9t3oNzEiKMi2hfXPHPjaHLp8baJm6X7URTTeOjcN
UHjXOfB6c6s0Dmqp1zkY122xiqqM7PWRhhhUKoqk7jV5/V9FX/n+dwvDu/1+YJyf
7c8Pr1n8Gu+iRPBx0ygwoCyUy+W25JiRFYBP9SHm5VLN0PZoL0+OD0nKIdIHCsTd
aWXO6hS+pqTOq+dSXffCZysxFVhyn1Hz+d7GZ3u7FjfajT5m6Do7TqdUIR6XrApk
iEFfkHTAQOgEdi502SgvqqsyoD4Ib707OO9uZmHzzWiUPU/qj9WFGHu5zrDVN4he
AfidlNZL5KaYthhqZNzYtgRApVQzZIXb1K/Sv0Tdek0qOsoA9ocFZavMr2sF+Efk
i2c8nTJHtkxCru4XR/rgJMh7JGr3AKCPL/hoYSX8ekmnpt8IIxA+VvdupU2/ry0u
HEEZ6RvOEHudNrBRxgxFU7tnn23r57xS+mDg4UNpjS0l0ISNaEBIea+b8ze1N+ff
i9jyv5ycN3jo4IDP4ZKcaStng+w6Pkgt5CEYAYVgMwt1pHf2Bi3iICvly31PIYxN
HB0J0JxpSFDfqDXuAGO8P0S0Gtm7yTLJveRaG1K3+d8a+Yo7znJ++Yb0VwdnetQ3
OmCyO0+8XL9noTcwTjovd0lIVF4JdwxA7bcM+d0PYyCPghx+E9TVQXAG51kOKjuC
AmNSmn/6S1B+M27vZtADjX1waK7tjdGUpnHahKNHkySpMyVVHDY1wRUMSX224pVb
fpaWtwS8sZaI2KWSfxT60A4450x3UwaERoiTENBVGyhWmHgq/IRRXsR3cGOs4UKq
BdVZy09tkNqhNwTCcAkQ+er9GAkdcFCfH5Hxwa3nYGf1sYoz9znTMKxlIpwZZckP
Oy3JSAPSug61kJZqBT9HXuKj27ui/tnPNfKTgYpINnS3drJzYhjYTVDCMtxHz1q1
aHFjsUE6rJAYRouT/Oc5qEMqda+InjIROjqBZ7ua6MQoX0K+7txKnhJp6SCzGNZ3
igMKtjovPVmPrDKhO94/PZvRE26hN1wW3pCvTANVbiRZl/yrXKvz1t4IVTH7PFgJ
8HumInbfbcdjKg9EtG8jeH/a8dLqYrpH55JeYFJPNEv8TVo/4wYuS5YmkY9/4G6e
SsrcZjmxnkIMPQI47m8IEk1Pvb3rnmmvKUZe8wlN2caOtAp0+uu5DtuR5vLdDthS
HyWdkDuD8reMzxXd/l+WkzRbeMHRL/TS25C2xzTrdP3rZckTWxNeTVENafVmZjsW
ihZZsk4PKlRFPXDvFa3x2+cvvqPEXDX54PDfcu4+5Hh8a2KyjWcR/sh6/QTZQ5Ef
ht7/ZOlgrEn70MX7v4uk6fWtkooY6lI/fiRNZ5/h+QV8t1wOPtLxkmhGVIaiRSxb
icUHvuHi+4aRPtpfB02HAHGsZ3r2gYgCpOSvZYZ1GFCLPMi5HA6yDQf34co/t6ip
sbhl82c8r6tQArxbMiIcxTW85PtudPXF06bkB1dDu4A+70Q318ONJRXuhDjMAL4+
i3p8bPKgthG6/ux2RBsUbog2zqN4ROp6Jz8a7sEuoswGNa+qBD45rOdPrRS/VgvD
Om8DeFtLoYDkfsxycgxEXpo0H6blM9TZRYKDJ9U1iP4AuuEfGvdIO2giCGf/9qt0
cvubHEJYZOsOAP69DFdo52AQ8msn0bqnZ9foNQhAUFVzBnT1SF5Fnzun0vkTkCw5
Img4dwycH/JdkVI5541cG/0vqFD267tENuugOI1IGSrmz4Of2ZdgowRVKeUJn2bg
wiTtqFEWuiOZrLGSX7J8moj2aH5E7J4qh7306HD+cQY/97T+xL1G3h2lRx92/awq
3y65MiJIKvrAHTPNPbrhq4MkHtANuxuRxfGYK+9qQN6ZnTE8TCamXsL2fjZuC69o
3sZkUEc99OIfRggoMCteQt6uqNGe6ulNPLIKx9rQ7uEaawJ+/vIrOTkayVpPqJFg
7PVwLSOgU3NOq0WBnnWPqBnx5fkaoq4U3YM7/i6RF7ALGFIdlywVri1NoG/amOwI
g9rWB7+Khpla+W61rvUkOVn+59Q/JzKG9FJzvLHmZQdgIuti/i/6asEW/mlcRT1S
zsXFm6vYH/kPMt+B8fpV0dhQAP3aQhbGgNB+WmrB4t1FRSIxO4iGB5lHYy2szZ4X
Gft5hv130yaX+7ilTk7WrLzoHxJtsiu2As4phvaj/2CZcnlYl7nWBoxRUjETO+fI
EErsnBL3f7RzXJgeh+bTICTnu5W8HLFw896ycdfWs3rUfd5V5kklB5uYF7Obt/t9
uc0zBu5yAQ1zaMIadvakyWAUK3Mb713/7iZ+hLJtPqGKWNMoYKg2rjqTz/n6y+uC
QjIQAbCdJAQOTR3ngEdi03Ph/5eeIfBPUkigPH9tjjC0+McqCl1LspEfaWqWmB4q
RWjKs8n36ZJFHOpg/aqrdH/7OKCHX0/CbThipqUzSlqWdpevsu9gobey3E4UEAJ4
bQQOc4VOMYz/kvD/l35wZVex82SnfaW2kutTOeqWL4EZGJ3tSzc/t7DfN5/O5gBA
SEgFpjF2hIstJolMqJkrUIEo06qanPSHLq6Mod6kEXrvNuRV8Rq1ussH9oaQVz2G
OliQ37vF8IRT2DZFH3tXAQcA9OyRh80BZxsQkk6MWYRSAvONe4PZ5DcP2jqa12E4
MkbhkP+j0KA8ORfGc5IhXlrGqj91eTpqmdktw67g7OAVWpoA/klUcCCICa7XHURj
NEx+kWuWtLee3REqUN0oQw4EIxllgI6pJaIIQO6Wk2E+MvCTpkRMLJ1Tfx6BfXPJ
EyQEIAu2nu/rwX1rz6aNxyCc/H5T7xs0IKo+Z5F3qkjeEgFyM9t9NOg1BHE0a4Rw
sFjjFa9b5nSYgdGK6VPqxZr/AmRU/XA6DuPgaBPgXZ9KJCfCD8w3mgDR2O9R6HhI
r4ZFsXNIgTkaGNGA8p479AwzwyYK7C9tmmz+v8xNY6zPSM80ntmOT2Ifu84FoDMb
05JWjxJAfejZSKXnB3re+Vw9vJdLvv2NHz6JFCBHn7/Y4xwt8gkeC/rb1yTNHhEd
1tp8BF9xFLCGeBNNUmsBGQRLyyYibGrGYn016CxhFosf4Dm7CPuD8m9EQpZLFLHb
KyKXyrVDU6CpD3N0NVp2LWGOnINHC/sG/lvVVyaqr9S6Hlip5MPw6ReBbXVwlcfm
yvRXo7FY7NhXX7aodfrEtzCV0vgg8VxGC7DHZfzsb3+j3C7BmtpxXLgF4jQpPkEp
2lYV34plnUbnEEEaBNXlYGkZiKqncabaCro0vFhxl7CuPydYKdQlAdKIpef1aDAs
L00er8z5XxuO2nTd5tCcsIOV8kg0ZGOmnK9xRfF6YWd9JGMJHIPF9C8OMqmSvuu4
lIieMUA4z3Db1jJgowMg0lbZOXE3ucLh417s5rgcvbLt/Xi/VlQJG5nlSIn3MRSC
LQhNtoEZdGIpBWs21c2zKEdSk3q/ocIij29ormuIcSvGtwCU775e8HILqydINy3p
V2KO17+wBtOwOHH/m8bsF2nv18U46tBgu0aAi+YILB4kr/4F1jj/A1lIi/EKaTe1
v0GxnFo/Q89Jae5LhWn6RbnEViWbQwh3wC/UIlpvy3pW9M3Gxo/AZottUTiyUt1I
vuyTYwSFN+lX+7c0Tq20CMrUTCP4EQyWC08L+tyaajFwdu1EMO4xD/KJO81+ZZkJ
TNoom0bAtV8fP4RL4nEQR/s4mv7SdfJJX40uqnOZJidKjiFfPqJO6WRycW4hYcJa
ZK526Y9tldHQ87EkRYaVqy6yKgmwODWyQJDYN3ME+LbkqaPho3EAQtLB7cTJi2q6
3lHBOpSNAP0owNMo4CVYh9rC07zxxZ/LZsLhmNPB4hOCKTfgsvs+5XkYm1YtB3nB
UYNnRMB+LuaRwJawxKPuDZZrKgnvLkyyFSRBDdTymYmXURJ2nLHTBI6r9UooWw7i
u/Ay/Aq7qSn6sBAGQPyA1QR6RGCAyJSs0HPVMSf54fF48oFhwqdgdTl0DQJvCkeh
DGJ0aOgCuWx4Ud/4b2DqONylrKxgMhY0bKGtR5+EqtH3V92mhj04ZqZK1vrEfSR4
ZzHkrf2flnJZsyAfb8IfVNZCx5dkkSkUa8SWt3lweHnvXjB3ujsdVW6vxbi7goy/
arRVmX0adx8JWY0DeGe5kNdtH35hvx7HPIVUUTfqAAgEfQBF4/nTEa8sO7YSsUyF
c2a1PGdFCxAGtrajHx9DY0vCkK/3ifZB+Qq02gP5NH0b+W0t0qcwbRK5wG64n68o
uBRLw4rn2UtgUzbpjv2ASoWS3iwNDPRRkkUTyL2sZBeUxyUNFAzlkHo+gmk4tlRI
YjVDS/x6ssd1/5NYbB36RjJ9LpyirvS/TWfVfIELioph26OMradu0hkM/67mmLsS
WfH5q6aGc666i0h/c87789Y5LqpvORoajG43KaxoftHnhKMCdRrkkMP5ONARiIls
zRmG39J1i/OXMh2FG0cSDFNz168F7YdKIeo5xeyDMMeqD67BXDh2alP07cQkoWgn
aME/MN1Q9/bDjhFb3BPRfMM8n0sMKhf/k3fRhRfSFi5filhsRyfjqvWm/9aJbJfc
kfH3hNetqX+PH+UrzQSqfAzy7PIV54E/owJpBmlUfjWXTg+rmzsYxwdNeLsvlDY3
BaF2PRZRJQO1vrq+U1TlWEwt0ozj2SLuJHt4bbj86uFrOzjnNsvsd+cbDNPf4b4j
jlbIOaLW1mb8jtU+VrVnQOROa/GjlwehxzeeXI6polWUwSABYHSt98noxnL41NVr
j3KMIUVFFAAb9kQrNOsblqRjmECFXsd8NGE/gKJxPlT8j+UOZ9P/7i3mZSyGsijS
mO75b+i8alsi1bBpsQ4vkWrMvfrF96P8A54Zza1kAab3IVGBKxV8Uzjlx/WIzDOY
4zxurDYBBDUmE7VyySpz6tn45u6JWlsZQcP204S1IqjU9b54mamf2cA5xAB6qtC5
FrY/6/F3NrW9l+p1X3y5uqYJol8QgJDAtYa5Ad5zKZy7JJql12Pycom+93vUeUl9
lC7DJp6OtOpxqGE8Q7fouJH+fEJvaxoPQITFrGaySnS/4PE9X60O4sjVSGxQPvQg
lUNUrX2z8voYE8as4CNqe1j89eFx3TUy0HcF6HU16nIJ0bphrqrYR+i2yTJiAjn1
sO5IiGZPzLa9eSmdIcWpO5IMUPdbb5dPeg4YGNnkWeKRWqPWmznOsrDB8XO5DCE+
LQeVo0KNo2b40/RlzxyqQ0L050ZgAUNyxwi2A5Bnfn9j+Mv0zAUsSXQ2WhzfHOql
TIV7Rr3xIZOuui7ouioep0o6NRsi3gDjB+kn8tcoYlk8xhvG00lgUlDvUWJ6BrFH
Ql3vmIAPccq7AGSBpV2n1CrNoh2rggrA+ez837iIT+lv7Fecu8Tx/AAyKn4Jh+Rw
DLtufwFF1VoozLen0Bhfn5E1YmNlRgGGbrmxJLZ+Cvyof4sP+NK3/pSm0AFAF7Nr
HiY2h1UlXRwLIrG2V/ng1cGQVVXI6RtTFc+HF41n3Asw+gXj5UYTw/W8d1gm/zpo
Zf9WUTVEcYqjez5JtJwBkU/9dw9jUppF9RmqckhwnUVGKw4Z9YEBaFwUZUZ5YPqu
zgczBaH6yV66fKRn3KmQv+5u4Ob5ze2cgGYbe35G6Bkm5/3Q9rq3e4na+ITNIZt2
yzE3cpznhf0M5m3HzG5xAYxbj3BmBQc/P/jmi6vwKjQRm3oELWH//5LrFc8YU4GF
Ee71O7msGdpO4JDermu/15OtlQcegmWt/oFPT0gdmP+IbobDgD4JJSK4V+zlTiRx
SHJONOEEKkH5Ba0d9ZwaWGL8b/F9OA87oTd1a+HQ+S3HSs8+/O1ojqD9mVGyC1Bw
95K7lBarqur4VUgTIDsjDrxS38p1tLE39yxtd/Td1+nLXulj0ilCkohIlJ84DlGp
/+jwQpgp6odDDzZyJ1jl7lJfCJI01xIc07fuCuXc4j2z/SkSa8xBrSdo4zjEWk4/
5drjnuc9q0wDtVq/8VgJX66vor1adrLt5v3/eaL2RqOPBjqODGR6+7QqnDYDmcr4
47tkD5GXrdFYFxiqWgFuu69pErBbpTrJ+ucRjBB/mArGEK8RziVqVBrsYI1NINY9
AEwBQl57XrTWyz2MBBRd9hMGSCD0SgYMtjmiQDvXv3kYx/LctSlQ2/B+GPZIS1Y6
TtCsb4aawz7D9xrQQVlooLZ2RR5eUHncEWSsiLUxakc2uUfiS0ut/jGGQ6pUAFES
U7lsYjG+cor9mJd3zDGIYlljKp2Qpkpm3C5JqJbo//pi9QObOvloEk44CrXEkFwX
99AeFy1TCSAzKwhLn3jVlp0zQEBapA0m5xdRvjMgj6GAPlVNAXi4rsWIAyFfJO6s
Mwkp5EMYJDdrKFRv6xYG4DQuorPMD/7aIELV6gq61xnXL4YUNzewx5qqozFHsci+
S+4uZQpWbxx+DloW8v0Jd71HOckqEcZLWz47skchdL/hoVyOYsJ2pNRoDOm5JLru
7UCOynqpmgQaLv8Qp+KVq2JU53R4HDzEMWgz5ZKr7OqxcNsMkwdxg85uLXSCplo+
ncbWrTiyC7Hvhq58gVQzrbomiJ8/j8I+2CQ8hVozgFIHItXrjHMZwvJF2JA/h5Hs
Wk0zYGSIDN0Kq2VOAJIsHyrDqX8ztlLbhS7qphSCf1u9OisKh1usaexR2aKWzFiv
dCC5kqqsrtKZ4KK7Hg17aV6T4OtCbCdkIaR4sctJZa/A8/58EqGuPagz3+x9SEtG
T+DVxvQe4qLG6uKbyWHekwbLKvidhaUVEcYYSQ7Hpzl3swEHL3T5phzBX6l7KKED
i8JVqXmr5T/SxYX7STbLKWPN+nAN0PGdOKyWppprjs3N7jO1gSXrBwgqCrPMXAjn
TANz9LVe4W5E9ODEVvfKRhjGi5KYguNex1dXRx3lEp8E1DvnM+evP6QynJIVdUdu
xaxasDDdSxFIcMQTJ62hcJDrTXqX1iv72qpHri05nWV8bmHtwgse/ay5O86vi+aw
KHea4RuTHYFgWAu1ayG3AozVuo2sikG+8Pi95BjVP7V2e32B2f8mYoeO+5Xmok+3
AK2bJ7LejBOL8XZMclbVTKILY3DnDT9KkHVV/b0Kzg5eyHyQB/N2LRVZfiNseieZ
w7VxVXkyQQBFs3zxkgW2ti6bqlTChXvVqh35l2mVLghUSEo+qIep+zkrsT70A3KH
7xpU2pb6z5JxjYutxvCsu8jLrwQA9YzeXlc5y4oRLhnQxcOC3aMQ9s3RWXO9Ks56
GCdSJhw2nMuyHM5pXetuHd125D17TNqk1bXcgH8OenYgxaJGyFDy1tLkkXT30mMf
nAo9KOFPJYvJx37VMlANZQEWrhAO7OgRsfj9wvE7n0WeYgWSpk3+IE8q7K+mF3eL
CIxslTdYRQIWWJIoL4nwU7sx6uYYoPgKQDFVA8ViRsYFf20RnG1V6DToHYhXigZH
iGqf/UFWg1cOQ0keYJ1DcjZEC/YboZG4DSOBQD0t5TwQGYoRu86MKCjM4g71rs87
LoDyfX7zs6QsCYnldjsa+plKcW4U1HjuoUnc8JtXiVFYHu5x9bEyGGTZ/Ae9dM6j
g3zZ0LNVjOVV2ysUBG1zT5bdMfs11shZfE/3hTJosFrihEuNovC+vOVgPmU5CH/g
mHpmpuua4e51ZL3BKCAILWvleZNDZQOQZ8iQayl078XlAEuhj7Aq+ZAnxyAt4NQW
xkP1vZfSGCaWkhslnTzSNH+/Qirk5XurI2olaomypQlWotvsvmvYBb4psETCrnDY
NbfvgGV2NWXSLhi3+4ITyZvOF3rhhS7+dcvwCy7NbEVRnohmQ1qco9brePQ2IUod
Z/fvkk0anjh2mI71xYlmKiXZucbO8RKcwOjwRY55BLNL0IyZAog6Uh13y4vCJe8Q
Csw3ljIKzaI9qakhIxJ4P9MwQwT/fDr2L/zhX72g+WXiLymfrvV/wZVSF2PAkgjy
yXSu/E8G5OvYASIdR0utJHCpWl6HMYxUIC6mTwtVoOCEqX2J27OoNP+3pNzi1iJh
kwK8fLzop9Xe1kB3FqMIC5ey6FgMvLy+twEzvGUcpjf5sQPBY2n7rxNuC9lJL1jP
YCSzMm86NWrCqQ+dBcNFESNGrs7G2ZECPUIJf/X//t29+UA760NCasXyu8ZPMreE
oiaITra5xBAIbibJqebciBQ/k+X749OfxufyPt9AN3GqHTHBFUa+Btsf0yAesHbD
4SS8sPQJNFIBmpd+exYxSMqZjj/DJYSVx92wum9rZV9mRUbJbWiSFkXEmmEqdOnj
2jlj6N6oBzLEf8s7jnr+QhpFg251ZDxoAC9XC+NSCWdhgUYjGlxq+Elwi0l0oIhP
HFZzPe81c3/1fxsn9TcBbde58D3o8HaSVQo1hHBdpM/lf+rNizuIyjvxevNYpC4W
JlWcA2UzEeo+MC/pFCqCki5uNUP82Nki6opPpDgxoxX1X/xXFffVfcGDXZ1iMUVQ
njwRmpHK/QYLCavbtYYawzEEPrKPsGUUuPhhTW37k2iCh0h61os7prVUFsOaF3EO
SQzFTtxoarERTvbeQkE6fbOZbuOtDGC+xgSOct14euXIwMKT/R5mQqxxlBK9ZOs+
6PLmwbS2YVdod3DtVYpdLpGpmAlWPjMErn7JVxiONf0CYDxHDdfg9P94edsX2btX
yZwz1Uv1Y1Dhf0kYTE113mT1gasQApByadMRo5BlExkr46r+4Tm8Ih8/jC/DoDA6
Pw24mE+BOyeua7t/qbq0H418smasJH+8HaMxIh9JB74XZFDeTjhR27MEi2IaZj6z
2Fhr8MPLEMuXtnPUjxAe7JSqV3cXFNv1wzIWiI44wiBSDz9bdVNiodrp8mSChTnq
LsBgz4Pwss0SPKObOvxtc8yaUXLX2ysK0gJdwMLDsHIPOjUmTgkjLTg7swN7SVf5
ty6jBQ3r5DvXECFILVDD7IIHE2vLO/aYsu1Av5tzko8hwILF8ER3qA7xnGkoYlom
R4vAU9eX1kl2mpOy3Gb6KODcIo+X902x6gC7DDLHeaS6gh1pDMdZQoMpiDB/tgJX
xzBjTt8h0mrwTTzAMzyOMx6A+k660LNlVYqUpnsyGpkpIiyTohv/UiR5t6h07coS
c/jphKMq4gm9MzRd/sdw3pwcsvZUMGIHQuyt7HUDbOHNhpg4QnBnU/PL+YRW5Q77
VTxsJYh7a+kSkaVUFwmamOAp1Ck84NjYXyM4/Ewb78KJhGRuleLQPSwxgkJXuREv
0JRWm4Btwvr4NLfPHLw/41tT77lCsPE/RASB6jEKNUvv88KH797IulisEEcglOJ6
DFsjYTWYONIhohfgqJh8bQDHTCQE1RsxtBKh5+wBzoX9e0dWyCq5xkH4CpavNKyz
uLoygCxhYdHIbsjWS/eKAYjR8ojijbY4eHWbzw/0z5+QGyVdwVmDSV8DJk1E+FWv
joAKx8IQzRl50s6+NqXdLD29K+R6lUbILfxNQy+zQr+Xx1hH4HSS32tklVpCMEeR
SWk1yMg+6e4c054GdF3gt1bx8CEoD7/d7Q5GiCPbemjydPlBpBuFlHyAVakLucdL
GbHsTEFltRFQ5f7rc6miWx/eS1VcKWnKlVmY/J5LzKZqd5WXkvKY9s0jYHnudHCx
h5x91L0NMlZ960B07024UEVgz/v9rGoAuwpUwfBDLQYPA8GUrWJ+cq49z9CWFb5c
XGL2fMWcYi69YeI/gdOthzKmCpLD20N4RDQcWnz8AVl5GQ2+yWItbLSFwDg2BAWk
47NYOLtnR9XdqAIdpLH3vvzV0Rusvwzaaan7qZtKfXfO/LhOFfPx3hSDT7Yc/C+H
TKHP9UXXNKKxKGbyDNx1Ef9+dqT3/I5O+ePJl4rNa5jdNIMjvP2eCB0kHObeUB6u
Y591COuixJdZ5qqaObGb4HQB4ncW+P8st4B/vl7aK3eSqxwb73L/jgemBIpti58B
ME4wYZ09RqZaljWDMxXI2F0x9yOIEHOywKP+kgBiiOT+tovxU4OLUcpfvMe0Tbx/
CPe8xjwjBa53jbI8f1sCEQCHrJvJkT0uLUMkXrJtVr6O9kMqKqnB6J9VkzJVP/+/
HvqMY0mLIHjDdCGva1+SBTWD8v5WlNhRprX2qbgJMJwn8WY4LT85SWbg7jjTuHQB
66CzNtysqFbqMJun78Vtk8CSkheyjFRSuUPzV2eaPfWFJ+XpWuJ6UWOgrP+TWxCq
7ZrFstI5n+B59ttNDxUOwTAU6/6jGtIU2lQnt8bH0BGda1qaTMKVJghuEt+GVFom
4PQEZg/ypODEyFZ85pVnghjecMSrWmTdvBewatlhdYkG3pqhBLAn3DuRhBg5nUAg
LRD4zjVzYnmXnVoBxZfDaJLPnt2O/82jHO6b2FF0u6rMTNjbzjUCgDyLNF6qlDZn
+lJvQntCXOKaJBzHOFvYCcvzFYt/s4JlcE3BiKAFG12YPEIwQcXN/oFPxYyCDzr+
+5bqkGUbHL9cjdZ13yb4k5c1PbaJ7iK63UJY3DQt9JgeouD3297WgKRd2MxnmNjo
FKCKJGsaP5yfSJ8Erk9mBYcump/hxn2Yl31h733eKCLVXDxlSIECohKHFaZIDpwf
Z7x6ZfTIoYApKESZEap313KJ3W7xUQxgOjzSdvheYs1FFDtK5G5g6h65XxfGIYmB
O8XUj9hctFmB8TUH77NgG/DFOzlRUWWNIXhO43OaythYrbivNrPWmFk6uoYJYJWr
dpWNr48yMDkwl/71659lBPgyajZQmIVCNQ1EZUG7MtijkpfyM5W/nu2p8QgSUUSQ
ThL60597SKYJGV2PElKo+EdOKnEuQtuHkUgRwtJ7KIAbq9+WJSsBtGlqWXTte/DO
skaTsm0qoZ49Y6Z4tIGsDd+p8Q0hjwkQVYdqp2lHRZ1OpI7SQW0eUOGnBbeELkEn
b0DUBs9pOATVIRdDtu+4naxVNetMuk21AEg+t8lRLgQwkLkjwXQxogXwPdo3FIEz
fcU1DNi9H9d58lDwQ+SnjUJt7J3ZBAsKv7I5CzOJMh9lJxeZool4oNnvHkGZ2urV
wPdB4wF7FMBF97Csz37xOG/lluj2QmewQOAY8u4Krxvsg5AUY4Klh0muhScoiHiz
zy0IwPBXdve+W4yFMzPIZt7JiUi2t81prCrforG7BTRdln6i1z5XyuI/LugLHj10
l1abC/8l07KV3tU+CDQn3AbEnKQlB/5EWpHVtJheQmgIGtQlzkZ91OjqQgvlJedA
fvqV6lqpXGBebWPVSAq/X7C4uBYWFhgqK5tXFNH8OjvFPJBaISSjMW/gLDRxCLwP
rUXV1C3ATd5IHPq0Zqdtflr130+iBtBF2g7OmonwahjGsXsGTttTTSzO+9a1cDTV
rylNuf6cqkEuwvWyXWs54Pbq8UA+JyxQH9gSnzlcvHbF+fsymM9fg4WoN5vQsrep
+/yyY7LZQkuJWC/FSbXcIrGb6enpmKUgMHXqbTkWTW+vOVqifhlQwJLemCaTfgL0
YAUswbFfpBo6EeaIgPQCZkZcQPOx3PzJl74IDpEIGeWDSY66jiL7NZ48nhnM2SBM
Yq023AYbavHXaxUrECTiDWTsIDwJOddlkd1wz3EINL333OobFwDcU4RruxKSGHuh
zgTq05yBsPnRpxzA+WP9mDsiy1SqOu1ewgb75gm1zcYotMNmXjxVFyszLFSXUf1F
mF3oG6RAvY44uqaFt7w+LlU6nBPIlFzbiOve7jltwxOhcfRLmKwltG7T582JcKyE
CdSH82K6qVaWrvWBdrGK6XJp4sOGEF2SX+OAiW0SIL7yGv4HGNbpej9CuCNNDPdb
RIdt9tGhKf1IS6OfIqTalUm1is4qqLLeWw3HZNjzahFCjRezPZvCo6l1oBMwvg5p
Igxlx5hzQlJgZ6HdnXNHXYwBVUcASj+LlI/ElFRrQN6CovOxyAFg/Y5MF1m+aRRp
6clpf68Fg10T7klBjircjxSHlbNHM7eOyTBaH0hDcP05o1eiizYiPZTo/0eru5gh
Gb1DQImCU0iWMc0rUcgk7yDFu0MvRcNM4XXRr8FNBxcNNIP+zmc361lC0+jRrMJw
nMiQFSLO6zaEkMR43VyEcr4+2E4VDZCoJw+DvsZ5HFC0ZOTrVksOZpJqn1R5e8WG
u59MG0c7XF1ghCDSqivgRmUv4FJuEx91Qe0i4rRT6ToMjUETe9S5f0Mrd06f6Wbd
HsE3ofbkL4e57dE9eljLuCnt7mgNLLbsNw21MK5PQqNt67cseOHUpkDwUezpLnV3
R1hDqgttnPwCBriwUx+p2jFNZk67198J4fydkKD0xdFAAXwunF7uwHSHVNwHvBsG
fsGj67ZuPZbx/xkrVkGl8O3BlGUgrcBF6fMx/HYDkh4rxQGlBjBRQxODVq/JqZFE
q+J3KzO8UDtnyBws0WiyHGu3wge2OJDts5K7Mc0JBSoNZcoP3ZdAX2AY0Adcu7da
44k2+sf3kk0yp6117tfYHV8sM4PdmEa/AB1SJDwlbJYKToOZDUFHTyoTx/b0c0Ty
Kl5wOEljZwzU0aFDgvCxhtIm3ineEzRNB0AwL7XWr/PyB/Has9wis6mrugSLvsaz
y9/o6/v1W2QYoyUjSyXy1SOkdivUbIgu2HUjoqhMsE89VNMnuje6OAhdIWxQK7/F
hH60m+aBiNnvTe8m3Zwa4vUtxzeHoZB/GhJqz/pSlXiYZwghQ4yBhuKqgxRSy62i
z7acKHbFRVjZrotIxdxVYZgWD+PMS0M/+RRfNoPih2sX+yc05dV6Ey6ab9RL+RmC
SrTmu2T8UAPJj4VhBTAtP5oj+MSBxopjHu+deIsaxuWHLI5Vq2vQvFTiZroaw+Ik
1diJnCiQHTahTJyq8Lsh3Rta4ar1gJN9J/p5fzcFTrVs6NQM0y4JIjLVLSJzNkds
VFfRz5GbA4mWpozPlKBWwa8TopcuNmKg2IUrUSnMfOMjJL3fafvkPHaDKZvAn8u7
CpWa20TbcOXIbjhSvxtWhKQ74dg6k44eHZ7IrwFP7HjfmrlixshbeGE7Cq5aGfk/
UVrL2QAIFVqaukq3iN+SLyf6ebdGuA7ll0Z56/6sQq3OP5wG9gEAVoO0vV2IoHjB
/EhLM6jCN0/CkxdvhoaDa5L0CvQ9Fx/2yWYw6bZJj+N1BL1DEgGSCcJctXt4JiCK
P6x6TJl/SB7Qx2tsmBpghhDsD3g36E6Oex8DHSR3MTK0IA4lHcXb6V2v3+TtZSUZ
QpHZ2eGLbxepOq48KF5OBrezWmO8bs+dzHFXvoM9Blpdf/kXN3QDbBvtR29c4/+3
tzWiDptR5I7tUBofFQ7RgLsVnHmnHA+A1hDkp8BrezoLsIYEsaSJjYbKtiiIPJ0F
cH8mVlqobAdbaGepjuIbeE0ypLPivH9WEMA5XYPtrfnI040GCmz0obHM+bdzbPyu
7sUd7yBQkLqP0/7xoTN4kkdsuwp7FZvLJlQyt3xe/+EJQvZGjptJaQvUS9aw12C/
kly6iSci8NQwnw8SsYqDwDL4U4s+2I7PYfEM6px8X1AGRnkUlg6PMx2jCyHWlmu6
/38xsaKq9P9PIxHz1AgwmuFdIs2XEQI/Pjb7qSNKxWTfqUN+W2fJA6JaZMeHz/o5
sD+7UqygEWqRFP0G/ff7D09Tr8mGl4bUEvkdvbg2r/NqG4vOl3Y0DEimUqezFbnS
YzwslFsZGp8BeqRLjS5nJ0KO4CTD3CdT6jCqUSc7JU/nA5wkDKsRA+xZK9Gy3AWR
64wqwoyJtySpJM0OPdPy7gpJKqIT/D/vrPIp7X1VALXjvo/0pfT1vQkYz5cuOj7F
Xo9bqk/+GnwXk8jrhgwD5wrQRX0Vd3pNR/n701V8RutLrUz8jyOttbumsfbgujqe
xRVA55HNx+wHu8mj4b/7Rocd39C0K1zEb7F51nRkOb903V1u5ifHIdNFDAcD2ike
xx8PRZriBp32fdb+UMSgbBm0KAaPiaY/xaar9SclZXfH1spaRUXJLj4HGXiGhNY8
TMJW5TblzDpLgi/MCzsBnjJSGqOQ7PX3SRWlCXepahkICo4H/NEjEmJOWywf0Of0
G0rDKtQUE72PGsmSghYjT5gocm0k7fRjk9ESD/lZOTSrzdo4nMyffC5RRhvE+KOp
ZlM556lnJ1jr1N+ThxLN/4tpuAHpSssUPCSf8Q9T4J89C/2CHs2paEWCGi7OyYhP
jrpUjeW1C54yw7t/r7eOJHdZUDwCjgbKfhb7nMWG6C/7eWWaweicSEY7mOcCng2h
wnfgc+jdzmaBcGP1k9TA5Hg3TVsVnKzLc5Tf/2PXGXpg5FJ8aDDl5/X89B8ncE8i
hX1kV7tfHqCkJanvfZcQUix6GbFrBZmaUYOXzG3MFV1ZDa//TmhMvTQChbYfL6t4
ZsFD/rA5bQcWmXTZvAEMbbv54QRw8gxmyK0KGDKww2tMG5dmvF+I/MO9GSe/z3I2
YWlAHcXsm9n28CwcHddV93RyUSZFcoYEJtdpRrDOu/4MiEAlKB58kPMlS8YriR/x
ldxe80rVEZdnp14ahgmKBqF506DEOIk6t8Nzvco18IYpD/t8T9kwTXxoNgOPxQF8
M/45G7KADo8+Nhjrrvxk+UjAIumIKkEk24W+a0ZSSWzBl6kKio6OuHbVTyazeHST
pLBXWSqVeOINPFHceenLevQtVWntuiK9yQKZj3wK0AYNYE3HLPRF3DUOqo/gtaTF
S3HayYGPcm7YkQ8a5+0xA23LYMFbQy5TeVfAYBQGE0vzUbb3RNj+Ql0wAUKZIuho
Ogk6eeKWeyfhpp9fcLuWOhvaIH22IgW+fKoSreaois1CZ9UYqy+496lva3T2fQoO
2UtXkhDcNh17Ewqvxc89bIM+Qc99wq1dxCwO6KGLU0wRs54YqZLGI7vpF6AtZ1sg
MOpQZC9T/EsCqeNfJtGdufnvSY11nSWpK2j20xJBa2UA6E4/u9McdoQ55/QC6j2j
gTStnFBxqU8a1VYsrmLG+BiOgK+TCr+1TSsnGLPSt2l4eoTf2uQuMt9drQPgmjg9
/sc0oPSz+HDoAob9mjYa/yT0dEJDy6kMI88mLnAfyQH4X/EWOoYvMYxEP97LAkb7
n6vsLmHeiuDPbhzpKJJ93r0h0b7N/CBD8HOPrLck5ZDrS2iHeJE8Qx8jnBrVExlo
ruTmprDAVRR+LYKnC/mT4DvEaE4YVTwtUJyZPmA4AJeyZSSZZimEODd8XwM7OgSZ
jU+YgCb5Q2OY6Zl9/30u7+56n+qy76YambOT24iP3UcOIthK8i8tT8dIHmxGDLuo
0u3WWXcNNnHIeMXSJ9XS4abbAZsB6cDv01PpNZJa0v5vn2UFlHg72Ih0io39UVwD
nJcIhQaKesBTR5tH5B60G9geGLeJNAU0dVK6BnK3iTOmIZIK+3XCc+whqck8AHlx
U8OsM0t8fr3E/7XnuEU+4gd/IYcyYJhdaEIGt9c+XyQfmBONese8K94NJfe1Y6XZ
nuu6sI4GSqQNgSlMCBW9hp4xvEMbS0IT9QW0i66AQAqc6ik+nLHl6zMM80AQhg5q
DTLQactoFvMkrq2hYvSuHYEm0Bm5R5Ppyt2Z0DCa8M+COFFPOQyZidjz4B3EukVG
8JiYEe/VQ0q5NL16QChQxj3MIeVOV0GgS9EqpriRr4f6ZP6MWsDTifHLh021ZQV5
wemB+vghJ+t+OU3MJR8j+lxwAVACHn2yBG/5aE6rrcsMzfV8EeXc2VKa3NnMW3/M
CBRXvxkTvlpRWGwf8iY+tAezy3Fe76apbTlWfA3wT82HoT1tUUi0AjoPtGTRR59F
XEC2GV0eiDtNZ+iV5bDrd8lOSpKNceaDAXYYaqsvcM/zsyWfRIr34Lv4mKpBYPss
sBa6tK4+iZRMZKhtv+2/O+cgHfV7Vkq8xSDyU/Z0pJNUoo7P2aXWWDrya5R2Hdpt
WOE0i+hJip8j+o8r4PxMNo7OuU4Z3FH8vL1cSHVsSKOmEXe3QGf37w2u2cuTphLa
8i6/31NmVFyraVLj+AjzV75rdzCCtQK6T4QpFReMZ8mTfkvEPZbQdQ+GXeg+jByM
/zG5cO4Jo+U1aNbJI6S+A0aMQvJ+7hK8tY5bnrTtxhQ+WvHe8BzSgoQXe0fiyUIH
OWLQIaj9iYRYSrifuP3WzAsjTbgkIouHzDV5oYND87QBwrWNWprqOHwtZTMvysG/
AuLpzattUaSP8zJpqt4Cfsw2I2dxrIIE9RDuEmZ/iQ/028DdLvwZyQppeHfoeBv4
tS4cjFxGInSkDi4/1CF58GPT0b+X4WlXLg43oMZtnc7tVrK9XEbHANRDzgo8ySca
EpNJdOnTjvM8l1VN9TlZHuyy6k5FVRHt1s7YAirHWSKcWJo5yLWCzv8+hjhri8K0
E+gAbV8lhRw7255XseeZYUj216/e00BcQbhUjKFTZAV4i2ym9VV4YGVeqqAsh/+E
gNQcHlGwkEQznombuMODu+5qBDhyC/rCE6PMowIRGwx/+pbAei+Hg7sqBA32NTq0
Zkz5PMQdVtpH5SeLx7vYbg7SE5hq80fyDQEJvA9vG+31f+Bce1zVvt8HUF2ny5jT
2YRQ8SIv9xswpLJVn4yyDOJLknSOPGQ4uqiDJRCa9FijsCagRBJctwX7y2rfmwgq
enwB+YTYSEnsq9qcJs55GslVXHrnQ/gdg1SYqrajFe5KhCZEEf8ZVlE6aIv9Dss+
XByLBvwZr71cgz3I0wlKDA/K7HERAf88YzJr8x2TUFjvDW9tdGWGFtiCnwFKgpBX
meOcGjV2R9zNIExlO/rmsMrAyoyafbig+KMNHC7S8xdZXEsffGUYmmWOp9m8E373
H6Vo6LREVXSzAvubtKioYd/riiftwcHmYRU+Ztyr2IFR7oslIBWxPhtZ8632PlDK
v//I8MtMZHHsZ5wnpyJMNP1yTD+JXQOlfQx1cbwfVOaPPiGH3N3QSvbLNE6OHMOP
RiiT8yIKHoakjUEviV9ruSh3+Qj3Epk2GVXgzZkfTQmtdESpOpPD/FUyO/X1u2BZ
6jBkqNlwM4vBvz+1fZGAF6+E6PPJ2Wxi9phNtmLOXH2Mfyro69c1E/A23wToVTSA
f0amguYVXqvqBDo8Y1kKBtqX52UGK2HqlLKQv/Kx8wbLUCErnw+odWJBqWsRlCmU
y0D+e1QLXvfeOTbZbCPP39B3/2Xz/jd076dYgUtyUb/zvV8MdrHAhkc7ZRIwWO8J
rbCY88ETSh/uunz+8daUsKuqKWdZPaGdqriHfeKf4V68tniKOjgR7dzusSyS9obG
yGMtRhSUzU1qT2Yf8xtZq5MaLIfH+v+cXPld6jgQf11IKKBoYAKs9JSq/lR9GpvL
QwMD8YCcAVJ03ietMSld4s4stclI6suXf1wMkvIKhnTgwKqopmj0ach8b/cQhacU
kRyBoVfDpTXFLS+7h6ku1ehZxQn25rEtpF5+nq7hQPH8Q+biEI2stCO0S406xM1Q
VeFraMd9X1xTg2xsYbyh/zuEaz+iCPbAuiI2/cYCAMGf1f7KponsHauqhCx1E/+H
OosL8aFEHfhLBnoys9DVgQc6UlCh/XofFFZR/bmX1/q4SOE+4jWR9yha7wkb/dJc
GOfPjFItuyaadFkR9ITAh6/0uo+2Zv6yRw0sYoXL92cDOCgXnr0NLJYjmNbPS+hn
qtnqRQbe7sDFF6MpOIlriw34xXJokyxwLnHoNtOzKw45XdOpn76E8iHx400thOQr
BYdnuuZPLldhq5f/7IKVeCdahMxjjpDbAj83uQiK58m1OsHO57kXxLx8jVtAxP3h
RbA622qniVQBjhSu5uabfTAAH4L4eRk4YXSow3kI/nr8x/fDigiSH1nv0xr/ZIxI
MePmweutMSi8rBp7Pjx4WTTNRUU/SVUy5giWYqyCXgJI3lnU4ZNi2GnFT27+jxqL
gdUYe3j1baLmS65uUYQSOD1Ej4OZxhgAP8qyYeYjgZG9FwrXmMlPzWelkFDS7tJd
yVlBDwn8ymAkesDBeU0WScXGYZW06AAQsGfLi82WGJaL28NiaIDWea/yn4byDZSW
ejdBxk33WVOt/mJOHR2QSygyel5zU10LxQwK+nR7wfoKhSWaspS0SJQCNWtlL+uw
Fgv7fQNBzqhUmU+wTjrn/rq5SVLOlgfsLzM1sJb/vxbw4K4LGwettJ7SGyyA3F9e
WOpD7bwUER/xrwEBvsQm/2ZOHOX8PPyX5FVGXmSB7ILLHw1OZ3snPV2Hvl3PcznK
AZJ9rAIHFJCDZII7tImZc5hMeo8PuvAEX/YE/AQ/J/PSA7alax7HEP+y09KAKCAX
LnxGhXDJpGHGt2Oqc1YIXonWhdSvM5tyUTlHejVXWaiaYBsg7uS5ESqzapKIYEHi
peD5EPyF2w6+ZAb9N3iqNIRRbRnAFh6VPb/JYcxydgFG1tIMN4tFz4mzc7F+vaXy
/NPZD/zKZ7jemc0D+OxeXJcsHCN8gUa3z1+jYfaTnXf8D0Jm0rQkc03n/7Qd1NgW
86VgOe6tzznP/sm8qMQr6CiULAUfgeb1TJ5jU2bv9PKvZ8gSx60+SLu8jxtzHalR
ATwPGT/P2EWz49gFeDb447qdjUNyscc+R40v9Ts4qzAAXoXWeSexbp15xN7y4XR+
c7AbrxeqH5zd2M4sdOphu/ThcVtJeGnscu/V37FKl/a8/WAd8ZDN5kYA3mlL/Gpn
dd/8tBXdpy34adzH1G3J/ZRmjBq8Eg3cD1aNEXnEuTlvc2wor9VlrA9Z14hWbTKV
a7GpFA6qSpKb4w5yYSX3VR9vWbFC9JlkMX19i9lpt4wJwAAfj1rza2yZj6L6v323
gH8YsLfrqiJaGO6A42rTYmrUkxh2GNZOBqdaDuSk0J4oCCSv0Czx+UGjUiRxJyvT
5hCsVgivmWtC7/rw14GbNEZtc2Wycf9trWbwyy4LFDHlhNMO4eCrd0qE7IqoAwCS
wxbb+/mhUNXaSXdC5QTCz1w0RAciWXAWYpeCc35THGXL4OnXVflx2rYVNOxIFY9u
mlb0uRCyDl1GVykptpwlpP6/IoZwqGrYy+uKJSGv3qvhxsPFrkKM8ebrhBm1obhb
QhmcWLTA3G1MfmE7LlRNWHB4tKUJWpXsyBQ/TURneSt8jIgK6HAl9hrWQhYEB0TV
6SorAjLs3tOLZ1OW5h7AhvoyweG9gR5fiwrrhr60Il5OsOhdsyjXVcB6WzDqX0Lf
VRWMot9wnMMms/zurWLanljsRH9OLRYkru40QNugw9XpZaULBLqsuZDHdW4mStMf
+NkFiFjrtuY9H7CouJ/B5NiuagRezDbKm3AFtddMBOxfAEyUnwWKqZVUPwNOBi/c
CBAw9xhnl5N4Q1KvHGVvs080pyp5eEA9PnyoPKWGMVz1cEI+pcrfwypEQOhrbBuT
fyE8BpkDUgMMFQ7S0UHZ/zioDRt/yCHQby2Fk6P+yIwLRrXcP20rERvXus4K/xVA
kASbbzWyZKCiCxbib01JWhk41QJ0Olj09eBegog49+coyKkAsOEG73MqScd0Yuyz
utbQkuJr+cTvzxPn6ZoUNKEcZTKyz2FHDsHNabbw6YqLh8MRpPGwI5vo3zrE70sZ
ciBmWMfIlBlLp2DlMDeqcuER8xHmNEB20+TereZxi0BwG+us/MtwwBBCQAvc2NIK
qZyIttah7D6RR0gh63nPUlUP4ReZ9OQRN2iM+xnhafOzp7h1UMtRr6hGZbYCwvDv
RceRJYSj5MUcj0rQdZWhjxX1kVXGw1Cvh/dDHamf6CvkTB916HqsAYnMK68olc+o
YywnOR8sOypPExvIEQ1jRg0Pa4eNFlTHr7DoGLWZlKySR9aTTa2fCTUZSIqT1CAy
smoDxrMTyP7ZPs7szrsqwiur4OhlsB4kBR+iGSzqblSr9rZ8i4AwQl/PgJVFlOhn
1ZpJqVWN84gOzMlcyg9Jz+8LTz9k7LBIEfioRU9t/wrEhe8nt7Xcaoy/Re1EXU6c
Ntv4efLB3Ke3QPbbbTV8X34br8zxfJAB3cB8rS/ZvvdaMTiU4dMSiJ4mNZXp9/SB
qz6p6IJG8orecYkESTKv/m8N6/LxcobxRrIDC6e/cHznAaHOhdDLn2MlI1MmIQkc
rsAh4wrfoU0bLXfol9sKyjdS6pyiqdRoyLB3HH2ItHnAF6Fwsgk833N2boPOMg27
ZCCzqjGMuMEmB5n2ggh77DggcwxJLNUlvFV5/NS5QW1tShIZaUXq4GAjMcvzVsom
ZoiwT1HtTR52LfufFxVrJy36i3IdEdcpuSqA/qwvb5pylzZVJg4BzpN4u29qZQpu
9iC4OfXUF8AUAeNT+9MwLLfkSj1aoHTXGJ1aG2YCjH/BlWfw/oISyg1RawYV5nI1
K/lHAD8mOadRgs9611ds2gulGs50ILtFk9pzVi21241STfQ+BsRDIS4UwtDLPwHZ
y/uuZOGkUwMhPXSbSpa35PHd4PQDGXmgLWaHNCxyISYqlGOxze3My0NLI4tmSa2w
UWGmLA5fkmCMCh6N9ZNMKrCKGbG8Bg99h9U839VbvpQPr+qr+o6z9hPG4vT6XwLs
BeAJNW1H5EpT58M7grfJzx9cUv09a029mOC+wes7c2VtfHVKeqKtkxVwHLIVKDtf
nXkdyBFFZ8e6ZJF7tXrPyf0p3MmuDetbauqSN8MccMMwzeLAxHByPdkSbaEJd19Q
PEIU3iDwfUCIl46pbFd1q8LGCEnFoDhyLQQLBUCme5rfpC/1EEllGUfkiH3zoGhm
DuHjjKPeLswfqC4u/rwPhN9aOMyS5czBgEtr5wgz1Jmyccuv/sULfvlEnTw/cKw7
MAbV5/Yfs+LK+avHS5cilJcmX1aUbDYdMgLO/qRohLcO/J0SAaip7iRMZQPd8Hwi
/h8bC6UnR8yqzb5LBjNW1T+CSw99qCKUrbmkjmSF/nx6ggdw2xteKrfrjZjpQ0O7
OO7E92LUW9HNxwj1rCvdN5E7XxWaQLr98SfXQo/yJnypr8ZsI/LpPGq++czki4j6
Xlcz402rn702dmiReH89A9jHP2o/N3k3gkQrBivtqo/2mvSKgwn+yLlKrlbOlwxJ
ovFAN4cvAwyeNWtB6kr21adRRu8FiP+iN5PfOiJn4Nv2z5rXpXRSuaqz1Lakf6ra
CtPQsUJBSLbo0WOy9Dl3K3myp3B0smBqlYPg9vIr+CFtuDCUkxy7+m+sjIqRNkrs
1Is5U621A44mHXuYmYFPXD6cD3LLLOaub4LpAo/5qaqg59DBfKIl/nBfKaQHPoD7
JYQuG9zZK3FsKTg1Z/gHmrvWZ9lDNfcXcSpAqVDbIlth/IAzF5G2geOuLo1qK3vb
5Q+HE+8eB5r3qbvKc1yi5f8hQPwFktwpBDG+doBiGWwVmgsTlqcoYAHgwmwN1d8C
dLhLVviOpIcgHVd0HX6uNQKn9K5B73PCzsqrU4GaVTC5xPLqu384BRYymLfpmilF
DHI3hTfSbUy+vNH5e+XD+ETdVWOvLPms5h8nbLwTMsxcMBKVnH7N282oqPsqj3qy
QjMlaEVVi6jVR0kKLG1yW/qf3vZk6JdxttJllYE8JGhROnRU3ZNC98QPNR3nyXSo
ggqgRrUjr7Ozt0ojvTAoGvf5hhKNXpZcWrjE8+WuIoRGsG2xG+yOOWTntRT0tdhH
8MPUq5LPsRc9P7eNIclKSeccY1NBleCiDj/bVRS900i0gexwb8XA0CNhtiIk3CtL
Gi6ez2PtPEb9QarE9rGG6oJEhL8OOkI7fuXm4Ub+8NF7sPOAeHLhNkeIMmnBryy2
yqrsD1yO2J5SpPAd5NvklhBuBqnDtV7QjhGS8vr6CzpSaM6Qi6QNcgj7Qc6B/22f
S1k27yZxPJfIdbnI0/nTrLY6QjFOfVzIIRtnpk+HzpH7rqJ/PaR0bLOyUyyRaW+s
I2CTVWMTPFJCV/r0kxEywLGZE0tJlXO6pM/DQYbNoZUNOKNfkbETgsccY/X7uN89
`pragma protect end_protected
