// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:37:00 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
fUe8wsBfgTJyJ1wGkkOm1Z/diUiBTIecZjXW1fglzF3UOgkx2j9QEB/oNmX+VV2U
ZkSu5tQV9gW8Bvv2oJo2YoJq3glHXrpOatZE2jSYD8yKtnnE/FdxbtdmCXR2Zq26
aRj+GPRjNcljD/KgNACiwFuq8k/xQ8ELL5sypk9VZlY=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 18880)
LrdMKxYVBqQECIbz/Qi5U+ouw1Jum9rG+ZgTZk2K5deyQq7/PGzu93R2+c7mpULd
QhnNAvIji33cdXkYQWPgf6llFO4iPSWxbKNY9um/lpKnebSJ2uA7KHLyu/V175pS
1HRUs7ON1DQhwWTLYaI97WfQPXSd63w3yNSo/6lDm3rgLCpWxD6ZxH8Ef2iKQtJd
58GMnCEOg68dbAcxtLXfRV4uuHtlM9xwVdTGnLOPVDHnuV4eXXB1AYFNAsfPgqFs
KgvkkQFwQXTkdMDpviO1hzbaQUvPJk74vvw2/LaBAAoyTtVP8NdqaIwvw27sLJSo
l6mryZV4Sltwm7MVtFrUPUQQ1Hde82aBuSAGN/FQciMxQh15pFpThL7Amqvd9vsE
B51RxYBCjJSuEEVpYunKZxe6LtDCWNfASVjx2PO5u+ij7Yy46a8g1fmyb1bYxZku
htLjLThQjjQg2VqbcCUW+mBQFbT54CR7ReJvBt1Z1oYzBk3vZ60hBxDQ5ccJGy8N
WtpLlyG2qFAnLv0H9nLiUFA0ACnmAouUxRme+iVKWBUmEHYyH0TJmvb11/y6rzo2
7vC2ruMjgK4TeHgH4iJ+tzMmJZs6S3r3lDHOFlx3aQsyW1UOloxLQHglCA45XSTJ
XQ9hQWOH1PV47cgwM1RDkdkijFXH5a1u0SUcDpL776zsHWNn83wyCmPZVv2u4/aR
ns26u/4OB1f+RMcf+ES+cPT1lp+F+eC3x/vqHJAlwU4bvgR1m2gjE6eYW5zxeloR
FgVIWw77ofy8lBOJM7ojORYi3jh3Lss7pvB9DkIpSsodOuysTzSgQQC7teI/PVS7
IqgSdTb4pPO0yek1N0KWr8LyM818t3zUFtfXqU6xK+KwZPh+fnL3uh580vZXZbOu
7y+hWCuOhJJai8NsNFalYPCPsDz30L7FvnabTJbYh5QuAZQMtRGG+IwndidmYY7P
Ia9DvorQPwrDhgE68LAJxisycwe6GuxTNw1p5vzTzp0QxwOUuAtrhmysHtbkJfxt
hZvBg2LrG1TKV9OYic1cUB/v8r2Fstq6gG3shk0p2RclrAJ3v8mq8xx6Om4OrXZA
h++AAMYHQHmWeapKrV9LFEMd/lEj1JptAwjCeDSHGCrex6hSSLjZSyllDpSX5JqB
0I+zLO+6aYmA77Y3ScgY4i7hznQ0F8URRxw6etFLAwh9qWgqd0kbgcTrLW/mZ5sS
CT560cv3sj6MWs0rw169Kujjj+G05ezGMfWB8aaipPqb476zGfZKo7lfSUXmh2Ii
Wfak3QQrez7WhQefdGTdUTrnYHW/Vj7vSnYGOmyMrrAD8jAuVQlhGDn+PUeiKWlh
XhNxQ847gy2IcgtG3NP6tmMxfzW9IFWShdxqtUfWL0d3btO+C3yeQzSvRjdsPOUx
xmZp7kMFhMBVMKxoQqhLAz8kSDNeCzFzDeLdj06pO4OAyqoNTAhVYv83zrLpEGar
S4iJaeNhbLy/5tTlF4V8xGrNOLVgUmYXJwA0UuuzweG1NZMHvdBKbpdKhnqKi4Fn
JfSjQI5R4ttb/eTsXr+U1f5PT+kJ6ZJPwPIn1B0+Pg7KZ/2OZMTGG/rRej6mgjFd
Myu0Iuey5qS4PQa3phXQXgInmSMntZ/n8iAPoBB9LfxBE6ln0w2HgkaQ8TSl4pJb
4ZRdxF3qMOlLh6PQ6drRpqRm4js0kPUSNpn8+jwItNSP4JfptxDxKKCySSGPev3L
creXoW8BA7GB6nMZm/O05CswqXUBIFUwt3NVfAeFWEw6MC+VP7Fglbrfl3/00B30
CMWUPIXgvpDxsqEBence7Gw09imcduJTZ7wFje3EX7Qp66+ScCenozknLT+oP7sj
9J4pk0vFEtga9XOIAKbiDkFO4uz8hWbK6PWSukdf5dzyxPKogHWrijqspbPzy2m3
Zrcc+JGBTXbd89zsGbBxMsVwsPOqlP0NuLuYvtYsBDxLLxHjfIAegldi41yBoJpr
+md6FODJMvVB5bpUa1EGI9ubyENlx7tX+BPFhfTv4GgzRseUBRsRMmByv577ArlU
yZJvDkApDykXhybJ00CB7abFPoN7O13cy0us5vAkH/BlTbjuNeaIRHZBM33SGJbe
aVoapNaZJHn499SfPF7p/+Ht7g8Tl5tAwY9fUNhze2dSFJqQcRs3PDj8dFRvzwiK
rlY352F1QbK/wi28vvVz+9aBVYIjTsS59tRAhm3rfXlLR1V5UvAEMtR+sgmo2440
PgR21mec/I8zYZbaa0aOkvuxEGKbg93fRbpRbrvezNW/ppOGCA7Mm0DJnIbRJeUo
s8GrL9gzB7N/Habco1mdeGq9VGItibvHOCf3nW48K5vMQrx5iTHkBFhttMmgJd9t
cWvZmUqMT0QOIWMbm7uORzyNH59DS0U05vl7mGWJoFjdCZwG4Xc1+yTk+TJd7k+Q
813PsnziEEdehNPutQCe6eXNtACk+ctLtcsjoC7HO01AQJhTtxNHSmt1xettul2K
HrZCdVQmw0mt/Z2uVGiuEXpDOjYw6HD3EWxJkBjysIXMkOCqsdWuSdwkoISw40lw
JUvbfnlB+T3uMG4ZsU7wy9nMIc4okLrBbh4fv8yqHBf2tW1olsUXQv3gF1TEl/nE
C+ltTBOBzLEO/0Qz4CIPxYLL/fyCT7F0dZv+fHc70wKnBJM9palajMETocni17e1
Lwev2uVMcCqX1+NN+6DfdmZMIbTkyxMUjpeE5yiHd80YDX4xLwsiKA3E/4CUBMuX
PAq9SE9ou9nofQSYADtdhTGFBjIts+S9GXe+VgvMwU8N2Zq1aYHMik4TXlNlkAD+
Z76LFquuwSH+vTKLl8GhhxDoTXGD7qahkSPeva/GIoOYqJ7i7SgX7rzll82pFAnl
ArQapMDfvZ2zf2kTLM/Tl2X2hXy0RT8mMjlQkganxg1vykTdsZnkxdkOrabK6WE4
0rayUlkHlK/eE9kB2H5mkKu3bG5V1Rki41d6zi3+OfHBpNF7L7qBQiM6skk8ivQ+
TIa0Iwfk1hw0zkCuGRRW5D5nWawzuDg3u3wxCE83ajYk2AMg8LX++sfS2tYQSJjA
eZCDZC4jJHEF82XryVjjAm7MisIuihsxAAS1QwosTsiN3xaVuwkZPzNSGHQtFQqf
UTaQhELX3rT/7KBjNbXCKHbp5MnpYIN6KJNxlFr4vFSMexruQdE2mB+i087ajacl
03os/MbdvcmwEV2nkDm0WzMqy/Duln/DVRrGxJOAt+sHWeE5z2CLCD7LYpZsBFaK
vja3SZAWQC1kKAj4Oy8mpXARyUgnGFQT8h6kPRijrFahIPSdNK0sZKeuW1yjP/DP
GBO5/EhTvtOZGep8w/718rVUixJvd9Gl/h245X43W5sgVSPpYed8b0tibgKrPlkN
WsQLjV/LfaOhrzwhYg/7yMpOPe9cUfPpQbRDdkEKokbT4YyDIkMyeFTEqHc4d9lI
pRgrNUFOZHKBprphbydp67FgAPkqLVdJvFTo7JGZJALPe6H04kc3i+ru7r4/anAY
Xw2SyHv+xCXnD6DQOQtuRxGspJ6GWvFtNrpiJ/WPKRdnLf2no5IeNnfdupwyeD+3
z6LD+Tul5tYIFXR1dORZ9AP6nRsvL/8vpfHiJBu3Eg11Q8hnwWSliWnA0i+YCt2Q
cFUMRiRlx8+T+eMlF1EAJUq5k6tO8QG51m1O3/uF6z1V863whlgpMvSqcMs5+LVI
fvIvPWLW2WVssRhTJtp+ESjSNfLjCUFcdRrvos2YX83aWZBZNFHhmgqvZPxIFgJ+
S+QNCesonTMrbqnN6B6UkbH8zB7sTOg/3bNCnDGgruRgv8cydvUbN0j3YaaiVerJ
tku1IXVS9SphB9C5aoQhwxAL+yMDaSPFYrWQmCtI8dfphPpu5qN5q1w+TFl7tG/o
lKm2pnypXbs5TMryx1B2OqLk1ZHJyHr2dhL/jl0KSIhHI2wrCvVDv+4FvGUs2ev0
ZpFv83GjqvdxMXIktsJwVl9T8PigB4dqmXhFV0mit2pBx/2reONy5RExReyDXgiu
rlbjhtD0rjt2SvrlJ0I6wmx5YSnMbHJ1V8kgOrGwtozmHGPQq5o8zQrTtg+KRwl2
LHsTkt+XfBasJStdO0bwx4S66kCWFC05Yw9oSao0Xti9Xp+X6eKP5FmfkOJyNAiQ
yM1eSLUDZOt2RfGdl4ZCDjAtdbPgA0nWmE+TndrYfKgPJpM2moZrFfXrEGXaVIf+
FTEPPFYRvLnDCGRC1QH5+PMA/0kyEqibUkZ4xDD7yLBudeHUrrEVciqpbrKQYZRn
8pODudyXKhwV7HAyf7Y+8eH4E75b/9xfMTya4iJ13wbgQto+r3Pe91QUdjkG88oK
0DdtEW+iJbAgttJ5y1WjNVHyWzWed1STO+JQjDvVg9vCz5dgosnKMc2nxsNMd2d4
9xQMRqgLJ4km4ZZ563L8AT9LMICIgB+lZxmSHZBFzpgz//ctQ6IveqKkiIaXeJJH
su5m9LgEXYpP+7PDS2voLSX/K9zbPAZsY2wzAqnjDgm1QrPSKcyYIZAsNejF19Xk
2M2piXUKDLLAy6ibbSUswhcJPwSS3QIS/Drc7tVXI0tYjhNH+b0b1u4fmf5toHg/
K8jQiTwbVC/qpJGykJQOpQY6CqrYdifApb7e4eo78fKLINBocXEovaBRPCBKAIWa
T+5k+vNdDOXh1e2yPW9ERl+qcEQ7V+J64q6fiHBbqnAuuNA2RnCsMW5EPYvNxgUm
BeBJPoAWGhztM0Ayj7Xjv4FMpxlRjF0ev0KGhT+iFZE2BQb6k+uncjdVmaoR+Ptg
wWPE4Iit0i04bXTUS1J5UjDwSkcbdiExiOWMHhCUhSzFdHAydVpPgGz7RdNjebdg
IH8d5g0gq2cNvdEKzFQlembHNUodk60DPs7WHuLTr81RBQW285trHPhUFnNE7DBt
dLggPwQcRH7hyqPTCVHZlbRyjL0QJ/E8DJTQkEGWeDO7wREl9bshRV4opgzPY2FZ
tpWgoWkN/F3MkuW/ymHgqX4CHnho23KCnQ5mIobn1GQ84J17ejFOkU4I8SblhJOT
9xn3qHREEc6rXX3rvJIx5IL/34o/qH7EeeVWfc04Z9pbMOy/4ZmBxaGbQ9LsYHc8
apVXlcXuzkck43FpVU+VaExSP+Y/vphYxJIKUttClo3Nb1NX3sUapkSY1cx2Quo/
RNNdc4OGCe6YKS6tNwWBPN6FcucCgV7FNnKU8BddKKRThDAybQ5kB1XKY/ld8Bz2
ktZIjAIaodXTRBz/Xb1SzOyL8bZRgrvw8hevixL2v8qE0bLu8Ef+1IMk3o2Cc+y4
TjWL83tS2zgua2UgTc9A0p3Bblyi4Uau1zdQLQfjn2Tl+JaSqaZG++U9WppXsOXU
PLufw7bmWPL+TUfCbXQK7uNPpS5ym7V3hSTthgCer6ZiJw36xaBjdAQt4Lu8BJJ8
+12HLbV3S1XxkCWhApQZr0VS/v2rI1bh5i4bQRiUy48YVz4Nr6jl6F8DAhGNU/cC
LZY8b5A8y8MQRzQGN2wCXifrDyDHeQU/NBolzk5gzuUr4N36RhHsJDTvNCZELSQT
MinwBk2luQ4gxYZ56VbpjGA3RlpChRC8D5Kc2uId+pzDWB4uUk6Lh4UflKquB5vL
FgsWU+riSxGUzIKbXVmdRmTf9Kbv35Rq47IplKugRaYXtEI4AM1HOqaP1xWWcq+R
/Wd7MKRfqeKFKxvIPNQgRiPc/QSeDx5DC1ZDoeATrcPCKDSaCRRP7Lze850VpmHL
OkSC9M9SW+mTOzVLvPFM9L3IkqZPFxl2U+wK/sib+jk09hj8QsYRfzKfRTzH4ORQ
wvBahPRcn6Y0QT3Z6X9ohJR1TBeFv37zys9LrZYBZDLtS4v0GUmoDvCDjCP3n1rM
wf2kEMJeE2OvJuf16cC50RFlbDWRvLl3mEyd5v4blDNccgcXAQrGyncjbjbjL1rA
C7RduNTY0Dbb0BU6a1DVIHZ4cZfBs8rrOYmUqLNrJA1XDKaHSwnwOOIoPGJ1q8EO
n6Qt7QKK9RJ1tJhdI394I7lM1skMr9R7mE/93jcJT24MtQRsWSZcHg+jGqsz8aqD
kuaP8NBns4gt/BTmh5mhqmnwRUMfJNMZ53BEbEN4075J8ghALo57uEtf12ZntaUN
YMDEg4phLRzkjw6ZKQYAlljdzwWPZ/gIg6oxj2rhSuvAi4qxDbnmqJ+LRunYOhfd
oTn0Zt1yXOdil+OXdptubylOQJY76JAGUp0354LMXDSwLzATtU6AxmFsCZajoMBj
r2tIaSjHH9LJX4jraI6qPvb/JnaSm4mCd+5bDafMwaoWb9FAn893dK3cm73Q4DMF
lOCvKk9Ltk7ohWHUt0e52Z5lgrVjfo4cKqdIVWJVwkzOM0kZ/hPgqGo6DWhwjDnm
hBVPRGi3xh//IwBTUwJUndWv1MiNKPg7zwRxwXV+i1/kzUm1O+AwGepPVMVnHOXF
VcCaJTNAl+gr6KQqOnEysdXk0qtSz9NSyuFNnThMO8AMXmYVNsHypIMpqC0mz2ZW
NTE0XNsmWn8Y3z/OnJs1g/h35FdUNI61w4BoLQPhz1C9xmguorIEwqnQ7cW8giav
XCnSLVBMqI5nUD2B8JDKzCMnUmcX8nGDMbNTn5aqgig30WqREKVdobsNvJ//J+Hd
ptHAUd7F9eSNiLlppkKUsLfWmr/3wOZRP82AavJNNMjmkiJpR8BsBKEy8q0iPQjt
V3h67P2c9VW8nX3ugEGOEzTb/xOSe2i98Rluv19qWnVp41zri/EJow1U3tgd24kg
P3N0BGdhda45olKblj955sQ4q/2ERELIhodPv2hDqT97hlHu9xSzftegUkHMKbAz
W+NIdR02tLBwrjKdJSe3hBkSdBlMhTRnJGRocD+GOpnUDBec8IyNB30SWc++dtAf
djsgDg6NNY3VylWOoTzeDumg6sEwqnBmzpseLrLXyaWhMHqMiOGnHzoMh8d0ZL/k
OHmyRvWzEWWluHiS5HTmW8k/KXbnVBSA6rhLrhwIgaqF0A6BFGOr6dmpEJRvc9dc
ylKm1DvV/s1Nm0N0qpkscfYMerCtgS4cJs5IxEV6lPRM0/2ld4hghv0FotCRzMHV
5VTFOLShICCNZCSyCn9gAU+d7W5u5CDk0mAwZ0m/fEmrkqZWtcIUeGQSM5RnZjAd
h2rroE51KK8XPzr6C6tyJ79f8zqq+341bCHHFaDW0efHj5n8x+eCiw+Mk0BBL6uN
oX4uPl9I/6EXA2Q6CwIrUJbpC9oq2jhPv4TT85S+Ne8Xp2utehheEtJPVLak9o9m
XJ9hewp3r0tqqX/+H9ryDcN7rW5HxXCtOMIWyomvgBvBhiLT9d2haeWVVEtnb07x
doDr2LV22nnxMmPyl/bm01w2kQfF7gKAd2jWLsyKnv1PyFqXtbDE8Tq+E9elPY39
O30PwwtzmXPus8ZjMljVVhcA4fzLD/lGO/1FXYJgg9Gi7Hx1Rt2snBADdPv8fn1+
aZdhnrjfcmfCm/xD2cKuu647FTvCNW0zfrD5IX/d0+AypIvsYxEmGJEIDbkebm5S
YPBUYU12xBCBTQmm4iOHTI+/rZOIcUg+eQVXkg30KaOFr695XBrFg5d17aULj41c
PrhtyIwr6pZI2Pb6+1DV7jwBUMdLlDblIAjLt2d6aV0sAIjFP7/m2/L0653N8vRk
RzLmIBzZS5F9B8YkShh+dteaHL6xw7Q8/Wx+9HTnqkyrEWuohMLGs7Ae3ogniAD+
68yzZUagxPTkoDLCYGEyGTHjFybARMalffpZB/Jy+4jIVIUHuO9n1l0fM8x+Anm5
4jSVNTwAar6xDVVE9+i66FdjUy5EgPlxjLA7mOMtUSLtDyy+XLBye/9hBBUPQ6N1
Gw+aXtxl/anq7q4kHIHt3gY2NtB9vGwfb5obC4SnhULQmQllPd3tkF1I67xmvcMa
o72O/iorcM0meP6an+OjS0Pp7ggeY+18olVgT8u064iEXwtB3OKfUknk/V5ec3jo
i30Rm8iRUwpsmumNxJzQv/FW5JScDjyQEj2/2Myd680fa0kiFGdB7kLhuOl4G5Z6
nhTsa+bzR+EScB1bIYouPixTX/haLyDxEFaEbZV9xvlAOU6RlKdC3XfSTqzJYfIn
vQY60tzheUAwkABpxNofB9FbqeW//DR+G/RF4iaCLed0UJxC38j3K9RGaT9qoVYl
o06NfNe02g0hoq0pHPC9ZKx8iLULAJl0IuseQS+XrsPNwiY1r4uZstyuT2YtzXuY
2yGyg1mZIgvM+6Qr/Yq3yEPSmZFKLViro7vnhTj011GOGokb36dJC1GXc2jSkWri
bQxAwbEwaCh/7R/r+MmmjVpvcZlpevqklFE7c+noBEsiYFHV0aW/hOgSYrac4T+M
OkuA0nGVdmlyYB9EevPlPw++xMYyjW4LTA8g2DQkG4c/xn5HYU5UKR1h6TYNJBfk
vZzK9qdIGapm2EXXqxGUOeSHXdNXI0u7jAWGlcIniZoW0M+GGN9TtyQ5shRGm7+r
t1YTqmTIrfsW+wM+mbX0wqPHYLSgyR51dG4rUfQ/uhAUwVSEilW24/1RrxfxPfGd
/iCh2WQvM37KZvuJiu1loDaqKPlTaaO+WncvUHFzMYAJjXpSia0qkafQTdOhp4gz
2zTxVsinMKRBpMjMxKdAE2CwXN9OuIcF601TeIldQrVkf9hdQ2rX+Neec0bj7e0k
AXytFErLJ0Cx2LLTHXc/xy8yeAJZr7qaR8VR/xASeyi5n3EBbg906/3MTehqf3hz
5tDNhymH8YyOl2iomE4asLA9BHSrCvKhNwSQz+WTrAc3dG3GaY9uj+nckGPF72BY
1w6YlNPY9O1yaSJgHpkn3xzsYMthfmzNb06W0/6f2n2l/EcYqTNIvpNUS3lL5fID
lwzEH/gbV+N537mYzMqF8dl1YZcpPBb+QdyMN32UcCctfSiVsGUwL4XwKQ2C0UBE
lzgb1fF8kv21ysmbGv+PFfLWVS6QEwnJ+CY5Iats388fYv4Q9AYGGuG54jRGTnbx
PJKoGgAtt2n8dqxmF8qeT6x8iI3dQI6iiFu3TF3SH+eG9b/1QJ/hLsKlFWW6WMbf
eRK91spFgF4UArG9mE1U4ZA7Qhrn4DvzObAgg881XY3iWVcwiVt2m/9En/a0LHeE
jqQvdYJHfOxsozF8NTgkNm/huEFhs5ZNl1jGAgPMy06M8BnInQliRbnxIC7BAYn1
XRGuPBXGq4wh/CLV/5jxuKdkMpP4ohJXnVuTk3Nx6Ai89eGui2RieRyxYz7Ki1D3
jFulJwLNs/5B1et0nBWORX68clmj5okyokHMrn9SnTT3+HHcs3tqcB2b0F/OUAsk
sKWhIgtg3iU//KnRFHOfarjACH9caZl93MHv0yyCqfkE4toU14p+caFyFvhspjB7
5/AXqQh2YQA7z8dVhEoVAM4uU6L/2KzFXetMu/78ZXvikfKyRLvFgz1/kHr1ehUX
GtO8guVImT4bwPHqLCcRMWZzDNBW8IRnkd1qhl7PIBc9pcaJf37UbUQ80UENSH6c
aPoCaP0Luiot2sSv+fPxWEUTOHZAK0jrHgWGfx6Dt2VnGdGhShT1OoRjVO994JMe
yRlWoB3vqbTuEr+1RAvALXDubASUaGpNp0osTzraujrhu0Ya6fcT154Fe+mTP269
xVC8B4owZ+cEmflo43vCIhWUaiNYLHoEKr5nPo/ZP/6DA8PrRujMskLC498Ea9C/
kERXAApQVy8cVDlFbJQltlPw33qK+/jeh+d3aYEGg75mH7YQdqA5ea343ZzN6nrw
uj1vim8Nia52wTDl9kkOBNGFr19pE5HvgKF0WA6NDpJ1eeSmxVAQRl+duupXaOWd
dXPBSJ89ckTVt2JQLul9QyREowRl+ShoWGK/vHXWgB+6rjBX+WgfN7bvCbifeHsV
7Lnu4qj8prDwLLW/xxxnqbph8A1/anjP/R7CxZtQhkzq5orOgmx5GshZGkeVud1h
5HgOIMMSLCl7Mr/EROwnA7XK2RL5pV6ZS0DNHPk7pvNXhYIW2WgdItkplxPCvbfT
GogqlS+w6o5HpcAK0PRSRdChYR/zqA1E2I52q3Nxql0jzAdgKWP6txfz65wxP4/x
t7MR1EPySBa6z9xJG5FDriZIz8hfIrH1GvAaSAL0ESTwlLQAvDOaf0EHTa7kgwUm
0HnUdkFuQ4dEe4TFyinpq328cWO7Ll+YXk6j1LWV1YkwYp4Z/9znDaUn0s4zH2rV
dSzKcgE2ZAShSkHdpJvTHbVgzuHtqrU0hH5Tc+TurWRdo61xs4T5n+Y7qZd3a59A
irJrLDbgQ2Wi/4uKsMVgymxWefIWAubxBhJA309uVWOT/7i9D5eIgbJzTZJJ9iP9
2vxmBx7Xy+oP4CaUItqHF0SWdG+Bv0Rz+WLuVrg20fqPdZUA+QDFNA9k+4JSrt6D
ouq9E8OtDgEOErh106EDtjHJqv87sEuIeFoeuwcrpz7KyuxYbpy6X73VnXLbpjiK
Lj/8xZvGZqaZei3u1Bq2LlV9lSjNPsvxzE7cl+LAysgn4Tfp+UwQTfxwrFL7dOhx
TcFQgFI6g9fgOaEkIZ8ud3XRV44v5tX0D1+4+c748QXS2qub6hhn3n56fGWTqV3c
0psixUsHSh352V3cw2mI2P2alSZRW1CBeWMOBvzH3v5911OtE1LPcpo6/Slmw8YR
SRh9N1IbeG7+T4ufaiyzePNjqSHU5bLHlR/S/HGU4/MrzsyW2CImUURnf2V+pFJe
NLzzlJCcYzlsyLOOZS8u4lGU8XRUDd1VJC4Aft/U7DVLSNMVscXUy3NFdwCGN7jK
uDTCZVf2ijM0HwCu8hI/rl0VQ6WT4tpBvkiHRvquLXnBEjFnM4WmCTJmI8nozzsJ
popRhQf84K4/eNIWWLOKIoXbYG48KLE1j7LMQysEP0fdcB7IxoWVI6jGMKbooTI9
xsoLKjBX7KiTBFy/UQnmbyzZIK5pkvTVwxRMuT5UNdr3V8WINlaSji9cOmZ632pD
bGuBIzHe8pjNDTbGEOPzy3An20LyNcDKR9gTlseenQfJjuru4l4BwyJmP3ZdU0Qu
H1i6MOlY3Zhvh04DXSLOo0h6DjYmuVr4+XA0zy9s4CZBu4/FQKdzXoo7SlpYTjIh
1/FI6q0QQUxVcaB8ZoWHNlcGucrCxkNX3sIypSPJyvSji04VmQ4iqxkTaZQxLAit
zxT5tSkToDwlgQwkPbV7ZOpjjev4OtsvRpdG9NBNT48/mkLt80q/a9v7lduAp76f
gasnICB+9L0GTKlbxqT6WBrB/wQNedGNdn9NHcSSpRkSozq24Ri5bpteK/+NKhoG
k2FJFlvBkbkeiL8e2ajNOsVxq7k43uFuBro+IdZPPFrZp5HL74PES5KPSqoPvzyu
KuSIvGR0r3VP0kEvhc4bOIKL+orCUwSguxfpgdOrBp44dGNayunw4TmwWbSD3vQt
1aYa+B2Y6sP8Sl/3+v7tiV83OJ6aeV5KC92y24u/xqvxypuZM7jdvQUbIJp3tUCk
FlblG0aRu/yo0Ui0G7z2KFQejC5TTqsKoNsIT7FBmI8j3wt2aLUn4SULQ2WuZ5WF
vf3/OqB55aGZeF+beFOKfVu/cvoFkkq3rzndsOGRIwcgN3Ed78iZUkwSPn/jSAeA
qSIk+U6nMs3Kze2gD94rxeLU/7cH+8Vc0Xsjhx3Iq30ADd4H0mmmvWJ8YffqYSJn
rhnoihujRS1aVj3D3qy84mVWx4eQii7Ic0tEqwefxbDKA1NvslTTE4k1U+Vind++
cF8Pi+eUmtMkzeJS9y+wFgj9nUtX1MncvEEw3tlJBhiIdyqzRFXrGKYTQKs+gWYI
DMcS49MjsO0xLG6aglNtTvSepX0jjsN511rhimZDX/6YQo6lfFnTYGI5aUivVMMG
knOg/eyshySvvXHO6MXhJi9Dw+0vNLIQQ03XsYBfDTma+1Dldx42Q9gLXLHfsXCC
ruKinWTfPgr0t9NbFRJNv56vA2LjKgdEqHm+WYkAxiZr6InXDwlSHhztoiCsODTW
t716YtRATbLzMdebRqzMPu/IC24JDNoAzMT9NBT+KU2tr85sYSmeCvohLH6xCBL2
5yOPOemro2soTV9CBHyfUmqGhSc5whwedbGTbj9xAqNqO5y3zYX5XVRDvUG7NSvQ
7jDEn6Bj92BXbFNj7pN8ra7nvNNWO9xZnwkVn31uYA3z3xv6CGjfwZuKUV+4p0rC
ImVyJzHwICfuyTzkzTC4L3Hzr5F1HzcmudaKOJd0rC+JmBeLOGZPXIsAPWB2/CCW
Jiqdf2E7LVAR1DgfLF440Z9lobY4evZzzE/TIkd45hgW325sHYbU8CMJc9kqRhps
ol8ytZNcww60QWJud9ZVBCK0e1QnAHfbdBOuAUmQw9Opl84S2unLj8INM8ykskyZ
4BNfgjNCpy7JV3T2RWWXU3AijkbDt+M95L0aeRGwUFcoFVF3ulDRL9Ioo3AWmcL6
hGYPR6v7ylYvfSILCSSiboGVVUO0XcX4Q/tXgZuSpHQNt018h3TYsC8JLKvTfz9a
I/a2Px5zQm0uQ6XLnQHoD949SnizmfJ2nSxOqIVIVzdPf81klMUKkYCIWlrPaneg
wb1Cpv/yDOoeGOrJv956f09XC4VMpd9j6hPeL/hcz69GoRe5VuWQ55+JLB+zC++b
w7V+QJrdFzNZbX9K4yiWtJcYHa/jXpgBN0hSOANl4zlq7+hkWdh38HvJIOYmBm8M
tClT3zX+BfXeY7zbxCZk8Z3z8ZyzeNQrutPuBaour8g32BOb1gHhNU4fpZjKWjsj
bEtKAmzv/wYB4XAT14O2TU+fV7t5NACGTRhgao+W7Tp8Y6COGkZ8NG8tabERAMDS
9JP/8O+njJiaIii0onegRGb4Qjbh5SQD/P+Tf4VBrr7WTzF2Bv+ZM0dt4j1Sq+B1
ZKWCW5l4a2RHoHAhi9JaKb0ijAoKQNQAemje/nHu9cxOtE7PFNBj4KjriUC4PynH
NPTrUxw2ZSTpriOSC4IUDeQHmLrOw5TItnBfToEkzWf4K/ZUm8Sm2ub+hoFgPIkc
yXJJTutB8MXv4+gyKAhrMTr1vUEexIkU68xxmI0eNc+NznY0jL2E9yujg+mK0pXv
kaohsSx5KsnA4OlsOHgSM/Hb1l/Y1mmn4IunQlmcAXZ1z5Ecfd891NuXBFN3jpmY
4h90Dy1rozjXb+16m0jbxUWD+N+5Cm4yhd0wfXW2GLJW3q2+KbJEcIUvIuT9dtrB
FddgW3CcQOx71l7W0I/W6tit6uKNc3+HHauDyGUtDwnjNakvZ3nAOldrCk8cdnLx
m1zALd4vKrLMeBX0HsKTay4EI3kgU3bkRrhnDyqbschbVXrqVIJerPuRzLmyp/c7
u7gLLOutGhmJlmeLHzLS6UhdDq80fhNEbh+EP3KkeqAzHvfXurfB+exTiWN9uyve
VYf7dqdfRFQLgQ4Cj1D+vYjtoj8nG9+x7pdd6Gc/Wvtmkwk0DYwALTNf2925AfjS
Dhwbl2gPgEOS3tr8lMMpWfxD/M18+7oQVm1FHAeqbRpL9K2i/8D9O7NN1474yt6E
5Yfu6xRFUFtl48gkLn+lC/XMmXXIFwAX486O2B+88WRVl2gYeBng7BQpS7nPycjj
2ygqYgmYrzubszCqlTHokIDYgH70ArsDFsfjA+t1+NXELzfn8dkU3SGNfuwI3PHo
1WxlFIrOAggOMAEnAUzTvBt/1tVuDjUVL/wroQ6ejXV30/SMc6aMyC6nwXTTQVxO
txP3r2pOTZaRdIdX/dPzswuP5DhX0I5f5SIETmF79zOW/Bd5YXR1m5vtqbC51u8c
rvm/4tOlF00Ku1bix8lBs8UAgGRN4UANwMpFoie8svIAk1TnXPtVLGIZiB9F/bhG
We3z/sD1pKgC3AYJUJb58Z9x0XlmxEPlNzCHtq7+wNX9yeyhyFDXamoa6VNPXmKJ
wDd9FqomBYbvosqt/w3deKBZwMVw3rY+6J1Wjmpdxqo5z2+eLJeL+fOLD+b6MQ3d
uUm+cShn2ARTLQROCRge4nghlOjT8YLQGyXzAh9cSJ4Ac3M3Xddac1I1u25qJZ8R
5pRTvz4ubZfb9rXd2z9VlQF6z+dYF/UHQ773xwrWPc94A1bSt6M0HShkdMIVj9Id
cNLQD52634DKvpQ4Wd2k/x08YSsVMutiVdgktR4M01lPtcNPTpRol0sCGsP2//eU
8+yd8cS/3/fVnbq2/0YGmL5a89TX4EkE+CHNi2wgMQhuqlxNtc6r2MAg5HSkylkb
36LDOxbTf/hZkKZA80dPjEQU8Z69QQp7nB3QistHIf1vfxBQjRQYzQJ4l/9VnKCw
mzPSAoEPLi4pU7cr1SNxO1MWuhRM1WkPex6WWyeqxWbI4h5JpU3HREJYM4PN6t64
fr+pc2p/7hgaj+1/5yAJpHuMSLkklmbm+QEZ12HxKNk6Ra3uvbsJdCzEO74GTseb
W9q9EllcAo5y1C8J7u534bYM+EpRnyKeWz6NhFkBg1HCYpon9wHSSBsroBp4EM1e
Aq2D+WEtjxZI4/KS28whgFV8rXrM3ZFPuXIAM/XnYOj2aaB6xHwi8d7EHUREfCTM
otveUYiOAJsfrAeOr8YuUgRwXFk/87D6JOJ09tVxB80Ihn3T20hw6gN3NrXDOFCs
AIK5B//OJ3QAdZZTcHWlbhWv9n5AWQozO1+BHrrxyrdpc7YIQ89d6pm8mc5Wyx0a
kbUIJs6Hri9d7g3NDx7+IrGzxRMS5hJ8x9oqK+bo/3Stw3l2VTyvtWoqyq2hCrz7
ujlqLL6L8ZVuWriid/DuiHs4gGj8y/V9gtFZb6fgaI4JPlOzaPq71JnvTn9UDr3b
TRtehRvUVSFiJJU0r3hxQTy0ED/Hmc6pK8jFv/wNFc7vJEdPfN7J/F2YSYr1OWXd
Ezp0Ip/mlq9pNfYY9ZikEk/G8HD4dShsgK0vXKRc42yeNMVvFs8hIi8hTDQQV8QR
zoUWbLaw89kdrnlVQUf80RvadpGCZejPaXtNkLVfIflg7Q5I/MnAP1MxUmrTNd7M
i703IV1roSwjSg7gAy5qoKaYo5eaPdNiCG2y+10cdvSx9P5ujPuE70fY4Sa9lCf/
dQiNqs75URY/joUi8f1TAF2X8MGrSTdHdf9K2cu2SFZFZq38eRzdWsxyCnN9nlmk
OtZ8BqQzDoOD+vpcsuJ+cvs2TQZaYqKHyInyJi7wi80yltIPbydTHv26TgGsGI8C
fmTJdKhS31wXzr6jRyvvSfpbGtQPsgpbtEvxdtFOONxMrBTFjZ4vNCM17aJR63GD
HOJiFPsf59ddzpuZdMSCuX9Q3lclPeB3dpsjpeRPAet0CdD8sVUj9q76q5JRqqFz
njHXD6EKhY054wnfyGgNygn2IERRFR1w1kxWx6ejCPODrN/uq0CGMT+cyCIM3NZy
sLGPO35CPE2S+9g5h9iUH/g63uwkNt+5SiAVFCI7Uvn8smGXAoBYdjV1d15V2lQs
SCxEI4Vey5rKD/kE8sWx9dn1BTGKlqhnTt3XhXkaNfHAR6OUZMKrLjkZI2OFo1mK
3SnC5+xZnZI8o8wPaUZvMxbp7wzEBsrkxzGCVlboBbiIqwO1APirnK4Z9cnnZrwH
TMB1OqW00sNJjxq31O0LzWJ2V6mJCk5gQU6IOjPbg3LcRRwOgmw6YWY903jDSw0I
CZpp0BxpS4/K50jw79/NRZtKz9T92rLirXvkHRhp6HL+/ulZGkGNyjnMhZzVRbvE
VtxsVWKYmP9+ytNxgzYITQ2SVPy2qhORPWFnWNgRwAh1lS7M4FnLhBRAuJ7ZKEoC
JMXYj0xU1v2QMa+5OhAzZaofBzKzptEsI9KSaFGd9m7YR1skD5v3MhU8UMLv2w6g
SMAey9y9nb05BLUldsu+9G+unSO0zqRinOE1dKM3wcTGBWRjJeR8im4f86Qz8GY0
3UFLum/3V3yls/QULUKO8YBQ+fASX+zEHTVF/lBRdJk5RG0GdbYUWhWRTW3XfF5J
Of6lbRwvH8qCMReRwzG9xndpTTby15HDVBadVilA86sc6d2QtF8khp+gJnMkpSsz
yiG9y32Hf9D6SoclB0Qp+sdrXQms2oAjUEFl4wsSQ4qju4eVtbpG0nUkqNlVwzPb
hKSZibmyCrdXGcgdBd15dE4WFk0DDc4k+Oia5prKCrsdtJbJ9o9qe54DU86jCSVF
Vluzikbg1o/4nDl0fbqYY6ZMraugYvpX0y/BLDMs8Od75fZv2+rZuLDhXmGLxya9
RWzwRExy5w/VJY9VYal2P9jRN6dxYjMyGxJw68wiNmud/tyqGc6S3/1H0p8fyZMG
BEvZ7ap19AbAMJPwj5Xw5zdDmZNT7iyME8aoi6jF2hGsuTvayEYGrikBKNZPcuGt
hKje+w3KugGp5HgDNt3g58OMaCA04ok/A8vnkbv6XW6RHKp/y1z5foACfU2rUb2L
9oDozf+41zhXq8/JwQNfAU8D3LClP9CR19aVeDuK8AdpWHeQYzyWGBzfLlqGDr0l
USIb/gsGINTvuaKEYRpeuRoCGg4zKVWr4DLF00RMA97ox8U3x/VMUueF93dMYN54
0piNo2dEqFRCi4fefVPrcfeUYx+j33X3DfmQc6Zx3vaGfwNpewYAejBgXEcU0x28
klbZAX8V5CAD712YXSv6klOEWKJ0/tnvprA8HmNHHvfvEVTMHLig+5LYfNneUnlh
Pv8LmMx3y23hY1S9ocv6zF3yBtRamBmTsWupfBrUxXqzw16OR1axUl4KOnwV7CQ+
xRLjBcB3z3KEytTI7p5EJ3ZEzrSuOFltqnTbFiKUZI8bDLISKnDpNUVZOiOmj2wn
Nd4uFg6HcfMht5uZLDQqs62WAkySqmVzCOs9HnnfThcAEm7QRvQzJY2IFqwJhCxD
q1wd1cj+X/wT7O3AN/Vy04KQpBhf7JmJvtf1xm03P4WNtntpv1Igo/gmVnY0KbCt
he67tngJEW8mJcWhMBZm83F7uQPBlt5g8j+OhrM+Pqy4Zb1LaIZNca3/5aWK6aYo
J6t8oPRys9VovHopv7cFyldQrIVpIiOMs3wGUcexqa3NZO7OQ3QjttWiPvVj3ZsQ
/N3BS0MWiVK1pGMpowdiCGVjgMwQC2efj+06WBrfpzjhiHbbLZG7MAllfIyzbqq3
mF9R/O+1vXLLrEP1gKTDFds2zZdIR7Jko+C1dahbwk8xMupX3TexRg0Ydus4mXBT
ha+wUbS/7kTLeaWfJxDanrqBCYgBMo6e73LQuH/M7vNB3e7FbLn6pdLrFJvH//XU
88yXD9Mp2eHdOPGa3FN5Biowm6jtBL2JHUuEPK9i6SmLRdL2SsdxBMHxQLoAvBU8
cTUQ77948JTG5A1PMuCKyvMwijuP7bhjWAqbe79RAeFZh0NWTTAzrF+FJNNJX5R3
pJ8NafFfhiKP5RCCNX0rpzm0+vrWfJR2hqkHTkADsOf4RobmHE7shx1at9beLijQ
9m4v8s5OPEc8PVn56ArDqmRPTrC2pPHypvaKE4iPDT7gnm+A92BuDu2nHTYOZ/sg
6xOsrzeQnsL91aTp/gldhrWpa8CHJBoGHHcK1cuX42D72j7ZdFv+BvC8XlXoxxDZ
M0s+tyPH3wGGSrASP7zsZVOks+784djSDDcRK8sPWGdCvZKn6dzzV0OYaCktWEgJ
TUEgFIrn/UCVzXxUUMGvbb0pnp8ca9OPN+SnXs58mzGG8Rk5BMMP3KjAjAZv88we
ZfKDjrR/Qx/EU50Nua8VjErkZr5IryOMNRo6eRLEsZChYqxlBwFuzULUOSkqXtIv
Vn2gPvyz8+kdS5dM6chPXDsawKES2qJ5l2tr8bOGEHqSkdaFHdi73cjOzIifKb/d
+ZH5B0Lb8lyOAkD7KU928pIIWhPeAvVrAM4JDff7bQBGnv5gyb8ByDG7FpDD52Xm
eL0KYDzE0H3zmC1rw7a9q9E2ks7HPx/kY3TykDspLF7pBHuJ2FBkjzatGL0wMkv1
E17qxNavtH/ywHlpgluunjNDgJCjiW4Mrg5p3NsAAwrp+uwxr5SA3Mi6BntRsgFv
HU9i+2lfrkqrpOhyBRQEBvOsm12cojgcX4oUpDH95kkbPpyqMId7Podd4GJ2M/JS
NOFwi+HgV269GgRN+66CZPBbCl9T00CQTjOGp+B/ZbXEHAiP8lUQl8M15XIZ8brk
o1VhnSQFwVXOwPxmZ3i69sj9Z319QHOhj3IDDc0fzjTknQGMbw8wbtbovpAzH7sW
Z3HwQC3yqrJlku4matBXvawmmntZ2SSJ75cOJHUCh1bQKM4XdSr9gou1V6k7qbKv
YPhkyXORQjueQdefBZnUyp4d0L3oxhF7c3+3zMfC622Y59EV12EYcse3WfiSHlDK
EheowJXGbU0sDsCm3SeYLFsafM7e9899nWWR8KJWtYPNlFA2gEoqPytww9m9dtM9
IQRbEpfYZ9JeNBc3SSBsC09ZFzqKQI3vwa0eEiHK/r+sRY9FnCyJy6wiVoVGiZa2
SxmXJNh/9utZlNuMrpJZNjeNomXlHrmH6L+vuN0ID2cps19bmeYOJAdLth+y+9tL
z7dqs2a/Rf78GHweucNWRQGImD7Yr0MNEC2BShA1eeIy0YJ6qyQAUdgMBb9fBiu8
zzfoi+ZWI6uZNP14Hun9kDh1q5V3eHqAIkpk3bZOvXfGpOIDaFoADM0F5HQcv1Mz
BLIXB4pFlW06VmAVf6FZZZLeICtduh7Hw6oBVMHi/oa1LO2q6Q10bKDXdJdUvTwF
i/N8zUJdOX/yQ+HuFfnspLf2xTHQ4Ej5D1XbdrzHy2AfSEGOqqmwJhHhkapEJMDA
8GdzJ+TOFuttHwzviSkr2fdpEHdBGxVkS7Kfq+xweN9Ct75gevYIqnIoZvBp8oP0
3IgvaVGy70c3a2Sw5ZM0y2qishwwNkM/nxCz2Imz7sbz3j612qvziUXZ75tgVhzX
PMheWIQIPmftAfnIPDyv7li6ubXXdEpDWbjkvVDtxDwH/e8aSKao/1YqO03l46B2
vF5kIpQmgKtZ96nFGd5zkVYp2mzhClPhdGV0ZE1OmPUCQ6Qx2iqo4g6EntwL6IyV
1QkOVCZ6tX5clR95BDadOb7kbPebMXlzB83020ciSFBH1lzx3Mwo/yYEmjBEkDz+
wIVOjDrhcZ/vG4lM6oRs4fWuSqrJzlqgfYJIbP5iXeqnnSABfOKMMn1NglYaFPDc
ldGLKT6k5zrcVo7M/4d09ZhonUq5n0sTGpgDDRXciRbAn3SEN2LyfNvNM8e1WBXu
XtfT7GFVJzZgOarRa3ZBBCItKFXGhK3pwaJbwtqSsIUyUjH5UDeGV4hjN2npxFAW
4q4A8t8sFrjhheD1wiNCPu/4aW8IbyEFl9KzAwSC0v60mXWMsYxJ/GX7C6RDG4ov
GeevFpSr6UTH5OCJ5+4IQzE/5rdWrvIqM6pB0vTOcwtdxi1bZAuUj9UCsaZiXMik
x9v6aqdv5II3RRrRWC/B1SdLJysKDQHH+vwl17EPeEKh7qrhtzNWG9NjfIqDGXk1
3rely7U5hzalhIyNTJJHexIq4HNOedR/aUew8bcxmnbi2McVODqhfgEmyNwxBWqh
Ydko5c6HopclmoGc/3M/2JoQguQNYOcVk0BgK++S3pXnZlvZ9SrF9tnlx0eNUeqy
nRiiedRmPPm+pQXoqrhAuj2eSRFR0VSdieJEV2bllusSUXg1Pro18X9Gq+gqoqII
eU+x3OMI3PKPoD1MID5z9awKXmwbxYHAV4KddFIBCTBm9JbVoA9jkAFQYnv+j93d
CraQm4cWL5jwUWfo/10OnnG5C4GO+YQmj/qaXHd6jNw2/hMGSNJ9gJjpHeWXL9pi
3o+WXP9Msu4c1zE6VGkantOphylizmu+ST3APA1u0BMlkIQ4BgU7OV8H8wYm3eVN
osvlgpjEztDKIxf5vDJJF+zzj8CVqVWB55fahp4oWn8QFCxEpNoEYWsk341ykk9h
qpsbeAnFpeXujAaKtz8I/NWsabAtop/jQaDchW7gTSMPlLmzTQB7F0xE59imgk6D
rUDxU6ABjcKKfJNPagJZz7+nD/cQNQBXfxYOvFtruoyzAlvb4YaavIguxtb1X9xz
H+kTkGBRcJvGLCRU7+Fq1kgASyOVfzBafYQkcMLAsLDZxZ4WcnhAPN66Sig5uNbQ
LptfxEIEbmsm789VC54mEbbYMvzMqU8MQX9fgMj8j1pdO7B9608gFyfF85dMDU7C
lGP7YitX11j+ZiGnmhhOH/Eibt5Eh//kt6NXPULHfOu3BjxMSR3B0zvkyiTJGJBM
5SHpeuiLPImTeciikUXU99Hwi7SKT3JhQWw70R2gxUG3TVIvqc+rtxxRGMb/jkeP
pSU/ZeIZNj8w8WYihS07fUOHblTgvo/FoyQWCV5KoB6zvS5KII0DWi6aOkgssR0J
EDORma3/PWrFrR49HiMhttoMnnfd0q4f5eUUe1W0u52+XO9MIT45lbPHca71G7eA
TNxbXHqEieJYHbfJnNHaUi5F4NZL5Rg6+ZbJFUYs8iM27lwUgMiX3A3Co/hC2zJ/
KaP8Ll63Y/GeYAgUvidAAME6MUPoAA4pxK7YJyj9AwgsN8M7O7W/So6fD2daYSaX
GUpl04BK4G2hx3U3V6CWC8RCpjB/Qf29aF5kpWU7+x2QXZ2jE6thbogOBcTkzmgV
sfcPjEtnJCiYIX2YcaEHN6l7bXiILjZTCCjOGTGvWYEH6trXZhyRFFU5etRjPzwv
2v45uxa5Y4cJKijZN/miTp1IMJ68HfVvsy/LO4G37h68WBhWNQ2fzolWnmtzFXxl
QqcRbun0zzL19+bBHTM7C5uhWB6xcAiusbbAdQePtRyBM6o07P86I+Tfo6OQnQaa
8opR1ImILNrFkscqn9ezh0PvdSG/9lCmmjOgCKM4QH73msI3q/qJ5g1Atm1NJACR
wbKz0Z3E7VqV/yRm8ssqvSwpj9TpzdirDe2Xtvr7BfmWtGDoLphzhyfEaBUQBg53
wVOIRfnwz3Exgb/qWxoUx2oaUNsqCsp3Wi9+bIvcC2O1uKmX7LyvD6uXSb5u+8bT
OPcqUs3mKMy8SABjv898SbdiM/HzcgLxN6HC0gbTm5BCRszmPMMqVHg580MCHgx2
V9nNVJWfd+bRYAcGGD2QUYH5Irx28CoPdHGhPCihiq07Pd1ul7mif/gMsxS0uzPd
ia6eSrgYOhyTRMQ3QPjd5gdMiFp9g2WcuJlGP/no5P88j87I+jQFDSB9czFge/F/
FdXkGJwFNaBumTZhtUMybkg4VcxGwT0S8TievY9dfr44+ne9++t+StkiRJ/rU508
kfPV7K1Oslr/M9gTZ0LHBIu4GP2JUlWz30DJMlM2Fl2XTYhWDCHmt8dSe4/s0YCk
jmGuFNk7KbSqEB6Sqqg0DQXcEeb4RxPWJJ7irtblBAv03DNa8Mb7dZdit6mZTY9l
jYAy+zNo5bj+fSozmsqH6ZvX05i4PvJbjlNmdRjAGkK8yomQkT8H3z58NoqUaZ3J
cCK4MBjyZdGpUnaxy6pqEHs3psQFnMAcsmdo/cel8AyZJChkPz4gnfrjz6pnWdK+
oaX7JE0Cbdi1Wxofc+4cY13dZvdogzePGOxTttWcfplxTe35vFgmVnuWpO9dp7wv
JXLoA4HKk41c3ZBLLvZKNNMuZr+Nz1JLKjJDlikOP0ywFoMq3en4OM0JMekJqUDb
7h7XpPysdYdyyG4AygPnqMGYGj02uK1lgeND65SE8Ogi4sfpIeJ7bizY75K5a1cV
qp0FCEpr09teklffSFYshPJDRXQtswVj5++07ev5vy38vJHwnHu8wmTmesdgpjmb
0dPIrBuZTaxoCqeeJLYS34xDFKAOH7yySMil7wF8G2nZ5/mTNJ0KmTFCi+c4eAVu
baPP6xriWjCTv0hd57u+S4H6j7/iYbOnZGOfJisbS9HPzcFfU9i2ytdNwjXHlOxB
2dVL1/PiwSbIB0k357ai/SO3fk7/XoLSoMzUMP7zdnHu/7VjAAAcycGOO9pAcFb3
34kh4+Fw6ELFmBKUyQzoSF+H1Ov2n1FsqhBfKd9QyCKbL5Ej0oHIm+H2N9JXbgsi
ChPPdvMCQ6QZDdaQ6CEtMstupwaxxOCTM+mdS/zeDGUnxKrakCEf3ikE/l22JD37
GoQRCwC+1ky4a0HggY9wQ4/AzrFR6UzdbRAPDduFUjCyUh+ZzTJl2dTvLFEDOcFZ
SRMHd0BzcKoLbQlXdFIkEps1ZKGvosIE11X3yD9Mun8V6ubJ/bbeklPUtH5h8l5+
jGG8oBeg8K6myeeh+9W4xYzxDQcLzD3ycKyG5Wo9OIfiCKYyvaMJyqYEeMlWjQKp
mJugXXL5Rnt8uoD2kzOTyBu/RJSbApIiDBeI10hQqniU1NAC47vd/gD/Toq/1CTG
hkbD29PMmBdWOnWsgbBSYIkOZDD1K9oY/TtxKxb4vCk5reSxkX3gIDvQU777MHuj
8xF7P43ZbetNyU5wGmfVKXOi40TI+htk89XSpUijs4zFzCVG/64cEsdaNPtGJmGy
qLPzkY0UGBDyju0QLYrtmZ+Y8q/h1M5xOEMtmUk0+ieyKfC9oNxu2odtprGhHFxy
dxywD1h5Kvjh9F+ysG6yLeBiOy98Z5UaIViCCe0+qSASc92fHy9ixsjAhg3UH+nU
+eLLBiblt6nwI43zgkFs+siS6Ejy0MKBj/8/mHNnmoeuyqfwrhktOqUvdNTOjC6E
74hDlHAYIHwQ6dkSTAYEAGbsy+BT6Qq+mckHj77JZa0KhN6m9lJwEyENBGCFpE+K
j956bWRLOBljUyMTfgK3tJ5uHkkEAlbfSkowK9bHEQ23rKQnXevi3v4b5Y7qHYfc
4tV+KDYmfd4jFu/yyJ+gGJCZcWbLe/JoYVbyQrD/dpP3iI7fcwxWfXla490aj1Db
vyS5FQa5g1al0JqSuJBcOuw7sY310cq0mJ3QNjfKaOfV8gV9nPztMSZTisEQjfOW
lWnd8sAm1UPPK3HRX/2SRnpho5cCBvn5eW2lfVzcXAJf9ehX0e8Q3IathnIN4bUV
mTfyV2IDekGv6CkN3aY5TnXdaUrP+N7llSrt2pQRIzUiKlp2oZR//NWKXwpUzU5m
cDUcVnIyjP2GQyMBkH3X7XWzmcDksPKElFC/L+hgGrd6leat3ZN/Jbyv4GT48MIF
lHbBtw7TlAHWnSkpvfTwig5iyyCXgDEGqzjNbfBqczCCXU76T2ZuQS45aZa2W0b7
MONtDSQeDalr8izDkgg99ZJB3hZwIhPVgiT8OeMflaBOjRfqTDMXCe7wbR1pjc/7
6xLya4hohD2egLDHV9d/gFpceze1w9MkmSqtzQoOeQzFk0fWFtwWbKbBdAjkjybc
iOgeptA+swoxsqdueyfo9D5m43KRwx4zzt9Y/qq7gv/2Wt9svByPX7744fiOevTf
0sHwCPPkhnh9m2WZd1dSPp4WLp9PFKX3caJBnc/EICmrbM7nMRQp01aSwjgGvE6j
vRkdwNdDwP9tYol76PwtEPnsBBF/UHLaYe/4pHIP+SSaAexoOMQ88RsTxhjz+sfv
ew6TVKDwEetwcxMqbJAIOHU6h/cb90mcbA2AdgAcR6MZqeF+rPIeqlLxK2+50GWE
JNUe899hzaaPcUm7h9csFziuM8Ex812BLozGSq6BNR9Bc+E9bYOk950V/p6TtkjE
KVpEnLbmQGgmi4nyAbs35+weOEocN3prrm9yLCNWn5+SKSrGc7XCI4UH61+sv046
fMqe4652nlRes7u7TapN72U//F0HYaOITCrJA+Lsk93sPcxr1ACmGvAgbKjMeFXJ
dybYQa0bqPcJnmgegDwApDDSxnkxjjJ3LNZW/WMIq0INbZiB/p25RUjTAqzvyQlm
ZfWH/KclKIjU3kVcj7a1wcYsJBfeXvDKYltTzOtl7JEmCLPs+ZD5rTznoMWk5wS0
4L2RgjS0v1KiCpMAFkM+9s+sFBfaSt/9WIWTXmh9ltJQ3yqW25l+sr3a0Axt98WF
SZHtyQgiGUbtdR6rh8gW+S4r1eIkZgNCQwc+kPF12jgovTfRLd+SkR0kqnt9WV7P
5eKb177kYUPXhsDiLjooXomS68BlToTcQ3kJ/1LTzGYtys5o586ju1PdYWxysMcK
Yu8V9HHQUmb5Ep0HdX6fW5isGIMjIp75yOEjPINYy1puNgIXCdieKj4kwZT0N3Il
Z/aV4PdWU3L0+WSCDyGa058cpou2YNaqgVx3+AiR7u145eVPZuQ785BEibZ8Dxtj
ECrfp1NoP33OYwymU9swZ0qliMYHvlpWUm8VC0HM74MDKsB3q3ghc+breF8bSlZs
jy7BKSNUpSc6xe67rxZgRCXKQMhKdT0chk9N5Vsq+NKP8oLfleuDT7v5jfiwnkZ5
8cCZFgp0xepJaOa1dZ6z26x8fR/JGykCn2FBWEzlDMyshSG/yE4kgYpLbWSUnJsd
LjHftzlpM6/rp0vFiGYCN/Jii+APRonmHdujTbgA6EODtN/T+CnDPMw9np4WXH2Q
i+qRa+vB6fFRdL42Qp2+62glP/2UZWwLHNWbgXykzqSdo+zTVFOWZJ6BXBPb+eon
CdMYEo4tXGMaoAekHP87otWJU8jdVgPaJVLDZd0eptkNZ7WjO7g4fOi06iE+EYj8
AQej1zWFIEt8bxxn/JAsCL67207IM5UjSpZwus5/NGiswLK2EORlx+gVl8skQIHm
81/GMh8kCp5Xf/pnQirTFbVsu4M21N+1QC0q6E8iO5Ah/7Ni+ZaXa/dYKjwJA8Rl
9VTjB48iebZeee1eQw5nvGMqTMfSKuV4NEqgwcIFIM7+494zyWHgic6w9k7mb9H8
1iKpzy2cu27a/aIt9oK/rNuvnjxz4iWqzx0D11TfrOobHRvqLh08UfgdtCcJK6bN
kF14AF2i0woTQeVGsI6qtX5BAcMpbkCkTL7OmXgmT7rMRS+8KRU2p0OSF5jJF3Do
SCeAP0ny38l8AG10SUzg+oOIUNh2Cms962XSkJuDpIK2FS0svad1iQoxYQVJf2e4
9q4XrTIEolhpm1ZZ7KsgHaYvt+Rk/t/HfUqO9g8uktqyTxasnjJ8P5sEuSdYa3Hz
gxYZo3OlBBlzRkggKIoQP97/VfyGT2g4RO0X9H7L/MPwVf0IqpAya0qf03M3nwat
gW8fjcwDSTGt8vajL+MWfA==
`pragma protect end_protected
