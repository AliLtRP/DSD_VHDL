// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:41 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
robS9s0SEcUL972hrAVu/wdE59DCP7NoVGAtYc2i1qz1+e1BXUxN3XYyT7tss6BI
Z4rRzkPyX4wPRvHRiz0b5KfE2C2mYWL77w0ceHO6c6li94g+ZtShLCNHD8YJNJAQ
KvM74yAgslCr3mqOmNjNz0m7yNkUvViYo+MzFwTAV/o=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 9856)
TD3rcfY/j74WFoVsQ4p5jDPpIfHCJq/JkMnJ/atXWhDeqeVl3Sq1pProzge/KVwH
nCZoaqq6leZaA8mP88nZipplf2Z4jmdqgk9SKQW0MiQnbv1cP9XOZ7H+rVjlvb1x
rmkSuw9N9MqIyeLZ9hS+IA1qzRToe869ZhmqNXerOwLBqYoCUrp9NIk6QGFliX43
GKbQnxWuUX69ruLgfwQDzTq/OEgPp09K7hqnk9z8ix+VIb7B2Q1A93vAqnP1lCQ+
uXH6HGDUOufkfDx4yhtsGWfuBtTS7UxMgsIxc8OGoWt1My/aY/pgg6KOWERhT+S6
py2z8jZzeIjX295OQ2Yw+UqOnT9rz/kLdt5/ZXMbxMIG+X+rA6xVm64gtEGfnKxL
kezVedCJ8WhwEx0W7Kxjq7UzkNkReWwmsYvyAE/hHpg8yftRVW0W730s6xBvvjxy
tT+6JPB0zuZL8J827B5ZDAmZXQSBBB/gN7AyYYgOcNmyyrZGBtEm+AvmuUHnVSo4
N91kNrygvt/gNMvzyKGKTMRlyz4W8gGyV27CSp6Tw7XPi+xRov9TbORz8XmJv8mC
8EBBEwjMJxB4O7l3wq/gi9zkcBj9EPVIo9KQktCpYrH3Xaz5qVompT9AFqE5zUHo
OgqQddVuYPGelpb/g5iJGL165jMVO8WOhsnV/5u2PFTtD4IrCnopmE56gwLnhiHr
sNhcMP4k5CagBIs09hWRmwCjEGgU67ganwhKovNVqr96zUf4heBYgnFxJSQAhYM3
OTjGWP3cglbYrMRC/cgHRWsGfv45p+WS58HvcKaYC8/yX+Z0UA9fRy/PzaMla0NK
ExgAitvZcaEXgKBcNe/dzdT4HXOArmo5neAkWyqEd0KLeLgaKL6/9YS971Tlitgr
qYySLywjAP773Skg2gMCOgTe1wchawJOSZQ4nU+gXLVSvxKwpaeiuRGveFeS9ugL
4gu2iP1GEnrHmDhuZ2O3AWVHmdem0Rhgr8fdcGFs8kspy+r+uBhdVWMo9utdO5Zd
ONbKUZbHIuA9Z5srlxq1aEZDodsKlkWMqEZ9hb2rjXovC3Wox58RrtFmeb+7xbrV
XyqhwnjI4clf0GGcW+RLe9wSegVqQ1B+p3fEQNGCNvFDlL4XHIK8t7LPLR+ZubXo
AAvamaX9BSztUkf4AfScNtsIYQOHieM0FvdrpbiY6sqEdbCjVSv2JJ09zTJ9U+lS
lJiuF2cq0PxtKdLKXCZjRMKhedvy30Vnf2tdhtv4pW8g5N6LmyGoKaY5MsWi6/jr
ZFnPnWeqUX1A1P/RrYefhcMtA6ushJOW9MeWK8iI9fsg8PbiX7hoPzTFyWrTyr7t
EqJ+e/SO06C4iwn4jcBAuoF7b8wzlB1ClTuTWeGEyMhSaMag7L1/nGV+XqMqhXuJ
rJ4BmbcOtNueXklVL8xAbQQebUkyPNgC76pRVsATJ4//jHxYzyy5X1SzNM07yTGL
PXNGQPSGQw7O80faZVT5GH8l6+L1U27NxTKrgQBMhudRvUMn2qbTpWfQfj6fIvKp
tK+zehn4gNL05dywvHh5A/yymt+Ve9jYeNzXvqKrnLfx+yUTa9h9H3PUkUQ9Ee70
btYKPRYoJHMf/ejl2XP7RwBMCDUw1WPL0oa3+JpfyFW5kwZldoo9of9aT6ysXTF+
657cB3rRJ7o5yMPqDT9bJDERLPovOERP4cw687kOWcF3AFVHxZ2S+KJXewzH1fwk
eoWmT2hW1wkBXxOXrB7sjnNc2+47onjV6vjrs/HoIeu1TBTXJ/aBNT33wqlNIZxa
LK1geescJawbPj2LQt3s2YXpleF5xC8McKPWo+9MypsSzxh1UokE/GIzKVKJ0S32
Ztaor3Q7iUp8GAi0AD7LYTrOmndGug1eAqpePLGPDxQnqQzatuTm2YmcVMKjL7J0
MYoxIFIQTfZNHtj2XU14A9xSXITI1GddH4fgOeE+CmQIiCcfT2PBbMQuHGZeVHTi
wtrw2ExdBeJU/JVK9Lgvimv6VWZiM44dbSDm88WvGnLJKSl7nOTj960vTbxqETnb
jGH0WP63bSCzDr6IHwUNwLLPju8plEDOJA9lG08i+H0BbCxOKQwgSYkPpjBCrN/2
k8fcCNvh1LRNDwyzY+kU9+kaivHlesCjfHuvCA93tSezbVNCS/Zue1q4wUTFoj5k
pwXnb3FTXwvTH0ZJrmsAEC+uQmei13W8EOQhAwjYgkSI4azFEJYn7EF5Du/zLkPb
0MSuBeycijFcFyW4O7bdvpkWUX2hva8//IMfnfDbJWnDE5/BZE7x07Y0lVj2y5sr
J+5T3wPHrxkwNNJdfeXu2CFF8orCaFNBMuflMCi8rmYIGRA8ST3qEsCldmbMTYs8
vx1zVIN7H1aGB1Hkn2Rv/JZTulfdW06SHsULZQ4uuvNc8oJPOOzV26XZQ+Bz8sBy
WqA1mAm22eet9KIwXdL0vHzjbg4U8kMlORMI9/+Kirl4tSJAaYvjxWmxt4f91BTx
Y6vB4dfjh8xZm2Wer7NWW9x5Mi/tgvtfH2kgcIFG1PG8axKY+uTjrfXZdeMB2K5j
NRl9+Yrw+dZ6Ze4v/r00bQXcy+fIYCAePqmvUeGmyBud7WfM81aq0/Ocs3EfTzML
cb7t9++tLrInZSuhkU4ugNilbdvImXRalyCpUE0LsJBAV2o22R8muF/bvh/yN8xI
QyQIU8aNfvHlFWN2IjyFRCMCiJjaXp1zzuhMpUJ/BWwWY09vQmlhXvFfTK0u+Sf0
fvXoxct3l216F2J57aH5X4XCM7fi9iZpCLkhEGY8dQtUc5pheECFSpit8420jV9j
kF6MkxitUGSCbDZdlZshPoe5QwiTLujN0yQmbXYmodntBxra2lYKwhga6PShpoJn
XewP/R7m9jPkiNAZZlNlXxLYuGqc+KT7W/Mnbedo/LBFQ73rrxYOoP47iXqSw7it
9uow/HNz9p7GxEb96nEen0aXzBM2Ivlf6rlxaKXCxWJE3KcrrkSn9Pp6Oj9B/l92
6gRSloCDRskmbHosyQC50KuiK5VcLwbtoOXPibl0axIYzdd3vNOqg7HoxL/6n2s4
3rrV+GZkVzBeLjkIO1E02chZaPWUmku1Oy2vKNVjVUUFBnqMrcslDKtWfCzI8eOL
q759VfhHHlQ+rkk+QyetCn90Nsz0zsWLcmmy43I8Jclu6ylALNFjVUJ1RABKpXWt
SOtawpefLCyGtnGLAPU/scjKAsLzXTaH8PNEL4iVDhiKYY4RKbEU2XXMrkknO3Yo
ItJQVvyzfdgvz4dOu+dDL4VABXzO5GvZc1jJsbrVT01ZDulgwTG4qcjCUQasorbk
l2bgVWL1G/0jTPSdwo/r1zY9BPNf2SgnATZHPqQ47+bV34QlzayK06hp5ZRJ7GA5
jaSJcCKcwhVSFFqftzznYrDQ6WfnH8jzpdCas9Rgvoew6czr6SOZMeYi3vBcxltA
3rXeWUWXz/TtBlA7lSRjCOqHsuJ4sVyKlEVfq5+rI6wtcHl/fxBQrrClWKlyvg7C
Zc2U6fkInLcu788DZDbq6XpEn2PREp+M6+3PQh554tN4LIJ7PJrTgeRHaf6ZOr5A
Cmz4CXRq3j05fvIYPF1KsJgoAU/VZlUow69C+XEz9kB4UXJTwic3gBc4OccgJSxR
wpdDStf6BWUBOFmaQUqnGyyE2iTTtsXL6W1YcnAGE8/meroMGEyWmJNCrPR+AiBi
b1pIpsBAJqlwtomaImwCeRDpOr4Y0f86IkRTMHgFwS5ghYzI6IIiwUvPkBXXU4HK
I7szdUKrx/eHjIVFBEIAFj5Gdufk1p0h+S1kamy2sA9eHdOZ/O7KLJf5BUZFTlCJ
BiMKzPET84O638/G10/3E00WU5JAsu2e7AzVL6fywK/kHYx0xrlrAz3PjxVY/P4i
URvznhoTig3pjJh2MDztPQkwstbmeMMiCFjp7xZVANIbzqyzVjB/PGqZ7dN0nLk8
HHri4mQsNVouueNWXUd0C6SQX4esvsRxgcaQDW64ZOqZBsB4aZp4b48YbmD0Grfv
YdbXQ7E5kTnkdFYlDbiKpxInbjNWAbomvQ5+oxYc0HQW68+671DhSRDKH0uVcHLV
DuvbyjUXIjxvJadneYB+N/bKwO5eTyfbOdZepzV3XdwpO2JKuM1Ggx4DN6n642hw
1yCM+LCVNS+U5S6EqWiR5W4YfQvTiqzN92SkRSes21nU/MuTiKodzZWw9GvwjHZ/
cxJ/tsgRa5ooNFqb/FoXF6juxevWMjD7gITI0ReDFL8GVBUNm5+vGWXCvpi9YYV8
GIk+S7G3G/8a3qtpeXy4MEekWqmtcbgD6B0Syi+e05x10+yvcf+xHSJPV9899i30
s+37X887Lk5LBtlKShURL3bmxaTyGJHqKqFdKE623wVD/Ut2zlEJkDEx6w4QANeE
Hb6uiMQumAUprycQmEPVbtUYh6/c35YrUC308vxn/d8T9Ny44DiK7YQDPTsD4p7I
tDUdNGU8V26qmXtWu91qPfk54e/CcSDTXpRe6/KIB9TyRnipoTB6A8QyaVdXU2c2
BJxQi0jrCZzyDFOzGgC0Yi4b/sINrWP0FPPQOq5L+B9sfnMJhbAjQnabCCigCrbC
/NoOMXzoLQA2Z29F/YL54pIrG4QSArOPKtIYRaU9//laCgoVO9mxTjr5aj0Av0kQ
Jif/gLhbj8RArRO7Am1jAJVsZYHhKX9nzhVZQPPhBCWDds++1O195QV5v1uAFykl
ZBkN7AK614a0lGIYZbonaCJADK/fFxDfSMNLGgQ5nAtdFRjZmlNQ9G+ekxEKq9Rd
B6ZwpXw9jjQZe7Jv1tu9Tu/RxpVlCDn31M3zczsoZpBACk3N0RPUEUuqn6gLt4in
0I6Dmiib4RgdFkoloudRohrctjnxi2/95Ud1XuPUvPyz5dD8hHgz0gDZp8zlG+kq
4uIKLV0xJD+89t62HjrDssfZnCloU71NdK0m51R91Z91DiPVOz4uhHcAxipHMaL9
g3ONsCtUdhyS6XtOS9qje9VQEsDBIAt5T56haki8rAOsY3ecGrZHOsJZuFnSK615
crtxIWDBaQmhHm15cXYUNlMCjqPsacIVyZHzC8l+Ilwn+z0NoGC0ZlcXacxXGoRM
KAnQQWbj6OJipYQk3zcC9eaErjHTBAjFLEC7tdbJJaPvE21O6wCWpeRLQ12ejhm9
KaFgJv2zupVikjZdGrDTZsyEn1fr1Woic+x1PSLTG3DvsUJp1bPLw8+oMmAfLAXT
R3WZ8gGANtM/mFCqaGZVpjSpF8hxBR4h+/pz7ieZRttjXbKEUci9GHC90G3WXoY1
Ev7qlSBZ9d9wmjNmU7uL9EcPPk35CvRlfeh5xGcPrypJgWr7R6rs2mWELvn4GwHs
8FSD21z6AimwkwhDdIDOs279GwVNLuqy3lsquCxXLLBDA276U4gYDqDMn5Qu5ucR
X1h90We6qulGo77a99UKKUf3DE7PS5XKEaZruQLDUugE0G/lqjFUggDT+otXeaLC
HJD9SKgzPwLkwlK9ohY6FSntPeBzfHwks51uxowa+l4i9yr54lA3wUGRU44DlXWk
Tcgs7pr0Y5ceZQ4edQojNdgX1qLMO7DO5mMscYp442YFJzymK+b/Oz4yOGfaz6wB
gVnl0zz8YIA2T1PDcnCwrDX14kucgu+bkhnmyD/LDKtk5i94FDYfyqIKlpmkcg7d
f25V4FqScNYVzLCLXtmW1Wm8DqJs4klZoDt3Jvo0OqXoF4M1wMFk7Eghqol8wmKg
YhL+Pxi37X7H1DhCvrI5I7l4glmPSZV3vOv8ezcaqjHu+TiBarAfR7cfHyMs5S3X
0rHr2ref/toQY3hObcg6MhxyUhlbcRINoM2XfpPwb9VwJHA+ut5UKXGgdTjP5QCR
YmI3bik3OiP5yYDJXjWQFgRMQnY1q4o5ykGRoZmGegBI2FY8SmOP60ZQcABCkUUq
TvfaMMCLtKiwcYX8CkYPQ9V4Ms3m794hZbElwMVNhTtg3Skuu5yTFqEnDUmEPx7/
BaUQdOqcZ8tjfKLV2TJ9M0GVh9U65RhlSJ3j0KqFefvomF5aQWj314opWo0Zc7Ly
COd+qtqP4mqyxm1jdIAV1Z30hPnCLPIdazzcshEiWj6WAtt/lexlxm9ymWO00NUj
H+TU2fIzHGvUGfayifIZ5yyeUew0yYt9HpvTGiRU0dtgZsMgxeQ2IE1Bf0js6K8G
zQSrkjri6M0gK5yz47tE/5U7NXcHYkxlnPFXRBUiTl29mqKynFPxDue71YsfYmDC
Z9zqCCqTIn3Y/Ph2EXwkPdTvuwLnUVm91U4DTWseL3eNF8xf8uLVXhSicBBnLrpS
dIL+jB55zDpxCaKfqUCwMyg+Gf8aqcBFO7SwouxOYT5o05ZkJN8nwbMI+U29HX88
ebeNcVqWa4agxFt8KLEXyCMUxPjQwAHcHuPE/lywkdglR4evjz2ECwaNXzRRlgxu
YvqRagDbG7POk17nBRhmonoJmRMr5hbf4/o8ENLy29AfLA6pHo1O0H7zsb4/5+V3
Q/vYjgTHbWiCenuAx4TVOWG4HD4UiB8Ob5j7r5h3MCNgKizSKwN7qUAmuNOc9jFV
PN6EADFmiVvETq6Xx3JGRv36oGyH0DtjXwB0GI+bQRt6IAWp9v8JKikEpk5W2Ap7
YNWoiLNVlzib9hPeDcN1kPGK5a8s2/fT18szMX1gikPAhzyfWCNrolAqNnoVTIHK
CPzci37K8DfP2CP9c7zNNU4bnYvCzPRqRIiJh0eYcs1HkiZUSLTjTfmRd1XiIb7s
98xKszko3ktkDlWJr8x0umCzdXW62OhwcSJKZ2fQcXe6wTQP9YvGnW+NezRegyyC
ri5iLLpzESyuMDEJVR+vxjmWcflO6mAg6u1kh/wdq9+QK5ZC6eDUmYu2Egxm2Lvp
sKgHjN2rf9gKiGwzSwUlYfYUlxRGr/FENtabn/J30es7nmNeCi9dsYytO3Q4ACSz
Bjc0rWz0i8sVOtNdRVcfN0PjQERf3LaZcF+3cPEHuG+W5r1bazD81Sgtlit5lg7U
DRZo2GOcQBWbFmOcjbA5E4nYkWAn2F+PYJIErgYzM3ABAUKpZqOzfF6wVQEpDn+7
bDbJg/FBdT6A1U9hNLwEY63DeBWeo8jGuP2PVRrp9dr5Pp+FKAdNFjYkY6Mz0bp7
ObfmEYkULrBq9JhqTOhy5r1huoQ9aiMLUjBJicz3v1unel+J9S5GtM9bEAehQw8g
wzPu8U4SZZnSVN+CRuJCw0fORQ8CmKF83TMwL2y19Fk+BVq/nmHJN3Dv9T5AakEv
qfWQNmPXM1Rc6ppi1SWKKJJe41/4ehSKSxz/hxlr+go16q9wtH4xsFv1kj4fSLTp
zEJDSKswOEVoK3LASIGk1Aes9xmcHe1/X1xCE8uFEL7cfMmaJo6VQp3ngchsasUg
cqlDBM5XfItIz2W7xkii2M+8qj6NDt4WTE1BNtd9EX+0UgOg8JO59IiPYm7LTY9M
AuS0CRIWX9XEHl0K10zIWHGnAWnygICn3p7chKCAnsffbciaygfU75deAQ4VvypQ
YXZzfdyOsvnefVOK3xf7foCRUN9pnbFWuAiWrSTHY63QtAP3mBqyIabV4086fjrx
nNCR6NiIQhnS1yqU8idXQUKsPCMrztjNTiyNCIXlshdL0W4/P211nnuZMWDsViaP
pqPmETkJnSIs9bWexSyKPu40WzrtoAsl5JV+LjAr9pbQOCG/dOm8h3OTnuNMDMQ3
ubPS7N4HB/+//jR4sn71r4bgQqfC4MqgJdEUoUWMI52j78fWr91paEMTYjG0zVj9
/DDbwVt21auNpsYWcIF8ePYbt79ljE/ph6pxLGlXrqRgn1i1/j11rCMmqmhqY3+8
TiVUyjqdw0DZhXpMIg1nBWJUO/Eeib/xkrqwHe2ojdNGwan61CL1Gm4rXKfAe6eg
CPBfArDRis0vmZ0ZFpBofDFsOcpCWuWmlnI1AtONIX0nNhXciy/ZN98CjfjmHdkH
E7lhRDWYiRP0UKLtDAkQCATtO6ecP+9X3gFjwpxwXvgYs7vzZ2OhLOQ0vQsmF4MI
Xe3wjTrIWj7Sn/MMeE31wPsH05M3x8sq3ft6fXe7Bq/5tw6HmFKbQU4/F/iP8a/q
eG6kSOUFC+ilb8UyIscGrJZl46EiSVJViyjCwghm1HMQ5pfbfLFvWE2Oe22GAljh
XadV66UO+n0SC38aAVxNusxs+QGK9m6WuCnVLZCFbidpfZlzeDZNoXLYi9Yd9+/I
YZmhmS9h7s1uEHaOHuXsU0UZPg8pjLCpAPAPuI4bWaDhGZu29gFcZgbeQBkUMyOv
1ngrX+zWY9H6TOskV9JpLkZrc3raBXuFjYcTeO33DQY9i9krzAn8KoBD9JcynTY0
WUhkhrGeOemlV7dr6jhFEEPlJ197UrW/6w+9BgumFH7p4ihr+kCJSyqgxk5t32Jk
ikMzuaOWBBgMTx28cxkfr5OuoRUZntDCecLanF0S+cNRGPwGUpXXkLWEQCyiCEUX
+KBwp48qmaeZak8X4qjBXkG8jP6H7ZzKlXUwbahCZJb9syiyu4HvYcUk1SRZ0i9c
+jCJ02I9ZHh1VyOV8dQsp/Ol7jn4yx+QkbNX/334WpVFZNzjw3xUnfEZuWBdzgh3
IIWCvxB/gKY6JjsZkT5/xagGgnSd9VIS8HTqt/DZndyw4/ZsF3H13a/HbuKN0zzv
K5eyE8XXt4Rg3LkNyEnCX/k0WDlZEGgEssSLZqKwI9NpMw8gnnwTOYQra6FUh8FZ
UpUT5xzHelCRHQsx67apG99+W26xBJcwdBdpcBX9UwVcpoh2yUY2eL263pU4W8zf
bcSI+7v1QJjyDcOh2shpQwM3Y/5kH8eJWB4Gm3qKqXx6aKQeDTkJaZsHWI6HueT6
SE5F5mAOiQjqgt8deaKpb+IcC1itjgyRqmfv94L3XlKil/XHVZyYo/vpr5L1aZVJ
MnC0zWnPsGHJ0INizANdYo7JMpuwveoc1RMXt0rKCwgFF8+1ePxHJL5IKWexfnqa
cU36DNQLv8HGnmCVOxHg0sRsG4oSm6tUw8vOR60tQ7Mfkf1phSEJYB7x9JnjUiou
a0JG4jAw6NaRj5Ml267fS4zm0Thq5OC+sOXW2V3ulUOPtTox7YwNm7ilakHeG1KU
6dGqTicYaBIPclN6sPDCx1Ar6NAjq55jo2YrzZbJKTJW5PU5W7sBhJOfXA5nbT00
YibO0X3UYf9DlM2k/G2sApNhr4QemOjb99eNNGpo+aX6jJ1RBatEjQNXgGQkrsc8
kXqKRyJsEjauGrTaR1E+tn79+v7TxoTetDSd4WZI41s43A4IhbW3WD5gKNKr2q4J
k/uOQVachMeTHu4aeaoNQzkauscwdkVKS8fwL15J2JGyoQ0K2w+O57oH+lKap+y2
mqrxUIsEz4ruZpOeW9M03TpEXrFqBi2vA3WyBf5HxFvExY0ztWaToLxpAthz7aEU
iRx7Vw5jNWKtqu4V0g5IKd0jUXWjevcWmFdGSKlvCl3/Uk7pb81wG8KPVJKXRYt3
SyELnDNDdjHfbRHSQcLXz5MJgcJ3Eda5zR8lLPlorfK9ErIMjrI2262a6slTkfoJ
SPe7I/yyO+kBEBSf2Yc13dwVBI7/qKM3dxkxjOH8bLE1558kRkHunU/5vDa5B+yB
9AaW2t/i1SldyNcyoozdHdnk06faidR3fINlf8SqdOfoNigtO2TqX6pw8xubO7Ew
n/x4c0zgbmkSXI+SlP2iN62njtSpAMhjmfoZdSr2l3Qe03qo+xM5d0XcdpPXvjHL
V9QAxYq7pZ+7+Wap58HVQDOuVz1ngvJvMjvkJ9zvRHL7AugQmarq6w9g40XAbM/p
t41LcpfCbwat+U6MQ3QHOM6uY5ru+56JiF1/zDT6ACq+x00NSpGXlgfomIgRyqIJ
P0IwHD3zAr5nUAB2nbsmdRSg6pJKz0nk2CAW9Mu+aMhJ3otAfFFEHyWz1zXfzjgJ
LJExNl22r1+zrSVU8PhF0sSbIrw07ALh+f5astkAHKNHQ5mkl+JZ3wqmsXTdgJFg
Jq5hXSEPDmNvt8GdwsxMyhSHrM0R7k47Zx+zpusOm6pqQDp9f9Bku6iYCe7PBOkL
0xzAxLjsu6BA0JOAUGOWD6Mr22ktgX9MJb8WsyqDtXajiGcjQtvo+x2/ah24DC+1
6gb18sUi98mvfB0iFMlApkt4zW37YLldxy+jdLOC1cih8ldC6L1K6bV2JHCB1xKJ
BbU+W/IWGNFX40Hil0txgcZaMEr6bpcVanz0kJeyG2RKtZW6eLUPxEb4eSxGfQkW
mFWfBsEeJmAM/s2wHxZkwGfRQ0fk4qR4h3r9OseIQzt2E9h3iJoQzAg8KhhqF3+b
WHRC/oa2VS8MRr8iJeMgW2X3rQIqLeZ4SqWQrWuTKR0Ba0HpXAZroCguAL8Wua9F
B3DHogPyZW8gIrAK8eMPSaojacFV5kHYMNaHBm/O1hbfH3OuBfQWeFZ36/X8TsC6
CyCHAGc/RUWsyrcDFn/3C7VBdJMAbSgigR77alOglCyUMOZoopR5ss5qTV6u62iY
86JHlX8cjIA+/hZ88keTvOnUBZel0DcWaysuMADy431yTxHu5Q+lm2F8490sHi9e
IpNO/ntvyMLxqWipBm/BX4yVE1Fef0NJ7OZUgJoIEZx6diweF+pKfSiaB9MoiPA+
7/zzZReK08pSfGibCJBlJzF4It9GJd/wJyllawrzKf4Tse8juPKmoz7apk+ds8U9
c7MgbMGHEc839Eu87LsQVd0exEj9MKL+4rxuGg+iNUlm8TtYi6hz1V6DFnw5K879
hM5wsNqsEsk/I3xIp2PF5pfwtHj7uE+cxAXN14cCKk1MlprdiO3CQI1T4etwyNhL
yaw/3eNqx5ym88MueTl1DMHHURhvVy/rDnP3OGeau03SqgdKjNbASYLBO6AmCcBq
F6ypaKdzmTTVWiygN1RX/ICT/EtI2gWSJBQtLZDMZw3asjn9EnICIDfrd2PmbgMZ
Px219nWKHzJ2OOZs5hFIeOTPutsbtZe3urqHrah7s2wiTFjelhY4zLTT0SfREy5w
A9gtcf+IkKIUXgQ+OGPG9zOtd+0dovQ3fUUfncWGBLEntJaFFkBficz76EiHMHIY
49yP6uwUOIaPToFTG+J/dO5KLmw1BMwKose8+G7PYBC4qiyjrg8Emhdi9kzOeq4b
c0tK6gRC8S5bME2LlhHgp7sFUR6QdHjE39DcVvyficb4pImPhLRK8IamR/FcPVNv
C1XcYFVAU4HY2GU6D8OCRP/HSKopMXil450wJhhn2on25sruF5ZE5KDYPgp/W+cs
B8AtpVL9CkQ96MinYHVxXYrDJNB4lVYC5W1N0XUF7aqjy9iwL1XG3arGh1Yz+jiB
ZqGeQ80yZcSwtT/ZYCVuhdqy+IKkQGo2rNxnbHeDwH+tHiLFoGT2sxk9OkKkFOkx
PZjeAKHEz7LngWjvnCLWsjhmVrTaJkcIhOwhxfWqFhzWhjaiKcHzF/xxa51+xH6Z
WZ6hiMagZQkgKMG+kWoTWkR3azSy0zFbk6B8CDoi4jL2E60jVxmWa9AnZQo2P7hD
txDB6DpG+5q4+7CHWeVvpeuSSmfeiCVZchk6hljhuzCpZPPU7hbVWhxLcV8ndEdK
fzoPvW1Vvur1MaBlOzvP3LrWTJWDBMmM/Wk4Jk6WltjR5LZkiQjbq9+GYPQ1wFrh
WM3TlPyf+6dl5dDnd+kf1OxZnJngdhBMboPBBKAFAXy4taTPSAWkFhYAZ2RL/rxZ
N+RoxyvuEX96aBVxlw7H0fuoZBwVZRbkiu+17cb09vRsmzR4FFS7hPKvXfPuwqo/
EF8Y6FT63HP/PhPdfWr8GzNv/n8Y5AfPKlMOd+QVH6iV2PWqsZPHT6qdvqEnTHxv
+nw7V28ejunvlprs9iJDLcQCWP1T5HnECSppiDaTbXQIaB66WbaHeSND+T+V6ebi
J6RxooqFZwIPlBx/8BHPECDMm3MBeJM2u8CNhXd2jaUFpPXf+F9uHtC8XAd2PvZb
38a8n1OlNv8mv6g9vnAWowWdcfxS27tJimt4RW2S8930K3VR8Cn6/YCyKijMUcla
5tBiesssBIdM/M3sdF47yN+9YbvBKmmODdiY7cQkYnvA6S8t7l7A54mxl8Mg6UPC
+8rGlX+KWfrvnVlGuFLd9lvMvfP2ozQTrAGQ9kwythIyW5AowbEj5higLqposw3S
8ysCMSnBYYmbxz5ejxA3ui49P/SCaT8tuPs+AjOvjrcMAeyDgMH1NlVAQHB+YwmZ
dyJizv1ymuAQfJvy4wJQsHUdYrOvekpQ5f78zvVX9xp2Nv8SAz2ozKC/7oeCQzoH
ATFAfwzPGGgsMtxPhHxtWhRIcKRVjuseigN70u3AI75MSU75LwE0VQ8waEU/P01z
DqdIErIqsfO1yxuG0c9Z76db65PJvX/8RUCS3Cieu6NugGNn/RHAoG4B8aHDob5A
Wb7pSTgbnmv8BOZXHpIDp0uy7leDc0B+o8A9UO0WJxmZJF2R2PEwMECVZzHjlCb8
FMSyKlcupUmIY+tsu8wnucS/9LMBwmjAbPGNn5sWisFoNxp2da2HwWTewoNK7gLK
CcZtuueYWmKebn0/epW6mDFmU32BFW/Ovc6E4bmuDvGboJGOBVsQcznqzH1g2rEq
8FSZyE8Yu7/8wM/VuG7QsRU6yxFYbi03aUuhu9wPDm1jRJV63BV9lxrOwTk4rFBQ
2ynmgw8LzqXEKqZv+LdYza3CmQi7uFUYTjeCk1PHxDZwAprv3B8mCT7Umzc1/Yjc
zLP94Eg5s5+73ieRAIriwfwFcEY2wp5ojRmK7oLN9NGDA67oSsiiY9xlo5nYuQCq
8xI/t2Kro7xahZn6qHba3b6QzI2I/m+YDqFweJcXr+YjhKQSxGw05ZjRILF673/v
Iwty/iu/GJqHg8ZedyghWXNnUOD/otKW29EnwFkNiIHxRqSyl+I1ILQ5tl+9bCOP
Wy15JIwVjNrRUQdECv2bJwNkk9JXengmUQy9grm/M2oOT4cTMSB94I9u+wN31YZe
+NDD62R6RFua+5ausD4Dp2ln1ux0Ng9IJe9LYuxpsPiwptW2pFIuom7uC+YgdTnV
j8otyZEhzl4qA7fas29BPw==
`pragma protect end_protected
