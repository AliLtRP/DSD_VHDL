// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:33:59 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
mKw368i0Ycl0z82xM+XbPo7Xel7ksp+smOnJwk812cv9zQndQYxTgVra430hnlWi
4/4wDMgEBII1KsOilxAiVuldvSocT4moMpmTepeEHbrrdeOgQOc7CINyLO53wCK6
D2P8o539QnGKwgVesDF/orp69kVdLOu290ny8fRKrPo=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 9216)
uDbR6ZK8OO5iFZe/ycHesb53EuYg9E4t3J0Ipp7cmL+GFS5WluMf9xtlDftc/axV
0LPCS6Tu3N6quDyQS5Mar4tjXMnFeGoKiRE+gCMhzQtCxushIFl7m562QUCF8lt8
ScOULl0RYqZutCEer7DKpjMVBusQhK31VjXgpbWWKtYPW05BthmlgQEPSl2VDxUn
Qd0Le0QVrFKHoKAE07y1d2C8KGFOw+JYtGZcqED/lCd5aaCQOmqYt+zW9Mj7QFsH
uXads2ID7r0mdArQvNi4VmuHbod6PFnMt7fytFopdTlMwmjm20zObVNDjcwQsTps
kBlTuXTlHwaiLqbZaS2TcmKe1SvIFOztNGkum7ZtDAUy85L2ZMHkZXvfJIh/0oVw
57yplZOv2lDw/S6fjRqPC71CmCCOEDzeoQAJmKf2nkQ7ZkCYg72RnkOtWkdObxEh
2GNAOJ5dYbactoWUqKBY0D0YqOgmFx8V6UAVpz3/KJaOBTLS9ab55esSP8bxfynw
0EENl4L33H9UDf/akqeX6c2A8h1IbXbhg8H37aVMIeQ8DYwNEukgQtIYOJ+WaozD
Z58VSyLQwYjWl+9Vsn6daJ4PuO0yzykNjZ24oslv320elJvHmnaNA9NjBm5BSKVx
j3hLlx2wroHDZDZ1UzfQ12dysBHpkCyk0/Lqowpz/f9wTTru2s4X516EdFffTzMF
WpdLfECdt0cEMVYAbLu5YXZTCs3yCVrEYxxr/abNrcQ3hECPg//4CChTl+qEisAz
CDFAC5c1HEDIaMFe5PsMbE1c9gtP/j7pR+LV6DddU7Jl3XNmL2drfYh97FV+9sS8
2cxfjXW7EtC5GUakxlDbg5DzqiLS38qo2M6Ogm+yog0+ks1mQfJj8IOhTg4EJAj4
/nFu7vm2uhn0bX1aIQsfpGgsu7QWTkx1w7XObTjMOEp3hDYeog7JD+rotjUP9oDg
tRAJS2H7zNRppcbAeW8uV1GTj4kFgZflweSEkW9Z2V/FD4OGoF+V/O0DJV6syVuG
w4YoGVpplE+CS3Hd8iweiEgv76r62wbsuCJhacilJqidYXfmVXjYn7kqHDqVZOzm
wWqZuf6+SE4hZg5a+abzy0rIXDzWf9G5HaRHTGI+9tudjC2mPWy+AtMVQbe/CmSB
zI70gPn14/SeGwtOya0QcP6gV/mg2V77Pc90sTrTPfpR174mdvUag5WuugvMOcC9
cPaln+3RFcipSR2XNNe8ZhVglruzRgo0INNDj2bIaGWMNJ1/ggs9Bix5BIko28gg
f2x+NXPjtInpf/RmMhYLjDc6gDSnbpeXUJFa6YyAsatJ7TlfGE0NguqQfnsqVaCE
kLmkr+68aESyblqMFl/IUGO6UhUlIH66w6ZgmiUn5+Uay2Gxp/yCu7XFg3LvQwun
n78g4NBwIgCLurjP41c+wpsntbWwt1yTVLEo/9hDDblGJ0UnKgWs+jbFlA1O7Jd/
Q+euB8gmCGULYaMGZAzLNkwZ/5ADSsDpBfWauYtSdIVdvUMTGxjWHlGaYKCHpcMl
gy41O8PFY0aGRMeebsgD0a6XJg8z/Xr40yKYtT/iaLOdbq+clAODMePTe1BXtN7E
POEc+hxnL8r6lHIOgk9DlMPdVuVHrgKzQtM/o489iMf8Tq3m0GB20T+K6HXz2zjz
4IQ8Q0uNQcFL9u6Uu+C0x89FimiwOS5dDj2VB2fqnHcJhMn4g/0ujD8o6pSO8jEq
oMwF2sunSUIhiwczJchnOz0zw6gruWIj/g75ynXfUnw272+qXhuI+4avBv+Rs09P
s/O5N6OTGOvT/IFZUA75Cg3C6ahyJWbcGZB31T9WO6m+q+yuSyE+bX5CaiIyPViC
/b3oFlQSCnzhCuos4ElHaQOOeRdkTl3lfsMcmKaJvXnWpUypD6qTZK5uMOvrnFkv
psrISWQs88QgoPr355i8hMkGu5fX+F19UrmrqVuRTgBRUu30Mb0SHmL98lJwh2V0
mQnvmObjDd1bOP/QDXRQuJBUT9xUxq6ZUTNbFnf7Aca8s1zYiRMNT3Odai9P+SCz
U4nRu+N2DeUckxg/MVWiTCQ8NO7RHBN6t7G0jAbz3Tm5KEK0UORaa1RZzTQaQvIA
gMcfBxEBmkZ+sF7Vf3rsMGzTXe0ZPjsb+7JX3Sb4vywrsnAgTaY/p7BdxXo7cVXW
M+yZxQzUTCfDF9q2q9W8K93uH3hA1dxRzwznd4VAmv9R82wKjmcHE0N9CcTwq5VT
Q+wxxlR6wG+sHx/ZN9ojIQvoK7jm46Q88jKotOMirOxl73f8a7f2eU/tsCNaFRY5
5UBQvuacvp5/uSF4feb/gMZr1uWTts6U7ub1S7zNAdD+Lz8kaHOERZiIghQjZF6i
scpNu9yP9ApuSIbr6ZYt/WNMZH0CyCpURQWtRs3v46jp+MR5nI5gmghZXCwYC6g+
HVu6t9m58KwlsO6CIXr6pqmqdMg/D7PoDXVEQcDvfRY4bw1qMbuaiI36PbCQE6zV
l0OICtU9Yze0U2VRm6dPNyCsCCQ7D8UM0Mnq4lpvmpuvPZQrBcMeEjklFzMArDE+
GSv+LpJv1vmLV1HwbdJdJLlEh5XpRnKRihPGMk0BW23IMfVBJ6B+VBATdSBy378H
Msnig6TXphTnmjxavszKe+g0iMxzpuc1yO9Aag054Xm+Ty1YiMwNcdf9H9wsi4KV
cV9rb13xEZXmGui02fSysCVjRw35HGpzTVxoKT/Tlizr2obY6cRJcomRagk00tce
E73corTQsdUvitZboHwoHMQaC7+LhmmdAcwkRHCpR6hzakZfw6U31rzdmuq8jeDL
Cju5ZlLpCo9WK2dEChiiNEiFUbSq6L/iUThf2XRqHUhiqpeR8php6ynJupdXYSfM
y6+lhtitDP1fhIrRw290pgxSq4ZfMlYwipdtjw6VDYmEEvcCEtkWd44sTfTFr2SM
FT/nUscwoXKooGOMddfB/no5f7VaOfej4gZTNzXmZ1ZB3jwd4YzEBT5AhzBIDpnI
RVECxwzAfM3Cu4+0bd1PvIQlvz5gh50pWf5dEav960cgpG5fr58oe6zxbZliIlDS
ZNwHW7VHkc5SqmVLQUGbYfyp+BI6qySrbvA3RXGEwvyH4AHrXw5JoeCVqlcpzo/T
2XdpZvVF/VnZ+M040hztnI97XKd7QPbpPiJRssU1TQswq1G+CKaqD1FOm9aPzyy/
sa4XNi9F1C6MH7z7cYGeRaTd9HjW3SBYHU5dGCc501uE45b/blEOGjuaaAyWVTn3
Qn6Wt93NhZVXzODUmTT2oHRaxFur0eJFj7eL5u22Eb4waKbBNs6HJMfGwxGlRdqS
99/5KqIt0eGY9pV0kj4hYZfpHQkrXkJrzsTojkSaypxqbX36iKOOdJ3Ws9TC9tR0
lgJHQBVGkvNnVwui5dPPBmYUvoK8oHEWN5gTgAmEt6BvK2h3MGabvZ+/GAQALeCI
fjAXwAlKTJh1WLGwltwx4vrNo75Z0XbQUOeGHcZtd5CGNZIrlhY1KkTviUQaF9U+
w57gBRc3ZbkNXJEv+rVYXPhOCMuv435w2fjjt6b9RP2nWm4FdyDZVpDBJiiLdt49
cbvedv9hQC8/ooM8FRcF0AAfon6a7XF2qC3F7kiS+ntGjmtFB5XJXGC3ly+/3+uT
qEraeIckox3vUlnAiIQUkXOatztwfePGpwGyVbpkht8oV5UldPsAr+/PIv9GhbnF
1yKXfRXKWV+nr7o7WtCOiLfJvbGlviO9YhPed1EhLi72YzSByvZ9GTz8Apnwu6oL
gkA4hGwiUQ7k9lsutRlwp2/R/mae1x+T9HQmjwp2HvqCpqckiVh4gu1RKH6YWUeS
TTSD13cqmKqzpqrXe13NiQ7yShThVQNkkb7lX3/dVyNCsSVGRPHBL5f8rw9Se4qX
+MVIq2nLi0lFw0NulZQaS177mU2UwHdzoZ1bdzsjah+uBbJrHJzbhiY2OFXQb9MW
23CJuaqC+UrdIvMS6XDq6K53K3iV+ichbuKd0v9MV0IdtmKLYXk0gJ3sUFOlhDbm
YnW537vgvFuSt4zHRwFTFs2eqmh6HHlb+bkB2P3mGyuaK9zp3oRVaQRFuCqu+1l7
8zMJBpD0qmBNlxXyOOIeplBoqoWojw3qVm9xdOc5hZKRu8/0zECwiDCnPIXhcV6z
XVSelZScOvwK/Xcda2EqtvIN2eABZDN4ZDaZqg7mxbCLV5QVjkaJtWfBflUrfAed
2LgYy1Ugt8nUpxPB7ESci1665gvZxl+vpJRK9vh8lXC6ZWJAgBHaEiJTD3f7dJSB
vdqM90tQh4LwbIzESVYkWhhU6FlvI0Mvij5JWz85RsQmXbgcgKGO2anJm95Fq5hT
Y179zzM/aWTnjVUOLUMOmNHHm5UAQ2opm0DCU57bGFWFmH+T6DhZzQe9AX2muIbD
D1k1v8jlrg9q6jrNsV3DC4EDzhehI0TB8sb2RUSXW49zfSE7YzkqW21FMZPOFkMq
s4CM17kIo1ATSvU7pOG4F2zyuWjM47++O8FZ786Wwv5x2gMskUzIzRIvPTaFg1PC
eMvmPsalCvqgB0GZndxOQj3ByazBHEziJ6B30YfmiSNvG3NmfJCkAjBDNIRc88ps
SQBrqDZIIQPgarW6G3zjzQuPDrgfV3ZPV2hiz6XThmDcUNDMuz/m8V39LWnifL8w
i4CCTJtNjiagP6d3hN7ptVbqlxAIdouahmGw5HelxDoHWPKKEQJmCY3om0vJZlvn
BYzmNPH4gnPujtkv25MkmwNgGUf6eK+9B+DcyR1PdB+45Mtdzc1zfuxzuia4fz0B
oLrfpf/wWKYV7ZVvJcT0CnKEDOfa1y2YjNHO8JtCLtnp9BnqXBMEg5979sbav4QV
kshQvFJPgPn0q7d69Fgi1XIkYzfCFGNux6ziYwwvkmdJh8VwomVLpTDa1WhsiMiF
ikAOV7hRZ0qFPWNSM+BdWTCrSMLy8a05TpLKx1f7BzJUJZ7qHWHTTshMOG0mr8dD
AqJiZlnB3h9Kr/fRmbBH3e0slioP6AJ+u8eHtSAzI6Lu99Mr8VPAWIyqo9kK63oc
3AD1VL23o17gNDfRSUbDJfQcHbNM+VJ3olK3QuBOGplJKEgeR5jjOnrkv/QHa9R0
Y+WXkmjElvY9W6AkGaN2rzN53vsbL9vsdGM+4ZU6BtVBNNOIyftImuvWDFRgkQc7
rNyZDeg/+xaV6OiBdjaQEGzxcRvDexmu8TXDni96oAFntQ3DfUJejk6OGDKDYBdp
GlYd9IPI6FZsUWHhqnwrgzZfBBSKCUmV0b4WMzce+S2HIxj5noY+84OoT/0QKfyf
PrBUZ5r5k606bo1oIJaIOsYLYgDSj33+fsOSiSGIgST3inwcbaoqNyMcKTJZZKGP
eiY9a9kH1SWliRA9mgOSEXSF+JtZ6H1ETYwwr8/H19ZyIunHsnya9+wm+2/Ek5tX
eld/SlKX6QJDL7fRe+yKZt6JOlLbOwBjlW7AqTQe1BoU82UWyYGk4plUmDfrAnyI
+Hkh7CQFBtGY7RJOCzWFO0F+jpJKDNukyZstFpLIZul3gg7Bz6yxfywEviPoW7Ap
sKuuq5sQ6T5gJF4KxWIYzW3RsYGt/WD1mQoAc/4vpWn3+9i1+ithCGKn+Gqr3XW2
AqilAo8DqvJGGKUT9lvgCXc5eDzOy8b1lGSYEXpYNC4uREmGnS7rD7fKn8SJWnHm
3udH0YDNMLn3YDXxxJFiQv1Q3neyeMmPHLfG44V7nZYT5p+1qVYHpyRgaUnR9NbB
ol9O/OU0cyMUZt2YF0v9CsbtXRGyhiCZ5IMR9POi/jzDc+nYkheYx08kO400OJVS
XTNcChAQqxghz1pLLQdg0ceiK/tJkp8KfYwzYzbpVhyXbTWQnqhoBGsvsvFCZY3l
ei7HNZrBdgcZ8b69dycfiZ/EQlnaLlIUJ7Sg4bOOQrDNi6iExwle3kM4oH7jG9Fr
7aT3CpWAnHZw7b6OBGtncvrLsv96MwlTp3eIG8tQ8dMMBC7MEFWiqVPQMp652H7H
1UVgZ/Vf6zHdT54svJ6/hpdAEn6rZLaCm2Yv8PbBORv4nZfIyM/6LySiTml+b8uN
pEPCUswt5sgu33tF7FhDd64xb147WxuCqHjSS4r6QgAqko/v3d9j0lj/LlZ6COxJ
WRFnq1jFRvqsBZMbdm/RtxCrw/XGWODB0XGfTHqOKPpEaOYcZdAXwWJgS5KfDxBg
5IlhFH7LIOh1l9KgSc3c7x3TOnyI4RNMGcFcs51CXxZunKm/hXnZQ6uek2e7ifBD
/pbczrA3r62qeYYuTMdcdgxG0GploYktRjNyny1pdJh8+HkVUCBz/PbAR1sW4gbM
+XUtuKZEPpCeonoPwEaaxvCT/FnRXkr24BDmKVX+keBkg9iGqATqn4BB1LnxIUd1
1NBGMYAu5mcqtFeqOnuwQuD3swVN4ZnwKdRjy8fCqPQ7b5CeQSAg7pGBPnmazA++
oU/roRTnbBMp5skiFun4NQEh4PCi+NdaVwXOUyoHVtDPvTPoBpzpfp3PofCVN+tN
bQ5yTAE6vQ87uIFrpPgamskNWmA5FYKfv23tpQnMr9ONVcGyPAa/UCreOmrrOe2q
oTP5zudOS+3p7vhj4VnveX4Aeb6N616UbGV7VxWzJ5bkxMGIlSW/FmaSFLynebHZ
3EGhj8s6BExY3R+c3SYTGsfDuH1wKBDeSI24necPAKMxVcVMZPXcVUXRST3HJ/UF
fo6siI7CybLz3Rm57vfs5lS+AV/3T8KEumUnUQcyt0lgImXEGQtjzVvY1Nir4IXf
dB3TqYmr4lRH8beAIZctk7hjZb+NwUW7AmIMLPTse/SN2l9rBmVGEQgxyfI89PXv
F+MZ2aQibF7tmgwF3T10KcPUXbZrtdgFczfUFvccoqkCTQ5mirxBiJzJiMEcxR2c
R+59LlEbWEyRwnasC52o8cqYggqIQCqWepf/tpCsaT9HMfxIK+ksESpJnoZ9WOno
/OwB/CMGg03kuDeZRvbncfBse2g0mLBSyo0R5pyZHR4yEBS/eTDUr+UdV+I0/gR7
R7dVnsmLxG5Z4t6A47/9NOBlGxtkccEwisPQQrQuxyPFs3YQI48DcQTw0GSzhI0o
b5TVvpGmyWgb38tZoenHv8ZPPbazWBDnJHy7uSB90qUvhAmEPt9rBFW/8GTb+S8A
4jA5gxAD4B3ZQVf2eSvuEB2HGNZDkt7kMclZaQkzYB9GFctsCyuZdjV5WaHEDIUF
Butc0B/qXmD3gBHTYsRLZ82XkKhRAFE/8xJjvrFcPGXrjE0KfLj8ixBe8SpcUO+P
aX/o4Z5Q5aKa1BkjCTI4GFaHpob/JCFWmsl606exUYb8hhjdWGnJkpgaD605NDl6
oDLBvJRDuIV0WyKRksQFjVN/jXQtN4EvlA46UXtTpqAU46uAOiWxnZizZDSdRC6R
iaJcEwgkuCsKy5sSkjqKRSF96lrFCkpF+OoVDjnvydQLnlpUxiI4to/7ENrMzBEn
YeOeDx6/wMbUFMOAOIYqHocuoFpAxtXtWDRgbPDLKCstqdwE9aIizoWAqMh/cjTd
JPkfwZ7YmyVjqQ3WN6nJhGIpmhl+F8prQJsT5pPuLfcZghX+BIDU3AB/NPRpXf2P
A987QTRHQblyas8ajkd1UrUSlENIzNS4H3Mot8TEl+wpGBwoGjgXDiFEzKWig58Z
LtNjHMgkULJgpMX8qgaMnJmiHjmrVXWC2GVKDjMMNuHi+WIK4U4gOP/r5vaKpfHD
Dq8dw+BmKwwStzKNI1yeUIxng8F9QcmH76MKX42Lwc7w86fs9HPgX3UR9pRi0P04
nXEiN4x9EgLDMhx2NsB+VGWi7ESTT/C2kD1iB/ToO/fs8/Pq0wNGtl8AvRwPPAip
Ygi2enr03nl6FT5mejcuELjVm7Hi6wJotuwysTVGGk0Xnsjq2pN4IqLFiZLBiSFV
6diIgmBKcxvQioI4MA4fhKbHukhFWi9vSFWyXa4ipM4uYfaLvc3+Is5JBC+62YaA
uedG+5okoSdtA9D8RO23VT57FDt0CdqGMwX9pu+DGRI8lN8qQVZyj6VhqY+0rPbv
XH/MRUgY2neuNw1DVyf2De4IbTsCaHyceLhvSLIm1yZgY1X0KrMF/FpWjS6QXElY
dXtj4UQHUDNtl5UCc/mqpPZsRc7rwaJcIvBWukOKEMsAVzJmWv0K7ESJMxXhh9hv
1OTbrNFjD7hLFi2nHFsxPPPavEaxk2q9yYXVUvjW8lUbJnKOvSchFHlzo8442mxS
+u2/z+oFb9xm9sY7UjY/spzAQHujHbkPjCUArJkhXueENsfA4sAcy8sZturn0Mmr
WuiFFcJ683wKH9lP4UEA1j1f1HGC3AY8JuNraf+PL3VzY4T8GfSPVJU95jhF0FE4
hTdZibEBifa65XZhsMvf01GDp8vRKWWWkadFQOYsNtuI6iGWUkq+YhM4DjLS7i79
zZ6ECWcMlkkqclWIGEVPzYNPH6brQ2NFr3ImSqEFerMojflU0RW3+z/kj5kZ/zln
N/vUzF1Lx+0GaOGH2VwYGZkkfT3j5wQXFrM3Od1FJiEY52i3NoHKC5r6atHY4EjC
xNz7JrwUQBYcTHaZkY9Ply+cZj/leikNrwhVYGNrx41lyo0h9pKQmBo1KkrHEiRC
6lAgliQe8ab0dqbeA9szGjgBhHiBAdHkRVt7np5DHA6f3xVUvTCKpga0gKW01O5W
JTEmHER2lkwDf3CwRhhUstFAxAc1Ju2c3fwWjskMXyGe7MqXFCjLCx63jnIXhGos
CPWHs0dt+9HIrn0urpUFm9xBaA08nZO8pRFKhubi87m991v/pKI1Oa3vzlNzbGxt
ZLjorLw2/PcYOV8kwgpJN9V/rV/OGkZt9tgCDyac5r+JAo1WtNTkbhtupRDcPibW
g0lJ5Nf1/n/x9yoo1eqDR3gyOHW7oVg6dZ6l0WXQqJ+JTBy665DJytCYxNNXdINd
k3kZ7y+EZ0Cna62zFiS8RRc+HfKMSS3b6Xe5mr/gDIoSI2f+LQZStlJFbl+Sn6aS
40ObOupIwyadD9NgrjpVMOG6CpQCBw44sN4mk+8fmRE0aMBlRyNLR8KRf3amqQTZ
wZiOuDt9Klm7HT0eKdO1z4i11or9ESrXOUyDmceagv8a8dslGtbZzS60u+5RizmD
VLfO6LNeDO1s3eW1GYJV3Lsn9S3Iet/jf7OtW2HMLv0ZM/YpodAbNJYqw1dZExir
GKDDygktPlYZPN5zme808THwtIkuP6fVHmDkzdIM/QSjBu7E6xZqrjGXV9NRmTYw
qFfcWVJm5t5/GLbvbToiA2jeTXvtI5TbNsU9o3gHTX6OaLyPh8UAMXPTwdXZ8REb
TEcA2cb9v2d0L9Yw1bOL2bIEFW2MatqAogKachT8jwy6vC0Kv9YxWwLZkb8APc/1
u++pD3JcoxXWp5PjuYQwluLKFjUCBT/iQNp/pedEoYyPlgUqU/Pj81JSJE1vNMRj
0OYq3Jc1G67tKITL8VZvrLWxkm5pMD558Rf4NrXcB7TBsuLS59YoTAqJtFhe5q48
FfwRKJE4bB0yg/w0FLobH7gil86H+91EuZ54iTqwd/ozo4DhvwDTjDr8AcBr2+P3
5lSA8ICZbOf0rVoovlPuVIHaUUosY5QIozBxofwY7/X2x1Yl928MZzsDOOtZf0/D
g2fxi0097KPlaM+Cp8BpIau5JIU1sOwv61Q1fkYUbm8T059/4Kost9i8FgHzBEcs
1rPuQEnti82C737pBcZznvnWxKNTcNPexZ5ZSyNbxarMa32X9tDyjkyo8TSF0h86
0/GwFYFKXY6kvfOXyLxlf/AF52oFxcpKgPmlyj1623rhX4Q4EKDcH4R8BGjzw8iP
6kn26u0RUvIBm4XcR6f8VZOjvgnJGUcS2ORC8ALCZ++L7yr7hCBr53wRrvmI4YlG
QFzslLYyAwsZpqVpJmTFRxijC3OG/FZaqpVoDQ9fczdRCsebgxn51IoODDzZ9RMh
hljC1L23p9xCeSYK4baF0LR/KFrIoS2YDbtXVeo2kVijjvRPxrC1A1XK3rcdm0sY
7WfEJri8AZzu5FM0ChNd7iTH/vu52shQArpDZMiwikon0Viq3fH1VrSag7iG5LO3
iVQRJ2cVdCpeJPfoNwWH5Vno+lXiibgthNf0KUN0yC9aIYXWICB5pUqJtJ/bMKwc
Lzw9eCR6cBLoCa692lPwMvavZ5+CzcWI9j5Gkmw1mzFR0O01iBwH9dN2U113jQ4n
+lan2i3z0nI8J8Zo/CGa8+PB3cheLZRefHTPIqMFc56e62Mf0F8PVsT7JL3dAd7z
vuz8ST6//0gmSLdjpZMR8VEZ5K4jStRjJUpx8Q41LQHsJvD00cGYPFsjbUkWo90t
9e6vE6LI+uK9F+HOILfK58VnzZ37K8JrZPenf+pRoUO32BLNb9pGhH0lurLTHYMH
3uDG6OCk+P6cvykB3VNHd3CkrPQ/jCd/Y5g4kN+9Lvt5mcKFQDBd+1tIMeEkgs5i
g8LOp8lxv3WTzrYszDY1UWDZKaxWjKXMlgP1LLYwbUVc/pPy3+eN04kYo+RFcxRY
fduZ5pot9SGycuKN/AGYv+sZWG50S4de/TTnq7oa0oAUbdqkRnacNrvgHEr9vFY5
ojozc3sj0AuxZnCLIPVY4fXyLsusBsPAowORtxLwMJEV3ndEOdgt1lmWYFi11j65
/wrMR+8/LPzhMGjGhcbArHuvwhtQZI8gt9gjdxI0d5vqhf6/eO4agoe1G1FfHcVK
8b0NE5vR6y2+jMGNHx+molldNF6XQxMzzVdzpRrXByuqU9TshFSJOONTPsN69ztg
f9fhPoBIoLCrjW6p8YuIcfnrhA60Qi/w+xB8knc32P2KSSnNunPQWGctGrJX0OWv
9RTa/C5hMAQZ+/jduyBAsi0uLgNbQNZcApsQ84xxU/1Xb8uNxNooorKwWXCxin2u
d8wR+ldwNRYhYorWq+uNn/PBFNg00sT/U6sxpo8D/kVb9ng9vZLt5AjqpQBAof+E
qtv67S0+NrWaWaY8kPC0aGLS1aTb8RjYXDsUehDBylv2HRxM+vSEw3rNFRiCv/he
UXJW3jk87IpS12cHW85sXlJJk9qjzzXRZIGpnM+9th4rzdbvAkwfectM2jLpZqWd
H5B77/ALdB7r/2Tg5WA6gEhXBQYdbqDsf4Ns+35bJoMHHUmgf0uhYzYFLFj7tlJA
KF90bwO4IgpjBFSBsn50gGu7l9dBKMyEaRAfqteN9+m7DAsQJib12cw2m00po3pa
u7ID/4RzHe4K1hD8x837/Y1OO12ekQOpWP6JB6CNBeVpjTkpnfzSbBusxxYCt9hP
ayed7/JOVFwsGyan0Y46Lbhb6hbJJzV6sd90TVQRrTP6Je7KWVN2RIOA0TTSZFgr
ZedfMElMHx/1XtS6C5kttT/qYvjT12pgXsXliqKkr5qjnck3Tz412aNs+mWJ+X+a
0TfnXlzeBh1KXbbOiB9v3TwaBOwC7cke7UGxc2f2I2r0tWbG1fNZTy2P5t+4wrvw
ouIZvSOsVarU/DbKZCgQDUMagFdlpS+hpu0glJcdO1/+ZqJpQR8H2h8sUnnPHnjL
YgsY89GdE/84hsDtiSO/Oypa35y8wJoe21yuXAUe56tJa2ROYDebN/vuRfbySYZB
13Q+m7RUhsIlGnZJNIut1W4IlapMU/jJPzK/MuPc7/3kWj0F+TGQ0/8qFqrp4/1S
2pNpT8TYQar/YcBd4aHJJUyt8QYmrihCI1bn6DMN0V+HJQuLkK3W9IwdNcyr17Iq
dwjeUQEEQJrLYevD0HbmT4OzF3rr8uxVFMFpeh3Vy2ZsxcrxnEfjg2Wr66TTO952
8C1TLaAD542OHhX2iVvyor6mpAWsEVqPK1rs3Vh0E1f6zeRbYz8gctieehdKfe9Z
vWz+6XDVG1Rmn5hzQqNZ+On028m4zTkzW+ahsFiid29g8tIs/OPEB0aJB8HoYpRC
80za279pUM0alzbuJhlEkkW0FDfkbrZT65IPq2kwMQYQVjPzEBT/YQvWnBrtGMs5
0cxQuK6f+6gWX0Ty1XU78g0btm83QnBa8kEnhV2AOtvBzAOTQEb7tHx6xGTH7FlR
roq77RbFe7D8yOZ7yQSLgd02Ww2B3cCVCWrqHThp31h6oTBFYh3Zi46BZiGnZrvv
2ZXvrjCLvC333gy9SSRLedCBhUiH1YtaruP4mRY6swRmGCJRjHutPWa1DFPa4FNG
/KWaqeraBE3N4Pkp+bLV6AZUVhJ55uqFnERb6IRw8pmtQGEZZ5qAayDmuXeBKIXD
`pragma protect end_protected
