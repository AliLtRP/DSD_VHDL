// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:39 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
eIFbUkUGNAmmW2jGKTtmG+PttszZSGEuZjF3IYqAgjqOKrlXZU4i57+Rj1xlvn0Z
jeDob8Nzy+x6FO+oGv0jgUukjt3/WUTn8PLhWoN8xvo8b7kSiYfnLioMw7Ut/9vg
d2SZp6UDfj8ehhuXoioqca/PEmGwn4IRwtmrUC3Ng2o=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 26032)
lgoTcYW+ByBy/3forjgaJvjWChog8T91Dt/1DhgiCT1ZlnWd1sU1XeQL0M+z/H2C
WRNP6+MSAVdfJAzCVGhqRX3bKnK10qeiEYKRce2ngKqmUDnB5ow3ksBF+2lDHybw
F9kDJ8hMlvwnuK0q6054vN2vmXKgjfxXSj+ZzL2W6pMXJxPuAcAXUHQDB8pafCN/
xLhhbtNyRvWydp0lZ1u/ioO3d2Ukp/lraJX5/M2odMGnMinZWG/IYB30EHo7ZXKa
60TO60d7C4M8G1TC7GWLlXfjK6k0e8/KiHLa3pZhdJ1YgaxGzBA8hdnWFXSc+OHV
glRbM1Wh2dyT1pNDit0DV9eAN2Dzt5WgdHp0zyoq2p4l/ZsDRw2uIEKF9ItRpy0V
ohQ0yIXd6A5obMCOFWhsE16UbUQfw+n9VaoDQR9kJyxLquxFJdg6eQIZICUGyUno
w0QtbGh/K8VQ5qo0y1lOmXDO5pYNSCBENwYcMuddJxODj1S6CrQUJcZk1Nb4+ThB
MhAOw/DVQIUv/79JZkIpEV+7McQ+5jainJJkyx+1B8FAr95eH8GlSt161aS1nY09
R2+CiDCm+dqPgewhUfRyLT9zeTMRc5nXP9PyMQ3uadUUWJ4AwieLF0LusLmT6Aux
8scBBUsCjJ7k3Tz2F5ybOsq1pmTYmge+gZDww7G8bYpBN+sMsl2CeVclRxrnWdXk
XRfBYaEMZ7S1uNFaO9VfUgFE6BkPtyIXhcYASR3i05o26if5/x8LUzVZCo6XKpNt
myYTF4dRFBp2/ltoz4siCTiizGRVuZeJ/jYkO3lcpXUC3jfxUprbinsUvCFezBxW
JNUDWmTSPY+X3X67SRDFC50JvRI3P+0LHpg2Dcc01aTcyT3u2yG2LUVBXJXs9wKE
jDkk3CJjymTWi7ro+5zK6HflfXPI03U1Z5wTvH3+dEfTTeSt9rM6mVEoLpUlvLja
dSI1Mtx3Zq1L+8MVRyt4FOQX1B2/LNUkHyOr2oo4PK7eJ27ip6aL+rV5lM8q2cyP
iEJqLSeVy4nOcXy9twRq3TY9l+A01mHWGjoiKBlHJJ6q7Dzl3Purp5C/K2U6jFP0
RV/hpf5gJLzbXlVByGByLEiN/rPaL33DyNRvcv95ndxnPnwbNnfSCidf5wDCuZis
50mnTLy1UpOpjkwr2Sl+Bpu1I7w9AygXcBrK1Vx3ItsVmXZvrluBdpnv88t8PtXq
vex1Q9aG6SH0iyOYcf0xc87EShWu0U2smAtj+4KNZ6CN7muuKanbdhNUZQ74fZkO
UGahftzywpwmOO6NWWjjWMRMLgw5xeVhpJFGj4jdki0sO9gg+pcyorxYBzYr4ccs
04kGjqqzuluhbIgYZ67Cs9cwix0MHUJmkWDwKWlZtxuxIdAES6oIz23ipVoOhTOt
h9ye4pnXvpVA/e2+rfvnzcMt5R5a1N4tbCfKgXj8yMsDUP9V+LS8OS7bce+2gc7t
xYr28CaMUEbA6zfZyQG1brzTv3ZWeq2o54kVs4iUAhtvFZ+rEbqjS4jaEFO8ZkSr
RvkyhPSQPJt+V5ZlY7L9bNOQ0CSMpr66ui+2rQ7TbkiTFid5lZQPX+NziuGXWU9E
fqyLShgiLk7jH8oWRMUbPJ8l8NyOXi/TP2fZlI8E++FFsXhzMz0nbcjpjNcPkZ8N
ghQFCoM1VuDR3Uj6r8CxMwK/tnR1gD9/WvM9XWNRavkIZssvRvhL29uV2sfmj8m8
MR+EiR6AJkUUWCBbVS/7fz+COPbMxc4WANzw5xET16potf4gZ0MCs3vxVyMZH3IU
weGZoPpyTklsWTJTuFyLD9mi3Lqb8kaSUZPwuYsGcVJL13hNji3+MlMExsvf0vJ4
RKj8PK1QXv3lVGNaMSIWVNaVl+DkOoiX/5+QGzvuN/icaByR3Vkbs2AZWM0Pjhgx
p2y7fZJgZAYNmcYj6WkHxR9eW0H6Re6Thanswn5LEKSPbwRpedw2ijfmLL7kHfmE
2q4M+BmEvNvIur/rqQ2pihD9XeP6VwzuQeIS5/s5Rz9cJun0um1MjNlJ07mbpeQn
maELjVvtYmEmRw46lgsvTi5nMnPxodZh4eS62QkQK47w4LWxKyuSeaWUgs60QBkY
Cpr3WyJMKZRIs6qwJ3f+EvlP0rfaBFuV8iYmt+ikjZl4j7IHvgD4rNn72ar5INaQ
euExhdCzMsL1deBbYBzmwZBFyNcQozlY1VsvCMAd+GJsTdJGCOz1EnOt/XnzEkVl
loptFr9r/dZ8IYwY5gwy3zErqRVe2+kbxDx2quQszsTWXDDr/WSM484VmIX+Qj2Q
I3qS9+Nw+P5vKf9K2yP6v97OinNZKyjxPQprsZH9K4HNIAPQNDVXBJflUKT64dNa
zaIw7yhjdOKcdauDPE+UhKKzGiy5BbyY/9PG2O5eKTeSbIOoKhMsNTuW+Wtce8jS
XuiFRL7jSGw3xH+gXyedj+nJAREoSjcdLYCuGANbeIVmZ+et5F9ko5ffkyU4Gm5r
TBAueFNltx2/3JYsE4AzNV4xdJUWP+6jeh0IhhtHJLdXeC59tgBnc3g+X0cIktA+
8JD88QrV7CGqJrvFrXCWHyhTJO6gy83gBrOPthAeL298jBokFVeI+1nxhvdBWOz0
JRPYmqBybHU8XubOzB8iBUO7JpRZ0NVNmA+k1C3wPjVwjZ9SFHxzUMDXYDOxf+uw
r6XKA8hwGlfwgMmeVCq7eZkthbaca+H0UcWFdil0kIfIwanMgqQ14DFdDeShZbHg
kdQmPTKz6MO+JMDXitJkkA/g1LxZ4WUHnQ63OTFbCqOrE4/6Ph8kKOgm6Q09ajIr
ieTG5tj58Bfnla6xw3FFy3DnfPeK4ExMmxSs0MRkDIucaZ08i7vzh9YfmbaTH0AX
2stdrmFpjEOZmlf9kgPwoBWy7ZM+svSduEZSlwKCbfxaEITRNarVZZT6MYenzpYR
5OC64pzC0q83pZFNoGfUqD6ix9jvusVP68QEG3BHbro4aBtB/QbPivt3aEIwanVi
cc54txzdQxVhyy7OIO8HIa/0ndZCrhDlU5JOdhgx/tSSap2jVnAtA7kRUtTRDV9s
SuQ0wZTbsNcPJIF2KM2v+nMP1t/XVv9l4V8t1C9uaeSQ/pqMEXlLIrzdn0UNm4HW
34RA9rVYHBkrXb6C8Q2uhgWHbR3/f51EUL8isZMfANGGPWaH61R7Jn9x/vHN3kn6
FEQ4ZNZWR4a83p5p5L1yByiJDBZ4kyvq3cuSt4B2PQMGg+NFSjc4T/ZDskJQkKQt
LXdeopj386nuSJua6ACXkFnt6yUcGS3bXNwnWIKKMIgcwx3buxrAYVOtOwVSs799
fd/ffF3LWWKxwza3FdH/9p0zl6RC92Nz0CUHwWZKueQx/rdFZXXJdgZ5k98ODkE4
+3vxwp4SEO9td6WjUAZkBig5y2nQA4p1m9+5Ex8H05KcjMupliQJr1DkeFGFxq+D
8dcMKpoUArtr3bscfN69+t5JLdt6TV06dujrvJVYRa7IWu412rSFsp9cWMd5WVXD
OkM8SQcw3+kfKOlDCYX/NkdVmrkPdmF3WJml+r+tz+YxEnB+/aI/ztTijdFf9QI8
V2HMw5c786tUX5/N/fX5gElemFPGyHM/MBN374xf3eOtB4QvAbyHUqQQJyePnFQy
FichU0neWYGF01fTwKDO+Zufzz9t5n0z/uP2rCpfjn8+XNVas/2qX+8OoHS9Vyg9
2ZBO8CA5z4VNHa1TqMYfEuLHtrIHVEbwbK0TwR9tgbeGQ+GL0ds8iYIS1+cXbliV
IgFDh5YfAZB7YQLwEz3QovCQPApZICuzeNn4ES16V11RyVaqWa7aaZjExkS2XNVY
GZ4t8w/cCnswRiXQs1IGJvwvzqGU9T8xMChWcXPdklyEdS9SSXHU9R+iBkTfP+lY
aKLwjXr269w9V85NLqCNM+A1ARt88TBmOLF4SOUldhom0uf5yl7rxTy1UKtnZUPc
2chVIcVu/9fJ1NL4w7asj19xJRyFqPMGIkqniSL4tYyjeQqTYcwU+uZEwLJw9HDR
OZBEROALWDSMEeIG1PJcyoRe43FmAdYcXD2Z+3FRwSLhrCM9FgbVV1epoFCJuzqS
ge6ollY7ZiotepwcC/aTIp6fM+Zd8TDLfxm+mCxqs443pFnjO+GZWsbSy1Hyh2Tf
vQN0vdh3zgPviCIYeX0d3BxSpSL9n5z+NUDkaG2ifAq2UhSkOjZseX29nHndQpxJ
PD9WQ2sIh05XGt7OgaSErIPf5GQvr2zKEDAZrqG/g8RD40iHubimnaS3TRczmseN
7agQBQFJJh29CSez8cy0108riMScH4ZXeE3hJiLMq5WuHPysOUBJJuE4Qg4pc1bj
3wKsv+OfaiBPgK3WL4AcKj3Idp/o+Z/EwBkxOteDKhqxDsC3O1xc4wNhkCa+09dM
hxCVAIzjoSUejJcDT1NEx/eJfgky+IrvioB1scwhRrcGQxxnLKhy3lpFO2I52aZN
oUCDGGLxJn34T5FSg1P9S7cADcDubjLd+8+5K6UX9pHqban2bAebj1lQuewInr/O
DP1Xk0TNY992bA60lLyMK77KWAoplcEv6jhP3V9c72mPGCppDj8nJv6viKDpMi+V
uFm9UDNKpbmUmeKcQonxUrH02gXX2cPZ5c/5HcleVPtM+cMHNLabx7EhY8U1EmeM
/zZ74q43UAekdlkQ0wSAv6wJnt16YjwFw/GfyCOONTI1r78K4+KG6yAEMfI/IkoP
ymSfZJnvtSwQ4gVbrfltQy7Lv9t0tDYYJCwmQesI79tT+ccpfa9IG4HmbAZr61gU
TKpfa9lKxmfOzYOSmjQV7wai5HfdbrxrmLzlO3fXbNH0MiZldGbIDAoq4mTg1fx2
WDQVA2POMg2O2DHNLq/ZGLCddTRZPlA6p0CchLvcqmSC7zSZ80CczsOS5SaJ0BAm
U8My/Dt99HV9CG36RaplvRClMRdqH9RT6AiZAHX3iruOfgg9pkmgSO2+K94QevCt
u6l5czT8h18ySMalSq2/jFoTN+sTJvlV3n3edbERjX88C0OqBTzYQAPsUlnK4BeI
D7Xw/aeKF/C5dEmBb5P/n+GkRbgtKBbmOzcOwguM+3PPwIa5QsA0MpxoDF5wZs1c
VLkirGcZ0tzbguorzX4YSJahnLFguO9N84hthMGZauuHUvE11IxLC4KP5DnBi7Xk
pm2MQBrsE8p7lJEbLq/mONb7q45aYopQNDVUGwq6l/QISod7QfrXuZ01nMdwL4+P
/nGyy3aFxTPY2dEyBBCeXq8KgI+o73UWX0Ajclf2Uvr5XM00mF4PvA4EBsXUVrYj
M4z5rldfNQ0CUslGu4nxTbedbSEMv3H/VGMSaujQkrfNFRBkOx64jhp+doYaUAea
jCvkIZuoV879x7bGmMUjirJs4w+AmsunXxPq4Cy28fov42aEC9y4GWaBEHVP+IUI
QwzY2eBAm4SpIx//f1sJCUZjupuxtYn7ajHc20cuqBzqL648iy6Fp+ao2jHjEInJ
C2wEMmiyx9sDQq9B0PWqidJcVx547eScC9uBgUhXaneapxub6LbYoXW58xGZg0J7
ICtUa8zN3Zt8eezBuEElXW4iDbpCWyPBE6itHmPATs2QEiFyWVepG+w2BPWl1JAM
3OtxHOyHt8ZSRXCbInumUsrfPnCYtIYrc5/3tiAUg/2HEW8oCuHTieyyVN5aUkdv
iP5auJJdmsiBZHj2He8Bj6FS8AJmhyp/RFQxNppp2WGpEfXCwJnfsVmZ5TrwTCgZ
CC3P4Sq+3eMhG/NZ7okhwObvq93/WvX9D7zbCMoekbd/kfEzAQJFGoYBrSgeThSB
wQ6hxiT1Upa+obxcG81HCiFojdW+4EcgnWLsCAXg4blfFLN6vMM5JXtlI6M6WyX4
30gKn9BnP+cYXNJroPYVrsUylBmfWBTf2Sick6Y51gqIVGBQFkifMGAstQcFXMGJ
aJGZWZZ7dsH6K23u1bYkFOVQbW6vP5KEfc6+7qQH3G/xbLfMWPhSYmT/dGYwjesi
5sHljIQq32Vm4pdrGDXvC/R98iRfjjujs4YUG7Nu6mrbUIZonRjIPzzE12MXxPoO
bg1soRSIuKhBcNvskTFPbx/hI4Q2cVEddatKZ/ToOGWpJ3wCeof0P725k1lldmDq
CqG2l62eSDLRwv0sNDJ6ikmXX1Mgm8OrVBehrh8cLCXLpQsKtIOf9czmJ1oyteuZ
otNprLFXn3GZavVlcqcV1uLai8HEdUsIlr2NipKAZfk+IyJptN25CotVy0gk2AnM
q2vFj8hkRVBmHey+XVHn6+fCsH2EMP2PZGU4YLk3il6RJ0UetuGOd1z17iXo6djX
1Z3pf/p6ZTy4ChdU3Oq8CmdI1AvcRdH1GvmmVus6XYmZU5qWyerzOsmK3u0VFihM
FsWI7AA3O+MF7p1DCu+zjnztRh+laWy1+o7BB7GlyTH4DKnUKBtt6xWWsZCdERFF
IooQt9bjtqN43GqaCCdXZzl3FBHjrMk3REJAdF7/SCot9EbKKC+zn9XYdcfmQw+4
eCZOE226MP0dxzpp/cSBMxIxfojPlFAXo/DR4xIroywIMMX+m7RJ7Fb+XoxnwEmD
6+su3vjpjYqdrCAnq94bdA+vX533DrXo13aV40mT01aL0gDqu/Js428c7w5rsbwK
QKB1PjcyZUvRo+hpp5rW0njY2SvlwZ7F9igMW+9w+ODDXdl1SPUKsm1gw8th1Ylx
k+wyWPQpeHqTsdMVpZVhjOM0RgeECmfp5+gCQIvLMX6s8mJrU6OJn8dEDUmXsKWL
j8uJycIdxXmnarusRkfIQ6OdSmIkCteDXGfaPBlpNY6tM//7pwc3qBkOG1/XJnAL
PJe1u141DTKZjDj7LblAQT61tNzUmkTNARwtQrBpIIkMng/RGdOSghHB/DV8xsac
pWLBMpj5i4DKqOl76LJ/muz1hQRzE+GYfjt7ItYQTdAQx1c2vLnru1rxTkUQz22j
VwZGVoMxP6d7NeWfimyhPdyu1KefL6anItPZKW8OdR3PqVXq1crRnlpKjFi27aFW
j2qqL6Yy5YNyFdlRallZR61LyLtizIt59kjL0vTREJBWyiJ3N8eqqBcqOcjOr9v8
K6er1nd/EK5iNMTTFxbWF+OSeC5SO8rCir/9pHRvhuhLFha55K7PtE5vHjV8It/Y
mJzQjmb4NCgaeUsYRvxMq8f/ZETKLxzZhK8XIfYx7ZeVB7ANbiNRNYaVwR2u9sOp
S5UM2XL5Netgix8bqTLYPIl/wveX4Rm9MYsKFBdL8xg5xigDubbIY6sRg7BhEzJF
5rcyuA7bnvR8ug1kZNaDcLKeRsz68f0vI7H7yjQsA9RhRRwX3JXRzn4n51+SLod4
ypiIxngE0yoB0rXP+yPy8KmN8Ix6mBnYZe3jv1P6GdaAuoNvJesTZuBPSsaZStSg
akjxAGNDo8Sjb2kd6GVgHetX0M7vscMsX1nKS6o4yZrs8vGeDysmug70j8jO+mIX
SKWBmcKHrdVQAIQip8ouv2vBXX531LnLqUxDILRcgzAvLQf7yZzjoFGacKDGNHxp
TsSr0ASDmlN86TvkiZr6CU7qpYTYEwhhOt+b427mkxNUaT7wgLxslnwanZKztT0v
ERJEyuJGgpIINu7pSEt/hynsGeM4oEkjBwWERPiIoN0ryz0O+4xqkdJHgo4W3l6z
9NoSw6NfI7cs76GkvvhqG9Z/k3C/36rof8+V/d83aqnb3IneuLG09qRl7oRTHI+e
XwF21EM9beuWMmPa3TFExbUPRIYfmzmXsqrr4im8ldNfxavjS+ofWEfq1ILexOIj
4WjFx+yXnFH4A+gNO64QCOxMMxe6coTN3RJnHTV6AUZ/w8J113X8RuN6npg4if5p
U3FAB5meybFRZg9uGpj8RYDATmB1yNwS4seeAoWm0pk0ynqozX26vCMXiCyBMjDL
1lw6LrQDON6aNE1oVmprOUY1rSRkH6nuZu5eDEMxc76WwQExhFqe+em40jlGmKyD
r5GBlVgbU9aYICcC1FHr2SuBZkeYA8su5dfE4fdxCD2AA1qRHo1pmQbsjqIMTs6v
HXNep0XDDJ9CCHcI9cFLfwPGuQhGfKPiChKD8tFVsVYAR3mA5B6kcOmIAhtmEm1w
I/Fpe7JbSIxZmO2Rp+OpCFw2fTCrp8v3mpvZ61AdOOE+pvuRskRTnruLai+ntEFf
p3imqeiudtpce/fv70o4ggE8inEwPaPQACp7khZHltF8Md+9yV7o0oPTIAbVqc6J
uuaiNKtL23kHhETpf8Xr/OBD0G355ebrY5v/944qyhtYEfrz4Xw5xw3GrKNEUXID
bKViATpI+EvAxzQgQ5mi9LFx7d1iRlhocXFhW350/iVCAjYgGvqYpNp4LSGesp+A
gCIARUQmiTMj7GZnTzZY7cumqJONOkhsy8LhsZqoH2BnvDObse3A9NkjqKkCMILF
dUW0b8K6PS1CkHaW/8S/oqCLL58601+tr1ydmudxr5TxJTo7/ttSdrVsSiQRyb1L
NB+NYgdOWaGhhGnQO+zpSopBYI5G+4o9czRUNaWvVAP/y2AG/io/LQO+vFEjZbE1
toDe+lIds0ulf3+ZBs6S2EbYx+IE3c3J604/hwKGMsv+Yz12l7KCilEbj7ZlGYMs
xWrvAPe6P/u/6pvc/rNdgto7fl1I2Qaud2t8sYv3aF3ZQAZjpnM8jS/Dg3r0HkrR
1hmtGLQT/kV/6qo7vLfh1ommskPm34J6SJGvuSj3jB+LQkSplva1MdCkATORRqsm
SIdIrDw/iTJGeml9jHX/rzuxW+XjTD2IsB7g2n8cHSgiscTdVO/Aeyj45KE6LDHm
bnkRrf7QOpViIMTgDsRvyGrBxxCcZSdaf8zV1i8IwgNjLErHH+dK6rCK6N0hY0pZ
dW4ZJ9TS+ytrSk5iLVf5etiMFpYQ5Typ76FYWHxOPjc7IPdk0hqxZeziDojSB9ii
RgjdKs7S+R4kHb5PvBALCe31by116qiUh73u/qcG1z4Zxlhy9pEXPRkvnGlyN2cc
+TDVb6j+3p0kEdSD12LKZMXbgsByAugnSsxRL7qqqoD7fsi9UBEJ/D1wlHP4jo5v
9YeULNM+F7nSToDNlqxvW8a24WPs9g4WoS7DGUpyLeLeU87Q8olna47joHhqKrbu
ffHu/xZFDpZsdjr/BS4k4XVTz3/Ia3J9XinuCCc0iaZxaF4GALNu6t+e8mYmroQV
DDxK8LSAF9JZAOl1iPT3aMOuYnOxZaaMwDaqSRXrMyhyW5+ZsVgdHGa22iOPivP0
eUHReWcBCyXGE2WjawivUdIbh4WpJNyMC1gVDcWz/7ofYp5ckPxeT0haP3bZhlHD
KxhNpIxqWW0Vos+oFo4uTCbTQQDtVAKmo/rCwe+brUAucaT57CNub/FeFC1JIdAq
q+gy+d7yOGWfNgaQDxiKXgSA99YRXIsvJ02WxUbDVCt6UQRdPNvQLZw5iZWRbQMe
WJ/U1JhTrFlXGRSckgQkOAXyH7E2x98xn3JGSqFXyNuuyqvZXXEcjAbuz8lJGVh7
PmRSfXGwQF81BKoYeTEBBSFcZ/vb68BXn+sRf592SSqpmsgQSbmfXsbTmt6sXplf
XNLlsQ4UEOMA8Jwob2bTeFWQlxu29aUrFBr/nll09jx8v+1hAORMY6hxg5u8oqHS
FpzJQtse7Nry53BKx4I5DBewUbgbSU8q7OyGuz81628L5x8wMm4cSlknMEzfwZ44
EPDbq0VUEzNZxSM8DT3Gink7Sm2dBpsR1ciqazVYYFOmhNTVDynX7sXdxQ/crE7D
tbFpfaYKBYNy6x4VeHGUS8HAAPQJWaozV5q1ib+cTQYHHkEyyTb8SdYC7etG8Um0
ruJJQgliPDCUFZVQ+UWRhO+ou6/m9KvRHnJ3hnZ2bytAyDjB1WYg7/QrVpqbOnfj
LO715xkH0cYPlB2zaHdS4kILHDsOzUOa5al3j1N3c3f3GWjU9395qm1dAXxzu9Fr
WbrDAXQMZXrCaOExzhx3t3MF3J1kTj6XeZtYUkA0LC1n6Bb1vFN4me4VS43n3O/Z
Hxqjdc4ZgzXtjFhCHlyBZDmHxLfFlMQMKOtkP3kawSVMiksXOLOtJsngCpM9dCSg
D5z2+HubphCWJ4QgyNwhhR6eF0iyNpkK4FvXfGdD20BIqqGu7psUJLElVnzgIJCg
bR5+M3TOVJOp1RWLyt84tMSa4RGuPwiR/rsJOCpgxs4dT8jAXVlIHxGCcIIg6ECN
WscQnmOX18nazP8UveDltsYmQ9+kM28J9H8XTWsKNBpZBpw19Q7dIEtOIiuT1T5m
Y0nMHxraBTJPunO342t1u0kbG7Q6mgsILe/86Ws90tiCH14BreDcexVDJHO0a4P1
QYpm7/iAMlZLq/533iX5+A0zKnU7p8yayS7inWU0/AIqo/GFrSSnfopWuKN4GNPm
CXKGSYr9G97z6E4o6IzIUK024sFIoqiy5q4GjIYZq6USynxN0C6kk0oGe4ssuJqo
ns8Ey/ycQHNUEbNmH2iDLOutcLT78C65E7V7IHaVikXvHAfbBcrBDvVY5YZkVILL
gHy1h8iT/mQ4I4PRHnAFUjdrf63Ip+wpZYkIPjHmjESFzxrpV5zQQ67ntsLHV6xi
22aiQQBZUVamZjD2Qm8WCEWlXTw420baPTJtQyIYtkhHxV2cc466yFjPQxgW/Z5+
7HfnuarfAbKrNBmJRA+3i+/SDkmhW3pV0YmQPblnvntoDWaYZ8uo+lqoOGosKCEQ
cm/fiMPlrBqqCmsgNVkpZIEsZiTc5owJpOZtaBzDS1klP75u+e7nAqlfgKMKGXmS
LU/G5NzsrZ4WTUn65TjWtE02kMyg9c8OCPvEwtuNTO8orjpkv6FmnDFnytbHRm5+
2RmcWFfZoRfKfCybcgATmHan8MOvtATNqTtO8145a/GvqT1Vc5Gue9rfRkljUBsd
dGAZgE3lGyM0x8hqsNpfUJLyS0bIAmAU4spyKFgPk82dZc/jwQJ1MDmkLAbvYmcl
kR2MRPRcrH8aw79h4Njc2wIMkZN0wfubd3OcU19zMJ1oy3E05etoxK26+1g5KeQf
hrwwH72pzxrnDqNC1qzGukCwh0vMTdo0ym69YFpn+OuXk9/v1v4JeYTVgmdJtdmY
B7Jh3+Hy/HaVoKfFgCUR2L0OXhvuwGIZhcDBmvJbE6JopR0/nRi6DR3HQjrkBE9W
0El0Wlc6v5SFBJgYaloYbdBjymSR1UcqbNQpWznj4GX20eaWPqS2LcX2MUL5zGRg
KdEN8KPlnAUg26SjxZ9Wa93HZni+u2cEInibXqcRqedna1RY+L4ZYlH9ArLbYN79
w7lX2BZJnf69fvDsnSBrgknOgy6KP7hh1akN33NqeJwkkhFQ9kDJKc035dJNxwgC
TPMIymz4xV55LpFeaaktKy958XlOfJiMCtU5FNFeBsjV184ENyOkRG/3DHf634ZJ
0kuC8jTuGzDPVUsCAIxaSIHLYF40E6Up71W0M89ZbHfI64GJuxByfCzdrTUlFP/K
9DItiAv7mpNTYWleRmQZsMmIV9ZHJeX2YdlEGpkvOMNQ/L+bq8fOu7xUg8kzKAwz
t/QCQ4WuvG/a27A92rBChyThEgrAD9t0t1NiEtF5klF1269SMlqYNuRo2P6AuxZA
W+wE5he9qxHTz2XESMdBY0PVjIkY1pLPnIFxo1yjxBtkq8a2g62QDwnfT3I53g5K
kz9dOri5g8+M6bMW1ENRpX7vygfJvOWbd6WLyDVzpeNbTcQOTVlbt5Ktstg+PTQs
gKmsiYZF7PG6y3yv1/rtn2gbX4UERwPOwdY7pKtl3w8mXaa4W59EYHKpHRDzbVGD
2nSE/MZ/xtBOHzqpgnHY0rmqdQKXx8fLWDdvngTQaMVePSbLZqu9d16jQIbJ0pin
/FutrLURhfE6OPyWu/q1dQTnhDFrdkf4fUH1iN07zXyZint0yfBDL0HNhvBoAdH6
WiHg+QaKS0ugCyxzXTy5ldpu170zuCEm7Hm4/1bAODxt+dD5drB4kiKzZvEyfM4U
MA63S4XW4cK/2V7EuKtkLFwSn0xkrW299vwgUP9KtuLWW4yXBZ/0LYxF8E7QEBME
169ruY3rwcYuD9MagKHPuz6j9rxH7DBISDrfel9OG93X2CB746cBZBJOYY51Qf5l
ru1L+cBezJXivbnQF1KmNmvaGVuvyM2HyHjBC+/ZF8fc0w5nc2lUEcV+R2oAGhk2
vDv0coBD/ewRq57VdhCpXiv+HDmrQty8ea0NtqdkXOwn0mdoIkf/lJqKr7pWOt6z
0bKD2pzySNPBU3dax4ULX9FQcixNWmr2I03antA8eygPBlrq64/5xQ2zryK9OxqX
EMjjDr0DpqsQf/X6M3Ew2KmKltiynnentltm2S4Mbld02v4GXTRnsDhtC6DkIzpC
NcQ7EwhamtPkpxLCnqsYW1jhF+zO/WeF+TOnqHl1C3whzLOwWYRKsNAaBi8vn5Bv
f4xg1fkq7MELUmtrs2iGLDspDkJ9Ll4qV02gT3Qf8v9BP4PLvoE1p6l0IbYmMqSu
hwduqrDDrCcFDkgMhF+52dPYbmoXdCUCJjX50Q/dFjNlAlz0KjOfh6bzT0lSyOs0
f7WdjFP7GlVUxv5BURvHS++4iiT7keIgJ9sU3idWAQStyGYq3Lg4IZFK7v0HJLGv
R64qxDUkuRCVH4i0jl1Q+MVJJgWWJckR2P8/sEyqNOnu0jboaDG2I665Aqf8at7e
htXm/nwk04lesmS01U1jFjRTamWp4dDexYqE55Sr9o8cN7onTewrVLi0XPCUxzlP
Qwn3zjtWnaR3J27W5pu7LEbtH8kRjcL3aOB/q75BHNa9tkC8yW8fzxwMFTykCbbm
z/4kUlKbJPUP6WrTGFADplq3eCJAHpFho0nDH2MK3d0xio+wPoRjeaexlNU1aHZz
NWfvqVhpODBNdvUElvOVzdrFcGpgbWwVx0rklo9idZ32Kizz3DhPqUPaH7PXxhU4
jRVkApTcfnJHlBY4lVvYJ/K454LW0oMtiJPbXO/pO0zKFlAIJkJnY84lbOgz5uCl
hbJq5p7qsmg44/6wdVDVHZmoMm4F1jB4lKT4kVSiUF/zj1fqpfEs9NuiCNoses5w
IGrpCZUTCXveACaDJ7vwsr1icJtfFW6beWlhJcTrVq2TMZVNgn8QJhuj+qL+s+JG
m4hb0Ro+tw09azHRS1s4qLwsg54STkKcnkOsJfvrPqwPWvgVFLVzePKY5Ta+/LuG
LLavl+zGhYRdTg0GAUtF8jAC5t1Wmz5Wn5rxSi1tqDreiMauRZiKwxgDv54Vioo3
5rPatqF529GEQw46xSFbQjT6LODwRf8vnddsBIBBtoiYLTzRKSJjN3oA1aSyUulK
bJorr4vwznu85zdBlZu4rWMxXwD5bucLarSciSSqLtvcnrxT20b+AAXnokWToGYI
zCRfrxqj/yyXlHPT+SFPm7dK8TNhfFz9ejMC2tEFBBWhX0rufVtINCpMwKaIcaxt
9HfJ9rI6Pte/a7Kx2eB+/dg16vcdUQ3uLJ9FqrGbjUH3hVW13Po1CDXkntomGqk1
CafsUwfVYlMO2jS2evhwLjW/wTG/K4q5qd/Hpv5ReClTGIBV8u73QBys+jtulLQP
k309ogXsucYRRXp+3k5hDT7cqMRiSV7jkKKrPxeiodr3YQIcokryUYzU/nca33sH
2Qzj2HHIRVXc5vlMA8kGUtDcFBzRGaWLokA2JksY5RwtF8dWkjKuZjhNWCVvXJ+X
mRJgKXHGW7YDG6Z/oq4N3Wh/h4YsT7H/jVWIVIWyrlYLYA7YfMV2q+Xmlm6abTtQ
PRI5ru9F5RJXPFuC+G2uWO4a1m5xLXLO8iT1IQSzlZT7qrpZLAkMk65uNwNT1Ar5
sitmdYJXIAYImvV03Rkism4NWuxWuksBWhTGbZy6ut6nm9Reva9pBj/PJ924CBiT
9mor6kwchpksEmdTGy1BDeOLD92fok+rFZBR2wZFvfvyqMv8YXEUG4+WuRtPHYoG
pUGits3AsJ9XrxW06Xtlvm3sZq6+h0N2hZxpBTZ6ujww7c2QbQsuyxmtx2+PqNaB
mz5EmpBT4QIC0XyiGZou2wDW/HdsfPDcNmqHTHSH6jw4x3LsRmTfKwhBzllaZIvu
QPJx33qlrbmf60lXmzaibgP8f2/mVI5WfKClFhdzhoqKcgSZFMCKRl1poQzWqDph
cZtEZAAMCur+Zx4gFjN4CzJUX9fFZJR7Dm8soURg5wa/m+Q+VV+6ff20gu4qG7L9
HNtdqOYaHWT7pyvutdywztEX+qdepoS12QxBtHhgI3HLeWTu6beY4EVu6Q2fMUaf
gJY7F1QNZhdnCBt/aHKda8fb85Of3INT4hVyn93xtWAM6k4oKoJmPz40T4yOn+SB
T4iDQ2O8oY2Zt52sd0NSB0Iw/wC2qd+H97RX9w/A1SJ2uI4ibYCO5U5Q3QMF4xx5
/DQSx8DlCe44v+F/PH6xDROH8MryJ9+A+58e+AOizeR0X/DHUd4xUonZsrWebrBz
v0wJdF4oorQFnGQSyjwtjpLvDvS/HvvA5Qa77IGk1d6HWS81v6GXC5KacvY+Z0RO
kdCbhI/XMOM5YNAlcZJNampoNVnHZbW3mDZ4er5OejuXj03buc51v1NcClzGi6I8
Wwnea4/1LZ81Nm/LroPPdvwNetebg6WOVA/BIve9R4PM3IOrjH2MX1Kd8OkbsJpH
DQs10mBzyoFCJlpZRmXrZJfLPX/+WajEy46XkxCYBLuIi5ky/JE1cpmLPbHbFKD/
k3PmNvvOikZZO8iBCaP6OZynbQv/4R4B7HAuAb7q0ZpmeBfc8wG5FnPZF/HUrEad
WPx4+j7TMf0rbks751gRvAX0aZqeD1zzwAzD659oCpophPnZYvkJ7ZnJ7hUJE5D5
dekSE0y4djj78Hyd40S4EMsF8NByH1nKqE5WU8VU51dj0oPkz/yj1TcUm60r8+6N
Az1rX8x9y7Dp82qyJuVjZr6+onkYE66AY0l9sm6s7mgOsZbvo0IrpilBZpn4uRtE
8eT1QfyMaMmqX0FS7/JVFNTXftIts4+cyG9wY9FdZOLSeDIT6LNqyYXKiTdKpSQa
NTfLb+mIT209wXcUY6Kw8n3M58BoisrrknU8CQZJnKu+mLLr35ouPA7GddOJseCC
cdzQdVQJRNU4cDCA+fD/OoON87UaAFAQ+HuUIKsxlx4iHEEGSwm0HBlI/UqejLya
ySHkyYllSx/IM1CkeAE0YAAGBPoOP8PUxl1b95fCjtSqf+W6SkBWlzUz+ijr25zf
rYEb97Q00xzc/5IR8QOTpb3zTmv52p4sASiEpCHYCQ+Vh9ABz0jbc0+1Cko3Bj/7
LZWoJzFZeP08MUBStXMFL7I8NdqExrI0sgKMC0lBCOqi4gYmT4qnjaRO6z7Kx22q
bLbsrmFlMtcN3hqBF7g4wkPwMVMjU8w7UHkHRkaXNVXw1as5zbXPwf/2C+PykHrd
I9phVyJpyeNhEKhq/hkFncgfGBr1U/0bGayqSfYVoeDU6TCdOfASOnDLWjmRwMaz
bW9xucTFAKF8h0/2Yd5ZaI+Pm1OqeMtwJt2l1KD5rBI02W4WLimIOFwp9cawg24Y
m5j6ujnv/S2GR/ZuccnTmW0HIq61FQQX9b0ZiqW52yp7pAGzciSM+oCZ9zsOptKS
55kLFMUHzb3bhjmj7wVCX9xVr4u1OB5xg4wnPbgtigdbcl9s94xP4/hSkarkze/f
e5lyV2+Sl+1mKzosG84yxmj4DnJ2x+H1/OtpMic1aAFHMHo6nn+B4Y+onxqUVEgx
jkP46J2dMxDWxM7vc1Te30ZwlvyGsohn7yGSfcMCMO8iKD3M4wljYtgwU3sYocQk
p2EEKUCkbtOg9I7fx9Cj8SIt+cRwoYF4ra60Z553arKb07T6Z9av7t2jeOJDKoKR
sJgXM8kZeQ4Jji08SGn1O7oQ1vxpt6knTv1PhroIHKDFx6YtagCCWOF04zRVWE2Q
nWsRmg8XPHGZFrKU2FFBSt4uUevSzRcy8UfGcwa78r3DnfOnp2rdLmDM/RF0j9n1
SESuZ8zUd+xRuo3jQ8UkjRKqHJY2Llwzt+ed3wUmDjSf1SOI55Nd8JcNmWqYb1w8
zhI7rLA+UyI9i6lt49hoy8VI5/sE2+r3iyEuY0wCjQlDe17KPEh0TeL8JSB5OPnY
cH/qMSEIHmZijuQkUIciDYiHzfERNHIXDdp1+drIrVVg1IgRliK7Q+5JaFHGbJpz
5Rpo3E0kAMWK0qisHGM5T5otUY7XGODJQm0tEu1F/skul+bApLKKorYbWlWzCoXq
5I6Qjia4w4Bdt856vNJe3iXXYJKKFp1dos1Cty97jXdfYvzPwPnt9cbpKQrB+gAU
yCX5AjO8p1vH2Od0eLTXUh4OYvxt8fUWpbpM2OMQ7frqDhqNkoxI86S+fiK+ct/w
zQNOqlCYMcwQ6Osk7GzqwzFPYJPDR3V23lmj+OO5CnvnyQ5crS7cehBgLKfF7rso
7mU8AqeOIb+ac4DdrC5LmOLfUcspv7m7eRVJFPSlfOrB9aSQsKgTeL/Q8TApk/VH
i4rOnf7c+uXkuapTgSc9PnYwtw1No14sEf7bm/sAvmPtWdkRNGhsiKwU2yFQ9D0M
PWhFBCrULqLawQvWxq3lSiTYhwMAeIQLLmPdaivLGYSu0vwSDOSi7P/SvP9+CkT0
xLvxbmo5+Z4YrcOtkf//Ez6EdG9pPYRAm4tqXkIpz8tVFMi6RBtaydM/ynzdDcle
YWqQ2F1ZqnOWdjOOCRvDCr/XV6+Cl3hbFUJvcXhK/aZaBdjPRgUMHnCUQiQ+FtWw
zgi4DxqlW1cc0MlUdDVNGrVUFcOtldSGiPPLxmhEfcOoRUusM6ehxTzQHSCqbrlr
4gjgfs2tQSJSswFXweYqdExYAwW/6YPpf/wu4US5QVY2RQhMLiGchew1gIXFcLkU
zfQ8NF9rusAojjdk7AFuzvrX14NBwgnPxDLLvWlYrd2qL+JEts9iEh5+jcowvk46
4/eLteAH3IXnwC5hnmYogmOuXakXvNafNt677yQYLjyfHZb1sg49jG+ziapKxqvW
36CxlAT+qeMZ5pCMjx9EC7h/boa4yET1zCp2E1z7bYKFvVUaJHwZ1yzAxO8JjWe3
BzGxyBwr5cLaaaDRfaJq5Q1yHpSHK/Oep8DLlvXRTE2uxmBAHQ9DoXg2Dpj8oq3h
1GNbsNi01EavnvfGs87J/TUN8AG1+pH05w3w+X4KIWlwlmFO7GgYYVfZtYd+CUoF
vTCOpQkP15/uRffhIUzfNBV8iGgkWVwdGxCSibvxuk+dpK+wwGheXI7oB8isa3eO
gK/FhoqDDwv0XfD/ue6Mt94EeJjefGM+yr/YafzU+kMraJR5kUtN5mcd4vTeWTzJ
ShY+wA0K5rpjSaRVCnGE5qbZqe1cLOEvwKHtfbhtQhGpMptEes6S5PJ+vSGhIzRZ
0hlb1Pr8W17q1zLTMlNHH7dJl04ie06kz/6OkNX5u7BIs32fCIiMA4T1agPyLuQX
nkvvzaEvBderVIqtENuQeJYvDPsBLUGyNWCEiX8C2cfsQtLi/0c68Hq8Fx60kcId
50SRbQ4s9bIQMiWqIum/VupKFWFcFHdzM8OHSpFTw1Mlj31sFhvgj4R2lGUHgct9
KWZLCKHE3MWOTjcuvlxZbr8kKHQiCmZlt8BSLxye59LT5nbF5TkBd+uGtAcAPF5f
ad9r9r6BQOQeJJ2PL8fJ1lOi3nqJzgYsBQnisQYiIvuVRrjw9Uc6DtXoh8hASsdX
o5iAlWCj8yYVU4wJjikvMvCdS2bjy859uUHtRazB65dAGXCJbTgSKAJhBqf/EW5r
QGK74daoLaSLTdEbrQ3ROf3NdjikDX5MbXTb/cmQjJKu6vj4sirqHcqzhcKn3UZT
7UR9mI07TyIeEz0MLelyMMqwzNYm7TTbUoz0kJvltAd5tH2FXSYmNCZj6dfy0t4+
RNzqUtOX0DKdbt/ZfASkr8A34k19iuzE5gx0XuIVTUozYdXr/BjQv3r2dRq1VAtK
aaZAJ1bV7ryoyvT8Z7bIQQdpZx7WvtyP6doPD2ae7i1kPdUsBO/DNIhtWdH4fXGY
pju/w4zwNMa453aHgj7kclLMbQaTriUiloB37H6mChabkSa5RyMbnbPwUbjLkWmJ
eAHCFt5tkCyyX0sl9f1dITA6H/liOU1ohZEtcDI3dNO+vsYgrpa+EZKHOMr6YTHJ
mGn4id01/f79Hvap1GedOslk4JIpZKJVty5PQzGskdVaWu2ttuVIu2M5cNGCA6AF
APFQVXf+T9y6FKu4GhSaM0A8pe7Eetvv8lozQRHV9oh/w7dTlUwAo8P/wfbjZFys
w2A6eeE12f/tkWrwtfGqGanfv1tSiKf15V9v1+BxOafLFAijjVXOEDrC8jpJ8ROC
/rPhsZAhEozXBYdHXlC17ryA1pZVH+xKV62LxkfcE+VDZvIkN3UnvSePkO2qjulZ
nuzQgZEsZlE/iy5VpFGa0D6uS0Iaq/D8GpH/g8FueTzpL6mcJHmeo9xy+NTReabm
CgWYy4tRQrtet95x8RobBIHyAH5Rw1NrS7kgJXue2IyEpvanR/VBlrLt8ltI8iWi
Ym2Cc8j1rkvhc5+yirKE/Pr22z8sA+R355QgDVCdpqDMS9LYdhnRvrS+VGzXKF4r
X7DNwar1pRBRnWjfJSc59EgAuFKutsSpTiaZKUeZA+Sj3GQxnwyIowxeHvQ7N3Oc
4eZmhr6AHWnuVwhMjEMbifYbmMxL8/Ktzb4VXz/RyNMENZXc85zskEohb2NLIAlp
NVmDUPepN8ojsCNYKtNf5Uq+w9OGcFFkozU5DYb7N4UjlOc968ksSCmb1eLM54Rq
eixrC0ODK3EimkZ8FDf01YYtBvhaNUiQAP4qH33ssYC3iIcyBSdWiHSoDN6A5GzG
+Om4ZlD2PugdzJ9mSxEvu5IFJ+7u/OLalZ+c+Ci6pqIqB8Rnn8neTQ7TmPngX2sH
xeRojHx3zFmqjAIv5Y7Wno0Ect8L0Apz6UGmfU2CTYN/UZQ3/qfBlAopRYRMjcds
P3kxmyy2h72TKkOEbEef/VqHbtQ7Ty9wzYyxZu897p+oMvUNCEcAFaEEsQHU46YQ
uQ3OxJG+vabjhA3Cn39Pvc2+SRim3NdfamUJMSjvAZo7UB6sYtvI7g7C3Hp76FVw
R9/0ydZUjY63TQhCEmp6v+5izjVHFdYEkms06WPzTCeUwqVrSFN9gIxQwKjsqb6b
Okq/VACO6TKbMEuwDnLoxSqYbrkBBQq8HrYX/rMdDlsl2udj4luK+MePEJi03oOR
gbarI7Ha9YgH6hKcTFlJhraMOfpWeXMz/9FoSoBGnbu1SnJWrjqzbpXDd/E9AwrM
yW37b5iaK0HTxAJGIV+82hm7fCpDemr3PlaG8F3uPn6/s3qV7j6up7io0kqMcIWV
J9HJIrmp4PboK0lnx0PzF9qk17MtJ8rqU7XVQRryqmFYLkuiE97qHweCyHKjOb4E
1Po/Eh2UahVdij1cvjxFKj4LCgdmqeEDbYcbI6KcOdZylpwqNs2OKbuJmztdDJIE
TKqas6mfj6UzhpMTuyK/QCnPTS01ibpDhNASiUnoYZnJIKR3eIfPgNY37NeXNVRm
ArQ3/tF2kn7+KBYVt3sZU/CjnOV7ojEzyTlnU5ux5vsClVIiC4aJD3RsNEUj0zgA
SOku4Be8Fr7p3pfATYM1Hd4vfyksD1Hdm8ifEVjlTilkeDpTAZc5b60pOyZ6T1bt
MATGzEIRiZqdkdVgvKULjGD7DK7GR74eOnH+sqPd4rI8FLKD3Qes8LxKtYNsLuM7
RFOJV30FVi/yJJT51VnlQFM4j2mGarmTsFXLew6lk2RgL5zVmGpM0LVC96afI0p4
gyMst9juaipbRrjnWz5P75QjwV6nJPRshq78iZzEH5Xc1/IeTcaeGqlZOPOlt82F
+sBhY92RjZl4QH5G8PThd68CWlKqSS2E87A2hUxc1ml5TAdOi0DY16fy9jcXW6AO
q2enaJcvLkahmE0QvAarpzBhJ7x0qWyafg2m4JiVoGw3Gto3ffdNUKBR0zQxhYfE
oyNcZeTWz/hiPKujqWPuLpRRy/ScuWsSN3mgVi6ZcSKAkCkLwe635LR3depWngtC
f+D3+yjHU2fd+BikPEV0uuILih2d3ccJL7Paeo5CusByWGPBwPJyF3S0Zk/GoTFh
/uEwOnMfcIctlVOwOj0qDqhUki3uOffza8NnwrMgyQ8hIU1g1WHVV7DpEsI0X12Q
5A9j9KwbIY1hCN83dCWA8c0Wj3ZbAutnsLAqkTvdVM6s/dBai/GRgVI/lW23l+xR
5xbBaZhhTJqqBvGFKXLBrWpy1+6nSbD6S5SzI4qUzXZlBYFQcxg1jVTX/B0BOc/9
NAkeG5TNC/G1y/DRCsCKxxASWNZIQoBUmW96owp1mA4cTgjwWOrYpGWcwVc9JpRb
C02aB7GOeU6FRER4sIcMFUcc9pL+GLpY1O4GqBBVmRtQbHAexrrmd9CUwd0/LciQ
huJtKCQwYnKXKUJKNuxVhQrouZAg4vZTMRRQYg1WVMGpphgrgPoCXnuEu5GIPIe/
NAENzV+MImLpVg3txZ5QwpoanuSbmGdLvYC4dKjI+UMZAYiUYZaWziuiLwxcLEul
AyhoQXcBAdlOx30+IazxlbsBRmwpmhTCri10sD6cebpAbjAXdVL4ek3GkgEcGcDP
OlSYHiyVcC5oZgO/bJjwhkRADzcysll2UmVMbuips24qIvT1WVpCsaQgTpZtMaST
xOCNDJSGI/3dbaF7vmqXSq+2g42hBFULpF0PAEtiEYEcM7nccd/AODf1Yk14JeLs
IX/32ceP9PmkiMvhg+nNXetH8jZmDRRESR3QTUoztl0aZ7HfAy1pyttLQrHseTtZ
2EuMoYdQ8VQAHEQLfHdLxZwX2yBNtWQ79X7u6297xkZbxq5AXmAyfvn+wie3oWrp
/R4ttNO2BpmcOfBUdotZzc69Xf8Ngp7Q7MKswoAcbqBLUpu+BOD77VFmRC+SXOWi
vCfnAJ7/LkQsrbRZsqMuMa4Osynj9XskHTJjq359GdjFxSKgzPTpvKtzsO3tcO3j
4rSpDlPxhZlFwKHN9XlLN+X4vFsmux3dyRw1x8Ab9NZcCstfHv7bPuW3nuETeoFn
5srYr7irq+uRdHXtbFq6BVqE9n3Q3ke7I7rCrFV0CFdijIl0w34NBzuM7k141wJC
5NKQh6ZNIGM4QkZasHNmNuCKmC9/GdnnAv9JMYHf+0JmvAb9WIIGyPnRHvemUXsP
iowIVZ23OZd8W8EDW4/wfhZagObQ+gUbiXGCUIQS9vaN/WSUKZvJ1ytMnLfqU2n1
hm9kDwTA5obl24jhRO6PVsD+I04raBRvDZkc/xbchaZ2L1Dw/OouvAsc9N5PSWwV
AAmPDxpstOUFoiB3DZz42jtEO/fUErUXrT7v5mhKqVcoIBNi4KO86zpX6Sy5aW0J
MVr7iANUECGJgn5iXL5T87XtbW1ToUhBHc0CpnzbsJwv4BwU9UFUl7uNGs95mCPy
QWOF1fQVsXAQdfwiDBHcYERInOXV49ngFzcLEz76WaeyY6FAKN6b7yTDPUyZwD4o
68gVpNiuKJ20K5rS4krVG3FoPTT3UuPz0EBmA/SIHFGIQ48Jsx/Kpo+FSLcjqsfN
DLjQ0JkjvFTwKRUGG0Bfa37Sy9fqZ5BVU7V0cu0yIc3mXO62bwfS3rsnG9P7pMVC
N9UNhcTAo7BnGMjEYEcns1u96zdQBfmZZ4tBrsdjqhE+uj4JIEzNBXJQ/oT8sPyt
mQMjp5B5m6RenQJYLSUX6eVeH+LfIG3H8o/WkDtwrZ53s/xvMfxk42Dt0kiEJNap
GcoqGkB8odpYJg3rmF6deLQuPxnEO7oIKFfMxTxTCsxabDhHiEqtRM5z4Nam5XNZ
CHJCApqM/KhU6V8Y2le+MXdX0dO6BBuUX2bxGqv8yMagGhTkM1yDb0Ho48IvL6g6
Q+IaoJIouuNz4xU6yqj/sEXqCeb8Xpk373VvJ3gEEa6RdlrzCTMX02AGQ6t8MCW2
jj25KWoI/EIviYiEMm3d4IXhQdaxzs23098h8V2DOIGAdaVGZfRlwU+I6/b+idsj
Bhjius9MM2GrkM414d58jQBhWuk5I2Xfrbg4hsTJFgVp16doB8o3RZqTQnvmRoAM
KDP0xAMsezFo+Vngwix+J03ORSFkVW0IOpvX0FAMKoZSgJ27jpN3Kkobh1avZ5yZ
TRUWt94YbgjCfsIKwcMGp7eL8KobsbP18O/c37PZpiJAVXveVT/YT/fNJHi73385
x3Uc4NWUBE4YoRm4Ed3DopuDWRCmPVlpCDurt4Bn+VHxJN41zW8OmkaqXJ9sRBMc
LUWdo3pLgK0H1qOkgcYrB8jd6PHcj1rw9/Z7EzNjoWzbGynU4cQ0RpDZHa23DnuE
TIsNfNpBrd86tzkxFUDHgW16s73oj8VCzfXLHjgieY6ozHxD2c09/L1PQMA1iuhN
zLjixDmXCnQFWPDchcBQ38Hc7uiuCUkrH3qeTuisqH/0JD+SbYvnVK2bPzkRCMF9
Pb4PuyNRF4BraguioexWkOIlDkXHRU3TnQM8o7Od1g/qoBzUCERlDrTodAADzyo2
hOb5AjOQ1gznZ478ZLJqMLqw2P2WN7zdi9Xrm42z8UIWYiUfy0dC2/Qi9/BEIOxa
1OTOaYivVp/0j1t4vF9Esd8bwRzbI5UX4OVylw2FJHxtUVPK739lBsVa41OfQf1Q
ZF5ldnPzrQn1baGTmu0wtCycAe1KufRuNQMLEvjGC8/GJ9SVdVdpARY+AQ3m8yr3
bzzNhzBNFy6M4WJUMRcaC1VwnlqSCb13Gk2XKa/C/MB3OHypQMBpu2K2V/fiJPj/
oa3c9aep8gPX0JAMPfJmJnTjVnjdqeDokgyzmInScKoa1RQCJLojXJVgD563Kk3u
RAELPQS04uQaOdVcRf2eV1ur2gcpJdU7ZvnALpmUq9oWov235Ted4WAUX5C2GogF
cMaQu1ncQO35v+nqUWWdXWg/z+OUZZMTjAQcw81ImTrrp6g7VA3M95xqHVamPOgJ
AegDpr6mQJ8s9KEr/F1jjoTMqzoUqHLfXerkMr4FdS+e5GPrYj1bDLPXkZgmYktW
9NMylABhcSmUNmj17OdIAxG0teWpya/7LfkMT2pVUcgQ7O/Jg8qWO9Kj6/s0ApoS
sagcBHPC8gufgIsgQKwN88W0G9YraBEJIHy5sdvi2g6agmDL2RW+LxgcfvtBSTwO
ZwE6PR/qFXb9V4hVSJrym/PKQbB/QJAwjQK1aZZZ3SKh5DFQXkJwBXTM+B8X7vam
s/TPO2mUiBYdnB4x2WGhCdDcVbGawMWOpuvvVFCvxG9xfl83xopWioC8ZAs/Dxb9
rzwpP+xjIjzzjxBxHwf9Ek3vnH2TRCvPNveldq8CJqKNXwHvUdHk/3kJb+YzVtPe
s2RjT8YNtemkajwweIpnHSi35envcI6NSHwGIqQ0TA8kslpL/JQZ1XUWqH/F7XEz
HbiH1x4hINhffUU6jP3c+fE/jAuIyjF8CR0p6soJ86+pwZthQpuGYLuPsak/cPd7
3tnp3Ck2MKWs6FxJ8hTeadKkXyoVgIWNyzaM2YIGQ0b/oY7L/ljXgRtz1UWhJ0w1
C14o7BlYalL5Z1DmQLrd7s5N2LMEd4iDkZ3By4CGqd8ehdx//lx/n+5LtwzkegiK
6hhdqrOgZMkbupKYIqB2RCKQYnDVIkxGy1U22EyLRC3lcNGBrDzcFfpN6H14iLl8
yGq9Rv5yrPODxRfCgXft305A/XltCspYHUfELSBqYcmkSn2qrsh3v0rYrmEOxg0N
Oh1qvHTvY7rl9RQd1yOFODQzNa40nY25xsKkHTTxkKnV/p8hfEyuKPrg3gXA8ZAu
P4aZpTbODtsJ6a5aPRivf+xPMKG3Vdh63ZVvmQTz+l60so1rTU2wEDiHrQ11jvuA
0Gk0OPLcaLoqVn8sSMBNQQdpy2bbZsDBj/GoH+LGsnMLwo/t3hPt11M1yqVViJVG
fQ+FtImOmX1+Inn0hIEJtiCE1L75lQ52yAnmGbT47FTVOYfD+SiQIbxiugnMObnU
XI1oFDzN1O9LdbUsXew+HRT1qn97YfwrTZr9MQMkxRNkFvnlmL2lGpwaNR0eBEqL
cV8XvjXCRCEdNacKwXJfchOjE8K/ODYRSanSWJkn7CUEXf7mY/1P9DhZPjluNCLj
6u6kJAfUkIfHnKRAwEEgmD6E1yZzAKbSdZeWrMVRhZGHni5/RyiKQVnDgQ8+NGuE
LoZXjM63J0We79PO5SnxaAvO6stnGJb9DLVf8Wz4+ENxAU9iIq/mqmoZ8qcTAHoT
G+q73wUL7sGMivouUyFRpZhb8TXKz0GN2UufgtDjH883Yw3Hhkz8mSXvFA+aOG/A
0NGVZWdmn9dftveyJ9uqF8QxxNxFtloZ60HqrboI8aiwAgyIP0vCiA+jATi9M3wU
LQEnGlCb3A+cEuw901iKgvkXoYmSOGRHfPitBzSbcSANJg+E5FUP0gfIYEMzeDTI
P0BWI3UCkkfj0Yj+cDLLjRApAym26Wb1FOHuFhjdLKo3u2/2EIQA+kK5iRIRRoH1
UqMnOgWZYBN7cK6sxL5Gbe7zloY6IZJGk1nQ6x2dBaoknc1Y5cyaUaUnyHlxyWMl
yUDvr5+z2o89utwmsuuGorml/uXEuSYb9bSis4xbxk2AtAWDoDdzMa2q1ma9Y9sv
sS5jmtCYyUYbrBEUHLchQv0CqFX6hWSPPKGQbgeDZhjWc6pCP56SGzu17cPaXYPz
RcE+FP+qYeweM4qHaK+UMUjGstIE0PKaIeojQMMAbsdAmFCqrmOytZsgMukUb15M
5plV0pGIkw/j+Cv6P859ztAXJ9H4XZe3fvPKwwlulwHM3pG4Fq5QsZQPqDcD3gd1
Gc6d4OKQ1kokzxgOMO+GH6RGkchY+1WQWr4B1IUX5c/XRxzVGsIOVnKoMeKG6fI3
9esFRL0hAytFbSe+uyfNdpyRNpGoTuocg5WFxl/3umTFkB26ETBT4xA2MxgO0BzJ
DX8aXZxsbimmIesGqCy2pkj/Txu9LFXovqeGHm57sd3/vZkCXctDXtWpCwJ2DUzr
KQAj3Vn8YL4Sh3YgZN4YYhu/wiEF/6D3Lb0fhRy4iJdUgXe0Blg1nk/pXB3Q5jAZ
4ycNWDyDYh1Rd9ENty2YQ00lvTc7WP1CoHVCD+GYDoNd0wUM8PCYDvn3ceHtP1BG
pf/ELpB5KN+aO2Gp+sLVHoljKUU6jeclVuTVP8HCLm5t7OyxfEW5ufnTt2tdWRFY
8JR2UAV/Yb74tgbeD8UIZbHu4TuoDKZa0WLubbRJSZLachJJ8YMU3CtfJ7sEqLdU
JXSVivR17gfXhwgpIGh+qxfkzepQcKzfKe5081ePQ6x5jcYZ5YmAQQUQv5u3swrq
q7GennrdFbj7R2WwySCMIuUUPNwD5pZ9tvtkfb3AYO3PoPmWll0GFiWCEIV8rp7v
RsmBSpDNdLE7VDgliDk+0S7mixnt8264LLo118fOlOklbr54lvqJOf9kiFx0DK3B
NLjl1ypQcO6dJAO97irrwtRYRVi9AqIbDAR0rlCbsD8OjdD/mzLHww84emHWGgvx
sTwChOUL22ulahwIOn2WG7xmfhfJ59boQsp/03pMbo/9ETX39gP+fQkXyzy9f/5C
5G0NZb4+sJI+iX6wZ+ZjyFwTYwPuo5Jw8hEZlUb3J4FctOzEzZX5H3p7fUdbu6Hu
yrYGsN62TXHOHhX7/ZEnDRSaicBY07dKSXccAvOBde2/Md1giIcc6tJQ0GxIShM/
7vV5Q4/wUMd1LAgNJGvEm3J2QFrbb9W2bEAoj27dp2w+ExwRYiPDK/92XahCtFl9
EX4ss2ewIztih/RRY7lllOupkV25iylmz5l5jyU85PqKkefb2MpqIkHOqD7VZQHC
FDTxl7QbjE5YQeJwW7td7ZVGCY8vhl+dayWNLNYucfEeDyK/b2JOUEGLEQmI9u8t
BAHvC3hJzMw4GtL3xTIa6kaVk8b11Xm3T2J65HvWU0IYTqg+5k05BzBwJjGeDHLH
kPgdwJ2+Kn/jT5yhE2hSaHGKvZqo3Mxox/NnsC86HL+n0K083EgSufW154A7zDRI
5OFl6u09LDj3THw4y0N1jRHI4kTGw4zZ2IDu5TbVtLj2RwRttI9Tc0J6ctQkroau
h2Zy+WqP2Y7Ia4Ld1Jdo6QSIt8BuCQ8bRVPS4BJPhgTHNDw71jknsuRNrL09akLB
dxvJYps8wcBCqMBjFvhRWQbpra9kG7FqLFftZXi/+E1fUERNczU12UUQTjsXbXOF
ESvrvuPAL84XUCM4T+Ezk/H5nh/OVSZGRwbSgxm22Xvs+pUBqbSu/rn8v36rFKT7
SFJ6aVSWw6PVV8TlIQfi8A1sLuo7wHyBEZZ2O/zEXJsT4t3qED1NdP225oEXDJZY
I6P/7XJ5jMKRVGaiuFbPXaOWAOd/zFm6+wbO7C5Pp6LZZ3kmBFCHp5BMIapU9QxE
OcjOOHVX6Oh2qpstPPQMhJjuCfx5wuuLVheuaj/tI0lO+tnaxbX9065ffKwShwWp
h6H+um4JiorxUHY2H8iPIxBu6yW+GMwhqqlEl+9r3L8VI31nMCMhbTBnE+C37Nu1
Yf8JyqI1r+ZBUoZ/YH0lCm7du3XA5AMQxzY9AI7LPN0PVWN20U18q1yNvj1ByCvb
RP9AMcDjnlNLTXhXXAu9/6fNZUNWa68ZoAVI1mxnS6Do1sJTfmz0iMEjDTOZnZcV
mlZ0l9KdzCwThQ+S6+p42zORLpxiEbjPdMS9PbImM+Q/bRr3wI5IJzkagmoVH8QF
pW6Ga0iit2qMRa+labZCrd5NVJ//EYq0ZAaaNYwGpYhLDQZ+JK2vudLS9g14pke1
8A9PiNQT4k5GCKLXw7GBaRhxwYVr9df4BCuxduELg31VqTzusXFJVNXBPR8IsQbu
yokCiyKwAcGoy3A0rNIkv/w3L5cqGjTcbF0R85pb/51/ieGYWc0G0a/7c6NwIHNW
qEugeCnZjBTqdTiJl9WpxMUXOLtIn16RfpM/DUEh6ZHu4otcV8MlDBuYyG5uAS8R
QpKzODazOdvXLup43o0+jNxO8Y5yHUHeBKlOkLRVYgwj19VSYu0Np8dEvbxIBu1+
HNTIy4fH56sKb6vDhzgZhw6weQsSLMGrQ/cJW7vBwX74QEarpSgWXz7x6RBX9hA0
J2DKcdqplLgaujNpriUrCSZZuyTjxhFoitgwHKOrB2SjAsgzmLae2Z/w0yjLzDcM
+mhLxYHRWXTsWbZJ1QvBkdwD88PfINBsHaau+SxT8gVn0MwANo2DR7qtai7VUavv
NYUPu8SSaXzXRHjQZsg4EoJchpjOFU0hqIJR3B9aJC59L4T0Z8N7QB0fAsrsWlQg
J3+iMg72afkPBD51yxs9yWk0JvxWHzlJKYOZ4T7225+t2b8HSQydGspoF8/VyQ0v
Ft8L2Z4F3eZ7qLH6gZUoO6vkS4ISNvggVMPgkrJehjqUKh52Dqqyp3i/2bOK2pkL
A8+UrYosTwWDKMCI5Yc0THLGcUbeGe5wK1sbVTYhjpivKe5vRPcyhOcVwjTAk7pc
Uow9kS4PJJ96vo2atcuPqCVCnZ52PTwiP+1on6tRKF7Wxb1vHqN09zCR3q2tkI9+
SUS4rM2MYROs1O8rFaUK/9Sb17JbSH0IIxllbxrCobBllKveOTgUaLurVreAHZon
F1MidKLTA2o8YSTevNSO3TCMX1viUtlMQzRlt+3TTJ6FfEom0NFt7Ugsj/Zm9vya
gMRRghPBnb815T7/Qt6a7Ex5V7M+mtf9z9gdC5Y1HMC4m0Fw73s1JET1Mc8J0N3l
9/E28JU1G/mlkeBHeoqbtjfGaPqF1EXtcDMnCGBdLow7lU22+DsyO19CQ/EBljVf
/h9Yx9sXq5RJApIQf1NR5kgmJosFocwkMWcXQ1Xctt2NJ2FwEXSZs5Mf0SrqBTJC
L+V3eV+cU9gyxm+RPtzBCN3cjdZg+tfq0nAX1in/YPjfs4jfKB7qDVzCyqDETmBL
sh73Xnk+L0Av1H1mG5q2IGRjtE+txYc0C5177szfLPvkAWueZDUssr66IFydrRaU
4bSfIqhlA1fAEWYnbadf5TnP3JvoW8T4ilW4ancDMQ3fLX05CedtVwm8rgBl0oai
yc+XDfU/NCsIRep6DRUqdHBHWdR3L+ln6bKBU5SZfIcyxkgpsjeiDX9lQl51vHSh
O6VTrEKbot/o1Gjap1EtC7NFiPrGn4xzhcIaN1ALHr3hlPGlXDEPv2sLW+GqJzoO
SPPqhdXQERk5Z6TRmLQ5r6mFJNtSkn6J/I4a/TfYyY2uwIhudgSbHseHdb/HxxVN
zdLhQlmeAYi5ye9/1U5SRZgTfzAgwP29VTd+NCH/7EoGfw8INl/QRlZJRM/Mdb1p
ES1v8wot92H0Wx0nMYDoidgivg/bO4xWuewkBbXLcH1j/L70OTU1MOJX8UTqRuuj
4H00apIudigH5R8Cdz3RrsWwNXz2oOk1R+vLjXCVM57XJo2wQIZRmOwBnrUOi7hG
paArkUiokoBvI+dUK1aINdK+oK3IWwwI+BUZgXuW0eP6ZFROTMj0owTM2/IevTrd
IwJJhJkoIlFDkf+K4p0QMrR389PwtHDBCpPDzY4Sj48GEg9mWvf6U4eVC0bRxMHe
V5zLXh1db7RPE2mgF0SUGgAi+wSPWyFpGJdNsORqFQN8ghV4u1tTlMQD9p/SrjL8
3Mu5wwvvF2/GTlkNblJH8jJ8jgV32QRYc0rTuDvE6v092COJDBKKnv0+MLeKyXPb
3TU/yjFGlobnnZm1ZOaSF0R3qCCGSvgZZGHswXoNvtCG8Gcu58k1p8iO3GowRVKk
k1WwF3lPsp1tmwfqiK7nRoBox2trfp5mQFoZAPtRuAPI9wHu780i26TBqQ17TfMT
eiGCx72/ghSYU7FAbXydf+ySSwkb472xmHrR5f50ZnlK2BVWbkAPRkPyFCwG8J02
NR2bLk17ymsD11J6iJpMdypYZpPXxrE7FWIroed19OBnWUH8VQnQfka7GJXzqtSi
I5dtCZQVP4NDwOecGDxRBUoi9WsjKKJhDY6fgi4/egJBY7ZsBYKQLVhOBwmrkQgP
sNpfTVJiuG5/1vBJvsZzsrb/IjA1VAL2PXLpvswOTnygx64BgL38pk/GH4sd/fne
hVB+hCozW+WdfY8D/Yf495lg9T1XMcbAQop755Yoc0TEPTK45BgSOv5pGHjzpsex
lg66tk8OTxwfCFaRpt3ZSxJ3hdBxzaI/nJYqfNJobpDB3yWYWTY/QmK+U3Fot2+u
0QbZGe7WqoZCsv93RU0yIM1prkqx7ec7Er+gmXZknA7mJwdfa6dzPwdOYX9v0lO0
Wsctx+Z4rRfdQvW8G0P6zjcaPe2X2xz91ZwNW69hnSrplsmr1VyoifEjhja4Ir/U
jErV9I0Po4npOKPqGLKNeTFIGkeFCsYR1RAqQlQaa7OrDeahWxY/5uw+Eo9hQTaS
K6bFL7HGPuQ+3/JjHnHBeDJbhZ3y03qqxePMTq6bLhzwh4r0r8DDN7fafVW5rb54
Cj7heou0sf8/wRZCmW5H7xhk1QI/QnFviqUTn5g5akjVox2oRTBh0gJqG8hDxKw9
1t8hYzRbM2qDxU9cvIV+9QJ0D/rTr+tLns5eAGC3/AG45PYJmfj1e292x6T3R7dU
f05QHPgubG5TnegQQIV7jPZnkyzIgLxKsCFkxX9fFZGE7RPShXg6+xsGVQZC8CzN
ju+RiJBVD3CA9F30JAGW9w92MREUYqMOCCFkJ4xPWx08Rf/NMgl5nzTYpOw8Hpg9
aDmFgWfHUsyVfdvV0+M8KrFh5/wjsthf0PYHzS0NkFhKUezttJfPAkZfgvNnyOHC
c6UNJsQ8ThWuzx4U3Cdbm9xLm9naVDGq+vPFrgILVlxcGjbUJXOjSQ2D8IOgG+ks
/4oTKMSGs7lwyjgfy7feFUPSqdOq8ZdhDUnTwZVaczP5ommDHr5gZ3Xh6sqr2UXg
xFT8geerUeRjPhnAhSW6bAp3crtw7+6UIuWY7ZexyJQMolE0pc8bO+p5MRCuQuYp
fcAh0vslnyV6Bem7PDKYG+26un2itmtA7C8zoMO+IEO8ybHuOb2q+goFo2EMZ/Ye
n3tTqWtJ01Od7zLxCzab7lxpTHqBIV8BRLzUmwDKN3LlFSA9hEoQlXvg+cAsc6Io
dKG4OqrTrPehDDjadWcDkHGvysH8nKxU3LqO3VvwzGkwWuMhacNCKmBtsTowTn2c
mkuPqxaOg+sIjplrtxA3+b7KX4MhylQ5AGB82C1Hy+ds2sgEwBqZiv88ePV7jp9B
lPgc1t7SL+ZMmUSaWUvgtltGWLO9FE4KVNx3Rg88yeICrvk2bLPFiHU+dHICyyF6
gLxywrxKMH4Upc6q7L8u2XCe9hSzbjPlNZypVmpjTlr6kXeGUuXD+EfV9W10dcXU
6HUAvNSw7RZRzbpQpY7y6djc9cUkuTGiTNelQaGdhIzeaYncvXJpZDlnE9nzzNSz
ZmQJAcuyLQn+jAw/M0tVtLCjoNKpxtSr/23d2ihMxLIaAL0rSWe47WJEiV5GUiIZ
4SLvXfJXIuUvvcf7G5es4vSBJ5A15GIZ8R9N0GjR+BnB7uZF2RKV+BHOc7GxusXB
CclC7yl7ZWNxky9wqnj0lBCTb0UVbCM+IptS/NDp8shTqiEDy/9aktMgzmWB9g2q
AnDACVpghA856mUVbLbanQ4rIzrirqDBMUIsXp3WhDHoov+ehqGHxBjdPZmmbVsl
OCvZygq890E+FvHcEOcI2bPWpH3wiWDlIMIVa6C4eahcM+S4H7ofq7GaMYEOw/XF
bF14O2HsVg37CEsiomZ06ZHsHchu0o+JvbW+DcQ+2VIldwX23dpUsAqrB37iM1WC
qmaG2JIK6Uc0jruiD/JBnRMWG5EIMruNsg5uPnNGyIqEVtArpQsWEH8LD6mYxHXb
JprqZ4iEpCeZhC0vlwp9mQLKDcrxcf0oFMsw1Ir4bMs47L+2AK4p23XsdkwEelJe
8iGta0R3yMhhS61z93MuPJYcoBSHQauPIpjiFMDOb3RbvicKSdrSpr1rldxrB6hQ
2pZs1gAv5wA1ta6MgdMEXKd2R3fI+aInS5DsQilhTHMeBynNoII1ia/isuxm9Dkg
7nnZUnRD8rpb+vo06bI4ltXiAlHpH7gZiJ8NEwlqg4ZkcvGkcWoAuTp/fg4JHvNj
C+rDCqPBBhNMJrM5XBQfdPtR9/9riecaP+0xusDEbHzmXUVQhI/YwWnKUhq8Du7d
77fl/Nh9oz6MVpehUgz2IE1Su92RiTJjZzk81wQ1nHeEstkiIh2BgHJPsN+GWIhD
IIITJRlNhNpblxDzzElGG93FYzchNuP+8f7OEcIG6oPV/sTbN2rfs2LzYP2lfaVr
YJqiHsX93h1FfG/MyiVOE6a8K7bLxu5cR4A0w2nIPbjfZONjScp/GfJWemdRW2t2
JWoxtIOZci47DRv9qwWSkkQfbE1WlXGjIk9nQEt16njvPEp7QvyIn7b/fg0l/foM
6W1fu5Thrh/drCRSvpoV0+QD/bWOLdDNuJ9iSnqkgcPjM30jqAvFh9gUl/i5ytPw
ObduwVfGikdtaZQmp5kh1xkdyQTesxguTujYXjI3hOfagks4zyzfFjQbMy0jukDh
nus0oNlmJrPeDc2iCRKh8lTjlGrZ6gE5EYphzQZnMMRsPjQ8+lt7IoZTUIw+J6JX
RFRfZrXJ6Tr2Yz5BoFBJz473XDa3EXpXOvX+iT+UfB0pmIh2zeCr3JbyDfuA08+6
Ts0v6t0gN1fRnKKPGGkFh1lQc8ltC5aYiXy7WVj56tw44hL1AG4py9o9hXkz3lZc
HFfZhVM6dvwODcOv6wTGSlKXUvfLnPxPNDgno6ocNLBbWqeQu+P1QTyYb2X9Svgk
LMMjN7OGb1gWF3/oMVMYMu2XBhNb5XhonjdzCKKFdKVMiRx032+drU6V2zLaU5L3
fSmRB9CK81lF5IlBmKx7CQkMYtJYa6FzVkXF810ZfreSQPeSKv/eWt2uAMRCOOcl
PLnMOBkthSa/hZwP6YavyMgX+YoVKYV96GS/Ma1dVWu5X4j8QYJ+sjh3Ubzo8cFz
Oh6j5sTnb7FyXSosqiWPD+VxafzHU3+dj3TLmJuUt/r8cckoSkfpINoVI6SkkJpN
oCdLUAjiL+Fof3P983uNmC8zcful1hwMSNXUwprcOZ2XtugCub6VdSL73wAKbcRG
QBSGcJ+dI28QWvdckPvTe59QP03Y/MXjUP4XCFcG0a8qA9DmAQOvmcyo/5zU+2Em
bXvkDYlNUH4sLIse4TePwsVvIOswy2y8IlWGyEOOvJq+R/vhqnfJGHh4sFkXv/9L
qweGAujrjGgRes7IJ0dnMVLTklEoCTkglUCGrW7XqMzZDQFkx8PPmtenTBn2ruxC
nSKmbAVA+bRtpMVikLKO0nnwP8mBes76ZSYpIGlvGAuOnH6Gk++rlOYy/9rj+//5
DugPcliUPPpHG3ScW6E3nvFHyCgFPvEqtCvf1AV2fbQASQdmCWBuBD32YC3Ndqky
xF79Se9ueI8dbw51SOx1y4poJ3z7lDh5e1Fft037RpecvNWzeclKXoNEJeTyVOsE
SzVwBwaYgbXRqOpLEXVN5ZNgeEJGQkbVV7eFY/4QwahoADR5PM+HWIffR3cUq1X6
3oaE6zj6CJw4oUFaviGAz33poKnPBs4KhHwIzjd7TMVzkurfk6LQFvDlrdvoXkJf
s067HQPYwGbqeEoRUDynasJ/12SyJZU/J4HP2SgGM0EBeKJPwPvJZdPAmCtV11zg
W5Yi7DBQL9i7750tHPD80Ns1B4jdbBt0vvMAUg3JtlXuD/bZwW3sFBWHzQBdLXvT
WkVof/hom/UL8fT9L23mb2YChCbFV3bVojz4tV/Gw5K3HarIyiyJg2Z45YeFziis
/VwReIa5wDFxFCwEyiwR81VA1ZbVa2AsJsSxIqPicQLHKbG1D6QiLhXYftopuwIL
R65tMPWIvZfYPJjpEP+4vrZU/1qg/D5qEOao8Ck1ZaLlfcvfh31H9VdaEGfcyjva
vjO30bvK5yqyV1CbxRBGpwvPpgtgb8/JohwI6Q+aWGu3bb6pD5ReWhGAbzJ4Ej61
IRtyg2muZZBNoWjzSsx4S5RhrL9j9XFMAeyX3vr9fbuTJO4s16f6aVneoZA6ih7t
O91Ifdy6GQaKKt+mGRC+y2B4QYaxsudvidWyGzjBYIso/4x9vUTBlrT7JPAIBMWH
EZV4u0PznmaClE6Fwh386jYqZHU7JN9YbELQ4DxFTo7SQERIk4y2vTJBdQqDYg1P
84qOrrqFbATxniFJuARrgzKGDXMERn2RtKG8Rb/Swvi0+UXBaOFMtfWlJhmqniLt
XPxM0ghihWuZAGmw3ZO/8JK63Yn7voBCsKgt3D2vQatTb50CkAUcmd2xW8Ef8nBm
o9kbJoO8ukJcwsbSUgOVCdwNYXEE2GXdF5LU0ULbyIdh0HxMLRVjtzMfsJxLnR8p
mpilT0PaxZGX4hU5rRGg1ZPeuJx9VRxN+eXsJ7Z+UkGOJzUMnI3GyouU8LHOOwgh
H+fYV2tqxdFk87vZpVPT0I026SVo7aSUiLAHolHWb2oa/1KSKZxy+rn9PMulFcMN
YuIdFmCiqkbNQXlyQC9UzlZ3v1xrJCZOch63x8xJsdWWJeY60t97U2+9lutRB6oX
Dk/5SojLOTKt2NVojJiVroM0kGoRmnaSLQBlgJbHj/R9DAgIFuT2yGYaBt/UiOI0
1cz2XUR1cVngWJ+Bm6Ddf+R58ivBW7wSIpsh9y2Uqb05dXiwUXETQTcxw0NHEcTO
bWjnGEWyF2N5pDLR1SMWvbWn3MsPXvxUB7Ldi/DoBoAXrLkAgS39fHp2WDy37Y0J
TUtWVV1FfBwKkmBbpFPzCv5WCkyaxs6UQ8p5bjR7cyqEJGKZDWz1ZAHbZLY4RIN4
U30QDKCDACdnFXDgl+tTYZ/OBIw8C0VIYtVxH+MvXFFPh8V9VBMeWgY1hDC94wOG
cXYTt5ftH6TwT8bogrcnTuzbh7CHdCB0dQf01e77t40Rrq2Db3Vs2seuaa1QG6Eh
9YwIHLl6GD1soE3vEgoX4ynILoSqV0teh+/EPT/o0MOtc/g6JYdlZgXXStDCNu0D
Zd3doNvycdjK+3vohb+fTMuecINkisZ8bixLlnMMRExCNNjkfSbpFn5mB4Drs0EF
MZAeBSx7yG2TfEsQUaU81N4IlbZQ5P196njRj9wsIbzdihnX6dEJBqX2WVk9C6Je
3QCPCpq2V6AKX1PXDr7COQcyeXdpEtQB6spHb6+uoIpPG4drh7iUc33iFed/Ab7p
487234xoV8FjY4LuyMOrricVXa/0tH8wMpr9oOMv3AyDiLWVYoAH//ZOxNIspZOE
YQL1FCNMXMism0u51nz6/1R6OhqCyaqeUMHxHwF3XHgB3hSR4+piZ/z71+EPleus
t7RcGWCCp2/YUZlFj8opT54Z/CuBk6NdCY+7OmZ3nRdNJqVuw5CRAXR6Qr8lNBYn
6kE3YvpH/EcKgp3eYh1xM+D9Qbjztyj61NSCEeF7RIieQyAOFcSKjoxa4OZF/2LY
RZpWxfbDZKQTMEDGga5O7Q==
`pragma protect end_protected
