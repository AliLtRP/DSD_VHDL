// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:50 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
bJb1lod9106qySme0/znC9xG+QTClLQ/rCf5FqURRi7ZSKtDc+t01gXBnGiYpJ43
QhhEiHIpDHHt4tFxntb6NJJMidSXWjK5KZeKKCCFdi0SYkjhUGYgRQjei8f/7oCN
IYYw51maww5Qjem78dTrxeOSRJSbFuPDZwQj+dhMyoI=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 8960)
hFnYbvR7auruASQhLxHo+Va7Ar4hblsCi8AWnhlUwhlwKWG6ZTGr+PsLMPRTTf0c
CH/CBfCvVBRVdWTzFIii2c3D0ejkXrk34gUqa5RAYn6Qg19DJmzTWzpC8Bu7gGeG
8wjwNvJbfVInTCqGfLU/QbTvrmlsTePIvE0mJw/eKQ5lvhV40vFqg0Yh9f+AhIAk
uTGfut5RBayXXbTuq2MgIDzuFFGgzPw8ITk7K3HJiiDKPeU0+zUwau56/FlwDM22
ONP+0ul7UT8LnZRn9NbVm/A3oue3LlamKJaZEDMVKHGihy+WRPdsIZjGrgjDinTU
L+ZWY9uFKHCPvnzhN8jvGEzPzQvid1/d9x2HWOTpbK2HW3BXyvHRG2x+Zm0fzjC2
cUowCYm0OEGh2hleMzM3Ql/MIhTy1zP7Hd+CBGpAlKvOc6b0jNLc28hjJmTsy9D4
1dcKnST7ti5h2TjKycWFIeLvX/i/O/9tVNQOnbXjXCWwOnehnVYqF/ZZOiCru5Fj
tYDxQQCObNQi2BQv7QF/89ExmeUw7T1ka0J8SzO15ajysE3Daf1kEm7TSerAW5dA
/JnhuF0V/zqH19azuM3EQo7/dtyfwMjFNibBANGcd3SKVGUR8/N2shQA31mf0M4C
69ozC0dqc0S9RvHYaKo6JaSoqSZYKMNAqbjs951JWYnTVGC029XJ1/epWxczUBZH
y3Z7cKkpiKWAJrXmveXg63Pi0Po/4Vraz2rfItFPH2VJJZM8oVu6Sy3QGRgpD+3N
8VJTernJNODEOkZVgMOGH/+gnFfqH4zIKX2aUrO/AiV2vkAnjFxpEoMjsybhMMvz
QzRPdglBgaSKRlT0LTx9RNBEV+uB515zvq6hfoH+4nbbJi8I3GCtNYmvXoXPTmv9
/DHDeiFaAAmWJCnpyTBWkjbbSuhjLBjNnjQ6f8EAvQ0XC60zP/tO5FrFKl66vbax
klvUqXPy2O4cGU2YfpsMlZTonBsiEFkwNldc017Ke1xfI5ev861P1Lmv6zcm+TnL
yQeBngoqMuutMB2rjJVZ3miXltLZhWcU3atcDA36Aoet/q/N/07bVReKYB/bBAfl
fQzxBBlEK4fNXx7jotmRMIcvagN/PR9Qs4f9ok+V0uS0wo9UlUzPeX5bRL/XY1Fw
25zuLi/A4gRydBWsnJRqMI9hH9fjJwSxlyG/c+vgqZEL6GL6FryecY1VZi0PqG33
VU2szbDMk07bMVfdHpuLBNoTK0pFQNCd4w0Ih8/1j9/dDaIRs25qvx8Ejdgp+/eI
79TCAQwS6Y3vojZWhuSNTT+iPL2jvlIrlYwfXoDQAShukN43LiJHSv54OI7jfOBy
qIqUYGscIok8n6tfzj7fpxh7mDyWlgQQ0auDF26KRnHttlvzo0LDyEbW1EtJ+rhf
cCkmcKAKEfY3qzJpphvLxWoZJ3kRlPaH0lcEEjXXqtApUEoSrOIvFyvrncYGlEwi
7qh1Lc4f1gT4h9cFMfi+b0DKhnrmNlwELs9LDOLRFUEdRlUIfyFG0om4KndRzFFy
B48kI19LkZW9cHwBmRrnrVvFBSlNeNz0FZ2w+LPk8BUbklzUgjMrg40y75/3pao7
1Eqar3UmLsdCiVGYrWadJLhqxqubkFq3U04Av6MdynYq4e5bQbalkT0rIBBAsfkr
NxV0I+kXlw7wSRKyAHtcxQPbkuo8dYRmYJfchFBlA7rRgYh0yMil5zVu2G8VKGFw
n2jaXQj1MDG8J56aQtAdT2yi7z4J6t7NYpYZaSe8tREnZR9rvgzYFxkUpXCrtul2
Y3BArqYSMMbiOj+IkGu5XToOZe4/ft3CMjyVCRTY4rkfYs8wEHviZoMevIKJ+sKb
R9TTgyg7iqkdVDvGcoueki/UyqLoezptszW38JcT+Kv0OY5HrKwlbMYy0x80gCtv
aitQnBIJp/92qXWUboWdA3aH7r01dqz7ADX8CZsTsZvRhI7ffQY7hi3jc6Zeg7Tn
/f+Qa1qLJPD1NAIlpS9pvYiazFnA/fhSRmuaIlS9H2U0Q/JccJIvpSU0BoHyv4je
s8VoOZNX19L2P6OIrODbVRQn14/Iw2aZXOm1sTxlNukZV32Pa1Ae0zw/oFsrSupj
FNsYB97y1RM1bDKbiZTNbtnn2YpFsgk0SsJMW1DafLfkKgLlGmX73qxYEw8jXGwp
OVKfRzj/RJpGpI+6UbwKDcmfnI8yMkbiZEQSpezPfnu8DzsHN0lic8ITAef8ZIg2
aFF97VQa119gRTU5eRfRGVbQ2F9joxMqT1upjrJrKMvhhGbDtshqjZt3zRT8pLOn
JoWMWsasLihyAFJ//TApVSuYNLRRwmvBGM1IxyuR/bzzDGeXGMl3cksJ8SBuRokg
Z9gF65kldlQUiO700MvWg4ISaIW3YNcJ/BU2SoFuv8/nRtoXuR2V6b1C0tidvpLD
Q0J/woN/4xZReNEju2+g6ygnXVy7hL3sZNd3xX93W5SBVdJw9uT3P5HTnrELsVjt
SQaG08Azh3kAuZNAUwkU3dcZ0t/bVsI6NHY3CPqB0ogJMsV/HndiJYf4ZemfZ+fT
zxT2IZaGjU7vqbolf+DXcKMvAPK84MlIdrez0M5KY6f7+pGWjKawPsGQtVoAiQkH
Iwxju7kF33uElHFJFq47KV7j13gg5gljLnskzXoNb9AYeMo3PYWqadG67RT1bMmJ
mylfAvkvhJlNNLBBmBMEMI4asLBr4eMzox3rjSv2O/hX+Ma9upm4NxEKttrVZlXq
8ezqPNg8tbLrVt/BF6oT8jK1UMaqYI14b/t1HWeB4rwMyCGapsYT8w4+R37LFnZw
apjIO5i6Ajg9x2OujjIDAka+rHGcfOPJYiQHMl/b0E55iZhXsA+EKZCaTR90Ik3h
pcqPdAXE2o+ryh7JBpqCkVx7ecDF9xCQPy29BzmX6XlagLH2W1x73NR/zky2tgUF
u995p28m56/mewZKsLLb/NdJN4mCc21+x3GEzygXj9Yw+s1maFUh8zzh97VhpeWI
qPoG56kjs+6pYvdhI1NkFnkVZG0UOmueYUn2BRebDaJwNa/AU8T6hYvXY5QtpDV9
HkL0/XqawH9DbFmDe6qwNEpF27Nx/DjmaHvWEGQVhzDXPQTXTZeYWABuvbAWaUzR
C35UZdwnkpoeWumAutDx85SMyVUvMTNwLaryKLyq0U5EQBnKiSwps94z/xxeSE4B
G2vNkzP8XsdHZYSQxZXu4v+QG0CFapF2MUX51kMw/uJNVZSveg+XncHwNZHW6cuc
vhjhI3Kr96VV2lQllxQLsqW59ihRqwffU9w4Cy2tM9mTji1hR3AnUVpnIHPnWFvh
4nU03YMPSJF/HoXvroW3sJ5lBeKcFWaD3BBWV9ecVjwcmHstdCSZFDRY0UF+9Lyc
Hh+Gc1WoGoGZeVD+U2RN60M8D/Nq23bhcFBp5ORrMFFkV+A5YR9dU/ygXViQ9Bvs
xnZArB2dSHIzDhZg4m+s/RrBSuuaOFMleozav+EZnyS08Fxc5eYVidEZEisndLGS
7YNur6mryUdqeXLFO30ZPkr/zPWj5WeImVWFLmL7eRJ5kPYxX0MoBoVE02Elpju/
84UggWBrEURrWfSs61GBpbtdaHzL08F9xR1owbQw77NGILwaPjRtdIKqTnTakDWw
c9anGA1PgQfiHojk5KorawBheC0amOtZhkZpuHmUh7NBqN0gVODgttZBoIQUWNp8
qk0V2h4whL1sXQZ3F+ql3YfYVAq3HiaX0NGvIYTsfs70GhS6HCL7IULbuuYajXlD
lsmyNcvg5S8V+xrnoxS0XKW0uXi7tAQYB5cm18BSkkJtawAl7cVc+xGI2kdKNgLi
X4VvUXobRlu1dbj5lwFhLbWN3SN5Jl4cM/4Hj17egtFkO2p3TcXTBtOX7TccMSlN
L0InmtlsxK1K7PQVbcAUgebEcFrC6WRKXkKGzRarx2X1tXpGsp0LC0UxSZQJfvOK
D4LY4No7WSGg4mfYEeYhxGqywPCAp03YSdw8psjbVD6RDgPyRA56FiThLQjvy4II
L8El+kMY1PYw/0RH3WeKkvoC2d58dCOakA5s9CtbuVayFdJuTRPSeOh0fz8mC/Rl
CLsTh3n9vl+PmuESnIVZiNfgCtMsSpK53kBcekf3ySJLzpP0JEBE9K2QcIXB2q30
4puX+HANUkzIzvHMtH1YnkdrekRJ3Muwp8phVKIxs+aapFeXA1+miP1QkmHGVvjT
Y5DECgCR6Kj2y2yxAovbkP9XDPOH7dBzWQNq5SEev4IgY8VXMtY7ftAZfDpAyZnX
0aGmfXesfksHZeGvOGbfodau9v6wDElbr949H66kZZgsj1Zt2RZiRqx5gcvbeKtX
1AD0pC+MlpiOTBl402I2F1AXQjs3DPovkn5omT45N1lXVmlgOstxHL/S/5prCehQ
O5qH5uSrsbLTaAaCwPBtSgoZ02Kx/eETPdoXrGWpqoU9h9N6P/GnaHh67DZPIR59
iphD0AFDiX1BzBt5jq84UfXX6JdDBDZznt5VnUlMqHCc90fKa8msmMZqku6KtBjF
pQAFf4YoxAlpA/HHW3215MifzINS4umV27+JCPa11e6MZ+ODZBFqR65lZCXbQBMP
B755T48Svd//+UPpPa3cD0bUtPw7qzT9K61v1cmig+qwebiOtw0m8S0zAZ4pZbn4
b+0Mgn98D/T+h/nUaQbnsnzE8TGv1wVWKLaqW7+8AEv9vYYMYrY7wZR1Y+52AyiJ
CRvr7vkujL3mh3QGyYeINzcE5ygFZw47jPG6Le0jENyhpUmD5wQ+wd8agB5iL8XQ
g9vNOsbPSUBFzxnZ5ad3wSOYJZZpbVfm0nZRUebhWQK/xODMOUblZfG+JF9tLMwr
+rchEGJriZ23aqg0OLhMIK73K46QAVvnmwisLVBC13tG8jKlZEOpVVM5tgo91IRb
gsQoVOp1lkk9u+d+jsy79/55zG4IjWhLzGCmjOyNN2lyCrpbBYSdMWbHdwWwVkh0
H5L3pjdkgn/9C/66q6fad6/c84ergdDlg8i5nCa5vo3rBIBZ0gmzKcv8IS0HdI6A
PJs2UdE9aPs9fGPtK6XlhyEQDWMNis4VntQpJRWtjmDUXzjjB5paBSYbWL09GrcS
XdvWQGAbjbu9NkqsUj2PfQuyJWul47WzMmGS4Lxz22Up5BcDJlASgjnqYTXyjFkv
hseCCi+vGa/F3oKdxucl8Vk7Hr2b3SaRJI6QehmwzJMVgYf/u8k9Bk2O0v+rZcPi
VNbi6panQyopseg1zWiIn8cuGm/RpWMtjZwL/NcPIKAajuZMrPeiNb4swlEuBUMP
ykdbY0qTMoQ16rOCAU1oobLwGtvx4borBp4YXB3nRxk0JktqaMxZksYaazdo8ALG
cxv1F1VgH2/FdaS+qrMEkmQd5iNqrt30KOqeOLw2J+aThceHDB1EYLGFJGNF8j/k
cNVDbyV9BymJLKBkre/lezOshmPykpdZ0xzFaglI0hRVa6sXuyR24yPTF07m9UsU
G+epC0K7WQ4psMVNuZeMS7arNi3TRI+rlC//lDzlR8HX85dScZ32b2UnU2PbnqFf
WDeJZCHcBam5r1bTeVgdJEKnutVlCgwO4bcXOA2S65VhtljxGZCXu51nWefKLw4k
ga7c0na+z6Idkl2h+v3XfziBY6q3FaVdJmRIirNE1RAT//r8fbVYK2sjtlzeIXpQ
cAUcUm3PPOSZ/Rqbw6GKFghveZgE5kXswwBGhMzI36RXAlG88etxSKLURkWWFMEI
fjRoxGM0GpNMurpDGe2Utw70ZH0zLqVGDrND65cJuFHBDE4O/T6wDQ25JVvLXUHD
vsgfIMSc+334SagM1C3bfCMmAAdA+0MMXNwQVm2eaKU4oE1rs0bG/2LXORoQ5csa
YyJogZX3tqmxKWV7pSe/820oxljkFvOLrarIkQKGLkMR8/ZDOH1s6L7PX6Rpu125
CDkKE4MJHYL8VS+UlW3UstMQEGlERlVKG1QI36NQfxsuSaTgrvUZfQr2Kml+Mjmj
d10WbAx6ww+0CsfTRxH/QFWa8fqJofRNzOIwVkE1uF5M21nibUc9Qvf1dVhEYlo1
QQh0MVWUKWIdyRULjAh5Y/cn8CwhTbLq2Ov0XPTE0PYRKeTu1WhGS7n39VNzAhVI
J12YKtm5jHq9leRpvsQXVmmnrI/w7mzRL47ygvrK8RiULnYBuQrRxnmmgXmIB8wW
5fNBuxK5TXD3WOmjFLoweg7mC0D6e4nkZ/kvwhzpWDMRyZPEXcg5yLjfoj/3Iazz
KgIH1os7hYYsiaUcW/XJyhTZPfXRQ1mQSORvMH1FfivKv+5Cn9BL67GBMdBc/phS
kyfLtj3Lofsd8mf2XojKwnSG+z242Fr30m0CVQGBt1Wyr123+0G9CQp5X6bF6QvQ
rcVrJrnViksGELI1whp6/n2Ant9mouVbU823NgpHFG/amVI9hxqlsDL+u5YEfCKu
DNxD/iOBsF7+NJU9nD0da1Li/40/mP5zBqOuG4yqp2m0XDeR/eGNFQS4ERp3+r2P
JyISCuzJOqO2S2F5PpQrWEjJHeFMdtnqXpk6wf20Y50E3O94+p8+rFAKpPBPURP0
87LCdKN8Rj/mdbJi64RDcDZwTDb54jTyCUJA/wwFffTRJmGGHz386jK66y/0wu08
H4+ywseH5EHYdsKQAzZOEIc3laOnxlVP6mnwvjIBFG/24LlvvYU9h03i1j+OCXKz
2pFkhMPUQ+7CH+oXPTzlhpLnI/ChqaOhWMkeCbnC+Lbl1SOvtW6ISO47C0ZFPTxT
0I35Qiv5vmEwNViRYwaTuCY9rN7/rogiI4y7fpM0qdLPhE9Um0LKzk4zD5or7szV
IcBX/KzWZbVY2K5ZGRbNeOl6Rsyz71lOV75wKYWNX6EDVDiGlJQ+DTnMOHBoQkDc
X9MHnKAdmGRmjUUBZZy3rqxQ/nA5MbPgOSp0DuAMnPeSnPTqswVMnlylmqvzGXtQ
llt1yIlHUQ4ntAe5mAQIywiOZ591yz7WX45UksbHTbsaBfIpmeotYNzqPY7BELlY
IekopRh1t8S4PUXYd9RfMcAubJcZz/foWyAYN+Tk+FP3voryfv8/xg5t4mmvj8Nz
V/xwLoe/r3M97RzIngQlpzWyiDGAqGzCqU8RiDk6mSyj80X4wJH4Vkk8c3PmUGvA
Fx9OgnBJre/kG6OdL6U2QbN5o1KwPJS9/WRBHbmXwiaLUAK0AK9MRvvXI8KvFmBx
+LU389a6T9dTNuK1MCPzSjsTS2Mz84mecVPhieRHXCGe58FgUaK6ym8I04GlV2xX
Wb39+AoA9b1N6rixMo5lVmkvTnoM+x4nRuhmnsrpzLXZuGTmN6XORkdrAjawG779
/mnhKd97zKm+WOHHWPFbCZkQbqqvztvpkjwBsbPApQBLrYf/u6bpe73uaPbP9sm5
qSk3jK5PPIHRhxtcfUbDTbrSbhCjMunbXnqPK9JdOJZHCRP8B/ujcDRIPQIjEc0i
Ea1FGja7pKEuQBeWG/kD89dbuNnv5o8Rut6ScE0g1WaQwgjdLdoycAne+mVvq9sQ
rD8f5UBUw0nSwn92VduxujglT6nlYd7tVqdQXSCdpuwHnmkd/nOrx2JeeYZWzX5Y
8y+Llu8nQo/nDKm4f+PpHSRsIN0x2dcgs73O1tdkfdM5ocR8O4E46bSk4faCVzjG
p6MWhnhejw0RJEw/kpu7aQI+f4LoSArgLUmDBBrgCVKaoNFnBzd2rfrkDc0Xl5pp
Zh7LPNwK6CgDVvfAawswEBWhceB3izPxAu8PPz6MvKRRn2tVQRv4Eu5mk0Od1FMO
RrbiwvGQ9IV7uvii7qjHXDbK4KTLf+RGygLnzXziRuC9h4B1aLv5o+vZz/H0GHue
2xpsXJg1dxUMUVYrkziD1t+AXeZvJ7HCXptkdmimEMO/QG2iqJwLNUexKkajKQpt
Iqa+abN+ZCPLBfKaOyFeQZrSlR/bVsv35/XItNTWsShVw3QD7cwQSX4hJRamuqav
lQZYK95E7jQ5paAlq66O/p5qNZVlD2iL4zCsjlFUXKRRR5uULnZ9bpKOE61SyZKo
ckG2qdoHAPA8MQiAlRdLk2SdgcHd8UaEOEhf5UTFgYTQUpe7FtrJsjjrlBYIQrHk
AioOOpW+xRTNn1E8kGTuQCTKW+uNz3QpziHUyesVAl9F9rfUlloTbkOJYzgt5yqM
c6XrhnGGG6ljVUDwDquz4/n2dDwUSb5ROw99tDtiCW+Koa83j9h1dg3msp+lb/x0
qE/d1acCJzbsz52ahWtIKvnLTK0LXCk+Cn0UnkFE+OgbrqqjeqTtoDmjmGZolhP0
KyPCijWxJgRJyNtCDtCibODdWYIZPqmCTbbnVAaB9mYuf0WhiQ0KjOiFdcud8Qsu
GmmdkSRVcHdnfyZmrUY3aO59Lm6jU+LF2pTFmccnxFHDUU77aocvDvsMYbAYW+dN
16PU2qg3LwKiOqhWi8SK2QHM7oL+tNKoLKwnjP9VD9XWl43GJo6cZhk36Ko55qx6
XbvijrI1ubvIEfFytt2AJgB2xdw4dtwSflgnI2Gc9AIfxp0Lq66TK0rk5XIwPOyg
HWRTDD1FoyFi4YT+jOImDTgHBC+WZtMDlIcycKdDAoLhjM240HUjEeCmAcZjsf+C
PMymck26OgSv2JHV51XZbIfTTKsNrmBPFIXtwNaEEErRhPAWZV79pICG0SGU1pyC
atxcfDHZ1ylbN0DzmsyM8TARzksaQnt9Q7FXcLtNEOMr+xy8GAVgrls1TkEBDEBV
+NQ2m4kRbeRSL0U6ZGQwLXB9I/Jt2vV9Nx1uzRPIEYc2hjH28G9WogZfPU6iaIyS
Hy+3iKbmB1HX3vM7BB00+qntzLbA7EWX6vmRzcXnpq047d+3o7Q26CLQ0oI0UAGC
zSkzXm57U/HVJm/hEH+t0v8oRAlfvEgBB/XgjYyzN9uvG3PJhPB4tV35GJJh5sIm
vKjUoqrteOblTQ5gV7lJ+PY8iicYwGZe0G3u9g/SRE1TqRIp5ZEKDJqSTDVhZSoJ
iWqrRFI3hXAVpx6ZMVRfi5lmLrTIb3gpGsGE9Xxx8bUE8brUVaJtvogkMtr8Q/Dl
XHbcGsQj7qHPuSxIX52cwv7IaEm0zH4W2rVKhYva0NeHlfsp22w6TcCG2isujxtG
1QYff+8b2/yMAL9hsbfGxEX0+ibW1H5CiJhD1sKYECzmP5tQUE3aW8yWsm5D37wg
hEFuQVvAQR/pHmIR3w9pALK3Y3LgGiZTHE1ZeJYL5IooYfw8blEc7EdrzcQ5vi37
2Nrucu9gsLy3o0laJ1z4W/GGe4wzLiNePQ34NFqcjZy03BWrwsrGrLkDkPVGdI4M
g4EhiV1MWauhxw8NlcHIRMHI53wiEN1xM6PPBlrckqa+TUSWT1QrbIXdlG5KlJBi
K1A4flJP4htQ+X08gO3h1Ev9ChQN8TURtaY3ooiphdRHOIreSGS4sPieSMqHPz4S
uGc6nsl5ZLOy/Z+a/mhL1LwBm+d+jMPfIk0SCLOOiH0vOLt6q0YKrxHFmPCtNwYD
JLMsqmk13of3Ojh7M2Qjyyo5NcAr23jpq8krSQASPQL4sODfojrFFNSS93ZxPTRW
Lt/Ng+uQP1qF0jtbi36gy/mWp3RoY4lUNSoRLJoHZrAW0JUN7gZkjtxfCR/bwAG3
g1iE98I1GqgHwaJuzjLAG0R3LlvaZB4RBtTJ7fhEOU6kj4xotH1LrSE7GXmZfYFO
u1E8PVIxdETHcaS+smdGRekQQ5+SDv8OH+HCxH/gTHuoxus/l+ztx5jWWvqktfwy
qVOtVnt5HCmHtQ+ksFG9hji0Rlv1ujXTwiZSXLrgpKAsMUW+1tmSFW29nv7+w0p4
ZFlSpPXCqz/LS5w5KiUFG15OYREIPOVdM7/gyf9bvOFKyODLPj0GJ/stv6zNGm3h
4yWr55Py0NqgPuO547GzbdPrVGg92bz0KfyQNHEOngtrte/RqJTnH4ADoryui8pN
S8+4LoeBE/XaQaOerb3cYI8MWCUMbGWJ+Bk6IoMFrLvLtlfhxxCewkvrnEtkWe6f
byh+5FHSJPFgs9ttIB90bv6TmC0QKOnmGde/sbKGfTsfQGbL6lbxafXJEyia1Gdx
+3l+q6hvLlzCbTY5ZtDMvvdi/Vv7EZWChkxLgzktoIDXzksPzE9H2r3IHaCWYDU8
1n6QMoOoyNO+2azBABfM2YTAytUBde3Z7u3yoK9Zgnl7ZEesixCh6oVifBjw2am3
Fc+0C042YFPVCak84BkCmewSFdHGVV8J9rFyTDP12A5TwaE4C2MSJSNIM3/lcuOg
3FxXQjQfPQjaevjZ4q6SuJLLuxgMVMdsqsXc8x7LiC2zz2mDxU/vxZYVql0iEPTH
ZsZdo8vanFq1xfvFoV355rTGooIUcP9dIwuyPhv+NEXPnodHIqtu6UDRblbIgRxO
993QoEPM1/yk3TgUOeCM4uk5X4qSTqMc6cYvqdhow50tvfxCSOKlID6ti+CXT6TH
RxC1sx0LzzewtoFCa2UgoDdxXwJetdPVHttl9+Sgh+mpXchzePYRAE605G11Uk+D
PTB3JskHaPQygf32nDyqgfUzyv09xwk2GEZhpFz9d0lJSJR9YsM4OprCDBCRU7VJ
Aa06SY39oAUCZ3Whh07B3kcYL/aX4KafZd04kzcGFlRztiCXfkN+DAiYynlVsONu
bFrY9LhiUTOwE0Re+gST6azHF+rhQVf0B+wmt48aqRd6VSwar3hSZA8x0wSLL4c0
+RDGevSo+JSTgtzUai2ioqnzWjcX4XEaT6j3054XvlW2yFLFT2UPEK5CtM4odtmu
u9riI6gzQr9uEApVXDrWTm6yzbGCIxocJs0UtLLObQ779NtD6ELvomaSFWK9hvaM
rPGOVEd8KW8WVbu25fS+7KLSMWLpJBqEidRIqtdcjrd6j064YLDaMY7Lnge8rgiz
5EezZqyWHQN87trDB2qHxFb8ly9TK21fGYf0SvvFsyKl7o2A9dXII/aZOCYYJVrJ
wiKEFTBjhkmwME2kZPAxjzvPSqWrPERR3hUBjFRgy2B3BFuXJt9QOXNmySkVudQv
Bo0tdogmfq/B4CRYCfN3kOhGzxMeouB6YJQJ7PDwGoIprfDOP5pDbTjZkGy/gaiZ
Fi63m4JzT1j1OfviYKqGCIzmBtXbmvo4QlsRlNS6WU7NjekyhRoIJh8HxKHyzszg
w8/hXciFblUzHuuu7LI/SArTBH43zIeYJVWWG/+62TuuFnWUJ9xk1iXM0pbEdycB
vpoSBf1viU+FJF6jH7xQBDi7JPIGdirIFncVREq3A4kV5epDUSXZ/pEQ3LY+HN7C
SvjtszZelzMyQ83HBIFiZlTQFoObyNt22HvT9Ck/BJJAxs0BhIATW8L3doWve4ZT
nnEaudbW8v+bO+juwvMeSKlUOAmIuVjpCSgxqI3xS5xVEl6gqWVlReFQmPf3klc+
Bkj8/q8rSITSkQ32MtNXq3NiKfQqiYrenw/Np+IUc2yYbXLGrM4aGCRTcn5YG6Hk
gvixBnuRVN0hedd9UrPxr1X/A4RDxikNfW8qTP0NGhcQBY2ouFXNW2rLwNq38RTQ
lEVOF16tZU1UVy3OcXBd8tw8hf3bkoherQuLIO/mK/zIq5aBOKFQGBcweipotmIV
WaGhlQtyiAhegXR33pntg+QaJ0wqrvaAtl/DeF8IFfYrEjgYiHA4O0xwN5U6aV0i
t3WdQC5xNaG7sxSWss6pLlPVpzzyItBk9Ge6x+Qkn4pGSuC986yatD8lR+f+OyBT
MlDhLeB7C/ise/LBwblHKbO4P1kmfRYNCcASOTfegJ62M7wEGzxSSO2ik86QENyd
4viEXzXnELbY5nQJy1k1UyrSMrZABCzQevHy8Rhe2UB3hGl9L3pyVxja40T4CJwx
TEjCwJRjzu2jUrOnVDbi/kE2zsxoVXI1bE2LEv/144s=
`pragma protect end_protected
