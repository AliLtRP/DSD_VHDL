// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
UHxwYbKaJ6HLDYQ+jskUzLkcmoDsSfdubIfrYSEKObsL5ndbWORlANXg/AJS6NFHpqUniUowipf0
Y5BFzPwnvDpkhJAQ+4xDvks7LGuYImybveeo9oTU4omb7ynGxCeCiiUHfay1icOtrdB3PYW0g9IU
IdKP5g1PbxcQ9Nx9zE6qNTfKZqlvimLkLlOURw6LD/tfFkgaohpnSe/YJeT28VxfZ+fAHRqIk8RA
AuSJ9sq8e/jaWEC1+A0M7DaA/A85XNLlhBFy+LGgJHrFoYldYDoGkt/2+4mgR55vz+IkLPHVdPNP
sAGyu2x72Ht7QbNbso/hidBQmOncEl75zS2ofw==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
TB8Kr0Z8kT2mu82okstt3bghRQLiBMBaypflBIc6cDAbZ5lXxryGVAO1AJStrEux/PzctudC/2uU
nRR1AIO6ICYlt0tMrqcRhwGMXBVMaINirxILCllugunE9K5hl5QpcaN2+nKjzGyDSy2O52+qOln2
khKPMym3Vd1S3iQjDw4RekVCHL7Ldm8V5961NbkZok+lJD7xfY9PPKa0EItiBvb9AjYcIcficSRX
Ust7qFWBCDFvM6snNUDoj6oOUEcg1yR6AOnRWGnP8OqzXiGkpo6eQ2+M5gI18F6S/napoF+h3YJd
zcKQkcCGypYYSuVQEvwGJOjKS0Hlz8q6afHhPdDp53XL04VHkt0Cchv/Qb5PieZr7PZxEmaPWxbE
ZOX2jKXePb9b5i+ptPuKxoYFpKdQt6ske8u6kKIsDRSPywI8M+Xh6d51ZvguqLKJHFC9ZV7rGei5
NpWlltr5zgXE866z0lgmcpmVDzosHVZJ5QpoiixNSTYoPxLgVd5Qkm0IMuyjxkDz3c7UJaK5u9xL
vtQFd3lFO/rvLjMmtiEDJ7AULLQEs3fWwHM33HiKUhRM0CM6KzNfBcAxt7AjCavrWeu1OUo/oeMN
dUY/6oKqrOGKzn0evKyhUZzVyHkKFTrbZqaayU8d00oOM0cneah0jErW4mDVAC8oE+mq+wHQBJf3
V+QwAe1RGz7PPwXVqx34+OFWIJKrzPSDvZQySQMfTRJbDjb9PnT8GRP0j9O3CI+n7u2KscGAkdMo
8i4DUvzdcrbeOivrW0tZqRKym0aGYuyxd7MoIykxyORoJKhav1xZ/X9MYMKK9RWynM9zZxQMG/fM
1zWC0H4nYzEqTf63IPsOSDMm3jp6A4MsqgeRXG4a3VrLSu4GLM59qC39Mt8DJRxWjePFASTF8xCa
+kiQefI5gUQz7L4K4AtjQpv/E9pv4YW1pHwzdhns2tA+EcIp2doShnhJcKNnFwAzWq3tCCYR/DTQ
P+jYiJ4VQYGgPDag9fieM+x6sWsmRH55rAE1slbHmcxALQA9RVbmZ2i59ZhFyk5JYEP7jg1Dwy7N
DRfpz3MHahH8/gRcjZ0zjtWaxbEmYVW0nqMz/bmdE4k3eNwzXOg2ZE3+jYnLn4HdVAB86o8i6add
nDWPiQ9mLuVRzUqYEYwez2dks8UUTRGGIA48/GvTsmQRLPtgyVMGhhD7XZhLjqBe/g6ZUCnPTaLa
nHfowdwf1TfsHfI/0JEj2X+iTS55N+WX/pBM8Jj5LKWylo272OfPuC+gmhabLpxbTOCpJ6LhchuY
IrDyybRW+izU+JrvHxbdLNmFlxG8Q3WpMuCw2tvt5GA2ezo221YJHwCZT/DshGSd9oYBthYtkrEv
n4M5kCxUNG7f1MLWYLvJZJ3Ky3semXmkiIDF+b500TqJxrHCYpuvjh/nUOYQWHhHweYEyDV85F2O
iBJxRnlV8uX4473mIFCYJsEvG3QhZF9FTFy4Mgd/7XJrpEL2z5ZI4TcetDDC4B53+iwTmkYdWkyB
j8YEwKC+kdB1U49hy1SWUSfZ9XiKwG+hTXpf1SarGPNlGe+sU/E6bEuYb+jg8vizANng46dW8j2R
8IwRG7uSeU4LkgYecWcos5sAFnbE8BPCVUb9i7z7q8WqprM6R+0n0cNf3vMTPmIg7ijbH0ZkXo6u
ibGNzVWpBHrs58cJZpQ+R1qKTN29Yn+EainUqPeH6odJV4jyzX92jUUgHNCjb0myOp4ST+o2XDwV
+/+eTN6Fpr6Xiat92BygQSVr0vI8wIqz4ePxLYArkYgoakSOjUXG4tE5V1AE1k8JzQPZqsyzHTza
ng4nCHYpLsbVzYw9ETckqBBmsoHXoK8VS4WZ/YckBmV1xDjsqzcs47X9THbxPlZn37eXJv5mg9Fb
VitNQteRKcPlh3kV6ZOrb573wKIPGqUMemrmrkcKHHG/mERyK2KrngAPJ2vU8QE797mnyaMeDbXd
KYEuZorj/veALkhvyEijt0Ur5ONijh0yzVYtoAGLhVo4OwmMrKCmARKfP8pfwW11LP1dy7jLotMp
lQdING7s7Yl5h/iw5lPDDKF8hX4ta6ob+07VB731i+Z+xPKLh0CZL6Xi1B1PygqyKolt2gBE5/l+
/Y4LqelsbSIV0tau7sI7+o8OZ+mnjGIOj5gpe9EAJoO91Swm6s8wgK3Mf0hnZznb0zSWlKKNKi3s
YLPHEHCT4fP1ZXS8JWMOWM4zqK0RFduWN5Etz0dtQUZZ6vw/Q6QdbRagmPgPobnSPDBQu9KPK/vG
L1a+JSXiUExnecPYsU0a/iM4HZlGs1OU+QCIt/BK73nN2Kd+vV/GkBOaPAUzPhSpoU9PJ7N1eWpW
jQrtRT+fcNjbRG0NP9tcpR+N9iE4A3wy6t50UmDUFrjTkNc45DVvAKn1iz8Kj+KkdglR0fL0dAo/
y/FxUeRkUTXKMTQlY9EzWXCvFGhw54Ze7bGSq7u8waxdpyAfyvnh7Ug+Y8RsjO4RXhi6XysKMGc+
f6nx6rukF3C/KFtwXWJfUxA8ZdLgzoTxTtk1N15klnQsxwoRzX8DQ+WWs8bahGuyi0uxrOoi3qUt
JJTuTjsncbNw4c96mEpWK5FglXfQFAAiuTh6zVAOmsoxHfRPJbtNpiXmAL16nRfpLrJAL9TirKjm
LcNqyNOW6O9s7VhqyTqLexpNta0k/jv7qR7dvayQXFk0C4TJ0OoXKfd0RtI+e6Y65MmzZfebX+fa
vaNzksG5V+e9bbitYjnKaRolTiTbWTyvLpTBFGbjQEDYN6ftRt1pVEJi4C0KmKXyrjm1JDRAuNNk
8Kfj2GTkStrU4AgKqV7WxoB+xVS3YeLOKdOoS3RBLSVFbUbhV2EOUK0/NPTCCHgrksmAXHvuWdPT
KQ4mF35kFd4u8tOQoc5Wg5fj7Bb2cSYg9g7E5At0BQ2aIR2A0C74IuyduCSsFbuDGpJyt3ZYqnBg
7tBuInloOOa5SfXIaV7vDjKA5oPAlifA5T/ZMPrtXgyK/2t+MbUGHOClaYnF/Yww/vZoHDwaiLpw
CL/jEls2yJkyhJNTv2wElXLuPLd8brI06uot7PUa8q60QvJPpyUjS6rt0Ob/2XcvRc7RDCPHbNSB
7rxKa/UylJc4jQuQcmQA+GGAaiMS+3CWCSSiuLs2Kq41kiCFS5Xjr+1zzdvYit4u3WuFoFgkvGX5
x/TEvGVACD+fcSg25nk27J3YR/3qXRDM0/DcG5NIuhVbbzLDcowwDclmx7oQVORY3i+D4gejLU1y
hsR8nezCdNMi4/ewMOmSVbYZwyYgFW5pVefFV7h6iEfBBMd/vBIrncAAMSZvUPJWuVj0Dbxm5iyQ
niIX/5WyR1nrNnA+ACVtMZT/49uMRw+f9FSxwLJGuwfNsYU6EMVy7t2FuNmVq1akvUHsLQPTrZ90
eYxV+Lul8BmS6GJyhM8RTKwZ5618TmynhfUGZ6ZAP35LacUM97gOFlk5Srq8xqSagzmhWUgWGIj+
g1EPP/DmzBYiCKkV/a94bwdJpwhDn7uPI3/dqyJ3zETy6Px2m+G42fCYDniqpUXqg1F4oCggLiMj
UeOhuUAADY1zV0f+cR7AsufgsZE2KTIyaf3vh8u+RyFU42iLs+c40FbHin4m3iM7rZ1NJl0nE3qk
D1wMGuX9lKuk14gaRvBE/g+nt45Uf10cC+Z39TCu723OSaj1LZKQQyOxzUV4cgmNGsHJ8xRH7pGA
Cr+4kmmn8e7sASiD5fx0fNjxvuBi4ZMkwfvqS+W8YBO8k9lzLexp8PE2OTuLHHMfIQtyrDxWpiSk
DkFqPw8OJZ8tHiLBTJ9P1r9TTsNBrc7lftq/rU94/1SS/zP9cyX9GR4EYlXSmfxa3oo2/zUa5DOl
+xcc3aQDGSvwoy9w8wu049YotlKzF4NUgGYzu9oeK91jQaSiC6948gFXxMbY82t4H4iEapxKv85t
IsK12HyCi+mn3DQXq66JXGgCxd2skOEJVPxiQYS3snrms0uvZTiZdrE46OjqEXUYVoTp2B/MCZEI
hzn5+jQq2SPMms2cj8MnQ6s7pmMplGmMeioRIy86aeAlKT68SSnWpZkwvCS7hxLszLw0ovfZzv9m
lwcO7JEonngHG79QNFCqiplUNObX6kYwWqssrTacU/Bw9XbM/O8f4ZMOFGkv4krqPiMVypJ8VrR8
KM8c9jn+AjZfGffTdq+X6ALz6JkL5lwvGieOvGEnzV8vONEvapon/hJcB7EFogMY8C13+IV7x/Wi
mb2CwjcmeGq9qo5JvxLwfRXu+6KSPZAhGERAyWZTujuElJVOmTilBWtrmSplvZvGapVAZ44RDwQk
tsnN3eXnJ1dtYNg4tF2XXIXxmKJTyDlUEeC4cseLSjkak0rYUcGKY0H1v7oJ6ayAxO3ReiSXmfHF
eaoQCIHk7OEfvBslRVSAUQhnTXdMztf3YWkOETNPyHehzK0tz3E4CMEbq+ne4GSXDg63HDNlfFYj
62Wlz0D0XtAtFlqUUOyMr2sHZjgodxdQ/TIt5mNHg4EdKvUuJhdl9zMO0XiiXkfhrCbNgwKQYZct
BF6rKMIGhlousJBpwLSj4lC52zsqPKVAeLNYmPr71ETJ0M1aTFx6Rzu2Z+e5MDqjUkxiDAZP8QBy
RN5MFyfak8m/gvFHS/zQg8qOKaRaokLD3IA22E29H04/kPa8sulsf5TgjxdFcqLgjHf+/hHfpho+
p9yK7Z30wcHiGXNmNMpPlA8gfhtrPk7Zge5J77IZH+dTLhls6zMKPDOEPDwv76O77UhZsu+0SXkd
18LQOWfuO0KR17GepUc/s6H0udnbhauLBffGx+ScvVFFLBjG7w0JhvqATgNLDzrVlP1lXg10ohne
em4Ea8PDFJm6AgfqDWBR1YJ4RuRD+4JcbRfMUVwFiMLcon/kwTLv/t/tWyxxPxOOjetWL6L5mTMd
VHnsPULp9NzArdaX8/lgwGX3pET9q/GADq04lXf3S4LsqBGt1+Ncz3aa2dCCRTdunpDPgQgnF95V
I6iz/J0hQTQBZfXShbiZp7pYKJe/S2Y7D1jntYugk6O/5oLEuiJ1cHG49fGe9OJXruSZiLNZDzX7
IEmTJ7MEUd6ssBvLTaHB4SDkoe1gztgCZ1WzXyoPeCnGcNJhcYxdHpGQEKRc9UQ0DstJ68lBC+Cv
Lh2rguK/LfuvioZ+TFZd/3W0lKmq/qtvxDI7D//Rs0+jz87QhzKGtmXidqLFHsJs3cKG98so61Tw
QX16eSeAXZILWa2Bx5Q9N8Zu+0nzJ0aJ/uUc+xD9HzHlekHxmcdkmCGfJscpJCZ/z5B663e4/xsn
5HZB4ujPAEdTsG9gTiXa54bhlVoKQ/dv7Eh9X1WCucGipdm6DS3SngHN15e4dvyqMxXEQmO9IT/o
/gvG9TgTKtcd5ulIMm/ZDsUG+0SYNXurxgn2uQPPOK7AN7ricxerZ3nANYxh2Ayq8c4qo5qxXtPQ
h00IEiRN2J4fHHq5NynrINKWCO41xav7G5MUYtl6OGBaeh5XIM6fpq3URls/TQCw9Et+Hb8qgu3k
TWt8/aSv+SKAzGXySKtABtaTCgB8hxSRR58DhKdxD49Igc6eucQOVvtC/ROYPbprSzlM16jUwnPm
8BzRzbjtXdTwg+a3DGUNzU1blIS7CNjgvD0/0+Gyru4E+LVvpVJWM4aGBhrAfi4krIZWRNQYvi3p
IWIGm0+ccuco63xqvMP1+MNmBRv2OK3oVbljdMjleuw3H6SJdq3AkPURfhvjE/YAWRhhmdhZXjZq
3gaooIMZ2qThL/utbAzpmfwTjZsNmlCA7V1ipq737aJsn0VbhiBi8mWvzFfwC65sYiwTVxJuqIMd
YyH17zH9q9CND6hdFArwrt6BS6ImJjVH27SO1BPh+MTLdbFiHm26EtfgGKKrfKowh94DsxSQxIKb
1dVx/VSeBKz5vXu4hcm2CUTZDUVKJmm9jtdNiA2rve5nJgccaGYescnzm9ESkxmyieijg5bvoGuw
TzNS6IgKTZniD5p6ifEDlC5WMVWoE/14mCpbvUNKekW1jx1ChvE8TOk0cyd3ZBIw+jonG19fny73
qN2q+mM5r972QuiwES97hjepYhVOBoKYZBc2D2SP4HqSp5CehvVEpNYtGIMERk6uET/8ZS0nnGAV
bhiqGvMV+7CSteLXabGfknTK1l86WRI9VBd0/RLxFRPkR4GoggnA7IDK1PYwS4cz6toNxmMv4Y5H
yezqaAfBF3QnkQ1b/Ejw5mHgCpRay2hr8XpY/4bZCEC2Az+gISrdMCCdUUfZNj4nkGakJdGCdTBI
F5lv4f4Vd9mwx1t5d+/p+Le9V35HNHHDkSjAW0BF/f07Eusu+kCovUE8oYzjc7uXg6ICmb1fh6Ad
kljLF0rJsXWmEPYzrD1UL/4J7Vhb/XVfC5VCBmVrQDpW4bsRor+3oUx+lcOlW49UoE2+0YbU+JYI
1ARt0oJTC9GXLbABYWOGVW4yzZBqg7UkgMRnicuHexCkHydIxtPvudFPvf7jx/xbz5oQZnnpoNVv
0kWh1MAPUskoct8gkxNb2oDrx9P8pWiZvKg/M5LovYxxYBkA3KH1T6A/KGQEmc+fSfKWnuZnynDI
ykh7Cd0jp4rVGhcnuIKVQw93eMHfLhZMA6prznYxtouoAce3T75iM605oqQsvitnIQyTmt5O+U75
pMiARAHuhTxRCmHbvjVFwLK11cH3SgHi8k2xRnfd+OuIdPqdpcN9ICEGXf+uQiFmOSs+3UX1vPcE
fQAOvsHRgBn8OJilsZA8xOgzA5rsowti+/xZZlMhOAN0cxGj/UFqLmJ63mHvyBgqNhyFMbfVNch6
Lk0xyc+YFKQXIpo87OdOuwk712RFAPJf+1eRvfAYM/JwVEd1da5wpv6gP+0/JlTvE5X6qvwmjA5V
zB6+P3cIHxoo2X+qbXVQ6AC/t66kXL/3GmOBB/+JoPaBabZSSI+cEODIhJczvRNohxoff9CfXHJG
PPuY4CWOM/+k0ZZJKanR051O/rac4AfqqS5D5q9xlVgKRVcmF2/yHF7Qx349jVOrF75wGBo9bL7x
L3BFAndtwpV0tPI5QZghZZ9gvA5U+2HJVpRVJjkAVmGQjL9d/GVBAGeBvL3a2rTysiKYxSE0u4e4
Xw9JkgSoPTFQH0Ddju7GY54HsB/ooTWMIVmsuetQhvglVDfAYmqi9px7mn03uQxdeZuglYOoidyU
vw0ACOY44F5cU3G7mv0nnKovHQc4KIYXXkCWobjm6avUtKjDdPNxhWEzW78mdU4OdiiyAUVvXqs9
KLtFQ2Lfzkj3vZnqpcfPlbpCoAr457qfK5LU8TMoxAJy8yGTlY2mAhw/vSYNzRRpeIHped1cuRiY
Y09TqpjjaF7zMK4qOczrCEinsXK9oGT9nvhHOVHxA+UAMC7vZfGwaQFIUN5eXd3voNNANAPr6tb5
u9n9K2rqUDUsJ7hHca2DWPoxSg1jXUb2+cZozV3fn3I0eobeKq619FsJinwrQ9gKgnxEeBK5KOyt
C3jmaUW/BefiU/sWEBz8VR7RUBQNRnTcegmilBR8kdYos7UoUuW/LRssZ10rI+SgI+t0bEUskH57
OI4jyRatfRVrkLSrLt2IiBko4Awh6Q9yCUFb4aDmcnNrvEo63A9umoyjQFTfubyIFnM8tsJhoUui
vkkGmTuVzyVDUGeJZmvxi2VPZqrEEiEjq36ZwWyfkwPIA+q4dPOP38DTt1nUEwzgFkT0SY/CntNg
HC8iQ8ST0yTN+iHHHmCowP2iDk4B7jehF/cHfXD1q63dJQl+dDInbSsXfQOKC9/5a5ucxbOKMQNq
jfjIGC6Z+TWpNMK5pfpsPEM8tYtUM4IgHQMnDpoCDt1WGP0qywUSIYSzwBaw4156OQQvl2yxvcc8
EbhefFOSMdoBrxELcMzFNrd71J5HqVUnGFur+zsX9XMRv5XGxaXUEolaTu5uQKUFvJe6mK3miYWc
dxfcfV0JluwOqdOnTInKzCtsDRj4gjRp+RcNVbm1oo3A8TazvwMunE6bO7WXX7RiyoY+uVDKm06v
6O/wH1ZKxUwPErvn2R8EfF7Ht43pBIfPDdZe/1KU8o4D0seXVvcbF8HkbaVerFqgN///7USzdlsr
P5HLQgZcHL6GGfn4rWfTNFNJ6dfmDZOf8UY/BkCt/tc6P1mInFwhFKywZd1McOEjO3V2AMa4iux6
a5QDUZjfFw0IxZzwmR7/NAvMpuOf1lNi3Xjn1Hzg/MOok3pmlmnpA8FSriclE3/j4EYQZMuWpEDy
IrrW5yiA4rB3fnfkNc0ipb3KnpOC+ZQ3BiDLDrQpHOvJvEjTp4gvIUrkj/COSg031ARb3KpKUOF0
y1eq5hSKI4hrY1UJFwV9GT0M79NM9jIToI1cOvsUeoLT9KWQ9vWg5wB3x1Qr/74FZbeBcdCQMUb3
FFkNJGAMSDzYBwV15a8Pw7ZI8GvRPyqowirUG4mh9sCqxWZbZdBeQlq+c4c/3TrBBTitFQ5RwaHX
cieXianWAJzxQk3DCpKiAdIjZbadrSh1sSTKqV3CkkaosRCRizss4Lrno9c3rqSmy9KxOY7luSIA
XzRj6ieU57hV3kUYxtdtCsasfyRShguonU6nY9BowtoBWVQg8GfCB2zMnGwYa8xQ0e652mk9URCX
Oz82PMZx2ArbOv/RbQaiRQc03dhFuBDfWJ8S3Ns4DdlWQbSVCU7n4TRPaEfQx+rh3H6eO/vBZpQk
oLUwx3nhzBvGlaJOifCUSqaIDL399SEvuaBT+xknMrFiFcz6DR/HwpaRpB1vSZzP55ZzMzhdIr4X
HFOREgXFiGyYtzliZL4j3CqFSIf1X3QO5cbPhGnY01AodOYRNP80rBDgh7orNL3jgmzjCMILiPWD
ZOlwQ1Yzkik3L1X2HacFtQP7HIcpHNSUb4UPHoiIQQfoUOIgEY9zIbjvTiH1sMcsh9+YNPmqVcXP
RKyqz4/vGTixYJTmn/N6wx3iOir/8rskve4MptQZeSBuXfDUKfxbhu2ot35So7xO/+8xMo7nbbZ2
MeyyqOgPt+tDjKxILPpP4Dw0yhNGEnZY6G1DsGi3jzP2RmY2j/ef+AWunAx/zl8DqlYEkt2FiX47
TO0FjTPYvPpfEwryM0eDQKX+EEoAKTrEooKLw1FRqZNSotlRoJiIddFsqmi02EoTz3FVwO/+yqvM
V5ZAIyFNdOnZK8revpf/51fmv0kBDN30M+0Zj4hOF/tkOosXWz6qXKzhy7DN1XgwWOhpNGrZ0phR
Q9ZJ8y2Fyns9L0pMm8baotP1gL0GfHOQu7LAiraSRhE09oINtLhDZ87XoN6J1s7Z13c1L6X4GvNy
hguTgQWQOuYidUTGOVEc+mEvWGzYYTrAc6kggkYDKn85uH72I+1pskfKuB1dGoeXALp+6dp7qQ9x
MDwYM8i/nNdpCcXoxFJAD0Av6OWxIY2mNRcR8IZJRCieLCYj6PvYYeXAfHY8EEq5EFJX0zIEZByy
yn6oJdThdGcEBfKHXtEwAGJ+ZJvEKr51WhSNiNhSePShDEBmso+MtymO9/YB7aj/AWguE+JwE26R
ny+H/B2cm6Z1pLET4f9nbajRpghvDSxZdNIRODup0sAH9WW/rqlTfUdL+yPy1o4VmNm9crRpvWL7
MFpSLnl1fnXSRqaLMeEJtcolWmbppTy3AVrk2HXSDXl88IaNyMWWr3+R8camGYwitXkYy+EE4t4W
182Qnx/fMeX8rGT5MZlqTeP10oV4pyoLp1qqqboHLBq6uRH6+zf7DHtoNdwZJK9Ez2Rrf0VybQ2+
/f0E3Qbg/cziH7W97pzrhB2qjgiG9nu8OQs/kOnbQ26JhzIaVO8GVzVptwgx/gYsAs+S+p7wc39/
+495aXvqDItE3zM3qexYpoyBRJL48qUeD/jtONBUDMs1ea2E4hoT62t9pUsEzt0CorDeoIclavC0
ky7e9onpCt4rNc5SfjVGrVS75BlapPNAgbubGnpqm3JJDdm4wCesA6ACaQZvufTutuEsY23xn/4F
lWAoL6TVB2pVk0dGu+QLrL1muuUfz0Qe4SmFh5OtHAUAbuNv2pzQ/OFLVLpry6jf0gHa5j+JvcT7
BYgtKnPDyc+gdXeSw4BzS6iXjlQhWWzOINry20nxHsStGF8WafX462YNh24DmSXCvlH23vDXEXkN
G7DQeonjjizC2NUFWnGwGAtOZLvKeqC7sNWrXG2O5xLcO03T+DtDNk48tfz2XYiNi2VOPMicdMLN
HEmnBkhl/9p8orDtJW+dIbfWnoD3l+wD0u+Cn+b3ARAh8Yofs99fqv73++k0e4HdYhKrsM052of2
ykDqb1uTexgtlgX/xa1y+HYBbi9s2/7dkUF6rGKerPVmVArdH2GHosoJ3lwG+vdeUQRCVTOX2KS+
dk+0vZodxDDBJySPlGFeDOj0xaDk8FEq49RozLU3ItdYhnrn7Z7IDhBJjDIDYWQO51jXAUWhehCc
PD+8wpddc0aqLgLdZJHO12iXdSYkEcV+xqIKHJJlgOA6W5Yj/WJX9pW499VONnDZ1hLPIcHIjiIK
xevw9j4ZhakxluCoTESsgyPqrM6dd6oUa4yjs1D0bVqcZ1hTL52OGD+K2pzBckbyaZYZGT3+WSIg
fV4ME021IFdkamvzJAXY2mynKy4mFPupxtPLJmpQxbGrymbC+m2wGrHJyCNCSAe9NE8iKfhm7NjE
9EKHUO4YEeRxsLVl/JgbLNjVuZXfbxYDE/zjq40XAiZ3vQxS1EWlBM656c8YS1S70YcFEh4sFbci
Xl/z4914Q+frfemji48hvrGJha0qWZLas5CQ5khLSegN71wzneHTwbZOV1an0IDm4RYFMWR2SnOA
tkS4xLLh8LGhyXIeWnE0GbpllzerEcoe3ifP3ALGS7vqEefdjP1oQ/Ang2jQTHUS7EhaAjhHDKfk
f7wp96umsWPWt8PZpjegmNWUa063XmHr+7fXG4mbWJmoPZMdqcomKSxEH9DLB+hwwMmbkDlJcYex
holo8smufOHQdBtEEVb9VjteyqL5K28vTJJEzBc3PKVGekS5yqdWAEQW3ISC9rsVMTIGmxH0/RGR
eKbNEoMszlIg7r3R5ag=
`pragma protect end_protected
