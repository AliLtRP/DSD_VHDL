library verilog;
use verilog.vl_types.all;
entity four_vlg_vec_tst is
end four_vlg_vec_tst;
