// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:35:44 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
rB8+5ZaKSsYORJz7RJEp6KF2dKVrQ8gG3w77qZRiK1GOaTPrFkm2amobluLFM0w4
D+FlevFYYjJFJiBuCgFqvlAHRVr7gdC7qusw4D6LtqUrlTkSAay4rF7D/eKBZs4L
NDRd1pNiBzKmdgR2+SsoqGNy9OxEPm36yNgNkthzRqw=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 13680)
RhDUmUAeCDsal+zczhG5CyPRtdFHrEJkqWqgRBAJIqg5YAMSrTCRh5UEz/2PJLDc
77vH9MH3XXhFV5uCfBZHBVnIMx/h0+/t7fFKB+/Tr7ZitqthMXzJJLYQHdXfx18O
J/jLua4/BL1Nwo+fBlAuBpm/jqyRY2FD9oDEaBCXTXrYxQTvOq7IaMtfwQQxK2TH
jf1kjW9+xxur1TeGPBVkOIrWfw7ref6nVTEPV6YBnUqr7SBX02IBUZrYccJ53BMj
RLYubnjuRZYCtjAlkU2NgqAi1VHISUaB4v9q6ZeSKeUkefQAFjx2Hz1aDjJoRU8l
Tnu04jv4Vc10fp6N1aMNfdXc66xLE/MqSRYdTk68C3U58Qgd6kE48vp05Zf9T+C3
snDEuvxt3qzG9jQventXfepiQBSw5lCzltWqraq4a8nXIPtyZXidwTiHwSSDWy9n
ncb8lXdfGf1ZvHtvmdkMNaR94DqM0ISm2MrdAKTv5GUXHbFiwHu7vY4gBALBpRN9
y5goEp/He3KXO3E7hzhlx48vgh49j3qokxw1l1aj6J253DQLfCx3LAYrB/AoEJsr
NEbecaG92hcnzlAQNJOEa7Q/fV8rUWT4XYSLCif60/aGSeLogqFU14dYPTE5eH4K
Q8XqbUsB6MCRrD5kCgjF697HZqAOa3F2ZsOAxvAdNuKobKD23PSeeNpSKTdEaDI0
WNEk5/Z2nWK4Qvd0gWJtABsXWkeqL675T77ZYzz5k+fspPbVpM19Bn3U43u+ncJs
WO8SvJbckLY7X6rTmqA0no8UvOPefDuOyQRQ7IabIYeB+trIUWV53iUM9mmxpNeI
5jsCDoMfyPfTCONUcTm0lgsP5OjEiIfnnd1urxVva2vU6OUzFViZ3xuZuGuBY0Pr
FEXTPkL84zbplNjzg9iI/4bXQcban0u2bYlWQmUN6R6cGo61y1G65/rVcmhULbU2
tdWK5gS41/P2WxhcqLeNDgZStzmiVDg8Tlx8uElx2xLIwqXm/kfB4gIxWZRVAKnf
X1HOoLDTxJu3UqjvGmDHlh0tJTYxOXeqWRCQ86Yc6xa6+s3lSQbXLhv0yQzOD5Ha
rugSWt6pEVHTd93z2vh91PJSrB8c1PaXUtkDso96o000eDrmwB4MMNaiRCnP0BKF
Z0/yzIyE9equYvCnfG1fxW//5sWYijSMhXgbC5MbVVIXsvWqTNRIP2EoSkHzHIcr
R5WnmO4a0BA4Pm+Epk0nrMHmTGSn7tRRygWCDhsPYfViLFkgo9kKXlaLvZBj1ZDq
4evA6rFmhUJMV13puXIIUfTh5MWa3Ba7Eb4ZDp7dAhNSyMGVkRBUk641ZApaP/UW
KZu2rcU1IjDUoqNaQndST+xO5VNEyzrer6Nn7CpfcyBPld3nu6POQ4jq55fFRhH6
8rEgOQbA5fXBpxe1bRNAtHPfvZVFjNqMLVr+f9CAoKtkGwbYl7V5SaUCPQeWWe4D
OYuguPSF0hTgyic/eS5WnEN3n2D9Wi5x35ly50Pd0bwShztFyMfmf2aebNhoOhOW
u3Yx48df1ZaLw8IsJVZOz+3rZrljIzAlP3XgYIDIVQzWlPjOhkZzxJRN4Jfa2MgJ
qrMYAzT3MV9rNTp6D0RZUx3VVA6kr/yMW2Jzx1hw++phCs5aX5/hPdba8XvdxfKR
s2ALRDxhqyaKtPi6EEgIHYlIyw52H0PL1703xCm49qb+qEJBGQIye+6o8THtGVyF
aPHDPyyZFW8sbtJrbjFrz51CvQnMX9+FHmtKmOwRvx8y7/NzRm5aU9dpAIRMKooj
/5CrQSa7Jh79Hipi2FHJaZ9+Z1IVEd2Iszt+fy9qzgZPzg0TXXGAGHkagdtfFHAh
O8GbCkMlsImq35ZPe8I4OWuNN5h8OjA8SAZLfUupyjJ1BNBFN/ynx04cpNSAXRRk
VgRP62DwZUfn2ZpU9VxNf6jo/z9YnZm3F1GyFAiIQRvqweJWgcmA5t05RlrubehV
kxpHYIg5XA6T6FN+ojX8mW75U7/q22QyaSaAZu4ke+QRXeXvmxa1Ecp+6gpAJYG0
sG9ew7mHvRep3ldaARfpM+wdh1tS2K0UF23cNl9l8PCPCeQ73Jkz+Qc1ilvHc4u/
QS6StnPbq5qKNqoC0PxGruZD5ll8mBc5j7l2Pn9V6RmQ6J6UjrOqojUvPhWGsh4U
veRF57MpQo/KGGBSOrjWe7CFGpEPv66Rw1LYX22e0DFKh8KOdrRylUGCmozf8HDF
uN8lV9YsIj54jZutRDykb0cNDFyQ3VZgNqdegHQ3zXzOwnszQBN/n8klSLDgtR71
plhtvVYFHic7FU1R3a3vneUrAcHN/de/w7UyVUHQeMxaShGWsR9LExq6mCcIODIS
qTRqIr4MuQ1lFLigBTouCFC3OnzR3CW1VMsEqlI/GeEaElGdKaGCqD5/COwStszE
89B2I1vRHs+EauQyLsDUsDCgXunMkX6c4e9D2vFjmpgqqngPua/Ev+NcqmOJkogd
kux6MrJke2EhH3hwqhza7Cn1COInfCO6s2OiLZKOoxY0xjre5ZKZQQquPmIpihbx
rTNiqy6cXYjd2PNUwnA3o2kxO8diHcxrV/BBqrI5oaduxkag82X8j8Y+Fwucs/JK
NZtxqWR7D+BMVK3+qdmPQtQj2WGMDdEUOWsgOCfIIaJUTDhSpwD+t62VtCUPALQ7
T6JmWuNT4hFYAn5/9EblflWDtGHQgclA8DjQAFdedyBNAhoxW3cT/nXdYex6v69t
Zqtg0gN90VU1vMAyhodxAm+d8aIV7EwJQTQLwLprqBhqQj8yDr2GmafBIWEjfh9X
vm1l8+p2C9z8BOoaIxylhRfM+F3xpamDYotnOaVlFYD/BujOizJ9wQ859C+bJgDL
h3/ioXw4TYTBFkNH6xoDKycz7JntlYIR2RRATdSZYINKkctYzbOjDOpL09/W1N7a
w2YX44NZ/7faXqPaevO5ZV3JloePdoC9vK3tJ+xT+sMZNb1Ff4k1+8EnqvwJxodR
9v8Ukz6NkSQWXobRZOCfsWngjlsWBwhizLtKC6ZR+AHAAPU0H+9+yjaqB5PN4Xkn
O913oH0XUYGSX2QHc2X0geyAt9j3N8pGsWBqbb8F0+KbwoHCRSo0X5Vh3HSyUn1m
zMwlWYLvg99UVom6ovelq0P41GxDdrPCUiySvkRRbX0ENDY+3XRUl/886mv8thPo
Vobde2xM3uO7YgamP1zGnSs398gV9LE8KwiOoJ1Iz9535pHRa8L4dvN0fxBxDLJW
cZG6hLYjE9eoMYmlwWBqZkTzy4fSONbU1fkJLM2DayyxebEW6yeS1swDNbJyUntL
KvrrIMh8Lnn//pylW4qMBwZ/eb1knkERhQ+FtrBb/YsdGoVOkD7WUqN/5TSe1J+Z
gy4iSUSnV5psjwLsphtg9U0TEyDeGLxLsBHZV6SgU8+4bitRs8gbodTEMMKQTVzl
7nflePqiHsfQYaV5GW5x1W02+OCQNhaFpMy4Cqo0oT9TJo0FAZP16PJr9W8O/azF
bDN6VBzV85WExV5b1JWaSIWb0qbQEjmkcMR3om+b/DZ7u9E4O2RdFry+Agi71i0x
+Qocfd7Kv5LTVZdmJIBx+TYFHpTdwbkDMw/94IzKaJlY/KZsQtAXSWtW9mcqh+2E
GGqTIBEjGDdAw/MqhNzB3q8CloxE//RndNc6sTQXltkzpqZ4rKgPXOXFtBhevx70
PVPi1us9MgFy2X0LWn6dyr3HKEXuFxA32CjvabUNVmdoVJ4xlgQyCFKJ6KvwVp/H
oY4WNtBgS8RGpXM0BqLumncoJjQFrCPMtzGg/CWDtQvatlTVcx8svCQaY/pK4hzm
s92tP2Py5JRFrTaelIlGJIZEv5oS/RAB3RWcNgHpS5ESJGTgBRvCgUptxrOdaANt
q1JPyGoJ3Q+Y3GHJP4I4ibDg/NUJ5nOuIZ1mtxYG/ynR1tKZydjge8XgYBXKTBGm
bI3DRDT097kaMM+wMftGVR2fYJe608y7GDQASlOXVYNO7Srycv2Evh0JCqCZsOPF
xko4tdmTDHLOpMHwBXLSoAUnC2hpxs2DZIcEte0qym4C62RYAgTErqt7SBt30wlA
ZJYc22Wpz7suPMIeP7HvuJ9/gmESLsOvfzGkqwumfJudYedJMWnEzanMwPfDaTmF
EQzfsh3HlSl2PtyxIZF/1LiTmNFuJ5TuIy/bniFw0s8LLGxA79ZLWekouDiC4Tme
7PxCwmw7B4Jt3k/uzgAAcnWceDtKWd1MS5b0eqyQ7pGqliFiBDFJ4pwyxMXcaM5y
F407vBZ+GqO+u2QiAWJ4KdAIx48K+TWZ2HCA6ApnZdJoJwF0EMz4yzFX72aG2fb+
nBcjohzccNoWezNUPAD/GckMWdCzwt2DwdhaX0XOGudmd1Wukg0ecN3refhAAQ4g
cg+0ROH0F384zP9oHtVM3+8xs2/Vep2dNhHNFuJmlOuvGjcfsrLQzgThpg36z6xp
V6fdwRi65dgpGKrD3/NTohd/vpuIw3Usf2gFzsBa/TGICAnRlJRhroFrUKEHhVSx
dJx2MACPxUnJ8NKf6idYU8t0w7D+U0DuGdZLdFnUSaqoHrqnVgc1IOsYt52J/Vx1
JgQJ7g7tC1OmgAzii5+cKa7QNhVcip6fVlFV+6Min1SibLXnnpHDAhU7/tDgcp7d
wlNSiQ0fgHgd9pFZOgYBeZOLKOz79zQCE/jYFZaxQ5GxVZjf/ysDHim9FrwXARGp
lqWs+Wta76OhXq0TAB4ekaYoieKy8ilKO9600qcxDYYURmS4hVaBjhPE2cwFyOv0
dhY2eVhbCNu+p+WhJskDQr2DP6CPwheHTwDWY/31psLkthCUKWAWHMramlQlGFMm
BO37o2k2Fu/uYC/1MEAJ2zbdDpKul2X4YkSfL3FGdVIXk6lHHOdnCXeL+NFg2BoR
gUwt7lyrng1DjOaWR3pYU3CIwFuB6DPq4KuQ1ReJgayMaBKbbhuyDb7cUo+wi9sA
oa7TeK1ctRLo8msCN4sh9yO3MBOLxCYldzI1WVDmsWfAmdiWClVTRiF7z4WYn8sd
VzrG4H/dIUraZ7EJGPFXQ6Sdkd9xoBf2JzxDq/EfBM+qMEPh45fPKnKf+YbIIqZn
yKG/6k95Ymqr0bqNOqPcPXoEuX3Y+GVPZWOQoMKvkm1SdThBDHoFchnMJPiUZNcZ
eHJUxO2plN2vj9KcIbmuoDbTs7y6s9IRmyIJBkPa0q5B2kFTkFI/WeJy7dxzajeT
7PZU2u+d/tC65lSHtDWrplcSq4wpjHf850qxCReCsNCh4xCPl9+iO4jWPP2tFDyt
JPTL2h+GWBVq+7M1pbl4cOQMF31CLjXUryU82soqwnr0q7xaK86emADJetx4UCvG
x4fDcEAQN0xHuICrxUOUSrOBdzVSlovLqVG+msBmLu9AwwiFxgCumZziOdP0y65+
cx4XvtMattl0UyWPdv+pMje+dlAdWZfLXuiXXol+V1VCUQoz89FbyompdqauTMvp
sMAeKdrs10rnHmAWtl8cG/qR5foSV0f8VEoXuegV88EOmeY/qDTzpv1Qur93J+eF
bUmt0JaMUe5BhQpfA7msWe3/8VO9Fi9e47DeeR6LiIa/WFEEKsO62mxDt3Km/ktr
zOsoWko/PBnospJjx/uK/3VwJmwBNgowKdsfogJ887/pt096j4dphVp2aXtai+4W
kSdWvHhLIHbqxbdcHjbhAQZ972DOgXUM5lV/WzX113hjdfzdrUay7j0+ssYYqkSj
/qVy0ACspXfsOkukoYn7Hml6AL2GmpUlMUzfhWjSfuzJPlMSN2oqZxKWppgVJIaM
g2C0Yv34yj5/RXRzC2CyAicee2jOzg5ewyRTwLPypVb46o6DX4HK9LFVAxoQXY6b
sPavtS/FGh5nLefmwYmnjl2bXhjIoaB2v55yvOyLQkx0F7h12XdpeBdU/IOCvZpW
FafqlTbf3bjtoHFHizBMspkBOGgIBDm0rm1bw3H41CNq1frwwxxKPI6Dp+o0clVc
RaPoRk5KRp+Ge8QMBtREjicMHZy4o8Ey8Okyt3pF9jR2D+WgQmqyyKXo9wLee/I8
cgMLBM4iWaKMeUeStJSfoBO5H761w06PTj+Y9ZOovT0EmMNqeXXU4nHDzSjYjfxx
iaj3WY3+58BlDM7iRKYaCtZEuNMY/PwL/CJXOIt1chM8W1VmPCfS4952vzdujw1k
7gCnvQYadKe9+JjN1y6cw5nkV6GRKBk3E6bhk6aRRGh1ntAJ+WRVU+MWSSsAxFQS
NT4DmENovHk+D16ImLmLlgLtHI8YK+H1/3SjbOJB0w163W5YBeSdsPnvu/UrsKGC
lyJH838fpUOeNqu4FYBlvj42phHkyJ80cTu/P9h6IwXMK5cxYQBxu2R++f9UgOH2
vUUv817tYBFhpDJOsoyl0cC28zS9oUvpu6Z7SECTwebggVtAw98ZZWBxsPdJD9s4
9Cr7Q1AA5IXUpRdLf4yTMjeChYQ5bp1VtEuv7mGHn3nWpmcrTAwecT7BYk8hjHup
TO1HuOIrwkUHVahgcTdj/ZflhpbfxoZcNUtPYaB0Una3F2n76kp2jCK2Ujn4w7lR
SCW4cj1RTyN2Glst/UWtZKaYgkmsSFWl3i/9lbYn8ThU5DpyhqCJfGBx9ujoJfGe
mnLZ4MtF7MendywxVxPTE6sf88BHfhTtxzq+Pif2TlpgwhYrdQVkhaAaRNk0o6Pb
7lh//hF/JwCTTZw3Rl85kDupU9rvdTKx/1c4SwmqRydU+PWoulnwB8uib+5YMu04
V8d77WvMh9hm+Leois5hoSr4xQGXpxuwsMGrI5kfAknNdIFY9Xs3KjE4lw40oxPI
JBL3K/yqmPRCmrPSzNJjXwN5cXNyJmTk1MT+2lv0Ox/o3ZUZTOKRtAt9gjyndvEm
Lkof7ZvdWU19CP9P+ItYpx3jnPD53NB/x6uEqeT22O2EPDFYAHyoFW6x5dJODYGo
l/YrMp5ZgnRkr+HQsOxDNzkWoIv6tFfgSkULUhPXMpXpmOiVY88qPx85K1WnAd7w
rR9p9wn4FlP8aoA0LAwsgUSOKgYDQu4EmckQ3OVS76XES12prcTI7mrG98YDO0kG
wO8hS/XexQ+GhQ+xgHWVRNewbV9IX3DVwmzovgTwZQpdo8/KfRMfTeEoreX+gS7p
If1GcIN/ZzYw70yKVt4hhalNAr9dBfBj1cIZOOVOcrYxOItSsxhWMgOJqjiVji3x
la2u+1kDBse+cvJ0HdwEIX8RXQ1OOYbQQdC8gRsU2nGw3MUzBKi6g3ldMXzMgUwE
mWt21elIUKmS4vdekcF0DbQxfn7ZZJG91Bi483202E4oed9tNQeY32zcG04/wv4J
m3IOR5+sX9RQtXITfCEKtsaq3qepnSaxzId+7MljvKRUCdh0oyWiWJ2OVx4RJwAm
3fD/k5qsWmlDWf+VR/1wyzWOIQAoC80p04Dz4Jy+Bpw13WFrWvle7YTiP/Q//2yJ
Ij028pKZHrj8vGwON+ACYKZKd10lVEqWCFmnCFPJoRH0w7l2zkB+OUeNCU+FaIJ4
o/UIewvmvFn4DCq5sB9jbO/5YLu0kKTEWj0AOlyvNWRbB8SwInwG73kF3SdHffFo
oogcFQ1XN7x9mN7h9LksSFWmTsGWhEr9H/wIpXQbdAs0Bn7QTgXKVX16fW1ahBgn
9Vbg4gAMb1dS6RkucCqf13Kytd1fQ5mr/WCPCruznLbwzaXAya3RhvCVbJStk0ys
Ph4biqEGvdUwKnaEWq0jHtiFH++BycC79QmaywMX+IPRxS7aEEeqWXXr8961xGzd
ZTIJNhPCHBpKMlm24CKEcT9I4MfRdPixIKsIu6fsaI5j3rIn4AyHG0E5deis4ATQ
GoqrS6uoix3CiKBtjS5pqDsYAx8dNpslrGjUAfcIrgQplBYDZSWnlD9Bsgu+hm3E
uYuI80qAA7/a1Lrz5qO6fqw4SesH6rWCriTMZgY0d8oZFQJcSEU6iqXHS1VWZhBX
994OtjG12KcTDBLUs05ZjK8Nbt6f89Alfk3rh9AAfMnFbSBE+L/enDu8r25Yysvj
fqTtwyc5zMlj2+BSrmKVXCoZ1/UO41rcmmUa5cjK2WrQ03kCa/qsoX4ddAImdhay
Gz3VQ8xLzI9/oVJ/Trds0Dz/UhqTDginccBvyXsE0zMVMIltZWEyzvUCN0JMYUdN
PSafWRK1y28HeVAohrEWlxHxFgw5sQnBCzzYtkHkYhG+c3oOn1I6WDXEYfLD58bi
nGUFpV2bUlgf3StxxT2ZEP1a0MYpCK6jC/aLQpFFq48AnUeu15+YZbNQL7FYK5Ga
nylRtIFh88UK52M07U4fpeWWzFzcD2kfGUzZKwQgmkaeG/BGZU0kw+hajRCjZepU
1wm9aqgQDk4fU1+ox6ZwhjIX+DPq3aOr1SHbVf9fiYbQlsG8VZ6rrsWGhM/WXV/n
Mo2V0hMLH9g3o+f8rSkSilB7bM39Y+ptdG9HLzIT7uQin9z6nTgpyT01DcSgnP+g
nTpThZ5lMnqvzTXrPs0XbqPahCodjA7oIts5AYhITKeq/aAAyvS6tYgEDLzoTVWk
ktWPQZkJOcIdkSOAT2y2jESrNMEyP4XZgfRtoG34rzXYrU2ZpjJhmN3LgguOjaTN
kotIvzZY7nPEOPUdHpnodLGnzx4vdEfpac2ocskRETLO9MQkBXMoEl+XMeoah14i
ejmtKl+3sYBmio9iZECGzHXjPyefS6oaIncCZIp+Bpd6OqDpzmKaQB0RhJLAjNwA
FKZVYncUx9yTwdNJFOt48IKxu6tzs2HOT+1+sqZ+rdMrQh0dUyLYXM+IJJstDohC
BktVkI9IKOZZpIWwGIErlAyD/KLI5HZImHhjigmS/sKuH07KLPfaO3qUYJzsNZXO
mL6lTD6nttL5pSQeS1SvoPZlL0QW2IEL4yFfSJq9gbSDPwyBY5R+ODd0hlVRpOLl
mA/bz6EVpuio5rdDcX1d6j/LLc52Fz/xoNbltBqr+ddfKSnPWAHITJySFBeSPmgs
+UgD6vVERSUksg99RU8/41bFBk6xdFWioGCDTP+oJVJlXYQ4UOMW+Ykehb6mVtD1
+l3F86tZ70K+t3/HuDtvun6d7TR+PyuuFRO4Ef4LsRCQfd/o1Y8ZH0qEobTeXwjA
e6VHr897aCnR92chHPRZ6CxabUmp+uuFLt5vNf/hPO+EwAssvHeJQi9QCQ54bCMy
0PECmeKkNJ9MVlX/SStMid5MXS28MjkaAaKzC93FgjMP7tcjBGFqLxdRf/bqWXHD
fn7rQQ0gKhy1jwuoce33vzt5Wj41jbqlcsdhK57JUI6MDnyQ9giKrtEl6wQNBO18
wvUZVhM/v4DePq5qFXl2qjoR/I/mJQlxxphGhiWsFWuIPJNzdMrsnIbwtGymBt1N
UVY9EZuJgEZORJ9UvCEO1dCI+zyoq1ATXpi3QTspNXrOx0RM8wU9tRVsP2Fx0YCQ
xL1GTOigesmI9J/o82zbLydSvFzkoEJR+ydVsr32VlFQCyL1sl0Ck5/lUooDlJWm
sG34RofQymOz+YoiNiHa9/3wwHyV+nsEBmGtDKa+SJWDnKV26nH76TIIJqupmae/
S7vg7rB3TeE0+ubYz7U6m3oNmE6UHebjtNiSjpXLXVTfciZP3421Jb7WnbkTFqS3
QeWtU9PYMQU6dH4Cva/Angi1PO9lWi5BSNg9lzC8LyJ+iZlASa/dctaOIC7klgzI
Yw1UYmhp4PDbEb0kvkaBSxQwb/kvbR4afuqtO6s6kRISyks6m0BSTho2Jjl8ZtfJ
33cxV/b7X8A+AUxbIXSpRZGGN8A7mTrxuJSPfQw2UhI68OAq+KFvlfOpOjq8csfO
0RPlBm6Tt/oCvl4hbMbYNHdPgNpnew/XnXu2JrkwCw6848i3c2lG5Ssy8DT0QLfK
XKDuc36n35qP2U7V9Kuu2F/ojdlnvoeaZpN488ue0d33gtsAiGfT9DY5Nw/RapZy
r50nEFGsijHn0oNWZ3LfoaqLuMiPy9rtLiXKXzibL5IM2CKvNww2zm8jB807jm9g
8PhUH+/O3LRnNccdsJbATeHPYDc5HVUWJrhRfH0yB+lQE9X3phTQOS4BQGwGlxrq
mwVQo80ChcyhskbGBcugbTCpUBIcYhn6FAubn4myDJKvlw9x0x9IHAMHx4Z6vxq0
I6nPjaKdiXECyP0O7JNouDXD0BqsSKYxa+idVCC+68UnX1YmVsbID4jATY5d8JbH
EmHLLSQ9AQQkHbxkxeCUzGBwZI7ovgRdGsJVJePCsb4Q7EVU0a0AN/fHA0QcpSMr
vkgv7f8ME8qE9GOKye5PCf/55mooFbUGYsDfn+ftIrnzjErhyEWWcM495Rzon3LQ
zSrYQCPT2ZN83NqsHZm0aSTIcbQ7kciIFCiy2NMs4Glk8MO6kMAZPbYbRvEst1LR
EE1UP5Wr9H//Pxs+17ZB++F71s/KljL0+TzSy1htnbM8BFd3FwSCnl6taLM9AkKV
fwWK7+KTHC/C3Q/q4PWPKKQMtTb15DZLQGRw4wSVddPuoqCttToqBcQ9WSGnOnDJ
y9jFawkjDgOGID3YXyAtYgefLH7A9vwyvMTlGB+VWwptIBLFG/S0/1WwfH1zG9eT
nvLH5i3ab/DXzxR1JZmXXgsViU+LjRr+hq+QuhIF/F1DuQJ/VLlmmv3mS9aDdGad
CYFwT17K2Z04Hr+EJ4in6/GQcCK/fj0HEAFVMxZEqvxZpF9+MTV+ZFqX+qp1eAl1
L0r0enkuTmpe1aHM0oKf1cMFiALmRLLBMzAW+83+XyO+BqSDqtgqopVAzBbxjxHg
T5r7go/LEkm7sslrwAMe7/BiuAlyB8oG9m6/eeg3l0zXAh/9hYEemtBRuCQLbUkl
Do9LDXt0ANm31+cV/jeusdBhtwhlIaSaCjYZhMmappWNwTryDEDgYejuE/2YafsY
i7GFBLro5puEQIzSCO6dvEbWqLeNZp8RL4K1HWq++xLGneg+J5njAfuDbFCyGXlL
C0z73DnWDI9yb6TDixj4DH9Dr4OaWmPd6eL9/RsgE/pOxo+zmUdk0rjdHkuwKMOT
V5RySAT4z2CiKOj0A4B8BiahaRTy82mZA1/Jn8lY4jiQyTV7dp6SJDrdW6KpeoFj
0FaVolWhcFVrauyGZ1PMJLsLplyKvy6QKcIM5y9MBXv7F+0C07fjU5m282V8+fFr
S3zWuibLD74I56vxajqw42DPyS41x/UFAn9j1BF4gVffUcPSsjQMzG9wCkUO/PNx
q4OCt3limDnrctSV9HWWjYCGnbXXxAcgy3Mh+f7kBo59MQLqCnXpgYpncy0TWJJA
1uEVwlMqjNd80/METoZdmcyoN4rQBLQapl9OsF1sZ+tbxMbGKqfBLmUDI0qhXUDH
c6dfaKxFT4mA3EomaXE2sUUXaXf0oyviKLJb20yu1tAo1U0NLlbuRHbIl9KjM2rc
xzcuyB/gsAqok3mY7JtU/Vnd7/ojKlLxkqB9m83g8Ve/SgD0MbxYUOsC6nqQI81g
HJEPFetsqFiP/B9QUHZMy/rmB+JE0VVdhYSQFlu7qEgiuBxk9C5Yqo4y21g70ymq
3WmPgdO0fIfoctvFTkDAaKk0j1neD48baci3S68yU0Q33fpRVEnKULwf7ZgQIIRm
ms0a7XdbWEGZcjqQ5ZDur0xjFMLkY3YmudiuKFouqHtyF7a7I6Kl4KnWumH6+uTg
a/Do/i0GjCCa2fIe1OuXVKXf3oWQTso7J4qhSj+/YHXwDI8hVlP25I291nGKjMI2
oHHu28mDP6epZ8nV/StrO1nkuTaTiwf3m5H/68xNxTVbTfFZvdL0N9v+3PfXZmja
AyrlsxMiCWeDMyUZLtB8UNOdonAY2h6ugKh214h+MmFiBB7vvFwPlGinpQ5k5tDy
v9A1/M5X61iEdoBDN+uJBLFsTNcKs+2GcV4cekTP3bhSGYzEZzMaKC5Y4PgsaQVc
t/9RU/nV7S5V8OcvInfSo9kTW6tMD3CkZ0BPYyjZoxba9C8R01+Qzycaar4yIwOu
xzK7+FsbCe+f8/ViuK6bXDZasrdvV/3zSUVEToAX1OLSa8eoZUcQU4lC71voEgmp
h37sPkpJ81CvFSlgG8bhK9f76lA9vqRA2kqG5CEQlqWnidKjm6ypzsUAiciJftEz
ixsJ/68ZCBfyDMs7HWeakaNjooHjC4Z2SJRq/Z5x4x6Z0qCbiAi5aTEGHn8xstRO
pFTboEAmnmSlXoqfCi9mfsYU19FT5cliN2ienYef44YpcsMFQlqkfQkyAPTrw+yG
KS8SktcrrFCyG4OxAbiIVx2NatU/7UprRdeg/bWh1CJALHmw+6pPzh37yWXQjWzk
nI3zsfnGQAt5CeTJjFzLqULMTanWhtbzCY3T+sE0KXzRNsRw3N4SknagOGIKn5hd
hxu8gYKHOzPJFNk5/L4H/6YwyCdraLQ+Wf978ndG9gUjQX2bx03B6wDmGfFFeDTK
YUIhPmJGE9nw01juNDNKxgzC0pMrRmHuAH0TQee1NuI/eRqaOrT6PjXcF8b14F3K
djRzqCn4bb/q4g+3+fX+Sq8ErEvctM2cOH3/dI4WTVdxj9T8V3X28ac7BeLjwQ9M
IN/scf+u3Vg2+tMm5Vcg60DjM8vyHIRFe6Elj2LRRGiFC7rA6OcW/WmbshbTezcu
uYaK+BfkK1k4Loxp0VSY8UIz9bUBry2ITLTE/30vFuZ9z+RhekbaHJtBFfBZoFCX
RqidlyXxvYR6WaUpCIfjj+REbYrAaXoyyPAeN+wlYndXq38TIWU/IIS/GUrL/FeO
h6IiZF6Yzivc7e5QrkkCQgpOA+Ii3uTOByJ+OHAR2BRIG89NlbJ9gxEK1pRbVoMD
ftfeMDlyd/w4Y4PeMy+DlGBAB9/rPk+Ty1I045IbRvDydh1pw7+JoQN5+eQeXRQP
KLZNe+4kleDZfFwdOU9LkFKwbfpkJaE1ISDzXvkKGBw3KDaYGd197KnZpZxfh/m4
eX39c7gDkqFbqdayB165kHZzeMdgQErx6Sws/0H/bcXOaV3nffliIxu0WeIQhwuh
fTlQfZ2uxfLtzh/q0WTbhAFncKWzY5JXTQ+ZHByDmNH646ZWbC5xRnH66Z76/Rgg
1HdXCfRd0YO3oldPKE8YpnKuBcpF5SR7+8OsIS3APMd5+YrCMfhUdePTYPHHygFo
/9/MFB1fpN9YsvoXcvEH6x7f3VTYefbrKHnaQPvFVzjdK0w94WXJawmhCzlejwmW
66GQ9SogIaWiBaatH1SVo6eYIh68I7MJv6iey6uWnlSfP1qYy7UCwZRrA7g+4/bc
55kA8QwvhKRpayfyl/YUaQvY9DEL0P4H5b3ILOpcP3QGnU+/a8Sb963MJj4ZTsj6
a63fiGTRqos9ImB/di0T/y+AThYwQaSjFjYTZdTXGhrgy/ek3f/P/+IjDCr11HPQ
jluObzPuSgAmwcLIuJc7qdQgGgo3wQFYJZp76n3cjryEsS3jmskmWjNc7HI2zfQ1
bImLAbrUDhrUNGKwcCc6SlJ/Tt+JnSqPTp58XamawSCKtaZgWzI/eb7TgrhIwpdb
KFd63Q+1fVVOL5cZ0tKBheBuI+LqosFYLGdkI4CHlpKYFMQz7LHR+DE52u+ov0x0
rinDoSywtomcyQEhj/YV0L7l1NJlOHAcHlyeF2BK6gTPdWXofGNOhNaYnJR1USMP
r8vykKBAvd2nCrV5KSbVyqYkaBnclNLM3Ta4546TcYCJxiklnekruzCRmdxWoVyF
fhCHhweFJhAC9pzb8KfWOAw5HnVol+Br38kLxbUDjw+vuFcjc0KO/xFKUXUtCAgA
qm5rgFkS2+UIjC7PPJj/SOi1IYHCql9D4JQnPsgt2MV61r/TpMXIA3MysJirPyCK
4IVFCIzcfYnjcRAgBxs468fz3hucTftMUddaND7cBdaXQ9r/vQVymqmDV5NoQP8K
vQYVOiepIUomBA/NsmJRkwXGER0ug4rRP/WymAvsH2wl/8BcrCwmTRPwrgz5HeBD
if8hxHikkHJwDEBkhv7CJQhSKR35+j4eTu8YOaWTYXp0NIWl285ffzvAUMH2gGQh
U01OyNTi1Bb9h0as3EHXUu3QSVd9iMg1Yg9IUJmpwXwoR83hv/qzfa9A3gO1hqEH
W4sQM2W9xi82Sjo2kVEG7m27erlHEXm/L8Xl8tvkzx/ex6mmUqu/7HmQUskw9Qks
bSWCkdlbl1Cvfm6zNUC4eVCeURNFZbHbngmmCrXyZKmkxwmikup/3kpoMrhc7GGj
DVX6M6tgevowgdPH2plCdFcdjAPy+vzZzdfE4zg9tI8s3I+VxGYBz9WitcIA1JkQ
eWqb6/piYlSNJGwL6NBPBzYjphpXkmN7d7KN3q2U8DbkIcf+rGqpJYcrBpcZc0Y2
wFQwD7lsZ+W1j3pDZP03tDcGAQZvbL4iOEMgQYC3SwLCs9QE12pPx67t2dSD2Hc2
XJckRPb6AfDjEJDnpLkqPIQkOzdO0U9sKww+1oayz6pKeoJMndoJu4lFW3Q2tNtl
G+gq5Dk77CPpZCkNSNYuqT96svLD6nNOGFjp6SatickyT9kAvsRcjE9jp4basBO+
NDVsp/Ft0NmiG6Fo0UN6rZL93wE4iNLl0JYC3KCl2znHnJ6dpum1gSlDbs8L2WO9
4HMm5p+ISb5J2CiFwJjTD5YevMADerkwCgFkEXky9IW27Nu+e6yjDIQJq3x1EC6+
KYj0VemxQXmjNLFtoSAAKXPISnFUm47VWj8251mb6KzgzpmGs38bGFVpXM/wD2Qa
feEgH5KhUAbK23ExpdW8tKIOwh5uf9S2amTR/PO9aGdFngk+ZAGUR8KYPHTs7KCL
Bhgoh05pS1HAVNUO9QVi62nraSblyXQ0vjCGljDITxjIbpLQhR/b4/rHo9IpjsGM
erfiArCvMBFCRkU/b2fs/LGGBnIOPmPzGAqLa7eN4NM1AMBCav68/eSeUIIE55QM
05Jq75E+F37k4s7DkdSPybzx5HapVGPiXHbocX8zq7ESLS7iZNLBaHg4Vn6Jnd/S
7YbMoGH7l7XQ4XtQOv4NUiw3eKLX2qvGuGalIEnjaLZYBvEqcVajwOv0cS9Hxxeq
vT43RFP6a/PsR/Zx6tNlpWgWf1RBPn0ZTC+7JVK1ClDSXJ/7zqPCwo6kCqjjgp0P
gHTgiZbroWzog+RQyGJDDmsRFFJ3BaXCJ+7gcbwWjPCOiuzhCMiHbYoTJjlh0/Fo
jiX89n+4k5S+0aLglQwsAot9ySRYEwFzvEUh/pBLHGSGv9FqYTMY39hFxRd9z50X
kd+joRUMA0wsdmJzvBsx+jwCTgi5TnmsPKeEfB6FFeeYruZJVxV4aLFDax8VDkum
HhYrSFUneLQuDiuY1G8O/m3PtHJwBuh85Fa1yGrAH0xag0/V+42Pja/6t1jHfG8U
WheolK8ThRM76HAs9bDbSvDM5eir2MW8/fiA3WBHUYo2hk+LVU8qN68DI+aKdEgr
4ypQxwIXj3wWtnHhgkjc8Z6oSKq7SfVCXTIJmBNlnFTnbufRzPa8e6uzEELDotcv
TGTSrDPuxpp6PJS7b75vbzaNB733SaOPzLCeEbO5rb4Cdhuh4ikdqcPwfQptUONF
hWC2pLGFhBRCTqY3zNu/vhCu/PstmBFp/f5bJK0PXKJ/8wnlkw6fBnQhL4PE8dA/
mjcq9iq1cs8PXUMIWFRrzytx/Tv9dWq67bIrM3LBQGx3pKFXM5VkBsEB69hVIoNz
sAQr2GXQCpRo5ZQPUSs3dTxBBRWX8GMmPC5CuHDP3maUxfXkGLiqVcgenb8zdAgH
VV70KB/CKPG2+AuVTh1xHBa3w1L8JDIMtG8LDQg9LcBme8KRY1JHAhqjXHY8OlRZ
dudD4gu/y8co1WM0fQY7livMB8vzf8nnfu3e8o9mDe5NxJph9J45/tsylJ+RQp2x
4+Yq+Mgwk5Zhc4W5w5HrBs6TClaTh5xOr+MsRA5vZcl/k5BL/5/ra7efhc1zqAKb
b6hw35NoEU5Dc95ocO9+XlntmE+4Gi7MvOPS1IL0uifXke+1iWJrfqc4rylJIMnk
Jbx5ukFTodLudROkVhbpibO3XQ95avmIRps1/tQSonjk58uarkAk2uq8lBM38lhu
Ew9xsA+n/jBsQwFx4yzoiBgirLrBE9ijiFWidYwoBerwJUwasEYByN5sm3l1xunG
uaXh0fbm9WDSlwWkuh3d4E8JtA9M+IjHjtcrr6Op//br8g9vnKRvQCeOnMmEp82M
Nd5KKVqzFfy9/oTvuQV72AW5WlqGD11Nfc85Eq/wM82Gp37dQpKlKksAZrp1K1Uf
PA3dA/Jc/at5H9xb9obextwq7lW/03T1JDg/Yul5qjFErAeYeyBODGEZq1ksEBFm
HtyWOKxGIK4MGd15vo2XKOTp2B06HUzKkHVDnhQya+d8gBBvxIX14NpzfiqtF7GL
2ekBSAGRYkFAvBed6QkcU0SE4sICKaqMzlyzEOeL/HoV4ByTSlFzu7N5ZoBCbGI5
Q/mNazG9NZf2wW9K3FMIb/r7hEJHnEYcGlEYqzZAYLolCCZX/dxpjpOxSslLFne2
5qiuOSUQPuI9IvgIfnP6xCe2nU6rjgPtEUAUidac7VmIYjAaZSaE1FIrThd7u0Ux
hYnqOw3HF8YaNhpTkDz01sdSjo5vn1ajxtxL/zMUxoZK66ukN4FEFRwKnj5GGS4t
PgaJex7QdL3RM5QWUgqJs2woer/QGyRPx5ZG3aSn/WA1aPt8LLfZLmQUp29Od4uZ
QrcopmJ/Zum7jGKDSTSMzESbzVJiUeeBmIVW7ChTC8IvDYJEiDtyVN+1+2qLt125
xBF7nFr9Jcvshqfv/+FOnGg7432VoKQRWAG7R3mWGdEzHz+hQpDIUG0vRpGxqzH/
yulcb+R/e5Ap/oZlMFs79dS4V+uknPBKGkqJZgdZt0GQGXSvc7N6+PO8+luUs26P
2cA6udkBtQSaB1NGknGOEgmP0rnNQx+W51rTycL3iOqkFazUxgc60oCjk5LM/mqz
P45DtWmT3f0DK/rnG5fGzD8D1R1L/rxRnX63UcncnRNSFJ7fiy7YSho33uQDP3n/
LhOT54v2Bj046shV+OiR7mTTdNEithGMf+Kl7GqvIr6BCqNSwMaI56ZhSGhEEF5R
Cqp8JylkpBVbpXLb+ZiHsAmJeHvD/wFzI2CbUxw8k/7c4e4Cwz3rTpky34A+6H55
JJbWSnAqDZZ67NCUJkyv8Z/193CcXA31lGKsOAJsBpJbOsVlD2lJOfkWbCR2iEv5
4HwNemGQwtYxtrypczljscFCR7yWZxddU06y9XtGEp1r94qGRnGBcuGr2nQD4Pxf
7VMJ7ohdYcgxsd2uOZ+r7rMsT+8QYxMdWzWppW1Dl+aqbeoyzUO6DA4W2vGAmBu/
bUJ48s2cxcr3eW/8INR1N1gJrvNU4DRemWFhxNkwM59Pj4SzJzjY2ROQSetpNXIV
jf5lh2JyT1vENRevY0bIfd4BCrEC3iZpSrNqrEigtc9vorB7vOzGLvluDLFdQod5
Y/9Yc2u1SVXIJaVz6jkRcYwNMxb+Iv33IVSbi4haBzk/HvvBqoPH6qhuZjaZabpP
5TKZznpxikAjpX5AavyI1ymiAmzSFM3m/5pRevm7P91CotuJ5oZpt/uchtxI0gOh
846s/2SttZTStBZXh2S782sMDIfhEaRjsOcscGEzqARW7N4xp4ccc6si/2NYTjnv
w3KgUYnqgvsalJYy+Dapc7r+CEeRXyKmUiYwg3s7nlbA6JSY2hj8Q0KmbndmA2Uy
s3CLoBLTO5VucOle8yf0DPiwbXWY/XDyNREEVBN9mg1WSn85dwO9TyfIlsTgtfsg
4YukFsRg07oyrfWpOXKFCzc3NyvwEKA9EUMW/Qjm5/SlI08Da9JCJtlB1Rnlbers
bWyVUS3etJA9+XInCBy9MbUZZHvHGSs51c1kdWkheM12Gfm8WiqHFpCY3UFnOLdr
+5H1kr4R9bwWRxV23bwRg6rqUg0bhzFu1YKHkse43jzSMbOOfIy2/b30cVIPfdl4
mPY3+h8r/p+ZRihPZgBApjMIK1pixTPXdNaXTVdHqL98keVpBhUMVxLiXNB0RA9Q
1B8yEE8Vbi3IhGi0fCmNVIpOCL8VKb1d1KwmMxqx9wu7J3U9e5Pd3xE0Hg2gOuxr
YwiSyLq0yO2HP5ZUiXQ46LJQH3gi0FP5e2MpbK+Ml7jPPgKnYm4EzQgmIbGkYbNm
`pragma protect end_protected
