// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
SIvBD2WzcKktqaQ+3kXhlioJwgNZ4sOIkD7AUImlAn6YO+Ou0GEJ+PRxBokm6xZVx/dUKiNbuA3y
CMR37gMiuzjdpFOSRbjp+L7ROSjpKGMnCdirRRnQZCnG+EyL+FmJcqtwtqiMYXQejmLDwz4PnqRB
GK7FHq8YCkQoIJUY4syasaqx+vYdtPuex0e4yPmP9ebP0BL2Vj36AlwJ0VPqm0szQdvz+9mvOqAe
fjuQSSRgly3fjcIElfXlW4+rClUqqGgOS2c90JQaYF61Jxuw2W9mRUuzyVzQhxjssBb0LDrbuMkd
pvCmshInf9mqZ6brBPIddMc3ukjW6Fk+nD55Og==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
wlUrRcK3TZYaJwE/hUdskj6mtB0+1016La1XCcVk7n/LTTh+Ln+1/11JeGbERGCeZq5cNrInkVnX
bUBMuzApH/o/AAOaSnM5n6uY4nwfmmei41RT8W55Yx9tFiBI8hMvtb8IFFG1IRDU6BK6uWiO0seG
IEK6t+PXWRRJdKzXA/xvZ7fdn+jEp96+E6jkSmsIytlOc/ggG0iX702Mlw0129VN7aYQcl7FEOEx
ewYbO8gmG3y/0QrqRwYnIbGitVTTjDHbyN1u9blE5/mmmIEuLVUy1p6h1uyrlp191sjaCNvLsBKT
CFORZ68UUUJhFdS2u0Ms11/MgK85JggXgIDTQFFhD6nyTCr7qfZUiGfCs5YVMVwL8JC+HbevPzO/
l+xkM0QBEI5/WDvnQ0Oh+FOlLtNVOkUYvVgEl5deVLuhwswv7Ku2czv3Dc2lFbOQYYH0WhYDs1Wt
n6dnxGGfDfZp7j1FUM0DoSQW11sD+iVVscqyGscWqIK3B2G5SeRIfIW7/1d2F9ltnk6h4RoEm+5m
o4aJ+lA5xxIv0EMRFc6+kl56iEM4GX0s6D6nU6iTYVdbNHkBnVqHLGHL9DirW9JHQhApTZqkrxQW
Tg1o5sGjzjUcXdkyEvmZZOIDx/gZNLXP46aFofDfljq0E8NwVe2Nvu1ptX4V+x6sNwwCX93FFIHT
75L2/dkBXjZnN15NV7jxFdffPHc5gm570JxzT47AAMuucJdr7qJsWsBLSBfud6FzmTHhLsXS7g2w
VirT9sdNsT3frBAcwwYVv9NJi80r2W2uaQH2FPaC3mQryqtaE1F5+oSL4RetMPmXv/uq/KWtuI2v
NEkieT8zgVJpy0Uzg5V8gL+l9hUOG9H1nJEbWv3Qij1XvLOcMFFS0epBY1lUTXsmFqbue58/DD/i
mZCq7DhCnPe66y42cMlON1JuV2w7HmppTKSQMzp2YegVwWV6wxUHecFU1UN7T1bArVGQE92PQMTI
FznmMK9G0a8ivy6XvtcKtmuBU1YVHRgP57lWYkg48Dz4CMYj0VuoCEYWGD7tn9ZEqkLE5hq6m+7J
r+4qOtzGvb0whJ8F6V7DfzmEM/R0Zufe1YV8Lg9imbxSykxgL9zuNGXjxUbOsgmPVIDY4NLEKA43
pZNGGZ4viBV9coKDZ6kmjXSaiJfcwU+i/4oNOWvdvTCWKsLMCo3BcSf7p22JOdpXIu+hIr7KFbBx
CfLj8mzE8NKEjTKtFoQMEngbH0wyvGuTLqkYGTIxOTWccdLmcFS8dhKq7yO7096Ct6KfowVfZseB
NIk3mVCxvrw4NL0b4ZLjAh+dsx2uZcQAuhGzRfPVG8tGSbgrpRGBV7YQ1fdtUZDUt7JUQIIFIhLl
S5q1H01YDRvtpjMCu5Q7BahVKhcnzSxEF+WAJjhwilkAexilx/zraElMkGDPvvI4dVF6pWWA1y5m
6E8MO+AM6WM2BUBi9Z17qvugFvvPB1kh2iRktexGqAU0l3+eUxQRhq9KZ9Q+CKj2D1eFo3+khWgg
IYjl/AHBQiHRoz4hmisV/3G+PfcZKgNV1EaAUkflXljP8BuYiWPhpi4++yC2JbIRDXxFUiB+Uebt
RFrhb6K4/X0FjzpP1fQG848nMnYhJtsdd6ZfvqG17plt4s33VgwZL9dkREEAIh0qyva4xOrY3nE+
ltpqtY+dGnbL9Jsfg+nWQZqQAmLGqgu1hf1QTTDl5sIiHdFYQIhznwTge4b2Gt+ZK4Ha+TLiOupC
f2aeouBgnggZnHc4IGwMK4TyvBghVtWQOSfV+bJ1O87fZQW1Bi6ox1XwczoHt9hPgN3WA01Sq+cO
R+YBtAtdLtR8nriZLYIwv2PB1xCTVodc0N9lPCZJ1gXysyTdirHZ9iq8NeBJ3VxaUH+gHwMmixif
hLV4cj7CW3rcDQqAr4dr0CBmMtVUu08ayMi3IgLxaIgfObLGYmebQJrfN33ehl8cenvmGB1Bqlcs
u5NZQV65chl3nhOCepeq2lvh2BN/MwK6q0eA4r9QFVXrWV5tI/+ZuxrLIWKqUJRRSfBzTtr9tqaa
uZyvut+QohnWqHhhrjQ5rM+4YnGFypnsQq8LwfXTLy2Eyuo9ymukdgdF8iRkar2npLu/BSa60WlX
B/ho6E9njHj7kXd7AFYHzOuFRxvq+WkGPMz7x0qHgbS72o+b5+2xGSWNiHgOC960xL6UAbYjYrJD
0pYGbZz+vnG92wutJTm1fVH0cnY2beguZgkHl08AvP6miO7ugzHcCeWTdPSd3SQBlgkX7SksOWqe
svpu5R4Rc0ouELuxyQpaPNG8351bKH07f6jPyMuLkb7hEYBCE/rOLmMZqt8alu/d3nRmlrOme4ja
JtjO00JMnB22iP8yLwyQn3qipjmxbtHnuL75aASN0gLTJjMFAUW7WrOq6anZRTjLkZ0nCfvEtRWI
RR4pA+o6Rlkio1qu7EA1kTDT6Wz2xwDFpheViwBU/nfxqtoB/eAIq791pdUgdL0bMwUMYZTlmr4A
jkTuCJUebjaU7FQbliqMZI9Lo9UBJMyxBwsjGMVuVe4/4kUryOQjHesc40aOKbSweTGOqL8Xa2XA
T3eUDvSzaMNRmgAHNisZoDNMHI5FBpXQVyWL2GOv1urPp37FjJNwIxmyBxQHSaKsCIoAQhCGSasd
Qg7PCdpQp17BsaciA0yfvgvO5/L9N2S9057Kpmqhd6nIKP2uGjknTuNGSHd7gACYOnpftumzryfp
9rZstJYIkcufaOdhf747UVmCNzC8t7EV7UXxm3Sx0Y+4DKWZlsPE+2g0ZJ+YtSQSQG1sZX6xCWxI
91U8SN3HoRynUngzQRViqHysxFXdlbqvuW0lbIBz3uyGZfbvAu2u4udW/VU7pMDZjW8XITzvZiBo
dIaCj0zzqIjnJPBtStlKMy2EpQ+VI1TDqBwezI4K40uQknpdqWYLeW14vfEBiOcV9WnjU1vaCKhQ
Lwd2ulxCjNY4xybxtVf/uIb7YgUTW3CPbjo3nUUKtbBITg1azFg+T5HLG1FXaqmfxypg0Rxw7znq
EZ/cU85wsu4mo2aoAQe1BZcipq/qGLUinAFklmsIvxXJAt1I/HD4NKAn88iF8Pu/xCr6v1SRpFcW
eNgt0bE3KfhVbu0efEhfdTDAuJV3a0QeumI0ScICVEgg5TLEF1uXLPfNkjXC1TWRAQswCzsB8mr4
87YwavoXXOA7PiZ0ZwwgR12lFQuOpLoU8FCIf2WCXXElxnM+CaAGvIDOx8HWdv8UBeZs+jfM3xzA
6fsRFQ0gE9YEyPbHVfQcp8EoW0anIhexZECSxgqjA4hw776eT7pZXEPFqXCN/HQOxVSJ56lSWgec
yzihk8PB+H99aFxLitkpjgeTYFEy1QOT4lW4TnOFwsnz+DefrrYncnPNwZJqxMndNpqlr5e5AfYD
UwIvkJ47hPy/NETFwSViu+0GZr8al0cfCP7Pe+JvbHglTl3AYaDZ+r0SHG2TMygvvdjAzXbYcenU
pXfyfTE/NgnnOAwRiKolZTENjoEkkEBoVffHXxp4vprnJbL5Ioctbp7HlcFmKYj6WTe+NW5Nw8b/
ObSV1vVwAWOoFmaGJmZiSeezSm/LdEmQBWdNVPkF934kxCfauA0/XRqleCCrkQ9YaZP8Y5kjSz6W
bOUXuE8DchRQV4XOcXUuHFlyrCtJCFNa0f9VCqYzE2EGr2N4DYLR4fOGp5p5xsHgssgpOvLW7MQT
XPWn+uqCL9DAokn1/zb7QqORxxfc6Tm8Z/sZWGksXDwDX11Ez7Z5bRa2zeUpPZnBW1BV7pFeMSdg
Z9Xv8F12iz7Bm605ieyWEz+FE55RyDm/i3sc//RuivxNO8N+5E6ezTglW7LsmhEaRPCKg2hmIHF2
XoRfUSxh8P3Bu+w+k7+88JLW0+iDVWzrTYft9bBLcyVp6iobj0szzehURhP7Y62DOkDu9aYHndtg
YwnniTfnUp9nDjxjIH7SAwP59qycQgdojwodyyVG8QzQDbsLldDF3xs43TpJ6xpiBHkJv1q9JCtt
fl6UIphLKyIX6l1mQqN3I4pBBpLndiwxNsYMw2NfnTzqa2+JAuB0QHr1ile4noelhW9K/hjmTSBq
E9uh1rXuWtV5wSHNjCc4phMKFWR4Kxgsolql3OajsS2/se8Chp79RvoUqe+NfUz+H2WWzZaEtYBn
SWUluP14ajgaRrD6xIxDp3+lt6VUBPMZXWvKe//7lYhQ+lIZq9OsKrvJak/WCbi00QmxYTcu1m85
TyO3XfJyX6yqCtAjvsIjxcM9DcHRYZVACb351RKcCkVT9EHjhV7jI/2Sc1vY+jZPpalCzwD9o5Mn
M2vrCtL7yT2eZQnHjABSu4Ixhvem+h/FeMCYYunr0I+WgDncxwbectJI7Rl0TJGsTbivA2EyzPMc
BMG0Om313u6IfWkTncEoaW19xvl4JItIUOR0G2IPMKPQ0NEUQbPOw7HswuZZjOGftWH5jZXAGbsL
7DvovFPTZTwX8M7F7mE/MlFMJEnHLXwM8kw7uo2SX7Zsi7LOeFJez/SkGM09XSuar9Mj/kIzEocm
WrUoPr9q1tduYwrgg/wksUvr+wLxbHQDbOp/3jcs6UJhHH3k8N2SvLlI7ZUhWDIyiCuVZ3WxLgMv
i0oF2KvyNgNZ/yqp1Kl3e3J8F1/nHr4NidIA5bGX69yXM3WkJkrio4YVIK4+KbK5VpTQGymmlXfT
5qz+cK8e6ZHjiObqTHVVz3MsEzhurUwdsINtmfFGt7+/9x6IcBRtGR8dmHZ2UQXOWZlvm45eGkCI
1j53sOxtGV5AP9kXsoLX76V0FQgLGhVGf9NjZpcBdaBbdh+sbvJ1kcs+wj0StooHLvsj8yQpfTDt
EX/CJaCUGJUr0yttVlvQCEWzL4i3z+2WaJaDDtt0kAKIcPRnXVJN5b9uNq4BQ7WvoIAddVAgd2+t
P7jhfF8ZLqqT6zK2M0AeYMVWbhOxJQ5FFtCtAQjaRz0pujDInbmGl0ZyOG54zO/dALDaX3V5quWY
ZOWJ8y/edbnR8QjrfvZ8+m7L/wBzPXag+KKQDOvXdV3xBAcmgoKZqCciuMHzS59WTZgAiwaoKx17
hNEGRB8kX9uwMjVE1WP2+22lRXFAFgi0UhfAuaSrWMVgu/U0cTIioqhNe3Bly+MQDUor/kX6mOpU
wekZoDw7qhCE4Ky+KnJTjE7LFF8iBJG7jWAKtsEvg4LmfJWNelw+Mk6IJIfrGTWOgs3pJezFFmZq
8ps8uSBAaL/gdUl9fe2h5tvsPNynIUd7pYisTbSYs44lEUVmyBqAAwOnXK0Dh1WrV6WWsxAKGY2l
DXB4NXzZmMYdhxs2kfrsMzBUZ681yMR7B0dbQCd4YuJ4CG04UOvZaMCXSThMPiMzfSL/Oyy0GIC0
qMgqbb5orysekmkO4pAAUkb1ZBPaBTB4Pc3wFVCjLYOqo7qCGMUJMk+ufrY5OCnHODREvrauuz8x
ypAVTYhsbRW+XzwhFcZMbJpW1xTjIp2iaxEeVpKJVn2t9MHd9gw9enu+o0PSL0DygHP06b2iC1xh
T20ut7bJti15Dy+pSaUaWaY5fKdi+WOqUneHWVRzjIRY7bSgZhDrDN6VU+7gi171euIR6MlAlNiu
TQJQYIYeAsWPzQzBxXOW9GEn3mO9XbP49YPQA0IiPRZHmt4iUhOuDPP71lTSS3TzbFjq+w6WCN4c
zyWgai4FY6SBlNMycMeiBqIG7lJlr3yZ/jf+6/zWLMa+sBSkj0qVu6Yaqik2EHUTJc8vRggULWtw
OTMm9PyX0D7mXhGcjPmJ+bq1Inupu6VDEMctwvnqsWoGjxOvlvwJ7lcXbDEpCL7sciYhidgRR63m
cJHAI+DqwwmekIt4FUK0bJC/FfOT+hR/ZuO/QCwBZXqRdWiVolLWs6Jx+cRo+KSvrix/Lbcv5Rjs
GsVLzbnb0AqWE2qL7s9R9r8Nuhv0P3k/KB9zI9q8dcloxg==
`pragma protect end_protected
