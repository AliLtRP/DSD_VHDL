// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:43 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
MATHSsgexLNkVduNFZSi8dcrPafZ0tMNCqC1b5+jQW8vKxIIEdnCqqieW1SNPsQo
itt4wIetm7lKPnVyFG31faN5IDtRJO54jVYkJdzsT9ccF8ZtkLu5tb4Iv6Xn8yyB
97C0/j8RYqQovt28ouT+rG/RXmLKfr5kH01OZ6Ldq78=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5472)
JuQkiFuRd7OAqVtWO/N7PtN40fSZ6CZtEIREMUC1TtSM0QTXeikJapALgjlyM223
/eveQn24zX4gyLM9uVs9GPI0dx0er3xaIg/0Ax41akSJIq3JdCnqfcHy+Zmup9qQ
ob24uJhkHJ5NJww+zxLxBNqIjLub8ioFAgcwXCw4spamscNQUSwMCuQMXJnvYB8x
JNfkxZQS/Dow9hHokJAoBmAqxsLagGXYD0gBGXrz3XwJ2llemUkO7ezY+aQKXwWL
0vIePG80nCHnPPiaGxA4hcMfHd6n3Ire/dX3iuP9CVzd9gOcTYHIGEBqHNIqtUn5
j40vjRTGSzeprzVhYup9TmrvHhryTDmA2TdKBa6eGrZcAzz9wEvdN4q7OOgykF8s
KvHF86hORPSBB/ZMXCWi8bzhoC2Af6tjKSQNM1N94uKsDzukqQLAlm0neqPrPmlv
tXf6735NqPNx1RLQ2HUJNwAAeGbEua6TY8UdAn3NRhAP6FVfUN5mriMFkYGTGiXm
qDhHqtXGlI4NTflGaClHWHoBru6VrTmB3hOJjS/ZwRPywXdQlNezNYTa7x9Dokui
DkdDkGly0A4SydwtYi8UliO12JPWzUd0/OVvmqtKStixGIp27b6VPaYbH+V3NXGd
6DH9HRQQcmx0sPXahDA/nko73fbif+lfs7cZnssP+E7LDylAPU1WPVhqPndncopq
MA1OotTItqKmCoF7gAiNrxL6h6z05faGEdem7Jo1niu7XXmGAf1Mej0DhKZT4alR
UF3I5270fOQkSGNwyDMEV6aa2KRvASdCklGwsiGgMk6VlT47H3LnS0vSfLpl2Abl
O+OUUGVpKAJjOpdrKylV5VgK7vwJum7hSh29fEY+TVTK2Vh2NkKWdNE/dAS6yA1e
rHY4gNpdcVVYJFipHkC3GSm2WguuCMnn/VsOgAhVZPclrvIXp/xbWapR9sZDMj30
JFJFzs3bq9kbJ7HLcuvUNrjUNEVbMGHO3kqQVDUX62rUQwRr58kJjA8l+bXAptGi
V1SnUStKrHpmPN3ZSUZCOQisH0poek7aoiwlGaOe1DLrvUCRvhuHug5wgpHPmvDo
EslYp6jB1XXHTJue8C6IZIpZxsOIM+Ck7JZu50YUdRT2qx1JkNo1fg8g0BAymuz3
bvGPnw58QQEQ2tmDrRC8NKB41R3zYVDHmCQ5oxmsdwv18KPUPRhnCxaD9VG/9HsH
ltCu355I3b7epgYwSobIoM9a0zvd6VjGOxP3ogQBK9jp6pH4kwQ0amcPqOTN0iKu
OSmo+18p6ULT6ekrsnIIkuMEvtoZjIHGBqJc5kvGR2ZgLLp4y8whD1uWFIqKKWFY
j319xmk/uNXmhsIK75gorgLh5IVE/iWy/qhm8+O9Og/MegfbGNb1RRg03njLNhNc
kPRY2awh/DtGQICpbflg77xmdF0FmroDIk8Mq1426TQ6o3kGh96J8x4+Jh2SJg2Y
vsOSFxuvnxA9wMeQ34Nkgp0Q6O2z0B508d/4xvxKe1Zd8pxY+hVhdlZB7Qh7t7Ry
RWkmZDo+GLaeIB36W0o/AqgRN4BwY15a2qE77uh40NdRWhC7mJvwyYjku8M4Z9NR
T+BTEMDK+5Z6JtbUgC6WEUEeE45NXAqg/lv+gaynjAf344xeD6La6mWJAugz1ZNw
f1XiCxRIosAwwVIFy0OvyVMPhTq+hlVKwHRoKaaamEM/ufUkDoDHzlDlU2fgd60w
DHKSm5BtxxiybFmjY8IplXZrP1uG9SGZ4GTpaXgI/RD0W/ZbhAg97vrElGXYuLe7
QBlClF/SzEmYZ0Tz717hh1j+5Aki3GKoxATFMrE5F+Dr/5YyPEJkL3yiOI5HeL2+
n+STnVEDkfpnCSVnZI5WNQOGNf/CB2MusQcZIxr7skv9t5Rowvv/3ROneyISrXCn
Wuaef3/P7GhjznCyF1vLIvqkr8cqMup/gVXWQDoQvTc0Sgdc5LrmyQAqZ61OeFzv
mS63iZ6OuDkiK6ajfZ5AQTvLqajZhmpLjYd8zVOShz7XHY944u/V6n2VKnmTV33G
ycx2H5pAWkjH90aUDI+NfPwx1U8I3aOUrfP+kuZaF1zuDbP+mFnJfs92zXqz6fid
pp8gNe/PIwJLnA4E7G3xAuVfFgvfKF2SMG5iHoHmWxxntJMy/q2t1FS1RkYMG7We
z7V/Tw1JFJFAva9GvdUMTXWqDbLz8YihCPZVJI/AslDkjGAq2aPQLRGC6LS++Jnk
Jd9dP3qvw/fWmF1rKI8iSubUEHzyqByy3dSknaZdC+N8sAlzMQQ+BmX6Z6GBTXZQ
hjNpW8EvB3GD+S1Xv9a+6JnrMtzXTqDJGtL/h+7d4we9uRlyeOuDa3SIGKon+A9v
GSXpg3oVDr1t+8wDjBMa9qj9D6R/EwgwyV6lhO6Pa34r7Procxo1blwa7GmUs9zY
O4dfU9DWvorAMAXZOyPwzoqoWxceox5JeKj/t4c+VpHmibCSgAwVDADxstR6HW4j
Lw9mZwe/QLd1Tbdte3kjY5iBcHwl3XaXK+sasAQa1pGvkTJ+JuTjmH43qAJo/oGc
wZuYaBqqellXte/Cf+Bm1WoRDvXuVf/RTyRbYYecyESQ2RASyQDRaKXwnI1DjzFw
83XVWTuwoF00vpyrDSuih7h1AdfjMa3EgNHIr1+c+7A07yThb+KY88WArIQLsTo3
pnTqX7TjB/gldn7PqE7rlNzBUhw2G9KYTaFYFj53oLezT2zIFuF1Xb9TYjf1mwkl
46+b1CNa6/jagPAVUjcemrQqJSp2GVTqIkzi8wt+mtHwaecpEev3j4IPbJSrmpAs
tpsr53zWEhNhOsw9Y3UIzw1Q+PwpveIkjfxqoi020DR+F9HvblW+7FW3WugpJ67P
3874W/RwvZaWz48d2ENhlq8tMB9eqMG7uhYxPz9WSZnPBSI0Qk0W0PKXH5Y6uCdn
OLmb3D0oUNHCPZzPvP9arl8DckKMY+EOpTvonm86pgxfyrBZgjXvQKBy796qDKFW
4Z6sqV4TuufBh2dypB+fiJDPaoNDT6eSENB+vnx96NnjfzFaHrOe5bUvXEa6PbID
rLeGVTukNobjJoJuzx1SRPGTq0gkGNsS0pWDnNlIM1hd8hhlKxO490W3FYEnXqaf
3/AOGsLexa2RijMBqfF7t4AkY5v7mB+SHAPwPaEnn5N5WlUZwJXidtlAzD4qukyo
ZchR08x9NsIKHvCMdTluk44669W7f6hBw+RhHlo79UobIPCDkZlkEcwWEt8ycoK2
8N4z4NbTS9oB0BaNo0PWQkdmRO+T/zmsXX8wrgSehyg6E9E2V7ChdWralQzpOO9I
zebfUqOI+hTqhDk7iULfPa5G+ozXLNrBIxg8KzTPo8xv47CquLFWbCimh8ENDcfs
990IzrZeoxLO1xDVhYjj+lEM6KII5F4k/TBdl4Aw67CGLCdQNmVpvDCReEOOMFQn
dYjjWkNU7L6jGndy/w2KCQsTEImD2YsGV27Oa3+3NLg8Q6NrZ8wCO/GZfbTGdfyO
bbddGOvpCakk2zd5mMUwprWdkqxvbCKrnySWLhH1/d1r7WC0zzgml4Vn0DDBFnro
UEgCOObBZG61Bv6zYj+J+++K6D1d6IOtJr4mNro4DPtTLHQm3wfoTOm9ria+8Jr7
OrmKGkCq/Y1rBp7AipKMYcY1bOEer1XeD8UgjfxuAtW2jqcbylr/7dd+dzsnSOb7
w4tCrKiYj5jWyMKfGuFFv4xlvqjYKROPFY70xO6XP4Ge+0Dq2EqWiQJ20zKZbdZg
EWdDuLdF3hzPfAXVcygBU8Ano2pscIpypIBrWpdondNKV6BVjgYIsfHpm7SoOeEl
tDnjntA3E1rpYW0Hp6EKj6ncu502+VH2hA2I3DXUrzuyfbybdoeKLMZQwGc3f7Iq
VOdRsnBMNc9mdq5c85fxOKvcBpwW94g7yTvrYqcWEsOkbyO/zQjFwXsS3F98CFIo
YiS+EcDEOar36ltK9DsJQ8tj/2Yk+fdxREvicdfMUspI+C2SpcASo9zPxPrRvaFe
cWULZjDmH5+IrnnNaNSdpL5szr+a2DrOIQIavtKCvxyhKbVYuu0rrPDptLhX1ec4
E3ypQ+EV/nZwJSWPjUeNxg/7XfUt+otOTG3Xu9JYu79oi2NyZP+Jo4aJhxgCbumC
bCOqaI9HhJMXMGWq4MlfhvM1JO+d9m/SrJvs4SmRjiHDj1aUSTE++4Pkdc4h1o58
NVXNhfuPGEacf6UQqBPOFbmhsLAHvxNj5SRZHqmZ2YWVCNo8RpzCdiDT1TW1C1jo
cChJs/hg+lR6bl0v5PCMEyiBQ7IXWO4QtkfCUsLF9dVtJxQ8KeM1ij+faH71lkcJ
eXnA5w87eIrcHIqzWatdOMi4B7zf4ySSpiHFp1HNUNNE1gF9tguNJ8nPhFe94IHg
T+y1zDA87c4h5muUeKsrWiFlv6grTofpDw1Bbstk2EpYBQm/9g+pg/1zeVTarZXu
+cTALGgkn9VgY0x+jwe8xrSNtDHHVbCIB2e6jaxzmnzMxf+gZYn5HQkw6RuAA7bD
gy9r5+GYFC80eiMV9lEGtn+5HYZpEhYTUsrDVov+gPl5AgqsycPlyFezIsBokkbi
CPg2VasnVZclfX3shu+MjVwYmnFIUcIbNcUxRUqeXKbl1dFK5GN3V+syVVmlVSyH
ATRF+Y0DLPxtZs+KOZEGzmAWMYov4mcYsend1vDN8XoaGlsMqRezrfRcJIGuyiim
NgZ179E5waud+wfqg8iPsjAyQFoVy2mmxJy6UlPRtdTcd2KRDn8AoKXG3yWknwSK
vZsx9Vhtbmb4wAYO+aJ3tpruYuU2wxC8OGwt32fU9mSO/NhlTP8Bb+7ndp25elu2
EI5wCB11p8tEVYJo11DaCq6+1jJAcBQ7VcnOd16/PRZOPspR7po+5IgEpLREs/lV
56iDAJ+iTyQO/EY1ShjabqtlcV+QwcoanqEARUzd4u+s9aLGdJ2u0WeBh8tCYnLE
YaKH/Ti1vU/X76tetFH+6IskAQ5ZhcVphrdaVQw/d6VFruH+KT8dApR+Q6i2IDoC
QA6mzqcGfN/bjJIsZTk45ZXF/G2aQUsOzTWZ4TmD1Z4uTPKcb/Y52t0hZ6EhGnMJ
oS5mvWMiDuT104B3X9yftOtb4/ARjtPZAvw/XhHYD0DW4FnjJ6N77yA1iit8OFmP
x2AcgXsou+qeKWr2JIeqnwcZJ3UOjO/Vud8UrxqzeYktcpWfTlnOC94mhDw9UvVo
YuxCs5igdJnRMu9jFcDr2dQgIMAEH2Pg4uB7zoyaBDBKR7+SsAAka0Q+9YtFA93/
a6qKiIotara55PSlsEvzH047e52u5DmIgVlBjUxr6GWaJaJ99q4UIjI2GyD6IfTF
lR3rFHZ8R9JFhsXuOmXtND6Lts9a3r7kDg6v8KqiwStWnt1WZh4QCSZJJ7UDiAOf
5fduPdYoFJtm7JLs48an030ix9HHWu4dPvqO25EhOSq5li8F5bYniHRu9Wlw++Y0
WEdHRv+LD9P7F3cM6Exn19V2wty4MUOgBHfLPIqqoe6s9xAHHi5D4i9TcGMPLSEa
4MBcLue7MKw2UAgNN7ugmh+vTlfX8AOBruqVbumGQzsvdeCgDJXfZx0Kite+UnEP
uRl8Fe6vt1Ay8XbAPndytD/uhrfUg3dPDR45uup0sis6kTA15atyTaZKe1uoIrDa
RaMuuPUXSaSZRhtu8EaHeRbUDGnivtCz3nDwybmz093BAZ6O69iolNfOAszv8T3U
H51A44qiaLKtZwtrswcmxDWDQBMnGzzLyYv3FN1b64uCIq/ZtMx8DMG3TbfZYs4J
YVg9iphNNuTXOYFD2aZ2/wkFUUbS7NJSeMkpKUDQrdDB7aRiGQgEmg5862+fYTvE
LS4v8dMZcfwlUGvXwhiptoacHIq+wRRVogVRocz3FW5nvgaeKj1bDEIPY1S1Vir8
9uAVs32d5CdA0LGkxNxDo5xtpEUzwrriJGE/GDb5oJzXwJKNtvucKJ/FfPW/T542
BRYWs3rYlrasTDVEAolWuWMjcm1tLSavIayZkepUlwyl8OkhibaMmlYii17aNhIB
OPYYRw8WrnGHbW1OSpEp4RxUFMktUOAFKcZ4CadJ9poap6ocv9bMR0JuGikqHmXj
gKmLELWkLvyuZX49fMnGRnl5DmWTBcU6nICaWwu50owv2m75XQw4LSbffrUNLS2j
gYxHEo7x0Yi73l/nobVDWld+ESygxOxk45XmMAdhkeYzVYhWCHRNKPKshoXTGJPM
CocNjH4HeaAxAQrr0DIjdF6APKlcDuBt1bfiMPIoggSThodgbpBh93SzSrRp8eAt
YpyGSdbFfR/mfhOY62YWK82WvGvp+mhTNh+VFYFYPrs8pEaySV3x/ukQ27+P/fUD
5tOKRqqqaaUXq/8YMhlpKrbdQCNbSrLhxeK/gM7v/zBBaApiF0QaEAu8bs6bAMn8
tdqnHZZA9i+XIJ0HM0Gop06gt9OFAJdjGNWHSoJqIaiTJnS65FRfZ5D3IIhLvSn4
ow0q3jChbBBCg+OdgX7n5lbdVWJfO+zxsdagvnZPyVAvHhW1fefLo1I7yISxMRvN
HsOSnm8l9b6PJNu0I8hvRXymKxQkGBEpc8B9OvEigZguPd9gSlUStZw4Ofu9IlCl
jBuFMzRK4S1OcS9tFX7PX3BE/Am/sXeN2JK9sBHdkQ3nBvMLRktv+y5BXoIKv73k
9mrOXcWh/NJ4Dp2/70JhV6bNYwiAIjTfpxAFdSu1ygmtsJVn3WzXDaCfvg/grgun
PGEWmhTOavggiwc3TKF8VQplyK/b9jgfzgcG95REDtSlvC/W04b7blp4wQJNsMMs
Y/VPiIfytMyjxU4EG0uloBR5fqtRcXjD2kvTMLGY+UIemKpKVYvb2GQAiQEPyWjG
wdkvr0CFTuSvwUh4ljCLu4cSWa9KhpL2MivSgzxUqU4hI+N0U+Z+Wp8l41c1T4/0
YjKAQ3zgFkR9IPxf75EmUyTEK8KGxLZCyJi0Lfmdt/SWloe0EGLHMss2VXBOGrnC
85lYix1cz9n8T94bfI1m37Z0qR9wsng76pLeKEtnu0KRJ7r8SUbDf806kXmo5Hxx
x4WMPPm9oM5iQH5OgjdkkCjmoHZMKIRTJBRW3Pna1BMb/DVEfIGvM965OplCaGT7
dvgilZ1kKu6j0mQo45XnGsLaTYM4brdOeX8QhPcqH0LCgvMpMrvyZZh4vsI218nx
uM0W4GvbAq1yQuClXTiHFDqD9y0EsmCKnGRvHOFEM7JxiNd2kv29Zwo6b9xfan2Y
`pragma protect end_protected
