// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:35:33 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
nzgKmNpZsIcoBbkNw9vwqZblevBxuYHzqz9IkIs/3sRMUxL25gKLaQmjF47pNr+F
bq5BzAFo6ab+yEZVatT/XOipkpO9f1yPTN+PHi128aQtoRQJ6xglNJE1niOH41NN
7CAuZljvx7b66+tY6TVkkWO3C/LJvwlMNxlU19z1foo=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 2656)
M+cWzck1jDDwAasv0uRx+R/XQ1Ogf1mRsWuoucSozo+NVlR0t3A0XppC3x2iYwks
XOGPij9lCkiOtkh1eI0lMWFLbFOk1dmQj8T0O08h82HU86ICjqRUiHogssH7UJ2p
YPR2CXh4uiZtGxcRQrQ5NF3ktd6An7DOd/jC+vmAa4IgKetNIlWMPlKLmEeTrZxY
CouXuRvQoFcbzuB5gsuNVx38NNMP4LINaoltVh1oVUDoCjiVZ6QA/WSe9FkKEp9I
2b6Ao0L9wiwfwpuaWeT0rhCVqk2X+pk+GaXF64dxkkU8nwEtnM5k4TJA1y5IqGe1
gRwiFtyJoC7rNFBt+rRAzs5Z3DkTDxBXYtHI1EhVeoNozVncCnCpD+bDRAHrKLF1
rYnw9vmdjuazVHypDeklEPd63WzQQP6EbOUMOvgIT9c7IfhAC6vtGJ4m3YhzVdlq
aimlAh2k6h76gp9KP/YBcH7X0Kr7rqiwV5wVvZ011z/a2hsZMC4Hr2XN3k3dKesc
s7haBK5MlH/tTh359w0JyhfVs+c9yDVEFuyX1eEifzJYilywc5PQr8jvs7LTf1o2
UYTBSEBmICNA6aa0Vrex6sBy4G8JRdf3Th+bmI7Yi3AR4qOi0ZNqcv8G42II3Aq3
GM1FpEnF2Edv3V5FMwGiufhkpkvj9HnJzvyZpsRUCY99cebxmDqb+xEoWVfs8xkz
na2b3XC+8ZBpnNJ1Gm8EtYsj+WE3DE8lAcdQ6jOFu3hDXRsvlsLfE7GWPMhkJpln
X57bSw/MIOo8E1Tur/9vhCVhtEo4fyetmEAkEijtCElcDLTM1nxzg7tCwDbcGkxg
YGaMDKA28EvV1cKG+h83slQmiTP4DhnxLDyQHXqT2pf0QLKHBu8Xz4g6QSmyijbw
PndSdhWPMhkaZUCZLJF8xW7c4B2Q6Wx0AnljyIx4xZkKe0eD8ybt6N3IHXET1rU/
RhaQSPqByDv4wDhC4+TCOjpoZkCBL/E4CzSyqIv9sWm10D+s1OXX/inzhAGmU4Rm
/qK9faxVVvw2Fjzfy0fdrjRYh9OsfZqb5D1Kh6pOx7vSxqPhofEwDV4gc0Vv4nnZ
i8IyC7lfCvK0oc5E3dnNdhDY1+xyiFr/nHfJxOnXMzMv4tpi098CG+JqNLBtsUCs
2KGPgar4S0okc51cAAwitLB9obono3PFA6nueNGLM7N59+gW9edi4OxVz1HNAddx
9fZ2ARP2KJJRRmOM2YXkxQWr1QbGGztRPL7sHzKwhlzY8hrA9UrDEj/q6/pm9K2f
64NlGXymxCHbHMpwnz5cyx7n09Y4xHmcDgAw9dAqwu1Rm6qf9twUu3IGoLbegtTt
8bHjZ/SIGH6tyABpQs02LcYE93vY9A1cEJXXCTgpIn5qj26NeZYuAPiM1QkR64jy
+Z/bMemJTTe92y//99drZFjmPELneB2upWkXMPoRrd7ewI5POOXsMv4sL3xEJfk/
FEiDHkESOlSvRBKZvLEds+JBNIggvvJxotoTTzR4Z9j1Z+5i1xhs4OKa/awMm1YA
kdOQxqxpTYqjM6D9h7AIwnQF3v7/D/JLY+d0i6l3w1uXXJq6ZMyy9XhX1c5kOYBd
7FX1Es/7wsRu9Shb54uJHR1A3xD2OVS0YLxceIYnMM6q8Zhf3s1pTJnJRv4Fa9TR
oJpFzdJbGxl6GWoSZJFpMubg345VvEeyH5UKLEoWCzz4C+YoyjtKFJN+vrXRjXvI
EivAusnTaa/P0gOoRY4i8n1jdhCqqfzRZRJhw4EEF7TMdPqQanjsBot+ZwKc/XNg
jMpZ4a6tXS/OR5LINoeVQSU14idqRB5WmY8XovIe6lAHSl5C0dW/CqrSu912PGnQ
Qkfy67FdFm5lgEV2f3WKbBZ0pGeiHaMMYxGobi7+/hLQFPOIUisuwa+tSqHk+nqw
IefvyjTDhf9hEdnc017fixQSQm4ZRui29jTr1kBmgXN8KMum6buBxb1qzRrTaLHv
g8xv609ox2dKHlYxadAEqcBqT9FYLTV3YXEjU7WozCvH+5JYY3p3uiKwVgtVTTMX
Soo5juhm01MMbB2W7zY/2YY47/y+9XQfCosvtcjXmwwbA/3IBjIs7471qh8RpcnH
DoxkLg4US49g2ZYlQN0U+Hm0VpHMl/sk1VmW8pWmx1RHpXcD5lw5PFWPAKHDonRW
11Ylp5yWYKJxMiTVHKjgRz7+vcptvru5If5rOO3s+26s4bysmqjIOp/B1p9s9EoP
JLHH1utC7JouvvTAO3zYui7M8QZ2IRQLvkKnbkvxqv9Oi8gTg+No/aer7+ZTPqkb
IWx4xU0DY/BHT9ltje5+GG/kQZMT+2eeui5hy4JZSy0miKztPMzIc1rP3Qf+EGTQ
yC+t6rUwLlPiDX68Po6DAcXdR/Cw7+M7vnRjVghw8MA75h5vMmn4tSO43z13phb4
x6FMKOv9WVGzlGKaMn4ITO7LtdB7tvxvefpYoKypiX+BJ9d6lcIDsysrHbL/wwh8
6sIfpm9JIcGMb+p8IlMyaegnte98BlfMXOatyN9sg0cBdRKhr3h7NJRclJk502Yg
p2bah/mxvTMatkNRwZH3YMvgcobD98nIFXfCiXrl6xCh2Q5JKdrOZlKIku9V2Byl
ZbtvrPXi9uvlmiTI0WrtBgkgPqE3haK0Ijx8WpXZOIXkxbMzhX+ZpmL64Sjv5MzP
d8ZQZIPvgUEU3sZLjBZbLGZPinVq1Iw3Gq9S94LKhDs1vie/PwCzmOwaUTEaaiSo
1fFP4U/UVTqZbZE1ffYhcHYJ3YpLsQPfwH5v6bmmVmI27Qi+2VIHjbnHC97Fq8jO
VBt1FhkDX9HZC+zVZF9GP8HzDsR3Fo+SkqA/WwZFKiPRrFquT+wgSud+m9LnQDNX
DEZZebuyBt5H06ez/Rn71wpeItboXRhsIhzSTyluxRBxAF5Mvi6FxQxsv9eZiq2M
hd2gVIs/m0UlfPzVEAev2fiNf38BranInc1KKCv389NbN70O2GNJ1nfiaURS2g+V
V+8NPRjGuD7SOj5DdHZ0zzuM5mSWLzB7HvB2GDbJaW9Dr+DEgSH9FQOJMgTmjt6R
4RzsZ9fNYKr8laYUo6sLLuSdoECA4jVhACeh5v8pGBYzrgolyrY8mp+lqnYHBDWG
z3RjIzgjYR8wOyCKPrPW6xaeFOCJVluUdeXI0hRge7wLanxTX0U/anPqE5QojE9O
EJJnJh51TkCz4ZUTaPlz3wRQyWmCoWF6OJKu42T2QmzkzOVPQ7sam4dZ9SvqSlmM
c78TTExg9A7TowNWFSV/XR4rEV2iWMAC9wSWMb+LVUTJEqK4yOhKERUd/lvR3jgT
LPk50fV1DTeykUWxcrCm1Xu4qK+Ocn2hHhJ06RPg6NpmAxEVpvJn0Paz0+oDDLoa
H/OjBcMZRqcmhn/hZLCLES8UPTxmZxUnIR4DJhaOwPCLCjhbSwWlcJdqYsG3KCBM
7m/O3RGQJEEwLZS4S7FUILsR52+sRqUANhO53KlqE9eOgqw44N8U6HceQu0ZVBUN
w8TZWGr/RfEPQ+ndD4wQPw==
`pragma protect end_protected
