// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:34:00 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Ara3kciqIyAf+lVSTqSCR2wHw285fq/aNpWqVu0OBLpHXU3nZK5LmAiotxBChhqe
dTl2aYI0ZoLakf0DzenaOgfoeS2SPWd6nmDYrLp3N+bm5yO57+fo70UTtVuU03m+
qPcSNX+5o/Vmb9OXpOhyGmS48uXdsc2136optIjMgRU=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 34224)
d/2s0AFtSK8JR/CjsxJlsaY4ST5GOSbhQwNjRKayLG1csW/RF07y4ndv5X9hvd3i
PzbAoO0IyKZG+9h/p60Le7BK4xOVAWBMpeZbzRZx8+XUTYuS1tMkF+VN6FamX53k
IRmdleIasq6VcIXN3r5d2U/0b09wdIrivkZupc23PWKHa+2bIDIQnGKKQVAwpDCT
uV7Gi3sQSfp0fAFptTnn6H3p5Vp8rNHMrW79W2yWvlfahR2+71z1r1KOOnHcuIIW
eufY+IpUfPms5dSqkWG30oMbpW9tKpeyBowfQLXrHdw9k01bXnAeYq8aDfQEdLtY
s+yrlJxPchkkPyMZ5XHWAQQu5R8H99bhsyHTf3PmGIZ///fYIZwjY9c76LW5nPPT
AVRGh/uczRo/xPka7h6XKDOab6DXfBuM1dsg+RL4bkA0naH/VXopJwLoxb85mpti
5BUgN7gBqLfEUDk0+v+yvWLxlmKQYPSuL1ah4gK4QGNju6wYIa2U7DmEdY8aUbQM
/HYDchn6n65RuKtrC7J4IbCOnWVw9QBgp4pKp64+ssDbNAeC4vUq1bdwMtBJR1oz
1kzRJIkPAayI3CYnmW6BMoZlrRGYPv+9DNDENcpGW8mvTvEmCgOuNs/WZgRvGQsr
fSQg2ss2UfeXgvfAQt6Xc9PQ/Z4vspFhoXd2FNCi1xbrnHtjhb9byOWs2V/zy8ki
mXK6BeyJOhYimDFb6pEdozzMrvrrh9Q2JgNaHEjGH0nuFO/Lcq4aCkHrC72AI2IK
BlCEbXWIeqsVO6G8kiwZNNTDgP5EWRdAabBD70F4Sxv/l3/XplhF4jJItJLw7US8
N+P1xnTWQCQ+LxzZ2GofHYb6qhZ1wH22itz9lB8yUmshgt0gHhtrKYEsIno5yPeh
ma+6Aca7RWY6V2CKzhhXJqx1EkWaMnQ08pCNlm6+4fasz6SueHaXR3fxN03rTXjx
0gLCH7JpoMZQBiD3fhnhdANmavfNe8mlpkoz2b90KXK7EiC59nKc66/wFTABmobn
x+7grOq0n48bavb+IytBMkbIgo+hSLFIXa6gKKO7d1yMtVrDULzuDoUDIjxbiKcu
ztmxDOU9JVHXhzzuxqznGi8xTlU0yFIt4atSUQYBl0tWgtFdnszLWpfDmeLHGP+k
uNTY9XDn4tMEz/5XS5XegL9r3IPngSV7TBf0ajkpEVylYNaBS51jvP1Iyit2OjfT
uvsmysfeiL+zpMe6tCH0Ru1b94EBHeLqmmQ/e8KTwIH4Z8TcHBnmyzXHC7KeG4Gj
HZC+ZKOim5K5C7Tg5IhABkhtRQDxX+d51/zOFZ7NqHLUI0j7Fmi6BXSvshRr0xAC
zeJKjoDlxd/s6yHAMJBtdO0AsMjERJp4Y4CKQ1ykPbrtvnou885Ep/AVVCOxVd5T
4BQZZjXNxoUtVVYHigdrG5rPdD58Cgl+LdsrR99xM9zpq+oxGc8KMTsmA9zuv4rO
qBZcH3ZTyTEchlpdS0OjZxJWjLNPTuiGR0seV03oEiL7KwxIr5YFaJ+X+ZqGcEgL
Jt5wmoZD5UE3cLXAOt5bXklaGVPLcAqI1jet80i6yck01yQj8otF293CXgKNOzwP
dMfjUNs/Ee5UQMVT4BAKjHGkhaA+IYjBwsjzPclvPp/0rkAPLeFLQOduJA9iipOh
+f5XC9DOV/vyx2ePFlyS2qpVkCA+60dXFoFGdK1elBhSxZU8HCmanwk14FlXyKED
MVY65lkKEAWBC3nLIxj6WljEq90MJTamgxM5sYKOIDjjNFEDU2xm4oV8irBdN8V8
RalBtwHA99uyKafMHlHpm4sOIZqVp9jm3Hgao8X5HjaWb/gUUUmXlnydA6A+ay4K
z5oLDY6OE7aMakKkc2+AbrJqVvRaOnGR4ZRrieo+45j7sJrITuuiMZ8XhKs7aCfN
brWFSW9MMXOU7q3GBoVoZdY5qdO0acZsMioM177oseTLn8WWcc1N+kUn4dWk7rHt
qQNT+kkqMGBIAldNntZSo6F+vkOio+1BjdsPNQqbBrI+RLmXFH7ro4XfygWROTxZ
32I63gocQe9kS2J4dQ/CS2U8QpuQ3le57QAm0mypg2UffTKrGyeqpJGMGZ6Neeop
aPAESixJv8+p8xcpsqCZ3x0hfA3QAPHZbCfAiwzcto77Mz6sDuoeWCBu1ULjcOJ+
L6jgdrtsKH2GaVhIUJvUyKu9YFbQusV6by3+kd994Q9BuW531ZoAyjCDJXFsE8YW
twWqPrZzyZ8Hc22TThO4DVAKaso0TpVHoRMAyPt5JDnLMdFlURy15ZTTTA96GRvW
3OmOjgAFBPyZOu4eDIuZ0U3DobJpr5rr0oeaxjfaqO18rfeAbksfUUxiYltkLpL5
m7wKMTR+9/S+LFZQAVPsbhwASX5fAsu9vsYA2lINnmoaiu/FxbpPBzo+FCexLrKa
rzjNACftKSO/pD0I421iwgyvIRAjywLNLNxJXY5p8LNytJ5hVka/hKF9i0jN+U/Z
K19/P0SUI/HeL0xvT++4p3+Ter7e9d0F/wfw4OYoC13iiKSmHp3REzhpWnc7lNN0
NYFbHdagiguWU/9ehy6UjH0E0DhT+uGPHEZCdGtkQZXDKQ+74eSWFC7QpThbxqD6
z4a1mFuQGqlmRQy4p4zkC+SPI4WYknwmrl/HKrQvyf6/C2myXPOMTr3hPC1Ld3BF
zV6F0X1XwwHptr5ZOE24lHwoNmaMPgS6vfVPPQs02dmo5C45wK+omGEx3XYouUGa
oqAQ/KL3jBiil0ytHn+PJ5yOVa98vFnqOwgIjRH4WFaKysKkf7siUyrC3xZAsKu2
nnQx0+4cdSkalEpf/U0S0lAotcaswmqllp3oAienm6IdJRtLs4PF42tNy6AcR+mK
Zy1KaSxfE+C2+b/neapD+x7DGTgOaknuEcozZJBBD7lyfb5wwbZEFDe5waFntWuc
/7lrlewdFt1wHvfeOax2I7eGctavIZxEieGUp8p7pRPrTnpXC3cCZgPS3/HC2Rqg
rh3LTb8dTSHTpKD9C6nkP9rLoqaYet8aIurYKOiZ7JLb9CPZk7xD8Nglegr55vtc
ewCAY7PUo+9Ff0vBdvIxFaZqxmPimjI214fa8PQWU046O3IFD2y4BK+L4TboKSdW
BB64tqXb1yqBAb5K4FkpDzVgPv0X5c7eaRdybOQYVzRONUsecgWaEuvnyIT86G8m
qFQocRDb+DLGOAziehzqTYjzdvz38i+tm8wzSgJ4KniPRDJvmXNPPHNeB8Bv7sBT
41LvxsRMUjtWClX1E8SbvEf5u8PkUKVN1j+ElnwuEXiJD6y2GHM5eULE3IOMCJD0
Llj9L7TzR9V5k0I7hJtGbVHAQs0nQoPCI7sEZ9r2HdnygDvicxVIOyJl5oA35R06
sUF6AWNEdzPJqdGw9A5bXPu4UOUtt17gwBMPwPZHXfYhokrT2ocD6gyMB335lXqP
zmb8BFdlM9o/T9iBeTtdTfnkqmGgufDjF5LlMm5Cp6QSrecorwRPe9KHLvi5Dc7l
lxjKVGoRasJcIb3TuB0+p+hUP7Q6v3x1a9NVSltSPnuAGfd4fdQCtIFcPfKAlYE+
t+sd7xRsgfvoO1HhJNzI0q9quera5Wj9PjT0EUTHUK/h3xmSbOxfm1GZqqi3UA+h
wN5BZvPS7sauJxnOch0bLg7XRpMh7iLihTEx1dD4mT948avnao6dnVi0hr4jS6V2
91in/s0QSd9wQg+pt40n28raZc9CPTxzWqm2pIjVMpmjcsAlqmJdwMCg+ailWdvI
ryDbbDArC8wwq/J91XMqEDvKSJSGC9MnepCREymWMZxSlzAsukuFMCDL5I0OvJKs
F43TOFAxdnUxlraqc7dJGTTJPRfRBT56cSEiQTdqOP0pRmCkCVBFtDjtNFHulaPc
1C643BpQHdQlfqfbGQ1VJjxpL4aiRKQCSAvmkrbln7b7kMo2yTXrAPcUR2an0UpU
U6Y/e5noPuNVWJF4qyXS/pJko1cCt7njvixWsjMcYf5yu4+9StXPITz1SKXWV32f
xvXW3d2cSTucC7wE06I0bCZXxXz3ApggmYNtgnUUeJck0D2QC4Ki2cDq54NvTQFS
VnmEA1dwqCa0VjlaQCgYFfFhZ2XwbYo0ipT75s6i10UI0OswecR5GUZG8hg0MrL6
yJtUQHooyMCkcDhWvur6bqZ1IzD9KwBaMeZWik/Rs5GcNJkjuPc9E0b6grzVpDUI
QZe3EHr7MfubDIGZYBOD3rt0wGTzFnORFMLQR2EHnln7YL/Vyz72TFFB9wCih2qG
DOuun2/gUl9mIXssfIAzkAP2Tc0LBk7JI6gKFnx9U8NsowuPUb6e4gg/EMXsPg3u
eeM0wShVrCJ4TEDU8+BWgflDLnqQXRhvlfgxKzT5+qgaN1OXDBdG0SH6sJnHqahY
qX6Og6/Fqg2NLbd46v0JLUlNjBMTZbqugLOAXwT53ppcMg+6QVC9wq9/s+7mWYbo
8j8u1bLRIlSj1YRHElecj2usNPrWtY5g8TUSr+qTeAC4RSaP49FS+4MniP4+A+T7
ApyllV1nYfCiiXteREGB2XB030LW1GldtJPSRhy4Ncg0Z7vKLnEjDYxpN3864A/T
vAOR9Lpnec5w46rZMAl0Mb0Ns1+SNirAxrFJ+yF44TNqt5l4ZSWF6YYuV1h1GGjq
ZpBivBU6sBDcCCKpv5BJbwW4MjSV4eC3xy0v7LmcNpTwKv2SEDQQIIoUXhg33SX2
g7b4Dg14U2mW/UzI3iXEARLM6WJkUpGnzmQJBK0n7x0zzz+2MYOtJGyQpHyKQuXJ
6zJu/ZUcAFOYIFeMwELxRUUYS5JQmC5BekTsvrBmqUbZHfZWMSvB7xPm831Ca2cM
SwsbeVBwY7PKvEHwjVsq4pN/PJTwjxI6QxO+PXNGmVPGpusKXJCfb4yjh8l1YEmc
20n7E9py8h5NZ6Fi9fJq4VHTI+umH6fBltJrAiJJPh1NKQUwEqjSfeyVHnKLcHgH
7iZwRwD878Kkz7M2X7fcpswSiNFpRt3IH+j+ilQPo9RNDxOLznIhgIsvfiGZFka6
GWc5Jkrk8sUtni/s+ilY+DjGWaxtoJpFe3qRqfKzrM78O8v09Mb2RrDDchGwdJMs
TjEmWLwYFdXTND+hl/VH5gZuR8ckcAGqbwWwWtiXhVzAO+hHCxYwxKg9Gwb2Rj6i
ybSrIqUWGLj1bn9pDfTqqlvfynuBfindmis5D7b90GYt7tWpdD7EYGUELsoLDLxL
kWr1fKgFL/zjRjMD2tdyXXLG4efpD3emmKgsfXoSkVBsi/JSgDx8hngQidnM3XFK
OShZeoffSiSY1L1ZZ7If9bgTq2cUXdjI2dX3rA/Vis0uMiTuMl9wg4+r0JtY+9xF
qDvSqsiJ9qnKWbKCfOGGiro1p9X2l2sJYEnRL7tQtMkGxKMkfcWieL8Oj+A8Y0XK
a2H6OlRTbSHjsQZhWD03NY+WpDLopieskA0tjxsU4BFwLUZ5Y4myAyohHFlm7MEM
b62xaJ0s5R4i9GKgfG34EwwwXc6TpO3M27XtxSUvJAnG2OeLH876rmgqtgokhpcT
+PTNEbXfFLqjAf7rsH0PLlsuyj6GkuNyd+YcSalDA7arnNvsysMR+rk7LCDJcyUN
Qb+sc+v5feGwUQu1JhNzKu2GeDx59e7GUkQUGkGOHRpuZ1xzXwROcXrBK5DdZCf9
ysI07ah+uBC8JOV4/osxIg6UM9YQqt3/ErxVsJnYSRrdG613HN0IXJoJPrTjGLUb
LEQ3wFRuuh9q9A7RZDUvPG37FNhfRnvL0jQYzdGOsV6O8Go24bhu36/VNgOVtkyN
ZDg69Mt+/Ffkor2e4KRUzO5/6iIp+dmRpsi93etUIhiTFQvS9N99ItFKbiH4i+sh
x3MoH4xEWyk5TEj2ka9mOD7ajE4RB5t3Z73DRqEVyN6rRuXoAF6QZUC5xnZQe+7G
rBlQZIdHoKKUMQ2jHiPQfkFhjA9BB+g8diWXTFvYcpXKrvpnlVWhEaUlJOx8Yqej
PD6WCh+BmWzOe8rfDRL/0G7DdV5UZQcwWdWy4pGFVJjNnc9LOd3ljvEcWLCZGrg8
AUCaBqBmLc3I0CSDamUKX4Eror1Becl/LoPZr6j7mOidfNCcMLBLgwOyjqEg1em4
rDOGhrpU+ra2r5GDUG7Lcbta2UHHd7gFEIuoW24XLbAN5H1HQsIovzysAmApu4kd
33yxItyNmDkzlGpM0EfnwkRrboelyrpOkXUj+tyzK21rmYfBIf02VVkWzj+gp/mj
anzJH4Lx5ubstcf+9wAKceXYKWecQKr6zVPWD34he9Ylobjk84RRCoW9XvCoqsBZ
T5FiRwNlRCkENZ16AL6wbuE9SRVM98yW7SfXKbV8qZh9f+Gl/9JXe4cHx0UYdkTU
JOs7aUitVZXbiAFtWA5NKfkPYbbiSglerxisrWjoijxBodzm3YS1CMiSjZckbZlC
sRmc340b/+gALv+4ytXYaDUlzOoA1sOh9US+OqWz5lLPQjy3ysXCC4If/RQej1py
KZAiT0E5pJ5RE/uWWjE99FsRi1oa6l0sA3o3pzFWRjDC/lKQ5d4OpUivL5w5WGHB
zMjY72EZNNIU8f6O903Xai2Oz222HqsndIB85HGwX7qswb/7E8z6eEYnR/Ob/VtX
kEOsiqpw7byLn9Aj/7m+lpRmHhBGfEk2dSpHcPQr4f13gTMNsVZ8hnCi/3boVykZ
r/u35OMr8vim8AxvL6GJI9WNXQObiNWi1x+MrMz4DDwbm4dBeYeV/cK83wFxNpLI
TQ4brI0OuqOgKdehhrRGL1aT4F3+zxMaU1CjmyppAoN3gkI6KyWxTE4CmK3dxqJw
i43mflVNzCdXMtBLyEkyLcMwZ26z1MaGSsie4pvsHzadhkHfOmL8Vd3fwebZHHop
M30E1I/7L8DDhiCRax16VQZkdPzYfsDwu8nq2LXSp2fJ+Wx5/63rrNHVilXFQzwB
0nBGK1UqwYzT32SZ3H2dZrksuVsOwl4oosy5esNU/7jEtrMOoum6FYZqRoqfmEZe
fNRkxCWtpv2xWJFb2JTFMWC+8s6ssUiky6R8fjZZuMY3Ta3s9MF/RUcNvoWeGd3t
9If6dKPdUUa2ia8dzInMQOubS1jjn7HbzN+AmVShYvP85P1pCrzHwo8hiXzFPjs3
qUaqFEisJrLHmULk1EsjrbH5EXbY+QJAvk0W5x/F2neYFH2Gtf0qN7tyAD3ejZyV
HCLK6UgH3yGqRADL8K6iPQd3m5DL8W0kkPCocna9cO7eWwOFwThbl751X48T/Dqp
moOvHjRUKrKfJOaULzCqldn2Aj8mi4BQ5PxI8IYNNSd/oyy/xaUWps99aRXR37Ig
rRO7H1wY2iclYgFN6q98O5kyYMC5AMaQVd0RXrEbOvgbjKa65+K7RdV2qRnaVrrv
+xb5MX/BXOyqyvJ3aXNBD+R3vxghChzkvhfxudQsLbjyNzfdaHx0TC9mHmgCanax
GTBTLis9Dgpl4wWWt8xtdo6VA7bN5yCT8deERIDpLdwtDOhoOa+iemeOdn0Qw/3t
ipLpCDity+k/nVhZVuQP951W33yEiGr/+E9HEfElaKOMvqL0SLFXslrCuBZlr+Uy
RnnLCf5UMreJ75xXO8wYMbm2jlNeg3ysZ4ygR23WRBmgg+wy87q5EBuaHdPnOXhv
vu7K1Dp+Xn95zesD1Ml0odWAnUjgxCmnWw9W2QBuV/42pjrIkrwKkLKAcCebtbEc
ocLyRz0fhRRipr45f4dUToFVk+Gf2k1SAd3ToHdosFLWceJHwxH0e33JgabpwfNp
XsRVOGa1c0tT8qyK0SUDPBy9U/Nag40US6erD+8fE8qHvkC5UiUiQhAYogr/i/5c
EH6p8akFsN7x4G7WBgDd4qGN3EgjYLoiyF+hKly8iBVe3ufclhfe55coLDlyTniK
e0UvDf8aESkpU8BdvVFOIUJoe4MHjBSa6CTUM46i/U/J7fUcQxyCKZzoaqEKjvaN
BqdANSCC0x7Asx2ug6t2AxIbkcjHDZkc0EZ4CxlnhksghtdUjN2qx7n5TN+1iswu
FiIiKHbqFHersTPH9StiTW0s/YXRFWcjKAnj3inZDVuiB28Gn48b4vlZ+su6PtFq
kGNIAPa/kK0TpK4pZDGXybRPowN8sdo7yAEwdSdg0ep0Sujl3DWZbm+nojntikTS
DPYjfOwbaMfYjHmx+wK34DOdWpc+/6xjd/+OE51xJfwpSSuOL0fZRFehvp/HRzaf
dVx7oN+4VDRej3khJnFtadSk1LxYAjM5q07/1vc2O8eIly7uOR0gC0xdxrTo45EX
2JpONkrtJqe0CD6VbgtY7uy5oPzi9dtPdRkc+uqA0oaaK6QLhDaYRrObMxiMkuh7
y2L7y0O81KSofiT4NhEMW5Cr/GWRZROvf5MK+y9AHxQRlEDZhL5i5W0Gj3QWFpOI
13V8N7OWnv3enEozJ8l0E+d3y9s+bxPY4/l+SN1lcak7bCpuWD/0kd6l1K99Oro/
FVB+xZ3jvSF2GujlHmYjEA83KADuuT6xaB5nwGhpdHO8gqKUD81j2+7HiyInptez
qyEpdhoCJysjkD7K673jdmDAq33xrLBN86jhshobWlOeErWO4TY31bG3eeckf9MZ
FsHDmIOe2CP+KPoWo/6cQzWlivxN0Vp7O78v/28Ikkj0gnYe1cozu0iAQTrSpWkj
AwrIQYFIlcZ3epRUrjBIaU2sK9zmrgLKpouqzhE6owu94kWJgF+R/dZaYaUMKmmh
70mOXWQoDtlTjXWgZZ6/UMYVebxh5dFPXr7CD1IFOpKNWTPHYolGQyHHs/rCMO2w
hK7xMaNlIzjKflE+i4CM05jUiS+JU6EqdaSVSSbBBiWRVINLC9sZ5K2t7rqFPSxy
zDBhgmgsb49l6F6i9lNhA+gNwo/5290/ipUIjWRF5m1RT30YukC+7A/Rg+Kk0her
YPEo9nYrFHr/U0O33sfsNW66S4PrbLrogIs/lq50tldHygfDGh0eV8dlAPCbxBJZ
TeHYlWeTnnqxSJN6+suir15QcELJsHz124vHE0wWeYlmVUuuj8olAWrMHTFknS5k
KFMXuEz5DLydcf/5JKj4UdMGR5xAJlpRtLetSXXIUoO1tu2DcD7x0xc56HWFUOK1
4PcmLMor92rloXLncFB+dyzNfpvd0uNwhD7bokTug6r/4Z1qfJ3Hf2pJPtNOuI5R
3Horn3YFVlmjBFLyQIJo+GrCw1RWMfRAPqVmVV52QNiez1JVpSV3g1DAVYar3BrF
nffTNr5eDnph14BvOn1i+APd5LnMFJEJ1iQw3KewR2j7ca+Yc+6F4Xdet45livEf
c3MyPo66qdRB8C1Auit9dEES13Pew/RsVfIi0YVVxu17zuH824aF9CagKBNT2X7l
Nb//zbNm2Cs3pOnkqlSIzLIM9Gem3NoxEYNLuQ6pJpR80Jji2Me9YUcpAHJw/5mS
+Op6ND37CS/1Ca/ArImadEUQCzBpTG4EwnZMusSRtPD89s9bRW9muIGrtvC+Fy6w
8NE3FqcttwJmu4JeI0HYB70LEWurnvG4HFXrU3gOlLTYnABdWRgYjpoVdWImbZFy
CpHPqJn5raIaMQOvwmhX3TFa6FF4SfMXDp8+zGJN6O10cDtnUfsuhYv2tb/hwkY6
N/eTWrkWTEOG0qnrEI/lGLiJTrldIwFLxqryppC2jM5VKaWvJVDQPyHOmC4RYy9b
/DVBYD3QXImk16Rp9GGv6mwioInyuWU7sFKqfzmGAz4FEuphzcXF9ilPRTqz+OTV
1sLLfI8ikKDVxwgBNviOtrS/3iPzXAraZVN/M27tDri1l3dPcBUr2wjGz59XohdY
ntI8AKSgIuVUhI0Q4WiwFLMHgJX4cOIXhmplOWNqKEFgHfG3cnNY4jaa02is0h75
otPB5RMTRI6OpgWQ8b5vOweIqEG7HiCXnfMGa+awZ7prp+tOQ3nidgtL769bpabh
Lo1CeaoVKqdrq/z3gv2AbRCLDavOfUpr0zSJ1TWbvkPzUg0obiG34LaOinXXWX9w
w/RllWSFSpAnKtBLQX4ouQrK8qAbkuDRzV9s0rwju3ZmWosXXGsL/TEko9GdtBF3
ejaQB8iMi9dYZ7/fLScNGpwTOdA6Irh5q3r9dJ+1496CXvkvwuzWTtW3TZO3uaAg
tQP1mb2z+XbGoEElugMAP+TFmDTxtvoNSPHDMnqt/87EnZ+nwzUWtBVxaw3X9rXX
6b/evBCLvPr9yr1GrVBjr84qh3/nNtUO9VWjv7UFLtyoCTnHL0xmE8oJ2wVCgu6s
47OOaVShWM7ZNYE8dmfSggJcYIRemvcq9i4plN/HlUlZQgt0ezFZGFax3fB0Zogv
FWt91IHCJ5iLFuj9RyRRhNJw47kK7i6fZPytAKnt2SB2HtI8mZg+G5CcGZSePrwb
/clFwdL99V9yN6Au6/L3sdqbthMT1+JheDNEsnob6hUf62tpMpG23UyetjFPcDLS
7SyQwHDV7RntSXDmPMyLSF8dPlRjf4phyBqnhqiXcxAdHqiITmigPvRVELJEQ7lY
ZKVSMrkdh4thkehUWVMefrcFJdUvgfZSRIZfF5dODY0wO/2XsFiwX9yi8Go1Euj3
pWRj8B7kxl5znMUzhNn0PqQGF4z/w53nxwQarIeCF3UgaGk/kqoCJy4ZyrgqjSM3
34GfE4IFMURsK0+5htbMK3aPh/OXdysT9VOXZvLfekHfo/BjFiJHDSYfHTX3Gw+1
I3lhEPvTFWeYg+IWC2LiupYHwgPdds49xHUyYsc9+d0359auxvQLTASKHnGKRUlq
C5yqBDZXcui0tbhstA4lf/sXCnYpFLYHzv7cf1mq0LC6kGJnKGb2X9zWSKgpAzw0
qOaC4mNRCf0yrvSp7uC0bft1K0ph46LMflK4hOVxWpkeFSjhxBtI1u+ljOpCfGpw
0zKG63MypbNW371Iot/+lx2+FTi0CeShMZqQZHbFGXp5rvRG4RaLv3hRXAis2hjr
aMVuPJEHJALIIR+1prlH/ZJ9Ik5BPM6YLfdyuJCL5unZzHWCZ+owxWT/3HpdIoDJ
NkUvtpikeasRf0nq93by7Ue13KuUZPe9saMV7E9+qygwsypBEJY//fSbZme+kOFm
uOa/yjGpWwjy4JJb87eYiTrSIZ2yWzl/bqBQ+dtRE3n8HNf3XeJTgFAiuWtVB+uc
Z5VUZOltJVnRqMK8iWL7syJKuvUVXy0oNlvIDR6enz617gj/RikRx0CB7prQ4iNF
o4NfE+ZDFKkAU1uEcJCO3hBNlu9ruXy6MkdLLWUjMRqRxi3FzYk7V6Td+JbMgozq
enPt3M7Z6MBEWdd4AbAF4/0IMQp3IKOWiqLYEyAfWmi0xlHLuWZczEW1jfrKJyo6
5QfuTLRT5vNa2eNp7aHRWc7pBKNs+TOHWvhop4daAliRApZ/e2KZiZqm1VdWE4eA
R8zmF4Dh2fnVi7da04gK6kkS+1lkKefhYHGy1kwr0SpnXU7q6JlzdxhbXwU742JW
CRpG+sHXpNqxDZXSRDeEWYYOIvAfNEc8DarxwtoV+Bn8NbJokCtZZRaJhXxgBrMG
fp7iArClCU3WMzmgduMiSR5PQfTfqTAjleeRO0lBqg9wWqryWcTya4qy/zR22h1I
kfCY4SB3XIo6irLfUh9Aih2T4PSkGFYvV1JS/+xOMF61a+5a7DNQsuKC/fr7WbKV
RhcoyoxstS54PtDFlL85ZGqY4a978Mjq5a6cVuI6/ZH0tuoTGdwCm8U+cDK+vTIa
/5ZgRc3V2eQFv+RMA/uNp99CBq0FyaCMC+Dl3TGI1+6i0KxLN55Gr2LtXSOaWYJE
o8Giv8GeJqf4WV2e/bCT273bxJvpPPi36T0bNCVOyXnRjJ84X4PGbNjL8SjWsoSc
1jjNLihI/NPMFeIe4aPUI0y8UuVDF5J24yC+2ALrpgg2B8AGBMCCKqP6/d7sJFt9
FijwpjO52rQWYKxpK2qpwgQnndRlwAXr5HTzJsFdX5eKpTKfbxDuQ7s1VroExU5O
yhTlfC1bCBjhmmPtoYtp9qO1r4YuG52ynjgcS5dS3rM6wxhBPOBy606xD7vfB+PO
ksiZ8CxHlfJT7w6FSS8XGM+stmeyiB0Dz9BPVQ8YmmzfOPqoOvFtJ5Xi5DOUgF08
4QgY/rm3kv2jpU2DKoCl0oP75LlckQBHHwslXvo5cXilRHEfUV3G9X7VB3AqHFNb
MhEUZzY2kxTpRzOGFvG1rZhw76fdNV56HEGeVLT1n7U9SicuTHWFs1+zmE9Rzt7z
/30oEvlgo8GAOGpvcGdcRUwGtNfdMlm0PugTndWqVwKxr1L5if0gI/Pbxgqk/Utn
LuB1cl9Ce4aICFnZ5tdJpuhKb8nwXXZh5PB91ZcC8TdjBN8p920Cm8YSol4GxwNH
sBZ37tZ6w6/kZ9A15WVpxHlfceT6A5FGCO7+++ODozUN3gZPcdb0mb2+pa4AoLrU
GqcZcj3MkbXsOqlQoz2ha70d9mY2qBt+09MVz9ErIdAK6yn7BmekYNJbhY+SIESg
h/TUUvEgSt0mC0PDFwt0huUM3Ou39Td/PfRYWUyAE8TKrEDk2ghEFKvV7VKQAPGs
Mm9xbG8DQtSNdSPdl0iA01ckEmNnjDWZUalnJiD0aKYII2ImaryCqDIVA8LNWZ7O
tR59GQgGttlXpdrR6mGolYNgMOahvcK9tS7zQ4jAeUGyJuEXIV5LLXF7JsrWjc88
x7Tww5xNnA77QBkSDjMqbLWD1LCrIWsVp7Iajx/YFAIQZmQuvRiuH82QAeF4bXAE
ocwIx9sS2gBrw73IfhPj9Xhv6Qo+ZAIE409T5NCaYyQE8HU+r+qCVXTCe0PhEQbW
cT/T/VPIvWh9lro8KtuP2/X1fco01jTIFlQ72TjGi7h5yrwSIlZeF7xvTJxBQONd
0w4nwCCChGks4n8HE2oF93c88EHd0BTgSoJqv5ZSSyltLkeVThpg6PC/ZedStkvw
HyhFUydW5p/ArjU47IJL+WZt3HJ3BTYa+bVdzq6cyNaCrCWw0L8xym008R30qbKt
QA1m5fkwfnLyp/5Tboc4XU1YMtA/1QHbtKg/b5CYMWqFi+xBaeoA6BiTR+UieuIL
fJ86iFkm2/xplH7LpmNUVCyZddHKP+CxbqMOxJ9jjnOTYXYd3maPMFr9up9dzept
6UnxTccMqXhO5Kd9o/gS6XCCHjL+ScLo5+ofqpaAj1uTTQ8WOynfSWe8ROgdupMK
Tr0Pb3k0tEQo60254Wbfy5DQxUSRkh01jaXE2uXlEPxEExCDnQWxnrr8qVJybwVH
CZ+T1DNyJXaHoSAiiBRNC887kmU3f7WGNBOd2zEjqEk99KuQNcn3FEAEhP0d5S5J
kxxjzhyKs97DwXjVGWezkJuD2dJ146fIdZ1k8MiJLqFj2Lczdsh4jIr6jbLEV8dy
/Gq5uHGL492MpF1m0KG6rS2wpdqpX4gPAgj5ydY0xcMCZ8aDgxBiml71aoPHEkhw
9wfLaZwBldy/OfnjCR76AFtgmgor+4SVa4Em7Pd049e7nVh8+k4G2z8EnSyEL/Sd
3UET4xctBsmDD5vpRc5yC5y4z1gvZv8l2xcFGsKWdo6CAYG8d/34ZYjxkcOPUPEs
FybP4edSJmq0h6MSlowJePJKzRZ5AFCnHpPihhwzonaVIRqPpazCwz0KY/Q59KwF
CDuw/2UUd3fdkt7sBKamh7pWZOuUN8ikWr8f1gprXT/2ujAwJTQ/t4vODh26UeKN
smXJ/Nq+CWZX5xyVdRwPT08/+P3ZF/Q3rAZ/gxsrBNRKlpKmWOhmHqZSBFEb7YBp
9cRf0/avBlGg+jKva1n60WNMK7TltI3ciWlcZyINoAsigkuxn3gAQvr0VBjQ5/fw
5C1tKiuoEoM5XNz4DMCIFZWigl97UtVmKKASMSdaxavLrl+0VsY/O0cTRxcLJWMP
3R9uskTT3lSvV6z8ZGnh/RgPW4sZzlvfHaFhWChUU5oZrcaicHgEnimnlItbbGZ1
dYLwkyW0FXTBdc8LTcOkY7wzMQqcbcghhZamv5FqIZnwPvz9AhEPw1jcLxY44eg5
OzkZoI8QvwBFBftXAHZS5km2zTSDIPQKpN687f8+kb66WKhwudlXngrWYz6pp8yt
xvpfQfA1Xb0FNvt4Cy3HxA/UO6Ru/ec0i44p34M2padmkSckgcadINBlrTDde1aA
FiU+BVAD1kRdHKJKcExHfuetEQavUrCFAkaR6vrfkiBYY7zc3s7k9MzvD14hXOsj
1STLZ9z8tkEzhN1WhIAJb6Gd02XfkEVOtotqJgk7EyItb7klO99hT6BH3v+zMkKS
wHG2dhzp5trgkG+Bf9WSlUnq9v5aR20PpyK4u5MHN3G0J/MnHzPuJiYQk+bGQgt7
0Ty30SeR7UPG5b+WSLmbarq0HQNWYWJcJuWTqyOGCYRD8uU+S6RmbsIoBSDUl/gY
Ww/sZbgoTc2/zI/7RA7L1JhOm/Y50+XakFOZk8hIxy+wKrCJixDObf18FQWPGE6S
8/gHGV8v5yhf6KVUQvfCy4ir8+uhDHvBW6qhzJtcbgTYyXQZXEcUJVY/Q7FKX7U6
7t6ZhsiOBSXLyXrgBhJ2cb2yTEJMi5aDWZltiJYBHpjXyTjasvdJ63N+i5vHKeGW
S8AHFigP6stLL5yFLLHKoOEUdodjQgSWVSQlV6zIPlfDh0tA4jw4XA4dyc0/JCPP
AY5IBUoJyb3jO3cxs3p48vqvUjN6Zhcv7WN4i98c6xzbYm4jkJUZLscHULIVzTzR
iglo+gTe3SD5+p/qWCDvXTfUE1IE1mkH+GJJzz7NoU0TGF4X3WI5VJ7qrO/NjoXD
kFl20dwlCS+wtceNcWMRjMd7MdJ9pQJ0DozcXl4PMN01OjbKnyXmioJ9LH48orXl
i3bhD1FFI/DtqY16uD2rbgrDo1mFCodxgF4I73p4HYjowttUdMeUHY9PE6jg2MBc
o/eD81idUBGK7L4Rim1EJjOtp/Cql3eObrnQ5fEdOF3vq+Vle/pHEVkS0dvw5bc6
weKejBYK8z03rQUaJogQ5ho1RHMhyEn/9gK0M2ul1ElUIuRMJrooDS6kZpy0C+Bu
VapbyLqu3Eo5UzLQ5ydBMTOC7q5ey+X8dDYEYQoFKL98iGGCIW7VIDTcP8izfSHl
IOM6XdC6alLZcTj1SFiw43tWXqMiZWdg44OB37iWaQx915/dKVM3GYSK47fVPXTC
Qg6jb5RPHEEQig1MUgDsJQ7Sj0g2xsXLc5Sgcv7yyVugDy7y3jMnPnlIZSuOskyS
qh/A0ihBfLLL5HBHBPoIrToDatjWfOgaZKnSAhVVxp0ZeVgFe1pCcDi/CPY9cWjK
oTq4CvuV6nsoEZXQ50AMvZyTvEV/Syz47DmGdEUqKf73MKwv41uhcfPIi+TxY2ra
Kx58INsQsZdJe7zwTlhtj35BY7t18XQBmCunGm0QKHi1XSCodirwRCWjlh2uD8r1
2HvR/c93DMnUxOH50ACFajEeBqe70yFzqb99RHWaxHi1aG1UNRGw0iV9V62jh6Sq
j/o4XUsIXLFtygqV8fj0TDdUxQMJhFM5FM7r7gPdyia3XTE0HZD4ez/uZF5Da8sh
ir1N+Bl12QVSDeBLvx0OMN3g6QcQVaXX/+vWAzOlcwhvXyX8BlQ+zNDWgd8avyaU
FJTXso2xYPNuW1uX33Za+ywTTy/3etEFOBTm28TAwVUsffS+9+tQZDOgMzKpzdYb
E1fpmw0pCRzINgOV8uUgFG6cehGEyzAyjTWpwLFj9ge5qsS+YN7e9cvVxCUvNR5d
quf0iAlDYCj37NSK4aVQz5H7fXjIuvAAcX/cG9vbvwY4TgNg3pVBJe9WOJIwOor3
4f99axUoToR3D45mEllvyPJm9ETWjZw05HZujUIf8B59gM+1VayPnYnxK6tMhxNZ
uQtpbC0qScdV0st7Ud4FbmBfwWnX8yAOhkte93RgeV24ORfcn1vNWOj/sd1t/pMY
d7XpvlCW/Vr+RxwUWsLNYD1Mu3dVxuoFzkNLrEj8gvExqDECSHpn48N/n1jY67qV
a1/9U//nITr5FKiiGwtXNkHac6PUB+n+Y+YfVAdrV9nNuBca677u5z+ufadRMtN0
BIqOas+dSHu9ZfEZPT0pGdxkFrG2Rn7dLZjjvFAboBXXzlKgLDj2qQxTkZyNnx9T
9Yaokh7NebhXu1Ik8tt/5CeFzqXPuUIvvNtUxIToRw9tLe6bDCqCQwRyYEV5Kqp6
c1gzqsShm+zuM8KxspvXAMlsdqr8xyquptStJWZQIYEjPPHVlC9pNzb/Q5zoZf7P
MdZPod+6nAADxfk/3Kj9VVn/9Jc2M2K/W9m3Vs2kYsxo6weq42ANLPWHp26mcF6l
uxcdCzmlL9zl6JL+YnkqYU9m0aw2R/1iA4dGNAiJcLGWxjRMHNn7GTh0lc2yXD5Q
mQMsTpvGPnq3KxazqlmjlmqE0VPIkAO2RqdPaHvsOx2zwz6URmv/BAw2qUaZcpZh
/HQDbT1Lpcgkrze6vi0Z2IeyzoFlXLvFAfSg2ZSuWT098U1OsAGqC/tgfs5vNArl
goFcXMaTebgkr7FrDcZRIz1uROsQJqG5erPe/4heEMMJcRdyQf8PUAO3wVP64/NJ
wZCg9VzJp2UHwcBbo/BzX5AT0buEzzStDBMUhcZXJhZ9S7qVZwIgLJDDM4GSbzoG
4RDHwE+mMi2PHKKOQq7f4m+LmF7TjQWu3gcXFltT/cEHnxtQe+ZOKX+PM5/okuXh
1cNb13OqWdTmv6KFU5lPxBYfNN6ovaschfEPhd6CbPf+tYvxEGpZXi0oPVKKldkd
yjhGZ0RCtswfxsInwCRRlbFnUlvw4de9A2TY7Y6dtGKBgs6Bq4eMP2xpKTzHL7mD
iT6VXfqcKAia/V0RlSDZ9DJjrzQ2ZHGC59z4nnwgQOS8xqvpbWIbe7bZcriZqnbn
RUBhT4insWziGNxZpixvYgXzt5LdkigTYrSNl325HlJGCr2jPj51cjDp46eyh5lv
YIIcjOj3qfy4LEz+tH22wVmfM7E5WnX1Ctq7FuaSTi6/r45hFj3Kw7syfRErblJl
B0YuBrn0Or6Co6rkaOgz10+oDzjD2SluJU+SA7dhA5xkuxnu99JEq3X9D0mO0rh0
QJLaj6Wm+m83LqlZNqgB5z/9dF8xTEQmUoDW8I/M0U8eWrml52YxtA6Syh5sVmXC
ah4DC/yFo/j+s0vjckmuKmW4NBnVdsrS9nBWHlaWWw8/tovf5KIE3SwH3fFIgw8l
lskyLCQkZpnw3/wBKoKPyMUmE3/Oy4PHjyXP4gJ1Lzyw4aJ+VJhj2rq1Wynowicx
Udp+rnaSxxlacIjQlyzGgsSP9sAWt5P8Dvj4z7Y1VprErEsVELlDh4R7DuJM/ez+
nGmlwPz3BFLmzKz4FyI+X57yr5LMSqLQmkE05EIxiayrSQB7F8Ur0DARFbLmMD4g
08kedPfCrpKJOoiFet4oHZenr7f2Okgci5HeLh7UlCXbEgodQLTRGQVM2p0ySZJQ
V02dOkboi62EDUuyz1JCMvLe2ubH+G6RNUsq9q9mVaNwWc0fnKO/QbG7qNJl9Bsf
pUWffWTyLb5/x7zoBd07yyAqnaqCnx9DbMPra17DPLAIsMvNqbf4enuzZa2njfGB
O5Ftv68zEtL5i6Y1N8sYMU2omGHRLAVcUnyh7WNIoo36m4luZvtCrXunKanBMWXn
RPccM0+9ywK8Gvs+xGCCKzyKpmdsZ2q7VPCLo54Vw/unCRr9RGiLmU+9J6viZ1jS
agEQm6JcFHyZTOMKbvENbCotyCPg7caxJVh9CXxyZdZP1Xm3SH2CKRSJdO3JAYwG
PcAp9jzf8IP9wMy1VbiiWAM/UOm5okKFPrKKvAv70KuiPUG2ARbzkbL4Y5dTG+XQ
1TEs8WbY6LVTVqFvnUA9l+ix4tYAYvxTFBFwVWeiO9W/9PMLAn2DSqRQTMKbbzLq
1I3VIM41y/YFJ4f0m+ILaW7VQ9q4xwai0OyHqjVVpl54wZbLqXcxXnLUjfIKYLax
y3zpNnQvZ1rP4LXdIrMV0cDo3VCSMkWaO9oQolZkGqLaB2BRhw1PA2Oh/YAKD2Nv
RLZZyt6Ra0tAoH8XIarMj/wjv1Vz/gr76DZqJbu4vjg7D2XHcbLbRyYWI6J+RbSe
Fm8NFLu9jW0HsPbTbWTpZsX2uyDNEKqZwi+2jfZIx6l6taInP28T69g7v9KckkC+
lIOpv9VWHrVykn+wunnUU2lZCMlI5aIET1vVQWQ32XlcytxUL/kTUy1ZOPyNOeYz
qKh4prxLdN2cHiLa3HOFqyB54zURryMSqFA1ka9OH+P32+cWPy+9AiyoxqfVU1kP
nl0XVmHiToqo5YipPdM5qHHhfxUX2EmkOhrjBsqpedupb57r0nbWLt7BYoREOneZ
xcKqn9/9J6O3P8nBL+TMpgVEXgXlf0H0FBYYxV1nJ+GWfPVUAOhMMU6Qny0aGd8N
d2VQzqt7zEUx77/0A0WBLv7ETc3Q7fro/ypxGFvbGaQIpdyDQ0dK6f0ISii7u0gv
GstJaA1IAnYUbfmPLReMLSXQWoaHGQZY3aQVoCZxY/0E1nFKseaImu7kcwE2VHQZ
H+8eR3qiiM/4EkqLMpFyjKhr2iV4TFYmCIvjJyJz/FkiW+sVi4oLito+PtRvLjeu
LXwCA557VgZcBo+ush48FONdn+goIZN9qceaUKrCZ5G4XEQgsNmj4kyH4TSd4Q5h
AxlBwuLGmC8Ma2Sw8OqnyqmmoMepk4/Hpb4ydb0LZyZMh9wPqY8+N0gwwOjsSi0f
jvYjwWaB3EgnbfY4RUEkGyZxvCMn43rclVgAxDBSk347EIM1WPlgcR+g8DcgzxXB
rHrjVsfYziyIUea0AMSq5a2SW3eSfw8ceK+D7CzP0IMW10RBQsCmM7DOim+HkYqe
yYVLHxwV3fBc29qBgRi5cQ0y0J402z1oNXUokPoUziboWb0Y0N8vNHgxM8XJw9m8
q412uDMgN5Hk+kSJpYVaVS91bGjl1FjI4tcAQ+C6OVD6NAcwodmorxXcR8H7iRzQ
7zz0yMx0ACBCkRm0roIq/UmHKEDccFpISUXZYrBML/xHhcCVm4/6yq71Opt79B00
sJ1SPjp5D0/UsqAs95WM9SmGSlVW5k5PbNEelKCk6mfLu/N+G9JtwSJ2ksLc/SIQ
hBM1CC9jHjteR+4tkwe2Qz+LeEIUPpybU1i4g4xUVDDCZTZV5Xh55tv18HfsIM0o
tEcizOZsVlQpNvNvn3XBxikiAGmrP7oMHYY8l50MerTearbreauO4GoDhUHX5O/Q
8SjTVmDw18OSNpdkIsqX6xvMtNNYPE/1G5NXLQimkYSLW+3szI6nK3f0Qla3rkD7
DQIPtk0jDcHRc1vIwayiZvhDr/CMjJWyuwtGqX+13E3MLNJs6Fjidq4bvbvcLwBB
YHIdyAAwzgsSZyWIhl5wimnosKjAWRb+FMp3GiAnHX2b7RYp0ro4Uv3Q7nW6W/Mq
YFm7zA7wqmjqqR/2D1yuNm46Yc6OYEI27xQa3KuCzJPQr63W5FCyfEMXl1ew3FSy
xlv3gbFZfjJrO5sNTMsiLqNT7ynXyvWjlIuKTnXP6Okv43cggDcPJNLBN4K6iGs7
fUe/EQ9JTdX4BPppVOhDO/5yMqBtoma7Lqqalemr9OW+K0evYLksG4C1/hnQcgmh
ZKT8ye0cnK1NNL6zwGBKzapj7sKbuWxGzKqTfhA7eTws8sUDlaPSt+Pzi+srd2lZ
cVHP6v/XSjeLAPwrnBthZdAMr8qVa3GxMYpEWnDXAHowIMP84w72znS9UZUU4/nJ
Xc1VBy7nH9p9c7TMgM5VWGdVljaususVXh2STBx2X7H/h+67qzt9Ppeqfjk+s3/h
M9Vt1+lRz8/aWxdjtdhpbea0ndmm7V5dCIussOm1ld6k+j2A4Grqc/55oNYTTpbE
sS9SeDvTGHMs+dEr+3AWsJXr7qtmeZ1aPqgxXiHJRe4W/AfT1H/i2YsFTyXZM6CL
58ESbsCEoySnUwz/LYUW9+lxDd+EO6TCVC+MYd6xef5ObobQAb/5rSAbiSzyXe3f
kBU5h0109DFTyilmxW5wcBoV7vKi3YHzKOQCI4SPVccOaNCxkiNz/ysiGfYTMQ7x
k2LZQ8HHvgPdi4O4tRC37zMkJBUnfUEZR4yzOH6NUfn/PxKjOYE3PNhvlHVK3TH1
nIW9PjpKJGPY989EJawyz4vMpu9abO2DHq3iTmvcN8sL5YLufnBJl3zm4OKXgBKI
j+Dq55tbm9EU8mM3IGogyEa7iustp1Seot9jAAHgefziDLFFMUfCTbotKtxBj1RW
SIh8iBavI5EGfIGlgQLLOuZtfcbq5RpUD2VLIfRfQm6FTzNyCGk6HCcM897TMdol
a6RWAdzmeUYcWRs2P+expnxRBeI9RYtoC6Y4ubkG6njb+e2fvZhvOWvShIfITSOo
mt1bvi6FurCILfZHu2XU9JqgbgtZZbeIN7L7uCM+jsNE2+budxtQOIFe2WZzKEGi
7C2ygFsLTWvSG09wRBUkJRiYxEEFQ4U6WBhqFo/zcXsA+ZwwFUrRbcM5C6tX68hi
kgijbQPl3x93dBIDc2aDrLxcNa6Ut5E+LgIl8sOuzrUWDEZ348hiVmZnZTMDsg6F
7B0e+9wf8EvQAGJkSusFMhEmwXeoKcoyO1UKzxa/GVTNKjhcJc/dEJn3vIHnS8TP
+Ny9dJJSuScHFF6ILdUtaui1kYWTejVE8BT7iSTsO6x+/ZU1akffd0+Jfl2XwloS
jmHV1tklll17/ygkUe9Vv6PtH2rOsMS91apr/qVm19TtGkEE0I2FzhBwzuzxFMJl
LxzrCSau6TgbrVRcGrBB8OTVlv8Ip5/+fJ/i7CTxjPyalQxKj71mG24/EUck6moM
qYCyBMe1AaRtGFR85K2+GaNvf/JB0ZDmC6H7anQTHP1boaR/KrgI0TaH4wkwAv7V
XwYDKLDqE0h6UaDDbIYEompc2ZwLbzWi/rvtGZ6eIcYYnIoJULC8Z9x4iRKuSEVO
/zd1zrg1x0kQdB0cX8teVcWBHofisti3hVoacE4PEisQZPKsrAorxKwd0DsxDyGA
5zTDQz2pdEgpXY/E6CfqX/7Rqiu1iLSmd3ieyfUd04f3pucw/YZ70+AX4f9ucUJH
rZ/9/0/A7XP4mDefYFOtFsEjbpKUorbk76zceeCOwdpeN2WZcZbmBxrgv78dwVQG
xAH7w0t6O9S4UUtl4NiZ9VddkftPQVqD+/Wn33hVTriSYNAK6RzxTSdUWzz9lV+2
ST8GwVBVnzJuGCL0vR5zROr59rymhrtXvgXffqBNeMNQp9pZt0Yo+05BJB1ed+WK
1zHU0J9k7mIvVt4rem/b3US4ml4TjtXeZ/8HlL2Yt4UCg9bXNgpNNqJSg5MBX1V+
Vy+z4b4Lv8FwagCkZCLj8GvG5xOXdAzraLpXpwmGWnGM4EqDQ+XKR7rnt4yZUhrD
9YlVGaWOR0s5W/CSrwZR9qxfsCrpgmRmPesj7LduN0GawFf3AFxZqIMAOyx7FCD3
mZebFRpHG9Z2H/4nRlK7TY4C7mO8v5b/NWjbzTxBdPTB1t1wX8FIbzaoCyioTApL
Cjk/p1bfr/tmSPJr2vvL90AAEv/Hk/j9BCD66/UPi53sCpMfh+kJ0O5mXRN9bJil
XboVwTCR630Yf0UAPRtQJXnFdVtz4EXuVvv9hrIdR9Y5YVAtQR0AKGAlkDZQmUya
e/114o6b7We3cjRNkzjkHZw1gTzt/60dDV6uIYVjxgiVOXNOmm5peG1yBXKO2R5D
/qsHgD2LO8EpsPwwrB8G6d3tgSvvG0pOD7K9FGNmhbKgeySSZR0RXLMaDAuiJaDs
WEJdy3Ycrk+kjwYBeE2hjTW4KFtWdpSebgBwxnvuEa157KEs98EthcO2DtjHhjJN
tWPizwf0vzN18YSe+ZUomAZYXlpPKuTOz0LCO2tHiM2zoqYnhq+QeDNe/9VL8qEk
FZEhV0j5wbCtpvf4JM/YpaWxErDFvjwd9VNyxSHGlUXuSQcBq4zgrO/fbCiff+5D
FKKUF9Ud1hjZNsQpWREWXlA1zuy/dcoaounItWDXVSAmwjfJ8ax0yGaMzYT6GG8j
QmklP9ynwVkAFFg7h70HqD9zO17HdLvsuDu/Xlnhvz/8YrRAJ0SJt0EtiVrUi4xg
dcV+o4bdVh7sC0+KBc57Z2NaPGvqYaJG6dIUrRrdjJ60XUTCZ09jlCjPdKUIF3C1
QQQooiaK2tUEDVlem9NMeWuGEbZUuCJXD/Hw3DA76UUt/VaEOo5soJrHVWapPt2i
GQJtBFsSoqRlWVnAqoPhn9bT2nUj9XWiNQApWAPoI9NpVYvTy/BGDluC4ngBl6RB
Ojoy2zUmYo/a7otFfzWm1pGr7ZJy5uARf2PVGPYwKfjtGCQ1jO/0cF0s3aUKLpjP
LBNj44inpcWWtc4A7EPzDxtYhN7HRR0u3xg3xa9LQ0GhWbvhsCHbQ5h21GVOBMjh
bCK+lpBl9KGr+kpQ1Z63Tslg3JeYT5769srwl5EvzB+5U5bsDEkj1BilKlIAzMH0
08EgxCr0jjEQZOCizPd/YjPbYe95cTL0vWbsHuianZtecpxwIOwaPRl8BpTkDYMv
HzizXpE7tQrYQaP5MUCw7uKuY2qJCBpOQYwgE/fh9antYbDpHU4SCixWXIYJrYYx
h7kGpnW+VGdBQ8EZvjahfcyIdoINe6WaBRbQd2UXHVO19WH9AAM2jau0XArULV87
NKYEO7+B3QhkIZP5cx9s11eG3/Pm8vl3qFOAbL/TWtA4cffK8xZT7M1/B5zxDKhg
Dm+RogyCY9+XoaJwd2BBmGEPlzQyW8mIEAYz4d8Uj3KKerfqjUmlPhzoN4cFrND9
1/OswK+zQiUZalW6iFEhjUpEaZglHoJV4OfDy60wtykZvdWycw+m5aH4LLsutpjD
7dl9l4AAH3g6wGuhYJgQqUUWisdARLq0JW6AxFjOAB9O5krp6NmLqxmTcVEpW0Pq
NGNj7PQADWomEuH/dZVlOHxUt51wgzZVaTf9l30qdvbT8WYGV5QiNRvO5lcnyZLb
0VKqyNSFh3lYMSOe1awUgbMgtDmIr9UfYZWHi2h6j2kg1H2htrc9k/bx3Y3pgnmO
M4R+WZsBAZQ293E+/YJ96yev9+2q7nxSHApE98PZaLDab9FPaOIUzu1h9besx+xM
dWh0ips+EYg6b0H2pMkBQ0kQ0GCtOMUptTJNnbiK5HQMy9ci5CaxIeF5qRQp/J7q
tPLp4zzoLy6c1+wr+Fh2l2wcxLGpbQ6gFxy9UFlL6i5Q4c6zDqv9j3+Y1Jjw4nLW
JsSYwM27UgYUYq1+4oMeDEd2L+SY7SnAG2+RB3BelI1NXn8GbeR989NhWO9k+SLF
ElXblKGKaKg3v5xIQwiNJmRYI5/z5+v3XiDmUXVafVjWxw4eMoQruyZl5K+I45PU
+PLqxPItpntgmPjfa16hZAi/gFInyr09woMsjifW/q39mRnCxnS2TLI2eeUsHUj4
Vvo651MAvhkHFgxoWglLzqPUIqlYbqf5yGf6cBk8KkMk+wfELx2sxxkfIpEbXtaH
iaCsfoYTvkWD24iGX2HWELG4V/7G8x1jQDgQaWDaC5HHrepLv+1MW3sZ0qVUCjQU
x3E8Wyu4soW3z9m6K2JqJr2Fe00ZgMd+WP1pXo+cdOBZ2+WTJBmom5Zf8gQ42XAf
LqAn1o4acbwDgbErNBrU1TSoB5cwAw0PZDATu/ombzE6aXcvWLETU8kgQoCzRRSX
qNXUlY2DHIoL45ZUj0Xec0sECdqqGvimQ+N/4D1sGMjT6BhrDgnVE8o07dbf2GnG
KZki7SBSvLoySf/tmQat7aPzN8l8glDTuz3s2XYUt2WCn7rrInIUogcuzKCwXr8G
f5Tn1PmJNSn2mppaluzRy0mICbbp80iGQQ7najHYNQNrCNkpkrTXiXtMEx+671Ha
R1sZFPiS5WEymlQOOd1/r4eK7+eJsnNH82KVa33NNPW77ibgVBd5RZ88xfckOUQo
/gTD9+d3KdFBgSMX73slYe3pR9uK4h/FhERQKKyUaomznKG1YrCYdsUK+IGW0ezG
KxaJd056/uhczmdMndJ03CAxBJF9MbULwwR8FRqdDGhVNKta0Q7YHyY5VG+8jH6h
AYpug3XLt2y9+odCIc0ieup1LHoyPWBOSVdNrJllbPHw5TugkskieKz62RBzlZ67
coiH/f35xhSNwWPxJACAaoZ45a8yOFYvsHIs4R9aPYDULT4IbwOOpWoYwYEVSGoA
jgAVKQfrQj8O2BAVT8egS26FGs0lacDHXqWpvLY6F+BU4lfsGIfH3X3FKPMjsxQU
t72IA35sLde2QSn1QjmMS0gas8kVlSN4AihA+0fOxkqcHdkwl/GYhj7iDut0+iWs
gNa+LcjtA4kTAsrSaNF3W/8RGKGKhoonreRIEt2S1PWUZFAT3gSrEbRFSS0Fw6MT
wq+js6nHNleYYp0FXVu9RAfWPUp7G/N0SlJhPTAYJQNrvPAy9LGqaL8ShWfjMoWZ
fjcA9kULgzgvBr3LXfWM5krcKuQWUbwKtaL0MEF+hRgd1KGCtKr+ZqGt9oBUgc/p
DribZm1PH/b1kP44YMhwETjmOjPYMrgLSBr45TZ/0LypJ4ZQgWpcFyXLVYEuo16L
0iKJughwNgMAbMzPxblmZpHdu7QKH9QL6FyuVPYkpmIpg8e4F3JAq4qnLrgnD4yP
JjYiOp0q2eAeM3ShMlDN/Uls9SIdeLFKl5vF5Z+lcU95N73VwGUZK5MbI0Ej+bpr
nD34lHyW+AGrPkXDDzJbJplL9pESTkJOSTr878j4t6Owaz56V8AE+liJBwEtlowt
yvuioQW/4acXCkZ+DH+Ycqpi3LH28Vsq+AhhF+iCLBMRg20L2zXC2TgtnngS43uD
gNac1Hu/L6A7++DG0bCbGpdF5MANkmZD57WIAV14vuPPo4rc7eaRu1S838gKPY8c
FDvfPaJ7qV1tAlnu92d0N49WG+ItCDHvMJUmvccWa+wwNKt9+dygDHGUlYPYPv6p
ZRvueTox6VkdJIMkYRYDTfAnKSylj+EQHRJk16zx0jMFU1vduwggUpFAXrIt4pef
NaI6Qzp0Pbg3pBH/tud94JrQXWxLvVRoT2pFYomjKCEUSc9bhXJR1kaUXFEviO8U
0HijSuxe7ZhhNIR5TCI4brrayKN18W+G+b/TEuFqPk/7yHoeKPl/8X7Q46drfc+/
u89GXYpmC82sPu0JjP0Yi0Z1B0s+QfiGdUJQaMVTz8v0Th3hUwBAhT5t9TtpvXSA
jcAgQV3mTxFbALbjB7yGxWJExHUlXDkRm24IgeYMsxhxdocSPLA3MwR94OKOHllF
ppVSpYIGEYJJjxJybLpvOsjlDarQBarB+qfHhBulliJUs9Gz11Ve7EgDi5j2SfBd
sth79SSty5B552nmDYWKozOuU+MFpc5WjQ+LBNeESXfboqnkkfc155WDijAqETK+
PCf2U9igxxK+zMYaQ96ShHcn9xCY+pPArUWiCtbnSTsxNEE0LHYuQrzN0ELtwogK
gY65aSc/AqqjzsOoH1kxZGcOnHVcNZzEzZX1Dz8MQiuUZhCTwoReZQ18hmAJvCF0
qQek4woRn6f5D5saGtuFWlH0BgvUFiBpZu5LNnu9vGZzemwR9Vxhfq3pdV1phlRv
jvDGdst5AftjXNHA5w5+43BIH7ikeP5hk+FPGYTN1eBfZoXmoiKZoKQ5EvA1/KU4
W8nCRmA6pPY8EPRHB5SkPnJyJx49CoXM4X9VqLG2PCByVNjzCiCouNIwX9mKK5I/
+90AsjGBx/ATAaFr00lGc4kJlvjHFxDwp820kn+NIriq63+e8zm3DO0F0WOiy1/X
Uk+oXLyho0VrSXweGR2w2pywBaq3v7BHqXGJku1BGYQ9MyjG1eyPxO1O6zqXX/f0
KWzzkWymXie9joS6JusFq0hKD8dGaIOmUeeHK45uIdiZH5VV0L8E99WYl72YUkbe
mTYizW8l0YEiRs4DBkcbyJ/LbWCX4BApKIuD4tyfyZSxlgejRwFjh6Vxi5hP9l6C
94mMO7TpRDMzr6Bco3iZQBUgus7yt1ukR4Et8HVk2+3rjlFiWX3m8orOT+OcOrRo
Azhfyb5ERvV4SamGEG9v5OzeYn2Pf5hbN1SeJ68f9eam7RMYPhqUaBeGzSFqCsbM
NhF7llGHHpHBorv/RPYQTYA6RPClhiqvqHy0Q0NIrUnNSeffdYQuaUBHr4nMeJHw
oK4txKD+cSnt9aBgBb20/5vuQ4w2dzLneMVadyN+vDfOb/jGopGFIdoDI10xSKrY
A5y3K0+C6O2vmnWa0Yk7ByqDm+/6jxhE6mbKopbxjNWjgTYTxdbO86XrojI19JpN
/i/EMwuRwmyNiqcQNo2e2sQ4BnCVAlknGNgsNrmZhj1YCaJ8TQz8P0khX3BKnvG8
kFptENHKZCOAMGQVDzgnNL2jKAwzz/n+1Cyd667TiZMKXY/dbrm1sfyXCyqyD71L
Vz7vg/qa+3n7F8SDwTi0pQQGVoNXVQDWX63lW25kykvh8TgNPj2DxYrrunQRzKnG
LZRbGYPSJZg/YXmq+CsKaCCGsXBnz9eFwpFJkYmsz+hePv/FcDR/0VhAzvRMR0Mg
BEqtnCKpCxWah5N4nxG/eeAyyz68iGVjPCIVo8XGfAgWKxiDFjrdjfmjCUBXsdWL
I61eMSUoOHwNbLiRgLznA8octioJMMN4grWKrxzDdMdh60hpBWzW2jvLR9Jj2ai/
k1l1UkxpfNppXMd9Dv7JM2wX8SaSl+Vj1Qhu6iKOJQooeTKMMhrWPhxQntESBQMy
FIGxyct6hboh6vYZT1WMi3jzSdYDT5hNy505lCC9b+g/bNoaaSiMoUWvQsaJ6CRt
4RED3PXsaST9lkM1xxrjqQJx47m0P+RkiH3txvYVH6bnLEz3OfN0Y91vWKmgcJKO
Qbw5F2okNnhLu4Y+ezj2KymR6YQUxv91P4TfQokRR76Tgz6rq1bJpfazbmQq3ua+
25OG6RxUpnH3ok7IGt9GtBUf6KYKbuK/F+Co43D+mrELh5Nyy2ZE9knUDJp20TB3
TCK8DQ6HKhiaXPuySlEpU0NJyPUxMEr0d1DEqSSViS6At3cGTF5cxZvx6X9ui79B
1ByZtBdFCl7wik5gx9VE7Lb0S/A9UAVPWpPlA+KDdCSDSCGNQGRzSzhVLvSKL471
lB7+W6i/AomPKrREfFIlXM/63jF3+Q15OSMNzCKM3xfmttvDu056t8h3Eg9PKqIi
+5WjICvt2JbR2gffR4J4J9YPLKuiUkL6FX6n7/3DjIEDZvxCRuv8Tqs6K+LveV9V
obgvXeog6ePvnf3EWCHkg3oAhXDzwY25CjgUD5GkRyTyBq+a7oRW9dF6dxpvgItF
te/GnJt812kH9j6fCynnJtWCpuXCroF4xoatN/TsbYaZegOL42El2cJWBy6YMKK6
kI8VtkOUz6uWPf+sD18ic+fsQwB+lnkrY1xk/iKXdDtQs/3XITtobibwYGbDX5Zh
w6ramlMAlms2nhO0WIdaqQJ5qvlHmMsE4gOPYzaVbnMbcKYChAGee0d3YXcU/hvv
Nx0Dk7zSwZMZ6te7Q3M0WnloUGmCntHe/hgJY3AfOoiwsxeTZ1Q02+sdp2q6G8mv
QClJjlAVnVav7tGgM0U3TLaH2Nk4r1C56KMIPwI1iMHITIrU9BCBI2LNiwLIxWXa
EFAPsVAwO99y+TWIQN449J4NlDPext0yevll1dGtmO79mv8jHg5jT3lj6gtF+qA+
wWy2fxCFUflhCtmhwbynI0nNrkncSXATllPsH5uX73r1f27u4XPXK7LNRu4+q14V
GQ9XHPn+4EMgwBPkJY2NlSqWsUu0/pvUxUfgOeExqjWnyofv4ruODGiF97/sG3hE
neKtN7q4kUOrh499czC3HxpL5jXVjWQWLS2mUtTHF84UPbKE1NcNZG44pdF/wg8v
j1N/P7TQ+awAZ+lvD8SwCwFeBXCro6HvhsP0BL+cuv/NDgsMe9nobtjpNXU2Vigk
Nxri7CAFhigUXBc8Li4ZM7O3Et1XbIWLkMheHIv1m1sFJ4XEYnD20Lhj3+u96vfJ
6HVsHn1KKU0kJNcKM+5ie9oCe667C+DJnRSPt9oUKCHKImv6yGa/2DY/VoVBPScq
bHI28RIuMigfZP3TGP094jWZjRITxd1QlteM2xQlsKvO4/CLnpVAGInDZbkuGsYq
3C/Ew4J9Sq/CIrFThw0CqCsFqp35yR8Z4UKSmxrSrrOE/X9s7402vrSgLxqs+8gi
e+GmatHWdcs+UEyRCTU/pnhkdsN2Lg/+yrF92ID153wrHMS89nCctXfriFZyt5RH
vWV/fA++Or6KWsVJv6yS+uyPNXwOrZGl8FE7MJCessg5eNS8ergvL5X0z8l2A0aL
5Pq/5J1XBXnE+qTCCvHZXKhCGC7L1W/lbNvLbROvqDXyDc6lMWwzkyz2RMHEtq27
HOrD7Nw90uxGSkheWDEYkj9Yy+UZW2rGREZCqfIoYsXJyM4H2O6VMKu6/UrjJFLp
8RifRF7NL9IyeAZHxtQrikgsEVZt+67AZWiMiaUsqfttl2T9MguoPAA2emQVi7R/
CQD0HLYns8GCcIOGBmbOZ3dA2rQlBPnjdvoArkOexN1LVZpCc1QXBweCLogGJncO
gnQ57Kreb9YElU1fnpb3d+C/Gmnm+dqQfEHrxRTGS5NI4SgjllLKLDL55jPmfrHt
5IlgDZKkjw/PmsxzOoHl0l3m6PY62XzUiDXI4ligS2HeT5Um+hkV6tSXugxSctRn
9I9abclqabbLINxvcL6we8MkMeYA2WWfzCV/m0ZPbsYRuytd7pacrdSgM4D+UPgx
90zCRXihAGoCT6daLkSFrf1c2GNFkeXZfMknsGA10T7NNtfERLPkGZaz8qwkuo/4
foQLePSwQzhK3gWBGIkUUuuRbsWTTx9vTVFYgQe7CYSNUEmwOUiq8riEK1PUX1Sk
ieExzrdfRsUeT1lwVShyPuIF82HwNN+eP8x6i7zvqVRhZmQeYU9//oeBR6/kuUOc
32N+cJPYJKIVLrtv3n3cEC2KHruuHOo3ufGnhzstYIw/zfT02KSudU4htNXu7+e+
KhmdK2V2pvOge+HXGvqoYyd2EbrWWRIG32UhfFa4AROYFIvAh6Wj6+1VokBVri/S
dEDTfyPW0vIkbdAul0xZCSVlWksmndDoU+ws1bwamma66WpG9PURPlEFefKuZzZl
CGHpsD/yKR+0wR/KBoOEU5B8uLPRCPyichSP3Q0XKCNxh6I1T3tReJtb3RiZbA6s
+kd1vN66M+o3v91MuCpPVxSnJxfBzBKJR13aDQP7t/CVh27LiM/EkCrQUAKuAmn7
SQPRNafbwSzWN/2+btdf4Tkw3Cd2gsNDPE3tP5Fl2GINwBEIe+NuJxlZvy9H2yX4
/M7a4qVZiYZLEb45WwT+3PI4QJ4dDWeh3N6MeA808lDS4uWE+nz4knVVaCCQqR0B
lM9JpKxO272YwO4QHdNq4ohEUjqMFlzjTByqcXosB0bvvRB/4kPwtzuolvUyBAxR
2L3L5g948A+CHaIkdWkNrbA6DrF91oTjoVm/KVmtFsbFCGgRG12ScQ8vyD90KPmj
+qfY5FImVxLmylJPArC6dSZDW5lw/M5gH96GVQOnmYdh4GLm2IklMwbrHeLygBsn
uYj793XjJMNjhR+gLV8Q59S23Zq3gccx216nufwfN6uzJqXI/uRt5V9oSNBI3K5i
2aMAuC/yw26sSunOsMn9+vTpuOQc4AuBsccEUyVqliVQHrJLh7EhFyCkKm3dVwXL
dzwau4hUS0mIXklQzluFoozPDqlC+CK4vfaTF0UAdCcPULgwD5e2wWRu1VYpQUVj
8gCvbUXuNcQAcQW8+tzCBcihuXMOg3nl5d0Pi+iec9uPnhRNHev85yoTSTkTKZzs
BMMd7DJkGRwLXSmjxVtEKTpJNQcDjro06RQ20S/JIOp2sKpok6N+3jgisPKWxYwz
kzxETipxQCR3j5aCG6SnpdGCG0j4l3BH8eXLEmgrKR481vGAuOxL9qhs09fk1SDv
tlt1u+kcrje4QCeEcjHv3g3XhYcFLLW4m9xukkLDnaBJQm9ghbUWxZpDVeH2Mb/l
3tZToi2UoNOOqPGe3ybLpPy+Cwth5UKn24c3djN0H/xlZKL8D1IRYFJhsdEuNcMf
x4jLaJMiId1d1ldZ6m9aWx5xNbk+KCce53d+NSPCvXAfe024y/gh11zT5RbNU4MK
zXkjimsm8glnffvjHVAcFKlNccV/ebdzfH/jmKkHbIQkFr0QaBo3JeUq+U9ixLe2
Wz9MijxExi1Lnf/JhVw/rTAOE0sRooEmw8sL5VpdajmkTvCs1WQpyle8Wq6rNpu+
NS31fw7Hvj1ykh+gEMIEj6Q4BeK+u5rPj6wpWoyKTJnS7GOBma+TbHt8m7GpK66m
cefn16+CPsdpe+Tw0TKNeH0Xc7AGGWkhtB60u/2Q8ggBOmnv4xhtbE2YhqEE2FCs
eXDT6SI3e4YQnNCtSiWTS0tOWxCKA8LgmZP+fIzDvAbBc0PIvX/HR3YdyWccgm+t
nI5GG9GQydLU5HmWgLuQMLl7HwVfk35jSOzyT4OBiR93QGsU1Bz0LHpZisKSxsjs
czupvUS+HmilX7koAqv1RrPabn555wdDg4tdteBzp9ryXPbQX/1+s/NqnT8XOu1C
IGSsNMsfwAbF7gXUMQtrYyww3A85Esj9iHbJeISWB9uJtpMjZWtaCLQkPa53T0tP
UTAAjrz8hVgzAy5c6XfzIjbWxJ+oYtuBpufInK4ILgO3NfNH2JJa6900VdCK+NYm
X2DHWSNwvd7kRABXGyEl+3dWc9AUZlqkJNIJIlZfnsTBj/NnSug2bx8dpNdx/yjv
krO6xu9/8vnp1o3V24njAPtACDhs1sGnd3TjgR3yDs5xgLCgRqilBtxjFHgUcnVX
KSQ5+if7b36/CY06TyEFM8kFlI6SXv+GbFuRMal/kKydqeVq/ZuTMadD4yRHYlgt
rsEtuP/m99bB7ERer3upA0si0RyD123g8PqtlHuXpso+fNOz+eGZkDuEWonqpm0v
r5JAsuW+oKwU4UaWYD7QnxBs3SUuS8WHWohgWlHkkiDhJuG+1Ov7GaYboRdpkmvT
MmcwjiFp2/zdbbrDWEmUAzK9w2ooAEl/dNGwOwgvXY5jZq0z8HwAedCG/8cYVGlD
e0rgQQMaeOsx8z4T+qKq7tIZ+RibdAWWEiTNmCPpBr6cKEH6kzqk1Sh8qqkWs5ut
U5SuhIVnDH1mnoe8dXdtwen7gOZ9vYfYpYi+HK6gu2lfCsZrmHCiOVmtn4DCON04
H2CQvxOJvyioZHG7YXFkQPlJ90jIkrBrnY5cFZNsiy8X7W0yPOvR3iula5Tv5htw
YJ3CY1ERgcNUs16sMOoYrfB6JIxh+lQDxhKCQCecSec+p3XIAP+LvM46S5gmkJDm
XYlKSVraPmnFARmB3q0nJJZI9F6yjz6oPpU5UIwhOuiMgmqfqVZCyu8czQyJNIJ/
t5RicZESK//ZukRod+bEog775v1BPsfugZoLI03fubsmax8iNm7qglFq7sGftaWU
C6sj7F8pBYKXG7FH0Kk4ihRFrJLW/ZGbzL6R9fpfEtdCO8aeKtXZYHM0uQIopo8o
h0AiA644kllDs1tpb7ggG5bPMoeap5yVsrQouMMcGIZc9yKtCL8CumkFoA6C/ATi
hiA9S6J+fr/N/QR3CHF8qXesNT6x4dNdHvFowWPPK9nr+R/wAFCm122jAVWqwtDL
Uf1ij/jNoq72NQeZfGTlbwxRcLS39XQTWCdI+iVUiKiS38AhB2p/WPPFQ3z2VAki
bFNnCOoFBkKNGA3wJZA7lzYlSQF1sDFj6FezdielQiB7HgVMSIQdcsCbvjnvdXVv
XPD/ANjKlTFm+opGKf7DK9L5OKH1HY58fTRLnMq4VFH0ylHsT4MaE1pTBhjoEDyM
mVcoeSuOSLb2kPaUifZkWDs4FrrMc3EetNxj2xbECycEOxdWLhVbTxS+V53lFXKO
Fa8WF4uZYVpmAgP1uN8C6mDSHaHgNtds7pECzy2S0SAriB9GouvMuYunECm79tXO
Pj6pf1gQX14Iig4SwU/JfA5riZNWVdLudkG7kadpvvOGE7VNjErVXl2JrPKWvQfA
SffVX2l9QxIbqabrrHagc+3ujA6JG6X0kKw2BKT0+52EdcPLTBUCjeGx73HeBTiV
T2LtpJvcqC7VCUVX9DTuj8N17x2hfdhV0qVboHFjnna7GopaLIfmSY2Mtz3vEN6v
lTCJnQCHvVUD6k69zw/mEm1SZGpMn1WQzE0IPC/dzEYDasl7/sV/raTI0+FMwi9M
xHBjsjUoXyRU/m8Cy2u7n8aEaKRhRuQJaVvyH/dz7pgeyeLCH2kl51BcMoNap4TZ
jb0bSJqSpt1FUb/pGPw8mMHW2wwYpxUUOkShZYNkbauKHXL9yNzTwfZ7B1i6z27e
XhF7GMa3aSyv/phbbT+z7Nm19XqUjqyEvPT8pb8mZFRKKnh0rnTe/0BgvQeLaNY3
WC1MaABp0UHch0wGA9BXvy0NNs5q3i4czBk9s8rsczgBzwvHKixNCyl69znprBrO
OX/lSUrpuZSURyfFHV2BU6pildKmXKIZMRozKfXQB0kUxvjCy2V8rEl3fYAWDGR5
9s66DF4wJvpA7OBvYaizp1k4vBR8BLIP3vxfzDPvZHlbU+fc3EwMlhD3mXBFLhsz
73xjjKzX4AkaHiKI/0f83IJC10C1VPlrk0Sg/rKolulKf8UazubfFQ5Ul9N5RomS
3LmKBzGa2/2Y2wuGAq4n+cWttOBT3+YI8boQhv4NmNlJfp9mKubUqKQHevX+XfQS
uY4/gXI1Tn6GkZjar9NlcJWsCPbBogqmar3pboVda7dVyJwHncFkQdC/KJ+0eXHB
FEIaqA5Vatwwn5IULb0cxXxDJWafUtX/pClXO0gLg8mna9tXmVrjyCfQHqKASrE8
0r8pfBBvnJECWeeTj8KPuPAQbCDjmcuI1YLuBpZdb86r0CxGIsgHDddL5UpZ9Tev
AcNtb3bbbbxdxpig7tZcCAlluqoOmx8jV8MVaZN1Aogz7ri+jBlrBroUR0RB6568
ICSt7FDlL5XosKK2FRvzhZ0KJFifpMZZsKHvrf8Z2HhHHzvn5MA+gyagb7JlDTDR
mrxd+FB5FG62w50zJyAimBhKNFcyJ7blsAZOjdq5uKJQkfdRp1u51hdOoLRfE3ob
t7d+izNKJxlZ563DXJMNpBFiWWPHgq1D3GqVXzFunvZqMBSIWwtzfIxCS+sKGRRT
2IUBfJMdXsqdE26ZgWpysT4sIOD45spuPWJr5Kq9HS9NPUUTA1CJHY8ZbUgN8ngI
j8RbkvQeLJY2JiW6G11P0kGN9b8Yfhw0elA4pS+ZkOs3YBUV7NxXKzlqvKPNUU6t
GEaLFZC+BwtZ9H3SsFRkz0b6MTwDjoVOuovja1r4ORc9pCTjxycuK9/3KQeJiecK
mFTI9l9w0KRyClxFCThSXoVF6D/vXrc5Mda+PvJuxyFdNRviCa4OlEtBDWVVdpLO
t8SII6k/kVYNUbnYxCPr9NLCIlW7Vw2MyxNt8Uu45zDnQvcaDY5NUZBiQLy+L02u
Co9fOsHmqVFV1h5wQRFJ9nKHiw51YyufmBkDlkDk5ZeJFxcomuN4wqDqS0IpVfkA
wN8qHLTangYLULNDoRrGuiglASD3EQeUA/u5dDl4zmEqPJc5pVmfpExJbwHEGQ5g
cK7/Rw7ZCpNBMOZ99ICKo1DwCoB9Ish5VX+6SrNA28bNdZHEZVqsWaQ2Clg6KfcJ
lrR+V0W5nSifulFmrilodXOP61l1qsM/qGuyOX8vI5rNLnYN1oLbci2RiMfQ3rjj
eCIBo8ZKFyd6sYpsQfgg6D+LmxiYWnCmjJsbySTj96Fpm2g7rxsSspb0y5F4YQU1
NetPrKN9hOjG6h+uIkX6nKlpaiHzWGUU3p5LE8b60tkSzjhqyIxT+cT8Dc+u5nDk
ZVUjUltmhjTyAFgiN79ThP0zG1QDQeAwYN7SRApn+aHGmgv2R6rajYD/g66Ok1Mp
j0K2PK3s6TWtt0yvK5pk1XNhHdLO+hip1WMXNYlzlXtYha6Lii2Sy73q3aObNPVL
uKktIwYjTGOsXdCPDB+i0f2w0Q5HKNaRCvTvqALuncMU9e/+7L7lP/RhVqNLZCuU
NqwbBZMTMeKMG6HL/KUELoRmNqcTaSBoguRAfypU9rh8jJB0EHgzUaedNptynMhu
rptBlDtGve4Wj0+Z8ZjZKgya3nnFJblSNCELJ+5TESD6qf24nNjyLUd2R645JuWO
YGnVE5GnCO0FNVgsGd3xYd0GwfsxGRgTzL0+w49+dvGH2Y3JFtGBp8degHHCefum
BBD/MxbdUpE2G4QbFeSiJO1g2l4WDgR7Ng4j5LK9hPjvYStV/xu4J3es2YgEJ26S
UJZIpPwlhCqyhIxdLgk4iKNq8x7h0PyKiNDaykmZ//rS594WLc+Pc1Q0Zwu/N8fC
ux+wGO/YMtRSyW5FnHAz5XAFnHnNvOaihCt+8k+W34Zvc47bVsKhHfLUEl2ZrEQC
TqhEiydgW9VxdalRPTDzoAcnT5qoGxhBe9DrYb9tqtPraudHUCTnlfnHwTDUJOPH
0AWIjRt0ZNDasy2ygkPnbROOJBp+7As1TdWgLcoadRo8/lXwknP7ZEnNfPB32cAf
K/Pn46Xd18jIRg+NTqiSWgjmAHw1oCXiwK5CuFCUM8e2+YWN+RZ5Yd+NPXHh0CTl
TYiSIfOEwvxt0GU+lhS7GntmR5f5kdMcwlhPuKr7KyFT/hYNwPNHXvZqYV90w4oK
Ndb//LL2GezX3FRx1wz+QgL4db5JYhbdaZ5bKn4ngYdNNMI4ZXekLSp/BqIRW9du
YKZP/jAjv7A0j8q68+PXxXaNeUnPm8vUMdmY4IielQVcoDqiQNTEgng1IAfABLHs
xxuBtkGxi1Qx2zO8f+6z/ovzU2GwYva6baygaqXqg72n16NDlZ/b8t7/4K2Qp2Hv
F6gJvEU4X6PWsx3J6QNJPQt10AHLGLn18YUzfCtB+ieD5xngnEencRhEyDRwX+Fn
temntXvr+d/Pm627AO3SuX2kb+uBlevjzLHChHgO9ukr9D0a//yWV1YUsBUUmdFA
ILpLg0d8EkGspZFDNRDwJlVrfI/QhXJj/qmJ5bd5mOEZb/wj6qb3GGrSSK3Ba++h
yhuyYn96BhZmhs9b/Lwz8agyhrRgWdRjrxojXuHKh67WWma1EwMv/T9k559Nz05x
OOa6ncpzj6r6unYCoZ3kSyjaiw5WBzb6RtQ2RukhipTye9bvNauHHZd0a2DByM58
xLUloH0f9mWU/UC5sO9q0oqunWAhDgmxfynzIO1DiMn/feHj05KrDHs9DorQA6/9
ssJFf9EzZLXDd9qZeXcpHbuc94zmIcOkp6Dv5KOo2203HpBVPRuhtrA3oTvIJ/m2
WkVI7g7FrRhnzZ0DXMD8OSui3N9L94LEJ7c6YY336WZM0fbbHc9POgcZen63VObH
aLcZGJSpzf9VuZ41q5+NEwLWTT96szYKgj8EO4dfMKYDDj6QoDBCaICwMyM9xAgY
+GoVQNIKl5UUZcir74sNW+oFr2lQslyLAhPs5jK7ypAv6yAbtugIkiYdkBIZASjY
OcOsumsp47qCsgT3hX8LNlIP7LU1azjMbxSE1oLgBEi+tmY01cNbocZzeR1bszwE
KrD44NIX5KZRt7CTmXBQeoAvQqqLXp7klLgU6l3uoQHMjNF3FuwDxgEf9YPYvvAU
pFUh1EXCLKsdYp2pyV6b5IVT4QLfus473jdysLRH5fwdtWTnptYurbzDjeo7A7KG
DK3qJG8EDmsbaFyqQdYHVCICjmTQ4GBUGERg2qb8/Sw3DRFPH5WxGiJN1tEVGFQH
G8CCqCb4uP3yhqxBh6EtnrwkX2CEiG0yVsISyV0zSKcZcsDo5skaPAn5r3WxxeTF
xnCnTk57NGS7Z/E4x6t23xXob+0Z9CiJWigmlvgiXnvg9PNxreTfCrYcCb5XXZGs
jlgvHD4FY2LP7aINUfHlqoKtyI/wWzeaB0QC4sWQQxweZTRQ5HkxDi/06k6wAEmw
uMSs00NVmAWBaa9KbL+y80fUNzjY50UHztfsnrlwcueqq2ehoGBWJlb5zAu67eVU
DMnAlkuhLWgzNyJvHDRwrE/DXjc6ZEZiHip3PZtoo3dNMLDOT3vdHdMv9xhyWMRE
xQ9OQ7yGTv7LG6FPIar+tFiosvCC0J7xqtGeQdmR3ES5sCL5ZsiQ9A6lE8d6QGw4
dEYnQM8M0eUl0AGlYeE89TCVrP3R1GtNbLK5wEeZTyk//nqzQIRqNR+XH/9jrEeB
Fi21pKNqHFguqL3QzgyOVCsAG5cVF9sshYuf+8pHbKTXCXieZrtld46wCpUb7yi8
1nzWQRZfGM78xyD95V4U+oHuuW5K3QGoX2Qfg0e6dLJLqeG5mPpcFanbNaS8KODw
dUM+PoPk758eMmzAB+OAzK0mR6HaN+pECQXX8tNjDuxOHOU1yg3q6Tgr7rcjObOv
o69ifPKvgDSNz/I2K1VD9cYi+IE+a+wItbX80WSkYUNlYk3S6y4ICAsyb4bKHxFq
c9JJ1kZ43EXyo4Z9Yt9/CvpHGw3vj42uH+hBPDtjgxdhr9FoOQkF3QtTAbSCozMw
yEApHRMvLXYC6OxWfrdcBsA8se9DReGehewUKGYjW5cN9fpZfy6V7WFip9T37ROE
eCsxUQ6pbzxXko2qu2YWidJ6OiPbc3oBGRMNuPLwapQt4pIkD4PQLUx7EnpKh9+7
x6nPEmSLlKW5fI1vMVZwc3lBvphlF6r2frSNor5jHNwhbRfVLfcsjobRiv13zLSV
1Jswfx56eKsjCXNTGDNhY+6G0B6HPf/SBTnKgXgZlPb+5mMaeOqqa0M0p0uDxm0B
8mrzXMNEvsOtdiqjcbx4iAGR5b5KLZzwT1lvNb52hpunVY66Qk99Y5xZMhzFpSuw
sJ1xCEV7wvf0qJa5lcZieBYSqRCXVQ9jaV2HZFONO0igQFnGtvsN0Y4CA3Xx9Fns
U8Eahvi42U3U5ExhDKDGr1SEA9OkChStKgbwkc5ng9Hr+HXtHZM6UcsTW/yqxp90
DA6NR0uOENON79H95EJpgv0lQHCTzhKdhx0/hqVeJhD4L2uz4AlKSpU8KgNZY/86
26Ysu8ia+kZ7mioRRpOEmr7avos3KA68lmiA7vPj7UDjb5PWskQ5iTVXAixcfvbP
b9bwnGx3rkierbl9pM/4oIpNICo52CAW4NdVaD1herWl3UxgXyFftqy/Y1AQZJ8L
UKBepSLXE3FnvkD53MIpGyxfI2jQGD5tGIiTFGcYIhmOyAUYEYlMFPBxcs94uCnn
DnaNDpMmAsXkmd+1XWTGcKcAevVp4qTOt+rKfX1hLgSoFWp1yHuPBnap5BcSkpI5
OMKHES/kznAERfoL8WZfHPBUveSDXO1h525m7UqosfXllJ5DlUSeVqEOstnWuFCP
+pf9OMyrgo5RSjhYSEZLh0tLjcWH923O/XxldSt7Jh4eOMkIs0HD56Nxtod3VOgb
1m6g1HvLYvTnK5n8PbRsbhDBiECSPvduzAIsWIHAT2Dw3IVSN5RsK+gTeebFZTR6
DNnGbnPFu6UVP9iQsxNwhNIEcnukX8Rg0qzgJbsikeCdRcJt1seBmuQjH7ZgYOmQ
CllorNCMdj+bpIq1P8IOcf53nm+aTMyGuQ3PZAFK8aVUT9+L9eDPnIQSDsWdz/yI
yIQcNXewzsezk1nJo9qWSCpDA8fHhHKdmixVwpec2Oa3MDAnhIpVeAdXx1AIDx08
0H1x2GRGUGUSLHmjsi5mQaGkERjSB1cPOf22P/y0AohkrJTmSyAYk6H/FXw5lKSm
4MMDrV97EoWiWHltoBoY90CdbI1P8IopmQZICd+18YSwy5g7Q2U4cW97YM4VmugQ
bEFVVVnRj/Y4A60uShgMKtUwkyrQsrfneM4ZHMOLNAOvWybeMZiJpnCPMBX4d2Xv
bWPgO4ENGjyN2xuaThpSL9X7IRVqpeWAVaFXWyJgUjWsls041yDXXfPE5D0a2imO
7GFO5AWsfvovOINyhseOaGPzaaYyOE7ifOJunz9YA5UnRn6fI+I5BFZfUjXE5y6n
65lrm8ncuBiBJ54KF9diFHfmJI/FSoJ53WVUgJxeho3yNACcyPhVJ8bhYo0nDgo/
Himyo4YTtZfEl/ay3mfn0D5KA5YbQyjEVU2IoMLNT0MqKTBTpJJ4oKKoS/BkmCsE
OHbP3LICWx2qS+v+Bnm/tFPXkEdd4hamAzG96E2BFwrzTkO2iinBwUuljsAf87JH
kGURyMXgOD2MqCtgbb0ndR1e7RLQa64+cT4AN5cRnkM4WDlfrLlicIcCiVzn9R35
uzS0MmXOf7gaZX9cN94AC/zJfkJQeXrXpt9nrp7Xq7m+QDU3PDIe/HyWU0JPoByv
PfTafj3JfB2sSuWogv4xbpXVjigjI5XFC9R4WDxiOIzmfWbqfJiKR8DCKvSKnjmO
CK697d49kHyfyjdo0m+dmYrClFbU/18ifCCaiyYJBZusA8LwXqEJT+u1DdIenPep
zUiBml7EpKM4/C2hXooTKDCF/DK+C94cliT+/tlp5I7sbRC30Fq9MBf3Ul5Y89xa
b2UBihMDUsYBx8bDuVmZiXG9OUs608Cdm9XluA6jsiRcss2D+1xEzVg2eP6iLxnZ
8Mt+Mo8RAxe0VZwQZ866X/L55eGpLm9ka5n81H4Gt1O+aQ++omOPoBrvz/reHY9K
qJxttKX59cmvsXlPJ/qWBiJzQ7xUpMR12TyA6aT6I7EGtqoWuC6DRX3Q6dKHVe5U
2xNfmQJ+wct0C0fMbGgChIdVXcXGRmEB+WWGgX9IbvYDyNsK6pFw9raID/FEdt3b
gNrrcUsbxlVjLgd56TpGeeJxbMn2NAyFvRE9T+BIUoPBGPdNg8vRMh7sgZW4TgbI
91p0snFH+i9e5sWvdbbUI1ZTJHDThR+ztXkT4E6HJXnVcRNbpDOYxQvpD8P1mdjv
IQ4K+PlW6p0CgFnkMmgQohY0XasuyNFAz7SKe7+BRPawPdTcPE0DmWrqk3JkgWhv
gT5zGRcbY7jlCwpg/3Q7EiqN+LBXLf/hY8wRZlQuFNr0QshRVrsplU2CcHxfDuZ8
xPZCvmsW2fDL8HKW3VPVaSn58twZ0MRk7J/vRFWy4lZq7CZOIprnBCTYSlHrIrOl
+6l7G/vlGIXfu4tD7Zc5h5AVtRlgIrLmbYKQJssY+THrB46Ke8eL6b2nnVi9CDJM
RTdPpPLNwXYmemC4vawo/bul6EgXvGWeuPmYc9+8J3YsuHoRnXsXDl1XtwXcRGFN
7Iw8OWm934Qqlo3FDORh4al2vIw5+75CVK7MNNtBM13wR+FVgHif6/uYph0eyjrJ
VnKBHsag7YG2+x+lRNrH0gUmbmc/nUIC/GL10ou+9BAP0dIpIIN47R6tjoSMCH/d
8dD9LwVa2wq10K7+g63AZBknGfM8aGtvkUymDawOZfEemxXgNodcWQqLMHcglPyR
tgGGgJYFCEkZqqtlyH2ed1p4g0t+u4knh1/f8EX1GpRy47qHqcq7xO6L225TFBcF
pBjv5yIMsQcbH6CrR72tiuSnMV8oPOpjZjvqgo2+lcXCvzM2ruyogN/26NG3e0VN
716ibib9HaKbic2/8EQBcer95L3NFICMWSxktCDihsQcff/mmymVyYUxDhUcdkFM
V8SdhrxRi8/sCL58WzY5pZTkMpXzuAul9KPWH0BRzX/ckmXqpqEY8FeIQF3GZoIP
apqltbqtcZFyGIW9R8c5AgJbjsLtdkCZnFBDyANTEQvXU0WqWy1seWBNYjzcFF9t
f/RtHhftsUrK3wUzMhG+K2UGViPAm6MyDplTn+yQxNN616z1BW0LYuq2q17v9Tk2
NgvbdWS7jqvphBiP5+jZWzYa4PS0oaHNNVE/3KpisCuZTg6bs9ZdXc4EzOzwbTm8
gaXgKGI5b+uFbYew98BFNqRZfjyKGjfXp8llFmlCAZrqD8b7NWIt4ese9Otrg7Lf
pS8mcnk1VPfoaAf/kOp0T8Ssh8ZPZmyixjxCJsWQeJIwpuEEkyo9IlGdwAy1TVXC
TW27lZsfbjVDEXh9eJiRqMKCmZPCBfY2RBebpc8+bi+O5sVCJXp7DO6/VVgf24nm
LrgvT0tsn0FCI8ztSvYG3WD0+0aJSZ8Fg6t7e1taZN3JH1RDZB9QgsYkFNFUfUdy
8ZKuUCj+y9+sSrIxgPCtkyUDiSiXmviThOBV7YZsxurnIAfgayaQP8hBVIxY6fyN
jaAcPuZW4GZ+LnNaO0MwhDD1gqs8cGPNZckIbYSYYHpin2ik8iMUnhW2lbNas746
VLDKBteGgJFGq7lf3D3f0csH7gpdedc1fkahRXmqYkE8jLx+6r5TIucH9CS7I4/o
eINrJtqM8zF07AxfEwuVQ3m9TwdqyjA3Lx2lbvgGXF/QpK9KIQccBMjjBDN5XW4f
A6aUPVBxBmlL/LG2rHzIvLDf6Zc49lm3VeggULI4knSbP+TjkRjhkzlbtXfSc+SC
X3HOZGjjaYf0vvErrTcYDxBEkE2voJ1JuDV11JXgceRVHt7wy9/LHvpwauN76qFI
kntb87pAM9UU6q4qM+FBjCI6Fzbr7fHdAQ22l9swl3ynCJbcKZLQGq4qpe2Md1IF
NEP55D/9scQlLlGOdOIocCeOg71dVhQODs1KhxJ/S+C9LXN1bLZFBpyrx86KvPZE
7fKexcNzXE4Q05NJxdki7JeKXQ9mzUpHW73alZN4f2nwymX7T5cXkNqd+fyk2KKq
k9P1mVlYUP6/t93w08/CqqevsLcYc6lSWsu6AUsbC9QVBaMzGGBYlIQxsfuILz24
G+FbFpPQRdjSmeVzUllE/6h+6wSnJOc51iSYk2wDSn3vE3WlBhG5zAUgt2dExhpa
ElBRPqhP6SoR2LEfoA3tN0q6hBQtO53CD/Ag62XBpOZ72RP1bgs/AQQKJkJna8w5
dRlB5rSjfYnZ3YXcDQju5ruhwSKNvNjzrO7qp5cXXFi8Uw2Fs7Hx34JgpbE+tW5L
BIv6u4mcsucewKlkTb1iHg0bJPLeo9qBElOQ5UaVFnJU4QHHBDoyuEKxkmleABqZ
fTq4r5A5ZV1AGo9/AK2mAbWCsPtoWKXRyxA4xGMHAtzzu5IHroA/pnr2mmch/i4r
TC8ErE0UKZNVO2DTbD0Ymo7W7evaPatG8+Na9ZvqdKvq6PyY5wROMhtpfbbZEUHk
6JwOjtyy+7pOdlOrH9t7/2ts2YbB/NlKa8vt5Z6h7mIIgS2zWm+Hhakl/+I5Q0hI
WpT1b/yp5rNzWBp2OBDLhfMGoq+VgpZjgVEDLWkhi9B84uWD+SymKOrJNxOrn0oZ
uVA7dkg4tF+t2h2hTHqol2UNxsie7Llc38IoYviqMSrxElBRqj5/z7cEw383MPB6
bkPFNedmVMdr3EnajmS30PgC7DtQaGjTzizHBHnYlpHBsI8Azqlr6XK+Hd+3p1sR
OmPyttAVY9r+tgAXMSSu49YF2X00IAl9pEi0qphujjnCdKomvsXhWU9V1ST08WRR
HAzHS3WBaws12eTpO9jcm38Q+xzTbzdoTe2rOLCIV9dbw/UTAI+VepMGqimDdO7X
+3LX8rxmgQZNXdcEuFcgscZyqmuV32Ggj0+rNihyd8lqxF44SbkZOoEJJdoQ5eok
zARLzX1wgnxt3Wqi1zGCjlIbPjAtOrOXzGa2EDjCLrlLpDnXblabfjDbvjMBZofl
QmoKoilk4si0K33Vt3Vx97J2XyifKUUhoPUhQYsd13cLxp0/Fg/C+wJ3UilsC02F
726Qy+B+Sbd071BygxQtSgUb7PTiLZs6nLIjSVhJiG7Oyzi708GcemCvhgtn/Dqa
rEz9/LjfOf5bS21BTIeI4lUEYGHT+Qbp15drX53AnjWSzTHPXUArAE1lJ+JK5fWw
137E6Gf21AfsAS7fI1dqFbreRNLq3WpXFMEk+wq9OSItdFidoAHeytELpRLWPCNh
l0EEKjiOuvnfWRe7g5cVWt0tgRuYvkmb3VJhpahqxDLz0pNQmVSZcuSK2huUQgyf
K1ZK/4BX0GS3gk4VaCQRCdL8s7FSSYIZd+vJz5bN4nGypzfHsS7UfG4a8oRSTUO5
SiB4BVf0582DAG7NuJaoQma5SQcEGr6TYZK+etLePazRPCwxL5gYUZ4tYQVr5VY/
4AqhCZO8ARiy3VSYE+VzfGPCf63b8D6EQSMe3kY8qUyQDwEQGPY6k3FPPw96F3Ip
SK+zhEb9u9AX8xgnaD8w3GjJGyxDLnm94VDBNX19Cd7izMd1iOb7hlDkMmTiV7l1
yCCofRS4C63BbROR2R7CiARwA9iSb2iMiZg9lzZf+rXEBZg85KnJ/3O9P6Eb+wZR
V0mIhSPb1ftmUw60u7kaIJIApm6jRkRIXGoVX+q0ztUeHCkmwW4tqF4/IM+ErAa4
DXp+q3j68Z/5//0BGgkxPfM13MY04rWv18lldym3jcGXQPjl2EqNLMG8EKI134Y+
g8jh4feBDVsiq0mGdpPjAwhFEg1TKoeMTiaYzP+zu0dy+nyv5ezrsPsKphloWCgZ
7Hvgh+l53T7ob5GYiwbWqVBcrdiUBcghQKyY93xihOvuNOZiVtPP97pAF6wwcS1U
/ZlKSHRRwOehUyZmNHClcewh5z17m3/eYhrbQ8V8FKemu8qMN6nQJKdsD9Vlw2BD
/gdCQS4eydduyBh/TpmKoQ4YwftQnAk4srkq+KtPNzKNhdrk8qXVfqv6L+rg2NlG
D2RquvSWjRJSik9oDPa5mBX6UV9KfEG1CRJOUZbsnkHC4heRg84BjwizhBXLkVq8
cdRXPqtbUahqQXnleTbTPRPI/Iup75jqyJGX8t/dZU+zsAKZ0g2vw8ygjHVxTchz
o6m3ZLEQYfY2CyO8yUQtvG1UXiA/D5UnPU7yQHXHBVwRZ+Y2xWEKW9ALKSH8cZTB
EBzc+l+eJv4sUVZe45capZurl7+q+3z36PjtRhjzENa07DvCFXtggeLbTVa3Fbvx
CbPtq6otc30ziktBHoQt8p9tPx/nTyG0TZyawkuZzMD040Jbh/zwxaZbbP/QZvYF
fCjutoi0j2Cw40LcOfAm7V+hnEgHdT45SPigwqNjoFsrr/ViaQ6SxOiLla4A/Slg
TSRQZuXx4/e6fFFGUpcDZLhMciLBFgiQDb+QQ6uHjkFLrJ+J4Mu/z73AeYINGR3Z
y3zS/YjFeZHJa9JhQ+Fh2VBrQCP1w8HvjjHRPt//TKOS9yKuCweWXbXTHH3cmRHH
fqQCwm4J/SXi9XpK3e7ePpAWUr8fKAh9mfR7pNOlHdMAxlHbBr5KvxOJ2O9Nq/R3
hZ9KxzVoGO2/HRgb13tyn+CXL17AW4ZrV5EnXtuRiUv56e5KHeNu6RpsCyXr0tRg
TQMcIocqV/AhHnS0MwwdbhXlvXSOL4CwFrXTvMD4XmvX44ankPn3WQ+Pglh2p6PP
g6to0bapqFVGIj1/e2apf+ztff26drtvFShxW2MjvU9osX+pXH7TDYdy2LE+RrHi
p63dgs3foAXUyELkgL6s/TO0R4ON87QWyQ20tC/izkjfYITjnnFbZZItdzVTNIUU
35fVs3I1ppmLXAgrzBM+rmhJc3iZNzLgQW7zBgHrbogDt0C2WijK4nTdiWxH9Yg8
kRCAYMgiDgjcKXsbY0lUvIoFF2Otk7R43bO3UYErbf83LyLjd+ANg6u+tlzthp6y
/taipjyePkh0W0xXmYb//EhLUcjn2WNtFX92VBRfrx8x+iKkrdVhf6BvMUBQhffB
rkmb56AnQELy5N0KuSEohzF8r+J8TdCJvDJZxN+n0IUXlEUmtvPhAB1LYmu68JcA
8bmNaFAEmRApSPd4ij31KvQhz1XifRl5g0G01x6XAt8aKR50j309aQ49QsaNf4Ar
YbgE84huWdfMfTQUFgx1n9oumGqQEMv9ep1eltdtqwz2Wg3wYcAU8dsx43b7PNZa
EuibCBtrFJc9I4Q5TBT/NWzHSRLcjpFPz/+sFWrYnTSlhxfFaEB3cv+h0lIUFaHB
R4bnnnHYhgPsJ9UsWuyICuKuYKX+nWeWTFql+YPuT6DiQ8CdhscagMBDQf0elZcf
4jhL3bRpR79n1LquJ94EcjsCawwNQh/dMo0K67LjWvf5a0LP0/QRKraaVF4NcRRp
E6G+vPQSqVXnbXcIk+ncNs3mYKFHaDovlEFHcHqZ8KLyRcQ82/ni1TkHRjHDEusG
ZFg6oLx6O5uYEhYlb6LWECJfXThwk4o9zAigDfP0J6zNbU37ujzimnXnBLmyNt4a
M0dgal+33RKyPV+hgmCVWhVAwGwlvzNa2Qov/lgofC7TxH/Dp1xU4Sr/SDZHsLx9
Eh/RnzrFSXEqR4qsHw7YH1ge+oXq456wsgnWMJvqdAJww7BnnLvigRvA3DBb/7f1
l//5/QFNfqNuxaMia80Bmtz4xH7Tl1hERda3OZSymcVCkuPYpjBlu5xYob1V+HUe
aYbrXc6EI18rK9c1jssOhVTQMOL+fIj1plNObCT0QNX/x8IzDV4yyzAaG6rcenE/
JJVVmxGRhDkriblLY2rcIu9d3BQbcZBlHBmKHuBwf9+TJbxP6rHue44gIdo6sVmt
o/fnG426VvqnEVC1JDbRr02pLknRTf8kUkzAvDA1cdGEzgamJdBYtlISozurVfh4
yRK9PgdtDbIpWF8TJeMYy3M4WoKn56ipkzc+WewtJCu+SG683ggtf0mgXp7/k1vF
dhTzOjHciZ9NIFgSVs4W5LibnQzvO6X1R9ZyzKBJUprSFi+G1R3v+8JF8L6Px0g8
YBIXoYQpbgFmRbHxYjXjC2vjdi6RDNBwKuE6ZaHgqBvjs16m57WvrvaNUJwTSQoq
XJuK2BDET5J7j0qewWRJq9HiFMS+hiXS8+iBnWsH+zoYgenSFQOttzAiLmUvTM7C
ZdtK1IxUbpnJcr6IX3yE3M5Bu++Twal2tbRdWM3p9ssj4tl39ue++1OtZt6sNaxb
5dBGmpaDCi/aA1jpHWTC2y3QVELf9EnLJnwuvpiNpvDJNcIYV53aIm8qf3+xXxJO
dTxrYe4sahGrdsH9UyY0nQCZF/Azdpa2kAw7ivgSSyf7ISoJfOqNedOhriQUnUWb
Gb7JQ5oureCqaGrlkOV5bk+v7WL+lc5Y8K3OQojJgMgpt/lfptvyfpBAydYvJ0Kh
ESMj5SKXaChQT5k1muPjixYEI27X+HExMjDtmi/m1ZlL0WrcE9hb8HN90YbyU40k
BN4Tnq9/EU9kPO+HlSKrmqdycfC6E+afIOrociZg6EmVN4TmEeVLv2V+oCFpKRdn
kkfzKzy0k6KOMQHaY1ZffJHMSsnA8UA9Z6o/TQsUOYLO2QR/6O2ReIwE6zMpgBEO
yYvrj/GfUYwT0yQz4F828SWldZnCnflWD3lDK7QMwPx05jGi4sVS87wWu0obdXTz
`pragma protect end_protected
