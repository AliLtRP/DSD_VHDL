// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:38 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
lW4SpQsI5Bm4VSksVZklZlXNrVz2C/ffb55P+mn1p2y6YHoFyFWESBPUGQs0zHr6
4CFYkf1yqPpU+aa5kbV/KMi8w4Z9XosOhIxlIM1crlLyv5/mqbRMQysHhMG+Xm50
lFDtTvy+TMclzMldutR8DrGUIBtPpH21rd+IfpEoe/0=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 4736)
Kyqc0a2XobmnHiKPALtqqTfffsb6FXF7v/C18p4tXTKzDdIxV9Q48xtAi+FMMpQz
p/htl63wzQi6DXWNXPEDSk9xYeR2yIqZcSk4ksf8NA32uzcDPs2MAmQttNSZQKPO
8f6TPLjpFJXJXgeytQQX7qZafnKxaN2ePwrklOL7l83OVAeFCjqG8/BG+R6QZoBb
m6PvtHq5K+ml+MnoBRZeRroaOQYWXkntFaX+Qs/bDwdN1BMONiSEo0XsF1k+w/7N
Ur8jxEmV3dkHIJVhcrzPZ1x5YOT/eztjjmpG/PN+vm5NPdIG9Rsx4JHiKWGwz7ml
XTggCdI+0xGxjZSHaT29Qxtl8An24norPmAbPFx0gJ7vdX1qBiqcajErsOH9H2MK
2tA/2SyKOQcSfoVLEHw/vdmbkMKDJ/wWhs3cvWd8S6RD3eMVCY9BNymEN9sy9Z2I
aIRne9OmGH4//VVkBLqq22pMi2az7ZgxVqN9pT2t3sJJQggrPXrKXYQ/0PYDl4Tx
Gdy/qoBVjXTZtfCUQ6dC2nnvYXsKZzEwn2+4ItBWEj6hxyFhszvPqL0PGaVAggSC
NLhKwwDFaf5jPCwhYDKTWsyJfh+MUnxm19cgAzbWpcmEcbxzfo3+gVY0jOFDYdPD
mnRfobiHN2hcBDairMksbvc2acJkH31wDzdPur9nYSyy2Vn3inwpdnyywNxCIl09
hVPeixhH7OSXTiHlZid2fGYgq6whuFaY2npRKVzS6jQSw69+1y3nk3bRS0iU0kQq
13BvndwDMeuiFgtNc9OcNWJGxcbdResFfCmK3u0uAaOYbjRy5RYcbaFpl8HbMBwT
ykwjv4Z3m8ueiz80xS4zpHyECJEU0lu+80Rk6I1Hbrgd4dHZeQnVypDvXaUJ946q
24pl4mxARk6Mq3uy5rSpA+FddFkNUMFmw30xUjDZ+2IrrHjbhMWf6l15UHP3JHLG
mCGHZXJZT9S/xiaYKpI/3KS3V2iJ7jz5xTk0vDjj2sY+V6QFiVqimaxwXIqL3Egk
NbWxJwZ0625zbmpwR+6bq5iM9EmuTQPLmoOSBaIV5u64YkMJ/siBmi7twGF1IlSx
FU25p5SPRKockicmu8FLTizg+0Y8s9CVfWMQaC/UR8pVzDHNaASqEpujqFTGRK73
MGXL5uDouF3uyZjWaeR/q4Z4m3tFw1Uj1BjWDhcNgqVtD1++aUCU3UJq0B6mGQtk
bG5PI8nfAio56wtIFzKrjGbWbKQu9P8ApBUVwkZmBgYXfXcoCOyRhMymMzcSDfB1
44EVCGR0hoWtb4vAeqznZ791NyYbU8794xifNzT6G6e8YiyQ6Jmm/nTVMnamjWhJ
VLL6cRc95KqSVYAd2X32R5hbopsR//IJPQKabRmO20txVlL/3W3b/D9eV4ULluVH
0APXYvtoTIPIcPa35OURhd66nfnf4Ft7lxSK/nJ36U3nPXRK3uVeExVjk2uUzJxs
rBZmDkZDwXLjQEgaLJWxuxLL/4mtZWA0UENjD8e8FwegQ0FNdcfnMLJVzlKd1vfJ
I6vBTWH5bVaFddS3EgIqshugt8nX3fY2Fy7y5ST7hclMEWYxpy17gKsNoCKuYAMu
fgpdHZwHQY3gi8tfhKGcAEPwTWz3zvnJXEHwvgKjQbMwV3DrzC7hZJXa1Jl4W7ey
/MgYNGjw3uwGXFrA0uDKbM9lKwyBIp1C6ROIa417v0rK0HuOFa2d818pOi8QzRLv
t81v8AAbPQIZS60n5LazkuG4RFhKlkWIa8xp1piOXh9hF113mFWOZ6BXITI4Krdv
+rrPC9OH73N6bQs4hEwuc/XKrnagMrQVOS49yPrCL5crmV+vR0SSZ/PiDD2hyMbk
ncWaoFEGVIKLZrWgCNw5YeAABYWG1npo39FxP+JRDT1uW7HvYotSjUYLEcffd4AR
4progpngMJUg8843nUdzBUPMvSnUa+N8eRVHJhz7wKSti3QYB3rqY3TsMIkZji3d
rzpxLZ7vMwNAfXfT4KpmSOff/ZwQugye7j3Tx5wvlpkt20YtkbZ01Z2cnRurl33Q
f76aaNnAtYVL3uOsEzv8qiqI4SHCthcEgEqW8/6OlhLXbGawyGB3wIXyVgQaQmaB
8ruBu5iGZpjmCu3DCKXutywj/zVTwCW+LdbuZS0Rh//fmGWPBcZLT7BeqmT419KS
7GsntBtoR7xn0XascjsWXsH9RBcCJspefIEQlVzdEEpr1fpVPmV1zoRsTznSFgvK
BO2N38us5gag8QI410h8wsDW/0VkXKUpDS5pY2oBO3SflxagO8ckBOAUB8JryLlF
7a+kLI6uEIX6iU/WyS7uOtGlp/k3yuMLZY0jeyES4lfg6VXlj+cE6OSjwq5lOvh+
m179qySAh0krN3NSzwePub/co0PnCKddRcsY0QFhw0ry7otliMvAeoF0PIV7f7Mz
CudMRObFWAfD0w/LMNgN/kN3Zb6wgGzgf53cnijYqmoIPgK6OhKkLOhnHWH2vw/8
linPn97BAqfuRZb2HnFvC0h0DdFIW1WWhngNIVmjKZYmZc1nr/faFNQhzV0xDqSM
G0LEDfpvX3YToRYsAkDzym/ryehcaPlecTSh4HnqBGTsjt6yUP/dr8WFxbsyEF6h
ANSoNM2//Xht/O46w+GJm+v5jBb2l8WGozV7X9jbi6hI9TxKPkHF25pn6peT2aD1
ohqs6uaCgczZjHn/jj5fgjr64wZn29R0GFIZXzG0S+daF7guCnI2hTK9Zu5Vas08
dTLGUuPvMHybhw/Gsh9FQFp3GuebAKYELg3K+PGnkhpUOQ566RSKbsVaIy1wfmmj
UaNWvcMLKNfFlzROedqL4y4Dr7eWyIWMn9oyByaEttYRlzdV1+b7OYbkjsWZXCh2
hNU332p38bVZsf/Dw+MUhJtpdxI0iCHLQilxnOvfNTOWTswYxooar7eNgWmze1h7
yHnLLGBZyamAk32rmzgNFlWGACGpK6Vxrt/EnDSGUzwFS/psgZmAAW/6lpsYnHhs
WDZOCX2pedF8EM81JWSPhOTPVqazc5p0bKTyJ1l7t46JFGsIdVutEQ5D7rgPGtN6
aDLr08IEdmh5Z5xEEbBynDivyF9fnQFHFQjCHt+rQEio8EO5F5psegOq/2flysTN
iHYgzNrYi6KiIttI9tx6dHb+6Xg09ULjSN4afQtRaiijzMpvBWSc8nbqdP2Sz2az
Jbd79DUj2zdgi+LkPvlvQzIpQDgTHjs7nIDlkTVUr102JqNd3+EytBbNPxTfOjUe
2ZJyWVXyNjjD3Ht0TdTQxHDp6Y6ScA2avcEdmgYjEdtUVZ7DQDr3OEm0RQ+2xQvm
6FDm3JC2jd8XirJldX2MY66/+9xmBc8ZG6LqPNmehy5RAqt3RyEbW7uKyQmEIaf0
CyhbdMNpig2ZZSh+ZxJnNpdnph4Xrik0KCBKDmXRG7BqfGNktD24+4GPmMoKYk0O
39WCDttGmjWDkljzlLRbCXlcDjpLpAYQEX4xx6qpXt5GlcJXU3keEeUix+eX6T6y
fe/Bz7AkFbc0YDDaCX8F1CYqkOnQ/BSEcl5SM15pF2yEMisanOhjdDANeyISq52p
ShBHuLKj45YsBKaoLxfzLvx2+/qDqQM9BghjSSL2U/oO9xK3JCrr88Y5jX6AGA6r
J1UVjpVtLwB1JpDre3XSLJTonPcLrB4rSTIhQXT0ruGaXs0qsJgbcHM2zgP500Yi
+fVlCmsdm6T1mLWYDJWuRe4iSQdZwsIlYwCQBugjStUS00mjulPH2My25J2iuBR0
YMbs0ixv3z5yoyH+jx9B1+/hvf7C5QBj0XnjdN9I0JQM6EA7eanS0EJsWmJnW2pR
c5jFX7JQa97c4aSRK74ST2WY5O+7ehIHFYzOaUmwljf1Eqff9ac2YAJPLbeZgfUp
w7i8xyvAZ4d5yG9zOXxkXCDBwftSSjL434YMm1gjb+Mik8t5ikLscwnZvRXGUIw8
iNGHGsWHBNSMSvw4TxLCvyUarAlj5Tdfjl/7mO1mWn8z6gXuXqBbuejtMMDHpF1b
QwhJiYYg8U6fMo/5pvb6lQazLLXscRD2ug8JJuZWjfoEoX27oGhYzvy3NqWjGx3t
Ojq0UZe8oRc9r8HR/ovZoBv0QkbC9Vb8fWEE9fHj/GecV26y79++Zmt7R5IfgKxc
PPQSwx8Su5qJ6VO/IPPvS41WVTBE+h4Pibj4gVFQv7rs79cr/LXMv+rVULQuvpC3
zucAKgzsv1ijKgaNzlyku5nlOXg8MYvaymPMHPmZhBxNtTnLOMOsQHHUndVD09d/
SrAV3M20V3J43NZ/GUuWWLulcwoHVIxISwhXyZidhVLK0in/zWU9QTSidyj+a7PY
9BmdNQpIZ4LkvP1nD3um3aNLEN7eN5NzRfvUkaqzJsUGa88N6QxWjlT8ZysLPmP9
Kd4Cyu6hdiB4oFhkjl5w2E2NFhiOp4nJoxvFpmbrd1s+PJdXB6ufeF5PVxn5aPMy
xnOiMA+nI4HLxawrvj4Qcdjtz2cW2vKy/asuiZF1P6Y25NoLjT8hUSEr0J9B489e
K1884x7qs41sWDubE3RNKqpAfPe5RXm81DUVAKXEGXUja8zLQfD73A2wOxGyC5Mq
2snxnJyD/XK8DHzspaYvfOhfPh++Bj8VznVQifCro0YEwxeSsdXf+tNdsP3qWBLm
x6lRaAba9wd1Z7wLk9iSUu8J7+C9jHOiMvm8ZBmr2uHubm2Zy28eLLUX3DN1/fEC
K2XrSEWYRKk23b8uotjhFOnC8DuwfWtbI16DH+lpvDHZe60to8nGQ1VeD1cHeTVv
gkURJkDj3HEd/I4vuiaHdm2fRraC4OYw4yUB1HsGir5ViVAOiOI5+jxXmNxQcRoO
xb6myD0xkAePjlg7KWfnZeC835/mPtfwCCIQyaF9l/8w+Wqj1x7MwhlCStRSxSQx
vvWcvzKZjA7LPZzqp0oE8pH4kY1ncsGSmCj2ogVHfDtT6tmadyPqAomVoGqrc3FO
UNcW3qsBzL+V8V6arKLVjJlQYLPoOt09D3RCg2W3Bfp4UtTm8O/ayBCzF0SqxxlQ
/BSutPlLNTwTYDSV1DwW6hMaXloYRDp2ey+vDfTGTmz6m2kMdfhlrZgtozXBRWcO
YevZw6kLfB4Uyz+wbCeVzQ5GvWXjWo8XNA5btFPXHyt8BqIy65Xmm90eBfS8GltA
BPwsLMO4ZXwwaanPzRffbGtUueGboEuZNriqXoKbeRvY6eeBCqxnE6RLk8sm/ExK
3+nRkQ60LixnwOcY2YBtv1g6hcVvQxq2aEi7cNPvuntrW5p7M6Bg02n2Qam6C1V/
eulVqJsGVtwkujqF0TUgZGua+lWtpsxeZuNPqLV+pqfjVw42kh3qrzFUfk87l3VX
ryTgs+DdmKgn3I3Ij/a6Zba2Bvq7dkDumj8nvDHuH9mpWCond43POZSjctKOTe/v
iTPAv+SirUAe9FFPjyaubTPzNoqkMeQATviTHvaPvwEkDrNbaRNiNwPHI5YZN63Q
9Z+IR2/dDOQjrygSjr6TVkRMNPoUbh94W2m9tCcdsvNpHpWsOcKmh2W686Bobonn
qGBXLXSx92ldq01DtKzYTWYek513JHlZuZwUDwErLZTU6ZDyBvGNd1DiBdjoiD9r
hAtN1esqOOwgyVytdRLKo2KQDdzRhWZjvbqNE2XMjZeqyKjcKgH2BeThRgHtFIWz
IAbsHcfFDSKUtkHaZR4hLDM8npqu2bzCaB8ttOwmaTKwtAEIuTkJITrkjsjOCBNf
muBHByu7HUvrVsiPl/Dycded6E63adroo3Fu4DhrSZ68NRzK2oZ5KnJm7sz33el/
0oA6CUcnurNeguOpOGvLvh7xPKO5UD30yjm/Tb4QrLJBnm5fMQ/dYq2BDFsPe/tE
YuPGGF60GQhIMnhAgJgcIYVV066lZbDGslgKFxRTHhr1EB3YRH5daLC2Z3B5kBur
1lbshdX6Y43hFzJq6i4jFQ9dPH/8MXceTOnfKhEmPTWt3BmuPp/MmZ9qMVeI6vLM
sMDYGym2vbIXR3s3ql/EYV1kIxgiUdt8E185yKKE+Tdfw3eiWcYJO8xgNe8JidFQ
sslUiD4WLuNsQ4muWQtxHjIHHspr0RSfC77XuqxgMsntcxnQDe70z/V3+xNBuqQD
2p+F6ISBVkAhwo6EG5Fcu2lUpMQI8znuc0uAOux0W+yiIJxJxzS0bE4fTyQUUrml
RDXl6P7GVnRf3EcDP1990OO4TwatHvlGH/6Aj+NK0p/4W+8b8m4YL0U9sAqYiQS/
/swRuNDpnR32O+n6exEHxvwts4+N3/W/kPlMi8oH8+M=
`pragma protect end_protected
