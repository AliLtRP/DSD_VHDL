// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:40 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Fos4AD6DT13b3tP4cvcM2JDjXEwFOhHkrF+qk0ojRAVDwF8ZtltJad8yULNwQUyj
axEzKyYug4iLjKrHN7sEjdDyyXgTYLpEep1PYuaF7G7a5ozn127on0SHVpSde2M0
ZNvMCXh9x2IskUULa1sZgFQaNT8Q4cSsSkao1QOareA=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 6400)
aZpTOaXcaahIqMR+XuwsC17QELsSwS2y5dUD5quH/Hy94AG7IgQVmOqceGgNgwtB
aumlTbvFfos/+bn0vRf6lTlV0Kh1k0gO5hRnnlVGp2NKZiNciMOFgT+DhQp2XWAt
8TZLWZ9aPWY9YiNgnTW9GTaAdIYEytYkyEKp07rrInqLKwGZ2BhsDP1MHj19mb09
rRDWl+BKmHSmsHR+QOp/YnGlkwG8XWaOkKBLIBZCzlIUXbmC/t+23WxCYJMYRQEv
axW/SL00xlT0G15sN340vjeBXg0iYzMpG9zmdnxaqHrEu6b9SmbHsJ05dAzcjqXP
n6rsb7tj0wZcdLpG2FUb9qZQ0cvfYBAAfG9bhDkh1R48Af3g0cSINlzISCO8hUOh
bJlJVWVGIHfSb5XViiUVm6hO5VPgDPfEEc65g1BsjEWnQWJuf+NcbXUQnp9vC9QK
l1G9JKqSC2RjBGHEmXZ4rDTtwWEzhp4CkFaiJeg09R+jG9SOAIFWdh3BTpD4tEmh
V4hjtvwiGnQMHzbj8mWY7C6RRqHuAZ7IhnOsZVMRCe+aKP8c4Bz+G+THYE8EE8dL
PQZBO303iJn0xpt/Xd4rZHXfDK9/7rdmpfVY5uWU+nKTucZqKI8Pkeqo/AQQj0fS
EYvyUroH1sO6gfDtLqFZeKrkWzT680TAlQE360sYk3PrME61+sPCLlB7HkTRvzoq
VKmELf/LRzIkcwu49aONV1EDJ6an6XAgwf7UWAiHqmW5FbTJbMG1P0YiECH1wdr/
gpk7njc/xym5JLJUQUf1udCx7KO8mGE9A2kNBNevgdLwQglcbRZIlngkkpgECIFo
W4XIhqU8jbF7TxGXzCGIaaj4o8cFJNAv2tngzGPCUmaZpxcmJJ5baNecH0T5Dv66
IEuOW/x069fY05Ee58tz/w/b1KeotY0pT/ZKG5Apkxxa4Ahp5PIUJek+08Sbihnr
14ZEUEJ6KMD4eIsikHFV2BROCX04FZ72Ced5yqy+5PY+guQlj4MXH8pyFFk9KLyV
ublGDAVLLct3Q/RiVXa13DouSY6NbjvC9KF+CKJDpYSetFEepGnQCpkY5aRPs8xj
pQguKs8qJ7CCiMIybejxzN83+q5mHfRlmtJpu2pTWcWyo02NDNMK1g/C4zvYCfyr
BIg/Wwz+FdRkyHt0YrpXDe5odXT0Iqs8NxzIIglq+XK9KQ0AMU22TexApRCiDA3L
JD8oD9Oir0dJmrDq3xfbcbm8R1UgV8vyiEfGi+doF6pq907T6uYhmX4VIfaqM8rA
Aiv0N8p0dVIzuzVPQJUmoPM4bey87TRSjj31KfvOEa0zbXNSf3DJLgSbLc6CO5EV
AGqn/j9pEC2RKJyaJSnE7nLkWv8ad3Zw19GROCCmXWKKIZFjVfKhrO3LGDRVKi+e
QzbKGb0v/UBS502ZEU7Ho1TDyS1DUif1IzpPKCA6sijUgzQj2iUTU8fpAADybwXO
Bfa+R4+r9AsHZcq/1T9uzE1bDB7wQISdwHSO/0XIZz2XuaPYr3sHeheGOa6X+TAC
3u+du6Og928s3qJuHNtcLtUbuIW0IXNg4JG4dQDDSNkiMpNtq3U2NfdeRV/eRpBY
aLqhJiZ8P4prZSrlMlin3uq4fc1xsgMgWV3W6IUNYgf7dz8PSAmgbNpK4FI5u9v3
cpGcj4YArnIngLXkTdS0pOWCb4SHhtUxAAX/Elc5X83MntSlh2DXMtZJHyHmQ+K5
WHrIXnaqssy20q+F3/0Vr3Zeo9rcc1usxNvNE4X0LJ5Hr5x92qWvhtsfyg+yk9M+
z9vakkBiclO5cBFjOHUFnamYG6chFvzntLVjnfHkYYTfi0Cczog6/kYorFV8GcVO
Jjb4/XryZr7eMIcBAASTq/UaoHai40JZlvqEIg/WONUUlGYZ2M7dYZXGFHFzE2WA
vjK52p1eQvaVCmDBy/agcKCRikh+/MvTvwEF5iZS1on+81dk5SNe3tNGxFyHvO5A
A8iTf4Q9i9l/OtuArtmh2XNL+xoo5qYqCBCpFavF2X+0FyuMFFfBH7quj6lzh1L+
lE1IDXko79P2K61CqB/3Fl6K4F9uVcSvrHFsJmP+3DBsd5DC71Pgwbu9F4o3AlzC
WL8g9CaXoj5pKc7B7p6TtLl98RIloIXjLweTY5cBzr9BqDOKKiwgiKhAtjRfmC0E
TsVeVvRqfqVXNmMbsW11dW+p4nnUzhrxy+TxQoo76jgJ15+IF/DGIuGBc5Xxz1Fe
SaAKUYDhOTOQ3dsTL5Hr22NRMITGqhLVckCUzdeF12VHlQgC/RMnQZwggaBuGrNv
sdIYpvyShmXfw+8G9z/RP23FKz7/H4FHAoe4B2I/3AA7IHPg5l81HNmeE0IB5pM2
HdLc3sra19zEBd8yJDG9sr5TG2m91jdj+T0pu87LcexMdkad8NLaWdq9R0k1CYVz
HjU5cgAeTGcQYQopmOjFMItRCDxHro4wALcCYiYxRT+gtRoIO2KinkkgU80C9SDE
te+KqAc9UPf6mGYN/17KY3nuTDlm9VwAceIFE8lYLPVWnrREwwP9Swj9jP8IdSDK
wKPr99bcxjNRb/yhOpm83k5FnX+pf+QqM82wLGkClRkJelQIVU3QdMk0okA0ZuF4
PU9sB5Zg9q4L0kwDcUlCwsL+1mWwlmLfKIHaBz3tMjoToz8rZ1JivMaUydcKftZ7
+6rOgJ8OLnyeyzcNXNkHEkdFVGb8rHap3/o+9SAtcd1hOcsNME8AzMDQmr9lRPuZ
UYlsBEPcZOfElHvjSo3NJUC40p/GwMoFGe8ad7ZfIOiIm7Rs0HqOyfWsq5sDivhR
n1Hxcmjlahtj4olCk5yn2/iim5NV7mUxhRSrQak3+b9TIMfCLv3wzbxMr3Quvrla
WKHi3MuGWDwcCqXqhhBVIZ47N12hGF2qIWUTiQccJhOngu2pSct1/2XU+DS/Q+Zp
Vd7P2FyIw7S49fcrSwENKMOrEV0D8vtr8mN5YaPZC1nUmiOz4/lhYcqdxAJDJs2e
eSKaHG+xJhVUGJMnHjck8rpUYTPWc0qlN4wqZmaynmvn5YRYCQOef6VHLbYk044s
zgNcNbB0MZdYnrzGaUzaEQG1NBa3oh1k5LzSyq1lCKTiP/Pinl7doLoLqatI/B63
OSWAafNkRNZcQ1ALqhStr47+5cpqegXnHzhEs+8ekwvX36MOayEHrn4jZktHqm4C
tr1a6aVCI+aTgnPe6IdBofI9qXnPfFpFF7y+E2SdTzT/X9xSHgYwnZTVrhnQuEuY
A+7u5NpzOqoiNqDwkSRWd7terjp2UHi0tUpiKs2+FZYrsHrt1fqmpw/YEOotY//Z
BNeNQ1zQJ2Oudbn2g2BWl1fOmicWE3wci1aVqeUnGu4bBiEJO13DTTlhPS/1JIVH
Cy7WOsFk1oAaYF5nEFZYLnNYZ4RAYjgqmo/4p9D5oFEXuH6LoraedFBc7Z8pXjTW
ubLlGJD3lDh0zaHcuku33cJCRW8TdikiDT4AIdqmIwA0mdVQ6JjIWh3d0Acxh/hf
9+MiyLEnCwBRQXTXIpdUolRRF5wM0qXLY4AdfqtbWY0voVvHKa2MU8Q+GvOiR0r1
m0PuvmdYT6zAKMbbqHsJR2utTZrTw7x9HkQJbK3bTWno4vb6drGWU0tPicqSosNb
vq9UJvWYiSOSEi2lYkDpDauVu2jyMlt/J9n685qeg1HR5yNvWdk5jSge+u57u4XM
1UUyuR4R/tg8qo3NsU9pZ473jvSj4IViSmWPnZaR5d+dFIpTo1YFPeDbjtH8iXRr
qK5pJUSi6MUZfXIgk4V7gQaqU0HHdaPMczwKhglUJnmEOIRp9ryhGaC8acnkxtbx
eeDBGqA6vZpiTvVtUquB5AaJTZJbHF0uvGVEhC2bfQpPvLegnQq205rplDGS0GJQ
25PdG4CwTfQOD5jMyVTqCHKY3LpORK9S2WQmJjLsATYXFFSHM1ys9m0jJK8Bl7SS
t2Yrpx6m1Cw968sqUSl5RC9/G+DhVv05O/caA7CY7pnuu1iW8zrFHEYQW85GGKgK
PnFHzwfK/pEVv4UJS0agVrZxfAyOaVu5X40sCcUExCG0PW3TIJ2Z/78eYyDGCEMo
W7TgguGrI2/gZWSh5syNyEin0ummc9M0lgLRZtKw2f7KS51CC/WD3Gooq5ltFkgf
VBihMu6Qi2QwF6TAhVpE6G33ASWAIOVdQj5uQIePRQ6WovIougrLpfI+dlH+Dpal
jB3bhV0/gXi2TL2nkuwbS1+zVoJWNh6w92PnpRBnNF9B9x8uSCw7NWH3rPJ99NFJ
mmzAZGQ/UnjiZO2bt39R6g260iWFXAkelAzZuKBYWGljKdYYPYdPSOpNESytEfWV
X4H3p+q2XcBYgXyAJmZrg+MHEVXn0QnKF5C54lU/T64l+tGIJpjYac5C2r0vsiRV
wwTkGj5enYArc2sgbT9nwnakWkMm6q6HrFlvQIkHhAxZBFvis1bw6b/Lo7O86H9G
hYAYMaM+Ijw2YuNti+yWxFHL17h/udPlSP/2MKJ2NVQq1zMUX7jxHU7KKQSD2uoU
+GFdXdlsQn/YqRjWsyPACXDRbEMwz+UeV9pGCl+Ed+6WOQbsk0A3CzULOwfp2Kgr
SC9setkHpjo9r+/aONW+QelM7kGzyjX4atMupG0Bk1ekJqASrkUrMuoqs3tF6smp
ac+0TFnTVPrnlglAwDPTnaQHwMm2xoHM0sCfgTDEHpuYnOPKIcSZESLX+HJ0uV08
+DU/b/mfEqWTkgyndXDYUKNKZmnV50gD0D6/yD9fdiBQnroAwN5WC244UxjQBWZ0
cgqT1ERCxvDT98gNqrqCWQDhxI/EjJBjiZyItm58+gAb9vPLyTwsDOTRibvkvIqj
6AdYME9GqrteINu8SjjI2IxrqrgnaUnMaQNrSR7HKXOEmNCqbJyBBXLoqqpKHXvf
IzSun5kVMuwV5GmA4hKzMWqSe6uNJiX+V4lUDQCd61q754d+LSWD/Vbg25Cfm8yJ
JirStNfIlC3270MWVdi4H4blItZW3Ojz8X114v79Pns/r23QjnYvkyHINYMEo0nc
0SE5NIsdROdYC9tDpHz5fE5V4BSmbft8qHPf5OON/PdrtdUmjS9q5CUfFSw1l25u
KLpxvcCva1PI5kWyf9m8goeO+9Oz2aNCfc6htF+O2n9R8TwOtMnNAPVvtDbrqINf
VkIyC8r2jAKZ2Y2EEhTpi2aP0WvcciyYe02aOslp13kaXJ3YsTFpR5bP7T1jKVsh
9KaFQBlGc+eH9l0Cm6DQeB13vvQXqC7BxyBskSKyi8etdBA2rNgBdEQkPoVwva9w
MkGgGHVkIpt0tqXn05Jdx9rVlcmnXqd2bAaO9EteckVoUn06cKH8O7pp4lhkZew7
SNDhYBnQVt/XV6QxJ7dnCHX+LNCrFSYyvp1plWJhN/VsLDddCdqkBvc7VJk4gAzz
sF4MmVdRm78lmOahNPTUjX3sxqPyzX8BUfT8y+WEyXAftRIR6RYWXEHA1aFqvoTP
iqrALTQyBPVHC4vjQEZwNXUCz1G72CfLN8mmSTtsNQpNKcD6DxsbpBF2m+89+m9O
B+ETtByfGtaH7fSvwHdA+l7N92A0d1EXBDYJhU201/s8pxliEiU+WDqhGYftqEVc
TqFer4ezeeVOU3QpO0ZXf2iqo1IvsBG3Tp1fozqBkjBbKygmpk1LJSltdwlxdHew
UWnrvfbTIT/pHtyKSUhDRUHxoHEvOSUDFg0gxELMgU04zau6+zXmn5AT6h7H4Rfj
qmXQwS7RtJGWvQYESQhSE8/nTytpyB5z3ayjAge62w+26fbiVuQhjinNyDTldffQ
ZveNSdEj28zmJuysqCVNI8XoUz3JQHqTr43nBIwSCQj7VvHxVspsEmvkH1NeGNMu
GU13tOkkhZlqNZYbSrhNZ7nHmmINJY/VgKKMmZjtcXmPsjL5CFsOSWuAMlwoWuNv
xL6nAPxmrBT8K5Ntkxrb/jhU8AdJBROG+ZJypE2cOGg5VEf5J9TdoRVgCWZx40jV
53ML5q7RZDXYPaYUyPz/k4pttzdK3zdFdRM3U5vwAFBGw08UmnKV3k5O/p0y+qPp
fO53G945PFaADOHjU1QhLpQ7oxkHb3dwv+NWzYPzUrXkxoKO5ucanRG0rdTtgDds
NNTmJKrQyGHhYXFn85UNDDQRh6c+YxiISkk+eLGGuMirSsPeteF81QqZkaDhzAbR
1DRUkPPgpeeI/1bHDc3iCKWkQeelJxa1vDncekt7ySDuLQWNSlMia4k5DYwH0lbv
yJ0HHIDM16BBvLSNASFpxhr+l2I3h2awuqISRtugg6WPwGpHGXfDeWBfsLFm/Q3z
1TYU95XRDE5cn1hnHaj7uYD4KYBenQbgllmgo9MrUVJ5n1dwool4bOfAgOadrYbR
zmLijfiY3aMTpQWAMojGRCVHYoW36Cbj125dC0TCB47dhZ+M9w69QXbpj2PxyCKJ
ELiGsPOW+YMqrFiMXdaNo2ghSHpKOryql9EqKl1rVsWF8Om6paelHyNCaR7eedzC
OEXoi3sz2BlEEKWRnzzbyVJZ90rbsV4I/MVw8v/tl9Viibnac4wLTuDCagEg0EgP
Qgh/vGniMvlwMO/US3DgJ+LOUoNE0z4R1n5t3XgaOFAzAgcFNSjw6PbAwMsK2yNq
x1MWkBOI+rlvPFvmf1/0hJSGAcOu/HbavLZzOJ16Wz8ARILyL9l0Y8slWcc02Dtx
mTYRgujNOi5AAYGmEV4OWJ72k1hQ7Nr2My+Un5ffF/fJSQtVtnBiWUkDJJJ/7m7G
2JEEg0mmweQxfIwjshmqWZeYm5MAw92ECJyNMnb299PRsICn1Q/AtmlrntwI544+
lP5aJRJ9ytr04sF4J7Iu8ugGH0Q1/HHEYfmvt460W7qfut75lO18xuykRIMebJxr
xO8jsaWx2wS4jM5yGdt8V+EQXNFNd84M1MNR4767OHasEKL0S5seWe7GLAy6RYJP
YmUnPCMdAU2cbUVGqFc3L90hyEysvIvB0CKmhKJliaylC0POAaXVx/7Ub2ME2baN
MqD1tLIoKrDYQWfHFDshOWyTim0ybZUimPBMwQEPIik+PUxJc0UUaiYqGRMDhDiS
8Sw1AiYgStN4V6bTnW5j4VpygbDWR6X4RXqTYoujJxIt2JRajsvkDNWyu8x754w9
9EHgj8Jx7BEFoHK2IIF8GTgfhpoazGSZCAwxbtdXp19jjOH3kCV3aFU2IPjXw1+m
/YL+Z9DGzijJzUcuTxoZIEnwPiGA7u/xeQ+g8wPfNcpHGyTqWW9nv176J+RfO3Sq
RI8mNYWqGtHLyOph3tV+FH/+8HYbtM8FYMV2+MixQMolNw6o78ORlWL6rTjn06PW
wBYBT5iLdK+dbqr45hKq/PyAuCnVhuyd4RTndA9Kfqus6OCqbeVJNHTCDp0x5xGg
mpYZ5zu7Jx5NrkjEjGLbZ+DoilLRaqY+vMMzSPsadO5LkAZiG5y5CC9UReePHlEP
xIufqgIh0AXQlSwAv0vjPbICk5FJGjrSSfmHy6zZiI95TUtJFuCpxJB/iJaaxShk
CbwQTZO2AJqyLHkOlSBQC5JC5VSZQcBwO49wBzO1ojqgXMevW0XLqfFVSrjBoM6f
+SjpxC40KCZxC7DzVp/cZoeRwN8Svcs5bZA5oTmnXcfml2iCNFB0cYb2ln3J4kPc
beFKEaZsw8S2chb78UaDxdkmgmgGljZlLguBOudRz6lSzicRK6qiwL1ZVcm1ANos
kh6bb+YgZoInoBiM0zasxddwGFwUg6WHuiMUIHuGDXRXHkVp/8uSHRYFoVtItmEi
rmKFqnjiTAHQxLZIgF2A3KBogwntTZjcRJDNL7Do+w85iDoCQMVlGE6kjVQMMrjb
s7/diDhckVUASmbZPCyBXDRyposIS/6iPHm0H7hUhG+j5DrdnLddBI7FcXIqo/CB
LZbjt+ykFnlngmnyVNQtYYrrt+XEjkd3Y4jhMVUMxFA3idcDFXr31DipCYAcNDkj
oMJI6685GsbhlrUUTgCHMmY0DWJpx4BoueJKyqmag0hVSgDjiuBESlUXG/wD1kE1
khWtFbN45mo2vOG2nk1DLbIa6N2nyyI6ycjnbcWQGtSep/Y+Xr1i1KfFImwWNZ2m
kpJOtqP6KeMIr9vSNHgUWvCGHd/IPnXM9SckQ8Wyqob+YVD308sXXM43qfJScg21
pI7zZE6ZsePd5FtxQegtldJwWFYyDGCJaK1L1Q8b90UV0aUAo5BG7jg45FCCTibv
7WOL566kQhKM0i+SJK+9JaC4I+foFw2kDK0AYT0msECXjWvHrl9MriP3nwV65fU7
rYzZPGZoT1xgcnK0KPkzF+70hdkeq8KIwR70LMFXvSYLO90dQxcwUbrAMNa6SoJ8
IgXCVtVz90YOxHM/zlIAiTzeUSVJZdcjnzp1BpcUQYNE8SFdCmmUj2QEdDSLGuCX
QIo1dLwF+Erorx0IoMZmV3GQuOu0Z5Qfx4kpByElx48kPC8Iy6kZllJxW0ltFOOl
T/Vm0gtsz+YoRmNlInJGvg==
`pragma protect end_protected
