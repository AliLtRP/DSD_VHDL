// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:37:20 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
PIi9E5RO7JyvK3wBxw7HC0trq4gX6ZsA6fPmgcSSpRQWXCw771/hw4yFspqH6G3N
3GlrJBt77/D5IrOQG+i1Idwmw4Kkz4fEf9caSL5qqB4mCzXTZANTm2kN90HS+6Iv
PccNWAejyqYjzaVVau7KW9T7Tg0dTgphn2sXwIZHf/Y=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 7872)
6gohzbf6KT0t0LGk9UuaT3lZ2YgZb7KTQFZucT6MZ9RoGpoIrDGV3zhO3mNYiLwI
4t6GJ6SQbyxalm20ODnYcWT5QBiwUfYXvwKPKVJtxbn4RQWVbwlgqbVfaxCAkhJ7
Mw8BqzcU/qzMxfIpTSmV5eIopO5+jGFiSwy4jlgA+/KSOwE7gobnluSNqMbuh7hA
S6IKsh+xzsntHekBWjBw+itnqwXNDPCLYXWaUZR+OvWkKC14dussTWkPEklbRTPH
o0Z5zjQfOplwhxHd+gmCj+HPT5TCPTOSnB0vNyBNMia8fu4A0w77efRb6mxmSbk2
KALCoowWjPHVXRgold5n50rjcOIVzc5+cVGVnQgThZXf5xkH8aqKxh0LAN4s8NLe
BZUHTTG08Pmko9ZXjcNNQAVGB7L1dLHoAVBXvfT52UalRe0z7MHfgpQE4jR0Gfun
5I3fsrPUVBJCY1Kse2bxZKx/ZAm6Sp8x6J7zFno6vcJezVyvGyB/7mGoYu4OAbII
9PMVu4XbYk2tzt2h/Dqwp6ZgZ8gwDsG6DdXNF/8g9ktxjKcqe/0lalh1zpRFIAJk
V4hFlHPu7IXKgsK0WIFGJWmsRRZdWqB97EaVpicyvE6FJ/ZD5fW7nUij+tjRBys1
qpwC2MdVt8ll9+odFXghNyyJVn1jCjg92sKq74yhy/49xvOV+QyfviGVILE3vZkd
8GdF3WVgpylBJnBB/oSY0p0yN/JEpoF6KpHCLJ4QEahw5CurBDmmLwiYoMFFZCnR
MSkhwyn/bVF9dRBs+OzFlljGBSZUJ8RVls8tql8GzYjf5UPHBF+oJXMeKSeGOOGi
gRdiPAnOgnIvcMzH+yx2EtT+vwuX4tujjQk59ERcv2an4B2OS01di/NzCI3OXlUT
usWmNPvley+P7SAk0Q1gEBmCrFKqm4DJd0NyU1iSLDkRmkkbPXl8SJKPqXl2hiqi
S4tmetF4l3MWqrlcJxBb4Il13Ey/bw1NV4eC07h0McqW+6aNWBjwhv956mHvCc2s
Nrz+kmowHM7tF8ha8w7xlmuYtewK5k0ISNIsxro0C9k1IyHgaZ6WMQc9IGarLDhY
gYzp/xmyuoJaFKK2Ab5kGV0Dv50TzgzBObcYAxtKSGXvVx/cE6Ec1PIgzhBxLbhg
7jhhBf2y6wgvJwQJL4sgZbC9dDVq2/yIsCLrGfG0coL40NLU0PY3S+YyNeNifJGN
BhxlTRP4Xi8UlBBTRhW5mBnzziR3DcGsIyD5WtRi/Cb5OSjsk4H64vOgdyxj+NWg
HG87kb/lf7eyhSUMBg5QPrSqeE9lfULORwU03Yd3DiJcKdH6xU9qgPWfkd/VNAFb
owYwwpWVV3Sb9rd9NPY+QfqLCUgdpYx0fwR2vZUoJwI0PkWHCt4NN8rVwQnm65bs
kZf2i2aSv5LCICwQ7aJFClsPxVCybvKuiimE20XKWqq/4BpXd2w/ENndYpFFT+3s
/X9b6dAlc8Jr7ydGXbTsSMlz8PFOeSgszGmqTiGpXpL6cIqzDNBfo6M82xXbGCBz
FlxZg2uwwm2hMv11b2UX6wqMplgSiI4hAL193tQrqhIh+qEog9880NsnzrXpwkAC
7fbd76FKPI2fi+lBZonf2S4sm1kEAbQBoYSCNs5aVz+z0sDbF+19AoJAROSGXMVf
z/NEqC7dEBTKd0xSD4jj4ialZ+WXGEEURgh2osesG627YUhNQa0v8Uv1xQbUv3QE
aOLwkDqeXyE5CrjVDOeAPZQnoL5Irvn3F2CTh296KSwpMYVW5lEWIH15ATMeT7n3
cUUYRH17BC2hQ5YIC5I1RsUO71cdFG/d7Y4Cuyg+pN//G9F3FPZNRaS2K0N3faUL
7KBVIJulim+CFl5CRSqCbd5vsiWteAFMRIdVX6AGhZH4jn/LzwEms/NpzYj7eqfy
Zj23eN8u7w4oepw2s9sRg4dq57T4EmfkkYJyUh5xhnEjXeNy53UQAulIg8XDukS/
BwB3qlAMUEsIy2EgARbViCBWvhViS/EXCsc8X735LMke/RcTJwHJTft8fT8J1RGZ
ZaxRf8dbRvg4FFIRr90pW2htqIibB6T//9xHcxC6GX7IKYnuCUPe02gXvcyWq7LN
gSeZ+FigI1ob4nrlhQpFnx0FVlAHcWOX4gVBj/9ZgNwZuQQ+g8Kt3Hmk+1BiTU6M
YAKmvYskooRhyIz3H23t86SGr+fxly4LtxNSTQxUAxhHOrZY66oxj+YKwKhJyfpr
ObQ8fOEzbOFBPtAUpksWvKmDqOGTGkmqQSVe/Z4ja3sO6ME3spVTwF81FVdG/xTu
tjj+paE3f6kjcTjmrhdL4bRs2Qxs82fTaRvufERM6sPOtiBJzw9EIz2vsLEtN3Zt
mG3fkacNxHow8fhtKplnbC7KkkO11022xt9sPAKYs8hggDNr9d3qVE40Yj9+N7Bn
h/I831P0nir1m8+fi7cHuRXz1ElmgrnYFiOaxr123vQrJXMvG5Bm205rL5MuGjuv
k0++894OZT8BfhzENwcsUSjDXJGUFczGNoKa38BlS7DLwBjuvm31QBTcBpOgwg92
jDJn6X9W6nhaONV4pH07mSvwaYwGNUocZO5owPEO5F0Jt4Q6rrhROPeSrF7OarcT
gxJ7lOJeIQfJJlTutLqm01F3kWVX71nRPMYocBJ3rpxyi1nbmbCIS2i/QejUYlG1
ew/eoPIV8VFkrPqGaf9ueRunEccxRVlCRDp+Gii6VSK114omege6Tg6kgbPHAbxe
sDhb8HD2JZbm2XHPsB+TCGhTdzME45ibIquufB2NgQpAupjIIHao0dM5IFrCC/Ui
bNgj1W2jemdIr5obt7iz/lP2Rr9HQ/T/Wajv5fHnvcZnEo11BJOx60ryIUfDUQn3
lLfxphZg9JKzztisJ/EKrhkTwE7oszGdq79sHCqd62VcShz16shtkFwO2N1Wr4p7
ZAai1O0KOkWj6NO5LgAUMR+lXFwnKlafvDoX5bkudEGkFXYh1WKc/r4B3PdbhVVB
xmpLU+FQXnrutX7j7QcyNcFxGJPlmWcjaGqhHLe2Re/AaBWj6Qcjk6JtfxYlXJ1W
xvBBA1o82ZJyysvwHMMIPiA7g4syKuAVxGcVonuP8ahMLHL4pG4L8k04k2DMhzf5
Fue/2Ko/5VybjZrbIVt5NE4kfOFaeQNVFQNje0oUqLkTbOeBx7SKIUJ14tSiiS1P
5zVKxm7MIDmnrlrL1gRiVQCoY4tDdXm7Xsu7pI/xL0yLXr6Imn4XKMvY5X4j/wSW
oJ9a3m6qQBsWEAAgRV9s+ZYWf4dOLL6xaSP7YJY8d4ZY9ZB4Mh0gnh0CawDqfTvc
RbxAm4ipqzVgYweTQe834W7KbBnw0C0+u/E9rQ0QNB7SqgEOJpLgjs7l2FcD093X
8z9U/nFJ1aM7FMf5Nh0ww9V6l9HERma9AVQr+wdPPbry346e8dFPODfsfJe2woCB
xqhZ9Wl/SrLPSgmsZhrGTKihq/dmzx5hlEjIlsMVv2nIRCWA6mKpacML9HzLsX2E
oZKiX61DNdwuf65Evnt71Wa+XrjVS4u3prn1Wnq1DgbScBiklyjeR8p8DHmYwQcR
3N4VCU0dSKE0N6hmLVgSFzKpYeG/cM0KcOXGe3oufPyyiIWALFPneHr8vYG0VhWj
ZUIZhDH7FcV5e08/DUkNtBge+jAqX9p4nwJeFYagrfBuPVhsrrUdFVlInB+j8Rsz
3xQ8OY4s6K57eL137ZK4CkOGL+Tsr/+USOG+LxaVGMjOycxxL7mOI8gL2AUwloKp
jBzqPI6FCbqrrUZGBNkLNTPQJ8rMoajerZRlV+C/ckkZQM0+VjbWsTngfKTYZUXg
0duq9Yme0SrvTPSiR9hVYSWfpzVkeYgrptdzWKbhQ5Huyb1YTy5dcRMEhu2IQbCN
8Us835AaXU2hspICmfif+2ihaQ2uFTOB4wh/snAcQtXZR4foM46P0cTqXU44rRnn
EBBMLdWRFlYBnw8PE5zEsY8u9K81N75svKKNI8lyTaHNtIQWCDyHMrdDOGtDaLiO
uCFaWL3K7M1Wa8pPbr6ZFsCOL9cAhomSb2M8zZzAld3XVNF1XUNfjTUqrIEsDF3m
btNugyvLXD1oUdwME95cgiwXZ0900fnCvFe97IOR2KgBm3GMkYCbhpipBgq/ooV+
IMVq4v3k1UPodEWBD7VprjtzIGXF5F848sV0DR4OnKyItKWz+0t35ztCApZtPrbL
IqZpwpmzbulzDB4+gpTBxwe7+A0ku6/A64QSVJdS8KeCTkwGlQlPOmGCTuZLXEPd
bYMQAWJnsAdv1ss5ll5dy2a/zCUKou3YmYuFT+i75Vc05gJpe6i0E8b2LVynIN8o
pwpI04qszpbVBjGTqzSAT8ZwUZfuYSTtbx8Cr5Gs5PLuh/dOrssUFhjeZ9zR4yck
OczAM0dbfMCWoME73rrVKqbUyuX5LZsQ64CbKRics+7+t/JeM3y8lpGxDl8TdlG5
8VQ+XS3wjc/LPiwk/MoL6euP6ryI6Po5h5djjjFx9jPezTjmU/TzYZEbRg910iXh
C1L5wvIKC88StN70Ap1FS7jVaH1biS//nFzMzA/1/Bo08rRSuWamwy9K7p4wCUNk
VcEPuyr8IU9bXaj7DxnzH604nEP6QyOE4juUVxTKcBWP3vHbsXD1QP3X7Vo/ysct
9tzMESu7c02N9zxp/lOf/0P9U2sUQvx5fgoDWM9Rc1QACOAjkoLGKlhizusU1Vgo
2fU+7UvyiEk8amBRZvU659FHzrGhXPfV/jCqMBrPEKW+KbhmT6pH3CY3K7LboorL
6Fh3nORgVAMim7wbt0SliyXQG79KxEuwwYp2O+ULSdiuF/kY05AMxSV5aD752vt0
COHfcB8A8vRRKBJep/OikJE/rEQBJ8NGBYK9LWYZwwBkYyb5ht0m82KBnbkapBZh
CcXplf39R3v6JINuBSJ/lFmMNu+hnE5FCNYJ0ebRtKmlpMJk6wMblxQhcQhdIDAd
JzgKLihXBCT3EOQ57j25CMavapeauW+CgKaECBJgPgrVLwxZQCYwDvHTrWaPQVkL
XA0UZR4DNDmgr19RJqdr00ZeiRi6LLAQrAE9nRxjtu7ft7HtMU7qTtTvOveSxhHO
dJjPuHw3e+ta1PBEQb7xtr1OX9ojYU8WBsNE+X1aEkK01CV2MBHrHSPctZVc2LnZ
PE0UY4I1Rh4Sgj+ixXVYE+bjlqz/Rd2nRZiuqktzHf4rXBd8L9AP57b+ullpul7/
A7F+61LwJeNW8MyZnx9pK2OxECXbs1Z1GIr+nw44EzoZR9k/kL0hf+6olJrdDXTT
xeiZMaEjWDdwCwdyiwaF0hBle2zc6XjA/CD3ToPvg+g1DG7mXx9BdFS7amJUlD7V
Y2uPYTovh623oCUybStjlzkvhwmeermKH1mq62CBhR4S05p/OgfzJgiwnDEPDA+t
kduNx5Q0g5bvYBmwFrrOXoxyghcz4FrH557o0ul30mi//E3AT1Kxr8jxrlmH3SRj
l98ccQaA77a0+KvGC9OiKtvqPu+lac5Q0G75yCrGUsG242KAt6WREvHoFgxTh1rk
8AouuZlnhUYVI7orKqFsT85icjQ2PbKaKGSQq2Pp/rz4B9BBkrexqYtFZM90jMo0
QfGTBMuQzgQhMuYweU566CdNtMOw7AFD9fgc58GtyUKKg0WihF5ime+aSsDx0dyO
AKB/2O02l0vMWbxMajhiWGiThp6iKqRD21odhDB0mGzSzuG3nGuZ2xWBRb2KeFRP
JE3Oi/3fSRlWqytLZEG9JjePM7iMqIlB8XcRmH7adp5Rmyv48CT+FQ+wEp5xcwU1
Tsp4Q1X5GVJVnFvSoNGE8ZipwNd1YLouNoFbTp31Gd3brmcK+/1i1s5Wwcx8rkQP
fUjrNyc4IyBgw/uv89bMPp/TldvYzmXrkctiNaYn+xd1/qUTYV3Nu5ZEcEGUeXNl
kyoMkySmVQpglZrKQE1kqpZUH45kJy6pWXndZa9eF6zFr24pVMFtRUCw86qWoRlr
ORJniU7bTroiWvREf3dGiMhksIxp/BWgPnm4rHSXvr+4l0dqicKr8OtfbIuy5IQs
+R2MJxYCJUjDZeQbaAeuDJjPHaOQ7VMeUP3Fk5vafq7ZWK5mhyuyebb5aOIcSehe
3QjxfTddpFu4GSa0m5Vn622ZJMJbSoqyOalx7vjs/Kly0Hr9LWmBVOKAXxaxFeYv
yKQkxWAnnOF0jBw5CWO+IKH7jtya4b/6/M2MAB3nhFhqcsYe1sEBswvT/UpKnJHA
jQjnN6VKT6WKPgsHWhA/+9qF+cf57vc1+gGb8qCVlgAPpZJAR1fiNDOjT0XCAmwY
OS6NXVh0MXhBBiepDtFugyZmeQ6YnbZJN0h7yRT7GMGkibsIwshkmHu/8Lwj7gT2
g9jcfM+2jCDMVeBffUxd8maoClH/S/VJWambJPX6rdbBnPtWcxft1vzA+PK4SQrh
xUJbr+6rJrdaUxgZ3302VELi+/d0HQGMUFpG9MXeIVJekpAhSVOS0UcJwQvQfXnc
yCvAWhxC9dJ617RsemoDsqtHwG9/BJ6KS5Mmhp5x8BrVTFzHdyog+QkCkNx4PVm2
JO7JURmvrs/VvtR8naj9G+uwQlPcaMfAL9i/MsRP4DMwtsDGtTNAXd8+WDbaMY/A
4toPxxic7gpNUlRE7n9Ye6YQxzb006R1BdaSiRFLPVWZztgnQSpKdA8J+8zyMEbr
JEZlcf481n9f11NjMcgDCmasKwZVsQnoxkLaJQ86gzwH7SuAwZt/RL1aB+kF8PG5
E/N2F9hSKUENT/MI9A93prHNcHmI2a8NAtA4d/mXSI+ptyJ+6ytE2gdc2YIlXwSR
y9bJDPLJWaOILsgjzvVDLpMjN596TMzRQz1s6N6SsJRWGEiGoXy4R6FdGVtOeo/L
Un+e9jaQ5cbtRIFHZKgy9gqN6chaMg58NdF4dt79dPLTTidvbq8oRp2py8Kmxj59
hpYVwTiS3h1kJb6n4L/sWUUJgT06Vm4+F3BHXNklC9mkUQ6z9y+vbVnAAhVZ5PWR
mBztJ05Lm2Xl0mYptvHKbNAD5OLQ+lr/GrW0E5b1hu7O6VuvaKDdz06ijJJx4ojo
tKdJVpSIjc/FVk+QS4olxwVZB1wcY4OJpEn5fcK30K4R7fTHxxTNzHJW0IvqsyRe
8bPzYQkOF/BwymXDuP8ddGSaZZi60o+MlZYNFkLGXgGb3Wpcl4NXXrXU5e+tZPHT
2Rp+ODxO7Newbxrvpp60xqbyTO/uWtnU5yRQt5UaMzWEKXh3+qJHQrTeYEfhKkQ6
XrK5etnGIs4eg4kdTXLYTG3Ra9n5GUW3fqqr4c6ZC+u4w3oxbv4cCN43M8/Q77jK
46ohUpehu3o5C15NfbhLD6jhQdQl8yubZTKd0kqbriYV3OwdV2rIl6pnpMBIozMD
8znu8wPM4u7w/kCZDxZrlG9vFcyYOa3CNwFkDfqW8wpHHaHqcrOvsXAxtF20+xzC
TgEi8M5JvVbM5lZt1Mo3toB3SeoVh11QN/h6Th7BO/5ZD0NS8a9mw6jgseu2PnTg
mtdUhYRx62HrViFPX20nNPKxaoc0Hiz9h3v0eMQzK2W8FUk4qe+tm31zWWEN6r0V
zt0o6j7FMewzwhO704Ylf3mj1s6PIyh87EYPyDdtLnydr/3OMNeYsPtf8x1ALUO3
vX5Eva5c8N/yQHRl279PVAgkN1UK2YHHDqBmIG7PX0bBTMwIQtkVEBAl8oBuKeS4
OztiWAOygF7SMTC6Dv2UX+pNT+LA7RaQdkHRCJN5KO1GkdsV8BjNoRTIh2woJUnS
ptmWSxwxW5lWODmEbfaHZxCKFzP4O5AaASVyN7Il3kXIaK72hn+9kBCOmhRosPdc
JoxlZ467pSrVddk0etOSMj0xkwhIkIXtSPCQ2xsQImtaMGPppScWZV9iVbjIy4f2
O6uFWoOAr3/XY0+72wqzNMRbQQOGzkowUcB80eg2JOLhGwbcQ60zTXEaegswYrbT
uMF82gNSoMpuRuQ2NaBwtkwJQ2IQ0TIuuE/wfm7MUVS4l/AG1nSYP3kPot4EJuGO
ZuTMvZkscvhchoXq0TGThBM6TmR5swnQYX1hEzOsAke2bT16hU0XvOkLyohIltXE
+7RzKCqPYZeWG+TQH+3lZQ2Ef6wUqioETixOwk7Dou5vwOiZc0KBNuyAxgu/9McV
o3d8+Sys25oUxEtNN4lJcQQhMFwUGlEF9zyTD0aM3vY+bHbMqywecbb1cjtFMr/i
O4cEA/hVqa5gm+MkK0K5icsbNuDsmwlE/7RnD3WUT8s9zu7juewpd7y0qntsmCr+
kEi1wPaI37XPThnX0cpWaD/MYUurnu2d7pYUrG19GlYfjR0b91fgDTzG2IMyz4bH
wmpSlT+9bzUTi/4npUVs8d+BgOhQvUyB/rUPVbuILKmKmfMsv4H7q1pV0Cdi+W4R
pK2N2E0TW/2aRHT9aiQ66j5Mp0gwBXOUISRy/DtcGYH3kx9JGPcEXeelMpQr40Ve
lx2K4yg97DIV5fYBvijAkGyKXHFlxvbhieBK7ZutFLVPcbhrdo1UBQhA/p5uraxe
AT4S5ZZ5C4SMoSTG5lysNFyhBipnZCzrwfUx0idpJBeAjJYYX+wb9TlX37xlTxQc
GF6QJgQJjoczBQf9R5j8Hq6oS+ACgMHS6Koa1zPFgVTkZm6Gtw6ysD/TFIWGYn41
9s/UiWHXwpiUmZ5/wMc1GDhT+nJRvNaPK6cmLdBG+ZG/Za79Ob596rXkpsV5ghqN
XPyqID4zyhitNJDJXwa+KhYqWdWJCrvJNjdYinn8DvBmQIZHXZ/CgMzAClc2sl+B
mrXHxUBuYLa1nQ36qi97diW9E9bB/Wkaq+2n0oGMzMU5bKhon1OUxYLWeGpuZp2y
Y5yUB/QF4S+5UidTezANCqg5kNRjPc0GmTt5bc+2bBf5vd8xTk6TPjaEwf/xJxSl
sXvaGaEcJB4Zubaz4xGGOkpXvaDNr5smn5fPK4bk2QsMr8WGROKUTVIx++Wzh7+M
FVnHWZdKebiGTLb+4Mu8fQNzIKElWP2BjBfGUuFsIXaDMeCxdv1U/YDLHxH4tPGK
8XBVycVptND1jUt4HfiE+VJH5aBWuf6dLSOEVGRbC0BmZfP59OZwg5oIUHQFLqiM
0Sdir5xst7CA14MFLSTlSa0CxRDWx64mPhp+4R0wmHEhWFkOJ1Cj2y/SMPp0GvLC
7eiGm4u0v6iFip+cFHwA7pRJCS1n9PzHszRruNipFlU5Ym6pgRjcQc5nrBinx9xh
WR1PTZwpgc2fCu/YiLw/Fu7hDjOv/OvsO/RqhQ2lkMdsWbG//h7G30+sgtKr+ghS
L1D34gr4ZnLEMV2qM+dhp+AJfm3C7QnTukNAW+vR1Q6gBoNlwyns27cOxEyz8gN1
BNFLEdYCmb5EUBdCQQoFFcJWh3JD0xsLkW2M6LZjxfyjskIdgggW3KdGBmh0Qmn7
qXu522vnWWg3CTP2vunKgyLXqvo0zb43NcaE/gbp4PAwd6Sep+3A7orYaA7qxj9C
HDrU0s1L3EywtTLZ9exiUezI1e4nidInCxQHh6GQyq5PW9fX9lfgojoi3cb3eAHU
nGTWpA5mX5vAZYyJ2M+6nCstk2tcgTKQBeaUylY/AADkePhEsGFKerbvd0ggRSiw
LFYjQq1Lu+/oPmm4Zxob1DLEwKVTTi83mQrkM22yfxIKnjOR7hgU/hp7ugOJE9pE
cAzzwCFA/DEp8dnmB3jJhIPVB14yAGAXNRVNrnbGTOSbErO4/QUcF+jphQ6mKGQE
3oVIEA36VF419rEYPLqZkqGphqGJSij6s9WztEH/J5w6Fj9/F4FmbZANme1NDZGf
/ssTiV+xvL3OnYJQd7QH0293ZGsBy+D7DzW34M0yWk17wIiYqqqpIHezsMnmpz7H
XCtM5lOjo6o1Q+hYJA10fX0qi/VsJq7i5rr1uAihcRFfj7CUQ4r01loc58K2EDI/
GYdoUet3UVas+o5kAw1yAqXs+TXrgTSf1yqZ2hC6dltg1rQcM0cBEPaD2yHFJsvk
rBjxmAVwx/baB6diVm24Ho1LuzOgNZSZl+TE9XRvxaRGJSKLDWbKhlgTFI2PgJ94
Rxlg2ehTGAsGc2cmDmhLUJra9hO2GL2QuxCkKaMJayiTnyY3f1QXx5z9RJSBRUgc
hDHP41wKc+kSMz7vlaecyfUTBPdmYvQqoESigRDZzBDJk2c8N1akEA+3VI9ZHl+K
Yo27OHroXyVtA2wjyhP6l2cF2HnkF8reeJj7XeSstqVR40VEd8Qt/38YRYhjWc7Y
I+U5SxJM4yVrnBhi0l0vNl3bkiMjLYWsGBhCJWYYBJyA2F96I9mX7iWewZ0OjoI/
C9R4VMSmRfoEXibFxZoQE5JDbrncFM0Dj46msD3frAroRhQaufE7sX0OJGSRAfq2
oITshJm+H+IwTBoeM3FxE9P0jCTqJ22vwzufW+UChu2Ln0Jm8guU2Q5xN4QIwU7W
`pragma protect end_protected
