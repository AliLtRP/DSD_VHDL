// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:03 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
f6ZKZiPDG8iExl4DAVwTZED5vL2gzs8es8xMhvKRHt4nzgN9KP/CyoMugzuwBMid
qK0T3WiRqnwTxq/MZJ9h3mxARrM4TxqFc9P3qj6TJEetXEdgx9vB9Nf9suWK1hP1
eJH/oUbyGDqASEVJmD7rsVl1HUgXJasY9rnrF0YtcSs=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 185408)
GZsu5w7KDNO3Dy8fwKne2ZUEVe8WFh5mbKlT0VmTNdZJswd0r42am7q8eItZpRgZ
sTYZYLWKQkIqorjTYJ992FOwgYPN8TTsBT/dkPh81qRd1fS3AOcLulXEI8gEufV2
BrI6El/XRwpHmfkeNfZRb29Gi+DtSmq25Oy3QfBCqIlRe1NTjFUu9eFU/Co1oT7q
LWGPqI3QYeBR4kDWnZ/K3Z2u7izSIai6rBi6Mkd9qTCciBSkUMFfzXeobXVH70jA
jebeGA+WP78GtWwWOaS2nc6KTqBcqg3yqirR5du5nduC49ZEuEBqni20OHOCQGuH
zTpzn0xfNbORLYIgq3BcVpEj2yxN7+57vehz+RXjp/Q1SWzVWKmAnyXGM4tA/J4c
IpaZ+jd/nAXsrcqZFcCLUxczKT1jFjXqvJ3sSpPz4t1D7yGjdCDNqGir5Rn0Xx5x
VAl01PnkW/B7MEwwpgmfvrqhLepKPZT2b7oM720+m0I7YCHkmwYjgX9ES5M048Wg
8ElIsKji1+ZlSihpJSmYurALEttOEMczQzu0XAVsA/lZm8FpUxDBK5g+v83brBKY
OOtFUgI5TOsb4e7ZB0DdlpAFL9Ds0EMTPULOKgenGABokMR7AOp20bXLCfvoyejV
eXaSgI3WcKfLYa7kmRMVdv3UPZBIrsXWZzLBC8dr/U0MQUH8v7EEGI6VJESX3zn8
cUCMMWC2JqjJVAJpvnjn0TApPtOr5BrjsNA1MjHvAZvIJSh00ZLhZKGOkA1yjUtA
rpVHfG2d4kSPExpbYz91hL00zb0KjZYE12cPKSEeqeloyDlJOCBJB98S3OkaLDMY
hu05edu+a/ZveRuqXKTGfGCMnMb/gCpuLqOJSlTbmmiwj5gqN1nD20zR9KsUDReT
RvB87P29z8qU6jAM2v9Uxz0o0Xxios1pgx1JHWIJc7dGiefpVjr/Iu6ZRBGxLMz1
iWu8/JnM5rUFfHP/KOpRcXcTodK6DxQsxE4vXo0zi5+Vj5uUbMcag1ueCbS3RCM9
QbC1hb1RW86i3ehu9DgdkWGYGbsms6flEsxASghixPrKGXRsIYScr4gSJ0EhRQgQ
PO05BPxGpk1d23z8pfTQvm2t8dtEVdNgjgAK+fvLRkOp0kUuSYAez2sXf3GnO8Ly
I4MYf/bxLZ9UtTmz7KhTeAG+rLXgaDH0BFvsjTcHfGRZw3lNWTSTcPXu3dd8BqCa
+LbnMYNBYWAtdI49Mv/pjQZ5KhSMu5fltSbCISdc/Xgpf5nF/YXT+KeHMinWSG2+
wZhFvtvtjhtY1SbHifZxUXlN3TgsQXzwnMKzFhLLq39orA4rkk5eUBV9tRRTagvx
ThoPvgkb2OqyCAwHC+VD8t8s29xmFs9xzvJzxpU4KYGp/vFrCeN6TXIsTaOhCZMZ
deeeUY58KsSKvAVqaB2SGzCf37Vgkr7WLDMwbn2ieqd7dtKQok2MB5BCNfHkGBAb
nmQ4p4F0t0eT4VAF74OBf0QqZBFSC2/FaZ0aYNm/nvVH+kgR9zFn8buHiBc1FJZ6
DoEmgN7S/SVx1VxHKUoGICxni7xmMHGDtfSF/uSQI8rEzeOPjqQTibwNLlBupQvh
28AXY2XuAe37znV0SOtzrQqbhhOAJs2Q8i56T6+H/0nFyb5XD78bmkvRetjC41bX
Nur2QWh+UdNqbw9icqlRiKSyW2nterZpcleJlc4Dhkjh5DuIU+N++HgcHGWzhM2K
bcP/cQ9Nn+I5CFnvgU4lVUgi7jN38uQQnpTCk8fzEf+E+iNzWQii9aD2Lb+6ZD/M
2E04R9fFCngCX293f7wxXlxVcBpfNyHbNAbXQaAmXzPtUANY6ZUcb5UJzV5anRd1
eOdL+LssjYNElFdJLSnNRFxYtOcJhVSRdMZQCa1BqiWnv3L8BUlx52iaePy+0w1X
m0+R+TsE5EFD8uN+shRDC1aLGlXscYoLRqHWhWA8eTsnqgp5Tpj7Ksn2J+dxGUbS
8oYOsyV9XdwSEGTcQGkqK6ZwQNkcCeaUrd3LWSEJHGK3zld/C3FDpue9NFhclYMY
lV3SK9y2MA5JIj/qSepvppZrEMpeXzcRBfoO/brQPnc9W4IS0Iv9jQIqLJ6KP7qR
tVlCFXRwg4qVafed4UnDUsRKz3QuSEvUzp7jkesoF9Q+txJj/Wf3t58UCKFZ4XBX
al3x0wGBGUGqSXsP6m16yQo48IcKfc4CMfP/wK06lQfFUhpXV8RXiUGjkYpRWJjS
52ex2GQ/aY2aMwUd42VAgL5aTU3ZG1G9+VZDm0E5vLVJySds4mDOLeC15xR//xz9
d9hbr5aWCJ+gKK00HAGfUE/2gSCCTchBuAGfyJDo+Nr/6Y7wcntQh1YE3paS0m9m
UN8LNNRWwOjo+nx+4vS16u/lN1r8RDbttf1fD/tw5tIJMG+tMQ84Y4V5avttS7yu
FaGeRKwKjym8Oq/t6npgW85GUIxsmGR6a/AXB6b1kyf+9kpfAfpZ2fLp97NlyRK0
cQ+zDOORbFa5txmrGc8WowmX7HM+skOoYf9O6nwUVylYLJWYf50CzfxGzhUA0khP
zb+aF4XWV0+Ng3nVCit+yav6hFIdhHh9Iur26QkKbJKyEnqBfRLs+h/DINzl4O8M
PSfBhADXvfHS9DV5VYjRWHxNwZbvlLzYApMTarX6R6FxlB9Te9yUT0fKI7Uwc8d1
7dLS0cUilyPPcxfVcodvYTBDOxg092dA2wq2PPs0l0DUe64Kh2JorR5zJ75a+5ci
l5LqrsnFpC6d83IknkGjqSyfqyps+xEbcPQvwGcBZJSvqSmZu8sTAntPpv89JKyH
YPf33+mrM2sQXAiwYs8FmKi/moyf9JkiYK0e8JdwjnnN9Ez/WodaZbUgrHHXPhmK
5GY9nGNr9q0GVF39FeSThOFA7PnrjlZUqqgdQSdu5CfVCK2DOqTvyGoQLvWDu8I5
h3kmQ94bLHgz5xwR2vACAdePT2x1aXG73njnpWO8vJ0YkYPh+LGhQEsLpNDMe/eA
3uY6IUU7xhHDBg/jLzvGMb5dj2lWF33jivMEoggb/3hQ/FWPdReFAeBxXQm5SX3s
g9AxMQi1WSmPCB4VSi2Ux52YRDDgcSvAbycfbqz6BvzKZksNCZgmG2xXEBW0uxAa
C7eLGpnAk+JH42o/QO3z9uc9ifFe1ShkzQd/vYyNmUHk8i9aHV2QtnoTdas4GL3S
fbT+msUsGEMsH+1XyPiClv/EUz1pbXk9nbK8FWWenRSx6MBxaEVtJ5h0XAaXumDK
kMUiwb3VSxWbfk76vRe3Df+lL9snACRiLHSHOLVfeM9umjR8LoA4jqbEVFKSZHjW
GWjeRvwY4I8yo1JzMeiz/JaDZukuhM4MilYUyb8UkaQgn6SGQ6I82yH26SMFiUst
0NVWCAG91Jpnw1q0MKQbONFBqo1o6KlwagnYwyiGXRXtiQSR4tBLifX7IPX/sXeO
+68krrDJP7plSd02LEjHnegaj886BnGUO399oFsKIRop8sEc0/XUOqC/LwgkGaza
9RR/G6P4jDuVN/00iWwZFxtIgvzyQDQuCTWOKtP05VQfVmWLtWiuiH9PHKBAAru3
xSLF3py7hHjT20w4szJX0Egc1KTS+4qecfKcEURxBvATym+jK+Wz9z22OAj4iKet
gYoaOD7hfJO3JOvxSUmyOZ0fDIHJ8jnG9+sqrHa2xx9ShuM++2T+5W3ptTMkeGLV
+xFHPPbdOMXpq3ero29yakbz82AGWA03KEURRKZBvXRWZAGM7HqNN/NbLhqddl9X
o643ci90lxI8z7QIGXpF5ODh9zYPzUewKucuUitpTZYVSN3nuCZ5pv4t2e8VMTnk
oqmonibsL0iS/faFgQ5gn/y6oleEejBIPwwxMJcey/BmeMSTd8om/UYXwHH17nlj
kyaCDVv5Zq0P5uRMOTPGosj+1+LhjrOIdxTGF2ldrDmxm7/KdvuxsWFyf6a/PwsH
pz7zeYj7CxNpA23UI4dTD6D6SJhifYInlZ91uQ4mBKmsQpLzLjAf8JdW84BXVA1H
NBqnfh1iu5P/Er27LgY5grWr5W7wgS5mIxcqBHQKMh6DQZatCD/tFdqwoErlAwA/
Pqr1tLjQBQ91grMz6L/uk/1e+9kuDvu/QT9HvAS29PACqxHmOMCWjqHqR8AFu9yY
zSoCwFkGYQ9l6uX1z9te9JhXUMYbEqMWQLtv9oX7UpBq4vMuULefC9a0Vw4kakE4
kizXH7xKd2AdvrAv8Q5OfI9AetxxUN4wmmD57F6s0D7yEWIHomSZgJ9RuhQjsLAV
Xtgxj9pIIW3LeYUJiz5LjmmwRRYplMzVnLYyvWGuDYOMG19wySFCn24f+049+OTQ
/oHNKGYspNxNGQMNElNDZk/4J4MZpoSAvGJ3MA7cuua7gRgxqS+vO7rDf/OvUWRr
JuOG4KXRW0OpOn+B1NAdQNFbfn+8ID5Vk7T7cLS82olpV3RsEKE/9ZvjXTKKeHuY
mZqeA+vMSUGOo2IPp/I4wezOULp9gDDBteKzLwvCLu8681ZZ9TtLhYV9jShGh2Aq
13W3tERc7zh3tzUTivOhZqgCyjLYFuzhwig1NaktZMklN9Ic9siHbBtHrvNIcPw6
LNco6g2du2/kYdGBov6Lk7q4jaQ1K7NPMcmrf7fXpG228gtNq6AwgX8+hCjLYgaY
D7IOdK6qehuuEx4FzhIvRb2Gx+7jPsn6HQyhA+jNMlAGGvCxhmUmWljmsr4/PVEp
q9iqXNCdup5vyWssleClPZLB5HjwfjmfvBtZMJmKnSbGqilcqHDPKu6bVMculvwc
+rFXlWIuB7s5XcIAQW+Vzo1gwFJXn3Z5vucMzD4Hs2zsbWEQmydmN/jnRV5CCnRk
2I9SUbdAcGxtuutyhYvycEbiM0XugJMUJdYzgVxLuz3kgkMj9pkgsD/RtEz/j0//
JKkMrqnlywO2o6lnixb/y1CNdoToP96gwjaTefY7DRbed/cPlWhJ3DlVPqWkOLga
bE9OYmWPwjTLqOMrwKey4tNtgPsVjOtq+qjuNKqtLYaU4y3iotakT60sdb/RdSkr
m85H+cSF8N/ZcsPi2lQRQwVUKCb+l2dgeTQMeI2n4E0bCyxsnwgX/hGZfMjTYmYX
91seXMglhpmkdqF04f/Dwni3MvhbKwGyh67/zw6IMzun6ov9k/QDYH29bE8GBhi9
Y2Rb0lr14fxk1ySse9xiQqMHvZA0aOL1ix9DB5ktUNf+Cs8bhFT+AKsjq3sapF6A
87uhF9W4ymaaJPicelxPr6NERTb/CwtyHZyewt5f9G3OhhfguFwS4XFteu5YQ8fW
jfMTQrwbaN5E9GgNfLx86GNxIG1EwdrzJ0dDUyBJD4j0ka52TCY2UVkwbw0yAZlG
Wz8JeSL2EKHKLt0VVxUYTc/XBXUrbkzR3HB30raF+4TaJitT1kF9A5mQuejagPhm
DuQ+3Y2yUyUXNsZyHfsybfPsaRi6CLF2nDou/k/HPwuQtztiHb+5d9LBEb5x06KS
rRZEKZlX5vEKj8YA1a8OPp+CcnPzCiSq4B+pADdmLhkzpTVAqu03Q1hcKaLVgflK
5OwHCSddrV9dax0Z/GYgsu7A575OGpcqI4EEt7qmf7lj9Ke02TrmETulzO8F2yfw
YwIzSgEKSg0dldYhTFwpQD45d+RJ4f3U+2j89QrdaIiELtagVbaRoA1a2fxaatSJ
BSNdWXJ6vpXnsBN3MBIq3nfhyICiLi6yJgwEZAwyS/1Q7EHTv2t/ynTEexxxF362
0v7pds47fLbT7XDeswQS4NU4zUHO1N3mslsrprv42EA0bWRprjD71E1w+CtlfgYy
yUYsyzVuf6SiWRepVX0uGb8nqj30dlLf/ZljOi882DtLfaCvKuAlw6+X6VRC/isf
9tKaQKV/B45MoQcTI1YzWdNS+ToLUWKjUhN87a41Ivi5o9wf/kZh/uiqqHjHWeb6
mZQKjl/PCwvf63gmUaYH6++aYiBeQtjFbyoyszb7QyLCKQRyGFyti9Mi0/2e6FKo
XGsSjMc0+K1B1coxNe52kR2tZSjw0vyHeMhgYdNXyuWn+aJ/P/EkBzliyjd6EfGp
wWbCSF6H5ntDFs7jG0f3Ud7c5IkPeDbaUUPXPB7YrKG6EFYFHbe1BdD4u02fqG6J
B9ka88bjYFEAePFzjYk/avQB9oEmSYB3awK5PQC1diEmXe3NcQJ1rNB/Ol6d/PEy
OxwyDV4wV5f7Ych2FyMFfSbkqPocP5WChwtmV98lSa3pVVNcUDAUoWY/I95G+uD6
YVo2edauDCfwIumM8PBATbI+E9w+d8cQ3pNG4uJO9o5nKTs8tK3YsyHpm79YrLgG
rQqko8d3IYGACohCotfTxx5UCRx1/4kI5VT6d6HlMwCIy0mUoxbgceoCSUjab6R+
TZz2koUH00TvznBp9NOO6EDamG9eXPhPtOCrmB6RsBGo1LV03tGA2a2Ov6vQFqy6
uR9dJWwTYiUR0PJtQ2VTzkzLlCTXZ5Gui7xEp053pmUeiDowxCW4vqLvtGXnr9c/
Dn3zgt992+1PWuCKQ96W3bHN0apwUFC4AcQ/xHK9gF/+Mw9PaYGksQ2Gy3VmMTWx
a0aR8GsIqZ4VPhS6dB+iPfZt8l7tR0cb3rzwk8Jjs5QaenGJuk06ZrUQsnvrO2Jy
KFkTch16WttKmveFRzRKtsRjEU0whQWyF2gUUSuVwIPnwwnzYP1cGuyKeqa/4dSO
UyQ7lV1T30BYn+pKvr2BR152394+XrhriXGrBhrJdb6UrGqJdFw52mDSpEcUniu8
EvgY8+wljPdBqcH/O7XkM/NF5XcrQOZeC+r4w6lP+ydRR3Fp7GyzCofTwohLB8Pa
rJwgaZREUHAdzxnbg/D42/sxMzGkiqiHl6ftmwzTzzlAFFDD5eHetjDxvSG3oKw7
PMkpUaMzp8NwpnsjY09Fq6IVBC3Hqiw3V4QxkZXyK6i9PervZfu7UwjgqQd2+myM
fl1vNVr5BMq5+VB5nNscHTMpW2wriMndB4OWDtAiLSbpWjgH5rIlR+ieEK6si78N
SZRsTIHq+SsMX5V7mOhpQvmbBMQLmfg64CWx3W3x0O5VhVxeoIILsyDTBWtKBrAT
PFVkGUhwB2jeA16PigqlZNwpuO4uH9tLF4ijUyToHRu2tWAPBuAFNZKACq2ic7mZ
e4M1WzG/F5YJFo5JJzBhPeLUiAuk/8Y42l2gC8V+YlXZkNaK1Zl6T8VzDbNiDUsg
82WD4UwW43LBxpcJgE+WkqSJfJfg8yvh7c+gFD2+yUCAWrtYcGK7u4s5IrLTEIfa
wyUsJCQOV2dbo7WHLQFc1jWkQuJ4YQHdwFlT8J9mLpyju9Szj9BKqo6cRLIWZzJZ
urB13j9dwG1x5/cRhCWo+tzv8rTw0AvmYtL3KvEqg2e0YczNtSIA/kAcQ9p6gDye
5RMYX9xfkDVmtX/x3isz4FEjusCBXphfKrahSczderYLRBGAnwTeaRB12CnDTvgO
6UX+t8ygT1QxLfppcjhQ5E3/OjREwHt/0tSzHHp6WKn2GZwKIi+TGjnuxxuGzhua
jW7NgqyhlbEAVfpqac5qqa3cnmjD3fGd8OtrzgAECbmH0ZUfc3huJVcUCGVaP2E4
1VM6xf/rldFSio8bKvUPqz041kmBT+HN4dsOiDW16yo2YJIpgP41l1TFfnPZHwuj
06DH/b06dN21y0bhSvHlxxKkInAuAL67Rx0vEnIkb8Mb2UVOlUSmz74WJOZZFRRd
DiGIo/3J1RzWwIaH+4Vv3W3ZqpUYEuUaITPaOL6gKsmapZfk1pe38SnyeFL5ZhjN
cPr6CtV7VeT0+PU04APiHRzAqIM5UMAXBYHEWdK8G4yl/alzhlV+ile6SXVh7OTc
OLr2OB6ozZvOehMEtdHWothIUVpgEsXjNEGjG8CWYhj0oG12PbYL7Mn5Fp78wJaz
gE7LqSgbT3NnfkuiyXtmfPbG83tF/7/FxKxHxmcx6SJdia7FG9XD5XYBsOunZETc
BCawFjLlJKWyUAn3nfwnzflBj3rJZsH2gIFX9ElJf1k5gOYAs7dps4B7nnmCVuXQ
FzdJBAVEk7g7NfYC4eEbX3d5qOqArKtsqCxjJtCglZroGJiBEfhYxpxXRx466rF6
j/a1ht0sLVTzjar94Ct0hX7ASiLG6+XoZ9FZTYWp8/TSKxftAXIEtszgV0/YGaZq
CLP9YUdcXmXa8W8wSV3xCgrLLsjNie/65aI2/21r7FWh6RGsOKRqjMAcMv7NxuYM
JXFgAe2P7Y8xNgJU7w/ryEjyK8xeWwyT19fo2AG0uF/TEQOgWkfiOMbAry7im+z4
oXc+OTnUWAN9Gl10NnYHc+i7DF2vSl+fLiyALX29U+CKGx+zhehXznS4AV9+XMRE
8r7vVl+Kxm2LDGhe8fapuGq74yK89K6YHy4SXHAnuqOYm20VUhTgH0FSk7FHCTsZ
iYief8MPdiY9SSpoCQdjNvKFd00/CKf5iCod2VGCOxLGinFY7PovyDLWsn/awhXI
5beBtWqHipW2Tc79wIQKOWHSU7gZEoptWLAyIorzLpwMmy/ilv6p5THAx0YKI4do
P8w6SzrK8X3UV/AdGU+iB8R7apBdOjmMZqL1GkwhL8/0KeRCHcuKyI4YVdlShYDZ
BrnPV1Fdw7hKC/94tubtLgkUUwQ5KMtWKtyLgjRuJInxEIVCAUyn4aT82tzxal4f
b5dh37UEKapH3r80xxLbd2pHm1H3OOWn9yWfTcxInlXKdSSQYawoVJHwXcG5gNL+
mCfPiw+7WQqv7Tb6Lk0gvvbtiLFWJplUCJtRGCNxiRshde1J5d7Sg/SK4IznwyCD
z40KGxw1u56MvIAsu22mVJ8Rm0/gWBJXwLfO7o3HqjWiVsdTeP+/UomHo/Ypxy2d
gdRqe0iQ7XlJf4/XywS7VMHAQn7R2wTzQEhhc6gTsRqaMQo5nc0hh6Mgt5oVI7wA
C1rwWs08K1QItcuExH0AlAUrggiNnyW+eeMb04So6ay6cWgix6D+sPPK9TdpSiDQ
7dFB5fa/EL9SZ1G3JF2RVQ6/3eAk1kcEsbMfwrYSKz0de0QRj24+mPP8g8nzYAvL
AfPhs+ydN7ARrkevVPaAu2wlZ9m3a1y6lU0tsCa1A8OUAZYDyxJP83ltwJtJhszk
WpEXWyi0zkRj//uVPrUOLZqAyNlol908BVl7TUx218mTCH3Fol+upsBdCfZd0wOY
K2oKxnOmgtshTJ6UfwmE5AeK2XnnQZ30Htq4d8h6R4ZlJAaboC12OAXK2DrpWvhY
9zdN0j375lkUNbcVsQPRllrjkF7H9mDtQiejL8oPJuLLYsWnc3BfwG6gX/jZdPpx
9OoG4BCb8ZH4ZlTm0jof3kMDTSaqekCyfI3dEYQ8q6gi6tUbwQkICB7QCMd61Owl
CLNuelFh4nIWFhADUdnAqSxNj9diVRlaE6lU0+AAHCVfHhPQxgHNxT9U0H/ughsK
bd9Ik0LH4Y0FAL0gbq3nz50OZc5ziQm0u7cbf2Cf67AFGl6VltsUSafCBV11CNY5
Cbn46A3hi0ooMncp8/PSs+ynsy6YytNfB3MJn3dbgg8kZi1DUD0Ug/rAXllfC6vF
BuVnX20Rx7ZneiZ2Q3/aLsMiA9aZVV3Iol3bKqGacl/w2EPzFZeUVW9ipbReiaUm
aJHWXsx5Qqex0zM5nAvLU10Um97KNxGftNs+VM6IrV9JjmqTW5gpSz4FRw9Rp1oT
ibDdWj0y3Obv+rLFYoMfEOmaX6l4Scu4WsG1F29MqGu5FauMz8z5sutVRvs+ibH6
/EohZYj6sPRR7on7gqfFuEuqaDotj9zv7Kl/NPRAw+G6AD8zNW1JHD0rrH+Qgg+4
nefv/umpv1jUrnKLAuWQelCGUsyOpIhV7EItzq261i2ifGg8EmQqJJ1ARQedpuVN
NYWvChfOWQYCCmOspuBDv6AXv6NigwD517DA0CMqGU4JWF3WxNRfWuW2/X8yTZmD
3WJ0ahf4vMVUpRbBeLBT8ZS+jlLdaZIgutK0CKnf3TldAslb7dFIEsXOSHd/Gg5N
1K9fPGvEUKVzFPUeFTiVxHpz+ghtYjQiHEah/0BoaIVLQMIbsOdXlkQL4D5MKTXV
SJwopfxMGIfJHWa3x+gp0pIR0OM82E1X+QQoEJZifpedrFvcNxc/nf27tIzJTFWW
2MfOrxl8c0XGiHo2eU8Fxuhqdms3vlCABX6x0cHBLv8GTgMbPCAbm5PbHqJYG/sF
cBPSV+VLQ3SP5eT3MlHlpZKqZaU2q5ANQ6xzveVKgbUK47CB7o9Ze1JmOQ2uOkKC
7HeNHqJCfg5+YMzjXFO6GriMM5xNdtKvoVN4ccMScPMM4WN4tjZv3rGb21/aQ0Kf
D+dReFI2iAtt1bDixpnNNxFsKKx/CG80YnHU24UsvixcIrP1VotWckuWhjAmAt/S
bgBuv1Zn5CECNBSTEqfmAl+a5+rm8S6fRVHFC0gsfYyAYy2enAgNmmKM1jOvRbL6
Rry3L4DLx0lBJR5y6EMeQvEjuYHy74pq2pfO+KTBX9jh4+lieWEEpxUaCTt3U+je
9kyyweSdstekH3ROoEKZJXfnTG8pJOURrHTBhxhI0YGPAcpGuILZG/1ZIcY2HBip
p/DyPWCV6vCfvvqqkKFUdZSyrU6h1DkPUESZy3r6NUR2PNEZJcbnjEygcEN1rfqQ
Mfd84Vl9vYT43zQF/zBUAakRowJk434DPytX9vl9SqoVpPlLqhjKbnGTKaK8b5CS
3W9PB3XIGkYV/CSO6wFDj9VP5+HiKbrnwySw8SbhX66S5bml1icFXk/WksT5jNtf
EQaHGd4uUx+kg1VSeZm3fotYLEgs0hOfiMfnTAhVcJmyCNrHxiARFy9Jqfu0NwZ4
31ffPNMxs56465sA7jU6+MTy1CnHk3JbsSIQAo8unuQWM8I7EIxh0RZ0GmnL7ZkX
G74A03lj84tmEity2FRzfzzZXNhW3782xQyp0o0DQvt50qYaOavwl+Xs97lxtHIO
3uO7WqWmfDUM+jURmZqVXSpShCzYyHuhi2Los9ZZ7bPo2eRKF0rSpbhvq6Wzrnal
QGlItHdpTS8/wdk/HvBA0WxB6KMGnhTjzGOTy9/oFVJAhRy94U46tFm7DpVpPeKC
mv8vau/lSkj8qP0GC0zERjL629fuJ5Dg8orj14XpOoxt0Ay9yGM77NXDCtU3XUby
6M6hSOmcGWNpjoKzb4O1rPJLPRtIUYyn9aXfdsaKWk8Z4XG0NvXIRRSd/Sfe10vO
GVFu6aG1Y2Jm8ljoE4+jDG5d2ejtPSLL2pI+rS2/qEiLLjCNOwU8fscZFGSiu5kE
x2Mu48KltQzfFJkhlgGtjHsTiLlSo1SE8pnYPKUs/U2Fe9a7KsjZTIZl7+rC6c0o
sQWqQdBbj9jP3tE734izdfBsfC2dyi0GMdNoIBqbeZoy/cpV23Cew+zmR4mwzaHG
DK1fXpnS3ZW2FYEVRN7+UsCPflWYzEZgRYOkaIpz6W2jnQlkSXDFgLS2AnCBMpiE
F1GRa6dmgdFtn8of2PihpR6etcuc4eKEgf4eI2xuJfThRXHV5Vz9IRwJhVDl/7qa
g/bGm0meTD91PEXbSnOgLaIIVEqHvTCzSJzP9qAeXts1Fw5E4Z7j0IGKEBuFAz9v
x4X7+KX6HT5xkb1aVifHQtTWA4tgiT/sngxGqDkXCCBcxc2+ruQqwLT5AAKYBMPS
Ren1ley8BhQUPE+DZmNukTBjqeF/UIEnHSOw4z/aFmuyTYtruzBiiYt98sgXqhky
AZZkMc/w0lD/kZOI14zD7PtLK7yirqycRBGGFgo7Np4bkFdlQahiuZwJ8o76PZ21
7fj9R0GYhPvibKIpYWjb5doapN7z/ueKuPzk0HELame4hPnQCjXfo05wW8jecEqa
hzgGGSSk17Kk+xsqC8F0S4HYzXpefq2mN0f/2BDs7akVsx3LB8UHziVABfJnEgTX
aEZGaPnxMPOFWsByoMz7OVbaSssrcSoDHtt1OqTjpzNBaOLYWMB2ylbB8PXqVjJZ
07lzlYBZV3ZR16Ff4bPvuQcTqVnPZqGUW8Kwcc0eZVrV1VgC79CNsKeUCcrr5uMd
kuujYpuDOLRvfuRoJBoHx8tAdAJvN5QYCjXbwRu/PXK4lqN7v1GMU3yRdzkCk+Af
NvIMwIl/fDZa4JQhuJldR0EVzZO18h+TGRo7oU7Rubl2opmIA6s6PVM37wFuKYLh
wX5zkSrK0cfeDmqWIruY5G24XeCFxRJOv5GhMxucrDSzxl160qgoFBSTIBKIYDTD
BrJ+uZKLgLRi+HRB2E/Hgbqh7vSUfh9H6NUtyrDaQtWFED0qWrw/gGd+XrLCa0Yt
08Df5X5mageTHDc6l6eTkHoRbGamOqdsaRZeNP59xhfLwf2KFy26rELslHUccAGo
jv6wn/y2c9EK7e+ZdKBQxTUXYSaleFVa0QCuLsDkdYWDO9VxrVb39W+bATjliCKJ
HUgp2oW3JYy6bFFS2Vqh2ISkq56WnZ5BaDLiio9hlKpLoMt43OZCi6ltIpFOegcn
e1Yg118Ie8cpHn2f/XAZAuEAZa2zwBKuusWJoVLdyHGeNV24ApEuWPNNKsd7NtM0
uD2IFkSkkAcvL1P9oaoa5aeYd6Jw4krHFpLH9xq5bjjzs+ikHRcHI7+lqfhbXYQm
E7jW+ozG8xgXHcvo6vQjR6yXM/PeFH4TEP1ja4EC58+6sKxTQZ4ssYfMPUEFRF2A
a+1I5svub0n4hVOg7IihdhxPmoH5kJE4308BXo1T/YJ1Ri3KdIzCqvgRJ3BRTq32
mExAXC+OBJIeSFG3WYMgQVUgEqVr3jVs4YaQ1A9Bv80bhqDcuGDBdhU5LbblgyNK
Mx2oP8NEoCOJyw2/gjF1VFeSO/iQHayz4KctBQ+KHibHhxGI/NnfKdL5Lvwq8G1P
Zw1FGX57KkpVgFYkaSGV9ht6EDBfHJUdGKu0oaHNXl9NT+rNe5YPD1x5A7i/bhcb
Ijp/dMbbhM3XTtkE9gt6qpfXHyCozy3z0W7nPGx00MaV4yXrZDUaEGr4GDYdSvk5
NZuMFVKX0iWZ1dncPWTkWezwovV3gF8tklC9Du3wJg6LG54JmHdc8JU1spZmjamk
mJdH/LTBikWidtznyu15Rt6fW7h/AutfRZOhgitccoK63LxRn14ihXWs7KcH78DF
c5j9Uea1YW/LAI7gXVjhDiVD7ZSik4AUz4bMYwA9Ynw4u2mYwUNjJfnBsLhZb3w/
nV6RMmcRSosud41oHD3014zRi3sNgExTpj2JW31WToa0YOE6NGnngkpoRhK+3uOb
qvpF4UPtoMUx7TlxmvVkLFivsBHooRFo8ThbK5c2sgketxtphGTpRS2ZtfP+72gX
+g18bJ/xzyCB0MMZJEz+Q7bM/IC80M60+Slua1X2BbowP1ZqrwTwdgsDRN0IF1DD
44LKVpTYWXXF0fLobx57GcNpxrrZzC5WHppbU0df54NPATjJazs4GwUFh+fadQHI
B7qQafmg3MSyji+191eo7ivWx6jqaHjEBw6LqBTLU9SwhP5mveIG/WWu1D0vMAqv
rW+qzUc7QNUoTrckPWuIcMMKDir0iUT80hTPJ1gtQ5q7/oQXF9t9/dgeyLRNbsH/
bOoBq+UYf+DYkzmvD39qH3QZozvZO19HcKMCihPJTiLeiaqqp0l9Iq+zuii0h60k
VpOLwFUU0Dbo8KAQoByzdkcNbE6gxJJUn3L1GbK7bcjyLWnV6JuOB930P/yDKADs
Z/1mgQWxWmtCSwW9pmI3rmsBVleiJQxvuLxZXQJbHBmpfQeQfZ4uwWAMWZ9GA9mn
eRLEpH7+Iz5+GpaNRIycCShm2/8PnVaKgv0fc1Ar6HhrSRGRQUUn6DS8HdEwKyTB
4mnDb8Cfb6Z68IfuH4w0pkvg8sqfmc6SDq/AcWeKArFSOP25pzCWa+91eo8BUROA
pDNrLEkEI66X/Iqwr5klo2b405JTi7wO0vWbArMmn3ReNSeVf4sMLvgm1E6+dlEz
9/yNoxbjWYXEux1lt/00JA7lsfQA/Kqw25g9KKBt7BZ6tE7grlSnhd2Dx7DM1RDb
NV1dqfhNbZKB8O9RHr7T/GDAjAhaIeUuKKzoGqzgTsKyy7qULGmUJ0SfEYKQprke
pEHjvjSV5Tp6lLOTqygfrO+n8uKBfaRTjhPEtp7xkcCFeZmrAouz5C6Xzez6qZjS
Vi4+maSg+0jG3AN+DaSru2JvNqKGf1sauNo6mPTdB9Ix1zRNj5pImNlBhq1LoHNR
28dmsl4S1YfaB9CFHP96CHPSuri+9rWOWeBC0Odl7e1dizkPYg/1Y1eHWjIcdaII
pgSz5mfeP1BRwtcsOtJK6gGi08vClTxGgD0sUIhq91nFTq656yBMbNkZQEcIiIXF
6ajvVZoT1BuSNN5bMGLOIW/uKjQQdq3YQxUgdu1V9dZ0004YouLrsREPV6dteQ7u
p/Ts+wz8LM+QgtvjJ5j8/H2HlTLDL8ewcVOtnkXja+oU8DOJwNmtQbH7JnoRl6h8
MvPFzjt0xGnD0BQ+CTYHgg3BceO8ry2h/D7+yMEYTv0Jm9O9e820yk1IQvCHHyr7
ILl6hzz1PINR+wtdQdel2kUYWGTmKyiT7RW1clEKErSRTt+8wY5d56EypQ6MnehS
Yy/vzfZKTYBIUfcD5u3KLlNvxzW9sviWeY2b58q6dlSJSehlyHrKSdS9zotrQcN1
cJUjoK4cpqo7FcizMsmmPBVrcF7x1Oh+bHF0vurArh7sV9wJUlez5tFS5YKivEAE
ToWnLmO3pZvedYzEudsXhw5AEQgLld4mk0pYzQ+aFMJ4rAnIf9in5igsPm46Lr7t
Q6MHHCFPXNSbRdUuIFrBNmOlm2Lu7RH9tKUPM/OMFTrFGJuzP4r5XMR8YuV71M3p
r5aVGWBxiE4I+AtGsmQ2ZM2viqweA0pzxj8wivDWLn2TbOXqvYpDGlKTEr0tzPez
4wTNP0QY4N2/1/szvGxzWPkCLGkzo0WhP8Ddime7rrR/TwTMQG0FhoPC59uuGEDD
p8/N39zh/1AycSDKEl1ziKNUh4E/pRzZ8dyEr3Sqj15AB+kqOqwr6w3duE4dlg7v
fG4BCCCmtTtAxkp7NYD8OCRIrvTTFhvgPW/o6JEQXWrluPHVZpip5BNQ4WtrtMWF
cUaWFT76y1OCQXnPDBO/IFOdVVqkpc9W1u2OmOo8VMD7ixM8hqDGeC20raH31r34
XXKNnTQyAQRiw1QOQYzb+9PvfHIBetYuTJ1Q+i7Mmyzs5J+WS+ntQdoyF3KI59yM
1NQg+HiG7YkMNlkXs5S2OHk4neRwMcHNQImcur57phjgMIZsHzuncecWMjJKy9Cc
ryHvdtUU1eh/+zHrt/Ne4paUzEj1cMYGLB6ZGR7VaTgmp04jHX3du7yKgaa+r4xD
ydsKk8a/VJahe9OB+f+vNc37biieBLDXvftBjkRyGZ0w2/Stnf9sveZEhC/mCaSP
BYrNRKnmEK/F2j7VytookFC92lImizTpjoLASd4H4l4qSUDxptihCCgSdxzLDTBB
aaXn6Lwte5YYi+WslgPOtEAf9Ag0eZC1+jEznwxwZp0z1iEqpmKfMhSMCfcL6rJD
LDgkxiGJKj0suaccTgeYQFnEVM50o3olV70SboSdOQLg6NScBh6WZG5FpSOYeTJy
wrBRf+sKIVNTyaDAS0c4qiv/pSv6fgZ9IzSfQ7q4m7Nwfwvr+9Y+oAdCz00/zgNd
Hw1qnWAT6iggxSfEp0+pUQP7olGa8z5OA1CQEn/AKgUhHq5jI0cFvj+HBwQC0RCj
S9BiSc00ZHXUYTTbU3kdU9JwJyOJ57GLPvysLuNd2UhXhE/Ovq+d3fRVC0asuIYV
gcLbZyFhxYMHHrhxGB4mmQoNvkViqFlLWX5vHk37TAzBwuC5H4ZWCVmtb8pTu/nQ
KkR4/v6AMj+OiWnxveQN24V8QhM1ciAQiyFWeRiWhiWX52sdDxgG1CS3soeJmtT/
N8zNTaSdpU9u9qq5+WaNw2MuVoWQJHnZ1MNBvNeNskkCtRzjs9uJ+9VePU04gus0
U8OIvLQ4BEElEdTfuMBYSSrzwHhRken8OAD4WmulNQvGx0cuBQAFqvB+sLga6zzI
zHeEFhcdDhaDu0Yw2O+r8rMzOOVtfh70AFmyNRdWJGiBzshTiB1JHJUz4p/LtFMk
mJos1P5mPF11BR85AK+KsBwU4Wcx79irdnlnTbPKqVPGJfhiyDiX4Bal1t+dDDnr
lF0u4pKcMLMdjBQBT0tF6nbMlqUdMLOyCAD19zgowwbK9POlNEDVvAhpWUKZR/bs
OJDR4zSXt+W3XA1HEkOx6JEzrgfBGfB/HcqfjA+WqJYkrYeqtjg2WpEukEPg/KtW
TDUJrRfLTqw0VWqkso28xQ8RFEUUrQ71GXqv7bWP0UH11smWRpBh77khouRzFP91
p+uMqMw62LNTpopt82TFug3gD7pksR4j5yWs3KY3Uc+PGvaXRjDSBmfxWj9jgsr/
dxDkLDpRsqgUrsbOiML8QCQELRh/u3WTqm2fLBx6hFAnd7Ca9yjDGj3MOr4l3hrw
pz09QfBCMZFjgtnBoaezQUD2nse/hMKD1bhb1BkK9YuUMxx0U8CXM8Pl2Uq/DD+n
Tlx+lYhlPLE4FNRRg51yWtexzDdRxy2Oa+o4Y8vCuWsR+8Q3LZBPyvjcLWtIWzzI
DF929Y17eboV4Fnqr9UQnWtfthgYNFVlaQamtgkr3oIhU86gBWfBNPxRs5ZeGhRz
HjaRK9ct4WlzkBRkAOTVVXRPxLYN0cUnV4clZaXBwgOLXVr+VTKRE7Pfq9rgKJWJ
na27seXcXe+JUztPP5z0XwCh+hx/ocM5vhJ0QTvYfqWDOIyw+TnynVgEfaE2nm9n
HKuvb93qnelwLCKlLBo3a8yfQmDawXIcbxPtqaSPScRn6HOUYUw+HSJm/SCwM/Jj
bNvakEDtZmdhl44Wh8oZwtKrpr5F75FRjjrobrEsJsnz5Ce3/LiydxgCjWIX1E71
r65y+TCUI1qT4fGf06a/EDbneJYqccfoxCmSANoqspbInycIZ1sYvE6khkC269H/
KlF1kLW0oA80i0IwvmLVccz+p87VYcHkXXtoBOFu7gXM/7ngLp95FhusCby0zCDe
8Zryb6LLzn8jMtRHsQNoJ7lRbIgSZDicG13Oucp4S9rHHnwSwAhAqYuxtUW+Hqa/
Bri5ENf6qzOaFNpgieoN4/cd4CAnpApdVqkIJDMFFteDlkKebxCDkLfVUQ9DaKOi
BnUhFeGsqcOqf94qM45legyZIubeNUP9WU7BpUgmSqgPSYgx+HmHzvGcrM886Rw1
gyC2Z4rMfyIizMg2OIb+tAFpIFJQikz2mg7h5O2Y/e3jXYnEVPX/yq6Gs/Q6Tj5D
L5OvQGtT2QDe1JB5EBM+MskfAcB0hDqlgKy3LXCy7uesboCjHlJL/C0m2SlOh850
05gTZ6qDh7xoE0/4zvnjjEvJYb4LuVsD23XKTmh/Jv7RB6Rr/cy3XxJE+hxlpQWJ
yepfBjopY0wbMolVw6+Io4qzRsk0PyqzBz9uD68GTjC7xnOZhEq7d6AFsyVOn0Oo
V96897w+5ZKip40k6vy+mPafrujmw/moXp+gE78Zz3+D7nVWZBegCnd6S5g1KQou
cdxHudgbszNaXqigH1eduj993CWS/hTUv6lWnbPKqoBuPGIHYptHUGo2KZLkqEJK
FUb02e9x+PkEnP7YV0dOxqLnvU4PZRSy5aVaCdGmahqLyluOGZ7y2M23u00MWvJw
bkfghhc+wNJYA+kR1qOl2K3skwsiEvS/msIZuHH9FOS/7ykR9/X4TNJrvYqLLw8F
BteEYSAQfKR1yuRzNCj9sPYbx1b2QG5ucOpzqsV/xXvg1G0o1GudMfjh4o4S7QMK
8x3Z5OmiLzUVRYFAmSfNvbSmqJkuYX20fGRMknPi8BJNU0z+a88UACrZbt5fLHKN
4BndZse3dJ09GHPxcS2LtuUIGwPy8KtjH1o13MhTO/6A3rO6u1+DQ5Jtz9Tw5s6u
E6tic8gKIt2HoaZobxa5OA0Jb7nl9qikgym1IkObjw1UOJ8P5IFEsaLoUOxeAxcX
GnnqJr20jihQF4mKdIDtz5Cc8p1W7oSGVOYTnnG7rvJiKnxefBbugDfjp/fuMkEt
VoGeS43mNwF/WG7LHwtMmUXm6fcRhPyEIeQWgKRbGieuoxmK+82x3DoSnXadwOtA
6nDrsTobgJV6P81+BOmZwEWhm9J7Tlc6DcFx1qE3E68fWDzhIwGv/yOKs7dmCAjC
HDhryZqAZKCQp4+Lms6z5KxG3q1c4EhZsEaIMtv8njozv7p3+fGqHBgmTT2qltpe
wgw5xjyl/bn0r56RXwQ9Lv1fq0BNlqpTojf6waSbEm63DJaSkqxFQjIuqyPyVrgn
VSCIc3ZVoaHgkHtq9n2dn0/1EA/P+odE8ke+SpEGoIbyynHI0oD0g3OW8irs+dy9
Nv11RMGdgHN5oEyGjYiBOLrxAI3PVN7P3AJ3kJJrvMO8XYupC9ODaeisunlgS3yU
3KHEerm+GZO7HC3Nb5kwo/eW+Njdg8eMBQLWgE/IDbwkE5x8HQltTLfIb9QENOlp
xlRV0laUZG98dByzxzAayBskr6xn3RkzPczijT+juS6QI9lC8juZFgGuHwwGu66Z
hLFkWFwAtb1hGC0PphBwOwnAFu8iRG7jiAkpqi8K4H02CgpQd/MVMqda+uwODnHI
XIBf1Xy8d/PQocAz4uYW+yOCv37xQ3X6IZFO5auWxWW9R4tvRomOleQCh4EvZz7U
WjNjrmqPMs5vuhJRl8M4ed2Kcug90I4tZd84+NSzDtBhZDTwj725f2DL5BGmbs7M
/Wnr9OWNp3vYlsimPi70a04/p0fzziEPcyHDMDn04iER1qUm2hiJj2uD5Y9+NE69
QRTGOOLKF40/PbYrDTrUklKkK2jb2Qjm136JomaX0Xg9rTSVIQfJuQdcwZyOT/Bi
IH9EjFr4MxumSP9Nsq5TUHDEGetf1VqxUkK1L3iY/rFAwH9jkrgdFJwJFbFnclDA
wwmXTM+gH+k7FWCYChYoUubOSOA5Zc3G8Diz0ow763yh1/RvToZnwWJXn9OtPzOU
47v0WqYkUR5YGtFWetAOgQL3lbgqhZLOLUJKG/jevfzQKQCKrA038Cj/HbjweRNc
8ifmOR7+HYBPcJclsHH7k4BVbEmrruBQJaNoBvqyLUkDa0VRRPUeyOtbPtjjB+Ac
QALau8QjF/KfRVT1y2u033cFV/qB1OCcDoTqNOpzSTrcc9XZU3P8jjVhDM+QGBnj
PJnSInwYIRQbqjoMD47+wvLvioWLhr72hFOcVvejtc0SShwDAxLCPG6Ix/Y8MxJM
pp6RSvKWqdIIYHDzdaASF2OWJTHzCMsbT6EXI6bPT8R+et2EsJ00p6bztXNU7/BW
kauD6cRAZjYSBo+LtybNzMd6SISUrbanYl8UT/octyIP9hBW1XM6lIS0q3Y9ccBV
5+FhpFzByyeYXEqjHvabo1aAghLtzlxS6wwFN8uJBh825iTd22aRdho8YkNYReKH
1t+zov+PK1fHWmNZHVJi+e3TrFzvDGN5UemQD8VTA4NGwCIp9AFtjTavU/eXVFiX
Tc3oxb4TLl/Egcp/Yk2YvK4zUBCdDsqvEmtsZ9cx6MY2+kav5rngYaF1VINCRXHo
3g9F95/xOT4JIIsZOKklB7pfZkOGw9pF5KIDKVvdOlloJyNxD7wLND7Yl9IkET8s
6lHvVXxlnoVtaliIelKxy4hwy5ykKOboMlHjULsFKxNu0uNBfCOeFOHy4SIjjXNJ
CanI/BRV40UF5+KbCfQNtoaKko7ZpvuSc+bT+93MFUGYZbSxpSfXWl2k8nx5a9JC
OKXgPzOwM+YnLdanDDRzgEs0Zsl1ULVIPIaMN2E69Z0jv2YMxJ3czqaYt8LZDpuC
OLptnCD1/yJ6d/DEJwstIBa7YMOJdkrQrMIh1Ie34dQnPWdWIy5yuSm5CDyK7lNz
Pe+OvEZVxCmnIpjHNQDaOWr11WEr4Xl5QLkW5ImYODiS+PofcIuy1DoVOKTlhAsy
JEfMEqlvGif6hjPvqA4w0Qg3D7kZWqGD+CRMCMHFMzOjPWfJOnodC/YYpyhQdXLi
lCaPj/zHsb6gaWlWJdtRNIDHasEJ+36arZRsgkmrj3arqpEb2JCSd4pVNiSQ825D
PF+3hET6GYP0KNtV3kurx+ml4aEPA++pF3eojMW1grd9UNKfszEdGIwcyNPCeFV6
f1AKLrcBGCa5XQs7TKcZv+pyPD2aPkgpLp9q9dBFvOXX3TwXstIRUZ1q/tI+vTbs
lLr9dkyHlGU8hCHSqq/3uOO0x1agGYSSNqtkA9duT+h1QRy4G0t4XLlMHw5cmMQZ
K4jrrgleF95LJ/qdKi7b4ol/c231VpplRFLmZqpCbqBOy2Q/T3ohsfafLQ7u++uj
SpCqb9wRYt5Hi43R+Erbh8ltW0itduc+RiBkTBmLX19wyXDF+CZj0W/mPC6ziT+F
6gFtsluWhYvydFtz7WT0T6OOwV2x6J/o0fZ9N/44hOt5mhpQq9T5Nt+O97dyB6it
LuYv7yZkrxDb5vQGgO0+7k9H06+IoxuI6q7RLbOu1PfpJrmRyYKrh7UFB5BGHh1h
0jTI358PrTvhg12OlWOGmPtMUQJVuLwD7ObOrb7eQw8v+HIhexvISMoZ50opNhuc
PCzCnX5KM/9p+5PaRTdg5W4csokEpfSWwGas7Gh4XGkXHD6DkgQwjge1s4SNFZkk
llcFYTdOZMa27hm4sQueqQQBwRWdGspF58fQ7sMwKigO6dNtnQE+PcWLenvFHsic
jWNBDx8bJvTaNlLjDWcKHtgSGcatkAAE9ajqtFkv5Ra6oZEtXYnGGvxLu1QulyzM
RDA/owBbYuLuL1qYN7/yrPNG/RNtrNb9s9KEVHrbTgXP8zoEYtaU1pAzfkxdBLyz
zpANUD2cdw5Ny5W1k+bHN/J9Emi4ug+p1n9Mw4Zl+Ibrw9AXqNQ9InKRqXX8nRQc
YMoJllMq6LaCSTuXeKiuHGjazi5fBY4eD54CNEY2Vdic66u8iRKOD4Kj8IndJ4us
5mkoAI2CqjiUp+/r4lww5iWhjhaoOUgplGnugbY5lNSIZ/3ukLt1QZ2B8hMPX52j
+0V49tyAK16X7s5bw9visY+ZHvs7H6RVI4DhbrV4AkSj2lDTMTlgYlbBQT1jgU+T
rpl/VN21Z76CAEt8+byZ0GwL8vpYLqMyDGcBVe7bY6gihc1LKFyjqI0yyFwVLCBW
HUWa7xFgYR5T4sDLDDMZNNVyuYhylTh5zWrwzkdeVUnEgZ/axQQzk1fkvkwohley
pu0znnU4p9fmNyjlcRGP+kVv8B6Bv8+KJFM00dbOX8ABM+38UXKEN/PDDZRxoGJX
TquPRFrrDcLHtBwOUxvx65i04vrpTNr0vj8V2Zd2M1wo+xWXGpEwgXUoRaORLD6g
oTGay3FfHX+s2KAbk2TfyMvQV09Oej4bDoATW6wZoN1QJSC957e8AGY7eHz1WMcv
mZqYIxfLNTcJji5yY74kFrEuIi28u3gk0RaoDf91LJAh10J80uK5RSUf7U4uNQpj
KzsnGV8MdiUrKU1+3lyYHvSba1XgXvRN0K/ir27Qysjtvqk3INnSZW+eU+oWZ9pP
y0ObnpiJACYFNAFvptONNyb51dVsx6jhhu6HEsXqy3D5VNyloC1CKmbz0c5psq04
+u/7j5YnhGHlWB7q56aIXK2MS4TGU6NHaDsllDhflI9vs6ezAWkWISKBclxNfxCZ
0igo2HG4hWr60tsb4NHk1WlVYlqrUgiMDZxBybnJVaUMgpwARI9hHMeZvxH9k86Y
IDs9sJoWhFwbVc3MVWBZ73+M4LXvAntbWCuNEEGWQ8g/MaBp/txEQY75VA1BeUbZ
KabJ+bLrDk3uZ0F33ZwvhL1fpo0JxQP4z7i94H0hQNccl+pql2+HDepCt9lLEhd+
IMZWMXi1bpJQh7E1E6SJQ0m1Dmzj/59ekn8waIeh4to5UVeZ7Kfvvid/1c5IaZq7
bQM586DkbiyIj6qvRjCsQwO9ZXl61iSiP6AXMlEazyai3XJlR7H+fseyBbXlHfC6
zkNdD25utomkbrDp67JFfTliPAX9Bc/5qZ/J02fUqV/j+VRPGdGyGIBUjkNg3XI+
HHs6tKCkxbeRcpNQUt7BVraPnZ2k6eUPtZ2kmweAogSht49hJey3jgrMvJUbdfxu
qqq6gcmny5aqgn/SQNI/VSXUhaT2FcVTJOO9moqTnF45OqgHRKjCQwTLySosdgBe
1NHo5GtcBmErHKzcAlagjEboZoTOyewG9mRx3yjKFqywLkrMGdxX1HaGRqjZbKQD
l2T19Tnaa5NviKwIWlxs3l4Bo6Moqw2ljiqeXF0+xmLxrwUiPv1QSPpAWYgUqiEv
/QtPq0j/+QgJF/Rb9qvDCHUE+H+709zYzM4vB1ddZPUl/A52p+RdVl37UmBMOcr+
Xo3Z3mK6fRBWeSK6m/CcF67zAvogZz8mICbRGNTNiZSvJtfvJwZlqeKwpn5TC4Zi
H44vLe3dd9lUS/+3tffdEI5GxiRM7zOiU/0afxyLarj6esH61NYNQA/MgMfHDpnL
TNmOfPtE4APNRkkb4HNqhkLKunpmbUuWtUuWxATdcuff2IHFSVVNB8+3cDQ0nhzg
j5D04oWNaa2tfOMg+v7544Y8KipU2d6LQ5sMNGl6I1c86R53Ah5S8FVUjUQtty2s
89rYByqATBY1nZm6hHskKtO5rSwjFQCb0r6r+TUYtVbY26+vslk0yMd1SsHq3I6t
iBnbu6drrcHB+ZncTRzpJrJ/EXCce7wKwgJZfsfOc2HJbHVkoPjuLMx/b47oGwEa
g2GFocP+Dt1KfVMH1nryWwlaiBZyJAUcagT1SW+aYsEJPHXhO3MFKuNZuzPsKn2e
tv8ResPOSlzSBwk2Yfyw1thLpCAJqGm8cfMX8Ic6x8Ig2diMSELfYpI09j9GBxAd
VomH35ueheN3pk5to0O/0/Y/mMV3U8pRapTBySQjUy/AWfMkMFAeKDk+VoViiRLr
WFEOAF/ih1xLQ0lcu5o8SL1eSU7PagvRh/f6Eo1olhBwNi/uguAh4DlY8mPHpr0P
ak1nO60EN8Cn5j8YGgafrEiYjeTHLGCD+ZnPPXmTPsCLKrq0scb3Ywf1WTa9m/Wk
Sjj4uTbTMkBhdtJpAfNt4NZBrhMllLi5oUeGDEIikOChj2JayfXH/Sf+XyArsLBI
DtY6PdWLnU9pRA9dKIMJOvWoB8NXN/KZDFclwxQ0p3Z4YbgmzGDPxKg5Thvxina+
ljr/xZ1+FWqcGqw/TkZCSmnF3Q3dSh2BEmIfs6YKEu6D0UpGqlrwMBf6G8a7yIbi
Xz80+RlTWJ07r0z5bOVH8KbtCVZ06BmJY24ITmz2qwGdE0JDq2aqONqzaprE/17I
Jzwf2ahYTaHqOExYnPeDVDBiXhR9lbFCRTsZVXoXivXeaJrDk9k1eL9MNgJCnJo+
IHwvDrOCx+n6inEWVQXYmNGKqm0w1q8KOCqBFNDISUIjVdh6n+oyBQ9EjAwO6zPh
Lu+eVpALwB2nyP5vdYefkKXtdN39KqxjHWxztihuVuDKorSvlLpN3nuUd/gNLPdj
5nTQaHruJlGxlJ0fLeA/8c31xk0++5scHpo6GseYwd5hDqd2DInTnPdrxBy2QgR7
JbOEkQw68HaiiekYf2g2aTQliF5SnfURSld2coo75qYu3psMtsbvX6/OPmtNwJVj
uN7G/nu5f4Yi4xDWTfUPWAKFNPcznLECHO575lpvixUmYBy6NUuaThrdM5ZV9Wke
E39CuklEBxV+pVMKwAkAQyyO6eE8c4s5Sr1LLmQXIp9FGSZT7DzymXTeMPh2FcXt
227MB6Owp977QKVQNy+FsUyMF6TEmif6xRYA1LuU+0LWQ7+MP4wwJq1zabat8u6U
s00aFpGCK8/V6Iz1I1sNjqjS01mFc4XngT9QnewCzIcs1V1J1zRUJXRomDxwmz8g
vrMLqVZds/Ee6btFQ6z/bGSYZ0veyox+3/1d1eFNW3dvodKpsHWfKDxaloDGk0mc
EeYORcyWdifSgBXrtMA5x/vy1lNPRfy/8P0kapodihRndjrxumR17v7TyDWBqTSS
iXh1iqHQlW/4QuYwO7kQ/7VkNfLLcfdXubDlA/lh0VrL5zcjvD8h8Mx0vsmX4i/e
zsw35y3baVkxg54F22G91N/DlwHbbSkJq2PaeWa7UrpDof8M0CTpSwzlOPunAeLu
QF0oaRlMRLjr+xJ52gQmH8javWlpBxc93wEayJB7MXvL7YiAdI+1GLzQFPAjcPBe
hHBu1yap6g7wUs8W8/v7YlPG0wakf28uvBX9yfDeRccd7mt8tDZVe8W+PF9z7bWS
dSF9AKKzHItsFjp0MquAcTLJSz3gggTWo4FBT8RHeMrG2NHup2+Z6xy8kWdIkv7o
b9zLsp+3exYG66gw/W+2Lvt9o8tfAeVJujBdKS2MqfiEiGwHRpaX2RyzwRkN/2u5
KE+DjSZaQpMjQiJDpHdPIDkzQFdLaQ0zxuW5xpN37lafgBcy9S1ys7zlpN4L8/2l
r5j8SiCZiahroMURifi053Xb6QNcDQaED2AsAXIEH17EUdWRS+AQE+42chNS6PE7
quh4HB1nrjPYLHPm/lr85os7+qLkU6F6L6bls8prB5wJk7cj57tuBrW/MDCJ0Pv+
n5m1r1C6N7G3QxPqcDzX6R74xV2ij2xOeNZcheyLvLBjQhnGSUeoX/kF+DKA9Nal
kCHqAEDrfu2IbECJ/2juDKW9Q1/vv8X8pUXjfJqJeIWIp0Dy0vz3dtuSHC04k8RP
f8tcUF28l2/WQ9EwksPKLeM4D0ymL59Neel9HdVRTCG4feYctSWVn9guOsbs0SD7
fg2VB3N8BIqr1otAxqoFGfoAVLtG4zAR/vLJtDMPgmo8xcLnZrrblQnHpvEy7uVx
tVVsMkzg5hl/cvv215LpXS7habzSOqF4hdr5qHj+mS4M1UvsNicqAvre4BQLx8ku
0r/8gR/64mAOvXLk+4xpxJtdGk1/zUk0CjclSvieArMnk2C2DKFmQadnm963h1DR
2DfMosHc7A4Iig+flewhMV/RccKZdnvQu3oyyZE7uQyk4IEOiboxs92e0Es5UXOt
DosfH67TxxQqvjw5TFrvK652lo6Ija+9kAGfn8qd+jHkYB0BD3vKIHMvWgaZNCvP
W43ACQguj/rDyX0SGoUNyTgiUtMqQKR12PQH4j7QrkMosmW6/aDU2cc4tumYUhC8
XKKePRt9k+JKx8F/laaqusIMnk/bG/1tk86EbJB+k/Z2YS/e0wSoScSRItfxBEUf
g4KdfQrt+h7B351Z0ZfjGDKkQdjjuNwYKz8zDY2E8aPV9FbuAawP+NbJzWEQxU6u
dtLIsJp866GfpNSxOYhmJ8tU3ePb6VG0YiSJbMB0oeZDm7CBFwIBaq2C/NNrqbkj
Zy+t6sS4IF7zrFWHOqYqdopEOXC+91jo4j4kNG4V+iLznLrS6ddTe+/6JZalvVds
KPo0vEAbp2pUgmIgWlbOxFtVcMvRomF6/qPJd9w58WgCD0hZwEvWKuuB95rG1u3t
MggAHF4lHmSawSukgHRblKUe4S5u1E62gMfyE07XDdSXdnKiLwT/R7GD4AnOgV4x
pI62p7AlluHXRY/igFTYlSjM22f1FBArjzARdgPZB4h9GwTVWHBpkWLDrwQxf98i
6Kjcb//ZZEoCz8WJNCS0vMztBw6OrGpWqQrff6xcGws3hlzOnQcr+XLYSPuuCuzJ
9kQaIuDXS/wqXjx8C6atqKVXZ6lZydJp0XBU9ZhXNuxGVBDSvAZ8gwrk7+knzNAo
Qzh0Akxq56+RpuKmayXaJWNud1uIEy/r83hkisI+whJ7LSwF9pXTMnS/MfpFyq+0
NibzjiDoQBfFTCvGqQXoNkeD6X3azshQPzjl7QMFr8nf7EsEa9tuQ8wJ/D6ZR43C
fguz9bSDjiIPb4NcrhPfzk6SUM31fSe4PqT9bCDbPIctAKi1kXG6GhwqZ9ICLpCR
RhU0fHT7Ql3x59MkgTjGx5X6d5W/CWjde56fAkQhOHT+Y0/HBuGheRW6Q7bJWLA1
eWjaKX5VCe7u7ZJdZ2oOLN57R5WEc7ZCs0//tVgNYX+W2f0Oi5JtrQ+hlu8XswX5
onsUWt+GyJMEA01xudRIaM0KUhqMxkfln93DvERzoPl2cPjNTxuTlyG2coE3mi0C
BAM/XbqEI7TzkjxMfQdSntHU0fwnXjQ6NhdpyfKfaneSx3IlJcwGOnyEV4UEoJZt
w5aiWYKDKOF4/400g5HPHaoRyudPsizYq0nWXHDQYnEO1drDOSdIIjFxLTQTCkyb
eQsLSwgEZ8Z7cnmey7ycFt6idZdOZ2HSlhML3VvHgW4K9jcOl9s2B59k2/mBwk8L
qitzZro8as5aWHkNYGpDv+FAedl2RdGZBE/Ps1FJ4JCAYL4BLm45VJFvq1wWdNh2
kagRgeFIm/MZW1Zurkjmsclg80jWN9IoBzDRqZvMx/pweo3FOXfzj3mgqHnwtq92
CgQTl1OH9qJ4wsLj7ORt2BpstEyjvJIyiPtswZ7b6sAgQ/OEWANktw7zRWiUwsIl
FLCoO2+u4FJn7Rp1UtgKfxn7Rzjib38kH5/VU0jzLU+eKculrEW2XybLrUiWvpWO
6NlMAZKKf1rsXHoNo1SflZ0D/COhrt4iOVCTAaznGxvg1Y4avp5uyg//fil9sMFz
2NTOLyXKHwd7liKl2Yk/22qTyJ03OoyHBm3N8NSiPS1o85lUlm6HUcr7DMqpBjaq
B3jgK9UcvdcTM/146EARVU00wRes0n6Lyd9kCBmkjL7vz9S2wNBuPSc7scTtfYsQ
AZNDiNw0ZQlXZnbHUSJ9+b5hzgl0Ja7JRt8rbTsBmBYBooQbIBBCdGMYi5OD2MP3
APFz9rf3LpndoFIiqkRGHuua+nubSRc/lKAh/NGNp1vBUMfnNGMuesm+pqFjhssh
hiUO4dBq0Akhyo58rfmmTNWCiAR8aCTLc0W7od5Gb6naEl4uJqQ+68V/dtl8tx3A
XPaQokXQOEd6VVTB/tMhFvt21CnfrKdRLs44QEkDaK2bIzOJjM/OyHBD+o1ZhaYs
qknQ5gnr5xarunP5bnTV468LWmVdG1FbMVSfaq2vweuVXWmza5vQIWh+DA4y06pl
WTpLOBiD2uufcHzelBCWhBHuEqXI9Hyy+Po9BhWX2a+BQ65lXp8w7q5VB7xcF4AC
m9MPVhoL36qK/QHhV/eMVnwuQS5OJch/uu7/YnBMEFuhNBlIv7M9+EdXqYvSFq2x
gw/XYqCwXBTXDk25kczN/QIwSFPh6JePgXkyoDBvSH35Ta3RfrZsYW48oOLlnPzx
4xNOIiTNPW9DC/p2sBUNlyupU5xqDj0vCFuGnDlscX3OwthpzxhH9vayQxbD60wQ
+rl4KzuV6joFSRPhYe9Sme9hWI3HhD2j3l3lQcREZYTMTTEzd6w/0F/GzpX7v2MR
JWP+pfDCRfI5Fk+35J0lVCEwpP+dLTok/aUKiNuouj+vjxi+R0PTyuRRw0zLZTU0
Z3jtLSFJlSeW9SsVp+YYIFcFd8hbcn3WDZkWJobek5j6vOIoo5jgGWNj22kMpCfM
sZnLwYR8iizBJUaSzYdVRP/pCul9UmXrbAX+CYnpLsXE6WZK2OC5mQLKqn8eNFEe
jjirkTbskMSj0ZwTbn+YI//DUPz+EYOWwcmntwKshgg3g8dZhx8f76aDa9m9bZjJ
OnqfFscUv3zed1AsKOH6Sk5wMDW2QOCxGMgZRTLygMNo+RjuGDmxw8R+heVqiUuM
QkynIr4F82en+ndteI8DK9O7CHjvW0mNZ0qZwddK5MpYn58bIHpTKNe6CKp0CWpP
mh+SzNtNkazrSqBuiJAPJbnrLgcN9mId8yMnL/hi0SnaEvWA5uFCkf2AHdt3WGU3
nRZISxvvKuv2CHtMfLroUtd6sw6QAwun/t6I0cBzJk67Jnz+l3WpsgAuzxAIJ9pi
UD5mQg/yoYt0LrMdySKHpfoDMUoIQdOmv2WKtaFK3iDPOrfc3Aevf+qWXxABWAWx
89xY0f0PflHjmJOrn2AqzLDnb5zdg+xQSpztUL67djisdcGUw9OlaR3vv6QvnyX3
Omg4K4EYcOKIspyOJSq0Aa1CDuw5H55WFD9ByN6j/BBNp8bY2/H7MydyNnq+7g4H
Af6RXynYM806B1jFchgti2ROfXoU33Hb8aXFAkce9ZtNXVvZv6fU2+VebMzmGVE4
JPYYMWq3WmIM1BjWdKriF4u2z1qJs9igdHXpn2IwTB+TaIhLNRiKQxemQ/rDLQAm
QznMpyQDBRMz8uPVR9GsJtLSgi7FzCRgtI8dYh0g7rV2NaskO0EPtOkgvYtf1ecz
7umWpsdMT52begorh++x/1xzUmEJfusnExvg+WN4RLKKfxwWw5slnNUKBtZ5lZ4W
sWjrnuizeJ79cyEnYpcEaRekhHnYNjd5jxOkosVlA3blHttk+UslS/voV5vGWCiW
HLcU6FCXXs2KjgaqQhknlquJnoQ6XYnutxF/+hBJS7iHLwbNHYae2sCZD1V9lJ+U
dpqi/cFKofdza1kgcrmX0XW7suARpdrjk5FwUJ8vHM73vVcJDX1CVXgcNlwKig20
SwIkJRnleXX2jvCzV8eoA4jfadeV69K1M3uABHZWw8ju83Jz5Ee1EQ8kUIAassAZ
ZOmpCyu2ogRaoh4+PsQkt1p3vG1dCPwSarNHHXOtHYF44U/7wYhJQmyKtTGTBQmF
3sTxXCh2JrkrkAEaMxWaTg6+6I4A63aGOfSK5YFvEPu4d5W0wm9sHwVCtAf8L6Kg
ujAqdHuK0pAcX5i1geBWrxjMQ2uGlVTsUeSykLn5vSh4gmkR+cynYUjgDWRej5VU
MoL/D6+iWJv+2nIGXNwM+YG/SjClVKf1rt+RpFU1ocmBLv6HxBETZNR3xPopq5Sn
HHQW7OjLByo+gMrU5+IWtDpMUHpfQd+/5l552eFfRAYUDv6IYZIeEURcI9VPPDLJ
5wAN2r/23qVHX7UKxrIr+uDxjBA/WBo6sba73xWGrPczxKaRfCbk/y0ORG0a7Ab3
O0xH8tzga3I1k5VTGNyXP+/TP+zq0bBsHDSj4k7NDUmCtSRD6UzEAt05cE8cYp8e
pQ5kz7fxVjk3s97WBzMEDHhtGz2D7NGJNC8Bu8V9xkzaOQOEgRCT6WIrazchaMXq
xhBJlXdBYtdBwi4O1sq2E0bxlWzTfsNkv8YoxmEyFW2/TOMqBGET5rwA81PmI8My
g6vk2Z4Tq1pMKtnsd+LVicggTCnIWGbQqux//mb6JunL6a9xfKjMj4Uu8d4nZJxK
pEjUkDDqjCmaGWFbR0r/ftkqAF6mmsk+4xda2Md3aI/04GMRZcWuVm+m1bdavhuK
XP6bi1SBOq+UnHSp/LHfDLahQMaWsjyR5iD60QENh8jrYgDUQRzv8ZNP4KmTVpUS
PvFeJgSAR3mUgC/TALkLZBRToD7f8De6f7nX4YtUQB1B9l6vVjqx4y8trR3Q2QR9
52zpcyPEdD4m5mRvyymN0X0RZ+Uz9e1uskmOb+WtX4QHccnWCTL6x77G5PkQz+X1
aeZ/X6vEDstqAC78t7cIgL7EER2aQQf7pWJBVcry4iHn3UFadAzt1UdyfV7d2l1D
nXIKYQ2AxTw6K05AvT20bfqkTWzVD62hG4O8xQIqMFTV6wCUPDdygSNk9XqcUA2P
rii7/QPSLiZ3Q0UAkov9p3furo56EMzAjGpV7c9OGm56hU5Fgy+c1WZ5PmYsToaw
s/Q2OLem5Pp7ZvxueV1eZmmKApdOe51hFEklENU3yMSqFM/aOB8Rcyq4anNQR4Ln
0PWJWnbRCHB6SElaAAfeR4GD/xAr13QzVlGovuf2jECkeFkbwywNkmlvINDysTYZ
BvmLggdxwcIAum4LQetFBorHWYiacjxqt6vB3wh1T2dw/oLuwsRe+TLGIJjFYIcy
v1V8nEW1LfsZMdK5CFsW6Fb9QfMwVG98MpTldRvkkn8HKM87j0uYlgGPUeCTbQqX
ipAZCm41MypTIjGXGB4eOBKaN3Rj2RYFSFJ61+CivQhPEpgi61ce6K9T7Q/+8S6a
mmXKXGC8C+9vet9oaejECa+aIcP7IMWocXVVcMefPvVBS7rXTU8LPUaLyzf2A1xb
c+cZNlFwOQLZ3hdhYPnoNRoIQeZwk/dTzg9MVEwY3IJebrWvbWQUWbaii3gXW1A7
6YEECEZCizzj9OShfPoF7I5SXmhNnvnLeTU1nJ8RRHYfObUeANJTZJRcfyBFs5Nn
mQdgU3zhxA3LSK9M8VaWg8tj+gr8zVZHjSrRV3XI0eOilxjb/sYSihcgHkwkAnwE
0AX2DP4omXrIncz8hrp6+R8WNA5NQAsXvX6RzEoVWL+nVgt2BZp0SJkrXbbvVXnm
N/JLW91/eejQI03/ioSbiooXn6UDu1+yYgRaWi63UapvPiqwk03qPTDJYswSivAZ
AuoCkud3Dr5Iku/hcXVMfcKfNCyTaYTrkOY3B+jwJqyRXWU8+owzAE8CZzqUYfz8
lzXxyxII21V3Vsr0hyUVviK9jTSPHwfMys3Bab24M+d3Bzg789Svlg/jClqjYJeZ
2ms+tyqEP9cq7/7y+UnKdudWLJ7W07B71xuwby8MAzIm8KdUS1ANWXDepGm//hiA
cvQ11rN5EmsDG7/8w+PcHpkRdTruMC1R80rBHq8nTSsiDzNw84GACdBkuWKXE8rE
gVZbkYfNfuJaPiefjNqLr6sK/+StuLGhmffLVakyPfht0BlCP9JOgLr9CuZ06Wfk
0BTgV4dD7jmY/OvognjQ4eaDmOU1ECt3WRxDl39s9UtazWPr+ozlQpPVYaKzk3kV
rTINQkCvgbAP1macnF0o3aOt48bLIFYj85fG3VyxpZwe0xQTj8aVHXiJLy5S0D0W
dzrOJ4ecF0cCa/JySf/oKBHVMC/r18SgIH1jJz4ArIyHRy1c6IQdGCfhPTrXOZOZ
XpCVtqeQRiK793t1mfaRFX+DN4F/euRsR550jbzxeqFDDUZUOamoyofcKaJWB2ry
Jy/wolItLbjFitYZeG61j+EDiswqYPgcDW/bBVOJYGRspsqmq0ESku5OcEZUhwT+
7WZAN4d5n7O7J25m+f9Sia1Gfn7Cf7pF3OIXaDpfWhArEB1TPhis1yoIustx2bCT
4NRiFErEsWWLrc+ns4KWaNQtwvBQBINkNF6fhJKmtBJTGliZn6g6ddVcdeTxJsPv
0yAyrMJXTgYEAusHIRDADXZv6IwlsYEcAKE7iDIymWDuHxCbofgnPIqedRgI4u4L
nKdW09DesKI+cFbwqCat4nPm6i0cOKB0I26tGThbZhwMXxsRvC6nM83XQaFdNWxa
i/jlfq+7WmvlSJS4aybPYP2cJtvyoOaRIn+R6R1JXhVp9Twzt+Uq7DIJQUFHEFJ3
q38BK1HFzSBNbvO6/PVkHTNC/D+wFOoGZMPs9OmgIY1B3QJd5lMfoe4w4NwmhXuz
7djT6ZddFEZd/YEeeBd2oMfWMiKErIEsAKOITcKHLmj0Gl8qTQveZcj7hy/I9gPc
YbEcuublT3BejNUHMpH7PZHRhSkR1wRj2jV82r7xM9QGDcnyDEfMmVAjiOemCF8/
PTdZua4QwvwLh/bx9seskVpxcvnhM7sJdhBXUCHkkFg14CgJ9AXQyeQKT/IqDvEX
0JkS3KguD9iQMoIEwyEpkWoczViSBfSFmEeQdHUphqs3gljxGrxhk+EHErEhHkHk
O60F9TA/3wCgamsvZ5lraWIuZs5d92BrT3XYbd1lqU2lxcGklQ/JcuFWJHgcmYtF
voUi8k01XxkLsEDibv/2Dt1Q3XmPq+IkP86SRBhDRIX9ihJoczjC1yxYjTj/MMFt
NCdPoI9a3ruELj2LMkjJ/lEz5HZhbp0rDS1PK8xYsL8za+0JYKk6UpD0DVYQ+W30
nbE7b8yPVKwYkvreQou0eYjf41uWvSXB3y8QPU+Zt+jGg01+HDKw3t+tTsLteLmO
ApXWMSPeQRKs+aSeoMpwG+Dh6mkXyMk9mV+C9qBaK/8c56nxO6FwmSzNbGz/PjXN
ONE4xGyjz2FD9OfSS41+Fmdn9wcEYKM3uymrgG2f0/xbsO/7ZZ511DRx7JQVfz7F
7ntxn2/KWUY83FTsDLn4giRb2qk8beO5VBXKyf1Ss6uOl6fTjc1Xhsbz3Lu1Bs2v
M5o/vsEjzhSDEFFwOjlT5jpqSAv8mF5qL/55Idxbl6x34fJzKaEJDry4NEM1Nln+
gBN88UBaeVZtd+pLIVuyA1e5M/xXFQ72s4L0upEqc5wjC/9nYtowJxyvUTUPW38F
KnBFt5FYkStGaBaG0//Nud/Hd9uFMsIX8vyLrs7pqe9Yc8dVgJuhLa/WEhctJ/Ii
RYhp7XYDZncZgOky/GywhndonRtaHt/rOWXCgw896HJihqP+fSOFGD7QnyMvQNJp
1aUefh/aLJmio8/GT5QgTSs4XULf1DXHPJB05uV1MttrncJRtqNq8ewZlrxUsR2J
fxDrQWsQjk052DrXFmgN42E73zdhfEMrEEtDIYSEBztglixRsONSWDsJ4hIUCdrP
jTW8jJR4kVq7Q+kZTDJvprB78Q6ddt65M8qsH3dS0Z7fpiPLutAdyeaCBgaLTtM4
YrTs7NrZzlsbkzyFcgSzegx8mzIBaiMnPQth2uWMYkYN/A4EL0CdAlB6uSGSec7O
IZn1BfROL0cJ9dY/1hu27THeZ8JizC5cqRQR+7LOkEMhmVft0F5donZOprOBlt3T
y6Wd/1lyT6D/kSykvVQQ0KGoIhEyMz/l9mMNyQwKEch/L2PFVQt9XvS+VBeb/Xkb
XVtg1/AMwAZpmhclu2wnaYyJFWUTXH/RZZR/T10S5EqKBrrEREwRScGNsq9RnfvO
5iOWrG4vwMXHO9nK+1VXcZUtQnXuCy0ztnS6KFjSc5UtcjGDkR/NwUVSq9xO6R0Y
CQVQ+BnUokoBU5/FT0QuaBAH6QUQ/Bx6ukt58c8gad17mVV3Lp/CyVTXAoBHdKga
qiZ5BEKS4bHLEbHs7oP05o+m01NJSv5BfHYqSuvY5+RMCDUwwQIGlPMLCDqsvOrP
tvvE6CqYuJPVvj0Z97OsQXCWRrqJi+vX32aLpLeZfMcTwkg7yadduRhAfTA+8CEz
WB17Rlf1UcmV9tAp6aWgEqZnsiSH8jo6mTq29T9lYZxdUXYWEJH40wRxWEIw6e/7
gSl0QJE+43eAAXQwTiCyne9xaihHJfdjFXyKlmIIWbPeW0HKkMLun83SrVZbWaIW
Yc760u7MHMulWfPT+YRzvBDk8bspOy49DBSQ9a2X2NV3gpsjU8coqkFSyuPhK9Mt
0UpBXQIEXpvHLnvJ5RrW5OyOu0XImoaXdU4mMccHPJaDMZAfPRk8+Y2beB9gdcqs
7G6LststNRtwmwah8Y+Xx9azWt5BRZLt9dqQJlFO+C+yAPYaH5CuLDv3XT9S8MoA
Ha5dAQbMMVMKxnYPAYDD30TILL9Ng0zBFBJEK49AxE4vzLlNhRhduO6a8sy/EY3L
5MOjeAsrzxLA4VJFIfmCNF7WNmdoLkLboCa1K3pJkbebfRfj3pRo5ejkJJh5epU8
laKzEpTgaA7cMiWbyRgw46kfACNAb0uraUXQAB1Ei0BkHTIzsdv0rm00M7pNqLyL
64sMiFY2nrZUKIPmdJUroJVsoKGFEyA7COLZvYTRCSoDrnveDO32aPvibttAa4ib
laaZlQljXB7vB3dkh5q2+7dB8r2ip3Yursqtg2txZjTYxF3qVSxclixxOCx2Flp6
tRgPTimRS+5Qax5N6jQUDHi31aiuik+M83P2XQJqVfEmaGwgrKt+V6zlKcDdZx9L
1ScCx1fwDM+Fs/+GAP6IMu46Qla7RxSk8hLr/3/bN/HTox3E0cKFCbM6UhuDXK++
PdLXi6EqrDaZJcuVwezKu3adr/snRS1yfKZxCcmspbnv9uYJuEMZK5ut/Gd95a2K
M99jOKmfoI2xSKChBCzkwqJTCBDmL7slyaAhliKVWsrU9J84zIEGSfXP09cdJT78
U0s3S3O759hjGiE32qX7AfXpwScd0uehkSykAyJo9/AaMaTbH3xSWouIgPZATS5c
un4Mi7lWa2Lu0JE/JC+6s+fvgTk6DeX5AHMJGhQ2b50XES3QbQt7tllJ3PjOVKBR
tiGba+pfIlBLhx7ojwz0KrltnpKlbFp+W030TrLX04vw/E6rn3StE4q/GuUBnPC8
vx6KkCEwSCVFot/1ZBa+WtWM/B++wwzy0kE97VI5Ak6Et8AOdIvT7e/+QPOPkN9h
Bq306iCerg/dmruFJVRHaUYoNcMRTUwCu7Xy5WY/o3PNZU/0zwD3PHy/YC73qvl6
XxQBJANpCb8XhY9xUf/4zjmfvqock5ipUZFER3xyKjuSnvYm6BSscFn1tZAHvsVL
GZRmLdx3Gn9/VSxsgN4DSHdqaixflY3JjmbXM/i3aPKntNGEeU/0xlc52O3WqP57
iAmCwW88pEwcQ//z3mfzqL2YDUE/LMd17rH5PUlfO0l0ygHTr3OHHetQmm9j48Pw
7wCnBvKWvxiwTeAr0wbiuc/SWkWNoKIfQ7kmpUcK7h24l5ANS6DLiki/3JQIccUi
qcBU1q7QEQWpqtnkvM78nnpB+BCAUiA9gB9PwE8iJTdIFv2kA+NVfhKZd7ZZpdk6
qC6ic6AsRuviRfxFNp2GEeTlqx9UtxskPBZ9zitqBVX8bWjbnOLYcrzS1ANmbM9d
Dg9ZPicE/hPdeIeJvZrnlbtfinmkSwMxoBWsknM91yaKR/0hAO5XIbdceKc1bvKR
HrSbci+WzCCbzeiaQrPt3pOQvD8shDSz7u1G2MwF4SCqjWo+fjFDJwvfae8VNnEB
M49t4MvlRXqw7POw3WzGP3+8I5rZ3tfsZcQOKv/qpcXJNG/U+hfGI9cvJSc0OjYB
TZpnMRq/cFHa6MHPXZNmfdP+z8NSFu3wwe6lh3Uvkr1ID/k4xBe3GMebGzBRflg9
2raLDo63olwhpRaQ+fsbxJEut+oeoNByIy1dFs3IICPiQ80U45BhDFn266nK8HbP
DmZEF/hmaOl6yTWQr+Hd5BZH2ZvSsR8zkxZc68HL3+rljKMZlZkDyptSa7YATGk6
nvkxobkHJ8W95WckOTXSSlel9pLTMKBLpJuAT6SN4LyPs09o9Wq6hwRks9hzulcT
g8P1GidTxsINXaAJAgoXVkNTT5XRZw5rhnJn994Rbf8cqdfQP6eSoS4keMrmuV0j
INB51hMgguFaPs+PgRvwv5+ermXxuQbqY2nnMjer5dzOG/k9L5V/wObZoMZs8vDE
ahKEac97tmatNHEvYj9gHyznnKz5ahYT1PT+zJbN3KMMh/vgK1xarI2DFBKnFei7
kGK0wZaWCFBxqWo1wO8rmz6/vjiCE9qXNk5sazWI124KIntDFMsfQgek5L8TfYXn
wXQlQArQtk49VJDt6bDCTrbFE8XY8C5qzP4tIVtdqqMb1o69J8QGp+ucVzr3mVD/
9gQE0/7fSr61RjRWk4yCf3snMTT56tNvCKpcovUTf774F3hgsZ23s2gS1whAFzpQ
2g8coeNrIeYvsgRMsgazID5QZ8HHvJ6kdkIvW5Pd9ffjJ1/q5KTREC6TVyVEMPGQ
UWYqySr2EbeUuazs3xpYIfgHv/CUDj5KYCuJ/AwGIVFY0CWPM0OxVUXJMo0m5tfN
7LCqlvxUt09/DKcf9solfC+/wkXlALIaQ7UOAnRUMa8lVVcvQIu7n2QJmPh7HloY
RH3i93F2MqesfFWVO/68nW/82KpSIU6MOIbjvd2oXbvPKsSLy2QcHTv6pfR6sJJ3
4IPgEnHFfDLrfRGCBJCdyYu57W14hGE3PnAXE4YGau3Q0a/hxCHqXtaMCXAFt8wv
dZmq9nIvghPwD8uKQiiyy7DfppYoJ6COzKRUiZI1pRKAQUIZa9G72+2AuQXFkTQs
e2bp55UD3pAudd/cOl+0fyu6/bdpBbqkNPcSEMB0Kqo6sUPgICTEcCIzohuKzBOq
M5FqjiUbmJ/KksImTG6cgY2/s3Sq2qj/TBb8HY940ZpPa2S4KJmmGnUj39RbYKgl
svK0M+uHi1elDF4FSPP8I+ChilfNZKKp5T2ycRlY5WHXVfEWiFFFevvHUBa9zZ+D
r83nSsSBtYlvJ0ycXWWpST1jVucP3n07uT8EBDcgEmrG/GOb1S+tzepkMId9ic2f
n0s5VBzUW0ZL2RRHyfe7Ly9r+/EJ0ZVMnN26p2yhzFPLf9f5G86e8KYQr99qtauW
ORqjfw6Z6gL27A8xmin0rpzClFBfV5APQVSzaWg38sgD0JsIZdy452Hdft+ctcor
Up0FzsYvfxg9c3BtJsB2H+Zn/X1IjpY69+tVaX/xjLchA3dXo5JQBYJc6fwYMvSU
cH1KI3fhAT2qTRkte5yawMIRy+h6GGTwyO24MoJIjnHly4TL+/a2Fd/S7NeGCmFY
JHjyYo83S5zmln45O0YByRuxjEidaKnYVZ5XzqeJxfI6ndqb5rQl2tjx1DixGGdI
BK/ONdNN541gnA1Ai08YgLn8mzXrIAJjFHv+uo/PkqXT8hhc7LxaoYWMQN+AmNDU
30bUnbD87nOO7tLxuYFGIf97vU2+fY5houy9AxPEtAsIy525eTqP2VZOeuAHeK9B
fe5zHW/63Gn+A30EmRegyhJI4d1qqnHYW68NL4zkU9G/0yWXilVAnARdqXrPzBwI
gw8sn9wvWKPL9kQCnFCxuf8j+brPfQR6eP5y0PXOH05hHel3P9Fe0m1chK7auHBs
RHzQGA8wZiJKvjSyP6lO81OoYSsQYr8r2A/5R8lpEmdwwsw0hqWDwPqP+jUUTCtq
g8DEatdOFre/xF7qjBlvA4YwQql2y87Sj62FEXPv0zlGZuqFvBXbfCWTdDnjCBA/
wHOs5s9F3GB0HilaTGOmMAgTntAzbOLHplr9qBf5nz6mpfUlVzErcm01cOsimg0F
x3Z19BIQyET4RZXXKElFl07QpKUG/2YWpi502UgwgHL7Wsk5EsT+S2Hx1sKnMaOg
+D/HV4deUsH4fAXu0B7qZerSPsS9W0x5CeL7Eh7BmfQtXs7ee/+PGYspCufwgom1
i4cu3yHzcEWEnDAWo2FhNGbrAKCmH9Dnx1oQjrelHKnCcEk7Ck1JHrDJ5kh0FJdm
vOZnd5fqwWAivWKnvxZjc1YmaxoAM8Ea3wTTMdDLKTPNLcv2YFF2NfGtxdK1ju0p
0ln9Uk3RknPZCQOFIsN88fOw4K3rF6cb3xRqVz2MZuj9JypKoRcYin4HBdg6eA6p
CqhC7AAvlJn+6aU2tDNSHVHWtGoVfwXwnks5GQa1XzuYRKvIxfo1PQcXU+at24cp
ioGalWJ1YqqKsWNuTz/3pFHYvNKx4VYfhH2BbtMymUtkFyBMToSRJu5xRUiGyr7P
uCj3XgBDsFFT5Uin4SEL1+DqSdmXlcilD7hj9CtkrZkLxrYWVhQgZrWggR0ZYml9
WGz9Y+f37wBLo16QiOsnO+r8JjPETmeroH+/5HUO6JMSlhGuidPence0mzsFCg1q
0wHei84TExxws/7EBkKg5MlrYFdTbYSMQ+q60Y0MEY33fjyapPSoLOhr41SnM2WJ
E62JKkHQ0bDs/oHR8VRpITPe57886DxLiYM8PXoRXs95fWdPQv0CrK9nDLDVg2Fy
LrqXTp5cFekAKI4sfXLhi+n6G3FQKdICCHpuwHJzyD5lByx4EZ/CrfvF7Ya7+Pmg
ADBAQx1iyrnJTRL33iOBkSxg/pnghR0ZRyFUlnlwIkUX4AKTRG7nv6c0wq/Rf3HG
TBDxqCsJRCKh3fSmwCa75z1qKOMgBz/NcBrFaYKutHWbLBxPSSN1zfCNlXXnY/Sx
B+b8yb2PyaW3uduT9eKF011xIPGcyQ4l04mBJcEUZWH6Ild9oUCBXVEX8LoJoqaa
RSpOHpfeI6GVQK4aQ0bZlzZpIiW/r3PIDk7xfYKdYTA+StM1RH0v5SFFPwj+CF22
HaK794E6Hq1J8CYFYpnCg+7+aQB88MJWqBvoNVr78JcgmZ5Q1GFA6YCRlEbHVBp0
MHClQyuW7aJtYt5VjGq+/9Z4C89lda0BNejJ8GgECE6rKaIL4xelb7+GE9N6qBww
sAwauWH+yRpTlmpbh7TFnxrma5gJdun+mFKiWt6YI/968JDvf/KZS/iJB50zEZE2
3ovbwTvrn7D/FxNTbsWfqKZeDi8GUH5kbiaFAj3ddkAD8UowSsARofBgUM/M3G6Y
/Mm8PdEu6g/paO+76pELKtcKdspsJjNov0zG3A1Drk5d2drtHutXd+MSYB6g3N4B
skoF22RtQ6PdE2ZN50SmlvKD9IdCENNKGhvYCYh/S//6X651eXxOZ/BgO1XdheJK
cgHEgAxqqpKp29hydZ6fCX+n883xRQfdRaB9W0v9zO/gyQ08masZs1lrJGQmQe+N
AQwK6Qc5yKtA1pzX/p44ji/IwCCwWXauWBMNi54Qi6YtbDzgDDqYJLsq4eIhWgwS
KhJUaTPQjjeCreE3LulZRh06YNfIYItJ8OotX3uPmYcAmInrH4o/irI/faPzXdzx
Umy8TFaD1TwhYCDoCaSJ1irshwVHNRjjJnVVsOJTPI7zFWHJiwDUFd7HyO4G4Mpx
aGh7BtmBoWrFbtQLjnFupIh9z849ewYVn1fuGh60BT1hd0HM+/gpWqIhaCKFw/5S
iypAHcfmdNkxHyr+s3dXlR6kamZrHQO7nxfpfVBiL/DJeRQL0AsES+BFvwAlKHBP
fN1TJL9GfWNYD7p3BrR1AHpkHcocCbcwB4Nd6z1UelcP/0bYrBnhydcqt5+0acLs
xh8Zigufczmu/5v/JFjkIAVE5XFjfNTd/qusU+O1qgJno2P5Kew7h1BSlzXGaL13
kod5K6P3r6RlV9srRqkyzc5OhZ4YOg+fVsdEAcOEB0DpeNoqh7NMCOtWUiHU/EKs
tlshvGEpMev+8ZBKKw7ctxu3kb1KlR2zsAsMs1eEDiCY0O40hOaFU1ms/GNp/gfh
cyZfXZfHmpGvzmABSTHzS/C2kuePzI6j7OJa6djBGRbvrEXd0gg9vsPd85GA4b/U
0+P72T0HyqNfPEuTnE8kuHAcf/kWNHQFrJHcbdDDHM5zjJWcTn8WXZUEkR3b050s
95ZW5b5kEqsl1v6KNElvmDgZUyZREH/PApalGHYs7zlUYnp4/x+mzsXFbnqpCySB
CIx0oJmvxyUywbbBcdnfZxrlSWdBpc0ctSODVaW14VYg/k8vcakgzvYNIdYWhY4j
LoYuheotyaQEfV2rcP1Zaztpm2heb6nx7tTt06+7u0R+BHgZgnLfsIvAfhP/SVs4
2ABLpSS8x8LDgu41LRWkN3YSuX9EChiiuuYiNZTK9MvEOnYNRATJdzzE7A9TVRun
mo3F2eyfTaQiVkPw9mBCnzLufO+nF/kUYTRN3p22LfXEhiDAbU62OwTzxuUHW/1J
BRrieBJLU2IdcaO3OPhjKMUUT/8GpBTAspdx0cEIwZvRNG1H288yJhZYYlQmyK8B
DB1CjDnz1SbgBa5MG/NPG9apXGZlji+imMbqRGmG69arFSAjtTlAms54TqP+c9Ev
tYcc4hzBrVMHHxQ/mtgChv9VTWbsr245dzGxxmXo0WYbSIxNCIn6yQVLt8HY0Fqi
6gJtYZK9PZtpdNg7q3rvAeTiaQsE9PJjefJXW+SsOi09tAGJaBLOkMJWtQeTFPSR
MsvoYBwD1YmRFlO5RwDzriH0cPmCQsoPgEo8oHMp4JeGuYRpC2sUC9PJ753DMeI6
8hqBTkHKUE6SP+wFO2Yei+UkhIzI7HnHCuCb77aThoxxaIcxfUgMUr07l27mQ4Y2
4r8XBSyFo8NlTXpQP93K1KuQHmC8sjvwh0XAV7cnT18galDaFEQ4P3z0O2ciMKKx
h9vF0SHCBnEHQeXcxPhul2EdfCg06woDr5y6DfhngPwQ6U0dLGDWaKKWRH3VbJgR
V1FlczZm3Z3/hy/72cM33BTqo0dEVu3L8yIF7P+y7SpVzw3kCEmBBA5BNmmpnvMM
eu14huGfgkb/LpWLxJzigfe1MJWDicPPk/xatbGPcGthxx8EPnWSzSnHSFwLS4es
H1Xxg10kV08fGRjJKqjnM0CUPN9gwRy3Pa5QtL55ubOeTs3eQWAFBTsb6P+8cbIm
e9RGsCRb0Jvgtb+e/4JS8rfP6BVbVYfEZ01NfFNrHQ7M/seue4tv7U3a4mVlhBLE
pMyofwaNuduoIZJkJvLwkbOrZvY3KgzCksEqtFeb/8kcKi4Ab50FwR8vSX3pH4E0
J5vHTSyFCkSRGwzerEsXV9h08wAeieRjiIMAKhYYECaVQ3/yDyu0l0tSes7LdOV3
qsPbgwhJ/1NcLTyoCmJPyeOPTvJUmxim92jkix94P8U1rwbFZ0rpMD5O0YMTW8/V
d6Sm4OG6ZMqSwJ/ITielp19uPOM85A2l5AhTAckgmpDDcrpae+95/coo96p9lird
6MrE+c0eZ53o2325BccYAjPdDEE6TrJnDnX0uHrwU6fLHgMWK2eVDkhoQC+5K30J
MDUX34e1UGtgw9M0i3KUf1qqK1oMiGAGfa51Py98sC+JVjyH4hD85HEUP/eIC7WE
Fmd9paa+qdgBckl72QYbWdO7B05tY/XLqP+HNLC7a1SV8/QmQS5iexfjbNBsB5ng
qIDGXy6npRtOZf6nLjUB/E2a4w15NNc/bkbfZWPUwhucd6A61XRznnPh9XjmJfYI
92UxbBAA5PD3cI9Z0gRpVYq5mgrUp6pzIfK9HT6o09LWjFbDaZxmIjZIJOAKQ2oB
791KzQN4sIZraTlFE0MXUBGR1UOTv+1iGLC3gPgfKQfS0fv97qn05VSSnNY7lIwr
lOycPFYfpMjMG197AbdQJvDytrR6TpBvxzx3tPZHcT9NoNzPKjf5OF1wJovsTLor
7ikP9nqOD0st0OlRLbwgfWqa74z1YV+uiy1mwsGiTCPQe5lJGZ4nMt6yfm5KQxFd
fs1g9P17dqcLMJg6SjKlQOLS1KRPr1YzzR/IpFerz2KhGacry5koftrF5CfObrf5
uTjJQHFMD5FpiW8MOtUIHbcRzYQ94y57becQHomi041MRZY+Vs1hEKdeo9Gj8GH9
4/V4JewIaivVeKeEhYgu+dyq+477k8ij18wTCiWNhNXIiI6LsGNHJSNMXSn46L6P
ZO/vUa+H6kPStQxBdRJtmMgq6rds5bUFHQ5f+o5q968ecWx5STqnA8398bK4hyjP
ScRPJhGddcAnjMujGr0yfJ/3Fax+Zy5mFOkuywz6O6sKsaQ1BZ8p9TondXzC5DGO
fxF47etIprq5bDfgHy/IgZDvL83cwgoJboHHW1AtTZfitGprQfwxgkpO/BZWaC2y
cu4OvzjgyFQPF9tMdSSzBUuRCLvSPPvsiOE0FvZeA1HBwYalCBnCwZ+4mgt7x/sk
72gmq/F6YTFKT5LWJgPktqTx8zfh47f/9Vw7Ycq6xS3P2jjqRCI+rx9eeCunJO+V
BcU13YO/8L6NbxYAf0nMWF4r3Uv0VdYIOPY4jphDXCjij556f6lHcHzSqwCb+El+
mJ3gGkJZLvXvBsOiiQ4j2SnaYL/N50rjoTH18Q43pLjYuUn+TAv2FfrtVqNUCM7g
TYGhwbHL82nxihSe5UHTfnKxJI/UuCGeLzN3bFA3Wsly/hzIThihZfENCoJFdfwy
wdgbj1aoJKsMEg7KgVbcMmXQzxkH+ed9jWqNA4M0osSGPdmode1/fmA3y/Icx1bF
6tT0Ht7MwQU/o1ucLsH0ncwYDlpotHwCsIy433KpCvOurh57YbG5nbYJlEQ1N6CC
1V6ybA+7I5FC8UtMAe2QyrELf3DQVyVdwZS/UbSwmshgAdYYNTiP5Xrnc/gkMZ31
z9Yx8l2pwDWK6neOBAn+PpnP2e2ch0iktzNoXnFUf4eqoXqpFBrye1i4I+A3wg4K
chuoo9Qopi93DCtOZ4QBuS4mkRuJYYBdFILiiJD0ZXJm8bmG5ab/PjEmhHIIVAV+
1lDIzRZKvKpzGKzw7RJpn5Y3EICYf/chVRaYjK31SiatreBUI8oBwd5ro6rPJ4ui
xtOwVipsXzjneba1M7rFrUoP8SYdfjxeLU8IExXZVQZwHuaxf9e9SMXmXtWSu+V9
sRSpGRQcssJUCN1bZyFuYreG3Etohq4E5IECKJMWqeNjJ1T2FQxwLjn+vcvFwX7a
yXP+nF6lddYDkrElpv4DOg0BSJx9A28Ly+VxXPC18G/En9ncDeRiDRU6c3QEO7Dg
yMbTJBcG0p/Ldv1M/x7nt6N66ceZfMHw3hBSNIhhxFNzreDU/cwnb3GAwgvQjAsi
4g42NI5buSc3ku3KfroBevS5w0v9g4OZWCNXl9zHrLhAntm+R4K94H/+iBaUhMOM
NpH19IDymJRpMB9YRifLbY+X3ngaz+g37vEa9HbaY/+KaO3/Rdu23ldNAlrTUmDM
uHu+khSFAhMv4qxZM3QpiNotVSjCE6jydFKBP/KSNc+/phkLCDdhT+1ibyTNLKnG
hmjYND2uucaQbfw1XRWIO+RW+C1EXJ9JwLgDwjiAT9RNg+qR3xLNbQFdZGk4Qqri
lvj5+zfUUvPjF4N7Uq/wLO2xlMP7VR21T/GSb7IUxG0gTkzXv9dCQi4ZC4TC83O6
JSoOPpcRh6IteNeCF9HPpGQkPi6zLKu5VNCP62Ypz4HmXtmAPljN+r7O9gyUuHB+
qeZDETbKWh+AdpdCyPUEkFX89qyrA+khXugCzeod+dYgu5fONR67TTxk8rH6MfWC
BWk9GEsGIAyCADN/DZoz8Qc+yorzuHSSs2Omrjlfx3k40nTQYNhQaACe2IAT6j3u
7EhmAzzh+4kadWGt7Ija+3f93VtM59+yIGdqbUa3RNfhnPl4ewTG0RkvpIqLGX4P
V5W3oBLMyQtz9Nk1oCBbAwChuiovBIpOd9zNDDXvaOJIYA4L8NCqjbCAw++kWw6C
ZO7LKWrFajjobmx0ioqzvfEBMt6grcs+2VS9myGXEoMxQEp2Lb9eIxLpC2U4ky1e
+QNhu1r2ScXO5BKUJRaCFbxHP6b0URGEI3XgBVkDzvDK+7wW5FfkGCKAC/DY5YZE
P6tsJuycVC/ixAKKP5YVP1fPvA2IT1Ydv7QdEo1ZgQmVDg7BdKjpjvvfaDD4mEn1
LyguKd7Pw1k8zjwVRknTvPyGGWBIlt55gNdOhKwVIJYUmCE9gSeulZm2Ff9dy6sD
1P1MEs98u+9xAGo3Jn+3u8We0LK8KFFLWQWnmMtJkGiZpacPE2VNhZx94BybInxg
u6KFblh2hIoDPWSDOZSNiuY8ictIRHbqMJWWwGc8qQCVLG7XRRhLtCM7dS8kSd43
q9PXFNt1L4kmeEFYXlZmcCK9RoN9x1A9QENJSnrxuAB/adrq0XXwp1nQJ3LdfFNF
xGbUbDrkiJd3mX48y3+q5ndQakUBmMKDICf/jv5wfYBiH62lERYB0uZZgiASqLEF
bNm94rI97ShoYMkKnb/cGSFDxI0F+DnrjVLWX2gjtfY7oLmQtLjeKbXtDNCF/xQE
YRo2IxfNRopxzKoSGIu5O/XMOvjp1+jHaR/yOxG3yG4w8GzQzy87Iu5psYboNKfF
157rnoGMtw7i6V/5E+QTLgUt164+vaGrgMiANK4PmY/+9BHWqB6Npr1HJMEnlTAV
bKnMVVZv7xXFq8EeznfTVk3O4qfxz986aigd0jzavmWTabGphGA3c+2d2HO4xJ89
/YrrnFU25lJi09GT6qj5RsoC5vOtd1gEpsEpPZPCvM5onjEqN7odykQm2zz5Pd61
cb4JocF4g4s2RaUGz/jgwpg9ZKWkQSu52WJ20c1atMHiHvZE2pPAse0mTxLqlMWH
YpqHJzMi7y1SlT4GfNAdqEDNpsvXqbKHukMvbbaAS4YvvsU8Qk49/OMC+vQaZ2Mm
GwIfv2BlcP7jhE3E6dyZVD+v3rluyClCX457/6pCf3/F31LQ+76BoQfKBC3B3npW
+YaVOK7XdtAZohmipmA9wd52ea1gsF2FWntT5iTonWvIPIyGdEaiIWgVrnB0LENB
gL63tu0V1r5REr4YGcb9Nh6mDZJ6rWfCwjmmjhnN3JTRz3ZBt0znYuMVXiA1/6Db
zuJl14LXxLeeK8lG8GPzH3FUt929JJINi9A+bGSQhV1z6awyuXQ4dfBoVNaFGf52
dRRCeOEA8n+oNYUCdW6v/5Yjxj7UgFT5TMHxAfoFa6gRDaHU0LWvhnHen9e8NqUT
kOjFIZZK0+JvK3+QkScBTEcaiZqYIJZY3ubPtBwB0v+wRMy78v5Kt9wL/hnbGWtY
3XrvVcOG1Vu80ywGI5DCPKP7CmnCtpUjT949RIgF7YRAmgMdimhpqYTcC+ciLeFP
jVddRRog7Xt+GofLklhUBzwS3JHfEczlTUzVxm7OUPm/Ac7PI6xwAVxo0i43u8WR
Js6y7DqXnL2udHraiGQ5qhFt/NFrE6ZaBrykA0a9ZPF82m8hh3I1NIB5wboZjWlf
R009cPOdnjDci8+xTZa8X1lJNLCVikVEuqKgQ3/gAcqalYt03BY3pKqfRM88Md1Z
zjTYcp3eZ51ejWMx/YGt4Aw9GrGLX/UHEMHKBMAPyBoehy/d5iGNr4OJMTVZzRKE
YSF/cKkVxQ8jSM4xqtHEWllc30Ww5nIh5dV52JPNFjM5Di8TkfnVxnlb9Z+201nT
/DVAKvlEX5VZxc22jmj5+Po/EEsdKKWbtwYRuNiH9iX/NaJ8BJmTW4pag4Sf55wG
zW3TO3X4oJ1YsIBdSIeUCi89do/JUJ2rdqoS31tHlHGo6GV9L6ZLrVkd4gpY04JV
gv8Wuenbkat6qB3MKtUxSDXJdD1AMaXjqqRST/Kg5MKihgprDP2s+vhvYo1VpRKa
+i6W+7UK2KbwTGchKx6tn8TDecWXGDOAys+npIc0sBija4+Ur70ujKBoGqGadTYv
N7WNhDKT+GdBMBRHYF70ZkXkFt47IILuFBIUvkwgn+QA6RawAUG56ffbA8Q1EwIv
NjxRtoC40NMy4xdqfFI1Oc69izXq8fwEo13cd3YpCMjguQw55IWjtSNiK57YeIvf
IDsQHdNwlNTQjDYXSkpyMikt80riDqpZNg+FxGCks2hPnARKkTeJdLcoa1FWbRaT
lMGmlqRyHoMvHEzJY0BFQHrhQTxQLlHgZ01kfh1cmC7GGeJPrFD2pjoFd7f3+kw5
0s3aUSm4cBrLidusKMjlUOcC2R15wYBS/KKUV4eaab7zEcEEKmiaDLJ02MK+UhXB
nVrmq3/w3dnqEGAVAY4/5c+YwOpxYWcQxA5kkY6Ul2+7euFHqhBNA68Exvy2vHQy
FbDfTPIo3vMsNyKu634BVifmqShVAnLXOt0dV8qj80RzVUn2xdhVETng6oyNrdQU
Jgo+xNvijUhL7n/5wYkFq4MK6gPQ9yXg+q6A5rcdV9+vharh6E8f2XpLU6O2FDqr
+0AN5N5NYqRLWu3fZlEKO9RuSwuYeu+pj9lgYJzFwOVWlmYdUBHYFz1dU2iruLuF
v36E4n94iNCVuj9gtkdMDtwn1kLBwbw6gHh9AQiM4VncwnBCMPVBVOFWDhpMpB2d
+EyL/YOj0HQZA/TzYEX1cAEKsvI8YlKAek8tbsv/xJtF+PAXCkDpTOEQiZ523KKh
2EGbVp0TpGBWVypV9oMF/oFI7Di9LvA3hHJHoBXftP7iLfbhlTbNuCt0MyqzJBqG
iigzmcTJcljO4t2CURSaheKpE3I2HC9LAH/ui1kr0s79bN6rnBsJIikjbDVQTUzR
u56xfNKijIShV6vgrCPpCdicOfWEW07WdnNAlwElk9CuMMV31W6xmKeIu+kninfw
7Wddj1ZqDzYzoCJrG9UYVKYgoY70x2d2BZjsFkQnPuQRJp1p8mwEDvTbAAtxF6e5
rc2hZJjWtqEGYLvR1NcLCILpnrQtd9iPT2IfGAnm49Gh+3b6ijB04F1vCtey+apt
y2V8tO+zKxwTwYf6qKaNKpB56AWUYKngLz4RY1Y3ioi5L7O62IVYishYtsJgs0th
al+y2UOcDqDbIE8dXpC8LP6h/9V3kabwY+8S82EnaqCk7nA8WAargw/b3UwgrQC9
oyK1yNUBrnlAizJAIJvZSclXWSPNp6Enjo9osfapfpTEEJBPVRD+Cwu8keo04Q76
VTCWYoUgqMWD5MdyRLudY22MRnYrqCZA8OqTXAr8IDxREBNhN1BKDpjlrjpHGgMM
S3MzFsQjbWspZSnEkhM/ZjcJOv6C3uFYzqxEboyEbkQWp7fvFg1ftfTJSW8MOj4A
sU5K924x+kesCE1k2UyNptx559h38tMxYSPpyWavA2LfKWDkYIwmUIWa4CSSTmbc
04Z5VyT5XRiE0NLBXUh0RG/7V/lVMYVx5uQKIECcqrrS4cvklzgjJ2v4t14X+lIw
sHIvlmnQlBtDanEtG/5XzM8RWiMBMQRGDDCv32ql0co3+xzeSVAZ5L6yO1QWD7gG
jVCYtl8rTOTtOE7kqlzdQuK7foisHvvzNQ2AvnA3631cRF8ZCYaAHtW+aF+Yez0L
bEHaz+5EpjcFdk8zkBKH4K4HYT4AsZbxPZcbYLn8TKPVSOpyMSpfZ9WJ+4QBRRpV
2tOlyg5N7Nl0VXD72SYspYrkqq3NNRReYgfOEKkWMnagWMhL3dXA3/wfU9NKhHGE
85KRvs5UEWl8ZKlbaRMHhMQgLM7E4DfU9lgBQ9Y8zHNwrK6RQ+/hze9Ht+rfPp9Y
7i/52g7NzD6t5/jAAUBFPE7pavi1R80QBbfmhO17MZ1vpnvqZDjs95BqJ7TryBPF
qKosGlq4Dk7L/RSj6wDJ6Ud3P5PJAHEANCf2lgfmO+87WG4GNpqDvLTaYi96fQqe
6DquFS/Ztbyxsudxgo1fcAy0yv28i97R2FaQ1Nv7nam/pLEexv6m6nc+54iQ2bcr
thMuvSxVL8Qg5VQdf7UT5Vrd6ZRnfs2eczsjTXqm2gEmiWvIlwpz5N2ryHUpO7CD
6XCiNDwxWfYWlu34NkdI4jl5WZfQvZFEx7dTx+iEgFMG7HXA8URPMXeBEuo9b8XV
fL6d4/8oLUBiUNx+3BTpypO6dOIx7DqOgujCQPdW6Ib+FmT1hujcfEapTR8r4vgG
bJ0N3xLH3R1SZ/0HEaZK+NalPcUBC0R8cEDopAWHxfoRn9byHYQVfdehuKSPyXKl
c2JXkX/dRGwIE6yJ85dxth9ajtFricMQuQEwyk6gy1SUblOMrBJINJVvAVJwc170
Zlh3wp8ILVLc3xrQc6VxAoH4edF26fsT6dvsXnzbpqgNaB734eumMqSUZ49QQ7wg
xF0BEaWqtWhSYLshN/CWJb+EofrmqXThbvEMD815k83l6GyhxDW2jJYogmcPotxD
5kwpdLLXYCO+gFESLTaGgSm23tRdZyZsRS83VTNSejw8cjhQfXBPLTsp/1gJ2/kZ
l6xVnYmgVHfnhjjDE2xfh7sKzTV5MKIsZonRfgPBbFFUHloADYpXiruFuM0nxuW9
ipVsSNegbTe+e+rMuwA/LYN9wQ1AuQCT8Uzs2T6jXjPIr9llSkRSaQuRVCqqR9nR
eOLh84hwJ9Qf8Uf/OpIZtJ69S98ZGLVKc7ggd6Tu3+FgHHf3oTiVeWgMLJefL3zV
WnY7ZjIqceoP5yWaOPOuhF7ZqHJZWnQwdiSe2QA8X+jMJyxyhx557hszt4rqtb8Z
skiPXCm/qPvzIMoWJbtZfPqUzecf9KFrRZePuPEqhmZ0R5mREbXyGBJnCPVPwc7N
nyWsV2b9d5c1RebFvecQdDHDbTEGH9J+QofE4r9vQidzzwW5dxWfpr7ToYdyWM7L
fVCbP/pDbIUeaDhxPSEKLqWVG/Xb1CETFpv/ZF04AkCLRRPFJcDMlAq8dcul9XqR
Vr8nWi7dbRmTS1ot2AGCLD36ZwaAMQfku5rAJ1ee8xUd07Twf6E0VHlL3kE1afVS
UWjxPPN0qJdM9Ibcm9Qj7oqNxfMXA2FNTYNexWQrw5tfE1n0g+mHgq84fsevCye2
WBiDBeaw0ZdAevz6076rQwINMNsXD3hOzOp1gWZlkDu6a2rYFTiToSWCVqFixPDy
dgAJ6Y34Uba4EE319cK9G2Ml/gZB1QVdFVGGAOYgMqBnD294dLxN4q+EzNtil0/9
tsLa2fjpXkdujh4/kw8ksu1/TIGnFE3BPHpV9O905zsgQE+uAs1nExB5LXcC5aFh
phOAdgfwMCSc7CmYWaqwZJzW2HoMG5yuDABoMKDxB+hUyd2u1sEwch7ygLabxbnc
vFLQPgiJ8PLtC1yPcZL0zaXlLB6nW7SVrEQatNxxo0jdcQhpkRxA+iewFsUi9DPa
QBkQ/qv9WHNepqQWn4pRHzG0uXbQP4TBrAGX0LLLW8ly9l2YBABwTU+i9v6QqdVF
6mJCYcX0MLw/z0XLTJrf5FGG0+6OLaz3kZCKFIrU0hzCzq/EpPMTNCackM3Toox/
VE4O9hde27JP199jkJjr2pLcVnaUYSMqsRgKrYVvAG9h6DTrttk/RfOxwbFEkKG3
KVMk8Jnb7Kl0xnJ2YYNcH6DBNvM1TRNORaaAXjdsU6J0BxOKdXOJPJW8ghc4YCWo
xN2Avk2WJCOqn1lH9u67G09ubP4Z+ozVpj5j57Fklz6eOChpFQ7JdKKKDK+uumbW
wx6hfiWjUu5sENXsEcbCBn1pZpToblaf9lEttBZJE6teItRIPBsUvCTfsNa5Z48H
ZKAENPuLLRCQ38ansDidzYlPePia0D9tIr5/HpTQ6zbUw1wedCnbMnQmegOHDZ1R
b9CA6/hWLDFnOdts1Mk0SmHTOF5LPRX8EuLUQDO1r7tvpBRMyfSET5+l4pC3ZFYb
5eqmrnSmr6ROHLIne4oKa3fPVf1WBgqmmUAJg87b48jDwH60OarsjpFe6bCQtUNC
3HBIS9EM+W/URi4DfT4d9UKXINz6R3KHRqk6Yiiw/OLFX8AHMLxFFlNpozXv0hkd
+6CQO7IlWe+F8ZVZT0qYZHWtBNL+YQ23J4voa3gzeG++pI7VesTC0I5B3im73bhM
TNvrLwOcbRW+jcf3GRUDi6Brthy36oWuVbhkzN4/X45n/+CEIzYyhOXHROQGOJc6
nexmaTwOjizJ6RO4hv/nzKEdN+0GtLE4CaDCgnCMyKGNQnQwOorPi1ePZs5Fg5R/
NXhk1SAm2PF1ceyFRa7LnAUeoktQQvc+zilFYQpmhmBZ99VngViEXhAstewpqSYh
mksEJvnme6iSJlpqgELaMNdAcQZTWgWwvRoTCatdMDmBTnC/YRS6lBOyplB09ynU
caK7yJveYiylib97Ml8MeC2WnMIPxVupTQxhRXZ5POxWr387cQ7hio4JP/rF+OMS
Ii9Z5EjTXvFwfynV9u8jvrhUxDa2pGuL0m5v/H608WEptf3j8HH2YWY7YKtgWO6D
XtBKhYqZwkitZG20KeQnXaifaZXc76jYFRG6ZkKGi5muoIaE1/B8DRc5UTQQcKjO
TN4gPoB8oDelOItJTHkJGp/T/r/OGS3NkYL3wifkPT/GUPH7ITeNZqgCXwgtNfZh
ON8gMtO8CRqIbMlGTKBzQ9lzZIGI66cUzuL1g1VQ3vj7dR4gyphYwo6iP652XIjC
wS6Yw/f5h4YtpixjK3GxQ11FYJp03OyUty6NxjhgBBQZhMn+ZZ99UoCywIyTRsT+
g6KmSaF1d1LbXz+KYx1jCRzRWqJeXDLHjFzOnmfuLjQuvMoywSoIraeVfIRP6C/c
r3EhMgf7TDUS/XrzYTbwqxmJefrmYXP1apvL/86FGMKA1RyKxwHkcGO5wvp605V3
MycWOl9VXu3tChXo9scOc8w24b9pkZ2Lf8rcfGo/ruTfxScVutQU5iCbJJTwVvGb
sGht1pQFcrMTTwwSaeERIy56AN9ma87HfC920WPjZH9x9t2tNeEINWWJHKCipmXO
qinyqDvuRa44yk7S2EeGAqP7ZHqL0hfGVaaSykxqJ2UdJZaWzjRzXBCmUUeoiXqD
EJCwKnrx/KmzF24DBfyszGjQDx5JGe329W3XHI+trDtlO25XJf7PwhHhEeUedjYu
DPxCuSwswtPb+Y/c5nfU50KwQhTqRM63TRFAc5ZgbFreCGffLEfqjaBkoicZAyM4
jhcPpOy+KSc5GI7pET7B2TWQnr8pNWX0QffvWs+LZBzK79CNBQM/Y+nI3TNm8bvX
bFHxaWVmnIjBnOh4TPJyFVU3JrxHeet4tDU/aAZcgqBpD1C9xLb+fOGMkIGIIE4c
UstLbnDxH9fplWuAh8T6FNgr9f218jKikoISmF58KYsVKC7BtjDfiU5Luob3KHsp
ioEakuk9Jlcbjv8rugsPiqCczClCKb22dVkN6inWjxwBWazmVuZWKLHA5wCsJ28R
DO+v0AD8/byVaEaAw4FpxZsk6SK0p6bjnjo5VR9wkSVPl9sJJJhrucZb4PpEVNnO
rjNlZaao2Agb+MB4W35FXo5gVvva0PvRqy/pyFbS3klSfZDwjixoF3RD+g8IoVBK
02T4xDhUNH9DG4IrvJ7IPDqqtk/z5kMmvTpfQGyMVzcvDA9+7Rz92vLP5QtGJtK5
Q0cK1GWBkP288TSsCXzInyk7gsQjZMi6ZbG+3DXHGwuwc7OWakh0eZ0akNLmW7gG
ZZM76H6GZ8DB6PPc8jf04Iq3C2pFwcATrb6kqnl3SfRqy8k/WqbkvReH2E8N/AbZ
xpmdr5q1H3vCpNt6+jY836XDjnKj+cEaAFuZbtS+Lyrpd+KjlExZaliX6lWLafvm
YuY2zBtYHol7nKm+u43xbAZjevBcFyvER5DxdFBQ+rwblDzslc4Ni2Smn6ON8Mvd
hw06UNkHsSAtBtbv/TRsacKBRKiZPLjots7c52aKe7gy64wDvm6iqtDhVUUVGZyx
wPEL3xdH0ZDB7hA4f3QGeUqx4seHCKct1V9DqkSdyCiumMJWWNfp7fmDsNQwbJsG
9pAN130Ud4cnzBVdk4cF9mTyisUg/kcJ9I4yJszMORTENll8cyN2EtvW0SQK+9CR
kNAvv2gnmdoB9rrTXqDOAYP6sUOMU6XR1jKRpvqhCQvrXmSx+6Kb5qafKwZ21Qqk
+1mmB8FqDbbHmxYB7izuhpnXP8dJo+pbDQ1vuuIrBR7/2r/MgbvjXMo16801dRHT
U5JKUWKlFm8LMRcG0BtK6iC+3ifa0sgqsUILO5J/wZmvu4Efh/EJf62F3O4BI211
8IEyV/0psQEpppMO6MOdIyhWb9nFsnJ9sqCghjdxRMy2j4ffEzEOukqkRo8PHtmV
iTzwqV55KFa5mobgmJX/c/hZk16IWeDKEQRDiMC6PuhozpCb9V5P7TBbhskN++jt
h5Ot9Y5T5secPTlpRpnqxt9lqwYFKo/cFPWow0Fjh+6FM0lRIb5fT8WsC+nBAsap
MSeLqLdq8K+/pOlMXlhirFUfMj9RFd5IjykEai7WvQaudi7B+zNeQCozzZq+rmGN
yn9kJUEXiwmOx5LQkfg+VwZbd8Pc77nDY5LKhL3dwAFpBrTr0jWbV6z21+rdl+0a
nwNUtLEJB1gOXlz3FED9OXzxN4TVvr962/U+AjKJUsqvK8Tq4G3ekzL1UXic5FRD
3K2LIJHIKFM6dA6echgpMqR+jMDuSB5TxJCCkcobYy7gSgSNKynMTp8j5EvB3hsn
0Rrr9XQBHkkWTDY0VgfKcXNYAwBO1LiX+LwpCrtspkYNDP2daRA8qSKHoiFwYk9T
/1COtuoizexQhoWTJegsYFcGxRSuLOwmYeOZHeB0z2XynFtszKieWaOq0iVUNdLT
ACCxy1fHsfCQw6Oi2cUK1meAIwa2AEE3dOBUTd1rcyggkxh0srQMecWfb7PHfH6N
lzVNZi5jniQHpxaQ8+a6AM1pMo9H4pJAOZTi4QHGaMjjmLEtW3+yXYqc9/GAQgi9
1oOZVP2VI5QigYqDbLFdS+S2o96dvbO+drA5iyhK4P3DrLZLlKp5rJoZcbmADgz6
jhypi8s0+8EdjaHSjSrnolsJpdR7dnFheKzOrEmB4emeEcc8RRV4nmnFGxancID4
G01AoY7+rFsVGY1iJuUXGfpq8pN25lstvgeMxitftd9evQX2HDO3zP11p732rgvo
3JNbmEKtJyRLGKZyiU6In+Ab9n5yZrZDus0ABKmdifrJSWMnVHqgbqWl00CpOC16
G6/o/rb78rwtlM7+zz2HqE8SceREpPM9dHIMRzSccvuujH7e/oGj6xbKN0QNwgNE
/D4py+sb0LpSLAdnhWMrPDkCKXnN8yvgpffkOQTGBlk9sxIHmMado+ZMPjntBzga
6dVvI6P4yqE3A8eZiDvX5Wiwwt01rIs5Ec1rlyz46MMHpbz6YW0Sb+l2+oQxhE62
WLmtX8lP7rgrAgwU5DmL9Bmm0+XH9KPXQwW/LAkSjhxKBFzJe+NuAKGysl+PJiDR
KIAprWl2sg4bSCpyNxD+eKQmBvqjs+yWTXlMNRv/k9SsAECNDECZyotCNCsJn8os
C4vb4oDXVflapytQyRnDcThQE/pTuyqYetAJzHKU+e+rD0gPtypj+taO9h9MJs40
luSNGInAnqSt3y7K/YI0y+Ij1DOO7k4KtFd1VpkZb3uyFoghG/2bHpn3IdXOwCXa
O97BxATN148j+3T/HX3mdws+Gn2m+TnQauQ5V5kMKk+v+Lcvagl5FrQY7ugQyIg6
5RNTeDp1L18U9szz5pj2ay+bQPsEYjnapeh4BL4jHjADKR0J3TnZz3dxJlpwqdNU
y8WQvUQOOfWCnN2P/m+09io8PMGFbIb1n8TNchRTQPhQsxfb0vVGsekl1rLUJ5iI
rN4VFDZPdPQkF0jusqTurtZwQu5tk7qJxZCGBP/D2lL588ZL2i/9siNcPylLdZUo
TKwzQIKEdjl7gslB+TdR4iCgDLliPq2IEvbPjBJwUtYuDjYbSB+4Uv006sAnLua2
bqFmjwOEJZpxpSeklBfsdV4gNyeHYXZ66NzV5rUmNgGfixyrGC0to0sRHIcmJRPp
8mcr8oP2H4uk2PoFwVrJfL+KeqEhYtaM6uvfBdjPtZ1CCk5cRbZe1z9lWbhEqzZ/
uvF90LgoBW/xoynrQHlzGz7iCSWjoCFL7XYynRMV54nx6+WkYo+Wi96Vk9GV3msj
FbZ/XwxuokC+U0p56hkwr9uYzoAsOqSPhsPqi7npn0sJh/iCq3IUyNFPeU3Qa5+s
rBLZQut88h4VREowq7TucF2Ikiz8NIAbLMvOtGdXq3I/9ifqnqzL5fGudw0nKmUP
okzwCZeSYcevZW4GlnbZ7P1NNqVzxeVvetKsgrrK/7YBIeUovWuzpk9qX6XRjsIo
OYzH2MjD7Bo3RVedgI9TFLLBwESYe0mueIbyoXZYHiYAqEiIjjYSA/rp5LLvsILI
LkdqPxJ8Ug/CkMWLhsI8DO8qkV+8i7lsm6RvQ9bhIHMR8XatTVSJ3XgnffnAGiFx
FaUsuxDmhbYq+mW5yaavMFyFQhL/VrYamjAFHv3hvlVSSeG7zHluKJ+W2dkcz6L5
JPOAGIABTMSEwXol3tptqkJ4VKLgEDFpvrqHUez/t7aEoj52szTRRsAIhVUjkPJ0
QuOKvKsGlc36nZNwtsTqdhmcxXhLyVbrdw+u6kJZxRcT69JUGDJZMaGU7K2VzFwq
JcH28mjf5QBNV2HUwUKAvbWOX/jtKQd8khG0JBDbouKolRgxjoplXIlcjHgHTGYy
gHsBFhhvy8OHu4kfUyxmrXVfs8rrrox4AbN7sRl26WbEjCUFy/kcnu2OgDFrBBRP
WMZGV1m2z/K/5M7ZV7NDlwzjmfWPN2bJrSbDt3RfyIftmEQEy0ZY2nh6LnZq0cqU
r0sa+sVJz0vPcCxJ2/DONbZVuTOKdWrWoidZLosFktz3/0gkPrP+PxLjpm9sBtCt
UFfbdDaMuOSJxAqzJAptonxJpxave8FETnkqMbeJrflri7kuV2VC30VeQJRsLT5T
Ch5uaO4w/2wJC6VWT0aaMLKqImlFnq9/Fk/ciTb57O7H4+uhFct9Tnnftc2vaT/L
1KaRciBQBkqQBStl1/+Z3tRaEV+vE21HxIRQKXOrwDY6lyLuAomUnCn9/F7JlInY
DIqwvzngkYl7tJ2PujRW2F+8v4Iih5vxoEMMtZUkttCNTVUBRQSaNi3DhW8z6yeT
jaYxjqkxfB/ZFCDChLOYm4Co1UK8vRisasOvsIYGSIdXL6GRJJYQn1IwFjxzKjB1
4L1Kql/AxhyQkOgasyUHzsKCmiKd1XBabsMlBVy90abG1alGoEr7mA1/xTY9hjfY
IS1m0dvuAVnU0ZgX+AF2B8l6Lf9lREnsGvR4Cv+IT5hdve5DfQ27oJIbgfEcr4Oq
jpxble6VcZq0IijPN6djpl2MC2uc0LXDV8sQx06X7t59SoLZMQo2j1tAlEyohvWm
y08+OcRJzytemmph1DpQj+V23uyKji9i1yq1jgUamoY+p1xSL8C66nVXK6YUDYUC
aNHb7zxFBx2jGBqwiRpwKnIzVivZB3afmMxpOa6vw3eOY7ydEq4FdRBczSnA4iVR
lK+jAh9rH6NKh5bdY4A4JCfHRhRDz4D8CaImC5O0NRInkipwENB53RocR+cWk+nr
CI2hSpwmwNxuqo12MsHdAbg7YJScboffGwGdX63umTKv2nPtZ9bvt5plw1rqdBIx
dEnEVi1DjR78TMBewuxGLWDf/wCIGS3kB91x/fyzpojpJtAWHZcxBW/42fB+iFmH
ILusF6PXPsmTOhlcG7dlN/76O32R6DFa8AGHG/rsqZcoPwFvR/0tbWDMejjGDWBw
XBO+jPVL+Z8/ZCskC1i41Q5DAdDwLh172vmsUmGjXC3SOyR0v+I47g4NKlUYaubh
ABwZmlwvIcBK7/J3BKW9GeYZ7C1qCfUTps2MfTUZLJaX4FVT7Y00XeI6G7d5TLcb
nf8YqxAeYVcUDnPXYXeEAxKd0vMmExjaQHyzlsH6KXqQeLa9OElvwwWgo2j4/mYX
7ID6kCxrdloqORfotaKOrgjtnaSe/9zEMaHFvUMvY2eGOdhb1JINBhJtLzZUTc5g
/AANxmNt3aqCLyh+eIPyzWm+Kkmd38jSAkFz/akZXyry18KzsSh1oLakEkfJt0s4
X+tC/fKbwCWVfVsAJg9ZVfncKdZS6JjZocjk5k+rC8eCcW1aaKBU5CmvPNKNm6Y/
qRzbyFWIIvEeMPkkjZALFSDonb1bIZ9cDbge4guq15o1kaPCiSOaUYF8z733vh4F
GkYYV0L9YSJZekyi3EgIzypApmodcWAaZbOLcTtgrc4UZ0naAxVUlKAcS7IIt+Yc
eZmjG5TJdY/5c6IQef5m5UQfHfAv0nXZ3TxaOxJzeRAGtrElLlz5V6JJVHffBTdh
Vc/KT3L1UlAlnPE1Uk/dSMpkZgUJzhKNVAQCTsUQ4267B9J/2L68sUD8WCypJQ5O
aJAYPGItOWfc7Xw7Q2duTRVxTox+7kAjfAPSNXF56A3gqeIdAKmwADSykRa8c04G
WBEbwmd5C2EYRIOkD4mDrH0/ANghaY+aki9RpikVZC7perPwNCAqFSvg4bpuMB1B
Qr162As+gsZ1Ubp+lrkC8HuFBFKUzlbVBBH9pYHNghQCEkFsq3Z3VN0Y6pf0zHRi
SO6gUZ4BRA8QjzLBL7JB1l8A53iyY57IoNdLkYSgaKNHUCf1NvMPvQs56ap+GdQY
bsVLvXFd8r0o/vTXD42wWkYJR1pFvJFS29Oyim29/JmMbxSrnGwrAgujPFFIqzbN
bRmkw8Q8vv0+igxIOBaR32TEXTM5vSvVRznnGgR3kQp46I1UXL9lXC7ULGHu6DaG
7M0uL4Iorqlh3OjfXrVHTfhR4OYV4qOmc5qzWGJZ1Pcj3AmeVxL1pmlRksXqtw/G
kyyKaKytjtwNnjuMNjZfffo3iKKcVRc4UTJa4JdY9F5P0pCA4wo7B9SH9IeQkePu
dj8pzLctLfu4DLeo33ocSMFb6vH2rAvn0xtIjFloFuBIgDAU1YUsACncndO4JkQh
LJhDwlv8EuXmx0I3iG+kRx0/An8IKwdDoK07hcSsKWXXRtJEKk92KRo8+SvyGssr
xvCsA888OaEc+++LOrP30gf05t2RlH+8ENp8iv+XlZWOt2a2X0hLuCLPJpf8Whmm
wmnvUZ72rnTXdcKx7KWjRMRV1t6Y6yHuBqMiMS25WLsHVOFUWaLpxkV/eMxj72pQ
jUnmTbr9zqVoa4r2vkP/K9kYNA3lyxCpapTeBAXcRLMq0tj+PnoH6ILtP+DotM9/
nb2W6Xocl1rsgJDn0BtdQTwIiMD3eC2P0YjJQqaQ9xO0r5fscSWevS+Co1uuh6Eg
lFWHkk2SEGBrpvXf02HBONZJfWcBwEL/JQY2YfFeY/ScL5wQzD1ORRYMNwvkAAmw
HI1ufIrAJ6cU5jOzK3+D6Kfn7ATZKHYDNlSNoQamp+ApNFf9ztp7pThUZ0GKeFas
szUhNlvLguNPe5/3WTped+I6QoAg3zkh4TmsEhI2w+qGZF1/p96xxsbPdsUnWM7c
xxDa6Ax4XOSD+cDzO9waDlf54RqJvIm/v7f+0uFmrmXzcE9yVzWWYw6/WWefbbPE
F2KQSA/qcVADA7mcHXM/g9YdeWhblUGWb6Ku+UrDT+vM0wgEJNFJYcNaax2XA85O
q95Jz2gMmaIlqHTRDbMcN7RGLEpybYFvZQRY+8KhQh7FiIXrZKRJ4DDHRknX1Ltf
TaCBmt9OkEoDWYnGwDdkKXsYIcHAOIOF690UBz7I39b8raUP6dEFce6+/DFDlW2Z
Z0hUmaUeJKP9L0AvGo1NxynnYhseIPyLrwFQfmbzafIKOdN8L70t/7/8pQeznjjj
RsWAddNwN0amfAgTwRXw2x7stnwOtIxJqB4NlnH5JdSSbfpwDIqz9CVhspjMxb0h
a9WyrEnQgjkmNM8aTArUpwczMfGaX/dfT6oT0/PsD0Ub1HT1QBjRE4dpTYVtP2J+
YXElyxkpjDe99CKA5Q7tB40oFOmaZKOsbBSvzMAnhWuFOv15AO6IhayUBH2eVGWe
g0hklS8mmpiIZ+vGGceHu+SFzmUh+xvmIBUUqKWiZnCKn7BB0UuYBuA17X0FV/eC
YN5wbd7FxQxYpGyHI+dTmhOq+31hupDMOKlQFJn3/kmZiFUHSM7f9o6lMm1d1Fa1
16p6W+B2jSk25YLZwh30ny0KSAfLg/4yaeHa3fgkw7PnLUA5bFsvuWv95WoClr1w
16z/LckBCKcGTY4674u69ZNZQqK2+oQwojwV4LlhyFTZNMSyAvoCFuKatp8LwDfv
IhK7/rIy0FLImMwKwJnm0TV7EvsNjMiRjUf8+14I6LOcQg3ga9h9DYtSAhi1B3xk
j23Us7OihAZ2YZ1VNg+voWb6m7QIlK8ULIvqbAMKs7Ytsln960QILFQMhS7Nme8O
Vgyri54PNAJFQOzQhuzfma052XPuVGXja9pagtKi5SEpVTC6ikoS4oT+PYFeziUs
cgNI4Ye+W29/jXXEGbZBmUjYWX7yqmPWQ51Tw4BOQTjXPjHL2/W5K60CmbzTAv9w
aUDvlFD0u3IEIzUhra0zCMACJPXj3ALyMWsP1TBuHeL0gsRhd97oIMcSw0Q8DcxN
HGfHMhAtWm71Sq9IZJuN1kXUEKG6seuw1o+2p9le0DFznFD/tqhvWsJ0gl0Ejj7+
5I7bNLWvUDATlAYpwg5o4U2WJ2xk2l8RgFx6JhNEE6/eqKvtuqRgzm/Ybi3YeGEr
Utkpv9bJ6pbIrMAs1pDbU8TKNWe3buzEFGmzK1uqN0jYpGVkv3RZ4Zg0SjQIRZem
7i+qZg105TVInyqLMda6uEwhvtlHmoeUKMykAcbuiGntzf9g2xQwwt/pYxTk166x
lT/xXEGEioMp4Hg6oiz7SWA+/yIkNHWQZSX+ogPvEv8FYSO6v6ezd1P9g1sXtmNi
TOKfGPn1soXIhMKaBe2lL9anMxFvWKotuxrsX7oeSGClYia4rlh60/MJVFCiKA/I
O2kA6FtPrOQT85WeeUvTCz25YAWA0pFDalkT6ZGypfeZsRFyyQeJTUYPACTdRwLI
Rfg592xUdm1CZbliRWpgVOJtcPPMEaWvDDPArV75ajSpZ9ztOMZ08twxpidULZBG
0G59ajIkyazx2tqRFaVQE7ifYH+Sj/0O+2SIShzNUWorHLeeiB5kc1oXOMRxDaVP
lkEswgDnYTvAGqmuqljn7KgjmrgWZC3qF38qoMcQi5XO2ILz9WInEyDRLUq/ErRD
VqbXvNcCSzslpxIMq/A/oHvaCL48FqByWjuFVrP9EiXpEOZODD49unj1xV3ZDHXA
pcnrdj7rbuZin+D7K3Adq4tYdOg8FXF6KJxhE/pgg42Sk01kKJnADAMJGsnyQa88
Jp7mWUZgVucJ/6wzjGeNspE14QGIEKcyZPZv68Bn2txuqmFOpUeF2Ksim+opr5A9
UsaxfPXlCQZ3zPEByEfbkHc6baPiWI2yjODQM6pQA3cWLCmVwpo/n5gfWRELR7Qw
rDycd1zW4i66ribs8JpwEnWvcVVMbBJbMH0pTvPTIFWJExBu0TI509sq9F+HymNX
km+ZVoF5Xpgo5d10xmAbGkh1CusOR9DPrbS6ZO4GgD9q0KuXUfppVk8wncXNnpzA
LuHQIuGDwYbRJAEbv/qSKrN4H4z0SS+TuUFKXp5w2nm48T5YH6gmX1m0jJXf8/3h
EwCdtPy2VJLVuP6/4bg8WiPCVh7gGQXpbW/YRcUfr60pFlQnbwUDgunl+q5WQscc
oiszlbFadOzxn7v/jVaPMROeYGUn8cTD6/9Lo1xspVtltsBoVkBgshUk4eGF+n2w
7yIuDvGY/rK7xcsb+4k5qs6uv8I4RqnWN19YaV6ksQpvGYGzDJ27AWEn6hK05q0E
Xp8gNlk8o0cfwdFpZVOtN80VCsxxjVqcs9XTKVPe1wE47So+nJ7vHbYBrqo2fHoy
UohPfpoMmiVU0SWh302v6up9NUts9Mqn3iEv5OVEJzy5m24oBtRH5d8NDCLxf+wx
fbMvR4fW4vZVSHd06yiur/HIcWH+luEEydP+VSmiYgFz8j12bfBCja/JrqPp2vYa
xmYHgAZQeegtU0x72c9+O5wANWyd7Rpe2wyapiwPmOrjkWRs9yIdiUUA8MGXyPHz
sLdhETWlEJ4eM5HtTtwr8oq9E6UvQnV5b0IapgS35KA4MOfz3Q/AyDLpczRXsbZF
TUK7iytUuou5zuV8r6NKV3y58PiGsaZt+e7gyu5TH8ff/Btr6TlCuzRbNd3VIy9k
47pZtQ+cCHqc+bifdGwvB3NUXmXxkxS+AtAIZR7gK0fViBc7NzeUJFOsHUVUsmZ/
SvFSWyrzN8IE5L7pKxilhU54+bUA+3BgH0Vxklbj7BzD0+2M5eb7tnwvAJiuv6FH
WLdw1fB4FQkO5czMQNA101hCAIbjX7uLdE7YoMdjzstNYQevpnfhTDlBFiqEzL2z
Kw84KWcAR/nx6x0uinZ00EfSiOSBF541szSzHD5y+qbaO2jJ9nBxtOVbNLvA6wgB
FG9G85RicDGib9Y06vTolWvTOj4iPycZeFSvly26wR5ahn5+PMmEZ/5/00WALuUP
55xYIgBMXhW+UcWvG/DxRfGJr22tJduaGSGmhuJCXzqvPW2MxDXZW/s94FDhF9I5
DprkwO+KM/8MCwnrmCHmPjn0uuImvIfyra4CV/4CfOnkyTBVJdroDEGjTP174gLO
Umow88I3F5qdBvKpFWJfa4ZkzghWrOVVWlsX8VED4wI+UZq1asQi8LoTfyNC5EX8
hLGZvCicl06fWhu2GTG6nwfrXwfVxnKNph53aN33DDg06F3nE3ptz1/3+QuEB2Oj
0mMD4ZNhm7Xrt0cBvl24RumuXnJkD6iQFt7CX1di6ojSn4jXFz7j4McN0P2E6fo0
lRtCFhzH4kC8ObO1q5+A3rPKDuKX0i9BVANzSva21i210wbYW6zn3+U4LRYiohia
HsCnwv1fl5dtJteHJSdpPJjXbpMsdqm492PLskKfBR4ztfX2tMdjMjLsGeXLQLih
kXrvjP4Gsaqaqgnc7hD9c5GoOscAAhvrl4+xXmx8FZJ3Re36XJWy4w/3YFr54RkX
ujSvwmVFAZV9vVwlI4Fz7KjQHoWsGvDy5SQeAKwORy98GQl7gkwihr9DQPUbNZQr
gR+cCWI9R35WWH9zNbHCMGPo27+XKVQc7GHvsKbqwv4Rk56oEvNcrjna8tBirDFt
Mqex40x1eoteu9Okna+DXrRaDlUw9bLOuTT2KcyQt3JnbRWQI9b3d65P28lNcVoD
8+r5XgzeiyuvGySeQr7RyRYXLCQpWEF90ylED3+c/rJhEVrFgCeb/mmcmTSEjU0H
F62TzdUlX3/er+XQOrRgOOydBZHc6pnpWZtC/mPZGiyRMqLwrp+DwVxU78z0wkRy
vL2LdiEF7oSWY0O4FPgu3CF4aBZc1C5h07xKa4cO+O9URwHBO+nxTgvT4BHwsRbp
9Zf3BMEoTf/d5xamzAMk4YjgKtazsUrnrCBKDK88w4oqgJUAZcr/v/wex0WXZ1VY
QCRjfxQn1Q/kwpuDxaqUe5p/Nwp/gKuJFVW3TiPv2UoHsIkFhl3SGXQY9nVDVxrj
EVTeLkgwxQQQMlMJbyCfRebw+eIyZ/M76q7M9meo8aqWefHv9AhaBHkdLzeDcgXZ
8OhTItl1NpeLtFp8ZLAzgwKYHR72L6q3e+laHuxLrTI343w2cVds3d7TOtPIHfa0
TH15Ey4OyICSl25boCk7wgOENqSQmB5Tyywx/ZmLomnvcHDhS4KezngwkH3IsMaU
0q252AAl0ijqp/TaR8owyhL5rQK5Mvss/+fu79p3Ks+Cg4La+x2/tea99IgqgKd6
cwfDM0zub4VhzbrCUOQl1sHNRJ8B3EapEgFOTQNAqW4fmDn0EvhBdNUfbVBfaeJS
ynBApM+y3cPOiVEfgMyN4JaewQbsLyYaNceP2qYOD4fq9aE5Q1jOM7UAlyW2uf7X
43yB6pqj9lhx+/9Ja43ue4hmdqlIJjqIYH8jj2fEagcu6a8iEiqxrAP+1pwoJVF9
tD9BINLjhKs3lCD4ri/q/ejplim4Jw8A3aTQAHuUdlFudQznWnMsC8c+CRvC+XDq
W41Vyl9lw52vTEgH5iboZUZUp6QAgvLhhWrRzWHLPz3aftuUY0UCCqe6beTuGFHm
xCWBXb2dYQD/ozGFm/h2nZoj8zEeXisb1Aoxlg4aDgm8qVSPas3ZPXGmzkBQbzx3
n/hu2xedjfDDVG5u6K0h5CWckUMXdj+hqLrJB3w7Tzl13llg7F7rJFE3RVWzziJZ
9RBvX+nCRrULrLkwk/JwBr4K+GnXf90FxvBEgSjP1jWc8QrZMcx6ZkM+yxyFlZHo
x6tmnompdYLLVQQvle/BoGyJ9aCZG3FIHzUVNuEvx/6GwguuHyW6M1GW/9o1CQ4w
v5v3ORtrgJzIT2FtGnaU7DEndBYIi1Hf/GgathJZuUbBtIxEsEyc+h9+5SCQIJ4O
B8RqRvauWMDtccdiH4FTZWm8EpsAJaLuz/AQ15HTw14khyv1p29PiPXzxpJ60lNs
EW4dIyzcKgoYaWhPsfD1AbrF1j1jPZzVZOMu5J5Cdl6Z6b9Q00qkiMzN5652W5T6
dyIOzw03nOf1Q3Cd10XBYBheidAWYPcc+aoQUTN06UlbheOjRn7Sf7lIvNAvF3qN
pAWgBh8IHV0zfl9cq2WVPwrGkHEpzHr7wdnMV84Da9LPv5LTL+FUS4rJCXVvm6lj
1/+A2ZVFvpD6tRssTgXXX7SIqlv5wFaZU95/PK3oOSK3crRHNf6bNYYMN9OJZddz
6NA7dRCocvgqtF/fJzckIziwF/PIaeR3CGMkJxsPvgoLOQlmYS7nwc1Ek+PhnV4h
feyEY2P52DyGRfTTK1LOwyQ+biAHup16sPmwsagosXpr24TifKuyXq23bSdNIS56
JGhlESRXhlnKHj8S/I5FvUvwb+XI+1SuzVpJ3q0RbWuhTxYiQzGCBBQHsia43lfM
krLViWvrzTbcC9puyeVqy1aG5uCK+fWLjJTFF7ndESd4ocU7RkQsBM45eRS5DAMJ
UWmnrKR5pS2T23ETpVa2FkFiSPNTy44O0K5NN0YKqoPswZFtn8NGDpOVadtjZ9dY
uviHwGW/4TwFE/JcE+e73eHIMoCE3Nei3QM0w986xEDYWv+XUWfxVf0P5L5rNnRB
s9tML7BMmMcfW4v+jBWQRDOvPQM6XIjOkhm0kPWpyMUxJQVxgqUDZLlu7HwNdkr4
f3M03CMtiYInJavViQSv8hCwAwJe+fI68uccWV+QXMGrrJr+3EnlwlUspg2A7rsK
Ncexc+O7ZJiBh2DLVi74H3wD1RS60GTkKWZ7e+Ve3cfjuX7RTXHKdSwSHDaeob94
4hSZeyjpHj8rkm6uFE2zFi1rXr9WEP22ZE1qREylVAi0ael04jsW6T6W1ocobwcX
NFM5LcNJNySyJDkM6NLRuRkq8xwfw6ZzGy9koXo+sZBn2YZYAR/tAI2HNhFJ5YC+
j0wHqP6aGimco+Q4sh4A0Xb00bDoyx2o5ix/1Vl+y99z6BvX/ZZBbpaaurf/aPGR
EQQi77dV8chwT6sQTnoS0/UxNJlvExOwBfTUkFaXKg46f88PI5PDo9grt4MWWh2H
JEX+OscSNX0S6dCoBwnqz6tGfCbd4d2ENNpeyBlLBmWhJyxpb5YT4q+fSfh9UZdk
JBjS1ucNYDo5Ug10sx29KS84aq8p7KtATuIQM8+thXnbeycKsEc2eLkdKNDWvgju
9+xyJE4qhKrXmokBpUyNxvc7L6j/d9BKL32DVQ0piZoIB6hf4UTOcXtK8rxc8RCz
melb21tjrprGQR5D5PROh9HgB4jVNQnolSOJz4twhgjUbHodywebqhbmXTK7Sivp
li3KGZTi9h+f4o+5WpZCqmFhHey7FAiFrFpES6FOOMTC2YCZFlGb0Rnh8gU51X39
+K6RAT7v37Fq+O2oWfYwopgIfJ2OkO2lCpk1JJjIvscKoh6Xlge9xJoKyUfZjIq6
xuJR2YjesvQwcX6I3DFlscWlq4yg486glYr5Dz2cD7vfQmvw7tRJyVGj+6DqqJPj
SXArW2Ugswzu+SQfAHvAFI07NQabqE/BZmhH4mmiWZxhO6gOILEKMn0UmgeysKoR
BGj17NM0MmmuFLTADflskK5aYVVTyp6kkjZXHO9/pbf6TphR3YhPXGOSEww6Y37e
B54bpJce6kW258paVTMmbbF9mDX3Zd1d6ZhGn2HQihJYCaop9TuDNUa4n20HtaCI
8H8wfQ0l0VUQFdx05JpSAMt8aan3XXHKhv/6WQjAksuWWo+qqpl25juIYd3UIpDg
3kFRXF+xPLUV/nG5DC9EKdLghmECTWm5gXuwTW/xV/weK2l3AlttlU1/pVj/yJwN
b2v6Dgp2siO00wtEh4lfVkoydbRH1JskvWwYV9Ajlz3lHM+Nxc+u02EfZYPKM7Wy
OOtNNMV1jzXvc2fUNLq6GBCCDQrDE5rBz61BGlwVEJnpKmPmqN0IgZo6c3+TW33/
Vp7KzS5/OlN6vC8HcGluLZjdjMC9EBaU+yEm04x+s0iyw8cFSPNOXECtplqtNkPi
MFGwOldnSYd/f7l/cqZFuSYmv7yZAhjzaJ/HqWPWWathDaKAQDpmAFBO/bCvs9gF
XIYjekxdGQhGutAdvmCAmVyQBTct5doQL7iNjnQeq1pFkGfVJr+VV+hfsa2W0lvH
pPhQkhqQ1jR6KGkpSMoWNVsCQfSQzKC99hM+PBkmGBC/vkFpoZua49go1Q4z1cxY
8SNLy0UCK6Rft0X/c5KLf523zf/54o8wWAPLUAmJ0YZgUh1s+6RxFeSoMMSP9CYQ
P56VUnkO61r+DY7AY6u1Dbvm0Zq4mseC2mH9ts6EKliaNLvFHTPlWF/wPwUKF4v2
midK+JOqxmDbLhqaXwIinzkoSAwtUZ3ziFeEL8c5lizlYNw8vJ6HsEBAigxMOMvP
uvtobTgoqhgDZ4M8KU+cyNsYGs2DXk5TCpkhd4QSHbTMkELTxjYnHLTsx1+bPdEy
j69tknwRbT5bdw/giUlMFBCrOexAHeyb62ddM1Vn8Zfqm32V8e947thnx0mp64du
eWQNhzuYFGNGS4hWFy8ApMt3kh34gdKOJysUyFxXfcRUw/wqmZVqn1Hd0hPdxTJ6
eoGkAOBkRW1t1wla3kJZ+/YB9TIbDwwyCbt8J11WTun8J1zFQHY0IKMB30Lvawu5
uobO5GDja3WdwZHUDez10H6xhh5POPWpcPMkVbbcmwO2Ss+ADRwXGHnJgsLVQv7b
mMcV9ct/oeXjtIbsW0WdKwF8AKueYCr6hVP+HTZikc47+AQiHlwzBnYWKM5QJD3t
wuVX2N6TFMLb90YPz5lSK5xK9LV8VdBuRopg3DTBHZ3u1hoUV+AxHEutKjtoeyND
uUoqZU2Pp42079so6yW+icBMeERbiytOhzZl9eZl2YyYV/iW5bKdTUOHo/mNMEqV
Neg87giKIzQYcebBnzg3jqIz24/EObPbG5oXg05gymNqKfkWnGHgmg6hR6NS0arz
WjYyH0IPbIDjmV/3DskS4V5ISxr5hIggmuviqM1IWf8oZn1u9v2u+aT/DfTd61QN
T3EPPCwbSnOSb/C0IDg2TmPpGOQ3+x+e4YNa4WGgDAWV59WEsj3RRNJzMaezsOKc
Vsy9MFQReEfQn1jfU/NruHPh11mxUTPKLXpGLSRcff1KdB/qgQO5BxlhvNTCZ8J2
cZ1wzJRrLCPe7EqLRi0eSCOxG5bGEsIcR9d8Kpi+Maxej07rkTVaRcomIIK6xdIV
I1EWUGCUgU99DvfoMzHUfIuRYdijt8CceHelk48X6tC246Zrnv5B4+itBQxog3Kx
EP1gtHalYYn2i0J6Vm0itb8Qz1zAvf3PHipYIcA4K5P+CJFcrZuiI+Dx8tyX7ZlD
edguYBs1w2c+Dd0ArLs13Ali0046utgwSm15q0Rcc53+T2eJN8PWX4Kw32wf4Fal
Oo7QUWwW1XzqPuTsxI+S3XY25eMi5/1pUruDIEo8LipcrRHfgW21k7uI331nj5Cu
TC7lKtGOHHiDsQQGerAdPBRESOsiwJu5A+9SAnv9GibDC4siljGy+9I8/ImXgIwc
gM7KZBh63hn3dPpSfYfj3JdKemGIt1L30F2dBVRI/Chma0kDqRaNiiONw85Oyox+
eQxupge0CquQL0IeQoI1KV5uShnAm3dVXSKjkRIv2H7IyP/gErmssuz0/cc8nfAB
GS4C+qM7RjfPVdRA1PM3oXqiscISb4Bc55BTXLC2ovB8MJB0OmRxz4BDvkM7WSMR
J+SzPXTxJdEfIFFKVto6I4jjTuNpeobTDV+GXOGaEWqwauHtPYuL2K/qTBUP1Eog
uVLVDY6ZebSLX2QwKYVEge7RtipPQCu5cgW1MtJ9UbzekNeFbIiEhfv9ovIYle21
YveaM0xgdFwyoF8GwVSztzv0biX4MTBda81xF+AgvqptlXjW5T9zKjV4VFRUuQ24
bRPPktx5/In5DOa2gUfW+GzcVPnIQ46wE863NFT2v/TpjivOGx8zY8vBOXel1CFu
QZ3W91+M1SyZVXQkAc9TxTYMgwD0CR7QXFtZogsbehQgHOz9dRaUrtcJNw2nct1B
kPh9MShhbGEo2gdK/3S/WKGXe5uK0EY+YfCyJqmd7QXExRvLpvK679+PHFeaTrka
0llrfSZrnpx019hwNQEn+cnvkpV97SEIk83ZHpmytm2tteQx5x3oSdFtypBSVZBm
HDtqT0FsFPa40IAZ0J+kX+qH6zHuBCjFROKwsCcgxcwV7X5GTA3YJV/LWO3sMXXx
u1TKi8bySSc8PjHceAzY0HXPGy0qflvdy9Vetnow4LC4g8DKPqwqwx6XeEWgzg33
MV5M7SAHowl2Rwko2G9RLctmeS2IfAkUYUNyPcoT4a8n5gVxJrLb28oczIEZ3GTj
nhio4yaNOqGfmMPn3eEI5o2cbqGM+6Bzb1mGKljYi30S2Y/RgBu46Hf86HuKoJui
NUmPskpUHM7kB8yGD5gFF1y8CNYNEANO96E77mH4aS3vSc4fdwyrLcZhoDKpn7RR
QwdBUHNUMaFddXKfWo2ABexan1qN+mDgjSLGljp9J5tj8vrG/Q97UkMlIlHp+nyn
j+gz7CAsJjeCJG9wULCUFgKF/6/KTKKHGrOwnwMwLKb3Oyc8ud971eJpRgzBIpzT
LNkSy8t/gBpG2km6INEKH35eRpd7W6Dx2P/mwgS6Alt9ee2F+0sNsMEiun7FgxbA
KXD0ljzAoQT1aeMrCWBBgiR4zmMnjVCW72sdGy9exvP9xUPjWWpwGRmpE72g5FwB
H5wKTxzBubRDlgWHdG1HTGJlMyOyF1bRjLlDO9gVe4e8U3KM/q3hDW7/lDdA3wUk
bR0tzcvSe5vXEbAV2PJPn6Ja4z25taBD6OAm+N/nqR1i3Tmx3f7LfnQabbb4U+HW
oiSjTsqoXMLmCkEUXL/x6o8xIOG1BrYODO3rC0CBBWHv+vxX9dfpQfDS5N1PSb1o
BZSHmUrp2LUThBR8ePRwcmc9AWkRojz6/H2XCSvKTmn5KyqTdYfRsovBAPFgM6Dm
u2qBrhFdZdXJw+5tmlm+aLN68pxVbCN0B6ercx6QIz3Aby7d5ijRJnb8zZ01q7Hp
6IHNJSwp9bs8ugB6pZjJbJDyIotpcJr4WZ2w4rXNWndMXgQzfwoU1aO4avPItM1F
VdDJfvGof64f2pb+4C361WoizTkK/1YmvugyxRP+B20ofWuLpDasCtlDGQkKtPFb
PBtyh05NrZ1fAVR9EqnjsASJUzj+1XSxy2KoIh1DgdjLRCvhyafdf5PmVlIQ3dYX
1TT40lbJ7Hbpsi1psj8Gd0ufuXPHhOtbzaWvs1XAh6IAGHIE3HN58CMgq+ncNouq
2SZFYcXAXvLueAj96gvHr7dsfIFpqVJf8DNtBVIC1GEIuloRGEG3oFYL9vF2bzbX
ZA/rhHGpvp7R2YTYS0y/745CWzOJyTpIQz9jtv50ROGgP5vlHIGrzyJJQGOVYzTy
kJlor3koE4H5VK8jhsS0jgMqShh3ffIhiBBraZvVWSnVBKiGy56T1OOFBGckaogE
YioPYCRo6iOcaJmzRO8w7/fCm644kLnlSKtsheMrHtsxie5kQt9m5vMckI10HkPA
l/kfTnNgIEqodE9IjFI9QvLd3KYnKaP2pXc8pIq/81WISWotSV46IBX/ViWizIKI
ljZscaQgce0n33GkeZFy5hq4l/yrJ0OOqOEPuvZVo/C1Vf9q/eaGIRshrJzhlSV7
cv5MJ1UoN1nAOiiEyx6HA+/e3pys4K4oj6OzDayjegO37cOjnNfR7QN06625G8wH
pfg/wUKnb1k7RdOitQjgPHkbwkHfQfC8PmfX/UcWlk1v22AVqcZJH5NDYxfU2Yk0
lSZCrr64qefb/0oeplnrxkGlr2+RCR5tEpJP/F8gx2FWl3kWOkvUoyZMx+IzDiHC
hR0kNN4sZaI7GiEKMV/Iok/B4JAjlesvFM56WLEYDewFYFR2v2FOg0ZTYRz14mDC
XI2HKOtLMEZY/GUW6rAlXz+70PYYyiy69aZ+efpbfUjT9ANMezjYJMSkncRS9Z2Y
lQSn+bdvHNCveTZvuabxdBRuxEX1v5syVHTQlAALRauKzY1VoGHrDsGSPH1n8nbP
jpwV0xCsrt8XxuT36uf/SnR/COw45k2snvcbwrFHnKUAZd70KNpaaynBBW+VOjkR
NItzwTVBF1wXfsO7euQVWMhBqKrECAm1NtnaB7nhqcVItUFoEFv/fV8CLR8/5zwt
iJrazbZxq/sLyBJjDv6riYJJQDWoTeXgTeNdVf9/Tf1nmjWFhGK+wnzOvUXpwEwl
ZwrwVn6aPfATHZ9FdnBm3hw7qUx2ikQms/eEQQEoGE2NH2U3akcAXKy+H8ZRlIz2
xoQ+3yZcxnTXZxMGrqIY8o64pxexzFyRajfqxetoU1oRWRg833CSHD7ggsTDgNCc
Q16xRQqJJecnjkAnL87So3I+Yk3GHhofrAY2nYmO9oHtVArx4NAVRcTwvULH28XN
/GQjlXvpIRUHuNNVuymmLCgvSQ+x6av2rPTopLEJROWWOF7hK8Tl9JRP5fyv6mlo
2vVWyjjx1lzST6nXIoOgW4On53V1+fZm7b6FrEcmWlhVdJ36PWVDFwom9xuLWHu4
YxqPCQWOP8U5tQR9oX2EI83MUQH94CbirpPTXL56fxxroPSxcevGr4gKjGMw8T1H
OZhvKG7etE1GkgFbIFTR3gD9oClQVoxgJ3CMlqQqSccd4PZxJZhmf0bpKqsSfOT7
URZV0CfzuvR40idbq8NKLuispHuHLsNh7lMiUBTwhAF7JR+BfyN39dMYEcLFq78C
rrvWgbG485YXcM6P3f2BkmBu2n5aqOZN4Onf5SzzqBaZogsMtQaGIar5ZyblrrQe
2qf3ViL0Ikv+2O0uCeYZJN6LLAY3j5LfAAT7trx/KDuFaV+EZuFxuhNAEDNlKTvo
j+7OpS5L9sS4jiNmAfLn0RMbKphIEmtZakdDCh+iuxbSatGW9i1ylUdmC8mILvyV
4dRIS9St3WHnC1zqjsuMOTr+Ny3DDjlWQuUzUuIGubbVXOnDzTnFbp4x+yuvpHub
We2YGdmTg+Ebw/K3DTv+htj7fhus/+fg9qLgwTtSwt4Ao5goGYL+NIiDREo3KCYV
AK6Yaz0WDm6BDUQPCRmWd/hxydD+jQqICyfRv7AvdjqmwMjbAAf0OgigYVV2tnU7
IVezNTQsxUKkBkH7v1iBN+rB5xCg81gp0AK5UV+vN/u6bDArGJ5/vGvG9Pa+UQrL
s0VfGqRxGxSny6rlGRoAbEnDZR7MxI4mnYN6PgGYvO9JCvlC95NAC3pA5OnjqSfZ
0Snp935EvtYfKFY9Z+kHDzIgeV1PgsqPbhfWkwJeeKJaV2ODvKOBUs6x6govMvmb
LmMjYyqUhGvRztlV3bSEvc/9Z96G5lreoqC3PGfEv47w2OlylYjfkukFiLnKN+3E
vmv9g4/EtaCXaRrQj4WJWKJzkY3uFNqSiXjSOMepiFfWyArVy51Ng2igdcrVtwsq
B9vNUdV3+WKmYP7LV3WfvcTWH/LRDLIdcAFXsWvJrsSRJ4NGrD+Sl2vvnMiM4h+Y
37ULyUX7D8BosSdzPmI9uerKPhxmUFI7biBg//xHE2ZNGvjuRZUD7BthJeLh0JzG
83+stebatbsGEOTzU2tehM/TR8Eod5A4JPb+5O5Fk8vYuM1ejgwG/6rhXsGoWNre
LBFpQDAu6QfQjYp1j+jr3QDT25TCEqfJD0cn2UxPO9bcrLQZf7wAy9nI7VJOOWhc
X4TKvhvB/ekFK6sPyBEy3qYRmK/K7lWFj4Zy+IGNGq0F/Mh7FjNjywVPHm0CWLOC
9xDwVEcM7P/g+EGLlYz+AYXPTxLlsO36/SqIxB3TDXDUK3IKrGKaqrARPZA7fDX7
0AitxIII2XO00EEyZVt1PSNAWfcEyrt2ZwmAClhqAPGjiCh9dl3twBTGPOC5jN5z
enQuDqr/ZIug4PnpKlVBk9KBrLylrQ/kbEtYUA0pIxEolyqOFHeJkmEtYj7Riynt
vLfFmaTNoxtqxW3DBE9gqw7piPnVEE9cIO8e8Z+nS9XHL/yDXfBTa8Qtdi96/LBy
50GqQ0sulLgcXy5l7U92e+4cR4gujm4tNy7OlirmFwx0ATrHUm41L4rwot3NsUF+
rkeUilOt436CnzB7p6KtxL9ihXOmUAnDfZob3LS5jEsFTPwnHGzPcnkyOcksUcdX
W+nsfstsv2f9NTlHWXbRpH2zfarKo2h76sccVBbrLhw/xZ/QYS5RPRVzrb+kgt9y
cMx03talM9d5PhjTWQEPFPlHiOo7xyss+xBRvDOUQ8cJKu9ZizI8SIvlmg7UtRNE
VPEmd+MkNscUwsqU/65WhFv09zJcBbw2/tEcilUa+z2pTehZJXg/J/0YC76vSVGp
N+h2I+5T8f6LUN3FK4egA74U3IhI0L2I3TjtLpW3UgwmEyWYPx/meOE/6kCuDgmr
6R1SigqwrPQqaQEQCpEqhJgRDsfcWLy8tHD6GlpsThi33BfRB/1+5UQg2k6rktJh
mgLD71WTGS82jAlpH9Zy/0dX058J58jrEGxUhROB5So/DLFnpeciX0XSQdX/I404
fMhzrUJDdgGUvIXDkRL+CVsBVzEJOcAhIMKHUvYvdnVQPfyxpYtwW3JpyZnbkmVM
xKLpcJc/W6uvUOfyqgKP3+/E4bOHhegQ75SwHAjbCdofOKkLE8ZlQKG4thwl+ppl
VBfjZ4VcODKyHhpe/oyf4P2SjKzo67/zM2Rbi94wVVyhCuwgpvMkncR+RRhBM54g
B+9e7tXN/1dSzNceQ9Xc9wXDAMCAzHd1ONClv/TPUSjc75OZTKqIDxK0vcpDkYZ1
hR1m9fILuF0WeRX9XXtNhJPKaCh//26JoZsTwD84hoowGRIX/lD/vNv3YfAHaTGp
xPAnXioTsU21jGUuaDLP6kcq4Ykjul8X9kK0rJcARNQ/6q2/ZjWR1a4dOuIFh+8O
BED37USWNQ7KTzQx6oSxZpuUK6HbE97tS2M4duyx7FsIC/fkvaHlk9WjRQ0CnM/c
zRZnM7zbz1WGGg+ASpvxgg7poCIXdw8EftaxF4vLDNM0spy9Sv1BcbtzkVbxV9/O
UgUi6V+fPW0aFOybOZFsERT6UwkuGHozkWH6X7ueCPyb6cXnH+Gxifrkz9y6I/vz
g2hjCBrvjlJjXuGqbGUTpDX0Uh/M25XnG0ut24s/0mOMBdf+BO+ZK2WJjsynqwJL
pUaRYZklt6wqPdE+UPYCDKyoej77Ki2Z7hnzxa4r3PX+Z5xYqnR+Z2KCw7AFhQ76
Qb42HQJas7yM5dFLQKGwX3Y3Z2tuEOCowyXjRJyWCPcv/IZwedz398ekfO+2J2qZ
gWKTXNGoldsCacpTFnKjwLoxFdit+i+X3se0MAiqxnaLQuHRAX5KPDMLPdDj7cf6
lI1Qxgf1R5ibxeHtkJsvknxDS6KGFJQekZoYS2NHI1Dwm6Kp3DlRcKB4AfnD8CwX
Ew0F4XJWTATaRK3V8oKhB3Qv1Zv+1nyD4TJN1n9RK5WrjPssI+L+E01u6UUxzBVC
iJvC/unL5I4+7yBVmTx9yFeAyr3fppXZ6KmPBSu0z2uZFCIBo3kr+vQMH8m7wLS0
/pN56a3KoxorlTm0bEIztxLBucAxuJO6SejGySKQSkDTkt9FgfDmXWp3mv37eb+3
7mddneuoX/+++4hQ+xxwt1IzwtsG3omZYMDv18o1oYuPEVwB90ikItfDdcgyeokr
Vvv0XSS1Xki2JsdCjU7cwZoJEG21Gbn6hd6od8lBCa46RATnzy3CaRt2LaoyAoLF
atci2iXf7eg3J3xh4NLkwc1/54i7FSkskI7GAN+8MZZvcnxIbrAURgLcfeUjzEfb
05NvgQJk3qr4YBlym97XUd8R73TvGyCK1c/O7Y0mQ9DUGgNRfhVbHsQrAMP8dvAZ
WYuQwMjbrmI7Ifzjw8L1nVl8k9ZjqFndsySbXiwiK7J+ipYIfwa8Emr25q6dFLoc
QgjOSDAlpFgCHsz477oQufM66OJwp1dNE7BgiwqQKc5cPsAc17KDNOtu33hRPk5G
X3iqXebGNEsoy1MO/g+HokLgHeoq/mTvySUi4+bucQe368WO9zziQvFwQFtAGumH
7Ed8xuTYZmYq3Go+xQz9PnmCJpR5DWOCf8H8liFwyYRO3Q8rQ6N0dsqz/VwodmJz
vdm8R3PwhmXWVPCq6qikHHyljix4P4ewEiFY54cwRZjfWckR9OBtiFjr7h8vrQFY
WjydHebR3U28orC7XrDrPJQGMdcaxxmcARjSgF/N3uOgcw4K/rSzCPP5b8C0fYy4
Z9Qi/GyO1l737gZCOsWHtfzP8hKhpHrJAaMUtz79N5Gi15s9NguebL4cICY5yYqn
WuqxS6kX2wfEdTayW9WAD4t/GMCIUGExgwT0EqMuVFKIuzhW623ysJ1pUGHtX+Zd
HK5z0/ln9iAzOmLk1pY2p6EdaO7KSU/aNygsBPeXkg5GNTqlBTNACvukIlwquyx6
UJBiL2QJigXOWd+IeyhLIOCpVUyJZ1qXyMZwmCx9hx3xFTaVKeTTPxT0WJdZv9OQ
EjqnTj+EauqgJx2QRIhyEcckhZoHyDw1DnWu44l6Zm+cOh5OBjroQTxUxPcg/JAf
WOekNa+UyYTtPvfLTVGxprnWUPjqD4CZWmmU2kPi66zHZprfVhtlJZmDdoeUJ9pY
ko9VYOxyvl+jxpuaHKsCWT8k+9gBy9omk4Mg342zni4UmuPPrpzXhNPnClcfygSp
3WhWbjCrnLYU7tvVsMxQOBaqfrmQx0bcLUukMJMUkkQMravbiGm1GoEKwI5wd2OJ
FK4uZ4c0uHyTj6l+VcOZfPCXrAyLpBzgm481kK9ar4Lgkf3aJKVMO70bcAc+N9Hh
i7rWupwct91Mm9gqw3EQ0TFLjZWNEOqlbaZZ55IZD1Klk7rTR8Upcj2T8AoHUj55
NJZCg8Sor9xx9DBHrYy+Q2MpBSEe0wfKPLguVbuW+ArH17JLthNplJtdXy6grw6l
w9D7P/t4LRmaGznWCBLvA5hCndMxsQDLHk09xfgX4wodTBU9bTYUw66lSXA+/A5E
1jpapRtnD/yj1W7VYbrHrCkhyWlWMo1SLuZwg63fVuSlaxXDUjjTR3ZxB0jwZw9M
kursy49pFjlA4CcnoDGcHsz6RF0TnMQVCvoRQWy5yP/6QqpvYRywrc7pZeZf5tfH
oZO8IeBeMHFfqwfZNGWEjQ8mG+hFZ8ETg7S+THx1j+SGMrukKcmGql3aaelR9Hv1
rlyh3YponZt3ivMRTDqTPfb3okhlNvYwWk3rlA6rcjLPulqLuEamXcTqKV1PlaIA
T11eBylS+90edNJXpUPaUGxqxb84+MW6ZKeYWRRi8US84dpf44occqwuiKL/Pe0J
m0xIXPdgMISu5xPOU82nuXdFtmV8+QQISkfLgr6psYKZYtBXi6auR+hU75KPJQK4
0+y0aJQOt42wnRlY6TJE/5SVQ0iDGsHx3pFkkpRBi1dodhQialdF0IbUPdbf4kcv
fM/SPGNlAx6C77NpIyaR+GEcnQbQnCbMIEtLotSRhbIWyAiH/fRdpWZCNWj9ky0i
I9BkQnskaoud81KGPGKvKtbQsatDpK5mCRLCDNR/c8E74Vl55/FXLhAEtnAsmaSR
fUQbVsCnHC+YrLrcFnaRmeaKdIXcOnMSqGAzq4a2Yosl5rkV9tUl73zsK8dfjCvS
d1SCCTncsBlTD2GI1PQw+zT/J3rY8zk01bAGNZSGfv4wUHUTfBaNTlbtARcTik0M
cC3wBEA/EXnT78eDE7XOu9IvIYhCGUBC6G70gbjLC4uvLY899yKELKfNdrvZo8hw
pjQBd2D9SgdLbMyKHejTQ2vLfpgaIfR89IQtgaRcWgZyf/nHHZbMQQSApcyalPbV
bk9Fh+RuDV8+rQQkyIZBxJE+Q3XTQyCr3OEGKOPE3imyf5TB5ABEHFxpUVDm1fOp
EXSGnAaBmiC8ZeGcqFKgPFvweUJkhERY6yXOG7jMMfEMMKZ17R4SIMYsmvWaeG5i
FbaehNBXg01y12caoV+hlhtC7RQ/9hrTKwnfUzdIyztpu2xS2AbNf/5qTDjHUvFs
MMEis6lBYaHzqNrLKnZ6WaTapVtSIRZh61i9Xd8ApzXxxOstzHmC62CuaTkpEjDr
CTyfRpc1V3XCHrb3UuQLbSyOufhmGahNHe/o5XJd/h4wwacpJ9WrbqVLvZoTD73h
fLOzgmc/kVZfpAKFIzCff+UjtUg0NqppnVtZj0Yx6VeDOtmZT/UyDOJerjjxofL0
3gB1Lhr97NlrRQqn4mRCFIlTdJtl4jINhBqbGfR3uhtCOWdDM34n1WTwDGSGPVwo
I2R8JE6y35HeuzO+i0cuvE7swn0TGo6tLNMUErwImYYAXZ2h8By+4iIHoJfFuedx
i+sv78Az6m3IFzSOklj5ftU9OtS3AaKNqxJKVD5F+sj3dJ45+9LnCqwuG2FpPyiT
PZhJK+5E+zrcjIoiZp8UdMjqdPxFbjgQhEQzjoVf+FvknbDKz8pvQOYmNLcx7XgR
i9ePqICnhfuDhN0+A3bZAojNuOEMbe77PVLf5mdiBgHTdbeNFULMa7//TTHUv1ld
H7eQP6pEd+mz4FUVlZZYgEXXhDqvQ02uhwxbMYnMCzszT7wjzbQHdPfxfWHG9ZBp
N8YytG0gFH0zD25aL+TI7aM1fZqQmwR/oZ309xFsInvTNEMpKEf0rpWplCAiyv/Z
S/wb8hvjFHG2frFMhgQaQ0f8yNPf6MuPOaWoxuhIqv+0iwuHNpfvoB3ZxSWmJl7g
d7rKFcQ68xyazv8BJ1UMXxQMHJakUKw8CmmaqcX2bxznw8XtFXSFvt/bsCA5ruNb
JiYsC7qLUhjO2UIG0SxB4/iI16DOtyk2Nnp6zMHDL1SYbmJF/URwFmv4n39C7Wua
Nqo30dZ5L9CV9pHgIVNXHX/GLmwvE/45A3R0tByy5I8VVYbQmHUZ5MjUGVJq/lVh
hePdGgOIo1vvBk3dCB15Npwdly6IPNDlsDI0WOzXqAljvPG01len5ey8m5Se1pct
p2jwg394Twk0D8kvUpo6qIhV9839WedcQW+pxetCGtwSRKblWYZDh+szhYfirmxb
o3DcUTjavHKEgUDIhJKfXRyA5Bv5YxvlOckCycGXpWxrCUoT677AyuAK9HG+04zy
0Kw3HjeK9hTpyw5f1qBidaDF1Zc6Ttp6a7l4fPI3wT1viAwLc2CjOghi2OERV2II
KQ8ercL4VIqcQT5Vt8mD/Hsiyxgpbx4M1ksgNR/6ZFUKK7kmIKwi6X21h6XiRB7f
usN3XtOKkpY7yrzaB/96TQF+vRaFzuvqsmS1V9l00JYbqus8Zbqb5ewabM6eqE1I
q4xjvDnPptLDJk4U1V0Hg5JN7LVjMnWspwsbdbW9ANUFq3LLee9Mm8eZkeW0GsTN
yypduBvpCx1AYP0JSuwBh9RVn77GzPjXVJN1X8Kv/OWkEwViKFNoRJ7DztH4n9Sf
gYvkVcxQBhrTdAGKs7bYs8nQSMdHjcddwpZP5qJCnFzL47P5CUV/RmwN4Ct6Fu2P
1+fLMmTpDhRzIFMDncEJPulIO+dRz+YqJKufX1p+AtUGGH5Zy3nnyBvep49nohhx
eLzkYWCAzXzRBkPpAADk6rAJJAEaTFlkiBK4a2n8Ic7NPw3yn8jt200W198Gn22c
31aCSdhlW389A3F7ei2RMY8xXua048cTiMGzECxzl5E0vksbRv/UWw504OCxrtjo
YlfULt66gxwh4+q68thbUikdG4o4xgdapCBVl0uq4pGSGXag/yBGntdfc30f1bqQ
p2L1D+8wuLhAooKLB9YahvESy8RBnChXvXKIzWX33syaY7o6zUwuXIOEnUh4U5JP
bSYsqEJ9e9miq+eLPrjDQknOLe0hJTNXBeY0/MfO1tA9hKakivHL+YJurLf/iEyG
GyqT/V1LxrTQTr65+M7VLFmGW0DSovaWCy3NC2/W/aIz1R/NGyeUZ4ato9B/wfFk
3cAJjogSJpHq2xZtrUDmFx/y5iO34PRVJYsYW7Hpd8UrGc/tyipVVAlBSfgWM2rq
izwMl++dOMMcuTWne9WlLx0XFgOXjluoCBW2Ya+e/3Js162oBjp82g/FJMRChf1h
yfUozgC8JCIwIg5ysv37S1Nqb8s74n1E85XXPvGm5EaMwkAeei3vvMlJXVpLHytR
r4YyMkyF4LlbGkLUI+2ExR1Cm+XRW3S/uCmkCoPy/ByX9/atfCnVPK6wpwIfEYVq
uk0cxfulwc9Sobwxd0tRIy8VR2lrSVc0tYoo41P+Hwv4HbpGZKZTjWdItLM17lM+
UIZF+1A7BNtgABcgZ7aZE2YoOIt96JgtDUa2AKF2YLDBan40AaKvVz8LckW1VD4A
2vb0WK2DPDJUIiKzG0GFn7ABjb36slqHida5+oHM9rsR8Wox9CA+cJZ/4WKVSbWh
nANtG+grcC1ndJgO38jwb00OJvMKFs41hEIdCSNo4lerBFzxhMxN21WcqKpHpRDd
EBRsA4Ahn/s4cBkjBsTX4+NhZPtFmAnJ0AwWORnlMuGM6s2vsCLdzlR3d+4YHDFC
PpPjqKpxlcTwQscO3/WPY+ZmXYHkyWbEDW6NpSPQBAOJUB5trOnYi1Rl7WvY7VZi
nqwxtbYJJeR/qpw7YqxbnGsxpWwqsbxgZZTz17ZI/KX0AtmLnrE5Dw8XvTROpF59
5ntnjINVWJcPBAmkhPFU5wN6haK+prb7Th3g2Kpv2zPWTQs2yS1hL5rjtlhXC1pa
1+26Wcwb85a4X2jOU6wMZ4skYfDbmBLHHgUTPQ7tOcBTNgfD+3uV+N2fVb53D+TU
ae+az6Et3Tuspggfi8/RvGP5YYiri70gTPP5SVxCUV0PfXk29ZXOJPVKXZhSZsrn
7md3/DfqRHAKmkc6w5IPjldPefBrywNxmPelg5yZAi0ACabXxjciiykR0748aPMv
v2VAhQbD4gBuI/LrAqR7x8FW2XnP2VJy67/gwVlcF3atjR3IiqzW6wPEX2WCe9KN
QjadDg5ZPX8C4fus8PWOTQFOVJFp7ZoWQTNTPO9TfyM/J7GLBg3b+lQ7feVWirpI
g4BHgBI7NfRoF4gn5UKwQJSeoWfWMYEEWBNU4cJNRyypn6XShcFakns+qiEw1f+h
XGSJtC7AOOQwkSI2NJl2tP8/DqhDefGs94HRZtdinq9nYzIq00d4Ju5uwQcPRXgw
rnQ7RhVRmPzlWBuXbrv57FWPqqwRnZ/6BqqMPdX4vnhghin4AaqhJc+Hj4ft/D0X
x2S8NJI2NBLb73pZKsAd0ICTgfRxuUCDKpOpMQObmO76C4o6+Olk9fH/meeb5Gq4
kQ6muA9GuVbXkmB6xM4BNFduwxcJNeZtCLnAsu5zbwxe0CJDGGxLnWYnwDB1gjM1
Senn634Dwijp6v4w5aiwxy5PT7Y+b7NzfCHtK8hQZ1em8cVvOOdLaNatTCIfJ+gq
T98pCIIpR0MHdqd223+p8V7DDCaS+CC3kc+fEVLlQc8hE2NC5T+ABp6QPoNU2YHO
6Z47B8mRZmoKt7wqFK2aRQxtSE+TmM6zhSEsWWELhRrwfAPOliLMY2Kd6WGLqJYq
0Jh2cpxTDbiRzFb/EGoFDxTsil+dKoIN+bfy/tW6lvsfXuZ/YS8nZldMBxlhny8a
vRyqyrt5CEMcfCPCDB5ZIIIVXl/sS0jc+al2jBtW0TFEzbKm/7CInRqwF7rQ+dzR
5mZExoF7n0Gh5cGEjiGeuk6AnHOFQ5Y6pcsfoHSXbJqzDc2Yk00Y0Jy805vfzDTe
Z72a0RkPxTv9DR11OkB4ZlvfNNIrdmb/bDBsdG+0rV8cjsXQks+rWUd1c3IIaFP3
H1AnGcu+HCwRmwcYxj2IueW4ksukk8EKk20QURKTM89fPivvkptTHoYWWEpLjnHs
mS5HEtV6du7rMh0si5bIx3oW7YX7lLBobmp8PEge23Rdo7VUAYk0oM1JMGMNK+3w
nP1URcvHsEV3cDA/iFx3BKZW0TiZ6xMuD5xd1BYCWl7GvgS9kCWEv5cv/xbjvrgr
1EMjriJ5sw9JRfBuAgFuVffbc2A9EfRzA8EKe6CeDI1mJ1NSXLFFX3BoI3V9hkSn
KaT47rR93Srm5PyyTkcWESXul8SuWD1c0JFnwgHBtmnVz43q5qqNDKKotLPycyh/
zx4W0vfxi6ws8GTrpIyGopE5VCPek1vj+CWwby9iCE7XoDU8IB/nsJmAX6jH2tLh
t3FhO+V02Tx9dm6xweNqY6N6tOsGsYVMbzFtKmp6qoKXygQSDSWUj+aKD4zesUOz
WeV0kagYsEDcUhE98a3qKJOiQCG6WyAZ9Ae8Ez3OebotXOKo8mbUmHY0+rGDrIcf
Q72ovnj6JxAH8tQeYL5Ok8jegZ3lwo90HZjcniRMb8A8JpGyvcBHpwszv99JDETU
qGQBOwYBOswlGbIOCucL/7prUnfIuYHk+bHDR3Mj06889ka0OOwBewXmXr2iW4nf
Khkxr3sUhd4A4zotm+ODII2lpvhfBm3kHcqsnnXwaUcCF2TU65+BQan1OJ+Mw+by
b7xJmR7gl1o0KJgQDfIJp0/fM3241rnmjuJYjkDpRVrPlKUngOAbTx18RTpJDm9e
WaeJflbVF6OuEuIrUQKn9Izr0/nhOX9LjqgMXjEUwLJucnAUKzsZShPAf//xpOWx
CeL7uCR78BO167p3TGDwa/RdJtnEndahE+zUvRzWS7xu81CCu5wiMl4v+zDGvWy/
CyboKA5JHijiESZwqENId/uVMVvCRErBTIp2XWvIDTCVfNQfKIxjTEpO0w4dmupW
SUfbZr5zTUc5PohlM2JSB8s7CMfOMshrzJBDmj8/U49a77pB+obIJ/zykOOPg126
IBORi8Vq3ZUGi2Wg/tJ3TIVHRc79vHbrrxiq+XnXWq/df2uPTe3RTqn16JusLiMM
Q4xTO/Y0KhlbssNzgQQC2XqOoTWSb8UPp4UHhYLqXXj5FloS9qew6gm+ogLf2lus
/gykO0bTCCMui6/K8RwPzopLasiLTB+KHCmwUVMg63eY1CnNKNtZeE4yLDLmFgJs
WYalzLeLChg/BGCuMLHnqVhdzfPuP4/ETvbt0HbTDAi2BSzU4A/sNZKopsHQ6p3I
wxS8t0FWe5Ko7aE54JiQ8WeW0kpCQQZSEvnRwnYKQu9+oS1UsTYqGPCGWmqswAyt
ji2/Jo9pVflWP9OVxlGkPnphir0OFJnJ/SO2JTS6Y7KpoHgVOGG0x0kdrf/F6Lkq
J+wzd5yoV3kQMEZtI3vuWKbCk0kHpXIdsWxbd7QJ07sPrZtIkFhhB3aCLYvL3wic
zKlCCHRADO4maqvRGtiWv+Kq64/xe12iGOJKFv7kTknOmPkbOaYND5cgd+9pLi+S
zWXUpjaLGzWUCOEcyXb5UzBW+A6r2tp/WIzc6nJiXKKT/Hz4UW19EF8L7b028nFN
OD8Ul1aaYsU3wKkYDh06B9+zEUMyIEHJIAEIKy1QevSmxNPT9kbw74xI80BJjSJ+
esNi/Usjoj7OcNEabwiOmq5jCtdzZSSiKh0r5yfcYS3Wos+tmWXraTQGgPOSDMeg
A8M48/N6ex7ShBioNEWwvCJwPiY5aNQ4wxl5UYHPWuRGKt+2wKurrE9xm8IVZdnt
jtYu+TTL9RCSea/G94wZLwcPiDdctnSGc/eR0358tRNBSyRUAueoluxxEvZTokXG
wa0yvgABh/JvfVbjnIski4yZSFwKUbJLikrrblTuuhmxUlzVlIB0vv66p8DNLW5i
5OAKG9UI/1pyYiyxIk5N222mGeMWHMkbEPKiLnZNbkr7c8YTzcpqSQ49yCrILPI0
Szk+gw4vSb13hTqRUTPpbAE+ZTbFLxFrHpgl+EeBZaU76GbbHu0HPlBUmJ1ivXGL
tNsiOcLJY+OIo4q84tsWEpFOCU+LUyFKgTZEgmbEt/vM3B2uBoVsfqddvMgv8j0e
fjmODOaBclSBlarTYO0ctxO01n2UfG2r6yXEoUMBg+K3Dnf4t/QeoyJjmgMRfGNv
ysPdIFVZ2h3d8ISU4mE+4JaTFzZefuxBmTAlw/yOSIDG8asFJ1j9wnwAOMhJ98U6
9wQfk4Adlw8lnV53zHC+9yQuPiD3xZmaMOVMMWNna1eqSrzbvifX+V+mh1IQfXE1
3slHLGmgQGxWFM1vGaPv8PkkijZYKUWMIX/VaXV0PWvmgzPc5C0ZXrYJbW+FEhTU
lCbBwLLBM292c8l8/cyK/jHHr/xgrsUGvNBiKtAdEC8+8A3bqJFe2LKGcyqB5tkY
9K1Umsndfx+b10VkMvZ1L1vMyPGhf6N5BIvNQz2tdPNII9/TAcP9tQJUCdTv5SLH
M1AhTVxeOyw8XUyIted657FotdmPAXaP0TsF0Tu7pENc0ypMoK73+QWUbKjP0XpU
g5Z/xgAHxPVaecfpmTs1TbhZE3Cf3Ihstnq4Dw3SHnogISP/P3U18kawXAPu9zyy
utaTsdDByHnKBpHMjfNfOhblm0NiBRin/5QebSaXkvsRSGbDqlKMDq7/BHHFvtR5
TS7Jlf8r/XT4GN8vosjaW9E4/RGWZJWFDAMqsK8bXozCeXMoN2sIAUsoBHCqNBdT
8cHVl/L87gY/dI8RRzRbYeeDUk6/M0RDZrta7lRJzyaaLSEwYRODibA965TW4EUn
tD7tPZquD/AQw0y4etn9it05uy6a0Aomlsj4FVIpAUrxUbbUiklln8Wsb+7nln+4
f6JckzITaLLwZJk45L9JLfEQ5d12ZhgEnC1RVvY+wo24GaELAMNmmSF8WgfYH6Ph
UCn3q3hQ2a7P3lYTnGeMvglzMZVAZy5xJgg4He7v2Y5XWlC5mHFIOc8NOsgxdmqN
M1i5imn2EhyxerBY73ON0oBRI20yms5nNqU6bVvfk05hpdJZkVs3qrfU7nQTJKyR
7LBqNQ0DaORaWADk26iQGnndl+lcigYvdzNKiv1AOophxutesGwP0MrN9czvHxV7
zsUK8tq24PXlBQWALXdkgxxlhsa2Q4rJBTx0bzXKfId7xs1vsuLdhWYfQbM2T+ga
rwzxRW4pItY0sKcQNW9i4zrlf500VGnUEuEiSxKdL1iesyLjT2cFsYpO6kyUXPWD
+F1hzgLN1RlpK7tr1Fu0YvyJ3c1hKiIyTp+c+2cWYYEGx0QmmiyDCrYySskyB0s0
WBzHr+5nyGJu7nvNu7emgOHfsP7JTU9Wn11MA9RdYIhjsfpRbkzzcrUd1DqCkRPD
v9fUKA2h+lc0LowHsse39tuqHk3xhn2bxvto9gTm6O0qnuOJp5Z6TZ+BVkQqsYrG
Y7OIW9UG6GQWSET3+21nRK1bGNu2t9QfLcpbVgcSpjzRZkj6ovJw1ToM/nYZFLQ7
y5hgPWBmB4ydHwVXo8rnspOXDDWaxXDyUbesUj+WXGUeZbNro9P+eMPMp7+LNpAw
v5tknfZ78nSKvg8p6+Jwi7K9tMCzVszYHeHd8BIOvOi7hACUBmQRXRSavKY9Xa/9
ZC4UFj8H7pDPNUzwtXhj8foo2axMkjntOqvOiDPHQqL6LvCvZA+pyCjIHF7095Ji
lFJ5vE6tRHZ6Y36wCs3ij9ceqpm+9FQdPnAPgJHm3coKRsvcdVyuJjDDNtb8rXtO
ucqsFcyk3qkpipdLaWbkpa6mjIPTmTCtK84DbS1JHFKkKcRLUGPOY5b7VOlsmkM4
2dMIUM1V/XEapiHNHryGc485/4x5nYYJzN8TNX2grh6jSHeRQN2iZt2vMZ0LZujk
5ne3Q9vBjnSqUz854njJPVOBS+O8BLaopoLpawJ8YLa26IdkKMByOnt2UZseV8it
Zpz+wj/DF1x1ph8V/CGPZkKjbilITHFo1NpR8PglgQMqDRi8fRVzQO3cqT1w5KL4
rayscSuqbi13P+3T2+FALUfidw/wE+fFWPMqjtG1ffVuM4jMNwVlRd6EBluLb75w
KNBXk346Eag5VZoNkSzDZLlUnhQJkySRZLE919BZRpw7lyb85uu4UnRFTuL/uuAG
oqbUQCwWaprPDuk5NVf532tIrOU9qS/ixY+AmhTFnZ+PmtEt91t+watSXs9nVPgj
49emIbAlc8n5CvJ7EMwPwTO6KQMEgQ6H+D9bIJeOTrFqyDftOEtjvPiW/0+R9mcY
a4Vk02MaiorYugngM8XWzJ9yvbkEuJ4kb6EC7CWehA+TsRQCPLBU5tx72gruZAgT
qBoEkJfCBPdVuLxppbqDU0/ad8VPp9jgR+8n+zznQLjz/oD09yC7bKmI8C+vE53J
W6c4R2QMUTp3J1RemtJzAyTgjD2Sq01jgRlknZ7qT0QTcrUkN5qTEMbOr6SrPh88
Vt4TmzGxv0gfWjzinRzOSaJli5wGViu+0FTrnrwSNSHuK2LSn6a2VxnOi+Ht5OEQ
mDfjHPa86IffuStSudO6z7oQPUmQG0Vb6YscJQZ0czbZKtNzd9bEoB2PuCsKU5iv
lQZNCdh6MXf0x9MV4hF4roFrZobqJbp2XFOlss2u+ts7XnDEhS8NpaT4WFN9rw8a
CWG5RpZ15bN7osBJmkQBVM7b2xsrp7bbMf83Qvd8CcZQyBDImG5+QryaXYJTBAc8
XMSWmOpn1CNe0cLLxm2I1gnsdthYUuAxcXj+dRrFT3pVjlmHuchDlpvryitX/044
FXPd3IvlY7FV9/b6D5zJIxeEGR8T9Pw94gppFSoxnN1RgV7GzIEvO51Jq4UavemB
DJQ+A1wb52fz5OkZDyqA36smzeolmc5DjeYdW4n1GmkWTIX+xbve9lViZHLT5aFw
G7Q/rYEKOWr1iCfxkhl/cIQQ93F1guLPqvfdUckw2H5Mi2I1vlR2mU7tMbKf++/x
KBjUtas40gCb9Uxx2euNlv1ffLVoJHzJGWxkc4WbqOgHvSoCPsHcsZUSyNs/NspQ
SQIKH01fUHlJC/FdL+gfTfeE+Tkn/pgEsITafPhFg3utAO3IX6bpjyRFYVKfxJ0t
6CpaMfhEBk8ZicctPYUJ5h3W0KVaATuTmpYu0aTAi/DQ1g8SjTA4BZ/TtxeUGcaz
6ZSCg9skEpDleI3KclPGRwWHJQXV+4Y+cflfv/sHwrF4D6HDQ3tCUBCjAL/uXZZp
fRO00WEyNYz3FT0Eeu7oEt1E+F/dYfp4nARHM4hT8OsY63nIXCh+KmzU+coYFboT
lC7EXtzymCNy+aBzaOKdAc3LM6ma6bNP9s/tvNpc/EtjGL+cgDIRx0h/G1r5m2+t
H4249bqwDE9pda4ARMfX35/MHCkxR+AOvJMRafvPDbN1dk5W6Dv0bdxk5tnrnKM5
XfiQd4Y2Zq3WF1uYxwaQKP0Tz8jYbRmAZUVgZ2FFLfCLiTrTKFA3xcR3R/xHAF9T
P1NbrFObU1FeXxSyTopMhDoZlefqnd9gyRdxh6SmAwBDJ2ACx1tQKcjLVK6Xt1Vj
VEXaSqAtnQboXyxGEmS84O+wZ5JKTS4wCXotorQ5nyukBAhQ2JxAcbkOxB3frReq
y3hQ3kYCBhgB8EqVafYjwf2TvN1yGDffqmnlEmG2ypqEaAGP2iN+Ngl4SBa3ExY4
iSyUebJt9uOsB/l4gLZy1UWUtTNqGUqdwXlslI1/tvL8OkLUVJZWTibkEuyNKlFe
iUOzopSDk3CsWP9iEhACvim6bvl29eaDMm3N9XxBtwPMj4JuB35ll/+DogX7a8hf
TM5y7R4fk6eFVMpCJxto9jKzlbnbl8MAK6/pn8vy9w9/z78PGEtAL8pqQg8w7TdF
7oeBy8Nj32uOIO2oyMWQs1ctRO0R2bswAlSF1NdLS1rYQB6lcuc89Ft8uoGMCTZ2
1LkBrJ/C1FhfqlN/iP6M+WQJaBLnY+xlCP/a3AySJKm31LlCYLiNVPlQaJ9OG12L
sisw+aNtXAl9dpQZSNIYvm9FpkQVMNxG6J4hQFQ2moArFE/0vdqrlpQ3S5jjKIPG
/RqyVegi+AEVgBGSSDJcrodPD3kSzXuSdejm0rPsBMidgMLhpE1V3HAdLuPfUJsO
RBpSZUt708UCC5Yu6o7OYIC1L5WxTUICq2b9FQtobxwPV8r5aIAA7VI3GbuAS7J1
jbiVl0409vQ8AWDLPmVKsT/EvEA/Z3RadGvAS1cnnviYh4YUXIMRKtQSHnRQqjJE
5KESCzKYlyeY6Swv8YBpwzrhwyQOnyP84R0QoaaqpmMsDyAP+ov3Yd0XUIEV9ypj
6aEev4+Sx6Eize1JDuT+8KUrJnRDOa7eUb8nflYhoxZ2x6TjoCZhoKzaYZRrUFJq
U+doo+CE14DhXIhmJQZay3KgShenNp7JSGIqYea2LfffcxY8o6tVpjvipB7C55Hd
jHc2bZv9Euo565i971OM40dq5r4kcwIbsmaKUkKb31aKJI16DaQxSkxLBhRGzX9U
xM5WjJxVLVB10xPJjElEQjnVf1I2q/2lM6P1lVtSFR6/IAjHzHJOIpXWfuLIvbaF
xcpAU31vP9a9X9T9T/5jLU5say92eqg4YM+F+cBpMtjfn6kjichiGHslOoT7l77b
3Z87gpzxQh25IvYkj+gYcMiEjvXHP9kvHUZ6//CE6vJd/Ka11xQ2sdYR6P8oQhn0
FuO3mj6gy9DgRo0iuFgqU9NAN5+BhgOSgBs0LabNz+UodzJ8BGHrpS76QcieWhpA
hKOu9QbdzGhlcuFmFHFqk7tpmoMFvhXgx4+cEixfdRR7eP9DLU45yh+8JRd6v/+B
m+R64+91n7zoDbUb5tc/n8vE3RJTLAgBu6wURr+6/TMHQmOJKbpLsLu60mtB9t80
AUuQCZRr7riipOd0O4YDRDkp7V7308DD1qK5ToV/dk5VkzvO3MQbrW24lLlzaAQo
VRhVYrWB612WO8AbnOu5WYcrafUagcIAtplsPlCYdZIUAxDTVkvmkmVOnflFZyOy
DJfCuXXW/oA/EMJXtRpIpv7HZKKCsPb25lDQ0AF7Ixs2KNFWp1XVu4WqUlXbNAc2
9gC+hywlVqR8WT9vfgMfVPGS82vGgbx1Mw5JxZEQjq/TIA/yuNbmsig6LBp2Pul8
UO7pQOlL6C0wj9CgWZ3EYKcXlO/Jixq6ncMFnXUUXKpSGjXyfc0BvVB2hdSe+9ta
FcxYYO7znBCs/AFu42xkWvteJZrWoK0lJPyt5bO5X+55qDY/BPUtR0MDR6nUtOMg
7PRtGo1yXAzy8niX1NV9QTkP/qa+PtJze4eaVTUfm1N2aCVAgfKksr8Ir2ZiHEKW
wUZ32poF1uM/H3Mx74bPKCIHKKquFLwAARf8lxWyf2p3ZBymVIXJsoR6tEgSGZGl
NJiYlwzBl2cPMxy26oQqGfG6OkxIvzdsDkWQrZiakgVbBhxPhR3zPoU2DmmjsPwN
rbEGkBULMulz4fF2BPYf7ShqaWHRodpBpZPbmM+DNAiwvNuF2EwLLfDc2U5Z6UxX
z68p7e5ROjEjFGWKAjTcQWvoI5TX2EgY/nKsqoeodV4Iy2kpfs3Fx0BLonhgES/2
Hd7xHLL+2n2n08/8dZh5APn9+0HNWotIoVd+7LF3NenVRESrVbDWHEzVpwp6Bjlp
9hWAgvPCBU6hc3WAEm6puw5/nLihAoP7mHkUg2x3ZaW1/NnaLmJMT2X1F2DqLeBK
uTKYXfpO4WxYmYBuuUHD6AoXXAkHR0cxi8pkXQht8qmkpAcarxwz2iQiEUw/nNM1
S69YTgeFBq0l24e1C3+l0dVoSmi0JYgebUl2ENRTWIEGIB5pPmXtUrZ+PUvsvT9t
iFXqHzLtaASGS8CMs/6hXnwQcW0RuQXpeGkmhLti2z+BcOYNzbYa2deejz7S1c7m
oPTXojgf8ec5ZsGoO7zucYROLzqZt9uPKLQtklJBskIsCgSzaXuHW0w2L8Uieb8n
xmiB4G9hJlCQkJiyXv3Ht1T12vyCoGh2K3djEbDkT+sJDMzvGvMsmgVSBtXYYIk1
9LJgggAzoOQvdm58jYbpldGT9x4kjWt8wF97qPMkv1Nz4Dr0tFQagMhml6IZ/yKw
Pi3GHxXlwx7qHjiLiMgkCRvC2Hjo31F+uuuWdgCleMNoB8hQyzJBdi9Z4w+yPqWc
ZEYTuLApvxY2Z9BLhrPYvGZavjjne4kUsUxIjXc2oMY2Q02VEpWMcSs17bvtfjyD
47b8CI2bbR/rlGCQkTkvbH27oku4Hjh4xaC/6GH24rjTx+smgrTRKtgQF4dd5Maz
oKFAF83tASEGlDwuZwGo5qo3c0Un15i+gY4G5MXOmDOm9WyMjdQ2w4UjAXj2NRGL
i1qiOsESzpOnkVhyRiykNpotXw+FfDSZIy8Z9zC4WJjK9XGwG6jzIL3LJUdgoG02
Bol1NF14dFBsM6VJtvYW6gQIJM3yRD0QqQoDmQo9EwdXmn3aQ7dj+qvbVx1k2jQD
Gn7GMZa3dghNo9TWVzNuz/7xLdkoVLHVIxIUAxjtLugKWAmLMBosB3oe7XDdrSB7
lvEBjBAZyV2Io/PcqH/odyU2jQzB5rjyzP64WxclxOLRs2eJLcArTrushmgo0kXA
KV7ZW8/gWNyBBEpc2rYy7yI4A6zH/GY7ekuZItKylLvv3JMVK86wqFxp5bOgRKL3
/6/DGVR5+BZmk+C1OqGXpir0KXTGwPVFzz2sP7tWsTYIOIM+H7YZ+qJgn0IjhWQI
Bybzmq+YygJYWdCEemPzmtJz6vi8fDsTx4+liNtR30A1kXT67tOZixN4pFeFVqYY
28L77b2gIsB+xDWRJGqejLPoVRcNCxUwqhya1EZ22OMXqjtDkrMbQqh1gMhLCvU3
Hf+fEo4jJAJR0xcl7egzjWHEUEn6TUHQSQpeJt0tKMyImabXXQ6kY9UkZewVQVEq
VBpL7QYTSwUc0K2yrk7wGu1aVSlTKPohu5iurw4qdnxn2sfbrcDrbXkDqe6kqkTH
CraOZ94IzGrAmtOpMQDlYyrmFSnkDFc91a6N4kqe6GQFHnmL6r8HE7FVpbClu+Cl
pFw2Zv+h3VKtxsfg55whpS+AmnqN9I7MeFrswG8ZHvJzfCJUL27EtjyynSHbB8RZ
GaZDEUEA+t70ffGBvLEDgL+95meODLy7974EvpLHEL/jQkdHLOzh5pqejMzBKKUS
9zRGc45/n/maeCJyxymmgeQGPAnXqXV6EJ6A9bxzoWVeGt6uTNROxw4FEGLyDhPP
MKyj8csBz/lmyUcJdG+ZhFjDBO0h/U9PyTrZqond1RztX/Y7LBrBid53evD+DOHz
28iqBnbfBa3G1aNi+wbPY5Vu2KEEjOMRG9pFdV7CG+i5XWWyxU6w0r2oeibkklAY
9jwLNOl30vA3kWTagT2nCzlLom2F9XfanVoK+fo+CH3/w82TCYDRWWqtOacNnuGY
44XrKEsl0OGMc1eILOvJwgen0M9lYHDlspv+ADSO7XvNVlwiXlCdzKbEqsIUEC0W
ixXsxaO4ChGNomuq0aG7M4V2NPjTEIU7O2n7Jhf3GvdGakNuFtnVAtjcNCZ9fr4A
mL2HAt8uQmpZyuJV6JVVGhQGtpbF8TmiR3k4mN+A/m84Ph4XqZDerDFvzn3zwDby
VNhvME6yJhBGtz7lACbTMGAel7D5riOON+m8nVEUUtr9Ngl79GOi2t3/aXn/Sabn
mhph3bnYzS/UUdre8+Mlbiea8UtCsBYtJ2PmNEjkTzDb6ZeeaEwB0rwQhY6OUXnt
3PLQepcjDDnH2yjD4NQ9PU+6wSf0RuNLD8MSp117AoIkytCZ2JE/egm+6/bDof+7
tpOc0d8DhQEOnz64GAxQgAgtvpNdidg/a4gsvUaZWRC3+7V9GNIDblUxCHH2AD65
HmnVyVnf0Wr6HnWJ6hvWD97VI+fReYrZA8RA/dzzH/euP3epHjTyi9UN4gcpfZkG
w+MVKkiHc1gqcyOWX/LZOUJgQ+FnZH/gY1JkJSwQmURQhwsOJoDovyC6zMbHLpz4
jhdhBpZ6FWhJtiH8Y56t67nCGZUjuN06cpBOvlLiihGvFsl1568KOYb03qlrSMXL
i4krVMNN+NHtugqRO0dJwmh32q29MH56t6NShWj06A4ixIlx+NkYGxiSRjkdiPdD
KONos37ytMBdVR6wVCeY9Vb6L+N1CLrt3YUww2Obni8Io8jJ/O4VHaT0617mOfiA
QY2Fecge2LDI+oQ9pp3bNRmWdoPB8YR0lRnwXw7jiLQJ2nuZhsaEHYMBEGDXKEHh
TJvK/UWzOpsoo8TaJ2uH4VN0yDn29Ne772445zMUsjcVEg1eIaSnlk9trEr2iNgM
464BMb1OIdcxLzAPI43YyXQWANOv56ffwPuQ7JlgNkd1gD4Cs9lSxIdnvE8Lcg1u
aox5x46bTLo6DH1z5hiGXFHQvXsPNj+CbwS20J0yj2DvegQ/fc1COlpoggXa9Ecb
gS7PINtGdCgQA7SJ47GYIgowahI0jOQ6UbmN2xR/3vuN3RAX4lM/thERQLIIGbNa
My9Q+WwgfElqIJQ8iWhNAXR2DbR3TB2MsSeXPuTf+Xycl4PI4fFmTYI5x7w7oQG+
HHCZOaEJTCl4tjaLd783bd+OArJsHOdNjzx7ZCNhQp4OGBARitacB1CjbSoDAiQO
my2B5qfiDtYqcNCMWqCk+JzJv54IZpEAq+HE+Gb/uWD+J/hdBHwA9LxktwJzCtsj
8vM1b40bj7ggid4a9WmYyzeCvz15KSk4/XJK8ES963utx4B8FPvwxY1TQ/MwwstR
ZIxDcqyi0iGPHXUl2X6j+BQVDBzksE6ipflbu/rJOuFvSJT05BvfRImGEBlsh490
8YJ+yoGn5WncEe+xmw2KdK5tl508ag2utRAvRgJwrnk8PTykX/xrQ00tZR9xo9vZ
UoFzALkorC035Z866+LiyPrzDxzK75Oalvk8M9BlH5kW+/H4sUYOlCqMpuiGgWnU
LIJtAprOb++Fym86nPA6dSkhc8FXLPANn05yYcq/aHy80xGK/mN8DvDxP/LcYwBF
FXQgS1IwGDU7sWZjW7sP1iwdiCkhvhclobpJhlZx3jntx6ZppFwJxeVArtH7F4Sn
fkDVP9Cr36IWifGsp9dxGihFY8oP6ga11c6dwhEYUtfDyb1URrRbnJsXwWCCUQbO
XTcvLQQFfb+Qxp77gzP+buHdXvH2i08d+C0+9Jvm30vd1RZf095jn/OqlVP6rSs/
RjqfvddCYgYQyRGHmAPDRvrKycX+IBoVx4mMssKKsplebMh1p2A12drpY4y5swhd
kSkqCIpS7E1bX7ubswjlWjsTwmnNsGunLfaUUzhRWy+fq/kHtG77KwtWnGfVM2gs
6Z9jq3k3sFEy7b+1fpzmVJ78K7m3hNmnVKAm8yxnU54Yj+q96/IMMXjcdNOH6IIH
rNYFacdfwBHNyYyn3m8SVSLEScrv16eDBWFKaMp5IeDkPp/3gR7oSnGqaEpuRyyU
wt9TxhEy+mF+MQRm1ysXgnpit/IfgJ5ZRgEjjvjcXIrVX5QfSGqPpZbVK41AiYMe
xMMFc+NyKECrMFHFbmu/4le58JJIzv8V97+inyujRFIQoy5DDqaUctrSKlSTObGy
uPnl2kfNH+E8lrSY6ElpnNAQSHqcVz24boenMP3Cw+nIDIkH90iDgogVgkk86hYX
7Gqe9L7SexayA9/f7FBUMhOZ0Ete7j6ApzGI8bdXU4zA4g4Q3FnGCFwG6vbVu3Sx
hVxGGFN+t/9JVsH/sdB9tX4rufHM/pmFWcu1ily9XkedurltgjWlKQuEulcFpE+w
/mENyI/OLCLw0LVZjLpRONG1gM0U5I3gvgUFXiWf/yhryh1XgojqnEgP/xvl7w61
7urPCHQPhuFM6P+JehZoW7juIAhBVFwC9859bt5IdwY1SvVicv8oOw5YBNaEp/Wb
eRAmrXLSM6fyEZ5IHF6xwOln59QeIa2dqScOqcix7wjrnPedhphSqvR/54e2ResI
pjJy+GltAt+l9HL6glmVfGDI88C411d2pv635g1wzFD/MO0RdZOkVKm8HBe4sgtn
DhzZZ6eeM/e25rFbDlpJSRp5hCNTiorIn2qaCUA5Ru2A097y+nlpTVYKVMXZOQEx
qwWAQPNUK8MmLdvGkHXtNOnxTaVaRviytmSLcHHrDELOiui8XE3CLaImpj0ciaN8
DfvwC9iWiY8ootEBmPDhSfQgO4purXw/yLpkOLWWfwjxY/9O4vXJQTayVllf6BKE
/3pTYW99bSx6uKvPRIgyQeXEgCuMGL8DCjF/EeYtlEVPx1utA/lTtfDL5gVBOldA
2nNquJkLkxV7BADuBJnXLuDxyEwTOhwWK/CfbOmTqcWvNAGVlu62L/eHttVgq40M
q4qX3d2MACNhKxQlkQlr/ZPMKM6hEAxtFpI5wENWZqlP3tlf0KyfjP2SJZwC+L7s
bN875QGQ36IXpvJBWOalbSfz8OZhEk55V53/9rDkTvHQVdQKbrDw/PmwEBkzWWfZ
CWv6rk0UV8bp33/S6LvKlGYWTPgYC0EOVRjCnVMZRBW4CoDgNUo+qN19u+qIolVY
MQEkXR5342hND5P9z/fT0r46A7bhSqSJIopIYihBJcuYD3ud3vZeHWytPFZigBuK
W4OUQ6iUimdMlv2e0PSQTcGUyCL18m7Ur04UECccJ3OpWE+97Z/BtM0RBLuK7iBx
ny/Avt64IxLZfNqsbdjHAn9HqWxydIhl8UI6WrogmCSyiD9b+EegiU33FzyXlHjO
tfk/UPWFwljpsccMABkQealTi0V8IMKCLkkt3gNAKsIRWaxolgff5AYIG+H2kpmG
LkLfw8hpu6qHZGd3SAzoD9ACE2td7loMuhGWFftYgXgaBmQ0wEm8jczL0HStksuJ
DEEAsKauUHJ+HQqyth/89IYm7olJmhUz1j3ltt142kkbrZogW7AjXvK0CZ4Qr6QA
WFjkeEQnuJ5u1jN1XkiX1Y+QUWU63QI8unf27kFvFQNbeqTLxgHHJlNu6ZgIQ/xW
J4B1h2SS9FM59ttYCKfbmg/T/oJOfn4Dfb7NoFcuWlG51vuOFxaQ4W19vZS7stEU
e0b3ZDA4yGzekeGBeWhkQGqPr2gT92PQ4VA5qwjNcbg9iDvNynznrrPf9A+/l1ty
uduQCetok95A6dy5VWEmKsC+YP107fs+pEN5OrygqCwhxGSLWkmZDjOWKg/Op5/6
Jy/vxNEFUClhdGOyhdIAaeWecbzjNgmCCeaiSu21kiKmqfpnUY6SXUkGaZLOTcVp
EV8FOIyZvd4T3s2ckxxmcVh2ZiZDauPDC5tgFCZmZwQOdYvuBGvuteGQYCiGLQRN
8aDvYwkGt5s2zpQVhfXe35z7J7lFebhcxHQolpheEyN2hKj7gnyWzHqqgypblNlk
sdVoFJma9C8AmUG/XnXxXwovsqPQmbfnl3iW9qQUjRvGCqd6BwIxX9eGhILMHuMr
LGQc5ZDzyNxlmQBFgnnwJKXxabyXy9nGOkXLdo5Aizn4p15qXvHyUiY/DOZb4aea
MyC3TUtFQ7WazgN9EFexD9hx+XYlLVhAxSDeoshQLi3N43LHM5famX7wGfeOm9hw
DfT10lttNEIHi14ptEaCqI0GSdWhjALR/P54JkXAk7KqmzteASAY9gOg5VzOwLd8
OQNtbQX3PY+1MLo0H9CtmVC+RkRtyZC01wVfdiiHyE6Co7bm+uI3csWtDbCvSW0G
Qvahdwy5OvpHKsl942yTQvjgaUJFA3U6lxQAQPQDw57lVeGcVag7fZNKcXIwtEav
1TvwFQq90GhV1ID+oKNRzx7I54z75Hp40TRUR4UGzKCSAyg/bek4294/f8xj2zv2
DCY4ASq7w6s1tjFe8uSzUCs2knxZ76ruYL0WHk3deUGsPUpUcfGQcgJgC9K8OsZ+
586W6iax0uejv/weHDzcJkktjfr9RFhmIdfy7Mt781uFGC0qr+No1tA/qw3stjgF
E4ukPR1EHTB/lkMopaxu7OGcmv/vZ/XEkEI/gSBJBasDGP36BWAxZpzZQmKgeavp
DZ32uoDdUF8/CfMB4FWWds/DHPsPZHKpKy1r0wZaZ1Itxp136TctOu96NwQxKvhE
nXOnHTw4OPZBcUv65nDFS7OialffMiRYbYmquJelGSXLF3D2wBENDXOEUXK9t26S
+Uih5U10n7cLNg0xmTjEItLJonyTR3YM/EEVTkmRureOkNSnuXwxMIQjTqDQSA3h
eZgSVd5BSM078IECQnpCxvu4jZs1Cuoi/y4Y1gCkNCw6nDH1WnKO0GdWbweYLnO5
1lvwO2NSPRp0T9WBqaj47N48uI92mX/TqBLLFgILHhovwxcqRAfSJyfR4cxYK2uu
059RcH9ueQFEN+TMdmJjZImFw+CKMUQsc+l84sWYXdPEur9gqSblDQmVI43vRQPg
ibo2adGRdfiTOhG7u3P2vJNtG22ENviDTh77YZ2/8KQ/EjYAxuCUcvVf5PPqOShA
/GHqXWyU/KBFgn9ClInQJOTS9coZ0/HHHD+AKj2J1xFT2DzXU48x45rSzmERK13A
9jItLMZCFiogSXMcJOc4wkiTqLV1ArWyFZDCQCAuqk3cDXohfsIF2lmTwjuCuiYj
0J0sQbshy2qeBUwpeKXmd7nOF7cegPH2tXDxOk8cCn/HPX7wOOk3c9y2O+6vmhf6
NsrY3Ft/VD7mH/ZWsnr7NJoA8E+TAALqUCFBN5IliAIWIudOoGRwPd1ExYEp72Ig
N/ZAQ65WdHtP7oPKOBNDhSKgHZgLBXmfUXwh79aWlPN1Ut5KcDB9tK0D4FcmFWDk
6oCUfmbMryQ6Jc7wszSDnOPEQDlySgQpGv1m+m5OKTJy21FthGvzlPfhGMePAB7f
BBInKD5veWnfBdjJF/mcPEYcpA0UCzN5yp/GEDmmFTNYlmuqrXE4tirNYbYB75L7
Rm7UItDXeWiBjddUnhOJtFoaSAEyCtpe3l134QKpJnuW+9gWmToZ2LFvoGW45Jgn
h9Uy2j9xV/0RpRTjibBQgM5vFfLbWwmlx5T9UV3j6y9ACgAdjCarJBBWixQshADA
WdoKc9lPL8YxQdrexmcyZcs6Cjo356tSoMHkE+lfteTcdStMpml8vz974azNM54b
dM5iDSUByzCysfl/T+LzPHFeHhzmlpAfl8m5eV7dzEiRMpZRc6P2hH7XZXIH94XA
SKX2/sG4hvgt2Zvkw9SHUO1kwqJD3cN62GvWa8w2Ba13wlO8mXk3kXp5oj+/g0oL
fGS26n8WUSIzgRLVwM2tgY8CuseGB+8c+grtIJWpo8xtIvPHE2S1fru0EEHKu0sa
5mMNpMuw6TG6qtQcaW821T2NwDDbRUG8VIKsoBD+k1zDN7RCtgpEbpI+NTA+Op/J
8n98goQCj1smRYSpixyjOK60jVje47XaYLCEvbTspk15e7YPu9aWeG4QCu1Sn2y4
uLdDiuH+DkLnj09o4bKFal+p0kJ9bn8OnOVUwECdMBU/SvokMzg9DSq0GhIyTmum
ehkoWfUz/wZBE+o73wH3CsrwtWBSS5LAH+ns78ben7suB9jY+4lXhsl/E+xIQLu+
DJ+xadycm0iXx/5qY1IaNwEOhVDDMYbEhHn3A9Pz5gm6Fa2z3gBdOOlWDv0pZtjq
EXA1ed0RzQK9vAUwxvAq72J0mikYmRJyEI8oMKao/bN7AFAozDH11uDbJXKxZ4yB
0n9T6tk97LfrR66SP70zHQgod1cbrANTGHx5ZM5okF7TTOv9TVNW05/qotiKItuZ
nBSoDGj825q8ssQ2JFWs+zJX8+PIYsIjFcSzSGqP/vCXfPFMspfXPUBQAXlJ6m/o
zNODS6hce6sHAvw5GayhBOYt9av5joid1bkLb/Inb3PxKf/nUS+OTa/FnDbH5c1J
ljVkV116U494YLCtWC+RcE8eHtTri6m0MRew7w2dAFc0Re6bkAK02nlU22U3boqR
fvpZluRcu9xsctMl8e/m3nDtzopHWk2Q2xSH4Jpum6gMle0j02nQ5GTmv188KLme
yMf+8ztYlE0Ov+VCbhHTNI9mcY+LHqXR7jc+WyHGZG0UVoan0FXf/ztVmAY1kUZG
9GapjCj0tFJ6KiXf767iLof5Zqx34gBusRVxZZR2l4MNNPI3bb1eRXZydzFD19r3
as79UUTJUS4XdUUk/L+ALfO/2/0trUVYGBgmRzC+bTJ+wtDyZXjyhbDRTjQj+Q9e
ZKQmDZw0iJwChLv8AYiuKbGXeWBOXhkqTIBt4H4DU1vHAYX5Mzwb4k2N4ySY8ZA2
8vKZZBXAZwyORYIWp9R/nkM6YxLCGpD6HlTrX289zeKPHWM2XcNwvE+jmU63OItn
GeIel5CrZ1LJStGNUo/hndZBdddBmpTxpr40InuyiflyDoymKfYDCYoKYFtj81Uo
dgjXS7OahTmzum4JrZqlXRDwDCogohNtXb73WYU1p6f5wBTK0GGfVHyir3fBX64Q
I6bgiJaK14tMfCAtxSd+khlyuhwmp+dKH3Kp/SzAYmPCuawBWCK1w7dDaJ9IYD/u
sLvTyT7ps2p8+E0R4d4q7jO2apm9s636aQdFlyfavt7GFe8yrCbLEoJO5+QHCRFZ
XeKPN5ct3abrKSzmM1EUjyRPZRIBh7J45U7zFemEvT7Ac/3/jRlKeDIq4Zuq3Vaa
Ydu0QteAN6+11JLbITl+sWZUkl1HmYLyQvY6MM8XqMCkKSm8rCXO7rNgni3BGu6O
2EUJWba/4aYJR/cVErjxk829wy7qKRoIq8Rx/3D1G6S1ZLBlSt87AF2HeGU4c5P6
gwFbtDOxPhNecqzypo3k5GU/MWxGNOp2Xxtj3teMAMfzbPUXRjVObhh5seBd63Ao
BnOYlm+TQI4F2LGvRPgHGsIutlJFsYgzhKWCCMBEWv/BgiHLlaLWE7adHLdCQ6QM
k1HjCDpdvSU0BZZaFf1++CPRSVc0JkFvPy/eAglUixUg2adXGXYtSjnVElVHFQbp
5tob4vSi2HbyZcZQg9xaEVgZSEQsH2jaQLfvLpjqqV16lvRj9u7Z9GaStQaFMuW/
pD29iUJEk28o5Slw99ygnVYt5sfIgF896774vKOJITFAtTmabV/0XPwl6SCOzE6C
e1qhSqN5n1ekMRWiKDXkA5Km4wScnInwMBuL8fq+rhdhc+v8Y0PLkrxS8zuP1jph
SKyfokcZ/RybImIdFTWYgdy6GkH/g8ez1T7KRNFCR8QQSEx6ItUJHkG6SMLygLSY
to4aygDLmKHTEK7kdg/siASpP9sSpVlDnCaAOphqHLUKRSYCS8U5m8+bx9UeEeST
vQtaxlsw8ifVO0mtpymQI7+0E8jMrQ8Vbx1Zk9C72cQx5AQuu4SqylfXmiKdJ+KV
YGU33UEjPgQycPsa2ciEbzaqnHtnPp5u/6XITz6TbTE3rGihkChFnoo46r622BFa
u9jRSXWyAHL5qCy4+ZbPhkXQ+WXN+IGUjyYqt4HX0UyE/k+wFKD4nhU20rk6LTNE
x+FTblTfVYzG8IkBl3WCVxhKyurG7u/O4yCmFr6YbeKSpV2+YA6FqvKEtlGZ+Rbt
goxBPwrjUJE04tJh7ah9xp8GvyltQshbJWIZb+30VdKJoc3LZmHgWWrEny+IWO+0
GcLN7IOLf5P3SUuFwB7IcfqSRHea8CEumWfoPXSgHYL70API8rtxOrqhPCEJFmxT
EyzFWnjro9e2cJDz2yYLQC3V0LCZG0B9yjjTZBEK5SY1IIx4Y+a4Qct+3wyUsbxH
D26D2wAlkzOuakImqn/UnYv8SW/Hh4FwI/MDKUBafOF7ftP+dU7VwxrhSVda9oZl
Qb2pCffJLxHmTE3165KZi64jKDajv3VwKs0o/BCYevlmhkLgO4NFdxiL1PSqUD1J
AP2ZX5MCwc5sVowHRRc92Jq7bZ7lH+PmOEomDvDSc1Zyz1ISDDQG2aC1Y++xNC8A
QePJXkc7NclrNlhaKVU6uHBXI0ljW4dnPal3KJeLZDD9wCwrL6leep1FqG5fUJhQ
soOy3JQqhkWHOjiS9LD+A8yCoco2r/hh2EnnNfbKPgsHBEQrxJlxuSwfWPkFmuOr
yrPzU3QHURS+ikHd1SPdymJSzD1BX1YOq0SyYCz5NQUTcitjA9EDFspRzsIoRACl
0x9sI9OZeAwgdhnG36rYnsEygqxltA7NxQHiopFK0ruzjGe3q+dYUP/1xx13u7jj
ShyRJC5DTqeiyGvun8Z1uMgMtxL0+9e2N//eu/WXCk/wPoS1fX5DtCGsCy6P425S
ZC7bkaYKqt+asd09FiJdbfcS6G+N9daPPa/sLH5ljs6gSoPvElIzFnM0XWLI84u1
y9sqZaTNNq3AAW7Jx05qFpXhheqFzt9NMx7WuzLSiCBLga0vly877h0BsJYKKuY6
+BsgaRsLwczWmnFc+lv4j+zSPBCkVGyO0O7u4mgvQUxWVijGSJfnhQC7TpmphQhS
YkyjgAXu+B6ZlgM3X9yIlPGQmk5bSWABS5gpAfpECisy2JK09a+DyVMSkzZPgCB/
glJW2LT4pCUAxwGgahg30onDs953gBL8FYqJ+Vzf13OMxsatKM4a0/nyBQa8eM0N
NeJlz0XpTfEO2XYKSHMlcVhUo2gTzcS0OrQXdcF63Asjlh4w8z/xDqhZi8HczTPz
/IYv4VGc3dLhDGcRd6a6hlZwjgSZWzBA6dPeK3Kues/nNhjumumSrHwuUgcUPMBp
BK/lYSDrhWZ7mFeleyLWqa27Fx8unaU3w8Y9z/h8hrann5HmIvPLVGn7CD8Ky7FQ
RNmjT0IxpSAV05iMfqUKLB8gcpwhufR1ijWRirv1Aa//LjV/uem6o11+bd04PKRD
FMdsxXM67XODS41xw3wcwFHP+1tksJMsTe3ikEBEYJKYohX/366jbcXNHAzZ4wdR
Bz9GdDy7v6Q24Xt8+DlYZObo3AjaTt3PVnypDC+DcKkkUKRkZ9XH5VAa4WCcLSIl
3BaUCgp4Ur26mXuWu9eSRGYCe5WmW7+EzZBc1z8AAbYRNI/l1GOyWpZ5634m0e8r
64XbTgfxy9iAvcGaptAYvVdlkf1eIOZCYkGjtBqi6itFJN39fGXa3mKzf4zb42Bl
H2ht6/+2YEb5FcBJRv/OSXJsWlWJoR9HCCMC15oIrKRkaEzz1AwaC+ofxpCTgggX
xkiRuU0NjVDqI3ivwsCA9lvZdK6dCX9h4pgGUM3ox3dEBrdlfl5t/zIopNuie5ri
meCntIs+Te3HQFsgJtH28B0xobcwpgoHONIu9DK0KfgyMiVwepHd6ZSpM8UvZ+1G
RFZcZ0m7zrNiKlBY8WiKLTDAxHVeoEchBKCxbiFmvAmQMjQ2dRDsZpPfclQG7TtX
+ryNTxj0vuVfwSrWgyySyvmdh4qlbDzHBeg9S3dls58GbOl7u5BEZKkHVMQ7q8WG
0X8uzdHnHwR4KLx+MIas4wiCo9X96zN5hYKMxYHTev5oz9orhC3XqR59itzE6rMT
RU/ltEmwwKmc2HbnuijBye05ZDFRu2GqWFyw/K1RQslm+NUTCZsR26z/rcJUnxpZ
ZKpITJrcrs5C2iJmPZfX8TgUd0Z3cS5bKAlSfHmGSnTSSFRRVevhi+V+Pdah2TvQ
Rp/GXl2WpnHNMPbTvvUqPeussB50j+U3hZvER+bW900rGGS39qO/3bzgN0Pza0Hn
rnMARH48tb/RQar/Wh/Atf5Hj/c01jIMowsqsK9d7MX3/NfeGYDrQ4A+arULK8Sj
TCFFEhI/ilSjF+1IfND+v70WZAAQReiKr+hvDZl1KvmjcDMeKIq0BRTbrIVCXmEp
xrFoYHalmtHjAOQnOP70fGD6zRR1jTpyVfP/fHP7Ujkm19KHCYBl/jY/fZcJcEz6
dTeR3Zhm0j4AmJ3BQBVPzRESC87UdiqY1N0t2P2izgtDMYWHeCwLgA45ep5jEW0n
rX4kbsxgngNh75y8vBTHW84adfkBNBXM/l3qTYtoIqbjTrBewBCI4WSqJ99kaA3J
4hJ3vI05pFi7Co2OkK20nuge75/5W0Oq0FDKhP2gxN6PtGtshzsh+GC6MZeM9URK
M2QESb00SUO+jEXQdA1fTfqNKxp2Y8Ynm0bbWglsEqVXL4MtwK9y5QAPpox6YQAZ
t6i2cIIN4lXtrE3H7mxTEr7P0AQDIjKWIMSLQLiqHoktuCe57hLItmJv3e3WivEN
MKC4B16uPTF/QfasgnmPjA9e+c3crJd1nytB1oG8kl6oCVn+89Gjllyrf7BgXvmW
F5RIShNJFQTzlv4KT2bjXui7rf+ElKd/6l24aUAYHBzeNc9EuDNtCLLCLL5ER8bT
q59Qv1OjkufoNL1NA0EavSv94thIexmIvOzly3rqKb638rBDHMEQlvLkxspSI0JC
Nxw7qeWE9TsPQLiKUPxQ9XvPcg0iWmxAoAZXTnwD+9GUhgRfVyr0GEaUIpVaO+9l
KsdAXvSG1syw4QXiOV61ZnvzhHOOrkEAJjJvqvtKB7Ib/TuOBL4yvQ8ZMxqxrQoJ
ZQe2FvMs7lNQV34/oSPrY96ziAW2xZb9Jz80XhTpekUnUMJp7oc4t4qiYf11IDdp
APQ/jdyhkQ4xPtYb5fKmPERPtsdVQFcrKDf443Vv1+LLcL3wWJkir0og82rz/Q+u
VfbnejQczuxjGPJE6kUOOGWcr6bLTemZOBJEQ91tl7Ouaq7GRRlrYlC6I7xLNZZ8
DlByTOIDCAhlX34SCCVc1Ip57aQKsoHANwhxbKsz0y+BeZVV0P9YNA+63a/5cgXv
SjNShlMMcY7D65xr72VC2wCR7kAnrogI8BuvITYgEBSCsr2jT0WjGTu2/aFblOfQ
ckBP9bxiYrQGPOLFBtTi1uP2Ju/TixXFla0dJTlkM3TXBxFf9/fQ9UzV/j6IxnZp
3Vp5g+uGJW7NbGpkPqnyYejZ+D/Z/G3Cd9ekzTSdX1pOpWbtkFct0x7NDAO840vi
An89P+pUlkui38GnB+xq1HOoWbiYm0aEeAsq+XNsJP1KERVV72Rc0SHRPzTMXSb7
nk/f6IHeb21/hmRULMbrRA0duMST0YDC4XMjntsuUD3f+xJiWclCkmUDgOTlIW2Q
+6E7/WKRty2ratstgoS0GTa+EwfvxXHAOZpXLiLv0CRaWpCBH4x2lvV9MjF+z7id
0Ft+YIUyPL/kXAU+nC/UJBfLQtHAofgPnfU+E+FauzHT1AamqBM8491pDztbW1VX
Ra+ZbcQbQSetxEAFdkUvIT09ExaOFQ4hQr12435AgHEj617rSj5z8RR1FLcLgUxc
lvGJ6JZ4pSGIMNguaeHqwbusJXYfCQWXgVOAaCpPZD7zt/dWoNiIbZor19ZB6UDX
P0FDDnpSQRwUcpsrEeRtor5pAXoyIWxFjo0m3gXnTc40y+n2HbP4WWyrIZRxAzl1
b/gdl4TInmengQ4DvVmx2vWvaj/nT2yaCggjy8j7KBQ8B+Mx8WymDZ4tWs1qBu/D
EHknlS5I8FLI3xAEkDoPm+1cqC9cI7zfV0xlPu4R7vl+4iPQFothEMTENKMvu/yH
QcaBzTQg04ZGPiCeUJR/l9SF9MCT+8iZvYiEDQjEGhQCGEp1PZ7jr5yN2WAjZ3wd
d1IrSKCxu8gJbTmwN4Rmbxr1Ki59wH0F9jBAOJCKBqsYbGEmIBM5j5HCRmoszMCf
FNpQHarMQX+r+mHTsv5oG8y75tuEjT19HEbSmNAhY9JMvD+ycO1MFULpz60i9POX
OB2uRbIQ6wFYLuT0UmivUub13PKmdpjLOaCLw6+Lz5USbCfPSqJI/sGI7VfBSNEJ
WQzXx1da+9IBS2v1LUGYJTGo2qq+aPgJBo2KWyzYngKy+nZkfczO9PVM5JinXxmO
jUY79rRAfq0MSbkKjAyvP4u2kbrNpQPdM6jtGmbnjy/fzaXi+JqvvFPUPPc2i99V
stTYHh2L4vIolImVAHjOJmCLwM6uYQceQBrCjpnSSh3FlqRMSWE/3KUOGRwve9/c
pkETGxxE4Dr6YP0F0Gk8OEVQ3mBR/0NJCc3rWeWUz9Dtg+OG/gSvgfUHwB0Mh0Qc
OqrD1bxqmjzMq7AfzBdGNZWcI3JBx6I9aj7sg3I7K43gdnk2UjE0QKANk9FUmR26
QcrBA2gfrTAVTjcK3A4onJ8CC6ELoAIqYDw2Ug0neIqm74Mu447yTDfPuFgkM2ah
oMP0wqcbakQTSBW5kZqMt/zC1rbtAGhFxmtThStQtqaEX+298/rYa9j+gTpTrwvi
gVX1YL5Nkqjo7LnwegWxtH9cou/98ijCQZqCQZrdWEBhm6DGIIRV9h4fwlLeWut9
O9pQECFpRVRyE4KJYElSx+r1drNKiOyowlc7D/tyBhywrF1CGuGCLWYS0scrvVR4
vCHkqbtukdg3oxJ2LmKyMkzi6s1IoZv91z7H/6eHu87zjuufnal83QDTw8fIkjhz
qxeqh6zXoRQQvtJxTI4LWTWC725ipzay3FGKWoN+iacgxXyyuiUv4NtiS/FRIBU2
Wp/wx5NByb2C67FiVylAnNfk9x/VS8ImJt3NcoJV50TfLSajTA9hreFC230yjzG4
a6+yMxOunR4jy+nYYo0Q+9uvXMU6UuWELY/wUpM0uTYxS3gH+aED0Q6DWMojO6sz
sVCmAchW7jT9177aAB45iGP9mpOh4qDB6x7m7yFEDGs9OCN5T9hLv8pmsaRMQFv3
F3Woa18rjCPNh25950LVVtZCq3bhDxvabsoGXu6P34QxNxya3rgqpD8lgLTx+rL9
ij5bIUUFUf4dD+y8oxuw5Qb2E1HZXvJCsR86qZDDUgNvSreVYXrstwAs0UhfdOer
Q+U6i405B+6vSGLXQLU6Px4t2+dSWSI125PfATkU6kypJtj5ZKKTApDYFTKWKNRl
SwVO1fpoFkLg9ta+Y2h7tpBP0gjYcSOk4+bfd9HpLxKnLWS2JQkZwL24pX71hGSB
gbuL9T3nCKZvRtBb3hr1gjDPBk9AprB5fAv7Kq3nFCCFzgLY8FlSdpOW5sYolnmQ
al5xRgyWxfkspMCLP+nZl6//C75tCBHFXvkdsXWyUpnAW51M6n41kBSnjYUM/0En
Rt9q47ndOPvjhejsPi00XnsZ2ya9mL+ZMFuTx0+myTik4kUEeBxHM7W/NBeCW9cR
UgJalTTNPB9iq4VSxq/D0nvmKrJVKKA+bvkHTO86lSo6aIoU/XE7myRzx/gSK+Ka
I2g/g+hF+G0+T1aVqV3TYzF7K/pwYoq7eLOmjgT/F+lcXSn7y8ijDtkGNJfinOH/
KnCqUpeP37OrXOH27LVv9RVe9iCoQ350QNPq9a4q4HXu3KuocnNXN7pB72M16uUo
khp54zQTFFOuRT0mxlkR6zL6679lbrS/OiyyTrEN5pLpg2fhZg/ZiRNq+br4JO8r
dAYfptxKuAjVHGw1oa33MbwynhBN7WligpTU3FsXdtgmgWP4VOK6fX1eNZAR1rp6
ckUYTmVTuwf3FUW/HhJWdQVRzxx3fhVnfaXxU8VlKQ5lOQVDMZmreWEF6DG5iqdV
P+98hUtSH2BwJc+OYxRpV4/G1KGMrztex8ykCNcKZ3u6p8pfr4ToYM+dvV/TdWIe
n/T9pOiDyOd1lmi3rRMKGeasI0pJc6J0ZjFBfBMiq1+hlCmsnPK/Q9uzunsI2hJc
EugZoSReLKmDtJXHunNgzDHmaUBnnd7ThiJw9DKjpOMynOY3Z5tKPzXGUUDapP9j
aHski2xRXh26poexhPzngKSWR0inCtrEJL6C149hq9qFWZnAuqZVQATN+OO366is
jXZ14PcYtAjNknX/0ixHnU9Nf/mjt7dzvnyLBrhUCeWvYstTY043O/tO7M048OfB
7JQHDVVCnbyEfmbL+JLLUsYVGKZ9+ew7dLd8Pii+ozMAhIIUuON1Cn5wXBWefscg
w11V74z0XZqtu3KFLOrkBUEFuhwrfMS8OpxpneZktUaCRS/fOFPsEKHFO50YMeTJ
zDClPPWeEi4M0Z6FVOl2EQrhTgxO6jSxckQvqhdwAi5JDuycbVprP+gsb5zbCXzb
+axJJcNY3pbgJVkw8WI+nBGcbxy8u7gxuarAxrttrMR4xXAhwgwZKuA1IHLsqXj1
mprGtKMG5Jghw1nNM2kUj/TtS7g2w9+SVBn7MoKiojbrZXE30QLz+66OJsQ1H99V
GBHUHa8xDJYaJJ7wswx6Ms2Rza/Y6m05Lyv4WKjXV86OJQchGBjQ9XiV05QIRY9l
7TaQ4OtCGe3PzyYXVA4pWQAI08lAOeswgT5bhZIQHlvDLnZBAbKCdjMrREG4ZRZv
Y+oOxPhBr4529iggFrFrK1gtCVKS3XOim3bqVUJkD/fnCFVR6sQxkH0Pk/BuIeWW
Jm2zTePdLQmlta+Ec5lGtD7x4KDRnv03f/3gYKe3R2ZqW6lknyZE18nbUqOI0L3R
sbXWKvgv9ynUf8O0zbx7WNlv8MBt5k+AuBJ0zJKMFw38H8KT9lmX/Mbje3Q5w1+I
D0nTvyFp5t4NQlUqPUgtIRr2KKWvcvelPu3afWanRYIDLO4ZyR+cuj2z8QD9iRhd
8f81OdqqMsOrKMgK54fiZg96kF+pbWIY07IaRoLb6Jt32x0CwRaoFMF0QTzuw8l8
JWMYqKJUCp/eM0Hs10b6121EVIV0xr/cwd2DMuAFSNhvqr2ZUANi61w9SHIiCGIT
kFkl3dW37yHDUPeorDb+WTI6H9FiyoBTgBTzuYmDmpF11iHfNkhuOETRn1MGwXYc
uP9FPz/++0T6egVvO2BNM3sALcJ1lDpvGG1dQudsa39A3BJa1Rb/nmbaeGfgGoo4
pSce6xtq0ril9puPDIi1uWhR4Fh01cebkoNtJTOgA8RAJsEbnS4R58JRY9C1zlCt
YC0oKSIggeEeNH3gxXY2v4w3E+PlO9EJgurqXCGHhks76kbbbkEru63rpDEJkdbt
sFwU7IVUIEY8jHrKfgnasm7r1vqxRsDU9JyJ72Prn7sGdTkRVDS+lWeByoHgoVVj
5I2K6MbpW51AXJhW27TCzxtt0JFq69f20jnpGds/C/0JLXFtQIBcdMpEnrSW2V+W
nBa7LA560GYhtcVlzKdo7gPpyw9yjJdm/Uj5Zjs5mBXk7BQQs0FMbXhbOOdNX7e1
GeyMaE/ban+eccZE51wcv9HRNwwS0PXpKGfBviuX/29L5HGVZMuVFqmVFh/hDAXN
f3TaQJ7xi3iPBO7w26CHjp44ZO6+zbVF6Bd/Qys3fn0oHbLnt/G50RHEC/dHLnHz
vu1qrfbs8qNobvV/ff4lX0nyHoTtTwwQeX9xXhu6PC7/tYY/LVvj/ccQ3PHFSNjF
tYOS5pPvTsn9KhknUWxhb1N+UUorCexZqwi3rMRAzgUqVYObITlgkjdYiHLRUZXY
kMKcvJruQgGjsqJ3aDO5rDtFzatR2fFNCAbukxSw1bz+iMmkTzV8QGSW+BA9CAb7
Jvodi2YCsb6QV/U5069Y/O3iIoLx0vp6jX/K8hE3Jtlnr4WrTF1v6Ze/yEs8WjBo
5dAX0vB6r1R3vC6X2EBG1SRuTx7Eta6raDmIosaudJb7npWfKdS/ztnY4GVzolS9
MFl6EeBLP1h44EQOUWuikul/ZqvRd8y/vwdZaQhPebi6yygklfEFf455CytWWiHa
aFJHflMWY3Waot10ueI2xVGsXQ02Nyz/KWOEDi8KfDnxzWWWhXaqRNn5hgkz1ZLM
mOf6frS8VOQMMiwu0O1+Py0wcXxysx3aBHzXEeZ5U5asTRMbp+ILFdJN0Q3uAAVf
rEL0Xa8+NKtP1HxpANyMo4ROonuAPyLXfUjJxGBNJd5QHphsvXOJP4tVTjsEmXeL
QT6BZoTbMZwN4sW82p2vAscvopngw8zCy12afcLHdC0Ce51hY3PHEODUzM+VhYOl
L8vQBRNXd4NqYVBXkzfW/gfV+3U5euAK5GlHGw+W0RKSfjTbJnoVafFv6mYDPeIt
rkOqkDFXpUvqyHNzAH/yAZDl45PfRBFGosEfowdXVoBiIQz3ZLNzRCWnGR5ZGseN
hbQ6jplIGIeKx9F4XPzIAFch2Q3aFdhgVkYEqYdT1oZEcJap9jh7q8LqRWrGL2aD
HRzK7U59QVRF4nKL8V7TTYYkO9gwq5D7QqlHi1XYte9z/bp3tMyGjCeH7NgKZ1WI
6uMBpfS9AWi0lxMrfTwW0STotWVVyjLoZzCxQXSH8+YoSRC+SrwgnI6g65uEuEUT
/TRubMH+HbjnTn96raY7ebz6maXkZML6Y+DaRLLmpCMJWzO0iOCPyeE7HaUu2y3G
+2W97v/o363tthV7dZLcpzyl6bGy1oWD9LtNjEWsq85OXcukl26dh0DQBMQhS6R7
EfjkkSgE5aNp/RfabEZ27VgiLoi+qtpri5xvgYquT5acNjNzI06Q19/nBMXM6nAh
4+57KVZU89DlznD8qkINvUXIv4icpLmD9pLYyfSJoHeuTZZ5yc6K+sI7/druZdwo
E3YbjAoWTljl+BS5OfVTKVbo5/+vijuzjdj7iB/ZTyjj0wHebssJHyNIFiKBMvBs
QBIOmKeIqidVnF5Jrv68P2KFB/DiH19SioSLbp4SNZ4XCL3AShzKwf91OraTJrxP
zYner7gzKnY5BV4pVjbv+LxZGIOh8D7/LreDWaJNVTbrYuOGwgZDnHGVPMrZWR0f
eYcNdcxbNvTVW2gxghKlPbHUl0ZP/TKCjRSux5fgCpEzc3ZIBYGt3MEDm+8Z7biO
PrEL2TV0iR6RcsUzA73lqWLPLo4Vc/4NFDp0brC6t2+yEt8Lp2xM70Jz/1Z0prbv
qlvrSpaJISIwS1pO7ZZSqTlOFhkn/Zyqs+QMyv+KhWTOzqJQ1RuOXEN8PCRSEF6V
llA867KwcCgcJ3XY6kalUcui9pNkLARSU7dCl4sunlOrAxB/9qI8Pk+eMpOPBFbL
eZZBy5viG3E0Qgys3A1iq11Wi+pQZrj2nUdldpLDX9TtbytFZBrK5ObiDjnMwJyp
1uGV6jSR/KdlEwySGSlTy6TQsrFCpqzRhXb2aZjJ/z4UfsJYb7XbbgS7gbp4TjQw
iZUQ6sNEx8Y7wci5EllSHiHHOZflD7N4tszG6OXemU2GeI27D+X/GybbPagX6OX5
mhVa5mbxDif4+oKk572PDg6i/OViBWtx+SeIcZg7ybEhkzQbQXmEmZxH0/4TlSfz
A14WZK+ZO8VHvuG2lhrc6/Nvm+zz964HaZXAY+9ROKdEsl3ABBw61T5v81CRbe0F
/CMh9B6TXoVmdF4kbWUfvx3yYTx2n3OG74uVPDCmBzI4iDLtMJkv+tYyAGqWgOiQ
ZBwqTv2eMuSxGpm44ki6Z3ycbeLNH8pw1rMl6zN0JCKN2poc2qIXdTrkjdNJugtq
CQJAQl1I0XkL82ppCyaq9t6HrTXMEWVjDquOtS3dBXR+e/2uB6/fWBjl2arFyE5r
RskEszWSq6vQJASYt8HS+YbfEchrTpCmHL/NSOg1GcoRpcLN8xDX+rSL9ybb85HV
K4rp7e0zD5RCZEBrYOrZEKRCvkjPOdfzCqh+lkn2ykK0HiO2J8xpgv8o5WaLK5HG
GfMqp40g9Co8vZQ7JS8GPA3W5UeNZPWdYSzfKjod+NoC738HXfgv1c1TQ3t1ec9S
FCjRjOr/vnrCMSY2RMtK8OZNwaKGxUGi6eOtPQYEXso1OVOElTjDr2NlT31zDD4f
/WNWlrt8k0ap9AZmcXt4JfR1SUhOlPtDsWAm7HpNWq6EpTZXRtzxZ8UQ1kZFduz/
v1fvcRFRgnAXM0Wgd3XFPhRt9dfcpRw9JP3715zJ1SCmRXEybVDbNteqHK9HvxTI
elD3oUS0+uPl41p+KeSxJ1SaICBC/iSTIz/DnBvXgzYR3DHhKXZ+pq+EYcpPL4Pp
y+BlzqX3CsYiiJ1//3zeE8C9KpBSOuPo14+o2M/jkikNIGawTc5gTt6CAW/g4feM
rz2XD1sGLDB2eunzCv+VpjgUaobK4iLXVNJiQNM1qmHMiqkNIReNk00KLMS+QAKp
CZQN6CNX0bK7ucTEVpRyJVuai8QinQeaO7D/hyylDB8Yww4OKCrrBnaU3zsn8Sij
VfBHgcmgPeyYYN2VBsv4PtCh8x3WBNkOVeUJy1DGR8N1dwxV6Mz3jtYPkIvwf3aN
k0V6QNdBq0WYwoym3nVTnAehxP+ArUEz4I+5txY17GrWTnp/CpHCkXEkfL33JgQC
ssXQxk89/UPzmkaL+PQ67lLh+t0P53L5DFTudiztuw4SkooDHYuZPaS6nNmoeT3R
jyNEUsU65+HhsCUqWvQTjw+y2JuK4QjpxSrrLG6LATNIMig+ZVXEiVjbUnd5C0Zz
Sbv7tsC5xnUG1FWadhIp7/6vUAvKg+0mPm5URv2eAcjJMdL1P65Xzu5lVSdTS+Uw
/Ak6SXb1jlsl8YAnwPkOEkExw9d9rYlDZMj0QA14HSV+4XCS3hs+qXkZeeXEIPzV
+5VYEQK5TogZjQSnQISuZ9TrEgUkJCA/T/DiJRAd6S6Myr6XA3Ykar+kSIgU6lF7
jA+YjP2X25PTSvoOs68bFc1UJq2+/z9lNGgn1bS0A3XpzlmeHAvPi7NNuNdrecsF
OBS1nLE7qwgf5EZvki+6RN6IkTJhSmSpvw8R7RSz8gk2qKtZRaA4fNYQ4MkpkCNe
2JE2Z0rmu6eN6K6+/pB4pH6O1nSRYWK4aJMDV5IMjEfLLtzwOPty2GZ5Jx+aZ9Eg
oYrC2VLkIc4Mbc5FH/ZeDJvYQBVAl/IOfaNgZg+3VRRT8exlcs+X23ia5yCGnvJf
cBwvhApORQOb1l16f555dQqCYp1NJ8cse1V/iFNZEzIzUFMTRRfGE53u2hM4scrX
z/IJ44eaei+LSR3HcRW+wx33t6lhCzCoTXpRbj/ofioj+aeYde1ECaJqNI4CB3eZ
xb1yfEXosEcwlju/FDaOkS3abzH84OlLOM/kVfmYWs9hIvUofmKmqp6K8TfuV8dF
x/Wxxpvr91GmszhhGsyAmPo0UkRCjwIYDYbM5VDjCxL3oo+4KMUe+w1KCEqNZMeR
HZ744x/jt6nP2F0POd8ofGaWRSHMqS1vAG6ddQqKzX0mRhYQUOkI3Jgw6r1/+C8V
JOGzDdRt2S4Xgk0pI3dneOj72gDXUHWwnfXsNyVOzEaYAErEvFX1M/N28bIJHQZu
IwSbuK2qjVr1ytJ2nJp+PbR1lahzPz65ippEYbhHEi71eGNVbZSrEWojR03bmBRN
PcVMkiHyW2VlKr9pcQSITNRyx71b3p6eGTpx101NilrfkTo9tqtKuythiEI89jZb
o/yxl5aKv8d5Y/qpCA0F9b4gVvshLD2ByuAbGmlw7gToWXuRCEYYlVm4dHJB+dbt
kmV8/7nQaSmkvtqTcku1GSAzRTHlJrVRFBQ32gWAqEbx1Prm4HLLLw9Ik/OeO0sn
NagiAggJg1Jv/bF7+0FZoLZ/9PzBOWrhe1egAQALWJctGrIxxd/f98k6eZJd3UdB
O56NtIu2du1s13S7/fVkU5P4YMzGoSG+jAaLnXojspxb8zVMye/UxjzrmfS6J/Wj
0STChchS6Iv1BTuPna+uyzJHJRfoXHFTJDysq+JJqVVjYMuj6OlQLtqBWe4MKtPK
7d/fGR8Cfb18ULbOGB5bbYpvZ+xQLl0DepbdygsQGhCZT9Ytft6Xr6d7Rk1uzVkX
DYydjc8LfhRoSiEbneECjQluJJKWdQgzu8FtFwV8AbDpL/hqm73XiVIqzvSsA25U
QRpnpwuiVZ5o1IodvvSr6o6gi3wqI2lvliKz95hUNmJmJcsKAXF1ohtg3mz5BFea
lKrAPMcqoGKPFxh2fKXvuhtDshmG0yaEglJILuLcdQRgYSQM+Btq9QmmR+QNfOLf
sDGGR/c+b/4OoOXCcFLzU2TFDqkowuYLG9a4ZExeWl3s/o7IgGQmsPFIQoI7/H6Z
EWBTRAfm6Ul2QYkH8yOO2T/KGdkdAxbTqqWuHaHi5KqsGw463CCmiEUhgUEQSKlY
6iNS9dWkaW1LKS2NhW9up64/Xd+XmhpCJhjKq5/XyGG6hvj72NrTzDILe2n5oi78
KWAlPVt48SUt90IPaoQiGfJyLKNWPrszqM2FUMCg8/RyZaG1vQ9FFne7fRB+ScgB
WpPOexA+Vx8PvcDKFOg4vx+GGjEFb9HcOZ2+VimkN9EnrOcCNiBDlXIxRklNFClC
vhd7HXRO5wbUPU0Kyv9JgVdsWI4sXKd6PyZpuQAKEVT8adj4DkU3J2xqea3gTsrz
+Yu8oXqxpRqpFSi6nO+8rZ4EqkOktEvDscCJiQbKN0UvM/A7OsA94rO2bX/kyqW2
AlLwpujvUf27ZOyeGzFFU+7r7O8Jpcm5QRuC8Tc3vnlNabO7tuuoQc2TJhppDxkg
XPOxdeijvr0EY222Q8ef/5556BH7+qVMQM/T/zCIL50ml7j7lshGDGm0ZW314j9Y
6VVNW73VdNfzOJEqfYNY9gNhoWPHB18k2r7/75SjFP6A9bC7ps2BRcL5W1rQXnk1
N+RpCIaS47X+EtZvs/HW33bF4QwmzxA5/48JNJ2jkzNW4Tjk65hAQgonFelEjUP4
Y7jP+PJJvusAfm6PpzlYx4GDXtVGbFn5F9bsPtqEt1pdop51QaKJGN09IZT2EvAA
2VC/JcSqEQBqsWv5Z/lpniN64JCrzwiLOtWBU43Z2v0Dfch1XnjalAEP6ySRz5Ek
Nebgp+d/jI1zzfa1OjJVxR1kDXuTboErT1Zm4KRErhf/c+8fEty+KJ6cNhmuP+36
X8qo57wC+oyCh/VRG8c4Y0wGrubUcP6mEQXoOD2Gqv5EgeR4O7pSRVwjhDsK7XwV
eYmBj6SM7E1R6YhUwfxulQ7YR055bXuRl11xRh4QA2p/CH8ynZ0+GTwyt8frbUMb
UmnQlivmuPRlEkwiSYZXhvMUcWFd0sOC9wtxKMOGhvc/Pmv7VcJWfEmpedDSBjta
B/k5chesGFM3yOLzGIz5Y0R5y9G6LJMpZ56z5vHW56FYHabKumX/OGRUcfXk2yTQ
jDtiVbCUXU2J8oVeMdhvKUcRkYL5EbjZxVBL5OLaw/Y26EkNHAefcWGyh79n1Nqd
/onD+FpchGC9LzV6c2OLtnMcveetB3rJXuFIGaf8cVuJ6Z/dVqgYiwPbIiQ+xq3t
MWysqbVOCdCPK8d6o2mfy5ohCI71BvrLnc9SI5Z0nq9Ke5av5xmbD94e106RUGBB
Eb1vhLGSSMNZVpl//eKjEAgbOJ4Os+uOJb5n9oi9pGEJFSRsxcH2RiAP3+c8Jbxl
L0VB3ofz47eltqgJ1loNRh4HvG2S9XwgxomW4R9VoV4VdwzmJmiIg+YbmaulGPlP
TN3/8bBWAS3aZA5iBL2xLOB1aj0ehnSriyYEWrfvVLcA6pTID59bknB3MIdBqsFw
6/daXjZR7TAh1zjzEOKUr5wecSYssdKJULO344OBESoAteaZEc4b1jKhNRMxjBTs
tRcaz6KSC+0Pqc7IXUZa8/S4n/V8srGAFpiwwbm9T3CTIsDrxbJdORO7cIfgxjyu
o2fQjln5WCSoMlkedyMCXFy2OxQmqcFh0Ep/+p166huFyOdg0hNxZw142RcXMCJd
WblEcqsU19lM+AsRJDAMa83ck95E048BmHtUFphOS0v2ct95icBegaICzJ3mHuwj
uqX+7leDSo5FbSHfRDqLrYlpXTZjvuUOjeF4lwTsMD2ftYmrtuTZzJxlNu2A95Yw
WL0uUptEUkd56J4BMlW+Yq28VwFMSSEjj1YLY9FFXMoaBIBbibmzUDKXYx957yLG
URjnVM48i+Is3BHcu/Yv8STCnLbdnuevLu2nlznTJiULQKccz6mcd7cKKoiblQuA
4oGFszneDDytDrkhr3OEo+2r8nbZ6qZDN3yc0Mfls9mZ4dRBf219TzTLKWYj/+Cy
C82gZ7bMvyGAw1SOCS+ZpneQybvW7OQxqdjckoR8fhP5jVq00Hamrqyx0iAIPVN5
gpHFgZlX611XbvDW6ZwaQyEltZKDy+W3DNk+qhUOUghF/hBego0olOAO/OGsAmRj
oZAQ2UXCphmJUceBe7TrrL1u+Vloip8xG/qyN3S4kVV22hV+qKj2q23+iMnqQv4q
ILT+Aq5R84ntZwDU4YBngpkGvgDPOyXxN4yEbqoaciDvgUFZLNbj0N9icztJ+hJ3
FLtmg9eeZUT+1+LyTcL/OlyanFN+dkMxfWlgKaMaaWJYR/D0uTTiG7EYkTvjdMup
46Y0ZMw2VE6BtKXW8DVf4M30Pi3tSs0ngdIOz5RWg1S8XabnFPfGPepO3TqSCkWK
XsLxA22f6VaPO07V+OXn8wPO891lYNRr4uKoSQP9Q4L46riRgFQNrubTVaPEBMkg
jatbLOXtq8Sz+gLJ6alZFdl1WeblMhrCRVkH90oAIeEvUpjmvQfYbI/T+0s7fcb8
zsAGxTo6MYhq40Sk7xqfmY16mEYMLnD+BWcMYybS9hXALPfWbbOlppg0rfF8lYaz
quoyFB7dCZDXh5MzKr1jlR6co0tU4PhvmqXaElR0/gPYql8ncJ1hB91HFtWRTnv5
5NNnZ8KXrunEb94S7vFFQZHamilZPZsMxAu21K/J/Hzgw0TgaZWTvR+EVKg0K6Oy
RvBZqsr0FvLnEXeIY1qngGgc5RzJTenSa3gJcrGde91m7Nb2OMSdaFoaZWvsZEOL
G6jIlgZDNUl8ZpLxo7bZ/sHDEuymlUjc3VSYg6bDJumPKIxhmALUG44gPRoa9Pug
Ztz5iRN/WVW1a6m/pJC0TdQLeAILNaqDSm/x2T4mkXkmHzLHgEzAzjhtbEUvc9jc
iNyIUD1wQ04ofZMM6jrhIvrRd6pXckwHoPAU7NgHPnaQhMoISHk+6R7ij6+9EiFv
rIoq7Xgpv+Smrcanq7I22rJqZQ8jH6U6Lzp1Hf18hsiQ5NOjsyhyFdVOvyXwWeWX
paZwHQZ0kj1KoS8v1DIqxBpnkIz/4VS6PIr8vuj3M+KCckESk9XkuPL30/hqjSK4
wsHfAB6tHZM6Lcqyn4icGsoNikmtFYJO4lRxRXn66lnpXfcSlIrvXjbzWI0QMonQ
YKPiOCYVRubSJPVNgcI+4456XYIPaaNf0SUZfdCkyspUfv0MTH1loJmmXrUWcx1I
yJGGq28XXrc7yJ6DC3u6mI03U2YGioeWOW+bXHsJWbXraiYvC3WRSmDsHsfu2W5G
oM+CbGQzqdpLh0RuFWRE6YxmBrNujMOekCv+ea+h/tLyMs4qMqjT8ZBCQg3wKNaa
LvR8VcKGyE39PuIQPDBWD4NNrGGAbZgIUa3chU1SI8R7Qx9UgW52Zc52HZ5q4w92
WljGOe84FNXgYHOFd/P2iQaQpU8fauS0QQW/0hHo33fwOcBFopu77dDrJqO9DLBw
kVpP7q8Rsjn75+nsU/5qiEwCfMTioGd7dGeFV8Y6w0SeSWy425MpWLeYrzbd4CJS
08x2KbjK8MIJz55opfhL2Keb7s5qU0EQS+0x3dN6czuS3WZSkkammTMRYFmPQF/u
jwKYK5SokoZmS26MVN8HONfM9AzZLCxAg005lnbiRjFV6gDz8O8+d9fB9uMsqdw4
xCFESFtkW07VdYBVpFtRGmb2chkFyD7WyoH/jQo8bhNmH5sFS3zL2ACldEtTVo1j
wtNo9/eC+7d5OzmBUDAdWp2FkZwC/zCSmO0ErKEEhhOiFF4sV/pNVS3vH4kjiY8p
goZT/Vz+Cl4+ejPpLEEBGM3iHjmG1IoopsiCb/r8R+OC3bxvwxgNdDUPivwRQq5C
9lQs2Mx6V2GzRa9ly7Ed8Zbev1i/i39HpNmWXradh+2etNM0rR46ofDMtB9EyV+e
42FyZJTo1JSkrEZS4ECQiRkEjcpy1BclYWnmdUBmxA3KsdEsxZ4U9vWscariGnq0
79aMma/kazzEIsZ1zhZTN5qDNIvM9m8Htnq3vSyzB9eejsIPXPqTVbhQe2qMD6Ns
P+TjTwj1DbZc669ak+SgodUI4mKYUcgi7bqzte2xu1evcR1V1PYtfAL0tc91YhBF
zyFIs2bocKBxmmocCMrF3fbxBObfkXZOHsM0PDscGm4FpJMo36ZC6X2qL/WPU/CF
ZC58c9k45AfVMHz3QISlZM1VVTrRD/Oh844UlzQFgyateO3zJYFAAOXglpGjX1l3
coaup8T/lcQspyT+6/FVoGBIUSZEcZztSe63DjZ83h7tjB/HpDtfifeKVF9qGBe0
PgfjBczLKYHy0J4UTgVfLG/Nj4bMQTgfs4xJOk/jnJ/JKIviJlW7X+JpPTU6ZmNn
m2Ca/ISKxCaAQzAZx+G6kvu+Tc26Mbk80PQu7y5QFvgrV7DMLZTFi6RBVN74FhrB
YqxBJdbehtLkZPc3UGGFlmna/U8uvnsJ0LU1Jri2kYOxfZ+u+5MDo5zeEnkWje5x
6rSyr/cd04GbZ1isb5Mtm07vD3uaIH3N9tTy68iB/OrajVd2o/USzsSxCDyi2T0K
BuzGhBbhwryQgaQwzOeRkkPtKJew2Rx21ohFS2xN43S+qbJCKwhALx/E4FBub665
oTRs8Jdcpltc2Aq6dJL2l9God5Cpv4G83lTBRKP2onx3cuiAbsQSbWu6GsDf42YY
4FODERjUNMMLFIoUzW1F/rrsAVJWoI68aanEquNhgs5wABK1L6++y6fww1qXJTvt
1Tkb3Pdc3JzZ9NA0n28egjNWH1ZzvXRkuknho6TUPqV4pktKvnDNDhSsLPG+Hd9t
33gDRG4iAH7QeMiHrSQo3YYQkRDR7vn9Vovv7PnRw99kkxq3Qktm5opYOh3vqi3Z
NUq2hxjmh1YJrJWMX0lhbPq4tCj5xLRxxihHQNkk8JDHkj/VyzuNvOd/UX/aNHcf
pwBnZUlLhPB5xKrcTaPcyazbOmYcxugsHuoXSLARP30p6Yf6A7duva7Vrcjb4TqP
JeNhGdtujvpGrckMoS5XK0kanFFri48tgpCsF8OdSG7ejN2muVsiE2laIkLkXoge
7eLPUkk37+hYt+9/tvVYL4WV6unpsdWeX4rCNkSozuIxaprl0ngxjwAukXL0l2I8
XNIN8nkKKgPN4UprYaFHOOH+OKqQsrHa2bgXGxlqpf31j9b9QrAuKhB5aQq25zNM
qQ2nsacHiPYscBFLzJNuZ0RgMxgUCTsY8GcN+bgWCOOGkASlHF4O1jFAsbG3VA5F
OrQ7ct61z6luPvX0hZEKiP8wFJjPQ7MD+rmvAChu6VlPDvrdzccI5g5SrZBHt0HT
NXv8DUlthYaJsbPK5yvtwsPSKaDOZhzfxw9J0bhhh1D9C/SfaQyHwdYLqrBspdZv
tjGrHOg0H8K8Qzr9foV5pnWTIbksav0l6A6TPrxvI2BmpNEe9PDFFz71advNAFGQ
Xw2a0qHLnxslJrt+WvjUyaRgjgUzmscFurDle5o6nVUIZwQN/9P/nzc1j/1oA85M
VbVqRAzAmVkxjk8jBxjglAFHMxgB8XgJ89v4SsBGoKmMoVMp7cFP9sqHzBsBOfBV
HQK7zRNAApNfsTchADfUgvq5Xh7YdHJJeWAgNq3JjJ3iDMoiHGujpI5mUDKdAlfy
SONI6/R6rGy/NCEykhg0fcF/66qOB8NljCJwtaNYKinYqH17ToprgRzJS+2yK1KO
3asgTlYo+OGroaEl7yIb8loJm6wLYVBjG7K1rNM86WvKmjVGoYcLUD8XvNLqUiYZ
UgWvBI4UkyUOi2mit+TxSnvQ0taJs6oaMyieVnnK1L0ou9yffIH/48DMSkn+DmKd
vWRo9f0F9lX3JA/XVclJpvBU0zzQr+YeRtm1vm12ELxQ4OZH2cDZkk5tYV27tfMf
IfaBHxmTMq5QjSMRS7XPv4QAB4kDlzLBSsbka0FMPfEMMXUx7fl9Q5tg7xKQrRWn
K3a02mA6We1K+N3r0iqSfuIZ/nuFvak/ejFXrQB+3TMWirL3FLLYw124tQ+hcPxd
bP4xpft4FnuhLqFH7V9opdcccFtsD++VpovB1LDRhV4XRCJb/we48EohLJsmc10v
NxHCET84v3YKgzU5nT3DGbvvyMOgmqc/zogHEvQKJnMFbkb6nMLJw9Z/CBlRAyJw
l8BF846Md6F3OcCwUBfI2AkUe5aOqZLZeuZsUJHOiPmd0BvK22Y556GC01Fb/ZwG
vZyvAglgX4xuTPjnoRD/hmhIqZIgmYOd3AhvfmqzFV7LmyIwrE9PBpM/Yj6az1Nc
1Pf6FTBwxCQjTrVdspNXKULcb9XPlZFtozqkNTAY199i9DBfzcuIPAik1vxMrvvU
HKvwCkIRbnSA4ighwHPYi2QFcF2Jtgqps0hjVln/CjCZ4D+x39nPmTDOmV6tM5yg
vFwvR/0MjyvtXlttHDI+55V/qNFgI+esXn3i0I17nYu0wMzhJvCUh0wzwJCMOpvx
2bQcGvyGwgnUYrarHsaZiOwCFaEgQC+LgllQ9BxNDeS+raiexK733kHEFUQd2ZZk
8WT9kJRWS4UFKVsd4XsQp2clEDca/GwJjINRquwQBbgriiv2XoRdOOKQSiFhej6w
QyxqR6i53f89F9EquaZaPv41utw9hU7HHJAKfMnsH/AfTd/6K9/9XQOa6NA9cftN
q7PuzCZHZ5uZJ1+EVgArdRsBoRJqnJLTfyrAZk5f/ynaZjV+dNvlYCzUQSyU1pD8
qAd4vds08op6c1jw+ZYFVpddnOnvDV14cb2ZZW89lk3xyMwIxfLphnoSnEjMXLhF
vWvlHnMDSLWHYYoTHCdlXtHSXf/S9jPK8AL5S1zcjfsl80z8etfzL4iExwcDAE41
30B3Okta2zBXfi28BBeU7TINjkLf5P792b5QxpRf813ecTBvrOo3DUsTcXjJZEkx
f3IjjzHxtbunw5+8Ig+TqHiyjrwsiGMj2gzNjv+eOmWiM1yWC0aXGBgS5O9Rfl+l
9IosAdHq8oSejMkeD3AsIXCXKba5eSX6o6Ves0XTetUwAsfAAyL+TtD9ybxQyJzj
0t8SuYBfPr0i2yU2cU+9sbI01QN5NvX3Ht2et+jTNuU0FpEkYT0FnY0dv8yM1cCW
sCxmE4krAfqS9CHBKSVCKgwyVFBurrI8xXon5XRSpn1jJasRxsTA6c5e2lpRDcqk
dlQe5pprFeqmu67AywGTiN4wJKouACG3BNPCdejAWSMSKG5MYjx/s4D1KES2qdqO
SPdvRczJ0ce6tJuqhp7OYKVAbUKMJlTuOB0Zx+KZIueLqg4LNr2K8cZkP1y1qJBS
erVOcXsVh4qV39yz6DQH8wQXakFsde/Kn17iYGA1ATtBi3N0J6j2V+AG60ageM5z
aOxfanfx91gct739xF9y1oLdg8SgAcW1lTT6aGcoubMgifCwz6OE4uo+3dXkIuBW
+gTGpfl4/3gJjFNii1qHlhoW8xkS4tFrWQTBD4OYQE7HruQQdO7Xfa+WrbDVU/jJ
T0acxIRw20rgPvRJAT1QcDLm3xsjU/LdAHP5D3w9YxcCyyutvmo5BU6XKPuTWAsD
Bggh/lFxsqCiDCLwdleKETcac3hRxel8ilJd+pWyJxR1fTj6ywYaBeGBnabEX1x5
H7c4pJ8uUP+X9Qn32h4k5gPLdxAdM2VrhptMM19a0ea2D8RujKDtWULS2E5TLmvu
gmXBExzOyJq0V6cdolM5C0f6dsADBysHiCbDUaLO+4gksJAkZOJ/venI+i5CRPwb
eCalF4ctiFK3/jaqjAudyIpp6dzaJp89lkBHdR3kZfVHdgIucocxEXVAz2cal+31
aUdrxYa7XoroOpa6mdTr9oi/lduO9o1Dhtilj/D/NqwdB40w8zLLGjnixUsgLJn/
McS6tigUX9lo3z5VGRRwpBmKWKfHt6hUY0Nh6uMVYjInMYeoyjgSSV9Fw5Apsx2F
kmofju7CTfRBaukdy02r0x36NNI0gfhqGraV+PXB/DiD8bgYpssj20CvZ2eKIRoY
L+iwW9oupyBktDPtjLpV+V/X22+EAEmvtX4xT3d14AWOWU65sE6NlEwD0IRqaLxP
U42a5pCCTfO/xAcHPOD5t3i8X6r12nCT5B/yCcb+Dcseh1J7C13TObrIdqOvvBE4
Z9pOPE1ih/xhSpIQCwWg6p5uoFWcmradC37f3f+3946eVoGbx8rfkD3/3kPZnLWT
MmeEmjrpTn5cai8bDODODd0U3KVqpSyZpndiz1sBF8KJLsG1FTszpN9TY6Bh15oY
uXJP9n0f/U0g1NGL8HS+EhMFcWBVDyFCBiVTya1FztqSj9EH+yxFJtBixRWeh26O
ZcJfy8E15P047pxKbWxSwzIIRpYvlwGXDqFI95URo/qYjE88uNz4UubPsMYywdqh
n6yz9b0y7k1m3VbZNAQeqTZxjNpPGryxfksbhcp8A0UZu3u/cuUeuMIDm7Kmf8Wz
yGXIAj1DzTURMkxYmkKY1rICWvzOWrEcNE0jLjo+aNuw2KDoFujVyJuXuzM1eypI
nOsQRGq1t0nezQ+Gkm1i97A4y2EiSUOK6Dv+LTSBGeiovs2bj7ZezzcaM6Pxg31h
NU+/j+xuEHkKLwmiRMH3Z4u6Kj7YhU7co+2BgtTcXYEzVf/cprK6WJTivrkiX5U0
nYKXKxPYqhgOonHKXRjIFoPZ20198frMp6UCtUp8FoOUGQESmUpUkEURP5XSEcXD
jPGB6uh+qQbRnUfTYue0M943+Go6vzyRcsxSXL9zKMwD9o6GyoedBdbc2haBDNaw
Vyf+GTO3V8ts4msJ9AlgXKI6ukD0oVbHVUkDGuLX3Dh38QPS4tMpnD7TynqFeqg0
r8clH8mZpUtlkKjG65PEg54NCHNzToeWF/q+k+pjjHAf+gti2wCipGUP1vkVHDtH
9cVuZRQTfVSXB17sRadlaC8OnFJ2Jv9VYmhi0gtCacutLemlGEmbUm2sZXnOgimK
3yFWOPC6dl/tr322kDtXokFHZ1vmKGAWWQ8ptJ+Mt8LcTNOL97RCNPmnty8PqUjY
47V7UtWyDXKkpM+Xx5b4OA1m3N9BMjRjv2HR2QIIcJDXL8d4k6GMRf+2NPRuQm83
VzmdcoOTmYMgy1eIQtbPgGEttjkmec8jx4zQDZM7bop0RB5N4A0CplQQ/I2ByWSX
1WNwz1vFPVz4/cq3KG/ea2k1aWHv0+FAtCiofoT1HuTshl+GDYOOhcpKj7/XhIpN
TeLKSStK4OZew4tS4U7Ei1f3TRDqg4JzaAOi9DCKs4p1ErbL4DjWV92Bv4pmJwTK
vC8KgM/e35wNtMRYBckaTA19crui+L7cjZxbYngmc6ZQQ2/ymdFCi1FM1iXuG3x4
R1JaMTa+sgOV80k8ZdO/+9C+3o3Uiu1qggV6UvPMYRmMcTVSjNRtZSbraZwDhOaD
q5jLOYd5LU0mkVcWRoOgx2xhvfcKuc6EUH8XqxXPpNnIZJ29KwJyb557Eus8zNaY
1uLyP4T31OQ81o9fL/A9K6w++cESyIYKF0meUSjCGpYw6jwZc77tgZugLyOO0rEc
jOslTm5BQ90bQhm1cLXntcPSfWUNwosF4W1GxozNtLA1hol4i2wKjVtbEcF2Kude
5dAdGweK/TEPKvAIqDC5BxYbcAKPpgntlSMvBBchv6YClgGhrWsxQzsqGtjBM0Yq
+plZznfo2tnlVXzou0AFOq8B/KDNmjeRRLPeZGNPEtbRwj65xMDvt9Z91hKKByoS
4xv991XCEMlrd18eSP+GsavAQ5YW/m/JM+U6ynqTEHFKGOcqohefD125mF2U972m
dpQ5o3QW6PvDnhcJ1miUrTFAth0101pyJGNo4YkFR1hjJ51JULznFqPd7NQUSh8V
nx44NCKZgj2fdv5bzZX8LeymNcqaq7H/oUPdVJ/CuX94qBWyMZr7TUWdb/UdPFID
VnIGDTGhN85iAYs3z1SjdqkeCEI8+B8EbZ063+DXaEmwx/7gQgG0j6iMQcAFer2t
0c0Vs+I5CEaTJAlpiB1A07g2Kr2NSclgzI2owkt8Kg+EIcgxrV8R+1CmRW0VIM4W
Jiklf9xw0alUEUoB25GebUFJgEPGCJooXKkv4iOByxQITxuFUTFHSWA3wYnp8RzA
Nb1GVtGk4/mvqCdCL6mtUGs0U6tNL8+TT6+rOZzwvAQ+vSovFcO5PUiw8/ydkOI+
ofdUlMhj1CYeELUgCLOyYppoeso49wwc/h8EAk0UAMuepBFYent9hJIsqR51PjJm
79MZF4dsmhYvwUtM5EhI7fiG36Og5XJThywC4ZYl0UvBQVmSLa9Mw6sw3luTXQoa
6HA0ttgPASc/smLWQE+/DB8vr1TWOEipw27ImwC5Oo7AwCaHP40GvWt6NawEz05+
yhok89S9NEM+fvPLddT/gx2rxF6w/pVkr1+Aupj0ErdYxSw8RuJCxplOCeLTKLhA
1hzDKkuLTDw6DCNyLbaQ7toDQdGOSdTD+zBKpkJSdN7SBXO+IjVi6ZqbUyZ0Qi3N
6HjVmD3oHzTvGgwGNJ/dgJ4O43O7Qx7m21RihsAHxsNzoHa+bvkJ448kQlN9WN2+
Bfk6mL/j9j64SNCiFMjL++mDdWeIafBaG8DyLWuwnJyM+8s+oLy7mrUzEwptPXKl
keZVp6XenD/flXyaWmESbJcBYOM5JXLa//5Tx63NzzBhlx+DABqIsjnUQGfhyUr7
1nhARf4ucTMhR2fOSAXgXxmnpP8OmWlsMl5NycD7lP7xIJQNd2qk5gwXkBXacQhw
fJ+egFMoJmPAJ+zFf0c7Ax1XwMok303k6hpBlrxwWiUuzl0fmF9RYhqAe/o7omPe
ZBK9/MihTo07OF/UAHLHtPhbJCWfYr9K7KDW5EiS3XfOtlIHjQj6W7qWI0I11Bg9
Dp11wrdP1Za43BDnfaLYB3945chdJnEecBHRtp7Slo9DCtkxAycXiqKregkmsRrW
ilaZ5OkjaK/C23FJ9qlFP8rZ44IOcAm1qDGJYh8ONWKUoxWJa0uZde4jWBnxlct0
ecvohjnsCyjLYrH5GqovflSf9+iDDKUimY063lNEp2phy/kDfeILFQP4vw4brT3S
cU7ah/UOj3QzVFyKl/M+TzuJNqvKNwqbuM3IkLIWBwYeIg5Metd8tBBWRd1M5TGh
hJ+tX4vw8xSDdyE3fB+9rMc1QS65eNKrcRZDihpuF51GolTl4r61+z7MDyPdpEw3
uy8XUC5Ut4Mrr7WrTUsKFMyxB7DcHYJTqu4+wEkkPVSoMkCDOZTpLQ04ognzKZkm
SRrICMRxfy292IHLGDBgo3mQx7R6YJRt89YaCN4ExFZvK6UpLzIuxPyfM33WYCKh
Lnjg0jp0jbB3skDbUqKK1uajnEYpUyPiEey/hbDRJJHQXjMbhK/R45tvRJ9evlrW
q9YXFBrk8PYgyFQraGlY8OBkXbOCP23E0HW+kYOmcnijsmKWfZAbcUtD4cWEHLzo
HxDa60fcc8OTKshs5sECtPb4wYGB5Scb0FNB6acKPhRxAkOGgNontyfDrRHhIkGr
GTf93at8lUWG7AxNNMOH/gvI6nteN73twm96t6ZMIpsaQCSk7ZU2F0SzPT5gBe4i
FlveiOhbIpFXhFjskh6umne+p9udGL/c7Shrq7r0nNL303FZY8hJzMc/mWT6tEdp
U2D8g6CkJWR2GWNHSjDOnm+s/E9E2wwIQGyLP8eNSVYjfoRPAWto7N0Oc2JqdiYk
HsO9K7p1yt/skA1oBIG6IlyzX04tztnOTVQKJJWJmFTl+cZe6/2jQmOBitGkooVM
PHmz1qrVSgruWLSGx11dtTgEi50P9jMoMcgo3G0hCmlKw/IJp/+0yCMQ1wrTSVfq
qsWBK0EvzkX5AXePd87VDhB7ve8j64czY2rez0ulNLXMGIq62ARENPxWtQUgfOX6
5GvLwVTz+Fi7kTGGi0y6nSwZRxdgT2XPLiI6hf+SdHbUrZnJLGKEtsTNkwp1Sm/g
fHiTj65aGhPFNtrW05Ed0U8DCxCJhOr+btfgIrYbPoeVIJqIzc0t3Sm81MxKpjc6
kXwTKkCXArHXAtTDJt4JpUfiWettd1eX2u2IMp/EZU2ehS2zcv5+cUZn5qNf+YnS
297OlCDD803yIVB3Zbxtl/9hRSI+nzgRTdgQI2OtdCdZZdZDzBm5k2/fCuAI6MUL
dRYk9AigWMu4cVLMdky7ulknvSTyR1LnMmQEcb6gjhX0MKOL177XditMpvktKSPm
R9zH+GaTasa3REP9pUOM1OdOysjU1VdI1w2GMeKM7vz/20jy2mA0bshc0pqkrEic
5pjiuxs6JNsqBHXd20zY/iPe2Sc03fKFAyN9+R+dNdrY3/JyGDlvA4XdNaViR9zJ
gFtScee8hziTfChEFKM5DMwCo0ZRCgOAFWsUTJ4MSRBc/JcjX6yKVzBS89CblviR
yomF13mwi2vDnmc0IacRGtfhyP0VrYI4wqK9+4fFxQxVgRmIKBZMEFUnttHHweb6
8bKIFsg8cpzlW/8dyluRICOol3pyueZMywp/QsZ/A13W6mM9kwMn9BVVsClwR5fF
KTBM8vSxFnRxxbuQGLWvLZ08+NhGVTSvHoYsZT6/I55v8IEocx5jdwQM1+mSuU45
FWdItWY2iDjvZZMSRua4CrBmO89oxbylOjH7QAW8qxxLx9EH9++M3fXI8emc0kBE
hPcreLG+EyKxwtMieu+/ns1d/FHOZCOnrAIsrdASjWJI8OJdMP0L9Qv50co5k0Bo
+z62xiORd37KDKXuMsvKT0AOZooFITvyCFv8YZjp/ezPJNHL6LcXps8fFzmsIoCb
x59eTpJ2V372Km391vASRDeIBBmTFKMG4Aqi5ZP03rbPf1fm9f9AmT/E4uARR/35
3wRBc5x+OZFKNg69ir54aRGv0flJ5Z7iovkx7FbBchWjMkjz7gOL9E+LQIAyf+CY
GNOqrPDLXqWxdFEShlvpqxGNIRWLAQ8RDA/OgRzelU9HtPIhAXx7s4iu1KPSUKSl
hO0mqRC9M1O5tHxJtrdrS0bUsvUHVCA/YQj7ttQVcxnh+yKHtSUh9p1o+Zs1RcyL
8woLocaqaPJAr0AWPaMR1tuMA/w5lYnBEUbZUQzlJo7X7X5BWkSKlXi3+HNvYmv1
rjJgwe07DVfnVyvf8srWA6QFHqzXaivWr8vG4fEDIvxpWitLkiosEY76I4a5REyX
oWWaA+XF0p2et6EnGW9NKl8I3wQdGTWw0vLe2gbRoHsMZQHnqPfw/Y5U7u+bKFXN
L2XEA63rL9K/srSoBh04lF+O4T82c7OJBuKesWfcHMYC+T4gN1SKSlywKEsooa4x
mPfFvwOBOxnnoEZ2dnLfgCtqq4WHmf9rUby3UdZkP91Jirq7wGhd7kLHrCtoUjeP
c7JhNdHI9KWAbsxBsTyxzboAF70S2MMnWGaJDgy0lChNo1Lnxv7V7bt0f0rLIQup
xUZnqPRGHRLxoS7/cHsFqk80Co2c9w1aC9OjPWcX+H+dZecWQymdl/i7FD5dPTVC
gPvyHy4NMWGy62Wzm0IyFQHeEtre3gNc6h/N1ZqHijS/fkC7ERLb6ob5AEbJDnD3
LrX76YdvzQYobeXtojQgY/LiFKUf1jW0OxRdf0/d8jw8kh0SjCnFg5MQ/fCyZOGc
lMiZfHjy+wDEQhgZsiLeCQm8uTvFCZu4+GrV2/CDHhrlySXxIAxOxC/1748kQesG
5pW3OPbjcA3X/gaHawE6G3btUobOi68Ui886Jzmf75gVXScBLldrpO6RP13LJztq
VL9ejQku1yj2a1awUJuLtV2wRaEuNor9tbLkHg2cYOI9rSsEJ4u6ze2epxdtPLwD
YL0YEEbH20RA7eNjbom/vf932Om3FQQLqn5QryK0ms8BCwqqRW3irDggcqAQrO0G
u3hqkexiXBnB8R4AueTgsnPFBhuYuNQ6VU2fJmG1eQHUWAC5+9klSXA1hD6RmlxY
WvBbMBzlmCvPProF5INp6LHIhM0krA7RsCLljxO+u9WpF6aikks+ouk8Kj50BrHE
EM9YlF8eORLIwveiBwUeMabyuRv6IcZUTpdmed2JzAs/9iFbwVEVIGKsLYrghd0X
NnZOxyCuhzRaMm5/U5dkJJdVPcLxJ2jLFs2RbL3EJoXLCjOzCSMI+F1rO0f5hHw9
w7RTBhpnbr3W7vr8eZ78tlf2qLEDPHT0sobBZD8E23JTtpddR2ZsKLhAnC1AIrfA
XQ1g0cAmVQjBxMbDKWUdAOhsn9tYkNhEwV+Ak8p5gHgyct5JlKZxMHtCXB0YxG2k
buT8RWnnHKsvpoxrA7duCHIKh7q7yPYGe9EfBpID84WVwbQ2zXhiIwjsvEX+Euw0
bFyfvzoi9fvO80yA+0CggDd6ynsHFUd1sUrjbfHHmr04SpMd9QdA9u13tS8v3Ksj
o4L5jYHGFtZm/VhYvvaOfkgNp0pFRUrCrski6O9i9Z8vdOR4NzCD0F29Oud8sol3
/zCMPMlUFG1XPAIhnpw0rZ1VCuRCj/ypys1Xuw+98k8X4GECW6J0Xs1SQ9n88Tq0
/UrKzYnH2KTbd04xbJHXPEMJg6y5NF+aIXWRdI9g8w2SY7PL80Jdb4dxqDxTWExB
Ms84PVznY8E6Cuff/mHU1nLDngLnG3UiSRjRVBJw9QhzQsm6ooh0KjeOsEGmiV0i
gKkQ/HX9e3NfXacaDkChDUnZSX91qA0SgQTTJGgzCsiDndVwYLxjMmahMOqj061j
oqq0WPgmvySYStf7l5krHAzmEenY4qFVClP1B07754X+pIyc1CuUCK/cRmVO97WM
YWH3xL62noLQIukk4VB6sJwjDPh1QFfb1xk8Jt76xfgp8VlSk+uzVo52V6A540BR
1jJ/9iw9SBVZMmicTQt0H1Z5hDBbjTeKG17XWVuOXyu3YcpII7iMs7SmEjNefPAT
gkaU3CO6pcTTP1O2wrIPKrZmF15oZGYKYr4rcgS3cINZmtQ7zgwwp9lQBw8RdAF5
bC+lXFf5xkGu2NqLkEY3nPXhOeAUOIn1XAWtJ+YX6R5ZTlcP6M2dSmzctOwwXuyD
vi5Qy4WYLxv+l++gOnXXVkLAA2VZUIWOjBhywttC03G+DCTi08iD7gQn9R9lXYMw
R6UEXqQRcFSPH4vzD2dQ3OPaZFn7El1bMZhDHkvpbmdbaGkOXLPED6dQ+bX7zXzJ
bMd8TGIZKt91nrLRRVPnaerEAXsB/Zf9lLQjD7NI2AOL6+qke6P1ICsoX0kr3iSj
OeK6kUDynbW7wElaOBuQ6Wauv86jRmXV2FMwDbu2IDPhki4cSx3K4WvEy/TSa8hJ
SuVwGbhc4P6krEEO4TeDZ+sj3vnAtgm8qrKlxAREc+Bsy8FOFQKFgulAAo0vLRSN
TXrKgWoO1Zqye43Tak2e+g3rWApnX9d3bI65xtqhm95XAF13KlBewcQhhbuVLtDo
i3OlEXh5Ztpl9RB/rDZf/kEdvAWDI/Jw3o8j+WePm6Hg3407SS49AwNAXtmwTJnf
RrIHhMVV/rdC7jTWyGAblWLa0RPULTjSd92K7YfoYLUa5n7gpbgWvmiVTpWL5iXM
QXeQZ7NQJka0WxB1Ry3U1xwynmDsxh0bVge1ycxaFzWuRqnHkkSHfDTluVbn4Dxf
4JoouDuBZ/eO7Vggwc8BImp31fPv/aWGAlTSHm+i1cPdce0xD7+ZnZdQImjxXikq
xxdWTa8XId/8++ki7OMVINywNWokRwwp5UqrOXJP592xvFiVCPr1h5us/n4898wY
TRVqTiGCh4Did97lVQDmZs7Fzs98ekfewuWutobybjOAP15Y7sV8+d6tqjqN2AUY
t/PqAUtY/QYMohkdxBQDOG7Ufd+oV+b5H/UpS4a3T7dfZnfdw6t1qhy0bFwYvENi
WRl5zO4b3VRuTnl+SXuvgk3rEupEcfnDRq1ZE8V7fM3qNbNAAwEW31UMvfh3HPsi
rU+78PETvCwvlSSg/E1BMtuxWcFkqU0XWf9udIrkFddPb1ipxJaITPsEVho2flcQ
k91WGfJ2q6d6c1LAE0S1aSFlsnZmToHQn0oL3xfhgqFS77WNxhjNVu+wibxVnjNH
GZACBbqv2GqJscj4yA33Ifw+E0kojw9WuvypSssBWcFMOd6gv3aYf8JN+HYaldu0
l1ptplBka3XYYA4JXTNPjQ1U1TRYYUg7tMNO9ojrcmFJn1YqI+IDj4cXU7i1PhMs
7JPxwMmetifYaf+hERQTkyDyV1qPoBkdn7y6EfG5RBJExvCVLoVN7QtSvKB2Ke/D
+eUlm8V0ik6qQStzpzGPql53FDqaIs3kt9wnedZB8JD4qvrZGmPsdzdp7HfVRHd2
lEJ9khozb8yM3JIRGXEmBGmjelImz06Gm5xmnk/npLRjVsWKai2PuE6ehTwiFRqf
0g5A7VoxGIh9OI3nESkd+WjxvEbODzHGJ/4BX+LkPXXjS4jrdMRaDqub8MvWtf/0
/vpbDf8F+FfFo8IUjLnzwNHRpbb/PCXc6MzV56C4wYSvW7W49lW+kpVWCIk1NQee
RVBDvHNTyD94xZ7YgU6HkacCTn1gUVM9fGV9SoggEH9gbcbQsCpIKZ62sWSGH9EK
xtl2UmDYgREGJdc7JZlIZynDIo4mE/hK8WfcPF4Ach6V7wdsvlFx7Uaqzi4vZMcm
X9fnxRw3T7MZcbErmxdUrAtuNdgdhDHwhctJgPoBTy07IqXGR8hhpgxt4/IsCVw7
IBupgROYcLQeAIyp+QHcUimF9xfh3y9LrDlyLugn7RcC0ZKet6E7qhQX+cZJtg2c
/54CzZs1BHn7rveh/5qFjSqCvNMMjNdTEXeapMA3Ku9ghXzgnloviswJJRCoxShw
M8digsDzQbTiGKEbR8K8NMKveTRFaGRKAUjvEhVSQN3qsueYiAuUre1l64TLFzFP
bd8mcFPWjzAVHTuADCi+H3azk75wFqoaRaqVqn0z3y/NLFAFMWWDvPYMJTD6pzJP
zfPKu1nmSSLoKVhUk+hCRPXzE40eQUMVMkJFH7YD4bSChONULXkz0CYHrR2vPLYs
sL+ljIeg7vYP2yO9j2kyryUEjNy3WGbIJedkHiVzBsg68LwwQJ/YQtdqzhmBnVNZ
rrf0SdhRfwjgIk3zESdWLeSQ0g4zMPQgkMz6RfzJaZB/Kk3wgIMb8iY2YkfAvuxP
qUerl+fU+V6Pv7EOIzAJ/9NMQJWkcrPYSdkVK3CVFyTDnK9Xx4kF0FMxIMHYK3Md
2XhjbvPwVPAgN/cMS24BdYmjVDRfiyxUA/pJECtURENIrNViQMsD0n0u0CKMB7Vc
7UxQEtgQs+Ej69zpZiLEFLdQsPWlYq4LaaluoVmwTnKjcdYgNO/y+CgGY/Jt6b41
DlCdZQZxU8l3vzYZ5zFsGOqfyV1HZUMXZYNNCSLV+GL2kPulgAhS6L6plLE3E/kK
6yYfwI6NmgQKpwWW9NC1tfeRVaJ4ShyQREefPlHLIOmeEq8KjB1OjxqIRQUGRb/K
eov6vBT3tvo3nDoW9aTajkU0/udKOYM//UFeDvf9OkrZJp//uYnrCeKyO5VRobsv
HssZ17P6aZRa2RvFutRCCvcgVQcX/W/Yic5VuKRw1YzD6sFir9Ni8okvq0Kxl5AK
2uxwej2W7jTlnlAlK0bO1EoKfLw+89IxWtdb6VIBg5HlPxgKYYcJ+DWkeDwlVmvF
giaXv9MU8iBkRy3mr4ywmsiBYca1svcNKeUXncIsZyBk4CU2ec/Sm8++3/75Hkwo
xpIhHnynmC36t2iVjflmKst3l3AqmBRTCfT45VH1tfEjfm52s2qqFx4ls+Fh9KvD
Y5HwA2KelOaVWSO2dBKTfyT376SF8mtHDOH7GiZthTS88A0VTi/XapgnfhCcq6pD
zvt9kfGlXhARv2FKwGv9+nLzQLEUZwAWD31o499iEPKgCZlzYAil2bNQoMWAN00/
ucZDW/MlV+02aHqY6RuS1qxQYTVeqpPycuSWyHrCmyYfh5L4d/j4/nnOXULmG7t1
jwCFB/akCwansCYBouqvbrq431AfdCURCDh/V7JhypydEtIj9F3zM0Fax4jkIDSj
MgqOv7CHRm9X3aPOz5mTaA4z67ba3WRsZhYPbWSyBhOmXGeb1oHWISz57DJyq9f5
LqL72n5mwMHjdXvrZepYgni+1I1wzs/rpdLnbY5Z3EBewGshTQFwFyRzs/mSJmDH
4QApH/+0BU9F5wd+Pl5KFv0+zgwFFumxOmsahvh+JRRBDFUWEJSp8D62DHIGyuIR
X4Z1Oczst/S2wQtmjcxlGK9TT41hl3Q255votmN5cKSeJQ/RSS+wo5hayU+klcT/
o0nxfe02GkcyzDjyJTlDY3zyGc+OlxukZxSSeL7SdngjUiqb+EHg3Fv0JcSBPUkG
Cp7zCfHtuPKlFlah5/qXJ1SRklo3oNLPh7RBvQotL/EzifWQUHraBR1+xtsn+EhA
f4xyfjSxHG0qpNJHyhZz27Qjhw9UgWl/T+E8qMxjtlIrCw79aX+EvWDHtkFdqvkn
tC3ZDolk4N4vWFx2E04pvTmLlDbdlMI1Yncl4bd5nHyaCyx6Wf8chwgx2OqbGlMC
qeRCvhdHTxtR/KSm3TJlDguRW/W9ihAtidPtiYRJv8ybtQZR5RgS59wNLBXHx6+e
aO+A6pz4Nb50BBDYxPbf29aorCj9TkD9ZuXo+SJJY7KelEOozoAErh8Xoe5CXGxj
M2yX+rX5cEt2DvfK1rTDVonR6Ztp9GU4QkpuvLGP/HMc7yWjEayGdVwoFCcK8O/9
ORIwDNyI/zvkCGkLh+FBc7yS/a6MaW5xhZ5wfvKnbG+W9nGPh+Zb0YHa4bTndfkL
m2gOVsMgNbvxZ1rVBmbCMkc9tOo7iqz02sPf4Ai7nbqmU/iUBp8kFcV9khEDUq4O
6DmkbKHCw6zCcpGj8uSdEN4TuXV2ZDKt7zTuMgh7mmjAPA7jJA5W55S7i2YGSzhz
YH5UHZyhTJyRZCwrVg/Uluj1wBQ5EWEjGpzLPeFPPK+OdGtcMkOBV1yPbjS4pIPD
k8L40JDSl6nwULvMRnIfV+YDgcceTJaUpy/Fe5FjG2ZfW6H/Dh/qYQhucqdWBLeo
r2gAFQqW/m3ktm1Abg3ZUxJfdWDMNF6Afc0buivPHJ/G6xO6y+Wxu/YjNfGbOCKG
//30e1ANE5hzKEq/cAfOtb50KwbZrHRT3jMVYjolOOJW44yY282dgweZ1G+vPDwn
uOwlYakzTq7c657cpLHFzMNZXSKuROXtRQk4HBxdtdiqxJ2pxgV9cC37njaWSSLe
XUph4KvnJedtbw7Uf9Y2xcO0ksK5bqxcD1u9YiuxRIpmL/qxJ3Qo+Uf0xOgx9YNV
sdj/sLZw8acZiYowBH/BpWalfyWaZ6/wXqxjTAdRqv/D//I0qq9gP67xMexx0TjB
s8KCFJMpKP7uW0+BgRrWRHTj/Z4JhBQk/Moyagb25KEXkzMrSWThfJ7J4RNTYAWc
aBHdeZR1omfc9pg+e9gyi1H0g80wkd+23PAo0JZ0PrD0AReaLiceyrWyiIskk8Xx
v6DOvavn+A+V3IGPnFPJypdlHXKCjODCBmA1CY6d8WrN61wFVEjS0BaQfPLhGQ/C
w/c+gi1A69yaIHZ99jfzz/PLrudnhFAEzS5+0RTEK7Y7jkPFMIUtUA2qBdB8k+Sv
sS8K90dd9CI20I+B4fEct6pE9Ti18FWH8ixG7/Hwioxuc5O4bN+oSw3Rt/N4wXAj
tkN3s61BKoVIoHlm772ahowNfBsMcg7nsddRTgaNGtFQJ03g0KGdEKSf2S1dSIQT
dUpa0h++Ph6Bn/8GZt4vT+Mfx4CZYkgj00DQn4wIa69fmzN7IC7+SGalkktBz0fa
4lN03xfATgHcYRlFq0uHrhPmpWXArlePKpwWqFsgJyNEBAcHCAbEtS9OL4f///p1
2SupiqcP4kDiTcVkUONMmfEB4DErq2K7XclyySl3eQx1d9CKnMkwQSwJxhuMYfxD
l7060QK6KUGsVQ1JVXdAB2cd0960I7bUOPwxcQnScZ0mQWQWjVwNbKjhaYAk4wSj
2wUPWwLk/hCTBQ2n+i6Fa28loKnC1H/iPmS3krYxvg1DoNsT10yJA+ZoPIQ1hFfk
tOhYrH/YEfmTp2+G6bZxs7LN7oLUZd9jiF0D/A61ihHhdAzdpn8YTd0EAY+fTFXR
pfNGTkCOHvqkRwR6YMCbkxHtKZIVPAnUe/2PiWrL8TAlwx844Z+pMHqhP+/03d9v
wDyXiVPtfY1HaciJdj8RR3EObPG7ymXnbtS6GkgRK/DsAqby6jnBq9nQTj0KH15P
tt4eSt9nU+Nx0ViGexC/NJjkxjEhba+5Z7QKRTxPvVPSYeUI1PVCPcy7LeJyB/Fa
dhXc7sOWn0t7QEA1Md/v83n/a20RGSH+3rCswlj2cSHmDzrWQ7/ow8d/3W4bHZNL
pMEeqp0DT2z7vdcQj+DgSo6nw+6CqAHrsYM5Cqitg7dY+qnecowxpHMuwT1iHrIX
VTNo1q2vBuPKRsZ6mTt2pqJLvoaIpSTW113m1oabprL8Im6z21O63tyQBodhqT6k
/MSb5m6vLjrNSq0EMIt26cewS9bdqhBquj6dDu0Uacc534O62OoUhhtDr3hE8HbI
/jAql4ELyjnxmD8LSkOZxY9A/bcuw7rSKd9En76dk2B/UIS70rFBrKi6JNWI7QVy
AVy7S+NTDQQisgbLgH2d20j6PwUY5QeoahAdb3apdVLsPUWovnK9e/S7JGnCancJ
vMBzhUzH0pB0r2QbDlMCmqJfAfrT+SkVXBy5sx0BXci1rfsPT5qcsHITc5FjabYK
B3Dhv1JUKO0sXOpzfegZjYuP2TEsNXh7M4N81ZnxN7ZmLPluds73Q2il1yPtB4/J
c8aKkWdWvTsIvkAaxn9Y2O+pBHIDNOAd7qBkiiFacecQiQZumk6KTI7CP793Z943
QyCEmRmE07MsKgw0aUBQxhSvLJzLvoc1DGPDz5AgtsLLJFT4qzCBxniutWXexc8R
otYC36BzvrwdivJqkn6avitUXe9+DE9aYqzT5prh60UZ3zm7+/dZR/PGlzD/1Sje
MRe3D/XLpiS+eG2WGxjGdM9cBVZu53TrIwhRqL/iJcL9RG8u4vAjlwbclWMLfRx9
mbjY9tWgGXKNOYUvpIIrXBVsEFrxXMrV0tl8F1z3qcoK2UcJtYytQdU3pxJMamjW
ntuc95o1YhdkkyajdI6DxSAhZATwcmFrivkGcnOcCtmJamae4ENmr2oHWX8KC9P4
tY0h/qzPxOyG0mSECqfHXMf3gpCT9IR+3qAqO2NHPPUk3Xa2zXhcF8PlShqkueZJ
dIeKuKj+eTp/heOOEapql1fgahtLv1RY6sGqwPu5udgw/KDZiE3Vo7gq35hRbbuG
+1mQtQ+2t1m6mtBg9vnYbQVxZ7CaV5rsu+uTp1b6Gne291aRcYdO4520albkJZXz
bPp0p/DsTrWuIBtLUitkdhqUaA61zfL8FBztwkYkEL/6RvNoJv0qzQuBBHQvPDMf
bbJjOBAO7uBAMLJN+b+y9/ZzPrBqLWSCQBDo84oXfnUM0rkL9j0Az4hs2bsWqfyb
tXRcjVra6OGmCunSA/4KNmJ5e2BD91jfNvmmGJijOJ9k/mL5wbqTa6QTD4zoMSlk
A6N9ZdJ4+ol43Au+uKrXsKIT4KcDnqH1lGtqBFOr/vZukdR7by4uFo8ZfYAlYimO
pV482SzYG6PW/3QLO72H7VBxUv7u0v7uwzvbGq9a6LKkbOpTmM6xlwcc6dO3m/Jr
bfUOAcblSTKpadyaSxa+sM2kgrYEbeBSJzTMh7xw2cBH4lvvJ8RKyBGDpjYIrCXx
+HPe3VqyEPKRhvh5ssHl3mxhSueBnxffRZleVSG0wnGtfUiU7TVPsiQ1CAqYKTZ+
s/J/dMC1a8QOJdIlcTlXuRuWcJTbE2I0UUHdHrEY5FUGUUPYroee6aLgIOdEj7/D
rZKhWO9kEUb24zl9SsriBj6FECQD1sZCZ8RFWequ04U02Dwj998UnaHGLXj4Qj5v
UOIeiUbbysLh3P14Oz6kCcowy4aawuvSV/mP40amn/rnp/iluR8dwcZlMgxpyOmo
hf59wkN67FKF9mpzHS6M2fXsGpSjW5hSp24DuQ2/IgyrFn6pABj7DMLhavCLsAD0
20GU94Eq6RPr+87zkd9DaehQE74WDqQsRFF8+oPrX82SVrfFnQKsElXmMdLwT1Kj
MIvc2NxpapX4keSeZmX5LiTSc2MA92FbKFHcbxQu2EQWnVrUKLye34/ZSVJWA3vT
mNhg8QtsbBLLeC15CsYKFgn9wV9Re7EIbjrcLf8Kiu04UGPGCUC8JfHH0fvxFwBe
6CQfl3SyTjz9m2Dly6DHh2qOMC9iB0UwwqPpDYLua0RGEwW9iTQbSB8JrGOPGPf7
q6Sa6HEo9/aeZxels2GEpRHXbt6injqQFQs+TydHZSEaMX59V9Hk08e8Daxa3QdE
852c8icGloXG4Aycu3ncwhg8/15cKi9Nek4swSyBOTfalB3hiRAHvNAySiKMnOJG
IsLtnJ2cFqTDkwhFL5V654s2kjRS2QRAB5//oOXV+YIOWH5KTmhxlbt34s9sU00U
+ZufnYwwH8P80lMKuktkePX8FXRqV4pzL0JixjKNt9I8Bbx6IQYzjq/CCBGh+BfK
us9fGmNDsu8gSVw1q3BWnCYTASFOcaPr5NF2Xp/9dhEMK/7Mzry1HeAxVXk2o0zP
bb45LYA73o5Fj2mrWZCK5wMTxzZLYIbKYLkbcrnMeun3QdNHNDV9NSKQMULeqGKO
P6I6JSPlzFN+IajaA+wuuS3L4ARz2rXa0yfjPrEkjOoH17vpHqaPWG0WaeS8I+GW
v2krVwJyX8LOipxXKIMgrdR/lggGplN+Q96pPv5kDllb4sH5VNmtHIVWz0TlqEC9
O0TIty91xvqvrcRUGmWo6NeNM1g5HfxT/3t8bxD+vRGPCJlIqgPls3lt7RH9FTqX
KaT3ORYkJaDwkjmajtBvmY5vNLKBNd10sGEr77agr0ffEgRY5M1Qk25/A4J89Roo
Fyww1v06ZH5qdWuTQLPYqEX7l8C54m+gwnCXCcw/09f0zE9clzEG58xgV4mG4lCQ
0+9A88UR9umryfwXL9c93rlvHxGHujYFh3BwVSxB4qhSMGoElVRNsctdal9z4127
QQzoVvuCKhj0OZqCyTmFHgFNjPRbWbX9+Z+EzCR+hCbm74ObmBEh+du7WnilVeEB
knr96iUKQJzSH9BeIqcx/b/lS4STn6GFVk6IoY/bX9BRboVcb6YiJ1f2MoQQNhRc
icisedUP8Sdsxb0ElO71e1Bj4h4g+ZD9BrT44WTHaFKq4HJtANEc0ZWeNq4gXmC1
dbENYTjHNlpwOTH+z2appbXUpZgSdcZN7B98OF8cYX3wbjGPHIox31OarDGQ9zqK
TuNKEPIJKssnWKXCZa+Grc1QX3sJQVXT0CDROXkMzH7KlTW5+nYrCbrBhPO9bIYR
VeDFj5266zsrUspsUdjC7XLi73xjrOEx/MqPM6S6FZv/RA6ZUw1T+00YLRpnAFrZ
KI3VrKSh1YMIZbCyunbel4TOw3b2NdMPcwIbuMBYomjr5Tf3O1IJxV9wRcB/zhKG
ovmuWWIZ2F2oRTh6k1EM3yBHBcYZ+53lz8eXJYk8h2T0LosdRLp9IHEzC1M7YHgU
iv/BNWmQwoZsMQpCm58FSQR+lV163i0OsjIymud0H5Y8GA3SqtuKOpAbs/XuGFO7
zUyt9lN8D8RnBUA0q9e78NGcFVGQoTwS+jHsWy2sPVw8JJpiH9iXSRDVKJ5NuPC2
Bh+drXmnMZ95GNSbRrBFLmiup4xz5Unz6AsiziigdAIxoGb0pnv2fBP13Rj7s8RR
742de1eTG+iMeSxX1x8DdY2d0R1UZysT6ngRqc8fAP3XzJYVQTpSIR2fwUVpKccr
hbpwd8OlGfeDaD4frZyWR/u6KQcDhbIue+Dy830Ax+1+W1VHOffHSsnWksir49vU
hOmRgJNfAP8euF42qaCk3JS5+lHm8UHP+BITdUmgI2hjK/+2GyX/LRJgZ7GQj1s0
xHy2hKr/YseG6ndjytXvTAf4TbDZfJo6Pj3axS0fXyCmBakb97I4MjbioaccTg9x
NNm5AW0lOAAMBtcxVDb9tmczhSBKpXVpNdWVDHMQj0XNtEz/8HoVolxqieBWvm8y
2lbMoGzpt4Ffk8QHKiLDQB4cgyj8P+DRZS6lFPq0U8uj6ucfEuYBQgXNCILMjb7g
QRqsLSZUZAptZwBSWrBd459j4jCiHnczBBFX7se4/EcpGT6DDykCiexYdS5HwRmB
X1A340Pw8DqpqoRt9Rx6AIEUoypQejCApr6R1d8lTa9Yoj+dxkfxPS88lhm4otrn
GB8pC9mLJNvnjlWAu2O+97KpV94I/dDhdew72BpH0xHoOLmevm7RkWGHGZ4Os4Iq
ore7toQ4FUTW2RrUiekPmATM7jfRfHrml+L7zY3EFhQetLva6oKWl4dCFHrKIO80
mDjAo0N6LY967F02At63OIAhFCDx+KLkcOzGy8254N2ncwmvkr6/xfaaFAsbq5pJ
uA9GVa6+GLTMMJMj6IBAbM7vWNrfksq4TWRCx76N1OXjDjfI/g6S883TjcuN1lw3
j2uxPD1z4900oj08keuLgEOafeESrPhyRUkP1HFaeiFfFiYrhAJGBq1vF3PCLZV8
MQDCgPokhfnIZvPHWe8jg/n5ua1VmioTiCRGaYvonWV23ky0eKbwTRC08tGAu9iA
VnU3DEp325CMzJoBR4sUStS/dGMftw0h1Qbou5ri3fnbO+NMBVVezTbkiuQApxQz
7fbnWEGg3HIehOdLPh3aiEypecFBoyW5R8pJblT9aiVYFIluSwi40M+Nj/oQ/iwr
uxj4tJttlzgGCU7g/rG2ovYTF3u3bXP9Xy8ZRVdQ3Y9W+LOqa7RbBJKffMSGrJYR
vf5wOMOK9xY8efyIlfV/adbZYMK+v+DiRM6GVvEhUdHY1HQsPCwpQR3lgW/YGAiC
ikTfq8/tX/sNpb9FIXC6OBQUgDWgDXjCncTqbaCP53yP2/YIKDbuDy+y//mUBv8o
ksCnqiiuR4amEpRyz6p2y6+s79BvkI3cAQDOaBSmJUFCIShN7tmSvcq0lC7jsJs9
ABOREDd92+rhbPicP++Kq1Fvpn+zmYrV3YCnwc6okN0x85lWZ+uqLa4PwdnHr0pU
GXXziNZFtJilTOoUn/+moe6kF0CB+wfo9TH+fcwNTY0SgP/jd2lySlQEgMCoKf1A
X3zp1vV83AyE9FifKaAzQvvEo0PYf4QmzMm4md1k7J2dDGiwjHfk4x5BiPJx2ILs
DRt8e3qMHZr0ttCqbA+3z6lGHo4+eIpVwHNAinMHFGyoYlOmxbWX3MQpmCjf1JN+
q3ZBen+HULFAorlm2IhhylF4VXzAAn01FCxkCi+TM28EwEm8ZEbDk445e8H3bsE9
BkcA/d7kC3DuitKV503jthRiGJUhdUENeMbF/l9GTyG7gdTAIAvOqL89S8GmYgM8
08adiwgaxijRkjapRWKpkhJH0jwE34UciGjaA5dohYQh+4Q9skSY9Pdnn0c4TH1h
4Sce8I3dR6/BMw+ijckbKX90zxOSU/n0ZPkfUwJ3tDAD7eUdxQO5crGWR0r9EW0T
Y+bmzH2s/9auj+O5DHiZQkTF9fkL9/rcS0ynZNii82oHMJjwkoXR/FVHOTn6BQWY
QkGeBV5TG0Z+FieVBy/x6ZLUhKdPBfWHEROutO0SAmUQN9tyXARu8csgMc+pUPk5
lESMqdWLGz1iMXu1PY2mptw7Cc/n1Md6eezEq1ghRBtLtXTF8olnSxyL+xyBTnpD
N0/ebWKlMh14iPnwlhDkesSlxcVerC9wQM8SPpksAPl3mopefwWmY1cfJbeMyJPB
JsajU+h65v4RYAKNuHyvLMWOx6P/gT5hL06rVxjRtYfASn18Wc0dX2B9GNyySDo9
3DH0/8XrxXxhnDG9OVUgnTh9loyd/R0svjF4ODrGjxOahbqHsb5p46kbhT/RjJPN
OHhWbIC298aQs9iOxZ6Qqyu+Y2AwWJbAAYFBbdzHF9y0ZjspqPSg8cuNHQ7Z5Ayd
MxEsJ2rQwkohlbMJkeVQcqJm1FjrJWGXj+/TQHL0JxpBEAjqvpNcduiLw0B44Ue3
0sDYW8DARVMnjsn7po0VofeP644ap0MIY/W8a3x+2+2YX3izpqsGNvzTWmBAU983
+Hn5mzBCncMVE9mBLWgv9ydTLQcBPZyqbmbclZ0AaTriP1fsGw5YZiFIp7ABsqpi
lc05kK439HFRD1HzU4hEhGc8H8u7rPYgUZvaYazAdiIHm4Cpty5HK6tMzAwFG7jY
N9b1IVR9NC7J/rVqxafkhJxTguL8Meil5BHFJk1iagg2HoT7Z4WBIoyhnfv41ZiZ
JMdq3YtEnuNXyyeV1VD1qL4TVW3SH3my2vN7g4IMvC3KCFwlIPZPGaJPRNSO56S2
z0fdEqgKZMVw7FCv8V6f9lwxUzCz/yUceEHQwAS9MaRsfhNHBGRQ9rAq3pWk5DCf
Vb+0aEqbbH3JaB7mBXWRtJE/6jtAApDAMe8ou169UZsDMdvsSp0lBtkPF54w7o8E
xe2QpyyvhbhJ4Z0p5uQ6AViunA3M0qprCT+TFeGhcoAtkFEqDlgXwh5cT32WwsYt
1b2aGYS9khCnx7ku25bF83chI1M72AeExdLwhgL3JIOuAsX52gZHcgRqWV5rDXc4
QSXtExjmpgTo1xwvcxj5u393MdayQeG7SK6qf6p3/Z5GdYzq6UPsGlcbquGP4AA7
6K4jDkcXlz07UfGvlZEcFz9fK2H546DZL7I3vxtczFE34AtL9sCH5xj1g9fThAvk
QZVUhRzFk1Q9aXeuljL87M+CfX/oXNrUcrnHlrbLirxhWnNNtlFRd0yNLHpEjpVK
iiWL9839B4jntmb5BlpggdyuPbCBmUvYJ+8dPXIK09ol53TxivYZar3k1dkmtH5/
Zwae/U/mlr6d8PXRPrdHDKFg63Az8w0XDBIVgb3T93MJFg3/kBBRtYvKzUQrkMDF
fH8BOBf477mEZj3LJmV6bRicP5ibOqXZtl8c5ktcW2qhm1dNBkNIDKtOF8EyYy1v
BxEqKlyeMplVlWPGrrV+arlT9uLGD7pT4tWmzdiW4w0OnV8y8/tst9ZPfjd/ngDW
Ql0gLOx1SClnXfAT9cSrJJl5jkvqSdczJyXxzaTvwPbyJYB5B0hhm/06hU3dO7h/
ONRAJQTm8bxdF/Jpanf/3MaGMfV84Y6am8/2fwR5TCiACmoEra9QpfSELyYa5g0/
Kf9Pi1QG88Qkx2r6AAFEVCsPLch3sxNzZrc8n6CTSF+XFgEQRjDPvKobw2dcNCYs
1o+e3lJihMKaiJgFnUIzSdjznQFyhClzgadmjg9aBOHrf/KfD07Z7QFTMo2+fG6L
ZwVcd+yTlgjM+gyOJeaFlH7sdN8/rJ6gBwJSMbw1JPxcfO3mMOdl0n2hO7qU3YRD
uKvQoUNIjOoOlXAHzngDHcnXVgw0t4EQnQ18xGFx8kHkm28v1RW45VriX/fwkq/A
XH3f0jGTpXUe03sHMLlyhxonU8AZku/oLIgzXqZheDzI4dlqHtxftx8LQMAnIgtt
NBXYxlEjqTfNapgR2Gao+W0u4iZQLfxgQ9GYRKUZZMR+dHgwqWcmU1Gq/m/aQ+vN
FT8+Wljbq5LUfi22jJj4OPaNEIzfHuhaFAbZGsecHFAX2uzzB/oOGwAoYWcp5qFF
JVhojl9qx3nOFhE4f/LSmFdhNQjAz08P/geI8WCpUFRkLxJ/xvjSVd8/NjPcbwSr
Tfg6MekZQa0vSVAEqLzwIPv16JA2L3o6X64jJBeGWiq2geljDDebAfjQH+QTUigT
yKw0F1h7q1v+hMh8RV0tSQHsumBvlBTfjG5F3BCydfYOPzrDiJiLKh4gfGC86TSH
xa1I/7pSd/bhjZoPyMBMxTEx4T1viKNkVSF1q863kgUH5uy5AqBpgWJYlbS55w0W
RXCXcVmHlmzcPCoKt7Xe+rr6eCBUOgux2AnwfpH+/7apWVtYRpGRqQYtOGCKB3UU
b5nCtX1Rk+5rpRINKriTzr3mLqzAeMTDrzqOGqEZmiNGDFMLBX5PvQKIWHFI4exG
zMwbY8b5nYX8FskwAuetGQsPRK5cp8NxpfTOFelthO9VGxRFPntRTg7BohbBH5Iu
ktQz6gfT1K22lYUH1dN7TKzLi1QciGlb6BKTdHbko89kfazV1DLvzsNecday2ULz
bx7Y0kprB0HN2eqAjtDFpqRHkEW0qjZ01XoAXVP1Z74YQ/vu0gXa3yNSHxaxWwTr
fTS2963j2ByrTAKiD59rFWubw9I7UqovbwaaNyG32GzzhJEtH3H4A7d/Sc50ENwa
w5wYVl1uQrgQZXQZy+xZ83Tuzb8AX+TNeZYWHifsAo9jryldhLU8PqgHpUVvOn1T
vQfNI1cqzb1u8BYVa16s1JY2rmJmM50h8Ni9UCcfl+6jZONZm226C2mFQgxkmgBE
h9Om5069zpmTfEFgEdekMvDGFOe00j/N2zmzV8msvG8j5RLEnISXA1hh+P/H17kV
IqJfczJ1NUSgRz6DxzxtqqFUyocIURJ+GoqLcRPwos9ophmcoh36o7vFyPgfsLTy
E5ZbLYxw+D0qqbT9OWlylig/avMnhLLMsV4CKwcK2eRSrgLjyp2dp1NghsgVnANL
W77Ar7keEp64Lha6646/HiLVrTojJyCg4ioHVTRFwL5wOlxP/qKTNE8i8UqL5dPT
jZo6+Qk1TC6asYuApmHWtCy8HbHzCDMvsvfHPLRfms57nue3VyASBO1bVPEzZSz6
oYwuu+ritEcEc8fvm9U7EZ1BZ2rSsE0AnEs+nY/R0OEmWZH5O42f4rnZxvMjdxo4
r/A/CsH65MHlDNhJoaeqwFAfG9clQHmUlnxxTQMI0/C0Ocmi5h8OXBPuuAlQaaKt
9qbW9UzBCzNP1yL1WFlmYjCloKlXk4MjUl2+X5Od18IA0ikn1c9IJJWXLGp/Z1mD
D/b4TdhuQwQFMWle/u2d6AH/blaUERGaCoCh3ucUQfI8rKMRZigo7YZsktneT6Xo
IcZBb1NiWA9/sQDf7XucugHVn3jPDequO/N/ZxNKFovLvHKLIQ8KqtHjK4p24Laj
KmXf1dbWdT8rpq8zFBIHcZRMEdvufJbiZ02LBAinyM+28rPRNF2cKitAvamQJ6eN
hy3xn6xDNlJKe3HOsJCr5oEPEISCf6tOUHlnpu6xoZhv9crBIiIG051HyAsgtJTO
b5i3zUMEzBiVtvKacnUpkcR9kugV64k0yhkbbwhyG4HgktLSlFJa+RuUfzTvmNOI
SEvzepf0urvow/hQA5BVsFo4++b8/Zl+0m9jD3vdgcO0b+fXrQtR7y+5ZbxpsOZy
pqK2Gb8HlnUgPSLdjllDIZnWMqF1aBncK2rnGdDdYiU82BvD9bW29t0yIsGnA9ef
yZDTJMueFnm1aE/g/MrwWu3MCOLHz2pTUZhIg4xwC2+fU83GWZbcJeAEn5cSc7la
8y7QOtrVqQeWksw0s7EvspN9Gh9hug8eENvx5PIJt+s81LfQIEzWPrxoTdO1om7e
nkOAtxa/MKU7/gd1aBXGVl4c00K279AoJQvvSrhcoTOdDgxMtQ9w0ZMle3dq1qJN
gY1oS7AwKSqpu3fZZCV5A+u8taRKx5muf8FP2Gju++aB2bpw0v07YhQLcbrzf8Jc
DzSld/35/q+NdzSfkq59US07UXJCKvEvDCNJRy3i1Gama5yTeXfc4EStlfmi81uS
SiFOHBQ7mMO9/C29gMa+AljYyBwwIwz2z6h5MRx8UZdGr2cWDr++Mk0KezWrp0IN
EsgzA2oB51SJcYDnibQbEs+qfe5gtAFMH44dHrMd7ctNg+ses9kcJhjJZv3n1rgk
ek/Gt20eRU7O1g3Fl0AF5lvJvN+GqUyZ7rdKqCo0ZTt4dhzcoqRW3IsoUGGb/g1E
aeQ3tDIRfznWwiaSVjovSLQ6sJln4grq98BdV3p2/waP4dklwiYXtCQAuWnkf7Gj
VLOSqT0iFh+nLaHl3/oeZKIJ7aobAhM6/FdhxsP7SDK12tubggIh+A1gAcfru5Rd
W+iG4RiWG2lfcI4/LtdCP5CCMvnjLoGnpi7kNRUVRE4HwSVcfyxJkCgDwgJIGxKO
BFFScMJlnfY9DtKZL66dTZUbfzBxFfxYDBt6zUOecrOoIoZ+N61zOzymnaOyU0iB
cFk2yuGRP57uH1OuR+E2was8RMv+Nhk3cMHdtQFulxRX/PLwb3bPrQfuq4xoQjfK
kVZkvSgnzL9DVLA8AdlQ61ET8WeX/Uh02Kt68czPYyfFZsD+XmejeScrLg90azGp
Rwh2xNeWd/MNL06NlzpKHY+P7+4lGemQyTl3tS1Zioutf7tdQySOQVRq6G1aH7gd
2kvg9Vke9J5+EKZj8JrgjIyFkrZ+BVFYxSvxHoWUj9vu/+s8r0MIRFoIBrPmv5OJ
8SjYn5zAPMTfWvilQ6BMjywyHykdfz9CZIL6BjHgtv9E/g3iYAeAsRLladQhmTG3
JucwtV++p0jCoP5LqVrv1gx5V+io44k08ovfUwXKpkRKV6S/t7DEAptX059mG+j+
S2pFVccLuBuYVGe2oHBSW2R0bTElxopLfnkMzH5TYjMiXXAiW5IstRpJS9TD4I7M
f/tDhoCabP5k30R93yVqw1F2D6GhMtSbMBIE96mr6KIaor4E1OstHnpq6NEea8qQ
tTuY/i/6CCCw1Rt/mYTPnrTwZg3qeh6ak516PkkfkpATn9lGNE7Jatvt7b67Hjkr
EZIDvXWE5JSJigkvXeUbb9TizXau/t3CM4p4Gz+MSMcvSCaVXcUQPnDM3ULGQXp9
3m+ldH/+SDitUcir2fFtTn/uAx0fej7OkccScqCS/baqtPqN0KVk12mmYjW9in8Y
K84qhO9oneDOmVHlbddniRMWh972ACrsLzt+s16x9g99t3BKgwTPDj+iZitd4cZv
MpdcTSr8UNTKGWTMLcAo++Z8cN46kf8tFUAxZlP9bEBxW1uVISiD+FqHhJaTDCAX
2phe+JxT+NZwaHP8KL1tN3scTpzXhalEtvzJyszmNQ5vC6rKobsEZy9OD6CjPBTr
Qt0rHDhDeExITvvkjsA1lDT0N8Q069q79cCFhnSlp8DZGqDSupc2KZIpEoKqn2eU
KbGdqYmm2t9Uz8AIhhXw6uHGJv00xDDX3RkbypSrwNpR3XBdUa4ZGBzlBXhA4Xui
O8dWrZXoxgLqK0vWAIiT0k9ZpO2UZaWIFWCG1rG4wZZCJia0mh+8qC6jezzeJAzr
QFx5hJyUvV0/RKobcLLdo0r/daXhKAQ5f6z8WavPlV60C1jMNEmbsKLn1IQcEYcU
3i0/BGsr33cieTa8Sm6ROwCqNeZbngqN4FL44XHY0IoH+f25ATEBWyl4PjZdT2jk
SkcD/vc1KVcqfDTp4OPYDSGM8xk6jzG3RN6F+S/w9XbnuduXjZDAAgHrV7w0t/0i
gPZP3ZF3S5eIyMfLnl0GX1U1tiWw36btLANHf+H+crs6k8I8usfFH28REHNG80Ei
9oYII86sjPhpI6Pt3vTPT7A6naq8KA75JPisDZiwiOO9nAS2UBoqaZSwS6/V6g2M
Dkr1G3G5Ok9pAcf8593yeyZ8SRtkt9aCF0J16ZsYu0mGB9ZTPBuDqdOoUW8fN2/Y
oRa6C6yYx5bl3CUPYP8RP5kU6OXyhb603svtyCz8xR0PlkaNPBNnCzxfDOOLZKtz
U6NCx/fsda/m+sxKC3gKVtq/yGFAkwIIyNo9PxFQIm/8oqXiX4umsxBzQ3TZnT3B
zpiGiv8VBE7N9pVoJiTG01junQ5qHEh9yc6elX6zEMdUr9XhBxpER2qgXBHNoA9Z
r0TlAPPrI9zoSKthSGDm6r/POBi3FrcBGxQfyJA9TSjinEnXPEoJWOIwDX1ZoCNa
xtqhO+5v1yZU0m86kBUSoBzNQuYejQl0ShsaiZXapZM49MWXjiVyWcBx6V+FqAQY
tblIvVDglG3j2HEV5U2rjFGh1ecgQfRuOnHDqR7g2xP/dhUCTONDc7LNgo8cnnd/
my7Q0wrKUKZqMZa308U/SkWPSk0z9B08CWcaBXbbRSSUzVKdSq3YwEV3ERT5R4UW
3ZeMV+nXsGNr93abrfEACY9kZp4aOGh3m5mia37wCYW5qh8obpL1V0wTSox/PDDf
dlIpkAR82WWe1h1MkQpqCi3QMRjBH0/ynKScFDQ4C3p1ByZiFtl0nTs7I/7FxDgw
/3MYA0UvegzZIA9+jTfNTJY/xGguwb23SLbspUMy47v2X39sBJMSIWPIwc5LJXWM
l0mIYS20D36sGQ5oySnFa/K4+irl1ldlrhjz5sVVT+k77XBedYKXm0D6FcQ6dcgx
25Vb3eyYI6E3xd7yjsiMiSEvbLvJG7XU0lHzJkPTs2kNHZE+ADq5i+RAueKl5G69
yvgH9TQFLNAXAbwZMOw0cs2dwcHIvFVP57LPXdi8qoCWvOBZNr0sC9JhodV0wJOb
j9K7hnE8ttVTZuuKYm+kMeGbiJTj7ZcO0OBHAyoF9HpkifEkcL/IsGtEwrrJrTTk
Hvhe+56RL8IFOqBxg2CM1KORO9Jdhkj+wTTio+hIX5voeg8TFv8DLv33JzPeQjw/
QMm4WswawcaLFFKQCSFFgV96o1HLMYYaLk9GLt4fjWdHl7VTJaJSu2QnADgbeD7T
vmReT9EdSlpSIE4z8IVLAK81pzCJiE6nL4PbQaH16hDK27f80XMhLS7Yqxi3FLs5
8n5BLOWY4Pxz1zpFDCNB3Dla9JfTBiaByySQrsN89HgMlUf4yPJy3UYYeEY3tR+Z
yiMANcT7VXgxvSNn0wKCipSnJDt0lvkkrYWOfMB8yroQ9dMuPgC8tCDJ7IuVqGq2
D7TL1UPngptnuxMZhK43yfmQybJ6CCP8zJ8QJPZzIF+DmUnryGZgpvSbBrlwSlC2
Xog9C7FGFxM58yz++J18skOrBNTyGWd3+Vkc7Gz2sEHRMoJ3/ib4EvT5c8bGvNq1
Oi/OCg5XSyJiYfYW8dQuUeySAr7MuJKo8r2vmKEpmUI77X+3KJU7cTtid+ul/qYT
sBfIiDUgVE6+JIdCkXWy8Z0JbI96OEGjP8BsR3ozU9agAv7IQ9Y0PWDjKw7oRBmi
iaV4ar+LQe/L7mkscwPX/y1lr1o7FV5bHznRZUBn03qiKUlr+K2YlZHN1JcoF1P9
67sKKZs2+hNzZyEoKuV6zeRGsL6fUISiEAlV5ZUZxljDha6IR0GmlPKHZKrF4Cir
idGUxCKThYvMNTudAizm8x2YaF8zHjHtyBtB4D3GCOY05KG1fzJGW9gHzFPT+2Lk
KO2+63ydz38kOYrSvvRLtyr4e/jE4PQYgz9WK9ZnmVecK3dmYn/jM1QLomYcaTh7
gVWE4e5VQ1RDv7MSFSZ+UmgH8W8r1wh/9iqXYUW+0aX6Xwqv5d74m4L52wyXoEow
f0hJBjkf1laKI4rviJFMs6Hdhdr57W3PyiDughmQAF5BP3dcvVaZtEtLnz+ymyh9
hbTkBOu/c6QD+u5PlSn/h3UMHwLatnDqn/4QvlH5+9aRiILWrdP2mt26vKJj7pht
B5xLzVe7WUmBMFb2h3OmtaTMoHtJMwx5FlPsRHg6fBPb6dUX8jXPWuF7h5MlvXVF
zqZ2XBwA+50FaLw07pLoWr6FXr/wBLNXN83nGacGtxWrDo/MJft6/g36DvV7BVfO
vROrSh2dmpivxn20KD3FOxvNomrKvBbKeYA+gYtFxXJly1rX/4lBRSunPjtA8CfD
KBD8d+Gpr9SzARvCbviQsN2MxXmB1LnlMLZztzuQbugMq27OtGZ4j7e3l5z/PZXs
rAmZHq34p+FQYjkjng0eE+ZxIff5yR4lEAQbGfGFIUZAEqU1a/y1NWwxu0NKs7q6
D57CcELPd8erw9oicHZCwkKz01YWo/AIs5A7u8L1hcFAENaiAUi+poj7/6xYhszk
UIMUZ2Mlbp+zQsVxfs2rV7hMpXuPeTNQqi8p73C8/7qm/HSpLD3tf6nkMGE2wrn0
63vwYoWd0BP/rkHkje5yndPyDoP78PbhX9AEukwBr8RQgK+eoDyNAbVNttvKQ1ze
iMroONASLZm9iz6KUB+2UTrXGyY6JQ+6zSM/6/NyGYnUOGHHyh2Dmo9Kvb6ml/69
xP6q8Cu1CPi4+KQILkIN2veFrQREwEdxAsygZX3jCSxfCIVJIIisC6U9+mzah8fE
PBrYcN7LmAkjuqO8I1efF8i7No6CrQ3v7qQxeHv9+MBghwZppF3h7eLMh/pa7bQu
gSVU2gXKZLUtF4tJmO9qimVeGsAS8xlCuuu4zSyGj57BLGrZ8SbM6qNr4job4U9d
F/0nGlq0ABJy4J4GH64rUZ+zKDnaz6YIsiAbAl2Vz9fDUweZpWKql/DENUpI8PNZ
39rmvzFPYl/d6WzvZJzQI9FxosvKMlQFljc3kRR3RpfCOwqyqO9i+pA47putyXKN
5DrFNATmxZFzKXGQroXNZGz+bOTtGgP8Z0grNb9QPk8hW8rvq889Y8QsxKYNKg4n
Ik0MBsJEbvlZglW/QyZnaFnF+3FHJ2OYNidMSjxF/yuN5uyFRcMKTuw02/uaLyZt
MOUgGQI1Sj55YlnzQ0plcqdQqpI3MyikboSTkd2BVS9z6EaGtW6eERblxFzokG9Q
E0WHktUFJ1zWjdfsGAtDt0mz/IcHWzju5wUyJVpcPZOT8zS7/lppFAfPCP4mRBIt
3ODq9rebswPCKzWkyD5LVXJBBOdBxL5ZnbZ19O3lXKUQiunXaoGcd04IAtPgf35e
dp26rDJrLdw7zo6Vz1SxZcAtz/f1lsf21XCPzuqDjYXfHkNM3FbEI9POLEgBar3n
RwhK20J1y/X5kZd5DYpodhdMACaCwJxlvWEyEyC/grZGrM6NqCYGe++x3r5PAj2g
FWcryUZgIPeINWTvP/aRqGt5bAoDc+W8GIusB8n3Oja7H9tVXtfmYoCQGjuW6LBk
9jYiipAafXCnNkfs3LYWEilMQRobyiz37oIkeSyKQayXnROVz2V9Beq8DASnwBxP
l3RTdjLjS7fGDApNcf0NUeg3s/PWnob5uYEzRsaTJ2jhoPadcbl0zIQYVJ7otPo1
5ddldvk3vLsIwr+UGcZUEX+KPXcOAkLH9vqYbLI1EXi1Nl/QpBfwohpTBVZOPJrq
isGkCh5zk36EsD/dNQyT3PxQTsWo2XSaIpJNj7jbErZYPiH2K/TMLI3c1X6NEcXL
Eh7OBJR8gJbDl7gz6VO9meJWwouEh3NvPG6nrM8hEVu5UMXmPA+Q8LU5pNLl0ecO
hTZM/DtNyHEfjmNEeH+SV61JJD4MSk1EIfxT8/E4j6x+Tyb06WbXrGoSnhNP6v2I
L++Ypp975SXrx/e5f60QcsLm9PuKamxxTCetVoZZr1FgA9g6bsmPFgXc3feyspUK
8sns0zDLIQe52WMnOabTf3cRabVQzbaGDmZD2VICki+0Ysd5lvNDRPwPN7ShmhPh
oxiAs8s4pllr7W/rPoLlPOwnQ1HSW5jVtCkjCx0LQ7MPWTpQ+Y3hywzK20N7QUhm
lthIPCIBcDxL8xDO8y8BjMVL24WoAiM2YZ7apJ9g0VLZzQdlpyOePwHXZX/Fr9FJ
0VWIYtMope9GhBzYqeZBMYYcvYOfzNun+E1dFMzYPlNO1B4x1Rv4OJ1b3S+SPvk8
4UgvYZGC1wy+77Sw3C10BLbsBbe/sPRU6ZOHx6Yr8NyJz1zUpfPN8V4QX2PVb0CA
5PCX69EeKm1hhsEgeQzUA3Sqbmkl0OoeEbSeT5IXCJnl8KESHOhuW2bu+Tu1KPj+
+xdc0/chsmz8Nw1HoTe7ASTgPoJ2VHFPo+TKwRQZszNGFTsl3JAoo/f8IQeAlh3b
+guEPG+b1A5LPurK3NYeILaf929f0J76AZwiTbcw3qgRYKOA3/7ZnYgrTV69QPH/
hXY7gFgFtuMb6bRM3lx4DIFhGdhpwIvC8hwHH3w8ZBoh/tgtkxI2eZVA7LNtYRSv
aZ309X/gdrEfIRBCkFUesga+83+/ZMGV/hQ+h8kb0M7rSO3rQxxmWbd+ICaPP8PV
+cT2A6vFgkV2hkDVqFbWqobJ4znZXnF3DxfxnLACXldYQap83fm9XnytXEIUnhQI
qCYzNcN3CFeTJO+orzX6jrMLgzBQSs+pH0FY6OUl/4xNyhdrfYPet004dqTrqVcN
GgjBXt1SQHmfMwFLzB7SaE2a65V9web7d8b7o+R3pz8MQ+YydebSpLIWv7ytZbSu
ihvfQx4CX+48HmqeiW2ccxOSbiVDJ6cWRtWZLmGdydyXNFHnlUo6VreVIcD3gxh7
MU71NZNwN51Vd/z6YuBbeu2cwVA34XTAZ2+ZL4qzXXpL4k5u8psUQvbacXAmPHa+
lSAfAKgvdLWqy346fSkDUWXAfC2eehr0e3ZNkQjKsz2viHsQf9JPRXYQwwG9sTxo
+aIX0LM4Uy87Kd8xQavZwjYDfDBQRHx7HiMhakgEgIHDMRvRTHlpvVix0nHyBqbC
vYHX2Pw8a/duJ8R2/CqhxYbT2e2q/Um9eDaDvp5T+hUcv9Jjj4lTzX1EccX4PnWm
hESvvr7jJqLnf5oz8qhYyUfzriy3PRxCSm6TNIPmRJG8d6Dy/RLCQJcOHmMahbFb
//fv8JdGI5ni6WePKU9oEolCk0w9AqJEQZ/Y05YxngquHxR6hJzXPgmtYrfKeFVx
wbQAnz8r25Z3awgwAlvMmEyYoU6Ql9YEFyqWF0n/PGiL6hToYPqIfl1j2QMGpLqG
rofnOCMpS5nN+s/A3+MghewysPrKoW8zBTZjvax59Wk0WeqxPjE/C4X97vXQe41o
2XQpwtFge/WS6Y6bsr/XWkHphXyrnUl5cSsaMK9JLI7M8FwHXYT6vDBtJk38Rx1G
knOm9VPRpNLnkjgCGYLgYiEmTBRsPINJ1+vgOqSfn4NKJFFVu4OtXJfdYWYY1isO
y3YkMQpo5B0puzkx2ShrFKXIU3vktzw/AjcxM93wCyspbQOvyb04TC17+E3BcmR3
6UKP6gOciwZOTUnSJ48yW4pTG94TiMbW1avHSodF8BSTN6aGsA9ZBlaBp6gIHzFK
yGgu7ywxBZfOwfcXfC/FG9xwvyhMVyp/6PpknvDPqxH+h9Wbk4mHfsgU0ATdQ12r
snce9mfVYCX5NTO/8mluncaDbnsEs1R0DTkIJcDojUCDIhhY6fu6nFgeoMboZzM5
hvipC5uZxIo7ajPWaMMm8l2h6jrPu2FNrwXEMsOuj1yveF7nLMRgQAG9I3pi/LOw
IP8uSafOpII9qwpAMfe0414hx9Hx6r7IEPD32xXE3qSDpkmXJsUbKdMP/nUt5uKs
vL03qJoFLZ/Tz5qALmjkXicyo++ugwkNtcyyrPeeBa2kj81d6QHvib+Aq+M/u+++
jE3fc9Zj4KWeEYF9ZS6UWAg6HJ9mqLryWainj6093a1+wqLkrNZjTqHP3fMLT006
X910DlrPCsF4ly2fdKAlAOnsuKH7MfA4G+9KApRED+ILpzZFmX3e8zCA57UFop7i
XvqhdFeYGSBkjOxpH2m+h5Os00/ZzrCddTPjMU9UVoPrq4hYs2eFHaoen2UzlBy2
xMLhuBjNybq319E42ZJ5LF0XmPJs8o+Eau3PI0qT053cxhzhiZfi/23rlKR6/uIv
4Aukt8AJ6eLuKjk6nL7oCE//qBakIpoaYvhAVBfZ+ntD9WrQ92Ul5Utbrl+wAJEM
/XmxkROBWLgVVUbSESet07F3UHzzy2NKkdfnkamkGwW/4h4YxLvoCS0d+ze/45Nn
MtnlaKa6J5tXybfpQNof6bnkJSrqz+7xGEHkj/3vZzxt2ckUlIghwO0hym75jV/j
vm0MHJHSPyq0cGUhBi9cwhZ5xz+uD5aEpat5Fw4udQZ0jgaCquXBFlFDmF+B5N62
6no+eK6/SoGbxdsvdIwHUXpig1FXoe2ygy/YsX84s/P21oCg1KgGnHh872pj+pqW
GOLfXB+bWvuXUXL0Li+VanjBiC1Ux9ddkUaV4mDJWRsI2EAZSRUM+rtz7qQtGypa
EhDCuIGm3kdoDxZuKxaFiqK9ekQLbm6dHEa/XIyCzARKAbaKajTsu+fcnVYln9PX
GTE2QdfKjHU5uRGegLcP1Fm1rsV8UOYaU7WloysD2KJx+9B8mHBKt2jULdxm6wIf
ClbSfyArgq6Q1XZUegjREqAWupYHRd2S4/EltrG9Lg7d44XFNsJvfIrXRFpC9DVC
DrHZ7/VplxiJNvT4Nb2xJ5sPSD4DH6gLYAUPwsic//Xr+ooUsdTgh2+oJZgBHbsT
zDW15WkTD4lQX8aiLga7iTyUPqN2Y4XWhzYfsBhlTy2lUNNBPLrsptk5EcUX1sni
5N1G3X4hVt3ssAiAi8Xjh9Z7KpQdGUQP2OGeeIoGrXzkuCoGqzWj92lDmn7wW7qm
lLz83u3AWw9F6yQhf53Ivv1IX8ZNYju9KUeJEpudFNZWLs/Yf4fX4+k69CjufA6L
8qW+fMEfTnNSAWQ8f7SZpMzBE1QRuDAOyI4EKdohze11GKelWP6ftIH1H9/e1bov
+Lu5clx2XXNSH6maFkvk64/XTaDjlNgDx3AJJDpcq/goQxVhnqu4wldiSK525Nzn
paFxMuoa/DjYXlOu4W0GfHk4RmX4JlBf5EqmWhyAC3CAvfH4/vpuTOWoCVZ+E2Hy
RckUUNpS26cJepQz1e2Y8GPTsyTxYOZQw9Fhh98zTmjTG8ao57gimt2rLuAjQLDA
a7SriBZsyDxnmZ+y1mn2Xn4sqT9Nr1YB3mz8YG56ZyWhLFAh0YzkwXwiYrXQe3cx
X9Nhy/iirHs3Dlk8xIW3A0NdUifgKia11XET8r/k2feDFyTfZBY5jwwXtgiS9fhC
UOwIwRou9Qbd4e89LrQnrDF8ayX7YqDHpsyDgscv4B8abCtcwWLR5IHqv4bb69L2
KSe6iVTSwxMh0VLWK6nNUfWFrbHW6kdwvQENR5Qx3wbAeiBHygT6bz+PuzhkSLe3
qE0gZBtG4Xtt133NNSxfDk2I3271edyyrSUnVjSkUtY3Ksrr85wV0Gm9JQoVTAr3
Twjin5rwiYdqTkiJBUh4oo2jzpPFYv3yItPzGOqEasM5Cwe8WGRgm00q73FWJ8yi
6IlFEgSSY/C7Okp7VzFFT1YrfCWF8M9YXRNKX7oow6m2iAjl9EQqAOgN9Q2HCJO1
WTx+mEgNRSL+GMIFFbHntuyHQL28j+Uz4GexRiao4c+62rlLTVhLQ/Y1Dth7FfIs
Dh3LxQbDGHt+XvswxEZPoPEzxvQp3TDH0pAGa8a5k9+P43E1s2BAzPPvAnBWZcbt
XuX7eq6qNMrRDcOMoFTm+6Js6ajZgZxRTRl/9ABmjU4hwiFlDldnYoqRc7/dVp59
ga2ffT25bcnaDjmrIeICzav7DdqH40f0E1oYYreBpC/9TYh39PLzDIn1C/Qusz+J
dvMDJ+4LtvWmWfzaixqlQteR3Ki/HuIrGMcl89D6ZwIzjXj+KrM1Shi/7WHy+OAL
SZ78XW9bAPBevgzSlVTIoKFOSUPU6D3C/W4q6I7YUfU07va9mOVoCqt+2KLbWtU1
iGBdloHqKCFf6h2QfvFpZFc4aZIBrW77YHrUF8nADh1EY+8d+5uNYYYt8io14NV0
H3FY9y8imaCiZRyAmbcPpiCc8V+yaVVbSuotVExuAdep+xDAQv5clG2ut02o+X9H
BLhSAHG/NeuRvvqbSMulqQtw/lNTsTinVeWLtk4l8eJ50wZfF04TcohQEluwqTE3
HH0zhz0efjMXsjs63OLdr2X4IUlccmg1K1J/6vqAyut0H9vC/wY1s328QXtYjX3P
uZN3ePR/U+iXBDFeRAL6GpH7j4VWzmFXlqRNhUV9XdPc1UKZ/6ag1Ul3qRW+WwDD
e+L0VaGKYQv1K9bSPz6oGK7x4a7ccRsKz7ZSdOWq0P478NzkCBvn3Z5ZBgUZzud0
EggqxE1N2sZ25+ddWGfe/TED7mDbBd83/3pKtGZo6fiGCze5+N5FCAONXJs9Iv4a
6wpjgu/v2SdFvIS6kBNKXbRpRtWCQurjKD2tiV3m+7z1tK404cDQ5d1ltznKQ9/G
MVSBoD++I6GkS0dExrQ6DMOeHgh6ZW6ILdqhFjhBgtNuKFMZAdwEeHmkS1Xr5RCd
S5Dvy9lAK2x+okthS0cPshFvUN1aCZG4DEphFBU0VnPIgpxn7WtIQjp0U58wyaSC
kBABSXEo0W7XVSxRaWwCC6iY/e/xTSJ7MaaKJQKjytXZgSBNHqUsaftuS6h7bCvD
aBwpdK+i2OE1H2nMJ3S7RGXpZmDLZcMwKeO7BeT2a10Kz8CoRKbfXA1uF0v7+dAO
G/4WordGlrPUwkrt/C0QpqDuUUcR32TGijLn4ybSLNlpAXGuqyu5/LmFOsG/RLiN
DHhYD1RosOysDLWCZ5ibtCfeekNZRc+sAxfn/g+YEF+jQnrfavdtuXR+d4xYXpuF
f4N4qO9EOp91qQBoW+XHj3MDGy9YLtP+9jaTeh1KvisuuO23/93DfKuBNT6F0uAW
D45oSaFwX/QcPES5RMMK785e9b4up2sdz1WloauOJfXNtwLn3p5FbnWOZ8Kno1Gv
QrkVkPEAmefz3uVEPPUmq3HEMfgCEkpvdIFEfWASQCSn7FsaNLdVXFfuf7kEnXym
AenAdLCgo9s6LfEd5h87qC/QrAoxKL4izuG5VNFH82Cfu9q53BwD1mS4PElCnT9U
D/igs07UPqc0ZyAZhKg61EqD3w/GyjCo0HiY4WvoHKOp6ylsQPn93/TcIzJzCvfZ
jEmzqcoAEJk/e76wgkZ/7tIPYIyuv5hG4GvI/wBKXQqARewhCRjOY3JIWIYyeAjA
y0Zf6zXj+JF8UBa77UL5Kyy2n8uAjZqjY3FARO5AEqlZqAdY2w+NGVFRA4NBRIHW
1eJjcxcHiMZd2ubNDU87ty9W7UF7AVOG4yWA+JLe2/85Ofxsutt4tkUashYGoxLR
TKUWXRYWvnlGDF6gWLI/fc06aplzgY0KtGkXz7W07m9+I5m38VCoeQLASz/v5beo
RnR8TOf0K36umgNQFhH6b+MqmzTCLUzz7X9buOwg766YA17qKgS/dLr1efF2K7al
ndTbsnXx8HUYN92fumy9KNFEZL4mPfkP5cOjxN2weXHXA/2TGcadsfSUr23fUEL1
Jq6dk3DoZmV5Cyz+APQWk6Ljl0tGWjeMaVvfjGosSwkW9G0gQsSQ3cwll60ql1c6
3gzPLcsGnMoaYssB56RqJ0q7Iuz77OT/NnC/F8aIFIHWunrUDDqUlJXnrNgkcvwi
+bVogtihDas3zRCCHCFyj9IqpsZsiYGA1ZzDqzsGA9wqv6ePEQbv/eS76+6RpOmH
T0lBII+0cx/DwCja1lreZY3ECpFRQc8FbntyE1xu2HYz7f9rIH9MA+94IDDoL4Oj
DehjWAzonyLkFDdgIrn9FzP8gXT2TERzbsRDGdvKBS1Qzcw3hsBs+xzTHJx71X5e
B7h7jzyacnXm97dMecI1XZxWWY9EYT4eUt3PzmE+XVc8/9KHxwRIsRCzoMbA9YsO
yPPUIrBNH/i8sRo/it5cP2NV+Cx24me9KkJp7oHmvzWrFxn0De0JnF0C6OzhUna0
CNVxBfnRD/6hBQMncyKb6eqa1zTPbRGN+06zzYM0IXJFQT7/K1IyBg1iroK+Cn5o
/pMgXZ9Iuw4XPKSeJzTBTZzVzsXUgHou1I/l7bMSoYFq4O6acK3Z9RdiuMU+MMUz
swb5wL4AsWhH+iB2mFmPKf385UEz/k1aVM+t+KzTDH1PQKP0qil9I1pN9hG9R+IW
7KvBja0W3VBdVUxuJOJZ3zFuwZKRroOlt+n+80vNF3nItuzex6Yg79fcSDt5KA/P
s0IxPxMyAUOfMIEPYvSE2WywLfeXpJhQz34M6n7js4c/SovxLbRSsIo5NtPtC+a0
yP+9F4uyLzetnnvMEkgPGM827a/gC2K3HEooocFz4UQbNSxg+SIvc/HzDDBxZaqy
8WCjLykV0mfe+BUX9rlht5ufarvKCjtVPrygUWTrR1uk5qykO3EVlkiDgY43oF0r
njkGfbFgNAQELHI37nElyDV7gByRjiISQ7ppsrwC6wFhdU+MIxhtAJWwt9Gy79jW
i0LWwtQdW07kf5GW/A94kbg6HL3d8fq9dfPeEnrkgs7pr9YuTbEIUYJGJACptOO/
eZaLKm7Cnx4UAtVO7OEI1OIPfDEMochDHyAbEO7VWzwmqAn2xFPypR9gu9cSnIio
I2OSBXmhzHBAnQO/uzRAvYK3d56arXxgaACSkYmWGqVnkM8wp5eBUvRoz2U14MHj
Tjb5usFwVeWZioR8JQ6kPA1w6qHw0SJXiKePITh4CHWvR4Us9scVA1WsYuMMbnTm
RIvtXxWDkOSj76SovFDTQSL4uHSRojBSIFUrX14FtmfnMxM75npI8UoHlaQmDQRe
z2TrwAMvnfvZqyTcJoTJIYamDBCKB3V/V13oxcdEBmCyiKLKgk8UqBPOgTTpk6wl
VSNhuNs4MFVSLne9nig016liefFDMkRZuoPB5knNPYTdnyg86cZqgOBiQUOOCPHf
MsyZ7V6250cOUNB+n7pDV8o3MK1bgFVAre4LRBHFO2dcgJEIFljUtxhQaL6CyNz+
tpdimvSL48wAU+8svg3Y3qw9wSGzOUyY0LoiEvIqlCvENUsiJaV7HHyqa/k92qAO
/U0XwHTc16/6nUESFicuP5IWb+8VabHZwpjlaCFUDqB33UJu0bSNJnD5m41tnFaK
OYvO9iUOEcVeUgadd1NJwWNCpCFaICTU6+gpjzupYQ13MTPCJQ06qgDsKl1R7rus
Q5U7lsIxWdrYFVO2AEWeUYArjYnrrF51XzCUEVrHMT0X6WoDmpE4h2DiMWyBgr9h
FYfut6bbv7YW4jO6JKg7nKkQkQ7kLLPh8jCigpFEwywPW/Uw6XnIgzfZoQHUyZ+/
WKlZaJzXs6xrd6Z2+E07CAO7ccMvM1CJFqULh94VyBRdqaG6vFtdopC/pv/cMhpK
8N9+/G5g1xGq2NraOwzG63dlt3kqgh//HcLtmlaDRnDPGuCs9JSXbrps9eTVE9Bf
jLr2vpj+JChtF7RWtbu9xi1E8UbMx7v/v9mZ4u8rhjyPw2BcBC76/rnB1eJVAfX4
qSns+RmulPPL+UfwG1mN7l4HSh/lZtFJNG9GDkw6lz6zEk9RdLVPEQaqVJBagqce
5NrcCiZKbZE6BwvsgD3hupWx1UnLfRIQgstaFEeI5wPL+dESFGP1TT0+5YFrTDo/
GaBydTtc3bWo1WotQ73/GCyiZnhzRrL0uobYlWMw23kuFDRrT95IyoUF5Ptp+w89
nLGZztkAxWULrsLODhe7Q6SjFVXDvUewLUbhB4MMiqlpgxKsstOSLNi6nHEcgdr0
u54HlVu3NC9b1bW5YI/yWvOW/gC8u4I5K84cZTDEWDB/+TT4jhfzZhlFs2g8MSRs
HOAs6gDvW0d8jj66dRuXD4RM4Zrn5P3pOD53Hm1gI23ciWW001NhSkbW44w/ZlmT
QKH5n1shOQ1LmffjVEwdG13klYQxhsEycpBweFbAsAF0ZGGNwPMx8CU2NPdp2S1F
+Ovxzd9/JkuJ9ij7dmtXaoQS2NjNUeAHiNwGWqwAa68TPlGK0mUwlebCRMWsWGm4
Gsy7sKK3WYgB06kq7Ea3pnzndDiSsdxtI3UPP7hiHo6LNtW0j1jyrhTLkN8j9Sv9
KrWrJTEadcB6198Wrl/FncMWdkXfzpCsZle8QkUaLjlKAFMBEjgczBRhBZADKHMt
WtS/NlwloQGvjS5NMiEcM/+WKQ0HueLi0ybEwfBYHyiUhcLVue4tzlc3Rr30PVA9
6ejN4m9LL3EoTOvB/zHB8GNQs+am5V9fP3x3NpIxoNTME1k8jkMSUH6hsBC3pqiJ
lGKBijwODpK9bY0LCfEqDEhLQiBjXGmzAsAkVvH6BFm8LLLfEmQ4HhQlfDDvvRyc
Kz/pfmRXgW52ax/7rKIvlWsoQ/S62/0uwwCf4iRCCmu1A0dL9bP9dpUluyXBKb3C
yf/wgURhA7ii1MnkkMkaqntyysWvHap1cNHVbAZmcedt8cpBUerto+F+PWSANSAG
EwNAhTgb9/CMeLb/UWqqiBLX8WHWP4WHhGfBVZmTNs4imSh5+IrCtpYtFlzL070C
7NM43NB4nG8dpA1vljxkFQigtX+/y+qxKYbi3FNIqIWOlJsMQgz/xyTmtSdrRkq+
c0f7YR/kF/J7NuOpyQuYnxw0kZqaFsnFy58DTxnAOnrcK7nqLkVgD/IvG9SvweN8
opl40SCIyIrbX/54fDgMcm+3i6D2Fj4TbxC+tUqqNZyMXdEgPYgob84Swu5vMeo+
OJpW8LNriZc3OdUot1mBjDXg0zlEIPSNMsuN8fDsMtKPngK5DQ6iuH9BcqsSszNN
MFx45ECG/K8Sgr+MEzwBBAwp62VVwaV1/qRTh8BfR7NLFAcfiqBVEMHVCvxW8pWP
8LuvXMO2oQdqsnnSf2deHiFybEy9S3YYu5AI3wAPiHtMzTl1ys3ckmoAWREEZgXP
g2ww11yw0x7flIWtclbTrMaZk1JMNdBgL7lk9vLrVLcjvDoVGNANMHUvcH1rqyfD
wfmyTVfyxVzuT/JrG+BFtv7k31bsWb58obrOVw8HI2JdNxt7kMrFrM+cVhPTShtT
EGKbu1tlc5U7XlpU8gkEv5hWuAPQ/pafy6PcF3ltMvZ9BvXxdjBycHXpUX7y/Qvg
Jo6BNVrL8RXRH7E1dZB8H/RAOSiVkYX+xOvcqBhof7DbheANkpFSwlqxerYxIc9t
dgkhN+/lidQV4yR+TiLnAErb+KT5b+aoV68wfxVzywlrUWEOICA70AMIqv5ixoEw
blCGmMHdOXxW0GwiSMgiZMwFkxxpghdvgx4+w6fM0EFCk2H9tGl0lxZXFHXqCirj
cLkcwFi/jW02Pdk6pzSjfH2nW6A+5w3ZjN3RVMyuW1wZJ09jhVYt8kXQSDNBJlQb
FOuft2zl0BJND8787yGKXlnkHJ3+laWD4alDKRCVKoGzadPXk9I6AQ/jDpF7hQZx
hYRTp4KFTVwkFeCDUrPijITJCm5XOn/y9vNK6q2159RMWgjdCYbRHdwsCW9AmTMu
fU8ENVTPrmDIEhwGGpLfixLcCIGqcSHFIVCPTo524rFsJ7wFQ+bBnB27ocBV8zIm
VcjNVOpK0isPExK3he+5dztCGIEpF96nXhoMvXiiLFppnm733SVCk+eZ7+TXnmjt
EZu8mrNm8HXfE7rWLHjSXfTbwiVDVM8mlpGgDZJbpBXMJsZFf72/6twf6JEQrVft
7YYxYjtQUMEvYfcHYeWDkBbUlVJa/900G99NNYiF7YpLpP+9O4Qa9o3VVEwMULn0
Rhz8Z3vIFAhzLbP5gcJYZ1gIxfVpqOoxzvUN9MjP8VTMYrRNoGHkWldDfAYkIrzJ
5S51HruZZvmFMuec0f1OFYo5mVRvKPP52Igtn83aGpMzFCJPKymLfteufNMfjofm
Yo83JoeW8moVXsI6wl6bU+mhQg/nVufAw4zAREQQM63JN5knUV0a6KbVdnMEgsj9
rKGr+1rTYC1rqDNRjcKnlJt56DGp4mOq8mMBqRAgdPqca7nr6o4sZEHmFqENZJ0z
yyVtwh1EH6pWS8E9JB/k/WzoiEXGTwmbCTYlU/x+N2h/Y4/wS4ryGucit9mBJAi6
NBQ265loGwsdwyaR1Z+hAoJ68Zz+1RmGu9E0gDckNnvSxya6diYRwQdHPh++sGQ8
elNRfThK+hqjqjIRXUr/w98NsnLuGdUnsL42uxCXC+0KaJ4rlxpg32HW99DAvsPk
pUZIiY7bzXd/8gi+ydVKCRdDQ+50iS2oL3VcoJSneh+OBeu8lsxTQx1EOYLJW6PK
20cwozmusBYCDPp8z4+WhvomU9DxZXZmh4ZoP/H4MC8XiMv1UskPodu2xpHZU92K
3C511udQLy2+HHmpcqkVtba3VOH6JsVlHf8/D2Rg7IiQfriXEpXtI2zUaQulZt7T
qzgcVaSo/buhu9scxBjK2WJ5k3x6f1J+o+hWYaLG5ojB33vwZLH4/fJirsV1VyLh
Fxu4M2vcK5hlJaF78P2z70iIxkRrdm4Y8GHb0kh+BuN4dctf2L0ThcHMoAFC5Npb
ba9e1K+GNIO3HGolD2YbOsAHcrHYTeuVy2M7r59+Bfol/Jn5bq/ezvcZIR7cFQjV
OPKOZHKBT0NtIEVq1WUCk2+hu/9OWKufpPQbf3vKDDjQ+0uY5BJzowQ+IznV0otT
5OIpihO7Yvdfg2L8P1gsW4z5nbs8hc0m8gMWH+CCHfLaoem1bFaYw/9B3gl72xyC
agSCOCy+oyvGhuzeyd532vMGtGTx1qCKgNexZtqQbypNtObQb0hBGBOjKE5JPMBG
/Hkelvi8iaYzjrGK4RASL5GiGCzat7M4JEjPyklEDd7Vjxaia6B2nDkyvcDGvOnX
EqhZuqP0i5vR2pXryOLSC9ffXoKSMT5D25sfXJbjbFTExlz4ZPfGfbpy/eokg/mA
y2JelWHVbZGvBAIafePeE72pSuG0S+NXRUHMElJB+u/Y7KfHq2DAalFEfnHdNbg8
xQaL1rukVbw7CdWoOm5c5jQD2q0C+0zg2JELYGGXe/xeVudyMzv9tBRdE8wgvmaX
cPp1a3zMTi6C+xlphrn3uUaOj6KMAqUh/PMwC8elWQ7ZEnt1eWJvEaAHcUK5q1Qs
emj3tDc7fqaRL/FuSc9KVER68FMXqGYWQys/Cgul2BKtxmUB8wyL3wcSxkG4+m/p
tmNRJunfoj549hrQo0KhVpvzFy6kmNqG8UrSvakW9eaHv1k0ekl6LTKaYIH+Qdwz
avZ27DPFgn7UESDb1CNYiG97rno9ibL78I6zamw66LG9XV7lGELbxvMXcYg+XRzz
EwG41LfTZvCXqo+py8vAp9RTeV+yr/7ZkTM0aaEvsJiXzS+TdWgHHqrkrag13hJe
dQX2QoT4UWiy4P5m/vjFlLkCiSTcP3TBrzggsAZTJSb/YycpfM8y8D/UFuRdGcGl
80B9k2yb7fbrurtO6srhpeiXAu2VZ0+f1IcJ4MSRQYQfoj0rSuCzS9ejUVrF6Mcs
bmQNKeXHLS44UgwKRXkXSz+GSZ1BBKsg50eowEukZ+jp9dl1LKc9Tzc48y9d2edf
YDJn2DazhjVx1qop+tpmUso34daMr9rxOnvUvfajQH61eWA9PAwI1oMBzcBkiWut
GZ+MB63qfj/IptDfsblHXADQnanGr707zJzXi6AXB24Ok5+Ywt3ttsiYAr+h8/Ki
X1y99BwLweO+ABTxAFY7MTvksBUGtYWgoeEfhfK+pXLGHR812RdmFX4/cRCnJyeI
/a7zVGh052Hir/Ncuq5pahUnvAWv7Nol22QIvOh6KGYt/f70ukC+7FJVKKLXAiR2
gdNA9mDDw/ew9cAQu6oJMm843oIhvXcBgNNbwTxNnXXoTlRHaV8T9K+B96ZEc8I4
SI7G6dMO/0Eu2w6ZPQDd5cYRbxkd0obIuspbmGkziY2LpbTkXvdjppyySOIvL9lS
1zNLkWk/7vEHu22UV/jrPm01lfg37eoVYfM6uZikB6o4k3KKM4+L481rBCV02w3g
kC2UwshPVr4Uw8SGEOLP0O4ejHV81sBQeQwZSKQCMuZnk20fkPege7iaEQqs2V3S
mNV/baD49eWt9C4B3RQq1DPDqENXehxrGaWwHVi1FqKcQLVHXPcTO/ugrBkNsQuu
CHYpiYf1i1yJmILOtlh5tbxaToUvsrRHrxoRDkTtt+E1DLEL72GJ7s5fg3gwR9zl
14LYqq8brN1Q3kDe4gj3mT/xpAD24OduVAJ5cXHWbZQ8mWCFGd/+DdyMDirQaXsU
AgeFrYMUdVe6hlIvQr2lRwKZfDplUAvJsvMQqmf+rLSft7y/7nPsOwQo3BgAwaop
9bs8yDIX0+moAKLHJ1Bi4xD8OtNkLuoywWT/7uRA8YineNpH8bybSTGs63NHhP/i
sz6tXKNoaZq61nbgbhWsi83rOH4IWi9LPKwlcINlUag5mN+p2i3+FbZzNagXWyGt
Fob/XHdIx1NuTlDf/MrMPGZD4Zw6GOYr1qayblUQjLwmiVhjDYJmOPHZLTmewvnp
ALiDUu8ws71QkXLejORZYszr1XRFHx+ExlrpjG2letXxuYKQc68pPfVQdKNBMZ0B
5fB+wshYCnq0LwU22rxbMdtSy9DJkrNfr3PpqIoRteSCW/tTJwGF6x0sHhMoyWIn
CJ3ocm3fmX3G0f2ZK78P9QC8eeBZtBEShhwoAK5S2dppXoqHaPU7+5L1uSNdTVra
jQ0qNMgqM4UAYkyOsE7dwhejZ0nAUBWshhGU+WkLZ1Yk1DqC8UvQ6UAOqW0FDaiV
B0O516CAvl+XufVpsYFS5Vhd0qW/E8TO0+lSJnXT0npFaZuH996zDUuSKJAxpW5P
aC7xqPwWkWJSrSsDfDatPkz8HGu0EDIH3ehfbKsCeiMxTOvVe9NJhXT98v949B4l
A3xr+Gka9zC+669dJpGJX1vBIQR5yp8Il3ZdJRSDGmx8OiodaR8JE3SuWuxO9vnR
9cGNo6PZNJdIuhE/0BY/4ZGpzgYnTnX5mgownPJ0HRumnP/+W+Kx+9KhaMmL6uT0
ewO66+HSfO8bMRJb/iRK1uKFW9zwj9GhK1BNo+atjHLaGvJQnStUl1kXKd9UMm/j
TDhesRjmmKdPGdlbrkjebCBJCQEfJ1O77xu3gpTj0NnNGcpNiFXpazUoUHS4KFw0
xgLmlDzGizk2b63GbpSmRSe3h+AA08jHTw0oCuX4k9yIjlQJCseoRrQcAdGtt+4M
jxPtoWWVxvSCYmCGQco2+suB6MYY5Q4BAWlS6OQ5AjW2oCC0xe5Pi8xbNlYX/w1U
RxRMKi5nIY3jcS1e02blVL8ULUWGlBHeF6yqyMioL1dwVerO0SzTUaUykfAKvtmH
fINSJYD0OOVmUfPCPYW6y3GkwKvwGdOymWbc7+AAA5IGF6QxUHjcc/w2Bb1Gbcul
L5qBQp/ONUMG6j2XlmAKAyyqqzHD2Ev4wjIWDwHSumWz4zwzcHxL1g1yFDOv09kS
E419dNdgOVM5/aJFR0ljtbUyKJO18kVL8GW3H8uJoHfHzW/c0pfUR9vRQqFhDR4+
wKQadtrDivnLsRtiNWzPwTCwwXI6zoTNfXnTR01hlY2gowp56yODyWIsm4mTDfGM
1WijDhSvHMRuBOgK5QFkfAzVdvvDrUMdd2MH//HEmPRZqOwnX8wfSBXP7w7F8EV4
FTFdAuXb9ITRB2adiXn0q/+oFfwMyaAfIeghjqe6LYYVlKtSzlU/WTSGx0TsASXo
ii6+FS+OnTNdr1faBOm5kbZDHHI2DBX8EylRlnNZoD5TE+8GNKmitTygu8GhZJJB
QB05D1sdjIkSjkIYb/tw7XeB/QwNNelW9youieTO2UPrtET22LrkSEpaF/r3mlE6
VejHTuE25MWm2bxBKzZ+dnoH7wu6nDpd2P086wWPn45YEo86ac2gaCNRg9dcErMm
7I6PxlLg6qyUh//I7c8QMjgFV1VSAG2xnAspNMQHQtLWxkBgHk6w818kx9yF2FNO
E7iEVpUH4oib+DfzX3rS0xGWaja9eAm61LkRo16L8PZasFBYMQsdVS7ulXvKnsq2
Z6+yZuHf6NgFXHOKk8u2uBMvVfRmEM3C3Nclmk+OS1tCEjsuc1ceh+k9FXhyH+x5
OXAdSZ4wYpnUq9SlFBAzhx6StRl4hdyk/ae/ICuCmMqgZlZ+qv9pK4e5AKtA1GvH
jLJcP8YczYuR3mT9X71XKuu2woQOhFir7tGA55nCqt+/0HRYLRyBWPXh59CLhJ32
d5qUkPzaYi0xefkCsjmAYUcRf5nlqmQ2zOuUWe8HhMqrdfy9hht6L0ru08bnrUrz
G8+GHdZESgivydSmkL1UnYyl7qyJL4ymYalMmsuk7c1UT9Pnqxmgevor/aMdNfX0
NN3wig8yTwqB0I8jN2orvp3ESnCriE6jmmANyKL4/dt7ATw3oZZ7FB4tJWEEAYmw
2JKSicV1miNXxkYuQsF/1YYJXHSvJeguhaSCPzzAw2wzSa5NKfS2rtbhbwmErRlr
3uz/LLtZR7ywjy3AZFQh4uQLTxZrrfUKKbOU6OVL964FfEUg/OpxWAXIFZIpMohc
vUAHF1KOFbXZSyqtKFD3RuZ6oA5QJ8wrsQJMrkSoR8B0XmCmx0bYCJGfz/iqYPcY
ag6kiPVgfqVtEnsEer8U/i4tWVqu1ViDLXT+JBKGN6HMTn3IAu+VnHlQN9wveyQ3
AUG9wxjwaxp/ZfhXqmLj/VHhzeR3yiYY85moKqcnikd1pH7PhuWZRBBP73NVsUCN
tByguix2CtYD5vmjzg459fGSa9AS/aaheLXO/NZsp9+wnZP2EUMhfB+qP20RmWHC
bGap5gvDFPnWnF2JQyTk2rkAu/3WcJLveVeop3FQP5dduiX6MlVzOkWI1ifMlJBg
3PNzknD9eCEaybFBTN07wMJkHkg0wLQ2VhSDtMBI6IpRfMHQIaIFjeqYuJ0bHo+s
FWlNreOuhVz0py6x8D4LRfAlPsPvILjyGkpAeOwnA3FrymiRPxvpe/eOzvePoVXx
fxtaQkUj1vx+vaWETjKKNXfCCVc5mAt4d38ZnlH4YQWY4ynsX6ryAJSAiWXzfy2k
nXbBkah1APE7R9mx3i+DLyHDNQ+0jhPvsO2Zq77V6AVhD1BXhKcDKci0R+INDxzP
cIvhcFRoW4mUdvlv4WaAfVxO8D1BExdMSZxgAeNdYGNbyy9ZR0MsYCMmkJJqPPZS
DKPouKk8X4KuXpYSOvkMa7lIQm/eAbi2eHwPnyT1JcP04m0kl+f7v/6TMRjgGA+z
RxWgkzw4NeQBhZGLipfHbsgKAvupTVw+MXNo1oqghBqarebDo5dsDQI8Jo5IK2o1
NgqExFesgV6rClhj5g0QovTYDBYmAeJuqII4xt+wuDP0EOFm2taGnGs+lLvnQ0+R
9VYk83e6k7tFWh6DF8ICFWckmSPG6TrcKPtLkIAWAWWaGnSDHkoEylE4aNsZH0X/
It/5o7QaozM+/eD51Oe7Ogd/s1R0n2S2kri6+2jzUoaHyh5hVDUyVFq1wxzRbZx7
V9fBWIScfvORmeM+O7sUihfcZrnXwQSW8U+/zstoaal9/P0524m7/1zr1uqc6uaL
vlkBEnU5qvMeBQcna/iz8WtBAl1D4cOw4LAXbRqhysSjkKf/4iWQtb5k4jWYubPw
U3gdGg9JzUXGtiU162wA6mw71cQzBLOCdcezal/12QXeVMDYkUoXzfJr1spuKVXU
3ST1v37ilorleLxDzR3zLnmblTNBWl1M50uL8ZZLi5T7p5DyoYvItAjfb37p85Fk
0ZobODyNmDZMVtFarkBLyQIyS4H8/iARGg5ICDuXfR8BPk5ugLo2Dv+Phowe4Wgr
Mn9NrtO9SpX/rXznD/fXv42AkhAwLmlbYDaDnHVi8FAiCJzkVoxSH2NqXyLHOCL2
j/rrK3p9Ljnz00S0gw93HyeaGpVGpZlGvT2gqpEV3X8oBO1KBSuuns7K9Dij28IG
DAT0CzScCH1WhoDADEVBZ02C/QH692QuYRZWPZx1zOb5grXtInqIQep4nF4cQapW
5sgZ8l2/weMzlOM3/drUYZ4hdf8x86R3aXiMYSuk32i8tf09zXI7GT1lMjcvxt3I
Lk8/6MF5allcPpzdO7uDItrvtk786BwJDIUratOW2fM+RicqvuefCqwphVFU1kib
h1Z8N/ivMDdrtvC3oAQ9xA5eW+wxo3NuPqFmnJOFWbto4HoH5EkSvSaJgfburU/j
rmwegQoluZuDyUPqfq4kW+A8crRxAg5JMYA/31hNQH5a1gEBu+4X/VmNhaoDB3ZD
skpTOUMzILCRM39v/OuTo6KoP/xeFgvX7G23hraqLc48EgmTlGOGEi79IVDwFaZ1
o/OjstalK1oXGSnr0sxwzbJpltjwe7bMVsQeBvAVx4AFm0hD65vE8OAr0uyOUgk3
t4KoeFdfu1EeD1WzXmuKk1mjvOc2dc7WRf4paNiabtBwhkfnTMvZ9Fv714OVpGlN
TXbL1RvXdjDxO93v2EKIIHrAM2Ieo47xTP+2BUmXR5DNIBqPdqkmczf2DyCLURO1
hnc42AE98dCCt9MZ6UJqyZWhNAgo+WaTDRWvPXVrsvj3eiEt/t2j6o/yVXodDz2p
br0rZ/t0tn9kY9jIS55RVYkhwDmZsLjfR0Px2wA9sKnsy/yHQX7bzaPsBR4ClCWU
iu2ekl8OmUuDHO0ddgZrOSm5JEauxW//bGlssZQHJrAPeB+/Z112YMT58KzG5YSl
EIg+W0A24I/76XQJrc4ni3F2YaLzC2ihyqt6J5KyhKtqZJpNRh45mMo27AWBRyTe
DVzP2/RzIf+3c79HgaFT1UBhVdpsu5TheB7xEZJuN+SY7sF1RlUhVKU/nCmQgp/h
XXMyzXtOiA8K2rkF8GWikGRs1phtj9oL62cPKLGR+yE546mqW4WZeTzkOnmN2Wg4
eBfTk7I+wjUNmcHX25XZwSeOu0Kbbn7+uAillL2+98asBzhupOWCdbDjYmh+yHAb
b/D9LhGusZQw7YurlV72w2pvQdZ6C1fgxmy2nxjVOd+GFeQZlgMwDygwmTnVjTfR
ETZn3zYByWrkxA3n+I5MTzONQ9k1Aow6+bnyjaqj9GlQnugXXbnwoLAYlOexIbzC
spmCqQDRLtvYuRLh8PkRXBCrQDYki6KOcNCLLjcnP2LSU7yWivl1sse9MSLOJ0Es
gAx/tg4N0q0FlLlV1qXPX3tSm2LlWmYSiY7s19su0I0HkyV+TBXV1ul2d3v03QYy
Zn9FNpYv5p0F1OwDh+5R6UFIzIq3N3I59tjx5h21REGckIy9zAORsLdtC6tCAfV1
I9JZ6O6gOroJe3jgXcl4m+3+aVpG2wQt2CfE+y3KcPzlr1pVr20hVppiTjcaWPhf
y5H+/dW8jrCj+G2SsiEv//n5hPjnN5oLhHR3L4M+ncuyN8V5Q1k0ZKyPYT88fnyF
rOVaxNzxd4vgt7Vh3+AuoguOCiyJpOTXTkISmZ/2gLHfY3RHwcxn14wi3IsrR0nR
X4XrKjKkfc1Ai6XHrc2ei3X4qMWjvnR/8qkEYa3yEVLgvn9vY0edJPkHkh/BPuf8
JqffhuzDdGDdgR3s8O2GLwtx8ark1QO8VvrZQsVvqjIUFOkv9EmvpoYe+lRchGuk
86sLS+s1D1JarnJ+IiOsX81CxIrHN4KI+VIJ+Zf2VywvFuNS+yO6TH8ZDQs4cd0P
S5Iuo78XSw3K8T59VOe6qylPN4vvcNPtvQtyWCSspJWlcwa/DkvMVejF+i25yGD3
rpg61skF2sqbCTiGnHr1kly57rJRDxt96rKYSgzx1e2BMd95g7s0Ii3AM2EVyVUB
oXzCBGP7vLly4oNyFjYGoL113bqREHkT/qume7DRViOLwJqSIsRtV+p7FCKeYYMj
jPMNIoOoRYIHwecJ/hVKs2vOWhAqYoJVbuPmH3TQtUBDj87C5rJSyftC3xRXQzm2
9R2TC70RJ1KXSuWbRu/ZlbLYRwXJh+aQrRMqkG5bE7kkIJPzzZ0cv7YyBoF8FxOv
PtpVmgYL/UhAmcblK90R552lHqDOX6kaw34SixY3meNH581QIVLiuBfAEMUbYXxr
vl2HvE8IFXQzCH29VOsSeAs2/3+7TpAIF/EAwV3JY0fPckNh+7oaB8nwWCp4IcXO
Ax5r49BkM0UzHRTFVu/q5V0Xc2dlxhKLBlez+NSAHfC/0Ycvdt87R/iNvA/3Vu7Y
R/Xs9RT1xzUhHvVWK2AimLBTcZWMmLhqlggKL0x8IKzuy3OSeg2b5wWh0kw19CkP
jymFcZvzDrvP2a8TjcTk1r3K13enUynslPlVkDjS0Q7cH51RQWYqPeqBtCOAMR4K
18/6pvQHMea1iecCDXPcxlpMYj/vsXHNA+8vvJNt79IRU75dRjau9TPDHCyBt1GH
4axfaN8InpxnhP75zPGJeLmlmV8Z2C3OUxQoQW/adpPREfpjrVOyakX51oQ1C0ge
n4Ihc1Aw6WDcvg5i0+nBRC7Ged0Q6oT/kRUdzjKaLSDmSnhI7cQVz0PZcYKj9lX3
8znusNWpM6eidPb5NfPvrrppHwOc0thNgdOOnw6wxFmDi9OK66V+Bl45VDgItyhG
ZArrfqATWPCPTpUK4ZsEDmP6nOF15rzeRe9/qpZpBjZvByGtzePXxy5IJYOjb4ON
EX5qa0s8dNTfR3WGRmdrlKPB7izVRaiy9XnyT3AirjiMCHq5pMhaUbhh8QOPh0rc
fcWjy+Cc8YyRjxWrT/EF5QNTU/rLNI+ymlzxXInk+yPq6qTj2ZIXk7FeVfJC1PY9
Kss81yyaamIkAxVQwrsql+xcesVfdX2RYlYkwBKiMG2Y/kS4h7jNc/aIX3Tk2jSH
PQpqBfFSmznkLkCgpHKoSf1YPtoQNDokWKaxhcAYN7HlkZU0RJJZ3+QYFsOUe5xX
r8HNQLNNqH0LIpJbV3VELj/gn5Wx8sDLImpxmiYn+EEC2e5Tyf6h8hkq+WfxV2st
H0j0flzKCXomxBejWX8iIZiUpnbhWBUivzh1Nks3S3rZMbFqA4+GgKPAIMarwetk
j77UiqUmcFzIcD3oR8dNOwLekrqxkpFJzH6jM631/5Q+aY2c59U9W4XaNZWIsJvA
LrM4nPupyiG+bjncxWsmMSphjU+0rEgH8U0y+Fj+qn/xlYowzkEvwstCK1yqPAPj
RAijQ78iD009r2zYqdF8SU2I+A1izgn515U1mm4yCKSWFkv+bmDMep152RpfHMO5
EDyfihh/TMzxZ7p1ePjm7ndZMmMsvYh/CcQSOZ4u/eBc3GBv7K3zBRuP1oS10VeY
h2V9dTFnJhiSLbDexnECiYzWmkAo6hctcc6uv2lVvvrvij2HIkf4wi2dZ9wWvD2Z
2OmhvcgoHw6hFAulv33A0alg6Sja2+yFwx4XzsJx7C7COcYkAX1uAe1m1V4YgF5D
/6uSo7Th99w53GFTKCQutahcoYQqKw8IZWy7QVceE3/66zhBYk+wvCLh9NxJ7zOr
nGCeABaGupJVrWvFNkTCNf12GWI7pkhgzJSr24C9Kba8DgRN+hUR/sEHt0W8Nx7/
/RILDHMVKi0CcaGCT//YIisbpMhfb95YjHDRQi0eJQnuTt20gojjlz2kr4M2XwsH
yNzSd/2VJbnO4tYnBbbG+TPxHS1JI+Wm39gOj5FTkZEOqAULAZVZJ1KYl/lLSGEw
y/tkjXjax6/mNzphNHCsbSyFMYYuLveCzOP1udXkBYczIKyFPGwy9Ikt0XlXQWHf
e8IlL8mksLvRstS0Y84T53EtouL82oBQ4GNBts6PccEOcFk10uE89rXDlvStI4X/
8bsi3VKUsK8hML6RZivhdYmmevQ3Cz7+dcgwLdxbQkFDimO0X9xE3vuDWLcdPDgF
K/VcRErDD6LwPaE1X6I/8iRb5SgoQ1pIrH2VdGjwuNfzjrgZufXsv9BpxUIPZDB3
Khpw5sNzBgV25OAyC8dhrGf86x3dU54N9J0CVH2lrwlVnxim/vCa+ZAxQ4UhbF0u
P8fbpBY/0oAavcDXSKskF6C6HmMUovuksQZola1BKKRrMBROqztrr8AtCmGB0OsL
fwy2mjhpHHtAQbSD88OFSgKcswGKGVJllXgQeQ3/Nq53gYGKJ+e9xRMNnOMiiXtX
rDorqtd3JBU4ID9c8NsTE3h9cHZZ3hEPFo7QXQk5JqEalM2z41m0DRTf3si06bd0
/Saimqd/QUx8GKQS3LjjEZRHSKSx3IFu9RVkfsiflhxLwic/KsfYmus0XbcdlMcS
kpzWhnQbJfcnpDmKdJiwvw40Wqa0178W6wtUF9abgB9q3p50toKIc0BqyFjhCqFn
bcvqCcrIPRRIeAGTUqiut2fHgZQ5zTishQlkTJ8SBAgYLs1Br224dosr4CR83a9a
CADtAmwAPy4t2JTwy0HcOS0+v8DoSAT4Q1vf4Tl46/tU0Dc8F1w5SqA6vs8+q9T+
RGYQxOrqFkkI9Rs9cauFvZBXe0wFj6V9qRyIICE1jYGSPXyIkm8iDFbbTEDfyKZ0
ZrG/FT1hqrn7Mb6DUvrmoJl2PLE1WagVbBudE/6dXDD76w/amf3/6IHdD6PK8mAJ
PrKKeGeZHNEzpotvnvuSBdl2O+j4OWZeFQbcRdDV/MYbSVKv0VkIqVz2OWqAKV+y
5tZxpthG+b7QvbbT3TYhU7YtjBEcr8iqsjz6eMMeJpN6helxeobh+xDrEWU2bLO1
vI0GpeIkEnO4mvrM0ZYSQPuOZEdESINNpKSbVAtrAzj6vs9CYDQMvSRnhkyNBtaM
eVhLd4QaKDrrhvof5ojhHNRKJSnnZL+LQW/HzKdEjd1SNnafk/pEBEGsKj9vKqa7
qNgsYuiWPII3w58014wkr8q4IIcKVejztDQsazeAXaA+88g1I1ruWVYjTM1hxhCh
hDOPOqn4jI9hMJ/eYHnEP5gUXphAChd13f6WMISYbs/xhETbKSviwFgJjj2boLsW
KJS8q4XwbpDBm8SFMXUP26qPKlrk+7N2+e4PacFdqICWOoyOt9DzcCqQT6lnlPVZ
qcBdYKB8fXsoDvn01u0W0w4XZPCEXFKsbCutry+C1pkDoOZjCXeBWyTCmft9Uksa
5XlWimZATfpblJ8+iR0CIQ0aZa6etYNwmGaT1PFn0a1p0twsd5WXyLGJYme6f6Jt
rM2TgR6bFLDrTwF6Sxfb8OPF+dwLt3zZlyfi3P1FR5KjnLpoHtfECU3Cd4jPLtk5
7AbQqdlo1B/oy1sKYwrUIlUsWnSdKh7qSzk9CvRCklIa6cOpgY0sqjKfdBp4V2R8
naTyO0IMcNN8s1Bhd6MbHc9dKSUVOv3cGXCMDbhAv488Jh0E0iyrXaO1x1H+42q5
luP7BtRc1mD4xfHwci7zsh3I/onhUp2ejJ+/QdCcxgzqshtQwbjKL1ZkGmjsvvzX
hjWgGSBtRsufAGJzOypubcAw2n8I4arRSSVVI0oXTKTjxuV9CNoshEwuFtw93PUa
RU8esEkazxapJHSeDfRqiEsjJicOJi4iiHYqu2XhnL/kVIo9/OrHhDdN5SU0fUBL
ae9P3sdwSOBuElGP37Iz/sgySc55Hfx86hXtVd7ZSidSObkN2d/ifzGjtdwNeSyj
RiucWNknOqKGQCc03rQaqdTNZaWTIBy3GQvPpdABPUWQSzCWqbUWRYE2nn4g78Hm
YwAQjdDpRNe5hZO2/NKh55qqxKidnT2rFpSXpEgMJC33Blno0aD296IOMcsD+Xkl
adI/VtmYE47S7TygpR7BtraCVc+9E/pgbera2r8VCEBRqF4gNB46qfpuPfBQyEEJ
+/riZe2JFN8YbwsJQ8l4PkF+JBQsNCq1AEZB8deqxHbVIRg3EhzfevNlFXvz/c1N
DeUvJdNoxHfTIrHaZ6TMVhgghP3cQ3KrgS+MJkSOPLLtS/KgRkxmijBP3Nv3Ev4V
m7yTqzL3J0Fph+fI4J0pgwPIjRrtaIQkFo/o2iTV5vW67voY+OUcU2jK/z+a8Ck+
Yja+/OxRKMgQdJYnAlybf0cSHB94aSlwCY0fwhxLjBKCz6k3Aj+GMDJ7JPi1bvCy
SDVR8EYYU8omc/cjrD3Z0dVbMXmE/Vvg4xNljl9sts9GegwAgH+SoEWJgvcV+I+x
heB9scTXeNP/1IwiKBAgH8bcSX+kPBjDItQ9sLLeb0f3FF/yw0ylp3L8NxB2kWWG
zsuMTD8dz1hhzj/dNiMyjM4QX36qNfK7clhiDdttN7BlkKjdDYplbEaIfQ8cr1Wt
IdWHKgqwP1FfK2E09ipBSCrt3+xKBfifEf1vq37t6tasJIUW0+h5PhA/jH0QSXlk
FIvVJs6Mtqgj9TOYT+7XFBwBwsRZQyTIG9Y9ItjRGbAGlHhkFdErhKUuG0g65xvR
UAbuhhEg5YMFU0oDdkSoiZyD22vNlqSDt5cDsoaxLv1AlqDMPkdS1B1699XHE3Cy
xNQ8mdgvqS+mGMY05TfXPzJ+fiCr70281dDsPtPlcf3YJsVMzMQ4xSWF0OUkHM0+
A3/gLPz/DsQNdwM5HXTkRkc4cBBlzZ0RII2+4wTPBbtdVsCa37M/UvuPJiq+V0+g
6O/Jha7H9+dk2odhXFUzL9P3Y/2qfkqmVNzptfYNKtbQ5G3G/nRfSX5Vr7TpZe5Y
ykoAGlMgVDfjj25cSnm3bRtvQUtNyQGYLXwpB9SdYspUv2weErIsAysB/Dm4hvE0
Ncb6hYfNpL1RbtPvVgQ2gcE4yfwzQ9hdwXfHHbvxLXET2kIIGWHXVUNmKqXNNq7y
Kfj6oSF/tJHq4YdsRpbmqKKZPKT/lRwiHsF3Hf711l4LK9/zTqWmED0Ty4WyPmuF
F65Oeu3Fi1VjX9xwo8pWkTIbOlYEATSB6SWGe4wnbi2zbll6Kip6YNeCIwP7bAPr
W+9Xg1N3Fi+cS2TEjkeEFnLX+Rxehnd12scXGFsnSbEiVMjk0fQmITjwSi1BIUY6
lFfP19/rO7pNp220GkPU4KOs5I2tlSOBWEkDKrfdxkGyRPaPUWaCDBF+680Y/sdp
TSsxSBeu0Bzv312foyxzERrjGOpOg0Jsqs0WiE/FmbfFV6pLydqIXovQPYfAGE27
HHgDh66f/rlWY4q7EsFnyYUKm1Ta4VmLI/o4iCFvu4SxGGTn233SvvWMEAE28UD2
ggnOL47OefE8BfymmLUBjYgDR+tU/gJKx95oaCoLh8Gm3ePPBsUMU+tdshsEEjoI
o6J3qs3VHyAifLAlbp+OzBduOKZkPfGb94WOSRH9Y0ziVOQM/2pbhQLGhpK8QL+y
oErBC0YZGjh+bo1NznYtbw+2lJ+NNBxuvrDEqXwcZNc4d6AFW7wTMJPtCAVK0mXx
qbhHCBNkMTH1qeUsGG5coZxfQ6mstA/IesOxHwaAFnQE/NliAY7LzSH0rJq0fSh/
7oJhq5O+Yisq5zvW87yYv1c4bd/UT9XDCXnUF1X2n6HK5FSLkT5Kwd5FVw/N7fus
I8oi9rpSlua3e4eoGY8WQOqMA2alnfbmUcd4BWOyFlbMEi2BMS/O0ohIrk+ZATg3
M3PVXeZ5C/wrjk8+TIScqi3FnR/+ookolS7HJcsrFB1z6VYgL+f4ZfvBWBikCeFq
QAXqVJSTguGh66XUuty0nP/tuDy+dfcgdbeJa1bNv3WWp31fcZkiMBmZ0AsHGUdq
b3bnc9i3jPA2qJRIbtc/sFTRdAj34L1kSnpOG7RqMLMITscndr7V31QhsrhqLj++
qOY8v/PfkjqbFCnnMVSHUhQji4doTg54kgGASeDiNazS6jCoTlcEo/Mc7sY/5D0e
SJw759xP5qhI7A+LTFJScGZBfrSvW8qoqSmDN6WJhtOPZDVVGT8rfEiRc37CEYkT
L35gSC7j/SOzJCceZ2+MwljSYb/pR7h5eWJTR/jEOHcT54O0JDsaLIWaA3phsdr6
sO1FzaXolj18RNpOuX6b3OeRdoL0evartxUC1mFfkp6vKvpRQCq4KPPJOAeB1fFw
PgadmRRh4lKiP6kFG9EKqZ+4bS6N3HNHsVSkH23GHas9IIRqiiQnopbqxh1n8pnC
GhTfMu/aYrEww5E2jnKXSgZBc9itCK6AterAMRNkJYgl/AiRK82we8zPtif+Jqny
kjASGLgiZA/W96+d+sk/1biOMNlxDw2/gGuvLLMwyAIOxfWXrCbL/6UXnSC3g/rI
VfKFWfVU3Tk/4l20EdI7ZVnTDA+1dW37SmclNQrFffaVXJX1c6t6iNFnlruDKwKF
MHmRC/ArnafaQsNYPoriA4rpO+DcxEjuI950A4tmOzs2r+/UsAlX4lrNAXYaJDcN
646NQNHNqC0s04kB7gRa/ARY8pRH+CpR8KydiCMEsCtc2gFiwV2KBPyABXLTHGcz
yPMUjUFrgivMl0y5r8fHkwAahc3yNvKTBXwf7eexPyz3H+p+sSVhrhHAp9g8liVQ
5j7qw94C1p0U3p3Fkg37ioTOVKM0rQ8mUSaYeS+NYNXr50/4ejHbZp65z0dDuIiY
zw4gOX26q6QZzay5EQXz74QkmTU6gFt6JgeFZycRDT/QOJnSUBgRBHWa8848aLex
yNzFJxa1Rb2H3UHhOO/gFPc530FEzE4E1lA3J+GcFr+2/fCt5AuUaZSuweN3XqrI
jsmkypthn8i/8CT6xLSLzb2mRgtKycHPK3HSFTL/aBEl+6gkIsaroj9FPvE/kdK9
IRz9NExQnomOunZlJaGi/O13XTtGAJQ3ymLqk+MUgXkgF4HEm+joGn1onGWOGL44
jEeZ9dvNWMw+ZY3Ed2vv3lLUWgK7/10b7SRACE28mFyZh//CQJ1SJePpVXcHXQjp
gYS2vee7YA4ubCmYAetKRdVXazUqCp8t86NlqL+l4P92K28gBZUBzqwRmfTvA9tA
+1xGDSp/iQ5U6bU5tSXMl0cCrPBIbZ3fwAOD0PDmKWnlzjLStwo1GcabIeUsbSEc
KkQzNzpyZyvvXsjjeX8LkAUIy9+SFQwdsiN92vivqT/jDJFKmLK6+wZPgHKNBsq4
HWsjGHoq3voudkK3NA6kd2wsvqfWB0IUCxMLoLlJcsRKLhUczuModV+cpFQeoqPS
OhLuANkQk5rCcPPPaPkYISWIqFvrd6GQX+/TMvcdseyEHBDVsyCB9X/Zls2I6vRI
vzh/I1bKe5x2f1yjR2eYZ+Hv4cjpbqPNNWtI6AF9PHoG/L9T46j61RO2wBMkYW08
4DS/VyrDKsW9haoi32cB4IiunFj+hD0/E3ro6dRoCpP2fIIoHnQyzdID8QWorQhK
OaxljQNRehIt1d4zD9iGIGksOKxbfSGenoGFNhVGxD6gGK6nrVzrZFQ+Z4gKk67P
EsbatdCuXKCam9ruDotTeTK1YW/0P9sHqjqDucLrDf4s0SmxVBcz+1aIME4kjjlf
7irQHcrjiiqHVPlcmacztW3h+BThyXbtlWcMHrjJqyr+bpttCNIMtY63vktStg34
lqwNdhp6ztA8Ic4v8cwKwYaXUiHee/QvSx3IO1AwHDMgJEkXD9cjkH1iKJFoBcrl
zMJVtMZluaz1Qq0+RkeHErPwZgUfJ+LPoxn4kD27MM4K2jWdHcUwxC1PnXglcezy
h7Wjtb0J0GWaYyRet3H/uEEZsUxVyV0u1oZgVDNA/rq+GLSTg/K0sMgVey4RWs3x
xcwKz6X4xhpNHT890jMw11L2RH+vTp0lvghQ/r1tdbgiVmcyJE1tpc/Owv9r2kYj
aUOD5bKOj6YdhFnTvCozjtZoP7M0EN7zbKfjRerdIMqyzCiyvNW5sMHo88CKb/+D
QDY855sESKSxw5E29RjXRMXpMi8UQMSyy2t5PqztBUFwFbrZKiXjoNx6YcYerP41
IbGYIVAJA/a7M9sutrmvmtJFANjjn0Z1NNLtqLrwQGMHdCrl+qTsKgrCuZ1WnrK3
IfQBjOvXpAwE81+t5irajboChPgP/d7m8Z3ymZAYkpeBG/2uxmE5k+U6yU4j6kZz
oj1Jo8xE7LFuBq9TGvDs7qTELtNPpjZU1al2+QHcMuaWIzMmdC7v7w55/tT8/G4/
0IMyJPd/Jfq4th8wZq0TjEh1haq0axSDJK2Y+q5PMFdDNPPEec37wD6mPaOkceKk
cgnCnXnKhqDB01t2XQN0I1HAytc/2x+wVdhhTv+ZJ7U4HYtOIiJ41fGBZJyw8RjS
ss+3hhHk6sD8/9dMAENbnSkckKc5l/xlRJS/lWOQlEz36cC6kJmo6WV3FPHCYqwy
cYfNl/ApaVUAyCvPVtAaC+TJgdL+sP7PAsVjWr8wD2qCBjOIhBbpRsKNdQSY3tjT
BB5+8ZhZ8hqDkfciO+S09xs2BlTqpAWdDoRIkbF26HRA9vKhw4RQNEeBrkjog66A
GK63VC5tjw8XOjdr+A0meOatfaZkeqcMwqSmM8oEQDDe5fuqKZmKc7wVnF39mtnk
WcIwLlxr6pI4PoksK49ADvw/7T4dosZfwmV9fDIluUvYrmSuQmTPJeXLtHTgfj2g
SVXg1vq29TBpQAnig7s5uWTpKy8RDeZd5C0bBGVSp1lh/hd6/kbiCIv126na7mIF
Q/+ewvJ8iJdSNXtlUclht52RGFQvgxgdWhXjZL9bghmZarncWxwtewZ2rRfL5EI4
OGfM7+PgCJMNXj1dWhs3J7ePwdVjzHgIkqQI2CpV9NvmdN0siIhviI4eD6DIQhEk
U/uPscK5CSdkah8Xg9fDU2de1SlAexb4uUPlHgP+e4Gz6jbjKWeXYzB+5wGvL8XD
HKvu5rmNma+sa2w5jsmwhKDdXc+qyCNnOJ/LEEYXDbRcuXHz6eZNFKk6onsPNQN5
TanX3ujdVjyAHXfaxAcYge2bi9RiaIlx5wjsptcZeQlh58eXHFCvh6vuUwIrp4Ak
gcdMWLp88RRvCElFFUT8Iq5Xub1k1YwByUJhU9s6+RhOceFKQQqkA6WWmkV7r8zy
kMxSd3gkHnmgE3tILCS8Q6f+3+XXVhYDO3WfXLhtKcKUu43qqtrcng1tN8b2PHYi
eBLxg+ErCa6PrRzcE+YAChu/SsXkARZvGoe8ObP7cDzJ0/4ips/NPRvNqJspvoX5
DqlBSVCUdMTbRh3A2ytcdEpWNr+eAPipSpyvs76h1dpbyjZadiXxj8SPr/6BGc/t
oZXI5ILfgG4q25wDZdO4Q6+3YpVtcRw2gI2cao9/d95sZ4FDNq2gs2AK4WfDxi0/
t5Ye9BpmEh0WYo/5h6GC1S3Xjy55sguf/I5QYN+3nvzWioWu5SaYMQGR73IZjCeK
3P+2l3Hjn2oAPStjVRPcHZjjwkUJ/4bDxtY646fsO0PpUYMr8lhsRg/NPQPDuLro
os+NXd/crGZaN8s4E/HP9KOV6gE1SFLcG2P8Nv+mI7mFQcpxz9iX4qfKg4y+0ffB
dLib3O5m17A8ind+mw6KUzFlTQrcm5phQL4nSxnJ9jmHDCGsQchQUW9xk5cCaCjh
Za8fBa1y7Z5STwU47LZFLs5B0X5XVcH1gXeZurrXSrAb32ACcugdQfh6oGwQ7GtV
UIBkgamA8OjlL693zIAxqmuH4JvG4mRA1Ol/82PXb3FhgddYebgGREwF7NHRjOwA
0xyoi6PFauqjGgnSp22u0+6AOusLRxfFKl//hS4hTlqj/MrkH/62Vjld9fCzKv23
7i2tsm/LHUT5bBv9X5Y7VUlxKHSggLNSxSGOdSJWsDCGNwF7nqgmoyPcw3K/z2CF
4beYzyCaHFuxoa6q4WBRc+kH8P45X4cJdLD/mC1Vp1WubJbYknSPWOhDhPDFGFFx
MyVMMTLLl4DnoSTL7f07I7+VhWv2UxOinoL/LAq8/BgHnfikcUXkQAD4ubUl7W7m
Lx40NDigQGY0oAbB/PLHiLmuw8HYdzkMmDz0Z9XyCam4dmfbRZjXcj3k26SexXvR
RCSeNAYBB8TmGH+oZoRVAgyfirIXDFkm/5wqZFUcsQvzvcQ62NlqGhRGCSPg3VAf
AIzK816Zfa9cjHIGvTdYWCtpm3prKgTX1Fq6DA0CeA7jucm0VN+Y9YVqEOw/Lmkh
ystzJk6X/PlxKk23cYVjVKPTpPudi60WRQoceYLVtKQJD7LLU1BBOL4LatSz6oJc
bg/MPZxWQlQ31j6udaKCHddBtrJJMN156efIofpf+XSk8JwVr6AgpvsoJZPtW9ot
1UJDwHakqH90yiq+UYh8o8XDQ65J9rMvKNhV84pJmpRJtRGl37KdvUnAaoRkM9Fl
v8tsI34A1wE2Xl7OKuIP8Xfxs1/EmdWNs5Fdx+5schm0k3xkfc5hDjkFskjXSRcE
Gqq7JmIalhbHcLPVJRgmC9yaN99C/v+xhkqx8GclIoCSXPm5KIUNMTfaREP8U5SD
lhK+SYJ9GSDINNutw1BDevMfeCjNulcE6JKm03JA6xQTWr/tu0MR3fZf/botUzc+
MPJ0jTqYXy9HmmsCgJoVT0D2wLlk9IsIxEXKL90a9y0Ze+IRU+1WMQkM3MajzFJ9
dtO66jqAGBH5C+nk8CFeq+mJF8PCw498qRdpk5yrqgdqA9qbco9gtq0uOwSCvTLc
dvGSj2tFU4Aa7VpfkxaJ7wiSqgDgIXxLqp/85L3jLUh0szC5qmn6SNxJu7O5IHeV
0jSvZhjr/op+iFrXYwFvcPedbWuycSF/L0JArOJddcYKIaJaECsCP1tKCuljE9v4
3BEyDjwQyBToHL5YUDpfYpYvT7s3yMMs8RtkTECbXWycwOnk6enS1T/jpb91Zv/3
BsupkJo9iARsKiIA3c4p/Eh7rBAqivUJC+XzdpX2XWXX9M1HErQeraVkLqd3PqHv
zCehb0g1tK+cbB1sbzGECChvRcQ7v2lQF+EMHdzWjYUBg1ALSetoqeDcOLrrI4/C
Z+QQNs/EnCdFw7k9OK2q+hRpK3fIO8S+f9ST1WKeys2JanH6Y07e1mv/xfzw7I8l
2duPBcJrcN1PHl77EudNDeKDiyKq8daoowOu9aHPLqzh0V2UNEM5K1NF65rbqHkg
1bYRMqTlGNX5JJHuBIvgO0ek0XuWHUVthi2+uN649ZBEURrNS77tbee0Xj8AC5Tp
Uxwy7R5apgsRQbyl/a85dnKawV/nlW1L93VKaB4jLIorddt6decnqXDxxViZK3TQ
T7ifQfvIN/J8Npqo7K3vMjp4dP9yiXajECmOIJRuqBktzfS/uzy7+q20dtQi1gpl
LfLAFnQzAyNcZaMDgRNhR2aDfiRrttefukHvvf5u42z1UQQ2dr5L/oZsHD/cEGUP
15whdWGVR1wGJVuV6D1H/iII0k0JmivANdQrKOISpSGpa0TKD71t2Z/NkF5jKId9
2+znmLPyBQs1yJINPV/9aC7PK1/SUirBy9TlqWVUxlLgdnjw6UMS+w8hmQyl9mdj
3+sYV7g8DdkKl2+O8HmqS+b/EzDWgTrPCRHj9VSJHU3W1+15QOTp06c2WO2aIYxT
3jpwf26Z1/kHuAjvveZZNk7RpKT2dmHv4dzwOpdVmsunkDVbl/OOSWU1FHCikGOv
wbtOa+hHbicNM0z66qDcpkFwW3YEQDRNlXm23fzanQD3erKLytgYm8sV4cZWIvgU
Cgbs8FxDtDbdaMTX1CxxKGLVOlbQF4uKLzkpcnUaxTzhqagO5RwK6R70sLr98ybL
qTnyFCBIpp46QykArSVX06FjaLK+rd0LUAdpfnfOJscGI6RMy+5r667TP2oPb02x
KN5jIo6cf2BVJmIRovgPobPqe+FrfAJOmWJHuJwnn5VWm8uZAKgBFQqtEk/8FIY9
phhl4di/hlB+3K1cZXy4Apq1unwRECsxauFKffjF7zwly1qA97UOwLN4nTYvvc2q
3cy7ZS+TdIjf0DgnVKAzZECuYjMbomzOfArmjWWFjfvkT1AQr5cnYrfyx1kX6LAr
pGNzu7WnIffWXJQTc2gl6iasCZRZxunytwmp2pSO/7GFPwE3zU18x+5dZyFNQdUK
QldC0AeCmo6G6B7mGqXq8EEbexQsK3gfqz0bEUkcRNRfp46L/mNz90YFXTAJLsDR
e5Mys2jb/GbhVjLtZyI76KlTLL5dM7fTbFzP4InKz1UzJyEx7JIER8uBrILOnNFx
jXTaoZ5ROS4biPQ5IspyUtVuNjU7/GYvBAuiAgY50F9zKdsLDxHB9baedfTdtINm
BMAHovSzhDEzCCHoXWv+YdcVd/SMWnGsJSGAuPnVI5r0opYdj5OaHlMzyEQJk6xL
meShnDS7Ujpqo27lzr0VKqxcLaxSU1aXjN0sjBpm7XtAZ9ZBH4jhHD2RUpadFOir
l9SQ3dKRXPwhd3q5zhAONrZ4vMOQdknLi8Cm+ph0RD/JMm27U3vQiAQSG00guWOJ
yHzWKStmv3OSNNjrFxCULDijb/Afj2OAAV1Ik3p+PpJDT3JgjS2AbHkZNw+S088C
n7jEOKhSZ0eElAhJEMIpLwEOADXw5uTVYKGE+CapowhL3xZASdDHkxJezTU8Kog4
WICSz8yeq0ZTQYQ2fVkZNUZyDd1e06EW7Jo/XZi4m0mXNIqh4uj7BwqT2Q/5usMK
ijCLAssKOjAJRNs5PDkuQz7N65M5oENeiSpHyg+KarnIvPnck6FGAJU1luxMsZYF
JiHdlPlkO6OYvU0tyES35l791IMy1qhWW9cuQ0XeNVrnoiWuaKBTSNiYD9HALv53
M5CfNH+PM3UvBr6PHNeW2OhW2M3UP2KYNm59jjs4OCl2S5hC8Rd/YEt3nZ558gvz
Utk8J0OPWe6GGW6sZ2/bDni26tmyqZjxQpbwV1KTsa86t4LnROas+BTc4OMTkQcf
x8LlO3HDV80a64BWcARqRQ9Yo/6+1XoS3nXSVJwG32xzTyZUv9UmCN7XePLoAuBZ
VJfhFtm8Sv5hd98A3u9iHQtYNOvo6HAJdDTYg3BSV+Bma7XE+s74OX8/MfhkjHou
3Aql4kTsxwZpZaTQY/s1zSKX+KHsKx8jDH8PpoDb/aYMkLE/HkL2iJ0PjO2Mptk4
IU6qF/Fj1ftwdUmpHMUIbOFXCT1d3nCOcEOoosZzGrf1YJ4ATWPVh+4f+oQcEpA5
ep/tNyAyRIruLmv3BRvuQ2DZxTLiJqWPhV0cf0EIQywO+7Cr7spQLdP8lDvHt8jO
ZlkC/ZE39JlWK8JbmBp1YMNcyvYaV4ExcJrRhC7LHTZNc3FqIBuRdQME144P62Dv
fjih+exLB7pGzyQA5QBMwaC6Rv9ZSlR2I96rQD/wqbFHpBzRTvxQ2VYBZ+ZswL21
mle1Y4QOvpSikbRqsl2XFQDj/VlTA+sGpw/ekTupIwmxcrhql//Bo8a0eTxKih96
Jl46jIRjip31NMjWiTDIWQ3F+fExhGiBv/UKLrd3Q2ppsME5aR6Fd8pPLnG4UJod
lPBXOPwvbzNbwmcTkCJyNSAodqXM9lu5u3MCw6YlgDUnMcridJF050hwOvCS2oYH
7UxEvt/xB+5bDzd2+Cg6EFOdaNkdUXLDE1oHV5qkqFjEtORSIvJKg1X491wxGchS
1uFG4nI1JDIgzcq7gjI2qXIFKJ3C1XyAVAcSoMEaShMWk5sw+DeiHFLA3AtS4Z4T
BzyfPXtV7yx4dkxSWmVv2TFZT2eMTA/5xV0p4/vfo8x9QsjBXJFJL9vhu8yL9rt8
ta40RREKdmz9vP5W+dVm9xrzZ73HA2jeHqeX+qb5DARF37m3UQWKDtnNQHxb/Y9o
Mm0imtsvJIRRcPEkJl1XSnuY+Cz/XlI+CRxS74HNEsXtcJp7vpmyGHXWvZ8Q0nXB
iTWLhxFDLaB9zO432PvAJPmgPsr+EHz5qWkDALto7LM66aRb+TrXq6E/PQLzjCH5
Jq2bPBDphud7C2V6jFqxCEhV4d4NZAobj7SuPy74Sn3t9BNhKEcAQSaVywyef79X
TVfipwJyFh6qcW19Mxk5NPyZGNFcuvMT9pKC/SHvgcLeopQ0mZVmuY/vVvuOOiGi
EyipFBv2zDOxn5cN7j7iYNCMR/mdAtXFwATr82WFnBmOHMn+c4gffHzJGPDaytM4
i5jTEuLn55UXy8nZebBy14TstDKr23bCpS7hN87nDD52ID7rVkMKfOvEA1ZoZt/J
nHnUGV46kZhK0C4O5hJXE2cGn3mT/4gx5Ofgw7pSdjMVJCZf6e1wZ1tWxA1cTKdS
O3GH4P0qioD4pzJayhe0YuS6MRnPQ7LgMsHfXuoCOnjLxbMiz5gsHqLvxC+hdGns
z5O9/INqYwyPapLQNnarst8UaKUnz5e08HvTteGSvnQ/SG1rJZloNGjDLLZS9XxR
7p+x6qEiLla00HtJ9JI/USYzVrHPkxcFNUz/+MSP9RHrcF510SmJmHRN6zLZy46g
0opELtq6xCGWN50HAZ5Zf08j2bCpF8naVp1Gg/HPT7h4cJ1b7DUp9HkMHflMneBD
711hZtrf4hO+21+5wKUU06/xh0gtRImo9HPHacPdMoawPdvOfkfqxGY3afogDgIU
uHwMxtmUKZ+OGvsqr0Ml8xZj1JOj1YXTYsixotVeuEFremZsucVNUh4Z56/JzIOF
P9kXwL8Z2ClTzT5Dx2jwqWa0L58RnV6KscV7RTKSiTYeIXJb/fDCYlUvoJzAuo+v
88h+xW+KotAdpltpFppu07MLcynp1wIFPbEQoOZ61A1GidOY6/xXtymRp+uAOJ1i
ttajtHjKhbKd+vDzYZIK/stz+U0No7cJkEPWWvuE9IA5gD1myZx7Ve7G8FzC/cUi
ghzaAcF35WcEZkoYBbCUJlr3j+43fDZ0eDjg+UZQXr3ntuX+T8Y5kA+fD53ulbs5
IiE+6T3czgBoi1iSP0jv6d2HK5cmyFsNsJxBIFFhV848y40YhCzUiaQDPcDFRJ0F
PWqevQR5YDGw2HTlQ5umNQEGhI5lNkbeAPnxBIsVyM7y7YbZX3GeJbbLfdSaSaDM
8od/A6NOcxhepRfCe3syRa6EkvIOAECjEx8RH4EbDb/uFuCjNRXBjfU46iFO6QEJ
KJ5pkBOMR9mqhbaF/r20oACJ7gVr74X1LPP8I/8siU/TxV5qRpM47eLc5B+mbiLR
IWmBRJTvUf9zMHBbac5Ac9loNQY0+WGVEg+AM2ycVTA8pIe19tV4XI6IUO1VhwPF
2vD+uWWVxgPSwNh03X9GCGXGVQeXyIeKGydSbIOzEah6A6MmdACO7l42ZDl2WO6l
a7FsUN02N0gnUxWZJ+X1jecR0iTLmf60U5BsgMXeWDBsn6KHkX40StPTQ4oolFnu
adbjkp7Bew4PKcNtvSw0N6mOPrnY5kxf3TMt1JBFCUGWwkbQKXjmUKT5qGpOVUNp
4IDbeDC0mV6YD3WumrFqqwcYloA7hJkv4gA9EkmD6zK9DbhgM2zvGEbxxusXtt/i
hlaHVYTNmqQgKWw9YJf0smnXWHRmNPL0qGTejrmIr2T5zZdSXqHSiBG8tS24tLrg
uL1MsqzlH7lTuZgbjlce31WDakJocIcTqj0BKhxXxE+KfjpJvRoKS6O1BmQOOns2
4orG29paKCBv06IkoKbYYG7cbzn1/uXszonpd80YDbdiwEi2UwdNV1oCN1qIt7XW
jVWKfvXQvOlhYm50qbKEA7l2vRxR3kFtVKrygptb+fU/TowwjNvghKjfzCOHPjvK
Rw1QKfvq1B8Ipt3DHAitDHYFr+39+JZr/WfgrXROx7du3XuYFVkL+26mWFFox2SX
3vMmspdWmVMI4rRkYynt/cCOGXr/r44eN0Ehe+013cYnMVlMcm2OWVoV8LJheRTx
AAz/yoO+JSta/5d5w3kuEBqHKqYRzGSvarNNV22znlaqOn2eC933u08088Wq7ph+
kZa1BEPKJkH581kTNPxWv4g87y3k/STl5tRZBCF0v2xQy7IKtApD7OoD3nklxtQd
VPzKMQ5LnDgcGI+e6rqoLsZtYyxKoKi6+9iGFG72VFQvfX5Av4YDWIlUmXS0DL9c
rpSJdeZp4u8hkfw7uetFeED9GnA5C5fF7IQ/iGkApnY/gMfVzsQzulguWZx5MCmZ
iOWrmv4UPdMuYkslvZ3nLbZWZh5MSfsZozgxoFEWQaaHObEefgXcvYpLQRKMew7v
4CyRmZcEPORteKY6BzLALwJecN9WJEm+5eBFWkw2OBOsUsIXQTqcSokI66LQniAH
9RYn2V3DWWpwzy4RTaSyv2nV/gM990O5oQdN3WkC8Ml11xB4d088IqRT/CUHbbeC
9Bjxa2ocV0Q7iZGjL65TIIQMw9XiOtGctRyMMYKefTE6qFoxK2y7/MPD0ZJqINEe
Z5yomJDM7MmjdpispSSKNScQFCgEqMDoiT27NcZrc5w+aoqhWG6T9o8q7ilwMOqm
gIlC8hhShrik/0IGujC3bQKgSCDBITzScUZgQvY5YTe2J4lYlTBqqY05Ux4Igm+L
M7s/8HdEUa7GGbrr4CTAOTeKbjZLwOgB9hFAOUOvapcNLKFTjWDMhpGBve0ADv1l
iRS+2cyjyLamZikPiYmPOJRHkIyh4JLaHqM/tY5B83NeeO5MMOg2TtIURiL4rG7I
QxSQAe2ORAfbXKp88QUjdrELt54Tp9b3IJ+s7q73AP6x+lwNPkvFK0+vN4iGG7iz
eWpdrA8KY4W962on9kF1Axe6Ird27RfsjB71MpfeuI8w4hHVmO/LoPq5bffdWnMz
xH9+EL2a5IcZuK0TEoBZeeXOTF9edHTqEe63pDBAghEKKaNPic1NJWM8d9gkofcq
ntJ2nX1WFbkjKBi7cVjJQyZV9By9nwFHwB6fa6nXY7N4toGqON9N7fXGXHu5nKf9
lgz3MkdymAMKN0mGclYTr0xud5Uf0wjHA4z+mYdbFJDrjryRCL3YRmiHRt4Y8nZB
BLmRqPdUB+Mb7ZSrMJ3Q1j/xhJpis+oYHjIOp8lx1Oo7+AlIIoJw7lWsZqlKXQTq
3OwAup8igM09e40YLWUZQz7DW5TVMGH9PqTFEIV7XFcHhUE/jVXX/hLg8Ft1Nl2C
+tbVap7g59eO5OwVMDtHgjyvjzTd0yzsmkQroKXvrxDWdzOy6Vv7aocB+6pgCBn8
04xIxiNAaTFZOtJ5Y/sqsCYYxJkqDkEj8eaB//c7xVTW2l2ORxjEYY2m7v3fQIFi
yJmDJ/855wKANlHMlWMVUWraaZXAVkAparBNxcwfWXFUdnLANVL39G0O2d4CRsgj
nDdS9oRhtAz2qhytMgNWKw0nisPckwWlMUyTrIGUGB8Pc4Gl0FVl5lhCDNZVx6t6
BFLQJzkxcWkoibfVcjbVUWlDHv59YzsMVMecR2hhVTlBjkk71QJ0S4fkOPzeBmmA
CJ2Vb+gBkHtfkohJpCE8dlzyCZjLLeay7GktN+R2K/rMyZ3R8qg+r+jPedBPpWhT
v1SArrmaJk5qrvqnp9hsKoWmeGp3zfMLQzBldSXyq/O/6EQb1UwFjkEWRDarMDpZ
U55i+1FFoiqekjBrci2CVvr6+Q2Gbik7/gE4SAH5eWqOxcSU8+076KIjoHbHVr3y
blnlOMsUPyYds/5MTNNGrqk4SPV10ru5q10tnDDOSFWAvUWV9RlODNoiIJ+A/Ars
nmYrUycoee5wQQVkmicticPimuW9++jCgw9i8MT4PAtjIHgCEAc9/uXIoIIUlIPZ
s6KTTGHxW8+Q0iEk9AKHPDFphJo43ldT/0KUzJJn32zi5E5+levoCAwqcKBHtS9F
Rdlutl/Fa6whLuNjGfeBCzupXBdoRoTDQG9Nv8E70et4O0Xk23jQzTtlEcB9DYd8
L2yWtFon6Na52K1MFkoaAPAetl6gYf6zI8kKn/wIEqs6qIKgF2mmKK+89rUQjxFQ
tz04Q1fI7EPwsbb1nQp+decItwjoEUW0HEkQa5iat64rqn/yQiYXqn/54i1zU90q
ihWzxg6CrYmot1h1xmB1vFKHzCdKiQ4zfY+w8Aq/2VLiOP+UeMF7olcXPZ8mtbUy
P8CU/zSLUmNKinhyWkjsoaSqw60YkdbIVtdFIBNAg6bmCcxztoyh8ef8hgsA/msI
7txsJ2YsA20TGLYJViI8YLZeJHmamvLnhPGxAIHTsrvJqKbJE2WhvkaPmeqq2pUx
KfwgIRHO6jPdr18ICtJrHeKZ+OT8d2Y3AkTCtMsvU/yDNU709vrsZeE5K97vhSRx
swgLVTbwYfiuBPf5pib6ytM9oI0r7RwDn/XtNQpGwUTkbd+51V2TqdF1IcgkZXeZ
fYPWemEmhUrPNzjN/8i31XTGZhOBVDxCELLHvNY04XV7l96NI0rHP1D+XAgsHZC5
8qqI/KhSXJGZYp36M7lT1if1akZu/Clv4zh0R69fG9xKEuMaoa3PLrzL62gRHyDz
nmDdVILqeOcVlfVES5Tg971aC7tRmPJdzW/rnAz+K1boH34m650oPPFIaXD2ruPE
Ek9a528OKGcTB4GvXsuPEtMD6xxM4DuMD26gq28WvrHt4h1fAUbkfPYzdbbxQmOi
E9hVIFZe2LjlnV4YkA3pOoX+ffmPO0vPoBPMsnkpOmHOvW4k4VkRzPK04fUJ0+hK
jExmCRpsZf2yhkCDZIJuXUn1dd6CKvLOdry1DYGbOCLkkuzkPpLcQ2FInSRiaYiF
ZGypCSX4PvV3iLhwzC8Qh5Gq/IV6tE7kT6dWRg+zSgdptyna7zIvGoxspbRro88y
6DrKcwBPH9G8WWfE6ksK/g8meHVssgI1ULH940yp7scWIrytZKvWldF3Gm58tAIc
JMxW5mqTGPW9Z0pfcSAThc/Bg4ZpL9iRqIFrJ7r4GLujaQebLHnWKb5fG9iIf1IU
nodi4f7Xc6dscohhm9yZsjyd6F7ukwdh4pSFuCld7cC3f4fqmOg++LKGDt/JzHMx
GfMrRtSd/jwq9OxuuMj3u38KOFD+Mo92DA1D+qiMaS24orQhOW73W5Ttc9UsSyCf
PLLLIo58r1hFt9d/VNVPNYZyZMQE2bFf8hEGC/iSBw3zHEbf3/fLQ/Wkh9rUV3Z1
PnZtNa2YHrLak8zbVvkU6fAnOPi3nx5bQu7Yh7T1KKvHatPwXXFq5wdwZRp97cqJ
bCm5MPg52WNYk2+6Lj+v0W3UFmDRwaNTffUdZySVMTkhgFqdSOPmdgx8R8vyDrOX
v7DRqBQXJdHFOECJQQhFpHtmFm9xnPOXhaBWuLGrm7+pGlLVfhW+dIw2kKepr9l+
thA+z2s0tTgixNLZtxSUdOSvsue5GhIQAO8uAv9b8tkTToDBIo1BqVL5tNRiwzUD
S87qCIR2eMOmbWMkIU05hRekZyOYGZG26YFLH9NtL9cZJpJrYxVC1X5rsOIiqfYI
eyrzc7KoT01tPkWq25cXZpapbSoYNilvVHMhEMlUD7pfKx7Vn7XuWBVSgtBw/YsU
P6wU3MRyd8M86/qv4hWrI89D+UsRpZDEQusPIvBDr0HmBd47LSsmPvzrbR0oa3/t
i1xhsz6aJ0/KtosCJJYGNFIxuMCYHyjz8fs2K1GBkKwnMHtJirhDftmEXHAXtel7
/SIx/zChBCD8ReweClXf+K+gWhf22G09gBeiRfHtxyktYtkITDJ0F5VGVCZxCthc
9oot0kl11YQolFl3s2FH3OPdOCrgnoxka3s3dtp5xk9y+PfdtU4W24Al/cF9YV8S
3MQMubhFSFaM50lTNBi7dcXhmkI/blq199QCquN2Wpl2P+MrvlRmkRlcECK3miGK
kJWWlYRMnlpG4MAa2JAXXTh4BsngGHLZrluxseyVean0YeaI5KPBztBvJGk3RkEi
iqPrqEESh8/M/0VIhMdR2k2bgeBmISz7grtajzs+DjaHF/faJ/HmSiIK+Kc+VZr5
h9g/pKE4QyMf7z+Vx4R4r6S6vkuRhAIOAOXu+5I0ToTP0hj6al4yiXV2kXhD7lns
/0rDLBVmbA6Is83jcSoJwjhi2YUwvukws+9y4jHf7J8AZD7z2HKMj2AWDGNiV5YD
ohkvhRqOpr+wPkAAEZifVPfOboZ7B92uHHDUC/CV8j1HEa3BO+TQOXpwzqNSzU+A
gu9DQNfi1c2h1gKQtIiJxlU9h7Lj+0Okizht75HPvLQgVkorLrVsq78rnLztz9gR
dZ0dILfR5PChedR0U1vaLdkl3ObJfWrOnl5xmDP7lkzI8BhTXf5iih5KkccJ24ze
eBb5EFnY5i8cctNYHiFFCi3ZG1N2nrOM1gNtT5EBjIjTmsxH5RUtqx27BCO2CnI+
QBE70ykxDbjoqVWpOj4hJZLKE2ooX+74KGIRaImST2JOZQUBEDLoq/sjnGLpPZxX
o/GKBdkYOHE/uMaCp5wrEk9DKHDEwXijvn/jnu3qmbADcuep/GcjdO0SGWucf/Ac
jRQExe0H2Dw5hYLaJDxOUXL/KFp9GdchYgpjxEu8XMV/KEhaMxbR0lzxvVF5QVCG
qoSJzX5Gfq705Ow/Y+m0TrMxH9dQfJYAMHXs3Aw26RtgnLVCgoC7uemOqePxTfQB
cHNB3NrIZ8lK+q2wLGCH37tgtzMACGFs8Zh8GbWLxZkdMj8RU/J2gXqj21NvZW2Q
whiaung86lwpIJm0oGDKNBGfLhFJ9VGc2MWc5PAsskvttKuuOmuJQKN/5WRMNkSf
ZOAB+ifMQ4fQEZIhMs49uFUP/NopLbUS5hnyDu8jGgfDorrgywK+EKJbD3MQkf8C
RaPj07KzIXBoI97UMPS4Mfa6ugIw13jvEBl9/8GVFK9T6YhLBqJqhJCHHSMnYOjd
SmVij62IjUDavvR5wfCYVpnkL6gIrwPbQRW3dX/4Gb3NSm/cPp758TNTT1wq3pcy
NGRD5+X1kt7qwyC1L+M7nsJrrUdpqF4aj5Xhlj1Ze6GzOindEZEn/kqmpYjBYcMl
0ntP4EFCX2pM+shRUq6kW81cp9ArGvo1u7n6BB9GK7YLgIc7malmwpRP8moDFBGe
/7hvJpULv+zFKHzx5Pd468vgr6ijLYm+hGfkdkxG79JQFcdXV/3PWf3wY9Xsu6UT
/XCzfQkAONwRX/W6fVqiSfPHpOQSBIcqPrCcocAqJjdsnwJJCVKfzKhBeSwqKioy
E7LXdvJgFDqYldzeX2eEgLs0HpHImEJwCp8oiWtUQaTiP1ii8IGlDcw5EhWLXWeK
vUicMLcK9Y6aRMvnfaxrqw8ULIerC9ekwwt71SC2xynRpR9j7UBpC3VCqSHruGw8
OvE/sXr5zbL5EbFF+KjjU5ijYeC2P4Gx3NZEn64CIgCxpx/xkVRwIUXVLZU0aaAp
fSZIdk+OWIZD341hic8oyFoWbBv14itwijPkYRyakBYPuvO6r2SJIR/KzwkcdMoR
PFG1HsCFJZzTzCerDMbaiUDrRHaGX6tENEBfj0uKrtD0lf3Msd/UcUfLgmvJajmL
rajj34VaA3XPR8dkoJ0L4LVmYYZiuo7SfqLx5M1pP/AWlaID/9bpiYDR5CBCpuSa
h6TK98+QTy9XZs2pjyRJ2Oj+1A4Vt2g8PEQ4b557539CmQL4N0SLgvuKBW3Wivw5
w1CvRbPX51J5cOS94M177cvalFUvjX+nrKZrtkRmzKAuMippoHIM/uvcE41Gme2k
kvMdzg47G2IorJwrUx9f09+Ej3E9lhVP1pdgUii7LClk5FdlCK/gxnClPmqFrGGA
dO2rsNaOa38vBDCVGs+TeOfnnXY4hSEX8uGjffYMNhHzGytKA48lpIsAC4dawxot
Lov0wd4fyOodwxqAgN1ghwi/0jF21YTz6a3qYMKA1sjA5QGrSRM03oZfkLK9V2ET
TuViiaZBzbVkc0k3fa2+lpSbcQpSHXPoexSnmST1YlxLGxfTUCcAxji7cM0GAkO/
xHrFNKFlWnnhOojdDSUbq0OGFyf3PsqrYUT90m640hrbk/RCaVuhcAOq5cyfg6iM
XTNRHIFdZk3Ubvhuz9s7S9GXDhvxcCrwXoTEB81C4E/v44dPeokR5RxO/E+/MLFw
x70DPKvV2viF+b81ipkVQh71bTmAA+3Imv9qWAzG5BV24cZLI633WO9GXBKDz2Fv
Qa1KzMULd7DSXoj0VdOwBzmD72VcH0fvSNrARMwy/jrXkDP0P/2MxuxR6eYQe1UO
ZksK+TnTq3fUAkr2QdqXm2aFvkWQsWGr0reHZABvkDgR9gW68OZ4ofe+g28PbmxP
PO/4F3uGCVrQ451aR+LXabLqK195/kD6HFyoRo2YKIryT+Nfly7yxP7ffF9JgvC8
krA6AafnBbAKxMuQYhkC/Q0zyZc+7K0HQDxr/V+JGIre2MId9a0frLXnJLwH4fR4
NKBhkXHoakf9cJ8Q1f+pMUHRZs2iUMaI3Okox6IAsTEgmurMg/CZkjdNWxZ4j60T
yzYTh8gAcfF+SujAFVyVIShQLe9352gIHpjAxngWVbqis/YKXKiMsK/CJ42+CCEf
jf/sXyXbfkHStKdd5jxGEm33XuAbUzABoI7k57YNr+M54yKkR/NubXWyNvPwo3Gu
HiB2skJFA8+FiR4VerAt6JxUrT1c41eJdImDiokteOHejjr+3PTyjdz9VZpclTfE
xWvpm8KvMBhzIIdL5GnVXl/aMmoC1ND/XQGfth0lL0U/oUIzFPx7YxyAsOEz8h1f
byGJo3eVhMhoNgxTWGuq4HcRzbd4xPpuvFx7NHbqUH0qfFLCGTCx3Jso9hPIJSxk
EdIWPptxH0k5/mRsomccjHElIiaDTMcm3zWHEuanWVTcknfbZwsTnanTjFNtbk8B
FdYA25f21aPxt9wx3n1MqRHNnAYcTqr9MWCKlUZ7uDsrkY7hufVPF57XNDPE/b4I
A56dzukdMvEQj0Qz8GqgmLfz5bny/HCgsvsOT8qgdilEAJEER81a7rqU7Yd1sXRi
NVrbGkBWZBYehR5i76Oy18dYgck/03K5LyOas2MBBa2LNsrnfPCzhR22kDdiTq1H
J7vbUqN7ZAFFPHB4ErhMihrcov/kkn9U23VE8XIQz7j0XXJxxC3fOfg+18tYxrrQ
uy2lxFbOJ4jV+glaCt9tByuUrzyv8FG2oUYvlpfaMFUy395Ld7/n49c0w/fpyz4W
rwZpaoib9FLH/R9RZx5mOCcYwj/sFMCdzyld9NNC4SBHBaaUG66ibctuhppZ75Ga
ReWj1jekYd4VqtmxyNVhaPVilEM//MN+IiXIq6CFI71eqdm0Rij1lVrDf04vQtKK
9UrhpLRw/IHRpmy7J4g6Qp1hr9HGflnTQRGmhrwnWMjxG+XDg9XfR4oM7vd5vgXC
6PEo+A+mX82mDptyzE3BmT0cUT5MS56sWCaHIPv6wuBEkXESrk3urWM/BHzymSfj
U2CVUhg5rrmW9go7Txl8lwH9MOshq9Ml14cbwWDckTZM7Bbd/vn8ZKuR9ORAZmFL
csjehYeb+GHr8nSNkQMCjvss5Q6BUZRxHuQs9dM5Pt8K0ny6p/gWT8qgd05EjeX0
fZSx+Ry8SPgAlw/ctYHuKc9rUOa59eunA+dd732xzgerH3j+ztVSqUKkN/lsDIDi
HJyUy0aiMqOd3i4PXA+wspNoV0sbUMTmUJ7gOkjcJFPSlRZ/GdmErhllJR8WBUrM
unBbKxW/YqYUpMUmIq8JSk6L1A86Uy2ng6sOzBO8SyuDOoRRhG/WDx313+aZYs5T
IcF21tfMfg1ZOWo08NaikjddoZ7iwiShCetceBknYj5DtFqeRvb5RfIc6W4dZc8Z
jyhyUHv4aLDDuJgqnZMXxPn37yWVpSZzPSS8hfcg7vU6q8tsbUaY6k9z5JDejGjr
+1y+njfG6eMKrMy94H8VhjkRFo5qzj2XIupRD769LcjJp2A/kOnw6VgeOc8XIU81
6nlL77EgKPQMUD99dKSnRj19KKlX3ZIGgxlSvD+qLWcHOCvUViiLN9mK5jOAgrNx
muH6c7nM00uqFrAXhBS2kpqgHOfEmgPE5g5PFGm3tTUbYajRJG4iIbP/sEBUYaKM
ceOo42zdv7FX7KUq+zRg0VOW32y0UHiZWFuheF0w31c2gaHxPfn6l4JumSiLoOG8
fwaMZer8D8EQQM2hCBUWlg3g9eLD1ge+gD4BJbnO1B8s0poIIILs0VWbbxBdWPWG
qiEyu3Ks2zlIojmEM3f3ArUYXELVGdG97TwxJ/F98aTD3ZO+71+0gaIDq1B00+SG
p1HEJb9bUoKljaZZ0J39/61/z6lIL2cTwzwrqwM7h8kwjOWBEAa//lga19pimrUb
wSkAJsRdMiNPUUrRiCmAqbUmKcphonRZHlPPiNjLQJMG12fIqKbrtRJ8De4ZJJkY
0AzwB5y3UqP0MdcDQyrCD6v2VtxIAmt9HMJxvwdUSYI6ekB+qgzrmXdE6HPvgtuy
ekqQhYYKADKYPljjBvvjPFJvak8ouMKtrN+kAk8JATTLcDO6YJ5RehiMz5LYOLiv
UhTPoo2nOvuRVPjC8Tv7Om1BhuTpQIhwYXFBurHheXq7QYaFC6KVI+aN+/OWoIBw
5sA4HHuxrLHLfJbuP6TzVV5cD8nOS9oWJAA8ilaPeYZndz2bW1tgDIoDRDWcS6hH
x6PFRDM7HHRfMIrvDucjAKSZW0tCW2KY0NqfYTSR86QSGrevz8U5jZxMvhxPLfN3
NotD5T0YlE6WipJQsa5aUpm3KeioQHLJZbhZdtX20pRYxx5hrcz9FEb9CKyPJF5j
0404kkxH3603mbEy+TPTpRUk7a5twrQCYH2vdvsSQvZgMomrep3TIASgg3kDCSQH
wvRLpZ0yuulSp+GQa8dzhQSjrIsyWyv7gP8/KNenE4tuy5c9aIu6WfZs0XyzOWKR
qyIyXHKFFG76P3accjzbMLdF9//lXolvLiRvwXn7kJ5FJ4buwhJnkkBMh9QdQp4B
O+XWx1Pd2q7SkbyHP9otOTawyjiutsmVHSmB1HoaxVQ1KlZVLBdMSKgmwU/HFXV2
3uUbfVJ9l58DimRlM+Vi/gZ0gh/3LmVUsWZpNWxG5GV6fuvpbjWADWJhx/HXMs2h
zgWEI+aL+v4vg/1p71I1gjKHHyFE06ckkQauO0Z93Telj0074gnSQHBRcLsuQxu1
65kc9LBkvwk4olz51eYITmYcDC+/Gkq2OyVK75FO1+kSloV/xT/+8QWGVPzIVsWt
iaHSJrXGtbyfv/9xF1F0ybwqXc57BErHbKRBI4vzj9SXTTNdEFu2sv+GQat0yzMo
gVait894ub1MU/8678qvFEcf5CxQUQDYVSQmPWl43a1KbT4aJTMoVwX7CJqG1KTS
YyLX+Y27dbIxWZbg9d8OCWrFhMRBeyrLXqoDCBN4bKLwn1Ec1TCe6xLcLj9Uv99V
c0td9tcEwKWhtA4hG8InCOlnI+3LzFy9LwE6L8mqMpCLO1Hhb101I1Pltm6gQ6am
6XfBl+jk3nh+lrA2Eu6qeSmxSz3PEYfdfDsnavS3hNKAiESSd3IObQqlyBMVBPkm
RTOLbAWo9qonCPBJWJRNuu7kQ7SjOweFeM31CTD5zm4Ll40FmgbVRNzY8DN6QwCw
aj6DaTLuTCDaacWCZ48vI+S/5IlqQH+zWBakOa4FMW3TvkE/9O85Z3Dg5MYvi1Ln
8b/K0rqzZ5Iht/wZ2F9PWl1i7vNrnYSR3/PHcO3txjI3/vDi6H5MEXpFe40mbfb5
rMDvdpZVCEpwA7hm5SLt7Jj+r+NGZVslbkPKhy4sZkM+hTZQMkG6MWLRHzX+TPL/
yvmkGK9fk9UKh+3yIwJ0QCxzI9dGaxrpJA8VAe/fN54/2tb71gmLYzguW39Hf9zC
wiQciRc+6u3/zX1gWfNa0VYPoiZZcCLUsV8ZfaZXJJHnRK81fcQIEWtK5i+gB0Mi
QXgHXNqLWc0HYBZ+Llme+ZPW8bvOyiShm9f3np60lG+rhBAaXQI4DqTGUON4rELU
WBnLhOkUYotqmAqJen7hdgyOb+ZAj25MQwH4IAMvNTqjyjjqlD3wZ3HqpdbRwGDL
mVImUI1aZW2HspoDOKUCrPIHZQKLo8yf0XGjNDQh/RIdCGZzwfeSF8ClXJcOyll4
GRA78cojIt7TjKNIh2ERQFgw7VPmNFTeTYqDq/7MNcxFIu8CGF3L29KB68Y4NxJn
p+8aPeNrB3QIRj87CapsAg7qXNsqS2X9IwMOJKqOyHhVDR8TZa4vuvp+quOU2f5Y
zbNwobrDd9zhp2uTNXR5Uq6GIkv0X+9Gk//YCalp4M/ToWuPJhik8KCYFXt3I3Hc
oGyPOV6ybEyGxuC1rfsg38QEjtiriRL8yif9l2H7VpDF7JmLiOsEtMxfGZKreVkQ
tkmR+x8ano08aH45S4G/wwfcmwh3C4Bpnh+nzemnp1XC2vRmB8UEtp3EQCp0ayBY
FFtgcv8+ST+E83DDCfsa9RGVaPZPSQpaw0/12HIoqcdt29xH298MeXF3zOmPw1Yv
UtKqdVVneefYJzMnn2mA19u6LopswM7oaIdl1ZtZgCezhs/1otuZ0JHvLNW42Xxx
rBHHJY4g7mYWVEFmCe9Pmqk/Uy53kIwbtBB7B3wXOGPpwpvGd1QOQ6JzMdw83CM6
fvOHUxUR+LTze9z7VsyVA1L1Ulz89YoSFXi6ZrDBiIw/tTMxpvwbDOrSEoQTgNmH
hBs7cO6cjnviETvXqiRZv5zpcaebQf8LfEKKuMSjwcd//Wk6HAsEvViB53YYYKwL
MckEMNXfnY1TCHdn+Lpqlczg0+1NVb8cVutedqLv2rPhWv99sF3EF2dERAlZJMdG
7K4etvuNXZmMC9d6ZuMd01GupIWiarxOJLCv25DAk+KayfGtgRMfbH1cGH/KyDpF
HFXTZ6UgPFNAQobvQtODwFfOMGcvnJepRmICntHxHeAv21iIT/za0zwEqJCxeRq1
8DIL9hAQbjjoeJxCgVEIbiE17yLbaNbJFocDQgc2XuKynL8I20NjO0oXY9vguccf
8yJcKkj/L4ug3X1V/flasdALK+4eNyG8rMsSTNa3p8Y12MqSdkPuTnACnXEgycZ3
CO6UBTd5jCNBacg0cjXBkSaY20MK9rXivYRAdXuXNVs3b+pPKT61C/zzkL3ubqRl
BsKprs1l2Zbf5Z5SILw3eKI2h8xaX0EBJl9H56VeZExfk1ET0VE8WOCRz3rxVHxO
Ji9JFcQC1ajrc90rN7VKp7Fu89EBRGejtwAbn99gnhd3stfhZVycVFEQGinN8WMm
U2+SeiTphnJcKuo0ymqw4V1pigTmn3DlaN5o5m9zTc3eQnxknvEZdu7Edo6lhRoZ
er8jCPl9DEeAZ6IzWaeEJgV0W7VeXXVMoSpFLf1jWE2Pk04cY8xrt/Pl0M/XkSnY
KYZ+4RlK6PbapoI0GNDeXl66/hG4BFoYxOSEaQOoNVuaMwKM605UioBdJccjEQV8
A6GVs1cFMqE3ehxK4ni0tTz+iE1JC19mJPa22VjHn4k1ThP3zGTHLAFv1eK2y7jy
VMHw21Mhf+YxAsHynxew5wYljUgC+HiZd3oHXeKW+anwplNzv7hBSzy+Uf0hdX66
is8bQ7BZgIG1hNURG7TxovswV40M3NqeuI5Eg+tQ/A1oR2iF4bhBlOdY05rsSkKg
cIpS+HjyeN6QsJgYAXLqH5SCs4/ak7j3bUxlYBiMggszOjRhmziPsQW327TlSucd
HDRGKLff1f0brKE81JBJtvCoXoAy96CMsezI8BJDRBY85QZKUbwtipqfOpbR9Myx
8xm+tkEKyU1lxPLX+ZW26QIzmBjwGa49SANzAoxoQsaOTA8XUgLEa4UqlvDfApPl
Tc2Gz0P1FVKPxX1NyXzeYmTyp6DSVCPHiSCBb2EE5/zKcz8F5XuyAIEA8iXOgyH6
1fJPfgoXuNxqrIHXOspVxRBkQgj06JEwGSGsvlqOvtmTHCJ0Y/ENU/X4DOy9JSmK
OP4tAft8G8ybMTlobVJ3ayzKOCrimdDQ7Bmne+nyfXwnt8GYcXm26obeRq3/+BUl
syC7ArqD+fWBgmH+3GVTCnkvHW2QR97ocSLuJ1f0yVZIU4pjt196jARFmRzQaMLD
vod1OL1FeAdDxnAUmCDHh7aogVvHWEvHkP1JaaKWCY304IV7sHaSE7VUO9JxWdXC
0Eggoyy5eCroDRF0ceYEgTf+o1fgUZxrIe+ZQ4HV0CIVGCZrT33Hl2ajr/dIfuls
77uwZiRUfek0FTLoUOl90dyzYRE2RLc/bVKHhRG+kOOocGsO1xAWjcbTpunyIHKu
Lc9n8Qk5dUazm85kTZPfbN/mDZOmquI1LSvys7AI7I2gwDXIs3IwapTuiE5TFOmH
kKXN4npgWzxbSWWZ7wQm+A+IkZ+KN6mJlYIBVce3amyTSzn8MD5BCKB+xe1encHq
gqD+UPF2+5go6wJzUnTH/qTm6qyir2h002/acL182kpd64LGvwjXY8P2Q7cCtxma
NEyld1M29RFKXmyuf58hdw0mof2eDOTNyKD919uhhkRsU+88p/D4/r3Sa2DmB/Ei
R/t/ascn/agi4x8USEyy8hNeFfe91l9A6RUsJ4Yjs/qGUIUveuOC4tOo/Cre5GMh
9DQuVs3cpAQs5KHR2+38/A3jRJGYmkS2l13PkcIQ/XOeHpGykXedwwqKqJ6+/oj/
nSk7/ICYeRIAlkZTRGE1shhmgdo7nA38wVUjtoIWeMqpXNv8A5nl+ienHb627gMp
EL/7Ck23BtlBvFH0jc3BiILtTqg59rmaoVKG4hd7PaNZ7l2Z3vQc196VtUDmC0TM
rviIIO9wMbQRJEWuhi5+hl355BMzpYZYnhnwLnzAHNHBa53gUUStN7dK4/dhYuiN
Zo78nDDVLqf/b0K0gg7fR0Nn7TePEvwyr/26pNQTkhfRjn5ui5/Fxr4MBLe6tVSa
MOzqaXplomU+ZadrHmTlKuik93ZvyOW+pXMhZRjkKoIDQJj7yUKHjw2bnc4UUeQj
AQ9wpmwes4vqGJEBGydUBbrsQ4nHYJexVIYwoLs6lDcWZuaAvFEEpdk4Q2ZuAUuu
P8OaD+i4b88jw4wEiCv81be5hNYyEDu290wx+N3G2AqJujsLIV+u1aDsYuGnyp7/
L7/RMa6ERkvI8pyjwXp7Qbcr1DXixsBDCtnlgXW0jIFFbpwNn73Hdn4Vxf48gxpJ
A4SoyDZ0K22eOzYginYasfrBrPu7qYcsyn+V10+Ey+zKpTXNyOcKGmryk52nLj+1
n6g9IT2Kf34V1AmO8Jd7/4lAOkXyah02PmqRf27L/gsV8dHyYKJApqBo2mNNRy0t
jqGZZLN1ZRweHWXOoPQr2Ecbizp5l2YGCHmPAtiiBn79VaJaehYKUfoB5vPL+W5D
QIwf2z/L8oGJAjITESjQXHFC24o0rl/eup+qqzU2B21rDJ2BOZIWmPQM/sScyRdq
cDFgNbUVHiyWXiivUsmenTrwqOZP0TiuU8mSPDW8UZgqpCvql0QBhRQnL9phavOs
4pTXjsKn2EJbf/z5e2AuEHFW6k/Uua3yBsG9zK6dAKLch5MEJAUI8JQweZUXc12D
leBpYoJK+T9V2cPd6Zs9d3Rz/w8LXQV7/wkollc1yxh7odbNFZmM5B389UxNsQM8
pLdgYjdmutdJPVpdSlBw16fodsbYp4txk1OQ4oPnhegbQlrtyKX9zNlDXy3sFEcB
fx7nGswjMwyi5HdOkKNmp59AWZgf+SBh+ASknSSDoYHAGh3g3HnYOSlaQqpMcxRN
gIWhPzHKyktXhGhcR93zhoqtunk6k1FEuTVNRunm3Pajv6lgUtT70wZmsNPdy85H
7E5MVdP62pwC7XHp1mexxEDNxMRP3ArWTq16t2kLiOLi8q638UBt6BumHh5BnPtu
HIxT5B1ERIimLvwO5GxpWJeZLuRMLVud07EK4ZqJ5VN40DjyDzDbWXP39xOb5Kqh
Y2pQQeebWeGKY/2B9XDn9YtAdNXNEGuRwnkg+GI6gmpkcP+C0+ACPtWrLXvNDDG1
9cWjSG1H3u8BnHXynW0RhpJcPBzN6hD7JMOI9h80AM6Io7FxWYLTXKWVURHF0RKJ
kOSI6uFBHSg/ap8Nbm7XdCms52FS8OZx8GtPrBtZl5G87Pe1N4n7Y+Zx/ilQiRgo
FKHr1OxL/KebP/pZOZrI67L3kNYsLHFnBqd3/B+eVT+XhNqSBIIDUtaUXV9tCDQo
n38HY9Lr2+TvbtxVtjI057/J2bb2OxmdtAErcbtLJt0WQXU0bCkeTesQGTOHBHId
zvkPIRky43Gmwv/11yWnKylZsyfNXNo8pfFsJ1gNIKvKd8gcuQIT3QPuFWUjk4DJ
U3MgHFPp8iuyv8iEKUGoS5G5BvpZWoeI39Jttd/N7PH8uqxIWHGaNwQRh/ZuWxdR
3qoOiOJ/Rb6ZMLL1GpfdGGNXSwm/k9OPx4vjDjNJlg8aH3GDWFxUpLe4Rzav7HyE
sFDnOqCqZtq+Z1G4eODrrVu4T+MijeONxFSUmxqslxIRP2tmfdGekah78XYidJMp
LULWDbcyKwPWB3gDDyWPLVInspIbvHJQrOomhGdAJlceL1XBvq7jINxqOL5oOKcD
IEFu1He4Oi6q2PYViCpofMHtEClsKvFn/sgszE66khKoh+Vd5rH3C1uVzftpapFz
1OfowLL4wHCetuNXKaBra9VUXw8XoDtJsQUg5OhYPMvahDqhf69lbYbj9PjhPUEZ
eIjLcPOiqsgeODwcLXE6KT38+9cNO2ZkwAzyveTdZwRBzpu68lotqIQQov3AIq/H
3P1a+4cCcPl/lL+ozAtjKSDBS7cCc13/kiDGlBGBbY4pRDOyzQI2JDbeoWtPVfQK
UAw9Og4nVG9aTyQdCfHCLHp3mYVXtUBGCRVkMKVe6zXP8CFBKyFhW2QAnmiGC3Gd
mqasZ7hwVwhb0ouVoX61XEkaBAtNpxQOznVjJ+fgBct/JLHvJ+JqvnD56whUM+qL
+WNCSoMaHh/PfIhSR9v4WQPfdwpn+zYDy9IYu5Ih8eZaKRHoR0CzANzmRaTmk1i1
sXMg6JooLKS0Owjflo9owKG+t8nvJ/QRxj5p4BJjDUL5hN/on8yFOxNgznQL9AE7
kBOExNR1gei73/zz4eTksdODqRL4RjuiqLk9DgKJuot/bqyqqjphopEGqNMiF2e6
WK9Hm8j7uhDblK2oE1hILAElbKs1STtCkTIyf8NCQBPQus2w4FQySS3dFKUCAN8O
bA2eWLZYEr8dvrUDTM3FoYf3c8poUWUtZdKeM53xZ1K79JEUXUecBaxSlZdkODnN
WID86fDRjJtMi5mi1c5SsHBfC0i9b2AV2gIGVjJ16AXDCSB8jlSP9EEP2/Dh4Etv
oqPFB6fi3gfgq6VD4R1RAKuxlU67daQmkLCb83rCEATg4oYTI0LiCSV5NHgcDANy
KyPfodfsQo8RTvAr55h3JBRgaM6702Oj/7mol/Tb52Nax/lRouZHBEw0jhEa8de2
/KXgWrpjRcfchCrNGyZ2bDPMfd7/0FPW3fjtlMO25uSSfA3UDBRC4S9Wp5UFFpfL
mwIwDaeUZh9Tabc3HSCFUdWuoMSDJMD0tD8rhhDDkd6klJXFtCbnANtWrixL4+kU
STeN/gpLd0Qxr2wiUWI1PZRyiDLqJsJrsK1XjNiqnhxNvuxVsEmjdEitV2VR3ZOL
FmTqEwri4yLS+gcfNU3id2HjQiqlOvHrJH/Ilj0FUU/SqDeifgYUXhwM5Ve/D3ui
GGIBjqGa18TFU2VEQ8pMVB/UUgVieO2ayDNn4/8GYa1E6ymvqH6dUVFMPVpPzLQz
B9+Hi00MQXAEfprcxQpFdxIANDqxwCLIA4b/hXLu7lI7vuUN9QoAUP+i8GIte+y6
CqBjKLFnUsAtgKbqdenunnoBfk+X97Vjj7FvSX+3gmOY9GJi4ZgoapB6Qu43Ksiy
dqR7U4uOLu2dyChxEuQcLaFhYaNEKKY/2IK8z7YfKiuh9MwwK7GqothvDdUKbxfh
yNc/WtVgcq31m7T+M1Mm0T6vK3BzuY7nK7nqYqpoB0pJjRQCOaTY506VU4ufvZMK
PqLgpP2A2B2NfyiblAaHRYps1d1+/B0213Y+hzZmQfxkQ+nwiQ2JT2CvD3UX4wdj
hq42abaGDAkKo9q8gurl6v/CtZZkWMrHYnRiJhlkgavTEBns3sWVbyKxYgJxSc1t
pMYzAPJb8lecUec/Czme4mjZDqzeqRMI0zJ0VS3N0gGu5f/YOSAXhSC3jkBI3TJj
AQeZA6ek04h0QzQxPKYn5AH8sD8Pi8yri2yJD5V9sszsj7p9VgFSTpsmmoWEqN0a
0waY1fzfjBRyKR2/x0cJj+k6gDqsdqfH6iKR4HmZt8/DHsMhLJcbWGcZiw6J1DE/
86higysQ+O8VZKqxlhVg0YQ0Nm7kN/1yyTS8reFU9LejJSdRMjeXQfiAHLEM5Ckl
yfLnln4CnLslDEg2+X04pT9TgrV/eIDtRR2bUAe1GgCnpJGWcZDLKMZBgXRS8JHm
vPcnoqpY/mTgDnxHTCe8iWoIsaRNz+Oqzw+nB4eMgsmG5i3ZLuMLJFHCV62Ht72s
exkrvkOhw3OcPANlvRSoQ/WFoUvH6xZGjKaEvzRq8vHmgnT6N8syHgkbpIE9n15k
xtodXAOQai4fcPLnwOarilUXPwwfcPn/jH6reerQZP7gadsY5mrqK9uhN4zsjBib
MJv4wvfstIpp3HtCtXSFpwFimv4L/2rncsub0FZZ4ta67qDJTfkCOdzaJssSQHzH
Z+Em4ugW/ssh8FWsYgchtqryJbXBDpKW2PaQxehI2IfHOq47xbNCt6NmYfFDcSpv
Tu8FY//SaGzmeOJSkyyhCzLRxsROmLF55aiTC7xcOv+CtUfKKetnLVMS0WSCI6Ky
s9wOZMA3I1yLstJzP4GmTYfc57npoHA/FHpzZFTFIw1CadVeecW1vRyTc4o9C1DZ
hTQklGmHbDF/6Y6i2fr2UnRnMKxDowH7l2DF+CzYEOSAMgvCVEa9t/3fk78nUhDW
uRsRR6s8zwbCvttZVeCjshQ7iBPNIwexng9KpaVSY5cW0MsuJBS8hwqjKIOxVImN
kstT6A4V7vpwSKQlvVJiW7nkcJB5jpzy4WbYCtdaZqjCX5np4lx6Ns2cXhATCI24
4llbiSf6Hhj74hWFvlwpouUnDOnau8s6TqmR8+LSpm7I/rFPCzg+7KeWo6OldDtj
qBQl5MBU2TV3/5F+/3BbVbyq0pDwUKPNX+1K0zUgWqmgZfZ6Ih/7QWYiWSM4GLMR
TL9rqUf33bDWs3/RENAT690I5Ql2tflBo9ot3BkdzK0zwDY2pyhYIiBDGmfZQ6tb
ByGckul5JCsXUso6MmjOHU/jYR5KUA2EzmuAMHeAV5TfJtjQYR+XIF2d6+V1rVwB
qYMzZabdHMVX6EeezxLU74I2w2c0VmSRkCyTt1ggbXoX9DdcDbUxKOKEJIbYah3D
R00LSTj+XaL/Q7U+Tu7lzNr5r1HYhe4uLqIGlx8BOb5Jctgl/WqTSFNbK1kGyfT2
2jrrSTT6f6apMu4vGT4Ii9uEaNCq1y3bLMZmsJCcZxgPywWDDSZyjLLro69t3Fm4
8guTm95E+mdW/aN2S4zwcQPYIqLr+ZjocqMR9g0T/xP7VovxWplGkUGtH5YawGiq
8BG0rOuv4O3j/cf1DO4w5o8w06ueV+XpguCR7mh0z9K4EKLpUb3eW5hwWg4ra6CR
6vcj26XKAMa2zXC0YpZ09mFacqdETONdfvCd5riYc2FgnqaP0zt+Z/AaxrwiOBmk
SPvlX63mgP44a1o6AIAG4RrEo6GI85SwptQzzDu38by92is71VGDbiOYQF4VXW38
R+tSuszb5ANfkYvYB4sCVG54Br++LiHr6S7G6nRKXa1O34jm5lq1lnONqvZX5yki
F7gc022dHw+KRBfNt4uQfcRltOFFadIRVAonlMM4545rZTDE4TzcTTMTpnJYsdQM
hxKzfengvucmCnKAAD1Agv15VdqsHjzOTL/X0vJZaGK6R8pgnGwUxriE9uN/C+YR
ZC/ELE3aHC0zxuVOV5Le8BDmF4DyX9trcK3vX2EMJkSmMcYWFSvBqqveqHRLkqlt
OeYN0v2GFbLl2Ad/9A9IGk+ux0Ic0yoOwQXNvkXcYpvNXuqDeer9IFddPS0VBibs
0oRWPWhtbrwyp4bxR/ZbflQV/chRrQleoWSDKHI/AVrsNy9QBT/x6Wkqvn9sfUD4
VrOM2qXY5HykyBEKRL6Gx4S1S6m7EUFVNATbdGD0uJr1t2M8QSlOgCijSYtZKcCQ
yyMjiYMpMuQiGe66LbtoJFbk6gZW+TMclmwT6SHjlRxSQ0ke5rU5oUpO8d79FRc5
nrXEl/mcYS+HxWMeU7VSuhc8U+jhyZKmXnRFVaQ1UriiF9B/RQxeRZkFl7IM88Dk
0rkgVTnjx6TIW5mt155QDX3rUV2ILNLfdGzDrac37PUrfYn14Oy2djY5YWl1pyd5
pO0y35s2psYJOpQ0THvhUzcVaUtfmxub+3NbxAaV0AErIiqQFTSInvzpXhKgP4Nf
tcbdNC3Q0eekgOEk3uobpErNWNHmOJP7TknAxHYe+DYdSzXgSjevXalHsiO1+hjX
1vK+EdCVwgvd4c+5u+V/e4qOG4vb1f8IAox9/zNYoQp7njymlEpmaWCwzIIm8oSh
9HM3/4Xi7CQ8JcVr+a2h3cC/mwMp/mefCu5CHnlUuh0CBIS4m29ZU/egihBsWMuP
PTwxIcUrKod4ks6f5mSSewzYS8PvvWXdPCC+bVoGcQ0EoPwiF3a6t6HqOeIq3P8L
lN5a2z+r2/P1FCfeST2gGpZku2ltamK0ppObnNMJpKeZfAJkm0LSP+c+8Y+wODx+
K72wUlR5t6+1G5kHueStn2cZGdC6nW2IC+5A8ns918Hw+lhftkcky4rj6M7w1rjf
zmdX9wTulf1MnW7rPsgV9zFztGNy0x/G6gFW3NPLfH0gUFhKaUqdEMQwgSqokWWi
9aD4jiWpccOkqoTgCt0mjouGJNHVtJzoKXyGu8yI15t76MOv7L/fUNvH8DZWtfaM
91lnB85P5kJM0qiOAgWw+UOH2yLib3kcrgTn+SkhjpxocvFsm1NfKxrmCf/08Bzc
y7n4ycfPGPSypIgeosdyh5kWSShZ7FQlIUHadVVXbIsvLX+133mAD4GclquD/g8J
5yBiqZOPKczlUUH7bEapwrF51jXD1RuAmu+62i6v7jE6+6yMBx165W5gN33qN/9M
mef1Ca53TYGDGUDbqN+dv/FG9FZiIpC8hnITc38cHWv37MSpEhS1N6estaNGsDa4
mD76gpE0ltZaV/+zWmvdtBJ2coGaCAGwtbVcv3ijoCuv8sJVU0E+c2ekUBKk2Ft7
Uy7Fgdkkprs0jrFmj60MmeCT3JuwdJGSOsTKYu/7KlwHgaFhX1HehlTxzpz2pV0R
CpAz8TqGNNtUvmqdoveYLpSxnIfvOJT49xYgLHDB/HN75nUMnXEvPjxjwEPshcag
wru8Iz4H7o0YBZ1bTl2fdmE2Gp7w7C1v77hddonE9vs6ainm8+JswaT7Xnp78t/Y
UpuV0Pfmn2qAgi7H+k7UQnFbe3fpqoZw8mtY4psC+Wm/abgZFnTCMJtGBbcyylq8
jPSSt0w14WvqPGXetxEagkgYRRLVuZF7KvbVm51qJWTARSqiTXKE7zEcYFJ5vqed
Px9tlp5wHEhmndqe4/uzDVDmXZUmQH9E7wM6G+Wmh5KFCS/Z39EA1/UKgkgqaSBK
rkLXKOkOsPVTrwx7lalFECE2wGmIXeSGYQg5agIvh9WxxwIFLIQUVRBN+ax36Db9
f5S4wZDuS0kBJmGxqVPEBnNFrvXINsyX1ideFWv3CgIVuSy1+b9ilGwZmjlEUoHg
eUTGeSFmjqZ3AcLZpVrP8ULmMkvD6Sv0V44p+5FJvF577NMGz/gZ4ikfBtd8QKFe
Zby0i/McAQn4SyaeJPGaQSyDeJsvprsochkExKw/yFq7El2OEJSOk4gGOFTGJhhM
wCHFYgRmIYuR/I0Ud9DbtlCNxhn+qhe9hO2iGXE6VSe7oQPxrxrbVSUrG9g/ggNp
0RrR2sPsr7HHqGfQHGMM7HD882OeCWKPOKl3NUGAXXCcQJ+MQyMBhOaqaMgKAZL7
QwRyihhCmPhSG/XfNTBlmBvjx9+oifkt9mZMCSzDj00n3y5Z55NUOXNEbW5fS3Py
1Pknis877i7KRN2O7+e64bHrmSvVc6Z1Df0hjx5AyRPf9ZZ2hgGzySg6lxpe4uUF
U1GbhfvCaUYwYQVdDbHhO4RkBUfZ+19ql+Xh4KH8t98QldokcZf4S6rxiSPz+VCd
iHEXtynCBYocSTBCpfUR7ZpKo8ezaUvLlwkYu989NKNgd0VY9nyxv9ol3pCKHkrs
bQnK4PNB5LBqV4mdB5cVHP3coSIS5f6bx+NDpGN8bB7oB+zQnq/JzL6tkITH3Gdr
/cshQQwn4GykGGfsZ+/GDH1Bbbm8XYEJOdDMxRbRLYXsQ09xJWoRhpbEny4zZeDd
Ab5eEKFv5s8af4I8qkNOZPybDaqlIbEZL0eXhQaOS/D+sEP4mx6oJ5KqaY8w9DeS
w3yM/wFBuW3K8Rqq6Hcunv/YELPoUe0f+eSWl9pmM3VYDs1/Qw1MUAbTVGB5FEzs
N8zAgCOdEECJDb/Pr/v6pFHdBDThhaaAyViKTwbFfDAsg4J4LxzT+4gej06WkEyl
gPk5YBB/o4FZ6OA3iDYNalJ9y8P+/vODdYKlyXZbFxCEz4XrQSHg1aYcDQa0OM6t
LKnNuk6DpB46i8tELlRmx+c0HsGOCCMRzqo3YXi5rVHMka8Dp2YPt1oYxjW4BYHc
FD1P1oHu/h1/zHimLcKvsmGAEb/GrveE42lfmNPVDo7CqTc//Vnz+U3eNETWpCbG
zwE3+ZO51HsP+sXIo7BPy10EgfqmCiqtXJIJV7bfCSOGKf8NrbvqfAr8P/GRxDMT
cO6a09o3hVKMTK/f0xIQDjagADEy3RoAK2ZrN5q/h60oggsrl9bwqMCf+Ugnf2Kq
Gkkw+Z/ijewkPQ3kHjiEgqLTr0WFkGt1eX/RRZ+tWWGzAdtPaYM3yBBdani30caL
fjlIEUZT2lzBKhp61EXj4VzsnuStsC60gNg0NLjV8ti74txomjJVgji2ystP2iAD
TR0UanBL3kQszALcGUfu42VZuEPNDMAWRT4ZL51PtHLgQUTqrXy/7U5emCE3s5Hn
9SLTsBtFbPuoJFtuDIWGSk46dYfH1wxtS1X1Mr10lq6HjmoMGPGR5AXIAdTA7XyR
siI6OsD/gYe6xiPNj8gyr+/JRCNaZ2jVRqLN0kywgW7aYaek47gfz8cp77KnPfiy
+5QKUFCGL6eeDSAo7EOhTpuLwQSVfgQCthQxLa/neqcC9ZdnKrmjt3JAKi7KYRCQ
jU2JcPLp8gHowavsxMsc0WJf1VROT/9UYPQN7oBr2Lzb9Fu2n1eszctNQYf5WZ+R
Co7Wdj9W2tbVRCBnNu+wWu1igumb4ksEFT2TmVpWm3WdaJBhnyixEwv0rV/3G+Rl
Dt3bkaOScxxnZeBhLXuOIuEk5gfttD7tVZ6nYlIflJ/aGp44yK305ZGECRyUr2F5
gm2TjUjKQW8zWKnbjVvNboUx//E7+VQZMtxJP11hCRJK2rbWwO2vfl2ZGmflPYNk
NtM6p8QsN+2GxpOTWqQMjxOiY88YgWNYJAT0HgUvbityIy9TahwXxfpBmMNrmXPL
HE2aOHeS+FkUwEOgu0xay8omoZ4TyoJ5/fzKawUU5/SRATIrtGEP6V9bZlxzYbCV
8RKDmrKodU0kmP6l84vEsw5bRnNLzj8mKYawK5v3G8uW9lfoUOKwZxtkxpKbIxQG
0CPRroOGTCzAREOS+1wcbrvSQb4vGMNCMFfzV5DrLLN1AfS2g0M9Bu9ppK7l6XAP
vKuOrzxqO9EFzqPHBL9QeViHarKuyHlGW61z03Ylswefpusn7G763EXk7SF7bm/Q
9cuDFdxbptY4ztI8yvF+wCR4HoPu+wGh3SfjjHS9VjZONw5t+KmLJjwZ41V2R7es
li0LeEYVXn/Evwo1Yd4IEfJuLFaO++ZpUt++GCyeCGZBocAk+EN7qI3UO1SzTbiB
2Zcswlb0dmWoPyblJUEEUgewZjWIvFCSd9srmXrmI+otQyr1C8P0nKoaJPQZx5/E
E8DXxATLxxsvQvOUAJkf8V4GxBrSYLeOkhhmok1bojOotHwpW5jhgI4+AXsGADr6
P/+vFGebHRKhuoqsJgC6qLF0lkDq2aKuj+jc88HMWl+jklkSQ39cLAPIi/fzP1mD
ZeFfxUrWQ9PCXW4K9N1ZGpbKXWnB6I/4HaRO4NE63SF2x/riHBd545qAz29ECa8e
4HvAL8qIflR4zhWE0lAY6Tq6MoLZULWbDG3vvf69OFTNZPNGyvrmrFgR3PU3PYzc
en5MLKlLS0cFMSDVRrWsSGSCYD89W1BTyNmNizgCO/LSe5ZSIvW3E7DYnYR6uy7D
fPMVjbxpL3M3XeZ6Jz0jIQcJeblgcHnRw6x6gZqWNW/2ZDuu/872PfAQGPfGHCW7
LMWlQujuiuouiwxATRfYq6bFbSYwH5a3xjvSd259DGv2xsejHjWSP7scqnOq7woB
Vs9DIBMdlKTjgzZVsN/ZlJ2N6nPOv/8oouGuBCLGddztTA50eC/Cp3wnwUIN2bUK
MIznEXyJQTVHLpaYu+b5aNWF8VDbLuZ4eHFRg2tTWX+sGzSZ3nedrqBEuHKdvHZ0
IG1/aPc8U7d7Rdpb8ZTTNc33OqXg2SbHpQ0C87wkRUzSzimJZYLW1maxwqWBsO/9
3tSSujiXN+qLZ228xIKSQUBXnz1Wlbrbbn+4X2XvmUEaLr9CULPMRF6+yAASI+eh
lX9XWHMaKKm0pDT5qPDDOfb7Cf2K3WBZMpz9rPCiRiks9RYnlEElvF9bWhWHq/OY
yGRs/2cMn/FiZ9fVCWUMw4wWuknPADIgdTo9gZLdvA5T87S9pz7zbdutw9LoZKDx
eDxnGkHBoYvYTXgCUkVqR257MhXAeAnJMFOlmOSVhxP9jXfpplD6dbBF0whouJAZ
Yj1Jhi7woGk8hrw8bScdbGgEsGUMEdtAZz7h70Ut0/+RLlfJTs2Pg+/pq8jWPU5f
kcq4JhKNxIV/JI2D1yiNNuoCvbnTrbs1ySCxcAGxeP/pJgjtZWso+737CGutJYPZ
OdwCEHIz4nsWwfC0SNGGLUf1u+HagL4RNk014qRuOlhfYVStJKVhfo6VRxsalscI
6+uGbL7QH8bRJHpt2fAtkt+EuzG1Dwm+uEO6PNblCEVPvCV8ZGjOw+U8endgfCrm
t1qP+3KgZ/IZhQYrfwCi8p1TBBW2dEy6t5N6H7PMg7DAyVTJ66BNQzrDCSen3KYz
O17PY6dktj29sPWN6rQ/OqX9iZ2Mn9EfljGnFmQnKLL7jZrvNGcjQVTF6rZgYHW+
3/zoPzGnA1H6ssSVrGYNnmDMkMv91/TEeQve9Rxn2RDY946kNH7LoJ9wKfu5olY4
er8NGeijUdRD0b01RKdQOUQfsA7Xst628nWxTdW4ntAyffRXKAWFqBZrsHcAItOd
VCURNXNLxZy2uoEYO83KTqv3e31FOQj4uPwjaQ8OL63fvdpnTq9ynb1QJSwxjDBU
Ro33IKaieaHqxaerJUrxIh0gkljQgDu/m7UiXqFxveuO+Cs/JNCv16T/Ph09ltJh
PbawXOokzTiHnQKby+9ikY4x6OLCRC/9kCDbLsske9hvgXuaLHaS4tDSjdtgNCVp
x7kNpVdqtWwfxzAXPHIGYhBd4/obgi3y+5gqy5Nk2TAIBlwud8A7CMjp3ZnNB/+T
a10edn45gYF9i/2fAe6f7bWPTPmHq3OcBJ0Bit3i/pioqFBT1Wvu7DKqzsAKCUxf
AfSydcjddl3xh98b73fcj5aXsdJDcD9v8qbYvd1xaPGvfSaEuIRlEkxB3vSMSznW
9XFRaiz8wG99wf6MZk8lj8a+CRMUcu13fO34bcwgQTmvjGmfpp1LOdKMQsC5w6Ka
du0pj6HKW9INnHLuiese20A0Vo22jWJGs4V3u3cMA/pqhL932lxze8Ui63mkR0HA
YdeH1nVYZ1HgPm7GuXV3m683LAVHrT35aJBGcTSptjre1TugnosAwJsdGoNwa+lB
2i0hTYrdOtL+tYlR6Vas3BCuCBp7jI40ACMp4G2tCijVIccmRpXBfba6cydJ0nAz
rCpSxLC1GAE/L/JbdfREvDl+drPmhpLGbP3AFzbbL78L6LdXzsaqpVZKbXFKsQ+c
dpgLPOrUtLvHgeWBoGM77tu33dydPPRJGYnMSmDBNH6zZsfIkxvSqYl5bokDP7St
z1HekfqaKkdNg+IA2TNpZcabu6131m0KS5YSO1Mb3ffPWMBjpiGZSbVsfzWfiXkA
Bh+h8IqoxKtRw/6VLvRMC3rgRUhnl1K+yuisolpcMcCZ0AX1fdMNDT0OVUsg3301
Pc9Wg+C9aT3yRdaOtYlhoUJbqSFL0DNyO39m1EnHfrwMfxr4mzA1+hyE2+yq5GtR
zK8qHHLMs8AS9g4iWR/aFc7Ay5SM/U9Eb7d3Z3tAppI/5iZJhlTmnmjf4fN0AoQR
g36kwsuAeW9rK/vNPwsFBqw7D1dMKAZw7+oTmlpNNWjMyIuMktg49HdkdsfB4AMQ
xAyrSD37avzH6tXQXMpyCvWviJciZKT0iG4ioxgXtrU1SHx79W54e5nDUBjV+FTx
6I0NPHtsMBZR1+1OT34UHy986S6pX89yTYRx3Euvzo9XI1BmIuDxfg+TEj629S3C
Mjz0GEiARjnGOb8NJ6VsQiyAfAQeORhnj4dWbtLn4j2dr6JXew2giNXz7SaM7An7
6eik5oqupfRPqg298wwWNSEieO1hnFpgx2J+A8LDxFkNddc2gVSl+RjMBlggOdgQ
JIFiWBEbEQ8kJeHUQtUVJJA5jp69ohawf9CLSI82knuRSEpjuuu/IaWLBS6euXQa
EZe2//0L0Ekiqm3ubu+eCdteqkP2nMBfFfcIEXWK34nF6m2Sd642h/NiyLeshOfP
b3RFqPmnhLZqLPLnu0tjhO0LTULtztBv23oZjeRsQAUZh0Jciu21x26LCZujAbBG
WndSo5x0dGz0QrxX2fQmO+3DqN9sv49sP8Z0gW1wjVgWqJrku4gWo1sQaO3HkLYQ
nYOgRLESrQ9IZRZ5ri6JxatqPugeXBxZ1ex8QjuhZ3ncbyPt85s6B4nx0dJMnfVL
3Nh9+SCnqYUa67WUnyl27L56YIEeuKKAtSvqcFanL2eMM1WotfsnQfZQOOdD9STv
U0y2lRnz6jLti1aHE36jPHqZ9aBjIq0D50OhArF6qwUirRud/uKk2HSiInrU4Cii
xv4vKhqgVCy8AOr6rA/y+vU3EORhDZG475sMCdoKGoV8jps7eNP1WVy4aUC4YsXY
RoOIRXNrW8EW2lPJc/1xwBUuvrqZE+89BrDDYj4r4LvP28J+Rr2wQxPQHTRyH6+X
lTC0GfEzIz7CmcQ0ntQfLwvoBNMLtBUQKoHgzdziWNdwsEBgYG1mQi8dwPmK2TvB
D+V4Vog98w/e8rPC0KXxVSfgDBXbt6WB6l1unq+Cfv5w24NORdHgxezrBvcimOHR
DSYvuVr27OTn7W92q31dMYz9OAYQdA3smbGhD8Y0Yx8VJlF12MfIF0GpvxXehHhZ
vauyiJOWCszt8AyPudKatoBhTAWcMPzm7p0Fkx3LZ/IO3TXRfVyrasSAxHvNlJD+
y0pTdKc0sw08UevSJyJWA/N5F6Fflkd4fBFJy+We1NLBSotDk0kN/5shFWhgW4ZX
MnXHueZwPqmFcIF0r3ViWCLVVhejZSFUWyDZKDxo7g0/RFKbnGZGveEYLpG4pdQM
LDnRFsGGeiGoiaU8M2sZAc287HBVAw4S+e4UiCTnglNLUYUIVYXloVSZBQ70B7Fl
per1jMsMFbtbF7nAevPO002SwPVhOEchgveHysDzOChJ2Bg5F/At37h4JXyoPZOw
j8jxvK1PcK4iLw3+1bUtFuOCz5w7zN1K5dd29MJ3O0V9iRWAi7E6hBjtJa9D6vL7
czDwRVqVnEozBcXlxk060G+kNWzXGeFBKu+yPq9a/8S/9Oj4aepnAkLRByX5x0WI
MhZjxdVTwZL6PZFfuhcwkJT5uyeA81lJgZivgNI542CEUyRHM+gtzJMah+MVMhsE
8e9Yfl5htC8yAXCArjluJUc+A2OKRrGujNL8KB8psCVdW55Njdhv5WJocTzgp6kk
oCAZARHx1bUxR7WgD85djgItT8PXvq/ZbkOE1D4Y/J7bDHNBDMU33O+miskWakD1
1bTiZXK9JdxVpYSXgXqTxjeJvTGeQe8vVDm3AzMfvWc6lOTHkp3DW3pcj+YK/Akj
jGF9TGEQgls7NeHZLXVl/MMcg/o49Aw7cXVSTw02GNLW0mewQPvjIjO+Q83xZHyT
lHuhDVTX+uh6zrvRs+WsRjtpoLZQmR98FjDCmGdbXJyV14rWZZbNpZjKmybLQ/sG
Q3yw4JOVXh3u6EqNYINs3qdSkFmhoFj3LU9yeDruDTuz7mM1MHnY6XzK8JNhqvNn
3h9PTvYXULlk0wEQ4moC40YoDsN8BpdClTSmf5uz5RFIaV+iQuk2TNvvlAAo401o
EtN4IMm4U3G0n80XMCgiC36tsrdqDYurylqUC3r/WAiXSJmdKYNFgFWMWRmiojuB
kcgHyc17WQ6j4CywxI7vj/j69MrjoDIrF1mjNtkvPjhvvMTtq9xSyBgbVj5Jf42J
8LfLbRpoyeuDUCv0cc8rsJiD5WlnmByuJQgYyudz6dHNYM7l9XP+DhnK2VzgGpGW
U4mx9qsYvMVglh9+/dEalclMZGwko0Aa4pU3j7EerzoHhlyyDcepGATj4n9dn8o4
oXvNyzq5l/ZI/qZnIo1EBScd0sObZkcNHS7xv66eBBoDC198x9Ez1hesJtyYp4ap
QrKS4ERsUv2ZkGBjg4kO/2xs9bMibXqXf1Vx3op+sULUxXJrPD2RPYPsg0Ii/+//
Nt3CR4Q1X8dGbl4kXDTpMBwPFjtN4bPwfQCS2oNljNqgNc4im8neTvABI3vaNMjH
yiTzp3AQ+f2yrMPfvkLjRiYcpboibdxVx3lP+TGJYhWn4Jj4QxZoMTr8SgD3le82
qRp/nZFrDgufavOJAITVdo95DIqm2+MqHKY7+WBanb0dLCRTKaXYjok44DVtJlgg
IyvPMkiV8s+QW5uF/vRZg2VI5PUDCQzuzfC3S9EKFCp1Rnu+/IX3X8Zd4NeuQaGu
tX48ZlygYvma+SDxrS8151Al1pY9mmEawSTkQ6y+6gE1jbPHtOS/vwiR94qa0G1m
9AuIg5DISBWOY6WJdQP9AaCSqZtKAtqvuhmgNbKEI+47r/XD22y75n16LdRbvsrE
SaN0AR21hq3U3Fw/PvjvkgeJeRQLFQgyzdQyxbnwmj9ihqd6B/TTmpchtofnN2u+
kxyXoLR/d8OqYcGVZxlPV6cn/p0EJ5w9B4zzQdkgUI8ejeqQujPbqyuTE5yrHG0k
/ffEs9B3keA91WmFFNeutcXhksvPPfPDTBYX6Rgx51H/VMPBZin3EI5kmBCTUHgp
4ZrzbOIchBV0jrDA7J2FVcFETIbKTS63Ik8CWrBnuNEcRB7WHsUGfhn32N7NvUCq
tIofrYjHouC/nbiFVypFBKpbTX5Yy8aifhreL17lIu3t/Y+zh8ez4e3Ii2MOEzEx
OsWnafWAUoPiWlFULfj5Hnv/BsyISfHG9RWMfc7SuRNUWOyJxkI87osLQr3xel0G
BBZejfzCGIeevl6itxymy+jq0G1yugCtD50jxOpRYHK9gRbRjHUdJgiLUri0LjOD
7C3+G0lmmMGhBh8SBUW0DoW4BdUmJRUkEvegEE4M6UmlxNU5mxmNjy1ifQx92ypu
BNimM8ukHHLibTGJ49ilcVsqcGUhMf58j9JYYd62ErmOC8Ydl+WVs6xVcL3/0EUX
qbUiYZ7d90IYfS7ojXq2IsieRAaRJN0sdpMk8Y8QV5BTkkmAURETuqMZ+ebbGWiF
SWwfyZmIy0LsaldpZA6IHijs3VVZ8cuOEhG0MwtZ8ZFC8zMJ8yjflqR7CpMlI7qT
0P5ymjka3Jiv4xu8uZt1WKgMqti0QOqkfAsQfWhbBPOZrdpNap32AUddti84QeLN
Ecw04W5xgsAZyZOtgyx3FCaHPYJTXA3cHB25t5iITBZoRt3K35h8K3+J2NCHDyoR
XmXOx382MJYLtTWt/9pzDf3PauIfdb+CazrsDkhN6GfQ3UnFwI+N8QM+uKP+8A2D
LHrHC9m1D6cCLCxmVhnQdc7GNk6iUK72T3JgLdn1uzszECynxYiOtp7KN3hsnHdw
3kaDLQTGyiclAQhAtchoku2HPQcvcF2C6OVWsnxztjKESL6z/qLvkbDxejln745n
EZbBCG8dhtVNPDCq6cjOS6thSxfRgEz++oXINaP8QKViLwDdVWY+5BkTExF9rPkP
UrwiSmItOamf9K3rPXvH97wrd6XL4tRBsfeZHk/q5vIYdF+0LSysHhCxujBbihDl
7URbn2CxueEvliD6ZhMRWx9WTWG2dWHNZwJb2Ir7oBP/cSg/efZHkebjbWuTnFmg
c9uBpji6QSWG+6l/8ZkjTBMgCBYjOXZQz6Ux2SjXzNNCvM+dBLfanur1Yi5FqCCv
8Nrxw+a20Upj7mtue6Y47VuENBElx0SGRRSRAsxuGUEImFnakYJBj5wnSJD4nMo+
u5R+eX+xR2rDtrQJWuMv9tgETH8bk8vnyKSThV7whuOxB9+o/cGuV/qO9f9YgceQ
LA9wXGr2F0dIQE2oBaVqK6sa6qR0B8Lv5LiL+TZ7Fi4n6tMfqw8IHkvdb874lkVq
pbAgMGXXswNU2o8HjwTCUrn9rIM4y2EiDjW4+2K/f2Z/2xzEu6MBpdNRMb45Jd61
ccv0UG0rvPuQgDrGj4PUPlW+QK+Or2m2kNfrjmsePAZUrEFCzQeRRn7KBmA+EmA1
qAtgSU7o6VDwoZ07+v2PX7mQ3AgPxFgZrsLM4dbEEMU5fqhZCagT5hddLixhxV+Q
Z9VR2tp5IPUqM7+bb9VOkt1VQdv4EGm4fWSai3lNaDnP5EKaUwrULSCT4FK/CLlb
fV6Kakf7Ogu5sBcX4qIH3O4UY2DAFwl7GmI6Q25YwcBsA5/F+iBYspwjagLU7+mW
HbAiUuZNzi0fpHBzXYSbDL3hTzVuCxeUhdScd6wK8sMZ8WH4M2whXR9hHzkJY1O0
s/UUePnFzYW9JAdCj4MZRSqhc4dV/xqw7g/muZW4Q05GVq5ktl+hSzGH8yiJTBc3
CNUANugt1yECdBCfgirrFMxMpdQmAHlnJ1dG+TCmoF72UCHHIglnjqPp8ZQ2/BRX
UqWWJGYJO/V/rUsuIHb6pSbYQOXgNR5/0tBbnJhDwb/Cn/Y73H56BViOrVUJ9gsh
8ZUdlT4sVNfIkVbNhQQCDvjaXzF0xIZgJM3ghk4JVV589mK3LLIT/9y6k2GtXOT6
NFoTmmKsavW8zvmhq6UeUsSAoCGlaDfZgXHgvGvft1VjrehXlTcHKM59xHWaINSh
Oh9HvMCVHOfiHmFlh4gU3+g8P5JNHfMKe8Lbh3t3TFH7KYh1dOwA5M1gLg6Pcuq8
bItp9mWNKl3xIrVKB55jKtmUMNJvBwfFusMhZVLntMYog0SdZ5vLhCpmZudDa8pD
kR98+DaETUtsHnVzI1Q6/ivDfN0ZCghD2yI0Rk9cFHtxY9Gcy6RuYpyyo8Tsou01
jku6uxkjt8z2ysSe3tXWEa7caE2BPuX/mKR6RbwQpgiNTt3+YEgdeSH1Pj4mbj8r
PIfJSY+2rwx6Xt6YBXeIbrOirbnLLlfHWjdaq7IPavJGcIsqBhtB/T1uSCBXVNgh
zLNU7ufDXQLOLXvCz0GmWNWTDQNzaLHxj6qCQ9A9Cmt8Tp/1JBCLnuaa9ma7VVLr
ZpQdsbuSgAf+/FIiL67fklGd/AeOjFUk+0yJyw6Cr3yWwk/o+4DHn2GPU+UjL8oH
Q/jjgxwEfXSWscOYnoHKxXLdl8WEVNbzzR+m+g+aFwibgAuJe3LJXoU3wBPoki0+
LlDcilTnVruKYEUCROT50TN2iTzlPK7FIBM1GwxaCVvHFlJKm8AKrSWAkcOTo50I
DjV33ADBltvjmDzQPAI9GcgT2/TEF+Eegorg9FgKzVOOrl9UsUghGOIeYq4PsxRY
Lox0/6JN3tIN7USf17ZtaN+LritJyu4mgx5dU0/EiOyZtHjbxL/QpuybDzVagRdB
XRKEmp8imyWJn7v2kgQWe1EFa50yw+GBA48EDq7ip/WgiSZ1YZY7W8hTlU1fBNcC
fknTYhhs66a3VAJpX1b3P/90mHjSQOqm6E4/atm8BTEaZoqhjYcCBSZ3VqFMUhT7
oOO7onSeH8oXzroHGnse2m2H/dpC32NFMbEg2kGdESsxmNQXE615h97deTlEBZgE
67KuGuHQZj0m2F2/HhX+ud7fYhnkP+KyDFIbHUsrpMQ0WFgznwQgJocIUxKryLy9
6GgWYc4cNmK8d5q03rfBW/jev7Nz1n7ilrf1MZPATVcOu3+V+CdzVjUooOPPIlON
Hpf/9ZuW2XI6uWeqxLDMMNwf7KFEmO4ETbzB4dtSvqKBPk0CJgdrnrwclrUtO24N
5KAaozZEdbT9KHNx0uJMtcwXtcGKmE+JizDplq6XDZFSaMhByCP8AY0xiex4PRYw
3lodvIVjuD1PlPPwfjzmzMHWC5KLj3jlKJh2To5o4rWDGHB7uoH3+jXaO8J/8OMH
hhl9EY328E3NTFCX+/kKRjoQrxclKamagE86xkh5RMmWlFxWrdui0iy8MLCZsXgq
iZaONOh8L4ioJiCl13F8vLi1xb24S1Hlwr2W58pI0PRYlk9+K9axqlVLDhWTH1xe
Ltg3hG6M58IdvBPa5e9k0ij03zRC7vp9BBfIk7BT4WmRjiz4IMCbaF06Pw//pmsj
MFp6P0doG/5bjGKU6uX0HNZn1aoNiYq6uBoyFAg6JK4HVbvt+MVieZFaXbLQbq21
/A0IKH6MswzMe9xCMTXhJ+nVvzPLieWq6N5xPjKYdhwyvWjCMNhmnZZHsUd+yiY8
hXZazCO0oGv/+vzSC3wUIDb9sV8JLN683y2kPQsKHffeVmCsYZu+PqllXxsR4Wzv
zALjnn3ntMA+I2t/i4a5MKkIrVp2T/o7X7hLzJqISvIwzbvwyvTd23ua6Luymx8O
lml/Il6bZJMsIYSOr77Vn4Fj2U513xN3FP9Sg9VWpgJHXQuIed+xH2SdQPWPnRDR
t+pfd5yNZbNXalyko85oz61aQlVpCvyZQwbsyiC446FuaeAtI47mkrrkz8omLMV4
4HBhG7Mm8LqFJsZTbdmplRrXcljEC4BdTAxEScU/dN7PQ1rNod6liqDUW4JlZxfC
AEf1bY3cp7F//SeDs7WkSpux6XLut3g3flbTDd/PiUVSo/hB+wVKiRi8osVOoGXJ
xjGTntRFuDLMS2ZjE5ji98NHLKrOL7/IzKVuHKzGgG06iXHeWdc5amrsF9JRDYMe
TKpSYRz2xe9p/r25k7KAKJ4vokaM872vHxlIas8OB11ZLOAcaYaCUNpPbKXKYjrJ
8jO9cKYJ8HAmbbsJFxDYES84U1ImBBl7XHjoxSRzxWJOf2Rg2m9kqSl1zw10O4qx
bnzaxDhzLrVUQ8nbdTpcEm6tfmX4CfDMpwJr31BZ+HH3FpOV3oQQzUTytppl92TK
3H+IbY7VkCA/S8IlIs9NxB3kofYo8RX3A0YLegehdNQgFM++/LVkTcMOp3T+fM3d
YircndauYejYo5Qqz6rRvAOdJc4C4wzuPEHGtApMsqWd0SQxEgYkW6I62JR+zjD3
eo27wtS5jIw+9+80wzyqmJCJSPsmNT/YGXpXjhz/39KAY45oh/QZYKoJmxaYv8m/
Q7TdLqz8gWNQpyA/8CeBU90nT8vCznLwH6rNOaYpVg9e1xj3VoimUQJGdr0g5JB5
GGpdONc7ARaZ6Pm3g0487nGu78bLLNTnRPvX8i2bYbAxtgRKxZC4TslLyRCrTvv/
yeUAKTkk+mAD51rKSlX0xZlaPAuulJ5PnGBBUgHJSliwtc4wcCsRCVAQ5bTl9RI8
iWHFyUZ0lOhkssC416BBQvI43+YBd+Qiq67g/MGgognHvOIPNE3VIoUS+tyOnwHu
C2mZ9xS9iwfaZ7F3aev235l3N9zo0oUTkrdq1r9KEo2J2p/Rzbfp+dgtgn2kMhcA
iMKG62YKyEo+ZoybBBtN8hafU59I048i32cpCxp4jPR7cvTt0XZeX2amdU2Ijg99
hGE2tfu4fOpUxLWCYiyXRgT4feLkqlhnblPhkY4rET/USq2ERzrb68Yg9Dv9eo+A
VAgPRr1yLoP07my58Y8jUpRSb39N2sXuM6+Zqps2o1W1zXIM3OVrwdygjbanwxtB
/KPiEL2Jn1a76eVQIrQHIvlemLLT3RMqdG2+KF2M4YF1Afyp4fndLXbUYidzQ4Qi
OFft0nKsO7a0kELEW4dYwCGMXIAdfnzNv8/W6obiWYOLOcKNe6SOQp4hENOwAiJu
HxhaL7ddF5KnfG2fXinvyDcqV76XR1m5sD7D/orQRV2lnJR62qVOmtGhiT88E5TE
053UBxGPfq9nf+CGMU3gmZ//hJFh3eLLET/zVlYAv7m2kMNzCjvYTIG1bNfpeOcX
xD6lBjbn/vLqcHa23he3fENOlcMdxdUKYheXn9lS1izIiV34wH8JW6qar64l6CE2
lOSqcnEzA9sqbxBa6Qf6CJ2gmlaDmG1XsOjMwePSX9ktNqrs5bonlBKIMVDtLje3
5oaqpXAALScJDKbAv56zSTGQY1PuQaKS3+gvxr7vU/6NRSAU4ztwIJdQe1FQ1Z5x
D54tpNxRMhCrbkwbdl61b9rFegQBhJC93tnlDELM578JXuEFaGZ2JvPAy7EXhn8P
GQszx7JITrLMHzretpltnZ9fwQ607oKjiS5z0nCVkKD+sDyvCj+NgrFliuPn2iwt
QU9yWCcIeR+pS/OUrfp+EWvse2yclSCuYexEN7Dc9+WBxYPPiep+BRHzzz+lq2gk
qKq0hLWvBvyzSEn7wR9ocn8Lwt5KSuUyAMsQW/IPPi2AJ1eoBa7UzIQ9Q4RTjq1o
DeHkE+WhiJvwsU0A34FdqUt5M9KwjgR6Gp27P0RCA1MU+W46r3M+1gaVGldVe2XC
YSFkQySUkRKkhMGcodxvWcLuI1ifDEObl57bG5RTjY2b+DxKZD8qjF/PAubgtXfc
xKhuNXGTBTYaeE7/qFuOjoUnOsxNqGRaf0QF8WPnC4r37HiwyJirxKezB+gAqIma
1oCX+oi5bHulv0EahPmlBnthM+H46/m4wvboZAO7SwmK9S9ZmmUbAgdGDC+E1uy4
0pH/j2CyZc8t6lTLpxaCxL673UnowBYoj8LEJPcnkNJ9G8zS04AOYUDjX5tIzvZm
JMm0JTO4rN9+n820PXG0ALRBh3XCrwiG6IOvRe2EY/XMLGwNDbMp4dYxr++sPi4k
CH+BIRxvE5TV2Sk+RsoMthxeg5sd4nV1az5g3udqY0AMQJJRD9K8AEs4y6KpjC+M
tT81j8VlLACgoBkPXnv8IanQLiV1eBQ33SOQ6gHF3ydflVVBWbe69I8fyY+iC8ok
Q4yh4VZeondE4B1hJHD8XwFrpzNsUOGlgdl7JejyE4CjEZTJbEz4lL/0ydfri+PP
isRXeGmanENPlidCHq3pHqPBjetPKcdnNZCxbZc7wKgOFeb1ROFTKiooHBOKdGIm
re0ZK2LN48oXpxxeBvxbRRQk+/f+UGPmd3PCIL8nv+NQQgUzfYcTWlYBA2vhDDX6
hnnTu1o5ETfqZQZuQx45hNNZdhUbyR+1pVn/Uozf+Z305kSzSmfCqBFU2CbZ3Cua
aHqY6yUpb9vlWrxONyugvnSVwf2lsy91AYDMmLixgnDKnOrgv5G99sOxwNrJsA5r
dkDfAWb31MbDszPCHfvPhJpAd9TqPJBgiC0G5e7AXpWFkUkkz4Wcv2/rHDm80hgt
DusWnZaidfXpt6k0i1SIkAJiylqVm/KZoq2mgy2//xhdnCp8tSuRvgnCSmj1wESH
iqENU1jgQwFYEJev2o8bxuH1Zv6k5toLuO4r9f0D4eOSN1lOjmkL+z8ia962q4py
U2xFSu19UPMJSCnAzigyqMPGYV9Vb7g3fTCUw/whjI7eKGBro50pFMzCUPtH7KPt
9VriwfDWdDtbppt08h28DWKpYN1cGRDUccDoQ51VlBIZp5q/kmEdfxldHQOQwsuH
/2VyMYmCKO8OcI8aK3tSjDUXu2x14Ej9/lyCuCoih29R3t8STp5tsQyTI46tNOrT
ydaqHpuJ96ugvv2p6n5Swg7hPcoGMXxMKsEJFiFq5gQgdhG4Ti/d8t21yjkdaLi0
wMPG5Wv2zJnKX+Pw56CvEzALrxhfUFaLAB1gDmRvkcJiaA6mi/XjPXSe7zGMr1Fw
ljthgg7ezV1xD1T/laDPidx6+1dgwF5nBdzhZC/FtT5PhKbAnlzZwdi188gs4SeI
+hVhCd5hZNrIpCd2CZ9fACc+Cowtp/50JTw/GbD9Zj/PiglLGCMw1r5PJ5ppC31r
v8vvsOw4QFkjsp5ZgM0yKZGma1rHIsisWShBFcSJhr+myANY5kkiiGZQDudWRcfM
Xv0R8SWjnl6+b9oMnzoU7rSN5qM7RbBxMQQuvUvOUn9m7bJq81tt64c+egkWpnbY
vJEHeK8ga4d9najuiYE4NDapXRqMkwPk1HUmjDXCT49Py5mjvLytXY2apuQCtZSS
L+ixFEJNnOPPX1W4sxVGWSa8dJAiUDoFZc2S1cAZrAjru/iAjH7RXzzhOjXwGwsq
md6dOTRQf+Rn+6IQbOLuCC+VW2GdaoFlqshM3U0k9sDn5dR3T2Ihf/GYkA8GW95r
+zej0ua8A7eMe9Jx1Q+sP9Hb44ranoh8ulcafVzHNeSb768tRRauiUWhi9xgwbaV
3wOugmPgJxbj1CZoFjm037PFtiJFGH1HsiXSuBoJ4GMGBAa82jdbZ6ocPI5rHrXX
iBGP6phHbPogL8gmzfeYTTPLGsd8I6yxq8PyEybY9/odv0lA25/ZShP1E9ypuycu
jyu3XgPJ/f5L2V6wWkymIS1sONtBXIDm+KXCBOO7ML59N5RJAlU0SRAYsLhAMZHK
QOu3brrVLwBsAWPQK6N4zJzGS3E09pih64z5egXMMGKfcB32pfoh0tmVj1vp4x+w
JaGGVy9TzaHS5wyyNMH5yytPzc6yNjb5u4pY/QGFSNdd1bDs1K9iT5zRYyy4oqD3
e3XUpMnKHu9UDHV00hC3deXcVQIwYy8+tSsLV5r5d3caeF+wBovq6RX7HBPvF5vT
TnOwe4CUfit8vEqynNsTm1KjU3na2FO0xABBWbuZGXF4Z4ULJZ8ZElpXj1w8jvUe
yTbJ8OVTKBEUQtQj6kSGMO5DxP8orlfnz10JSmAtjIJH8XJZdIEiwRJQWjWmxehk
em0L6OzA+ZZdFmzTh6GLksEhZDiMb5RT0NgNl8Dm65XYAzXsk8cJ/CrgOta1wruM
6YhikoZiDVwviWDSmdI1u3dXN95Dka7tDH4bHhKaiHtUx33Q0fncmY2YyAdu4ouy
5Nq0/rsOW03qs1mbU8Mc3wuAjnxCl9nWqoahBsetrNFNp2cRfbrH1HFhfGoFg36h
SKATH3Xavw0feToFG6XCfIoOj1FqB7ueUBx6d7CpCtWluvwz0BoJNVPhyGrbzDkl
4F6oU5s8rFsE95Z5oARqa0CxBinqR9IJK5v0FpCysRcTwM+pwHM8GWWr5TfDLcto
k+rlF2r5/4rojye/cdowmxaNtTmbeeMyvKm8+eWBFOAE2+4eQ1W6sEg9jkIKd1ju
tn/LAIvxU3sHqQRLK+PomriRORQ+9x6vRFtjvrKGFUu2wyapFROc+6jBB9vPz2Os
lFbQs2qx2wEBKYsEIjpzMocYxmFZ/V32sGznyV8SHpybyLc/sKRLUNOGY2UafQo0
O4is2Rp0dJ9JVBzoyys0SRLDHrljxip4Hzj9U/gIRAY7bezP7l+cJgufTJ5RTD4a
tuygN+VckjR22kNDiU5KtSnyih3vvIj74gMyxMTw9wOw2oP1JQGGMfbkNtmb4LBW
e1Dl4IlKms4UMCWFjKtpAHd+Nk7P0GnSkAmMdy6gHcY6ize+F7FS5wWCyrSsEnSZ
fHZs4mkj2wwgNgdWTQn6aJYNSfiw9F2LWu5VltZPyeNKaGj4EsYCJKzUDuVKO9aZ
wrCr8gAMEVP8DPc39SrkthrNkxblTwpPVgu3Js4OtnLuOJ2dBwIyzuaxSkgV7lvx
MAUiylFy7HJrV6gYJXfMMe9NvWDHBPMkeM1YBEzMx4Wka33z0uPmqf6ExC4BAPEt
OX3SHJS/otUkuRJEMPMvwe9bEEcG1MjBiEbvpHO9HYZrkPZFXhR/W4fvJWIqjo8b
ZxhWPeXJiKsuVicnMd00fs8oDtlL00NC1CMk2VdJhrWqGsaud2xuqAy95v1oi0Be
GbJcUtKV2KiDvhAGMhwOMrFYCszjbw6o5X1/hMSuCu9G+Ysu1OSUYodf3Vn2XNMx
uyx/czadoX2+VuqBNXiPSqtyq/UsYx64qJOJSlp1CZHB+HvBotd+X/UDdA4pkePv
5FOHiKbmQuaBGHiTe3VmcfE6ipsiM8wzDAvkaZKwUe7x49+N2mRZqUureKsYB7CX
MNBjuFsOoUFyY0TMSJ1+p0wjt2r2snKj169ep0FFSGNnUlrH+0MLIwGqzVEk825S
H66FR5VDHH4GQuSqYG0WximsWRq+3kncbAE7lA/mcrGdVmqv+RKoO+uemzzibrmx
nAv2dQ+2shfjgQgUbCUBUJND5ji163gD9Hq4plM5h+4lAgo7Fm8e0Q/Y+mOYhsa/
4XqrboXCiNJiiEyYvYKLf4Zw/oa1uXdpPE17PyAtsmGyJyVCR3CxyYu5DEWDEmIN
MMPNjRW4UO2JxT9bmoxJcPmEeh4MlHPr2XU7m6hfBaQSHmJ17WSbDUSYv87ji4Ot
E7Q4cKN9HgZN+scolLA9+8H2WRpWDqNILziYZSD1dooldg9Ct2WPrkrHKd1yz4Un
tTVF3KvgLj1Qjz0eXPnzeCLbJCKcVtg9rH2kdzhwkKqIZ10xnGNogCwJDhT4eHhH
4v9pJNKdS/OgfZE/y1AuUCYxJD2p35daD0hyfs4fM8JY1791WH9gm9qmrtvtfvEc
b0jxejBCilLQqzIZ77IU9k9kgQBsuTycpcED0DT5MuVAInM5jmxgiVRt3keITRKc
iP93G3DvffwILEDdThm8r9yz203x6uDc4XI1wTpBv7E/45w0JcgmiubIhdwsPmjO
hCtwL7h+DPOWXsOFTkZK7lsdyn+7qG52krrXGdx/dLmdb2mT/pNJS4HTQMw0qKWx
3zoEuR/9jXEmJVwwa6Z55rMSShxRHB/Q2DnG56eDH2X+EoWreTuoLn3zxg4v0yN2
+7os4F113dikK06lu0fh8XUFIj1jt4twdfWo1dcvkHlphMTc4GH3EZEqNvVKhgPK
bfcVNL/gSDhUbBcjnR51BrlF2cKh5S0qwOaHXTy5hh4KtehEB0lt8K/bTIvrCMM3
fcqWrrdsy7DHoQfS+8aWfFbJSTA/XbiOFgc91U6Vp+Ca5gHm0psGGnOnjL+sMHic
p5QuR4cDFLCrnm+1qXXHxE87QmjSIqJeHOJSb7PjEixPa0bvZCXb9ZHvERsHHiMD
hlHhrx5NAQQ6I0yJSnx7YqHarsWFhw95lQLV7gRoIsyj5GkjeZrbTqVh1t441/iL
CyAg9IjRZu/siS8js4yUja+BLOxYkT+faBLAnJ9ga8prQZMM5Vr1cqG4NR68ismU
FC3bPW1JE3Ck1zfFJJASUFcqPc5h36Rnp40zhc6BAn/F7KjnYog+Iu0VvGnTkrTm
uHg2uO96/wWe55p4XMETS6s9DObBPF8bk/O48mYBVdnaFo/P2OMvqEsAY+ibveBh
71Lsy+gRQbaKSBdhDPE7C1WqGmHVd59TVrwSnEWkeyem9HbEjqyoCpprCwZCAACI
Ysv4N/yLKxSgEVmcCLf/GpO3GdXq2ZcLm5DxsfojMRY0GyxtejCXRWFHP3P7vAUh
EKo6OWNQgWVj7lQAikcENYNPJHwzox4f2N/mLfiANGWI2KV2IQFiAGMJzKyfYz+G
/85d0vBw25xIUdpKH3iumtscbkfNTtaOTRjgBYKGQY6Xubs/ElvqCEA5n0Fl17Wc
o69ndMnYbEyVD5ivGl1xGgetjvoxhPqbpvLlIje6NIVi6ShycNBG8DI/EuYNtkc5
Vl511yjRwcGMd2PgeEoKKhqndw4HcAe9cOF62ilW5jhrQ+j9IbOj9z4XIC3mo0j2
hMdwfZT4y5pU7wAYp9cfBrY1daN0nbWPxfZTRccLU8kwg1/l0L8p2tBQ/uyD8hX+
WpIa91WYaX04uCT/2NNu025t2c9dHcZFQqI5y0okTlBi1DPNUSidcfC54FOWFnxS
myPyKt+u3MZz5RBkdJKDIjSZCOW58h1riDe10BgzTWicIgsp3hlYWnvcqvQUWfNt
2ykYGppaRJhwKbaIO8WHO41iKWPG++Z7Bb6zmqr6QTgDs9vaJyeBAXQ4Rf9wPekh
SMNIKcm7bsZJgP4IJMTYb1LoHY5Wvzd0XeVCNCTy0zalH77kuIeKaWznucsoWJVj
PEE1J3n8ZVq6LFJ6VljH7d6Sx1M9CCcIDX0lQb3zclLiF0lIhnpIKItMceqwEebj
2IQxmJWnTB1J956IkjqSt7ANxXCm2dCCUjx0u5G8yOmTUNVrL25fHy7yrO2rAeKo
M4ZlPgKOZlwIyzhfklWZYh8JEUVOQcvlItGyutG06suIforF3IOo3QNvGe7LNqsQ
wKPfAfdtAJ5oquVWJ17PmriX4HKxJ/LLVWILA2NqvckC9o/6eIGciT0EDvHx90Rj
xcdonymLVIQ5gLcnv6W+ZM7xipzdv6bSIHlhymOIyu4+HnnjmV6JHxZz+m85xqvx
8WuVAcdxfVwoaAg3szfTonS5rs2WTnmbkNJoLTTcxFXsuZdas+/VozC1PapOZNJq
NFQmL+Z5OchlsMPQRohVaR2O87SNo38eUIBLZYfsl4JlBRRdc5oH1iGV4YOZZvij
YemE+nLSVdOF/m9Mxy6Zzy2dP0UDjwgqIqOv63mYhzOrOjESrBHqLmOM7qWM6wUp
QINNa6nFHh+dxoNnCbEhKKtln+WoQtiJCJxaFnoc1XG3ybNnViiiPDtHY13xGTXL
lAqft1A+ojP+n73mgiacmkjPPpUvRabAEv1F312TTvzrq1sH7iceEg7VgLGGhsGT
SifkR4lIt2RTHGM4GEQCoU2jZr41D5cgD5rbrS5AbCDPRLBIB0ioN0VD314HzSI8
bppXRlBcmtbiN/tl2kPEAjtHJTDXPAukt1MWsf2ySY9dGeywGAf9Nit/xFgOb7PT
6OamMQav+awPIkSSW33jshrItcNqMEw5bcS3tzQpuN5sBRa5tVaCvPkJwpxE6B8Y
TiI9wMgUVs47RFgeiE5KpKw8+BPDsknBBAGc6UpXUtUNdf46c7KuHT/Fkdjg0/4B
bIS7iWlTj26Z9YOJweZpslNms85uONyRD9jNhlTNRQI1RlnnG4XNgJUiLhutG3OI
h+4Sum9v1S/YA6tR6aSk7L6poUhir/btlqT5678bmW8Wyj32p4KU2kLPH9LKCbvE
XXKB37h8F/rx7/YRQSE0RkhdQDxM8ORD9rWfUANtbt5WC8XM6OWK395haKScoQIs
gUVI4rh2F1ScFyoVb8WXUxQQ/B95l1mQ9Rc/FYy1cYuh4w9C+JyxiLToPSnP9/Dt
zt9B6Aq0B4r4bh/hLveeZEzDh4XVGJPW5xSXvToktdzMLozdyf+u1uAykT/zzM1e
qoQKsh7LBZxSticip3ENoZurWMtYms+c0xEufkBmb3M+o3AYhWW8NH2gP3Ffbzkm
Ba9uX7VkmHPth5SxY69p4XFbrE8mCNH3clTxCeDxTBOgLm49BBgNFhUI44Tyl0n2
QRuJqn38z/3Q7WLMog/t8Y/TKsOB+RpM7uB7KYJTpImZ36XniFvVIZ/VzbatjKQl
GJxZC/cSObOobaEnZSOIKuNbJ8IcxGmv2u3FDO4HmKFXQBYiMvPeGfH6oqL4Cy52
JIa9wlRlpuc5tVE9PEzrkO2lLBhZERF5sxwNIpL820KoFfxVL5PAxDl138DJdrpP
FesJHOtfe8flPFwlX39vGZgKtK9cLWM7T3nYtut1oviOIzYbfT/5YUJgO1ZJlkr/
UpFVsk9TqZyyDShRa4ZLbrazluyZJY77NGFhSFVDvGa2lJP8y1uw7qWoCNrCwR5N
89A20uDVPUSupXiK4GmZVaBpeE+jsaXb6KxPwe2FL2e4Bvb4TP/gjXHXz+F/VBzb
alkm9s+dxA/t45K+/g0eLsk4tPBWSH5h8hLnJKDeZ9PK3qvvMwePuLUMio4RSex/
lFvdUPIHJlUbaoAJYbHXKtBzDv38L79uq8JcoWdSEMV/rGyklHEpqHvYd6yCGdPU
e7rMJwLlkAsA2csoQ5hJATBLQ2+vsPJif8hbh/dXhtiYAxJsLABqXZAVrkkhSuR3
KMuFrf9IAzuXo5lBM9yQUtYITJf65ojIenwgDPOlF8W0u96dO7fvc/UO2MzUlByC
nmMmaq21NkJ1dQ6EjPZVl3SDY+h6TMlDt3OvuIIzEvpT6x7RJTjPVrrpiTMzsdFm
KelvwCBZ0NK11oBqxadASGiug0+StgJphPs3PzxFjLE+DW2Q+KIqj0xR8liH0U17
80jRRtrMzys6tJYo9mPlCrBzGc0eNdSqID2p6yfujPXO2UBuGLal2ca3gETMOJGh
MDRyprVLFdClP/1METOssuVDj5TG46LUJryyN3Yo9AShcBQFa2uvH1S4zAR8Hq9t
FZ0psMe6LlgnpmLxAc/x6dYqYorIm69xSmMotYoQ2w1ATStk0KNa8GA2jWYV1Sr+
xyqJRX5/kcADKSk6tmTfmYTbuBOqJV3YSh7b1lpQh9s7Vk9EsiqhiUZ1lljwXY1Q
GCCbZSfkBZ+SM5rSe0saJIjRVBzRj3HsBE1rATfjM7RO/u06WhbZDhR/SiauaAiI
YGCALVseZKdJ1tW2aJ95d05JJOlkS/Yz2jp+ghlDSkWm1K7vGUTBI6c5ZiGfVpCN
ONUbhLkJgxB8KmDfQGgxQ0O4VYLJ2xn0wPeTFXTSRlwg0dNd/PJoMgHe5le/Rwbs
OTjsS5nWmMIi0eya+M4YkbmN+1IiB3hiX8TLzFJxKJVx1/fiwEcrwoiiV93yDfwd
n0ZRJFcSCGeCSmWmcGirhxquISomfMaOf0aGWQDb8O51eqyeNJaZgjTirndEcOVk
yUA/KIOFAouuRG9o6LLjCHGYuhHC/VXysdd5BaPu6ENOYA666E4XlIDPdDOnXCCp
7cT+E1b6ZnxiOZ368Px0TZCwPs8T0pjroy3BW8I6cY0FgyNcNdcLWbv6xjZ4nv+t
EJeK1RjyHSMrQgU7Q2WRBpLl+Od51o7WO9F2l0NxYz+/lEcch1E7wqKcOXL2TfC+
gsP41i3dgAGhVPe9jkRSmJVZelhBuUjnzix8FfKDnOfSCAwURSJkEqU3PwGV31mo
vTeP0eny9JylsUfmrpQNB1pI6iC+L+VGb36xGPceaeMHdIAGnNf32ofMGzw6jnco
a1U30uzmd2HNexeXl123/PDUV0iW3f+VgeCErvEzVo7GknDSSxlUkSWreEgPerdy
qT6uVMhpLDQc+04T7qqKyHhqptratGjGA/lAeMEjX1qmuWj65uieKk4Ojyc6cC3e
uA3c/g8J0KNk8NRm7L7Wa2MKXVWu2fep+GKkC24075Mh4EEHYk6uwdgyRZr1TaN6
8mdUYTVA1C4XQr/dr8A1Wr69jOqQXc4wLLm7MtIs2r1p5zweKfAAalTky5rFtS9x
2r5VUIQeCggZ+oV+LjtIKIImg7hBUDAvv9er8C1T6fHkVweJ6ax4UEfz/VqJG7oQ
PQgqYviHMbleE/XBBE6pwpcZk+zKrq/zlShQf0wGCLQXHdL6MxV/gHHDcRs42BuN
Z6wFaYQVYwfZpjySlgRVfME8uxRdJyJ3KJ7AXrZxskiDbEkOa6N4uL4R9JOVUH3y
12OOeoVEDu5DvPlvJ2nLagMYajTqBpAr5q4RTXKL9Yy1OUEfWH14x+XGA6SX6tz+
XuZNDgPrcUDNW4nUtoCfj+APvCPhf8X9EygNXKvNplKOJcTuRxmvB3+jg2qJUAw8
9nhL2yb6NkC4UtYRdwkqnpn/3xrNpfWKrRpc38Z0D7Z+sAhoFutESsvQfllt4xpz
y9MfyyxfikMxgOoFwWur+/nDHu0jzzeFtr8oNASGSUQIm60OF+VKEuvGSma7Jv2U
BQ4denno4alhLJUlKhFrqQq4SLbOaZl1vgNfJL53yO+17MiRpKcIaVwbhcBS4wAj
BAf1lfXWNLCew5MrMpS9NlzRGEtAgtFQ6zcJ9AoyCCLcjgc4LVaM93C0i4qWi0Xw
j9qt0pZH+4ZirrH5nRB5lJZMNKHqrNdV+Kcf+/YHmyvEWKB+o3l9zyIJSR+ITeHN
/48rdk51ZXUibIZaBttA/VReczC6r8NZJco8tFJZb3l0Z4JwN8lWmDmrroKkVOJ8
zyM9fG3Z2fIAoUOlGikRv8AOGCOxGswoPwONWxhL9t5U1YBteXYeLzErePyOZFX3
TqUx8Mb0aZOiLqDdzxjUVzNUCrDF4lIrU7HXHV5lGBtECH9UX6Uy3Ohaxjob3p90
ATasRR+B3VAAUIH9q3bzm0AA0FRXtjSWl4GlFlPPCtJU8eHJHKuP8kaon/k+Ze3U
WJ7DYoN5jpuq792VQcPjVcG/aoaPJnqC1gUK2daRbHr3h8cuIJZuzGbU4uFunAEM
mlN06Ho7tjT/1XeWmgckuANj3q816Djn8jiXR40218pfKYQHSbHQO2HmRoziNwfA
EIBvyQUw/cRUxTaLkGJ4FGT6wHnRW5WT0TL+7oPO9w6LcTCL26LsiKldEzRzz9U5
uKrcVX2yksLt07jIzh8S5ef6dhiwTVMwvGZUEhmve7Xwcmd5pZ6YaPkI0YzYLHiM
no1+3c7JlfRndXRNAGiNSBslhSXLg9q7+qnKzsH12Na0khInI37p2oOge7qeMcD2
XzhiufUxYRn/4v59qa/nKeFgAQ1yRBflDFP0wbhSjbpPOTglNNw94udq+KKf8xlM
pDJNUZn4pmf7c3r2tzMCoqDsp8/vE+GMXmslvcULEjk26HgiyROalfy02phxYk71
GL7YPkTE3m9o8yf232winnLzor/1kN8rsWUSu2uC7Gy48nJkPStkJVYMK1mamBAx
RlLn/nH67D8TSGpFxi/v/GuBFQ06kg+wAR7wM8WfC85Bgz/bOlLXUVOw0CyNLoJT
Ds+VCboR0enIF6KF8RNQTf6zB5Z9Z1tYobWnoCU9nKrCx26Es+/iF9WSmegcAW7v
fOfTGL8i+WmxM6z6X6kKGoJ4AWquGzCSZVM7bTzOdmaBk3c2co28X9lGTebM8ryM
1oObKRVgZ01tVKSg6dMvjAJAh3U6JYw3HKJ0hxshtOwIw08TWnNSCGPP0y2eebvW
/9AfkVnn0H5WOaheLu0uhn7wngM+4i2C2Ak0jTXwwy+RDwMLE9eQu1GOu5nH4XWv
7CzZjNQeFS5kZAVvHr7hPHTUTVvR/As58zrGITJPxLGTI0uXzYOzA936tWxTTvKa
AUXQSnsVvleDFkrqAjV1bERWpDGZUBNbu7UoLiLxcnkjhMIGF6rsMy6RnSC2RdjF
oVFMQPq1BdMZ3qORsURfI6B0q3CDb0bM4Qbkp2HBWDvETU+sW/o3BlK7ctYQT43V
mu2J1D8jYlT0bUKEl1yewTQwJ28C6gdA7wlZ5i9GQ1Re6crkHfMGznSgyIehkd1H
L72KW9cXzAV8PmPHAx/HG3enXCa4n+9vGAuQFaykVAGTv6GgqxCBL6rq+/x5czkd
FXkwdrCz9pDXVPTQVKppNt/VDUx5HUd8peiQ2YR0ViyUFJzBQ0E2YX88fzcq0oUk
hwr5jstEndO3g8Om459vb64OxhDaSUdK+5tGKUPipulksPNk0lsvkIPS7bKXzybb
OREjKzt3OeRlRHo1hna/35Oj19CF4oikWwHpp/LveSqDYfgETNCXM2rZtpx7vVSg
T4rPTX3zCqOEr8HeXZRXR7qXliK9kl3ZHxmNV7jYpkoxqkGKp5w+N/DW/+jrPCUV
hqgyWhbCGTEbI2a6AWAZHuJGpLrwdk13oAI0zfpUm/JLOuoSTNE0+yVJHLnVzJZ9
T/Ts7qlV/m4fjlnZ5wlfzo413oaSYTd8c7qCdkq18UudCz9lUmVWfuyWD+lIGz/w
0/zzyyUJWZhc6vc8mbstsznAHVGQAwIKtQzKTj7Lop5aSm4cf/+VaF4nLkymxjbd
yjnNzhbDwNqAImtMacW6onkfMhyQjElodLJQrMD7Q4IFhoS73LRRT66EqLpizTHc
6vnYAOUIwoI7ZX13qxFnPH8PvgyI51P2I4DFEYz/5IkaMZxHqxchD+RlJxCTczHH
pvqCnEKoo7pKvY5qwqorBu+wiCMTmWXWtlU1yCYuUFhFMmt47lFzM+Mqec0ZulCz
P//NBuMy3vTGOwIxN4KPqq4KzXRCKdb2pSktBcF20siUpkOW62mJJbcPd83Ox5xI
UWVtKLxOP7xBtMPkEbT7ASQUD5z6htWkNiMc4kRiCZvWTVB4DlqBU69igxhwop7b
16fVXH/poOufCg7O34v2uCfdA3QtUNCZ50day+r5MQ7SA5RqDvG8eOizuuRdvrvS
eCbbfWdCG2uxKVzrZ0lPqXeSwvneFYwbVgZ0PjN016wA4163Q7X3zj8rpBwVKqkm
HYL0MAwIDar1JrXp+Npv+NyxaEFer2zh0pkMJOZMCgnkD4p4wwhIZmm8mb+wl/59
w91UBBHPXYVStQ7C3mgePwKwOmARdwvJHbsnkHIQEtwHRj3OI46VvDzrT8UPUg8b
kdcZ2R/EWwHBZ1ubzwI7J/FZs9bt00ekgM6KWUON6K67zkoYZCc3vohzK6McQ7ke
5BItGbOAes/g4t7Mj5DU0KCBfMq0ZweJKDpxMnkZoX8iW9EMXVKpWJuqU5hdPzGW
8hyh4IliLzfv4CzjeXVbiA8XPl+tWlYMGoI7BczGUW1SvmVr+Ac4zHabZ+IvBed0
J+RCswyYsf1FAVY3Mkvdx36U9M10i0+0w2AhougiKhAcW48dyKCuxd5CSKJ9FKNM
HGF6Sdc2pTBbzZ0VXw4knvyO4hrB6dbQjoH1/8+ymHrOJclJAXxXH6jn+fU4QlFk
2tdzGBIJdgLMhGVyhUFxkxxctFzHpiIrpOACGvrdC3wUMHgyItZW1NA5B3s76L82
fBNN1F3oSeNdNv5Thi2DEiXHp/BsIndZCeFZP25km4bkfKs7CrWKGz9twWnvu6Jb
cRXB2WBZz6pqVa5pX57nrVXi3mt682NBOJ/6LlbmO1QmdzVRDm4m+pBOcpjVYvja
JTsm68PavpfAHZfXBe2CdfxZEwcSt22N3zQuRVMWGEsOSviQYLUsPnZklYt30JwJ
es40PfX6qF4CtEIFKqzuyQQ26E6o46JjQ9GY58I+SPdkwhzS4sdYRMDQWacpLjUo
UbGeeDmkvbAH9ZE+KjeMnVYwZdzt1jYjHHb0EXIvw0p1W6lLKDfKDDHLYiPbduix
697DfOPYFZkiP3wTafgQJoxRcn0U6eHkCsLKgnCQXaRWEc8odOqahIIsCU4lsOaC
2ORVZ4VtULWHBzin4zsTinSzFGrcsailVdWvTzfra/dD8c6k6JAtMSwSuepTooHQ
TCtIIXhhhuxp577Hxy15/1FNAy+PBigmP96OBGmZ7nR1QfnodK5ko4bAAdXwCDnF
o5ZuoZ1MHggZvZqZ6Ab3cXb2nvO7M8HWw1Ik9UZ7Mecs/DfQgJKdZTlchirMceNR
dIz7wtmbPyzybofDNFEaBEkxXwjpQcZ1mPcFSTFh39vXgviIooualP9l0gChb4Ux
HOm0Vl7zFac4fzhLISaoLUYQ3/Pq0Q0txGUD6SvF5UDogTIaBVbSBSwjGdiXECzx
PtzNolbgFtl25lNVw8u9EnMKBpWdFbvsEhL1xXCjIYeApPp2jn2wlOtnizwcqRfQ
kEnh5/fc++t6M5dHpduWWZdpkKK2A7w8FWkPZuUXOdtApPVPDGfJSRUCZLKjANNk
1qtitIfjYnSPokzyEOPT1n51nldiH0AH//tOvNcKRRCXI0Ru+i1X0qR+8YUkLGJF
j+5bP7G5mg8ms4ZAXgpfxyO2Rk6DmasIgQL5DOWkOXxWFJxW/tLkEPytzvVmCnAV
K5t8uNlbL4eeq55+981/vCYNhJ9ESmOEx63QP1UgW04GwROkfBdPUpgE/h5lg79K
wTR4Kd+3VvolxsED0swlB9DnewPnYw7nUNAnfbLXHft9wkA+fS5vm2xcWqm3p8yM
OE9u/EonnXzYf/FjD+A2hzX1ExG07y1Fgh21W2+NAPBknWm2BbbG6tEjCKQmIcxa
ieYqtFiQDRyyVx1p6pFZBBB+q0kodNNWNtF+0Q/HDFvmKKbAcfMTqbsoHJCI2zgz
i/rumH7XF6Et4WfAN1DHN64q58dFE+N+9CBLj6yuI63D2A/UqWoDHaSTjEhiwJd7
QXarPXTcVXHaaROFRGzLGvC3sAc5JLjaBZsqbFVg0yDEbt0RJMp8SpO7ROhhZseh
eK5L/UBNM5HlkFrMZreDVEPBejDTHhH4RMPdJ/g0XFfG92M7WHGbxDcx41GqoqTX
y9bAYMPCNCJshHQEDGiEJpywYYd5mxaG9umVPOt3G+qY2lnWlxT6WBxrwyvWTj7/
A1trtN4lvIQZcn/neAmGXy2KRxLabESayH8lVsi04Rdntbuwa+amUXaWxLQZKXkb
0bru/vf7Jx5HX17tObuxd/V+k3U7Q2Q2fpNgo2sqZu8BgnqZ2e0yN1ZBjTbGoOwv
0A6GEB0gnrEI1b2XKBrGyVrEErPrr5l7c9rHu8KTICrtUWNMYeJ1QBxOyXK1TKaY
VyGkXYMiWTKKJVcTpEthLBUJvfVH9lqq/Cs+ZEQvWKHloo88q6sAYWRQaiep1iBO
xrbhNGYiCdcjWM1NmKMM6OU5dRqV0JXQTNFDHBcNo1VPZegsUFu5tVNpCgMdIa4o
s2r3cq+gDoYIkgFXgAsMnH7cUqVfD6tpOGXvsxXFuzX8IkXJpuJWBIAc6I7nEMKq
DQPnG+aTyvpVwmBYx4r5zJ/IuvC8f3xbZa7juau3NOcwqw9pPILnoXMYydsAbk09
Uye5cvGUkF964+2WF1A2qeY9I/mTpRk3RlaPdEMfC4gRPgig0aJi6VceZwyGyDNt
i4Tpee3THNuA16lWjgw3eYDuez4FJUOP0M9I5xlZDxhBq0GMV4VUBn3aLBS6u6rb
WgAx/JOK/cA8vEaOoxjAW/4NdD7u9xnXMSgh7NWHWDGbz8rnOo8rQV6g3yyb5B0N
lZkWe89olu2SeeXrT9+cVXqdEnnuGJSXW/TJwZVryB6CS4FolBlHIsSB8n34z8w8
6a9KjTxcLiFZzuGu7/HH6fPUp7D0OBJeb8YUFGxKPJYw1KLM0jc/GJxGobSJj2eS
2OMk5PvHDO0hcTTH1a93gwj1jQQNNQNxtbnZ/dc9amc5uKy1CWEXCZ6xjxpODgMd
VrdfwdRR490NwwsbujqY5vpVqEqa1W0VaKjsFKmkp9dlhqmOaJKpCBm16Apb9TNt
39vu2zIc58qRGArKR9Z1DZ+iqkpuICB10vQo2mMp6n4jilGIq2PezKNN8+qVAUwC
0ZmJLtBcdRU0zymd3/21zcixmIEN62ub9B7MC1pQ1hBfXeWigfiTdzO7QM++cIvK
HRId8oMrPdVx8ich9upj7IruJgYwX57gNEHAbQbllRI8OzSCiVFKGCWKi8Ayejmk
gHo+9t2JEGBBU/lznxKKPgVC8ZXkCO5YnCvCcX1TzJPullec72snINY1calEbIYi
U6LRGWAMjBVnT7yTV6T/R1Bjv7fENG9QNF9IeH3CK20gHc8hzlf/zwmkN2mtsc8Y
40IddUVjAkRAGu1r/TAXrcGx1JHKZalGQVz0oJYyVu2opHccUH/NToRKGf1GnjDl
KTZkE2+1kB/NIdz3HT9ShhLA06VjpEmH7aVGW+nVasY5V7V0V5wb6KNs61C5SD9R
mZ/cEwRPWZbdJ2A9+McNYKvDHV/uhk7RIJZ+/H+GOLV1fBXRu+4WlnfTsgcC89R1
SwWfLtlAg7IwDrwnGoRI+31Y1MresP74XyvGgFet3vNpvgw71VAlw1rTMgSr/V/w
T4A6Ko44CJ7PJm2eK3odbll5RcR0ZuzHATIfpahbONLOABwN/xPJCOEj7zuEif1g
NIT8JNV2oMVbg9LILRcJwheVNmoQHX/oaZo0xh27oF2UErC57YTyvcAxOq48NUo1
pEcc11CW3PY2ysz96t4uJEf3D6Cw9fLtacNIo14HBOkxFZ+VQgNeRPdLREJWQ3dj
LFmgf3gYC7vsa30LiJqPI3X1AVlttLDMIhmLif1IPz5pq/punNF2A1H9feabJ6CR
1830FQezMY7ukw263mLWi1NYCBMA0BQ1k3raoS7mwO+d93RtxEKi+255E4Oo4lgd
AwYmb6OexdOtcmVvtwbWUiBLZlgT3fiD0Spns+RGtJAoDW3A9ddHRlt93tOfhDHP
cznzXE6oTSEVtMCohpo7IG5m9hBBzY1sS6H6/qow2kaszIx9wT8N74NzWmZtOcfm
oG0M7OVXV8jGcTYmmoINBGHHA7oGfymwMJCQdfvKJjkHkeUamdJvyhuUPu/MOrP8
qWIUrKwWG2pX7TZWfIDofeuh9m0SvbSQmwmBROKLq+goptcWR5GfQ40WvaxsQia2
mtZl9+rtsMAu2B+0do1iRJfyzG01W4ub3lw1UJIo5842Wpf5JfpwF1VlmllEfhy5
CtfdJunwR7+s0yau0nc0Xxz+Nn84N9RLxW8T+nPM9kEqib3DMDfqNuuL2yi/v3x+
dIq6j8XGs/ok4a329X69Bf9E645h5yizSOqCZwJyOrBRO9VdiE3RP07MtLGdb4Mv
ms/M52vJjitOg6gTT2Z+GNK9oqlyDU7VkqFz2WOl7VlxLfHnVKTBAYwju0ItjHNy
fBUDW4r07MnsnhWVTqV9expURKQ376CAGemNCcT6ZOfV6lj0CMKBAIISSAiWIacB
wxt2mJ+YHDfQqi93zwnMj4gslNn4wpOyX3nB0IdyM8kkmWEw8SbCD2+14s7Kmc5z
tPgbYlXKrdpV+acIpiz8cQtXfwJJErFVSOxyxljmSSBQtSO8+F4NwHNjW3RXGGnc
WT+QkJ2J5qQWHHt8zmPciUILhrLBSGh6IrDpzLz8YJGoduSkDxNqPuKGN9rF2T9U
eV0kwdncT51eCYB03c+4FQ6TlN58pef9YzhhjdWi002ptaQVB6YQNHUqiPw9JWWF
lPgeCsYIP6F/sGvm1k4VyFsRhAiw5ohwYhQgXuenLLxBffKTFzAVmC+LUNTR8hu4
TJz+6EnQIu/6t1A5jStI1TF6v0A2EvGTw0hLZXHmhO7xxHmbJHOskJMwIvjyS+77
kVWEKNzJJobGpz/ah3ua6Nq2z1ynzUrwKU23b2ChzHSlWYgq36rlQBhEG9gtrDSf
goEa995pOwsmA77PckaVHiuFYLN1RPLcYVXYVmjg4c2DWAyOsFwC8rHuTFwldGyA
XsYgLHCj6d+iSy+5vMfA90fLijMbV4Jnn8yu3MNqEXOopwE5I61VcFNXdIjxElOq
UipXXxASaeDjW6Be1uEUYfHnmlrJP+4AK0RWmsUpe4h+RmxN59oSRq1icm/jb1pv
Y1ezjq9nmXPBlUR1+ynJD8SYu3m+OnAsnmKKYiiRe6s5+5mEVn7dG9rKQf/RJtSm
fVIIG30iw2AhbQ7Nit2sqnmTZSYntex/2e8MozTNf7pdx8qGL9IuL0Us1A0D49dZ
1LjFqqj22p2/BsRoxYkdbzggkw/dZC/Q54cVp9AX7EV7uRkUHWYg2d52M9Rw0m+Z
xlDI/L4gPUV18jg3f4y8XBUTOSAFfrq0Kj/5/43kVRgtbUh2QwP/BvAvI7FecA1L
84ncyF6GRs4lv0iNj9XV3QE0zqkZM/aIhA5CJc5xCbB1jMOFdIw4gSe6zQXKRp6g
Qi+CH1XVlPzozy5Zwz/Z0Pwfc1FFh5GOdScI/NjuLsSE90qK1kTLBTIHEAZgG/pK
gl5Sfd3YbRpKVnUXNP2yFO3UgSpyrUq99P6AS0cy4Njs975/ny6sZoHXjTjHl7Vh
a4/zwq02bk10y8XqWZaNb4pRsxXbv+tYaV2bXCByPE86/pDQoS0tb9L7bQv3V1TT
e+w7vh7oXZ1fGWU8jFFHGIwozyi2mbgJ7GWI1f+RJT23MNiEVMxKxNls7W9tSZ7I
55CdhNsj5SOyj0hqhz1TfA5/zfIXus650nXISDnAxGTZDOHKZmRFOlngLPmBxP/9
OZfJeNDr3P4EFZYIw7ZU2475qDFMJO/UVRx7iXWQmZ5Euz0ao7ty/JLvMTDDH0EO
5gFWf7O3xdIfKoiTuw8U1wzwMRE4xYQ5uNz1Dq/OWGkrPXjV0OTbimtXryhxM49Q
d/scKyQl8DQUr3Tbcu97IhImmiNzDdFC3FQA96DtV4BNzGvp5u4CAT01FzjE1yWH
6y5L5I7rnOfdcXinReeXIIT4G8t+C58dp0kgzwHs3z20iS8qVoTl9mZn/6BdObTq
q8ILGXMZkWteXrXR/Fg5fHEBJ2aMUDDzlhiJmiaffSFHpu6Lftxv1bW5IUbnTfCC
yM6rQ6FSGRmIZPOSiuvvN46SEALldpBqlJUGN4CwI2XwX1ZW1XOHOBBEon3JSYFg
q/Rzjk+RqgiWQNUNyQTJ4Btv52gqqHQLOYDmrPg3hwLDrs277wvTOfWnPptarlob
4D1l6QFPmJp73y/iFY211iXrIHM5/xSXvK1hQRERPv0CTyX9ZLIQrjx55DGR5y4c
yvbaxltB3x2kd/XYI0YUFKEBQnslgd5n6PwMubA6CHNvlaVOQojrI4Aixgh0X2+n
HZscPI5YsBXlifOFjBjQpG06U1E4S0VKummUqMRyCDNXLF2J0qVWwzODTiz6F6vU
sH3ph88KTUQcdnwR+PGKd9mdxUgexSvjbbBbLLySxob+fjyycFmll7WaaPEd5yEK
UXn4D/XN5l2ULCaq6fJ1w/LTYGAX2+cipU1QZQ1HYiZK/nmKSixvJdCDVhqBAnxr
ocwe1XYjYJRIYrVVxH75uJkSP4/seceUz5f+ZkGFv5TbccxVthNASgyNydW8mG4A
CbxvzkoTSvfbI5E7sPvPhtBRPSHiA9+N8gxIsO/mVF1FJDqqSeNLBUeBcIllSXdQ
U4PNCu+p2mGgGMy0XvvOhNCvmwWgpWfflBJXZlIgIqVBgTeHaXYau4QmGMw0U5AY
8F/2OSEIzaYS6wh1ZlFPvyfORF4tt5N6zyuIzp2C8TBL0Zy/Q7Th7Gr6ElJcsYe+
BKxQIP8issHqBCWUBFrgNwxkWUx05maXiXOQyuEuilTWGSUOsxYqBJ6oXIOQ4F4f
GlsUukO54wwwZoRiEdrgap8W68EE23cTKAGy09OqGWKN0Gdl66tGxea/4gEWhoxB
+9twcf+B4Dm/sML1fAWZyi2RtFskQ/WZr5CCbTSpIAHLphjQTpOVqAv7sksPeGA1
ft7VRGEoG05vS/7jGSBq9l7HWqoZjwPLcObKeeT4NEHZMozHaBAruRXXylYhTMA7
gm5QOLQk2i4KArzvGdVhzxDUjtUQGZ2A0rg/b/rXWN89fSoPWNFBx+VNYgOwlxZo
C2OWu+8+HjvGVEjl3giqvTkXau0itBCixWJ4iT2oMwTe5B6rp5bIGFE9x67heE6o
UtxXbkEC0fun5ce9ePVwLVdY5wpcNxUBv3ndsTsSGnAt65SQuuvCoJLB8ATwuTlC
Ah6TRg5pjMNtTg7qhC22xbV3QBLK9+z8DBemnulyviTN3UqHG/kd3Eqypv/RMSfc
NAVFMEVFZ/n0pyCu106alEP/PT+SzopDI3+2qJqw2bizouS5/+bd8aR6DILcSXcB
huYIlIPrw7BslDNarSA9BFx+FSLyJOmvMmzMlNmlAU5QLmNrjQ3GyEBUjASMNJVU
ahVs+vvY202BEVw3IPpdd+HWBhlqo9BJAsdZh6hJ3rYcx6YxQKSsik6mVq5dGltb
d0YJQEi/ov9D4TbZ3+NzDi5dWOIFPygOGynj72sXkPuArjHedIaewfV4uJJuhum7
B5I9EvVaH9Iz0tEv9996D0Rwsll5VZjCHVnV9pNSL1fwIzv9mkBZVHvsg8+dE9YX
PeUR8lcexK/lMwQFvYOL2IugaqCuVQfk3C+NNYom9Q9pfdhOOuQk0aeIvrZ8A0Ii
Yxc28og4FvnPtEyI5EhF40iHo0wWxq+rOHltK1SWzYwA0C1Do5rusdG+KjyQ50QO
CLlIowH5gs4ML+GDSESfJ819KBfXqPbJN/7JjMuVDSbvujG1DfItI+yXZm4jglMk
ITd6kEb6T002h7EDPt807eoy4icfWUH+FWhhhX3/XYPCj1lOMTIopaixXEuaQr+Q
hlpwLOWbXhvbc+WwliljjqmSbqvy7jpMzNCE0a25JqUBSBFXBjKRpVHMg6P1Uj05
bxJf8w6f/LpSnXajq2/CQVH/9fSJ8YRh/TtaTDTBjszd3IqujoFpQlBjLg2ugXfo
YQfCpajaX1GtLe5Z4iHT9oO6oTCOeVRy94eL34KAVINfaKpoZGz8udKKJka/CNmX
23sPMkMvM18f9TaMAUfnikIRT4s5Rt1fmz7914JH4XshKAxYnFmHd/VmeISEpVEM
tsEZuGcvLVN+lXAQvLasd6FJ86rBIvqs7hKgAmZe1ig2SiYvBgEKoB/NOzmdcr95
ztIBJ0RcY0R77CGdxsix5TpEHDL9bI53UV0b+vGd/aekGGBwfH8tPZF7mbo2A0aq
JWRORZYnLjiB52R8q9cI80U83oTYl+WzyDYqIJXp1aMfBAA5MAlIRyTEIRMk7I63
xuJjCjo2Rd6RykB4sDvxnqsUOxuBBiXXRK+BwzJlhb1IhNe3dQo9V4q9HI3n8DVi
0sZboA0hR7MNKT17tPp0Q8wdQP9fzjgs8Tona2SOAkJkvJZEBAaGMyu8EA3omZXX
ReJHiYxJ8Ld2KcqQBSnC8k60JpHZySSBhB60UdPgt/Ilg013etVIDqyxXYuC0WgR
qgAm/FEbtyrvPC7rvSTVBeh9UfmCCoTwGFG6nkmiPs3Ma05f+xPHRd34sJhlMUA7
UUYnxV9CMmop/mIdrppM58GO8nx8+lpqWzLwAv0RGbaPjIWsHWs9n/I55PKES6IX
tDEhVnJPxOHn7u8/feFqMroohN+Y8II6kJrIGHbtyPgugDfvd1gVUDh72RMwtYSb
u0P9vw9tjXWyO1UL6Sm9JZdorj7z01JzD1AGD39olNQ9MquhFxnCMIe0oWWvLyTt
1h5+37S+evgnCDSS12PHvDUTe8mtTD24vSreeyKmMkd0NCul+atFOxedEElsWQbI
MrzNygwidBLrxGjvW/Rv8kbP4lC7zC0nRMmQ2C8hpsM4UAXtT+nemlCazcr3pbDI
7XoFpbGVL8v9vWLFIV+hNjmPy4LbL/ssAvqhYsD/eLVXN3dnyuUPaEy06sB8hrO6
ueWBDg8g/hsHPinhoI6+h7FuB9Byi9aWM/O0p88ly2IwRQHVx8nzclI5Xent8gHQ
XTNaVIXVecWZoFysGeCgCTbNC9k3K/aZOwQVHlU9+6yrDagEjiXYFVX+iJOwhofp
f9UG4m3kzFoa0EI91NiXApCLo/5Jyng/P3TiVwb3V8zC1vA4paCoEcTbO5R5+Rif
ifUyhqnDD4+sU+31l0pgdJlqFQTY46yJqjX7zyIBaGUwTYZnRWc23rScIKpjF6UX
6bnZf4FwZS0JDWDgoNhaHy/qZS0bsAy66RQbvcnDLIB1ZwdXl+tvbRyo6WoJytgu
AlGSP0Dr2I+BZbWMKbTQX6erwNxfl77ZfQfHuzF3l1qMd+6i3P7oNT7ObAZdqlQw
bn5d8fen3kpCXLkzXv9D4YZxW6ezyjBGbtfeTZJTSApahKu9/JpfDYZardFENSK8
CsxrWgKSZA0FFuiDt415HutXME1MnZFYIxwEeNtgY0zReeLvkXipeccZ00pLbJGH
OGVUACeFdpIQ1RZhrpRTm5g+7t8NVJoqYnggZR86TjSksE/AgJKZVoOqkJsDkaGZ
v8dhOjjNZ2pnQZel87FTHi4BVsL7T3AK/zMh5vVHREww8IqLOLY7K/bwyYOM2vCT
Iv0sipfH4AYlN9qhzK3vPtBBFMNsqTfopr/FplYLlG3aXRSxIyLRGRqpsKgS6Qo+
AqzF+9KsciEl9jeGgLJQaxgB1if1CR2Z0Phisc31ZlzwtavcQ6oKBfV0Z1P1NV+d
81dLPW9LXQKNtGk2dj/6F31ZrPURF6zUfgr40LO4v4UFRec6M8lgDI+2986nUZg+
959aHoQYgGFbaRi8JCW5wnp/G3tg0rpgB13F1ul3zqfnCDDAuzOkQT6JNVjlqjEJ
jU8AMUIpFnKQt9EKpbt1Wv5GDcjx0rZYHxLvbK/14i2/MGG1Qk+j1wKB2fFTRGrF
IdbIiKS8i4MkABM0172PmNNmtzpCJ1OaCZuqJ8RSmY78WhJl60R0D752mImIY9zf
YUWHrlCcQtCxbU6MYsBeqk158ZZ8RZgaWOv6DRvkfqAOIpUjtkM+kVlG3NBqq5SI
FdsQ1EkqoQi60Xzl1Hy9aIEC7DVu8wU5Ml8vZejMNXIPvPTHp16nh1isq2bVz1dn
jZwVEn7jJ4sFQ5S6SgVKeWZYfKcRjMZFVgjmDSvm9Zqlk745XYrHQ2BaG4SaNZgr
GeGx+bwSxkV/6Waqcrk4blSy/BynSwBWW/ToYC77LI/MLQytif0Ghc6z8X5eVDt3
VEEH20XiFgWtLE1WZkZRTXLTleWTLA0xe/zyWnkJUUPiQo2AfYSPQQOif5DEG+7p
k8oetbOuArXcEXJ0Krz+Mya0J2tDPbXHqu1rcUYUf/7ce2RCla1VDyTLl0l2KC5f
OL6q3u9Fj15CzmfhI/Kr/OO89I16EwhQ7hcw8HzsxTB4Nk/cZB5yS41re4ZoHIs+
JEgp+GKT1uGiztomozWsQzOKqgVCBtpVxLWuqeU7bnXFYr8UsMC8cEyvLIWbUsva
RVYksGPGE8wR4OTg6wrdns+RbGog5yT8jxdh+iSZRoBoeUrcGlggcrRD/KSGz/l4
z0bmUjzQyOG5IC+tsQCpWb+Tci/PjmHlwADpmR+1OH0wVfvLPFHoHTLn4WHUAytg
hSJYbDJ81rTTKTFVHGyKue0lPsfV6Pc89Zyf2KFNELjmlIxB4HJPbYjMORnREo0L
4x/z3P5H+RUp/+TCu8cAxK7QrlljlDklm+n5tES1REomjJXmG6g7vA+4/k7keK0w
Mw3xkc3PCGfOjDRrkeOEHUmdfgGosHnbJc40V8VaIBtwAQrr7qBPRIjtIZnNHtsZ
EICVJw/qcCyY09s4xEF2cdorRYdtwxuQ7VbzR99I5flpkAKKUDqnynCRmonSfp4B
qrZlDQYlTMCE7/n5PaKBmCaJ8gJc2UodLkww80VUYhCf+aBrKI4bZb6GnYT9aP3r
2qgEKYhikNZdM/Se/2/hbMVV+yCNvRekalDnHbzetWbnAwxdDAhGHOE7SnO/UgjA
r/u716wr766fNl3lwzVtKey+DyW1C07CL9i4EiWnBdVvuB7HksOIKyBev337oL9O
mvdnLcxskpb/5+Ok8Pds6ZDX5r0kILzJVhN0DnaQfIkhgUij4mJeZmzbQTmUd49J
65eWUCf1O2vh+Z5xGQNsrvh6ULE/JKNUvOXOUYYvvmTN0aTh1W7mEuoeiKbi30Bj
5xBpWDpP/JfWTJi8QaIpxo3T2WJR1jU6K8GFrjUfh7ZWfNCi14+aqrQ3qf4wM7sA
ev9VnEm/0a6wSnVDhJiXqYnwkC4NqN6+vL1JXGoPiaVu2Ffj/OVSYji83iu0OTdr
qqhqwI4z8iucLpndmGMNodaqES+R1s5J6Wmq9d4bY+sovLCok5onhAgtB3srzFS+
LS+Tu3jA/yImsTGJt+AsvzNl9X8KmniPPr3m6QDEdXG6u4E+Wfx6Nsm1+tR9NybF
LFaYrhgg59eHgJrtTq9lNhFT+mq+rywlT8MLWp1XeyHfOoK9E3ERGMaQTG2yXo1b
CItkzWH6yMn7RWyBqGUNN+YTvGBEms1hauINj7ygA25lyuHAW85KEXvShav5Qmph
7HNaThgUGDjVkGR77CnAwAdj48qEG/XGuDRgvLvvndHay8ZiNuI8gTb/tucxpbem
x+90crvxutmBJK5ph2SWMfQ/w1Wp6mCPkDz/F4A8fnpHJZqMUXWszwgZDTHkY8ji
jZG+Lwf1nvWv5QwmgLHZ+/3G9r7NPUdru8wYMVMptIZiFB06Vx1QsoK6CC44NIyd
5vhdXWGcThFAzVDTGJx+flDuzaKaMkT+a57eVows3Za/klkVndd1y78HnvJRVDqK
JcUTMOwL/F42y9ADD8neRuQSYvh9BlQvV+eihPQYBDa7ep2VkDJ9vY1+eeQJW6ID
PCysjPvLri5/qKPyRczDmxcSi7nh5YXxhjXd5X4VJ8ilF8mqHNgFx1T/ZSrTdzaF
+XWb+OR6RPm1gYySUrKQrmRFONz2WWZmftORxXaYaFILXK2AHVE8CLQcpoPDasTM
lGbBj1J/cE+lx+mBqO855ranciURTWpN+2R/EoQfLyhsnFSK9hO8xd8VWb65CIMI
OxB49hhP1kKHNcTXOZcYei9EmF4HF0LDYU5EyAIexNeA8f4rsoo3MLKy4R9gpmVk
93kib9DR//3tAP4nvVn9hbMnazxjIOs9QT6q6EedI+gSESWdHEvM+w+oFYYK/KAG
o8llPqntRAxUmK/FwF5tPuqHcWtbaUwz67dSb2wpKiWtDV95pVJr0P/mAwHA9Qhe
ZQSb4shWYIifJH1j14eeg7Apw0eCwGTxLrXKIz/borJqoOFSWw7Dov13AmLQiQO0
lnt1GnJDEEDUt8Tb1zuUbu8f7V3aHNUx3laeNjLvNgW84e6RxhL9Xa6eopQY3UwV
zrFtk2zEDpu4qK4Azojxj6FjRZH/CTY+shqEK5q2bpRXS5mWzki2xmSpTFx5PPuO
LXOXwrAPDZF3ND5Hlo9X9eWCeTbTBbAYS56OtSugsJa0VdqYfNeGL1jYX61hDy6R
BnAYngLuk4qZxBi6giJ1AWsLgIUQSyQ19NIP6Eu7dE9rUw4OkjWdW6V70Rtl+KY2
vyp5biKL3jYsj95LXtFxKRockYz9emC6kKAi4z5ErJHDT9zAPzrAWuKtSJNF09H9
wiYqE2lEEA2jpDFxYkmQMA4wFhy6vP94uSUCOV68qr+78Ijrcg0/KAzMKlDCSUyG
2CYvsB6S5X6uCSSB5Jt80uOWNM1eJbywG7InGrQ9a8oEqYRLEUe5YxNMneh9yXWe
FaM1VKr/zcfTs8nzI4NHgRhQEmmlKNfyL80aLE49bwUfaAQf5t7qSkvgsXCifiml
lRBBqJAI9u/gMHVtTifnTMqa4BV2+3hR2pjdVWbJi3C6QH0Qapsz+sEFNup4T0K/
jBxap9+H+qTtNLkY58BVifdcAQ7GTJq5G3YJMnneCbhD6SBS0gf/hvdJQGlKVOLs
TDa3yAp6+ylrBvIHKNZ4nejAsVi2PZV55eGtwgk7gpvVoYJGkW3qMSNL/uP3DfPX
mPoaZPwYqbxRwIq/yu/OoTXLOiCIelROjwkr6fN5akTyoU/tV0f8xuOH/aHnEewi
ZrDSDnaw2uQ0XwyfZ9Tvwpn0DO+hTLbHx+QTt6i3bXwVltRJfoEaC52OFcoMcyNA
F7aGWUC6bnbZPSw1rcXOziFGJTC3sDbM2LxH8p0ciGfGccrVZICIsYcsQk0hoxu5
tsx7AIeMVgol7NTVs5GykiwQSYvxOiXg4VyD+oaGlgfewZvItpHKovULR8ALWfgS
134HBN937TlP3g4vlDj66aZJdJosxRxH9Wkl/EKAeI0b1K+ahY175yzKeARj3qQ1
U23jBxYyctIoM1/HwOA7n7Sdb86SeDDXJtJAeWf+nOAQuS398jz2n+p+c2+lXWBq
UtZDtIeZncYAha/qA/Ly/AIDV/eGEDs/+DgaJl4wQN7dqWb9lW+JGuEjbjfGvmqW
DJUPNeET3EPTxMEmPAseXH53Wiop+zyAL9LjkJdgAF8avXgI7/EnEWcLo0uyTWBb
tVlA3jL0Iq5ieuKhUuOiJ3UU+I7PB/fSjz2A2u9dbQUu/0JhwNWgeps7eZARxS4Q
lK1aghtB3PyVGjMhT4hUK7heqUD4n7emWGRC+CbJ1XVdYqwSVhN+Yxn7ozshfCTO
arOgoxNd9ZzmbLWi/+JFzvtd8acmqkJu/CnCQjd8EBWu9oGB94UkCP0h8VJa3Xxt
6TnbYCTmelyX5lmvn9WuH4NSe5rRDYeXoPGXEkwA/IX5IVKtzZa1SBWbM7XksCxZ
k7uFukaJz8SptymaCiATSkZcPJD3UD9Gp8FmhF/V3XCrCJnfEkLiWI84c4BiQGrb
YjQK0oGJBydn2ZNT4ZekUh581GY9w6g/2H5opiuMEevqsdvmXf86B7QyhuW2gr7u
i4Y3JAZ9acc/OkrdxKEl/tMvjWl1RZp4IAB2nWc2Ur2mh6LJniy+DyqV7HVU97uQ
we81jVMO8kkuvhA0puseqHXGTQGBDQMPNCXsd7kGSiwKLmg9ICV+8+EbzoofVPcH
yDrvvhK/prSo3KB93SbOheLR2mumcHmdm+10JfXO+Y2R+FcFyTpVfYiAx3RFfUuG
/LX8tWU+3x6fDB6CXUUyxuT9ILUJh7mI1ObrWWJtNjJChBr3XqjhT3CgDcO8qcGp
dGLCHNNuq/PVWEFDubsD0DBgFF5vHYrRBE5qxQTdDKwQubFeyh31yfTWnrsDFuic
EX3i8PQTRn9v63+yEcKZdE9BoXgtEITKD9rZ1+ODf0MdWvV5PuqYAkQgtfspMSvE
mCjPC8klfwwA/TOLTlO0N4S6BUsbsiSIbwVfhItr0cZQfPrSD6pBDzdAkl+qZ9uH
kTsWI9bSwGLYgWpswUQpr3FE5vPMYt4zc+FkxtCzLuzLOLKbRYe+H6r/0lPLgIw7
YNLLtCYYfHtBaH2cQlQO4sMM8HfAwYA3CUQQLnXkVWSlyW9saPT/7ehketx4r9aX
8droYtwjlWT5NWsnlyKKc2JoKfGpzQVc83NEQp/YyhvqbDVNh6P4FNcYpCmbBhZE
NaBVLdtUoK8wnTf1NuSxeEAS0E2EIUZfW+e5dwXVIMpQeBnIZ8UrNJbcMQ1H3QpF
RSCVTUScBNQO+TjehXsYI9hLbSaywNfw+cfTAbaLo9KJDIvJNKoiYHcfX56l2erT
r9cGJ0Ps+ouBW/2wsvGtzgZ4Yl7wPho3d2l4ll6aod9esF/OJFiPGS3q+cNmIP/o
glTyhxZFLcRFVFNrF1Nd+VjmKOdwigdeCTeZ1rayqB2Crs2jiRoLexHGEwAnpgOg
c62s/5MI5AXm4Ywn4Rja8w+KG/Nnk6/00IJvpzK0HCQ+slmhDu9daDPT0hFyr1yx
8NL5oqY01uJEisODy8xa8MWYm2ToSPS+Jq33qBWwHZzShplhbQak0g2WkTfaXJlC
Vt4+mMFxBqiF4Z/rgAyyfLTDxDDysg7X56K6Ec2fbBEikTrbVvEZtXqqdtTxFbOk
3ps0iUzzIfsmVPjauJ4BcAxo0NO606nvAuWCgP0lKGkA2r1BkgR9EDvqfh1VQ+qi
r9g1KC7+I2x/2U5wiv4NSj5WpCdxLnFl6Lofxv7lxmwN4ryO7RdXpUESnJnRfw/L
J4LoQMN5qPmMOWlZg/A9wYWyPsIvjlfyof3J34/NObwPcG44XHzB+JdIAY1iylWN
H+FtVlsyHKOokVw1eunkJ5tXqhr6EHecrorfiZVIad1f1fJ5T1gntliY4tFszTXY
Jkv/ny3TOglhYB2AN+WW//7XS6H4WB3A6Y9i6MIL+1C+h68HAncCpVpQRJxQhrMx
aDiWzv56mmJjK4bSPt5FX4JbS8wQlMwsosABQ0e9pBE9Xaq5+3EIEZ+eySDVwYPj
ymQjLoUbKlMa7w99AVGsi/KgewtRgUQdTJrDnmLiXwsV/bh+S1z6ghhwGJWY6Jed
OXZQw8UPBwo3Ch3CvDlAD/Zj5zOiNRIAWQMsKGuPCTXqYnzeXjGOv6Ewwh4Wk9MT
eE4wOxcAX0qji7CW5aphoBlX0XlFpjS8NXoaTDe6GQABn/L55LBi1vmVurc1g6P4
clsv+2jazp7Cqtf5Zs5+Xj9E4oh8uzIx6mLRH7AbIOr3iXLr9YeOkDvsKTUNOspf
n051fuyo2HRus2P3JDbfwu3t/vZGjMOPJ4VKPM4cupvvHZNKuPIymOBsyShwV+5h
KrIID07GB38tasPt9FpNUPec5G6zHdygAFmbGKN+FY/EFCUBdM4npUhTQcbRNKFq
hGXXwtTB+p55jwSBHMvco78dYXeQScG2XJRtCaShCZwHCL7yH9fAhgPR0y1O5f5a
RZVid7YNQCHKzjmRCmhwQElZOJeb0YInD4TzAt+e38+itDAkngGeaCfY1OyoLKRk
249cCur0LnMjjobladQ02d27B8GMpLcjejJ4XvlRJz2TL4/Q4LeimBnBs1y7FlsR
jwgAr09rRZl6zFIpD8IQkWOucOm4g+oDCoGaZKrrUfwDrV3XekmPBvMjswsAXyCj
DeCzsr/Ws3hsuXntPeU3BacCKSTaniz2ViUzcGwkeTzGF/qKDbqSPwJcsj31me7w
elwHzdF8Hl5oX30yglWcJCf4qExctUnAp4IJhWwdHo8ovgorYuEj/zdMZYo0t7wU
V4QwYlp21O3i6Fu9BSEu5YUbyVgHW2q5XQv9TcS2vQqKvohJX32mQu0B9Xyr5GVK
PPqObSpCRGMrPAJEsPdz2ZQSc+kLg8nCPiWW0++03yyx5EdUoZeU3XHCgDIwrqJz
/ZItk1EE7HKvJma9ZraVtq7hy/Ade2iZVNDQ+0za9MPO1/bMJ75O+Gpj8cWtu37y
bhis6jrxPIRkHlSkQSwbyAvcfab2mQ68az5pGoUhqIJXaxczdtb8lHBZ8gY4lPYq
ZIZKR2f+xW1EtXHGGGk37EXJjQZ+7IEtxelie6AwPZbi1kI0U1IB3aUQcMZCdD60
h8shS0+uslsZKgVYbzTex6W0rC2Y5aSHjM7K7IvSNxb1z3e4vHv5sf3eCNB4LO3a
3B35rgBJi27WpV42JTgMC8pdut/XyY2K/jwDCw2B+/GeJ3TrXffqYtwyCfmVEZHJ
YiAi3oFU7GtFPv4IZsGLsxYRcpOmadGyUc3kArIEEWIhOcCFTddr8HxcGWMLtnPH
85z0VI0wQKaYK8wuLd8EC7uE2bB3ox4HHOwGf5GCyM/FGYo/aQdkGpf4xJ6C64hv
Hi0g2t1GHHXO2aKDvofw/KsjczC2nw31+a7YVxRmlyNu8cMhpEF26boYqBC+N9av
cetZxfoZtA+ciUcKtyYTfQDdAad2oJgzy8Xm24NW+o/siPToG08TcjhHx8LR9vY6
EDvp3Mx7YY/c/Q3K3/RCXYqxAEV3ET2H+/r48CoVY9lZSafEYZBYSp9fjwrswVaa
0LxatJy/0uOsZHj7MryVk58slSG89iavHROM+GJiCySMftl/kOmtMEamF937b8gH
uXPZXxIJRN2uT/HzuE0qYJ5Bcvmt0exAiKhTqStrrwudy7KEFYUgf79DxmezEZ37
R0MLWbHI7UjgfDCaEh4fr0pnllRHbSvBWiceQuGYmaFPK5Ly+Qfv+iumsvOvvuo9
vJL7rnXMfmT9B/1fs9Myqe+RqLEOraQLeQdFM5j3AVaAC2Xd5XpWYcEB1WnsAfs6
ztxJc1ELKwXLprH0+BaTXqbSKeGwpEDJm2ywyr0f6LnyNPLMDgt/HAKFdLYl0I9j
Or9BuhjW9VKPCTbNB6Cg+r2xVtFeSjKuHd+b5FW+X+Phzf4HGYJUPQ2a+ElomAMA
ahArhy1nJkf/YsKpbCVAb9qPEEEHYolnKewK7fRZjZuE84f9cW2WAGc8+8JIXfAP
CE0vlyr/vTqOtOybU6bIdHInXPQJbpkk0jRtC8QMvqi0qRQzA5jarNfxT5IFRVte
4KJOMSXgh4WbDDNPQgF9vU3zBlQ7lXRF2u4Y3gYDwLnGIShaoiwVVOGrm+ygjMjt
5HpXYRgHwCpQR67Lh1x2zf8eK9ZKcIs8v7oejJDGqTI6d1nIsDmVR6vYJ6kAI4X5
Tc5xGirT2KAo0hbU2XrBLk3IT1sU0Nxwu2CLn9aaqoVU+dhAXPF4HDfYd7SPYmVx
cfWblWrSg+zIra/pWp32FZ8mRd2HZes9ZYyGqsfOLU5Sqvixa3FzjYnUkmL+uH5u
vyK58rTdwbGapkkOdlrhKarMZzQa/3oFVpkPaZxIcxvc5khaXv3MV0RHCqPSg4ia
Jd8i2ka46jESw0qvsOlZy3HWY0QGRg4T6RCdUgrYx4k2HrWhn6KzWxKFTex0m4O6
hUtZF6Y5q6W5J6ksXEjOuk4bIa03/Id6OYtRW8vzAQqRNlhfgQebnfFjzo6jqLiS
RkQapQEy7g0zjx20pAgjkd/y3ADUdyXc29996pgr5KsoSkRcSjkuMbAh8uazgW0U
6Mg/yTRbwWuK3996x01qBHHM0f1sQjGUW/JJ1dXKX9YjBTKvbIjYeau1VYM3xKJR
+wCRLd5qFjYauVJOFs2745bayHjQoexml4umhWrbK3Y1YMub8IQXKsF8zfRhEgA7
Tk69DajRJDWd9Wf1FZm99WoIahzgykqyK/qI1sU4sNtNHTiVSdRW7b65n6UDgjyn
vaAWVMxvsBvNPyw2vad6hsTvXQrKdzp9CKPoMsI3tnsx5QSOzZarg/r2j/TlItBp
bMVTohPwtLO8CuFpRSp4OrH0alNkpU10rv0SG7/POZ6QVrYjRt+oSKRYymjGzhHu
nUV+QUnQNJGymiy6ZnIJlL46GaI6EJdoMIcES7ocUTSkTj9J9BzxPz/BoWotfeg1
LBYgeNA0SK0zipHwvkOJVlXBhKEdaZBw7zO1J92wRAim4TO5/ZmeJpRU3d7alZ0G
c92jC32nVivJsgrO54Hd0LHImwdWHiD28HtopXJpcGKY/uIytIr/hOKujhCafxtN
wecE0AUqvvFTQ5k+UOt+bIWlza3mJ6twzj8IhR5A/CGA6b5P/ein++8yB0wuQbr4
dIwuOcHn3lf+DcvJWtdmKc4dPNAycbi54Iz4lPGo8DBbNm6OvNiSmhDing3zFXiX
/zpCE4RdBXodAJIkzzSRtM9eD40fgwVqNcCal1kZdoVQYARpyt27SdgwLZ65RV/b
tMwXmX1NDfDtoMFfAUTRwF+S7jv2i+7+puhA1UfBLJT1AlR6Bdw02DDOYJG1acg2
pjbvikyS8IltnRo4VwiJvbgBP8D1S69VrWjpyYwb3ykAKGHNvqgBOQ5YuyxIK/Mx
6NABbAxJcT9R4kCErjHwH1aSIf6FFHcmfyY32as9YFaBkNB0JVt+JhbT042R6g2B
gsWmiXN0ZHgQm66KOuYev4zCk4MYOS5nd+xfxO2nqrPJ55zLjiUAEqzSL++6YlNp
F4lvs5zEx6mkeKC7T7EeYbJg8GjCr1NrT0mnQ+RAM42rihtc8aUOgzk3m71Ir3od
6n04Qs0L/pGOwiZrzUeMm/iHaNkOUCDCPWJw+cufvVAcUSzNS4WbbL9XaRLu5dd3
KZF3fTyEJhbiGHAkj1sS3sgXFXpRyJgFZ5ZsZSUcyGMs0M/cn9lf/GBX64MtkVHb
Ttr0SQZtjwWCYVoN7E4gCGxGTN2YUBP00jkXc1iHF7TjPwqO4Qx2D6ZG0uOC8EGI
pcd+sNCYri7rcyff5hN26IGHZ4Ok14R4FswtlxR2OK/pdKetfAbn/iAqqcwXZNfi
Ea3HcQ2Ptsj2Sj/xLgHyccVl4T+2fI5ZoMAEgpQCc5wxdcaADFdbLSs8rA7toOea
Zp6O01GAYbPihlJodq24jBAXcxiRl9zBFQaL8tqIqhLUfZc4WLTVQUwZKv1aGKNf
UpZA4GXQzN4rBPbf2UvIv0siCk3yz/t87TqsLvt9LLAcU9BhHNNonyOeeRkvXuvz
8Gk4zOUOU1Tjg+FTTmLJL8n0L0CaeyHxtv1/bQPiBcb5LMjsbWHUBU0XN60OoAYm
5g5F4uc7KEsfiG/6DTFC4TbXplzFJT0mfJN6jGZ7HSfMVhtsRBsaJEZIGG1YKGfm
AG/AsQDq86OkBm4f/YNjTSg4zUAKJKgs6ckYwy43Nm3icBQaJbzoInhNQI7vrTpG
oUMVi14cKE9qTJXiy5hvQ44LyR8gQQ/rOU3/VdNQ3y46obtBr4AEwqm3LupuoD80
ywLfZ+PvLLtOUNfnatyIiFQv910jykeB+KJ/Y8ggQoNmsZx/vGF8Nz+cfpc6wQ1X
EFfwiQER+l18oU+BIWluD7a7n1TQc5XyhusMBRyjpmqtTxihbE6HF8qYkZQeyWRy
HxYmb5EyS2gNi+DV2GWEPFOLXUcvYjQulfyYz8LcNetqXkkR3DFjnscON2F8sDfH
imrfUfsots0ZZyJ+9RgIcZWDOgfmhCWfq//z7wZo4BEhHWnApqEsMg2FvnE7mXVK
joTc7WxPOt6zJntK+vwEzFPVJaT/hQ8C2vDli6h8dx8g9u+DPZLE/gNW306itTkq
5RBTjcrmICYOzl2U9sqaLfd2GvmPIvpoGf9jreRm3jRqXU+07liXVrwsGW7lU47X
U6OeT2+IjJiV21CCLnSiFkH8q1ZxP3I1Jk6BQEdZ9ulslwnEKwQ3aDaRWfCbNEZo
7KSGaj+1pa7ZYWPIWdA8MnxwfrNgrJ8O8x+ahwaEcRQsGSV42ptILZpfUodd//Up
5jk2ty6qhj54qUOSuYw+Zjg+xzZI4GnKznpsyagWZ0phN7+GC7EDXOo5RZVLzmU8
jDIc9Q9gV19tldAYOgxX9UD3cojdyCg+qbQ7VPJ5a03ZUUg73GjPBp/4mU9leCHW
wFX1Rqk21/fdE7aVkCBkDABRfLUctekPCE2sSDiH8UZJ8WJcdDlXkibWBP6NSYcm
l3WTMAMrutTCbFLVLArVlz1EqWupFUvnkGxM+BlZZ9WUKT5Cvf76kIVP9UsrJxqk
kihdai4c571MxFLTkYT3ntC4kyGubou9RCMpXsZo2knKY5mEc9s7VBAgB7S74foI
ciToQH62nORT17xQdXo7/nkLkCM2tiEOEruab+ul80IO8A2NUZU3vbMTDuoFViKs
sg+GdpwBQzct7ShllGgHoM+Tikmrpxk07MFRPwAnL6l6xcDfKUuyyfP3CyzKFyb/
Oh9hUvGIqKJWK8WdySjAfeXkUEADhhHT/6eDG8qDDjE9DmVLczKUvJQiEdXC/ctN
2uEqxjiHjGivBCMdk1aGt7xpwj8ud8WsfGcaThO5GRBx3Y9bh11i8jMhvhyxiEP0
gFhwKKsC8z0uzQkUm07A0SLK3AcXW2aFzpwSW8k/T/GDwzYHpsFfTO2yH4vJbQEo
s/A5sMIx4duuiATHx1PDO8G3HHIG0+dprmKs2Azk2zu3/1rYn3PfVhpvxHMMaxtz
t07v6Kl3v9IzhG+RirrfX41/Q2ktGtQWut3u9Ec+336ToG3ssWHs5CAMnJLKbqHN
ncSD4fsDOHeVQGlVWJKKbBKKJncYyqFuUO7+P6Qojz9L2G22L1DQXUtzHCh5QPw6
8a2GRgUU1LPrNrQ5rIsoR6fu1F+5MxNSEKgixYTEqa0VOGdbQWT8e4etTz6iYYAK
aa9oVIZGVJ+A7We2hCsE4KHTs1uscFXJvmkYBjD1jhrpi9/sVf4yWKmHmHEzCJ2q
OCKgJutfqdRKc3IV63Rx1YioT6yfSRyrj3zUTEeyLrrSSPpwehEmlWZ7N2A+0tWT
gNHEJPC8QXdnxx8dhtVc3OKv7D1F9H1rmvSj9pyZ5fHU8Qg4le+hYnhxr74tae5O
Xwe97k90Uo846wrDjljq5ihxacNmBCl6OzynbMAoRi5nXqrlpCKFaZmDS4Nbd8nf
ZMXciq+L1bjnOz30cn2HkUI9YwBSLzBTCVbQhiqd2JVfgm8jEYTdWziKFIsS4sv7
/X11eH86ckYfUSwYoXdOsmtSAIqpPllBLEYayhAZZbXDr4DGq28EjLG42KfjSL5I
lj67lKA/9yALxwP848u6Lg3CCj5gIgDOUCkS79doPybkuixCmUDCdZqAZ9gxiqgD
708zrSTGOnVBLvG/I1ZiqXNIA/+E2Lp2xn/qWjwqirdl80yr9gNj9ApdHxZqbJru
4oro00rHMp9b7vgYfAdadwUgUtRlEm8z9j85iJoNcm+kH352KX9ymYrL5BMJEuW6
OPmOnuSXvxyEEJ7XVs7smTW8Si2ym0WgjTGrPQsn+7T0TwIECvKFCla3QBmbIvnR
cxOaoYEj+bmtxdNBRyhNemZW+XNIcItd/DzFeja+zFKFVmR+4AGl1PKByav/8qVU
LgPT11N5vd9+ha6+qyGUMq0guopBszPMUlkHI3rBvE9lmZq5EqvYTrCEusaeTeLG
baT4Bq9xRIIogWndwN6WybU/OK1ajDZwEBcWVD7tEDTO+AkkqZXFYG0REZ6gi171
zwj2dSYwY/nlYY68a/6RZH5PnYs+5VFoVyI/AkicbbgJv9isF+ufyp3WbMKcP9mA
Rg42AQthjhBvtoj7sfl1X2rR2ePZGuTANkh6vtCWzDSbCAjKR1Z/kb+oRjY4hWBx
Y+zonn7wyrjy4wHkbtUzfy51ud2qIoJrrYiI3jtN9Ojyy5JqjbcdoqygXBJ7drbw
Uc5CunIQb4h+Za6HYaO2ef+Z+xxTK/NtK1lNJIUWrsTxh56kOOuy3BM7xd18yTzI
9ffQPVCXks6je4k+mXM5ihwyaxh3BrymHwk5Bv45dNkPy1IcykzekfK/qacH1iQp
kIeFlrloae1Q7xEnwW8Wc/YsgntXz2OPZgUMDHM/2cJp6DPqfWlRY56WcitA0w+I
u/mGLyOYPdu8PXHoM020CNgpArXp3IjrlUXNUUFAjT2O4ljFn4iv/p0Q5Em5vD4L
c6aCGR3v2gzSFOTmSXFco5h0MLoiCXRdGxvR7iOFr9km0J/kSr4OWwe1321rbybm
nibQYXjedcKlBw1YS6ziyvX30pjLwmyMecZ4/rD+nke/p65T6BmCD+P0j6o1utn4
cLQQAG5oTxS0FED9mXFu9tP+RS1rlJAyAHsLX2sE+Fc6fDnlZ/kkWhLcsNUr92CG
GLmCQKUEdhBt2y25JCjyGsZ1O8VFZKDMbNMjGRWPwsIBn0lPrb3kZ7wHfBwyw5Vh
yz58wVn0DdCMMdcAzffUxkbhh8GliQiAKVbTI1IwWNDk+PJNgg4JX4fywEl4ZmR/
P7000B3Dm3vOU5sDvli2FKQy1YD9eAh7oDTJG4CYEagVWEqnBpmgo8IFoX2o1iiU
DG/EpJ3c3K1932dnNJzokeZXHHlkvlJRLylLL+yUzucRc4+P0i69wzwsoDHY/6Fz
W9MVb/Uh4qsBqH4wLcqLp/5eyOQbeS9rMQ1AjzuC031gQ9xJQfsN31/m1uJf6ys3
0Avxuzf4h8AKtJjd8Z5suCikJDB3WwUxE6cdJJWrZ7bX1nSFlzUERf73py55IrG8
sE6s8JD/Frk0QGetvLN8NNM/KWtJhx1N22XecNMzxqkdrhBjDGElM6+E9pbC3sn0
3ehvDNNTr2MohPitMaaF8YFF9QWQHDmE34NzfEZgr7QrGQnl39YibIwM+fg8/Cpd
WBVGuXdNUvP8tubE/DR4+iaCsbJwTwPnGsbwmR+PdMFhx2HkdlrS/jaxnGypka6s
EBVdDN1OxpbhwR+kFesPNXiXBiCKewThYMTgf+qy9QhbCGVxm7nHv0CohJ17o8nq
q2rZ7ymk3MLdxEe42rybRiYL15N/HfSeak9JMPTYa7otI9GOrRk3hw0bMaO97Gaj
nhKjn8+a9qVDIMSpEjzHxBYPOuW5MJcB278Km1rr7C+AXzRdGmTBPrYXH08XEh7F
Bv2dRm4k62jWHTypKjTIQ+QmxZIu8PRSYjrPlaqnV8xC2aF8RhBusqnM2x9EjoDG
VM31FXaswn4jYjZlrNnS4hSsfPxpjftmRAfvIgHIIsAFof/zblMo4or1JrBeRzsb
tRmcO4Bs41kwerQ5riahHSamoDaTZh1Kqab4UqNyN66gsva0c03C4xMGZdo0wHbp
QvBxbjGw35fIt50jWvVVYBjZi7qxnCR/OZJBFqUvW8kZ4J/A3rGZyWeGZUoGYDip
MFEJ8s0iky8ORcp6pHsLsvFDDPIpQBDyQBjRB1KZStWEtwksfyzcKuD0jttDfQqR
0Cb/9pDmkk2yK5DymRDR/k+iashXEdYv6VsCH7nGnq/mG2GmwHJnsAXhnGbzhwJG
jdmT0FhjpvRqhPPrj/uw6KzzK03F03oynlXmaj0UY2+yEAe+Zh+fqrAc+1tMZaCn
kRbc4zOZkpQC5d54VklLS0azM/Z3JEpVdD9mW63q0Qc4fZD0kOqteGHKd+xyF8yb
2zps/5yMdV1kEMvNO6GE8s/WO5vmA8zzqNR4AwDHEyOXOfmdYG/sAo4kKMbNqJ0m
nZIRno+z/DUi+liOTPHkO8EXFOF6HKw/Uyn9oa02Ae1PVfDGxLOsTLO6sSqAx53w
z7I0/ogKzXE1XeH57BMRennXBdFEIV2ArBLb7j0rQ27CQ4Sf6GVGXDCrPniJth/A
D32El8VEi3rmBXyYoI11PqQ8OZocUbwV/oFOwrtO7j1HHC/Rle1r7TgD7hH2thxe
0/iNxkDQr7ElNzHmgLhqD2XBNuM+eOcJ6NMp9GHORuC93r6J5nm1ZxXGBZkyjUxP
Fz63r8vHOHLjKr+cRHWzFcBmL5cIkUEiurrVOKgvu+g5vYVBs2PGld4caiXwftgi
FBnC2EFTkYpgfV9GGHN68VFOGGM9RLgaZ8I1v44RSKyNI7DK3F7kwK1zkw6W3Vvr
RdmMh6Co2kmtUBtByzJykHQHkrtrtc95Many4Izi3EMPA83Y0yy74iAszqUH5SJx
KzMcw8Mv2IX+XICSbIM4Rj8TqqgBgPWRuI3+JsTrELiSQcVOcLFH7rthRTmhYBlp
KsbuX9i38ENty8uptoe7Kh7+0bsUdPcrvNUlLEG6Sz1ygSpdMety+msAi136UADs
Z2FYvGCN/NCsMWflgQgZgTvxqMLCbc3mXiszH7s+FcE6scNJylLJDm7UTiWTJyX0
HkBKrCLV1WaKXEyaKkqXu7Eb0rwk7eaisqbvABNsW1uFA/EJK5LiDNuysqrK1BJG
Cg1+DEpiXe4Jsi/KHXU61Gk3tSvUwlnRxoVCRejWNpPhv52+yfCI8rdSUcbYdlCy
ZFR2IxPKE2cg/nNlWIHiFHiplUy9ijnnS76hA0Jr1439r3lTp9nlDdjvjj3bRvSQ
4cnX5aNE+4ALetA8slzo0ubWEIllSJFm8HYElHNi5xjHs56yrS4XFmMIv5VmqEi6
d26zW84fMLJTE01asc+qCSCjDo7y6ARXJc/Bx2Xf8JVml1TkoBfOE6cWtZpaTvFh
wKyWiYOd/nkcT7kPils8H58XGpf89jdw9Jf+w4jwel13pvgBdCli5ok/5W2nFsw0
x01rezT3Jvf/9NbGIxLmVhu/SV+a6q77F+greLpPceY+5UwAEH0qfewwl5erMch6
oAD/UU6NNI42vFaHhbNY5BRXDINDgoZ7dhU3w8i2wQP875PYdCpIjx7immsFBjai
wS3CqCXzE9aG4NRALpOJK64Uf9RjmCFwC903cxu3EXyKol2yb/C5r/IZ6FuaVdi3
yM5gVXcTL+LNnDsK82Tc9Yl/SNpc4ZtUx+B6SiaX81A=
`pragma protect end_protected
