// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:37 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
MrTrIZWo0X/6Zm7unDG0jfav+CHNpvfBueujzsxyqlx/MbrV/iR2t6trBKd/Elhx
97soLqub9Kt6qq2Hn4B1YSy/G+bINW5acq5fHSkFJtCSpg0Ye78cA3gsY1O9xgys
kKOhSzcaNEA7OcBZFcm3nEAJ3gPhEfWqbW40EMah1t4=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 34224)
BGwlnnulxrbx1+hpzxKLQyvdk/CfTGcjrWqKbI4AXQYqfmhcxaDOoGb0zNdfMb37
uwUCNWiyYraNfTxXS3BZxIDTUwHlcnLZgKFdTREyiRqeUj5+irXAATgPvvci6VfT
73r2oLYbGGquOzO2EZC3uiw2uzobsKCY75aZNbIR9r/GsWVou9HosQ6Uha0ghMtc
Qtr00fgYxZuCSbB5cVI0z48fgikIqGgr2cnThsIN4ky+sWeAUcZ6POBESY96n3Xb
eiLeBEIBXn7/qC3g1B3bAePakCBUey2Gw8rJgYZM/gWlWWejGDPJ0x7QlkqoeA3T
rUIyOD7OJ90TUQA8LqL2sJfMA4ZoRuvsvOLMsSd1x2dTNKAJIruePNP8AaMWUqIJ
EjIvI2nVIK351i7+kZOe8YfMWSN8b8cudpVEomLLTz7l+If6vTvuB1NEEvCoMPKC
SHFH1xzA6xmE0GY7z9hy2OF8JjLi69MDA2CbZlVTA2dSC4q9e3FyuMUHgd2tnSKy
dz813Rupmyqn4Gv/oFJcpmDBDjE6QTnv6cr4L2ArQ6HVJVRbZ2pFHD9D0Yr140sy
Ycc8NIvZpONFR0Xx1IYS7wpB8so3aYRMA0nM5SEn6Cv0iYi+iN0h2kj9W5lMnv8a
YwYN1w4s+AkFRtcuAxD7kUtC8Rq6zw/cyimOmLoPYFR4sjT6U+O+kBHxxleSyOyX
pXqFZBauMBMPsPtUk+U4s/xX35/DpUutOk35ICajuwo2IApz1kAU6TCUHNwOzV6Y
D2mJyrBaLM6uPwRfDgs90I1SHoeOtphw9fIetcc5gzDvkQoWg5ut41eYo3sabaRj
fGTZKn0bjhdaRZeWhs9gK0p7JDVmc4M82Q8PCz4JUAjiSTjNfFeQkjVi4bbWZlEO
/E9rSgK/JIdfeynBqCEBxJjMWfttXDPg+qF+azM8039WAai3xoJLZWif6adE5p4S
9xQauA7SaBEYQCfiTYqxZDBGis7z+5j8PE9mFIJWeNbTa/H2zEvD4kzSBO5FtxoC
+oEBGh0BAVuOlbB2l1UieuJKDGza6iGb4yxleIe+Pip+LW9oOOIsSwPLcDH+3Brm
JloYI3IL8W+Wvf8Zh4HBEgU+/gxYuwxTX6mV7ptMp2RcxCb7UULh+1/Z4+oydZ4f
kypGHKmuSlj9te91BWUKvjJ41k/1KV+6xGjOQWCJlg78I1a5DZcWdnI8tWepvjH+
Rcg4GphL3cjPt/Ze2QaXPDlMnXE0cVM6gHyt4nZHoGfoEeNW8iEPdd5G+BfcfAHa
VOsNIAIR6d3awlG8WGbzT6ANc14ti8AqkbsN3znzjuLDXzIoUJ97RTNGgUwYFJhP
wfpZlsitPmfBQCRkMLe5XfQjCVlbdk88ySFZfvUAiwL6AnO9CsirfaBNfT1viI/j
Y9TPDktARhiT2et4oGUvhikUBAg89qBqpzN2YPlvUnp2IDLkBsqZvMuLbWILUGKa
NSwDENXW4Vy/qgCam6epaMaUjbA5IkJ3MrT0IUeYdIhU60lzEs9+SFmvpTrApuvn
ZJFEowGsUtdR3fWWlMZBLcDGX3atmgkOkeEk80FPtDEC74VGdbfpcjRNDHFDFl2q
s/dwcl8WQ79P9c5d7yqmzq8D2sRz8KEJ9i7Nl0C/myLNZ/WOTtQRysmtg+8HnqI7
WS8xAeMlIbPotWr4WGJhazI6J8LXa16aTr0vorgEC8lNT87Xu9lv9TuYic3kJ3gq
4AW8zEJKX4MGypi7YusDtwInVqM793cXOOdndy2brF3ZvYHpCJZWtfsS6p3vEtUR
aDtGrQYNtq5B1SiSS/vfWbuxuHXUIl2hxreRu7hCixo1g8YistKeiag7e8/Zf7pX
XAm8RUiJMZG7hZ29qlK2iena9TIswIZsC+hI7MFIvVCN51QmmEAc7G4od4uuiCek
EZu3t+HMK7h9IjzGbcz0Wc2vGdeXMqbCsthwtq83xYMsde8VMc3IEpVw/rcA9GNt
YER+KifNx8aWby5bOE8ViVvHhkRXIt9ORNrc558vg7g/zv60A/rUqCl61ei83ZBZ
vGwejgCwyDSTeQS7ZlfhuQ8GXG4UmemVR95AyfICdElcJxIgGK/S3/TVqG13f+ax
vnwZnE/9z4XrPhkVvX+3WA45K4CrKtEYKcdV884gBQpqY5pCu/+UZyapk1jkt+Ba
F33mBlwbj6jvCKzLs0O4urZ3QFYAo0kWTi4jfqTfb/egd1VXFnatllbasXJMvXbY
cuAaTk93kkekjd+uCZFE/3PCy40ZJmo2+q5D84Ie4uj0P/tUvnA6yUlOSPn5QlBx
4TuY60fzQ8Twaw2vu8YkExKQv+1RXiYyU8IoFWd7f8keAO6Z1KOTIdYlfJuo1ZWE
4hADrWgp3mxaZJhutNZnJ+4lFOLgJRQYZPOFkniKNtDitJRqfG39ybXd2R/zqE3V
oJWs7nW5vumAPCWu4JZY9IzKxKCXnT3i5VZccUza26gZVKATiiGK38DqfDAbDL0g
sEGxwwbgxz7p2HSNVCtzF4HIfGpvkJrgBzSf5SPBFEhG4o+KzRA6QtZl9ut+M1JL
IpcLYz619e4XPE/6WoY8V0voIYjTH7G2nrogo0PoMZe7BvP69GcDdG8dv8j2xTLf
FeJ7dEwnCdzF0n+L2YHzQsimGHB2+AUI9X6qAC0Yr1PRv34oegqnR1i0SJVUOKav
/2sf+MIuLROi4tr26vmWF+8EjtiIXZWd005OvcIoW0E4m+mUa1uLEqu1Z13krfxe
Q6hppw0Gf2/WpafTuRpBtTEhrs7lXbJH+r+LM3NKdwrz93mObQLntzus2zCmY8ms
AKS/J+R+vR9Uqu0+iuJPO9u7Xo2W3o1//XxO0W9iq7VHGyiPzIoTKbT6Af/zi2yl
9eDoZUEBUnaWDaJXPni+FLfEGDa6paZfUzOZdSJv0mgCe0Bx64y455woY+THaW1U
6UdTuyWYMpoUniO7SHYCJ7WE18Qe/le5YP53tMIOdmoRMZrp4E/hjcBQNGL+ckDm
r1PjdvtyXaE4Nfa2eqhQ3AGHDUIeUPQaSOYh3aIsMIFGSsNcvWzdagXWUxhVKJMv
l71OlfRdMIV4LXJNzs2FAfFIVH0SquRDR95FcuQnq2z24FZcIEvDHY5IlEO915rb
/3l59oDHXItfZjQEoctGfRwwh/xiVxqdM82C55uVM+hM0Ob2uq8CABIoCrk/9Ag8
i606ZWq3/V451b4dses2NwqyOKEuM8fyaU7HQNtP7DEb1u4LrJEPdkox7ZGBCb6i
Q4tI7bb8gTTONo0uQq9CrvJfiGMfyx0o6l0Woyy3Mea3btXEaT7FWoXCQezgDKZu
n8DcSfbFp4Ua/bCWcclzyzx/pxnjq+mD6/XkQ8/aHidC/DfW5B871g4oAiTHPQhz
e99y4XZ2/oHhL+sOYfSh/u5ar2ySYJH/GUu4AbdkRolKT5hpQU4DoswEysrXPCKI
qN22N8I6/cgVuK8BGtsSl1G6PeUmgFoQwSe+WGUYrTOIG7dT3dhJ1dKsPfpTIa/m
qev7xGWym6waFbd4SH5lesOnPIcSOr/xr8uULQEsbrJsMZ4vkPhUMHhlm2iVOcDG
gCDyuNV+mP2Kw7E/wqDrDXlpQ/LGptouwRb3mbogDX8nuIWgvHyopg6Gu2oRXa/2
VPcI0MNPQHZJAzVyJGObLGNvmsg91JLtPaGJWbO806LsnzaAOiQQIiuLGTzJ6qSo
18n2E594yFY01HYbeQd1V1P3OgicFF5Cy1pSCMqYhQgwDR4u5mRfcJqp3BZNdP4Q
PuItJr35lAYpUV6ubzKsa6sG6nwk2jPnisuIRXTW8YJVP057lQozPj/A97lyosXv
4e2z5aMoTJWPPRjKn0ajuA5Gu/s2nzQdQEB6iRIiVQnQylvTaotYOhi5rRBWrqI4
zrGAb6NZpKhn29PKp5Twquh/VOEQWsBq/akE/+TnjP4+1jQvkWpQOICRAKd4KQO/
xTjCZ2S2Sbny9nAb22j9ExAKCXpO6BlNkFTf8COinRoJv0YRUngv1A1enn7U3AP3
gXGKSru85t4OLDBgUQ9jb3dXx5X+rOWSASAEGtaH8fc0Pi3FEuFW/tV3qscmsAaF
2GwdqIGnvUDsRoLe+pOJCAYLwmBlaENCvnhUOv3fKGl0Lv1ezQAM6m1Oy37N7K0j
QK/iP+K1awbd/vP7AVir9B5/JVgY9XMZWuRLWjICfxj4w/8pydq/trNv77kMSA/e
n4+XIjebXZAAzyxSOIlsbIODVkRbTB23viprCsWOgULqBnvlg/MC8Gnw3K8grA7w
Rhi6ixvztIJoSG9Y9VUZaKEf0vWTSlY0WYXhsCrzD/5ijmRfacCCUDvHqyfjJX96
sWxJMwelGBtb+FFVjxRusXDQ+TLwKs4EKpqdGanmI0i9sgLfBgGNcRYAs+SeyMnQ
Yj/QhwkbbDWASMWSZA70/Xj0HGyDsPdaAnxg32eRBGD0eEUqDLg/0uLGC+RIJlLS
ZqAIrwpYlOKIhZK099tkALwbhPRgZWu8tvOzlY/5aEgGc2KvGsM6ehAQTytTdYSD
XNr3YsN+pASIhiXnNajIzeEF3f9HvHaGP2mVTWmNFKb7a3iwQggHaqD0zg6QS9ct
TE3ebQcofx/zF6dYVD8YZGEoeBLPRp4vafVhx9hIalhqD9HnP+wv9nUp6mEWs/tV
9YHoupvU5tZ5BPi3uta1EZvOHSXs3fTJEspaCSsZ/O6lok6keyjkW7XG6KR4Q7KV
8dbsx3kAOq1bQG5ItNTYBXAF/56Ky6yjbsgV1kVKOowMYphII3FkBW7j+FMLFbPB
Rt0xGBYBjoS1ZoudhTsiQKJunJMhzFnDu0dqymgth8RpAPyWuNyeYwmnWkVhyVlT
dpNVoE6FN4snyTJaXZaz/HOvfc6ek75cLHUQ8rnATMRTZQAprO8vqvG1TSeHQG5+
XXmtVHXcVdqbjFEu9jLQ0q/62y8A4RHObj1vOaa4G4JS2Gb7lTBLp0xjzuSMlARr
q+zJ0Y2j0CEXkcJsbU+DrY+tXYFdQQnE0CGT01vMTk1IIM60luhwAyyCeL2J4hRa
xKZVZcHQvDvYuZn9fkUlP4aXco4oQw9Ogsis+G4mQSHUMWNRFpj79CZW9LST0KD8
XHYLnAFvtBS5A9gdQKzg6hsHUoTJMM7IhIZxdyoBpJ/qEGTLVXbV6ciRPv1o7QPs
Pu4bQrKFVLIa0o0h/YJ5Q4RYj1d60duDu17l9WeCR2aq+T2+t5V5EuDBXxrFDmdm
I+PDYMfkeRhtH5TAzjlPJbADbrSInSoWYzfAKGgmXPbnB4/W+gJChSn7hWy0wcN1
2Sqd/laIuIuo5X3pzaAVCQCFC9UY/TemW/NFgZzoeG6jvJZ+XN618evt8TffmIwT
eJUkN3MgCKMNGSwahQWV55iSKydJq/Ek5EMj4qgRUVViL2NhKqedVHkn/kTS7mZQ
FPbJlBnXjwU8Ji9MHOUPPFEQ04/xue0vRnsifLwadP6g0xnwlQyxj0//P8MvRH0z
ZuAO4Rt+uSV5rBhEOxjP3mcCgDyOUSedzrN5nKtUYEqYC+g4pq1zkrxl2qY1+8VX
3TA+BXxt8RKBveHrdfR/RsWEjFIJ5niZFJCtc3r2NBjfTWl/xl4RYsXgqTNVW99F
FDOPUhofRE/EBZJO7VRC+vkZbyX25FebvzQIt4OsqA5luuk+s5zPfIe+fdSachxZ
gYINLKy/fSihVFxpS5QVYZioh0YYKVqasbJ4KWOi9kZop4kNfGBbf1z68xepFBju
qILtbWjbm5BjGhBUspZkpMZYy3RwUAJPatJzY9ErJJEfI6bE6OFhxP7y2g0aVIe7
WPjUGtNKiXVxk37UI1HnP6IziKc0CDr2+1uWy5ZooHrYb+PyWR5r7+sZuVyjj/Hj
8Ej+CWmQDo5AgwOFrfjkFKRjU85zQDOWpU+cjAD8i/Bq2sznnt40IiFYvEDlKY8B
fdVSJKIGBlJyLg0xbMIKdK7dD+SGGQpuxU2chvKFtbsgj2qXETOmSgMvPsv6vdk/
R31Fl8ckKU0WVHTuQnHP9RuKsnGOc4RJGxHFgdfEoTMlzLAPKVv3JWSPcoQjd/3f
N+V92kDpxPeJwkAxqOwbxWUP9XkGd21xL+QR2Xazu3B41VDEk6IMcy3a3bICRpcp
/+jUj7wxTEa3kWTqRrQZGeUSALmFz2/bmy4duKSIuXJX4j6H8WpfR5g9wPveAbUO
bbGNS6/UE4SlQuStMVSaJTCqqkpHgA9wXcEhRpu64K1cuLfuAhXNv6xcjvEHBW/Y
fbd5feCUNWe+kL0Z3xID7Ii/7rKU3JyIkvHfNKy5Mty4AaqL563Uc5gwzvmTLxZG
3JjGbiqV/0GnvL24/hyly2s2lQ8rJ8MrfT/L3W53hdwMrthPd9hDEO//D3s8+zF+
/zx242mqLuF3PIrshoVYELKdPTuewFSjC/XEJI8X6zHCuXeyRIw3V/wPXnX9IIEK
ke6HKLeIuH9Tylw9Yawk7wklkpGHinq7ELFTZ4d+Q69uBHzUPDAjioD2VuQI0E9u
exhORUiMGjQ8lnkONIx+j3RSS8Hy8BcUQ8EqIUJWulaaVmU5ra04OHYwHRYwfrh6
tNTvU+m6cN2wr2JkAJi8cXcy7L7wynRNnlUqR34+C0q1aQqbOdaJVMs73yfiC3TU
NFMo/DmFKZuv7H1zutPkkoTr16DppaEoIWMfUhOWR7qHDF4DcrusnC1aCcBdNYUN
BXoqUuE7Ra2OzecdrXN0i3QgsxkBxujIxGrljlS6T8nWcOXOUB6y57bZKM8h3rqx
LRiYMYZJrn5v9bdnmO7PepSOL55FtE5rP2KOtAn6mH1YCnTNKa8YtnH4IBcMylp2
C5bjY/7P/EkjasDMyklZDO6HOdJvFifth5iPejPuEDYFMA8zNUTuTskGV0xnokTG
nT8oUAfX+Rz3RMTAGRIsW77PMhqlssG9KBZJWf0QP2hiKBI/cMYLBy2099STjKEh
KzI31agSvt/5s/ZXxbmVdMcKmWIUd1Z0kUeT9UeT6c7V4nE7TI4+T798R65iIYFB
QMwVga5KL2dp1UJMO3kezrZ5GBzGbLb+18BLrVs1uQzJIJS12I3m0trcTq8T7V7k
j0xsCmd0KlKorvw2joEV4zT3AqWpQAcCpdZWe8MG8e+I+aPHHZYBw02W9IRouyIw
BiQ1kS3LXsDBYNMZKrGwyi9VChrDwH2mNFc4gUuKHEwY9GkmpOmXvE2HJpMEFlsk
yrQFuafB7MZryUAWUgCYUF7h7Cp1yna8CjGBnQAnko9HgcAAIFAIA6lX7Dl0knBP
8Ui2dbqITYoBrMRZVhUhxUH15vm8Kmel4fPi0VZQO+1pelCsx8gLYZUTJN2w1Bax
Wl7Sb0v1wDB2+isekxCmtBcetk8L7hsYa+eGRFVGbredc1aAUYqrKjGy9KNgPWtE
eZA14hyKf3zQw6r+DkKrxZL+JvheMPFLSO5NmE7KQPItKmu/VA5/GFlb8VlyPMWl
VhGFzTRUhDqm469cMEMV8DPTp4A4ofi0q7r7gTpl/5H9WswS3z/1hSYwYLCicYIW
twsglFsfLRFznvrDzyXYm8pma3iLjj2TZewIZobdYKXR7AtzOBCLJ3lOY6U0fjve
XQeA+mPyei6gR6ZjzRlNnJ1GwMQ6w2WHSvQ+uZwU+NnNcUEOnH+NmGUA7nceTFfa
nfpfbTpz7uIMZPKOtbkd2IddVHCJNXk9rRyEz4ybBq+z4piCRzYy9O0tPa6zJUgp
SHzO92v0l2ai+yvrEQVKnTvW2VKN7dLkCi4Y3ehvajgaasekzLxrZs/BBQCIw5We
aYySwjI8OyNrcTHeMqikmaQ9vZE2EcD7Apu1XtruD8N/6By9yifC9v2m2XRK38W3
MyyadZjUGjAQYTPrfSS9r5ZyG+PsghUD+H3u/zdStUVwBMN/X0PlcuJe/vGNFUZw
daWk3jkZT/aslhqsJ+k5kYd3NkczcggqjoABOck5jN4LuS92llF/31RVrcgxtnTI
aEeEY/eglY1Bch2mWpfZ9T4YtKOCFR3z7OXZZm113oiViRVQFE/tVNo56CIfJRT1
BCOdtMZHTnAV62Os7fL+tLglEZNgmIaEZN4YJ3QPgRY9GJ6AX9BArsbR0WN8D2Bb
Rd62aSd0kIMGImuMa5fMi9q2k1P0r7uEr2FcPSnaELoiXV3Mh+OZdvXYNhtjpwYk
nJD38mFnUrAozuyw/upHAujQfXDNbjIi4PjyImb48FaD2J+udlux7U3UmamJbKVr
sTP4AVVSRUTrv9y+LvXpa18Svtj5ff1de/dFo4mC0PF6za23UwFC/JXFhRBjhIFJ
04FqQs9sdjjIf/F2GrKEAaPhzo4C4z8cc01mP4aeY8WofM1G0mvvIPIz1FBdRJ2M
NIuo2QMJfNS7KLnDZN7R48NC5q3ePyY7dEdmWgdLmou9E37PVueTCRMa1i0viyeF
bE4re0arXuvqS9zGMxy/k6HBkxZQvMgwbubDAnIli7RmOtbE7WLjJFIEKrccSJys
Vp+Lwk6txHnthExXfcnB7Axt9OffdT4gejPFe3WstQVuOtBwyAtP4soKn7oJ4ShV
x/ug8q1IPK37JVm4L0jdSTsb8DJVkcvTD9qCOIR2zu/vgP1RhyJH9evTU09OrqJM
ESEXFHD/x8JbGQQj18rwHVhrDbW07ZIB6WgkekbOp+HMSGgVUyGKzus0yZfdEL21
F68spGXbLSMbY8PQijkro/k1Ln8Jx3Mcf1EjR85Jut4Tm25s3ce25kfw/EccsNcm
Mw7IYuFrBD4rLwB3EBOJT0lQMC3x/mQ6I1T96KDwLCnXhPYBrI3pBW7I9W/Hv0ZE
P/R6gSc9waZnL6iEKU8clhUgEQ66udUNhnefhuzOQXb/4oy16mafrRe8yU1I151I
lUXm64vYhY/acQ3kYqFsWsDJ6UK9x6QH4mVv1EYiumdx7jHVZKw5ABLcm+ra/F5p
UpFlIsqZBBgQZ2R/aTejC1uO57n1rLWSIILxMYiRb+NYCSaDWJv+cKrQeJRtjWFh
91CkjGdcwlQpRDxTPqr7qXZEKvun/FqssQJVsDGsawpu5WBoXLBgO4OGWx2p08AZ
DO1gTUUpNYwJqPiRg4vhntqJHl+Lz2K87qlWLg3w5c3OMEEvMGIz5RRKQkUn8CB9
R13S+aieEUq7xe+cPIP3blivUryF3fv65CohcgpijLEmk50dEpiIjAkQVG+C5ORz
vqg98UQaKmTq8zNA5yc9bYPiWLqaisT647Cqm5+ijBXgm6Kz9BNdh7Ym0EFNyTVt
2EPYr6RaWt1rFQbl9Ydw2ZuC8U0xRk8fEdRCIi5fkh7S7fzZXPI1JWEKArKIRzL7
otbTzX/Ncd1C2LiR3tPFnv5zI+U+VHuF1nMhgrye6xZP/x13uzM1KcLD9CD5lp33
ge6cK6egiPmBNSR4LRLCYEekoPkry6G0uIYcxbx6cSLbMwMsy2m9Q1xe8V7KTmpU
IwVsV+c8q7umVaeIfFHy7OFOrtXXKwp5CqHpa9pzX4bjGhv8Lkz/q/Baw1rjmlmc
/myHi0d/7pOGtbIFI2HtiOZbHG+yPOP3RLdWR/8GOipoaTU2XYtHE+BmcSi9uVOi
NYyM7Y7Peg8URWpoCSWdWzMxDfcLr4ZiOKLJLE98VDrjExX3T64v/hCUdc2rhXo6
PCUyAeUUsdqKy/uwscffgsxgc2zFb5mDfkBtihfE5IJrEjhbwFWtJrYfHz5E04Rc
vo+lhzIZiFz1QN451aNDfBkSqMnMsMIxk+NHfE6F9+DZTHBth9meUUI5TdN1kBAb
PhFpe6A4NL+9DA3EXVuDLuRMKZ0DwGtk052jljLggL03mRGOlej7B+a/h23Ofb0N
CiBK61V6yCW9HSZ+FHkKnsODqek52hao8QG+PRNF5gfFGzkQYLsMeHF36zC2/FsR
SK5lmXADC86iJYOD6QB2BQZMamPKfWnvhEqEvDFv9gtYesTS8WsGz+XjRzJgFytj
DW6kNHjS88gDiNgRAPQrAQzNJYmJwfC0SCWiFU4mZOHoAUVGpTPC2kKry+p9oHVd
H2kSHVQQpJ1PDh8/T0aSj/+M0oeoKTIAijT1SfrphWha0a8UZSm6Jk86iPLvLY22
u1CGOtX6UWVdXlkT7vP3hbCngNRD4GJJetmsKzwb7GmMOcdzouwc9hZoG7312kj7
Laomj7kBEVuj7Sgnz+EpvKjUopTd1jIMyLgwsfSRd6PM+nfEFDg4UjuRk0J61r8Y
wQqAHqM/vcaeX7NArjOz0ZMXWRkV5vVYq+5mHe6paeCIK/dl+pdjnUxuu1rLdwzY
NzEzeu+DgIbXxoWdZkBxcV7hANCCPJ2M8aFeBIVEJZx0d/geYnlmRPL8yG8olfWk
gUZ44YRfzwv9olgjK43+gidhyZYSjO0RoTJpshgwugQ7IztV1zvrMQbC8vHXixp2
HuAa51eq1OGw2cdpDCexGSkwUrUKfCQ+EmRnDHAvknH3hYzAQWZ00Mk1O4/fPeyY
NJaVMFPiJ+vxwg19wrjnSMH5Z49K4Sz8dMPXJoubUSQ59LmJt/GrMGXPpSIef6vR
UcaKLKRmmG+aWD5RtQ6uEYHCaIZ4PgY2eYWdoHvsTcdJMNvprLrXdJ0x9XEqL3ro
lpzJbfdsbxCu06MNXnwebpRFuCzrx6kz2N9B6U+c2FNNemNyPl2KvvkOTdViNJ6a
c3JpmVa25PJTyy9hWEqH1ueOlcOlIXy6J/OArtFxdljXqmM6kgSLYNWDDfxDz9Wx
cCOW8JAsOh1vIN6KprgkehPMm338S7KlmAdJ9NtFgeTvrzQTntsOhZ7q44Z/nOns
YINlQ+GC/B7GKyVjYczGfa0wZrEa21JEAdsTSWj3YpL/pbSW3L5DjQgsWdebPTKk
zRvBzdYv64pXa6VtAelJp8cSvMC9V8rTDdzQEUa7x4GAWJpFp8Asj0gwO7VVYPN4
EZ6Tk+JsQ8+Z/U4Rz6xI+b+nJJFqqOusnN9LGTzyUaMdLEc6Bnh9ZOgfqwmU7YKz
BfoN1w0Ze2nwNlBj17xBGIpXadeODmet8lfXFu5KSgdyXJ5Fwj/ys3I6LtVigPC1
+n6ksCdIWeBm/paxS183ITStLw6+S/qOZPXqy19pwok5htpyO9SxZmIEgBuVRWFC
21bxowJx3oVy1jbRr1YYGYRTlgpV9QsTyhXKCtsZK895giowrefu8tMmZGZ6dan5
tr/Z7DOg1emvB06y6/rH+ioL/LeV3tJOweK8+QzExCgKBGEjpPjhVG+OAJ1Y9IMa
mTTBxrFyeOiBXnBEHQ40TZXhFGnBdSwteDLl0DAzTEFNpVJVwyVPbswMD/OFUi5x
pbggIYbP8V/gzhGxg+XAjxT45+yvVeyhEE7yNGk0ntE3/wG4a/nTz6iXuPmvfkhc
xFE8XIp1F8YeC0lBjZ9CCVszzDry/3lZluqMgo2oyK3U735EA5v0qTekIKS9sY7m
UCOiI3f8HBxZ0Rfu+XExsCoZOUS0QieUwKmUTRuQMZX0yy2uIKQZ9qT+nqCSVak0
FMXliHrIN1fOH74RgtUnM42c+x0fE00v2GGZWsacj66bEVGVJL+IaLSOpnW2ao3m
AAdraOCEigzeXlqRePm6Y2E74sZuSb5fbhQux1xZGQyWZyoMsjjkmXuEHLrTojso
FdutUwsRf+42K/xqdWQaJkplCeLVdZXJa0chuLaR27ItFY+Dhw3qqmPMb4WWz2qe
7bMwQsWyjNGEM68coNZISP2IEthSh23S3Ako3Pr6kYpvfZA4ZsPm4p+/7awG0r49
HZEwP8oFN2noP77+q6xHGTwLYVdwfBOsVnTSLMxQaD9QAFp6l1oIJ4CCAC9JemwS
M58NMn9O/OeeWvL6uTKTKzlhwk45Yy2v0e39ijIG+/upaBPtyhvf5HqSeKs9HFVN
vQRaejE6085tSWNYH0FcOGmuwV/4El5KyPz6XyMTe3+6tdCrQeLijQsSTYMNQqmG
2HkzqTzY/vHyVNj+cFMiAuiVSRt/GE14rC07gECY7ij9ekYMoP1Hsf89yXZ2t0x1
EvcSn5kFYXjtOfNC3BEngY8q01kZgmrylT2Qnv0W3mq7KOE14VOGYe+hKdvfxDF2
imkDHgs/6g2AtpPLwBJzyAnhfNlRKbkLwLDo8nDk52iRUsMW0dBIjgwyZM9POfWP
8kCIt+Uj1qd7nEjRle7Sud51RS1QjdMLVA85TeU8F/h6bBvKlW6opgGVUysNYXLx
XBU7SEbOYDdoOp1jNgIYYG3rONHzckv6xuqW8KkKfId8CRsSQap2w/XOR9+WQe97
zlv1BDGZQhz5aXGen4HVoEkbKdJkFro/z3/KovFFVzxzOyTEFlUsFLyglDqR1HDN
mx7qn21QEjpeG2kyC2tpplLAbJd8e2+H5MmMQhK3DJc8QOravqfPjuIL2ttALPAB
3+KhzHOI34qrjl5Ep8i1r58yiOSPDE1N3plIvM19DorgIcXfDVwFa5LopIzKdHkH
3zfHyvS2q+YiQmov2sOokrx41V82hMi/1HskSbBZc/KLcbZrXe2+SooT/l0ROZE2
HGCp2O+2O5g66/4MtBjnifxM5svA/vnxKCBZHSzt+A9HPE0bOcYZTzfQ5TkctuzO
Kje8f7p5fhHYeGWEnk9fmNZR7qr35VKEAA/Ro6Bq0P5fr2yk9T8Vb7IgrcoF9EpP
GREIlwmLCEnJHrVBlDGUYBktAw/lpMsCmNzpVUxFvdGumD8N5bjdjgS0BpBcJKAt
B7J+8C9ekioNN0z7zFqMuzZjvC+LlcaVGaDx8ed6m60W4CKZKCy0A57azcq+E2cZ
80YNy96T2Etw0DIQIHZ/YBSg/iGl6y1VrmgAmXJgIyGEN8JXqzTD+eU5PaiJMCyu
2DkR4527wnowuinbPPBmpwhyq2EH/L2QTissCYAG8LEk4za4ehoRwJJWO0MoQvdv
vbzo4d62cchNPwjOdLygyxiI9A9u8p9eRUN69EBV+pPFhZkUZY9oBM7XrFkm4uVY
se7UPzVfudvvLgqeGDEpatjvrcy/mB6UAwWF9LlRxmMYM2XiNUTbO6hVgcLvXaOC
TF5ENofBnDX5HkQ3TMSbhxeSYff1xY4uyzfYIYErAI7Pi5dapRmY851/xlkU+ws/
OX1d4cAeb9qnr70ReojXFTx06eaGII7n4KXYPuCz5GQAZXgzWyEJ+TT3cMNpol68
3RRguBwkBIx6e0QDrAVtYumUnIZpDCjBZlrLSWtlfgqkbwjHutTNGqWTeYsiqQ9k
N9NlR5KUEOGpmr3Tq+PKXxSJiw5rX3Nfj4CUdfOqT4ZWge0nZ27QBvnqa3YQyreS
KLl9kABteNachLip5AuGqEezJKoDMjB2w646Cfh04G/qngcIQbOGxA73SHIUABD1
/IUIs5BZJW3MVGrgjJKFi4JmdDJ2pNCMUFmRBa4m4e+CdaNezcBVeRvmbR6Zodzk
+uQIPxHMqjM0lU1Wmo1+Nt3kq+s0iez2tUSzPsS4Gh3LxFoPokzJ2nX9P3bOHMtB
7n+aZiZR//yG5nYvexYLSNxCPjLLutG/QOE24icul/NUsz+s51zG/7bJsnAc79o3
1FiF7uxNJIuL5Gcm/LrV4+pj0ZyE8GPfU5cELgSO8NOkMwTQc2rd64omEVk/9DC3
QJh9phHj28glv1tR97Os+9tQFGJfgplq5KjfeWJJHNP04UhRMNsq8j73fJ68OqH2
ADg2ELCcnHfPbGsTu7HwGZ0kEG23kHadXkErpVdRbrdPtteAQikVA6xpnz80RH4I
1CnbF4zY2ZMf5jBBHLmv4C1rUpYVcaK8CeQjqzIDCbeG4cCFT+QLH54oh/5jXuJU
4g649shrJQk6nwr1kzrcm2RsrObbOjJbWa4l5OU3qm4oN0RPVStggpZRuE7k1c8O
eGVWxmsdv39HvhjTRKPPGmkqHA3xNISsNPcwylxLNP4y+R0h1DtsiMt0GCvl+yco
sfAy19jK9LKaVUZkjQXzoSr6UsdH7DFNPVZCb/EnpLdgvGfphd9WrkQnjrwwOGBr
oMUHB0tJ+rNWeO5VfUrQqWYBJCyEAe87rNQ6wm/5vK/0895jA0FIR3UxR53CqUfC
QD6eeFaTXchPKS4AP8mMFrWnrD+s7B2lru32XrEcfJx5T2WxB3ddWzB1Rg34m1i8
azdlq29V+FmN9lD1wBw9ybqIYoFe4ZW4BCxV4HZXgmmacdeg6sjrZKC/arAAGlIj
6YzDaXvEX5WxPIvIwEStmau1PqQWTDsh7yh2nc8ioF6uTecAZtDKT64cy6ZZ2Wzz
1aRVVN2NpPBPYtLuvJsQCSWU1nxGJ6Kn/eUVwZgFtGITt5AS5/l5hnoGqPaFrJ7j
Le9/hmKeuaFv6J/kDSTHfkhMmlXiDzV7lYRrMogTVFacIidPCgbQQbX5t5KWHtyT
nAQhSnl1Rc4XDZF3X0PSboSE0csaWQ9g1vZKYs2hQxzEO7p7+9emDRo3c0Rykag1
9kPbYNfQlcXUQgrUKS/3Omc5seVd1rg5ZT2H6q41XfsK4xuzQlL8CG/bHmnWZ+Ml
473O7CzY67QM2XmpL5RWhKL7QUjMCjAbo3ybjsJJctdS96so+H1rVWsKnaRtw2LW
owyVW0esNzXhFX4rLGZVKWH7Tijz4YXmId5bO3ePOCEDCfkzp+VJ9Bq8g9XQNQTR
Dk5oVH3EgYMVPXKHN0OoPPnTRZwYgIIKp4jsQWEm5liCvQYOq3iB/iuTEWE3S461
art5xKn3e3ipSkmdzL1zX3+4xFb1PjwXetkxOPkLU3VO1NA3zjZ0Jfq70TvWwIbP
wh/DwfL5MpZNNbbfc3RIZGiQmQ873Hfl+HFPEWe78ZH6FuU+pAHHRst34/I5TdLf
mVEvQsXXtyQ4vjoEao+vfARrQLCXnCZB9v0HA/hYYuM/HLu33QdiZCZvHYwXBBGA
+IZXlwlwzJYM4Q2vi3ippKbgD5fZiW7+lE8I+lLKVEO0/0NyIRCbc3Y5f/gxPamP
STXRAefbyxXl86CSzUWcCJc/zVHbyfCC4SxCGOzXUTV9xTfY/HOIobM9W8dQ4jXc
XJTZL/2ci24ifuRNaWeL1oByNABSEuYVQdbp2wig4rGA8hnS0on8eA+dNAWD7TOA
ULsj7zaqobxdhv80TGSwuMJrz8nAS4JAYdoRQKwJ5yzdUbD7sUdr02PpZEKTJdjp
dyif9Lkm290fVGzPumJaprPM01nkRibecMZhWaP4tueJoACEqP8ggs1le7HpLX2Z
nFJ5ey1VKW+YElkD6ts0Sd4XZew8OERO640nzH2HjezK6sSqA3mP37lhelLxSF2E
Dns1LdTPU8vBl0+0sgU/5ADN4RHVjXO/GeXGjyZrDPCr75awVGAQE6Xf8B81M48z
+vtSxwFneAB7+Y/0t+XclTb0neh+xiGoKjHJqwzQluUukSDjNbM8O6LccTmY1DSq
wJTc2yApZOm24uZ1jgUC7h5C1z/i9qGL61aKSmmYrvSV+RkIMbmDOy2as7nZYl5y
TlD4fd0Hpc/wH9VY8kaALy0Dqdz6jzE4hzKJwTzjcKxJHIaohnN9vufte3bPwCPl
i1OTvktD5OxPo0IiMLg3dp1bkFfr43s31eSwKTzxKVq3vvwO1iLwZadGEeP5hoWy
QPlRF0TzpCKIyiqcZNdOeWe2+nAqdGJBY/vfFvccFdI+mU4BxPLxwkUV6GpeRXDU
IIwHGYwg54l/FMSIKjZfLQi8vvL350gaQacQ46FHyvXtbYu1A+QQN+zkwom59Uat
8oG85L8CQA5U8GmcF8t8Ai5JT1zZFrJ3PgnPomWAYDYPDPwb9Axfw0PU72PLNezZ
E32LdbFigDanLaf7xJ7fCKC/gfGQZSQ/TW/X2mUo+vOF2MLoysmNPyP64pWmL6E7
IaOinx6tRM60ePqPu5bKiKFnoLW78DmgaOlQDdTLF55nkQvAC2HJy9+vSysuLflc
1iXPtxVjsvE0l0ngMWLWKX8RKynlIzkW/4U5/okO4WcuiYlgUi0y4chKBfN/03a2
zBrjcePXXyq6OJPpKvWbXMVsR5shD2tPBEOEO4Y7+ZT/ZtjioKRMV/Nws12w96E5
14y8s3MDZgPJYGHL7zVbD8Hj4J8HPTmP4QTnXTJ2BeimkgA1UcD25+grKvbM7YDY
HzXm70NVqe0lOSO+8Rei/TNIEJfAw5HEvPykg0ZtgT/x7Sba2Qa+M2JolxfmCmcZ
fRr9E4mnaE+JIGu9JAxsv1DPVQ0sevJGp8f7ebwlCd1DG2W1hwPNXi85EcgDcMnB
D7EhzVvWZm0mb0z8HqHfeZXqSqjpu6QXkIHk5ZEfCX/OphELCMCXZkTAmoiHtbwJ
XP5wz3k+CV56q+JQysQMCAh+lv++Oz+iI1GZn4Hcej4+FGyFRFDYo14eARRfjtMW
RgoMSmzIlZtdbf0XcJWwkiD3yF0Uy8miV5EpwOXReD4hKoyPrd0o5tYAs5N28hM3
p3sJVHeN3XmZsnFk/UFk41tHVlxSvDYlQdARzXgYulWOvKEFtaOuTHa/NqfC0w8h
hHc6rs43M+HBic8xCViw7MgqIHZ/o6yORuGr+p3H1X83Mr0AdJmlRApfACGVIEIY
Qb+Qqo6vVy/SwG3/gmcxJFKX+qAe4AIYWQtAf8nK1eIqyIVXKR13gSRYFRAgn7Hd
NIdCQLAQ+UpPgK1O2Bkjgi08GRsnNAfqbB+fbm/yiht5Z+/Ot+PIxq1vwHpAcWVE
XfwyrHK46231wl71a7f7x2dnprl8C9rahNhL9SpIavGKblOxlDTz6McAgAaDckLE
Vz7k9vGBknjVvLneHRlIOn2ZaG9V4w2XAlejjowE0BLRCYQGrTDWVRMeLAU4ypH2
XgIlmU+PK+1WLy/61uQwyU8Nsywem3ODR9+LX1+Ch1fJJHr04mYsfBUpiVdt/aUl
Qs7lbb3x1ikUmh5gtaGGCwGq4tfQZUngYGD2qCLNmWzVpHvLG8NIsbl3JAY9OQJY
Y84HIJuBOzxPG4wp+hoTOcG3kX2oYoT4Qxe8dkJzhmoYMJKgeiza3Kr4pEwCnUMr
cZDBEmIrhzDPFyuUfb4vb0jC8BQUuBvF87dG5mUQLCutK5W4SVlnk+uqfmIUHfb7
3Ml7yvm4lyvkAzx5eYBPwu1Ds9V2idxuD02n+aVktZUBUfFOFjt0XZB8/Lg+8SEB
nbXbuTgHgpfxlbWRigbpMTM1GGp6EpNnIVg8OcXdoa2fSDiT/Ah1xoG8IvQhCYzx
MRxDsC769UFPggOuT5OgqOtATPKD7VLsKWrG+aQdk+27VyGuQZ27wCwwT8oArZ3C
QLkPRI2OZxcHZK4/GCWcN4tws/B+C6Vtnp7i9SjsY075b82dJGeUot7Cc8DnVEz7
JWaRdL2v7ItW2j/77zXmdJjVm4oCepz9uYt7zC8bSudPkXGflqKqd4CSBU6KP82E
s6VIuL9cOdnGHWmo4BhK0y7q0MXf7vqzJ6Mk0dgfWhBG6Zad35Qe/Ti+8J/9K1ck
MfU2dljnQK7j1EZMcei518M8Z0xXUSO5gakOrmF8RvzSK6fd5XBoIfuVIQ7TCvl2
NF9M7O1RdKOLumiiQDSAb6orEwOXp9uOAta+2oFkZuXqYsxJBseSMBQBn4/Wf0xX
2KYQGmWJS4UnySAh58vws7T6r2Kmpdp8NIARJgSLOemRFI72YFk+O0CJxOV1UCDV
rmBi+yDcwRMdZSbO1Jdv+URwQweN+1ZVI/t+9sOkFHNXkpKlTqin73bsxnQo2a6c
fsJQUBihmi9TNyPoNBePmdRJ0YdrWUge9F+1dDbvdNCwKzhvG8ZPJO0MVA9yIlKk
Kj4/UCqrjU8ezxkSLW1e8dFx4D26nJGmt+JsGNl4D/JKY5hKWteuGBtzFLDIyV8k
cgMnct6NnKNSAnFX7yA0h43xnY/UnWzjW1kxQL1e6z5JblikJ2/nqPcanbSaPT7u
ew8axzgXKLjS/KiDTyjHV6E0PN7y5p3dYLvg1TbbPH+TRfKuTRMuGsriGD9Qxvoi
+Qt/vtZ24RNZtC+sVyMUmkqM5soR7fwgrzwgP4w2hghN88xLzOoozqAr1sU9URsp
tHPHuYsQ4XrYsAzNGh8UEVl79xD0kQSa6KSFmzBkL9XFRES1inReF02jj+51O0rp
HTMAZhI9Kg/FPzl9+zMODWxoUlWryDHOJRItJc6XKQrblu+JokCdRq+6KBly7HR5
4Wy8vhozLgBs8/LDayTDbIIO7F3aaQ2AfrDRlbrPYzFxQ6RB4gpbMvkAr51p/OgC
pvln7pVbgVe6HTn88Fgg4SWmAMxMmn/VNTr40JlTgXmaCkaQRKA3paLYvzxIhyA3
Ob4ufhDzw/mfsG1Zh/vcR6kQXiLdeGp36Gxs3LjG0frZpmPA2u3R3PtGebwG+yjm
uvGlzDK2gA7AAk+ySwL2EjqGxyLo2GnDw/d1XkJQ0Oj6eDzgzmpRENttlqFI1YwM
z8HGs74ILBt/acMjZ/7OXMuC9wsQ4zPL9chIdF9+qJ/X1uJMBvBIGScnePN5j9/g
7p6qQGhmdV6ltzf4poEnWuckixjd+x5aKWSg6880VAky6D6r4PrKlQwb/f1a3Tr/
eclZFuCbrqxJZAiccmV1lIZHY+lfnQA4jmYBcIVBfvtOWgGvVrG+ilBY0xFeQz4a
4shpYBTCGktHLIeA/Ea+9ZAfjIsVcWY0pvUtnK8/k46NHT1BN7Wxl5TtMb0x5aXX
8DKWR97IM8uYxOC3jzx9cdfyffI5PGTJ/r2OGvUDDiH/Ho2lWX/7WLEyZfhVRiFk
ks952k2e/CLuFu0u4uQk+p3hjHdK+UouunblkHhORe3v9xaqBmSbtTaclG0Z0WWy
Km3nS5eRYELBzNpxH8ew0q6BQmn5BHq5E2HapW2V3FYHBIVnT+QFbe8zJrLySxhw
G0s9mSDbbymprO4qsAx98BBUgfdrBxiMq9xS34AZhSgdyPk5Rvmuanix1qPcsBEd
8CjLV9tKFwuosnaa+gBhr/rgO4rkvQqG4OfteZC5Rkt2sbhM8bJYwzTstAZQd6G8
cRp074KRvgdbsgL+7UCPWowINcDUmKTFWnf8bVI8l3RyaUx2QMADhtABjjFssxJ/
04OY3a1JkAMYoTqRkrVXEmLKft9OzWbtleJJJY2XJk/U3hsM+JCv6s989mnxZthY
L+sK+Bmj+qreWDQHP9BXxoVkj8dg+KTypzJVOyL9IQOAoSvnMz4Rb5lhk3VptfHN
ZaGIh5V8vpmilTod5sDlKq8tTsZYaa0NYL+u6kEDTIT4IrQEGou4sX4FVj3d+MI8
DrBTJGTUPSeNx2TsYPZfYDH06NrzmM3a5bijZwp9oBJIqyHi1IDx5gD5Ds9cSpfD
OGBROIEf6U4O1JF8HQueBuzPg11/PAEzweXK/kUE+6/ZSMY8FB0+BzDszs3AexAY
qWPQZw3otB7MgzaRezJSTpG49REpyR+wQ9jeMPzDBtobGdgejWwEeZCvhrPz09S7
5KomzkyJgV2mEmlSblYGNT6dSqCDg9OHWh3nlE66m9ZmBodQI+YCSX9aktRPubey
AHD5/iRkPJTbuEKTspAySpM7PGIoUXfDBPqMFQpx7BFa8o8t3qSj3tmejMKt0Uac
Wq97tagu0lk2JGOV+JB6WnmOBVE8Mhpjwj2hzehRDRIxPwjcPt7+4XlTf6Vt0pKb
MGwO0CxBudGhiIGRTNJmcmiQwWM4lBQwRDRRQvzBFh883ThcyNKVekpaTT9ZceTB
xUA/OulGZFomk8zQtFefE41MI2D2/szvmYVLMkcqeJZjD5jnDPJG47CwCr6OHTGr
+fsn0yGt30j48oJWTW8TdhK1z20rKtlNEwGm8yGy1YCddeg848cQUht1eMfJqhX5
ZwDU3G+8PZXEKbhFwexgcRzlLZt+kFLH3oHaBiMgvRSMr6reSyCB2T1RW8Y3xAvG
j+LLSdn/OqP8BKC6jxgcy7GjhZUSaj/NTtD2i69JuqfslCRbSFabfDuI5o99/7nO
UvwVRAl+MefUxLupltdh3Zd8WV14XydrrMNJr3/+jfp6SfYHC04kOpccRP0jBCW5
3o6/LtBNe+Tu+aJGbUcyW0Duo7fv6AQUx3QQOxGzisjfFLqI4CRvM5tHkskqM8M3
Cp2yXjiKXsNEvNdP//TLc7JxlbDiBdGmKc/2/HKMsBxwPPbrnwVxsHTY+yVmD/XV
HVbzpLBPUsRH80grzsv+bi3+dk0wE9vVYo4E1a1haVjTErlBg39E99FRGsTY8mpT
dSuOYQh0gqL6WnGIupFpVwDd5teJi4ywa6nHKyksur6rL/rU+2OqZpQBmf4X9p4w
syuIkY/nlZhQlIv2MlLeDQHLUSHWdY+kZXaYk9NdzYRfzlW6BLz3sSuzrh3UiJlm
gm8CGSI3ev6GETSM8O069KEwRjKhOOSJBgwOn8Ovdmx74jCKDMz33BCJ7ykO61RN
Lx/H+l62++EyYe7lafnWSbc08cng0qFcT+OQiCXVhyudxe4alU73HwCLpRfTdynf
4KZYYQUni1zisPVGNggJ0KOyA2KHvAEtZngSV66XNhDWl7wDC4KF2ZeiK7vyPNJ6
n3193+CbYCEHVtYKFK4txs4gyOfThw8zo04jI7fWcVt2n0RtFxDwVvTqb3eXinvF
LhW7jD2Ocy/RNNDZEgNRuK4uMVo/b/Gpv/78gMFPkaAnJlgD7xNpa8YercarODzQ
oGhRzDTtjBv4TJwnAwfiwlsoZPUgMy0qpEC/9MRxCqSfeH0kuFTbOxWnNlTwYR9H
BCNqLeJhJ6ydnP9n0xb7z0tl+1MM+DiCj0H0ksEfENI88KXpBmAh9gxDdcnBQupv
INvirrsPJ88SU/rBd+4xI65In9Bim8Z0V1nKdKe3CfMQUslrLV5GB59GOeenzq3e
jegFZ/k5jP2/cUYYrcYKraia9xsjjcmZSf0C1TDqaQ3uJE2m6mhz6+B6gTNhn6zJ
hXf2WdBw51gIet82P/bHE3g4/83EXxzt04M96vTusZ+dth+BvVc+Bwuc+rAxRxgA
8fvx+vbczyU7tByqYtsy1OfcsqmiAeDIp2U6Rf8SWxgpaHyZ9lmCm3HY62DR+cXH
7PKzZetX5AgfTQ5lDJm0qPMlxQXl40SUNo+SoLFEeZx/LtFgmk3q6i4QADfn1XVl
zJ0lQC4OhbhAoU68VzkQTCanfnT6eh6dGIyphq0DstrUQqW+zRWzuHGYZpeAX31C
Ya81NxU9s17IPApU0Z7ZDYAzKcyJ6j/irFmd0Fse5HhjF7p1TJk4BJcaIAkfVss8
aBWoV25gNtDnAMM8hIafSzjd8uf959uJAwtmzdyavAlP9xoQEe/D3k+duX0T/8JQ
YS/9YFPNDkTh9gw9ahtMBo5VBW8Gb9HsmQVsjuuRnCw4UcNTBcUkvY7fs9k/5WVH
S27zpjX18sP/ZiO3zb42UjkSL6/xJ74Zd3STHsrroJBar4cBRvKtygvuRF/rTcZI
6w9mi77J0LuXtoMdvBvkiQ6ZexNpaXU1auwc8uyKPjI0/4BFmW34EtdaYSEDW8Aw
15bvRX3StGbMqtqNi+AHLHHuPp+eULwx+XjJrjgEhzXK6JpmwUSSnpqmggOjSr90
J2bdrghBfG97Iwpb+/HhDoPuYCcM5W7t/UCRHdCwz3cv8lmSIlLLtt8ib7yIhWB6
DkDj68RZUGrGoUF1Hqt1EEcpcA6xTciOA1CoX79xnEmONedOdgap92RRy7TXqU0Y
ZUvnlZDmNoEXDGbXURg/MYVgqj3LwF5ykJQOEykVXTvijMhsfzXsfpWVjld8sV//
Q7/gnY41gQdxbyS7s9aKa2NXy4xDXvWVkAJYYK6wOBdRnmM1TBTpGJDsVTrBof2e
ArWJMaSAPhEkipWf8MUexi/UFSgSPwDDebSbCbXAtyq9ZiUPNJoGedoSyd7wMYJd
DA+Sb+DLpLRu9p89wA34Iq/G5La0Dg9CXYjhn2KKV67IjcikRMEUeoWZLWgPTk70
gtLGxQIIAKE/WbVNURCCIX+ryBM2Z8RYpIfaE6uphL405mWY6QS7NIJ/THQfqa7O
0P/pBmE1vjH1lZ52dzUzJw2MIfLtaheW9nTQNhwe1UXR6TN6NSAViV77Y5i8YVKC
lE7pnzc/YvxQQ/3Zn2tqC3cE2thFkpI/FXapnzcTJfpy6WTMdMiohfs8uTvCYJM4
IXjTCRP/ZirCMXLNjV0UvQC4WslBOJH2Qr8881lSLIjUZVxUYq1XUipNDpkxYaRI
LA5DtM5ycQQ4JhzQpI6N6hbFknGxG7jg6QVz+fFdmYayn2kjAcIr9+LJ7Px7cmFH
cYqL1SjsPGZTH9TWjkWBPhjKT2AJigS38w0czwmlx2NkK9aNuAPf75g2i29jv9zm
kklK8nkBVXQEYiURjMVmw1OuAmkPT7XXLqFtNtGYpsvuMsQj0xf9wUn3A1cqLw+1
S0LPEqMI3PM/fYQKHtcpJyFfUfyAVEwhe8p1tGHs+2vnVyLEN6C9UZUokLZi0RTa
/4phZMPCRZUDz9xL4l4ZAnAutdrr8/6LMI4FPLTca+Z702fLhC5QOuC/o5rKsgKA
k7aeG4H3l2pAUrg36GBAGlYeG2n6marHkw+0qUsc14vATR6BFJ+XOPq5M9vuGeQT
WEAik9ZJNpEFb/vdYKx89PgjjGtJWEGZsgKgzpDt7YhQx13iePpL6yjrl2noWk8W
YeZKvD07ClduVOjyzftY3d9i+MUdZ84yvEoQOWIgbvmuBpi1zUz7XjgdHw79qWfH
biurFoY+jkfE0C8WpKk7HSZTz2Glicw3P/7Xo3hZzFbgweIGNWWhDWC0Y9K64Xzr
KSN2lA02yJx1SxHuhjZxrMpmyGLg9n3FsfI4SvmiabQ8BeOmeWQs6ROD76A9X+Ao
Z94x2DzA3BCoLThrOQMg32pOSKYN8rqdUBHrVG/MCpDFsxQ4BZNqdPP60yfMdLZr
8NE3EHcoOF6APczNDj4Zq0daFR/Hf4BgsiNCNtomJB5LCNcl7aFodntDIY2gXB3T
pWygxBKgxtqB+3nMv1R9vvFKaBntNPA/AkIA79jjITI9QIp+catau8bPnbGpwlg0
OHL2sBEpIML23m2qVVrWuPrSBRJ7H8b2CYVn/9eA5SaOVvuIHvsXIHGgZmcKovOT
vOt8ymhtnlrqzvR+A115v7RVtMPLWBJC4ZevxVYZF/0lWBFseSgENzOL6GbvUMez
JUw4Vje0WP3baOwozHbyo6xweenIPF+5vrcfGJO6u8NgiAcMurHEfHpuG0KlGmSB
/Xnw4K2hDXn/VRESEOkZ0ks3h/y/6FiZdaA/oZalfQDu8eAyQoPnGUi8q3luiucd
8BlC71tkNMzWr6ayj3WKPk9yrtTIDLoSnkBCNOf5AW5rDumXia++tZdQpFhM4r3x
z75UH1sqrAn4WEjZOq7norRwoqG0YDrKDLeLY37hARh6f1/E6Ar4Iab8MfMcYZbe
y5Xnp9Wb/RQY7l4oNpSZ974BVr46co0OSULkmEIWME8uNA13zVDr6//uykamKB1G
R/jOs5IQV1PQfM6xEWLDM7tvHckw7A1ogGQ0n4Z90zdm2AOL5erNgvvNh6yOzJaK
g5K7/RRQPPUL7W0mTYCjX48ArKyOaFhLCIQAdtfYlIUTKkZA+Hbts0bxyOhWkra4
bhjDq2SSl2fkujGCW+mPwkpobchYt9eyW/WXcJ/9MtYYUJ9BY45TzKVkvb2z66ZG
HZSbGExbizKorV3qoQ4+WfYj1ST7N9zMk+pNjcXhGqr5urL8XX31Qq5M/x5OmqdP
cF2SLIYQVIPyA0GxeqQPSY5+k32XCOmcZdixQD4EF4/4ZY7PVI4H3RSwOoGyVoZL
FRi1+TpVafNB7676QsCcuYyCMtBfiU2rTcGvmIRfKoc1/UAhVdm7z66liJDxLyYo
neg+qfWSKbCsaE7Tb83aOHz3+euN2JmWg9XxgppvNu0MMIo+jS4SjwYFQE6YX/qs
eGInjktKykEnC6Ne/Spj6JFekMSnN3CvtECwsXT6UWILumMk81ibzrqSGirPa8cB
IAVMcgvPCuMTk5ApOqteeKB277y8jO4uWFarcogixSZNszpjAYzPs/Bgoi1jvcs4
gS5lZX8B6Y8tu6MVK23FNA6yMH5BALKJ0zhFXqPfsM0GtEKcVurlOJD+6i+YZSc1
uEao8hQWVtfUMgNP0NQg+fq1OP0HRZcNhEYEVz8LcxYP2dLYXfaRhmDf564WGofo
WLwsXlwFNqEp2fVmGqbl7dKqFy3xh3Bgn/26JVcq3hWKOd/6vsF8Qg88ZAECbcgP
GuEU0GyuAcVvZMomBrlE2bq+2Z0rGCC8kHdqhJMJbVeXQ3hfBJTknl1CEffrYQY1
DnfFadd3vDkKG2h6k6/03ZFlkWpQp/4jDuXaOLeyEObi20RsD06hvUgf5sKL7WTo
hkyvLehdVTPSNVCf3HAvMLd4AKl5DzcxyX9hogdLfhUBeU7n67QMxrFRzPO3pnDO
qQfoE9Ede0iosjZqTpIICyTWHfW1zk6RhaM+9T1ZB3iAebBLj4JLWAOV8ylgR5HF
j83/IqwCM0RWBEr5vjY9hkhwE9qavV8o/FiKQE9d6p65tiEzX/gCfSNKYsoRBtny
3uesy94diDGTNIA7QXU+ie3lTVEft5KrdK5tLg6rKtL7BRR/4ypbIytGkLFdWjtz
p+Qlaq0uh3wq3HfIp/K+6hMiOCFXDuQ8fJfbXEOb4ZCse1aluOQmfSfE2e50zU6C
ROq5H2V2QHXbC0gMbq11Ukog2ZsMV4EYd9KIsq5bVQPigvuKTjN8f7UOI+STtfE+
p5TmbIAV8THKW9UjW+jHiZCHCPKNHyvtwDNbExVOI2xuDEOFZN09KhT8/C9kY7X0
q+EM8XRywTrid5SlOIMUi5C6GadrlnMgiF8/aUYcgLy5nAsS5Zb2E24gR5A7axFM
4fw08RzJ/uZBzQ/7rUi/Q/tC+cozajDR8FsCdu6anNBy/FuZs/FYg3dRKT8wTn44
jywxIXKGnQE+gUQ0xiZMgs2jGI6Zjmm7ku3Rcw+YWfAK3clTEcr6gDszHpCXHEiy
KzASQQFgIiNKCftsKia+VpdSH27/cYzhFlpG87yvFnuTMJYlmeMq/K5SbopSYTNd
7qccpTbSEFJc6fIfGleR/D2/tG3Y4LDlTH6gn+PGNjA/Pu0zAF815TA7riR3JZvT
qhHJJZdsw7s3l9J3qubSAjnJVrsVeSfbdoiVZxB82g9oAWwzQaH6FU3wxqx26qC9
89v2ufue84K5BtMSs4jS98Hd+Iy+jHtWlE/QeYHzziqNukzzK8JimDj59Ei6pTH+
rMBy6e1hb00H67TxwDc+uKJ1huwrRjmCLJfKAshWpzmESWkiEu9VWPr6wjDkFSqX
+/cAekD/gLctfZD3f8BzasJw2f1L3GhB4B6M3XFHmTo/v8mRpdVtIgGa4m0ZCrBb
xzYjiyqXspRYK7fA0PERasCObltH3awGWuvEvv11rUnqMRisHyT4GmoaiA7TgmK4
aRG2Vk0FZW2iIaF1Bp95O3KNDntS1x41P8+ZnO2lNlC9eBeTIipUrd7Y6xPUBb7H
75Om61YVgwz/uwoAiGpocSCacU2FvKwuG1wW4HRiUCLi1qmOCpKAbf6TYHuKhPFH
jV6hvb50oDadkAS1/RPWLJv0NOAkSASQS/Auv8QNK/+kee41ppwMZU14tlFLGnAt
xIMV00o0Z7OCMXaEMbBpUYNIwARa+7aGGZFrkxZ/h12qC+ZaZbBH7PeB6Y31k7Mz
G2cAmEyibEjWk1D85tgiuc8bUnsuTX6aDDFh/02UgI1KRij4tLTF91GTu9BSAgwP
6zV8ZDsA3GFaeTbaW66GbBe+haEzvGt0guIjK8LKilw9k4JrhwIZGpqjP86FFXxW
NK3m6PsjZuMEKKDF9gjMGTMRszI+4IlV/e6ZB+AgzmVzhEnG1IwgAglxM8dxF/nJ
1+3q/iQFHHtx7XYCEpX6BXH9kDBHgZf92ovY720vw/k7JedGWFuEiDVkxFOs1Zgq
NJjmq07jdidPb6rOnyYnh0tSuP2Rj9umDJLOxDdfOdLdl+DiCDheHagpD1OfDT1B
98MP9jtAT64lU/VU/AIoWtzcD0k7JHlUQ9IwIEcFPvx4i31033YWwmli2MKq3QSa
BS1vCiONi75up3HcqCum8oMTEMreATryDMZY1kVJgFH9tNt65Ta6upPVf20zwbIq
EEvKy6qMRpZeR21YnweVScdD6jxB1TeiE5ruP+0Ea14t9YqLiCHJ75wMxYuf/NtR
si6UkFl+3BPbvjjuAplbV+vx4uwaCt9CzFAdHY0LbJ8m41OtnfR/ATKWZlCEuLNc
l8ML2uN6cm3dLvUTaAwH+vkDEv3NiBLtishJSAJfToOq1hWLFV/Fafs4Hq7DARRX
w+1jwE01pWtwQ867IZgP2rZWET9X02d9p7xKV3NGJ2BKduoXZyetPI/4yaBLTCEz
tsPFaQFZFDrexUweReQPDQgdsD77qR8WxWR/pVhkhr51jyViexDUJRx65szS9eTS
rKRgFx+/CX/kL8IxvrVZHZ0Ud8wHiDfIm70s23wC5IrD+240irATJ1NPJReEFxwX
vEogG9RWM1lgKuTPQe6a7ydXMwKRAXATAs9lAC2ua/j3uvSuuPwxY9tTcGSiYbFe
x/7VAXKYyQdHJbDgyl3cP5ZjmqJcIGmjCWOYqpv6c1dRn/e/47kkDYvFqnMrNNPy
ilBKnIjHb3uvyTFrUZOn41agqpGZXZ0mEYzTr5H1ljza/D3X6ECX2SteAkC/OJQ6
l2Y1MsRf+he1tRUFURvhRdh3vFiF8Q7bl+wv/VoobJioEgPElwx/RaWX9XZ29q3w
CmFiSAw1khwSv6urut3iqPsZwWRHYWAFPidyWhSbmIzDL/+Y2Myo61VIlNloLUqH
3zYBlnQu6YKHH3pwRStdqY2b8Qdv1KIJPU5pfgD1zcodpguCr55oFpkcTGUWMRTb
M0EIYQNrrfirCVEgLx3cVds4nWGjpld4viaPwIP3MNivsm9a6t9AEV81OT99H9kR
GWKTWTAhwGz37gYvo+8ji7K98dtkuECoyLXCubDX7B6TYaALimC2dnCreHGgvud/
TJJ9kQWyk7F2Vq+DgEzO36KpjPGnEm2iDJFc6d3hn7f93CKESCdlcN8FnNwA02+P
WlM6XSZ4lPZCKNdAMrTX1qvGrVJ2qJJelSMunFNhVE2+vi58jPs5FzN1K+fv0xQu
flgGAV8uhMluZS08X1gX4r1nEFEMftp6ropQxhS5XZMyr5owr4me6H2NG71HpRqw
RNAfAqT5+w2jx+cyNqRpWQokwTQELPOTpuWLNTvLjr2ZgENWkEsZ51MUk8diUTM4
2HvC3nATzPrazVg/jltPA4X/x/K63KO02xc0t56As1kiYfeJ+62IPuXK6ZBkwfct
3skxt+dZpiPxOvwBUxGnK7BYI5VN8P9sjXk0NCLhT1ONBrHF6MBM7SY6BwyorSzI
22njbM2Gtpa3kemJQb9mfsLcppx/E9ZTzL8XEpeGwYYTEPs5rq6Afxu4cf6rqTNT
txwzhuzsfTVW37J6Rip33udwGXHjMR9mBoizEOL6O6yThENoAuiKwG2ccEC3Qt3D
8pZPXTT1cgp/X1BWhEd7IX3WPmSD7xKG5nkQWr9e2Xb0fEsf50TT6o9/qnJluDAv
FClxiCL/ETNrIY9y4/IhK7JOLzavFD2ehvPu/uLZTw35yspa6nms2E/MqzDMFZ7Z
ZdzQCaJpbdK18m2pTDRzl4BDpLtnQ7IkRv231uz3YeM83VEODzuNEZ9iwlYaAoTW
DCLFhS472DB4r/PvTKYqB4CL3sdQgaFPz9vGZv5WYorKKrrNGtF/eztDo7XoqBJq
qTNSadFkjjDXQs5v+c17G8MBIcJkh+prz7iqgzlqdXeEbyumSIwrE+0onwZRXYl8
ibeJdnPTQEBeT8eiQJLbv57MFfDWqkYtrIKd1Rpwj4NvcgGcTV7DgZAhMvirQlvv
LGpW3I/rph222zLTAgswy1RkHwHVx7n2nA+rwS06MCkcdY1tQivPIvBHz5vEEeFH
ZNZFPKVwq0EmxbjXkkKoVKsTUYhgCWwqce/OH1jYaOfTCrAqN8tO2zmRKGrLdQOb
qs13KyiEMQg/unF0k3FRh+Axty3LArWawvVzjZsYarXpa9+PmZkZKnpnQG0y8ct9
CXZPbJy5RqaePzmN7n5uofeQl+xwUOdpYRfK9q570rRsMKGQ8eGUBRhPFQ6YGz6o
A2C+ejAFrbpI4ME8YGiT8Lyka2ftff80vBuSzsJlLNWxKWsxFqa4aQ3yUzLJPrVT
jefJMQbnmauUFVrT0EuPSeWp0kuY/CCsna++OhMJ2KfM4/UbZXInD0u7O4BF5mnL
4/VFznXqY2I+E99/RVnUK2G+Q0YO+lJLQs0W0dMZC8gQzZEAZ3tpHEELcOz7+ujn
chr42j21baMilF38/iJEUXwjT4cS4q2HIO+NQ0eS6H1ORWfTFUk/3Q8NLull2+95
VIXmG9U6n1bpCtdWBF4I61cBDe2nqMoDefQ0/nAR39w9eZITjrQLC7UxQjTGtvG8
kVA/JFNjTIZb5CbKeieCXxPIe/P8OMrnl4z57dne9E2AMA/JHtpHOm5bccnB0n/D
hpooKna6XJd60QdCIlJYwIpgTh5gLIqcnoRvgRHD9VedaP2O7nkR96RWRHuxMFtD
bAWYpQjmUiPZP2CiDLopaiotqwf7gmXxyBaf2pRyv6qsd4a3rZ+ZTdX/zPXFF8w2
pju/GXbCwbZxK5e0MxPoJIyWGsrgvkW2GZZQoN3kp51a0NFNO2JERytW17TUEfXU
0oANKiyBDn3fe3dEhX1Re/f4Hbo0cEQiAYkO1xW1Ml4Z/7ehXCOUzwB3KaFzz393
ixwyx2CqBOF/ntlm05dWcTxJrTYGBKHuJQPl+bLvAwRB/MB6Sqqihi4I8OJozdOG
zPk1YzAZMhWXD225xyDlK3y0aD/u/iNVrHpC7BIq3Fc8fpB8+z8NYvFOxLqQH7hG
dpTk0AFtFeO8PjIZ+p2im3Pt3GDZ362p6YRtsWcl2DeZzxVBGG/zPoeaT7iDu4Di
9VUcEAY3fhZlBdrB7tYCVEOY0lfgt7avWWkxoOFZDPkxx4d8tt3p85qW1hhRkb/q
t0ZKrBeYvMtwyd05r89fWPxQM9c9bec6bX/xZb+22kmw6j4hyIvNlWQc8jEy7CoO
jH4pwFOH5TrJaifFh6tpYh0hMipmDyAm42LVZFeskwhGmQULA+NOfy0Vdo1du6hu
L5ely9jZRWQftRK8wlXb1hLh5F+Elq67iYZYPy7IEKpUuPDN1VEeD4njCb/Kn68z
GvTjNG1duclyVl1i6SM/WYxbavwUcHkjlS9T86jGr3YRVcXGTdmKSUusXHxgXFHJ
Ga7z28v8t9TRoG2XInNHBltwZ7Vq3T6kN86teXAGNB5/TrGog43rdOXeLf2n9yIy
6hbDvoS/AbYf3lYmOXBJo95LQxqpiqNvCNIpLYBOJV2nJ+fSrKU9RK0GWjBeMb9p
YukbzktwbiURyVLl1VSm6k0MxxeF+h9vBOIdTQE3Gokkng2yw2/kqTWeQDZuxwEv
syCgB6zTk+LekvNzKf/OO2Uf/O7fxdZ31SYYNgzkJUh6GCKTBmbJW2TpZtZNRgXo
3VQqBn0i4ca0C5i/t6eZciBRF+0eJrVjPrv1tmyRMTnS4Wb6SZZbnDZ4j2rpiBqf
0MlatIHho+tAcLh73EZOlXG2A2WFUIP1yRKLD6H0lw27ezlpwY/6nfkitgr8gMRE
TW90uyNkOraoEqpuz7ctnvEqLlNscbymsZGYfHfrOkhnsnDz+7JDDF4fL4/7jcRJ
6o82eImJPv17/tuA3hwJ4v3Cx84c146/b+wl43SLtI1tXTirR6/Tv6aGxopyZbto
4oEajVkijvDoLz4L//lXEbVseQPchiqjNw0zAlBs3wj6VsqJolXT2QdgKG8OHnt+
NCoAsrTp0KQbAnxTza7xA63oggdAiULBgqESOfEHwqVWqSrRnGituPehEcHCJ3Nu
jWvMlwSCSiOGVG3hRETahwV0YqpY3r15aE61AAzCp0/Wltrnsj7cKYp5AbQbVwbk
ed01wMxpcBYbCSz0xr/e+28ECZfPgtTXRaZ9jZhH/p3GcuLtjZUvCY0EsR/3fEvk
AybNSLq/7yqbyAh9xERxDkbSE4ZjmONSZY4khEMwYFkAVYAEPQKCEfSNov0niWWJ
+pbDg4dkLwnlGKjKL09PwX1M2VPN43jV5rEflsA5SmxmzzTh6R7SXhP3/odm5Y9T
ZbgkrLuLcdma6qXlrq0GP5f4xNw+IKUau4c2Dk35Ogde7zzBCFH3+M4UgVAT4Fxf
XNsnI8e+TIjsGiz5MwnZyN4TlpD1crPKJXvUHZltYAyL8NpyZ5fzNPW7I65fmjAi
052C8eX9Yph2eWY9z0kfdYjmmp87oN2l9SS+FfmytEPIMrPf0VsvL7NbyBY93TzR
IOiXvr+kN2BrxH8IO7jGBdWcTyvYmLeDQrOHecmPY1rHqajcE63UqujHnuCL06xv
0rt4ujgtjzVOBAIZvI7hohKaNtBG/SFTEWO1dHUrw21ANrKeRYSxDaRRlnjg0Gpj
ZM6AB55xdFUQvSS8YFo4QYp3WTmaqoJUzBLqHBDiXqk+nIAPE3ZGxAydoJbe4ZQP
4pKviFnvg1ruHqFz/66FEqda9h5vEZwYZuPmODX5IOXEcSZQ23iGX+VqiETArZQ/
BZuzg5642mcuJhNYGCvon9R16EUOxTKVtiSJORLQh+wFsy+Z4wwMgfV45cc2JILV
oBavefb2uVT+izR/Lw4SfnLoKYP8BNyfPAkbMl05LEDrc9EYtabeQ5ycOs4EON1O
2MtmueYKANmUufQF4NAmy0Qabu5G7apYHDSnWNmVcxaFVB/UAJmBG/IrH1CRAWed
wH6m04OqXBRk1djm8C7cqDRTe08yZ7GygbVp0pm0ojBkg+5U4iNja85n+IRXtG01
D72PrHS206FJGrCQ7dufxjvtL+6iKTQYin8ZxGa4REhZnUY9aQbo3auMfaGS4CLS
QpmEySqAzIlkrFgdl/EBOSjEBtHPwJo+QZkOeiE157YR7pH5HK74jKhGKOXlbj8a
tWMrvZ0BiDOjEek2MbfE9gPQQHZh57ViRlyZInb4oWrh/4MOhnqK9PiBvqRDqa4T
vYJJ67fzSY7enOxoMS0ntWgY7z9JHZ2jiQEQgRUR4c1YfyGhNnrQqDx4dFZkcVf4
6XjwUFI0SeycU8KboXvgwh7LKbOwLCdtMO5/MtQOXql7IWiWY+3nBoz4or2IITwl
owQF8NgGCuUZye7qApBN0PTybJI2/O9KhXJARrZsrGJnvRgZ47KXNxPkeVm3uiqc
ak80/R5JqmHEnJ/yqXgZhJQaHy1L3zT3/3E690z+hU2gP8Oy+hX456ayPS+6zTsw
KyPic3sv7kLyksSlDKQwE1X9YQpe2o6SCWKly1oMkFZlG8nIFt69HYTiV8iN/vBT
Lg3krYnCyMUiIJAp0ekWBF7r61s6I9GrlMOAiIOXmWNkLTRXAlqcbW+WsMqOKpAb
EjfYpwuZtndnXAaLp9dWsxYD2Uh7rQ8hAGCetgJE0yZ0BXu7lQal/MBOMuFqWS6U
6bGOHlqH5OV74egkKd+/Ay0voFTHDX5fLITqgLapl2N+MaLdB0X5JAKxZht86YNe
cdkVis/3NitUcUwwHFfw+Ar09tFRVK5AYY15TgnB9Eva20C6DuJKswAZ7b6MExzC
Q7YBQGdf10DQB+v1cs3GlSeKijQ8xJrf2msyjd+nklWQxiSx729dmhBYupo9lhzx
uNYuGXbFnAIF1Bs50mQRqVHQU2W4Okne4LbE0lZ56EmEyTS5UjdUMVfvKXciRtZg
eQG4dIrKeX0dt/U5aT6mOM63UYDPcHkdVcIUPTiWgPAhT+3fgP0LXR5HKa6tPEDT
JmQIK/sTRghzSa8d/sBxX7XX/ONduaS6BYeIqNxC9tfI9H6K6TDw5ywhO/66yv8u
gNT+L7kqdKSIQLNUyt1ngHqb8tWguJaDeqKa51dDb3tu1GI238vkh8jd0r+z5EW0
vkv8+LYtv1VKcSv2Vl2CJJIOHF37tjJVaac1trFkQV+eXN3qBrVis0Gf3Wj1klBB
wCuppj6cZXB97WV08Fw4qhQWp3ONOWyQt21mYB5qim66DqPJ2d5EmJgM5xYXiPwL
LJNoTx5gGiRrOGkevyDsy0J+RFNIGh3/tff0CwKXRIsCmHQD3gywhLKb/a5GwjYC
wsLpQSkuamhBRM54Nqq9JJZcl6SOus0xnfLHrA42v0Lf1zN/Z0PTGjbe5HDpjf1j
1tn92UyUCCTwuCf7iqAUP13Xl3iEn8iciEppYv5qVcqTOeA3dK4FDDNvKE5XnZFv
Umi/DOATYs959zrfYfvK6xMakDF+Gj5cFvXrDsZUvZJf/ibYZXt7kskcvFfosI5L
fPtDmyPgFFf5dyTrAH/99zuSDgZyHpksCJYZ+fczrVqHKC2nw6b8zGeb6lsdqz2+
Feesc7/8JB8bH6i92A0THexDk1msZW6HDsKRrLULRz8Vdds2FgQ1vKy5YjGW0Kyd
Sqo/cqocD2hwBHrmWSqSWpxpqhQc3oE5dK/4yQC9xY/9YXPnxNmaSAgND/4yBrWU
TmNP2qFwbZZuwL4VW+wZB2Ti89JKI24U7xZP7QhLy6DLhTUr6JLf/ZjTB22Qt9i8
nFL5iKQOHvhzDGO8qs6OqGUjeC8XvLbLn2ZqEeb5//qLSBYxY9y0UWyHJI33tkwf
KFEbspLHlAvXMqrXsylEpM7y/rBPcDFjmqKDwYJSJvSmtCnVvXAwo/nOYTiJEa8t
1nonfGYq1jAD/rFSMtu+gUqOPZmM016BBL62y/m33w7pSE4YQdw73cXNsrWo+7CC
/r2spFgtSbjXAm+jozA5dmbxT8Fg0ziPQRytcoSVmj3Ifa1MeTehzKgW1GwiLuv3
L/haSlTYo1VSBN3tMJKaOzATGqxGRTk7YLuhCdxXSxXXymUSXo4YJG5VX3kP66H/
H4wTtPACPnxHPOnYfWM0fta8Tt/dOf0Sp0Wnh9Lz2XQnhY/C08NHhkzPW82DmNYP
ilVOztoJQtg2OEZ+jq5B+AgRs44xt+rvyrjhey1PYk5y16qzkT+4n5RE18Gooxrk
hKicCETgm0vIxszaf1AqsYqQzymsMafJp21eTofX38M8V9ThSgdPbH4mD5fLIx3B
B8jtOqoMsGiVvci99G7z5p3aC34/o2ssyMriQ4lapebMoidGbdwSgvSHqZ2GR0jo
2+JnQzNAV9c3HKwzySPIhKZXu8HbjrW361rA7Vr0ibqMFPz1J0Mnkbe5C4U5+BQD
QteC4/qvo9MA7mdQwX4hDq1g0iWSNkoODpf///xh/Ab5KIsUcr4H9YjOLOEiPerU
635esD0M1ulv4TKkhS2WKONJFGuq2+GTWiZcI+4HL/3SwK5BedwKHmvhNfyMIxQl
hwdC90876JunhVF4bY8gpvyjoSIzSlLZb87iHfC7Z++K1K1y/IBGBjH7HbvczYhO
Z9C+9HucfzS44HLVjXFYUxNZTNVwpCNGEHo4509LywQWuPEjI9ZY300X4zETZlEk
2/I9+OAoZZh95zeairzZpxnd+ctXbrnLmkqCdlaHvC2mrF739i0V0iwDAdjYycUK
e7s2TTl7R+Y16lUgyDuiBxWqcRb3CwLiTu0Iip4XGROTEC5Mz4zGr9fVKG0qdOe/
Sk36ZWrSeMkI4q7PS8mJlj2shr5tR+1tc0HgxSSmbCbN/b+Ht/SHoyMo6aeHSeSo
O6XMRQV1TPL/WNn1iOO9GIt8zrCFok8t7ofIfOc0lju/DDykGDondLamd4kQiIy1
WrAqlhq4MPfE6I2fmv0MPqhNXmyC6/PNR3L+gj2OH2atW//edTK/z4u5BtTtOLT3
vLKsKVgosJnoe4ST+TQycqeBPKLfsciE1hLKeVVH6H7sLYXkOI/Lu2Uu9yQVf6v/
IKztETn/UsrR/eVkiQ9YlHgeRoV1FarTVEnbt0loGY/SptIU2oSrxQgA6CM01yj+
p/xYEeF5/57ck48MnqgwztxeHs1EMJZ7Zi+yPLGaPPkXZ36oeLUtq/vgoXL52O7i
zjl26KkjRXSRACICilE7vjRWIIJz4JqIYfvpnXsNbO/P4uj89R2CAi7swUiZxa3C
24Xh219HyVAyQNFgWrexQWLtT3VO8E80eisrXjHVm7pBwTaLajTuvE7EQmg6Apcu
w6uVeRqnEJRkbM3qa8Z+6EZjPy8DQpR/kEkpz3C7QMuzFKJLJFpM9jqeF+Xg2sX8
mLJLHGDvYVsaDAi/pzezXBywaPrIb+sKCzy08rE5F8XmnAmo5WsIniEkNCSAfIR0
EDq85H2Q+XFFKUy1VzZ6ai8P160KiTErl3NBYI227b1qtBgRCgoVy/JwpazFbJzL
m9lwJJi262BHr7+OJhZ56JydA6KDNOsh9tzDIdr4IOkFW2kYhyAtoIcCNVMxK6M0
uA2CdXOvLpNpSADRa53FLv7gVa9jixA6EWud5knb4kViArMbSk8CDOCL0FvJVA3h
KXgZ3PJRULVTMLLWI4Sot+zekYOav+mlRi0bCFON/KUvChDeL9EW0JRWjbvNFPxa
Rvk318H7dYCKeZaQBfYO+EEjvbW+rTlliVLXevct5K9Vt63HKy7xRFS51NOKDawY
d2/RinyrX8gfd4Ukmme1y46+4IZ13tVqWvrxkAvb+OYBiAfdsUG4z9+WBX4N1N/U
n2cLQ8haX/IE9JWxTjOp+RKktLXhc6A0cJPRtEqlKNRxDz467QMA+TqL4mqQci5v
gD5ZT/JTI5nePBzxPHlEofTdYRWNABGgPoGKdzcU4X3/93Wp0bXeTEcziEMufLTW
5gKEMTtHFUuJitWQurIKnFd3/Dx4VO1ppcDfP3Z+Dy4uJtZmO6UXqVLtPBT15dHr
rtljRFDxyaT4j8oNNjN0r1LLb8/1oU5w1rRItBXsgTXLDl4wT1MvYg6vP1zWb+7R
bLj80VAhFqAZG3L3cMMwVdrtu4Ygijz5s9c2+893KrSKR+o/vl7P7NKjmV38CHJj
fYPS3fB4NhEkD5fRiRRcH2eajHw2PPWRBjQzucWAX/1dmNkHgsC0DRburFoYinnE
lFbdlSR2sSshU6BAICnyJabsUvh++gYiro9nFNMwV8/PtNAvRFQu8BXuvKb8VZWl
dtMVqAo5SoBVYeqCIwTt224CkWVwOR+zLGkSQnBrThsywwHUWKJHkgUib0/xIh2+
bopnlTsP7lIut4umbovWK4H13eXhYIG6FBWEPqTnVmZgHPfG+VGv4ZPRBbaipvpV
wqr5Hp7+4hvu9XxfhSCFe8p8IPIr95wT7xSUtchAERGiuNXqHpv8jA2cScRBQkZ7
W6Dwj3AcFQ6eRpWDe4W4yXcTSLyqDJ5oQVCr3s5JWd1DDoYNeAKvv9pJ1aemhzdo
39Mbtu9+ncvDP01e/LzpDnM5KUn6tTjkagvWYR1yAJ2c4xMWZNqpYzolkWMPhUmH
qope2dpveOmMAol1ETg1bPE5jjYAZvf/4P7Vpg1sgU7rgXfXXbPSzwLFa5Q9Abd0
lXd0NQaF579D/BvzluyBpsNBjjabRhyVCgEq+3cKCeP5ZsIsHvbSAkgXIw/QMQkb
46ACpAX9DFwSbg3EeRs/I6gkeKC5+Hedl/gfncRrF8ehDNnSszesHwvQRH8JI5tS
vXd5ewK9//wBZTUuv8PxNHuPn6pD6ieuIMe6fkb3rFcFKvAGoG37PnFshaVJ+CHh
Ey917PoCYhN7nbASYzL/VlZJYZycYUMbBRr34PXwWOeQpE5sit0Zuyp2lB74ovEv
d+MSqVrpBY1k1mclDRz2GBnliI+lXoaY2MHgO7vcfqpNjkXtkW+F5L2K5zXFUN/I
LamJg3X2fcbNG7X/jKszf+4Zr16c9mEmYF0T9Ix3IV7h7RixBpiN2jCxBegv3mgy
9auPhsUfqL4Z8yjPQVb7sGBGrVG/1ZoGKVXRxeK+nYMa32gLScAwP1B01n8vhuED
05gdsqRyPQB+hCwXwgjYapoH+8vbEvyi24TyE8yh/51eQfMRMYO5qYQokhFu/Ihc
eg0BdJLc8CEl8U83Wjj7KIe01nb7z3qg7a0vNfE948ztyZQNuG3lXU0FBmHwYGdc
QbM3SZi4OfQS70RxN/rTfqQkKfUZDwUlJ4XMSK/D4jzG30iqwUqbY7/ZK9a6nq5d
4ad0lVBremMhmo6H53xrBkUX3dYOBPvWi0O8GzgPSbVTwKODbdOVLbc5u7PIMlpF
keRbgjqUQRXFitck3rkXIjUg77uy2jxOd35Oc0nX+rJwm6Nn2hcrbz/eukRc8Wu+
JcTETuyK5o4XLAwJuXOKxbVQhXPO+98zd4CJCMnaiyQJQJdJQpqa/6/FksUnZkTv
9BIfFR7AxpfLbpE5XYV8+MTkDTNZ/WvY+mzP43aynfQilpE5gWAkASKOoSATAbYt
XcBmwrvqPFR88bqvT/jENle6vCDLvYbPHQF1RLebmXSlmEu1o7NXh1cKvzPXUJFd
UmUPr3x5wGzqxQrGEIpFrnLc9dKwUOfXnMoUVrrO3LY8f2YhVJSM9QQKtw93SCBO
CK6Pd8h1WiXjsyIVVPqHQN5NkVduEpy/sKnU33SkfUJ4FBE3XqkQQS4Yqy1tYHgr
w4zEOsfo1Bj0fCv1TwADpH0dB2oQIIJnP+yedokzL+/EepFcONRZc6oTpapYqYsV
ii88V+cLaYc+x1jKOTzeiUWX9hXN8A75Tta6s8P2aml483JhNXOWy1yzYEQl4j32
cXrtZyoLbBgm4LBu8hTr+yZBN8HCXbEOY2nb1aarLqOHBRyt6/PrpiSV9vRcHSNM
YDcd2I/fLFSXSNDdIThnlKX2rHbn8r6SlGVHHBbJazn1SVP0IZQaH/E31BLQfMo8
zeo1usAtzjO68f/Jm6UIPkPj8L/Wgztbp9Q0lbFYLljbJIYbTNaMRvL5Hj0KH/sX
xVaOzGQM6p6B2G9rqNOmAb33eWkZ1ZZVnWg183Dsal5idIx7CXM7zqAZcBC0l3X/
Cw4nZTJ8zDYx9+WklCnBvxoXOZDKZaMtrZtbuj0dd8ylrZAW9PuD/p/ut3TVl0+7
dP/8S016agS1i5bytznrbSni09qKxrnN3f0FLs5VryUNhcY/Yry8AzE8UgnINipq
l+qjjUivnh52erTTnkkBOyyIXZra3CiJkI1biJd/sUgB3ABXV6cX96PL2c0fiqXw
RcyMIYrLhfzVHs/x60wTDqz2yurKwR7L2thflMq3U7rjY0NO9cxDIZdW2QjZsEmb
YiJv7J59QqxGbDG0JhTpPhuV2s9GQdMZcAeHMBcckUDA2QYALDfHBmMLvciZi8bv
DChJ5Dluj/R7QNPXYjtvjNYBqsppxXnPPeW03MxqGc+05aG/nA3ndUKpv03+9iAr
Q6scLL1ckuyTIBER9cTBhhwZ8Yz9dAY/NAQGtfCCtk6Qvl24+tIsVet4IbaT2knt
RipR1Hda2B5Ik7Bize29oMlx8xmiGTlKGJ244eSm77cTSgI+Hkr1bdvb6NDpGYOy
IiuSYeEOCSpDcib4k+/wV3wCQR0TMVM2KsMTqOjMQnNz9lEW9TJa0Xhu0gls9RxL
IS/Tjx7Ar7l8hhHE1jf1lSkOtcUyBtNF2rh2HHxSilZWmPxbM2R8TukRghh6PE06
QB6FM6gFYSUtZZPpczKTpXPqdBve+xGN7vEGcoEwq9YtDY/fnhkyRBHDvJC50foy
J/k4nEqXMXYCwoLLiyRzSxqUAcAzONTcCZHHo1dAYO1+a3Eqk2AmYPVnWLiVrqA8
Suj3GjvrcaoqAeHHppM3K35TtkjoKLxqYNCR9/1uvGY6BvJo4HHm020gZByb3c77
T+OUDDSQeBQzJdoeP0Qs4k30iSkZWeN3uggfs0U6ouQUY5GuVWPNFtrM7PR9SQIB
cFa47FKo7rkjv8dLYi1/H7nAOi7SOOIcwM+UGi+CCzLQDsVtQEF7OV2DTCk33UUW
3fBivGW7/TxVDPH+VLs963DyhJS1krvyRpa79clFCkbCzBRAENOJ6CpjtPpEsHSr
QDyJh/Zm2uOI8JYCW+qVAhXGp3XCYsSuzXSwuYQM5k3y2z94nLlfRLW9jtc9PFNZ
zQZlw6WaeWa/kEdRl3ngX84xV6SHq2WyZe+8KDubmfLT5JS2Rz1VNEiLu+5YfD6L
e8R9U5BPiLQkzmTaoUDJbS4Qf4prF1z68ChMxh1kc0vnfhRCDpEEYLlOURjvqkcE
gqNhTR2Lx4SxAb5gxL/mHl6tFn0/Ibu8yccbDpjWQveoxw1F81N/pQ0lj9x319Er
TE+Vb4v8yiUR+c/1meE4XV2Qw0jbLNY1DXj626GV+Otv8euyCKNKkErxjFzEUrA9
6484xNATDU8rMfT885i6L/dcCkZ4+QsgjStdDJXWwemT3giogSu2uUP9NVglaXlv
ZHa+uAePM8l6He7UBCTJpkMyN+g3GsjbH2JgWFcKKiqJG8XFAcq/BXvn7grI2OUz
obEBHFHHUgOVpaV/Nuk+667EZia5rK2lbDMpm1O32/JD5B1ZZzL9MZdvki9elbZl
Xw6bkMeUkPLR8J8a6zjoEUeZt3Ci8TLvn1rQ6SXh+f6xMGNLGUYb8sYiPKI+ccy3
Pliu5xmzHz82Jk5mkuvg70VOO91SLvn7mO5EYRNXHFCth8zZj9yjKo7xOgjwdTmm
lWmg48Cz/B7Q3h+60Eq7JI+dzfPUQBuhjAT7tTxYF6A0oWZIvMQ7P/kBb8VX11tl
++3/6wJhP7+IvcbBZdoRtjZL8x3N8Z3TatsTNisxDHS2kYZNF9oYduIpKJDTaztL
S0tgGUDHKCyvQbufPZ+Kpmz8TVZq4dBhM+FJunsp7Nsr4MdOtSy0osUor1kveadw
oxj6y9Rjqwpq2CxZySLXMaDOs8rqUxsIHwnZxrJQiyZq/esYu//1OvIECad34zpc
On5c59qtIwGXi42ljVS9m0s9zR6GNJ4SHkgENH++2wqcqgLhtRJPxtrz11cp5Z61
+tY3YXZ5au4gkppokcxSrkyEVbNww78EcBiwgmwpGSZ0pzOQZcNepy4qhOJuLGxI
jFIvU9lTFgldMox0SpSGLaE7MxZseuoaCHQK+Hq57nPgsAZfdpMh7Ll13tMVCkGD
06sSYKgfhQfiXMai8XEUwwSQ48uvVW1oHqMaVtvVo+8y5Ohuolg7MXkkXwdK/KKH
p3ttLvlPC67zWKg1Gvylva2PL53ZODJMFCnLcGJKshm/CAgYqVlhPYSSovOTcSL1
J3mX0kpP+5PiBCv//P1Y66+o+xLUqskCubbWXaOa7hYYHR+eUz2SVLuoHoaV3cpd
43crBbwF51PyQD/V6xO2kFWTvxd+WiWJWApc5ELScFtEzz8QoO4TFRAZHSwDQnGI
n4kAZDS4yLbvSy+bWSO8RX+cJLq50Jmbnnz6N8YQ/ofe7WjNvgyuFy0PjZXKlXs3
BaZK5PVgrrnW4PdiI9eWdtsd5g5Gb8hiwDaTTriVr/6V3Yf+njc7qr0auFvbIxC5
ZhtggXVak9R1kPF4NfRzxA1FFTUs/kPQr/0ayEQHdShmqtRJYiIntrLnM8YC1Uq5
wPc9xBQiPcXHg2zGnRmgEpqxs9ueU8cTKfI9E8/z83kJJk1JgiIJ3T62iMhIzZKl
cXQ6GaXluM0bjQR0rwLrj97lLAu2cgwOM+KfBcnd3dfnqJ+koEIBF4v63UFLtjWy
xEmFwXaQMt1DwZ0EqzS97GZQ+YQiTG6sNyZx4mNHhPVxgOcxalTTGBtkfJ7Z+Mex
4c/VwISRGHBR7edz9gQTm/8eCXf0d2N6CKI8VugcD9mR3Etp8iZsHYzHsnRCe3wh
zuAGHfBr1RseMtJNynP6Wz0X28fs1xf++jirN4kaCb+wUaRfF7f8TLbZJ5BPQpIP
QWc6dp94BD0Ld/oplTBn46Glhuk4XCfVQwB5XUWYdQ1tzFSKcjrgQAX+nJ8AqZOR
3dAc31XxW4uU0d+98Hj9TY77WC20fNDpG8crgTdQjri4JeNUf6GAPlaDE+NY3xfx
VtY8uvB2I6dvS/Cu2a2XI3nV4viJKU6yfNEWATU3Wvobl2Pq1UOq5jsQyaQAw77r
ElH13yIrdy6ffjjdFIPRPryPHtqnJgkQKHwDOf9R7vJmjBxPkJ5avr/LhC40ilYV
wavbrYrVNbLz0hsgQUbnx5BXBIFu9j+xbh18phC3S6Qbv2X/YnB9eWZLQB37G8EB
X67wPvWe4ivRWoS1FeIRB2Qzx1Er59NFEBsjvwxpQVduqeQIlkqEa24U2L3Kzygr
urXXwAoBN6Y7HG3A6vpHEshv1P2wiEEArlku9Yu9kdz+IVO/azPsM/v3BhEIudQY
xz9Nf2qYFLOjPXAJjV1aQHVm2gVM0DoH5JqYYd9DQmzNiawTIiO+WvYo/NZmZQcN
6P595g9bVsphXNbxl3SjtrohDWGGcD5oKRw6mxuMGDHV9s7BBhOtWN3LeiVFKVxI
x9YT9AYP8tdh12IdK89LhEnh9eRH0xDBa4kcLCxRGa6NuPN5+dWS+nK2LMqFEiY0
3U50hIKcLo6PZatb2YxVqlQcW6rXvE16qb3Zd6D7Wm89HhtA1Pc4HxjzUIB5TLwQ
boTTgaorf7wIxBG/fS18Ee9TOQigqTDmbUFBolv6EziUoulNFwwEDqbgZUWw1WcO
vWVrT4HKwkg9dGH1oPsYN+LiukljLLgvBMAEAjyIh6JTh21q7c1iAWF02CywkqKG
i12OabHshMHH+xjaeH5H0rA1TVUlnUZuhyN795a5Gr1KGbSADeAY3YdYkGNL4Ecg
sP0wwSJiCnOPLkSRB2SouuLOCBQLSdkt97Wv+WziXDNlMIaXRHl5jwU9cEpXDo1V
hBehrOS97q31O8Ik6juJkvZ/PbDUnSpS9i5Nz8zjMtP3iRUpNMj0dLUAQa4p1GBm
sTqcOZ5aOUJDDbG2J7yV4mo+NDMqV8t9Gsb5ux3JwvLshXBKqj8BCOToH/sFC4Mv
gcOIu0coll8phi2OoVpdZalzz0oellrOnBM0fi2v1QCvMzTnkYlivnvM9ZQOeAQw
/S9CMWp/p+vly8hF1a4rOVqBNH/AcXlNcwcaDo2htGgPeXbgPYEt0EdTFRpnYK35
L4OY3JG9paF29ZGW8W7lW7waoT+h19sEKhbx3ZOo6oydtovccBu5FrVjnG/ssUTs
LRhdZeW1AeuyX/Fq8Rrw0WC0vda/nAZXCqcYz5TYBqyU/V1a+cwrTI0LHRExhzRd
K2DMlaDT81aMQDoFQ96+HCDLSDTOgdFJYTsJ7VEZehuqclFGpF+i/yHf2qg/fDy6
qILk9XsoRbfQuma0tBawZQ7Ek06N2E2DIol9PM6r/AMDctIh9BGOThSE7fTOglm/
REpRBLR22bT4dcKVV8mYjtuGftGYOzNnXlJVr9Jc5B32+dIbMwPKwVkvdMwSHH1k
OG6WTUydT/sAaplo9WCs5tVgLMctPWRQXeYbKr2qfS6q16NYLMkHwy3Q0wBmWyih
glTxxkrBrMI1lDKuGfX2snYYhdgyC62kePanJcreJMvSZEmykcjMJXIXMLBw7ery
BAO4ZizRFeI7v43Q8WBb7N7Wi2Lz6Fp/8PUPCt85yEPAPM17JqD3+J3sNb5j1fVn
huAktxVMJtfUxVK4r3ScPNmBHBCX1IYfTk/VJewFALqDc74gMFy/MSvzVaGZg4EP
OVyvJw1CuANprTvyQ9xSlHFkececgqZOtJ7xr8VCSLSxIAVKzXGXOnnfGZnglFu9
87KHbrOKy7Houf2VxHA5R/y7rAFyzlmzV+7lFhOe1BWCT2ojLi0b5RgZ43uu4Uud
OWQeNo9GHDScgSBW4dSRLrjc83tY9jKIj7O2oZ1OQE9Q+l3RiALLru/2ZZJE+SwX
7X15rnXaUGJmtNkEtwjY8gScRcQ0WWC6+bF283DXyGzreSQreNJH54HZ4CdcC4x7
srLLnljiH5bNs4LDb6OCHALm0Y/7X1u4xXXk0MyTa+eaC3a1jFivmIrJPN1pjLg9
G0+4g5dz3rO7ay2CAoK0bYb3GsFrF3G2LqhNm3RxfdsRAsCdpf5vIPTzXZCA0CAf
AbKknyvH1dRx3M0U3sZuVJK22DJlHAnbu6KVM67HHDrA1v3aCn5EE02n/yhwbBem
yehN8m1xI/fAoVOXoRofN/2Z8xxQ94t2Hqk+82AZbXJJCHlGKopHOLTgFMuLh6BY
0dZpBKEYJbpJ4lZHEpb3ONN445VuWDJkmMwrr2Rt/z8jdK2i+JMjebsZWkjAk4vS
AOTli3rIqGoLcyVSu4nRPk7mEnODu55hZu07ZvSuv45/E6Ys89g6itAn67l+GJ7w
QmEZJGYnYcQb+c8/tqoWY6rSjwUWD0HIuzd+vM5W+MOB1CzQVjvc5WwM/pD/NxVn
eZYTXQRzKAq5R1nC/BJnXkM6LW99QwtHRlhtYxMH1MXvZh6NGrE3xpl9Ercixony
IrvNR33rmpubUDOURRWPYFM3fOIMwyOdE9g5c6ewEDHBjrYYBxJJmiJr/s59AJ06
yMYIg1J0fovoCDVdRYfasKBkVnReYPge5MBKD8ndHj6qJGqM8Dcb0HIUPMNB3q8c
UfnmvET2p6E8hRWYc0QpSR4nYRnRNKKYbv+V9p9IAdbdugTdrIiUitmn8c8WIwz/
GnyNmeoCXKxRCuhmXM3V0GzKzu1je91dagZfb54qMW+1o5Dsa4LoBaWjG31ZIYxn
c4PbLpPGE7NBDwAuHLDNNa8S6JzUuAX8BDE/s1KWNbet9t974os8kBt1b+LYtIDi
GYZ8Qy1DEw78KCg5ZZv1/i2g5ufMVsvU4toUTKjuecfI0IyG22m5zay1T6y/UkKM
v5BXHSNturEz5HebqfjArL6TZypLFR8zynAWyQtu4rxQiJR08pmjrK7H3+NQsD4W
yj3+XsbYdwJ8CHmGtsmPoRhB4b1CJlwdtQOcuaA9S5QUikVrArfBS7n7eLbaQuWw
q7kUYn0NL1SUlZsbZDs9ny+M7FTH0ZuDH9qEm63un+3GBSs8qdR9IGmbKeUu3tqL
T/Cm7A397mbFjte7VdHVf0g1X311mo5bgoY1piAMa9IFdmx8z00PKjd53Z59PuZ1
nk/g7NoB9bB/uky153Lp07uhItt/hFysG5pRXxY5JGNMqfrj9PNrmIpiD7venc8r
U/kqN17XvYuvW/WWTGMO7yrHJjItssHEoJ3EZ+MkENaHHTyD+1gCj4ztkvZ/VUut
RlGXzovq8wV+aDWaIHGvRpRC8KpmUzocluXv+UNz9CRAMqToXDxQMKCKYydeu5Zn
qe/aPabJhqFtFyWKYyK38OaiwX19VKVIs9pMosDYrwpaZZd69OUh0lOQLmQQVWrB
mwjwCKLzOJtcIv88rQInJmLrw4LKcyQZr+NU06pN1Kal8AyuyphWGDDRkxBbbCLW
ivHJ43TLi43396t/JrKjVE9g3DSAERCwMq5kO0WDy6h45TxAN4/LFhcHl32opYJ9
MAPJg2YIEVhIVZ4fAFqW8TqQnjTXuM0WL4IPHGMkz3yxewtanywvVkfHjfBER0B4
YvsaGQSw+aGC1kLFBpLVbQ27R0xKHtsxK05lFTTJnIK9eRHUyMMwca4MAW//LR2T
4/50ccQ9BNIrKZHKUjJ78KTYzQ07ZzsRFl7/PuFL8vej7iPMmrOfdmu2mKdar0zI
uDo31YX51O7yYLzTjuJkXNvJLHECl5U3xaoBGjwoj0V9B7eLWQ39YFjm8btLnEnK
4oWLZTYQtYDT/qfkp8EstJhPO64VsDhsVXaiF3vBOXKZTl/lkBxWE3TKphMdKG5j
D+OHURfNOu1bN1p7l984VpVNrPRz8imc+AWppHbQoLPbhJi33S14LQIEl3oVfIz5
F7BW2RFxIdt433A4AEcySMN8sWZLNHB9PTVUdpWX4ZlwGHi9ACBSohSMS7HwX94e
dBVXNO8sF0TsfPEMI5Bgyskz8uOH2vaufjdBewGM8rEO5MxhKmACuDUClLVV0cFU
yL1G0Q7nBADhxOvU9G6K8wIw+7H0jPuZPTxN4CcxYxaKc5HHDD/OS4KP3IVvnbjn
owGG2LMxtB1xmM8SosLhWBB0nwXDDtMRTwQYMIaj11PWAl9TfgBU1QBcFlCsy8qN
bwxZmrh0Z+U/z8Sg3hFPYX4BfGu6w0Rh/b05c4Qa9hcpOKYa+GZlnF+TuKcmmlXs
nrdA9C+EGVv0oDIIXMp9kqYYnIO4MTdFej9iuilH+bXP2hW09oTLBSh1BVYgcA4j
LppuGjAi3aXmXs+YZeGK3jaZi+xweTRU0RJfAyo/SSuVzINp24uVhHqxVnXUf7v6
fFL9tLrNfbCVvYsBlIq8Xhaq4p4dqhjEUFDzjuJZp9Y+/NlEv1WAEOXKDWAFZ9oa
YaQ6GCAuoL+oukT0oBRoMP7Igx9bSb1R3Hexahufp25eFBSsrMgy9JGT2vAOpNLK
AbacynkBU2UniHiLHSreq4fimlqPNmA3sfxgZ48yw48WbYSCJBL/cki4hjaKi91l
dppq+nBjlNAHAYdY9wWE+6EG8xgKGDih5NC3rJC4WXOhsbI492WuespoF3mn5cjj
J0D4y/L/p2uxX9JcKobuuV6R4tGYqSvBZhLERykchAuPFQ07OfPeAT9doJVpsS42
PbazPLDneboQJWfuDuIAWIGtHF/uAgC++kTjR0mGoo2ueK/0DsEmY8uFSMOydVTB
x3QDDpYQYIGsA84HfJCwaMC7OcfKnpkwRGKAGMjPBl3jlUaKx/0zfIK5BytUI8M+
/kN75+81GrC29P6BFMY18lQYKYMGvBiADKMF3KRr6/GNQgTXx2zQiWVRcVsmrDnD
iYs/JIvvxE3190dMmSVB5+FTlltDQmxYiEtUOQiJzqy3cS7bDKkJKx6f4JJC8eEq
V7phOOkYG3NSZaIMwKginRrcAXTQZ7zNLHIeqU+IPyPPKHAbCovoCDXOpRgIdOuP
pmNLloOaRoahgTV6yO2f7zltlxWfgrE8nYr/MrzRqFq9uoKoI88Yf2533ZpHWI0b
tYmK75yb9BMI1GQDvDkf+Lxl/jxSbEsLAiVApjvADfOaSWKgUj5pqFqOKID0usl2
K1rwn5+stiiMa29d63+pfXqWze2s+y6AvF6whZzR3ZfNT2zVd6ZQT13IH8cdwSgS
0qff1rHudT+l9n4TNterRzRQaocQjVDoDV5Iloi9/LcXZZ9cFl/480YSedKRz5M9
ZRd28pUYcTiLC9/g7v0PGxd/ZSGGsepB6gx9QAlO6eVkrD9juZa4qWuqnIX0I5wG
pYRKuPxLy6ZIURfVlYu6sfMpe2VDsuMiS4mTf3kfXRnTOvs+JZhnBSwQKO9QuM4N
frRHk4BWW+/YSTYEZH7S1c5KFbJaUln4CB62GLCFQyKsmgnYBLQi9OiATi7ZeGLX
vH2ZwuyM5EG1448vWcuN3m2/PcGyPlYwDDXJ2kkqSJm92BvhMtNZWtAMIHsXKFKp
qrntlk6hejMntsj54/HNVQxBjlYWQyE5cMb2QZJjuNvC5cXuP+knPEPk3OAYfioT
6h+FEyfH4PLXvLhBxuA3ANczi0iO0bTLfH3fURGy87UW1CwkjF9xPJdAufOd1xls
`pragma protect end_protected
