// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:33:04 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
nabHA0XOjLgjp9NfxYwX+nfQWiuMH77XlJ/Kf+3Doi6JvGMPBUE6UuSqcS95jLXT
zEKTHwYtiTPTC0/a0O3l6tXaXjZMf7yHqT7ffQrMZpwHr1SL//f+UFFMgKPIZZ07
Y29h3MlKf7xKfm+2O/7aWbLr8ETlKg5q2zZZ09BBD5Q=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 6304)
MDRp1v5AEcYhFl45qSnI53UpJF04ngFkQAChHyoTzNRphairSQ5PtnMlTa2s91ks
u+CoIN/gJUZTjuef57ZzDF17REBRszd5Xhe5JfIM1IojOTXO5y1MqB4AQhrumTdh
ziJxrClF8UJkK1h70L/2nv4FNhJJK0XnPXrwJT7Ahzj+t63Drd557JOaNz8eacEy
z7beGMcGZ9lZCLDQ6l4xIVdv3+6z80tRBNovrDK6IvsrgDB43bB6RC1UJCcHHCpO
ok3osGiQfydID4zkSTQHEYMkfwV8cUYrheIUO4RCZKrwmS4PbAdxKT354tAwwAJw
y7p4cM2vTpiH/QVVZ+9lWFOOEfpLqGso/tJISkE8K2mcrF7vEifkeohWbmseWhB/
axpQuxAhv5Mb7v24/WHVq3rUcXcHlOHxAs8IfoTLBdLhpmgVGEMAX95QYAyGGWNA
/H8lm24ajFlrwbdxGtcETlAZ5hqPZ/kXMfXb/mwm3w9RbgNgPEbTMdThE9LJfN2r
kOkZamPDAtoZLf2ABhRmhvcI0QoLjNXILpPp6FHHlHKx2mclE70+SHIo07f/YQzB
kPsGGfCHBBWsR+wfbG/MOGOzAeqeU4aG8WpQ3TG1WdgK/bEtSJ55CiP5Qw9b/Pjn
WXNYnUxs4xR+Ynrejy38cEc3fsMSwIQiZnohk+5fz74jfTh55kJTnrArHSqb3PHT
TeZy+jxvDiDWhaGn4xOHefW0Hmv4I0A37DJv/VLhktbzAMdL7CRuFpUNr+cU5IAF
/9lQ+rn9owCbCXHyHMKgOs6ioxIYwbL4pDRRI1+KZ7X4p2T59cXUQVtd3F2la51p
0ghHxojirjZExZdYPVLsCCiRd+vdwul6m3Jfwz0IeJfbTkrSKN/YCUKFrPr/Z4Rv
6MAFllHry+1PJU1M0c6B01P1Yc9EGCZYB7bxyImTLYiX46+rP64/8K+BNjRC3zSc
i29R9IMahrupy4RC3dZcwuzkzbtOPyjb4l2L2Qb1TW7gc9m9t7e+xsWCJJH7BAF+
nEFj+kh79Rxjk+o/9zP2b4q6lTd4iuyP2Isuc8FET/oKblPT1c2SiMDAplqp24yj
mVap3JVe+4l64jDqRmfqFrVd31V/e48dxoLluFXbUwC/CRJRsdqbeKj5h7Asr/YE
zbhcMC3OuOxQh0L58Z/Ag6s0PH0EWUOOIwTTyatuK//0BDd09UiVq3EknOZLHcgy
aEyONAU++9ut9LYl8/gfqNx59zDoKZqm59vux7OZOX1K/OIadc49Qqoe+NHQaHDO
P4Cr+vjzOgB6wnzTVpWsIrawqK+K04gI+NiJCmDHPAHaJC839B7dRFU7lMvBDkmC
0xVs0jVvPH1pHlQlgQiS7UhN5/mlhvKLhwe6v76cQgQGWFBjfXJ6gN36I1vZW11B
jgXFaCmzG38ukJY4uacoK2eXrST+1Vund7TBavgY4pu8VdQids8/ol4/47y6PbRw
3fdUm5NlXktcJ4PBsjhj7dagh83hD39K8FL4FfzbD/mfrTX9Nj67czplyAuHXTny
dQdfIdAfNnwiO8eVjZwNmzZW0dMIrBnJf9TcViwmhuS6N70umVGVXxl/z7k3TNKP
+cbZv7cLY7v0VT8fnM8XyZL1dq5srrTe+FbS7zDoYxbkBDnECPuY6Acbvsw0EVkj
brhqqSKk0VFfUCwTsdzOoflQZWHDncMPyqQ3kH4vJxeC66CDOqJsqfSWpvWuu9S5
bEW1qVQ7KVvuaBX+oSTn9AXplUeFN6UMwm4ggsyPIxUfFa2nIzSDa+pbg4BzG4+T
Smy4X7TFm6zfmb/pBuYI1hmXHGHiBqQE9bYc1x8hChVVM3kSWqq3//LyPZyX1a5n
bmWFW085Fg87UoAT9+jO3LLUpJDo/sfKUa94YKYO4iedsxQ2Zshxb6ai06V6f/Ex
j6KjYVP4lU0OwgMaWLyL0YYtTIDA9/cO7s8Cep3xhQBEp5S9aWK81caLRcRSefnG
bQYgJ1YUcgrLkmYimIFXKxvZtbOptUxNTu5rWy85TgTSadWP+xUQeUQb5yR60onx
jXQvgbiLTxoU4mJaJxlnVe/FXimVIptImJuFiB/NkHQcbH/7aes0zWwDldbdbRD4
fKTCVIbdeyX4VS+QJEhlfXpaLNqzvnlXoGjV3a8BcJ9pgWXKUcxQzrMi6LGaTDSL
T07JLxFzvzYQMVzOZMdHarNZGgO3FVn8gcrG92SHdcXykWZm/Dt1UTxw/Kwy+cyW
aH7J/vIW+t2l76EGbbFBYlihWYkuY69Z1Wv7x50fTmWF4NUOpqnRg1Wa/Q9Q/dvk
d1MGMcuyjwZcGHUGQmejOHgaBlU29TKAUHgM0RN9KMkxRmIPVOtjKlxCUnfp2E8U
CFX7UeqSAxad2KoVO6z77gz9oN3iHQXAikxXhhxXW5c2+E2AvZRIP8+PLd+BQjOh
O/wAvB+P6XrV9pt9eY/YIkSHVtRLdo5JGPmcSGv1yun8wlhX9CNvxLlyL+lbweP6
wo4rooUDHnO6OFu0BuZZfB4y6BXv/HIgT098TDz6LfRQowGRD5DIqKPh4fgljYbP
YHtnJrrXT+hKJqbnUNVE91/5NWB1Cx4l7U2tucW+s4XhgQMxDIneEgae69k0Cp8h
xzlLHDCf69YROnm0y0DqPX2ZYZpcSUKrnL3mjDYQZH1R0fJ+9p/AlFQT4ojSaaf2
tBDhAGQtn0Qe88CvQ75lIP/DaBWHQn/xagIRmzmF4jZyym0z8RfhcQiOtg/As+7L
Sgl4hyAg+zXG+XL31jHPyySVhC0GgRPk6c/TtJeT+jCIizd9IEkD4CIVG5NLfLP/
ArEP1gp5YityqRYF9cr9r6CSfjfYbNITkv5XbiN8vuMjuU4NbPxaiSPANE1VQEe0
OWi1gmtvT3iWejP4AzOGCuwikMtxMXXMhUlL4QO+WqjiLB6BHskZAv6gqBh1/sYr
HXXRNMSRKbNiLWBZi/yGgK36vE1BiSSEZQbRPts8envX+WQB9GyYgIk5xlwlqrFR
EsZ4dQvyDETa46YWOon+STPTGB8kORgdZutraxragblZKrQZenXzssn68SfAv1cu
nxPqRfXH0Q6rmOaw1Yl9f2SXsgi44j4kBetg2aJjnwxigMZX3Bx7f6rC/PjpsHgL
iK5r08gkVyy0tKjJkeNDDnAb6e5F8UKBmQynEpBAik9N6ssYjjvFSTc2eYtDuZKi
sE83kh1zU+dgPOUhnhU5QUJCVLVJoaORjBzjE12YqeMTxLj8erEnpXcYdCUE9ZoC
npGQqV5LC/stYk/HQ22W8CUE8BqTNAl6UPCZRHe0NdO85xKn6NeyokplH7m6GJqC
+ZQIHTGTMiYM39D/CfvFzLJhnZPVcnWuMcefMbeGwgr3HorIA77YAbXE8GTK1sU+
cAAUIXMgtUQzQXNnFnOiNQKoeukl4xQmfRtd8GRbSgA2UACXCO54O4dIASO2INbg
WtoRzDExhC2n/9NW+V8yu177U0LlpGgf5uH+FoildhxFNV1bXwc6LBK7sh6WUt6f
PVOUa+fIL98gksakRKnWAJ/NpbX7mSbWDfvDpwsxlMlso713TnqjKExU+V91jVly
zINr99hIo+n99QLgPD/7CEenBSUu8kI9yU897Klpf6CclepcndA94qGYlQpDjIK2
E4ZEc73hLPT/LqYQ5BoxJU8Yc+QE5WQRfjePYGvW4i2SD6EVw48TkEjjjm3owsA9
uXSN5tT6j4kmn/8h1Fx2qajK7bYNwUVZGmLP7qWjLQKe6WDYoWnJwBHX4HMnrKhl
5d2ct4HQGQk3Uz5gz24Uk0yrxYk/7LJTwj34+YK8jNEUI6Ru99bwIz0sGI3VVLDA
8uVhr/9oLo1/wP263V886+mN6drCp/GvlwZE/WLd3iwZpvbmWTUMNYmVaa0Mzbd1
HKOfC6tfoQAlo8Gj30h4/lX8HbUETj6laMFXCeSIVIHPLI4fhtVeLpMpKqKHH9j1
7pcjHZMwH5sG7TD/tfYgea+ec4PyPEEY6Z4ljfnG89KSO3XH0lDXI0+G8oD1CzuF
uFoxmcjW/WTN/1OJ6i4O3fACNtbW/1eovaZSM4MmL8tb63tty5vB6OvH4DCLeedS
2iBIp8HvKfZBZQKej6k1sE+crgJnpeEw/PI7e1Wy+y64T9g6chXCNArq0W+XV7lm
euvfEDKVurTEAa5o1iQZ25mn5A3QEOcwn0u+11BrKUpdz6YwQbqGaXM9QvWa2+oP
rOWe3w61/UHhQhR3oMlXbQntkwF0GrMWwOb8Z5cu7U+ltdtrqpvC9iRNifpM4gyz
9r85dK8shRb/aU9NscnOSQ26MuVK6mABEGjsGHjI8OMCEeDFuxic/G9yny9xWCpy
KITgFiqmnPp8H/K+yqNXF4KwLF+P7I3ueKZLQPSInnxIHXfYFvK4A6DI7jikNmFp
fCY+8Cc2Dqr7PVkxJrXCJ5O7Le3j+Et5uwCzo0M4K1x6yOfgOGR4EvlcfgsTJEYm
JvMkEC4vITk+0lnoAkIVrdKyY5mLvLiVcJTPWfqTT0dritxWdT+zuBBbzYEOTNA5
I19d4NJ1WPIKG+8n0+orncMK4J2VGPb1RLAE6J8C6Mk9toToqOnJ8FSBsOZEuykH
9i/mZj0FCL1cv3dNftBQLj0jLLBWhvQopEMurKNGXRaK0fjZmii9EachZybibgmw
Bu9QUb4h14IjdRj65Nm7v1i1tIPr90BJ7mP0eIJtveOTa6HWaaueFF0w8I2I8Gec
lvDmX2+/JS6QT/wOWeMyymjKFQBUc+L0/lbkknogO+zGAh0ppRbd/m9S/FCFk35/
8mwkPtHEXIfJPAww+xrTggl69QsNUOiYZshrfrEWzrQRAD62hO3gpPg6rKJf2iNw
L6H34Q6Jb3FYU3hSVGMkRGhVbbFzjSNwm2R2An+q+qbUqZDPvhQ5D7Rpyr2tYl1n
G/LVJ5Xx8RaghgDJM2gxaPP7T+WIIuj/p99Z8yzHFtHVvxR2uoBMAkMmGSChWOwC
mvEMwSpubbQqO+ydscxZ7nukRfZZK+Y5Dwp6fias4MywZtlbTIkBWmdjAwUsBWSK
54/QZVsrElZPyDyQ3dOFHa2ihZ820aQNahR5f+VdElPP+l2Hr/IQw5UDGdcNp4YZ
v6dK3raSBecgbRV4sYonHu3YTw/yrUOORY805LWNAwVXkSiM53A8V9RSMWv/Igh8
0cn/vgnb9yISJ70DCDXPdWdcVjKIcOZpVfh/B/V0FGuilMWh5ZHzM/L+O2ZASDTV
Os7J7jv8Mc/PdpnBtnugpzWmAzMmIoJL8Te9UvTsMctsT2tAKIWpLb9dlFlpM83U
YQcn6ed3eztJo4Ccu5WNl15mP7iyu8AMytkJfhtHSXvEsZC3P9FsFGpw+aqSufZQ
vGAauO37PRF/5Nm6EctB5wO/ThpWzRfzKmHnJWpA0q34Ow378w9mDOa19ZLN6Io/
vw7UHXcsCxHgPm6YgN9u6NZRGIj4StA9pcjxy+8ho83UyrgZxiajOEPwcoj1NF0/
rUTuryatM7QtG8jpGhUWFw+G8wo1biOp9tEmUYLuQ2nLsw3qu39kBPU3hg+AAtlV
zvQW8V+2HRnAL1jkNZygbqNP6hcqmxgyevVVDk8XQv7RYx93Hv6s3SvLpJ0KIbmX
jiGYjNYJOCXT7LgEhCPiOl4CShLUp4FakWddbmti/YtoJUG4kle2rAMOxF7q9sFF
03EPbuZstjTHpcXfk8Xy2wJCedxOmQ7F7NsL73dbY6+TuZjjSq7DChwqORhcKCeP
6yl0gwbGA5S0zjSii/cRfrEbQrplWN9m8PcXKzPLRKxe/pDnkKUh2VDjtE5SmWwv
B2di/qpszk5Es+E0ydwQmmWs8XQFYPpG2Gvmz2/lXi5q+Jlk2igg/q6DABvxRcfy
CTqF9jaTvh5tZYvTuftD3TYv5YRx2HeU+ySu0XSBrmAgosQnMMqUufNgjO4OnKiG
3Rna/QKaT0Vyy9fkFhyPPi9mzGdefwPane1t6cksZV0VHub7Rk39jAOdRBpMjmZB
BIJVr7i/NCEHIbVZt4K88hgTwla6APJnuU4ld4IPQBeK1/in+iT6A2G3MJibDODW
cU5Q3Hzl7wfYc/e8Dfu4Yo9iACrptUs144ILUSPi/4cNJMq0e90CKgl9+v03XcP+
T4mq6/TCIKd20cVNHbW7+d+knEb+er3XigEmYbY3zOquFa8DGbJJCkgOUSSPfZCv
BfpkuZBr2NdT8sKGsf3wrY/1ebRy1hZIdHsvaV5NTrHNWrMdH02mLX5YaexnEw10
Us6vRRt7ilPMnsLAG4IYL3uZoesaSaCzV3fJzcVD29jHHhNhHNLr1S/XkX8YX+9x
+TXk1YGcou9utXQUKox3oGqUAJsaS2ujZbWLCLA36F5OyzorhhCE1/BCDbHdLPmS
UM5sgEkPcXPo0C7G2jP3+nDkdzPRRe5mgVyyNzlR0hdrvESklrqV2JjY9NQNY2Ov
yerAKWWA/PERnH+2m6Fc7RJk27794PT+mbNWR6saXojuzpBHjh4psXrjZU72jIoa
o8Qfqi1bQJ/TkoibH8JZkOZ3oToWSffgN+A29oG0FlC4fVTJBVHC//NJVgI/y6U/
2Ek2KIyxu7uJ+tA4HfcaUv3RkXU8Kss29zK7KVVhy9QGyP+CKQyLU+TmKg7hFBTB
k1oFSuFGNAt5a29j/J9HpWTSwWLh0FJ/9QsaENVEJaIUfZZnQ4gtgW91ij7P1VWZ
R/m2kaCzQyuwVliDY6w9m5+rpSg6qxiNauHTD5SZE6gPXBR8tWAecIBL5+XuBU+O
Bv6wUGy13qcVUbc8N2K0bDAXKa/tBpUTU7czG9TYHRKGsfXFUXypXbTtv6sSE8QH
Z67E00PpCIMYz5cTUMV9JWCDzvvjbcZiKgnCwgtE07NapBxaT2eXuwCTrn8aR8w2
SHq3NzM50rsBKFT6vW4S7C6BRWLQ2afr+LkOSDtj1P1nesJweJ4RGqUJCk2wmGG+
IyC86ZfU0PSpfA645XE4mdP6CdT7m29lINEHiuOEl3HysX5MUkGWPSktVkHXZcLL
p4MwYLA16rKxDfT5ovB+06k4/RJRcvB2eAeDxKnKh0mYtmXwUxtRQ88b/sZfFgYT
m1eR+j231Y8Mk6+4vd044uB9BJ7hrGC5FmjnXdub4uhlb7VsvLDIg8HCY4c7ijQP
D67Ori+cugQxeLGi1UuN0HbcxthhJWpguKMBalVZYrymkoZm9FGbwl/trW378mMj
Pa+BCB8R+XdbqdgcUAS4yPSzOQLKzAecYUEywPL1yyrpP/SAuAh9Zk1KAwZDt350
4Ke5MdIoG0zqSuK7I9k03+ynEjd/2545RIvlvwLs9Y/5y1wKyFDqDflsIY54a6El
mUkqV08qfFB6I7+GX7bdqmzf9a2RFflXkZvqx1dLaqda2xgpM6IjQ2CfTuTF/Orh
ohaz0Uqnv95xhZJ2B1vJECmXxFdQaxRtMcFrtb5HYNsOte0P6cJidiKYECUxLvuF
Zyqy8civr6Q0NFES4j8ZP31qSfL/0LnGhOdhWc0ib1NbVrK1HOQQVKe4lX4c48QO
bqGVNLgcZiSinahb96SLR/SHepZDF2lO1yjOevfhiQofVqK7QDv8m+lfAUi6ocLR
4a/Ve7u8kTkzHI8PSQonjXWZ8K7dqcjCUEfRC7RxJE+O/RbRmHNbKm/qhuDHK9aX
DeEGPbHgPQDTlOpfasfB8ov3F7F9AeMEoQh0e7uyRWfL6o3HOmXj93OizKYWJCcH
Jih0Uf1kyAxoWTMzmjUFqKBMTTFtWNNbvSlldyMzaLO/ANDIoYLo6N6uP1Qku5D0
kvzZkkC04vWlqtDGPBtNxXW5vMh38QZBpyjKkTTv7Zd+Wyo2P/zQNP1qkkneGozT
vL1Zi8AuF0YuAdtWfmcBzp8tG32BdOL7AJpw2/BgcmEf5z2NV0ZlcKvOnbsE78Jd
aJBW95JPxa5IE0y5dVIWCzVLuxJJ9UZ8Wr/gu1WbGjCGAQS5XIacKoqySriEeN32
1Avq3108PJpadw2SQMajglTg7BXyL2C0ICZOeGFR6Lr8tSIbOrxqxrlDtzHXDoz0
/XFgn+bGdgtQCEKn3p5JWJzFhIfDSdXQMcvNfqQ0J2pbNZjD2BQk+zTOTeWniar2
drZTlmLiS26G8qhwohpspOBzbZ8iLTLuv2N4ClfZ6g+Pm09qexM3B7hQA3d0Sg2j
iTmwyza3K9aNgkjgFDKcpFGfbI5kCU+nUQA+xlKvn7yC/l58PbJJ6TTmtzTwhSXT
7deURjBsKiEsWNgI/I4EiCriak+cCWMWWlerviSt62fOhsVHv3S3wqOsoF1RG0Ca
NeJ9c2KRpOqga3TAQM1Oh62+X6MK9iLvx5jYHSKwtE/Nmb3astEtJdQKZQWaIiB7
78C3FA/QSA48DjYNLa/4DQ==
`pragma protect end_protected
