// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:32 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
foCmDMWgFO7lzgA4flalrsoOkmdpjUjo6Snt4cpQll3pCB9GS2TdO83s1x6YGdfY
jAjuoFkfgcEc6RTgMoh+gMIzmADVQQHRPbmhX9vmKgUm9he9ziXfgcr7g4tTfAe4
im1IoDahUwwDjGUS7b69DZpb+62qIspkWUrZZnmrnNE=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 61216)
T3whPvntkZxx1EQ8Ugeehwhdf0mRt9EuEoon/QA40gQl/JHCXjrgilLHEx040EvP
SIDxnul6RC6av2A4nqZ9tNUmosmO3/rSEhGRwbMW6BN+vhCiX0fctYoJmSDjCRRP
ZxoYrwGC/1xvPkbpuV1miZnZRD7wwwePwDl5sRQeV4j0U6BVY6dVm9aTbGyg9Wrm
xrUY5gYhrN7lFT/7Sz7ceoBksiXPbJuRv+lmhvCLSi+Be8rdHBkt+IruKeCj6cEy
YK7bDPIDQKJGSLsxw9sCsZRyDvr6i7nOuczwprVuW0FWtqvyEkzL2UCiR5FS+IIb
ztbnR5famPSatDyWAWzSLeCz2kxzVHubFZiYBNTS4POWiS0K9IEF0/0p1ul1G9fZ
1gKj5h8yO+37YlJq7wy3ypAT8TIaH82E0AkDcCl6m2BX2B8Kh8vOWRJmsQPeWhVF
CBGzK6Zvt1RBRmooO4uRx18HUrf4Hc00HlrLJ/0FISxDZXv27eYREVnN8fhHXotO
6kEp8pISg3wEfr33EiXekNwqbwCDabbH05pR6qH9OoC19KuPZVIuJZ0EZ7VNruZ3
6kiSXVC/Zzl6cLaoqwr+z743UAqefE8p5VBtTN3M648PSsK301oujGZO+3158L3O
fiDNoG76eJuKaCx/bwil96G2TSOaeGMTK9fsktnewOwlY6j9jWTP+XlzMtElvGJa
UVgYlUepxcHx5Z+bMk7XaEnZvrbbhWeRISqyXyssozdZJR2a9l+tC6jU7FogKhNx
euDmzHrnXiE2rh8SgqpBriRmtQWfnkBwTGsv9VBa+i/oLlliNNGMdoHN2xv9o5Si
hHvzreOzygnQToySpDtgY46UjeB/sQtMyW7WBh67tGovXnm5Io4J/eM/LjKI6No8
VPsfxQpbIgA8zc9bW7/821egYIIzDuDL9SHVNXfAoVTFhoyz5wykAyRGoi0Ta7Jt
bz9o5yGpA4oETbdncjccs/skBUW3jfoWY6PfzkUNPxTJ4ppWa8lQIPzVFVlLnPkD
2kDuL7CGFJ23Ev8Csy9KjEXuIyMwnUB6KyHJQlLLwxMFxZ28uq5VCmNrDOuufnrE
ohASJtG5nsoU56kedBh13Ct4qeg5XpOcj54at5m11mXPBYJwq/mebZ2V1C7zVd4t
KN590iyHfFY3sLo1IR7lp8OoefkJvaOAh1kzk6+2T98+syf94XnQCBk5PsXkxjXf
q6J0Ff+eiFKvQfUwNFzd4L27d195MvU9TSnBP//aMYeBbmL9/BRGeuQ1kXIonT3N
FBs+UvXzsFOo1YNLd38XM2SOxTP2pe71du4pomTheZe84d3H5uBaUkH0yiON9HbP
U/QRnH2/YX9UnKwyri+kQZkS6OatlhaUmX7OJZjmeJBIzlla1pKA9lNWBQ7rq6JJ
SzgrdoTOju4eAwwpcYyvMRhPnZ9mKwbt2tqtY+Ht2rgbiqaBLaV6HIO5FpjxRk7c
SGw85SWVca76H0nHa2aC8VAYsWbLxBK6NSXEYwPEoxijpP01OJsIJ8/XewVofGlL
uHAlRYA9X05zsZwXIcQQGCMk2oWUiB96aB11bRC2Ap7/x0j51NSB9hVpg+lgwlph
LAD+PTCUQuhDObnIU4R3Uvm6zgDtW1P6Mz/j8Mwtu9CJBV0rkl0QuORp26gfFnes
P9DHRYqvzeohI2hTuDEhX/30SgCFOjeeFQJddLysi9OF0h4Jjvxi2+upxcspoj5u
b5TjROc60k4M9dp2EIRTGWvKSx44KmkUfbvcKsZOArncVFJ60gzamnxGmgw3+uqq
6ZUR/7oXT8UUqUErW0vFhrJzOEuAjqKbZHQYxBNtB4qQrqNIMsbBcsF6aLUviCkd
TdSlJmHX8kKp56y+zS84ckOIV3/wBdHqD3spI+b+WcmojnRbpFq5muJ6SEDGHp3f
a2x5PGx0BCG59sYSBpTBtdPW4HY7UaulKNyGrEKN5er9tNR4+VI1Jkoy+zWfJGDX
9Udo0mm9uEFjde2kZYJ0N9/x68s09KwG9T4mCrkucJR0mCO4fQa5ZFYXc4z+VN2U
jRNkqGvSc/Nyv1MtubnV5qm5Lotj9ntVL11NL0UTspE6swBkdBXlJccdK5Bb5+R9
RELgwa4+kdFlC/6pcfJmIrv5ZQ3RIzMxRaKWDUL1916P4SNDwv7CKHp/YS5SD15b
/TWdTeYnawBnxnOp2S2CpXA1/exM5KrLanKQEpj11CJdrS0mQSy/5GbinBbwV8wJ
t+frxZHjPBY10ZuioKZiIQ5huwy078RvdvIRBeFu4L/FDHOJ+FQFl7fRUPXBJ7fO
11ot6bk8248JAQUX28nl9BEKJBzMbjIRWkKNzXZiNrMtwfyVv0anrf0CRsU4Rk7g
0ZYQfozkvu86ahC4ACqtiECmk9pMCJL4S5RdiJU4AUFwvwECRiNQnhuAjcUSpLg+
eivjZrGxrm8PDWv6jDjtm2pqrk8few0uPswNrTq7nNt8EViTwckUA8W0X+6u1EmX
7kir8USvWfCx9ccC60EDHSP4f6xs+EyaxgH5aY1Px+SperiCEvzwMEzHwzqP/2RE
3DF5RhoY/EgHVNSOKA3UYqEy44mGz/HkAfTTPvac2YI9+1QRiah5llD/lNP6WUCv
OgWkoPds46/q+rL9SaaHGXjXUdRxGtO3r2tgSiVXwTNRjoK/lETfO9KYGfoz4bS/
+UVnwxhRsFjEqMcCbJYa0cs02Nkp1Lqcx0HLR6skEQ+kLDbyUj6wN7fw4Z/wLdfS
E7xskSwNVRr8/Bboqe27Qd72JBVgSQOyfsNu6T4dPBg3hEvLsDRkTje5yA3UtV4q
Z2p5RSgotjgvUzcicgF9ZDGc2IbxRjrjGC2ihGGkrQ2tltz1yXRI9cDOLK+zcvdo
HiXW2NM6mWpAHdag/yCc5Bwn+adTpxFYT5nf+QrGFF6IXg88HeBPqTtoE2g7qFG9
su3SU9ih6hiQlL4KCK5Qsg6q4i3j+CIkqUt49VjeJBbOx4BaMdqACL78mw0Oe5zk
BrE14aJ4eIg9DqGmFbn3F111n8yjCrulGm6rFUXPUDllBUSLv2bp1rql4u1u+QX9
lET6rbf9/U5Dj+hWtIyHW38q9LDFdPnyvSn1M6Hrl8jGf30AESf8r6vtSYaV/sCm
3lQZIkS0xhqk6DHQ7TCMwV2lKBxN8kVIdnNg7ve4pfxzQ6FwiN7GKPxqPXR9WEQi
gHZu/IJ62vKG+PBlTo06tqByEsW26hHE7EKMK+RdT3sXvp/e+kaUJJcUVu7dGRG1
88aTuEfz3gR9scIwMdn1SA8QOao9TlhJN94bbRIgXcFs2rYgDLe1m/w/arR13uiJ
nHaPRMwGzoZ0toT7Zyhb7dxg1UKtURJG6RT0izZWfF6im0pUCbw/S6Oy4pVeaK5v
ECZgUVkdY603uCTcCxU6U754RmQoVB1T+g/i9qFS4/s1+wAUMoux7+7QHehGxKp8
WlsOeR0eQQolJQXorF9c4M4nflANcHlpVmIKIkTl2WuN32/jgxrBp6gyg+ol9Ybj
7tfWtEMvw98vrM24lruwHiQV59Qn5sCPgP29/l+kTEJibiqc46O80MrhfEN6D30Z
tadYFLsYvZQO0aRfNSPPGr7EdVZIuycH7TkMTX4sFFpjeSnzLqomUCLvLNP94OBn
Oj0i4tRRgynOFxezACuXGAmjjBGYs/O+5s8ltr0lj5cP3lZQL73KuJT1VBkVW9Jl
k/ErrzEpbH+RlJIC8kJVQXn7fAzzYAf1GPscs62bFqeCwvbwjV3fERPEY1ySA2CG
OuMnb31iD/UbBFuuJIsk72Io7Y2VRulO2oWfBKCFAfer5mNtng368b9mFK1U39nB
7poBAkNxNlCsUchvXgluhV6l8ORXdFlJXUtdVwdVoQgiraG8FoAUfbGgxySn/P+I
pt5i0QwEq2Y6iAKhML0b3z7RahSwuAKyqTN4DWUbuFil+L0psbRmZv7AEiRvtCmx
589PvO3bsPRnnsWxMgVl6tG0VPSxYIdRTXhRpY/A3TGQBjGORQ3c484O64Z5AtHP
TrRW2OBjAFgtGgpG5qTOGF6N4DBpkW75CSskQOxhOLpqcXUSXa+axp0MhJh9UDdH
qXvuOoHg6mJle6QwfAPwzc+hjFGUT+e829MXrO8zO5t7lgpfRGGxP52Q8S0wAciL
mDe4g998wxsGGAD7vTB2sKm02QMmcbTnd+Qfb4DHzVWHOE61GdFeQX/Exsr/pFVy
5JxwpRnmgfZu35Zl1V1jAbqb9s3GgLtL6w/i5JaXmU4RPw8tNuFbgD0Ii10PB+NP
bifvdM5emkzBMg7uXHNPWt6iLKxp/A88vJ5gCHAeQTo6fbSXnTpwzfdsCP6PaIwS
l3BkLf8liCSRobdOZG9pAxsDj8Ncekg0+U9ODerGznjAChzoFDfrc1u9MXFMCIC+
8CgABITgVJgcbJtZu8Mzta1th3OX30q2uvfWPLRkgh0FdEgntlnrKqtdWJGcYpzz
C5GKa+RPO3gIwLaL5fp9zjonm/tSq7pL5KzmVoBlwQtXNdOFL5Kbin67q+5vICeo
ZF83i4XuJgdGFOo7qKOcevpJTqpYSS+QfXQSwA2XEEpJVhlQFSEHog0Y5BytmOMB
1QLWKtbbfnbHhasSvHo2AHBGCecB6te8chjR1RXhByi9bLBPL82RZO88tyI7lMx1
2wqcdIuiQl1Cjqf1a80YmQ5PdBdPFV1nN5xdHIcGPk1GVPl+V5xUeZILL0ecQOpo
reCxep1dlUWF7CzD0RY9AIzsp6rH9LmyYIWKgeiBceIjjWsem8IaRfaaCSf3N7QT
sc/rndKDFmJY7OszuHXsdrtGHMx3EnnGMyXNQAGi1EqrZ7iuDhKCcF/GX0bO1B5U
u7RclkQV4pRLPn8HLHVCGXnw35FX3ej/R/idT02VDLd0XPuQ6ynvlzOPTGUJjdTk
XnmiQPPauRLBAUc71k1qLrDUeMvUGG0+ZuHFOX6E5P8gX4ewbiEOoY8eSkfyCR0t
nW/ftYwEbe/LlAloOBJgfZ7T/oX8givhyPPb6n2JzOLJE/CtcuuSNvlqWTcqQAMO
bex262NiICWLszD6MNET/N/EJWLE6aGP+NCvRq1zzcA4Uv+9WqAImPK9esagW43L
v5VwZW9KhpyLy/+Xibdd2+PtZqKMtEw8wJ8zHSa1DhV5qSync2SHDm/tftik8LTb
nz5B8dUh2/z9Cgh5GHcZCAuunbBFzisUteSe8iZiqOwXiv+/SkX6gOXKRm7l2oR1
MtMmEA8v4bsote5OhFGoXGE4iUBYqVwvn6HWsLYNb3Cwekg851Ago0mNlm4ogQLh
j5zPUJtALTUkCoRJ/mDaAe6JvKNMVY7TOWW8iMr7Yzy5RHPwhb/zQSG98t9haHoD
dNVVUYI6V7fKn7Fmnu/O7GwfOwmoRWWw/bovEldX6OSAgAsUnc8LFouO3+35uXDq
Gk4AYspnb6MYuBgNUHTtQ1wh2bso3t2sHPpGkb7pFO0oOiK7t0LSBg1PtGnPMeNw
TWPDRUqdhvgLEcK4ioMI0ifadotg1jXuS+xz/fZ/N/1Br1X84eZjuxlrtk7CEtLV
ZxNFXweWIRJvUNHYozvAEd6NByIRsaDgtqyzodDxyC205p1//fxNAPlDthdLwTEe
pgo6sj9VMv+zuTdydOmH4DeahefdsL1EhY0/eXoYM1Vth5BItvg4MlaLecjU+fsD
QKf9Yn510Rg7WVocbWkhcYFvEc2j6EoIuP8s9ZSjuc3oO8iSrb2ZVVzhTn815hiB
WTXYDliV+Y8zWwhpEZKfyZ8+vh3Nvr35VEQpLA7MaXrum3+1gz5YIUlCYoCG9TRi
XOVth3Mho4euKQ+n330vNpyZzKUlq6jyX68vXecItm70R7nDMGSM+JRSJcQCyOqT
k4Q0MJR6LTmIvmid2uF0OQnvRW3kZyZYBdmGiYjgIT6k66hAUOnMq9BTWYI/F1FT
pfOMoiIe6FY1UZcoxDB3OaY8Tw36L6RmkLpkctxiolG8kDYsfAqUWbpo9gv8xu5b
O0SXBIPk/r9GmI5WlFn1HUlQfgGloiMc2Zke3XbKZw8o1/Ji+soyAGjRT+3O3z7S
iM/JGzUxjojYq5LS4oiNNPR2HGtbBxjy/AlC+brGiAmXqCJNw5wcpGMZlrljsHyb
0poK99ycSYxFD05SbsHsy1v1u6rWJxrawGpraIV4Q1tGZEY6eTEPQ9HdQlY3rYV/
qnlWN87SHFmSv3Ye71Q7fM2XA2I2yz1vBSYE2lqy2hDYEyjST/7Fnz4n7na1Y1v/
wMQWNGVSQH0eI5MmXMM83+/17mmBWUV3B7hB9r4eto9U4vZLB0s0SawdZ2WNGQUL
HExlNm75pe10f353nQ2lwUYgELlB2Dg7yYq1P4VROZrTMsb7TUsZknmVHjllSine
+eahqATqPdEJ+emAeABAErinRusDjGhDmRooY92DSNVrxV6govVNBEcQs+/66nPG
NGaLXug30VvxH5UPoP2Sq/5oGaLsYWOgAfzITggvg/xLNT1kXeg4e58wC8tanSq5
rhRcRCnm5ayo6C4DPvkPIdmLM5FRX5KJCTvBem9kkzbNr4Ickj9BCnbutvkwVCRW
zrKzPGgI9CTmOOETflJ5C/5pX15a0ZYSpfpPchIFu9xnqwnWdPC2SY/FGMdF2T4A
qMQ2siKnP/Y1WzEv0V9j/XKbMXjUHOY2QvRcKvsH32cGFg22Dd0dAk2eDJe0263L
gYQSFMc+92OFnV8Jdb5/Ne+c7I2dlfqpVHNP8XAhTlV7Zi8S/xhIeq4BzMQkNQEN
Ys32xwQV0oAvMMoUuGM4j2BRcz+IceySOb4UXKjS1mqRKqKBkqxak1IQ/V2kfbZG
A66QxI3VExOCLuaw3T1UeF0NBHkiVeBLZSn7Zgne0KZsvInMTQSR6k2tlVJ13W7z
Xay/dye8ATnf5TYDgaYi6TBUMBWMO9UhyaNSgMPILTyrtwiT6FsPDWk1aQddDrFj
UORA+NQNAfPj6ko9vm6VEQAMYuC7VdkzvZS280duEeKIUmpsqYfA7ILlNEgltRuY
kLq8Ono3i9e/S5oT5jpaJGAmQMqe3RwivioiIdbgWL9e8FzpzNWgKE/nMNpl7XQc
AQECBQAepo+LkoARrp8TmJPQCJQcaxf9hYRkAtanErE4oIa5o8lwGpkG17owFEDL
lZXCHLCpRwCOmuR00vcm6j7b/AitZJsWGakN0joCqLLQ4DVG586N4G4Xipet0GF+
jSYDkwSbuPupQwTtGYqUjURqTrBNEA9BS7C18fvCZer3JViw6f/pkGDpVYpA1+Ys
7VW8GTM3DvnD/YzgyKjHHA9kJeNM152FCTXa7hRTHWRP7MqFfHsKbPEFo+/iHfbC
RZSbinT4N6OTHGQCw3M4nZsBgiMbpcwETXVFj6AWQ5BRs21PXSg+ylnq+raZXC5t
tq1kK7s5PqcLHSQwzfqQObPBxUsml8eg9cyRy/E/U6NkYjqKJiQhw5Hnc5H7Nyz5
XDAPeD7a87+Vkv2DUKWmCrkjAteGcXb4ZFMS847ScAiPOnWWus8EBtK2npt97Cn4
nYs+LRk3jrKqv0Iak2wKIAU2e98D1GqRS6HAL8fH568/NrDHtvppn5BmwwaToy4d
w79GasV8+jry//s/yaxv9LyHgVJ8Sk0fS/bwDpXkWCi6tFS0maxPTcmC+xNLom8k
x1ZoY/JlCN+4Ih6H18yzXR7hXoxR4oRuKCX//QM3C37Lx7d4lek87/cM0Nm0w5EU
4ALWha+d0kvAwrWFPC16qkmj+miMhTcx8kMI8IdgYSxpGGIz3l8Y+THynk151Cfc
PO0h291TMuKMcI3AJMkWf+PfrtkdioALz8IBcFcRUmx1zVHpOg46i1crO/XFMjvY
/ga3oNlTeHyXGbokiTgpkGAMRxatFkmCNIV2XU4hQmJjqvD0RSpgXNMMtiWmeqoj
xDxybQFfWt1u5CMPg6grItH5aynwlHWzs33LhFIMguA5JIBGO4daiGWHfCf0lato
6luZMJ+z/SHAfR5Jrkm8stYFaVmgIfOqOJuqz1/+DtUnuC2ldgKnWQYa7Lipll/v
4cqklq/ZQhx/oiETH6AzmuZt5BxynMXuPf4WrYdTqUMQKtoWnlktSTiAhslfHs9O
PThhLWL0jdqbTekh9P0BRCQmgQWTOUn+Fgi9kjE79TbdqIRHwvafwmOtxcG7OsAS
pQHNvodg7NSpN3KfI1426z/RN53bEdDK2eb9EbAD/u25WGaGKyfXjDgKGIh7Vcge
UiarOsIPUwRmucuZ8ihP6XNIMnhgOyQSb5pp9Z4zFM3EaGSVf8Vz/IllipB0hnVi
AQlOJ3NJvQ1SVwQNN0qZ7D5SL6vsaXoIBPx8uCiMnn4yXlBxt7AIQ5/lqAtpPpLr
mRs1cReBCBrCyNSatwV/3L9UlCHnXB3+g+o+gcHZhIfgK//8Aattj5PQu9zfm4eW
yw/R7tkxKpuWsYCFiJMFQzd0p8VsEppjxBVgedDhjwwQaTubnVpo/Tcqnbusv5y6
Qs2IeggX5ZxZ6YEbJB7uOBoszG95y24m/cpLmA5fF3xMc7CoGwYAH9SDSDpApx7x
xTE9SNfd/d+CMcV7LfFLG0uew08i9avmGVvEt0rlJUJeW4nzA6LS9NUsem2OzWE4
H8th+A9zGOk8jycatoYv3UGcSDKanmyZqswkZN7P5kVHnZko8ZhX5yezM5nPHMvF
aGwCwvRIb8phnQCceEdop69a5xsEDW9dfWSImG6rnEjOYmiIqYnTn0nS8ryKYaXE
qq+/5tgZNmy2CxihIo0hLvZFMFFvrP45CmS9l10sm8SYFwYC+smv3gazIpWZnB4q
9y6IHvA/ZWaEINSQzghgnX9XW6gBekOheSlbBKv8NzqVASvjUauwELvZNHgpDzN1
8TGPg3dgKWdju+8OweOqBCtlRuqQrXPv5DqJSys88witYOodJ8MmIm4b32csqPIY
eLC2vUpAD+AsGQjC2s+k7iDUlesCJr+j3IJMFbwY40h961bSZ9nlb3Hti0NUTdl2
/6MTYm4AV9uUF1ymh2V4CksdX4oZgKh/rrKXO7GL8MNzQOupKohCCKs47kWed/Fm
RJxBQFbkal50X76Jk+fZqrRusjWyTuUv8X7j6mg5BiPaVCHCMFkcy9N9R45g49/E
OkSglUH5m7XH9mQWp9qOZIN0uSOfXq+bHove2JOfQpVI07YuvJVP4jQBOxWoHA7e
iEVwT+P0vLO7gVQu6Krxx9W0SdU6d3ciia+k0W0NGwHwmosc6mU4h2Hf/QzskHKh
etVb0t7JKX6C+r1JgYgs6TMEtQQ4z853+PFoIZxQJjSiu3lxH5IPUBKuegS/ww8K
lELE8F7bg69xh6Ngq/T8/TkReQt2E3DZUmuwhi2OnXpKgOFjxEYufJcCtG5YtwuK
s7b0nLn1C/p5ggARjpzctuetW7onkBA79phd/TARTr9G+BLV9EJdylF9q+4HHkl7
fMkbRanwjWFaHC+aFEHCv1x14cGooPM0UhPecgoAtfurQis7Tp44GntHZEZoNvHm
goldSfoIwok47JKv5U83NqVk/I9qm1mxXCCcEs7mZtyFr2fACY/6cGxSdMpupiCI
XE3J2Fu05BtUDdcF3b9EOF8ZNtoGDoOwpGgIJ0axSGADCH9FrjhvMaSExtvt2GOB
G773h9ccdiVuqvhW0PCTDiA538iGAEX9JkITD+6wH8ro/S9fP9wYmganRAPYFNXw
45b1qQ+SZH7Hl7YOeMbTKFbcCGM7pKV+t1jQ7JbAt+kBoPNhbB3slHPYsFUt49NK
RjAp9d9BuwmEnhG4VjmgxLfE1ff/knIxhhA5SALx9wjhGndAyBJ2uOPIFsM2kAmB
RMDsBTifsbe2Vw40HlQgWrPKhaPw5arOTSsaUUwkGxXWbMitofEvngXnNUwThH/T
UiAz/PSyaOgetV64h/cr+8pmG6MrYyLQw/BC4aZRQvjRKTOXbDAJD2uMRAAH2VM0
rHefxRfBd1Ro9TjNYp+JQVvuDk0607Rb4ZlTaTEDGD9/mGarw/wEZA283DD7ajH1
5HcV4BjJkyBzmIj72sECpC1Vo/moLmoZ9Aikc+Xs5tZdyRhdXPbdpR7LnpwtKIn0
flaWsF8tedNE92NlVptW0583bSNto3EmWEhdO4CuJU0AUPcLaZE2VVjzd3ohvEXy
7WJuAQR7FdRhmEYPSD3PaaG+ICVKrMzdbZw1cCM8TjusVZiKSpLqpicEZwlX3dCN
3zhVVPwPNTNAS8CUnMQB+/GE+V56Omk7XuyDU4b1FAmdr/N7Q313tfrVtRynwwKz
9ZII/xyzBtAssEsrFQoyiFQOazVH+ZRkmzxAhSVL1eJRHYuiRDXBRvHGpebes0nu
n0Dxd0kvWuXujs7LNzv4oBzmkxqeKwKvB8cysHVof7W+yYKGvKUjoWxUNbMOazxC
viCupLpB2bPJrt9A7Ab4YkrH9TLqsfdU5qu6DIrD8Rd27xLLaukNBw7r49D34fau
1LBABhoeT0tGEWOTaEIAhymJGt2utlcj2A2y993+yVDkagmCQpAwpm6lM0HbG+u+
V2zm8mhncInMzLpajVyPAWFIyaIdw1X9pFwEqmtB0JZPtntT/Ac4IB0JITz1H/27
IbxV3is8+mTetk1DcKplOGM5fpctG9zhOjDloMT1BTtZ4W3OT0VJJockqjNgsWwn
6Mw0OC3/+VhVQw2PV1GL/bd8kULp0eqLkFoEWCjsF2JldQMDdeeDIPm4EPRulDkk
4d4P9LeGHx4NXQBXr8c+PNId1soMpAzEG2DehMp39IptvKq0odofsqHD28188fbV
BRq1300ZTov60AhrCjsh9g0WDcy3eRmWBV4DuZz/oZblbk3omFc8q8Z0cAMHLlXS
OAxB8RCBmt2VvrLg9zV3HfSCJ4GdjnxYFZyAFV/d54xPuGSYl+DcpPsPbLHR+KN5
+TLWM/XVEOSuMWZiLhYSJi13qwsXRs7atPnAMaz4T2DXxbvKr44TrGSoEMS2Qcwg
qt42Z5RsZ4kK2//zKRSrPRATm4Q5zndr2AKlxvchASL1x6gnDl2skZLcslSH2N75
+NhFL8pMPDRB7NLB0ZpCCpN7WtpBMnDRIlcijnQ55zQEFqny6a+POzK0SdP5HEJH
myAY92v/ikO4UzaZEUjFtwvz7MaJM19CkRwmaXUlTvh9igQY5U61Tl7tCA7nQHZW
gqjn2Nyji4MBYDZk9TW2NX7wuR+xlvcwLRPT5eheNNNaWq4C+ezvQR2sast0Q3dL
w21Ik4PPXVg0ho3RqmJILzRDuOhrLagzEPuUNBdhrNmeOoSKuiQUkD2nJ/i7dJ5p
6pTcCLxtNCJKO7VTdjJCaNFKVimpB3IQm6TRvKdnXDqgSyLbNCj6wFOknB4RZhD4
o3ZjSsRUQhVTx9Q/T240/tc/09HcBOrJWfpbPYghbkYdTKUDPHmgHuv8d7TJOxaR
RQw3H4XJ4stVHwOkO4jpft3CNFvKMyJBEKi9Dt0SMAbm86w615TVZ5+iEHlxtbEe
a7anxX/gJ97DA4hjCeaU55xWlrdHAo438D9NyA424Q1r4ix0xu3XloGrJnHeMPIw
/jG3FYCv5ZUXktqWgpSoQ1JWM8RaTpa1Rm9Z7NjcK+yxZK0+5KOAco/NkyB8uyTl
SWlCRmUIJfmT5bMmcr5wuFcGJ5TsCAhh1SxJPRuOJr4rBlDGbpXMa5M2oRsi5Uvc
Rl/iCJO1djVBEE0kW78kDx9ChvkeNVbKVSSMWrGlnISXRsezEqXJG/ROLUElhbKH
c7MPDdyZgy7kFsYBzGpNcpSE/Yls1MmHhcdcNeSb1iZ2wjV3G6qB7WNjoHwv5FtM
vJDfnNnuQqM05UAri+eoLlT6gonLsHIEY1RBuXoODmKiC6Aa9kLWonbUsOIAbC7b
ElohfxOkWJ3R2zlwUy5VdAKJh94cHymEputVFr4r59t6occqFvQEv0L5i3ykdGDU
YT/sugLPosTsw3FYPO0g82VAhvLUb8MNswO4ptstTEwug6EdP/hvIBw7NmAPoQ5k
7Ijx1xUjvs8xExEXnvLUm3NTNGkSdJ6rEvjyI9C1eTW0JZyWnjs2jVtss1vPD4Ga
53G5RqtVEexXqy8CnRwOsCE6EtZ32Bl6oq99+LV22J6ZELZS5PfG6kF3y2kAp3sm
fYOeNRzru34jCVHpaCxuBgTqxXOjMbuI663kgg2FwMLefggUdfLB9Ow/npr3oZ3U
9GBNdhAqwd3F3bEF5j1AY7Waeok5EUYFfTvhUg1+/vFtDp5Ue5oisGkvl7A81ukn
Ei9S7x7mC2j7iuvyJFJrRazLQe+/IWum9UHsoGPsWJzP6ZC6jcMQAT+quTKIK249
OdWvzN7BleYcjhpZ9jz69Tu3zJvVVXXs31oFDVG+6mb5Vn18N4jWmD095+2DrLlE
TGUS9McI76D4Cf/9VaDBSW/8UVWcfYXF0q/E2wv8kRN4oiE+oUWGNbXVWIqB4Z4W
36XEDX36Jk1F5QX2Q1B2dmg1Lktdls2eJ0hbbcn8C2/8+8QNGLKvYNHJWC2/MZIG
yS3P93Y71PJaz3Ofmg98225wCm13p2i9XoquClJLYmQ1kcCmGqUnggJdyT22oYMx
YgOj9M8QK4Bu1wIWsUJ5fZAJq68i6bIK/LpLBXSWe2bwlzI6jWCGbGiqoshaKNHf
UctgL5TO1uye+VHlJOV8i1/HwkYbs/S8H+LnbB6HGKXWSnJ9BVaVnqT1KDfHj4C3
gpEtvRMM81Waq+owAGn62yxaIpQsVyxU4atLk844d+Fjwg72QGfS7ZXpr36o1Gzv
eagxWZbP4v6faCAS9xUkpYoR5XenRoCGU6tMZGAW5VcNQpB2n9iDkSevK5v6mcsA
OkcBX1esB4+uAbynnOfcbDcixK/v0qOxD2f20OIfP8CX0ciy2riD3WYWayjAlDBT
UD9USh7MTGl729sXnRV0Ot1TADxTycSdlpMLxp6NgQDPDq5aJDoH85qIwHTa8QpY
6flmx/yjz5TuYS1FzVNdRh3Ml2fGXPHsnooJCTR2jscHB75MYVdZdihzpeE/ItwK
ydRUH783Do4bjIMs1AkGuQJYhs6015eotWvi6aoqzPJpDVF7l19bc3G+U7jETLsb
VDTNmHYpkKdeglZW6qQugOMJIYSdnUL4pu7Fqz5lhBkQTNoky5XBDbdC3V7c6Ysl
J/lvpiv2xa2SSq+txT3ByeTlZ/XMTRuo9uaWTHpHVnuQ1dFH1WoRACgmvil7S8Dz
dFFw0DrTgvnpg8KtY9gAvJ/RyyaqftNJ8HDjLexSEvZtNiUZMyVjlawqv3HArglv
m46MZ8TWAHBTIyzSdWvxKVfF4/SDnyvUrYWij5jAUfei+oD1e1l5xiDEKu0K3OlW
l13uiJu0hxlq4wmdxNlb9hf+zcDymYDwgLeJfYVLanZ9RwqFjIskOv4dVFJGxz+l
h7WAJFmQlN6BEe7yn+v8yH0WmoaTwU6Cyz8hi/jZkpW+RPlzvx+mgtdWBRCdrQL6
ZM3LVXeWPNeRkqSnhsMZ1q7hwbYAiqvkmA8z4gTxYTcy+64CBObFTmjU3OkOZBHG
MZvMSYE8gDIXiyDwHuHpjySSBiDYaTPCJ9iPXUJDGPxHg1xElO2wSsJC6uEZt7Lr
KJt4XYH50raAMxD2mqo3Xu+ELsUf5M1yagWGu4BSFamatNcoD3GGZRc/jBI7+L82
qX8WZXBAMxGk9ii/D7K0QK/3+McJ0/ZTdF8XxNvA8i3Aa4oMimdzkYLr/gRVKggo
FqIALiH8vvMG0LTbmmPWmkeqkhhsoBYsKD5dFJ65WHmnug9pSi6GPFwN6PZqPtb0
ROboy9ISekK/vBeVd3zzenTsi/v/XWnSehW5RiCOnh3qBU/YcnVnLpQxdk71IUsd
MECOraJsIvsjxGODzOy6gwDV2ouXRh3/6Sj9B8Od6Mq6KmnWRkIyqtaIllsYYlvm
TYENSIt0P0v/E/ciuXcv3TKq8Ui1fcPGFbxC2peUqyz9w8P6K+7avgBiwvrsr7CR
ZNMqmgUe3eJBaskWlXYi8M2yOS5nuBjRSbegle1Z44k7XZ/qchZ7nZiiIlI2M/Dh
6Ayb36Q+YP4JC/0tN7wpV2pCs093PiPEJR8JRH3/ov975j6eM0owz+UYtyMX9yIr
oDd+dMlGw6DhZPkLy+79FX3oAqWKqZ3TpjjhJZKLxszPEnNlx9iDXvpEm0sBUl+n
lHYe1eU39tyuSgprNwephnWDOgXKjYnQeqHTDpJhKgd5NiIe977lLQ4IQdXwvcH2
I61d5LEiFEjibRN169chopuJ8lnPiwjtjBl9aAtRm48Pty6LG4W4879nJ8mX1Coc
uJxWY1Cgxg7HRykMcrVhwbPaZwQpnCid536H6mm603CgE2masJfYSyHPcNkCABIC
OWK8U8IUd/xCg/Su5by/rkxaVO6DbdyRdFk4oxqR0Wm2YAcV9NIjdYXvu+fQXAy4
hT9D9l6R+LrH/22WMI7wXt5urJtKhxI+UQ9lchmlsnIVGksLHaRM6pBqytJNoRuO
TOl0lH6Qq6cCBPuvi7vv2NpNW4kgDXfZNL/A5CHA51J+EHsKquiV73mvpTWTzXWV
va9Elvhg//1nl9kASnKpmGnoatDyJ4mei7xGufgueTDrCZCz3oRqHTaIHQOJlxEi
IzQPSUojRXF1ssM366571hArObAT7rXFTto6hcqj4gw+xA8dtB61ZQ5sqtNUPrRl
KhIHP+zm2xZujD2JJ9pEsLxGBLehdS5SqB0ED2++af3yyLgt/z1O+1+6Pypn63Nq
2L/VMiaESe7jjFiBIQliE65tAAoSOK9LjfOQR6n7uE5RgguRnQofNfbXHvKuwi4m
tRD/Mrt0mmyxt1sT6zjV4ZVorD8A5rItLRps1BBjfnXcj/E8DWHM8T4Ux/VstSAv
1noov7X/6tX50m7YQaHLnLxfFJTLyKCog7E90EK6JrQPtiy0vZv5mylHVNYI38PF
qjX+5NXM6AZSPRJXj/AE3oJeLKdEyw8gjcjryHKFHIT1oES90mE/ZzhxveT9EvdP
8lTL1yJ3UJ+iabpMSiw6aXi+lbrxWgFhu/HpTyUn9wHLYDYphzTrOHJOkeEMjcJk
m5h8umxVc7EYCdzQuoH+3gofhMtB+ksqqlSwzJIskfyu2RGyGHlPh5uwggE1Jx1z
TtAeEF+NvDM/znZr7LHPIWOG1h5ah/KvNoYWLdyNTMdLfmL03DO2ay665GMqRBBZ
YEgso9w0c8yxSpbApnYOcxW5qxl1SeRAgG6xJwWPHCgaoLeiAvYo1ReRFfQrgljR
1i57OKoMAXp2wRrd0A0+MbmdSQYqqqVLSM9hIhsqDnVU5faVtmE3f4ChWGXyxARh
4qtegFoBwwETDbfLtx7gdKuTBU/+EVUyUa5PywVo9N3s/7urc2V2phZQNSCD2XGH
6zpcsUb2rfRVJGPIBRGQNDvw6TPby61aGfv8NdO7MTx3PLTt7hpTOIgVb7GeUVEM
dl26uQ5DcuoeQrVQF6OvN3ah80i5Jue+ER5a5gyVy6++KudDXSQlZoYOdC5jk4XG
kw5ko9iAyQag+xnGOu7S9GJv6RmiUfn298Nw4t9fcxbJ9EVh+8bopNLZyM1BGXnq
0g0RT+2zj0QAovAxgbhfTQJ76kp78tE/mTamn2rA7Afy+CKvfYbZZvdmFwo2hqQ4
s7du9JH7hT3Pnmw+DaGPM+3vU1udnLNdO/BiX0GhF0AQnBoCc/VYQ/vtAaSLOJsZ
R7OswiZn6I8wiDx4f1KwC18Gl7NuYEN4Yrecoy5alCFGR1tEpcmzQC0+vxnUC3Hi
SHLLhRcmga4kUUr+Qge3cggkDQ0KLYYWWs95uVOpr4z+aZQi1lVpeR/AcDaQsKp+
1LApWAUrAPawcIzItzuKjfXXwkBl0IGsCIQc1fRBdnv+35IJKY/x85nfRrW3I6lh
wjZPQ0PRXYqM+Icb89pOQoiVkK3jjhoEXVI2s8zyXWayPJ68rWFq5yNfuIurWTOz
g41FsRy/J8i3ZDSl3fmZrCLxUTM7JJtgxg9g5DaMukEaNQRceujulxMSv55r3KeM
bW/xrIUqccGFLAzdGlOcVvTGZkrB1rA64QFVw3QX3+rLP9ziMDrZ2ZCHUG2WsIjE
bMrlWMn6/0Bs+ABZi1O4tNokpFPUFrf0ybOw2juETMzHOEGqCZvLQkQwm5UymYNX
s1cUJUcvqwJb6V1Pd3RP4zLpxN/o9ntgyABNr4br1i067y/eKjktS7/x8M1J8vGR
8mDV7sBDM7iZyYQMZ2tFov25V9E2HmGgK4IzP3CfPdENq0SPcJATMTsVDDqzv0V6
E0flHevbfrHOKASLPsfE1BZ69T+Jk4sLqWRVD1P5xXlXSwt3uF7xZ5LUwqmpovx6
MTl3zyAmmKq9R1hRz2Q73wc0UO7F8GvkLXaR+d4yDHqIvKg8I6lJSARumy+gnq89
1cjGUvItj9fXZ/wkiYu6iDTN3djOCj2uCigPgWLI2Gcmd/t0OZTFs+NVmtsLHpVg
kGPKYupNyvhZL0MNlC8mtp50slkO38qijDFbd4AJuV+hW74dlRz+KYgsEi7jwKXA
54QHvCotgX1BlotUgQFxxoQpYicuDA/IgpnLirdXeqlVJiZi9Tl3QEM6iWXYr5GY
aHM+RN8qNW9hDeXcUqn6m+fazvFcTD6WGuop6g8epjOJQeOQBc1or4QWlZ4KTBRv
Rz32+/yQqibXOQACksKvMLYUj4GZYpqN0+fxgwaGIVVilO7fm0UZ9ksU0FM0iFI3
Q6uJcBf0m0uJbaCXc3t8nAANvIukKIdAWd2ikSXy5G7XVCKUbK3USSeH9TcgLm0k
uefAbuSlOEOsdteJWIwj+7lMoLN0+CM4R7nnODQuwtzWp0Nv0Ya/ScdFND8puVbK
vrDYB8fphe3F6rmCz2EIjV5qt3TIG03y1IylG9ZKSAas+i1Zk47gO3oH43gfz8mK
H/odKe3fFlGQizNwqaY0Lk4cMNgxQQfM82DJ382Wb2omnFSKlu14Hg3IrsjbBQpf
Ty9DtCLuBfMXsTzgcyiT/adP74JvwPL9p0lOQXB1CVic0/D7PnxMvO+Uj1pgfr9d
/P1zMOlevGQsTVW+GEm+sncpTmcwdf3D5VMDZn6SkEXBVWpBuWoUW+Ij+YlX68LC
i10BAYQHBO/e0ekatHAkqZZdI0PtjsEx3pAzAgvCm3vsHM8W7T1GuiEVYqIdTKfn
cx+EAX4QjN7x7iLKRQYHTwcPlsiLuWsJmtbHmIyvK6gUVNA6NbiyW9iHEL4GAjaI
FdX2+pTNTM6zT5MOqjE86QuTkiPNDdZnzafWHNwSiYs73KhiFujooaFs1XlfSwRj
tZ7TaDyNNJl8/KSAXbT0WGZdaWJg6M+DlAbFCZw6+ssbQAbi1MM+T2NWPLBoLhzi
b/2/X339ij/3HFe84KNOEqpYZ6nkM+FOozoFwJr1GzIbS3g1ZwPLJTxiUfKsV+Eb
S0nnVHAR7bh77JXVd4CtPzdm2QLX0gdd4+xzxNAfrASW+cBncjzDMgjsPvBPYx3X
PFQrQ1WpS3a/OoevfWF49soszuQ8cSs5iLZ4+TrgkwbUiVmDO6RrUtKZaJAJFiws
BVGvbnUeQ45CV3TNY1IDNTWlZQMf3xSOh2xcoGilb3P4Kxg9Il/f4AoZ8Dh1PYtr
ORHdse0AJUGDuMVEfap5qbw47lBbnoBJfotudfhL9tk8IR6R/pDx+FKmZ0p6h9F7
v72Qk/RKsbQmaQOI2WA5DX7xq0VU+6KwZFUzNdR/hW/l9jORGA2n0kZ/TV9KEYm9
YIkqg/CGavq8hy1Ray2hkko+MxJn1+OVgNU3yuFFnW8h/gyaxVoh59e3tOl+XEnY
Vfi2ROSuF4tTeKVThKR09f3wkxNYuzOUw7wtI8bi2xKT0LWkXdG/I0RxxptCcCY+
uTfq6Ai1vgIqrQAEtzJRsOvBb9zkEixub2uOotyUb/rMQdxhkPuSv9q5i4rgs6Uj
M6Z6xnJ2U3j+364adfBRoKVAnA1NOidJFQRzpWZMzm2qjqWX4dI60UF+4FbEpV0l
gK3IR88hFpyvzqFsy1fcO90O2O8FkFXIHpKsbMAvio46DoTRWIVdTLC4AfUZRd3K
mSh/yCf3IXiKMz+Y8um9mxjM835+MKQy8QGywMmslTgDKhUP5LLAefxYven3UNbp
j4SNOle8V3VBqe4O6yuoR2/+KiMWBO20qZ+38HyXc+/M9zTJwbVV9PaLI8Bk+KDq
FQDUcVHZvlIs5XRVxMPKMTMpihQTA4ncyd40ODfp821O/K9aCpAycTOOXJQgO6Ns
LH+A+8JIYYF822cRc27xWkqRCRX/FARVmqEGJgy+C/NPYrt8ItWKIWnUKCW/Mcv3
19Cl6LW60yzjGYmEkUo259+bheWNL0dfjlUSwUK73oDQ9VC8OH1mIsOneDHoCLFW
ybkBPnXuV8PHQ6mnNJ4CzCKpgG7pEXMOk1HdMDjhS7gxuI423JfjflqtmNr2IAsv
8Z9BG+dVSw5uImPaBArhhgwFrHEwacipTlOG1yJWhhK5SqJHVKQeBa8l6+irDUlD
7F+oYX45QmdBsMzHpngnfPmekxmQNzkpUlOru5kPb6Hdukd9pSQmG/9AjnKcJj4R
INz4Jx5H9DRGeIr0W8nft5z41bUZqpuSpEHVOMwmLw7EnlZEkPyRaNaMo8WFqc5k
v3fzGfeZLBMeip4i9eNG6Ha7IwlNHKvT4+PuEk2DcXdsYzdLzNB06TbVgxCAD3An
W6ABvgSb7gQPHEbUnkcYBLHP7uEVCRUt/a+2XVho63cWxbHO8Rqp0Y/hNdVDpu3I
YEoeW/K3h3MDYmooz9Mith+YpF2u7plKWpgt7ce936ekNlhuj5g/vnRrIYxlPES5
5L4XzokFX5ipEKHkkIHR3j797JZgHpomqPP6CPu/XZD0kk6rQ4A/Bv40BH48hHVd
4y3UqTK1BMQp+KzLuUXBJWez14gcIvxsOXdpSYXhUq06rRGQFLeeyD4jlkxGL1Rj
UEF52PjukVISbnfaBtrGGqkUCfiQGmLrnB4s6zwWGsqMODjsl0N3jjaEvkcjDCwG
OmhIIuHpUQAqH73LFhkv6ov3E07/BLokYUkoXFjDYbO6ZdkFFbgWyFHbx92xa8pT
4moIb0sluTv849tUyDhxhANe1VtYNV+EaBUtL7J+ZUrBl8gnJAuAaDRb+3fPNsmT
fJcDJZqJebvY4lYaGgk26L4qRb/sveawNaLKvxvYnAU4xZe+/TjHfocb+MtE2lwS
5B8sgLzx34DPKMT5EMphugZP72aKmeBEQygd0jDh7KiZYwvasXuXwepKIDl0Kzm9
D8deQAOHk0qhnkH75eQmIPUrS7XTpuw+WtTP2iVWpdvUDkYuojjm34P4VAFE3QcO
tO8+FHwYvj0VKjICj82XyiVeyUL3ETBWb1z4NCQWQblPz9a27vu5P1JdGbwLwFBf
O1hcRzqeSJnuQs3/PZ00vnxjx0mRQ/hrs3VqPLesRR5Y6owqrvNHyfPWYoEu040M
1ZEBQ9oNDjNUBmt5RLo2FBHPcX1TFWMkrWP2fkFOa+CKHJziKg4A6i65w07XPocm
ndzC0l8JwvsEeZWngrM4yHOQN3V17nF+xslbxH80yalvv9orXymimlsA4bZ30PtO
roGpYg7HFnJqwPxQvV9oBDr91poFTYu0E9OqjN/VaPPDFI06yiZO7UvZyfBiotUy
f26YqTdjRZt4erKjWvd1e93TjDzHP7/t7o8xgE5yclNEAjKeVYcRiKdo3KiVBTrt
eNRSCC1f1Xg37pdQ9/6p/DqZ56TKhsikmlKR7wMIzgCQpszm2ntdaRGc/2m/+EHk
1rqBzLgJ/0YeGKb/dy6hNXbjgM9n3dtsnqV28E9jZtWv93Lsfgv9OFklY4JMe+CU
vQrY4lOhxGorqXSIMGNmjnLghyqmlZwPEQQ+jdLoxO9Brcpa/fwZ+i3J2rA0rRPw
84KU7nMPGlm1oQLuJPkes1iLCIOWG79WZjFPqTocjnho7oARhVA6cjqWQbqeXoE1
bKjm1kQk1GY3Qu4dhzVCqMsoSh+7DSWfq4qRVdNjP+bM2CNHMd606pAurh87mj+o
lq2pM0D3YX+oBoh5E0ReTfA0jEjKImoJLCix7UVorCAfa7zk6K5TumK1j2yaI+r7
2nghLmaX9qQmFP+2UewHpfelWx0pZUvXsJW+/61fotyyQCRJjAy/GzKssoGUCnJ6
aKUd0OC1BsBFJsJppeffcGPlBDmJkcJ7ETEXo/ZSE2rgpUvsI3oWMUuXGKHAlvus
JJW4iercdiGABW8iSWRrCw7V7TXuhy/7d7lm84q1cLEUXcoa1oWItQ7Fye5K8eL+
eEFdogIGhwigmdMTyIuWHT9l5n2mzvY4I9AZ6l5NYAkVwG43oRx2Eb7+ZojSVjjx
aVKo/582CAdO1Z86tUO5S+UFfvf7G6qMwyBRTEMTJNMBaWBHE5HAEJixH5i1F+mj
XUWbR3gLRvqP2hrHwonDxd0pWVv0AlgHD0RWpp0qqJkAIpWXiDqASK17sPtw4qRN
YQNf3h1MgTza3MSC8ZYcIw7Khhv9QdgHwzJV0GJ/D270NxLz82UP0xqWpsGT/MwD
EXi3ZKllRGZy9bZCtRg+xnHAjzeW/1xnI4Xm3PY3oUMLKffzKcOB8qGRkLEF6cUQ
MsJo4s4KAvp1IvtPh/yvhohlh3qJKkd61Oxs51zNgSc+2Aq745LKWaR+goMjDiUh
SiW3hJnVIDNnmNqJo2sRW/6qmwLbfRGqbIvJfexPDdJqHLfE2C9u5FaSuxAJgL+U
tONcQL93MTKTSbme6bL5OH1T5weSUJ7DRbcoMGq/YmyNaPBHxZWBzopI+R9AA1n0
oQlPaWIKtRVtRLlnFgWuiT32BAIRCrl2IIY6FxVaO1wHbHaFjZQjzvc3sUPuyS3y
gwbFMtw8kMgQjFhbFkc7+Kn5RDo3EBFYqNl3qqzGy1IkIp8kJqorsiSjOKdjw9K1
vERqElnVYkQM1TBxZIfadlUxQWfhOjZBoRdKOCveBd7sz+vf/nS7J0BMIrk9BSNT
ENexR5XHdWMOLa3dBoEHFwnn5X6KMbSh08QGPL55ZCGuQ2hf8JT5/b9Q0zzcu5aJ
C+c6MEmfbiaI39/4uHWdwS5IG3wJt09gYZIGfI6A3n86a8JHIxmK7eqhEU0KOG/6
OgkOadWkF/xJS6zlA291XUAB6oSEhEosLJMO3/OXtnGBWTatOkzYUXA/olX2Bq21
cyWTwXDnXELhI9oyQILLIHKPU1SPFUVicAsrRJgxwKaOj1XwFac7waSSRVVvfhZ9
A+hPaALENwopl9fDu/HEC02BmVWQ/Kv0v/csgBYLYQlcdCNYAW3L4UGwzr2HGyl+
otvLzmND4Dlnpr4R0rT+WpNj3M5OF4GS7aHU5DcduAllep1GlQujW8Cdj6MM7dDl
yu7XFEd1QvhVMigWjY9QDwYoSY8h0jr44OzotxRiYi160/5UVx3V9TssX+SgYGK5
RJUPEaz+YgcIroMFwc3A8rwxRLe3mbntAqLEG7BPHgRqXr7Psq55+p0R6tjaeSGQ
NOtiTrdKeocVcYDRB9PvQkMUSepUKs+ywxSUu/Q0dUwLv0PdsSUTrqh53Qeh0EUf
6lEQKys/ogLBSxV4eUCf+euoSaOEElcW9p/bNCqLf0RWLjGliznG+CkvnT4SyU83
6KqXawvCLnscZbVgmeBsPFq7CghHQC3+5wpF8TL9T3KuzSt8dJH5Y8eQo5ypGw8V
ooAuflZhc02SYSxQOkOuFqXh4UlqkH7QpwdRcQQGfzyM7BnFQJq0JgeKdlLFL0YH
K4p+Yx6omCIT+7GxEihOScm/naY6OXpfx9LBDDy5MOw365xqJ2wyZiIFIS7cmjRU
NiEW5LBVVDQPYBvS56nSyYxs1nEjQpK26ze9CMX7GNZAB+es/bwp12vQhPFNXsR1
hyti5Ph2AEEz5PWhfVYpMvTIoNhvNzP7HoinHEWRuiMwsFy09cEw8NktwVeKAzcH
UFxaGJTYUH6YJhRP3qt+DOUkvQocKqazFy2+5ujNoMfylI8N7joAdGpQL3YcTKAN
ZgmctFoh8dTwUYinb7qzZuGSS8OUGpjTt464fAlZl/JxW/4x/lO0CS3ZFojYUvHL
NyOGpbvV2sQX9rsoZHX2WpZWqZOqDGCEY74NlhO8TuhUU5h+o1eLDyCB6HSBZz6Z
Z3MJmGuDhfP6o16WKFK4wcE/KKh4xN7T9OgSNQ5yRilwENB0ZOmgJrJXbC6p+B2R
vcWdz/NZ+kTE0Ijbijviljfnz8wIqCUztsMJiz4pgcoAZQW7A6AnRRyZEDF0jb97
6cnKt2jM03pj5U5JOxeRLzF29XOTj1ZvT+OBA9RhFI3DXZ5+fGVoxShRgm9knMuo
LaI0r9xvtpf1SqlJ2HxyVKTMuNGQ3FSE69xKBJ3LOYAYLg4dRR45VECzT3WiqtIC
jswAGpmJEk9Um2fM2VzxEqpW/8Vxm8Pi3ZF31rWGDuWUrGdrxgZjwyDiAqtT1DVO
Ds3Ctq2nYREPM9Rr/urtwgKzPO08MB1BuaHG9YAwcbhtnD8abJvREl+1k0NW4MyM
9lJD2yuWPTZ6ZyAhmCQ2KlKR3t43QwrLRuzMb6GKsc/N0rwW3R1LzSWkrcCyWrV0
amW16ZB44/qnp53a+iWvAp0AwyAg6VyVaOyON1yHZ0gDX8R+T8PCWYvKNy0UoLnk
2Ei05oKejf2pbE3mBvlxOp6CzymltW7wc18aJjPe390iJbGUh/cf/z/U4yZhWQa8
b4vHmHXYFSokbOtwYhMjHf6SCkL7SGNraR+tkM9OSQr8R2525sCt0SjAwzUyvSow
5CFcbtkJLRSSGL2KmWzLyUGApfuTlngBqLXLhX96RW7nWxWs/aYKtF54EERYWugP
4J/n73p6OSzaSPWlNDlgAY/Z3aHcdIaFKHITWeL2biY2a35HII/jxs9mjZDOMl1L
ko5ZesiT+JlEhiikz1DN91fFNMTHzTSltEMDosNGEVMEqTVycr+Fod6KzWcLjmtu
wCrq/5WLtj3n05VYPvL/rmbTKAKcJmOlPkk5bsvtByl1MdT0H9L9lyz/F6lkcJ4N
JPnhgbNqQYZrMnVbzEMHRndwIIUdXzCkwFjzEmsRvnwBepktdbJlpROvU8HqjVcb
6qR//NHW0rCJwgKkpqdr4OlLQJrhW1zuXbi7SNYiw/pLrCVd+3RDRYvLwXV/r5ry
7L7kG3eHw4FcFWojabsDRpZzTOITP0VygLjpYgG1/qg5mgCTnrREAkxExVrm0Xhq
+TaE34Lz7xYItoM4/Z6mKHUzvqAeiDxbjEYSPlzv09rgjxMLSdSRBsnEP7VYKAaq
42TxDUx50raoL0wMvMCeGlGMGs3JNPX76yMa2ajIduEEf/iVTPdNpf5m+53w2Dpe
kgqEi1XXfdHOErjU41NHDsk8cH9xj41aUbwzYig9p/Ir0jZ2p6hL1TN/unt9O38D
xwUkW0llVyBsmmhnvmAEUEWPsSJlZeh6W3kFonVQhOxxtYMjvqTtHp37BIBdwQRn
SW3UhgaDLgxzD0knFhlXOePl4/i9n2wAyzKrtGo4S9uQEM3G6BzsbEZQcNyild+o
Sp8Hc5I21QmUUckSIGCohlVbkf0+MoY6o7Y73iLFpOVpYblSbbfTb5OuWbSEdEwJ
toXtRCc8ABBCqoU/Vo8nVKCuYTu4aTFV/Nu9Xi/NU9Aoja7e2Hqe+iEC9mEhUISb
/A47td6U9ZPKgN1bkTo5Ehav/lJvNVIKgLXr3e1qZ+eTlwoolezDCKpO+poUDDyj
7G4KrEPmlpvxmKLoCr8zYDreQUCbXquXemz+g5vzj961nXkXGM+Ff4dGZRFK7XIq
lCeDukPhfF9HtCXRMGJGubQD+uhcnahTsvxNQn/wsIn0MMqPFgiYVKB7CbvZrBCE
66XsN5pZK0jYzGa6GwLiGPjVwRxDuN52J5mPMZAAjRvPU3GlEr7w2e94I3XhT0Kf
m3ZxDDNkm+y7IUL0S+ur02ICC+ZvdxnrPYieUjWd3KH/XD+IS5R3bk1F/9S0YXkK
CgLQ1cKcijIjVf3EbkCJjD1C1u9BjfQE6Y077TpPB4gCjxqI4BAJy18gUQwfKkMA
0sD9bmAd0NCZP6U2z3rVEEQFh0MOSNTDlen0ywi9sUSHseKDIS7Fp0OFI6h+V1G2
VFV1jGlnueNZ4KHaiiqNh8wzWPc3z/RlGS3ESCuZxg9ORNl57uXkVTVPiZPBUD2Z
UfHLgsanN618QucWp1H3YHQc4Pbgy6YhPBOWgEnw/+pFP7cfCDJWdZW2N8J1GLkG
l4Qu4xTtbIGhrpULbCq871mqiucVVkSvNxFdxyi8nrr4mEWfRDx79yv+dvjDY+ue
DMhKQ4pUO18cx11/MGFx8nFiQ2eBOImXDX3yo2RxkrO7hLYvT2gdWh+5OjaNLvwl
6AuI00dz7pTpiP3spzeoMy8fbi4LCElSTivAZbA1/oXcgUKBkHADetVPMckaULMd
NN4nHy4hk+WdlvSkwg/3veL5Hl0WkQ0Agwj8IqfDjAI+Sqj9+uCJF9aSGh0Ft6lL
htuZxQWZoLehpvLYBCfL4YX9AGDq87xYItHBMdOzEtm+W+IcNdzppQh9uS2a3bbh
qxdA6MIgpTaqFD9X7IAkwpN/5NXbcfctzmBlmbKKK9F+lxLnaqJrUzjsEfWleesA
UCHnM8IUP5gEMbV7QNdxkZRBNieQHWy+BLlQoE4v2J9Cs4LdtOGZL4YxLdTKopOL
Rm8nhj1dVeugOQzbtxW/rUz7eNg8PYHPxQT3ik5NReTMJ/SYQMPinT18TRxFHys2
28xvbSeMnjwbcyQ9EM3Q5zkkep3OizRBFy22lLR+I+BokVNU9f1C0rsext/PhSsn
9f90asf7SaFhryk2TFcZ9tyJHfzVXLlaidjqIdaujlvDoMCfwZCtYHHcBghaiN34
wPqYQCVxt1fS00GCJCtl7m9jxnJgYZOb2p9Wh53UUNlAJ0pTborKbrLlQisT4rhT
WXen/uESozVIAtD5O/28DFCNfLdL08gqXeE0syZ9BonMOoghO5tlt6dVgDU/2ZuG
G5IWxeCISqHZ9p/ZFDdPgKKlQ6TqRA0eJrSy0oSGpCJx5/binAupwPDAEACiGIN1
OtiHTgFdCTpAtZaLIITxyCues7WHf999UCmsRXDaYkFGHtqoPeHXR9LhndXVAwNM
6r0Oc1xhXeZKcKZqiU5Jz3a5WMSJ+GsN3pESl9zpktA7pYUxAY3n0w9eqSLfn37B
aWBXGqx7rCAktgF2UXdJYKOxSFCmc9rRkJ7/IVKlHrzzwe183hCDtK0BjM6V1B+N
jhMCgDG6VufbPZIZSen0rE+L94C0Z3Fz+af9M9zyr0z5EzmETkT9eqEKX4w0ajrg
7YJOndij3zbVkHKnyg3SN0hF3f8XuKkpRI9atfnmWvNKLNoxGappFW7QCTEuODNl
6Bz4TjZ0fcLREfom2YaWnNlnlDhXKgAi8W1Z0UPBbbX0R7DyMIdVrQ/TNtMBxFVC
+GNfCEN9Nn1Xbs4Nt7JW1R2+FqEVf/gwFB0xpRb96s8WxDcx3aIcgjP8i/UOPWaG
7Anzd73rRGT3cHl/K5iTZzZXurWrCl+koOXTlXjZE1XDFqRdiQZTMUic9yTVQVHb
2aW50Cxv2jjYZCzqk33yaJY9Km4btpZK40SR65KJkq8sU6WPXVih/5pQCE1tLefM
J9ELf1BsUPR7tc+c+wdbCoUfNBCPTBbu4TiTF5YXSvH8h1oglYkpwaPmROqbeg5E
bsWpuqwIGszfCQmhjeZBPJPBMI4td+6V07fpvBLDcj/yzQF39InuzXcX0ZYB8upi
6ANGvNwZeHxWqS49WHUGmDY5ulm8szCb02nD1Yv+9ANg+sCfN/RUm3oNxC+d75qo
6Q+Mjh5HynFoJBx5gEgtdZ3NxcCuc4i5kjrwNT1K2KSf3xaf7DHmNPdCCguV1GbR
SW4r12toN9jaJFqSVf+HwQhlzyv1f2Bbp/hzfL6u/tHs/yUESl/hZ/kjVPHD4lGF
fZ2q/ZAlOXnG5PkhyIMf7k5IusSDSw0qBiAo9zQTwk3YdMp0BVFK2wGUiOkKtd3o
Hyi/MqHHWBj5OlGPo3P23ePBr9SBHEVyWK3/3OqT/362s1gIzzCNANVOSzy+tjJb
vCCTl7AInVZL4I67PWwG55NLAq/nhmYT3yZcpgFGVz/JXVW8N93Ns9ikDL9ebMVV
Yz/nLejQyX8V/RL8ga/hQL5LtWEI87N388HMfstGSBBCFZFuOFgYYhhJPqt+3b6P
5UseeHhUg2tUzT9fPgPPZL94wV4sW1vLCuKOKFHaZPUYNos7KRqb3GnxKsktY20p
eEu2RnQ69z35ppWCtE4/XPbuSDFRb4cTp1RvTrgzk4mm/yuMvPhg5svYvxBuFZvl
na4L3UtGMbLynKgjnmdWDuoXbEIQeUEDwu8KU8Hy7JnsBC/vpXlfIqzJdBOCU5Uq
z/BMhrgvP8VJoFozWMiNHupi+J8ezVS9grohvWj68uCw8v7LNrNnjO1f+G2e1XTn
w3iyvAAu+HVdksGZtG/jwYgmAmOnssEUvWzY0ZSEOS5EzVBMz2mlB3l9Wu5eiFvN
rHh6BX3oV1m/U1bEYInV+5fWmMbS3k3Mgl8agQNB3J6iLOgqU1WyonCMCyKyFFe+
lAAZIvNtw4b0EeLyf1kVgwebLTIWwY9Cvrxew39fKoHqxDv120UQXqFgBrJl7cJK
4gVkZlql7py0vHy1Ud34lVBayDHOvn9dIMBr7St+VT4BK8PqeeU8uXfTFuJDoi5I
eec4CC0aNHdV6obN8FGfjypSyMYODxsyf60jd8HjahCpWQgDchsGs/aBO7lxOkFK
HW6lo3u0SBB2G9JOUiHJWizvuv6IYiawRaGZTZIArvFSAmWbYEA1No0QvuUEzvKg
CygUc0OWZukMxtdXC9jToWOXRcbRb7AZKOKQK3YsCgIdV36cmOBjfsptRJXRO1Q5
UYo/vpLi/PYnP0KLpJU070u0aFKhyKQ0+gEEj1Y+l0kWxnyICuKj4XyeX2xxQPDL
2zg8HwR6OkqddbVRPc8FwIdavjBTO+ydkqW0z1aHT1OisDbF4rrRA+e8avxXtwcf
gG82+J/kWqtf5MZ2MPIjWGg6nuCFsOeV1klEi/FwdtHVi9ZHPT4I5b49N3bw0mhS
XnUcDJIhSB4YUZQklRW2tuNKUGFT2RgNCeRLHj7qOvK+7vVtCnkVVV9c0MSw6qo2
vKYMJKb74TdIXlRbYnrIhmrpC5zzDyiiNzrM/ta7cIRMUFKgXQ2TrKs8zubEySuY
YG/WMtyTiTGHOl6YdQrP1alfODqEorw8eL4HrEwhQiO+NqdYCsYBaD9hC1j96Rwo
kAB0e7eCA58vFfF4+HZrLno021NBuWdE3y+9H96H28bUOO8jyiZlDvTQrt1uEt2n
V9nxJchWsChP/8Um7JAcAs/C85myHH6NEwuRnacil7v0AcsB3JgAi5vS4u1vFa1Y
SCqwSsBrbNudIcGbnw4EJZ+07Z1PRbOlH8dcXSrstPYGLFQO1RjUmM64NUssDfbz
5XdR67Ynh7OJPypmqmlLNZvkFMGXyHRKFwRUF9PnXVgV4BraCXZdQ7Xy+4+sLU2b
gaYorxPWvRigN2JxCgNglKDUuisJA9dXJpw0precW37FFteKAk24aegNVRQoRXi1
M3l7MQAeUAC2euKPtHucYTb4QmlQDI19AG30vBoLlSRoXhW1ZEoZglS1qm+NYQf4
zWG2ZY+JP8R8XY+yXSofbrOKNvqoo8G6W1GebtykUbvdMjzffn4drqvg7vdLSsYR
8iRv/lkByjHO7HZLY9LhEKRRdOJu0yvEs7rsyM5EW183PWWccEL4tRfSqTs+BfpD
7y4t0BvNisUmeuv3icfRRNJKzmv7GWT/CmAkc00MdcVE3ZX+/DnDz4pTOB8U3v38
bd3GP4RxHJlvoX47fP89ICB2DbaI1VxBxAJqmoYoFVPy4qqACISteKoglgE5tQp8
PYcHhwb7HzGkNutX0LAoBSNOM2fr4q0xLutfHpsZZnYJn2XS2QDDuSsZntrBfyiu
vr+U7LWNLKYssHKWrav8SaJBk0wrzw1oEVz7Fu2tSdHIRbbwtfAs3N/hWLs4E5Ca
Cqb3SKnHnGJMJMTtg7VAR1AkN7AbifHghUQJb+nIG0IudlbKqCG8FlxsMCbEbZkB
b25KncDSrlfWRwuKco+T4loF66gUraPRM0/LTRllwJ4sCniYGy1WwxDp3/PfBiZH
7b/tKk/uFO7tWzqcfF/xVLm9+hEM6tfuyy6xZk36BnoQyJYqHAlT1G+Srs/1whce
kB0zdAv5q0llZUvs0EZJpUQG/bD21pTJ5U7GKw5xm0+OW7RUdwgf2FsSt4WgHAlv
zBy3Ki1zx6XCJ1YMCx5xj0rNwIpL9w++O3d51ej3nJ1Ia5JAnbhfWNaUIMXnM/MD
tO5T9pVrJitdGW0GSdu2xUV7FWluxTB6jIhASnBsrLojNqDM1hyKCdYfjMGU1Haq
fyBd29OI7LjjyFjOuNyHN2tzR6OplDaf/asKc6ZJ77TKEfr6VMQCK4UVWUjj0YD8
SxGxgjPJSJ0h/NrYYlhyvpxbIYCO4yR9ozXGmJof6KwHZEoRjMyrkvCbVZjgMnfR
z0xfh6iwDanZadmgfZGkhpjO15thMMO2SPQgaoCbKfzxtS3TzG8QYY4IiRT3ipO2
YaG7NQAVrpAghdf4bJli8uB7v/atrYERKAun1FwnFjvcdvpF1BGyIclYjBf97N5/
zlsvgb44As9hd5QcW4nIEHVaOdOTq8el3do48O4j13sAEdh6n3SIcQ2fPkQgPyJp
gLyPQud8n2VX6RP4T8S6Jim9XM4oPUGyNFRnFi+MdU3pMMLOMGM5uLrUW970zpkx
UkmBGMo0OTQgxfbywmEDk0jkkKIAKZhYKe9RbDZOJ6cdbCeSJnYF/XFESGBqhKff
vSlnFv+rb17PgdXWyh59bOoMaVXLasuDLmmCl/vFPY9zb8G7/1Nt2D4XchF6stjA
PDrpE5eZuhYPT1B4RKZH5/I8S/2t/dhThMBQ4E9gtOAQ9ml1/I3ljVr7FlPrX8Xb
tc0a+XL+sUyo77nwfKJr2hGT95t/LJB5EdA76kX2XxhnJ2hAKkMwBlchhcfceYjZ
vkBZLjrOwYOQprKDY3J0/H5lqPpgzVnrmr19ckcCmmlVza2F3Dd1Z+Q17CGhD30O
slb2kAyFFFHajOX9eLWvBLq8mWM0q5qwT4aT/VDTsPVDdxktOD+nJAmyUg62lwMZ
XaFxiDQMXX9L+IwFV7YppwI7EmKJlEs1HMNrCzbxeRvwBLLhKi/QxWJ+9sM1U9Ig
eQ9If2tfp2N3wxsYcdOcc/WRzZ3a2X/Obiwn0l+xUlyo6b1VUkoiZ8bsC2O5J3FC
aR92S/p2C+v4rECTYFYH4p/+jNFRzyPl7lm0dkrEj93yme8TSudbL1i0+jwzFC7x
3/Rgzcwj093v2Z6k6oErr3Dr+1NUAKGoXjnoUNJKOV1GPkpq3zTjgzXVlE8OsBQA
OGjII0Dq3O74x+qo1iND7axE5XX4HODd/UTSpOlX0DBm1KiSA5h2LYQQVsTSxnzP
Fo7O0JK4Ii4FkjKEAi8vHTrE3ePm5g6hJFgk4g+sABxgySLFt9tqGfeZxo7u6fDU
szJRN00j8fYe9PDQDqOAUGYNkojYnxFhVOZao4Y+kqHPwQaD9wWMtQF+MlOs2OYR
pHCdnJLLusievZEu7PK+frvYkbjGOuDp4bv8wXb90Cl3BIsJMbSbeUXLHAQhqOFE
OoovDoLkZhsk0ve7lJZJcISNVFkwWK/BwgHyNh/409v6dCwistxQUI3Ao/5Ntqf6
IvItZEMI5eXgI4+EbCmTUlJI+2QrPLDBPLDhcWxGskiJVvfiY01Xj05m+wrSm69X
PSPM7nVG5IhwU+uTphNwIdmAXuj4mlXf+UCOvdPnObqRsfFI9EZEC6i7YgXmLIXh
MckHn8PPZkgxkA+K/ealOwVrYLZ+5/91PPxkTNZ9uFSpOrCjJecxtAQVJKlmfykC
6/YyKMa8BqeFiH8QgWt8bfGWTD+6NV45SH1140W3laoYUD9bNBt4JplZEQ2SZdEU
8Whf1yeVfo15JVl2Q/L+T/dhtd0VerIQSJsm16p6E0pM+lQJA6iT7l3nO3ebES09
uRCzRIC+20DfgWeb29YoYSUjueFFcCmpmSUFtdXYTaXr0kT1XAnthY9rd9IUOt01
kt9tVH2bt8pICwJsy4QsWmN6IM3wGEa1Yacs3XMmTvMv5aHxx9KlOf+KxdWbdkgA
syuGndcYHRuKfxKr5IIM1xF5cKNQgNTIdxD8FFbiFUIQZIcMYgr8sjJtJVXZ24+V
jq8OdI3pPTRQigrNjeFlKLbp22VEvCvMVN4gNFnURrKlyq9XkGWAPf/+hoFan/tl
IYoXshvXphOCIFtxkLVA9VcNV0fA4Ji5YcbfL+S9eM2Jh3o1XSWYwHgymBPwiS1/
rObG4aHUeYUBcBIXKDab5BVdTcmKWLUrFsGLnhdE+7H/y51Rv8NAU9RQJ/z2/pRq
1efdz57GEVFFViU8NHTV6hwGrpTI2PqMTh0o2lUex7VfKXEJvW1EjeLIWd/p05+h
GVhYw5oBjpQP4u2mgw4669rinH2dOELkLKGBD0rY8vcaUZsz0LZq7vAdXtM2cBMP
O7MiqQJ8OM/brQrHlK3OtNXfEbl7y5QVyPwQFxoiPcuiXbs7Mb1mkIQRLaZ5fMQG
UmXAGO+Ub3aE1EAb2C80hnuE/x+R1X+OIBhFEEzYYkL1MfK40kofP39ZXmWeZiLc
sLLPJRTvqzH36rJd7F897B+jMla9/wXAqIm09qrbZcIkLpVRTRDLRV2sYCYrKiVk
exiqL/gKHAUtLdOE5HLa6KqCO84OaN1Dh+H7hQXSHwQcWDSXICB1ERRe0btvqaa7
tAStm02CA4z9rm0A9UrqBdXgXVxC4jzZYInTJMMU2N32eNxK5b9cv9bD3tXl0Pvm
SbUfWF/2wEXeLrh27jf6O7wLjh6ujI/Seu8lA1JkkpUhhWFHFA3f639Kf9k0wnDs
bWmgwvUIVcJjQDSCoHwAJPIoykesegGwQeVadQRqL6PoZtj6hsajvYyNxqHUeOyR
HcFLwYv782wwZ3APeJQcU/MU7r8UMNRhF7BXaiZOuA7FBFhIFgCLO7ErX0RsDzyt
V2z3/SXQI/rmT/wcqy+uhNRxMfMXw2I6MyYXuLZjet1pBMYhOvUVWCwzCow6EWft
tc7uTMTQFCRoGk69IRzMUy2WeirlaJr3id11U6EKbOb+Vn6r0Y7IgyVSvhDOD0yq
PJIGKfpcG4gH98OJZrVf2Ki0PsVcMU8vhNNJfpJVRut8vJX5L6Q4O4gYx4nRMz11
t2PYiRw0axnByMp1p4N7dIDmEr+u/3+oefJwWJxfr1ddWPGOzYYF+jbYRAYrnv8T
u73Il3ZdWLnsAvsl7iPkUn2j3XmHH/MTRnllx7cdM/ROT5i8zEepapORmdmI2I+6
4DPtajTcoU4unaPTkaC0xBUyM6hYA3JYfcINsA4wTYmC6TNj49VUuoyJERn0w0g1
Pgiu/uMYvEU9LBsDYOBCTPG1UpMUuDO8Hc27qdtGzz8blw1hX8L6mQRTnxdqoxCQ
U5JixatdanPNlHjafWqZuocjKkSd+Isc/lJPuhX3iIA5LjdDNIYjwCJSXvN9XTiG
qLBUIrv/wqI+4hY6Atw0oEmeJV6gXNdnX9UyTbnuO9QDfHaiJ3PoNG0p/BgLg2YT
hSl/GXoghxpa48hJ8gvoncTaHSc3RttL7DhUdH9XCpgwz/QrEell09Wh+CF0voGY
brB90yq3aCCSDZa/HLypunUmuJGpQZjnQvrksoJlxiIebPF0VaguramuAXKSdxzJ
f+ZEIJBzQ9qMeNqwt1Yw9Xf3nmFF3gOW0D2vTaGtlyoZztD47K5DtLnpGSusKfIq
xgwVvliySQ16iUpaaOEgdwmtnrl9ycFrF3LJVltMBoAONMd97AyNRQBQtSKsEulR
kTGBLs7HtQmPj/EWmRvpbg+ohKWcmD13NbjzByeGxgedKpe//ntel7ShoroyKQXD
3qhNoqRNUoNGG8Y/fvgaAYhh5fuNdSxKumNNdw54KMDhe4OfCiTDTrq4yuZynbKR
gTJUyLCEyJR1x16JCmJeFvi0bKq7Sh8h55VUtmXNamWuWxm9QTwIXcxmG42He/Ls
oHT8lTmPSbn+SmUzE9hcc2nZHpwRh1g3r2Mff6ecVvclgo0aELGAUg/uJkd3nZ5b
32HDFqmA0Y79r+LqPEioOTpFeNObdbsD6GUdKM+vzaB14wcW62FuMA2HGiYxn7DS
8JCLjGhV4tXjMSO8z1l22t2nQyAvdPYjgS17mRMuE04boo8zWAqmJGAEpOASPQXf
1rcVXxWA7Gn3TbnpFM7MY6nZ80H0KCswWHMH8vHZSqMtjmG7EPU+NWzY7kUAjlOM
72nP77w5oFRJniKhqS6eOj89bi+WYSLffxq9k/6VzN0fCIR90dF8c3Z1GAOb6d7d
ELV/swGTQeiihH5nwcLjHQT/EFsB5uJ1OiRTIVNxKPuRTtkxMe+yfWZd77Pto0q5
0YGrSzyoppARt/6Nr2i+GXp2HLgLy6mLVfwiUdwiad6o6gBX1CO/7HTfKh20U7PO
N2hTNkG0NxrEFAN6pt0DXoiWSLbO+ALgd/NpKe7ppqsD/USA/pl/ZFuFuyBo53DU
Cx4lUt2XhPQg1WurlJDm2o3YSNjUcmV7oea3xTwBJ7zEm+15ZfgaQqamf6c+FDCU
+yqXAvR77Mkvv+NtGnLUDOKdhPWgIOBiLHscujQsB3FO0JDtLtdZt5fCEN5logF4
cLms3CLYjYgg8MeIb703JZYwThqLa1JZ+CNEchIWs8sD6R7sJiaoudMkS2EvSg62
M6zU62P23ZwceeEIriIbrLi4cP1mJ6s4h4AQC1GT+LHEb89GCZFr1rB78MtBeDpm
7C4oVxyF+6Xhe6kXa5uWaPVhj7pEQ4Nahgtj+LMUZtdMPXDx+tK5K1eEBeQt+QNr
NPoxLvh8xjpnN1QAuG5OU9nfzvfrZxpY/r3hKLhhX0p2xwwA35llsuc7h/5JC2dj
Rkfpl37/oq/sJKUNPPFEQIYi9b+IdzKNgjxLLYwBKmUa+mQGo3FvTBZO3opYU7ip
TTC5AIkk104tOtr55hKwMe7r865ggmuNfNeQyuccRUAmmRFQsFM0HMil17SlUlrE
axM5JsqYsvkxf5YvXeYrg2JtTSgd5UclDIOkuhbEoiOnihGz5UHiwgohgYKrJwye
r3nvGg6UBBXCE751eplkkwHcP7NUUdCEZOwV4SAJbAm/ObrWfxUQX86fjlwYhnqL
wjvHOIa+AW245+16MruYKNNVWH1R2r/lL9TXK2ZBxdPjrh3RMs9bNp7E7ZRsB+E9
9qP+319pjP00q/Z8oDwXVQeXcdytVNlIiWm5zkU/h4M4C20Xm3XfLwo3krGiJkFv
GlA8+6DsP1AIavjqicr8SJQhYWNsp4ZARfEG8n2lthApIaPU6wUqmxmTx+b/QyQ0
9WJGHPefmjUc5nOxtPB0iqUTR3Xo6b4BtuGUMJDW192EdTzFD2r1HdVGUy6aoaRY
ofhBUquNk4jJBTf25wPtxzChLlzys/sWYYG05eqEEMsfc1rkrjQyb1hQrWFxTgnk
Zp3YjUzZgWFISaJ42kyGFQuaq1+h63vLSunDA7IsJsxioX9jEZv+zt+7MhCmZKnN
KwNT/KVjvHGTsozxk59HgPo2scA5k8mNhF39Ax8muqQL3Id+wLzUHbjMf9rwEU9A
aqe0d8/FSE+BIqG76goTxhJ5FtsJKrNJaXZ6uzeYzWCJM3HhwDkT3jyjwY1Dxr62
BWBCXyKTxBKVS1U4bomgF09ygQ0lakL/sg4TFaQV/M94909iK3bzEJB9Pow5+C2I
9apsK7spEZ0gTJ9ko1KOjdcozi1zVAbHXxUThJJ1BiHTjQC1P7R5q2ZjEaAbQcUY
7n/NCWvqe3+nW0cI9kwDwH7fdg/4wWzRJBaDosev/cyfxRP8bzb63jrJ6BbcVMCj
olXqGch47nKCAHJq9MunJReihtDIV6mlRzoVHMsCqLEUU9bfsYTydD6auEb02t0B
FKN1ig1N/FG79khBxbf9WSoST8DjN72v1/mAtUYouEE3jUVcKzFZrKMBWjx4dMYj
wtEI1Q+ZZV4Vhdy52uxd/ohnRjY7GLQp6HFFcSG197hWOoF99pjylZKpRChSv44u
dvF8Dp4xVTCpPFpDwF9Jz41h+swqEz1OrZKh3yLthK/pcISiEKUcCbsp0Nj4ak98
lQ41yVkaSU6lLd0DOZHml0r9VYk1UqOwx2RFwlDjUXpoj7b7eJk1WeVEHhsXo41s
h6CA5t9QLe1peJa6ddnuXz1OCF2FlcBS5FTrLkpZLR/3B6heeoag7/kqna8Q8HHB
7FfVn4wybdo0BI41ynvxhyM9nZCsT1mEeCtj8z55lktLSJSgUpk4oxKVtQfMA3Pi
G/qIA+Sr5rbTfSU2Kc643JeW66/jVlxdZXbUefrY3FFTYtLD/AD960RwbLjjZKAt
JX7ereyzkBr7JDqZOC8MMbLgRnIbueLW2rXsGA7+h7gdt1FPrmjBrxetFqO37+pq
1XmgtIfe/zkxkVZU+1pcfzd+Z1FSOjYHb9LxnpCKBJrjN82rWY5a+K82I7uStBU+
95uC2renw193EIZHc4rEP1juhD6aeig5PU7mtvTTq8qKI6vgRyubV53PMxKIyAb9
1W6GFZkzfpV/osYwQEzXINDTnx5bwe5VreyyBMw6OKxukwafpcBNW43CMZKLgqqC
E7NBAvXtCTb4wLJ34C86yqvQWsX6pox7rW2iyMT4fW0grf68LFdSxIYYlHBr8Lc4
MYlTXxiiLVa/+ip3vLmQ6Kmeuv1sCnDrcP/h4dSZU7yxrWMM/RgqL1It0DRWgmyI
T39tx8DqZSUv0IGnbqD712WdWFm8SrWgqh/TjXzK7ijawBbv52GL2FxMGoJRK1QY
VHSPSTCq67v+N8JU3Q2ooPgu4xv4H5e7p1Duy8g16LtJ6iJZNKyognsSQ5GUWjZn
VAt0+tuDZY0KCBKjbhyLZ+ylZ/EXdz+aSZPmKFao7E/ZGvkFdDv4zhmhTA8/fcD2
ZUCW761sxDnMgjTo6B0fa2gnyYh0ureqyFLEUhV+OeN8afCJO/mV5TZIVREKB0Lp
RV1F5AsPfCPQqHHfhEOsWmQuAzN1xg0kzHffh16xAedhV8xS38OI0MzwtpTtQm3U
e5MyjgnEQg3aTjt71dmGdqKvBJYBMuqgktUM/FvBknIzzUn8e0vZqRIohc2gRAbq
uyNKfYjwfb77MCBXGRpVY0YYzmsTAWnU8Hl5t+LzyhD3rkfE/eGxhlyzADwTtqbQ
rFsreNA3tnDFzEp6pAwEmgbbDGk03Zt7vJ6zQ6YiJPDCC7hQKKVwysYD2ecjqgNX
58Ce/CQjO6FkRWs6OOnMhsR4LCo7VL0mFNkq9mk62tOngFHIClmCDHMH3nSOl+TD
GIVL/3MfR01xp/sAjY6MKvm2edaV5grPbJVTspU6dtbjWKZT1SB+ubLzs+pr5n5+
cFUhQct1auXpp95nQ3MlO3213gsEzh4C4uAGJqcTYQ+FU6HpMsbnJxpKmTUFw7ok
P7pwG1GbvgnuZemFB1qqtWktW8iGAVYIRJ9tTnmPNzIFkO+3Dx41yIew31jdm+9X
76GSDlf4DYl7XvS69RZrxAbCj7Acc0msK1N3R4EBwedA9bsTXB+wf7b3JPbNJTnV
kkTMHF2DdcOfD2iJIgSJJ08C7Sp5bH8Fi9KgGIyfg/nlT0NE8OUbM8Ag1Ygbh0lP
66GmvGAPJvc+Qx6D4QBnVy02CBxHew0YFsSwWToF+rTV27Q/Gepf/io5Qgi5TQ3M
b0G2iTEQeW7Z7dIwR7N/RaJZ548z5Xi7B0AAxZ7axRkgO5SgfgLTqo+1cvQramS/
zcxShdzX6gHGXIbelN/mNH+uEpRwaunGEEUEWsDQti5KTY3TbOEx27b+G8pdOOTi
3boZovwGfaADAoTZxTwBCmcDPlnT+UtlnFW/1K1lhOSVv0ePvaCzeUWS2+88eanV
zMzTaYhbiiU4oFr++54FzW0RTCozvqa8SM3ZWXAnwgyrkS4r2Xh6TtT8nNggkwIu
9mag8c+f2g56LAo4pzsuodQS5SsNFiSLKwW8WHTwm7rinzOohfMrnGpoIgA8GMkR
vjmqxRV/gmItQ+wq+nlXV/cvk3lrDkmktixynOOuu4q5/oVGQpTgWxYi+srPgzF6
wCFpfkPnxQf/0YrQ+2uiTFXyuboGDR40r/JyKT7/5Wwj2ByrpwJHX1+jH9xGZrfg
rNrgQI6DvmshbLuQQFtKeHR1bQRjkiXhVncuupz9/SHA4CrNxzSzg+jypz5fsDkt
/Rrg2Lc24AUxy2lAdeE+6KNY4DXcaoEKZVyCQnW8X0NLIApLBBBiikjLjgpTBghO
eu+g8+yIpX6Alwnh0yjcYx9anS5Vr8KQWs0VAlZqOgIdwZX3YkC+zD1I940fzRt/
p+ne+Xif/lzFvJqRbOgz3alWiDAAIkmnOacjxH5EkbO9zFea45ahly/RZEptrCbD
xL0ePBu0c9I+QYgy5Yr12VNKbzjt6km6TI2cDPQ8Zkli39j2QGGlczfW8OQXRcbc
KGSBB00ig60KFOOdL2Okl1MU/9C1gVCljlhqKXG5EAjPxsnSMRp3QR7oolxDWCrb
TKo9VQ5+I60s7ti19dPe1ktzlC9T9lo+svTaWFrfT8QZCM5PMZhquTBo3XX2Evpe
Pzzfw3waTxqyemvb9GB9Ftk9JD+vN56kgO4UMfmHj3LSqmRl0HnWVVJo9slP7PgA
hl17R/FJ6TretRpANcilOC+z06YJA4eydvf8LAB5FxoKDIEl4ANyW6bwWYxjaOEx
mpHZqZHAz9jJL/MnSX1IpfL7IRIb0rJ4taZtSs0U1cY/uo8FnIrob3pVcx0MdTji
DhvOxANsGK0LuTc/gm17NeUWJw0X+zs4WZ+XiGj5PyH7dFBGT94roawhOD8wF/T4
7CYsYUssXzjrOf1aynWPMTQfv16FtnZiDU8SC0PxMewJlu7LNd+57pgke3TrOMsL
J36VpkUnlmJavemjwURX0NJau+U60WOG4O0lJSobEFZX2vqTbloqeiHH2cWbZknU
GpI6AftLyuCh8mcR6EO1zaB5kWV89bUhMm0E6mNFhOy4AcvE7OfBMtubfA6FqldM
8GSNCp7Zwd284BHlaQR6fvoTsVAkPlAkDDrJAYyGSz7TT+fCEJbYbyHZqp+8HZRr
fM2gsgtETQQUCmYR4aMEmMq73QUj9/fW0nHB5cxx+2H/vIjV1fhBGPIUitncfO0J
1zoSUYZhDzr76+tgdYokrOyhEKQLw9EV8DIBBUFe+Mna8WlbfF8wC8FJmo8GRtvB
szIZFuDTwavKapmCeEzuGlT1iaAgTH2cMwKBgdvNRtOzUbNtpDSaLUgHEnn4xVLZ
7zjF/cb/CDtZJzvNJapiR/Peh1gxYNAijsJHHbn9K3BloyGfmhSvLWy7IndEX64j
80S7d5TV92WVg0/cn7UM4XBgywwGkIc1+znM5Wyc3D2TVRX+XZR8ym116497xuhb
YgxRuL3giOOkM9xg+SnkjThlISEfIhV364wuVBoQIjWehASRfdkY9/9+7Rjin9Ls
/2mFGDlBofQGeK7LjLW3+9md6MayIcfWFS+DdVBS0g4GvoR/DzQ3T621Ber7HUWN
4PF+/QA3KCf1KWvvwfYfuCDd6ZXZVU7jd+h8eq18FYEFci5UzhRnpyFXGPkBm8tR
8OibxV5l3TgPo1CbJlrceMXFOKFqv6CCccSjwjoFXS8Ob8htyaQALDuXsoun0Yyt
L/s0nTdJFYGrSAIK18ycY2dL3+I5pA2ggCRvjlN6IwJzC7EDQ9n2k3unpVacEGEf
p6j0fjDnZg4j4H/VLhFsgTQmbJMETlOP4i1v01ekS+h2y3VYCVJAmzIkGaGjNMEf
mmj2gS3TMMATZPuBA5cZZ0bXiGHFi7C5yU1erRYccuMHk95rZ3h01s6kk0UhNsKZ
LY3GnWsOISmPFG2jYC9Np9dzDtI0OCKI9iG8c3r/Omtqo8RTaucNz1Oz95r49HV9
qKm4uklYqvbe358BIsnjM1NbryqKS2Wp8SaBiMZnwlP5qb9I6fLTYJzJrpXMExKK
WwSaS3QH9Xv+gTYmXNzXauve5A8oqDm55nnAmXB04YR++vByhQUDNnOOIx/VcQpG
XEgmGh7jEH3Jk8pMixWc5dyHqTJ7CKGsSi4ricWJL4ZGZI0KRc/6Z8evDdHpdSPl
PvGQIL2oxKyEUdh5z2VQjOGoK/TNwv3EmCrVyVw18Pf5ysxaLcCnIsLTcFO5cH5U
StEZ4jm2/6KLV7Qr9+3RaknRz4mgdtxS3nCz8brqJR1mdalubenZ69MiHFIJfxyG
0sju542F8271vkRCpdWzgPLeoX1nPSLMVc/qSB1pbUXPWLjSE5OG49BkUksAVDHK
1XVfPfKhDGfuWiTAfjnISuZf4Lg6TuKJVgbR+ilE+qgFO5W7MX0BBCo26w4sYzfD
9WQF3JoXwYtqCzxoxf//OcvXo6ao6hlCHzCX74ls6b6lxYZok3XL+xepXVG+T7qw
iZ/slWPRU7KZBWwMYACVE17S2uZPEyQ1F3DydYncigX1tDZ5DUf/Mbb1TNH9xSif
pcn9E4VF0Hfh+Z4Buy/ajdQdu2fLYKpFvCAxPg6WBd+fSM0lQZz44SZeYZ/WNG9c
nAxcruWi7lEVXBOSGvoOdR0NYP+HoN0YSnIYgbLk28JQqtv69OjYELq5Tqv7dH8W
dEAr008eZ3vxYzi9KyigqZhQH4oKX/21Dlsz2NKMm6ABUQpIOVIGzfSTcFZq8ags
V/SjEJEJbR4SUUrsdY26qw4RlRM8HwIFfBxybcNhsjy5cqL9iA8c8PNcGdGH54po
azVx4vyXeKv9NB/8p3g52OWiiBPnaSpZLF0NeLhrzM9QKINP3XqF20FptqJTW2l9
at4HF8N7qm6t60hVd482nDCRXN16hJ+0ImtQek+SOWq6S5LswlRIbJincMt6zAVn
65PEcfvgnTt2tHsRzP/O4hB95ypvdo6m4DLO+BrLl4MpdFxjOpz/yK8rNJEsDTUP
FKQjYJRSdL9HwmWgpAMsAEh7AzgBsCEWA4KaUE/J8g1RjMH53WXFy1TD4M6RWxDY
3/ht+GYxypUDWJXCKsN0pKNVImN9SoDP9o+FAY9f9HvhGHDAzX+u9c4Nj1XC5uuZ
Az1+7l0wU9LS1gIzCgyH1I/Ia7z9q5r8xVoVKBdj0A+hrLXhtandgqQRtvjk48X4
7VSzIygMyndm2AotgRiOE5F8GMC79720RFa7xtVDiOqee/0rvzjNMtKPM64foS1L
5zyp1O9q2RpB/gys1mK30Z8529p/FYpoLFD6W5clR/fI8COaQMQAXPSURq/IoMEO
YnK5/3YC44rRIsCI8lTYP8g2CbO6iZIlAsOpN51+KwUqncWkAEfosvAKwQSfOM+6
4zH2DR+Fbht7Wt/TvVGH3xA0vvjc3gl/cuZUroMG/MKL/yryfVVPkczeJ1GVha+k
iMV0OH2VnE/IdBhGDoQ1BpNV8xAQmJKxcODHtJUDlRGDHVoB20Wvwo1aoWvNGsZA
JL4uQBnGHY5l9I7qljQldZ2bDjKIR5FjYfxvuIWOwqkOP6UoFMW2rq0aoCLnhAMO
+76L66nHpvcXBWAZ5SYg5RPVUztKq65IFrTDL5rP3FNHHmqAM5V+NC0ijExukudM
CFRFEkWxVJdR4MffDQ2jKrSOWge5KkTSfiwiqank1A7a2StXn4YIvCBTpP2u32hA
G1mGzdqU3vQtXW4W3Pz+wHxzU2KiQPqlBm4/maRxHW67MVMggYJFV4p0t6g/BD1Y
etZnMmg+6MpndMZ0wJquUVoPNolf9rMIL1HDjdVcVu9QJxsACcv4WxjKF+Ts61QM
AoyRjXox9OHyxzYd5BCKTkJ05q1JvADQuJvWjyoZCtGRP3bZwaXmuZ0yE0ja4gbp
YvHtUat7cT73xdx6b1avpLGPVU2Ix1J0unRZ1LRPcW4Hr3NeTc26UoHTR09ckG1Q
YwMxsZIXJ45Fi30UrsKtT1r2ecztSaXLr4eYYaUEqMhWadIWJDmE8nw6WQ1S5YWF
q6GrzemFk+lRMREVt466t/mYL8FZ+ikdEqwkPixEqdv3X6En5+Zv9ADx8nlCIpOO
lv4oIy4dErdhDwiptg/2F7LwvNoMG48kCNBGVL8Tk/x2f1476D0eFLMo2YH0m8tm
SwLLhgs72/SXa28eqF8HYoG3bysLRdmMc9+cssSuqgYR/ii93C8qUP6+VUN/aB4z
KZSLw/zHD63KSZl5WyWT3JqQLAYuKinobOguYWYHeo62cWVlzJdk537pZyfRL6W8
1tmX0msS9301WPmkzZfaRECT2gA0NklkJLUNPm1PHgcsOhf1Q55g9gFSC44PHIh8
SkiLggHVzVNl+IKCC0b3kRdWPZKE1wzbmgHQbrSFIS1QdeewookroQALDLage1sM
MFy4alQ3N63TGTkstyQWKn+prBJ0S2HWGSOb+Bqy+Q6pAmCo/ueDmHyW6AhOa8Gi
ESPx4+FnR/C5MiRM+IMEAYHBeL/4NZiARnO6L2OAS3+DOmdGoMm9d2HmgXxSFuQN
ycyNW3h28yNWNgsTr512zj0DCOR993QORE2YCc9VnI15PRLyMHEGCihRdxvOfUGc
dODtSCun8wrxbq16uY+pezoKObp4W2HPLjTJDJorHfJWhumWAzc0Gqol+vXbStqE
N/z/S6XdyR2yPlFuccMvnbaZy3VYM21NoU/0DiUHminv8BQ3O0P7Tb4lyuBINlbm
/mP47NTWzHByMxqC+nbaxX1nz/+fGfPshJIy1mC4Y0lvr2NbW2wn0U9taQMDbjOw
u5pBa1NnTt0+jKLPiwuz2lo6gsoQBofyDmr5C1zW0HduzHfe3/1g4OR+3me58nQE
qIZK/2zZO94nLI6QzsAJ/X3eHo6iIpFuIfbq9bw4xuPOywJujlDSia2KFItFR+VA
nQZAWzqerHX5lEPqSMWZh/GdadIUXyi6sTJpzMVZybvxAWVb5k7TSsRT/wo6SQn3
5+mk7aXl6mVQtRmZYWD6hIhO0UTzus0OPs1u2SlekuXuxw2zl5iNCzo87Eu/mdJY
a84Z6kDXCzNtJaDMFZiHHp3yxtcnw1p+vV+lfF4epPrnVm/L8kOqrEMNtI791rtW
lRB66W7lPVFntVCu9qVeb37ljXtgTLSc7BNh7ZY8xYH6rm5fl8IECzaEuDXFeWGF
Zv1q6BnG2nIS9kBmBwizdUsxW6hobZhDVj8dv6K8MPG4NEwLCtCJWTVMvnTrjIMz
w49Tjf1w+DKk+ZcG0QQiPVci+iVmoLv12JlpKMf+bR7ei0WdC1NL0wj7cha6rC9c
rupOyGe7qi7waJH9UeZP1xqJxixNCAxOQvhduX6MMFnBDEL7FU5eGID5MmiIdsff
UTfYIsFhZI7Ntxa12BllAaoxKzXFmASquDNNXmr6tB3Xyz8ipJvDOabwMAVbMiF9
vRH+pZxl4XO617cSf+7NdTTixUKROFLRPR7P1Q1BnM17+ftp6Rkzrh6tb+lxbY0V
2JONjpdSHdv1uKqqd8zwKZH72T+l6394UyZvg8WytVOm3o/fwOpgyGnMQaDkIHa8
fCNmX1/0UG5o6HjOCLo4GWocrD7w0ojhhpiUFF/MJMIk26d5Jve0+++2toN9Yqme
yQEW7cA3DEgBcePf9q5DQAtfhbS8zo7T8zgNp7y98eTkcYWITWGMWaqmpHaOOaEV
ymKk69JYaeetzRaAKyqh0HMQSSiW9Rrs5w3H7Ty9vXko3cPNczT06CkTwq3oEreL
x8SmkF1mxLyQvm/3ibZL8GyAu/TXWauJC9TyzfYaZhpsqp7JEdNfDeGrTzHT6qzw
O6oXmt92a1xcIEDG+PF2SiT+raAgSJ21/vIxZ5tuvkWbbqeqZM1Xwjw0bQ3MwhS5
+LMDmR1GFhRdAhFIcjymwPdA0c91CQltcINCyEuxe27EZIUy4nSA2Gx8bS/Hlxlz
qoxWOKZRclrRdWTWmW81TDzb0Gf+NHuqEz4KAO7oIp+ySHBVGin8ZbhPJJaPQU1S
0G/+o5iSpmXKJYsMrnGkygR3ZVNAcrnALq1vr3HLrOGPUSBs58mgx8waiyxadjC0
lr1ZzXz8fbveCtPJHcOC2z6VM1Ce5nj1RRYGBiX2QVcPUbmGqPJcBCiK5pc7bHHj
LssipHLWkvTHeHvspUF0/xgr/XZLeyc7BDaT23FgQ+mR8qVQnva8BtNQrzrE94xg
YL7wnXf7dy/eJBHDWCnUQRGJCA689SRrVuoRc2vJTMoSWmzFisjIZojUrZe7MQtm
dXjBDWLp7xkGhCiY9Z3/sP2YqroEfWRGp/ij1+h9yJdK6+oZa54jvWrVe3HJ52KQ
SaqoQ/HGPCwKLdMRAHsQznh9V9rIKc2CeC1uXBSQdLpoDKFC2xVdHKE3uI0EEB1b
y3EiHjGMdaataYEVnKkjsUkNS6nouQnkUoXwwtZDLa9Gpx0yu07gC47Awc8NGyCK
MMAgRHZer900tINYjP9Xmok3A8hPbF2NJ1hDpgAwk4874GJw/pB+ZYDBsHesIcw8
Tzvc1fXdtBVUS+PnylRZarAMC5hbrpP4xiNXkMDWim2B1lJeOURPanzKhY4GL8uS
20MrX+SLeQzvfviQkiZbCsOPD+C+gktOr/oVCP55pXnv/6PxMN6vJVXLwSpbsfCK
Ky30V4X8w+RW/quDI7mIq03PmEThY9Wv06HKOF5gd2WV2Ho0M4r+5gbRVlk1vR5Y
Oh71QyNdOM+kIQ/2J2Joyv2A9o1At4oQjRC6q8mnfQIy28mx8taBDovyQU0m5cWf
za5/tV9KLWR2z4VC4I1jZM2l/B4P5t12qNtGdgEx0fP+IyhFmztVaXTevgNsD4TU
NY6adu3OUly7fY9sQsbkgnFeD9H8sWgaj+gGZQ3TpnnLOuOd8EmwdtiYxAJHvCjS
sHJE27/LKFx6Ga9HapiElNjw2dSA1zWSFi/HI+aAWz8QCpR+MPeN1vF5saj23/2y
wfnatipPE/I3IOT9WRHThIT2EvRbT6kkE289xvydlecTRwsLVNQSfIuKXq3otbnL
sfMsXT3usm5xC0F+qRHJcx/+bugthVkhTkbdfjiJmQ6AHszjx2VpeJQGpOxlS06D
ep6eUl0lu6lIuxJGzK9iVSZXfoawyJCCDNcNwNc8Rkb31Oc74CZdG6GUNB9TkcmQ
tekqqMwmsYReOKLEDBdGaMIY0yTt1rC0cC0oaqhbCMHga2nBsyjUoEM4NkvN+Avy
jEill+ueJrlBaaeRJAGCIsM5Q+TSF+mVILFOeZXXyu16APV1OuXYVowU2B4J+o3H
wjKtjTB7RlnpIvh/2BLlA759qjWAq2GAm8+GPUzG5XZv3ZM12PtQEH1a+K95gBoq
5DZxf+374fucgbxqrvcYIcvUfdskSH4tHHUBQ2TnRb7G7sKARZysbt57Pid0wldz
7uGWeI684vJ+s+gzWQ7uWtb08rosnJ2hHohrw6GspkYEPI282HDBb9icbFwgFDO8
MsCBSjmQ4C9BeKNMMocUtl57l+Qb9HKYS18vwaVzeAP9qbiOuARQC9dnj7dVSF9C
aFmopPViuitm/iLL50r9DE0KZkiR222vsxAOx3qp4F4ovbZS4rvi9klk9gBZnmbM
fCAQrh13RSCZb1AsWKVtHETo0evj9V44To7ozhcN7TfMwcjO8p/MMBKh46Q4vB0G
Fw6wW69mCDzIyENvgNSinP/ZV1TLlwwstcugR9Rzrb/fqpuUzLiZ9QP8sKntdjHa
UvRvQFB2+NzRNbDt/ggr4f3q+zyoNp2efPpcqm6K73JeT4+i4dQdaXA0Mpr+2Gwd
nUeS1XUqvgkdHCcospuBKVAnnKAp9adWxchAVHb5DpBwI5YLqnm4xi+PBKzXgviW
FzD9vzFh3ZYqWo+0gkaTJ7pUbJOjQ1NwCeIG6pZEl2JaFnAC015YolyiBQfuq5ab
tEC65jp4u8LeAnxIt8eICdvGApQV+rX41W2IvJAvc8zjHfP5XsZrXUT+AzU3wTR8
clxsqbCKQqs4mldng+uUkZVa97Vrki4Apb1CpFjdmqxrlqdFi9lgXnb4BBsq8gyC
VfGjC4mS0RL5zQ/j8Lb6zwqy+9vpyxJeMmxnz/OGk94GzKFEicjLnZKsQALk1r+t
kbxu9wkZWiGRXJyq8CA763tcKrMM53hQJ/G287yNW2RU7J2V7DykrU3jfrD+5TNl
nEK4UmOBPElDOVF3Q9cZEMv6tLcKvh9vaig07+9QtLHL65q9bjynRGW8RkDovzbg
24fmS1Qud+DmTWhIt8TF8kn4zxl1HjpI3aXKoqsVMUI6NgF6huoVWlcTY+FmFfW3
zpc8iph3T6lcIqE7Kgou9kO28NFrK/Z4fR69JyH1tq8fLS9YCMhPSXwujCcuoyy7
9Q050ZCTs1cKHtLjTrP9PfNmvtqXgf/VT4lS00+ugDP3w8ggYPSEvuWdzIIH+8ln
TItVQWQXhvLHzy0aRp5jsJLVR2N9G0nHKomHayR7v5T+g6CMQsWGl4BdvxRY1Cnq
7dnt9WGfQzaoU6u/G7ZDso/5MVjQKH3+LcS/LPtdS2ByGC9mdjtbebbN1asyTnS1
XR1O9zBqolZ0dXQt9muHWK2W9l5XWJuxkf12PtLeUIneODnldBsQ81KAUAoRTKc3
mkUUaUIpS0GHbQoKjWZJ/fNhk+oCXg92+Wi6ClaZfHpqQq3DFK+zZ5aqFoY+TKJ4
y/MVG+QOC70mZXHK5e3N5e9QiaxmhhgUx6vowr/c1+v+hFOX1tmsmD80umSkL6ja
+Qs9BuY5SqJ4TAgqpxaRyRPYNkZ66o1/ImCFzFIIC4FLgL8n1RoDkzzkNJiPQZnG
bP2I6azkw2fiFzOOI67WqAMDNxsOd/xJhdHjTy5byUFS/hh91DHJ1lbvvPADh8t4
awwft8eXpGUViK2TYXVOG3VvGj+vzi82cS4K8NcCVEOuMHJEnn3Yd3WZ6jbQC0od
GOF8YNV9+QMg/jQL8O2UQzZQ5+63Gi5JpsOrtONRrHR7t0vHk4HlxWQ+9R3xPP2e
8RrjZFOI8QAY/AIyXV3ba2EmijzFthrlsGmhuIhvUT+RqLyfmEKwVQzEIdkBblDG
+2xZzRMylCXv2Uz4RP/52iXRxhO7i+xu43YzQOSRt5saBj5Hi7611CH8m76dyKOV
82NiIwd48gsCVMLclVEChm1n1EXIlxuhjI1Scc+TVxIxPiA1RdFhMBitIrX2LzKS
SfATcq2ZQ0HbFKDMFkKBhSEbEgiPqbkTTS2CGNIKMW51YjkiLq7kB1MeBet9tun1
Tnwr5k2swcPdY1GzRyHJgyBifZ9415irr0ihmXhAz/g6Dca6VoejjwKLvcgAmGNu
rp1LmgG+/ktIIuPICYp1ogHI+W5e5uElfyUFk2RgZJUy6tTcS5UK5qEybPEpf1Dn
GuI03JBi1Tn8U87myt1OEj7jClMKeS83S91+JO7wQ5mwFuxw3WzS+7tVbXYLFm29
7lRdQdN4xw+01KmdXml1fGxKzZiGGbU7YB3Hy3xzm8ZF/0YuwrfiHU2lF4INGwd3
4W7TAQg6Msrr540GyDqTYXCxVOyJIRtzmaaTEk3SlNtrmTdLGpDQKr25u5ofwZ8x
/Jhl6MF2sUMfMeT1Os99smf7QtBsDAVVzA+2qqy8jecMzYFlf8qUBjPk5cQdb3ec
Vg+qUeRAUl5nAsf6gCaL7m/pML7a78tPzT5SUraTA1gpDOqgRcVFN6/2gmnQxp0t
Xt4ZZs3QNVPVWN0kinITpQElPPEgO7c+yblCQquda0EEVpnxjrBISfxH04IbA2iE
xd5gDBH/UQB4vHFEiFy2l+4GNqV655G8g7jIt8gUSVbkoQQnniiSNPM8Eu1k5Jwe
YiWo1EydahrNh7g9PHysfTqhl6YkFbuPVqmC8eL4pv6+ouW/pDoBYp/T0hpN3Q2H
gkTZftdi31bog3z6ScXAy6HqgVo1QlsTUCOUSY7Yd9GtR/7fQbjyf5xUqfNGy08d
D4U+7LMo/J5/a6NfPQPrK4to3EAG4qSfEXNU2OXBBxcgeqpSFsJ/elYsw01JzDcW
ACLGQibNfw2szmDbDjjt1Gx4ZA/tqLXY4/h9O1DALlgvoQb0H1s1e/+wzHZjf/r5
gd8sYUdnEkG7EgtspAwOGg9DFcORaQ/Gna6VViekAcx4YlodWS3U5KWybRnEtDzL
AVpJD2O6KEK1QhYn5w4yllVP7r8igBlNQAk4h578ZUpv6FomgXL+rfDX6tI+B3mV
/xnw+aBYms8lXZPZPsOvBr9ECH7WvL+1tuRclRaZBBNXgqsp7OIG1RtIRjb0LkZF
2izBOOC86+4CUltZFRIJk7UFAeiIXAXCLdJsOd5HRnXAANW6Av7yVIN1hxw9vUQR
j+gr0YamHb/7jmp68b4WlgUzVIS8fNos/0NWkZH62/i7hGvPJmLSU3OBnCBM79FA
v9pmd8jgEK39SqYuVvSDVk2NewrYcdHej95OtpgpG+vngHp64xHbyJZBZvOZGZ1R
5A4G0Mgu6fcScbLFj7ru1IDuwT7wWs/FGJzPtgXHOwHbFoP4RmzuZUWL1u9bmuCk
h6Vg4rK3r9pI2nrG18MDO3kEqn7HxGq3lD5y6V02G2ROtefR0GmVX78Sozx4X79p
sCK25bYj/LrRkDObnPZsgeEhIKJwsatDEr7dsCjPbXS2/qJnNsL6d3SwNXtIUcRG
ajjPZnkKtS8BLOH/nXy517o1+D4/Xve9M7EwNbzyqUoINJK92r5z/F/xA+tsKgDk
IDBpFOM/s+uC4qWyNEdzYHYqCYdTN8tDbxX+oIT8fc1krK1zuuTksnBKiqu4p+Em
wqS/F3ASyngy0nUJ70hiYqTOu0B1BlFc21SqW8t1g/NiHhIckclTbggHsY39E1zQ
EOPzwgnYNEuWdrGS7b/Q8u2nIyARvKrQO5VHh2EaDMo/ICjQSJ/9BbBqk1gc5/sc
jnCsYJqMMvXumiPt8Wv9BXsoAEZMzT2w2I8ISh3R/z3ydW7MX3+6tKQHrS6FMvUi
04XUHHz6b0RPvmTtvhXN9RjMAUlNsEpxdYQ7r7RX3HBuXjj9+A4DmUBGfieKCr9h
4udHg5cb1eyb2G+kxeEWQjjtn70pPdYoUt5xhG46e/dV4pVXSFA83B1IiCmsR9UG
7eHs7v1sYwAWPOchAcs6psK9P9iHniS7BJqdruSwik/AZz25zLKhdPLCB37vHbyO
UuOjkh0U641qODapUNc77fkfuchtKMWXudoqtfzQd8Tz/N2sGz3KRX7Ew1fiRl1N
gh5rIwU0QiehY4Wnzc+D78eJO9+ig86Z+lbpo77oGcjPm68bJvdTN8OnQyLsjryn
itTZKDg3BizsOAp12uZnbQ5b600RIjMwQ5H025BM5vdkycgghk1BYiR4lOY5H+yi
JbcvJO0syNv27km/XHkz5CPpF24xwqvHbrgdnhHWHfGApGjQexMMezYEbTIH5z3W
v9JLghL3uxoqx0HZxB5RGkFtotxMexY+43bAStI7AJ/61acZu+hfGPOB+zo1juNM
+ePsiAM+pZQNLrrAu4WX7NVWWkGOOH04Voi+em0NRLRU+gCeBD6nVVI9bGdTaFr9
cXfR6uEVDiRLH5q0Gl83Y8zchbepmNOMMt1gLCHrKgbGenKh3mqG+eLxcVZj5Z2o
H6XuQk0s5xj0XGZsciGlWV18PR8RGMHkVBL9X+FePPMNPjggcI+j60QdtYagK4+k
/Ayb2TY8eS6TxslvBvPrH6oTGD4TnNmtBPn7BoiHZDQvVhD5wBxEggrc/Z/C/raJ
VWiWv4ztOtM3Mc9036z5eTr79d4xCEEKyBEEA4btfwbLEHHRr9F1gYf8tjJebvrz
KXg3fS/koQzcgBYYCjvVRYDemCXjjA48Wadny1T+Od3gCqMMN1GVOZEIoeuzhJlr
u6xrducm3S8S86lDjIEaGFkpGdcgnONv2T/9rKYDZdUG/V10QXvV3hVcffDa4I9Q
nMwcnuHKd4p64330XfHaMiuMgbu/P+sbo2mKcUAYPZsnHby9r/84X/fnlpNYd26A
IDeAUWlXs2G8t6WXSq6o8vDHywR9qtdaA4rv4mcOGInKrsDOXxUMhZ7af+Vc11gU
NXQk0MOU+rd94tsy/MzKKr3VTjZXNntnF5KSQb3nrHvzwRiTAMTLD6gmX6u0zXWS
yhX1vTFI5KztN7HqwfwA2ktJkLrp9PhH7IwC8pPfrYL0TZcFQAriiSKWgXzHaFvR
CxzsBpaU+g9HxlWTbdEcQSTAe4LbZ8etjbImkeHco+LAP2/sc2cWah/zFbWfOgha
hUcGVv+OV7g6+N/F+N+YjItHbhcXikP2uN6M3LGmys3tEqrpVomt7XkWLHYeKIs9
NVfPGD3DRkV5qxVuFx6D2CL/KZK5ZsQi/jI9KQqFhQ/9nTZZLToHvclbIdwhRVjZ
bApOFIwF5Jjld2Dajh+unx7heG7ObafVNHUzmpxUl4WbA94t1bHsjOauoxhyR3oH
xZyDh1k9XDIj23oFYShnQHtP/AYDUstasLoiTcjzoTx6x2KK0JTodvg302vKFceA
MrKjyt7ZnBI9YmjV+fiuXeyBT64xidMiAKUwAMFYhEZUEe7qWWodl169ciyWMNKn
t9ho9CPb82VQbrHdbWS7L5BeXEl7De6yHoBiWmYnvVHJtPKDh5nI0A31FCF0zSiz
4UkRagUsXOaRBWsilWMQoVqPCRBTOFwZV0Ei3zEH8vC8g4CV8HDZSOvAYlVWVyE/
ayl58NQj7US1BcNu7w40qIihOwpHnT38IWxwl3gVt70fPROpnl/CMm+4CMMPsBvC
pcRxTP1qoQnE3b6zXcEinvZp8Ni8RQvOJ7tZdRipUlhDM844xdEoLZCfLwjYz2sz
eS68FYDaKvmaag7wj3RE7ExcHL7vANy4G7k5eFdl6tzCs0HmccfyErZfaIz8Kz0L
qGOFZzE0lgEyRX0xLNt8bVHB3rYMaJnmJz2fyDIG0x4C+uerSpAZ4WWHIC6BnfUL
j/yurvyl/gK+PuxH8Leef5fPZzXkzLIT/+PmNR+JBXIJjwMeYtHkVKJ3VmInoN7w
Eh+MXFw1WCQ5KU8lY/b7be+tciCCtrRXfunVPYa6mSHy+yNj38D6ff1kH/UyegVl
LuBUo/MyoceMTcQvvP4zwT/9K/FgPPfHG9cyll8YDjRijlZslLuNaINdYRBcbYmE
xacaEn+Rkh4ZormVfRf4jS9SBrVz+Grm59+tNaRJzeIj0DLxVjJYbzdJVU64/WDT
3vQodwZe6HKmkfZ8tZM3TjFz44uPR/jVfcIGR15sWPOia3KQ7fug6IDcaVdwS3m/
FGRuMJQ/787cBrbrtZ3rLugy3Pp1BBxemoByQagKiRWe7twkaCwr3o+pHdfRgAl2
w/4OX8+rGzNwIjiDOC/HUYErarQAkQnMw3+YnWAd839pg4CLjGQ9DkzX0Pj3nzDc
iOZQcKMil+zCZO8YjWEhJHxnw2wXA87G7lW4Zy899FbUEkan2f0cB+xB6xvxYRZ5
hXGjJaSDPix1Q9B+SL4q/h1ix4KGmbKIaUXqATi4ZaIBRHHr3GCPL9xja5u2ryue
Mf/kJYjaI7w/oGGkP6+IS94+3lFVJs54S4WP7ib6qekH5xMLWD223KTX2Wuv/xCB
7XfDAoURuGsV+LErtucGjk9lNUdqEbsuGp9OW+Pcz7zJYcwXPX2sDUT0/NXlZHSP
hGZAmAssYle0DueJ9FV9FWM1o51SzM5U9r6DO8lHK/3uYwQhy3xyhULGubUjE4cn
jdh8vKa2s5c/ZTnsuLrB0UWli3rpk3C+kpNCSoPfzBTaigLNx3crxH7/L2kRf0NS
yVErKX5xaqNu6QUEBA+zbLq7m53k5Km+QSvavOt98e6zrvuVOqfY6rBKpkKMuhcJ
73lDvmJ+QVILsa5GJa6P1cwOeKW2D+/iAGlTKaiOOPtbiZ/D2W4UBR/gCsELvEdC
scit6m3nEvHnLL/TsjEsSGzrW7/RfZMb4KocyzOO6qEybive+d/39ySoCetPmDjf
qUDonopCgcpRbrb/LKlN/vxZErxEDfPAPkyL7+qdMG2eWH3QuycdA3ExxWw4oYG3
ces4Dt+VyA5jTdpLf5pI5xNMVMc62WE0ng2HDa5azqe9lMu7cj821yH5sR/VeSJE
QLDxinwnVOoOV4TCgZYk3x3NxBXWElWpvGp7uvKm4XpSebXERAbjs90jgRXP+2/6
KmrzFbXsh26C+aFjFzC8JA4wNHxRJxOBAcW8gvC+lNYblupunxu9O6WsJQ+lR38z
msHNQcXn7l0mnWpl0n7LTIimTdEUbSHpZsnP4rMwhPU3ZEto02alUkASvVqx3UBc
LJm8q9SeiNbJz1imG9+uvqD+X3yC5UKVPI8wtQgKYRi/dj9AAVA3/Qck6Bk89MD8
Veika8+hVt7lrLfD9KqHz1kZ4PKqJnbFhgJyhF+NYj4Pytbwu0CLg9ctYadFREut
tDZnXmT0AZCxCT8NC+bNIMARvVcbwAaMuU9QJlp5xvRAfhhtnpvrrnmPTMuR1SOP
lrJGzgcNiANoeJVSOKXHN2KajVxiyZMmCTiUyp9z0vArfy43EVAoL7q/a2sAyyxT
s82/EMar/GBNOdjA0gazNNBH9sZVTbk8rhLPBUQiLNAh+nyoLjXIGyN6NemCZphB
xw4h4UzCWDez5j1u0Jubd65A2++AKBuDnz5GQAXWhywfQ1/enwD6ddGJo3h5ymJ2
H5DjXwIIQqTzhFs3gPVcprbxFwhiqHZ7euOCXbZNWJSfgqFIgT9dAMmljxmosRAT
IHcav/LkscnXiiMVfVulLjhD6caYu1Cw9VSS+pVox974W1TvVU/pdpD8/73LKclN
6eUlPUj5wjd8upF5qIyipuJjamXXRjHiRcd8H0CYwxi6SQqEp9Y3+6s+rPuCwoA7
X+KUa8k8ox/jdlZesqIdrf3TcHr73QBdc6vhGn39XRim6IuolfVS+SVT2h25XutS
51UAQYCg/6HM/ITdVZ9uiPTYnjw3OnmlvsKeCH4CuVsKj2ixpbwCeye4vddvDsOb
32ywjQUsLuaydX5jGs8MR3fuL3HNCxZr7+OHDbxXfRbkPAISInG37AS4cgsDoiNH
MBgHVc1RANaGXhXWM7ChAj3Fnji7GvoHXvmPC4C3GU+KzUC/yfiDVMpp2q4xfzY9
o4kvues/XYDCVMOF7xfKKiP3TU/uYWNFgh9DMBduuNdJfy5HUJ+j0tJU49InDFWH
5cNIoguQctf/yOzCv7IG97xCZJKMYv6YPODJAC4L8iMFtlBgHb8AxoAweNWWqw1T
R+Tl6+f7+pvY3p3A9901Km7ZRgKYNLXCVAWI9ZO/i6fpDsFskWHoIucHH1FY1f4y
ghh9WxFTZ4GFHgdRB/zE+9fHpabcGF4pLqrZOeU1EA3naSpUwpf24vbhBKqIkFUg
heD/aVLK4csFEEFRB66jv6dYt6EIvsMs4FQh9mNusHryVzp01hILylhXBjzxRVOy
NK6KdaXJl6ykRmmyD4dRXeaJ2KlByyMfQzKXyCPsZgN4Ag57Ru9tqIjRquU537fn
W4835mg5KYBEkRzPMylWyv1e74A5d0S6YLagYZeIy8UWk63EJJcH4AbIHXqTi2yw
F25f0iL5G1aoYVfY79qu75yBBwEVMDsHhgFRlrdXOYGPsflJqApcDc/4bj+TkcCa
cpLKrQBO6uf0LQAmAqhxRQGMEuwCze9A6FBj16azGDd0S/O+Ac4nTLNBtYYCStRO
L2XPCsIEpPM3M8w6rwg2iPejM5W+zRrvcVxDRuZWVWVHTFNCAG8jrw+wE1UhLp2D
lwkQ8D+YR4ivTZQpW3oSMBI4NdJPeRYEEX/Dd6DV20npkXYmolsP1UB25O5zJiP0
Qu/wbjYxkY/L2G+4OKP7YAS04ecO3E5k8ahMF3DxwylvB4zmj24kaGe/nVttqOad
j7OkqUp8wloZKXoDyr+F/v+IDZWFXX6lwkcjJNA5p76FjkByp7XC33kkUOSRQWqI
rLWUlJDMXnJYsevKrm5eKUXRvQweZ3efJMmiPp8P3+aEL7YDFPazOy3H/UElsSS1
HgnG0NYhgVoKQIs8TzUbSoeX+2fC/JfLfGx0nuzSK5yzBI0U/K4Zrb0tX+qAAyPf
1gwTLZqa2B10Qud2UgCssUgyX7cmHAy5WnxutGBlHCt6nupsuFW7fTLwWfOv3RMS
BRC82Fa4J1Si4jcT4A1AR48at3E560pdeGZLCfnTqm9Jr6SKoYz23HNdv2JaV2E9
054mjMsIYCxNtq2SoOjHXaNqUdpgxHeIcDpCopE0m9biZrF91RUgcFW3GshlOWO6
adGqR6BxiXPuFwkbs7wglVXnaGo4kUi2FEefU8UpoYIRsrIdkZ0jL/h3W8EdOFlw
V4NVTIB6jNCKzpCoRyVuXj//itIVIPbACUagnedTqztyyE775E9UXoIymwc4RjFK
YhdnMj9AuyV3soP44DnFGwbvQwx54iJOou0h3bBHiIrJwRv6n5Njc05GnmPWWYmp
nP6qj6X82RNBSgl/qRTE01RB+82QjrDpo4Y0aQC0EMMAZV6TqnaTq5AgFQTdVjlx
5l09YDwwKyl5X+GRXK8WfFTwSi6C4ZJDf1R4xjSD19UYd9/mXvmRhUwQxKSTu5of
hQ4Bo44OWtbbvU2pZTYGjRB0qZDDQM3vRKMpJ28qqtvZelD28hSeWSXUKZpB/Ucx
TROw4J5nmt3PdLcUNK/vV2jVWB98eHvi00FNis8kNSsj7J2Pd0qyLpxhR/0meOGA
KogohhfFr81a2wP1LT/yxPSqT2ua1MuteUHqrvBsFMR+cCMtC6H0hzOb8UgZqP+s
HQDN+m5QpjgtyL/TYgEOMgS7TiZIM0ZvFlIDcbN+PZ6CR3dfjg9ao9IBv4o/k87U
XK8Ru2dMBPOt/v1yPfxdvX+UFZwvP5RXsJel6i6UvNnIUG5Y81YITHm7CDXjiTa4
5V3l6W7tGaHncbKZ44zUr0hj4X613W0HRMVszzCqPSLyv+713wD7gyXvBmxuTl5h
NqiS6bBx/eFo+JjClJbrtj8W8oVsIoOUQnVylAoCQZPauH0XcuKmF2f+n6EkuS54
sRdg1Bx7oglyK9ipiaadm7nTksvX7oUsfwJO79DpoddJzAKLDVe0ef4Gf9sEK4Ns
cnHg4Vb+JF6hdjcGpep03XOitrKwAgT/IgiAUJeT5lAely+1gVzn8RhHjzo4g2SZ
FuYA+Gh9VdYmaRP6Y9mbVsfMwfyvlhYfHYuA8YHsepM7ppsiq40i/vx+rU13w76q
nC00ybREneqKib5eD/lHCU/uMpfXgriSoLguyHngt5Ew8F3BLWK1Ch0DDEGXzMZ2
0nI6H/RdyUTF0B8MF/NOyvbdohfCqPYI32n3Qrwbeuak8CVeglw/ekwB12bCFhGi
viXEwbsq3fyfEWP8sk6fty8hI01N4P7E8T3Fvm23d5+zujQcx0OfSg8RggVvRL7/
jJogtF9JziK0V8aJsGeycPSUKGJmeG7+x64od6zUQHaq+/edhcWkj8bx+3XFdvSU
jIaAV95cc4QinoLp0tgeeZw7BlMNawUOOoWGL6Ueo37IcX013c6eH5jV46KIXY1w
pNIBwMEz+LYanEIn1du3/+QWLqzyP+eCpFtHcqXQYrSRWZN7j5GIzfErFmKv+Gg0
MuF26KeY5FSJVn5vkqBB80gZXUUpJfKipF/KL6GLLJXz+ptCAtLw4O6g29Xdo9nF
m2g43ermvSqwuz9rYT2jFstG9QKvZIkuVwZOHxpGxbzPgGU1qBhsaRJyml1119ga
AgmvjHwDcoJtwThqPxF6sP8ls1SJ78LSquvpuWtIFcLgg5+ufsRiBMiIQJDPqpr9
WguFBHMwH9HZqRK662coMIwxo0AD6dFcDjm/zGhnViqORWk5KPDRfvw9KKyOwZEy
mikzTvrqEz4zYoKyCr9+hQp28voJvsFg638n9zpnijlIQxWHu7TAObTh+BibWHHO
DlO4+B4gO6FdkpJmlYn5FYpBwvdc2IHVkUapWNjPRgZRb1o985UD3zmI4noxn3ke
1l/qWXsPWjvuziFJo//6yi/fS1oRqvlm4lxNXKI++a85CP2Y7OtACGqgCzw6tyA+
OTgUJe8KHN57CkPnaOCOr51maCoMluvbXVroNOlxZ5vej+Tsklonwqclvuq74A9W
oD/LcDucST1nZy/8zxxmN3eCkOb9/EXjZgXmCeygrNKaTNrTAgxmiJQSk4l5g+ob
tgHBTdU+8cSnAEmO2mOexkgEg7EuM1V6+TrcX3arHSaAaWAldUD0nfD2kuTMwwLQ
IvKPRFnO/Fcya2eArGgbU8qvaKx5DsbBTCV3ri8kyV1o8mAemQYtlwq/bbiw8FEw
hBVgN2Ab0UFGcfff6cFocKkxOFJklDE7S7BeLQFHDDF1KwGy8ZvJRhiJ3D2lKxzM
Q76Jk7QGT1R8QwMbTDqPWjC3Hmmos29mapXLyoAERS3WHm4z4L91isCSV5S8HMFk
8p1C/4/7QzX2x6839QhFcOqO5ZorMIni9mn+VX3VnLX38yOK8LUwL25gTUo54cAU
BUxoAUPsSDhxCEQmLi/dl+uMpW9H7slQ8YQla1SyIXtiSB7/m4gkWPZ/LdxtxRQT
bpWxTqRYo6V2W3UXk1XPNzssvmpE1JcoB2R9jn+2OJuXeXbjcnZjYR3nbj8a4aDb
k72GuD3zYI3MYBrXgt2lEPS6NQ1buLNuYze1D/BltBlCGvWFQwcfINXCLPYfzdek
Z+jl83DvwCsI8R/70EcvJeVjO0SXxq2QIIxn4ToOWetb9f8JenITmnCPn5mXR57Z
L9rloHMwnZp5etWiV7B3IS9cmfm27NXcmxxJGMDqwoMeBvWpYjV50lGgNCtu+Tat
sJNUHEI5p8KM4hvHdoXB844VOkfyt1iXXgnuxtMPtczuazKeYUav0zL6YWSZhM9Z
iMwoOTzqLQwJnbC0hAMM5kiOTE+ejIRYsf3tRhMEHNkPpyLp8HqXYXcaA5Mraxyl
KYb+vzpAM2SKY4cr85hoywITfogx0RrWfNlagDVXPZWXAUhHX2E3HPQsoSTy3Yi5
DxeUZ9VA10Mgbk+pdiQD5P9+UXdMmPnO/PewxQqeJy+dRw1VxhHWnpMZJmS4DaDb
K0zY76mKpGYEiGibYRs50505hbGwiUViaDAGDWOVS6v0LvaUurVerIZBN4BXRax4
HTQ4qqaffngFwGW/rb21HIrwUxLhGbGZsqhv41wR+sU+aui4OMZE+y5wSVQu6pkC
Sy3n9Y89d7QCryIsbfcegVFtqBW0Mdr/ybP4xKI0YqS40gnrVVb9fwFvk/NOxMOS
Q6K3YPzf7tNPSdhoWUAcYpQgeabLNPfOytFmf4p6xvK566IPdoMUvzHj3VZVu1S0
KIeBaffcdfJ4r4kvRw8W/3GOTYvsQBqE/PE92BAqfTZuQXJtkA1xi4pItnwke8Ou
KOu/j/lk7z53A6l5XT54D5PIKaZ6k4PjS5V9LOEsf70szMdQ+hA139MIPnwzUaCH
/j+0/tiqDjJCNKD5YO+HvHeQl1erRedOhjzWdZ1vas5HcatquuwEuwC4E7bIEX+Q
XKTScqXp0dbOMN+XDrgcGgyMl35KS0G1YvkU11f0ZPjTJdw0nbK8NR/PjVBt+gk0
npIR2t7PLQb97B9efuKUJFcpuX28cbs5WhVRi/vcgrUTIb2D9GFXYGmKP6JDFF/a
UpYcJ/JFbGVRD/oOy5jCvHu9PUQj9GYk99wOqP8HaIGyd8gHPJvpTXnO3nsEjJ45
myEuxZtuFDJA9pwtz4UdlFA4V7ESsxuWhxicTJZJcm102kM3XRGlCetMSybQcGO9
9WqJJ5Y4Mz5teiLGb5duE0imtf4vaW384ttgRp0uMQhlfpD/7yg/jTYkPNPODUH2
z6JZ0OidFuuR007arj0tsXvHUOpRqYIcf7kqrit8zdcIaBR1RyCToJafg436VIPe
iau63s3xr+6KEkQJTT+m0G86dm2O8abBUt0tjq1UVpOCbAHfm/lhGn41DQhxj5tz
/uCyx0lSCrW8GzuhNsOcBkvmGFNMLjnwtDqVjIw6Zg0rBq/4eBpvxkVRoMdxNL+K
b4FDqmFUlubFflstlKOW+V+yTC7L8ZlyDnsWsGS/L7PbT2Q5nfdwp5AmF8NVrBVw
a1A5laf7BGxRH7zxc1Mw8HHR6JRKgeVWnIF8Y1/PvjiaT1U4fKkl+IDuj3Pp5QIx
IBM5lpK/ZJ8bv1pUh1zZXYMA2e8TevofKfct/vKOz08lNH1mHUFMlJ0ytMKF2P+a
LamYPdP0Em56fbwLzzjk6ZfYNSOdO9RmSTGE7YqehGGWZUW8ToU3RwetAVkv6yY2
PbxY140tSC8CUC1pNKW36Wu+Snir6tBDO+CNQXWp2+goDMwTS6rWSJIe8teTD9q2
TRcR1CPvQjMpbPGs6zetJ92F/H9USkkPe5t56MSN1s/nOXn6EYHpcZt9BLrKCMri
fo8uuXmckx+fzovsgLTMFy1AKB4gQ9PM47Pvyy2bwdqMaiN162efazOG3mMUqni4
e8d/slgYzM8pe2TRwqITqis6YBqo9WLdCtw2l7OzblENdEXB2BV5598qlNSA1vfd
Zir0AQwxQFFm8FjJaJ3ko10wmyeITQXai5oS3sdX2EfvYWIMssJAcgjMFXEMTpUr
pQRgy12ZeT5IX6lNhIuG6Wx3P8FPzcz8Taf+Vo3ZSzJEoBgEm1RZ3t8Lp+xig6/7
3LGur/xnE9+4SuCfal5YUfCCctQX1uN7q7IWt/Y7vFepFU6bXKHXdnhXFy34mwE/
hCAHd7cmTZTr7+47M7svOr0XZdSRcX5whOte8eFe+4eJFFlVOmoIvqJIj2Xar3Ot
Z6qLIGH7eV1WQ17g4QLtC1R48VTukVQGAFBALpxgRfJy7CfX1974/l0mb0auWyYg
Owfd2liZkgkKlzkvf/K+C9dR4BPCZFHA1Af1oLBOvos9nuyJz2v0NiJmv8Ozuh83
rNv1YeDLxQ0OPetpQ0PDSZmbDX0LcR0WP40ORdvDuFDDGhaammT9e4gHiK86nm9X
aJt3s63nONPhGMnPdvHPrqIfoYH2p+0aSSo0mJy1g5a3wwDBaZkl3i3jk1v/33je
oxI0BpFflSdlHfan0kDhJfNS9owRqqAF9y/v67f85iiluaw4PCAwV9jmdSiwSH9g
iTQZGLl4ByDko9WcRzukGcLnKPPvYvO1Puk2abFVE/diOnfKka+Vyumun6xtwU4i
gFQlSXMVOCnwRPtqM2fohPPzhUWmUAXpgurzayEYYpPtiPzFGja1ruNAyDhd/I3j
ZMG24j354/pOOWXy047DdEG7bKUZGSoqF0/UBj5JpGCqi6yW2YREvAV3EpnC2YAD
WsuB0OMoB/5qk/pNbQjkEj6nuV1SgJzxCoLW447XYMGzu6fAK6MLgJFV39HILjrd
Qeus1V7jjRP07CBzfUZ0H4E+xs2jSR+QrA5t6r/CNp8kNZP5TEb3joYEpPcXeEWg
jXnQRW1fDZPUnWAxGJMoH6tQGsSVJLICT8GYPzeAXETdkXqFqdbRN1ihjdw414V+
DRLSmShDohoPClzmE+6wvdBSZPmF8x4mlLRU8iuaElssj7jvN5HmO4X11ch2rrEO
b2AP7sf5JotS9dTpFuAXRLsLR+YKKZY5dpvJRcM83vneH9HCPJ5oWk/j2xdXpZY7
bo35k8XpMpn23A8WozYYW0/ID6HIhFN2CpdOFBxW93Jr3zR8Hb/nXoVNhjahrwfr
E1ZNq2jI7QQNEW5vYvxkzyGsZ9QrPYd6+iKSchrBNp9KMT31ivnJXoOsLag8RO/R
U81+xt3ax7BcZ57IGydhjBoK0dcxu1AvCwVKYFO5kHRozRMIik8TgzT8QZL2bhp8
vIwttxYifruVZViaDdxkvyEufjvkR1cR4SaNXvrel2nkVeR6QHyAoeu2tIpt+WpK
D1YSf1SJk1UcyMAlCENlF4iftIjIybz3zmRpD/VDlbB3QSS9Vqw6PHUTDm4fVFrV
gfsnWh6/ooBbUj0aWzXpVnR1Um+ekCB0j8HYgdShQKYK5Z2QwXrJzdQq/FV00j2q
TiE7552EqkvJqqwDtmzu96u/r0B6xaHt2LZECRCk6X1ctPuM0mTVx5jYuynR07Wn
cywBpeEcpZIcExwbI3jSbjru69lxboiitQwgfBZhYPZEdRzttT8905RqfDWjTUai
le1Gjvdx8cjiznHtrg8XMmTOaZR5QzEfGB6MgoUYcYmcIyTlVRev90zq0Z7z2+Ks
Yor7JRSxdGyajhbV303xf1Ze04Zty5EZNNx5+Bg7wDMvPF3qCj6BpqqI6Hii+TUE
bD0xUM17Z4PpH339qkFk3piaxHqi1pJP7/0sGsAhv2K04n2VnhJhLr8wpKRUem/X
xDpGjiZfTQSsTsy6zM/xFV49Y2Bj7u2xuDJNQq9dUamX8uz/m0FwP25ECPdQe9+R
6v5WcMLMTxFdLedjaM+3tzdvD5LBoGs54xFRs594mfhZ9PcJXIZbfOmN5DcjdGUq
kicpZ/2XkjGHXTP8VCAgXp/O/qxc/TS9HApzMTLUJXX/UZrRj7oPx7x/FSuNUcLW
v+zxGJv3Q5I5HwJWsGboCKlHiE++pDl01X3rfES4Kq54vtJPDVf1ldBnwTVWmNq+
AGM0c7wan8/RwYfmKx/ulD4ZgxEWEZqa22OAMWgB95l8k95uH7tWj7z+WlTsrfrz
PVRQS0zLrTJ+pqFC2AUnmCvXbQbcfBE34PrP2eZSWsNGlvrsWmlcASDK5MU5jtnE
l/tMS/qIiz2PegDE/dydjHvFu+Jt66eGfdq750YpabvgMxkDRlDr5we0C0yJrQD7
/QHxhoorlWxppFQr8fFXFWktHULUVZJK8aiOPHkzdXAS3BVtVOQuIg4fOMWoOYT7
xuvA3481jq28V69ePLewqGiEEUXxsTCTX9jLKIw79u0keyKKnmWMiDCqZvoN0rsh
RRYt5hObRWPxo0ZVV5HwAtIPtGE9MnYuMiPe6PScvY2OwLnLDHsAOfC4cBN/eCac
hU51ncRPyvrTwS3Vkp18LtxrbDF1SlFh2/warhHM2HoAaRCdC6T6QCZDF0qfOlk4
mKa+vR7pbq8R9IdpnVSD/MGUlfvThFWViIOsD6YCqgV8rrZsX50zq9lXykBDkEsL
IF5qbJeCVnT025dkmtxticW6+CtlDvfWq/KSCy0oCE4a26FteMH/K9ExXYJmPcH4
+NmYT+0a62frJF6N8eZu0VpsOMNqXCnd8pER1PyKmfuDiZG+DBj99PC+IcSevWCQ
M4siLaFGP/kqA6uq2EjvrhVpfoBv2XjbiUBoX0c2XVlv8NJC7ZUTi8Z6uJ9CXa1i
Wsd2COBzmvcLKDKrPGUTNy76R4suPWcE1oIOw9mC+Mm7fwwMAo3Bm1k/0q1Y197+
f8lFFVJ65mj/y6hasWa05XIbyXgjr7sQE9640ny5OAGeNgJb1mMPIM/im7YM0Gbj
hiteetGu6eF3eX52sbBVvTuyiT2D9d+zlpPnhSkDykQzh2GV0OWsIAaK/IUZHDk4
UMOHENNUjAQWsFah1I0JTs43v/K9mHdhIZqznJ6uMiJDaVqbETTvrnYI9SuBFn/9
RGoQZAWimuDbL78LJLDK0WroTQVVYxBcD/enASAT/jBKGz9CNzDQOk7DOVKhdTN+
1Gg2BgVl6D9etIiZki5GENoQuWfWXsmvtDbk9oNBC5tO++ON1YOkyawQV2svpxUQ
ndobdjSAXLiDIyIxG8ZamX+dYojrKeSBn8/ZZ/2pLWWFtL5W8Er+AEJtaY5TKRdE
rokBbCRiL88fznVxXU0MiLnAoyt+Ls2wvHh4OvjWNhsT5U476N4Rn51MkjURZGWM
mBWFIgL8wpef3aHrRsiVbY3eSo8sxxEfhc5Zwk4nPSfn7emV8BtrAK+WbuFKaEN3
nul3S6BQHktacRbuULTANlSzZEiX+HUiK3EIRkMhsKtcFVSlyAQLprzVa20M/7yb
n72rb7XCUS2MIchOjqMdPu9TqXQeg1y4XddcfXRm91DKCE0EzY4aKf1pWzh6Du9q
fzAb8AFyrxuNNx1OfYjzIhuy3hTdzz7jRbSOJrDVtDn8GECPKwp0jnGsfWXPkC+5
PNPiAIpkIBIuISwnmr0lNa2zNPBeBhrGnPPt4Rp1gP3N1mZfZ+weUW2970JyR2ki
24g7kDk0B7Y3L1KYVW3RLzZckVs3VJF9igh0QI9OsX6/L1fVdugBGfQL6bwseAdy
faoB2tOsLADVU/b8mMpyFAg/DdEsZfL3bkGPWmg9NUKtq9g1SuLUl5yHtYQLGFAp
CfYgT9AM+xqEXk2ZFsleCM8d2xwZwqj/3mt4IDc3PVynRxFg1LR+UB2c7Vka6vlZ
fdx/dQ0vk6eyHPezMmMx9BxqAlFMY9ng6eReBbAfJWCdA0r3Kzjgjsm5fE3saTR7
I2bJ1FVEz28/xxvhXcJ7EYe5Ebrl8XjqZ30faLSkTYLSz7K6DKAf91cOdsg74TMe
G1GeYS5FJhvhjpa8MzT9g8W9t0HMchFTmB5HUUtSOjNIob4//lDOsJWI8+rWChbl
58flc0+oK1ujPKvxlRkbxq33btXeVS0IgaSrfHAffIuyd8WACSAVKi1+gp/MUkFU
mBOKG96p3NUdQCcH9IgqMjL6Hxy0ROkuAe18qSXOlUNpurtPWlCdhh9kRSqJNwM/
1y02lywQZ/ORYJtJ7z8k3560Bv8iM/AOGo9fcilkiS/euES9zIv3S/iXKudJuaZH
Qw2HluKisFkUR8QabGEb5m9SdfOa2WaB55SrnvgWUHaFf8+GB7kSbZz/TGyh0xVx
Akd+OyyAPHSr4OiDzQYomXwMN+9mGG2o9QKlSOL1sZ30ZXMVJ8jFLsklD1ICMeCF
duRM1LX73VqHeWH6aWAQCvj8+Pv6MCreOQj2rpn8ccstO9xqfKZx0PuNLpgSag19
qT6tqfRJwptYhFvDTppAp/so6Ajuud+oQ6i+B7xVLMbaA3dxv1nlmfAlO682+PmV
FXCQHQOFJyIrLQPOTpUcD/zQicGSG1xQ6zvxrFbdvcQPKfDGj4jO0dF7I1UiU91i
ZqzzrCBcmNBoXaA7pzTG1dWEbNdF75PRhRO+bgmvjk2UlHg+wikQ6E7wsPIu9AWy
baKW6TohnhLllYHcETcWu/rHZUkwCg3C/TPh+TfP7/P8qWFg1fRSdJxFpxwIFYlX
h6kUkgbxMPxwdClx31FW789xwLWJHLxG3/R3FRGK2ncoa0yTyZDsc0jVQGfpyN+o
bf0eBvtjHsc+WTESdS847EZhS5I3+SWOuRfKw7z5l6VbE6rs9Fe+ITxKO4F+6aiB
+wXQH8dNeVurUlF9p+hojk+cJTi4O0Ny3iEeeOW+Vv7iQ9xOvdeY7YPf4T50lr06
vOd8T74IdmipyAh2tzrhyKqE9mamBo9XFZi17+S8vVxpjFKy/VoNQQn5Q9KRTlfj
943coVCetq26lpDppjV+X0UVh9J0HAoBAG65cid5dRU7Cqo5rmZVLdJKcoYrjmhT
2it8a31bKtFAhr62omG53MqrsP9EKm0JVjvbsGRbRzxfIsvSwxXNzv01/9f4cN6m
ksLWCz29AGBFIQqZs42N6PhjdDJiO7FVqj1+3vIsZWs8YPtzuMv2N/xzBUfwzyFl
xjYCDfgbIiXyrU8wVdu7YTpXRG55KYwG56XF3xpLLEuVWyfmQgedfoHGUIYlDC3O
XYHJkIHo67qmKpQxxVcQGXs7FZqpZLr8SwUVoDhZdKSYuEZnYZ+VfK0Ygu6SFtDH
iE1d6zuUHp6kAntIdCMzmo8JOt6BPDtGqjhCmbm7rEcwJiK44vaCCGiIDmszXTpP
dpqzrF1F8aaPuoexLXIndza0JOuhrszcPlsJH+bdr3wdTBCFr0oQBwYwNTW6W6N6
FOHDh5w0CurE+Lk2Akr/qfvZejj5NC1TzpQOsxc/5Dg9DoA/vC9taTGRWQhGc5X8
aG3BnqODfHzZ+eHavhS/k6O/iVA7lumhBI9yjwBMPAj3L8m9QIc+cy1ffIEp2wQ0
4uhojdKyYjIZEIR1NH6WUq5OLxSGzrRflxfyOAjt5/mu4rlERU6pFQklNltZ3Wef
mfewcZvkDpX+U1t+2QZjO+HEjb7G4xLFYZ7XJYZng1N8Liei3igXlzXDs/7T4gSp
OW5+x9JC+JqNdpyEVGii/L8TSOCiBnWBban5B0EOyM/R9TjKScOjqVVARbDyWrAe
DtCJ8bEDr2MCmYGy698kc3SRBW9hBqQ6hzVztT3ev1IseVdRo8StexTUMSZG8Gfd
R4DGz8AP81psRs9IhjC6tjwWtQQN657gunihfRvDYgjRxxi+BW2d3mM6ZjNu4KU7
li9s8sC6IxUCGc256RXqrkzT7x0RAJKvGC9kuVYqlznRX6mVFGfzdEOUSqOXbhlW
mQC9wz75tfGxzkCx2ovHS3zAh2ah9k3HG0WrD45UaFQwkWYOwkyowc5dlyhDTpS3
lAEdPRshkQis50dapiB7ZliU1yc/Xt84me97Gh7SBjmkAlWPxrt1nOPxS3mt96/C
zUrnlMoFSCHkiWEcZ9CbJFedKEvP7nZMIDeqUmKYhxezYKPjJ2nOO7TXZVm3VVTl
tIoSWEj36w39CsNxXRSJC7Z0c4Z3GSpUuy8P8vp5J2Z9ac/ZSCG/vSjz0d2GV8Jw
2SJsK4kycgiTcEvz9PVzCfwHS37hrzmS8s0S0KtV2FTdP/I837higstUFciY9LjE
i3sgxTSzhPEt6QOx/I2mtYYTEDq63Ae0guQtNr1QY4KO1g0R1u07SPUdlwibBZLG
me/ygU+65ZyA91qOLCVoh6tyqsZnNHvwJqiafv7pBo1vK6fI4iiOtf27ZzBrnR7n
4sCH2LcMSjd+muNVtQggcRLwQGz87QJPwrUrlWLH24ww2+zm7qhkHeEoAkNxonFS
BywtikI5HEFl4CrYc6WA6kgbBe45Bt3hyys5f0Azglp51mtiAufWPOXUUySFCJ/o
atqE5Y2dPvwqtSxYkkpb75Zek3lQlb1KCWopr5p/8wlZKJRM/X6Iv0z2xtAXUN/1
h5HPyiRsmJZ50PqMZauBrGn4DHVUrXQ1r6EXoG5yHmwPonjQzEmHlsiVpoWM1a3z
Eayd6P6JvOCNNOqyhgJzXo/mbTnf6oVmzyDzs7ruYnqLUL9ed8Fnax6aHR2YsSrz
fd6B9BQcQ4faWiBzJoxePq+7a1eZGB/8YL1M3d7tgxkVYIE8H7Tzdyxie8ywzNJy
X4/k1a9VnRDC+cnQVxOzRP5ufw/5JYXmOy9QAVGcH1KF3bfb8gKTUtAs70Z3Zc5z
hEIpMLehgcSrl38GPyv9y4xbNFaoHluJorUKUNL9wC9fUcBDeVR8dE9elYUqwp5B
hGkTPqIE1lFcLKc18MPqn1LNoYUrDzyAPSPf9eKNhfIOQrR6FiLhezX1jS0cDFxp
P4d7kI8dVS+fOWDTV1ve3Pa0yOOiqlHy7BYfdakWIoYegoCD5H60SGaGpVDLr+gL
s9n2zp64gnenFKSEYp8kP1Ul6WeOVQhotnBcpcA5/JdeB9ES+f+iQUU3QGyobljs
cy529m6wg0WB3cOxbQ/y61n12tnPq7jgZEVSjxKa+wDHHlNfF07CB6oRhGQlQhoO
JrLY0g7p2vq52n/ZoIbYTCl2I9u0V02a7SDIWQgfBHERwTBOrRq1SVzrz4kGT+nQ
+e33IqMLXJlEDtcY/is5bGZD4D8oOSnzNzH7qXtMwwQ4xf5p8ap3kUz+VptL+s05
rPXm0C6lPYJCMlCHv3zdRVfUAudmH9MtnzXUDqLY4bNnou+Fo8exfV+TRlI4LC2A
eiK5uzdSUotNnMbKeg5nCZdG9yN/9TzOD+X6tEkTqTJ6baoftvO47wVirwZSESju
HaLDGRxNAUNyKzV2D2+SCXi9eldog/xJt84dlIVJNvHqYu+7a6yMJKAlEK/XIzy6
yzQW7FuPPf+BozjBU5bZHhuxq/0TXAbKwtX37roVhbLUUCQUoy3ajLEioU46U5Ed
wZAWZ1A0/ysbGIDzj0Sb6+AJhyb2pOqqdocoLvKi1/D3ft505K+CT/UNn8h2aOq3
7j4b6X8xmBOQLfib0M/1vzBjBWXJljiSwrjMVvq0fuf+sRHWz9cXmp+wQzQeuUFj
n39hblPC/07xt6rdSjNq/edoocpGIgg0d1EZCEBDQPDJwsdvkiI1A4PZ7E3+DOxs
ZzJ5My4EGCtuarbF3cVvkauYyJpmNTiWicOjxj0ve73FG2c7A1eAwWKky4hDeY/8
L8iWic+Q5D69g2eZ5y7Az4yvo6tZ87PLdzEpRgnPXIgp/ARJDd8S+rTlipz2iJki
0WJ7oA5/DJxxdQNep1xUD7BTbSAqla0WB2zf9DcI+MM+1TOIxjLUO1ROJjPXV6i1
JhylaAeWfE6QgRYN7zI/uFWyPODsjAh7zLX/g3WbfDiS0QwnOLjT7yzevks9ipsF
lEU5WrCtapNWCHEF8iYWR43OA590OQ64odgAwK7YehXzTbF0cw/EGJp2JXEwkQvU
AIMKvHo7wss8KwRZZewlTfEyM8MKokXtk7fMa7ckobgrW0mthP+Lhsw1XHupkwMT
Gz2QyRcsRctiIuA4xdstem9oji+fKSiGR3CCCQcZbYE3FEJBjJd62/ot7v+FCMBQ
8qpl06uKjTN/aKVm/zVfo2+rNt7EXmpy29+AvioPrmHh55ThJhP26Zz4/df1TG/U
IjO0QT5yddWapH3BO5qwUKdW7oltwlM1+j2L9FmofhzZCDJQ90HiI2q0nUPMwxJc
1wekXa7EbJFNtE1w0rhxSo4Stid12qGMeGzriN4DXIxanyD6MFLXM3Bodj8eOO24
fRNhnE3VIInDhcd3b14D0JkeJAyT7DWVVNDdrQ7sngWWQGQwtckMR5MoP0ZJwWT6
56YMLqMyS3MOo8U+RdPYWhXwEtKEUF0F51ju943pfmERP8+VRoCKoXCu7p9Aw137
JDPYJu0s7x8LSvFOGlD66uKyTPzxBPMgRN9SORqEYVFjI+BLIYqPY92yXve9s697
sI0+Yx2xtBPdf2s/tfR7SoY9A8b+N6+EaygcZKTTjm5mYN3YAdSc1PXTIHQwXqmW
As4v9N49eAWkoR1R9q8dlCN50nv4K5aPNnA2C7yd800IEADzeyXVo4v9AAybs8E1
8Pcwos+2csN3ilG3/BI/WBhkbaNrtf/ZMSuxhnMrZW5zG4Oha/i1utZS7HH/J++o
ViCIT2E0d2PGQwIcGrf//cx6jH22obBZhJaNw7pXW+9JjeZaWQ2x37p2b750vEQ7
MiPmtDj7GBRYBoFiV7cuZZ54GrLMiUM+y5dmHugvLlb0CoJuWRTI0mqCWqYh27a/
ySdbzQd5emNuXydBTsSkr7ouISjkHHAdFVotp+yOhd9pzEcs0bE2gWGjw1SeqVe6
fyGQGi8vlTCeD7swH9PA9gq9VlWzCW3niOtbyNzlwEoTZIf0rn8fY+/oqfQTHowr
AOuNR6Up8bmf5ZghIZI9scQXs+O0XlBs+CaC/drO8zCvWz6VQUJcoVDMc9P06uGA
WrDI9GIdc0a9QNHo1AmxGi18eEcnTqtU5iw53IlHHQzFGrzIlozimAdNzVxFGKOp
+LnWErryEnVXB+1O/iUqngk/2wIvVVhXSCiR9OC+y5pk4uv5B09YVLY3J7msuMvO
YSJyOt5M4nSHN6eYz3xsdr+SXHu2s7F18WC/Du4tcZqfyOmvk30N0fXoPu5q8Ioj
g5VbY4CHw6qB5v5a+MG8XNGYHGxqB0ERG8knzGM9Xmw3anp9uwcbpw0nZzfhF/Va
0CNDEyNtD3KEx2Sq2rqqYT5X+WjhhefQ6Kzshp1ZvQNrph+wUp2Rd1rG1GWF+qNV
xjZ5S/kvWIwMCtFBgg8+TumRrH65MiRlMiZLwEMU38fmT0U3EZD51eAcPXTgIU94
6CX7zHNDCddT1ZValam+xf/iW0Qu3W1q49fegewHGuVVXBLqn08jpg3lAiwHcRSY
8G5qV69ETJ4QwhfQ4pcmOXR3XnmmHuQZ+qbaMv67WQlwks2V/2PDzjAG+BSd8CGD
vJWeX1Y2iBRn/xDnQDqneYaigZ7etp1i/0TQszysVvvtsBn6miuF/fxvIhfabsBY
mRfOhq45VJOTDlhrB90fmd0x0TX8SG/O2faBa8LMWuc1j+4/XgdrK+ynTtZ1eM8B
cBAabGRz3lOSlJSbcTgp3qOVVazOTHyG9fwxW1yWZvLuGn50gwYgnTu34orPdAgU
xq8umJbIZGlb26Xr7q5EQh9JhP8AshDqU0nTCQ0N0GXUVb8TYWKT+XOjvkX90qDI
UxatffW8cSbkBjgzSWtfYb3WafsYh1JlGzo5f3Nvlzc+0y1dvihyoa2hQlY2WFpQ
rOdsZtZKJ6VTBlJQuVbN35mo+eARTORck3QwS9RnehzRviwvL7c/1/fapHjeWHkK
tinZaPbGXnqAtdY/SQKxUpO+nwzZ6kW4zPkz5kmU91kfJlQWaVoLh8sTAa95vMOn
uo5+xRSR22o7sGqjF+qQJ02WxvceL5YG6Ycl0ZDBLPHa77X8nLtqWhJW6NTIDG6k
Lhk9nAoT8VnH8XVTc8pHR2lVu1hOTcZOZRdJytkgL4/ue/hObAYD+Ww8WfE7p5wD
JTLzML3Ujw4jbJjlTJroBOBtjLDpsKdLR78dPg1EcwdEE3HZCfZTOhT9frTSL8Ua
d2H27wZVALQjJqpegaoXqOMqmARi5ki7cEihka19EnY9VxcDJqXmZsrj+KHu4C1E
oxocPpi420/TqK2zYE+9yg448nssB8KIJqlQkyMbexhtR2o0JupPROz2RlggX/df
9uJfnv3aENNwi60vZ8TmNiNx/XEGKpISvCM/++xYuDgUa4zqUNv80giG9+QQzLbo
uWsvJZX9I60YRkM22AsdPIBUp+rt11mYeAtzg8oOtTKRAIAVopwMwAfumyAJGG8u
ThTZobhV8grXiYyd99K8eosB1T2KC/PnFftbCdGNu6/D86R5WRQHH6mkPvXjAeZC
knNnioEx72Aar1DL33uLYwAzodE0VPLozQTQvV7TVg6bwqGMN4yorLKkAcdkQC04
EjAM/1Ftq+77/2Hol/AfxPbVXDKB6XyvKHtesEP7DcY3pZFXFmznkh1BxdG7PkUk
I/f5XV46MevmIr66HGrPvSH/LdqwQcaqTVIwFgr+Rzjm6Px17tOP7QVa7YMB668c
3Wea/Pst/TWz9YAkZVXE/dxCO/hX0VNRD4LZP81b/uLkntoPwbukiwwQO3ATdjvP
A/45jJeYiHeGJtokmysl6LSWrRt1D5z7GiQ/YJDP9NWDloNX5nqyeOMaWnWCQ54H
IY8EY++HaedFf306LXNOQS0VSnLihta7+ne6kTBZ3nsRZfKy/9fYXNqhSYlNJsdh
DQuK7pDe08P4Y7dHoskPC8jvf3x98kkPq5Qq1jTPDc0BV+oxd6mUZDCBaeemunKu
SEyZjbs/SA5XomLDqTcMYMGQoDQFxVOddYF9VI8sq0whBro14g8b7To4j/9lp0gS
twkT7BswwQQKJP8Ioy1rsXqw84tPbOCGT3mVF2+vhP4fIQa7oJjHAgLU6sbha8OO
YajVgwRMcWb+WafOvluqUKO8L12j+e6vTgsCMZCmSv43F8NE9hMiJ/PLLG5SG7qk
pFuUa9bg8ys1ltd7ytYMTEIY1Gow9heZI12zenNdhHbyTY/EkJPCoblQ/JpZr/sb
LMu97U764aEHfNklwhts3qa7Ri7h3OPc5yFazooPn/kwRR55KGawFZTCYYNvrV46
8BObvZStx9pfsDHy7y0ZcKpBoWyu8YrkHzlTMEYI87QU6LQ60pM14aRHTWgnrEt8
HlZYKMQRrchzDVhuAxGytzBa1B8ozqO4y99uuggfWh7+kIHX2abA97dN4TvgbzB0
vsqki3S4gk+MrMRtgACMwPByUBe5rBdZz3s9LNYzpOy4zXPeHN4eJ0N0Pt1SXImA
aJdGoiqP1s1yESSndMSYzLVmVgo9jUnNr8ydPv8c9/ofAMOkf6C59A5PAuiCXB4N
MbKDh27hIbX8H8IopJebeCMMp9utoQMWlCu1fqXeb/lE0Pt9RgWVgigA0XMZpiNA
wUcirlamNzhra355Gf4IkurPIfvDjram6Aodm6LDFnMJ6RspaG6RWzR9nmGTd0Jy
wpU6M3ycMYR4KtYGhQfzhwkWbyj5uLDHfy7iGnjiF8rrTlquGHLulS2rStxNao20
A/+hn3tfkTc3v2u6gqAmE05WOaHH9Ew19a9DBMnYSlAu3tBZY33ar8HKYbXk3gV+
tf35ctK96OMvf9W5GT0VUhD/nv3LEmGAPiTCGY8opWujc4S8y+0+DQmRXjzO3wda
hRF2aKMSZxz+2U+W+vxoLuzErdJZiqPc9vQEZwCzHHsw4mdX50PZpYrj8ObcLvhn
OkUclZx7Yh7ir8Kb1dRugG+XAc79iUXyt/XiiFJJ0DPnBt5TUPDeNexesU87wwM+
nfVPoCOKAnGliinkoh+Tmjwx/s0NYo2ykZauLoDvPxn3/sIXRgdRZddVHxJXFPSk
vGVpqBsfV0L62uuIpg0GVXP/Ykb4y44uzAPrQ4JtQ+gECKKwfRnCaY9N2skfiVMj
pOrXZGqoF7Gsk0OGADzMwTJq+WwKkyTSoV03D2/t/sHI1vbtYHZJd4sZw+tgZN8a
+GMOEV4khH35fO1z6cJVh3sqhZ56MO9fWRggxLtoZmH81VMU15RQo4XgesEOEJdU
19IKgM5vtFcumlEA4TmvTt7AiRFJU/sJTe8cQTY3whdJxcNTRsiRyF91k7jX8A5v
vtwhpN+ZF/fun3jjla99XBiNfZKxJ9oEViNbQud2UfFP+VEAFiwcwEgXIPfYjPPW
fSmmuVoHD4/pF/BlMTu1fwurIenZhBaM3nu1Ad8gNersRiuD0ohI2rCKWQQkaN9l
V1X7oejMhI9j0L6TMv70fIOTsBpWn68Bc8tGbUu3wysWmB/DGpih5yPiVzKRYEa1
gvFs8YqKCNs1JjbEa1Uzr+GQVLsXIbx/sbaXFSfYYBFkKtRbW47HzENmJaIeVdcd
XDBQVOnkq3EdnaTpdQKivsAtitb2M5zFyGfmvE6yTo8eH8g56tmuS3KE+msmkLvA
4v4Iq0a8RNpWSrokN6dkXCu48E+0UWIFfLwfmuRBaA6PhtIquQg9Pka67OXyeVxM
4qnTgHkchIKfVf9orJTBsOwGlye+wvvOf+sDrMI3Rd7N289kEizyZhEMz8b4TBJH
WTQ0KsumM/tLDVnVBvrL2swOfKUrKKDb1+MTdLp5e+b75iStZYfBODWk1XeMVd0V
38Dcjh8ymOmj76EQxEcQgrV8GFEtU4EETQj8FLo7aQyYzgj4+9jqdmigj2JnorOY
ya6G7IeXefiEiwzx3JSJrmesTWK2vgc0b2Pcd59RkQ81ktYQFAiOQZuQH3t2IE4o
16IrqmqxDcIg5NXah3eFh+RlXY/rimpGPhIo1RerSajnlFdZrHCkAZVDlyk9HRkZ
rQ2s/0l6dfJXYTY2h/0aPt/SVuZyqm2D5cTe542Q6YoCAiXvIBLap2hQNzBt3oRY
mPWk2yU/l5Ui2q4z2oVBizd2xxYqRPJx1K0/0gn3b95bl1/MnQ+u6Rdln4n69m+W
sdfBupf0LsGiFegKREGat4SBAnYj31nJd4OgHfPeJtR0ELFUaYnyrj8dRT1GjQSs
FfugNNArnBtYDfvYi51RIToR1y+Y6JemFZJO5WAfKgMAR8DmPFJ1BWOvLoh/jzo0
6FnK2DHMuh+6EM6kczTBW2LsV37WhXetxGZoOXXphTg+wIumjJ3yA9pSnID1lg+p
VnicM5xR8K7TUqlee8uB08femi7tdrpVL6CuInds+bW+2v4QM2dNGos9A29VvaPx
2rMTmxaElP3pimV38LtRGcaTVAYMbdLv+qmpcRU4Mj/R4wmQiRu3sqdUgq5/7qcx
segKqJ9JLr2BGxf+mmgf5RGqiph3QGiL+Ai0q6+Cvec0dwb8HxVKMl959c7bIiM4
sRaSZE9vtueNnCalCeK09dDRkvn3HLKB2mbBXK9foRKUrp+Cbz4LLhJowZtqgm/R
gM3HsjXewpXLlGg/VahHQZ2P1dOXeR4xcolNCzBZL42TMUWTS14NvuFd0IoKDl33
N+MeYzmiw13jIXs0VIKiWWRaP1oeAwWLYBxJAghnu37B6kdc6Ykv11mGKjvOFY0K
VZ5Kvbk//rNjWcDxjamEq3s8gR7rffAc2f6ugFMBYyFcLHFmm1PvTcj4ZF3Imtxv
8O79IENCEoa5nGWzpiiWT5K2Y889zpE8Uz3H6JSNVKzO6kbHuQ+yBwW89iY1UDw7
ILt2XOzNeTIhnMHH/SZ/utdBPkfdY1lHi0SUNnxdqLzIOBaXcxpPreNAJ35VfrQG
Iq3RHzClDmMZlILlhb0A+cLGew6aggIMbsmFzvikmBdbuxo7IWBOOzqFvwy5FHOq
hyaiOSaVD8b4ibVd0yCun0YnRQcKWy3oNZ4Y33oFlzSSfhu8CGG4EfJF0zKLMBYk
3hdzxRloRVYiJkvDV6szSTNrVSa1keoAECmtHj19BnG5ElMJu6/F3uhgsfZS6W6t
sOTOuW6yDp1Er7gm6ogtL6KNDTU4zzy8GxnLPGL4GVxhSkWZ1rEGSfTmLyTHPS32
tGYUZVmSVDvlcTZlbhLkYXZKF3Bf2o4kPJP5gtC3gqepbw6iAlpW48pbKSqDhuvO
1dV0jLQZp7Ed0SSE+IO0kDhMXC41odoC5NJ+jlNtZrX3PHeiKVXBPVuTnTw/fjZc
DRCyNw1Hr/JA/ZL3KKCNPG4mDamfoXPcXHkjn280fyCw0KKa1HyJ7f+TNpEe6BzG
H4obyuwMuWUbH6KRRe7FLXu8u9bbtPhH62mtDgQKPc1g9Bm2fKNHpE5pZx2KErTu
e2aCnbnIx8qnps6yxZa43e7noHBY0PciWh36pxDui2EcaUO7rCmWHQLYYGehjvdC
sIyVsFDLn8V2c7kMAJLz8qKadLX8ZsA9buLFLMqeUPG+CYvcY0+mBYcNhSpIN6Vo
uYLweieJ2x3McWMWbKbCUXoHX9MfZDS/vT0Ah584LaVcAkDIrf6pQwN2zUBDURey
iYVmA1Hg3zufgbwhGj/H8mKcj9tiF0eYzCEJ9hWkrtEocBb/WzVrSZ2NatDA+ErD
lN/5eGARvXSHqzcYLYbomqYpromGh4XXuWEOobbfGpl706czebjNgDYPRL2Ht2oI
4cddbybnTjKi5/QiJsFL1R2g+a6srsCclsqmUtI82cNeqrrdP0U5t54/OwLAVrGJ
v50jED6DNDCUc2hIff7KgwlAIHoC8i6cwjjCYAMWBXPS2YqDc08Wg59PtAM7SPo9
YI+krP7nqgHmCApfQ7u7/6Mw/5WJHq7sllx4FWm+OPVqfZe30NiGTbtNmFL9CzRM
MhSkyjrUZNgQa0xh2f8XZqu46RjrL1Z6/4fkYUJ4deLewvJRa+djHheWyiGt/FA2
Woz2zzj7Eq1Z/J7WyZZz4qMJ1INuF4bt67NMkLjSoV9KPycPHU326aBiK2IRrCFE
gx8EZDqAZrl3mBB5Pr9/RslEYn5moLTdEsxmELQI1p54O7wbVSJsnndLw1GmF6FZ
a10xT38PNY2z8RoMJ+tj6n3JFCuMXbbQ0lNN1qT07HgxOixz/3phNlmOcsOisFsg
YrywIFpCjspi+RJQCVgrfFFw+CCw9jZ5y3nP1Bp70H0k765pS5rdTGNJbdTucW1M
iiaRiXvsSFk97+wg32inAjkem7b0TYHzhLlUVod8MOqYGXxeS0VQm7MwSRWdsSbU
MV685FnoORu/2OJ/tkb+uWkpkcwKv97FI+OsLFuGzAFo2J2zhn6b+5Zh8zf2I5vy
qezjf1l/vJbU6VNubevseo7Y24eNb2ZdZCSulYozjlu8PAAc9mfxA4P+EjDzULjH
lhU11NTWj5HJabVjOpaeWz77ebXqpxs8VvbKoN3HODO9vQjmLv1L1PGBTKaORKYo
E6OTLfCBuk75BRhNlYP125c+otBTesv5XiSQuNYoHCt9gBM1a75HWvQcFBZKG0BL
rwuD6SKWkH5a1LaBeV/o3XYKkyuR+9FrXfot3eo3Mwf+sI2usJHgnB4+c7sjfTS2
B73wZHLWkg697bH/W1KVIg07/xtQy+7ixoy0wyIadLRB8ZXZgQE5Zfmjv0iTRCVy
El2CdDqhkDkMF5ChB2GAeyVqvGj4X+o+Znzqj2GXFPV+qQCZ+7HAT+wE2CHTHyrR
Mhtwa7Q6DoJxBCxrLh0uLc65XlYdfV72ARXV14lrHWPC04r87C0fu4WkMP3Zy+g7
+P1pmuDQahcOHzXKa/DghLbYnSB7GWqc8f8Do6nMIHl0eswfcqN3BGknZ3Oxuak2
cEBcyFXLX/wogWQRmkr1f84ufiDZbtAvRpFQYLYsL+1QiRJC+ZJoDs/XKjgs6OEu
kjeINSk9pCPIdyjQFZ+vObRM0GtN2lnYAa+B7dXF0Tv5j1ANX2CZ2KOmGEsF24pJ
HhT9DvbevoCIlWVh6avVlAjB+Wdu1diM0xpabVpP9QCKQUcU1ue6rbSuirNZtQ5Q
fCc5R1CnV0/8VUVfFO5TXWHDKxWbs/bkDwJKiaP0xhWDOLTbHoOfjzvMZZsGbdt4
rB2O3aClMRzMc9rpTdtEbT2erYQtQMzLNbQtfNuxN4HDN5TP6uB48Ngjdgw0911C
IS3AB63xNMhhHnLVJgqjv0UHOobqC6fi3wdHarq1UXY2Xg8IIjvgmKpcuA3BAMKc
Y8M5E1PMPPTX3czWCDgM8g9hRZF+1R43Me4LIBwSWmy3HHHPGmQwhQAJi2T7EM4+
qdiFEbI/tLTa20vGWirHQahcILEbdV9FGzK/7qi5QkOC1RswS13Y1ugmxGu82IUC
bYmoG885kQ4VPV9FI3bpkPO3sZ4fCj8Babi3Dtqe/sy3AoYKWR5YDtHJPaY/Zyc9
6WMRsP/3xhtTOstFhjqPwT0ludYMoc4LOrbDeBu4Y+LjzJT0Onq7Kz03AxhaM/+O
0SR8DbMJ2Wn/JjLXA4788aF33Opr900l4UJpeSE5ux0xxIErqJhVJRkVL5bTpRtz
U3FW6KyBv+CqNikfpcgDttCoZ+xaC0BwRJYlFe1KSVScP3Y6h5l6nNpAu9fG+2co
xRmNV4N9f+K+Qh7zTI1VpjRqKOrUNpeTvwUKRpv2YHkL1xqO1mzjaO7CifERefJl
Xz4tvivEhSfgm1whv07QmzrtPvmDRjJSwQS3uXlSZUKk2LYXm7/Azrqq1EK8DsxA
6IseGN2ZCFbruXBVcXibuoqlYBvf0JRe5pv/Qq7qTPomeGhdcJGX8ec4obcjJ6Lc
9BSjPudGEd0RAF9ozkNV5LPUwDfbtQ+Q+UlcjapCUT4irYzRX0v/QoXD/v4H8Wzz
B5C8Yhyr3qtwW+DNQzKYRMAQSCdLpNx1X1Vj4Peqwat/2dlD7AWHqoT6re8p+5zn
qzRew3f3ykY4YkacFPA0uN2fnO8PyUz1UUj+muD2J4tw/vhN6huX87PyvyPppwrT
hYIUQQkhQKsN6yIC/8xS7eV2aPTIn5Ks/p3B/NUTRrIwaktbcVSHy/M6AV4iPTyI
ngltOuBTA8YwT3nTCMn7hJxQmQw+BcLpFkeNxljf5nSFJmllgOsjNuba3e8+QodO
w0b7jO4uknvyjLidG8LCfRaLBunhOesmQ/i8PDPe8F4IPogkNRRG5MAIcNBlqCNM
n9Qm1eISGE5sziTZ7eUiVuI5zviEv1JlW2HAT2kcIYbMqtcsyAXB4PAurjbt7BxA
OVpfBqPQ4wun/wVMUaXk7Hrs04A9RBscrXsok0HG0VfjvG5qVwUr5jiEZqF7ZeAM
PbxkyYPNyPL1d9I43EIgi/GzUqL8arw9w1QMDtyOckihhgQz6xzG6UW+/CxNYvr8
loX/sTb5CXzA9TRuZ6/rf0606AB1cvVhk7TkcXcSlsg8mss+ULy9PR9jw7Sp31ME
uX+3cp4qO4w4dSOcRZMQ6E1goGQp1k8Z/tXF5WgCTi0Qr9SnUV6VpR5hlhI7Y+BX
CRLOY3U9XJCE6pKzytjpwqE80fXkMVwpJPINvDa56UJiiz8IHQN8Tr9IxNvwuRlZ
Qjtqk5rmBa1sxa3VrI8JlxDvGHjewcWDg+ZSndtBkSASpfmoteP0Xz6uGCaGsurm
xudTrBvN2ytHgW8SzqMP26uAA5GYAJPO7DKZ8EhrT92ZtiNDiQXy9x67WyQFrryo
V1iliueR9F4pCuQoaLW1RJaS3d4Om7bgy2MFMJLnzMNYHSv0r2XHiNR1FGscAl8F
abFAIrBFSSyVoktX3fAyGxWA+aAyoV1dTnsQopFYHpK2rxlTa4upXxHxG7llncQI
Jvv28963jBsYBzJ3Liy/Wm2EGSBwR5vB5OFEkP+o8Q2liRsWQOQR4f8cWKGhIf5R
+JQhfGLS/TinkTx8IGZd99rlwDnXXWMcF60ISW0k7ZMgrDdth9DedDVWZPao0p40
7XXjG5dpFvysk/XrUG6lJmHh5FpInKLdhr6zvl1rb/3voRkdYbHeUIfGXuniXe6Z
9iSbuXGVaPmphRpyY6O/vedNp/lV1V56ic9WjRqz2PYDxcljo+kGm8E8rKheN13q
fYuqvvjI42VUj195e9yVNPF2og1yr8TZ3L9z7fBnmurvJIeJUcFHq1pKUu0zB8FC
iImO3IAc6xGIoQi4HeXWGjySlzRKmTfaZbA7HOrLJTkWHG7OxD5gE8sMaGCqRteH
53pS+Ifto/F7Sppd3u+KfNCQuE4evCY2BqKwb6EAvm+zlNmCw/sjI0uWKe/WikNR
hXwnYMbpeV9FKJehv8DNPT9BRS4lhJbTma2b35X/8l2ztV5Mwvgo/MgoUvJZU0/R
VvuScErc7QCBNtBguw5w6U79lP7UpHBbwslm6Zn58fxm9uBuIzQbaS+rg3zJwbeQ
m+0TZdFMS3Ko1MW9Za0+/FmLkqxlEdD4FIROOJKg/Bp+i2kdGsEv9hPJeJ/ZiBYp
6QLPc2s6xhnHPj1DZDzeHE8eoHRD0cDyUBADYOMHd451WQ4NLyaj5/3rrteZfA83
v0MZBk/XqRVTkVyN2evSTBE03/hWe+fRZ0p23DNyELvrwPgsaDwSQbJwTDgMYqU9
tQEDXZXFT3qdQOtOZtbJ9SCRETOzVMLYCC7d4GpsmLKWMbGJl8sK23FFo/HZvzCT
pMJz3wYscBvGQAcqJKzhfJ5N0tB0pPpgqQszMaqe53tu+gCQjLXDVQ0N4bXF11h0
HS9RyOVH5OsPxh6LmC2RVty2JGVzX4Pv9BnmwXTgDPH9J3W7pj2Iec7CBn5+Bowq
5MPsXCAFAKoRIxWM7TEBTibN0d9i//8m9oj8TIfLDsPuDyDFHlmWf7nOCmebAhDi
G+lHXHIYompYwd5Au0+Yi7Qoa1uCsyV36rcUYdZWTUy+73ldr0u5GWttcrQOr+vp
z7RbZJ0GFgnLwd8ywz5fcG0JR0UGYEnaaVJbYXRq6kSnBWDzLROBWb5lH7Apv2jX
aRPmoL9eURpVeASWfVG+qG+bz+KclXjNqcyQLV0283Yg5Ii480Dn5vFe6MSt30E1
QOZidzis/aeLHFfqn0XPUNcH/VEJL+lX6C/7qm2HUe2PEiuIqLA78a/Eca+9/0Yk
qvNvdh23U6FJ/VOR3ei4YjUKw+0Ko9aWkql+m2aWFKlaPQF7rfCQH8RE11tKFzQ1
P4qozWsh2RHQ9DW/7dk8getghGvJy8rjNAK82WkMZVePam/rmHcShzd63Kf8PF7Q
moQQF18mSvEjDAe5sWo9pJcklQrevGXJ+hwacICPivuEYpRblpmuG+2QlOHgg5Fi
kuTx4Vl6DIXKToEpum3YS2s4Izw3xEMtHuduvo+AGDSrisRn+X+nfwEHAEHe8i9p
hLHeOmMiiy+ZI7+kXM56+khZptrcykyfCbMdr8jk8D9MYQ9EBxobOHqH91x++jS6
hNyuB+R7wVPvGXKFfcp1Cx+gqGlotqvV1W/Ai1c3H1+ZQHTYGUE29vnc8aAiF8e8
ks9+q02sJCvgAtea+7z81eTfl0I1oaYTUd7uOfqZouJ/K9SJFHGWFHwQU/S3pUJM
xQqR4zigKf8T+PqHAQdvqQihBvlBUte55CDuuar2VnkcgwQn6dOQEDs9Q8t9ACjm
0LMYIe1uh40qShJGXHhLsR/+vJEHy3Rj2RQZTkLHYVIRLAz77YTTNpob51b4fjUp
FOISXZI+3Pobb5nA+G89/WqR267UIjA3OtYQOnw6K/X/8Ndf4Vgr3B5iKZ1ZpEzA
WoaLIpxglW7VOVUOF7g9Ir9klpmW6vu1RNXbrj2fNMrtkFTA7NMX2wXEEF6wDtds
l5SBOmIX/Y4ay8z1iglkhHiNT4agPh6BFFvx4q4GNf2zH/FnaY8l3iDKQg7Dj+Lv
vmufInhfQlYIO9QQN1epYgi5MeKfdhLMTNOyxSdVuMv8jex99n1AnAHVnUqgM7hl
tjRpz1oXr3q6VEifYs4kKfC5sjxFgtoZrsbtoAU4hMN9ofiDgKLWWYbx/pCZXQot
hY/UhGDlRZgNP8w1Ws7ildUirmMDYbp5ASlCf3LrnxVLD9aEIxcl819KXjlXw14V
doAr0qM3Vfsbw5Hzn+ryWseglSaPbi14utqSqk7Ka3tVhDhqPCP4b9/yRdaLNX1S
kSGiVVaPwqZYK/vjVBAm7/gf6toC2eHCrUeBKvITMUqHTJmaQ9Q1dWVii4zVrkme
osm9MvxQHHMNlgyX5nK03Cv53gKsVNIrgEmIs1B/DZTR7vEEtUHPWfjiwCWEtfoq
5GC3Ie3S7SJ0nYoejymlZCuajXCXBkFWCl4FcfJTNi/aGfy/0k5fwoA8OohgQnP6
x5Dh1BIgQchwIvydeFIOlpiR/bfmxw3HS5pnmk28+8kl18lX2C/jd7UR6KC5m717
unj2Bb7GGO1nyP9p7hkkx8FHmpjHJG603NlR3JUUAn2XlK2qVCIKbljS70zISlAd
Mc8VPAHkvMcsQrFX7I2VsrHUJzihMrZGXIiHKJO075giQpF3HI6yMZgTTUrBMfr0
b/N0xf3vnm/Wi+XxQU+oP1zCfd8vbhwELmn/aiWOIb1A5Oe24kFJZwmpq94wlySK
1YhQXHfgjCttERcQHMhF+enIe/vQgEfHZwQZwZZPcm63GCkXtd+Zlm/cyqT1+3CE
WsA0XdYJupO18Fc6iz5xIysYXWvI/1c51phkDEKEDdPkcwP+2mk8cn6L00lgG6Mm
Dw3WKkOW0mQiyFkAtH5CZC6bO6TaI69jyhxV16+Tydyoe830oao8401cq2NjTUGV
XkLZEIOLXkmUqnEZNVCaLnDs8Nq5aVfr1p9G4guUMv1lWkVBtfmEwJuV6YqoAojc
4Fac2wyuNg0lLfUTI8UJzBp7rVGhPKo+n0uVMnchfUWZXBYH04IfdwuY+fVlbaga
5Eu05G8v0DCxk7wfA+rdxCcUpPLYccUdKTPArNWaCYFM09hcMsHyxZqshVEKYXlq
sFTUYNShDQ9SG5r86ZYCWsAyBJj3ARI6rl+UJB23Or4y9o5UHvFNMMWwkcWaLewW
tzRafv+jJy4sdA9qsggc2hDauWnx4dIlCqRRaoH9n5i6RHwLT2wrFbSxB6KaYizJ
v96yUROgiljxwACaRnp5JQk19eWN3P9qkb2QI1nAA6xG5QHPPp7iisBnYWPg9xJ7
qCgV9Sje/mkw0h+lCzlDD4KLNqG/O6OcEfFJLzVPMU8AiWl8I9roZdZOfbQkwMzL
QO7KFLsbh1RD+EZxlDt4mNN2tqjxu4cfHON5USmsLwd/iKeFDeXdvLp3nibPnjSh
s/bmgn2uZDJqOEOcrd5y1p2zwTv0T90ktwLUX+3iaGwWbyONlbwdrjyzaJzH0X8n
3zQ7AP7HWgvXKNZZVf0UBdOLT4HGG5AsQL9uw/4//Oh2lQpOTukeYCkoaLwIFciR
0wmP6r2Lel94wjPxUmlNNNTc44fA2pPkhZYlrLPFoX1leDfnHRgN4MTa7E0Yq++I
bPvCG4mHCvT/CiC6XBy6Oem26lfFZWduDKtNl88RRfOSsY3phTgGBD8nUrA4PhIi
g32nvK4fSA7lNGCzbPezNjkb2Wq+FoxvRxPGzBR16cPp/14psAY5W26zO9atmG/9
Ngymui6xkR33kiN/ciDBQsCgOdSDPioQeKnkpnuOUQvsTlR5w/qXjM/XhjWw174Q
ZrVYMKIKwp7ciXGv8lrxJj5O9R15t//XEDgvNZmzgVaanb5qqElBLHgWZ/IT/Dok
IpJMXcwMOwwvW1MV+TWQi1lqB3HmTYj26zE6NkGyrMQKxkdHOR3DNz+fTe0gblBA
vnER9a+kKrDzNOCIQPAOuCC8u08Io5TgtRZk6o5SuhoGkAc2fKyBlKv/cLNicZfZ
Gd8l7ecL7yL5jd+91xaBXo5JyDVI+T+CBHpq67ygEHvAjc1vbsZk9Mp9SQq2Ie6i
PKpEwb1PzZTk/8aRbm1jLpy4QuUa2c/1lmokfhNsjZ3X8Hhztli6kLhyatKTfXni
acliqV3hZ7p9MSfTNZ/8h22RttBeY3mdBq28ersol6SFTWQ+A3Ke7Jp3m1XO/+9M
jFE8OuCKpHvjAcZRanR62A/IWP5eeo7eoku3snp0OgD93FZ3sF8DoqALEOUFbrp4
qU3nODY4Qe2jNkh3hyJk9tPt3Rreb4j5BAjLUeTuHM8iUP+wmdTc8WKNqZN67SB7
nNCKZtR0ZgJy8x23MPoflWoZZtVde6FU2cP5cOGCAjsOiWi/ezGG20yhBAyu5n1W
mv75PCi0cdy5OtxzhYpcNjdRyI09VxIkoCsdkbj9vMO9i9nZU83uL7wApC2SB1as
WwD+gtTaPLjrdlQy0B/de+0CCSCcg+C4VKl6gfbEWXm+MvlCOTZEn9UuAMs1U9ol
5tkQl3p/Uccm2XaTss1M0pwBitObQkG32qg1BE/ciBh/lQlr1DYBBo72N3P5p0Ug
l/WSthxgetWWF3VMx5buAKnRvBZC0gfuYKLgETA3QaqKGTzjH4g7lTfl2nC7C/mQ
sslM8vhgmbElnQ3+ZvjHuPtwpf7Ehl5bBlmTUfJLEeagyfqMO5SzMepW/SzWCcEb
OOu7DVNWp0CkHaL6JT9R8mZ7E4nGegGyKv+LVN+uCJTy7VTo212h6vGcMJJrowF6
juUllksx2VOPyZMmj1JKw6gnf/W2cGI7UjkahHNZ/Gphp+V7ZvMwRAigTHXWW4X3
EIVlNhI/5Y6bLAucFXezHqbCoEeMUKHOoP5TJg/GC13+2t+ZnLu/aMBl4KsxEL2l
l9akzn8L3zq/gL9S7/PQcgvqUpS26X+3e7ct9ZHYMQFsxQsVFKsWvmnmQBvMfDaj
cIsVX1bTOoTImQ6JCZvKAFNofB/QTKU1hV5rTeLZqcU1JmIbM3XBuQHBhxZFWQIn
4jrgBalG67XQ0wXFtos7H73HBoRNVDEjr2+zof/JrkMLvOr/HcMZwx3+P3MKFq0L
kB7KprWi3bvYcz8qf5y780GYGQlgVm5PDy5/vp6sB8cRCUY8NBlgW0BGrDZ7NCvY
kRf4es7XFRysAmK+nXuaeHRNDmolTjHXRZPYn2k/Zezw8sXh594EbMAehMw/alAC
+AYCtR6hEN1M1Dzi1Puxza1GJWqbaLun2vhb1xmYJutme6agi9PkDjXJPISvPNHQ
E0qh6aMQVCir/pR2tZBPwcTSX7I+spyXBGkt8lfArS1e347/akDbdLnLsHTnNKRO
oWWrlyiPofCxniDvnNPZSvL+zCXUgs/Xz62wINt01okY3Rc7uIIQYsS3PD8ayijB
nMbm7fRHX4sR7Fh3wOguXnebnwPOvlkqnsI+uBLXPbo6AVyppgAxnemhGyNvQ2zA
4NGXsHNbef/0fLn8fjp00HNJvoDSByfAGbZB2qwXN/Wxjv9+FHI5lv0/qBVmSIf5
IxEk4WQToF0hAcz5j6iW4suv7EZau4e4bu1ajeSgvwhFR5hvTaluDmCepcRmoM12
Xiy2ZObqm9y6QlAJO5n/9Z36j09dp2it0waNiY9Ae0nmP1aczZPNg7oyVnwFMi9T
WwU8jPy60vmiIzXKDTZlG4dDTLtjbC7UR0oPC7KrhSr5r93SuHX9H8jJ4Gf5l3+F
fa9eSZZgZye2ijDRkOcK1O3T+YJyB3ggz00BeN51i8qs0VJkansjMf4gdnpEmWlJ
xs+nVeo9SPPKyty+/nGHYJvhA2Sj967SKo0ZGq5AvwhgB/Rrj3Q4qTmxLwJt2cV7
xv4/BxSb4BiPnJb1KgA0QIdq9fUypKMRoVN71wVKCHTX5+N08kti+zw96jUfmxzI
ia9Jo5jLDfaGkAg2WoIWPp5l/163g7IGWL+N1LDWr+rkSoVTRuhJBDPjmu1LMJyX
Jx9wenrxDkNBOe1Uy4RmmrjbuldBrl4+mY1nd3zHs+yRGiqOuH0y2AjNJz4LrKOI
KRkDsevNpeMqfWtbFxfOX8eD00VJhIc2GRqKc/4pTWEv/7IkCNOO8bROGpJ1gZud
1ck/Xea4dYSc3v6SR/nE2esg4o9wRqTQUgUZn45T2wJbhZ/nKTTjPsIg7lVxlvLJ
We/hs34hNfuwGkthB4zi5vcjlADg3RfXo8/6nZkTWfawhjPZnRwYy3jyGUlxeYJE
VbHce+ONRktXTMZ9tXtZ8XkkBEeyz2ZgscsQCU+42vEX9ULLinvr0jQRHxmuAy+Q
45nSgy67zJDHdACUYI1zk11H3706kgL3tMdB9KEJ0DQDzdwHQjS3MdJC4U7C57BF
/WADSQXpNfOkfSIdzi9i1vCcgMTwx/A1gwJC3AqRZEAs+jpobqHHODHErMisg4si
gZ0d5n65jk+jzSrGcughrBDTYQvxAx/ZjPLNICqiGZv63dNZ+UTt6AQCAoH80vYj
AvLHgI0YBy+yjs9gtW03tnthyscnP2HsOJSI8A7ZVHhd5ycQJAuP41tuUXWt2GFX
2pO0EW1vWBb7iJn8e6bPvrEnXxfKU8HhKySnuKkgxLcYz1+PRv1V3lZSSWRiR1de
DjUj/AK/NBXPC5CixWxgln+Hm5UvDUuJoH/9y695BWz7PrIsAdss1YrczaVeu8Be
LpQ5rtAZuCjkMXJWBaLIwPIFe2OGJTf0MStPUbczQrlv5LAMBvqqPQvbPt57pk/o
+AcaaRMSjKT7/SXTz3vKOdEQtzxfUocex+U5HQuelrlWgm6nJqX5aJeqZ6wUm34T
FMgd4f2ALuC8erJ2Wl1PidHzHCUY95HjeVUJUSKyv1UbPNKf4hSw9tu+fXkMX322
G6zvz4XCn3PRLXJQFJ/IDCOnzRrCqTIgwCgyPy6C/R/uyA5yTTSeauoZqoE83DBu
cwSq9Kloh/HoqNL4RMEyoA==
`pragma protect end_protected
