// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:31:43 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Mfuk5y6eRbHJS2pErrC+pMkbYhdi8tvIPA++L/8tRulRN6t1ObIpAA575cuK9rQL
H+kny9q1xcBy5j3Csc170ACdjPXlS70Wc9DMMXciDBwwyhar011ze+tOYJXopAQe
r8AuO1pjk9cIVISHK4GeBzSdjXw9NEjY3FdAv4heGxA=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 8336)
LBHqh/MW7tdfi93H7QWDMTBWCKkCqygdxPMi+vVirYZ9sChnwYtMc6cD8IUCIepZ
ml1yws4pid1ei4xTfRL9vGR6/HFgWKTAo3m1BUYUWAwqEPpWj/T6N/4Dnr6cbRLL
MqYdw+wgYFrqe/BzzfFQHnf+I3x9e+DIxPLSZrJI7M9oAarKm9tkp7+DlSd1MfD2
hWA3MUve3N1TGsIH3cLaAfExaE4NfB8V6n92Pa2a5EUVqiCEerWteHj84pFeJZYP
203Fk5K4rr9Q995VUU/5lxy9NbUHvZw/XkFmegCQxqBKBT9A3ZklqJxpNIAxl7Yb
zt0nodCb1fWctVLyECPrsBa3yHJibOon5NGas4wsymOVsdoxEN7Oibk+q0sKIdAd
cNG7rvpBsJuEbnOVkFSmRMPAd6mawIOJLyKw+KlFbYE6pMw8RxaOUSRSAP7mrkFO
A/c6L3+iHlNHrqw+2HcsPdNiGF4Z3H6rrcOToQfoOlUr2wWL962qESlK0mfsEYbr
B/+eILK1wpVmjclpi8NoJpUmE2R/9c570DwxsHYab9O583trSG3N+M/vHEtZCfHn
tog2cugS4m+a7eMmJG2lRvEzXlm63yFtwJL5CS/6GyWX0Dp/ID6KsxiyI8DDmLq2
ZQjBexk0V6F3oMOTqdnXWB8pekUrMwPEYZFQV/a/Ftdp+lir/H/G5koQ3z2ChE+E
NQrdnsz+WbMij8JRJh2HXhfcz9wWC+peCrpS7LlH5fCfMjzm/wv8iWtET5HEonkl
jph9U7E16hLQYS3T21CusWf2dl4vb7qWQ/755Tei3Aeeo1lChPavWT7U9KXtDoX2
yctyom1gmepzbH7Y883+eIBict30pu4ppJL+iW/idJ45uzCXPEx4O2ssghpP9WJ1
8MwB60YyQuGspYlLwDsk5tRe3deB7PFJRRtSvweW69mGnMou574gb28zTYjSFN0D
GgtELb2WKzz4kQz7DcT82eyoPZKd8D+CXTtKKHDd9FDyAzp+tUimVrg8cxYIQOZz
u4tUq/S9ZUwtilS49AZ0Gwu8X3RfjOEVlQdKAKaxhcxC6vGtwi3iKzHsNnGcdpJO
Fjg3oiTh8pbdcwulw1xX5gqzEcc5Q54ecraKSJr20LC+RYjpOWLe6Q7HBIRHDqRR
0GeRdMgbHETm/QT6RrQw5qlcPrAkjHkpSlLfrBreh55ECdtPjU4hlfPRUHSOfHOe
sVL8D4xe2MQM7NHR0Czz0Op0Km9CvB9BGXlWD1NcJRs+xHKb9rIa7ma4BVz7WJSl
ISQG33+xnGqxOYN4QqO2Wqclr9n8w8EwZv/gGjf4k2kzU9wS1IFy1DYtEaC7NwKG
13YcGjo3rqirmfVoeHR5cvlsrxj3FE8EU0A/EqkhjvxTEU/xbN1Ej0cF7WCp4th0
27dqq6zx3ziixhdyyxaFguk6Ekn1StWBSIR/kQRxlXWvsXOE1fm8CVsW6OOYUcms
ufnJ9SCreie8IRYvgVM2ymhEovRZkjh9O1bmAcaFpVZ73IY5yPtGl+ilYy7woAcU
hm/G0L+Cn/+a+5C4rXvbziQGwu1YBzE8kzmXbl2/NE+nMeH9hKmbO1+JWj+CtGkb
stcWCT/KyeyyQLokwc78Gko9gJbrBPaSbC683B9ZwQ6syJhcQVqjBruisK+8qtgu
bO6owGfuZxMxn1RLzBDJhT8EbfiveHdH5bekpWv4SU5sv8Q+9DpptSKLP/ZB4OLM
pfsFPgBWxx8mmI955ksEnUTrYPkhcsVaTAvd3STu/rHCSxcYGP22j0jXa9rOJkQ3
9XpK/ia6s2OSLu2Dfhla48lxZ28k2qRf3QBrY39RIUqH95lbv82TpSC0nx/UvbdH
Ktm7FoNlN/ngHFYNLc8H2jrCakTdA0xioSAoSFs5VpFrmDyh3jf33Yg4eil0qMhX
FtWDBQRm/V7+rX2oWFxAJr6M6G77lnMsldQWT78J7PDxPNOlUK/BD1Z0VO0LdIpP
OiNLnYxzRash+D4/el/8fD29lCOWRqKAtRZAiYhlfji7Bj1AETjYEH2gCggmvIYJ
i1wj/X6gMmNZ1XlXqk+ZxjazDe3lACEwyuYvICNVrVEZtAPEoPrRHRW/3NHExxJp
0aWAYHhJWTQ/JMJwWWeHdpJqjHs7VzUaNwxa0JnpbOQlly84V0TQ8zfB32ahg8Zs
YWYDxsc5XU32GKei+Hvzlxb/LCi5E8/fXaoA3LpdJ9orzPlIfNIdTB2yTYwU/am+
9gBV/jKv1Izoz1pTMBLx89Zw57//43LP6iXW3A++8LReNbMF0ga4rU2RzzVkSpV8
4mbHfAIEbbf0Y80s+oyafs/FvmY/hQZTn+JM4xc8HOHW26lMCkl2UlZkiXVdDGVc
x7/rqhZxaWSEyL2QY1+nE1IeDNDjj4yyU4DTjbcc97SpSyoWA//hIU/15pYkg3zC
O+IEXHUgbt/On17vdtsx4fKhmQqNCckYcxhJJiKChlWxLKIqAChcP05TWVLQkITK
7zSHW3ne64An1ZJBBypj1r1JxV8b9It+xKtBNPBMgD0MvTXk82qYGPVt6MTOKrIA
HBB0mjtUy8cqXg74YhZGxIZdftvRWzzp6WJQGofCXW9moI7apbCnayCOwtzz0Ms6
RzqXD3jU0KCmYpn8BqUlBd+1yNYa9GJdOzlj2R5+k10jbH2l6nVkmV889yWhNyY1
foQcDuhpVWj0YNvUOL90C1uWyh8TOfQ/6YCX2c4mW/tPD2ZPIQf5QILGA/2/hUrp
0uPrnBlqx9X2pGbGEXhZNniGjN+wmrFNwYwMeFi+7pJI1SN47J2V9IVflAZFU9Xc
Jo7026Zayi6LAEww60xJDdTvNtH3vrwcYXnW89wE1yZ5cPYzPota30xZlNgSNvvP
GeAeYG5LGWe1Srydd/ZL5gn5rrnqXgTg1bwcHgD5kxRBhcvSCJP9BDcvz+19NAJr
Pue0GLAXeYe+l8uJWERm4AhZi5zGp3ldU/N0/NVUw6IlRl78vzwKg30X1SR9ngTJ
r+Lt1vzN9mcEd0z6obxoKkt14rZnoffgRGLEzqHaOYvQ/iDB8IT1NEKV3bqbWGa8
9ffEnaWY7MXPqSoIazPzewF306oaotxKb91ZIeJY1civQP3jeWYZ3xelTGmZ8xX6
3CAaV2FHGO7gW4DSZ5ETUB+q7w+FzRDebBnan0wzJpgX3ZqRorZu0j+xGvOUQ5BI
/OHBH3+VWVmlqUPLRysTviHxXpv/VGpB9QRa6KBsNF6swyytPvOkGgQSCplx6YKy
0dVMoMTZW14NZUWq+18cQ5xdIN3giU1EwwKFVK4fww/xIoxU6jdKTmAV0T0jsIFL
Pc8K7OB1uAvRznGpHrQYowXm2OoXj00MlQ7tJrqxMJvk5SWRZPwM8cN7d/Otdvod
Ucsla9HmK36v+LKhf4voeS8gAIY06u1yy0eLLuGGq+OxZAlMuTq6Ay6kG38VBaAl
GjwHV900b5NJ7WnEXtZiok//8ARiGdwKz1aoRu7AmlfT5Y7k4T9m9brS8dXS7BMj
/B5pRHI00TsRoc4qSBAx15NV7NAUrkYGBbhY9044GrEax4wR+muM2f522b9sdRqC
CJbgj59x/5PyF5LRkdKZm2ToPDFzwak1ODLQMAL+hBU7/JBvtAXvGk8IJ3nt7ouH
bdrLtVQU0n08tZaQecoBprc/xLbLQuBL1VxLR13gTemqvtxZ4J8UihOs9fKqm3u9
BQl5WgKyIN4W0z8PjFnLhbZnw/pse6VFy4XcWhvM8Fi/sidnJ2KD1Uiu9wyRrwd0
i52xhT5+3YgvcFGHJfF1k+e9xbpvayXa1iFG6FORQ3yCJVVFP4025BMJDdJPp/ON
n0I0pDgyTE7YjBjoYlZEXAWFWUF56jzBVJyIkUrgdYaf0XX6heSJwYByKrqv9qBf
2OHTr2qvpQQWBYzB/HFVRh4fVtp/jLxMst+t1g9k0FAie2U+4deS8BXXxlR9rcwW
WXfPYQxN1HbCD+m9sv3Oul6CqGkHlht5rZGXEreN71qYGreKOwXXZCVvtET0CfnY
FX1YB09oMAKJ2t0Sx2duqd8xoxSe9r+/+ylv5P769IzPliQ3jU3Qa7MbJvusrCpi
l2kUK+c7Ua9aRsnpQm7YcLRb56ZygA8v3CUfIxw2rnmMLegvQQBUeQI6T4jHavzB
b91T3/ntJbsgMYZLnZk0Gu101TAikorsHrpT1y6iyRrC4meIFPDRbIU3R3aaVdb8
rxi5USB6WVrxrz7IxRynb/qBzskssbo5EIz63HYTptmJv7KB8Yawh5Xiom/gGXyx
r/Kc7MLIB2OcM/bGk180rQf96Ir3FBaodpCELbQv+vtEpR22ru2M6rs/vW3ZOFKU
AiZz0Hg1QYBrd8V9higjURWF1PhMLOtPAmcmzfQzpw1WgUqw3Wge4+A75Z255aOz
8UJluXGp0ASdLiPm/pXL5XZCXBjcklBIDvJIMXT++GdbNqAtoDJTQjsmTiOMj5Qq
i7YCDkINEzP8yhJfIZNfHgckJyYLs0YJ41FUOVVAPVvRylBFH75bT7kUueJ/xLN5
lsMpVxwCBYuViMoDssOynyZryDks9u13oOj0AoUabCSjQBEzkHfMtzbGMYzZ/69M
3q0kcXfGbdivhqhwjge7pXH26fx6zWORPLjq5blB7t4m/X66QUxeZJO8ScSpYQ4Z
ypGlKKLkzlOF0eB0NdKCUShKNFzPOgN4HC48peKdH6A6SHKQ3Ze3kX/fC8CT8p0b
F1PNfjr4ERLUDMwA+R6OgNMdVVCOlcQEiYz8R/SwIfdVqGFnbXrI5d5j/L82EIuE
FaHQ9NzHnuB4pCBDf1WoqB3fZNpZkgjyxf1P76OTMJvzr7M9A/Fdp0IdaH95jiRQ
hAou8nBiC7c+29QFXD3tYXIelaUPwmPxxneVvdqweMOS4CKlJcKO21Jgu0gLE1nx
ykazgeuX7KHiRuXZCKfxJeFFkRnJaKd8SrHCgHfS945guDI6b+o0kaIt1PD/N4iY
088SuJesfHC6xd0wrmi/hu5yWm5RE9eyC+LO8yl/fXUsjkl860rIgEd9CU4yXODV
lFYQ99RVTQ9dV5QCf8TO1GY7qVcb2K9dRZdEoAjcyi3tVJT+gCoErXL15F+A8QHr
bY/aGia4F3dBS7i+qGN+lzT9S1e7HO038nT8ltQlarNGhkDBzbviR/SXB9nIKl0Y
nSHRdZ0LSU414v3W8mHgR3lXKl+h68fK0VjjWrWnYBI9W/9gR1kP+JpuO3wI1fYj
vpHUGkIQ7FSNhi26PGoPgAwlyvBoW14Ry7Ms2H3INOv+rmixRxJzUDGcFyoRMmZz
W2TyipmeK+/RvWYcp7lNQ0SPE0/TUqawgPmORgNiUIdZDXjj3manNvFDDuuPVIZ4
ARxNz64C9KlTujCAWIKyYW1kbmRyJ9y1Sd3PbvKjOCPyP4vHj62/cNWD+5ytC5gU
r+GrF90p9Yq8xCgdg35bRPka4Ak6EBwP4iBCwDyrIkLZFsVkVPAylZffjtuHI9OK
Q9+DoceovBFNOf/BCerLLLy57J4Nwvyx9TqW8eRbSWXKGJPmXPjCA/qSRDueFS1m
cgMLN7JvUcs5n3P1UpoAcBgx3gOKBjYRJZt0zibvo9XlCaRdLsU3a0ut7vsCJcBu
2m/dVs4iayo/KLESEC6UuYmOrBv904OFE+sUCDjpm2mPLU4ghY2sahGVkG0vqro7
V/foEoQYNaOMJ5TIoj3JDzngNlNIs24X13rOb/MRG6yaRSYVgmnYcdwyS+1zMMYS
PnP8RyGDHBw1UkUYqqNyqNJK8mTsVJAHf+hHbNkQ90Ng6oMGzcvqiBY0a9tBP3p1
xpCWfURQIA3jUNnxuroIBe24QbQbFLwzc5DhBTdDUkY8cUjztc4LNbjfe07LTFga
usllCSaCnRh8CUrOHntfFt/2o9B4skxhB6XpWfKxyuNAS4wJEAYrcOSNwYTYbStI
fF2dI76La7xVrE0b2K8LCbYoFnB9kYCD4rqQWpZ+ug76azd+7mGcXeOvbtDTG2pD
7FJr6Ftrv8mmOHC012mlyFybNBT6RFy2EhPM+1+mRIynKvOYESOyocNE+p9Zzxc+
aI6TblBOeMY5n4Popx0cJ265lR0u7nEJjeqO1szO+ZCMCuzin3i/KyfqiQccORwG
ol19ewPjFqw9VREWrnsVPqTeEl1ki6x2+BkuXZKSLMuicA9HQ6VPvSvSo5VKi/tY
Y3a5A/IdNurYtgI66EDM0e7iZ0jMyAUJPfl2iov1x7lTshxKuoNJhwJNL17Tr8iW
8PlFPikIrxNLPPyIH0OqzCgWL0RoAFyIzKnFAJMTNXj6s/D/GpeCjLDeYB5SPhXM
6lzVoLqKEVnueHRdTt+Uw7f86C8Th81yII63ouXyUj2Ay9mRZKPOq2wU3hvw+n8/
o2orbyH5xkZBVQmrrkWYhM01U1zx9cUd9Q5oInYpaZggDpAo82xyDtX8IlGN8NVe
3439stuKiaAndAhsyEq5vkkLY9umjh/x9Zi+CqEFMQ1Ls45nDVauNtODsvxEbcZy
Uc4KGTw50laf81SaM/koD4/bUJA7OjqpLN6QOMEellAwspK2FHEohWu2IuFAERYQ
ruyiWFtdCB0MHkLX7z/9F7/lOTubcvhwzEsSHKEE3Qe5+r8mYq72rOYgZJyF0rhU
AILomTFc4W87FkO68cFydCvqqEoe9FUFMHjx+5xI67Cr+X5nHqPT24AtqbC6uLU4
zRrE6pwu2TJS+3ZPmBZ63sqoEfHrYGasz1TQmxVH96SdOkeTl5v8r6209sf6Lht6
YiWuzKho60zVtCNkS879tut2zRMDhz/89MKrac+qTkYD+McJpSLv584BwX/g2sHE
2tX2wbVEneXt+85+WR3rfwbAgo4+cT636LHsQu3+C5FEbPkvZzufxsWRJFabjjW9
23iftW9ac5SLK0vSRKksW109ozwqpEVwPa35Uy5ziV9jgafR0EUuqm0u0IrnYwQN
rSrnzWsE9nHu8f+NK52kcrqHDa3maU9+9gSBFl+gEvc3eVS/RksNQFNh9Skquou4
GKXS3R7b29khy9VpSihUEfC9lmYpPWr4pSJ9tEBraubCNrkE+bt7o+8iIuVoFb1v
08zzvRtFtersuqBgtgfMG1xdY/ZJPMLGJDjbUsoaW2JWH+C9mkpEW746LKjjzPTB
S2H9b/4Ntu+XlUFadhyoayExEqfFZMd3e+acRGpuEoUECNeBN0DLg9Xw1wnCsMpE
a0xmkINfhSSk6xKhNvUCPbn/3XxTF0K/M1BDO395ls6G7wJ/7somnh7QU7dOHica
J5K2Df0Vn+3F3rPIGszmaTtPz3j0wopyMat2viMpTfHjiP6c2rMXAqlUpMfqX0A8
uwPEdxVqf9iLqYYl+ZoshNZDQUBuoQd46XYXOzT1QN5klxAv5Jgl5RKE0YmpSUTh
oI6kkt+dT0LfDl2H+2f4xEOtecZj960rA41AkJ8n6MxnJWn5KMRlaK/EgXmddWgU
5jaw2SjhOuLrDDMNRmq73aY61F+ksz6eweeMrMBgi8O67GLXh3Lbngqj2TgS0D4f
k7ZH8ePfz62o+kg9IIzzDbIFBQmVGH8J1bu1rJwBJacA0b8BSIMENzYH2HPjhriC
enjmFyMSgA74PIef4W7OeDCe0WOG8uB3A+NwD4CKVkTUm61DbJz1ErgC+NKY833T
59EDAGYXFUq5p/HKWfipcFOPFZmYSJhjwd8HGN4JtE6GHjMh1ir98LiTSrAsd8Aa
lLe95rZWyng8+y3+tEXzRofNLWBS0VAb8N38NJ9ZjMqx2mRthnvx5IwIKYhiJHBu
TPltHWu9h/wb5qXD06onm4cS1er2E82ForKJR/gv2JhwMxDDLBLitlT1RiffGNCK
8b7mtLK6GW2DLitDir/n/tHjHcnU87p+/Uuzct31xbRbJ0XcduAV3dOe4c8oduig
Xs0giOiIr2XRxIiCbCPpbzzdNQi4U6lb7qMTBf6mN8uXClzdQ2okwAsmXFKV3Cr6
z5eIttFBUIdRLv1hGVd0YNi8qcsFpSIsgpY+2me4m757tunpRFFYm6ZEJyni0cL6
BNaepSc+3QxENpu4LTSq5QivLTPx2ur1o1TYYTSfpoKuh148xJ5yPjRweiTrMgfr
A9KusGaVtYSoh7VPLNGauJhFNm3Nu4wrCeuLKzFLDxsqWouezf9jsufW1H8OKvVt
IWrbeDDqtIkm2wHqg1zRNS7BK6QTIk3w/t69QgQ051fCmPXmKOIsmVnDmsvZtDwk
vH6fL2HrGDZkNp8WAnCc06/6WHaBjUVuATN3fezoKTBL+Ix5IF07hJj9KA+/6uLi
NmvkoqNzwPSUn2yVXODpINOa4QEXxlazAlQeZuKqJQwcugXwtDllvGNuw7heGn9u
nziKj7IQZX/Sl/KkJbknRL935R/nPRUp/GyBWcmDcN8HBvDtFrvEYS3jPpPXxhMC
GwZNY0a7zBDsVWZC+bHKohnMH5KHAtkNNPpKEXq4oBtYuWIBFo76m+dWVNzi+9Lf
zF+4czmoQWb95XdFSvTITT0ItNQOOdw1mJpj5jfeZUHNivr0aioRPMw9hQHS/97e
k5NB50jw18AeYCa/7WskSeR9OPOOTpt0SBBuqx8RSirECZLijGuSSNAczoTRvHqv
wgm7G/tMX3Sxl4YtCiWAeH1gIXAbLxq8eem1+fHN+Yr4w/6oC3SGgpa10KqY0Clw
QMfTwEd8pCR87ngRfl1xDFHcbsg88TPjpz1S3/a/OeFjws8duvegGQ3ooP3fxU6O
0sijlXpevA1xyUTn8vXHhAD40khkLHr5kNPO/EwC9vCPTy0SRiwhowSvNBIwWJdv
MMbl0QAQhx965LLcR6QkR4bBdkA8EHu/E/F0QQMdIQBelJJTHoiTjOhjoQBzz4Wt
c+xbaVo9KUAF5beRtvq6JLRimb3BTQiK3q8MhmIJh1V2pPPTGeTUvrHQ05o/ppXF
zayw7BZVMqmqD+IttRHPtyrLmT9luojzpWswTCZdNpxWNVk0MAbNMzJtgftSIbeI
dhKSijNTntaDQpPBc/AV4bD+TjkjOH+C9L9FCZ05l3sedaDoxyPepYxZFt4qAuCe
tty7DaZQbYEEggi6A0Pv187dYUt5S6Cxg4g731AG9HKAKdcHDIoAUdMlaL8EPn1D
s9dDALAuMJ9V0p0KgB8rIjWJrIZujL7Fz2HMBikLai8NeeD9K2s+QKu24gjJsx2H
lSRhVL2/STSxZqf5ggxeLxyv+xxfMcDqq8WfJuVbO8AiIUOdW4d0F9lwq4LvA0ms
cqtgtFq5ZB/UiqP4uO9O/zy/xPM0S3gaJd0eTK84WHX92NsE2XgHu3siEO43Bnyz
1xyqVPRwKuAgnTRTD72TpMch5WGyUr0Bc+bEwTG30IzjNcOPj2GpcKoDJTfXgUHw
8903bbEtCUxZUjohlE+vy9c1XRW+21LxyX6yDF++V9Lq5nPfvJMppDsExD1pSotg
bjG119sQ337Zr4f68HRy50QbVkXLZI+DZllwgUY0Yd2n8uFLpt9v9F4pY9yB38DR
2zMUWb3Rse50KSlES6ejXpOcNXgcSA/VcBVQ769T05rUHAxnJd8TfKEzoMU1f1Zr
+4s19keonAP9dskKnz77IQUiyZj2fs4/B5Y9LKuri5ZzVcJn+RMMN9JaICXEIose
s1iPZ05FKol2Y/CNYID5q3O5GYyTpdjdaOCfXFUQ28Uf4YWrEacX/+8TI/K3p+CX
yh8FNNAevnk4igeI96YQsG+C4f/1NeGNhnSKxSfLu3OBk48fkSbt9x1T1v2K+Gq/
RtwjaEgZKUK6SNX6VO9UKDhvA8dPa0rnQ0nEfj3Nn+qYg0NAYpRE+H4HI2sDUb8t
WyQRYZU4BNG8RsAAyFueo7541Udhww+i1p1UdLa++DYkq8U0vqcAo1gW3ZxT4bpo
VckQOcjV/9m2px9J3HrIYJp9iVrCv0M0WLoifBOFsQDdLUlpnQmjaTCYE+qZzLDy
iRPIPcv/N/BgSTFjvqVFLwRVoSrMCS7qWroyGkX7MYSNJjR/7Y8NLsXnDrIZ6acm
ULyioLYuF7XpBLhsIYRk9GAEOr526C9r1hTfhWWPb8eX3IG90ESy/qmYWJdyN9yo
xIwBU+spu2Uc1rek/iJtgNqn/vEg1kPWq0BTELDDnUc2+LvEiQzjpkPkZhVdKPBf
LTmHBGITFvWud56b/W5r5gcNiu7mpkEWzXVQvBY+l70t9mlO94xFh3Xoj/lpImc3
KqNnsDkryDwdTpXafxLFV8JQfwhYVQnD5qJDYGbSH6wfj14QhuEGOTLXCdiwhGjm
bLJdlXVXzO/4Ab4S+0iF32AwlG9HetnpXSjZB1X5ReQukA0Wj45sUG6WMTMIa+Dz
daZPSdmLvojFrIDRU+O4QpcG3xbkDmGXt3AjzYea+2T3qdV5ucXesdCCTbQ74yUj
Kk5fglMnuLK+g41Bu4inMvVvA3NG+1AMmbnhlvgGGRo0yrk93tCQQ7H9n8XHUC3V
tHRHZb6g5ArWBWLLbBZ10HsEEewlpqSSaakr2IK1MrUfuKNR9BpnR0i6q4/VgDYY
Iqor4pk7UaTsWb+c6TpSwimFZGpB6rAQ40m2LorTQdLvWEo3VHTBojSLDVwI9xDx
jsBCNZiokRfTNDrBQHp/naVvN3sjJd/c2FPl7QN+APaFiVLycdn5efFQVuVSMw6M
0GyN/pZgjDyang96uq9803Q4DT8UABzOu/+TJtW1ZssTLEnA830Hik53q6G00H5p
8B3FI8rxlDe42faQE1iQmEGU4NJQ0h4jMf3NpuVfCKQNAgF2ru44DO4A1cSmLHJq
ZnupvjuMXyExdCg7Q4n+LeJFtNIzLpfcVCuo6tf5aUpnx4JkpB0mlNZbAFYy/lRp
ll2ejkCJ0F4oUmjMr+jtiO+TzmDdQQdoHbUrTTAVC+IYCuXZp4vfwAeDSb6a497j
Z0G5AAVu2+jqyRmF0Xa3iExwrr6zqDEO+CwXTXXiWh/9oVv35oLkuwYaNZQs6djg
1aU5jiy8sxPkrkj//6UkNQ7pK/4ogL4k29ZH+AQl6Sv5Da471R4pkrbDEij30t4D
vSWVcPW4JC4THXtwe/5B9pmWnqfu3AC/CYi76XvcoPM=
`pragma protect end_protected
