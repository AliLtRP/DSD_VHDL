// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:58 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
slb0XYlXsG2/exfAkfNq9gu8O0vC9vatFDNBCxj/L7ShfyHYy5ZwXsOz7KdhDump
Q7PDTQbDA3aeQn7wDxwUwU2MWctZuwZDzzx+KzBc/FpEuzx5KtkERP00oWd057tb
TJHHdBOFqCD0BOoilNFLn2Vm2c+vtrnfRfnzM5I81Eo=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 25520)
MLXSeXYyQQkrAsLYKPYtmkf7t/A2+ZxmQBzWvqq6N08FU02LKSI3OWHdxGN4PX65
Qap1pYO+WYaIFU7dqM9vhabtBoPp6/SvHOUyry24ezX8R0+Gr6QGxIb+/WBByM6M
omwuX3Unocf2QNnZuri6zBqdVOe836eNU38L4FxCmWpdlsgaNTzpd0+66Jgz99iT
dGAZwAhE4KtVh1ogDpu9MW9Hwa8rmicaCspJ9iyuNPVT1o3p0BXG7sTIOYDeO0pu
1RZE2prFWVHJEbp9Fv214UGpsE/T+stL4VXhiyx0xhF/wjmklxpZ4Pa1QSLqSKWu
5UZP1PM+in7XkHrD/sjbvhXi4blnBLzm8NkKdTHQoxCka5JYuOA5W2V2ZXXmKHjP
0WIyGPs7WcJap6FcRSXdhpEMYBYTA4mv6Olb1B2tYX1iF8zxG6kY7BacPGhktNPO
sAAd3YtFMTWjpVNzQ+wJ9TCjMyXpkvD4GvKSYNfvGUByBn1qSlv60pkwb0WWysqk
U72j1qB1+9ifJn184SRoUq4+PrChpMDHI8WX+uhrVqRYOrwLjcqzMqUjMGpSF2AW
+jQssqedFX1SckfvDv+PbZxlB7NZEI+85dSNs5cd14LQ/VCXC1OkWs2aSjsdb4AL
D2G+CGsy+cJHjbmSzJEBEV6qM6kMH1saPRFBIAQC1z9p7g9B10kUsM0SiINuJDXo
D4LWk4Ii733qvY9J7HR7W0WSmTGqQxlHkVla5Mbdz+SH5QqBQamVLU9ZOJDweA5K
y8f/A2RrnS9SCBRS2vF1lnRTLbgbsOvbJeyGwQWNJm6g8iuOjmkdx+SrEfyrOfHJ
tIeQm911xOfcJr3MiZFj4IHu/rr8+fSM8Z3dQedHvBRUy4h5VrwYDB7WXlK84uSw
cYFQNiUe6GKnwO7RKt46jPjes2WpRjwqsSRx70jg9eroPLTBy59e5sAhZ53S3Ubd
6NyLL9DeBKcOH+/Lu30kXWS6CEapyP0BsG00RzZ06HF5lBFwslIxniezy54wKDo4
jBPugKL0VeLMgIg4stQTc1WiuQvuyM433fvG76mnMovUy6fXbFoYB6aNh8PEpHfH
YrGJFlfdILbc6CGBcPV6C2mScwqeDnOxem6cAAayVwqr4x9nWCs09LiFTe9F4UXv
TOs8r9Ev6m6nGBKq42Al8+MtC50DxFqgcpa6+MGIDwxSCtkeQthucJamKe3I2u6f
0IPvRRmPULiewNwuTHfuaA75XVBZikCVB5y1fIoUGaiuCphL8NArKMsgCxPWKP+O
FxuGU1JRekcKN8hHNkA2jt9z57S5E/IYXC3JsgvoriP5Qr8wJkiMBxURtIKiSVhS
B95JWN5z+yWME+H3T7KLMy8uKoa6Yldw1Gq8YLycdWuL+G8rcuZGhtEPHF3ZaLe5
cqo4vge5QKGuZEtSA++In5j5oW6vEWbA+QqoyeyBrEZDHLr5fTPJLtRbIDJVfr+j
zo5w61cHOdPHDKShNLjj3kGU4Vr4p6VsEk6ITSXHHGp4jB3lNwnO8WfIE2DDDHT3
XAjb/eYTe4J++a5LuI1KwXCWX85urGvh4Xi7O1ZJ7lIfAu4JTy3gRele1pZ9ngAd
TmZiHUDTlMO5oCP8CB4B+YJzGeiW1JWaBzU+5iLPyS41Lx2EVNjkixDohOTorE7Q
HthKXOUHi7Q60wq1TJFOogdZcOQgYEYQwyMzG7e0xOsSaGPW5gcjq9DbeATfv8AT
MoXp/w9NOsnIbZPspytkJw13g+q5xZfG+IK+h9TJhbinulNMcaFH+EpEhyMfTSEC
8JBpwEcjoYEQ0zVj2gxmxn775V1NWhU15w5g6KQeqqJAoSLEowEJ0J7mQ4hk+h62
rszJ4wNBRETHV2Sa1or3WLzLGTnm9sGZD8oaH9cnwV/H0OSpkUfJxfwhjEUv+Etq
beCb/1uca95cEW10kjcJg8KkvNQ0z0OWGZe4bY+pe9yg+jT5SQxNhPqKr4WaCCiu
on6dXR4LxU6Le8wC0UPk5Jq5tNgug6zN+hkU4OazMyZ1no6cvWTSuDOMV8QwQ7HY
/RZkCNq7mhusXQomB9mP8idgg93L1W15EHtsPTz0dVv2Ed2eA3hr1OyBjxWSSV/n
k1q7+5xUF2dWV8eWqknhLr/R4gBjZOvtgh8+tsWhfwwREpEpf49wxA9dD+g6P4av
aLWMspoqYApUyoD0SPTyA3Gd0hd37ZI2CsAiK1syAxkZYAyQfYvD+VwGIJAKywUB
puTV3xE7LQOdM2soJWVZekIJ9Pq5Vn+sPTlNVBr5h4xyG8BeU8JaZhhDmXIlhnaX
/f8hM04zyObIusGBfbnJdUSqK7LokxVjEYzhpRspQW9nFkv7aElpOSbGcuEkDPzV
S2tn2mI4NTjfxj9Anwe6CEc4lUm+VH4P9i3i8FnBHByTWNZ4WYNuozZ7OYcnERYh
w4mvEkDKNgmuXl+dda+TpTD7sYmMJFOl7KIx0H58745M2RxkHEiFen9+jMahUIlU
jZ11Q6lpsO9gPuowruBzEbZx8kvxa7XJ/6Gu6Rp9RwPBwnE21uy4TJ/DnTkZhx+R
fcikulSfe9/rLYL7JQ4QG83CGoA280yIfXJPYS1RUzfyFqp1uvZydPmQqWDx3cm6
LOYnEWfe372UC94crHvLRTI6JyAAwEHPDeLdrHXR6chdeHHk/lLLtTE3coWqVhjc
XADK+i0v54pR/FbBwGf9fkd3sfS2FBZneaSSc2K/ghqe0zD9qxveYEyipM0a3oc3
/b86aaeOdSi+yOUZvzi2Hn88ywIPZEqh72qfTIduXJY47nAL/6I1aJ2qFz1Guda6
lVWmyYFYIqdvi2J8hqd7tUcbexVrJGseeMI62yI+2CXdo0no/utWgBSiiAfa70hf
PGbmoR93WhL75NZ2ZFH3mgy3zQJxsiVyVgd0c3b/riNbBwf6jc/GtcFpnxZxTz8V
/s7XD2k1DOz8glBmcl7hiCHDAn0ynWT5tKRdTU3ffn3PSEG8H5zVGMo9SKe12YEn
yAH/2SlJ7Jv4LXGLpTkaz8VRn8ZGeq92HnC+0MpfjjJMkU7dGRRAlMX/EZvRgSv7
0o03CD4nKFMrZet0UGPIA0Yf4FnkKJcH+RArGQIbMXfUlhixbbnYRiBN6cxrcpuc
zmRZ7+y5doX4Wy3Pm85RzCjywj5EELtQzqc6+6AIX+lHsBAyRiAZZlyAd0XmjWqu
ASD/K02GLLlYnNaVt+9mztlVkZQwvTSN3mMt+4Jka+9Tjoia1cU80bzwxHXWTjTO
NUJzYjdeGxO0pzQcflLOkRt4T4NyhoXQgnISDtdvwdIYjcZCQfvW+oBIfKZO21H9
1PDfzzuDZUieBNm8+gQNHqZx5jr9rk0zz06GGa+J8gfhJa7/TVTW3WtCeDLeLrHO
xGX/iDRhPq7pWgIE65N4YKfwRwEe0Sz5M5FbHB8hquYmDxfu72Z1MjfXaKVvKMJ1
3qvevg0Dk+LityAO4Xc+jLMTsv+7xuecv4FwUKem707MHb3+5h5MRTgOdQS+xNZi
QFGkzypIB7QlAzbXHcWbb01f0mLlyM7cZFmFHSobrS051r4wLImutcCeEYJy6Shv
dKiDNmh/jEBhSSrWGPklIZZ3xMyMFJzABxuE4mlD0J6r1S3smB7oNFrTMF/8FmJF
HGGHKMCvv61im6bHe/Z184UBkQLZPJskgtm0UwOfUOeTpF77b/KhfFMKhtQxXxgB
Mr67812kh0cwURDtv/r95uZsByMBvZj/9K7Q92Z0U0TUZc7kNhh7pBfSFsUTBpXo
fIagvQWD/Wbpmb454WiTm3nbocYjJcEdkCSVdnHdu5+ukAhznLgevaC0BSacH+uB
mTWVzSKOZoBrYHeVqh9JFFVmvGXpET0ojW0jWkY/MyscnqjkSukeJOSOakIzB7B7
Ued5CyTfi41g/WBfv2WxZmM4pQtVcw9HkRezLhRS23K5zAU34anEQ3R4Yjm/2nru
Iq2wWtAlJME+1RW4NnK7106SOsG9qmi/Qs9Ws8k76yshj5sHiA97dxYDC981Iypk
ZIrpVxnOnr2uAkFbnT6gzDb2bK+nt4j9EO8M20c3IloOsesw/dAFMSuYxdQ74doo
gx2qtCAxQ4QPUmeWoHlaxmHrlJfiVZI+pc6Qj2DX28CgM/vyHMliNth05NFJT/8s
Tiaid94yTq8sYtAZvQmc342O2kuJpI5t6xobplrZsu86hK3pqajLjBaqOwCEh9tB
36FQauPnmH9+Yg4caAwn6kY2PiyalWxwX9d7TDSxRpyvZ5ptzPRnWxjR4Lxg2SGU
OeyoAetH+D3wLmd/f8eeH+YR9gUs68bzuwqHH+cq1wrGSEjEH1usq0mV0nHezvUd
YiQq71hTTE1VUlwH4X9eWQd0gdR9R8DsWVcDyznCkUjc8PGlXoIPy7DvCgA/135H
XA0NAOF1eqpds4bKuQtc/6Sx4dCFX2VEO4RAv6DdgWu83lue9xIlOIMkE9+2YpIV
PfyMrUHSjRJXhZeZlBtiLniTthEmyhGx+MDKgQyaiZIX6waEjuXtTL6n1z7ptmmY
scT4kn9TCgpdKUUejfTOpMGl0ZVtne3PvC3lqIsAvJ+t/Rrlzdu6mhiSxsBu4gph
IDIqd+UGU6bdcqGz73+10BYg4FOB5aH9leZl4WB6v1FWUrOXmx/YqqvRDW7SwW5l
jLYShB3/K9XIxOvI7AoahfOo+hHVDypEdHLomE+E34uBaimGrO4lTkV8TEgHaS4+
fSktJeaJMeU0qMj3x7mdwIl2PMzy3lzJ5ganM8ViWC4e+GjsYN9+9WkwMYYlkKlq
EQJIQliagTK5tRnek9RkWifEP7Mrx5C5hKjVWUGa61ySvryW4LKfAbleicSJ9aEL
df8d9VBZhQwhhBAFnYESeliKow9zlISas9hF6TNBoNJRRaFVeiW0ONcBquhWLrMH
M51rJA2EloZS2K57REjuVf8VKUlD6dZ3hPVKsKJpB5TZhgdhpLVUaQ42bmLvdX48
d3OaAxvogw8Otg7K0YAlfRgZp1ToE0CbvO1gRyLIPfA0ysNukhkOa5frGHT+dlLD
013QXt9T4VBYehsvYcQz4afNqvHpgB50x5C6ed2oMkjXZ3qKnjCIaKv8J0rw4wQk
ZtE9FqTsqQiMrcnaeXPdRVfpomClekr9emXN8RvfBDBD8ksLpMKCmt8MupJlm/5I
1cf3ZGbH+TO/aG15hwcPcnUd3ssh3R0Fi6kV8n7EJY11P9CQtTCbBFuupKJriDXd
LkwZKxiOL3tSKDT68CDuMhlEC4SANmqBgakmDQnKloMLrINAe3wuktBx92CWqXrf
hDX1MB/EpdI2bVgHP6Z0gIZLqPErKqNJ0KTg49oAikreTCo9TbEFTDPnYbbeF3J4
aC5FaUHOM5/MMOlHRJk4DPqlxxltb15XJBO+awvudSkmXoKMwfpKI5AluUwjEYA+
vBL597kHSHVUCpj2keS9AP7IzRRNAANYtGgQtOK2pwGzWiP+xGRPtJyp51+dhkVz
gvS1Gx3IrtxIkB6qNXv23U3ckDzEuUnNDIUfebMaXJIlm67su7VrOSPIjK4cDOWo
EnK4gIZE3hOAEf7xD6WjSkSU6ZbgQwbQ7VwoHP3fb5OR2m47A6qopeJHAkYfda5r
tmaypy5ZC2zxurVYRrkFpF9uLDqlfQ+18uwjVtpDvWEK5onIcm0sJ8+j4+C0hy1v
Cb6MdsSgXrIke6OSZDVqfwteKKrCQi+O9T0dWfXTVa9ZIX6oeiq8/EVxDBqQn10i
R2urnUxP+7UNI4xJm3G0+bnnmarWG4X9ResTmscpdfwIEovVe6CcbpGTQCSHgs3+
Z5N/NAr/SKJ0fehhPveBjnqq1cF3fOapaRzXBdpSS5suUkztRdtHui4O8c9DH+cU
J/L8bu1bjy/SIHvgyAd9xWgLXAsMc73Xs9Xxy1zBM8IkvDFhWdfKQXrpiHscTcA6
FtPNlWZGYQ1xxlNxyIgX7Yi3c/fguVUyq3SCbgjIusc+YmIb71txZAy85nohfARk
jX8pWkbo986ZiUtIWBxBRpCvy8pskIThBj/riwH8/PEoJPpixYF9RDkkYm70F8Ue
Up5fyEzRBOk1iV83iA1A90Zjxf3ypU/9F7Jvb3RlWwTFGgSlRWIPwyzu+3U9be5/
oYY11oXL3fO79oK6UVWzaoRR/BKdSjV6mLAv5F66eFUgbca3U/M5Sy+fulsi6H1k
NU182l/CC8dyWr0G5o3c+nEEcRDMh+3r662ytsDBP/4P+ybwHs96O+s5yi0ea1ON
9sR9l1Pn17IuyxAfnrCGK7HOlwW1gjUAHyrYywBAUwQDAWZ8tvKjRsMLRwJWpAtz
7s54DSJIsGvsVc77DvMUopQ2L7XZ/0c3DuEBjp5HgQ1QS3E8KeYxaCzz7p/hFJoJ
GZepI8VjlRmBQMBMv2aiGKRG+Mdo5qDky2hEr1xrwepzkOoYODmXEYJ/CND5DNIz
veTX17aVZ1QtKovT5Bp+Jlec5nDAtm57lgiTX5xvyEm4aCKClGkEp63IxobSV393
QZdlKqQ/VdT2Rp7GcTANwyhbaPXCpbkN5ZShYcCHVAdf7VGwcGgctlAi6tnxSUtj
Sas6IvnhDKeK1YEMg6MhwgswxW5yfpX6z1Ck59D8PTsKHRudJrdVOPTy7grzecXg
8EMJgCeGvIT2E07LRWqozJx2LgwJ3fK2AANypZRl833YglfuiTWwFav10KLRbm2s
IsUu4fJRCaV2u7pMBFPOjHl44XJLJ0VcLlOfewW4ojendl5T5Bb0woNs4A+W5/9Y
JUNTgtyoO+m6rzXIqLE/Kt+zUqhNRoTY1NWjBOE+hCghuXHroJMSWsjGxq1MGHl5
8uLCcatlS/Bba11jOvjYzEIqhgciHvu6kILuhzqLi7IEnwce3W7+1WRdPbms5Ds/
Ns6aKmL3wQimaXlOdL25Zx//yQImy+krxEZqw1UdnA8fPDHOCptoiPoxqiY3AToR
xGl8xCTYcjYITffeW9IFA0MeDPz+O6xhh39aT7PfDkbfenlfGza2VDmEITK/c14Q
HrFBaGyZmIhRzM+srTd/73oKSLerj9vRaEl0CUcTkEUDclUUl2xF0rzYTSunlDgk
/pr2FxcHTi528HOhu0TRIo2SCt11Nktd1rFPOXsaugKuc2wh4331G6W8YJkCxgKz
FF0+yzzk8DLWRYPZe18JdvRYLpLLR49OA1im3Q6VasSz1t+xWD6vtTbUAraxZuLT
EmIIUhdJKZXqrJ8fAyjB9nUShRfuZTLrYW84yPXnSdmXIsoAa9jCjlpA7RdXdnXs
KHAXViRHi2t0lA90e8HlDiwlnX+K1ZUWd7TdYN+HTDBrHEUwTFD270DBFq4D8ZEc
lBiF6XaEpQT+jVBPZ3JS1bByWvp+u+yNXfj8YGopBXGcK8HQn3tpzHKg3O3uvLny
KbkMS0xZgK89lDBPv9FjGRL8dJZRiiYejoasstygbEu+X8dRidEIYj53De8sSMZV
dpoDqTOrHobs5XNcln2tmwHDX6bXJmx1ishBUPccImcfXYVXZhc7eOLZ8hYBKZLJ
PHEm1+k0nAFMXGQSq1/7Qar0VSxd6UN2Q++VJ/9hhEzk6zh4PVG5z6o2QN+GE7HU
k+0V1iQN/nCXJcJYfXZ2Ygw7cpcuEFx+vdxiQHK51QlCqjMqdJW3dmXZVSV4NByE
iofzDCsAA/We+tgoJelqrOQBSwB0U1QGy7hVgIOWb8krPfRf2biI4PJWALLUmjTK
Mw/HseOprS1Wbi5EAoijN0/SjCQ8ugR5vwH/nTLEVBVHsbOsPbQgNzdnkTIb7A02
WUiI82gpxGvQ4rK0Y13c2JC3DSOdyZ6Q6O56JAY6msSIJonbmpi0QG8A5/z+eG/G
h0rpnuyxD/IlAgv4NvXwcXrHskr8CBYUa4LOxeK+JrPaA/9eDcs8BFZea6iBHW82
LsoTErQ6jJ8Lwi5tS8VNy1OhhysJ1TCCq0KV0V+6FGhpp0lfPJnZ6IH2NdyxQSFD
nbRWKO7PjtrlAAPmtArkScSKkmkwOb5SGGfUBZzgZA6bAVA5NLjVQqewoNDW9pnO
vIDOqa/g1s6lg6HWEEm7RQs23NAK7mQc8fOAqaf2FrDmEdNY0KXIGAbbBJ7BAv6R
tMp0U/7MxLkKZg8+RUeJ+cPSZ2Z64Ie0X/+wROFngGzan0RKxJaKV1VrsExZN+gz
b/4gIaG30KBKioLO3aJTOWvFz5wV1QNZrxYrK2R1AOv6+qrTGIefx2ex8vfBg8Fp
ngY9N9F21Oyz5sMexfiwcmnIs3rsCioC6z4Rvsmj356NEL9dNAQVr5Af7TXLkN4e
j3IL4EUhCPLBwM4rFZYswzNhT44hKlOwf3Pj4EbyQrcjTzTeoVHWjbTq5QLWwvsH
fRJpFwNG5sK+Wv4UArqZmioak/dGlk082CNUHF7LabG5QoisOmI1W20VBj5un30R
JcDWPRU0fhHaSJX/N/3aB19nucWrh7giT06ZvjZpy7eccCWMwvT7Wgdsn6zr7e59
ow2G0x4CqAT8Xlxm1RTjINhoYE2sd2GP8stKb7Q4QQ1PTE7zzUbYTIDSqZmCF7Gz
jnfNKVuKYbjR+2zV0NuCIxweGUjfw/N1bU64BNVgy6wwX/EcmkLf30B2jRncEEda
bZPSnJRB36qA6WfI8qNrLVUjIqer5PVxm+lnmCgQGGZ+IVQZXOhH89tkIWzNgl7d
J/yBkXSO6ywMc6xrbmdu1CWXQhObW5cQj6sI0kFmjDwNzsD0YkXxqzKKy19bJjib
hConC4ltnEYhhj6QTdVLlbY4sMWMjVRQQXL4rZGZKuGE0rQpEOANCSrQRpb/QybS
8wACwTZlAHLwvl+tj8ZneloDI64Tj9A0NjeygNEh19BSZmyJW9FVNP23kXOOD3aO
GW3ZAL5A6ozpm7Z5AKNwRDdSxD2CZ9D3utaalh6soogAqJon8T1lSOoTzzyZX7LF
i8f/D0sIDd4Z33M+4S6UbFh+P5NxnCMoSbM8f+c6yyUlW8axBqAgo2pMfUhGiUWt
kEPtEzswcZcY8iFFjOqfHbfedM6pEjGfTvfWpbqv9t901T+1Fd+Rok6qsKy53fxm
rX0sQ23Kc7Q8eJJ4mbq9raOYG8sYVDhVLDfaullMxj0PTQhvYonBEn6G7MnebNjC
IssNLJjtcv576HgLfaZI2dQuw1dYPi4PJ+f8xwxZRRZiUg6NCH3QP1PVlRQUcBjO
ZYETngS6Ef9xJGNZe2j+NnGxKO/Gx/IiGmMBx1lEwNKB6+JgZlFG7047oOBSB5XW
IC9teYUifQWK1MD8Id2dFW6j2ZIyB+lExbiJtMYL38NOCNdDf3Ccjy1vmEcoWvis
he+Db50h9/gBoKfsDOd/VhmaRJzqtcA8CLIdyPfdEd898Usg5GBaDwdRBBaY7Hjo
h3cTo3Arjj0iguZzFbxSNe6YwdpAURUXVxBTOomyPbFlKJ7Kn2KDMNg1RmaW887Q
QdTTrPmtQxUUBgqXmfO3Kw8muMj9dAbwHSkGdfAw/r0JE69SBh7jJ0su+PMNCQOj
aG+yJcuxXu+9JyTrXlsSjLUbBMCuFVVrJjnL9cHWrIhDzzAEUtoz+GXM8BMaBy/D
AwCd6NzgQXiqKltMW1D675CVbWB8owtSWMaWIeb7Z1mw0hJFq3HQaDuHHoCT/SJ3
jZD1bD2guDuhcnPYHydGJbqFnvaGaKbj8uXaKWm8JDb6XfBr9gxE+7m14CKsAhWN
9nFcY1hhHMhlmXmapcOXcITLKebqOS98M0uhn3xudI06XdQXqdvFJeYKzmwL3n/r
J5uK+7ctcSvpd66v+s5dF0bBlp568K6H39IKcofpZnxZG+VsE8PEq7z/g9ALaoYf
O4d/FGDEslgbl94dVoUlysHT+xz45XM+vqsz3al7KfpXMVbftPG+H+yLkGZDugCk
qbl4I3cd3nh/go01RLmk1Dall8w6MT8UnVX6gVEu9JA0l2poQtFuXRRZEIcb6RHX
QEOy8YNv2rVwa2DnVyjgx579UKfYAZUWwjs9cCxnMYRMpr0lsZ8Qz5dTD9p3r0vG
7nbrfWwWyU30iDVb13xnDE4BsmE9EH6oLhaZqQv+2P4GgFCk1CJV9C+QnB6byfRQ
7Udgpo32TzvrrIKtDFb1QH9E0e0rWYBbbkltrfNFG0fX2fo71dqhC9CWa9KU8QOq
RP6I2TMCJRo5AJMCF71Co1tdHv6qdDBGixIjRDHrDLxrDS3/LSTEjIWZpETzr2Fl
Y2tmHycoIM3x+7Q4ZDOf4r0myR7e+54JVBd2JJaosoPzgfgKTi/JL/NEm2d4xzFq
FsC9IWO7PfOBJM5MUg33M70d3iD/R6ZHxSf9OamP9S3+4jNyDhbDt3i15f9P5n59
0o3eLYtqxilz2zWKJCZ8ffwma1AV0HYy3cea0a6uIE5t5TMDBS3yyDkZ2GwcGDi1
wdM45nII3YC5WeXq0y88/D5G1BuYDYZo0leH9aQtSypy9QWSOvJmWa6uLQD9Wc51
gDBfl/aQjdvMUGjjqqy1NKadFAQnq9t+o5BEDMZKQOJn95Y+x43XsrNfppkK7RlF
gz1N9GWOFkdnxMKt/M1poxrs8xZF8G4YFRVYUhclID0bVCixl1oIEFT5Io0tprJc
h5vo//YBrxn5E//XW68hldXpcg68nicyi72MR0XVCDgIoYa6isor1DkzUGNQ8RpE
t+3CXwpa2TDuA1NqQbMSiKIj8RVLMj0l+juoEiBgYv4TWrjXQzrpWBDlXi0tr46Q
hpW5ibTfb5kDAPsyTQ//Ujw5wAnJ001b4hR6bvj+zFxHRrKxHeCZuNVX/24uNyGm
oUqujj7ky9mhs4z9lrqAXOjBXn6q8DeYd4guQsSUutcXWM98nYYF2VdkxbyHJFvG
dZFK3kkfzLNdnrqFIzkmLbv+B+UfJcfJbeZI4BF59GTUYxBRDJcLrP15Fw5SoPTq
NNvhpbtlLWigYnrvvNp6YsPVeVPKMUnWHNLEGXrzywZV/5pWnO5Uxqg7tHZhdL7O
N/uHTGq8rhTalr2InPCISNWFZfueyuLCSQIaI6qEaAC4gUkltc42FggL5tcLbL3y
wsnnwWO2m7zOzwEgTDlIbJqreLqxhusms5G8N8k8iD8spvd34qMM3bBGJflAzP6d
KHLK6AjlNxPKymAXxYvu7PJnRb80rInycs8afLKue+vN/UWCH57DkN0W8TXJK2k2
OVryYOHf6iENpstmp0F5ienrtAHPZsZhjCOnHi3S2oQ/De8ORr2tng2Fpp9EQdPK
UZZKwq5v4zK39oc+xPequAcP1pO37CkW4I3lSg63zv/lk4qaACjJXRvbRDnWEcuu
EVIEBdxANiQvRBpMnRt0PzqJXBrZ1KpH0EqJqHRhIsXrxxfJSAFNuS6SJ8/gbl2C
IOn2B2hLGzLgPfwQ7ASlHQ5RFYo9FU2AB6H1hk5QV3ZIoDLhONpWUkBqAMIhVVJU
NgC7mYsOcSKgRRtgsNd4Pqe1XjbHrbzPAplx7znxmgYxdgAfdO90TRXQ1nWzLCtY
Ja+W+oxVFrRCIZ0mnFhHOp/M12Y5WhKdZg6rfnMiTtg0JvSAZBzsYijRS2WMq02P
qusBi31lEZP89vWJBh/n3VIe7Zbf2aRU2/EZC+nGycYSwDotMrrn/PADEC66yaHe
3RBdcJPy1OeJvwbMTtIaeqJ7/9UhJmV4NLcEHCyt2tSv1uCKX7rL6OTTBNmghZLV
FKz8lg8PK2pDdNz6dL8motzE9VYO6An/ynOBhzwuY0L66XoPGfB6SI8SdDxXotaF
nyILHfhVxsEA4pMVT/o/PwEAc5Ss0YRAcYcKGxy/ySZ2rRSC24IgPqhkB8A1uAV2
4QUUK42PodVuD/3hoYgBQ8zykVrl9S4kBJbSsigb9A36TNMOmOdfmz9LTKQXpanC
JfCi7dVtcs/xjTFydi8TDwZLZRf1eNWb4G1GjGs1WUXOvdcrqkr0Ndor+sv7tXA1
BXd7h/OL90u0f3nDsRBZMnTUSxBY2TDmdMXUrIIma1J53PoDjPZ05ZebZSydrOoF
eN5rFaofKQGqBXYhQWp0/OWGq455IgRfxv1jY47fK/zWONczj6DL0Rt5gjGBW1mw
kcjMNBTtfmevk8PA+HMP2FL+fxXT6uE+YPnRegp5lkqUR10v5gguPX+TesydQWJK
Mj+THBr7HCotX00q8mNFuyzYg7M1LytOBBsAXHqoitVOvkz2mIU1zJPfWpw55A+D
l36cCCM6pD4lG3fanzuwiT3d4J0EPkBodeJmJ/viisxVxKIegaIuJP732Iae0VAB
Md9JiJRqO0NjvWYeuZ+XPZbXz5lRceiVodVyF5JAsTsd+rgjJi2xdFRYGfBK3nzR
rDmHfPGj8LlAOI6iaM+0mEF9ujiOfVC/sdeMehTPC+5noGnaa9hUR/acFH6zDdvb
937zHbwf38fk5B5MPNb6c2hjcGWHXqoDRoZxGtFIPSP3ZYKwU3mu5LIr3Dar95Db
tVBydOTKpQT9auaU4KkckUYJXO56QwaePYKiAcC9ObsJmy9uaCipeqQnrBniq3Om
lFS9vNS09e1uIQHugPF0vP3JVBYE+Qqd2oyjNv1YrqJfiGcfn/6WvwUdUzAv5MI2
rDL3rQhsfXB2ImkNZgLBh92JtHT1YK9EhkfB/Oeb5JXdLUhKYEnbz4iVAuWGZhcV
SJ54DQ6SM26sKjg1/nX6M8QifV1vZzAZaXkfDGJ+hSb+NXYvU71C6PyrqZ8xLnhD
wiqcaDDW/C4xAby5HPQrmiGGT8XCTlwx500EOxU2Kq0lmFziYpj7qTltcyFJJN7r
yyv1zTVmGJ8IwoFVJyVOIGMh3jfsRAkhfoNRwH+f25B/FeLJrVZDB2/1O8vjaWaT
HjOvwNFFTOt0Cda6czE+Uo+vrKb9Nos8CoMaGW/Qi4F/vQWxlQ71Y5fAAJ/MSdb6
c3aKY2cCK2VmfYTyYNqsNOzbQVFEqbm2roNhWlFX73I/im2JkAcWJHuR7z7pRnG1
5l+V6qYhPtBZCIxdswrIFs6txvbwDCPSXdvJ4U3F0W9Sagt2cQCwaaBCeYLHTabf
IQn1sbEyTZaRySpv0chMdJZbiQJe5j6coGqkzJau9tjgmJtt35aNh1/1cosslI97
e08ytmheLJRKPLMcM0GawXj7xqKcWDyB1YkoG1rtuortdQJ1qemc9Z8E92mUOqkI
9YFlVcj0arF2REBJsNY8PYbk/61LfjbJstu35sTXbe+PgljY1HoCsRF2eBY+ua1F
zoG/1B1uD2eWWBiFvQNOo0m4fqj66U7jvhLWZ0adN1ig+XPJN8laVdxJNjgSRAUX
CGf1L4jxqtY1xjywLia8fKBdlhWL70WTYYd6gfDm4DHSqfLrQx1HAcRbwPxn4kkL
bfkNh/TXnYUixyoxgWpfYoWqfY/NOpj5T9lBKSZ0Nw/e3Whw1PRSRLqejj6SrzJC
1u8o/ce8xzEJjEjZwxpzbCcqA4KHYl9Pwi4HWiOlQaTCeJ2kjBVrp1q3o+Lp1lS0
sgoN+B0kn/G490kwyUICeDTKmxhhJMrVsGvKCxM+IKPevD+9ItPRYxNTe0l3PFOZ
L319u5E4pEI8OgtieMRb4MxCzd+JaQ/gvzAs3WxVhyFLAbxMS39o9ZBYu16nZFWj
MKmJk4D8GiRP+9zRtkIoVtHwEv5TYsXIyGqAyNwmPHT+tJmSy+/D1aLRT/WrF1jK
hbNqXhwqCNlAyT4cOJTvy8gtL5t1hdLXdkXEOmbUElkfEHN50poOLLW8R7o2yIw8
REVc3GhX3bZp5mcr8GMIdnwoF8APf5eTpY3yQ9QAV/7KQvi3+I9djxSNoEZwKOtE
FhP6RzRZtgG24MMlTclsq+9mphbeZiUaayyKYPTHUfG90De5+z/vsSO1VIvK/1nr
+0f5MiopPSsWEiPuAxAPAhI3SMBZmFyoYmJ2ZaI9CLoHhuHn8ZHP8xi+/aTtGXhy
q2oJsZ/OHKfMdBs8l2RSJ0GSOcJw0bLGe0xB9c83JzGN1RmD4xzLBFM8nuIqOmxa
xTyvQu8uOHInvQ+nC4xF+UTeh/+fLiZc6keDuOBRjuAiRBGFwYJWONRJIQYsMXhs
kA27j3Dwvlmv9Kez8rck0MqP/3XZEpI0qFhooXuwKLnVgmnjrfGgOI6XaISHvQyz
UboRx1IZKrOL/06whSHQIX2J0OHt3AXwZNXBWCVZ8P2ifiEwKpv5hUKW18oTpcNC
okyS6wMtQ1iqqLjjw+/LnuMumzgLF3iiuKfnQ/8H9GxF/Qg/pBAVomLpN9JC4yZz
HeZaFKLrUjMGTI83L0uAM02ra8iY0gkGOW+ExphZLKARODP29U4vp1q+/PbMC+wR
HOOrCyJE46V5bZiX9tYbeYscv2ExiJYcqIVur9DZRO0kylDK4RBfRdB1aWRDcef8
vSHn9WnZMokjHZ43oryhSSkvuFnPikVVj8vbqw4kGO8IJ8f7cu2NoarWuYkrfb+1
oRIib4QdrZSKaROT74Jm0PxoqDZrGQhAkNccCd5vBkUjPOHxP22WTHAlqOonGeAw
9ff3aW5rNT9boubEJTVLiYnSUAllegGEVd4DATd+bDNVWA4DP6iaXctXTdBcqNn+
KDD/4ypU+cXl0ylXNoHf+bzbsM284ulAfE4SxmwMfKRLpChZ+VW+p1LLZVdWIJpy
3BWiy7CG9wN83QOneBe4FMqR0PxmubYfFauqs3/9C8LQsdCvA1IiqKxU9rET1jir
lD3YDPHaIjXvqbYD6nVNpKjm9RCNeQ5ByiNzXZQhnUdiN2P+ujHXwgz5ap3eO3sd
hIC+vOxwBrVvEiwH0qVDar+eV3tln3J78xfPEA8Xeryw8TtnkNY/GvcTffT2R/CM
ZfF5nfn+6UWxwxfWGorxCx/GH81X0ucMkuxtSeBGpq3/tRotPEs/3opkF97Sr5oZ
6cu58j2A4Vybqi97WJJQWnPsNE9xHYEYP4y7XIDTxPLrySUgLF7hAv/sEb1p9/7W
RB3W4yCot43XoOoBqXmKP1YvNGwTIqDaH38JBHDpztP+xK6/tD0pNUUqmkjRDa9e
aUhENkCymYuJC4UDFrOR9nlRCMaeJVhgPET5fa6arn24t8OzE+dFz7FmsX6RbTWa
dTiNRYbwZySetAOpX4EkZpxz27yPjkfQHZRUYdqu6qjMYvXSCDTXP0E2JN0l6pWZ
XPGvC+1Vp4xfVsA1XB/5kvBuh5/tmNQvlCwTBN1kk4k2p2u0KIeAuQJuE0+Z6mli
mcbn/4+efJTaaxdH2A5SGH72N/Y0HCvfAw1v5JGcC82TXwImF1RmPN9DZh2oNj7Z
ou+qFC4MQPYImbREmUZ1/v7IiTaVLg1Lp01lg4wVdkLtw/JWxnMfGWYVCvEqbjmJ
+Wq2inSQsQXmcU9w5hC5vdGly5Au6wRnqS81rzhjYdvx0jSpWktNgIQ68IhLM8Nh
5negOUirFgcqpY9KP/nt9PYOy1muJ1VastJYtKFaQBqxapitqqTAPAFoDeHcd0/4
bNWZKAK7cfnXhqEJV+3AoEPYgHegelG8OSXj2+eGelegK6OL4jH3Dzrt6mDJnVGm
jFXKLR9OIP6jWVQxDzIzWroBGiDL/ij0ztu8COt5gYag5mzXnRILZaTRzvD4kUTc
3rCVT1p307ZiwYPDQiRJ/ITNQoL/RU6mGCACChjWpwyz2zDq47iMgHtTli08Wxl/
lu/0JzdYn58R1MHoG771ZMSR2U+pd+aBaznRHVlcajWrBKNI5zmvyGocMC9a37yW
MaxWbKBnZKv7q0MFmRxan/6ZMFzykL0eagt3QknMPpn+4/Jv7NMJ0M+mhETyLGQA
lTKENydzT3/UJ6nutXCqvwubTAj0XAVf7NMP13hW1hhUoZ+XMcjiNeZk6c/vk1vi
vSp4qy8xsyUQ8+SMJJz2rERx/+Q9+8RnuS9VCztJhSjHLFQwK4SNXh41cWU94phE
SJxuVGO/0A3WLZYjIk7kKEzZbDJVty+FvdV6y7bf9BiWXdPlIDuzGMxJWbz90Uu4
wGfyZe5U5ws4ZowC0CWf89WAyS7vLMk7mUERnz5pEE5WCVpfefG9n9hp5432yjzW
NMAiWaqJMvqfZEk9HS+C2dsqDLKHEBRvn+k7kqVtFM4v0Emtgb9vYDVWi9GVsDga
1hQN9Vf7axq0oYq2S2VUG7gHdQUoFhVIsCWWvOq8lCJw0tnRMVCGde1yvLWgoxhA
gQm65QoaEZHOKvFw2RcS6aFtOAvtg3itYXPi1Z9GCLoGbnegKM8VWmoA5qbdf8cC
8qXMB6mX2ZSUrZ9VUNiwbl3pOzvZmot3fQPF2MK7JUo90j4fGJ03GDXPLU3LKt92
9dkHpg2ZS345VATlkX/GQgeSm0nU0wz4BzQ8yO2lqjl/+rOtqExs/b+igTpNC2qb
ppjiqJK+SMFncu1HV4pkMfZD6rdhM4arZaiV98DJuD3ERpHanPzSq6TtiyxM0acP
MPsb1M6IX46y1BANUh0ka0EDxmg2x+Sq2ERMjZYY+gy6KnQBLL3sWmacXftAnESl
GdH9FeHmPCTVCO8TF4BaX63gG9j5LWeUrGrvZetrWElcN6c0EMmP9EdVWNrbXutF
68qcmeMbMHe9G/MAsKkY7KyvCC4pDCT2qzUXJCN1y4HNh0T5U3H8dwrWVH8OLP8S
QjeRKeq3rBktYYe/CXY47VtOecXYFSP8/tMzhXQa4wHIWtpgO+fCc5yj536BMDWU
oWTOOpwA2gegMhDXg7W/j7M+qo8avxEnK5ix0tX5OE5FyowpSkTLWtqbucZ7oDtL
Rxg2kJafMqhSFXUQkHqfxoy0GCiUzm82mZrS4O0la7g4tv8QGcVklZLmRiip8SHu
IpmoEadpHk54pE3JhEExXNrl/PkHU0qok555SpwY6jkQC6dIJ+aqS+7w6yWHvbmk
nvLo1oBCBGOvA4LJOGiTDcmv3taldtsq31PV3wRgudf5RgoNbj3FdrM+onjzwl7z
sbaxw3al3fX/1jjCCQedjU1NI8EqUSk8Q7e893zZKDzmJVkWibJAoKs0pD8M+Ciy
O9mYOxoCcq+8xsKgf+wqlwtCamOi/At1u3DhI+jjN0Hcs6sKHl9CweT0fYhSNoj6
rC5kvVU7C3PzVZLLH0X0ndJNiSxdux25c4PN2O9e2G1rpHdCcMw4cHyzYfS3hCaS
ZXCz0c7Tv9ifNSLJ3uOTjMsEPpuDNDPjZ8aQF1iw5fITLOT9TUes/ui7PeO+uEvI
uZzBs7SLSX1D3Oi92IYlViPeRJlxjViZYihtqXn/+O682kiX+1433zo0jB0tXgJ2
cnFUF4PP6iZxfHLOHr+t5B3gKtNewHwlJw6g5FYKILfCeEy0E1aTeJe/sJdYVB9P
Pj2uOpQWCWl7xM+Is5W9neD4wMiX4AVg+v9tOtZsed7tVsZjOSMv/cvnuUVnmQUw
LWWxjkbv6ImjgiwGCuQHzcYfWwOKJWhmhbIpas8p18EUM1NUiVyrw+KQcxxaOEFG
bUAryKA4EnhWspxv+qxx6yJ82GjZivPKMt4uBdk7PGmzvosfldY8dgIf+pcHJ9rW
aTTh0QS393buQadl+0lZXi59VeajC4iqcaRSJ2lWfUaLfTD5BcNysuz1e/trSB41
PgQCUvmJAlUEW1ZtG451D/+lcxbXQCxsIuN10zBLW/u9bBNukwCC3pS1F04wcPoq
0u1TNRARU/3Ne/F96P3XKvDkfmlr0anY2AVhqiAe0NADtjYvppdPVlzRcrr9OkQw
66ZsrK5lHA906PjIumsvEM80C0/lv3ZxeZ5ofMZPEeGtX5iooHWjgXeWF1mDZ36u
4fWb/yw5l2ekS1fzgOgcOwjISb7sWnAfs+s/Efa89j9hWhaE+UE2kH7ct/qoE4hE
c8VptByitOgaemWqi2GlNlDkCHw+QiIBI6GK6IWfrJ3upWnRtV3jIKY2HGyB0NXg
R3DPkXpF3HrypDmaXjpOVdk4E621GD664qC0as/x7X7pRbLLVzv/bCiRTV0Gq3IT
8HTb3H0UXFH7phEmPS7ahTEnc2SuJAG28fGVirSDxhXVjbxa7PwETvPD0+OCl6JH
i2+kMRjFR+XWbR6yBm6B8dbEf+Y7lglhB/jYo8BGUGG4FIMPaoyRt5csD42gym1f
E9Y7kW3ZrQecjqwl9ACk1OLCuZNG8vOx2Thgcl2wGkFRCkvDYDnlm1Ytf2y0VoJs
8w1Qt/3WFZDZmE7H8IvAIMvgBDQRYPi1CU8DtmeaWhfjRhIDVERrfgvv+CrDwbTQ
cOdiNeQWKXrlVNDSFTouymp6N6ZHvgPbHSI+A8/tO/zgbDgWCfNiKzS3Kp7fc/pa
uGX/Us1dsCNIxLcofyMh71puDrUoma/faXM7pLnhQbUusl/cx9GF2UJzNOEqBBYm
SbcFhTiAw1B+LsdgvYAxS6UyXe5iXHfSc9Z6umN5ZlTd/pcs8n0+9EZMLr9ggccH
Zqw1AUEwnYOD85YPc9oeUQkJA3G7yE6/uckUqgiHGDsnz8OnN5Mjryu3U24YfPa3
I0ozLPqysQbRSAP0nIADOieLedSAhIHWGHpJfjGnDwvbtaEwwwNrIy+KM9DdQyGA
utePKHY9yrWQYyD6PjExy/QVfwRiCD2vWaxwV83hjqnORz7NkaLpTNb5R8CsV1bO
zum8pg+wF1A1PP6RGFSRB74LWYDpkNBUiIPEDBJrhw4TMaGrt+0/G1AY8CawDQd8
86FbmeT6BEHX/YnzLabo89goFwCB4zVLlW98NMi70c/En1fNPy2W8/vblNcPS4Vq
WlLUud9WNGTrv+mbD4Y2QhOKPKzDEPV6jRy0Fa6Zb3/QhMxcIfz5dFikW46kGdIA
BDwbn3rCzkZT+VuOuMxRlTS69np9/FsObfpm7V6E+30EP4RSETbJrM4hKkbjU2X5
8s4l1iK43/bAy3Ij1wxLAfB5WtXnlL3CUC34piElc2Bnfuviez1y2tVtzkB0Z9n6
2JyApvnHkeX4a/2pB/CnrlwNxWOdBWZ4K74VqsE/sXQQLg36pJlex9JHQPVx7iCM
5QBPdevCc5a63PBuqs76Ymslk4vkKRoTUqpyZrubgRBg91zNaqLiZp8vtvEPvi9p
b1ktlfWhRekeX64ozjo60r8FxTbLcuQNe7qPObdaSYCV/aIZu+Rq4bIdwA0eYHF8
vQ9qCOld3HMtmSCZzKLpR9nTn7Q/gEfX6pBntC6Y1h3lFcfn3AZxgVh1koSRnyyv
Yn5H2I1VevDC+QZv86gQmOPRqcGbAqHd/2ItNEYtOvjIRvkOMXhQzOQpxghtx1ea
7pk/vL5OLXnEOHt8nMFemBa4/SuFHMcs+0vlk98kQh8h0lbdudvuwPKuh72HYbu0
k1PgqamxTBOx9/cvDpkWnLwpxRa5gpCrmrAIs9i3NH9u7EHhejsqNOqkXh3kJP7m
FozfcG7qETCaHxdL9pmPD8IN+h0STuN/1BDdNeNNoPGcaZsngUkkkdFX/HI7ibFs
xf/sUGUH8lriFZVQx2pPar/DYMGUMARdfYQmz6dW8zMFUONVIbT5u0vncWr/C4AM
ja0vq9nrjkZ6AP4+JXO8hhl6L389TDF4pxgInTV+lF92uZYSHaibX0lfNuDEzVIO
znMysggGASmyMaFO2x5jywpO3V6cmkoBruwiYGwK/7eUmxWzRpH/1qakk7nR0y7P
istrKYlENMGyCrnORkZIIPHTByFJtjSfsl+HsWEuq0Hwwii3Tn16B5z3LMnyWDtu
EB6v82cuzj+edRxsvJHajovTFfV9uflVa80NgUky+pwsiIdeLQOS5j14NoI8wjcy
/zxRS3gnG3vz0S9ITrD3S+3SgrybME6W3G8aTcYfKLYJkM6kiJssZQN7RKzNA0Mg
81RhhOSY+ktOmun9xejlj6lP7OBDADwU4EcxKQUeHY1AYM6qpMrD1E+fucYycXsn
OfmzvQUjsn6TDGdv3MMGCcovm8Q9uSXnJMbHi6YhCx7d0zzSaeJgO/rZ5DxSADHn
xmJE61u7aNBKEte+gAmrPq/FflYTFUBEciblilQQZKRQeumxHTil3CxDer3N73q7
5CswUAhqHIUCQXFXqPi7Nyn3U/jwUd259wr68i/d9OsYSIK277KQtjFo+o3koFDP
zuwjTavd2nrvT+NazVJmWDuXyJ8MCOlRGOm4RTJ4S1GrK+FqRrzlWSlwBQg8Vkn0
crdilXSpsHvEOtK+/BQw0KioHwYXzO1ACvSY7WUuP//E4Yzy1tF0YHpzJm2GbNi0
8kw6OG2n9PpO8SN+e0K/WOpK84fSZBkihAlR4xHHaQPAOnRunODsEuqL/nvF8Lya
6MBmeQLnTjBBX6TgM9/i0B1FBuX5/JAygi74hS/2MgDqvXa1BpepuGK4rmSiIuNQ
AmnIluN+8MiBylZnkm6PCVHh4EtB9XsI7xfjXmKIRpLmM+D4oJbwdFKaRv/jv3us
SDLa4SvCuZNmjBR4zHVHGAGmA00bGMqqrySrqfHEh6UVVM0MGvkTndlhPJgRdFx6
AQPVlDf/pHA8TUBYpTT81TBUQt+n5pLIcSgoaO9DbikDjwtRbnFcYvViMOk50ruz
JE1GXIgLvOQBG8Y8msB/RKBB0metsAGooHgY3JgGgW6KvNaEPjjJwy1vCKOm+qKL
gbwKFdjbhEHWP6eZx/xEAernvJrwB9XhRPHyWr+7n+vAB09qRrUESB53pOATdHow
+zXzxWp5OxlOEYJNaOpiamtfk4ry33+yuWXHeQYhOPum3h1IIuwNXqG7pWYfYe7v
VsC/K6KmyOkSrOeRmpAhwaiTCEn2RZzevZwh76pfQZ5XrbkaKnWR4TmTu57NXheI
r7c1X4rbRhxGEZCmFwPdIQUEhiwnO1had3MBtw0ubE5hVco7pEleZr3raQwyejJA
J1IoQ2aqsVBcRfOQdsUb/7voleDbxxZFfIJg4GdA7rOQmvLrRbdQf/irQQ/sWyIs
sBouiMEzrCfUDHw3yPPzFKc+jsOlvCc7rXJo2U8xd8vvT508hsqEkCuWjckLKWMy
FTIXkTmgLyZZ3fLOtn0Exqh1PFsHDPR39KPmmX/4AMXGhlMzZimjF/6kxe7Ta+Y/
KUXbstTXadJ6E7zmVhjrltzz0KLX+TaxKein15cCke+nH+PK5ZaJPojHCYq6mJuU
fK0KRI/7/pAKAprnBX2juwpAS5b736ERGL41GzcHO8tiFX+V7C1hSxGUyIy2oFgf
/L3iGRvkbUOJ8kfnJHUFeJsOmuASzpIjulwo1AuSRXnAJAe5xg2aksV29Pgo4zTV
vahSpJYt8R9rXJuNvJ4l4fYcdHsw9QewsssnFexYhjMJ8reic/n+TlnQqWM/75Bb
/XbIT9P7NGmS6Ca66fvXT1AD5WULW9ibRnRyXDvqJZAae31MfNocnxNN6r3EhvKi
79eHKPiQVUen8IYpHMugjUV7T+icq88VfQKI/d713pAwJB7DXMjglpi9ssJJf4EN
SL+C9/NEU8oRwTC/xktkBBdU8+NxeguPWC96cwoYEWDkaMzB0AOAuAFsEvDcJXLP
rmm8DjqP0S2CgPfAUUl9BIMwhar96c5jSHkvpi+YSYqhPQySbiv+UNZjakjoneYF
q+/QrZAGuzy7cogeu4Th+7qXUkwAs+kp4Rr62oGF+HPPK0FoIinFm3qWL0H7s6xu
t0PBIGL4WZKSoeX/mgXRtEH5uz9DDF+7kj+/kF6mqkIqGIB6fMgSGIxyVs4uCq0I
h9JUr5DQm3LEwGJVwHfKmyfZp52hzpeLWslOXe3vDsyZEgqO9av/x1mQ3LveBKAE
znbjTFwCG68q5PiSLxBpGsislQQsl4b5rYaikZAH4wZImf6sNjaXw2OHg/j21sOJ
F+5zvJFmnNxzq+qkFWBMctYfm5MHnQmmMXRXRhMMU6pwIbLGX0SW780J/AJdRp5o
XewZop87BrgKQZpHdfNL5REecbzIa6ETO7Zqqn6HZ1hrAefv1VFmXX+5ZNnQfhXo
OuHwVdTI05fJKgBY4Vd7p7QbVYWiFvPEm5Ctz9Skae51tM7/cObIcjKPXEF+NGOl
SxUNqkOuSSVERGQ9gzyeohQXOjui9+5pwJgivGWOE/6rDPcp660KVg95EMOw1DzO
fhJXL5U4NA70gYRsSYA5ymobipATLEEiRVe4o9IxHbbsfYRaN3KGGMJooFwHQgfD
VWL93RguynswkFbm40M8qhG1hHKbB3UevK5ByvSDYwDyweGJDCF2HyoAd1zPkwjs
QkZm7ZbWGnHHipZBqNclSvzRl9VbQDDrsynuxbVaEGigLuoeu0eH6FMYyU21QsF3
/GUloAyA7u56umG+XXii5GwoV0UxXvI5a9yWZiSnE2eL8xm8k5hNNiezxlxgTn9Q
eY5snxn/3RrEROnkLggw54YixrZbJ7JqjsIlinCdCv9Pr9N3pHUIDxLiLcm8i9RA
DpO7WTJDMrGD+H7OBPhEvvPKPFnwlUwnCTkV0He5TlPfIMOmp5WrhpJ00r2OqDuu
nrY6XCf3z2tmNoHVShiJ1R0pyIIctloOJaSU4ThJ4soT8JW4qQFXzOk4WFA0Tf5C
iVTziOr0+8HH6kU/CITkorL07oFYYx4v3m/vCmudhIvWawhE1oWravdB0lbnKS8n
1g6SbUvKTnjFNNc8wJEGacJf/Q+kpWsnBXZ1dziWIDMO8nwAlCsBO2OQnmFGn39z
XmhLDcpoH1lT8tXWSyI1hvSVLje4WxVX4zlbRMwuX34Tx+o2/thv78UIeb+wxwNR
CnG0NEF+N3zkO9IppzbX4Pv/SYljkpZL1crzKgT4TW22Y0Ptn2WqTd/unzreOJtg
bz8ZiSSf+m/4kytml4QIAxpOZxTw4vQul61L1tqBfWCVJnSOODWAKXLGAfLvRZN4
R9txIK11WeopWVFeYAcu07eCTzEB25Av6MarfnXmTMi8bNsNWhIvorMmiP6DzlyE
9FTZa8m77fAa1fZ8gmJA2Wpuw2xvsLJOBDW24KVfieZK7nmYO4XvTjHkpx53tVsC
FasdJdhX0vz4KhFnIKt4ZE8UFZ2kIqEWTsIc0mpyiIIH0wWcEkw5j4FXsGjzP+xh
1PrMVbIcTrfgM2LC971cURn0vu27KEym2nbl0mN3k1kVKz7ZkzLhI9c74YIO5W30
GS10lzjEZtUqqEfBPcqMAIKBfBsMH0vF0KdELgCEJT4wtOQgRv7ZzgwDsj5VU59P
lVZDLF+4AcWJEc0kGdkiyViBhTswQSwRATTCMP1Lx3lFg0MkW7Axg4F2IsWgborW
zEis1NCAwO1GgzMVuxq0pmb1/uBcduGrCHJY448q4zGQsaW+9U2APuO6X7Med7xS
TIU5OizE2grNMM8tbNnVZV95UB2OvtbXVlHevV+lhhbyb+kPp2UXtqCqZTh8aO47
li4sEv6Zr6rn+FOrU6HfTI3FxIi5c95rqFU4w+zxzYHsH1YI5M6mSk04prDH66De
UXh3uvUyw/4a1Exdpqmn2wYXNtOv+nTeLV+qyoJD4dfakCwU8pck0mw4ZJwrZ1FF
hkJVQR1a16lHC73B9HzbwohS+m3Ya6osgFlIHw+sY1XrH/Fd9Odoq8UsVTfemMdF
Ab5fcUInbONbkRpySZDWHVuVzslDDHrgU82Uq0qrL/X9UuiXIcgaYJQj3hbcHTNt
W634wZs0Xnc9a56JWdr5YU8AODineAJkIfIcKGL03DAOfrCEJhfFOeaJcuXlqkwx
AabE890x1OxdfRxXqf2DkSylUCeL9jBy3oTq+3KVjJVhT2gewzvBTEZdRkQpwC32
/5AE3BPQ1BuqwVRS/H+Pdew1MFU8Xng7rRDO6J6y03ClmwxuO8LJLoTUQVRyAiQ3
RDtWTePnucYLBX5tDR7bzQNgsRkvtWXE1FWyYGFbh27b3ooXZgyqKNl79n9XceTC
8AUhIz4Zd1C4WRKx7ndbXvJwshn490nsmI11P5xxNd+jydLcRitjTioRJb4QI5PN
SAcHr8qRikrCz9SW6B6Z5LeFMYcUGSdxPG5FTAmviH3LzeaxB3wjS5ZAfyj4FOYh
AycE9u73NV3iswWCn5O6aGLV5Y6R5441dPtYg28ly923gi5yGrUEsUM7nNQZlHVh
s0H3PiZG0FQEmP0CHkOTv1kO8an3WrQanzZ3r8LnV6saxSKYLbcczhHy381HCJ1Q
Ra7OJPfliu63NCOWC0KlJH8LbK5bZJvVR8ndMaHiCdNDlGSHZcIigrtVqKQoU2sI
/Gmsm4Yaz501+NOPEa2mgnZccQjxtffOo4JZbRFYhZj3qY1Yv0T9/clsKAeOLEP6
BqsWs/L/XDLqzAqibjc6mRtNNl4AZF8brNdpT/+aFL/rpA7hnjEXS8mvrFInzw0B
3gbSx8urFeU7rqpTJEUaPHc2vJDlkU1eyVTVu7l827FAoCCnmFRac8t/oT0hS1r1
+qaA48cturg9IniUrkf1QOs9/YG8iqozIdQyVo7BCLI1GmuKHB+Ra26dXZ4YUj2d
1oCBDm5yJ6ljfaLa097k0MA3SBALqyq0pCrkYhM3mTStZ5GK5MAwjdshPFUegaUl
mdZjqnGx/NPCq8sFA1emJQ2Pdw7ZsUQnIkWkZt3WL+pZx5vIz3KZ+NE8y+neCmh8
t4IvjFJc6DkUFmeuMFmS/RLoWOiodeQrULq6MFVg5jmaGgu+hAgO3IajrfJJ1QsL
LREKsp1NfnkmHmTgZEWoHBRpAN1vjxw7aZWB6WS9bS7cpMJj92U/8iozCCl15uTF
EOqoTM+yLANAwi0psmtSegFL3GiMkCcT0cPJQiC1oxzMmVwPMiibxqE3aA2d/ltj
GggwIW9Z1l+jkR5a6rleJfs21tFrk0+FPCxaNTQxv9WZi4x+bpd+Dwe901DoZylz
yS+kqQPZpFHOPtfkWNPv+QJ5/C8V0Ke/fP/gb98qTskJBoYoopuwrKcgmvOxU9pz
anaOSGqPUzpZmF6WKKq9Pj8kWaDvR2Is4ycQtmuTGm/DlUgn614vxftG1mMnwF9G
tkDLqYxFA11D8F6Ui+NOrut88CGN+lLT3l+Ex5/WllkMQ+udrT9DoneCHnaH4qvv
t6HRi2gstptHU29LpRYKLKeQ5MO6sHsjgx0felZHSjWT16bCt6T7dSd8gYbA55K/
DqqiwvNYK6hVXf9NKWjIvXeieG2rbUOFJURJW2Dn+UTIkMnA/cMwLC+7vTWEQaGH
Jmqs8vqRH3Z5iVCTlrKbv0kTa8s4igP7v+NvXFFPQi9V66VMox9eluoKOT6UQNQO
kHGpmZtMsC//xCy63SZiWepKfibgHetudZBzilkwTRiw92Li0zfNHB1wSu6dJ5+n
lIUvoDCj1HxkPeV3ctPgywp+LPHxFK7+aSkAcvwz/z2bkJvLhQBHaseOnWqx050P
OcD10H7O5iBDnin/mSUwojfpVwKiqWWMGlO3IxXwsTV3jHXiDRZvwq5vO+UO3ys7
5ttuCyYiOj2v5Zh2rsdVhX+tDCZXCe+L58a7vrTs6QvWwnvWMLFJJAO/ugy4QVAI
ddV4r1DpscgzSmJY3sVdWumIuuG8ia33VtkYYIFsVABiXy1vsPxtxk94MUJcqPOc
uVz0dnYwnGD329nqgiEBf0nktcMSyoS/3pkDpILTb4Rh4qUXpOat9qCFmxSBU59p
9jKIgXSG7/do51xsGGGuJrYcHeCAEu/NLfmBoHGcw1tRnAT1MvKjZtjFdaim+h/I
HpkMdJO14sGfRQeElP4kL+kknMxIPLZiO3gbC459cnx1wtT9cXpXTSTkHWQsF3Yc
7QkPBwuDxm2Cp6D4WWLfiXXP+7izNwbngG5ngsiGLuYYaVMr5dWgPsj/i5fOzKxq
+DnNsq2K1WbpYldm0qHd1+XmqkVt+gmFPeAdm4LZTDux5aFIxcqbgUrzDE30TPvo
ZfGiBtXqaainRVJjKeTFN2HfgHaeCxYruBx17W+uprmTbOvexyq2f3t983ElPJyV
PExwQFi8Jt+X8N3TlVFcK2Mll01GFIb06HoVT6YmYha9zuL3ooTNRFGmOSaqE6Db
VxHRFrx5aLshc1h8Rml90fZ5PtOL1urIOKzN1eBZlZojpPXQcvw/U0ua7tM+xjg+
wsehK2rSBzD26o9GOPoxk5lMqdVSezet4fajE6iCKaw4cqMajUz1eA9fRuhzs45H
1qLaZQlS2U7G0ekEONGQwWezhRwBEaRmQQB5L9BD65RBmh2HRjJ3ORo+kKsnUh8j
cvTtv8hJ80dgf4kD0YvFvHqzpd+HQ0o1USBWITEouhKEF62l9hn0wosF5p83Ofrn
mOKJsJM6Y8vR9LKhWKazn8qOb8yJT5vqXQJjeCEkmcbEgRjWPZiuPaIExf4a28b4
Q8vuM3N6muPxQ7mjh988s6gfVbMYRFp5PcN717bJIYzUh6FORQ3SUXYdEPBWmF/3
Uj5gL2PC9asYzhAQlMfnS3GpjKYRIFQbGeZBWn+2iE7SVCorzU9X2j6+nyej9RKl
gBenGq61vGM3GK095ygr8sc/nfJPe/X26VBViBkw5cLiH2+NeFF8sl0BN/vzx00Q
bUb2H51+4WSZOElZdLwS+h63g7X+AmDQGt3aR9OlC8o0PIgtSBzzuzQdc4+cFVye
4Xqu6S197P+5xZQtMzKiBv7LfO37KAxaPsCWo5rsmJg0w755+dAgl8Fm7eovKR8W
h5IjFE3esyGXV2mZBxvBdGb3wqHzjxwV3hjSHX9ax0yoWPjdgYzr4qL8/TjbWFMW
vz4yA0OjK/YlzmutBjGzSA5ONxKrdWI32r2ZuNdU+mExVjguOYgzLXSDA67yZChA
gehWFtmSHzZgCLCEiQplTOx6vXfLbYQeV37pQ4PettG7JHxNyedb3gYscRsDSw74
wQrO8PRTuDz/zKo8vVRcF3zDn+FYr8WSQyO2k4axSuWeAQUhUI36S+GP1u4qoa3f
18kt3vi3JvjR6y0A1qG5PVXfjh/YIRaedKx+ycirAB7aVmLe04Uonz8ALp10mEpR
PR7oRRixlACywJqc6tWwXRofQOi+sWcFu/q7Oo8oZSdId8gF5bVqpUJo1M/Nst44
sDDZUYYGCWvT8uPf8PDw3a2zwfWOGxR0Va9s8t36RgqjuDz5Mbb3/Jl7UA3AycF7
fN4btUHLF0SwfRcjDgzWk0jW52nSoL7v6pRKeya7SUzTDRUabCReO4s+qfCUocCL
DZdwEZBlumsWie/ss7HJ90Wy9qu0ESkGt8sZ6+GO6vGmngDGekz2v4N/NPVrnDDv
bJEXYV7ErNFsDb62zaykG/tSP8rxNdgXif0IrejK9NkEYyOdYbCWfO2Usjs6VkF9
Utw0TFzfNCpWeIgkCpfJUW8CUOofi/1i9AXgTNZC8ngL+zkCkUNm4KNqWnu6b5Rh
8Aq75Eq6aHsUCNDr8rw6q3Wx+h/zuyzIeZHcaYc9qImOL+VjniNyf1w5Ne8cIDed
ebPdMJYn9T/Rkj6wz9wApoqmEvYdTnFOA/mBzOjIb4xJRVaU/4jZblTfc3jXB8U7
GJqHMHKJrWzZqU7l3O+Yb+JZJnZseCkSwBJCK9CEaPXrVyFuJfG29vNPD/603Y/V
H6t3aMhlLJDNMfxU/ZEi7pCZ2P5MzHErJKpXiHcWAOLrXSNQwxbbenvr3cQVH+mT
bpmELE2mprI9gG9i/XWK64jY+cr9Vxx3DcQHJovvkHcEOcJEvIt56sZ8mZMGq5dN
zFvc03xpGIF8kphR6i++UYjuBomxhGjMqVjx1QOFS0EZ8XxJ2IUuzDmgxvC16L9E
BH2yqNPsgmhSbHM4z/yFa+pr0xylivNPIB1pttbKlHIPSaW5Pg7ptjxDzm/D/D4v
r3s8tYzLZIxHZolX8DhE9UH5snbyrGV50hf0Ur/uIhxkynHTOYmC17gDpea9CMdl
Xh93Ni/hj83cHEtMJGcd2x+CRi3Vh4zK9Re50EuNoNsQRZC7/m13YMO63NQLdOzC
Ni6SkL7dPU9pFZybl2ug+8i+uIUJSPH+JUIT/OiJ9RHQbaP1X4Vd1r6pRGQeGKi4
ZR+Tq/fhRFCi8JKleAjkOEesa93ZvbAN/RYr2sjT6S97VzKIOFW7g3jMWiOwmEMD
58Jry/6HDj768lFknkvd3EIsbMCu2WqFFDStihOFQ5gQqSl/jR53T0U69xzCvwXh
Neoc2NjJf1+Qq5chCJjvjSxOCVGzNemJczwbR6U5TRYwajnYhhFzWRQ+Sa1Ujl36
NBZmrNA2dbkRPOmirrgdfaNcdb7ATuDGFPQQ7ZwlUBvotMoTntVf4Cf5PXaFbIqO
y03coF4sZqs+WYc9ARD3sa9cO4Nj+/t42GAT2F1ymeUk80CNPB+BOlJV0nj0cq+o
d4zClePZeIQ5EKqIHUJ6XJfdpZAmYhkjX616nEPjA2LkPots+R3DsnmwckKcv2W9
NJt4RrJixyy/OmHQ5wkPM4k0N4F1zOXIZhW6QFoHDcO6mNvgREGND4+ig8qlcCL3
nCPhasYrCHMLvr+i5HhpaFZOTGm8m/QB+4g1YRc/A7RtqSuNxjzmM9yK7Z9IuzQL
dVr5Kfx4Cue9263iiDkUn2JiqWCENb3tob9U9F3pHzv4xulYpp9cLi13M6LEnBp8
mF1N+VUOJwBf3HprfqnZ269r+0kMhFS9F36t+IruW7u1gQoWCQpUsgmADlMrz5fE
+bMoWAILUajoL7uv4KdYIMCE+hUjVAZagw8PBEhpLJPfksj78UL8cAhAFX7bdRgw
CE/Kli/q6sdOgfaU2/I7qBe5U3E1p9aRopRt71kRxwp08DxA0Gxig2/5wKhg2B1O
hrR2M/eJkgabDP9FQCu9DEpLrfKdTZoVCMqXuogQM8GgD5misOAz1jRpReJOv3ZO
QUkgrYk6zcnI2NLVhlOMMonnyQ3nQpwg7BBvBM88StEMgzGV4rWKypcqjrByV2qB
pTtN2nxbbwbEWxmUQUh3Pjswngf4qTDdFezz9Au8fNGjgSTuTat9ebbCOkdySfdy
qICd/SWeod4kNUY2zeI3KSW9w2YzG0EIEzJXMNnuHdBKNThkFarzmSk7H6axNn5S
xZhC2/DJMgt3d1J+Ausf0myxv4uwsa2vEISzBDuXhTQ8fL/LFK56Ey1Yp8L/Ck4m
C21R6icwmE5cpJxnzX3CcWipgG7ZNArWrcOJtTdsitVJNIp8BuSK5Z7857j50gG3
hK6EKjFW6kSD0PRGXDWNfPHLQwxZdLQQMfkQw6lhPNIcX17OCDiONxDaAje8V2yJ
uSBvqIVckGcW6HiY+Z4HbxlonDhxUfg6OmElWBNhj1vJjFlObx3oxl1NE5S7lAYH
X1e7BcgcVpAGZVfwoXzLloVASDRzYNt/ulYA5nACuIH+y0Uy0ke9ZaesDcN9J6Wj
6vJAMVsVxOevM8HWev9IpFg/6xZsGLIvJAfapcmDMIuJv7KuqwlMMW3HjuGmRhGt
5b0iHkcaHbwyP/+WFZWB9AhSHEgfo9aV0v47AYoDMrdwFCJiCF2TNokX3P15exEs
5VnxCyAnMFqlYKPF+H/szU1ntW6Tqrgo/V352fc4DseM4Q6P4h6jYsDOs2cOk6BA
U/PjIYaPbcajN8YwH/X+8FtgQ3jUvWRFX1rF+XCJi+FcjulU6a6tqy6ipB/aeV1+
t3WvtSCSe4IXm8MiZQctdG9tZnt95EZ2JtBmpZr8RJv5+9B0n5Ly59z3f5l+8Im+
/b9MBlDq+HxGbN9M4hJA8CI6WuQZF3xh1UQNWdSrJ9bxz+L3Ajmzjmy1PILPMtnP
Ch7OOJRg3NOFSWqAJHV9XbwOgjbypwEyaE55AgUNaVUMi/jEsvdA8uhLoilRWHDN
zLH0sgnOx3o8kJidXW1fPD8sqZc5G3csaZfBvaIQ3PurzTPu2iYRm1dWaqHJowmM
ju90fxMxMswOQKye9JjbO+xPlP2X4J6y/uAdHR4dKENFfnN2EUrLul24bj+ekmVo
KbyGJRmsXJdYUDwRsAOY7Ut46Fd9Y5YueG+XCh2ojuzNL7z3y70lUJW8l3Q48H0U
imACXQen3MgjeAPBr9hRWaDcMMkWwvpfElOYUZjZpkuB+49gqK34U+5Rx2PeI5Bi
97yPzVybtmRRg8eI2rTDKZuFqBptC553scX2bA41ILylgRRyA8Tfh8vPkwM+IvOT
IwMn1khgdj+DSWrBiNUhgf1k2af6B8FYc8WSIqU8uCrzOsWJvZbM0DRMonFe2e8f
BI+Aksuqyasb0hkdrtdpi5NLsC8MW98c8oFWSQiILeapslP0rVqi4ZsD+7yymj1i
aUABL+uBl0AVe2+tloTAuBIPhh82ZLGonMSTBHMHD2mpY2rHoYuuB09XyqbuhgbW
Ck2TpIAR1qdl0TeXy/kbbzipO0mIxccgCNMSBmcBT1RATEhNCfxC/KXTHE+IeBFe
mjo+IZCBYzu3Lo8m8+hanYQPDKjVzbmPMad5xv+QhQ/R4w99VGJG0hgtU86jfLDU
zUHIcSL/+tHj6cCct6dK40tuiIIvjVm4Us86+8QpXgzUjnTemaRsQdVxURLSVxpB
lGKHLOmAQWAsmK8UhFUxSVrvQU+oRfnUXmKtQC+tyoTe4/pbYrezUT0hPkswZUHd
5otdfmeAnCiaHzsfAy9YtHW1YLe27ke+QU2wQkt4ekjAUcbjm+o4MaFTQiYXC7JZ
cGzBxtCWBJlSA4Uh3KZVrV8qXOynWHsKZBLzkWi7wNJTYJFUakt0NKMdrNOTF46u
TuYRugB80OLp1OnS1UI16RLD8xbYFz03z8sv2Abl2P/Xn41JiksTmSh7AAhOtHYX
rETsZbdInz/lzBF0u/5iEUFH+U5x7+phgFSrZO00MCWcQxOJ04r1payXTeCbRVPq
oCSuK/Fks/VkOqmwBgexSPkdhwPE66xd9n4cGp1rWBaIKvk9HcKBlAewdJYGywjJ
oMv5gNgNKFOuz6ql6pIFzZW49fHJJVIwj2KIJysC4mhcndls4CDLMNZujuVGDX46
2Ibua15P6HTQywXaZWPPXhh3S/Tf6FD+2TZWsx8S8tsOUErLlF5dW+r70sk5BYzf
ww4LL8rQNO8P28vwf6XoB/i1i1tPuUHJ9cmgxzDBF0qhHUfVc7SdPFB5kYnxree2
OqRqHxyO60+0w3SE7zM8qwgJczBfQKOzIxkqbYp4Ex5bC4VqKtAoVqB35vIM7sCJ
fKTaLxaWYPUYsEVhsOs1X/DpteD1wxDPaeNbqQCxLdVNsPweBDZvCx75e99sokRq
eznDrbI48koLYzNJIhbvf8b0Ai/YkCbl5SGMmVFXVauttNRhYj7RupU1No7jmMUC
6xfL5VCsn/JcbvLlmocp6ck9SCCwc62TMxkCTNtgLsZ/+Z1M/mFQXBZfd02dvW2Y
a+EBt/NXsiL8I4DcqSZEbbmc3kjP1eam/2B/eYJwXQX5OXN/4PZHpy6yJEmJo5ay
K+ZZB7Wixr5I48IyBTRKYm9FlQ8Jd9ORU/HME5/VWuPCMLTFOEUH2DSNxWTGGAnv
Jt/rqITe7tzUu45jtoQMqzUcSMCPrKLl/hcyEUPuC5hElk7etn/zBQmqtFrE4JCN
qxnmANPwyZ+qhC4XpTMpjjY52pUeC+AIwpcbb9h/W6jA3/3vAn6Afv9p1s/v/6MN
TV9yisdthAboZ6q+MB7dhEbSnwr6oid2lgECh+G0rVzlXmLfB2PXLEOpoB+ZabBN
44WPlrRoQBkjD4qsdPwxbBs7RwfJ2UHMCb1hkBDLJuOLDCiQ1FeIAw4FUSsDMBOX
Sx9htR3KePJjn6Yuo2H7Ry+v6Kicyxfnj1EdOggqgI2PRUT0dKgJcW36f3g4SS1k
wV01/0YQn/buD1DNwROXg0rUBjQGmCaEkXzqBSAGKVY2KaoPp3Fv/pG71QIMJ3tS
Bf4gQdGSVy1b7Jk6f4p9GzhEjd2sXK1gFA9pXVelk8vhSLSbdRKie1MwFiQ4GIvy
OhBQQx2X5hCrvaNrXByHvZjxPWNUVBfLn5E9LmAn1P0IRLjvOyFkgl4sYzMYjUow
GeAHq6wkoAcSQBgbb0cUbyLNSLTXdcgu8sThyEZP0xRzEfp+YWW0TTF1FkTpfSK1
aqxfatXol9C7okjG5WdoonWO76qrjAnoIXB34gDs0eOdL7s+I3CfqhyDF+7eUpJq
Rv+oT+pMAihJzJ3Qyp46mBRS9PGC+xLo0Zp26ShYQBQ2f/RnH033WJ4TWnpMNzJ0
5eNha270eNLteF6xfs8p5qr3NeY3z9hG5y4itnmtkQiUumbo9GFzJceI3/a8wmIF
hKoQd0k56KYD2y5oQSmiEeX+5vNngAwglBxTcIctCKU1ZkLQin5LBo0Oim1Hw1gS
XgTcVg5fiboz9zZKifVNJm/gTj5vFd95I5fcA5F6Vo6HIxGvQa9g5XfkLWFkmKXL
XNXV5Y0+rqKZAKfOWLOeW2Lmn7rpgK5Lx4gBRXH4hKtM4zr5Rp/puC2Nyg+HUcGS
wf4e9xzGUJvOOgxOBVLEgVPtoo590ZjfDsuu+JWj8PrZUZDc5ujJ8+7iuKllVDqX
GspQnYxgdaL+hVIBObr82mUNXUFaqCHLE8I+KcnGyHTVvWAJxBa9Nf6C5VHcfCTK
qXpMl9NImc+K9RX5M6/3EYKBWlRfC+UBKHiW/sSWC9AGBHGi+Gf4+a9iq0UoSmwY
LS2r8+KQGGaEOL/hgYJFL1Y2Z6hFmzVJtXxC+NCICOQPVcmtudeNzcDHQVqlDxF5
6ToU9vioHF6IUG6cFCbkjfDJ5OL63mVvJ8mnGxxFFupuidiZ2+jAl//XyrknHEWW
5PZzFOCKPkivxROE2uetSXlSUKQev/pnu4VzAbjQwN0aPtl8NXL6z7Jlln8zOCj9
Fe7xC9C74GLIySeg8kwhM6hdGFF6fCA8xFwqNXbpqZ21PxCc4qHSmFzrzgaX71ZH
5TUZ/u0XoVqBwzngJKIj8DwfGXL0xGq6Um7uDestXjlxkxW0cN6oPZu+shRU7i+X
oDTUW7dhvPVSc6ZWGjjRHJVYxp9nIvxYc51gjAMnfxdikZkh1QbqR40gIXC1rQKe
xxCCIsgJPbv9VsSYYDYBmG3d86nDaANrG2kZHy4rreDjvOzomvrtH4p5TC7AcYMg
ObeHfsaA4NtC38XKnLX8eV0lt+rbqd43h4usEJYE4DQTDeAYr2Ec6CMrEJSUfr8b
E1H6nte/g3fXm+WZQ6C5OGLY641CWhWh3jWQbM4ZAxM+FZzuHvZbS5Pcya/RAUWr
kv5o2c0Gug9eYCZr9+nPLn021CLArVUA5w72LknCZ64NYxO08vskfz++wI0ogZQa
00E18gjv3ZvmYJZRcpK7P+O8eDsKrr7Ih7QjY4nZzMHOnb+hKWAPEN78t6lNgZrT
7AK4+vOExkOLgB2oeGsBOolsP/emVoh4YOaytDelSvt5iOvuAIHg7v7uxngvensZ
dB1vdvTKIjORWZIvz6TLzdC2WT7JP8drdUyWvqlChepNbbrRQaVf2l5Zs9fEjGtD
QcOBuBa8lIspwJSfbWfj3lzhxYjlEgtpdLXomwBR03PfkyMYTGMLmDX2il3D+dFh
DME/njAsPe7Zu0VajFNnTtaZs8QZu/ZpIHUn0TrrGj/ab9bzNkESrGaWMe2PtKx6
uwvDgIJnFnX7t3luE2gLoglCKCm/91O+jFymHAoh2mLp1uwX8wuab6vUWvqJ1c20
tS3A7iallnn3siJs648NMM6iNEKINXWG0gmyEdwnQSL8pseVQjN4qsNgtGBUaEKB
vlfNcmMl0auATAwbkgwUluvIbPpbb5mNTg3GZjtcRudR8f/0eSMLSq3WNmjG/j5d
7ZBTK+HwzGu1xolTUm6G6JLtchPuIPEuiqC0AFq7cAuoy6SF+szXG5g340GQCb+6
8ja11eo03qUT6OBfCtbh6ssdt0ahfsoMz6TCwRvAdY/yG5GhE7krBizhPZm6vv+6
ClFDEo/zDtJsht2xTudzoDE/jGRtpIO+ZLnYwJh6xbHCTO9ALRahoN0B0ErQ/P+9
7G9i9RwomZI40B1xrpCobdPPMkgDtNUE2BDPHpFO0tWTfC3DnfJBrgEFuuySD5AI
kza1d5gDPOTPDrykapWp5Q9fx3ISCPPmiegM39PGuiY=
`pragma protect end_protected
