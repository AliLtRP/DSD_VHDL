// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:37:18 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
gisjBgF3TEXkNx97MdWspMHZYSsEpEC6A8nlcDwUF1Aza/ZvhsWBeQz2EHM3qA/I
kDwQFXCgN13klNKduhM2CSmbrqYd/i/3Ee/XVJhCcm5a7yc8Vq/GvxA8HfRcN9/K
9o4ibOmDfjyoRN4t0Ha1IfFRzCgt8zNowLu6rOznzi0=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 7632)
LoUOok7nL2989gtbaB1tLcYR8ZSyyUGHg0BbdN5daphUsQWrgvbmVPbx+HOoY3jw
i0KWs203L+MCQLmdwbI3DcG1rXBegNiTyGHDa9Ud0pMpscutclhlrr0JGihYXftr
yBzKB9jarPrmUeJVbwv8RjNDS8p6FJ/1lwDEysqCANWtFbd2bWPgOgD/ONSGxa2x
EThvWrmaGs2/0aRf3TapB2QMEQY8YShED5etv4dgzOcbUjNbTHa7DtI2ype5qCJS
ixXqNXYzT8ItJqCpg03gqAnW9uosfUFbO39uYIekYnQkhCL0yVI9dO9OTHDyivJj
A+lHpSsCr6QdFq+7BbdQPNydcv0glG/Zkk67IX4gl/LmvqnwPoo3Ts70Ns3D6vdR
5Rerb36oQEHCkmh7N9So2v6/pb45c/7QZ2AZ+cxy5of0EXkzU8ZHerCW9cAcD6ov
Xv/tnnoy3ljas96/VgHnGYygFJ3v0s4av2GwpHxuog5+Rp+vaKehRYMxochO5H+a
3Rrkcr+cqks3F0SktJBxVouaoDtwVW2DWxK/w9dZZEdOtupenf6uMlrnJ8MKoH7n
fpN0nJxe/DHdTFgUMOQEUf5ch50DXoNg6bQ+ULJI3Mi57+dzEPnKWMHI88Iw8w/B
8mBqHrdy1gX/cEpHnjOQNGgg5tZ0dnrdZxPTdVXMVqgPZ1wtEkqzq0Iiqf5yeZKm
lp93GTO/vjyN/vhQ4XpkKPBbDDkHmOGvHFaQng7ABwQR5pScKboPFku2hDcBaLWq
8L4KOijpi/4UDq7ZgM24b4JQ+cP6YWjseXZJCSYU0TMsfwhG+1N5XNJZ/HXuzUI+
gv0q7TKncZD9dLRsl8XR6t6quyNwZXctoK+NGT/766byi9mcm3I/rR0kI3zVxwN0
cNKZ8gbe46uCw3Gkt4cecQH7wMauEir3/+PRhE0MufOh2lSjvz25jaGoU79yiwya
dif7Fdkj/ypQZxA+Ci1Tffw7VpOmLUOI36S9htvj0HK3xysTQt640QJ1MiQlgKOL
iuPe+PzfdyqK6rJy6IA0mM+KKqb7zQFmnbkK6L0IutKIQStfhAF93ogIl8oth6k8
HFJR6UFQDYqhbeytjG95RVVWvJQI/nRok132dS/DLQUPhmQqm1L4n/gSZMAnXkJb
3kjAlnD0wJNU3rjFLRHBXAIeETO7TbwD37+jnxfNMAgXw5Ajg/K1Lr0b5uQfbRXJ
QCnlOxJCTq8P8bthdTeCO9d157lE8mDwsoMgfFv+gM40GYpd13DvHEwGABb65U7C
/teti5YCaJssgXK+RTtzXOE6HV5vYHTCAhCh6C5Wz/2GrIpogUc/ivdu3d1DIikp
OWMp+kKikTxsydZsBVR+87PAbrkNUYivBjDz4dqipVjZx6BiB5HHwbnW+uQbLvdW
uvE67AqyTeucI83yRM2BbuNbvRQum/2uaD7Zr8da7xejbdKNk2Zqyi6xpBA27KiJ
j/uWCf135X2Gf281XlSZNrlopS+yJC5OPCiqREvVT53ZRcDNIIwO46rxWFGUsAFL
tTWaHeubk8UeCC35zpmwvl0Puat0N3VVcWjQgRWEUx0C2MMeSScVVs2aZfgoEzGJ
Cgks9ooqQnK6Jsky3RpeQkGVVTikmhParcNRzAlCn8aAo3h+2UFQiXBR/b+/wuVV
7DFmAlZ4NIe6fCjrXBL6IZW/ylZ60rp2Ixaec2e6aqC1MSsxBBchFKaPbaD0gSGS
oOx2DfIFMWwteKUAhL1+qSltx7Xz+DxcHwbTqDpCQFJSUnoMmg3j0+1raZW+zLrz
7fGiNPisXy8ttn5o4CAaeafk8KdzGLfmPhdgEpzyBUtLbJj71kmr1aCgxMl8jpqF
Wwxexw2pVZ5dbLEcBfGN3pUmHmpFJRP5RMkxxANxCjlNLkA6wd5CxItP9eibtBhq
VEeIoa9mniLukHisKXU3UYw3RSz9REBI6E2KKGixljzrscTZvoZkps4DkIxboC+e
dSeXMIwpOukYEJLv18ZQzT3ytcoH96LRZvMqpRa3gFSfDtmi1dtLITtLu12bijht
zRhxxb/GjlsdqyA3P6ezWLPjUPEqXvU4atTdugRA5BaT8RyFcBpSEuXdo/fYcbgz
1k75mijkHLj036vShY7zd4KEfMaXnYVpm8ThORmYp/xILGPYsGH67PXisAeIdnYG
8x91he00adHc0LNyAy1MnQQhgdj5Skau3+s/I3VvGqHX0g5W786Xa8GxCTC9IWWt
eY14SGyDFHzIzxOT9/bzvfG4+0a0/FQc4usTWOyH/36AW2Kfc6oxwfjLRDppAkis
hFLmEMEkdcKwzgmCntaBzdw7CJB7yBHCK8jbA6SO2i+OgKPytik2OItbWxCNPPoI
DrT/u3W5Wh+z2go7gJdd1NtHZVWyQ0F7ML0EFCN7xWoxvpFp2xYOBcP7lgLg53Gi
7NaRldmxgr/oIzomsKSE1FTzwtfE1x4RkcFGJu46DSkT8nX6G5qEQHRZ6KzYhdqL
7GgcvdKAJj0tJsc7c0cDVwshERP2JFFniICE1o8v947sSfTgHGYtHy46XDHsmiTh
b+7mAEH+0AjAldVS5Ies8cr34Hks9mlQ8CMTeEAFHEPGVpPjijRmKBhxmRFsWKjE
7Ejfe6Fu9kIPJ5fTsIr6G2bC1TthMWp5saWgK58wkv7LZrjTufK51wSqVCX1Jkpb
vGy1AafZgMewB3XQBri9qu4pq8uPGNHCk8eQP/ixnC/01v93hrAaY9uNGCc/qSMW
P03M1+r4RpUO77f7nMKpseetp4IdoRqh9mfBnMXu55vPwMK9pOhMKJ7CiVdbyFWz
noiWtn+eA8tflI8iyVVogS6raObitXvrd4nv1J5mIhRTOtigQX2j2jjSVy2UsRPX
9PZlpqsVH6wtQ1708RvJWxIQHxIQ4jwBvEYaPTzWQoVX1GRARvxQ+3SdLH1NT82k
YuK3LV46DJ5VPGRKu44oB3VfUgt4/cUosjXZKIO9pEk7hF5EniMCajkqT68fibPX
21456Lj7/aqAu4gbqDup5WNKizmK/3c0ITXOCeOQ3na8WTRj6ucZJS5pr+eAl4uS
r81sQR6TCjxy7ORiRWytc42dF7Z+Ct8zsKCJQk5tEEf+2eAVaEDC+Y/PgqqN6Gao
wJxHjRvh5nwszrLC5r4vUOvmQuAM89dSHCyG0yhiq7u9eIJQkIs3w3RgUK16cTrD
IejZ0b1wpD33caZu1ioRWlop35NuO6FBAmquNAnqFA/46TQSqOkwzt/4OeqfUKrt
tilLvrBIfLCn7JS699wgndinfWct3TUBIFXHoY6ixu660lRf9JB4vDTAf0UJFYFt
yXsiWgimVGlp+csTFAE+Rw0wrqjzq/9YNwiOC9JTU4ksKIgBL5v0Xtm43X+rWu1H
/mRq/MrqQOZAoov32LU1nvbKepRx+CRnq8xzlSK2/ek1bBqdFduCXQCo/+VwxVMr
mMDZzBaWv8UawhPjZRUogt73RfucHamonlo3VYZDdoglCRgI7G6j52o8WQjMchRA
AgqhVs67C47uDZcX5g+Ixr2C04BBO/rqegCFfrEtaBrbxigiQZeuX41tcelPm/0C
RRxJBMdvFsRnEN6PETMAKVYkslCJTkjA0I9yVhDg7Lc5o/3Qn23z+AuMQ6XeFOJu
IIhOvfbkOGYmY0uBnHB6+q/YKbpjieJXvqKCBjFIvvhOGfBjhwkcbEApc0Ktz1/F
22Vw93+w90HxzfBqZ9rrmdipbh0NuuX6zCa9up+zoqJV4fAwMU7moe+BAGEGmnfk
/Rs2FkWLIqjqAGs+y0zRzSPgQ82AtoHjuQRtonsz1PyQs9IuATII4RRRN1tFFPpB
EGlUhFh7s6FzmrQeipm8jhRQyqJDr70emSqhvbP0uRWlYD/mJzaCka2WTsOHDil3
BsjTYumb3QrM1njm6hr3HryzITDlGZwsIfJ8tNytq0J9mwHoF8VS1eZBd+FBjbZK
jTngCFs1CYEfTz6dk46YsywhfUKge4xg1f6h33mMu38WjOTBQFALJ76RA31ucpBy
3F0+plRDsxMNtb1wR0lnUUbU+0CaMutuDN9RFd0qknUEn73xHB3Chz8hB0zUXMx2
oo5O8JFNA7mm+vdYi8IBjRv18sxsashCBOYxCcBrImOh5ojx9kWutkYO7TusoaTY
cJ5gqiLwGDsM2Rkcd/S8dCKpf1Mjrun8mI+U1ZVS6rCKbf/LEM8uW1zoiV1r/uRb
c7tv4liQG536+/O59eqXn7h7p7C7Tqlf7rPgce1f+cs+4lPJcDq3UdSdxRoOZn2/
989uLk04Eet4r7k4QwUDhpB0v6vmPi3rjF1qEMZ9iiluZuGKIPvvQCuyPPOLKle1
K3t7KFAj8JVYmAeuUb3nO86cJotLcm7mvgovZGYaJ0+ycataPSrxkDosO/1J2Z6p
IsWS0hG898trfkEtglMsUF+VENO2JWBgaH8/aBttAqEFimX2AdsYewjD1OzWbvCB
3/3g0/DNJ3nU7g7WRLtISIdjYZkbvg8ebxqajQrtbEjRfM3CYdq326ygp+I/EVUP
N4MuHE3N+A7WosHG+q7fG33tZxXWSCqXHMLSICGN46bQkS1bElbirsClKgEPMbiF
I6MiOKlIet4klhEgXnhUH1INHm7DJszKceK7ixNAbgnCGv4Cx3yzn3EXUcILAwnd
y6rJi9A1t0pBOoDeJUlCh7QXcoA+sHorc27mOeW6ap2qw97jL8SLq5oIQBSvA9yd
9uzt5GAFuRlChb32ahBPPQ2GbwQnVDXpoXj9pZp1w5B4UQw9iN9nqO+JyKaAGtpU
n3aitgoy68LoPDDbHOVfCq4xepCbrwyyghH1nOQfrp1PPp6s1Ms+Ajevd/s0hlgO
plHOtM12BZzO3YwB+ekxQ6CrGbHIFsXWqRB+F2BgEv5H1nRL5KCNt49CM3L+Srpv
JIAaNh2u8q8tmIrDP1tVObxHZ6wXyu6g72btepkLTKF9HGqPYP3IxtkrxseCscLm
SFFf2sS7Ug/4frs3fbGOKRt96JBltTGWEVxfosXMQwTi8q8EjE89nWXyVKJnanaB
bydyZe1qs68bARUF4jptYWkJjbA1uNuXx1n8F6w7QjAAIEEO9qL20WGBE5ACqOdN
WBiyYU1x6+xezjDNiUaxPQD1NMZZxoQctYnSXFOgG7rnOXamWY7ttYOENLMWGcsL
QdU71dD2MEeh9L6L1IxcfOZuJ9eQVpHdCgdEuvwhFSlPHCS9EPJVIKyp0sngCG6g
cnkaEsjECHBYw1aPnyQ8f3wl8TboiJGcGlmuW/ksAjGr0VLAXQ+bo9p6iteQzOas
JNvnvMAqvnVRqBiERJuxFsc5FCaqsYpbpcbeSMLyRvcL3ImqFpXFN3Fq2/mDercO
eRXd1/BaHBtBGQMPVIaOMK6/OFp918AXsj9v4JtS9VUqycQmRmJqEEeewu0p4GWw
tk2G3pPX4+wCMDV3Ytpqwt2fm2lHL6gbHwnyJsKW8PPpzoCWR06JzxmSDFENjccx
mzxqDA8JgIEYXXzrgcpf6pORFxUWVrYLTHLDrZsUq+MtBqRWcP8e23OwmMZKr5co
YwMClWr6qedxDVlXIo1+BHfAQ6ASaAEOF9CpZRW7vuzK9AcIL52fp1xGAHXhYVr/
zoLtXkNBPN611rHrPviDai9MqkH/TlnNlOT86Mb2+v7kD/xTK9ILLZ1gtil/bojF
b7HtlHjOMbChjrqMKwcNxnNTLTilyVjZ6dsDPLOSt4m9bYUReWmHW+KOzW+cr+Fz
ql+EYsL8oaj7SulOJWCCJT3t3yAF5L39IkTQtyO2sygC2cixPeau0FqbAhm/EpUs
NgUgvBb8V//K+uLasPsmzX+J7eSyCNVPQI+Co+4qbzxTX+A6aT+mbilMVkgQ2ECM
5UcLJmgmPLmabgQ+0OajjQ0MYadUrJmtYkeIPDy42mU9TKmiGpZcnudAa0Zfobik
5il+v05nl4nPM+oChtkC4WOsEh7GZy3CW2l2l6qCKxAXN+cpwn0v55jO+FrCiQ1p
bOjwdPvrkX+IngN4NwLkRmcejilg2lNHvDVRjeqiHcg7Pb5kp6LoNHPYwRzy1heV
E2Pz2BjBn1khZ8a9kpd0YriZIv6ftIPe01qdFEdPssFAA2zleIaQ5+VVKRz0qaRP
BBGKTF4ozJnx6dly1kHLLTH5yX9+Bk3hdfJRg4cLaBM63vm0grwuLMIL2kvYFakT
bH+EFBOr7THp0BzTYsRPJVjNOmj4dYseOmPxfV0rv+6Ul8Uvj9pMprMVCMg8iHVN
jnM9fNKWQlY7G9Lrq6dDwCDWBjL5KRvct3+StrxNNrDnzfPU/ewjsu1DB0vL24QA
hZqmo6K1GUGiPofPw9DSw+ODnOFJiEJMohkuYKN6hm24XTjfqeizdkmnhitLm9x9
5R4tAckJULMP03X15RNhHoBu2YHaxO3Zl5lyKfcrkgbN9b77Q2Hyol/DwHryjRLq
iAqoR9o9/HbMWGzZnEmfZpX0FSiOmJB/uDnJG0fgCWvBIK32Kx0ut20UBR19DaKi
Bea3hakL9z98pM/HTpFXdcMcZXkCDp/VM3vLf62bmwHR9yvuveFI6TX0JpFiuK+a
f8D6jSJHq8iFlUDLaI8B1/rNDngWBTuH5mIfF+Fhti6s5cEx9XRXH8NCXy5dIohz
hWgftx+8LiYfCE+SfMf7HGyaMImrRYUUn1webS8dAEsTFxXpGNf+07QKg8LH9pSJ
Ow+cCvMWOBdwQEP7On8jh5cM+Ka3WsEJs9j3KAIEceJM3hNvpQPHLRLMqj8quK4k
vEeWrn4HcskRGJ4SMTalH5551ZRSY9v639kPEQ52BouvZJ+tHysjgSMh/HAUZR65
T0F9kS+1ir6deQEovc2i3mFjFlLfHjUrfvX95P4X86W9W2P60lZneJ6dL+tz+usM
qDeTY8BVL2AUOOiEzgsM7FJKwG4BUOexo9ftx58fzsZ/V5vEn/4ma+v1LDiu8u76
QdXuHmw0eciQRLYiNNkl/cntjs1gS2gn6b3R8i4ym6Gb6za/s8Wq78e97L30iLEI
STEd8vWFhS6nOYu9Aqi4CyyaWuRGqKKM/prrXZjS1vrTTSuBajlgrImmG5BlrKLn
JNp22BpRK5709w2+OvI83oFjkew1wN+HdA/Qq0wrPJQHcNXjFcoc/kwl/WhOHiYF
eyoXyAWoams1/0VEYCtTiTiK1m0Rou8bGFIIrBDwawTXxxAQ9ogd7DNUpwCz0IAE
yayJqahp5bEXCQaRmX5aIgd44JqMogzZq7qLR6kCGOo4Fd99e/GL383glqN2BfWv
NbZr4iJGErjYaM+uAdq9uBtVUcMD19B0Jxz96Z83AZE8nuFOzh4o7LigEXAe6Hjf
ZIlU+ZWUXpnCBM50YP9tHDL57j8qoNHREY/Tx+RTAQXUhElPfqWdtitlXXFx4OdD
6bHu6tH4XblkLmtZdVYrFiY634MiYBGJ1YpwsluTvJd0JQKBT7reEuCqSqtCnkNm
N8Z2DdTpdAu7H/NYHX6lRQiuXFo0siu2X0fhoDLlzM0mR5WPpNccID/DysJ80X4l
lUxIc/FPL6S/ldWANBzs/A5Ini5yu13SRzE8jYP0/JQlRMRRWevCudz5xd4AcsL/
wMxU/mS7SvifsErxMAib4iWAb6zRplY8V5NFBQnBMjOdvv+2rnbSMN9P4G1WLMRE
DJIMrxH8CGHxZF8TQDb5Wyc16wjZBLi9fCHZnZ2fycW4DzQ7F87kUbHUX5oZsOuJ
Be8+G0HFdn9hre/L+PVqd448yEiCJhz+5KYH0piUOr12bAXTI3tabb5gVBrmFMCr
Ap5VzteK/3yJndf8JUCQ2Iok8lQnP4grcvDOnIZvJfXEzE+jyqVgwLlSgAgV+0CT
YT7WHq8C5nWkSCu/3LpiBru+loM+tX+u2TSgjIE1QfQEaUAdIcsSES+Ucp4zSpGQ
+iAqF7edD5WljkH9INo87Nsk7faRXJCSrKds5Y5iafNMtiqAARbY0SR7pEuJ+sXn
mIodkRm1k8+BwwWR7kT9mUkdiOskL9EeYsU0W+vo3znYhE1QXb4jM09Id16zvNkq
5Nwj0Ro/p/JSyPqud24/F2GKfmX3ZRo+tHMGQob+oF8T2kFS1wUyTsTT5cUATAvj
3DcaN2kWmZcM5ocZi6RGNa9eUsQy7CDgFLnmxFwbwS3BtXwk0DPU4g5ZCTmsIqIR
lWjy7tJzPdeoYZY2njIAh0ytkpi/OJLM2xG8ynvgO0gkI7+OVXcipx0e+CHRVjZT
IwuEpahSMTQBo+CdvUrv8Y2drZDdbTA0/Ih/tEmW335/me/9hL3P0EkAnzvORsPJ
kVn8UksPVNb63s0YG2QrOfFXEcFVH0Zkav7w68ms8FkRxiMlTwOHFTZ5cBk6BvnN
u8RhuT7EbW6S/Z9oX822PDY3ndAo3nMDU2QDzXMSHP4aiV+hq1MfymwNdmm8hdIN
x3iZTg+/+H0bkg+DXAwtW+0sZEml4KjgpkEec6RwN+CUExVF1d+D7jFZ5Y9bumBe
uno7Fx9WMJcohz4qXV7OeUVwJi/4+vKltiV/MXsCEm4s3BFZyewnRMo8n9d2BpNk
y7d+Zfuc1hL7Ugp8/m7aoofDurxHTN/3xGMzsZlO/S2rQ974MWnCKO/DGLR5u1Me
YAr/o20lKiyW4UJSWCYIf/shiGlfF4CUyWkiiswIDdP5WdPGZMIZ0Rm3ifk1higL
sStsY5QJZ0Q/jc0WynxzFFbJ47tGwd9+bIQxC8J4f8JKgcVjLT9D0EDMHR7eLmnc
4x4/5wAWERMJi/6jZMqriN6zsfAitfmLY9uQM9ky5/6+nHvb9BW1l/cVTOfL4mPX
dsDa3voM6CdmBQCZ3+e2fd8/26aDnoAMnJocynw8eY5ZMhCTB7rO3dP5Zp36YUy+
H+hT3Ij8ZLjGQf888f+FX33C7+Apq9yNC4ue9Xgl3hut8wGpGCA+XbZcmxh8XT9n
u1YFNoMqjPGutJEgDo14LYq+gBrq5eTkGDacST+HFWp6o/3bgWPalR+A3xZFi4a2
v45s9ipcuIeq8tWUlbH9AYXGHAxjrwOABymun61uV2jvM92ShODsW5yh7LFKp0Yf
JPNSNUmbezlZY0wjGE0xYe/tM2a8hqqtTph7c1akNBKVusr3x7h/B7dW9LZYhGg0
sH8RnN8OwGEGVoqIh3uRErzV9qaG+tHaELtNDGSIC4XEgR02ZE5ouZrTyNQHSo2z
mZVF4WseNDNW7GjrFWKpSQqnRkV8hgBx9gM68nwyu8eaXpsM4qdqeDAfdiwW/eBW
ccBr+UVOr+zwMJfqhicDXbGDhJMgKQmeyrng4Lr9gTYtAsE5zvxzeeTY+OZRSrgH
5dBjJ6SjvF1lstsh2pj6Hqny1tr9MnEpZdNcSsYNdLnhzJ4OdSai1rT/+IoltM9i
Uolom2Z8QVc1vSiO/0RnSyocFWvXHsHlYetBfswLGPKzdzN6+JnbW/FS/oq2aE0R
W73DnXuxmDNQ2N6coQMHixKFq5LRIsPGpd3Y/KQmynj7FsH9ftlTE6RXNBKj1PBC
TFLOx3R/jSZj1Ik8kwZ4JRDCqc4K2ei38GLVGT+f0hzL6T6RmnLMzRA/2wF8zpx3
+uewObOo09JkDdi1SYsVVGLhyBA6UTFq/jbTytNMoxazFLXh3jxps6u08Ls0bkJz
S5VBKgIYBLJugyzd7ohH/L/j4BuB1kP4RS18ueaifwQp9Ww/u5grtWPwJUw5Z6Im
xWhPOKGH4e7/DLPeqnxsU/jJORtUT2gi1b/lJhm4Yu8vb3QZRhsTMAlfIsO8dq7i
MHnqHf5lPKWZfXV2rMKXlEsqG3y+yhEiGy04bOs979bkVLWyecO6lSzmdh3VwCoh
sGV915tOACpPtkz8YC73cgX0oc58NBpepTjQ+N8+uBLZBssjkBjiL+YUFWDZ0i1G
RPS/f5CkA/62TxlF18fGslucEn8DwwINUFmN48TVwJTByoifsPVtbXmyYUc4clIS
+Itkbxf7xiTs7NA4ZzFcpRPTeYUH5bhTXtt6amCQiOCp7YcSEgmHzWeHDwQwfUmO
Fjojf33U4LP4qlVcXnykxfvjhHGs+WVRUaR9n+QGRROTBj0DcWLpVfEJ1DSc+/rP
gFjJnJsAvrfxjutRU9Xjj5w/jfVYywON5ZEFPubMPbWVshu9JZNAPrVYf9v0l8yI
`pragma protect end_protected
