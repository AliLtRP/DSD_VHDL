// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:38:25 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
ZWLceeZPkwWeKhdUIJSWQG/2DMv8EOmH6pUcjV1bEE41GjJ+rbpYQgbZA+ZlAKfU
qYYKmxjNktCXdybhBS4ZIhUaOLDTmYkkzo1kzEAplUUwYEzTVOu+jVZUCmQ8ZW04
3DC3s5hyvzHLsv4lK92l+eLifrckxTLzGGJcXA//4ig=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 9920)
fMGa6dkvP4NmQYBN8YfcvC2zBHiNxNu+2VYZ5d1XYa5CVFLN2o3mZEffcpMkFTPH
HFg4o2HKyxFvSOwRcm/4jnObFsV+3PJp3pFZ5OkuhS6c9P+RXtsnYzBd+ZygRTZj
jY4o+b/5/JtKejX+Y9sayul9ZUVVPpW/JOgSqJtxKf8YbiJTuRPzuFqKjrx7VTUn
R4M9p0I0BkfJxDOGRCFwibTX/VALv1zK6jvOWFNw7dfMU+dq+6WNtlOJUoXgXVcG
f4l94dj9DHL/RzGvHZeHKvE9uME7tirLTO4OEM27o90P6Xuf/H3PUT7GvWFmLmfD
mhMqIWngwoRZ54P/SRznWrBkrGgnp3zmh/PWgudfjiVo8nu9p+nKEA7HoPqQ9A+I
R6QNo5t/Utz+XD+t3xCP7ufB+X7veXEeSGPAbtO//bf0iroiYrEp74WZ6kxwudh5
2aJT1F3EUERNIy9Rt9ijnEhBysqBSDPaP9OIPqIEPvYzaxqLOFqWck3V05eWyqjJ
XqfLlzmwKaejspLoEuOFjAHidLLgYNWJZT1uVXTmNrhwKEiJ/gyUiisLmNPtQxD5
HxJs1JM5LUldX/bT2jweHyK/yeW7o6rDYuXEfeyla1qts05xqN0J2sNVSSEDp90J
bR6bkJjx13BwpIhKjWnpm4HtKgFvrTGg2jxtfy2WtNe6TB1QumfjJ1hn+xKoB9d0
RL8f83p7J7jhfmgLGeV2xSME3Oyaxcyxkg3QcNMEdOpVwDpMCcpVEWoGEJmx3Z9D
Nv+ASghW1D5dq0UbGzF4I71m6U6PcIo1jqd19g8OdGot3ogz3SWei8dWBnsX/NR8
SR0v3FhAS9olhp6dutRPdgUEwLZtlY1dU/R5toygkUi7/FAI1ocHiLDj2HQgKwku
eU45ttmCSGN8npq+v3C8EGIn5kTixk7MBUiyB949DMsWunNmDiJB/y47cUAuZNV2
uv5jLeHL6oYWFJgPrC6dS3hhluLrfVo7sSskeqcWnasHqjv84KiwY+nIy6rdg0OV
WjIa5007Kd0MhHXWti6IcEVV7hQQGwo4/noMU/6PCenQ1pfF/P7Dl5SPmVhieB/U
QOi+xwSIiqIBhLFkeFmQDW8V/USLWEnslCFmIqJVPu2W08939inzgSt2JB4iOoy4
R9hepfIeAl5cH+D7aJky9UnwJ7LCBfqMKTi56APqpYY+JTSq+Og4oqzSXxR4Kvmw
6cRfQgDiyAb2c+r1BAQAfqTQZOFfLn8/1UQI21zeBrTw9fVB5LTo933UXwEL0j7B
hEzF7y4nCIuEpuMqKYD1lB9+8VEV6/s0zLkI2vwt2SLMSDXEEGaAP2jARU0Sfht8
YwXCjpxrStt07wJO382l5+T/Ps4bzrZ2gZ2BBdeEwpWsgh+UsZlKw9yRQdnomX/r
pgnmKrMFvE+mOix4MYswZiJ5cnsRjIpHBpOH1fFjhA6qDvlCVUg1HmtPaxAbR4D7
Vnk65LjPl636zZeqcW+zdcYLUNFpGcf+utNwoeimWvycYzlg3IJaD4N9qZlj0+JC
86StBsG8QECh/LiVHB+2SunfB435nSlDdcmyq+LIXPB6xSq9niXHfBVgAFI86sc5
lR9ScopG1WdUnf1UB9BUNL72HNAY6L+myre8JOX87VgMyUtswOwO1v9V52P1C/H2
d5ioPUfWukGDemfNhFsgZSV+isHcVyLggL3L3nAsK59kM9CmpYlbPCc26Sh5AAN5
82XEIDfsTlpDInDD0UwJoZm+voMo1nN5nK/LtGcce3a+YT2+5C/DaX0pqiU6rgjL
cC5CTn28eiVqv7yvyX17/RLMRyqzRkUpFZQlT1MQz0fq4bZkBM69P4qDJFqDZR7V
708glmWHURVmoKd/KPjseT3P6gb9BaYHe6hhrOevH3/70sK/j+poIFbj+ZO11zvx
Xyv8ciZlSyE9J4GIA8usHdQrhDHIkCSbcP2NwTG+JUQr1lx5CMeGL2AGhXvSA+sd
KKUl7pLUtaKJFTJ1NBYOQBxXHgx23xT5w1+FGpGugqyOd5ogxTu4gnFSYqecIo7O
feucxi8CL+D9U8UhIQogN/LBimWc1x0zuXAS3/DICelbHGEJJZqW7a674Fv6cpfJ
nX+Za0p702u9Mnyxpn6gwzy0wmpv6I+QjCOpLfdNJEBIZW1JadBgSEcUvMdZGqNf
lIJKzCgpusQWTO2Jn9EZn/6Ka3THzlBwnlkrA2rX01tP2B02nuTSyISQSHr2HCw2
4bcW1vgfAMA5JRy9JpbZt9HvWHL1MDQbFidbnEegvvbi5TK1EOqHdOCR+d8qaSoD
WCoIFvSXF6SK+PO2d7w7xFHKJGrIEJUr/vlsp5D6OaKnr0Lds76F/QagbBGXHIxS
MDauvePEfvkUV9drGCJl5wacCyX8CI27VzfpB8Ip4f+Ks4BZsgn4a2CYR1X3/q6N
jZYAq2Xgpc/kevlQwrw7YeiLiOifT51s2Yo8HPb+HreDtnf8RXJMk6jAPbSyh4Tv
bGxIW7TsIc8ubk1pbB2M9MB0bfqn3YxzKLURz5HbxVeSofSzGyo/r8/inooAb1rR
Eo3LEgoe+fNkwxzz+t1vNGK9gButWPTyKkLp5QZdUPmqb/zrLujoVXu0ga2su0oC
Yf0vQ/wanNESt+4Swl1vLgJ4CWZRnODMEvmgctjLp9nQOhywfILgXCOpNxU+joyx
cTvlMSXSugPvFTFtsYFTkizlK10Pfb8m5K3LOEGYVcyiuh2Yyy0vVyzTbeQ6AzCD
6t1q9XdR1p9HT7Kicfx6E9Ca4wXh3hpvp2MhVc4zceUwdaCU5SXgm2FUxNj1R1fh
UixnyqKwtZkFYotUPx+0/OIN/8xdBEvH9l72aEDNEgW0xSMcTypc4Hf8Sh+te3y1
fLJZg8H3CQoD7uq7v9PJKNnGQf3BIRNB2I+nI1/o64pSKhXO9n6r58qMRZvXYC6Y
VuAEAaqslAthwnDmD/qXEgvfWhl60BQPz1JOBhY9sN0Ca0C+noRg8f2cO59lu5/e
LYvkExhiAyTqYjKtwc7adkPX0i3teFR2uUl7OOfHGJodjROlL+Xm1P32RXp3c4FH
icCkGjnSfmEeTD0jXQFLSBfk8I2M5JixBxx7RHXsyCOVLv0NYPpJF2XZDccbzxEr
vJPR6yoHV4fsXK3I/xXM7HrAh4n4pP4Y1rKi6+6z/BidFtNy0o3efjhoRd3xldma
WC8jPiNR9+WAEQGORSVFnNOsrxDwk/W7cMoFqwO+f/CPkfUc4t6bmMXuo3cyIz+H
CriylR4BKYofwyGUaKQ6IPb2homIuw+sYLL2EeDwB4Sr5AX9Ra1jmLKZXMvLQbl5
yrrHDRGXjLm9Oy9kpG4pnGwkYA5ikVJXVp6ut/sOWmN/bwPlScSYpKXGw9uzjO91
EVfPcFC2Me7luZdQcWpqA69JODSP/zC91w0o1cuNGQUBN4S5DQCt84rY8JHz/yzW
+E99RnG0ywv8mswSPWP3DejlimToJV6xY3PWODoP1DrG1KNsXyE4A6W+n7THCl2l
1J6GLj0FJ6Ia+2EPnzz2PPAqeKIB3GD2N2xOoSsdTG5gBqsHjqm2R0DI5kW+j3Q+
oBLS013QPMOffW1sCxQUuLRS29Oc63fFid9f5fr1nng1FlWgzmnnlZknKbeRYAYJ
xjmANMimA1iv809n53UbR38QEOGJjTpd4WwZpRjtPq66P+lTaIonLaayZkGjtpfw
oslFwPrScg7LeYtng2shXov9yjcEe1LCGYSTSkjHatFa/Ard4hHD1NJMi0XYxjWz
Geh1AlS9XgL1RELUimPptQqUaPMFryOBI9OSkoCuLLa/p+gFMymS7mvtVHJOJaQi
1fddKVIxz5cl6boXk/3Bs30dbTE/h3blRevugWDQALOmyN96NvA/mCPAyLEGCMTR
UozeVY/PFMBZ3kvs/5za+talAm+Mv+HL/OzfwxHDTSKe5dw6VPtkiJbsbz01+dlW
89uvfehGwPL9ZmYIDeab/Zuy1k8iRXjb1/4jdDtNd51eH664Pcm6c91KOlBMBg6l
asCubYnW61+jsHSuhUghv1Bn7nqf0dMNIm9+pZj/E1QYVEdIj+poFaGjYRztKJOf
7tl7tAKt+1VjKmmaMNM6Bshf7GWs/qC47iOThohs0KIdhm4dgjcX3a5g/SRC2jDr
dLJ2wgGwzAJbZQmKLxk49ZVCDJj1r9Tj7HuL3HHncYYoWYOkbOkOIN4cFE1L0XjY
ANsNBh4jVWQyc18BxI3nTTr5LMoi+ho5vuGFVlOfPvqrGdtDXeR3Zt1FG70bJxBP
ah+sqVryBq2O3O3q/LqXCLaPTUxsbBEL286TqpGeJ4IsMYjLZbTlzs0SE/W8W1z7
JAjhBNxLqsaLMdrVIcr081e/QXV7AdGsJ6RICnVlPIGy48xxVFr6vCXaLreXBZwE
UWfCL47+hGVYJZ9t5j8bS9bmpuHIk16YB+ziV7Lpd3A36asUpvwbn+GosBy215KT
UKfLMaRn4wVCmA4FQRsUDju6jgVzsSlb9WTwyp2dqt5zlxZzFX/WdRN3xzmHQu0W
LKjUYJ/UG9Nnodq6NJgqGT++uVcfdn2eT+9awUoZnewI7qneeBVBvihBAn8TqRwQ
RKDyhP0IXco74QelkdDz6fFhiMMf9nP9p/6cx7E5O1v9litDChs7cbs9MljgOh2J
11lQPBDrf7jFfd0BX2q4uHIeS7/VE6DYY4piuz2/uQHQ8oIWg+8h2qk6+9BjC+os
OUEaYrFVmlse7U3Kj213v4SB2ZXDpbsv4i3n8hkiyX33Kcr4a85ptotZuaQJTt0b
YxBplwS6Qlu8U3vago4SMwHut6IRnuE22VkmIdzBl/KxSqKIamkCrPH3lGcUYNnb
dSkpNhRT8S7qXI5es3kupm6qS78mBjyMJLKm6sbc6APx5skdoGWyE4YU+3hawq9N
KbaaotLtOVHw4gG9cOxTpmEarpX4EUsty3HlLuic8ZKOplAUQ7ANVnSVghJ+EDYB
rkB8Pf2QiBo1sKN/5qyk7XPMukwXc9wNrJ5rYUrwYzWdZxr8pLiB5YUwqOLeGE7Y
Q7Hp2cJo8dUSKYvVRQ4zZMiqOCBF3kYH5ztvS5l8McOdprPG6VpDejjJ60UtS0MR
GxOZq2yHHIx4eIursAHbslUUP1TVFmrgWgqkkS+TXxBPfyZMM1M2pYQQJvakuU6h
uNQdXujDcl2zJPFS5aLRx1pmfqjhgdF04DUdTvvPkjgdHccwIWzwxPM9ScKj+Kej
eDsqpZvCV+whdBC36hURbE48Svcb5p/V9Azwmr54FHOhv2IiVT+YmTxq3+pEemRd
RTmpcwqLVKcJPIxVS+tZstePADQOIJrmCbflgYlkgG5ToFOU8wIAMGQMH/P85dl/
vuotKGiZaD7QsdtOI048NY9R3IvffUrIwtIipvxAGTGnDQq33FJ0hBOZZZMKLtuN
CMvaaEK/NiKPArl3P19jKE18eIDyFvakCrCHMB1hYngzbCG1iVKR4SI+LvKoRWRZ
RCV38V3HAC7aaiNUq65uMauHMvUTaDaDhUeYJzUlvKGJNzcQYayCcSGRQbAxmD94
jdOUjx92ks9u37KFy9MPHf9/BM1Tsk+WTzdbewG4MCQey1UDkjpqQ6pCR/bYISB1
OU/H34hhu3PBrwFr/dUW5DZRt6VPunCSJ7khKSSpvTRMUZqgpgomlaCH9b1z0wcg
x9uQ3x2LE59ijiPkYavIVtfoT0J+zuXgMq6RROjwK8t4TOtv5ZqvYqNY8nephHhl
4WHdgU5H8c+nq+3xzv3KH3tIqnNp1+pTCShkPRvHwBOlhK8gmmat0OyM2bWoHCip
MZ8hhnKvhcn4m3/qjhDbpP7QFXQOkmOBi9gEny+Z12kEVWLlMlol4uP3c6HP7fUe
pUa42kw/b81J43OTowDXQzP4fn7/K/lG7hbOdLPXGCvhFzaEoZCYPsLJ86S0E9gL
AUbtNGXE9SGXJ32VS9rm3FT6tzkLz2qV+MiWEJ2L6cH1X3p6ipt49cY1vmrzW6AY
U5AXsLxGRwno6U24INeeS3vh0gsRMsoVHlWPcGuLdlmJz4idSOCnjymtCfDZ7IEr
EiO9rReHyB5FCtZw9srSCSk2b6uelmZt7JwPke9KaYv+TNfpJRjX1E+0d19m9oaJ
mGx8E81Vj1lYhZ6+Fl1DB9XlNedRAGKPeEb85jd7EzXBeNnITKV5e5S8E9SBoCPN
iP3uuc9AGrgIF1oAYZgttAlDSeG/x/wwg5rNNmJ6H3rxnE3D1SaR2VdkClWeSD0r
r6js+EoJCQcjeRGvMKPTAVSudAlTfz154pyvgRAin606biEf0diz5vOTRkVG8f5w
0ir17I2b5mpihiY23rcK38ZBSdGzJ5qLwc7dsPFYt3kwv6A+fKbAVvvzkIavSWY/
KttDLa456bQPTOpOXHaBtYej+B8iy/Tyfjs40sIUK3NCMEJoHIMmmKcXJ/79Wwv9
62sMe584favq3UaFG0UaE8io9nlDODqcKgt+PemdPqguQ++2RV6H5ZFJSx+LfJCm
jlCeK2aIMkh7S0xDG03hf28r/p7vKW36rpGqI1+pJJKxYG00kNPZQzB+6NAEJYZw
9XA500tFjsduTpI0Jf6mBC0HsCRYj6hdozFo8olp1M8jrPwGpZuE9Zwhq5+pxkUA
F6l+8Gd7YzFw5etgAJkzv3xzcEqxs9muHa+tkypHiOOfpBhbwupUDdVvhsKpDL5X
scGhPE9feQeGE50T9Sss7dvHH/Q4UXcSh4wmYzIC9EasEH5vk2ahoCEG9ZS9cpjd
ty7Z6GtE8dqo4TCouo+bGfn/yvb1Ty9bpwcSZa7qcjBPjmCSO4YGEbSdAVA551n6
dJa5cgaCuR/N5tYyPo4EOUVuWvx6DkhyjpLbiY3ONLRHYNqWnXYA3O+b0Y9k/jXK
z6aXnk7PJv4K4t3iwv2QmZDS9RYPEGA4UoQ17ED1/7k8IyxOo8fPjo0ccVllD60S
BtHmaYsVNtjkD1ys2EplFfPNXfCz5lytjw00F96ccqVm4iSrI8KiqThe9LqYjLAv
r97odNUflURdvysIp5QvJaKXM9Zn5pLG6gwD/4g/9Lzm7Z4kZlMr2RsyBDuiM1Sg
kaGtAx/qX3w1Yo844/xCm3zXg5Yb8lRsnUHyT/UMau4n0ZMq1hZLEuRIexwjelKQ
LE5Q0CQmMdCxTocWa9aEi1yHkGhkWMwf3Ep8ehoqPO88rGowSvB4uU7/nrfWRJJt
/+1IPBENLHe6rK5kzsttTgbFDUbYtRf29J3pwT5rY4TPBYiVD2T8p1xuqspfMatQ
AE/B6W7UnCvcUEserN9xcqrIspUKPJ6RwuTD+1eV56grz0lrrcdj8tXoogHEvdn0
EpuVuqYPDSG+b4EKXLZPnqUHMKpxAZGv8O3y0JgFC+/at+U6wMkU11FnahvZGHuy
MFeHtbzH6PFGa70jpkR+Iz6KHb4tTItJRr+2XlsNxZHRdR8no3DpyT2bLc0XMb9u
Q6ZmcUcmRnn35V/zmkwJvrDqgm4I/NbU6ukUdDsdqxBbQdZCnQitOya2u3rOyBnJ
Axy4tmdsQgTn15NrU6EbNuUbX+6qf/kjV298vjk2pl8JV8DvDgRs228o7b8PFzyS
gadg4yNoybM8qsuVlRYV4d0izy8CSEvP5UFwBiku+fM2o9wN7S7k6cLrutpMY7r/
c2fUGxwdLHliAEEzioPu3JvvSITy6w9RPRXjntwwk+57P6GrpOpC8dRdMkIq/HB4
lWMrtMOTrKh7VFm7ExqMFOP/OkzgBYZFSxtg/1kfZWB8fFClHY0cZbe7QRhFzZ0f
XEPKqkxJrmO0BwtPMVH0FAf7cxSlK0HeFZ5e81a+guEeiPNdWQ44Pa6ezK1oN56b
akR08SQM8V/LiRh6JVPKYy7y5U1uWOeU6OGBXyKhqNUjuh7pC3ScpMynnMXBYQcL
Ms3VJywjPds+sHLMoNKNR2NWU9MROj4QccO9ClaVV4yCHPnVl7GyrSbD67BPvHQd
NjnkW56xbffhlUUFPqyqhdCeNmAPaG1lZ3WwYt/Ofa87ahYG38x/5Zgjh5QNn2Vr
15fhNVXDLAyx1BnQ618KFvuzzbHxxBPCnE2jJ8V6udg1hnSHxSTdE750qq6Xc8tw
NknXiFBVYBtfTrfJRWPoa60+DwK/Ne+YMqaz/3xK2zTjVBUFtunn1n2v6DEmr+QS
1k43zt+bwPWkmWRcxWmtKfjXGvey1HAoXJBUVcaqNfV7difGUY/PzUa7IkO6wOoq
aNim4XRuoULtTlQ1qkLHF3JZ8HK7YvvPxcUjW+7ZgvS/i9abcGbtny5zggQay1HR
xXjAWHiprw2xy9NE/70wWpoOANHlorKk+Lh7GUxudTGe+lRLMeSbnNl8aakks2hB
F0QoSFdezR9+UeNLOIBpoQBlTV7il8ZnFEvhFMx/pyTH6AIVHL7wiC0two7HS/tj
p2YZZxyk7iykFU5/HubMVzWv5AVMD5XgNH/ZyeqLDJ7UO4GMOa0RmR6MRJOHlbdr
tWVNJF6wASN0ekyllf5IHdgIZ8g3AVT337ncASm7TJ3WUU4I+hLZgverZf0f/qVD
P7TgPhl15K2LFS6OPLY3UFuovHqi2JMhTPGDD8HOUIECBfGse5Tc6G5GPsjSftOk
EG1vsFtTommajuk2SI0Hd4Rtn/iwzLUKp5LA2TSbh3xOPHpDhiuN0INjmoEAaQab
o0KZk1fOrLdfO1IsAZUoHHbhEaUiUSfd2KltQejVnJkbIqpXZORQJDRn5EbrjQ/U
nqzVHxgmPpYNPkJwzqqjTsC31SYlIJ1elpT09kFzuRnSZ4NuQ/Y7WTyc+ehsy2pA
B8QM7bw/hOKbA69WeGqyfaS+zBGXIWhhNj1m2vsD6/nv1CiPJQBCWf/oD7O5nTxW
uopigODhBZKIjD+M1yVlMK04gxiy1OSv1WUT4hLgyEOBYQ7//QwPnnpvRnv06YW0
9nzk5PsE69nv7OqUcQ3r+jKWSBp5Vzft5C3MkS0k1guEVLiXIxyMs7KyJEaM3vDv
xWakYeCaAAorv0P27AWeB+LElKxNbw04K9ua506GNVYftQRBBJfEklvZdEfoJwuL
a7/nQ6kgi6qHI+S/aHYjkF7xqe9k85wHGpZmV5sx+i1AUiP0DwF7/4rU+oodN8aI
paHJHNJrKXqjKkTzNNcDWwynM/6u1LInVSKtiJCgBZ8RJMUju8zmtmxsb/zwx0yB
pTYYidV3mfkQsMNlqKf6/zgVOWPFw8Q66fCGE6fEGQdKTeOVOWm0aGMWx640gy2a
iLkFJBFtmLyw81+aoW49ajxIbeZRLMCo/WChqSHGoi6meOeM0q+I/aoHbOyMdV8I
gLlZzpgNsl2HD2Vqp+ChlVoSMcfU2feL8cM9H0PgjNcQjEf3YYMJQoffilIoM+Ds
xnNUuozvebxSyftRjFrkdSzpufHY80mHw/v+dwmvHw1KUI8E4zkOGqQB0k+Edm2U
MEcfiyyPNNpBUytrEU19uhn4HEbTitNcaz+hM2Oj8vGwI75xUTr8cj5bSH+PTME3
uFbLI88AJG88CJeNtZ3EvOhNDi4oIZs4UpsPbzfpJY1nckPu4GMH0l3zNuSeSR+N
FNoQwQ5pcGSLe8Dlso400nuzOEmL+ETqXFm8n51UDrlQinJ7mIZaC0flEgzSzgjD
+VUxzUxGJTM/Xp15q+2zn2GFKkejTooQstMScMmUSyOw/f/j+5smsJKpxXOUChBZ
0LLxGfMUNZMP02kbYjOO6Fhve/0WQYwU6zoNe01pc4LD6wEhk/FZWXHgYpNUdxsL
kEDdZJ1uu30ZyHrnomgzWY24TqT2dOLKxESfk3HP6f6+ITGWw2SsaRMiBQHVCpLm
gb1ujZ+vw1xTwCQxbaPSkx8aGzgI4Cj+fucP75VqB65BubAGrKK5QKlSj5LPm26J
bkJts2mn10KMpXewCi4kSl5zCNy/oOcdDIOsQKU+rR/hCSQ7HczGd2PXittG5psh
/I9FYY7ZRgBH3fk296WqE9AoWA12gqyZWqQPiW5aLGKec58Unjj8C4W5LiNWXx13
hbmc4VSlc/mOm5QdgBDHbhoJo4cStdzjY3rJF2txXFn/iegPoH1AyPozqo02pYVl
kpZ0osXWXlgrC5buwE7JBYpdJSCMuwZrsHqG5TftMiMsvPAXLbWGv+JaxLENkTQX
l05ppgdkAiWEgOhzUU/oKWsNzzeQD7UYp2ol8yk+fg4ldSQZ/V+52OSwIfT8bJHM
Jh+kSTmMg3j06+sN7r4mpHVlhbAjUTxOynU3K+Nwqi0/kub6Y5F2rY/Y3BX67f+F
vMLgji0aJtPhjoH4WlWQ0Vqgsph4XQVRw0DbVBqBhUcAwJpkktEcX2vAIATCgs+v
NafV3MN4teuNbAojVbgewclVxOeT6RshkY74NQzM+bXj7GC3pHkOqTmtvHTGw4ns
h5t/GOARe7kHUfKpjxhJCL9LSPjoJPyoI9q7/hquIqj2rVf1UBGAgHhF7Ni35ZPP
7UVvaVm83ejS19quxCO28CxXkZqBtGM4xZxI4Q++hveCGk1Q4KnUNtv2soQsoVF2
xPNIYihrKMbteQG5EhGfRGL7px06BEk3gS8WQCAtyzoihD2aj0KmD7gcZgJH7zid
lHwQXKS2tnoNiagUoEDiwhvqoMujgOoqpLptBbvUh8/D3nJhoI0jIbQsuuQ1adJ2
v0KSdtuMiqJMp6Q+WSW7EM5/cNFfo3OqUOKJLJYRBIKSS/0A6afAVvS3S4Hj9al+
VJo5dmXsqwcchykCocmXAcB8yxtxngYOihMb8LCA8QvoArMYwJFK496OAMNxmIbg
9ktzCJhGmRHymlVn3SJk2AGwtEvkX5jXtjO5XKVu3X1SR7lxRuWSfhrPpoYWQK2d
e/o3JwXzCTDDHqbabUuu7jJtpLST5d03UcOc87mOGk/6aJRsNbip8AYio6+MlIP/
VGnB7y3SlVctBUs7kNICvWrXVE5BUusq4CW7DEp9a8JsAXg3L/Ces6sX5HCQgT52
SgVwuyyypkeMjcXe5l/NrtgY492Hfd/JsYVbTavGgty0uFV9q9ZTVVXthmvq2hvt
Sr+Xt0cxd7goGl8gS7XM0rVAGh2C3F2fBtNRULE8R/DTgC6Tsr0qHvALi3hfiPZv
rBKw+RGl3VxlbXMIX2Fa96aJniLD1KlBQ+LDZdMfOUI4PA67sI6TJ7tKXhnlGihV
FsGKlH1OF0WvMfGWMCgWOJKVN+KSpxzK/lRbWwA8WsP4kmZZXwLR2qlKJX0o+73B
h58Zcdi9sYQZkZgoL8+OO4IwdtXRYbtOhVcsOFz8ZEYv3cMhz+AwHndOch0LAVUP
b7AWKbQrrnK8k4Umh/x+1eZDOUVWZOAJIHvaywvfVIZRXoh1JNMU3Wr/6CSMdBu3
qPxbhHzA+A8h+Jvt3nF962eqJATyqT5BfKhSvkJHOupJcAmFFa5E938lwORjZIoz
KraMSNRWErgA0w/5xvOd2Az31heS2zzAiJY62kR11rQWtIESUPTbZTFNYhBCk81c
uMdxjPA8meggn0HHa9R15n0CGXVRD1OWhHvXIYeBgTSHkzRmjaMMLPEwATfbtf+D
pDMUoYNXhKTZM1cQ5ru1A94ACRlIBJClvArCyXnpQs7CoA8hyqXxJh/UsdVbt0ZW
MITs957e8l5dwkZ3NOJC01hqWeer/eKUmnUkJqCM235v/bSX3aN5rDHYnSy4l3Qg
rzzSe8nJSKUob2uaN9Hvuxdeh/bOkb4w/1cJ+HXWHSzX/+d0Tvleku5abnlzXsjB
sgyuEDNTxVJ8v99MBv3Hq2K61/ZYRAng7ZRNSYNMQqmF0x6/ajYz4iqTuFEeuew8
EIqCeJhToLxo1NvsMBxJ5YIxqbL1FSlgyS4oAau0f4ypogmJITK1YO4uj3M+Ss78
Qge3xP88UE2I2Z2lNpPsLFATbu4Rkjw2mwBagl/QPx0bW2mJRgJRnAqlaYExb6LD
qRDIpYSpM0ldPs8v2O2uqU3u8uEQW9d3SeAtVnSSwrQG3TcttHAiwFQMli42H7Qb
Vc+wMDsxYozxZ6Q8DJ08glXC9m5IUr0aeS+aslfhSkbIyUi1eTke00Fov2Iosajr
eQrWxCx4dapk6ODk/dGyknd98s4EaAYZ1bJn8mgTZlQJP56HyjTiz7UtRnRv1NnR
MdTR/OxPx7nbs3NLFscWxynAc4i6MaSrPKdpW1179TbMdyjNdu/TSRPxA+vm/pXv
rV2+X/2IliMk8CXTYo9lS+8njT7EDUsjJG17tYR5nNMoiCkoOQ9Xv64VvRdI5YUK
Itno7V0SYYEdtJfoGIOOcv5j82hYSjfvpRFGeiHheTDDd2GyUZhH/PL9WjJOSQBn
lHEDfNRSH+ylN7+oKUZU6FM9fPEZ8astozWYCGB6N+vppGqc3FfipmC1TTchkYN+
JksD4XUtJR34WUMJKJgNQ4HbB3rhBCj67/1pOMDivflRctvbeZBahg0nT/a7xjfA
iCG2kI/6pW5PykB+8KgBijfxklHsiTX9fiKINAT177iuHzfgyqOU4qVA1DkRxIAf
+7dRKuPkrme2xSqDjrMl5Qkt7/yp5gU97jbSDu4+EtAnMRc0NFjsIVUTFd6XQbGR
+RVIk4jtJSj+zmpGKQFwHmySWOu3oeA8xGT6eyg8WlOdmdQLrWFoHuXV74tCHyJk
IZ8FozzAA9g23lJhA5/deqguxHZKPBv7+B/d7bgnk2pHFd1cnGBfwfYhabMjSUPQ
QVV5tuAaZC5Wysdj5UMGjXue1xJpiR3cUOuzGip/59T8VSvPDKrrZ9YTgUGphAe2
05cDBmNkE2hYURSkh3PAPTOelfLtYEMdPG65Y+CPnnstm4fvSFXlD/ekwhjQ4Bc+
vK683znCWbUVCtElNkR2gh7LJv04W4COhSul8vK1/BuoAz+MpmfOywOOE55W38zI
m766bR1esfqP8h77+1+KmdS7RFYIro5wJDGj6hanPqy8SyEn0hOGZ9Ezf8oTdVg6
g8Yiesf4SU7H1FvXwB8l7mjz0KZj2sh5IwMLQjgRoTelReQpczcCtkqFHtcU4a8n
mVM89olzKBCzs/jzIkse+Yh9rAs79CoPauhIqUI2sL7QXR3lyG7P9Ikf+jkW2WlL
kp3QlDvX189A/G+XwjGtO0IH4EdsfQsYSf14By0KbQPjyfUeLNuW3mZr90pwJiKa
lxVjbk+PHJNvcYlLi1bQuHGZ112/iikYprGBpQU7UBY=
`pragma protect end_protected
