// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:35:41 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
PHbBC/6l5rKdXLlwrS/abeP1SSLC90sK1eh7PX9xVCHmpO1nQUfOxo1E1IuZGkWR
/X24OJceIgRU5QWvVcf3S/2dhjH2zkCTy4aQBpL/CUdsLWHA+3olvS/tn0kL5lHE
DgU4yTuzZlc6ibbxZSuIiBKSjgo58GGstGNY/zNkj94=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 6336)
RsHWJ7MO+pU7Er6caA7TSqYMhbeaQB6IFE4u0IOwU92JFeD+/PtxCOqiBrCxcKpe
4N3LiT3EOE+0hjX0P35X92wvuudFcrI9TtNCjwGpakSZRZ0aIK7f0tBma2PJmlL8
WtUjvgzXQQ/VKL6F117I2z0XXUCYIk5twVQXDylvwqxlvXUdcNRbDVWKBaUUuN+R
OyQn7/8gMI9etBRzXMkTCiJNJTISz1q4xtuMJaKTB2L8B5zD8NrwiDPGaQkF7Ck5
K0KUJ5MJq1HIcP0ti4S/CsOoaSwX54YoeUzqmW5DPGOqF/rqoqzddTclsrDyIki2
2EeHfx+7RkhLT8qpgjGpCDy0zBjeC99wT6xn/hsQK9QeiitFoP720J6ia6XrnScm
gVR2konZHhjmFMUhS2y2cfgLS3p016NXst8amFQs1922d5HnkvtyHb26vKfjDqv3
wRPGnNGDve3e3LlbM226J5R9exVbTWDWrWqHGUJ8Arar46ioXXvJP9u/imshx90F
vXJj8UV2xOcbAqAaB3zhjE/rsqIfpexhRDTaFecDXP0KZvjeOH5hYsT/EkxelNAy
s8fmBLqs925OZVv5BvWxaFa0o+Wgbojit+2TC+mIjFS/zo9ySg1SoKqmIXacRx+4
T8NyAYrEYY0oR7I0+1NDCrRFiKP5i5IBZWRHieLgppcD5jX4/P9kcL9vblwOlhBB
3cXa9s/8cF9GcVVtwLrsH6bTG4YTOAaHzpgVg7hVq7rchMnYUP49g8u9talKpupO
uRJ6004DuX0ZiO7i55NH66mCJwScR9Ih3vkCxcMgNX08sqTw6oIHoUQaGA0uW8fK
0KjovQxoKBuMiQthtAdYS6TnMcGRkR7qpfvYv3rJ06L6XXyf62HA8+GxCk8SaPta
V06QTBl9LMQmzup7JDgNWY5VDm0RJSTvvoT8rlKxUPMygRUqj7wYnxCWCoV1KNFl
QmnSs88H8gFfwatE9JmIlmHgg8vbR0UXm/0XViDMJd1BM2kP/eCW2R7wQrTJqLbA
+x7fVoUmeVxhvtnqLd2XnyQG8rDrM7TWS6pGHzBbrnCviWD0Da+OutoP0Zk67HJI
hkk1UKG7GfQXB05tB76qGkHeIWGU26ENsSOgGDX+7jCz7I1eYLnrchnmhVQNulig
8LUyVtA574vADt5dfiQed3IVt61w9isEOh69+7gLx1+7I/xjsLiDGn6a17wY4Sbo
UwWTsunWtrxT0NtkMv7VMqNJdaiehJxCD5aPv51B1VCgk0AqQGYgAiM/AhMZ0J2C
8plC7F3YoxrrUGQhfg4KEmFRZwHj5vscf8JX2M7Y0+fOq/Jln1ik7CiVoARpmnZw
1jpp0TBuv79GjkmFBpdcPXDah/HBMk2KhUkAplfnTIrlDaJ6yEgnoMl6PMjty67Z
FoInXCCei5udfdLmi4RV8yf+oFqrS1WSrQhwYkP/E//X3EIzeT/JQO3cxo4iIdDW
xF5/KOoGldekzwnT1dei8sVnNH0w5cGQSEx8Xj3zv7lP87ZmUcJ5i3XRWUYAW9/Y
kNi3NGevyHSefvgLhmhdgtbIWJHp2ZdaHm+tGRLMFBU8Gqpf93Ay33m95/Vh7oH0
RezAF9WTr0o1DdmX9mHRAFgy0ZpVMuXYtCfdjdQNz4jw8JVOloFQFdU3dX7Mhab8
DSdn6qb5GFvy0TvtRsNErwV0qHgX0PpQ81kPpkVgzuA7mr588WcugIWkeD3R/dDw
fWS2INsQ4K67DVrIoE4aoH8ef9PlllvblgHiUqkZwLgWCLQHQjoEhnmz/+AemkuX
ouFCQrCidYol8vI6pNyB7oh1QEeHqux3wHKd2xq8eGmOPvn+0EO0WhIEMUOOO2Np
5RiTjGcdwNF9WyquCJF3BmG2u/g25H6hpoHMOEn6tSZ/MKRMncc6/P7MA3QHuM27
DkBxunUVFZ2U2X8SX5ahPIdDCWzMu34BsoqbEy4aRQBHO2Ngxfw1DlXtYi478J8h
P1JB/s4aGnjhDS83mOL1octPFOgQ9CVu5NplBe2fTK6woMQfBBtKAlcT1u8wYyps
9Sn8cSk4wNj/+xsXeX0egUlsHBZeixtJUtVJvbTAJYSOh/8n36owTykcPrv8Rt7K
KFohFRvvAHS946HCyjfmYx2I4Dy6PRP+St5kr0mxRgCSCtDz0bkeI9zEMuOrinHh
8o5+7CvGavqoz9YgewN6fhv5paHTPQ6p+DOTIIYXUOvAlhmhmwkqpTEM6K8kVLar
SULXkfuvK4dR2+fzztM3m0eNI37F/d8qxxy2qMhLsPxitG62kZ5640k38COYtNOd
7W+pu1XHOf95XKOa+Q1MP7ODTaKM2b7BoMLqa84DOi7CrrQNzxmeBlwiK3Nz1zC4
jPTKEwCrsha7hvNSy21qTzXNfVb0rSH/mIImDHMtRfHTj4lNEgPfp7lBsc/EOCF9
bv7LHjCt8X9DuclZBIuWfRkY/HOmtKibCccbX8Rk/HUhT1dS0TmKriA61u0UWLvh
iCt+mNxS5GjXgMyG5irPcAUGalfV46HvdqZ0OQ7sXD9/lDdD7KKbRifjLM9835JY
67AofExA7NYOi+DzJJCDyolTCHYaK/leJTpycyUUCs2cTpzVE7LwqVj6RgU4BkJ7
Kwtow1jXBjaOQqzYLiufbXDUw6WacujmhyfpNgtzPqoBnx8LuO010sadayrF1it5
5ABJxQ3NFHxY1lOEJUyRSYHHP6JwXMmPrPgfhhWJDQyEK5CAkL5F3U9drCbjR7tV
8CbKOwbsWeKfJD3gxJ2NPZYgnh9mC41BOwC+K2pFl68toBNe6IuIBwICwYZE0sIv
yZmsUkd5403L8cfw4Pf8Ib9tg+lxrc0otnQ3JRTgdrG0knibQCmHcunYXkjffPS0
K5uL4hMY70ne4D/G97mCWDE6H0cgum+K1lisXp3gPrX4qYoZrmGPQYieqW95aL/1
3mgp64HRPHEcTc87dgGgTzlvu1FAigd6jVt4hACU/7bnQy0F5HsDKnZKYZrt9v6f
gLKLgPXRNgX4vLwQk8ycMOlM35gHLAO09bORRpwPoP/uzY99fntCPb61b0O4+OKe
U9uhrv+CTWMiRHZnnGYBGn3HMPl/Z4OfTEYpFGvrSiQRo17KUIFn0BAs4wbSL3d0
N5+8s2cCLLDPF5uEWpOn0Pd/CzdSQIEszXGqY7UjhPnw8OAG3wZVc59tY/zkLSxU
V03Xv17VR5/TEWDyrutUvjPCuO2w9X4ic7umTyGzcwQGi2vv04+ug5/SbNItF7zr
gEjSPJnP8W+c8pzSKDUGG62ue+pmiL1mlNYKjs/3nnq/5Gnzz1eomu94n6NYmQxB
B5SB/MdKUEBd9o3bN5Ji1Byki8BeAdJ9NDL2r479zk035SQF97H/AcO2Wo+sNBgj
pWjKi0iM0JAlPcw2u5rNXTlZWbXkv/zG2XswtLN5rYU1fjDgFl1nctvvOlgrBJCX
+A6r5esqvyKJ12uePVTiDdlGGqaMUeA8NUyy9/HczEk3tWHRdPhm/X+G7grw4xo9
3aTeh93PFv8w5zXU/f3nocpw9XLdBKT+9whNKLv9ffHNaTBLHqmfZZJVNnxDZDO5
SEQkTGQFT/pHswPVaSvf3UxFeTp9XOVul0jBdd25346ZqfNMyS9eBALkegKu54RY
tjFxllNhYCL32YEfoXbsyAVg+yX3j2MxGCYT9Ne1A1yYdfJ+gVk4e2v6ui6DPLl4
hdoKY6dkwrCEYKO30+DjsesARXwiuT8UXIItA7JvebJ9sdKhNbpPR1ZpLEa/CDGd
6jCXjQN4QbGkDsIrtmWJLEgGOuCSnQbMB2j6TqYyN6Scu3EhOFvw5y8Je3jwjHFC
W5wEy9rG0ltz8bGH8qAYpQ2DmRTvFspImDHFTeYjspa177HPQQ36ww2QSN2fxhpl
f4CZbem/Hy2BZpNuDoN2AkvxX9dP8sQ1CgbyanfQAMn8TYpfD3CS2Vyz6U2LycYQ
m5v1RThPbCvnxx1ZacrCG7EMB/bVyHJiN+V15jLCpptoRIq/Z2AGsIpha5WBJsYQ
QSaA45vOrJRUivG2qVdsWvG98YzvRgDi/Fcgg4hXjOsy1uXboun7/BsqxG0WZx3k
MtnjpqGYHfNlo8hukPudzyXRxlnpQ5cDR4ObIGS6JQhBXX2hIZVaC+TmFiAOjmUP
Y5U086yjcQko2iO/aKemthbLoVSY9kDTPK5L7DhP/nOd/fS6xcOxONN5HngOHb8n
D2e4KXandQRB22cuk4emMKuGrCU82pKw1wgcBDcJgQnMk3yVsZ1st8I6TNwno6Tz
FlinqIc9BXA+FpTJD2HdZDTg1x4RURbfMRqkUEeet3RSaLV0j5ocTz77qkroCr8G
imqBCyA1WWalewviIUu7mNVfEU5Cwi/hRfpA6ruJqCEojGbo0TXYiOGjo2X+bVN8
6X5zP1FmJnJYeS3EgDq9+QdFKz9I/SXatx9x6Ep2faCPCwDXSIIAaNp6LoKaaa0u
EbMvme+8CiQK9EMd7k7ucpDWrgnYo/H4hOQN9VWwoUXw/IuMAZOZcWWKbkusktKT
tdmTYAnkyAvtRb6FutWchi01EewsNlmZ6nD6SCmg9Ui5fArMG6MR+KPHUda61Ojz
JS9ocB/EhjJ+dpRA9Gi73YS1lNdPuBIiripNd5wo4LYELVWFWkJVDgu0q/L4aSLf
pcCsTOMgp961A3IC75iX6pAOZYejK6RkUAIUHrqWTSjcqxAE5csE40WDXmGNh8cJ
8EQwHSB4JL039lRnNngBhuJ17T9IgYhnvmm7M0SzXU0zUzT251l/BDgIx9xC1MLi
TNpTGraJrS+MvlmfE+8DJMXzn9pu4h+bzSqzwqSwUS6qgXJQ/5hdFHtYs/bvj9kO
hdbhB1natcqwvvoMP8fD4Nr9oYLr6N00cVnXz10AaklYn7kH3vxbP2UR9HeQLwOo
2/HEcaQN+ARJmD5kUdpbVTMVPjPVcYC/mYqsfL9dpn++hgp52O577SFm32/XJHKB
+witmDb4zV0ZvhVZrGip8/HfeoZZK823xb6lbk9TEIe+RIA2awPEnweJj72DQyQG
b7YaufyMqB1lnkvU1GRYOdo4b00npLrahmkw1fFFvoncJyuyBFe0Kyiz4v2BEFZw
PnZP2zKzUQ3251AXXkJ0AAmYZKgrSVBh2QgpqnNegGWySKl2w03YFUEVcjlXyoHV
YhiOMsocgtLPhkIEOP9FVRUmyQyKi7hCs8VGPpejnsHqEL3bLde+ZupKQL8OfIVm
GqxGWU3rLqzxWUsOlMSPpKgv2cDjmYnUXk/mrA2a2eKOpxMAsQYWj2o4KKlcbxhn
nCYpOTGaGuXJ9pdBzEZoTbDv7tYdJEKZevMJ4EC8CM/y1qnu/h2cJU+hj4pLAKr2
DIM3aS65Cnxi5/MPnT/83VnzMW/NeIesAct6DbEOmg09SMDO766UdTvEEKUaO4MS
3EPSj+3l+eRvXPZ01YpB8dnob27ieULz4XLv/B+/u3Y0NYfYn9YoPROtoHmmtc2S
jyrK6jhL5LSYeTaIfcxQcbhFKRBqiydrLrUv6ef/G2dZfwf622ORz8zpSzVWvJJW
eB7FTay3BagO4wcfgUU9bcGvYwyRfkQKLHp/sFlTbR+AqcZj+fpHcxK1H8a2X69i
b2SY98/NT8OcSZzIVokv3ezBSmd+Qe/9tOkK7fDMsYHHfI7T69RAMgav+xUzLW8y
/2Q2Vd81jc/V0PAo9UYx1xe1hPId6aEU/k7/jEiIRZ/dbp/mbwa6FYmieyV0mYhg
aBwNkoFG0vmO51qK6092aHwpgSUcD039RePYm2So0M1LflusY6MkdCWHwbrQ1ELQ
uo3TivGWSf8apRgZwgt0vR/nG/uIKhXQ4CIKFsZigXVPQPNbBh7f7k+asWm7/9Ja
TseamfUB0PhQvz19I7W5B7vSeHohI79fW+/c786M2Qcq289paWSeG8V9sHLHep6n
N4+fhi/NEcm/hqRdJyji0TQwmwZ4GCeXXvSJO1k2D9mSNd85aAfq2g7vLALO+56D
jPrlAttdaowJM76ELNFbao9bL7pQYJPlYTu2hu4yKoX3I0QkxPrTdiSd09b74j0K
Yn0FvzVHXhqtO7hvk7g8Tf/pF8N9+6vBvnPp24Ikkcx9h9S7QDjp09wYyCPA6d1O
iStX1BFZGo+DF+lGWw4WSq09bJPy3xPnJvMQ4gMiLyweecX977pZqrso5OvUOe13
saOog5fQJPEel5VXGLrxPYvK1/jdrODhXEe1GgH0HF4qq1X61fIpHVVhGdXQqhDT
uGWA4g65SuWyLsJ8Bh53CVKm1cPFBt2og2pyn6ZNKg1D8WIVnrTd4Ibk9r/8fhp2
TrqiIyY/zLoOXI0RF3xEBZSSuBrTOowkiyByDFXZ0+D9I30r9UO1NOaNdUf6OHWM
/1LkNexysDriekNKPOk0KS2uW4AlI6MUhzuDdf+baufLUctYDf8T7r48e+jEfWEY
76qV4aLpoT4WLVnwK6twv1Pad+Wb5qdi5lCephtJMF6SUs+H4AXNPxVeN0LpPC1S
T8OGZ+LtXOpBWz2XguahHV31nd1qaQlbgizHdXcgzoUSI5ZzoDWCKvGQ/aqcE8mo
jTswWfDg/E4ZF60mCk2jPupkFlHEnkUJtrTqCa/nSPYb2qFSSPpPz1pnkAYo0zex
V4hwqMt7HJDonp5rLNYt3znuZXeGEMKT7k+ZvJMCZA1s9tC75aZ+KiCKiy5OmwGT
jrhGiIa7FEbDcWdKHhAcLG0ddMT8tVJUx0CYggOq817RrIFcNGNtpVcZE4kkhtBY
ZOuqyDh3FXYyhwyhxwf0rTg5h8NnhQ7CwCPqhFYmndLXQFXqeD0pyHe2BPUA+jGY
WFpUxHhn5aID5WWoILTF37lX7eVTQiZwSfx5O0mNwubD2zJgsq9ebZZ0scwsG6Bb
tR5O9k+0RFYh3ItzNXCUn4gaMeOMvDE0ZaEs0rpMt4nDrwifRPS062lovsvf+zMe
vHWOddRDh2cFZzF9nf6FwfLtF1oOqAA07ITjverNcGTJOOA1/bVW24ByQM20mmhB
3thN00I+9Z9yL8vig03o15leWdpUfISYsdInnWg+Umvj9PfKldi1gFyWGl7x9cDw
zMriMycgscz8HbM6HPN8/ym3D9eOVdo1DhRyjTQMys7K9ZsDe6d2yuWbAvJZGEiX
bsG50j1VDnky0elogylN4vD0h8P5rTvvkP1nUr3rdjh6n4dpe6+CdSUdx7e8YPTc
c1uWXxQ57wcgruhsmIIfHjOiEqfDJzCwy0Shqo/72D3yw1IWT0nP3UIeXY9+W4QY
dRvsE4dp2JoMHrsH2CiyEGHDrfnE2ACeKpQvzqVM6DilzvWIMlIo+s0l/HiZKQnU
OMgSi+zfGWffouoclFKkaDNqFq4oOtMPZxg/711aNZ8zHHk/O4iww5uCxriHO8ov
2q+wY/D8rJ3z2SEfotfuhAuL0Tqr/y7HhwE9b16fQhgQAjFPYVcFZuVn+rFvz5CE
JN4nKF3JIf1lTgC1KpzS8tZrb2s79Si+I0553a3umC1t3Kt9lkum/8D0i0NtF8Tl
3KgKhT+Mf0jd4IYn+9y+ShCQGV7J3q2lUZj/J7gf727paN64DJ2TjxxDDZEDkvyy
o9TBhV4zp+7xUwmwoepruVwjrbL6IS36q4r+b0UUJZkO61BRW7nx/TjF5Qp4L6jJ
KfbzFxei0PTxCnm0co957rUgCcHM5FHLVnylefmWnxYm2H7X+ATbLpAAvRtZxg5X
hbEFTZAfYPqW+rqzr3BMbmEwaF3RfobWBtcje5GpD4XzyXkj8R6oFfDbO3mnyLY0
veN1Sw+BCImZx3Wv5wJ+3Hrwah1oXhV4r/dqaAFr+YB53nBVoX37XvXZ325xXLTT
b1sXrAox78ky7bghHuj/SPQcUeeH0pBV3TIKEZRGrhtxyk5Ak7gWAAHICZnHXL5c
rhWBJLwMnZy1ddhiNm1TFFDzPvmcWHICXvWQD27pAtZWTYgQ211TfMy5ZEv5QhhR
3YKDKVMllWMZi4Stadmpgt7S9LZ5kApxIluhy3wyNQZvxhp4rUDutJ/4ePuDFkjS
fDnd4m7o/u+4a0GPGppNwUOzNW5YTljDPwSGvSyZKEQ6sWJ5ldiyR2TbKAa1Apmn
JyaDLGFXf4I1aFQNMSRW2IHOzHaR7wIOa1HmSiiDvJVdSTGKDdxAcqyoKCBKsFZd
94bw37fyefXizYXzZUcctREIKly9V946eCQFhQeIGtnDmM9Lq+I2KSqhccetSlhN
BxZPYrzQ4Q7EMJ39YvgQMXi5hqbeXq7AskcGs9tDw6BFQfA0zrPsn5WkdJ0cpWyX
F3NOLatpqbOHXU6wD/HKIjV5bAKq0y5kGRQG0prpyZGFl8Odr0PcVEfME+j4+beK
4QjTJ0xPzwu76R2WP/HkJgPCOBQYaHGBP4BeRaoUsuBheRrFJLtSsC28zR0tVLrV
`pragma protect end_protected
