// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:32 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Rz7+1HiFVSzTRNsEOG/tk9Db5IB3+AI5W7MQbc339cjaZ4ywDU9lbDOkbUpGVm4t
4A3JLkYNeWORSyu7UtOql62jACjuTNTwujewB9tuVqYwGyeCocrSXz+HwEx6664A
v5S6h2zUVqV6G4YP7SLXRKtu5QHaQhrM3CqDVe6jPsk=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 19088)
4kNA2DLRr6vaDbywXluTYz7x7VwqkRbaAIiAYI1BAWqgJIhkeDDlcPVaZkSmks7p
1jqu/VKAYOgJCAQNtnoJdR5wZYBLTy94qi9l5Y19uv6LIAq3dI2Q2vud0G6dQzvm
m0eh1lQ166q1s7i6dpRiiD6rhg5F60ZTsW01E0UFJ9SE0OQ1S9ujWKScjPbDK/1y
XpaRsdCzEDMip7mU80T2mq2LG/VUsxXcrD8DyTkUWrC/1EC0jfS+ZcqVWpZY6WkB
jNJzYCn/ONEmQz2C0eDyVxxM8gWjarXVz97hcBr9FPRHfWlQMN3TjLute8RComKl
RDwGFLK6chbKodzjk/i9TY2cYusIuRh6cv3JbXAcpe+Ag2kDXms1ZiFtrU3z+xPa
tT2D9Ga5TYsUS0lW3RjMKTmvcEAEkzsLTkzVN0Ln0tLnmq5uergpqKZnmMYoUYBq
DTIlgZQwzMe3m0hWZRQF+hadqsPey2zMp71O/8VHwo78HL4Itwo+3aVbx9yUV6wW
LVwg2/7KU3e/KexIMMeo0dqOQz60xa8bCSVxyRzxqyaTKz0PNURquU+Ttw+1TH1y
DTbLl4cAHnn53zLrSg+gRPjY0Vzb/FlSs1jnwaore910XXtIRmQMLCuUMwCUvZ94
Mfpa+3kaq77d9vUoXFKJymWXMv++kN9hHJXQHDN6ZBYOuagWR4hipm8Z9P3B2E1F
1XQgy6yg8p40uMPMsos684wPrnxbxK7FbDcdvW49FxSqFy298iKBL/E5VjZVO4Ay
rP6kbYWO12Sj0QM0TOhimp3aVNoSbahkSPCtLJ0YtpUWF9MJjRVaLYPfYXMW/BRs
7yI+EJ7mI9wBwqCMzAjzDxx+sKjheuAiWPC6QYmcShFMRdUVrQlu8bV5BLe5/cJa
D+qXGUNLzLuQ9DKVzNBI2etunJjWwC9kMbtRAVBrg0XZI1EWD7NpX8WK4AB2j7pi
aSrFrZ7+bj+Zp+DzxQh7FjY5NIh6p12axJNPA+zDJuTcv4SmQr+CdztPpaIg9fgn
oysiGgJzrYo5MaD7+VmA0lpfLOlPDXPbO3nwh8TpswYQOEhKfkDsFm6jMPEa9CHI
kgvtX9hf3rsdb6djonBcIDZXtJL6MHT2mNPB1I8ilZ4BWD/WQq8lOmlIBHg8VXXK
e10wwUZH86sdfhzNsM4ZkYdCq8swBNxoIOkGOKv4hqbqBaR1ro22KbLjEFXZngEn
BdFHe845ZMNwy8787gORSC0c+0XhGvcPl8MCckTsuymFC/5qTrEcT0L/ezt/aRUF
HtBSUfjxhwmszyUGSHxpqUgSwTGGAtE/xGAwEjrcHD0G13UmBou5Xy8av+AA+NoE
Np2oLpcX+DOb8odBHoPYLD8G0s/v6afnkMDE8CKqUDquaL37zGWym0QCu3SbY6io
2F3dzJcrzRgO+I6jW2watfDJFlUwHxtbHY4xeeMQW8G63p3a+ZWn16lzq9LB6mJ0
dXp1/Ce8DndvtlKDiiLqwml9PZqviMNOCdTz0CW/xqSceZC6cZ+T7gJ1i00ewskO
uYqDaON1n7MPVMOKCD1X2YB9cUt22e/aAJDDuDpgt0Zgg6+lB7Q3rGtH/q4ppBbW
sdmG2ae/wLoMh1ySIZ15TUGIpnMIcg4tQFoYrnLrbcCLVV4lI5wSZ+SUhdFXA5mG
89GN9PW7M8Y2ZfUl3SozT514WycM+/OpjJQICfR05ItkPSmfghbStcULg9kut26w
+920D/3KTFHqdRwWD33zBUEbyPjKG/ACqYfHhAtr22c5EFt8H3zqJjvioMd4taEd
NtM1TdmWof97rKeJ9E5HfjvYUnhrzMJZuO4JHHcZi6hYbW1EIK+9X+jyRLmqkjwz
LAJQeHJEp6Uca1ME4jUPZoYkplpkqP40NXmwgseLsa39PaKInG5F36aEqjKMn/1a
MOfG6t4H1JKqnn243vnxc20SoRDNM5gyCGHZUzxHlye8tiw2r3QZBsJCsNSVC9Mv
NWTM9PORhYdjk/F5iXs9eI/99UK6gKwZbjBi8Lbf9Kt53LptgZswZdgLUGEzwGJ5
QODmNFRtgEJYG/J5Xd7lXIM6rn+hl1b/dF4LrR4TQRamhyx5NNWL5yufxLalP8d8
+KT0pMASpUdnfyoGg+H+zbOdfCufN69MIsOI6oGfgDVvL174yZk1sMfBA+DLqveu
RX59qZwbAR3QEZU/MIZBSqrw8/2BboE/y/y95SLjNo9gd9VWsOkoleD3xmDne5T0
uwmuObBbBYmsafVKqlQc1qYpSAYL7NRQkmZn69lds5KZGMzUaZRHEPVqcevgl+TH
gTZ7nhls0/qxSzNuA5uymz1NzGRQdAPJyNdlelrbzEU+TeMK1lp8x3gMvzBy24oI
fbIpfg6PIs0fJuL5Dh+L2Vev1vjr2cljLrZJLsIznfzBJvCJY4E5nw9vG6HuwX4L
pxDwsPCgB1XPrFJVn+K9xCV2uQGIl6+pd/1NZc/pwGCMOGvatDwjF+BNLi/aJa5q
g2Q0hfi7QIBPyrCo1FrQ1O84xcGEEv0K82Wn+6l2pCae/qwvPxeC9GGwmBMXH26l
EpyJ8NF67O+yedXux2ENyvDqMW59Lqp+rYg9Z+T2k5CL+6LHY0h6JzQ3DET93WGX
STAhOKeytvlB7ZfnU1WP8QVZA37uBXoeGhxIVOFxwaH4CABLWofFDZ8RAklB7i9O
WDwyPXv8//c/33fQdiLcyI3or3rXrRrQuErlvH5yrDG0jLigX272KTc6dYu8Iogz
rAXv0Nwz7nAYPptx5P1O94h4s7vNdI39bKUaOx6ZjcM1aW2IcKeUulK+S2K2aBUa
QEVy+8KO5S5QsNsLtUdS5mD1TI1bSr4eOLCEfkyxU/AOdkMU7NUwJOs1ElAGiGwN
ISmzkKNbnwskaMJ/X4GgDOzTndRL5GuAjDyYsckhNRA/mceI4z/rmmvgdaTotDXO
L/ezZ8QilwVvrHSBsGqTB18fAshSeFxKf766VPzG28xQouoBGrQWU04h09h3dWfw
5hx49EtYSkGB9R+OI64y2PSi+wdMF4xFzrMux+GD4kyBvGT2CcxvuaYxxrkmsa6+
rsDgHCMkHlnfg2NNI0IxWK/4yP+Gpt0HfmKQeoQqias9Sf34YaLkkQZHdFBc8urm
Y/ojWWYzdWxf6702pmqJa3sMUu3xl4joGVu+Us2SggnaYZbHhIZaLYcAagXp27im
WTbaQ3X8ScoxE1oYl0rQhTdvxEspc1IHxz06zaTJbDs2W++uQ+ef0Tk0/eQuzvuj
2+F6+/5B9XkLH0oDcI4X77oa4s5fM5ZxNv49VS3wWQb/v+V7R7FOEQ3aPWLVZTY/
eqV5nZdqlYb876y67NXz3q9fikeZw2X+zlu2poC5BzIBqfvWkzsO54tNe8agdVVo
Y6mDfNXIud6pED4Y4//Kh3s7vcbmqJyJzyfG8xH+W08Mf2m7edK/dnf/uQ6I+ySI
ARLpgL7EcjGSRkF+MBTH7Raa13WA4VLrRdDMc1jN9eLOtK8u0M0eD5jSOiF0zuEl
XgrpPbba0QRIGu2SR1tUnD4I6BZOfd5HEfgkf2GrpMzr2/aV/ZalWqeY/nbd9oJ4
/XRALwAkFANaYo7gOwKwRTUMZtiPwvNsXzkPKo8w99EVN+BnTHQjgrSsZMydBQoF
ahsxkpVTnx7h5pQNbunFOtszDijQ2r0vUQOLySXxNYRIMF2SbRYaWMDkGvrwwbfM
aM2DoWmJ1QsuYcaR/UYQ9gpskx+VNAK8bImOJFc5PDQXxPLDqRv/xCfu9JcoMNPb
WqA+vBwmYR33ixkuHMoh7iyvsmC60v406p+grdDMlsHvMlxNEJu0qoyyfPr/SkZi
HKkwNFXyTYsW9s/64SHuUuPXlfLRhL/KVCtvhbAzmmfgW8psQJJJTBVUgNr/+ox/
LdBxWZTw8BnUj5V2ld0NfsLYJwhNDNfSHQcIV/v8QXYPhHqlBvLOf6Zchl/1E6Rw
ylCDosLzbkVuTg4xk2qWnJu8gt+a0XhcCdZlc2M0uKWnSEDpXiBnATdShkvp/klr
q+yeYQ7ZaHzvhgwIThEW0xqr+wGr9FLaVeaQdk4g4zLtJU7GAKjVCTadlQOarY2D
SdFZnswxblhHOHpf4xOpAQ/pmDd09ZWxiS2vQ6/tVp8cEl5xB/cLYVlOGSuOLA/1
oocDP+b4S4Fci/c+PjboCllMjVyRw3QJQ5byF2j+weNh+aXeeNfz+QfHOoHqOE7I
jKRNHOc0St/zLllL/O7SfD2V7nA8f+rGYR0b9/UYsjLN7/2bZhjg/FuO5+xEGuYO
j3nC0ttWJVthYT+i2aon/ZZ0ht0oqRKxZCgy/OmIPKdcWCSzQrP+YccCtcD+uUt+
xvrxFa+FmmtZz5fuigqlNFTrnw9+INHXy5yfQrB9cHPy+6HzASL0mOnpAUAqLpj0
sY5L2VPEoQQYITIXVgoQgUoopSnHSqe59qsKsThUDU63/jgCgEfFFB9n9weSp/+8
v6ENLjk9pDvzwO5UdlDT1D/EvWAy7YGuSa2tupdHrYPRbF/wcD6fxCcAc6Awe9Ke
W6IbOOv07eI3l5alRO77kXhK+UY0Hr03wpnSEUxh49RvSAXFntUjipN4tVYPlhFb
oZaVCOpJlJcvO5IG60F9hW0SeGNoOSnEwfAE8Ib+kpneWLolXRKAkvnoF6etZG6w
bK3n4TlVX/1W+G/5M+okBbjdY6ZWmDWenKECHi4DmUhJS6fFmvm0/h1tjXZca3dc
6GeJIivaOE1+taTtqWQipIA8GnSUxn0KFFxRCnLeLIvdi7HPxiRs5SqAa3kSdOni
wPexSpjpbt7EfzcRrD7RaHXcy6WxtoJWLw0vJNVSTkJ/1U/vo2kOhcHhXzhiCLI1
tVh8Cy98B/OSeqKQHaLXCffspdpYbpGQm6OZxIoeWWilSApNrbJlVf8Z7+l0ztMH
MfBw593LPoA8fWoSCv4aHqDS2RiZrDENR6MKCaY7lPvh2s5zR9Wz9MkQTPYzuWS6
2/e8TXxKtP10WRGoXkz6l9qn3dS2oG3krRBSRDKHEMwOm8G9SJtRmT0EmIl2/BAV
1dw7ed3q7wUOBA7U6a5ZKUPziQqJ+pHoirRiJa3j9P4cg7qF0Qps100sQyLhgDdW
ROWfHcT+X04szs8ibs76ija9BpfWSM5rxuP6rZuwlIytJkhb+iAvS8gO0L+tFgTn
6EEd86g5OBsksrebL6Lz0tKdD0eRvBwcd/Hx6tN4rlqpl0vAw9yzNtp1fra045MR
LSD8sZUQUWMo50CPkuStVQwyAzyBoeMPlspMj5FsJYmOBg9cQpcSLoD3ElCWKH6s
N9gPAa+rV9pIQBZg2OxJqw7IgpXUPQycG5tyW8/PTYE+jhlB+TD1iHw0yNNidbIT
Eg4zT1GszSPS7kE0CFeAwaqDanutlNtzU42Vv8PPa8x1BRgTq+hyOUEjh+uXDJb5
27+gqvIkEPm0dPAr8cbP8Tnztcci3l/fVtsyTTPrLRVNeUZAx7SgXROpVdy0lNNG
4rUarMfhSMrSYzgdiokBinWHfMYfg8LPU3ad6KF8fGHZaJbJu/wltFYIm8TqVPaA
w2hHEZZIFaGofIHsFevl4Ml3trgptG4Yd8uIPTh7hpIoOtZWYwHbRCJKWqmCJ4qP
KJC6C1RfvApeLO2v7j/ln1bveHYyU1gTvlxaXQ/UEelVuvL+KO8IsPNcjEeDajo7
azjVO3yjTV82to4XKyfPpfMGuzcxRAx6wCz822edR1ysAUXTa3N0KiXCL/aUREqh
Fw/dB+nE9J0EgccXfy5Yng8jFnsM+gjyS9BV9ldb/F9c0EpTlgOADS/369lVCONk
ApiUtnUxLaai1aRiXmPUwamzkzZbAGQ8IRgkLlNbxdQ69jbFIotCornnJcjx1TxW
hOXE4dlcQaYduIZ3CzgaLlGN9P1a8Elft670MP4stCm2EWq53UqE1wEamaOjytfO
KgdbHNejOocKENaOsa3cDHZ9U+C3iQBY3R2G4d5qKe1URjXNnTzv2qnoNnCLoaga
vbBDFlH9EG5oG+obdEu5i7/yS4eupBoDb4+MYj/1NZCRLppY8t7X1gTjNaLRBp4Y
eBkCp3JlbupLBAak6GFJ3y4DqnTKix2MgnPeCp/pfFOrUI/3B1c3iqOlbKBKIm+K
uOOCvCUCH632NDaXKcLXEIZ7vjIXr1vSoxhkuMTO/PIQCqVPZhSWwyy/MxwPAJee
lPIocVm4teqv3O3S5eqhsVkOX3R8UkrHYPHVwep8gZ0MzKAC0dgXlda9FnnMvilM
N7k4m0Es+foMpJWwkJ+xmJVrCSAb9raEw4qTKE9EgJRfggt0Esn2o9ZYc0imsluv
Ec7/y17zK/cTAg3h4Sn18gg8+kV3cGm3Kql7X5zDS1sXQbjz/AaKf59097xs/Mbk
7ewgYUPAI6/8ljRnYfI7hqA6aGVOupaPEC9IDk/lwXYnEtByWqKrhRUldx+om2XT
2Fk1aWj8QTeGQeIIgT6pD8fsGKrSvZEXRCJ/x3Ljn+jQZa9GRcRhJBkWTZ8ucNeE
Z75JMssodKOKs3LnGELR2YX7pjDgkIISDSbEbwVbrmnzI0taaszlQAutICRMGSXB
wbdINI5sDOP7xLA0vSe9tWRzWrg7qpvmp80vbaysjA+gLEGDsT+Rp2QmX/EcQzsA
nSyv5+E0/m3VzirmuYEaCWzj+t5KL8dWZl9PEvhmZkhc7PuTDSWvCoxly9nlRFYQ
R0x5KB7IIRnjbxxxjDY/I+V8yVEzEl/PNw2yxknO2FkeM3wK/qXHvKzuiN+h8KTR
cYNaCsDzHrVza+BxrFIrT1iSkEa+2Q5NTYGgaQpZsnLTN1ODd4buDTWCqs5bYgx4
sY9JMsXdRZSYa26P7XmIDLd5Ck+vrYcEUM/sr8OkdQfBjHcGB7hmXUylkhAzub+U
SVjjEsXhyqDsYfsL4brjIWwpY+eYrIDgEIL2wuf12nDPDFdoPF9Y6+plaWCqDrZe
WlxkZOMvU9QZctkJoCMQhD+8qLsRiGaZkwP9LAEs7hszzOXKYJnSeQV3SB09LxPT
yoh5ENUqfPh51CgIOvn0dMWVVTRTz0oLovG9zsYuEa5weZo/tIDheY7qJxpwMl5N
fK2HF6es2sbrWnSTZTglr9c8Yyf8iqlG7AKsBYf+R3Jt57LiYgbBII2KPR3SHKhO
fQEJALl/IVkD8/Dq838A1Q1jUKHmhW1UkEdrEZIvCw53mEh86wn+EFHBZjU0Cr3m
unu8t9ap1NMO+QiGr0M5dCds6BfwTE5fjrykqGw9J4So60sYqdTigq62dzLbAlUN
3uNNx7V8PPXW3qKEhquQzx9oWu5FOCF1KJzgsAmHPFpwi4eiH9jgGYVWNRqgq+W/
duTN4oLacxz5aHUENNsi5jzSXfV7QLJiyvKdIHFLX3Cu3mp3EHMCcJfVCVcy8PkS
CM2OoLPL1g6W4sUr3gp6Jh5iBpGki7m1YQ4g4wwBj3bxQu+HOlctFigNr7EYhIfZ
4AC1ESZa61Jh2OCYtri2rbwda7w8UHQpwprvmX/s9Ra/kwtUHgsngkGggHcfQ0/a
AD7cL2Qn4MaorL9lyhQQzDxfTo5jZL8RcT5+TaPQZcnD/98w8qoa7W1KwB+TfhTG
Zwlgqhikj8ruOpV1U23pFa88bKP4mPUevNrqPrQh9map7k6fxZYS8crxz3A7Gpu1
/XGF6q4yakALKebb8qpm+kyP9Rwxn6GCWImwXW4DZYTldsaVCc/AgZtVA5+C5Fgf
eAfzxNakE2ePuslxL/z28EUspWvY3kQS9A+qsh8fpR9tCenSqIS8KbPO84ZlN9DT
mMcz2BFCIM43oqTPKHscH8xnPovi9YsDJYZL8kkTc3jHT8sQxGxd7UMJdW6ubytT
/mWGg1YOOig+zKj+vXnxBRGzWBrMjOF9cHDJR62jMbb08TMoODdYhzSL5NoagfFi
0+cAA0u2hW4kV8m0PaYnuR/bEjbqczZmycUIXvrPfoFoKYsQWBmFo4N4IjCw+cnB
RL9I5kXKW27llbdd5kfx5mqxXogCGj68cbkwsOccCLtr191L72lUO+DSbfpvMxhx
Pd7ArUgTjWNhcOuf7UJqlZx2Z9q2dOMGaxi6jI8cLRkAcBq8s1HeBqFcEr2T2r+x
LVc7swruR2QJhk4ZizLC10kH7rhzl/vRN6TuIkoiYPGTx3kZz/vKOuGpHqM2GBF0
1qq7bXLRjYureX2AoBE6X9X4SbQnINb9HvO262NUkssWhkD3OJpv9TG7dHct/hxc
txv6rWcXiYMNcJ4KvCUa7rpYr/ViCnTIqTfWREGkFCBIYTQDtirf44UIu5CWAxAw
JYnkvusBE+KUUlKvWU/EL1qAeMgzMlRe17pkVYR6y7Cbx+ZozduKrwVQ50On2cQM
IUAXFFGWjgtJldD30WNeef4iffCSeiGGjIFvvxJesFXPjBF2Y+IQBiLLKP8EGkIt
NsrwbIMN33oTnf/A1TVRSt65FmW2UE7VcO31D/VWI6mF9Vat0mwKuMUNkooG1Smu
jAMglVnjP4lkrK4AJFY+kYb1QSqYtjFezvPCXc+E3RHphYxE7cwK4IbV0vLOnUaK
4ob/dMtAamCVCgoUXGZp5r878aO/QMiIFY5L1HkjWFM62vqs8Jow1pNO4OK2WRbr
oIIHoTlzuE3fi5VsDT6ZFgfMEWkSQWJ/pbcHEGm+8asGzQ7AYKWRBfbThN7eBKi9
5zTRq/8Wo6lruK4+TIcG28KUxK/2+kLaEM5SG1QrmCX09jDb0XpiKGmbTbyY9PVd
/ZmKti5bPiCRIpWxOiJiO2BYOuMICoQvlAVQVMdqROvLWmTg1pAfAv9EDkm0rSMi
+JP6wwiMwVB+O91cPK4Y1UJSwZ02U4jtxx1o+tK3ln15Fk9n6QYl7qpaNqS05KLy
eMdu1iQj4x5TAYE2s2dMbYVdiPWH3G8GZrPG7sdu3zsJjwZUfF4AwCRYS+QI6OZT
uz3XZS0NamVM7Rco5VTKPlp3tym1sYsIeNus7yxB4XvUo+9ygY6T6tPC/mDQAwwS
ECsvkM2iduOHmEGt/rJCCqq+KCD0DczZRJU9zUanf7q38C4095WzJc3/lOyy/b1d
WnVTKMIgg22BSTVAnM+d38k7IUaqdttjEGuWQhYt+ySe9N5Ba/lfjDxjKhLlenNK
l9iCqYK5PWPOvnYtGNA5TEz/Kvx4bNXhaqCopN2QJH/j0Itxqz9/u9st4Gk/UYyZ
XQhZoZp2D1Efv3b0YqaDf+DIkWD7fGP0FvHSVIhISs9ae8fUUriK1nz8Y2ixuIFA
1fqcYNx4eINjIqQivz7pq3Oj5F88zMYkG/baQp6cAQw40EYDUpd7yTKgTz6ZFMsA
rPN0lWI3o+Z37BGvQl/HqkBjtyzGIMHBCWHP9Av7YuZickZszEY9HXYUsgfKwP8z
vy46/6jkWKbeSBvMVhWWTak16kzFY+fdfluno6g+pqkSUQeSuf0XCbQYjXAcV8CI
zzozdTEBpynbnI8vH37Qmz7UAlEkErzF1BdLhzyALhPfSb3SxkfjTYiGyt15v4tN
X3mTBRX8kUDRjUtP30SjUdAUWg7UezKSyYFauj7SxfcubPocCFDuYwYJPFkUuN9K
Y7QEypHLbxPiXMwXWsoD7uwatZifpMmPR1E+6I1fO2VCSTBdmP7y3YAgukgRCupu
oCotGkKAPeJywajVMejxu5C/i+A+ydEU9lIR/ozaQhLzPCKK5oSEyaymoTO2Gk80
0+iEM4sBaDeNyQSzzVGQxygd+bBzPPe0usUtiGB1otJ0U1DHcLJtT1JCzcJ6ZzWw
T5uzsjlyScNySt6uL+9S7Z0ygZXfVhdb5NANC/zIReI+hQYvZPq6jyu8KwuvQFNC
Z1ZEg+aG60gxeaTg8/09MzK6sHOuhXpT48XjTLqF77mAHv9V9ygbi6dYxxcF6092
c1ztSFxnoU7fNZ0JM3+yPMvwejDpXoviBqjXbsaY5nvLkq+EtXwXpxhsL7mfI7yq
lBX9p9DqF/RrMp7CTma0c3on+bQ2pX9c49zvyujMEnMwD6ox+oSMu/o88ai7+Qko
3/wH1Ti0xJjK8w0YlABD03uGc+rLxsWtHJm4Y8IfF5k4rxZXBe5nlFrqOUDjXP7f
trE+BM+uAz2srJLcASHuWu4aO/xVG/lX8itcqB3ciDI16pQK4m1tE8PhrpI9FpMN
oEpozFfjrrF+6yeSgqOJvIFVDH8fMkJ0wyk1XjWnF34sXnSmWwCs9T2U4XTXIyvX
QwFUKP3xKrajC36RX2B6Diho+kvbn5ZzIKjTHnGFSc8uPwpDt2Qx2YCaH0Vjyxrx
B9sZALy2S4+rcTnaUJOml0A/+C8Ae4KpsQVNjYxzMbXdQX6qAOidpviHtW6qH3eZ
pPDgqoIEpQq8Pi524R6Nuv3KOIvT3Xg+Pl1dZdpU/EMTUSd4b4n3nm7OO86/DM6s
xuBcyPCQWSYnmOyUjhlUPAsuFkiDHjS2MkbK87ndOUQho8EKhuw4yJMwEFye4Sc7
7UHkRj0cXMafHbEXHHZ3u+VFpG6nnotGRPsYOqo1k21KVTYuiOboHPNPiPJAlHph
5FyO55R5iNXeOQg1aCSzSHWFwDyw7Qm6JoS2/cqJzNOzyH3WrzeLPLk80nSftXXZ
I4Cr5eTGOgaJRMenoOvbqRunIDiKayDo1VBgvjqYgYGawG0bTyPRVq+5rCy/z7qf
ovwkDeZXeFcOzo4ODvDuj9lHFrgmtcWrRUzy6wytBVZQeLAIlp7gCoth9OAoL7Oa
h4lNu+ozFsObJobjbns/8lDYMzjuFmDWA1SLZA+HyGWwKRSI79Fd93bMSwFK4104
XCz58Zxa5sWNYKFNBGaTG/fmA15ZHfHTxTbymGBHsFSThuYBnbQirnEit/OzePHg
OoMv1cbr52hXTcCb8RS3S+axrT4ZmmR65Tp1mVR7Wkkj7A4vFUkUTjR6meMOrmhV
L2nZLr9vxikMgvv/RuLkYbxGkYxIjCPui4RxIVqtSASjSXBIB5VGniC8hQPiMMKs
lt5aqxOzmikTgMwrtWWTQnCWybmq+So43Er5rwyDcayFWv1jkI5MlE9yxg9sa6bZ
N+PYwx31j5s7oWhNyuWHRgYnh/MkFkjngI8vP+OKIHre/34FdlP2m+RcvLK3cEXE
ljzZ+ntyzNs5jU29LXDMRoH2/aXt1mBpjzrc6shXiCpjYk5G9CKi+jCY5Gqzyznb
RaGZvWb+9etqwaUrfggnnA0c7K0qVMIh027K4EErARNradZV4jJ66mPs5S3MSApG
O1LRSC1OSkWGVgvaGcfSG7nepSbX12+RtUtXhN9vd5j6X8jaAIIVcGjJ0E+X04+n
YMz345oxm0UEb0R0R2aj3R2QFFavpl1a/ueouDhw/mw4FEc41XPUrqk6YeJYkTm+
gA/CZPhmUJnTe0RnyewYtK4YgFSLqTOL+5ehVAWZknTk3IZBS9Q/f/fWnQa4zhae
bFK0rQvFWJ72/tAzbkIpUCJeCJxnGt2GOA4bC3D4CwDpQJKjfExcyXbH7wTH80Gx
87G1B6R7/WTFq6uCEDQ1P/hE2JQH9EmumfXLWNsmUW9k9zUi0eQGP6PmLy4y4xUy
N+gV4xTC/y0h7p2UeaZnH2gV8/NbNAv/OXe2yk9iUPlofSyqCGrWlC6drdEUb3Kx
oNfQijuieZKfNBR1csSdohiBQ4N429oIkRz7bMPp3yAg/ubXRRKNQMrSTn1WEPxJ
IXr51kTkoMUUhvhplHI7QrxsGaMpQYSI6qir+hRj/X7SQpuvuPfKW0J5I/DvmBPN
Y6Y4OF225GK1SoiH/nIZyLcp/LIHeQdlLUGodLiR/0tuu3D2FCBuMmPHREih4MED
4AgJ4QGyU+nvOo3HDap5Ek5XCOahW1BHnZp/1pgDaF3QiXthyn8GVDJqpsFhwzID
wOlNFfJhhFdGigXPvo48oc+q1pXCeCf9Q37vIrgQgAV9Qz5WoQ/Vk22V3j2ZMvIo
jSUDz8Q6wGGqtWUU4u9pOW/O7eY19ng3uUCnh96VmRHfcIf3UxQRkHrOpnjWvFOL
5lJwo3CctsToxOB0GB7WIo1Su0GunNEYGKqWpU3/0WTtqhzw0qwIUj5PsXsbb1Nk
78mKmv2jv8iRHjLHxffXrquDpd5TZaurGyHgmZROz62linRn+NRAEptttoFYZHqN
GSe/7SO0FdmEwuSZL02zsm0wADXFPpgY0vQCgw0AhWmzrYbLqhBXYlPGNHV1Dw7Q
FxOqmKtz9d/C7eM9ENIK2meaCuNKRGqaoOdV+Mc6WlXaWG4MM21cSWjaPn9qkeFO
rgukA7SSqqVlMwKYzqF8Ys6hZk34UPWU3aIHVN/1GCJ6R0X/hhO4fEDdam84r+NJ
/ifm8h/qMxxk3LWjx60nnzm6T477iei25eK+BT9SNGPJlxc9WoNq3HoOhSYjQCFA
5y/Nw96UHUW/pwsfv0qOJdxD5FGsLR9jVttHZ4z2R1kTFuki0mPTvVhmZG6I6pbC
lyIHdYcZbxWtZtI+eqmIG+EF1jSLAw0fVjolCMZhczfeQPHcmRvYhuG91BUeNw/3
xnqAUbvYQprSM7etGFmoRH17CmQobmPCKBJSO8Lr7F6peLeGxlL1Ue5yWR/PKNQQ
NYNLUJYUmqNWkpGD0GnCPd0ujO4KG2GgYjVHJMM9/90hi95Uoly+JhiooRR1YhhO
fiURFcKWj3Rj7h7BBWK5hkzRxgneZt2fN/jMRrXak+SBcRDZgb1KpW3TIOPOJQZS
lp82Qw4pBGdC7KYQcppTKK/6g/WlFmI1Ih0Q4aTsRRIXi9xWhv4YkQmgyN4E/aaM
MwQxNaKgh+uiI3iMfS1zJGkhTo4xMuHSHr8RDeK58hOABKxuj0BWjcQSfkZIlEPh
BCJzQmvI6XCRG/cevXndtHisLyKlBpYAkqrO/94BMNLlTzuBgr5zYqLTDjn+i9Ff
cr8WF8qvv7NvlIx1EMExMY12MGJHFQXPbMZWSetXMLYY8UNaeQ24jwlzZOja/JWj
hXgtnweVCbO75MkbbS7ETsyuC9TMg+rzhIn4PDLW8K3ysHCLid2MTAtS1pmscP23
4PbMmXh9GLjO0bPF4kBb2v6ZA9bt+ytd5FYAT+5efRb+wM7jM0B2zMkJCLvkDkIV
ETXkyQU7ha65o5r1MXQZ1bT1RUqy4gVvZqRye8jBcOIxWG7/FUzc4c1Cn4k2dqyq
RocQaTJyCdsRZAvNol8+QUwRUJnVRsvBNbqC0KXTqbax1iQf79LCnb9LW6glCkPJ
562ZQAXdGTQPNfcoPWgpgghsuUDp771H7cVHWh8KjOBL2L8g/T/jwkri+pWHQdqa
UusjKV6NUbqJBIVZEaZF/Q0On41FrXwD8a5JTwNdZDyRDZq9+c4eLzcc+pLm/WW3
LhcQh7rHe3vcDRKNOMxuaCHtFh0FHF1icGpsYJaEf9B91FbeUUOJxzylcCIEr7lb
FwiWeycRcBzo1eDbqreRYpcTQqqkP6BgCAADLjPPqf4G18FS+I/u5tGcMjQbexlf
7dgLXap9uYG1MX+Jeo4CHD/ZQeg1SZjsFdItw0A87UxjZRdUSVvzfb3vOWzxWkwl
aVZ2pcHF9IPhIWKwjB+9cqNrC3T856AvanoopBYZcZSQ0zIQe9PVBjI9JCgES2gr
BpRg0cOnB3l8/5m+GWuDL8ixaV5DhNH4nrAcyqUPzjupkJLIaAd5O11DhRHVwIEH
+7qrxlMTGpxfMz6gnJKPChlmmHjpgCp5KR4ZWzLqj3VMyBK+7W/THRMzrREW2E+U
86dLw0LNWl70TVMhJp3eqXmckYbL/1jzQuuOGPPa/uS6OJNlsGtxHge95yBPQX3O
7WpNuOJ8i+BkR54lEwgwjQEj4rpRthmxuT7o7qOOR35eg08cYcb+WV/I98MTcQvs
hMQsSc9kmfl96z75deQ351NXjLeuhr7grrtw28G7IpVc1Cv2jueOnkIpwDNW819B
iPLkzVGiN08HqSC4GeNjplP+SXAZ3ZLctsIS/ExWU6MG9uRODUtjAGSyMuiWXXzt
eNDAAutb2PuKtvOq1M50YrZG0kcFli+/4ofQg3HOFT4Xz7KAyGxmOUU4EqoCcVPJ
08RIvBUmkDNKFY9g2xzFc4iKN7uPMWa+9G1/RLwumSmT2vsHgsxTRxLvjYrnI94c
TCSNj6osrqYg5uQrC3NJqfW2shxIRXa53GDRTKDc1NaDzCY06b6sUNDZXEXJcI02
tgfsR1YYk0oO1FGHfoi2kijSC+LGqKjaJdqviSnF0GHW9opoYNGyv7g7Ld5WWIzR
aL39z6MdfZAbTmVyIWccI5Cl9QqX0SYxe65SvgzZz6NXVrESWW4kto4vcjLx1Qu/
kjjqSmcRV+j966YiPIVhV4oOh7Kx0vWLGVFAYvbN7H2Rah+GrdjcMnmyDF5aR7Mw
94nkqaGmj6nL8p34h2F702nBs8c/4o/qS7plVJWsRKtSJhnQcKy9wxDuQWnkn5EP
I9fv9yI8G4mhws3EPJQeehpXXKj4pkNxAHvemcAhlGUPXrVHd4Py3R7BjjMU1oq1
mnxb9nsrcdZr1EIMkxr6q+AfZzvw3zzMx2h8vrN0pRdqwPl7AZXskX6nOCjzkRjM
PmNjOVMZn9pGuGMUOr/5y3HIEBusJw7GPeWRhqA36NT1qtrVXhXcneGSPeRHTtF2
4NE8dNd2HfGO2lV00Qvg1OnuAd4dZN1sy51xGr0VwVYrRPy/7ecu0PdAI8NCRkTK
klBYxI6JKpDbtPIKe1XBpF3fTT4bPelS7zZX4ixUuKS5L9kiT6oUt0IDwrl+qvuq
3xHIly+xaUidBNYns4POxE7bBkH33Xy4VIjaEVfQNRaN5mFtyEcObId3ZjnYJ2XA
KN0xwyfrtUg8fPHljMRP3/xcdcpW8IbDEjhXILrwr+E8YquAreoWChqrmMLkupnv
G3+zaqJTfAQPMZgPjF1baCN6QfbKJYsrwwEQTIkI//e1PilOTomHYoH1IxhQYwvB
wm9dzDb3meql7ndRKh6jwauHRRN0xVDJclHOTFQdgneEpa+/8x94YDwgf+lTTDoG
4UcTT/3JRkzRjc9m1rEVjgkhB/XdRQgvfQFqxFmrWm+wzcu3808yJPHfqcMiZb7n
3OUmEmarYzcr82XuXJNyvOizKSN155Z6Rto9vumACFRwCxVj0lRC82j3ML/W8jou
3Hohz9ktObz2N/2ts0nxTHLJpFPoGATfJM6jdplmBenY5tq3uJ54q/piI/9gQx7v
Z6ksoVsfmQoMMU4crwKyPN49TLHNMCcB/jnrXj1mI0CteR95c7J7E9lDtkOrrDax
kzqzHtLTmZqDrxr7T+jD8pNqXULI97y0aWNSdCT0g5TxRzc9vBPfSpRNXCP8aQtX
wv5yFC6g+m11vUo0Oe1ccdazfYn7c1ORuUDzkqWmlZA/7wYDGn28S5JxAzDKG2Fy
tFvL3+ni/AujWwUFeTKtGNjmfRMqq8rjFyxLZ8Be3qFDM2sD6acn55ViwO4BWddL
O3Tiuqpm6ReqsT5DXYnAVZ7PcBNny+XMz2Q1vvWy1jtB3G7QVndZq09/PbWFZWt5
V/Gzkm+p2mxtVBEnPlKiRz/82+inwvz+fSfgTB1ctlvjdijVBYs9jOzIWXsufvqO
+KqWaTBy2WWSeLOP51Ggao0uGabDRaEUM8Zj/7XWqN4SoaDPtP+rVGf/7+7//PWW
GTq5FyjhoxB4JobFtNGSir/4flg0c60JUQ/HQGP/GFtI/mVowG//iBogxZx2kmQZ
AcOUwB9PZux0dOqVBPbqc42rDxAtvZ9clDR22DxjWCecCqu2PFN9xdrm4M0oZlMH
nvQKsxKrrIMa9uW52sT98WFaeuwN14BT8ISeObXBxtJnYK/AYaoCbLci82Q49CMS
Hso4nZK5KUryNHsU35NJX4m0vg4da7IFtLYY1XLne/IyovLOfWPApTjUJutBSU4H
O3A2JB+FZbK0L314kk71BuwLB3EgD2JeZ8QFpQBQPfKnDtkQxJhGrx4l2LOOouzC
n7UGWoh/6V9YFYfQuo0lIH5/lhHpXI2q+gsgBApmM/G3M0fzJ5jaWwg1cfWzIq3i
c9qx3JbV895aX3RQf3nj3rnE6mZ3saXfGoI1SzmKBT6MwvUG/5LjlJWfmhrI00Ee
EQlaEd+Em32vLKkx9D604tHBjDHXW3jUdn9p3kGlN0MxuHQ//Dn8kJgX3p2dxyDy
kyokj8/zSMjKun9GfCuVfqeUmv6jRSLnfwXAeUQAEy1W1lNT2cZaISpWVCpA53Ff
ScMGsAUPCmBWH20sOh4gf0RJc5+EaXoDj9QrZf5FE63fuCAs05E9+WJ+r7QMk+wn
SIB00OFOX5yPq5RRW1DVALwcWL3ADFUe9/hxi2+K7QFd+jU6qJ99eLQ35eNipWCd
gMaSVIAszBfF74LUoOPPMp6DQoZgDIxjNzoppCxSQSWBmo+Ytm80RHc4a7VnBsWD
Ey3aEfWhRo+ihgiC1iPQLODgOrhssTlMXnvhzYmQXuaEHvpHz0Lkl7ok37mFEIHD
4pOk/MIhcbz5taUy2nahFScMp6uJb8+w+ri5bbyLCEq03Y98tG/PWFQrM9jEHvpI
u0roRD1ofQuYTOGqXvsPnmcy4T5H4SnRHS0WjnbkFh82MrwQB7E/braSXuNbd/il
AMO0qBrqBbwEPq2tzfgZheDhZDY/sVBV8j6EGlwCwo+64p5Pa0SoH8Q6j+wViOmT
A4Thn92Qo11OdjuOVD7HgTzDYXPhiyXemxSPRFFAxUWGXuRzw4snA08AIT5tCrd1
HWg+HYTPvmaoj7FK82kMRkOh/gHPpLJvkDeG3bFs0mJ6HZfh+JLZiht5C44UIKW1
wNFZKqPcEBHCfHrMhhDFE5kBr937PszVdtGLEXuvPsdiv3NRG0Vrrr/g7mycATdr
F6CGqb2ns3jBby+bFfmH/JR+6h2YIRgXKK7i545Phyc1fAnGJEJ2dP5/+Y5UmftV
C/Nl6Ywlzc5skzbc84YYDtonb/hgpMEpAoD42bg9mr6KSgEBQja8QZU9KUXgl4S9
NDd9DMRAfO5eFlZtuyzaxjFZzcB71wcJMYntJq8yqvoKmnKEkPRGwXjYVivhrjRK
WfhnrMwDm7YpR/hDX1SXbttA7CX2r/I5X5o3LJfNMFwD8ABh+5JcCcWtrtGaErVk
+2rWSDpIJlAP/X0z5uzgdVeOcuJJ6pDM56NMZwfvFMsY4R14DH+KYzaE71WZJQV6
nnUhJ4HTl0lZnBpoNUKhIwyyQdkRWhAgldjCm9Px0tgAYALzQs6sU9liyfr8zv3R
+4b3+eEbyjlPpczD5wK9eqBni83HtXjbVAcWmuOaPO2HUtbETNZiOM9X3FASEUA+
uKW+L0N/rOgSoiYbkTlMNImDq2xLfgKHvVbo3Ev8eM38h5cbuSAsIfzCUBZZQejd
l9oIwUhiMW5RgWiLaWc6ePCMHQzgcA53dnWqHgkYDoK9K9YYEenDjRyfhO9EL6G9
5J8qG8pJqiOMI0pfJKbWO4L1ovuYlaVxAnwEuVI9v0IbOHxdc1Lg2ToUz4XbT1+y
+ch5pvejfGn75081BgRDfj1wlq4AgLpzrPbrnbyBP8fUWjF4BJx7QBYlI7wyAWej
XnvZ5soWgk7B15GJPUeOlqo1gBekoKCYkHTG4l9tMchQ9wlFFsOjax5wllvDttZp
z3u4ZK3s4a79hyU5kcmjADZmycRE/eBAlUXmgIBeE0u9jy3o/EFlrwFyI8xlxMqK
ERvAXecwx/6ey/4zXXS2t3D162NqxDtiwCgTmZ42dor9Ui9/ht7R8jVm0my9Au16
+C8BLOV49/q0pPxZmhjTcwXDJEKpUypqJlMJn0GZgadO90bP5zU3QImH/qtoXp6D
KF8cxML2mPx8dqGSB6S9UbEQ7g7AdG8d35ieTZlkxZwl19SwtG/3FZoPztE+y4Z1
ywo/FAnTgB30bb8IwNSv4b5mqo2UTINMqTwyIrPoFMts8G0zf1wLZbXrGoOaluw/
s9H9iGQLwWcSUQYnOLCWaIok+2kE5+4ucSWevpqQnb0SNWMutnSfEcAD0o67lJOg
UT+g9HwUIwylF3pSEqDGcxEGdvuj8IhYNHtaaPFyl53kQwv1wDTOqndNZ0oHz9F5
GMNexiHR3dB3yTIv8YsdMoHCAWhFcNV+QaFpfWpFACkajfdFSOWImjwZr4cDM1Dt
fvM6rkRpaB+VmmEGqYG4zJvndNTabgRDzW2am6R6mp7MlsJXKKSopJkV54RZtsOv
ohuh0is1dGLq7/HJFQEggAwsxSpsNjLTWvB0r24Th0e5MRgSvHraC18GFA2z/o8Q
IUNbokRnFPDBWdbFKl8i/kmQb/UzLbn2JwMqPQfoiPRXDyvuFvBf1kH1ILDpSDjf
w/dZMwB+MsPsT5ocGflUp13+h3wi1CGALlvyX3NU2iM0Hj7O2rbOGKw52XCZQJkE
p+4YYgBkV7L+Z0KqJuZFEI0lodByChGzZXc7mz9w+7NFxdxmNkYY+tzAAZkl3CB0
DNCCs0XIicT7uxojWn+Rn4XRmeuk6mI9fzf60yiWtbb9t8AmlZwgsbmX4d933jXs
SBn77biALDBlzm9D+LTbDWqJ6QLQaZQwHNRPx1/WpgDuehpFRB8t2kGSC+yA1BNv
QPGadT0Y/Gc0VluQau01xFXhpzkc7j3ZmqxsO88hL+50/6OaCvP9Iz3fHB1Eod/d
ql0aFh9GzDxQGn+2yzMDEnon96Zn0cpf06qgfqwrr20cc08kxTmUYMoqYm//9G+A
amr1JDEabT9UUn+hAw58lJe733PY2OXBzjs06yiecude1mO2876Xb/CxqfeUOs5f
BC50sDsnsjmA58lwt2t/Yn/Kc6LcSuNSrVWskx2G/I9LAsmBxK//6KGpQcjBiwaH
926i2tGTafzGkrRVLJ3nyIqEYQXDSnQaJJwgjXOwWnD9rGxijW/Kkiz/fuwhwQDY
ZT2bbPvZs9/cD0JK+jLYvXoWyr4hr/yvpMm5eQ4LdDGZIzMDx8wpd8hhP1p65+cI
uLaxmBKb19mAgL8xB7eTQhty8o9Wkw0SVUe/dMp2v3KvXM4JCJZsU5OL9oGuP4d+
xn1nnuJVlS/b0as6dBLazVrde4jSjeXhuG86gdKmoKkvR6IvL3a9oAO5NkKq6c99
KFvwv8RiQ90ygruWmKHaQQgRJrfmIy5bMhkS0F2SAnqUYYV2d4pBN8FO+TflJvC8
StsZI7yXHWXN9hteLVqniFrauELeFJI8QYpR5aexbj3hL/Rb7CApr3SnJ+v4S91t
+0K4A5QgL08XmvBP1Fmha5+sMHjbwRhFiPwGJ5TMeNZ4dS5YsJg0Jupu3PMKAdc2
ogKlpOJ2Wj/ZUtPUr0qi0csKqYBBQMzax4UmwBqJRNUjaZaSoYSo3Xrv40EXsmpO
K+c01jVAacmGqzBP9ZcifWVRAPMJEaZ6Xe2WpBDOSuIWvoYqUtyg+aAj1c3z5Vf9
0KVOQGXEJjES/TX6eZL4kmb+JdaemMPhkw4j8VU8FXHtkRhQ6Onl8jnpcBqgVUG/
YJfU0HCzeEiY19WywXt3RnA2zrPQzn5iGJPe9AafV/w1ynGKq5brqi1BJg63ROql
gOcURihg3ewAkBy0s1vP/xaMc+Tv7SJ4ShowUm436d8lUV/ofCa2nouqZIVWm09l
5ncuX8R1MzpioQKO9sXwdJ6JI4GZhQQa70qgb9Nuszgj8d7o93XjRDGMtKFZp5X8
FSMzCQWO17lLnjntqPb+NDDFIUfVhlxvx139SdqYq3ntZd5G+zKXI85ETvVgW+WJ
B9yOrSj1/PbG7qcVUDetFIdj4fpJibj48KDYCDyr3g8srxyvAsvqn3dQoUQ+dSVJ
LGoT5mM9IGamd5MqQmdyAVq/2K+Xg9zx7ZpNmV8CCtXXqq6fDSqiYyHQkjvfCOcb
al9ChTvM0dNFxgt1Pvs/hHgIQw5FiMme9/MlqBgm4CR4TwnbJjF+PQGhvxIMImEz
W2r9TnRyEqtvq37mf+RCC0/4BAJO9d6GIDHP1MoytcKBy5GzGxzBf/h/1zhWRNLa
zPg4vsj33yeazfRUvZ5H2jeirJjelO1l2yqCAU5GSC7G/3d76KlHlmuF8o59dvpD
czsyPYLGFxvoy6VJdyk6Wo5DT9R3TQU+Rkz6go3qDIs5XqT5uivBgMOeP79BEMC3
yXhDoYYxgneDalAaERN4Nu+9B9f0+Jlek0rVm1+qwc7dfz8YPZrkbKBHeTJPBMnR
+pG71AIPiH7pIphy/f0EvDNQiOrnW3lZaobB2PfmkghKTCoEJp/IvZkQeZyl/m/N
WZbxKt1QKD/X4sQBdTsKT9iR9gSwHQ9dIdlSzps/H/sInEEPP24es1aPcN1Eejqs
/ayDC/iUOJ3sv9BeCJftpP5aPUqpQsFKC5sUlnouzDzfYYoCHKNG2ZEx7eAnOScD
uKfhKR2xmc2WIhVBgkxOzIc0e7+xAaLFPJdwCVwQspQWqT45Na24w4y7cXmQVdm/
9+/yjKl8M40ruUu8akUnBSc74WzhfvO+zUE+ay9xzJrEfJND/n0EWDDzJHgH0Hms
o+Zwzu6Cu+dYwtp3KZslVmUpyhL2+dzTKPY4B0LCeeqm7YwZfV67eBxX5CHmTH+Q
ffMcW1Dr741vO7nzAdHRTMdBupTFuniiFqWKOFSFvbt95qE1Ala3+9T3tBezQgBv
+B9oXydxXKBQif8X8QggE6wIrkUQuYsZnWgTpRWNwL57hU3M/gpd1rNOYK1kpywy
qS6fUVzGimkDs9leY6WvwnTMLaBno9edrvSxqpcbdYX9KBogfUrapIeC0d/mtzb1
8Qo1y+TMoKgPuRjdhAGBaDntY54FWqxDi8/LV1fO7JG/CdHQLrwyHl2RW71CMwb3
HXDgLyMhjI/GzVxXCop8QcuAh5vYPs5rApheKCLQIdA1z7Ho1WUsiaxayj4FNqQr
YohUsTDomfsq1BT7HcOhqrEs7lece08xkCLZQTXmthcdGJlxL8y51+BgBrSjR5dR
W9BDQ/aOoQka71jPPtYTwxdy2HaE3OCDtR2IGLdQKWIii05Xj18wLLZaGYNVgC3n
w5Oiyx7W+X80Jg6FjFIQCs8fTMjKKfr0Q/0xpFuJQB3Cp2ZO9zQPL8oHGhXtcLqp
FkHa24XfUyRyAplZZVyt8Qtmf1R9LsjRHYhcWt8Bs69gOPRwfo7NOjeilriHi27W
gmvgf3HiFNohEyB78vyMWW3uZ0Yg8KDnk9mEx5vNfhulhwbaSrawZpsGB5ZlszX5
ftBRB9+e1NnWfGHMUMiT8So1Dsd+T3S5zmbE4RelCipXcjP4zGkQXM3SY4Afg/qi
y+OfX8MwnvdxPKD9rVTufFIsV4UlC6mf9rbsWZTJNksLnqlKWNOmgV/5o/feYap0
XRi73BUJlI+DmFvAR+aoOMKhn5dIybtjNUEpr4j+aCqAuO58OXzrAl6hATAwCCgD
NaCeZilR//BSXd8Qufhj5mp0HRmZLWK9R5faHs1wRT3j6rKZifcGdFwV7hF5N4r/
ECV8ulQyeBJZZHMZfsxQ08UX3nER1Lw2L9rbkbskXVwhKffhOmSbWBAWfMgVfVx9
O2p7DMMx7FRx+NaeGVQNd376x9uHUrO3syRKDpz8HuPwYQ42jTfBXhg4U3NLZq7n
ffjzB2c6shp4ZGFoksFtvkiAB7CdIEWH5CcpmZnnpQYpU13T0inaUHT8j9ysTcND
kqBOt8CYuuj+gauL8MP7z5sd6yFNJ9E+F/f11ijrlVEcFuTRrAtXGlpzPc4QGxph
DQCzxF7LF2MXDPkqZ7MUbGztRg386ZDS2mVQMS727zAYsrHoWEtHfgYXf3XKAXAD
bv8esknz0Xlk9jJatas5yk/riqqFfSScDlho2TcqHsLEPVNDoRO9k4gqobXp3Ii6
sXzZePwdLqw5qFDqMRzQzubO+k4oZREzjRFeHS7aPabOduZWyyCMnE811l7yfwrx
jXZbBLb96kuxZnSqxzShZRiS3+Yu/IQWkFsICcUatT7rcf3Lw6psgVc/PiJekJI6
JqONdH1iWOLzNTIzuLFhiv7iK8i5R7FHRItQFD63QbwEctKPwifZB1E4NUbwZ2b4
Hf3lxGOMf5kYm6yG6ZKAK10igtEkZyHDC4+UFJQmcwzJPusGymiv5BuCPHlykE5F
ahx3cYzagu4UUvaH7/mKsWABvhhA+BpU4FoP9ZGxnaJogp3q6SxanIRVlQwEYyJK
n0V4qbAu9y5n3ppBCqPDmgNx6/Sdc/JZoi8c2rEoApRzbxRiSl01GDRqPmrZzP0J
gtX1HnC6AT5R/iNEGYYPM6skROgRVuM4TmnQeeRCSv7iqqWelpfyCBAtvQDnBj+/
BTSykNlIylzL29VidSiRTbF9/QXknabyOif55t8vgT5AUdVxA2YXIiV23pkJMklB
5QhytfWWew7CDjvsR0mGfkZ2dQ8MVxskokSnzYettKQuK4lR28wSuNF3rKM9X62g
4awomluxr5EoiacmMwNth1QGEp9n77RHq4suQI09QtrPkqMpxaOcKPIueDv30FJ1
r6VAhK/RtQfMkE6XIePkxCi5v0Ry4w+omR3B+Q4UxfXiRqStsqh6/BYudjJDgiuG
eTO3FMDR1BwmWqxBTDPhwZKQMpYYdGZS+4ffcjQh3nzo8zS3dplIX5Dp9PGVjn49
KQqiljurPUjYceJ8XsyhLzmqREAmkGxs0Qbaa2ntlKAqOxgATKo5MSX7CP3Vrfds
0GFqqIl5twMhagAx/vL500lAP8evmXJRQridcI/eeHuisvy0yuhTvQBhqjIam+RB
wE90+BVI+oS3hvSTmqShvc+lWtx7b5WY8PQ8MJSIlToWVAA2VgvFlJI3u2p3jvro
MtwJRjyPPipHZRh1cUbCUHfguD55X2zFodzTaJokNvVAtPUejy3OylGf+ngFNUke
yifKmv6HzGVcFBDQoDzBfrH5BFKgsgkDNd//xoNgMtWxsUSVgsnlXoD5Di4NI3R+
YeoVRKtA5uDH4jzUqZhXXAZT4xYHHRmHme2lMldv34jq+RT07rukHgspjlXU3ja4
Lr5OTRNYjPnu6PZaP2KPe91Capd1++aTBTuqxDiOiZPFKKKBnv2Cxh20kwWDGq+I
5QgtcJt0IISSAGKKVm8yg4KLBHPDtt+JNogcuTAfTpunWWeMTWeU8WFTKqrEdQDy
Hp0Bwz1+CWP1kO2y1I7NatTLZSGw/B1KEU8nkrTakof691clgFBg3FLW9QS+5G+L
EqJV6ops6/ZjitaSNy6FqemlQSvHYnXH1FMUnhHRXE3ud9d10YaLwxJz2FDi/xZy
fna2F1gWTEhysbIsFECjCvJXVs2XPwIrGH3prKTvX1oq6KA2pnibQFTeI1bfzf5y
HpdtSS3os2t/VivcZzStCW9uHyWOkunPCSdtVmz5fnLhdnalxVR4gMHdlCXxJ6jM
Q6k5F3GtQceXfl9cvTSlR37lKj3STUTapSGz0MzEUhsuqTvr09ZGaZ3R1xrHvgUg
hGXYjQNzaQfUuF3w757TvGAo2AW8T9WRKNDo+WROR0RteTkvBHpZMCukFPyx1T93
vTO3du+M4glIhDXkKGFCBaRyuKNLmAQKbLoa7jq0FHimKKPsN5crMeNZogFVtrI/
kzmb0Vw/wI8gOld60OX06uzEnxKJ5yRxxpWs4u25P6DIYd7W4/29qWYMBMxg2t2/
4X5cE//CBO1p/pBT+t1zZkJAfA+jebpaPrDSCoFecw1symvWZ+CoLZOV00gSD7ND
/tNE6nmhFjeypMwpMHZO3DpW/RpGnc87b4c3pXVOfYwNhd1o3mSoyoeIxGTk8pzd
vXlDTDOdVy+i7Sm9/xPIrGguyJQB1UHsf8RVRDkOH3/cV7dKQYBxgLwQBgsZNHa/
1OstPAFvVJ8FvDiM52S7Px0KncN59oBWzVlH2ypDiD6qIjyK+NDKFYYEd+KGHKfd
Le0TDoc8d9pEvAetyXlk7wq8ozfKUvIX2sJperDe0zlWvdFAzTXCET0GU8FLIjzM
8dTWl2+VOUNIlSwHDtgpGnI0urGjG3jRhjZb8fPCbh4z4zRVXXkhTbBFoarmeu71
0FWIRtJbn4MgRAx7PL8zd5WrYF/wxXG0PY05G/58VmawTIrKam2w7Dl9evfseeZD
LTQ+p4A8nqYVGjvWgJCfQlzYoKKtDgqEwlx/bxgxPHwe40TEs2cr1yYPK/TAuySJ
uh9RG8XLvu9hyDBpOsrK/C1dW1vAUhxVkzl4Hb0nCCP+8cf8WFCCUMhaSn4wEm9E
KO7hoMoyPtPocQjy6ANfwh3XhAuoWpy6rXGiCkC9kVGlrWoOBTRcIpyTcf3eN5f8
JXThXQ7TgFNtQ54uzDwUov/x7BgyGFNGCaDocsww2LxE3s5naBW2kcoJ4q10ai6k
Bc3MUgceNYrevzgFVoLq1LoVXylcusO41VSevtBqHLRqabZXzGRaB9LCZt875E+o
AT64lITTgbMkOx4lZHKtUgbbLAy5oZ1CMKSinR0eovGRpwXIrvLt+2Ei8AYuO1ek
v26OavIggiSdZMK7zle/kk0A/MF2ixeyTJO1QGwEsp2soT6qPv/mvecZn/eUtHOZ
hl3hg6UX3UYr6hO8kUdGnIv4+6Buxdhh4jjcr+QwdJZ5Bn07+D3lAd/tp0xRNvYP
d1ATIdSFZHlY77o852OFxcucJrxCPKvGMoIn8LFm3BAf3zidW6LCbujqxqOHfvhp
YYyNmKqioi1SzjA4CwXUtNA4FaCm5fbsWoBBVHxAByvbTJphKDdtAfNOd2R3rpfw
YTpI/ESZBG/trFf0t3Oqj6zuyjbYx7RqJ0ufRpf2hy54jg8bGwfE4faXhHyO691T
SUeAym3dqBbbuVNzJBpZCm18xtZ+4xCSNvkUlpN+qaPJEI9rCK+p1kcX8OqQ9lWg
f+BCrnfoWzqhf0WTxcuudY/HsPZZmdA0+HoRCrxk9IpOwNTxui2CzH3r/4i9oKRq
tLugyn4WTR7LF7bJ8zQ+KuHa2CTxgqqg0aRZt/oLxaF8/6E6sTYiXAB9X8/0B+IJ
YmTxRXq6yFFzq0YPEd+pFxwOBYK1Z5SFN6/tfu5/F1SJ3dQ0mhGRDdTAWi0+6+cm
+Tg5gGEDLH8OP+8RBWjFfyTTP5MZ/wzHz9W4v2s1xHqqpKe4jLgjj4LhuFVIq61G
yX9yHGijQVVFIVtpc+UF2CPkCgYFfKY31eAKI9cIGxaWvrIw+m90gEyyc2ZmHk3A
Yc7UAZP55DmV5D3eCspNcJtKDRrvv5t8+7wr7dFFPaMpOfJ5g4AXaXeeWZavtbWB
wiJS/ukYxBEapuMPB8yW+eVDbgmSVsFEU+MCvozSz9B93DeuSDiuUzwUdU2BHZ3G
gdNbmyOA18HXVGkQa2F97tpgLI7WhSm6rMQYk06NllKaCNtCYnecquq4dRwhJ7Yl
X9YbNXW6r3b3r3lqEfeHDoAigD6I/KTWUW3KtlscNzU=
`pragma protect end_protected
