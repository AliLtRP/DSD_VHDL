// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:45 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Pja02OykX3gOgJ7gz2YMhNJQq0w7hCUi3e7Ef7jONu6yTlMCdAJMHmgjbWGWintk
pFr3irGLGo526n0lgSPq4NYTVx5lGcmnRAnYcixA1mOdvYzsUQIBQDVy1hyjKaoe
1scjfqum/+FJ3pCmIX6InIiSdebKzjxYIdgMqeZeVD0=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 48896)
xrp5rOwbBVrxUjxxVuWozo6EKQ43f+NtSMSH3AoRoNOZcsnh2+G6HgFhoUA52WfI
tzmCILG7k75usgwAfkL6axBxQnCcmUnmNSJbmYoniuTc+t6zT3B+hwffYQBbYBWo
7FrbUJsTlwGL4N8dYGg6cjmKCBCTMKavWq31993t8SdWpUAaJM6lwT57cOQFE7yg
XQ8jTPKtcmMo1gboDwT5ABmNe5JV0PKzT0nVrN9BcaY895Kml7sM487ir9K+cB1L
ymxSzVgpE5WP6lJGDzHxM6fqMBnzDurBXLADR/GvAzknQ8f6ZT2sHrZqEpwTuXJQ
Jrf+Zq3jqVDNu7OW1HNUQI2Nzf6NIbbOBSDzS4uEOjDKG/zHic9PykzSrtpSf66C
oTIdyLBqtIjNgo79s8yEOZhfg6yFCMgdpyvjT+mfv9u4y/uHHx1Q5XK3NlZ1+2An
rqLxmTOukOZlQnEk28yRCUViqATpWCONJ6da+L6cmCqm8doMQpU1HhG3CAIDmcN/
QgGIBRxHB1QVtcqNFVb1ZdDR8KGZfHRUi9lzIej+qosbMDHnOhlvEQlc+EgqpiwK
jKWAlDghQWPsonbik0XZxwIFUgIHBy9FRjDrBPh4dYzrsfTzlMdwA4YMUyEjVjJ8
JVfO82I5Rnv10W2tPKSfteaUaC1giLF/jonugaPGKLg+Pf1rDV1O4L2737kcosYU
HvDg67izlfyfl/s74yBwnckttrTqBgK/JPZYPy7bgsnPcVVVOC8V6wMe8mIPP1Qg
ivaBiOY6YNo+b7hMSm9jUoZZmHUHIdJgNvq5CMMmTTdxuA7qgA/c6ryJSRl27eAm
JMmcf53NVK7K85ys23EU2RYxSr6Ai9Jj6brPgNZY4FDFxdnXCv21w7AqbEmCWh0v
3PHwk8ammm/r65fB9RqlJxAPu1z64LUnWmMOevuhQcOHsZPq9KrL6u0qcth2Oqh5
yFT4JlVINr/FOMFDkaY+al7nYwQfZIT0LTB7Qsd1CH4oKG8jYSBUPk0jQbD74Q76
tpncsY9/hxkC1gulkVnHCCu6X4LOHpm5IpXE8U/x0foe3Ji+dR9YwRBXRshTSCWC
FPaMmyD/qgr94sXiHVz/usgeq6BVxljXs+NKMyCUkte1I1M3czX8ovTAoncMoIo2
GfJXwuSb/X+oLHEn3E5CJ84bo0lMlOXFffRPqvbhSu4QG/wl+I5IQbmojcgjTgiA
cc+S6ZlMCqZHCUdYlP7NRgwpl1cHuqGJx7Ked46OIu+MLHaPPAbimAGW8GrbpDJH
3b2XQyaAJNMiG2iuxTYcSBwQ+EO0b0XZrXvh1xlzxuKKZf46FNvyGVN43dScb81I
0ohOiRDBoj+NyO8x5JJ4lYUp88O95dNUq5CBCBFDNXZuYNaj2SpOm4No9zdsigzr
YBez5/xKW7i1RrY3G1fp1xP0h9YYU9/XqnVjOT0Qs18+aLy4uKpnTuvuZw++GEeZ
k2vl9LXv+rqOtczfbpXj9SEwhsrT2PvNmDk/rZXMFul6Lo2Oh+wee8jCE3ge+W4J
nBCTLhf5H2G/nFAtLzfiZrV0ad4ZRL6xRg4NE9rd9MofF8O+qhM1uEkJ6ZXsLAZs
/+xEWAVwkF+e5Bw574vKgF+usMWoQtifEByKcK2iTdPreM2dSBSQKeUArq6JNVE3
kXm1H/UkKh9eHT/kN6kpDXr5q/7oO3wmTARL46qgNeddBmUwYj2YUqfLuRfnviFH
zWflGDAT2i6xNO1NluuIpbBB2/YTUPfkI1T29E60hgZXapd6jpq2+KpnKxPmYp5S
G4BhqxFerNjt+AhAR5ktKB2Wc3Lc0VJGtSlxnWuqf2Ma6z2v0JKCPgB9eYK32jno
omtmx8tiOcNkQzs8gOe+dG5cJzH9ISTLEOmSV24MrF2bvbaM+G2BcA2wp207LixP
4FZrojkJhlPnzwBBesl3sX43r39OUzV1ISw/q0TBs3bHL06Po2saFjf16CF1s7YL
Z6k+aKOq6cZuPPlQEyZLXVuY2i3kJ2IJvO8n6d6NJZ/MLsXkT8BNr3twFrOhfMrV
FyOxxRnk5Ie3FjIVK7bKsMaplzQu4uGdkj7F1ObpcfxxRk5Fing8RUxCYSstWcNT
q/NgGBA407h9YwPu44kS+E/ULSlt1FBfhuIoc5xrG6NL9UFqGOLcKjp/Psqnn71A
HTwT8rdAMO1E6NAp9tUrhVVmuxbu5G+50JH1eO2OksbLGYPA/h203uDBu2zUol08
zlxR1A1PhqifqZsapT9xUPpWJJGzVld82n7Jrbdw5F3D4zqOrTweRZwgw2ghUCmE
sbii8/NqFW/omqxBKpMscyJBR7DQzadrg4PT+HF7Kdm/cK126rOC7y1vIKt+2auk
C/FmTVCm+UKRmpmh0p01xjQcGCphoNSZsMvYYGys9CKy/+tPyA8C3CPkLh2DBTaY
etGOWkhWnNaqEp//97HUYL2PMecxfwlKF8xWKMoGQttGLgnr1TfstVWKjglIB6jQ
fGO4q1ZGTnglnDXut8/8x2r+jp8cNrkJTy0D9D1xPG+54IxH46GVvrBLwrw65T/8
FElf5C/djm0MnhW9/t6gGyJMQTGaSMBfAKMN84WlymPyO9018fVudyU3iwbguCPV
Xf+tuf6hN8XGUde/xRdQNU6p/XiYt21GxlefwF/Fl/ubiV/8hvugjwkLwdhvISDD
mQav11c9f8kLMP/Xpkok6eRIougxFTbIhgl2jLqAkVnrpqTnWhs8N2/nE6Zxv2pg
BqkKpL7bzNFKbjQXQKfGCt/0aIvwMT2LYSNMA5KkNysHiLOSlOpMPKEpdlHFle0+
VkMH707Y630SHJFHa42yz+xlNn+PB1/Nz0c00rTE+De4Di2FmvMyqpiMx8Y1Tgi3
OBFBTi+jalRz9t/sbQjsztEpQgdUvhJ1MGzm5lVMi0B6vXzlwJa/3oXHNJymU5/4
uMl/SpgH6FNuOaLtcMxnl82G5jTo0199It0CQDFSjrkB3eKzRZUTghjY3QSUKTkt
bcW19HYpjQp09ptEOe1f4oEzEz8+efZPidTVqP5oVsduWRx2vh68bL06be2qEzPl
FR/IsngJP47b8hRkuqr20LTG3bnqGl7kFYj0ue3ttJl7DVZ2Es5DjBmbriNWKIRi
sxcILGYkO7I20e5jmEY/reokPgGu405nkms7Xvws317ZAVG44DUHM92tL++hWpsx
sktMNRZ66FznA0u2wT04kcOtQxEy/ygivKwiBmOp+l104k1juG2b9ug1QghVqoXK
7N1VEBkAtrzY36TSy8ZnqoyEfMJbHdnNufgRWY5VAN2XPGK/D4LFpuRzdfGuABK9
iBcqfCo3e/o9aZL8YYyBdnD4CO6s+ppOC2QzMIyEUiWJuOnTKzpkWwXyYgEXnjTO
ku+X+nbW76Uw0YSDvPlataj+iUAtM6tjzGS238tCFu6ExKN4RfIA/eb5iiGkWUZB
9n3MdEUGyJ+UCpY5OyYVBjmT3arxYtmv/qIp2iqW4UeOAZcHHMg4++KltPd+FL19
M16YbCnLdOq5W/hANWlrr1X7vGRhr5pQjgJhLCupP9Me03t6Rg9djgTZtGt/+Xl4
8FMJI/YeugeuuXSTd/W0oiEbmL/cBgIbZr3+Ldt3+JZbVW5+DQddmiUZmV0RPXPh
OQ8O6ghw5FRp7SUNccVegdrAmLEBN8/eeVh7K4F1ladVIeXvxPftpNmOrV9y0X1B
XqtJuVRh/tTdSSq9YI34ryWmDWskrbHkIg9rVslXR+uAQcB1l4wWslKX1jJLvcpD
WWi/IkUkNPvOP1FBFyYuKExXgLI4SXa+YZriyA975cDFVaE5THLYvZV2qHV80zH0
Q71wmT6j2cAkGFkm61MgfrzfHCjFXCEod2hhvRu03d/mJ65Xq8T6ruWNuNzR7uzQ
AEipe+TZfnwqQnGvp7VhN3u7n/pph/4o4vAqrTyVOYpxP8UVt9AlgBYQaEyX6H02
eyGXhegA6B9ry07FHmnm4gTkFdw/sLAVeZbf+FrlEm1Pe7WotXgBgFaBTD/n4N4J
98daWLhAkErirGT3qnFO8xfRshZuSg5ZrNgRjk5GVnXDXUfhbnmlrJDYDJha/Bo7
Fxs7WNaR7bfRB6uY7MXuxqQwRoVcD2ehAQ4ZMOw55mA3gUG1hPQoLAZzhyir1Arj
U0nhjw1fIzmitjnM22PXugYbpM/DNVKXYmBo9yzCySLnY86mFDIsIjh2TOo+mTkv
gC4NPfkOKOnbZYDizRnqzAQlUJjRxr7wfN4x8JPS1PN8H1l1YoxqtsewiShj85Iw
TLFaTwdpTnIp+IUqC6s0Y9JMRNb4A1aOqPk6cnim3iw1yn5Aw8H3N9lZZCKuR3Z6
IWoPwf8fkDo2cz4ZJO4igw3Atns/3gARr542s67jndONLB35MSxEeeZ02gfVba7q
6fWJYMmahpZunsygi/pRYt76e3MvRKGcVBySFSCGd/dyQNFKoTA2HqpKkFh6zjHk
Cmpzxd5QfESe9kEth3ZpZ27P/VqYdIkRn00aVp5FKNT/MOpkuf6gwRya9oEhW7Cb
ElfBkKQWMAFZS4bA+asuZR9gMdWPOBw1SWzvC2JyD2h8Nsri9CSroGY+/3gnY8/G
R/Aag583uLVz+uixMbSX9dBOLmbIfLbJnHI/xpIIk8LwpvGgmAjWCcwA0gQP1O6O
wSj3LXakok25rb98xjfBbha9CWEaNFUBms1LSNpIzZfiKsV19FULhOZHNoYRd0GI
eKr3+jBDa7rO8b4Cj0lytZoxTh3Tt97/WtCsOLmydy4CPT6i8ueNKqbAdBxlxTjL
5t2SQrqbzYRTnrmJ7rlEFNwMuo3rhN9kAGcF9r7oBWfkxGOoRgOyeOayU4fpSYxA
bg9E7aZLUfGNsXyFQuQEcokUyHxkqvcwOdxAZIs0AdLcKpCK1qfLtnhWMExfY76r
e5BuzsjeWYebo9y/X6MejIJzaHQVH+sE6gRHKPdvxnjE0J5HqeE6MW3hyM1/Cd84
BYnMK/2We+shJ+mRtRYCWLgxT78DhWMVEMlf7OrzPMeOZMwPLoZPiVewGpue0yhb
hugOCpS1C6gKAJOUN/CT+rSOLSqNx5Njxdibx19DCAlI431IF8I4njmIlDuvcAx+
xGvVyWso32kQ4BcFYpy2zMcdu7rP1kERFtMIOC99UqWx0Hk8JBTb2ZnAU64rP023
HaF4IoUekSZk5bo45AkXK8Kbfj1TjtQKQzGRJnFSRV4SNcMhqGEQFv7Kb7sM9ndJ
RakXS+r9Il2K7EqnLWnWjqOde0X1P2S7RbAdzi8AZwFPgob4SLvSTgD/dypgQN6F
HXPrwKUu8EbPlVxqQlCCisCPXZ8tvTkhurF8AnXPwnd4UOHevBaXwN2X1I0bwfzG
SW+4DrcswSgsy6u0yXo5exTffZcsh6KUWLFYC2BtlSAbgn3QhkEtA2/E9EByJZv8
BTKS7c+xvovDu+eRWz9eSgNPgJ9zc2HFIhsbX1EzfI9bhCVpZodaTqZR3gY0tPAz
7oxvy/+Y7pS7xr5lsiY/0RbJOZDggt5hkyzEtWAXWhjtF54xYbmX0jT6ngRmdubj
iZKP69CN00DN0I89JqqLcNkSaBpo1mv8F6kpptbw3BBkTgM87rnkONU6ET+ZuKU9
Dkl/vp5Zgp02ZrGjnR6I3rxCyyUM64YNgJEyWF8taeYyNq4ckrfWULJe/c97KSE4
q9a2F0Ph1ABwWyQvyCuoD4pc+Xihf/k22RXXTKaZCuavA3v00bWlaLVcy4e0pwlD
QV1uREetxjFUU7MvqoUDvptXZlVepFCATnPn2hkxLOb6K7i6cpUSdzh7soTJsBwn
0odx2rfnUVAZXePYy6hLYvX6rMRpPe4TER22GHSP19vgTxPtTvOmbpXxHsGmJkUY
4xSPQ5XY0HL/ZyLSA1lLOOpZwyOLpQSdGIStn27A2om9HbABfZlUguuv8LIByFa9
tbHkBcO9LE8BdI1hN0M1sq7z3F7j+wCtf1LJngqAmnb+Am1Y+XngIXMgp4Bci1b6
VB0D/HAdvJtHQqSjWeMpyOkq3P6i4Kh4nDGnu/1+UwGPq40rPv62/Q3dkGDBAeyZ
bGhkEX+MWEbU1WBzPF80jZX6m/rgr9Sb3F64TToR11drDC7W2NcAPsOPP3FSA/vK
ctaFme2bfECDlRwJApykXZ0bSuLuAgZAZjjKXzUX3qtfLnolYjNUsRSUyRPb/jOQ
3A6RuFMrFfbKA1BfzYWlbvAFB5QnIOsONXLcTAc9sUlSH5jD37ODxdA+nkbSqEhS
2uMeL9E7oGqUxsrr34e4gO4QqlVEfKt35L2TIYnnEHGi/WIC0N00hnwNuNbbdgi+
qkPXYWu0Xjht8HKeylKuzJcbxy04E0Qo8of38amJuklN+/08/YXBQMP/dMklsFlH
kpJ51DWvgtZO4F1wo7mq8/OU/zR5Q3L5vvhE+UvVhLWvN2mr8KNHky8lEHdBy46N
3UOod/7xQoN+cZa4A2QbQfg5yfJ2Cf+5k0p++KothsBhK3xJY+vxB2hLkP8VpnWU
93vWfrYhVCTm2aTk8RmZzU+5fyYkDKe0a8vtrZYxXkFTRuOrz3Txybx8B9Jq+kzC
jG9Uj5b3vlZUo7imrXdI13j7wN6gEk+M1nxxBXoa/aY4cQW9uqjW2gmZLc2tZIGb
5cBGOxL6wPHx+8W7zddgex4ie0QZs8OU3HjlEuod3MvQ1GoMX1+mzRMQQTkITAxc
udjkJXQHRavCLb754dlx7HwuJoVJzCvhLUfperhR6gFAqzcuwiuVEuUN1KivLb2c
uO0ozL5FV92YCmENitF090yR5us5sGZTKa+8ICx37cJuvRUR9WztvkBfelPN4kym
wpbcb5Vuz9RB6Er1Y/D77SGRRX6H3jEEUJcCyG6Mn9nwKCQeYKSqky6NBq789/fT
26eyqOjiVVlwTAEOb9Hly7awIx2I52vQYxs6hFZu/VUXiX8tFPnEcr5+TGeYG4ij
ZETSnBHkXqGQoS57E50m4GL9R0OMHpsBzNVMdAO4MDXvzTTp/L2pt6FQkmgaZ+/Q
o6Wi1JFsNJi5CtxNmrqhjdLvaKnUSvuLxUbr4SzodLm+5B82qKnyVxbeXahYmAqg
eSkbvV+K9WWUBVSskBXtf7Llnj0eGaFnmx/rj/P7Kh9CuIIOvHEbN+f8KTYxeqWw
CGPHM8dSk/vA3rMpnpzQeJpt5Csl0N5YTaw+6zcZYHPT8526qVaxQoC5F2RCGG0U
ZYjs/izeOwLpkGUJRflPUlrKcmNUjS6rIKcGXk5f92zXvXMzkkXSo3r7OUNKTtnE
0cvom8nqb41uH3vqOHleTRsvNEGz7jJlqrsPWoy+3tMe8RScDf8fPopdBa6PkW1O
xN4y2DeCGj16EB33jz8hqamn60SSMMzdLHgwxGlj+3DD6/PcLha7ZU8WkUMSD26L
8/tGfKxjn9yQfLUyVb4Hq9twfgaL+mJMdIEsqZhR5m+d4aIfbGeGSRAlhehctd70
DIGek6Jzno19fxRuKTG2/j08ZMDiSL8U5cIdRYF4Dt4XDAMg4OHsxI2m5yrPb+oK
xwMxmllBYOdZy/gJS1mxRh1O0bdze3yR4WblSHcIYfTMsAR5n5zJU5CPomCfx4yF
Up9TKF5kgyc9BjgbrBaVBA0UOpqQa6YfgsMf0xZiaENF7kbY0fXZAe3QskuLzp67
tjY3w+y5xdOo70MdDbfJSldEl91atWs+YT0YuBl5VSCh7aTxzVo/przH/+7mN5B6
Mb/durwFP7KVMbnBNJdwGg5/vhLj8W/7fUFJJSI2WhFu3x/aAJY8EH4hFvYVH/sv
62pAD2LPH8VO+hIOOCoZ33qucC2uTNi7c8Dodr3DecDt8gLoq/DwsAJ+0Cq713+d
gArjU0vAu5JccDcjFY1YeGdUu32v7u11hBmXqQxWsTyeaFLGrpH2nWDTXbS692VG
Qj2zYocFtsfxn0S+zmLS2fce47ul4FaLIWKxZhchbE/+63M1k8cmBVkv5OANbkOB
2GXGErMz1TgVj4KMlMZdTBMnTptlC/C0i0crlL1vf5ajtL0fbfaHu9ndZeYegYM0
6bfWNw/z/oer/Jq+Zvm02U6Y2reb7XD/U4vCdFzB69r+JpscujpFl+B5yaq5viqO
ZRdXIOsnKM+JyQbLwN6tdavC2BSKLgG8QZc02gfHG7iotNdp06ci2fBIODSyJsmo
oIzty0SZaNyaeykVhGZcaPEHqOi0/xShDfT7cm+zE3wk3cfqt+tZG86dSshBF+1A
eaQKENW7XUCN2lXD6YRQfovu8TxbClgeU5kLjtTSgdfWE1RXE52SJnLnpNoaoeNF
E36m2rpGjypmRgRapHUV0/9yck0H54yXYfVNu43h0nFPBHs5Ho+7pBtp2meZ6o07
oeSBw6ry2/SrDbRTIbyilBmJuMwHqYmSd9R4P/Rbz2HKMRn/sj5B66BFGYhWICs6
lV6sNYSKXQME3RrZ2KFX9oxb6WRH88HNBjgIeSNSviaG6yxi8yh0fuTdrYPf1SMf
XvL8050HxpCSzhi1Row80rAbNxkW3L+OiyFlWRNcqrC80d8Ps+R7ZviOjMW7qky9
XDzjLAuDZg3Jpb28qASQwDRyMUFVKL9c+hUxu2E3ZT1FBzV5Y8SZg8Cq81qO9B0D
cbti6jkH3f/FHi45hAdaSpVpGF0+g5eLc0/YpbkSTmy5MqzbqelqMRCso2bRwv49
BQ+XFGSaTJkEz4HpL6laSnEYNgWBihBuuwqw31u/QiQPF+KwwYpqoUH0Xe0hGs/o
Mp+EoS+oN+tvn+RrmvtQbWKleh8R+SVpw0WBy5X6Zocwn6DjeRs36gYddnwpLlYN
1xuqER26IEYWS4CAk12EdlikY+416R8/Jel7uMwLDLICQKkyDdSGfLftJWJUcZcq
Hg6JjpEkbmNGQHHZjXgD9aAaXOykI4B/o343ZqeM0OcpAtKrsXzVnV3syZSBNJM8
1vM3xcSv0JgMZv6f9YsXii3XptfDhNCjg9WxPXTxiUX1mBoSiC5kIXTagsQHK5Gj
fyqEmd9FK1IyvFK5Wmb/v0EH0X4/nrclQxRQA4MnesErpu9lzelJxC77oHrcgInA
I4Q15NJ7rT/0P8ti0gLNi+ZW39743Q8e+xkz8PUO5CiaE89wN+C8TCy6AWIBEEkR
JvZu6xdTo484i7x80qaZVhCP7Jwqoh8aGgeZYl3F53ABTC54FBfZXg6yyE8PVWIo
gRVj+8eZBfw1CcDynLK3baG8lZj995QNq7Zkes14PMhIHEAmkL0SagauHgl0vLk9
xvYjOXmJJDAoxamrbn5JduA36h0XDpdkF8Xmv50cKQBPH0A9UhcxUD+KMwsbEa0V
h0dISOUmvdwEcO/W24r508ZmnOq4y6p0lAjCc+8f+qbGqO3BaTK84UOT5s0vwCbp
Xa9ANFf60keLQcQnJDkYEWf3aNacju14zstSA38O5b3Xm1H4vt4erwvGGA5QFQ1K
+GFbjVcMTwXY0gzQ+0ag6HvqMMLk1zYLnTqGBtFHfigBa8y0/jPNO+0EZ2Jd4rj6
BoaEupLR2TuZo0Em52rlkuyHzeRhAfx3dp4r66dhzVhG2mL1wUQSP01VKrnUCWTN
33o3EBzAhqzd5B54W4bY609IwKfXPfGDPcP6s4C4u80QFaBZB4pCQ0F0v3TlYjjI
fo5g7PlJ9L9TYt7EtJX0LwrIzRfiPOr7BOoo4cZrm+cHtr97re65eo4ajCKu1Xas
nWaqyZs+P70da1rDwN64az22m5XodADgq95X7nDmRmSJO3EZz+ph6CWKWREiefD+
2RjZ+NxI+OqUA7jPm22oZ8Sav5U7B/s1qdOkcoEJde1wPra0bRFim7X1edFPe2Z3
gK+7yRSCKQUPmC+5CHG45QKS4DxWuhCrsE59dp0kjC6hwebei4sGKXQ1+R86oGAR
RJ524yAXwpeAepWPbJg+mETJXifb8b+GQaoAC7fv82vrxthqh6VRjdwoXVZcHRSp
/a72Uyrl2TZ/0eo/wg0FS0gC7b3ISgkcHtbF5LSoxbBgVWFLxWGIeT+YdaRmsjxE
JWfE6rS1t+ZFu71K41tof7pRnyGCsSuUgkdjhm3994EqaD2FEzoSWEHmTA4wrhIM
4XYHK2DKNQMTAslg3ZcmZktRiWu+W4HgH6kX0w/a0HLPwPZPmQMfyGDeMtObBnV5
EEsrYOMzgy4TYlOtNiYvT6IFAnKyUa3oYbxaDG/f4sWN/pcyAgdF0VUqwK23q24U
9r/cWwqEtNtqUUCrqSb6CHIOEF2aPNDm6wGSp8Nz0uYNJ7LmE2DZtOMnvAweznx6
batc4HyB3RMBtyY7/E+X0vZtR4fMNUjItKY8YreI3yM+KtjxVDkpRWYaFSkoB5X1
/fI4oRylDjtKLT1Ik9DNWzpkH2Qj6mgiJBxD9jv8GmZIDZVQEZ83DP9nvfV9ceRE
7TX6KSC6Q4emAYHY9SnNxxq/feQM3SEFb1xP9CK9RS7wxSbM+2GvP68m31CFprMK
n6ik1eg5DvSyf9pnCLiV/YENvWsT1tRPUgC++yj/d39xkDkGyQG6pr43pvM11LSJ
l5773v4+kDgkUA2NM8AJ7UOPkih7K+tayswlaWtSl7tqAL29EtcLDcSTYpidwG5z
eJVP+9xyyRtgzSsJR3PM9nMIAFS+4GE+X2L40RVW1Ugik9J42roBxzAdYYRXQgUD
fUaNNcH8HwurfJr+I6IsrHC5QuRygMY2sGAuA06pt6dExPvpeuJlcCyAExf+ybGl
vYc+WoVnXluriRNnGmMqr/IREOikgkeDjh9NRiQknzbHXnJ8lcq6KKOFRUd9xEEm
wVNWaGa0yhY1RC803jXmCnHHWzU1WB7Mw6b9lcCkNCtrmCgEl6KWpox+psJS4LXd
I8utaz+Q9v6+/uOfqyDG15HgKO49AyHy9sIGxAlCc8XwnYpbZtJ5SJ3f0y7tkUfJ
8l52qz14qkhkKFRRxzD26gq5oN1lhsQLzmzHYcNqkn6BL5Hiw0DRMsGPnu+JXD4W
+AvEBehmVzClC8POyOrNUnWJll/tIvOZwsL6rNH21V2NKJW28vUmFM0LJJASp+/I
sTEBFzGxLY4/eGcV52Uv40583Y36xaQivDYkH+QM+9hgzyCTjJG5wgAug04bXdmw
iqTV8KgkGwt+pxEOqvGF+JN7+Alp3kCswM1rKan28kSG9YXXDN76v5mglDC+xqc6
GfWioW57Fgn8n8fM6CqaQkVHJbvoNQNf+JYz5TWK5iaEWl1/rguwgSGN7Gm7M/b2
6NNKuKzI8r4L40HRkgXaeCHL40SYl/VviYTy4GNQU8IP/1vP2Qm6M/QDwzXIR3wM
+x6iZjBwXMcMtUn3XTwzqV24QwWRZNHNf7FxouxGx/2wctmpDlQ8CpoBu9JMQ6t7
mzctt3G+BKZvolgtFp9eScJicgzH5Xs1gqCd8FCH0dMdN3JkNT7aHLEsUvwl+Q1/
eUw54rP+yT/OdFovpYmZsfAME60liBiuctSqV+uYZ5Khja0rSjiuFrA9Yp/Ly5LX
uSC07CQ99hzMzewhxv4f30OmRqmecFb0OeP7VR4Szct7/AqBANVNBuUV7bwxh7Ff
4vmUvkDwULOcZBOLS7NsOwgcdF7WBnlGASVTeoZuv/cSmmWlCWIXpvsTOKpqy2Ru
f75EY+2RhE0l6W4grsAyoACfCniWBZa2LFtNGxPF9+UE6qgwNppAUku3KxgKqEeU
nr/Gp01AQ6bxBQCedwE2ca11HLhrpNItdO/ne7/+5hizMqX6fWuuzU43JJ2diUVk
HfYcB6y0qyN6nta2F3KRL5frt1f+shpBgV64hpOZSKpLaHM9Wd9pifJ+Jqr+eBgY
siCyOC7385slTPiYOaU70EvzTNUbuV7BL2/FNAIurdYeGnnPKf+8yXY5RB/Pn3D4
7PUghGxTxHF1yLuGE+Bfnd0F/J3GCddVLdPs9+FE0IpiHnyj/WrDJRwredT/7BzA
oVscMqNpcW1IbQbLuo0TvrCOsh3bL5+ehqpkbi+BmtIxzhUi6H/JFg6WkLAqr6ay
hWcfgk4WMJvXt/w9wmPhRV8clLjSpeKt39fmQH3GHpOg3TmE06TPYi8sCENFjMBJ
5jT2igHtmU6IE/ye5xaqcV9kWrUH43OjCvYvkDFH4/s6Dtj/kMP/VePCh5OrXdJ+
ntqr1jNBqN1T4pI8t4SGMsWrf+lsuT71EENbhuwVqvkC+pTrdR+EV3UaX/iWrFHf
ox9m84robBnMoLF5oUexjWUIkO6B7tszZvVsl3te057owVFmukOT+5IQ9aDLVCSN
xa/afTj356vUIMyx6nq9HKy5GKpagFAPRnUFPqCJYoAu33yVw8Znc4TTox9srHKu
rtaf1173sSX6iyAPNeqZzZsW4avhs7ayMHnxkXcCc4KcgPULvbLgsIWJg98FMUHM
p1kZEHvFCxoPAjK+D3+88Bhsq6I9mpyUCkYVLp61TUmkPQ+KuorE4YjnMcacIO85
ijbE+HQZ0IyIfbhEEoJhIVnLbEXv2jYHVyPVd/B2CJO+KJN9+4pE1YBAhsZVdi7z
HFuCc/ItJ9pPJhDF8HKkE7wEJQo4QeCtWvgG7CZEwPV3qKQiT1G7shq2VCKj8+8e
kVYsFgVteQ5hzSRSdgN3DjGzZF5Er6izWrmzrwR1MNKAL43jpyDlwSLv+YBVrkmE
u+GewS4//okxtkomN5/XzGnfZIUS4Fg8c1udRTxquzB3GzX6FV7eJvrNK+rKyuaE
NfUNgpQdgG700WUteO5WZ2AONTx3U8pWRbfEyOPxxqy4VaSS/3sVzM5/sHCi5czI
j7nlCtWbVfWte9wRj1R6aVojJMC6jCdbNzq13FSX1kHfZHtHcShKao9J7rW7nMmK
JUGgq7op1SF3PV1MN5UffKzY0UjTuUTCn60soUaIJOQW0ZdnFliiG4v6Ogj3Mt5j
/UxLU+d0P5bYAnKBvh0MyWAunPvwb3QnUWN7xppDcNS1grphF1zuWnEUWorL5j1h
Ou5f7A0c1HZII+kwgENo/tZ63vBe4e9Us/S8xWTFuZp3pn4qv7UtdMG7AKj3rIjI
Ylpdc6sZ78/iaTcFXXAdS7b6R4Avh8vmnRNTpybY6f6vMzzVpe7rhTxDjBkxj6pt
AGqwLwSQ+a+xDMkogiaM1J/TaxwkR61796/t5V0y8AzKNZn8B+wnqX8z8ZjbqncS
dgpqkQTuka6jWG35D3Kmx5YRHAYWkbd0tGV+PvmHmPCIYXMfld7n5aY7/cS95JD0
kdzv5+nTt4Ls6MHqpG4za6lLthaUwLc+0qDdfHsrQDKIXMvE1Ii6H6FgHluTXP1K
2MZwAsju7uXn01N/DBsGU4NiTJVme/zYfa1Cl0x0gcfT6wNEC18g1BzmJ0NDbwKD
nA0QhJHJkTQ4S2XXvIiuE3dDPmhF+Uz2Q2nKwdkHzXdZHhkrKe+BUSbi6MB7VSBH
nCTr+4OJkzDykD46gh3qHZoOZr0wZsT9meJNuM5E3gfgCpOXL0OKREVe7EfCbSkD
OjNc2Urn+7p/QpReT1cHqYgoJzzmJaWgL1o3babmg3EAYLtzzldpd3v7isj5Cse0
AOoKcbSoU6rMrTGxW7MDEYdWewazOwkBzRnN4iZSKpiheInL6d6/8MDtWSekOMuI
gqtA0xnkUcGO1FAEL756+AExK8bHG7neQMwTK2SHIWFfuU7dSOyPJdmtvXc9M/Bq
90JVRpHN9x9tm3DW0IAqWGucmfXYdpGomRKXwiTkmc6dHcDMTSHCKapycLVRaIcP
fwGxJsYEsw+PvFTQMfchGswVSd4U3Ofk0jO1wW9ZdZIbARvaiWxrpQ28rllbiEhL
yAlwTeHJBtrxU1Mrp0iV9T7dcDIl0PMmIRmvRMylq+SuD090JMKRpfj5x5F8Lijz
uK9UgqFdnm7IeH2mzxL8TPAgqohAd3f4AKddTVSS/tMEZxSK4cuvdf/I7fG7hXZ4
DvtedrCcb9UMKsGMWDQF4ka6Gd8WrgmHFBTZs770fXiIKU2Q/6njqdrCl1ITe19M
sLcK8gX+cKFpBaklgor1B4siY6BPuHgElQIvIn8zNQCWT/xJI+nB1mvR3dpsT0IP
BSoXjxnjBGyN6dn+lJMS+Y2c8gcu2pUUr9fO/ovOEClK6MC1r3FSe3HkbY4i4gQm
sbilut9QL43PlirIHPDEHxdaVbpNmqSkI7w6+FnGC55MDBF04RqKY9OrlO1pWBdf
tXz7wsx1E2KhzaE0GH1zUUra5O+Zlz9o1QG2GgEl9VC746XNFYiEeJhTmiimYQbu
MM03QiVbfn8H/ykmMfNgwK/4pdu54hKGwiqG1eHr7nB4/GUO30fk89y1PMIHjPus
rHmOaa+a9rg8oQ+j4Zz6Vr4Bku4HD+jiA5kUlcZBTHIe19ewcyIAa3AeXCCRVYuH
NuTJsnrGnFkcv7aKGoZFvOSdPki2b+zDEuOrsB09nIIUl8prp1txNUGkKVgz7U+D
IDt1yDIAQ3B+LmzEnUfoZJ/FrbroYxv+SczvbQiL4tJ/3RkUHveYLqc1Td+RautD
kruSj6lf/JCQeZPDLdU754bcw4xhyuxc3bhS6eoCoiuMPFJIyhYE5P+IzvTNvVN+
wuWL4m9Z2lNlghzMX3hUOWaWdBpMm34ClV5lQTzhb5vtEcfPzciyIyfqsDBS69zk
NYgq25x3E6NCUAzt7jGV4gpBeqtASpaiyR2aLXCF2oAn9H6j/jHpvf4QyT33xs1g
rVxpnnOOFfCJ788jpuGt+pNanBjeroVkDPMWsk4fp5XmBcqemaDzWthjh1YoEnVW
332YPCkNGk9VO6gupsWyfmE2o41UApN3zmYFZn2iOFtji+zF3j0BL98BmDx7GlU2
TrJQLjJCXD9eWcWIeUp+TRAFEjqT6AYxLcPowMuRm9KYXsLKJzgTnqp3U5nGDYUw
Ee4U0OCESPFGl+8/dPOv6K1B9HBNPo5TwecXtc0G5uXxNT30OUlRUYqNnLKW3RNL
HCcOSPJTngJLtz6tPsbCyd+k2b8775YMgY9V+weHb5qxkFFSQZmfyLv1ckwYhZVm
mqsoZ198pnThlsi7U+UnZzZWH2qb6oB1VtesR8egt5imeCw/YcCgkYuhWDyOXdfw
TQT0SEA6mXCciLl9SbNTX8pu5+AIJuNp0xAhzc7T2CD7f8ei3Lnu3hpgxtm1J9Hv
KGzY60xPJ7YkUzrabarfTPuTuDjnxaj3R1qBbH+ZuO50gtEFauixsZyXK923qlIA
j6UVgfkwomjFQblmupeNFvoyWtnbiioCA5krhZ6mQlWYS+rzMJ/P0WMpvA7wgU7f
6RV4qt9SNOH8XWD0O7ajiKAQBBmRiE52F6cbb16yTLpn6nRISPyJlAUbgKSPcc5Y
4fnMiX7CIYGREDJx3CqGHrDeqdouRGehsJvEMZp41L3mtRk7a1fIgiV/lX3O0d7E
AWZqdldVSw7EKgcQrJrPUqLxVtqbvV+6W/eImZaAskELweb9TX9+kE7Edwha9Ycb
dQ8Rz+Ga8tcxKrBtsFFjB5D4YIQ2+BEBEajImxoUulG7vUDQoj4gSGcmo5rrUrhq
koucB8M3eQjPdfc72gtqm/EE859SVeoIWyqjTxrTxP7DGEzbCzPbS4c5Lgl3782Y
7BMvPFCjDgWcsMQ0K5VQVo8r2wotjFBh9hKTEgMzKkB7nujzjOQ0f2siL2aMXOx4
XCyt7N5aqp3cfKqLIOEPh1n2gTx5lw9ElmOWnQUWPCBDqNea1oBd9ad1XHdR6ap4
1MeMvQAiRRn3vBTgiVGTW7yKm/zaJfvVw4d+WwLdwe8MXyGeiQJX6TA5fwWj+ejM
iXU2l+TxX9GlaFgyw3LDR8kQs6qRSITaDv1Z9DGMP6wB3SGSy1vxPAyOXMC7uIkn
qDIZ+cTN/98RDLSg4R38n7FzJQm3hDnzo9U/xgrIo/VzaKTYDvgRy8SFrWGpUhKR
BEm9dg3qga6f+n+EYw3CK23gMg2DuozOVQQQ0yLOEaYCSll2sphcvHxE4KV3YzoW
H6vnBXJ3BZgqiSn9q9WZZgtZIPu4xptgCYcs3PIyWK1HHtEh+08BRtfjVWeHrEch
Q5wcfknHv26aolt+W6SfEbN92fv9daBqZ8CG9vCd0/Cf2n7U4hzT2Hv55VXrQUCD
L2j3yIdUA2pCxj68JdHmpnOEBXYPk4HrB88kIo2YLWiSldvGA6kXL2toug9GMdKG
YEUCDHBhm8k/Q1zfzU/oClGw3CA6JKhDiEbX4jkw6ku8Mb5jQWMd7rmsla8C0RzB
uubwWooBx6wKtswDcsFnr1d7CMBE4RCNPJgJCS6xMF+gmoCzrhQ4d4qiMjHBSCPL
hE7ZTpZKl6dKqkul62IhF53sSUSCerjSxZzwsD6bqPHCszeNoXUpUQwLngwhYVaZ
95RPDvMJRjPUem01/wZ2lPBodXrVYO+mpYtWylF2rMUHoVQOFsM8QHezmGnhSeUB
09eihDLm7nZPTe8sAUR+2E5AgIoc0fzmm7O2BG2XvCj+/y7VdHGxOv7Aax/w3C+M
9itTwPyPW2Zioz03WHIs1aApbVChGZHkRF+igA6dqXjxB3H1XJ5+czIhOk4UKEXl
XuvYIcU0jaK96AhGE3sjV72nVnEa81GioyHlhXdan7Z3n5g3QRGH6J7wVSGuAy5g
iRsbjKyXsrARrD860WazGJkKMIAa/+0n0HAeVvTCCRA22v+ZerZRsjWvJnGt4IIJ
rNG81DZLWfyg5kVkc8v1tTujzMJRi4iaTs5A5kR3gGRLeNJ5MXfPYcf5B7zdjd8s
iztIdXT0PC0OByILuVOUCdKK/ZFkcf982NRpI0nZ9jgwfuTBochtUZDWFCtLR6r/
ZOHimujZBIduxS8GIvIx/PQ2C6H9ZFeX4U0JPrI6RwYUs3F+fq3J6G9pz8pIr1PS
S1x+bDyEQELWzdRIwt7xL/aQTSj8AgQYthRPhShXeeoIPktmUXB2mffdhMUARCm0
AZsWOQd6lxegDEcU59euF5up1fzb0Su/LezE6bWTuj4NOSgYf5nREW2aKiL3uX6Z
5jFzugWVRD/LqhNh/4nxEevDeDoxwMowqfDcKlF3tO/beQvgqJTLXt0aK8HSaRhx
jttWXet8TJPLAvVvx+cb4/AsHwNKzX6QRL2rgDqm24GRr90zN/Zb+YGceAcouHuL
wWRDOTesncAJh7zi+ye1eA+D1fDLfTCcqGGo0BjGQI6EwgN6tcy/mnShl+8pSMbl
IUEYvUKuGYAd9yZIJRsi34ik5Y8FbbwP2+TsJ+PkH+U582K/ldciqidlOQrRmAUw
5F+Mr/mfdLtKPSvf1mIt5lPpcZ80DVd8ixM/azCnQGptWAxbBpt9kKuvLWJP28PZ
uV4D3mRYCs0nCJ6Ixcyv2xiZKnJturgvfqmvhrHPGOM0asEC2fhDx9tP0iT7U0Pa
FIabUySQKQmlaiFCW1t/P2yS7silu96xCUFdOaGy4egTv1kfRwzm38QCUyDr6ohp
z4ijkAy6lQovacvdQXqsu4EbcI3z8cS4x2iKq8kqir/Bngoe6Z5pB5Qnq4S9H0rs
s/D0eNqlbIuAUpSeIRGWAYi/H93qVNzizIusx2VRDo4LWysANcCohq+YIOigv7M0
EYZJCI947DkYy9KHqG3s19yfBvLhQt/mYialF8MNzTRsjir76wSAtu66SsTLvhx6
RzbOMV3iq5ANLL+OWJCe6GJt+oDqawRecFaoL2hRVX3Dyb+Zdr5gJ/z8HCBnnbyh
RdVm+UdQtarjJBdYDOWyvyAjzT9l7KtjJW02DvDt0bnDOl53yWh3P7nD5YSYzzM3
djr9HWTSNEUZL3nv2oLlUoJKuW4sQ2gvguHZsDvJvT9WEPu6sOOILxvoQ1o50Y0N
eLXcCQMnNGMWZ7oatE+wKHKQ7sMcjTWTOzXdcWOLMTD+T7pfqL0b6RwdMB4amqVn
1LYfxh8WVrZ3PGiyFUnSa/m8rU0ly1gT1AoQHX78atENSCdtw+YOPUJzOFAQEU73
agClZWm0CUBlLSpIXtoFJTybPTq7/666+05CTTSNq64MVjywEcb7kUNPp9sFNs5V
a4tselEH8s0eVcK6aTH9iBDCyMH/Ks2J8xyvH2D2lNSwKIzy/aOHlgqCdZWQV8o6
bLjLWmbZDYUPkM3AHwwruEYnV/xNHtKS7pCfWx+n45rMdQPpjBRf2z5i5FSxTCBs
f1exvodl0NzZ0g6R/tPeec/aZgnIHlLAU6nKQaw20lQ01wbfpqKir92VXekLS9Mt
jKVoheQqiM1lvv2ac8CX2PWpx0v5uT1J9fX+v6obqmIkHnfPHL17zri3xMJcvobY
0EsEF24Z2XZ9zr7GtwnrGSE/sgz1t/fOprALxjboNeDzwsm21yjp73lB5im2hIDp
/XvUw0WdpgWLyUmmCMgIaA4gpm5XIiffAvrV2ZqWgIwbebTtrRziBVuxia2Exwtc
PZlDaR3BYaLA9XH7AbIRebmvQ8gEBTxJr8+H7mmpiLMCU0wkRJGSGn2oaSnoHSSO
4IFJJ6LyErapgcrJPRFEPZhxNqb+TTvBA2egh7S7IJvOQJ+6ba8pPUxdLPYM4exw
sh3aGBhexIsAnUe6tGAmlY+2M5hq8IXhDH2mGyk3e/VJcCw+cmN77ZeSrpBiZS4j
gO1QoLXYkQTQTGzQwG7HcViSHIns/bUqrbxKPrSDf5QZaMiBUm6wfJGsKFe0pnIt
7RVRfyRC+AqQpK2mkyf6P9PQ5EEG45DpYIcLEX7G83HMP3/HZ9AjfdPXQAN8FnEJ
7qLGtjK0d6PyLCDgDWF/QvhYzOwSvEHlhBt/b4pnwUlztCp0VWH5DXTxE9mCDhs+
NxBcx2NDivl9czLaiyJsiqXNob+f7MxTgRIn2Mp6sXZZ6KRv1u+wmLEO5PP0aWKk
Ukb47h0m4EZvyq523F0txj2Dph/nwRiRJBmGVewEV8VzuHheoChsGiridCB8fBw2
CwrPTII2SR96Low9rK0Ia/g6nL073kcKOo9K6TLKVD1oc78FbbFj8aR8ZmIIqW4j
c/O2aOscmWdFtIH2iu9C9co/y6W33RsucYPWYeQDSR2H5+N+AWlTYcRFnDhCc2/Z
H1vtSQTphks6x4ZQYygY/MJsZAoKBrAy1kMyUAXp+mQETyFgc7O5LCLGZIfxt/tq
ce0W6RAbdjTS0PxFEM7Qa2iZrGHgONZttWqxMyLSC6DcRs0uXuhul9a/MBYxdX79
kjR/kmSlb9k0YGmhsf2aZAbjHMkm1xaXk9QHq/sP/wKlRklW2hO6VKcvqhnwKMd4
Mw8gHFo+hgyFlTnUFIfRjJ6SnlFmgvPC7d7WGVo6LimTqypH09JZYurYjcr8SVom
UQN9osgzl3NQhU+9WqpUlGO/pHgLt0Peh9q3gjvy9BuyEuXwnG1gAK2xv7pjeC3T
2I81Byb73MzoiRGWsDBBOcW8yaBoXdnnKN9EAUDbLBUSuiJ77AcED5ezoZJ0R/eZ
RAfOr6LboxhLwVz08TcLV4DUaGR/HS63R9aGQMDCsBVw4FgCXGpWEoGQGZo5F+iJ
UyIxpmxZschC/HFTXcjvCx6aSqesa6hVBn49NU3VZ84AulJch8DnbUxEEcOy2lgo
V02gVnbFzTOf6Mbu2dqTjj36lZs5CHHZO+uAfVk55OQpJVXbbS7Bak6Td9/QHu+r
VTSiLYR84tNvWKFV+jj86flewRS+hWNS41gSvdC5SYklqH2/6+Ufr3zdFrr2Tw7+
4Lvk7bxM/WdY3Q5wg1YQ3lhqG3i1CVJDds2sQe1Wn9uYjpR4T7U5YD3tk9CbnLDD
TKa47jSRqFuaQkG6/xvUbRyjq79UqSV5+h47YGXKE06Tm/15Lfl73i0G3fCQlYtH
S+tfA3pWnxeJpBg0ljYycZ7gTEzVOfMiaRleV+B3Ev8t8br2tk2Xqc/CghAlIqyg
uqlhGBeTUey3rogOnrVWsBUABU43vi0DwzvaPcSuNh12e2hFrPDDaeqZ4wEu6VDt
3RJ9ahZEv/M3+j6DwmpxyD46gHloNZdrV53iEPbQh2m5t09LPiJjv5o4NjO7Nvvn
x/MbySqxfQbbPopSkieK6eB85NBDoz8uoSV+bLfej0rWdGgjYNdETMgi+rswPgRZ
VkFnk3esuVemN7qycCNGpkMxlK28UZ0TM1pyt2MixcDpJm2wGSmsi5gPIhD7yLq2
2/8a7ejOmXsToOStLCn7Tqru2AmoWbRely1GcmV6vDyGV3lEJ2Qg+jOUkv1gMhuQ
VPmSalxiF7npsde55Mw9orJQEtTDdFHILChjw/MfMloSmdgt1sX7dluJyHUevp2o
S7v7QeaG+76tqtxd9Kt+ZXftIvOLDVk1TiuUnoxoAbyJUCFFLgEl2sOxb4hRfFpq
DzTQOPTSA6CEN4zgewQTjaXlEDEuASHg08mng2YtpPw2RYg6ZL7XPhrmyD07wd2m
qdSrnxKmrrG5KzrWoA7zFjnGPJB+16Z3YRIrXEovglVQ3/vtP/SVSSae+8mZ1T69
a9aFK7zs6i6NTMGoy5XDUZdd6d8slnLfjgkKN0zavca78O9URo3MogaEFQFpw6UQ
EUCqelPWrtCVoMZbmQONbylHXP9q3MGpizs1wRvr/90nSt22PIVubaAEEpoEFy6F
gCt09/OYjKwPwQ1nV3S+LWJOsD8jCg4cc1KLX6P5f9grQMNGDIXOVNCylQoTiMMP
iYMbYVm2GYUN+a+Z3P8HgdSJBQriHgsSK0oKeXae09fCGTkvMfWagfleNpZ1UEnf
B2RAh4vrj4UN58gNEle2BBUJku+UQdf8XHrnibo7dAHv8bTjrSV8heiHjs8Qjjaq
H/igPOKdvoyyEVH9PCeqSfe2Itkg5NUwHb8LkC/M9XoCtWSOlw5rksw0KxKzQPha
kYOexHzfZri6NgGZaTZx8Wcyzp48IfqC8EfVSskJV8k+1rZYkCvdQ1QXdBMhnA8o
LHJQ8gSUrYi6NzwQg5r9cwBC5Yjgq0Wuzbu0KylC6IVkM9N9RhMcZrmR+4Kwj/b4
AhszJsfOT8U0IZcNQQjlzdlcxkaDuv3QdKVa0yc2A6NYxoVvi71k/uOTQ+dGiVmj
L98evr55sumQ4UO3EEYv1Cwg0ks89rY0ZYQeDArlu81WDJZqpinIkBEPuhtEjpiw
50ecJlRnaMSw+f/fEJj+V08qFq8+rfK6SXnYHfYXUI2PVLMFqfoOZ9UnKpRthW6y
VLZM4esvIpA/XaGgZ7g0qEwuHJoI7zKWYZ9B0eazdwrvyQztJPJk5jqpgVwe9V5p
XP6eDP5sl2LWx/nZ8PVXmmgWtqogSRFFQGI+i9y9UIGDntYAqIffVhLZBX2rpsn/
/mtq0HmebZWxKBdNmB2BNtb75+VW8m04X73FmPnWEeRZYRby6ZPp5JR+XJEXISX2
haj5qHYRHAIVq1kKpmS18jpG6NdONZJ48WYmxH0Oy8mq737JC9RtquDTeOFfgWtA
SG/QaPlpTdK7fzte4zS9lcrEL+JVV0oC0u4IvnOu+uCMuQZnhWSvVJNDCIMfifd3
l18MlgAcHjuKOvW0/GD2ZD0mgjcznyGT+8Igs5MNZazoBIpofbw6LxU7rKU3pcTT
puzWGY5JEKvOeQ/AejeHv6yuaHJ+F4Qk60hqImnUbZEgpJsGPP6RSQW7Intr6js9
7kNsFIhhWJQKDJ9nuEib7O0Vn3chyez2gVesT9ruPNeboTa/xJ5cQ6Ky3/1E8Zck
ikcpyXZNvJU3d2nMGrNMwGDvdqvIFCvlPlnICbyaFiHHneJA3a2YIg1635cJCUqn
JTYajhB9sw/Naiu/VTkXyYwcEMLZe4RByeX2ePh9HX6c9CGGMuezv+XIFy8VHXJr
S9DKvYys+JIGm3KxTr14OsVND/LZeshX8P/+fFdAW6OxYuymFZqNb3xn/Mb2zEKt
DmVv9jVos/olsv4YiVFJfbTVudyXbOjA6vvjnQ9KBUwhiV7H536oiokKoGhAInr5
Vwl2tAXCzrUssmbeyVRhMBu/9nlKAXIPHTtJ/sSXri0HLkVaGE+phLL+r3BFPU06
YXH+EdgEmIjmD6cPDIW7UVJW2wrJyQWRBPcl28KqLWVEqDhCj2lIlVge3caKVVwc
JI2zfCnFwc4c/oJVY1Lywz8Zpj/HZEowJAcJJfaGPt6DGP2jcYHQRLHME9eWjw4R
dzAH9EBZrBf1K9FLKr08O1DzzByDLTALT6rSUKQiiatOPLJiSzK1od7pdn2RHPqw
2sFA5HRqA+2zeCNsVOpcKHJwtIk+1MUsnZfwj9fcISjswyW8rdcphbO/5t+W7a53
dpB43vTm399mahVX4d78KSHkDZ+xTj93m8b+oRadN8sZzsBQoLsm3cxfv3PFoigg
WIUx7KujvZnkl9wTyatEUuG09xH+ZgqsdFeToEbkUuVGjBvJhTYG0hVKG3gZGpcR
gE5XX12uPU7E+piPGuKU8Uy/xLrvOCQPXiOS+FiAEFSU3KJQyDgagODcCvfpX7BR
4kjyE5nmpziouadjQXPggFC9bIqLq1kVYoKGytzOrvP/qlb3AHjBZVP2nqVxwCQl
n7wB+QYX80IKYT8iMh3a8g37e81JzqGtJt6JmjhiFjrGlNasfbSDmR/qfahYSS5N
6m0etadfMLpfJoBa2SEu94eC+B8XoSAUBDBu2xeGt5Z3MsHAt9MHV2lDjk1C3Myq
PtIXLygTzlTmz95lSj6nq3zgctRotQSHI+xReb9sCXqA/YUx6Sme11v7x3e5ro+6
lz5oBMT+ZhyrPaVU7bHn2jYwfaXHiRQSWCMAHMwD/Wu/qNiP8EIPJfbAD4qyLRl8
5x5/U3FsVr4Frhy6rv7cxNZe9zHG64owFgxwUltyoXZDiBlMkL/stBVyCHWyUAVN
gT4PX6OlqvkWigflVXb/F6c1J4YLfQcOH9jMxYhxmGVH0STE0oBc8rb/V4Wmd8tN
cpGc5IUBi75bdBszy6ZjaKkpvZQHch0B6GNGVBGclXMhU87SsKR7+c0BQx/8AXDJ
CFeAVIvDvTG5QMGP8P5x88pzF3uCsG0zAoEobwPIkgBjHMAaXiUzbbZg+cdlXDhW
TPztHQWx2YtBqI6Vm/zx6X5O8HcRUawEFc5lywvZIwKYVMU+zaB3oZfx/53c7sZD
UXeyyQZA9Yc4lqDKNJDh2k9mLvh3SaZrTXjK663iaclIuzzR1HWykCwYLQmTYNd+
L/M6XQanxItBHvKGl8hd4rp4vZvAq97ZuTQi1qmvOPvc/6xEEWNJ7opEiFSvC16j
IKOBIQFrzYs6OfZncJzLOWVurszOyCvrSORLerpIejI3BwyQItegUcloEIENoKqj
wIv8VRCHZ8BDl28YNmW7+7+/c3GdCmvGVAFBdACh9EPTRbdm6QrvwhKxqia0WydY
4OhjfmBowqUBYMksz9sqViY+rS8tF8U8dxDNSmavEqqkl/VEQrueW1TjP95p7auj
7vTMi0FxXueG/3p8U6fzQtvW4emtO+Yw1tU06V+HnHSjaPZu2QKvE1Q6dv7TCzZ9
oycUNA4ZiuljRsCeg1CBAJ8bldTrURf7NJebBnJSMr31+1tPwvhQ/lrAEVG97ps1
Q9451J+DgUhRmdy2sYH9cN1qFRExUdvJHQgPZM0oTCvxPOE2uQFRv0y2ECB/7aVF
YKCFx4WuWGm7WOY1HL8iJc5vPbl2I3tBenytg2qF3S6u4L73i7NZ1zvZJpRa3Df+
EkJofn21HvyCVFvfdqB9pv/2CleJAqVjgnmpp+xL00riTLDJ7CZMpLW3VOn0WQ6W
aU4frwwge8s99btS2cclE+5eOOcIkT5xdIhxQFbjxGHf4kSbHjT9l9E2usEadWpn
bEka2umXVGWCstKE1skuJMEcEGS+7Sq5PJBryaeRbNYYC0wdHN80LpzR3TdJ71tu
SS9vL6/CDuYiWMxlrHRvqy+Yxdvpqj1mVHJesYV15IEWiQvylS2G9K5HIQxpNLPf
TC7e+mojr7ty1XeRwsTvU1p9WaoyQ5f/prIW9w1d7L8OLvKsG6iICnxQY9H8EdYQ
liEtHHxM0K3160QOiHZ5slT8WCnrvPNmC6bpVbJV+FIv+B4UMngnyTbPpTjFd4eL
7a5CfRTD21o/SIIkDfiINccfLAbOGSzU/ys0Xd8IohY9XiEwyuuLgLL8Nfo6ADt0
GFnfJjC4OILtzWnz0wbc6HTvwltczzJ6Vab7VKLPn4adY4JqkRACyfVp1YaeznTs
lMPKH1mtp7wqpGYuSHK8116mzg6IBaBXX7W3Xw0x8VzwBOB9VTMqZuXugdSF5UnZ
2zKmyS4mksvhsAHfIf/p3xaB89RFEd6/w/xSaQW7GrNc5wYOp4qepSJ41xEGoDa3
ughfIgR8KAZyf4DsmlNu21UddxuyrVPbHOJRlrnru+klquSKxKzQKfPmpeSLyFtI
Mo95l1l+m0GXueX6C8zw65QI0Y3+3Fg+ZbuQqfwn7drKaUXd23WEtfwP/JNmMZUL
geD2SUqnU9ER/pzlZStU4XrJcQMhRYV+HQxias3n/hFMTuEzNQbmjQogNoTr3/o+
57eqcylb6tGm8BXBvTCulM3bj9/aLYE9HYiENmNSL/dZwEPTHLRUZNV3emTMiLP2
Db012PS4WkSPVZVF4nxcFCx8pVJEOSsKzYlR4ofHSXIW5dR1vYL/0MIndygdJ9Jf
09sR324ykv59bz+kpFk55vM/QHv81I2PFRoT2lZtfi4zmSEZJOR+i0/1hIVFsBml
qRC8z0VeVLWMJB40/yaArt+cjKNnGNP7+qSejpR/YoniGAUCX8IcihLHfcRLK1aA
10Mnt4kwQjPBg8kZNpSUTGkm5FUqmsjgt2bZHvZOwt/IF+nPcQzNEMLfEi2h/zeb
enMt4qkFf3AyEa6m8GKrI1ZDaMR7rvOu+JPI3pHPwmOsapKa9JkNVEJ1I4UVhwuJ
dzNyyAy0Lh1o+jEtgpy6QYusekc+T/ghd4QWGcmeC0tx2MG/Rsl98iflDBsoef4E
RSXmh0kX+t+KdNZy4eV0vFWnQbEGpPMOK5qkFBajxLp7dg/IkGAuLOo1bQU+JkuU
1vAF9Ehbj8rYqpCW/QfxZ6T8kjs/CLNXX0rs1T4trIQX2h4kdU5oEH39IejTwNCJ
5WbvWWBdNGBFGxycGCM9MUwTDqaKgOHq2UwG32KVE+7An2JLmrbAMcLgatj77Hl1
gc8MMeHIDa24jCFEn0kme63V29gq98EtbUB6ZwYWrynGPwTWpucW96/xl0OI85TD
BUBTg++qJf6U1Xsadn9jUajF87Naj/fRAJsvBF1k9iy7fNj0B/OmrzZyYmQbp/Lq
bY6Ovnm95Vr9jGafiPd2x5HFmdTLIB4g7sdt4WWWWDaquHKOdSDeiy61b0Okz5ii
9uY8vAo25JD6bJgU2kZE8z+p+J4rGcfGlpVNmiDwipiv2nvd4wfKg58cvxbh1KAd
GgTrW3NEd9pLn2x4b2YCOaC583otJmxdIN5c6Pb4DkKEivlTLDlPQs+KTjgeD4Ml
DhUpQvwvRcgC0qm2dzhroiHlueG5N02AkiEYiQ3XFoiRrzjxl6IZd0LMJVCfrvdB
AlpnC1+rDboPE3FajQj7mX36RBXPlVO8vYDWgB2xTSHVxWnPeKqLw/eOFLypS3e5
xVxCZx30WNPlRGUNFcGm/LwE/nRKZeJFK3AgafGK1IQB/r/PE3FEseuRdSjM/N80
axHoTbGFfzc8dGAK8nvSD3yLEg7Duwk41drIY765tgPMAE6Ys3dwxL5dATtqNLMV
34fVrcloErqTl1puIqkOIGHMTBMtEpNHgYtnlHZuQ/ZGe0smwbemfeMgvd4icyXF
ihFH5RZ/VSH8BlWd4Zu+EhPa/twVl7Xmdg3VT6GhXJD+Ql+GfzJ6IG5LKkd1wdCS
VlCMqD6/ET3N8EBIL7w328em/pHSVVN2DCp3tdkz55RpLhLzxD0IlwvMsXX39Z5G
4jdTBAq78x1clnOXx5711rpPF/f6kB+JFAQ/cva1jMPGM0taHt5GkFPtsffN9a8V
RCT1msyTl9eaVGKADuCotWqkhYo3oh7vwWy/uZQ9FtGjFzkLujJceDS3TuVvCbwE
z69v5vFcOsC/tAYRd/F9bm9HLc7vZDWNmUG29W60q0XMdgqsg67bkoRfRPRYl+qg
JFqscKmIiTCk2cox4PVKQ03BfsfA0dCeZZOlro1+XSYwE9jlMtpbGkv+2i6I0m7m
VLSi00braR3si0ftcLayQjrA5IjBhrZaQT1U26xJbDzIE7FmArrO3DknbYKyfyCH
ouRGremBfrYYn5xVLVelmVlw77Kejlh/bVd+JubGj7cgG+2Fp7MOnjKwBq9Ok40U
Pfs8ROoeUkd0XD7FyY0DYtlWjrjkAZDG2ut6e6pGX1oO6OXm5GGlrJRkY9I4eFwa
YssA1vy/31EUJmk9PfW2AfDDw4SomchBCO8cuJwdNJL+GUptZZulsueus2Q9clrf
E+sJyBixV2gHG+jKszqFtXv48DbwNbQu4z4HaecA6mTDxKJOKlAnSoJtNRs9SILx
IFco3O1Ck+DTVnGWeLWSROg66KA0Sgzw43P9KcRtBEkAXa9NT00sNagvjDaHU8n4
+55Xlbxz899nKlNxWBlJQb537sYtNE46eW7fvlBlx409BcTw+xeVuXHbRFljAcck
zBRaBftqVizkf9ENtnDfZ+5WtMNxj4vHeqa/iKBwsV04KYFekujQpMHixnHYOZJD
ykzsWI3HPJkkR4xaGpiVr8nXN4LsuuCiWzz4dvr1aS09pVKhWWbF3yFJ73uCQ331
na+V+YdROHeKdvZN+ODiO2+GmxwnFlafmpIFcTwtkR0R21gwC5fvLMXB0Kfb3S5B
z7DLZ+VtgSDi4Ab1LM8E938sTrE4hsjRBDzCsxDtUaK4h02geAhrH1TICMv+8A86
rFp2vdvBnE2Zf9Tz0oKlsSmaCSKXPfJh3RSvUxDFAIyXMPup/pfthFK8uMbWvVn0
mlKjixCoTb7s77A5nMEdEC4HY0ctS9iye7rVssgFBcO/hkN/vOvFGcJj3njCZ3Mo
p5TGWYXc2QJ+ptDocrCgqnWNGeB9TtYLyL1WYVTptkd27po6CvKE3FIGg7kiM6lv
Qm1Vk2gOjlW2QehlVmarhk/DR8DAkbX1hqgrr0CxyVC3dvRsSn37G9hQ9r9Jrkdm
X0in7Z1+vTzh0Q+xo+cqCqA23kVOAQ40IxhCeWwqHYa7Wa61UJBjtRy5gCcuFwHA
vfSD/lY3FuDdFgNbyqNZafFd6gANHYSZ/GmCf1SRD5KrRuKyr6fH/bNoYXZdltis
PulRB9EX8RHf+FmyfcL086GObSGs6XfgeXwz9HS8GtxbzVOWQZJpH1+beoj8W7pY
rIxuWtdyGh2kq4F2/AY7LMGv8lzwi+2qeB7XcHttxnK4FuUGHYF4AD0Yq9PByygK
IFbEuTQAYVbP9y6421F5SnaNkOxSgHfCInb5s8aJ5giPYkXUJVK1/ugnyg0IwZ4M
zjNrtqzukgEqUvqrCgUH87+FIrV/CQqCUYSxL59cgG5EhDVsqTn+ksdEh28EIyit
DwCSSVERTUCbIUmN6xa07LsrA5i55VS7v5dgfMeXmhR4a0dgjf7N4V1uFoZA0tRh
Gdg5krtSHugHzZV8ndiUEOeXMe1jXH1R9zvNEW0Ea3Bv4hTGNlaQFv3/5VfQ1+dE
e1/NOg66mJ7DRNVT5Gc9f28XsL4vhf7+JxdiWnzMOmTC+1Cey1q7MGsoOL5fA1E1
1lcGt3TTcqfWCSwyocVVjAZ3v8F89IRTg29LhwTEIK6t2rTvBwmUiro67IAzbfbb
HrrjOJiUmxZYOWf46DzskYJt2Jyxv6FP4HWFFQ83KzqJL2A6g4HlUlXiXCWcPqKa
1k4xvg9FnyouhHX+L3jzbx+pw72SNQ+weA/s+b8kwOsOIC1+2xM0rCad5CF5vz6o
sL7Sh+uRDO465UYBhxQCtTHrBireopgLktEZEs0kJSCBCcegWXr1Jk+knYhurqUT
L+oP8CZNad+Qov64DcHQK694gpQ5SUtOl8gDH99CbzG1xeRljCljjOwl6ygVmFx3
essT5xQH7rDyJgwDILFF3KLGMYz+xgE3wMK9GhVU2Q2DnEPuMO5B7Vw+RGEiWlDi
FOY4eirIOUpv4zqNVCGB8Q+qfyraYJlK1APj15ocpnuxsbxYdvxxStyeditAz9gW
mA7mizOVjUvE8K/UydwESX5C9rtzSQP/HrG4lkaIBHe6Tji4a2cEuvCxAfYu/Rbc
6oFiI+Sz45jNyRdGeSc/D0pMOPhQkK0WWEAGuHtnmd9vFEQUdgCUDua42ON8M0Uv
NwNbfVPuRcOI9yk7nt6WSr6d7Fz4kQLmg40OASo+vLmC+HSj6AckSXo3C+W8cFg8
6BDI41Jb2SybVcEWzptkiPCpW5HJ58lhedTdeIxQlLDywBx41jU9HaaukDxLf/9s
RaLQRalkvFuY+xQRW1WIrErHuCfOwykDP45aj0Wonz8PKc2lyMqXyknpUjZtyVkn
UCfmkKNXVpEtXZ8hdxjbny884FyJ3vJGZNM4XHmL7vuROcD8KcuaSLCaTF+CCJMV
gABalwdawhOVDa0jNDBaFdhhfqd7TPKEpQxglC6NN/I/jPdRwPyniY5IvcE5BT8z
sI1gm+SfWkpJpjHBmS6sSAr1MW5lfa6K+w2B/1Jh/lRx09cOg+lSa7UZHNeLfVGV
R38904t2QTnBI9T89WwK4DEjpLbJORyGbrbcFpEPOUDpby1HJZKuoFit52rf9bFv
rCMffH5GhCL5sB/AjeiAF4Nzgu+lr/2N4SvdsthJmcUp7g4AnHLTqF328MK7jP/A
peDJRXSFxVoWHIqhmd0wtQUeOReTJIrXfgfGGGc3UB6tI+rwgcZGcmeHEOmAtFPx
J5DsN117p3fpDuODmr+7rce2IMvtsalARg6LlsMEMjF0aNV18PzurYIBkksBnN1G
XRWsK2Tj5xIrYKWXcgkR5aPBRK+CN3rhAvx3/nd0wfv3NeV6tB39vTU+iWNqsexp
NxFqYPqv4rr3Qbh0OsadbIHH3h5Zr9ZT/ldKSRn9/scAhepSmhjqPvYu42IQqZUi
ATM+d5XjOXz6btmEjk9no2hjVEf0F5wt9RIYLPcrzXHlVJz2/aD9pST0PbkcvSft
kBJiDSsVTfQ/imRG7dt7tASj7Lmmoy9LIjktNYrXNpGF5JzWMvRLr9r5z2eBBgh9
64ICdUhEWFESx9eUR1qQhFVm5Bgosreuhf9XpDFrCClNpT3I/re2e4n6NVfL1LL+
7uBbMXlj5XUxPrrywarQfs/YjVj6ux0cQ6tn4CW9OcK0ghD4wVPzLc1CwRNuZGAG
AQhQPhOQCEa7MPt037syM4KOruHod9PeQu70lxrf8wirVisSpvJ5Iay0/2x92yuw
Oc+2WYlI4WpvbObTLChiWnAqY2aB0ysrYGlgnnGgGe75krHB5tRZ6x9DZp67xX0y
6zF4PQ1v4pQ6n3JYF+YUutiFxlzB5KlB7yiFAQXgNnKOESnDZ7whc7W6Qr/q7/1T
zXVM9LWWcu8p7l+sZdog5u1YwU601mSOmLog57W3u5AuEjc+S/I4hq0dazbMcA2g
OVC4txO9mKeZAg6bghY1zxIH7I4gA3QpsHCjxXvHXn4DeeBwpibGfJp2NNJ+yMnE
1wq6YF/Ciih1LgaQy9oHBRHe25WKkHfU9m5mOn0Ny6HdXpQ775ZvTnnWVZ/MrciZ
XyQpL92jiZEJLhj0wF53JV9t8rFo17pO+z02WPK2nNkh/xPK0pkzvQTaHHWMhhWQ
y8teJEIQoR9OHiEqp5iVm2PqsjyHibqsDk5jxoB7kmIjCO0OYMO8STW3K4Z0Ys0p
OzwYa8m1RT8EEfRPmQ8TzZKu0/sZlpfSxaawvaSAaqc1hMZjacJqc1rx+ABO0uV2
BFKEFM/9i5XVj0iEQ7WFYjuB2a/uq7Jkzn6HS7O5IhPgbQzmGC79oyoAYJOZtrtm
KeRS5ZWRMN4Mapnd5JQ8kN0ktIV/B1wLbt1G+115EJ/6FTWoyPxIHMPDlUSZjW9K
IjPXdaU4t4N9voE9VUVjmDINDlHREXW3u237zkjxZ6BU2uIWJToDkIhylJNgWvOM
6AdJnqTX0ZmiTTTuwZzmMm1jJl4LSldFAKf0NCAI3XHpcU5ugM4pl0PQS/2aD8KR
atcWeKbx5/KhV2jArdtwz9tZpPs5LISr6XSYZ7hTpjwnA7Ut+MJfksUGlPBCKl8E
i03O7r5352XV35nUu6mBuVjZWZdvEo5lgmNVgJ3Oy3EAZj/3mhMwJEkMsEGKAvio
IgmLBnWEOxNY3epe3nXShSZIXxqEsggqkro+WhRwb2uXhb7uv7/Wap+1/he2j55Y
zZ+CQkboLiR79LUqXLAQ5EYoTa3IYFy7iJB/uhZShqbkJC+5FumojuJYpUcXRPq8
D3PHNIxjy+e55enHKMfDIYlRm+rUNrjwU/nidZw2LvnfweQPN55icoYGFPs6Cn71
+pGz5efKODsYQQHjCwL+/YIUeNliEgL2wqWIm3RfTkuovRBQH5qviY7dTyD2LxFv
cBpEJdSmcc0PRKtNEZm+4phzrRgyd8/0pPksDFDeAL1lNJiyIpFTlyENFG70c7w3
PNAfpF2+OrtGDbhe6Yz/y1ybzCW6vnZ+DGdX5GavKSPfap5ZTmP8diQ7yZtpAktm
fdRzP9U9mGApD7LnjpB10we3MFyAgrpT4IMrCNpThWeEKOQGIcDoyaVF9jNzwZ2Y
3Kiabft+WVXXFowfP0pdBVrwCcCXvBNFtYKPGFDraIce2zXZuRYpfT0neTvjaVBV
uNOsPv/gNlROvCI2Wk+zEYSwuI20rEMEce0ShwPIMtYManToT6zIlblcEVhUesSX
tHQ4v5p/aagkkajcDy2LVfrylBL8SwR1yxmNEk02h5swacyQdkijGLPRPDunAE6u
G+QSp4XK701jPSrMKu6ZXuyUaYxF6eBfNCTSMSTOU3W8XBsVvPpk/edBdhRbu2/I
M3Q5fJhffL3Dr4crA4aGX+DzOVPqyJ2hxrv+tnWpnj3xjq2U6L+CCHWEUG+GlTWE
F42QKXDBD3bU6Ieaz2irMHBFHq7QjzauHBxOVy1UP0qkyGP49C7QHqlobAhzJhjZ
Z7of4qaAOnxLDmmY/O+bcir4eq2iniT+wlHW/fw9wwgHvAnT7AoJh0MuvJvqs8rA
HbLZlf+oDu103H8B7kwKOnT+Sb9Eq2ThA0I1uPX3Mtykn8d9o+Ngu3e7UkPjajJN
6bg2XtrLJ8/Ru3pmE0HOAVhP7b7YH3pbi5SbcnDUQkR0dmtT1Hmrgwqp+stNv/F/
GEJg95D9MrrYeBqvgaKJGIr6qHAqk8E++3dfeudcg6J/4TnE3HYZowufDaQONSXP
mvMJhTHrEtE7VWMuRJUmIJetfr7N8zmhPtZanXk2c8CyB9ka8uUNL8AcUO4rr+un
dFJA9Qgc9AN7JUpNmIPHxV1v4ZU3l0rii60dOrP38TjkrijPNZ9mdAHlE0MtczuB
zuCf0HKoSyPgMy9TYxqV+qG6h7drFDOcwqWAsrDZMBU/+RU0t/L2KgDkxkf1nr5C
IsWwCf1owui8+UDonJ062u1JWkMpTyzUIULd8owigIxTHQDC10wBncJWdKnQwesa
pfcyFYJgm9Zxtz1+/lG1BDMCX92yXoucsUIo89ken33HMCTXamUgKNU0LStm4rTf
JmCzXeustKBP7JyvBZ0kRSzROHOls03pdAgGrDEjefL2BbZ4GMdrBMTQWUuI9rKt
uvHZz3M3xzxtulYwk7wE7VeVOB8whs6mv+uaNsuAq7XQcu3dtaV1yZLdzEEJFPxq
ZGdscO3DiU7tK+7XwvIOFbIoIlSyB3HlH335WZMUdW/e6FjcWsRxdlw1QonaBiaE
OXHnc8K+RkK6PrVl0wIwrb3pdadUud3lwhN9LJwmDYQRgYfscj0oNwoylzX+2S6O
iQdCB52aMZMYrBVGJb11TvRr+4jLbYdschWsib0W6tFaCD3QE/Btl2Q0FOuyb4dd
lKpeRU935MJvseXtF4EmGV0cqgVP+wBUXF//lwwHjpZiB5xT65bjiZDp0hv8spzd
IbInLOzQ/titiImgkXqeLya3cYho975wkT2zJB2VVEVXq0o8kFGbEL4zNTlZ/1Kb
QShgoyY39y+9DxHJrWzq2EDI7ngC+E75I6qrVpcxzU++6vJEQVlxEeZo4lgIYmBJ
G6fjrB0ftKiIxCKCBYc5hWG2a1mBDgs0Mo8DXeFKcpApboFU04GmShHK7Hz1Ck1l
0RVxPiJBO53mb7XUVRBTfrySoDJLf6YFb43qyZUq7S0biJvq87C02ZlktMBIvrm/
Ep465JgI4rRQo0dTBxFuGNbTOB7mAzsDa+OkxPC1RmfjjC5/CmxME4No1+DoK0Kg
TmxhOhs30YG/Ovw3DM53GVj4rOJQ15eQu7nMZJvtjsYlRyPbK5paUMo7bSXaboG2
CNPZpQVXfI78Wa9ZnIGgLPgloAj8GtqZPz1BhoHrzpnran/Tyy87tjoV0lzLee/h
DGvyNeshe8OvCbMIw8tzNyrrruI9RmsV/F7XuAVfO1/bgiFMii61D4bkjRC1ePPE
FT9yzC2e+qW8pHEie/zwinFYWmPi48CrNMg5d+eeCk5YKvU3zNoryA/xjRBNbicE
CD8WEkb+Kp76Q/qHTNAPhmeyWye8hqLByxIH6iZGBCNYlt84xv93k1NwP+FOYcr4
yOHIAIzf4aAGX0juG+R32+0M00y8Hhh/4Dm16336lfcTeNiBf9ea63hVrJvVNoio
WY76K1uybDTes3crmB60pV4zxhmusOFpQon2o+RF4HUgYOfEr1sn3kvtf00LbH3B
od0WqdSK2GM+Edtyh0ZdXTQlg6Apzh7Vn5LYtFcj58xWot99+FdvQLC3Nnb/kr1h
T1wmdUc36rt7dw3+1ahCraT5r1mgby+FBofny2eOTG4glu/uFLoIbXfIUGPRrOi3
7Lxa0ElN/HlWbQmGx9quyeLasHmO6/FtE4S8u5r2UeBz75rmevdG1UbvkeavPI6n
wuce9CSmWBkiv5kATwvM5R/pbRMtEZXiuNMxwS43xUxjIKe8KJlrNFrtazI4/voR
axqKyVCB5qSBK8bgNhJQm8k2zA/BKaFPrJ8UO9DVhtkIUxy28G+xVQWMLu+4E3F7
gg5SLLLjFDAfHIoTevr/Rz/y+akbD5f2UKh63LIAhpaagQRdw9BlXbZQ1eoi0f8m
AbBHRUIMt/t7jZ6+p4Uh0fW3o1LO9eqvSU4epnVsYhTaAwc4uNfo3sVQKgfi4KqK
fw8YInAtjLjPipGkg7hUDqZLqplqBmKPLw0Ng1eMUHQSD+nbCq0zLasYZsJ8J50c
j66e/GoL6GoNNEHFI+yiSo2kvYsochk6sNcYAxgu4jUg6Fb3F/RIRqFDpaWnDF0A
HnhyMXviXHrlcXTWbA9Ew52Xud5fP5UM4YA3RkklYk0vxLdFoDfeo1biUl0UNUTf
aeTNMwRqgPpEK6BKyCXrqKWrZSjAGVr24LLG5l4xvaiNAwMfPIM8AHqDZgge18du
cDnrp9GQGd3GlR7hJ7gQfWxLb3phdGcl5HGthP3kiZNPqPt2f5X0j6aSaHVXR/s7
/FF+GA0G6v12o+2WFwZnyFRXGHeLe8X6xvY2twimVppi4pLzaf55fZzQK+DVsz6V
L3awdEnhXmjk6B5IO12TuesI4nwZvGLT1vdokpDELAWQu8lpacvGrzxAMq7xK8eV
Yr8yX2GTuPHt6K1Zx1zVAIx605MeU3VjV4TBsBhJryWkRMFqg6PoR1oAR9MjZ4GN
9BEhc+ifqfdLBIW4R1lTXYKQ4r6vN9mVH454fpq1BWd2iX/c0tb32IFVFlxdXY3i
fn3rBY/XY4BqZjNm94Dfqb6eHN6bCvIPycoSQ8B9/fm0j6OXlO9k2cpLy2xADNcS
oNDhzt7rrhg/a/A5DPgQyjklK3QTngYiO0y3LKZ259Uo08y7N6Z3ycalfouVUZsq
SSWbGhx9cr5Dr0Uz5LGwPKYOgRav7DgZqQjT33MfzJsmGfirquDEXZYaSPAKicUL
LHaBBr9k8+bj6LvtntzavwUIT15xyVFqrX4F8E0ovwegX4/vAnhpSZWgiz5IIiul
HksQR0PpFGOOT0y1W5qtErFRJsaeauGPqoWdXXyDY2uYeYhXYJSveGe3wDXReBol
W+FVK7KlG5N2gOUNLbs9NBARNWNmS7hnrxUBycSMjG/DAGu+tiD/Jcq5rIa2oZEH
GlHIikWuKXNgHXoBNtjiOH1SyQf3+6is0oDrZUThfcSNcZ4ns4jz19Omlzl6eMUO
8j9lGXTgkC7MMrCJBM2fHjFolxC+KkQXqqxHMHu0UprlHRYG869v0MNpbqzLkkB/
fvuqy9Dku6wqLAAqbHiH+rU5VxvXfCHcnsVGxMkpeAPz1TgM3Oai/L04LJVfJszW
63uNILphk+k9Kx0vbNGor42SH391Z/nnx7N1G/xy6OtByr/vl8rMawqAMHht5Fpa
FGWcp4HFgn8ytgP+G/2/aYMi3W8aZh5ICITNTbefsgLEVubeIpUpem93PDAXd2OV
ikw5T8HivHUG/EX83N+36s17stxEvXncGvQHiHp1MrdOjMfFxpoHbEHZ/dmbJzhX
JBXyTt3sTAbNwtsFRzx73t4mICtaUEsjKrD0kw3iDdLP+S9KOqRwiTx+UoXs4QCK
7l6Fl5fQmHN2cJGjUMV2eMxHr5NvcY1O5vfAL/gfXqfrCw83hU/wuK/lREGveadh
cpzChTk9wzuk5FCISSMCoFo7xTbER4T7RXBstmU+Kae7GfrKIWkcMNqXsHcV6GGq
iFvJTTUnpQdj/OWtYM5L4ZQghCGOhjqZYbRBHtgcJcyGfFO/+Ofke9UqHNSpbT2m
4ruUh1nYG+4Hp/IGG4k5FzbDqA9EkgD8yylIMS+cmE8Z+S7jZ2iPLuEqaXvhg+Ra
AvrPuraW/I0tjS/nKx/CQjpRbRGs8/gMQbYuel1sLoRKqMKqfkw0vwUUOLjqRNVK
uQjnqG4tq8Pwx+VE35kqEmed4Q3qSrHGton0Mnh3U45jQXssJciY4dn5MSCxB4QZ
/jquU+qqHuRiYdeaw2z9b/mHE+FfziydRNz/LMBsp+c+mUc16c6gatBVo1vUXK2+
e+mYcGgj90AksaQKh7NwXm7TYPw8Y7lrQ9FgxJLpfToExwcdkRp93S7AXFF0kijc
70zJvZSoa/l0Fb1l7z5VkVkb4yperYsUwm6uwJ9pypWkf+ZPQsqZHybQWP5sU83X
UqxKy9fk3aVdbxRMGxB5KM60vcvwnxiqpESAm1D5v7qFdLC7/gh2grB3XNTmCaZ/
Q2gKYPN0MVmOXUqQRuoWG6zTs5MjUG2MSD5qolnwsFrHwJ+Oi3tvWKZFq0b5Hdf2
YOg6w38SwoJUm4i3sxtn1bR1Z947XLEqjMerKwGTmWaMvQU8i678NBYBK+8qJeOs
Z4o5LfdOnBMZ7vROD5fxgjRhIBxnXfMFBnOjofhUHbUVmTK2LrXle7jJgysnLmCd
/aQ2AmmrFf9qUD9QBPpDei6H6PGFgW16eq+nwCGFom8lezqa3T8S4p+OayvIrLwM
94blZIh3QEwjQf1cvDfvDMQr0VjdVobJWMx7wQfYv54HQVRII6h5nijnd6SSXofW
F+m4i3V7oxAMb5qNKf7tnY/yKSPnIky1vgHiA1C4sbEdt5V4dKz0a//eKpTob64l
iJc53woEYxm0X/1tIuDETdJkFdwEro/cpxh9oHLTsxT8PM6bk0usrxvvDl+2Otqo
1fMpMsgRDorTzfddqZxRPPeuXwRwr8yGMJfh3U1B3X5la1XBkhEPhjIrcBjcsQSq
C6SEPJ1f3f0BSpwmwzHFVxI/F/usL7j0AQZQFG3gl6CDrNQPzt7vPFqZ2jrOkIFe
5ulO7nOTOWKNqjl7JOewhKfV9ysBsvE2a3hD0z0ButrbozSCgI45XjvSPqaC1sVM
IRNADHtguCRjvK2jIOepj5eG21iM7c9ggC0wp7qI0Sv8EplcOmR/LPl0iG/pjZ+5
AeXZyP/iJOdzlmM4NMhkjfLwtLyt0eZl1s30Gy1BNl7+1ZeAXBFQYlUMqcTQfHcY
g18Uu06X49qxl/7RleV4bhaMUpGwmzE9SbpqxmQhO1YThofUqCT60MwTJWrL+TQ2
kGG35F/7oXZGDto4vTtWvaqORMftcGDqwNaX3DWqmr1Vc44V0O/nUNm62j7eWtBp
XZpmDy19rXlM4FzNyFdOg/OKY7IIBplf8ZWOireqIE9u0kGA8fyFe2F+33xuEicM
jti6MGjCtTAe3w/2w8yWsTYDwEq2Q0KkQYTb10v0is76QdIjTmdCDzz+kQxuXiw3
5q5KzxarI3kurRxHu98wk1AKn7bsUroROnuLuMB11uywxqyhKZcPhV5/Hk3QzaJj
AldRV24ZcGcKL2ocEJf+/E9tYIObQlfX2Eka+z5v4ReID+xbS9vikdvx/jPx682B
MYVi8riL3VTlCXVVevP+Nw+uUd0hukQoRdchThEFKcCf84T1j5N3N4yZzAPHe3A3
PwI3LlCZHQwb0+CT4vsds2YsHw3i2p+H+IrG8pCuXPNfHzF5sh+ZpY6e/RHoP6g3
PeKZXY+3CS483Mdbq0L7XmcM0jT7LZuevmoGiwf8vSig6UbDeoR3ol/OMuR0+BJj
pz0EcY8qFP5RG7Lg5nFutKzPZRvp+g4mCBPBaWHIHHY3orixHu56rhVJHp0WohuN
wmzQar3duwEZRBrb6r6r0Z0gbzKGJOvbig9UMXReqTx5Ii2LcfjnA3Lfu2/y2m1K
BQ/RWm9CgjyeFQScREEcgealxEK/pCUGbhob53QZGlvEpRnrJYAVvxKECX6SB7PE
kMsiiUqPBPk/WjSexc1jwrcWhyeZkjlQgWOdp0mG384R7O2tyjSnmIxRb0deVYnw
GnYPsauYy9Unu73VQ3WdD+LblP9V/mKKhJmQI4MiO9F4rJjyMxAIUMY0hFekVhDP
FYLYzTubXRddxw6kR8wk1rj+mjwfUsft8H0d6LBabRYV2oRC4o2gTc6fJxd9TXDj
2ETklV6gefwPzwNdnThuxkutju4vxVhYqp7Cz2bIcJ14/JcQsuecDdxf39O9mlnI
Gv0pvV2d4m82ys4Qyj4bitjJiooDMO4n6spNwYXWWmObro0lKYB0GqYUXdV8kmM1
lDzNmTSrS28pa4gu27HLz/gvTJrj8W9m7PhE/BKKKZI0XEz2yQsJZjM85KJnjDfR
WPRJF7Fx9ei0XPWdiz96/IdHoNaLgjVNKakuZsxwdy3hTMAzqrvrvAllHpZm7zGl
agvMzVOwFUwycdrUG79QQ5zY4ewoRtGtuE9BkO7eHiNiUKrbacWGhm9W7W9Udv6u
U19Io1KULoK1M8pODsRh95+likKMs7hY3FSvTYeL5gRXDjye/UAd9OZTkCTNI0oO
Yt1a+aT1JXg1uegP+Oo5DIecLsImfoAhxqs9X3jKxb66GfbR6Ahc/D+mE8NrQB14
ZwIkjWBvvUCc4P2jCH34VtrJGI43ZruCh72acu4bVbKGgNDqQcUEI9uiDOMY03vb
FGrOi6KTaFnsbsdS2uWxCWmmNLIU4W5k7bW9Q3Qm/jECQ13EjckHT4VTsc+lobh9
gRGObCovn98ou7UwH4MdbVD8J7GSMmjJXZwoZA2eTMUxxkfImUuyDwyagCq52YfW
dLQ7L7MFa4gemzqakGrTqmWrue1BtAgxkjQ59ICWpI+1VsxB4vckmBrmKH0Rrq/n
HPr4Pycb/AurHTQZ/wpspns2zslyg99+WeQO72VqS7OUranBaUtwWLK6gQ4T1CpP
ZG0dIDcwKk4qnZsdltjkHCzrVnl2Y9xJtQMiGrNWHc1smwyH/qMxiR5wbqmK289M
WDssx+IopwOnV3Ic8a9IjD/f/Vhp1xyXHBIWea6/85u6Fl9YkE1OkqMB6mr/NNam
Mb+IIUcx5uaBOAnadOIbqhEK214/ukuteQYPIaX7sRMdmYKg9uHyauudhZIvlQ5s
6I+5dg413R4AsJCbl7V+EiBTwuNK40x+yceGOhwbOCVdt53NaXnFk62YflnMjVTT
UVv2teuo9kUlstUrp/ww9fNa5TLVgQ+9HhP0I/7hMV7l14OtbbHUojUDsIZ2skg/
fvmxqzIO2b4tPk7ESkusRASbfcuQEnKlU/X5qJ7baJsM0pH0dR2rb18FnbIods9+
Cpqn2lIRF7/3OAsHVjF+0QPhHc9FRegcRm8nXqp4YbQosFXgsjWnAosN9aY1BCYT
TpbnZPeIxL+sypPGPG47V890y1yrxjaCNvMJjTzw/8kj/dwxHBRHGDLEWlPu59V+
uNznOV7WtKWVyRVb3/V9lpCKT6XUar8Zcdu87akN+08p046evE7lQ+CFRB1QDIyh
AlvP77pNIj6t2L8zbhBW7dcUHHuu7HlmKGrdoxA4kEl+kguplyrqiBt8GqcXZaAJ
TGGZKN2Wx2qvru15hmRL+Cp/Ut+hFZbHsxmKYMmiaQCtSPscBEPjvQ+z8LciItA+
HC0hkFUa6q2JNUBQHyPIl+kK2NioDGISG1igEyCbE/v08Lax1rXFZ3lTdobCqteO
BRn3NQ5BafVmuxFKqPkzHzoANfuoD0//GTE9W4qr5f6+2nOCxUMnHYe7rqBSHDPw
97WT0uP2V5giy9N9kJJL3yNs1r1BlfVDOEO8oWSsr7bQU45ni1Bk3TW8XbvvxeB4
43KPonBLLGqCuyZr1J/l5O1GqtTkpyyu9EUq163yvvfu126h+c3UoEdW3Dj6kcp8
pW1crzNH/ApGvSFs7uq97Mpb1hg2aQZkT1ULbyW3lGPvaRmwemDqMSL1i2+CE6DS
Oa/L39i+QeWNE2Cpc9MQQzZQ320/hxp3SCIRrvVImOfamxl6ncZdu7XIUPy8R+Rb
rzhVnv3qjC1Y/3WC5kRLGjWq9jaN2tOAoO+LqQahAX/Cg1q8SGeSINxPr6TyzYAE
UT0uhrA4IZfan4PjZDjXICcAiVQErHfzlOFvwhxe6o8O4gMENViy0baKlJA64694
9iqkBkxP9p706y/KBdcRCmqXRsoF3hVTpPaf4IYRuzuOsZy2kIh6pX8ARB2Fn+7r
vw1r+2864CD4sPvyDQpXG6m1LvgPlkitopiNcojTwXdAlO3+v5BbnI98KU2z9Ze9
OzFUC26dfSIlatGqxBzrhGE8Ac0SOukva0d7LvtWYm4opzBmPFMI0HN2IBHiyp4E
eHu08WQ1cS8pDVQ+ys5gvSoHEZWfEgqVhTkyH99dFb2pdckwk+YBFItbFPQrg0Es
W8PdQS7YahCZeBX2psdh4y6uOQnKNQuaQnbXoTSr42cdVKVfoCn1OEBhYh5KZNvZ
eOA3XoO0f7Gz0qhfePwSKk0AgQnuw5Wmq2UnofAe4+8HaZC53Dh2vhxGHHgT1qJJ
YxUfUJXWr6lc6LVN/BFqJGhvpItgzZyA8uWE734broy+CHppVWUKyFQCrO1peb+X
avhvqDoaGTuTuXyojqp5/rZRTWD12Y+5nsgIDyqxBh1Y6rxtOx0vDajlinmCAZhi
hPmzjj4Gchh6xIVpTk1oMJhMVQGxTVF+NuyrT3kW8OnVfXwe+VB7uokmu2ZMQdrT
yqeGWp2U0GJmvyIBo+vquouTzNeirP4KCpDGJZSY7ZRUaEiDRvd/j/G7+oeTgJwE
MEFOof6iuldfZKSbv/m9e8bHk8WHt4wPvh2PzGN82hY0Aktr1QbNYYauXjeVMBlu
bZgpPi4xRSIF0oxg/fuMS+wTmOxV1Uw0f2xC/5vE8Wr6f2qpxDYJHTZlI1wlJZF1
3SUdZiPk6KLFi82DOeloa+Lb6tY8hLLsz4v0sMMFrU7P5VkEvEwATHSGcqDdHD8n
4ga6noa9j0ycP9yaVXVvB/Cs1IeINbqWOR2s/xr1aLxM9rxLnaagOHHlqLTW2Vjm
Z8R6LxvNbFu3e++I2MocP7kWUNryWnrO9+X6IixGucZ/upBMIoZsOdzYw2xTX4qF
1fElxv7oTSDtAlVy+aVm8V++YVolXaNdQSybzHuEe/SdqLW6uhBY7pvgu47kE3w9
jH+KTdaeZrQjWAr05qQiQWDPlFM5UcXwjyt3DBAZJfeFEVUsMMZvKk1jncQZF4Vf
abjYkLIKlfJSzdlWygMs0niqGoHeR0y/S8+MlEQtvcR5F6RdvbMD1qU4lXmpkn0f
GZlgDAjezEAj109stdg2zOk8XWbA+mKAVlJcGTOrYddBfu0dq7jm5XXmw3LJdttj
qncR2RT3/P0xfg7cHXOmgDCOdrgH+HFxLYDmSEgdIDS3bqQHx5KuO8EnCX2yqkre
Q1SVrfNJAKDzQFUeLy1JLiXc+cecSRMs6KWul+v4OLLQJutbvFu4llmZ2y9CZ/TL
cfLpoviqu+oYCOfzCfwWLC2G0Li2dsCzfqzGX96Y/Szg8bTM9ol8zMH2oGxV5YrC
0lgF9RpvwWJ7gzOUcQtWo1jLDPYNcGLRPGwifph35YEwHXhnVeVEUPhNpcHMV1g0
B1LdkVSL18/FZyztyo12xiiIjXNbEdwvtKEERFGhyPwc8G8m1NPUDAyvW6lHTZ5+
hTjFIvQssCyd6cTu1ECLsb5+zD+5qVP5y3UbVdGD9g5hekb46qJbgULY3TqJusI8
d/xo0n8EIR+UX8Y8cEbhazPxAZDpG8J5mivYMBE+SLVaIR41uO9EE9TKGq46yhYh
iBtT+I5TjjT+u65EiFv5OKK0z/30u0w+vRcfp2xTctob4TlNxoPdUlO8h34ckzNU
o0/CP7KGnBTceM9nnFV4oE6MyqLdFbeqy9eAKFEMMOg+m7OlbpygCdbIdV16ZC6J
JRe+plS6e+NKEEbzS8QIs6l+45OF4OqpQkQE90ZscysjgfLVejRaPBoTdWU2+ayE
SyJq1Dm3Gx2qPeM3NAWOCIm9DeP710OfHyot3G1Lvt/8vc+XNiwVrdvH4jY4kG+E
K9aQZ/3/OQoG+n0Q/RaWvN32E+EcHE1C3vm+Ivd0j5YaUpoFZhkhcI3091xN10Y5
zuo5kZ6ZcO06WVn+Ok64Hf5NsOzCRurTf1sZ9i/hFCcOYnApAz4hOKGHTCn62cP0
zJZAT5HSptKkoO75MydeGmX0d9YoZEvDQIe/AbmZT/Ucqs91Wu7ZHEOd0L5STbw2
rNtqDNjgn57m6X0TbG/6XFjrhaKEfO7XqnJg28/GrLskpN47bTaBil3TLDEDxWQH
COAE+sOSimp6S/80tk2mIMpNlrJE1PANrEdqYNAfBWznbxkV06GLvoMI1sCvhYwl
on643R9ky1IQifCL6oAKElZB4vr+6EVnFsqBgNdXuhjlvaGEOtITumwAsbsrmTYI
HSgf0mZ7nTgG9w3ipP6E8zHr+uUwBP1q87NmquxBKtVUvYEnmkxJpylgIpaoI06e
7/x+DTAau9SIBggP1tsQd6dGTPDj5rZZ0aN1nU5D9AlYPLZbIs5QRnhUFmQJnURu
iCtZRmHadLyT5IXi820niOU4QVIRtqXynInEsoX/fkfIiND0tR9rat/fhKOJp2Ks
KbLzls7G4jQPovrkQDU6R9HmIhCIalBu3Hn5ATd+PbYwMjORsUr7E/qr/CQoZMPf
NcoblfQUdIt2/twPKMJuaPzkGF7efG4+RUZP4P/vcurHmL+567XApcd1xClZToio
mZVdMbyOpsZ/eVic78OzDYPQVH1VDjDLeksdYZpnTzmepcx6JCsM23+1IwvOujpo
w47GthJ1a1TUsnCnsHLlRr3xre80HtmKFbQv+MhBSnXsriOCOvHScnrIXAnpnfsr
ziwW4HyOaulu1RtgibspwPJ3jIpOF4FtIBujzAWaPFjtgQMiBeefq16zG20K1Vw8
0wZbU5Lf3jCwBxU1gzi1gXCkjtjCwG1qyuQUm3epYMVS9MrTcWkexjb6olL53S8y
1ldMpEdS18pnKbm543gB8hiBLqU/O3jjmJ7gpJHqcSJvgHn61gD2nUz2pLg0jaxP
OVl+xDjo1/t5kTW3OH8tQWafbVd1kv9gnKA+N13oemlaSJPQgfSbnEReg4zdRC51
E1yVVyaQeWUYN58oSpPhAbv2vrPLEHpk2FCr/XgFn2uLjqVjiNJdhT4SGTMYxX8x
XRItF8uVX8gfXWsq/zS4+ttA18LPIO5iKQxO8J82r6SiM3GKB3kHKqUFwKK9+cSU
ry6Q0zH1BE+6+0ZbVgeIjqCVFAPk6fiS0uGTh+eg53RIwltfGO81Qrbx0ppWlT4G
A/5y9OK7LnSGExrr2eIAFnbo4I/dNDNg8TTd3Ha0FoAtdcj6wk06wUjsfVEL9vcT
1IkfaopVVjNnIKgQiXk9HdFKH5fRlwcnla94W19h52+0+A+NzJWCX8eeNkb5IKzD
NfeWMziOC9p1MC8uYzpsLscSEJiZxEVR02IV4wBQsHqx2l25Ky/yGRX7MQNzhrvU
3Geua/6VeszMTg/7fli7H2Oy3zaKsHp7cUrooKB4MCF0idtp5BY/MC7tvDGrVsqV
1A3QO3qME3ueL21bD6fDet6LEVOkfplKraWwL34ah2hz4RfgjvILi8W7PVEhs3cC
YF5LX3lQ2EnZMk1lJwV5Xts/LLRNda6KKG8eT4cUJkO6dYmeP2qWAu0qvJ1jiPjP
IeqDmJqU4b64QAn2/BjDgkO+eo9TP3lmDsYWXM6/Vnvz7siZwaPpYUqO/x67l0q0
yZVTVWRtUzDs2lrIrk1hQlPq1r/3tLgzZmmdoA/RUBYldh69i17Go/TcWn+dOvdD
izy8dZLbz6YBQXffSMOYDUyHqrqXW2xM7dxvwwD2G8cdgNn/qOptNmkt50PM3sbb
0e7mwpLAdG2oZxEvHTqVJRVSKbsNk0igj/G/leMvrc8WyqCMsrX/B6ii6W5kl14N
S6nZaprTbqyC8rlvPfdt5BPmz1JsbzeKkwQlay3ZxtvfruYlzYvBJAM84i4GM7a6
QlnNrnOxV9zDuikk+LPhFphOXq7U9lPU+TME/tosAtA0lVYeQUWKf+pHQFCHOXnQ
pt9UCIyNHmfXSmRS7pMsOSUVV4bOCVzvNU3/D7iMIChVP7IPqDdW4XkjinM6mMTh
vS1+/k4sIR26vzVdeNcFG16vL/13lG5b6LtDY9ARMYylWfCdqxcJliuOWrvier3G
s3B7t5zRKMy4kTITiGZmVkusTF6b8V1l/cU0Rsat2IxmAeMM9zJaCtbjJ96o3v+b
yKBIazm5BUdJqmhKOh2RUGuqWcG7LjKHy9RGI5pBikkjoLiSCzVd+tH1XQNXNVkw
N9PwLgWJSwHJDzoc5Y8Mnoj03vLG2DQjQZe1Xy3qp7t9oBCSPdYIxNHf3nWV9scq
EmEuUfi0oGBPKClIHp7sJkLQL2fMTZEyG3/3AGO3ewJxzV/e1A7DF0Ib5D2PMgfP
m7kTdmQh88mSYpNt73rTMF0Dz1OGpJR/ODlP6fwZs8dlYNnwng0b3rPunF5W6tM6
B4KJzh8egXZnz1x3bfQ+qYlaliDnMXz6Jc3Fw8u6YVyLUrhmr4UArIiQBgox8f+I
MvhWwhEsPMQQ5wtpF0INWdD2gkNch5Bo8/YHK/dHxeAKNXd1zGokGUloBhj8Z6lP
2aSXHqgLkyAZge5zay5sX/NadCpIPIauA8v7q3tDQpO6rcs5qumJzXDN2KQHOIsy
LKQKaRqsx5ERV5xzzQ5DTeQeinHrfsL4dBTZojpzmlH64CsqUf1XO0NsQ4vxsI4r
bDnvLmi+o5erzBB9EEhEfetngYc3Q5F/1880ncYZUzEMLojCmH4nf5ZCPyorf51K
tynvw9l1hzVVd/avr1Ntj+681/nMdf1smDMx9ZJU/BfK8owbLYWK95eYjMIaVvYk
NpnzU56e7gh2PXyBn17M1vN0AThlLJSu3QMaKo9QQOwAtmrxsYs/47X2BPcynfA5
9iS+L3P6t9LYfwfHe36kXV4mlUoEM04xYA/NbFWGgBLSI0CQ7on+c+MLDbCYJ3rv
xEQkLzzJwCEzpSrpQdo/GIDXTLVfajZm0ZjGb3yUOFNOma7mQNuiVvGN0F7oTanA
1ykIumpaQ8DMEquOdpZS5IsGykwzkjMgaAH/8NAWENWXH//Z2Pmuo6g27GP44urn
/NauHWj5O+qPNbaxm8Xya6BrAbo7AIFGKqO4f87faeQm9lA6ONgsc3gssahXZ5hz
DP1+Pxn6g3MHNO4jWBH2bWZreOr4a4Mp89phBQhbnOcpolZSNBRb3s+VQjUej3yM
qmZpUU4hE5CeFX5EkncImS6nq9a6BciyU0OFDd+ptGYGiEpWDAjjqC0YAstVChwX
itJwr7Lxg+Ego03ukYgxYRvnYNRRGWCHE7ZozY6QIkZFBuL0vRm/kAyTGZJs+6L7
xY5A4AvKDMttzHRAhIHjwMaW/q8PyKVfEwg4QIcsiH+VArroxRcoPyGUkpPALrRq
kdGmNFy2PwPFCFUmX6xja6gQBwLzAYghqiNCgMfrf0CUyR9Fz5iVcNmLHqGiKSXb
PjBSuQZeXAL1uwA/FbKCuxc21axf3+MRdN2qOzLz0Y9kNPh8X0YbXvg9dY/iXgxN
h200pbZsaa85AORnnG2jjIrepilP0o8HQUBi/Dl4KhZU9l3Djflpm9Rhr11uab7G
Lt8v2SHQJPHWCaybIvW2LoPVow67i+bHXuhDhVgObFQ/N+6WdNzQO3FXgnXpbuz5
WigasbwPDhGY1mj+TSp8QyB+uexewSWkBOqZuQPJaSXwC9+1IOfeytwDAV0ttL97
1M2F9Srfngm7f0Rt3whuRmg9oZmi+LDxdwuopDrqUor007zdZ2zgR7FwpffaXtuR
xPwHQ/53/ztFOYT8O8k6x0q2mhG7cB62eIh+G598P4rWI2UAwgagmysyHdG9unel
3hhogau7wdV2cHkJerozygynzJa5zUeWI99lwBwvDar6fRYl186CRJFh7VZFWeDq
s5e7Jn4IvM2vIbMvop6sRzW8plI6EGPFFsIDz2+5o8Rz2AgLmHyxIqgj+RhG2dbE
+efpNJ1HmBLHySwvFoz80NB4cLiaZfsOVm/SGsBsVVBEg05FxP0ZDeTrMsgOHQvK
lqnyEDoA17JeOS35QYlcsAitrqcYahaY6wCf+ig0JhLvWLYdys3WCd0VnVwH8HIN
nVw9HuzNp4P834ZX4olonmefN/GlJTqnSlK2LRvcoWTwSEBgjPOjeyy0iuxJOWJD
9tmKNJ9IwF/4jX+UOGPRYJf6dXC2dv/9L+esMgZb8wJUydZq0yShaCCBESfk5pPA
zmE7wXkt6Nmb5yqLpylS9NFTYAVEz03K/zOHYwKwc9Fdak7WSL1Zejldcmyl+Myj
9NHMC+XmbDA/CSnzGzGMLbBd57mpOU7xUs+/aNgpDfMo1tbWx9VPjsViwfiUWlRI
F8pJ0GplmuEB7urtJ5zm3cGEVDY7gsLHJWWaVZOV7l6Y4K+I/3ZPq9HLqZrm2AZn
HEdZ6H2MCt7nbyyaKLJX0rIaRu7qaT6m2kNjcZYsKB63HdE351hGq4wH9W1f3vk2
UAF0uxqg+EDbKxParG1vm18Bzvmsp4Vg4mrCbuRAEKGtjgaB8+ECzSCR9ma6EwBv
En9gnCK71QdyXHsM9N6wokkdxOrE/0sklsXiIQ0NPvqhXuNSUQuR1nN+XzZG7QW8
6uT41cfPpgTki9kyAi+yDYEUUdf4HLwjtJfZGWi2FowU4r4OpxEQOSo8rexLJEP0
Q7Ody37VdkyTyYEf9SHv72I252jQ0FT7fxh9BlcNCAJyEhUjp6PpoP5+nHzqeoEI
iNzCx9RbgEy4SE3rUjqgkNVVLLWsrf9yjKB5LJ+2Rgsin3MdpJniL8fDCfwia+wD
F/XXt3V8N1+GoiFRqjO/Y0AnjKFlgEJsrGMpZ1ZB81nlDmRkujBWHmDqNclVQ3XT
fPhxmG4bdZLk5QjmjkySPEaR46K/tK3xdOnFhvyAGveeSOAr5JrqN7878BuXwgGf
B+zJlF7sLjFH9CuIBhHTyydEQJKxhDIYvyuoROfatW3Bb6orX+h597MlQBMPiIhq
AcVrwAsoaqASFA8RU6vJ5At629W3B1xcTMMbVCS46MHkdYPrsGHWXSK8z8tFBHoW
spEdDMixLmHj4XjJ2AfUOO+R0zG1EWZcwj2pm9OSgtXiLk8YffBN0zQqLey8r1V4
DkxSvFMNmTTYHBD35zmsW4RzLVed7Oc4WirIvwpcUY5NaB5p8t8Ej/0SYlabc4OL
rt62h/jjKX/t1SyzeYFX7cdjhyXDsjwa9C0yv1gVdgKX6psj42RSP8VQP6NSNm8W
rYfrOsIzcmZzTx3SWOmYjQduBovSwih+OZDBDzxSZjStzoKan98xKUovcFVTbR//
PKOviby8pSu2lI7l7eErRahRdNwsbqvNRxCtYcn/Y0ZV5DIGDL4Q0nB2qq1Uia70
fH4Pdksxn16CQrvRDKuPx2ZxTm0no2kpGLuUHCtmO2dWXo9Rmvi/F6JfbeNnYEWo
sEG0FSocvu6cnYVyp8YIvWQs6d05KZG9OlY781yjsgzr94t9locHdmonFXhu7sg9
JvZXqOwWAgtxWDobuuJPExvZm8/3k0YNaxxRKgWRviPlWZwLyxWdBwJdv2p416v4
p4gSX+tJj/nUDejncF8TFudHXvvp202Pw3pK7bC2kQ34gDH6CM+OgsuIRoLGfcZe
9EugLza1Qj6QPfUkUDcfSGgcwfBNGn9vI5aRSz88JuRgB2oBqZl4j2h4eejc4P5G
2Gle/1DZ/NDkO7X2eTFsxVHVevLQMw5lEu4p1I+fEL7//grFSIYfTU6hipO0WSV8
5Hacyy1OAmjgZ5DxKX+f3QbtAlhnZtr1/WzRFuS1Hqxbkc1QYnunXtEvCCBYT+u/
WMJhsbc5Cn7pxfQBfdm5PyE+XA8AZoC9akP873hZjWIQUh7AHn2rAy4LnADqbp68
XGlwtEvwnaqcZDAn+EPuK5S5GZxV5Y6FH5ExRB5Qqvlzyl/N7okgpwWz2joUtREk
dAfY7BDthU5t8dbJX1DoUkqeA6rcielBfDp4XtfyG4KAnbTUOQdU+kbmOdVI+0v5
9CzYa/J9yrSGVvvcfxGmhP53pyYGi45ENnLZFMro/2xOrHSKswXxwfGYt4d5QkbX
ZJYINzrHR1qsX0A+Uw0e+zDg9ySL6JO+G/MlyXos2mVqWBevwA63rhfsmkBQB2qX
2Vd8w98VUD+9iSGkyfV3HU9MAFOC7QmtMvzJ5k7r5+Pk/uHx+DMfCmvuBh1phsmG
1jrB0GBmhNBaiRJsN82rXzacrYizKjYspdZRAOPpXBMhjAlBjMF7vxi2N1Nc25YJ
O1M2NKl8ci+C0jO/FxfVxHYX5cnFHAfmUqPrpEmXAGvKgXOrbLnerB75LgxwnC5V
5iUeQpSkfGGPSVD3qH1P/opo0EM4Dx1vx+e2GF2S15tBqKlsFNNUuIgeG5T/eNip
PQBVMv0US2baf7AmdqxY8KaZ8uZXp/e2aly3uNEeBqTjF8om/n+VgpmOfJFhjoww
/JiE3z/NMoYVrvRe6KwBPhSWvoqkOioLSElqlCWRUZX+jyks4nENjYrIUSYPtupl
EGF29Rbp6rqfsdiFRv+cxP55SLij5qpgm3GpBKy48PYF9768WVZLfNoynnBckcPn
hW+4ajsOl+ylnr9YBJ62FLV8O0HbR/cCqmvFo52fqXRh1TQSKzKR4xObZL2byQkd
xAmwwG68u4ooLrWwKmbXHh6DN5WpLY/3+q4iC+YAEM2fe6IMsnVB1IotoXS3nZqd
7VBShPT+Wflu89nSFr8rDAj3mouCH+BGgZTBedg0YAaQaIpaZklKFkp/EyTKvzN/
e7dNW/ZN4jAw3lRbmy9zGIMUDix1siKytTMWfrF/lBxEsa3v60cw7f3bsueeL8su
8wblfy8TOwYFZT3SKFG8jCn4rMJLK+FoD73IFJR+fpJ21ZM1Gm+WhRDATBzB1wzF
F63lvpAwheAx19gSF2IYu7G5XLrRQmdoOBNX+Q0x3IlbnQr0YtEriozio6UE2Sbt
hKvGcBdATDoTxhP+i1mtQ3W+vN8aFQNffI8R141jEpfhPGrxx0tKOZT6k1D0s/yj
fn3prDF8m4YXcqLyDnLHbo+To0UggrQE1lRtz1iKe/Ac+YvY3Un17Vl89odGPU3F
qsVUkiBXWYalQDoXGyJxz12zq1gxvF/HzCoxlUkxxAQrl5sEsj0d/gKhpbGM9Kg0
byL6U1EKKZpBElgxPDwtraMv9pQSv85zkQLNdWaxwDm4KH6poVXu4Mzv0LJgc2kT
/YC+YIS++/YPQqwD1lhXrM3xMfweYjycm84n8JzYQqUGX5/2pGYSmPJUIhTWXl/L
EaA6PUSS2C0uA1FeoYTbMwf2w2BPiQijI5EpsXbZNR4oo1jVruTVI3oMDGvyEChU
e0/9P2UU3imyFnDcHh01NJOI9DnWt6vhWFbvujUXOkFs67yLAp2uxJX/BzOvl60y
hvcW/OM3hf/hwOAWA7IsG3ZTsR58+IzuIMW5+1/kijb/+Pxptc7wTepk+r+kzINE
Z9pGlTOnOD9VlA3myzOfaNfK6O4B/gAYBQam4Q9Q8BbO8kvVc8MqKNxXtoLmeKtB
28cpay0m2Y002qfhX5pg0j5gJoF6skkBYVHw5gx1GfMUZnrdCuVeU9okKP+uQdb5
P0XC4B5ohme7uMrB8Y6/xtDlb/eyhNmThAGPldtdVJOLxvYpipdIn/d+h+YBle/m
oWfaVXNpczgKCuzG2kjatjIo9yD2k4Ja5H/egI4eU/6fCpH4OR174s4AhDR2CWxU
86JFyjmrBV18ROebQ1ETQEDs+ya9Skp7HfFONlfLXZ8a7wuFflM+iUk/0jNbjASf
/cy1iMGvs74f0Mo0b5sxMaoYDQ35wrSIP+grbd26IpzP5iw3pSgXHS/JaJmZrCnt
tJhthECuVppu7DnuoQMMm1lUWIPsqf373JyhbmnMmM7vzzIoAVxwraXn2xCx3TFt
8Wi0tePZzWiMAAJGL5GMe/5REdfNNF1JG+2pGd6DPrjaKyFp38HKMRbmWp7tjzMG
3YIdUoupzXaM5JRM/exlx/SSeUjfyuj5VckjiiJJ89J2WQfrbS2PyQyvyw9etiCy
fE9ZbTnnktWlnHILdEkiKOvxta1JolfBflCIjef34h07IdXnQRgOFhKPckISIRZc
g/CbWDugF+KL+YgUrfcosXNgWuQKYekwctNCn64TEzSw7h4eui7j6Le8aAM/8w76
4oSwYN1AlbLsUt3pA7eyNRaQxN4MQKjkdkzTSz9qH8gb38cAK5RKqif1KDuV1KO4
W9zIsyaqKW+3jMwd25zQXhQa+Eahzb06GhCNK5pNiVt7yIKi0OBFoOzRP0J5np3h
ju6Z61nlMZmoxywx6WMAqwvyDC4w3fZuQ7f3mCVRqw9pYSvcBSUXrdI5OnUevge3
q3semPW5zqK2Il8fzI8ua20y4/TJWGCHJhho6PDnFOP/XGAn4aO8c9hNscnTDnSP
Qo/maslzpclfqarB+HlGwV9/DKE5doEJewMn2BHGT9Fj82+rbPBUH/h1fRA+sUZa
5mkDhPzqrsQVhfKnUWNRATH8dfWe6JXV2MoadfecK2EiMDuRfgsPgipoTM/GZ0lD
2RQWr9/Z9Ex8uLjVPkZnQB92dN3kYfJEkFA2pfOCRAV8hP0K1vJV3o+6vB10c/Mj
x3pe4P4zC/BWOoF7w+xtEfzzUyNCYY2CX5XpTiRj6FgdLLnNVX3wIaGhSN5AXNZ5
PELGvugXN9H3qa/NWkDfYxKIgMcR08Ss0q7OhuP1XbExfiWLSSlzXBJIJul3vW2e
O1d0Jx3drjNts8s858INguI9JxoT9kpH63FJ5W+AOT+NyOWgbiBHKHmlfWeHLvzI
r8bN3oxKO90V8WAEE9ExhsFjS7XVGPbDSfo4pTlfKwxVikjxfX1maP8vrNUH7aFj
3msp6AqqT6NOdWdUEjGD5o9wGJfjiyH+msgYtHzLWIydC6XRC732ll64ggZhUQFX
O/Bxig+fpwBiM4k472iA83cuzYvvhym3WSGCeurRkvjiyD90nEVDyCOTN9SW1nai
bN+bzqNhRV2iAsF8bt2/RrzH/v7ZG+3US9SWnJDEkqHggaFBJrX6V6NjVjBdEW5t
uELG2iYN6O/LTe42c7nFS3fmIyNKpVUggEgy6Q5lluymjy6MxRR6LQ7h+oTn11kv
47om7gl9k55Z1rCS6sKghqAA71D0JHXQWak62AfB2y8h2KL6qFErHWrB0yUVzJ2n
0hV8AMLjWdP4gg2S/1VNfQ7FZNmCvkyIJOW02WlrQrQaQiC/As/wmV7kvnwtd97o
dUw0hST47EI1bt9zHzfTEhM/dcxWDk9b0EHQTOa/p4vumRn/Cl9NVaSnFteZNINF
BnZnUyvbsHfo+ixhPAVab4arD2YDuXa8+waB2GEjhaSc248bLcoOjf6TIEgb3MgH
Lf2Mpl0+mlUGlNYwAUvUOdSbIHQh+JmK3NKY+l916/KBu9QSecqiuDdE0sv2vHNA
rABFKsRZ1+49gE8b6al6m0+M65+cAzt7iIuwI1s+InIovJyTN9GnMhLVxRmLsiAI
VmLGow61Zphmu7JzHobwCrCKLQlmaHrkbFhmR1PImfUfiZdUrRzgL3h828XkQDfh
QB3GGvhkmL+Xr8GrXDm0PMFwqNQ3LxgQKRb0zbqD1IR6xglV9HOzaBWmaPXlmRq/
GDwswLSoz0MgdHUcti2KZjZbVN7ZZQyT5mKQKY34gqOjBBNIG5rI/QixO2O7Z/+I
L4X08c2PH6vqaJQey/YkaNRLtR9iyCObX81DmstTXjfjR5ihRbfN83Zho0Sr/X65
XF7qlAiLUuibuhu/kBoAkZnBKp9VVRcPiTKo1qq2u1UC3A50HgcGy4EemDO8vljp
92h/duBHsge1eIIamRBAFVlQ93yKdWE42bHamCKJuTcyTn2576lJXPDg5zxjU/aF
BU2FX+xJD/znYqgpouU7/mkfQ4+qPtX4PZhS9dE4dddaa9BQcUYjIOlZ1noIuaFV
7HSIUevjgdNhSJnZRjXL0D7vGp8e/dWimyjvDoh/rc+NxrrdKoqzv9GLsxGTzpUy
PK9+u5OdQ/vCRmuLrRLUBhW9FXjCnpodB1cyg4pLJgyn7VdA7rkaD5f141GBCuDk
iWdytQypQWFxu0QzS8UW+x1X9n4WMX2jjAGw9ls36d8zlkN1iubDP0DiKDniLP3w
d/wzuXnyy9B6LvpSFnT084RhN9+mP++7mPDkfP3k6V4DvG1UFmTrrR9q6npgRcZT
LjsmG7Pe4gyVMzo096FrJfrF8D4Ni75LAa358c+XC/0pf/cKyEJ1cS1+keK2Bu8g
aTWtRtuG1HYazItABcdkERbhgvwOLKgl4iro/ehLIzGnAS10DOdJeYcXxo86ZDe1
aDBLqKbIH0o9mfGYT4uwXwYsVZVok+N/YZrV5bJQbUsJz2nkBT/CGDOrllP2WSmG
Q0LxqvGLQeTUN4B0VzZG0hjr9EdCXkWuFOmaCZugnfhUiEmflhqkaycqMQoYTVB+
qrWW4YP8Y3sYNgnfueBYlVmKWncXIG+6ExGf1P5ruIoJBs4aNOlk5OW5zTfFK2Ub
3XsL/ddrghv0jJti+mW530qorRDMijIRsCB9v6M5+OqZn0Y1dCcDcOMOC37ule2Q
mfGNYkhgmeSh5CWdN+y+q0tIxbV/3Z1oet+tiprECrkrFgm555aUCq0xgtNujtRe
aNfeNdRUR9I38XQlWsEL2KiYMQ39L2gA8hfWiSVPqGqCO96yWiQQUqKh1jdE8pR7
IINMr7AN1y7agpLsbbNbZdgWAF3ogzSk5JcKCVBIOJfgOhdrIDsg6iyWlSu9X4tK
TUOnsab+23Uo18a8XY6krW18T/gqGuH5DZZyRKtWhhLpASPjbwd0+0HnQbOPXuQ7
c+vlpOa14SLPL8Vn9dqb99EeYqEzqz7TyvvoQ9l3i5YVk7g/QNVjueYD2JKNt6+F
fvIUUp59T+jN5pb6zpQPaEXb8PT/zXzQuSka7/xXSxG6x22VIe2k2bn3z6Kze9k0
CJfIvo79TL250gfHWr7zU7lIduAzn7UG3bxZdqRnBtVezErw1odtXoq1I8ZDVb/a
zoV9pRQLvPWUbhMdVypqVhXJYBLhZ7AkLfzqsRzA5jj8Zcws78ZuLHeXpO1y5mhX
k8Ek7xEgz9EC3nhwRDq2af/4q3/1Xxoy1l98Ud7d2wMXv11CwDbpVCnUAnAdA30/
284WCMCFWIgUF4G3RxuVxXyV6WxWyOg0EU/6YR4sCyibEnXRMeFNGlZpERLoXLaA
EBvRpRF/Ohu8FumLF+I13u3QnXGrNtR04J57qnKnxh/hpE/4BiVDTpMCRiEhELqU
tJVAfAEEntMh7I1RoYauzZGm9NpyhoEvGh3MIX1wMZ7Q0knJRcV3vl38QHXn6pGC
GahyS+6R4s3JTUIqToLAnmutwSXhBfeJfFeBSW8ceSeWDMtskn/T+aFU+nZFnuoa
53B2HlJ0JwL15s0Plg4lFd8oYcSoc1+8ofLSHbpw8KhyjbjHQUNm/HAHfCm1c/Fe
mmFWFDe/Mx4orZwbwMdbiFxwoUxi+9+k6Wm6YO8iaQ8I5qtJKCqLmL6AccPVI1WC
bBnVKtLHI4MlCk4G5nPVA6Ga2348LvQ5hOcWxw3OHLaGaqlQy5Wxl6O3gKyS6EE3
O2F93/bGZVouQ/1DFJ55o3GLyG/TQ5BhMWd+zszmmEvQqeFAUDDZn3faHimyexaW
tC9WYQSyukdOcLZ+s/gHGO9PRvN/30NKelECJXjlYEGMTL8CHlBLr7VJG0/OqZAm
s0W8MbKdJOwOkeZ5fDbsxvUHunDfxGXWVgRQGOEtBXxoUC0m/mYfDH+CxiwWyKvl
Ia5O2I6XfomU+7BCM2DdYCtLC8rERiH+qlf2vkby+n5z0XduRIHAm45j+rWcZ7NI
SJq+B2clJsEHdLi2vMWvOfPBFQ3BGAxdn5Lk8aDJOlb6YTLJANhE2CKnPgnPQo9P
Cclfqoqepir3HgI1HyrRbaeNNC/J3E+MKTXQ8xREt9no5zyNGVwZtOeBtQxC9xDB
Y8QDzjdIz4JfBcExDZagab+9GfaxkNpN2Z8BgB8xz00XNf0SIDYTDjw/QwBqTozn
rHcmvbTS8X/ikEdVMNQKtOHEeZotHKYhaDD49Cn6/hIlwJV+WsMm3nmYUjZxPHdb
iqqOWOJDxvyBTMdgJOVgJS4TrPN/eaUtvhseliaMgNjbTpynvmJPSIzoPD2hrB5I
FqV77b0nJqz4Z3vWF/QSzds9qmcBkEJbhcRH6+vntryBYfw4odX/3vHeT7lxgv9e
uRLUyO6PAMFsrtb2MWfscF3w6hfpaOmWzPSXZUkcln6yZ/6hEL8/soTmKIPuxTP6
F3rnW+HQ/c0DctSQnWyk4xMVmIBioXuNdHe54txZ1HrmU8inJfpbDL+JIqzmkSsG
UBaLBiBFr/u7P1xA/rfgKB+4JodyWcmZ9+K9hVBOOSDW3revFNebsECzJ0hRdMQ6
UBFlFB8LjjMSZsDftis/bMpqTWnTOjpCralJA0jP2awkofK6pRfR1PgQTpe5sRyN
AT9AGDvE9oO8gvKk1IKcVOUGBFKSf5PiNuxjglMcFKE6wZXsPLtapDteOsLTwiHx
q5uLlWWutdte4CuLCJgkNzO7xgnW0tGPBGN5w2dB8RgVYNtz5c7AamQETunjWRgN
qaWAdmHFhet7/UoU9pkXqAAJEOriY7i7X0r2gAg6fVnwvNLA40djtf98Rcj3rZlw
Ks75xBrAggoZZkaYSmRPNMYSQciWmtJ10pqjtGKuFlTnZ/L0LqV5yhUKozL8B5VZ
Zh9GyiU6sqj68uiiWnT8rfVrLoxShq4aVNN/NpOYB88D082Rb4jW+/Q1HsGqzkn/
B6Dp0Sg56PXFV5FRB1X4wsfg+5xU+kf2hjVra5RijsCwcK1N7+IL5VESsoqdUjdk
y4kMAn9nq6obMF2811KW2RPyeKwU59Miks45GKhrdq0We6XXMfsJNcHoD4PnRWhi
4LLeuxxxsArl6gLUk2YoNxH4LSBhXZ9O/13i7iiS7qeV5V60u0zZZGHBUIICPYVF
h0HAR/Ko0pYb/cS5FwzlHNTR3pC1OGZ9D1e+h9iVAhW2k8sIjXJDy1THX4x4cMhH
bXb2wTIKjqVNC4QWr5PJDf8K6aAAOpjpnVWIytyN3NCEafjhuOyXMi9c7cXIzWW+
knGwq7yUFwbE14dUR6W7Vt+5oOz1SzrJmCiUCwJAwpc+iAfX3HFNqE/BNB2Hv9Cc
0fImT5Em45Rk5nyNx2yUQpti7uW5TFGuUrkr60UGfkZBR9jMTAhYSiYCJSUhBpfj
OdPLb3oJ6JHBaKKA5cNk9Dx3FJMkMG6RuVTeESI2iUYlh6WT/GQw0HkfpoggaoOm
gq4A8VOlkA++1/8exGqpD/T7VCOhnhRLZISnjYLMkRJo3D2tyh7PB/9P1aUtm8+V
/HmzYsknUqokcHTXAK5syYCVs+mUgu67kEvkt82tsdBDgEOEJ/Rlkt3AKpnNCGEi
mvpDK8730N6MY3JXG2yKRkomtC5cCRaAOZ1bn44/rqCzipS7fDIaGrEMCqlC4ULa
SX++VavSfeiZLpDbkg8F2wM5BHtAeoMPceHn1nTuxZhp4f8LVkXFgfO7xmY7LhfA
9eg/hpK5g2jW9nwclQfGVFVgCqVDqOSlr//3sw0+Riz5em747mdHXY6dgXgHb8Kr
KpQrA3GoEVphwEEQiY45wOoiBo2GBPWCwckoN0BPmhsr/zqRUiqZsbPNP+a095gk
Qbx7mvuR2XatLdQ5NRezv9X/OpH1lmctjx/3Kv3tWctftUtJUUiIL9LrbOpJJfWa
swN7GGH7xdK5VqHPWBY7G2Q2d/EPnk9OZPF796/6bsihZ0vqvILVOGxbAUD/Uy0s
RYASb3syyaWY/6TKyzc7cp9/sPQ5SHzsz3ao0C0ZjuXvPqOiGfrzyYp6e/+esMd9
TdwEB8XIy/AolpIR0o39JjCTJHMpnPtyo9/t2xQ/IeNJhieQCUKOuem7Xgq9CyBq
dQBTugY2dIX49oIvomCIsas0LaGP91O3Cvq0pZyFIQdFDadi/XtwRUjUHTwuCxwO
1750UqYbB0TONgCxim7ZgwMOahI4fMxJ2l7h5WuLb08ZnGuCCbW9GMnxZVspjnaZ
wX6OliW/z1LUoArAPoA8cNDb0BABBYKNwQ/y+dsCVntmN/53BAN/d62b/b39ELQb
88Mo6+UNXxecoDw6lb6bPiPDwrIKY4k1Wujn6cockU5YlaEheDXMrGCwivzhiOHf
4QVATk0P7/hWHkYfF5A0J2KJsSxMWXalI2TisKzjcRrOwQRyMnNfSFH7rrfeqkmV
9YAgSI5ylQ5TlN5NbnD3YrA5xE7ONhEYoo8hog9QzBoTBkJ4fICCdsCJ4RXB3LTY
WPaMqJ/d2LxY6r6RUC3iga+64WX5dhKoPcmNhz6BuyP91YbwdvcfefipVfoQpyLc
57ZEBYtod1uSG8vOL+HoAJiBp4VZ10xKL4JcgCKKRfl5mbat9J64le09TQYAN1mq
M0UhRHLnI73eNaaXDlpOxJsGxXyVxOnOnYjTDJ6sVTajPsR95OY2RZ0JKUsk+4PV
1pGFqgMHLPtplUNKL+JUuYCrYAb5E187I5kGLBlOdqyBXuTDHxNrRiHmF/7BxLfr
YYSRjsmuWDgiJooo4aukOZAFBg36yviZWCHBYhYWeCJsDXQ7NPUwdPlJ4uL6MXo+
3cMbjgc6tVfS7PXbzj3QW4SqNUPnNGOKBGex+Wdl9hsModJtXfLKOZYVJtOPVjfm
9PDVAcMC3/JbZwDEbRKxIkIdMlqwrVno26wVK8sA/+buEJdLzIB9GbmgX9VNIsUL
bo9NA0AXgnlbXlfGjqoQiKxItL9jv+zREyKWXRcjcwi9a2isIUOuH3Apl2ytrqGw
WanTP5YdKbRmUNzntEKbT74mi+YcxBkW3HBEeE6W0OTmzOzPOIxl10jx/csXT5O7
oHfxAbP+8TwO1uyNxZC7gcK8spl+l3+zbvy5lUhixiFOGkmfyjLBj2QBwkHD26dU
ze7CJayAv1oQfz9PZLUAihu9OUxvVfCGr3RLm/54LG3aQMFOI87MD9Qwrp5xnFvN
PZVXcxzEsVsXQ5fwaYBzCoOS54iQO5iy4LexO1ZS/A0pXyHEJXPryxqBwAv+Vd9N
Js89v2xfxO/+Xna+foe8I0nkhZDFDVJWpU7HFLNTLqWpAsNQbqiU5gKxLiASRliA
Ajfxox+KLeq4Dh/9SjixsyNbv/hLwg3n7RhD+fIfZFSVbniMrEkze/7lbFhDz3Vq
iczIh8emIfbmsEw9C6no5wCThyKIBWU9H6/A29SxLhjftb6ocTcIFyyxa0ABg2jW
R7K7E1nurILqLBSqVasJ8WFANT5HHSuMRqDYHBSHehxY/P10irXU47h57VZ33t/o
ZuUfm0PLOJ6DuYhD4kGWq86KP9JPU9qAM4i0/9LobVZYs2/UvLwknWNSFuqYH91l
RIxKBMJyHxKHJ6kkvFYK0QiAoOV6yoQvrGOkiS2Fec3vo/iSnCvefDM31gZ7Lfey
HH7WXS2mtMLKU7Qtbr2biaL7DDQQuk6V+DD2zv9KhnfPgFFA/zghoqyezPynuM6C
dh+F74AZxR292oiWAYzXaIQZwgUZ+WSSwBMQv8V9gWFzlYquXOGcoDFCewz1PRKe
55/wwdn61i74IxbYEzweReM73qqgjUVn2+QuyFmOccdi34Qq87dLE92CZfvua3aY
6qmgJ+zdilMAROehyuAAA14BXhJ7m0hDa6t/F1QwriOZ7zYaA9/M2SIy6Zc9Hqmj
876JDsuDRvGwzy8npnWenoOKt87zr0zyAZok5qZVZ1qNH9SVGNR+Gfa+VbdB3rR9
DhdEA99m5NLHDSZzqJCR8jd4PKV0LyJic98xHs9/ZyquZGJBn5C0/pLoOaQXGOsg
jNXYfhWFECXBy9SHXrK30AGDaiP+TOJr/8TFCm4azKqw+Bttc9siBIZDwL4me7xz
eG876+P+ZqHWiOOd9SgoozylFdjzQqNa8EfJys6SYO9fY1xcKmkY+PFgMdHaKxMU
TMVyzoVc+WRlT9FTK2Wx561xmd8Pvhci4ZclWehILXxDBPDU26pNG14dRehLRs4m
B+5YogqvgmeRab/xMjIj/QOlJp5FuDSKojrxI5FCsa3rS/G4Qw7vUMRyh1XDXSe8
fiObVPeuMItd5JssJBQiGWvcp98shFG8SQWIhqf66bcaB4OwMdVxLasmOvBE7Igo
Titwgs78gsw1UdrcKjX67+kDuh3DZ6XASwUUfRE+RBZs9Y5LG5U3oV/eBgeX5Cib
h93dMCQWJ/ycJP5c6Xt/SVGP9lP94Il2oQUPKDVo9NM8JOHkPsV9xYbANHel+CRv
vSVgDEIOJR86g6u8eyowNlI4hpEGuSdd5BsX6/siak3KsK+7ypROJqIlLTLO0Avn
86mPRqF3is+3nVNZA9xRCzocdwjAvkoBtlTjQ9AVpvNHWIddVIOQPM4+cjjNziFM
aLkjiagtjy9wRN6DLbVYmGMlnyj+9Xes7pewvCSRm8xOtVXeR1s09W9LBgUmliKg
3sBABjglplsLB+ls7b8H6dbnR0z55a22hVnFQyp+dqPfEBLVrKukhFYo8LYoAfds
o2ENfwjC6ofhW9FxpPT1q1EEhsHkpML94rtZR4n2euaankxhn5yEf/lcwOUVzjP4
HmNLQhF2SAY3PKfSPT7j48tGmraxzXHWyqGsmpvzf3kP1JSkG+6XpFTcW22r8WoJ
e8UY5KehA64PseiKPl6s+V0QcoZ+UW8mNQh3yCJFXN+A/rpRM/5omEUkAH0mTATY
yheOXvJGu7n6HrhGbGYG60QrV8iHBMdLnntZgNxWXBf2v2zC2AK4ArnyhsCT1+eV
7e55QZHrVAp+Rc3ozR0c4Y/fhDYrBi5GGHo/tGNE2fKhNdCHxmMDnyvXDde3pKGI
U6pnj4mE/KfaP9D2wjgmx9MIxnDyKUfmMPEJwDpqBZgKFPXmu9xX1zppvvjwJ6Dh
GwTZ3ve1Vzlq0sojsgN/VoeIMjOKcEjlKokxjoh0UfstAGyOLohYp5s0lLhuz5Vm
APW+vt90JYxnxIEC0J0NkG526hu1UVz0M5OZbZWnzSLSr8I3zlZOlHRvpu1Q4OWF
IXqXitxUOt5uZx3E+k0Uq3DfGaqvtNUDNoVm7QJJoe9J+HSj+jDrGnJVBM+hDjLb
DHavWbhAhYY4meHhNF2qFKtPYaJKTvm2bUjFUQ7/qfG/jzJ74MWVJ1Z5ySvvgzIB
0qSc5UsbsxTfO5T0i4BpFJkMR+ToshXrFa9MPfhwRsJKtImt7RLQ6HGpia4oEExa
++PzvkGPdrBbm287wThEYGhUHu7vF0OFhlS76lrfT6LF2zawZa0PeTRMb++b1WUX
USiHIHwX35Fjgpru6semIxGMYW/1KfhGZv5AO24GEhlZvEg5VeQ1+XmE6hvXr3s2
mca6Xl+ZROUnpKwjbdwZvg/NfxQ+WMfIRR2f1fZQGtoZKFtXiBf1cUJaMM/6gVsG
vmjY1x+ZDGt5CcRS69yxy99O0aVQS2LHP4sva68YcB8PSyI3qds1DQYFl5ZBHNzj
vUt32XKFoyij6ThVsYQOZU/AhIGnKrx1T7VYuePJwAoQCV3P6hhZ8f1y3GxJEeDy
LX+Fp2CC4U+rCPO5IjKnqrWraZ0g93IHrZg6AV0xU2apYpoIuXl5yCARYhw3IxLq
L8fJE871kxsZiZZF46gtrGcM/QG15ptVzvC2957rXxr4VllkuND43K4bpQUE8p3E
pwHm8TvT+5SILsfc94aNVqfyYX7iRVpoZBzfNOvaXTU/bgXmEqSOicPCHQgRIbnp
0WK2QlLKA+dGaMdcH9qzYLwbjjZZGFZlFFB5Er8T4380UF8GxOwMYzLgZN+Yownx
B7JsaVOK3XDTRRqSriTIU0+kjbXe1M89JrIbfjyQzWkGu7tE0yoW450Az/z9EGfh
i6h+cTVivdiY3diuyznt1BVHbu5XZugrOn9ED/wTow5sLoX0jB+j+aucu9DHTF+9
QClCemTbaGGfWiBGT/sPoAfjc+50S8eUdS5xDi5uWC+N5sZOns2bCe89tLTOqNP/
YDuhYGETS2A9PCbunVN395+8Bbki0eJicSDtLQvyh2HNEiBQBWrrgPledWn8iIvf
hEENgkvTcwPTvH/v10KuQ/EdVQCKVkLQGg3izLvBLf6JqCS/yKjictpdurNXIftC
X7XZ9rFRhafL2ZQuoYqKUv76MpNZKhKoImR8I9quivHiF6KXZgms1m6T/GrbKLgY
Ei/FHpcJj50L7u+pb0ceKJcuLMo7XFu2mAuxd9Qkm3jskpvT1Z6P+d1QrjC9ec5w
QSWywVoKOcKlYoB7eBkOQCTr16D6bXNyZ3DhxOQx74cAmFwMx3QZPhWTWa1BYuQP
S7ymyRMJvztNMa6m9uQY+LmjEEA0W8it27fsZTJWSg1fiXKkF3Rp/ybaUqNALxU6
cYGJDDh3HSEv1yWN+3HC/Xi03gvKYf9aQPUhxOi4I5cRaJVLATXIFDXcvuQ9/xDE
g4EkEBWQ9SI2LNMc9Bmgs35VIEkzcrPtdaWDf9DydYxCxZz1f+L7LEwfqQSwJsV4
5iBaYjbBubuL6japk4qf2y8z7H1Jg5K4VWuTsT/eHR8vKfrw9OR3LQk1rL84O3f7
FfVnXISwgbZ0gaizd64XblzMCC86OYkenmzsonAUdf7J/XFkPWAYsaIZQR3ktsd8
dtomw4jFufiwbbzARbLUhP22JuVjb6HV+EuqAlGdWxLqri7jpVm35x2Tv5nE+utJ
hduNRI1GAbE5PvfGjj9IcEKqhff5CnCEEtoLVMkFdL/GfdfrKxAlIdYfYBBHrOE9
5kY9oDBjXwyQSnj8ObbBRPzhbLMw1+HeFE4xuTcdqvf3y+wGABYN09T3RONCd6CC
+BKyzGxOqSjyNk04TNr/URIBKCCigdpyr91CWptsmPyuvcQIibWsfaYgpW9oKbqX
jZGnxqBORX6obAuSMiYg5kWsRRlcKqm7E3pMVh9h2j0FDXgrYkZXajrG5a5gC0Y4
8QQfqTHeMCLYmW44rXbDvpgggAx+7rulAKAjqe2ZP/CzYu509xR9r8jTdxOv350Z
Je4tfnykpAoA/La4S+lM8IfvIfLr3QxnB7euFjjcoRCaoxLSCGv89tXr5PC6qp98
aeMdlz8teJDFigec6vxmbI/vRRRBt2LXOmJGYxwNRcVQLYuwr2+0f4hXkOSKdD8W
L4MgwIwDboKDHhx/ktzi1tUZ8fDtunZfh5eCFkBccXfKZVqNiAEAuEb0qiwgpHng
SDIoXfbMfrO0rkD50Epc2rlKbeFDYWh4S1vYQ1ukQCjSL3aJ5a1SHY2t/K4Y8meH
mEMHpKHBX/gREjlAW6bAouA+Tlm/OZbr4X+eHt9FmG4tbPksQVvEVq0KHp1LmQH4
JzDKaTGgOi44czmBeGc5jnTmvRH+eL7yejWG6gBcAuhk00/y0fJFcG0DoMJpZMot
8GKFjyTrmmrlJCYibp7d6g9rvsoyUIgw1oUVAUjH+87EstG1WkDDCpBGWVBP3m80
CNkxW50dy/ecf76pOSwtVUDDOrAMin9Te75uUCkBAbRH4ySUdOyX4UASAA+zTpqo
Pd4DEMffGhh5AOIKLvAzHHKHggLvKQ1ZZWIxukMlMI4Htl1UKEORohv7hN4W+Aii
TcLzIotTD9AnTKU1Eh3ZWvJPS3vxUnoF2oygysyum2sdusvXZVZS/jihBiz7xkGh
5lZvWd1KAopxtjbd2TUVnN8LqWWGk9f6n0zEsuWtBJ4MDEUYer7okMBgkISue7Oy
FbMCOfwAh1ekzWlI9N5l1pGI4G+BXrnboj+vXPyZ803Q/Tqmyirtw7I7pXOMAB+B
v5/WrFpg2zZb5B3boFSOY7KQYwKzB1OgDa1qbTlP+XRh2lh+2wIYqwCP4YqGzG3+
ky0wr0nqhL5x3I54/Zv9y8QxtbG/rE9pKPV0R2qL7njZHwth8mswNp3KZG+5YMBJ
oZifVQhnGeLSHNwN9MFZi1wW/r1BKQ7Yj9ARc6YQOXri32x7i5DbGT25A+vqo95Z
bytMt56/xxajuEJit4JcdS5p3kTavngHr1MjDR0pk5/gXfVpkx+ZEb3W0GDl+8Wh
vfGHPKBdHX4Xl35fRFpWs1W5vXucjPd2o3BLRhRo7FwW1iYQ5YEASvpmzt2G8n1F
c4x61QgeERB5qtbjBAi8qhaKQWNYRHeg8STo8rutQVC7V2oobi53zp71OF1Ag60U
5anGwoGmcLVgtMhZ4dKfdalud1i/NO757lU+cY3yFSA/tv0vLLTzH7ijwYFdYimX
GkqE8yUU/pqF9pnCrHnOIaxvq2HqUMzRTCrVEbDdOwJ1yRIo2Il6Vb6YIF5/mZ3h
v/5Vw7gu8UWAUr67RiehN31dUsRhj31ms/YkyjjMFneb5c8sEpiiX+75hqXLCUww
D9fpIan7rUw6m1kCEZKqb8F8PjAw0It16oGV/o1EMYAxr6mzH9CWJEltA3sDSJcW
0kwXd/WdHoeZwihu/PTGTcU3EDLB/CmdQEIdcnmbw+Il1nwK1i25QmFhJA1ffapa
4FPVTgZCHtKHNuElL/L4OJHmPRieo9LaKOwAurFfMdBZve0INuceY7Qe0YPz2hLU
bu10nGzBTX+3o6b11Y2+I8bkKE990uveVN6hRMk1Xj7NxOOkg1QMHmTnakwDBViy
N8N4CkHCdNuPtSCtg1aIdWzduvoGUaZ4X0WuTu1CEopKXEap39mk5UPXDlTOASLb
LvwAMYio15xGkVPbNmh7prHz+X6iTdwaZr0JXFzuu0ilsGIlRWRZ+nf6Ng3miZWt
rrJRc+Wjq+rT0J4ntqYzMalLyoINYaTRleINl2yL4VEDub2tefv9Fso6h/riV2+l
+HzpGsgYBhrAVoE12o68EckupXYWZj88qD839w3GzpzknOOcmuqrW8eGPryuUuyQ
a+37y8sH565HZkzMxGSOxqlIxYJciGrIm1bmTdoeL/Ewzeb8Fv6PQ/8LVioGTvl+
wSQf3FuGnMQM97wb8RkFCOnR+6X0morpz4A3VCNGWABC3u3kX7QxyrQ631jSepmP
Yu0xIBjh4sU4HctjCo+d1yYeDOz98J5MfOS3p20OGNOherR1yoWn9lPDcpyCL1fF
XzfViZyCC1x0mrdlO2uJQoT7TtXYD5CQh2T5oY+bqAQvLxhjVkANvAbJWPHDmbGF
YQ9xj49qHJXhWcbuiX10YQRleqgi7eXbBl6o7vjZcvpiGp3foEI86CBYQ3B10ehI
1S+oAfo1CF7s05wsTCiFxbYwNNIDuB7gq1ZdLmIngXwubyWINSsSSfexOwQ19xff
/VyDMsmVHTctUK5nRxwF4IYqi+hkXDFKFzVU6dTkRKxzrOE6snf2hKW3EXZ2GT4S
rDWa9YGTkGAKaCHrTfROfucxFr0QIwRpoMRnAtHLmkBWnpi0PqNACiQQ7vC2EwSN
JqKZwMFjr96aqcVMgWb7orbqDQg32BYjJM3TknA6E1y2NDntaHe+AWRBeOippr1W
x7a/qZwtYFEzLLZxepHWql70h40PktSpFfUFr1myM76INFnSXr2xv/QLbrJoiVwI
rXzApJhFjn8iCK+1mNt3HZBDO2nE3JZ6+VAOOhyYvX3aqkFtjd65UgWH0eyDJuOZ
YxFPURPgGFfIXBLCQ8gL5mcNKeT+kEp++v6h9hV5YFBF1EP+W3VdsimamtUpkn/c
APrArNkI1HiKmLotI4CCrcUq6DpA3ScEuNjduRXi9xI70SXJx33DPj4gorBIC/D5
J14JMDfshZuKhaGHSmHnCbtdVJbef6F2oki8oG3WMlCiaVr7ZlSYwXNikQfhac35
Zg8u8StZSmtN5K4wYEz6Q79ca6EN+AhrLvyRqrsVPGS0DfHzpe8lSlEGNcr45DOh
SfcqrAbsYsI75zAXxGlf9GgTqiqMjPa5kCnLzg+F9Ck98EvuA0p+odGkDr32rsT8
gaSPVOc8rf4dD+mb2VIPo/8CUyIkDv48KN9ldmWAufWwsoE+v5cwJty4VDbUF6J7
njE9BJ3W4NLc3Is5UKyxZ7TtfRVKtc6ysvd4OUs4rMV3VLtsg24qYgGkmsN/w0Ci
3qyWnEZi7rP+gqBmBHnwpKeYXtFuY91gRUytTjJh4LSd9NgJ1iK+jVC57KRl6i+A
pH4YeV7NnoOLfXa3/VfUcsQq3AwTMeFrT/lO2UV3w1dfmW8PGjNGbYF20OxxmEUC
yPyXSu6acynJ1y6zVc9+jD9pFUX34e9YRUHxwu7myPz3j+3fW03p9Ji4e4vCYKba
SzwNRAZrir1228N0+bGCECPQo0wWm1GqOhU2583UusHXG+ASV5o9r1Ww92OXPX7N
G9iFsRJJqBom37kco5spa8A7gY4Y4dihdKa1cjOsocv942EnXgZxTrpfnsW4JpuC
2ithTH9UpU7uGorLjUUMj5WHHJGSVwYODBn5zP7seoBugzlKh/Y74bXsHMqSZ6RP
E52T8Po1RjGqoJSbXjiyIjG24FE9YA0aiQOmqFaOfCYnin1JJskRrzwszFdSt2Pf
GLILWldPrB8Upgd48Yiq80+oEI76VFhn2Hif4S2ztmlAywKGDEzN1/RDYeGYDERG
biTNXcelcKMvYNcNO7JYuFl9+BGGEnfhsinDMIAAMMU+od12H51zgFimyn38Mt7t
fntTwSSMW3/DAqzmXIonxYyNfjPLbpK0L72xEB+RQCKdyq1cw+5y9/WlteK1N9nN
ZTk2yydf6k4Zmb0g2EtINUTXhdX4rRo+4ON6W3hcjGjWx5wKm2ErGcedBCRAYwwU
f4EM94rtsIQSoI/pgYgOkYMou87mX68J3RqANWfb/rgFYpdMCvJSkEm/Yd3YHQtr
0+n3bToEiCH8PVLFWVr3kSqoRX3890xRtAW61srB//TApaZIV/ezrSviRcXYmCXs
S69NIxtU88IBJT/lwiJC17hUoqqJo8yhWAsPSmr3BLwMvWaQ5iee5hW33j5TJHrI
B38XdLqIUAfJB+4TYdrPMUEp5fmdLxQ0jcJ+pkftU6lVN/0hrDaqAPsi9l0fpGLh
+jN9QGAoPD2MvIQ8rBJ5Ecn/lzSp9OjVvar17zmzGR76jZJXyvBrxwJGWI+BqsVw
AGnZszoeR7CO+a2SXu94i7wqeGwdfVT/x9LtbMVZqG1aLk0vj5d30cAUYqDDuLLR
2s+gUYgtiVyneg1M4Td/HgBsXFbrVtx4rnFqQOi0Gat6pO5aJxaTrniWcsDg5Y9c
8KvZufXcAIHVAgNVb2eIqJ+5Nf/naiBIsn0YREQBkzhYrSU6JaNKKt/17piTpRVc
3PAqlNZ3XvpoJashc5pyVXogDy2OkBPF6jQECmPQK3ecEA/tnx20M/sDWoL2VYad
QTxnVTK7UufQQo8+ua3EbI3OEECgOSi8HIYRMixRcpxJu9NCgGjbdXWLgsAMgQAG
fSYRP9r2F/TtktyaGyAwSphxrBXRb7P5//ajOJzsYZaC1m6RqbYHhjlgEkeaJ4Rb
9V8BFgeEAKOoqdsMe2hbdS0QO4q8fN8AEubA8TS6z6KB6fYzYGjJNUiXbtzSrNC7
QUN/gYFJhZ3EiE/rbDIcMl7Bff7GhAEc45C92zOW/aORzYtO8kDt9iJiBZin2QEF
DXhL7MK7P8dTqDVTVj2KBtPoyrKnKf6M/rYLP0FXA9PflmYh1OZ8l45yUPkIm8Nb
m0bGH9zWOkhH+GzpVoNjbMLw9Bimhxlptikol3UuQFE8xqOKYVETnbl55WoIz8lf
DsVSmZteFRwRSzrA5clQljxr6NFxwxhHuqge05yF8PnSlBDU834Pi4v13VFFYDEO
y5a1L+kd8wsDBhNOu2YGA2ZWj2JuDh5hEajxVC2jfW9FbmQIvvOnHpu63mnqn05T
SzZtMfxBSA/WL42zBqHnk1k02NvJGo09OgEh7ZqRHWtwz9GeTYB9AQURVcwN1Ags
ii5KT/bA5hfx9QenXUxeXgC3HUIDQzPhbMzseV9WkA7Ny9lMOt93xbCRJs9MPPMf
CWEFagA8sYM/TQx9aDmVNJwZ8UFns4xfY0A1YB8ZonDUeoTeT4It3iBo8zJdr8tU
YkrMvHnm3L+fzw9DUCy8IcflPSiqUqxjX1jAA3+nZtQ=
`pragma protect end_protected
