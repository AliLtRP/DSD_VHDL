// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
pqOzrwVsuvy8eTPKZjnOcloBIhc62VHmqK27tGDYNE/9pp7RagBrRQ4QHwKcQiZIqGC+50td+PQz
inUiOqbuuOZMR4ZvDCuKK2PAKG25D0Ou1ZVRC4lbM4qIW83Dlzn7ZqxxUQlBofBpk39FlidXphLD
+v4Dxg56WbyPD/HTUYWeXhbt1PHv3hoIOc9MdKpXXwNjncGpgb1gGghINTMTBajadPAoBzT3Ydi7
FXbbi3nvinej0l7PGxCD/YoFrWgjzfTn6p2fpVU7i7Usm6jcKS7/38ZgVt2yxaM//yA8Nt6ALk8h
yfHDWU9o7273K4XH6E65WsgtVBzhkutiTsIpgQ==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
qvfBbrzheqN4Gof9JSavowdaF6vXpzeP5cLccy2Ji86S09u7ns0RxYad36Bn9mIE591E5b6ceLCz
9azBzC00sbUmoISc7oo6icsuKZAf3dfwzyz9qNrC88FnnibwCThCpqqzQ0mfu4WmzpNb6+YjOdnq
dHIOVIbmvGzhTd3ib2XratAsSItQHTTj/n/5HsHGzylN0S18C45aEgPXjg0r0eFz6vkYPoVDo5wk
V1GyKJRfTk7LtEc9zc0BZmcmFnxUaeBW4fAVURz+7E5GFyq1ocJ8VRWaPaYe1+aIwA1aHjBm7Me0
VKzLO4CNKIaVswVIF8vjgQMS5AA30sd5HrH/PmHR6hUOkvPXZEaJH96cPAH6sjLkISsC8Tq5pqSI
FGWTrDBItwALPInpNQCbnaqBjlyjR9ifb56TRpJ4kwAUSvIA4KK1/lF8c4OgWBdOX0XdY7Xw2nZT
8nPFuezQ6u27LAInSIlJSP0RnaH3NkbBvZSxoaKJ0FZf0E9v0bVfPNOjrv7MJXxLH9luvTjhj/VH
BuPZobr0ST39Jlkz8nKwGq12/lAzcXm7kfJaGeBa6mw12BWOlmNYQpdqsv4d9v02TIytxk2ccCuK
r6Uaxptq4+HCfIAzbD1o9+hU1U8EfKYZORkGczESOseNt/ajN0j7lKq3z9PFjXCddYeT1nMoJs2U
iueYWT239E1ZZ0C5WW7Y9X6wUhJEyGUxS0LckHUuZbou7Yynb+DElCDX9Rkh0s34DCKlR2C7whwr
UVACFlR6/DUjX5oUj3YaU7ES/9U/9bnT88jgLRUWTu134v3FEhAaXSQt42AvQH/Utam0GhrKy30B
3pHrnFNFSpth1vaSn3XUi2Fy0KBtspTBq5tzkmvG6TM9FRAG2Hffg9nQQqUPo872sqAjPQOggZM8
z2dY7iXEFLMCP7+gN95T+5Jl9Ddh81kzJyTCzIIDIO3HK8RqOSw7uD2kexL9aiOdnew6OhVdw9wW
i09eie7ngQ8zaKF4sMQxIHyM4nAVvRMemcqzlDf77FOxI46WPQvXQSly1NThwp+HdJHaWPnSTIuj
r38d5oTimUUj19DMrioxaYJNZaRd+ju1smvDZrBeS7UU/kdI+KSDrstMEsBeJ/XMA44onKmxCO1o
eaAwyUfIxnf65o4yHbchAenHTzqPxEUMDDpioxlvK9IPkd/d3o2UYCgXWklUv89YazITK0/2D2Q+
IM2yRmqsFmSgLp7pcxV6AOh9Hws+a0kWAbRZZl23WH9Cx+iiOqcydJv1DDnfeHHukFlu1F7Dq/9c
Af5FzkVg42PvV2a5mk6NO/3hsW7uqb75ZQ+dbcrf1ttoCd9e/TadC5oKxQCta70rDjcnIAX/a1lb
Kesioc7GsHzOSAKFUom2yVMZ7RLUAyl1LZ1ESIcmK4ZDKtR3vQKvdjoBCLJnAQAA9g6N2uaVBG0w
jJmKzOVrMyDQev78Nsn8H1hH1hqIz+5OWKo4hpsKDHLu9HhbWa6Y8OkV3ovmUvk3qN09USHQQmyn
eHcBAYlPRiQPO+zAyr23IaX8au1o/iUyhqwJ1nZ+/G5bc25l3U9mOMfGfENK98W+P3ehhZVgLLYZ
nBcXo2Mq4LpjWzy3qKQuQt6+cLIN5JAbgXzvtjQ8MbXYfaybun3lndzeHLhMQqQTIEKxUNP3/rNM
+cgE4ffo1xLw8tO63vzt+cv2Woz5n3vNnoCjck9sK77655jEW5k4eXCUI3uro5lzfu8XgXtfruN5
/ANfZNrKSt0+FnbkiuWQfmA6a1KHAbjXmFFZ3L4xdlzsksBsv4fHSJ48vu+KhZ7uAarlgOfBYGNE
q9D+MnF2xB/BumWko+B78fWDYEiGdboj4SxYPsexwCHYWP2v427b0RD9nhDcCJ83pvOzFTq1J34t
afbHLSXNWWv7rgJo48vRrUpfkTY6n6+kVPcNB3Ehdbx8NVBLG4aTvlsjD82Q4BM2zdQYGZZFhV3m
o2MBLl6vrlNAQIgtJ3vperJ8Y0FUCIT00tDEAOD9kKFHcCm95PYu3FMrUsR2JFaxT9H+XXD/qY4p
bA1P2UxeDHktj7yl4d/Gh7MUv7EzoJI+hv/Exy/qA3Qd2ZMGuiPpwbQ1onay4u26fKNpU3ff6WsY
XfUh2R56o7C25TCRqGDbPrQyEa57d0L/XHSmeoNtJuCS+7wrsWxiTtCfoJdkbLD+SkZW2mWE/vI/
N11aVTdagR1oOkMPEs5G7roo5xTxMOeb6j5BWnUEOd6IFi1pHK0xaXzYdUfLIHyJJPtxirqVy9HS
gOvpchGHFbyekAr4yb3Ppx+MUMKQxvlyXNNB2xKFj0EW4wrIfcbgA69i91wFT91Izy1OQ9ncXoLv
16pFj/5XCWWw58HRVVvpSRn2XDq9yovm04ZuMHKpY5+vDl/nE3C+nhPDST5DdWGqz6Xzo3KZists
ETpUc0VRPWYyQbmyiwggJv7RbyV3xTHijcLznN+ZpHgMLiPhN+wlTevDrTHaUDPUPRA7a/CHgMB3
h23S+RVCLDozcnzQ3rd4ho5miPAcw0QcxHTJsGQlCOeNPQHr0+EFzjdN7DPqoLpcKltMmEK/nHzE
aG4Ryc0tjUFI3gUZMCNPZCSQQSqZ6qAF4HiKp9IwRzKgvh4NDCs9VhntNV+EzP1cEVcVlUuxmSKS
F/EBXW6OgCLipKz0Ul+xUL8SrAopUaBTC9N853spNkC7W3JV/QnMx3P4wPldSDmPbgl1AetQjA6j
0sKo+x7PHoxAUi6wXnpqQ9TBn/chj1B4qcmpbTQqC8BtqAjem3AVsZP5gXLrv4zQRyOi+U8VYmER
O4anNK2eF1UpqVfZxrE8vjnlkRkIm/Qv3Cfi1a39XJFJRWddy27I1CWg+hXZCgWWJeiM0YH6x965
L21c20F5wiYst0VgDiCyxp418CKFC13PA8k1ltOgDgvzUUBke2yvWz4X3RQ6/bOibupvn8mS4y9L
w9kQoSpsH0hYbqAPWFbn3RHD4sRWWgdawMmnXG1xN38N+YiBFcT358i4SiupWBo60LOnifo5VbNi
hmBEAnqaLe8k7toD6s9alsLhNcUsZO4bUjERacu1esSHZAYOhxKy+u0AlhwGpLilOzzzigC2Yz/K
bH3x5/FunafQSmFQB+1H+0jALd/zY921e1Bx5/SuGCJTiSEMQ4m/r6AsWkPaqESx4Q4Ks+iVlZeW
lKKToUQum0hxxVh2+Q2tq4R9TqAELOXHBwUsFud6nBp70o0DvEP1jtYvsq3SO+c3k4l+7/p17UqC
0RPCbJQ/Bkcf/mzL0lubsZpq1/WO7mDTX0lRL6sTMxgaPYMR6B1I4BVTr8q8uJWuKIMpjYME3U9N
Jb0TMhBvNai3ZL6hcP2TxsFLDrduYicxdE8lYCIM4JZdUSRTySaaAe8x5L6ueYbZrZz3CGMbL9h3
LcUqUPm389VXD01ysRQRLdVq65QoHNNKPJfH/h2799VKjMH+tEbxR+nYhiXOFnxL64w76luO1zsk
3cZdvR0SmjKWa1ZC3GoCi+0+RUmcnkbgAjWot+8fHkI8pJ+xgwBoX43cXJNZFIqlaH/yvJmRBRAB
mRX4wfzEptzMhnOrF3ZOLX/rOkdiWV7++6ERtDymEzh3UDBwiugx/qkFReZPRV8O1wCUlzquVK5q
PcjgfuLPJHFGgLggTecQE8G5Hj3H3Pv/+MpKD77IuodCIOUiBq45+LeQ5qbkzFHimqCjoWSX6KTs
8thwZDHOE1cmqWNHK5X5TOLyoRYvzzaOzpqgTYD9ASmlYAmIulOuWieJeFiaRHjRcS5XUsC3pwz9
H3ixMaKC/hLlVW8DBB89hzEdMOLXUyInM1ohFZld1MYNfDwE3mdq7cn+8WQQJ3KDJgy6qZiLbzEO
4wxGuBbFLrUqkzm7XX79b/OQgBz+tT9yhXYOrHt0wYZ/xi1WaekGK8fkAuX5f6lBwdoTqv9adFEH
DaxWKDm/JN/gZOqMEHmCrwJD3xcSjWqQWRlujCOTSG6vJs9DqOMkEvEzefGm63uhGFyIeuMen5Vk
jZbMrVtnvQPBJmvJ1eyMdmP+D4wBDjwZt9bDIgeK1qeQfYgc/Z6n6685kREbi4DK4JappdHAIM9f
kbXHMI0RW4IijJHA23LhocnW35UV9asZd4DVCnWsC6CNz3gSpwnqmlZBp/3Bt91s3cFe0DxYSObF
c/tCwvQuUx6Pt8/i0DaDUpCFIx3v+idKP7CvdpfssGP1vg5mbaXr63Gr43EWNJtOGAcZFDWKpdMY
6skJwx8/1xlqhKTY8YdWG38aNGoRIzA1LUQHkgeACpCwJCZ0MkHnZKbp0vN4DTKmm3Zi3DhOfKoG
pp8+jYecuLYXp/Slq8fdC93Ba4Hud6TGYlqbqOsJXrND6Qi6pOc/GxgA5Y4SVfFfBJcPikqxeobV
Oleb7RH+Nt2E3DxQ69x12/WluUEGzNczwUOddrxXf3PSzQuZzO7JL+AaY4fVXLNoW3nP4vIm4sQX
Cp/Z6nq/Oo8rbGTzgymt7EsLCcKQb3hZbuKkn8LI7dM1auXau6f4n5qSASMrsmCmZLMuGndfKDXA
KQSLjKESk5T9sljS3fRwDp1cgUxjTc2d7qudF3QVWiggtBBDc+r5Za1GiUC7Nbkzf96on9DARVyA
ZL0r874ZF2mfas9jkEcdEhPZoTtEXq+azmDKIq+K+ild8Ml9QcJ3kShd9YgNlfsJnvmelVm+pl9V
a72xMCniHcqSdjjOA/1f3vEl8SiFnMzP3C7NS0DH2+lCQDq3j4dZhCF+l9OqN6EU8+qSwceRqvc0
/ROHL2k8RCo6GytCGUHzSpRerXlpt3dJer1+gA3NZsmjAEjmPjW0oCUhFO/Or+p8dS2jq/lJ6Lgc
M5hXSgZzdqbttGabwhTsNpfh5FbQaJCxu5nvN6HNSfR7Qc9475xmoFqdBgVS6FuGrOhuQM1p18by
MBbC7FzMb20/BCyKVY5hx+s29ZsaJPWsXGYiJQWY3JAeOc8AlAYqZ+6Iy2qhPO66WjPfkVtREhZi
mhMYPNBV6JQwJSXIeLToRMjXmCsuVIaU9+w1oKMz9y6/LKc3yyoOwDIgJ72vh/emwLpleITUFNeh
MGYFcfJediV8SvwboRJgyhPZoyfPWb+0P1IQ19llMc0SoRayc7KkTzZAPrySsdni3ZMIuSHj3BXF
NSMv+wrYCaHJquLvivi9nu4o5t8axvLqSOtCXW9STE9JB6Vk/Xn8fSPst2ffIZprH/Gj06W/D3O+
Sl0WZA0ITqtLmxt6FqcFzZHjw8WRqYTG4Rhzp3TCa7zmdRevauwZxvbtEQS8w0U9aXhuQ2n4ic5K
06mLUr6JGbFtSDpXdtLMFCVIAjoVEYytR1BpzQEKnsiGn7Racw+MjA0DIJ2nARfc1wG28uk+jF64
SJ/StuVnSlmhDxkcHsDtUy8RRkmVQz1NLqP09FowlcakFPkUNNy+xs2t+hhuOq30qNxu+4nLl3C2
cmDcUonDLN2x2ieWdfvmbp//qtNFtiKIdBzLDby7VvQOAtWLnkpRXQJ5WJPlThBjqSXUwoYzf2/X
ZHzKMpTh8CIgGmuN5M/UszPYiYet3O8/WDcFZ2AW7W+OYAC65OZMpnitPjg//Ec5poPjFB8UsZLC
MoBn8/XYmDEbVNkuR4Vd8G9OMo+oj2wdxsQsNchFiWlXcsjIPK5H5FjOS/QJlN920LG0LUOBVki7
NmLHKszicdAcAEQ1CY7i2+7fyzbwg6NVQtvQ8kIMA+/shjWdONlksPMwhAHqZxrHUsgjuGuXuz1u
+FA/1A3OCvdQsAm7CRhy0d014jwkMS0MmDI1R19+X48yQT8ps1309GNf0mVKS3y8VyuAMCFn6XKI
BSfMNK6anSy3au+lzsod948Ag6VFzfYMSQPsXNgGZjAyfKqpxGewXNUQMiqYCFHEqG3ReaxElvs2
84JJguGm1A97MTGr1cwVgTvuzRGTTEOfztWk89V/xDPw7fWqVtdi3DT4BuQwzCO5x9b9tWFLc5Uz
csPGV/0s+PHFTr1df68J8eNb1MwGEobEwQ41vk50R1Ys+gdkPSWNm2TD2Obnkqz31kAhM/Syhv35
tJFUWKtEe2bBRQAzW2wWlYLT7GS+UIdYFSHkgIhQLfd51wJUQFsHUW0iUV04rbXKUglDLuOSSjz5
yDkdStUkx86Hq2ldlHHCOc5JgD8QE5M+/dKydXTvuGF1vZlffitRfxwVO2J4rDgS21j0uIppp6YD
YFrltCZkvg2493Bf5VMZutpSI6yEORr5VFXzeRZnzvolP/1TeETSXZRpWCOBr0gkg3uH8Uf5uw9f
rrE/LrNVjz2Nnff018SYGZ27/dAcCix/zsAiurLNgb5WmLX1nzwAeRv4sDMiYblJ3dFWEpVk7py2
L3YdN8bi2TWX1MPN1BMVzOaqq2q64xspPqzKCHS/656rBPJSRSOWsIg/Of0n7vrOhoUP13SVF+ZN
FZ/fNMT7AMiemvtaH5Rr1V6BRG0DP3hwf1c+GA3lowB9BYID09RB+6rNuYdZ8TZw13k6SqwfpnFD
A4AtMA1pOXAtsgmDFzrOKr4zBBcneGlhH0qolizT/EppJDxV7yp5FR9O7FQTT839DtWaTE+f28T5
NaguDLJtHPFE+68xNjVqBc9P08oAmkcATOaZu87xqfOiKebvPY8LSVMSxm2iuX6uRLRWdrI+p8e0
dBOtbi0fU7D7hIw4GOOsrICY8JySJTAYwVACI4ERq0AeVNuPvykE22GT9os9Oe4IkEVofon9izv6
7KF0tiS6IyiB9uIF5UJPleeeHt+uMXyBV7LFwRnDXdYb13VW7pNiQss/R/m5CfyOSQMI667aJoke
lHdBcE6sNsqxcV/AKltUu2r3R3vYcWBFGp3jnYGvQtIkG671y0RvEBeuqyto2Co+BH3fUmuRTBY4
XxmtRobqNVUDM4X12sGmeLTvNWxDt6Bs3XXfdzpTqldBcaWBXKLlQz0F0S5SSaPIGUlbouJADZRW
uDXNFxC5Ae3R+CvEgbKjx5wZwDXuEWQTHRax3L1u/417MWemFoLZ2rwkxrjbGmCq66u7/A1gHT9h
sGHTFevC/ES9jWHcLzAl9uasw2jsUkqdYuFd4Jz/aA7IL2+VTZxhyi26wiUgdVZFH/DKcYtPpS9/
28vppGsxRGsaClbZxLW8GoFjz2e6nMhl3ZVTbqSUYpc7vLlL3c86FmWGtPnDc0BXEysd4teqbg6w
hLIV2ZDfKM2UoSjj+JOHUGhZHZdulmZWaA==
`pragma protect end_protected
