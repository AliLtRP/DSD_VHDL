// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:38:24 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
RHiXYnhkLWBocmHn4Yt0tTcPH7sPKZI9cR5iSu/GCFg1n4/fTOvtlSF+740A3Ogr
dc+4jX9r62EkVHjoxh7biSDTI+HgtLo4IbAfeaw4fO4Y6S/ZTYDc+H4A9C+iSxhr
xVdphsW6ZkuQTo3GOUgb39sxuzvLC/ZU6IGxDSSvXTc=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 11360)
V7lDIHpyPE9SpnGX/Tht5DZhBqj/qKgOWpGmlARVRbz6NFel8WwtiL3TcPGgva46
71mItpJhkM5IQCenkIXSBNbPHNvgSswFWEwQcjOTrVewn21CLGr/rwSgqHni0lru
Xl6x4TBweoGGDYx1MfDngM0KiGOhHMIhHSpr85ajt0A5jhDnFH6Wju/THDGflyGL
kALq0/gX3Rg87hHmdp1ZIpoqQvLXEDWIk/igQ8fxVFoSgx31NIVmCIa+h8lOUd2S
HdH2TUcxVSi/Ce//vxKbwBUgQxImTPiTmIZ9SxJsMxQTWuTSNPjuZHhV91swVz3D
TNE5li/gF80GzgjkiDw4glEe/gqYtGfnweztSHh462fxQTRANrvueZQ19QWe+AQc
LrZydieHEXaU6fn6X1LPPg4+Edi8n63AFVkiCxvWpLl5JPPVjpWZk/szCHNwU7Dl
jgOr8kVHz/3DQMBRriXUdTq8mqGiHTLNxNyIKro9ZGu3dLvv6wZyRVbEPrzv4ZHF
0PMWj3eGNcI2GWZhYM0tx87OWfWMW1M0Xg+Pyw4AgsY89MUkcfQ727VsPgaewiUe
mMslMxkJ0zgjvgyVHo22Mj5dl51j4zzxfC8yBFbssMSYc2WbMrAG6V44iQN3hq2x
1aCQhx1m62KSQOX7MPujIGWvil/Q+aCow2+ulQhROxPX/B3fEzmCtjAUO/zuq5i0
LORv3t8HPAGBHVSWXYFAstWlLdN17qWCj10AAg6+5yTEwYRvDSYT5jCJC3B2EBgX
xZ3Aa4cdVyvM5aMO2f6Xy5pWeVxgvxT/lYXKSsUk+7i4yROw79TdCC7mryTixwlv
xva8ibA0JxicCzkW4MFuivwTBLtzJVNmXW6hWxU/gW1Bvk0Hvf+MoSxQMLtSug79
JufHMY433v/DVNElS06pW6BM5J7FwFLQQsTMhUW2o3sWkLdCNdxRyCYci5J8nVX1
biJ73Be1qZuRG/j/CSWOlb+MIr95CDT+XXNN5CQ/wBwLuBClFct3V6H5IwxcdY5E
nfQqHwd0uKKt8F8E4wNEozf9S37Iksv8TPsnM7two05wsh5dETUpYBur2UiS6jq0
Azke3zLPNpad7Vuk/08oSLPaHNtDKVJq2bEskv3lcn82oa/QnAsPvAxswIYuBEh4
MiassuueDA+12zLLfyttYoAoN6JNk40Vluuevny7ZP5CRrNQjkuJGwDizdMdHL4v
vHb6nzIqa1DffSuhdK2r/QqSxPlNckNbnWbU7/w75m5sOMaIpI1Ndf4r4Oaimki3
PWQXXoMOH7oHZuctMcfhliagCHGbh+gNY6UNP6iVU4DJYKSAtK8xWNDePDAcx/HV
5jiyr9lS64DwOT8zKnSy0Y+x+0K3wYsntDzq8MvcRmlwMkp/+gEuz79CjGNptRS/
H24w+9ODyfkumlDlU6n6nb/LVe31TSJn9zMsDYcHgIU1ApLKWo1InAJZyBNbZzrs
xaWl1LxMKpkVcJbQstJYSha8sIYH+n2JENC7Y9Lum+BFmLKhltMUOLFKbwEIB2or
TLkCIyPFZr0jU+OxCTf/RUg6tj6c36BtPfRfb9hVw6eAbWOtdoYvlp8hhdP434sh
GxBfgCyqOL7cVsDfB3Njtjc68L7y2LXdKmaw3cUhZt6znFbLY3I7yE5sTvI+lVoN
qEin2CBbWpv6lUav0BMyjsgBHI/sCD2jI3SkdcUJshgx07nmxJjcIofAX2/+U6t8
tvpWA1bsvseI+9i0E85qQ/0zxe97qB0e/Xa+Vk78ulktdXVGQQJsNgQK2EmGOzfW
yD9VV48UBp6CVY/C/PWxp33J+4SrDkLmiQJrBfHYo0P10ILLJCY/c/8nn+1ilZt4
0zWYoT3ZRVoXiBRc6QdqMh4tBFND+F91hcStqvZ+gSTfnvNbyuyZ/tYeWP2BJ9D/
qcI7TQ8CdEayHRtSM3YJZLy8DQbI4qZl0gf3KKBO9CMv5/R4Nm6D2aSUKtjNeK2n
NvyQzP6LrFgcgI2dCLvNFt0GkLM1zhZOoIpUQZ9BFq6w5VqqLQ5nyX9PHRenlC6l
C2xkudKj8/BsMSI0H3jjPIRsiL9Zu/cwHDExfSua0tXne+2KKmbfYbbjuiFxo/JY
xa76LoE0FEY5VE2nE7j2RpRcoEYtAhOkY4z5xa0O2CMt84UVoCcztgP9/ooeKhdA
AxYmpoMvl3k1bEo4eanF5kIZCnFeEKGW1KpbiUPkK653QEScHNOCKVcuLcIYBtSZ
Pd5Nrsq+62jPIvpwnPiAOe9r0rKc+XEAmfJQFofMPDSE9sfAER+1p9h3YevrOsBn
EcNUvBfl2HVL+7wUyngjEttAHY7tSu1pvX4oD/+5Aw5Jp+A+CeyoAbbAwjAtv9Yj
HT8WiL4qg9QaWAI2oYEYFY0/FvrsOOx9CkqTlAunpdKj8UYSn3W7Nl+bMNx+Obvt
/fdz7UYUu3Kt9qXdoPScWBuT+8KIwlsKCCmZPtdmbacdxiuVR/WiUTGwoG1flN3J
iiKLSnEabgrY694nFfIcfnqmHwiPbAQJ1rwl3Fkm3dOYykHjMKYu7dgJfD+kxIoo
dQbfI8yg0KX0AcCRYbK84KYaGbWEj/74pfxsW2Oag/p2FHto+qFnckJggCXGh/EU
8qTDw3FjyjrOcTf6BrnAeE3yfoov9Bvg4SqXGaWx7nhiFHndmQBpPhpaa7WZjrP3
gbbo/FvsJP2WIVFL6OvfQFtbNfoqs5PrQsFDYgp3Se3iRWgvQS+TNT8dBR4V1TB1
lmDm17CHzf4nTcT/StZOrT8bHLbyPcJrCidHH6N+zVeceBBkyRJRR0dvLbBOoeZU
StXmIi4kiJKeQHwElvhzAFFOgfDcJoEGJ4cV1nZpo9TD4n30mtPT/hmkApbHgV5M
ndg9V+JLIzO96K8gB0tk9A/HE+dCG3dZ9xFsH8h3DWC6rPjwN3FOgT/I8kGgLPG/
jWTCGF/OTagntOeWWSgxyijDhnvu3TSpraHvqLRWDj5fs0Amo4NttbY483XorN8w
ascp3oLgvWmQqLpqGER/Rkjf0MmGoS5EKvVmhoV9VmX3TclHNMc0wFph+h02hMP8
wda5gCZeV3M5q3QQ/dTB0aIJlE8eXR1WpSfkG4/mOzarsQhi93SxyqLkIJx52kHB
UWBCZ3YqZiA+Jty0cw2OODotbQTXevKbjhXleKZk/Xvid2fbogEZVbHU2JtgNOel
MrAjYfsYHck9/K2d/LQKDt93ehTZxn2CFR5+tvjIAg0Y/GPLcFOAKRo4qO4qbatV
KVB1PEo8rGs26cVnSgIenpIPy4SMf7mtYHAkXF/5RxEbe79Psbh1OHX9WCPShS7m
B6LqUkouWE7OjaQEMsxWInLyepgzWzEigKBnRZ+8ccYjoPUbqrqSLe3swrdLuy8Z
DptqcpkTrh/mQNbRJywiuyggMlpYBmmVLdINE+2uhybVt762jHwhrDo1HM1feYgY
IKsfkQfSoIob+RxIsn4GTqx4VWnh1z3F5l5Z1UF/0TdWcduuHuPlasnqsW4FFaV6
fGywHdsfaxvAwC0ajL96ATWx7YGdv0zA0PX0/ifE/ITxFgEzdAJ1TThScQDBCxTP
t+uQfqTRVsJRwhfnnBL4b20cjnuxJxVleOJvar3L+GPRIybIU9fhaP+HBMgzEIkS
gwRyrzL5JyGtKlMusVAVeoHOVTsgoNFvYseIMk7iz2EEyhppXvlZU3LecUdypGbC
FwCl61IUToeiPKm4gnZd1vBZCafDKBnDSBQxaw6y0FRjsHqlteu3UuyIg4L4NGrg
5KmvDVCwzjj348PZfz2o8v2sp5tMFGyV+3SVpt2LCBoPWuesy0JYtr4l9pSAVb+i
Pr5cSbdeiQmaxxiqQ4kL2GEHJ0c/6s4rc4s/BKLybamJftVqy51KWxkUy9rADznN
eJ5JK8p73x/rCwKjhJrriCHrMHww9rMDg7BExGOiXKENdEXQkth5JWGqtz19EJco
buXgroS2ntRziWDUjdQgnkETXzrHUNErSn5Uf36UedU/xPleK2yyX3sPYX/Gand7
O3hXeMRTZ3Exc3p/lX2xJ1R8cKXlCGn3rjEIlwrfiv5Pyh9+6D8hbflszj9swUg+
4flwIk8whu5OMkqDSUsJque907VQubF12cEpuu0wzQmEESp3TtTwhOf8rjHGysfn
qDT6RZ6KO66UC9EBLIR1blcVbb7mvuVxGs5vCiyhlYGdRl5+hzetjZHFlDVU2CBQ
ZNNyNQMhbOO1lTcjLR/t2H3FfNFeZmtODSDInfk7DWuwxJ7zvmJ8nJAM+RnWi/zg
xoLcRMSNLq5D1IwvstnR/ST23f2S9j5td7DFFYUz+7MWg4fBQ4LyToSMBXAA4ksZ
Gz9sCYaNe8J6vmrh3+Cf/La9g3U4lTVXjvDVJ+s0JLGpJQUITFlPoXfqJvZnKqSy
hc7T5814Z8TEFiJy4Q2PPtwqMeKcBbq5ULzTs0wozZI73pJpoAg7FOAy+FTQL7xF
XduNAM0zWD1q6t0QlJXZ4nrXZ+0yugJhMF8bjFul9CVhad0B89DWFxsoKVhUVAbu
Q2GXn0YmZd6Ulu0HC3XaqzUdmfl3Tv56LFHEfGyKLzUGHNXsV/ZaBbUUehzgCPR/
IUCR7fqZo6Q2E3mTPUsIi6n0FpZw1gX0QWKJl762K8K4+t+V/yhbnbIX1PMsqWU5
AmHgzgfKk+L6hR63u1y9T6Bsl6GXIBmEvU7C+4V+y1rAdI+robs9yKuZvxd+ynMU
4K3YfGaMYI4HpsgWHArsoYCtZvZou3okjpDg5ZM4TqXoI/Uk3KkRXyUncg7IfaDa
rWrjlhe/N/a+UEwZKsFahTQVWseAE5gu0Yifl1pQ08PQTObDu9O0xPWV43Au5qWJ
bYOVuUpdOS+jn8L1I9usJrSS3Cu5EQh6+79ArgsLFhmGSM4kAjkt9b2fkf+3Lkbp
VwL1NBKoC1x/87OCr0mGL3H92JV2nZboqblZX1KekT1JRvZPdlGTTo4uLTryQ2K6
RWfAWLI9NVWmhqWLwtkIpLDvPWSpOxWTyLv+7yOip6ZUFXsaviukecABZWr2NRFG
auC/WEuai6ulkcEQI7/PMOCpzNum8DgD74eLLyWhyKVY+nZjhAo+MxIavHnJPjQ8
TjHlt1ORQXbPTpPa2xmeNMt1tDdgm3xni3CPhP6AtdUiIe+vBvPntmCzeSP94xJI
V2HisGOTFxbMyKA3ocpB/GudNrOfe6Xh4fDd4gvLfqBVxmQqTcMQSe54zUe4wKzc
A4+TtVA6oqE8/MwJUvm5+1GAE8oo3sFGTpezlcJ87MS+0mRgMLFFES7ZpO91NTg3
vr/p2Qh5cKWCnEZPkx3ArZZnmDzKpar/KR6uXlBmEBL0Ympypq33QFzTV476zaME
PcARiawTWtEZtMmpv5WvLqwR3289xW+CkfUlhkQWWzkr5SroRBPZ3+DY8ijZGfas
HK7CCcIKzeL8tGooBdqDMYenQu9b5ee5tGWcMKBinFvO5I/qpb7K79YoKahLINsY
K974Ct7kM1mydX4MMDo+Q/lYWgKpQPKy+1RX4FVOwDFt21SW6KcwT96tfj0Q+B4i
R2dgVQLqtaHEmJJBqtGCzdndlE2ZHQjWQ+RKygcl3f77CQSDs7vbJB0bZZ0gq9g6
WcIAYgFvtyn8qFcB50kuRAxqBrwQisfaEG9BvPnKyRWu+s1l5SNiDbmwLJuYhag4
Ovw+pI+sUh0iBZnOn287uuoa+xEqUc8As4sInUfTTdkO6CZFxlYIjH/7qNY64lQH
a4GxpSovOjlq/w6XAt7Ra24KCPHkUywCpj4pQy/aAb5phHPlQLxxU6qUMzZscDBC
+xJ9gJAKXMmQUwNdVqCsiAW5zsFM6lYOSyYlQAwxnFRvoZ/5UIgoz1kGF5rkI6KA
MqPIvh1r9xsj3wppn4eUlUtaqyFNRVXyQS+4ts54HpQVxxbeOYf8HEXTDd6EIvm+
eX2PDLBRmZyhzVcanQbTHNNTF0deR52531B62d/v5e/g0xPDt1IUej7W1soH/buJ
F+kdu/7gw/LHNqMWiPlk2vjJ3Kx7z1Qm/bhEuT1PnEp5z/8AtAysmDWb4ulT1cPC
iV2dK4vsp2c0rlg13ziPUAMEU4yKcB0I7crnqrS1HUXESv0sosaIfxekIG7U8gOk
txp43ni4VpQuvNiLwxIJeFL48H2EoKBNj0ZVj0A0bEDS6ExsnTLGSg4hN0MyuL+u
5ko76ritwiNvj2EMgF2JJAX7mshIuuIl3m80OgikQIJPdwbXmLKm02AYhqO7LhTj
z3vVKyd5yCIa27AP4irKAI/YM5gIXd2ZfQDP7kQlODBxNszu3fwLU5Xom1EoOdqM
oSlb/14V1ElLkYzzDx0k56xhEfJ3WEVOgL7XC+xsrF28IdHVTgaXpiu73SuHXUl1
KCJqM59LNiylKYP0X7r9p5KNDI0olUyJA0s+1aEV8+gOJerA9wmbiUqmLT+yfuvt
6YwctZ7K2PFhDhlV1a/ct5fNMaTawDq7chyeuxyObsk8pMjam3DoXcvpr1Eh92Q7
PtLG2PHQN4zm4jOdeXX2bZncoExMUpOVSq9v6GFqMv360x9GdtQpT3lgI627a3nG
whVAYGoguFZZAzr8I7E0xCW/bf8RASO9mw3b6xlPp/37flFeGGPAjTUX51zVKZ8A
+g86zf61cbqXfAQl/qCRwtoWTKvo16IPEqOgZb2F9URcPiP1ml2pI4ahQzIBhvLy
oqHQ2GeDWU/OHN8fsdQk975/YyXyMLQAokEdONLoD2X4YZAWxcy8kWntF8Cz4Tyh
jO3WQDfPaoBkZf7McfqE5ezZe7l0SOUMxF3aR+r7vW1ne+QskDH4huu2MzRZ+Cnp
bWJ+ga9BWZDzyCtj4tJLpUyt4wDDtlGrnE5qfHyIvSTy+H54KRsGdbFNn1oQMOED
NvQDBwpE1bCIKTAhtuaFGBIt0ilFRyUFCWnGefToOJoe+gF+kyRSwnNAMvpLXRLu
pxbF3JtjWLtUTb3XvYA0gq1LTu0bfFBH8NJdrcwbOcsjJaZMIKfDWWegzgY8p1kD
ECfckqMXm9lEaAA5VjVf+F2Y/LwL+imaI7pgJ+XiN3z19vcHkH1QU63mOWExO1+q
83nbQrDi4QuWNGFHaiCqkTS+JdazSXTC4c6rftvdRoocu61tSv4WMia38SgEF6Ti
u1Qu19lQU+lH8Tz9yhvLu85VqyRqyr3YZ77mHqUIza/SHOI9lqtLgdSVHlJ5VoCq
0U1IPqIDPDN4svXElYtJiZ6W6xDRx450lwCq8bY02qi3O01HbdJE80FcXngEMsSx
hRyQp4luSUc/pRPk+6psmubMcrU4sGTdpkjDJpmAnS9KhY6ogy5ZjPg9DP13+gcq
r7hHf+9y3BKjf7wlDFhd83U4nDOW8pNIR0pKDdpL0KuKjy3VI27O+H2EJR/b8PRt
eapoxZ/LPMknPfEeongZBEPuJ2fzr7L2z9Iqn0El73FXXb3xTV8/4HLTfwlqfkyU
gId0LzxR62v2n2CLrWfccprUMw3Cet84b53B7WuDBwlXfdTDqtBlBUe7j6yfAV6D
OO67yXRzRAa229uvFNwE6toPehtEaVlLeYtfjp6AAQH5J9jNjECVFlpXtKt9fld2
RYaPmhs1HwyOojptl33pDECUojmfcX70Kum+MvrpD73NMxiSxkyCCMFpkUZgI2YT
RaQQ+HkiiN7mjJsOYrDtmWiMWUMFLb/okMsIW0qXsG/f9iHf8U+Eqnns77pHQoaV
HRMnW+XpuanFRonBT4zIeud+hF15tMl1QagHOK7mmHzo1su1VhYDvJqDdrAl8P3z
hFgaVqRn+ILeW1Y55j7lCWQi2dnK2KpPTTFsr+pLe3Q3VnhsyEStgUl31iy/BBmU
miPquwP/q7+BWnBEdI7VW/SK991s/hg6lLgNNYlJ8H3SjcolKBAEdXz2YSWZydiQ
CCYrVhl6XYwxKPxAwO4FRydpZufr9kBVrp8TxwXFUbjH5L05CaaYRxUlFOyJ+oy/
NIxFz3bfVwITcmfkd1xMxSO8uHHrdxAAmG3qtxJiRTp7Zn4CfeYpCg2IVury4Z8t
T/uo8102P7HFbsoi3mwrO50OKn6sQJGq3O/d9WpFtGaiStL0dlOLkslFbCh4RlEC
R4AWZHJqH+NbsYHaQuVPeWn/3qCqbpCX3P7j2AsGVC4vM5ZPwXH9/XKdg0LFxWnG
683RKjDWl9akrly0UsbJ2+H8rLud63gtEqDblW8BM0hM8gQ6CtUOC58Ubp0eGREf
aIzQdYfxhEckJ3aDCSv12mwRwr67OlpjwWG50R4SiskaLCRt7zbwMUKyYZj2SSuC
QWcIvBfY7QxykhSEMt+cXD/boOdwLBe+u/e4/Lr9l6+FclBj0ObXEJJh6FspxYoF
r/imOctfJPiQA91p2DxnesXL7NJdHt70kL2a392ekXMQP+CXsgccDMQNYAhC4bgE
PJHyebLhzF8MFZRzjrqYG0ej1Z5AImN4kETpqgNyCnfn6tlEfOgvvyZrG3NdKsF7
Dv8fc15wlPiwGzthAs4gVCwLDMjZ5c23mhz+e2QhrJw5YMEPPNcu8e339im6k59i
1t/XxWnsd1Gb/S1iK1Kn1fazM/Cp6VEKqOiY/inIwwz/3b5kuXN3vYEVIl3das7r
hfgBSDEmW2TcOjVKDlNoJ9Uy1O7TwKGnacV0bEPd5vpr3wxQwTbFMt0b7LvUZZkz
5DLYbh3h4Eb7FQ6C6ba+Jdc5+ttv6DqmsWHq0hTng5qcfMlPYv77iYvkub0iNd6e
ep0UOtyLG1GOtvPajUWLk+G6T22W9NVsO4gIlKvoOPTfWLaBrvi1uHny3pU1oDQA
TPOekPJPkQQIWxq5yCaJixcv+K1XkjpV8B73PPBD5Xl3hrTshDbByBOwWkvF7Lct
EuH58Wj4bymUEKseU+l6bS2UvINPB/pf9Fj1KZreuXvD40kl8sZLHyaCwkLK8/rD
qe3hxhFawRk7bUKCvhL19PPd6ujxiTHw/7leK3Y7IZ03lAES9HrT5fGjpF/hGhm9
Cl7BIMrvh7nFupUg1MHj+fJ+6/WzPO73pYK1kkvk1GNI3d8xOA6fVK199wcbwuqg
e+z/m+0yw/HXooZ45k0+RJtZ+G42QG5mw/ibNEV+3Ek/mUiF4z7F5y4uAnyTcwjA
JoxaY43v+LKVQ/vjyHfmpA3iHWCQ4vwxda6BkyuIUYYs0r6VB8iXz9sSXGrIwCOt
BSN52Gad2fBkVG7XSImPEvvJnFwpWRqVxTB8Hb0vouc0HUbSWdh0xGZ8DRiTag46
4pIYdfcX03rDeaVJ6bPJIX4ydPCLfFfanhCMmjnBKpZejSRnz+V1CwYekCV2vz4w
2z8LH7PGtJxtShlPDNiQcv3prRbWdeUpf7AVMavohT5xgm+r38HFUdBNpi7eN08Y
oD4XM0Y4FMyKp5gHY6kt1dDJsrK6Qt0HOrwLA6CufeLxswbAFe1eI/G7tNzrSMJU
4zcQogMSlew/aKIizm4r3KSRkfU22VezrdRvX7oOv57cdeXVncV7W/5yrabhOkmC
Z2K2TikJ64v7KYKQIcZHCjtmjdsOLdGv8bq3SgsSurfN6w9TaVMFJGfEdqsB8Qfq
UlF8vMGZEgRZAh84XorcxKOqaTJ2Yfo9AwEh75zJeNzOGamzRvDlx+7V+0MlSE04
slKhQdaHbjIXF1RQDYlXyTi1ugbEGxD77w+Z3j84OXVg6hDHjRKbUKsc+0xMdvJz
Iom3++LI7i7Z6D9qJgLQKZXnz9aIFQQbrMdQWK3SJz2WFh7RKK5eTvPkA5vkgPlK
q2xqSx5WCBSGL1KVXSKY0KVtcoq22nZ6/tIlF0a4Ow8nWAcaJauAZXsy2LQy/uBV
qOOG8Whp2t+GzKly20vPpj4W2bhN6cWk8YQ/ioa2GANVVRA4QHeXiUclPS2kzxfB
m8vPcyRsrwO3L94T3fRbW+FvTSYy6SoJRT2H6e9JUPiacuOpNMo2+DhN6sUiH2Ps
HZ6vvxr3jXJpq2Vej9odArlS3cycqn0z3wTLWh9JvRt8TLYIf3UuVrirVq1ao+Ys
gSZ6kqfHWrdu/MvvjT+fJB4liQ0V+V7davSzHe9/Nm4SwisbS2lIh/PgNI+pZvBR
C2nfzz154s5Ho4XhwnvjycA6uoJOqhm7IPbeJwWN9yRJeBpXX9zxBM1y/E3FmM3Z
FlPdU82erNJBVt/PSdgsOmVdgdh+wLMFmulZEuEcChNHaZ8rYiE2buWthqGaFYUn
M6zccg4rtaRE2ZzzPwnOCjcWwFmO4FnrLMwNGmO/wP7oi3MsdTq7z6HQHsScR8Oe
AaoUsoqekyCfy0YiwocVSrEPgg5t5jQl/NG/SN7/gEPe2W48Ttv9s6q1lBHlR9AU
DH2+M4gfaW1pe5oZWvf7kPT5uiNIzSfkqWQHBzZcb0M5WGyd8TMsMh79fjjG6EpX
AV6ge4j+ierMqYJ6BFbqE1ITmvyvcWVKua1N0BOeMLUMyExiG3C2YlxWgRmfvUST
BucWGtwNNNDNJy5tZcUY8HpxbNJw8zSxbqEBcnuCaMuLhZBGOo5H6rxcXZzz5k74
Qto8I4/l8xwPW2h1dGX85pZ47sS2y4HtMP5ObYO+G0EaTuUmWgEFCh4I+uk0je7k
TtRO4zkgs3CE8jJjgL4y9bD1cIFOsAqoox1QEIrloeXY5mVLf8BC8em5gbsK8Djk
DqnwnSFVSv9jWgAgSGF5M6dTIVVhVV79HryQrsiqiWmlLmrAZrR+Z0Np48PcwWZs
HmtQCPknKDfJMiAU5IgZBQt8d3Eqp092jUjln1pO4CSGTlSz2XoOpatwVSL5ZMpf
UwQhW9W/BlvWmmKwaY+BNXoYG9YHiaYc4/GGB0MHLmrelxd2x1IUtkHuo+iXY/wC
kEJymj/4TiDDvKpGhOWNnwHpEAd6Gl4n5xsg9WwzyMax6ND5VIT7g0mxyaeRHR5X
bvWZobvAQ9LQytaPQ5pgS+vXbGXvmwSVwQ7w4DFV11yIbP3B8Qmub7q23RnpTsGV
Ump7yiNd01HbmvyZIk8o/HOgtbCtm9D3+sy6kqILCWgvImCSjjThOb0gjcFtGLkZ
CuE1j3MgLCBy4SSd1trN+EDuYyqnT653mb4cZb9H34zdyXcqlFK0xfKzdMo8de6t
BEgAyFd/zkwum51z1FA7IPRiqzBxNdXRgfvAdHtPSRruzMaD45A9leUutt7Wcsbh
NcXZdzoMt1YTJ144L4ejbC2f1MQAkLsoxCfGgJ2lE2V4qasr/4wwy09TuUy+uJt5
IiqCJwcQDOaA3LqumPagQRQyF5Fh0odkzU+lKCEBznMgnEpJTEhF0I6OY1wjnw6b
GYyKJkG+bwUk0zDCmCMybr+t2P/XOWRnXTwLH46+o3ra6dCI7NfBu3DK1j5mVLOr
whIPY/uraJStRsGu8K8a+3K991USXik3zc7VU+mg6stutlUtx0CTCvCECsWwADo3
o8ec69FcKxjVF9Z5sCK8sxq6Zey4DNU4A4A3WWlq2nejH2B7k3RmqsBJN4a4GM4V
KSVEZvC2JoalTFDv9E/tDk11aPEDjSFaWhg+8U9JVFLkL1ov+Mzzuobc04m8Njb8
xHmt4M0dH0dpchzmgCTeUEsFELXXarkiEik8fLZMDaZT6//PMM+BQPwqUi46HBnu
zkvSPL+RxUJW3ze18I+sOn9RwHxfmxG97y+bHjvp3SecjCtt7dTKx6N0PbWkx6zX
QQmOMXCv8u1LhvOSOo4YFCw5y6AjeT3LLvjDRY2AMCfpjUJQ+prNC4JacUoNCwDF
nDzvH/0FVX1QZ+iKorUyLdHSTCryLy3+kJ8ek0vfkj8Zyqw+TTs3X+E+BsL3IPBX
dxdjXd6rdUtCnnfwnKudzrcmPplInoA/WSBwlOfwQ4BdwFBeRHaBo2QL1XVXGaY0
hXftJ6KNuWKFbhgeGPDbu4Ok0WSgYGNkwh1S2BTkXlf4Tc3hrcXHaAUuXoOfDuXi
Y7cMdzM5BF96U2rRXyfty16B6umjZsqqGCiC2+YdMeYaMFwsUlYN8rjBqF6H2Erq
2SIbIpOjV2uKIya6UygvbAIKQour9EIGWBCKfEoECFIZps7cuQx8LoEpdQs/Asmv
emOJGaHyk3X4I4Wqyss8TB/4uq4K8YvqQKET9SVV28OMgqYEk2gxQwgUGo6AjDxI
LAoeTQlIigOhCMGy1613kSGuSoEiVXvnRuX2FDzVQD9/P2zpds5wUsA66IxAhEfi
2OtSqY2XCAlQNTpOGQiHkoD8/LuslmpM34ZM9Ff2K7UHS6cJlLRqQ0K3xRaMW11k
Mk3GiVIe5yDceEmjexchrogbaTTZ8vU/qNd1aRMk6+46ACvRsZYvJVDE2Ip4tow0
OynQhQwI7b7dx9POGYu+FJmy3dyWYSkSObl45uCvNUpn50T3jNkxenki2S1BKHbN
ptSG8cR/1tHDWDKKrD/34hZbB5vDkgWskMbogR+R9Ey8W1PK35lssEEbBj5gGyOK
7Ogsi2uhS8PGNptnoCcHaGNGWf3uiu5pGa8thXAC/+gn/Dtw4YOEt699e6L4rrPK
UhRUmdvyuaJ+URTnHksMl2IKrzp5N43/7qF5XgKFZ6Qqc185akBGczDmi/KdQKgc
Gl4vDhTItqjtzfnSQ67Jux7nxRWKVO3DmMSi1xZVlly2kZMBHsNsVNEzBevFLuaj
KiBoFGKRrRp41/8PV2NWqb/x9QX5bmTLH17QGW0RFYEWITSfTV0Dk+82vyTK3+My
QHzngSz83JKfTw3Wr2xYnoHFggriBc4uiRMsTlTJUzPjyTiJEhmp0+O/5tozrcy/
qJzBQ0Pce8Qc5NpZjNwDmC6aUKvfuxgRk3cyQNsszHG2nK3EDgzhijW4yDc21fuF
85g9KGP3DU4jFWhUM7LntMC77dEYLiT9ToMBEi8KGDUJHDrTlxKMhS5GwY70xe7L
LuB6VG3C2/BTcFM8BIr8vVEBStnTi9J6uyxi3SuE8ZWWjBk8PxW2hCq4asDTRUD/
KB7AwnjQMvrQejNRWoNbCxOAvBw1ynco72OR0rNIrC9+WEmlDoH9Ebr42LbcxhZW
KpkgK3Ewm76VkHnVGZwqWT+3+eBt4wHnlQhMci3+q9TREj0OAI1O8ECYoHPOZcZl
peSYBYhpRtRUDd25I+Swjc87WB/RA7O5yFTL3XtyGVyQvXrIxtkf3/otYwPkUJrG
4///No9wjqEN61Hudhfu6q3r8Jl7TVL57YAMiUvjHMfyXvikfGWOE6S1wu7QAVz1
Pwfc3UcrtoVEDyL5MBsSjfI5nNz0CDbzWmc+qONrQlRyZ2rKxVezDzp15Ju+frte
osyyf/DjCAt9FgqqM/lgcJPV1U9m2AAP28k7f04kdJv9kVcVuuBYvg9x8JFQfTJp
SKL7AUEFF/GCUD/w6PHV3Y1R/hIMpV67RkQK6NPrMTjG9ZxDhkq6GbruG+GxpHgy
4b0DN0sHgVeE/Khs4eZDX03XAa4L8bqssSSRmfggXpdk4Ihr3qDFsjEguP47XhuP
CpVib8RMFoMiXCK6DDVHycADnnelyO2JeUguFXIVlEFdJex9TgI+G26qjtht7Ppi
qqbbqntRADTJkAdUS6GcDDKpZRU3l/xK+ng9BmofuZjfHNu3tY2h6kSwPfBCnD7e
w8MaSaHnRkDJL+yAmam3Su23lPGmCd9IgDJa5e7q4Uayy6970yBFwnH7q0GLuJfC
BbWzoGGWuGViz1SiE6ndC5fCsNy/Gbn5exJXoYs2cixZb5bbdKq5Zlhgm1EFBqdb
Mw8pVH0U5+eBmgkXsvdHoS9MhQFbTSp4rYcqKXW2ZXEz66EvivIO/JxRf0/UePgw
DTsdCaqVl51EkJTmgvjqR4uviKvwWANDH4ayWrxwCvXkGQpo5wMBymzboW+iWsaT
prnaat+fCYNOkDo37NNFQIf+N+Bjyo+VzNSkUtkj430h3Sq176wzQ43ry60PIX+7
Favb/6FwK4rtvuSjqvyfE8hCj4vJ+cahDaP9o1W8qBsePNf0tVabeyOAT4eBRYXh
yJq+gjANS67c4E40L1gQfx+Im4X32n0OkJFqJgo2wu2/DnQqduN9KVX24MSqWIie
iLA/sBgD8D+PagBw+FRDBjToziQTgg1Fawlxqt2KSvSGXSYAFah7K5Tb1xDNSKnz
Qhxv+bQ3kaDkkEIzuP6GcfViHxvosLNZGwmhymOZjYecRcPu3hhrapS2wdXU1340
1VbUjsoVBUgiGrVUXdfmyWKZ7w3RqqmNr5LdwYZobmAEZhN3uUdtIknRiB2NWcSH
0ouOUGLpyi0CKHYrhAGOwJDz7u4zO2rsqQTIAn4IAhNcHwO/k4pIa0fe5pgky8on
Pn8UTCD3TnDr0HeODKFQQhZxvd+AiNb3CRzPh8JFQuLVAHEaHuBNb6pljzeUX9hV
mcYK+XmhL8sPouLCqbP7+XTsC/UDga8c6TxaRNbWInIsoQjO02QGYQ0nmCYYpI0p
hmCHHbmz+LrTcH0/8ErgoB+WMdmWBjVeao2guEK4TDTkXO0NVHAAolryerfbA2vk
5I6ROZR2PBX6G7STCz+HD6Ou2OrLGV9DP9u52BFbzObTkD/Fkq023DNcbXwyLfL5
EbbEVrUYGxR2xiU+aqQd7/keGjunKqpfjWgu0nCtNSQzDIZBE1j5T4n8QYHmjClI
btifEeFtnNl11tTk9jCJA0Byj5ZDpx2rxtu8OkXOjxrSmBBwufemo6LYfTdUih6a
e/4qqPJ59Ixl2Cz4v4cxgdUXr3wyhAtNR6OeTRfiMIyRlwBn9BozdANOKm5op8HE
EJmO1A48mgcBq7RG5EDNtxnChB5rQcH/tYPozyVbyg623q+MF5eC4bcezq0Ou8u8
6CHBVuNdq1PhdJKwzCzYUSCbEDpdeqjzwQkljqSuUOyN9TQNKgcZGuHdIqh1A0ZC
0q81WuAadblJw2RaOtzB6OChDdTPHPpB46/2bskx+GVRNTWSPc48G/nkOkCCasXV
5iqqcX/oSxSSYSWToTfv+3olSOvXvXNpDZxJfSEjWXeSXceOie7Sf4Xg+dy51fDd
+fQjwwioR1xOV2xMlBZExYUCoz1XRjtjKG8yZsS3gZnA/NGs/G+v8ipo/PKHZsYE
fkl5dk7ehyToHNOYgBJtvxHscqVyPFJDjQjdYHM34zA=
`pragma protect end_protected
