// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:48 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
fxKdjdrRbcVtHBX/bdJ3Wik+fLmXS627xqaBML3dD3UGXjSBuIT3zbpG/JMLSrD6
n07FFK1MAduLznqNDVNQ60tX+uKXsaJzHi958RC89/sS1r81XRnWcJasXOtgQPbq
EHYpLx+NJDl2EhzCeiTLMBvn667fIKzd91Q/XB2Zy/c=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 22896)
yotP+rhF0zED/E9lT1i/1wQuGq56kzaTPVNR+PfboWKtvbsTpG0EFcX82FLkm5tw
KQEUKtv5uoFcdsqPTaX+DZeFy3jA6avLqeN27Q4MKd65QTip955NYLdtuzr5MFyz
u9aDmo8rScGQypS75NEeT73KuVqkI1Mc3J0BNh4ufUXj+n6cxxvE2NSkWkfd9RRv
f59pKWSmkmQTLEnN8XbgV+hg754iX7IleUPNIQtJwEiGUujDJyIXGhlHVcKh3e85
7Na3m7Q4Iix0dNb83/lIrWOsx6HPxxKqruyD2VNryztRmPQiKHmPSA300znzAyYr
oQM0nXfmXltV29kO5MmafI14oMeP4c1Ku+bWoXqAyRz/jjK3fZ8wuepQqMHmBVKP
BWFCj9tolhiR8boX9yXDeAYlhT3goRTHqUL6njOiPuQu9FL2nmFDi1vc58zXH53x
RqUVoRCO65ihspbIbMTR/1VTr6ynizTLWfmacKBor4nTDJbvoE7Hw3tpXxIY5UI4
vUrXyC7NUD/qU9cZfW9FmIsJojpTio46tKOQjPnkt4tnW6+mhtuJA3kq4qyT3dgZ
JSz6z9JE23HHw91F68+df6DIOsQDsc1LDP7p1iCrt/BIW3FpfbKAi++paVoOtMsp
BUooc5Xwck6W/AYarZbCDJphfetBZBCqEyLzVPVravSu+ydWzmoJ/kW2um87tdqy
nKNHD8oIaYutmOtMORUHyDAZm4AYWKVq3IWmy4k9LVpekteeulLZFd2ESjMbLay3
4z7ya7VL/Yyg8fbBUx3a5BSeFLWj35y8tI2jRSMHqxRJtfdPOOEP1xZUJeeHduey
Zm3OHZCPnq8JZs6WZq159CaIaNZIJISGxYL9eVA2XncJ/uCAaVeG6tJUTkGc4hEM
N06WSwFUBlF3+Cjy8PGDg/c7bKftDSTU5bA0zV+COnZPxmj6TJVuYD4t9IRkHL+o
LAVuTuBeFRlRrxEfalBwA++JX6c+EXPgqrCPzW/OMH0o9Ze43fkU58edV9TjNgpb
eDnQR/dOLpldDfmc8CLEpMCkrHQL6Dq8yh5N2Z8dcw4NO+mAJkFvcvjnObQNO+We
biUjUQXTjoMJPkzhpNULt1MKU/8NwRg/Ltmo/eY6mAbxEkYTz88zdAU9AJlar/PR
/ebdkaWAqT0PsBpP0zcESeLGV5kQL2TR8U3bhwIKJn74+ZN7S28Emt/QPn/unyrT
60YydObZCZBjmfibgiUKWsn71GS49l9f8I3UYS/1JR0GgIRa7ol5cRQyySSvKHDb
qsh71YLwj5buf1aJrNqyZAqxSh7fsckX2D3f5u1stWcXHLh97EjQHeRlUxWSSOBQ
WoRdxlQdCxHjqDayXLMhRWqTVwm56mp4eX2ZczEw4YpCO/iUDRJbGOtXD45vluHM
q5BhfTqiChwDSMCebdzF/VeOV0MIfKeBBhexzw/ajYBbGszLdHQi8jcAxcZCw6sU
U5XAf53pHwg2q7iUw4g3cCuwEeBH6qCkYB6in6E26w1Rw/lo2hlxZ5LG06ZGl39X
AyjVXbnlBGhznqYPibs/L43Mb8n5W7EWOVR7K/GYz32HBtYGUfgakGySI/sRN5RV
SSgqkKSbo4HSQENTzR8bsG3nCvAK4MZ2f6+Ebbefd4zEVxoTHpl9eiW/P1f3exyz
AC3gLq+/iU9lRxq2n5X2jf0J5XsYy5vaOBONb9ziIiUD8XG/UpbuPGn9z1fvJ1Un
K3enUmUgX1NmKWoy3/siJIImGhTlwpYcvS4Z+LsnL7FmsuIvE0sfStMnh/+lBgb4
gwpHD7y3WLgdzLoJLrWhRWGfeVfpKZWHkMBZQfP9xl/uFsNuoKnCXW7ee6aoFyE3
PVwLa+30b4yTBlO4bD62fUTZccG0oPpRudEb2uGQtUGJESSTBiO5gkchGrwSEMXj
pUVQ68jobc1Uo2tf2gKQlO7zpp50BqOHlTbRC8jFGb5PixJor9Z0IhnYQrxEKRYO
K3g+oWQMMPKzhVo4oaGJd6+/fTOUpGnRYGM+3n5rbAJOzJtsjmLlkgzrJ2nVIYAe
AEk/TpvQxjUVAIKlS0n68eNmmq6FRadpodCKSpmhQCStuS3YKinf/Ml358xASTLM
gFeAy//jBkoAGM2Ymyk+LciOqaoSSR7v2ud+/IXuNCe53xIkoMjeXFOGkCwbtewV
XhDflTFuovpF/1YGzpiCJi2SfDPg827z3GS0Qm8dhqi8UPVcDe7qyRivprVw0eL7
vFdyu6JcUUB5NWSV2Fl87H9r7L7z12oVJ4bxmop/sAp4A6jsU8tUJoa/UrHJ2CdR
eDpta982HRnbk6oMxvmD4DjsrtmFweS3SHw2R/F6GHQ9NLX1dk4Xdmf6oTqTflWV
JH0sv6ZgFUHC9Ph3RUkgKvzF2e+p7v1Fj3tjnPt6BKnHwDRL9sdpMP1Cbo0315wK
+aDSOGidAIGSLdVjJ/9RMW4T2gP0DC6uyPuyD/AjGYo7nx/XNec7/V2iPjnfek4n
tHZyrwbeYbNTAb2YJjVRhtNjmotWA26GgHNNdU+PW6n5UG2u5gbcuUM1rG7MduuA
eExzDMfw4rYh0IIxoTGsbL3UkM0eQjpZMB9IxdgX4t6xKxtuDebsmlKFhrCeVJnM
KPm+QptkvRe3X+NuszwZef6Jb4HX1WKBJJc/978Xy984CdGWDcMT5vQdVzzwi6Oa
O/Xke0kBV5umvnpO1YogLbSuCOlkwDYqcchlyWti3kbLNmklpSa582lYJ8uTwwqy
P36q5dlLgDtNZBwASqW+uVRdtJb9TMdQllDBTmQ/iDxjxzUf+vf0dqai8VRNpmeo
kpIExTVwzm27wXiFf4RtvY1/bqbTbWfAIKBCUgxnLeXo/3HMkUpt+REt3cUi6R0V
fG+I2nWyOr3bEQaxj/v93Mc7399UiQ4kd9xiqzn+YExwwplooTeHn+0403M5qBRH
EkFU1/+2ZVnfKWVdDShtniMlUtgbxeVmCmbz8vFdC0yHG9EVlIKalHcZ6dD7xbxj
iaNkJW35NIyKpWplmUyYj3ZmYMlPM78U4FhgTd0DJcICmqgsYdzhoFxaQRmuyA7K
cMaGXp8dQGQRqQfT/o1HmsgKuiVzfHzJOwIALWmAhWHKm3BFLzAxvME0sn+Qik16
Pr3dSh3XXsWeMNRPi2ogY6CJoWjMjS8AVN2trkQK4fNUXP4HTgAuwic04Q1lHE2w
PBTMuhGOj1hsPiJ6ErqQF1k9aHfbpyyeVC3heTcC9UngyqdMkskmKC9ljXtE4f0N
McFca2nstMXrlazBhthc+GTa6IlrKyH/7Pi+2N2ZUEvNuQ55VLrWLA4XC7r0bWZ8
XPBEq75uKRfg3ErPtsc3a4PmOx64vXbDR2ZLsSNwIwLjkPvuqMqMHjGYOULxeSCB
b9hCjojmCAYVOiRISf0JNXb/3lVIMe2q9NL9SLC8rI42k3x0aUPFKvLgiecVBhoj
FpabwMuA3mODxzlSVrqLy57uxpjAGhf/TIr3DzD7Uq/UWTJbjYKFByAefgUYNwpq
l0zkC6XntmRQtq1+mnccIZQ3o9HtW4/VUd77TDBS39xd6+4snEczTqdXkNI/8eWf
UkzYKKaO7jefANpM5qX0iBNy7yf71LrlEH00krKkoPSJSqvJf6hVK3dxlxuBowAC
1QsyyOpIwq2Y0ZlwozSI183hkd7B6VDgiCa5PGx6urkFqYtAcawDjCz/2j9CrINf
3VwRtmu0fbj3CjlU6mpzSO+GBAsBzF1Yzo4FDG4OkhCieLQOG+6SVoyqMfxIAvJF
jPiwwS31pSDaDYc5bWesQ1IlqkBHPZoEr9ZmUe6ASg+EyoS9LlyGFb2CKr1fQyc+
m7634aEbPC4THt+bMsimIML16KmpyK2vwFEJYlidwfRl0oM9xg3rmm/m5aW91ium
xVPk5LnOVjncYjb1s35MFG1ipa55guOvCioz2u3hz7PLynnuLi9wW5IGon0sOGUd
NDeNUyew4vpE61OU4r8HxayvtU5OS41KeSjDlpuLkmf3NQWvjGh7NFI3RlVmuXsr
1v4DmodqdQON2IIE5NsJ6aBZKNy7SB6vA9pTlvzMa3eYlehN/20pBgzQ2fbd3QjX
0fW8ED3+sptRFGkQhutjJueHYRBi8vyrzDxmlO9SH5zKIpS6Dr6sETeYI/rzCtSJ
u08okI4ZOSetBwBLUmlmJ64aXU/U5T+Lnn/1kvIsLK+k8bS4IgiThkIPpVYYPTNK
ybw3dV8ZPeEetdKRwZ/SakMttfMZXF0II82WPaf91u8cPJeuzJ25IQClh8LrMQEy
tyMsD2gTCpZTa27XGAH90T6wI17YvlQNaC5yrRsqFQhGFBdWky637fhSQC+GG7/z
Fn7RI45L2uNFKPnH5jlSDpLrDRE66cbnLm19jS0tchBmX0QKf5ezjJid9bnPggXM
egdFmNFJOtH8pMs6yD2zjvKZWTBEheHSRHfXbfdbI/LQ+yQ0KynaBJw76FEGNEiU
kNR+CqRifXXG7A2OeE86m6R8ucMRJCvnFxCVpFG/miOTVCf4tENgjiS60Opd7kGv
o52kM4fBd4JVgMlCsgqf2YmqknKSRdMZpbbZVOqSdYSaxxHZnYR8KXGyq050zx1P
tDuRiZBRc/XrBUzeU9++s57t+fCz77u0n/EnsLADjlZdhpcJTsLN4uw1Hh4t0iH5
tDtoomU92iYTj+igEHTGL8ifyQ9IJNdvBqoP1GPcEvDht3wwyYKk9Bvb3lkwABAq
mDkyIAK5hP19fOW0AcgdPXaZC5J3p9ZCHvWsrmykAfCTlODQ0Zye5E4fWUJwJZf+
HN73/BndqAq/J9LxK/M/Rvd7+rLneBLSnU7+9TTsKIc4ViF3laWx2fPQCLmMrQ7Q
S5duOGZcCdOEkR2PH8hH+QXtx6NbkeH/i6olgHQC2MwXc8d3Z8Tuwez9Pzxp6F+L
wquolX9p6VxN8e6rNWFiiNkyYwzUIxa3mOJD6Dk2pSGHxWgyDO2A1KnxZXs2jECx
BQx4siHo4+Zlt8+UmYCBEQY9QjAPQ1TXEoaUKr2+PBfvM7zXOgIxSfmV+rlwODbs
jTdVyLccKtv8xrWo/1qQRvWHwFystvnJO+juoqX6/aIYwJsHEVHygFerJi934fDy
TF/cxoVHDhToUwMS7Ot4dArDcsOnE4eB4HZpxud1Pyw5XGWd/fBE1XyRnYBS8j6u
da4uy6b26zE0QAvBSLnjruFIro/TMXe+mOjilG/BLWmrilXaXF694ZxRyRmIUIxI
b4KmHDpa2/mSrKjF1/mt1cR9WsMjxMZclr+lJCOOzjaBAMTshOMPKjkEP6BPE8qc
0wwmhBCECsb7iF26SZhIHG9aSyKXq/Oc5fMH6pFLjakedS1xvBLvzLFOgIGopprS
+C9X6QcISHQwkmLht/7wVB7XfsCGZqfCQ7pYFEHFI6MmEXRfDyE4//jZU1D710oN
Ep5+c2kQIufRF332KXEn1LUzs+vUbfkL845oXsemRF2N+wAKBN75yXoXx/BBTq3/
zKbSXFsp7LawIxp8VQ/aGISMJGzvupW0XWxWaO04jL1wR1REg+QwWxzWz3XvGOy1
bGtExGgxJhwXIE4fxvD0hMbpxXKN3Qyb9HM53HJDeJPVXIt44JMnUwQtAE135ObE
RIxV68HXMhLDV2Bto7Yjgg2i58I7tGwaWL0aO1paFYdSq9R7nXC68jGJTB9tm7AZ
7l8N/cYEU5uNgfER3kDIiAOibl40khVb6mZMTPs5s0DVWcTTJFLgv1Q5o8VHRPLi
yHXtOUD45azItYCqFZagqT6G5Q4rNei0gcg+OPXlQNrKSYFcHgoTBxNVnFmIZRl3
ZO559fO5F8ujkDVB4q9lRarHK6/jlZy1KR6vlUpIIBGp4hxFq4sAuHjFQ44x9u84
m8bsd+HUnFYGz/OM+1/9s3qeMRQ2GsdkfZXaqOJedmX7Ox16MwovZ5lz33IGcHLu
FkumSLwsr8e8M4GRzThydhC7wVxCtFb/to3vnoMynorsdIpkBNFVcQuh108lSV1L
0DXj8LCT5rMhJXEmr6pM0X9w/XZaEHy83DGGxPdEfT4cL7FNlc54RNmMpH16McGs
kTP28qo/tWa4AKsY9PhlfDkpuh4TYVUnVkSUw/BbBCiqzvsbORm4pL8ulEZWGsCE
W9lrqOUg0SQAf8mRNR+GtFcPWpKtrKmsn/iIH7kP3mMBzmMSYVt5fr4QCmpwGtMp
QBi60BKlqCraXdaKx4QGp7KzhqFqYFm3rsFsFXq8+R7w/GklpxX1KGLx6iqtQ6qe
pKYl9NWMW3uwbqAa4OJq9gDAUpEdcDYqSLE+RG3NDVg4amtNtUBxgRmrUKe9lWK6
kHuocBpM+OgHk2e5/wC3dvV3zkiQv10KHBqTCASVyQyNx5qj2e5LWetKwDol1HcF
nRJhKViLrsFOZxnfbLuoXZW8dVFLo0RZpLk3K+3P21dT/BuxfpIgQRN2nL5jUc+x
6b7c29MhyVIB7SnUMp/aPuMwxo8T/WLzwWCElr6VmYQZC7nirzdWoyFgSfEcjvmk
/ZhFW0YeWU/CCLKwm1nhFONTMUfAkyyQ213U1M0PzcDdTWQ5TMukfhLQTQEuwTb0
p1azv9lPpLWrTIbRUAqtZCH9TqzTXx53GPI+H75sU5v52Tbvg0lbZQft44oV50fX
OvLSqC/V+SQIbl8xAsByL3fI1fsvbY/YTtinNTW0JPx4hP3HdqPhwXeRwcD2U3P0
X13+54MYWDZAa1Vq/8+gKLuH2mNIrcjJz3QoNpfqwAFVfJol/zqtKD3hfxZl5QGH
tP3W92Njt7S//MKQT6roso7jJa/KyX8OLRcWvZSnwprqDj/8jOA6I30rXvJYz/pg
cqg2zmwq/X/fC4yLy/HQ1p+MwPkSm68W8YievRcpnQJl2rRCwFzbqJokkwrW1ywd
b046bMX18sNq6hMTEWzBXAKTo0XEB2Hd8t32DvNRx4PxtVKelBdPKuomXCNsGlfi
bnIS6QdFc6x/iZ/08MLymm4PJoRP2UFk1SuH/4x3J+dF+xmhtG9ZXmo+CF0G/egV
L5Mk0ya0zDWFUm9M8hXIfOV90FA28gyCVA4QW5Mj+1X4xAM+/T8jrHJ+91gkqK1m
G+jhgx/X407h5xEQ5FgDD1NlsU4/+LV/t0l6gS+GATBTYxaEGMCjC+9s38L+uoJ4
+IeoooXwfNHckblWUz28zF5wkHHngD8Z8+mkm6DJ2c8/QaFO+8l6OelLMkzbhrQm
lFLO3k3BEYyaM0RZ1eRfxaewrlovDjuqgINJaVcBAkjuszN+e0KDaGlujU7otAoO
i/eo1/127Nsg9T/d6F8nVpNcOkBBLocwkWD6nurwg2geNXf/QFSedFKpDGLmQ255
FyEZ23LHib4l8ktYbEHNWYzP6lGQ8TyuwBlT24CPP6h6Aol6a3IntX3WGcD5Lb4+
R7IE50fWo5CPzliYSHtZptElEx02cpxK52NWhDGX/muTtTpr0a7IvWegQqOdS8sQ
BuyFy9hCCY6gw0RdatCLhX7SwW2s9WN90qA0S2RM5SLSv0VfENLkeYQd4jPqE+Dg
rzxM4gLEBBzU99BsB1aM2YrWAB0UexTQxgAa4VKDnhWscGoLtWCbLjAlnge5DcOM
UdskLakvk0fPop7iany8lK0PRvVerkWhxRfLQ57/Fn7+NjswWls1ZcNyeKjN3LfB
evb7cRQu88VdW5IRQW+TZqawOcC5K+AYHRoksW+jaNGDpqhwnfpIqpqaNn6Yn7lG
zCKqUPZz8bbXDcIM5oE3Y6aZaV0yx3UjFEyukCGcTq5t/go1FubUvGT+phXW1mtT
5CIQzo49bwgzkqLKEseTc3JJuIuL98DjB6Y3lyKw/UEEGxhOenf4agxR476ehSfN
Q4db38m1HBiOs4ipA+kT/b3R+mGU+yB96GfWS0lpnF8NAqbx+Gu3Ev/TOrTjaqzL
ASWJY2vBE+AsNFheSH/n2u7sPfNGNKH0YZE7Xh2txf7xq2kLBu2o0K3p8D1VdUVZ
mqIYogm+VkNWG9IcrY0epWc6JIjUXi7b586weHP+xZJv5hurG4TKczY6V0TbEfEj
LL7rhdPSs/DxdyE5MjEhca3HF74o3T2/HXNO9rHi+VaWid6zQAXyA9TQNQh7CSME
BahPip6MvRwJE3myzoyoHOO4FlXjxL9cRasbmtlJM4XTWmkXllNWa9yNfGbvsw/y
Dg59MMgXySBuwhCYnuTq9Ut3fCu0Rtcp9icckHkSVwiGGDjDs0jpm7gypmQ6SkwN
fE451chDPrjQ4usvL1at1B/h9itsVL+3NSBTczVtOeD09pUv6Kkt0ycag++bw3RW
Ehd0yZKMqx9rlKAUMeYTGCA1INqHAwSn6MGBldZOkOPpw6ua0iyO9OoYyFSkAfcQ
8CNM/iYmp2e0X+XC2vLiy1wwCrWqHh9QDz8v68nY+wJTwcJArEyOLbO4tVmAD+NJ
jAQkibIZaut10a/rF/q2rOd6hRSWqv9l8StG915PpwV1o9yaHUOpxLBvUt6qZB11
yEFNHyHmjt7BN0KQiMSzmD7F8bRsiBw1BAgjKUVx62PBCAaWdfHYsg3YfkeOouk1
kWTJbc/Rq9dw/PgeUhUlV+Xdri/CzQD7BUVqUVwzPFkDLlHp+E2Dzo0fp4pLFQPh
kgwz5mNGUvT7wiqXdjvg2Gor3A4u35C5s8fgDpBnN9kH1TTGJs30rfQV7ni9Xyqi
IONyUxzuSR+yrLM7OxWelnKS3BhfNfI6ofR+zMVGTyXYAgybhs20QZ+ppcffdsmG
lrbo+ECXHkcu0eHMD3sdDpvvY63bvUnKPea2m1IwVYwV2xKiL4dUNn/4V6Q4w4Ft
GxgGBeect7rpT7cUZVn92LB9Gc3r15nhl3+K4Z+I4l4oZTHFqbdmF19vmiEJ4QqU
6hKspPLS99+S9nx5RG2N5tNEPKMEvT6DPRJpXf8Q3U/CRLskrco+dTBQbjmgD44R
PyQiN9L2nB5bGHz9HPg+uUseEvmyl+VXQwyOjqjvkmvAyOuHTikVkRFR6W3TXLeo
Uja6GVyOYhCJbSShXxjQVOhhuQhTdziPzUxuJNUH3kG5zzlnPjdFbiAwBmWAshIS
sloQ5tcd/vKmKl7nwdEUeLk+hL47hWypDoIxIale5ap6oF5k+UXaSZ+DZ+SotuYX
jZBkDv4qjuDW3sMmt4lQwNP/yf1IjuOixsfnUq80nh6ERYFkHJOif/f0SVfaeBFU
jxOONzphccHJ/XTBhjrJJ4YHa9mW4xIqKalGw+38Z80qSbxgVSU8cj2ARgL6S9hK
P52fll83Rbu46M+PqNuRG1gVQ0SIYHvio4adFMrD+YHvXErLPoxmo4vF66imNcLl
TNh4op88fJEgCg5z+Ts/eVOzBkcNnSkwol1E43PBTKXQnA9Rm7M0ykkP7DTprRm1
0EdHybQCs/VWbG0XGzqk6vXBK7561RLY8Fmf12r42Mk4yBbla31L+6NhXCBElDtN
M9fTc87XB6RQKlG9vN8iDQbJCyp7pGOJaganrweK4xZy5avQuL48bVvwD3tKYMlA
7VBQuol8eSdT3dMPBfToIsBkOV8IC+wnJykQMpbOPJwDfzgIOqHYD7j6GXZWbF7e
gT7eHI4RChoKetuUja7Af5lrwM9xbbpdBp/zeqJqp4O3YYIapnjWmE8DvzH3v8Tb
WObxM6pfsDeXmfPYNxMCbPEOzykrWO0IrsytRInLKsp3/IYXlHDIzmXBOttCeQWI
7sv0S30q784pV/iBUJXef94TLu08MN5CDa7DOOFb2Xs9dulWm2GpCcb5FFCH2fTM
QjratVOUK+cu5lwos8b6YuFNquO5XUssqv+EW+7pp5RUW8gNmsl3EUEhZZfGENy4
2gndtyDvjcuciBorM7ac17iwo571L+UkNI0HQmEt4vypmg5L6tXLFVSz38ONX1xF
KI3owlryrM5dUZfeleAvEMwYbskVJk40qi26qJe40YT5wdh8In2xxzhWnwn5xxo2
JgZpZ+Zm2uPP2jAuGbdlqKF9Ddk1w2Efke6m62lu8tXUljO6xX8h4sYFIXjqxIYI
JadKcpc8cEzirvwwXJzDxrd5ns6VHBUeMbdM7sRy80ZifOlc4X5Uf37zgkGJFTaD
Xf27GOiLWrKdXy46tIAOaAulutqZdFQljFDM5YM7flQKuOUAcwTlESqH1OIYxVY6
kn1WhF/duNRO51LaC9lKkDav+xqM9Xj/sWMr/TYNFevCjaojMAe0lSsw2gxOOAUp
lXlbPnNf9Ohj2lxZUJSSZ4ww5ctUeHgFa5iULWfAQWqt8U0m3QnYvjkGlYL1GA4r
4SMrALXBdnyr7hby9tFKer2CUWgvOxg2KRp3oB/vAey0DhWp2Uvnxj1bhqQlncIr
mHH7+RjnpQZrx5JtK4McLi45IIIxpmYK+nQZUziFZNrVyEp8ULstOBz+xhnFTJgs
XtfPQT3WcMDl79606pQ8f5DhrAn8rBlnpwhk+PHN+xG4pL0qLWDKw0iXTsa4gXHJ
oNhNKu3vcB5I2ekBY7H6koo3I/ij4qyemV5lyF6qMgQSOAce26NcYURmA4ugt71k
XWdAsQjUipT2YCz/yUmXvCX95AkgVb8p9sGv4UszFPMM0hzxN2MoRD110sQrF6BD
fRUFLcr+pPe5aDo7n5pYPXkmio/xyng2Z2JwJmtZay/5XWQWHGpGdboYOAUBqAFl
OwvMRIELvqwX5BjodND9kMzckxuSk8klx2Hp0zjHaQOtyAKoMwKqeEaQxR+bZPsG
ifZ2czxaFF9W5ez3ez/EAkV1p5GaymphNMuANtCBgQqBqYKtFPbFTfpyjTIK+wr7
wvP0TPlcWoyMGaJ9jnrbbfKHb+c4T2HhDxdgutKIR6WmLHxUFlcU60Ux92fE0Q6x
GEJG0m9xzg/juBOj9RI23o7RQjvlIl79Dk1U1ximMVTc7Ow7QZbVm8ePu+Wq/xRY
vIIXk1Y84zznh2Qd727Nu/v4zY5EI6d2JwFnWYQMjxZ2F3FNmqSMUZGXrAYeWccr
QraPKn9KcKX+S5CQBKnVEvM4z8804Vcd6nXCgdXSSNzwRU55zXwtRLz/V8oBCK1J
MwpSBNpgU3j5fGcn0B5Ij/TVYOPj5pziQJlNJ9YPm/szXDCTyn92FCYTBTK4QeBp
PAL0ohBPBaoFNfWS7bKAD3echWvWz7d/36b7GJTtVpNIVY4zFd5fwzBgiHu0KukJ
K5ZC9PSe+SqTZTs83q5tDkzyFDPdeTMU6jyJSL4j7jBUNvsrpHBi0UnWtCbc73PU
iCgWQykcjc3yIXHzb1Jx/L9eevRkRDopaVg8WEduSJPB6W9i7G/sVXbZo7RKP2cs
uWj5y/GRgYswo9fgvT06/bzff9dtx1Rr4Xjv4btzqisTvVI4Mwr7a+9J5+J1O5Eg
YhMfATqbdm3IXT7vbOO9jl7kQd3GI4Py6DhISg98GbaCz4SjJ+yd87fYuVPcmWC8
dGpGWDbkIZMlXSYiphbef8wfCIg4o6w11Rb8BYAKtJDq3T+FUDPQjkjeXrVXORHu
aB8P5Docb2CIqIdF2iIv0c65CB3zEJUPHIK9i3TFi0AxIsIR9dfAXTGgUn6jMkDn
6bQ7AX6Vvm0D+getxEquXyJ32g6V8Dho1i8fb2+TrBx5/qZkB70zZQxmfCzJh2Kj
KFSoCQUetsk2v1Q6l4FcUclBjOfkvbtKTijHkZXE7LqyLLHMf5lfpzn7Ctk4X1Xe
SeWVhknQ0DyZlSz8cj6rGrM/YMD4/83HX0tec2Zx8uARJcogqWQ0DkkHf4+QLB/Z
v+/P4kePKnonsw3rApU+9B0XDizjahe4mGboFaOpgv2W29l9wQTrz7mUNoyCM7GR
ImAcVXfr9e+Bt68QzNy8zxkzmtQII8rpmCFrRWlHsOhv0HEzOLE56qW7BCzPkAFV
3AG+1tcfYqNRG+jRV9P4YuLj5JHM57cv4nxeMSwhuR/Cl3R6X2ro3IFbsT0TSAXd
ATnLHVLgO4y6nMBsQAXPe8UUoaSOj+eBtmUnbXgcs9/3DF6/apJYE8dIwGBRUrH7
rFtQuOgAnKjVayLQZZ+NA+DC7uoVRuIQcMX15kku0vwFeIDHncuESmzFmMjKl1l9
6bqtjLR3MrptDbPryW5eaMg+Oc152r2f0AX4PrSciqZZlqVXNHf+WsmvkpIxY5Rj
hXd9mqjiYlbeEE6rSmHESbY8MB3ZQe8ZhyJ21aAtfbvd9cXU+k0lm9MrtKE4WHe/
s5Xo+UCCBnie6uaFWysANri0WLnpbGMdHJLkMxxCF3/bmtDnN9exLi3weJ/6za0n
nroxDbWWfA2zF8bvsJxDLI8mj+f+9Z9G6hOaJdFGS0ffmOQOpaFW/ZHEHwfhZDdF
OKBMQlGv756z4x4m/rRiky1h82ovLra6AMyqW2zTr8Qhm3mYnTP3m239bHzFZpvj
9kIzrnbAo7eVQjeY6iJoSHPuFvrqEUz2UHhSKInc1pITlYTdsE3sMDscRnE6YOti
l2M3aYciBomWwHh2SB0uMlgAqRT2rFvBM9mfBbmJZz0yhSDRYPy2CurGZXKGSqJo
9NIaim66M1xirnVCm/raNdwAHF1qmMYaAXY3NKwmkt/4VQ/1h/UYlKF4T87vN+So
2kdZxMuFvSbG0h3gCBExi71QkLNRuS2krUiwPKVYUBFdfgw+Wbw3tDdtSQj3fRL8
73Df0VAsNciF2gKDojBmnpXbU4y5Wwwz/zqeCPI8JM2/w6Omz2MD3VcBYYTRWxkO
ZQWNwbeWZBvZQ/++YqIAChHKwoLpqvUdtokhTb/Ho/rsGiT0a6Vlao/4pD99b06S
i68Y3H51+p9VIalfZ3jhTeOJ/GoDnERobCxKPESLndNX7mFznTReKVLFgmKXp50l
cvxUE78bPcIHCkdPTs295R0oVDq23hwObYaZwIIyx+n31n4mECWxp41JXKWYcs5s
F7/ty0GrSAzv5IA3ryu4Ueqrf1le4EQ5wSoKmhfICh0CfaMIMSPLAXbquywRYCgn
XQQfGgp+uG44cXXuvyMgWffmPV38ZbZMv5BQQPi0rfpQWNRd8g1/uJak0ZGT3Y2l
5Y4QKXnl/ZLCeVnJ/zOparWFQWlADvoktpvrs439pxcH3N9Yl/wE44nT6znSY4AX
uz0WxtdUg9+Hvk3R9Ki8H33OdzX5zkMW6UX03lgGGy8So27HTIllWb/5xMY8YR/1
M+apuN36Jb8sWHlQ1tnwa15gvLnoDW6/bxx7RR7187t3ozlWV+us9nCBEYTFUb1+
ljiF7n+PE8NEnJQR8loAnHQKqWEfCp2AISKdviPNE1dvE71bDH42Vc8PfcHc5Dyv
k4I2iuwFL3n0P7gwttElZwVIS+vTJWLTUtwsyMs9+o+FUhO7AlA8SqdbxKSZmJdF
ObLlYg3paMRzhtYhvftuEr+XsWrik0ruD5Z7QEqqlZNlWcwK5tlONhThU95h2K0G
zJ6L3rqYG3zE/HCTXJNB+z9VS1mdD66Tv1s0/0cGKTRF7aDuhMWvXDYsdFeH2CR5
ePAVpBQWjx4vSwLmsj/4d3oh0BTEcKA1Xd1pb8UCsRMNHb8S0qi5NnlgyJauYI0H
fn7sDQ8KvD/PEtfuNbV0fwrFJZxqlx3lj9KL0enFQ1idJUN16CIj5s0Kh6Syq6gz
atuqw4keeEsFIeNS5xVDbWfV8RTrt2KcZtwD8EWtK3yVG6tHLOvs6WYQfNJteLMZ
827nTl4J9f8WGyzkjxh5l31douxPjMe8Tu78IH2EdjvEASemX+3My1E5z7a0vkxt
L0huvAxvSIb+TLqs/0wxpKwapLoSUhXFwyVYDRv+uxxtlR9TwKlaD/nqIqBIN+x1
kmYbyJfj/DVBhnz7z0gwMIDNgaag8U8VyYkk74Nq4OAFvVbHHdpDMymxUtWS05R1
zkMx85PXWl+dQ9h+ElsQpJ5uObW0JQR7KoJlf4f6gRb5hvEKFsy7E50vId35HtLq
4uHGMryU74RHpssoB2otTqP5+Bhaz27Bjg1Omyk6Atk+J0oVyxXmqRZowgRbbBud
ZMyiU1Cw/rXsWjVWtQOCbUhUDZyDVw5F1urXfsuK4SzWbdFNKDLRB9Vh53bnztCE
2xS3dagcM1CwkFMAqumj+C1deZiN76apvgkTAvq5rDGuL2F1zq6KzDHEFJnhLHIe
RhoVEVU04uYE2VXNi6NXIkZiNJ9JW/1NN+LCg4fKUf+XFHebbwh6WrqjXcNBojoG
8jkB14Cos1oIzib4nYogogY3TAPWf0bdZ/cB1ECoSoQNxrc42tId+tGCSAK+WeCG
O7Q7NGVkfpvQ4CrSbRxUrmXfSbdvQbP44BKchBR9dEmzBp/X3bleo0HOyPx3tM8G
RinYYf0AOY0twQBH7zxlXGN1gOLvZYu0itNbwbE5cHnotxGX94zZgTlP+FVWpq94
RW6dPQSM79H7zL2hqlsAVUGy/tMMOP0fkifdajPJvwLG5c5CZF2BnMuWMgD+6GRN
6eYLaGhGTnFi3/wqQPYCXklNRZ7DTGecLdkkHJHbLuZzJidlwEtEli5C7ap4ZmIh
qVO3OhUDn8p8BC21xIMs0dUsJcQGE6b/HV4k7bwqCqcYaVAnHI/gW4Vfxp6epWaP
Uue0CYC4YPyBjpmdVR+Az7fNhyquwjlaXi1NMGtriHXb0JmUDITxHhLSMGFZZoZh
v67HrNVwlHnAzw3kPYg4/13BzCzYWwp8kPhQJJMIbXvzng//Qje8WYtRJT3Xski0
2VNpVihD/9s85yPzP02nC3+spmqMLlO1oOoUrVl8Vrt8qFgo6osVakZvt2hC21iH
uLC2SaB4jnLmFQrZxlcu3VESBfemI1DhhJFuLQHFFCf1tMDrq6DRCUOHGRLZi/U9
01ZLb2FCLvB6uKJUcI42cmaEIMPFDYSGr5t0ySUWDTAXEBc1yNNS1ZL1s1w7WtB0
pEUqi37fZ18qi+PAhkmwCYnOqFdVG5YYw4YoR16h4lwEWP55OlNIAYesdFG8Zdei
2MZ0D5ks5VvnSZG3WDYEMvdY36ncxXGR9DNo6XSsqS59oX58C0hIJHhqvuvxwdUq
8dl4vTgr1wZ/JxdRSzwTxyr5kQzGBaKT3zWQqyud7ccZ7GE+dHEI9KcNmiwwhtla
B6EUP89obNonlDTLDQo67H0cB8xc3EBZ8fP0Dzv9gt16yEGdSXIGO4H2ZiTOQmZq
mR11DMLCxPnMeBzyqQOYUtzNQxBOjXuqUa9YYh7UtLGx+ykRBt+3U9vlz9MiJbKM
9X3Vw6k5WnkZUrD7ufjvCKSbmITadvGxuhybJ7m2EM63A+tQrAJXb50VbeUSczld
G82QFlMWFdAJhpXMkD01qJpu8emXIGSSHmkBZsaaQyki0w1BYXsXEGZGR5tmlY8V
qXV+FnmQ6FViDs8sew/xcqLA6zpL9Sc0tS+uXIdN1P9mSQzzDN1XrWxaIlKavZly
j8Yd50jF48++rRljeacmh7zroGTbYCSQz7ffggcvAzlZNZ6SZXtI547fdsYtvwFk
bjeDlMtvmHwqye6T6jnBwaIHqVgEYSVS5WmItrGa/Qdit1qIDDPaDg+gYztBbn9l
VXRAANuaLkVuAIDqI+d3OEmCW3oJjsyWL76RNFu73GFVMqvoPyvfi2gZuhTYC/8R
IvKmi/iScu2cwlNg6rDpKobWcfXsksWOEu0g6tjr6UZPUJ6TPN8VgOjOGMPQJUqN
Lq2aieLU5vp2TbQdGPBPgzeco+nN19Xlygg1j/rJ40NSsn1L8zatlc482WBFe+03
LGQyJ1beLvVzfyafk4QLXGdMyS4wdP8vaKBGF/7zG4Bg3vwbbEhSnaUaK1TaUi3E
9jbECaSlVyE5yjhUWkW85pDBmvHDqpYc36c/ExdTYhu9kQ1XdjacN4Y2NguRJqh8
stFOuaLvaoVxXpLCfnccOYuIsRt0xjgYXPyLYyb+GlK7bh047jv5055oUJClwOTo
2goUKaq3CJNjsVEWvSOQ2B8/zIz6VV5EemTIF7Be2OjPwhkY+LuOo0xspxl/E+1j
JKYeQTvF6EX5uXTxTDhh1FtSmk0JJM4jTGhFPoqlcs/0i8ASWMhv95CGbZ+2nAwp
sozSOOTxjkwyu4WF/J6uW4k2HhzFV6Q/EwtFU9wwo4YoVApAFBZDXOFY39pMsmM8
ZD+lSeOYb9IexuwxTZ2Va31s8mdT3pIeDLUlRSgsM4dvmRbcouYfJvdAx/vGXZ1D
X1bM1nCHbrLFlLQKgFvOkNUfzX42VkrxZJGifElrLBimHlsI5qipFoV1doZlogMJ
zg/A3go9oBsL8OuVeMXc5fk8EfcaS7ttN85USP3+6AzGn6+2C9bpan7oV1KpY6Bc
C3Q5B4jmA/unbfASZTqJpR3ort+hGWvmPf4z8L985hlebaTVE2fXewmvE9WZJypb
Rys7fXD8T8sZF2NlEvonW+q07CX9i1hMf1RnRqmEb60TAxWRFFs47DzUr+jjxHzh
jeZd/H4pT714zWdr+Vxv+AKGck1npwH+Nqqvnoqt8diHUa0JQ6O2z/FONcNGmlPS
juy/dtZu/mYbt+kN/x6WcBJRMZHRqJBcLh5TrENTDXNriTDViFJKqx2Gx8M+2s4U
J378UsUeVpPs/RtFORyapFXrp7KglI0OYEkfiOz+MangSTLYM2oNntIa5kXhBZLH
SN2zXT6AXxmMqbohJNDZrHyY93VQNYHUmPFdlC0pNEYpWJThroF0jFqKlzi7a7s2
zYNlEj7dgD7oFI6xstV5aJtIXCJ3fUfqpcc+Qk1XCWZjJ5zG/2tiYL8nrCkM8YoY
yelmKyVsnBMkCOjG31EBPmBWD5Hm4KKKdgnd4ubUATMXZnNkOwSELRHWR0MdssP7
ljXjHv/B/C57jLoL7sFpztZmKiiOd0ePNqDyk5QM2OJMoGItzdrM6o+Aar1u10EX
B9NkCSrFyFmCbVfyxWDGj+aD+mJFhMWP87MJ/kZ9OaQJeJUpSzoYSqWzva2OQlUR
2Pa1vyBvGAxZbqJqhXGQS3wrRo7ReI83dLSdCKYOl54t5Z2O7r96EFWtQt5IGMf3
KY7y2enJ6sRaiI5sV5ZYiDF06i6fbDcD83U4pmB0DK4bhw/fQAs1DLbvhIPmHvah
BcvQG2GBIUf8dPO1woXJumKh9cr+FJu1/+zFRyuC9QIOOl0+xq9vU++ShVApk+Qy
6us4LBMesP53C71uVWgYvjAoZIkG3t4RIacOxYlTGqj7Kcb1phd6XW7VINE1M3dM
cU/ylfY0f822dFvrNQxZKRlxk0hlh9sqFgfF0o7Oz5sXhWYSu2cgTrC4aqKtdR1q
I98kZcqCfO9xcbZKVX+k9uuQ7hRqbJXHdpsbd4s0Id2RA/QyMVkjxi8r4iONg34u
+FuUJDFCkHkQEzbUtLX2uaYA273A2KaesIqBOhtfaCJJ9EgekwmDo1TUgVEbOA6F
qLk81Sh26BySqcAH0kgSVvNMLGmCfkWBkO6lpK5wFqB3mS9k8AkIodUOVZ+OfDdz
6VKLMbs6/EPXhdHbVJJqWKFLKBn9xOdCGgcEMtqKCg5POw9inIxcfO4vSsASq3Vu
ku2CwN2tb5EorrZ93YWqseWYV6IMVPH+Hx8/qmhCDZ76UEybZ8wX2EP6wZKwB3fI
gGdzqHX6YHS1+p7NOu3OEt7UA0rYL/AaHPQLh9ahX/fPIEfzyScsWunO1m9s0EaW
dJqjscPsGUSaiQNNSPEa9Au8cl1OW8fc2jn/EdBn7Xh50Lz8hgvO6KymQyCODS40
tf8gkcAgCcUZZlP3IvESwEVYKNfJU45+08B11SYNfk29aMWHMdcfSrB3T+Z0s5Ju
HMfCrJwlqR3RPd7q/TKFLCuZigY3c4Z7R3VVOI10IBOMftMXiwulHia9cW9tdiKW
rhuMqJizNhik+FKGbqap28EbGx1KncIVAflFXkeoQ2Mg+rOqBs01Kv3Gc3Hy1yBw
JdwKJeLfSfW2fhWeGkjPI++I7cni2ZfNH+lGrSBe8nwWLJXQJAJT3255bXoJG80+
7Mh6sGIR9p+IV9g8mbVHd6DmSCAN3P7wp3yOKJAjEUHV2jFu0UrDUSGvEKSmY497
oI6s7u4hCE7VkhvlAdHFtBf/aFP2RLcbJRidEIHSMeBfS5+RYLEMDHGzXAUO3MrU
IpcrUN3YZbrWL0WwxmEIkiOYzmPWxj3bfIRO+RpV0q+b9W0/spA+nKc6d6gEfSim
V+qWCgp2ogzyOUkHnqcUV6mWKwIgLdkpAwC2XvW6BUaP6cGExCLzcciHz5Q4IDX5
9OKnIv0txvKbBmHqZ4zbKzqKpy7BKKBGlvzHBzNEdTewtw7XrrfTbD3s/LSUFNSG
p57xF2b6406AJxrky54b+TTMPRV67XIVzna6v6dTS+gKoYCvhggs04E6Zsh67ZDo
0zxh7/vOe+O1BqL6M5gKvarDM/OT4+T2q5nJ1lrNlWsFO3bs9Q5Yn5UQqv3U1cAX
mToiBTGQ2iCyriM/FR5QSdYxItXedONj838jmZKgBd3ZNjmGs40ual/QdXPCwZSL
NmKTURr2bS1pnab/CsK1ooQGnDRAsLXpz2V1etHgg0522mXlF1Lb+5h4TY3ZOgWY
sA0qFw4PHjJebVLq+sFNpTIB5wNvaiZzDjh1RCuhGFEw1XRkIcvCQSbOxDP9hl/O
E937rCGlizGp0MO2Fxcb2ZO9XTf7vLT2h2QOvttJz1KpCIIMKtEAOj+75vlHkYKp
jFxUmXU/GkyuY3DqGglglBMc3mveb0la/sjqp7h3bHFprAndhzq1e6RPg7nJBi9p
dLPA8KY3IHIH5TQSh0au4MK/d8Jhrzg8xdJ50vGCgr+PvwCch0f9L2ZgC1rsmDFe
dtvAkE/RZwd5jbuopInJ5XwcMC6IW744pG4/WB73s8U2k0lgxAFa9yQuOoV50IC4
OIpwihBZuOPonyRZoE12W3v659O4I1VpRVtzZCintSBjCEX0fRkcwXazFe1OOYDR
t6zwpEAsr/0AcDfHprriGX1YqMgmBrOmPZH2UgS4Y5puZkrrzsufqdRHTT/SucdS
NZKycPW5zHj+Ql3RaQqNHxBQBTzizYz/l0Yt11yYb6ZezIqtm8Jb+DHTRWeq0hnK
r/7Y2D9pEYhvOX388y+9EghU85zc0aZ7Hju7jCDjGfREGg9XtcdeT8JRY4SA9C3u
ZYlOpMoUEx1WttwFipfY06BoueAOgyv6+qyigaf9YHR6Bd/bUAms3I+qRaRJag3D
rN8kiTLqBZh6zAYKv3cui0DH7yuGcVwDrC5xTxYRWBixZZa02zbZHgHEjcLoGgN5
tINOGZCmx+Pt1xDd5TbBIHIneWfaiBPQnmMxz2Z8sszrdNcmSvWqIQCVkKeaHXp7
lhQTViuUXz7aMq65wGW9GumfIIpgGlxr9E4AWaP8g/khkNxkY+P0177+TC6+FHoA
B/z4vQBA55QPlFt2iCKVIPqehlfTaS292pohS5SWY6S+w+X/G12TqAMqGgV7+N7g
ujm10KYC83ACEMQQ9iszWnjVag7T4f03IdJFUQe7TfJLMl0/ElqUpAq4RqcCyFH2
GYdMBEctwYWAFX9bJG3cF/QdUHUCZnUCI3vhem8F7fJaC/Oncqgz2FBm5U/wExfJ
YUyBgs+uZFAzQd+ZgFXlWzfvc3CYK8FEBI/Xz6a3euxdfcYCpu+4cIkMU30BV3I1
N5q46NoMZSq2euvJTTM37vvlWlYyMYSRK/LlxfSq36AvbiMU4cOdzCW4iLMcpEuv
gZe5IPMmC+IQjjBydc48uE2M4UAJmtAUqDrQHp+O2GjQC+sk+4XyKr0leUShw/Lc
o1xONRjteXkKCq8Ltrnd08j8EFMtOmbsMbNEGC6CpggACLKlnmv5pDQvp9YlAcNJ
kYbdEg/cMd5wCBKGeUKI0YDZHH2g3B8W44WwXTrS4VO9mqw6ngLfN/EMLA+RAstP
qZtQpL1OKMtcR6rQrbXVI88JiwmZM0moj9bHgwlkg2ST0Ajk30KqMi4RMhs4PtzY
RRqbf94vghU4FqNBkp6NUXkjo/wthRWBvcEnl+DpQ8eXacTvySQuGrDSivws9LTu
mCiyPMjoBkEEcdM4/90e89e0Q99n86hePlgz1ij/onHt7ZjwLrZTtAR+4TZoXagy
IfaOvjcq994yUbj7Bm10kP12ExSNLBP6xFbPWEqdOshadl7qcxpiAH2UeGzXSJ2i
p4L7aL9ZotDUOL2rzS3Qlz8tU/C8Ub1qX0Dl07W3VfiAmLLdE6iW2EN2awOYo/aJ
JllEAgwnPvQj08+8JxVcWON8vJrHHchCSSg1PJLeMBPvQQEdBjaMq5FdndrTdz8T
wOjP7CeUaSpiLe7qZVq/qUadYr3PixyLsYTPz0d20LxJphfOm6WMFiyKpMZauWGl
Hiqi+WSjz3K2Ojs2LGUvsCCCBzPtVHqn3TOSWeLfJpddz9grqFlRrvAN+12GJeua
r044w5Y//0dKCUKKcHtMk6Zq7CWGMYS6IS2Y6eOR4u3F7lqBqMjP070Ts3pcFK40
EQVdcCmj8k0VqLEK2UGz+RQ9+w79st30cZd29fo1FZ7dwe6DTEJ9D+y3r96twESU
Im6Qx3WyA3d4MlCl4DE6y2XZFShglLoKMto35YQLsOXbD2nZLgwT2HBxoTBgJx/M
uylJoTuSOsXXgfcSmj2hgm+oCLd66zBK6EhCO0WfeuBIaPnphjqZXqXgkG6FzPOj
1tKUaJ7AgQCh1qr5LKR6WUIvkdhBrPWOn4Bhsi3iKoolVSqMlNIb72JcwCeS7EDJ
6uyVC4nSl2/xcme+2SxCxjlMVAglOJCI7TA43th8L/A/XQjjoS31UE4TrHC+9cUr
HMAsAIIw9yssQWX8h9gTMXzv1IC97nXlt/aFGZUL1Ari2htziibJIcEJEA16rISM
KjlrNkl8ODsgXHPFOOTZCp9t2fWE/XjF/PGP2nGW8Joy3wGXrIGZHUiVh0ga9fB9
oeszmpy7ntaDuEhfqb4tX+rMsZt80mi/H4VXt6gLtkczWn+rUMPvUIkjf3hrBG4p
YuTAf23VebS+eJy6BDo3ihJJpp0z0b/HER6V37DIvi/C87imQxVFzDbFPkj9r7uv
MagO87HXw9rpZ360USnzQK89TGxIo+BSOgmA0WEZEOejoPuX4p0Y9/CjZgKzo7mA
yfL8Pd2uLS7rNnKJMdjJbNuo0l/FZp+6CCFYataVaZu+HpS92rIOKVVhgndeYqrY
pNYVrZrNk/kFrCcHh3VpFSbOA9PnEsGa2H8Ipbrvtcepnv4GcWKzo0KV/ceQqBLa
Ou/dVGD6B/yNsiCwmkWdQ2zHm1YwPjw9IGn/HmU3EJpA8jMFkEQP+p2GiwryCArH
N9qHAJblFS0EOMxXAbRF2Yv9bePWBKrrAcc2F0Dlyx4mGP4A7eVATEpJILpajK9x
RGYBL52IVW4yJ5uujDmbQkpsckDCcMtrRM79rIwXxnjRMO3EBO9XnvdhMzaPjMI/
Fgq+X0FfI99g0MEZViwElR/U/o2zKVaaXInw//YagtzS8m7vgwhwX39zWKwgn82N
by3GCzVMI48yfp/+3aKiUfy17uB/EL8mBZNSUf6X/G9Fb+zv+zR65S98plTGhn7M
YDb7PC4SViqWBspzXyBiza96nCskJ4Pej9IxQlOB4YCpx2gEWt1OHN3ABbMUsIHh
u8VKgbhuopoAc6DWLDlhcjsapm8hbUPVSnssnjcwKIjld0aafUB91i8np5DbGYHh
GDrJqdWwPNAmwHXlB09qnDbLdQEmr6yRseeVrqVb1HrugwWNwoc50O6vK6CmNANK
CtvMe/KwZM+ljtLIZ+JXosplzowUsnuRmcapjklcea1a4o6Gn9mVIazsw2o+lP+y
JqFoU3fXszLv5t619NM4ajQQW005Bx4adcv/cZOjwWgy179RjLzTTBfc1k/oFkO7
lc4tSagdUtij9pFct1gEpfaKEQ1xHEr0mx66EWm1VxNovNeozwV5vpSW0H/4USnC
w5cAzJzRQSE1QtA0MSP7sHBpp7onGZIeY7NPCKlIBXhallniYq7TD6c/I5iIpqZa
FdGaOi0QHHn0Lkdmw9d+kOTTq3RgO+HHoY0a8xC7WzD5ejkKXhFHHBJKjpVQWqo8
YoZJCJEnLQ5yqVvHwjH9HRdJYhtvcde0jFrZPiXK+FrLRivESTZ3e9dGhGhM3wwM
KiT6Tv1Nm307gXfvUj/AWjzJk4I65SaRTTTnzGaM7+fQ6z0KTZs9ZpR/GvkmkQyB
lJj2J2CWaI+i5vdFuK3AsmrlOorEhL3pdlDH81wHSxd+zhjZOmd0mMv1u/ZJmJQB
EmmmJsvrkZJHDv18cXlGyOEF3Kn/NHFLdA0BOYKbjVglImwG9YpHcbwlK8eecy2j
bwBrXJcebiB77lfAff5FJS/VPjNZ4nKZ6n+q2ZLyU1vCsoLWH6KkjHaM8cxgLCmm
EnR9VuReEKxHTcIEFCYQ+XoilV5o5GV4O6pvvtwt1vtObl1vtD4XwZ3VYtSCPgPt
Yce483I7dSIql0BD5xVG5H8yCEaqkn0sW3/rvyQHjgYF2FIycDzODrU973IJqtdH
HmHEikNxeIJtXbmeRhcBVWojUSrNlHNLheOs/nqEEelGu8lpteh9nlXSH65KV+2v
IdGrf6GgeZxCoCWzR/Bwve+/3zK3mzeADxVItKcE0YLB5q8EUAJgGMyHfY8nSE3D
rWd9Hii9DJGgKyBaqdMWY81+2zjWGIuP5jEv/u1Irsyl8xaaHlHioingx4GKSPmQ
69avD9ygc/g4HEwuVOWig4H46enfYJHLYJ7YinzRO0ldHFf+Oc/Ni+4BkyXl1vy7
f7ihWRQIBcvlwxJokTTiqCBocQgi36tQfiU5YbFYBY7oe+9b+b9D3GwzxiSQG/tM
j7RTPYqmN3LEiEpDy2Okox9kWhG4466tAVVTea/nmMIRpI0pI5U3Albjh3MkMlQR
A9RkcxZX61d398ft3mFoNN6M6VtBxYyW1zw9+GnxEi1vi9f7bRsUkcp5gSkBrqSr
4FvR8Xpevp9N1/qeBOt07zSvOj3eoSVplYKlBh3uDnCjAnj+HWcQ71xN7arBz4gl
T9Eo3cVMOQK/JQPdIbrbOmtZXa4ElKvQP4esXjgE4h6IwLjJTlOB4PqFyWOdiE85
EhFUqEL1SUQlI0SZyH2YFnDccRkqaPVvanaNG4HMWIfp6lmxGjeL5xERwpv79grz
1RR77bB4HNDnJjFnVRgGSWojym4wPm0FnHEn/Aa0Gv85UvL0+iN5JwZxn+aITlNC
flFgS3QIN2RNlETFMLWE0dzjErYbfVXgPASvjdoOg9mX85VrwVgjNkXfb96olq+w
BECpwEvYR7jViPXpDGoAJkXH3iA6KIPaMi+9mflTjg11REvyqz/+v5VLgTyixpUL
R1AJWOpWzJxVhYTfZX/wPtOexQGEaTw2Tot+hi+QX7+PBLgbI1vHPSHkqpovCIlu
uewdzWw6CHnQH7E5O59Lhv93MK9qvQzN21GLnGVlIvWM1A8FyL9M/a0P0hh1a7wd
yRf++aREsHv7N/dpiNMTVhlMSkyLysY15XvkiSnAJUMVKb31H1B8c2R3KlINmkNG
+yLUYSedHV6vJ62OCIyedZ7e6Pu7ahyFMfFKrPXn7FibuG5qfnz2fF8XVNd5HqLt
rXhghchQFInet3iYKDRrm0bDNL0kK6ggt7jQCLcXGUQ05TSvqX/XWYjY0Qs1jGkk
ozlmoEhYg8XpML78hsEfZ60bJO3pMgrP5QrgI1TFAWF5cs+N9VLs7SCem8vLkI+9
EdPRwXHnBxEWWuJmhX9sJEdu7NIrNmdu/ZAuljvqTo9UP28Ki0rC2UzRu3k2gxYb
e22MonEbpNQ2OrEUmW5ipyGOnS9ngkDyaMJSFi1t4J9Hah8RaS7JqT3Ro+hVnpKa
Z+ZaW9tfJk5Ez38jcSaQJysKL39xvvgZUA6M+rIU2TnGi7N8AFdQaA8FOdt/DekY
6P8OOXCrlRa4lAAgzMVhOMIS5NWhqmOtouIzXWHsSJiExUF0lJGpScLxoc6xjMHN
Op1DiM68ixEdgeMVXZRgS/eEnIeOiMLB0nVlh+C+tEvMkwkvb9fwsCLVXrujBStS
9kDLDBcljxQ6actwmLtK+f55gp0XDtVWYVH57e6hLqh0FZvFSeN4YnvBHsJrFTCH
ZtMksa41JELPFPEnsMMNeweLPsZ2PBk9Vb4WJ0c0eBz6DmQ3hswcJ3ZV/lcYHFj/
5MVkRPzkJSK/kns6ORHRhR4ad73qhWX6z2oiDJmaudJvFrSgiI8dzjolCl41yONs
aMroLddvb/f28gGFTn0M/+BX/WyqXlffPpTYIRQKuE7UJiQ/6hxoxpqDW4EX5TVq
5OagY4FJMa4zG8S8NemtkjIJgJEc2SMRJehKOXZHQ8UJU44YpisPhRBRxka9Da1/
RWizl/WWDH2j9Ap+xz0MK4DkKyN8X8GUCh1DkJpAI950ezs3KlwKENitjyKvKjvJ
mOzD1y2SkuM8Ruh/VItQgKOwYE01G5RFeSy40aC9OAfaTxe5tm7dY1HPGrhPyl5P
OAvYv55hWQXgJcxDPt+Cc6CxHD9ECp4uOtrkyvnL3mm2Za7rdrPi8Tz6ZzKCVDY8
7EUJvXbbMIuq0xfWJ/3fBOWQuX7ZKTMchh05zl0RijMPwDTOmI1O+JUgCF9rqaxf
RT31rTwIAvPAjdDn39v+N3nI8ft5gkI22ZHmGu5g+QA62AVBiGHU7RDrqUIpWegE
tc3wuAlkONHpRJ6KnNk8kbphuffxEFDuFM2eva/trXyCl55O/hPGAfJ2q8k9y7lX
xaujqSBy0KT2sk5KxnxzkFTwh6hk9k518WkbJ2k0ZrhxlgXuAcx/ncEWquQZYEl0
cPVZ1FSqgKcwjpNHqzMjmJR8AjJdv6jfvyFQrtQn1CSg4DsGKbFkDz1Bw25gM8m5
dg3P/V96MSzWQJ4pioyYZHwIJ8YPvDXAB4XoxF+WXDpVrQwZ1O4VG94pxSy8v/FP
BMA52rMpbc60GPlpgUAAkVHhIKIFz8IEmY9Q83RArGX0GJnsQq3X4+lwTnTpg3WD
q/F63OcbB3wS20BvRAFk1qvS5+a+t1MKGhyuwCQe8dQ7LIXNQGnIFJCoU5pzPHuN
iGdgpwl2mD+gCEn62vJMhsr80dUQFdhkvacoWyeEx8XQKUwQY/rZRRNuzFL8CxQM
L4ZJVz0NfsJXQlEuEJadGev6O74EcCe60Czap4GpCfesHGYkj2KzpvdBEQsWm4ev
4uZw5Kq4CVtvRi9nIH2og/vn7h5sTqf5A3cHT/J0dvu1XLF8p79AhgIeMn+5SOIq
9cn95yLlVPCbDgcU8T65zhL651o1VjIzafWdxZWCz4Okx7o4qgt5qzOqtoY771RT
Ub25oMGXcsRtiUs3QhBr/vUT+JyGxXnj1FcXb3wZXLCANquT4h45T/iwIXiBKibX
RiN/0jQ9FncRuJYfCUZwutdxdwpQ5MjkXZmfqzE25rM2pc06C0dCKkQKvXv7wfSB
sxHYhAkhiabXPY17z03LLfugtu7Q2WLcaJWc8camUWtGE4TVf2Da/C/i/OEwuz11
Z/GoGU15bwX+rNvz1g2gb+AdpqqF2jLpohPzgWh7oCBFeVPgoELxE7HvvvSQg3Jq
/Gk5OlsbuI+U6x+i1mtqJHxfPZfiDAPOFe/s+t3wJEEUWxe2+6ohbsV4NOlCLIfP
WY4NhVCHoADCasHiM6mc8Ba8Judj08b8zfN2MOfwM5cR5BTH385IFNh/Z2EJ19CO
poLAVw9xNITJz6a3Q0xbelc6zG+PeLOoBfg7FBHdN3BYL7xYoBWm0WjoEdWzjz35
gF6S8D7UD+JbO25zwexWE0LhY9wBEi58+rv51O8mkpTba0GtVXBH5MOD/iGHjcqB
tjIHY9cF0Se3L2xWf86mHyaEfEmdoH0tZIgRmEEGj8w2MELUxBUi4jAn+NRtSOQh
uVZuwbgVccanQZwrPDJgOmMLma3v6Ba/RKNobA653359cRIU62T94fzA0t1NcfeQ
qbWuYRlfHhfhbHJLkbid7QjqCvGET+prJgdTmkHr8Rf0eNfyRnqOWnpulQX6C8XR
Z01OKX8BSLsQxeHuTbF3oITkGuRppIf8dd6WBiddAD1Q4Q/AKEYN/nwv5+xiw3pN
WilDQQgCzW/6AK+vy/GUewwFVR8ZGonx11p0Z6gJkMEwzRgE5lAl+Z+XlMkYNqkQ
agb+6Pdd+ng0nPZR05mVyb0Fn0l7KDjSLM2azaCsMwOX5k8sQ2ZXZB3n/utTlY4s
2kcwMiBFedUnTXIiNIAUs8eF1MXNi/NEgFWjNF71Nu3kbt9d8KBDEyPrT2kykfgM
kHXHlUTf5+AaX2EAwaYkUP1EeidYi2Ov8RKmT/Dj7vGnMYS6rC3FEZe1QKm3tgmv
vMSzyMhI7TbznzdC/jCz5YbxJJUbYdeYwKL2XpEqAJY4FTv1y/P/buDFUD7x4Pe0
tgJUvarhIxD62DI55i4hnuWLWjpa2Cr2cIknpRJ//F9v/TT3mMQQkDwVmbMulecC
vu24hxH82TqesZgP3750H6gyqjAEtRfTCdihHF28sQOGEbWSoS2goTpCdnlMVySs
X4SYVWuSK4sikdjj8Rsxrkx0QaqnLb7D3uNG8gBbWwzoHfWl1voY0fdz2mqC4EoD
C34AsLBYB/ztJ66tt4tHeQO6uz4gK8SbjH3nhLoNjMMmu2z6V8cjizcd9Hjq+owZ
7sH/Hq2nRvmEqZlu5e7OumjSR91N0gmqAtAkUVJ1XiwwrvtrxhPO9F/8KA5gmjeT
AP50Ra1IwAzbESUzMmFE0XDVvlKoJk/MMmLE6yeg+EbCiqh4bdADak1OrWrF1LMM
ZclKRghVCkUHvK5cx7MWPHMdehyICtL3bVH0BYdwpgavbWKhiecjB/rugKLP+7rw
J/zHeHMbGHrSMX5tgln7kwrPmNLkYD6PXLCep/HQMfMK9ik1oMcZ4yori0B7NziZ
e4HrocrKaIyy4fJdw1RoArJQ56Scr2b0qwiGqx+iE3xEHLMXaXQLM2wlXbJ81fop
2enCyZv0sFxjDVgCjXu/m2QjHehj8bxg9GPxnrxG6HE33o8Q8LzOAKVYERC6RUS0
fH8XxiXdIfvYiVwJs9gvPjayXW5YrKLSEzwqeKIR/gtJ2aLj+JAysEIaeqPixg1D
q9GUeD2aP3eMlLCdPlMJdp83WbcCzgHgCQQ760T6oE00jrMF8WaNNHz240CtbKXZ
CH3p+GBmdTvKW5NTuoAPlpoy3QlMse5DhooTH6CYgGn4CadE8goLsIytpz4Qe5SV
8MMDDh5H9mfsV/6J/zBThGDOTHnAyJvcezkokCjJTj+XiD1aRYL8xo0c2SiP3HUE
XB3NN9Us/zcrLqmu9aQMiCNxoVZzwEpq20GQW5YYHAHwW2iLMmGCJfuDMi+2LyVx
sw2O4wtZH2UviCpFtbPJuUc5/OnM94Z9aEknUITRznEf4CKvv5lsh6Ga9/DjtOsG
s7KAeOY59UcQ1QzZM+CwifIglc9ittOU1z2sAo7jb9VL43BwOtcjZs7tYico9iGL
gHYjYqmDGgBEqG+opWheHk2F3IoKJC2GJn4xxyZgRnkIX61mQ63RC9jrEetRpOOH
spUyfA9hXXw0PbkrSOHjIljzMI73zywrXp8xsPOJfCpLRiqPbX8RrbGqQxRk+vZ8
g8+eFb8v1PcztbWgiyuGWPhYRJzVLGnijbAwXSj1iCnYLi8ZpYYgB01OfQ6GgRNK
3KWlB+tlk9qcCGEnfgv+cM2CyLXUSn8rGYY59Uk1JAX+X1fczX4p7D9arVka5Av7
P1VSSQWyyAvy5VtbASBVPzliiss1u5gPZL0k1y1wrmioUcuBQFziw16F3SMV/83V
oK9uxgvTqUNbp1V0OpDkIDcZJ+Pt+TuBJOeVZvjtVrr+zxmwzm5GjqWKK5MvCSuo
DOvA043Y26bhCW66fn5aqTkLQHmsZxkv1Ec6+j2uUUuBk2KCH7YmXeOoT4jBNjBc
kBnMhplK2dzQ9GyvxYEYV7y2LDJpT2TvUSABxuX9TQIPntAIcs+9fve5fpIJeEvK
hzN/qieVceboT2ip+M7vxO9igD3JpMXBLQPFlo7hDsDf3Ccx5+JarMBfZgduenQR
LLgWeA1/g2QeS3hpM/zoAoJqvf/UPxzfxahx/7cmy+/X65hoSn3GikBekd43f7At
SzJ8nyptAr7jXHcfo3ayLyrI5/deCLCJ2pj0TeHty2vBm4uYH+eaNqjCM7tfv5c3
y/7WNdvw62kosp7fwoBvMcySC4HlIz/iEB7fBXZvFLFkMZdImkf1b6by+LRCruNF
/XxzlzJ+yw4RMDGk1tg99gn1EC3ejiwuMQs5HLzOfUgCmMVNUMKSquHLr9HhYd71
3DhF3upfppS105vkaBZ+g66JvXBWDwuPd7z2S86cwamShH375XlXXqvu4y+aSBwC
iBKdflw899AVsjtIbtHbLJEVwzyMi6e7cMOVnI4rE/1DOQ1niV2AbVx0rfDfz3pr
hL10JA1AVX/LdrAkPCYVDkBXledlkDr322++M7b49+VY4IIVUxma5UFC/zQMFzFO
hkaTpDdRvOysnMHRUlItadIzUPykh/qbpzSRGCC+uSZg53apIv9sZARC/QvJwIFT
YZ9heE5DE7wQVTbP8NMLj7ADDOYEU9v8Q1ya6y2fIVlvTe8flzKQcONF/Lk8ZRnS
XqdetcPD81qJsvvxjI9RsquNrLZsOy3fAyUtX8fOeCfbpk5HyBiLR50N2p6mRrLR
hvRIcC3nBi3s++uNYn/r6CjtaTBlp6KDxLdPeATUTxp4fT4MTe47j2/Bnnp2sSl8
pwoOv13pBddfTeQPzsUwj9evko2IN5QdhS7hYIvx7BhEM2fvxxn4KCj0XGKocDJe
vd1+oPTsLjEag0bs/w13G9sLTy+m5vdjm+nWdmFRc+b7EPbMyfhMgtp7Co0LTCgG
HhChdHznoVR8Q0Y91kh74s3+qUY4/2A9bIaTffx/qhkl2XisOJTgT+OF6GkZucPq
Mdg1HtOwjZS3PO/BYZxKjW52Z2N7u2a5XP/OzNQJMcdFBgiNknzAZhcke7lNFunj
RjWafndW5jnchUftvWKhN/BKsnCdPntM/aiIRXTupcZLsCsdKkrIuCuhNastushK
xmmfLRM8de8k9LAB374pqH6pxNflme9andXvmxjlfsTm9BbfhFG48sqywxaXze4P
tXeQ5Q2HGdGZBW0XMt9Z34QScQTcNb+at77Z5Y81F7s6QCh1rNOWcoecdXu+yzhy
44t6fJb0U1I9gsrUPij8jrrFIg7BH7288UZ+dlphYn6YYyZDQBKuVtsYa9yGh2dR
jBuFmP3lakRP29f/8X8peCSM9C950uiQNkhow5+iF0CcZmd457xruuZr2XTVtezq
N8woyQTpLWF5qQi0Z/i3/IYtOATx5SSW93OWv4FjapDbpTVZ9/Y3FG+qq2Q6ytXL
VruVCqCJ8Dxs2CHpQmVo+LIiIujv9PN0pHlloWaMk3KUkVnlKFECemjiSuD04rzS
2EZ70K30+kC40P6wmE2W1fSLJZciFq+2F7McWtnpW/wudPOnJlWajSFNjQx8os3u
qGG5de1ON20hIowb0dwnGtfVZzr2gSviuOMXYGn5F83bEyik97vAElk8JzyCGzrY
PM83M4yhQpJtsne8U+wvbKVPJS54CCCUFPCEqk4EpmIayIL+Q/k8hdfNUTGUKPUi
WYntadWx/Wy81o/nMo/pFKXeFv+FUbu/ie2YZFn0g6qE4jnYC3b59m3PZmOuecgt
sYi1LlSUO7Wcwyr3Nn7gCuwsXsp+fJd9cNjbzKjE/rSOOaPwxzE/Fa8qIpWBdAgk
JFiWxo+TxfRVqL94zA5RzP+hZjI1rLrpoTv5qSiUtri1Ksf/YNwGBUt93HFTAZPX
zYaVjajJzmyKw2NOcrftIaPnCSzOytEBa/HL3i9Y+5hbQkARazkcMwNtYqEEMQj2
WMJFGHdyzYNyS7BzJ9aSriI+ASU9iUQ9qcIfXJRPwXU919lFYdnN4mA92CacdXAk
wXXrmsKE19Q1OJQKk3/Cao5bNgRoEnaHaeiPRsnEa+GGnhrAWkKYw+6xb4cj08vp
MzpaTUR+KJ15KGEoHYQ6ZMn9HXHuC1V9RDE8WQ8ZhyuYd6J+c2w5H63dDIGWrNmZ
K4qL/GRrlagq/Jin1GdsHpJisB89Am9WmqPnOHKvwMTm8kY5ALFoBc9YS5zcMy3V
2pUSNLWhyOCz96c7kXmn38BvOk73yrUhlhfOv9WawgrODS0D3OUy8qxlHDHHWdqW
7/5CzzPyvHn4pcr7ZmTgff4vMmGPnrwahrtHTpSyJ0DgpP3CGn/UkXRjQEtSFRNm
E2WUzZtLQeJ5QbIR8++vqcF0zB1QysVibAuSS8PGixQkr5L2336Ln/T2FiTPgwOd
Xt2uP1Q0Eyp3Rekbub6N3JmGWX1NDmB5yBgIm8vb7ZdVMcFlGymzL7Vwtc6tSGb+
Dw5Ew8ricKjzQMTI5GSAU0gowfd+0uIrGceseTTE/HtTh478zm/3n0MO9pH6MtYk
`pragma protect end_protected
