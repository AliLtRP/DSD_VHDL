// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:33 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
hmIHv2zb12SnJwsCo3tG+/4zvTJw7nHPF/tQ6K2HW3T+wQLNC+3mTt0mphWPIHW9
qQhLqEzH/071WKo7ZUQS/MEJ+npOhHdkPpogR+qMg94xj3+qi2ImXOQbCycfoRB7
9rXtxB0epbB6UrbPdz5z2oNFvIMg+UEDRrFlz9F3P+I=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 19120)
RJzqB9QlirsIr8PN9eWYWu31O8LchhJjEB4lwfwCljk2pXvl1KPmc0Ro3mNCu5SE
2YYXPjZjU+kY7E2TS2Zk9TxbPDsZ7cGyj9ixUX9pxBhdBnuWN+x0k+hURY+wJkMJ
Cr0rEsmPXm1yR0kRvvLaan7p33E+1aAYtxRLK57+uzlXRJTfRLias2xATHDPPDXa
4qG9tz0zk0IRuDxIhrqhRdVQouq61ELbfcCG1g2As944aorNVrZquFZcfM3x77uh
jYiZz7JUy9QhfkSaMsI0Ov3TvTvVjFRQjN0rVdAbuEcUop8eGFl35OSg/6R3lMMn
ohP0bZEpAKuBsxwXqNaBPpPf55Q0dLZLxudZTl1li7G3MG6szQud79EwLSM3x8fC
AiWQ0iKLzVC2x8VxpNRv1mfH5m98Of03LNprHpLB2SrjsW1eNkHyVBtuI3V4ehck
AbMY8vTgCINyjo+sQJ8vptA28vvhOpkqm8auoSkf4ZbP5BD65mWcTSKVZm38e2VY
zGRBYxkh+aym+3Cy2EpPW62v0Nj/mQp4IwMUtc/mMmRVKS/ofqWtvwCyvbkIYboZ
T4B7WrtRLeyYazS1kfTmBvX25m9CF+8nik7hLEgiyrf3dlMLKFh/7DQdbNqB8JSY
wwEPyxtJevBRvxoQ7LrBuXAfMj2LTdrOsRqvQeG7TPHGQtzxhrJwwFSNsHSmKHFA
dBzZ/I5xU49A48vX7YUiTuHLMJzvd3WgthWepQBnkfdR2CFuLDy0XUdPWrVFrWCT
T5rU4NVeOQo2afl5XL/Hs84O9wZ608HvYq2p7LHjii1aTNxUoJMvub5gxpwvSvds
e2jbu2nz+09a+q80CQuOPORLlDcQoE3Q4JuGhtmmyoCMcuTVqzap/34tgaUtA52F
k78tUqB8Fw1SbeLhzJwv6mu4f9mhYtcrnFhuy/PZmbXXMYHgVYVF5JLpCb5PPHGd
IYIOIO0k7e1tWQ9TUP9Cz6hJw4JhBmw3t7MdaEt+f4gC0YnNMuM0/iXFtoel1eEw
bAZXa00Ts4kjNJC+sFkXBd4eCct/ahauvKIrd1Mu7eDxssVCajJeXbudTxBve0y5
wGtCl6sytcx2crCfXBdMctPZLpcHq3XyCMDGh6TxZr8HvF/IfHN3zjBewrNXIFES
3nlxiLQXes8Zqdwh9O3jCfg0+57Yh/eNpwvpHOjXClqObUcn8YeCntxRDzO7USdy
2GbAVqG98zRFnRzysuqsqUab+LBT8OeYrV7UNc5iPtOCiXoXAx0u41W3uwY1t0ja
2lmVe8WtZf39+5k+EMEA/Z0/+OuK4CHBPz+YLKPy11CTag0oSp7oAea2UoBZNUZt
1Wo17UtpHCsrcgA2fid6ifF0Axgm2UtjQshwEYzqprXPdT7hcNx2QiDfx0t7HBdz
R6YNorp3BzjMv+IBUqX1d22R6kQD+pxdeWGJeU+UOgda2zKkcs2T4tTCIZ79YFOg
PvVM5mBTlTwFSnEzAfSf14cTRIWDyAQnvCmthMj/Ga6zErXB+ke2HJQOSWksNlDM
6hnSzFNm/dqPdNRUpLe921QEsLPAO1JMJeStu4lLtWNI2cnUjyogFXQxobWI1Kip
nkXDzD2j00WAgZLDNQq/5jKmIWWSf3EZxz47bSWXGE6dAGwcsAj7GwJjvlPEUsJD
JDnva21Zpq4Du3O5egP/3D1vH4j4pf/83TEGYOoXroT+Mz0/0q7xifkkk/HOZeqE
Tvqd8sf5PTvTOsrgEsZ8UmuZE86ZC656ouo64kmZ1Tj6aj1u/afOTefq41eyIwRC
DpQGUeaJsLsMoiaqV9D68/19LV7bHt9HIrmU9o4/e84fU1f1BTlRv0/C8zAFrZdj
8cffErSZy86fp1LUMPMvNwduKxfE3Cx0i3E1w/MTt8xMM+LOD8A7fEmeR9DIur5i
JWD75X3QyQbui/bgxMie8c3GhReBTtXyUNx1IkPbdSweZXywl74pxIw5UGBdR03f
j95qA1Nrr+sBjv13A61lY5px8AnZLz+1Zq5rJPKlM/N6sps06Blh1MUD+Yg6yTxX
f/qrqjnYAuCKVoPettMbVm+kYWjgsOrE9+MQr3Is+eZ/1p8bpBI7H+mpcAr0gK2Q
ScOSjM9D9L+BtmzdkRUV/7mim75NynZQTs2vLtpnQann3e1u/UD2ENIDhSP2jlBe
jqO0iLp8t/ogm4UVcV03qHRrTc9PlOWCnr3+gX1H7PSTEFFXwZdqA7Jq27BpOMrl
xhfXxhG8XKCwjF/RcMRRHXRJknAq+JOZ8elvpO6jRrFyqxJI3QapvrmosfUFjnBU
ljEu+yCdpKIuh32vCuYbXZRf+1+ZrmPLrCmmLJZYkWy74z0MMhXfieS+5W10LD27
3izOJ9AUD4wydhELcwjz8acJXGKjNe8/tnfCLS+3AwY/5jku5n/6ia8j+Cuu0gQj
GbdSh97ccxIEnpztZteWUMXsB7nwY8QrJ6sF0nTVLeXVf7M/Nbj3y1h8h0+gW6pR
SIf5NOaGYWo8MeU7O+yE1i83bW/8v5PYa7Gqi5WJJAoRmhIA9hc2kUWOxTI7A5bW
aCtO5Y3KK2ls46ZQmU476e5fDKiWcTfJwyijtzPmW5eS7KQgwKqpuq2nVdysIU1L
5/VstVCNjPrjT+bN/f4BolWFpR2Hj6IQ/ZLAQy0aX7m+rHxHUHhCb1+uVuoRj1X6
PdIOb51JFpmhpqbOb1HdSAwqpAkoSnRKhoDX9lyXIZeSrjSDeD2dDLKAbOBctnG3
j/7/94e//6L0uDi3n0n1it0iVD45PYluOhA5ZWodqt/tgbaAswT9dVJXl60li+Fk
V5c4BX7KzbNqItx6xafOMpwNvwqvpmk+x6dtlg4ooibzVfdZ3z//EiV7oYsAGN9+
2/oY7u4LoDJlSVUBJn2E5t3Gw4EhbrNfza0GUEyyDbTTIv8gw74ZNWoJOnPePj+S
4uz5UMPPl35hn2rW2BT2zeNBvBlaYvkHGGnr2beX6dwMbuOw4cE3D+NbAN+0gNlA
XWISUa/1Z9LJ1CVbmY/6z9VZ+musQye/S2BArrl5uSCn2EDled1Uf4whS6AqPJaP
luVtf1ut4E4BjoL9UyVeCL2Arl5T6qDmVT7a8ptYkGjOkxoFUgnZnrsn+3X+V/Y6
PLStz86tYyMxoDVDnKy8fdrdBF3Kz91M3Ptn/SHImJ/0XZ5KmyMU36cE7IoW+DCk
YuiNP43MeIVOulOxwZxZPXjj2RnKKeeUTWCCYcj1HNgKP19T7Ucp/MXeGoTel7mW
b94nV1NK5bFHbSFdk9MVcXC7YP5CCaEUj/Isy+48IXJdkXH81qsKsgygUWlw/xuf
q5IvPXg5R/qeH9cykukufJs0SbMUV2Aw51Ta2xfbi2U6yfm+QFxRsMjcDVrbVDKU
3K51TkwMocIpA4YN5xq2JZHaEInQZjDb3CONOBupN74FMQrqL2eV/aVnPDm2jxxT
ps/3AxeBhWYYYuC7O0lGtQnJzOIyXF0zlbfsFJM5MkjxfXwIx5lUmCJ0rs2VwvdY
fK30uBWW3Qvf9WqTGPzZ6r4AC1SRIidYowJiXWcsyYNsNnUPs+FvWpgSVrTf6IdR
HYUQ9Pi/7e7nV//+QtYKxvTa7qteluTBDg4zz6CRDVIYfE3iq6XJZggZ4CUOPQtv
/ml77Q0AEGrN7oFVodhkPHscggA/GYXFiyTuilM1OVlIb2NNK+p0DUldNMxZOWVa
xg1GvjSvInqrD1F8O1axd5yI6Dpyb1pWvWrRmUIEmFZA8zUW6nJJ0b6O2JmcuaNk
PgoAknTRJ/xs41oFicMut3h3BHYRnsBb6e/QsRYy5taSOEB7T3i3VUNg7ndVy80r
uiwcjH589gxYsvCSyI2nxC2b15RZu4Q8xsbDV8yFfcjecJjnDotHZqQNPwpbZL9+
VTRZPF8Nh2OfQZH7wSmh0rxNVnPbYo3Qu4ItSOgPbLjGD3SDpSYPlFACyugZcJXe
T8WE2sd3uBwXj9ZmdGt+g2lC0qgfd5LbYeoY7dTIu77yWYuJzVDwZ/y2LXzCJc1V
mRaVfX7iGbqDnUnLXAOQqpUg7NAr8pkPTZNdzQwdpdEKhIfE2mM9whS7tolGTugl
+W9HsWzMq1CVbUNEKhSDNw9NNabBv2QI8DXopGBT7+qdyweBfQsPwd3i/rJl2zzd
u8CfXsO9+GDkkGFxS0yNA8Wq7UyA4PfgbjK5h9/98a5o+59pS7urWopHAbsaUBrQ
M5VBAIIUpgmPjnnJ95zS5BXumY+1EARx9V3aEhAKXP7DQHQZDUNPNA8W94MpYDkA
kiKfMmU9M3+fY3HScscPDshzdQSVORD+OtaSAqhf/lwc0o/K07p07Me76FUT3pKi
rZdwieLhfAY6/7eaHJqeFO/S9LZ9zWgp5iY+bKFOIXlLnhUDqRFyPr05xAKvS2O4
2lPhOSn3vxRoJle/ASi0DTXA9hNQ0pr85eXVwrO+h5RO6/+4eLA9dJBroX4Hc1JV
jVNK+pEgHdDPQVN12+x5Y7WE2ds5oBCXeLzI0ET3CYe3KcXNgEJaRscNwWIX7/dO
6ca7sM7wEsH58PIJiyq9YkNmdPrjKWl5tAOsLNT7fMHvWLPPy6SGCMxAJhMxl6ht
XYcy4cjlaOMT8SUoWlIdSiAMvUgdFLVJiQnTxkxApEMF+2pbU9K4tEEVlK7+U/bU
kLF+oVoGZx642Iu7xcYSQKC1yKH4TYmUVacxArL0fXy3+8d8h2k6tOhqgmK261yd
tVIXeXDmTfX9v4BWcrqJpTDEnazMT2VC4qqeCz0YeXlkrSCG3TRpkQSUGmj6Ew3I
ktwE+r03xqSV+5r9MwVudq3xapPd/s9GIE1h4shDvZkuIV/2qlpvj9ruBQgu52cA
q8F7enuf7a+5QH0m87EaZy1AzaabNIcaP4tC0AT1scZJ8NJHeeS/gaZT2/ByT/aH
EAriLk2lO8XQm/ShKET92CWX2kbwDwwc/1AIEy7F56VX1ADJ3Kwi7jeTu5nDV/9r
46Mnn9trwk9UICq6ANLCf+HuuEGvGPRvccZyXMb7pigZ71RmuseI5L1gtMRz+aP1
Db4FfQcrlPFLtTdvgHjU6M4MM3ShkiEiK16q0SKeFxr1WBchDelMZLhsV1+VU7bg
zc93G0WXJ2jXnQnWXfbDmijInaAg+QN4DHDLtFqlZFHWTaamXTcZ2qJecUElDp4F
N2vR2GBqcDoE49RtwdcgvF4mcMUF6TwHw2yKqzfniKfXmo1NvwY0Pq7rYZI9yVsW
4LjZLvNCVZaB1qZhLDPDlTVQBQPPN63Bsi/19ln+zJryLWDZRSuk+T5fNHx8DIqt
42QGFxc6hKnjsxpESewweIIP60C121r5lQ6jhoa07ECMAgi6YJu0uv7x7i3wcH9/
3WbIoBXDURE2xttUHYzwLFKq4PtkfkXffuc7F1hJ0xux039O22GWqKMU/UPK3Qs8
FgKsVgDZ2Ke4Oe3ou537YHebKFXwc9TudUWxk9m1rztV0MznP3wc3D0hDahvKJu6
enRxkeCLLnD6BUCdOOB5Odd4ZtF9mpQxkAx2aL3D3SfZ/WxysrSfkFwV/0Tt0hI+
X2NHCa7dTKDeIGAOqKqfp2wBsx3s9Kuh4QdKG3Vp7qKkfyZUNuE0O0scixyZFcgl
0nRWF10wFG0J1/m8xfm++wVntCuKrIgWJaT6YApgT65rY+qTy7N4HpZr3ZeoqVGR
wBis+nR+i4XaKzfiB5TS7OafeLDZXVXEQnjTR9BuZxsULuDO8eYKJfVCwysTE92H
ZlodNSD586cMv/6pOOQiRjXQrtdV+VmynNpNARVMtXwsSxrA+bYl+J20b1etmfCq
yxZ1jhepVxUMw/lk6udUE+rhLKLZfCwwhQDyaWpJR913+a3VMNz0tyOT7Y4f3hFn
dMD9W2XO72vI581xuJsrzJyuxzhfx8De9yTijidDFR7yKxXHcalgvSS9qsKk7GV/
IvnHa7ICN6ijNcCWajnHL3RaatJL39dxLOL4zUmJnIg/Pmvmp05A5Vx2CAYpTcaT
IJ/Y7f1ABA4DHrmUQCkbuwcE7pt2ISHILRJi9KWl6wpn5pSibIBhyzElooMxkh6b
4LBCpOzZ5PSjZnhYrSrzyeom+2sVXoyn2ZvkaEEiqGoFJYHmMJ/+6hX+DlpFiE+c
RqoxFd+UfFzylzH+JKla2XAWDzXNpWncGXwhILOFE6KwIgx+AKgfHhUUphK9MlNQ
XpgFyE1pUJ9RyXI3RmRHt2NAak0a96VsVxno+efe8bA2p1Bd+wn+2+MW0wMFuUpA
kn2o91vmGzDB58uoQz1hHfir1JnlTJqU1bDh2MKqEWTTygCQmuREDzinvaux2o7q
GZAMXwxmfEugCoIxc3hcb+r9ADx6FHtTYNrUcnfxdU6WlBRRPt96hJcASmmeYRdg
6i2zkXnaX7+aXYq8ftpnHQadiIKwybPkGsrha3oV+l2IveTnGQbDV+BxkEJlRjVy
RyezvGNu/LVW4C92OibUGoqODfzrRNkSQ1wRd/gBXEZ6fQM7H7zYzLuJqMWmpplu
I1g+JaBvGMdhPOTj3h0eDuFD/mI5wX0VcKZWgvGwZGSUz4GSlnkpTu3KvaKRM/yx
i6/sX2RKDWdB5bvMZCX4FwccTGlj4uslED1aBCNkBUukTMaYwKaL75Bo4p91aH6v
sDHRwAgktXRGZ8ofdMN4gI1ZD06Sc2vm99ZLJ3BgrlYwQk44NZBwWpCsCVA93AD3
lgMNWZLL9GtVMz8ohdILHYamTE69neGn0UEzAHcZRXoGbQSsY97d0bwpjnDy9o12
SVX6XB7kd4ZwgoiXERyQzuub/SoluAMpg0694dR/hEUoM7M0p/RcvMCw9FrX17Eo
N6uRZMP+U8zLIa8OlV292KuR+W6+JY7v2GFWQlERJWufnvoIJ+X8witPgXQvv78U
SdZThI8kuNPhGTE1V/XLtX//pXtLj5s1Yn82swmLSx+4ZCm915PJYqb45JMW+dwe
hFO1Y4YqtxWK0rnwk+59/G1SbdArqsTzPNkSWjuvRujCpTCrJ3J8ZTIIJcYGWwLV
22P8dUrJJVmuikVi+fmlZR7ni0xwm1gdHmnU4Rxut46kXuCNuGbmaog2fDRbFLia
jDQXSgTAJXWJEvORO6gaIWPXOkVrkxk7Qg6RSgeK9A215gbyw2+Dz3gTVS2jRGLs
oz65G0KjyWtHuNrLdZQ2RqHtObjE+WqL5dIZYc1mPDJo+CirU3BFefNRFpojJKVF
HbjdZ2XJaTjf4lW2X+GcsP7TBcsBvwah1mFheu1AM41RGPSXDotmN1G6wCEX5/2q
E+OgatiMqgaWyRMNIDYNloqBFyzkH1dvBL7eCvn3CimpfOWMXpma0OCTjLrR+Q2D
fSks92z3fpmPp9l7zfLT41Tn2mBIWYkdQPX609wdJJtEMwZQwSSqs5fR87GxzeMY
QMXAFcC4O25hqTaKanEo8HadSooM2xyjmzkrBPBSdG2C/nWINUA8uDSxIl1xGjcn
fkYMxq4TmHrShtvXyK1iyLGKS5Cx0X5L++xtqugCW8EllPQobuh70gn3ftDMaE0f
z4EUnAFhlga5k7ekXgy1ZDcFkQwPyW/C3/1aoOX/0NkmuPOC8SENtRb8HSX81B1e
Ly9KblzaDmrNgUYpmW/rfETp8OVzpciM8WijTnG49pO2j4fiw8iMdVXbhXihc5Ov
NNUkL2tSFvfbWZF6zHWLeNnv482DdOFV3rhpZA8WN/6iQOSRJ+V434ljB8O2yeIW
SbKMtIV6JNiMfPH8j6HK+n7b+O+UYl7EgCc1oKq7Ik4Pr4q6A7wuNdpvYLpsRxoQ
s+2miZV/Sbutbsk9FimsZIJl83307BrHwEWBoZQ/4BTpaGT2XJIwkRE1ZsRLYYiY
zWWxvEHw3BTizdMkGhZvEoCiG2/giJ8Igl3ZVxQeJ+6GDY2/cTLIXDB04Qj1LCdM
KMRpV7bjRhNMOBPcM0tTbtEW3XuH6i2COlDH+1WgPC943z8DSY4ZybkbU/2/MwQ1
sB8QKSVJ8LZGnltuyjO7BTOaRfz2yz2a3rPWLOe5U1W0Zy+bXwHRpXonGQXVCqty
JBBJo1EWPlN/pr27Ewnu9SD61QLZY4V0VCsrBAuuNSOjOmyXCRcBuHRP02Clv4VF
ohi/pNJfFvGE8tZtSaEqIBd6lz9RqxhwFP08Z1PlBDulTpFM4B/VOcUp/aIfvAI4
3gt9p8e6Aw3SwVahwWum09IQkRQ90yy9R7ZdAglUOB2iJIRuN1XbpOC3CPp11HBe
Q2tVVfUIGpK7cMjbG9AJ09sOkjUSCxqMzWcYpH0k6k5dWM5QMssSEuIpWhXc/Fav
L1ltRS0d0/WzH/dz/LacdKYFs71Ri378rln5c+3MBLpxfxyZgwbiuEZtmMovWis7
YXVwWvSX3rRFcqFGrv4nlOQ3OXCg8/QKMaeWtQzDie5nCKiFmhDxfX4sqeaFtRcx
jTcYo1xETXmwSQ83/IcI3baaV5J/EILV0L9NvN2Lx65kD/41C1lNkyWj9Xv7Lr24
bleunTEI/KRQuScMYEF3fSxL0THHvDTbgP4+SgqrEU9YeFZ+hv7QeMSco34hxF7x
oiDQXw+B8mPw2WMLi5O8xOfImaPUQLjyRU0Ubi4eyVHlxPWPrLy9EVi8Xvy+7JOj
jzgRpAq06Kyu6JIiNohlzdTqT7Ph+/3RlMc7B5vwkyXOoHNvEVzVXbyA2apw+uqm
q1DRCtrpV3mNWbTY0RrqOH9izVmyVnA5OUXaGDYEnUZeu70szCixpe5rwiqQBGJZ
QGjQyrZraw3hR11s60G/UGYqv7lzZ32Bz3E27Y6H4FYBxZNmCHiTiY6P4zYDxDly
CJ4idLZO8v30ojSzg7i6T1evkUg53Th/6ancdmTSzPHOM8kB/L/BSGaZTx7HOofj
6gKkdm3DxOEx8vz4qKKip9NlVAs5rtSIIZtaJffCdwx98fXrXI2W7SToT7KFzN+V
6kfR2xVS1XHsBw+Kw/l++xvyYEjRjIei/dahhcS+9T91dlKhjZ8lKu9cMjDH/12x
WhiTAcIATHE/ZBlJWUlFcEvNkVdX+KKEq4C1c4DbcLRjR2NaXEWQW8TzG0aG68Hv
Rg0DbrTp8rcQljvkKUm6442ymfu5hrXXUSFUArr2mfD5b8PWQ4a+lvNr4fgJThcc
i9C0jaoTPkV5j6jeWjsZOFrxu07SX4V+axlAvBLGqIIH683ICb38SCIspMqkgSFM
53iTppybspoZk1bcAeEbmlCfbo/Wnjvq0NRzxxVmy6hydEAT1lTNRgsrZvvbRwkV
3OzYhv1VOi8lv40SmPNdyE3LVzQFWqQ/YabqF37aVajYil1yxaESqA2Bm+DMtdhk
hV8q+o3OFtaOe/9RjO3K65zjntENsYXJzP0OetcPa5UYiIFqVUBdBKpVslvJ1Ha3
isrPByfwAQ8whuzjxxA2/vV5qjoC3oWIpbns3Zmau908oXrMTZ74zNOsMKtL5PRD
AvlNoVcB3sbICzyI3SyyC2kj5O9K5sOuA+g+XUzd1wan5K8uCwQEaBZ5Qc0TA7si
8btJajTqa2x4/ZMmIBU8ngDu50XzMkHiL0bb43VrFGuWZW93aXir95ZkX6X1PQGO
ZuGJtcKDvcjAFYlUzTAgteBKl+CU6uRUCNrtU9fhfeA9YFnzo6AFBc9pVl41y7ZN
3d+JyNy5O9ibsGD4HUYcgnLzEcJlrKhsBidy5Cm3Tb/LP97itEQp+cwPIP83IVUu
fMWTjn5NolvJllxVp+qzUp/Q/+E9DT+MhfjKZSpAQQQMl8M9zAwpchhU/5h+YpyO
66M7ix4Z75mzJWyOcBfk0Qk4UQYNpgK1TxrDHyCgCd5fS4qjMGqBD62Mr+6OhSfr
hjGOsB3k7Xi2R2E3EOmYInH6B5zUs7YadCn+ULMX4/x2+omZo0/bhY8qKPVmjBu2
2anKW6K/SU3adJEiuXDgFLSY/4MVr8hjjwy3T8UiyFJnVeJOhrPR1qM/tBdTnOaX
tH7Eq3qp+sCRnKDQPF2llvUyrdWhcM4EIbRf+cFq/V08vcvWsbPtW4F/02MD6oSp
h7uFMcW9v6GnbAgRuBMf0OYID9P2eG8x+V0G0Q7VJ3zQ+CrOQeUflegTV/Ac7RU6
gKNfx1uLzNMSkO1NJHMqcuK0c3AExzxUk9L/PcRlVBSJj8+Po0GMFaNNs8cz0s1s
H2jrXWkBbNP3sqy/eAzzA2IqqlWix6aRVIpuh8V5TyHa+yLugnIdk6IG0mdCfHin
79hE8SXHYhZ8VbrYBAJActLaczALbeFjwYz0B/Pll/bSwm0402jFZ44VqfrME1MF
UjbNnYUEnJyZ8YxcsWakbU3HnuK8BHWDRPNUWxYE4nxS/6V6UzwXOaujDLCQsiDf
831vYTuDkxeihKvEoO8sQlCrKj8L0mZ9VgJzfYoWYp9Hu5PCzXF23qCUAVIikOqp
0g/fgpgBN+Fasp1KSGLjgcuW1Kc/9NwhyzmY2NxoozVD8vFQ8RVyxjWMBrXgyyc/
DjiBP9O5aqhhvYpyzPdaSUdh+kPDrKO5DAfH31QG0ipzyb/Rsb4Qu+JRn0voLAEA
TI1Sqpc4hty+P3bwWjf9v3igb8UBCIt+0kRm5Vm+Z9ySj2qNeDAnO8KrbMiCwLnj
HSNv4X0iBQAtwjc+diMakjGE/LFtUySICv4uWmyZkeYT6iT0rnJg+0Nr1/c+GZe9
Hj6pePbs0s9EIDR5QXQx81/io+Jek8jpILM1sp7xfsDuix/LnzYycpeYoJWxYeMq
NM+6Q5zzB/lsxWGUTlUdQimadhSe0ijNIjDDz5Nvqj6utTe6lYwGAr3hA0LJCXaP
ScovvXot8q0Vx/fpwrkIom4/BOLb+yQLdPGyxn7xO8ILmwpxWBGotKZzDZolgt3m
k4fcWRNd4vAOBCVeWMuxCIhADpbxl0Shma1l3pZy9U+O9GjhItfnBb3A9WrOS7wN
nKPTOxCBYEHQJR+LltaZcZSbSOe+TkWkgghVYboX4BZwytXfsoI2T8i5vx0rRL80
YnV6tPcu/3OOEK2dQD9woLPOV3ZuLW9T/Y9YyDlBIqEuQlixR7tbbIrNei/DOMS2
VAlcByADJT8OvRuuzyM01EEONKcSoG0JT3W2eSCqx3pxFs/hRDukdzH8C1nED8Jf
pgGmB0JXeGkALBKCIwgcPNhfBxNHeDe+hxTUnnziBpN1aPKbcgjRWYvWAOUDlBmI
MszBry5zgltSYl+Hc9S8TJ4RoKavrP1cMWP4CIb2Qy259WGbFezJFhpjj7a6UxG9
QPZbeKKlQYwqZ8DfVbQTP7e3cZZSwRPjvHj9CfKLJqPgQtq+LWbpWEx6ynWZFU8w
3PlUxwZoghR8qQ8nOmxwYqeXR8SQRRl1OIOgya2OKMznYHiG8zPbERRniF10bjuW
UcOc0BFYvNzUOcsYxVqci6icsx9o5YcJAUp3yo9PwfaT5gdb8mgCNPM7meJmFaBY
DDIlZBNrZeaTLUOxpWJ1cra5TqimWEy1Ha7ZiRFY79ufUXAP5Mc0eakP4z1qoF5b
thndmIUf+Lq1AO0391XaTGqLMW8ouyqcGQePCmAPUiesgnJbMIHG4fDijfCYZ5zK
FrdeGZh+krhtrjA9n2jpyyOPx7Wj4lJPRO+dRLXcEAB2myldLqQwvG9y00z55ohM
PNTOUe/iu5OcL550NzytcFkvTSyDoqZFVRP+cNioXVIL5Y30UlePeM01/HuWG6Gv
WQyJ2uV8gqHf9S6JBvkQMh2LGUmJcX5q/VEdKoZ+EuUPfkuf18+Au2pr3soRsyaB
xUxuahVGMwa9g2vSMkvGTfppcyKfBojS+UyE0V6sDb5anwYToJS1KRPVoWkQ/rBZ
I8XV3thUpMYzxpTrEXnvbjVYQea1cbTTOfeVX6I/76xe6e/ahdGZahBgZX2dHA26
CtxSghYzhGqtoOGhDa06GlDzHwWDHaPiUonvM9DU94DKR2r8iGHVdNUtj+pzlyFw
YpxC9CUPqj05N3m3kH8a3T38bJ+O/zXi6cjPuXyhSlrsmOrinVfWJ3xXh0DTiJ30
Pi1I3w0BagMs1cj1IQXluC5bJanHd67S6WcO1k+MgAAw9qQT4sA1gWcWT3pvFrHj
5SDh9INn0EtSchayD/AQUmpctTDcMELZ+dAvpNukFpiwaRYk0jFZYU2dFsZDa4/V
g9JlaY8cmP5xsKnPFlwfFJlStCLPxwf54qvOaydq0z0wrBpStnsJqtYYDdcoKgyS
fWH/ZI7ALlnWtSD/XVwPVx4YherqJPD+LfrnylnV12fY8qLU9VRsAiZS9CJVQ/rs
NawYQ3W6zFxQkCF+VOPUN5sxVb7jBs1qaaEJgE1ElamH8gh8JcaBS+W54/cIqc2R
VUiwazS4tozNY6pBpm3akNULOi6Hv7oZ9Bmtv87vJTlju/pxPllYRu4+U4ykZKl4
L3mlgUTodguc1KabH3ok6R9lgoaj3x9JpsjPza/MWBbwHo/kBF5BZ0RKCF47hwAF
aD9L8dUSyMAI/edwr3zS/QW8u4RV/wcK7FcYou4KiR1AL4tRMMk3cSCWyhp5AqGT
8mUjMimVdi0r5TGV/Zan0psXbyvDZm7f03rAEXqGAegXj6JLc2GgKZT7jxHkFWiY
O2C48oMu/yCHFT28o96QNxbR/I+OouduZMFPKLbbpBnH0IUcyCIEY00m4L56UXNN
EWz32hUfm7UClnVZytM3I3I8wKzCdXjg76/weC6GoItFDmGbuXtDZNHOtbfJwuWZ
m1bAQSaOz1O6Gft4F8qnUyaAv5wpMKHpahBxV5KWVMhnejTSf5Y3UJrBmCeXSHOS
+lXQZcbcLgzKQod0RU13O6o1N5BYO5JbfJPnhdyJ6fiQ0i8AlxcKMqzY7BVho/RH
Go553FDrdxiE5g2yzPcHMQ53hVNHNTYd9NqszUyxMyLIO+TH7+LmiFQvZQXubeai
wCEFg9ou+SBePYkep31FRqhds50c6TqS9P1dyBsko1MUBoeiJ/+DbJpolTbhNB62
zYDDh3YAaW2rLww0RygAVpCwgzOXpmu8RtSb/bZMTiXjVnqeIYQXu8VViYBwbKUV
6q6kkVb9aMPdTVHzlSynM7EJQTBOJstGQZNC8tIBcV4wxnb24fDI6SQMxHswSsfF
a5lHAzXG1//FK04Sctz7zhy5V8H4MeEzsVboI+dM+IrBGpJo9oMLhEvrlFhc0z98
6Js/V8RIVJHH5bzX8E1BK6F0DLW09O06XpY5V9+wJ3WDUTcqAWd87dGntdd5/jKe
y59ueiKAqPkpPJHq8vwPEwzQft7p5tA87AX0izFBAU9ASMH0WUGQmXEOlnSbfnWg
Q2s9/TTazLAAD5j8IxdThhOcl993GKniLO8p+QvzYP9nUqGK33mV4uWFAq82E9Bk
fAbSaTHCMKkvggeJ7RioKjOhNfUBRLdjUHLR28jn5gUD7JmmSGLfu2bbAWFDPcjJ
ojDwV0l2YjpgdJ0YjwLT/eS5l6sxx28ElAqB/U/cWcRLoHC0WNvq1L+ezVvnKwuM
wWa1SFCpxc7mGkCW7PTIJBh+HUzX6m8gv270ax1yjHGgTZ3yzHlvldFC+x99g4tF
X+8yqUuhuLhgrKavD27Dtn6YQG9cylzG1VURZfSKGIFbGEFk58P7h6MqgnVePWrT
a6ces/wZ5ONdjB5L23Zy/FOBuZsJDsNFcdRwKqjVlEtABmhB3SpWlI4gmXi4i8DC
rbch3HMNxIGLdOlxONYxWEsotxx42vsydCtraFZSJuPaogy5JpJq/CzrCYWGQGsB
hyyG3WrwxhIUhK3UqOWzOsxvpyDZLrMBqada/ri1rgElYGSGn/iT51rP4f3iBOqI
A8CYhDBWy9FWiSXiGR8peheaqq40hGAptuZDM4ARKCL7hN7GiO3daM+X9hqljSfl
Id3gCCxVIZ/2Awc0p6HYmmzR0KL31QzxYnngIuM8US0EwgcqSul8Q7TgIjIL5ae9
mni5LcF9Bf1SgNL0vLPoiY5Fvmb7jpn+54xBl2bK8afac1S3ufkRkvfkKyDaRiTk
f0FYp9RuoQT6FHwrpa1JsHr1If7HWdwr16cxNw3+HjLdkBTbygbLsLVChDAScBw8
7JodBjBV07NJNYgndQUWlMRfbNamsU3Ba+qdcZmIagcytP4wS3twUigAnD/vPjT0
gr/ZtG6Nh9BAibtT9FfNgKijxAqeo/bTT/VfSwo6Ddc19gHfeq6sa1MKCjevUp3l
kAMih+zHJY1QhOFzvG1qDSTRIvSoWZQr7LNc0oGHZ1+p7XO5A1V6/mln3FjF3kSL
H7KtyCFsY8sUDDN8iyoY1PvpLnebaVGVs2cpRBx3NlvsbFJUDE026iRn5Q0s6bNe
C57Z6x495oHfV95SOoPGd3Ilaiz0NORQcKsiUm0ik1Hiadn4XnmpKPtt1u41e9oS
hCujJVkQdzlI6QOySXR9iXkpjd6zh7+5nrvdeiw1yBXRTc+O9szotGJVOTCUQcrO
5DpCAsP6wS0+Pk+rqM7OZeQkPHX+eahwMgiwVqzrjYe8X6Aq0AmRD1R5H7gLMcye
lcjc7bOqxqyQR6GAWZvUCep6XELRQD/obc3rfbxprUUi7fui0HwCcXjw7oh54Lmd
Xq7fciGagGVqMxnwHXGk21S/t7PWODwDoCuR/O/420TcuikBOJdZxFXft/yf78Hc
UOFJakQaKVSianLSxvpVFWpIssT9yPHo851PgYrLPaeHQMCi6pvZDdGhdnkzz6IO
PiNFVruIeq6DRO69Tip97aD1Z6Ucgpp9puRSnGkmFwZ5yXv7t5G+cowEMtYBiDCS
LGAkxW8wpqH71oR/4s2idyZjlp2LV4Nkzk8V+CLX8f3aumLpjv9OWwKHSIRgXpvA
jk901+SJd4G3vMsz5Aulm+dTtLZYTv91wg/jO7LC8aeAnTRco8TKrQB5IKAJpmu/
ruapcSb/ugqp9f2Q4MBMB8Za9/uY+n3w1FySYyB6Ttwj0gy9lblC+Z7GmY4LTgYY
GlYWNgP9srvj1zGtyoNJy79B9zdi4LtztHa8CQQ5mXUIAnvnBWU0QZ93zAOPyNYo
Jzk0EdbVA1IkPWVat2o6ic7xoVhtV+t3R2oAvoLp3Rs1q8avsx7oTfNcKwYfE7Al
t3ayAbLH/tu68zGfSBwaUwZvCANyPBuvV3yEz7GnaVcAMKP44KYF041g8J8VeL3n
i3CY1Bu2C6VBrLiuKOoL6tRYjK5LPEGFE4uGuOTBLTn/dqar40F0kMuwGo+jkbsd
2zs3tCcmIa1u1XOUeW/91vyjZvn7KBTJyHuPsE7DsCMN9YrGCacvI/6fcrzkVx0M
5xnia0fboPSVwqQGNWixnCMOj2tSKdNYv2t+WjT2Eb93t6MzM8SE31kUpqUbVhY7
QfC/gDckGoxnX3athVnkgqWwsNt1SuRPIKCqUyFBsHhNexnUO7nG3ssBQawaGzoJ
35ezzQBY7aNimVA9LWZSvkiMBG85PYzk32ZcYbOl2TzLPTCCvddB2+7sV8DO/7GL
p6y/kj1Du2Eyk3UIDLPxKWS7aYOHl/SyQ5R5Tg7jWvG4UVheDu4zdKh2BykVayTM
u8pul2VyzB6zNdBxg8gaVAlSI2SApP9w1dzQtBJrqStuwXI6AXJAI7mcrw+S2Ria
t3yR9nzLUcw74eVXockxKlbSppQRY+RgmoRfHGbeTuNXgtMByzcIVRoYx/MuPIsY
VSKfIBc0nlTCkvCitgG4FKohRAQbAO6i7Ld5XNiNRRMFNxwEB0VQNFlpjDjACo2l
4Y5buK2IF38chXN3S5HO0rbcpHa8oS9kPcn1xaJhJaa3MEpVYT8kboqtBGe0pJ7d
yJKFVM9nZ4niiogOBqVtvfZfEBg4NLoWu0SFMjje7cwaZCadaDD0lugcBcprCu7a
Q7nXjn3+AX88t5bQAGyHu2RV7xuzw0wBcJp1APi3aLmlhdfCb40qTERozoCKpvEF
aiNvDvCZnbLeoslZfx5NSlqVBuI6V49pR4SQWY9E9c+hq2lwskD+cZY9IhfN9PwN
Hh8hhAC+Fpn3p9z7dO3s91pKSRsUzyrd67E64OyJr4wDt0lXRjhgfSNParHM1qjd
7jJDM6TpotmngaHlKh6otcvXeHgEnkbqxM/Min6+A1PtaDMvPzdryoPtNStl2Mal
0EmLJMSEC7Pbb2ph2dUF4A9GNbNNFky6jDWuXIasab1LxjlMQs5x4PUrsDAZkePo
ilkqPn9AV94AKxMr6GwH2DUBUFc5RRT2DNIZt2oMgtJ7sHLWKC2wr+SVYfoyUez8
k+OT5N+vseX4oW6ROpovT+LRs5d5zY+hUibnWhUcPDaBwZRyaLn31sH7ady7HPjw
t7OJJGRcqPIHjMQBNYSqDlsrwQDn0iieCI+aq3pzO1gzQO/aqTl53DTd4qE2ZKzp
EIuXJM1LB+f+7jmkuTaG9wDQ3pir72vvtiT9ap5iEfIhtmpmSt37AU1xRz5JbU0v
/kBugrDhp8LP5iHJuY3MXCFgZRkDur0IeW1UIL6rXHxDCPWuEJVU7JbA2d30Pl7r
8YuSNFJ59NGJQWZ38rLvrLTKwslao/lM+uqkVaOYYMStQiPSjILYJd8FBJH5h1pY
pBjZjUEJJvx+YISHLfq5f+zFeDG4TQ3hu2bSl77lv6cFD6VG+OoBL6mfZ8Q/OSnR
vEY5dpv2sEn1SSEGtQ2qbiDw+IlLsJB/TMr0kyROAQFUSTdTZcnaPg92dKvsP6mP
dJJ8kSl1hKYncf1mwAFmatqHXK0J7b/XopBmoZTC7zr/PqQKOU9I1fPssAgZzUXu
2rFS3zoqn+NBHmB6qSIO8rtb64nSJY7XO9JG0q+ueDp+B73rEXE6zAXlmmCzq+3I
byDGNdtn+2PN55EaskvL7sY5tp4aRrIXWyKuNjEjlDsLYc+WFYGcdNcpF/i/WSMo
EJg/l/GdkIX7wYOXM6YUOtFiTB99csW2d5m4BJigdqK4sAJaLanOoB7Wy6x4J87v
8d+ok3rw23qmL6CNL9Yi507IaBBz1qPib+S/jx4VfwqFkqJ64ZyhwD8iR2tH6YIw
sqO+F0UK5ES/qLxNsx6Bc06Zneb1x1bsc7vWiCewNHw85nSZEeuN5lUqXIsmELcQ
EhXlzniOw/2ncYShAMvRshu3x+xqhmMOkEJTxwwRoLfbrsxzLj2wnmnJ4TzYBZs4
TCZvje/iO8d/sXsofqnSrLUKbjr1gHP2NH97nDwvTgo9CR2EnTXVFYQlWhO6/uae
L+OWmwajsCzgfoWCrHDFCdcYQ9u71QT7hnnCkBKBHqdxgi7F80v1N3dI8iCsOHHN
L1xSlXSO+QJUeMSs/5IG6RPRLCynjqmiWTXbiBHbAJGhecaq+fChl72y6b5X9uGP
Zr7eVv/sFKFz1f3kKTkw8ZftunblUYEXFX55OM2m6PcApMQJP/mY9Syc/B3lZj+H
nXVOgjpxAB4e+JZ+Sa2iKvbZgJN8aatbsiDmvm+y49lacAyomtM+h8YJEOJg/Odo
efXEz2M7ZdLokS8n8WqbBvppZPOdnYoQcIPhhgSVDxRDOsBZROAEQnsmMQo7h3WC
ao/dYW0N/L+SROmuThGt5k2vwxWVVj9YVsAADoMREMKjPrhFbUbexYhYlznf1qqg
xM0IM8Np4bpyymOeVNO0SZjZl/SkVJRMab8v089TIAunHQIavkYsA3kv3vdnr0wL
QQ9+PKjCF+RKuStviobdDvdhq1bjLiVJehqZRhhJ7jn9JSwNuN/oZgiKBcFbC+o4
4sW6Dc51dlt3+1W6NoHt8zSodJ95pBQ0PNwrCkfeaoqCKnQv6pn6AolxqlIUVKgF
kkVDeGHEA1YyQYgxrgbmocA28SUwyR49N3tbTZ+n9zg2TotYKgcKLU5eGoCyY1C7
E6445eI8tUQ/RjZHO3jFtVbVqCY2//z3yF0oqYXbqiE7OnJ+f7H0NShfDEwu02Aq
42Iq8yqDuldrO2xJGoGAyY1dERUPOP/rOckHIXiODpwal8ztoEZm7Q5/Anfw/Sw+
qw3Bp5Y1ZOW/bQXyFC5tpVwoqJCSZdFdG9hNQTUhNK+AB1hgOQeS/W7Vo9QQ6XtN
zh0nMT78LguqgR/796EoD5Fu7ohhgC/DIBGw9IHDmfBlP57UmtmFCbdl22TYUL9B
8rOHMhT4mw/v+JnHoEVLtZyugvTtW7UoRcE8KTXd/ogDSi2hdPAHyXQ0ypNKgCDX
e64YYC4SYBd8q6irU2vrEvaNMI+RnX84YObGjbs0HwebS/DvvZRnK0xINMFVVEt9
orNzBrIwPolmdkxndQoaL5ugDyjULmBpzPV51ktsnkGOf/OHyvkgFpC7pV7K3Xeb
7THx7SO2ZNSRB5TVUvPSEIWYMCTDB/sFR9rmk/PZeORa3MsszI6ElKuCle6RCoud
HaRMm1NYSO27/Dk6vIZue/ExWEINnldsdfF7Q9w4dU7eXMQb5aWwNnHcZK7wF4Vt
lBPltN7c6z36n1aK4TFLAfJlQuQvKPGfSMKxmEbjk/UXuQ8oOX636Cz4qIbpoSs2
nOsSmHsDIMtGucvXdDaeItjsDqeNB7WDP3ruC2RPXjHR/AAhrRpg+JzrlMmBy0ZQ
jZqBuQ72B9zrY1b2C9bYs2P9UnZHmW0dWP6+P0gmrdxLYzSFH1PHn3/Y+wb8/H4F
DFx6CQLwvmJ1fyynq9jQWvYiDH3korTVyv10oy74TzO1gPFMdjxBvA44BCRIK/SR
1gjlE1IEnGSlEy2Oj4cGYfe85WYjS6mcCoZNMDxzI3xlm4hX6QEEMdVAvqtqEz1G
ICI5FA3xhqT3ypoGsCCMZPAMC/qvTENOLEQX2JQNlIM8lz16UjsZRT6sKaD7BTji
eyrv2net56eTRg6Y2X6FtrkUCUPeHXt9z8xj62UAJ+JcMybZ6iUDgb3xBepGlGkY
DGvmYKxS17RlPacPzhkE37I11iUXKQ3GGUUqL0Q6IfuuZGuqyp1/+lRvNEn1rncL
FB3RvmLRqc7J9aWmNJb/kxpHeCUOTRJz9toOLvPWzMiHVrBncsNbNFwW1NmA9MAO
zgx3aZrELMLb83+KcOfiL5uHSgQVN+g/mNTItT+ZQyZLD0EZ1ko1pqKAr5G2V7o7
gAiLw7w3Q8P1vMKB9fbe4F/XBieOhqbZK9MPi3s2GOVi/jNyITIiZ7XECgbGHEUP
gJXY8TV5bF/7Cg5ILiQvqncivJk6uySbcK8MNNY5EKpBAouxjDk4wLDem8MFlONK
QaD6FJ7JCZ6axgbLzlMgzlKC5G9oIHTi6NGvaUmB/WDxkGvYC9qVBRtA0CHTrRC+
JpnhR27h7oXxhnu7FQzE/VUm58jpTFIYnOJyXXzp/qv0WsPTYTWqHMV7lPbX14xn
9i0QNfzj1qi8bKADQ8UJ3MBQhB/YtSZh67jCVyIBE/N5eWNWpNPi/CGL1XDZhUfS
HVbN/+jEuGgNCGiG/w91RZ0QRybGAV9/xcPEAtvIW6Hv3NRz9lHqjHXaewU7gSoO
JMf3M2xS35gTupQFcmr5D+4TR9d2YrlDF3FUXm7olwFlIH50ZO0x8G3q7vsQDCcZ
HLur1GQaP26oFKWoZneJfe1uA3SES3Gkj9Akr+l1H+W74iYpwnHU0Zx3gMbrJTGi
ORJP+Cbi+AXV1fV5gEGdkjEATldC11Ml1DBCVQvQXnLYjfK2P1w4Ckq7AaAE02Ci
qP+uqmICpWB8rR+Czp5A1zmsV/NICu3OXB9l7zXVCE0pc6McAAHfckxyou/Kh6BS
wD5bL0rBPHqT3Ayrn0kvE8Ke2r1iHYr6zvG6IP44uBNUper7wHQ1lQQPIimCNP1E
iUSzh7YwnybZnmpEY4getHROuRRcGox21FL+Kh5OOhZiq3Is9VFad628iA50cNCm
UVoqpjLBgEtPc4efK5Fcpx6l/VgzUjv//zbRiwpU/86CIhbqaGu5Q0kbFSa9oD6v
N0EFjnCQBAElq3Pq9uYP6z2Gwg+rplcBdaBVZrpNpVjJn/2Zp/9NTpNGDudn5uCF
JkGUGCVEaDX7GF3txHKNtDwoGlTLQFVEFiJlXeNyaqI7pbrNEicCojvihZglEy9M
OJ/EHr/loyCpEWmlN+qJdy7RVhuPD0vTMYkRkl5iGLIcYrrnZIN141C2NWaBTy5p
Ta5jyxZ/KzYZO4AaQfTFh9JLc7i05m+6A5Y4nGdiIH6gWDtloG+Em/hbaMFxcFSg
z8U/3XBU2ecYPVLbOClH/kOYmbmOlJBZcJkPXSFDdqyrJZNgkBQiXRs+0aXCj88Y
709HNMdNjCu2EqU1Q3d7+u4Cr2NHsTnLRyWTcOgi/ph61aD7zDw1XBlCW7GJkAQr
TLvdDTdb3ee46mnhOTkNUxh/kgYGWA3sOzH28nhGF5FY5zkbf1dhOlFy5tTmHJy1
rMyt74q3zdldThmL3uQqGifc9FwBSb6GjHYSDJAPZDI12m9fCdpXLbu3/b2iHmP/
zTXVJhR6NNGkWRlZdvB6ehLdZrzk0Pa9E5Ovfb6/2PaxazOgxMa9BV5uviMsVQBP
H80Id3Q++8BdrrLGANEPGH7BOv7hMEJyu3dEkUETirGrG07nGytDVKvQCpvlZ80j
q+y+Se7lDz2NbdnpZOOzBKsevlPcan6XljUXadtPyh2n9NKv018HzyD17xmXTH40
z5EQl+CcvnhL2JhCnOco130tDGt6rI7iW/OAosnJksqaSEhvCmliuZZacPAyQB8Z
ML9b4DAnFvDtE1WUKiRRtEMYxDyQcQDqqklOR+k+7+XHtJZVPWgspJkmWR/UfDPR
1HZ21o85vZdJucNsHAhvubOCbNIxdTPaBlB1l9uyW7akIDwX/3CTp34C9bRStflO
npoo+rTUGAfwRVxw7JJGjGQgt5V7awLddjemjm55EafCmAWdYKWa70nVGL097uK0
rwMVRIjfsoi7ecoVAGwK7WUoZ7iX1Tsbsy88dmGN3eNy5A52r/ntqamKxmmqHNkm
tyvkFFjDwKafbC1tOIM4f3DSLjTYmOP90YZzaZPRdQN42UCMj25hoJZLTdUWyyUk
bQxjL6j3QgFGHGXSlcIzMtl3R3IIc+8MUtjMoAY7ZJaUDHfjuZv4sC8hiI5gOuWy
U0hNYnxjRrcKT1VmgTQyLRXf5U2thc5nLCmYUzMwFQqoP89blGvFRzFE8ZatoRsf
wFf6ByTByKANw29l7eJgxuUkkm/ozP+Ff0YhVqY2zWdpObkCkFUfE+gcHMuHNoYP
ZRsIqDLdktclhoph18GcB2KWR6g14ZhgVuKD+Z1Og/o4udwbSmHTLcnmySbBVH2+
6U6iCulDwR5XUP8nNQfElYjRj5qEZPcSzLqdPyqx9hqFA8r1jt91x2O74yZ2PTJX
fhly1QC1I9wf5dlYxYn+nLzhRxHnpl78GOZiuuJGvw69gsFBCOKOpL6hX1VQ7m8v
maoRUr0F+2dpIguhSPT8qlrTi74AtRU+c5O5CdXGNSeYW2EOmLKFbI7/l0SacXaY
olPUtMPzuZVZBXwVT8HeAFiE2UdOV0eTxhrDeTZexVBnX6CmO96Go77QdQdinx+Q
oGl8yVz4ay8FeJdX5i/6TllCyICyXDNNrk1XfcoqUJxbCJWVnY+7uNdqfXrTg63v
q6MUJgrN44L+lp8t+pdK/a59NLh56ntgvY6oF3Gnl4Xl+K6gx7RjuZtgd3dp0NlQ
bF4ci3ZRr1Sko4W5MV6ey0uTbB1IFnY9NSCoyQhqIjEk8g6NCorjhs/TSG2oDrmt
UNz/sqYmt9zpnToreo5u+otTCnAeIvo6Jio7MK2MGdBa+QIdGbX/3XKElkRTEGgV
VE4NDoV7Hmzp1eDT7Z2deKpC2sza2ow7LoQIPMHwg16P7oYb4VKmRBRCVcyQwqXb
W+2V6QJA1N/ljlzP/mE/MAw/g+EjMJamAiaHFV8bo1Cox+CpkXfYMSCGZOdMP0rj
nmVamilQO73/amkDkhkqEC/2yubLry8AYNEHghgnvNIAS/SQ8q4Zmo6kYMeO4nvm
m8nq1qLIooS+q0tEi6uDqt5WWjelqBS3uet2Xat13UjT2ZMpqYrqnxQcvxcb79TD
0Eh9E3ShcS3LlyF/x/+xfS/+FxhtwDwPIR2w7BCPSgxaCeD+PHqyn4fXaZV/rJpE
ADkzQvCbk+o2Mu1coHmpp2fIMA8uBXI1DHCYvaXJGpWeNT3lMkJ0ld/Uc0s4n2iA
j/A+FanSpGAoSsmv6ttVl4joDJrkSxNVVaFLRu+ikePpSZws426W4Tl4gnRw8aqA
t3rZtnHYd6bvjVO0R2J0fDQ+sc+Y79w5otqogsTQjheqhFplxkfbYM90qSFgafeF
PegGs4v/azekclI5YD0lI7g2Psbfl+QzQPyhhSrPCsj4gyz6iZMoVI58Dn6B6iI0
sGzplLFZzLD3H83xnZHm3VFYJl5iTI+kM9F1lBRAQyLQAP/8kZMR5/ilHt/r1ONr
csTA+s5+b9ecT1CigepOG80NnBR8hYo60PB1T6r6E2aV/B9w5h2yoK1pdlxg7pSI
A7wt0IkE4INCPLIwJuPE63D8Yfc9X2Yfv1KcrKSTjaH+19AQUuuSJVDro7GzncWc
t8Z5ggPWF4ozw2hLwmQGrUceijyT/zhYlnBE++BcoU9Qen2hSBGYYayaSt9s5eza
IK+Bng5hF3Kshu3yk65fanK51lTYh3zn7sb70Umpc0XBCGkLpyB36XLtD0evTWiu
+NMk8azsB/p8ulCPbxGWKntsOaB5dZnlC4740YzMPKyAatVylUYd5ceOr8lWaKar
ozD1WA/AIJxvTtQOjlkwx16J2VUgbSV5XxCRqNcJi3eckT8Nrw2rGHQpRhhNJxjt
B489rM6mbtksw2GCc/9nXsCuK9mM1xDdrCL7BjgLOqWFhmPjpWvCecZw0oQVK8xw
52E3q0Jc4A9iQW80RVvUN9Mcj5aCnnQoyaq5r5zkLQkIl94K/yA9EEfj2EZGUMU1
SwPEce0UvM80xKph8K7RPi2PtgwVtfffTPz7YcghciwV8chGfIWDX3VlxpwxHg9S
HnO2NbtFgs3MZxPZ9EAtfRAGJeZ4nb+cWBbCEX8bUv5QFOgVwy4hMI/b/SnVm8SW
XVs8lPfH09nqbrRnVkyuyHzPeJ3cLcbhA9swwD4nKPvOOMXQ00yrAMdN6AVSpcG7
7HipRUaoYBJ5ywRULafC5fRHV/txe5iUfCghpl/gabqGm2ZjBWK5TRI8MC7emHjY
bezBhPX0LFvaipFaoLgKQy6phUimpAKCpPhflKBPIFkHmTx7xQLOGHZW/ck0sJve
jW5ejalbHvaA41l9cy+mETTtGuTaIPAwhLghURDyovpnJQG7xin/A9nLbrUEk3qL
c/KhF6n+LxdkEDITBKkTDkekRJMXV1OebaTBZSGCuZG4RSUwc0dK6jVyDcmIsXzm
kn+ntcGBvZE3xK+UJSug9sY8eTq1d/NGyHf6ovp7jCSRuhgo+9xji79bEelD3UYx
cSzs+hkR9iKCsV++KBdIFgiYnpb6B5a6LLNJ6E4C4Ph9FB8t8Hju3KlLcx2eaQlP
roC7FCA3Qz9nJ2sgnH+9yRIubZtu0UIv/AX04e97vtTAN9pj4SqN+KBnXaJoRA/2
YeDdHQu2MmoWOWK6Qem7CtMjfu7KsKpc049fiu+7moAJ/ahZ5kIEuznKIjlWznFT
2JRrC+pfw29tHUwbJUxnf4dlxTSPDpQJAMNA4yrmJmaLda0bhdxZnCY9k6vYGqd9
c9/UP6k3fLsrVNFhYxxsaVP2E0Ebm8mur7qiPj3Qa64SN8UUiy4OQC7x0O1gPurO
o5IoOglHbx7O5JTWPbFWA+KyXorODgBfeKrXNnCamGlThmM9BzLKEC41nDS2AEed
pbOd5CGKyPzdYg+NYFvQ/oiNPQOdApNgLJl12DHWt6FRW61jFhGPBe0eaFohZcjT
Mv5k7KGtWqK7iuMifIZo3ANN2DkjWPl+qMvRmmp6sw8Xg9theDGjUTWLSztmETY+
BlxYcxo/Xez1mmAG/k5xGlimtorZfE0G+/EoNtBkHt1Q3ghXn6Z/7GEwX9dxM7l0
MXlpyLCWnutxP0GXmYwuetHdtXgkCqmivh47FLLYwmQGNEzoDlGz0n1R1VNtLtfV
hEdW9Lg/oXW5b4YDWMA2i/rsB5AP/1+akYqOTlXpS/n/iYcFzyBS03znrh9hCeh9
CxQfLzsk/q2zLcvFUswWL601RsXy/ffOj4zxHJv4ESmVUy+5YEI0QHrE8gGuRZUL
plGz3hir5u3gzUvIt8XOejAFZJMA0zG7BkFHgJFTjEL80OqLPyPinXloQtP0g0y4
nbAmP9pTQMH0Ujsl1aqtmUtqnKPDiR/6we1yuYcnNRWew+/zGd96rFHA4KZtVrJ4
jnJoPA635oGzbVE8X+kYXFPHVB9P6Tjx0zerEwPYq3LGr20HTYr1oYYd+0Q70N38
0KoxpA75A7ZS6Gafs3aUNygXmopR2wnt/fXGUYrMUnO/XPHeuFvrHfvnum//Ov7e
ooVcz8FfNnY7PUh0jy8pCq4Vmsgt3USgZRoPSSAvq44M76CRwLFyw/p5Uu0MhfhI
Jx8isUQXHBLiau0a2A8Y84s5bvCKyK6v96pWnbOGJYrl54Us+hvmrLOjUg4hdBAC
tNjLOOXizrsaDwt8f47C4DoH0L2QCytOOyt024XmmJ+dHKXJTE71awNfJB1fpWAL
OTOnNH9tNNKCWI6JV6Yf2gnqbkTCTC6gv+ODnXUx2LNeypYvYcVk8QU9mss+Lf+c
Ra+Gru+0nFM8l4pzx9kq4PmKDl9fbriDCaArC5WuONo/CecafY+8nPLhCxK6Qacq
70WzGEJZ16fSHsejFXBY6jc//B2J+8+xay7Ujg3YSVvOj++pazeC3w/YRlzzrDcu
SnhBKYVKLT4pT5GhdvJwdQ6ZbOzuFqCz50nYtTJ0WTGv/MDMDXv2i9xlt2xDlkgj
dIDcaRQ9yxwrr7LdgyzCWBFCWhrxfUSrtLqYknz8d2Ox01dK6OZd1OjrRJXUNn5K
DPUl6TGJm0C+7q8sf1DdtXiNkthUDOuStUeyalJWXXj1jTKiuUmGbkuwP6XO4STE
aeX1ZXkMF88kSHHIRd+weL/KJvK7Gv3waVoV0zmJQBm6IBInnfgb1sP1SCkht7nX
a3vI+1nX5zePxXQCu33Hta7PX+Y15PdDmcw9PBrPL+tu9p+8Y2o7QsP5T3deU+8t
KwSpakRHSKI4mLVemNcrTpEQsyABhNb0PLyrcNZAQ7w3jGhRt4rLf/dnU+UDNqQf
vFuRiWMaA5P/ex8V7Jxbw7FgWa5iOkpTkhy0cMEoPUbWRmf2rvAcIAnMBNYyk583
jjmC3AIBGV8rbIjXRDN1bUNE7R506Z5cNoGhrjDyKSgx9c8KSdQixNPf07/SF5wx
bmGZFMA75qWZNL1Cj1I0mOTFU2pmV+NxBYPETEgmXaJ9a+SxduM0cNK4qUnexyPL
8c4BQ+IYumDVF+X7fjS+jcf8BLPMlr+B9FbY7O3ELkicOTerFQyqPoLiKNeQb2Vq
4kxFiORhhIhyJYFCm2DqKQ==
`pragma protect end_protected
