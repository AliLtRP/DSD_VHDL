// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:08 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
QXRXOv51u6w4yUAZXT98eIcFWVmpzVa8MH3JZiUDCYVeg8Gh2NhZBDrTcnkzw0RN
25Svm3mxTNhlOCFRAIlC5VU4B7YXKnjCqmkCo/pkgJiLAgOzTGB3mtJ2Q0iiIqos
OSOC0vObpzpd+M4pbCsg+94ZnHGF0aYrs1fw/RC+geU=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 19552)
Syvl/Z5rgZQp49EuS66e5cQ18Ukoi2TimtVA0EnSIQeCA33GZ9RQ1XC4L0nyxKht
0DhpsCPM3lGte8hZyALqYHheubYe6y28b/oMi7hB8Ls2M+MunnWWPeh4W72Ij8Kj
KCe5GjdGtZ9pGqO50/2g14HXRJB8xWyYF7WrQu3wNOEBytcVyOaMdU6YpTBmxdm2
ScCvMYrvIo+3fOwvpYS+G1awfhX+EWEynW4mzr93C+vq1pWtp4cFcdUDNDw6HoEQ
oTx3eOWU+jP60AtQbzrwQ43z2CjIFb0dku+37aWQQUDWv50yeQKgXVNPRxvxXFzw
gmKYkN+wXubM7QiCp5gKAePelBys31ighV8qMSW15SxD1OU+9JSRhnh9scXRqzio
/Au5rLqrT532hSLMfpCl3rwgTYQgCkKgOaFB7W/qlaaqALyYQ9tgICl7IC0mUIUQ
VOFESsP066P4qHygfnM4IkMRrZjBwrEn1mQkAb+RHuLreKV6EsNBEeHks2RFGoNM
2xBZyNaz16LTET8YYwHuAUauipDzsuTQg+5QZ48wIN1ds9tgPBoU2fXbsSotp3pP
ef/Pq37Z8tDJqZG3tkiKVYKkbSruycmtmN/VP17fv3N9x8sTseeokZKQ0g2gdvaF
A18cTVLBaqu1+lzJQqCVjzyZ5HyHeJ3WHONiN/qbk7DA8vaANIYDojuOx2KVTKH9
xuAFYVr5OsDV3OTts/uKEKRKswLeoqAfjEIYkO0ZipnJ/b50tuAp5pLtywsaClCi
aa2E4NBiFTqvGdj7W3pRTcxNvDsJIuC3em1YgYkfTUEwRYivd+h11yhP91c9IHxC
HIRfzZev3TU81kcfHMydCsrB5mhjGVc5SHVW3SjHSy48dBbt04clN65D8VQojG6g
FFZZdGIVeMx14k/ircsjkLU4O5E5yyLjhVCCX99jNjRmBoTleWVLsTlK4MCYLjdQ
LSoLNmNWb4Mwc9O7TguB0Ee3j0IKnI5yVDuMarg1+ZYXStRngSnkbWg4MRkd24SG
4jrEAneWuoPTp6QD8GfY6NE+rtOYkzKjxlqzmmhNuK4EpK7Z9+eyCzAR/UI/aT33
KcJfpa5hsGrVWAc1Vj03VrsIT5yylx3L7Np0gCadlKALQQEH6eIf65u2jWdEThTK
yCR2Ub8rU0XZa69iW6kkT8ruYR0oGAy1TtAilh3fFfZn69l/kvxku/uXRKeJHBUU
iHrZ0rE5N7U53cv/oBLsNotE18bsmZZphJvsOZ2JDvjw7XVmkc57xfZTt/H/4G0Q
cQh3Tgbtr8omICv5UW/WHUsSSlrEn4WsZZHTYB+T7ClAALVMvZpIcqE0VA2M3Ey7
uvGr0IkFLrdASrwQGkL+faKFB1EHD49RTjuAO6Mf39SzbX8ymbJ1S9YUlOKIsYSZ
ugeiMshgh52XRSjIc7Y/ZGyiLrJLVng5fwEhLxE+Y75urctIXMeZXX5NYPM2yCRC
wVSjUWLuWNvCMG8MrO+0mgGHLyOrDjeTCFOkZdewTF+ASOYC77VIYpBKVJP01qJr
avT3lpB22gv6sCbUyx51LHEvPszUwzrrsV4K1612FgHijR8xXM/tIV6JpIOlUZj/
kRoob+NMhjoAhKN5k3pyAGp/HdQ2QRfGIVQ6+AsXb27Q2nxKn/8lyM5AS7MUjeuQ
Tsm2RNzGu/jZ9DJ7n3WdW8p1XHUI28wpElKron5KNinqULVyzK6xkcFk5gwXiJ+j
ohF3A47BVhnhfYAPL3T3P9Ppw8G6PQl8TiJEZvL6jxiP501s5rKouip+r2kNT+oD
TNM1vF6hIEqszrOIE7vrR7BRGzhdkGNPKKyhG3oAxfKl79lwUcTaYv/0jdyoRXYS
sAryXEEs8QqBrg+eeNlqvRlNbHCtd+mxtjKjHmLETLvxBqmQSeMK//lou4bFvmOr
pkwKLanopOT2IMsRKmxHD26t7bVfBMLIsl2hrSHeMfXCy7ucl9FRGhXGhSXBX0kK
t5R8kieLbAUsF0WWvr1xlE2A5fC9e4f5+Ev4k86nGwToE3F/DGulGCuyO10UlleO
DeuDNQC6YDVn23ecqKOYmq8dQil2FIhsbRn2mscJWBGSHnhX7twAq7HJAfEQOHim
wEIJ7b8hOwama+3LEsX6h+0GqFovpAE+FbXg90nROW4U7lIyNAq+zRW++4Fbv/+s
Ly5Uzz6n1A3At6RySJGpWBcyqojgkUcwysuovwQVfZ5xj04iR765Ff7x9+LWBnKo
IUs+j/LUZCP5St9xaa8NZsmAnBs5dgZ3wzNV3n02oOzmYPaz9NPBMw6dpW2XKHd3
FtJZsZKxjN47ZcL4b091k8ur3KZ8HOOzbOl/l34A0vf+c4oWDqxVRrb2eZUMDhSz
wES6XZ7CTH68ik1qC9P1uDysoYpEBv1OMfrd9Msq5ZYAWHtwCDfjykqFcUPraoqZ
Zu4x872n3TAAZ3s50WpVz4xwq/O+43+QxMyXYc+hwS/iqvz8C3BVkAbgdPGT0LOu
GFu3luUbyA/hxBkZ6Cfu3MRkJZ+F6KdnRIwywoGP78sfmNr8vAGUna99VpiiQSwJ
/343wFkYKwF0aYHalex9o161q9EJnmh00RfB2Vo44LE7wL8ltwP2GZQqgD6Vt/fH
5TJWe3jYuM1oTWsQ9mQI6MAr6CqSDkvCf6uDvcObBCMTLIcO6Kq+mEy42lysx2Sq
qTH5UmXrXpgJAOmnDNFdpfQJjgvZkuEaeln9w7bEP+stZXfGMnDTsunJbsrMclM5
0dP73d+18iskKx8xRP5G0dzAVfbpWVWKiB8obOvNDD0W3ZxYjmIa5JCARiuoHSV3
aIwFpcW8KlC3jIHUJWGqd/vXSrKyMLvznkx1qzAfTGlyvxgTUQLNqd4/rR0Hw9Q1
RhZxGYJHwHr027jyZtykCdSZ7+w7igUexwwcZ9EKCdGpoyz53/33dqJpdtHzA8lU
YM9j38BEOMVCEx05DyIh3/X1wSxhIv9uUbc7Kk6ko61ZBTQRrdT8HAC4ibGgg2CH
d/kA4/UXPfxk/FjsR/bJch8fwf3tRuRazq7DJt/obO80ZIkuMvuo4AZp+ovIB7t4
Yyc13vhYzLGb3XHb6Gg0zb0mDTVc5B0Zrub9dM74DjywE9d50Cm+3yWdAQUrbssS
hANhUqmA3RkSNkJ/xkMCjaaPycBS5DorqwW8qTCbUVJDyTZw0yILQ5WurE2L6xNa
7QbJpFIRCI+pC6EPFAvmwV9oyz3CcHTtcWcFJJylz/bW+s7sJDmdYW8iQOaetsZP
WKsoGKATamVCTPoIoTPXCZxE0LhEVDBruR5Bq+nnC9r+QAOqgEdrCQQW3voWr14F
1cmemT14olNjTaD2ikRgrVMVC+6k4LMExi3PrX6JIB+KKrrcx7EyeLh3Ayi6wCFk
j9XedP6JtRn7Rl1QaFv/qjnVYwInxlGVx/Fmlx6x4cIrAZtVy8kamfWi5HPOgwLi
aFA03x7oq2kHC94jDv5EOn/oC4bkcsFDXm6ijyky3CblQDhPAVjhtC43QCys+tZx
CNS/KX4BR5f6L5taxieQlsj0Yv6suRsh2Wnx5fRnqH3UNcEqW7/FTMFa+5fPaO45
0GdGCJXRV3+OoSOBWPiJRQIVmN5deqYHRy7aaZiuIIvbHlFsy56RSY38f2vIoCcR
Iuq+Uuwj1RgqvbEzh0N8DTCtVRJnLbcXcEYEwy+UQQcR2IBJ69sjZkgwULl7yPro
ZBXYNTGHqZ+yVbvydmRE8lwvRTpV1cyOoNDypB62AQWlHRjnSC3iB+0+kE2yyKiA
OoJqFk1Tt0QSXjlzRGpsOg2sR7ZDZBOuA/8rUZ/O7cUP+EtdKjcYs9QaxSHRRgjx
CGk22tYJxvZ7OVrIdkKkjvMOOQQc7utMm/aW0R6XLvsq2SfSChVCxiKBDfQ2S5c5
DaJnYz2iJf3pm5/FJ2uEI5agbObDrKTq5CwnQRlW/8sRfeHqq5Eyfto6LLsjdQ+b
g69Dly9PmF/qgWYy9Tv7Ggga2js2zA6mp7L+th2h11QaZjV8T/fGFhEwqt6+ncYB
jUlS5KB3bnk6RZCYfxibMn3EaoW1QSGOozZdm7jQJ1z3dOhywzrajyxQJIWmRgQ9
9HEW/Y0VVE3N+GiyU1wyfi3Z3VCRnMhbqn4AkY+62JVyVPrT3rLHfakSgHPmJO/7
YH/rj/YGCQZ+fQWVpgj5ljRnrZPIFUNKo7lDrVIyl8QJaV3+XYuNyjoUifd5H5Sg
yQkEINWq8nSJHAGejLb6r353mQ3QDPzRENP1s942nIAmchDIeoEL7zhJfbwckd1q
WMxarQCUHndegl4dZ6m7DLskh4hJ9LAPxCvDpox91eY1Rhi3+idk97UqU69gsa1Z
6Aozhd6vFghR/ePfdtgQXmdkKmgOHZZ+O9zj/KNmI/bQX0bo/OJD2o0iwshCnRbd
EievMB50GArZiMt8iU+zcXHHzBLUJL504UuQm1fb9+96CSgzl4jOR+ML1ixQ+c9f
5v/oRNvS7B3F6RL6s3zwstz+h3SNeFEdncoU27Kavq8OyU4CmYxQkQLQjZ+6BZcl
fPX3KYSTiwYPMxJpP751yY9mlLDntYAvn4F81JyhMW76d3l5xrwmXxcUKLzKUpda
AnhekbFcSJzrBB3Eot1VEbAy23dHx1QlWQOK/SpuNbSXe8vMGBODo4HRX9GSm6AF
HweB9M1nLBIBtmtTK74uv/h680nf1SY1R0s8vs0L/vz45OGcupLGq0kygQSTUjoz
7IBV4YQcIBSigrh41l96gcokK7VoU21MfvrxfB+hJ1RkLUz+SXADYp/SAeBM1DwF
CMps5kySy5k5bnIGtfgtRd6QeWjgZU0eMq8FAihjJZ8ql0rSiBTibmS3ukJiYieR
PWOfugh+fUAtNv+Y6kLvdSgo+ZOXLDhed29D5Qd10OSg0/vDYwpO/kvsl5zZYByH
zbO1VbqEumDDPjYJJQe7RjuULxuHSbH+I7ULNfEjIszOGYJUFkLYqGxIfTr0ZJf1
uk4Y98ke211PcVtkIFyPA2sVEXlbv7/2+4IPIzKkeJOk8Ya8wjv96QZAP+mkQSvs
n5T5Npr/ffhr13NezJFm/Im6AmC8wX+Kz11daQHBSUZvAGWS/VBe5tGZW42T7Xj9
oEL2DFspIToJp7idTeNDkx+IVVZnArznvVw8Wpp+fySgYCdsmGgsmlY5+9L4tpQP
mj0vsz0zeJQqtpRvh7YyDA7CfTdR7acApr0j/2hjzXVEA82l5zHJvtVbeUJpaOU3
PgImWyY0HNxj9Mp2nYL0WWePjG1lG/iLO+HDEEvv9UTNdITU6Mtbhiepx96UANmp
QarkobHpb4MFzeG8NqPeASMBzhCe1L9dB5JgYkOxutW0bPNZ/9UGOxKESMq+HVG6
QKD09W+KriR1sUyb203ej7MFJW+Ag1O2aYp2hI0lWZnoZRgfy+q0pqPY3KEyhhKW
/nkrAFq3VKPsLENAel4LbCt9E7sWglyfy6CP1EMP51RgESTj4rdtDEnxApPXfC7t
lJQTaVouF67L1GrsfomA9C4yVHIXHZ0Gwb4g9HDrvCs+sr22r3+3D/0YrjFGiUSs
drDapNdo20Jty0wmkJb3DFvozPQTWg24fplyc/6JAjVnjkmI5S/nma2BCL5Sl4Td
0canc1saFrbX6Jo3v+oxlVdNjwk/yQE3QRsA4nnAsEEjB+8FI15SwH/USH1rrspQ
0Nhr6wKuvo7/yU/F5q364Wf+zvFSuUbufq8/iijezMAxtNSGqf4/soinyKVMTr/j
/bfhYLxABPNdpMOW73kr8xxiC9La1DOzkwmSxnTDRhzOwYwpbTebrLSPM8aCyzUk
FbaPN6OeO4j3uCrUoFJ+Qx1m33JaYw2Gv/mSFE/cYah0aCsYcGZCll0Q1s4IKoG2
/buLQpQcHDJgfj0HQGyCZbSdaQooVsUpaks97JEoBW8cQ/GnLamjZJkkbliIBMNc
G49VkdD5JZoOAnMx/BRFTzYTZVymWO6xL1w2GvaT1Rl9uIcNgOSBllK74XCdNB+h
0gHrY06qgQQDY7NigwHjDeWP8ubfuEEmbZ6Ia4dxF+DedgCyePXhhsJS0WcicgXZ
7rcEk7kxlSnl1Mi1KB9ThWPmT4sbPNdpIjz0U1FFFnMDpfDK6U2mWdLvA4R7rch4
wQiPUiJbeo4m9IrjIcf5LiudtazM17OW8J6fB+mdB6iHQu0x8iJ8iCM3q9+Kbab2
SW8BBAWk8XyL2ff4XXpPtiGE5E4n1TuiXXZoa4UgFMgTWSSTIL4vm8ZYXEIvZ1fa
32ubYqpkCpidPV0MOJYqIa+G8ed/iTc/GHAcgm98+YEukLbO67XeMseZ0rMH43nT
3XXDEm+lRDe4E9i95yYT2YfjUsgjcUyLoz3woE8lT39j7ZMFU6IY4k6jPN7/w9DY
aHEEHUJRXVsT6WpT/rdGfaV1fyO/naS/o4LzvSkv1rcVUr6SanTkratpkJQFRsPi
98GBg8XaiL7Sf4ISuuufB7LneCfiouycl9exfjgNaHLgsYzgp3IWR1xnqvcAFZu2
3p7+aSLuRPr8qi30iDivwqBfLx+LNAYeZLeWi7lYZbMZOkcNuAZ6HUCX8lPaF8v8
/ybdiTO+/2/rr6RqKpsCT3RYpX9CF+oTE5HnG9zwCN25IrA6WwoW5BJpL7bpeT1t
mlIoz+h6NtpzYARuGY3a6kmaYjgoOZMB4fFacNLU64go2+VAhXs6eyUwpVhNlal6
zEl7zf4dcIJcr5sAsGvnKIXes++Rp696Pw50LQaA7tWRg8yBYNs4qpskHtLLDz0B
5oiwzCTEcXfZe8zpJHo6BIJU8Ly3/UrvNmTgrmZgLNsXcMwgBZzmKxTbghAk9oGj
zNAN1ZeI6UmfvQukdr78AieCZ+I6yWYAGiFSEFv7Iu8xFpIMThSaodOQbXywDjJI
ce8f7Kt2sSvfT00zz40tNZRknaW2s8/FpK/2Ich3B29KvbxtNlgFTJ1JiKTV3yL7
hK8bnzH1VO+KBk3Fn2HolmGwVNct8SUIgY44nd9aTFAK9I+sLFAK8PRtKWZcmf/x
lmwK5/nj+uAbIb2AXFcPHYaCblhkYB+ib86CJZJYmNKMOG8/JU9MO1rk2ukgJWBe
6sD6+Vxguqx1ofwjVFG74RLNbMtO3z4iELK8U98S74/BiZEoh1QYvWnkDnVwG7GH
MqwThIZ4S60uflQkrpqqNNHfelihgWpD2GzbleCNttnVI9nFELSgBiDvCF8eEkZM
2bJNkwCZiow0f3/6VNAf6s1YsPUaGrmuSpE+hGWp6kihobcFeqESLgzcTiRoK5WV
tawL6htFbhDJeU4VxWb7LwRFGvKjdCvz+mCgx7kJ0Ir9ygrB6KxfEj8VUbHPCdK1
PumQZIPzEG6xtB9Eo2l/7eIufhSlDxteeypzP7YOaB5CW7HGwS/miHWy6taib83X
s+azCf6tGDJE+QxQkSAQiwiA8RduYyp1aXw4eDVRQLi0onoHVZcFBGi/gQolozoG
z5PDIGBBwkBfhQ5E9lyydwhzm5eP5tc8uF3JK0cnMH4Qi2TeHYVFXiPEQTc1mgoH
G1DRwnPDkm/eAw00/QztQJkp0rcortC8O63zTPB1rXWIiem6Vqko7xf55HzsME+W
pWFiwh8QcgiKb64hId2jN4gTNdLZKsZ4NY/zhnL82S2BSXPsSd666KySe1KGqCfl
2r6ios6dwGSCF17PrJJru0a/AdMItG9PWspzvHPwIgCnR7EDqLCXXRQaTb4e6gDs
PoQ4fit5QMN6to2wqHn9ZmEBB1HMI16mzvd9FyywfCzGg5wlGbAGZdybzlyD/oLI
h+SriV5NIRgFBEoZT1SwCSQPZAqnSf6hYb6i+K4pNCdmuugx/LfNMgrqmzQHdum+
ATk5cwgc8fwK2W6i86g2dAt+q+Y65kWkQZwmnl5Te1oSkHHN07Z9UXhOuce0aBUJ
6S2npneQXddx54hVxFYN9r9kFefc52+yUeogcdz6VKQOXJBH1f8Iekjp2sZ1QSf4
3kvc/ZKJr4ywKjhLaKu8ccqATAHH9rKzounFuBEyqKDq0AucLyitB+p1NykeFDAm
Evi26VrRgbqYmwdnVwj+Af73mUqLpGOgxqY5UFQx813Iu8Hl5E4VeB2UaLkOeNPX
adDcdeWLIWFCRF4MDMn3M/BY1nkSBPgk7yOdyL7Q/qp+9HKMQtrK5bd3onHsCofn
70lrGVuHcQa9fbcxCNMzB7rNenmBwf30Sdv4SKHhOfjublWC/dwZsAgl5s8E5dNF
2YW1zO5bw0dZUZBO8quPg8GwCp1Udw6a7Fr8EwPr9hpWcwYVWw9boejZFp6KrpkC
IBkaQ6uSRSrrnDS4h/pV7adNU+WMpN9RsU2quWDMVyksVlK7fiv7Umhxv3mtM72J
WPq45BeOl1VKMKUIuX8ZmbGBEVlb4zoRCKDptKm3vPTnVeMtd1IGM5b+D8tmPcDP
ni2fL3DzKRdbc5iJnP2MOIx1H6vTDl6kV632liVV2u2K9Oo+Z3XAAGC2CMwch1Rt
Ugkt8iiDLxGZtfIjWPRleJyrkOqjz1Bt4K+IwwECHoKNauFzcw9YbkFfOT+wfD9o
z5yCm8i3+fFwnG7+mGi4EQ1oxcS422hceEB4BeketICTKxTUxbsI1Xj0foGckzCY
skumAFzyxofWhvalk7ih1i/sANaqewaAz/9HgvCnNNGCqgTwdXPgk1xT665e3mBq
oGJi/tSK3sP0m2eCZM1iYRaf1Q3rdKMk3SkSpUmYOn8iVbRfjhRyHYLr5jNxUA1l
s1L83XpPVXhmqosdDtoL1q5nK5sW4EYPwUP7qceo+6RycqggGFIrpbssZvSbchJp
2FWJM4PbAo6dMf29cjaC6EHuh/dWjw1WFkwPcoeoDFAr1OIby4b5VPhdSf5Bo2Na
11JGHsJmyt1OrPAwD926NJIXCZVA9M+lxc5eEkNDFjDTo1Jl/euiJ0q56low2sF7
cnTurJKhpv1VLO/d8kpwWJikQrHG/Qk1yw30EJxiimmp2mo4+CooH8Cjasfiboon
LfgcUUO/e4zKfJSjzpS5dZoFq8Vnhexe4t1lYMzvbkPEsIhOKb71AuLbSGQdoVTO
/GCM9shDdlnmmbcdqeQFIJ2aebL8Am9oppZl3IjCeSusE0ALpHicyT9HfSxAgBVY
yP9R4fGBlHQgWIQC1+2bK9oM8k9aSux5ABhTIO2H8B/foBXEPEsZM99UQe4SY8xc
tUz8aLJSI19gcYu0CfZTD7eXwhfG7dQCG8QbJRV9PY+zan3kvAlQDxjmixymPMM+
Mbvm8GFY+1d+P4DQLNpVF3TW3WEoqHH54nE4zLsIxF0DTZHct/kSt9HG0gSUfpau
37sx5F8TsGmG2SY00WpTfCH6AvznPGXznKoho+YWkHGH2vT2CWcmQuKSH1mwQPsI
CfMICk5mZ1q+ktfIgzWvcu9pJl9T8S+3ZZfJgoxdOw7j8mO9Nmipbg5Euo3E4x6Y
0AVZsqSXildZo1T0edV+PjYu76ybsNQrcpiu3nCJx3POekC5KZRoiZhdiKR1nd7m
72AAa5VgrsKghWjiOjejppntthZI142WqhNEA88c8valJ/U8I7l231LuRJrcd561
qVE0Rtz9PX4g7Gk2s8HX8wgzpiRjmwBVovohsyp93ZNUnICaF2PxVgRbOzR+pQtp
kBxNf3BJ9HaTUvbNMrR7ecsIlpMkgsdVIQ8k5mQCFxmLEOpsT21GdRIeD1pjoE3U
AlwOgvHqVxAyxNuGWQaLxbxq1IsVybvcTglnOROhC6oYzQwn0yAS9i3xzaLFCxrc
51DC9LqvHQBNBn6M5qKzsRuI5X79rIJlPeTFj3hKptlRvDuC5uiC2FW8YI/oKCRf
BX+kIoCZVa9qbIVi0p31NxSLC2kYsFRzkUpE08N/TCXXV2flogRF0Ytd8h8aLvjA
+sEhvg2PWvAWt9Y8BgJFF3MFC00j/OXcGA7DITK/eV8X2pTL4mLlpOEG5U0uEDYL
8ThO6P4Nt6fY72dnA7XtOg5KgK2M8hbwzWXJZYShR4LETrVicNB+TEW+wywasMoy
Zzi5p/TuJgr+GSV6ANtf4WPQ7J1F2bsUtDFFSAUrqYyw1v/qjX33jxwfozm0z4/s
dqYuRqIsARm/e4UWAX2jU29f1Uv+xtPfFOHxRgzGVLjQ+/Twkk30+PIATNeyslH4
VNuxpdCq9tQVgSS4bzAXKziWMIQECr9KUZF8llGyIkBTAjPqwi5bxQUKO4AqLgw8
iqqeqjnGbCy9Se6ACNpjtMGQdS1Znh+HIbaCyyJ82RqUNcWxNS980csbBlAGRZix
k0drLWrOlfI+ZhGiw3vhRf9xUmnL1MO7En/vp/16UhCyu72Xrsbo8bFI0fsB/Rbq
aQD2+X0uYq0WHuC+FlTJOAqDFhpBJZD7FFqmOs3Cs/UCI7FqMaUGxsCDxKqeZmMW
D9i6c8LBmn4KlBS6nxq69f0Rq0Tv39g5p40gBAnSav0KSdd/4HBgEuQe2/S53xcg
ua+STRlzi/YIPhJwRAoCxA3pDHkj1whLtgt55Bre3yb7lx21SkKbCJzr4ooc8JAB
6ek3Pw+pJlCOyJ4pq5r4Z9Y7Tvop7TPGCMcvcbAczLEPSg4G57mD9umhkgbki2Bd
mMaLKKkXFNkhAZtT+h2FOdCaNmzu4s6QVZ+9gflH+hCJL3ATqiT4095TTj6lNtAv
bp3KzqvChXAWO+esDX7oY0AonYrwQrd0hg1qsXMY8QfLamUrq9VqL+j8+Ly5B9d0
AyUngl8xz9DK5x1y/owC3J4C0qO68wdvmoUsuU/fSn1RO/k0FCpSNjA9dx9Vpn7S
BZzlkpCPOwn7peKGB6sKPD4mO2zbxP/EwgpDEiR0govJMcNktndjRYXObzWni+Fw
afiN3r9gmO3OvflQfFAAxiBZJZlE2D/M/Im7Mb2ddQ63HjhZ/lKYglIbGyAHCNW8
gesjrK9eBlmhmdjTTaRiM3sJdiPjcVMtGLGzDlrf09WqhFzKYXZjDceir0PoRmd9
L+LUSpnzLcMa2sjKry24vHb6av9Godo55mYBQPYqMOnSLDcc7U8qU7VcWMygiTku
o5j97+XGTA7ZPigQXWagEq4U40zXvDXnZe7I2xhxyoZWRyfC+gQroesMSCsKbRlR
kec9UwWVw0PZUleOYVCL52EU+eajeU5TWNYh2lRAqp5X65A3ieudGVBW3qTAdTbG
ueKRrjc1F5hhQY8jkAdwFLG/E4+njD2D9jDo8fSwed3l72e1VHhuUD4Ccm1SWTuE
5zvYY6SHsCqRXFgcfeuAIESX0qluDxp+jHB/2TQBJbrKmK2MQT7Hmz/clsPwDzQT
D5Nfjehh2KQoNrgA2uda0Ji9GiGvoXDDSP/LxVLPaEo86yif4ZAp4NoT+gaFQl2N
fGfLtuqGZAM8PnJrIUf3AQO+iEsjKzuzbIluQv/J3llSU9fY0YvTcm6BXFp+xVoH
Gvl1XiIl+OkYrHjNTeKXmdK+pyaq6a6hEiqeZxUFiBhMT+6b0SnZBsPuNT4hTEBY
9VeDYvnX4ViRaepjoaLRsD1FFJMIbLre1IcLKeVU0Sy0BKwZ53mg4iBTzYq2CBdO
AjQUO76A70g5w4ivrj+UaPlooNXkNoKpbHzWI+fYSKWfNvHG7fnj/eltns/Xis9l
X2+ovSdmU41Fy+fU3nnlbnMHaqJCU4PRshgGt1xgGIbPSKGSL5kY5jHrcNgb7lHJ
3l63bXdF7fdSTh+CHWKoeHFhsTHbN13028MPH1gtkDOOC9PEtWePkCy6BYRP5SHn
8secZC3NAc5g9slScGjHNkCjdUbIBWW+XkTFLjSfCXBEDMw1ypaoVNFtx64GmXNT
zvdWUHj7T/7Z/OV5ZNqi8qxwDlHKakaxcDovr5sNTrEqoRrzT+zxsrJNRCohiao5
VemNIGKQF6mtY9W7aqxrVwRW94xDbQBgQjQp0zJt8YMY5vkHrBJ3qqoRAPG7rp41
OOVdOT5qGKwGy4jxYT0hoIcqrjTphvX0/9aCftP47Jbne9EspcCDVMDsUqw4Gfao
cFuikESoFmlOSSNdVcP6FJMRALIkn+E4TtQ6k5h3vwwd4Hw4Sv5dBPasJLXppmhm
f7YWADemWZuq+wvZf56rVtIK6AVxswvkKh6siwqUPJfgHFBrWFDBDr11hTs8pcos
jUAKIoesUHx9el/ojmlTw7jaaOqY7v1Kt5uddIuQgtI+cb3Kym80ra0OW+GSbbhx
mYY6MFcwfBI46xyjSNADXS3BwCiH7kIHFat1AAqUAl8lI8c8KlfEAJ90aW8CE6wL
Rss4MIAO4KuHc2Dngo+hVAKWixDpnyixXs1hHh+3EJLcEgeXKnC7lJ51GKhloqI+
7ff3vL+HJCZpfTIkqiK0V7GylD9s6QIf9V5h64nwg/DmuWP6HBYJQWolsXp3OfeC
4NcCFn6GVjLlm9VccOaKWX/TeppUM06xxyZeVrzZsRBYda112x7452PKl31hxprr
Baisjv38XncgcDVdWTK2DBPEG7tVqgW1VRnFNh5rkmroROKD4yeefM6uBsKPGNHW
3nW+o4WCdMx1QCq3bPZj82BhJllJrgtGgC2eAKONRrmgIFmazp12s6w61k8bM5Be
YIUjY3xF2XhCuZboJq+QXn8u9BZ6DeCufRj00kxN+LW0m+FxUXQ1b036Cf9IpKwb
7Z3xIgRVFSwhi0NKZf1Af5gbfR3i2WSN2D62+38K2N4tRtn4NYh1dPpXZvxbJ32m
qz/vWCcxC2AFhZfTHTSQdB2DIkhZSgtjoNlxP5tC/sGJSgTuCGJqGEzsrrM7C/IF
/VSB+M9HdtjlOmYakapstFRnaOjPZpzCdCOvKviSRqaJaQ6xXTBPjc8yiss1MXOI
P282Z61zILNkoPH2vxiM9/fojiSpH73iIc0WepxXWZLgY+4oW2Gm29WZKHMb8wR0
Wmn+HmO/LKk6PIpMTKvfp9gR5Zg0/qcYrfH1MSS+64pHk812fUsFjpoAKI8BhlHQ
OqUXB52twuAwBpQaWvFjqA19mHherHNplXCtwbDztBdZcZHIIIFfWVyRrAuneVZi
LGOUjjWeG63MG8MGzR/RYP9zEfBx52ovAelEOuBH4kByxHhVqHsPtDQwtVv8J9sC
NXndo2F+UGmWaemuD/tiMo9gYTc4QH6Rv9j6UBYfe/c7isqNFLRaRcFhpgiPUvTx
txnGJyjBmzmFnH6E1ilLrU/zRbusN+XNtnhsW0DGXgTWdMnJM09Nl+USqbJPYtLK
j1Vazq5gUoBombNuuivObru8Rwqafy21wtn2YLyvmyFiaFApGE/OgLQ+ztrcawW2
u8dNS/E1aOlakpEjvGqQMC3JhSvMhkK8SzDze2IjTtuTCM5OwQXdUB1s49U5SQz7
hO2eZ7/Vi4QwYnSBfVBroPuEKTXS08uX+KZUErTCNV3WSCFCxGq75aQzh+RnNN08
1wP0lrOy5x5hJIOK24xampKUr/7pFHsa746kqbxtv9qRtlXX+9ZtYxRVWS2vRsu0
/XWA1ItGjUs9BkwFR7s4cRffPGByDugNQLUQhsI/mCgoGkH2leNN9YImXAD7ldiM
P6ZewyYyCEzpAtGkjHqQIjYqllFZulNPcxnhU4xjfAnESyA60gIjUk2s1M1cQ3QE
/z/O93fwQvnKhJ1lEfajjiTq42UDcIegBCBWo5z7Q1urGybe26WgqEQJ1PdsyDCG
v/T/FKZ6f2k+yaxCFz0Nzh82QhyJkLfHhtoThRhFvpRN0x6Oqlq2uUf5f4Lt6ZHw
9nbqLxM1lhPJSYPis6MWHYXxjILyHel3a/hjtfL75sfSXTLg2EIqASi4jymFjY0k
A85ApQQfP2AJr998SXZZymKBTt48GVkC7Ti3Vz3hSeY3RQGxm206ofTaNkTLf0xZ
D69x5Er8lvN3of5a4AKj1/AFvpFA7SSr2gU7jBYPcJF25uSt1WwILowJs7f08MIa
WrKcovQ18hLb55rxJ12dskhdQhP3XnR7aoghVylC5NWZTSujYEYyjLmeefuTZJlC
PQOTRGosbPRFmU5hUXv/s0dE/2aSmHAybvqqNvkNbd/1ZqMtS64SV78HBhJXfXhV
hBTtIuLvQMuDLws3xs85OJt1tJbT7EX6QJHA9TDqyMcjdQrpIA8dX9uuL9v47f7B
htzSdyH7p1vuQ0hdQCGRthy5lYQSO35671cwZ7UdZ8HDhbG97iRL89h3bJOLhGfG
UMmXwtIUxT40pE9+PMPEL8oCmsj2aQPSdyVcP3gENRavlat913I80fDCm1LV8MAb
yx1BUoDUdtLck5cekROt5Fc1HXMie4COfCL2w3ullzD8VnxhsRujVRrQeVTMcZ1Q
IO4iIc3aCGyL+dYcqRfi3/1AzkJSc95Gmow031j/WvSJ+caqLoN4Bd7pkGQkxjmW
R2Th7zEcAohXSgGYS2Qxc1CdX+oMV6yCmPKCNKxFfQP3dDaQv8wzPhH/N+eHxg6m
NCSfThr7mdAbPjpqIq3N7b54hzLGXQJY/dBmZ6XR0VJiHCtP4jzg1NYOTnRXpvUh
QT6N8dGaUiTNIeI7DSYIIOP3yZzY0t7CwllPtupcpW7zDpjvWVp5MKt5aY18eTy5
0kRi9QoI8F0nO9NYM2Gb8A42VKNO43Llpqch2ml+kN0xO7aRg2ErzUPhvk6g0Aec
jlbI2MyVlzM7KBpNcAeLFSrYvzkmN4w6EkDAkOHBJkOXUtitcdMpdj/ckGOoYYRe
KDoyOx9Cg9YHsf0IJ+Dw1RfMZkmdu7VhGie1uxbwN6DLM+zAn4jjsr9e3xLLBUmh
1cl8fRuUm8YMnRWABGlPwIEFYsfLaB2gKXHU1xdVc8WC6uAvFL/wu0f5DGLQC3SA
3fPOSvu4s4bGM864iwrUUNdiMpxUiKTn3wKUSvyOKeuHL8YikXLXaDtnZUYcNE/+
TNcnhiKu4PjEC7FhW6xbPClazSrvn8S7oE8+ktyAvZc5dtpzRqK4eQOv+OlfXvFF
Jz1ULXNtWbTPNfQS9aGymW92PzCjrWuAo82c4N+7KTJ9Y9Myjgo9GadZf91Fgzxj
s2Hpis2mpaap5p4y+Bo4idp87yThUx5enruDu9b74gvh13M+UovBsY/TSRXtjoVr
ogonkKvjxDOIyCz2UmJyww46fEfTXqAlo+dyjcn2rTHX6kEhuVaRcVoRXVyYKpSf
3CMoniJTbMMBBmK3ZLF8yUVu9APtlbUABcvZhvgBuBLu6iIFdxFI5HF/wUXAGfi7
aK4TClOXD1AYXCNmH7ifned7anqdo6aaFhSCAMOSX35T3akmEwbL/sKFhXc9qSx4
ff2pr0wHAOdMHzvNOpnng2Hefpj5QwgPQDlzm0j9sD48jx+cqx6AAxxTwWCVQ2Ei
/WLkDqNl8qgjm1sTdxLX7nj4sFR7OG+Ls900MLdZuPIzUmIOZOccawtJfQUXWOM5
Nyq4wDCkKcBhtsaDjX5AZ7bQTundMGDVI1pVqle3wg5c69FbkPjUqdggb9Px9EU8
85EUksMaq11dijEKBgz/MUWNbgdgM3/67SVksX67cYTTfGJcHKVdMDWUFwsSR20t
wxB53s5lPtr+iKVW/3zjBXeDRoOy031KubatdK/B1guz4W1BsONLO3x0iD3VrfxZ
5yQLR0x3zudFLoe/EsYzyzMYNDWepjAgHS5d4A50guJvzah+qh0LQ34Ucz5mcTkw
GtDku48W6Urylv2MqUizLVK03300SnhTZz4RhpDTxfgMO8pEliM1BdE4dzWEZ4/l
G0RsbKz752sAJjH/aEIhspHQEI4S4E0VWha7fGfcS3cBK7wgU6YhE03MlBfLIu4h
sTo8abVfbM+CKaznN0KgRdhimC+r+gMlR7jYpMjoDudNnMY2emM38j0l8wsIb45J
tNpA8kIaHpfOykPLYvTfGEJYl+UoK11PwNgMIvMgFhLJEMFmhdxlA+d5B1qVSWIb
CW5sbL3rtdhroeEMezX36iyee7QYVMtQBknRLUPmQYZrGy/1ynwC3QGEYce0f6Tc
7C1LM+eNDO5Geo+LThYKP1WLXI5h/BMSj8AKwmYeTNcN0kiQ4y9kcrxDUIOkrkSt
RSvvTN695XFQue1OWECegRKYcrPxrl4K7A+ZLcGQkUOopiRm8fuGQq1c4ZeEDbLt
7w/pe+SGah87fCbLaUAnC2kfuYpMNGJc144P2wEbWSbRlHqqko7vAPoHVc3XUdCs
a4ftHNy+KmqLfJ1jjpfyJil5DkjQzon8rJl57UqrPJjhn2NTCg8nuRwlJYcFe5oM
XwdhuONt6EXFYr6ZOHhnMIG3FJot2dkwkP0hKhxEmsTYete5afVzHNXvjFntkSLq
LrVuFheg8jmUg/QnxffnngyPwiqcazfQx6PeDanWGgLkLcD68S29twg2wVlai+0F
529ueP/Kv3wwi4toxyUQ5B3xNnKgW/vA/3XDcqakPVFubpbaYgEwoAf5pcHM30Ub
dsFPhUN2qie054NenfdIuLrIXxL5Rgytq147pXssKC6f/Gc2Focq56s2ukwx+scH
vRfxO5MryrgIlonO5uy7QnivzmeWIjhaSI4KHv1+wufypm6YpDFCmRvyGKWGrx7J
k3UxHtVqjJIvaCaJgNDew6E97kR4pR9ThIEQWaFIL9Zgnfd8MHMRFuTBCmWwqAFG
zoAuv+Lfm+bYmjIZgzAlvByozzbs9DE1cXaEmVaIurK1z0pDI+Ga89/pcPhwnOOE
3EHTKy45Ysa8K1K/qwRRXkw7QFHbdPVUPX5LMRBn0MupNC7ZrG0GtKlmLSgeQEmo
fCHW5WECLVKbv6XNjaodSWfBHlmmtONPE5wo/bno5xlrMK1hSFuvqA2FBhAmp6nZ
2aKO3lU3Dbs52fnVrriO/CIyZ0XTqtFKKkNkZPecRuDKanRfteo0bDVyEvXcM7+q
il7U/mF/3dPrm0Q0JXjZno5cZa1tJmYWWGVxUGVRkJEkj45MamimwaX1r/eb9SGZ
OXM7XWWBLSaXthsoBj9cCa7CIgocaw3XOL/NfGItG1dlqO+tdhUuA4Z2p0dC2MEX
5CT3EXn1vFDmK81S1xyBpFsg1n8/HtgRPUmX4mq8nPs/VrK4+a8fqNsWfpY/XMdI
arJi0mU5c1YHZ/joDnbLCPHzgqpO8B9nxxaE05JBqOJrEQgIZopzVUyFS38Hg+p9
7+xN+ylqoalI1u98y8LJ9odF17kxp/rLc6O5eA8gaqADuLyHFXYB44VdFVarWSFa
QPvAOtBARvTnDyFCWT0c+dLJfWHndZwNjgER6xkMYod9iAbEvepjikxwU9n3fdAV
a0GXYry7DlsANCkyB1NBt1G2bPIzefrqB3QFo5Xa00CI53R5AKXqn+TnJT0OKW2f
NhkLn87hcI0rON1b75gDNQjkvaBLQflyhjDSIvdK7YDsxEcXOzAPlqs9b6+Z/SZ6
Uw/J+X+qUwQB/NfVDPUaQKlxt9peK7z/TU3dBaJNrs0bEw92MHE0ZI3FhDtrNiZ6
OBLaLQfjScbS4sSc9HYaeDkgt50OpuzNJqFELgcxzo+UfQmwSTfhIaX4WKZHQqWu
epEL/tdOoSpapFz//8XiIDk8z6QvloaD3T1cWGq5EUP2Bft5O+o5PxEprSVBLyNA
gfA3las+AkwpENkrNyukQ40/Uh4d0XH5wFjpvGtGyLJNYgXZ8fsDQd+XHp7Wowc9
v7AnF5FBr2WbLpTvlS0uwqSsfSOtQ1xg6kRzazExSO9fEBK8ZHPZj3+y+CBXEnYh
18tlaQ4vF8wJJL5vN+Ne5G5h7EWiuWmA7UFrViFfB8fcX+5v9Dr698YhZl0v7uvn
8HwJZPgbXSYSjlDf7UahMULOborP5wRPVjpCDfbRjcQ415/0AsXMrQ7X+EwV76qS
E19xxWEj5q99oRyQh6pep7o2eoe0XZfhArj/m8YEcbPLbp7XSNbtELmT6JM3ifYm
b9qQtPFb0DFDppR4I7XR/T8301vu1Vda/FBzJZF6xau2n+g3DEgG+8wi0sp4A6GW
hyLMaVhWh0mFrdBfQQxQhrM8pfluGH7q5Km7YP4obxr1+fd+ehkERA1alj5b7teU
qdil2WgsjRM+n5ujJ15aS9OmpZjUjxgB6voBQFA8YkYLY0oyRH0rwuXK0PibgI8O
vlcPcmf4ANBGm+EDy2psQcl/YNA91UVFxGyFhMXHNX+KJDErWN12vNNoRZ5o4Cm6
q4O7vO3BT/QQ6kYBfsUi043auXNKaRbfdP9ajWiqC5EuXnFZkbgjV2v9YSXRA/5A
m1PTzJ1R3tjj5QqNFUMhdYz50HWG3N5N3gqsyqGMmC/rZCEfXMFDjQeXPOvzxQW2
j0uSOHRDqD0lmM9p4OWj0/5Pl9fbmOGroEiexr3QHDTmNEvUig/WP0ktpejA1R5r
7F322S3Mr7Rn3O7SvcPs9DuPLNxsajGOOspCiIJ3Ezue7bJsRwCLcexcnVD0JMDe
Y/jTybKISVRUjX0VQt1pyDlO/ZwPWpNMe6YIxmzGXSCMz79urJqAfpBl+Hp+66t8
9mIPWNrLrUSmqvwVeseYb8BBG3ClHMWcB6JSSXFo+L05mlrVEkKgfJcVtTmgqMET
HSApWvKumsDfS5bHMUm7Az18cTizXC4xs3p4dRom04nUgnS+COWwFvHXfizs05iE
9j254A/qmRcas++rC+369Ooq4js3dZImvE91zDaMMKRJCOGGOGC6RpH3JPZIyTxB
BB/jXl5LSB152wvWKYZ4zLWPMLZl1DXHK3K2dOe6rwomOdSTI2LvNwxDekNd5qiN
uUb9e7AlQat7RhvN6iKPPSdGy32bXixnVb209MmdEcRSKT9BNcuk2R46YUnpQJxR
ipx2XeQVuMTSdSa21G0D0Imue16zuswgAMy99brYNkUwxRQLIHyh90nntjYQcUQe
se2+wNLPTtv2HWgGjrnflCIO4xBg+Y21RufJ7zigUOJ2z72NSxiTMN7srOm6EAHD
gJzuacgAsFE6/0QGAZcVG74d0zJq45s8Cp7HX1aScE1Vjm6rXSmnv2wXOk5CP0Kr
kvcJIO3HsJ7TNIC0lepy+/Lg07qP7q5FgqbvjDKmnGFclBajhu5AO+tdbUR6V7AD
WL5IP+LFOJB5iBZYg4yI0yyfs0eyxYCcp5hp+7B9ltfpwdO4x4HF4jm1fVh2oSLv
8P2Xy6oYoJk2O9+70n5ygz1xM3MPniUEIrZMkrhVwo/pUNfM0j+hWBNo0JvDju1G
v7iCw5wO7l+Q3zULH0H8uh+ADpKvFpUGRcOEgwErMFbsy7qPzhEGWuUT6eBDVnTL
ZeOBqlHbtLs0M2rTZxp7G+LkrCg46W6JmLkJuKrAKy0YcY+JT3p8bwWGM8OhNpS4
XOdnPE/NZUeiY4Mqt0W00ixe4W55ykwRnH89N1jh/aVtFS/imJF37vpH9ZBqcvhe
BtrMv2rILqdQXOZGNg10P/ioxnioGuWYsd7kbAi2/oKcZyGjoiG93smskfKUYPqw
ZiRNoiiVAWZ7g8EBbyxsLsnqR5E0Hw+0rw7akm0+I6VEyV7PHCr1d1TppYq8xmGE
19s3ELfJeBS7LFMIuWBJ0Ha5Z3mqhgYElHCBY+UyhcvGOK8RIkWt/vFNMGpzz2gK
okVgmfZeT5ShOH/ShtGPJzvUvGvMuE51v9FBXYwXwQjqB/xcwpfQHZn3n/kyKYOh
ZxEo6/k/YMCtg6CGwIs96AmcVv6xIS+7i3grhqAO3pZOpb8GpkTZOv7QBLtG1MO1
dfoMay7lVrFz9fWolMye8Q8qpudiZmjtwQf1RDre5LxVY1fJXFPr7nod42wILIdG
SHNRbeCxQa47R2VA9NBay328pBaZUFSBoBCKqZ1mVUxy2zs+VuElhwMuIPJGehce
WGYeC0RzrFqqj+5awvmNxx/1mbgeHMq8F3tWDaSAklqHtwvXBAFW/1u0Kb8mYHCi
rv/C3SLlebET3pI2Q9FczWfIbKSIJ22+zuRk+Pm5J03P2PWkU1xyqY19l85+n/Nx
CHph/xjMToRbQ7Jn5NL28glfRxVNazL/0VP8PbHUsfYgxlgh3NiBOVhY4EejRTvE
twY3bxincpmUeh7ACVR1J0J3zP7wtGU5yW3YcKkkXTPgZiXpsr684vGboeLEtt6s
cK4gMGawFBkRLGsQIEhS57E7/Kkp9mXwSvUERXFZVUlXET9wtNHNNGyxGXpAIMpd
yDvkQ2uF21M+PCn6P3MZX3GThY9EVZybkm/wV4tZExw4Mn6WK7FPVvkmXHq1blvZ
BY4c0Hz4M7IjEiznRXdTVJolVp95nuQLW6g+wdJ6zhRUwv+CcmFgarR8w0b1Ad3I
KhClsTZTi6BAeWp3MEBwSc1De9cNxfda0USaMrqYnkhP/hMM5HfFp+LHc0lY+3SK
tWcOtMtdL474yIo4BWugxVi9E5GFd8IY2MQD9C+PXNZ5AUcEvRDcIuPIq4clS5K5
AQxM+Qq0BcuDvs6ow5JbL+wJ5iI6NeGFNZFNs5gW6MXpSrLdgDYoT7rymF4jnUS1
QooXDFFWZ6XvJWzHdxNCa5mGCHJooVCorPZjxNW2ZRjW8zqIBz1/mfW6AhSk7mjj
iC0YP584+nyXHXBkzA+cGR0BPdAtbD5kYIHX6jeX4+QdXsIV0viVmo+dViZSqqJH
rnslHiWKPaF6CPuPzi5WxIl/9xsXm10EdXPyg09imExizy8nssjge8qGw5YwQ7KG
dfI1MPbm62c31+af7LyCS3S4QMbltlFxHPRjg4sIF1Vo4L6Xg0GkzMzPQKv/ineZ
CTJwBGz8kCmN/O9Hv9K2VYlKN93/gl6g1o6vxWLfvvhfop4AejRjLLjbhAhB9UkP
wxifwISeD8hdGrv1V92XocLdehXVMt8DTXPOh9rsE3dbZSuQeGNGD9dxd3uu2QXY
dhCMTgTo/N+CijwiACqbQHWqp/w2AbsVad0dH33yDOkkG/4eCwujcMaDZb2srGlv
SIfXVK2SLiyigszVjzcmh5ClW5ZvoZErHsMVkj1a4HXHJGLr1thj45N1A0Pf39kg
ur3gS0i9WVsIBWvsOfObUJP8P5CNx9D6JcOcdctYj37dILkF9FnPlWLsyFONNmrA
K3Y9wAdzILP9X7q5kKUwDOnB35HRSCCmDqeKAgBqzx+avYuNbGM4bMPB8UuFrGWP
6shNd1P5rKJ45mkgtNgPAw+QdEJdd6ErUSRAXhJLkAmi2R9A31WQAe+Vnvi8EL+l
btYLvHjixXdFXizaXxjyrUdLi9pbzS4WBvpDmtnCprVDgjTjO+JmJQdZ9R3KsT03
UBGX4aNPIaYjpA/K6dGr5NYdzAjX63Q2MuPzVeNfsDRwDsqQyjQlSFoysQC6TV7l
xeH8miMMMDyejQjdVc+MI5ZIPmOBGwQ9Pof3MabxUfbDD8Yq5H+ak1qYGDAPG1u6
lC9yaSuEqFBRJnP/uNyt9ZLTQwLbaADXcpsFb9IstubRweF68E+W25KPMdeipd4S
aIcUZCCtbW9eVOTlFkxwrF/w6L2ITEqG8WoZrd0Oixyx+grJ3nyafFSLHbiiY/E3
8ek+Ps0izk+pAUy+GOUJED3NMCkmO3MBv9ldooPFx/iCZ93JXb5MkSzv0JyyNpRu
9r4XVVykbmj/e9hsuDZKEkhme0KzC2/A85RmQnvav4+zmayU3wpnFOQXENO3rqHH
lVWQ9Yw4lxjMaPZSGPmjNL1KwNRYvEBty505X7r7F43qvwiPf7pNbhMKLLOaNCHm
YGhrrC0G5iFzhQLTmp7LQmcQ/0EdWxFK9KhzIWARfvEYULxYgtK70ey5MPunlou/
EikE8kPpcn8ZmSgAt3tj60cLKvcrATT4lsMcPHNRvJWQEUJb2Bsv5lcRDvvlaB9U
oiIkC8ksS4/geMQdfRapnEOtJNqGUDzHK8Oteew298sqeaxkFILpmVeE0rGOHYfT
TOtqzYkHwyLBRMfiCTh+q6x4MahJRDQOe3UJInBsj2l0HSLXntLQYq2L52Xu2tmz
yt1T3bX93KtZuHawiZjgkWJkHRDuU+61PLKsRnHB5EHxf2XAtoeK5LRW9YJxrRpX
+uOFpbQXeBtq6fOZjR6QWixTd/7F8XKfW1w5J3X68sr4MGc9EV1VvsCHxJyVBmu9
PAE7CVmH7w8b9te2V5QRKeqfVBG/4c8hZ8Bi34+/f54N9GO1OtpDmlbT4S/cICh9
ZTmTVfWVyy3JcKP5cwQ2Pdbsjm8Yvdy2amn4oK37x+gvW9tOnoJuqUpTZCx0PKTG
KChxSquw5SrkNF0lztR7vWbuAASE9lzaXBNGmB2gKHRUl+G0bVBrIGZaFoZABcxA
zo8vWZu9Oje5cNh4UHg1kpqJrIJzzC5p5Avmx32SvRWTiPReTpHO9JaAr8//9cUz
g87uU4T6zKNXuuQU5C8AQ96zn/lIXb6HLmI084BLZqpQxkwqPK6HcN1tNDBahC55
emnxDG181BrZvW/HOhg+FqKdNTUEm2h93GRqok9eNs3IXqgrnPW6zmB/4GTmLjzW
5Dtty9G/vu7VQ9NBCCUyB0qFeKFBUeiVektpEZi5FSONG3MgdYAxO5SbSDY5DVAb
hUuxBnDyTznpB+71JA4mTbEhc9HQbY79qIa/x9xd5hTP3rtYqDU9LOJsPE9Q7qLQ
BA39cFNPVMuWr/A8WEJPlxxHyqkJuY5bgo8kv8h2QvqHI0Z1vPZcxEX2elRzGl0M
r9moVOG8okHNcmu92PvM7td+D3ZFED26zOxr14a1AvaiKa9vc0NrcZ5Hgt3OeCtJ
Es9vxZ3yLZcF5DrRL2pMiUJIG2SE9cU52Tjl1wcNmJA2q1aWMEaIc10PqJqXz4ea
yK6XskW+5oDe3oxitqzr/+ziNE1OXyv1ewrdnKKxnHwmgAWn1weTBz4YfX/5uijo
qhfNuSFL47EYXmE2so29n0j9xwemiPZc1ICPUQYY+uIdTxJ9Tn95BBDdptVwS4nv
xfLmDTm4n+aiFx5m+58ZDuJKvQ8YPbgYBVUMo4NU8sjfdFYV+W3YDkkF13KW2vKf
i1ObSUC9lo6gV/RW0qb7JcmKhYh/4iymigNBkdzSdpkTWOyD9OkWNd0Fkv7VUpgk
zmE+3fm4ohAHtCb9H+gtI8upcsX2lRdfdQSaVU0HBz3EDWCx2OYYjaWGS5fScvdh
5lBdwNY3bMkeIVjnhgqvsEi38g3KTGMbk+dbb4vNQS7Rm8qdRrHzUvVtia5Hlzd6
IddQ0GJQ9em8obUKlTUKnXNGYKfTN+pLUuWuWrLhvfHW62r+5Uh80nmpjVzeLM6S
mEvyOQx24HWmprHTJW9GnOPig1vpbaUfl5sq4r9Z1DTZKmqX8QAyTlPHJUYQ5YtJ
TJ5pCQwHjf3K39leAQkwEWL2xSKHkqcvL+VJH7kSaJdKoKuJc6REKyZchY0cdwAK
DJf6RcsONumMh5vMqpa0m05qRbkfxG0ip5rQoXIjXEIol8StAAXgaJz7nPp/5Qhq
sucCv5nis8klazZmoDQAWS73ykaraiLF4mRSDvYG2eFGP0d1L7/isTmg5uBDR55/
qfBGtsNFDrv0HW7EWGSfUzzJ613emY7ZqPLj87TlQ1EYzyenyHWV9DWGFL8cezXi
qAqEXSrlq/5SNmX9ELfu+HZutifhyhWucKh8bPlA9W5jM6o6gSZwI2C0QDxXj8s6
hDqq5DxD10UFll9eNkSjp1e3daYnPbk81Vs5/EF8B0zZQ7GZGH3pFWZEbTgRws1K
VaqoXTna5RSkd5M5s0EEx4PilpCFE6i5gWqGXQNx705onASf5GNKwEZIE3t4CobR
vcJQD9VE96RmZgfE3PztvByuV3x/whIXdfmLyOR68TEddJCTKprb9Y/1nrM5LDVa
gh85U2AI4+mfNiQKMWSi3YkODgjRfpToWGADFPrG72GLP7/cNZQjkcgFHoSZZLol
bHC45GQOJMvaE2wic3B5U8PJFQnerDnDrYVEUPAckqjrP7itSJel23CByV1fJNoT
pX1Z5O/YeuBA3YGwRExu4fY+K33mDhG2vzm3nyaU9EBkjb0PpJM8JkZTeKdfr3+6
Wjl+AuJftgAw2dXKL+v2hIRIEP6Crt4ZolkNec8Oxq9rvjqoepHlxz1/EwqmmGA6
PFl9M93ICKxQr8xEmiom2++WkhkqrVgZ/bnJ1ZOgxoqzTeWJhblrsAtgtpU10gqU
ebaqX4TIG6h5nQcXXBP0SVi2ucjmLwh/FrhoQO7SLjgNpnt2HmHiVjALG8Jop3/y
5adIPaSNKhakp23nVjFsCVUzb+LFzZJ6ZXG/LjVOpOeya65Nk83qOJq8OmEwoUC5
vFSfy1gsDuwxXF5uklBle3zzh69oFJsYwACvxXfjycZKVECHkbtwqhHvDmqAkLPV
ChaYlKrQ3ThKCnHxfJtsLwVEVtDVGMCIKt37uthpS0uK1JfzJuH/y5bKH86ebx8d
5ZjxC4hA3Qk2z7r3VpKHBsA9r4UVQxBqDZX6LYDX8wMr916y96vr0VSdBfne3hZl
8c9wFHJ0czP0fF2hD/NkSbY2oa/feJwUS5W2i4WbcjlNjGp/DvNGEfdtgO9PLpFZ
6G5tPFsigiakjM6Vlkrz3HZA0qGOUkhJ0QUV+T8nL5dbUd11Xo/bEKB+5SwVYkLI
js5MXDb0Wa7FF5fI26E9IlbT4kHNRowQFvubJ4VL/4MsKlEMWXUlm+2XmF7lGYMD
cAx0pneX3c9iz+EmqkosHAjjdLMdc5Op5AAJ/ywzPgH1MsIxXW11mkTJT+yi81m1
kcJUDcYRFGx1Qv22r0QDJn9s2Hk1DYL4LQdocH8SOvpYJAdvWFwTH/SbCSQtAZ91
Fa1Gcz/RJNkQi1598G21FbC6lf/UIX0SQrKd+bE9n+PhC1nEMXQPTq8ymhuj8uj9
OLdzNx8kC//TVlYOrQHdRZC+65REtuZC/CVljrSNbcgQRb9eWUy7UljXQf38PsYh
tbhODzHphCVlJXyx662roNBhY8fiqVt51Sfu0yyKbu6hbhyKwLwuF9bCgLHWmJ1Z
SziqEohTUfWVaBKiwEj9DSY9eFV/t0fp1b94/iuxyisucD/hlmam35LkBtYx8slk
AQgwo9vwDuvgEpCQtKJfSOcyRzIFJIzMYlDA8SjCQe636lMuSmsWBzwp+1MAUu9E
FbBEMgMzOzLoIcOsHD0H/0gG5ordN74sSZCIBkE19nZ8F9eGCXtTlpUGXozrXKaJ
xVhzThevgfnunizP3vG93gfBqjZ8538GT/5UiEF1ZfF6YHlISezKx11NAarzw2G6
WlrWVc7jpDNQwZFuR1Rm8Pgnq2vZwlZZSr4l76YSMxGxSVj7UzDjDW+KppMpgI5V
06MptLHqP37lrW6tMLmX03aKptRGyY1XLmR8su9VgJpuG7cxx2NyT4e+HnN9pEUY
yiL+4TUAsDFJG7n6Z9GDY5uOwf2LflSjArt1AuXtChUJlKDcjvhY7W4Wcx3O90e+
sHsDtKS/sYnK/T+T+JqKK+213Xce8LinRtXINrp/lLUih9LA0cyC4Q2SDZyDBwRm
GxUZqBugvzXnSTsM8mNLmnugqFbJxFGdn59ITFKEcKl+ZiVrxGK+g4wa5OxWFcJQ
hEiIk2jxVKMut8EkxvYIQFUQ11nQifqi/Jqw7xYxBVMz4DFx545qJ4faTThs8rfp
DO8mSUcHbpMho6fZYnPek930jHC0kz2t4U/xnOv0iaStPcWZoigX2O/Mag7IhqaC
AKBZL0ztHwgIX8uPJr0bVdHYLl65s0qpOeqxywVsQFv9Nv0QrKYl59GBAHxeuC2j
jVtKbjgGvDm/oWLPGPo5s31Q52c4rvVZ5CVzIOpR4huW95NxEYfT9ggoMHqAVrIr
mZ6ugV6JA9qLs96eJEn+kgUyv/5B3YOGgOBMAXyOl/k1cR+XOB/Z78eZxSQkmOh9
Ky+qx4u+ZrBgByzzU0rDscIP2VFg3vSKBXiQtwRVNC/S/gqWUG3azlKaW7ikWU0E
l6kCMkl9pf7K4VOCl/Kdl/7i1uNTKt6zL+gNuYzDGnMp9TDxpHnMmMDHyR17Ty+K
aNB+pasWXFX9K8u3i7KJYBBlHGaekA5lSr51s4zxadY5oiA44ZDcaix70Y45DhSX
dFsEwYQ/RYAPi7RnBXTvIQ==
`pragma protect end_protected
