// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:35:35 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
ogCrhGM2swGWIl/Of2IWxEI9I2oPGUxMfnNhsHZxxY8+cIMw7x3obWmJCVB2CF5+
I79hvzUGLEugv6adid6RpkJ9WvGAo7XrneKahc+hkvndPnM4jmoef5pGpGx+ezLW
xbcmuAUxoBRbfgGJyIB/XBeNMVJF1kgGh8sYnGQItSE=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 7600)
WiKSpzYA/5P7RWQ9/ltvWElMVao9ig7HgQc+OH32DykbOmAKc1KGm6XpnHdEmAO0
3FmMi6a4aHy4WKsQFRmGadRGciTywQJrUFQjbJtsRa71mMtT+7oHqVJ2lWfwFRKD
C1QGJXyP8i1Hk8gzzrGFRdO1oRLccllCQzXhQSuff4XrNn+rw5s8IXLE2uxhg6q1
+Z4o3wAaW16nPHpRUbGPpnR4O7l0ZVLacgWwY3qI8wNk8t6gppgZvd95c7v0fa6l
r9wZNpzw34TgBLIawlt43gLP+OBtsEYoi0HmRILSik/U0I0tEtVH836QQhVG63Os
86XCpYzpOugVZw+jVfOzXjnyZaeY6VrCNTHbxW7FhPzmGfal6avAkuW51i9vuZD4
1jmmUfx1VxYgx/WFxxAwxfiailLGO5IAQxXbI6pdYgLmZLTSbt8JKXQqdubOR0MX
SNjDgmdB5KV+0PFiGTuLlJEEem9dClUy8wxwFoYR8lcM3m4Rp92vGdDYe6MmYohd
YatfPJqwCkkHAiMWAtA7/B4cSJaenm4dMs25ExYA1EdnyxULCV0br6hEaDRRU3Gv
8y74kL6h08KgrgvI+Ju1h7Oy5ACNJzk8SWpgXKbj4Wb3gNaZ5IGhMsaVYeKeSADV
9EMjsXmSwIosQq0CurbBGjnrslAAJYWD5p0eV+90b1My8Bpe/pbJoAIhbF2EMwPs
hlwIV25vkAOO/e/mGFkMGq316HevxM7qh5sl0CcgLK9m+7s6jfUruwh8IsikvFor
+ziTYp7obEYW8HohdmH7x7blBQjEPd9Rwh0Ne3JXDw4OK+wwZC7X0XxflAcFzypi
Fznf6db+gzFDR2SYL6dKg2MitLIe38PTK92BtQjMpseh+rN7QQoNElmPWy4m34o8
ai7SQWn3HDDI3LCf0by8bfMZ4Sqn8cslfbBImEUoklT9pHHNSNdvSXC4V8NCVGmO
GDvxcKAm7CMmrp7kErqZWryZAIM8eu/xZiyLLhNHKAyzVEPTN7fdiKzR8s9eBeqJ
Wrkm38PFxEyRSd56eZv4vJ7J6GkuANTYWKfp2giQsyhixZ/scDUR/NWfdZevP9Dp
AoN2OVz624cdZc2cT1DVy5r//uU82yZAYsqm6PrOilD0WjqMd9QDFs/lwQX3ndAJ
W6gNQAexIXx9VWcju79OG8+0YDR7aXE/4N6DQAbblaO6DT2IgR/nYVOJh7AtCfHM
G+O3XeF+mi6DtoP6E1rniDZUrBpeFc0a85TfsBiIYhfn+V+pui9LfuqrHvaI0rbc
/0+WCuPCaylkGtMEUsR1D5BJfh06ifF+CbnHWGXCA8+JAdFe0mffTboxmg79Ra5Z
ZLsL+mW5ldQqLKejTi2Pc8A02qNV48COKxI6A8ejfQoM7rnxeSVcXHKCGAI6+cUq
pxnSem20/J8TIjnChHhi+ip1PQx/vV629z2qujYY84KvV4L0N6BwgFHYD6AJMq79
fEZXmRZzfZu0LNDZdJhQLQgqgJsEbO2wMqTFxizAZFhlDs1uTiJ0sSLBzkIPUm8E
tlQOSfXVmOgPebWZ8pH6oorKielkYBWpaSkZv75yxUPCevA/ee8dk0RcDFMRpjC3
REPbTQHKMtrRuYOOgycnvnxhbZIMDlm7a4ZbfKffVb0vw5aw9oArFe1zjQsJypoZ
Mj9Oz1+etgyVK7Yb/WenoqcBYpLqYetL/OpDI9LtFKexUJTVtse95JJCnXewhLW/
w5Sr9j84PjdNwRVEIn6owtO2/mBNdp4Jdca+TJ0G/DcAecehvyUofiVCsXEc61Hb
ffpzDZcCJB+JUN1xrdtAXUXTY5bA6kJ0+NxUku5NyH56++iviGsLEiTLkjgkxmMu
eGgXpPTLQX8pYKwWRL0sDEUyJee0hsOi4TfZCxsl6yKU5YA6vDppn00BYCS5jVMh
51tG8bt6MFYjja7aIhBk2vQAe8R8Pyp2IITO+s7N7PAnNvWzMBrOxLMedzU9xIkx
o6EMcR29zmP8fE58sMwNaII+3ND+9cgpbIVYVme7mckBHrbkCwpblfhZ3AJeRSXu
SJCYlNxs6icrIRbg54ufElRFK4c0nrxB+yysjwxOY+7qOn0AAOjkU/3/0KV1antN
zAfQNdz4UpH+BzmKmlODU+eFG2B+LwEmT9MsrguUCiwG6ZCOHuOTFYNfVZC8V3bX
ADDIt94zRLppbFek9M3LDN8iuVqrLcI9WzFs308r4jrMJNN4O04y0OjX9u8yhWoj
WYRQlBhCxlvYdEbv7YJvakIrGU/p2e4BimSzm0UFNg0/aoKFBfHU/tqvTLDE0uTQ
C456Hf5+6MLoVsc1lTpukphNcja7c831FRdbPaOMr8as93sxzntBaMPdKeaeZhdK
FKYsbXIHjTwot097dIVpFtJCjArKUkojcEX1s+mm14JElcWucD0cg6s/WYg6j8Bu
rhRcnrjASNx+Ht6JSnIVdDs9sJUrPgAqsv7nOr9ai6/7xR7YkME1MAQCi2jQRMHR
8aAsDtwgiHV+pBEsc/p9xj9nZlGWoVLvR5gsPWnAP+Q6osXwIiNmKHJ4eycPYjlJ
CDg09S4L+cfiBls+Fw9aklIM4OOrGnyxEuyNwMgE7VIajxZ85rf2gzPJmnS4g6Hi
Rrd4Rlo7qNFrBhq5QFJhQJjRzmPUi9gHDZi1GA1nD58u+UstXPtqCIjQIJG09Vw/
jqE6qkOfyZYjkFFJhlCClLJtESHqQgQOW8I7BrVf/FdUI7aSXwAXfKKSdq3rJMJz
8l0EDBJppKLfNXt6/vgq6I1cTMMSoThRMUDeFgbr+nzE4U3Y1nYhdZV0HuXTXhlm
AZUwVY2+VLRr3TXXz9vmDj0V3JReobTrN9CCaAWgb0JLN837SNHjfsvEDQtGN6U9
SZUa+UrFUfxGhfDOCfYBw1dO3C8S37n5OnszSNgwE+xg3/wnxyNDeWWnWx9FXq9r
lP7LfmTyjvACZHUdskZG328x2dqVS2mCk2lAV6Ukl4YdJwq2Kg6HR0B1RHvQdoPQ
XZngVEI+LtN6JAtGw2gmBeC/ZQJ4AYEWjBx6Y0G6pOt6nPXqovUVJFxUgho5hO/n
QU+KcLzeuV+lExjNLQnXd0enHG5aCS55XGpH3xSB5lRZ0NhGu2TS52zLzFiUBW3W
qF/azV7o+QLEB6oiJixpkK6roIyRdU40lNk4RKh3ln4ucLdsSgAtFnpa0GBSXpwg
cehdb4E2wftjUnwgMAr6YYPSumj1kVq7yWJEJnqKOVFYwbN4YVjhiivLsCAU7VWf
b3XMU8g3ZpiX1T67StgybDMIahyDfJpOiKfyjXFjY9iZrtvjAH1RKhWR68r1QILv
zI3UGtzVv7ePT4vAY+55Ua3uJLRCuAWUwDeHX7bX9rtvdYvRWR3FAGR6FcdLKr09
jC/M0k+K2pQMJBnrN/Uwu+RRVmF+lFtQ+d3hwEY8k1u+Atw4ldwtZ61771S7wvhR
e3iLBSQVQEKaOllUEjU//iZj3iE6u4OCvPppreNh67NRG5LBBmZjP+9ZJBvaOrcB
Dv+U6P9RhIzUpTmWBkNBQz/4cKRNLGflY/6avQWcHEVFRDeQV/rYQMJZBhVP7XvP
SV+qtTjAQ3InLmXBWsVMIoOGQ45NMEtjLkFsgoXf2IOlAXdcKL1PSt+00Kdc5xaD
ImGseWj4wpTD8gzh3uauyITZ9CaE5EOpC80n/LK78gdRC3yBJvHe7kIkFRh176dQ
Be3tvwwfwk5TppYXhU9YE0Qq4uOJH5Qf5d6i0VXME740lh3FhcqoDNVaFdH9UJyW
yif1JvUedZTpU6x60GbxttHL2IMb+o4ITINVpdPZQlvmoPYd8faL/wF2G4sJZcD4
CoebOdj/W/RF9I5c3PTFIN77wI03rQyd6CF3mczUj/piJkfFqzGP+VUU+uzV0MC5
sv3mFnvToe/a/nr+c6CWsZUdiffSksQW/JNsNsDM5OX4FJzQXkkYQBwSXCWDXmYc
eSfEAi1tkQ7GWP636841hABiTO4quNF7Fchu/ogwrTrSHEauziO5lEJrj/o87/6n
MmKJ05myCi6mJZyGCBi2PIeNXLPgTVf84cgA+C2ozgDHcj7Iw0R7HnesetAq4n7h
IMcPBUGHyZ022l3pSQaBEsCQ28KQ65OLUK0E8QA2VpfzVQcmsKSbJQo5opEVfKhf
gAasbnrkeaOaMVGO4aFl+ewKcNyY8awak/sVf5+I9y4sCOIkMF4hCcTumQ4P3YK4
5jWJMpaWV7Yt09DJTV9ulJ4qZG9jW5oVmgY6TORNIjt0KgcHAlQxHtoh6P5csyyh
ETVTZ4ME1mS8g1UgQkBNViRhyhj2feEQViMdYfxseUU9vHh/cXWACto1KJd2YBFH
sPsStOVpQoRc6aJHvAi0QYLZRkLqU1e5A/94wPFy8Rb8DAoLnqT1Z6zmnv19YWgV
eZNdSYoErO5mqazfjCLuMoIKJbluMUSqLysvGD0jFHIs745OsFE74GQ8vwFH7qw7
pOaRje57EQSTwz0D/bxyuz4bWC273bYyHp80y/klVfnk0gaHCBWQ5CYvNZ3mi7UT
d6IXeTeFm0eXwJmED+36GzO1GC3opMrexCaJOwBpBtEoc4ie/0SH77qgAeQn9HHV
wTle2oo+Z6J5afAHt7JsZ5z7W9TJo3gPQfoLikfbc+2LABgLe1itHne9kpMKAM2e
urp97SM/gzTs34Mb3LsNnm2DIxY7ipNoc5TIcNmF/AG0jFHAnzvVMOc6Duk2WZX3
L0XpKH5j/jv+NRh+jkvmZWnchbqqvrtoWuRYwAwFSrpSBE/UzdzNtYCEJmujVAs2
DwHr7Q1KiytM646WX2KISc3mpBUaD01KNE+AlvlbrSpGRZ+iivze698BO9PM9wpL
lRUq3l+y7E+Eu14DNDOdH3j8BEv7/6K+4XfQnHfObSbsMLZOPjnzfh3d3NmiD2+N
cNADTKwPdg5jAvEm5xXcmCUM7zU9gizs5y9PUOcXfRYnK6gG+DSrCgVADdERXf+a
KhyJ+CaaRQKzvraGHELaJZ4BSGKFGH1pDLOXbQewwpeJP40iZSqasX5ZnLNpQq1U
kOg014mjfLaRAas7uASrTqhTSx5tHSNJC8ZrhebcclIH2cIxtuq/xfHS2AJQlvR7
nHzREmXaotLsp90d4wmEDVurz8jDU5oyh/D5G52LiRf87KvYMcg+IWlXHySTLcB8
pTA26smkM8cA0MHvpAiCbCwEyjJXObgJLVOZ4LWCBO3hR4N1rpfl1i9xBT2anZhk
YPYNJFtVcui1+DBMpQ/xLrX7J/GiTYU1xVNy+wxrYeWigPOuQrsTHRvZkv/qwoqw
3eAchtPNYzXTUwNQZV/0Jcvs5Jpqv+fqNpnHbbmc8gBXMM2fwaKjy+NFskVp9BS3
FsOE63dE0li8AdEFlFlB+gK+kuScyHAZfG/cwyvZ1UfHjVz/8aoMo12p/PF97jyF
ZYoffqBxqi9DqxZXCpgMrLD63CoFycNWQ97Iu+2/mmXlTZ2iXQCBTId+Z6LPfsmB
uLcjfracRAdcQmm2GF5gYL98TAQAhT29ch2MmmfADrNg9EdZtVbJb5ZC8w4hx0Ua
v9Cxg14Z6jWoV2YkMx5MUliTYT0rAMXO+TZfykqdRYvZ70JiIa8JVjB/sYf/JeAv
bNDNSfDNo0huUsUyZJZ8DY55cvjEXnsi+zkX3WVE+gdHcO0D8nk5TzoH+GF1o1xP
/dijhxqeCwUbgqFaY22odCseMZH0uFWcKkAds7UU2grUCa/9f4J+ET8JN7iW25a6
ipCocV4RwKrJbqv1q3ZHLIa3nLgmCOWaGC7xBDEXVb/iL1WNcxG4fOxQwb6CNoPx
AxQx6KQyvJFKakemtlSqWTOtBUied+mkRrY+L4reC2Iu3jsUn3FbjE8mRQedLLzy
1rqgJ3HcCVzQQl2ZKO/nNyd7wVnqh7BRFFMVcXrfOZOTTS3SPzSMZfW3iyjxxOcp
oRegRlQFRMbOjb55pqzjMI7R6yaguc6LCLB3ln3g33Cv2Fz3n0KbrhHz0xe/8nbS
EyWJxD3Mon/X8qCZNMrz9r5LZcQHCpAVMDGpDX1o63WoQfWMZXLXkz5xfnDUUIjd
0uh+yFNLjcQbveY9mFZ6/a717H9se68MnKqs0/7oO3d06rQyAV9SvNTLsGkdvhV5
CbUCgJSnuHXNCFeS5sgBA9KaoZLLoPbvs34rFerb61OAx61H46nEaCUQyvVCbAb1
dDRjIkUURpcrHdUyInbAdrg4Pvco6npmXbTBLDQmKa4ngUcAOpTq95TIquAo+DMl
hMPLstzdijiyWOQmj2hrJBZZSSe2skokLQLTe3pRGrjjM2+Cj5B7Xwz+4wn5p5ws
CnTAhqFPmndgYIjlIgZStT9y2e9KpYqONo8AMLqFueEcoupATc3Ir5nzaYk5bn4G
8CL4v/YtvrJYJOYC0fcHoyiPAwQQ5lhgDCvb0mbf4fwjhgsChNCBeRqlMZFrygEb
lroZDI1P8va3rhW3lf7wUiJtNyUMYDWaGSS0zWlnkYoOb5DLhMGBDEl5boqFavbF
BfydKqAP7Bfn9c+CJ0+Wux1DJP59bv3tJV3OVpwJ+wnHvQpKMpPaNasq15YiClnh
9hdmFPw9z5FVx6vDsDsodWuYrk9vtBySLZiQZz/YRlpyiwtIBkPy7bINlDaUYNak
gbl0zLE+Rohy2BOEHuX4axD4/GbPnaXZC8KjKCX+K3ToNQZ//UvE8tFAWixf3WRM
r7bvxArQ4ZcCD6TzRUJ28EeXs7p1aEP7scIIeip7s8jKO4Ql12I8iasS2Wex/g7I
LQtXOsmD5iV9Hc/YztklnZvchofyjApRio3KRgeZkmWwfVd39uSNjMroOyE/8egy
B7tY/35fNiv5oF0iGowkgaimEN4L60nweVbv23QghIiynUyOrFTiTpAgMCTRNwWf
+1VV8BF2IQSGobiiL3UKdJ0TZO8glUQ+WuH/HVcvOU/WdUmORUsgsMXEt1yDQB8B
YZs4Dpt+OoTnPjNRw6+5iZESniE1mj2DWldDc3qmk/n7FW0HIgYm9mdT/YPCZ7dH
I8DWJw4GhRkPqJRzjR4WqmIhwhKrfHM5fXBj+s1guJHeVgxwRD87Bde2QP6+ktUR
a4DO3yUaaZYDZpq6tfAglB+4gVKkCiLqaC2MJndqsOEO/hmLtrNb/KCGnbS+VbWp
lNTFbRmEJCUATe11QbfNlq1xxGlHtQa+c9YFXfZLLSaBpfOBTEft7RbzXuOKsTYm
OVx9kFo1Xfptna/glIC3dJ43rD1nHy89eoSlA3AEcZUOqivctuFjjLRG724Douis
xz2NHx5MBZGwlpu8v7InQ2+z5206iadIJTPDpJ0wHtd3c5iNhQlVY2yqlmVetVX9
W4ccywkVB77I0TvZJ8xelDqIOd8AMCWQ8KipAuoZ7N0Tti9a7qWhFbsDIiLrnNyM
IKip+EbJ8d0irAt2shVa+lB3dWVxNiw5Ow6KvxPEu9+oBkOGmIYyEjG2iKkRBbpH
koaOIi0xphLIoQJh+RayM8wRP9OZC3Nj/fY6QN7udpwcEpw+H0G7BBOBFfG98+FI
x9424XD0IHTL4eYRu1yfPuxeBxBI6tW6azFI70hOE3iZAJEPGGSVlUxMHnLQmN+C
w/7bisxe6NzkeOa3flpBmtK/fdzHiNnNDYAyYnc7dJ8X7uFnSRyhlg4l20rth1wl
zZo6viwkp0fuhHIAG8Ilo6iC/j/mKXzdowgCJwvKYEpQz8/zhWUPtWAcbABXZC2I
0zmeZ6haTQJRzOiTr8meAEyx4yEN2PZ7nXf7z2NMhNQobhOL3RRhYrJ+BYXWosFl
qK/gkYCdMIfsMxlCzHi3vGHcG5tIacZrIWJES08OzG+0X4tHqdWSKIYX1FUIr0xf
Z591iqUUxu1vFhAdb9s4T6AQd7Y8KAYC/PHTlLHRG7uWnvtIYhZ4Ua17D1QzxgOl
L12lnCO3K0SPqYC9c1K7NZPK3pmejJ17igpk1Of1yxuKlMr4Rm/cNjtmTjhmsnep
CH8S/g2ldBqwM14ivv0vv8sEqsb/5JCTaS8pRUqPViJzmsxGoUrM7I3EwG6rJ7oi
26b9M1jteiA3RzBlKyomrhkLg9L7YxVwG/BZGJOw8TVhtSturZzY4oD9qru0e8Hj
NiKBZ66UbuVzrbXzfpCYlgr0ioNHYUIHGXF9bgHXGoXcbOlAsECBGpM6LUN+KtB1
i8XyUlCWEfF+0lJOXYo7GfiU7n61A8xqT0ziwKHwuFpo/YqbG/PeM/VFEuL1FkWf
bTWXZm8hRZr7ltdJv4XJIr/c1kWHQV6FkeBjz85qpMhPcW1JIVYYU/mqrlJ/v1OZ
6C2SyIOrhFwO5NPR8KdaPwki050kMs0C9gMxIl8+CJfANasGGb7MTIQojU4VA1SZ
ZKn8zYtqBPQe5MMw3zkxr1z2QyfHRgq8kPgw2Aa8hjCrGCl2Zi6KLmRvXgz2srlQ
KbBfkNyPaP8IxKI5SeE0+yqWDOpeAi9boQPnNeWdHjIM1BXYqNh6Jv4rX2R8NjlP
5todGyalYjlQK9DF4RQpVjErj/N03xIhymx2N11kPcEDYRiIWzKN/3/r+A1hwlpQ
gn8G4mJl5Z8JWDRM/6DZFLFZyuzTIERFDtHXT9WkTrcYOuyZS5V6kAy42D4PRqtw
c+SnDKHo0sPv8Fv2nJItkGWM42TpogxQRjBKbaS3+kEORwJdghMIIG+IPZ+9DcOt
sI3CxpKwhpJKWLIlCrsTQTP9XowtX3a5qyBeXRmIlC+TblgHJxW80nH6ZYxbww1j
XPnCHqezErkrQQenn9LUpLHG0A5YBNt2bsag+jZcE4TT5/uRLUhTU9xAOfxa45ju
9qZT/EZyhEwq3J5bEsoUtgKlMkCPCIGLF5JQnNDOOhc3QHB7ndhwv0+ORZr7YXWZ
tuTh1CHSIJqSJj4Ju8mC1ykOWqIB4iXC2Hhp6FJBFCE2Mqf5riaaQBDVQab1HJ0a
1oA4l2gCwMZkmbW1Yab34Af8PiOBqTbdz/nI3cMxuQZFX6HrBaooX9Q69c+D/u9K
1utO4npzlwUr2EHFXkR+ngILWAmpsoJ5xMyikrL8ucoMu5dTSlhoFVVewJgRWTM8
koJELqOEm2/iiwkdJslRuI7IaNeHyTyEnXkn/zjBzC0K2j+uvLqbKhT4cxt0IrG2
3AHCIPQHGCRI3QfD3MSWntLoqZLEBGTHZBrcQsbzIOlIhtEj15C8lXgLQ2+ho8cV
Fz39xUpHAaptJd3te1xEMwRBVJ89wegYdRzb+niMSm86DG9Di5qFwZs7Qngbti8u
WFzvc3e4h4vZYJ5wn7IPY+4HWnm69lY2Utc7pw2ha11fhZ2HO6jOuToBOnHe/HXI
Aa+e05KwD1GChpXIUYzscwx0weP173CxOFOUuHNOp7AlxnUC2EFf1GHQgHLvOsPI
bvpmVLA0ZLGBeG/3wNrr0Ncw8hCTN6D7iBDfrlZ+4ElcxIWpUEsaTtGkk7+F5B26
8Buhnz8m1rjxi+ioystM46UrTNyyQqoDLbVn1m6Seva6bm2Tb5+OWw0GvSy2PYYA
vIwrwzFtXLQzjsrDitrFYuPXJzf/WvwT9Pfq1KUiGQpbFtUfiqXH70mx/SAmy1n8
8nEC1BOKQpSYPdqzztRGaWelW8hkejwJivjUeNFAXg5wp9wQK68Rx+dDqw9zk3Kn
e/KxB4+qmNJk9ydmPBwr898WIHpHBCYAzmfKjAH/QzGYA9dPHrhA+0KBtq4l1bR5
grfTUJuXIIJdkp1g6KtGDFirXSXMf2QdPK7PW3d4tgR6kaBeCYKnu2G1rDdk9Tjh
tRZxbl3y30/Oh0Wi55MSFEGrN3rnL85dGIFQZjgGDVTprGdwRTRiiR1TMcdeTwmr
vkq9OxpXfQk7/ThI4icFQWZXpI2cvAEWvRiXatYslBfVnmre3bXBHo1tlguu3/6f
SrVsg2zPRB+xa9YnAciMAOtWlpAZznkJNOsW8+X9To5QAw0udLELfQGf+iDa+Mp6
qNTVSgS+BnmpsSqpR9tDZ5mroZa7UdYKbZFTcMVMFKbBHqVPmlP6Mi1lMjrnaV34
+e+FIlfzFNo6wl4LOtMrfPE6m3lC+EZnILbyGl3baKPoGOJsaOcriAx/stgIp2hO
5dnkrtsInQagjhoQ2V7y1A==
`pragma protect end_protected
