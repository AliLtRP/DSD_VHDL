// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:41 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
M7n84OlCS8IPLo8cYui+nn6WhzfhKNg8lYVs/gDGGrVAT7cFqCmsh6tyLHzhTKaG
qKFIuJjhwK7TYHBbe9YI/9lhe11paqxuQOqXMtdCwpFVz7nFDAjYNPevc7iSLOtK
uRGNyRPq+bYs3GvEhafXsOUdQmenlaZCKFokk2Fdj2A=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 2928)
sxXiJO/LDpQ3YdGxH3CgoZrkRvTj/yNQAWkFXP0UUUCLyLEWV6Gsa/2lh2GZjRDj
EU3bvtJO1Ba87/y0CivVS9pCGZ3ss4I3Z4dGqwKsBk0CVHFJ+ke/xsIyr1XCx+Pp
Dd+BpO4WmAbLPIr3ClSxnTFlN5bYzbCmaP4VHHxPuKD3txlQQzt/xGLXMdT8VdAC
YaInf4umffN5dA0zrwho43Syk+C8qkMqiGm5A07D6c+wEy8haDeoykI/FiKcT337
twQv2daAFEyRIsnoPpHX1wAU8QVuUOQ1pQLVuJX3Pdy23quj0iUZe8AYxiQPO2ih
J09/DuwSatIG9ZqoaBRafjd3OTArEO1UeqS8nU45T6nYeZ5IJ4zqXYAy/lp4Qfkv
dG1qrP0cLcmGwT+uD8hkKd/SNSuS3lWFtk3Xvy7MWNRZ88wIJd0QBwPXmBDKiCBh
Qsh4iy4LOVnm0onhKCHKli/bEaQ9mCjntwhpJp+t497X+r+1FM3+3le2WjxsEjl1
mjzkXmjTgIGYf3srF82WqNp+eSntibRy2zDBprMBG68A8DXHIyidPU4+72PA6/Yq
w2seuWIuaNRtcURsCChmmswqzh91eFENSzieuN42QBvHBawjwQzpRf8RdRv07QAE
nhdYAUeJT3KQFrGCwrd/xu+6zCs/MR/WTzcX0FAQ/539YNbp70lmGbeT125Ro/BQ
VCyMfnFNVBJSFAx1jtbMrRAMJbSQ9xG7BNvN5aUViOmuc5cs1cQxRcMYoc8hqjXS
G2xaV2fEP7MmdlG4Kb9zRIrBog5Lpa6UYAOnoJGr4Ax3RdhHxQY8A9Ho4rDRVotK
G36EX2yMLXpJaelXoGFvqGzgziSXn1iuf/MmAvlZ938s/PhsEDfI+bbJ9RsGOXr5
4paW8wFzHiWykqAGDMKmVSnamR3DJUi9KVpdBVcZWCXcgRzPlTzXCAr4Mdsq3Akl
OAQKe0JWeJUjTThncyPlkFkGUbIn6gQTOXutMHpHM9YxjT4C7lypAISZ+68uUfGH
X5NC8Jz5vM0+X9oBEDyONPW365YWyXmn+UyudqqBdlRm+kQn2OsqbOpwE7DVTUok
ys+w9OpHZSg7QrFvuDMzz+kY/yPbNpBm/K9AV+RpUFzeKI0AjyAIFVZ07zAVEY6q
9sKkgBeXKYbn6N3WZLaQyYzX3vgFjttRKhZVMMxgFWEA8T4Mb/10if/WXREijIan
+xOhhB43W2J8X3BgAbvstUPYjnxZ7WVR0BC+l+8OE0ctWwj+OgQw9ZnqE7kxniHg
hINIaefyJ3CyGxFgpxoVtbLCpT/Nm8u54O6udY76Hyoogden0bJlnGUDy6nIEFnN
vsI8lMzgsLX3uYx3yqgZYfmN8rWsaMZH4rrRZSyli6ntdq8G2QsruONYa+Lpo1Ml
YFSbrDOFS91uIFXP62XFTLNWa9ZYyFaUbVNiA2YkijaLZlyVL5o/qzPW7dBLHk8c
rJAXXGJLOX4O6BihdMHV9v4fAQaTBtccf6Hey/uaR2eQxfanq8KaL8X+98K4NRcN
TUS5KueBfHYUxFYh0YjgzhPg02a6YCNVsY4/FCEanzJDODrep59pGo6qFG5TmKyz
TMZRM2XZzH9xFm+yk3ziAm5bjWLOUfaMOz0x0YaG7PdospVe3L4bUjOFG3S+MgxB
svOeUjmWcb3Gd37sBZHpQC5AINDT+oQsXZvL0elWY3r/8X9/6MYkcKPa8ky0Zrje
F8Pgcz9DZdSvAQc+Z8oAK2A/XXNoBudxunYaAtPw5s6CBMp3h2t3jGXHvVPjFcPO
ahwzojKE8VsnQPpUe0SZWTF6rJKuaAk8zFrB08UndFs+bgkFWbz6TYwWEQqFb8Hn
KXoZHmQt9GLpHXYQk52eKjUC/pfNVQd8+kFYjoYt5NxOcW919SUtCR9d88iQGmO6
xlEE5Oyn0RsyW3dMZRdrNtIT4lM3DRCWWfNwqFefqPHoI6aORt5vgoTwQP+e59sy
MKmXWLv5Hh50yZaFWf6AbR2CfYVFxAY87PsaSy21fcuNqxxxt1mEhUtkSrbnJvU/
B5Fl+8ZY68Itkbpcf/HTHCQi5p//IzhoTzFs0fYmLVGsvRa3P/xs1cw5b0NcT/0s
TwXFebnsOvtEcSNXoy2ronQzRPJy3jWKoM0hD4PpapFiS+wvpsnAkDsPAWfeZ8RR
CKa12TIor7jrLml6G1fUO3lu0w804QlJoKC28rEJaOWHwVRoCSoc9PVJO4Q9mVZ9
s+gHY1YUcyK2icb1/lo1TGpgE9ZhVc/ua5tm8hJSfc9oX3h2AyVDHEGnzEoQJ+Vv
nVhXXT8Hl2a+ojI0ZA5COP4TARE1YFYa7R53x2KP9sWGTnUK6DfkazVDef7JQwEG
u3WC5VrrKK72SB8Y5iOtvQ8UhxRhMe6PgljnVHBPvieAqXTnllTH90YHEKPi3KD7
Eoe/ias+PCFOwQAOmqAh1Wii7dxlm3RpV2fARoQWPRQrE1FnkLG27LtLb1FwWFyt
FviKdXJBIDqArJWLGEPek/Jm4ZKQBlskxARYDWxXpR67CwblMKTcEiExe4A9OVyW
K0ko1NM9lAFMlrU8As8CCsPttMLik+P1XErgUqyQezsHgx5gce9knic0Y1CBuR9b
OBQzdBZDZ1joGNtbSxJhZGgtCoz4cfZrFgTiq2C/ciAFP3oxlGJobQx9o3N8bgL5
GmTema7ws5nJyBfLOu3+dJuLrW2Vp4YL3Ks5ohq5SxawPD3nd2SY2yk77L20IkMe
gLsViOqUSM5vS2NimE+l/7fEyZFT1RHX1ZaFs+HwECTm9s3Ud/2UrkeZ5zLBvAC1
hPeQOyVQpn/2R5sMCyxqSlMJa1BbD+ga0dvWoJNtU17sYhe0FzryPCBVAYypKN6Y
9jHuHs6zpGoC/t773T66Fvl1QD0KXfJfWYcrzLGU4d8fEdUUVOKGSzuVE9RiHO0L
V9Oqv9I01slEn+NdX/guqecY63FpSiOdUyVjXGkqwyRQ6ioIjRrhQSn2tAi2rRwf
fMuauT5N8wJD/c9mPK1LNaLlauyPZniheYZmW0uMh+JYqceqpyiAQT2rqf62GsOt
P1A0J7voiLZK/qbFEiiZygtY2nyE5tpGU071ZscfBrrFDPhy4vyIERjPUuHX3osf
VDSK0HGDc2mDWZZ1MYpissbwOjlm8Vq/mXmJWtOGhvaXZPpQOzo4vJ3WytE2PDyz
XKzUWyw9yfxdM4XLwswsZoRPGtTa4ApzMTDPvSUa9qhC55A8gcg1KYMnBNH/A0dI
qYc6p2Jn+pH5G87NfTEO44n17HXeRr3nCtyRirq1uCPiHbSt+elCWGpp0WgnK1mO
Qvas/sv7dHTz3Ss0RBG6/sA4uNCILq2M2HLZRaPpGPH/xlPYXyZ0zmNC8Yo6YTie
mdFjTB/sq8ARLam3EEEPBha2KafI7ex7TFJuEaALn5D5mTQhvdn021kwisDrs9jt
Mn0E9+uDMzbEYvDNBAna5RGKs3vJxmkgeDA/2fy4gi73prLBdsz75Sz5uob2GM10
nhXX5+xe4sDaneCGAc74/nYB9FsAXbkdJWW8QGrR/GVxbn/hgXwZUuJoXdR9bn5v
JeySTf5smISSzPb4ehfmRTsLrp2fAVzjDCOn6pPZ3SatJ6bFfTOHCJI1d22QnCis
IONBdLwY0rR8IJD058fukdYskVgXE2TDubUFNrFrshMwZOKZoHsxmKWfKwVkHU95
NfOGzlUIBSB2DRFikRspYA+YKY+cbWWD4e0AuFoFMDDwUFVyYxvZjXGSZMYAwey5
14jXAKJU5nUuSit1Lm9+mUGM4aXShl5dP4TIYVReU+EKwWpwSMvz1ikQcMbx0OsE
A7hEl78Y3IrPUlJ8IGsY3Z0zw8lAQQHSiMbF/nCkuGCJU4JmWepAxGLB4kO2L/Mf
`pragma protect end_protected
