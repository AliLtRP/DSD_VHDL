// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
OwuYNL0OkazJtdhzAjPD6mdVGDI3YiOuimTcdp0eXkNN43zeSu3LiGm3vcPg9Wv878DKnSNHaVDE
xhh9sQgNIXFfN7uJuyvo5IUyWi4Vw4bLjGXcT/TPZpHqNm4StYm7j4zoVByXHVoZWguwjFCTHLLc
FQTTsFKik+mh1oYJYUdL5SN1IwtBO60WBpGPKmZyR3IvAahsi3QeUFJ/w87kuxMx1NCix9eD8Oge
tmkf8NtZtf4PTznDni5vK8M9uHEXv7KsLc6pNHn7MvRPuw2U/8ATzUdEVKAdTPzHSkyGoG+PEPyV
NkTC8VRKfSim/HHhRmz+RMKozQt62WHTtuPJQg==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
7sKxCEJHc/Z2+33WwUzW6GYcvyRgdUraw2dVdYaNTXvA8lFdMW4vnB9lzang0okgcIScyZvRBLRF
vWk/3WRdhpFg03iW5ciB9a3+eB/NiZwKkeV6ZWAlpLDO+h/d5sZKoWxViSkTMoQ7mh9G+GMPJ/Ci
mwkQT1ZPHctm4mGrwCkRq1l4uAR+FZ84xNhfCEBI8XwA+ODnRd5S/07IN9Bc1fYnnBUwMgQ6F8aL
7qssxv0XJdfNTmRI26H16iXJAqU6a/d8133gc+JZWrtRZI4oiTwpT3mQiHxZRf7p8pWz0CocUwVj
N1TeKXJ5Ad66SP42Tx3GGpHzpxEpkDgUquFOCcTRDnxjZ7FRszDDRkJ+bVeqhgqTZ+ezTJX87eFD
Dtz9iCbD4D4hhwMVjAGndK3lI+86k0r2U8n/GBWt+YbqIdF5BXsLydfNL7rZ6LvlbnTTiFzeDz9C
pcnXfVqQnIZMJBOzhE6KlaEX0yH9N8qSYk+o5zzGLXj6zNh02a7JuQ5B5/7ERWfDYq5AUjnCxWUp
FpTJLH605uxxCKselF/DUAA+OocwbCI0smPCHnEQbo/XfTLk3nnhaLWqr8SeF3r/xbfEv0h4aQri
UJYTZAk4G3UujdIShomjzrAaq86LcCUzYa+R3coyEG/OIiTJfsR+U2FhS33N8hxXuoJxSB/esX6Y
D0XdoN8V++89fuRTMXcN802hub9E8txiJ7u7j0SwsEvb0LhdeJR3Fg3oV3k8V+C3wKOMfrp/qXjJ
v8kqBaZD/jsUmRx8CzwE0B1zKA8Pd55c1ci+iqn8h4GYIg5CGi8Xbo62yyK87K5unETKae9DXA4m
f9lNUfyOVcRx2kqYb9a4EjkJ+AIsQfbWzl2OHTs0mxq9Yp8n8c+oPjD4JREvBozG6p8I/cWDfToP
wm6Np6RMtKrASytyV+m30nL98LJdR5vbNLcmrl/POpTm2+XY8B0ydjUqEPL7ZBpCRzZ539Jx1MSz
LBNKyw/MLCzN8yxZONg6MQTymWszFMmAU48WlW8E1c1p6+jRiRWQwx6S/Ph01Lu93FFxumHvP5oZ
NxMGraHlUm7YcYPHU2ouOQFNehyeLh+fII5WNZ83HZ8+ulhIAPtQkZC5xwl6At/g1IeqWYO98eID
vN0Gal1PyEKT4i3TEdhK9keIqwj679of628KZLMbm6uPPZO4qqoJv6ZXE8xNZ3oZdkO3+fHfwJOo
V8fzcAWVPslhaNj6a8TganwujNnKGYfmnCu0q+IxsmjwoimKnn0OKUgmaHeUQp6w7t/Modx7+RwA
cYhHrbc8pLlNcXLj59uEZbKtCpUVyg7iOFkofVno3rCaLBu0lQGnVh5vA78w28UhDMbLObD7HPWC
Gmjsebo0czbSvAIpj7SndE6cNsiLN48e4XzxodW7jbWe1ptvixgWEf/Uvti0aiKhEmE39UOMWPqf
O1gJO6U0MhUIRY3bbfxjHZ7wl49NUSmpDzMSLCA3WiSDqxkMW/6GxnI0B+an4KN6kXB210jTtpls
tl4odIODJpZRRPuIY/f4FgLGAmHOcYwc5rF8m/i6FaYHjmBOl+s3PTd4LevoJUmUfAtKzaKh2lHR
geZltqUxd4GFcieZm04qQxpG1Wzut9wRZ8h82w58V5NS3ZOTxWzt1nneJTqy3k6+mbexxdjzwUbU
v2/vubSUh7lHra3YHNFglGa5o5r1A30OpAFfQxMLc1t4v7RQzrf2GpFuepjYQXxf9CuLPTdMg/LB
eKuGllP9Q8dUzlJc3kMm2rlLlQSdSzV+e/+CS7qN/C7XUwh/bQ3lcLkCV4IUGFW+40sY7Uq0B+tT
1NxcHKi3prgQKIo0a1gLt70A0t3CdztIirgU0+suWYoEUgWKudVi3eKFTI+Noclp+lvdJsiCUZbj
YMLq+evSAxzs6U0J1JYCGPq+dHFxkdabedDFB3fj84BdDmreGUekr0d90kIG0Ltc+jzzWnbffviC
bD+zZKfaa6djGRoz9dzbJpGQsHHt+l8klmdaJ5enFfNeFlTCDs1GP9CvwbvGYbMNaxRMvqU0xNrK
Ip63jCJjEjDsWykB+8uVKDwDTpgDHtncdfZleLRi07eeKToYpZdn5UZJvGo+FzA9FYRhPz1V2MJD
VbV4320ptKMqFBYgatorLHEjDhgN1E6L9lFyZ7eEVF6ivjQwS9IliweKm8BAOQedoJ676i3tL2WE
xI/uj/kNtBjAnFls5m2gQM+wpGkAR9lo2U0a2uV+FIfEbGmiIL5dwWL8ahoUksjnQ0zWFAXtxBuN
chntRjxtpnOOBYqAK1fTZLmqh3rIv88pSUjUZa6jQk4QyHpwzWtJl+8jwt76wzETjUSOT8JAaPJR
QDD7UEKKU+3g/z7Npi4yofwdxGk5CBq4QLKPyU3SBAZyRoWvSgzlbkieNrcsQhHCZubLAQqGT5LA
hC/59vu47J7VuZCg8Ob81T6EeSq94BGKDKOvSKW7g1p3Pntnn0TPKGBtULT1NuGiKAzqGeLkjHT0
yiJ9ETZY3FiwlIaj6RtTQl8+31KV0o6oTijZj31ta+4AwJZOI4cj+T6w2L2t3iDBGTsLKXYV4sTH
k2bH0lsPoDrcswaAdD57jTpzld5Ie8EjRN2a6aqEEwMQMRIVX11dz8VC0nqrExNMY0GuMWaCc8HD
0l0/yWxKYQkVxIyYOH3NEbkmSE8TD+VvT5zHETniT2ElaEu1mMJMyFH/hiVA3zunn82qZhh84Y4u
dEfS/282DSJjC587NZ5pKO5vK3TfuFM4Pj6GO7uqgO/Sz/NTqov7fnk0ABpsEyR98jkGxb1UlmdH
pOwLW6NE6Moao5aHd544Yo89aaPXutwUBgdZpxlUiqjhW0LO+1L62sL5ox9vDlzJBIyokCw0crfW
3m+eXJAARACYhPrxFxBUe+64YHJyToRa2xo2Q6jmVC2WRte4/XRXWMSSFpluv6e8hunopHc5kz4c
lVb+FZwI3GZmJoRRZWkmpcC1D8e9YjWYe6xrqJAymbeUDD4hsFSfRd6ISmd5YsBR50n3hkhegoEx
2HgZ+aWcf4sggjcXmQmKhyDk/EtsvoxWFLAPq86UYn06Ri1+C4ZsMJ0ovDwkbfUV0OZV5WwByk8R
tU3ZE+Q8T9E7tpHXSMWrf3MGHHT0bAnaI3y3uEMJMrbbBUo4WasOSohmmkzd8vGnTX5BKj8Bv2YW
WaExQXkt45y9bSXV4dc3mURN59wTwY17CVXj6N1UAiuplUQRvD7lCmKU5f2C/QUYFd/h/9iicEoT
cRYsOfF09lwcnybarftMoZEeKjmJXQnHi3oMQJTHOZ2/LLjybpX4t4xiL2Hp5fepxUTBeRGC/vGM
wg1OA8GSnj3qk8/Z6dO7hab8cD+vu4Xy/Xmufgl6vDLNhRR2r05F8HyJoFjqYR8hx5hSnsjOqMNR
q8c7kKI9m4rTFQeEjpI/6NJ22tiQA+S7vvCXBFMAOLIObbneNON3LKkI5us12prM6U89KNLz1o7h
ktcOfZ1SC76ZXi6xiNo42ppPsnE1cgoA7HKr7OcSfrgDSUSwp5mo/jUPaMcoM6j+oEOVgflYUfWn
4W3CTw3ardFDBAvbuzgPDeuEABysY5HFojA3PVQxvrd+7KAvx2t+8XVq3/zWkFvf6ij4LlGLOCfK
1zh4pDDxpOFk3xEBzVFwAAvbY2YT7HsvEIl+PL1fgLqAoM/+ZDJ3JiJN3ZjqRY9L20fDM+dQvxDB
CbtmZbrz6Gz88YjSkVoe45Gt0i69f2tzrC1hyE1iYzCd34V/N3k8ZDEoiUmkli7UDSAj+D09y5GF
hPpsKA6DwtdYHCj2TSLtzgRCT+686ONhuOheSZbj8niNvb+ic7aaIwnFdM1E/F1ytzBIEfP1cpw6
+jQnUorEEllBTvnB44k0nn/f0HnMEvwoIkTYsdkWOmuZ66y5nE3KdawU7JMpLx7GoAdmmj8fh0N+
uNri0BlDofiqh7JTPBBwrs8z/jZFop1rse3tox5LRmk4Fw4sxFNy5BEPEYv1qX7KkFI240tHDiDK
kPBcf3vZJyAP540p7aVMppTO+U3YnE6JorSvYUXAI495nuX9a18Gv3FKZuuetA0XhNyuslfzKsZv
XERDab4LJs0bqDW8rYabFcTRbmBWu4Nz4lBzVK9GRNC8BHsJi6LAzv/X3yJpVEI/07WNepAGMu4T
l+Ov69dPAPNcuY0uERI4Ig+Fa8ngyx56HOByvQyHflXcJVGuRCOlm5kZ84M711RE1s6vHYKV4npE
eksm26L7KFKs7FiiVerLT3yGnLnkLlWzbR888WMqa5G2lXAUbIo8helZ+f4nO/Iq4zHgJ5tkThzd
3Vu2gPSuAqWu2AP3q4IoGS91ZGI4+6AlwoR0lbUtmYuQpsmQHr1urowVdYnYfWhR7EXChsg9OARb
VVi2b1Zrom9DtBAgd72iH7A5sZ2Be6qpGVw0ZlSo8DTRpNzjLrH21cwLzV/q3i26q93qiGds3cJ3
UyI+7OWJUDJkpBg7gpKr8jqgT5HzEs8p0Lwld5Qd8DuIhipUGHldaEUBRG4tNUad8xSYWG3nZ6wx
x/cJrHJ5gAfEN3NeH+roHdxiq/uL6dWdZ/t9IYY8nyfaiGY8nnZrnW692VHNIy423DY0Y/2DhO9g
NK86HZAPSVlW+LGhPhXhS1chzFia8JLCkYd9vvELyTrv1enoQpylQt2Mn2C9Jv+WxctfBCWU6TqS
XK8PClWMGus6E+noG+7amlhPo9J3l2dbn5Hs/KBvXSNpLBizWXuvDPsU5VO/Qfj60iKma3onwsAv
zi0C+Qer9sMF2c4hNxDAyrMux695Uz1EKZdaG3Osl6qN3hW2EO1PticQiLssXxcaophgVMBVbFDt
VL3o8EVHqbxLJTl44aQ+y5DcM9DP4fzi3AH7ly6PTtpVoztpME2bi7dia2ioetchxoYsU+aVNZdd
7i1GpeN/27gQNvaw2MMAOKK6F/4KU2n/ysA65gCXaZdNGY8NnvmXodaRvBIR0+2s9FXHp0Cr1tkH
acqSCHetjV1DRaQjn4Byccs3HeDpLI03zjcStzqOTpgP7apPiHVx43L+/1HlEWYK2shB8+F/iLxI
sg4jcuvtbmVO5YcFxo79LlSR970CP93xDI66zNSQ2PUywAvdZAJhvRtac61qzNudOZveVk2gKgl+
XGMJ78gLuc6NKfYjdBIKm9NRu1+dNPh7q++15uNkrYrdsB+k7QWU102pH5rEzcLNHKYBy3qMOdw7
qlBNm2Qk6YuaibGyxqe/pbtck7an1XIzGYo42RtuomkWsOIIt3noQF3Ko4kSGks2dcuLifaQh1dF
UWNJ0vbD6eScQpuL0XhygKNcKbt2/2Xjvleuf4OIu+KHy3eRvAe4b5I11qQx4FA79vvDu6AAvM5M
tp6zZ3EPUnfJheVvZOIpbMF+yFQb1MY4gGkFm1sogc77WSd8Og8onRWLvzqdXCDmaISxyTAao4aT
/tZcw/GS5Jzly9Ukd1ebGQ4HGZinjzhxkreYdnC6dQam+sybxbkPMevt3kcR3IKh/1tIUn5VgYhl
0BDXCBj0251KyM3GBVbPLGARicZqC2BYFJlpfCUZIfJCGjLIj0Ofg+qgoKBqDGG3YkEukvVZyPqG
Fgy3gHeAa4IVlGimwPSts9hAMC+LoD0BZbzrKJ7/QOk9dfDdM4DrkWHI6Dfkvga9i5OCBfFcAv+J
bHQIc8MMcEoQGlotM2xU7ynKXHb5XvHStlyMXEK/X2p9ZFfcSUo8Tu+vjbnpTaQQpi+T0N9xzSp7
vvWPlJ6XckA//j+Y4TD1YbZ0BLImBd+IdotDvmAJ/VWrpxVw9rWjREvsAWmy4QjtZvpbFYLHlCjq
Vti3dFaOe6Y6HK16TacFDAvLfYWU4SADud6EL2mh9Owa8z0lS0kH+jJPsiAyyF7oKtt0QcHAL8S+
Ux4t8bPj87sTI3BJ0S2DN3ptThSpeig7R5hSkfwQH/jfYDLPUGNMU2WZ0XZki1+4S3gEHE/xB6nf
PSjY5MekvMxSLhNdGrz0QHi9J7mS6VfvhSMa75DTjsrFKcLM5Wi73YDmJQXG2Q6L0UyCEWPmJhBi
gEMfePYdZS2pxECqlClBTOvhZM+KSL9OoUaGdzBXZ2amOshB//Nqq2B4tZBIps6c7Ch26nolDn2h
YN8dDXAsZElY6MltjCPd0ZopRF+TADVEANYR2UA6JqARz2YDFLdEfkKPP1GQ0glNykiMK0Bg8dPK
byI0LGaLjTdOsbx9vPYGGMcIOQ6hMSh69LWX9ZJ/0UOG8hePnKlPuIjG24e2o6hU5jWKitR5SC0z
+S0Xclw9xGPwbhQ3qEC/aC1E2p9aVnBEJBWim6kkc0U7VWfCx/YD+QxvsCEda3KdC7Lt48kAbnoK
xScGtAOQlcMJuGNoh43mPcdd36kxNNX/NaqdTNvUaxL/tL63wzVwYGO6tJ7CKkYHehpTWW+j1mCO
ajcDvrFDuuWeH/+mFxjsR5X+xEyFvYE8Yei+cSBcCsUxYxj10jcZRLT4zz86JkNSJVGZq3N/iLCu
qiMBzSTkmaWFH5J2k9vPoQQKqdq7HJU5A0zod7HNwCOnLpW4GJVTFxmGKepq6wbGtEt9+VZy8WFO
Bf2Zl7xWWyMHqtWh3gE1jwLLYLdDf0oryHmmY+dg8PRF/jtX7cGUUISrgV4LEOdMPv5VKt7vtX6e
qy1IuFk9t22vwrseYj1NXSSto6l5al0DSg3tRV2r7QMJiBRCogHTcuwn9/zbddpiJHwW6613eIez
Yyh2QqTwsxawWCiANCQlQBzOumQMMyOVcJ/WPkmTCEeVqokjxKDXl2lOX4+X+Zg+v8NA48MtJExd
z4MBRIvXESBcc0MGADwxid29XrTnEorNqT8J6ndy5x1gTJfSJYnP6ARzK5AEXBSkrLTQfELno1yK
LnwzpRZFYUwPkPETcH9z+E1z32A+4ooq0cK3QTRyPpht50IRFp54g+A9YpGTmFqWlUWskHJ/V3Of
a/qy8qpRcZG6bpaLtPJEiX9+/kh16snosnR/u+/Pj8BifzNIi9aJ6wHylz6YTkATbBphwlei4pva
cj8rFPwOQ/0zc1V7WoVUJf2KPKKExLil8n59hKZ17Tn97BnkZzIINaOC9QzQ9RX4ACrDQKNAFTxO
QFFwVvS8x57kqIyTV+XMz91URzeTAKct3RVEMVvZdV9r8LXM8JscfwPW8kJWqR5Wm/h4dPnnfysl
yQEKp/OFg3OZyoyFLDpxwTwH54srY/JfLD8FRpeEoyMk4Pdshj/JghiriM6RTTaPzjJQ6ukWaWW1
oF946Qg66GYqlR71XB4HZwgp15eQDq2kgY8oEhDcz+uXAMM8Ml+G10RaG1i/HCbpiy59dnFLp658
A6xuAPIl6XMJF90ja7BJm5JcscAqLRYaNo5Xe0ItQcGbLx95CP5peg7l6Fu3UEcVIWjElrIFFqDW
ZMFvbZJqnWOwR4Tbnr7IPxkIm67KdF7cfz29Ejp9YcX4igLbGUaMxj4G/Y5TRZzUHebuTLS7XV0y
WFxWvOGj0SvMc3AarVy8jlDgfqVAFbRMCMIIO5fi8vhKaV1oXlMrDM1LyDxiKfBW907mgfHBuDVa
ZXArsj691J5JQjhjoIRHhOfJ7O4u3Va2OEhTGIFddt7X5pN8dtSA+xzRW+3LM8UKQeZKcqytMt+3
yUEnSZylApzMSnFKUxVODmp4SXg7D59A2jb1gMa9WN7iDgCbIbIC5cift124QiyqS+h21frTCa7q
k0Io4jA4wR+Os4ddjXG7dLTMKy+B+SbCm7uBuPv7pxm9cJ7WR4afh4jK8tJC/1kXKxy5a8lcZdJ3
5hsANp3WqVfkXZH6YFNUiPU9GXNfHVZWZqBEXQqZ64QXRF/BEC1OP8ZPnGuR7pT9sU+fOSr7aaRW
CMJssjB3IRWqgGgtpq0VzZuL6cAqWESSCeuIvk/GMbDShL4qLZEQhCc6mD3Rl/LKithgflSKLRB9
Rntz+n5VNVsOdd10HhH4ZzJ0TuFcM0DPZjbORo6qPOFsk0PjEX0IV7Fx8NMDyDzxXyCR5pk08rEj
EdYupxNyHZZeCvqm8UV7Ymz6TAGsQBpJNHOOpc0kuaLnIJ7Xc9erywwxo/Zz4C3W9/vc6t4sAzGc
dKQSST61Yz4ijlzrjA9P33TulqCj0G+E0CBMsJsjx7LC6HKQ1niX/EWD4DsoMCao6W6IPX/zjHcc
A9E4OCkQX7fZSrhO4snwOXZthOxGifwJy75v9wbRG8sAMUWDQvDUkPHyqvzCmKQPZL95SQ561KFd
0pSCoXMp9/ppcBq3g6/moiWMbxHxAzrLcFmo+phXMzX+AaKgC+tztro3hPQ2Movi4P4ZmFyTlEwx
gOrnyU8T4DTGOsH5LkAyoknYn51OSUn3WdNHLl8YM/VZMw0GaqTkUC/jywLR47m7FIZHkfniiIFF
7KHEKe7i1AhXP1eLifJKUIihykuuWXkKh+yIjOO6dlkt78K/KQx+lt11TTtFUQMCfcJnA4euXs5S
o4BAKnBVNFulr9iZ+Toju3vpVIE0mGNgSArwQWiH2s46Wm+n0CeeyeTuUQgbC00FLBMfHTFyICA/
TcblAV57obAFEaOtgumqaLc2c90kxzzI6cUECEyb9eeAArUJfXGx+BAqaUDwlOBWRJDgz/uYTHmG
S2AKbMEQ4QqCWopgMbmUsR/ER6AId6ZLbXtQd7/8jsqFWGhyY7g3CDzZCpjWK+994KhgGMfDBkcS
HJnhd13WLl5p3E/DaMflamonj+RqzjgJkdfr4cBldobw7KAWETOXk1kQMnotBkE0KON+3xWCItEP
yF4kPmloIT4jAO8tPzeHCzpea1PuXxk94tTz1vnf7WRmn59kpj1iD6OogOUHRAw7Qd1GXsjKGdzd
Xg44xkIlyMraWgPeXB0PwYEBU112UbWflRXe2Sg/dVo/7wyIGP2at98lMeiMgNvZ+C45CrVAUbEU
H/Y9tHQ5EWnI5urrSMnTN+CZ08Owz5h6DgM4zx7NLADPSkhZLXEX9inBoG/kj2uYnjCIn2bVwyjZ
/euPPtLUn5t74tHJ6Hu6ncQm5Hjer8c/ADNuHEPs+KRDwF95jjOUSJDYEFufE6+kAbUg+rQGi/tp
Fst/27qFTZlzd4H6TJxHOTVyBOPHyLDksqcye7J6BDDo+OMgwjbsnV7UMILQvWWRxJ9w2s0ePCjM
zCb7Rkp0XYfd2BaALeFdcD4PSM61Bnyn/DNEZ9YhLZGt0+KfCAn6HePXnjxu77cRxI2mf3ZNXKOR
8+5y8KwVBMWEuilzDc/4eqZo3EJP+qF6MHR4rzEsRfQCOm2BdZG6bAoesgCKOTtL7PxytSUx7gsP
FKUghJmcpGlkF8bAbzV40qgGPWRj3mNZxrhUqG3mc8WE65yUSfaoz9W08gtMNHdtiPRGywnz2aLC
jlf5pqc6cdKa6QaxiLYO7YzpHJQ5Kiiwo7lmKWVR84CUQ/AzggbGEs7ElPoa85rs+K5ThU5XC04B
ggBIeaw17GsbRhW+BQJ69AwYRSGMxDuJ5cRpZ+ZLap15quuX7rHiM8irGxzyIueQSa2pHqV2DVPW
SElQYMbgClWdJQQurOq9ZpQg3HfEkNcqP6pVSwZ97El13oHRNpI2APeqz98+B4pzgoAlVPisilI4
WBdtWwXYSkf9dgxTeRa0ibz8qlQXzNGUUjV2Bt60E95tl2E1K4jCjjEzTEHguvNChsgc/gdI/1Vh
KwoqhIurboOKx3Drmrx48NDEvSIzFQZfba4afVJuSqYUY6F3a2l6eOB9qPu7LkFJFDU4h0SV8osW
o6wjHLcmF+CNA/0Od6HMBjL7gg2NyFgMx0+OVXf9UJC5Cqg3PD21+ZzxkvT7/6ksOIbXZmSFcjK6
StG2CPEvYufmkrN5e7gQdabcykNhCVx9yyMRozvRzFNCF9N8vXFRruBuzvrO9JqAJQYL8zDylyT6
yIVwdynX6H4T8O4hxMfFWdUh36DKxPl8ZPBfQUpQ4AiuVY82XrEb9zRfFGUhcdxuYr5K4mZL1Kli
Jl00W1c0mezPjjW6MlYSZVMM6nX7lqYMAXa175k35ldmzyHg+9BIgI0rnzFNIEeNx5aiVCiKF4UB
/sFpCil7TK50pUltR75kGjLsy4ZOX6s36HJm/29XdKcdHN8DDoVKGsyDVTQFMXDWkZ5gOpteDRFW
d28MDmQC5OSBVoZ/fYRsctGTJaez+ztx63IwLcEXNotDZZPB0xAkqm+qPo/QaYMfaOcdSLt4326w
qD59MoJWN0qkLBrFm8dejMP98RmqXs6et0Ieb+R6szxWXrFTmYVXaJKnCiPThxmr971zJjF3eXmU
LV+iBJmbx+Nl+/X+OHPK0qEeNtKUEIWIbpUIRGWPE+QUdpk5nEgoCv54kFAysCi8zUhLX3RIRZrK
hXT7d2t7j4pjX/88vyYO0Ql0B6Eq7Q6iV5CU2gaS9/i76qAj48dxgC0OQbh4ZNzcIUvppPNzvo0V
JLHicqt7AwCeVbSkbBgoTuuQxOSa7NQVKS629bDGla2j7zsWzuvkbSnC6Cy6q9M9joEumqK6mBmt
PszxjBqGw2kHe0wlvwBVbtBNlWdZZn3fN0BvY8WTtC9PYxugIq8kZssP0pxubarpbhOhYy0NVnqd
rwgV5I7jsK6+DT7bDJ+Qkf5+kKmnoeffshaoQAMVFagoGW/mLu4lqgd6kXlLmGNbANJPvOf1yqLx
bVDPPczgSuGS41Pbiy/QlmfW/wvbbw3OXS0zee1pGYyUageAyOLcxAJ9hL6+R5Nys8tHjcuKJiDM
/Pjql1D74kOf70Lz4wijjrGjElhbDAz1Fhj5uhR15P6Axge8HxYM7wvW9Li7JXL234L/rfPoK6EV
cyJJzpltwPdRyXVPwJck/KX3dJ36nfBUFXWMjCleFtiSXMqAeTnf9hXVttpdiQp7NQ52eou6JvsL
wY/7R79C62G21aTBjQtaOQejac0Er+sgqESCV9ABGNJdWPKIwN3TkNP9mBmgekj606BqiUepVLWO
TvSPc178S4Ex9BOM7yU+aU1Lh4cF+5N6zbDlXPj07YOMngHM3lZU3bwB6aYSNQifXFTH0gCjynfm
YdYscierNrItTjxAa+TQ7WUxger2MKptx3YwJtV+txMdSqtRvNctnEQa5rkXTXxtS3GCF/Ef0f7u
SaBTWn3sDWgqjM5bjAv5S+UtSmzbnizoFgsvK5tXYUouiABIRBQFfOkXs0hiu9U+gWixcG+j42BS
I8bAkpCpUfIMhu2T1HlCgqwiJsYnzrr6h0ePqYJxWcw/W8Crw8G9pLElzq8jGMMjMpBCAiyYPzWG
Nt6wZqMTpfGpTEVj3Yo64Hd3rf0XwUq4am0jJkGAXj1s0Mp9ULja1PDo04jZdLTC1ImdA1VR6ilk
YTnryHHgs9OjE1x6F/z5vk5bwnLLmH9u/U93Qu/yZj0L16Cg1lYm76n1QeIrk/OYrISMag0yq9GB
bW/a/XANIxUwxwDOuBrfeumFoL+tYlq3kQqy6JaNG9u4T/TbuqjxdPrq527Df3U6kiV8ubzn7Gvc
N50Z/LCQATqmxSTADwue/Sjblkh5T4FGGnK5V31HpiGC+AhtJL/cWLgYP5piT7OjNkOIOysQNAb6
c2k17yjGPmidT+x5KTivOuZ3bKlBfCuLa7iGoKeM8qS2cXBh7en6+tPbHWqPWi1KkbzpXUFpf8vk
m+WeGFjk7WEU55ousn0jhsdXVvtDSHKwK8/PvHrkfiXrRSIe6PjKtmBHiCOuSyTX4WW71vT+52iy
Yqzd43t6xKyZzdigL+ofEHEYr9GnqJ1HoPtUv1fO5Hx8IT9nCLy/+tJKJ5JUWS1N88VjGESMCsTG
dfBiS1hC3jjm8B63hfe6ro47XEhkEAsso2e+BWCXQ1Y/6WETKvTIEm7iVjb+OX/nqnPUeCqXs/2D
2IOKtUcG8gTZEK6VvlCaClKvHVlAgt8hYALTNctO0W4lkn4WbpflQte3GRRWScFRGFSbtqX3jXJF
fIEU6xptSXFyZnigLf9jjHfqaEbusBlN/hiqaWUX1BKKgIpUfto4Xvt0BxGqNiUck7Scz1Pu+6MT
ziPkpXBe0qhRr2RskBe9RNoHrnuDzuPENzKDLNFp+FSiVMKNlLKNIDwM06Bu2Lppe7nAognBWQv4
E2u2XTWm9+7zEdyBoZ9nl6pu1mwIqEvz8p2ryRKWK2rQZo1JVhL+d3rltzSVTzDhW55QJnDqn7TG
UNgLYtqVZs/KnEg6LbEbyT/NNbhnUjXpkf8fv/39UFvx9p4Ic2vwyKMkQ5+3955ktKcVcQBk8/uI
pVhtWYD7zvALjFuG5mmg2uc1fSuPfzUY/830KwKgs3dph4yGxqivBGGypaAY616jcUIWsf27ml49
yc2HuB5cHj63jXFmguPdPGoaav/Lq4IRCisvpObai2qLzyY0wPiI3WqaFZIRE2fj0Rqjj3acV3UV
WvUYLngZK3hDcA18gVYabA6fig3sJYi96ZAsD8h5gcD5Clx4Yzh8d91ZZSNx2dE7omuC09BsAuh6
h8eqk1Csl8fjcvDSevu9MhW6lZFsJUTvt/4/HfoSgNPPLF8wriewpPgbZF0oaAYvJU3FRCKWSew5
mOyZe6gkmsEo8ht0TXiNFojKZxAU9SjnFbhye5DyyRhs0Ckzz6SytVtgHMM/Lk3IbR0E6FLtTlUb
z9ei4kHytClIttDS3vLqzSCYXmf3rn+jMxjOJYZKjCxd2TzGmhdwboqxhnEm0/NYcDo+VQs0w5K3
bt44Phq5NI7ryCh43cD0QQtakiYbeBbBp0kRks/JaI8lcMMSHSDWWaaCM+i3AXocaTwPVtF7uhd5
yL/eaW2lKd9X8Pic4RpMYlazS39EvgGLHCCAlvijimPlhrlGShUs5LKom5K4OklT07ArXhnhcAQW
I1MzjCPue1MectFJ64P5IF2VaiDqJS0MXgrCwDgdxjmAJyKxDgXzMn7ycbUia5bmS4xoi05hPfwR
1rxRS85u/tKvWNNeCbPX+7xBQU2A6B+YqXzbFP0ssf5TGE9Y9Qrg5gJ/YTU1CPVoYhh7gfABigC2
uqOoboQkMgUo/44R8uT+fS+xnY9hkZbwZU+GPLTzI8bfw46EGBRfQ7TQXn3UinJ+vYYtXj0fp0VB
uB0yRifNu7RHDt5Y51hzpInvNLwpEqB143v0ngca79IUhvSw+eCmZBp7eu8mderpj9dMGuY4z/QT
ZVdj3vTsYYt8wUBHAnrBHfMzOUclBxEuVVoQhdSlD/rjjoy3hfBMy+0rgE43lUlT4c8PrKeih07J
V5kp8qtm1nVLk10jzDj5DyQchBaYKkVOan/E4l8zFUk44fTkRm7vbGbUdVh3sr8VrVvls1BYJBcf
3aqmD8ovgu5bE9E3pBeWI0QIiWoGU+ajR8pbwrNmmh2Ck7pL8gs7ch5CrS55jXXiC/0IRXCSHVvf
NYp/2pbNpzerakb2WG7fhNyp//Ct4uxZQDgAsPH9m8G6XxOV9YMMID+Z04jzuAkJs9kasz9KvT+A
B6w7sbaldyZ27pFdEtX1xPLto2gVjBr4lQ9nog/S+Suu+3fIQH7vy2EnsgYdL4xIC4iyNpP7bgY3
elfRF/XW0lXgHC0RrWSpLMeRZKEgw4zl6fVic/HxdHKofcy67wcx4/adtaNwXaVwwQzCs260oKjp
J6ie8Uf3YqvkqEXP6NuAojCE1xJHtrnGDIictn6DSD9E/xm6KhBFOGKO2qlVFXotXXLxgznEqppb
xYiFFuDJS2e7rCEgl8x/NnzuIxvZPIk3Y2egNt+QeyeHk/VxHxr4udg5tDMO1bZtiSNQTSuz/XYY
a/qSfYgB3ycPP70yCB951QhTQ8Gx+RXsQm1UYhHzRpNpWKWskDBDEOZ2nXhKpJOq2/lzxWSn2UoG
AY3khbXW/2p2rQw3HRgOJxbNBQPJIOsgiJ+igwkYqdZOo4aU4iSjeCyo2XRH+wvbDHzbPpX0wuxn
NawMHeUqDv8XNpsWwXM/Ek7bgEUWOZmlm9M3JjgbbeaGsT4SLb0rzEmj0YVM4E+KEJQb8Ui7c/AO
fA7tte4f85mCnKC9DAqqQZv7FuL7QdpHiq/Ep4witc7sI3ivz3vEXoCmQvw7SeBYk+/sYisOCt6e
LXgxr5AMDoqK8gBRUJ92zebGZKFfD4qF1M5menNuRmtZUFlxFPeiHLjs/b88qRFsJ+mFigeZVlkL
JXyZe+kWCP4dzysr4lglWws9HRxrQ4XeYCm1sBDkE5uEQawOzJyYU3flRZkzPmHeinSF75Sp3d85
c51qtshV5JpZwg+XKdDL6ixvBenGANqubcrmUSMQLQtIF5tcnDnzC1CfQCLev9DG1r00kPkFDgTm
5V2SdkF4Y5VvlEwbRVG2BxeKPJikf8AINw5sLcopBHIkziWxMF7p6x2v9+DkQ+Ut+0VFaGWWH84H
DKFTLkjxPkc6GbxsVAq/5/m30uwT3fAJrd2ltjl0QwyNh4dFQ4AR9jbJpOkWt4jjog/YzHGFARyJ
MqbLyTe1plzLltNRV2CvIO0CzNBzH6VC/7CHVGlpthuyGZTHqQsMKiMbtTBVXaWgElBWZQrfUt9p
R5ZJOjGzPvX7V4aaYRJG+usoBJl9hepcip3+vRJnU/ACKM4sfcAn3xf41NkS0q39dae7W8K0SOxw
ckmXbwFKWgFOAiZVyWx0/vDENtc2VwAYloIUKqXUlXplcrgxwkk37K/fcFJPhzxHFVHArfy996ZV
sQRI6owKSF2i8SCxBH1qvLWaztJsFaFlbDGXYUre5ovfzpoZGdUztc6s5Br3Ruhq/MBqru/JfpEV
4hddGZtH2fmT4lAPOKQ6CN78Sj8i71Im8vpKn423eplps+nYl0HFz1jZc9OYMjW3M3SPkRiPCQdY
Ogiq0CwvrLDnPKpLrBaLrenFLKC4yInRoW49LgNxj+hJpN5LtZiDGBv5s8MJ19Nxwsg7p0VCjCuF
/xVaP45UvqQQS7jNIdok58PnVdoJ25H0R3OO+vuoWrpSSuxJSqU0/JNhxZpFJAdctQbjsHP9tz3F
O6rGeJWzhpF8EvEhKUCKSfKmDlX6V3OvYRC7W2JzCNxQAfV/fm2wo4YTupS6DtH0H4XwrxzJVouU
oKmWRwSyBD/QCkOgSGE4AVAS6I9XLYqBtoe65oJGtgnkOpcsCmdaVf4l+4spnLE7PB8rxbmM60He
LM2R7XGFFivMXCOkDDZ89/82fFKZiB7DONTdrm46Z2anr7QKdxztVMkZ69d92tECL2Bmh2GKJzLe
jb/PazOak7X4LqweeyKYM+JGAQ4liN9JO5ykUDh+B9yhlQ0DsmPcmR8uwva29i7Aaasq4npgA1rG
Fc+7BU1JU6qa2tg5C2+COEw1wxdQeuu8SgXLqc6UV2ifvzoknydhDS0CV1EIy5kE3OoXPfDWp3Jg
fPqCSKuku3s6UjYZjN1oS3R6NUM6FcGm0KQQZDMDdHofuwOz0sFb46bmRZC+m4AGQkPjLpfeU7lK
b/5mGlTerZIGDzW+dWRJAbbIbDgcEuttzunNRuKgeEladJkJ61L6Hpckj3RdNYAq3f3q/IIXrqOp
s232jvvHKlC5ybmePOC8STd/R+wp2hMDSWt+5fZc9lgulq9vArSh2q/8OSgCGdfeEx2EiFYeZVZR
BkaidnlNn51MiPrJfFftZKbxKbyj9LmOUUeqGDUEZD9ru5QSO2GUlDwjOiEhWDmzvyr7qMQkOXfJ
LbfE6Mqjd92JuV9CHt+bAW6YEtk0DNV8Qbl1uFAHnAOQDHw1z3Tf0gII6oFL/JDR2PapEDZv6l//
wEGdAA27P49PSbZoa4T8Wen1muXWuIFMKJQo81ae6/29ya54XsPFloXFt1wvb4ZKincOKDR8L2LT
f6LfUU+7As6FQIcCcyGNFBYs2vIMC35ag+m7o5Bokzvpn8uAfPfWk1EkGqaqitfbsSe7mPRFUMDy
M8Z75l9v0AOi4tee9KwTdah84Wl7pyuJEQEI0W4pgIgqSbPq3HpymjySyYBHq++SsnYdXSW9o2UI
S3mZ73SK7yUDYhz4B6xXxUOhXrGDLV3SgCUPJC+o77i1oc+AnG5Yel8WJU0wpZlxA5XeEigf9evB
+Ftx9IoTPne7FMDF19H8QZqKSAUMxigvwi4MHvHQ9D2Q4Zbxg2MNokb5RCEohtUhpIvQGFlaOSyY
ZfdTWLWpf0OoKUdW6TyfMNRmZnpFA8glx0FOZ1aNv+Faqaks6SbyhfCumtTroeYicPuFBn0C5FCk
tJGR4RVj1NyK8MFsVB9k3hFE2aS9FctYwo4LnC0n0Z1sns1yjk6NF/wSGPWSVpwhVXZmxGkqzls7
qeN9VB+Kbzkor3c0gvn/31ioSXg/lehM8jYaJYsu/XPrgVEy98k13RBNzetAg63yFZAN2CfASDaD
KhrRgBs8ECsczsKvsCB6ln+o2eWfe0n5+8FTFukaIoywsm3y7a5NntsideYrYoc3g06CpMcLJUlL
qosucelFZLkTpsP1UCz0Gpp7xDNh4iiirhd/RxV8iV8rfqu8qThThphBjTBJLsu9UWi0kYWsaXru
tEEIqIjn4FwAdbUXOU4QXPTfsQyX+njxOKHA5p/94lhEc/MHOGpbpUQm4Nd0eLCwAygzCxLu0RRR
M5+DIN2FTlW1p/oiKJMfyzkT5FwU0T7Sh6ePxLye5ouiylakk3yG50DUJqoAeqsBnfx4wDP+HwPY
EoQkFhrbwNCinq+eU2EKBXXb0TydGuxJfS0aORrDTUdm+Cd9X3PW3mBMTIkfqsRMgcWelPILhN9l
r1f66/BtvdZP2DNJmL3xSUBa+OONb2697qRz02nHxdbKs01ST11sHhL9TzOsX4ynexwn3I4WjkKZ
PEpMfV1RWlk4OX/Zc0iOj6aieksjeHsb7ts8TjVMhNXEj+AeOMRuYf1dAdONq7/zgI9rK7hJ76X7
QAG4Q1sHk6uNyI/aMHD1fFVGqu5dS9WOxJDukdSFNksQZXt02tS3oXFvkBQJ6m5i7km1c9Bk68kw
RxNwxcAs45Iv6FHZv3zmqJRq0X878IagGNkziyxDLpR943aYzaH3slzJN+eVtJY5qWGhOb3sPOqZ
5DvgasmxEp9gTv8nNx8k8p9zoaOUkPjXaMEaTOUuQ9dRKktNLcM9Xh1/bRickXMr/G9xwVKh/hEy
PKQ32X2t7l01EI81/b1a9ShXNuffYlZogdMCmjFzeISBxHHTroGbjHsa3I5SKYvcehGEVkqbLPJC
fS8n19AlAdU+utoxjSYHIrlSZxFeAGU2X8s+ApwKGABqJFtzbw2Vlzn9q6s4xOXM2Bp5+LAP1e8f
zZtJYP6TpfNCQnxdiY0XxwugJ5tfehuuYbyt4KUCzXPn+FBHl8a6XzgBc+21ctdzeYP8qNbx5FKo
FDRTP4urCfyc2j3TGeLd/Ex0d3Jyipr/ZmjIPRQx6nK7EZtMSUEyb4PNGdlRIsE1V4it64auX2YZ
8cfqHdHprEwA4YwW0cS/Q6c6ZFpWOcAN0ceX46oJR5kobdi2xqyk/7mfk0MWuQQOXeiNUTDxAn8V
6sUn81AqgPmxMbh+FaRpIFdML4rtzjIi33rPalZ1e1KzhwWp2vRJy00/ospMj+LVofK8QlBGjHNK
fRa3Xb1kTEpPKZA4pV3StTUgzNcgMAuu/55POXXBwPjL+d6h8zeXDlN5vhlvBkCKSFvGON7BtWqd
sjWcyMrz2uGuXtYPi4YNAsqH2wWXPhP6yAt7FOxO/mbfiKpN4ZcK0x5hPeLYgnUmT2E0pAtyJddc
lhnpxoJT919EG+LghwoggyZwOqnA33RVEkpefFDPZKoHsDG7vSbIAJQ/0kRmZzeKmeVb29WzDiiq
mshfOSwHOuYFaPemRi6OKkAJfgxGaJ49nwuv2ypJ8h8UKhgKyRmIS0avC3BoIqSqahSyYrl808K1
pYQIbsN1mAX/erTdiLyGFQXRfGdzURSf318wdq9eQemcreZZwkRCwWWwbUpVSSiTDS2o65Qpibwr
JKhio3FeeKBDO2ZtF/nrWxSKqiB4ZUeNBjeAs3350TGl0H+ldMUw/c21Dv3p359UZOSXR+dVEmQ/
vbj2fZFTPhPWIzwfDk6e3/yaUpTs3/yQR4rZJaEQjU8ulY5q6tk4/LDbhIYR/giMxi7oGMfDrHSZ
BeZVugIF6nmTCWrb++9OoZHtuL4gefpYdN/xyShKOn8ozIh/wRhKqAXE9o4+vlytj8wrS8IfwZuU
VjnpUjUdbcBkTRJVD2RexHbei35KI/1lwuGT9FlnvTvj7NV7Y5Rxjs78wl0/x2qS6Au5Ts28YgHr
xIIjuM4FjT3yO2DUM5ZxdmDeTo5+iWFaBGI5/jfGdvjn/MXKuke0MDjHEGXxEkIXjQqYZkYSpMG0
KSa359MIGNG1AxcZ1aJ41qmEZbycdjLz37HdlwoLub+ur8KT32T3ctKoLflSQ0dAnloR16gKMFx3
e0pPeNWnMXEiV7M2W2AdyyLf0S66PVYgOVl6wk8cr3gJLWRme2IAjejEjvxx5GTJrGQWj21zrEna
0/6uctgM1JTxG0HzUkXKD6ez/D830bBCwNvRETpb+pvacjuwlEYorZ6ZBeD53oe+oTvKCHvLGLg2
/hh+kMsK2Zi1bf2FgXNBl8f7FWfxndS6dYgHQR8rplcISI5Z2dG8V7xFF7E2RPJq3TU0PuIqwHjN
CVV9RFq/fFwLYEkQFpOuxNAL1Lu5eVVKkXHqBXYlxSygLQ8gVY77a3FZk+lq3uHsuO4C7ys0CI1G
FCdment/GbDW8r80b+9k+IEaqh1VkJIfQ/OGZj7gMspINOBAmvLrcFAySuPPQc1jdkxHstVdwDlo
3abHB2+iM4ln8pE3PcchHVd8Tcp/U3lxQ87meT5ZE1m2RA+J8FU2s0BAXtW5wMipo4tmwnbhRMwZ
u499WFVGjww2mRc31vuhwnJGqewsnLIMnDERtOHa+7lWbJ7fRQdEkvwEz3rAQtfpz2ht0d1tMjt3
oPbFfPBxBfmH4AIZ5IZ58GQ3zG/w3wMXPP2Qok9prq4i8+PaAAzQxHar3tW3v5AA9Cd6Sxf7nueu
jDsboYBJvqon8ODFs8KWd8fquaaddXV4nUDsL61NwvR/XDnGfptVV0IAzxq67RpyIvTjz+Tk77tC
ntLgY7MiA7Msoh9HgjwrNZg/olHiJ9HYgI9HKVx6ftwkuq9yCISRc+bQOeFJbqdDueVs1vRtGbI5
pIjuhfxN8EsrmgT3RT9PmnCftioxPnFdIMuQFtRXABhMo6gE9mGv2awchxpv+66/nlTcT72fXxUP
WRW5UPyW1TjZh3knCNa0RkekTeqiMRT/Qs7HVsFAdS4CDGuENjntEb2ao8v8csVjFzq7jRJJNoJb
geh2ms3PvcrXqCMGN5didyor7s2WfMYBV/h4egw0m1iyTiHBqdJ8BBztFST+vdeg5PjfCJp39Wud
DPgRL0BX6bCUEBuMhqaaKr1SLIUavffqqf00GqEnItNf8Kwm30UmlxkQi8aAcccJ+8vTDkrQeWvs
8JHI1yejZsCBWv3XBPPCbmjfvQffi/d5S7dHwTbeZg0ycKX01Qiuba6nubmLVnKWT91av99AGOOf
DcvuifRif0APxkRidH/jKGZn7IP8lCt3J+gU87uOs3MuNTMnlo4BYMp7zKQethPGO3zCru0g0gDF
0dpQIr7VPurENYCuQL9Et36L/NqfC2vGhoB8ifnVQmOkk2byCfs++YJEGnNaPqC8ZKdQkYoxvy8t
lgJ+6zZVl1FZq1r1Kgw6pleA8cy0lDDnlHGDsDp9lpd8dtToVp297XjbGwu09+aX9T7nb+e8Ubsx
zfGmPhMnrCpHnM/ly9GRRx7Hm/25XHm1GZstKBrSHDDfaWdGUpzCIWSTTP2AnLuHUbEcY+mS/oCJ
InkxYSgnuzXIGFQCzydBm1UXs8596/vDnoEwDFEPRI5SgfNWPCbAWZluKNaUv+C3FDMfTiSd0/Hq
u7p3DaLpT2amR6YAB/vebg9uAM7bR87gfM+kdNEYg0Z8kiyIa7JPcUbMecs6dynOgoLS8XjNDjxO
l7VYoUoj70v27nZt22N35QdsKXPlOUNRhEUfBbFe2xo5XDfXLOtptrvP0yhoL3uSp0fYaLdqS385
FsGvTJpBYKebCJJJM3wAnbDzxACaA6rgC6O/XkzeROwqxPqZaeKvLJA6HyFmJo3lhLc4SASgbBnn
+eMTcyh66yHfnFZ2O3/5HARJyYUjH8WUNc6q2xnNB/ofVDKPTqwhnST1wFbkjc3AfvZbscYmij9o
n/KpspOn+wjjHpGeU06uGWnTytVXvd+Ov0FS2otbDOmo980OjPrP3l2Rg6oZDxXi6z9NFKRUNFcd
0CxJUX+2YD5FC6yCx9DFOFzNgjvRiutWFuCtn1jZul/PtQszkl2PS7TeMA0GH8f1a6bDXh/yeJtO
FFD9bGbx0ubisBkKL/cJnlSRHa0VthRjmU1IeUYI8UZY/cJfOQ63yE9zcjKt9kQyhUkmKMlYVgjf
G3t48QH0nT6InD22oZ1CYSjC3mg3+pY35MlLO92VquVPWeZccgIjOIp+so96GzOHM4+RLzULiduf
R69aNciBwyVDdzVVHGkAjkyd0Kl0dSLca9P8RyZ9ywj8R/Ntm2EthxbUPIKOBTaLl/QkVUPp/Yaq
XUbFyf3EYYIkfuVjzxgxWSJ00X7j2CWk2oAKPa85SSPJugGWcqagmOiLng8On8rIbjqhhRcu2Y0I
Ef5yJzPQC6fQNHkZB3x9WqgGfST08F1gVsnqjhbxU+XrIZNPwfoz+IP8dk9Mp+HnMz9UamApfTgV
gH8u2iVh5qjsy9uisxvlQ6J5uANmsqHkaS9EwuIQcgyVWgOQW+KBKYli726fxrL6KMj/xIamYwml
3DUrttMXBWf5tnR90lrTuKFKAWrZIKmZMlusR0PnGwxOBzTBE4n9aScuvV52fibFddal1PG1C8FJ
n4wpPnClpWf44f0wluSXPhaoNIxr1pE+ReRIzKT3MC/7IZnahK5CzMTID2rXnIkdZDFGLCybJmr7
flfHlQ1fVNH92/JH/AmpfNwajbQ6FsXopY0BTmGshAg0XFVE3CKpx5MMQoHMAqROlbnUniS5wsRO
yp7+vdbo/iRq9sDTfsNy6mueCOQF+I9ZzWGdZ6eVn2fQ4lhxmMFUfjXDMewQi0Ul0qSzFEsmUJKH
SH3L8Dp8HMOexma7kYb58FOkVbsLpy987oB4FTanudkXdUaNNjQRr8iQsRaDp2m0Zess0zeAqz7M
r5wMEQDhwGsb/vJvxd4Gz9wc+lxDri23wYV/cuZJDvI+8rASwJt5bk4vVlgEDVXogUrJo0siWEVz
JfQJlbWPtziAcev+Bl0aIZFDSUFftJ1wLlyIsQdvs1Xh5YuhuCUuwI7Vwd8QMJbi8h+ylAK28/vW
9M7KhXEZqvFzJuw2psIiioi3+xsLRgT00dkg5HTqzDCQw39Pfh9063BuqtRcbgE06h98m7lO
`pragma protect end_protected
