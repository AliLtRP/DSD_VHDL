// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:37:17 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
nAj7rUPZf6H9v52VkVOa+4/rS374Of5mwGSu4WWhc7JykOK1RIUHrupwpgHRK4Ls
UZqYMbvOPHLr6OmQoSWUkk+v+sRgnIhzlmBxcPBFYlO8U4lz0f7KYuMUSMDOYBmw
Arit6vPvWXzXe1dIrLYqkDa3CiwhMQGH69+ofc/GzWY=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 10080)
vB7ZDWCtmZypel089IDW2/rQFCXH11duuS6ocMYvGlN29RUE5hY9MjDqCmVOoHci
22mH+M3BMEO2i9tD+6X67lttpKHbAwoUavGOgVxpNjxv+bCJOC3WtjgOkOxv6j+X
Pvn6JpxS8coMZqX+tXTffZIg9AUuAXsqkRxxMT3vNw5HhnaV//blP1VMyWbSEi0U
RPa0Ip+23Fgnh/5McwkVKa/AVZiB2LYXGUZajXv8vBeJ7fHjCVUiUkJKsEXw/Iel
nc849YT1O+0Rkp6auEM3xFROvw4nf+0UAL2k4wNfKmOpyIlvfUFuITlcRlOiwFZ/
X1KgB8wJgHtNsci94vvw90xT3iXO5ZguELFmrNp3cB4Jsfq4spYGqDgA7xheMxrB
M5QrglN4l6udFVUwQ/R2mIHK2uA/JypvJ07PSAlM9ofJj3CLShn3xv6q9BRLUEtI
TheeTwAKTh5jomRj8/s4opMNFCJYXEfFwDNhXYEsZoGbzpjWo55qC/iUTB3nwKYv
uPpJ520hKwB7OlJMrpZJj4fu61EJDo1rMSJDr2jh8SpkXsUh4XYpk7T/HUDOTaaL
OGov4XV3zuFOuW1q15fRAq1pmmRR5tf+af11vT+7HYpBosRZi3aA+PF6fxkPB9ql
U7RDts4ykayYxC4Jd+EMX8PFDJSlryF3wC6f0lxsnq6DHHyMklLf75M/PxBVEj8g
WCp9RJk5+h6BpC4le2b7RZ3K90RP8XI4vitiz1zNAJKZXj7wvSrItlsYzVIJbeLO
eXsFKcZDbt3zQmf8JcGdiPgbMcpJEfS79knDH1ZJjRV/AKNYShLT60P44Vx244kS
6A6StlEbEzgG4w+HQuY7RQIWYtK6PpJ0XZ3z4iCdN0JCe5wXI+oSXazC57/+1KtV
nxVVboTz8RwQX0wNjaAXzJ6Ex3xAHMtoQZX6IGo98Nuhe98r48M5BUHnxqUm6FtY
TvCVRFcSVqGvKZAFVc9nGlpCjeJMGNK8JjMW0ZYHXnXu0RqqcLSGWXscBfCai0y8
jUllxoUYTef7rWekR2dznF24J3yHEpbqTxpWtJD79oBNXWjkl8xIvNDe/SabnTrJ
pGafucveAP1yrSBxSWBkN8tlxLUu7B7R6aBVxxQj9Q6sNyvI/v2KguYXVas6D3Si
ZUXsS8XbalAU7iIkeU53h7tuzd2fkim9EIPFk7eCkJPrxEYDqiG70yL4pRxrg2Km
MVGJE5+iCtcbp/W9XZ+NGpcy/FwDGiQHYU7F/0b9OZiI0kjsyvZCoIM39aqPwcgC
Uske1XYLz9+Rck8Y98H+258CIGJWijFgJsNEojAPjVPBkwaiBkNua5axmNEV3Y8z
4EcF3Ar+3qQBTWaEfYv0kdprQltWahzx4QHMY3VR166RGXsn15ae4zgZ1FaolhvW
inHoMb/sNiliebkKBQjAzTWOj1gTW5Jq4PnjwDUsc81XLa4NdY+MVLE4FQ4xM6Y8
jU6+N2Bi0QoBiZHzc3K1iqVuMYW+LDq8FYyQFPJ4RLKosc+fPBNkEy46FAhsWPfE
QmcePkJVIJcQZegJ+u2AmACjVyHVennikYydbBnGioJ9IDieAkGg4VZsa7dyexgT
5MsWbDmQ5JTsuupSJYmW1CqtKHgY4Xg5j9BehWOYdaNrFz7KJ6Ucz0HuZlXD7fSZ
FAu0T8dKFFpuCdvosql2V1T0XLhEVVFX02PAPr6evm6y82NZrh5AzCfOxgWlDIz2
gHFH3XDBVz39kpaUO97ayJm25q3EDwaMBfzqmozvMMWLeJ0JWfl1AyAcgZ58CTJG
U0cUKilVjoiu9p0GslBo+3d6zFWZbFVImTUu6m6MC/bPONDZwmxtpvjKj0IGaaJs
uiLIeIXMgMG3IX3GYBKXtfPdIWGp7UyPORL8dp/Sc1XlejQjOjugzzPnnoxOUenJ
1GSgNftwFI5lqFEL+ZOQUqTRWE/43/71sORV1AOvtDdUyP+3aqUL6EDMbtb8fpgE
2BanPmN4G7YPtYsbXesMPxKfzQBt64+2Gl4UkfoBfe6neoQeAlLvUOiar87QbTWq
weplWG6lre8TW+nrGgIOejw571q/1jKNr7NqyCJkEVO2Nzy0RSxZsWmeTC9DGBk5
7veUM+gQlhaH9cbpWTRtTTuHF5OLlXjC7OXGL5SkISVjCxhK7BkdRkQHK/uA1B0d
dFqP2FjbaU5LbRy58sUeFlHzTl8FhVPqboqcPXA+jzT+vzKNiG1CTX8wlbxZRrvH
EjAx+G31UWxjY0tzP/KPadEZ/6P4uElzey48uBoWSGu5Ytmn42hFTT+7votNRRg0
zAzIaJiiBolUz/vdMgWzJsjgpqGEfNmzJcoYYj1V57Fj4uv1h48phf/2MuKGgS2Z
P/y+OT98ZcF2LfaB+JEqxJDLcpNimvoOyRYrpFWkCi6ZjtnbPt3JTE9AJBTuY0Yq
8rMU7B2tCtPMc6ZYztPWwoDJdLT+BZPxkGMnAyTjqV5ZQb5PjY8sn/nCg0x1uay3
TnYxUYLGNTqEEjUbDEiHxKrqdZ51hSob+myDxrTjc9qZWminsKsvVSacWz8R1vlj
HY5fEnRQxdW5NRYaNE+z77EN6t2x3xvIBiXH/mb8enODz2vBhxEraeNc2js+r/Ko
+3m3C1IPxh2Of7V1LxLcYzIaW2olN/EpDJIOdHVyaOY3SfOPhj/YMwccGD9nn95O
GCSMv3zjeDNeCHUScRTgnq2SMEGxKRf9kPDmpdXZIhH2GJi4Tko7ZuPqFh1BfqqG
xhODswmBruuyMBsycornOy9iP2eoT/aXsDZkjmkXgSnrtiL5rdQR3c9mrgUwvMlB
kcmdZtF1LNPfXlgpUs6E1sukf7UTd6dIxdDO/Gi/AYmGdTjODAKz7vF2Yl2/Uj/1
Tmahy9t2Xx2bFfsPTbShDZXu8Yt0YgRnlr0y/vdlr79tywvZox336JUNQyNtnSRj
Pqf01mCTcTUxlkxnsu7hVTj1Lvx8V6bdLwGYaePPV1hIkEY2e7+z/xxFi5JYIAl3
P0EJJGA5EfFbPUiDhNDGnImuGvmZxTBwo9bupfEkhkzkjJm8Lb8uN/z8tt4iUfz6
53qFKEU+8wQeGaMwL4O16dhYsr7C5Y0Eoz9+uUsLEgHaigey5Pfol54kE0jpBub8
pQaGXRgOg/KTZwkDPQNVaK/3O3liPal7x9xsACWte+OyAydkRq79SSGRMfw+xuza
AOWQHg47Idlw0AhGd59CdhIetEKiH6Naqh1zsKGpl2SQ3NOkY+rtp+TReaLt3GGa
laDO47Q3IS6iAgIrCCQ31nArE0cOF4rsB5zJ8Mxw7kaWY/KljWRXEfIN1VLp8Zj1
EupKu30dMAFBMg1JS8oZXpEi4m+6owKArIbJ+ehE9c3IYaaP1VCtMowwI/hZcEfp
ug9lsWQ4FBH9VrT07DnpJdAVxuNtgnN2/ivtUp4nleQQueTj/GXvCMTtlthAAbz+
G0nSNB1xGwi72IaELoSKQjoZ5XeqMkVnzXA/mAGQbpeCVImpAOhzDpfIcwd/5PAS
Dz25XlVbSMpdNqrokO0+grqv8/G2m3Y6BZ2Hnox4C+xYbzHCxBsrxobGUJwDwRho
RMNR9EB5lehKQzfStwg6Zb6rE8c+hoRHObengomv//lE8PnhFdC1Pjp2csumR21f
++Y5FSDQ9h1RljfeSmEItgQvHRE8H+OxtAg+4qepWCwGh1bAmcPJVzUMIvLHB45O
NJiGpI0pyWjgPFsTWktaokSTvWavIksFfNyFAZ9xVt3uwnT8Sa3vni9hkwyllW1T
hG/ukyXo5lIv+vtKZqSZqTz2VqZlyv41NBqSej/Dt3WGxFiqbXWcaVnxMEklDEEz
WhhXkaT0Z5ByIO2PIOemV8THF+OPRv0GF5BN9r5z9kv15NRsLclxkekyib9Zl2Xc
+WTdNDibSTch6ynYdOBZJQoF2qO8QVr3ht/bnJo9VnWFUKx8vLPhdVjPO6gU5nN4
OFiguuqP+k88FcJBHInctSxuBaPICG6VKFiPL6qrwpPFL2ljLZCGuWIHc7nOawWf
IPsimgTPhmFDOcucDoLDKS64k8kX8UXDm8P8ETLglvK7YUWK/Rskj6nKnNUhtHok
ZyExroE+B7DmaH5ojfqiNCDyeo7fEY1/0epP1AdIdYVJo0ay5w20Dn6ps7+6Y/8b
dVmtY3f0IfrYljr06tzxHDot4aKvR4FndAHr0usgrewRrXSX8fIq1PetTxSNMCPI
dnISmQ1BkOmKP2z218TqeR2QrHwhcBBsVX189Cp3R4WZ4bJH9aN/qnjv5vvOfxF9
pDp2MfE4K7XqMBEiNTtA1fWwoExRMV+tg+bHj0SUZcBovl/LjFNi7DsuifggLB5y
1onSiW38lNARxiy1bTbb+m3pRLQNsyWj6lVaINRaCJjQcqsGHUdSCqmMKrO6N4qw
jihhvxR2ULOFnbugk7yWB3oTR8L9PhIdJQYD1s8SyjvKR4ZZCwUgqRuIB8MtPbRB
BqZLeShD2TEPAFzsN8RMRAuXdSPDIanUd03du/ihpKo8bh3ROjxQagD1XGeHmzUa
mIgtFqE82qQ2ZftJzx8boHZX2b+en6IQVqHqALvtiLamtAzR4aZ3ocWeLLZ40NLD
4/a4LLZzfmxM1BRv19I9ZcIyZAAm0A0aCxq3fWn1uGJlre/dO6DYRPHxvFWE1alb
Lh3xPZYoX+monrt70LLqLNFOFFW2An/WnHyYkEzMu3hJC+hHYR7UO4cLBX5X13g+
erMWXQgRWTmuU369O5IlBpvTx7jP5X4zpVLDaqAfNi4JjYifmiNx8vKFRe4AeKN4
+2qMUfXseu6E2PKtiX0biQ6Pkob0sQ0T0BSY4mgmNXsc/UyREY66rWg1/Gbyf20J
d2KzfUbVKjQNbIksQrhvG6i6xLKKfl2Sg4Jb6EKvmckpjtreYYsj0PIwJBjhyHkU
OnE8FfjMNm3uQaLFDQcYnn0ZwO83SS6PvqyWedqgHO5JpavhZJorOPksg5Lp7Z88
Z3yPGEuSWe20CG7TbErg9aUzQoWKohtOVFEV6tNpx7ZGezNR/1qEEkXuy82AITou
fqhEtDfgPQ6pHkT++vOd7aBE8dNBJdlCXDAN4zHJ0IeZLbtmOL2xe3YrtF0pUHtB
nA0drjBlax8TcLSz7q4epIx24B1Uh6rpvJfMzFQyAboUf7j3V1ToY1dKKdfD3zcu
/2jThq+sFS2axNAobFtk7V5Dp1MTL5GnFH02GuCPLXscBQaehEcBN0nLTiCtUJh/
IeCwLMpDgKzapK855XPwVbSfgl10Dma66aDXHCsJ/y0ybk/Dx93uF6D/m0AZ8HSj
/ohRW1eOoICOy3G4zZfHwVkjbEwgUiFtxXBiazSW3x0AMLeru8tpOMfL0qo6h9up
nPsvy3JOYyWb5WcjJj737ceVpjIz/tIgjvDxAQoRWf+xGwWGv5EA/j3GvBEr2nxc
8I+YVkPK6lJuVYx6rr4BvR877lMHom0elgOLCjPzg1DZ+w7O1XrGnsMj2tnqaLjj
jZVjujFRb0xORgeVx2iPWkub85iDrmVL4QdkvosqEWOhmv7vGbJuJe0eMYViA44+
4gjdnWEDqaaSajuqwDruvJVdhud6LOavs+FUieiAM2wzKH5rRHUEGcJdH1Ie0HpI
PA3bJWeqZy7oRxBvbnAR5+Hh5B1S6X8lLuDJP+q206+Vkdk5jW3JY1iHdn7Hvy9R
vW7abtZiGoXTtwYj49KdqhR3+0j055NpMLRQCfZatv/HNPVMJrmFsTwVqufld9rm
JrWUVg9T56kp3C2wKcpcUnH5x3w+LPTzD5ipo+XicC+rq0uoKNJydk9ubCJr3bk/
fcawLUHyMEPCJKZ+lel6Fup/0yQqdyIejiYEqzNaGUBDXaXG0OPcHrieK31op665
59onByitj+bOlbNvlhFVF+YV6cP7t6D+9a11tPTfZIhFZXF3y2QjHcidi9n4qufz
MkW/7k6d0tyMhkH8kgckuynhaoHfqanszOhb1TfkE94hQCTzyTcx1mwWBpI/Fkvu
Y/QGGzoD+CM5Lr3w8evCu9H2HfUXWQ5mHeUMLJzzgjPI9YF1uSykj1CA5BQYeQF3
Hh+72LyvI3PMt+eot5Y84NAGCFJ8wro7ZXeH707+sdLnf/qrU90ynMlJeb714+M+
8G5MWm+PEfgn0N5kTNgvsBV/4sAB6w48BsGwJKG+Q3sIGboEqjAoS5W9oJm7snJR
1+vPNlecO/H81c2HWzllX8+pirBGC9GELjCDTtDjs61VJGAu3S825HyhPZap7cBp
85uut88megRk8vx3cAm1CRLF84UydkPQIqqy10v53NSag3ffp3gTk1KyF/U1ARRN
AlDTi4yd+UxNjXO0gmvwdZR2bVRq/lN607TCxaLfvjnGAzlLuVGnOAdLmXLciycS
nex9lWLpNrj8+ENk+DfOBBZZm+1gObb8GWbpxmju5HdMHLXUUmLgSs4ponEZOTuI
BZY69p5GRk297R4Q5Mf43Zd4nWivIXWmChsZMMT1kBJD3oz6lMZ3+XhSzsdqmZ5l
cKc0XER4zdP8VtRYdIn2jOhbMIJGIFSPpHpjR4MxuwIu54eH0MuENlNCbIoip1+3
UgN1tm82CUbbFaLl4iYm9S8Y5lGs9jCYRxaim7REm5++q+p2u+foxhz7x8yX1e/+
nvnZCD9s6l5LGdlWRom+Y3doQaHt4LJ1lQpsWXSlcwCqjRCTEx0tFiWczGemA/3t
hmf5ArsIfuo6rrP7Yg9a3snQrm9A4zVOrC1I2Q5sLFFawXPwOQZUA+CPkKDF2lUm
scSU3KzCJABePk01zXC/9sOuUQ/3mEDu6U1/kWrAP5Ql+vR+XWSNU/KCBRxuMYt1
XsZjzFdfhE4CNYQKNe0TAqsHY7aPw7Gz2vcYEHIZWnoIirp5pE90i2ygXQkl+gHV
dl+wazUnl6Kb5eW4oeTHheKlehuhq92B8ihCK2b1dkFv6VbiurWBMQTHiH8gJhw2
hcgRZCKtfAh59+igPYtU5N1LHUDIzLvVzFkF3SU/JYoNPA2vB2ARueNrxVTBf5K4
FaVzYRXvvOmeQXmfRADqQYLHCcmN3IgER8O2xupmLO1M2U6sb+90a9uqAAbxrzJt
ind/pqLdeUBGwCMTU2iQ4LnYTD8APGLr9r+wuUlAq9WV5Kd8IX8//VxL665S3WKF
Belk3rPJmU3WF1Ss4beRELgwt4sDA9DgbVTuonkCw0AYNhrioGOSWyzumj4CLS9K
2tixJMrHai9P071v6N5w/U5KAvWPy9bDg92HSQG6JIlTdYavebKb5raSh3kYVZtU
H7pblJpsXO9/qUeCSKs99B/3RMtdEsOdDkCfMjn/sIavvx9yKGt8tMCQ8wYNZF5Q
rnOzIb8UkcWWevG9HZr68Cx2+xCnfVFw/CgbyTXTbcBhJ5IhAJxeu0yymqvjOp5p
TMs7e5h3Dj49kCnFZD9uYg6Y0wHEj5mz195oze81bbIsyq+VA6iGqmgVrYpzw8Qh
qj6lFyfzZx9jArwKR9TgZcCHNsumFM0MufKFkbcxvUaZ3SeKALQ2+gTZHDlgqu2h
FmFEMFgyXg8MIPBhltZsZYuAN0sx9UTwatLBOQcBTfIp+Wt5CAerWfJ1S5XdPG3G
cwvQN8+KwCN8mI3/TsTe4uEv8tpz1tG2eYQ0IpPsK3+bbggz0s/X0YXAulwWjMjk
oSwwaE/1r3WUC8ClUWt+smG/+FT/+J6ncJrBwE6o9HYG11EZq3gEEoEyb/njaixI
g0fan+jjRPsr4w6XYg015ZWtFlUYswSOOBdTXyUVIfgmzlUX7CdzK9Z7+iF3dNi0
/5ydRC+FOEIIx7JKS0//MUCPBGIt/hDkTQ3AD0vTXd83UxiD0OCA0SmoJDxwYU9L
jJ4TDTVCEFIlTQ/8bhg+u0XtmdTdbLRjVEtcg/3oZZeFQFZs5Mj2keXp1QPvBDnF
+tPVynekSKbhuH68bVZWmBelET5CFThmmi7zsuurnYrS8AvXFBgHQuOjPKLyrACz
xBoZ+zDvKBhQE2QP54PdgrsdDT5LGTjJbhWH12j3RDQVidhib4yg74qe/C8hNUJy
s50/29LJoFl/TroY1Q59VwvsnvQB/XzpkM+bAuVp9tnkNZva8yuHTIp7hTX9TPmi
iOol3X818+74QrIxOVfzLBkAcDopuj29bp/qi42cA28oBAzNj+zXo1px32awX6cW
7LfQfHTHFfEjIureEBGV0hAAqz6egWS/I3wTOM2Kap41bESX9wTVtQZTlTFyv8X4
TViJEQt8Tz/3tXt8QYVe9G6eGIGeFOLH6uVX4VUE6i76UjvNhPS5M7vlKPtn/Ls2
SZJ6/hDvRJO19Rpt+0sEv0Ah/nvMyUEjqk7bPeQhd7A+bzIqAdV0SqTPiaO5zwJK
Wjs8o3nDuq6F38ZbUu0/g+L8P6VeKlVbAhODTW3AMbABtM0NIG0PIax5COr9acVf
72Ev85LmGYDQqqvXY3Yh5tD42NB36jEZ+Gob3JlA1HXrUuPfQDSDEWwxI6xStcgv
8zjliMOhII3dfI+UMXWtiEHnc1z79auwawc8JplkqjE51n62SQlyyiF59M0ehyDS
Zb4AKFrv+3RqalcF49QYdOyIlOCvCXHRZQEypTuDjNqn7Fq34qEd6FYRGs6niN3b
4Kk1uPD1r6FzKpJpIJpQGRwYLgUSR8DbhbMcdZQRPZq71A2UUGW4VNS8RhJO2a+n
rrVZdqJ/uBed6Ls5iA0xVjCj2Mf04i1bGlNZ6lzcTKiT6GWDYBXwUTPchJkcZ/Ee
6q2hRPHvWp7i72MM9b4AJrq9qNfKYVg/xky53WbCpZIhlbDY2xZBhmRWpppioCFE
VjoXu+PiIbyzf+myJgzeRUL9Y6pZRbi3AxnucETgWHhWPteSZ11Jix8zGpKoA//v
JUol2VRzAlAqPnXD0fP61hptCYOquE3NCP+9yjhYIVu3k747br9Ee8dLM5m0yarb
KKVm4V4afHYL5P1UGLjr9gpVZfZHIULEozB0yub4zJbvCDq+MiXUYjFQsjDvF/YK
Y0CUoUVsxIlCgKuqAGPcFnbWytPBqgQbZjbFTzhczCuUDZzTJgj6DT2G3wkE2mtA
X4YBUyBd28TfUP30Pz45p6DHbu2JMLUhQYKKOcNryFVKoTbCSeLJ5qf2yaHhSW3A
tp/z37YGABv/dHbVC3hllC/ospy0arO3x0NHuA1SgR/iDKh1dt6A/oHGUXRFRbdz
6s+CLJvSOQdB/GepBQQqoRyxbEa4VTnwgYJzpa9OpV0ctqUorqNUH1zZHHXiA9Eb
ZX+n4ChtlMofs8Lefvj4QilBuulDFf/fC36mds7ghJUcLZ7cMIZu8RQT9i9y3D8j
wMFL61eGBguKp+amqSpyJZL2vS5med7m6tEiiQ4wTAhq9McwVtld254U0sBGXIvR
IQlvhEKekP2gXCRinCF12jK70hjeGSdU+wbQvJozRJKVObwGDB0nLhTIi8AQRxKj
g5KlzJeBgX1GI/tO2jU0DGCei46wVSz83zEcYaTP4/Q5qurjaKbza8Qvx8W69bgN
H+bKZReciCLJ3qZpq13My3cT4GYspZaIVsD66Ql/z2wEHcXOtRuz/iesDVEQn3vi
Waj3AGebsir8XbZhz8eaYQaATl94dCKZimiFfgzBWxqllCDiWRu+mpeqaTS9YYTW
NLBVqPUUOJij7tWQTQO1tRizPO2fO11OL1ULJWPuSPLFmjI0AjVCyCG0utVcith1
rYsEC++oAwfzejsvlnNSz68nOetGqqY8WN7QAaX/Q9bxXCAmdwmZ8yOLKUTRp+sG
hHvMbM1GCQSFgJsYK8kZ/E5sRzJj/2ddGzFkRbXJE/0eJcJgQXiFw2iX/KdMy+75
l96u0RUeCD0Thbfy5epC8OWKGo45UC5BvWjR+eFY2Dk13ufoPTUPoMhn6r1OVLTP
WP0+n544Kk0xDdrEdzHrSxcR9mkAnqzUounw8ZB2dxAZsTChrdymlwPIG3AXvjWT
/p1Ng9HHT2qBZOv5kcZGv7G4/qzt5Cf+v1Z+qN8wVpNppUW0UbxiaeXTf8o/uHhI
cstwV8PXHS2PJrmCBBknJs9YKkoOYb2H8saj+jq8fSrP5PmtLtITWt2FKMJGXiOP
ViUwIU7W0IpL784dkwk2CY+9pz4uHhwjsKxPoRQ5qIWuH7cwZs25EGGPx2yEaXpX
soIqjBtaksmenbnMJV0cgvBezegT0zQeEQRf2YgFPUxEAT95CvRJsfZ9KMMh2scp
onzaFOCgcuBI6cg4cQhWVpgZnsemdsMce4XOwBgYiV4AkN3EnIt7vbMg3dMOG8AH
cwvKwLThHDlxKiCgi8ZxNwV5igL4GqRL4TqUsSUyrYjqyIDn/QWtsIvE7En1CiMQ
l6y04jlJiLCsB10kk+CE9noQf3n35ZuRQhP0FrCg4y3N8AouGoS5wj8SCfUMv9yv
CeENWOCdCj2hi4SzY92hXj4CDkW6Sijjosg9st8gTfjrDsDNyuzkAsGxZZ+AMpUy
x2sA67lEFRutDQmQUDZOy6cqyB5L+YxJOI0jDtqFWRKWtT9ZV5Q48mEOY5pFc7xS
8zKPAV4dKl8qVgRW+z+N9k+8gwqJ0bDdXqTG8RzkrtVJUQ+sS7AynI1PXI0bL9kw
bxF+iJuhM0X2lKhYVV1y6NwU35Swj6fYOzfu5q1UMhqKq7EKjVR/ApRqKQv1hJ0X
k88t5EMqtngRHwHf7JJn0vEiiTecVYlWKbqYK+xibaiog3Zug/0KOgE8EY/y46fj
fsqlNkB9KhLOD8RR6btD1cA+rfLJlIYUlS3RDLKVLs7aXxuaVrMdaZGtEiVg4EpI
7rENR7BPBrmoeQQRcptCqWZdCVhlGWBhtLm0vkwJBSOt3KYpy6Suju78dP/qkw1O
bGISowhGJ0gCIzOAFSre7svNZKlJKwTD1wY34G+SKIc1gxmQ1PuUefzbPQJdyqxQ
jhPnzC4hDfLQ9F9hWdhBdLhxAQI1LIRA/PdjuGcpRqn+EO0ucHo1PYJuwN6TpKN1
MdwLCdHdzzWt0Sb7gVfjV1Uf7NAANpNttrxlZ+kve08kh2esOf46bYHsJtazpj0K
O1r6tX9VdiagFGB+H9gFwCFKckuWuIGHfR+/bnmCsV2Kg5NxFQYBGX+SN/EWWrV1
+tr3womHFzqMY3RgyZdFI5PpN2PtObPQYxkUJr0Hp3xWOjFm1vMWSZ3UnaOVGtZe
UBGQKPjJWVgN3/guGfaJxjYyIFovPC0hFOJlZtxzPzry6MfiiP+5Ls0pzHReqyhp
+trUqKscq0UwAtsF3d1u7l5Lc2hwsv1vup+cmRv0Ctr36HjcVOEVPBTKAKGXItAg
ENvCNStHovwFMn0Ty3pqUgWqWSf75m//6O6JJ4UHbRmqc6sE6ABBc0XsncSvugx0
Vt5rwyt4m4A7RyFCTNAXBpplJl7iaLb1fvhw8I0110VWxbgfx422ypqTI2zmQKI6
6PBDA/EMUAp5oodFXf7zGz6Qq3jU+9AZnnGhAjMa0mqJyB8arMhSLKa4M/jpoptR
RAvKKyg8CeCT95zg60XgM0+cqaSEonBfVCpPzN/pOOZoASrDN8Ev7gdQIR3M+wJf
wlQ030oXQCfjFxISCKRmcjnA9kJ8LBc//05SXWlcbWYi+p+QGQfiE8Os9sw0+JLT
E9YlBdBQb727oUkZ0FQp1IfgTRrrRZoNs0tTxOt6WkoBrt01/iDtB39lsA2qENzt
vWfQnG35NSgPBv798jkFw6h9Z2028nlFh80zJdObksVw+5lwZ95dIxvWCRg3zcKX
LBbc+Y+7WDDKvpnpIB4jqOtSBc5cRX1apggQH0FGfmpY6UwtdjLbM0G9W0IEmS87
iSjgqoDt7cUc1+rs4pkp/HnqeiVgCoweLG65LBzBJvjM0k9oMnFI9YXA8a9AzlQT
VCVRPApItpgLYcS4BUFOqhuQc3V+yZpND6YuR0WCqe8CLpFpOIjEwu3TynRzdfqL
SUh6EZotyty9/kb3OtQmMaW6ZrSgoE1Ppd1icOnOrKO5ZVjxbH/GMKvgeBDvh1m2
WFt86Z82Yr5i7eF8LuKHEjozqwl4WkYxRUX/ORNSEhHXfrW2o9gqAj7Src93wIZM
rsD0jh4At9rxETPYHv92Lf0b5mD6QxIGXcXMecBKsjh7FXUT/gUduKuMrT9N+F4P
7GUE8xsk96s7cwEGlNkUvWLRfBRbJy1Nt20ZgiJOHVd6K5tGJBI6/paiC54jallc
65FTyO2x9nhKUS091rgXq9Vg2EFB0WHvoaHg3of9ldrDaNSes/tMUxLx/diRz563
vFyjHt6o5b8aWVkHdj/SBOUVWqRBHYWlNOGmUWbcUdFaziZgfyeU52uo0ljFseY/
wsJSD1u7rDNabdoFG1FcLsJ0v4NO4f+Um5vUfEY8T2azyXyJpz4ob8XNzLr1bZW2
DL9QNh62IIiEbuNYVQgxa2eiYmIfxGmfWx2lUBRBMfGDqkHTAuJWgpy5To1qppq9
BvOJ2Es9NuGn7CYmu05DaDLQHfFdMzix1s8fpPkpD50J/jZmzYSKnzSTCBhwqm64
8tVN1DJv90cMKtKa31e9j9Ud9LqWsjZsDbfbjoS6JfJrAol80JVe2MarGW6fcu/2
wRjD/HgVTwjh4gXOWSlM824e+dNkCDYPR5S5FfUvFXBXOOcE87yxI/R/xVMcrVKW
Mozz2x/w9CSNg2vcv8reOegIPCUFj3o1CrVgJCOF5wfqyz0rHJWyPGAoPf3e2uHf
BggNjbSmlEp9QeYXnb81S5m/NEi5+/5RhDJ4E88fnxNh8qmlijEzAAQnM6hD5PZ2
bUTDx6pATRMbaQ+xINzun1ugnL9RQYl811OMzOrmG9hkbBOXzIf3R/D+7dH8xfmK
kWQWSC8zhFp7CTv+JiEMGDxsVrG7MSFw5oNhBnDlDlSIKxPVfCHOSpStLd6ksblP
TS1R3fy7AVm3cKa6MSnf+S0j15Mp/cPmHyn1sfNLq0OfrnqpprNE3yxib5/GBsEe
yaaovU/qC9NAqXBJwxlIgSS1enNZM/dEQXotPD0JRGyhj0lLzTB4DPq2BANJY3a2
II3wqS7o1+HmXpvxCYVcq6HQ5ndmA9sMSrk6YsIWep2Yx3hM9GrdxHtaM96o9GCE
FZd5KjD+Y6J7G4QNcYoAMbohLiG+rzlZ2hApVoGnb8TO2rBPKFe/hObWDF8M2Suj
HYrG6TXwtcerbjmL4J53xjBqxr5lY5xK0atm8AIW0E5KI36KmAMf9YbPFrz+uBZE
YmLO8CRFXvcKiwJ5oGfb+WO7h6q7CXXgetPMix8NcDSOle7EWCLbEKMAM3ynxnBN
MSVr3zDBMdPJwd2OCKNKVEPUCsNWsNRU6znluppxgTFkcni0ibezcMO44pbL0znW
b72ySsWQmkyJFP9W0rehmG+ZSUofsHS4BgXzeonzqbQ6pIN3EivnMgMURL+TtZEW
`pragma protect end_protected
