// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:35:48 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
nfuc9/uNJsoDQNQ25YEWyp2iHaIf9ryeBdHNOVD6SnuQiq1657rnb8/AMKfEwf6c
R/IJIKfC2LH+Y4CvJhijNXDdDuldqFtj/U0q017+7gAtHQ74mq7TIv5y8Z/SGGyM
mP0awWga1oKhNRMutEn452RS9fQZQjTBiWu8+505Nbg=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 2448)
WYzYa3qE6s8VOzCyXpSab/1I2n4RU6Cuqb5+mjr3kfiFDGT85psN2z6wvd067evR
Qv5zcLFi9YEcBgaOjJIyD24e9r9Z8QWKSGJnJJjsHXRKtzU36kOvj4aKNKKQYTfF
cA/I2RIQF/g2CGopLDYriP87VpLWPLsT3MN/6cu0T8Kecx9CsVelJmT9vjKrDDsN
Na13IpimqtZ0fLYoX7JKXyi2HVgUMEi2TVrIg0KO+e7RAnLfA9adUeqDT7H6Ffgv
dkYD6dE5Db7OU0mmUPN7+zvkzByoBiR8puZYdgr9eqblWO/bcO5QlUHI8rjgon3E
PdgqiV91BQi8IIPk0MWlDDh7YK6tKlxJvGkoVpIEZ3RZ8DJT3w+/kT/YEoA7zj0I
W+bBA3+X74SS5QStZTJpTqAZKBkiYN66mqP8d5k4idpiuXnu+jtG0myDvETK9Ie7
H19yVnQH6wBKF5u829ObGkALO7opOZqbuApSOwkbSVdsmZgTr7qcG/chVb4wCvhY
hZ9n1cPDwzKXyk8rBAPgtyzHh/zuMHumBpifcGMWv1MBbuXmza/xppQPPphvkNPs
vSsBlb3pwFZIi9goIhMasVaOML+e/GyTjg2DLty8hkWtNrgUR+c/4gbMXOOhzJoJ
Jac04fgyfXPkuPkWz6S5aS9EcHS52yruHbmRZiTsZuhcg/UcQE1XnBXg+6mVI2i3
24a37+A/kzbr1O0StTjqW4M8DCyIkjoJE6ZoBznl4gC3FHPJOoK23LAqxbJXJ4NQ
jkRrDSAZvRAm3onpW1R2hYWee4B5wR9kggvXYR7+O89WC7tT0GoasCvuLK8zaqz3
vOBo9YGWvf8MIetdJcBxlZ1pEg4QnerUHo+s6cNsIfTuJM1r6qOGzzrqdrghZT3N
7hBQKQWtjm/+nIqMXCy5esVHUEHZBrfTn3Ns2Q7Kjy7CVIukz/GYU/f/x4CQeKNZ
G0BswyGmRj35cdf7XA+g4lNWXlb6sd8WJDjV8tJTDqIDvi/wt3O0InH/EkeDfC5C
axl0W8pVhLq0/u9e4Y+girMkM9HYdnLrDvoiYuRq3qyTo/9y0OXaggLQaXqqqDPy
RWyf7zkZflLw/enrU8FG3rnky/kQQQNw4wU88L/4lfAG0t4COjCt17ZeAhwNXIZ1
Q9Tg9Ai6d7W5/Po3j/TlH5ZX/M1y02hreTs9rX9gF2noe9reN/Awvzfga7qKH9Y1
ikhK7yct8h75pN1mep1VWi2A9bpatr62A7fZwNVq31wyW/knjjgzg7pWM5GZrCk+
JcJdfm87Z//+HCK9BBBVLZfSN3C6slGiJJ6bOSpcUFswVEI3wDcennu1tPzw2uea
Od3sREfruypenmtEcC4/b7oq2hXJhc/dSynHy97scGImg2ntf9GrhV8MqPl+Zvr5
2ZoAZxey/p4391gn61IS80c7DyN74nwiKRZ2IXLTSohk0OJx3s9RJkaiwoVdol7i
fahGbkVCxs6bi0L1lKzHOAm0ev3ebO1cKQwlaUNfOasxfAWJbjA0zwMOy8fm0lWD
Pofz1599pL4xF4Y8HbiJj1nBVq5XTNZNPT0sxcKY2/S2krqQ4tiuRfMfTBCaGwph
ic+P6sZOTFC6Y8DqmbCeL1laFQ9QVFQ+zjcnxoJCGv2cV+weeEoKX6X1qcU0cldG
spAsaozxQFlLkcGXNFOX+tzSa9S6RvzkHu3e4WN1iGTGKA2LIn9e/A+i2SOsXER4
jAW6ecUXfCR0DwmNgr1kEDXlyYCIiDVb1gqjqkJVONYZKYmi3X6/euZ3GWiRrVoc
sDTt8bFe+7SzkD9g0UeQXddFmykllOq70cDxIGIQABrTdbxEdEWBxzcIB3gVJcVI
M+39d8cUDKQHSpfPFVlYt5rs7rMQcReVpGuQU6HMAvPN2GiBQ3iFTZVTFdLC5b7L
geQuTrPrNc0AEfQFbxsk+ErD5n8VJfiiom4aEaE9eXOcICc2dcwstCFc1ux+lcWX
MDS1d1gvzrMjx6gcaT1Vr4UV3LXipcGqfhbHChOoJZ0Hkvr28JFe0xbpqLlfJUeX
yFp+qng4U01PVWFP8s7I2tpBK58lEm0MJjOe0rl/aciQiRZniCM3XErCQxWtvxuF
Mq3by7SrBpHuSz4/QJiV+ixqN1V+FhJG2ky14UkkA3cdnWufjKRn//KS0Xdq8noa
+3CJS94k70BA/GfCa5yiVdwGhdwIfy/aTSCO2we6KoZ2iyV0SpxGeq7n6w+1hVTd
lEt4EO4iw5pVmAptRIK1hLJx79ShqA6wUR75t+fxtR2sAuoLAZxu9wY8A6f/QzJe
Npy7ufMj+VYsokO1XMTh4BbaIkRTJG/8WGr3tVIoRm/5DbLTw73cRpFAZyZ/bvdC
+SefLfs44IBRPGpOUJUt2iUt9iFbAznNiT0SiONq7lSDfG3jR6XtREKMfGXbusLA
iJUKN/GR4twG1c5TGnKJeha7B745ab9S3loqRTOwPEdvBqQe9696Ern6r7NC+SmE
mXQ5GUchtkdyxGORGWP1d5JSTKbU1ux1pM8EFhtbM7OpEsMtA+wTCfBnGDG0VihZ
39aIRhtL7eE0Ylc5QG24FaYkuYvqT3EQlcyajWhQ+FwCswjz+LDEmAx8HhLZCtjx
u7pqcgWutfbU3YOyqSEc4ScxF0CzHOV5gmXUAnME5T9vzbFOo2X00Su2oGrcGB+x
NGTdwtrSBHCAq40kHqqLxXGK23EjjLOcKsBpl1Pii5fNhkYlu2fp1wAKLS5q7s69
+6c6pcRHR8GZ/CCEV/p60ok2XUpwUihaSF3dcwNBWoCcPx/ZfQnefu+/m26rhhRr
u0fWA9LO84diALByYHSX1KMlDH2C+v4hRNsFbAoTmh8Qjw0ffV8H2qURUXRYdGdx
4crWGunph6w2Z09Q22e4wtbGVAYkzpNf1VTtLCbB8urGcKWywKN9EkVhjfo+1GCy
kN1yDp1OQFTzDgn2Z5IF9s6zDsKsThibCEUL0sGX86oqv3ye6ymJ0gJSyBhZ9kZ1
+sHy8VkCB5WgN8xku5k6mhEjtmQTlVMkitVH8HGSiKj7M0AJa23Zpxxo7ZMZIZYn
2dcmmj0pCDGe7jTsfe/Or8J9PBV3IROW2I6W6GW2GmS9D3d49UrHotV+kgFKgBd8
dj2yvYPaYqmNfIr+3nxMl5Wu5rJXw1y5bdkYvlRyejU3sAjvvMEnDTLo4n/esoBH
Lj1lgaiQhOSbxjOf8uogeYTcljJ3+OCUfMwLOKxqvdVFXA0uDvaZ3ZVZ4yUG8ntK
`pragma protect end_protected
