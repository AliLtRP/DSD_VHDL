// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:45 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
IAT83MQzf439xiRJ4UwNlJqMGEJpNsYtikdYVpU9iD0eHbR+2EtAjbo967AD+WOb
d9LubccfF/6vR4LS9NtCfcpnNtkrdcjhbaWphOpS1P/kMFolvmQxkyFK6BH/xVJN
rbETDAOOTSF4MsudIcINX6YfUwEptYcfx8jaaOrKFS0=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 43152)
77vwysXHUxTzhsfw8FPRlhoXRu46W4GOLWbSHBxTnzdXp/VV+DgbmTMOq3OS0Mnx
gJvA3I9HyPKk9EaoIsEB7NyuWXGbBPx5I8WzztP8U5HhkTbeE3tUfVYt0tAaXKBJ
3GeWFDhcw5CJjNk+fER1PjQdJmFjVom+95wPSw6X8KMEz3Psd2NadrNVBln6OjDL
/6i2dsbBIwh4DD8wpyPo+Totpb92nCxdf/2IQ2Vl9Lj4Mn+UicHvMgRv5p1XWqew
ljFuoif0Qb2byzp1y+yows7ApfmthvUD8qWYRyEdc0WTKqIYpFNUE4Z07xSXQfXx
s6xI6ZasqlMiCJ5OB0JFG85tVZ3/8aDZlgcca5htMvQYTwfby91FcSZhJV2obd/v
7YxEYpE6j0ISETtAG8vkJvLETo0JjVmCXvrNcTkBJyr6X9plBC51Lh0yAvE/h7eK
+P2EqCNg3c0V2TfOt7lcLYZ1uDV8Hke8ZN0XFZQlDWFXIwPWduiSyWrzofOVOPnD
xkr7DQJzxAXx+8uvq7DIZfiK8IsUizkZMEYMGxH6nb/gzGQLrknFYATD+eXwzY6q
TweqkJ0TqNANxEmdVn7LW2FOE4q2in1Mn6ikBzraYSNbppOrsTdWvcdU7Y8fydag
uVoAMeb2Tz1oTR8BuhfBCJf7foH+P/tnF87WmE7op2ZVxFYcQuovBN5r690fsDQ5
ZIcNpqhfJSmTzaZknK8cqaoBKMnWn7cpfduR7rsKhxBcAj0+MgCLbrFfmn+4UDhX
Bzfp9wxXC9Kh6oYgCpqLYn88t9qC2sxTiyqxhYk4rq/C6hDeskoiA/Zu57YWULxs
VsdkgUECsXrVgBjkXbtr4ZcnnRprKYvAX/OTiYvm3pFwQmZpWn4Wam/tVLLSXwUq
0oV+AGprDC6Po29JQVcAk/hYVEhUFUEfIJOiBPXQS4F3R2ihLSTrcCeXAklVQeow
PV9vYATcg0tOn0J1dR+EfU18mvKZJNPHKe8AYVDAB3uw81u0y2qyUPWGwLVX3LYm
84+DAH/QZBu9qxgR8rX//FCANQ3Qq/TuNxUNkxFUBBYbwW6C5utC08n2+l+n7mh/
ZPHoG5kMOc6+iJPZXKMcodjIEBfJfCjHiybOxGRaRdtBaoQtTxb6MWIpSiSm8kGA
uRWlivnKYcfSqHMmXsu/r8cOXltM5+21tc5vhKJqu4nKSn3X+MypXH/w5S6ZLldl
Xbqtn1pv61MrWjZtZ9tX2pVrzMrqzBVKEGaXXK9EmbcKOIOLliar4wUbXmNCcoTU
UM6+qV84UipWas5i1D3uDe4vwuTABwWNCzeGunNCgSCiJSWdWgF4jzT0QTd3K4de
bgbNZDivMhzFT6xr9rkOGeacU7ZkovyHEi3JdrwJlOKKHq/qn3G9irfH8TEfogIH
QouNErD6VZGpU8E9jXGqlyKyVpT0jDbJOh8VvTQE0YttKP69w145g7Qh0QFwg3Vq
Unsm5Hw61naJuLwGvjbvLQmxLl5LWzPHmW9/Ys2pXbXJfZ23hBb4lxvzGSszHVOA
H6YwttSShnHQDhWYGHUdIWdiZ+TORpZZnY/ukHrtUWu38S/v6zruFksL/w0S+vWF
gZUpAytxG9C4TGp+G//F+SN4u7/mI5bbac88o0QvY28reEcX0dgFyI0zcnChj9bf
jxFviTb1Sq/sWESP08qSsR3fn8WfSMrDz6N4st2NtmlRE6R5g1lTHdetIkYIfwgX
zrVNlxO0eNZbopkkIKaB9LI923NeEWfGO/Od2TXrC0EgpSCyaAVcvaqJBO1sVYFD
gGOWsxq7gh/i0DCO4JWHSF/OtjCB9VyAP9fX+EN6s+ThMBV6/U0+mIMhYs378Mn1
1863mvunHRrKzKmVBvj6zgOXokmkIrZyO3lBZaQJvHVqQfcqcSYVajKo75Jf0yuJ
9vqE3rNi2XtUOmYlYWRzYTMRC+oVuaTK/W7U4W+ROKBfStOor2vtBvo0b2mK3gu4
8r8X7iz6NjIytWdIO+v4E1GsBBqMEmJfW68xjugqP8DYYevgfIb2lmTrqztkeixR
e3Zj7FThinRUu9KTEi8gbMe9scV5311lI9ThxS+dV0+rP5HmUGzele+pIwKy1If3
AGLX8R3xm2u1qAhJFmAFQlG9ipXnQddYjQhBfkD93lx+3xtE8iw7uEc3Ib7l+9nh
UmXYiw28lGXK2WyU4X5pNpRXE6kxAQFdO757GdeZ/rDjMfXpeWuF7ZcFa0G2enkT
FBlvxzvo9EuxHxAyXss/q9tVMlXoeCmudYTv5wE+5gPi9H+W4KXW6coRiDmbO9LG
YIgy6IRq6eRVX3XmNWmYSwXdYtEoYVWPYHeqsDIUvbXpSaFfLHpgYFvPrCwcy5XP
tubRI2XKNHlxFwe7YKk9Hv09DlPb3XcrzBveuu1idgLxk86CVJjyIXTlVqUTCoXy
a7P1M9I76MChnO7hCh3EvUr7lQfJiRiMgNypEwKM6H/YM/ZNY4ZAKVihFXQHos5o
ioN4x4hfZSKFatKrtLBjAkEQx46eD4BkObn7TbmYK0y+nN2pqonzji1Brk/6iJ9X
Bi8rhrafqI95Xph2v6b7RZ2+nf5z9Y3TtS5t9q7HFMuPrFnoNyxjadyFpZbEcFYC
d6IujabA4SD7tjPq11OOXqXbrQ06hwTMkV2uRZOjf4AU15iAJpjd5idODnWdxInU
djX30Hx14lMgysaLgS1sFveGiU7+ZQAZGgiEz6sHOT4EcRIBWzqjIMsLOaQVqJ5x
4HiCcNv3RM2PJvWmLozbMA5mSiZA82W44NdtwDXlnERz65q5Q6IQj8uZ6kpzqplN
ODoT4/hmoC3sqzlOTky5vAIXUC0K7JBHloodpOLT+dpKwdIlrITg4TvXVGbMkOgK
4xzLQhk1f2LuW6zg2vsM/B+Gl9FBYpcs/8gKgV5o16VlxjXc+FF3vskpjOdccuYe
k7OHJyYhMcJESRVlhJXbPed/fSxpT1Y1gblHrYc5yUZzCHlvYTCd3jsuqOBBt5jp
1Fg01nXNgzcIcwb8m++m2SaNPFrvjW89w57WAORr+bEnBXpcUapYLKGgFWVFlXUc
WIEs8g2ZIQEkZ1Z7HO+Zd8VXsX1QoYyLz3c87qV6iRvastBTGji112IomuxPD690
JpOv9hLP0PqjjH0wELkkdb0dUxDTYLY4/rKOexoE8K9Dunp5v1PUi9yfjbwUo9wl
ZUOllujmEry+97t0VnQFJCZNERMvpAXb8DKa3k1QAkhjadlIDbYXfmfOHwICGhNk
T49Mk8RmtEKvu//XlxhizEk2fiGC3IYF+Tvc+akEiHhn8sSzY1/1aAGpqQ8AZpOC
yKGfpCDyS19azbdF3snNJ0lJ5IODtrh1vGdloGRTjRNzKCmHdp6x19ScyUubw7NI
Z2CHPNl2Cc1zdOmGYr9wJyohYRXhgFE3gPnDfmNa+8UYlqNyxwMowLvvX252kahV
oqsmlsq2qZIJSDQedGgEoYrvJtU55tfKsBfBzjJg0noVrLQh5uqcq8ptuubcg6SS
fMUhqtaOD1O5ZSjEmmkAqxMB/NTpCtXm4J1xKqzGonvD8UGeSclHpPupZz3QjC7S
mPDmfuiN5LmGXPtKueA/8Zlo+YzkQQ0JKAQw0pHS3QY1qZs2kS4mhKwRlvtJrzNs
1/T9p7jNqiYG45sRJAQFMy118LQoVhQ/84rwHdwSPbH7a7mvBu6GIYcxFTre0hRA
op4kzU6EfvgSRLYN+ZajzAHpHfOfkPBAcFKr0fh3gteFgYtOtbnPDs0+TeYKPhmi
52C6Tr+M8KyPR5nrjW1W61j+yFh4gDxi2opziHlHfmRdH4nuKrv4SQ2VJHiXy7bq
gco/mUCBkiBIIa0YYGIF2GxsNVHOXomYV7OBuGVqpi8PAGZo5kwryc0G7/q8mpdm
MQDSmAoTicAsG5nLvbNQXZ+lytHa73SAp3EvkMgNKAv5aWL9HaRxnZzCcJTv99BI
CSs73t6w+u+WQw6zIwKGnfoApRmm35gi5ifBLFBOnBvu/PkX3STXuLUdaAQbaPO9
ViKOzguXCoADcAPAkrd7DlDqOd/Z5z2cqNuGVhuXxWqU7boMafTCjrJKTssdGWSB
+CfU39q31oxRXgDx+clqn7RBr1xl2x6aJxhXLSn1Q4bU/p3XxDUVQWdioOHigEvx
ak1x9QMFVIrX8D/2DzP6qVEnaPjKn5YODo5+nIvMTDJsnnhs0tT7zKlOOC6mU+MO
o9fo8GG1LrtT3nesyi7DCpf4HbEoIIfx0S6wzIJF8WAcHageK7+pT8VhyzSSpvy1
iyU4H6v5uqxO0qm+VWOrL8yqqxIwNxnnh2F/yJ9O5GelQBytIJv0Oy68gD2ey+i1
+E1HmjiAsRyE3MKoyC4lmLOBazytfoKItZWAx1CCFnin1Bmwp4/4LBNSMZy1K1aV
+AF7y0STbvvPHeGQyHVHZGevTCKGr8yDzsYFuQztBOjL4vBOgdQQVWbWnD0z3G8D
ep7s9y6rWkDB6tuiq5O3coZF1oMmFzU8jPt7VuG4kQb/S0E6PDeE0ZkTpJPz5FU5
oCIIsMvlZPdT3qcvNevDmXFHEigG/CioN+dnmM7JAvlFMGpr+sb9vALX8Hnv59Se
0t7xKK378r2RsY6OfOy6FsFzNrtGtafKLZfYWaPseApXCaKhRWJjSuRXgvYyLnd2
CItOImVeB58IpmBxLkypZs4/GdngqOVvmsJIC5ehNZCdDjy3KS36DAtUQMQqFAbx
mGKczG5sT650FwYOvduAFnuJOfHq0drdPU90H+gGqOPlOjhDONXMnvOqNPcFCzZG
xG5UE0ZbQiSGCxc383aQF0N9a1ySn1ASbgpLw9Ho3iEhs0ziQPK6Xu2WlVms1hk1
emLjlCei+Rb6my//iBWZGsSdzGgmSHe9ezbYFhUP94meV/o7XeMyxrnLIg2BeYFa
JQyGoo6aBvBArFC2N3FK8HeZHgMrj2z42xp4v5ntvSwkV3AJSUDUyaUQJCJ6dFFl
bxebIzlD0gqKCDRwW5Lk1kUUw/pVE83WlCDV5/dHIMl/PGcFgimcq3tuFY9GXtj8
Znbx4LuJ8ZorruCFDq6TAGjk0Jvw+KA//cSTLBa83t2aXGbD7FZmKC1miK+MZgwQ
cmSw1nv/jmXd99J1xAjJUKsaAleK+hlDdYs/7B+hSr0b4Qfq1adCgEPfu8UeDvxl
B7E4Ef9lw7DWuYl6IAh1FT0Wmxel6oBqhrqoG5H4vhkulxBKJAKZExs/GFLNKZ/b
L/p+780stLqu1x80tAtNUtVHnQoKbAhQMOJnZ7iZZ0xaQ3L6FOK7d1e1YKyJQgOP
9pLyG9L0Re6FeWFfQFbZ+I8PwiUcE1V/bgRVweKCp9/wPZ+RZlQkyHNYzHCmfRnb
lbStO+0xGF8pcwvDOsMg/swOu9CTkmYX1XQ7SxCxVfCFfEDxv/NRCCmm93lepxAe
5ZoZTYAjrgnu+nYf9OfRhOIYEOWBCLSavSNKg3s82ROK/Jbr7lfv9sFU+ZMsvFA5
tAEUQtkpMaMgF7PyJEzPlKmsh7rLAe1sKWXt3lCa/o223NSlwb1O1ms+Toyp1xiL
AgQui4sLXJRHRMxjFsGprjfiuEyQJCkZ+8Sm5F5N+zY6aTIZIN+tItvXcUYDPD6k
dBt4s97gIc23CsNr6J7OQrSlbzszFod5q66T3Zq9YCxvftwTkBqiIESL1tdZllrB
XU2D3LFyaVf7DAKiBec3uZduzYT5r457VNEaoqAA+YHIM2uqCZAEFXhdHWvzCAEw
fnA/75NciHuHOK0uu7ksHPV/Lx0P56Oova6lsiuYYYXko+kze1jAghPvyk/J2SZk
IVNlnyWx+oQ2OaWNyzwYVPNytLD30IuoMlnOboe4GxAri7iFD9J/S0Fx6gWLIbwU
Jlui/NVV7tiMzA0OY86f4nb/LM5XPxF+Kj0hZN32CaLnYuphfQNdLzjX3s/stD+K
2NmvNxaG+QnJeNy0f+tqom/gOAnYtDy2gs2Y9QAd0OumGp2rHhlbczuqZo5p7G5+
PZCtM1xHaRa17NZLMPeKlN6NEQqII8/yPD4StLk7uUd0NmYEtJrWJkjMypbzd8cO
cVYX17VhJ+zypocLHpMD/58CgTWPZ5IRMwyErfA7yvvkhW+phHXjDs1AkPMMHVeW
KNUKlywZztWMsO3HryayYtz/ptiuIcOjWx6bIj3JtuZZdy0difloHJoytgEgi77t
RtRFUeMqDlaQxX4G7UTNdg3KctBI+Z8cMBm1444v2/e5d43XN3FN+Uq4/KFa6h9G
MBudGCEAJ3Mpoc9+4T4OGY5x8ZyBySCvC3LRT9x4b3ZAF16bp0JPqNKKXvswtGLE
CGR/ahf+KikorDrL9b/dX+XXmZWamWgcRmsoe6XmV+6sMPxyELtz1w0lcASfuQ5N
M9guj/TFd7RthNhoI12PheeKxh12EdDM5uVOVUcLyNDrGGo+MrC+ZFVQNWSKyiLh
dKDFShGLd3W4fD3lV7q5lA8JPhEdsyRR4rOXj1MwdUCdbzyaOsVS9KDomPLha7XX
q6ZY98wHv/fpB05XXdQlTVHBDgHX5Ptp5i63XU1IvIuXAq9shWXLXKsb/3pMCig+
SKO1Qni5xV/Xj5yhPcyoNvKaNBh8tX+PJcs5FoBCPmA9K5yxursxZ0Ubj7RybbV0
g2OvGUP5+8Y+trG+oiEQH6WYbuQEe/UkidUPAjPwOQd9f1TKdzEIgoVywh5gk4hf
BjZOgCWlbdhss55YrmhiHbBDIWeWpx2epTvExdJWDz+XCQzeuX987Jq8Ae6lyfgc
EjCr5pzysCctsG9kh+B7VX7YvM+XH5VY/pJNY9oWyx3DDserOysCuniscKJ0Z9m5
DWJDCKNcasfz7/WZur4gkWT+pTorYFsx9R76DMyIR1MQdhXuY02FoYMpOm4znheo
T4qkWBmGK2IKkULewg9B7s/BJzqMNDdKFIOD/Og/y5DNlMq6TKALoy/Kjb7O4OB8
UqUgIx/VV54KY05d6nY4E3NJbSgAHQysIrXswTfVNGf8BCyB1e0GIAR1ic+ZjEoz
cToAJTlgvZW2M+4XrZzzL6MYvdz/QSqj2PCPM9JgtVx/lET1MPdkFt3gXDghBTwZ
ORonlerzGMRGRCGAIKBFAIXQjuZ/ZmsTvxmSluY/yzIIyf+cED8yh2NWckBRpGeB
lKiUs9TY3rdS0L6ktyJl/PNab9wVORCIm+0GhDcUc2DKmVhlO5TIUGA2yhuciTjT
JDIlisqbLO6LZgGcuxmMYkJ0bHXzEPr3ohRRIfWgK/GrMzUsgyv198MVoyTw7yoM
PGL9lT7ImZGTUCXGA45ve/tdO3jYa4+J9cW2tRVgizmSSMzH76aARKNSlh3qQJLv
DaBs3OQxvDOwG81pqOOp/fhCNsWZgu6N8eoh8HIRYSS4XvtpHGbiVUoSsejyy5Kx
AAOpKFsURTHZ3KDfaXdQaWC/pjITU9jhVbRh0u+NJYw2JgUkT7Hh7xhjQVrUUISR
beNTuoFe55jbNoX5bC3ddDtobHK4BYiCQy4hYjAZpe1eS/4eO+ArIhdmpbw2UPbW
wWXEDOlmVoV1w5oeYhT7LNXOCG1QeqLV1W++yc9/cyUlFKAzeC6GqPv33q2L3ZfL
pV/EEDiMgmsjRE1O38VUeXr5pRXU1VdQjTc8yRTzow9z33DwCS58NMSzwAtpMGSN
puSfKVMKwK7EXGPMzlMEhNhr3o8gkDZGO5mWvWuyBuPItuNbY5bQohDrgnjYxyhA
LRf1znUMTg2KTbGf+gGWD97Ivn8KOF+au5xbDG74VMILmni2N4wevvXpmhex7Dpe
ubNzZgFTOkNEACyNVlEC3LwH27UTdFq2ghQNJZGuVsGaCAaXT1bmLWS6INw+bwqn
e9HKKv4JspHWslYvHG1KcAeQBvmJ3GWjzazIyKEOAt3/kcbckPXLJRrg6cHwv8AT
OASXLW3HDIHMDhHecPM+kgekrNxfEg+6VWrVwMqzzXnYRS7Cz4Js3/EqbRKY2uiq
8IpT+VazSxEkfeokJ+BKBOqIWDuydj3hmrhvvqMJp+exFocyobMGiyGzrgRWma8t
VzqAdHoNe9CKijC49pohXEn7lwB1ooTE7tE4BsmukDZC2/YyQ3Ev2uvgMq5/BH05
u9Xpnzw1W4/OZr2Xt3qZM3t3bph3Hr4NEbRP1j3Pgg23xttuZkkEPd1kw2GlhN8q
z/1SjzL+BiWgQifvmzadlGmT2eebtFszgnfsoMF9xoxsG+ihYM9/JZufgdfJwnC7
J4AzAd08ibAOIHfE3ZM4T3qsxo8oqKKlj0mCTiogJcgNeTWdSzCB656Bhms1b/oE
mJMhIVG/MqHvSd16e1iS8IdX/bY0jjpTp2E8D75JK7Qrp9BXmUuuLHrzQ6NwmLoT
RKTzPCaxcKkbTKxbgI9oNDduyZzJ1rzpLkFOuJ7oJJpDVwMK9b2lRqjUx3y3mmZn
L7XzSjgkYBvGlwwGLc3Ok3P7NqlO/DHVAvhClc5ZelUrUSOAIcB+iOlKW6U/qeEa
/eCI1ZE/t+DbAZBnniAPGXfNBXE/Ar88cRb2fXw6dNlnSkHbpEv5VvMI1tKwTtoM
sV6rGokIVH6CHWMq8U2dcnUwVp/ntXprjZmJDuCVbRopLJuCdNHZUbG2jKAOzgpm
OAXpW4cbldpmaWFEX+io28MmLbMh01Vlyynu/ieAcozkxAlnDThMfwasw7RMpjxg
ZccjRssyMqdQkOCDmXSOq3fZ6hMNNHyBL6Pf4aljbgxMakz8Gf6AyAwsltT8udSC
msNkHFvs0o3cRj0Tt1x0YVa8WeUvnRPNsPBGm4u0tWgom9bfoCBCF2o2/VN6/Kwq
69/WBmqn5Xw+YJvtRNUT1PfFBdMpI3zxMHzECqyMcjlBKydOg2erlkJYEEWkDRYW
Vj6dI9EYgVz/Nocg0VfX1BMiu/0SvmkDvT4Cd2SZAZGF7Wtc2kpn3BlKE4VaoGii
R+Svf2pTSy88Rob6jcWL5yd+86Rwp9mYlWLfWNRRd2yRjoIY3LVTdxb/4pJvYqEU
RFH5om2BFB0j9a/Uy8Ot+bb1dc/Q0Zs+usbd/+C87rJqJ2w1iPVMcx7Q6dqJf4Jb
A6OldA9d5ZBASTdL0DykzkkEe/DWrL8+v+7nwx5GtYEfZub0iHVr3+bI7S0YR8lZ
YBAxA93Wv+4HKbrDKqW04Sjas/32bkYpqWiwIvVuLgKwnY8ayqMoxIexKE3agIfy
h22AoOrxNBqNIDi2wivAE1PyNj4PKyqpf0nTfOj4Fg2UfGK0VoNEoLMVAlmRRGOu
gJ7SI0b22bGJuZmF5/auTQU1OoJAS4YQQrsHKRt/k2Ly7f/tRI925QIl/o7tzXEP
TOwbpuLS+Z2JIkD4RO4orNO/Yt50QYaK6bF48tBoorIMrgDRi8FXFfUP7kGyqeC7
ufJpfWR8S1TITXypePb0M2qRO4zQ0gmBCpa5reBjakJsmEYqtSAspZFe4x6AW7z5
aXrdNAGga+7WLYoxUIeuqqTf015dvZJ5Snogb/N0zvNHVw+Vpq0nt1dU0ZLgZfra
wc4jH6PpruSamXGyWeNK3pJbt3rrsU1S8Kot2kJopZgAKwPaxdM5d3tk61KH9Nuh
BF7nw2y8K536RGy+fgoNNa/jXwut/zvrkoce1kZvKfu7lqBgZJkA/++eVGalz1g5
jl0o/bgWQTpj/oMmFUJ9JTAildpaNWbXiu29kpeH2Kvu3Oe+w2J4dYhoRDfDwjX5
z8J1xkmNG2IQPerZC/LBsd8FovDrmFnTNPwxFRrODo2Yf6VUDlG7oDF7MTm1shJy
jOBYdrv12aRGZ/lxau1z8vu7GRPfrRZyiGcjsCvDy6D8soDZm1azKL32ns/OLxJf
a66Vf3gnJStxqa6/7XzHiH23tGvOGRoI568pm7Sf5aNUg5wDDJyJBlpSHPKJ7vIU
HDCavQIDOxf43fvGKLyMk73BbnY/kyJrWX7r8E0MHkbJYQtsbBGukIKb6qaOZWBq
6wmRgBWFArLkqNkxXUHB1vWkMiOcKqSUlO1DCjco+MBgZ+x3vgUWP0iZOZBtN76M
YG9h8pVolllY5Eh2ll5v0/zr94NdBB/oqjDPExEq26TZ6iJ2t8r8nWzcUD34O/Sj
anF1Rh8lH3/NMy7up1qOpr5I7XkrUaahTNjZHLCOFArMsKx3P2Wuk/7vbD2ERMx7
Yj0V3WVb4ztN5EHxN5/QFXEw56rCHOEvmcPXYoNc8NUwwzcj5AHG5E+LTVC68zbn
AJlTEtkN6et4fxyDYTwNzUFAaogG9O8yxKDY6t2wb4nlLez+ikgOKGFrmywpuI5g
eFE5uX/M1yGFg92b7hkojZb+nlmOkDS5zRSjU6QqSLKLb8FX8UKyddryQ4BqWyhP
r4UUccRP0uBXanC/IIkIlPFPHsRIKwGRKvQowDVv+rKB/c+G3hUx2/W9IKjJs1X6
FWhYVf796mpBBUvE3nODRBdEcgpJCFADO0lAPDxqid+LQtGH0iLmODIV2YO67b2W
bde7fXSolPcQnNgb9T9ae/BS+JaZjBnlBoxkbg23fk3Ue6AJu9KV0K/ts/mwMzSL
KLjmpOu8qA97+jUassKxzCZurHizrwZEk3Gr/Z6MZdOOrorSVMp2mr/hEbTPe2FE
DSjyLBuQvXkeJEavaC9eNH+Q7kD+2/k1yWcIe1YWZNxK6DlA7UQ4cARCHlIJ3yBD
OG9XYqXZROHYDhQ0nN4Yw8vCYVP1+6tlpwxkcCoqJ0QIv37Cq4hLJZHKwA6Ka0iT
rgATVzYECggLEEhRH3PULspGGr+1saBNHvhp8yFL2uUL9WdRPiRo+n82e8HDBfYJ
TvEPQk8JHqXOtWs+R3WC400/TAaYbPWyZXwsToPducjHEaxTSjwdGRq39/39Y00N
7Oy3K3or326vfJArPesVJgATWuL6O7SgWlkXga/vg1+8HXKTil6WIUS1BDcxn76P
gGcwjfbLiAM4Xfcjahv23cNpFxuqpBSuXUrk1fTumrPlFrlM4Ldh1/lDO5aQN1H2
vuNI9ThoJXmcCh0A8Uyiw0ZWPQiV773hWpD/w4a8wkwPHh2APTZaI69Ue6qAi38l
4v+zv/GYy+glxJFkbbUSUqd5klCVjM42XpcamQa9ASjJ5tT6/j1lFguyGWjKFFYc
Q3QiP0YqTj4SMT9Kzx8jyK3kjuAzOdB5Hw4cAuNMhm/VXy05O3suYtZTBLNvyGqO
dxUsMokZrCdii5lOTPZn863U+TneJMQl3XwBn2mFCmNobPGKxmqPzBIcQXGgnr7/
L5il3dXE6Jd+2uzM2WHcZnWHIpP5z3Rr7U3kYdYGtu0RKIfoW9IW3xiyVPkRTCzS
xGDxb2cpTzTDeiMSNJIf3xJLiZVEWbPvxOi/Q0nI3wDh2oTcgPGCKS9qPW5Z1cu1
KHsKy2aRm01zt5RznAQ94VZktooo1mVEJ886YDea5NPa3QA1BlEv3OrjuS7m3+uF
b2u5xQuBclk96y8On+a5NjD5pi5dI4H01joSsmF+CwoA5okhCo6jaKjN59HQFO2U
BMjnkVb/d7dMXRFim/RZkKR61j/R5xPD/4Hqvqusxmiypb+qLoLKw0s4IKVboKdw
1co8/y4Lud/XW+X5tjnJ78pRHGLI8b81Ak5xeHeuibPqA9yu7WexWD+aa0p43lJX
fgpvfSWWudGwkmGcCYZyWtabs4Gw39gdTdyBRr7TVzltIzv9z5i2b96e2mG9Irat
rX2d+eQenibFDfoyToHhn4Sp08kk2X+wGlZ9lX4DQcEDdljvbtjNURSf9g7Zkv0B
mYtzJ4MBeZQiwPgSpK+6rZoDDrKzAHjg1+KbxvxJ6bdUrYC+o39MgBfLicDZ1oxb
2LqyCMKmbl4/vlNrwN+bLSSr5odOb2hUMvuePU2nGiGPZNe49bvKtJgB/ERlP+wQ
XCsyDG/tLFj6HQYsfhwlg+W/q5TEmlWFRQrVhblsMWJDuRsu7gBAlx9xq8mDjHHO
7wWzWjWe14hKN7qFpfgjsbm2gLvQfSEEjgz2AsceWrER8VfpCjgopJ6A3HBwkYE9
24hG5O95bGKCMi+crspgpwPPKLBdEcuc/md/6W03p3GXVYAIwD+xrXTDnmqWBOOk
oGAP5N88mKPO6DYpWQaWPK4iSBJmV+JvaZ76WBmWFfyWQAYvEVlKd6cf2dYChFtC
TeZu3DL4gET0jFYOWhZHqU8LVhyog+3Sq477Y/zqOO1CLdrjCAm5TEjhEekHELDk
/XCMPswG5A2X1JnLA8gXk4Rm0yx4/dWe3LC3srF/p8ob7wqTxMzkmrVvCxioHy8O
t3x0YfaGkZgBzpbW76iBdIU1KTt4QF0+qsmoP0A7jWiJtJH61igUPPIEgNm/9yTT
P1bFRHusK1o10ixxjWt/LWFr7OHMvH9uS+KA2DIV4/oR/iqCFeMF3baOt0nxgMYj
sqe2dwiGHjlx68ty9NMjVlqDylugigexztJQ5gG7H2aOMP1HjJS5/41g9+oRtc9H
9M5s1CrYKY+w0piBVxv9jUxAX/5FK/PhlcW0wrPDJFigjWdhmsjYJ5WYIs8lecs/
+5AvYCg/eOj6r5cVBbEgjuAHHNaHwqTeJ3/a141zPzTxT5uJnLNQMFyF0a/wUmDx
vLXKv5lV82IRMisdr7EEIdmjMKwxyM9uh2z/gh0YiAS/NKH+e/9RgKlqZM+rq3Dg
klpLJp+K4jne2dro+vKJ560u+6gcpO1oO3sEIayVFIZT3Iq1THcHNwmT9nEZu7gb
9hzKY0c4w17he2Sma5c1l6uMve0DdsIETgkMDwxr53dkZz3KleBVsTjHsQDfDgE3
bhikYQp3dkhmYEy2zEt4YGrVf5BGEQSd6ZOoNVVMdF9np+urpJWU7SQnau00BObc
kZ0r+xCGsN7La7yEX7hfOVjN6MtVN3ys9vrFgjTag7nVGoiu736TRT8XUGjo9CiS
gCGJkXwENrgysS34rKrQHTf2anZwJ250e6MvYknBMpIY7mzAhQ455bh5OzgQasKQ
lWPKrRoosaSxUAwhDVhtT/G2mdGeGsezzB7flk3S0V+vNGH1n0/VFjRnl0hZXuFc
01ovT8yoDXj/Yz14Sn5rvAaXyfFG/Ck9ovOwFIVy1wtylEZ84UofkTmqDFNJhwVv
DhlFa8PqcbMa3850iDxe2OLXHRdjkcIrL/CgQtc1bw9c9R5eaWIRjHp5QbdfOoEx
vU7Yzf0lFSIeNjbwQ4xBwsYIcCfVrbxoomkjsMfnPi2vT4EyHPAjSOfL5SOw7yEf
rRor1DyUYbyafbQPkcsHLWA6t0UlpcK1P9neR6sSYXFGJsgQ598nj1bwYUtw+J05
Y3tkKxlRIjaiXLYHtG9fUS0Mik6tN21d8scRsGllvMYWdZPIomXEMUr+bDbWspJt
c31u0UTDskzTL39E52P0buIaZOxztTBKFWCl5J7guEUf0ZOeyt4Ds/vxMTn9oX9o
5R5WbHBKR+6rdzBuhZkw7kFytLRYEkjrKuSsi/i34kVHKdhNWoSj8WtDIPAxMnax
tYgG4nQv/UjbCCzJEQsZsG3bkppE9md3L2mMEhtAJpA6LkI3txHpSStEO+ZXOv06
bWG/Effo1hTZvDecI0uYYLNqekJuXBhGEfeVGdpFeda0kJUto+IZ8DNLVkQIwijW
1ewiZ+nsUn/sPjRI+b18Faw2/o7pBq7f81kLvEisawHUG1KF48i3CpYHxxYlXaGS
MnjILhDwxWRGIQDeMRKDLUjiAEYoZVpjPRxJrgdAKAeRn5keeOf6HJQJuJrInAFw
3VvLljHm8tvhz2JKUKayKm/fWQmiWndue2QcQ840mbgHJu0pUvSm28KUnEYMu/8s
rF619RwHtphqLo/r5Aq/NSui0+sHdx/CVaj1FPQjgtwMtsQCEndlpC2oCwrmthC7
+rdUK48SCoaqIoboNdNK9oO9dYG2mtTeXw/28ih4rjFeL+2iupQdAt9NGOBt8kA/
wsGefLpDe09ONu961i4BlIQKLNrJIq/dxNf2Aqw0GLX4fpf589zT78ZCtrOhbDLe
w33CB/K9BfabOnml7fvS+l8tuzBMGUWYwT8EDYz/C37DaLUlRTs9cc0uWdLvGlS3
qp8Ye8sbyKZXBBTWJQC/tIBh2f2rwSabkEda6OeUTIDxo9ADuuTMHUzfnV2IUtN+
SNf0eE8iZcYoTsk51DCrKePA/737Lyb0axdJ+gwlWzq4oaRk7l84o5cyk7Kw4tBK
lYQY4DZxZhM5iL3uLuvGbqyUZpf2ZF6JpE6HzmrXElODAkc3WWvazx6Hj69sv+uC
U3+q3RwjKoDbCuAb8qU+ewJwz/MX76ISzdVjJ6Ov5tJwPTmZP3XUAgeSIPV3xzxV
RQ21xczZIpgj4YBEnprhWAfC2JWAIj9y8/xX5sh/K+vmvjY2qMDtd2qkX2sZultO
MOOEq2iLiFjV3Pz34yluefYifavfVXnyYh4FVx8GC3mdLfm2MD6jAQy0Z4J+S81K
40uTh/7+VOpwm0gcN+pl7rIGLahVlCK3ACd2EDIPkJIhG5b2gr0Tk465iVK+zPPV
hAg6Ah+dWgGIcc+kWj7+fpLLFNj3lp5P2UThHqe3LH/lzkQ51oIB8QkQOoEZSckG
hXJpyWiHAHPaR2fvGvUQi9IoVeC1zZFiTPc47pVt5Vnpc90HrBamtABn1zEbZyt1
7UnOjzQdHXFx/IruhEQtcpXB5xYF5+TF0XVNfn2tEsFxrEuuts/sh+KNsL0Nc0EC
xnOOQ+rlWhualz8XMcnj5P89Fmw+yctau97goWnxZ1Ev4IZVslhdvfXvDmAEYx1f
j34lc0cshRhWFAJ6UfQZCZoPHLpbhiJ3sEkiBHTDL1bIk2w+gPl1MKR+OLSCdd6S
l19R+R65+DBUFJryenTojUE5uK2FizbQnPdQMV9MUs51D3ySU1ezXYg0zeMJg/gF
SyAOtIag1mnEymwczQLkdhDZ4/nyJKVLtXl0NMGmr8rD/J73E12chpQI3nHr4zGc
9c5itySt1IBpcLhsISJa0w5JPb0RYGXnHs/wltzt6FBjgi8sYAB9aSJ+6vcyBDiF
hPa+N/mR7U+nM1joQB8CgIpmwghWRIKk3NnKBkV26vaurMvWxMPadszV5MQAfbzZ
Fql1F7utVuP1RllyP7/Hb4esoYNfEVlBLm43/c+Mn+zwtX8AO7yb7u2MgCDSO74G
fdxMPFcSQVqucJfzuO+kPmXjitLKYriXFGZolyfZdOUXBRU2BlyuJemZa8NJZqG5
cpndLIDI82X7ojcOcoauh+81SCPCDPAByXs3Bsy94XhYIXivTTL1Ph3HcdGcPCh5
B6K/F0UNz89c1wo0M6yicupzFf62EoUHXb/el66fZJQx30Cw4tbfgJFrzoGBT28X
Obfhact+v/riIzr+BnwMn2U4jvNx2IuxUgYK8BvmWQ9SVMp0OfKCiHuhik86ffYm
edFC3mVV46IoTgdI4QH+jLpgEvEHQLgf8lFTrr+2aTTpTSuSFWsyGKxTFvcxpwk/
zJ82cRyqmqKva06fI+CK0B0hIpFN28E9YToiaDprvWsWOJD5E+aFt7F/v1t43GtT
MwR+wN5cOals80q9bFKtQusLWcRs3pw429El+pnfdWVR3vGwNws2WuHDS+7iEUA/
DVecBty3hFAhbcVimadQv8hr3iLIOpVbTvMyj6XbdlnTLnweTDLPqiKYqEiA3k1/
CdRfldHdrgcNU9wCKmg3G2ck2h5c57pyiggqrO/DX082FM5ibSiZHsSUTSF3VBba
FEfLvsh4K21XGEAvox1VM7MFImfWsjxEV2Q/Efhf7+7Q++bXGxI+t8wXTkcUj1mP
wbEcnVruyvP919t/9koXWl27fHxujLs0pcvagnpA1l9e1eDcyXXECXo88LfV/8Hw
ZhKB1LGzuAk8UBO/i8Au1lfaHD7kjwwMi+c1b38IMIXzlrP9AHGqQdBHGUH8wpV/
eBWbRH3po90BXELi2XZhCUqcm1uNFpjtW7ucaEKqqnrO0BSmviBOG9zltRBUN98p
0aaEyJFv2+RnzK0BS09x9FZtDG9Ui+c3Ny5G57SJhUPvMIP5Iiifp32q53eimFbF
/J0fJeJYQvP7YqxOMsU6mczKAyaaL0p1xYGOQDtMzuWa31P0bYMSwE5vQ+0aq20W
WBnwBTrKIOJziBJl1egwRvCddEwx9OZHFC33PZmj8WxCeha+My6ThObFQTzspHYh
jgoFi2ajzZ6w/lz63jnBYNM0M1XKx/aTCuhuO87fGdpmMxIOSbZMKJm3SEdtJ3XB
AZIUDjC4A/TzYpYzTr+WMJbZSLV1Zf3BL6JfpV84jmKfQPNF8MNrao68KjdpcPfW
b3k1ldXLYhrak815uAWUQhhh6LSYsA6os4uXQQ3HsX2pmtDsHOiWqLgSbWcNqJvb
hoF0Q+mgsS0gzxP2tvfNt9VuqwClfou6fl5n7YhC+17gTsxTX3Q+vZkUekaGuyUD
F2RB0RtBeUW/25zoS0MNgDbwvaXkGyfWBLMKdlklTD9124A7burxAq0bkZH4oWq0
bvPukykUD0UsLs6rISuXK87Tc0nwzoGO3yLBU0TqcL7UqyPilfCG40X4goZ9n15H
k/j0ifYKTMEjzCcbHhRxdgsCzKTa+xZl+gkfhqrSAxIs+rvIFkiJfFKL5N9TGfy9
oEkhPDWSHCJOsf8RiYYMiSQU1Fc2HgMVcsTCJbutsCEE4vsIwrkLs6tClkKfreFk
M9TaR8p+ngGGMmGxWDBuPpBZy7T7t24Tzpimg2amfpiNp+SwePoVaN2fmElUhvC6
wbKwT3UDCdNRSLZvUXHy52QU5pE0y86GJOD7V0OU3JCMN82EydO8eijI4csSPp0n
s9bAZQ8RzxHLjfn073Wle5DnCNOdYVeCoePZgJ0BJXeb5vtnL5C8uogQ49jcw2DQ
vEBKYWzim1ZmUETD5F7H43tA/5PgsVmuP1yjvcOTzXq9BNEeWQLa6oUQwmKEgklV
2LrpSCIgA2kviGQYRBhE4LJ4CSznLtG00poGadb4CSXh01ZDxfRFFDNGCPGzH41n
5C8A7Xn0sIpmf0FoYD7VWZpEhm8rBnQkjivBjk7IcBzct9YMUObY/LyLBQAwccfT
rsiSPD+3849YvXuuZU6oC8NmZtBEkOIIipIfip9z9mbCKIJSE2GBK/aPuPi/Ogdu
6f4FpZNlXtm+J9IpK6ZQSRJA0l8hHgMJ1iDC7DcmlvhvJRMza+IJS2AbHnJCJ3gL
RFLokQIpunAYk6kvWFVmR/4PpaLwS4Lgua7m+4OwzUxcTnQVuSif/K6w+foHahfK
jsnOEHQUTXI1KIhFQ1qib+8mhCY3m/oxIiYrG2cA1s/lwWLIx8XRvuZo694dLgmf
dqFw/4Tl5AyV7sTeF6ppwOXR/wXVFmegIOJ2fLbeaBCbDstGu/FWrs1Z18ykXlD9
l6CDowKh/MI7Vfpd8KUBfxS0g14eyTEkReYJEhCW0GEWUgOlffyCfZR61nJT0JbI
iZWkVVil6KtybqT4RvfqEpSMRv40PkWORXbD2gYSjJMl/zzcFjLWDzYKS8gmWINb
aWdqFxjmnsxlJ/Sfpy0xn3bp9MJoovlnCG0mgo+Uq1ez+D4qcer7fRG9bQP8Lsho
qgAD2CdEiBinbce+/I3jxgwqwXF0VaZ0HOi3O2VV/BhSFxGcjC0rijQ6fvrRXB+B
d5MR2CapNoglnO7XKEDNATmA24OCYkLGOBRHkh/K2vzVWm+IQB//pi9jiDFx/ztV
JFBi44CCmjkMN9RPkDaqBtMRjFQClO68FM28lbilS3XLONeiHI7VLnyJszKj8iiS
l0Kha+GQgdaDLxUIHrsEcENZj411yu+J6MB/5ZRj0lNPeweqxLWfOAa7FWyzGnmY
zwJO267LMXWGd9I5LFQsXH6tHgW/uYfbtV4FvstHIzbU/XB8/Ae0B52OuWvvI7aU
BI5VxjqpQL7KjXsuhBMTxFUGcHWwju0kySbSug0LvCu0VVBTYISnxYJRv6DfjtvR
XsRc/nSrY1HombUHhJbvsL01sya2aNyw4ibc+mjEF7UTZAtGSFdwhavBysYhMoxs
XuGtDkTM+mDkP75TKaARymFON+y8BMX1CRaHeE5gTxSedtmgBy3knjd5CKbgG6fF
s0wSGFQSZZ7Lfy8Tx5EZgjPyJzF+HCVtSSJRMyjMHDSeVxHw4+J0e1j/JZ9F5niC
UediaFJbVVCT7bTMrcRMPU4F617hCLyyBlaYSkQgPDFQ5iI9ZdlEZBAcuTgbl59G
Fabk4KnpkdjSnZ4gnFoVrZnDrhKks58s1+4oaHFX2hzsjfOG2EHjgpUtSKwYoMQU
CBnBtTIq8nSz4uNM/rgrzSYUm5xZm54KjOCAteqOzCIhVuPgNyLZkfdT4M5nklxu
p60wVp01UgVggfCC8NUFJw8p9ti9s05Tp/zrUL8bRjeqY2ZoJipnpVUtTvDUk99f
nWSXRJZkDYMVqOVdOHpJhtusp3QmYsflvyajDcWzTe+KR/hmsDXeY9jl0T/6+jeM
BCl25ua3wUXBv+jDW481kWKBe6yLQi4ZYF2jI00Oj2U4xq/f2tyvmMjW3vR07Q0Z
pOxb+2XjXJ+a5W6NILr5IDI1nu0VjtsekPbv5qgKMlVz7Ae8RgoWVDdPzhv5w5vB
ndA0/D7oTeQcvEMT1QN/lBWn8R+V246wQLmDYXHk/baQ2lr0lqjz2yioSyGUrem3
57VPTbdhj5sC2LL1quY3tzNyO7jYVlNGUgjc60l8ekbRSPFgt8GFnUpqEPtYK7Gg
4LUzaQMutRuYjwpzeapWK9cc74YsflDwJnZ0kecJbZimNaODjKx1EgkHc54xGM/N
1ShSZljIWNIj3NMQ7RfsgCg9NwifCrHNGsj3tdA8d583F94uOMyZxzr8IUl6gB6/
qAkdezn7cqV9L7VUiQ24VOASd5vAloxgyBqa83zCge8qRv6OMTbdgsaf03jZjXDd
5IVPn0e7+7hbXLE1il6q82gdtl5vS0QLRU6B/6xWIEETsFVt6Ltf9iBgbFn++0qa
1yPMS/ZQxs6bPoOOmTQopisRYg0djoaOn/TvmDXpDlgop+zFFYLfPGEwEt9gPz/p
bEFa6iG9Tgc4tkjIWiI/8SdL/VqSd5o9GPDBedXc6+LdbhKKUfAtQ7xgBVDIV8JX
Bdehv9I/00HEVuEvF3/lUo84IGKZLnGr0FiZrfs4wZFxgj3KMrheE9y3VtlDUuOo
JAAxSOmf1lqEOn2HOiBwXs4SvGymLX6GUFHxqsvPB6aXdlbGTFWa7erlJObVDk9Z
JKAVJpUMv5k8JYLylBVYwhKztNo+pL/APgPHk9UXIBBvCZB7mb7e/bL/nzE/iyIA
9ixiaGhXjhXA3K1b3vAxUCSjusGkSoCQZtCLL6PZIlN3SiKf1vQTp/nQROeL5JBj
OG1hwBy3gaTJOYXrsrKLGkbqYO6mpigdYVl8a0ap+tEyRuhqc/xmaT1i9vu+yjcD
HVpKM2TYYSdh7f+Jflhuge9Nm+T50o2GU4qxc9xO1SSQveTZH/45sdATrGoxxgmL
+FM/z+hghJ3/s8++cB6jxeY6H55pYzlbmLgSM1/OZj3KdvFEIsrqGEih/i7Jswb3
Q5rgOWcIipdT9yTPYLPm0V9Lr99dKRmYgglx5DIvCDPXAXbezuBdrAKKfwKQIFmO
mooV9JLlLufNBHJASVDf0UV6hVvPzbRvW1VNAuPpnkPLyJ4O62Uq1O+4rzQplVZ/
4Ivqgs/3BiIB1AvbK4MnqzhdSdP+zsnsjr0kV+4Jg8QMKZhY+AunQr9RP7Nvsil+
uTAQpQQgdvOYJt1F+65MawdoMcSGgeVbR0j69Ooq0ZH/92Fo+32B6TMg6wDL4GY2
28esM1KTSutMCG9y1IGki2yAT+AjrF3nWoy+Z/6ls5ki4LaH8EAruHmXjJbOFGUq
PFEqecGroGU3elM60y8AGqikDT/58iVCtXDK9Pe8903buKMVhBbcetsxJBSxunkB
iOZEwh8Rpp2tre0LghfLVO0jzbKOvmfpTCq4li3aePAOwwOl3c5WMCvfQ0tpWOkh
29es39r9ddLW5f8ncJhRsktCZfykwmn0aPaT6ATQ/PyjEnaaQKfU3f+NuXBWEUvS
61SjL51BCwYwej5lp/14JKSSFqtz5nY6yHhkQqPQ45lZBNbS8J5a8Dl5Guqe1QiZ
giszcSMbJiJ+/eg3PytOvT/1K95d3fwCPPKVkPM0L/es0JP62IGU+8g2c+2nwzpN
41qdS4ZABEf1RFkXiiaLKi/HhMze8UN630u/QuP6SrKFMxKsA+Z0z98Od9CMNO+D
9K5wUVDZ3vtXUJg+ObJ1eZo7YphSunEwbwFCjze95cLpMb/lDbjAumASpUkih1zk
W6L5JRMO4m0Gye0ffyxCS6+6ijOO/77N1s3wGbHQ61zO4bk8xJnh3Fb7Hnf2GqFk
byGExCS9pzoarsYdPAfy/nYqhEvQg96yA7BQaMP3jmTa/zIwgqG6RschCwgoUD2T
B8R4f41K6FyPZDx0yrvW848q/swPh+yCbL0krDbYQN7WxCV1wMOrZiwvHCcU+Dhq
F6h/3NHHXUVQyyN270JdfEtw0OSmDOZHMcoyBRn9ftb/GDgl8yqHtFIWF9w1eLOr
DBB6DF34oz0CDKL2oPl8CEwWCcnYImdkJ9JFm7yV/z7CnKl2FBI5THUIWrn2aYby
2vuq5yfhSb+iKCRrmpIyjxFJ5n4Pd8Way1HEqNtqWW6D6eRyvD7vZm0ghuCOHeab
ER41ZTbitO2Q0YDVFRGOHYiGc5ztbx8Ctt33UYnUDXX2w2YURmaK4N/z5rK57SmG
s+yC19Q6/TSsoT0FepPy+VnxGpWnfiZt4w4RAqUSX+d4/fuVwcJ49t+D5toOwwIX
JAc6afzgCUiAaHAuPZho6lsPD2mKeX2GsmTzx4Cn3kYsrsndO8J2uim+/O1YKYrM
M0qXuX21tPpTMjYJL99WeJz40OaZOuDzc7ExyY0GCsJKERN+48F70x1hL7IfbbLX
OsajhSP0+2M7cPWkkVUJ62JGt2feWffHG+8bOLW+5NBWuplzuEB4f2Hw3n6761sz
3q7/LBBtvE99lxioWs1ezrgpKt217xIjtwbYoEUmPVFBEMZeM2HEULIQNzmvoEq5
jGMvdgIHktBJLexO57iyQRE+3eeZ00s6DJYYJRvtp3+aeQDVA9Pf3DxjLeICZdu1
kBwZojEgx3HSSox4rZOGiCXD3s8B7PH1yGwF5eaFO7DSrD4wj4FUoXq42x9Fum1B
BO3PNX7o9NxaAVYtLgnlqUI7JnubeLIGRju/xz4HD6/Zw+U0MNOp5Y3GVM5CjJ9V
CYiRIWw5+7njfdzirToKpo3OvpfgSI5ygQ/Gvd2RyClV9LAPrcYdntF+yxIMXr91
/Rh/rkSPrwlauREzSK0cb8qqUZuuj33peXCLZgUxtAZBlTDkC0StevGKhHJRHeUi
v77MweBftM0tcP8Pu//q1mgMjNuixmi3vub42BJNKTADgyzfgRfzxsSPTBgNvPw8
GSzAJfV19k5l4GPGxFWqK+zTTM4GFkCQvdboBb87CxbClxW567Ftn3W0C8zp2YRw
f0ezqp2gOWuQDQeQV17lDTeUUJNx+s8cEwObDo7qyf3kAv+lo2aijMwLkFRd7mwg
8LLtW26eb3z/2CjelM52vfWfILaUX28lXyIldF9ZIW9GcYoeA4aLbkvL2ofCRO5h
HbYT0A9JBtJuameqBx25TqtxamxgbHZrZo7LKeRWwprus+yehikEVTlhLRmDPF+V
o317/jRGiGEmULCdThNo6kTliE1h8Lq8cN0EgIxZKueF/6LB5dSbYLRP100xCPcQ
Rlsf/jtexO6rm7eo+Lpg8SS/q4ktsime7axc2gupZ1dpcPmj58LKB24NAofcl/hE
G4Va+JBRO7D9x4worh73zCH6nkA3WjPsVe08eNYFYu0yPyJthr3j65fXF2oN1F+b
WIU+e6Nsl9QHsb99JxEskArgzKiLpBLiMW4RkzBkrSNcTwJDByi2y/7RBCaH94CD
Wt2lD9UXBToDoN/TB/JLzphfoqZhZwWuY6jbwJYzXYlpwchRRR+q9Q4GHFtvkotn
ZvphhjdJ0e+Cm/M1GTTtDXdk+PKIIdoDe8Bvq8ym23Q+QvlLtFEuCmUMJRgPqOWv
vZCXWUF5cZtYNLeKLm6370KlRokKOa4IvqW0/RoPBzA6pCY7Pu90urXcDYxfLNRX
bRe5RdGVXC1ZXpnA6dRY5TOvUcXpRi5AwQSw2aDDESLv4dk/rzhgjb4uWoqASZ8n
6tCyDAM3H7twDE6TDB0jbBIDgKwiePDkUVqm77cy5b0Ad81+oehtcrJtoRQ/X+3v
8G9FMg6UyyYczAuSNdpXukHJxn9KBWYufKkFPrsP2wbB54i3R4sH83b6ZCV19jCG
P9DhRD2Q2tYDmXzdYOfNQDV69ApUtTGGhueImEEOQPteRCnVOi+pJ10QCwKeOlzu
b4y5TLY+0mnJh1bOIJrkNge+TAX/0o4nAiHJZRFw2F/ojcDcINwqWP4TAeJ3Yuuj
efAzPZmZ4aaHSw0oT+wQf+6px5UMrwYj5uSwFnxLDtA5rKuS54VUtblI8mgWZnnX
sdsMrCVbckDDIB9e4be9zvttIM68Zkos6txRQ5uWWTwn4oG9GaQvc9cjcrbtUEgr
mqCewQC6CB9tOx+5I/f0mAkGQG9e+P//9EMnNWCMfqzT3rFAxaRz7o/NdfJ8wkiV
R3qFV6WzhN22quWW2oKjdm11TYmIDbfUj6lPIp9BGkCkc1zkYgZL56iTbWowq1nK
t4rjmkTM4awHflatEhriPCpzqkkyo3Miwc9JdNYK7V0glOlxb7t7O2+v1y1FPXnm
yyu02wfjKEH3LYO/l7bR8iGEescaoUMss4bPfDDTRjGonnlnSkUFLLcIPG0aLzdX
5yNuUaM22rKgrf4tSane9T6rC4/Xm33uxD+JQDTYLPX1zM+YEkhethrgV9VPBAE1
Jo+e9e4iodIQ0lxERBKnSHLvttMmcCCafZFngGbfkT5cOpoMoexzEMRV86BLrKZa
3k6pqd9bmfyjpm8lsnBZGMhkGebDExi8G6xMZkWT7W2KNXreDfvEyN+mk2NnG3w3
n1FiCkfxEpCOaIE+4p9HOPTKD8qOT8OSIbKiHp9sZXv4wsP/wtD64vjlnRKmXgD3
8CLt8CVgdF1EF91yOMVGenaRWF1Fnt2J7C57fUUD5DeoCJxe45ZOT02gDqf+rafm
8c7+W7RcOlqu7JoUTT9gLYaEFK6nPvpfBEtwUBhYRpmwogK1eWUSNjn3NltMYxds
oKIeq3T4pB4xgKL+YV0Pi00ZTxU0gZryiXFiEokWb7kjXqv99sbP1mvwSsQfU/Gn
6mVPtta4f5cXTZ0fDcUqpJQM9bCswmjX3eucjJXpj9i/n/eQix2jXCn93fhM7Xfv
q9mMgfdNga7woOp8F9r6Dre/YAmNk4/IhGxQcG3qR7rqiKzt2QpTLVZlkG54++Hm
S4bXWSn6tdA2XBEaoQFk/iGhYttajpbi5mk7G2q4R4p+Jwn/vorln9JjDRn3pqo4
nbZkLxp55rUsS1yjwrUdScnJgP7Jj092bv4Rb7Ap9oOi4KPFHws6wEZGdTfVR1uM
4eIzZN2L660t1okEyepfEeATkPf+VRMQzE7f6gM6Lr50LJVjVqavZtRk38fkEjFh
n+B2IxtD1VHmiIY2CJTD3oh9zO1GnzMDTdn22wd6WJpamE3v6ziwbsC3Oq6uCx+q
MA8EGzDY4+50hcbqOXnAcwhZVGVkTiqmGDhYVvS8I2SpwCZ85yN/7jff15PiGlGD
juuHZjyfLY4FooXdRZ/O5QrXJG9IrZk8yYCoSaSVjqQ7KnSSWZRNfpPuU/Qu2leS
Vox/iyshyAaw7aONuLAyVgq6NohhUH2loPAeDZcUJAWdL3Xz7qpY0LOfpQsnL1gw
qPzmo6fyp9x/sEmGCGi9j3hDv89WIm/Yuv8YYJDQ26GdbDozImrbrra7FtF0CKz6
lg80OrIj0rm9HZGCLXlQ9sxlAwJ53DibqK+lXYVJ38S+CSYr4TOcffN8osEmuj70
J8UMv/j6U2tJcWFQulC3chiR96FQC+GvnQ3bZaPuX426mGm2FdDEgTSmRyxJNOLy
iYjHKuaOGoDtbcoKdU6IHOf5cXJNehsTPN1PNDt27cKMaEMlo4wv+CsbFhfdyTNl
VlOEo9dDXc06V5jw1agTPaJ92lIvlQVTqL/P/ZcsiuP/jf6WCl1OQsVNcKpTj5tg
0ZvEG3YYR+n6FfXD24dQFVp8xwrGN9I+OmrUaXLeo4y/tO0/iL9+Tz7HYWcYkG7l
7RY7elYXajmWnzsIIHGu8Gl99jUeYoI309+Y2PygzMvhh3rfpMVRKbNd+3BILE01
Lv+Xvqx9MFG0iRbDmOXrlsVG7cqupMCdTnMmN0axGYnZqy6yLWWnrVENAw83M3CO
T6SCBKH9ORYbrOuy83i+mraJgfFc6TEOYStKF2LhplXdhpIjpeYb+WPwUsKrUPr+
pLcTI0b9mQB6Wwwb3PrTCD+sZHBlzH5a6p+PPvcYvqPwXZU+hokDub6Wcno9WTxk
yGjlhlz9MgJVp7r7AZGgAxnYNZXa9JJIEBb88p1VgTNDqjHF2dPh7RBl0r4TCDAg
WuMf+cFkO0gc5uMbPK2gSdzeixkLDRAgra5BsjEFyML4nA/RsHvPbfaxuhD5qwGT
4tRHL22tkGUMID5PjV6+hJMQGcYtkJbIOojZzYzOB+gH8iW4sggesTdhQgEeXX8E
cYKdWcWFyHhr4HqIhFQW4SpybzSzNvEpl4yIymn4BmBfLxn1mNtSQ1tSt6CptnKJ
IHKbKmPajn54EnPAZUd/Y2ZOSLthOBsiXLLUeN1wN9IdVIYfxetkkkRDGJuktN37
WvwIg5ywnbnAN4CXQQkm1/5UEF3laMf7JbJ94IBO9P1j4xJR7pHQuUEP7HosVZXg
nqfDfueLkxwz+iPWnWMln7uewcG4rZ2t4wCwQ7CpnRThL5cuVfT8gnR8dgYA2NzZ
ATrf6oH9HXwn6TUyjWg8/19aP2XwNzU6Qo8Vyrj0W0M4J3Kq2t5bi7jU5XNmPh+T
PGn4E+CQu2pJoNA8OM0BzySsf0Y4p5EK1jURqFh36FWy7HGGcNnQWx73PKek2eTv
MtZUY6/aHo5tcSAIoPVimRdAHDqmEv/+5PQk11xlHIA+VA4KuwxWvXQajIIWB1j4
DNn6DYMK1X+QKvXiYF5ZsQVbCrEjanQdUqQ0Ho5DpxhEvSnMBxX6LB0Q+P3eoPou
vJDRyOcDLQi8a+Dp08xadADoVIStLt7bQCLQtPaQqpuT/OnjwB6HMTjDIsU+aR8W
9OknBKXSsSsAqLQutsiIVD1qJCjcdtNT7OYEBusZ/D7pPbNQCBHiyNmdO9Ieq+L5
Rzeiwsw6M26MUDQY6jNCJMgYXMEvx6UuZGBt23N37MMxUPlJ57ZwGC8iTrFN87VS
JTB3LTZHzzievErC7KrEthqdoRoP9x5G24BYt0vzDccOuDxNqcZr04je1N70WS3B
ulC9f0tz3+X6KctmEEst0eFSGVzUv8SbDQlFXYIbnuajczaWpkcmKChCu85ixuwq
+U3Swd4arbuvtavjhqdEhRRJFaWGAk7O65TB7H3OjLJ6/32B7MSO9zsUqT2Ihpjr
qjYjFVoZQf42Yofat9aeO0Qb3aWbxSmi253EZOoY/8oec9G/Sp1/UvTogY0sAn+I
ZooqlQAq1opj7hbrYY2oWyG3AX0wRn7W/2nTPPBXZSc0QdS5Icduljqjahs4pOBN
xnlRCXEFxtB4D1qhab3HIaV+aglkAh/6khlbwvZPXKVCE5TVLwg+ezLhUoziwyhv
iU0RUyW0bQ/M5u5ZUmyyrLzd09+8yTD3tePLu/Ba/cLUAeRo+yJOTkokn4U3ULXU
m2ux0AiSG1XiMJHGxf3L3g9CadM2XxW+ic+REL1A787lD1YCg+LrLKXaQheV+MKN
95z+j1jp/CDRzdfUSD9y0KvvBvsnqM4IO7iSiW7IJLhFfYLIXN3vHcmGa2PTtVY5
D3os4+i3b+Dzs9mybIP7lPbTclJoKWRrjirtA3JqwQ2oL92mqiKHiFaIB0wb3GJy
dk0JBO5w6wtUPL3VmosIcmqrHAmQp368SKaMRu9spTow3IfUb57MpCIVDlrKfpGV
V6oydGiY+8FHGbdbL0ve3V0DI/qdRgkvEMZ7mRa61KZjjnI37QDpLNCBmWoSLGGC
xywlyzkhKKzlQGL0/Zx+7i/6c2VTQGaRuJ/iFuIui1b325UMP48qUolwJhkhS0+4
jjUGoxnYX+Mpbq/WkmBOfTiIEcO5Sk8DQ4L1Sf06SjIh5iFK09ugitKIpFeKLL9/
Lxke2vNrXjGGPSc7lzNByflgoYDYLW0P6XULg+knmClU7tDfWmE3O0yBRhtB7wLB
Sh23S6RgZkGdJ7BJqT5VYbSQ8O9FZ+OQsM+egg9CLx5DThwkkSqtouLH/Ns6OBWC
dRhmNTIAYScsr//9pj1mQ5NXhgC8ySWEJrA69AaqTs+FsIG0YLNPgyOjfvAqsSfw
uYzaWsfwGgzN+AV+i99n4vpGj6RlQa50HIPREYCYwxa9ph1u1Ucv3hSz6UJIsyJS
DGZqlHF4xUFL0+xdkcgL2+hmtRkReteziNWl2HaCUAZvPi8UcYzVhNAar8CHC+WN
pPvl+ct7bUP6cW31+CtGlGhiyfmjk6T9ot7k1v5NHllpXKwYOMYB1t2ipRM2hOtF
O8SgzLApiDeaOC0osvv5Z3skUdyhOIfwuUHyA83s3Gatcphjr85VfXhWRBXJLBkw
5Fg2phai1NAdNRVPGcpqt+6UktKPEgAgvAPNULRpQX3lFlDZEIKDZi/qXhRAZlm+
j2XTcSvW1z1ZwqpR+BiclCYUBjpK9CMP/rS3sdAVll8gWrkX42Uylwl6bqps7dSO
Idmx9fQh6wJVoGjO98iFCie9kTMFBl9grtapJXqXger/GjipjNZQHQajr/gFGJAa
cAB5uYJA6Wvqm8JomjkLp5hpiRbJ3lISzQxgHpeQBN/x2WNxjTOHZT4LFd4vjQXL
5NRrRswPKztYv8whwl6zT3bz4WwmYIVvJqZjDU55F5aYhBUdaOErn3bcZ8av0Sk1
q2FwxmbQP3FJN3ppx7o36GK46d7P4aGUF0UO5QeWmVK++pWBs9fEK9okADF0mh0m
T9tIt5GLji2d6fFsZOJhswWcdhZvcSj/eoI3M9iqh1mZlz6TcXuG92vvRvexmapO
akAOg5wC7IotK+bEdx/Ef26FQo2IKxR4R5A1K/gxIpKXqFAeRJjc0d9Qra0CIQ56
8Q5ekSkKcEaXXHcC3k+YKdkDMcTJyB5GhroqeuBKyidrMr83oZWQa4v8uHAfY0iQ
c5DDoN4QZMBU6wgp6HgwPsruhwCltaWQit51R3gShvte7L9KGy9gRkUZJa14vR7k
YIciu313StsVD51AR685k+6Ml7jCBpdqqQnwuW9D/hE+SJPL3VOBiJG1G7258Mxt
WwU+SeyX7JOT/PBatTLGObLffiysP1ts1DdURc2EI1n4KkJmvVm2r6tSNl/7hlaU
jsr+eojhC8OUG0yeNs0oPFaOvL4FdNvw7S1JLwuB/JCBaSmYlx78uN8uaooPZCsv
mUVzl+5wHY5O/0SyPyHBgUtKQzLHuw1yFAkqWhgWDal4Z0og8LAza2h+kL+AsHSW
obevosqOfnPS51hRwTOqIU6IT4/GZoolvadZfBnCFzYavLRWeZRiSzZoLfG0KPuV
mV4VVvJk9Dod2jfEm9nlUhj0cGCjF5FoZENOmcKlHqP0zm06R0IgtJpKg/XQn7Hg
gWBQxIwtC53WLCHr7fQA1vk4gfi+4OdBUhSfLbxtjTVkx0Q+D1BRpgd2vZ21j5h1
W+q0p1GquzRzLMOqslTPxZbx2dLdsLTFbtWbUaAUwsx8q6anGw+nAkhX3VANErvT
y0rkGu1eww78ng/Kq2napGxxtGkrRJOqJWv/PGC89oDvp8V+Wc4xE8B4TeezHLOZ
UDetHxr8C1ycQ6tMjhblDzEqeKtSfNLdaf+kBN2728NhEP0cfQH2DtNhth4vrOpj
3PABvpvCsDEzeUnri3N2vFBBKcXgalmK66sWMPRsuqoVRrsYzIlAa4Bw2B8L4QBt
opGCz9oVknoBbmDhDm9FuzHnNeVst+iBkBVUPJQWz4I7wuviAJaOzj55smeKcGEa
a7zC9PJISUmX4GwcB7R7CBI9uu0xlBSHq6HZFA96puwygOitKbXK2FDudRN2ivx2
FI/WbxWA1UGnc37+eytqFRo+oh7Fm11LI37JNF4+REw+qcedITzLpofT++exe0at
8c8N/IVgkWHClSeF+AXedDINM96Fl1lx+JZ+H6Ng3/vpFAH6WNmnhgaPfjuv1N7h
MYoMvVrIqpau4eMruN9P4yqEX8JMO51Sx0zLLcCn5nMwLIpVOmdJ5wQt7QUU6sIa
ayeNS9QAISXB9YGdT7A7cD0qLa62ihbArpzrhb/mJU743IN8sSZPaJw/2iADzVwz
RKTiDG6t8TpP4GFvIxQkVsyVeK+jRJQM3AXC3kJSUYg/SDnlwP4EHKZG8dFxHnRe
9pde8D033Tp5HMESNeaxFgoO4hjjDBNhCsNjWGsYNa5rkHXNThlFN5rIRWYDF+Iw
V8B51OJpP0Zz0S2ChnBCCrPkp71Rv8Ug4TXCFo8s5+l6sHEUHZIj8gcFF79uutjJ
gcfKyEYzWam6UOeD2hJWT7B2hjcPqAwz9RMgK/mia8mTNKZv4L/2SDru2kRI0wLR
ohpJTym6DVRg08KOaWgoyphvfvp1PEDGIiAoNVEUVWhmDUiMMkrh0xgrm9M8i9sD
MV/OU5JCqKI8HcFLEzSblf3URCncZdO1gt1SyvCUh/inkTcSiLRV4guzuJzEzikz
eSd9556/WNXrBwieGMZF6AnC2NVE6aCjjS3+aSTFhCZzN90tuCJ2eIE2da3XO0Wo
utZprJ3qBnd7UvTrJz9EfTQw4VEUoxn+0EvmXNRJ/GRByx0uvRazCkXJtdzd4dMt
eOtvH4W/7m3t8XX/SGpwJnJHxDKaaSqd/oJo+2hgOtUNyBisJFghRurL/daoXY45
kbrvUxqKkcNlie1MtT3Q4RjlY5F0jIR9wjFrD4hppw86vYtpUUax0asjp+Dc7jOZ
N5s+8R7CI7mdxj3i5i4vS3+KoMvlMse8HB6eYax2w5lZttIlwPrgHzQQhuTq2ikO
SMsH4fKktpMjUsDxw6Yy8HXN4+bN6//fe97jintD80fsCR3H7/UhGRY3zot78XMr
gaQcORPZVJELAreC4gFQQK230LVyVMvxutIVMphci7F7ZF+NUnzas+ZM0fLakJ96
zg6d+7tZCHWRd4HK7DVsSvXWc+/bi27rHlfmFxcN8XXb9mQoIZw4jYu8xNjn10Mo
3wsH6CsQiBdDGzqbUqMM16eRXR+YMKs27AXy+Mo6Czhp4hq0d6ek6I/nUlKqVCSX
xcEuQ5C0vPIGfwhYQsC+LHiLXSYpLIbCl0RZBe/8/BjGAG418iPYzqz73mkpOvFV
3Vcv9GIq9XxyoRXbUQFq25kkgbI0fDXgZ/RAqn+UOXY7z0LCKfDOQDwrIefwRq/I
xCZXiSXRiflekXsyiTEipqarBtyy/jeHonanCVXHII++FU8YAYQ1OQrJPQk9KLRJ
k63HUQnYRJ62fN69qRea+PSO+oqfn3dfyR22L6aolGcj5aaPp8YOmr4mTZexbpt6
GbQGALqPYm3utddnzaiQ4F77yKumdbK8ReLEO2uGffddWAFBWVCyvJnd5QT7ZuZi
yMCaLN2UPXdeLE9WP3IPY6Kv0X9Hq2XzcfeyMM0skbURphtlI3b5VwS6uyL2bla/
AbEv4tnYuDOoIwvVwldwDJkftci34DM4TOPisS6ezI1By1fm/mHzPw+PvOXiPLWv
RSBYnFxMiGd2L/d7NhkVtBXiUHGOvpY8k60FSz8dmPjz43uAYSj/TsO7OeYfuPMA
wYGo4sktDrr3J/mQVNYmINhsM+t6jOE7Xo2LEc2EFQH0ivuIqwb5WKLEn92yHqxg
ULR6tQPozmT9QKYxAXgI7tsPBCVQSn+LkVr/Gd6xBszNlIUhz+JC1PmE94mZG3G1
d1uJG4lkPXHT+RE7LnjJtDeYadJOrJYK4QR7YliElZ+vu7F6M8a7rFpTiBddjYoI
iquM74kuYhcjcntnFTofJpVXTGJDNs0uLwPiD1U9UZU5YQFVJxZkxf4AI+aIlMPn
CQ6XL6kFop+RILd2GbZJ2EtchgoYxI6hQnqj0fXJnuWARuf/zIWxNS+sqhoGRwio
AoEykkUdrvM7JpjXSCGhowiT9aYDWUZJ9S6yHOk7gJdZ2lrP/6HkwpPRVfs6GgYf
tpUTuMJ1M7N9ygQq/cUkmFv86/VDkr4RCupq80xRjChSvy62gM0eg0UphAAFEN2P
KNqiAx2NBB+pc9fIk0Jcg5jUZxdUpqgWQ5FoZmrNd1/EuEQDAs5yXR9rpaoVFPo5
uhKqwZfbqj+1XRwRt94JrHPX9ftnOeSuYZHajkohpG5Pj7KWJh66cducbrFjnlN7
sICHgC2OcRAKBxfSw5qIGUxqTGktY1AgxUynnwqSIvr7VRMvpTsWN3gVFAMDUnYi
lLVYTzNwUuqzvfL0b9wzeZFVh+xXcXH6bH5ftJ9UZwUNoINOYIieDxZysDXG31+6
R1GrUV/k5QfnNoWncfTyd3FlngGs8ni5F7Na+Mspn3hQrXzuUMbd3fnoXcoLkvWo
2nf2dpmN9e389GGNZ6a3vQR/3cvdsyIi0oCKBjJvGJKgCHdg3OnXU6QH3EUGXZ76
u5+6TtkY3CR1/5Clg5E16L6W2KwUXlVxAeS1Abywm53+OdoSI84UMpQUFDinpOkf
nhLbvrjUNbvUC8eP0cTleEWayZTAkxgQ4zJllA/l69JM8Qda21NU9GIsLERUVdVk
qTo9uZ2Hr6U9V1VO7t/SiAx/1AIWLwvXohk7ZeJehSKqk/eF3vwzpvaJSICZmLBx
VkpwGCHzjLQIaHS2hTiwAmSC5TV885jA1NrEfuMzCzHDo6O4+2xDkmKJ4rLiSN7+
agEqkyXYNi1oAjvrzcD0/KAj0dCXjo6JGlFOEehdbpP3cMbgrLDJu9L8YGHNWp4u
oM0NSCnASPvBzuikmd8ctPynrw3HvTJ+0auzuqiPs9SxtoWPp4EDrGT5SdFouMfu
6FWjEelZDWUfdioQKSY9uUXQXZ2TBy8hjp/hyCxe8Qq6XQYKcHLrDlINwBrXC8W5
tCAbACQckLx2ENCtgQeW3rZ75xpUIKJpDhblgX2Bg2thu2p9cDkdu+f++hiJxMtF
j1z8FMtOoiEaHBmGq9Uw9Sfdt87jubm0oD0ZuJ4n4RnTvaKA5eO04GPUHsCdhJNn
TBwCIe5XdqJQDcn42b8TFiEWKjGKxilYOYVsvKAOxTJYw4c3F4i4zsFWamZA5/De
SfE7CcqVti//rdxGkLKPsItPqSWjI36F3YJY2+yp239++tRGsd+0TwM7JCXBYcql
OKb+TAZOHm4L1fcNIteDTwzwrUFkoDKFGnLX/Qaw+FGz6U5w5VBkwPy+miTtnQ/M
T1gIYocj9mE8HVKfOLPO2F+M32Jx+RMgUcd3zLEf7AVMk2nMnyg9457nIDs8na2S
OM4odSX+4WbHYlVXJGC9/kPH4q+sjsKkCh1d9AAjfA78REc7BZ/e3Py1Jz3tFIvj
99oArat4q5oL6OE5qbBK3W4Hr/gcQxvTdtr0xTIGfIW+PcE99rWQ9NyljgJ0+jXF
55QmA8ps91bqbJ177BgCDnHmf3MIeyls/H+PC+w8l1eyagdb26OZZX0QXiGKHjj/
vTwcMMFilO+lulC84X6EMJFOk5msLR1URWfEsrLZETe2tTD7fEQcz5Whq/LAVNyy
aWSmby18fxhX1x8JuvWJRIAtdKMHjePX+Xcq2OzfzeN7dPD9zlf/v3iNFRRJc0ne
s8wzfOA7bTGDIHDqhc5VEJl7styGCyJP6NG+agzdrrPWbBHt+KN83jGak0ISRgwK
G5STaq0bHcfyr/UDq69tqMJACoSxcNdAu/EUG+H7llqpO7UA6U6FxDCjEmbKNbq9
aHJ2XFkYOcvV4ecRhwzKyQEkw6YcEJm0DyK3XpBWpPEum/LUfV3rUOYj0bbyBtRd
39AmhB1Wqq/L58Xr8b5RKoO3ACShqaz+nNYUEFftA4uOZ5Q+i7n7Ct1Nf4lDwJa/
oKM5pUOSKPeGoKEjESq+IojZfAwixkRAPOP2QQZEWER810zmTSBDrN0t1tGZ106S
HP5YDRchWdsGyZWF8qHuAMob6KCm20rsecOjCntQRyseQzfiTHV3CHqQUunJDHLy
GjXQb5DM4eFN6s6+tiLBA5i5/LuFdY8vAXJv2fU1amLhH1Jihwe0oiOL01tSY93B
Z09Pm5p8mQcs0bac7ZflHzggcj4pKl5RnLocJHgzjyW0/Ys51wySiENeadvDd+PL
5DafZHQekFNOR9rSFhlIv6stPCAkq2r402T/JM7oII6gdi7xaIi0q/1sDIW0MxCP
aUGJ95tozYppPn2awNNmyTcQf6MyVXFW3k2AWAFaAzeR+gfH26iEF4YR7jhc8OsH
Hn79ybhL0S6Zi9inEmX9WHzcdmXsJIXGrALTRdGj0cDWldiT8A2komEZl7oeLxUj
aNquhP3L2+Vl80Y4zqwN7qOkvB8SjKBFyWqRIkhNYkFxNrJXdI9Ay7jsyNnyg5bz
woErBv3P2Kslia7VLLE6GHQ2UueFs+4hR2qo62hwCIPCN8oh06otIdqwl0+beJIJ
YG4lL8KTqGAYKEIzBobEPnebjHW51sZXRJ9c1pAnVGwCFPJFh+OUbYxv/PntE6Ly
QmTLbOhW+dWfaC/9ZjAuLc2SmezskB+mQB6lgxoLUgCO5njaQJgM6TpFc9dQGkc2
MTo5RA2adxgiieLTmz8BI6xaNV1eL7quHrbuuw9f6+oxUfaZOWiW527hWIkJ0llr
peCwxmYcCk1iSVdn+dPoPhFM9SJ91pJdXn1zerLDzkoEzmKKegULmTTZTYmOuHLM
0KyWhOa7Km5vdByf+YJCqtfXdbHj8452rg0ESR5asvhIX/w0t+eYrnALZJPUUisJ
Um2zts46BocbHu3zEmxjGQ0Tt83uf9rMcMKLcrMyTx5UwoX8JRg2G/KJ1yhY9Evm
kdnir31rK6lbWVpfUPwqAHqqZj8ZZUXwfRtLLEOUnC6UrCRUOgsYB0lAehXnAml8
hk0kp6PoUZa1Z6sKQk5xZKufbZ2CSwiLC7YKK8j6SPmwD2DAGTOw/rd05tTsAZ4t
h4HGZcyzu9SLtVl+O0S/YKRSRybC6krg1q31u+UWv24QG0b74u9cvDGC15pkitU7
F3+ushtEEzD3QCNIL6n54cZ43f7JMRp2QblZiww5mzi2kcGOvBecQZ9rMToWRjg0
SUAg3xuoWnUzmR1mvw9xpK6uD8UrBv3tY7V6L/dR0c7so2FwoyROUHoiuNvUPOHN
hoZ8I253pf1m663Jwkjp7E1TY22gkovpNBjJdzVWyQtm+TIWwudjkJYO7UtRUVER
aDOKk+34wx0U1BxtZCRQ6i5cyT3WOzR9l+BQqIy8dmc6LvbY4a48bY1ULjje93a8
5lKCFq2EKa/woK89VjyDiB1E8PuBsf9yNwMwFco/ZZUTAVdrTLu29yorRpZfr7zc
7okUsMmtCxc1TczfXmMEkkdII/OlrOxjAe8Un/TO6TyYraoajCJ+cMA2BVc6+j97
+nFBgFKU/bVfA7kk8RAYgtceW+g5n/dNuhfn0ZtybaONecL67NZvz6iEtWcTtXti
oWULBryZ2xvzqpahjwnKnWwsuMTefyUcMaq0dWMQd+FGzg85B/kQKONX1P4CbgUJ
Ykm+nVHI/gbcDCgxp3aNxxWQ+ih52dcLytbp4LMV8NG24u1iUJVXVvbPg35FvGOy
wdopeGW2Ehq1wRZb0b98+A+rqWrSeIJTNEDam1M/560gidg8rpxMx+NZZqi8kphW
R9dqEByoIDAjTqklfeq6N6Lp1p8TsXeiUi8o+jjrps3k/pHn3cBY5mwBog4jlIrb
1OA9dQ3u7PkeVhj8nxEi15SYYFtA+hqv2A8oCkd+8u319Kw8Af2L/ufmr6eQZau2
NgyE0zdnzy0XYS0nho4cWlsKfJqgpL69W4+/Jrcbtn8jaySRmskHk/gL3+JtoEfC
BV4nxlHoaLtSkCqJYy4cjblKWJVDhOEsoHSpEyG2L/ADeB71aGHr/ZPPx6ka+I87
ZqEKhMzlzfChYTRwEEjOtlsz9LzNzvWXdi2WGfRIS7DxlNxkThsVVO9ZsiY9wFrN
ofQRxhw88+5f11Q2zca31fXiCN61Nr22Gz2+e7L8RZKvVqMl2aAMZFufofEfgX30
kGZL9T8Q9oH9EZitl7mV2y2i1F8hZ/jLRsKqIy2RSbtHlF1wnBfNUvFFb9JbWlXQ
dqIUrWVndnjL1q1iRvRnVTkyzTBPew6YyqDnk0X0OX3W7KBoUUMel/mgq/Bwodfq
9AKUpULHE0OyR3kviCpzOnxo2H1GMNsotKpUTHqg9rJaevYHjW/Oyu1x9PcHyO2j
kveBZUsa46VgYU9gniCj+AJreMt73njgy/TqHVHr7oskTGvf9eQ14miXL0JGJZtz
rwmD1DiRbw3Av86u9pGvOZDDrWv43j5a8Zew/wZL84oZBd8aCdJEUxB4WVaBovbh
LUCjQ/yUl7lDtUWXpSLLMErr9rv8mSp+P1IrwrTFpHsM/BgBzRY138ExYITY7v7W
UwGLYpQnLTaIAMKhnZiVOVjtWbNdiG0tjqN5UVUjY0ZLNsCuEiSAnkaqgVI/4kqC
IDttCz7YTSoE0nEIzzm46cUaFTCe4BNVWu30c4N/11+LOBtypeB+dM5b7ELPQPMG
rkMtHLLsmoTWeC02TGAdsSU0DcS81VvPpUcEW1ORMc7wt3x1gliB9RMyZuh2Mb6H
ontczDyvCpUHDjKV027VW27a6dsRyjwnuSqUDD3gWmbFA4+hgbQwWGI8pJqUtVp2
WRVUqscAUQJnDosHZT4p4TjSkM6HHzVq/Ez2E7dg9vFEk6j1q8RWhiPjwAAZfM52
I93HoyoTW5vWJa51+opMKC5HO74N+WSFcaRHxKC8fQ/hq13tG0+02/JdP4+7cUEt
+XQ7Rcv76Q39iuWFS8lZkHN4X8L8O2r9xGFXoqZxUQDOtFBIjRLra/7KnEisuUBg
oW/t4A8fuJjiaNHQKxv595diHfcifENlw4gVncCE+8tmholrlOQi4+yo+oXPFFHY
+JKmfU3id09NlJbdLMvcgzBCx+szOtex4QgbINFJq/EHVIewvVXuN0d+9YQegGSA
Fd3BLIN61V1vXk1LKaqV3s7V1W/LtmVbcS3ZfPn6R/GjBG9q4XPskGeyU6xOfvhh
pGrv/vXxB43gKjCcoOVqBLqcYW+mqaMzzzgqHJlz4JcdNenxDKZ0xLodx0dqxeY3
FLY01wupBAK873SY4ns0/rNIZgdRJzC5VZWJEDxGI2vL63uC9P7ySUkdyyksBGAw
p1+x/I7r8OZdL25QZ0V6aGOMFLUnC5vIQY9r5K71XlXxUfEsdQz3e1PorVbxRZYo
2/2c4UREoRR1zdScgc5kG05ON5izsVhpl5ggzL/W/2vdBZ5dMmWDvnp0osQYw/oz
OaaWJdFAoJyehzDDWYAicNvvbUOoZ5VZdcjhei0cYfZH5MbDV+mVCx0kNXFJTP0Z
CvWnY6HhkWYC2M+jibSM6sCXVIS8AQ3h+t/oFKAlRrFGWdOlDF+L0mSMqkrADNEE
HDh/EF4TftAnpECUzOSAplyDS9y2GtvAC/sUbN/LrY43EWoQ1D7YDN/qJFAiWU0j
tBT0FzqInjaXIL/jUZG8FVK0Awx6EUvqhiyjf6r1CeqsquK+dGZ8aZRD1ni7wGJp
sclJGp6MBjKmDgWwKyXPlGYlQ5HtviiDH8LHuQnC2GGWWrDmXWlfjTQSwhGE86UR
hxgaEX5z1sy1Ai5rj3zaYTivHn9VEV+GRZMIcVGMul6s+SbSDFaTZFHv9wlUZtSn
X1PJeeyu5biriorPDHZKSRqxz4gxGWmPf/XpCm8vLOhcvYZUbN0iHPgwx666I/sb
WHL5sx2Ic5IH5bZFLMtGICM1g9xJiY28zrY/63CjONIqH/qTsGzQfGd2DANhSP/4
k1w4c/z+Cg5b/Llq387fkTUh0Q0VhSROBkeDvOxSwsMxOpZXFCQV5KLkjeQHyGxg
TcdrsPk+hIh2+wIlvMR2efTyYVgwyCnPynMT6LYlkGfn9/FcGMNiz2UwLKiOH6vR
W/YC13Bz62r5inoiT9fOUiu9MBs61HC1GXNf7a59NJrEwh0dzxszh9bxe9O1U91S
/kiweUI/E5y3ISC7ystg6XvQyzsXus4BlzS5wS0DUaeC9dylGFXICLp8oDXC54jI
QcUQs4ja7gIdm47XAL3wk6e1eIlXirzulE/u39UqPfxJbxYIJ8qc57TfyHkwfm92
pZbDei5wUuOK0cxERCaQY0666vwtCN3EFn90vRnaPNhH6xJOOHYhTlHl6/6/rkdm
jRghbhenwrQSTxAm6vc+WKIl1UT0ou9XpQPxFIclfZARDZ1CmSBed7tkNK/UAt1d
bRyvlnsH9X9fxq9YxQPKe828xxDkmI71z6ftz3L51tO56aKw0eeVyc04+gMcZpVF
c7tz6hPbJ78zQrocLFDEgdhxhm/H1zDda3+lXz6HMF4wYOp6cKLsN8h85McJTEAi
LVkspnOVxYqWr9jy1RzDBu6s8S9b4GlDF2M8d3whN3ioeY9+231TyPEmxb8syEhX
de39CH5srOuWx+qamv4qFwX5Esm3Bf7fFDXretTbreP07W2TdvFSziaCbUDXnOZ1
bvx99b9TbuUwu5wEpy7/SROWEPsnfQoULXDR5RchJKym5rcLmCG0ncTDKJHcc52q
XUbO/dYWUJG4qzZgozUt14qmooA1UdWWDh8g8m4ro950HljqfraLD55tXexVUOu9
m1GHsFSitkJ/kZIZ1ZFdaQTyP93E020jgk6/1uWehTDVPkHCqUkn30e+ol5ZurSm
alfoP4sT4AorRzo9QgLazSk8APyUnG6bbotaIYST1xTSNQApa520V/zXlkR7ZIIP
IyG3J57dDpLA8RP8gMEHoa/K3HcyIwhmjiHzYOzdCdH4/M0TsLcRWbTctDqj90hb
9fVHgsS4A1aU9czJZ0Bii7MSEyr87UtQ3Cq8dG9yQ6+Ab6Dgtqry2YbNSk79QsYl
x+uNq7/bAiE9yU+A/44alr7Z7vcjeymUbzbowcmE9wqd5ByRGBjnApG6uIC0jgup
u30r8gGqZ0U7xo9pm1rjmod9KHm37ueEqVoWBuFQoDNU7slALVm66xZFHn6WGTLF
3gYiXx+C9kAUtfV2DW+y/S3NhAldf6MDykNKpYZshQrOqw2WgoRdGXG8eaK2xOKl
OwbvJQxhzy+bYoG0K8YIk782utdi4/19wQnqUzD+qfWsQpa3ZWM+bqug20yzzz2A
9c3iG/wD9QhWVqL76UPpY2Wv+SX54kUKid8MYnaimDzWlqJpaZvWekoHTmTKe9m3
3ajTlLb4E1lbY7pvWNjGXGQ5Jp9z90yUBFQkO6KidI5c4h2AExXvZfsdWUYN2NYj
YuMG4upOfKcql55HYTC9lBgoGUFUQo6fYGVoiwSFWuCKaGmGEndChm8yzvlrIBbV
NwjV4NVpp/XSlXuh46CcnGmXSgywR+F9laalN5QeBrfKgSpO1kOxZ3coGbXQvMv6
yaxRnIvfNUq5Nss5W8aFm8drYuNQ24ih1FTXXUX8EUi6G5iKdphjDlxO5JldBg0D
2FqO/DHScEA8suj0pjHUVVPQl8AQm0DOxGGgDaXwoDbKsVJgqFQgqRV13Tl1xg5D
cVZXOuNExxjonBgDw3LEfkgPYxb3gCYsWfIlqe71LLmBlTWzr8qAQQkSVpR6S2fn
SYXXpkl1ObSKLQdFveSwCLHh0RMg4maQRUCFD/nT7st1efjMrm4U3SnHbqXnOanO
/NSTqjYTJSssdwS3pGT0VxoDybT2TnfYOM0kkPKy8E/kv2RysJ7UJt1RjLtlZQCr
iVf/U/lZ/NnlUQNhUJmQfGpJjNUC3QMawCnoQvU+TDekXHihSxSDERBZqUPzJCY2
lUolnIjCo6IjMT6qfr9WIEr3Gh7MtmwuhdfanVHSWH7EF30VG26bkNxr7voTksU2
ZqzeVXYdrie7ylsWskub8Sea89jScP6xMtG26jV9o8Ax3LB2Bv9foMc9oB7L5Wb+
ltbXnkYeCwHXcRB1bDesp8o/zYKStnuRol++kNKqNBPvP44QrFda6amz7EHRvv+i
S/K1sjYddJ5/Jgq2OvNtoVB46i8fKjNqufdM45thhgIPWA8CmEy6kMA/t/e32Rep
2E59IuqPzGfW9X2URsn1LDsXpMNWwaIL9K27dnVyNEWpQztKe7hO0IYN690aHNzk
cJS+EYIvKDFggCVdpBLShfMA+6+BvspsMK3IwUuoffwSKXUqiGxtc5n1/fD6M6tu
iGXGGllY0657YMcUmyr39eMFrs9W2w13d/V59b1+vskYMJvDBA8vJoP3QWRbdGXM
d86xYpDb/H4B/D1mkm5vVYWIBS+a5RijaJryjlVJLgAEghre+gYV3KFzgSIID422
tnPBLfloi35wfC9FZY6t/jFTh59xZE2R52pA+f6moH9MPeNK+o34aZkryufJ7nBQ
/tmpSIdx7b03YCxKWzzIrTZCZMDsn7trfpmg29BZK+6I1LZAjdYoTnz34qXrPaOZ
mtlGzDjcFEq75UtkfV9rsNzExc23SkbeXbBWwtqzk/ospWNd58w4Q70oaZmqjLxY
hY+OZjekTAGXCZV3pRL3lWxRAkknuPAOG0IvbNG3DY+Q1dNotFVSrIcgr/JYc1Xq
XcKHdb3WqlFSWx6DF3Dv7Np7i0Xgt4SP+ssfdDE/gs5xnYyTIhUy9BAM+4d1yVJm
2RZckV+lPX9+iHcK3IStklSj8+2hR1uG5HDxi8nhP+BCQKNaBDazYHsof4GrhRrH
TeJNBVThTyFC6oYyNS9uVyDUZ5w9zCOPE/EiR8QUCWEWsE3bd9jfx0haM1YHNopQ
qkEdrcpb/uaYEsx/JH/BCWPlb32iNjPI1PEIICBnG9cNPF4Bf1s3GXfsxXq5S2Oq
5n0dZs50WbHTjiJSLMEDX18OzS6IGbWRvqhvSTu5D+p9/oyuBXyPDj0fg5BBER2A
aXaNFhXXgxXwuZ3+MMiBiUgHdseSrt6voo7fpxAtnGRk84He8M/w1J+r0/98/Iuj
hJJGQscMcn2ovvJG5tt7CpVI/CDrhYa7c3OxVJd01VEwK2uBFNcFtmCodbWWAQfG
a9Vu0O1xVsXtIydyetR4aC9PN/KRZnT4BuLKzpcRRQO3OvXgdo22myQCwb9bB3+h
/lUVa+tdPVQ/BHKAvfhHn87/xIM/3i0oV4CTpky7dWZZIjkShwk1g2h5cd54RWCm
5Aw5rL/ETGJ+w99vGgR90/p6yHoSahuRQRJWMvrgcuaognkZCWwgni92ue/MDf+W
AKuVRd7y5lguhZ7g2Ht4ki7qiugF3sgxJwg8QjVZz3Gn3paqM9AHYVwpufU2kH81
5GapgncBP3OTWZIX/SlvZ4cBHFSAWN/emkGQQvk0uXAFA1vtlpqAzx/iGTRKokm0
WUunoSTZybOb+SISpxOY2+rHbMS7BW+EZv02ytQttGIVjDpUptJXJHnNwtvWTkGP
J2+HzOKFhPj6PtWxH/cQmUkO9PbUE6PU4FDQP/W5G4RYJR5Ama/xC35CJe8jgxPJ
4aVi1dVkjplRVNYgT6fMkpDsPkhjU1U0F9t1tcNFVWWIBd3WgXMSeRpqU/8MuNjL
rvLl0idreGXSfsvVK6lUA8P95SnrvFHEcjNv4wGqIMHuHuq1I4EQc3xS/S/vchfl
INkE67VFQDL92eoH7MKaAZKoYE/6QNGjWRbNRbFhtd/iZ3H/wEltvNUbX9rq6uwx
l/LgA6q3SkewIl/bqaR9Obdyrup0f7pdpKxVDYxm28xnQsHkNQY7lw3HbUW63Eii
lT7UbipLl6m++igg2DTDsjtaCFlucBtRX6WUJXjhzslo4YfjyphrqomWF2Q/IQYi
4Xj0QbUJh9ifdzFkz3NnSHDLbH9JvjATev2HUPiXBgvni8rJ+3h6wrTSl0t914/G
zlaVZOAoCTix3plRK9cmzOD91va8o1ryI/zOclzpSVx0gu9/mNbHPYvU6ijPjT41
b2fMthNaAVu5S9GVgsMrZZErxGLUP3h4U8VK+421Ds92HKFJc3wGdQ4Q+6KYraNj
CxzfTO2KI1+hrjuytrpxa0DLHrqftQaVaw1d5bveQYF8/6xBcxNEv6KzyVci+3AV
PxBdTYV2rOclriWYcqGTFmpepqw011ajv+e4kQnegpJoqkxIvUgDJQe1ITYUONrB
th9TVB7CJAMt77OmCWJ8gmQoLDWTHY0jlicyKoneSwpIEi/p35DzAGnfemFIkiZQ
8qt+tA5gQ4m9msU+B19VszOaDQ1jBTJBPKerU2dNC8vN1+lvYUST6rhl4O2j5fyn
uAUL51/PRiz222hdcfaTZPXsokQRKPYrSUQVjY/Pn+rQyowgZe2Bdvkuqsrjkqem
iaNYcB3hDS2CLoGlj9y5RyAK3n41CRlcULTmCyTt5bpQ22+FiUCLEBaTf9+WQFWG
EVsJ1J0BTNeDM4bFTapCtsy2sMrsBbxKH3nLhDI4yu/CH1JaWKE7TiSPJ+KDBPH5
ufOhmxzbKWDtlvwxU9vKJzTStOWx2C4dxgTxdIQlM/69PM5O9OK3gZHdkAMYOaoD
2s2JY18nxdf73/yd0acSeG6WFjPVeUdwPTbqxcd7Eu7XpmD2Bl0HXss4407N0YWF
jUxQrffuMXyZhwFMcr7A2Jth3KmPD3eqKPLtEFw3M/DdIYZbvCgocqVRKsJbsd+R
6tuEK3Bneg5T/XZMisrUIVGkZyzMeucFeoMYWQ2i+khGH3WQUen6bmOvey53rvX+
/tiZhz0zcQGXGvLNut7k6A/ianRNo4jZh2uusogq73YYJSsWd7t/O0SaRIf3TuM2
LaXNh83Rj0LxOk9WCq0p4ib5XPvwCJJiOxTgjJblPh43LLeI3rDja5qomyEIMccE
+1zVdHAI9MDHDLWIy+3RWvnhamOjKFgXkAeh4DQCZuUowtIeIHEbbAqyBVQSE2pw
fcj9h7Vm94BvhjuaKssYFRM5Wbecl6QFdNWtX7fWYCb+u8Q7KB64DbquuXX2qAgD
6NKJgmNlwxWa8CYshC1lpfUR+CO0s/LsfOSDMtub+12kbND7HXDfgpW04aMf6dHp
AFNPiamnnVCTRPbW8VrwIa5oA80S5GRAAuRUKPQytQf38GyCjc9gRKF6KauNiwem
dqVOq4lWsK45mG7Kl9JGWHnaCQedprt3R4A+CYnmZQlubW80gGEjZtjoeyp5CGHX
QivbfhnXQZ6lygAAj9L/KwL/1AmStwgrPIzYujqKXFpHO3O1vnVvBzDtGRIHKyC2
+NfV7rH12XYj/OaD6EaOCDgi6Cqji290MLfhcBmJacQSjzeCXNqTTSFg/Bl09CrR
K6YhKaKcdpaxhbWlm8UIbexXZlKlrBoADxwB28w8mQs93nrUrBP7SnJytFhEiZgQ
JfBxorqFYWydXUuFCwL4b8YDH/zIK5qyfYU3cf8EY7on+wy2SSRuFJB8nFxWpCnL
nnDYK/7HO+Gc9QxKaLxSvP3X/eW+YkJPKVGXbGdXGYp2B2qN5GT4p9nA99/Jdp8j
BS+JqdQ+wfYhrSjt/Zv8ZubNz8qQ6g3WfA3xPnfYU6LXDIDgpSvv2ZYy03ue+NxS
RlF8Y7Wm1AnE2D0Gx5hjlrzlqg8r3CD6IJm3sBc0zlJZIjd5NV/wMrjJgxd2CYls
znoiZ+KL3xJn/Evi/0q4Wh0w27VXHp8pESsO3KbY1R3Cfi41jJx85H6z9DEsKGMy
6a960kkbOS1ApP2Iy/OQ8z4t6rXe/JcBdSeZq8Vt2bRIO8Pph2Up4Gtkovcmgu52
7ZJQ20EDLLYwB0S/f281Ranl2Vqk4HLhDros5aK0isJPkIYaxVr+RZFvyvEOnTzf
go6fTnjlckitAmcn0MR/2zjTCD49B8W2wd2b1U8XM3bLXH6vZHRwhzZKbNYUu+bb
bUVeyiREjZtffPmpQ/sqbN6dMLO5LGgh4qOzqqz9/Lq0gH5oLsdcqWFR2U3IqBS8
XzoAcAmOprxEmvSIUsMa2xi+w6ca1/PhKLeHnb2fXd+ssIFWpQr2n+NpRTvPC00q
/aIGJnt1/sVlU3xLJEbZ3Jn9tP7WntwefjOjbxRIYy0CFtWgyAs797hERaRF7TXF
TtRaJbNEVdPqe6e4K2mjyZIXUd5pJjUX5cFB/wSDZ7chJpww53avxU73NpTnot87
JabLZDNz2EJAj+3nS9Sh40cbEZtFYvcJFTmYOdWTsAFpmY/JvRpjd6WTOd/cMun6
AJnSYZxH3mjI14dZunO1Zg8zJC/7Y2hZWO5BC0OwZ+TrViqCjVF/y2LSr9YgWSX2
M3VWdkCk+i3Bk2Mpkl7gaK/r2NWKDnmYzGunJqh1NxNFvE77/4kW00Nu2hfRyrbb
i2Z0RkCDo/f0Qr1kuQH9w6NlWX6aaSzFKGtNLQvqrmc4QT8cU/E0nbH6FBXZlUlI
6puUj4fai8ypmCzzByD7mG7CdrOAuS1kEVNA7cN/t2jnTCmoNj1aoUKQIH5jzGNn
3r3HrJ+T5mD4D8v3Wo/RpEkY2ErTVQTOfxVNkFWZ1U6ojCQqG+JGBRC+Uf4M6vb9
IbHtUppawuM6jwFU5VodwH0V3dJLcGYVnv87b4nHkaH+5DllGaX472boTSV4TYrj
T/EoALzmrvKZHX5CjlNjGwoZqtN9j/baiWTa1LKtauHKkAC4HbQUANBSFh2Ajn6h
9gdM53ikfYrv2v+kjd3+/yZMxSEa35zSNeN3aT1UH1v+tmHOeOamgWCu96rWqJ/8
qR9XeKSOtHMKxgn97BsMNRqsu5bAkh/0ZniWG+P5iQVdzecuJf7TZxLNaET5wxFE
gY3Jig2ByH5OxogdaoW8Ik2fErHnJKzdxfQ2mVUSwLQlh2vNH9ee+Lk8yzlz8M45
5JhG/UnM53oKCDIOdasA9brc+mn3AtDoLk0+WyXaruleA3YG73ZOF/jh2eDo5lWt
OysHXqiFFVy41Kt/eCQtwvBWnTrOoqVFf6mE4qkAInQy/UW64CDWCtUM+QwTDm7r
Kuwh/0K0Zd5XvQQsevpskIxcxOZhxAca8AIpGdBpqQsI386SloRWcxXtOXC8yKF8
aHIAdiwsxkOFGHxQSh+x4SeBOKRAo/hBIPWRPoRIl25t0shvUshXZaAM5TcVazGd
OGb5N8E+mU0Ez5FCa1VQUhVfw5U6pia58njDkdJ8PMLR1tf49tOXUdb94PUbKPSW
SLF4ZHEAZmnKQXFAKUmvpOKRN3l8WozzlwKZnZiGzXnCgwRp0ikUrd1Ukr7PhyF1
f8640o6LaHrvaNfGE6BCcWWAL5RvOgEJfWMVkLNvFkUlX8Pmr3eNEn0xsvLigJPQ
vviv9ooPhdNJ6Onc0FEd6x7sZfP/yybO4xjmdNs9iG5+l7yHzTsGAo01tWLFEdr1
6nk+gPDo/kBIdNsxGmwO3XygThfNw+Ja7YAMmxEvW/ouGB9s802G0vKGJg2WLiY2
7f0E7knwkloajemxzRm6hXTgrha3DKfnuX/dUp5XN3dsbw0mBmmQARm7yZYvpivP
owk9X4wZ5sZjN0/AUQEH8jvfD/yz2iScQcdz7N5Zj3q8mN5zvKALTOpyqF7FP7z2
5WRuxCUnTm9ftVWMIA8EfWFbj4/q/Yj9jxCvMR3SEfCTyBsblafNC/z1EnId0KZY
+R9nrNMrKFoNJEscNiSuZ/lsbep2Az4laKipGhPwySHp1FvVBaKHQAWXqwnmUtsv
QFSxEAaa1HR2Cmx+8ICpVMksWOa/gm9xymQUQPhkF6d9YIvbX6sSb4nSj30wmRJ0
17LGroXdBARnE4V3g1e0xBfGvSHbhrP9b2WlLfBNTkI/Yx07k3jphXIb+W4GHLrp
qS8Gavhpp4BPj4BnT258+ru4JwrKP/qeKTKw81VKNBpvz3bnfvrvf9zuHchF5lLo
+SXAwaalIBWDXVRxpmm6zhkSe+GH1GD2nrQHk87OgKPATUUqzS//CzHkUEyPV1vu
TIxphGvzRgnP92uU6z/pBCk92abl3V1SZMgVGjFN3ZKAtrODuk1DbsEcx5TJPWVK
A3vrJYfRBP6gv8A5JXWtOE6CcOzta42W7LpFqT1Nwm71X5P0lZZOXCXVqoet2nHT
/3j6D+1IUVnBQ2XFvOKmYccA6F8w73lLhyhOA1NJkV2H42uVdVAIsUfgXpJYJtvX
aitCf7B9vTySnPp2Svz8U7snF598wjm0Rlh/7tYET9928BDB37heO48F0URuQhqr
izW4COMYPdPhzz8vdCTV5VV7ID0O/tMmQ4Ih9tvC5n32kmX+B8zO1GBBjQsBSeix
PmOU/eNjNA8OOSCgKN7tnmloft8ptUNEykShwfYViJRsuyMaAz1cvuX4HOxDhKdE
fXoQhp1p1M/ai8mH6ptqioXlecz7iVI3HtPxEE+XsCAmlMg2HpqyZPDXwqERazNw
CxLP7kae83ppgiiExjtKz7n4awUjIO9ANMzmOBmRYwll5YPiCNnKFxWzYNJxZTvz
M1g2yyjgqC8ZprW/nEzLDIjXsMyekAMsR9cvQTmpHNJbmC6huLp1xEHXZoklFlOG
C+2S5YWBYSBbL8IctnCNphPNTrMrFKCECsvhOog5tOZiRePX8Wnuz5ho9YJqtcPT
fcOuBezGbcXmc8PkEauuHoWZpo4X35MI4FNLSTarA8QKTi3fWtoQvbVRQL+V1EEN
xFCrn6pnMxHFvQKaGB6TLiWQXKppMj+RGIV8DAKVtKCNvNLq9zPW5tzjRYCnNjg5
hqcwnk5pF9mREGgS3hI2GQyv/zxvpZ4uy5hxv7yQOt9yMvQUL2IAyvoZcwpnjn34
WJsuGBC4u4+JImB59lGDBKHndKiC3S/xigswdqv13ZNTFpvPQ+nLrSV+oLtZ2DPQ
XQOHPKa8EENw9zNVhg1zSTl19Ec92SsEsNzJuyj90F74N/bSJFKaiA3SWAJr+Ui2
BRzyDrPWuJ8jY0Yn8p1C1bbvb7phX62xoC7f9UlVuKisLI6gt9H3LdoCpjYU78en
vQGndNp2yIwgNohdCTvn283JGOVVz/2pHaSGt0U0T4CXqn9ejl674fA6tO8fOOIv
yrd/jC9Bdp5eT+1rjr4UWr/gHd1ySNpxESJfQ08IVlHnpsaTJMwOjYpyQwM9pIco
/Kr6iYxbfLx6Uu+Q4uOsW4ilNLE+uSjX+2ZREV8/TZKGZg+KRaBOm5NC4JwzyH2/
THD2S0rNuW+eANVfDEK82osevUVeTrQyO8bavMeK1uNO3UH6f779lWsdRvwsF07y
eaPsbCpnvSxvaQq4iS2xMJ5/olkvWo/wr00qdV6CIdCPje03oKUGSmQQaWP8Ktpi
vlgiR84Eu2Z2aKis0Ws/8diHl3IOLx9LjxG9cKo37g7wzaMNkviCbZpyuQT98Wqh
NF3JNt/p7HIOK6eGUeCTv/W3A/Y2aashqb46AxY0Zmdd4oLX7dJu8SFwhNvsSmKT
ktli5g9/j9NVV2q67GrBDsb1s5dcD3L5/Kky6sV+W1FeKq0bfkHwWegwJ4iSC3MB
jL9Si+WOtX0bhZk6yNCdOzHie4OMbUh/ek5zRTZPmY6p4FDe9D38fs7BJDvfq6AC
/3Cxa8ScofCPnSlggtUn8iS2RZqQFJrzLZdY2PboZ4drNnipFsklNcNYmqKJ3Gi8
PtuDkfiINNgg8z5sr9QfM2/WErqs9Qg54WTQtVFr0zujjfUliO7Qu+OP7b9dInVk
jMp+lH+/uicfYJP80j0KyIkBr4aaMZlQljIVInopt5j9w0TTAp4lEwOE/envlKiX
ZTFoWLmGObJfRzkKFR/kxdeJ7JhUwyxQ1daOP+/7qSCdyyLmbuSJ2QcYMkfVW6nO
0suFPH5kO0Ph/QLEJ5kys6DRfUfjS4S9CSKw4EsE+kuF9sILxevyp8CpJ9b9xHsm
nIuXCSyXMZyugyqIoU1JhWIpSoccs8e3vLqCdYiG0unTaPR45xSJirjLrog57fdP
e0z0BpqKOGI3V/kUqQ5bIxxo0xSfyXrWXH/iP9OtGZBZQKhMptycz5uCsqhorbiV
P40RUicy5oM63+dXaZI5kIeWoPOaeb+/ZVnd5cwOU7xMY7dRs0YCiavX54Psfwma
MZ/oOhRiaqAr1+RcEdTyj6MuSaEyXTpS3cjmpipC64dn0Jl4lWtYaHVC4oQYdLpd
NNbFXnKyXgcIriwmFwi9RNfdJLaRusck/QX/gWFcfzXbXaaR88Mo+oY4RVI00o9O
ytFeFb6aSxmkx/gDsWzxY1+iGH6kuqYoN4oO1Ba+b+irdbCEXnox0Ju0eHTZqmw6
Yv/sDInj9vu6YYDylYcpJy+YPYWAdvPrKXlUCfklcEHIYAuF+TANSP0iOhKGVatI
2WCX9/149q+jGDFmPFahjbgIzGY68fqO7eLk18/7eJDl6g7TxJQloGUI4HyAuqJ4
W5OyRo4xE8uut3763mFaD5B6hSB+FzqWK1d+owGPKV3uPvKPT9KyVbI9AOK1ks6W
mZ2/noEe0meEyzu819ZwS3uFUx6cE5Gr57VKEuGdsXdndNmtKDrR/TYcHGEk177E
jWTvTTMoeByC229UtRecThmCYXH7kXaPqqlDypcJ371HICWWbZlfhDYh0Wt+RwDx
jFsZBIMtX6w/Pdn3tNooYPAjiWcLBaUxEVp+4si7iuSpWZWg8QlaLweei1RXmquh
OEHp9lkr4jqpZ5zrQem6eRxLyGy7OosHk4EDGcdLzHI2id0e7xpENXbPIRwD2PJJ
Wrbq4mlYo75OBVW6ZJCug7SyDuK0Fl6dh5XyiX1QNwPFhLA8V3uUvVemK+HR1d1X
SgbTvIu8YB0p6g/jQAQf4mUohtIewgfdsVNG2o2Fyae0s0DxrDEgSkJU+w2p95iw
XU8SONKZM6Dk1a0PH9bAymf0OhCxkSeWIt/ichMGFz4+bJqx+yXO/7AWZD3sdojD
3dY0QrUrRkxfqAYioYOmjJ2fHEYK2ueq7BkNFD6mZQhnksNqdmUefz65T+I8iDh1
Qo9GF6GV/Z0BIQuuRuEdZvO0WF+kcO3z7OpRkvnHzduY10uHECpX3tVH+LzGy144
b87+AhUG1vs4i5M9m9foP6QFjjPuawL9gp0Mp2zPFl3bvGnXB2lc6V3Itkut2Qog
INPVnVk7ynHdA/bziATNN4yfPCBcCE6oDpnnEFryWFfZ/sXDUu2pG+ROxNu5qAZE
wH4reVUIjQfUUbYZHlzVEaJkK+KDHPK1UzrUuOeMSr20lJqufiwoyXylZA/64wFT
IhgUILkAv/341ioJQbY1Wo445Qkth4xouqlCWZC1DGnXNWdxt/bprD5FTTdtdX2b
j0RfjzK6+se+P7/KncZNm2waaQV19PqTDWs9IgiGVzPvtY29LtxB3GEvAlx9yFSV
5jR3+pbyxrEzvuK3X7BQQ6i8brRVFrT2UpVOuKTqmOjKPgn5qBYxZRn1q5h9wC7a
aR8GfJTcyf/4EVaWxoTbyzbxYfQ7+tghfLVj+dP2DsltGEVR1JxJT+KEKCbp93Gl
GWZlNcC3u0U1GKBqGZ35mlnSAguAeeyju+qVOgrFfZpdXw9LY5lIkEk14PBGYlHC
R/MCtamFYFGWlTUrPgdrhWQwomUfRagW+/fAj2yS1wSV59gVu5yEbXyP+zPxXb+M
4b/oCCisX/cp6aZl5U+qiB50g1KmLzoDYEMWmFV5BWXSoW9HGmJosYZtyBtvjPyF
faK6KFuJggXN7Ug8poObNnkbxsg7+EA39MW1X36qNQONbyZUOACc+e4TYu7qUsOR
QU0VaJ6WSuv6WBtCSp9lwExBCW5jukSVjCT7BisoENOsovJy5iy9Ro0cvffF8h2H
+uUeeXaliGwq2TCJpXLqEH1aFWS6D1hlL+mZ834RUNNr7mI3E0P0RVznaYlv8FRO
W9J4XoBSL+Z3cDPCwIFTYxMxa7fTXbV0I6A8ZmFYWBl57xuDfri/ZqJsvK4Y9k4f
1ksG6uBazkJuQnSZbRbSPyQJtuCC76qNKpESXQwKydFWQrAMDVN6n4+hBpf9N87O
Ikm272x61b5ZE2E4H2BF13wEmO+tPJXDh/WgJC4Q+ZpZM/atGalb5Fx73YJioKqQ
rcnM+84LaD0+zA6FFcDgv7KJ55QYcm/zwq/oo1KTmCtVSCeyuHjjQTzcXLNRWU9E
UwVPw6+eze9GSBXgsgaKPw+34ZQyFJhyyEpHbHQdqM8kGNa7lMX7aT0Jw3EdG/GO
hQYjBHckaJhpDiuAo3qjoi+o7TciTxLjcEVTuX9HEfHeIus3AVDYVUytSHmkwz9v
X7uNZ+mXk3CPgCXBX0WPupvC/dSaB0ix6wJ/4IgBcKLeupTHWzqenEf2iawu7NMk
u219Hix9dc0q5nDZNlzCudimOZtpWb7xpGozI9Df9t+ahVz17XSsr0azYofwwf+G
UBuPJ1eFQLAq6x7O64VlO+EHKUgMAlJ88O41niYZ4OddTcgNptwr5HY0fuMnxVop
LU4eWPGIxCMUZEq63PYQmhmGq1NI9dn47eOt9RMIyBUbJHkv7uUbMy/3Gm7TBwjB
YbnECDjAp16Ga40TJ1q/DzVeDS7RT3b1IrbvJ8+PU6hCDvE2Syz39yP+ivyCjMcw
cVkuON1xeu/yBzIyxxsYeTAwdchiNiv715jcMIXCQlbb/Wy8PHnFJ9faxVGC9Gis
3uGUYLCDm0Vur73MP85uo4SAARQ1HIvU6wohUy/RJ7F4DmhO+pVGa+iBX+d1ylUw
sGeRKkXnRcK0NCy5toVGYIzp6QCi5/gcdkrgqMP9vgitfDe7HwXImpzZpUOa8PAi
bhF+lteq/gsYPPzsRTvS2XHg+GM3e1osIdlXRMQqCshJCwcCcctzSL+zf/ZrzCIr
s0cKTbCLMpyGxxG+SqjdJH2YZdN2K3iu9S+EGXUf4IaiB3jACjqA3olo3c5M1DbW
oCer9z+5vhAyNqFOwgWZdQaWoL0n7X0P0SuYBGZp1yDuaL8cFEl9354oJx9HkgMX
qc3VT0pxbvog2+C/mrjMmFG68Ozk6jpwuep6Hraoln2ahxKD+uDSEleK9hCr1yDh
wVqoaR+yndkwfrd5eeIM0lgS/SAPbkQIizMWK1zc2f61nBdXR8HM8z5ZQUdgWdkA
8mq3KM3VOnIKp2J+xlAg7i0B9iFeGRYQqSxBJa90s693IFNcIRBoR8kMzp2xrFLZ
5+C0CFacc0a2HvXTw7h4gWx7A/BBkMBtAd5bC6Yqp16j99RkXUAhggNILRMt2F8g
ujjiunuKE75+Ry901geTQOzns/y+P3dDime0RpP2vPvJm3JkyCyLuBzC+yIlpQG+
804gB7LWXfX3EP/YJf0wu31ghuxkV1oOzk8w/zDAvT7ydmnTEqjw0n8MVSzzAajE
0Ck8Qo6whe2IUa0tbfSlFhx7RHTb9ulJnAU1SvK/fSOaMORMELZsPwiySblkiEMR
dpnSjAr2yZAFwmF93P3so+UYS8gDLv3IZbO2plYyLBUKv7iJUagbJDVN7m0BaCph
cf+VoDvrNPTHiRuO2g5BDIbVB3BG+w2p15jSaJ3KnuQ4OxS+zC9c68d/lAqpmUTc
JkfIaNubPoOzGWRavS0JUhoKYdG3kRT2qctQZF0PFG55Ly3xEHmVrxTlvgklUjHp
cUWaciQbZbyUjz1lRdlsDuzAK/cL/G/M23S54VUdQUHlbAJtO2yaJPcSL6HcQpdi
UMGxdgdHjnULoLnrzPG1ex5jpH7E7zJ3KetIpiL5Wpq5jn8awxf0doZzSo1vNw8H
ZuiAYnOyuB6u1IMb5DCJRGTu/qU1SKWzSw/YmDU6S85hB2x3sf4Pf+Tm1QFH6xY8
iYrTyr/qvjATDXjOTZeq/H4mXmpZsJ91SGS9JGsOB/T9E0Kk+HiB+tJ9KrWDhHGX
EFGE6l45FRTl8/U8zY1YBoaIFdClsrPqKW8I9zzzW8qU/x75dbIK2yWwNSjYAl2p
5MUqOBJwEBGer8yTq8QEfMaJrfIfLZKOqMRO/ZA3kzsXJL74srmn0YM10kMn+zi1
ElQsbKy7CPZunrzlqgDgya3Oba3gVzWYF8N02cQ5r+PLQsFF/ddJbjA0UfT3lZy6
z8OAgJ7jMuCUoRqYqX5Qp30yTac4R08PWNQiZ3F8z8aIthsfZWP+JyGPMMrVvmn8
D8pu+SLc8AfCResAEygtplXbW8+07oqrlTX+CmBKOVFnv5kx8v/btEgWtWDqu86S
CfWFQNtznK6EIcMuAJFDbH0GpzWYieCA9C05zmswU32+XNhFmJ0UlP3hmzHKLMoP
LyL7TVN8PEr+EmlJ0620CzwrZjixIQTxE7qpvqfQPDFlNXx8WscRlhKofkre8TzI
dQNSwQKPeIxVxx+eeNxVhSTvb189LXZBFACDOvpEWS+L++HroAHFIn85YtywHjo6
82G2iRZ3cTN/yShc2LAf0Ji/KJ0MQO6o8ShzfyekgiRTBp5pX6s0P/5Tp9A0Y4lh
plpOe3jIH2irq5PFdcv7uzmSyEyNM17zDcEQsECEw8aymxAdmtHth6U2VXgiQzQY
HZ77wBEoQAU2J81OaX386PIKymUn05JRi/gTVdjUEm78wPyqEjSPh8sFDA9UnuQN
fW4Unda+7MIIqBto0As/bshf64JBMywqMKU7MZuBFXtIIR7tL5yx75Ki4F7v7C1H
oLWpgDpH3qhezQA+yPPba2P07TZeGO4Wkv68mBwJcW/ImusS/5N6++6CcpJ0QpIY
jblZHKKz3W8GtE40Ypoib0tpR0GGV+XsvVXni3KgwSxeevTJDKbmLSYtZigC+P5M
xBNnkA0WuZD0bWfHWoz5OcbraDToaPuC3jnnHUMUkGnzGqI6cGUV5t2QP1n7UyXd
+B0EcaLLPQ3nwuqbj6JKo0h5svxA/N9tuN/DoC5efVfXNs6OmisZH8x6o69pIJv7
vZceBpILLgwbTKpCOiTz3RsJ38PIpcSMigp+NIK/S5ZFL3LD8Bp4/SC03KKab+Se
vQoh0D/eyLlrdmL1FtFa2+UZfnCueyA7U/YNyk4iR013ijYKgZzx/Z2b6ljG77ps
BaW06jvtv2wsvzyn0tSCeed0U9uQ2lJxSOkirepKHwcaUM8OXvKd2p3fV1G4OrAM
jShiyNSEQiwCCms9Wkk/vToBHztbxLHPM5ql1rlUtvgEoM6X/6sTeWirMSYe+prl
F0pGIJCYSCbnAmlWGH+XWnD4OEw+RKm4jXg4X7OpSurbkhmjS+ZwUIJlQef+8TqY
HoGXNidd2w2WjzveNpajIMuf3k8iJwJUFGSigFqaCEx8g/Ikfg6V16lVwDY0vAT7
kFYHN110bjr+o+1F4wjrfMWzI7CV+COad5K0QDsUB9kl0/hh9hmEcw4tkmtGGgZs
PO98kzBWzCu/WtxzNrqfHXO8tCeE6OmGGGpip+YpnAlul9/nhXFnqjtTQrJ8JCch
+NBbN5sbW1uyQasK5x2Y9RpBbSSRRRmJ8HbNVao3Pyn6oNmfTEVqQf03eFj0Be4O
dYXJUBTiuwRpdIG+yqOab6QhU7uxb5Yj/KnkIVWmBAh2s1ID5V+jUfdmpF1m0nV0
gj+ST+gHAL37euEYcvhfY9V/MBilMSBT5QEkfY7Fe9mMTpqbE+eRR2g8KMTuxzNY
hQxBJNa8EwgdTZOjhCBL1qdvH3Du+GPp1Npiw5REDn3a/OWfj/jyUZmbYt7fvLpW
GoyWljXzIqzXK92C5OMKDUypDkGjFFXWdKS0nBNKNZ4PtVnEeUSC2iMxY+waI8MP
qUz8EqIPMaWbn4JuSFUVUFNYRCe8U59qMiJI2DEbpGieia06/aYNuIeXSEQSRcpi
PR1PYEiv6oIJUkGM0PRsMwgdPxu1ul8+TE+p57+lWijcEQPQYnxpNfayS7s0Y5K3
XzO8srgzdAf6/2cEQ60KxZkfljcglpH0MJs9sCVvShRa4KWYfHXqUYLmh3fpsAOh
40RLoLL0MDc4SFqYupzxsjsWgB88/2HKNiyeylcYUr1iuC2KdttZ0NtmXWKTUcSP
3tU85knCaxzpvAMe//qYDgmMQBPwVttPQz7QdoMOTWQPYx7S4j4j1j9MdoWP1ymT
9IP+0tUEzEjFvcFRvTi625t0KXG+M2NcHIu/cfkMvAoQ6Z/SZPXXW45JETdFKE6d
GodNBgfPX9dDuiQLxDRj1Xb66hujJHrn7I1RCGN1Mzc4CKhzXFRj/QUXLU+25GpV
WWp5qs0mP2PUPpfGyUqChpmUYhkxRDColrAdRzBnxT9pQJOqagj/X2EIAhqqG/RL
gZGX23InXue0CNV5newGuoLKvQYHajLc7BXTBeDJUbP4K1zre3KVoUVTB4AJWeoS
IEGBEDrnUro73dvVkGYI1WHEh7dgeNOP5BSEk+YQCbDoKDdrM33tPUhIeNCQYPpl
xtN8DHOsZMXJ/DojGTlXkJy398qw5I7XDxsZs8xO/58cQH1yH2jxnWLT2nQx3UTB
Z/7miJ5lukQ3baz5/CHlc0GGAnc+MQrtnH6Xe6E1FlEFZkdLvXCO/L8EvRQHUNNv
2ZiS9VjDdPeJEePiMWvRysp6oC5ghI+P6wLox80ITexdIzZ+RsW/q6b3e8yXe7vI
8HjUeL6+ioLoHt9rUXQ28dibSLPoZKkV3LkucpVKbgBRnaCQezTO5dBk3G4OYwwE
vXpFmrpeb1MNQ9oLp9hDIY2W+ZZjU4RNcHOfE+tf0j5xUF35b+HiCAXGFtRcgpoT
HIsLeyfIngJTt3PLii+vDdhO6r0zg2L0Ox4ORNINNHxumFvpUtAyiLC+dk8PE1vh
3N5jco+WRSDB1spar6MK0ehd7kFPHmPlKRyhYFZzESxQCSYtmQBXlY5x03UbXrIe
4JR8gCyWO3LBN6K/FjPN3qRsxo+tz7rUir3BUK9K8RvG27U0Nk17L0NNgVsRe31J
y2WEOJYd2K23XO8mTIv8qrUqI8vnsYvJzE6KMLebxvZJqng5gdAD7xcURsQMHOG8
80oEDvOOdV+JYQ0n+aq1fK+jbfGAO1PjQva8qQVa5i4I1WYKAGgtexHZTBPsOreC
PpacvdZOvX0qVjrcjci6AAOQWzmTjaHaHiIBPLXp0sjyghRghynjZ9cdhjMGO0tm
IePr/wAXEAxH507hI/2eD0qx8/W4iKGv9UsuaYsW0jb3+P8pv1JdSpRAizUHJ31M
B21v4PdJF8um+yeAxCoyF/66Nv2VtE8QDsi/AG6jLmXd+4yDdnJoLgRnbue095OB
50WIxgnSMgnC7XaQDqVXAs8swFiKdiohbMWNIeBWMd4rovGtaV/tZ5zurpZv9NRr
F6k+tAsnZb1P19jwNmPCLqtgGVFMK+ns1i2rcCqnTR6mEKsbZyBx4wtwKMRJWX9m
cZBD7xxrgnOnA2+8a5pjGHO8pQ272xsV/A7HyEy3Pl9lPbCKqKEAOPNeMZ4jEcb+
HISanLz0cnwk+LOMmnBk3CE4II+H5IjjxhAwpsOblIGIWPqBUbr9B4v9mkc5TgHJ
BGSBePYyse/ZzssyLikqsLFWtdsB7maeIOXE57/AmSgiUExXAkdvwLXe0w3odZw4
HPck4f8hheeiAWHnyyzUsvb2LfvZPgnK04/GLHAZA61j4SpKWIkEDq+cNR1JPNHb
9h+lSODDtXr86RVi3I0oizgkq0+DgjVsXhP5Vrqcn3HyXfmLEw/H6HDWrW3Rvbyw
1IQfkZHBX5NfYnEPSC/pVD7qosRz8Nh+4FupmkMUP8Ddjd2kcM0Ys7g+QuecbhCF
5n6VImkStyO+qUxfdfdEufiVMpAPxu0tFj2c6fUcz1DsWpROaVw+zbU3MtEaQy7X
dZ46tUJNLSuOwUDBiA96s7qa8triOPPiNcMDJCPE7tSEqaFo6uQgdk7eVCbbkkaM
0Kv/p62OkCpIxG6lMM5a6t5dlyeiSTXFr5a+e4RRYiO/1KWf+FdRA1ERa+hSN/Ju
dXeLib5rt4Id5nDUejSCKdUqS8rI5CfNEdhq7A0+fR8oswF7O0e+nseVT9r2IZ4D
r+7iz7GH7w/exGniCtVTeQ3UXUpv9AcojumYcE/hjEuAverKuVxpPVq68u3yPvML
9iotaAf7s2msWnEPpVKadK4GO+QleY6xqgit0WBxrISz5+9PnUSactqWjRJ6dJue
rS3hKykyEPje6ouISSBOc9HCjtwkv5vNJdp3rIYZbCzje9CF5GvuUqK/V64vw3U5
EGeGqcPh+j8Uo5XXhBtw9ZggcJT3u9mw3bvmgy8AIIMUADOGpEbB7lljehTpKaAa
192TImu2cbkqiPQCNZ3q2aBmvez8nK4gTLmmN6cMlBi0KZrhN0sDCPiP1wUFpMXi
ofZ75IEQXlRFQlIU5QV/C6SECX2TEAR9/smkyVyMCiLSS+67UrSfBjWPLfNVff1R
CuEE2WHu5B6dZPZIgItagFbfWxFN6n2dNkWSgTtWry+cqttcpBHZh9ky6pf8AQwS
p4REyfDNCq2jiBeEUArID4hXhptu8dH6JBMI2GLzaXHOUDoWBT2JweyGmYnvj5Yo
fHQ5FTsPn88mux/EAcphLEL8rGOHz7gYRx3QkfsMU2iZ+WtFEvrgqXiuKAlghSJh
DIVi9J9Z9+L06ZLCxp7ssWeFIA0CEOxvm31l67oDSYtHx2d1P391SxHQytmah7Pz
V0yKuw5KfzeS+x9k8mlRXJIi6Mwt4wgt9z7Nq0t/RCQkKgXvGoF4EMCzYWoTMfFY
tGvmaf+0XHiZC6RTKxWnWd6H3QoKBJvPpoTP+mhCy9dbiJs6MKcytaEzKDoF0nyO
chyl6ZHcemGcJEtSVIBghiyyTk/awzizNC2+PAoO5CBkNaLmMlz4HcVeqUaVy9Ul
jW03xCy8D3mkaU/u0zup+zapjqDn8NuQ8hc3D/yXjYn4uEX1UNFx4lKdY9r8IT1v
GUKgnLtLxbLD4+KG7PKZkpziWmSJZn36R7/9uWwSo1nMqLwvldSwZQI1o2HxmbZp
mYylgow3tJ/sir9K1IeIQZuNZBP8dOGBU/gDeAOHVgG7Fa1EEvju37n16lYwQQsE
R3qnT2nRVYHca9npyoQyOClwALbCarQ3tSYIiJ+dJ3cgxQsMkRjmToh/u8+Qz7Vb
WAN4h6Q7OKP1CzaXsWPEanORn33AaGU0OExlm/oLIkh5F1TQoRlfXTUUA3s9o5L8
0KbySFYCVLIhTf+H1Otwo15hnGCVK21i9xtkOTrAYU9E972x9k1ye9/hdq+nGWLO
4UHARFWINmCc+uvTbM9lqCHplpJVcTmcrvnkfyxPVVJnfiEHMAr6FbmSxOoIB26y
f3zoGkDJdF280ZadS0yVJzFg1y2Wh5kSq0bIAyDPz2rocYlqzPYVxBfbTKjlhZUA
xRT7r16Qdt8ZOsFg15m7w3D7w5SQw6Qrpf4YK64TcCiH6KtJf5Wkg2lltJW328cR
gyaWP5SQvwnaUnUbEitY09N45Axlshyj3mOMT18NakZtvbgSJYby1qipfTwq8hDl
MvR863vw7YI1Biuc2LTGGxWASMh8Gk98HBgV9mxVG6tQhQwfSWP+o7YDUjndmnLs
lfJwYKv8DAMbB8owJUKo0294gdf4xodvCs2FD6L/Rl1GhMsxaXiT94REPW7Hu0Ip
7RablJGH4y24FKjaVntT+GMi+cH82PqpinAWsggky7vPA8VOQKBzLIQcwOCbsDcX
UqlyZF7jIMqlA7nRxI6lyTDYO3BJBejUaEnr6stHVeBuiLr1/XA3IxN6Gjj01P5F
7/leH6n0PKR9ZedeuE7g2Kge214ySl4mDkBzwIOfeq0BbiPhHUf89lgv1u4HwrxZ
IDsQi+sxKs1TOny+2W7q2Zy+hX5Lb4JiLkOWkIndQlga9hb5JygXZ4TZQsZV0nYz
1DK/FGJ59TuKJuDHwGNKRB0tep9dDWeqUOZ8POJhCb/UH0Ji2rhGrYQMb+PXinbM
F5jHyObSS9CSgTVzoUhQ9sQJWvTzHMKir83hBx7iqdfy9BL3Gg+VjpVkC4HjCCZZ
6f2uC8c7/OgUciiUTgoJZznBdnmeVLx/Om2v43Apg+ObMCHSgnc9V9RgQn8iKLJH
jhj9NyS3axrzx+vMLlwxGwq5QfSqxlmp3myUODh6ipBVLWgP8W9JQ0erouGrWKeh
UdEJ+kWdovA7/0pHr1NP/PrXtO7nSbpfYplA7RRkddhh3VJpDaLzjurcT6/GE/3A
nsJnrlvvLNvsvHEaBOlD0Y0WfLCTKffk07JsbOqIBNW+30deLnnRCmHwFnkOT9Cy
IR3/L/J9NnWVYIGqrzXOyBw1ld+lYRdlnozW8dkaECFuQi//xi9r0b+ArOakDnb2
Q+hHkVTZnzgGDhc3x3MKmFi+C89x6MVlCj3o1kkcEKteclLKjpHSKTpYSSCr93gt
P4dhaLaen4Pg0kevJgiPOWIJTLJkB+Fxxtu2Uiag2+hcIH1LJFLleBz+buoIl0uf
28ZGHjXzVlXpTV9b3F5zonvxnAMHo1OhHJq5qcqt3Fc069sH9T3Dqt/Ll2C4e4Gz
rwTESgP6NiLUuddOltTUTPwk3A/36RvinJeN/iaRwZCXLk3lpFtYYyy3cEbJ72V2
kr2IQ9M26FhpkZJYz/5zWatGfn1KzNyJkFSGHSdcqNfjYv4SCQ9ptvTnNR0O/GmT
mPmyKaydFdtgh35I4a2/7Yn80llLPFYBL+J6m3w29rK4hXlPtR8sFa5dnl0ah3Ic
OpR633aeBcd4ISj49rB2TLxFfNdNUiN+L7bazM8TnoF7CiEDOf8Ta9YWBbR6xhjz
Eh8tMsciDQDvXktxrwmnjXCkH0WxqZZ4NEqw+MO4CUY2yqKjdTdL8YRbANMBK+20
oz8k9rovtdAmkt8bSKmPiIuS5YujBYDxRCFx9VG6XWWTh9ILZ0qts12XNhgyUkZ1
puG2KGUpN5p/mcWBdFC1CKfOzytnJV9IBLgLcJ2/AC5U3eVUUBUWC/ytNW5G5Yna
nuzKxcgDe7xUAYx2pHXMoMkiiGGKzI4YGZxaQP2OVnMG0+bFH1p2lxXU+9sUYnHj
CRr9UuR70o9gK3OFd5elAKRAwDxBkzwNMCxsGGkymR2q8DGtBtRVDGSGKlw9b0P5
MK+hCFc/BOtghLLwCuLDxsRK6/nXi6LICyamBvPbULxieOhRYE3IVyB7GLbMVcF8
Bw27ZJKCixgKI1LY+dk/d7X7uKYCzWZgcmKV4lWs9VI/t0ROk9gb30S937xetPUT
Y1Gb0ECo97xcKHpZjxyugDDaFRVeibzKLblWyksSQoUAjQy7OPIuciczeRLcNNDp
`pragma protect end_protected
