// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:41 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
OKxP5gNEiGlNTQt/MDwzFM4K+L5R52nolv5iZvl+WdLrYY9jWXyr9cpB4crhfsBZ
298eBRZXt6bx4OmLIlxzCdkfX//giYyX9tJHvMqSGOzCGZxmr7BSOA4UU+eEDVN6
ZAqmZQhC1l2vhmhRAAkLE4Qk3MC0vrLyfH3mJZXuCqE=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 1664)
C+Gk7Ndp1xd66XbkqLwRbCRHV1Q870QyOUiQbKwqZr2r58CUB3vwP5fQ8ofADxFA
52o3ivJT05GcB9zUa3t805dFs4/V07xVw8QE0njTyKnh/N/DrCEVnKhfPvbfWUr5
KOExhZYku6aB9fjZwx+gpl6UTokzheJ3ON7GxQaIEo/LPg5UGs2HpUMT9DZ+FIEi
tePbMDWG+t0Kjlh3oxEVcyT3toaFODsjtSXOhCQLboWgBecOO7ScdYWt4Vn+xXqf
qvgQGxaIUtvL+85HgQ66lynNSyfoulxPYhl5ftOxwPSIibutpSFX7NmsZUNO9iox
Jx/LHy4K6sjhp56D2MUJ75y/nj9XGVgHaz0zhsl5JOevJzH/yG1MfcW/UxKHHs1R
AmzOGCuJHuXxRHqeSRacaL5tkAyDbuhdOjdH8pthFyQAFmdaIB6UcnbzAzzOrVod
VBOmQI3qlS1PcdARFTmCMCCpNwHLb2UnF7DpwULp2yGoresJQdUZSl910i3OPE/n
hCrimPOtLK8Hb6okz7gl3KntzhnNnEBfpFrBCZgxHLw8q8NF+Ki9tLQQTg7ZXRT8
XhSNVJOHkcKdiDi+cno/COP8zaslowGd/vGjuBs3EVLibjzo8XuwSRLbs60bbrkv
ZzRVKTN5iDXnOs7snPhJf5Iv490bFoNK0tTrGpiau73ZyojlmjZ/2wIO7nEDSCor
fphu1xIgWM8AsjgZHaKZ/rEm6s9M23EslNB3SeyuhlQvxrA1Zgm3iDGP3+wOot8M
WwH68fo3Q1nEDtktnykgVSvlgKI729FqFeiCmwc79MTrruPAkVTQ2pvldM4reRdj
N52HSmjtEcx/h2ikKY+PmnAZ0oe+TtzAy02MTh387feIg2h4VCuOQY9XLHsAMk9p
O5Zrx6ewjCuCvQHwiY/aBJACbK9QOza24KFB96Z/bodw3rMZHVuhUp/oSUeNviXr
B3s4I2GuZbVpWM0FA+G2NbbZtTKSETozGUR7+wtZ3wKCLgkYfoOdbhuT1wKdy7a6
qKZGeGw7BWjfJzFsltT8wgINIvKLkQuOgxkrRezaAc2UIqQfFMiIQ4qM+9aDNJ/3
6rrr6+gcfXm2MbjN4ruStVHLn0kyRZUukp2xP9pOHGJ2Tx7Z231/T+0F2NY1VKPf
pYmRkzXctKMXlhzq9N781m/QJAG8tUDXNlwl0t+WAjzLCUIQdhrEKW8qtZm6g0VC
wxeqiERSsSRQ8TV8eCtIlHxvSf/wFy6dqEkZE01+GjtD4yuRKDRMWMMy9BWAWcE1
lyaeLoRyfbo1cu1cLNBms0KEkHszpyxD1iH35XYqS9E69xFtzgC/YQK0ZGJxOe7g
D6OVQNZ0+zetKmQkQE0p8YbAfKM1SCIgSr8aPzh2vLDjmu/23JP7O7SqZ/A0yyJZ
UBgN+quPzqug17u59RsP8jUmg2eyD8CR7yeom+Xx7Gy8CHQhc52k6F2mZe4h6hy+
EkA+JBv2MyrXSzUZLzn/jlwCIJlezNMTgeBYPSN/CVceHEOjXu0yKhTLjyEYPF2N
HwEZ5xyQfmffwcpUi5fbdf5Vve/+TKeCmWfvHAw6lRR9qhPFuznac1a0Ev0RiT6g
y54WrJW6RSIRKlERTOWONTo8x6PKNIxG2sP6X09VPrnmGT6OPVkumYW3z9g9zRoC
moMDwORbbTKykylH2LVE4ojsSjuhHv5X6T46b+btGbTytBnovZ2LDqGbxT7o07m0
GLLqF6Z5M2Dfd01ojDraG2XP2UpF7wbUknulF8MjBDSJaLtxSPn0fhic60EVJ0kR
f/eOvU0XeXHLHkgGSlzAOEkNykqHCXc5dmu309JO0rfoh8DsMw0ydwUQS557i07C
eOWcw/HLKGHH0DJhOFm6iyE8UOq91HIdKUKg5YC8hmQx812BDci+YaOP83seaWq8
6dZVFmpKGqiHrDtDhirr9e1ajXy1A8rfo1zpKn4j40s3EihvPUMPJp2XL7O4g/pD
t/y6Fq0BL0tDIf2yI9Z7FJcobSCTrRcXhunVJ34eV479v7ZUZaBiHfXrI+aYTKPQ
+c56CRLd/Eq2OH4I8aGAdMmrM2M72ifqH1RGLhRnXiPkOGCXrWqsjKTC7UCf35Le
XCQjTt24h7ARvymhiOwrx9S9A4kgm6/Xg2J4IvRSkXjuLfJnHQ5BRsgP5Fnn9mtK
TVQBxeveV9H1zQkIOebu/nyZwHRUnNxFbjmQPYIogRM=
`pragma protect end_protected
