// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:57 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
PFnxDydNPn3A1iLE2sFgvqC+GDK7YBkxGGV0gtS2GtnPeVZ67MUQLLz+QDASvFS5
7sx9NGDKGLGXzDzkgGmBNNrJ2VRqOZ6QKV+abl8FSIPfJJTLsTrV3+jOQz2qulhe
ASjlBPhzV51Rjchj+OYV8BAxkF84q4odklyO4BQe3LA=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 6016)
o32hWnxrWLNj374577dCC3OExC2hXU1/Wxw164NkUqYOXvXwJO6U/us5GXZ6K+6v
eexVm56IKAy34IRkxDY5+J/yeEuWxqFDXqIoyq62vXvV0n+SldfzYeuoZd8n9DUM
YJOEVqeZ3oct5KvR0Aaca5r9AedzseKIa8Yl8rP6rjjdh+o9wR1nlvAbMGADkvfw
jA7aOKXZi9Sz61cjG4+zv+uAZ0Nalk8+KXFBKLhPd03lwg7rEFZmC1ZpzonXCqbG
N/zojXQQpUo0hQoWN8SpqKtWTN9s99y4jbWbzmSYYiqFk3AXH6KAY6DDBDZi4FR7
2po4YYZnzFkheVg9aJP34BTW+WkptV6vhcI+vt0l8NZoVBgfoUftJzIg/sOtG41U
CaBAZHefpkEEJT16BPoueIr5CIaYIVJidHFZrSHew0/fBdyQxZtggCYabZMHBlnu
5VR94kYgh9StGC791zmqi0VajlXUemDauYTqA1zaZXCRWkGS5cuoKvJJ+m6zKobb
fDqVJZvowt6qFBikgNCdhiodQeIVfLMdK7N94xeFjMs746C8ZbJNRdyPvEpdUbex
GocTGKOQ5IAtWSUZlj1o6vs5KH1Z6JuYMragZZNIqEGQ0JiUX0z88G66ExoYUM8s
Vd6/awtw50ShuSEDLgszQwpiaB+V/J+vPzMNe5CCu6NmkS8B2wKXYN1XTEOnkfgg
ckON3NEGi53chZ5WVbxhX5oqx1wbMfHumEYLYyxIADraxd8RYHMEIxnebc1Soyeo
0is2J3HmLFw7rdqvIFxqBJ3/OqKEWcjbfeIfaEltp7CbJ5pEFUqUE0COpNJQX94H
aqJwjioDbHz243ZwO96PXsbpiX1ZVO4jVksprF+cDS7/HD/J03kjtG9SdOLYbmq3
THHjixAy09BHa5GUsqS8ivx1WXsZY4R5rT8A/FbtYeuAn44vlhqwQRqBlCrmzAdq
1b/V134LTgCWYlObL7nUgR/xWhX+jwGmAnjGwnTkF6iG5kc7HVeZMuO+om+YQYKY
s8OeQ+u4pVrWzLuACLpNhXM/ykNbiiem8whqmdmdCswdvgQMpGzp0RXmXTgzhqOP
SDjlZRY8+ZHNzSPe8eQyv2Jm7IXa4x+HMFcZTOl7DoQJqePn5pENx7abzk9bY8Gk
0OVh+OHwIUOKIJBRSFt9JPjJPgPL1+rSMuaiL3BcFNedyxUwLUl/Tx/f2/fLb0E9
0BaEcIMFhxEo6eDsW/se9v9YawQYlNsHMtw+ED6vQDN6StyHqFYY98GV8dMYWHoa
xkzALS5tnZG5Gxux1DxNO38PSYxLJIbQ412ZBXoXBZbJQ/FoPuucByXHWozX9hPC
ceUEI5GJKNhUduddb9UxO0TN5ucTo8xB60osGtMteqwyK7OJ31jJtyF8ZJ1beTzZ
blJV5BLRefB2oZxZQMfkP3UObvSRNqpFs7GHCOXel9wiu2VS5TjzTPFX26RmoESV
yOIrablbj3Rc8M1DUwhsOco6UpKQoY6JQDTqcWDz1dr3xPawOCkhx+4BiQkzl4Av
YAKp2TU3EdSWTd4zRRLqkPfloQrGTfXIj9gzgbzK1wc/RElnIt5DNvtVmmRvYvhK
lU4uL9vQ2USR/wdxCgZo/delvn5re6JRKEJFpeVqvDiXiyWcSgamyjbbNeV46J8V
j6Pcpn85nc+G6rFCBX4CKhmLWWDHFwjG0Vj4pOeF4dvuMYfx0JlWffiukCmngbZl
m2xDVdwEgkh1ZjpWeLJUiboO3eBGd35l3x7E6KXlLUOO2d7QxWcwnygqp5M1RhfP
W7rWI8VdkP10aPbJ2cuxQGuCjZwfx+1p+F3CPfwAvCsstyAurphWYjIHZZZlEhsj
VIFy6Jd0Y0XJPFbmoYMNL69dCtKHAQFxQ5y+cyjK71u8QOt33+MRlCMTGooDGAw3
nHSb/4WuPkVeO/nY+gGiLvkAocUktmOo+u+bkCi+TPEVead1mKwgrduhpFaGBV+1
egS/1R6yW3a/ikabb5fpZWc+3nbO66E+7gbxCO2JNQfQHKi4O1yoiNb07BzUcDSU
BPteWhYtfFPR9U5vDywEMXwbPjEhr5GsJ9xJ8qHg63PjvJrpbC/tawoip2rJ6D3w
Rkqth7dHVOnW3bovj4Jj5zqmIVsZcI68pJiYU4VaUzhvWc3NdA6V67HRrvNW3OT7
nrqTT24OHwkmfF1irLEl5YcqxUuk6uihayDtC5QBo8z921NJlHFHw2+rRZPW74zg
o1Rm4Mj+aLj3hpVinKmVeFf148gvtAVOlkMb3GaHR+jSZ9QzZ9UYfbTz6b+8EKB0
+W9GH/E3Wefc9uuet9dixnICZWMJaohPMujp1o7EnN0/d8a0AZVeFlv6ihr8Y2F0
1opW1LaFi9BXFZ4YlFiQgQADN/3Gt7krs1wAtMsyD51vA/FJiXG6UT/YkpcV7f8A
RSSxsOxN6PKt2M4sMv/x/XmFFAk8KsVsL6YezQBelbuPQe/Ojdgsuznrgr5te6WC
xUMmeVcV9zlyJ2CYajRXpEDPVcwWBMHsWsNmB1CvpUNFZZEpDgGJaXhVqBgPEfDr
99n2H67YUAiLvZ1feB9VTbF5h4kPv4ilUdBxCr94IOEVUdO8HmfpOTxJYOLwjg1q
j1SyPcIDksiw58pZQ6EadaPMoGWg/gYNLs6iJzXiVDF3KNWS80gckP/8FTN9Ni4V
cI7pKaseLSzjFghKwHYjCY/LmXOGNSZcAGnb6PBIPndOn3u5RLd3BfNEftfhBdAF
11o5XmeYEmDaVvunuyFUiAaLiPT1L30/6+Yp5ORJLd71MqBgFkJ45g8TzveciCWH
xhqc+FvG7gIiQxvx9n4JgXOD+lniOre6LYSIjSYLzYUB3SR4d6zt3l67UqiOG+cH
3CvuFJ1kr5F3B9I1quGlxoz9wwqDOB8C6v0xNu3OpJ15gIhmVg8zlJ+Xtr5hQyXY
HEYjG0RUJGZ4emxFZ58hRe8HUK6SmrRJ3iK9PNgo8gy426CJ1jWIAyAFGt+SQwCm
jz0bQ6Z3MyUUHxKAH9Y21dCDPz4K4bHM2sXaPfAthttNP4lWk+iJDpf5n89GjOYb
w+XlK8HqKcYjhAbNi2dA33W/10FATbzArAfPpI3eesWZwgMuRG7s4vLcW22VSNsi
fKgZE/wWOZgW+tUjRSh3Pdg6UYzx3ri+dYhzMZga3NJdyEbO5tQZhXMjKkJM4CSV
uuJcdhB3Ej8jGZzqxrUvS0MVh70MN31A+Lw7HgF71ad9LiJem7Wa0jGFTQiXks+P
oKvYzLCsvD6I7UV6cWN56HMyBJ04n60dvqfvCaG2KZ5X9tXP/9CZmKnD22mGJW1A
SPzdUX0ug+jyxCEdfwcXsKcHg9NP7Oz5ZgcWVpgvM1ktgf0jJK0ab44JCkCLIdpF
eNpW+78IG5dqwFfGFgJZ/gwhfKzHJNl7/yJYXYepDkBBgmzEopBQZG+gku5AFZwQ
6SnlZ3qUvRM91WNQ9Brmav2OyIhpfvxcCjEGdMzreDZW0wW7Dul7K+0rz9mwBOYt
DMSHa8GBxfkUkkMmAdEbKs4ZqbtzOgzfZvkVgvjnMioBpAckjjN1ruDVWLmPrC3a
MiQr2jssGcRYsk+7MKlsUWqtBGDDRDxAVyHUbhFze8C2aVqMoX9INoCkLPAvV3i6
qZ0X3uoIgO+Bb3w0FgCJhzVq2qEVJYy2uKLcyz2g418A3Zj0h3owYVE0pjJO/Qm0
9gkhHN2lxoDO5/LlUdbUvo8+PuX1dSbaGJO1EWAUNBSBpCNBnGx7DZ3CR/TjNn/m
jPYKSPxtZInes3SnjVwYvnQ1dQ8JN2Ex02Ywz5Xd/WkNuJ0W+g5DvmMmBa27Mvyb
jpZKYHKZFW07WL5ieAICBNPplYxRCAQWG9NyWumIn6LFNPd1sE8SEkfn1/lzefsE
fT1xB+KDJ+DoRruFVwHusNFa2W1TlRWg9bgTL7Qp0bkKs2leJ7rW5fY4ekrDx9EX
ocubMU9opMWPHE+MuX0Zrqj4YFLuauQuIRuE3gAPh6nYFQToaer8XRtrEMhHSx5p
bFusfWfqL05MwxIRpq38cYF1YgKXLK1cghuytoK80Eh0bYq+reW2emp8FsI23yVW
NsuoRlvjhGikDYN46npVGfTdImU+ZV1K2BdKXFqtBIYakM7LoeMUHwTNNNxa2wlj
EcdSeHbvHsIrDxrVBXdSS+3RI5/0DPgUT8xlB5u/XPijXQdBabDu7XNX3rJYdLsL
dC5AXy8AquhoaHTCIMVX3a4XQMtQmcuLvvz1euiNaiIIYprGiw7FNt0qthjMbQqg
vTPytx7A8errnh15kTxxDRiEUKZd3E7qxfXPm2KM4oFko5h3/Vad6Pl5Tk/jkuA6
rjdm5r3bSyBIHmxfEg+tTV4/Ub0OLOHpay6LmckGecsIC/TjBvbvbYyOVSgkBuiU
RK6EvjG7vdpu4ekihdA/F1vSXeG6L3hSAl65j7su4824tbKDTrDMM0g39LHcdYsU
k74JeV4+KVGgjavGwbJeJTUSCgQ4cJtm8JYTRVaw/XsEt8/LHJqpm3JxMGwiOf5D
w4OMoDw4AJnzOrEWvxcHPi9E/EmNfZztwjsIVo+SOPyHjvlBI/BWpabNOZBzoFHe
hxR+SEwJPE5vwhQDNV1k5rh/uduFjG5FVhd6lFgNmb3LoVRF5V7TBrDOT3AyIbjL
oG+0ZpNT4uqqOFWN5O94tVK57O6UWXNuGs9wctO0QeYYBDDbnIk/iR6iO0FFWzxx
mG0Ox5T1X6fsSyLVvMuHOck9vEB1yvQP/HRrkMz0TAIZm7C6TquE5jTalQWwudFj
+uTG8jTjHdQ+vPLohZoJ2YM3kmBhifbcqsHnPEujV7FZpW04RSrZ8VvZsMr0S5wI
gzEMMXX6yOiuBzx4zKkoYHHOO7yKdUtmv00+01YdyTd9+SRp9QUu0TZNfQZADyRD
mdJiQACtqI7TVbSu5O+pB+60+wVgDYh3Bf1WSIs1gwS4uhMOqa13jnJT6T4s7m3M
DTmal4uFNqfnXLdOZt2m5QMMNOcdqRJF3VdyRMruDoveWnwmV1+Jfnswo4fyMYCV
S2hvJQrZXUERlr7PAZvOhCgQRMZo3BPaRGWjphbpWHy/Eegl9URQPks77isBEu5r
WcmcbbjChaEJuJ58BPnuRhATa/w6VE+tXDwHBpZicCjw+56FKjNaodrBsLdBEYFC
D8jc3+DKVx1bV1I9q9Bu88O8Vm85QGu2kdZhOvtWjija0UDlRDUT5e7+KfiPb3fA
C54EBATOefz388U4usU9B3Nihjh2/Go56vGIB4t3u7vfi5EN5n90vnyeke0g+Ure
ttzORM6sVeNSO29a0ZPUMI5866khqcNjNV5ts811su4LoiS+yxDExJUf5OysL3mP
HybDB8laMJGpn8q0VoQ4PmQVGYKBnscj6J1WnjDJ+vdM1dv01DbU9PFs1Ax8YX9p
H9JoEnHhd9uXpe86HCmHi0AH92ohwkR5nXQlsEqRAF2dDYNeoNoihS4pyt9Vvdd4
AhXaLQrFYBapcaRuS3szda8HVSVFDOBICgy2VQW0YiX+5NGerRV6TdPad/2ZV0Pd
GXJCGk95ehsR+yDpQ+Ve/s5AZmkSI2gw4O4Pu4us/ktGKTbz9LUOPBt6DmCwz8SA
JQv0kRLOCy1zefM9iTKiLmAweWHcz383tlTEAtgW9hjQKPUKxlqMUgVjrjjhVyep
mZxoyIOfJRODBJtLavh37sFeSd6r2NHqk/GEhkre3HfL3G3rF6EeXGHfsOymSr7i
/+1zMaSTWRF5pl3t0hQjctAqOhXGWUjHQ9471ym1mnl0tUzXtp7SdP8A5lyZR4Td
GanUFoA9srhspnmkJGPyOixspwA4Pnyb/GwMg3HR50jH79nY558ftwGNPJecWQOQ
SC0K6A0ZvLpYFmRjEJ1nr1z5I9j2GSP4C2FqNVEXg5EMcQya06JQ6M4B9prrOlC3
bHWdZUHVMVKReLkqOJ7OAtyzesNe8N7sjlmrz8BnW4waQaE/b+s0C083VYENiu0A
BORckMnYodl5UrDstZEB7Lj80Atq9/QpdlR+46CpMU/dwz8YqSPds4il4Jfgt+HS
Z18Wlc0nIvhqDepbBKxQPI2PXrYhiUdAA2oqBQuYDkow5iteq/l8/fmxABWFuIuh
ZoMzLqzQXHMDzSe3K8tVsYrazzn7UHh41cgoUTCvyF3GeloDlE9DzD7iH8FyV92i
uzZRXy9rdhU9gyfg8DiATgw3qEw8HtbPjSkbVisI0LXf7pRuPHg6VhzPrvptPKVc
P1Vj9mjYf8pEkuacsoLQhI1pAiu3K0H4jEJtjemcYwhtnPviS8HcK1QWtxWUmH3G
R/D/mNY/RJ4I7JyKu0XnaTcy84xqJQg32UCJOgvYt3jkK8iAbdpUiB7QdXwSNCTP
HA3DH+vIvTsa9cj9WkHEKcxOR0OuYvKoOallILjFsbnJUvyRHRkmv2XGKY4RnUr7
ybzJt85Q0oje4lF7bCjv3LSnSTguVvR18ehpNfpSBhI910VjyQHoJ0iYsc6DVrs5
zQRrPrG2k56u5wYCciKSNUULAV9Dd4Y8LtaoOWNTEY1c+Vs3hHN8uaJl9M3+dQGD
65EIhOR5rQoqgjgl5Ousp5NFfbc8cZkwkXLC+FnopS9Juqey3qSzeoCF+QMOla7b
U/eaSdqWxxpM56fpkSriwkeLFG6om4Js5dRvCEmOGDkVHkxCQz3FAmRokBrAhsmc
SsQOWcibCEgsTyKs2HO0dtpjxQqXxWfe918vpleJmgUHMTFc8uJqF0kVDbrKWkSl
t+XpS7NNVrGGoR5leUD6xeDiwmsoFUTFcM+rxLFTdGwAggOxiYnwhBSfLDPru21Z
ay0fngmXPAFcHVVRCLNrY15o0PthdEwt/L6U17gC7IYNkrEFM5rAYGr28bs38ZFu
thHFHhHMY7BfkjK8ub732Ea3auro4YetDyu3ixppdQP3UlW1NRPYikD2g0jdUNm1
b1oO4WeWcqnSPqFb5apqSXrklb4ZMKm7IlvDMHckQt/eJiDSTOeVkPqXcVdfTkqI
QRjI/ZzXGVI3ZoVw9/oNbwqSN5iW76cos7e8BNw4R/RM2SAbME4wA1+OIp2rmYsd
91dHINyVqPcUjfXvN+7xRdmg1tw2F9nGAkCR5kLco08uViC3AXcURBNCmIC5QIQY
FSjdZ1NgTBE72GCPL7BgCTpj0n1NW/H+Zd7hCOmqu2oTxdOIYziCVats4h26RTVM
3aRKI/MtECgbzFEvLA+/nLvr5LumfVpqVnLip3FRE1K/bzbKAki2sZNGDdBjaotA
15hizQizyy9qZomkIo472pJO7NF3VWP6clclwv4hMsDhQpbIvB3cB7wWykpxcfY3
IuOAe1Rt0Z9F+cgYIjmHPfZOJM8+Qv3a2DM+hrNdAHhXNYGELETPK4TIYjdnbUOv
xkn94v90OEEvV4GIriF55GlVTUxj926tho2oQvhKJbsMBvuCGsMtA1G0CaA6EWdn
wotZMOJp8vyWLbiEFCsJoSt26Da9ESItknPTPGE0J+5DFwuRCX6NBP1Ayt6mYejh
xbzv6b4HDF2C7cCzCQi+DhhV4k9Z8FBDUCdQJW+/gtx9AckxLsmScOzh4Xy6d++p
Qx8UJeIyGN0xJ4mi/g5fYQkQNS/CNTNkdiOr2e2z8kjD2c29GSzTcv6mectfFLhX
T1zxDpZyvzea3dfEp8fqOWvFzLvA2PBjH6KiaG2dtF8EdhJCKfDj0Yixt+8gwPko
erUleILAozfcxtQi1GQwVZo0JeRoJ/MVBm2YcE/vMDHxqnZXgwVXDbEe3B+krMKa
rCbtWXHDqi8p7wcY3syQEuyj4H4fi1CUs/cQqpShgOsa+3QbnPW+6UuJVIUSu+Ra
Pk9peIw6ZPV0aSYAn4OPOcO6vPuXXlrAWTj9PGN+iCgWAe9dqAOiUdOdo7M0PPjF
ld9M1bsh/8Q780Q+//NCctsv2IwJjRVFgTrsv9kAak0qLGA15ykqLtWruHxE7EVR
c6ZaOtL99qyvRdoiCjqhQA==
`pragma protect end_protected
