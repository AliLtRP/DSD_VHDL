// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
kkwanWbLKWQF73PulnmmKwHdFyts5TgN1Q5/VJ/Nm5LbWPmkUgOR4NTCVAi/rB8n40YPwkAjSH/C
ceS00kGLl2P69e1gZqQCv8B84cVnB8junadZj4ddQb9Xte7b1xveGA0TBPNQ38q1OJvcun9lpkt3
gXJ6dnhl/TIMIjIE4PQ27IBRcuUTcPZhbKHwhplaWTfoKn5XWkcxPfSbceZ3qzCIjDiUpSGzZ/jp
EFtql1NYE+McGdCfsNYnzIfuwapubLvI/z7u7jtXJobgrE/cZmNDaGW/6GCeVeUX4XFFcAeYbhIb
KMf5eCtN956W9avRQ5bVuN9a7Ec2JNUxHT487w==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
ujL/sL1LLcHTpcvVSX/Ys2fUqGax5jtz5nWAVOEAvYpBCvel5v41ijrSxAsKOu1zVB9QdRQDnK99
JaV3AL4AxOwDtdWiAqljyeo+/rMddav01mYtvL+QrcB48d7hn0U17mICHXX42raGA+eG0dW9MErT
O9FKoDksWC0ov7hjlMZ6c+5IwJnnCZQl5RStCGcESD7K46MyNeFiInZYgMUOCRKi8UUA7feEFj5d
NILfNsZtaPT7BFq2IpK0Z9+6NxJTWEMl/NaAGeOhZCfIl/RSK3EzJ3hddZsZJEmYWDgK2XASi7Ha
tQu2oqizeOwtqHE4knOXAqzkDnZ8RhVEWYLvdPH7dUu/6nOhPdSKRWq0JzEu+iZ405wyZGrVQv4x
q9KWX8WEHTA8mlDHNy14+0L3c5h/cieG235PkDUjlsXKUlVppUKaOiO9r7UUP35RTQIkOthK9LVJ
jCbjTAB7a3E3n2GsMOwnVkRMbBiJ2nMuusoD0ApSGrM5gIN+/KU5IoISiLnt0ViCve+UtPuSY5nS
0vdG8KXpPiwKr4f6TqV56sdTqIX4D+P705Rl3v/jIGeuRABS4B67Z2/sNsFkWGaEpCdqCEJAc+Qo
DO4hQAkkqkAhmUMM8O+YCkzrRIqzmTEK4obOozgJEz7i2gd4cPWDvmXfuVLa8/bH8r/PJU7gAdyN
8viMnPTgIE7Kyxrp1pdFgXCWWvMXKAp2cYWWSijGDnPZMuAFRHQTQqN7MwJHWzSA/lYp7sZDj2z9
J9C9pi7MVPK3PzUQeYXAR2oAOSaW2/hrbF7UB6idX4CDxkWRIcBhx7sToH0wIN3X1q/e4DLSY1gk
Le/g5fT4BHOnR3QBiP221LEe5pWQup0JTGu3zYEVaao6INxMGuyqyKUvG10N+5aOtnvM4gFTmggW
6lO6t59v3Ewr8Yhmc3zz2iHwHtAHF/mJNtslBMDuaQDTp0nDcAWUmGvL35fUE/9Pkiy4dFR/Z0AF
Yr5lalwikNKi5tpICHP+Aw1fVnTFqXhz3005bRFJFdy8VgS+r8Qz+5kEo/whC5mZ5u0Hm+WnqdAf
63/lOiUgaPleArHx2hgbJuphFJN0ufltEfpxIekYa4m+gp1ZBuUPODu8EE9LjUJ6vuv1TNlU+WKB
NC129JCqQmFwdxfTnIjJ7nkTBfnWqoGqj7JronlaBwEojTewhUSsW6uB1QndMl5oaip+JwdRtlVC
cXpnH6td2ATxZRT82xhrcascur1SkzDPf8wcEa2H8zJeMUTvYYU7dcPST9aZHW8z3de/fbiZCK9Q
on931/yH02Rugz00lGJv8RZzOMUXBwmLjfHTeVn6fSzjoz9SQj0PsfQqirEazg5cn4cOqJrmRa4A
s9JESa1oPESuVXIp8CbouRBpLEvNOvtj2Po4KHofV9y0qPU1c3riceeXPlw4cv+xrK/mRIfZx4xH
O0dcVe8NSpalO7vNzp1+w+MuFpUBR96gUJDKB8Bz8IkbDkUyd/K4mcEZpP9pwHeEoLKXIiJZusDA
OJRDTMoMwr4XaVlhZv9+KjK9vPUGmvx37LTxcvxIXJSYil3Pa/DI0IUGRkYEUkWzb+yBqvnupvlf
G9trnK4JdIb2mwDBBop9UcCcsz1r1dhmOmuItOKDAkaWxizIHKGZIaGxCqD/IatM+mI6a2EH8YHQ
96OE4JvEtdXhfQbkyRh1oPMRkcwmDYBa+Uw9d58ETzKG5Q51Mi8moRcJUwnQDRL9Sn2X2El4UT1T
ESIOE6RvBENO3N1Q/rQ/Zsa/ZypMdFqIM0ChbYQ/jP4f9VoKAYBQIDmzZVA61n+/9e2JOVEm7hLn
mEcgQ/LsYTCXLUwIa72bz7MhFVH4qH/i7VJ1m+5sGQC7+B/ulqnS7lJLcjqZkCBXYkNx6zG53d0m
HFKnAuaE6kbdrirCpg4eEp5uDJjenRX4RhDJ7H8WWHJlqaM7i/ibtX+yO5WbSnhAJ9A65LJB6Hw2
oEOdBOv8wLgp9Iq+nIg1dCsIvgzqWIFJCJdi9f/zY57ZrKAoRrBCD23n0/nIT1XX1ohdbdsfJCD5
Dxcxp0CbjkW3Lgp1surbZO6Od6BELgrFc20hQ8ry97t1ItyRFhv1CN5RCrNFjqtLtb7HN+QtNsn+
fGzv3swRaysnbVzJw/wpOtjpItTP2cJezVnTD/XBvKf678yr/E0zD+ofs1UYtCXYm/4ZTFwnFzkl
XdFK2+qcSxX7xAl+nLHcJgo4rRM2dxvt95LYcGnBiIC+hLaFijyEi3BSOYLrpNhDjGZuhm4qdfHr
CjxtRF+qMlbWwdpctNeGdLBxtXFhGcMpvZSG3Z4lY68rTAUkyYUXV7NTf3QMTkCr3yVoPThTfU30
rkGu8mbaivrxU7Si/TsOvelfBkV7gTnYKAbDn9yEUzOmqmN5encZ7Pl/X339W+JA6C6CRYSEJmja
hcu6dQ5ZJ2iNkdGdQS5A7wlYucpZgbZpMtJ9FYzN6b370YIIEO2Bge8QFMQI+4uiDErxwrgCLT8m
KB1x24L+6LaGfWMXWSebTjWnTV5xFCU2fRVE4c+H3/okWCEfp/RQINAeu0hfMWVLu8DtLWnChw+R
v/KXb+0pYQV15ISzc/CswpybwZD4OmFFZVf3tqNpPH9rbljZdLW4S8cEZGPIyQpbnFEVX+RGaYTh
g9RwvhidhGTYtXbM90JFkrBkqjfWpPQzfe36TcnHjJmMMdsI3Qa+AcGwuXVuM/uu4seikcaeMP7z
Nr0ygn4oMy+jQWYfXcuZhwR/UsPQukJzPEo3owj3iLRB4dncvsE988UHzbuTz6quMjOEyVQMRQ1N
cTG9ug1eyTVfuyYAZ3Zk5PUpP0UP4L9J4obMWzZncN+8fnKXFAXjYAa2Vv5vpTUe9Fq330evjlI/
hT5t1RxGXKdLB4kGKni4jdleAWyVhm0oOlIQoPYPrbI2+0b1Wino2lgd5/i1z1oGQuBjdBjQemIX
ORVWYSBs/9u5S2R2bQIsfKlHZJvexM9V1sks0hQqZ5mrJ3j5OAAUoIHHzqoqMDT37j4RnO9esnCg
11nMjJVq/054IqRYRKvTibMJXnMg1VuMvbDSTTdzkxKAVm+jbrG0a7ew46PD+8plR5t2J9/H1xmx
gBGLXxCZ+4Ttma+Ly/NNZ97W+4QqVAps8WxSakF2SmVbCb3KmMjP0PIk1jdjShlh+teKpq3/Sxcx
FLzHJ+jSBcE4S475oFfdpNfIF970CP8x6hjy04VaKSSQpChFs+7Gjb/MtcQuQIkIvHCX2nH8Ob5B
CInvw19LHwQaAcDTr5tFkJ/re1rs3X5qnRqJIWGuxAptrDTiUbR/lCiCWsU8U2PIy1raSjcI7bAL
HMZEdIscL7dT+r/oX+5kIIu/fo/JmRhzwIgboDiaVL9tRQlhrX/o3cM8j9wXxXipB3NsMlkWU3Ft
HnK5f4o3cgjZfRDxrosf+xYyxGh2cTStMCGNCmuub/h71B5fbkGzvfyz+vAzNsCbsRXELYfbJG73
KZfKiTTYcB7zGFIkbtsL8CYfPuZ+lBFC/QZuikxOPAwNvNK2A5i0Tx1byo06Uw7uxeJCDDb4iGvC
67CRD2lHF5Pc4qRTeujkXIY+AG8898L7cWCsb1alGpZolQuD1S3tR4FqPDuaRcg7SAbb8mUE1kbc
7EYwZV71uQ6j+WwlBy1f4bOww9hLcgtLV0gJqzhrOileNuTRsA7XKFfo7qOMouSTkIkf2qpuH7h/
Blr+7D7qnaoZFbnVFPw/FpPDtEDMHqnUkNdp4KcKgLESveSAA9/ZwQWDXtYlm14N5Y/zSCPiW6Xs
cHau0ajuiv8NjaD67GKDWMoLuF4hDNMoGdNKEsjKePtBKd2Nzxes3FGRsne2qv/oUWukdTrRCH18
BZRy5BEOM4O/RKJtEt8najNtTdfZcjkFbULO61gXtoJ0r1qhVRqDokMr70tjuJH1byFWbSZyODuQ
d9j1FW4tYqNRRNll+FUiqe/iLS2swIqAadytWuDQ+6ChRnhBsr7utRE2EIHk0goL4LATgOMICVK9
xXhDAhsIBIwI9qNe9bRPZbdDFTnECtDEh6GIRvNXXBobbVHNeZIBzu/2sO5sK00/WYbkSnse0Oss
YRMVr2WVu9R3wiyr9+0UB6Cy4XG+VOYbC13AbWOK3jU9VAiDewAiDaS8Ja0YrJoGvbewEWauO7JY
wnzLDtgV/BLBlPlFXIldonDOGdN19uQdtfzExR0QewN/LFM3uFOh59Duo0BIfxKwiO3dt/H9BAJq
7s3k899SJiliwCgAVGvYf7z6c1460jzt1coLv1nlh9Rn2TFlQmRxXxgZMR6Hr82DLIcQgqjEmRt0
n+9PK7rc4TyMBddpfWntcl+TCidnGYxto1X2ghSO5q8e9csIWCp7XjfKMu/OFXO0mMYUA6XjOkcy
q2f0VoOIiaRSYDV8MaZD+mD1yC5Gl2eLAvOHp2IhXe3gOp61/z5kkIJxEznEcETUbGJ3SN7K4iMk
SYqZdKTbZA+A40LIid2UTSL7Y5TF9nqcuq0s4971z7YjXULSXvP+uAfgkZ1cAUOIqbHt9B17DDvb
lEXeSObPM+SWuJ9Eomvw5EmcaEELoi2VUTLo+t0MQGvFRgnjzMTDaLmcHwRsIoApxjAyBOBESwYj
LGGd/NB4ojGp4Ows1NfN0D2VC7FbduHlxdFZtT4RhkSCT6Il9mysCDktKnDgXAc0VDsb8H6KbEsj
LV1+56JsMxRr0RFF+0f40zwAoxP+5BCY84oeu7ZHMnMZTLd/wobLv0G78XNsOo9Z5v29TEU+qiR+
cEXFcd4scq2WHr1f1wPltEMWee02MWVznGLL/UlARbZphICV6Ytl01ntl4PRPsb2Yxa0qGDFsleq
BlsH2ZR74jtg5+pMeCwQvgh+OX2QaICk3epM665Mc36Ygg6IdtVwY7b78woUfG42/naapmSCoFIB
cf9GbZhHfCSg9S/KG4S3KqRWQQTAWLqPQ8crPOcSpvANJU8u2U95v9zxoRyAmoJEwCmpT7TGwELm
DTwGgwSfB1jrZy1bV7dbtAVJkopNkRIHZuecD5riOkyKGIXgb4CooIRwvn2ZJJ7+OzTZV9ZC6VkG
084BzdmK8XutAddjScfDpllYB65c5jTa1at2/YXB4ZGkt1eidNDvHw0Vjuo3iLQgIB/I5ONbK7FH
XIz9gSILrWgbQh3WOLw6dXbjC/aWoBTABXcGVhpUY73+Xj8scAuoWEI9t3u9SHNJayQ5MOCNTLWq
JfA2kLDFT4trSHMAOLSa98DlL/8iJgbSmsXCb0Qfe9KgltszVZrRVdba2UjmVSpoMbZUpT9u1tum
f7Ix/IR9ZVkVAQSpjalNMpkYxn5OqqoSXnvptp5Q8C3zSHWJVD2fs05DKOjfs56KS0tNuDRm+GNn
VKSr9DIgHUbyM+xEONyYj91hwqqPUYQRZaLkLTA9GR9ZvX+1r4lxX93NvoD7k+WTugIUz3jxlmsv
JmLy6JKuZg73qWza4RzHADooXO54s4dA3or30f/9Yl5T2bsO7vzGwm6QSpbO3bbJCXfKftfNJKzc
ngzqsBTz4VjPap5bwtLKIZmnt8Mc4QDu8qQn8wfnJuvG/9yo8ny5C1VtxSTod3L1dj2HQpY9D7LS
GFWq+AjUnSzSzZBBa9uBzB1Yse/+hkBjNnfZcgdJOHuTkgFQw2U3sXroDf3ykj6uwiA6H2TvChg3
Xr3rGamWbJVGA3sdMMv7gd5XDrMqACyRJ2vW85dT7W27E7y1ax9f/frUX0uL25s9OmXTCrjTjPEM
mZHXh9R1TBh6TgBc/chllCcg7Jyi+nwN3x3YyrSBXNsP0ezXfMCwfnkIcyEUzxDcUKxNdBy+DC8W
VqZrxTrH/RRk2DlJlFkJcE9zK6u4rjdrgu3Geucj3seuZwnrfV/TdNouHbP9UJx3XRsURobe/IgO
U6vAe40Xl44hySYjuA9S/BNKubxFQY3834D5ULgk/MjOAyBZEhIkZ3YOUSXxvDRpEDiUcjFuPE3G
BmPRe3bMv7azYcA2lIXgfWJ/UfyQiUexgQ4YQ9fTVWCqc1awSxZcw7kru2WQWzU7N5byWUy+S/7I
26y/A3LYXqavS48EW1VwTiONk032xebc6M42RQB3wiXDIlrJWMfU8lAwgfoWhIEkInTX1ykCQ3sP
f0hyuCbTnKNtGeR+9/kxEzP2LNWmL/x/tu48ooQ3zIbC7P51Z4mAEMY9qJ9ZqlsZ/5vijQc2K9pS
d2xnnnDdDYx5+Q/n7z6Kg+aatV49y1ZRUEC4+eE2nfUHOEVatx/1aKlxchLzQanYCKELq4Uyz8jq
KAz2PMu8h4Si5mrpiFXUyS0zSyhx37YZXJhOtWjqb72en9uNLrYKzW9igXIE70LIJKrNmdJT3cSS
sOlF6OKRxue9iYHc14oTeeCXRat/wdrisoIiZiD/4pMCLeBdsa8sLbTAkLpeZH8PW1oTqGwcrUY5
2OFEQwBEPNg+v3fi3ZHVakV+2CXs15djUCdaxckwpZAZld9DTiyiQuieV2HUVsf2v+7yrYQxEyn+
STLNp3GfbLFBDOXzYAwyrG8DYzGJz7TkHStAjfPGilH4aEVUtT+ND7DnAw7uSZr0V4L5SLXrfAAW
mKJoBFUG/3x22iLUC73oz5uHFw6WkLKQEhwsuQ6fSXNO9otlb93+hVLskegvu/VOgGJVbHLK5rrI
v0HQGhnX5EojtwW5HbPd4HJWsFVugAhXfL/AMQSsxVz5urVUSust34Y/aETtk7DjOeJkPH2QiYbJ
bu+quQScvAxVBlW3y3b/IozFP5aQ8zUCY4LynJPDWZGVw54fCKdRhf7cZcsms1TWlT4ERgk9t9LH
FXdWYICsbxrG6aVlpvsA//kZ0hO5cVCopEi8nxLNjNNQRIGyifMhTjkt/+VIhFzByf4LQheUWcSm
xMDQDWxcLfD8NJAg9zlMuI+UWRAz4G8IZVbnGcFMIJSrPftyM7jNlj5/b+VCVmjhNpRyC0cgxAMg
WeY9m5kfO0jjLancNFbwkVmW6YbpjLORLEPGyZWLdJ9HwjqA4dMZy4ruzRQ/V7CuJ+2JMOHiFqMe
E2QmJp1iRIlLkp3wWYplZEzGUaqUdkTModVMdR0xxv/IPdtRywnhPgN8pA+Z5Md3PEOaoBY34wpn
c3u0u5tCU48kVSjFK34qUZCBtn/oaN73ijputf3XzehES56hjBkPNjzPyb59r0ogdOU4L7hotMKf
T7k/09avVNpAScUds87sNP4y6aZAptAcsgGNfeAZvDtVx0qmIjUr3ztOpJl3Mr+YW7KFZCFJWu7M
+icUBBg5/rEcyk9/ad5V97NaVCb2alTEDclw9SOOJFebLWDkAbT5B8sdjn27SrQpzusmEIVUAAUy
tCZL0pYKsxa6KlH11k0c9YQYMGahEH697e8uDYfcKZE5tIBC5J0C95BpA1N8cePLj/5eGPabLE6q
kGvxvyyEsBcbkI/R95P/xU4jeFuSqJV4/g13hcJHO/jwN42EsRxICALRdfCcuFACnFEHtqzccJLF
P0mLtAUcILv05TxDeEPSLfJbFWyhT4Amxa3BfaM6OQy4tuJnLEGuqyyO+FS0XbsO7META8A0YTGW
9P1mYl7yoO6VCPXHv3vPYnwCIOTyjHhrZZMBznZlDZmdEsQVxv5713XzQ+G9j6tIiWyZ9Zr65ptt
XeYKoSynFMLbzNKPIcXLN+/sqVVocDuAdGqwwf6H6Z3hxGzssUZKCOG1F0sI3XNKUG5Ywm1dWxxb
irgLSQUQ0FDAobIyG3y9SG8ezdOZtkdF9Oi8fki6HyR2l+szjVUPTcS37WUvD7MgqsnfMJQyffFS
JX4NDQQvgQcohi5T8ligv4SgDFBc0m1xccuNsabuPDcHHmZ2g1qTOMFmOavTkCoWgvedEkpwU7DM
iNDCmu/OKl1yNpKqh4CjXuL4xh6+G4h1wED3bpGzG4Msf6JAqQYlikin3qcHOxjO7ZE5sYuDVXTj
IIAhdpwe6QtoskKr8AdXz+hKvZtD/JV4f0r5TNsNPfJubEzDl5ZF96TfcL6X6ny9PasMQA28G7Ti
q6RyznYgWD69WKB2p1G0EY6r7XMcU4QFYFx+jxHotutZdga9kb+f9XVopWFpqFl7ZvKvdbDyMDRl
1U24wIcHa7WMBz6n1NrS+b9mm5AC4APSpMnAPmgFPDF/qpBNXfA445YpabKIVZPkjamb697jL0vx
Vm/1odSAztBPW8Z2L1PaDEkwgOnkO+yJ5ShPmOfi9f01E4PeoSe5mw7XQCR8TBjXxmREBZkTx5Ew
gmbMPEZgrZg6ZaF3WDkBxx5Zef4OVVd9HEBDKRGPfyr+bsCA1gwkYybfDePA7v4BcbJB1Afyg+2T
lL06ojKy3Sak5PzuAb4fMtQsyaJXVV8TdxR/TkdQsOoOevERe8EiJZPEOugxouVVb69hTvHqPb5v
B47q80+ZZK4lmFLJEWg3XmS2TWlaTfTkSDDfzUC6cQ12C+kbIBwzktJuOzWNIUX5f0noF6ug5lcV
CcqcIOBchgmVeIFnn0EjvZBXU5pb/7QioKqaNUjhkUf5wmZNRFHo686dz4VS9KZ+jikDYucw4/9v
mX9/q5CV8JdueVgWuZrUp2hixehqAR1AuJbg2L7oxI9PAHxWlmCRUusgHq+QoAuL3arXM4+HnvJn
PkxA2TxBvd2yG1OXF3pSoQLTSpCxzfExIBQIGcTKSkVGMIyqQrenx3XN3zciU5th1lxSK+fad1yR
XvND322NU6wYMWa6bZz/sLXyez7Glow9DBJDZNgqqlodbVE4tOBHXa9nG2rsCO7QahxzS1YrM5fS
XmKGVzZJptNLi3g4jemkbfHWEX6MyxAQfwzX6zcjUErZRobr4oEBO8gr98w7nG5O0FeuNwERWApd
WC7owLaTYguQ2hqkU8xz03blwPzYoc4D21sE9BGgNdKRGBdDPCByHngFL64An5uEynalfzzL/rsj
UnKJ3kmhHb7OJgNvW4Ggsuyshs6tfgT/s4MvQh9lIraBH0JOa8hWxaAuNCMHW+mF8lNIGwIqVoit
tK66kkc5SKyyDdzqKXG5zknV4v+5zyY4r+M20Vg2ZRJn30udyzi9Tv98asC9F6Lgzvc4AWHQAUQ0
IZiB4p2tG6bbyxAOBqdjs9on78U66WATrYSnrb1+VWkFMQ2oJPMt5gXaASqMMUmgyFCAJPF/JUkT
dAE75dDGnA3VsUyASehEdMDOUY0uMRqBba20dxi62r9h36IVKbn/BLwaLdtj159q2PNS4HwX9WWo
sDfPd7ggk4kR67ikQoUU0jvv5A+iCkw/nmDjpVGVxkIhcldrmWq17RkhJCfpSdBVl62p+CPHJ9Kh
NALtbx0vSpXl0Nk/5kdAciJB5c2iVAdrK5bk9w1oh+pqDm5nX8GxTTV9bWNjhRDAND/b0Z4L+cx4
NxdKau13dvV/jZ5LFiaZKx7AKvBEJjZjXrml3t0WZe8AYArLaQ1kJ66OVFkCVGnAxuNkpzC+8Oj+
GM0NtJKlYtkzjUcC0JPmJzZA73DFTs188xtHhBgxK7+2q0jp8oE3W2DtetNWTsKve69v2VjllecF
Axu9L1u16O5V4u3m+1K8SezYuBHCXg+lnY/nSgYS6+18EjIVpfpp17DUgkDVgydtwp+qwR7SOSZF
HVrOxbO21qoQLOTivYKet8c15XCdHg/khvqx12dWjPJfCTiVSNWfEaNaMTvWR5v6Sgm7vNUcopY8
THkcVCFf8kAwT3vwScC3aRFDT/3KRwJYO3czyd2ipsJGKaE2DweHbCXXV61oKslTyHoQaCosUapq
8C4UiC34wQXUdsO9cUKK87IH6rzDawEUehUHM683eIpmkOqW3gD0fG5SSpT+gwdOrBvPK70Jn9D7
MhQS/WVFf9hedg57TcSKniloheUocBtT4ZsvDrXhQT0Dw+oViGTPO9a0DwPMJPkIqbrKniQXC63C
58xIL/rhH3AJKU761M3PqNIzrmIw+1vflsLHqiGmGRc1ckyRSBahDjwfdIzyHa9WxF8dSz9ZV/fa
wN2L86elQlDYuGbEs532TBWgUE5iWEjXDMONM8C6D9IGZnCliUKLgO3uuMHoyPK2H9kSv5gHAoJ2
6FBhOhqwCdaZqCqZrigwpz5NbYcWJXFC2lUtMvCjoNR5GOhzW+eYKqyMvvNJR7M73Xv1JOaXk/w7
rGYb1ca+3eo9eGfJR5+jw/7sUj8QIklResFd7UaosXub+o+/xwvvRuh9cn0bv+1aZqJSX+RMFBcs
GLo5SeElrYsGuwjkemQ1b75Fs19pbbNveU7EqoifPfr6pwwLOGB1deG7rsDzEXSfnnKBOAnYftFx
OEAcvDCvZyq+5Fs3AEpiXOd3t0bhZ67Hbj0u3wJO0Wk+rk5QyUbn7lkuU8sn8+Txg87WD/YseL3J
K4ZA+shN4ndxEbhmoSC98EDsYe+aeYOFzPeZstkmAUCaiEUN2gwEtrF01oLUNT6vQXddAXUGPAnX
QbPlbxBWNSdmRnPTYETV6qhvFjkSm1Amx95LeDhHmMVFzYtTYOUUwe1u82gyHZxhE3VvCxSYH47b
99r84hWRkHyo1lNY9gX6E6JS+nlVAZLcY0wmWBhxnPWhHWvITv9KG9Xf/lM4zSaavEmmaqW8YC9A
eO16VNiwtNbDOgG7kJyRI2xgaR9m/YpPl6QTGgWduWPSHbJyJM6YAkFBBqbf1wUG52l3DG2VvtNm
4QnnItkDm+ocGde6sK59R24AmNXzFzjo4zV2vidFajknA1J6r5WHPxvKh72KKfy3xP9eS4tAoxhL
cWdt7mGeEBZqTkXStqcmJXYXeVm29TThuzSLnYOQf51RsZE/V/W6YOqO+3VMuZ+BYlkrMh4PiVfG
fbQyF7MeMKDa2Sqto/47L/1eV0o6HkmggrFhEpMpn47F+aL3kS66OoSy8tVA2Yc6rgfODRaRwL/7
Xlh1Y16KzlkGmzevRZmQIJ96wtvVJChxyfEKLSHjf6hZByhcxK/Jw174cMXweo11S7XC/lwN8qhg
SbfhLLODM3f5Ktn5x3uivtEfpx29o8UXV84flohYTTNmaOAI9bNT3SrMWQldZJYR5J6bpbT980mc
2HanKsDkujPb0ErzXygEWVfj6t30bMR6i6Zvj0GD/BArIE1xiIePzjDFzmMEjgKhwDDTJ72iTHW5
gLD97/C6VfKH04tvr5/dsUuAKLh9eSumw1tI5Ou8C/f/56LhOH3ag4Mu16oj2EPIUkFBxF/j6ADK
PqUtG/jS+rI+SuPO+hvfoPUqmyYz0jS1MN7OwbFNMst8hrOwrP5sNGQZpU1NfkRKGEb92wSD9z8V
oQefUf3rYYbwlo0u+4f5p0ZteRnkEAoyUJfs8t06ITbXatBmjYsnFhiM/jRm6llafpttID8iQ7D0
rR2ap58cYogpwiM0++elGomreAyXJt4NDx8jnmtWRLoLmGnYUlsqcNeZu1SSzQJIgUnWUdvdnBiZ
qkviMZErbdrJSBP2GRmsW31otwjLbk1GepfXIQ8jnWF0dmcb3Eyqf0YxJ4LbO4KRwbhxpcHMM6yf
sqdU9G1jXPdVg2rojXGG1ys/9CcTEVbGEb6SkN0Hq0p8fP0T9v9m5kBqiKTm2rumaBiyjT/hafjv
vY8NYMoGNgOTs/kqv2jWRpEKvQaAEkIlcYDtWsiL/huNbBEGRNrDivtzota2ewLz/rzWk4G27OjU
53uf4OSOTf8TCF5mHqTDw4wWE9BVaO0Gv3OmMlCwHV0mwGlgREtIgUDp7UfKokaFZCd+GZ7tg/4/
IpANPMESiK+OHO/9fCm0jdpU3Ge1kN8bYLt4AIUGLpr47sqGvJRdF6ocwy+WHDn/M2hLxdXSVEa3
HRnYgtPIifN6r/mBde4JiMVygDO6RRX/gplkyO2uvDutQFmPsq9vN7NIza2wnOPI4Y9MCG58Y+F6
Cz40IQ5R4cF5sOl9WX7viKBOCsvw5wIF4Pzk5TVtdgA32K9bTE/ALxauEVEGXLNUB/b1b8hk49eB
WDJ7N7Y0T9W3jy8FeKy25Bw/3b1mnIO7maKnNFtksT6Py7htCfpIug14UDSU5pUre1NYTRd8BpWR
tHlzylZDklX45ErhRYkvM5ZISNyVbLdijIC6Fvo8UTPwB2HVYNDZuO/lbZwoxEyGray/yT7f+zcl
hkgyrTRQ+sVmprKSyC0BZsbtWRDwMKav6H+KfbiK7I5j4+V26OpiVEKzYeoMr0TAoeTPv5bPlgJB
ev+lcTVv6MiGey4/7MQJRUq126iD4JN4k9wjd71hTgFLX+shI7QDcEleq+0krQ+RewAoiujwj7bG
IcC/7l7PhwOZ34xh8CJRxwp60srniK1bECYFfNxctJ3PDeTuHF7hR87IMSI2YcHHUnICYgqJ8ajB
gPU1xrdoIicIQkPz//AmEibDosBbxmHgKUrcSO5/f8Y7vdkZuRhxBc+6wFaNky/mZeYVHCEUuZdW
nSoZCnE73bvGfi+GLnx7hyqVH+SfTjESz/c+pFffqQ78FLPzdNl2NrXAOzp39p7uzk24z0j7jueQ
gJUdbiDCkGU/xMWi6/oqy1Si3y8NvfElS6o1LPwh9LT5fX2wAnzODgVxVcW99PWMVncrBrYhDlrH
t/nU5XURVilblChUqMmw+c0wkqmGFasX9IX8ctdokpEK9jaHUReR6yWQ7sxyEnIRqCNj7gCDFRLG
Vw8XCABSCMdkMvsQYMx1mjpVQXZ1EVNhHD7xLmHbvTzEpuzWKpwFQd5QWl/ZsD5ZHdv80PsiK+Gr
j1Bn6YDUPg6+nk1+RjPIynPDtnTdUXpyH4QOJsUCrz7J7fAuWUak7WLs0vYTZTLGJsGyuM7ieH5u
dGZ33tpelyIlvr7C0xoSQgSBzhOdpE3zzY0ulLwJfNpSc7cIdQqbnag44+MWgd0KK24c40QPmHiR
H9di4xV/NI/NJy3aV8RROM/yLCtGwDDzLGKH/UFyqoWWNuKEJVfoOiNzASFGP6HEpvemE5/LBzZQ
dng9kcooM/5XlM7vTp5kId5ZJH9ux8LqXCYfUgvWUwxVqKMGYd8HQVHN+Pup0J1anLlBNxnOVpkw
qm5np3plRmD0VJPXAhutgA8l1Exzy1C6uahxD1jANldKlB9yeEwgx1fWSf7Lbanfe3OOGelDzFsy
adDN90s4DImkI5aZrDsZbl0Ej2Me0r2AlDFawnHOqXgWGSzlrR/SIdDegh7TU/pwvHsuU5COe+BD
ud59nqdNWMOiKxOCG9GyRZpKiSOcj49dtD4oifutYkNhbXGksha+JWHO1IM4mcydvDbtxoYOUCAH
53R0M+leBKm5R/0z6jru+saWYXnHza6dLjehhFGNossn/9aL1AfQpOR4pYcl5vVnZMurPh0rIssv
D7WjNP1WAUZ97NXpdYCl54szNjiJ2O2XYmbSNg5eJBKTSRxiLjmN1NsTa2XHRP4GY2XxR1Kd3E/1
y1DMCkXXCyxZ54s/KhZSBrX9oO5Y4hlRdfzZz51WOXPtIuGfgXqSaDvT0JjDPghrT/uGdOkbKgj0
VL+TCxAyeZT0w9xADQGRn2ErHxDra+Ax89XN+1O3Ljf4JYt3ZV07OYOHLRFHPHPePEPzakEqj1AA
aAnWmBT9JKsNObImQTmrkGktgM/czpmEk1d/rptVnuR8eJYVx6vONDrD7qllCmZH5rAJdhVDmUoQ
rid1miSsKGaeXLWGnP6aSTA/uNWOtfCQo7fmxwCBL1HDGIC45Kcay2YHwt5TbRNyhfY8ntF+O7oK
jd6G35M6S1jvJMH33zJ3JDLpPKWKY/wI1US8aIZ0/1Phbs4yFtcezVvS94cqa8JmeHkR9Akknxnx
9LjBvBPw8h2adVIVmOdr4yk+R1UT3DvQN1now5K0wGCTOKhwsNe66OLK+cDjtxMe0b/SSTzubUZu
q0UJlKM6FOFG9ZV/0jps6crBLFSlcAj914FfAQmaEMPbFHIFKkTCOoEsvBZyHUb2QMLqgmCv0EX2
JdSAEOMLxPxpbUhek7CIvyZuC/E9DTx4WuFiTdC0SfGPG7wwW7KHkT3OY+dXkR69b1b73CaEcOe8
oowTzO4OxKJ8dBlskvbR4qSf9KOFIpI9O1/A59e19kCV3kIPj7kOzu74lxymHtnteDZ/apmib3IE
IN+M//6EZP/eQP2XvIegDJeZKQ8K8nbXmCz1XjRdQeXFkXbfOLe88nM3jAe7z3mED3Qy8AZSowYs
rVGXtf0TulNdYA1O1Ayj1c9ib9CwUd63Ont20T1zg6TpRdiRCjhPNuWuWdBFBhZHeeYVaFCx+hy1
SZqGpIdTu1zSOfeCPTAp+W25gAoSZaGxajOdrapvg3Iu7ln3P0II7zESP67rQupZISZhqxEbeZ3c
HzRtpfoFC2etsfI6FGtg5ZZBNMX2CyoNH5hQEpuqa3v09sovDWwSVsIZqBHwmHWELA5BAsm8YzgM
2TT0592we0Uhjk41ESIpJGZUtQ6GabSK+iVp8EECtP+qgEC+ak2jQErGUqWsdZhp+XtOKPL3hPrG
HRLS5ekYq3QxNXha3MwhSdTXKOsWDkKfe4e1BjxYfvxDpyOKjNn27vMGQnd43te/7uTUDdGmM/zD
fIyKIni5FG6hoLkn5tbpixydTobP9H6AOXTbPUM4xoP8f0eS8738TIY2BUSImy1yGevwjaS4FREs
f4T75BQ+Uk71jfOnTpaHY6JFiKxJlNloggZx/iCxM62m4755CBe/7Ibin3d2EteBQOrwPh9tFLG4
hxD/cHOzCukHrucxP5lzrGrM4MBADZb2maIQfaC3+D7JOANihNsAmuuH16JEQG2WT11xp+/bmYBy
WHgIARNLwEdZpzkJhC/JIl2rnUiMXkdawdssaOeIrgrHmgbIIvAtcGi0FLfPTJr3Rrjk9p37c8qf
qxFHsknLOIETCU7uC4vyadPT/B6BaYOegCQbVNgbFLa6s+pBZtIGNRrQKyrekQd0r1UcaHnEfCqp
HdkVFDWAy5vAKsfykJSvXK+y4U+rObzXGu48yK9J4fAfMMEG42vXPGPeRzL0vHZu0ahBZjEL6+sU
DJvew5TBkOGq66uIoHIEPM6wVaiLN/x/yoLh80hrdFPR2JKBPbNwdyFpUZbWPZv1o+RX3Kil3QPa
VuRRv6I+6A2t6ckRDnuzWxBgkgA3J3jEC8oTuflSfMesTDtcBf6pJM3QJHkWtQcUNqQNuYewcH9F
4HQQwrY+eIpTLe4jKwzzCQxoUfZdntdbkKwySCEvnKNkuJ74sFe/hnHU6YNGcQz9O6GZxfKtcWwK
0BgSxVTSffrZQpuBbO/xZFaeowKC45glkcPk3pdCemxCxfirWmS8wjGywPCx5niHiTRSTeHf4+Ia
blGwFD23rhlXu8pLv2Ri03n4/1wDjMoqiTGaLsO+uktlLa54gLW32DAlhTuNFrB4rkptLgh9RbqF
fnFKze32PdueOfoY7fhgQgcw9rlyynspSr1aEXrbjPBgrGjxBpEGQhuhsxNYHl47OUwnpg0NJNS0
HprL4ERJD+8D9MdoRthLzckpztezOzez90SPLCnGYdv9ORWrzlyk13w/ril5II3apt5yDkwVRH8N
8IpglIpiNwtXxbNNr3Yyg59BrzyoL/L68Trd4QQ7Z/cNqYHpq6GvctEQgNRT7DaewS6nFU4QvyYl
j/JuC/f9Zd+vHsS+TOi+DK7+8EW3w/TizZwD9qlyxCOljg==
`pragma protect end_protected
