// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:52 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
ILKgtPC086EcMxO3kjvgZ8Jbg8GclE/CGFVE/oZ+85RSkafKp/TzcOcKU9AnSfWY
SOz7Q2hHxwGCwNBRCpTxBCbjhpeoWNNDPC9dOs5Mnsx3Ij4tHedITDzgqYVMAmhu
1+vZAlAPzCsCKLRkMuBpaVCgP9nnCVAKAt4h67DaIOk=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 4928)
b0epZgxOheAy9JWyGPTM5etENZCdVb2EdB3jLNgqoP+G7ffspiiSegBHh0OUGicO
xgi0PLLtwuL4w1dkYMaabK8NGmrIBrL982Nob4xKF8cSX7+icLrGkhFKySvnAAZ5
5l8djSCT1/mYqvDMMd/1rn3uUrs5i4KlVgs4akYgXDqoCKetErWZIt0WUkYZTL87
sBaxDoCh4F910V9pXz8vgLiD3V8dm2k7kBh9k4XAObOvXKUmkoB6tN9x59ZrPTAN
3n2nnT1fpx20N8Z2fkoU/zq2cVHiyL7Zilu1v9Hjz+6zlL4lj2YzV+OEif8ujUEj
pu91PzfG5G1nMNcEsEkPrTqZxHTMIp1QfAzBqCKB+6G0ux+a19swEuyMfaOPAwhk
uMesNfdwNWuBKq5qdZqus6ZIDCuFQQ/tLNDgEmuEL9eamRpyyA9aU+4WZ3uCSv4C
CbgwKn6pwCEK23O9h10Zx44uP4vII6eEgNRUyhMQpHNZFFhOC2cP41LrS1eD9XQp
H5P5Pk0jA6PSHFYwqJrVCxYJLJl1/C5kgzjsaTH+Yxviouqyc031dBlGXF0WlLGp
AXj4lf+7dDQoPjh5R7OA7215Qo3M9rFc6m1+36V+Xc9fmTJaEnQBCsldqV9hwpkS
krQXIAjysBMvqz422+WQMznHLOn/3ukxau7IvoQ7Wy7137lSASwpFHZp6TlyOVAO
QcVPAVCkhqt8KzkRt99t8RC+dvnJLn5PVq7l4TLZIJrnqk/OYNfOCc79Nt0fFhzM
Rfg5/e4ocSbkN+oqB/Y0/O+kir2eIFkCpdnZUHpxSlh2ID7xIZM0bNoNXRRnZkhV
6A6ozZBv3otsUFrI2xP0cuSvagg2sEJ58tH+1bNTns2EyhiZ6sUpAba+AkTXHI2y
uwFMYFJvQjgrwDxnqENqcW9lekdEuBd/mc+IO8reYrigPhf18LTXHXfcbaoGHhXp
Ph+boIUIJfFpmNMrNfCh/LVnjW1A5SdrwcFeBvWcHaiW9AybjGyZbxc0sFQehHQs
AlU11Ysc/XZUxpsRl2HuQGcAD0JyDrV28KvXa04wE3w2LX2omiGt9SEdGIdLsQON
wDul+Boj4SRyIwLsLGrHvR/I4bGko9waueeFT9xhvUwqFBESYx+0KIxWW8p5otDD
Ms7jAKahCNngk4ZmAx7IomMYU164gfZh2Z3gUYFctblAqNd2llfYCU8u0x9US+2m
mVTt32+i/8YIG49wbvnDgYnzkA8P6Afv9Y4vYKZLOyCgR2qBlbrIyztW9nYbamKy
xMJr6G0q0UoYU+zNd2h3NP9t7qPFRbjj6Cn/Db15VvgNoIIpkimjjGwnIuUYiTq4
BzqZ7J80gqqaoAyPldRc+UdpuZF9Q45VP+PmgVg019buChTy4PPBwKCPbG5lw9kC
JZhhr5ROCLdmHP4beSIhRpaFdVIMAiQZ0kuYqtIioHm55fdM+hHzaSQAOXgf8izr
gw4AGA42z59I39ppEke9O8DxRC7u60HxJeRDD6wOwLSnAcin7YCbrC4638ZZ8gQ2
ZOjf8khWYzySE1anlEweCEqtTN/AdJNDs6Nw7rmbvj9pjSoy/Gl6ol5vnH38rBov
DAeycG0O8N35//s7dKWiaI4VABRoOWjx77qtvMVHZErFo+NyAXw0ZXnhurDT6Vyn
uIagGu1gR0Ca25uBwZ+rA7vnk+ToZmfSQucbeVOViSUZXPbsvn3scJca7MPDhdnn
3vTugNC1OT5z//Ws7qx5+ObwHrnQ0V7cG/RrzEMqRuYE63uyqXVLEmpTLVzE7sqy
4Asw8eOf97209YFWsVC//jxDVEVpr8qp01oZlmEswGzP6vFL/dMsP3ziWztNLJJA
kn7Aib2nwbrJy1/ej0lDUeqI3U2OCSSXyL2TquXtE1bNAr63limVN2zFy+LMh8hn
an8zPISGxUwn7jpK7IEtS6tsnz1VapCDOwbKpiEZ268Tpm9d83/ywvmuiVpVE4yI
PsWKxDCYncVNgp4mdVYNW/F+l54vnewdL8UKd6Dq+PbowXCRpDYqWqtXfHI+APO0
Rh0e/Q+iGX3AE48RP422cBfGT5rAJ9BSg8/YDf6tBssaC7teHWwQMe2m6u5RKSJV
p+FVOtzSSW7YH/vgqzjmIbDdzRehksIKYmpWQm0BZPFYtBfSdvuvjx1RasTptzbq
3ZtsbCl0oxgohGhCvV7OFvoSTXpuAKcWup47ZwHqz9OV4M9RLSMiwYVHa+T1MZlc
tcumSjDyCnAHcuhjcUgSi7St9ba3glbm2Z9CWxUrOe3EXS/30OzE955gl/e/2xGC
obvKkGTX28hPPDBQKACWlIm1T/XD/uZklKgxxw+7Vnlro5EQcL/NZKyVP7R8as3g
DXh7Z6k4+I96vEUUas1z3RzwHp/IwbTuxOQ3rKFzsTbPVBilntMhphvzYEnRe/Ez
HqaO15NLjnIFwvsJ3Ia46LV8NNMNN737TEQWCKQ8qnhwiZkUiF2htP18On8LtOUM
zxDOLt84QzxP28bpBfU5Lg4pN9EbxSQBV3+9JoCtLADuAgJM1OZqFZvjG7Y3ZND4
Us7iV4t22a6DCF3sCAGYo7YNZsVWBLc2yyu2YZXB095rDhC1H3r8mfFSEUkoS0do
CPmHl5T96FHq9wHaRmjyE9lVsk4QhC/DNW4B0hU+r64fe++QiFfCoUE5U3+Ni0vU
Hh/F48FuMjZG5EcnOLfNM6Vm3UkJREBddY+bBqNSLRR5mq5ZdqgntsXbUYCvTayk
aTE5JZpOSvJLAjutoBPZHFgU1Gx3onFJyTrx8t5dCXfjbnbS0F6bZi6zBAn1t/UN
WLSrMIRTFtTxGNfGRsbBqD7qPRjAlwOGhbXZXR9PENAFhr7VyMbTW4Eja6BPQ29M
ldqtDuDZagDVN5dgcqoLz6PZ8496ASfyLXhiyE6vGhmmNIXm3Fp5q5Ld/GY5LOVF
YDRIFcm2l+Sc0WkCIpwkuJ4QQS0Ko7ialb97DrzAewR61XSqIDaeyohyvSo6VKmc
d48sH0WLJfUDI3JcetKFHHghMY0U5il8JTTFYxnSKH39ThLQa/3sgRfwm5a5oogi
K6SujfR4Lj+NGl+UcVHfY9oEhaEWyIGWXaXDjrGVNmVkxR9InjL6ypVjVFQPV+ue
M+qSceugoKFWxZUuNwiSyp0J1N+aBUVStrt+t5sjhEAEd7N6O+8+RZFQGwr/V78I
hfkr+4AKOhAkezZQESj4KkGXzgyjuxm4stj9kfGVr0uhLZY61NSrqcvH9z45P2XE
6yuWJSuTfiJe2DWJVHg45PBDShqa+9UG/sqaBqeL6GShQI4Da6RhtkGKGiZ5dx9A
dEBC4/6Be0GfsWalj2lND5y9QHt+JlMMvfKkbhcYKjcuNcG/qYQswTzB6DyaFWFb
k2tpXFGAYceAScZM+76ZM5Lnfe1C4xVHxLB5IT/mJtccrhDR+yJ24fige4PF83tr
3DcunCOS9eSKqQYgXokbkLhUsoyrIJSbpOx2zoLqwQSHcxWrK6PDD4mSp5LKZYRW
xDPxCCzR71vFgg9ASuVuC36Gg17mFX7QLzkQ+jeO9h6yOub7mVAqKTpaZuxu1t3T
GGPewFXHf6QKJc3LWiWDyaSv/DGa0yXYTVsFzUSBqTOM7si163OF/YxUrhpD6eol
Cubmh+SzMaA6MnE0Epjipw9zPi+yMiKgJRSJp80Qvimv2aj5KfCvaGFRqYMbt/lu
uzoIKoSNwv4UGSr+Gh0AiZIDAFo7toe8fX8IU+YaT1Tms0FocsZEKKLWNQ0JdhYL
Hp7uoMVTtcsgWjUsTWXJpNVbS6d2j89uSFj7aVTndSSCEAMTjl3/jeplpm1mdVDd
KsOKzTWO1WhsHNCuBvP0TcGYMjdUn7IMXPvW9nir9+TV4CCityXEKIAE7PV/vzGZ
Q/rZereXvlhgaMYpzo4/8KjwKwh6AZ3aAU5K1MwpNINEikIRD+yysBvf9CUbqQdK
PdX+B1bxPo7fhfS1TFk6hpcCCLlVa1E5a6rw5gBS0LG05MkzvsFWA5nlPF5K3BuM
Y+qXc8/AfWuTYPlKv9XwaBvRcj5xFHAkNhdE9xlXuqNQfIcMAMmQY9tEFsL5OHGg
dz7OQUw/zrzZiAqrbW8ZTwTvjqVvYa/3sCjVd5/vG0a2JUY7yVyEj0mI0RU3+UiI
an4S+7NNmh6AHvR8LTdd+Hie/S5nS5AaK25AB9YaiJSqbItMFJ19pMX/n0TPlJWS
JDOxxYOsfR+EltM5bPS9Hy94GpZqEqT+cKvMFZw7o3ecGyqyJRpX8d5i3lt82O1N
xIH/J0weva6H7ky45AKOkAUGwEA6britket7xe5mDBYJCNGNllsE6GGF5dXwI6pA
8d8QVGiVi5XpRyvgk6zpiZEbP3jgee4VyiC8ffVvbGSK90hmYzob48/TN9hmd/Nc
yxzsMn4a/jiLLfSYnCzLhkf37zUvWkkdWZDB/kCRwq4emjOxNGbxAGBGA8+LY6Ey
NIvHbS6MxEwfabCheydHso9pT51wHW/ZdK3KMk/U+jjYNTe/dOZDHbBSjaU7kyqD
60h1EFHaE1+BtOnQU203sfDz/vRTYbc0PGeDm35+xAqCRfCmpOb5YwK7BVNyUnBo
yeuPfr+3FTCE7uHo04WPWlLddj/0jHtplQRQt3V5wNCO0/rCvnIybkiY5VA21sI5
1tBorjz4lVqud0uKAN5bMADcqqnsijlS8D/MMJxoKZQTkcmebCazcxqqhBGCse4u
LcnEHv3mBkPFcj8WZrsBGA3W7vb4AsUMR/iRLJx1mDN+vzZbDCb9Q4v6+wgXNLRg
ovZqbC+NLfVn+2KBI9Vn+BO11MHDkjzZfNPjxIBlp2BQG28042pN/yDNIk69LF9g
s/hIOFSAwZ+cYsb7AKkKLB5+Lie1SMflSuBC16zycf1sqETWvArrFf8GZNCHk1kQ
lo5sdHX4QA8TNMJXUz6QXSYqdrzE+cVW25cwCXGhBYmBjZnF2mASlkMH52e12pZ8
pisAnFJw00157b9vCaz38wDQ7AGmjLTeAZ21ns6F3qGdNtiOjQSsd2YB4ZKkXysf
u8TACU+OMe1k5DV+4C9c4NL1rEfyY80c7NJOOL+WFOo+CWSfU7OXhZKwWfyGUP9d
BUGoVzliY4QbJljxUfJ3SyLxNojDcLrkgq8nqX7iMJ3bF2L5a32tMPNQgPutKlih
7QLJjNxR3RtDjx+kcw7+wHmZ30QOzbqt1rDFVBa9yPYBwlKnPGSsz3iU6QTa0HuC
dZHwL3biFHr/sz7QcgKV3jgG2ka9KbveZo3Enev1Ln6JPtSPY0P0qZlEipX/s+rl
jf+QF9ZW9GHIbqm2B/dXe0nHcg/J16IW9q+zK3GIjyouncr5pYS5MvWbJDvGf1/U
sJ+kfBfgD+7pgUkynRVKsfHxzpmAms0IIggyh/Vpct6cKG49epoH5CrT0XBT6CFc
LJGeuA/IUbjZNwO08kYJ1/hkhTJgCmph91h0ggvVSYa1mq5fMIf5VuS4owjNjiCH
7CPtmBFZMhmwFim/UUqO3dOz8Ibnz+iuGyoH36MSrrtxi2hI0mJNlCiz6nSTqdtd
VBmH01RAmNpQQByVVrgA6IkKJpDvnbNCzn0W+m7OqDG9p5+cLTXvN6VXU0W42Aek
MKRR0p/un/5nrJilZRZFVAdafFnL7qn95t5UMEf43bRJz4O2pa2nb/hAbpmvzKII
S1NhxCl+0mdW7rlkSLM196WBgzNF++x/WR/3mMOzsZF+rUEhZmZvuVFFx5af1Zqc
PyQDO/+dM3PmYzFQ1kGLDqp5ZYPBppFCVWppgvzqS4WOHfmQ949j3UxTRJH6vart
pYCv2VLtFJHrtZqV1+9Xb6eA+DI+pVEzVXfllNF4jxAP920cNRQ7+HYB5i3SU0HH
GUvTVfeHeNIUCNcqn34O+9loa/SUC4wyM5BVnJAQ7LLjb9h2sC7HZGvRxckXwizA
d4Vy85ZW6+53HcJo0qIDCbz+94Ys63bZbB/9ul35f6KawX36RX0AXED/zhQNv+Oy
b+1pvOn3OwrbWRy4SwRulZFLQB5pE4wrdQE9y6rcnIWYb2wvXcPXPAsGB+IwZvOf
zxQp5HvcPmW6Z2hGvehRDlyInbKuFr+HzOjfG33X3n8b7gnaRkQ5hMP3Yb0msGx1
fblbU3VZlFuHaiEDBQp4/ySJsqfoaVwdnJUSh5KB7+YPDg826KXlilGBrGEqm9aZ
zN09J8ls4dECy3pj3EQVRXVijWZhA7sy4dcYupVJEt/zbd2F6KapNvQuRT3ESqJ1
MMcafS0F+MW52ZM4WNHL8gj99n6tGux2NxiodOsoBnmXjNy/q2CwILEnK65wZ4Lz
z/GAA4n4oSESsV08mDZgB/KH17MHB/KL8uJsvOc1gWN4XwoK4s6YaolTEf64Lwlx
6FOFPv0fLQN+c7k7LmLTOLVKzeuLlzIGdaaYDs9uqSlyP60HGNcEh+SkcxWCrBor
MBR/U851c01ZWW/9/1wk5k9pyCC0sEyaiplKDGPYXBfWsoyn2gkTPFiL7f+ZhwAi
wq0irylIY0IwwNBXx2rZjrTRJjiNrgAU7Mg4Ujg/5vQ=
`pragma protect end_protected
