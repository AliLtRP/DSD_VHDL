// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:35:28 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
MSxb6OxyUnML+MuYdhpFddA9W81H6oTc5Ib29/p4i5nRxA9DccuVTIwa1uzUwxW+
01r4q71Lv0Scxa6dWXVSFaD48xJPid6YrS1j3Ga5eWSyo52nvKlP1E7PFV5Wc7hT
QJcCRbmUl1FuBUK1MYbp0joejjLjwN0m1pR2Rlw5gFw=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 19360)
tNfMmjFECUWWAzIP1vnj9mGWxGZYomToTP6+k3+A2HPkgtyF20+78TXYmoSJRxxe
wq67Qt9kPTfd5fIpHmHKusxX9xKhaVX15605SJbd2EAWqy0Xuj3DTEOw4Z0lDV9m
F/486aBgxRQEa6YQ/STgo+DJJvtY3AtT8N+sNQgbNWHJlkH7dn4ph4oezdVlYoQS
kP0tw8Pe2zczRiZC8mCSPh4L2dHKQbSAy1R0vGWBWwtIzcx6a/nVTRVcc2glhrrY
y/dwfPsEWjLqMH3keRAw7VqQYc5Jfk9Ye9pmG67l6+eUR79dTRgrIQcirZzdNKUu
vpeM2YppFZgtWnUJXG/8XC8KkZp0beo9EvK7Vnnql3y52MNe6/LNFtEk5CyUsPGR
srhS1sclWJN7Vr7nep9D9PEBC2xx5Cft8QLXXnIXPi135lmp3dIIYCuebIA4970s
s81PlGoeBPyvQxUU1FMLkAjOi/4IiLisDo137O3I+wHX3RaiIXt9YzsiV1co9CRO
3rgp3YKQVp+5oCcedvRRdPumn8blCddtEJBkRy0fSeqGMd08D8G7XJxt70UZ9np6
ScquuQNqMIOTViMoHvLzs9ldPs2sVi59L7UJN7lkbOpYPwqxEIQ3po2fDhZ/o4u9
3wjjbxA5qncFxm4H5bTQkqq8y5U9vMLd04bS/MHT06I7t1pdLGo5rMR5TAgdkQyL
vGgrKhfg8f/0Jkk/Ueuz8GgHCNFVmymY/wr8b+Bty4fLpEawGIr6qmrb+SMdR9+0
Vki409euyihjuqg2vj6xiMJsGm3mIWQo6sQ6amTEtvymgni623WgMkrgsjv+XszL
NzZkc6NSMzJXebv6qvpSWkmkNd1uLXqPO4OCfMyytFBF7o9gP9BwFk0bfD+mYVj/
VpxyFeInWWECTgvNMeGr6IWaRxeIMFWs+cGKCNsbNyCCE/EBVNmRjlE0dOVyohRn
3zxiDPy/LO8PAcvRKXIVXHJRpvpaz4qT+3w/Evt4Y46BrMEwAvDPfipg6r6kyBqG
3DhFxdwTY8Obteq26Z1rmwp7FSfrcE9db4p3kx3NtHlz6K63j+p94DBJ/Cno49m+
tWc9vpauIa30o5iR68rzF50lGgfJyKN2sSv/2LOXZNYLBNEigaoRC8mC624Qa/cC
3ts+CKigcGqhLInIj9x+XCkQSi6D5DmH6Za3VFxDvupjXQDcX92k32h906iZLHF7
6uEh4SGANvtfrbV3IAOM2TW1cswpcWbaB3uZ4F2SyOT7vNvV6CDsbmIlkrmf+xLN
5T7IRGnBt6ERbkhxwvpELRGkuZLsrlbPgw65/kQ8oVFmROAIcmdb2pzHuXMGed95
s5GWoWyTSKNcyVTogshnJP82C0eC/YBU5KpcMyFiSdgfyJABI3mOiR5yogg89R7W
Jy/93H5UBRCFGFgesL2rX5elCEsP+Viyoje4EaprP/1nA3RqO1oxNbQih7VkEXn/
NOBZUa7+h28L6j9BfyiKH2Cg6rKuN/ZHtmtTgonXx7vac5ayIO6jaTshvo4p9mEg
Gyfhhbs7gyOZw9rL2SHWLYjq5cusboS7I3Q4gg9eSJtyEJ18J6g/q0KsG82wVGnN
VUgWXPpdJXZGXk3pw/ZoBIacAY7GBRr2ImDxix8yFSWb7eV8Iud1xqI94FSjMCYd
wUsLDAuF4H3IoJNUuow8mZyHeUv8CaTaW84/GB3pMevk9ir4zkMDro8O4MZ8mAK4
ZSPyRjmF5AyAUJy7L5/bCE6WZNxzad2YW6JnvRMQfPAc1VqaxhN3PU1Jk/evcdOT
qPzM55T645saLMx9dI92vVtN1e9X+TqFuX1M4Qi2SCQOy2yClIwNUVkOLqlaFe80
iSjTr1ZtRhlCWRg0vXy+Xys9PZCUH7V+lL14Yyt6o5sYv13kDwj4XuEE3XT+ZeJG
c4A6+tucerdwLnW7DBlTVTx0ieoPzZos3dzClg7DLu8KWTSr9oQNcd4l7P3XBvWs
q0V+jm9tmcDDUPIOvxlbinpQyeGPWz6U53tglD7GkU7EGQGn0bxGUfAuUSpWZvOn
JAencN/igExuH0p3OpqgEqctllvL23y5BajUymqRQuueQ1hx066euBq0Z11UwYCK
twIBCcF/lWlrmmSwZN5IvEs15UHPhUfKHamltmDfShjJ36EoWmVzl8hIZ6QK2gWm
TKsyC5i7wneN3RRoaJQg2Vs4d0jE2WjXjBxTeygdFZfBYQZM2U0TKqgNSmkFO6ei
GqA/FuEyuw5tO/SoPGeDffSoHFnjmf7MJoDPLJGN2x8AFU63UaYEIGReFc6KMaPW
ybFbJMJbW+VuIvQal9EId0f8k2GC7APIl20DWpipNl0LQc5UhsHY85MHmrmTamDF
9WCLcE5QmscPevcGEtKLQHwsWR1amNX1okl8WUTIBM6hx62kbzO0T2/2jW8wDUNW
6piwKffWhTmME5ADISKt/lh+2RPh2SeJqvH1GWqladuy2SkkSJD4Seosn6xNyscB
AeN07Eqa6OB+j4MNAGO075jiah2yNsICXgb3qbQvHXPZdA9L6G8r/XR/LzWODRXA
f4lg5EQRBhxkiEyh68N4BueAx4uxyCQ4cEcAnamep7qR/rAzFfxO61oJBWMRgWxD
SC7V+RoQ411r+cBh80IgPByUTCZZCmH77jy6fGH85yQ6QvbA8x2tKu0hv6Em3JqD
8lOEd+Mrjje3AbbT5fHYIE23gDOBo91KiYwFibd3SZ3bw0oypSS89hrTo12VEudK
uRjT9TYEjtrUbJNv3z1or7Q6DGvAjABUbS6n7/j9Fgt3iBxNngZ5s272L61d43eP
t4ZHKQk9h9kHEW6dOw/DmcgGIS+q1UgfL+BiZKryHqEllYPgRaRpvwjxVk2vrVRJ
W5p7Au2LnQDOdUI8LUHHVt1spHJux3VmyZnaZhfpzKtJrvc6HeCL5Jyvuns9YWoX
oEgoH9fJjozxezK6ofH1i4VgvT4Uz2wUEiAEFyHtSLZ9oH7VbcE+0aY6bIbolUOd
xcUwkkKDXnXaVjRKcnPf98I6yHSGFbx48zgcMCzC0yfkoHYBgwKR6MxyehhVILKw
3yr+7eSveVKlokTO638LI4EHHfYV5A9Z9QNCSyqwNVkRpye9u2/1BFd2th4CH9c2
gCati5N7KoLXKb/iBJT7CZps3HdexNQ8MAUx4mRTo8Fne/9IMmUW2GXiUOuSvmd6
lEIheZqXNac8bjEQ73sJONAmTMuOddkk8IFYlH1ob2qirmkzxfHY8NwiY9PDvs0B
3FcKSCE5xQ4D/my5+sgS+lejxjvHe0LWPAk/cuAQaMYSfimUdezmHRks8m12zPnf
J9byboBELnoeEpwUOrS/sKgzWPWyyTxnpjXrUSfdRf55xJGFcwIRHi4Kr5gOMarv
AYZ26v6maiFGT23FjGSJi4TroOrNSCb7GPdkn4HzLoOGLVwVY2LXkiLl4JmQIl/B
nkZVeSuqxwOPmwsZF9PoP2Sx5JjC5VIEt9iPDBkJQegi/x3xS+lr1m9GQQ12K44a
+L3+7w9IqIWebEEyVRyH/RKP1qw0+jwVpzkUhgHz0R9phFw3ZqBJ97vBoPwD6F2q
grX0TaPxVi/N/oWb9pNJqsWfPUw80woxpjWGHIGuG4LhyyoMVuP2XtPyjUDC7Vaq
1MEIE4ItJVsO+0X0g2ZuzczMy4d/cQJr+LvFqJS5RFEFPpNyHEB4xSlKdBpVHcq9
CgqZsk9hPVnmRDgNCrw7i3YPhqpOE/Zj0Yk72AisIzmcKOu0xXEUBrJ9fRuO9oJ8
5ofv3G2LGM/fIswJ0F4tNGQqd4d/0kYA+GmVYANjhl+G+Ipxqsbf7YF4adMXfGk6
jK29TdjpOF7opMJbx6hurNh8IrGjhJcqk8MA7HG11HzIjLUzGBz/T8e5C5EQwOqk
H1Nkg27w7Xh6SlgFgwL5sew4G+PqcX61UlOFebCZHyoikj58w378R7v2859Ngroy
loMz6Zp+gDX6sJ5WHuAC7iyxDghmUFpbzG4vrHcMzbSBHdNXJwf+u2RLASAg9WmE
rQAhHp7ujO64wiUsWS0oihoZuMx7WG0dF2sAh+g2PQQEwJL6JdM1OObJ9ApBL1kf
5rJ7OyJVtU1lMQV40VC+M+cgR7ti0fuvBRLSdinN+TZYCtxDevb4YR1dRYJaBYkq
Scm2Du5PyZy4QJ+xTAVELAqylDowMRdUmtxqKD3zyiesgT2rAtzpOGJmNt3+jk91
czk6oPDxlFd3/XW6osIgq2oZJc3oZBDlGnWUXMAgPvQz3C/RxdKXt8+NyadFf4Q4
HGiegOcOQOm5QO4RilRZ3fL7/5ryaKuJTL7/DKq+6riIJPgaW6AIX4eeLYiIxG5f
B1xSpWPCEzJn5tkc/Tm03SlXybEKKmVl4yAvBeChed4auEyCrI2IVxd5ixZpo/Cv
KI8f+6LmQAnmt8uQ0YLUsu7kIJQoknjksblzoHbd537Ik3AmH2UozY1KR906aACS
e9oVgb2tdXJUJSfDMoPR0UyQB6qpwZH/6wlbau8lH0FR+R44rwne2bru6EofN6s0
N+Kgb04uaQdGbJT2FGJBX1lkcNQrO8XPG2oWqU82cOdo/pf7hsH9RKsjwgIFgdHx
Ea2oPsgZSCoZ4w8Deo+6dlnXW/LlVjcoAXFqoIn0Jlotq56Rz9h1L3H/JBop5egZ
Hamm7BxT+VrU40zp2nQRwBuHJ+CRc82IuVUB8vLXLJlKIFAqAZFB02L6kK1HY7Ep
3pHb1LdpYWz7tYzKDCRnbDHNbMNmrmOA/mGlcfI3FnZj9tHIh2pLPM+bnaePMtfA
BWH2wNeUHixblWjbSyh0N7gAwcigwBsnkUzeQskm0Ij8t+1sQHUSN0tr67ULysdx
/vI2mkP1BXSDOAxlYbWomcI2MIbYDFN7ZQE82ZpIS9zleUwfjazclKG67yl88Dik
0hxMUquL8imglLhn8Ojyg7x/ElzXb6Xfkd7EE1Aer2STeRZV7ZRb3+RQuao0RHZY
TRtljBgRo1mnTg+MIbV/vFzz6tLiDWekpb+HVhqT7w3OC6pyMTvqJnjBOjvtILtU
aVI37jGM2qVyjng8aWIUBBPqW0NyyRsI4kB5l252yazOQFag8ihDQOMObEzOLkuw
3S1TxFrR/zTu6xfVEFaaW4AnPrIrjL3dSey69NF7TCwLtJxCoawaMcnC0lt8nhWI
X9BIDby4FU98T4R3U2+W8zrfCHOEsdhPdWZ7HhCJsy8QfeNozMuxry+rKuDi+RVv
PAi7DBz9ZbuDr1N9iogyePEARafs/xnXokfx8uO7t6/jTMEQqOQk1ovtaX80cHw8
ru5fogmen5grbCMFpi/4uWPp8hMhk9vO8cUxOJVls+A756yf2mOvPSXbCdUKGBq0
6lrtoIBjAX7tGZhuMppOkRz40ObL4xpZrm87yi4zDF3kKCF0P0fzKnqr8tR+JUFP
EiFHSQBMwT6hOg5dLEEv53ESny4d0hKPfCjzvnVd1LdYZuUlKIJC3SI1tm0HMVRQ
IQDzVgFNS5lE0IvFDc0Goktl1Ur8X+BUCvKs3bP3C57TDZNtA/uBVTT1fCVkXoqV
FxqNvao1Lm+ybRoxsMDd1uP9BBgsRPq73sx0wQs4PvMW92KCdqG/vHEr1TKZ3GCs
vcShMEy+Zh2cMY/dpfwbuTlTVbmXHdR/FiIWOpzR0dMsRCXFkPTM/89qqyFdJsx7
6f/nK8pS4+ALR8ZHkqfBa0Lltfmo8vdvHEMzAfXkIZz5IzUaKeIaSlfR6uLXekih
rssXEezGv9T1ooLx4uK53FaLZQ3lZXDR0sxKQHCTszI2/BxltvLA6GmUzPNl8VFe
V30R6ahO3Ln1/yG50JJXLmvmmGUFDUyuoybzQt7m4eUN6g33o5IHbeT+tKSyXG6D
h97ixCqVuOjOdqZnWzOa8Dw4ahxuzYVTQ+2f7cgyqQMxphJ6WkcE4K1lZCmWFLPm
N6/l9QTQ86QFhp9PUwGuluQkEPxYvSPpwYsm5jlssyNwFEqO6jtDOEr127KY6sjI
7uFZh1v0aPmj6BhImqlYjUmDqg11Alw0YlD/BkDaTf0E5MpBsot4QBhCv0re2/8n
L7Asr7MXJhvi2H6pddEStr1YmgiyWoOBFOCZbRhv9InMP9W8iu9xb1iyvNNG36f/
ciRX583axDwwhtcAbdOhB8XssdAD02EFGXsDNzcEgAWb3Ft4ExWwJldCM8OIca5b
q1QmAKBFMJmpOWDlc895SIWnppNyn+FIueoy5Z+uo8qMizvgLcY4/zuAcVsh6cfH
gC4S9StQSSJv2fElIANVE9xiVOeGjdEa/ZFWTQmDf51fcnbcwBPpjPt7nM2vglK5
tYa7i8R8Nu9qXH++/vePyxRvRRag919MSY68fVfMPWO6ELQfac0yaphrW91m7HjZ
DQQ6Bsx1kAj5TxkBWr45mgiROIwZxLZx09flKSmGe5SuYF/u29DHx5Wx94mnakr3
JTCmWRPxjEV6f9FPhpSgzET4drZXED7gYwCa4BLMXIMpLNRU2ttqvebuzrJGyWli
sORWfdNCck121/vjqUUqVR/9b16GjDZkpSmLf3cVva+cSjKwRDOMq6Yvz4xNvNnT
EupSQVUYKCgaQajCwflAf/ysAatRzIUhec3pIGqvAbhRxzcYidkUFIFQdqoEIpSN
RbpxKMFyDA5zY88DlHrUKiNdcQO8iGZQ05TqF6vw8n5CwY0FPjpp+CqrOxG/VtnO
izCU6CDRLRdtwyGBkHJWyghQNqf8wEnBjeCTOuaRG6W/K4zqSnwyPTKBlZ1NvEmj
ctSnrzipwLNkj3crYr5N+QL7lMzu8OAnHvk+iSIXCMc1mwfeYi/TuNo8FIKrUloX
tb1cjObNVYzi5801lknXeFAuFRNwxz7zOOxncrht0T1pyZTDg2pYalFKwyTJ6TVc
D655HyKiBM4Qf8vZ4Eus4B5Q/xJK6GUYP9N46fPK1SBu5pbIJORWHphlhF3dRtiW
60SOfj+ukTeEqoL9UkL+JghgIbns3x6Etd04uyazMjJRH5BFtasXNgtVQWsJwcJa
YiY3K5sdfYSNLSiAa8hq1UxM8loFlamaNBQy0e1NSGyD2YYv/DnzsRZbMjuzr6pf
KipwcoLSFQmg99Fkg3SAPa8E3eD1wZSC7TvE49GiyMCBjdCo8EaFwhP/s1MFxIre
CCQnn4QnFHRyk29FX9/k2iCqcVhqwOaT1g4YEy0ie/3m80udkzp/tSLGwS098p+l
Nx6GaVaOM48eA9bRQVsh6hSh1lVFmzDmre57X82x0nf6W5eMul9VnB0sQ5bMSUm+
dtIs7/o6Y/11LDpIbxG0psRDuHnN2uHxFEYimzJ50YD2glh96/833SHozZd2l1QG
jV0cTcjoF2FcvBsWAXC4/yyLLmzDTkjGnzVqURAtfc17YQPzujT8cvHQ4xJMlesY
buBnf8LC79Jv6LWKg0xfrh46mOINJHH78/n9xz1d/+mgG6XCjevyi7sFp12InQdf
dZpwtUSytRkcd7tyAxZxGz3g31pyElisEsRiGvv7ygAF1OKKq2ClH9SZAPjN64ZR
BqUQ1lvLvYwMA7NHxJlvoAjrjeAAVg6BVs5i0mE1IHYuoCs85kGjFWwZSFhzvNcu
gH4uBYSqXMcu3reU7h0alozTfpTyIhUJPm3fBeLt6PZRR/m+AjC7OEuCRckdVro2
lXfIiPJymUjMPzV8eewnv6r/ZyhmnCreNvMod8gDWi2MExz8VJ9sxL5EpsYVNNec
BimEzf3aOvK3d9e8Q6W6ni9YizCo9gv0q3aW7mkwQoOigT59f9/vDkSXZmGkm/mn
VQtnNYo6BbYnPTaQGj7NLtytvY5lwvc51tBYH3T083GxsQbvq7O0Q7GzZs/eo4e8
7fVSHdaZy3aYB7qmzLWTd/1oUT52uFig3CU83dOc8w9dzRbrTT2gRUIjLSSVikJB
Xi+ZxigntTkjS85aRksWiF44llUIQKtqjqLScPECA5FsS7Ee2Qhpb4+kuoW+wPpP
kLZxcDUXKk6Q40osB7GRcDuDcZR2cf8lsPb3DVHNlHXvXUNE0JsoQ1n5jDgDpVK0
ONd277YMsGqKXb89+vPxlMvxtCtP0jOH2brIrEPIVfuAa2aNaOseVQU+LQTMRqF1
D3v3lipvFv5L5ff0FZt5FnwdUZVBrObaEuPRsm/xDMK+kit7g42l+QU3W5Ra38bc
sWd4GL6wm9EmXrWNx4iBYJHn8/WeL0KYqOdA+XjdODXFEnRpm8gEcG1SKhGZT7Pz
e+FfmTN4OE0m3pXrtvHXck1xMbVcWTxZsfINNNc7Mx+NXDFQwX1C7tPdlxuc/D5C
F4+gcoqZFQSispOM61jnZKkcFoC2Uy628JRb9+3CLUIyj6bjgYeog3VB9RyXtYZ2
WiLoFs3Wcag/f19+8vvUZsIspnzKdln6nEZaMDxc651FxIdydYp7Hn02q15UA5+M
/UF9MIw6QGSIwtqX0eur0fD0KwsdExIMXBhL6C7dxkYlN8tRYVG1c/GxVhBjErZE
ZMGEL8QY+jZ7tzvLebioCa6ENiHGgZjOq90pFKcaOi5NbMzRmQWPlQgJGRkt7FER
KaDqUUD1I6Xnr9jKv5yYlwGf/oAsxDrYH6QIn732Ep3W0jFJ85eHyWmg8LxYaVqi
9sHqiGpgrV14yk8nzDFOGRft7qbtQvbpt2lgSI4B5ERVUpAZIhBC+rjymNoh2wqD
96Dwoa4mGUiBA18dAPfeZ8Q2Me1AbuOAzAUqS+V8VsTT5sPeLLbk03DJ5rS9sOqI
iBuA8OnrdLUdidHVXATPxR/0XlkqKpcAacWtfYEqO9xgIuquA70YCXIJfV4HpjoC
bQ0q+O1qwd3SzuPgy0YRI/E54htb9FmWuoxDvAP//8xs4XjCjJ75ANgwrDYy0HuT
SEXTAQdC1qyCGkP1NGTcaDuM2+h+aZX/zty+t65uw/TvGK/2TPjKw7RVK1J8HaHM
qGx5H+S7c0jsXQob5Bqk0b7sSZMO6BqM5tewZKr1WJ6CLpzqCkRBv2vqcOcMParQ
J5uP8jHgUrUCa0vA4hwefxPEpD9J/REbZ448HdRCsZjM2tPzRunfHkyt3I1VvTs7
VTXF4oszW2Y8SlXfzu5icat/aH7TAJ4YZ693QPF+mg2Av3f/MnD2xRiDa+qNCh+b
Ch9QFG3hXAX+gQZkcBm2wHoepqKtWLKEEBds88shyydx3i40fbUaYafBYfGZUWhm
yVSHcdW++DxMAS2VIxZhNCK+F9KY0NindgeBl5rn1yXCvq6ZBm+68jHAjzQfFYLX
aCXZ6Z8r9bAW4Un/CMh0EE8h+OoUwtX6bmkPK273dhQApuLfFA1kjKs/2av3SW7C
JuUR36Vzreo3UUx72CuxGSLmHzfxqFCmQYMTUt/W2XUW53dSri3b+bTFtygNpsS3
20h3ly4ppLtItPQDR675FpGwo/59ngcbQXefcXIn50jGt7BgSh7nUwv/mZ9E6sSl
I6XCXuYUvu/uJ6KuIPfdZlXgNvjcL9A0ZBPCAqCsYZErOSbSEVIQV5HqqSR8tpOw
rcagHGnY/b4aOi6I870wa5vOt5M5vNNnThPl+SQqlCHbSIzAKxp88hu/5j83sPxi
Lk8rupWzWK6aA8gjQrvPYUuLS0dWpn9JRqpnmBSPM+glc66qdUW/QBaUct8CGOpt
KnvNDRK0+0cHgCoX3qwsqsR67MHXgNRqPRo8OlUz4SqSyNfwyc+T3aiyX3JhwCOx
WMB7VZaDt5wGz0u55Io3fGyKdDN1buiRBSs0zsKXwjw1L/Cw2z3DRNDY4n0pnDjq
QxESZWCZIaYhF8oP2M1kmYt+Xukj+KzX0BMTsRZ+Rse0RYJa3SjpEqv4ttT1tJtv
0mrri/n5VD+h2QWyGsrrkfLQAyu6VMEBctXKE1gBGt6KWdZfnMunDevUEmO4ksW3
oCwu/OtR5ZToFoE5iWvuCvL+cLtKhCsw7ro/t/IHEO9nSNplgvMCFrM6DbP1HQgp
RZbYBnfmUyIGXuzDtpvB6lRTS6/X8Wemvy8kmAWqXV5zrw/Aff2jQRA5G7h0g2dn
6tOzEGlIsYkgO1HGFsX33FYUtRhv0Kpw2/p8424b/1wjtrvQw/HSwrp1hL9dm+BL
9Pwj63yxlKIfROF5JitwF4vZ4+jB+XCbHmJX3LModHY8robQ4OrZPxHA8ZYtMejm
X4++OsgCU40nd4l9Cprlcou7lxJBJMjLcfQm7Q7YmODZHI8G5fn/dzJGMuNbuVJA
PUfrzZ7Ts4dv9iK9vep6QWS3gzoXJP9XBG5IL2cpkU4iwSvmi/m5BRgKac1wMnVd
awQRWlE0OK9jyOFHXCcRU+ePNtyfaQ100fW1uIyiJucOQGfuR6aP5usHvZrvfSxC
nBuEj+yCO2kn1i6GACE6Ci+N3C9JIWAVwqjvLjVmeelRxiKa9ZpBxdbl6YbjvRNJ
BAKy3DU360MoVz4icgJlr/zxJTr/PqgoB64W0iXm7rs5YOZNvFX+CgP2XxdOypIy
1npx3GNpzIx8e9Dv0Tn+4SjNcnQXoKXyr5jhPPz+IOt5L0RUM57riFF2p9XccDTL
X6lGvZEf9zZzspeWRhdiYm45sp96f/xOO4sHaRzxLnkI7y95SI9cS2nOVKqOBLUv
IsOxnz8RKuf3KTl/9EMTyt5iTGgWnKogZFuhjYK4xDtC5s9vRX1yFD4PeLjfXD3g
/j8IeJHC/Ku3otYjPSR+Jh66uv0dRl9AVEaAP1CUL9wwIyZHJgBKXBUR2Jt9kqJs
kUYUeVqmifGgTX+UIS1GAJbVjGF1aGfYkyIvq11PwE2yuUNZmXuQT5Yaw4MYkzaM
Ch0cdONdrYmGKnAkxvkGXTlMaI868dKwPMCKoMJYNeuDaWlLO77GNmL44Pm87bWw
11G0dItYIQP7oDvXhTZomLvPMRmuQgylsUj5vbHu8uIHL8INtnzmsJR/H0c+HTRG
cwVqAqzATfmCtvnJMQ+A5SfN3BIkrm0EvSO2BKCEK5dNAn6JxwIvoaqcRD+16KFV
5lrC1UpqMR9Sk9GDwLl/UxT+9ChwamhcCyxV/ibPPpUQi95DmA1vNqsMQYuZQCE+
xYDj7dbluP3UQAl1gLX13RAc9xL+xPXAUNbQyp8VNX+flOGvSqsGLsk+cry5Dpve
X1cyJ2xk4KIVtToKX+hyqpGhNBfy4krjxC8KGk07rQ3gQUvtO36KeXo72CFCFal+
tKTYsdNTWkvojMTxkUhcpPLqaGQ04OnMJMplePJfNqgpxS/KgLdSwZE+MZSvvBRg
gFjWrpG3gMEX1CPPRLVYXQ9FqZLvIBhPWJpNkzGpe/fPpEt0ISYbX6JdcqnlAK2m
4306duajhkP/exCRvWEPWDK9Enx8esn4WlZ20DQFIDH7L7q/DC97CPqdDkbKncqs
Lh6woREbTQiGlG9bFIVpvkWwkFa7boqsSUVMhPXacz8zR6p1CerveR6q7JHto0d5
SxZEX83YD95bfh92uXv+7i9PB6Xd3zBzawjJLBMsrBEVtxwmhufVoqUXcWqcXeEh
UoOJxoRkiEJtPao6ylUeMEBXo89qwiybeY2IfxXERVnPENXxeN2EwU1dERnjm8Tv
RvKk/tFq9/Ktjsn7CQ0lE8aK370yq2oOX7H5X72Tfq1+cU+Pb767SF9RJJUtMBvf
ZRezsm5NUu6hxtPUv0XC0MNDfmZ6cl86pv2RRvA0wQr5R/vQuUUgc92F/Nthn2f2
UWJkyGI6nDBGtKcDlU2fwlMZcb004Fqpy8kxUubNuyPTUWw1AGmuOYvDDfjmoQw8
BTcFb/odPWE2O6Z+QIckDuLfTtW296/r51Fx7rMsdw8V3iJAxb/rU8Twji897O8f
y683IcDHWPGY1FPnjTwneiV/07Jp9vW/RIP+NAowwP+Wgah3lMc0Bu1TZ1OrrL+l
x65wdHIwdtVtAmwl5EttdJGM1WTj/XtDCn/OS9qUM2nmeGBGRLwi5T/7TSaKY26D
iWydqBXc4CxbWNcDopadzChY1hQUdG1D6+ww/AjAfLZbz9GkVAAX6wB04Cri62V3
ZC3bD08sYUDNEU0XTFrNoFYVGC1/gz6lxd2V3mKRnda+aqfDwMKw8neW73xrNVbl
E1UO8d53cXewQm1TRwkxQLS5HDPMRaRc5EVVkLcLS9aiHA1kiQRvO/xbOC6cDurt
mr5Es8EqdStnp+NDjPCklque+xBEnG0yp0P45EcZPU59pHvcRvHw6u6UVv3iFE5R
Yx2pjwCtc6fdE1vkGMsT9IoUKqM+WS0OTwB1rYeuW8IUUDL61iAFWqJlIZmnNgR1
o0JbHoPq16JBVo3TdqZVSJ1rRq3+fKdOSnsqG3fLhakAGoDHQYN0cZFQLgs2A/fY
ScVh0O8RiM04KnlSfVn9/32q/aauzXh6V6tqb2j8j3bcmbhPfnKZmZZn8TEw1A3o
cEKMV+F5qmCdASqoLP2N9c89jgVIWk6VXkK2zk/2DOSl3Vbz9VNo3S5685sngWLy
VajIRY4Vfh/6e1aZiRgR928Sb+cHR8bSb43mHC1/L73ntVczHYVelq20Q8liPwAK
SaSiztMg5a358DnhdsEv8FrA7964ouS1idiUKkVf4JSl4aGWGkz6N+DwYfl9J6/o
XDHlDWMq+p8MUUoCZ/cHoVk6/AGQje1mn/uEI88lOXRRXrFnziyjq6TT0hkUk/ed
T7VbcwMHWkkkj44ExEn2PspZeXprDxQwn1t9/I1LyvMxmfLenrBwi+N59ewyc1NX
Dzcm7c3+mLMbDrLu2tsr0EwdKJSJPyVTfzSPrbPbhNOktCr5RH0XeGFnUTSg4n+N
OndHIQeEbC2r7dGbsE/0ZBWaowtuhbcp2/Qu3TavZ/CylA2Kjyud9SbI9DOiTz/M
KQG6nu3ZMuUk7DOdw0J1jDiIY2uvpqNfuhB+0v9n+PitHYWOaYhrIQtvbO94EAmg
yUI9th1GroajA8xs54wtKvSBSG9kkAdwDz9Mo/osahnLcsAn0EYKVfucX32tTcwR
NoD/B+Sv9n0Ezf47p8yGZefOppzV1M3zuiX8fSFh14NUfDZxVA0J1B+KU4w/Xrhg
XUsTiBpeR25ZPl/aB7N/1qa88Nix6IJSaiFDBEaF8OmbO188vFjqVwzKq8YdlqFQ
4m2OiO+z+L9AGrOVNwmyYBipk5ZSLuuAcGJYDqIYKZMwdkjRkzGfEEE9ceL3AXxW
CPUuuM5e280jPjyP5m8668sjQBsZV5rO0yiYIxACJXBot0b7yI7VyEUIdnoqlEZV
J6jrvmkyz319lGv3LwRM2GzN7bzcrFEcUDjJS0kX9EWmn6nnmXCpA9CW2xcW7bUl
y5y/gWiDr/fGZ8YTlTYMbI/V0OQu6HHzpsPC/2FUkYYgS3g8+BmzeUS5iaZ1VeVL
3O0dJsHmhLv8i8YU15MD28AjvuPdfsA3D7H0GFybcmrl24p3brx2VKikhxSTdLph
mxuAdzxPeXEPgbdDLwhwVHzPO/GKg+m3QqrPMuYhwR41zfFb3YaVGqZZZDBBLhVx
xfHgBQ0Q6t/LcE1gZFsEa6NYNL46ehdk1/k8nl03pcB4yylEOzT/wk70QDP+9Bf6
JdiQx7Qz17FMXPRiU8YV1dejMRNruBxsKz05V/1+0v7kdmAW8p1sYiAkgDjHlc/W
GdFS0HtzYV79CsocpwMGcipsg+5vwQLQIfqsRITkZ7ZSK0GSpKMZl5wJ6zk+xoHD
7CiVhtgjxL4Ubb9Y0ALG4sVsTpxm7KvtjYABFycKevqfDwSVkVoQ5pZvI02tnP+3
MFLZ3zZV0MhjzgRk7s4MoBog5cwlFTw5F1L/bKuAxUZ45YevwWYhDUdXLPsHBSfN
3gIs3qFWY32O3bpoPTInbcFq12stFDk7AdnN6ME/U/RSRXkeRGIh5WDghKa/az0f
qijtOQbov2KM1Q5IJ3B5PwVNlDl3SBwebYjBJNETLxDwOT2+VQVJBfBBhETRre5m
mult64TjPbotAmIH58ywLW9eFG9EoZhAvoMzbrTW3noUPZCJyMjDJTAIDWic9Wjw
8ctdH+7Z1h83aQsXZP/0/2KqHaKR5AZWebhvv6CDZ1aaxRroslqOC1g5mgE/ArlW
6n9XYrsRhTZ38klh7x4vQRDs7ikBCe2l7O44NVQ+RdHSmsWxIamuUboOhBuRvQKl
RgtcZ/1wwj98hmZwSoNj2ZuvyKuHKv8DXBrW+N5aoZqci/bIpKR/tqmzn0aZ27Jo
/9PSEWyGDZAcrKafYrDbrB1LM8sod5REMF7lp63gEDUB8QO8IFBEqGPHk8ojQjv2
Aa0rnhAY6BrBbHhWTlUEj8v47T8QsFKx9Cv9lDI39dWxMSIUUuE/z8gOCACF8mt1
RiZaBPD1RVxCt+Px+bVeBYUNwj3iC3F95FsFQ2oHwtV6X+ZCuxvrAAtCEB5Eq9CF
ux5B8dUqvtpGhtq/GV4UjCKkM+Onl1mf2uS5/V9LCm3MwdIrexBydhUOhKAYJicS
KFOjuYzgEeMIfiJ/oAkuJQPyBdYkb4+6FPm4pGcfzC2U5EpFDHvgGxRq7bgwaM74
EypebSRldr7Oj+fXX175Z0Wy0oRb2Os6WqFYxyzOxuLvFaPjuog0dXCqolY9Gt1m
8EtUyoqliW0GcaszcKdLGc0WwjPEYKqVD43hY4lZVgCwGg/vh1lYeHaF2MZ0VoQ3
Ywt0hxrZ5TiVpoeNAyh05vlgpLwoVTs6sH+ADRy2MDr5pmb1hgBdfN4oqjatx5HW
jq9/51MGnFuuRpQ/BilgDn4FsnTaB6mclJrvwsAvCqbar8zhp6fxN2V1rCUJAskC
MM1LGeqE6SZAopKJDZ8O/XrJEGvLNdutOc8JBZHinYNSYiY+Zd/GPB103y7C0a4W
IXPWCptFK/MALrItf+4jILrVhAwx5D0nfnlyW94GYuG1fKSwzRFZtpNLB0dosbXb
17PCgKxtKOpifBFReo+Go9ipWgtzdQuvoek82WTsUpwyl52xTnzS+FCjgOZrKSPF
q2qhZPwsLeuCcKhgLSK6JzXEk8OwmKUOWhDF+RNdaod/zaM3fPhc2u8HDEHHgnc7
K0F8LOCHWmWTId/2Ihvim7kkfdZ7MiUcUCeSY5BBYvJsuBkGn9EuXy3lx3lC03fr
SiRp2h9CwB+1stdEBzec4ASnmcM11bXloTaxx7X09G5pArZvs5f4H4hk/bc6Qojt
V7JvT0cd8D/fnqTzdcccXOJhWKVErhAncTgvgr9tIC1beQPIF3H7ZlPRAAUIZDGn
kGIMqNibtQwuMS6K/yC56XJHkLq7GJRifSWjJdf+oCXtn/8DHcRxJvfIti2ZfT23
vGSY0lm2dOd6yH9Yvz6Mkxhe6Nkek7CjUscV96IOjILvSKIoab+pYo8ccgBo23OB
rcocfoBuTxLKTXEFvbjCnoHu0sYS3yfKdr1REZc6OAqM6ohrULdEY5GwUBqMvPzR
uuBWa/JZQ0NvNrrWoJMSWs8gWDgklXQjICPik/f+V1iz59OUa1g/5xCAPXBmD2Wq
bQ/Y+Yh0G2XmoWaTEccYdlU1BL+cD2Z8W2Xi+9Jo7wBY71X8iXpNAhEw6+CIzz1w
TunfqZ1Dhi+De+Lsnyppat0PMg2G4YdFeHAlISpCyAPYD3cI9Ywq/WupbFf+biY2
r4QQkyBRRl/5gvHDnPXIyC00k2QH7HVaK5VoibPh73ejjP5CQz4tHTLqDweAxfb3
mYS2WNmPHalGpN+LL27tBUM7PpsNk02h/amb/yjxYTybls2yX8lRG8YvXtXVrafV
JZ/18VU/lvyRDhCV5SjIKWwleNy9QfBIjRKOB9sx1qwCTziqZKWUh+hZz3+PYcfG
aiNRpMukx4wZ0OBtcuFvsPEfEnoIoOogelMfs8Zkesxn3FeFFl1xsVoxcre5MXVs
Oph++u/+C3e+LA8W/eptkcNvGGZx9xXsV5ah+HrBZCZ60dIzomfMbOvllnkr46NI
8a1VAYzc3PNCNrNFLthOMU8MLkVeVCLhP29+14vYoOR+WAAD7d/QOLg8rwVCSsUu
UOWrDpjJd5lUezV7JaaftulkELX7c4u1XfDOS1YVnC9P84beVZ4xzwqc2tqclzL3
sOGeZkS4XZ0ta4UWWJ4iuFN5ELLmrDi1VJOwN2h6loWBcUvoBZnsGK823fMHIgxF
eciD7sniHxqOWThSJQWIeYE5a166ozbqO39e9jXcAu+9lXh3BbiU/ZlfVJc4FuY0
HvzRe8xcgJrBycwDJS9xhhlyGlybNdbSeQGNU+eX5xUU/418BUxsEOvYZBj0YYsT
WX2V5Z0csLL04jgkiG3RbT6HJMs5MlLrOJi31YjA2432Ye6d5uwdaY+BNi3XetKi
yUosW7b52DoedAcK8iV4vnQdwnTje/2mKOAZazRYBjEhCUETpi0LpkN8iS8ERkVX
jTYvyXp7bDB08ms1DcXSmCdAHZidls+khmLAH1Xm318c+e9CGTeOvH5mIfmKOrrx
ZKcL6Jc2gqUoQ4rTIdzuzNvVeJwObeEXM/dxZM6Wc2+NVqW/YU0F1cIcYozc9egZ
8oVT/9aplT4rkWPaz1lbs/l8D/YsFoGcp58LUuMJHY7Q4VSaWS7XIgC8Q3MPLBYR
V0Nno8ITA0qKgp1UU2L4vnzJlkPOkVR+8GggBETpcjQndnDlh14M9ey6+4dHi1eP
cm+1SmeKimEhEFDVYpdoXX3MiMreoF7DTZbLLVCrpfIzUIrtpf0VLsQWC9yLfZSc
dz4ccQKc8/TSuzzydjtwU+mpPetVRl/A8rsFrbk14iTIic5tuuwxGw6qJaiLoujJ
3EiT08QD8FNpWlJwNW8CV27lfc3RsHBrc92YMY62e2a8Y3507vjFQ12IS8yvLgLB
iXTfcaFYSiFU+W3N4SBoN0iWvb5KUaaKLhcpNUfXbiyIdS0yHIubQjxFW/XW7C3+
xsZpinRUCJpa14Qym7LYLq71//J0DMPe03FRiz+MARtZFpfiG3dG7Ynu4JnGZysZ
k4cc5tMmD0EqWuPLiK3hre8rc6SGHBM5dZE6LjHAwqPLWWuZ/ZKNUDOWxcYo0pAi
bmN3jw2m2+XEUwnn4HVvRrlMMlxuxSAmjpscWLQuqPUFAWJIRop0HqgQPCl87k8U
17qGBEXndCq7VqGexqoougitfElGPzyfWRlSzNUN5CqFPACA3ST0Fod4z4hUHPcl
7D6ungCwK7EKTVUJEz+GDmwCve/X/mm8MdcmLr04rRHsQmTXI5TICl3Y2slODGjy
izzKhn9eiy+x4WiJYy0t8Z2GpWQRFWgA4cCD0b9BoX/EV99Y1eiJZmcXCBnk1Mqt
gMpwf2A6cvYC77PRFYLVJNUxel9YSXIWumw4El0/GL5vxnR7fanK5vZeKF3S8G6y
EarqNfgbDN13aj7rBQK7tC0Mums4HisA68rMuoe3zRBjtWyPPh88gssXlLu5WSu+
M7SXmvdXf3lhC0lzIl5ekPRThCXgp8j/2k1l5IEna8+OK0icigzjCoYc+uJKm5n0
4L9/nHrUMsiyJx4jfZUnkJX3sZXwPUWaO6xHkOMogZFSpPHu0lxuAKPQFQnlp84u
+2PjuRnPRuvYNTa78g+iuU0M99Z8AhlYRIuwp1S5QyO6FtYmAUGal+k2jTGQkWMF
429yPFyPiZwqT/VwWoGiYgbNBpK0XLyKD4Fe30i+p4UCT0Jrr9OKRd2NMcY1jUlR
Yjy1zZumuNDnyQvTl3a2m2xY+z1bSYzVoqZGIQUC5S0yxrEk0dRbvLFcP3OHYM/R
V2O1SREpuX2SocsmwCuCM5Cp4U8tC1GTkwhk/QOWod3CbLS2P4auNxP26ws6Dx83
5/cPUEI6LW4rMj7b4zp17Db7DsHB5JFZOnwzYOUl1PFpcaXg5X3O1FMaUTm/FF0Q
PPq/ZZbjJz3Obot3R5jYvYQAngLzbN+Pa3Xwlg5WjglmGLduJiFd5tX5POM/hLvF
b0PfgMTcVXnrg18SxTQZb60rQrpB1Em5RQGJPV6Kh7c7aRz1fh+5KXIrM1WVWfvM
w8lZG4UAO4N73OMnfpt9U9bvgF5pAMsmcvmXvgcK5O21IxQnFy7lN4AONiXAFBwr
MrBGZXPEXCQTGYR0dYjVecIA7rW7RsZ3pfkK7fQdtwZl1+3a37QEDA3Fo0CZib6D
i9a4XycYguhf29brMBzdSZnUzCR8a0rJyctCh4hp+XU6MSnPlUdKBZ+xsbU1v1lL
//OJf9XzCkrL8DVKYI9LhiX5T1QBb2J7/DEbR+ktHWOAkrGFh5oiLBL5APQetu7q
2RaIdKm+BbNzeNcEEzgaVtP9iiq+I/pEhDmPBD/4hgva3ox2Az91alE40vzdsVrZ
Qqa6bpZXz0WRiGsy4e3zDGfl2+bEPqz8MPeMwbmvjutyLI0nwXZ7cL+GkeKFP1GP
8VuHt+Ymtoni5fmosYQ011XyqcljpPcKCQsahHDDt6B73K22R1b/JZDIx9EBSghH
1y5ThDWgHs97w3Y3Fz+61OBIHujWJZs9LAT5xolYxiPYo4s4i3oJYshEBp5NkR6i
2Ite0BxzwXqtwiIxx6O0WZtq55DYA8srDlDw6z51lYORe/cTOrVzbvgIcdL9tAZy
oiiI8XO8uvi2Yqmi6ffexcWI96Bu79GJMkBhcV1f7lFv0tUwn3yEaIxixYvF6SNP
RiXJgZoMYvSWzqX0P4fxxrV8EikcgY89BoPomduyr/yPAeoCuGXVqmktokeIhczJ
BvqK2RSa0qnIRuo5I7vIpdV62JwRq6lKIRB8jvAQX0NcIea1cpZlIuxMejQ6QOAZ
F68o+uM/hOgeS83s6tV9Azkedq3n8UPZW1a006qubEBn+x82wHJomqkHwluc8Rgf
C4n5lJyKSZwIskqXmPPOiW4cM9AQmit6pFnJq94UldCkR+lgBXKXUI11oTvTCPnF
OEVxzRBARYiKROpM6vQZht96A4hgvEGv/NDaA+gdLhy2n1Je+LXb1N3o9+t8XQJP
xw09lx45e8BZBAT10YvpzabsBGhkWB8eRL5/0qk/ZVPYKD9KeyJnfsDdD1fddl7/
iWodTLU5w0pTiIv3XM+Q6nQzyWgUOxJFv1v2ciIqhpNZMiQYxKIX99/s7lheRvYk
h/oMRgFl2gqx7j3b+g1QYTleDMYE1JRZL/elVXgaoLCLE+BXYrNemK3hWhTf6Kn9
ruswRNPds5YqbO02F3WnZgsBu0b546ilfS19gP5nQrq6B+VeFkrZsAZQ2Os1V1Sy
XAFq4GlaYbG5npPsUVNE6oi2wAfIeFIwLzsCxcmYTLc25blIaj9sc9nIYaEN+eAA
OGlcSWphBeqeQnjDheufaXaiv4LxRi4j3QdI9bjgusnQIN1U/MoZ5rcGTHaqFruL
9kZNBuxlSMd6WIfzYns2XilOYOHVV0/P2VUyL6g5neHWDBu82OzTInuvKyTw39mG
wOjbWRdXPlIzgw4vXV1u99NFwrEZkjv4KYGHsLcImzOb8j1mlQrkZzADoty1PlBS
sR9OlNu5gqhLUPV9D2l24CVSWxcN9GvTo5FcS/al2BMRUDL75TczG03ILKW2kjvN
aIyFNjevHyFPhidXCUYn0TIkTg1f1wWoY7NRa2hUp3kL2On9xHluRa4uS/HtJsCD
npm7/OV154oIWXu09Unxl/dDQ6jzp6omyfmrM17J5wvPBf2FzVJiWCWaT5E0trYd
FTBxNQlSwmrSdB7YwpcrK6R1BELZy2C+ejyRMGVIfLMcX+KrG1g9PyrmWO4txZmb
G5RGedrsx0jpRAAb+kpYH0fjeMo03VJDPpBZmohv/KMPGQjTZO9s5zahvvuYdSc2
Jd/PbBDKOzxwkYOzp/Z793MqYCYylXiVliyPnWYRMSQzXRJ/u8o1uK3m35WPVm7B
B1VnZ1K216MBEnM9SsHGLabj+iQ5pahGdJqi+Xjnd/0nLFbqwwSciQLRkJnhFdSr
qRIs4ciFCLyynk7YbhgnrNX28D8AA3vwMsaEFWp4KyhYbQvZ1ZL7ByLOYB8wGFPt
JkcnOg80sg8+swg6FllVvPaf0OR4+tkVbjh52TKVWgeBMtiyRDxoq56hPlhwG6w/
bkfTajJk+TCPkfsOSfDdi16x80ZiuWvijz1Rr7cT19dXw4OUdV+YJmcvD6PPRJB8
nMes/7nvELKvYMNnGEYwrCgLKFDUfTAen4S2kqMiPQv/LiPzUOEbVAOF2QMahCE+
cyFPwEVOCjZvKC26ChqfEj1sKYm1dVZgYAyqJVjwwSA/NY+J/PdMqW0ouyR2+np4
c3+qVJeESkiMCdcEhu5rdRHCQjawpA9pDwvL2pAJsJo2lCctCW76N0RbRsBMFaC/
qMC8NwtAgnZoKRjOea1qH6kPWB2PrY6DLov7U8nUX23nKwoHuHRVOppu4Iixpd4T
R1eUW+O9nuRRdyhMM6ecgExm3niPFZjqZfE2KCPNyCKWn7hGsgHDd++fKybAnI0X
c8opxAnODBFxOazoYUIqgJ6WZb2UvFD7AoJWl6i7v84xQ0qq6x1A6VyJZ50yk16M
9YKhVYmVt8zKQxJB8XuYGob2Nc5OG9vGn4M/6cHkpM/DNxLz90rkCDQL07nGw8/5
ceARQgHlh5XfX8P5Au8Ll2JXTovHYzXNr/s1z55rviXK6Si90wYbBE4Qj/ETg9h1
qQjZyJmFcoHm/WNs3DRikiwClgzo9gylJMI+7m+wFnWDSeAKEFN2RgkrughFysJh
W7gU4LGvSfRJzK1ovzlLcOw+dcj5bMcWcJYNCm3LACtxl5e9Tqq4T78remnuKEqa
RKY+1K8VhqaEfwWUtnqn4iB1Pfh/xh/wawpP7Fi+Q5LcjwNgVs67ZHJ2t5gqfJMn
VXKpJxdAZuWcin/XhcdFChKiA6swHxSGwGV8k3Qo1jJesVhEf9oalaBtVBlP5sAA
EGmfLvf1typ3nVdWNh4IIE/RLDzFPRZT+Ds2mUyajo+l/2Sg9lOryataAX0vNU5o
bRJGyaSshh/HQNBYsT9pBiNpAf2d59IBIXsq1nqP9AJMqlM3kvTtnhSuXHBLjYdx
q/gn3LLYIIDkXIniUBywTjBVUWSmUiyA8cgBfR0u6yyIxwJuyBs9ioVrvdwi+YOe
En2aJqINNvsvh7fOszWO898LsQejkV6VPnrTH8fh6i6SWmw5GxHNbtLhqsIf0fI0
nLNnSG755thtXILtwWPlBWx6QHv+SPfQCcCP8IzvvQsavHjgv9AcI5iECPScFyAB
HpoTp6b/zmQvo3zK5+X+Hl6Btb4kphl0H13H78okg6FLJQxWGpMKJw2qkNUNPOZx
GKpDiD2EgqeK3Yytxd1vObUQMMZdMYZApExODkvirtnN3PAVtJC/1ZVPgK6J/2tn
QcZJlgDjJ7/BL0/4RfXetZRZZZzP5tVx1L4fnQAv3OGfk9Z3nontLiY2pqyuM6EB
I3d+XZJcfOJC7grJ6+9KVVHcHDCV+utxy322Mfx2l3KUEWMH0FW696jLFhKZ5iLq
c73x3luuwWGLBd+OSJVJp+EFbkhPXx9TiucaXWSgJ8OeTPtOU5v193TVuOz5Ni3X
PnfCIZYj+wlf87hhHRBz8iRPz3hM6uQlqB6CaTzTYe4hRUyaO7hWMPkY6psclTVH
aav1HqbBAPsexJ5bxfR1eSe4KyDZilBCJF4eWU5fl5NgEkX1qCcgosASprRUiOsZ
xy8x/kIwmAbSVBgaB/bTKSw09CZ9IXgIMWS9WDaB+4W6CbnW4X0Ta8rdH7z49aag
V7l8pZ0NJ9N34tbXPbAOHF0LFVkiymmPbJc9PQ7Eb7/Hn7F5nTSAAId2MbGEWFZ4
VgEdEhQLk4PPZYsSsS/TN3lMd0/pIc8xJJoqUEE3n5YHyy7P1h1OoR4IHgmBzFpn
sUwTlL8qM9Cw/CbC16Ol4Is37piJzm43tOqBnsgHDzItgH2Na3kvmmo1mUPM1B2x
r41pZjp7fXHar/t8IYVhlItlMDoAV0s0xImnJLsr3OA44Impk/ivjK2n+0sfcqYr
p5ws9K/x5QSkes8BdA50AMDmYXctEHdojUAFVjwWnN+ZDOlmdj3DL70DfJK2zrgM
eWrRD4/OuSICq4JACATT2gnFEk2gmbVCT3j5J4lSmUsVKI8j8Z2vqzBtQgW5WELs
V10RaSWMz3ylPQenGByZtozuYAwdzaOpysThxZFINTBR/sRNzlQNpSRUS1Z08oJV
fbsFf9DQ138Q0HRAZGfbaW5lf6go4xZzRrIvLMvXQPbcvihX1ZhTOg/EOvfBklzd
z91GUkaSBv9E5dTMSXs72367gAvFDk5f8od3+4cyb7nXNjG0BNiMCRTH51m6Y6JP
zCLnySriGMnxK6ECmlZEWJ64t8U8Bkx6Tpj9mM47hbTbjU5KVA3Yn3Smycr7Vens
Ob43Ntw49Z3mu4vk+99nL7gjnTVFzOPs0+o4kEp2M7Zpnolgopg93UinhfXvxy0+
CF9gdmd6ijaF7YuO++Jh00DHNmY6vIlmueVeGKKxOvRad7RSsLnsy1FFskBEzOtN
p/W09ggSxYMCm4vcMcr2fcnt/WdJVyJfE0QXyq6tZ6JiikBgbrjDLjDiP5KuQsJP
h1LKtMOHROIm4JqrK8ijfYb9aG32HqM2M7++181ZEOpSJPOWQm/EvI7N32VjD0In
akJIY1tQVundgN3RVCLfAL85XuWKZN9yte0IEvJCzH2WJHQ4kZgWLw3mCz+UUiQj
Ks715FjgWIp1dVQNXc5ak92todmHrI7Z68LEdo14h5bSjGw4SqgrO+HF8rHM+y6u
13xobcBeX73GaiD/jC165SzHrgHkUBqYPNkuyCrMRlkVYnotAlbpPWQhDdCz8cqn
s6eAY1yQMLKkCp3LjNNqIPPEdbk9843a7WYFVTyS0AVq8DFtiMVqp6bwAowGQx+C
S184NRV/+ahgRQAfYun1urxSK5mDNvG7MG70v8tNvK41zonnFagdS+Vzwt8sqNkD
t9PqKN5oo5ITJZlxoKUUIY+j/g7f+78T5rXvxdZ1gxG65kJUvwQRvs/Qs3ApzunW
yOWJi+2XR4YI9wQMKoicrEZmey0oiv2D6jPPtfCnuhz1Df9+MrLs1VvfQJbmuBnW
f5z9ti1Ri4Gb6zTgTVvh7N9ANvwsIPuT+QK9jhJ7YHZ66buxpN5Iw+eHjqA/sARM
JnbWsxdM1VHGUNYyYVataLsRBtbYsvo1mJaKsfC1w+D15X6YUc0FAqbTQEVunCNE
UWo3A3F7uKqC2iCuJJgfZmpzB+w+8zJtyBm0NuwZ7nil2LPCRM4yaMWcYbTeZmB+
TpmI4Skp1/k+0NBnkUhgZPBrSqOg4XShxNgxd7fePfwehfeGHyS6ZeUh++1r7QGP
97egToTv23P5mIyvaEAez/vdAP1jn0QfsJIwnLm7FMKPYSZRhM1M0anw9gVZMoNT
bjfWGryK0oGQMja8o6MTZYm+yds/g6aqHK7f09k+ExZV1SWY6y2ayte7VcS4Xsnk
zvvEm03Rsuc/p0V0iEw/Es57mGHHNMwiURImC0yZcfsfR/Bj13mUPgVsjbE1lGaj
veNvcxuW8jnZwaRs89d9I/USDxyexNPvF1ic3DtzI8t+OP6ouvOsogJCO7+AoSQG
mHjFuoyUXkMEtTODJcTipSqKAVpSg03MyigQEUZ4lTi7Cj9UzsTEmP4d8oOuYahN
Zz1h7K8hySuUovP59ATyQAoKbnz2Gv81JqD9L5nTBuNBavU4P8IxGg4GdxMXtpwK
SZPE40wwYsCmoRvMZrGPnyS5VVkwtjEo3miwCa19/KsJ+CtPM8NF3ooSnpOu4T8j
/mZFHS4IKESs3FtC7zhBs3juuyni4KyhigGAPSwzUR6lQ1DxMXQHBZNqrXeJFfCx
HcoS3nG1guX9FMQA23DYS9sERKZjWbLBjCid3U8DH3rKrDVFdYXHpZGes7UZ0jPb
xfENHemanWswlhkh+CaOj3U28sfOCmgkETEhZ4LgDc87MOctVWzil2Yns70qk73F
nNzjE42+VK36vexLtdXHSGFRN4zH1IkQciFXR9VPCz9KDdgiSuTlEFA22rUQSH1K
TNanl2QjeqRXiy2U3YG+jNh/R7iS1vPGNEHvyRfSsUMBKMDCAsCCEZTVlxw1cTzA
MfdmgDxa6ZXq+q/1Ysx40dH8Gu3VQAS7lnhu5ijCIV5ehVH2Yu2sIm1SJOuEN6hk
zHyjzAymxhLLXU1dt572nP1Zf4wkQWS0VZKhr34T0utHNlL3UNAldl20SxjWCu5M
7GFRrZvp82KleEQlorrn12nrhmc+J6XaM7Io7zpE7+ATuzZlrLoC9+supnewBfwT
1Q6AgT2B91urTsUnE8QJBRltnsj/dbP05LIO3CVlMawQzC3m5cXWeJ2aZNFkf5vx
cjvMnD7D7KEiuHhij2SaP8JuJryf87QQbn+KZLx8aKlD1YikbaLrh7cuwY0zPAjh
UDOc7SLyF2lGQZvfSxuVrOqq5dLNqLdhd1BqMWReE4C+1wCx9xtK/4Sok3LLMT5D
zvEKcmMV4I3x/RDnHBTHYO4WsUgrVsUQzB6fqfmxtYu8FESX3x+sVBgjqRGh8cMT
7WImZ9frCv1We23UqeVoG1729OzAP0lCocOIz8DzKSVbIvqXGtYfT/BF/CJGszgF
A2mU8WV+YaJSWPgvHWansWden4OKTVXAP6d3wUcDTVMesbWziTNeVmziG5EC5WA1
4uTJAIoyj3zGUTf2YA6PJ+XjzHfkN4H8CoyB4f5DnWAc6VMVTh6wj+g91fk7Z02Y
cc1d0F9PAv1ozdCqDPK56o4sIh3qq/y7/HrAwpKbgbMSUGn13ZlgB7wsTlFPcqaB
k+mKI2zOtqoF8++TPSNmuw0oK8e6qaSo20lLIHjpc54MDxZMWkFnDFW0fzUTTfJJ
Mwu36IfXqQTEdl2QpSA3yx04lT82OzMQyQU0moxJawnPyIomulkNrb+IeTDOdUxY
SEBayZa8iyCPv5MYxllBdZGl6FsSKSbSkJRds0OdyC7IQf81ETJbBiDFPmq4VCUx
7c1iKtxSiPB3/BRpV1MS1rfYgRUYuISxTtyLQVLEKSOTzbNSyTsuGA1wF0Qu9tui
kYOL0iaw0Duu+U7tSASgM6hsOZUCD8UOdWwCUtqKwtmoJfQnzvxnHgA0+Fq9em0E
EBvPBOMao/tl98CBgB6k5KuaZZVukdrZnS1UzxcuQaqiqlrc+qmkU7Mwx/AO234C
nxPJU/jNSEndp97RB749uLPv0BrlOQmqYiSa/e9FTNGxpyTbksdNSc2SB3mslZUV
ErmQNuhd5h1xs+zDH2AAdAj4SkmU5gBL9zZbvvKqtHs4Na1hGCT4pzY9vr21Vs76
C8glmOBrpKGZgs9s8959Zjk2wbsrtEFHBDTldQ0eA6b28eUFFZ6H+SXl58BN37XO
n+CUnCXAd9OTemVQKQy8aHBIAKHzQnUf5veIm5vnfm4+rg+rKh03L6tXgU5C01fU
/EG9ABhstR3MVGQmJ1/HttADvLT8UEYAhAYaIFlGLXRIyp8IW4FakaanAoSFuZy/
0o8vh9z9CDbpAI9PtLHxBGl+ZbeLLaOG2QQSI9DzaQS1bXWaUI91TMkZ1UHk0pfm
0lKk6yOZNMq6t+mXpgnDNVhW0fV8B4avoqu9CWlGpXJx1/yxusQK24zN1J86N73W
q2BqueFQw9rLbSUskXItn6XbiSIOjtc8AF1A1SxU5/0vR9CtUQcBUxiERZcwzHsj
oHkQ6H+jCTrb8EyH1yKfYthzfG5/INsEsnLi4mdMK5lQgjO3bQ/5gBFn9mNJHHTX
dzd6dpTPvNipkkNMLdRsRIKts6/Mucxrw0sOQSP7dThJjFYxH1gOlyV1Nzb78G6P
RiRGeJ9RrulSShf4xblTfg==
`pragma protect end_protected
