// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:35:29 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
pBzDz+j62uhk6HotsHAaeaVSuWjpO50n14PDqOz+3HXNAFeowDSb0O3ThnncnXlL
WWfxwcVIzFLOf3icllL4OTNMYs359maozTCvcoz/5MRTDlFS03KQL/G3DnJMXdHR
96ln/mMRan9H9cHHbtrLEW1bYeJKGeGNNsK/ycRhNCE=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 10384)
YPtCXDNIpEpqU16Cw+KC10ashn+CNw8/LdP0WhKWwOGRaaOGhpNb5DVmiQJS3F+V
wNHt4qpDywxp/DBymL5CgDvMrSZ4r62mdtad+k+nInpzMB7ZeQcdF4v1N9ggk9Ij
SZVf3nxD5aktyWfns3iXy3K9LNHnt6v+Yt5Bvkp7JggqlQbouZ0T42dbKJSU78rX
nnETSS98/Ieg9WWgAEoHI0y5KUG5vpE8OClVIwh8pePy+WGQZ6pUyIvDvlzJYUBg
71BCXeAw5Olb0zctJ4fD6KcvSDPjBMlPm35zuscdkTLni/mekBWJEpxunjn6Wa+p
rwzdENfK8M9ldGXUL2+L4RHa4Wgps7trF/GBxU7/6fSmr2Ayb/IH8myEgzpVEN9i
lzXSekA/UjoRpSiNmL0+w2TLTO8ZbuxWHjJOgs3uQW6MgGidxdF49x9SL16FZs1P
jlRVkX9V7U3/xVUY0rPEYrCMfgFDZsXOlm9ctB0x0jZhdIkkEZ4v7RHoVhiYDVgz
RuuzGPbqXxXlXqxDX15D0H4gjDyXvmregnqxDkE5PN045vZXBDTSOs+bXZEY6fji
6aXQnnqLZor6mBZQ0QcqawuB207wDlQu0Vo5iBKERFXAFHW6b8x7x8alBJVEFCZp
NsejzvDcaiOEvfhoacIDqfc3sjOD3rDaJa3ZMW/Fj0ALyjr0/0JcUCKEwnGUEscF
5P4vnp8rpXEgYOtlCQu1lhr1LChPVvxiSt0mI4AqsEYCvpAd5A46gsdf25ZbRS9/
8l+YK/ikI3CD+OjnsQFBbdlaZH9v2kt1Z+NUVr8C0iCV4i+21agJ/t4sryPPKGG/
oXA2ZrrZIDlXcffcMcPSov0KpB0Z9gprJbreO9H722OTT8D0DPG8Y4AeHWVzDpAZ
a0lfrj6lVwNOlptv2121Rlz/E6pbvLfELnXVOAZMgOFBhWoXxzHod8WDhNeJ529w
E9pIQyfEfucvDvqo1v2+xj3ZTeRAnISe/mOXBKbI0rYNkenpZNrG4VmX/vDQJa5v
Une1IvZhwaD9XoDKOL0Sc19PLxZI6rfk8CBgdD4Oe0Nr+jXqb56r9g/IJnaqVYWl
qxHR1SbX8oP33MuByB59CrQX3p5NL2H8HYkL/JhFmPz4eTIbZ/jkUaNduHvyRfTz
D7nhEETXy0JepU4ceWPkjiJ96zScsQabt3rk2gwO9iT1nnuBakJM6gbfsGyBC2kX
3xQT41oRj8VIf057wjQplH5xJgtrS9xC5N9jjwzDTZBDPaTVzS/RVlEUwEbFQdVX
vccletDe3KzE7AiYlP4g85ePiDR4Vs4D9aKDjTCXoQruFGu2ejHDC0l1LpXbwm5r
Vb2q+2JF28meYKuGjEN7E0h27pirSkbNbKU4Jv28sU1X1JEeK1x1+c8Gzj9K62ND
qnQYNw35IJ6k2VZAc1RSWhU4rJsZx9QlzGzV0CyP5uXdFi3cv1YMxUiqadU1+1mE
K7HfFU5QQiF4FK3i4Ts5bZy/SkQf0xQKKMJhDZ5mFZ73ZbYRJhwFmQQOsrFzMBwU
XB411lxQzhajPdT1BQyifW4xgL6Xd+NwNh4UAHXksOztyksIt2Ev1Vlxnnue9mrG
rzONb5FCPgnEJ52Ny4vxsUnQ2QcR94QZ91naf8/qOsTHD3xqt53jmS1UGV/51Efa
JINO64CtabP3UTOlYOdb++TKMUoDHcg4CtwXAXJ4a7n3Aa+Izwdvo3zW5+4IHCuF
W1UU5bJ4hrxby6U4z8ccNU5XY1BMOII1vJ/dnts5asyMYJFVAITY7ZXwzKg/my9j
DLRmzz0p36FxFD2rHKBIB4CF5ClEyBAsZvyqXpAHE/QDY9DCobvbjyeyfpaEMV9N
up7ktEUJO3rYtZ5l+MQXDziFBA9AaoT5mkpccb+dDLUZXjYoVP/Q8ZuF08mxsUuk
auZ2zjk/R9DoJ6+PggoBLiMtxPsrYaOIp7fgXJbnkUKoQwYVf2ptREsrDCwPZbBv
vNKxE/+zbP1qHuhHPy75Vt4pCNOt9ohsVxhxAO8Dg+su4GA2qbCqCzOJW9yTGCvi
Px/0TV9Rad7SVaHRTyxs7wzYoSD2PZxpWT79b4/f7+8IJI+clpcZjraBqEP6shoZ
PUlt4/qlGQ1iw7yvmXLA7q46W7oY8A5bwYu6FXBjV3Cnlnoms65gMHaI1RCT7P5L
vKq0wfzb3M/TZayXDHRtBDDO5ZoXv9DHAUluS4M4abamR+kZ8j2mLmV/0whbDZMP
FGnIAxjBGeXchItVt3Bo8rr2KPfJaLDF+AUpHXtqBcB44F2+38VGSuevTYQRW5Yx
WWCfTyNktYm9ASyW0U+unZa6dl+7fxTGgKCwcBLKhPRjJAWppV9vg7JkO8Xu9XPY
2FgsnlQJl1rxvatk6Edgk+jUDdMTM/jvjaZR98fb3A9/6FhOE9WnUoUm7M9woMU7
OtaZCtvaiczYzevtOy399K4Y4DLW/Gdixxf1lPK87PbX/xl57M/2gAQpu0FU8oaT
yl+1ZMDkcIE7DQzxXmwfC3M0Z022/jZ/M7voKfzqf9FK2kONJLvs/JR8U8PxmLqD
PlJaxindWPU/MKroPOBocALbpStDEIG6xACUG/svAv9jOpJ3ghxv5frS8nm4SLX1
8YP7X2HmSvGVpCEinWQkA8xeVHXGt1UNNMDFqVMX9NT0uozGG9SwBAECo8bwSZ+f
NxaspJsJJMGgSEX8/w3mJPBBaQ9Ga6oiGbjENXcvxNLqcfBf0yVDgCwJgh2knKxQ
Yq9s6YwfqcroILwfJOozXA/pM3g/j0kzz/7xsgaM4iZiWiUgbJ0AD1BUwhrx9ra8
15oWH+589iSJHgJSmOnqcPB4GEoIWvK3SG9PYGgKPwWC3h01hS0n0020z9wA6vPa
L8xN/6SCZbdsNaF06uD+88ODlHsmRB5bUAjkR4X69+310M69DKO8k8KERS6vg658
Vce0G29EJ9ZirOGAd3BVRDW/p0O3PL7d22hrDQ8XnGP7h5fqg8rKX2df0XaMDa4x
P9b4ZAIzoGGRlcpDyeAT32D1BNe650+JW7ckyrlAE8z7Xez3MZspJzJHA5/94I10
1LDwzuy2uOrSauG2lqLWyrZY+m1JsHdp3I+KPMfWPEU7NcvaMN1XnBGxL+bXi8Cg
GdQQSl7mvWW2W9m+eecab2wxMmo5k0MOiqNWwYujczIjTRm8KFfGHX977NtwnwY6
4hwMju1u+I42TraAIyx7Nn0sasszISyug1yikZ83P7bYWlkqgWzdnMVUTyjeYx3l
Qd1299kyePF698kdd9tt6UKReKgqSrYUAW0kc7oAM1yampgLNbT80xx3HVV+IxwQ
iYsqrSr0OxMs2Oik0SD48eR+Xte+QPhZpuTBr8BjVoqQ9mQwYcIULzfjWHq0NTSt
9GbR2CikUtCdLrGfZCgx1VOgM/F21oQGQ8s923nOQZ2/9r5VXr9m3B3Tn6PFECo3
llwIguxbq06T08GbS3JoHCa8UXVrWaIxYjYSgUB0WXP1qNXSSxNa1AukTH5bEfIY
ZnpYFknmzhxAlhqSTXoBsokWklVd3oe5sVDlBevt+zQF1R0uD2iK8eBYFRM5xStu
OoZcEVURWt5s7WkyiraAoo9SPKm8ftpawdsJ84TviPdP8s+Mlj/VDDZidhyvU80j
AIJZYrkxCh+yM+/XAw5ROZb5EhsXX+2Aj18mxq9q2xNFa9G+eup1y3eVSjI183gg
GXj6XU6GOLc+QEhohVYgqEwwAQXRLGMcjh0SJFrY3xruEDaq+sdZwqktAgTNWMmY
Un43kTPa85Mrd00qIHqPejc4RhPoLcEh1HthfaOcsFtka3+O4CKS7lE2uwd9tjFm
31m0/je7Hi4JvXxzNpBfOoVrZcKmj/kqDVuwNs8kCihfI8L1GSfzA79URUPcXipU
Nt4ET4LaY0roaumammq2U6mgSZRAAS2C/ARRJyCgFBMrPPdIPEk/WJhsLDzCxGcG
R30PDdjjFDhSG10HaOJzQeU1MWBXooy2XNUVylqBTAn6GU+SiI4Zg7Dngarc4FJG
j8TFj5VLJovSmGJAEfFgcKLJH7rfz8vwalPejx3R0uMLCveiKhwhVaRQE44594wr
AMjO7OGzpld847LobAiRNX3fjnbFNAJCE1+S8XQyZ+RTXiXq9tO44eYbQ7ixCXAK
fvrL2Zm3huVhcZU6mheXT8Pqxkw/fYc0phoLWpYFwJYCkR4hgJiixgzTa85BCeOP
Pn1p1rqhQq20eoFlvmMzTlWWdv/jOC9G5DlvLIIEavy3v4+bZVMK+pQ1Y1LS+VyN
QMbCb5lsWvZjtS+NdM+krEC6cZPFxtOe8w+34mUvVcmp5/9qKrPJD6W61v/P7YiG
kww9pHC4gTNPprI+6r9oloOh4w2jYrPz8GAPqfSvpipBtDJ7yeXthPrt3rvmcsns
LFZbVPtQhrkwCJxbwV4J7BihU0vF8+PUWw5xVrInZdM2FkZsCgJfx+4MJ83WbTuK
NDYVOK9mr0cP4D9V0HKhTjeidBoFcB2iOm85YX7QOhOxZQc8O61Wz7Rm6pfOwa8G
PMxFcd0wBF26IpVvtO+wUaX5fMNWcOPyJawXpqmJgLOyj+UHIi0Q+goZchRa04Yj
Ji6GoUaPej+4+yaBK2LZlc6GqaF8+IwDIdrH1u3cyh+sul+agztOSk1oOg5w6w6F
kxC+RDNRB3vHsxN9gZxwuOwJOnfXeZhEQB7IHsVe5a7A+SNvdHFKRegA1U36SaBl
afBYLuu1K8NzPw8mggmNGjFULceBOWydJB2E1qloZ094tDU8+hJKEZkRn2iLNav2
KBA4cPy3oGiZYgCV1weE3B9sSkS7KxJ8dEMTrONFZaFahUL/Swk5YPg60O0zrW6N
UEv6m7WbgETikg1pz851OUh9vJklQYuTWTrW/88YvsrYtYlhAJakRO9b+ZIGXdTn
dPM0jXVdVyLa79Y99TI+OjtiSiqe4QPbcPQwAWUN/0TVAq7Ed8ojbNaMko5kTwgt
ocN6x9McaiEyC6NniN9DlBUzHj5rLdgyGtQ1m0oqKrBpak0oRmKNH+Ah5/L4ohd5
SQCGX7QeupBCxiT1cRIsS2NaTpdx1HRjEjKvaYY3InOd8VYQyySD6hoRhaYVyeEm
qAxpH/hUGopAf5G1cT4tEALPVcKnr3iLWlK9oed0u10lNhIuix2ZdM5zR+8ZmxhM
f8wEN/bvDygth1ILSLbPo6Bn2jx/jb7gTsYmjxGBf6kwd3DVpoB4fGBeLddHHdNn
/MV0qo1QkZwGnWSeMbNoG1n8kMw0UauJXBJfoTMl1GvX57KJizEKAg/yTA2qre1g
Q3LGwqz0oYIFzxxmqW7kjRmzg6DIGVBCYb5++Mxjb0gvbMfWE+tqDXSZD6TE7LsY
jphK3vk0Gu0ij3s0qQUQh12JmyOfC3oMXoGRc3bZNF3R7A0oXHfaMpku6SjeEC18
le3c3QVSP6b7hjU45saMRuFaSSNQHO5YvusaqQResBaaC+nmQpejImNa/XJPoJJ7
Vs6d4yj37dHD2Tc03h/FyF8CkzB2zhKjNBs6znZv42IT2Kl12ZA3HkVJL3aJLzyV
+teHH48Z7qQ6Y3cR0XFrKiPieo1XH2+O3dPUje52rJLt2BuaV1LxWoA0sOkuBjDh
JOBjbe3h+8tb/eN5ujP1yLYi283yCXiXEnDWDqs0TbkzsXf1hhfmxYIqgkEOg7k1
UUpRaxMsx5Az3EhgQeI4dh07YIxtsvBH0AZrPdtol/5LS+/vENJyZCFqbm9fifdg
o0rLjoMAKz78hCG5GUopfQty/w/Y73YSmrvTVWscEpZOmvVq3yD9migNaI40ttKi
ax46nBaDHBlcq/v40NkK93G+KKxkGvWG5mpA6zcIfSmeoGr5xScYtXOPAJ0fhTKV
XS9Okhud+tzavCQ+0lcxYUmY0uQeHgM1V/F53X6EB2wg354RIbF+yafLyxqZtS+o
88wFmwNJWvFTk7o5ZWla6Gb24HWgQ6YJGC3l/I4NcTyjmJDKgeK+r+4glazQq/8w
3SPmi3k/LcK4MaQvtPPvNEsavciYkASgs51y442XbqesmqhezreIUYzBnLy2pbZG
bq3OlDbg+3JNGTxZnC7Gh2uHJb7r2z0OLhyCyQCAcc1h6BJJmOg1mRyGG2xsg5ex
pDEwIcg8+M36oXVD2d7eHYKVyH584LyfLmHjvBBrnqitP517ByPZ4vT7Vwme37Yy
t4PX1xaVkinLifpR3q2ozvJHu+2gN0zMi3sc/1LQouOce5PhVlC7/LDqbmwp9pzz
Pu7KUWdfzFWw7Llbo6MPvBVE60l0QCUDdzghDMYWFW1K0O43WJ+NSwZsSdZmgYQA
hmavqtgBmwm8awmeO+uADXKLBJkU60LzeFDzdBxf+ArBFGndc1vXfhoVwQ/ysAXZ
/RQKqlxdHrYReL9Tu2RAzWzCt4vTdgewV1OJ312oFERgX++w8LkJvwUaWVi1o59h
QjCHnDC0yEFWehuAX4u0KqyWXVZqQcHDBZ9PCvklKIYQBAVL1/dymvictJndA0jM
2x2pgJbP3vhlhYaQ+zIt9AORFTIhkIcmasKxQTEU8AYQBmwgH9JBtJVQxDklcJZh
BegdfNLA7nyRttnmcHPrfX9kMr+9N9i+sBnL2VmPpVQE/gR4rjHPZXXKVL3Zjo9I
zSNOHh1n9HkTaZUkWo+JoGcnAlEgFNClMPcNgANVV0eII0il1hPLi7kSjq4h7vbo
I+DEqj1LthiWG0YRMsSD8p5Vhc3E4KQ10aqXeKbJuij0BVlUR4mr3E4HNSFX42x7
LleUmHS9WlOfgyffpc+nIyDeU0Ck6C+fAsfngzGRn4Yj32i+35Imdc8dsEjrADG7
s7zqnRS+2f+Nr/sUGaefdZIxZhkk/lX++5sNAK/biCFt8tTR/tWo/eFVeAMqbSmF
cJoP3NTM2PtPS42R8G7MyU+jwFL1dQEJePI0+bcERdQcfVyGmUoVAJpu/0Uxw6zm
l3HMe4GsMODFUciANI3nhD44eJEP+LntOaXCH9acS1Zh2SGVh56PFWpodg0XtuRq
j52B2vvXy53JUSRcsib8UCfhKRZyaRKoqqLudhHwyqndfxyNmpinHYKZ7TUU3WlZ
jV6NhQov3nLsGe0avB7U66bxr2zFHufxqfYvJaXbRKXH8xiqntGJg6YomnTcEWVI
SI/k9g3AJlrvfnmCUbu39s/7YPayQsqwlTmqbvyng552ocXa1c+Bp0TyezDjBGEL
5v9Z4CsDWm0VROfgsB3VK5x8568Qg9+WJz34MHnzut+fQhmUrXR1kO/65zIpcpR+
VFIpUkBVwzfWcLlAqlsOXBPDLjejpkAaIPzZCHFgGzb/pHkI4xapxKqJAE8GfFgE
u4Cd3l/bFWe00mOz1LAN6iyRaAp9b7P1RqoKM+GmNsFL+uP3dkekjBCTPUZakU9C
IBmxu/JKuEW7p8u7y/Gsqx5Jac3NmQ1OQz5Sf25y79hfb3G3sqUTfoXuxi3qr21Z
DU9010xJdQEtHaxSbAK8/fI97pzYvshFT71Osq6XOaG9d21WPpbQwXnGmoyWxFqm
oQcPXOlxotixL2C5AHyDftNhWM20l5awV8bKoj0Q9dPU+4tGUi9YnjBlFhKJWmqS
NJI1FeeyWGyb1WkrS2/POtqr52zM4w35Xo8namILlb5nOBJpQSSKxzyYQ0wTXtiB
nARs3VGix4OTtKANc9xlSsFrtvuqHEDdmncUgLUgFQS/HNEi+KKDAvKWiNc0y+dj
0h4d0xysBmC8GOCaYC7u5lIUIluXM+RGPwpK8cu4KjziXOsrjQzzVTlTcNl9FLzu
B3uFcPtXqxiYxDrzIzp651JnxIVyibrxwgOAyJeIN3IDpNfZ7vhIjeUzT0F1K2lP
kzJR3dQOLX5eqbA50BMXqV4fgLcCYSNSvLnun9FXZM7kUFrfCjizeTnM1JpaddoM
RUH4sV7tG4hZ5Y0TijLYdTK932Yvauyoxo+ARNgHRV0338vKzBzHRU/Ljp2j9rFM
CZBjpkL3wX+uhebEmXyLuce9DJ3LFaCDVm8h4T+1rXgqpu8i3faUvSGKmgoiVIpM
2cJYaTvKr2V60cKIn15QZn7Yj2rq9dIuIcUG3BW6rNBobuKmuQXKoy640Y0dDPBU
fUm0I2FnhhByXPUqG/k8tUZPhP65TyESJ8xBoLAEfu3ZmdqLcxRww78pTRSEjkJG
M5i8ca/gd3ky9YvCJ6xOJOCY6F2ZRHWSn40NBvUthrfICHJaB13Zde7DiEtPDgNc
uLMZmGcGrictVZIqFBToeVGhWKK5iYG9qd/aC8RmRIn31z/GvViX330qc8SW8+Ob
JsrfNNM3xBG5P0pq+WetdvLmjgJKdSdRytwugPRtHPVo0f2y2xJfnF5tvOo0flHM
uLoAdcZw0dRI4GLrx0b3vGzZ08XOR+Ldmux96HYvlp5HpPJelFUz//C2OpZi6cYQ
sgGYZ8+6oMXldfjvptvt49Nke1XkTGxwFAP2xE88wzEr2wa0xpDuOIsw3h4D5Jn6
gXqAEUWYw88I7CIzmiwlqdxOv7qfUDwh5ANh4zVT0z+CpoNiSJKGt2R3NsnHMzPT
+2MceuadxsOWYZ/s/00l9s52TY7ttcGdege5KMIq75oosJd5nD00M1ecEBaW4Y9l
sxiMRvrMhn7qa2W3+SNDQCXWhGYJOXPrWhnq4cDcFiEUXZLGMRSjtXbmVhlnFmj9
KjE2wmN1Gjspe3IxT6VLjqhJGEwGxLsDA2vvv63mTG8JK1SmEqGvMu4z5eyd9fnZ
0+oJDIXETIuxj4B0V58yKcf/Ry8HisAb7i6hrzEtfF7smcVjZkBOD7pmYG55H6GH
ZNnfxfPiNI6XGzAnlWAo4fSgnWBqK5EPM3jiX4a3VALOhlOCYi4dFA7HHUjRpnJX
8/RTCQej88glEMoL34e2QzH69znmXC/Wejh2IU3D5EeKvgRB15q+SVllPv7jXmyW
JfnH+1XuO460ILnRhTa4tBXGl9Oz+fhp84lZjaMS+NEe7qct3WG7PwuWOuG8yp59
dX/aYUNXfUDNK+jwXY6GVw5Fsx/RB5l9nF0Tux1rSX+FK5/O4cHk4qdVC4EuTMgb
TjQlVeo/C0+apvnpyra6xvIN5W/5KxxsbjMTBMxoqumOjlUEWJ62CvtE52KvcTKY
rC6wM5lvrc7tMN34SHgt+czmu1n/UDrmxjhHcf1D0CWXezVqns4bD4Cx+z5vG3SN
gHt10s6ei5+qZbGKG/v/sDeE8pHYOlFc+xadd722PRMY1U79/W4+Q8f6VV+yW+//
PsRQRwgEl453WHJfyxThE+LGjx88UVRPhkTihAGHvZiEv79fBKfR/Y6Xoh3bxJ1N
xKr6wEEVnnp8JPNpnTCVOx67t2WpyJ4DR5olgYwmuYzlGAHa66wDNO0hThltPc6Q
EZsJbNAGWjIcYc9b69QW+CjrDxVjZK4L7nozevKr3yC+QIP+NQUt4GrjnHidw6ue
XHNgDUwQ3703lAGUg4NQ0++c1EK2eB0V6Dpy+fMlwE3btiX4Cpzfk/fchCPwTgcA
62ulr9l+Cdkd5TnxBO8MSm1qKi6sosyXyoWifRRQPfU4D09G7rNEbnh+rMi5jFGS
ggdC/vcbpK1m5wH8UYw+qzQqjXnmSUN5nwCcsuua8PuWEvPwXmp0HLuvi6mF+utl
LHiWqGVwWveaf1A6jMRUwcFQv0XzVHsBfNdDgRhIpuKcDtupexAf5CAG4fC0xNmJ
Xg4C1DfJe1Suzh4bunJTS8MT8HFmAULFicGnf9aU4qwqagZpGR7/hC4l73zbYIDm
JuOqM+vhC7+odX19IC33Sp2QBWyTdOe0OC/xpIG3O7/MGL/xBhzHST2wTXsMjgiz
mDnyekRn7hAD6XxaP2z5T7syAQ4MQHqKwoOE3XdBKN7rxiXxh6RCg5cVchdrt5CY
orG3PpnoG1H2y2I7wK5zQ4EJI45CT6q4MHiGKQ4EtgOzCqwkSt2H6BqhmLc4KxzG
2nn0s3gKOkyA/kz6XUdn2DWQAANuWoDVs/eB5aNa7hZaOjZxgqDrOXUFMh3lu/ua
5xhcdSgjncFSAAvnyFgr3byNVTvcs4UNUYlFJ2spPeAYWQwPe/e3Ct3ZoLa7alQz
AQPHWcZIorpTY/yDqkTYxbpQUXKYBkP3UiJKipxI+Wq1SIx8BQ8roQtlTY8aDkKo
YnoGLqfbQ7Rrx/JrvTOeiSac+2r2yWDouPlhCkPVfG/399QVJ7emiO3FTJtkgDOY
1pGj1ALb78nl+voQd/1zOyoLV6aqubFBRRBoPHwwX+RyqbXnH32GrMRcEkmqLOMb
SruXsMasNjp5GkY9iR6vKC7VSyZJ+WkJPSBfCuI1sVf8XFEn/1WXtAUHIj9QlNRR
Gl0V2a2cNlcCojwAKF6wSS6DZCUpUX+9Xtci0whcrq/22+XJE8zrYULqx3yVzrby
dYK0RaQxaUHFSj70ivb+OWoCFB5Y1v7HblE39bpYP719rYbrSwszMsb3YnUBhQE9
7PKKXVMSD+3Y9XvGUFVvR4mKDSc3kFYIupCQUdVceTnUg5UloG+uZj/lm9gCKzv9
sbIG0+yXcE8p8ky3/m3JSESaGYLdrfLwXwSkVpjKbuQ+BqDGdl7fuhBm+wawODv3
V/kgI49rjvOtcANbd2gVw0I37ib5eyKyrkWUTl1gCxt9WMFycYG+veB4DOpJgKRY
Z4AMZ0KdYsuyWz+hkbTqC57s9MsgYfGM+zkGwLUioM9CzwRMoohNssCReNll8yvz
GI5iozsT2nscRxVoCgrgiluaSt8HBrIEoskkD/4hT9wlE3b/kgOMpGLdXxAyxHfY
h6uliCW3epQttIQvsi9fzOEzHOCcpmVVFpYrBcJUHs+k4lZZfeLu+38lHTjMQuFz
9Tr6pJGGOFv6bsTqXItj1LiPRG76hd9mnLbo25aiLETcSHpMdfdFA/tn0akYi7z8
LiyXDybqat6wfB+D/Pb3qp8K/6LzL5MN/L9nPvQDbzt9ztgg2oJ7AAgsnEXSI1ry
oKZpZ5wLdunQEAWlexLzJ+X9fvw1mzetgcdsUdX95SnroS4mRQItQmurafbXcOws
6HuB25fR0WPlrNj7w/EcAZPQ8EFxkoW+UMFOEO7JboY5sCsNWN1JULINLnTcKYqf
+KJp4zOiOz4Y6VwZ7hnpy98OdUy4J7YCbCjq30xq22Ec8nzOHnahhph5H+uHRvUq
iBxLtZ1mU0/E3I24Nd6iLf96TJKNEfd5gC3ehrWvpGrN1fBvJynzehyXUzVla8VN
QMPuYMP16DseWqJqiPd+GDDMVvh3LdyokoWgsyJ6akRmk4jgnu+eTvp+UHKHPyUa
A8U6Ub2DFM0EJXML9KysnNuFh/k6R16aONP5YTSEHhB/gHxVlS13E4rHhujr9FXJ
N57GyrOZ6QThkGVw2/aIjfMKUrvjwyeKxS3ggUA1kCYGfMuILLrYrMmT0LoP/16a
G41KCbGcAlDxvIxWhFjfSkObHNKikyqjbWasKgp6Me8bS8q3ZflrS55nWHkWayD6
4/M4PFtH1ah5Y2xleDUlUfXHYK9U8IX9oE4XCrPlhDDGmG5T9tL4P0xojY6VqjR1
9kq69Uh3tHjfS3oT89PUZK7D86uBhmPwTcBxH7K/UrjiJQ9nuVrJHg9Hoy+98w/0
dC1qCylcntwRpN5dkKDrkECF59yAG9NxKJ/mUhLdxrbDsEqbmwUlztSnQ0MTydhs
5oWAL2tME2+iNASzRLHE5WTwr9y+J/XPGt3cYFQn+U+xcENe5H/cfZf++9DJhd40
r4DWQdOQK/DYrhHOJb5wEaiWFsDVkjZtSEhSp/HUVik32ScYh49fLrwi5Dnmndx1
h14T0grTYY/rjgEWn3jZdY1kKRSPO7XZSJC/ml1/pGRZ/j03K7u8idKCbWbZ2JVJ
YHThC9vXR2xL5QOIRD0hXoTSxeuyphX4Im9DnDDLUbLb1BJvbGJTQChgWWRukBZU
r5rB2GojAy/661Gnd3TLY9QDr8duOxvN07cu24Q/oFD3/jHvZIycJrWiBvgs8Fqu
2fX5QqN8jPbYbnH6PGtgsaYdRt97sZwdZr2x4BxDDjaA4tJtQZMQotTl9t+2BRhR
CHVMILmcqmLFjkuBFTIiUnh17FHjZavAyspaXXFpk52NP52d/q7QYvDUtcRLoO0O
MxYMGmFtHpV11moNCFX+n7OrXkLrVKxTYZvHuY5mEG7xCbP+ggMvTi0PRZ9cVGNe
NhJ0DVw5dgsLef4GgdA9bMBEgZl1XR6zNsNkj+qd7qUN8C/MhIkcVDTTjMbzRsYB
XMRnaIXJrQtuivgZtMYP3eJGlBJINmQPUSsX/06/M5K9OzY9yfc1nUTWaIcGLMY7
i7SsUFV+dwESHDKv7N1TfVqQ6ymmkutRv3RBDmjR6s64A9k+9bQMvwPWuVGtq9vw
iaqktM6nnxznvTyoq0XenUzycbi6ru7UqpWyuaJ0qq8LzKmY/x+tIlNaNmXSdaYa
03VwF+jRpD2idT6K9thACcqVjBzw4o7YX7NDHeGBNQEQOx4tp7nqt44Ur8QXWHN8
uSUheeU71Dwcftlar8Tpuk89Z85n0mTMJv13kntxWZ5FF28+HhmfTnBFpmtUxxJ/
SVyZRCclbauOmivy3sXvNm/S3nQZVTAlUYnjL21N8B5Vyuc06zfiNOLa9PRnav1k
QOfBfwY1/m6wqRcGFZp6t3aKJQtFG0SDl4XYCZL+Ebj8Vg8GAeJa0dZSi3kJGo+7
UsxIcvBpcTwk2Zejs+4jw+NAWfXChGQWvj0wiS/C6fYeWoGvp2Ezyu45PKaOzbcf
zvQrGESXUaNNHnhptOlR0W8eVbpM23DcVHsMA3fcIKz3QtXZvAjw2Y0tESF/bdrK
KFtI3dPB1K2VuoblBHvu5YSe/6Y3Ia8ntOVanVuDARuXOTB9z1fRpI1ACot1sMXS
EnCsXf5+eqegpJ4i4/vi+5hHG0dAmb8he0+DQB9v2IXN1bTtUzG8nKxnGqMtFhC0
kSp1E1Yw/c7j9jKylYRMbblbv3OUpI8/mlUArbSnYI4f9fyMRre0mQt2x72AMJlF
52Xq1PV8HTl3UJEqI4jrPhCitYhFHZNPKqS9SBr2j7ip2SeDVyGHid0KI/miMc9X
u3IkyX/xYwYBerZg8L1e8/nZU7M5I4PuDHlhBvgudHfflaGSsi9AJKqEWjvl7V20
RiFyDvqyS0HBs4GfvLTJ2+k9Qd4nLolS56YjaJ5tBeZggubWIch3Qg8FLi95rwdT
nRnOY5iPiJT9Y3CsOzhyvXojCL3R/m07H+5c56TSAuZyLM8UsixOY43ypLVp5zaz
hxUKoT+tDLRanrOAwkZOQ1Bo3rs5H9bBtK8IjQDYo2DM1uMygDdwnX9YHG57qvp6
N28nDdYwvwIyvblzpUbbDKZ+4Q8WvH5jxaYFneGQky3oC3kzHmLi7WF3Pqcf2N1N
2tm8fjIso1dVfNto3zBl9YIeSzpCw92VDSTTLu1RX219SU9zCjoBknC45eQjGvEz
VMnEvwF2RtC/Vlvtre3b37OktFk1Keidbzaxo+PY6eEwLpqeHmiEzMaPQALOPh7y
2rcOKgTo6LQG3qpKgFKYsvcJuQZyG7XIGnLRtdsMLkOttja5aIX0qWsYV645CIcL
RKZGfFDLrjpffkO2TjFYKwzu7ca5fZfJIEYSEsmJIOwVPo5thbpCuFrP9F5Sd+WY
vzuCy2Hum4XlZnB4PHdUYoxm+XRxi0YicQ2CjUaeLJoWABWwMXD+xwW/UqabkJuW
vwLsDaCLb4isl0oTndv2Qj/xPm+FcwoT7GgSNoQ9N8Jl2aD7VTWiDHUMc7+c4grR
bClgLHgDkTJmSVkpruhKfQ==
`pragma protect end_protected
