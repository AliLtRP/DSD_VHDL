// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:25 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Mi/2LTE/V/Xpjd9UhSnG2L7mJqDrkkMEPvovRDVctePoCEK56g9fq65WoaZnIMCv
5iDjCwT2IVCrqZ2sJiUYM6s8QiiGc9SVMPlt6huLqEuCHE7HTlblYvfiRPhEATdC
8TMDkYEmSTqKyen+aN8qo6xnjFYr7DXIjkyaaVbmids=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 9728)
dxa/UpCbJDprhC4TaJmV34vyG6ZOMjQR4m7dQqdrco0LXkCifEL44l/E14OqqHwr
BJJQZXDSQSpcivh8G/ov/coEJ9sBGL0O+o1vm5tbqqtr1MobzjXcJrNECGz8x1Pa
OjAcw2wS0JILgdpGeWMblB/asvLxIdY0CUcOIG09Azv5dc9iIelbt15BRLOtUp9K
CiLh7CkadktqNPiyXv1TcsiNOlRTQEh4kXYdLnWh7eIRZK4T3qD0nLX4Kv9UX+Ya
FCe7SsVkncPtvFqTEh6TK1q9SdJxq43DOwUO/6ybMUhuyUCX58dxGSleY3T5yteq
FoVJ7AXfsvP0EMryMXDR/gfCHte43dNHbwKNUM8ta02StG886lA5WmCeuGV3H+hT
BFIBQrkFTb+4JtEBubZw9ruk1PgSG9ngszR5kYT+NlarOZrDFNhCDN1ug45owzhW
4yUhplxw0c2eq44z3llgiw9QP2swwAvcn46fWfdb/CjTR3xwXhuIaKwNcVBRIPow
mBppFLgB8A61iOOfDb20P/LxgR4xei+neka6kc5U8LIpVhdrFiowRuvVWNAexLAg
ROuDtxuGkxJMY5rhB6TH4bcv7g4T68LuMK1hGFJB4Dr7pJ0F79zIYuG1iR6psUdY
+QdEyHOSXVaPjcwCC+rTmHWaNZIEpAaB6eyXqhovD0axFKeJpRSAZhaInc+towa/
TTGVTMdQmOwTJ7DNyVs2owiNHJ0bG9jPoVzn9EiVOFMMgEX/fuOLqv9N3vm3BnWu
b0IWWcRP5ahxTGVxpNaS4qc4fGebmVdZXw142Hjv5pHLSEVGVoMTKIxOdilXWM+E
+MfOKz2CMtu13dnl9lBx4gR3vRrLbx/nDBX+aTkmsaxIXlPSVFssBHI7g8a7IV4U
kvd/F3PdXpU2z3k1Wa/lYJLTkVaTPfIF8zHdC5/cg9/gCvovxSbdyKkpBklAaCQ3
zbSOJdrvNMRREBkwsUVVHuk+2Do+Y7HkmG/JwPfMX8RJ4T5KKXd/+mBdu9eXiWKw
6KTgIUX1BouQY3akyuxILtb1/KpUEVy0YkSdrSW42STyGL6qmM13jcUrqJwPNjLM
UOkl38jErJHqDe63vi29zg8Oe2kbuUKxQbLOejuTqYQe4FIFiwGTgLiNkLTgURbn
aGPqXBT/vEOFh5WrAszkzFcLai2A9JW6Rmq1xUtalq9w4cJXRljJlkDwJb92B8QD
OgSt8RqIrdl/n2N4l8RsE1iraF5UfGURATCBUlJGR38YehTxWTk+pn2vrWTFY4fs
R1gP5fN8TGbuwUhO9MV1PumCAV0P+f+MhQW4lOQP3BwyGbTX2SwCF9/c4L2VZMKr
phFG49lYk/VMsW4+fkXDLm96GWV98y6uxm1VJB97N3KzZSG1Xj3tt9NtlofUcaZb
x4PuhzUhXfodpIaatY5H5IUav3FVqFpdEqd0xdnUObRb5rHmJ4I9KHE2F1vHn8Kl
2HrfhMxcjd0T6D2EJyr4xkaeaxTI8t5JhWyBwCynzaZVp2b5F/xwokJRxU4ObjmH
JYswoYbzfbNdYf7xqCvDEcRWi/VKKe+3TG/5FS5GrGVPgRF4OT1rs20Q6cj2SY72
NjqBt1hfL2aPbxyhl+SIo3iaa+qMHnQM9UX67SXPi9Na+VMiBPenTxnL+iYA2hdq
YJnlpB7o40bSESG28dBRTPIS/oNL+kUFxAIljKlIy8vx+FggCQjVljU0k5ofuJrc
riWdh6EXsjs1tqnuwWl0I3mrMpNXtG+0gtSKv3KkCzvU7M87N1AdhZqo2Y1+J/zT
7deOvnHr9UvxnhsOlrAGLZZo+uB6Afv4PM2nlsJjBWj+iVUTdihvkvKcq8HJBx9w
VZjjdu1oU+ObqIHR3lN/UyUdG4IM1yeFz2XToeMYeSnfI2VktbPbcpz/7tHD0goZ
PFoyqXbZi2xDyoxQf/OyNeEsuldn1rCIO4j/dfRO15Om28UECEy0Lq08fxbUH6q0
2Ky7+Vh8JSXuiRCuEsv2aT8I5nw4glwdqsnzFlsW1gW0btJnFzsFj4hRTgDEh6T8
sEV2YiwdxDerlhVZtk3RbDRPyTBPd/9Lw6eX1WbMkyRYkJsstf0dF4/na5F01yXs
8vTHH1vashlYl6ojEI0/GK42+KJoBHbCarGpEOGqnWIajzUdwA47OgFlkkdi3jWT
os/aaCVRY/R6nKDSesgF6RseCHUBQslN81dnva3dUAaVio14IVEeQMFBcSHnuFTr
dwpnQlnx4eZgmtAO1adSF7dINQvqOxDivb68EHtR8exVge8Y5aTy2srx82nSswYt
/Zjy/zEiP9ZhMsU9tQO4Y2aVgND1RxANN8PbnQTsCgK/xm2wKVum8v9G4tjGmZvd
AigYeRsNssY4c6BCQ3amGiXGXgK8HE93UZHZ6W2XpKp+WE8tiL0wM84q0xbSalKo
3WREtOAg0hbzzlwTU+6jvHwBOT5K9GMVLHApyWHBMygXgKN43SXhdtNUM0BsgH/j
gHgvHyU8PwRlP924GM/vw/latjQnpE1TMXRB8ptk2zxntzxk775HDC6vu9Hag/Hv
dB5ukgtSYkiBLhUVLJp2dGjG2F2h5Oaeo7GwLJvOWiDnEDGl9Wz5gD9hJ6Z/yL+n
1JgYrYZE/igs+PZlSVMeoxfcIs/Bwwr6JZGXWeiGal/atvCkKa6QfhyWCWAOGYVu
1rEta4ygjHikky2XjuwXU3LZwLJFlD2bh3MlGO8I3eWA6eSlklOf3kELSZw9pgCz
hQjFStt/uxB6ZKE9hENRCc/I2CBR7ZWy313KGX2Az/H1kmactBgfOdSePjtIsiiP
A/LC9i9AVbOCOvw6UluhtlkhXU01LFJl4XdKYNkakW4K4M/P5kZta8L4/BQPWXaS
NUQIirhRqX18feDChOCGBHy4YbG6j7FB91StuQ2MtHC1goNVSSqCkb1Y6ZZWhTs6
JBmAMTBs+BngrbwwI7XQMMzAWJvzGhiI8Tj6YHzkvdwGHx9Rp4KeDQfoD0Rq6tRd
2lYMmiqVWVB9mIegvCB3M9+f++wSgsAVm5dBqQupCwZFSMvFLUow4RHk+cZnp2Fw
641Vg2p4CXgy5lndH+vkERIeytyGebolJMuMK1MFFjy4EPrK8E5Ll6pZK9e+4lIi
J/L1l2ixri/F+ZKBe7gEW+lJiUU3sEWIDVe8PJYf1WXQJdbJVikFwo7jmJkS826n
UO4yd4xhREQsXrvDyPJcpLk1k29eUa25tfL2jKkLDarjpGBK1be/k7uUMI97uDDG
wmzTxRjg18Yync+gEuMaTNRNu33bSFzZulZ6X8H/asQ6GxtlJVGDCbnGkg0XW5IL
68bO66DmY84FQB63oxPZFmV8aG7bs1OokfgW1wMkMpOYd0sKKRV9KA3vdQOrUN9Q
+HMy6pJBI6AM61kGB5oApVR6kS79dGKpc1qXw+W/LfYcMc9P+NiYI3kHVFG1KMwF
iMTRsjx/QTK1aa26kT2YMdzYdQLTNDdQS6iCczw0oXpzTjHfBA2qEZd6Zu0xMWo9
Ipt88yxfi43AictHzfvOJnYgvVgo56j346idYgbRtjfFoN+E94xF/n8BZ4H+6jtA
NQ5pbxHgO/1jKza8kfbE+8C0ZlVKTeUatgr70dbfQV3rLLg9HKhCSy32bHIQaxLa
Ay1+kcWPuoMMRGOWX3hawYcz9IUDQEEax+Rd92Gewbc/mUkgbGzP55B6hjf5jgUO
bis+CwLJkbdiKEkdjj0LcM2mE4UinohjWJS8Z3HeRbmvG0hfzGyr1WzPKxLx8QwI
173dlAubYIs3kyz9OnRx9f2BW8LXtQ+eBmc1M+vZIxq50vjY5WLH61PAmdFc0NVR
5m9wgqG4BVeUzm/p4ghOkaZREvcHwlUIPqiygT3qpn1Hg9qy7OxNiNd2TqMH/wJQ
fR+cKeLZ6Q65GY364tGtOrrKlBGYlqFc6K2AWQz+lHre033X+nHyTtqRaJDW7rq8
TB6McGqT3zKrSiS+9WfGmvwMyMBz3BojmGvcmNxucgs8JjlCDS35PWfQv9Vqclyh
IpGGW6Jy0yd8h9ZSCcLjsrIinjbrBf6xrxI6TXukCxstOakB+jJXaCxGcsHFExLA
BZhxe25pPZmUldRKIIMMXTU4mEGejI9jcigZOGzgk3aKHBaUbsvsSOTg6MgTNJSM
tKzcErNrnnwhpHHw9K3Fxrae5hiuj6Xagp3Q1+Xmp9YwQBUCM+MZp75dLHFVfWBV
5dRPlBg6+3SCgKG+Jp9/RGpmgl3LJs3K/2SEx7q/LUwZ0ogFgCipWVQEpjoyUjDl
cW7p3hygn1+SkUV3IL121LvyHsOShsHwGsNEzJdR13THuVgzoIh5yFhb7l4/Spgl
DUGjsEismy8rgCRWL6PZePGyuUQyFibZI0pqX4/GFN7sf4AI8bG9jC866sz140vv
ht9/1pq5NE9w1ehHwPNTJQyd8JaEhJNKON/FmxQ4pU+fsOsK82SzhEdQ/lNUdtmA
AjkzqG4XRKS5Mhrwotq4nce/stmxWZTOJ19iIU3VTFTzRPVfyTnvsYq3U6sQPQFs
v9YSk6b6kj8JJ4wpG4vIyUk/Ch9FhKJsYs7WwYj9NYuNwJBuPhHDuDNQRfIy8RW5
hCvCLXzoSOb5x1xsrBzqxnTbQ7p/3oGidA2Jf7r5tB707K3yRyxsrERh4kUz4m7n
l9AclCzpiCPZ25h5ShM0POXt/0Sf00umE1c1LS1dnRvYc3QPTZe0dndwl9GS7iw+
5MzgEnhzbAahk9IIOhw6yUZMX9NXKDMTY4cmuL5EM52BCYdzaNOXFzobSu8ybMI+
dQpbUL1Mtf7jpWY0HpNAwNH+zpzNCtd4d+Euc/2oyfoNI9V9x4PFQVcwNvGk+bSe
XZGanI4Egi+waI2Fcnq0YWxSAqcTy/dsQzjqZ+ZjBQAFoSjyS4LcNByD4jmXX9VP
JJ+CZ60AIfUWigeZ3kNeckUU3HXZXY28r3cVGlSsk1H7IXLERNdkuTFAtyLEXJql
XeUHqf1QFYuTIZpzN6RLwiVSPzlHmLlZWolRMDAL6IqsW6xf69DD/bLBP8QiFC6B
5UJ3o2wq702j1LdUr80mFWiVW1iJq0JbRzjCYD3gK8P/v2EpZUjeVgWhn1JwrCST
0g87I7YZPm4v92s/OIgByd63BBxCwpS674nCLoWkqEwiz9JTn3l4GMV3l4JXibS4
eDCYg6wY5QrO0kDe0SewlVSyaiTUHxINoQn7slUUEqe6beqoHnvc2/vW53PrrTIf
e1ayQHwKNyxftxXFSZWlBPmb2B6gykoGT2aJE/pY0cIpR7p8+W3Mg0rqv7o1ZxB+
06M7EeUDbnrKn+xMYsjiYuSQANhqHiTPOfhRBdP0qKAQqwe9DvLhfv2TYVizHyDj
ZYVWjjpcHuHrTwuMoEcD9VfkKPeWQEdT06GwyQzr08iuqQFICqOcCB+jeVjO2X0j
YQ6ATpnkQCwnWHJAWwtQLnSqe8ye8n1pBoCWxwqf/MhEPSsmPRH0/rHNSxIE4bto
dPg+CywsBdpLklV9tvb8VIeYIIU3Dm28zITA3DAOVhf50MSWDhNe9W8JpKAbl6rz
Y1FfwzOvA6joghBQ7ae/9bEyw2lk8HZPazFzrIcooYQkaayeVYDcG4Dm6GP53i7s
Phnud+txREStQ0iYacyrAtZCk3nHG351UYLl+UNOBxOJg+JahQit9YpW26cxwulO
j8fXwUq6QMlGok5zoyAwSKFaVAgGny0GCRh/fpwlgBE3Toz6vsiQCaVn+9RNYQAP
7KOGf8pHrufhanS8/DFels4q1Rl3GAxC2MqfNksFEHxCtkQAN/Z7kqoNUJrU+Ko7
EM48HhLz9kRlJVqc8sUJyNVEqXVLmDgTKYZAdViNg3y4wd0PfJ7OD5M0/apLlMx+
W3xCmGFpRJlOuZgL5eY+Qs0PP5c45wBMttsIfuqBu+/zbM+1jZ18jPucebGTG3z1
nR0pypCX0qmUtOAC7YWCDfv7/Ctyfgrb3GmClHuyo1WF8eXecaY1X+4ii79Equs5
zABLZYv8W4eMV7px++foSdSnUBF9BtwRtFI4QbYnw/1RR5odTOPsevsaEmKPCz7s
BOQ0mkjJ1wGQ/uJHvTZ+whTpwRewllceEh7voJVUlWX/ExZOl+oLd8e5kJe483qj
rdOENjgObmosxHD5i+3mSdTTvxt77KopU2yMUkFPgtWmyaxmBbEN9Ca5bxUM0TAz
0U40BPAhmVR3qFDzuxB4zUjfUjEakWCyJlLLghzKd1NKbfy+RPQv8Pm8Q4no6+l6
LjgC7XG3DVSThPNjWUbGlUMXDqpul0DDxqJ6DBadZYixGHg0RPLYYRQiV3+IKyNb
N9x7uXTBTkYV2VtDp54LCflqyQp7Soc/s4MqLjZcK3CbNLQ8ptvzS3nWlg41JqW8
OX25NHypgYjdmMIXhh1oH/FaoRzrT3M4rQ/H+PFbGU31G3baPKFWuHS06/Wvg8k3
ARBMAYYifUzjnFwVDLJOJyeg07dLri30WjcwiS1DctpE8q74k6zttnok6hvzvWDN
Im8Lpg7syfeedLut9WG8i/6t8C/8L18kbonFRJPahSqguZjCx/hnZ7LmG4xyWLCE
yGLTIowzOw9xZsGgERN2uWd6A7aDn1+NVCVr6g8ZT3JzeMn1/XuGeHe1tFgMWjDp
mG1k7EXskG7uG642w1FN64tqNaPNHYhe3ddE4mcShGHC80CSIRnKy5vhuhe706DO
aI1GK46WxqXQqhcT7GFo831oLxf4FGqLP/zkZsPVNzj4XxYH/01rWGhATkOl5vCh
lCZUDC5FpjjAZ4hUEK7YuAW3TdtEbSfEOdeRWGeG9o/609As6HS3jBNMjd0zgWXe
y0VV4OoBP5hL00S4D04GdcEVMPSeM+Y3uGS9BqdRhmB5ALxuttPP8A9TMs8Gn4Uc
nfJaQFkkynog49xh6IG5Q0NJETE4pyeBUab2NrIUtzjE1ncVU7pa0FRcAt6mOB9M
zz+Uxjp4v8zrv/R0Wj6s++t3vV8yD3ldXT54KubPwgw/Hs4iZkGaxmPz9Tj/maeq
Ktm8FGK7N7T4XszKIeRKDsaJAW/7A33DLFOFU0nNiRXS8XIvRN+xf2uaz2kzzca7
joo/E8irWZC/gRiUx7ROMdruA2FpH2Toe7+xMbaVujEKMfO+bXvzmWKzi1vg5HI9
7o3tK+vdnDoUWFzrnS8KP6jR+7tM6bvrgmqVOtVMyY1aNGFI7Gzxtg14VayDuyHh
IgO+T0XLKMX1dgP36ddbR6yYIKzAn+jURH4zyfLzdhVUBuEBcY2QUfRQqteU4suV
wjYQqO+2KyVPedVRx6gGQOG9hBdTZyWvzmgAryKdB/trP5jo+UgTRvxTQI4j7CIq
bPVi8lQM25ZSun+zX+VZEXizSMvo6VUaa35HFMBQroyTui+rx6h/M9DUSRl28xa9
7z1eZ7WJNsTU6VV7qeA9EoLyvPDb2bOh0lclFEIIyofSuxzxRz58v8l/91xIu+EA
8kINs5RUCBa4HkVEkUwBSY+uD9GbmLt9TvIXj7H4UFL2TONaOilzu6e2Zn5KyA5p
DfWBhkaCXn8D8EgVoO1ziQKX2O9pWRjcgAXiLGLUdreK+Zop2LSvhLjvYR7Rm2Cb
tIplJEeA55sfgQJNJIDY3r0K9ALRxooKe9uAyqRFd0p8UJwpVVQC+g+warbYJ+QM
LOScsdV4fe40BU+qvn0/DWfZoDR5wDaLwGZeue0aU/srM19Kq6/Ys/ftPWx05YQ2
GG8fHmGaG/jHGj2zrYO44Fwu5HIOdblEW2P00V/rfEhyoMKM9ep3Tb1JPbPWiIa0
yZusNuuXSVGeBnw46Qcq44M2Gf7V3yMA8LTFMq0J0zFeGJ2zE0oLW33KNCEKc933
v392Hr9YfoZw1cgPQxQuvPuIaI0Q03AvvRKmoJjOYZEoZiqsSFwQukQ90/JUnSjn
/T48HWMwdp/m40YGjvajZPyieuSUdUz4qk+cCPHn+2ekpYvUyrRd+emwl3tZE9DD
fhcYd1nQnUHK1EUnBnYEVj7irM/j1iDrvDmuzG54j7NsVChEhmSgcc6unMICzq7i
T27DP79OP00HeY/HXf01r+en9u6Ix6TzARA1Ys3Egt/XEwK6gl+efvBTSZSVlpvk
9Q/BYHedRdYyj7KxF5Tot1E75HOvKKo7Gm/ARpND0iMfCK3hb1i3LlvkY5/rmITd
jdk8W6OWx9oLvAY7/RdZxXO/3Gddh+SYSG/xahJM5gyUUShIvpCnXsbtawbeCksX
9+8RaYsrkyoKdfK3gIymfdeaOD/HFDXsl3RCk5QgPU6etNCR7ksudxN1W5X4KHRL
xvo1cmO5OngVKKprP3iubho7P8EclMVO8B5xn1sRIdHxJVhv6S/d8hvoUI9XkYQS
tw/ICGSdQowohcMtvg1KfV+eZYF2UL4/ursxV+Oc1eUB8TJUK3d5rt7vNnDidmWp
jVNHjho7SeP6GnjkBmor0vdGdl5BAPY6Z96Rfqc7D1aMECbnZmbPGqRIGnElBr7N
0dwSP8trT7XRBxgP3sdNpSbAcCBja6y9RWUvZw9a/qLk7jtis3oMi1eRbGnRbtbf
SOe0Q6SC+LiK4oyd6cOsZpyYLw1HTxcuTCVQ9rumrWWgdWXRceRKHGtYSWivlF49
nZvawzg4flQTMy0Kk7kLu7yuFXXbC0aoyWb2MdvLbCtbdLm5lTac6KnotqIeOHYW
d71YxFLyM081TG5EAMbqgKXhMgSeFcyMdSqPN/anL7pEI9Tqwr2hnQktyGz/Gbva
7eNGmSMIjJ6Hlq0gUyMHSKveqIy2Iglcwm9l4UxeWztsO7aFENy5NI1RypjNG52w
+FDYL0wxBBaPiQdZ8Rb6Rkj5KgQWTyEkhYMSObPmjVCyAvyIpniqkbtFwHToHZhN
FICcZp/LXrr8LleklTuiBIGCrtUuXlPAnG9vsGaLgMfHZJWTgiRv8paM/r6/fTOy
GzSEvhc+toMBALFtKCuMeBLyjYMHfz5iE+fe+R1eEWU3Z4EYXFFw+JXpw/W/2Bzk
28qCoDFpKLX9ErsEoRwEjSE2dxqtT6qAcZ3hCOcztsFa8NIp/morxhdHf951CJPs
xI1XOjMU1R94Ktb3KUwtn5HHWh6aCxlZQnlxpHyR6fmos/UoHO5ByFCf2Pp6QHF/
pyb0zV90L5uo5wcVQuywt+Op6eDC5A2iJEuNjzxnXTj0HBwpHrwko8Xe28CiM7sZ
CravTgNmhp/ncgyFNp4Krcwe/OHM6bwRriGRV29sFNwGv4mYPRqwb30f80tSa6Z7
k1tB8KbFgUop75JwvVS3YIRjXih+KYL+Aw2whgNJmNONQdPqEnxhJCUQLcxxIfVN
SpCZXAoe3Tss2fpBCj+tym85wjsdLeyyFKRpYDkPSdRxPJ7CyRAhLS9GJtg7oDep
ojNIsQtjZOk3mlIOPYtqzOT/LlUnetlE+sR9zbUNM5kC5sm6U2CQzOdfwHFseQJ6
ScCKlxBj5bpBRNiAh/kKdkbOzFhAhr/l81JH8vTwUCQDbwUfu8WkEbCgitfe7WDA
8qniLb/TOXJIOxvwJszvxFAMlihxFZUnJg7mHATvMDGd6pXB/aZRswPe0PUXZXWa
orHBiQj1wGHaBv7+6O0W1aw6pGLKuYF7SGoRD1BHsRjuK3i3qKLBVIT7Mqbwdpmr
ZbFp/xqCkzPEglUKV4cjFNzC4p/Ei0s/a23fRtKyfXN4jsjaaoKoHBTliRQcp+33
7ZMGURDwQhn3TshLpPgGPraAHOYcSi9Fks0MUjKru9sp+MmSEM6OvkNV2dFkbcMj
sWHI7R+hi2PH4PNVBrdGTQE5LZ6PsKOmWgrISnUe6D5fuU1aPUfIzZ9aG7zjloGt
OAuiy+xa19Pk+tSB7K7BlpfgppPP4b3m0uH4NzwD8WN4qeCgRrxaYgewzA0gFaOp
p9azJx11Wep4A93suqvC3ETSYFhT7Xqljs9k488iOsYv8EiEBV6A39duPmsbKdHm
+PYfSNosQooDndUQyEF6yhTpUyi4yEAPWw2z5YBHfnBFevbgziNtRRem0vQP+y0O
kmKVa+6rBiJMzxFxQabQIlt5//OHTyajbtWR/rAMHHD0OxM8EXspQc3dhKqjSyKY
q52z3+h5UXdyuGm+IS1fvpNH/k8pZfWzO7Z7eyJo1Q5K+G7vU/nomlF6LLhjOUvf
jYI3i2tO2xArdnwCjWUffy66V2NXC7Wj3jAowySJ/fCNJqmIKQJw/tN++N2NJ4fL
+Jrkik9y7VcG4zQ9sYUlUK/wZC8q9wGrUyq0ofbFcXQCAnHDPwjLyat0zD+KfOw9
MF2XNqSGuZYr+XFFh9xKdgUSaPRNqOmWMG40seVY287FMLTChg4MeALdXJ6I/xzZ
JZX4xaB1V79EkdMIE66OIH3SW/sR/OvKy0LC/f/jGVVgZdg04USQG0ofQHE0uIgs
LikhzbR8uL+xvoeWKOXam5b7/oujPB9zZdnLkyMs8iTHqLWDqh/Q5CYP9Fph8wIX
nC8DYdwbgyUX06eJ3vt7dzuiocLDvplLiP0oLzhqABqBZL7FCf+E8vnX63T9604k
1NO01H6rzicO4/NkaQRWwgrSwSwBkEh6rJTLkjR1PEhDceNs+4bgbIgPOhJPOkv8
OarVPCCl8UT/548rBlCDDYeUliwRzmqtg+wfZzz5kGkmdORma85WlAZVW6KrbLGA
TpD8qHx8RLhaPEu4p4+zDMr6PRBEqmE/Vzty6fJZb+0ThoM3bfDjqzJE/QhBfeD2
DmCWTU6MXt1wRJ6rdbakmGWlX14nUz/yzlDrk/LzTzVBE+lCpbY0rtTEA7goPraK
W341G5qrhsA7I3Wn/bun08Fdw5WoZMpJXI13A6tC4b6O4rxfMNZAikkCyI266xx2
c/XRDI8l0iBzcTi7gckYu/82b8mePX7DmW9LaTPv5KjrUpv7bbAooYGKD1jYS6yu
a5FjdpcXLwouGf10D5ACtvbc+Xm9cNIqvezB2QtgY3jFMX7DdNp2UxH9b6GlSMQm
w3i2a2U2j4WlOIq9purA3pvmLaIC4sRdLGeIc6PRq+FRrhrgVGOsux0CqQq3uCw+
fEussIoFNAYd8D1tJoT9PjNKr/m8nMui0PlqdbUoRhOxMvmZRIVfYsOdvHnJfDFB
GqWPkVCj2G13SzRrhbIG589qaCci3GrC/oHhbpmcvk0TC0TAEcHLVzX/hE00Dkmg
4dal8/Lb5FqMlBCaiEa6k+ogwaJ+vfHnH71cVTK6jKl+o9gFkRirR6967TGiDprn
EUDk7yRUeWFrfxmF5pUVZ88YSax53H7Txpiz1mqgJxn4gdAaJyOUjz80VzR4a3Fg
j1wTJRZHYWpuUyxkXN2Vsv/LjXhQLE/L1Cux4CDiQQqfPuAH+ynhwP7iS/9fyKxa
6Z6A8rBgFU62FqrwoZC7xjcckDEUE1q6kHNdm5yt/k0SKg++ZtbZ07cxWbL1/d39
P97JWCrXvnnCg3saOIkoQHOau8JVZIjdPnZMXj09Y+upmi9xr/WHFRKPPxyh+mor
nQQo36kNGjRK8tnS4bEih6zYKjx685ld+8PTKj4RDZZ0DFjn1AhCqmULRj6+y57j
xTXUJj1uegT9TRgkObQC8+WSTQ35SEVqhcZhkdtkml3lPiCv/NOlD9M1lyVCG+8U
edGV9/0ItE/Hezw750S71oYlgOhfjos9TDcgoJX+pUlvgab5AVYxxMjhI6gbXi3d
ie5OZ/PAgSxh//n4qOYU50vbYLcTQuQndfaC5aYtrugEBbVben9tLRgfJrx68wt9
XX7D9vRMxeTfPWaDfyQlC97V+KS0/OxKdcxmV0J8YnfUwRzTPqve2ilfJrVYw8cl
GFOqjdCCfOhATyS02veoWH7KIEakCH2BvDhrm2F8FpxDpLstnic02rG7qLjgi/Nm
pu+xg4pG+/ENwXTmz/gPiL29PM4y7rkkTC6Xtz/7RuO3KJURfSZUrezvXJywv1Fi
J9NGC0MqZzFL1NmClPwlJUrhtz8lnYR3Z8Vf0mEPGIWjIixG1NBaf3G4NMFecPDo
AaygJ6RVy4FLCAe/7nTnDhrUlPLYiwNnT+pq3MplJMmG9FRwjyKEfYsKG4/FamuJ
c287Fw3QmekUOlreFU5Br/y7jtUnOF2ZIE7O9PWK1t000/TVqnH1E0goDnUGO92j
nFl2QL/ZaFF0l9ipCum1ldBln5ZJzJIb3OHjm+QQe/DwZJKDKP4f5BhPBFjL9gBq
U0k7VYWbK31Ssa+6jh8sFNrY/7S6KRtI93I5IzJ6Rhn5Wm03v8Y0o4CAmupV5WxH
ieqnBAfqFQw0fns7u0PuXyuHxalHHWJjHXPyFgbmVPkjhrd7feldigHA5pVJlTBT
OLn6F9AZveqvlf3OmMb+3/hc8hD2lXi/lgtXL7ZRe2gKvoxEH6LiqTY4KKavVIj/
Ax04X+xSNVFQEZ/4khcpsk0dDksfGKosGNIxlH15Tc+TMxgK/txWJMXNZAar8oym
oZRmqhjdhtwlxURby0g3mQIgv0Ybf3zwf9R98goHsngFZs8WE723asLy0PjZuxKY
vM1QioUDh3evVYjSnZdZr+q1ZFxeVDCn8L+tEpsZlNsD9xTAB5DQi8nQdCsJnv18
bJJl1NUW19/qcXjxO+wKW43dFc9nkqAwqM3fCbewlg00rzKajX2hp0sG8IJ3Yeie
baK818FMS8sNjh0TquJQs6DzPVsySgyq8BIoGNeHRXQtnEbWkwTuBhiesCHl7p28
GZjL8lEHI0M28q4YL+zMdVtuCNwedzZ5S/x+loLCsgOSGe22yAgV/MsugqFp6N9j
CFIWL6ntpXgOe2rEhx45aO0F/5PkNJ3m0DtWeXdSuXBqpzE7qACo0xOiTb7QIxsA
YXKaxB5/YPhSTB2vyjxTBHKuFcL/Oe3t9ShTSXIDWiLfEleCGPlSAilulYSLTc1r
CusQW1BoJmc+LA6yqv1WO6HV7F3VEfHXPLWljxgePhM=
`pragma protect end_protected
