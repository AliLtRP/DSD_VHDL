// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:37:38 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
mjSjUTRVrCdZJ1kKx1NQUE+3D7VrGSSfuHf1YuNN3IgEgX5tE19YNCzJbm8RP5dZ
GjZ41qG4BhP//ku/DK6gdKb/zq0GhanJ4wXqL6az1dXmOPsTtd5HWPFHiBwMI9V1
OT7+8kPq8gyOY9ToAoYKkec+LRPm15L3a8+VbTwVJWE=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 9520)
ZkqAi11PPQdi7uETgkbDgW7ubgp83B7NAHj+RdcgsfgP/pjLjJW5dboP3oop0P5U
p8V+X+iQUW3P54C+kFylZv39FYG9JRwy2hb2fxHwmmOML4HY6IvaCCs0RungJODv
7wNnIfy7xIIlm9JWysvc1dBj5ytO4NIQFqtZfeo+LSiYYVah+0eZGAsh9LD5z+3N
ltt2I4Nb9Z7WMnZ4y4T7mfW/CAjQuSq0h201D5ijyd6f2hcfl36q/9FCuNldKBe1
/aG0U94rOx9U4uaYsSaXkfBLjY3HXLC5HyT9u0rbO6dahaNBz/zUvxlEJUhp9PA3
j22hYrgNU2h2eWDF456K4EJL6g7EMZ2utNgVpqNxGkLZCQX+8iaArBe5B82VW6r0
e2vmD2ka3CeChjKXSv9CkWlP6qkSGKXJlWrqMPiohv5JOC6qq4hNkfQKYjxPlvq6
luS2TEvleosYkmrE5AhfJcmA0hX8CrbPbM3W324kuSPSqmFz2lYIAPBn86Tpv3+4
gJ7yZvVCK7ff1g/9p+bDmSFE6gxU4hOn2FoNTzWMR0Wxup43J5i1fHASLe3MGqld
VQviq1lyWGciNgxOSQsc2vlLPgqvmiL3GTWo7nQfGeEsH0t7bWPnVisGw3v6syTK
BP+bPCyGCoE9AkrCiQlioFtRXNlEP3cnxi7iNel8EfqcOT6jxRmg8VGiWpdFcCon
zCLY8rpdwDZsZiUWYgKYZGL9/NdmNHhBcbKO51QVWpgg05Ko4m2sd5vFmE19QZv8
txEkgm0s7O7HDrTX22N+uQPKhT6+gSbcgms5ybR7aSbktEhOu3hVtFgLXnax58fL
QeerPyriMQhyiXZni9QJR9SYwdeiCNosRGpvkddULh0JBMjGzKw7GzhsbFRUSn3n
vJbLtCplP6sszPgKz+9iDpDmFE8S5nY7MRCXVeMSonSeC3zec0bD501vVyvnDSmZ
4uyjFksubicDbzOS1dNiTFg3UD9ok9Ef4Tk0/jc5iHnvZmMTP9coNsHs8tXx4pmT
vQABBUAxkm+yqznd5WIK4oDcKWyE7yTtZtx0WQaySIBzt4I1ZPR8FPkQJK2kydj2
Q7A+al2gzAm49Nka9ypYQ0sBPHp/Y5igvy6bWuB9T2EwneZFm2YcN3PoInn4wnVT
A1Xm07+SD0krChMooRrlu9z/LeyilrQ6vgdBY7D1WW5uSybZGFBHTZaNFm5wfKiL
RRa2F/fyoDQObtIODsiQNuDM4crDwT8ltpraMwEhF3Lc8aoAjjnYbeJtRNFAxDqc
GoUt+Rvsm+US+4wnLt/ZKkAA6v+Ax+gKEwP9IMkfeBHLf9IB0KuRBKgPs+3XXJHi
xuaNbCKc0WhZnLCXH7k7WZ0j6ZE2TRnk1FFvZiaWhbq471gB9d4G5nvf7ruPhTBn
vSSd8Odi9KZQsCE71amcQ/8UwfD5P+WuL7/z6mPChNU4j4keJ15ygLyBE8qzqkoH
Q1fXcdN5xlxe3MNBgd1KTMgZWtc4gX8ScMLhtDpEcRbAL9c+IxX8FDS1xWV1gVgS
zVSVNkahpzjMRWtAduhQb9aCNEBgNRbMmghCx/gONQ0tIZQxF7ps8Dsg433x+h2S
M0iV/Xkx6Ozk1Nm4EKtW86hYpm706c7aiAs5NNd5R4Soq27eFw2P+IhCuv9NpQrn
ViAVYLRttAxmYkM6vAwnbckh495H+6HxVnavnezKpnvcWlHkD3rVCdv3S20pW01H
cUahJYZpbFPOvoFserShs+MXvMer0SOTh3wEVqg2/ARdjR+6WTHI54vPwBrQFZw5
/1tA8f8uf6ISwAbUluPCpb0hrOcOTFkoovyvk4gYcW2NT2GVXtFe+IZmVkl6D/GJ
FjhAWpMfuRN7nDK1EEzMfLs42GNqjvN6Lov78QT5YK49Jup/Mn0/Ga1jyldX+HwS
Jg2ZlwhnEvnA3eaKfQC3O57C/imbdQhvadbhBk2uPyq+qvcJp3jwc6jh0d5iDLG+
tE9RtZSaOVA38B3FFdEO2ENEkH2w4fH/op/A++lzEKvgbcjk9qcWDnq4x3tWgBf0
jMjFnDe4QSJKSRSWxIJmNpAm2WCUZpCOegrth4LoaDVjjXmiJn77rtg4EPtTDycb
5b2Q1ck3OnWskBXsO8WTt++DKi1axMkQoNKTkz2I4VRtYW9b1H/bu6b2T9SnYux0
EWNKRqv0qjCONFjLGfXeWcudmNSWR5wQVsmNr2CIJHXEAy8gDCG4aU78Xg8ki5Ru
oBvPp3NhV4/ND/4jzbR4qumi7mmqOzR3XY/K6syfxdb2EDT5aJT3dqrRk0w+CH6t
xPREaBcmIHB8XVyhThpqrmB3BI1vxigmXBG3k1fsztdre+CMOvd4lb1ejqf2mvpY
1mxiPoa+69xMMDqkwcsffsWl6on2Wok0tMZd+S5AASTj+jPPhGpnaeZzRQtgnUZT
GWsT7Fk6kTdmnOgT+Em55lgCqaDj84cM6I7B4lccR0H30HR0v1wGDMzaGZK2lY4R
GPDjT/I2mr4HjczTyavAgE6e6W0a1UbwF7TeZtxfSHi1T4syUC6slxnAt5ZHNvbX
7O/4873x4JQ1b/R85zgYSwJQ5a+WUZxylxMzKyT68ZQYRAc9xXZPnUpAvq1oB13q
sMV8IkoPg3yxmbuWEWi5ZHTIXVCqYlKUhIV4Sar8YVXgga+PAkSM6Mk93v1fk23p
gLHKBs5v+U/hXQNpm0Zcj0/Pf7zXdKaHJkxgLPyQtyGusekOp800ATFOLiDxLL6Z
tytRQJWi1YAwznU5KWn/+LjpZTFkahBIb2znNsszQUZo5c/M81Q3gPCBN97XbizK
MlDk6o1enjNoQ+JnF7iP0ZzGwywzOj3GjgHN0fLP67T3XoC8IzLLK1Q/ROGm9s2p
oue/jt7nVbBjPCr6xOZKYgN6cFNAWPJZAduGz4ZgdGJBkCLBVp8jKMsYm/zyT7jo
n8y9DLZU2/cOJNjJgisFRLji6d1FWCY4IC+Nb8RVpvwvP9MaUQJCSmQPTWZinv9N
lGIdU9T6uqJ+lsTfVdL9DOyUSMhOLkEzLe1RoFBDtAERWScM/IE/hzQWYUcYxMME
irgCyiC0xXcLtdENMATUoVGfgqMd1chJ4DtLE89avlEw8cXw+eyEgym1vBn+QRJr
ShWaHyeCQNOAtuW7JguKzAcyBr1GmL2RrSy4585OfIQC6R1KxfOd/8UFDVaFkiU5
MMVreNTCAJ2+cDI+/JhbQh0pI9tuP9da4eQpuyY04IrXg/ZoW8nJbUh5LhxD/TMZ
pqxabkz5ve4JgR4on/fcz3y4SL38JyWH9MevuajpyuoNIhNYKJkmviXjmnDaDEY+
rcKo3ZsPnRXWR3+sdeir104F8yJ2AmFBl1etpkiEOP7aLzfSEIfkS7QfnXWj2DXP
0RhwQKYDHd9wtmB8nxyvX8eMfEdmR0zKcV0hYmfw9bCRHx1CX67IkkkX2nwQD0Uj
mZ7eo8E5FN1eQT0SfVdl5M8qh/OxZmh7j+fbOr8cyGHI2oDLntE0IdBQZE8SO+dA
hnczstLc5DLUdOpuBLFVJ9jNr2eba5fPkkdt3IghS7+2wrO8ZwtKFuIfYkaUaOBu
hkfTdhWgQk1x0NDaGlHEDtRt+Yh7XGuF76LKQ9DZ9Kz91Sp/mTQTXmG07nRqprSL
fpGrt40MjfZ48800LRE9gWeBcq+RMUlZJGqOJVuaRhWqgSQgEIY47gSnN3izWXIg
i5KFLhMF2vbhF/WZmiCDW+yXaA3zzElCqDJEmXOHdPrre0PIS3Ry/wcZPFOIb0w8
2MKXH6BWgVPOtO/zZcziugWbzraqXKDY6tkz5qmCUzI8AJXbwKVXT6PUcIgaWNs7
/QKbbHWkPSdGWuVAQ/0cUHdIcKOeNGwNVquOjSo57d3VOouiVL9XiHmViZM0JgMQ
BHMXQ5rOW5V2L3O7cS6JwG3VZEB549ZUpUpSauxgi+ZiOgbdJwzUcZBE/fdb9wRF
EOSsikjY/jmvqEMWi3cR2celPD0Hqjig4UpqOKMDJUZt5lqTicQxWu/YL4O5nFtd
094gKqbYtvOetdcB9dDS5batvUJTAFZMk+mDALCsugSoXFAkuN7fXj68zlUY3tPD
NqmTWrbuAOVNwq9SvlhWoeHBmahcrcVL7facLMb57Az3RBSvn8AETlswHAau1QNx
FaQpCyj0FqSslmx0RihLxtCExWTdZTjW/GfilfnSylmmq0OQwCsFwHyvea7ULLkC
/KPY815beD7lP4CvqbYcX3Tfl/0xX4QmDROaLx0QrKDBadyEgXJQtqlfiZ0KkRQ6
Scz6edKivoBqAOvipdnyHIu1oOonWdVJb5gCvhLlzBZ3YSR6YLx0Ctxhj9WAVr5f
jbj1NZQlKahf67xwETssm8XJ7jzFYFlW/PcqiJvIXYCPZKLRsqv5Gmgbk89Fhgrz
PbIkRYiPQW3K0MPr50/inU7qVYBqCf7RaILavYrvBfTH5x3pNo2kOqEXSALEcQeI
ItSKgLQNQ6niRgsfLDMnp1ARc4FBJIE/B/Fcv7BIQBH/q1WLVco+UUdC/Y7XAPO+
Di/JL1W7qZpw2fMNyW6B1PoMHGJZfEvu/GinTUmLjjyFVMp39o4tNj0KZ0JvA0Al
pE3uJJT/dx6MQvLq3T1XuKusOS5GHTsUdRqhE0I6sHQlzxaq9j6vByphFtTbMP5I
oJtRbGZxQ36PqdW6E602xpppYU0pe2S26jqdqYe0TQCmlyTOv/D9Ec7bu8smYtMr
AfY8F4ezW/u16G5p/8ogEJbKpuXA6lY0KTLKb6z+LCeT0J4tMNhQTKqVA2z+RN1o
y2uPqsPc5BKPJpYGM443cvEbFNhyPt3TnPEKP13qWuwCLS273+8fdrSbTP+evriE
Kfz8qsdTAdGvs6RrZ3HY0cdGM8POijxPSCDVW634MBliF86hvvj+E1d+N42RZUP6
7ybNwe20v3aElvYMIVo7WmcG9zOhLQmViEJoxpe+/GMzQbjG2jcneTCi6J/iJEl/
d+ghjKxcDzXXGPhO+UiMEM3Z0d0BbIzhjXiwJRtBY/WhEFHWp2gFkNbcmdVdMojV
uCRbrE7x1t1yN1uA4If/0HAsBoZP1qLVLv697O8H8cE2eV0xm2eotuVvwyk6ue8x
m5RGVumOVbgbBWObqqqFvuxzURaazWzvNTpdCjhS//Cfv9LLD7+kyRwvHKTHAiLe
c/iV/YJRR3eOqUb8LUkLX+zqNbjWrMXtnxmKrHGFqia6Swa8wUKq90leQE1G4fxI
ANy1QazuwtKCoeHsAZAJsf7WaG772AiVG6klNiWgeUphmQDrdbxsRYGKF32gsU0k
obUIxzmfmv1/zO9Zu+a8aiupRzE+xp7C/9TzMSLt5xVALW5VxzX1J81uvzk1LBNj
zM1TjcFQGr5hwj3e6Rfe/KvSy72DD377fdBaRQO5om67funbpZb9l5QI9jKcBkOj
xmpNnpeMWc/c656x/KIVfpf4/1YJerV1tI4LDb+vFJHIRDgf43ebeJDnlXcH7a4f
9B6a3cCtSHu2zGRUOuclg22BOCgWcrhVQxdZzjE1TNP27UU+/uiDDzV3ZPuW76s0
d4CSI4bAIai5S2XYcfj3/CPZmna+sqkRCK9kCkyLAcEmGL4Eqf3SIanMI444Ssq9
7uF4LvQ+NeZHAC+z8jKylbMVNWz28D8KSRyjRbb3rS/HMcvPZDtuXYCdP6r/aiEv
Frve4JYo9hgLu/PaM26apzDCml+XoY+yJiisBwaZCJeolVi5WdjPGC7n0XdalUsI
tclWMaE2l0WEwXqsmuwi04qH4CKkuCHdL8x6oA2D0+DrPWlE2ktR16x5ZGticB0l
J6SNrO0eL0bjwd4CTNVWinKWvxKbCGVdx8LUzP3rVYjVkhnbe3FWLP55TEgP9dy+
bvClKodAt4CHisxtJnVR+aapKBbMCBZCnSWmCakiWl6EJ8q5rd+3gXiSkk0AcCwp
8grqU732tzOUAyrmzu3qOrUUDmVGBabr6QhC4lGQkgTfczm7dDsSB0npG7Hlebc1
btl0JpF4sWP8l5AvL3ji/hC8mPZ297klmSVFqmJTIDKmrZhUW/TNj79/g5eB6m/c
Fa25kWJtqj3nKpNU2bFOmlVCsjMtgSa18SBnPrdpKAwq2e/qOawggfFGOyp4Wj9h
piXYhRmYCoNxFDqhrflkQrG7X2/8YvlhuV0P4JjOXIvTQasHR9JpQHy1pEUPYSM8
SxQhl4JE0P7kP0UQJfzR+8A+gvKIVDko7zz90vARkQtM3K24gy9j56wtQH4h0ms/
BowJQ4tHT0Hd3VILp2GeyP+zO7k2hPUXFQ1hBMOlySYPmS/kwCgNt3Tss6BCgqYk
TFBT6OfSSxdYKGnvN62kKYF+8KTTAXzKdKPms3aiZCyW5sH9g+nSvDESey2zWS+v
/DeYbYZGXD0CZGkCKu+ur8VeyfhwRofrM1MQ/vrugaF8HlevzWUBg7BY2jQgYkPN
DBbuLLiJXjT5S3hYpYsrZgV9BdC5oMPTgPsVDLkPbQ41vzKqnnmgmt2TdK7gnh2v
+BmMueo+HkOyJYacUfG8fYjMXdqMLqmnpvZnC2FusNcgU5QaF5wCXw1bBq0ym2v1
5RDo8reb7dM2XATxN9tAy9A/ebHhbnpDfD8zBb7L0gkUNhdMQW2GE4dEMzW7mTTm
Z6JRPo3c0joPbcYZe4bkuKRHDc/n8PZMKElVGroRAluuCVhbJKGAIxIP+rBDbhuk
v028PPtFXvVV0zqfYXKBosdovOB6tlWMXrQv1wFSygdX73GE4PUiYfG0xx/lCVWU
KCV/Xi0ViHPSTUaioXquFeJAWQCkBHr6dUMKcizblTTCr+RH86izIZB0LiUF36b1
CSEHWK5F7H69j5WK34eesNEEjqMCl+DNm2t7UfF4vhF7LM99abJieMVRVhHRkt3M
ELIOrAReEVElJr0nmK+PuJUw3VPCB0O+48gIUTgngZUD+v4BM74zrTyZgo2MK9p5
6I0WHEkMMqfDQi7btAbVDmynSOiOKRLiraE8GtIyP7a9L2UT8IafGg5a4zTyVHqJ
Pcw1UekVMSUJ0cLN756q5gnSABnGAxWb35elzHqiETssthLOITpsLX7bTNV6hMlh
l7NjZ7NY5Bj6QjXLfN2QlWPWpepRt774HBLmgg5ByuqBvGIB2zJ24o/zblQrnewb
dUsaKo6grA8PqHdEubCf6Fs8acsObTV78gPv34JPvqX71v6SJZlMVgK7TLXdArim
oaiMRnkQ/1XMKvhcQIqH35imeVxUdRNWp2CmOblCAQ32bwtXBvfSnrLr3i2qHCog
wG4zy2rvoc7v6cKQBaUs8ukNGH97FMg10+eGnHhEIMUxDYQD8ANW1sQUnR2jv3tK
0KWYerh4/4DRklxx/1/Z3/8+m+Cm8ERYgtztXjko1AMB6p70F/2WsvTvrYtk0eES
DaSqVDIAOzmz5S3mMZnfPBRIyo5/hlsR6YnV4nHP2OgQ35gKgARfvO4kdZXmQWEB
750yF2gAHRKqvVxoJ+pmQK+gc7ajiO/QdvJuVRVIWnDjn5IyY/Ytm0C6Bz2GVlun
yIsb/Anjx4koCmKH1wLi/598DPbptIWCPFXgpzpZyJGr6E7KbgPM50fANb+A0Yn1
wIZZOhQRfso3xwurWPVrVkBXGsxD1QjC+CLy/Zz2X3w7bxBX2wzNCuOVpAniDHLR
rjIzWbjVr4urV0dAywOcCwjiYAQ3MMpN2sraNgV5DgiuRh4kBmchE9dG4NIDiqGW
sukGmCgB1QCjyAKD1nERCUAYA8lRqoxB+SpzXMy76UTLMFJ8q7dTWn63cJ2lncl7
TnXTlL4ReQVixpleyGIZjGEIAHZABRXA8t7BHSbBTmzSB8P7ngCgeFFmWsfAZGhn
WQeMM1p3SMDSXat35bfp+6uQ2DygyoxaLAc4wC3/ZZ+5cMPbjn0OwO+aHaerhJfE
a4DT/q/Mzg8QEAZ6TjokjFcdfgk/JwTvWTfmlviXZYRbkVtjysQjmQRYNE6WEvJ7
NcaEDetq2YP+pDUUuFv1qy7Di+HAMubc7+pArCPyNNZHgT+r2vHgYVQAJ3gU3tF6
P9L+rK4sRC5D6m+xSoWy9tKfWEKXFB1s/P2zl95lEMkmy+3rfvVBuLnXK2dSEMTm
sh3cMnbmFCFGG01ZS/YHuXRpXgYdnAWQAqK2mDqqaC+XLLeZ+8k+Q0y/y47LGp3o
7kn+mZZzCJCAV5FsnJCwLjAHXazEBEGy++Ut8/K9VxAoruXQ2OGDZqE4fkqaqf8V
A+8CyE7/kjEIHIrRnVz4BzJ8ZBRyArmda6dyJV3ETAcXgknc/yReqJHrT8bhgLqh
bWYHcjDkLs9dmjEaKuprcEFentek8Pe2r52z0IsPkIT+FiMcPFO6ie2cO4HI9eJj
ugwf6xbYjfWppB0Ow0YvA+BP6tL8q0OE6OCgQ2PhYDwEQXQsIgwFvmubyI9dJO0S
qOKSrLiTUDIgxa3noiy444ZQJlzdlCqGCvm80OUzDgdow5/kLeRXppQ25rAmldK4
TNm+7qBJdnwVVlBLgJt1TZJQ56Evkrz5pqLY15OzMgn7mpBc5Cuy4FP7Rjy7jtzk
vErrVeMXVdvTqHpxGdqd876FPZlZPlUxWJP2bQU0zCZJEe/mnrCyQHN9CPIbnj0b
/V7XFBB0smv18OjQbVIvf1i631mUbzKvrSrCf0/nPVyKFVc0qd7Kea2TKrpbZXM/
mk+qRbQlma61sz67bzQxfKrQ4SScnFXU+9YWYwif3leMAgRzqzdt7feUfCeDTGFi
ft2mm83hcvQw9UlxSheSoRUNCaKy742IDHIoBLSbtpTzmjY1hvXgtIqkLpfLaWUI
zefhbVxD5CsH/8gRIRKOgyvGPLJYC2FCfQZu8/2fOSGOiKKXqPVGRiZEqsyAvcMb
osb9+24iM6tS9IOdZVsjoim8cCFFghbYDnEEx398uumKsVZMxVVuO80nDicG8yfu
jv/P+in16+sEhYIgO5A1T7oiqv36lAG+/B21n3W82c+h1XimNRuHYWFnzD3GzfRJ
p3FnCHhs2ygvvOvc6Tfk+0vDB0qwEbPbzfcpYo77iEe8GygM6G81hbr/ODJSY3cK
3KACU9+11YuJKogNqPI27q0RJG0vTiu2wBjqV125Ybys5ej7YY083UZO7fnqlXDg
VFORox6d8Fsv5tT2hdZ4TJP8hVnR5k65dROfa7opuh/rMD9yzdKzkbZ1NeZFhMNi
ViiY7iboyopFupHzHOjejcLCzgzGdNtVINYJ+jYtfO76s60ABhIe0pNpqDX5fmbQ
PzL4Ps/D5u+MaAnVRwZF3DmY0vHHMAnr3Hbzc4gy3plGkiBw4Bet1RKyPPvhfHt4
kSDrRsZ7jrmSgz41EK32yZ6a3CVbwIjWuNgm4z5DfsBrO9GbwRLqozirCdOJIgi8
NPAjDLwLv36i92j/lDp72YhicxtnOgLY14yxYYa48PwOtQt8Xsd4JKDdDEcqE3W9
20z1DNnh/JAFMir6zxP4NV1L4K/HO+D3nqDu2TxV1RnWS/u28RoK/bzxllfzoNs4
m3B1VWqLvLDDuYVApS5dsEXAZPLUN2YzYnhtuwMnTzOXywj1JmGjA6voft3Fk8DX
EnpbEObECoL/ZsAVPItrwSQ8RhlDx+GneOtacMMU3dY5tsiIpY/ufFR3rJjOjDOP
OvW9ENz88g57/nJ1Uhs4mzklJKuktT+5t51iojyYrHG+c6tsDUOAwBLpskirk2qo
Wuo6WeCPU2wRv/VT8yMaMec8WzpJkQCnLgB7cD5wMiHFlMn+6SGbv/1Gc6VEn5BH
knvmtpFBN9Pj4naXlwby03+k9cZkY5I1r38riLEit3+aqMtWqjS88oC1/jZfzF6q
9jPdABhy6rQgWyQ1cpMWb2fUVCkxZcxIlBzshD6i6CS7v5z8mAqTQgQyFn16N2B/
eHMYXBYTsQwKP0K7c/mXTi8pwaVDaCN/Xx5I7WHjLV5KMdifJzignv/7O7dAq5JQ
obPWE4SDIYSYh0E3vcTYhaQ00k2BiF8Q5g936yOFzwlRLWmQpCaf4CUc9f9olzDI
02ZOJaV6vk63NiurL6wQyJuNSEu04d21htGmfds0EvX8/+4hQuupAT7ClFy/I/t8
wBaNm47g3h0uw6I94WHWwufP71r8lLMxFmE4VVA20Ti5J2DC16wa8YYtR2Wl83xk
hh9DX9OWt4nt7tXMiY/qbBkPZwE16huV20/+jXHKTOrPUC3Qzbw1jdB5G9OGkofQ
LCKT2ei0N6WyBbzjqvrMB0K3GceiBU5ZRoOwHi/YqFexK0QpTo58ec1HJ1GQRU4x
vs1aN2aBUhClcPCI+sFANDQ3UmeE59I9m+A0xUqI9dD6tOsY9INUgaMK2EP+X/mD
zghzxKfU3YLKBJ7LRlKjqPR6eBvLRp2ktYpRSRcRFaIQzS4QMqJnJLceevM1Y+pt
Ff/LC6JDtPvZve1CfXLyU4lDRvt1WoUHXc6JVlupF50pdHPebRU5ys2NVC47vwRE
PHGQ6AZ22Z05Oe9MeUGAbeTIBib44qI+8kz297TeM+AzSRSRjz4h67N+Sf6bPt+8
v8p84CZnPoEcqCjPUMH/ht3aw3mGA8yrelKXP6U93MHDVbj5YEzrhwzewV3YTvpf
3Efr4J7xc7tRtHJlDiQn9IM4dOXjL0QVPq6AQ6i23yd7DJVjfgAaQ5mDwSQGx/Qf
XPh9wMeP0j1lc52xQU7O5w7M6s/ulAvDl3IQfe0aLTaGidZH0ZLJMUNXzD4nHAUa
1e0lDxglk6mMJX+TEXAlPqXCPREOLwyn5Tkcm+Udi0JwwAoaOlmlcLGzb1szD2p2
p/3zSvW0ygwkieRMv91YcT0BvvDsRfnx7DXhtt53y4f2+6UGHDty0duKoQwjKFxU
XIzFqviom2+dcYccLAcUHtyMCS4WLiwRFt42DjOb9k2UnwR27eIMoDef4P0WXVZb
Eswi9BBTBwmWQgdGZcR2u6C0Ovalldurq+8KdyEuak7nK59iiWpBfeax27mwZdK6
inif0eriedg8m0q3BErTKCofkl8xiB9f8cRREhAXAjnYUy7sn4nmR4SccnF/9Uxy
zP4lFtaSo1jou0eALUK9DjQE7jXlJ+TCLchPfptnok9UqLmq2IRwCpl2mcyBIsv7
tU5qbRIPaw021GoixSQ14vOIazButaJBvpejbtdscmhFGqZp2vcylgA51T0r5aEk
7zfJ/WIYsvAAh1g3+gIXnuoE/xWcI9NYh6ckJCT2V0q09Upp575yf2Qw6Ka7KxeQ
Ih15f3hG6WAYoicigWuuoGvcqZCD+TjapyZ9c6PdbDF3ig4V7HmPlfBLKzHXzOW+
lWGwdd/UpTax77ezAYWFIWlAYxxMRlz7uUqJb2tiTyqfqOKyjDZPHUpV7QF1CfyJ
SJ9+x1uXIyRs0hRysgslWQIbAMRTyxo4eun8n4AxS7KugkXZdAwhSNXF2//r2ytK
IO4iYl3a+5rOg/xnjmn9SEiYdIvVaBa8c2QWF3BCIIcks+YAUS4eQXDHU0QD6Ua9
I7i0JfmOizr2Jt/f6JP0/l4nC12izptJnWCfEXF/S/zT2g0pzawFqzpVPP685xR/
BZmkBfayu6jF/n1p/dZg5HUyzu7VvJNCCRYvVXIiVAH3tYFQwTkVUgsZQwt9LgmC
Zv/Q0p7FyTUfSQyb2xy1CHqnrQMQoMJYfTi8+AGXuxBPCu2+7RGnG5tI2fpzP5aH
+Mjfd9s/dGsOfElKO0Xgoc1DumMAsWR9C6Hj31I+5VLFdP3Qcc8KHmYp/DLNSHci
wBwEJE9ZleKdWHBqCaipvdtF4n8LWB1SvQN4sp4cYv2/XhtCwX8X7doeUpVnjVwB
8XNBi0W9BmcLRIAD1+Aw5eP2Tt1lV2SJLblkFsTQkborv3Jvg2ZY5dmLkuXAJ8e9
vWCDotWvzl5VAAaDuu46cYtjRJpMRN6KmL9LFwJ6lRqRV6EKQ2Ox4rUP2c7CJ8fL
8/N0tmvLbRQurQl+U8ohQ0wk8aZScS/F+lEACX4sbFl8dcBiyd364Qut+3SqYfmp
Lq9u7Yc0r5kujta3hemTxritPzm07RY5XOee4cNu10rxnz+sBO67XHJSvvzV5c5p
j425UkWMP/wyv6q5pX9om0T4OpahE4WwHpVxNgoK32QXkzK+0qFeG0XvjmZl1U4w
W0zUlh387Q+p6VnUGe9hbYHHge/IV3OBG8rZj8K6ExG3b3WpayQgkpPHhOMIfIuT
V8NPouG80WQMvNXrYNqQKWSAPvUGZy5PrAq/wOi6z0ZEhbe94oSgSyor9PDskSRV
uZyD/LhQkY4j6pzACg8Cyk3aDLr81u3pe9fMd4r93ZRiZZWQJG1S4vtd7W993OAZ
gErL0nWEBjUwBXtHE6Gr1/noyXn3A4D0qOUKgxw6U0F5FqJ+h3r7lDGkIKF4Mqk9
dHkEdYWc+rD/nuGGUkuD7GxwdJV1/xgdiEg41aVaEE08LgvOVwpYlF31qUcyKroh
XSkYfsTexLFXZzyLyn8pKqzfqVN60iDKLs9snnAId72oYqIdNeDmbe/NGBsi1o1N
6b0V+elnicOyVYpPIyP/f3MShCGwbjHPu5FF/IMLdmWgXqyrf7c+r31fyByO9cZU
UfcJE41edU7uyX+Ij55KMa0pW7gw1oBb/MMHDSrDAVbREjrvZ3g2PBHyYLkqlYZi
6EL0pW8kEtlkbJmgHeuoBg==
`pragma protect end_protected
