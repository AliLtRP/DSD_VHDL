// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:56 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
QrRg7oErSqdRBZ8TzPwDyoauO8fFgn1+kdADDKD01S7Qgay6jVXXFu4Dc72AFNF3
LDCQ3pk5x2mYj0yjqIFksEvsCyLpU5M/CZ5s85XhaSf519c3zFC1x9voxvivLPBZ
0wfyy6j9XwWL44sRk3Fd0hwWauHqyThLj9mPr1AlYjI=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 11968)
KYmy4G82rMSNTuweZr3pyaH5eeqr+IrvOwb0cLcDRNxz4Kmdy/cPyWcFtFKww0jm
pO+lvoxpDuO4EJbbCPMPCc+6WkptHczSnefe6hVw6HCREbHieZbfKXOUUe+BjV+Y
yBnRRAqRkrB9E8+aIw7uz2Gs5McUegTGeBTL1nDFCL7XVXnt7b+JC1NpJ1qWdlQK
RU/UxjleBniNWF7kuvVY4aVedHex5ow8xbhIPxUZfJFF4s9diaBT6IW97aNHVdVw
KeP5kTOzem5vLUAqCx4ov0x1NLgp7h6U6gK/FSD0SFmw9kITG6V54LHXE2BkO5t/
UJZHkoMsRq3MPkvwM0BzcUf2f+VmD4SUmRAzAz0w6bk+pT5YyshO7Tf5T4sMBieM
IjpCFznejemwL7FEjNOJNCeArhHAqaU2KoxktCaYS8cmDE/HW4stBc5Qtgg0zGT4
mQw7BdYpjdTkj9yqoT+tYuGGhpYSOO7wqnKL7WRinlxYbNfTc5SDtYJ4QDVL8GfI
hjTI/Ye4V3Q0cpk62eMhsPJHOWlaTLS3o4gBbHcUyhZaPRhk3sD4NGca7EnKFyYK
qBpMK/bLrO0g70GVD7w5T4rZjA2uDujgOPM/cAdnd/eh+jtZtME4Qaj/IB+rHhzp
6aK04/klyJ6bxoDn+xM9ijrNztj1exjTcZdEjYNOM5upS7N4oImqoebakXoEr5V0
+yRFSDPFZsRIGzzF6jnkFEp7H3arpa3H5bu6vrujeqjVLg98jqPi8WDXm3GNVPWZ
ZdnOZaqFrIj1EzDhS1VI1Ns6Hay+HovcvEMx5Px829aC8opvtUDOOkZc6imkwIYK
ZFa3xu0RwibzCW2gkR3miVFHATYg7kru7L4FvavjncmPauPm/ej2oj/ztCqd3WZH
sUbKH3XQITG6a+/qFirpgOB4imouENKqkvkRNbPgFTK4Fgf58IaVEQVkLirP9PtA
UrLwfbSzCFYUNdgCL3NQyTnguk6GSAGMch/53X1xVbqBDd5mqt4HKAjjaBSt2KSf
6W/m83IPw/RgVqLR3wsGfGTBr8Y8CUfEdlKjW9Pgh53BC5lbvLEQQMMnMcvUpsny
H8XEUYdRVpzFCV66KjOCRR7JSr4HEJQkxnGx8d5PyH+KxZ85108CZvtUj9XFt40w
uD1PYdXihybi+Es2C3P6eR7MlMIPbV5mv27C6nVp9HDLa5pGCxO96MKXnygO7yxp
wezsX0fXigaAsbbS0c18SztFNwHKA5rHFYtOm57y0BG4r0dTL7DI596bHHLLKNvl
UErCg44+O+bgueu0oiLETlpmkj8XXooLzQHfRuY4pU/t5y3IParb4Xe1ij5zdjXs
2K7KBG965LBCYyBR/rX0eZowj53v5p0OMAYEs+rlKpmu/9BE2SrzhD39XI/Ai/Uo
MW/k0z3QslYYa7qxw14zYOGQltlLEc9YqxppiQN+7PQDcGtY+AKGxO3EFaIwGn7P
3HSChV6D+9a25afBXvXcsdvE9AgetutVdBE8QK5scwkvhMeOBZDPQ2PRM6H5UXlf
dc6G/dmfZfC7mpdBXE1fzw84T35W50/YEVDAPVl8ZJ5B6/kfLW4DrHL/BEwQUWYs
onPTq6He6MLpu8nvgCfM+aUg8Y8xbgJHtmRimvnk+YWZLKiDxybcMVkwz3MkVJvQ
gk/PI5vE05zeJZrwTI16KCXJk+pCgVhzRoftNoR6Hed+hovz0VVay/axd6oqahwQ
F0qYCG4naKayA+1AyIb5C1dghZ1jmqRKVBzM5UtdlnmjPslp/9v8RIDF/oypTmBu
46ocNwaxUggsu7Qa2tuVm62itJI/JfYoYplXRYmMTuEkG4KXJ2qdQCMR0oNk4dML
wvZNABkVIGAATtevvp4ECxv7aGJjAGUAQokfFbip0yd4EMP6RfqzoXbv/MrwjXZ5
ZphYCvXNaBmYJbkTJt69fISJ672QxfKmlCV5G58J6n+vQNaEO4LR9JfoBFN5ypKf
qBKBAvSJHoZ+M0T6AmGrgEFWMu1TQEVRi4gw+8mdxy8prpj7MW9W2jq7u2i9bNBj
abvD3TjGvgbjI95HHFxGc2SIW/PjO5iEhsFt0oG9LvbpDh8GVBJ1FFWY1iHJXOqQ
F4gza2ld2IMHXOr07Sk5xGOlF3AVDZOhEBRa6NPcErjV3QZ/ZRsM+upINwCYBfuv
HX2LeW81EJ/2Qpr6a7CDGMund40fARTDL3HDXb1Jozg+z3R8IjZr838kKTucTpXH
Qs3jy163wYwjoYEDtktc7vvUu/wcwlZVVYy8hNwyZESaSYcavTLCsgZSxbK5aIJ8
cex3XSBG28VUenGfreqitTvzny1J3+pqCvScigF+isiAN0VbpwnOBmxzO2/HdYjq
7n0arInRvStjevUHxjfuNPsyKA27sViEnZHQEHIuSUThwey0IBzKtL932PZpouBI
bDUVxVCzLOVcF8ayW93UbI6KdjBqjYrDIE8iB+N7k+2YvomccraHbzD6k7zp8uPx
HmCxZz2j4D+e0Wy1PySvTsvoFoBveuKgdQ1t1WmyoV3r0/dmLMq1l9BPaXPgtrqK
GYn3ACkB4BmTFzgK8P9nxBKYWv7GnUySmLeY25aQ8jGLCj6vflosNC6Gx9CFMKhU
z5O2FGcDeQwuCuD2WyuSIrBM1fwuDMYy6AoGr20Bdd6bWC76T9raDuxJxLhkyRhw
XvI3/OMfRf2DP1PeICZBLd+XR+/uIsZPvdWt0gfpggnG9F/VJfNm1iDaSivLvQ38
spMXi0WC7ArRZySlxIWUxO1ZxTADcgEZ9f8FKaWxIhBrzUFU1v5KpVw3cq2bL1qp
PJS0faCGIkKhm0Ik3B2d/mziedxrWQVATp9naavWP0iFzJU8ROib0TE1gmc9Houx
JkEwYXiHOg0ELpx7ra0FKx9ZHYVf6/UH5yMee3sNcpJVoycYoiOpgMxlWSXE9S0s
fuRMdxBQtbupbGsyM6YPGOKdIXoK0XC7bHwkKo49YRE8W4U30smCeIZuJK2aKnA8
qB+sjkpo/fUeTjfNTwfHaIjha5gjLs2Z4z1VYm5emZttXoazBfJfCz6SEcYqrfgp
oJqNo22WzB0WJSFnTXjSCRNdAROHYRVPjiLckgEBQoSp1SrAdvI9haXO9wDPSNFh
mjTNpyFMUoYCFm7/Ijg2fCgKVEqH0w3NTQZjtVGwwyqUOaubRNh1n36gl9OYzpN0
JxhEW4fMd0/gCOsL3nkQiwgp9auDYPmM+tYdq66iVN3pgRZy34vQ8aTH+4YGY397
v13QzWQU4+dM0vhvBnUzO2js3DGh4ikDkR8THBHLFthGxrEULo6aKGmH5XAA/IUS
n2h9QeQd6vH2c/lgNWcfTL0j4W1hzytAmrq+gmqBHM2m8fq7rwb4zPSnpvubBLbB
UDTj0wpxLjf2nO630DgiXB5D33NpA3GgP2lUu1MF9dM5cbLkcdLcXKO0u9rtFoLz
Q5IWeq3qkY3mXuKjsCTZTCKUSs02ThyH/LwniSNCFuKmyyZZ42Esy3hx9BpuKs5M
Oad/wpuZCnkLyLhCSmmQplgzt+2treHH8dAthsoHkdxM94uMOY2A8hTabLmKXxAg
PzO0TSBRWFkdLfE2b9TyOu+B8LMKcGRC3ELj1rPWThkiLLYiNFjvwo93Y9gx0/Kb
1AgQ4D41izeFHqq8qCTfQadlN966A1lyajWmWEv5Ac1ugX93Ax/UXUN+FJ13N9eK
bkgHipKOLzJTb8myn/ixPMaCPGywJatRaSq8wFo06UAxoV4cFcL8DU/RxzONjOvg
SSam7WOGblH6W7QxlEKYpgHBSsila2mba0PaAK8DzE20XAjCnCmpGlC83ay8u6TD
UyMQCIXMFpz7dc1BFyCAN9ouveY/kLef2BKDCRephfzX85YhZgjW9HjkC1s8+Vr5
w+y9fssQhW4vtaceOOZ/2oFAv69xnERh31ojG0xC6W6AxNoi6XWGnrt09/ikjT06
Ky4wAjII8kv5/XfYO0HvZaADJJUwtQTyuX6Owo3aWllZhBUSxS4s0eRrH7CxgYn8
1n0a26KoG8dr6OI7r34th4AvhtPHlxUYmEvzgG2cx9j8ukwfwveZVtg0iZlC2hup
ygtWgwtYOsiP1sJmf4jroKKKCJNXp7dXq+gVuzl2OYbNlB3ua1aj0gfpmK6O81Tb
2qYgzUrtav86cO9m0QAzV6A9dY3Ui55IzFA7vPZNCGo9bTEzciAFEjclq4cQ8+RZ
FGcYomLTSYNushDUgJQe5McFInCTdkxiowoTg8FkC6tkkk3U3d8zU/OzUZaqqFFB
Nh+ypyQgYpxFQZnRZdbpiLAeCLedvz5IqoGmo3YsBjK9DDoX+Zn/pRfWn21qJvQ6
ZTDTTvYzCIGP338iqVg7fImjdtkKp9ESafE4uOyvIlsJB2HmBrymhaN/sMsjYpAE
LwsqE8fqOj/53aHykFYK9DXPYqe6Aavm+uUqb+c47+D/PctIUGET5Hq0QS1znG4g
BqWW7W+R8/R0KXOvIsZDk8Vt0cL2bhxLoTdH8+b8JvBjoH898qSX6lCIlhV0Qyai
tPpjvNQaci8YH3S+lq63OZJHAUqWJSCJxpEO6B4Bx6YGU85Van+0nuJTfaM9ypY3
9Pk9n1IjRbn+GsTbhoFaLt1K4w3VUbjg4jpRI8RHDUquLW6xXhz5jFLvIeLAQpew
bzsuYo1qOcvawbXAVUYmNuNf2lafMH2Niitpqta03AqejHRPkYvVBaa9C2gF03Dv
yifEbAq6ZhGUTWNtd4VRsyV9gKNwm55cNvbcmw4vY0pWmmX0bdyeqClnE4W0nQS6
a9TD0XXt41LLsRLP0VNivvbKvHQwjnfKcOVDaTLhvHLb2jfIl1g0GgrOzM17TaIM
iB69g0oTl8zVQJ85GqvXDjE6NBcv7N0WG0+Eq90wUCYluBzQMBHWoyn0K75nn4Dw
6oQU39YNBW+PO+k5SJT7VB/8DzXpBPk53aFthCaSF2JAS8+Sjn21NMte4MuxkAKX
BBEoZUuhyFpJ9OxTpVSEbSoiGeNGC6cWQuCpkIS1lKdQzhY7Bxl1MJunTuuDyW7I
FE9HlousdI/ybl8U52EIS0nKwKYCh7hlSns/zewH1ztMfewz6fi5vtDtBPwpfOWv
0aBY2k26Uc/5FL3gYXivOUP6UMm4Pw1xPpLFwJkKBtWnGmILy/jCNp+DmtQxej3K
n2Rz0GLz4vGRWRASuzvw/sy+IRqgI/Ct9y6+fIliiFznY4ODhbk7U8Q41lIeFCMb
CS8vVqdt/c17RoGrE0e83Aoblyjl/1DkrpIP7l3E/XRfFsKr8qITJAz6eLgDK3fc
Mlp30nDcz/f+0+ZBAAJsnM+lXXjf5t9R6e2q6LFguWKG3L5IvKZGlMPSHUltVWKe
DwW7shnsB9ebXNnZXFen2JDcQI8MvfT+refXlXuyDx3BfP9fUHEhlKg8ZDGA/TbU
crH6CMwbleOBMvtIG5//lruWeNukWZKbaASKhxpzrXYGRFl1jyx+scrrtqkCJAIb
i3auUjpkTvfilNhkenkRoe7t3/f9QR4qznxcmoW3uEeHqFuI24aT2M+3JHiBJt4j
47XwDp1Ihee6emjtBNg0l2cf/7mi5U2+A80XlgLVp90+8afiVph/ltbVsqJagWG4
QoqvNaNluHzM95Z8FyxaCh0ykTusdEriUaHlVt2NB01dIYiti5sPvperUpeT40sK
X7brnkLtW7rbRTnY6qpCChdUkvVhyGi8tdWkVSzWy4xbK9vTK27ti88ygJtRs34k
YYSVR/qlvV19O6cTxrZ6rRCuQHBfqWp4lyH0EOLMJAx/KaTp/xiH6sqMFyXk84YN
z9OGP0ixA9GK+1+qlbzFK29turpk60i3zvkYN2JSvKiFBMtZFPeggMUyGEszsdir
hiTa61D9lvjk5nZrIpCS0a4hRGkkGK1lTj9dAsNOMUpYwzulQZySTzo6vHM3PNOY
o3InyEf1PMnHzBKyT0DbqLrKlZsa3oECrmjUgu2nmGL8+nMvVuFiuquNlpvYdjOI
OpiC22cl6VWkT4kVfKfJ5SHZujYi4pvccdm8y3CwH+GKZr6yYpoqNDAIHWSO//LM
fPI9BunrM0Ed3z7V6mSj8ubxisHs/s767dasDKrXsTz8eTIKRP8D78Y5I+wseQ6a
Fzv3w3gdBVtlie28qrBSBK/dLqSQZ0YSgojQ7sst1cBT22hZZqdqWQ9xhicHwQnQ
rMNFgQ4KSr021phj64aBMCUgvAOmVYP4dr5neNBWh6DZDGuq0Beu+zk2BCVKZmfo
iuIY8P3EAqLwc8ixgBO6TDSG53VASTjJRF96o65MD20YpgDAW4lIcIPrMyvd/sjn
xJl3mOWc1yUJXC4q884io2GxFx/L6exTaf23jI6n5VHEbgFR9A04EmTlNagZ+0Js
UsShJ0ngc4B12NIKudwDvobVQVQee9VambhGfpkrsLzOl0eRkqq1AWxFMoeBFGfV
/WuyLxk4lCVPjhV8YGCecPuY6KIMlNh1BVQKpHLUpeFk7O7chhlII4sfXIDEUBW+
ugiTHuYQ8gV6t8btU+66wfJPvhvDHJcYIDczW2uiikDt8g2ZSmAhsXeG+DIRwb9Z
Zgx72wEwVdeZUUF/9oCjP1Ya24oOzV84LHDvOmOyMXC2Upk5b0qd4cBFlsA9+32L
RYnXHCsEmt3vME+WZOM2PiX7csQXsD3u5j0MDtpsYwBWzV/zzg5R3aNyXZPw57Wh
j43ZmyjCwCRIWH4nW7JOFI2s+yoKxFCPBUktxG840OhJCV/+35WQO1uVCJykCoSe
7/ufCBEdLIJ4K143Yb+hZ153THFDz6jRmwqy5bEGILyhBOxtMUhN4PP0eEZi4U26
PsNMdcO4qemp+h1diKyExHd4jD5bDohG1eu5oet9iw4ecAx4ufHzpW5RSHR76fqF
wJocz9kuo6WJGy8Y3fVnpMrz+YLaSFhYFPmD+K3ub8wRgr+cN1Mhjs803FeMqVgM
7IQ9bbSlrjlInP8PeLhHaTfbWjwk6+uBuSD4FGKzF8nT7au1q9dFxTrL3B7swEaT
ScTeWdgBhlYhN1DkdmoQ/alzqalOfAZSaItD6rJxB+gpO30tQC3ZjoI1Uk2om6lc
nbyIZgS0c2iv2QcFEzHfRmeRL7bcVwwmc/EDeQ2FP8FZWjLRs3o8USHD24vivo69
WSC4jD7gT1Hv1LK/fneVni64KiG2WQ+LEvTE/MmUKwkqgXR03Lo18EbjV0zdj3Kl
SBnMzrn7CRjm0VBVq7h4j1pBsy/XMRZ1XxuoiAfD0ZqaZKsIzsY9DdfxJwjvnXIz
VpPEv10/CsgMqTKLWlweNCsxIQR4u+BGL/7ExGmPUc6nvlNON92v37Qw15Wq04Ky
7xLMBsU86Z3KwLQubaFGDb8WjbqqnHTkN6ldVUsQ0kbYhKZjS8kSzoc9ggMrEm2m
l8rIrJ4dChGxSuUQSdN/YcC9QZDSflfd3WgG1/v0t+D6miW8ofB3V9qYMs0KwvwX
mMH7oA7RsJxIDcFox+0MA1ACBWRi2H8icX0mETqKb9dpaDf7O+xvJA8IooLra1JF
N4Kvh+6PwALJq10GrquxEdUxkMMKh+xFqGFuYEMOnBwe86Co+pAI01Ga4nPbgLSP
Zh9pFrJR2elqGMUSsrh1A2KldNZlvvP8BmPypbYpzyrGVkuMtsLnVfnnN+ApFIej
vdumprAAL15J5gYWgI3+Tc0WfeS22iocdQabiPkGvsN5QvNCLj1SSHWnMgtQSzYA
SlDxq9Y2AVAREdR3XtQekT6p38iJ5OswSMy+kn/vhUulAw7zjfUGn8zgk6SGYqXB
xXFPEY5mY4ArFi/m0P9T4SGGe9aSWqXlMx16FHSdHKwSAakjchYiHAY+acii5Z8m
q3yOwTdPZssL7hi+vR1ki+rY5gYpwGOJGdoEl0JplLy/ZjAdfDfUc80Rk2Rld6l/
TTRO60wnKDxi0WOxlhvXpowEroHYdKafS3ocw2ir/xXAC/4W+Z6E+4t7qwxLl6IT
1rltqkemvyjJBKYyWYYNIGFkL/smO7SeFn2vF6ySvDGr6ysaXlqmeyw7BadZd10c
+FdIJ2fjKgtZKm9gN83oK4Z9QxtJ4LpesNgk+8fj5W/wbblAbhA+pfrgoha8WbFS
AQYlJNNTtAhNUSpO4vRsFhuvBy2WVe4cp0x5sM9jGldUTkAhdPIE1FIBKXgUg5ZC
rlciKPGySvBkjDkwfYskmCuOG21J3+lhG7FAiL1Mde/H2sw9c1GDxwqOFuEOGnq3
Eugz7tEjAQG2z6HpxuFs+xfoPiTwner/LcQ6YompaA7QULg1nn3z0yqmzWrwnYXA
0E5SpkBhSa2BCfT/IogoyX6cuxRaEokDl0nV+9GGbTEa9fQOybIZlM8kAoVKemjd
ImQO1lsOJAlqQzTMKlH679yJPCuNItAtbpspVUTeUCu6i6uDl5FfJEwe912IQNmz
9j1OoSXv1nytEbkYIxpReHDMQuzyeQwGhcOtg1+zLzt4QmchPdqm4sVQ6FwFqGq4
T7PrkZPa2256mk/xPJ8+oyP9qoAWJHYFFLUI4wC5iNGZc2fbdeNDeRPjdiIZcI81
3fMSq2kucq+U2ZJyMWy7CIctbD5aiFU43hYiaf046T0TfSOUp4/iHChHg5QFu7mi
0dkdrUd0atTPEWuY+f+NM10kpPdaxQyqNQbghtSDlKGXtqxZBRrdW2B70RkIMY4u
uPCX8LbOv9qyp+iHeAxRz6wrUByMCUZ97aTZ1pz/lVd/rpk4DTZT8Ffq84p08Fh9
eVbxQWq7zchb6RlCMOSE8vXkQptAPE9kp6tF9GT5A5rHL3ac5WabI9mvH9bJ08Rq
B4bswsEA5hpYxe6LCgP9E01wYxBYq1Qmwx6E9tqPBMdieBXqvGP5tB1dWu7EW6kB
hL1FxUAaUQDhnTQEZ08KY7BDP10qFc4d8iq/hwbWogq825ssO5qiEAPLdb3h5yAv
jwQVV6zoDBA/nKRZHvebFm8tf+6yHyI7Rc6rJ8aKNDKkLa5T7v8CT/O5Bvb9BVHb
KEkbzyysiB97iGq1E9k5S7Sskr8tkWfffOTaoLqW6cjhb7kUMkxSI+O6LIpw/N5/
j01GBedZq6Tn1+HcC4hnFNK2BAGjCLVvmB8DjBSmmk5GJv8yQrvKzVPN9bo666ao
ZIcNchO2rxwwRVrF/6093ljgqaX1TfKWwP2ANqNs4wLX101lyXAdjVZ7wLsoYANO
FZVARzcV1xrXIVFmysqaSpdRGcVMj3utmuYc4/Min4m1dWNPQvwirdJZptI0QSdI
TTnUaHf621/KUB1pRX+jiE+AQcGzaey7S5WpGT/QSHXmx+kYgVVN4zLrMOLZvVaC
TCVuAbPBKzA6D+cVLPLfrAVbAqLBMPSkDRuTsEh2FMuUsJh2yGjsxt6B1xtLkXda
ng6YzsTWP4lPkGYAeESMkAmsy42Y78M2ddQZZD3c+tl6O/Xemv5nX75VkP1nZeoI
v5A/egmXO3r2x5dE3Ytr7RSrtWPuNs/j1ZfN9IracpqXvRc5on8RiV3csVwSeTm+
Hawl0ub7k/La0GKpBAn8JUMrDFIo8/ZqEkJPB3/o4mu+/4ywISimIlI1pQSSK5s0
NbPpxqvi4keUahU37K9HZC5HVoX3onJVgyBduCO17EkedzKZv8+Ndx0KYuYJCxuh
m9ePqQ63W7Iw8lPUyEbidXDryk0C2WR/7d6ZkROwMBa3JOI0BujbMeGsTrPltnzD
+qgzH2bHBVswhtA8Vpin9T/SHN6aNd7/tm4gH1Llecmfbe97Z2Ht6AFha2XCcos7
rUJyvLtnufsVnGY0IMIAhFaN8CAxTq/vT/0aTJK3RW+uRh5TDvVg24jIT6LSWl27
xMoo5VQQGj1QdUfn9Ho/K6jpswzUjb/Q7bbLD0LEhM8DMKa9xfHBLIsUvvi+HZ85
07WOYiebQCICwDsg5Q7uh/FMpvAbU/JlqkL4T7FRBL1X+eBCFO8Rm4X3tfaN4/CK
VEmNyltBi3AOyc4gBjVawgiPje8IgYuNsSZmp+OXy91BIdj9GyOHNGfFnpmsJDJZ
eVzB6RBVk9TlYOZ+G7mJK7pwVms7JXlpQ4PWHo62Qy8kLkdrPCMBvR4JPh08ej1k
PPxTgFr+gP1hRoAXtLe/2/ObgQfftG2kmDQCOKfzYuqZprkclPgpwXPMGRcv97CU
fHDhThXeNrHoug22BUCHCz3hfFqB3rHUkWAc2m79lCGSeJ1Gttq7h+v+aIh0uh5H
4x/C/EoU6LKTdcgUifTu39g5ZNPSy28H9QEL/LJtNEpDnAJ+2gz4Zo6zQZYmNcTs
DzAq0kUy4werVsiEz8amFwkeIX0ReReEq0UdLpvhun99Uw7CxLymrEoZgn6j8eQe
Lsvj+1tVEsbJFOHGlaghWTYznfhY6qN8ugKRPSktyIVeVJ2XNTT9afC2Ne5qErJ7
90pk9r4DTrUtYP5RGrCrhRd7tx0tudw944YN3O6Ef058gIGmPqXIcJD9cAPVgFUb
nrVGhPkKimPuXr8prRz+VmaRsvQciDDgp8XX0WWrrDQFMo0l/JGzwtIipYnEP7OP
izmPk3sVCivDl6Af9vmB10kfCnkwnd4B/zvFrjmhjUGcXyuRbEmG3tlU0OP9xSRn
wJwLpZ3K3qeh7b/HcX/ltBpTZKJJrdbd3+nP2u9dfoRFGbTomi68gEKC+ZWa4kei
mvPrptuznPns/J5fNDIYw5GvgMZYaQfdDw1NjX2NqlyFT4g5gLFDCn32ZgrqvbXA
O0jxxRNZrS0p1RazKX0IjsK/jBrstvC7qU2l0AhbtDFWOCsIPCGDEzpL+BaNWv4h
wYnmUQpk65wYrD2nGtgnfcgsoeLfGVJsG+FSqUvAJLaXipoTtGxiqt+zskC9bufC
C7mPLs5PYUxjctgnxHwSbMAvi3pWwgK7V/dQkSpOO/p1ldnNSeaIDcF0X+ocVHLV
Qno5W1AC7uikatxwPQp4WsvcKvvYd01TmV3AN4ymavA5eqEQd0xSfs+ipn/W63xk
CAHeG0gkQF2cBVVmWxwm1uHZ0AOWm8QdM2xvM6Okm65AjtVnmNcj2b90AdphwG+b
18fqDE7FBgkO+kMvqek+lvtkUAtIkPTroJY2QMio7LP7W+0dcTnYR1mIe4Z/APNl
p+zxpru41vbLp/stYeab1ahABggsIaQhoOT7E6m3EaBXiw+7Dvmb2SsI7ktA1CAs
3F0bBCdzvuLCGU14NZHar4mqb0jPkpDlrW1ANF124EL5so5ezYhFy5graGfvhDgX
QE/8OVUtbS95QuUfj1QN3jnV/Lcr3W0IfhD+Su75i4T14/cpQaoaOG4F1wTazqOb
ZO1dJgZWFOAscW3xjR2W7dWRyUh5EkgxaMKdM8p+/VdDmjr+tFsDHa4Pqyj0AhKQ
Dv59Upe+wePnAmqBu9JJDIjhkkUgFR2nT52MX4LeEBan9ocS/Evra0YGDM7zy7C8
5iw0aoZpkJ+Wrri55bv+GoovJDzAAXoMO4eq1Ovbpl7qINe5xBOkwcCguJTzE0La
bSMhOSPQmyEuUAahg/zoqb8J1lWn537HZlaokkT87QssqeYQwRWkHRy4QNZ+DgcG
3n7nUsX27D3e9AsYGWKwXXqvroCSyrtko9QYMGV8a+ZnF1fB3VfVC6gCq5lRJnWD
4UAZdTvWzkb4SIJWJnba3H8apE+lc2oPEFnBihRLpqVjxol6isnyhjlJcmSdmFza
cglhx5oMpv3TGdcl200AZOe6sFvW8QcrnffmvskATJz45DWqGydBvB4lVgGXFFxF
bD66D8pCX5aUtzjVu9HEUvR172soNheQk2GBRmO2Z4OFyYbApUOLsgYRcuqOGaSc
3FkUCzR+RjPkqmxrABr9iHuCHHsGwRwDeu4S6fsuURsfRdPk/fpJSqKgHhsNlAzt
+kGnbFDAtTggJjVG+T51atirljWxpc/oZEFo841mScLaWbj/JfaIAJV34QAGr7a6
peZEatxAb4GwJedKudLW7LTdE+Ob/ORjxzzJ2zVoiiVfb/a313GjWnPUGSxmwxDW
t+a5xxTc/0L/BydQA0FOvcM9y8/4hdJVWGvWWfH7H+D0e/8QJ6SKy9VN0YwB/Fku
L2SkQGuk1uTfpH2yfM2BbZkd0VVk6cFYZqN6OUAGwHM/4dYbvN3u0uKgQVspzcdP
SNj6UBk3cJUXQninJQR1DFDigZUG8YDs1n1HSmVbbpBEK3ZGSoMGQbvA7atCDX5r
ZHxHC/aFgIBPkyF+qPuVHAa7uYT6ePLG8RmdB34hCQ+ugvAo2egtPv7MUGzK7aaX
m3qbx5m3+lt+7HnbQCvhU/v7ynNKCYV6KRuPfmOdI0gO9QwUSLyF6C2485szzDjz
VZgyJODOKDjNP4sYG8viPjixTcrYlJKB8XF8UuISP0uawIyyDumlwEWn4D5zVUAV
oC5U8Gqpa62qL658HQ5+QnT7V3COva9Utfwjra1zBjBltC4iQmWBwIvVoNzaD0g6
nHjxP5sObXpHaNo7NqqjZtnkZbR5GPQVc9RtHXttNwG1/TXldzCwgIN3I2f0ThZU
ISZCQlUJThcswg3YUWwHrZaAXtAfLyKhqNzYFw5cuSiaTAHB5u3Gs5Wjdakpjars
MSzarKMNgSxZsSVw4rHOQT+bHx0ouL1Lj+JFMZDxwbyP8qLSI24DrFBzadqRuoQJ
1VldzZGeRrRyWwIsysI3OhJeE+pBiPbzDWhBMFSMuCCHgbfGj8+O8chFERRKTB/J
xl1uxwo2PJoo4jbM2DcOIL7R/D21j2YVHKMBVVvvuHUfuv+EfHzxfbw61oC1XJGL
fnjNCgtigB3WzDl81XeSYQISrhhw5l1MKBZj6cFhPiddb+mcWU2yPdrHEgLVjNdH
AXlc4jGFj+uOlAuOSaOvk73ZH5Fzqo2wNfT91HbpCQuMuvjtGiwVKIe86fszhQPP
ZAi/7uxx2HQ2rqSVYUSJWamGencPFQDmXiArUOsEyQrbnsD2zG+P5+iONyYa1SDJ
D4BrGG6tDvQniTdLK8qyvUk9miS8eCDL9QMwlQGLYC5ccVUpp0Z9Sl3QDF3M2Q39
00lKuoV+xNeFC7Kd5ISOWcR1Un76NlCoH6AE9vlPCdrj7U6zHpfBDf+NFHBdqnTr
kZ1ujPEccC4YAm7CqTgBRuH9Jgc6u0bJf9ru/Y6+b6X3tQqC0bBaOaoGHyxCWiVw
OogXnd79EQpIaSNXFMA5WGIYnFwD1uHNQFjJCkAe0jVHxJojNfcZ4k8Uas/H9L3p
9/F2TN2odTqLaU4aQ6tkpKzg6Xfy2GWtxO1kEfhwnrqXy+WmtTpF0KW5mTyveLiN
qWlpU3+TCfmhnXDIMZ2oDUxlECDIU+kKxm+A/1N3wIzUnXzKhGM67VI4hluli8jE
E2g/csGlaN4Py4TCOjGQQLBbKEOwqO6NkVfWinVE4DhZTR464zWfJH08Ss2J6zA1
HtdvZKHmR+z5TEZFt48Ri8AUWbReKK4yQjQ9mIDbczTvzhTE6awM0LFBgRVsun6A
kTaI+J++FK3LRZdtaJFemv+fBio0T8zP/DH3s0s1mU+B+PC0UQLM106JUGuPVyu6
/atzG/2wXcH7FUWzmARJJkOXuP5c39PlhNr/xRYnvYxqWppHcUqsLXfTMR63nn7H
KF9iVQtVMzTGyynVcFcDiEZNphABczPgtyLhXu3YzhjyziDg/G223eMJEun695TR
Y/GimVsclMCGfYHJOna8VPVTj8MvCvYyKMKhmPY0UoOgRo/hboRR0fLcPhH+VMSm
aADXA/Av+7jwpz3Y9Rp3UL/JpXkklC/tA7ANGPbdwknikCE6o3fWzifirHSrWEIW
bRaOq0s51L2xfIiy4QZJj8+uM/lkM8eoqmacPgwqcpJnXEaiGQ6Nz6L8RJu0Erdk
JEcs+LEQJJg6JaEWTvLS7wg7PBlxdqAjjXZ2t8tBvMJM9N1HTTeF77/69SNcNfOA
BwL96t7Qrm4UcRm4BWMDJvGqTxDi3mUfXWiHpLa/JCYN1y6TyE8Ieuw0XOtSwEHY
lZOfUXYX6a+WrXhwlW8B5FrpOgnYMResNF7ovNo1IXZFGnPTC/+Cwcp1WvhXnlso
Z2aNmcCvrUF6ySkkmS+kb1q1oeYuoLBaWO4rzLI6HXQaRAH0lBZ6WRBujSq29OnJ
jSXAWW1o3f7BxIV8hJZIQGmt+e/eqrGoULL16l2YrVWHxWXcGCi/JxtqNNJ3xnFW
XDxu7y+/eyaojv8X9FU/Wq0vCttkJ3x3rm9b4gVQ4p0X51DH7vjWN19bA2bxfL9W
bKntDFy4vTYQCnoZoR9ce7zGqiLi7gD1XsWUbJeIMVEY9dGy51f43brbnEIZq6AW
e61mdwirM+nCnHtiQD44Pa6rnuHnpWjGuRUz6QFT2Kd9s6lnYF7C5le2qt/T9zuG
ucRXJAnhbk6U9GU99AW+/Ew974cnlPDhD7BaailB3rITorBtj9w8rXUhjd3EMK8R
T5lu4dR6HdzS/LCO+2gJG2lFA0/zp1zi6WZPavBzd8QNdjlBLFXNzuMcun2d/dB9
teLa41tmp5Y3Y4vek8atVe3e6P9QZ4TYMeqWA14NfFSgV7YF99137DW9sdN8GljH
jfxhSVvuA/A0PKiF9hZC+nOYFrYjh32K/MCpW4a5lbSPUeKV4YJOBalNIcmKxkpl
MgjfmBCB1vGAcgc+x6WA+WDQSNOzNrs7xzbMFzDd0eZRmLtixbeTGm6pA0+hg1uJ
LsPoqYEPqFoIOdzRoT+u/xnrYeVPMjRay5YQsM/P59voLxJQPb0Uv1cO6gWgWtVf
EHMgcMcV2cJ2g67Qu85179KoDqhtSPcPQasBrLXF+TOzWSRFAb3Zo5hexj0esvhO
TIsOfF7GBBeKQTcB85DBgSwB/w89UzH+Hfmw764WYp2+cMguE3le4VavVSrN0ZOS
BEUAuBSM3JKVtlPsm3QbCFncxyYqDaQONk3wFWJ9bBwNbxwvgaceFA/uA/rQDnCY
JjPhnQQDSmLQfiXCizYbCanjerTPQmGIl+cazx77RAECaVnZhG0v0lojoK9oixDK
ug0S4Ahiko/FXG6zQM6u9V4qkJOCBsJeRfyy5KwkSRknSISSaxS50g1qEkvDZdHg
6S30jfN+uJXwKIXFv5gT3XWdFQJr/GNJ/MsKf5TGjWoM0zdRqwJHIGyGYxFRZOqq
8eDVzUq/MGiq2giLfslUkZ5bDm2XuExU+14uBaYCgZ+OFyxuSrvxEmR0wK2fFPRA
9RIkdb7MGGZCCR9JgI37gLM0X9rZwRlvvcIa15GR2pFMk3U+IwYsbYb2FSte6TFB
/TYq05JPom1xwaeuXLN7Ru9Maewbu/tXoCXfcHx8N3/zMmqk/8qM3Hc4SxN1JT7I
jE4iHaRY1KEYEOKRehngYpRsljJ4yXDsbzgyOhITpXXZqZaGPO4eqIBV63KBGokM
0NLr3BNWM+bP8dPVFboaOG4YcRsnJxzNzfnGjUcnnpFoYy+Fy5H+/39L46zKF6IJ
qtkDpWNxM17BcLloppIGQ9kBQp8ynnqk+JVVd42rSE0/fY4Y27YEhb7h/BoIlOAU
PIKIZ1BnBni+kqqtFxZSpIB/jolWd/UGRMKe+C13jmqQMq4WFSoS0p0fzD24ITLV
8kz0Lwslxg76PMfBAfbiVzj4/DZHa8bjBBi7mnmQglZeNV0QpIPTB0Np6a+37OmM
Kz1lVMHU60SUim615vz9vlXyUPd6RJAPYaFTyh6VRpliSzIuSSSWztd6lVeO6D3a
SnXL5iYzSyuZe8KclgXhNfhc+u3O/fgtAAMqZNop3Y62H+J7aiESYFAB4fZo+d41
M/aScJzRgkts29oY1Lha2fZAfSmR9hf0tzejJSrjWi4IDuVFwrTwOgcJfFPHt/KN
K3jzIPS5Yuwfo+VXI20t9IPbBiH7NeZSMTAzAal/XmR130AYWGEiJCFAcfjGtchX
P8Yvexn98vokd61AUg3x8Q==
`pragma protect end_protected
