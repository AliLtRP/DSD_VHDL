// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:31:41 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
XcB9DqsoXAHipc0xjOgIEhMt7MAh3LMJ+Mm7k/qB5P6Tgf/8ntFZf10fKGOM5tSD
LinmaTvsfdb3fMhg885aePKDU1xo0mnw6sA4BvOwtBczgv0lrRjuJfwRyuEfvm/8
bywAcLCVLC6MK3r9cZHU8Zs+lWSeaM0HTtiPEkAjnl8=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 43376)
uX2iwc927zniKM4j/MWmnGSQeBIwSoR3SqDiDrsqF6EyvioVbNZUMaPf7j2g4lZH
iRvkg8S8XBJwAX/ur1y0WqvU7oXXfqF7kEgG02DbuM5DPqUul9nd28IcVV+cS1Ml
cBA+JvGCgN4mrEVe4DbvoZw3pIwex1mG6WHQGhtKW1JNVTP1BnqhbR+XM+jml3hm
2hvbFQhU9os3ix6kQ0iyfZrqE3Ef60gRVg9N5Fdbo2NyjUowvoMdtyEc1RyOyDO/
Z7YoHdN8josoSRWiqU0lCxCTfFTqVwsgT1zSghzaqYJkQ3iSsqmWd20d6Q57gih1
XiDGUC1f0BiKTLXC3aSBNvaPJ9/uhgoJN3WfXmLT6jPXiQfJOgj25zgAUHQpsQD7
3+u8BWBTJST5akKhnmdPL0OPIw/7Ai8XlV4x7OVT7eyuu8dVN++l5QI/nGYgE8ES
fFtWJEb7uJwKWYpmeEAecXw8NaF0HEAURp7we030FdeP6AcLskaKaXuYFPtDkdYi
MoOEn4FAA2YK9iQjEWJm/f/ComyLigvQjwaI0W/IK2g2GNYSHk8T8hQAqAtuVQuP
duY4UB+Hkn+vluP5Q39M1GWjqPYA9yUJRdL5vOaNY3wIzZMFWQ+psPn/hxeitFs4
kcC4nTfEwkC5jI+leFTqWle26eCJDWJltq+kxXcW+Tkoto9u4FJuQDzw//ZLEzOG
CVZ6wW7NI1rOQ1slGIzTa6j5ytX9wmkPl21eCqx4MSr7p5Aypct1epafA8ZWCY9W
cqIaDXCt3notDCKof6+lnOQHwo6sILkEHohMNcognchv8qMsvdKbUbeSfOhQ3eUM
kmZA7nuRUco0oOWUoHKAw7O16gvmx+j8Ob+BuwLMUcmyxkkDtZ+8cqyKa6I7H9bb
FQMChtXGW1tXjo0ulbO8h1ynHJwevM4z6/Ze2qojZSkSKBry0T4Qo7lP3iYfu7Zf
q+hZQAR31FfKwQ3S0NObkx7fGQgSpKCUE7XxcXc/f487kyMDxJBsFUpKv6Iv1tLZ
mLaecXG6kx9wercwYitLDCZqf+4QhBU4zm/INm+fJhF26urTck07atVYKY9JFoeF
ICqUFxaUTP09grIsd8qCC8QXASnriXIpAIJ/Lo7XtZApO0oDYKv54x6XOltMJ6RD
AEDtr0WL/dEjrBOjVyD3sDRRnlHUsukfyQ2i/5BckB6NgqwEnrKsyXIGEf4mks/8
MYCaxYjLprQpNpgAljHAUVANB8BEZEcQ5IJOonZJ71ZvsXqkHrV+puH4ETXfc7e7
1OGJJmMIOXIsQSIK6iuDgzzmhDGm4KvnRcrFd8QAlf2mCIRCYYbSRy2akmbR+LPo
PlVseOBexy4fGQd0GRZTwrTttvcaiN2ufaVYg7wfQrEvhbK0/5vSmZFmUB6AQtPz
TP7ZJ6XKmYAbk3u96EMcml1YV381txpNSjTvehwGQOhPhst6KgL4kNsHbLEnV4fe
dUvcOLSI6xPcY5iUXNuesBh0kHnlXvex2Z/o4c4V7rQ80TpQxJHgjvixbNZh0FrK
1+iwKY3Wl0kNuiKzDd5bv+vADlRlugsTb5tTPdV5n/4+RTK/Yyfcw4YNSNNuPzY0
7EHV2kFIZ4JOIC5vOx79wSot6XG4XZGGI2ZOTar92xmshh0wKj1mPj3bd7TO6Qlw
h3ZnCfinWZjPOnpyi61idQPc3svRo3b084A5sf8X4qWadLDOYzRH7m7hW/PcHyrX
UitX4I6I7e2szyWB31uHQWSK7KzBQlp6nO37vpYM0yqglzA0WwxralzyhJPJi+Vv
i7ARVnESIk/G1xuDiMCcZMM/ySxUxggLpFBCZVjCL9y+UxQlFaArblFNPdIUUkqp
RcLSSO7i4/CpPm0e9Yd58AGLEC8Qak0CO36sWCtLiMDLqNd/aAH6CrCjdOhf8Tgp
DFjSBw/zFfSGqwR1Yt+2M4oPvJe/h99ll4Xuow7yqVdUIH4vEO2+F8l03ok/fBNE
jTQYR3TDNUMPBHLDRz+S52102rd0uBJ1mCOr/tIzb9kLR4a2dUtNsAIaL/8WAcLN
aV1cwvcmLmLD10cZLLQZkgfk+IxbF7E6fmht4SNuJcsGZoKxBKjYWWcNnKi2kZy0
I6MXeGiQNKelhjGOAN3T2eamUAUKN4zBCVJ/w6/T4kRzXgPKg0ejUfJiCK2LdweL
0u5uTn/+dTXtSol6w9bUFdHzeh2MD47YbaxV4bOjD1tJRc8ST1eJo0res77KLN/l
SE+QCYGP7LFMsgYhERIH/Or2lEWNZdyEMt9e+70SrD1p6AA5O2FXTe3thGK6Rzqh
9PnDNLPp5578vL/qxSuvGTArVUQd/UdP/D/isoQ1mXuDyzdFd8hpjpryYbdODXYm
cad4XG1skcDNd+MIk+mqIyXy50jAndRT/QPlwSDDvmqalmc9QnkTSrOY1+XV1o4H
fLytpEucIMtJDQkUoeL5yVg/hEvJGaz1WX9moPNsUeDt3uGYyde8jqcm6xeogptS
jX9vUzTie5J06+ulH8MBd2no22JqSJfRsQXWTS4RyL9whEpzkLnrxi6KABkIpBZ1
ps8pgxZWvGT1zie3Ahb4WIvDPVBBt39JKpjHacXmfcAIOgQ/PB2JnbZqur2aRU80
HEbE6+WsUlS6grgTtG1K5HGvfJ7AI3v8t4/06ZILCO49DlA36J7rezXshjT1Od/B
2SGUvmg753x60NoY3Qh2DTMqQsMWAFVr15MdY6kJOcgyzuz3UfUT5wvCPGjs1cIr
jswZGZUdWe9kvEzIEt9UV4CWn8ZCWwQCoW2ewVfyj7cuqib7HeqMwkQP3bmuKE2U
EvIPo/43IYtHGjyDg/iqHxgJaAvebJHYwwxT4Uq+xipqHOuxalgXl3PuG8czGDhz
ZoXPYLDVV7FDFAFYntgdBOqcZCpPu1h9G88dUfrPm+2IS1r0iYV/1RJKrsE5C+3F
oE3iD/fVpJ7w873n+UhwgrWHgAi/KzFCjRNfTWzGWGPZ7uRfQLCqurAOWeVwhh2T
afSR7VhO4nZWWTKVtwFqaUCSoCvX6h1mGwuf0u9KPVREMMNVd4u3AxxzbFpeHjvU
x7XMtc/kCQ5/aBRXAkH8//Y+0yiFHYClqnu6GkYKIhRsyay53iZbdztq0M4T9yB3
N39BIOIplr0KZBXsGTl1CWadeWkN8A96YuD/VsfY4qePFuUe9hSIRWM1X0vl3ri4
hsriaSHKwfv2QyUQC81hyYfp7tc8WCTm7z2Kb+2r7pCqpDvAH1Ti0UgJOKz2Em98
loUP1jPPiWSgrOjDkC4gDphIDukZ+d9eKFQ1RDlvxE+KtQpIzdFtMvkKYHm2xxJX
qNrdjfCxkkSrzTQqegj25oZhwhDcouRQQc9eCw/PzOqWVraf52LVIRHoSwEmaU40
6l8pxdSHSoC6qYAH1YxwFGB33ZJwXuEKLzVAhfwzLsFEWWeyWmOjYkSvp5G3ZaCl
Se/mbW4LvX12nCIJN9KvrtzNhTkdmWXTDjjpsJ/+KOS7Lu04E9N6Q1nTooZOTCo+
89oY4fL/dBtnnNp2Sa/xJcSUj9jo5P6oY3bFBiJwY5WO2Dzzu/VTeX7/n0kNbnk1
UCUKORu5ZiglfLIdhczuuZ3EPwzgGqvU2z2vv9hzYP9ihm75DRVukr8KkAKSPNph
zwdqcakrO0k/lI/j9qnf4EFVCna+1WW/oE5YauzL6vfIK5riM5cJpDZPBfUtasxE
o5oVXIIyQV9v3vlyqSkC/zDeEmWJ6s1vIJdNNiMvtJ78oIOsEJMsmncokCaSC8ev
tR2BqStSvqDGcMH3IfHI7QpfMLsMypafkgk1PXdXTdE/VJxEEo1OQlFbR9rGOmli
G4GA7low/iMOUM3ml8ckPhkLw2LAHIkVeb4ER9VZY77zYlL+DAm/SBWNsDzaktVa
ZIESXlEDMxqujWdcXtZemixmt/GIjNf8trCjJyuq34hn6ilHgfaHYa0WQgHV1L/e
sqUzaGsoto83sMiEF6xullu3CBvzpMwpIE25bABCjGs+LFwlxL97sGySeS47A4s8
y8r3XDcRCesJm/QfN93TdBGrOWXdvwGXlsMbTbGT3OFx9D1xBHaU0XoolpiP/eQ1
7LwCvXBIHaQyrt1AQY7tcd8XMO6bfet8K0YrcAZ/Jdm0FV7tIRnoaHByZTLTg03p
6rD4FaCSjJ/EORpZ+uv760MNn3Gw+GDS0wElDo0kB2XvkJwzgPwdbeVSUGwerM68
ZbCj4R4uHNkBksfZbDVchi6GwcdLVmBSBm4c0/Yqg/nvXoFsrnWThNEYFWKcqo7m
jTEhtfmup5WJtENtkCswkk3OWLljx3DzTzuSOZ6SP9oa8yExvICCUc3+f4nMSTld
uWUlEcjcIMxM15YGpxvvQKbnBqlHzXxe/q9aYhz8J4L0ZUPK41G1OEVRlpQDaEqz
WFTKkJeo7jcyc/2QrUek92Ic1c5khvaNbaCOfXDJH/mp9lJm8H0Y22eiKk0auV3c
oxWWnUWAKTuNF3DBnDKdkWlzT9g49k44Kkb2b8lbzNjEvb0f/rg0HIxQsknQStDF
B2ydxkkB5n+NDIUamMoNyyZJkuM2OekLO7//KoVG6zPQWyT93ZssZBCc/QN1cMji
9Ivg84w69UZqv79RUfyIfNTWeumBwYubP30cLg92AmQyMfD40zPigaxuPws3J5iN
k5SpWnBmjr6LPdIJK0RprSc95dPcq1TaV2cz1x4EVc8SZuuQIq0icgRaEvtloEIn
Hk1tJetjzPcoLdyQpmYekKZsyMhUipcZyn+tW43E/Je8lEjXPdGZwlgSb8ce/ACd
vAtvLPfxVus1QW/IUOevnM3ZmUReWeE+w8Iuouwhw1aQ7gftIBTKHsr0AG5IpkmA
bgdQhV5qrh8zJ3ZR+S+D53GPyQVFQO0RervSFUjPCsoeyIeKHFD5HiY70go8YyQl
Ppa7VWawlkg1ivn1KJYZF2y316qUvA6T5G5TL34MNAUdCBQvubPKZ11Scv0g/62Q
y/L/GeRchvr/SXZQysuR43+BUuKC3YbEQwW5SmF2Eh4OgSzOwRTyadGOWCv65glg
vwItttvSRQ/sn3TF64Isz+blyByyni3Rictmg26N8Z7hFWcbura5frC8aw8nRwMP
VXGfgkgSKHPrU4ZoYDLixSYDunUiPihQTNkEubveU0MyeEsPKgYMIoJBCs+Mqs5W
vHLzbhMM1kAnPdM72xsVUJwVIJjs0QxAUs4KR4HV9+ao/56Tmgg9q3zfrqjTTFE/
kLjH9T8XizUzgbMMYWOLswznrESWM/D7Nyk3XHSnrOo//xqyKb/6vRrAACK0trbK
UExtNCvhgg//MBv3fYhaCUIBJtGmLjoG7UwcKjBuDVzoiLq6Vo+ZQ5AU/DJ5MjyO
+dHKIF7k9cG9CnpajnwSHYjt3pKfknpnBThFvlONgKfhSeHLtZFUlzMWvVoWRDpz
7iChRNtEzSkwLVprzPaWQmX2akZ9QsiCaNgXvma1V8cEzfKtDNJIZHQJEDgXvNH3
2CGyNq3n52IgXJooyugdodLjIr7gga0DA11g7SKOhUJWSXLvHWitjvAP6LHQb7wH
3NxoSSNlMiyXQiAfh6jmXynruaJlkfvz2WIH3U6trdfavLdJ6wPQwVQGqzO4xWst
Kj1we8523srgliuQiiZilgaP8rZexWOAQ7Sd/pWmtrPDBvRlwBgKL2jmppdROkzo
a6/rP6r6vnMQSzJTywzctLyLzurM985wYODvZTHbmwbmhQbwPujB6klS3pGHDMG2
evIhxKoOrxd4e6Hd+EafCNMyX9CGvE7J7f5UO/oejayvxfxHXOmHrn5i/YtiQGhz
VzFLxDPdUJCfc7M2pTVnAfT3rjLrrgar/+VZpN4uvU2HdbvX/Ebv3kEwUu+s94lI
5+xEPyvMAYOFi1O8g5tx2vOnO8XkIcwCakbgGFWN/q21TTT3dh4i190f4upkoOGv
40IeyOcKMkUL2So8MXUQp3ypEr9pXB0/VAiHmjPd0abbLPAEcT1kP4CazhEKz+7H
ct4p4JiRbt4dj87bv0NOo3JW4L6WhraeCnLxCWLpoBjxo9rQ/cMXUNVdbKeJZVeH
s/c0NJ3gG4xO/DckxhVJbRzcibbq5a9EB2SEBM83S8HpT3jj3Fvqb4VSsfLXYY99
ZGepo39oZEtHhjaJEXCdnAPn2GKd7aOH2lnFGOCBFaIeHISbn1Y3OAqDJltJamPi
heEL3lAGfTnKnW2531MsxTNTgiMWNB/WFt9xq6quSaChCzL9TxhOG5Gmg1pHn/t5
87DfFAhH9BVjeTL79gd0huLEk4VC2UxsXjpBGp8vS4JGNVbrRHL2xUFCi944tqMu
z7SiWUBhz0Qr7X0f1Bz92ibxm1A6mOqthpwEYaJZqU8veQ8WY8kQuRNYuHvcXikw
gYD0TCGORUAn3VUxHiNjIKRK/gOaP7xZzOi9r6YRSDjZBIl0F4vS+NRNmdZERH1d
Qr2gZMG+hNmCC4vjTY8TWMFyNNXD2EG0uMJSGT3QknrBL2v/68rUKIb2kD9LBoZ9
1pZuFJhdcFjnZz7GcrPfERxtohWOL9/6YKYPf7D13HBG07OjhtZyK0ZlBjEzpw8m
/Fwx4YzT9/0n5hWkgq4vt8bb+6eUaJBI0VdlKqW8UgAx6vyuRItdz2djGEkZOwOp
OpWPI1cor7ZegdNaErG2Ftd+/1PaJhOleinqwm+h8ZTUxkfbsSWxQc9iF04vJft4
60QXfNmpchJJazchbpzxmJTqAVgkokqp/K1ng6w1ev/UkgQ3GGuvAaBoZoZB7X61
qx/gce2pMzpA/tncqcoI9EjkmxwFgxP+KBF79VN1Tg04zhUN0a4gHc49WYjW37X9
De0PsL3b5eNAzv47Ldq62m0XUaiW9lFEMqVbdNyDcvJos3pol4jWPShkSN8oqkzL
22dgqAz1sBbagDuuel1pWTjnpXqohyuYDM+FDnvNu7ab6p8E2fz5tLax8knWN2Ss
YyEzTebZbYFOG3So95R+8Y4CTBG2k3dXiNCyVxZR3jl1uK2hhRr9WQ9gIxQI4+r8
AXTKQ9tfcVP2BFnM4l7Hxd0zHiwen9FQQsJUCtXxTMZD/w5fgX4DwYgPbiVKQvoY
PVtLdsyCZYn0Rrqy5IHSkCKWD/eUJS3sN0yaBxdVeWvYc+qrPVbhKcimer91HfAW
5+X0AKtL8Adk4zMQx+cpMD0fTZNP4e7sR5qk3smZhg+iQOfe5Xwa7qHt/SAZNrbR
ivHeYUMqF2Q6nlbe7UZGk/MkchQVQlCpFYyzJWoPfDcUlkXh+rHUN+9zCdUBEZJf
6sg4+58t4mD8Y34FlKKR3idtRKh6YTGGly3TwXYGuqb8hH2vo4h7DFkF3VPfvvlj
Km3b4Ndctnrx6wrifYyMYoi+drJAdQX7vxRq2QbHAN1zO+9c+wz4stgfzbnOQ32G
LWfQAZu61eyvjKt0y1F5T+/Ij8kodTq8Lj13jVFCPmCYi4R5LAj7DzNoXdXTCpbJ
zpdewHLsUbp8KnIdC9S0g9JO8Z0Q5jutBycIgrG1uMKHtgpmVS+u053U95o4S6Dw
esB9WhQlPaspLIaadojb6jvNu95TR3MQBRuIaM1fP1nTmFMZu/C1tDSNqwBflLaS
HyizrU2eLJC8cDQrXfpFam5BsvwFyVCRPmEtO6X++rb5OF2l2wYG34hHwuCIyu/T
WLjzFL74UOu3H5kZT3M5J4p1tYjA/1SKvCAC7pUB3eS0GZl9j9yblhZqAQNaB54y
VJvSXVcJo1IYTqpjDN2ihxEYhzhkaCFDAfADeYAL3ucQpxLi8eOdknFBx9yux1W3
PNDkJkBb2Ds4jJxZdKyN4mD/N1ndLTGFBqpuOda0HFkK1YTbV9rmFYxJCcv/za6Z
yv5DSnreWMS9BfR2WIk+92fp/gPw6S9hVno72nI2oyLmqCZKPHXfHWQUx2NZ91ny
MCZZworAtrdFujOgfcWPUHT5H1QEZmeGZES/Lwfcaxuyir8ciDg1qjW0IQGaBx0H
v5zDZOpW3ooAH+zKrmzVDlJMxL8jvjksbuqGShbcljvCCzWs9zn9A4z31YUTUTOG
XOAZ92JlHTuSwsvkl9UrzGD4A8znr9GjzO62UHSI5pQnseL/PB02Gs/EBoJhFk2F
140muWJWtbvAwNyp1h/L7gC6nL0z29ZlCE6qY5oOnnSgnqS3odsyTqoCmRx7hCEt
5rvBS+uFSa0W4prL479DsdIErGgBJdytLEdhY9aQYBB4e50YAPVpcO8ua31xyW8+
YTauidreZWEdBLpN33ownx7HFEh0i7/PICXMLP3a3pbxPBHMKHBcNnrxurBQluZc
xC3TgwekS6ooRNOEDUrORubEPXePlPpyc/CARPMMHC3dPj/VcWOA+139x1M/9h1w
tFaFInlQnpOuW4JrgsHkpupSkdVCcQQ+6zdZk+UK1pKWDaUoQ8dHh6ewMhzYaCSu
Bbpjq67jp6cXeTbGc22d+L5USsz3vHESbO4LBcDTYUYE5IqTiisQw5akCpzlr/BV
ChlK++Fpq6mPTWDrAOEF5b1DObOlNb+uIeBoXpp53HBs6eIXdUoV938pZKuLpYcx
z8MdD82WgpndKs5rSwzs8q9Zjd8pMMAX3UdMrKKrEOZhyx3g/cUGnLGjxLDo1HG+
o7IBx8sN6wrv/Q6U1V74oKVp7bZVLR/CREXz5YdR5bIN5QykCEHbOE1PlC5z82ie
STFq6JPFr71ZkDU8yGntvRkgJbxCEQ/hOUjrQmdjYClFuvv/Rw8DN7OlGHc803U7
SKGjeQuondVXNVPwzVy3Vy5Fl+iI+91MmN3PQd8/zDK5oLYCgwLJ2XJmRFUrKj7J
nmRQOfExn1WZC4nvFACXinzrnzRL6nXx0gv1E6cazpI3GblB5kAHz5EvowxDJm01
+rX7CpIEbTSv/tiwX2AG1lJ9EKBtRIT/czYawdet76Old8PsuUZY6sARkXPYbWB/
ex0lda2zeFSkg1rRa8A7W+BIhG9kQWJ6xRV2TgP4i6HYL4Qgg7aLC3PuFIUPlAkZ
juTFlObJ4knOJtv52UaDPArwCyxQZGMmj+8vNcD66f1yONOH+vMcXgkAm+zxavJh
KWcXYr1B433pdaubKWDvUx2Hs7g3EfdfZ31RoL/HZYmdD1mS9//R7GXndu6J+fsG
lEE2MoHUjoRvvLjoMjiOqfRlr119/3OJFUUgMo5yMTGw07gnxc43M/P8oJrY8x7w
nKmQ2GNARjNgEy0679WBfy+Ljf0IKauxBRwg/zUIyLcMXjU+ghzzpwYGEG2NLjD3
OQ8qYWUdTcAeEGWYwoLVWgr4N1dS9od2mmGSL+uhuZOUQCU6w7VFMc03HQlt8CXM
CvIN8aCmjR0AfZvfrPGgV31EtMwCRn4IApyFL14nk0enb24UxJQzYL4izBYPTXTm
BZYXYd8jja2WoTAmATd8l1wZMlpOjaH99MWbnPBKzF3cTKnBfVZ5WOq/GkrbxET+
bmmFxk09pZLxVoFv0hNUuABTUFqsK9IIcvyk/BQMQ10pe7VlZeSTOpIyR0+CDgtI
2QM1jAvhK/w9Ge68orclmS1/jyz9s6ORKxxM/Ki624iaPcUmrzW31n3JnNXn19AL
omKGGJhXCGXmzwAHT/upsu/tup0TCm60a5WTfxnMScEVfcwC19utfS+iMq4OTpsU
TltUSvInFRuhBIjsDH8KzmFeJQcHTSIjE16bcV+aWUlsCoBwIkhhsL2YbocPtMze
Vcv4JZrJixcKm9PSmSfRdVHL14TZVarMrw7wNK/rTeuk35ZqmMdeeE7tfPtMdF7t
u7EJV0mDKA0QC+9i2m/wlkY6VlGZsD9RcAb3JxvNe22SKhKgiBAnft/CkdQJluKt
VfU81ADLE2lUX6df843QUmr8S5ImaN5XVZHswZrdzj1a8qQto3eCkHPW85rxlqTy
RywpjmoNGmSn+4VQLGu+HcJf+nSx9eRhS4ywmMFm3hsrcHHPQHVGyPRh7xdP3kkU
tXPN5XnMUMLWP0XMDbkxSYv6H22YGTWXFD8N2ocxLnfnw6P4nI1eQt1Cc4P6nUe5
C0mIP5KQnlt6V/xMmN3xAotJJ7XOJHTQhfrwlA7EUM/BvsgW/g0JGff9fyOzosNk
L2hue4n4pOr4QDYnABG7OS5PTg8IjrQqRrGtecpmxPi07XZVnnSt66yEwivCvZha
Bqe9H3w3Lg5BhUblZBarwkdW+MKn3AIrjDHxHuFBOwmf1WvaAbrmmmgeGFz87yBM
D/ji4QMXdz0TTdFYxCK1DAdVP5YTqkY4ViuUciSQlrBzq+Nuamxi3BQOzHIqbFyH
p8j5Yl5ihBhe3aKuJD5ty2DAqJQmGErNXAi//bSMjhU7xG0S9ewDu+Qqam3wepFo
0t1PCv4LBnJmWTlwmAmfT6jI3K5q2At6NxR/1t5FysVKFruDCEtMeK4hnw0Vr+yC
AiBOQia+fE0h1Lo+kBYQBRh8/6X15Yqz2ot2tRfPVPv/W6GC9pBy5yl2u7vIqy3+
WE9cuGbiLmHBfpJt0vh7xNH4AsSGuUiLUVYL4/761yYGYakUacEyZI4KXW+uihkw
SExn+HSOfTVy0IvDK5oEScXN/Sacd2ZZUmSWleCflJxJNPpY45YUHTPnSE4XBHhN
7xMA5qQrpSHAtPVTWPMjz0e/RfrVvjIxx0r2qMVTMcdiUyShKIN+xcpjRVNWdEjj
LhXr2laPDR0B3GOjBhZctiI6r4qjjbaQ2dYSjEOWimcW0dKNKRKxBEy4mmV3niAR
8uSXR5tT8FoUdjwMa+IfmCRQjgN5yJsEPRAYuQr4ep8gyt3Vm0POpwUlVpnZFeC9
13iaY311dW20Cy12tTerRZan/VfNwZg5kxbnsTmD32Tmq8CYsZ9XN4xP4WsZTyfV
zuoB2dMlmtd9Tc+jYqRK4AMcJr9O0u1ZREQjDutXqZTccZGjijz7lp6cnRqF6Y21
Wtpk6xTbpPikUs75hXfUkc/E4iPbIw1PqRJCAhheLh9/CXDF/ba+ui0uUCNUFmiI
KMaRDDiJc2wfJbR/lXBv+EXu1Sx2/O8p0rLV8XVyirgGnt+tLmIWZBc1m7sr15o+
YuTtKnEAqFK4h3H/JZszDQneVJlmMla21zvxVXIt/inbike7sd2k4qBoy6/UJ0Pk
ijUqdvLDZbDhv2GZHpY3xu8dSF9yPKC3bNZ8WHWC7gw5zdIsbedw5fKWqnTXtRo2
uuLLzA4rsvZjUoFhqSs3kvj5vG8hL2GVUWphDabscwxB4EPgdc3+r06ZVyNhwBWM
H4nJA86Yz0jF6OimVbpQH0TSV1iSZCEsaCAfHJvv6CgDoVNDYmyTO3pFULMltwII
EU6sYdZBJBEbRh6Oa+RRGgmJQZIYUQm+lp6/XEu0KRKvDP/M3Lg/pspOwg1jwEx9
vxo3FPNKIM9SAhXo67GP2cY0WCLTikaTa9wd1MevnBCIwpcor1cQGWK6TVXVC3uW
yeBR0VnXc+QW7Wd2PTESIV7vZER9hvEQOmwOML6wQ7Iv5hp3A/M3vSzUjY/xZMQA
P5OSi4nBByXX7D/5CsocyKIh0dZDtiDM+zdmp1XJQIK+1WyV+odBFMVNmQhFVwE+
HHlYbp8jvK75m9/g4uQHXrpRWzwDJ7JlbEeAXbp2C/PHfFYa1blqQf4MdhCXMb5T
G3B4j9o/1/00Wd2gH/QC6qtuXCwuLSZ+xBbjL2XN1ulCpcyDNXG53jw6F1mp0a8u
jnG3JrUKhGwpRmG0NYzCOKiKt0S05Wp1UQlxKs6pHZ9vpuUrb+BBVw7qapvN1+RW
UA+wujVJmAvL2MropIQ+/igxhSrh7eqZ1fvjxpT9pkYgzbnYknl5uR/nZAz/keqp
C73+wqkidZCC6j9+63jDsU6jPDx8wAseN+PNp/Yn3b1Hk4aUwaJlsWzS0tO5KXNw
i3Y8XRwD3q/81BnPaEvCe2wOhKP4+PmkeUEqlmp9QcomOWY5udJtUJWpc20ar2G3
EMfLLMpZzZCw0IHyQS6YF9zyn4ALeTj36s029rzhpA1AWcSjkzC+pC4lk5Y2VcXv
KGIRuYTEP9V4WuxmMuR+Z1m52aDx/g+bKC672x9P90ihCy2ny/KqVdx+JMmJPol5
5vxL5NkqCrKDyIxNRHDDbyXUY6k4SC4AXxajme2qHX4sqXTz4Qse5rh0SwIq61Ui
HRCGy3K1ahMVNSxKcm3Y2+WVaq2ZEgtYQWtZ47aD3iDzQW5cHV7Y524fSeVAtmFR
tMv5kDIYZkdatsndqZ3+S65YFE71WeIT7d4yVMzvP61KsCy2d0gwp0PiNsCCziKx
RglH7K2QGJHk1UukTFX43WZhIIflLoZjyG5d88/FwaXoGWmpucKyMG+7URuzEzWo
r4HUnBBaCXJ5Ys/ak5fAOigAW5ZZVBltWRtbJRqXzKk5MIL9Ot7WhnW+E+JvsqOq
k+SyyMPbuM6Kk6PhtuWdm2QUjMmaeD2JykSXy6Br+H10avjkLp4OJ0dsDeNwZCKK
IrRTE9mmgaqr1Tp94IsrZbk23G43m3SWLWJ2Rh6aFg91CTnMu7W0fk9DJgTF0Bca
meEa9qTLCNycgThNp9ILYSuaEty9i34Gsosrir9SyI4SGTuiCX6cFkZbt+FTxS4X
DpEMoOaVoSQRxvaFc+NLktN3KSOxczx9Z34gqMu6m7gs1RG7nGwUyU6QfK2v9LYy
MQpgBKrNQi/dcutj+jgXVJrvagUYZQrogTHcu5uKFoZOX3sHiaV+dsFLIDoqKv6n
ilyzOh32uddAyU2kR2bSKQ16i+RYROCUA8Wq+12hV81PCdnr64ctLspCo6MPAz9g
TYFQXdDWCPnOvEF0JrgUKquterdhKKjZW0UuaK6ObnwrAjpBI88vzNgy1C5U+/ZK
/ZO97uu9aD0ybpjRCzxKf/DV64qZAV244yawtfKIvD0NLL14r1BvdzlcVG2o16eK
915+kuqf+G6x+Z252IzQ/aM0F3U998slGfkv0Lm6m4kvx3NL0m2tlKZ50uE33LFN
etHJss8FfPP0C0kKgA6rHQQpwW/ZIoG+b+pWbqQY9HfT+pAqnW25z+tECzouAClV
3FuugcvLRtsQWRXqoXM/gLto1RtMXByff8+jxDMtVTo5eCRy4CZuLMcAqB+DW3wD
rmrNMA7c5L/SybG2wMLXOh2DO0rHOD63xNoG7zedcEVkF4CWWEPG5awGzcL5oJ97
vyMSdoDlzkP10ogii426kevf5Igzjb8ZyQdP6/9p6dvbnhsr5Xw3h6Aht+y/D829
F35dlYTuHcu1+CVb+74FUdnNkFGE52X8+l8P/wNjGtvwnmQqkM5yi6tEmtZS17ZO
+bYTUolZPs3mcg0PaF4tXH2dsL7y0Gf1WHSjFHoVO+Qtd/bMNlbw7QEZfNKyd2EY
A60iWZDY8MP8Bg8acTtALRTzbFsyd4auRfpWAoum0MASnSrAScIvXWL0W5WBSFOA
A1cGdJ4rUr8c+JRGMW37zd/YU07qFIrgB8U4SmfKEuQpWI5q80IVPIY9E8Mp6I2o
21BrZ4ycUG/YWv3J8CMiapJ1RHuPkYMjSUC9jGZ7rOd4dt33ecX5q/U4joV9DLAu
y8VEGpEkI7yu5Zdy3P7w67kYnTCVxaa8etSOJH9YcR89kkp2MavP/tL39Ej44M2m
4n9cS/T4koWO1dF8GhZaBHJSTTNvb4UQo8XeUns6INbr48h06DH7c4UA/l18ORkM
a8F0zlbEZO1oV1Ag06iAO0vpjjmI717i/L9jg6rsZeDGZWs2lPCX+qrLDp9Uwp3R
wjDtQnyrJdvVTaDWVJUVSP8NmGz2t0R4lPKhdbP2+CEQWD+YZ2/jop4KlfakMJGM
BkPqFfYtvMOBqPXekiRUOiilY1gjSR5d1VQB74LB3YHuSgcL/WOgkRo8dCaGZpEt
kTtUeoggrzwr5EQJP7XYFUx94+zhH3kOi1+iZf+ZAurUcxAKedAI7BSVzcvmx4OP
xDS+thZxtRb/yCY8ZNgCY3J71SV/lkmkIxO77ApSdIiHG71fPUvFd3OJqPi3M+C9
kOBd0iMkSJYuINMsN4XUkm9jghzXaqY1Azw6OBTcdIVA1vu8Nq37DIhcdgQLcZVE
9eNjMHXtPHwP4PL7BQYrd+BMKXBNYxy0NF7GUhmC6R1ayr8tHOLHqfuPYbMGCaIf
TP/qRzBXEFX96k1SuSjIEzTLXrsqF0LtfOv3TSHC+yc4hfVjCYhcplbu2ePl1tu0
OHmNHygezL80nRk4n6eLSvKjLX9s4msGcWUL/iV9Td0FtXI7n3Z27UEi1QRg7aGB
dCNqxvFiVqy7zUcGic1WYDSjWjcQbyMHPVDiin0li73UmzLXqnpBgOKM2OzDBS0f
1ypYexIZuFnw66TpsZnJfTWO/82SmIXZz7IB6dBAmMdofS7nqhNudu/lug/aWocu
ncAcMpFojc3HwOblPUnsBMM7CROzTirNdlAKZGgpFBvrqYQ03Pdo4qNX2AksIRky
A9a6g1NKxwVYPKAnKaalPmql9dE1FF7t52G6wQHbgihh0kZgPW8pb+A/CjYOc8IU
TYFpNWEkb8nRvruaGEBJAIDO/e0mSp6mJGSmQXn4X43DH4F+xuWX0O+QVaw2TUg8
ubUVmMErnBXTT1MCF2h17ihEvyelVeRSCkavFx1xnMAVQ7/SiHm14DWIo7aaF6+9
mYUN0M3ReTfeXXD4twjsO+S1brOmV2E1sTFkYc05qK7ugAbFC3R1f3axKFBwAn3G
1Na/JhLbuMZsg52W46Pg0NddfFQyjYzqVpWIy8wfwpbfC6ZE8BsAD5Xhp7rg3X8f
/ckgimihxvfhPCDJjW9MFXeZS1nHy/7PJTa4I3qro5/YCE5tz+HW2XUTPPbYO9Ro
LPbAkTi//I136Fqcb0xrhnTklOJuOQcq18FrJllJcEpbla8NeSOBQ6+KLmZJUR03
oS2Xi9twYqAeQ/4g4tLq/Xz5L/iYy1wipq05ik1urD+qNtGKyXW2qPXk7WRHwaJr
/6Ri0rnA8LinAqkd7bZHlrGfhsRVHdwqJzjWeDdTxG56fQlFNytAT4FxASuULb6h
jFOYbLvxcWL7EwBmhgpr7xe7TQpkc+uGDcdskJHbcIeiBq20Ubgt3EQBqFocS5p0
ljzq2USDlRIOHiOXva6nJLP7ZRmmMkryr0m8v4Sqxt36l1SKhuHZ+aXjo8onj4zz
Jo8ko6VmF3uf8CfFTN7C8gnxVENhHH5KEB/EJrM2yqqAJL9YQnyuZl0WyG5OVTPC
QSRNY1K2DzYyvPlVpNFTjOZAFkir+eBojIJRZIIgyVNhOPGnJSAxNuVydNWvtrVg
9CCPIqk/gd7d4xhzzJsuOYsL484CZ6XGHFReJe3dh5oV0I9ff4d86BkG0xRNEe2w
D2I8ROVUqguWAPcfVoXrRysFZuFJN3XLNsqQqY/0zrSO+FB0G8GOun9DMe1XXt2+
k7W+jPja+ypcbfwO9B2tZTtoo1ipe9S6X4M+n2B2FyTp12fRN8Kl/7XjSg8hyQKR
oR/yRjIJ17rVhKNlCy8a00tD0PIt++r7RP5G2fswkwnaLDnHFQH5Aigi938eSx5b
Q0cAwqRRNb8Pm243bP1C7eHdXxM12bMmss2/Big/0xLMKMoxlng/xZyJlBwa7mcx
2qFTp6fBUZiYQfsf6AmOhqFY0aN3G2yGNTFe4lXVH0C4drybttj+iv0bJ1Vrg82g
WHW9d65y5G9vqzCLo80A3lMG/zg+Zd4RBAz4zR7griCcSNKq04B71D/P4ErBXoPb
bqI3W6XWXhZpEW9zBf6O4TWMrJNbluQ3fpVBxYgeYm509WEvjImTIgcx4Pk9G8eJ
IH24nBCwmq3kRFEcW53yB0Aso2SQsYumlRibIfxsoOT/dOk69InTncDaBztG0kMe
Ps6q7XvNPTEjyhfkA8/WWn+lT3I0YxVtS8Ecq8Q9yFkVJnogtKuiQTtDXZolZPxw
XWrSFVXcK7+fJuApL2JNwDs8Bn1RQ/9NUW48VR1p4MVCBQjIdlNLjam0xupjnTIA
/Lqa4nwYNhgiXzLSugXaCOWlRoBvilNV9v//El2tgo825ifw88Y1OiOWNZ6/MCB6
wtlx0f/ehUBD8IYf46Wmt8cE6rt4cfYSR5qFpjEIDBex1tjhliQH0d+a4JNOJTsy
P8EwDlZ7lMZiPGdgthjRpdmT7It5P3BaDgq2tzBrsP3B9OHpK7I2rbT7Y/biJH25
arnMvqSJDrwUdSLla78kH0ZfjlMZ9UJimX41NGzv+u7uh2caxOAS8cymS/QuMnb5
kNmYi6l/NmbWpIXC7cmkvSzdshBSccK0IgLP8WXNU7K8fTgxWMw7jZgyprvm6krg
OBvTmQf49tEOuPoYJ0+Dln0zTzYm98NdwyDiUZmiR1Sw0XfsHIm2YUdZzXuZnt2V
Yh/Lt33iU79wK6OyMQekfu/VcRLLhOqJi0XVjUbMcJ7erffGzAyZqnhH024ZhMCv
Cu1eULQE58n/Hoboc9DwuX0Fskieq4M+CWVIaHtnAUOivrIzLNJIeNKkFn87OXkW
spen2ISls4xzbVQT0mfTR6B5cvFbjhCPGODirrM+6TCOeX0Vr+nyr5nR+Ob5gtkg
sG4g5zSP7oSMh0Iug6BC5eJQ3bj6LSdO6aMzKSerrM89NUDL9xT2DiJCrkEtke3n
uUyq3xMJ0oQckfk/6tFxsF4EP9VonU3Rc+Ig03GSuGPqcGUZigOlPbgmckPvwtsW
YoZ0eGdWfQys5IH1//nUBOxzB60TwQx+WNWxT9xmCkQfWeKxDJ8BezMifGIflbMZ
ti0SCYlkoum05iJgLAIhrSVmNxP7hAw8egNyU0JdobjwxdJlaZESnK7wV7zGNSl8
KWIGz9hQxrA66e48ot9Ascq3QqS8w0g2J00SlW2U5Emr2VZuxghCQQ+JrWvy1xcc
NoVL9UbqnwRx59w7GzodsnUEb6myK3FuNHwFQgeOsPP6ekjEXsbXYaykLSncAkPY
R7J0iXBPWDDJGm5EVALNjTi8dqEYl2x/gBevsuEAUEh5sRWEBK+D5AZ6APXg+ABw
lQATHHMRYobvFOPNo/4hcszu0bubtmgqzlQUETcCy8WMkSo7cSzq53TS2+YUQYHd
5jr2ExDPeyBaMlOQWv62jRHwnIwoyHjCzZ4BSRaX12mJdf/QL9pCDDfX8jUPu1Oo
JLA5O81+4OEk644zgbDRVyzFqsD356+3Z12SVu3hFNBjJZKtUOOxCSw4s6nM5Qr+
PIOfYhgDI/os01qBuWprtA7r1QUXUXk0KJBMWnYrqHsh4jN5t/uMEg2DFh2zNwD/
TsaEFBH9X9YqbxyBKyl/UDZgqpigIq9vyKAj1BYvn18HQMSZlpA0KlIHwaWGMZLP
m6h8vcNGuA3fAZ95qup1TOhWNEfjSWKnOIsvAsqLlz0ZZzTk71YZsLAlJIsAemZB
cMkA0iA8/lmNCS3WJ/hTKoPTqJGWjDwkX8O+02Fq7AtI2138EhTNKA41VYPQPvLf
/8nxMJpFqlawXkPpfKHUfkpOO5cxppvCnYbUxxeP5A0XLGJADsFdG7ceS3keNoAm
YT1X+XNsWV+sSatahld/B5JqrU3G655eCT3EOPBKIw7yRg9t/4CoHydBtz3ah84g
s3rzL2nXkcoK53oUCzJmwdLmk2UcOaEo1C0pO38nWEUI53o1oCRmaLXvkamF9BS7
RMp4YG7vEdeRlZwy3IWXAUpIPoAMdUKBbShr8olDQ13bk8OFStfK+irWffYuncuu
zHVGsB6utiDLg2b8fPzJ9Ta6kO87wOxUa2NhGSosaFRzsAzQueiJKH05L2cGphPT
uiJydc3un36pecCcmE1XZZCUmMRStbTxqQNuXVBKddTw1X6iUM6KVtfMcip/Z3fT
aLr15EknH3vL5HfM9QtxaxHNFSpZ0ppv1HKaDPcveGGfEkvSamsiIJtDQJTZ/IGa
8MPXnSyNlHePRbCldgt7rJXyt/nOocXPX42ZJlKS1B0S0w4auvaNN+3pzqBqKyLI
teLLc+U3RAOp+rk363HIZg7YreyU4VAbVIzwHAroMP0IQRuumCC+qKbyWY0FpnMo
+yuBWcANHTcBN+iVjG6N5vK0dl8hWQYuosINQ3+kLQeOllBQjLEjzpWBl6Ru0Avz
Kg9WkxRKSNImbRKkdXIb2EzmJs0628IE88pQuEI6elSfhYEcS3CvuQ5LlF2H76ja
KCuQJSOj8kVInZSXhAj0Ub2BHA0h0+a/8ND3ythLh0BSenH6dAraSANsksUZxPNq
RCQARC/CNJm8aFIu0r2LeXA/mOAjmpU6CmIAdu7dWLC19BsheT/2UxmzaKGf1uSL
xzl2JEn1OkRGgdDn0XvXEVU0DY4KaP9DcwWd1/BgvpsLl7b5x0dUB9K8KFPaQ0v+
OIabXI4IYW2wmo/04FS+6QxafOdBE0yvJPewAXQLewhZOw7e3Hr9wBi6Tbcoortr
GsiECKnuhP6sHEzXYSqJ3T3M+4a+huLbScS9Ogll3fX4rWsboHbuaIYROAlrLTD/
5fqzl9Q1zpCfdcWLDtYw/CxRGCi0OX3HLpQfg3YZaWSCUigGkag4vDo43MupuS4q
0xeZ6wCAQq6y0YvMJSit2orvWt+FnFcIDOZ0OHRLRJvcB2mS7t68/NPSPbQ/ecLd
I82yubfQY3FCz1SARNfyUDNmCjO6tT79NuEJr0lF8Cm/M2m23CbSjs/o1O2r9+Ju
8mz+NxwWWsE+Daz4aB2st7bmEy+daH13DUZaMWUZsdqBo3zNCNRgLy/1fVIhm+XU
Gaerz2+riDZka6onCZhM040gBpmDkWnqYWLO5kkSEay69UEpzLWFGi5KFyKXEyng
xdwJYhnH8pcvdKMYUc/6xYNl6o6+wBwHIvmMU/Ja4PH71xA3mrdDnHWyumnd2fvx
+/PmPexh9yYSFjX1rEUh5Wxgx34z/FS6x3BGHYuk+GGr0B6p9RPjO/3YnjGsRFUM
Hk+iHdOM/OqvPwU7gqt7hWwwuyKA9Vo+KFSUEondJjYJ4HbJUnTuKt/mSmbG1oC2
Wgv75leYj3pmFueGKQI90jHJTeoApg6XOqXHq5wUiikx0eVS7BcOb7Ksx9zH5MOW
PUpz43JwwNbfEULlfaYUMrYkRKO9WyOpQa7a0WqkaxDzWyq0By2ZXTu3vNY9Ae3F
S38h71tGUZhTrdL2Muk993t4zxnoZmHaRZX4RtfUvGXapXPbNJ3uZDcb8ZoqgDVr
KOrQCdW4Da7iqB1dKdJTvcij9I9agNVxlqjvaH3uM43pTc68wdyMlAnbO6PPN6iY
oXx55+dj+DPWOJqY3Nvrx5biXrzzoTD0NdJNxCyts0StZsLIx7DGVJE/4/a0MSBz
Co7ikwmxFqWGSjypWRGFUkluNXHMkYlOh9ixY+40tSzEMmGa7Ak1R1zQNidwb89N
ttNZnPIM4ll3XdF+qCAH7hxK925Hr2loIzb8abNevPxBrrBDBxkkZzyJnZ/Odl4J
/UBXptfmvwiGFWbCxtocG38HjHhLzQZg3T/oopzRvb2qx8A6vuYrvS5f0hFfclT9
COWjF7gLhoXTmTkYVvKfqHSd7tKvox2MEnPU/EqzKTi9yjvDRQJ1Negl+RZyzFLL
k9MNa3sYtWtUB1WNVDnV5XH3q14QN+Tsvzfok2OH5FXkwHfsbAgP+dF4ptuCPtkf
+jpaldSfxeyrxBR6pWp70fI0ekSYIV5TNZVhqJeX5NasOcGhEpZEaXOKH0Tkv9Xx
OZ9FFZ/CZCqjmI5UzzkWSwWARN5ifc4yMFhZ/usQ3OBbTVxU31F7ymxnlw+FkDt9
+qxQRcyG6v00stC9+OGFiEe38fw6FL2nRLVRTwVeRHcTV7WDaPBkRUdXOR1Vy4YI
0ptQjQlNuC32307bZ2cNq/o+QtTZGtXARRnXkCk7s8rcDG6JdAFWJ1OnhpwG0//5
uo8UslbUgAkUjnBE6VZHI0b/lW+bBE+bIa1PgViXdFdgDfOOQyU7yhxYVB1ylza7
T4UG437muArofT9wXa6JMJ+9QIwQrwMK6oYyfuILmhtPaqm2Df5lPZL5V5d2fkFX
mwcD/bSqvMqw9EvDtOkgb6GtCbzp2695abiUyBdWwRbFq7pH/16c1a/s5clQ4WAP
6cDISYQ6cm6PS53d/o+TC5S+rvKvrsepVIR5/8HJEO4SRJn2W12GDfz+yT+XM7uX
hqqTF/jFzvYKhTp+btRbUDhi2pnjvP1lcM/QbjEiB3hAp1BPzMPT3pqnWfcox+dD
fQ6p0z0bikLQLPZRaYcbtQhGliB9wgjZAXemUdM4reTenRRQmWqhbcX/quku2rqn
0QJFzo1lCNoSvwt74Uj9rYvyHTF1LkunsWd8gNTbqwGZFUf/33FZNASpx4Y2MEmi
pZ7SEVmC8FrLw7909l4RrDbRc5hqTa4OwwyV+HLYj1RL/czXGXMLr8YBWDah2rVB
Y81XojpY3AxoM6xnjM2rHK3FwrrIo36qOAzY6gt/FnIw8XZ6B2RmeRa5BUYMi4gJ
w/6sXlfNBlRmW6Y0M7ixFV4YndBHlxd/ycFmBHMqSDEhMn/diIrk8n+6mF1ZvVIw
uU2gtYg0fjwxS84JeTVh/mo7RNJqHj9jLdmoTQiyeIO0oRvuYWFq2kQte8R2tQnS
BNfvQcPZv3UTUjbTaTuGyDfNEJBHjVpY0UkAiD8PqcY0VEh1ZOAb2xohmMDfKS7u
Xr+VWjxFWkDqIcJ5OMR6NPXh6xkga7UyhVRgUlKTuQH8N4CgxO1bSCqQ93iGwXFc
5CrAXgy6rku4o4a6uQGlmq/4x7ENbOD4LvwR5Vhf/npWTf6x2ars6QxXrGOy5bUB
LpG+hYakNSyTppXzf3NrcOUtNobxFxW9TVtImNbc0/4BwRv+kfjuwKWYpWq0jY3U
vitnlQwIJhr5n/jm4eApR6xorUu5SVWOVbeXpN6RGhfLKR2z32OtJvJPQmRPvoIb
WtaZ6Jl2pDMQF4+UIR8S2U0yv3acr4zYiwo6hBMxZWRbTO6H9HLw8u09q7LAVYuq
j0tuos0CWPKahCUlAlny6M/KQL6dd8mKama2naC+o4p0R8TXzQjhPot72kVyNw/6
DPizsVQMZS+im+P8dYpp1Zu+RpLZw3ALzSlx+fTxj3QTPrHGzdYL5qWMKu3+Z4jw
cBAajMGTA0cTek/SZk4os2i4I8rTfnHNlRhPx2/bmsxH+LJ9wPL0cmqYEUeKTL5R
ytQxB2LcGuXLCzTfQDZ617HP3Si+cSGoJU1PaZrt79zy9bb6UZ4euah8tWxCyI53
sKjDdtFdBOYBEyA0Xmx0xo6gdqnLFDSWjFdQlHnaAydvDDnt/fKfz0hkc/mUPOa7
D71RjYCbCvfkF1YSNe/RzgbuF0q3KnvtkgDycR22MMa/3IVU7ohWqTKh3TKhx5FL
oNqqx3a0b2AAggNO7VJ3wY+9TaBWEocB6rAB4Ixrq4QVz7f7s2UX8jDFZBT2LS2O
VE/UwuqJ1elbetlAGxprGapenfbEMKzYFei/wKNbMduPI0Jg7B67+khi+ZiUjjSt
dTPXHeN+kFseFGQdtNj73Kltcpm7NvqbCkaQQtL4YPcGWDS1gUdLqdfnPjifrtUx
jMZtFjq8iKGxW9apqZdyrcofmYOb1UbqIn3oLUfbfinqs80gqmbwvz/g4NQMIhp9
ThnbUbaTlD01s8PBef2T76+accdcBcyJinrbAD2zPA4wEcZwSxpjihmKv6bf/fl/
BEv/2k5aU3HCiaLQTf6hsAnvD+KnqQVIO175LRHbK+cGEXBbK1Ksy2YGL4CYGCNZ
VPYbN2btcKp+h/gf47yfTia+YAByelZ3FClmCYr2tOH5wfzM1twbcJogXelymABy
BJHXEmdz7TaM2EIkpf4MFvuvAynTqMcUXNNF0QY9RmNZJRMqGucBC5cJHCLKQFLB
Jr07/p8UdyMKD5VbdtYU8BI1fV2Nw3pV3+8NU3/BOY8MZnxsgIAwIpl06EerTKP+
Z7S8paKZ/Ffp0NJn13dfUwv3qDtZYnysLrMM//braQhIs5AsbyXrtzms5DnWqGj2
jqjk4T+NB/Bjup1J582afgkSXLvI6NKJahhhywxVzxm/9Vmaei1I3GLqiO5GQPvs
rc2ptLoCijiVZwhBZly5UnDcSPYOQdbtT4MLdWUEsVZRdr4fQ/FsrcdY/GRcMgeu
hh1DmKF31ipU3mtX7MpmAw4uxItb+J31oC/ftAEx2Qd/JwaNiVUwtin8SniyGRtE
eOtdYciMaiqT9XPAuOnd5CyJjwScePsAV/SbBmW9CHwmMcAHLwhdLRcCEJ2scrcF
uSjZpTqJYFYqmjCsnwSpFxzvWMKxamXnEHr41Udil3wIqmvY2FEE8dLQnGlvTQO8
c8v3lp7/11dQcYsUf5yzt/ISZzFfEAWbkJNZq12qVdII5EtvWlkKBtDi8xYm3ume
UwgGtPke+3ZXlEVS1/LKQP1dCraW8mTP95G5AGbTe2oE605yGM8RilExLCb1z+Fx
UFbNEhRr7XvRv9iE9IGtpAkmKtpFRCbQk5Q+we/GKFXf2Yz1IDPOJajoMZ+w0WAS
phf/pUKokqFPk0C3mGjakG93JI1MAwBN9w8Sn1D9jvpCrj6dNfOpjKuHedK6ZLjY
xadRRJLuIoXXzHYstGEX7ILZzHAmO2sh1xlsUdTCk0H+M/Ud770k9GFUmFk2cpUW
MiLpkAhGf2Z/8tZxdaXnrYpc0Zha8SQWmAYa+BFCN86MZTpMoTwrS+te/jXOQ+pN
sFbvy2WYEETNyjcZGUAj81KPBooDHN0qeD/b6wBdMtDPfX9k9EQ7/b3taRHxDU5r
9zXaysmDbIg8rX89ZOT5tZC8dTIqnq1zkyoXthBirzh6l3tmrLuwpj+ZbWc3qlVM
UWosuOk6IZ3m28nr/E2fjIdrOZmdvgOGkKCIz1aCYIQbqGPoNCGd8rWd1QgJSOhk
LT2560oqRNvzbVzs8PVZrSHNg/QVP+Q6A32CaTP6bdMNNTVv/ilnZkfu/5QwdyAN
dsz+qP8yWMOcz32HyTGUjpJwhVGuMjb7AIDAohrfcDK/Co2SgbeF1PFh0td2tESM
Mf3FKAo96uMgziEan2m4W4lKIGdj+k/4djoxuCYIEm0EWVH4/HEyPRwKD/ufQiOT
7jcupWIkF6r0Og97lZq5wQVUEsWv+qAmAyRISGcm9KgsgKHmC4c4uzncsasDIr1c
GEk/d+NZ9dSHSl4KCQq4NUXNx1eq85Z7NG0iWRDhAfzJhdN3LyZXnn/l22mj23os
8OYPOtoX58s6fpbiKgObE7FvVPSnhUFzsKlTTLGYtHs62tz6IOG0hlca5M7RYFq3
o5PV4gMt+kaWA0GoCUIf+JyyahL/a04s8okydyHLErQxGnAPEz9KhrnP08JjC9uh
c7ALVZMaQI1SDFFq0GHdp4JSdQMR1uINE9NsEWctOGbily7Edp09Ecaqxym6zO06
muCUuj+HGvyAcGGemWlZ+ZL9x9NA7tvwY7BllV6zeXESwny1Mneh7ptaOlMJZ8uZ
DnJejhiys7tNUsT2xmDQlfknoCwpXaVYLAykgi/zk92kD6aTorJjbWlhifU6L/xZ
2xp7efuikdMtTw5I99YNHwatW7vn8Jd8wAL1v7q9s96p8hxBd4AG+bnAIvaNwYWK
W1rTTQb7Y/uTGId+B6/vtVIObpdTuPXcb8o3rg4Kkp7jPdkE07VjWN+zzYZtppms
lo3Qh2bqnq0Z9I+QLtt8yHDoOolOgaZi+OvkL2BgxsVVAC7T1gDnaMk00OpfSBjJ
GmI6fB9gLl+Lh3uNsLB/0bXag/y6GTxCC8X8tSonUB4goVmZDOjHoOcQLXjdtLrj
a8+J35VOAzEKBvVr8JmPx02ZTyWhZ3luesZCwIspAwj6DkcJAx7jDej9ssWJ6dXW
imlM0ERO8g5vey52McArInKEZHxvmovSGXpH8M+FhKz/njcQcbYblZmpMVx2iebz
DHp67fBr+053QC7o9iici9Z+7zCaRLgu33hH+SUJ7tmfuKCrs3XA6QSssTwIOe5n
/OkTXa47KezQ5hs/B8KS9IqjP5Z1MP2JCfD+qaux7Z/Kd7q2gBagituAxSvHvtsu
x1qbYc1B0NsYzzMf1liqpjLkmUzYEcYwEfyC8A6lc6cfKT8KZCQhUeC5wZszBuzP
oUJXSvXWMfd5FugrSEWBGT/P5PquahW6ou0iBREGQaCwhmcTjJQ+UK9oRTOWLGpO
6fdjS6iLNoK9ZSfrMOWB/5neGvX79GO1fZ2JZK+U5VTFSEEAqXa5V/dQOJSFGOmP
jAS9w7ZUTmCPLcjJ5NViEWWuY+LTtOtwKoms4x/QiXBS6uTxq6ARk5fSmYoSIK4V
L87afn0lYfrAzRIZOjh7SJGE1eGo4PkE7RgT3bUuv367z7qCkpT8Jd2s3V6MJ9tA
xL+HeWzilGd4Iud53/TaY06qf8BrFuYegxWMfVT0T0s0RilJHAMjbqca3bNLJVWT
Vt6THYpDL3qxVPmfDqwM+wU7AWehDXYnODTUVBOqGm6QLq83BMYc8yApHC3ffzP1
xIlbZKprFa1sJ198mMC/7XXCoXMMLNjRoq5VMISQigHxfl+ZqrH8Lem7gb7SVR8B
TU+nwsC0bnT6wBcFV5xPxHGLFpofffqyCbepsDsB4SLipi2acPyGKDY9/0MaDv2W
3kDGdwpFgxLw39O3fo7hbLMp4VE93F55Xg8R4nLbYNMBEx1wAv44uwkl099Kdfrg
EeAFvLvHWIaLuaoa/aTseULdTQT+0zYGyj3MEPTRiiwteJJRgvP2socnawFhd+3X
juu/2Dp2GRRgKmAzS8zfdBh3qEaRl7wg6vNXVCWxi2vmEank+RfRXoqLclTYHDQY
Gz1Ea/pZ9yXaRnsXmpss5TaS1sY9WB0QTEumM53KiWgptgYkvQ7BcyjmtjPI1PXf
VP11E4SQlA5vkVfGyyNbMD+3mANE++XIJnQrfgVBGeVfLen6sTE+JGC4ZPa2T5PX
Zu9MLcmsBnOCAZXmGzo9oTQWbEEvOLgDir7DzIRknmoUXua/PE9JQP088Ly8Q+Tx
xehE3mo88kOiCdJWfznlWaYSiin2lf/vqECY5ZxRwdEnf2kUpyQKYz4dQuW+biLx
zjVlem/0w4Jpo+zGFoo3PwTvl5wjLDymyQ8qJMyjefZJcILQDTzS7Gc6IlrV04hO
G1b1644YnOoXP8qNr2ta7tPv073x3/asxZz2JguQxAK5GAzCjvTK0Z1cNDBD2Ba/
lySwTnDCRuq+CuRHCDF5mxDcRNU0YMkn54fqhzTsuVsw0GKb6CcY1plUOa0w/ubT
B1lBvvrBmGctzgWtjK0Ym4jFAjJqOBmnqTODOpk44GdaiKEv55VHmUrGURbene7M
SI07/4rstM8e/pyfhojTY8dKznPKdMYBavCqxT6SlMKc5IH98wJ3hclDL8qxWoch
kd8TWVwvORViiyUX3PxdkJ8Mi6GbK1DUV+ZvFvctyABLftlU4ASJN4R38SN/vpt0
fvXaF5rjNFAxscKISVSHwRp+AFXZP70QIq9xIpfB3+fVyhK3Ww0jH2GbP1SvpqII
jQEm5ImIxrDWEePVcKXmo2KYvOdXeT1fuAw6r4JoHJHPEQ4y++TdbiBKmtfsYVMs
IRJcWv5CQq6t5FT8I+M/xwFtPzSN3txn1VjzZlRlzSDu7bnOZl4r/eKLGRrHTH8X
Dt7bNmLKe7pq6rfTP69zPp+0wY7RGjnRnkcTmwHfCzSRzLzX4yBCdm92FnUDJAl1
VBIhrzJN7BqKhbz9qZvh1MlAuTp86JDEZaiVlQGVwyBESoifS5QWPHlQsfr+LhzK
op6Noc6vY2BbQQZD88q8rORHlhEAa4mGvZX/MG4lsJOwOrEpyZX0h2966C5XIcq3
ttvfgPeztoytW6272zlWALVvr2YnEPo3OgWUBa/xTHroUGoLqQL/Zqti00Liu+LM
pwbIc05642QOqCTrlToG2BpjuG66xuKXOPCG4JzPSjhvFbbwqC+DqCrF1mzano4w
WF54Kw9aBqbJVLAEL+Mqfqfq+k/RP4wZzLSO1CR4tOaHopORsmNFnA09bYol7Azg
N691+uZCjQsdNpw9j+2doxzSnf1yWjtraVCJGCjtiNS0xCNgoHC0QHckMZAyYTb0
L1LVKFZbhM79kmtKjBtEfsCaqfxTprSI8BEMoID73E1fyZgsk/ecdzfdCfMlkkOk
UaWa8bvsYm/LYVJHlCAOe1KYpyTRW7EcSYjvP7YAxiXBqDvxa3TKK6O2MAJVuits
PeMbVJePF4s68yjHmw2RZIT3L9rRS1OC8zo3d53L+u4fjiq74CU89npVJ5hvqzBR
maXBK9iGPAzMRBB9ycIz/FuYYKNXfdjIK/yO6lBXcRqJqfVOd/Xtzy8RfSW3yQ/3
/NJwP/KmdqgQ+nDIXuN1afAvSllWItHpfhEarbnwACmjU9Rw3rl/Ld0f6YKvLMGa
LcShj9BQDwaMBB4a7HMMBZjwPh6p6rUcCz5nOqNYPU9aD0ZuD/6U1MLF46EavSdN
Y7W2GM9dPF7IPHcuVK0GFrT3jKFKn6BimzUfl66ky+IQQpgFBZOUEmT6ccQ+5nCW
4n+Wm43gBz04UgUY9nEcwfW4MRoJrV2a9A2RMUK3SIadzlHixrBlZaXRJpNQSAne
rqFFAs/OWyVM/UV47dcDvdS9UPfY3KcgWSgE5n9RaE4hAxIIFGN1IufTNqTdQfEi
/N4Ny4zf/Qul61gleTs1u8801tewOt3IX4Rm+j/narf9heBDA/nYoLd7KtwAhtk6
mo3vSi1lfKtDfn8mJW50MzxFg0ytKZXjYo3/xDBKpn+kw8SjUrY12FKNrAB0SsbK
LdK7m1MxKwmQyaIG5c+x7WS0cMUoXnrrW8xU1arI2921GoKBlI4/+lAZhVdNKGIp
dKxKisBslOu+eJ13+OID/L90sMiu6Mb15GnPXcZFA+n5TmTuABFRMPNbXcvoHFbs
D21jlBw9W3GHg+Qb913ZqNHaLQLSgmSZxuNtRdQ4HfYSnBjTewaMgBOJk9Db9HfH
U3HXEK67ZzJ/pohsZvTkZCDf4r58HSYikEuoBWTWwjJoLNFFTGFmNNqh6/F+mrSE
nOJa2KLKCF8Ql7Mxr5nGIY75leaItDqLk/U1oVJ7F27UtN2yotzm7P9RZMh3hc0S
+mRdB45Lr2Ew/79cu7QIX0u8PEOS5At5/X04tEdZqzdTBE/W+AD4IOFMothHoG/V
XiOemuBQ3MaLzcoS46B40t/dXT7kmLlPugvphXyKANPWhxbTJyXQB0AXM/0Ln+nb
+cwOZJ7vatuE43PaFMAl67qPVvx7vwItTA2K4hfnUPa+cEHXgAaczPYBnjLF42/n
bkOlu6Nc/0mep3RiPULnnATxToPV/7JTBHwivhKN+4XqEpFs1G11BFbqf1iMy9uQ
aAeH/CipIm9b3utqqGQ4h4LkM+QKB8mJmROgArn7l25XfJkaSC++qCmKU0FWvfZ7
MfxMKtRPL5SKvZOjNIRrn6ath9Z5YbMjpv7mYcFgoKMv0N6t+Q4okUJbRK19Z8At
pp4wLvNU0aepndVx29O/sBQo8Pgu2EOGFenXNXj+5IsoOnQ7IkzB6c/yF3IC3ymr
fDHfvicjptOVT1vZKpYAVqL5udlYp8U4doR1ghbaqYzTKalL9wSjybMkx5cGTr1l
Gc8E4OjUWTyQcbobybIhyE/SPBoXWZxmXAEUNHjfZU7qSf8ZPAENFJ+SJ5b1AdOf
Ac3L98hbkR9rxSgZTnpJWUzJ+gbs91AA6FU6tEpWfPwHrm0sfmi382B1fM8CPOHL
TDDJgd4PKlcFDAHxssG45y1JkWnik2IMypHpKRBOgfn8/3U2ShteNOdYSZ3NE30t
9ghXEcu02pW1Z/xsApvGGPgILwBfcUVkALngQJL7ZfGgY/1zIEbAhBjdwyb++m66
KNTbHkwj48vQsGaVNyCSr2klmYfR/fergugB3JAYINk2v1zNunh3Ncn1OkCFzpyz
ci/+D9l3EyamjO8y+foYhazQfVHZLzGDxyr1/RuPSlFr8JT6eQ13S8U21u8ZtYy8
DKmidpFjAFEC/cYU1UgJykAHlvV7TNBTdIilCZ1lwZ6xvCdxnsRhfTKDBNmWPryu
8ei4amBJP560UgyLffYSaayzvuToX4V/5a/2+2yWw70c6l47H486es8le18RX1uz
Nnu9oP4Db3S1wuQNE9Xwa0Lr5mRtMATYhlpxH5O3fsIKUu9RNfhexbvp5x0cbLLe
7SO5D8czwG4dnmWkuQ5e49uKPpNeXSzmUd/RBs63fb4hVyZJebJ4niZWxKve95+H
v9Ea1ZD0D4+5N+q3UBDxUyZDVuF7qJkZ5bFYcfHtY88ktP9rwfqvHxuavGgGGnjm
mXEjja0txIep+5BYZa0TpDnAcTrdpXb20ThTxB+ELlEMTSi93Tg+avXbjGJdQS+D
vXdE9tMwrjUoKmn13hsEO0Ud8B9UnLTKgBrUkMClLqH2ZJvx6xw0secW4T8wWxmP
njH3TGEjUh/Ton1R43PY1rBOHlhXbCF4jpv9gpyscn0OWbXFrg4xX8FOi3UORhHT
cPbNNJhoE2IwZuPSNNVUlfU+gKK8sKXl5JkeHU2rzM9/UsLUyfUhu8zz2qNAI3XS
3A05Fb7/LOM8T/rbBb0kjQ/lKnfVk4RmS9O/FZf0P/Nnb1AqSAtRzDqBLwSfA2C7
dbXYapRDk0ihW2Rjg+gOPhBxtdA/x4z9w00U0Z+4+xmprObhPw4a14eEzPIoutQk
FqbGoiBhFN1n9mMOrfNI/UXwSm17GTunUyPMo6eUZsDbQvzfhgXKY6tY9ohc5Wv+
vHrdAHPxBDm/WmDWFg/99lbswi+hCQ4tggKcqGQq69hP1Ppusn0SXe5q2dzPDDYS
OAWNv4m5a7eDh3PQeMJGcf7Luke1pnCZBU2gop6qdim5Ob/IUaCfgQkqDhnzPsUV
HsYzuU77wontLuiU6NomycmWfyQdKmgRS652XQzscK/oQg52TEothZvsPwdHh7Xr
WHZIBlS9uwzXDNxoq5f/3SK9/1iZ99c4ZCAZGsPyIZlO/RbNMklv3nKjr6sdAedg
ouT9mOvhJ0+BiGGkuglJ4utYKtOd/8AWMzykJA2XTk451PJYXWpq1iVEeafkL1mX
N0c0ZBDJsBqnLIisv5L8veMULdXoabmFfmPo2gpYQ0q7RQ5AOZZQrLW+0zHzXWvg
v1AOG/922je8fP4XDDtATcoZqZGttwyKkrVDDVLQv9J7VhHpX9ZKT2ZgcM/LsWlk
d8WvDfuvX/tgTwJGqmxDsJZswpp5S+X7mBGoy1+28eEFHPAop5vZ9aq5olLXbxJ0
L8ItjM21lzj2ZR99m7s9xTjosmooA+32AayI4BMvwiqrmyQEtmnVaf5QZmchhXyJ
ecd+WY9X2+seZOi7DR2LNL5ZDF0GzdvmcnlQwzga/fUA1lvZ1WhDEk3GL0jpasas
uRb8G5CJjq2/LMww/dt8ulId6RbHC3l/vrC2jhuNuywEQldByCHC+45CJK5OSo5Z
81X5ZA4qjFWbEjyB3SBuirY1HDthj8IBanMuQX6OP2KM4Pjlgk0QYJ/IRAbowBW6
NG3W7n+p7zghOUuGxm1X4CdJiACLDF96yVcVKgsJuOxtAD+wUS8cbUxmKcaRIJHl
oM8ixo4TxOB6m8cLAYZK0I0dNAh+cxNx5ymP7HEw1e5GCEF3l40OTo6ZFiHzGFae
wYuAcwKsQkxOoJLkF3w9bukj/+MBLIOsfZah5JHSUMbKmve09KtEVVxdG6yzn51d
jJ05wV316XkGDKiX4ZoJwtbja802swwm6ZogLcV25WHWBWiEkSKhgnGVK9Ew4f5g
bDb/dEf5FTmGU8oR9bhujmAxQOMh5HWtkqQgE7H6soFpgqtULNyXHA+zfl47q9K3
RsK8qOXHgHaYAu8asBYkOrEHZNXjQFpXEzMJlWMMLkOwPcSwFlEoeIJf0iZ6uvcR
mlDkh7mOeI1YD3EvxNgy4/m+5OlVGMYemCabxIehhJ2kUZ4O4hMc+9VFc67bfaNj
iwmScccwXsS4+jjDl4sp53xP5Cgnn6uBdQtU+XhTFInU6mCumfLY9uEJcmCMb3s2
yL2niThDShr9jRfJHWoJKz1x0n+eXwRmdazbqh98VEk5LxN04VbOJtpnf7x5a0LK
6/edO0TcOclwMQ1Frrgky9UGKHvMzDrHmkANJCZ5QCDgpriqRvLAEez4XeFPs9Oo
HGojXaiURG4gjfTO0bONO2fPFfsyUQ1R3HZ3IlUv7DI+fFOcoNrE6Kv29iiDcVra
nEftHJ1KcYBYafxdMe9OYgJy6Ds0gCE7sE/7Mx3eKYKwDrd9/ApFB0LHPPjInyoI
YhlIAAHOVnnlOu7OZXPIFAOMnpvTotLExvF8pwjTt0T0Itj8Dy91qUF7M08gGsSh
TG9g/KbaarkEywoRsV2IMkdvHqZ+HcH+ft//q6oJLkYMuHK2npgPvyFLQWQSJ+5r
4lIyGFWCgOoVU9EhdUh0ohG20MiihSVf2x9nGKpK5VtqsrWlW6xffYOne+KY6HxN
VE7NUehUV/LouUHxHOFcUslvbqm8uMR0NLnVOfzd/dFZ0GVg8Wdjdg205s0XECJ6
gkIw+Y7dkxwdZ2a218dHp8i1mBJG6y4JD+3YICB9PeJlx3tYJ7wfHdVHUrEDAZ6U
D1ek7Z8wdiIPfB083J8eCTwxNPti8+XF0AlcrIdKo18JY/niQU3nqljsW8J6QuKe
V+SDprxSYAGNF6eercn029FXVOCRK/NoUJa9OeczQew+uiN9jqbAPIiXd+FARvGY
h4kwHSjg2ihDiacdUt6avRL6t6YR/efMArP3x9/Ud1n8BbI/3X9trUGcXyTQOgfx
5N38AIVwzYlYWhYaDBn4hybWVyw7MdumgtwUIudl2TpR2vclFbmFWqIQeKV2/kza
JT/9peSYfWEQsbEhgsx5yuMvUFhQzFLax+XlOCDiEIdpp0SOBYTAT3Afp/pKSfRE
GEkoX9OJubRKG5GAJv/r2JOlk1tWb9eHBJywIaxnFFicl0uGyJax9YZ0ChmJTxeQ
nd1Ar5LMsyFjUtF5/QVA8E8DbdW7s/F1UJGRUclrXY/k0cz2CDazWFwYxwtEvcsj
tBEzAAv+Wd6mwi4nzD4lYnTLZo2D88KAVwXit3Fqwj2D6UKbdErf2gJTNYxJ8N0c
fvx5GEUaO20nm1g7DxEFvoboWzcZhZ8JgOhKVmtwBbR/u//Yfgy+AIdvqZXChBUR
0vDTcflDq1AbKAHpUSRcJN+4la5/xvQQu5MRNwfHjHDolF6eSpLrCQzvUVHGWqVp
ZjQg75eIpOORYJZ3vpfXstZ5cpUPO4HSExtNprqy3Xe3nSfWSxvesqmDPPkXqwgA
O9mU58YVYEjK3KRWWKHWsfU1YNnMSJ3mDc9u6mUXvTHaKCQcAseuybUoTQbpEP53
EujrWCnY/fdv4dUY0LjKZ29i8VRtUKNSb24wUK6cMaMxiz3xlqxM+PYftEEZTpqr
36+WM5HQVl7EQxk3cDYnSSRSXgGDIjFP6MNC/NYB+f53sgeHWj9a66PqhJDvEAGF
hP8FMr3BvSs/srCJW2Wgmihz5gAolSxo8C5V2ZBg/E4YhOK9I96Gm6iWGMtiVnhQ
meLr0DXIoWk+50v5P7UwNgPSvxOyV95rVl9b4nMmYsYvH3teAak4vRG1je8jD0Nn
WSL9uiq6/zm+1QRwKxFvXPw/OroGYr+SgDjCEtC3y+vLYieDwnnQFBf31CgdipO+
JWn3uFNpBsiY3WedtIRIL9y2vOnAse1An5pUAVt6n/l/DyHsUd0dfYkGqKcFdRgf
n5+drz5rgxztGsiu7md58z8yjiJ4yoIriSNwYpCYMqM+3UYETf8NJ9ccHoYJ9kda
H2tUwNFB3ekH8QELDsRf5WvHgJqFTRQjaHTs9i2iQLcH+DCXfMH4xEXVaep/jAXF
6TQoIViTG7jCIAAfWoYbcte3eVidTAVE53xbckI6+LMv1fFbXX2R+nWcG+yPB1Zf
o7ENWEQBK7Nr+W8s9uboaZdYdddBx/Y69MMd1yojEpdZbdviZO04vbuxq6g4sk8N
2FvzowI1G2u27bcia13dlLceryzgrrnULezrSX3p1DqhVYQiJudC+I+cDOJoSwug
L2McjTco+iwmKFnWJ/OBq+JswoKAGF45ys7bsmAX+15+/pci+UwBsAYwBPMxtOPt
4Hv2FChqxG1/SjhCS9SvnjribCwEj/FULcCqPf8KweHpeaIH3wqhrO274sm1DMfe
BXj/mFFAfKgwqtEMan1vuXHAn3kTCAOvCH08J3eA2/XpRDrfWDvMucZB25tFyWYA
G7PZa/E7CUSe9gWGjmP/GPWtMZvqR4GdsGc3RpCci/fjvkvrWhmkIlHFM3t/i9Af
M/9iGDZjy1Y7PNSfwfnqS1UCyo29vmdx3v86HECkGJKelQogfDIKTvjANDSKKs2n
tobhAxExmCNPtU8uZxbozt25heapg5xXYX8q3qAfwMXfOgMFo1lDFfSjtQy/yaG4
XYG+0qo8huFunkSkPIPbyGBLSEoVEexSyki1WosFiQ9lliNx9tDA3dYCo4GXcYlb
zpTP/9NHkLOg1R+H3w7gbnDdK/wrGZ7SmMoumcMtTW29XUfmERDsiReCWPhg+Vqr
WnQFYJaUrkUwgfSBLpUWR7cEKfU5Fq9Sda1Ql/70cHsAt6vqaMYpxTKaRt+vm/Tc
a98YZSniJVQ2LXUveOPgA8XlkJaZwcrOnq60ey4X+4Rp81m/M5DLLRrAXpQ/khbI
NxMrznGj1FF1Xh0C4bYYhZyz/w5Ha0yQuB2scOdbEyCtZM9jjhj5X6iqKG3vR443
fhIEV63/jvNlBcN1fnUz+QZt83b/JxfD8c3JbmxI85jImjjaGv1rCnexBcQDlqeB
EaEKs9+BQ1FTIY+3etbVcDqoZ2qIWfWoNTAAttwF+DP+WB/uIkn1g05SBnAzuPUp
Iq164c3jb29R/9GwOf9b8Ni/DN7FIAqfIdmCO9gAEqnw5m5pN15p4GLr2ZhhdApC
E4B6DmoW3zcBS34HsUgi3vTr9PAaT+WHvRV1vTN0a4BK68RiGmuDR7aTRVRVJ1h/
SM7S1+Uk8+Cnhar8Wyarz25i0HhgoN+7+jX9BUdMOTVYFfH1+rZSEIj/tBuYVlOv
hBVIPEPnSSxyTyxzR/5JCFLSqlGJoWHO5066Kdd9NXkTOsH1Q9TSik3dxAZet7wP
7MnYYoPTQvhKnHEMgKAHsAx0n3RJ/cjeBlUiJRtGiJunh4fUW02AQ2656ko75Tz0
JsX4hrqS5WGPmS3pPK0iZLVCul4gVRVqnri77G2f3BEGvbDgTinF+72PcCa0w/vP
l67qUy4bjQ5NKx4jaQjp5vQTqnk4V4XDRyNza5sRzKiwovc56o2vHc0qZg7UAecY
1tCGaQY4ZKXRHTDYG4nG7Q4T9En3H/O6FuKFKL49DFBVEhzfVVxqX+c5OWnVVXTI
XpIwxTUi1B4v5ymorDyGhe2VlCKfY53JgJQVNRPHuoIeH8j4un8R5l/TvfCtcTQN
+nW0HCBamp2xEvxhdID6WGDr7iFQCB+t3Jfw64M8rjr7fFXlATub+DIKir1FGyRm
2W/DAmjnFg1pue2Ze911mw4/3y60+oXGrYWpTCLD3HubdooeECNpMQS4/tRrFMrz
L8OHoooUpHu7ps4fE0B7brLF5WVUVI6JsZz7pY9rY5Ji8f3D0xdue+qS79nBSnx3
p/ncVOvKB9Oqo3ZS1zuEsa8l/pVXsl1VHQgcG7Zm3DGlY4eBVn+0XqqtsKUh+8wV
LsDud4nLBz9SXL97GoskfIW8h82AwXbbhlmYKUbiBzfg3X35gXzI2XLx/dc05FSH
IJa8+a0RCEBUxe43fzVn2PNlrg/HEE5dit89KNHYxdTJJsUuW0/QD1IXLEZy1a/v
QbIxkAkl0MhcqkPHG7mX3fbO8CWIcyTfFXRGgb+rVshyB5SfG8MVP5zeVhyNmMVk
ZeSIrAfRafLiDq8OxMK1eONnEtY73J3VPL+yvRU/0QLaDwJIsT7l0b9wEmnPpMw7
Pnhgt0oxp29CK6RF7pAd8OZdetWH7cPU0kNQPWmOqf7w/LpzonWePEqk8L2FxZKw
/UW2ElgtvoS+zGG3jvMYcfD9QuX9Gz5sUXFaMC8nUB0aXK9RXlr0ylMfOYUbSIen
Cpke+0I+56qrbEVksNeN7jeIv7nVBe9tiRxqqhohGs87NTdTTF7m1mH6hghxkjwQ
g4p+mtDM/7goR9/A4Rn8jmkpX1iIjlCHjcVbiWdiZyI22MscFcrSo0b7i7Ppj5Vl
Xdimw8gBXY9Vh8/5AYu3rbHyd62hZxpWODU21fqtG7GuInZfJEy/HkVor0D/6Gsn
r6D8YivmjrMO5ndM7C1KhoB9KD33VE2NCGQk7MWAAPndwLIRBDFB8vqJXv1LO6xP
BJmPGMpxw8AS0zE06QlmuUrsPfoXbSAQNU00gTh8SwAqmWN6tC5VJ1K2ESfadPQe
owNzRDgARRM1ZZ13/2W/R+MLWcth5P+eK7lwu9SDn7pUibFf5o4yYmqseUYBVCjM
Q+KKy3hiVerJYHS/cg8hdyiJBpLM63LdYHn7e2t6G1vkzXigplx19C391niJaoIH
UvfEdvzIMPye/liLl6WPtXpJU5HARSOcST2KjF/X1mi2Jz2bgrYyR21cZfXQQsc/
xZde/11rHZhpS3VOzpdjWTiOitT/eTGA7pwzA/VHWkv+bB5Lyimw/WEo8mPNSwWt
Udk+jz+QfcMncFc+Nc88AAEvivv0ZBW1QczebEsKwD2iscQljrexAxlqF/T4cCuJ
f52fmUZEChM80q7UYArQzYonkVQ7lH+HpwtFtxdYWa2CGQA8Ap2gL7ukOJ+v1pFB
fw4cELdlkgWnnyajfqvFRwWhwU3PiCiqZFwkIJKYOCn/EN0eMp+b0SBeXhbMsHSL
gbg4FldNOUvWaK/9uGV9331H1Vwjz5x2j6izeRR98Gsyjwz7OR3G8baxuDHuQL66
5XdnT/TN0dZcLmxKDySZQInK4vbmGKSxGwhQ0/KIuk1Jrscr1imoT3Wqzk0sEfUt
TpvsKBUrZl2TKi4rYlempajwLvltclE29b/PKSuKgjsZWUdmEWpPEdKPzbW0I7xC
I2CTEWaXERex6fr6Pn4evYrVDrllxkpOCO+B1tm2nhqd8RBGta+GbH0mJbVifzSy
2T/4KmmhjDt2z8z24lB5eKjDPvurDwBvMbaetxC2KqyIleA0czXewTrqCzcH2Frl
/pnD7otTBBcG9hx8/EYtUdVyrG4mCmJHyw3iMCUSg7v9ly+appYNXA7mnlPRUtAJ
kwg89WZsNTtYeqznAuuA/5lAwfHU9/1Tg9FQ8rR0W8x/1zWBXIYg2BqwC4FT0m1m
GXP4doWbusr6pyDtQCu3ER4LljIyKX+tRxl5fzaLQLpa4pmr3ISMnU7O5V3ki4I3
5dyxPIwTWC4s/hpsQ6U73p66X9syZYn8m86ikwDOMXyIFkegdsOAPOo1aI2owpjm
11bkYTCxO8ms0n9oWZKQMGPpC3YyVxLy1Sh5bSPMB1S9vKIgYb0svJA5sb6IHhMN
NIw0agy++VB9rJk301/ofKS1r4j3sHWOL68dSSjH0wTE4zAl3lCT3b+K4Rcvx/Ch
aesbaE6Wb5tFJsqiyljFYvE5Sf7XWYzI+WmcKJEryNCes9Wax6A/5d/4Zb+RXx9U
tF7y+qraYluOECDvyOHOMCqoANFooY8xXw1a6NjoLy+hisVN9vWWPjednkZ/UYxd
SqdZdGqJyGmStcarRVVom7tEvsffX6CCL9kEgg2eTqUt2UUtC6k7qv9x695uLHm6
pLAbEcuf2GUHVeHgDtA+pGOqEZ8LNxUJ1F+AssDqTPKEfNJyZ8GCWMG5PU6yOO3v
rREn++7ohEKEVYFV5iTFV6kiZLx9j1m7l0ZG0N+rfusH3Osl7RvBWW5heYS9M6La
kM222ezQw9BYpL9b25AQLXAL8p+h4i2LDvXVrZ2ybBbQ+8qe4CazAM4aTYawdRlR
S9UQvTfFbfDea9DMChfZO7fVtvdEuAwOvb/pUxiF3jNs1qmve7dVnwuABqeBbGR2
NvjrEfF9DTXhSgCdjPc3sTMPiXV/yBzMI+RULYrD5LQTcT1lQh4qPkXuQXrMCS5V
n51M5xeGW2Kt0betPCb+QcR3ykrhF9zcmPGKPjmdE/ZP/MuFYyYXbK+XkQYQNzmO
Qpd+zcGHl7Pl3mcf8DOiVVwq7QqJiGwtJC3pw2XSJSdyWSbj6mZz8i3WPEzfA6U0
NVtjL1ZNL2MaeaH2a/3B+CQaSFKJvTHlm7SZKEUPm/lDn8KwMdcZsmzKNQLHq0lE
BHvDnKc6wTmvSspY3QH9RVyV8Jv0EOb8DEfLLjB4O6P6pI34jZPix4Y9L3hHtpZb
1p2k4wdsUFmb+tcr6clb9CrDAPPb3qgdcxFd+oyGsr3xXXUpr11viYdI757TsaHQ
RFDzvGGj1LxO4JxSGdd3jbRa3pvnyiWDWjhLKNPv5f5cqNXgAWKTT3h1FUS11flt
sM6Lxw6wOenyDS+kFNNbQCH4nCqGwV1qOMEMVrmyVPkbwVwHAIk2BEoNxY2eWOiF
faeC8zx4fCJR3JCeN24Lkn0xpvHG5MWkc4IsZYJail4tT0eBlF3GlWCV7a9f4o3r
zkfqfoRYzk0QiGEX2Z1G3FEmB659kQFK+LUipkwYmbhROvLj3CeSGi/7PB8oApzn
giZv6B30hXubLwPyiHXaKi7N9VDmDhThfUPyVXsgcXwOH1feBC5MDyhZ/2vecNcK
LyDHNUmCaURM+Jigc5kndQeorL4VtoBwKlhufEusAB5Zm+KPC2pxVXVL0/LABD12
YGxQR2Y42QsuW2GoH2Sh0EK8FDAXmyXDXxdxDa12Ux4HxkUk3ccAgG8C0wSwvKrr
xhh/W8L5XMDV6BDHM/1AOYEKvUJlcPC+/tc4rYT435GKuZE9OQ8SHRD3fa+Py8eo
YS9J4IpNfipYmZ8xzZR/OMi+LQhA8Tc6zSJIot72HZFPUKdy8Qcx7Hu2JNKockqD
i4p+fj4yYLuvZ/WIMPvZUU+MVaqV/CEKBjerq9CStYlsW2iln7Vns3l3KC/HaUJ1
YZyv7GhifRHA2nYqO6ySSuwy6wLglG+XWqRMWPyQBIfBrNM/GrY+TTfhdFJG5L+A
MbUR4tytmMHrQxTi3iaeGqqHU7MBt4i67vIgPstufLyUkvMaZU5k7BEDb3ehq8JB
wbE0zowYuBMuVRHp90By/d7K5PBc3VNky4uqO3jZDG8tyNoN1l/FjKZ7PA6SPO/Q
X3080m3XmYWbns6/D0Gj7Eswytr73zhPUNjCjmgkkmEeR8yehdf9zZA0bU84N5Mn
+2eOXsMykPvBEGsXwm+r9cZwJez/dArb0xujqo/ghj/9EXkTBWNVHX0UYZFqY1wh
avEEy6idXAYFfmhPDuv03zGM6bCBxDit2lURb/ZOCSvVdpQsgImATrqKHb/DdGiW
gh0+8i+Cogf92GfwR5sOxB/Rr8AB/tmf6QthsyKG6rzk7rZNOy5P/KPPvgY3fM8C
m7ztdV5AjUQu7nNNqYbiWIqeX4ORPIrh36gFLS2t4AozVjJCzpIuM169LRbeUaR4
htO3aq3b0uU88TMpidTwQjfli46OzUb+Eb4jNeoNGginoCaGlY6MxhPeJb80acLG
FT1GES/6pERRuizChqbtc+ICybkxryED3ClH5KWPMKdajjja8pBjOHiajFl/ap1y
WNGl9/FwGMFo2TaCBOjG0eEngC2yLTHoQCW8fFCxeEtuUFy4rTDJStjzGoDhExm7
QRcNc0RoPHrTnhe4/aisinSqaQjD7zGHGvaKBbs0P74vWXxX9ERprHVmBar4mD49
66PiOnymKEY9ji1LEq0dEUjixorN6Z5qGYvxf2klmYAQNOeRNS+OF59LeiT/pJ9o
r65um/tsQjnU5jV8ctcXfVsXSda0qTte9KZuvmyvyDUU7BIQKzpfT67DT3Jf/oey
iiJXA4DBSC4rHGyElTB6HFwakM2sSYe1BquNRWnkhqpnIa0nkRBI7CtziWuY1gXX
lWqWYi8FtMrzrxW2BMmA8igpsFH6wK6oDWQrvamb2lNkPvsY87Ie/qkwtnqQDALh
sRi/vncaw5uY2dpCo6WLHS9AWvjdgYNBMrNdyzBnI4bELRNBuhNc9d2CiCFbUKAi
Pdam7aSRlSzvuwcYSGn2TkNp9YSj6L/P+wBak2b9yuul1WqxYy0T/FmciB9tzypU
2fMORQeA335zf/VK0JKqd0v9ueUFOntUDev0zaF+POMll6zuKYmsrMRkYY65JXxi
1Ck96OEj3ie4KPa+pRJ0H+MTZxfyOz+ip+fRIWmyhf2vkOqlX44CnUh2+AVqlOc0
FIwoPM2NLPpDKpnwX/yBBj+iXHh4eiVzBXqk6t57PA6HaISCo93PpvtDUtEQMSaa
86kl+tZBxCpoWrVoZkh/MYVK30HCzLgqiEN8sKFwlg0Lk4XqQVqWGfF1f3VvW8Qd
9sVPPT59Fa5Xt4fB/DDezbcxKII86KQlrU4Znp2x6b2qL0KZcKJgz7m9ZQwZwxBq
xa4IsONhsnCMRBozMMOZTRJl6rnTyHqJucg7mjYtcvSYfyfxjz7fDfzLZgGfJr89
Kw7McenvUDoLKqv0hMHZnY2yelIqI3PkgeHB0IeYaUqVJHryrZHltaXHU9aes0Vy
MUF0xWHKIUu7Xr4ciBS/ZCPplFj3GfSn9akYZD/bTWn6eWMdMATeVzrjI62y6Cxw
kLHy/s7IQLY+j7jmK4bsDng+XFCTWs56xHPci486Ty/2cMBvJPk5aC42VEbu/Kol
7flTfz6LP2PoPfQ3uwt63zgzsua+D6vyeiW9cF1pO+cJftqUpJMNRYk6gXjaliEr
9auKU92G4GgCHQhTRffnH8gFBr3cmZbIPIXkIpG5QNEtsiCYluhjP42I/RelNW0+
Wxp7rCpKU1Gr87Y4tAom8FGF1fun25Xjyc/V/Qx5R5UMMibx80pYLKhcfeSkW+sK
40lUM1HGfHdFI/z14ibgBpBafktqI8X97gakTMWf2VUUOMJtmi27kGdr5/vase0r
z44rwZr/7uoqhDxjYBVmBT9tFXVJGuGlt2elsXLEeE3+BIfNzIFrreL1Wom8yyPU
2z3qJK5gvOnSgoMcALOVexmHPreu5E/8/mvk2NHmpKdEWYN+1T+DqeMuFF65TESG
Bt3evI3laUzHqoW7Gc9S9sgGrxNfsVAToLKDBaIv8XA+4ydMYluGURxGh9y9vNGB
pTA4Tfp6/p+gO9LFYAu42KzZ5f3LDrJ7QNvwJ84nkIcAmdTZtVDyFN4Sz+SmoCnn
C16JgyGXjdW4s8zEqDZJKNhA62nJWkDh+qbsvbanYPoARUzHdcgvWnsotlb5+Xi1
9Yymn6k+LF+wXXSJ80yyOalzgJu/YKg1VOcyDNytQLHyiB42X8OYQKzXO4bEDIfY
kD2b+ND8TLtxACI3KEQC6a8t9MkgQDHBUNpOSQyZHZN1wOT+qbgGNu1uL5tJ0QYT
WHpHsNuMFLnalMELptuEMK2LQUQTk2y16To7WNqjKEHlEEDDiL/rXYhynoJZ+1Np
8pklW7o5MWdsPLdbR5M1YbaoDUnEX5D/cC4/XCPvhfbA7tAqcbC1yChcgMW4zrF3
LgjIHuUOcPOLLtfs+XeIXdZcWtWDv5RXPJsZWaLfBSVvM/X2yc1o38T2sNjBpYXX
sht+v2XoG4u1cPbwfj0fNtUJuCGHka9l5wf9vW4rIKoGBwxr3TH7xq997b/dMQ2N
Uu9AvoqjcJpGZTfZOdUd7oCwTr/I06JZFjRzyB4xEJps7kNsourciuE7c9B09UXT
OEiRkwzG8FTjPyyYAaYsLnceDIzwmeMJnDv8Mhwf1KzlCvlh1YriElpcSIaitTba
9WSSK2mK4awNiG+gaX22BQx311b7ar/PIfORdYdUKcxqvYTqZHQPi5sANBtbxTm8
0eiUyMkiNEBXgSlvwwzipCAVszexDu6zXjBWS1LaDivxaoGnW60YSYUAiaDf7wQA
L+PA/XSzYuCvrE/LV5OAvdvLfiY6u3o8fnSMlGSbY1RPD0LNs87kuo3NeFONhq8c
B1O3pc0S5PiuuvcNFcGFRVjZ1vbcX4fizPpVl17sp1s3TtpWPZuTZ2ROFOTDCeK0
9/oTbpxHx7MmvWl08afJ71hARp5sb6f9jhq3DBi9eW6+ZseK1oF4YnEs3YXMJXjL
+jBuWUK0tJz39MjrJRaw1lCFHSkWBB3Yh2U87HOes8oIN+wgPgrKZj5CxbgvM+eL
flIXQt464E2b9JWJa38ztC2YG/fa0V+2buzpuxSozyUgs5jGeThSvXvSiQuYZKlW
2O73bm8yYBQF6fiZiaAaqUumyL3PvdrCS/oV+zDCTNigJnLxfOB+ymIjfsK/b4uc
53KbV5mH36R8SEg6gDTdgZXp8oYddIZY5u3ronGTIXKFRAsnEd1xqWq+3yeYYpef
0fmAtpMkH0hBNsvX3LkgvfNEK2d71lvPMMfbVfF+FR+GnlOQMsXxr6H/K34yGPz2
q5zIz+vHPitBX8Vvyj4ymrIs9vbgw/IkatfYHRmoZ870cSAD3HhyM6MePXMmsD+u
HigUv4eK4vKJX83X0+AMxRzNoN6w2cvfgfGdOGdl+xAVuwor5QI/KJhbid4qYLei
cvdXUYWmLa2Vhxt3h2sHjn9droz9y9aUE1CJZDfN/pmWriNbqD0U+87rlyfL5tI7
Nmn9exNBNPJbXROX/fD1WdiO+ZliE8ufa8Csi46WHZBp0OF2+CjHfZBGOw44xhWm
DtUgwKCTfCvRGlKtWXd/FKZ4qmfVk9ues2+YMgJ30S5Igw1GySnvPsa/rUvEyg9P
IKMP7nyKzbg6ctAInF7vIxYNVxbEW9ncV63R19UWSPF5bDGZy2NfGUHqA/PiwX47
g8JngRcJsFgQ9VodQfXCPr02y/20PD6r9/GX2PgWJB4w1nCdZATjUo4FQpp8nyEE
lqhVyNq6B/p31dBFlNQOo3jyJHSheFuKbIcQNbp2/62jDlNGh8EQw0rc7KSYvci3
+WmbPXTOi7JeGbeDa/b2nOaSm2DtaVuKtkBygQv3uJyJKRRmqQCME/UH/zedE2Vi
rQLvFl7TQubHfYtlroHFrhEaeDnmQaAwUTzeXivNGjVAK9MeAq9diQHHsbe+45Jt
GmsquO/V6yIfJInfATayno0qSPsx4ZDuy8ecNRh2zmFK7L9GxHMKR57muwioYTXh
M9UxZW/ug3BNJVCAIiTvIvL59T2Kl7IT8dqOguNGrlkH5q6gAalTTwM8V6foJgj4
Zmt4Su3Fi9wV6wR/4Yx9+9pZw6nk++rew7A9wtk7AhCZF6iIbR86R/J+/4M38pCi
Cetp32vNuJX/taEIajLvvct/4UxwswzGII67APvAb+DViuWxrr+vft/ip7aUcxaj
jR/FfOzhk6x/0fCTAerBFB6JbX+HaWPPmpVoQiG1492U65ay3LV9IOVnAGKg1Jnt
zFXC893XQaVr78rpdz+Y5XZ14sY66snrusaPU421A8kpUzA1FbiYqPGIh9AaYSSd
ODzy9+Jkg8JWaxnJTWqSi7y1P2ZRGcl+hFAR2H1tTMx8TBwZ6a5PT2ByLfP1hHhB
1rDSPO+Tpg3HrVvHGPiSzeJNLTdqYittS40mr3CiSw5CplaeIUstKhQ2lIHLKZ0q
CiQcQoi8nHqVBlhIedolDvjFZo+YNYlHu0AvehpGr56snltDTL9tC6+F3rXIyW2C
p6UrYPTL2DcPLfR/obRrdHuRwKD4hhcyn1onHyj1xc32bZeB7IizyQ4qNlxoznIe
3tdf9pdyrg2qFCfzXrZ1uEw531I9FKT7PBuOpI46O1SDShfORP8lPhV8dSuye5M6
FkhSuXe4TfZLurY4GpCWKIYBn+GSyJI1DLymY6zfOazKkrhLf/s0jIBBwhg30gZf
nrq8w6pb1FaeZfD6cL3Axi8GJv9gPxvZ7UFR9AOHKa9g0plr2jmSB4FAVEzLx7pp
w4L9Xja2qVSm1HjjPKXn/O0WS/NRf2m04WSdvhezDj1CmVX/FLDHBvEpAiCAMVT4
snOorAyyNPHXDRwv+S3rG9DGuK4sTuB/7UxVnRO+AK35sq3MudrOZYEbb99FVrUH
Ex7g5lfWIAS9hF5iIdIfStq1m1M2mcUs4ahS65CrGfLxQzX2xRTCBwQK8vdSb+mk
/QiOaKgxdtEfBfqAZghtTJosujys+OpTM/qupOLHbMInLU9KuSNq/2Pxj6y8m+Ob
/dY/BHv3th0X9rCm29rjs2dK/bfHtpKg61127xfTNE5SzHDnjwTOZ3k85bu6tHoI
kMt45m8mxZhgzugFcMmnP2+nyqu5SVEwhjgOSDszzhebYmyXkas1hf2Rl1ov3k1A
CAwDOm3QdTA31nx2Qxtl5Bj7uRX/UjIPjbrAa9FbuPdQL1B5sEj4ZCToVUX/+epB
6WvE0XcNb6aLDIXBluN/LGZtKFqhHaE2bcB5fnREWPULyXgzGk/so+uVRSQ9USLU
6/nwwHaCQNSNj/jRgarLKIiniAm36Sbl7hxBfcmepuQd3FXZjdJ+UsKnTAReT6PY
Srs/16WJyL0TFtFZ0gONTQLvm2/c+jZu5+q+MB2jmb0/BD2NWVNAtuQSFWjt2XqB
96JWc8vTGrFfQyzcwyDO/c9ZD5TYNsZQWtN/wSDJsoAX1DrTcO0d1y0ieCGh5APl
figWA/ZZ8uQbjjYQ/CGIA7HEUhuFcmElQiGFCdbVtC4jRzpAbVudlHFC5DDIqulD
8f6hwYJ925AjE0gJ4znsZdSpNCxac5Yiu4cDUU20Nhs/qVOOPAEkd9BbpDTuzKMa
CUnSVdSH7zf9XZIcnAb1ZuwBWQUbm3lgCZv7TbCoGisB79nDQjEFB29ltOjFg7p4
AaY5ncjTd/PGAsZ+BKbLOhYbZwf0Y2A4XD2i3VSYFVXCtezle9jhmI1KxMLPDyZ+
5jWiSZhK1DGUl1aBqKTTbfZ5kwz1k1JEWFasGbZeN40jNYjJ9KzingqCdITnITYG
ScdXWO1su2YelVmqKY84eJBB8j5i2WkJ8U1FuoXJzDpWzxyu8FRz1o/Nawl6NHCR
A9gTCoXZzcDgiMspp4cmYZiRPGSwxBwVzf/b7yj6fvelFdri3HQOUtKSzv88lU8/
t7JKH1Bupf0vESIDZyib7zreLblRRmv6y9NL3Q585PFKREdx6aVypATP+QV6xm6k
H2t2OHOMWXvqKj69G5a7FvIwtydOgT0OOBQKzJzKiUAeC5XLTOJ2lJeEcniwC9bZ
EOGsAkW9UegHLE+logiGIlDKcTf7YLj7XomHvJpqviGkbnxMkzrHycEt5F/frli8
YUsDc8X4PfKJ4vw7TCjcWj1jJhzFoMdkivD9NTvgDy/Jwe0cxjmr+SfUlcN5JENF
bgiMlS87s+8DqJ4/e9yGBHGGub86KjiCwpmE5biko8K568oSdW30sQkJXvQaDGD4
pViOYg2hSvQV8epf4mQ0qpC9NcDcnr5uiF/1sBxbbHf9MbnE2u8v2o4CSAK76qwW
svyYNVwn1s9K8cnaiB93VAMrPuEmrDATeTdIu4HA2k8hconmNY3I1hx6QwBp0B7K
+Yb4DmEWoPQnB2bJNE4W4lgJ2RiteLiDJ5Zcdi26MzzkLXZBxpXKK8rBuPMdE17l
okFZN7Erqa7U37KoKGjYJ1aE3VPCTBCBNK+qSZq5jyAIW1jjelPrvcv0+b1o6pBd
elzfygH0pdN/dizgFfHrj2M6hNh7E8HkvHYPYC+GLlqtQbG7oWbBcHxIuUi1cKfe
pk7V2YqtWbEjk+N3Hp7lJQ5oFucttcUDTeuTz3aKKBx83NDnb5GJMo4Vem73uvKz
YvAh0zDcNWcClPRQMrfQsvd4Ri9r7zeBWSmwmsMe5ma5PGJjz0gCvYGv7Be+2N66
jaZbLLRqI+28Fwev3QUmbBTBTgnyQ256T6v7YuowD/6w4Poh9bws9WHiyRpLni+O
gpq2XzOWYI4Q26AwyrJP+ZTwCDrb+aVPy9+iz8U172lxwy+9GmtbxzutTzri6aLv
5q8AjslF56xo+EuH38Bv1RCJoXlk5cxr6GiUSdaz+SSaBnp4OUZ7rNzsUlmfsIBM
1L0qu9mjV/IUqAdSWA3mGnmOW4XWJwLQr0y84HLn15RSJPpjNDecEtNgWLjqHkmO
r1PNkeSKDf2kHaVx3Ji3HBrATj5KsIl03p3rzLg2EllA+Z/JMveBjHHY7IC5HwPy
uUX9RCRhzaNfDacYk7Jn7qB32RmO2wmoO+kOmkX9FS4fI/hCnrZeIPKgjc2Yvi0I
RyJ3lnlyM4Fxj2mKl6aWeBdiLC4gA1QWTU1hKoIYxptGywBNCoKWkxs49nl7lSTY
TwSyqEcjibGo2lSF2ZL0pH9ZuauxDXYG5AMnZzaAhvzmTmmDh5xCjf49M9ygrYp0
S9wJ8rkb03jsHmSElU4hhbE2e0iwfQdHDFVM75J+gYGGmF1XfW9iPBepuLqffSKM
af/5I0qUbwkIG+8tjGbtus5TRU6gTq7Dqi8MQzruKxF+0m6fiFrTxaSjMs+Mfbna
icxHaqwHf1QCxlNc35hBPMf+Sx+giXC+DNceXiu4XsihgzY8foYxg93vcjM6Uana
YUmTqKCbPzbcCD0wDdTnGm4CizREnQMEbt7Fisvx4l5gKOHi4qh2w6HXBdqO3fmb
qDSx+LZqHWsd4NqZfHhM3Aoc1MhxxqEky478HMuSBoIAvJ33v7yrix+I5I+bYt8c
TVcoU1hdxiBAJqHNCP4Ot7ZmPBvFIMH1GchdcKEt6T0tRjlF1YWAhISpoB8i0ARd
r7QGrVH/f63w7kbWO+8lAs5AiDl2muSNiX2AgHMplf4ek0hfKrmC3SB2eaEfO5KV
NDFCI5ynk2kXbl0g+BL/GgwfnqqpNZPi4Ggx5tdUrtPlIUCXP/D3dLdrb63N6Ctu
8MucG/qzeBuCI8itQZwCAEBsaw8/pzfc4VLb0PnUbQEcONgEmP5nsco0tP3qYkOI
jdhDWYbKPjaRSqxMk1wJQ3REIfLOxnJjv01vj5awFo3+oNT0E5ZAcStXnI2/JunU
C08Nzj0DQot6Nqi+MRAI9/jNx1L99UtvTanYOzKkzQMGJijh3ElEcMnG4wUObU8t
ohSZ1/Z89lYajmWOhmdPaFuMJAHr6BZhyiCq3/SODoN2QIAfgU9bCEmFqbIlBWrm
z09uhJgUNKew3hLoN3FxfGQfIH6T4hS25IR69r6kHC/3qjWGsWI7k25SrJuHqPqE
+g9qd40MSz3pMaJIoedJOyH0QTcsEvb3MdULjfm93GAcAq+1KHWlrfZH7Oe9bnPn
7sm33CACFAB/gOiz1mA3axCJBNiNzKvs0R/nXw8EnBAxM4UD9tKf4yF1gyLZxAxw
a6BxGzuLHkMwIRR9eD8mO+UucYVWKDknxjfth3Sn04gbtnxGLs/KhQK47oQAtJBc
SLSlOd3TQHx/Ls6YgLk/ZA1RKjekhAhDcQ5mf558j1Qd3Xzav47HZg5nsEN4FVQ1
ug27qwwV019Fpua2JqgnB/e1pca1fP4uNrb0VuVX3wSBrVfJViiDaMw3l+3VOwjs
GvMZIdRur2sTaIKb24gRZmC3wvOE2m+fZH8Mp0DXv7a16lPCBqCaZ6TIHNeeX8kA
EoEJcOq3+/0uO+I5xZRGxvIxKCnHWM7cQDBwUet3prLBn6wUFjv8ZcEz6xfCfiXE
HpXEMbEIv+Pgs0s439lECkUiheX3qO6FQrNzHQl3Dd4+qsNWowEpXkZrAbDpLis+
BryMbTNAMyvShSJksqrbVZ/EKVmt1M3WnjGj+H/fpFfjY/HQPpRcUa16SPyj/lJ8
Uh8eJrCoIGRlD4LhDlPqpE7y842gR0HEv0L/JvfkHUjRbIkQupbgq1UQ1lQYrk6J
O0hTdljvlrN9vTqg5c+OnQZO+N3K4A2LJn+QubZD2fOxbEVuoi1tD33rNylL+4wK
GKWfbUrvuSfXZWQ6HAOQD/pM4OV/t3sBvJL0oItlT6JJNpLBpndUkJwM6sKmV2xg
RcG1Azz2BHeDtU3nTuibkt4TfAMWP1YW+JGFadqIkbIPvjjHBgzKmqaGcmRFJooz
SKS30XruhjnvWtU71maDJwgEJVLBBIEg7U7dJWweQ6wmztk5RuUrlseJTbiRnLsP
x9Gb0kwM7pAXHO+V+c1Ms68qYsFh+r9nRRm+6OoNZT/CF/5bWtBkm9kTnpLQIvow
O/e3G7K3DF3w7NFcSQ98zbYS5RfqZnFbDmNo+HV87WmLQcRIP/oVgo9xqcoMM+PR
HvPhtaALEZctKUQF0s81ZAGjokw67B9P21o1U2hSkdZJk6k2f8OZdJ8DF3VJyexq
GQN7ibvMKIjvzxDiTzIiU29NUb1cLDszx0/7924Z+M2ZV/VH2pbxJ4QxeciFBKXi
NhVnZfsWa1flcV6HxeOfWLxZoehgqc/ojy2xGkFIfzQvNyf/6PDsMCmYve6p+WI6
4dK9JKYg86KzRHPyEe0Xb/C9E8aijoG8q+K6YQhpVeZ4EEJ691ZraD5e4XcHPgvg
JSfQj3wHMHY2GPdNJXRI/1t8lPsjGKnknqSuoA4zHmNkhX1FF0GBn21D/FVHwCsd
v5cBaqLdS9oQh4ZxKOsaBzDlNQJQaUzNQ+G/iOpRLQ6CFDRhSOgfHR7w6FFgYZDl
7t4sv9P+7eivwVeCGjaitjM+7yk93v+kzHGrWDyKczCmkRHX55S5lrNkGzYpYiAI
HrSikWT9ut5QR1F2ZBEfQK/zJiqqF/WjHW9HgxZO0W/ejKGDCbN3whQfqiUJRywu
A6Y1ce4IWyE8VVAEbEVUyhjrVQGVEP88I8FjdZjq4HCdz5tbSrqBEukDEM6HtCBa
9N4MEv/keuD7n+VxM4V3i0ZEms8+AGddF9NORBD39qHp4sjQ/Qchkg3uKeHj/fot
mwlayJ3jJGCNQ7s506ZDCcPpn3UpId7VCUTGhutZqtt9KhuclZt4dD+WK6kJ/ArU
htTxJE4W42yB1SPhtawfCEA+WXXV8MTqfOp+0mx9LHDiZ1nY5u6sdv127CVUOdlP
zfLBGyw4c80GnjTdKW7H4D1/3vxxTZsbD1+l6BkrB70XFpRQK/T60MTwMweWuIig
U90DyT/vzk4OI4o62VqzDJWyk95FMlFsfYkUlh8U5KkHhkE+WJU3Y+4necFUv8ca
7H7LT4OtEr1zDDExncchlM+Ezj9iWWQsOOuJLFt3izYj3vEw1zVnc+UvHeQlaZqI
EXir7NTC77r96nM6COKN61ADyqpDFnRS/SeX201SAPUewKpFoasG9Dh4oXObjU5s
P79WGvRsnA9am8YzON2bLFZBKeeq3X+c5gwFC7N7xEVFhDWi+15OK8xkC6whyPln
efsKxnARNoiTPA4kKH2Kv1SY/AyYee4eueA/QVDnKr0mF31okz8GNHeveElIdAQ1
e9aBYW4igG33XzOgUwiJThNUmVFP9uHOFeWuE8+jrsOZ2CpzXc5YDs+d/9r724n7
ZjvWZz5lytyDpSr704QD9T6bh9ic7qMS3xn8c12/nFG/DxZ/5+C6zFp3IkRR9tnf
ld9vpbrs1W8c/EfHwzjPpUmNFjzpqSOK6/zZmhRjxV+tdRJFVMd/cJ26zWB8cn8W
GrYuX8VDaz1ogmfkCIDUJo1502+7dXhcIDAdzArw+EahdlzFa07IjmJ/5ADN2kHq
xMps3ITsF0Xq1KPVolcEoeQpORdPj6MQ/rzXkypEhi/m3KHCSpqIi7d3GzoJdrst
X/qcEGshMonemw3UQ9Xds30EwpsAcMu/azrHNs5uKLhAZcthCiEU5XhEO7zYlzEB
FqhsdotgY4UCRtYzexoVVS/N1T2dFUEh6DuxxsU8BsPCzcznDnO8E2/chouoW33j
NVult4csBZu0w44R5AXa28+NW39RfdwcUOAKnnJHckE5wob8aQo6uIxdHWCgLCR4
RqUD9Y2lpnBREOYW+tN7Exa6SsSLCXpHDoVEXpVY0Vewg1HB/VhSFzq+o/ZL+4uI
AB14kOUv1+nM/U6toUXNJNkldf4NsIAY/qnh4to+BkFjQPRbswNr1+hszMZdV6wi
l/LP7Nt/57JhNMGZw1idYQZ7Agpzp8346OlLRCVTcR/uOGraCTh25Nl4iVSSu6i9
6p+MNEaCB52/1d4umMJaRLNcoec7h5bWGrX2b37Q3MoWq4NZZHOp1Zj/E0xMCPqo
kY6Nk3RKlevpd7aHy+IxArwmcTZX7CCu82GyjWHXI1ONDV9CvokXVu0v8JIAOQR0
WWfz/r0Um59vPx59KcDKufFJ7K+1zIJqKOMPaH4rhppzWEH/7rfBUadPoSQCK+eA
5I78p27lhP/hxxWOmdNNvw0Z7jXNSIyWQS1oYtWlpy4XnCKB9qNqTCkmAovcOPm4
y2n0H6Ki+u1WCZ+bi2ImIkBoA5TKBsGqVvs/41JjYoQlDDPY7qwEqf+eiyKyYYtH
1nfxLEGh5OrilH2UT4txdX+S2eAVOMSXJ7q9KaIS5rpvK+TZj76KyCvdPaGcgH1N
kKHYDX9JddXGB5pmyDPTaZgXBSQouc1ugA5q6RSRP+lnbAUilRHzbEXvk2fKmc+Z
1A1FXGPAyejDoTMtJG/YtnwW54qQppMagat8nALKmp+tZRJA46D/z7y8St0+kPgy
fE5uLuvzYpvedFTp3gV5WY1AVyEKWdqF1xLb6YqRNug/hkBgooidwsdQt18ZkUPV
FqPK/9RJvrOPzYuUy9MIJslIhbNDbbpzr0LeM37A8gA8ltjTd53k8Jqa8YD+k7V6
hmd96bf0m7tlndkcuFTsGtrnm90M0BoxOY602BQUcGqCI4bUBa6CaSBFov5IOu2A
NLws4NxywqmAJwpRPKtpo01Dm8HT4FclnVHqJZodSo8fn7rEnf9HPefA5AUoK2yc
0CpT8gTLTu9cEwyWHAi7KtWILMO3T4jxuU5QJha45D9K6BzgOEvfzFoPMK8GhM2y
4GdmPlusNnjkn3YK+b4l7ftVPgCo79T15xT+6l+2aLcAWssHAAUHBd1o5AfXxsCc
2DjMJ76+DObvoRkTmfZz03CznfZcK1LDHDsMi7dRwnv+vXIbCnZb52ZstBIJcfdB
SIYPyTYfpXg0MYUXHM2Z/PeO89/2R2jlOQ7CWj6UPiuozg+Hn2Y7NproV3HrZ8FU
GinRl07QfzG0lBkA6r1aLdCVIE1i8zVw0D/gJbtNGuyCiIGnHtcM1myUx+yY949d
9q+Dqn9t85eu8/DXzGF3MM1/oPphFfbw/GlBkfrp1do7IeOcFik57Qo9Vjhe6c5F
JTuItHHoSgYobQ66gKC7A7c6qK7HewU3uj5CpTjBG7iC7kBPtWabAKOd70whL1nq
EJbRpk1VTJWwQNqGopC/Ul6pljldR7m60e3RtLFrVL3+Yj94GPWW1yzEWuk2OBmy
3ORsGzBNCz9LudABRs4vTIjmcmlcb2aq3vQmD13qJIj//q1KovwiOy69JPoq2S05
Lxr59jEjxKRzyESevVw+iaMLP2YWUH387Lv/XpW65IJlxtJJ3qA9pTWLLUgBzEOY
mEITE2oPH/8iJJGXNUzma/Uo0WusQuPRrXD4mzPczo6+bo0xjIzxNjA5adIVKoEE
GhKO9kSri04Wv3YJp8v9IibEkLhx5YTT+1+AA4onOxd9eKhjDDhswXipl28CoRAA
rAm7pnRm7H8Q5LfUvL8ZKKNdLnSHDY3REgPDLSVkUIdFoC6jcGw8Vq2D1l+hSzKO
rNHwibYpB5NUgtMTN5geHCYSycbgTWD6aQ4j6uuHn/RVmDRbIA2v5Tz2ofo9B2At
/FatPFlpytlEsS3oCzQXuLXHbKtxdVmoDgKUyk2YrkOwaeH7ix10QMOZwsoLaj+G
mF9J7hL/8Rw3aLp5c8bUY1XQ2zmJuVzPnSIek8CDUVC99IX5cTf+12uqslHQjfWu
cwJFDgfWwctMi2dj+A+yXCKLKc0SUFeeDV5kjiKM05DkLa7TuRQPsckfd43MRS2M
ANQW1331IE+cPi1bxpTuajoxfnuXzDGvqla89mTNu2VcDM8/xEnOFZaqEdzvxkJZ
NwSFXabuhsnJ20KUX9ZJy4C3hYLspB3IyqzA8YxOOQ0hcSkUat6lwYbcMMSKNaJd
0KmTnsS170TZpDa9Pohd6SNhssC0TggZ7k/LOJIVc7QEqUIlxAR9P+RPyfBqA744
7QYCpI8Wc31yMpMV4h+GpLG2GMEzxKHNPriOrz5+t46EHCShFNfNzh+8XhJYhVwf
YvkbW6G8D5phh6Dg5wowI3EXdqSLzAbpHvS5dkTfIeFcctG0a8b7m157VnnMI+l+
LLCsx/hZGiH5JkbMVtRo9He35aAjDkE7y7WNTJ6eQrSLGGk1eStAHisaxmgueUNa
rkn3ZAV+gPiuUZWS/VhRu/udR80kp18yt9hQCjJLCHqCPcToVBG07Gc2KWnRrSH+
3uP+5IWZP6dBMDpLIBv4cVnOwro24/nJYOeZpAmuJTkcJdFwbsbm2i79Xz8juHBr
M5LdsRAXUiVC47MCfdqssAFUZiy0sYTUQEgvs7pVDuAYHDNx3IwyeRlr4nR4klhd
rMnDVXg6F48owNnK2M5fruttZKTpEZ+XzoeDh5Wu2/OvPVq1U9Z8x961IzNexz2y
R77jatS0pY4KEIySzKzQv9orMCesAYWNGrQvnMnFg/PYx+YIpl6hD7PyQTjXhS16
k8ybImZXIgv1V59wrXKmMTGh5ArOa9IJhrUCyN5G2Us93ALwTahJTZ6B5/WQ5fkq
Q0Vl1GnJxKpL5FuZ3F7QjMdhIKxfNPTeZUAcguQv2fdTcUqTJSLPyVb4YXq41Ehw
AQpzONaruxyeuiBfuyFyY5ea+OvcacpLuwLfcKgTd7OnpRQY9dqBIs8QYMwgzmTO
AkaXYB5TY9wf4SEqhhH5hWIJOb/tgfCVU2LMGhkP86sGSBC4ietNiBIUsiq2BCqG
hZJf9UWfWIQZ3N6uJGyGCqIL4QMV6UUIr/gGh2nQUecA55CqsXbkWAeiEjof6wfI
IZsnY1sQ4YBF4W23iCHS3T71kFNFzoASr+BB22CgLBJpAVQ/9IHOE0Iw9lkjek/4
7aPZTwzP3HcBlyQw2wZOQ+UA+mBNP/Bp8vlqKB5NRptEx9RRUq9uNo3HHsYbDqF9
IIMnqv2g4RKm+SPOCCuU2SarsVFrn3+/GeTKEefU7JtaGB1QRw8Dl0LA7xBC+80E
t9kJDNMTbMBUyXRNbTc6bprrwAKfbMQ8HKk4toCRBAJD7abCOCIEWOKgcjSGhX03
fqNN9y3dULR0HkYieBVwkHymuFVzFbqRuzsOhmX0bMO1Ep45p8NaNJU/rLHyrNzz
hu71dgj9RvBCo1kf9Qwlv7CyACoSGgMgsdOCOT1p9885dlkZMpUF1GN0C3PXf6J1
Ak5CoBrGay8XjtKKv/AKckk70b96P7fPL1qJzsfFIFnhWaQU36ZSZQok81zt5R6U
NpnSuYrfcgkyqVYmypxBkLJI2kaVff1to4UAuZyffweo2NRubm/fyO2OFqn03vVe
XDkdKWErh2E834/YWbboJTvDYZ5n1o+acKpzNLytIE0NGeeU5pfEDAbUm6NDFKBK
f443lyuCQCfaE5EX98QPoeUnFRzRF8EOlji0VQXJIZtBVTTV3OSjjMngFpB+KJCA
+k6PAJ1mQcdGW0DfOcnEWzMQIId6jCmnazB7rJPTIULgOv47eYDYTY6vKdgch9MQ
/qUV8dvhDcHuxniX7elgddi4ZikPA8WkZLwOxxdZwr7ZVd9rFzfewIXFJUKmWAyY
ogVXvNRoqLitaM4g+0b2LD4kfVEMfaawMbto/ybmMTiKAZzH/g3JiAA6QGa8zHuX
/DWT4YrRb5DT2XGjB5niqd7/XHiIVv+UQUZ38uCSlYC0Hq0wORxHDfyr5OIKsuLx
gwN1uQnQtDlpcvnIvkLL77Eb2Qzh6UFAYHqrbOkdT+tFIQtXZ7aysFF53HX3rBqh
3uPGmaAxjNJ6xnLEevASMwb1iexzme9RJwMrHyYZH9Yk5uMN6fpznU3UWBMnOzQW
Vf/056ENxOnvZs3jzoGXTVPACCsHizmex99Af2xsDX3TU4XxC0JJzQqfHhAvJXqQ
Oun6dfPdRBTZVunMSei8QCIXT0G7qdqo0Iwber9YJl1fM3BAHayf9kGsbVbGB/FL
tIXrTqDKUm37Mwh/Cjzt0UMzDzhuSvkrqbXEQgzItGlC12o0Jg4QajX1+1NO+zu6
aLHrslicvR70ZuKfwTKyKWfqvWSOUvA20DfD9ge2x0SgCoYHkjua55ZlBWhuLCOK
YfD/ZuuG/KMrrgvGtXIbGZsy1Oa70b7hDXr/gi41qRHbolzS53gohPV20Bg54Ngf
YgHJoRhUFAzkQE5mM5mLsGEz2iLfKgSDrQdkZPuf1whtdzaCacd/9JVX1jPObu/D
kuoY8UynsafkoH6DbsoW96ndyai3DCNEqozQPKdulrF/fSncF3K6H3tKyqVjoJG2
NH6LTuZzncuSWaX/LmQDM4qybSAR/4UtVzNXLqmxe7513AqyvKh0EsFKpNjxHYKz
oZVDg4j8hfBSr8WQ/ntz/dzHFa5GLZLSYbZ1qeQOny+aM0xOEJaI8bM7ieuQJVqJ
eYBCOYcfZjVAzLUWCr9zSgDXLsUuchpkqcxPyeqUy+hJ4mcol7uuJvyvSpfHnNVP
CcFuH70hr320idTJMWQWL6pOGeG2+f/EohWpzRTGy2k8KihUl3qYGac/k0JU38XM
Q0gYQNzf8exAl+HoCYA5BvKEh8PsOkFIesjuo2GYF9Qv5/OQDlhJzW/sOSwvqAtv
ggo6TOQrMdojNowZ+6gKYJSGBG293YTgKEcyJHdTm0bp2Xlo35IYKZ6qG2ykjD6+
qKgTNNFhIeOY+Z8/YhCcBgWXFienOQJ+hDWIM8KkLOP8pLCpa5lUvjdBaRqYO4Uv
Q91DV0+pnhe+kry34zD2+NXebfPlTuvqYlh4fDogYvhsrwGQdRPTifP/q8Dh9wI7
WYOO647Jzy80ASbt1LiOeaSsNcIDA0I9ulfhkMHWQ4Nznspfzj9tpoPH8Xi6OYj6
xgeFfXpgpzukklwwy9/3gcu2foh2LYP0VhVO/z353Qz4ULvx9+FLLzhpM4fgLfg3
BrGJsJhrGpGECZSSy5qdmrWEfhJJ9cFgNSokHRjGkMXqPiM7+Vg52lQ3U1rwhDbe
kETLLlVgdz9pzSVULatDygg2Dq0C5oUUpkrZwNQaivtQf3w5Peq4UdWjw9mMX6og
AkzsZEjLN/zaH5fM/jYWMh6FOc/5NTAbomgECm9aeUz1l+zwgcB5h82k2nSUzzPI
xJv1K99h47/MjufS4hJiu3FDY2+j9GhLNP6PnjQ3We3ozCmewoijTMDaQ5PcbSQ/
7TKlfwyxXRPhhH3DL/y+OcAhTrodfgrgDVc+CU7T2IZr60/LvU6hABkX2oc+VEHN
GnYSnCyiau6/JwIAnYZyGVhI7d//Azm3d60O4vbHWouoAW+/9wBhpLnbmukoB+vH
RWF8TfrTLz+hBmn243qcOlDV/lJTlboMYoF4uWmUKcO+s20+PwQiOxr3a88qd1LV
q0vwq+GET8+gsWPb4Rd5Ihv7yzQS4eqUHimR/yHK84RUC7ipVZRvbluIRYeAz6gM
28CaRGCW4ZnatLHYetYqmbxMqmib3TiK0eaGXH7lpuclw6wZVQF+UhBrBeDuc49v
PGNj14i9/MYVq3SObnHJJGJEGike+CloPQKDjJoDQEMUUi6UHA5jWI+y3n+Oy8bN
DV9rWoJRIJH25joIgtbqU1mvl2gBThJCpTUGTY/BJWWhc5PHeflizTEvydEca7ZJ
/poXH3ZyWDLU42GNWc5MjxRQNLu7Ud/QhiLNDMEJfCYmH5nzebpN5e1uENuhaDW4
WCYWkVfzS0gAFwohUT+LYz0TnXtKyOcOsfRtnuAPpurTtOIqVbDty5MWqrRlQ5A5
oDIXIh/jKvBKCyLalabS2UqZzXgCLltZYUqxV/RT1nUg0p8a9sPQpl24O9toud7/
4ebordteGsQ2urRXBBb+Zy7abIQYCmuqzryjRR24WrEQ78/RHR1hCFQh+xckFXWY
TBwLi23aBFKGfKEKWc43ypVzhRBg8gIv7IxyeMCsQIbqs/yKM4DVcPyYM6bFd4KM
hg5MalpXdWvsWjebotHFAnWvJ6LyuIoZ43v+iLEJcTY3bm1aGHbxdpCvnXsTcUt4
0ay0epHOjOnunV5pUboYnDhQUiBSy05WUtI7LzHDGlWuvot7NLSKaYSml4QibhuQ
HR4J5/uZpdYVBa+lEnAIvIsIFEjaQKaH0KVuQVG6FoIeRMqWJo+x5Uui3FQU6tgi
tvIf7l4qYvkp42xHWA/3e/ptHTNlP/OJVaeM2wbXoz0g2Mriyl1EIggGJQ6QmwqT
Nf6Rjio278cXuzduRzUZY3uV5LaIxTCt1Ric10zPkUKHNLUTB6h7lnNKhwW4ANhh
+njXouuHrt54g9sbaVp07esq7lAjBrvXzjvffAwx+T8vactnpKqu3n+oZy3GGiss
YLl73Fl30okRpgMgpvL1EPKOXkOmnS+A+NQkPWW4AfzQQdH6LV8HHspB8EfhRkNI
5psxOnPOLExGAUSqJGPA7YsINp1Gc2D5j3sgLTftJB8HPbayo89JTrlHKfNacawC
XuLzQGkHdovBtaG/N7OhhEzSCOEMzUcBhRAtE2h4/OmEcr494LaRuvoPPN/0PoGU
5ClGLtWXqWpJPrGJEtaFX9K7gYdSMTkGHmD/yo1M6XzzFl4yHkCvcP/J/5t+Df9f
i7catHNM0niuQSHojMYZYTedkNPKF+tiNrjM0XSG97dh+OqtRE1P5XrEUgbm76vv
Ckzxa/eoIR4j9t6fLUfZQ8Q/S+V0caTc8E45PEj64aqnORtgksdZb+GzpL5ywyTQ
g4VibTPNibBIAWrquZNRICRk9zkQLvHbJZT/x3PnC2kelUJPKD3Vve7wjeNtdRl4
Z9TMYq3aefGbn7V7PmThY1Teh3he6Eldp+RHdyhiERNZElDzh3orXKI4/uLyrmM5
2qIUoXSwu+EqWCpUoa4rbL2uUCXCesmlGDr8aHhX7YcypPhZde+rP5YOiuagPVtn
ktyzvDMbvQKh/NOS/eQ7/SZRyDT+zkGW42RgaWqfzGLnXfX+xoeYw6VfhZ6MS+dh
G2r4o1irco808F+3LTdWi/iNQVNFPNd6iawMBIkH3Y7GxHTCg2CB5aAfEwpZq4fc
H4TOZHyU/8QR7zNnHYdtEUydllm9OkSI09xsnWeLfQaGn/BVNmIS2d9GjJfQxiSr
OfLS85AsERQzoLFo2AXUrrUsbVD9/fXT8iPLK87MuofgH1hSUuDG/udZbOPYtI0O
PWXI5zhjQEcCAUJ9s088nnc82DYUw2FsGXj101q5JLPD2oF2iCWis72Hr4TMxK+M
oX+vv4fGm88Y/AHU0rVm/8UyzuQr9L7NOuuEPP6Lfv2rJln/6MHCe9gsBGw9TQ81
CbaFPs42pHSz5J4KbK7Wbmu7Qi81wFR0Vu0EswBNwCeXlTz+RR1YqE1aWmAHYtRZ
jV3/95XPwNjFFZvOFsZ+UK32MQLtSjoh2fdoQnAnAb/4ErOca1J/1CsRrZz85XLC
tbQimknpbA16zFhH6vWhCr+pC/TFk8TMWw5K7IqcM5NR3Lt3xBQk5ReXqyt8PwHk
rXa4gJrlrU3NoChJWfaIwYk5p4w7w7G1wT+XAG8hvXo08JBmBb8fPpXZ1B4jq3ne
UHvH24gPbVY5JUru3rEpoMbRKMFseZsEDBN9t+ZTIGgLfaDmXJ8LcNIAn3kNDLv7
Dfl5CotoWUi4/eukARojY1DmICtq8GnOIZkGphi5iivfPExbORV9LbJaByStZL+V
rElQKHms6BqKcUp8u47bkYVNCLkTyfGd8vKP7mr2v7S6aZiC7/s3vNt4Br4teY1m
kN4HQ9yrdS9VUDBGkNnDxTOpZoAs0v5L1tmuwdSOu34M1wh8YC35XrPfTuUWV1mA
7WMhMrDqoG3ySi91csb+REJ9iv/yL9mBJoFlt9Wx09RrIde6z7kVnIUuIKPYLJNX
yzobWOZ6T0UBfY1925rJ+v1Tt1XhiHdsXFQSvs5Ogy2S8+RGtW6ZZuGn72XdSyeW
08pNtzL5lQyug/MKP/BTM7X87daI/+S9MqkLXszfj1w2c6W7eeDVYXr23vutQg5e
S/4IzcWVarqLuVWtT0zBcYGKDdVu0gAses3NP1r4V6IdwW/NV/5qSckFEK3XUcHs
bkzxYOiz6Wc/bV3JZm/i/98M0KeMQaMqt9ibbmPj6PmZQydhgamDE+y+Jx7NgP5m
4lkQAeI643eKukMd+HNUaJxDv1h+L34T6o5vFrQG7m5rm0ZcnTJWFoSYaGZadVbH
JcQaNHTKAQm0aZT+/LIaDy+V2PUyX9e2LXlvEyajIXPTYgPClZ6E9rhHpXKhAN6l
lbcx3sgTGwdU7zt3nrlEEeieYUz4X8r661FsYf88azySySJzZ57PXvQClgM+mx86
rJPSGpcFw8prKeWv+5LxBFCuvWzPaj/KqglOdHeb3amj0+420KoBOmxf9OPNEXb6
2aXSOr8n9lw8R/mI5JuALU4NW/DFYGD+r3wl867JcY7uEQ7mNRVBtIn6F2xMY64n
O38nLCrxNSO8aSpYjvXHDHASPfqToVGesJYgzpq1UiXkJOSRrgQ3RgqF5pPkS2Xo
x3jXHDYyzYZKoosIXULK4O05+Ei2htnrcIKr3VqpG/Zl4fT2kEgVoM6OzPW+K7Yz
2pOPZEgyUMo2P2YIhNWFK9ZVQ56mVmJ/Anw1m18CvSib2MoHVkYQDILo4zdwzUNK
KdxybO6SgEhm7ezZXtjTX/ZxYpLIpkO1RgDbhAiYC4/CA1kXNj4wLYUkui5zdTfm
DcOKF5d97emgv1PcXlU8SkIOMiiY2zuj4Q/KECxJMwq9AZpf39axX+dD3vJS52NZ
W0BiFTA9MaukQv87F41znadtEwx4deZuVQayR4TnJnHMO54GCJQqpH/flrbearVc
1KUviLA2HS1TafdejBlfLSKF51uwn9EW59w7JdU60Xdf8XceFiO5MBHAU6TGaDGx
BZE8HiPFW2U0CueYWaV1pzXVrlfUceLsW/ilbJf/qeVIr1dS8m63kBw8ysCQGf74
1WAJWwYbR4MD+sKKnMloJfYwEVnDWIerx0pd578pU7Y+SFzUPU7oQxStOZNSWUfY
3OyiuYEAQ5wUvZWZWe33uUdssDBzanDewwtdptgAMZjXR3W22+kmbLeDHBOLtZEQ
uMgkeNjOJNnTJML/87t3lEhAJkwpRvBPRjp34NeUNWeyVOh/dRvq25fvc3gmVHss
SoTqSH563xAM+O9F6wDiNMp6EA72x5EW3nLMYgBSyba8pAsh/7qjQS4s8As1hQ3Q
6dUnW54fzOJzmIQ8+Qp9llvkRDkOraucqCMXddiMH4Uzf7q5gnBevOWS1jVMk9+4
GkKFoa/ISXchYxIk4dWWWmr5JJBiet/59Kddmf6RP7dxHTrlHNZ+76ZoRZfmjqjW
JdqX06K+nOLOfOwFgptStBonlbIJuoW89PQKBjttDSNj8N9iJJlKJnPQThK8f0My
4JxayJ3m/kEiL2KAvS3wDsoWUsVQ33ND5Tdnld1NlRrZOxhmZRT5L+zEsRO/9PQq
RH/Nr6wl62WA1uBQcNegZ5fxjEWrO+CID7lH33vm0nn9Snxgg+qcMYuoof6+0Kuu
NkIegj8ZfIO97kEHlJsd+sXNpjD7uyVzCpTDbu1Y09k=
`pragma protect end_protected
