// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
C6u70iZ6e5JByK6lduRDXlzCh7Bs94QBH+L19AHx1mFN/na2XZeIq48z0Nd4C3YjE9cP1h2eNFG3
cqYgE0WFrZNthj6mWjgeT3FIpIiKGsP9EnaMvB0t8F7FFda6c6RDzqN+QMAV4Zqw/0KzSRj+UFo4
JOGKH2rse+CWyAxggGUswCAdZdJo2EutibzlfVRxi0cFnF3K4MpHZL6TFZILYusy9v/t74lsNC9v
uSusFhyA3DiH0W0KdKfUl78C+zKMwzeYaYeXVwats2L9/wzqSDUVKnPRYB6l8cq8uTZsIbwZi/tr
fVFxM7yOd5WAILi+xu3RNvlA4WP6lwIyH/NkVg==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
VvrF3VM3RQ7AU9FFkHFYsy0GL0FbMrDtd6xgjyVhN+MHfAdiPasP14FW/mlvbOBJf7lQ6LGNQFZH
jMTazVPLiX2tekqYc9ylV8LRzIRnxK77O2xXJHu1hs8yt3thKz1IAzxj4ZlTPlEDt3AcxrYgYXWs
BFzubk32yqb8E2PlJrSQQrymLC6WnFTSxEMTq2LXCmPUsMNh/Q85XbB+cCo0rsx67+fasybx9Uq5
9C3FKU0j2W/vDfgxWuyH3MBK8GcBeDHg83ySXC/uRpHgvg1eMg3KufYlJaytwfqPuLHUZ4UFZN6v
jHLaMOoRdeYHGp2wR36zYFBQ9M0cwFKcPJYtFkcXlXZFAb+v+SD09dAt6AwQW9lAIQm84roIE5l+
E/tbZSFeEBaCrqiFAmYHG1AcNKHLMKKEZxirxETzXNKeTIUQDtuEhEXrH0MZKAXDKW1ZzHus6ULL
1pzrByGUdbMB1/8BZsfJxKTYUg2TasM628HSfPkrNtWVYyXxm1DnZgGxWid8JmgIhYN+UsUVVBZL
ntCVPZMh9aBoaKu8me/0R9Z0ve1b0FtLihhVmnYavA6y18nCWVBD7LDrXhpCVkMaelNzZU5TKl/O
ZqAXh9f2LcLFRdqb2BGtWgrM4AeB+MkJwqT/FbSnBksJiRsUEVbjrESi50fhCPF7ljk6ftZdObv1
/hlQ4/28FYosdBWDbbQfoaHaV2KSQLaKTIAsmf5lhACGVa1wx9vjfJWUsEaoxj+2c5E5/R04SIdO
4ME72Gr0eTwO1BN3+I+hFswbg9pNY4UK32ctzCm42mJezzy5sYP5PNg6bejpUp+YjbqOC/hchqih
DlZIHLzFVKlwAfk/dgJDKtN5LwU33R1NIo/UG6g2iyJOnwMMhP/vDNXTQjeONwT/5igsPUlRVU8n
j1ya04+Hqxxqgpv1c+G3QQzs/YTbzKNZO+ouUcjvvNQgMASfpkQhqms1/DR0nj3QqfoB/00Uvs5r
V+/CgdBJ3BP5EBNM/CHhQhxHc3wXPFzlzsOtfnSdTfmoDgycZK00NnDKg4F7aoIi9OFCyvyC8NYS
l2DVSuc0PTej7Bb4SboWPSNZjSYUxGEH4SZh9rmdPpv8R2g27mV2bhErtOkTTODoAvuz99/vJKeb
Zi7CBwoq+b4vyDl7UDMExH6JhT3lUtOrxGMYGnEjr1c9g4lQrkI+3sXlSiUDwH4pfOz0mTYt8HB+
m9NjDA/CPZQEMbAlVdXC5G/JfzB90yXGE9uqV89UUy8zXkDf31+OGbV3KZCYFZDmyH2tdkLqbiJm
X/oQr9xcgsZ5cTI919TuUAiNSfQggNIQ+YpCgGGaam5SOElqjVMjj9F7WmWar1CG8VEvYzPMl9Kh
F3Do7IkW0qA4K3G8C9dWUeIctI/3gxyJgYyNvz3KukOUezhIni2nX/DPxzV5EoAlj36qfklIWWHW
7CXWxjmldjpZar54cPmwQgPL3U9Foqt5FOoJNlUW/h154BfcGPDlaeieSRmHLHQxNwwlwghVnTg0
enOppr27on0HoEl1wWopNUSfOdPP7+0YXtWC1PZJ4ive5+sxnAXpm2LUEDfGXLKyb3MS8q463lbN
x4g6NxisklweU7ODF1lOCUbE8Cjt9+LJHqiSO44ubRW08xieWLPs4XUY94IGJNWs4x0avl+OjkVl
rLa80fuWUvLXsvXlCtjEms9JtosYHBARjnHEvfIfdOzxlp5wVWo58LEXVU8O8u/48I74Xi5sCC3m
XesAIg0u2mPSBGj7gUfQ1+F8yzSMDVedjJvEvHlEJyQrf+t5XElzd6dfgX8+6zWEptXoK3/FV+FH
XHrD41NMtLmz1Y+RXqL2dYN8dqjbphFDcR70lx93H+kkD2XY21n6ZqBgnXkJPbLTe2wJi31o64OV
4zWEyY+oXxyUrvcVK5NdSGingQ6uMtQst98DO3X8zeKeC7eIdHy7BFmFfWRqVPf2IHCsIh6FmiTD
9X1Ai4iEiFzWSPsOUnDe1N28X0CAYQbu69FuT7XsjSK7McU6ayQDHuKjz/r3fofzQB+LdX4Y9ImJ
Wtrx3BGJlBQHhjAyl4gW1tAm+qFsDNx/w29hCnjXlEEFLZ06DjUXOVIr2Jww9ZAZ1pGhFKwdHnqE
xWu0RWy+roo+U8hKi7yfAq4DHqhzBc9ub2yTkQo38MJim0Lhq6DmiWMfGFAfoxfgTwjK6AlNOhy9
ob8CkynXmvwhr1X3UuxcG0O9L528QEd2BHZ7vFWaGsn/8ffAzn8AdmQU0/vQdT8LQw2+xQFZt1IU
ZaHo9ai4Q2SLgaiYPwKxWSVilCTingZwWSca21Yl1yI11Xs6F9UXLAhDgCcyEmGrjNbfczbejKrS
gOPACwcqR3raYsor1H3WMYThrhjtt97V4zLYCXlzbOzEp3laJ1mzdLpJdBo0LghgAxN7FbEHBIYH
wKt+wz17YNKG7AOH8HspBZbDvx/AoC/TI/3kmNrDvoedOZjINduyKpvH01Rtpru8PTtsqP6cv7nu
ZdhTVZS5edtSeit4PzzRyuYZyM8JoMsn15rQIsMlC4cjQSsbaanefFhdafbC3NjahFb9WCeJqYtQ
81WGgjVtITGwdF99INUZvjJ79huTvvdRUWd8XsIS7YWr/YoOfRBy9lw4pzaDMiEwcf6a6DGpRCai
0FeWP8eY3B1t+PbPjChcjFCnWDKny4CqxVjebqz/cra22fu0bf554x3YlzMJXugNYQ5b3qxJ17Za
cvvu+G0CuJ1/bhi5brz5CKlVLfb78CZPGI9uNdvw5sJzXA7PH7BmkQwfLD/RBBqGLTU2ITGDbg6N
VQzKvKHtow9Gi4rNeXdsKqQC32eGQZeMsthe1tcx6DuQQvpsTFWHfW0iZW0/3fx+z5Um5w0jIa+U
mTgPn6jIKgG2D/VjU0/xuyjBfkXwvA5pjh/qF3BVviZzg/2/9Oc3TybUYGy3yAbnyOVXQqp5riJe
uVNH9rrEdb2jexnmRa58+k8GsmXpZ36u4ehL35wf/NkxRLegIEg0zW/I9fntVagQEaH/CUxSV/Tt
tVicJn59gsBJPvC/8q66Q9VnQZXV7VdB7BeKK6TPtYJyyUsmHKhqbgESKMzmbpZ+V5RGS56xpBkl
E26kevvAmrTs7+YsspgbvrbVG7ieQ8P3Lvo1sWmthiXzDO/FnEAALkba7lSQcx+V1OXVtgV592ki
IgX7k+xciJVSNjMK4vpbxxRwCojcRBUWnpVo9FJMHrsEfVNjDtLOTJPoch3JNu56DSPhCPbu4iGz
d7dC4pilYQ2GAoFjS5YIPGJFQmagnUhz9sNu+ASrXcC5iP85GwaFfgLMmuKAWAsGy970uMOEMWMQ
BAsrdkgU3HxoEqCvxizhxkpwkvIVxPPp5/pRc6259xeKlVLb7IzX+vvAJnX1YFjop1Yo40zdmZxA
nPV2md0zxJ9wSiY=
`pragma protect end_protected
