// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:55 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
NChvJgKC5RZ4d7l4yAe36BMX7hjZ1UuqPsdwYa7d9ki94VjB4TPDSb+fHmg0A+0d
gcgGuUYIOiIEMlRGO7WwoN/Y0vp5uQnkEo15Ji7lNSSBMiAPZqEjgazE5aokN/92
8e1EYGK3Do5AuVkOmjermA+hHJF4QgK1hWnDJNlE41A=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 3184)
8qNnG5XuGWpY4nbYUqB/hH7OXyBeNbjRrx64/Iae02I4vKKhYf8LM7M+d2bVguH1
F5Dp1w+eZln3/eCaitIL7ylK/9pV2YOnOv16I9rjPx0f7Xbf2t3dbNQVBuuKKmhY
F9bx83hZ+hMvNKdRc9YQGiulKLrXJ0lLraXU1mHPZ3BA6Dqmss9ILyBY0yty2KHo
ZGReweH/JyZLf1h6FYXLg36Js6A5gJCTw+f8jZ3rhCu9VzYmEQzmrsHB9KjizKGt
atGKaIgwUVrUYKEaAUPKZbPDr5iea+qkkfY7uCjIjw3TKb8IKj4JKQ2394cLT9Qe
bcZttcVKX24+LedAqsRiOaRWoIfDe0TtDTJ7wGlMXpZ7zbQZpFqQx9HgMgNfgQU0
tUM6QEmWF43Gdn9Q8F5TdKmr37TSoMeo19elkkPS0eUoCDiUpMLelVRsGSwCTeGx
kZJuARGdZT8Eelyx71AgQy9w8NMPDw3KQeRWlb6BFI+5lDA+naGrnG+lucdO3A/m
L02H04nyT05inwApFeEYwf/l5vUBY1KaE4ZyMHDJT61ljnAW153OGNqyXyPlRH7G
Ypk5mDFC+b97NPs3TckqCbq5xpeb097fmdL3cujneKmrYdnC/fNQHHlzS/oqixgA
1jn71EUQO99buEcg5sNY+T7ty7YGLLLG+z86PcyRtcrDPM8h3URd5EBvv5mckdnX
9g9g+yi5C5gbQ6x5qksqE1WMYhjcb8Bw70fz/XI/F/3uzmADTMlVRD1+o7zTIGSW
ZdLnr/ZNNg+kwk59oOeRWfX0/sUUYECN1pPoVpKbyBs4as3ffS/Oru/dRsfVhsrG
6FgdP2fmrF7FVHPbMcLDN5HIonZtjiSVTobe56MpF1FCvDyyePaLLja8tOjyiCUx
Uj9HwL3s7dE1Ya6sGh+3PgcZR8GMLxigsK+p6+rknb4T9JbOQHm31u/yCWN3TvBb
7oXWsappcYA9/u6R/L5GUsuAZLnD/PXb68GjZpAOMnczJ/J/DVkugAChAvK1euk8
eVTj7vpU8Du5G6+7/fPWxvxjyJqr82UNRILJD8uDiky77tHO39M0hhoW3aX7/PdL
UUFpKQK5VLz0Bw8VNLOftUaVpDaPA03YilSsVFCzJOE8VJn86eiXR/DshDtPQbMH
Tx9ox4L0J8kwMQuLKxzsPHID51Dwfs10TaImG7Hq/j7/xg5sRluZZicaBMaSy2nd
in/oL7TTkkY9oLCzn5VTRWOk3F2Bn1dHu9sO2BgWt9K7HbZwIfSH14Ofgo+lLptV
FeBAp2pkA088LyPCPdk04IEYluPx8f2g/prjGHAtuU9k1BXRxck7xLiDmpWmByK6
0NwAnQuWX6ZG7kdL/K4sFyuN4RU3AnVIzWugD5yWIFpHVp+675QCtaufZepzaOcD
ugmm/BixMxAGz6uk/aWb1OO9A91meMpl3Etjh9vKtSeq+3JWaZXRWXbuA3mfnf9c
zUd4InAlvydqEB1d5qkBLmT4T1fk21DGJrMK5n3ECjxx+e0AFIZ7JY+5CG+bs54h
JRAOylxkCKliSivggD1FnGRr5m4HjR1pkPHFD/N3UPY0dvHhbBo5z/V3vsmWQ8WL
yDYFvq4ZqMn5+arustrLry3yd2dh+H8rRAtRcQPxuq+gbXAUNCWn5mUk18qyfmPH
jN4ZHImoKvp5hqpj1Cd5MYQgp1x88ebb+W1wEZ5+M/LgTwSYLrjbUfU5h0hOZq0c
oNGoWe3W882wllNpuQKszF19ZIFE6A1WhyZ6bqZZHfyd6GANIbZLczxiqcJ4qly+
Sr56+vzakARVI4xLQ36kZ1DHuxVhY/roE5i5JaXuC6s267pCxSfv5YRESswAB9V+
dgUVV03AvHBtNPH3ZxeHU4Txq31t+Luemp5Yoyi+K/u6jsp3aS2B2BQ643uF3Yw7
+HddPxSSuEIz+3NGcf6d99+4A9ELWMPbedsz+Vi/GhJIhSgFFh6Mmf8nD26q1fW0
q87L2zjhwN1R/Z+BkupIzz+MULFb+7Yc8PbglHevmNfFLcz3Ke4jVLhATpPQJpi2
bud2dm97uEPHKa0Tff7Mob3Jxk0KVzfzIkGVPZtCKqe0osbgljXzfNtUZ4kBom3b
RMmpBXG777PC/Ie2QHMsinj8LkpBXXR/+zi0ZOzlAVK6D7f0wShpG1+KQ1rO3LMF
cB30y1zDxjliSSfAkbjJ1pG/fdoo7pi0oFNIqzxuNJDbx/qq+m/7PIerdigE2DJk
TITAM5VL3Pt+sI4tb6vNEeJ1aNYgT+DpnyYxyq2IBu4vH6xHKdwDvlYpRnsP+8Xc
Akk+Gf7ZsnYPmy76EO/nxlmu5qyuRMfnZXKTB9vrpAFzWkaGD12d/TopJRyBonki
ePBbwne4vbTnQJEXCalIPR0YRQmsIKaDZO7+6q8Ne+22UDt6AuFLo3vBVap8hzUh
j3dOR2snOy2BZwIofYtR4ReJzmNFauJYW6P5zg6cjblwXZSHjQdWAkw63e51MDw0
RysnOnpgXWDiN4m2HRfXDjT20S4fzLmMQgoen1MuAdl2h/2PjKPRDh7YT9B36GpI
P8hKz84yAw4u8j0FjLrcaVE+vWv6SgyBZ8uocarf5HnqW8IzdwI+XBq8Enav6aE6
Vki7m0cQoBUaEj9/eAX/lQw654uLyU3CSA22T9HH2PIwYUGnI9W9jHMDKo1M70vm
OzE0eX86+BASZU95DJGXqEMClwOixcLdIlcurptE3esz58YLLE7/5IwQShXvXwl5
emKaElXmXEb6lT0bmtMpFhIFuHN6TQiKQowP6LSeCqwYIs7fY9k4nwwxpzCAZuba
eWCL0jclphUauosRya6oz0Z11C1PsRItmdcS/N7GFXEn9xFx0ALL7s2qIbJn3FTL
t/i1g6Qug/0JtHCF4xQi/pe5eKRTMJrS3dD9GReX+UedTeJePClz0nFmeCM/I6QN
ke4+tdvIVrcXvvYbbkzwbsZ9RP7hzn/2tdCPPLdEHDupYVJiDEsgR5sRRPR4ul3o
sHtYswpM5arRFcZwMksdvHS922fPQ3u40pSShtNamMzCtk7/6+fP6Dwo91xvmXU3
+O7jrkv9h3h6gCeKpFxxhP1Eqm7Szg8IoldX+EyV82OWV8HrzDe39GVNfd0WXPJ4
U2rFMNIDDetxGjegT1Js86l4sfThJqZsjbawwFcP+exfkFNgJ3fe6yTbISiAGbVO
EKvnC6x4qPEC0IWL/Uww2RYy8rjF3Q0mTUKZ6RuDyRP6+/hUZ6jUPwl1RcwtWTK6
5XiWRUeKRvAYhLO6LOMcrju7mm6/rfohz960PyPolaaPmeJfxZqxjjj3n/LeJa1z
ZgY/Hg445JfO8Dhjf3eXsMQ90N20CdIMj4WOTFASeFVqrSHiZ9I1nOUNQmbjgFsf
ToAIdWTt+9XPV674ueEvYOpg3MZUUec2hFUGqv9JoHb5LC0UpYTSUwU+sQz9XTIS
DOQMjTJvuiisYeFfcg87rTYtCZadzBjU+dMiMpdOL/fYtmXs9NXrAXIY+Ttjy5/f
4VpV+/tvU6r5ps7XKCKw3i9UtP7UCtYJtb/Zgs0zHvGM2Vk4bVr+l0r6NMpqy4Ci
sROl0SrTGqGRc7aFM8Wut/zNaWwgMVbAQS9u+HNVeI+se13KyFkwBok4GkEsd2X7
PD4M5rf8zCKWMQR3nVfI+59oRR5J+6DRYprl2OVHr8WeWIXodaDHyCApN7DGm1OD
n+/lJA63I/oLBRNhmx6OmMVq2wH7NiTs+KvyiKYepcbf9Hx919x9DIzCpn5VtQbj
OyNrXjtI0RfW6k2ODOLTQwF2Uc90S0ILefIuNxEtesoLznMT5VAL5PAXk3Hgy3E7
EAR5lf/S2KW0cwXSH7pEzct+rtJbLsOIFx0zDoTp0uK+QU8nkLL719syHyHvk5vR
DkzHgYvCT9wFWlTZUY0Z9dtpD9I0NSgv7OA9P07U/ARk4y+twfGPpNS/AnjxSDD+
zFPYW7QvyY9LsDmcG8VGryboBwAkhius+Nmy9PvPtJl6aC9pABHm6XojBo22tGpG
hmSXj2SoAjXGvY75ZwT1Xb0rH4FKXB0RXSXX6ozGlb9Zj8fc0HMLy52aYNTdTi1B
OnQO/NStMm5s/IyKOjffd5VPUrK41NYtWqGtC2eUm2AOTR+LRmm9GUZ3Z2p3ewsc
yt55Y4zs4PZg5mH2x16JOeJ6SAJozj2Uxr1DhE9kw83DfgzlCJOfHHrccU+d4tlO
gQ8eXZfyC6HBp+/HUmz7uA==
`pragma protect end_protected
