// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
tiu9v5F49O6c3wm0gG6zoQg/DdopX+V7b9Y2hmeBWEOiBmAGCSNXQ0yaRze0UkB/PYeYgYFhoXj7
8vRBjXK6iX2+3S/CGk4aNAXBVJLAXaiMtgYfHZv9ksk/he0w8Umyd6BwiSZiCvZaJkERwojeB3RT
io3e+Q93YIqvsg5y425QmM+kuihQ+fL2lCWRU3cPck4xbru0wB6cQCVpsTEsep/gANE/PfCtVtfP
xkpKqff7MwQkpSXyO4n52vouOd0tgBkYs7yg2lYq2jxIZYogbpSfx4e472R/LwiSfKPg9gO/2lLC
ucfD91nGI4Hc8ImFv/z1Ee69bT+/zMx2CMAq7g==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
5qe80C5vWiMi3Q6UeTmtT4cbh6Qc85wjdmW7FQ55VZYsYmGpFXRJQvjmE7/g64ZxbYvPVZL6RB9l
KkwhAVXII44ZYeSAJfaPToF7U+Kuo0I1EKg+LkD/URW/Vxivjz8E/PSD7acbZo7pv7bAwLohQ7rc
4GDhW0CUXwCoX9/ng7MRrfuED6f5eJd3SdvqdvhOUOSu9/ExwLDNbcvO0DBPco6sw42FEzuVPNfr
5n82FzIhxFj4axqkWU+e42EIkubMStSCigPXUy8QUKR8S/l6fZcv53+lDsURaQPTO+zCXkJTR+Gs
53S1noWgANqdDAPLr2r687Lnq6Az87YFGZq1+iq5D6jSt5fcY68qAnnn2VnytqqOFVHCPDxxeGbH
WdzBPX7gpiV3BcT1rAQfOetlijqD7Ls8tThF0XJ6vRZmsN6cp6Zy1lr/cl1rfWtS8lqMfGvX9lMi
DNad7cZ2Ed/wsXp7/eXJKQl0ioXYM1Z176PWAatffd/5QP3OcwcqGhvH1L3OtdlwL3zcRSGe8jLr
RTpg5fD5VYsvNU0NdCoEiCE0YX1br8moF0zO5dFWmVVp0DJljdwqAjLOBN+zx2tfB2g99Q4IlMlD
CaUj5FgwfU+TsDq/DvJ8J4UD5N6p3YV3U4J1OxOm0TiIY+TpQ+DIAVcKQZ1Q5+R09DgcjLnSt+Sk
locqzHOLux+1Uow6/U8c9lZH9A6bnIDFXUM7jDeYwFtEyvx5bf/hY1raZrrtCNrrHupte1YKygSU
UJZG1IyaiXaw5RqLpkDbN+HIVVeHP2dcbP4jzAsEgT15HGGi5FRoDR5QsKHFjxXxMb3o3evbV/Ni
jiOsjF+aqE1FnO6OgSd3x+GGwrQgF1OltGFdzTC3TzYa0snusLnKcV3KfuSHSGu03jmTyrHpv7Un
qWQsiuCdbeUJKPMAokfSAQS02B/rITtzlisVRKg3ru+yNQHOyX5y8vz02Qt9ricgxL7HYhE7cktL
pK1WUOiKbR4tG+sEDmjUTN+gRLQvZkyyEfID7qF1biYlZdkik8khLUWfjkwDnneXnenzSPyxguKY
yOFKN2Hk7D1G1GIhBy0j7QJBAfwyXTz1Ma1bUlOrhTULv0ZPlT9CkDFvmLwLFcWM6ajThGv/lXej
Cah50Jb6sorjMgmNppn1iuwUhA+juz/AEwh5lXbAKyVKgEkMFtJMn1K9m3e8KEXBTW2hmiYVQLwR
qOVsIEbGsJIGoeOb7yDyKHIoErwIPOlZ2640F5gLiYsHO+Wr+LOXNPt5vvhY+M9oQm4UL6eopsR0
YS+T5AhZKlhqFPouIQHdj/Ntk0BdW+FGEv95sUTrjGfND65BH0LA/mNFEJs036gUsNdd1xHIaTuL
tysM9Of3HeUpqSsOkYXBfliMxuYfjRrhdMDxvfqkErZZU4wqf3QjKGumaO8oAoqmKRcbOsNbnQ2h
NLj2d7w+Vr7uMciU6zbg0e0u/4xQb/bHJbEioU6RCAC3UfzeuVH1P4dvogo5z/fKIHiH4vqMXkEw
KtK8gwLSwQHA7h1NyynT7PkKJrGEDbxuFqJdWvMWSTh1uCutYwIbJixVjJPvpSV1KAEUj3/DbUXw
xKKpubdn0rF0hLZoueQzQen2mEsXjFZxmxnWNvqQ3g7PK9CAPfBmQRhstVLSkEmb6l8r4T3B6rrV
LBAzA0B27RjhnTx0Lmn+BKMxpaPG5ffesXQ6x8oDWUaLCZJaJe5YaHVEPzCzGB1Uqj1vLyJfq7oG
d0I/WmOsa2f8D+kFLEgoVXy6P2Ea0+5eLF3ocez3OqoLAa1l/nJ00EuyY0055oroe7aUUkw77GfG
vBYdNULs7l056h2x8PXbarvMwwoYb1JBAX2JPL8LJsNU/TeWa4BNtZMRdQ7WPCHSxgZK1liZ9KZz
UL9lE/j33LOBW2TxlkjZkE2Ab58a3gAIEGuqiYaxdYbz9GFQcLRcVemUfvaccaBm03XMxeXogdox
eKtmoF9tX30ymUxAmFfJbVLuOeO4fZV6Sb2RCYOoslOHDAIeW0jckjAKnqXQtb8Z57xh68QrTVsz
0Q+vCrBKVuoJBEMPcGADVmUa3TmT48KTmni9ADsDplfLm02092CcfTe7iZyYQyQDYaBR5WzZ3JNf
jvebo9OTqRRo8eTGCBNE7ryt2ugtewKqyCV1eYtTuSxsWxYFJRjXvp/bEaIdhqS9rrJpvbvPjWfc
2Xuahx6B2ZdRH0KbcjIeurNKmyzaID42Im8LSNQqr/HIJieoOLs+bIh1OtVq8TwwIe6Mqkd+Db7/
PZ2L6OKFpvZ5roAMTIrWCBQFlfH25qpkD0lHrfR1N1JWyDIfZWXOm2T/WPjbkM6yI0EvhVY5ThEu
om9De42jrb/jGQr078r2ilc+Ylwpe6N2D+zVjvgK9CQ2qFBUg2NbiMof08pZHc493Td4tLviEIBq
EV2Bl/VPJ+b8t56FNMtEpw8LnCxyKWpRG0R1ejKXuOe209waytevgcvWK1dH4ZWrvk73SQ08vvae
Iz7R9GgomFueczYWZrO1cbyiIR38umXEyBskeMBU6U8O3lK9CE5mxeC8qZ4f9TdBHQ32rgj+G93x
kq583se87SSavIlnR+ZFHRnjTQwDA0JCFvGGY8Kf+HRHdiwVVr0Z3N0erqEGKpGgydUDrHwjnuIu
3l7ddmcmFOMaEFx3TuK2atYmoFfjLkH/nVtna4Vx/Fqq0mWWyWCFmXUZna5polTxpAImmxHZi00M
69s73/ZaUncllOwf8LEhqB7GsR9yU9VYzMFNGePWOhuNvTh8A/pU3djzTzqUVNsaKizRyYHNWsa5
gXisLbZslJb/QHMT7lwzhcH+uMSqLoeo42H5TQBlMGPQ+f9ilbYI24kBFzumGMHrACZ1L/AELkoJ
2hoG9VtBBbTrFtl1mECffnTqKV24wDl2b5Emvyfyrnbffy2CwPh/UR5avIK9xgQG5FV6EwKy/rxJ
T5ckPH2PIULWAG2H9pJcDe1XTXDY9zuGP/kQ6lW2YExVzDc2gD3YN1QN+3Sxap8GfNLGw8JUeEZX
2Hap61LYtFA3Qae18EweVpSQNk+2/TmrStSHmnKhRxTgV1Bu1XLi1O8ik3cjmU9SXqN2TfHVy3vI
nc/kK29YuTV/lgtmPa+C1pURsrIENdHUtZ/8TvTQDm8VmKjS7oG58QsF03xAW6Doqg4JghNP5Mhf
CzPMvEDQRsDMlhzZ/qsoJGF1w9TOHBmGbpgNltL0Jx6a4yK3Z2drf4EgLWbdqCoga4vpdGHgJ90n
XIOkI1maFR3bJGTcLwUyXjHK67GNko7jqiWz+drfPfUkgru12f1Q7dRa55IZVmFc04ZPkm6sU+zq
TEHKaP8lNW5YIPFMPJrzk4g3nh3s6BHmmyOR6JJaFRQ+PtqXUK6vb+uAVwdMGC7EPPKSw918QZl/
vi7AurM/7WOSgOLE5YaHIN2+9PjxKGxe8PVQ9166Wh4pF6EXyN9La8LLjCSOOGA+PZoJ1Q2IogbD
UmFRKgmebrqi9DcwkId+GWCiz3cqIxujzT9aWlJzbrSQbMmV8ggxxLk1dDmqaiokq3zzfJ1EiF0a
X/aoYJH1/oQ28NIsCQnMSAzK4Fkli4jd075fhf45kb/f21DpiGRy/ovShUaqZy04UWUFPvbMY8si
C99Z9Sl0eaecgkP4XOeJpXsOd003kky1vVtVRoDHS0KPw4VVjeoKTFXtn8ibdefiyccVzGFOdPYe
Tf0nqvAOmjfK7x8qxg12TSMT6SnghRoS1pJgthLg1ouo4eIHGlBf5meWCZ8viwDz0rtKN81rINDa
5XzMRUgq31jTtzHsFI+GGBv7hlTivrSDeOvG+p+Njxyldu8HV/qZuIQ89kKGZpa5B2wMHI2EU6ep
wWA3/g+pnCIgyDsO9P95M6b8ZAtK6bzUWsbIqE4HWxQrhNXej9QWQy73LlnJv0UgyIR3PyhRpdsO
Ot4/8FcNBvHH8NcRaz/Hr9RGfkWk9OHRQLAAkp/Y2hTtQtY7b6e+wgnH722fGEfY7q4bV4JDCRpg
JefNnkUpD6mdXUBwzfajmrT3FLIH/HsUGHZDAO+XN7rCD9Fk3VeRX4jKtkJT+wXA+Wg2UJgIP8zl
x8YQ/KUAbizAH+KBjUyc4iqTDdHtwL5sjQDcEryGGL/uRYrDZvxDLIXXIo9HUkebJ1YxkOEv6vxo
/GejVQsNZeQRAx6tqvkqtE6aLlhqPvomPHt0d3gC0m0kn9pIrFA/aSHnbNszVDyZj0yZQWWLsCFG
L6kdPqK/tL9/HLJLpL9wxpPDMsAUtVKOihS9jX03FKDWT1bTUrz/2j6en4fpDPmXXIFm8k2urHVE
2lnA7fvR/iY7kY1XNtHqGoVBqm5+0uv6J2fyDZJEe3dJ9g8o8u+UtjfBAmjksHN4UI37Z+rmKznE
vhcAMrP+ehJSYB4YSnwzCEf2xkn2q+iE5Q4rIYenOf+fJB/IzmJOX91YXdFK7NHCJ/skydAZpNne
bC5bfkunx4DRBQJMZzMFn68UNZRNVNn1tEOHHVf3PL503f0fzCDpGRKoPGqbjCVd/nJO6h++Nc9X
BEVhfMAMoJTlNJPZcopXNRVtr25/yS/fbbVX63UzSOZWBuP3LOUTFrTcXuZ1LH7rEVqVGA24BHHh
8rxJrtiu/dfMkQF7VIoTc9FhanIJA4WGTM5FC4ciuomTYqAFNtRZLk90kUMeu5TNMD8L74elT6n8
YZghb2sXPh8cySt5lbrTFtUeuxf62L30gk7WpC4BKA0kDpfHNOEFVcuXFqo17LjLzqYJSdbpbalx
phkoD5dnEP5Ol+c6F0muuOZo3iKq/W+uvcyxGXyycmimjORXJquvsJsHWvS/WDKXoRK9yC68pJYv
pFycdRHr5iPeK8z/+mxJHXDbp9IPCt2NuHc4KApXuM46T/lWFjCYklxTypIbUQ0PI5EIW1FPVr2e
g945dkx1aiRQuh7mXORihAd830/oC0O15RcUYrJLEEqkxzwrisvfXA61hzP1h5YrqfoTbp03zsq3
zgpZuH5UHObNeXLm1tfJ5++32wGeMSGYdmOVErme0xUb4dgrtCwpQBeO6VzgkY0ARkVNsuW0CiBz
FvBxTFwGUVhY5xpYr+xJbGNLYdTMTco3ET1WmFEnApRRA8tYBaJpuy8l3S0W6MDXP7JYoW9SnIA5
aVwaCgy0v2BFw6l0SIXEu3iT6nrMEJdXawFXnLXrsXWc3NpTmKDS6GzFqlJRhpyqWmuXH4ywG7BG
6YO6A3WiUhKLih/Lqv5iqhPQTdbNn32UbXZPYYwN6veMqfANzDiqElZPXFq4vkKolMYKsU56z8mH
SZthiORIXRLPpLBsbEt2T0Jz9XPr4N2H/qAirSOpt6hNYOsjns997pOX0KQG+8xKm9iuateKv8n5
CSqWDfqWaPq8W6G/Y7UTIbHYaUNrL0V2gD3Nw8L3cBCseJnRXpA4jSyr0+1f9WtTGVCYnoBlzqOH
LnlYiXt8kCUmtGVe+CzJgGOfJeGfTbiVc1CWEuJm2z6HAQPRM5xFLfcJQkNTgxJbgqfIFHC5GZWo
XaqLCX1gnX6AOjInfC7RS/Hyy5VEnPzoamQTUTSgfgaFY7+itfk8nTtH/eUmVFN1TFfxHNVpTF00
3Qc1uhutwKyxk5SfuUiFKHb/wRXtZ4n9ORU9eKTwN17zAGBDLwhMRdaSVFGlPS5zB6JyLJKwhZDV
5/DCFNvgiUDiJfy0r3PIkXT5Z1L0c8sZ/mj8/xY4t0LJGpswoLGbl1EP7GIH0s0TAOErtotTF1CT
vKWYw7q/MPkidxjQf4U/zO80/zrZ/40p0gLmqtyG8DYnJE+rgLz5v1oDuMyaH1i/LdcEQoQC6Vs1
GP63zwokkasHVyMVeoc6EWyUzHmpu88TVlcheehHqD/qwPSj7/BtgJZXRbzxnIoIKbh3eYNzEbIr
UDHD2iJiXThMULXeH7heVcI850wPzqVgHYrr3KNhazeCBBXyOrC1jsGyBXijbnuqtsUpK1T/FPsJ
BBjDYRvPwBXWgp2ohg5PncFkIOHOb9Q6wsqQN3dtbqc2ap5wHdMIa7O2GbW2ucaE4wvA1pSWgraM
NgfGrogxv7g4E8ca2z+FnB9qsbp+D38NAZjdAA9DBBhChFO3fQRJNmKAvhidKC0M3rvmBPPNGg/s
WvE6oPF991mt0ItO6AyWtyXjfsjiT8niV9ciVfT6UAiiC9vz59pjy29yo87MpHH4ouQ9OLK1lSt0
apI0AtZFRqmvgapoN+yx4FcgKVbElS+yLJHOVskIAvy/DJs6jQa3J9CO+sDTKp5ihJf2P74Zqh/c
SZS3m9HKyyEnOtYMmYc6p0sq4WHSzojywWqGLmCWCOeertlsFoME7BwqkqS5R1EvMLFAxU/lDxSz
YwgvoNfhzYFNwHfCqDu3Tdulh0kNWum15X0Hp6AU80hJF7P5VWdrEB3bSAp+8GAWpmV/7GujO+rF
hzZpe6YURi3dTf4Vc+TbE4DHFTqHzK2vdD0qys0d9DSLqBPpo50YZL1+LGerF+3mnIEfqqM5t6wq
A2GyAuoPHrLs30vyh64Z2xcg31ci9x1/Eec7vQozAN4/TInCqhb5Fm6+m+5bdIGiVvAE/oVLADp2
8AS+tZ/XSBwlGH8wVdIkZzUXSbk8Hsfn/D9pB3yD3/9UA1VG0ZNTrSOw/PlTvFmq+aBn3FrR0OIl
ozv6n97DgQw/NnvGqKmExolhni370mCApCF3B3Dz0SbctMNBhkM1pQBmHImOcwEa8uzcqrSYcPNr
HCIiU3XIZqdo6RsPCKHQHInHpILbqPS0TZVIlCkkfcPQXOXmtANS6IZb19FQKRi+Wrlxe2mMGBh2
9gTGlotBDO4HqUTw4e/vf3IAnqSHFeAsPqls1UbysmnQl1NnVb78B3jZ5axxebddyW9nTpquLIOx
1P2rGE0GtS8mk31yW0fBOcNwjQcxewBtdsfZz+LyFf89409+DTfGYFTAQOASPh1rNQhwBogaFC75
XCXAxq4zoga92HdKJ9K72EgSOgsXYpZzjSqKEGu8FAFVU55G9dWnXWC+5xOenvoucxctSrA7skE4
z0oLIznrSBD8S+WodpYuF0WB/xHrE4SwSlogkxyFk0wss+nzp8agA5tAKrZuYs9W03CxiRqF27mv
7TBwLDLaUOjWf6mSfDsIdvHTumnibFHqQGcDcwU53bI24o577ud/Bc6AT56oKQzW2lRne6KdagZd
DpimPPzNSm5gln5VD9rXfJh8pIcXJdWZXlqowK5H1Ctqyh2pvbloqIPErsI64MDZL8AEutXFLzzU
YltW1RZkKhDFlN9NILzs/MO2nGAqXH66cDpkFqn4JtVXypZcHfHv6A4Ivt+05oryx6LUw+n/julG
ssIE8ZRZo1fXtGG5w3W0rzNX7uhezL6Zj5PP6FoCwsrGQW3rk18h77n61M1CxdySXgc53lc5wO9T
WY0a5/v54g3THQ21T6skaHXqxDNGm0wFaW81Jgjm3L9uHLIQvIJWLErmh/0UH0Ozc7QmUG+kz8EP
kdOnhqjsEXlW3Z718amXvCPUGt9TbPXnZm1b+wWyqGgDzPTj1avvdZdOZnX2ZI20WzxdDwP/h/Z4
DOByf2SDjPm/IYLzPvuiMip9Kzn8ImKQQOABZNBoEC01n3wi0zZrEb4VQg/blc9Il7Vf1LgMBouL
QoSrloZ6CHDbL4s5R2S0ZSo+7mNsh71DxuuBEML8mZO+vtKMs4Agk5yJFTzSd6REkChAep+oiV8c
Ls3EoPdeBvWRQsq7caJYBmizOJn3/biDNAGcZPOT4zeDNcA5rg7lgBq3x54Gbp5Bc4ZUjcEeU1kF
hkv4Ctus8mY2YXqYyY0WOEraUEONLm6fGC8u7Fr60fLPByb9jklrNnTFtgqFvPA3a7B0Pqq/1toh
VZ7Z9n5+5p5ra2hJnaBmXBXb6aiQRouQydR4xPl9FTKHpgHDFwj+bx6olUDTwC7R6GwMHoLA0jX9
Dy0evBgXHLzji0MZDbTTk68xZQt+ey6+to/OgoolmiwGbZ6cReO+sGss+R3j+bIbAfy+tjs2+9fL
rDocLi/O/Zl6FIOe/ssXB26zdz/IWGC5CTAXmi4fAg8ku3PhjFY/YIn+Wm/UmfZ104oHjRVHuaYa
xyZBuVutTI+0cK6C9SWeEUw29jT5mTfVVuE26X8bMtb5ShinGriVGlI+5M42GgSYCCCdh8PlklgZ
Y6D4vudRkqtEcRNjPEtabfzuRlIMes4cb6WRxhg3U8p6c2MLMCJi4VuxGDxFehEgOOEXTPCl/owb
mqu4iyaDgTObQCJzIxeg7SfkmaTYBunhmyCh9aA5Pvpgwgt/wUQTUZdm6NOILZZPFQKh/RA4FA5a
1UPEtSyRULsclIKoVLGVtSQAY6pCZJTuygJFNtT99zGu2XXkvtacDZJgApFLF36OA9Fshz0crFTZ
WtplTYnJRNTuv3pxRYD499XixPNT3lUDxu2QtwlBcWhbetJg3cIbTLTrbB4pBkWY9F0MCuIYMcY2
9oEOo9rlWAKh3DsqY4qUwHdoVQt24ppYOPeastd58OF4ORzoXYh2niZiy0I9hxDRvqnmHJ2Z0aVC
d/8VyVTgEXBJL8Hqbb/Pzf0rH2XE+oMpQCpQI6EjgL6f/DZ5taQWxVtUIXKeS8sULszdLQM7nG1y
P7Cy5mtPrHiPnynC5iATDffZZyO5qIAQVHp/ATIF1p7/ALu7poNwBj+JZWFqJDadqWuAnjlTiCJS
rlu9ELp8Vt7ovUT1kkvxVR4JVdLMRmjsXila7WbpMYzguAcdjmJGndCRKCQLyeeVfcHnUAA5WNak
zHkZZROW+L/x8qOzy7igPI4Q/eWGn4kKAHxkacNZfsgh+ypj/OndhpnZ8z7yTDs1u6rlI4F8fv0i
YWmsJrwSzGXXbk3dsGuaRe1UE+O0KvjOubaUyWjN1m+tcbVhkNljImL86DXJMlfmxL9fVJ+HkjTG
SjFeQO/NFGJob8rTjsUe3exzE46PMq2J1qSlMH/g/N7DQWR51MBlENsVjOwhE5+6MuYdvZ9X9iaa
Of+D+QiE1+mCL2bL3OjLXTe6gxTia0m5GJRa6luMKzirIPYIkuIIoYAKxohk4gjOUVTntp5JXUlB
9brpJ3vRZxpvPorF2eH+/eVJUzTJE840MeYGGy+V7qUwO3GECT+CmapWDW8Y9jt4EeHdLxObJOeu
iv/OdV5QR3m7bAyMLY+JC/Ptsgfgcxes1uQqiPnwxdT4p4j+eL5VJlSOP0kBBnDSNuw3Dz6HMdkZ
077Mu2wzVgYeCli5Vo9cDgInqT3jEbwyEzGvJWcVaBqhgkHHV4VbAQ1vaFVaH8BQzAVraTQ0w+dG
ACjvuUieT5Wz0mNSQ8Ll4l5PRt/NN1JkD55f2CDwrR8bfSJ4oQdLgxXfVdUJU/Tlc8Va1dTqzhMF
19fXbD5MIkGLPODb7Ghf5+URvcw0THAB2w+Z9He5fCZl4xTwcAHC/eIinNzuOiYSphwhe0D/QuvV
ThuXdoHXpRV4+u6ja0N++Cvpz+fcvNue6CNo5W/Who3y5V5Fc0tx9pqs1H0VXrtD+DILli7Ckzkd
66SPENFqymmPKQEZTM7DBfffaQLpUx+NI7Gmtl1IgYzjafjpfIUsz3BcSz7QvVgTY+wZAt/GPOpF
5epi/gwI8ZiAOnmhDtlGWRNe+zxR6dTYQEt+hOSx2EQQEyescc+padptxcZkqR4qvWZxd2pQHbap
SrijLTa/WxRaqlHP4dbmW/iJFQv1NwbZiMUmOuZtBV1Qhpl8qPiV0UO86gO4LSaA1w1ifXcMElis
VtShY8C2KOmn5XGsQbnEewsUp5iU1RJ/+99SXCwmPvBgvxpZA6lcZqSnivn+/EDeCwzh7e589vIj
EUgfJBCW6SDk6bCSoeyog2O+onOviMYyNhCtT9J/zf54S3oibBhHY9lJ7dfHDpUCpH45HkFHL6l8
G42/yOV9Xx9ZiLQmcLUi9fHKDLycJaHdYCAro0ffN6+0pC2a48NdMj6GW62GkIEm9nPvG8KsiTal
FpHT4nCSm02Xpme7xRUouEP8gLgH2h3Fm6v0kf122S1QZeOZKXR4IiLzIY3DmgPzeWqmfLz9Bh+s
8BsLzlUfmGHuR84mMm1K1lm6zsBiwoERja2EBtIJckE5Tgt2hxEMTUXoIEbe1J/gMf5gD2CghSd9
hAr+1+rSgCHdqassJrRMhPskD4cFGUa+nLgKthwZSCZhEck+0G28TROQyabQ0LcurQzsnELIImIg
s4CXmOZle/ZdBexAHdO2lP7rdsSvxmRgG4Nryq1Ow3RWg43iy1MTnyfNo1Uf1vZUex8OW8IQ1Tb+
0G5zagVeMAn00zv+lvtPQqnG4YCOEDrSe32d+5Pm3uCwoI1oFT+7e2o/0b1xez2XmzBN+DuxrGnr
4RjLQHJ4k7YUtckJdyXL1dIp2cl4blD8iQmvM7Itf2fowH3Yl1Mzhw59UkqoSLusj7OPgsK/k+1e
kMsPtnG4FKf/YnRr9/xQ7wj02A9V5tFIGEOwQ/9t35wC14zrgUaUqM84yIMWj72BolU8/BQkJLZ5
onz5ppJQ+NUsC7/3GNbQuUUTHG3Z6d797buGfddxhkeZv5BLqWlxr6d+CnP4Dq70/SnhMnyZ9ULs
wvbMdnbvimR0lTK/Iz2Yv2gXksK7FJlkGX7cyVh5mVD78wrUitnRcYhJNhwYNpD+/5mIfFTY74MG
MrnZae2iCFEU/9pNPfE846ljiTxFGcLUWqyMT9IfHcQbg57ntMIaf42V/BH6PTOAkf1WJkDZfqFn
vekEE6Y0W9x/yR35kPrWclssQd1TJvGSOxqiSScdVkw09HsL61enhtitqVGIFmmsWujcVXay4Isz
ddA+7Iyhyvc66k/9gszszPkZS3b2chnlq995dv5+2krX43PNHbfODsY+76wWYx/vLIE/VmZYsUQY
V35Ob1rVG+vtZxB3BEdp3814a/ED69gggJg/2ZNZ3IRFMz38jWhHUsaKU4+jlyldUpmtNyqa1IOT
rhXTTDLxn/GxWdR1vcNS8u1YQzFX00ZWH0NzuOCLSPn6DJTmcMoz8ZXDJn9JggJiokz7Vhsd5c/7
HVlZ+Mhvh/zUJykby1z3OUx/o6nBb5KfaGs4lWyS3VTx5XMyqeRbXlmVJtlNfg+kD42S9VnJ7yc0
6VCV/rBRA8YCZsqKn4DMuugB2Zl5QbPWWQrtIOpEUBS20fFXRXPvVPzB1foj4Ltvbk48m9z9XjdO
YBK1Ts711zwlCLITJ2GKcFzzExvUnAoN5LfOAl0hewmcXQy4ZAXs4W2E7PNSPpqRPWY6TOG8k6Pl
uvsnj/oaG72nioY2/dVy6zDcAKnFP+ENOllrW1xAaAw3waU1owaiEB7qBGhhDj2eiP6RRJOjp9LR
2ciqUQGfvTbogqmDaoWawRGhEUwTER9tFmJ1oPJ0f8ZMgH9ubTToWR3PVzvwIJDUkHxGokgCEHLD
CgCrHvvKrelJNSbK9nvof/w1pob+E1sThhc7GDAdhhTYmdRWTUFD1dUVACTsTYPgFmHEvGj5bwyE
DO4JWXGgumniuCrHytW6epeSalz8Fq4W0EPLlPQsrD5TGGXlUmnKWersqAKMLPkuw58Sj42SG28K
sGxOE135D6RHx37z66WS92Qj3jP/8drDdW2r80x3GVFp4FCXHbLkUM8rPDtMTY/7wyPTYbjgkNb5
jP/moRCEjzJMgVnPbkFGMhp47EKTC43Q2zcWvRWirYyXtHHLZR/hsQiFnRVDkjByTJb4IaL5ciMP
NlElAb+Dla8IB6LNlPvd9cr9qew2dBsvw7Tn36gMgJiqz+B9cCv6aDkbJ8MANxAxyeqGSzk6fwtP
3J6oH/3GYmWH20NtSauV9th34iDguQzSw1Kfqrwohk5N4qek4qfIwIaMkWubTJilQfcE+lUYEiXs
LR8+i6RKzvXTFOcBWi37QyuE0mFOiMLBmyomCWu7rEArvyHM46BwMdyQT8zaZ2RXsSnFfAdNRend
tOPa4KgZ16a0u4tIEXq9UYX1zdLhRXtGWwkqaly1A/bGLSstFV2SXnXkkkFEuiZ522sBx9Tq4XUu
wUpIkUNDB0uRke4CgzR/ypwlU8zLT8EcjEo+DlqrQz2b8nqcw7jT5TfDeudt5fco4h5Inqjpbtlv
5DzgtKdmK53RVJce0VKvgLPfU2/gW+UdsVykJGV761enSfzfK2tlGLyOViRiWp4+QeED5RM6vHBG
2HuSrNIrQ7bK8fDlJO9VpWY4+tg+0K3xUkQi6y/u6tLooCA4DnEk+UpqYZHWzsBUNx+3wzbedKn2
U4slgDUjZ8YLr/KdFg3rjLicXJ9tiVdw6XMHGM1kxZrGNBNEJ6F12HbuC+CcaN/QPQHeT3f7Wwy6
g+4dDq95riojrxrwhUxEUeAHDQg6KufxJ0QVFLbTAsUsyv7Jh3eHs45QmUyYsN5+ba2Yr/pckmI7
2weBrX5GQ8TBYVOgtvtZcb9Xh+sZdi9hwgczBVIfvPM+TRmIvZuZQeI5y6vwb6esgz4WXDkvx3bK
+JdmlaZ5AVFFR+FofxcqP2Fl6qXOfOrzb40BGroLkMQmRdo9cVZAq6syR0erF+Rh6wrD/SqXbb9s
AspgwL7LT80uV4BlEA9d3aDm6k3yiTfGCBjy0EXlmcgS82vGUgJZRDDgaavO7l/HE8YD/X65fvvc
irD5synRazMbGKODCuuDM7OElBbJ2zJ88klLvNaus2IRb2iKG67zJIgzVsoGJfUs5fYeDPAjob1T
wNRdhEWj5X9Y1tEd/oQuMHgtL3nknnw4Db4afQ7kCkYVZQnhhJBODSYG14tz7KeEOu2xI4AEDpWR
6869DZAVlA66u17HA5JnGBvt9ABZ++QjAIdFdL35o8mwyY8XL5/U+Qq4AR5xgVMYIYLYlCPkv2Ng
Bp35R2Gx3PVsvV/idEznyrTSXAzhL1mkRIdSEJmy6YdQpadXThrGcJ2d/e4iefRdt8XT6ZXuhugJ
GVp2U/Ur6vyY2o+izLpnjgEaGwLX7vpqLek/IfKLHDZtaX49J8/PDpkhhnLIcpFFAqgMQOFnQrSF
oOPJ+vQFWbZBD0pG8kM0QaXBU43/L4e9lca+AS1QRdmuMjQocp6W28U8JEZz7s4IG79B2KDS1R5E
0GKBBGyYFUnbRODYhqpKJb8aMSyOqMx+sACXd8ZHNGfcAeIUeYZRvA3bblvkCUYyWMeDnzzCcyiA
CJy3GRI7expwJ1lwb1ulSyLp7aQlM+7mqC80T9GFx3zeis+zBp0KsfuUk98N5HpJXdsNiE9rv5NQ
bgNi/LjbTArSn3J6TRAukf+d2nDCnWcDzKH/1zOcVL9BTt8V5XoldgktzOq/n4E+BYoyukM4O2/H
tSrllkOl9O28PZ1i4hYXKbQoijP8GAdVldoaM7mhuuGY/cT+GkHH4pO+NPw3DyLxpXa5JqGcg1uk
UrsuWT1taZgLndmfuVERqGSBtqUAexukGJaamTyUD0HbPqXIuJgSwCFCIIfPR7DZtZolquMUJ7vD
jO1X/yIDy4GSukr4psimAI9KK00vLvfmsqRKEY1syl9xfEn6CUuqZ7Sr/UPbLem/xDO84U7/Ligl
w+1AAyPEp+caZezYFyLXYeqv3xyqyEAzpLVpvrPrD6wrRNyB3s55BERjJhnWP7e111L9rZ/CcotN
l/WaNvLTMVDaU6TZaWdPuPeIgEELY3JkLJ96XrAWRK5V8bIRn3gU5Cl++3pOgGxGO5ahOpJZAPXg
gkaWiYxGLNS1sNA7LO0EeIbIudvg5smtLaAgvvItv+vHs26J7vDERE4JDZXiR5AoW0IScHlAexzd
4tjEAANPyzAr7zGt48wnwp8LFKZGyzAwV2W7UqAEMRClWuREF5jzyi69Jo72APqIQzxbaJg6ZEOT
G8M+Kuqp1+UW6MckSQr/5OlwaLdLBqAluYbAb7xg0gOwEJMT1QK2Jna0PIK+oN37m8AozidBEB3c
D6mybM6oqUAEohnGTzKRwe6zr9g3ky/Q6HdMw1ch/t2GZCl89wlHZjiQBW5MlHLvaxQYZr5bU4zh
BJBUH4zIUECRhKjE71bwP0Fe5LtyFDjSt4eQRng4RMnURDQWVGGjLAffeQdtnJidLgA1dXFN6VDc
kDWiqjzWYUxOTfDahszBCijNd7eYMwvJcpTySw1CuqLS5gRnCqKVwKcdnugPJ2sihkSl6tuHlV4s
X8iYhR5k60EGty5XW/BKuor5ce6jQh3P+9N2N1niR+MB0Gm1+8IT9K9BkdAqRoV8JqZoLb2a5Rey
pIkXHSUo1gK8OhMX3pnm7mkk7wEU1JxX2cNRr3+DgVycuzD47Low7i46bmvlSK08bjApY4STEhqO
rkWy0e2X+hjOK9mPb4ZfL1DNYZ/oqYwDCBKnuQ5/htsTv4ndjqQ4pH4xRaFw39eI3a1ROvZ8MUcc
Z7U2n/hZXZoFn8nNbWpMO0mGhfoKPhmf0ifr4arNmFP9DSm/P0nFs5xFQsXC9OyXaqcRLv2Jl5Tn
HHAheGMErNJbk0oehp3xMdflQw/L7FJfxy+z8JK6vBv24FcUJuuOLEhlTdJ4p7aiJlKsi/8/KQFF
DmFvNLYz0+9mHE8VrpGFHUEZN8RL5+UcRL38pB9xtkylnX0rlNrBSRY/JQkPFXXx7mRNmkliqoZb
exGRr1pnZcW2UNJMNmBtr1fnwm7nkGxFdrdfHp/xpqMRZApFnKDgQN6jNDvT0GPN/0ddCVERWj8b
EqnuFdD7AZw4JmiMgBAn2eqgqcbmsgmWzWJqfpOCQlRJ3gfeClWV0iyuAxFLr4w9tY5yOow3cWKz
56ihCR0uaaHxLDK14Qa+WdyeBZ+tpmzMR+OgK7soX9JDlh7E8Gm34fq70u3orU8pYEKedqzoa+8Z
csD5PPrcyFQKYvjBovygPfYwhxWPqw5Ebp+LONqW6jTdymDDe/XUEwTN9nhXlwW0INUqtlapSUS6
eDxy83QQCUKgaox4g5cHodHWD5KY5oen9LFN2A686LRU6U7E+F0AGP/6F19EyY6VRCEKI0RzDOhq
8nELbnBNAi8lI7Sd6V+TMx6FX1D+z0Va0TcEEg8PnH5D3NWn848jJGByubY4XJrdE6fNW+odeJ7f
IuY+4n8B1i5/bohEzKe/jkpW7QXYkU5HxCdyyPSzDF/ZRBeTuP6iINT8e6WX3uAf1C5Xb3mJL2EC
tYKvxCZq2VjHvvK3WASUflTlYQOpG8nEbHtxw9m5AHz41YLiEXsVNeb2WDe2s+bGfS50VZOLEgBt
9/qunaHSKUEU9hGmnz56Jym4YjFbuzHrxD/ga8gFLPlpgMsdsOLxwtLLaBcEHwTVLvQz3KVURbTF
0SauYBgFPdgRs46BvBmp7j14B8GknkF0POLcTDgWd3/Kcs7o5YCoiUb0a6soCC4so001HXyGhKpf
wtC1DM2SKE5zbH1cKr8GqE7QtAwTLM+tXYkFMbJoAgcxo2iv6crChvSYuOAgZ7ikgl6QcFtnIr6U
s+k+b9W02IE1FphbL3a+82YlUC/+jbRJxKd9OB+0F36mM/2RaVw8DT/uKDKcKkzmFqgZSg5d2Awg
phxHSyspu1+gFhaZO5XIqWtoQRR8MxSFFT94yRcyQitHoa7kh7nc3WGdtLpcizqWuZ9O6zgr7NZC
wAJWAqImg2k8G2YQky76Tp4bZg0yzlv6aBsMPU6/2r2jDcCCu4VT6eOrcZYaZhq6Wn+xPDveQukv
xjYwYM/9PUm5KzgVXlKGX5Asdy5K9NPrjsvxf/0RCTdYMVcFT+tQtgSvp9bQJ7c9rZ/j432K0V9t
gOW8iJfth48QN8t+vGi016E7X7znG9CYGyabV2yipNmYZtqF7O5b3eV7iz5zZ0vuNsSZYgGONUH2
L0huatuc2wPGlULEi7HyHo8fcA0y5tjhGEpYF8M729nwn9PDwlhk+ShDpI1GDXbiTzp2+xQc+6qo
50DVA1naf3poOXflI7yHgF6/IzKdQQ2OGopIaE3SdUd+xfABJ2nd+EC8FMiqhS+TjnWmdVZx8i32
+6oyyYD3HB7OmQHZexbaXxK0kTZucN5E7id9r4W0vs8hUu/ucricX31tI5G+xYu5pl7puO1fP/6i
OqGLF3xfLg6gG5vyuSEuBEQ9Mu8YsgOf4Gew6dEklBmVHS4h9nnTnxebzdeUHa4AuL2fXqKsq/bn
9DeodZiw9JjpEKSnovEGzfUDylge/lUOxj6lJYCSZS2G5+DS9RtQLFvu/dDYH9IOSYkWjGbEPa/9
lMnfNMdGTFQ0vkwuFe9SIbz3czOzOOCVopM+H6kS7Hg49TX+uzZqIRh5SIY9DkghgSI3Q9zAD4Et
TyOHn91jWpqeg6U4dw1m5X/m3aN4zKBhqIZRRyLNf2WvZ0EsaLE58C8I4v3Rkr0uSxP6ztbUm6fx
p+jGt/NkiDL1jZ0U5ygh8+1R21VwpAqUXnshyPfhPSOx1l17ToDcV+1z28p/HZcqQAyj2vwu0/e1
d8louJJXgLKaAV+o8V9fDSSNRun7v0pxWED/cQeGglfINEX9Qyx7qmyI1k1rty136XaZrE0VOijh
A0+pupxoL8NOTrKIgvzkraA3Dz4XB+16lpV9Y/Ju8R/JmeSJ2Qp2loCqqMWlNoGcxCDIQM2v0OMO
2ArxnhJXuY8AlHGAKoVfOJjE03bpEZLN49TvEJTqPXkwkkOTAI6A87J/FoIK8ug93tsGvECIWWje
a+Qzy5diO+YSv9Jzx85WaoGn2+aYenVf2NSY1wUgBufgpAspczEqo3KmIeepTjLYjSoqv1op6L2J
C+q6vV4/sqHLL+hystGZYubtKczOlNnKfW0/V+Puq0AGHgrf2qS8hkh9ilrR5OFUK8H9qO6P7pJ/
mRseiQquHU8jrtqolbtTerhspYtyyhDAmmu541E35hV5k8HZPiqDS8wBYF5ebpTzwNrd0bPmDEJf
7PVTEdQtYvG6CPoGDsiT4XJS9NI75aVTV72yzvcmQLUqp+qVQBqqqb8nqSbwSgtoYylHw2OpAJfb
tdVqLb0S5bQxsvyD5U/y2+ST6k4VmqQgohJzKNBTNkdEzKHID5pMZHgjh64ideLA5221rx24DKum
DH1Y/twyu55MNpzyqJPEzyM+X83PMjYoWGKbkzPZtacJ5m7THDKk1E09h12qW7SD424zRauot7xe
L/W+pVBfFpwd/Wh+MC17QPfQW5oAG0qxFoD5tfpG6ZojSohM02mW84TIe0gIfu7512KERMewN+7s
mbBY+suVp7LHMiM+BoFAVr7wbM2fG1gbtatSXNykFbtjg2YDrG4pinRfMG5Nzvfk0I32xBZQPlex
+exEvVvlvO3ViFcgNqtmgjHiTeY/SAZ04B6A097hzqbsf+z91/HCmnf6O/E/gUMIeRGeEFyS2kkZ
8HVEhHeM2OvAX/lPYRoNPVWLF1VhCA1HAePFLKZY2wflMWU3FUJwdF5A9Juhs1+nRpQH4QToCo1V
PpdFeZpl1H0yy++n8HP5gSVDC5cNj8dyhhPHwoX7fxup+ylqsLx/yQwm0wSmrlaQCDm+c9bWzOPZ
4zIC1YvS7qEpW5mR3DDzx0kUMX6HUef+2MVbC1VpTd2r24y/dwRQjBeFGD/rMoNCcKnSZIXJNnM5
BxcM6YcuEboKU6GbOV3fovgM6k25WTWQ2smZ2nC0Zy8ElSWho/cUeC52CxqdYBdEhTdF8GLXgaSh
aXNZgACLffnKqyBwPUqnvMAn+8gHQPP7AtFQuWVxIeP0ljMMWIiZzqF4llLFIS7l8kMT6o4fEyep
8kV5UuE6aLYF1OR1wyJQYqZV/5ctl1Qr5vvUNIBSO2g1CR47H4/mmg4ocRs0HmXT5yzKMKmKNi6q
h6JZxzQk+7o1+vjjxun7CZdV6rGF5+Z9OdlAefkv4nUt7rqm2iGybzkD0b0c/1pM+6FoawG442uX
DUCH3FXJocXpba7CFV6yMOeqLXv/jNBC5/PISNmVt8Q171c97hc6+FVKEJiJzUmeloiChJu4EEm8
eyuB50tpCiuQ1Za9zclH3hYBY2Czx0ADGSgR6gSWxvFiz8+Ll9fzR4dXd7d870ft2msSRCKX6UHa
ryAy8hA7vXfJcVdRgwUt+SWDLadMo8RFeTzmXknQIvTgvWlXbNIuLkRwk8kVSQJ8i4jAxnEf+JOH
LrxvXF03Ig2FV8rllny3REg2/35rGHGv+ATRlFStwKKpwZR8Y53JlV2hJuuZVx89AAstzSYiwGAk
Xu32afiRWhJKAsZ4QAXNKLVEp517kUwlzE7sKVN363Wmdjbst+XcHmH2VObbIwdoCX0A9IfDFkY7
FO9rKj9264M9JCC/sai+a3lJ6kpqeBycpIOuxhXPJ2eJWWMIBCb5KZ2oDombo6nZerOQwlVEMM6J
mKu5Lpd3PSLfzydGc8FcMdfldIssS4oJQSNJ06JusFOhdYzw5vwCep+9DwALEs28t8MoCSXmuFYg
ZX8hwvnfXtsMcTcuiHezAbFc7ciS+DnquvBl6GccRW14jniaBHYlBZfyTCFj7FUZ9MIfMCCfSoGp
QGj8VISg0RBVUU4JlRfYMayhxdwO34Iop807cZwBxBJn1/qlIBoqCpllYBTHCMj+xqFvl2j+i3hX
7u/CFuHPk6xsrG76VGBpB7wEd+1rIIoEYv+mSK0dE9FRN6VeaesovouAxXCXpzJn00uZPTgx1lCB
ZoQpFnc/Bmjc6LL/xRIvPusxnoh8wdH/RM5Fds2KPD8kk8LEbHmQAlcV1Zu42z6b+Xs94gD1lAkZ
8h80c3CYDuaSv0E4E5njWemhRpFJ+Jr20vGQzyrczPTLgoCFCdQQ7V0VVkJSPZF5UzjTjAFW5fKf
GhQ3elZcTM9sVXpc8CFpSJKLAfISGLdar45My5XcSYp4gQP76NAMMLGtIyMolvhfxPctr+Tddxbn
lmEKrHDlZTDmoAf+pGoheZepDK5e6Q9C2OXPbcWrdmPMSnkRYjwJ3CIoqwRKemoxEoE3r+KM0Ris
jvzfYMY5hsboCGU8OkhCZ+Nlshrp64E0AblaBtTbUZcLG41iyAfI5BRknk7YxS4tEi/n94niJw4I
tvgFRtXAI1FSWTMpTNeXPJcYvmml8rKLeGutqqsnxDBSerumQ1c1VuMWPUbxHUzNH+3/MGs5B0Z7
A3tlMv3uEAmQ+WCzFHh+T0xm9zVSTx3EaOVJS/jUfp14Hp//s07KmFR83Kcm9PhZVW7D9tmXQSIN
WMD4XEyHzEmA3WfjdXrLS5ZGiWbRJSCbvXX63RGq9hHJMuweANrFLc/ok8PVD8Jp9ElDqHMPhHDP
jW00+mC7OOQb/Yj8YReBqud0oSEWCembvflwCGCD0/8L/N8O538WZ3Bgp22rEwJ2URH8tJF7V5kU
pbd0P6tvbotGOZ+gIHrT58Y24UVSP/LG0wXB3Ou3QcRJwFzKc01TeA3LAQQ0d5CQgDcMfYsgMOpY
bXnSsw/3IU1dR1d9a0habEPQWkke6Oa2imL+DTm0FlTSQANcgDD1OV23cIIAXVifWXZtY67zbh+9
1E6xY5fyZABoN4kUq9yVfTwmcP7cVvlCBla59f8QT0blGNM+BKrodpnetsgLPm2icGx5LG5Y3N4n
MfulmtpvHOscD6CwoovLdyUN5XL3d+aKIQ4+0FZoLbausR2ueHWn0CF8yguEPg+ec5d5hXcp3vcq
Fpzts8V2ziu4fkE/lnk0tHTFUjTyEz76buzDmxxTw05QcUq9SNus1lZZi5HTzM1MXVWUu0u4kF28
93Anljv+0TNIfOXfpQZp189AnKbf8x3PiR04uLz9ADVXFq/1ylybfcI7T35ZEHbbkfQo8t9DMLya
G+TYvxUB8FWfvyc+Q10kICWMZsNRXE6LXgBxD7+ImOgZNSyAOHsfdSWCklmCV0/QiNkib7GWrXLG
uH5DUo7fMN/FN9thp2yGvig2EhMZxXhNi3lo+gc58YJurWkSdyeqoza+0idYa+EqpKtoRWFkve2M
sv0QklDZXBE/dhZiOuM9UziZdtMqSvnazKBCnry+gg8LFbiau841yLuOqUeNSXQfN7ti3UmhOVRM
clSsfRVoeZ89/C7CVtMNN2Yo+rAcpIDm4wXtdKb6ghnLwzs3sCPtLHYs52OSTZj+Qv+QXqDFA1Hs
x7cq4ke7CHVVTxiXjzzKZHTw1oM6KnQsh4fWB2eEO0qEUEaowWNfbK8tGSlnkpAmCkjLXop49kRG
LCyjtQLQoNJiZWwb79oU7PzNUrxcBx1w7X9E1nyDBlOVR0svyujlL//vMxk6yhVQzghibski/lMZ
nl/+itnwNXzzxmMA5Gj/jimkS8LsU+DeZl4SziD0MruKsiKgs4SxNEVasfqpitpQxlyz+YJ9UrMZ
Z2mU7ISFBCoReOOlvokE3VngtH5RIiH7bxN7q22NKS3lCsDsOhosANm0u7vaV1rVpqHFkqN63u37
+1qhiUQQARK7pDGugpNax3Swqx6lYP9JXqNvZ7zWP3MaVaIgd60CMNaoy7zOVDVHmf/GdMi8FUzo
OzZrNcGbOluBDsDCQXASVqJyWoxWA8av1NZdTaOGj3hM+r7v5/tWkPVpnCWzAsTkfnQ+k5R9Y38L
XHirUGHXNkjFGg5vZ6N4f4Pgc4C0C3TpH9og12186C9gyLFGixzyzlnoSq6ZsNRIlJMdDdZJWBX+
0b0ysPTnYFaIFvjsK7ICngIR35xzeZV6z4qVRKJKSwJgW+BpQBCMrTsh5rMjhq8Yd0KRAOCU4I5Z
Jb3i7DGoYMHC1Pcpi8Ikv048FU+Wj0P9yhoTzjGizRIumqgzSNNKogJtp3yniBuT6tnJKKUQPSh5
zQHWkTuy4isa4SWjeHi4skg51RXn+cWFV3/lxjVwyKleluABt1TufNjgZNmfLPNqcFYnEQen06cS
D9lWXJUopZ8BhFdslsd8lCBu8rwmzOQu6KE00Xm9/GvHcan5Dvsbv5c5Wp3ILE6xqKK0bnMxFZfy
5HDHtLcXhAcnpLtZvIZXcyG7rP83/ughhRVhVx3JUps7VfO4i47kAnKdnqm2+GCojhz3C6d3rKdl
4aaYx7FLdKXDUoqbaTl2dhETXnhb+rExns1XIDXVq/bLQ8qHx4EA1HitVWYltKUPFnjxXbes3BYp
VviwXHrvDGYdgF1LQMSII4OzahlPUV33/3/CPsadJ0m5hn9oCpECiDoU6w/Kja54zRqU6O37+RnC
4/uEfuL1BHc+H3YJX4eG10qgJoxqOgI4SKZ9WsQmRgtVSjFewW0NLjBXD0AXCab06ZNRSIfCoO5Z
LcaGkiiB1A0JgUaKHWcCPVty0CFs45sLCYjaVe3ElyHiJKb1brJYewgpTxPB252TTWhctqv/U2+n
u0aumNywq6s0dcf5KlQlC8OW0mRp/I6NBQJCvWy2cMHmdj30REGUBOwLUXTROyvGR3OdftWbDbZQ
FiNxAxhi09SuDIIMxly5XB4MY4Od/4X+T7o6e/+2m9DTkqfgYSQloHsDOVb+WgO3J5iryWm9FG9z
OEXsa3fI4J3x0TlvhyAlchkGOaSs8k/T2tflTXwIqWOjh/2WVLyskqSwgQmjXts7bCF56RMa0Gil
zRfzNFoDcwdmpdM5uaCmoM8nNPNppuMhepSFm/GgW7jzg1rdGzTudhGOaSbULn0NxSUoeL7WIMpx
KU0i4Qw54N6UCh47BD9f6diOMmQ9t9tR3xd5OUd4kaW985/60m+KskHSC9C3H3oMiBhmsj7ofI0v
8mn5cYSJ/XBmZZD+hptEHov5XX2z/OztP6q8vGFKlYXMYfEjVXohDoojMoxLysLXg+YPubC6kGCF
jobBQtfPwjpbSeGyJ93rLijSw7Z81DzQzuysABponIngf+UmNANqsQvjXCT+ueGr1DUnlgFnDXP6
HeJmG2P6ry47jBXEiFSmwl3ZIxUKp4bCZ9jU0Wc4qYs0Ire7w/4QxPyI9DHulWAodQ8fWb3d5yzj
yexllua76mzMiTUoh/SMzDD+dGYTkNYZ/5P5wDg2NlVIPfST/W0iDyIf5b2J2s+p5ByfewIP8I9A
gNy/3x9dI9048lNpdVt7iThn7GkC+d3KXwV9IenqxiAkrMnRCXcjtJgekS4BEyEjLLybsEMhfRhg
lcaUsV2T6i+LHGESH4o/Fw0/jt4MCqZhabj/8diA2EaiKLUczLuuoMiFT96WKyEvZPRe3/odo3ge
Fq9cJ7QhTTOnaJsHvrtRC1vKtiQ7HD/aphBKcU00RE4GP1M8JU8q/lZJXLlS+7zgEV0VhMTY0Ldf
Cu7v1TMIJk0jErxIQsciYLkAB64yqpj4KyeQqCp1njWxbPGcR1f3zAgftPJlNe6C4nQkV+QRISiM
IfE9KPfeff56/zmbtnvqKqyoVQVDLGk/ulX+KSb+2zIGpcOdmw0WPVoRzb9WaR0APjr9QkckQ/6Q
4ks398Xl9nvRcNhbwB0Ah8o4SMtChsvwSm96zg6SdPNynExqgEzKppPWwOHRs5/b01Wv/pCR0aSQ
wUU+3hCH3dB2mKYpTrPIoqvRBJ6v1HiWcsGLF1zN7DnoIw81V4vbQGq16Bt9zf8PJrVZx0jqxxkc
jrYgp9wc5diW/MdOjwGOik5um1PxsYTFLvV/MdWZiY4H9MGTwDlBK7kVgwb8Fxdw/A9/I/IZtqB1
W7GYNn7iEiEjA/6gCK3s1FhtFSxwpMOGG1UkzkWefCGZrqkZmOeOwZOrOuIoRxyKeG9xBaskedwj
57EF8hiodJG00i5FWPhDyr6CszCvmRM6lepqUWrP1RK3FC1j3fWjqYMgOMSPX+Ld5aBffXrCBuVS
V354N9qp6rvWZXut35bRWUZ3L5gb/Hla6ijW9l1TqmZq+kNFyWgfpyM/S5IwKQtjN3sQYiq0nNgy
mEShsDUVrk32BYS11dTUY/STryOBsI9N9MGrfVko4mrZZP4HlxATZERXz4XF2pe/qN2bIXufr+B/
FC00FD5zeIfX7z9CsRjjlx5iGNyq64fSr3Pxs6Q0aK0AuA/WyuFeN8jgdKhPf68QWF3E5O8CGx88
0Nl1aSzZdFdCHAKfv8ENG4GcgDp7kO4QbEyDcm/IcP+R5vrRU1KX7Itc30c42arYJRVtKvLAkWjq
rAAQ28jHsoDIB1tJUaDp54pmsNzl/7b7mTNqnPLiNcp7TsEHKlsJGblPI/ByNJzZwD8Hu6dDa2Tn
25HXs7pncqv8yBclcvYjkS0L+U3cczo2DWItFCf+CmcYTQ2T4U/lsJJ5sNGYKgXH+OY6QEm0dIl4
VAaCn7A9181bH+jpPExUXqUPNLp3L+5Pfei1wa7HL6NR/Rcap5Upbfw/MhDXGLBSDYoG2cFGXjlm
PnOtt0OsfNFNL+OwUAOO8cDT8J71Ihcq8mKnKYliC7H3aiUj7a8NmcJj5pnxzdyEOft1Xx5dHHdE
BNOYphl5pNEppkMewFVIuXTvQmkAsbQWq+/L2PT2I/0xa7dbHbtbFgV53O1xI6f7ngg/tmIsstcE
Hxt5q/m2pKDpecVcHB7ccqzYXmXfWPdLyqJjSMarnBYYj3UUvt8TAc7bCDZ5riqUSlWq1xQenuhv
FO0ajTJnxsjUglj1pcCVcqL6YYikPyZJQOLALXeCL2nSsbik6PbbLWpCb/ZTdSswuAeV/ELhXiTg
sjE60WdRxHYQFofGJZyzy9VKRQ8MT1hCTAwWrwADDrhsU4d262jtjVaiBVxsJkkJZj8Epr9jf3Mh
aWfha/k9zZ4fuk3RjFnO0sP1/vQB+u4ReNXS6udbhZaZTAgqlECW2oJXDFqfqle1TIRvl225Q6et
53PYkg4WM4voYaH2yDcgjmWbhgKHPDGuwKESlh9fDBrsblPR6Q14ie6EI18eLKwSK0ukm2j28Vre
dy6YTNAoG+0u5XEVPhnBw7o8uBFPxOx9+LeX3Ko3PHWU6amv1+FD2FsgiFDDe452ZlO3JBbYpEon
CFGJCiPykEuQ1n4vXUHkF+sqeDeblTfIMlpEke36fK4a5GC8XMG7e4sytX+YLA2EawBGdiFkyKYr
GVj8A7NYthNpKLRroR2y6HT8MpaCpyNgcHP2sDSy0l0K5FEZEOMUxZB9+gRxHMm5b7U87NDjL8rS
7QYP55IV9T+mye2BnuZY9ckkWOIWnPoEOrmRZItJB971Xrp+rDFRteOJxElM3opSMkDTRwHcLolK
WUmWMUv1TjROWy7BX6qbDtyfF+PeZozQsrKUGPb0obCcyp9Cfd8gpteQwIIdz9zXSYy01761mgZR
4oUIyLejh89OadwVAGe3emclo3MD1gx4UtlQj2kX33QwzYA1RKDPZjBjQ22a+I4GUimjB1pwhAkx
MTXaUNdb4XSlnxuiibfI2q4PiD2Z0dWb676Dr+qQVpmSeUcdWrq9qiywtzd252n//H3aPQ9e0pl8
xHfBgvciJCIki6OAUqkz/OXGnmCzHeoxkuQ79a2sowy4ROOTaeFY7mUve417w5Grb3yUQfj9fJQT
lbb7YKPMeoRyf3g40mXUt6gPVC3GTcFbZcAmrMmzOPlIskvg3KW48xUbMGyA5lakX2O0Z6XS8aDh
1c0Malhh0V5JtRJ4GX1BAToK1w9G7UOv0ypiKp15MCW3jcebCkRu/bW4N4zaCZ1UL6ynucB0kKmi
N9/ArQNOMFaH16WVDNwpqFMx303QZ+jc419mpb/xJ+siiM7kxLM+AyTJbZi33KoNgx8WuR5Pd9Lw
h9psFcdgO9k4eN/tTrzSDUoiH2Teld3IK4JZUxBDxyGuI7q223fXVLEh769ddONrUYL08eJgvWHN
uMXcoM/w3E4NBAKJlfhl6cButcMSSn8clroK28+BKDgEu+q4aJEW1puPSATeQQ69Lo+7vzYcFgj6
7+s++yN2iIzD1Nxcuk7O0uSdQYsJR72dJS3BzLRnbltrnKOml5qjhnSkEjScUKHZuWFth+/07e2b
TXBzbXqVFTDMXZH6d5R7eYvIetgS6ueDndqIx2mtYEh1czkRKjVmGe2bZ/XagMNB5ORW0G+oG+uF
EOty/u/G7lA7jKtctRMRsC7WPLq+s7npNSCrErEQ85SdvtGLu9NLUxYdyEy7E0Ryo2jFXEUD+dwY
/SFgRWQse3oakKUdsgm5q1v7x3saUr072Xx1HEWyf4GZ3XLy4Ybso77ZPeE6XW+zktbr94sOOnmw
4Jjx6XWv9WCihlmO2fzXrBHavrfj5wdLWUUnz8wIa/h7pYKOz6TERUwXvDE+SuMnCLeBf+k3OSo4
spzaxkAQnMwnUfMAxFW+fQ8GMydOTa/3NlZjd9vgMhjsEoL+vf6TGodBTSeDsqdsAbzkaXkIOwYv
RIHywxX9II6Oq3iEdkioCHduqwW/ZQdQiKH8R1A8hR+a8IZAUbG6x6KKDvizg0M8wjDQ3Ht2Ho9b
VjjcHy7lheEO42AfMkW6gY49S0QmJvWYnC3CnyXomSCpadRcZwMMSt9LB51iuhmbppa82wbOajhK
nXoOcmSNzXC2Az9q452XnD5Vrz+XpxTQgt4emGeL10NUto1p5nFeOoTbwsto6A6GvQbXwGBJHX+2
82YsSJ/DhLCuCbc7PLpPnPNjTg38Mxap0iTvLV5LXvWovR8WoPusC8+zo7fo7RkUEaOTR/eX/JPe
5SsoZT2obh0YmhfLeYgTtRXNUzT8Qm/8W0pXpE4Y+TiSfD3j0U7wJDd/dt68+dRVLk9hQZkXzdnw
Di4Z8BhppDj41mmhGQjkazd8Asa0BhcMW21hWxQfoS8LU9lUoCn1C5hVADtfQ0cH8vlQF9MmzVNN
KXW5f47Z1ZuYeMLAEuPiKTFKK/0YGQbFiJ/4q7XkGtNU70ZCUYRAGl7qQB/qOFXWF4K/GpNMP7iL
7Xr9/7ekaueworXAdzOtHmKCEiRzSkr5ijOWJyhrnqZeaLyJ0mMyaaVvjiT2TAgXrr7pnPxrebxF
WffLZNEfsA/1Iiy5rigShiL1eFrUWmf/0golxPmManu0r70l6YjaUebSZeU0WG+MWH0nQ/+glFqB
m190AB12RetaY8g258k5T7Zj5xyhV4UAkMY+2UnJlwlq07unKBe2OwBfM8ODu9U6D1pTu4ZeY7DQ
/mo2C0LMGoURNPN+k7+XVpXLfR5YMZ5KTTX+fivsSG3AbP2BZN8nZGQ52B8UA1AEVfCVROMwF0L6
yyrQhtx/+/vv8Z83nBihLPoP7gHOKMe56k+CMcjaeiksoOgXCefvNshBeFIcPv+3dtvgAcW6/1tH
cxMrW2Y1v/3jJRt8etV/uHlVj14pg0rrE501yjkkB8P1YDuYEsZ0hnnqECK7L7M4Vo33K9A9JCIo
i4vRWFh7dr3ReW7d/FS+EEyJhXyOdzAqzM5VzclwDib6xgwQAJJQ2clfdb4L4fWXydB48f8zmAw4
bxICMFc/XFDCcM/+mXX7XlP53OLm6lxZ5NZ/bU4CaDH4cb2ig+Lw6R9TqR9xsGCnlBpwMeB6/Ufc
yej/oKeJT2QC0wJ0peqCrDBcfmtRzC3wtmB/5pMbAYLGFxO8Pkn+TjYYSuX4prBUTcb9Hd/KzokF
3S5AxzKFqwim670vt4rtU3m5GkvagF5BaJR9XN7UOWThG/nra5+xAFbU+/M3GZB7Q2ka1oeWGFYN
jOUTPRlqiN1d6xu1+AFmO8XThY30/u5JCQ98dIG3eK09rKSBl04enbkuJZZVNx5VLUXZPp3iwIfN
m4BiJ6UcOfXrhTHV5yUY9abPppvpHGjT7c6CsmbZXq0FddjueVllmtByEiodN7ILwYYqor/98Oo/
AFxGRcSx2KCupgQ3C7PfSmEXaZfo/JoBf7r0O/5svhZ2Mjw9bf1SKZLqbFOipvdGwUzl8UkA0b7v
ixKTRFpnjQeiYCuceQCT+kKrTvgive2jPVKd6twa/s6rg98LiITlEJii8gM6YdeErmK3RaH5Omis
cleqt3pxdwwJAmsgLvVnPd9dQ6hYOhoGJN7Z/Ds7ID157eJSy7bOdhxHeDlb8huzcthgbJzNZJnw
N4t/OW7qf9oeANbufKdI6/R1Nwx2+WTptySoW/dHSoFJzMQfNv+p3sI+DxUDEkBsThXqHNzuxRG0
7TbnRLPtIu+lF3PQUPnWMx08yszgIzW4QQv2p4YGh20S6zaWpBkObIS05G5kW21e9E+RuI7mTJ4Q
5OmXZAnzzcIsRnaGFFom6jvzKEcqH9cb+XLSUWJDdAq36zhD+ppGuAF18Yas07XJlwjHPrfvc2X9
ws4iKvjf3/iLbhDIkXNTKkNmBrvwGqGAbw9YprKWKucGITb2URAGVQhR7XFpRGtvPpnQLdufc7x0
fcTJSYPfhXy8qezQacUuCIWPjoJ1lcv8CQtlhGTYiV79qVf41LWOeRMoBawbfvBiQ32ZpqwfonWH
J3A43UG81OIAVWi4WssQk/jOVK7HtrUdcgCcH2muJ8vhp6cgH7cEi+9V0/OwCDBOCMNKKabyIehx
WgOj2zSb9SUZFMnVpR/xQ1ee7pb1IB87YIiYbyovKFhPP9JMrHZuhS2ukbMxmmK0VYxaeVc0J1oa
/ei+mN+yUcWacQeimHo8yE9hFx8eXgIdPZC7x2Fp2doP3Wl7yOLMTQxmqvRDAF36R7Lk4yQY2bpA
I1/tLzp6LABf7kJbalffLAbtRE6PLcQqJns1MxRXvtYqvW7J+awQ3uB0zTgyqGmdh8+4/NAHDO4F
/wOuzGjxiYPf6GPmG/MJRKQAZd56p3vAnqNygwnc+RoeWeYjuDMMCmbH+iYocSN8/no0DtODGxwF
Fdy0x5EmLa7bibmhpD+GJDVBRSIkw9OOWTPwZsd3hTxB8RTZarOYPFf0urVytQL0OM05giUsCoy+
849/O03BkoLQ2mC6cJxRMnkPh/UC/ihqvIKO1gMbxXdJy9JBG/qgaFD9XLodR8glhhqa7tntTbFP
9n42C1UN+U7qVXDG7Bn+3UPfU3WAthiH7g9OeVuXGOIhgt2xQR5CC7e8z0wm3XOo0jZsB/blXaNB
P5hkVYjAr4gCNzPN/yrKdqC0qzBN5Bx4xto/irU0NXdDdPboBOOWRW1CDRX3Mk9pxM/24r16V/i1
9r7izDN5pP5DaHlUEgvpr9efHJFigiINL6YUdm97LPmQnzAHbsyyAPMY0aKhB5/oej09B4WFeSpJ
iHOniCKnNsp7hp8dqEQeVWrUUKJaLn1/hFAFIAn0GTAY8QzvGHhOZBMvvBoOuHVMj8Ix/Irhhrfg
cpsZLYK66g2SlTQtpF85Z6okH4oEC7KjHVL0wamZ5folj9hpVhQDGoIGtu8z+2ZcPgMFsRv9jXZi
VslVVr7JmXkOlmbEvIEfGPxfOBRxJ1Tqos/D8VXaXAzHWQK0pm0acZz2Gc1QSAEvgP6YOf3Vb8R0
0RH9uNbJhbP/Cif1Iw3IrWEXNhYkVC8cNaCVveewYya77jr1jvAReYM/VCJF31WMYuExWuC7bREI
SZsLVrNy83bu75Joc0PkQE5XaOOjk6MU/h/xTw1/jhZVhwvk4EhYFY1p5DeUcj1720UJt59zbemc
nh5LA3lxgt8tcck2roeyRXOtAUepUgI7XQtdNQs8VzzhsdrGuEfE3lR3OS15CIQPuyz/C5n6YTLt
BndvvTkfEnfdaby07BN1wllWETiL5gZjRbxKJ3/pyu57Nicu6OFyQX9/h3DyOoVkaFZi3gECR2d1
vu7e3dN8ohLbpAAt7jLm6psaY1b8Vgs9t9DmyKMiANkXjzKGMdtthP2U63FBkxUDI1jNeYRdK6oE
PY25T5PpCSDFFKBy7mbW64ZJ6uqtu5haXQl1P+/2xFcA2ncAaSsNOAjT3f6hQwmRUJH89HtYrvew
WEDBEc39g/8qZdnFOF3t9OUlVOOvkTGFe5b+TjOyAjORDT/64/jP8nF6OgE0GJncQFlZK/4r/4Lc
fiC2aJcOv+kuwRck0mcy0Vb3rVx1zSoNppLuWdNfp+dAc+GG/mQ42LUD7Vy6/hIFhToMgcwAktla
MTMZy7mmvu6n57uOh21yrcKuQvuf6A1v29PP7fg05iNljkDX+m9SjkEQbgyIXz0HrNPGjRSXlX8G
/q7KPFmxGS/WRtxFNxpVk+b66gnAmcMxrCDYmEpsiby2MsfJ0R2OF8pGpUx4bzG7S/q13ZBYjRiT
BN3H3IPd3QVxzWNh3+iXikBL0e3VOc01SU8jYo3b4aukfLKlMqRn/C7LVtAd5qbppNm9rSRHSh3H
JcvdXuSXQeWNdtlgG5ME+Po3n10YzOfn+jB9zaxhgniKslHUJG0qaEzRNyj2IdQcQEDwINXUu3Gm
wA57XV01aU+NbiejiLFQou5ew08jRgklbhsXg+PqbeFqRhWX63fpag2dFFvk7PVHhciwE9WNL6PB
6LY9w3c/AcAbBGu2MLdWmlb4opF0AwcJrCCl+XFfDwQjbuRmRpJ5BHweye4ObTRSdgpASxVdhh0S
HDdGj4jFYC4ZvvYLIozLLm2qH5vvhS8w3/1eolLpoDk9jRe9soT2c5SErOw8vkwsyZ3Sp0PPKRXL
Fc11mig4z9ZcSkSu/tqVjj0oT0Tn4hI4wgfjIeDd+/W9NinLfJa6+X/8u7b27y/m3dIRAKtWB0oD
CQ9WuFA/bzwBOnhuWJNmhVSJuEZnm/mi4lLH/NfzZwLDrwkk16EkubVm/lSAUgVHGKP7MTts85oC
+7ssRwL2UPc3JHU3zlGmvQ3wSd1SnQBYJhmqLv3+zPV+5+wCtrq7pEEFSFcj4itt4KAs88FJ02IB
ZEEHzuNDJr6s3kKISCMOdkN5a4wUFCcBeZCilXdLcIXzMe2LTPLJ/33WVlZdHLtMjR+3lB8FTgtp
9yrlAdZ/VXTp+MSALQdJFuODyCA8eRKfwMvDm/piUfy2vHFqDTLAFllIXl3wvLZ3ka5EEOpi4Uzq
q/6NhUOLaLP9xOeSJI2JeuMQb1ZuEJD1AdxFh+w9uvUZMp2UlN7dqtbm1IvKHlSr1BmiV8EwuHJP
yXMuWJSQjGLsYiCCRVCYoCcaMoCOVKAI95yHA4Bzeu3SSHrsNdjUUa3VxCtMvDkWDPBdq43g98VB
kQ4t8mFAGCsAZmH8U6vGH0/kSjzI236wh5wimiG6nXdj9LtK3nRyrrY1K1gwou+x3ERhYrXkAWb5
xtBhcik2B8w6BGOZM+eBewh4YmV7vBzZpeglT13ZoRI6UIkO/fjK8oRbgc7AbgEPIqBVY+PTLzKt
7TrFQ860FWx2unjk1sRmm8Tzzb/8D0v3WcZcQ94ZxjNb3CD4OkmQQYUhgeSlwjSu95eCg/HYEpWo
Px1djFaJg1tA2I7PCjMYTz9HE0+TuADQ/bQpUlhNtKQiLKr2p/jN1s4S1rFtZBl7RrHhLl+LrZpK
mNen36T9QZFq0tlMzgGe3oq7mhVNyeFgh104A4RzT1YUJZYKi4H/hrQX8FpuaYSKmD4be5PFJq9w
Rxdd1lZXKsE8KVgjW+HlTqiXhjj7BsM1iezmin22h45OMwUAutJHxuJNiCMTRQRbKq+KTMyIWTlQ
4Pp+a9rltGCR6R4/v+Cc7lCUQsB/LoCjO/IhxfNY51CMc9sO720T32mCg9RBO/U+/Ryyli/RxdsB
tzO5up+qWYYe9jVggBtIIdvKFF4q0B8O6V6D4VAAMLSYYCBh/l73tGtogfQWiNsrsvQKUv57j5Lm
P1QTJVCqfOCY3QkAsxzn+IBPDSDGZX6J5k8vB/j9JGob/nUXW/I5AZHHrcA+hi1t/RnhmjYA/G3m
tTopRoQVQYk8DDLe56SIipyawzbliln0NRG15dUu4MpK42M4LTbnBP6FNNiFhy8AyiboSZbL9iqs
AMJW5AHiswvJcMjv+LkfMfbd74IybjYRFifY0zeVa9/U6AwFFGByYzuqFNE+OChME32PjyzYKX7x
c92KOENmpAocErh/ra38B8+mi3x7BZpkpNfqxNt5Fj8dmGQ4HFBuNK4Tlk7r/7WEoiMnlpzFYXmz
GTxyAAbiVbNkiaKy7JFgUztEy6CcHl8aQ8plZO2XOE72CLUc1Qt1NfXKq1fOESuXG13Gq8kzQ9dB
/eUwv9/XVruY8fOLfkbQa/p9wnSvWVtfQUrh2NygUH0NQ5foWV3h0eYOMu8oJIbL3E732oJQjwdT
MDr0BfqaswFFYd+MQhg4UcIFnKnvBzkZCzdhJWqjLIsnCdNHzaesoWR5TpDWGgpMYaD9bMPzf3Hm
hfKSnWXkXvKajtL/JWSg9muKt6MF8sCNWO3I3Pl5VzZVpYSd0HD/R28z7FHEKSw2bi36FnUrE0rw
ozXhFPh10iGS9ssL82onXa8CJ1M4pPNyXHxUfeiNDP2zWpODfhP/qPKNvDM1X90RfSRLxgLKkD6i
fqA0culvcrl8rpHjyj7XReG1MuTF67fwUsi/Jn+zdPVZd5Em3u77mKKjBOVQ9tbzegNDquGV2Swd
q7XuYPOEdd/1DEwQcenxkr4oHn/PyiiSU1bTJ7x976iAcLYWJnBnpqEWXfLI1LWFPejmQ7VKtC1C
Up2fPNUCSK1+rU9JSoWoLpeWXxoy2gFE3nSHlJQb6t9wZg0boONHVwBGC0xATRuiWGt4i8c8qfwU
au8Iu375rq5KNAeVFCpuBsaLTCVcowD/DymyUqFF9ofWeKm9taGI2AXpdCUl+fPojI+u0V8JmeZz
LRly8FJxEtDJHmjguX7M/40FmKXlnENpsggLS/DbtR8AXFPkwIhqbRNtdZzYrnkJEz66QWx4EwX1
o6jJbgEPttXnzkwB/l74yYVMuKC3TqusbqMXqV1Vnr92Gb5PcXQ7rpQC/6CO9ujIWh05BZ3F3O9r
5GVq+G8b6ckV7jFP5L8Ef86OF84faNCxV0Y77llmWKPzKvvGWdHL3t9E1bQylBs0AUPkk18qAPX6
7z3tWMD0Hh3X8JWADkl4ZWC5ZAIh8QV1n4GE6w51jjJR+xOh/bM5Qbq5VOYC83cTTvxtRH7I4dvM
IuaJKxBbwBaun7wYNdWsqLlsam6WThY2D7dqg/OrxMUe6zGfaf59NeF5V379sJP2f0X4KL5EHWPj
8UeXB4WI4Q3qxEJYruUn9P9oouRxO3v7QHYiZDNZoK574/ZkoeU7RII1XQ035q0qrfezzRc+fQeb
eddR6WiSiKz9dRaGn/2+4zSwJ36lCmZVyrSV7Nbz7aFppzSX9NTwbiqXzWHwA1hMG2ehe6nZk76+
c2tVAYvim61o1hnSfvIbigrPJMn5YsDp4OtfjA2O2cMHC93xodunri+KI2QVBleB3Q7uJImTWaiP
nesHgwSiDyH1d8haW7LykiyJBjbs7qMIrvErNSa3+LG/tx13kvziolIoO3mlnXAJz4j0Of6RALec
YcCksrUGifojA2yg+0ZWb7FT/SlWaHoUst+aZcAQwlsmFDGrdG4BQZmXaYA92WiEVNCO1tn4uiOR
XbqMkuPqoK0siQzTRAPiv5d9IhyG7dqa5lmv44bMBYeXTJglnEgnIEgc8TntzBIh4837eOXg7YDH
2h8hoOJBbHH79roGrnpQYqRUBs6B3O8eBimTR/rwMW8iEvei+LTNwhZqWmgxgQucqcFTpZGpN8h3
hidBccfN4rDK19cnAmhMaJKiqxGfwITvvsvqLbhOs6fSTc8gcRBe4hr6lLwx5Bpdt8kBD8NDsixS
CS43mXdNBrliWX+MDvTU+0lvETw6vb+sm1ACgKLpgPqIKkVzvarTAjWvLWO9QAWqwvjt5IxAYLwZ
riEUa+wp8xv7qHib5NVgQGfa4ZozKsYUKI2okLqFN7TdZ7o8zp1qzTKTIftHgrtdWNoC2qwoJYUM
82p3oPBK/FwRES1BVyY6AOzd2RDAId8y9igeyqX7sDsLPk0C/zRNlXz+G4BcgAVzMC25c01dPEIa
rt5Pb7rFq2tnjPi1QyX0UNErEqhKEHSWKM47qNZBi9RQSyaFugtJM4SjTBvcnvfg2qY8/UhKLuFa
INVUsym1nZOZ4u0IQxzdZLttZ81RHseZ2PKnBv4VfVMbEIAIHPZuDQuR3Q5/oe+HSHl5oGD2dqP0
NR8y6YnGhJpsNd02W5L1fmWBk5wLagShAE7SxBurJ+jmBKNRa+dZ0rK6fDAWujgPjPZJHQwYTd9k
1D4BkgOB59va7wdE0V/HvC50i6tUzbGUqL+rpIbdU14dJs4w0HwactLS2L2dBBIRtCdXEYaH7hoU
oTzdbvwIyx+I3LBUP3TA5elTBn0eAxRUhGHrZMnx2ktphmsx4auRTVfvvF/uIPWKP+Iq7CZWthBA
G2t3K4VYjG1evDuTtxReLV8EleXRZx3sabQLuipKN1fk8T5LE6FDvMpTHXeQCaYA4VAgnk2/naW8
fNcS2wD4XKqM7F6II3hA5szOJgezyYnOXrmyGScY20BAirZTmRnNQQMoeSE7+nhWt2oIVPC8OKA9
/vawKReN448UiaHUDZnw8p3I7rSKRuZ/4X+wMQEpHaS/1xlaHA67i4h3w+yEAzHLysLm93kC8fQD
XrC8FW1ohZfDloCd4kMfZo5QnJfCWG4IZae2b5OXxhtr8i7Fy3vSigP9dGFkLf6rREx49+r0Bx16
zZ9dbqi2RRuhXbNW/QMQ519eB9BZIlCyPTf4sPQlZflbI3/TZ7VR5wvV55KAe5MTpBwvfRrnwRhA
fojbbA5/UEerL449ICIUO04QfkljBq4i9HG0jAMT7OPFFpofoReiUf7mWy4ji9YIKSh1BXESalKI
G9U076kQ9FnKu6hO5bKKtvjxV1EYuxbz6WUF0MJHcn7tptJgfwj942A8/tBE5vtgjKUBbXOtV16C
5e7MbWI6GpMOR2XQGgltQD0SMzSocFLxL5qvPWBqeG5oV8d8lFJfLatLRaj/aEHKCT6O9knLt2k+
jBbUepu5uzxf50cSSkDaS7Rjy773+AxUKMGUBNxC4vCU7buld085l1nIwx2YMbiQB44ZsZK1W83z
OOlFEE9bNNv6AgOaGfvlarvgVi5i2X1VeRCyo6PvSosM1scKtQIOIor3z7gSHHoUyPqSaWQge5Ev
lmyQn/7rX/Vu4kISowKUIQyghxxUPrzN9x8B/YDIRManN+n80MHfLAOn2yGtZbHdgDuJeov5p9U/
EZTzOpbyRNzhEzoDNrRvUpl9C1INx6iAonROQZ3FwAzarMeF7ym0gIa+i+zAWsnHSVACTgtivDxp
WVg73qSjbRW7G29IKlKsKFqvIXgMkNGkrO9g3LnhTBjwCJJLQFfwZcaXZotFlM9arvkutjfeqhRF
AwLAqJFAVVb+zz6yranJMlh5Yff2EHAk+y0bFsgI9FE9dipST4Uro3pb4gtwpS7qcyGWTUdUBZEn
MiQR5wJ9S6z8CBBirXs0+X1NDYWOt+paL7U0GEkN4MxOpu9rJS6gca65+HssxqAC/eVsHB7w44sm
NfJNbhJYOw4xd0YrphkKfy/K8nV/BOtdyxHp28zfBx2NJpf06kuU1la6JDdXLnS7wqAGBLEec1fS
BBg9zr3cvHPt3DFFgPLH4RAaw4a/mA/6DBj+bzSAREC1H5yTU4YmQ/uoq8Q3kOoYO2tWHMOpop1O
fQgVLKiv/W0ny2Qi5/qp/vuW7XhSHUBqTg06FKoqsjUcQCncks9aD6HLVPZ8BNvTEriOQHDKl2+0
2+41HXtaQZI7L3j1OUrsqlRd+a005j73psPvdCPGf2LW7f6IkzgHu+Dnsx+99MkcBanUkRxyqYt4
Fb52Ov9OpYfP3x0icGnn+B2GJ6lw/m9e8enumBoay2NNICqzWbJbZ3USjI4NSRQqTfscfc8YO+1p
hjfC8ZEPJgEO1fOLUU64i8TrS5KUrND39AJx/OYbYVmfK1yZdMT29HtU+8dZBLQfvUCXLKg5nt6P
Y8KaKWO/RDLIXbsdMWE5SoJnCW4Au8exL8ZJ+6nUs2ReCmhcwNH7hJrw1zqv2Z8/DHubbwk7HwMn
0n8Rn4Rf2JcGJyH4PjXeBToX0iGJNqBWmZK/6gVYIk/hUI8slnJmSEnUzfl+KoEyx5QqaHUkwxJn
xxU8TjrRo9e6rJuhOy42yBq3fOIr+jMZZvAjr27MvPgXQmix4a1b1OHx6zYg4k09cA6YueVGh+22
9xvvCs5ZA3bYS9gK95mI8cwOVrCmWY8AvEORpDpzFDHJ0qzD0ur17R6hbAnF1y0XPAouxMcYqyuN
R8L8JdPWGwxazG1TEFEGanA1XD/2BgQDlKytckKlMqgijxUHQ5yk0it7YZS/VVYtegcmIwwPQOC3
M40bpBXYZTMM8oAr3YVMBY6lQ+Mk9DdksuVcAWngUHxDqilpUpRqTG0IFvoXzr5r09oJceeejSSG
vpj3GKTSdZKH0GLZVVEKsnnUH0mNfbOeHOCVZVxlp+ut4ioXAn5QYnZPa/F8/ykJaiyEzF9uLxZ+
Tv9udzsDDdxLLqk+18NIK0ifDJqKZFBMffgsZtCye0E4y+0uOFXW1JMdRz7VngVV4R/6KQ1AKiw9
QM36A92/QdiVK6KZIXGJPZfoCV/CmPDYTjb9cQWAWxPihA4yHqwiFOpwCwn+Uw3ky+3vXXEwP8+0
cLrP7ORmA6jJcvjoEatCEDJzhG9a9A9TLFQHzxKgkNLM+cgnoxXvOWufToS9nHcvziokAp2mXoDr
8mL7WVNtYEPdg02OTASFGrOKG/8OBAuolGrNvzhcVQtOL36F4DWo8ziKTr/pxMytkIcTT1jgJHNm
bzxSTCx/WGNQpWYvzCfapRahZ2sv/XXV5YAp6B77kEgPMy0aic5ccS4TlnFdqdtw1HoJnSgLaK+j
UKZrb4ehvJ+9pKpOHUwlRh5+HLZwmiSCbyV50M8TykwBiagyAVPqInwcjcujb8xcJjZnYB9Y900r
oq/xRzarEtADrt78ZhSwtAIerXLV5uRQ1xRGXBaJ7suDVgqhX5MSmYDi1FGGxg3L7wtvx5EWU6ES
r0+KAFHVv+nanuTxuNcrw5vWmBwnghr7yduLiupyjgJ7os4cS3XGNPLhVu1HF8HoX2q2iMbmPsBE
hBV5L8ycPAc/0hUnaRmTqy3uupxboxzsVoNfCvPpuAhWtT9XmdTft7fOCy6uLpSNpdgpnopULCZu
XFpxiRfmeFaqbQwoMEDYqv/IFgqfMrp0+Du4VEx+bQkHvS3tBoUdw5v/Qsx8jCa0WetQszBLLCgp
lpiQI7WkiVHzJBUHlEy1/6bkNm2Mu4dKmYgWT0edBY2WlGupm/lj4zo/S5+Qqi/AgLxDJZASRKnY
MwcIyCItUJM9bvEOJIgmllHRVyYVXUazqGyNhfKCLOLJNN/fKlfzo9p4ZLF6Ewq8aEAHP8GHHhXe
UMN/RNz6Sy0r6GcgRvU7OpAwDpLFavGpmsm54YwCLl+wCm6+FuI8o1OAoMe9a4fg0yc37JBUd5jI
et+ekA4rdh9Ok5ak7EiVQiMHQy1w7npwcXFGoWO1uQJAdZYI+Z9cIBRGR9ox73A3ik7JZ5UamIqH
NVm1wpb996JGHTLAdSnHIiSWVuZ7iy9djqyohDFHIx8IS4WpgSg5ME6Ux8X/oFTcH2aiL/VAR6Vv
qtQQs+0yBTR0OROixj43uSpWpGyFqJbJzRpCetc53eapqFFN9JkzA323nRWYMV4Fzr3SUYODoCVR
Gd26JoK12KIN9H/E8X4405lLTftqcPoIccWlBvenM9arQldDRoP0ueDp3x8xXbXldxkChg1slD5F
A4TGT+3UsQvNCOW5WEHGODxk85nKXpdsn0/mtBL6EzLM9FnuDc2Wm9DuOKCHAKry1c1OSKphKv1R
dJUxUH+EMxReCgMd0YAIN+Q2Y5ujZbI5vyt0zop8Ri+5ytkPiiDmp8FXPGzbatskGKhMZWpPcYfo
U4ZjaPB/XFl1o4cQ/MByFhXprmzSaGlfL+DXFxIf0R49K0gyVYywqCZzhwm2jhYWYwMxcY01W9KV
VtdtRY5sEfH9t+BSNriafsd1GbCb/41g+QO0MUOBjFIT2Kf7nQlmlT39o/JesQH9xGNYhReASAqd
XVpOF8UOJuHdZkDvc9RrkwfdJQwcY2Le2jSwK4s4oiNP2DvmBievB0BnOkwNdmLPsxHAemdRUZC4
JtmSOLmloolWAIwrvIFcgfcN+PfbgvksvTqvkzYFDIETf6JrKGkOYguEIKMdnLChWh6ng+4O68ow
Ji6OGBxPuqlLlnOKP4LelRB/PGLGvaLOfDxeHRLSG7HudUujNujG/LfAnOqBdYMmhIvwOfP3v+lp
YY0Y5bNz1EfyirGbvi3MWb5wIZYJgkyancPcezb51vAEtpc8cz7b/8cFTMIJoJmlXFxHcbUSXZHI
4AScznqsCHnK7jTwHcL1cG6Pr7QjIATn1L96bTyQVWLTUFUeVIfnOyno0sL2m1gqzKPGBRRsNnYp
R26XOSbpjC+e3p7LkQQ0NoGBnYgmyM3Z9Gyea7rxoRBzifcSc0OTKfMgyMfO6pE9XN1WlQBvFbJh
fiGaa88eld7ev5CxlZ5hT9wPnl3rlyRNEeeyDKHrfjSvhKc50ZMlq+VNgB/Zlfvf7uAQ5kxVm0Yp
VCSgaqLLiTbfcHGCTHzBoH5DwjzPWI6LCPfIv3ZbDtMyrLVpvxNzsSsVD0tSHvKQhmXWNhoMTtTL
Bt2CnDd3JogGn2Uu+vedB73ANrBKcdASu58/aao9GUlUVE/4spsYoIQIcce9WjBZGKzJ5U73dG3T
kk+YqHsDftzSlaaze6ADblzlCHzM8Do9NnC/6bvLGgCg+8h4mGgFyw9E1FSxbWEmmWPo8/7rzYti
uFQpJtMldij63OY55agVCacyd+7vsng0b9+aBEVU0w23O1tcbwnWhHi+QVUnzBl0MYq/MJzjh9KE
AE+71+yMVB0PsaofxyjFkejwT1qT7eHlZzZQcIJEcYDnzFG0aO0RsSPaQbUT9OnRUNVhDvHocHFs
mbTqIRubXLl9J9kWtYoV3YrJJqMZcQVMmwbJOkkpLFd9f3Xm2D3+P5Gfn8yraFesOoFfahpJm0G7
ZuFfajyd3F1/770CvnAngW9FIC8CWfMlSR01+Rv0UQFDRvAbnGk1T2zgENtH24GJzNjtmfcP+ugN
fCt+/H8D4hNpV9/aVWGCP+9bHM5DXiB4SsBdTk09ErxRyaMBDYm1owuZS85ibGtC3ar8f+c0zJ12
AtRTHgdzhKJPMp6vPIGsrozEsv4zrjEYyfuUXe4UeNJo1Cckb+Oew2gDL79O+9jgPxkStaH3Q67I
/zuxWPUjWeQyNbx0ZytlSiFVJJIqZzQ2ALLAD3E4ulx0FDDa8NqLRB/TMuxnuLcU6GpYUI76SeEv
Qx9LtrtJk6+Vh+zSr0mHrjGdQYg1AIs7+qOfQDOXSE2tTS7qOMCnsdbhqHq5bX51AXSHw88axhTr
EAEoLEtEc1MAk4m+WHiPRTyK8MSY2ab4SX9wUclozLh00ZwvCwXkIShbVtK92FLLj8xQhNRL4NLn
w8L8mNshFq5WKRSPKGxGCPsTWcLm73ND7FHu+miT2frEQc0S9XpMx1HDrbf12M9LittSNDmQ/veR
/iT3DS/BSMvLmiI1TnQc6lOvi1fCjQleLV/jBlU3XQqeOlmgw22Htd5gXZP7SAvPVh6DpnTIQkGl
VKYgJfmyhmpUPoBLCEoMT3VW7Fh1GqXHkNtVNEFy4eL+F7WSMp02X+dm5hPa1pjvWaSNtFl3uZhX
jAtaytfuamGxgcZ5OJVQgnwwd8Djiu7k81mWxYf+IFc+rjClQIWGajgiqTQw6QF7N137ZzbjQJbS
Kll11GB2ui37bUpNvOYTSnSpD1OTt9tXYX1cGjyAsnOVyiRkT62fpCIqmPUMAxy6Zi4LYizNTJ5/
3ovRS1ogerj05zenDV6JZCFhQ//1bA30fa3+A3w3LCz+JNT9ljwf+MAsOJ0G2UTlvs2tUnsHuSUg
z1/DN6zhC2N9hg/TkhAH2D/rMNTpLOMAjtMMT9p+2o2WrDEyuXSHxlxZ8m2i86IGaVzhCDrgF9ue
hFWr/EXT6BGC9pmiBaGgPIYCU0c3ZPj7gc7U2I/Ng5aGZAvH/alzokGuqBJmfVPFawXmTW6de/+z
1Vx9/kSZUq3qM9vhBG36E4kvfMnD7DUKSIAMhsmI/5c/ghnfeF8qzi6uE79qUdMwWnaV5E659GO4
u+NVchZKwXhInCREt6AiwZSa45XqN4BhKfaDGXam18HUfBzxD3T/oqtuvrXJ1uFWmUmNTn+egbRy
bZwW3FOxBdpYJOtV1BfO7XYPH0Bikv0iTvaQ7ycq3XCNZ181Vw6eMLba7yg6QtE+AHvKL3/TP+UO
dgCDeNEv93U9BaT2/SNJEyqwjA6Y3zVm7+TgywHxD8XynkMhAUT1eeua+/MppmjWf6s/dKjDzR8V
8tPR7cDsHaHxxSHk0BQlDo5hRu78Vl1Mt/QpJmI1bG2tuxh1UOzmr5xSfvagW5n8maTU6pMApOpa
VBJ/WC/8PLLkbFQjkkeMtNg0tPHMb0VUr46ouMZ1YMHOXc2HP+Yp6Ng/qCC7BAJBGnnwFhn0m3sz
GDMNB+uYQ4tOfpl873zKRXmu3o2ZBZuX2e05B+9SDcWfux8tpfdUDhrS7Jdhulb3RFymLHfp/Zdb
8N4KWBQoigXl8ey6ZnWdipV/VVN6NdpFqsEMUF7l9Qqersd8O5rSNbikLolN4bD/l1wlIngqZRJN
KOYmJD6IL3pmujA8kaV21uadwEzt1j6J8DxWhxvww/gyCCmf7Zn/UT5KZJ3gllZfAO4iSLmMLqQT
qUNanIn6IzHisu7DwkTnmlUnv9pSx0IYUJLIp2Q0c3di5wDLxlG8dODxUfOUj3et6LBA/m10fYxT
dNz1KlmDU4QejG4fXrVdBqNICZ5T22eQlHmWU6z4OGP267ynmMxvObA6JADKI7k0TeFJ8j162gkS
FnsH/7dMxCFq/Qd8o6PFjy29LF3STDdGMx4+wEREe4zGy+u/h4VG2dSsn/xJuxUcwyCimopmMppf
8p6WD2/FH/5S4R4s0mCrLw7/c+8k76vktyfw5n+T++W/LtXGJDVLjDJDlim5dPfxy+oA+hHzUem4
HnDHyCy95D/vkmOjPPYAxL+crcC6KxSpZBKq1C1bugayVKmICL80qx6AMU4cStSghljwjSOZGjdG
NmHZwD2HLnIsEakDjLTZZRHCMnAJS3wBzhtHF+4GLVOnj/3mhudbfdfitef7XgXrkZNOZkBEdmK6
EklyvzfdEr/yNO5zJOjMwXiDWLIQEal4kKrjXUg/zMVp/OxwezJGjIHJ/teUmYSzsRBcHxirrqn3
VB75laBBFKKRNqI9qhZ9ItF5W+WEr47/8iGIkpauDgT+peuY2KF6Lgt2adsBzbngLA66aT6NbJsb
TkWABG42ETyJzE0ujk0+0Fb5WWKtWKTgX2iA+iiDoZDztqQeZg3tPMTgXD4fycoCBsVBgYlbceVl
kmFpnWai2nxZ1pDpNYmBokMAS5EoTmQ6e3E76c/UfwJZCTwkTCQ2ucRV1rK2TASTnCnMCC5zHKSa
n4CeraGAZeZffyTq7n/aUbjOEalYu3OOqikLJblOwh251P8FvrqL1/r+g4hDhVGtk7qLNUHu1m2E
TPWUGZsIGELtoup2hmG83Yzr6Jk4A7+9AiyT7+V00M7lVPBImd+TUW1rS5cvGqJRvYXrW2Ef/eJn
QjdUczTMB3sW5Qhb5R/IDzyaE7U4oIuI/SB49FV6I3qP2a/5CwXwzfs81mwNy7s5zDuVPr/wpHh7
wVFe3eHvwDCYFJzvyCe6M+jB7MrImQil8y9ortX7GSvrv+XtpYYmrMFgLN22DLmy/DpKPMNcy9aa
kOn8dL8PCddAflUJ9Q+rP8mZKQt8Etpc3m99AwFEMuK5dDDlGdoC6HAuZORPs3d4u0Bhe7tEzX/O
NkBqHrbjbJ/siDaDk/czQFu+JGVn8Jwy5Bc5DxRM/P3/B+kT4azFj0oM0bF3TEwFuXJZRSUUieK3
nwlQOIhKV/8mhVqfnYUaaue7Nn98XV+MkrA0m36M5CM0CfMFO67fhBhP7jDG8qKicR1G6EEt5h1r
m6DPrJ8gEr2sC9vk/Tzj9p6GiG7H2kkhhY/Aff6O/9hn+EaKzBG04cb14erYRKKtnPunDYPVQLpD
Jj1l04dP23tKdj1ZpLB0F+w7p8c71BJblaevcL1ejvbl7zLfrw2m7dy+DlmOI7mk2bLrtJScaAK0
fbBSOgW0Kby2Oa/hde4Qk/xGZmLWwDs1jHQsd3aczovVszCwv9SMp9bz7gm1FtTeodYaBSpDxApa
JmQYu2PzTH4HEY3dC52QwROnvxeU+ejtOTlzgx6hZhQJ3gn3/ixvGC6TNcRNGZRkaahXR7Fj6jqT
gXzY8h+V+Dr2j+wG5I+zdpemuiysv+B1KwK0rxqtCZH8cRzKRzl22MnWV+GQw/1s7/5zxIibgoLg
sE57sUGehWNMIPZ2RC8efbIjNI1CULlNzCO3ZO3nVz2Bp9ebtZm0m7v7JiaikPtyDatFN3kXobAq
vLaN/uH3p8PR84NbsIH5Lw6kz8ObsnOLo3JHTkm2SjzsfwY5PrwbC7czEdLReu8cfxgqAmO0Q/jD
Xvay5ckrO0Izgodu6dkFy4PV3Tv0hEPHZFm3zvWgcc/oN0/4Hl5uRA+J+EVZfi7e5bVrmh7RYxui
6FBvloW5OsdgueXejjnRLirgNrGzZR05fQzqjoqjF9XnYIloSDEhCaOh1V1mDiBuzbUnPwMoe/3k
uPJRkmdhgjOmASK67Nuu5SQfN4alptlYhe2LDMKpdrMV6VLEEIyJpIa7uwpCqQnDu2J8tqtnYh5M
kfCu/mnnTNaq/JzCspziwqqHbb9tyIqkj6HGcz1TyNsYCpTFMNPeyfXdvbRBn7mMLhfjwpuPdsVg
W/cR8iJVicRbz1zMFaXQJ9nD7+uEoRze+0ctLX7xYxpvN9a8XCYgsL82Wc0WQY7CnMuVw6CvmVDX
x0PXoIW2V0EbrHLYPHogG70NJ7wM7wsVsdU2D832GeFFHln3Ivt9yxHKBB+2GM5JBwjPH5RF1Y8B
uUXyDH7ko4+oJEfU3y93yEUZ3gA88js/KItvPZEBH+YDwy6e6TEdJJNAw1bKkkuTDo3QEi0iYSec
3cymKIVz7FFhLYYz0RhadmdaTSVn3GQ0vjHpIiM5dyPeRuC2Ja/g/eBIgPP0eIFcU7FBLhWiFXaP
iW6LbCcjOawwCckCGq4Ostos/LExWyWRiSpT6R7hKWxLjPjq48mxiFOOQrY88eWdiqqAcZldqePM
Dl7p3huiSyLMp4Z+aB8Rkl7U1Q1+In6hOMIZ56v/LSORMFSBHjhUOzrhoQ8uH16uwVWcmptfzuh4
XLNnB+tf1aqUN3rZdGXzSgLt5Q5Se5mPeMxHdAp84kn1sCyXM1Co0vYhtvyDf/PHu/FXPB6Yr5Pg
mL/GZ/2nu1ngeP9RR9dAfir+aqA7rh+z+82MUkrcOKpzxRNpwK3VzvLV4mt7ZbpKleMvrRNYG5HH
WFw+K+SBH7nfN1kD3//+6CqY/3+UM8ylnKAh7AewQGAvx+CmZbXeFaPUhsJWGG0z375opotfkR1/
rnn5J57/y+93HW5pZGoa1s1BQ1sl0cjA8Xh7S6pG91vSQg+Wlg7Rf6cSCfYT3DYgPWgcPms96a6I
+ss+7n7U1t6f0hLR7KbZpUwsp5iH1PTZhGSupN0woxVsDVrmiptuadIan86hd6f4fu3FYI0S4kmE
/DWrGUbXpjn992bG1iRYoCqyLjGoms3+AZL4RLU9F9pciFJ+Q3qtuJ5s57x8AjG4few4pmNqDw27
/u5/rP3tox2vRwyz83KRGPW2URJSPXcW/pfTP5ZRpzoP6t1QghDc2JX4MOC1ijrfuayHQ6dtwkYo
WoeSFb6e4SsOR0vDHkkqQmJpiyrWEUxHBlYxnb1Zi/mbN6YnMoPJ0YG1x9sKtPjFn4FwR/TiGSlS
NNvQ/ONmfiFy4eJusjoPYE+OjFuNAIxYWa0UzXjUmfC8sxplmL8UB6k6j+r1ZRsgPr9nXIxN2i+6
AZ11KaCOcC1o/iXEh6sZeyS09tQYaAWnijFRVrcTKcUBC9RB7PH/vsX2vJ8U1RA1ss4k2hQMEjw/
gGVCN8rK/+XKZPswgzHKmBJK+sdD/JClFNKzqRlSpSWHJysco4KwAbwq8FtBrj5vahQQ3t6e2Vi6
nDhhqNPawzSGMDjoT2qNBwkLuZM0FRwR9+4bszn0x+ymebcaFTGNrgIF/BRo8XD8/W0C7IaZeJc4
3EmFPolXwW92ky1cdaqBZvjtzQcd1sfB0UPzxEtI8GO6z4o/wCsbxQE6XvrjQm0alw0Pqx0Wnygp
ro1NcSo36cccob0rhMRlKXa/v9HPCCwG2ik/SO+nXe/pOwgxu4WNG47GS5ZgshTpdOlRAKgC4VRz
bJ68kjO3Q0EImNcWjuzlQaDiF6L4DJfnGvgELi6rykxIMJku0JUkW8XNgBouKVJrgAej7DZsmj5S
atqYTgMRccl7Gn8Gu/ThSzm6/0lBhRg9YWwLJWrjnU09l2bHjo27U2upmiGgMUJFkUV0wl0Ztaxq
7EktFSZz4aqCKZgVX0H44JQLZEr0I1AcTh1N92vRVBDqRx0PYqoZXRury8Gjb45u73bWO/XyRo7r
DfZqu8x6XsICaqoIf2hHLKMuEdeVNSKajQ0EVnDopRxJ1iS7NDObFbtgw/g0JrpNe3P5hv0E3G0E
HnSjsf4bc1lJ2fRLGfOBTyzj74+J0G9GRH3GiiYwD78tyjiEmxbWDZ7tymevg2GJ3fMkBPdDtefz
v/M0dQvF69bnYz0A2z4gchHwYtqW19cgXnAqye1VfPrVLGJwy0Lc/C2Vc+MJJotcBXHi4jokXRzS
l8Enq33NSjJrt+udYplEvlWwa3PgCY9mHRdBsxCQPMJflYVpYgIVXZB34ZYVotgd8mrlE+49aqnR
DuJyL+r0vT2em9VBMW+b1sifx3+H3XREZT+ors5WEBuV/TWChjp82XJv9/Z0lyJ89nFxk0GRahJt
AR5td9QuX+nDjgH1WFxD8+a1juGxxNXHZmHEFwYgNgj4rvlyXMRuoLx6yPGP/xuZkofdHao0Z9mL
jbVp7DtPKuo21jBBWnZo11427ibgR0qkuOZxy/2Wxp8H3VgRrO+Oe4gyV6ipyUMTCtDXf70bBu9p
XoKGQcLZwfkqHoZLOVARysQuphTLh79gtAgeANnKPcbWv8ofJ/xBXfIb/cRmwBv4J2RDZCJEN9+O
6GLI96n4LnHfRnRtm8nr+e6eYf8b6TsuXRAUk1OXN0ZCt95iwd3H9puj1VXhOLoobPPU4MU37Ihu
xuGAeNgl8TTfRC2XKEb1WBzNWD/9kkqhsZKpb84PkV9SSYBnN/mO+/zHwcnr3yqOKZFtyyBxeWuf
qRRFXIIOrlZHxjeT7/MUllD6+HnDRw+BBpCxpP8DP48d+bxGVVpRhcQ/HFiF6dEdLAMoVBod/ojK
UyNcbRUen+YM/+oib0ad0zINV3KSQWec29YuUA17cTOdvcwh7SuSAhZyWBBCvIB9V+3PmEP95PtS
eZXrgHCllwTTLAHtdwO2AuReUL0kzMGY2zB+sx+4uEDVsINhFmLwlfzQ/TP4ZV9JBqSVXGNTCm+p
FPdRWMX6T4cFd6WGQMLv4dh/Zh9UYOnmuwKLOScaR00DgKqZTNKQ0Gy6AtFy/fGv6kF4Q0P5SSzW
MrDNw2/w4oGzb6c/KcxZ8q5L/fkaplw7meYrgnB9NcWxaNLhy/9jNU6KIM59wo4FFpXomIERCnCi
+4G0IpcRmwqXvpqTdd4llRdKcGn6v/pxVmYVFtfMSbTEZ2YsiNqGgWABcLxKKd6Gkoj+PEA9CKrV
hEF4vztgGT0sUZgqiTWvbv0fQ2Q68sVor7oTf+e6uVF6E0Qn6aB6eIOtTwrdPYl48c5rZwlhSRXY
REluFvNx5vP/2/50iNp2A6s/wd9ZCCoQUFZLFNYQTecPCZlY1K4V0vsOPxSp/df3fV8KxxXmKyUl
WhRB7QzHiFmqYLuUkiixHDRAPVKKWf7YppYu+4JfCCl7Xyngf3p4j9eiz7DgEIopTN2RaK57PfgW
TC4trF04buw8uMqF7+dFZYr7MXpYk0YAlDCXdY3PQ+jlQu5X3cKwmMl+g4W97LQVjioJz8RuAE7n
aoN9wEEpiY4ZuOob4WaBBxxRzlndXo7n7ylxiOcf0bEk2kjWhe7kRB9T80TUbf6Ps+TIDSZSXRQN
p0/tgwoPlodT04KSc5FAEOX5BbSyrIHGwSpP/9QysRDMaaqfW88b2XgjnX4TXhLGHY1RIokH5mK6
AZLVrJCIg+ZvW+JC2nwfZ6ioK5dMw+oh182ZpE2Lmu3d/c5Y+T6NM+4zUop6k8X4fPAg4uq+K7VV
c2E9+lSPmDAE6eAV3VqUY3tZFsHcKqJJh3Zr0YjrYLtZiVKrlnDTOkLMgPrH260h24gVKCkSkXoY
tfWTmnH5OINSeSecXLUnpbv+AFzuG/CXx+gNfeqN02+h2uWhkg4BaTDapXvnKVKk3ewwq1B5FBi+
3zvOCrasJNgL4FuiVW9dHolo434k17/zTBO1mNZqa3xSQSORtgw4AbWnq25lZCsQJrwLu4JIQ3GT
e3lLfO6Y/ZYrMzmj8jtfxq5s5yX1y2GtopxjN2d+1/LSQGHLrKOuzxuhiJr/z/fFbUfQNLXG3ZTB
C53i1UTJ/z8+01Bm0Ewh3XfXz/8iDoNHpR3Rwpl25iM3EsOsGuJv3duX8qUMNTUYF5lrVTjRQ+7n
c1czKsA1J7joRANt+MTEJ0j1Jq8/HSuZSAWLw/ywgggDXTL1B226WjNM0e4M8YDTziQrp09Z9GA+
VhKcV1Av+tHG05WptIE+J22chbrtohR1Uupti7FFBQNNTmWH1rcCqvY++e58iQBoAMlFso0SlXZv
DjfUTnapLlP4F1Ur6Vr4p/vlJ3lUlci3KLYmM8W64F8aPq78ZHOtJvqiJdJZcQUk/m+tFpHxeqIc
7F6YnXUB3ILs8/YxOOgzYTt3Wl7Y4vZHP4Y/muReETZH6RRFeXZxYQ42PYeQl4+kh/4C9wSznuzs
ExIZ1qzD8Boyv8hLBJKnVfbr/+9BoiXePtycWBzPtT2yveCLjUwlJiy+B1fWxRjILOqUf+mcbK5f
SOIhq3ESn0dkjFsM0D1nawMNt4xu+2EHmkM5r9NYfwhOxYUUyBcL/nSYw9DQPkGtgKUquKM09dMV
Ro5Qtp71hean+KVODNtryq70wKSGdd1dahoMByQClZkwDyeMCGXDCcmakLcsyQWFHofxBQ4zPPai
aiZ4hU2sG8CtgZraXsmhm+a092ECbghVXDz1SPFt2+V9Fk9/bvQJ44zrupRVJ+8mbgQC38jfGvSn
YnfKdLj6pfR8aIrxBmo1UP2Z/WB6dRm2rKm+25IT8MthqRzuvR3s3YrGMSUclL00+pdTfoSkePH4
Yq35FZ0u4tpSz9A/K52A4BHf02YCr+3VQqOHRO2/ysy6KwbxddxRS8aBwbqY8OWisFpPGMP7mTAA
hTkiUbDGkVvyJAO7XAJc8qo7eq2K9RxXUfW945xletQdPQod0+DBLycVLBb+HrfLEzFz1rR6X8NI
EDYaBT5JzyNNdvFhj7w82vGVvJbIEuNHBa09SQ8QvStk4Hr9dcTVd2gszAp//rFE5YFlGJON2NwK
uXy7iWIPksbrL3sg/6u6fRvuyjczz4wj8J9m17uIiln8sn0mIP8jBejRE9mz+SpRelwVYO0nhKKy
wfX/MNEm3ZNMd5Ky+ts0ODOj5xaWNPT9xgDuRiXG5tPi4/enOrPz9W076Fa6FdC2NrlQ2N2lLXmJ
Qd9jLhn4gbTOWOMjmubE8L7hkGTBvh8ALsBLs/xAC31k4SRndTmxfZkjxyh5NTgjUbP007RLFESw
qtx+CZJxYTq/lemdCaIXGvPBga9NhQDqxV3AmxuhhCA8Vn6BkjMSrrayPNApThsOmxjd5KMOz6Gk
2lHubaq6gROyVrKtK/ZzCYQNPrL89u89KTBI9KHdZu2LnOUygBOK83UReMBTtEz03hsO8zRt7z8s
HpZbbkgMeUeyhxRgUoi+5bHIUbRxI7cPGa+Keq4cmf4vwk9fgp+W5lBPH2iQmCzkHtClibO9RTMZ
FMLtHWyns6nVVi2jG3iXFeogg1vpgLQrWYA1NzyTE+Eq9+ecIphafh7cr8JXSo/Lkg8Hx9Wziy6p
eKYSwGFtbT8U1S0J8lMF5MGHC/cX+hxVQAMh49nbrX0GmHNeloV1w7+BpMkUjWzjA9z0JkyrNXpR
MDBigChf2Y6EEFAft7wDtIwZNqJEJlgKSUpyGeOmRGOugs3cvqazPgxfq6MVjjXt7RQCmhGnj5hX
KSADYsSxxEDvNLMWCtuImETiipESb6gdBCLMfwRoUCfb5Dqz1wORrmz2FR9QuybC9/Q4gimAVfdE
wAIRzXB4DuWbj78tLVr+OHHMCLgY8vCLljdjnE5WxxPhDvOuSL0L8zlPftl9Czme3CfqilNjMg2P
x5LPpEMdP7wKg+MOY0GqFcT+SkPwS+j/3hma6kBGAkLKtn2GsR9ah/i4IDeUCSgIuj8Vz+64H9w0
8lgFug2ydH+Ja7FK2IOx+LRjlL7Vkx4t7WN5b6awqyEYHioveHmMPqAHaLd9xUbaOAUH5cPMebJm
3Onz9xwbSoOOSqig7vyUOfTa8woyTufd9TD5hsmgV2srwUIJgPe182DAoNQTeEcg9mOX3sD12kGn
PhJu1yrUyu5lc35irrgYcbtQqQZsiEniH2q51zR1uggM0Wltw6yk3QDSlml0+uRwe3AV0SIEcnYs
IlYqA66/jjfxe7j+/PBREeGwIE+UkNCvqnqbXi6a8pjMvoxojdH0VTmxTP/S9b5QMksuEo4+hUqa
0RHw5RyuPK9Zncp3sRyTkYGssKAE/CfVt1+4xtckKHfZov4EDDvrnENTWZ2JLamI20eRleNJqZiq
RezRAI57QCdiYFR7UGAr+zBQi1DqkRMD8nT5d+44zdzrXi4BuNu+k9cm+8b6g4ZfwG2WaHn2dWSS
Ovm4748nH5TddjcRmWBJVjG1coNudkiaekSnesQeskaYHeyttI+mXvTC4qbreF1jXgxlNSp1gKNZ
awqBLRc2Mr9kH1GP5AAt2eWbEHtWVS5lEVTy4at/vw0AZMykFK/dE3kM6+ArfmB09TJ4aNlCxgFB
SwColNRIqL8DC4QiE+a9b6q48vxw6m2O/yAdPdoZp1IyH1hE7n6rpqn4RilEGNoS/NeiMoeMsDSe
2y+FAfmRaHC70/tNfA/nZrFcU2eHoQAvKAKKrD6+bgzB98n+4cu5b04pPv8XitolHLV0Unpgu4jh
fubVXG0y3HTDbanTZJV9eQsY3DLGUaAFbS6PMqySqt+KvJ2Fhm8uu35WZN+/BriiBCNnMDhCBVYV
KU4G1UgU89fMhD4njXrGY3ImCyjOBZ3605czbaPvN7DHNGXJq+9KWCzXR+kvj751/WQXhxuDmG6l
UQ8+zwKxJ3SunSan9IaFSWAJWWjZRkJX4NIkLvKUXSf+MoWbbYsPzBgu/da42wI632o3RR2wlSuK
qMowAgudU5M7q2dSnnhRf1xjevFVwYoLH2jzlZc/U5dfdDkhUOnchq7b1Hi8QWRb8FGC+023DTS3
OV3YKUUPKE8uuybCqjXeyqDP/1sJDINsvJIBQ/QIGL+VfS5V0xUuc4Ad9Ux3zxztNEPX3RO/ZzfJ
imSsOmJ0CuTyUdfYx6eEoKpQrs+lwQm/sRSm0YPcp5H2g+54+OLA8XevFZf/rNfYMVsVEnqdZnZL
eXtRznzkLJFeXf1br5U82OI2GUhrbb/HT01kW0dStvdOBPD2TV0bA6y7kEpNV/x2no5kKQWmNFkU
fZpROx0isdOCZzAqTxkyxFouztZYyXZi7LMpW7Rma0hrBV+/J/ahu1+DxdSiwxUUPtSm+Kl2vhid
lC+p4FtKGReXmv+xugbM8WXSEI0hMYijnFunjCwVVuc2vI4J8/xHayr0xcjKMQiAGQz+7drgvj33
OhNPskV3EwRMHfGMEHO3ZTX8jRi+VsbwawDS9eycioOF7BkXEm2tdHt9azV2mY6MWvoFeC0Aaczh
3CLMDbMPUZ8Y+1SliiEfuTe6XuInIDQ21vQ6nLIcKUCwph9RNo2bIdxsTqxpnUWTxwY7+P8k6wUK
gzb9BPWL+zWdvyhVVu5UxJe3sNxl5cdg6/Q1yCIfHvxqJBMiTdlGf67aza/gWDEb4BHkP2F3QewT
P7Jc6unhcomOQyp+TmNainB/NvxIWwCLtdw97OHfldVHyOSwSDd4pV+3QHNXWvGB4ORO6sZmVcNc
kfjwCtFgIkJbDGxUboNqxJChvfj1C+iSQi1+NP5HtzIgzIFJast26Rt7IzTZAOkPGxGuF7zpVz2Y
iQpHlOc/P8XXGG/cxvunTIqY8Za9hJFloXnEqoI67f6C9Qx4x4JFein8sN4lGnJNHMg8+TmhCzGq
QJP2RYq0IBYFPUUAeMIz1pygeQtLS1VkCu6OaLJdQgGssxmMh2MOmcPLpLSoIHb2nxjL33/n9lp9
elSSYZcnpDBg83GuEhG/BvX/2kD0bArLpcByS6/uvRd3ajALonobN/w5/ir0GUe9LOlO4KdHX8Ne
hbDtlmVAooH0cfPewjJuZIFn156/w2gn1+ToB6jhBrUSxRHM143Sswl063J5w7ar4qvmo4gBQt5R
age7oETATdvFKxU5c1LukgaUum4OqPSTVj88SPPTCbfsOYKUh28eZacN3E5sJscTbpJ9g+t4e/U1
35D4IwrBCdI3b4pDeIfh0KluKKJiJr8dcpkDfcmZSgu/qIu+r7SUuOjNK0ofNILLVCYisH6BqfZC
YqXqcoFJG4ToCeypateBmWMchsFGQMDMOuRXqcRo4Wp88WyneoTzSXFDbyXyZW0NrJ7SOVuAWM7X
PJOvrwGnfog62IF2kJ+SMSjBt1Icv2BktbI70txGqLzZy6hTiIdcKQQHrtAkq4PaLgtwN+2efMjv
jvVQn6+Mdytmm65wDibNjwNrpqSvYldu//8GCNm5clVCsAD+6c4D6ayA5+OxYwUWxARTboXyaVOF
UdjfqCz0AFO7bDVLbU4/3QqJZBspIbB0891jvdTdIpEyzKSEC/6BK/AYs8aSq5YG8nFdOmAaLbKc
Gcd7z+5eJvFBiOatfW2H/YBfCzzIb7jTgNSSBpR/tGImLEf+UD2ayjYsUA69ocCCmnRQLMo7D2dD
6IYgIsaej2BW8v4+7bAXAHluC2EfbmUtKE9l1/4G+f7eqiDiRkh2uTG6lnJUB1H6jIJ7JjuP1lAB
8Y0llcofbWv2klyhjeQOiagzfvC/3ocbuxOB7m8l7Eu7kX+S9BNqQpEPugarLaRDxDLwr0zVUvyS
DjNjinoJg2j7tgtkGwJSrLYT6S/3XZNB3IUQ4dnwT9mZEUK5Pdno/GTcKe9ut3HV9pEkiPBSK4jM
6TcmBx2EL3w4nbGHJzuFWtWToisTaDEO95ZsNf1kKbcMywVrTCHEwjrV7ozHG4ftRhHz9hRTsLya
vvZ21P9TYxlL9XUKAJO0DGRtSB2K/HrVsnpOWcmLzxe7yksEXvG4KbKTGMyMqMdE5Dz3LxxyAPsf
Pc32oDZXHYH9tjoY91PBnVWuuAcCuUCQFQrKIumSFt8H9/m40nmTtwNekRAzyVUS1noURb12kYIJ
W9CfO1KFFF6yLm5y/OqlHb+bY/MZ1OIq69Zmgbr7O8gX0qZhc+wpdHHSwB96Pj3FvfugzJbSx8/u
hpOVOA6QCtAiXakpKNZoe7EzjEBhcTNmRIZnycx+cItR3fdnsbMaYHjPIufBX2EwdOED/BTgMiIN
RCyuIPwmOndT/vNubSiUxfvZs2IRm6AD37MsQDLxjrNs3MZULAnBtm+gLQ+cbPUbRzrAdXwEI1KD
VZwrkmSm42r2MNdjKKXzopjlRLCh+hvQDetUj5W7SC4abHB2Vs6ShB+9n1Lv2eNv/D1sLgv3D+lE
D64qePpXM9dk8oxeYTK0/W2eiqUZcrQkM0N01nphey+NTR+dwQ+eiv1KDsG4xzTeaHSnYmW76D8H
MTR0rM5XfTsB7aNKlRmZOru6n06IcWtuKaWFm2pCtUnnoyj51Fubx1S9OTMAYvcrFto2sd7vgmlX
haDYEbCwwOTqHyZzgQRCBRVlZT8UTCQ2BvdkqPCKKEPRhK7uma+kRubUY+HLDCfXf/adZh+njOlo
302vEvPzom3cQEhUFJjv2k3+9zBM8a+hhJOrfNIaldAQGv2kUWOyRQfEDwrt+B/N4qQBepznpYY9
g4+h7xScMWPmrfdXyNhwbPNr/kaYWevw6NwOxqg5A6+CBQizHgiVONjikL9g+5LPBdMBPIHD2QcF
rYTpTFcVYsfJ0r2Oozb9Ru4R20WQvmo+jQ36Gp2d8M1rNKZE+RsqjnNS0wdt6lY3T77ZBIHcqLOA
6XTaqcDr3jJoGwKZucz5siPYhIpyrJdzFAvooAlhVhKHoRe9gNRFp12jBLMGrkkwYWOmybYEtcRH
9P35rOzen2BrPOlMEfLakbL5BG06dFK3+FommK+Axl5sosnxEU2BTc3VPGYT1dRK/tCJ12Cct/ce
gxoicubU6tyL2KaNulFko1pADH9R59PSFnIONdylImmUO7ldhuuVYxYB4vpP1pyekQhuB/stz3EZ
tC+nvLNsgb+GcsM66WZrw2wAL2hXuRxKQKUZeenUmIy6CS+B+Ay4lT0vWQ2BynwKKb3nI8kXBJbf
Gn4CXz1pO+E6CI8jnsFX3boaEzv6bjVut2imAUv5hMD1AtdM8OjnlFdQ//0phO/mw/1kxbIbdSJd
HQVjmbdin0GDWmozPGD1VomG9n0E5Wp1AhSNJ5xz01mNzMiNEBfl1IITDhC5EsZVKWXo3qZZOx5S
aVD5E5NLs1lKr6QEkJQmbaA89usTjw9zKVTssjmN3o8pR8el8qZx+4c1SKUv3aRpGTVuJDfcfS7d
1VSmshqcdNw/B0D/ufL6rmpAIcUY75NbIxCRXc6xt9cs/pGqxdZ6ZcH4X6u752d/I+csBgTWzs6x
tr/MZdNxyYwSobAIjjTpGwT7jRG2nafd1tC75yrYOFhOcaMoyRs3gTnLgo0+O0dYGTZ+h1dWplFq
j8tCIX2tmHxMjxxSWHJVIOX+V2I0fsb43iethrnRN3dk5J8VyPyFO5LPGgmlVVTdtn/DOV5Bg22g
fe9DjWTMOdNVjnpzAPslrMCuvAm0K6jezIrdAteFZez2P/cTDHiO7HyAKMFNjLRBLBNLZOHRmocE
DKs6NugAm+pEIrplYCSCvjSGOoWcYkqnZe2j3Z5oK1f3d06d42KgDpyeywZbDskM+TSkKyDEu5Zl
M7nVasjeV1HxoLEHi8p3NnDGOJb62TdGU40FvmYOVAvtHR3lkE/xp16QXJS+HLxv9cx/lwU9FHHN
7Im/4WlIhpD7x8ji2d/naohehjaMWZsP1IyTxmp1agYj0pNXBj0wD3JlzDAz6bSPPzdT64BmL/g9
wnUMXvUiUeVjtdlzDmkg5MNebmeG61gttgvZ7aNsxJp6vXN6nW7GFUu7+a4FZ1e4YaIk2UO1UzJ7
f5+PoXWLDUe1GsSgshDKcJWpXtlxI0zmOC/K7c3XLoRphOT+1MXUkclB1afmO+ealpO1l7FMkiTp
1okWBEydAGIQkUImkeMy7dH/t63ze1EuNYkiX2TDS9rkYkuEQn3RbX1L4A5Ki4Bzc6+fLsxgh00n
2vzYKXGWwXLnlI25ARrsmwJIOvCpaQLuQPFssDZKL+NVg6MlDr9/MjeBW90p9eVsBQ1xgwLcAVAV
dVcu7EL8hI8RKjrzTr2u1vVVLJfoJZ7ufENZoci7dbXPlPdjKbdG9AjFPswkFPKbP5x47LUMgJ/h
Vga+FmF+VLinuwnCi6GuzJO3do47ygRb057fAuO5Q1j2Tr7nSwiSBhX+WDtsEO6yAjCUI4kvDu4X
F4239mAl+Nzv3mzNDA4Ol6bM9GwqnpH0lJFmcs/D2ofGT/LZsLTtmA7KR4yHOLY+Z8yWalozr+Gj
HD95hLm9tGDUhv6Yuh0Xl6wjeNFV33xeUdtXMYOQ/jUa1bKUqKcQz4yr6XgW8zMGtXlKxgY1Zc6U
ng3bg6EAsL9vb/k43bxuhl+yqkULrZliUU4HxGrzgzlBRAlHAofl4lu90uEazME5E+PuyhywWUAZ
ib85AUWMx3mSxyltuwoJZ1gawI3/PIffy+O+77BI55x8tOl3E4bwVzwLZgm8bv621UVKMTrXxW7y
kB/IfowdPZRypz8U6Z2Flmm5/qe3s6E6EEX1X17yQIQGEKoR4uyrUofFqnAvyeWBfyhG5Q3wW9Q9
0XiKenwt/KT9ynr7ogtmBNhukYHlCGHyWmbVQCXkguzrwuMpFso0ugNfTCasqiGGu1IPWv2CHqBu
axGrrGn3LzlFxUyd3aDLYNidyfq1NKvoH7v83P/P67P7v6lmQfVWmKTT4g5RdG+XuCF0JwedT3Dh
sTsfpzA300I99q12U0hQXAvHX83szb/murxw1HwvGfjrZKBQUnFPL5AV+l4PcsAxRK2z9Ff77eKU
ge1WIcRspCobpBphgmYIgJYXj9JePK8NhJ9VRl6Uc1qYLQx0Fz6gGTlFu2d55lonfSs0c2Zt/8NY
Ut/UU6LWlGwzFTflKavafQ+EJqXMdIL4asKi/IEngY5CdGBxaDxi3QuHT7PYszQi9oy5mi60+abB
XWEMSgeT4hToNj5RXH9I2gwdtrSBa5tUvTxB4+z+Zw9yfGUwyaN+6r5Ee+JJl0tcn3Kj4pjLvm2V
il/JUl6jV+mLc/5yX2ViNBvKpZxskyAe3B1XfSo86Q7G/V8hI3FF6Zsbm0POnicvPqJNEKyHKccr
NYqhq8mfJ5POfJ1W6Wdjt0GzyP2gFVN778Oavx7zVbnqWf60aCxJwl4EFDi9Lbonu9OgE0OkLabO
g9sT8cUXxRr8871kBeN99Msasc4PG2DCzr6BH3WWMsy0IfxYXF2C0AfY0f89MxMPAezVkDiMG//b
EJskf+wsveThMS27QPnSQrBmJFO2wvf+8FmJhnDMdzoN6tiAejfxoofG4EDClKiArJJxSqjYzb5k
z6nlXTW11iFzd4zSQpMFr2ERH//7YpAz2ipqls6G1mb3LtHJ3ygT2tzhG+c9D9aBBTC203/XQkyS
lHMQtvNhmLPdo+1fknm7hlmUiRQu3Oc2weu3/xIxGKGd6shg7VfUxaoU58INJoFHfGah7cQcA6sA
Ts5ZdKx6zqfTE7WMUzKs+CxBCUPIa12Ur+jNRli9A83cN8QeZFkUFSf4FwOyUBsJc+1X+cK7EtO7
cHTqCRQTjDKvs6t5+ZPNrkwnAU4Uq5lfrq5QJ7NIlXXMP3cvXf1zgc8H+GtX8jhzS15Eqvh+97gU
yoHsAqqAFGAK31ldi1p4gLufKm0Ka0Vc14ZdIAaoOvOfPx6ddwOMuUUyR6TfBGpVJjCYnVugmatz
hlBbGLhbaMmltXoRMS68UqbSSbrpyzVy2mhdTjqDsjMl5dvYDWn3bx0sAm66gJqXQ4i+5FXs7cbF
iZTifuSoOgPZTPeo16MuHRGs+HDG+BAH7AK1SZTvl9sZoMNf2VGVyOTrqpB13PPupyh40Na9naIR
p2vyzenRLPDqB1rIR3c+na3ldqHXpjoX+v5OPPUSOJPyZQvU14EkuRsBiHqA9tQS+UyagCp9Y77j
xnrU2VBX0JZ+cUh/u4oAriPMyRJAf6JF3Lf4b91It55E1lGx2iNzbmLqFyn28jKlYBIKwcvqMzuX
FnCvCJuEoP7K4+76kEinE8fUfQO0067nctNK+/4fO4KO2ouyjRjeL1Mz9hbKfmvxY+e59JqfElPW
cQ1zJwTqr7GDguOD0rCakz7AlQXwP56jRefbcjykHTL3ctsZUTV+K4Xrtony3OdrcpKfFlEl/iKS
Ta1fTSah+hXfVn9xrdTTcmmlE6bXRON3jVqROAEP7xumQk2eB65erMLymBY4ol/mFtDuJIZ2Ncx/
BfI2+MXnKY1zZbPDoftljAPX1V2V9raeRb5+FGpYEObJIo4KDDX+5Kx3r4Iqw3wCIlcV6bfdNqfK
atZlygwFyZ/qvxAK0qMHtiNZytyQc2j4OQ+nRsmrfmjVequhATe3eTqvloZD07LmmczdNMyBL+TT
+A+sDEgAkNlknWXINanjiWByo+KZwvUUyclaVjGby2OZEBLWoma+ba9eXBeB5Lq/7W4FYM2u2bEl
Hf+Z9J0Ymad1F2o3PJCok/Z8tQCCok4sTy+kBlTIG0FatrIQWwzph5bWaed8cs5JX8RW90Nkwh2w
BWE+QIk2UlId/A0R+I2CXiUk/+mBZZJnLkUhMjmaQo8Epq1yqd2Vi1OEv3C3jCgmG4F99jYobQ17
MpM+5ow0lC/tnulm2L3LrytEnjLs3Sh9nQmFF8xNKH0zB7cRzjLr4x/YRqpakSnXhujNEpOJ3RcO
ogUFS2wlTYLjDa11haOeflRX44xZhBKLKrAc0cS79ui0KJxCF0ota4+pM3a5XdHTh2tvSstEJ9wL
pSmsv3TtTn1K7lb9dhZCXUZ6kfkLAWmI3vmgd7fPeNkKXrirBG3IZDoAKF9pYdFgCZhKbLfxJ0Uf
taPi2PCNUNqhcdGMMDCZhYX9P2h5bO+CnA1bRhAUe96pJ6GGEdyLBHiDZq63dzi+H/SH6ynSQtzm
VPg2zHwQCnbehQmsUgGJ8QJj/DQEuZB+HzO+NCXSXcCD43JZsnTIyQlo2FydrjTCFdpx5A20r4sW
hwCcVF4AUVFFFKyURK7tLaQrg796EpyQvsmLmQ5/dzJEkCIo6FbA87/5S7NYRXSgW/wwZR9SBNo2
tTlIDUI4KQeFY99OIvtDfVy5yBvy82EM6A68Uc5l4ODOuxy+3DUFIQszLgFFIO7D4iNe5pYgItZq
SxRC8iR2dua8OksyYZ1ljFC9vvvKtbUGfyahOMf06aN8yij45xUyF+rNAizAzWG2iyVxkxyq5lDZ
+RH+C5r1XMIx8oHzB057kL5G4PVep11+6DbFEMdaRaDaeE6IS8cU27QX0MjuAjX98V1iyJjAM7E8
6/30Vavp30jqt++Hz4fGDv2u4M3rzooX6Bxai9JQ41gtiK+q9FaZgbu+ANh6EEiRBBHYooqiHDap
YTRYVQ8fwdIKt8nxtxze4QgzUdTo1eg1iSmHIZ+AdJ7mKJ/h7vf+xpbzTpQ68V+IXb64/RUZAjuP
AzhGgX82In9QoZrQWfSMRml8eZ0Ua4dOC+KGjUBkS+Rwy73SqqrHPH0S4X+k3Pzj1/VFpxm70dBb
uFVFbqDGoQkwKmcYECgVdf4uOgO55s3iWZnrkkopp70J1XTwi1uEhRVtqUce08Oack0eUg8jImPk
l2dlAH1X8Gkl+9lCUdA9CFHWsaZaEWU0iSnG9ztPD/SSboaiih//Him1dpjiPIZaT10jKlmiXVE6
4sWd3BRba0X3nhJObc8RDsL47U7koQ7UNRJsOe4Rb67XCz3esePu41hv8ceSkaee23k3Uqr5uSoB
VZ/Lp5oL+ItSkQrwFEN8QOKLj0RYPhd1raSMCyORPTTRn5L5gvrr1Cx6joBl2OPtnQ62Mn3H0Rf0
235yiTTrItsrGdvNBaQ5jF0YcbeeTDERwnk87c17cx/H5VD1F5ewUsMPs/cyvcvqdLrw6AQSjced
TfEvRa3BhFHN5N54yrOB90zpB3MhJVQPfKbSk0Co41/Sm/pjhz0XPZt7eV6ExfywyhCfp/yHKHRC
Jn3QVx+Aw4Y5iyRNdwfKWds3kM1xqc5eKu42ZgBtKCSkl0Dlwy48Asc8F/fNx7YQptQ3YKmT+Htn
IXYZfNdpyL+Ovx446EqxUHraVKMCMczTvcfQcRPKggVxH/WS+l+t6Nd7Qp+ZUo2yCECxl/vMGzeE
Co79wOmOy2c04rzV6iJeHXE5NKjIBbYRzxeRBvrZImpwWxZ05Ixq3A3eEXUC2SwudvGD1buOOIdI
JTKalcVg8DJwb4pBRo4bn5NQC0f1gQkdLAtxaVop/6jVMlag2EYTegr+1hgrw5jX/ISV90ENFhT4
zex5kyJo65Cos2oCXhmbj9OaUYEt1SuuSIgWx8L8hYFf0J1sdTrVHaNRY/1Xzhpzevo2zvCjaOvu
qxgVjARhoPQI7Gq43p+vY8jTX9GvAXk3T7g0owHL1o+GUQN5nyeQHHJyFIlLTt2LnC2mPZC1t71S
yPAzH4ERCTAg6aIN069h8tinTXUNTXj1aNvVZT1JzXpAfNaGEYRSJCT73cuVz+wFwhvOFcS2Mjzi
g1a9nc3rubUhBX40GmVf+rt+r7JaqvCBBKNbHPg37QDxvuTOtitIUa4sF/1cYlhz6t0o9QJq9uua
P6OB9SG00s7lVtCBl8TbErtKL6wK9bs/uEtOW2itZdFISgFc7PsXFw2bockGfV+Wwu06rBshGZJe
lxs+RgSR12FSEeVpSSogaqUXjURcepHAORXYXX+vwAdHVI75AK3pkAEX3lQHVsAJG4an9SMxdGQW
WPR9Lh/QMpKj3WCvj4ccYxK0fFxJRG/qrshWLMHrNOJtEiLa+nfwC6V7xXPEmbll6CUb3JBgLGLu
ZuF5r9Jd8a3Q/7r2HgnCJuaysVnNVY8ISjjTbN0rsPiTAb8PCjy0BzRpjp8v3yhba7f85mfxvXTK
JuH20ZTUUHC6X4+ljr4FDAnwmA2lP2chMHKm30AHl9tHLrJmzKzKF7aXcjnZi/L4vTKBMt+5fxQZ
AAvcsmaXbUulmOYy4zNB/yd8KtxbmaCcZdwvN1M0gwlG7Wf4ropR3mzNSPOSvKNJ2tKGgwE2JXWx
8d1fHx4c/BL0j37axIwTPVgcs4hHm2qjy+t6KdEKRETN+arnF5VN4TaLVh+Mk7D2cHz0ai908P85
XvdBiB33ynhZXcocv9E7cPRJHVs1qCWdJVXnMUk5MkvhkNZTN0nG1QmY/dzsgXi/wlLf9YuMIDur
YOceUqK6o4GI/mNurc7d+yaEKYod8BfvNHpJ0MtdNNPO0shoflzIV1V+eqTBA8tOjl6QaQrZRkFF
OjN5KFvQRMVQz1ZA/EI1rzhnggALYERGRiQaXdM8priI6UJZoyHPhyceIcHKYmS3TRBp0QORVs0B
z9i7HeZok+DLjGPQc9oPwI2F7zW+gCES1tY72FBsWnbikN3DXh2RTPC96fQBPtD7BG60OGxLzIbF
ZmCDFazoSyscuUYUb61U8DWuFNN7Soka4Yy8rM5Qoa+GpC5Gh7utqNAW9mSsFbiiPbwzE/7LwjnH
rOmyAy1tqluR8Tu8u4UOeVlQ8H5jEhLwfAkBdE9zkytmZUVlumJZtPd7yn1mvkQRo9Jov64QitJL
vSnJsdXhoam5aaS3DNYxlK7D35P2tczoPMVkg62MXiVVkUfcdUn0w/LKLypiAuNG5dYylYj/+MOK
KnHWMq96QgG10kGobw5mjidxMTgK+KOoyPwau5BnS2OY/ccWznwuj2bmSRzYxTkRIsFt+zIWIMz2
bMG4AaiXUMpoDCvfXUfYXJv7bK8tkgas0PQiPTG8USGhkm+ZyxIvsRRE/ItBZ7/gFtpL9bzGdtMn
pPGgPc97D1gFJuwIG5e6IWN0u3yVcQcEwaGzUOx3WBTvNCtj+Op1evL3x2xwhZr+2a7oRCW1HTbS
Omgq98KU/bQD2XniaIeJXDcijsZvQbz6pAw4w+jYacV+pVMa18S8i+XW17JoH6wPStaP1G8rd2pu
fPz2NtD1phEw9WQhXO7p9wMXoW1SA7cFZZQVJE/gFc5Fjn4L0F+YRBXAeeuASIfdoIfQfIC88Umf
CEzOiAXKRDs6Rn3DeDbCzP/Mj/8If/J7Wf+r9L2LY2rScpO77xyKymfutMDsjcDL3JQLplFB0Nbi
oFLJJyliyC2j/h9aRSPuBs1rCHZH70e8r97B64c2iBlQSOssEFx8MGy+y52ErqNfHBUhOgGcj7Ny
DYQtT9e5n5+dfpGK/xaewbopwpk7MYrhWpkX4SneFJvvE4xvd2FNKyTV5sSRV0oN1J1nkYigOBjB
YRvlgP/s8QSXfrUzbuk08f/EcmXDIlAbozmu5xN9q1EesxpJSCDyPExOg34BKgDgkK5GNBMSFa/X
HnJxMKGS5qJITPLZQTRsZ4YpwHUhv8vN04NceOlWwcPw9Ks/qIeizigj8x4sUnPxYmiYfBLNYW+W
wfDF4L50BDdyqVHt9YqIe/wWPd3B6RUgEXaK6nDGMMtvNf0m3phybdOfXhE8mJYD1glZ4eBEG8Ti
h4Wyal9VSB2CXwtn1x36WJTgUl0tuQlp7rvlKZwzJtMr2+62EV2NQPf0hQat6JNRn5PaCqkHRTzY
TWhCzrNG2Hoh3kPtykbtA+SNSAZYxMTAyfswxLy/kYm2fnk+TCkVrsoHB3ZSTQoHgeVK/X9ZiUq2
Jk0LtXjDo+yFXJWBdkpsX0JqDTER0a51yxg7QF3809ZxX7uBBteF5EOS3AgEJBGETCwnH3Qa5V5U
lRjwlgIkS9JHKHzKZZJUxFvi7rwgvxW9SRWqoUIwVwfE5qZMy3F+EnGkgD/42jzyhL63v4N9oIQi
GgU4GoRKkShedLKxZdUbLk5WwlkjNW+Nt3X4nO0XEMxLLNDvw9PhL4LvT6t7vkwLkoDlvjalv7XQ
LbbfCz0D6EX5/imZ9tsz7Q3vX4LK8hxJ2JAoQctooqPZJqlrVPEnZnMyoozAzCocX0mlQTl6Knhf
Y/Tduh+moNWC0RT+AEvZ4AM0rymVou91CN8VuoUOs5kY5eGFhPMaRdiirvxtRguV4aKCMMuqLcr9
Lg1t0rOD//H7uVA9MdODFz3cXvq3DVAhznYTOasHoeu70313mPIOI8SbUunp7Vk6eV+C/7XASztK
SPDXvwae5GUNkGKGELBAn3RCqwFmbLP4Q88TmIn1qdNowDaTWRSJWaby8aF/5cC47R7FvOC++2as
0ZnGS81NDA3Nr/zQewOKqSTek9KPrzbmzjf86v0+2uKHEwG+7yh/llRvEdJWqf0w7RZyHrGi7Ccm
BHo8ZhR97I1zLn9LE8rifjgzIDg42UKjl3z4o1+RnTX7/bPiTJN8ZjabnIDsFt4jotf1aLeV4lMa
mbCDybeDutkmvElztUkp03HlWKJog0yF1+HApKitfRYT7iIsoA1jk5++oi37U07cmOPQJmTZn+0y
y+BGD0aybUHnyRyrr8MnHxSYwZhS7TG0iVfbYDlIUj0cokajJLDqyRbHbHjwOoqhi2s+Bwgl1Xxt
dkJaPtC4MkUP/IK7psnFIMF8fmjJMIF4zF9jLZotNBnqZg7ugrHHSwYkmvfBh3y5sY15t0jTTG1Z
7IoSMDSgmWrOCESQVg5ggvVAk+cMfJ28Jedl4xb+eWCax1GR7P5qQtrSpkqgWfQu6bzNXq4rJ4ib
DnSCXEOOANhHvmCZPnVP/bvHbX35liR/2OImWpqkluz00SRytf6+qrOCFTg/ENlzFHySS4fPpL3P
c4bZ4rBlcjQhiJfKxJL13wbUnvlmmK0ohT9iJJLT5DSowm+7b2xmdE6kCZKIgS7gWb4r7nJ9vNQs
U+se9YQgbnJIox7lUJsdPvnUhCFYsg6psSSlDVBs2ayHRdybxwgKysXY9R1HU4B2wgNHeugvUfg6
sfaDYomqoLNb+TB5giO1Y1wDNaprqkeLcwGlNj5vviNxpQGFcJu20WuTjZ+I5OO8stkth7ScVVB/
qSZKhP8cIZ+kglXur0XuxGGtWwc8nuCzKbLKcu53t8LCuQPfKskZtTx6MfE8/e2+02hQSxDmJLNn
bzGxZY3gHNzmFgnuKO09++NjG1Hy/Th/G8AoqmFqE+SsADNA9CAh8+qZFb1/kkXAhJ1hvHve+9BJ
OJUW7eoY4Wt2uolnbEnvqo63Snd/dEiQyb5M7knnGDdlhXGwOCSZzdG3KNX5R7AKolJEdNM2TUj1
Sq4V33sQGcBrWkqZuYCgUYn+zRDPEOuL/O120qb6STZclOolWW176lXPvckS79lR0ItEmxv4n9QP
t6J0AhwRNJrHlRAGbqN2eYnLHm3pwqZXLI5l+3Uf8EIbWYzLi8lo1ofQMT5GkNohk5bhlBXoP7Pn
sWpovSl5VBl8anC7pUMtg95TB/Li8vTHVOtubAO9Y35BF1kt9LlxDV0hYtH+axMgWT5fp7jhEW5x
XVzvANfycUtQUFoeaER3A3D3Q6LZzvK2lEYzezDrSix9Ozanhj1aacryz3vuQ5DuEfz4eCNF6+8H
a6YQSFpUkIZB2ugTIJz470dAhKByB6ZUBy1nLxS8WhldYF5cO8FX1QNM38HLP9z8qq2f/RyNPQUK
n8GDyAMBSzDZkhcHgE9/Zwqyh0xTIwEf5I9EHCZ88U/UTOGgqte+IRx+lub6zT7zjcZk/cdeuCfL
EhdilGnbr8EQjO2zqFqEiNveXG7bHS8BKzctjpfjACgTKUfdo0GVdzYwyvNovkNqH1Xz/oqfOQbO
lZbYRBMMq8S5j0lMyKnIcprRpeKefsJNe3NNuMe/M5PCQENfDhnH5znYCv5k8LexB7vWYsnp5hLy
BUYAEkn3JQS1Ns00OXoqjm/jB6hB14T/e/twsucZJtofhmB1TsyKd/Fayxxq+kNtFxDIpUu4jXty
X5yiFux09ZgXUkTPpFdUdAfKMLuy48NDOPBRgEwlTDbNBo+PZh0dI3O4toggTRq6AhrCDJ82EX+5
XhEGaKVjoXoiTHRgOPPxJAv5UX2fKeeIBHk7G6WkQAXkA3o2/6QkGfPPMDz42oBtmFY/W1bfcPSJ
rY/cfc+F1W3CibkyEyK9nWp9X2YIOXiIvSD1I6qbEyT59mdmP54m8DQycfcYHs4YsEiECfgoGKdk
dwQARjXtFmrSJoD5Plj5TrYk1hUuRGVOTtUGk50oDX2CGrf/d5GxkZyJzwHN//7xy+T9t6kkdQt7
vT73B+s+9ajeyFTbD8ApCKD5TYdLmAk/igWex9/Wpkww2btYcHJ59UuNxLQVoz6rP38trk3CG727
7KJUfvqrfMxyGGntLeWOy0d2dsYhhSHrQh/3hiAIgHP4BpQrGZ3OyuX5gfgfoieOdITR7PAHgRKq
rm0CZOK69A+2ips5Snrrnd7ouU3wkDb6nRN34Be6touP803PFNkSvTwoYXJQFxcGVYDmw6YPImFF
fjaFLUdy1OZJbSi/5xQO96LzTmItJhx1sAKxlFHszQIKNnb/OqAx8akW/srwSI6W/xgcd0adN4CF
Vz3n4oqXkvEDz1cmtXnH8Ly6zgNUvEsCp29n5gOmZ0eJq2Vm4veqHTnjhjGBkxVAcAhDmVdVTX44
J+X9xV35aHgJKBaCjiq6LibpZiYnR3OfiNuMgwp9XMWYmtO5mpuA/ruQ8HXGb9/TfuscYRiWLzKc
c0t135UwpNpD5KfN4nvSd+atceZRysolfpnukkJHPgTDVPcVblL23+O36i8wWRwOCgaKVlf/uxFD
C9kz1SVDtl2fiENd4mAQ+CMQrIsI0q2l/rIXXQp2/9YMzQKu/itCuLqEY+LFEEVbIorK3NpTaR2T
22342jA/ZzslUOLHVQvGLGDg1HFmOHTA8tYRHnWNxZhR0TFYLk9VPP/t8vFj1imENO8dwLlC4BbX
U9wp/H58LmR83N/Uk78lgz56y1RbZLYYLp5ZHff49MyKHXN8k45Zy0UBn6LK5v+/76eSnxOd8ybF
/2OAA9jo4+lEisj/sqMCBRjcEGHOtdMAhHr7EENK/jvGEUedugoMWLAPxitcrmH9ymb5lCU1biK7
rsVmrvlohBRj8zn99EkJ0xLQYWkFAeZ5LLPNYwJNlnMMxSPx5WJnvEkP6pJbpqrgoYe2Sihyirwz
I2KEJUuvNf5R654+Yp7AmECCeMO+Sm1PVtXAeB4AtqciMLtH08zYS3DpN30FqmU0ltpsmJ1KIEXT
mioLpdyxqirqBKf+D6DTTJncS4s/AN+ojU0SvxFzS8yQnyliKHdjxkOu13XxPgDd9QBkIdhnbGVo
IqEHqwtf1K5IdG3rVNT3d1Xhy26dUaKIzEQHF4hHNfOfdKYkAH7QuAS1phOYYx7WyRRrF+kW7WV4
bEv9FLDCAhr5wIdrsS7yPbMXdsQobRnPhBJhKQ3isybVR+9rUQeGfw93NWN6cpkuPjmHce6BXOrC
8SVs3qEwV9IeHMRnWArfoUsbm4tGLleUXwv7si/ik/4dYx5DzHeaAGTH99UYw7Lf7p+bnb/dod1B
V8hTBpSh7+Pc8OPPVmcuQ/UtwG5TUuRfsc66pAVrMVZeMXipVA4gvbnkdcNXM0WOrEM1r1o+gi6O
7n2nnCmUk7ciSdChmIZPgLfyw8nsImF4R05nq11vqJFN55/xWm/zk2EhlOHaQgJOHU/vQV9zOV0j
mbMYRhT/wfal/1WfmP/ex1acG66tGep+MgU3wMOtJVOFKm+DjbKEEq6IGvVFOvn50nhiq/8Levwa
MdY5Jgyxg2qOsa2hY2VDwbb+Nw3HiU03e8jaOjlsZ/eXNThlS4HaODZL+dVRSg2iG43uesZfCfhL
KzU89hF0pFhLES60NkYuR1WIJlcJuBCDEHfQa2inYAYpAonJtbGvWWQwIk/QR1J003ST9NrdLTGl
tMpYOOjYYYXW3w2HTrovFdEHu0kxJhu/fNokCJS5fv45peGkgEBTKWMbGkP6kSCU/IO30z4Ubbv8
pcNyjgZBqZltOICSSeuvvXeDutoWsS0Xex1QHxWN9g4MiTXP4xbUuHzUp1AyViYrhGs+z8jrx/wE
1rpi4qjWNnXNO2DyDSqAGSNitIRuseLGUte4rzjfS5dLZQTbm8kUPjawaTsHldl9Ik6FWExX+612
6yvkiVAKbS30IwYJy9UgE6nZVq9WoYUTdVOVXW/x9cXDGHYrpLmLlE08+3CQnGNi6O3nMeZbTc4C
GE09bdrsKgIs/UjfWHWHqiEzfS5bRqaUImz8+nRUNpAQ3aN5J114UyAqcrtnKVcYE2HYmXyLTPf+
Ddej9bFCvxu1tKTjM//P02RCxEH09UzTjB7X94DfsJJRYO7YC9XAM+D8pe/yxT1bTN3s+yIrxWjC
eN5NuhHTX/e6qPqXl1cFEGF5+tbSno7AWGSYmTcq/WHJYqEplM9UKWx9xD0M3hUFd14gwPkXBjY2
vwHDT+/aoamooG76Ecj4+rNDvfGUNQWV9ev9ejNvrZEVukU5tMXmzUPeqTLeqfxAd931PX+SEKOh
fl53jcysE2fiPE6IfCxtrvDzDPCK/08FiSBEhcvR6ECXQvnTPxVXSDxkaTXxWzvt2DaIEdUEp5Ru
LQP8ofkyhYPGDpsMfDwiHNKbWQe7zh/LvpRuB3h+CY3CRhaMh6R9/5MxB6+wqXH0xAImbPqs+Ohd
jviCskgXk05bhQAEVBqhb1MLO1KAKR3pgU+0HsVpXNRDTxMjmri9MAp0csby+bRRX0kXv6qLk2DJ
69N9DM91uMLobw/qpABhlzJiJ0ag+n8+lgTr/wXku3RLUm/jSHuDPOASMPpoHuniOvKh03PxF4x8
mv0NMieUP3rP/FeBUuUr+A7hO407I5JjcCOZVaSgmaiEafoE3cCqJZGUD936OIctuwrIGyEQRssG
yl6OgpOQ79r+JvVy1n6i8NqIlmkSJR1QsFF/Yvh5iQuNpaOn9WdZCzmFgMz7etCfvOcwtRDXr7Wr
Oc3TPkQebn0AXIU1JDNNdlpHHgFDxFspJMRKMvKzy05wJcg6vn1k4pqV8X9xKJ2b5zgaC/Cc4u/B
VWpVFHQPB8/HBx0GhZIpM4J88OkmaVynrhHWKDwn8IdmL+As7w1wxp3rlzagj+/l+EvUOmTPz6ed
pyVkPWAPv7vK6dRqZ2LvQ07c2//nMgnl3lg56nO9dJ/OhSCV4xs7e0TlH51a2DqJcMoe4rG2WVZZ
XydZujiTne+ylwtckOi2hr5dzW/QYyianU/QoAp1dog6VbMBJtuKmdav9PGoe2n3+bKYFk9G8PMp
vR9VEZnJo6iPMtiLUQT4DePa6HTjrYSfauOYDZdLoj4k+op/D9YI9FL+xSTVJrB3NUzG20k3wTVT
Sye3EhTDYLIo0V9hFX2xbyQj89Nll66R9EAW3T5WPdOT4B4yY7JLsL2fyx/Jzv8tcP7MGci8KFSJ
vWf1BHRpeL/BJdui2K25E6Uo6gWq5UJVOjxS8SmRQ3GvKO1Z25uQqfZSCYxEB9j513rMwnFbOF1c
RAdKIjjD+LN+MRK0CBtXuA9f4XK4jHTJyA1tMZyRA7o+jFun0DztdSU4BbrOZKz+tQq7VgWX96zT
XhtbqL3Oo97qnBWG2l3h4WlEMPDhhmK3sJwjkriXuWG9ZSIoU1aCBtvnzq/bT3Mocs2bRyJZhNxM
aPtIGseXGRfRKpQAcglQs9oDF+VxUKLqi1A458Oy7a8lNG5VgWg6L0kG7JaQh41tlik2i1JxzlGB
x4z2krFFnj6mZvdPBLVLDSSybV+A77PyO1MzpM8AWrvsOhg/49xOp3hFDU3MbOr6hk1c/byyBABv
Dbpo9ZCFIf79sYofNFWwLszH8Iygv7JBgfMjrpiBNzthaA3tRdJ8qd+OlPeC/uaoFT/CQAkQTyE0
ZF2miPafrZWtROsKDkSR9smW5N6GkrAcVMfzbYtmLujK19LWugnTcuxx6fs2yLvjzb1QBoVxzLz4
ErqWis4YHHN1Z1dzCIxssKHfhoRkbD9cJ8o1hqZESz0s8F1Tcivx+1+HsHFaAUNeSoQdOFwyG1xK
dvUC2fKZXd2PeAJYY6Yrcxm78l1FDSUbYe4H2yqvo0+hMQLtPcLzOQwEItiIUS5prD52OlzhfZGv
J2ij/fU6Pj8dppjy8DEf8a9tPNmkOCxoBm3mESa1aLN+biipNNMDceOyrw6IiDXkTOBvDY/Q3HNV
gtorZ46zZ7/19VSaANcbOH6tF6+E0adAhCSvLe+sBZalVvYsAzv0hyE7uIZ2o3d3R0L1emD5ijMn
14tn0TbQGnQjTRe4K5FAVXT8UNwZF1lxnWhVIEwJjAwCc5ijCH5qYLBbUA7xBkJiXIvzQrQAyxq6
17Y7qalLCrCOlkOibOi0m55oYwl6hFWg1BHTRzNbgIlkCcREh4frFM/qEUn91DsFT71F19WcEn3x
RiOvK9AMkfv58GkhbBIf236S0KRRF+d381SlDPHGuV+Wbqg9RrZHhaIxIMLh8Ow2ukwoxhe+uKj4
NkjUNbe5vt+Q+Zx1P6KCAOgIQwmAIAck1uih331vUnOOj7g4NIJJ/kzcnUqb4KjU+l2xWC1eEFgB
NkyKHr8kIh9VBydZ2T/8nuLRnxq9rbgRAbiuoYmyMi45d5HeQJ26J+pu/1Ztn492OdqTLI9hsePJ
Z5eBuwk/lMFCv3ZlEkAIpeXdBYw+8llp1adBbgSqqcnRwUoB2DTCgvVfMt4UYJpJjhFezc8+iubG
kMhwRS3qLWmubnRvGL8kiygbkZWOkcTG3wRVysod++Lagn8BHhnTm2A+kntsxfUeKeaSVjXCDDyH
eJIEs4IrY8KoX+fuqOTpEYC0dv6k7oFFq7lR+l8DmzvjtmAf7Foci+6DT6CgvagtNatB8xkIsPcO
KrnH2AfS7IQO6DfIh4o1ft8FeVvERklimeLj5/wqw4w5YSb/Q4fwXLRlz3J7z8lr5PEnqwJAZcRG
NJ6QEIPIsAQV+FsWwN26t+GLY/e4W5yQtbECwm/M0VF4pjp2yRPrW+ZKHwkIlf5WqyXPhw3ep5nZ
o8n6WJDWLF1yfntieR9FxS6Iu0m9TjR2/8PVLnWfKBBCQYOOll8RxTPP/ZHIasZZuh+9LGEl1Gqm
dhveElyBfEeiHyxf5wIKwcn5SbXA4/cK98uPGvq5TTfK1zgBHOz+UZF0E2+EWqQunKFtWX7fkd7J
6ULRfvZQssbAexRRYFJ4Mro/Q4oylvMNTIt4aVSE6B6pU/8DJX8JNJ7CDDj5c3Fh5/7iIydOI872
GOMOcj8pdgwHbfJi0tAurfHdX0v6HJ36rPXFe9ThDKwsq0Iu5DAvSPzUnWrZMb35LJNBrAENptyc
KuAt2UogRwSu9bcaheVuGW83t0gqHxnWi8a4WLYMUCKbhpMdf41pkkov5snxrYwK1UeONAI7yPmM
4bv9QlNSzBYPLKcgiymUG4nmaSLeiWqY5KoC6B9caBTsHPAAHX56Iw7LgBC9yC+wXgnhGrMydtMt
jbFDSxc=
`pragma protect end_protected
