// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
eZILPLnGWYqOVACJxnBGQTaLf7bg6reZyajkn6etYq0aNZLWtLbfVx4nS0RgFMd6YSCFSKOKCUSr
N+XYXeu64O+UadvOvthBqKkQrceneF67eybiiatCiFzyatVzfpflwU5fA2aIl+yjz7miT06mQf4/
Mh6MkWZ8z0kuuvpOFhnsZabdaJHurgroOlvU9O8Q3t93j5OVb8K0+AQJqIhhgbC563Wx3Tj4fCM6
9XWk2QsJlTwPIq3iwqDdS0mY6l5XIYQIq5vwwNV12nER/+xA5dm5fBoUIw3XHLa7WkWo8A134S9J
aBpONFsrysSckcDFmeM/MP+a7F8SAsVHmJO6eA==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
vT5WlJvYgl/kh8GeEMn1ZO2rAso31o6PhJKwg7sVyuxfkmRTygYOwf0cAw84syo6+MxlINFvDDxB
jL+flmwRKO+6SzB1ymThVwJF3pw6Zl1FcfW9nSaxURnjs39HLPgwT1FePnOawGdZbUiNPUjk6ldu
wwke3aFn4M+9loPaRWmtybUT7fYmnd6OLUgPPZ45KGoMP/rVvvwqoDHzLTaAymC9fA7C8NTrcEjU
ghaOiND5pX7ulC80CzweUs90MZGAMm/0PPcymoiKIobHxi8iHx+kZU+7nEzLXw0iiGkRftmFmQPU
XuG+ZSJvfyABjdiMU5juKg8FJrzmRnnzfjg68zlpIY9QNcUmfTsq0NeTq23YoeovNcaMgLyh/kvG
odZG2Pn8luPvyxnlb04t2J6oBMX9sY6LxzHdgrAx704zylhbgk2ZWbY07j16Gjlyx+8wmrLG9ceP
054/BSDmSWdn7DMDWrMk2mgK/vakpzGWDco/Yg2gd0DvAjS4WTpcjhJTwku954DePbU5XgAJOsAy
CunKD6s1YipYIFJHwKZh0/CdB9886OtbFubUHncLnl90T41t63fQ1mQ9fgay8NZk3jXjiMjUoXHo
QaJpc25HensztGaf9wWXHb4OV2P6bHURtnl8k0Xdu3imnoWjKo7wXyVc2byqtG9u7puYgVYmcPdN
eqCfnF83ZUsrsrgWZOIojlmDjhF/KiLcqaN41f3tzRHoOu1CNA+8X1x1CoDGTwMtIFU2M1oIMxFn
UnVhzQDDiFn5wJD1liCnAUBpbF9TJYmTi0vTH87/06/yEeOImDd7v4fiMfTXNjM1AE7X3ZGPm9lk
plQdA8WA4t8lqmaT8ioRpBnRmmp6Op4OiMPf4D7F6shESlgnMPboLzNn0Gb1scgp4IcsUWn5zkbO
fRxq9W3rUaUhvyX7WeB0Q+vymaJL3zSbALsL7khl9Wa75bF7LwXzHmOEj1FY1Qynxm8YkKbh2iFh
h38eKoB1DLBBL9LKdqHG3bzWHGXxIpwTH7ht/3rqqrZDHokV59oEFVXojhaE39YIUVGpopWB3zBo
B/5iDM2K8tRgA3lg7WxGw3grH0M/1vUVDXlSf22DcjJL4Ug70XLCMUQs7230Zrr4doAMFzimuLxv
FMI6G4lSDfXVVOBUeb92gvunhatoOAMjdnTvYod8VQqdaASuP9vLAzZbnER7FBukp+oTwgcRQ+pb
h9t7UXfb+35b7BpDF7B4tvBWPHXw9RprxVnz4bO3EvMnaZMvoqXx6+2MdVb77PFoo5JJS+j39FuR
xRzcUy/p4L75pflYAJQwCSm9qcIciINRA+TvoefndwIat0+yKtQefh3W0yW4M9BL5YsH1J+Q83CG
01IVLQRe+YQxGbPXLR6JD7kcdlJq487wyOp9IC0OUlmTb8d5UlibXD9VINfwfpXzhJ2Q8sFO4/9e
ie4rSaqFndDIiQWf7al/2k8xWf/JcvhCe1g1Rl2OVkCTLRC42xH/Hxlkv4u8MmyX0cXGmMhh2Dmd
eBC3JrViYhbkR0Dqb0wkX6KF0hnUivNU2fqjZ+I5u64g2cR7Q47F1Wy8xxs08u07fC4KRrWkG5DA
cZrzoHa86T41doUASlTL8fbUO0eX5nyRlb/e1DrO4bNw2ZRpyhUBvsKKYLzTsISGeyVJhupXRxWx
+71pPvUoVhdKQoqkOgasPd+3Ea7TZvPL9hG4KzSWednKWSaWhIwP3SaNoqlKlYcs9dDEVn2ajyEi
/XLVxYVdK/cONutqJSCn/KnARLZnTSjotmZlx7Cp2BTt54HGs/W3NeVwhtSZ1uCsHHWSr4ThZega
shEotd4KUfls92thJ7mK3r5m8yFBH/2Fvfeh8rNKtEkNZ9RtEL3UPAeXbe/ZpXxaZbSoTmFJkwpR
AvnqhhwScDS7TIWkIb7hvA2V82tBQwfeADOcrT76UJ3ogj9V7pqV1da1vHfVE+4merDbFlbRhDJQ
1sDQfsJ4It7IKxABgw1njYw6Mn86H6clSrEiVAFISBdP4f0VE2+ypX38I+r4A6sRGS4J6q0chADA
CBA5qlvygBYyfPQTn3wBMYCL7vOFN8grYLzPmLVZnCVYhM3hboKk9O/jX+js/w7exRU+CJ11Uthd
0OpPNBxrZdZF4oI2FuwPJriTdi+zbG3MOvIedwBCOIdHQ6grzQz1YEA1qlY0xp/Uk1dUv714DU2D
pz5A6TjPURR/CCUDPRlwc4cwVh1G4SW5YhBgc1iVW5OrB+b+1NLmGYf7GCNVkTJxAgAleQZ8izOI
kiHNzUV1Ugz1tNLkyMEK5Xf5Qsi47XcIOMae+9vcj+sJwjLDNlgjpDqtaOSCLSub1RQ2dEDCgZKj
d/89iaYjWml85AGfzl2PINCNh04CrfEKwVGPM+9q0zSkuPn1F/WWPAjnhhLAcf7nSGutBRFqp+xO
yb+/OjucYgWmQUwsb308RslM3UimpHPVsfxzh/eDfQ1gDLcJ9uNpMzBYn8V1aGRs4sQsdHpbMeQp
51F/wmIJdl3EJ54cPK2zw4k24ZZS5hx/0yeAuyihQX1iPZPrY84xxz+4hMtIzkphI1Bb0BN15vFS
Pc6bDtkwDuZRCQgLefmtVK3M/SXqkHWzqjyKrX7tmVNfi8x1OAooFP474V5pdiuk4tFFh2BMsSoM
czZjG9u68PJR0FN6fSZEEPi1UFZnnCUq9bhXl4xdchl0n5xEkrVp9SjZdYvCtEK/7QRnjP6iYMwM
9U8tdwrYKxzlTqXk2YiTRT0DnGJmvsGjRpKDv1pLqz0JYPM6fZdeJC0BtQHLWchbZ7neCeQPlRZQ
/k1rehZD5RVMWLtCBhOLwVOpQWgVge1vXt8fZkNJ4lpimUIuJbcTN/xrOnCgCRkEDtD9cF7L83A0
s67eI3SjH5TgTY1dfJvetc1c6JVgNQSgpYi3iaoof9619bMVttxj+LzL+ug8VlmMh4d2II6g06Mo
L4AuIRs8unKXK45AzoNjr3MEhz9ehMD/kI8cxyT9Kqm7hH6IJf6/P3+8Kjibmc9MjVaWThz68IYF
2z/vcQg8D+urRYa/99CS/6mp7kQZ/o6DcaNBiY4prgKcIOof5rtYzy/Pg4qyRDjDdh6ijD4UJ+mY
rmxdE4kXY9ZTxXDV1fwNPBvNH7+oZfjb8981HRu+B2BLNrzHaML7PdPPaz5Zw7uROmipP4xP8E0+
Ol8P5UkMPDoAn4/sYa4Sb9bXFVyAvNbMDk19s64RDFYqrXR+NW81uEhI0L8+MQkbly9L+OE68S1D
+oNzlt8v4AnKAn9kdPiNoSfT744MH8uDEIdLyceKMtb8c2pnTYnLVxkNP+spc7rY9RK4FzJLrRh0
rO3eV6XwzgDIWPJW7trFz6IT/G4AgzomdDkNR/hoF4Le3SrvTO3bz5TefKVZNRIyAL2QjCK1cl6B
xJX9W+Tsqjmza92z9AHZ5MeFtrk6hLs/Q+MVpqFR3xHtGoGnV6WxB9HKXAGDN1tyiXd6Y5GxkXjw
N6/blI+cXCOPxI8fOrcPn5o7tNXjzyBXorH1v1ncORrr60J6QYvWUPu7bA3FodEgGGV98jshvxkW
CUbmsqfAr1fPP0vihP/QWz/pBiLSbb1LtFoQgl5u5oIuo3hmXlYTbbIX80O0nFiSQtY68zT0ZD+A
ODSnQ4o456O72lS6WX+cQIxMB9/OMTLOr34LSq5zQ4TcsoJboQ8zHOec00ibVNgdQWUXATrF5uFS
QRMCv+pPgtidNe1hcc/mCJqRLdSvCpLqvOvs5vup6NjD5WkjYWywcPlxVy94xaBJlsLr2n041ZWr
uVIuskmC4mngQrbzNIVOyACU99oVnXN0yx5uIsuU76ycGFdIBIXSUKS8QP6NdTz1OGrYXp7ljt2X
CUYHT9DabSDl4JF1AlynjB6aauJ98BhWMnrDGEqB+BR1SSzOc4E6abeacKe5VRoxA7gEPArqY8tM
CmVnIIpPnRBJFagDgCk7Jwa08b4rPulCgiWeCM6acVmRUyLeWYdv8OmfbKw+YqMf8iYw/HaEhcI6
7SAB4BUQxKfuro6pp5xt0+4Af2Wxkc00SwA7zg9s0i7Fpwyv09apwHg2bbo1pDFRo4UfYHqVkoQR
9esIFNM621bpMFc+cnj7T1EQVHxIgDN2eBVCL0Pkq4sAERAuwD7icXM51opsVBxwE2Lda/RbXIng
R9w4nI47llzi2pYTyaeuvFxKx2meJAZBQFEI8T1yQoRwjyDPf/7WHS21l+q0ZQzl6D6EMYSx4xD5
OB3XYsdDZqWTzVkih+t405p8ZAd2pcaaG+Nv0oh3kcc/z9+XADdwLRLbma341JVd2b8YlNhth4Yc
us3+fGJttXfi77Nt4jjtbSg3vSMeXfPQa+Lf/Ks1MzcT2CATu6mfBrmOIz6Y05UY0QDMlt1QG7Sr
x1+p9zgAQQyod2FNZyAbloCkNWBGGSMFjr65jUBhRtZ9HXs8E//Ekx0f2RggfGV7sGUZhKA8mRpS
fK6oOyXaYSTLeGo7WJkQT3KWusHn8PK+5z8KmONYp/QS02YzJc5T7aWondgQlIb2RBAxlY0hDoAk
7VL3nSep8uFxtwQz5i6Zp23Fs1t84tvk7JgECTrN3qHmrNBsujZcwpwI9OvCb0Ccb9LwFmduXavZ
Fd8ZFfuGCqljClk2PC5TK/2i4k8zqgZdhb3wkAPO4192vbZ7k1ErBtDuze4FHMJzmZ3ikr1wsl3c
h7s8XEbTKqKoOUzQ2Qf7U1s1KnezQ0RMmek7kCHh4rc1fe6NQT9rsqG5vpia9yqBZt3VukBI4fmp
7drNHYbvuM2XG6QZNeBL0XSRfFjIzFF/Bti8Y3zSJKsn80ENuRNjHoKU4m9JfyMH2TliGPSp6k4I
/PBsefpfbpc0FpyjUh3FcVO8EHrvCe4f4nZ1iBiHMEaL5Vtsz4KtX+xnCeXTBlF/PDFHEMYYJ2cB
N69oWXHahi6iqjXdFhrTPBVubr8IetTcuwcKz5XjjImrLLgR9xLfu5WCr/wr7v6Nurmog4VoM+ve
HFMGl1GDK3XEWxm+Ke7tUtZdQHFHyNNGNbrbX8zC0DQ10Tngl4i6wiuhy0j3kFIJ3igfkjFXu6zA
J0xSADbT/3WCBVK6Pt9WGhg9n9S9MNtJ4zPYPuK2Ng014QSPWIhFVJcDQSQD4oA9rQMGrMgPuHU2
f5mZ42zlRc8C0p0yb12oJ7dlsVRw9RkxLYl9xaYVGXD5xGY8ozUKjUjCcOsTGlIouZC3dDUWAMSD
yY5g8B3pJOMlD/9QMoh22z43bR/xKnmHgBQFNfN/4o0w7av06zLSYwtPLcITC9kZiUBxjsXhIyQu
aanoEnlPr1uzOUfesFK+2lfdOU2Vb95WXEYbijMO+PfyIBnTCENM9SH61+VwoUcukE+edUXBKTNu
Gh2qXHAODtNFtIv2hOW6nnrBujdc7axAqBkV5Vty01PXC8gOE2nGsLZf/oYvz+KfiURvL6JNUQhZ
tZjKFNAFCcFl/cxbSbzbQBHYvxeGDs8DwTDD/RG7IOkzZj2nwvKdPgOt1yFHyCHjP0cAE7cGxonF
YLzS6fi6AwBKHOvdmx1oFRyItc+sC1Avyr7dV0asA6gXMhG1FeCFIW1vFVR1qcOP5Dxdt9quzoeO
xY6Mfl6w5Jbm4+7AhyYu6xxiiidu0NqPNS5KKpahH7pDKFzgCjrawiA8q9MNrl7lgHn+Djk1kYmz
BTUod9dAqxtfSePvvBSGf3grVsEfb48O/6UWeryShw0v8nkDF0m6fORm9JEoTjHbXkn8y63KaLD/
w3UXU8FXCkYaTdp+EkKHFefULjE4N6qsx+eIBRXVT/KJnwfmqB6qQ/NYAM834jYTYw4ki7+WBMhZ
+Fg7npkvFycsdhGXw4mxE4Q/IKYM605P7T+gPqkkfaUB6/VHd7F7YCwHHCxUa0iOAukXb5DWShdl
BW0vQCf5/bwTVCSR26SYARtANnE8NA/bNg4VXWRPqmpUr+BuQQzIKhh62vDb9a8ACouAwO2r+Xzq
UzWHCTGQ1IHiZRxdtENWgYav27o6KGTt1nky+4/MJlilOb9E9XYlfSC37rmSSa8s5QlKe5Bg/kZ9
H9OzWDyQUZC4nY46I7Kvv1GitGW5aUnLiK7b5i2ENzmBkN8yVtRb9ANmYjDV06LO706EOpyqtpiN
eJYf+DOPm14bQ5MmXlIcM9DymB9HD2QBdSvmP+8Ucv+ZCSMKgYhcuz+cBJuvpA/ZOPRbOyliEBBl
a0UkPuvgDlLHL40dtpALbWRwtc6lZuokDyZAHIS1rKQdavgQ0w/vjMGtcvgP/Pg1rZlA7uy6xxZO
ttjCuLJt5QY2aL8p2/+wmWMzJ+mRmJ9bpcCxuFjvUqH9FEt+4f9RbV3ZCKlqEbJizihKMGpF1K/W
sJQM5EkkUW+kMCcjx2gLMtL4jKbtpUPy68xEcA6MlHVu/LMrjEaHRNu+9kA1HX11UCD0saXUSe9Y
DtLE7beY5n6AETz1yy8rU8Lbv4niFxBOvOCv6drc9l1GPIexGB7fQSwgXAqCLMeV4CdpUXDLKuTi
qjt4axYcyuClf46huDu2itx1b2D4VN01kF3QnmjY5xyMZF4NRJxmdkKJQcu3/Qp6+7j1VrGAtTp8
sTJ3DDw6efkaxwsGoCGVg96+AMIt6kXSp0+AYrNn4KyHUmU1L4c624JuxqQAkC7qT4wW3UukZ9u/
+yIJVJhp7ewivCmzTPIbNYNUPIhXqNrDD38BP8xMBsOEU8mTI2Qk0tv+oflnUyhRdbCTP7x81EqI
Rpak/omMg51ANkIr/u51X1nlOpPcaDXlU1IckGCGkEUZyYaHDoagbz1cyqq/09dsfxlSOf+EVMxk
qSnkAAQNLotU9QYJpHytpT2yXFqn8vIAlNm5w7YtCUgBxLmCEwmcxWxnlY2g+/ERDX7+6gVPX7ql
KSTIDZq8z1nkXoTh+Bvi8UgQPVG7K56dGcWk5gu5PiiIY3hptN7O3pM1OnxgUeMC66C0Y0l5Dpe5
Q5pMIbCdWPERouu+gell7BP6DZUWI7rwRfIdikraTo75f6Cmco+mZPnuX6N9ImmDCnYvJR43eX0f
/BO7/yerwK8vdLjvriugaUkXpXELLnhschBrCcXQ39BApGi5hTX5itooZuBw2bwMxB+38zR6acQn
P1DiKMpVBAtvcoeJZ5jh8x/vHXfAVDKpETxXU9ZUzMSunNUo/4VLglbu4weehp+8BPk9uM7KuPWV
ptoUIygAvzuCmuSp1oWOnqQmx4Ni1/Gy0DJsq/92HFLWpaK9y7O2boJXY0y/e9hd7MtCiSNYO8fn
9fVQoghmsa7sOTg0YxHB/FcC9PM13c+ui7IgGWF/ofd5G2valVtDO/KbF0XB1szEzaY+/Q6tLfMI
jz9emgjC7DvercEiqssKa3pI9S1Cp7ays72vMJtmkwXU7PZRtFkNKScb45h6lU1O5sVwYqhI1o90
dBLscSjK/EsZTANrSAAUMsVPtwMEXHR+EeSRH+xKwelBgA9Gn4v3WgeVbZqUgDhWjcdO7mRbcYqF
DPQa/mhNwUSEYQHL9EEW0Z5wZTjgjmjtlOrWN+V4OFW0CAoyY0HUUTJICBDdpJ0pdPdJ86++n9ZI
CbxprhiPdirE3Zxr1TJdfsa27IKaWUQ4zKkbLFGkPa+b6BxVzlNNNKAs3rgGxuTUb184BL2URKSC
eD/VBxedmtWczaBluFhe0Mn/SCPhDaMSus8o4Gl3qIK0MQI6o7ywYyycLtQf+Jr8TYnfrSSU2zBH
0axQiqP7x20ghviJjTmxzFh9ECFVkQyayQG4XFm5pL6GeeDdjOCAECDm6/Sc/q3DwjoT9fDQqpGY
0lMslMoibCA7HBzvNx4sxFx7BclCMgoFgxT7/IXHTDE4qwdMexx99nEMS4ug+gDPQuDcl2mTmnJO
CBQswYvQH2F74d5PFoOq6hpNNyAnlzPz8Csg28O/NxQM823jrahgyLd8DBd/0LP3I9hQ9kcgx1dF
0hNLKCCXP+tcj0ljyHKdqNDLXmlUT6DtkcOw0KkB36/aKCdGF8Xb0Ow3NUMNtny/ZNo+Kv2W/ArK
vZ8jEWLTgCB4IxSF7Mexd6Xw83KCYlcprtbh888sZ7ly+MeFGjAhzpegRaou1tundvFMpYpjxqK8
b8AkhpM0pj1MZZeZMGPHxDbn6UkSWR9DHN47dzrDC96k9AxpG4NbemQLk3Mt/fTKOjoQbdC5Lgtt
viNSXdPoEsqAY2S4mTSrYRm+pUhOC4pBPW4NK2zl029Z4X/YcSIcfcE7lVbmtNJEmtl+wRpwiF01
pvLL+unRzMGPtp4BlvD6xNxgYZOg1+bdHhlhwjgHcYwPDuZZhK8GqsuRYQioubtIWIkPNg4VkwcA
3jPd5bjcgGU7m4p6S3ATTZT5VPlWTUwypLNf8bqye5RsDoZUsgR1fkn+AoeIjXZzoALVl079p19Y
LQyIpv0mD++1pfBFKwplecn1pHhoNJmP81iVIOIKsTPgCpYcmNxjFWiolarvkVHklYzLZqPg/r4Q
P/iiDvM3LydO7LQ62LFo0dYe7uNnbaJ0+w1Ya/McnFvrFyoBnkAxi1LCCBDhuZoei+L6e1yEKeoM
L5Zc8hu7w4D3TApn6AHdriGplKp5lh+ON57V0x2SW9txLNIpcy4s4JEOt63T93QJVtqE636UooRv
sJvIU7Gtp00YIfK9mtTn1my2BmfG0H6WDojJ1JbkyvEVUIN7zh/+1qVYtACaquc1LsyIJ47FfADV
LamIUTG0oikpdqXw1yfRF8ca/18HhKr2Mu8ZRJl4VHyJUOguNQnn3XNb0/q7d4MxKoNvVbnuRK5h
GW9SRPwuxSR6OniS188s9yWpyR9DT0kiJ1nw+wCW9nskf2KdWZJXYIAGEyZhm0WbXt8+NCVC4NbW
PYGIUgKRj+9p2NbZks76GQ06Pss9mPoOaGQfxsYexkY0e+pcGMsLJmIoYpXyiqghyFZ5o81TGrR0
rWafrUySwSrFaTmlAHhSyJ5UXPvyE0KOMZnW2UqoRMa8whv7zFz+zvRs7lg0nHHatVE0O7BLedo8
kv1tgzusAC7nS2mILTJoe66X8ua/L0W8qy8WptjKOYcvszMyZL+bxOfVHPKiCazi8r+qM0e7tAJP
8YFlfIjkPgyL7T5JYrga2E7r++YO0vvbgGpCo/Vd7UG65FtKz2TY4Q89r0g/z4XnKsQxjXrgE0rT
8r3nZ5v1HDBCW9BD6yyeM7fB34zfQvwtl9Lh9xTfeRLV42AU6zPccQfl1j0KGhFVdO03aiyyhWzV
AswkY1KOZcTnpXPBk2skB/Icf2CcTe9vTaEETLa9tupWmJWzGQwofxe1rwqc3y+R7Pf5Y9q2pxE4
Xm0ZCm9sHuf7AErwxFkvi+bFe0sSUwQbZglX14h5HcuTWGBgncCqU0knDK184nw3pT+0GL5nRaNY
5W/AtjBRpCTYZrKAsYq0RVI42nugmv3ERizbNloC41LjD9iuLqoZpIizocAX/7Id9D8z9S7uClK1
6eIXVXxsd6QMtNAeQ/KZyoFwdXS3q9VjjaCzyGPUBQUDXDvFfmWc2+F70V0kV/7Kq2Mwojl18uE2
c4c8umMPBqvCLCWrgzioOu5GMb8C24V75YfUkpyPQhzgOfWEOJwBxDy6WTahAf53RqwYxC8Xgvin
Y6TT9FPrSRh+Q377JhLNcfIiBjYeXX1ONtirQpMkT9jGmimqKHF/BhcvR0u09GcNv7yJt4znFd90
GDaUKESQUUTq77CAtlG9RwHb2oOHr0rW8ve4Q+rkNGLuv4Z6HLBMpfJ7TlttnhYLxS+LqMYBFHiL
rWH4qEbjpvwV77vpx1Seg2WIAz+1PcDRH317P9+Eqy0neeuCw/elNiSjPp+fER2srReBxRvvTX+i
UJoBYuozx9hIwLczoeea2bZJLSH2RFwpp6fNzWUX5+KxhObiFBiDgL+XEmYyCcslWSGfC2/FsVqk
vCU1vXxRMLSYNjQfHpVEU1hNpQENLEF3eJl/I8doP80lJR7UkrguIbAxUiOSbVKmUeOEf6eVPKLl
+/j6pkG64tv8zH/lrUz4D3fLueFgftInCBwEWhu1akgH5olKLrlf97/uO4/e6ZLsncw4G8CNot9I
9UVQIFYr/Fpn9hxXP3wGYN3kkNCzGwu/HSfVcsmj5xb0r1K5bqJyZZMOWMBEGMq3K2bJ921HK/Lu
DQRh5PSrvHw2eQehbCMM56Uc1egoZcwjucuuqtYo9l4Fk0GKJaNUrBANGAeHzayitpZ0ANPK3rSH
20Bh3EiYdZcKTH7y5To14cb7KYHJhoPajOPTnJH+KLq7Iv6+XNkq84uVAGHMAwy4FrRg7Klang1m
S7wWuEV/a/OL4xV6qP+8WHtuwyF2D0YxpsueNZjNFokB7oyS+LQ+SfvoJiET7DcwuPGC8GiNIXIw
HR6dLGXy7In3hGCC/+hvjjMKuSuXfcIcdgyvmTSIEGo8gV1NVu7NA1f3mRplOJsSWaPpPs04dfK+
G7x+iRIq+rnL+1qVbbOhL4AjCK8LrRtj/FMrDUR54oegvQNWjQj1PhyuUMfdTCrhqV6AqbnX+D7f
pDy4rRqqEc5piJZlmU544GwJsO8nPa/3TugpKBe788yMpTgqxytm17j2aHA2cGxmG8n9qV3CsLrb
fKwoXRXHi/gwiRkFFFibIRQw0QglO/gjeRKpgkJ1EDJ6CGA+HZzZDUOVP6Vf+x+wY+Z4Ph5lZMOi
DfYg8LoYnlAI8Q54VGMk2k8j3z04rANhJqqx5dEf2YjJtNoSkABBkBKq8+rk9xwC3/kN0mxR7rxm
HzIFLmPmWeWuKiZGuMI/VIWuEaw3MkVqbckkY2OQnbTTECNK3STwu4YPpejpLhypXbjJ+xGKsUG0
vWtM8b0AVAeKPddYgmb3skMs3b/Rqc80MFQAYTTIyRzn6bTsn/eALN8NmWd7xefe3bLzv3ZAcjCw
X6/3SRzIX0luGET5UxFFzVzfwjRIMaPfB16x1C3IQaDBoMZ6kVx0K2J6+Y9lbUrmzChWEB3iFbdB
SYXTj4gLYdtHBfcd07GWRpJhgC79sQOUCyKjkyakEsfDOBHGcS9NlkOD1xzU2zsvrBqQGI8UX7UM
I/lsLfd67CzxaCxSJTPd/NUGLjhZV8IdjJ0Vy3AHiXf1P27RHihGXHcgVt8lxyh8I4Zn8OZxq8f4
QNWOOkoBweW3nVMlGEHvpsO83ERNi0F/De+EzPj/kUix5YI8Fsypfv+37ImmcKmndJDhmz5c6Oml
PopYKnM04muTzaRJjqiqy/P1PiNoet+54WtjFGoHFOB6JCfZ7E10SI83Tti7YGjFsQiGVCEvn8sC
z1vGB4lAjxNUl1GZ6fWEDdYGqoZZvKTG8bbIvDpjeskmzv+IfoPuV8F74PhTt9VIpZrVe4mkNNpK
DAJNECiPoAALONQQdCwBM7Iy01G8fxKF70KB4H1K7KUKXom36GAt6yvH+2Inr7cdrFyUsFDL5/0k
8JZNHlIkxuVn8klaXjuT+ihxgk7QJfXt4WYkN8RlHAq7JI2AVUDEJRi6SCOqIFJW9C72KetwIaRJ
2sce7gNJDi887Aq5R1950SGF7MkEBFLU8HgufQ+BVlWGYJUH9m7F/cuNb4Q+u17alYWgcWLYTMLg
Hn85ec2HQie5qaCg4v/MH0Nz1vk8Er1lWoqjTGmuz0RZPf3LCuOYSMUM911I7tl6Z3Dhy2sHhIVC
iCvnoYaeTxovIRaRtZf/brd5jfaWeom5FZYPQd/V7OwxwlIHIvJQE0RUYRIeFLbswxr/UaHiO16o
1zA18S+t1nBNHZu694XJAoj/waGXPKrDyNyzvSQiCi2ox40orZ7OjYNZoh+nBpB6hFwRaw9muLDd
lqPr7SGOQSlXDiqBlF+Rrypbmy8x8pp10mpYiRtJSvGr4fJ52HhTdEJs84FgsmsZMMRr2U8ZiRnD
wkw+2+SCN5djAOVMYZ6DfeMVRIQht+yWz3Jdud+EWYzUeg0JbZTsobvaRVSw8Su05RONJ8orEF1q
0RW+YkJ2NlLlsW/CdCVZVa6r7ixPU9UtxoT8C92XF5d7vzlaXeTkWBXwmG4kPJkYNViIj1hf/Qs6
VrHNdbf2qZTAumSb/NjE1yqrisbFbDXfYY4XATy1JssuTFjtH3TrK9co2aZ+kvCfFdpR4NNkuvPI
ZJ0A4Wb/xjURsiEWJaNOdSpKUAqzP+2tNT2st99KTchX/BUS9DAyDSjVze1lW1+8hQHSCa0qYWcN
jVGHOy1eZUK8iRaFCAFKcGgqA2pwIQGWYuz4fOkB4Y9yq3m7Xh7A1vw3K8ZJqeeKpv5E87cJbQKC
Ximglheu5MoCNbP3sBQ=
`pragma protect end_protected
