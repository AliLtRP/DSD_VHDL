// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
pbjvk5T8alvGPU8kACWtOiAuT594inOUpDsdYFg/uKjKpkBRYwz0+bMi8rR6bMscXoMDMKXBIjVn
dkZ6cldcbM8XdGjpDXJYNKDDKphOj1LE5uDkLkHo/jlzv6K0BVkW+Sc0Nde7rz+jyO55OGrdicaH
Hjd8VeORTp9B9bXfVEo4x7gmUUULsMlUuFBfmZRi99F/K3I+uLdB0LHy6VVm/mE/xMtnAClL8Tiw
1LY7bNpEHhh6FD8fBLUAjKeFwNfU7uiewF8Uf/cUZt2wpjV2o9QnSWtB5tGQLvHJpOAWFdm1ANEx
QGJ1085kQteHYbDcAyIfStv3+677kEJiZnPNSA==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
VJgg6XTv7GbZJZgZaXNOzIU8J4ynPO+2FMcJLtmLawExEoneYFDTkL9mQECBkY5XIzQJ/HvTLoc0
aQNh1Ga8C1jgFiuh77aiY5mklUCUV8yaR4OJeRWAux24FBZmogZempbUc3dB1hJQAtvE4igt2KVM
/fWmIdFtzwYYAWOMViSgM0lMqpdc9X8Ek+2aTwj8zk6RXSgoGRddCV0S7vLqHWOII2C69xxDRrkD
LenUXjR5g25miX8RYRhWybOol3sj3IkNNOYzKhuK3fze9b9mjw5p7tUPPXoZ7vp4S1K1VeVkx663
eZdcq6D0xBINOjJrtFkqMDX9AyeuASeN4bAx0B4GCM/5a149HXAwlnrRg219zzfFMLCQl7feUXjF
3e5XPwugMEbQ22lyJEl8UzMI0/P0yeBUEEEwrKN5wIFG7IKvBE8fQtQFyS6YFlxfaD13pHxSB+dF
f97Ty9CChL6xjpHLCnzT39OyrkD/xVuLi16VJBstUrQUcr5Eb2HIGSf/hZq0+ZcBezivep+HIvNF
o7pjH0rhIjAvg1+VJxvJcJ3keePquVlSBv3gErNlGVSHv6ga/7aONnkPcwzpvHzdxQ9o9HrW2jBK
dgTSoUGrga1jgNprHodJ1iJuIDpZ5dgM462P8bWr6S9ME8g/99pTsEy7ZpXa+tjXRtbJMWbYSCie
gSY6xon8roGbsntUcBLZHK5YlwIIA+1YrSOdtcaed4kHsUpWtZNtPr7T4bX0fIKsjOl62Xnk6H9M
2Ocef5gSQx48+/+rtnvZTObuDNzDLtGlchHStm6lAcatVGIfI/VEjGbwgNVGlTLgeQYvyGVxuqn0
B3tvpjLvjNjy+ED9/ZOMgmAeGP792g8BnCt2pQtsXuxYkJ124cTJ8Asd1fWKzXrgIigyJEQaGY1T
MgXaHkjM2o3lkal26nINuzrn6JUwkMWDrWSSsKVXArEDDRMtqRwicJkiFbEAUpoAmgeAZBL0kE8e
AzqOFRSa14KK8w/nOysKuXbU8n5159I43z0W4bKma8zXwbceYqF83LwcXpQYoHVeWNPAhGVugSFI
+YS3WlU4aaDjsMLm3lWfN3mXzrmI0Vg5TvakPhFTvfvVAztfnlpI5IzCd80Y8ZK6EbOVM6qZ56Im
5N1gudSDWYffWSisGqKSLP7Fm4j+jgsWPzBo8q7gZ/7rOForf0bGQZManBNEmtMRAST6gN0wiyAK
uBsLmOu85Y2psImOQMn3HzariFTTuUb/Xry4UJiiG9qHipJY2DF3gKCIuxXJrWoy8yOLNSDIzDog
s8xHPRQCOkehYHztD+HrtsKyNiYiE8WtaGIeEXMWXRkI205LevYxON24P3dKliVXhXMhwiFE5tib
SOgwt8SjoYypx69gLwOPZ6ObZM0DFQ27AI56F0+QgOWmBPHKCsJvPaOtzahTLjXKRxrREU6+UPE0
TbIP7mtVAyneX3iVnehgbJ/K90HqHfl7tPUD9gIf994FPkem8/VrhJJLHorJU6rPP6J7WiipwrGK
NuwzwLhGsn9nQrRxI2usrK6h/X9s99YRS4QyIghmgU9LePLZibOie7eiHfhVrmmAoN67dodMXNLe
rt9btzPk/+lnOQvNUFKTx41wlaOV/JCIsPpLNjv8zY/X31or6vwaiDzyEVt4vgGVlsiGPjS30fni
sLo8b02zBlxZQ4T2G4xD/e8ShMq01vuRXKEYBrGDMJzo4WNFkyKPhajC4w+DcN66z/k1+2WZJ/W3
EQ4QYw0R4Kj/zq3EgKWUTK/0oPKp2x08rWZuOEYIPX0E28LW6H6a8VZ+ds7BqATiZo8x6yOHJ7h/
2a6Hnfzu9Y5dxTRDSWTDDi8gbKnf/H6SO6T1E4ntbcBxRLtE53e9+ilWzZcPajD2OFQ2P+SKtaY3
QZO4WeGFNR14rK2t15FqJ4xh4h/dIiR/hSUlroR9kTl+UOawfwcy7GvVeiumDvKK0Pwap3Dk0CUx
FsL2da0dreHMsNRsAvQ3/RMeHFWnN/oxsWPnSInXKnMqeuRIDyTHtsUC9gMJ1qeQnNRtd0QXlXsD
Zox/udKeUvG7sNCArkjAr8SSy3IKXpuhc2o7+F852Sz3uWBqLF98qx+OtuUGZ4fer1PXcblWP2Zc
eTySfnRrZLbPE/EJd67Kfb5ftFBNhLHRjwwaaDBE57qJOb/5f1ZzdyXK5593JDWRhfB3NVpWyWa5
dbu/WjnLe1ZMbnGIfdRjtxJifPprtZbZl70dn/ujCr0kQ7qcIbOBO57QrL7smzeujAUdUVViFTx3
+MWv65sWaj4IvgLF3AYYglofOusQopH5IyxOVKHprINgmvnjxwWhbD/fGNltvK3tUvAzWfxrAsMF
6ilPZdpaI/jz+W1o0jkFIj2kgBsq7LxbbeoiU4jIewEoZrEQ7oMiPO2ZNAmi7diXrkC4snQg5JAE
CPRTY9XB193tXXEayn61Ft/0JeyKOKMgGCz2zoH6S4QAe/bgvPGIFl3TgjZWK7s1Vrm5rM+sa4Ho
54XBsOCb08B3k5yBt1HcJnEEybkdqg8iLWNKR/pAN24kbVEJCc1+JHqhi5ZB/t9krhCtUxcKRxyl
XR5Eyb1Ygk4sqCdmCA1CB6kNCEObBZvpZtnJQiPtcC1g9kKxMl1rsorz6fFxTUMY11XYhl1Bmoxa
8I+uUgMaDQpghdUqhKiKjng7BgaT6cM2afeqJHcIZEM8OUwt65COPvs5oeA6mUYDh+iVLUOS7kte
qZpyujw8gxDTamxebXZYJeLYrSu8KguGsbS5qKNVQEJaLTqUstE3Dh0wFn1m6+LQSMiMXrhoo263
IrtEh00DkDi7rBj0WTSnP4XJN0Tg5f3qY2uVnQ0BHPJ/eR11hmlI32PS2EFUQbcehwYXEO5mEaG8
ulkK2m/+f7H5p34MbhQ7iYsGItM3c3+zT5fjbKNjNZhwgdQlAOrFgVk8i70O6wvZREc3+yHn/OZx
+bjnn8mBcQIQnZ2f3DzSpixsQRmpDiy0PTrb4Hv1ua8W50UaQbxj0mNEItm1G09eMuFN/h1dV0lw
47lsr1iIkoJbrMvTYzbea9su7bBxdIKxecxKNjlsod+vOvDpwU6cwbThgCKFZaFKcmLJP1nJCZPR
jLvB+T6zM0xxhdk0GG3Cabeae7G8vj1sso9oxTI/CCPNl5La4EkktECJhiGuyxk1FthDRqQjxJBX
lxCPPwzjYao0h8Dd70VYt+Ps0g3v26Vkd7y72B37VfSq7gW7hY70Y6lTmyZ9l3LH6BY3exReyuu3
Niv7FxVjJRmNb5waF5TkVDYeA1k3GIFrvcRkkCUTbIHC22afMsnJevIIcP7Fq4U+kry9YVRQ5bmn
JkdUNfVC8rWkwo8fLlnXNuCHpBeAMwvx4lxrHpuZhAwUbBavtnN2pngHg7abfSXcUClWN0z1a9wQ
YTY+rg4U53VjRtnZWPy/IPLzuNF/m0zI5du+WAGfjNih9VaGn8wjHySnCxTDI3urw251k3TuG3nm
Xz/zX135Yd6tBAQFt+mCV1SIGGtmr4uv4GBYL6BNzH4y2RiNPCrnuiP937q+CmZZ83GzN8fB76xd
3Evv7KBJK8xcIJ130RUtwNPW9pYhV/oMFAx9xbbvWvMPaFMQAISRzGFT8vt+Aj8T7+tEjwsmdpl4
ssyThA/B68Bb0br9UQymHuf1Im9yY0BdIduz6hzNfxrV5XIx9huW4sA7dUm9GtlBmrHFP1Cg2dTq
Yfcm5obfrYNg/B5NE67BRE2MtCXmUseu2z/76e3lT6W0wDihao45q+fCDbBERfkSS2wC244CgPCR
yVanFEWhndMdfIjZKlohhZgkWlBka+r4VlX6VTLcCgB/nHDYCRJf3N1m7jy+8EMsdjkMOaVocEnY
N/9/sVBD/oeSVg834bec4uklj7vzsf2AT56nFlHpEB24wjgsagZiYQ16VHik67woNnP9sIeWmgrt
RMonAOJVUzLFla7GhpzZyACanLP07Xn3oDP3J+xyLy9MXAAdN7mfR7ipHP4/FDC30LtkMm25U+Mc
SHVd8b74B++2ENnr5xcqdzG6ZaSRN0Ru32e8BAxQANNyJ2XJoeXh8U006OUTra/xYkenlBcekn9F
IiXpGtsXDgcUqwLZZO8uym+zqo96/9gW6QxTbvjh7q1nK5dIeLBM+uL6dyW74s+dr1pr7vVGrcFI
EEvvIknuXrCnNAPKQeRXLRd+f9YY5Dg4oht4v22nYETIhHmLcnAfQCP1y+iNqvDj1XhnEcge1R9b
QfxN1zksRoe103+A43hJwl+SBkfgBIabv/iyD4I+rLzLUGoB6H2WuoHM0MBHlH1KrPwnSGj1Bd49
FxPwjQTaH0QqyQYIURsVjBwLWgFSflhSeYt6z3fxvGtVf6Elw/hXQD8r0WnXQ8rZ8lMpfxEaBApF
fX9SKqg2TEVwqU0FymINKQwLyiiUIrIBqoCYoB6qtkimra14wU/U8jO+iHbQHOWaZldPAuWtIlC9
XZfQv2RgWiXCK34OJsd2wS1vzk4hdDgqL93mqWabLOA/KfV8Mwhhu1F9BiLIjcHLmXgh7Vxfnq0J
Key7JH6UADyQ2NmwAQ7s02QJytEYpA+5f5gF2TmPFm2SVQEMposeI2nOB8YtQ89IvRFO/YJR2Ub5
1C9L79vhfTVBLVyKfxIgUwMjezWXKAHYFblFx9NyRVbqbELnCR70jod+CKm+JKwSkRvndneeBnzD
jaZLGY7x/nBqJUpmaGviPJdd286UY94u34ckUEPPnpEMWovREZlE8ZJQ4tOLazkHmQsGcNCfv0wc
tB1JGvd9BUqBqLdwqEwxsvBZDzsVjj1Gn5r8OWAFXhhlvyKDj91kcNAsU4tHgMn6gpge8ApBczGm
nEAIQ848ZsfpOOZzp1kBYB26Slrw97NWPjxG5sXZfErId696OduN8sb1hVNAUaKToYJ66YkvQ4Yt
Wk/XVXEmCNOdWdx445ftk16sJHkQcMLP1sJrx6Ioo7+j+K0ysiPSUNJDfqjSPOgkybXJlHHhLdcQ
I+SdkRZhZ6cUyX8TdF4JEoAMFnvHbFlu8HP8+609mkHJW4JFfsX8mANlQQwCWHdI1OweAmWXL8ry
PQnAq9hS3OHL2yut00Sp8E/WHmG7chwW9gXLxssA6I3NZr6n1SQ22DJVzXMRwPtiYfdCtFWWsG/R
Xo10wkwViEygamjNT0lySMQ9uky0ximPBFoLSSFKHLIup1RgtpOdGGsSRxTUq1cFDA6ClZ1vjkxV
WtOxLbeiL8qyNPw6DVM2ipazjYR6SSzVEIDXCZgEiglwy1r3FEsTiOc5ZG6Con/ONuWumfFUhIln
3kcAzPiJMHIgvWZ/mCV/ik+7iakwrdrd8wjw0El8PBceBJxlVK7rFRNc+lKdQSURXiag+rnYlEaJ
03edZYoaP7sFpVkUjnTtJz3q0miEUyQmaGUWB5KVP6mnHOwd5a6IwBeV195FLnM36AkuQ3heNrBY
eFQqzxU96OaYT+gFlqyuxaPQ9fxQj1fAse9pn11HDCX7V68izPbb3XUWzlZRAJRxjPuLABQWYKno
UV/e/koE48/VUvvG7JaLlM9FQmPB3L23Hh2aTizeU70VhJiKjWsaEdk4bTddNMLY00jtuU6+/IZL
Nmz2NEAHusMsBPrOZ/mQwQCMq+6K6bYtOudD7Vizang3fPjznfyLm4FwR/1cfyw161htbXDskPpt
aJUroB5m1UIEBe0gyWNSbFvgssYcdu6CGw8RfCjC71PrtrjCzidlmfp9c5gff1n69gYYC+tMbBZB
n11NMPiPoQYUuZNd67I5ZcFoNO36+M5rci1qy46iH1bRpH0BU/JFIjS9Iqu4nBpyURIoI6iZIMdS
6LyUpd/WTY8b+1vOdbfvNvNodxmG9PkZR4r47OeNU/0GWkKNfSN8HSfox5uIZJpyGAvsUmc5/HIn
Sb2jmR74M42qq/IXUCS9NAvqq12wl9bYmbyCdo+Kt+u/mZ+LSU82J/d+NVeFY4sS+i0M4I1R4dRF
TmhyHYsJmLqEE3xAEmd2BF3TtEPTv/HmkVU9beMQV8ImlahDgCyVjK4+mbV28XyK2e/000CDUVuy
ylBTtIJrunm+7vh212cxn1kgtOmBNnQSXQ2X7AHlPfEjT4ewn+JwvRim7XYMEcUuiuS0Gm99UXlA
0RpE9BdQ2P8fsAp5lXnkBaR41vRisxwOX3UuAHaxNT4NiF+AtkD53VRJP31LAnJWnTb0uRui0/Ou
DP36suX/Wk06vkduccy1sS58c8qjNtkUAmDFpUrTfo5pekkaHhpd+msTaPqHaZKhb/+yBQ1PPhzx
yJy0iD0VPSMuTNK+ZTxRjeS95HtoO6cSZE6zn28s2vfHtSLxVYx8Kz/AUFbRC4IIfalMM7lRoNt6
W6Ngqy8R6/Abcm0phrU75ZHJ7k65O7sacPq0gHb0HpcN5l1lxp/NHfxyr1ukYDUb4h34tC6ZKENQ
O5rEsF1PRJWXXQ1v0q4LDc0cwcuOJ9DO0R0UiwMLXvsTS0iI/eSs9lBn1l7/YjQzdKt7w2h6N/Os
MHbAx3XUXZUnMipFNhaNN+btWi6pkM9BNPk5lki9vLo9oy7gcp5Ha0VNrVR+U+ouVblLQYg+csYn
0dtjAph0cNLUBtiDLZ2YSV5G4GHfcpUJBY/TRsV/eXwYmlDV+kWNPdZJnoP0kLlGOUvZtLP8Eljo
ONa7N8/mF7efiJaV80pb5qf+0hXjcUwH2Yplsb5PWAxI7iMyp3EMnpgG5dRDcceJAFlnFpDbShSx
CHM5t+eKxtzkw/65r1rqjVE5THPIpuX5eoH39nmqzpdO3k2gmGWr287vW155PKX8hH20W5DQ5vUs
jndc17I1650tW8dIKo2JkmAQbPNQpoMgWKqBDMkSqvgacXgXt4JmnaQaoD6Y8eXlCaQRJj3y7rI5
ASA3PK3rbgf2iDyt63MCssZQsWtiJZZMGQkabWd0YrYzwz+5JT4URrgNdVDnv3SDifbyLoGaaGYO
NuOfH2fnJNWMPbQ831opFrqJVyYTft3SR4cKu35DUtft9SbdCCWoKpasRXx8J0LJQoiOSHywfdD2
JIAH0pIB0Dx40MiWT0T6GDjPA9JoBmhGT1wYYSSFPGxGQjw4xF+xkLbDeiDg262pLonAsqb/+RxB
9v33Pb5Pd/j378rJ7OcfwGuUsxwFk2LY92HYZzsejxLJcss1wPJ2z8ikKbX/Md1m9iinxRL9eo23
xiTqhgPTuAMydd7nuMCxJeljpuLOTYfJ82s0wT4IsY/5qrvyo/teUnyAYeZyfWKzvyO+v/X8LD+p
625lLOCPBeEwxoOCzlwIyMP7Ro1Vk4FskXD7/FfO48JX7Fnf6mRlxcXXZGKFeT7kK1a7Yy/JdyHH
eGc5j9hkEiiHdYj7bPesvGJPzpFwmMcI6sjNSeB3ieIKZURGTt/GG35AnTNRCN7Jo3qGKedszEG1
n8sQheWU7WIfh0ZmQpdIhUz47+B/1KAMLllTkE1Epn0CYNKaK8m3zVXMtI4HsiGrKGyW7l+jydls
u2O6r2t8DHiAA6JNePU7a5XrGN7SNcDQuX050MTkNEw21GPxFs2NQJCfH464Put94fCd+jWHdPIw
i5FhOYynxZxH+dyuRQqG3NgmRNm9YNNztR81MPr5cFrjHc7iCvYb65WeE7++5/8yVahkauSYwApE
y1odOLSIMe51ZZCSiXNSuTZXzGuc/C8K5sjZYQdPm9V6lalDF3fO4srA1nv4rcJyYPTu8Ozk/3GV
BsuaPUMzPwB5C47qVT5j3X8jY4qXiGVanT2v/pu8MXk1ulJGMQ80Uqi1Gb8ipM0U9y4x7rYPQ2eV
Vv7lFU9My4p619rVBoKc2ehYvB/Eye2USx2E2obFN5wTv/fc4NApY7203IdBI7R90Dnu2FbG3evZ
Kk6Bt5ttVZqDomq7MeBs0n+tXb9CKHBo47ivi4YaZbGDFHOQfSCdBOrcEcGURzMqAlhsErg21h8W
FDEcJKVP24vNdZqLmB4tm2BXhsiGWA/E6LxzPpnAAyPLQN+9j0Ei9appx1TI9t/sb3kZhglETX2h
JgYmH1dzK9ZKz2hbkKR1nQGAPmxldutWGrlsrSvlOUyu9YkZkjuuaD+tJ+IhECHhxpkZyUPazNqv
4le3tNDTwhYTCg9XMXBLZ7cfM9Lbz83bVJl2um5eGsSAegDAXM+MXgjoul0MUR8/qs/apVHwmAou
1JLzQ/iP+/cpPNHWqNGaFcjhsDXE1Kt3qLz5oeQMbo/fMeRqJiCEGF34g2q+3yiD8/TnmE9WB+CE
BvlvMhaHd1hRfeEfEaWVjt52E5ltSNF4GSVFftrpS6aynDiMCFsYSM5jTLYi7Sw91BdIo0Pdj0Sf
dU7t5YvIZQ11xEja8YuTYblUZtUcTDD+DG9isrtfn/o9wD5wZbnlByETDgLSajnl5nCJP/8z9b02
RTq+hvq6LjSgsr6pHjSWZJtN4+F40ptzUx6SF0s8p3/6h3bygUmMKYXOz82Y7EkL8rNw+clEOdcG
w1xaI5lV27rX0nZq1PchxhdBxmouRAuSijQtLLmbsyxlzzJiCAzZQJ/Nihpv4nVCL3qyo7Fl3WFE
IQeS3uag7Q8nRoo0AfOLzEwyUV198ybcrSJpJWgxyeiPthA2gRwbrf1IshvF2lIZo4mKCtr+wkuX
APjlO7UWfuYOglMOhZDWAvc0Uv3MbxaBP25chjFSUA3Ai7cDNkqnrwf3P/WonzdJsjGMjvHVJrBZ
rEQA4scD3ZPYoJ2nrr/ktiExxMlfShS8rIJ9KnthAZAZjMSTQA4CcSEJcPf+hSfBLfMikxXuFGnH
9aHYynE5PvTKJttfdSSwcn1A7L58MXgLsTbOo0OSZk85X6CU4hCHBrQba4bSPbJdn0UxymFJCg8t
E+Sox75AAyi8MBwtRyt2enGkzSeRMFRrJ/wDr4df5JLedCual7tFy+mwXPjpXcldagRefmgC0pY9
L4xg/dK4hYAJEUOZ/mi24+oRN8wDBbWvFC+ridzUn62S9pxrWmVIvOm3lldm2FXN6yJ29w8KZt+I
YKvlW7ZgJUPmmdaA44+VFmpqRDR9gZVKNP5PHs/PP7hwZx7jmRGZI9CWnWVABHVJSLawmhKnFkFi
BVZL1hyLThoYOY/bc+fL9/x3DTTHDc7//14m6nGUnSdSPRmMeqJZcPT2aoXWKTy4Q9lPMUdqVRq6
E+DwTB8ooYEgg7La/np0YOBfluxrO2S2ZWPNh6tyqzYcV3H5mXwmGCgggAfyrt6+hTbTTytI022g
urIwoytiR8CJOEHpUm56pEVSxb2s2cmPLGcjBML95hw42CNsXz7chZ8Scv1DZudYPsSOXWnR9StU
MY3tKxFaTuhIrLuqXufPZo/JWMo+UTp+/4a7sBl+gZE7kDkjSDRbJ/gh5X1szPbaJMBo9uQHqM3/
3fGToBmcAn5v79zlmJNIdCnPAT+pkmy6+1mEab86WRg6wBRw3uMTafSurgFTYNWY/33EfyYMztPo
BLtvZmUQ2JasV44HDiX/PlH0beowwFCRxbNg1DwnSP7giqLimWNZEpHkZ0AmWCZaNC9mYmsi7qyk
AWJsi4j9qUdJ9vESaTs/6bXozb9X+Pls3zOczTrd2gYJMl/vF96hmVyi5K7zbbvjP2nlueSCnm6z
e2GCRMSaORRVMRE5o8alsI+LZZ/f9xSwB03YAZ/pfyRuTtUSZQp7EeIUP9KtxBXjpSS9j0Gdxkd2
8lohq+573Au6k77p2k+eFQ2Mpr2dPjJyudUliNLZB5/xvZQV4FTS1IlzCnn8MeAD/3S3x/MqLq4L
Rlyc57ejyf/Vblk4/uFgwiE42ShIovT+GHdO13E/w+4eGwJg4gZNWRYponkWo/P7vvxMvsUMH5dg
Q/n9Wkcmw/qaZ76okBFhnVyOOYhMDW+NaFdE3QxA2TJjm7BOKE9iVILjn9S9CWf3lildsJ0HIBdw
W2I/JWZ4yzPZLtO0ApW4AF9uOI/MWbI1nHpWuEhzpkke+ljvyv93BCccrjwh5G+1oNOrgrXAtcgi
W2IzKDfLCRBUJQS3ZURdQuj6AU43kMjmXzclMfgC0u6PUZQV7E4oG2Z5aWKmd6Wic9WJSVq7e+up
Ix3FOHvjNcGc7GPJwaSCZg34vSLlIFujt9k6n2PnzBZM31NnI1oufEboR9OAbPNgmmmwX9ZFnu17
bHZOUh9xOJGF7booLlmAibEZ4K4Kdzlgw5aWO9zXtXurjJigvf98yJUsjKmX03YGlAQKUfHkY78y
16xfFd127Jvgbqwr1YJ91gCRa6HjeKF0t2ZW1Sw9t52+PEyOkFKirid1Z9gtzG3wUxAcd4m8CKpt
myO2vpo7xG/ECBwRRFTdl4uzvtxr/jxjEIIHFzLBqG9jWtavKFIqGDnfWirFaPAGbMzxZ84/olUZ
Db40nRgL0+s8is6aNVX8BKP8f3kE5kv0lygaosYfIlRp3sFoY2E+KgHapyfGg2KduXg9Se++mc/b
c4PjhsiaW0XlMVJ7pWYDB7ud6V6MGB8DMzcHGGA5Kz1dd55PNYIAn4Onz7urj2ZjsN7LWtRJc62C
vJ/n2fhUGL1c6hWRY2X5q9JEUN/tLgmQtpTzMDqQi0/yTQN9nhQPLNBUQoawV67lTjRRgvgBhocY
8atHckFWm4O3VWtc6JeIsCNUZNYZsouSjoWm8Lat/GN7oP5MdsUuDpNLftoCJXGIMX6jC1Herolq
eGYwTdI/PCcHC9wXPQKrNF4Zb3r9ooVaN95NRWvqk/TNtQz2u2kjDYzRn+anZOA/kY8vUIQ14WpU
13ZC4s4cAO6mxn/Q47tWQePMshlwJo2VlnhNQ/e4dOXXvmzO8fq4ND2n1yORGgKZQASQ4D/QAZnJ
GZ71GG1GFq/KuY+kFIfSsBbxaBKwZto7PiHkGOfbPdf/hb9UK+vGQWqUBW9lM9mxBko2vCLH6xZX
zbzV3Wtu5nIGhbRmEigyiQu6L2J0dSqi2dWmO67m0mrEhNn5BIDrmKjjwvtS8Fy7gKCjTwK08/td
Dj0OZqVmfoWP72DMc+Z26oXgt5XuNTW8Dp6P7kuLXKqJ752kaoIht+T19a0vpoR2p5a1CmYB88na
No6ipu7hHJzGFN79fiIrxzo80FLKNifFNYDw0PdD4Mh4dWNNYsMHBn+Em9nmFytZnd7Cw5206EzP
Cg5n21bHT8fgbp0gcQhDVK0TAlOEu6RZA9Rm0On76kDospjWUuYjk7JQbV90OCPEC6u1MrmY4pod
tpjSxq6VRU3OT6M1dsQluwCM2NnyvLEx0YDfcEMXLZfcyoppQp38vmEfwuew1t3rDHoW7ObJAS3u
JLbxd7gOrfrV8xZUuC0XOLa24mqvLGeNLvGAuICbFru1Lp0J/81ur+/KcMwkreVXLp6hsrYd54tw
sDtGhsv25b0hwd1kY4uo+GoTzMvFjZxPN9+njDnbsu0umTXANfrRxT6Dc9IH5DqPPhziV29yHSdv
H0E3sfB4JtDPMLWwPJB2DrMhC1D0/CgNMZn5bsnShJ1wFfM411D2uHhsWdKuhXPiYO4IzjluYS33
78rh20MUnsorRq2xFiZcxT0/Ikw77Y90Y+q7jirtKYSsCiy4MpOYx/9yioFEHrVE1l62LxpL4EV1
nkBfuKISlc5bkyILnTwNhRJ04PZ4+YmygnlCK3Y/ktLBrKFYUIEHx60ChilvWfXcZbtUOjYGZycf
gwi/eSxpvmPR5K8JEa7NoG/9rrCAbwdzKLdxZOUlOZbdw3ZmlpgCPhhA4E2Vhe65bg4WxKSbtLps
lXgKqyer+r1hnTwg0rz/CcbtF/KscNNK0qxElzm6GbTC1c49GR+jssgVHdL8aDlJ+k+zYK4Pc0id
ftdgUXU0mLBSAStIHFMFe76tBSF7YDZ4yjehBApCuAdIjpItasZlkZS521K8TkZghicE6CbJ8X4R
HN2dDxfjm3Dx/IskWmI6Zl4Q7jZ/fNKYiIhbOMePBWgydbul0f+6SiR9qS+HJU357/F4KL/9bIXD
Q4BFLVVR7XWMK8gkQdeK7SZSNdDeq6L4RPdZvbytuDeYfvVnaGb0ZW0gSZa2c8k0qHj5k8kMn0r/
jenpQVPHVWRwPVYCKJ/emJtOG/na83397XYFuEgE7GqBrdUTHR0iWfwWa3ZIlK9tKsf26P7lntPq
xFVJ1PCm0y+V8QqxeRmMPbAAbc6UiqEPHh2wTGhrii1Nou9DK2wo8huyK2DR3hJgk3QNxv2RkEoz
Fxp0L2xJdyGEGvf5S8ayGS4s2vn8FARz0KvKv3mymEePcONeEJpBygjb/2kz52MKzllS6Pa14FJy
MUN60JW2V3yGdS7lELKDWfostYX904itSFV2H5nS9exkmTyGD2S8j8twbWy/fylsI8/glxJyyS4M
q4dizZ09HZaIGWgXAAqyoH2BPzaCObAB6v5eQguOu4/6h7j9L7w04TO4/lPoV+pOgon+J1KN39se
Db0kt0GKGtqM0KyhwDVYand/1WaaAvtEcIxHp5WdMHnUnZ3x1NzhpmbGUrhdcB6AmK+DvpHAjKaO
b+9AojUrMtttnFPLV6bFn7vGn58zcsqkIyRfVUzisNmG41DdxeynZv0mSIhqBfTLzrMtUdCQ2ID0
Fh7rhZAWVdHLzviPebXRKdyhoLfDbloE49s9wVwxO9p9NBY5kl8SlTkZJhdtyNs9art8kZ7caXL2
TebkR4BYWhsEXPaYybD08eyCGF9Ha/hp4kHpf4PGnBJc+RSE5oIIKMgJZfXhYDvs4jnah44l2Wf6
t+YvxBHVwChWMcavqQkRhpRkG/n2iOgbRx7X3qK0MT1CHdg+UuI7ve7cBVUo0kz7A9ocWhcAeRQo
R7Pi/lYtPif0Ym/lXrVV9knBf6QIKGlOW24EbdwQH2RXiBFRw5jPhydDEOIlpqqunQ4sFCSaWBL0
LOnj5p6eohT3MGxQoZ4FTrTvzWylHSHAWxByYXBBYnnBbjLEnG/DIqhMYqolHltPbB0ERz9QVmWq
P//BuPyTZWikCak2s9A3yLtfjNSDGB4UDi6/xqk80uV6J0uRPuLoqPYMFkbBCByxxMr1Nn1Glgj2
D6k8ueREOOhklwGAoT86MZ/3Kzbf1174ZcCRDTKT3HBpZqBzgdmI25cS31orLKfa5csCm2i7fNHx
tscqWShGRWHcKM2cRB5s294Jl9DknDEViTjryiKD8ztA3eUFmb6kspmP9dDeNoKVR2UPR9hqKDmv
MdTl75fDx5yNnGjYHRN8fYJj4bcYSvTMVgAtNlJckd/qnwkMcgsNEeF763uckc9yjEBOXw9lx/X4
rXRnI0tShMj2dfomOxvFgRQJLOEt6HG6xr+pPG0bZ7Zi5rc0Cz1Kb+X83PFaU/yxJyNIq+6srlbb
Qx2HeFQG3UHFGXslTX048ddrKnRsR9x5TC4ptWOflHeTnd4YPxSjIDmc4WcECYabHr8IEx4L3AQW
VnAW+1pbsF1NnGyl9pwwHxm8LHqFmKxJTINOBSCjx1IZINd0v5C7VkH0xkuazUWVxy5E7bZQrQFW
ekHj9CwuPuBzxEEwSqg3Xjvyg7VZgB4+SqfA0kYPVc8ojAq1946HFTehgDRzwwXoTfVhKNSWuPdv
QGmTlrk5aWD43c5OM/HcGAIGV65jxh+9pDPAgRTzNAGobbxH0uK23wRXkVrr18pxxCoPkzWla6i9
ZBznTi8diblT7JxfxcRzN2egbXJ5fwq2QGUO2dnwK0Aqk8Vb8wdiA3Qd6X5ZzHMZsZ0WmKiNlbv3
RntEDD4ZEP63qyxvJ5+QSbuiYyCgb0KH9EOxd5i7BJ+EpjsxEam96lcQytS+e41PCh9hwEhijfar
Q7wB4VmX8MW0s1Bh+2XyM9aXPo6nwSCksZYV4bgsuhAtuewX/36zChepoV4/0fp+Z7o8f0C16BpE
tci98z/veAlKJKwppOdTuVoQMoEW7v1NckIWIR5m5HYuyBz1aMCXo9B1C2oofvPSN0IMa7sam9vF
EcxhLCKHg4ndB4ZxbabFloCrQpUujaX9AVACdFRxhgqg/i/YealMpb9tNSMTpFKfwLQx1VajFoJ4
d1FCATWSvMPKtnbRIx5bEOIP6+17AL2HfBcGGB2w869CfpfaOutPMVRcwKWBC7Zpq2AD2dHP005j
y5xpCuzVObM6TNpq/0iCBRW51qfoUpp7nt2NZ7vvyd3a0penjH+eT6kup7RFYnxImJWMAxMZ+msG
U5cq8HM/lhFjL6ARc8Ye2pj0A804QN7AV6gSzr3ljy4klJMoWFvPHJNgJz3BcVoNcRX37KIccGPu
920TlbYDW8CmbCGSa87qABMgaIU8l6tpP0KLJFigCxu+LvZhdujLlQzZSXNL7Cxk2FpVye9YQTzj
MImTid9vMeYLTVGNf0Dh+bU+r7OMVRjFMRRnEzbfti6gqV6D3Ec5CJLF7gyAKA2Lw979PLOlWVo5
Ldo6roRVHYcIM6Zxbgc7ZnUSZr9I6rC5pmFNzSube71lSqn/R9gB2iNySkRERHPvPVlUMx7Qr3TI
zO9l4shXmdxeNTfB9meqjjxdsmMxPtazZV/N06Hw0EarxHt41noFO7YwfAdNiZ4jbCQvPNcobmyY
pN1x/zEjPx4oFtxuUuO7pnqvQdLKx/gkT7m3Kz7JC7+kiecNEajVkuXtFnpbKOG+wjhFhgrZOhlP
mfDjAATPI10DsMhTYQm1+EPIFrftpI17G5sg6/hUTZKf5ZT5F4rzWX6E94IcbB2yuJMVyYp2v9EE
KWEXEejegobbBvDK6myvumCJUkSKMLs759HbINJLzlbRoSltDCZNkAzPre1ZS+5S0QlSF/R5XmlW
q3jn6Kgfiuw5umeUj8ao8LFZdqA6EB/BJCX9Lu9PA1PR7mjeNMmEGF2rgzNd1bwsLflV3gJp1c03
0ufG8xsldn+OsXwDtUNz/5ZOBhN192+eO431ZU8dc24X+ZQvVasNYRf4gj22PKLNNDIUmoGzIXz4
Wezq+Tdk0wtuWZamZGpLbB+yl8WebaM6bqEFswgIl9NVqSAdmSFVXeXSU5OWBa7XzYcIAtRjaN6F
PoGziBy5wwt4Atvt3UsXBR3DC/u57+VHja3kBD6KjO9Mrl1caXm+jEMw+hNZ3jug3kmLU3rwWLqn
v0O3L45lYtHeU5/wYv38PnEATk2w3M/pCx5DnzVBw1nDcGtTFl6aeipDZD9Q1x2LbuqG6DBP6okl
7AdzU0cxzsWpDCz0DiYjlBwtX2180UHloPTx+lBNwDEFtrC0Pay7CgrORoYAWjvQcoRdGfkoC9Uy
X5GtvgW2819SmU9jh4zF3nGYR9ayav5TOxdQNAphzch0CqX6V7PlcqZcL5aUOrZRjsBf1LTT1wd/
dlvBAid2XxWj2kx/NKFRiltD+jqPJSFhPabVUp47izPeFahmii+3oDxLlgbv1QTXBmQKUXkwBfe2
EbxlJB6oHXXF46SAJbAZnyLpCGMWppeODDkZymAPaenCh2TeAIKSHGJHWQM2EvntUPZMTXfXGzDM
VkVT3xY45E5y+DQm3BzhNY9ruzG6trqYBS1HXHiZ7DUZMa1YzpCurs5/Ofafrpk+I9ot+byeB1wJ
j22XT2HKNo8ZBhNleLB4iza3GbekOWdVQFG06ys7u/KdE+bZFyOi8hhhpOEEt6xF885EODJYD0Wm
SAutfH6XWDNXtxMCp2BE52nDPQ+WTXqotnHXP21+EMv8DKSwV9hRneTqb1tb5/X2E4gixUZJnOs2
FkNIiDHTBSH4kcUeNnVFXemX+BhTmNIz1QAv3mfCCimIkaTtflhsgOQ=
`pragma protect end_protected
