// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
VO5LX1FHDWth0KB0WcJ2y5HCTagLorNwVFNMiagLYiiiIXhPifqUjwo5r3F+ulfbkEEAh4pbaAvu
OEUiGCBBGTcEOp3vRVxwlhDAOkbfUNoXNJZZsmHM7jKuAgshv+JDwO7Aar3NTfJRS8oVOal0rfqN
yVo4Wi7d43Tlx7gqFlFGUQaGcfn5zuLiXC9jDJ1sxjKhKIxsnpH2JrXskA6VT1pPQsbwrys4TFll
SZX36l/ktRghejADGdH6pvkzb4CULSBq6O2ZPUXtfvWkMCQbqh3pM5o+BRlFdfMHnvcYwkAJmZ8s
JtK1f7br87zGi4gIdakbWNYW6Da9yciX+Bv3Jg==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
8hQNisUpTXpC7PbMudH+NyrgFHBRccb9Ffz2mpW+UlWbksjUSw0/HBjBL2qlEDxWPGUNvEqfojW5
4sG47BWe4Yom8UE41mizuBu/9xys9nffMS2j5cmkhlNj2RgLHVvcsHm8idrtYNYiWG4HupFEaZVM
uGa0KKLvkAccAHll0Q78LPExqEZuY+4O1J0ycHl8zxzko984u28BWJPdKUolL2LLRUKOz+B6xt2D
Eo3DLyUqJx1KLVlqP9f4yZuSSEoipWbWYEYUMGLszROZ9jKB0Sb8d9XKcsVKvZbHOH/5pwvaXD5w
GNYc/XiRIVB7eGE3k95+F0nzFUlJbeV/CKg7KMJfRbkpVPjnnOsUZzywAsrj9sYDHmVZE5LzejgQ
EEhlOnOUj65C0O9SFDGpAQGGLr685BiKFenXH48FbTRW73FFO1jxiO/BGG6+ZFO1e6BdjRgxi9vT
Ah/HZYC2UPdPTWcMKYryfBxrbAT/jb2MDsOlqem7PMHQRjiQTx/vU/Inx7sgObDI/agzdp2s3r9r
/vQ/mNu4OhIH6DfBXITkLul/JZ9ntVS4C8QLELPDScmPUheSJK3jkzi93ljIMGjjqGC4+Y9xug4R
T+pKYKOxNL2Jq1csBEgWc5HKv1O2LPYu+9HY1bXv6SChMJq6uZfzY1nUd1EprrW1FyKsasyRkTww
dq2tkHZCv4K+3g1IW8+QqgkSarTbMqwuXhpNnNud5iyM8zNChkbRgSCALJ3EYFoW01vN+oeeNpwY
Qd9jeQRTkXXBuRMHo1IOP91fNWjEjcqa2E/qqg+kMuQo6VTnszRctXWQtn3sFC1piJ7UdKv7Zgp3
pOi+vMd2GnWvu2zeCZ7who+kKLd06uwDf7IX3bi6BBacP3BjRU/5t/EI0bMxwbZ2bieRE/VPa3vM
VuE+s5WMHPVA6gUhZkdZK7iYRj8s8zs5DELzQTXB0YIcbCpSkHsHwm4ptqt0cUgKXO1irxKvCsLV
9JmV2nk+tG2ZhqnWvl2LuzgAPFtjIrnXBZ8c8FK9xlU0/2TKvepZBGimoIkx/NKwXeGypsq2jUHf
P+hZCvMUF7BI+Jy10n0nxt4F6ZYOP8pCKOSnVldELvu1OiNYF4N8eUGLlX6A/90JCqMqbYk9nhEe
c7McCob9aoJcqb8ngFTaX5n94RTkF9jmmDjxC6W3KToxWkiLxk1HeYHToFeHEcjvHV0gNno+eBKf
nquEuzkTUE0SDguEitUvEGBQBdrpuujrIagx+Hz6VXCiZUQTPH/e7LJAWjXUxzeO9u7ZmQ/EDq4l
WnYOTx//mJcK1quHyzgWZoesdT8eRhWIiETRUMgoJQCmOekqb8skcTkpgkJ7z1n5B6yqBqW+hzg+
JPIvqGElIbqJoIfQcjoHQEN9uaGp6eaSP7X9w2UUOGnWt1RigRyBPCxpeYv2FDRVKO45mFsAwEVV
xUc33nki6Qu85wxVrnoV9eJ8t6dii4ZXX15RnnnsYtDf+X1ax3VvzDJAjYq4qQffh6huzmYG9k0d
ax3EMtZhGhqBXJ/fJnM8BKyzym7TVvMIavNynMMU1+5BcRees8kxBDo2A2BuTn/akCTvlXlCmpAw
SgCA9fZUfaY6hi+YytPGzSjNBmVYeMEFvp24eIPGTvoeoIZ8k0StRsuwsOSeOnrjKhR0Is5tzbf9
Om09X2cn39TEXp0ySqm1R3xj/PWXQsK62yH5PLS4bCh2Sq0wxc1o8Ob6vVnsr9WaYp9yRQKfr8sF
2KFETk3/2X9kByo5r+K7dKHZE+q9pPv5IXCei1stbxdwL5wCjshfYPFKBWI8qQvznxl87AtS6jfb
ZwvVJyAskfQe+qlc71UZ7Xm/9CnM5vFI5XguPPe+pyUfHQBmOQQMnYpdY0w+G984ULSO5u3t7kcL
7lw5HMsyvo8SIxyhATtQDBrByjV2fRa1mFLlXrIO16wbOyyLBC6SKR1PJ1Yjj26vC5XO8WInB7tD
vwYIzquosUWg76JD2dAUVxRqlre/x7IMS8Ltd/LwpZA8mXO8z4xSo3KrLxlC/z+Fny7qm2NYLWT7
7uxShmn3CV1dQwWy457lAwwHcOKy9KsF05S3Fe5fxrBH0aek5mXC5YDsbul3iy/ZpdAi6rjZc3+j
KgtJwPuBjD/q1QTxAfeenHk3J6yjbgJ/+E2P+TkOxiqunq/xflJLMwt2Vqq2UamH9s//wnWQuv89
unwkPVIcYPcCfjm0wpb3WrBeTVvp//czuLRcoMhbg2AcXsMy1Iv0QYB0LvHf8XbvBMAiMxSHsvJN
EdcHULMg5CfjaFAODcSQwnC9qtCDOZQDGtwTgzkL3+J2kyNDIE3jJUXnkjvlTEvwQYt1/3FoahIb
48oX1bR0X7jYuYpuuKgoEO60UZXcFXwOaHEiRBIxQSYI+/z6upeMqUOd16E2IVNIxYoSkU2oyywy
rcDmHgRuggzLT6L10inlsdhZ+nM+IwdWS4qzSs+EOF1ArDeorEsIiB2WD7yyGCVT4SdOecnypdn+
kVCJRiOkl+wvxTxuaoKDqN4gjYA9Ysu7wf5TvcApFX28Ya//Tie7IPUaX+CFu6D07yAg3CpHGcPO
Su7JL47qCHAzM8LH+nTFnx9LCThbbktwgm+MZiLX6JK6BK89cvdsTD8+QBdBd6i43FB1hNzRgSAu
FkMSgm2bWFfK25a6DQ74V13hHxjfl8mQ4PBzG7AD6AZ5l52KpE2nK9K5WJdv9qtNVCOcRMlZnx/m
bA0vq+YvpFo53dtXax0ONYM2etxjf97QGIJsVwv0qtPJWMt1gExhWNcn6oHNk2XG90+7ln1qQtGF
Y9vrpXFO2GCBFZYhXYRraUzBzHDGLugAjLpDCjCpnUqr8TaxbvCYn5N29f7nfr095H2smb8bHuMp
hYlxrLOd4iUaTjO39tmi/EkPIwMbBg8DGUcA3rXdzfHL7EaAMTfaC5fZFjwkQOkY2f7N0QLNWuw/
wtBk4YzeEogSeeNgyQrz90mMpm9jtPsYq1utx1u6q/9LSA5JcoVLXcaGASptQ8f07TqR2cg0PZL5
AGk3SOwCzJ3B5BSFL5yBBRJwmqpN7Angwdq0aifEPI9yCAQY/qf8QscGPD44Pj9Pdc01tF6Sz3/o
peF1eOl/2dEQ+TCmcXP+cb6f3YdkL5+mBWWuaStHT7O4GNYuTWpBsy6fydtDgmNRjp5ZvpGbDb2Q
6zO7R9OJQqPr0CGV3xM57e3NPys/KqCCXhdAEHfDz5Kg9EnES/xjXOJP278N+cUq1Enxunht8W8q
VBguRyEY9X0s1RHrWjgmftPLK4IUMNeHuhMQB9pqpxpnt1P7PSKba5rixi6VhmOmU0xE339sCq1D
DLp7+qJ/mqVg+htqYYgShY/795kGXKAIE2DVgKIctnr5ZqR40dlPqBzokP/ypBTuN5rCBjk8y0U5
eqSdD0OPgg3iM3eOP4cOkebRQuK5ZJH1ucOEZrmaASKfLz3HuuE8dzOqTdvBAHu0tpvrKi0DeDwC
T9rR4vNKNyEZcv4Bo+hp/5MZANGQ5vnmJa6yaCNifSRw4DbCYuvNv+oYKt9y2aC9nZxor4bFbobm
pZ/LXELGtQHLgNpDOOrKxIJVEyJcEgIgDzeQUCPgfpIROgZS3TUMNaovqhEux3hlq1oL0MdGZHtn
iv04ToicTS1aJhE/vgoJmcCRie5UfobgGeTV2Ki8sgR3AXr1V3iypWS0g/cRqbjIlnDXeg6FN8kj
1FvijLQfzPrL8/xBVYLHdT89V9b85I6mS/iOysfC/CCGQXUnhvIMElCRZ2l1QKyVZd/I67zHXecF
+afEuhgTF75vySkwUWOipWPNX6iOeCiLZUBw4e9WuqXbdLMSDqe7I6db0dolippuNAa3uAHrE/an
E/nGfdivDhMwpBqP4bnKN0B4VCZnNKZLdX/TClBgz16boBYOV1EKpXT9uXqeU7zP1ZU1HQyyrvH5
ZrFRKvbZnubD3byU4tkWRX6Q9/CwnoPsyescO8JhqXKuL9YZCdOlYubU6ACwbIfrMDXK3SNx/PnP
TFxH1J/UxKNq4qUgv4Q/hk6xHjSvu3keQP6BPFMEZEO6/6Wh/XJdObgyc9tDzJfXYoL8Bo0yxYAC
MAV3J0eKSzLAxvfKP/f3J3Bx6sduQF/NcwWpka1cRQciYYb+BoKsD6scJno/pl0s+gLICUnlrbDQ
6/rCjFRavV68F/Q9RT8wG8ufQsbUYNMWTpQXpLzndek9HIJxSSouEIhM5sy0cUSgKJ8g/s0CpnSk
t/PyJ3ZAQVkRRhio2lbMghPvRWPFq3p/N7pcTwq9bTxo6x7kVyJrcctBp8cxFkiEFPU4i0/xGJUq
/f7Uh35e9an5unZqSOIr4FlHQtXvE6pgl5LOLErSUUi6FJAcZLjPL1HXCZCP39Hnhyh9BmvJ/huV
S4Y01Q2KbxbardQHkXXxZFz/4Yt71VNDrHaz0nd2eB0JqJGsOddKV73guuT9wKEtVo4y7R5u4mEH
buj9vitNuBiXnacM37MZ++uXeK52NFsbR+xSxbYWYyDAwvEBYVeg1RuWxMVa+Fnm0RspiVz1W9pu
mb7ywx7lu8J2hPvG25wHSh7z6EiCzMgs69PvVBztEEGQrsuhDwEck4hhmg8DzVKnM/SpYwOiRIww
pHrckpuB0fEgrNyHdtgf7PvalIo2mDcYmyRcc+WzUHCCz5zF9yKzrH+hpd4jm8jLNxv6E76YFp5o
TObyNCkvHePLZXNYxdmKKRGR+63UgaJ+/ypuQE0ttq3PAHOYTcBgh1A8BwCl0TmEjzKO1T1ZZCS5
K9AWajxG/ajQ2OqDRyGChrtvCtv+a/cXHineKtrG1c5A4r3tVoOJLmpSJxIP//pJLfK5cQs0fWzD
Mn1wAQeS3e5VKOGLjxEe+OuUlCG0tQYTueiVctBxC8AiwMoYYBzapjzxi2Z3eFYv7hErAmxX5q9M
wSkmd+5+m+OKXLii5LqKAAwOI1ltAdNe7leFOc8JKOAcv0dk86v6i9iE3vy69O6j9F7Bx5qSCUTy
kP2zG4u2UdqKhkO8LGfXgg/0Ero4xhDIWJtyO24zwQK49VYoxpck1N226tAqmAGdx7SiRQFw00Lj
MxpM+rsUMxhKb4ViShqZGmFHna585Oh27Zl3Ojju9QPO28HTFyJuCAuuTbs/N1vmGTeieU3VRhbd
Zx+UKcIm4xBbAvl44QhlvWJWmm8KAyyLyDjX2XdAU9IN1HAc81Y4a71ggRKZLgiSgAPYUl7geG/Q
Iq9/KDQZjKWVqyd/FdNdveDook13DC2+Q18vwpin+VcNGEhVUnEBswBBD9qtacg/mrD36bz6URkZ
4VZY6vB/ZyyqMZA185URFm2b0G+nYovvD7U6Qalcla6RTOKZqxmkcCE/ErRWUe38D9J3Ct8iCfKS
9TVpVdiL0WDb4EW3ipl7QHRsuloQUEBDqSbOt3tb59QpZzvn7z/uR2bACc9Ekf6XK7Y859mqCwpS
5lA/+u1RNnjxqznLWcT+ZFNibf1uqihlO0m4bgDbuo/nNQaNWq1zIbQcFZIbqQsL07vN7agGV/Va
giA8zwXFuact4qTzsWhrifRKSezJQWT0WmuuyzKZ2r+k7MKI/6X0rwrtVb+Cr6SdmR9Np/P4N58L
N2eqIWGYGIIHiqZ6rtIuvuY2mRoYdAcNQbu3SxEXfbq79WBU11xK056vR7dQlISzZswy+g71P4RA
m64E4oGWQObwbnL6wKgdG4NN4Va6VC8HlfZSCjxOc8GjLLjjZRmwasromOGjcJW+/YPIUvVBOpcK
9gPOd/1IFrorXdQ7EMbhnyQByEYsqzhAOrLE4NoIbuQ5/rPhwYfIi3nRYgG6Hjwp1lINKiPEKUyz
AMFspb/wgfHy9/eWx+MH73iEb5bdNmrn40xP03xcN4swyQ1cx85AG/KT01fCaAoWV0JSIcsDGQyi
jHFx21/6EgLpeSlkZnO7PSQCdMfx3XMfuLjUp186vg+Oem7yOVmNZkOwHiulxm1ltJ/IcEljB3H+
T2CpnPCPFa0swIs+ise3Gxt5ibjeclK3XDWucVt1Ex445Q47tHWJeDtjiP+HEEYR66wlqtvs0A8f
HA2ouVTRImcu5xaOTG7ypoOs+KwCBNjka0FtYIY4L60pq/m3qwHLQOME0Vy2faFAD7gcfGS7XQ3L
CwCOET46ZJOJ6vfheI5meqNE324MUeGBpUrm0tGGXBupBq+F3RNB6lZbss2FF0nlXSVON1ajAWSd
Qv7s6KG1w3Zl/5OxmMSz03AVUT35HeYoW3Y0fSfON2YtH6ju8XkbvayoTT/PTjtOF11addwp72FJ
d8A2uenXlAhUkHZqaU38fVJ4t9djFzUVYX6BgT/GXY9oYYfPdUrD+viDQkhpZNIYBjMDw+NlXAm8
ZhJIRP1cE81wk++lp+f6gZGLIGyZSjQJHGNeTv0Q5ljnow1aq8JNMgsrfbh/U/L9XlK4r/1d74ab
jTscGTKCA3pN/jsDibafALo3tacPvvL89iylPFSUEoMyD+2TJ2PL9oj4WfolkV8u7zXPrUG1HJGo
d7Cx+xYW6cwk8KKgH2IMh63yNpi22+F/cK9NNH9ydcC2HsfU10hLgG6BCQym4kSfvAwrWguNL5OW
/VvsmAX3FmhYooizLWnzXu/xSBfFSamBa4oPR7iYLHwWA/gVHVXd401+wTZ/tDWoWleyqyWYnx7u
ZQjTZTe8hCUHpUU1zeRdl5n7AAc+XRJUgKQXDYb559hR1oN72chmg2vYgzdtRcQwjEDx1sp9JgAE
s7nH+c/p4u/X+FqNxJcgSL5QhXu8NjHunftP++tFilzi/egKrFnHRAozaNRgUhxYJ6+J+/tDH4bk
q41mufv/1IPWQAfBPNj048hzB5ccyoni/sefeZdO2Fqjo6KBXInVW3VQhN9DWAxmzpfDt0SeUzQR
SyhjV3VHHgZFyXWJrprQq3bU0NKm+Iwb5r3YINjJHG2UuqQRalEKkwf/khY/6oQEkxEzQ4Lw7qGs
ImYKvujwXUx6zpzudt9UXpZ3C1ACfOaGF9K0cSUSZyjG3aWAIzbkygB4Eefz+ioPm4ZjB6a7BUGk
UBr7BxJdiZA+2auMafS+1JCC3bSjuno/zbVMHMF8wMNwl9YtJyZULq8wdT5LEgk7giGocXksV+R7
h/2YxjLiIdRn/jt+Z8KnFONLz4SqL222H0jxIB8V0VMpjzKtIWIHqlE2rJBwkZ0a5QAj106LDawo
tRdpa4N30Cp8uJY94enAyXXTdHKzt/umco3uLBClJxzjxV5tRPu0d40FR2crMywdFQ3vHnO3pFwT
1hRaNIewr5DTEWscr637ghIBfj473L46htWfb1ZKSH6QCp+7p3VzU1JwFPzpEn8b8GQqST60c6J1
5za1+T0LpgxWvmpAQQCVJWfkqERpf5eQvaXvxiCTtjo/TaF394pk1dTXKXiYdhs7wF9RgRod96bI
vr7Xij1VZ/+XW8T+FYOyRLVIk1DqnbGPfCCxlo0BufI6ZtIICzoUpPpSfjmIprqwvxhJVmbGjrbC
QnQbDJryv9CeV8XQmdSj1xTwfGdOCau9uAFmSBz0sV7uIS8JjUYeanEm6QpI5tzgx/lHzvnAEH1f
VmHoXQY2vD+ZnPQRfwXjT4IiWnBbsFVXtfLd6FiipCGUIWAufB31McCZS7Q4xzSEIonzO0ZITL2D
wrFNKE+C0ZsCEHQI5VbS2/KHWnU8HudFcdAaCO1UA/9A4/IMfZRjax6ifWgEN8d1IiuPBq7ifOWc
Pni8A6qotj9Bf3RZ91yRiqxH52PDCT+WaSEmDDFuDBjKcAz1n0MSXpG7bIPgEZ5w5PBfmryCSFv2
TXTmxHpvP9Oj9dSEVc78P/SaL9n4XT6+M+TwAHJrA4ZlsgE9GHacFrG6o00jkE0f9nPn6Kj/LypB
K+zgEsC4dwEXiMSH6tQVYi551mu+Vw1pq1JULwFBfeCEMIpbuOhEl0FYdInOw+k1kk8+GYEnTTTv
Cp4LvKrmVww3P3ojrIXZLwYhBELcKu9Wa1TwaHnkujNzVjrvEAwlpIN+AjiSTmUwMpT10RD3b6kB
gdj8AmNcSwSswZ8hz2yWjQ9gbHAIIzQaE7y/TxxsOL/A3ZhnKoK6biNjzF+UKTxUTUbSAh594dX0
ZS5SJVKAhu5UTowq+3IqI8dd9dNGYREOXdvw6ZFZFfJqNq1tOB3aL2cOweBHttssXQwmCJzuWtpx
K6hW7zR4YgvjXfFCjLa8+NGUkApJT9nfKemUhEv6NbmAcOh9BDw2AAuQjqig4XCOU7R4sICtny6d
KgdZJYDTCBfJrwSzkTQCDw3h6BywzrFeMD1ki87RXJZKAD1BbJ3VnuWUybZm242AbSOm1o6saicd
tvmMr9Uqz4g8hfCzmo7tsPG2b83b8O947TdUZxDfwAfd5zacoW6y+8z9D+LAJ8wojv5mtLXcKfKq
AXgG2KyDmPJrUr1/rgQLofv9mqCOXxbbPhRTjwnxf9j/M96VLldv3MGiO5CEEF2N5RTaFpOwzsQK
Dl2/QrXsy2TxNUf7KkTvgn0TLolv+y1DZNlm/arC42l/VpaddCaIVa1lG0DwWsbAMRAt1f66D9aF
29Vo2GspAimkKbiPZYrtJYSwl/ZQvL4PB40Rrh31V3LC8MSCA97WYhURbQ1RjxdwlPswrd+wcnuc
wM/ZsMXLMZcNWKxvBkEZ1oH8kYYnpXB74ePqSRFxBvm3qw4ccQjh3h9QhnusK5XzF4birH/Nf4lX
gA+S6s52M6i9j39YNJiO5IEU3LzEcpFADCfEu5wedkGL6+8CXcrS+lFBnsViiCDQYEmuOQc0VItd
f7vnXWhfl3DogEHYGzBW9V9ipaGbfkGuW0T90qM5ObUQqOGKNdlAyLCejOG2/fxols9xocIkLZp/
7qoA4J+hytg/avsWjrfbfuXtwRd63hpT6ngh6kXmSsQjRrJgHbiQogVAE0ucD97ydOLNGpwGjWv9
sofB4R4yeWAUl1Fg0lhYCoayWxlUFfQKXsq1nuT1ZZg6HlSLcyH0nk+VYpiGHUMxdCsf4hFtwp2J
JoBK3WcbW/kI+k/Vg7UsdcwnUUtFe87y1Ei6QZYRp5fl+GHGuqkYjdVsCbLhlckHORC22kbSkUcv
0uI8iSgcajRUnq1EdXRq9W7o+GADjDv0JayZ8zpWHa2u2I05ye6tNUop4s2++yTpRyiGi/w7i9vz
pPKPi+/ox/2CNVS7rT1qQF0m/GlBVTlmMlSVGIMtuTyFg3yNV57J3M1XtySb0XU4xT9Ti+U+pCfI
kXEVK7jv2Qdo9XJjSisBfra9/tlKnP+rID2wwqeR7NJ6U/vCtT/P3bpLHZC/YLNerviyLYx4fSH7
h8VFPhr+qVUVQNBDAWi1aARoU3E7hq+pYNZmSotgFwjfjJMcGsFqfgkzroZJjtYyoHOVVw7IwcgK
gb9i5ksitbqP5WMjVpD5D804e1TPE4S99/UQBUD/TgHBS0O44IoXCVz2chLHDcgwflEoqQmlalre
cXKQLv9CddZEz/LAzflSe1ZO/EcbMHTNbfqWAvt/4P15hW0xYI/Na0+uVkCfifbCmGmZbywFZR/S
BMIDen+W0v5+jo+MWVhl2LIAauOGtQ3ZYRDat0NJblgPFPLba+TVjYPUnPOwbRlxPWXsn+9wmsPk
9H75fT1+16ir1nlh++5EOXl+QDMaCZXswgp+RQPZZIEyvv26xtI4nDUoXqZti9k5t7VwfIVpD8zV
zU/jRYMgbGVjG9XSrZIe+apFjUfUwo9nM5ltZT/LoupkEQhOovCU7P4McQipB6tXWb1EZP4XOUtj
X1SSQOSaxWuiC1PLsy/GoFNTQn6Zo+wz9fsiC29UpfDkmsX1M7DXtjnJwu7wtVYsRNDaRZl3JfFN
fz6ixAZKEtbAxPtPf83jMRRx0isEepy3JQkaAiUk8+kzEbvvEt5xCNZwDQ67p9DLIAXKDCUsWW5a
5EAzll/JnWkHBYcXD7PLkBqwUiGpEpxaAhao3tXatJqO6rrcI5+nnioSko+vz5lqIuOvQTGFYkEm
UBkN30HSoo1ABHyZWwM4BPFKxRQpxC5zl0Sv0ciBm71TM3G0q3XRxczRl1zKph6ZHMA34szl7yqN
aIWC+qOAbzKBeY4OlnZSAQ2ioVVjvXqlAWg+FYGVzA9GCqjAAc4PU+QGdAEV6uU+iXVxfoKNydPA
yaEVzM9k5OyzMX06FHOD28HqPNRq68zLKsvR/Or8hh17cmTqTLJltFbXmw6jlSxJeM7L3xaByP0p
MFnq4xUEL/sNUIMgqOF8D8x3F7DAFeDvlm2GnUOqo7VoAOa6r5yPU7dzyZV3nRda+mmexmqQAETq
S3KNPc1PhAq3a9kUXiSN5yByrgIAFEly1+whcKQJtVzYXqqQGlAxmeDfpTvUHBb0ylas5p75kpkV
jWQker5a6VTmHcGdVK50o1Gb74L4L4qT3NifM+62rfwzMwfak3yPC6P02DZVV3jNqOpveMDXc1Pk
niBnAwPSJmdMPrxAXuv6IA7K/T+AVO1iPPQzrwO+/oVWhwB4rWohaCIyuTUb76nllIquuEVoK64E
hBNc8pvSLWF/rPfOyuY9xFqfenD6PQP29+swRUqKZKr1lO7uDn8NWinLLYYvfn+Z9xkdirFsxqbg
NOtpJaotCOZOSQqCNBNOQfszo3vLwS0Xyy4fPtNlReeeKblCqAb1O0ENh+8XMHJ1iFSp/dcr+DPS
IXVN1+zYDO2EiVnboT1ICIgSyMafQq3vkMwo+f+ht3Up8cH+8EG6B/MLFK7E9dN0wjLp+XRHxLVA
1GnkmBn53SalHm83sd2M4ewdJhXbaALuZEhKFILrfCNka4I4nrxRAAWZwV995hiDkYzCJYEI3OMc
UQOspYgHJ+cN/yfWYTEH6Vzr6uryCYtHBZ12NlO6D3EVwJEV0FF47/2vUZ4m2ThVnlveWcU3orUn
MZUosAhRwNaIqQ7SrbcJdVXxiNNIThqBUgGh0qu3lwNF0jnFYrOQ8mcmAfO1bgh/2E3mhCDs1D+B
AdHYxMoRIYOLNE3l/enwyB4LniFcCDaujEV59TltoLPjAwIK4JrUmkQzkKGSQGz8oW5KZwjtpW+P
aFZJ2N8l4N/XGWpifgG030t4/xDgHZza+sUH5DcoJzlgL5CrRyMJxKJSl1gatYZBPaOjvSLnvCFt
VR5OJqMl5O4dYnqzKXxUBGGLxGSdEtyAfpLDt8s9O9dU2xYduvsknaOZE2HprWHYNsJH2LsMMnED
63BqXMzsvYD57I9C3IHF4U2TZ4shVE9YlrYW7AzlRcBmmMLgLQEoJnVIfZ7fvNqkfm4iG3E+ayG5
NGlywtAuDwBspWFk3SdxbQoXQg+wUmfY7o2OQVzbUxJH2IypOOKxvREnk6MBYzt9i225JQqQ7yBH
/zKoBvUZnkoKhzlhXkQbTtRxArwjO5/4ka4c4t9VKd8HBjK0KslbNMdLSUbEKsBYVfhFkJvGT4xW
Hx/EM1VgD6LfsyHLQDsNCX89TACfEnBXirRjcwDi8n/sSfE69AHsTI907ZKmoB/xj+QaNMWKFlHl
Q+UlSrYAkHmHXvOK+pD1VpVub4XOVvVqFNi6ImJoEo2/o+SzkZc27WqU1oN57wG4awFJqjoI8HlO
pXB3iFriQg/12m4GIsSF7fvro+7axu5a08WpTMwNppB4BCbEfAaWG+x/fvcovsBcjEQPGjIllq4g
4B7RJZ2OXqtZ8/WD0xJmiPORWfPoEkoz/Z9/1BimpbTHaq6ipluoNoKuTd3wWJC+AKpK4+UuDlZN
yabaNPB99RB8NprllEqoAykuKmQKblxoB1qVKp4YqiPDMa487pWFu97VN17lrUiiiDPAIArJw7WA
j0NcuyGAAHOGyTMQq0zJ7PURlHrzbZguP41fAC8/Sdb4EWU4bWEtxQxPJ7/xZCZlw4dPhNsO8Wsd
DGR4TmTKOLZ3Fil5C2wLuNCHBmLdqD+wOs7Ac1FH0RYfkELX9ZRrsPnDLGq9DYi5W7sUTzq1FfsZ
OwV9LixTWBcrHGRYnV+PNULYmCyFz9hJ6tLqZxjA0l1Cq5FoMEinquEeTBcvMpdAiMQ2JXSDsCjK
ZsfSgsRMwFfW7Ew7t3XsB/yHy6KWckIVoKrj4VEg4Ha6HEBb7ULmvT+ELQkosxAghuBGOQNf1fOk
VZo6qpiCb15SjuPEHAvzf8kQnNTxBYsdtrk1ychflx7mkiUmNPPSbeDCXRhIBaN+EwtDRlBRSWlO
Cb0ApLX03cKtWFLRuifLIyLnFZXdNYEdPlyxS1CGZBiEkaTk8lhgqu3TotspaxmLGqZoUEP9GiRC
dVgUD4jUtIFRYRnSTeK/qqpF15eakDOwUpg90U9J7+OFf6/aC4GceNpOT5YxLg8vv9IOSZEQsr1u
R+wU65XKFZ34J1tl86F+bF2raNhV74EcrKwyAcdtgfBjxllR56dZZK0R3nECzey2WOlB6zdhYwK5
FW3J8+LnGFBYuoTvuLaNms5Tv0vSKlbo5mKgxlcptrD3O1qWKvkOKOYd5cz/CjAilxQx+AZALl0q
lVhB
`pragma protect end_protected
