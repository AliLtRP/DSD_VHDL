// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
XfTbDOFeiTQgL+uuCUgqxyTVzahpbxkP8TOsyOPa16qxP419USBjyPqoq9pC4kMIpPtGN7goBgQo
0Hvt8B0u6J4pecc3SfXM9JO64u9geP8fVGIttgq/6ucUslvlh4jXdSUZr1r38GyxGbmkbR2DYVhb
c6pNZDGG4d6qeYDb2Ld4KEu9k8TB7HqfJUUPr1VxOYfAY3hE0QAQPaeYYjrEUDF6MKBDiuS6x4nH
2iT5FjqnJkoodywda7VmfJKATW2zRV8FKGlSX/Vv502zxhJXxVB2/dbdnDjkZFkvrmqF1XNm3TM/
Msn938Vv+2jbjI6Z9TIzeaxz/Hjp+B87y4BYjA==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
pVlUCtHMuiOHgH1NvDLiEdILG26SnoeulqG48Qeqnu2O0SIbKtP7lJxVw2lEG95TjOiOt+hs7Fpf
+FWXVF4lE3nmaa6SWmjwFSQp8lsJbemYRWbHfCInZYMGUix0IJjxfVrO5Hgk155g4AuAWXvoYv/4
r5YFlRARDSpPsVZdIYzCLRBSpNIhCWDBZepe9D4K+TT5kjZ1t3FsdLa+0t0xy9eDINUCMr+OQYhw
fixEcGPBb3QHKPV+KDcaG+1m9zV+0AAaTO4tLLCr5umEsb/u0zc8bwuNg3xp8P+sACM3DNkA0KZy
7Auh+sWo8DlSR18od2TiqVyU3oEoGy8OiyMPyvwglSIB8jWOsNMMNssNmB8nBFuMHUkikPxWIGeb
pP0aHM1/m8JmyLsW44beAuVEn0xMM/oLTsYDpJ5FqyuHTwhgf4ftl8QuaNzNGsVEMswPr06zvQI4
zE+WXjTwmOHC1374OHAYzf2SMGgSvoE9viT6HDBveZhnGUFX3t1pudvG+b52O0Sn27PGHR/xdXKE
Qp4DGEDCzYlWmC3iNdOG2sTr12e6vprsSIU3jZwkOGXY4lmQWTmmFwdN1hRESSBdOiQa+TRBzg7S
VGFoFD1gq9uX46QKtsMi9VpIZk2t8fXwvSqgVmKDSZBZaZRZZjxCHDn2h9OHuveqAS09WeazurgC
gVszgIlz8EghHjltVsg4x4Oho+evqohEEzAvgi27ygNTzPjuGB5NspZ68JqL0lEBz8I4+xzDoHKU
/gQVmsTBh/q0zGRVZ7IHzwiInrR2Xp1DWsxdFmPPjDmGhkJoTaIyQJfLF9yU4dtI/fm2r4dP7Elp
gLyqG+HDXV+Uzgipa9cifCCJcvkif/vwL2zH/M3UJqfeNrlFzYUgThvyOtzrRE894oUWRX4q8mmA
8J7c016agVrzmTj0gkft38+0VPD+CFBJ4R6ZxaFqP4HZp1yLyQY3hSx/iJnq0s40OPbPOYVN7gRt
wwrpsPy9YeXoBjWma9CmnTAdtTftJhl5VwKxNkKRfBA6y33nDnmRLAWtwlNx9sDf7mzM4Hsc2Hm/
3lF68Uwut5ED5GDf8x4sBOFLGuPoqGW3paKW0R2habqCQb4dSnfcCshnuRO+EorOI0wtpu+WyI2E
QYicjV0fWfvrOjQ2VpMPPCLCS32GoSPqEBgb/RMtNG3n0IOwgkxcnzMSEWJbcFM2Ft/6vPs3aqBD
ZJfV7uSEz/ZMjCUdTwECSbpYeIxJaFuVgdSJbK9HZdeti1HGGDH7f24nWJkxbhGG0yumGirucCxM
Ga/sF6BnC/N2TcIpAJZ0fOCa3UJXUBXmEQ57IWu3fqv0Nhxg57RccnB5VFPsijmG1gR16L/0dhpu
A7hsV9jQZvjzCzQBrmCPMUy6KfKaTFXAHnZcHObrjpIFmaVxItBMko4C6STkNUySG7kKKkE+XTQ7
Npnn0wSqhdzVCzEWqvyjWT3CrV6C87vj1oCGCpxrpaBMdnQwPbOFbQ/JFa4KhFLJntPIgrc7xWVm
Zj15Qz8lbE1XqJ7/oc/VAmGuWQV78gcCnS9MUDlwuYhrhPhBzO1v1HDcjyuWNr7LFl6RuHgQGjba
KO43uuKYjW1nbee06s4SMd7qSLujRMxkU4uQGAdvc3zBueahmw3h+50TJcJtFfsAt/EncgJBx5Co
IzgWQTH14l7GhoJtm8xLi09C03epy8FfCLQ04Bs3jq/WDFq7NeKj/IKy1hOflumTAR+zuzFVLmv9
bxnNIgvkn+WFls7uJS2nFqb27L0bufaflY+NRzf2/QqRJQY0T+mnBIV7U63cu3u4u8kLX4DsZ6Dc
DokP9PMF6IBA6jBeXh+5Gb/0YBRokxK6mgbifWggokEaW0mhPjnkHyxQxrvA0WxMsgv+dZLCV2gX
LVffFb494uCqsg0hVZTekbmZuNKcnn6sb2mY6GfjwpUvcE6hqNViZj6uew1diXDDrAZIXEiStbSm
ghysU2oxftNRlcL6RM0LI+wXMb89L8z4dekYeEQfwADavMsPoIvK2pF2kWIEB5bvoA+6neTZei4z
nnhzX/FTvJ7AX0kVgGqXz9beFhOfjg/39vYJVaSN9SpGN+TthefNOFRTF+489vH6dLpt6kmZPOEm
TPYGeuyj5UANc0xqSsCl9WMYzGu45gwc+AceeEUZv1xI5E7TSwzRXKWVnD+cUsicpwEfGnY0MRFC
ipoiKaeqIaaFIftU7xNZp0Q7oEGIsCnpqu/bePU/88ue3M99KndDAPCYzlRxqA0i7Pyn1Fo56hyc
1iZpRJ7kXUZGUAS7AL7a4XUr3NyiYEWNUp1+G0Sjht0oxvRZ/DOJ0nZFqcvQNcbSoX21g2cu4rcS
aEKygL6ofixLIVaeI9yx3TfFBBTkGlFZsK1lAmPe0k6WGVKL3EbPjQ2GIKyHiFj06ah2Y9uml02O
cpqfOOjxmstHmtJ5d7PTHA8AxV4iraHVa8nxCBTt1/NJ9vDZcP65ewg/OY9g3vJrBkYYPr9tkGL2
bpTOPslOv8iKqH+r42DAq5tVVSNuendLcSPsji3Mm7BoWLmFyfY51XXa5KLpT7BPQaEC7VrvaDY1
BY1TO6qXtH4AUocRPmo0kf1cPMG0DbsC2Vxi/116RaM1xW76mtL9yK3ETbYK1T4161f2Nc9Age8x
tooviWBr2cqQloW8rtnrUWSRxVUcwGWHnXmYbTtOB3IMf6O4r0ZOl+XWKyCqSznPBLEYb5MDSqyI
0ixsUY9JDgnTg2xONISskuiKCGQrQ1YDR8Wl3v+xOCNoPUDvb8Qnx5jFsveBQa3QB8AcVTIesqob
oL2n6mNCd/RCSlpjhCzqLIf03flX8MVmF8KNy7neveK4PeOZ5zPanc54t+SWcVyHKqu/jdyjfdt1
TlstDo22cCyGftKTD+Nyg/8vcz5QoBN+AG2BmPN493S6EnXs8GSth7dyL75H7HV2MDpP0b1hdI61
dTRo8UhTHP/ogqIl/GZ4sx5vrLGHv5ZG//Tu3JzxlYQuvwrnEHOkFCBqJCx7a/NevQoDsQg+ygyh
cJDIU3NG0u3Rp1PzqXZTImtDG/9VPPp3HSMOd86RT5BpUCkDNyRFM8HhZFCsWBpu44Cjm3xx/NLe
sDogpxKZ5mjmUCKmTj/BxcwJ8um3UB2yEHdnHcqGXFRDoP+WpZNBKvTJuCAWx+x5BhGQsrqC+e4N
N5Evk4rEbkW+2c/mt6U7BSQfm5rcGkas1WaFhT6s34BAuSfa7ojDloKzeANc0wJmz12YA8PwIGJY
gRgyfAL/pNxpjNfpVbE37QsBEqusFKdb+O/JR3lktmdp+KHUJLshU6Te4cb5SWYZWUCpH9l7uTEt
llZJFqaN/genRAAIPpmczpJ5g2cJvBSzX9aw7mAG+knfsIjxL5OesoTbugf3eLvU6Ceeeo97XdQi
3x9B9Y48k0l+LmAhQSXdK9Ja5aH/SlRXC2Nua4NMj56dod1pB3OvY/AQEYQUdBuCJNBAgkBWFjrN
6D8Gxpfmfy0Zg2IB+IG5Sw0fOJhxCrsUJcEiliA0nAPRPl7N67QEn/Jwos9X+8EDOEYtJbYauL7B
3iMkDg38wBpqHmmlVUeswIgqtPwpMWvZefpBA0e3O4u27AZ0NI8dw71U3hgDow2yFli8egU5srQP
ZRwpiNJu0Jh3NWUxl5Amrlr17mquWkdhlPawRPD+G2gQ3QKdxelN7ounBdZ1h5zFoGK/kJizD0//
nzmn7D7nORxfLBCRnAYzYFriKd0ir4q15nRk0gE3Zwt7yWAdO+bgeVcQQeuzbjPfdgbjtUpykdoC
xe0po5Yvp6G4bWwSSAgYaIj+6Y3GC+g0LYY1VMnDXO5Di85qJRAY6WV3MZw06Sx7TudJxmsfQkJk
9RcYj8Jq7GvY0jfi7fnzYyphY8zgptuCx9GD/c6WvxnUx/2iu0/sMZSCfVmctDXtfcXPds2lOQt0
IBe63Rfe+LGQ1pOzw2ZH+DbTh1FjBvWFQh5PH5xRNFJTtqfOUn9X2MuGnEAQFv2TK9/Q1Y4P2mf1
bH5Kl/9OibvfYyL9KXY2F/fk6LDH+P95kziQHdbgLcke5HyROeebQPMcmkSngkIx/7tV2jbxIEGS
8LMAkLQF+3LETmy4bZ9oyQboZBXLKS9UUC2ks+5cMsHFtXubyZAaY4H8L2q8CdjqW1081jGM/ix8
kB5IIgRCfH+So8tTCBuDpFbMu3oWh4394bX8F8lVtnNTTLPIqqdPjzKulwNwUHYx1vqxHSFM/Ckm
UmGYpV06xmI71+921ZVM6X/uFJLwSLPS1e7lmY4PKDnsEp+2AGADqFBBlyanokXhBw0C6LiuFbXF
n1RG2ZQOQenbEdu4HNWkteVKlTiHCZrZcqBMaYkTwdVTvxudWtnhPF2867h/F5qreSRLS0xHFHO8
C80XGQgW98dWeZ0uvxooM526Ck0FQsB+dTRJ/rBPUUaamSsyQFyEzUijTAHsWt/KSNMqy9RdygUE
el8QVC/3UsWgffa8A1ZDx42HCgH3iifsI7z8KdVGJ1KVEudBI+yoZBcpyhRsrXFkv0RqDlrHhzG+
W7Er+xD2jowZ66z3TFDQRkJhaNm6EXisIxWbTj+fXoDa8U2J9sY0DbItl8iQaIEERz7wrvRWgCVu
IijyZ1Ln1P9ojF+Cs6f7IktFfZ9s8Th7q9XCQxXaW2qXdv6PSSB0CHe5CJPyIjczkjR4QLzECxjR
SzyN5DmQ7qcE2POk9xz4k7c7e6ZHegyuKWQKpplmQxF4DxpUvEV2rNzPOHtS8f6JD2nLeOn7FU67
v0ALFAaxscx9aG6eGNDoQ/yEbu35jo7wseq9dafWSYxXhKX2PE17dfxt2hFTcMKnm0cydnjeUdPg
QyKyFf37Cwl6BBWZrqBiGJhnk4diAqnAbyZhdAWI+ITYBFvgSg/kRAUqcL1eqqEwibUoiD8eEYrw
AzGOEF6gOJxxTK4SGXfsRlAmAKvEceAZ1D232Kppj87O50z3rsxEBQTPmZpNfa/7L1ayNesAjv9T
ad6U8J+K7JjIP1FaRbjMlDmKUGpUGVIvLxyjMTVWWWDzx77+L1O4pWIf+KbrBPY2vvizjEkGpOVW
z/jNqWpnsq1dUj5ACu4DTJyWBJKgegjesgC/G4eJXCadcSVdnYqS2NK7K+8cRwdcH1siq0aAWWVO
a01BbSdemvg8XvxApzYBsyAiMY4Na/oRsij0CvGEMvSSNeoqIpASsx9MWSrS9Y2Lwo//+RffdHKp
tC8X8iHTlyHoaKqf6+TYjiFnraj2cLbY9ivEUMM5tXGJIRGBcUcxyrzwR92IzKnhj9hqbGavamMh
rbBGrQhXH5hupxtyrBa1SaSOffYw10EcDd8Hkdjn52aFbpe4k+liStxYoew8ZTQLV/HLrAtAiwLb
pggsMyLnI+j5kE46AyTXIzeZPzBFilLJgRJxfbGT+487RyZq9UuGVBXzi6fBPuIRwxaQ2W7PqkTn
NnZuVf2jh+rumfQp+jAfZM++PHkUBqf8yonAL74DNcaSVBBoF4VkREzNLA9YvIchF//wWo7XCod/
YPO13EGhUzM6M4lZaJ9kDKH4nMyWaklbUUdP/Ar1zncDQlLxjAq2NeYqRpEAwEANImFmfMgPx9Lz
qftUOMdB4OzAF8UNIHUMCqULCzi9jp+1oQk5NcbIvU75a+B/+J9jCBqIcCZ1rVCmpy/olN10j92U
aCyxIy6SefU6rr2BGvB6MFNGR/l465owZWEdTze7uMCmY+gh6iX1TPxP+BCc6rgxstXaO4fqIE3j
+SEySNGRvRhVn5Yy5mWRfG4RTrBUVHSXGX+LbBKolBl+ZAluCzjvsS2+yjQ+FcoNfi5siZDf+bEV
bKVdFfiYZSk4IkDbkj2AhZ8ajcgS7nyWqoAAN0Rlt7i9MrvILnLl5GTqA9II3cUvTP7eKyH/a64C
ZvF4Lf/GsWUqnz0W1bzjiPKJ58yItgETuD+qBExerl8j5I1uLBg6PBQQXedws6KWqVbEKGZt33uQ
lDZJ+OnFO5Wm79/lfBYzjYSwnLKcRob0nL1Iet1FQvlpmGmvZp+3OElridaxAHtXaSrmOXVk+VSS
VSmH6eNC8NR55JQuV9V0ozQa2hT2qthrZeBOwHIqo1QXJaAKJUDhhVeLZxaR9vdAQmGhY0CbS/t7
vnXN6skcQESabLfS8kRoGRXsHbkS67v9degwnRTlf2Yej0FxTHusS6MbzRbFsa03HrQOoM9eFtln
/gdRY96o0YBAkbm4rrD9gXPoRy3+S6iv2b4HH2mMBKd5arnqbLNUPbv5VmNrkLluU3pY7PQ5uSNb
jMAvsdIZ+LMso8CWzMkYGCLcJLX+U0/fCUMu+mMhKXv+HJXGvM+2ZlMeE8CXg6oJ/I7/XZjgVbS1
LpG2VPOZUcoGu4uSnu3r24rVOHiaibjS3yeHVoPuCNHwFJopM4Yrwy2LpeWh/uYgC1Ohm+Whxt6J
Lgf1kI7b6WKtNmsWwYivf14ckvQN4xn3SfdnZvblJYsFx58E50xDBoxOwAcvM8Xj4pXeI27GtQar
a3o7j1goR/CUA7kLrlk0DczvQkDFeDfxK5j7Bv9GHH+LZRnau+Rk/pUi7ByOSEoK2Sv00tj8gHCQ
SFA7kB7CQ9O1OXP1ThYA1dzLPsQ/vL3PUwa5xv1vdeF48ht3hxEC9ARqQ+7ftCosgeOGO+iEJEGO
kjhIo2MwFmoXOjhK90oesmGfQNZ8qHGuZoPUnJIJM8iunjIDCFk6aQCLbVWL33plrFER71nkICFx
lkR4jalEJinv8uAjhjvc9RpYGwg/2WytbbVsI48StTTQ3kd4iQysXpG2Z8YkYFdZkAuAE5ug0QGL
QtmGLQ0earf56PLxWi6zZUW0drR17plfsA/D5zIG2akFRyvs0b1TXqJu0g2N/RDbU8ZscrM1lxSL
5hx8K1jJvahB2/zT5sLVlRgOIEZeuZrU7pC5OoD+/L2HOA5ohgBnVzo8ocdUT5UOaBn3XnZJVOr6
uWlohkFnrA/CwCyz3LvMj8ICX5iwMF55E06+fJGfN/+WoP4ZBjVg+rxpfRJa5VK5pOGs/6yBaTFO
ioUdcppSbVYVIK7nXM/XD5Dr81k/VeugFAggq87uvwszA6mYM1j4NboQhWg4ir1Gj+3v1VXPJLUB
/vrPDVOHW0YdHyJZfurDh/EHcus23uW94dmf0EzX8hLp4Ef43q+tPFdCDzEzskThppkDqiWCZPn6
UmnrFAa0gDEksfikag6ZLugVE8XV1FhM3UNWAvPHdeSn9J3hFbJwZBzYk4m8zkkqyXU9HFTUAe4B
AoDKTdjcAN/9LIb77QEvN9r+pI0krwQrAhbfo6H0dqtDsvc17TPEz0sMZZDXF5mEZaP48KfbeJoi
l1CjJFIApNOz5ibbjyrET1QjPnjdhz9EfRCjSsvgErUV687y2h0KCozszeGimRrqAur6fXZzNPjs
zudUspUkTzmvLJVTzxBXyFx738ScKnNpp0CqgFGImbW4gkelVI7jTsNhyUQ8d8GHCA2fWuMx5N5u
6hnpCpFBLOlehFeDeDC23bkhjDDBl2vqzFChvIvvffzzbCQD3uRuhLc3yVo9K1lAX3HI0InzBf+g
5eSop1EaQ/XvDORSqr2w8WSxKek5l1mzUTfYaRDGgbjoKjzZ7RY87rhwI0bs4rfJEd5xpKR3gM1C
x2WJkUTzGymfkzDTjTqngFMyaTaP//c5i5/b+CGRUjOaqfbUwJNVMQCnmMWF0Y/NmVi84fsEU4Pj
47dZuLRpKWdUkR97icOOV/4JvXhJApbfPDhciUVhRH0lP/zRlvhlGYmbdn1hlXgRkH1lSwYL0sqo
frWo2hFtjzDJguCpmeD349AgIU6QmSGWVRT8F79ZgC+VgiGc9lOt1+X4slEydWrCZNXr0V+9naUE
nQvFh0kR2u+/seDNIPCv2P5qFU7YoC/xqBYGvpZ9qU4cSr3ZahbEsDCRU8zxf/uMM0r36FFO9c+J
iccG8a+eacbo682OfDqWpFjNshSShSf1eWx+n3NNeP53nsVLb70uapvYHgDe6JEDUYppGn4gA9c6
Q2RhFUoVtDdYMxC6bhEsSYS7QwSXyQDKee2929XknLk/vjJmPacPDcnzW0JDRzP8FWzdp38Z8WpN
XbjwF0EgVQLdAPwq9ZriBXzy5jSpic45Btqtix6cwG2QcXYYtsrHJ/IV2RngU34dixXac1401fxP
6UhMFJQWvEA75i7O2ZTwIEnqAsC82noXi5VVcRhxW+IPbmEEn1ScjxaW7SNcRPeTV6KCMCqsrZQ8
sKSTb6AlnJZ3gnbh8ZETpPVm2WUVGFwwDRxyfHDqySl4Lc4fbH0HntZNRNi7N425LFINOVXpbaAi
fMLkbqvDFsHJ2Dwex3Bw8ZUgS1qhb8AmRfAF5nTv3D/2CVgbdRqrAUQihft1OTQi/f9o8Z+1PSWa
qXI7mfq2pnUuqYpla1drPl7zlLDhBD3Ear2z+Ox2za0+hVFstSkbFk1UEwFbRUx2vMgEu0JCQ6c0
X7+ImKGRFlw3Fi814gDKHt4xz7iBT+N+7+0DpXqLl91O9GdOtWxuTv0Iz/Iqfo9KxmRxRMtbMj4z
iPZvgIhKKNSfX8ny/yZMGFRZdyTUh6eopZnsnr7h9DAda4bAHUb/4bD045B4rjAmMln6orp8HQvR
/Vf4fpYWLU+QmMtlQluJrue/iw+tF7da7hZdfXxi5kwv2eCfvb8fa7+BsXv7qfFMnBxJei+txrgt
FNs56iseyiVd7oWVtW7cAQTL1yi41/gtBQ4RBvSgwca83IpIhuK43sylmv0J5lZgeLJBXvjX54z1
qg2Z3qsrsl1wYZaTS6FyVT3Y6x6Jd9B0e1oxmzC/klDgZiVULnROCM9QZtYYb/6xyTv//RCiqRRq
uABMcwaaQGCsD4w4TEmjUcYUTGJKJSm5XoeaGB2u6OPvBgSUQwwjFBYAj+ApljnK5p8BdXn5VFB8
WzZWlEumbZnf2exDfzRtvGAJGTrRUbS46LoyYL423KvMUuFnY0mc3yNIhRRpVZ4BK2wgnsSPtnbk
7Rqj0+hRNiLDb8/s0TI93zoTRrf+vrrCnWhOAo3vKodJRqcKmx03DWVNXk/3MJbx6HGZ7FFtt4to
rhXvToke3Iv7+BzJbjoqaTAVWElkqUi+0DFnBHODm58Spym116IGgQOMX9ZIOd5O89sQlqtyU8rb
vahVEw34wi/nxxG/oDsq0wLCr1OBl/ZUfqmj1tDprktegHF+u8Aw9PuuxjctQwhmg+PwZ8ERZ2ad
dgGND8+jvHT4vW6yREF0MS88m5kg5qFhptSX3gNpzikLg2r42g+dYmhPMoXRYONlAyu7L6fiPhku
IZLJpGCjAnkylkJSm3EGQ1a8lniYmgoenaii23Lg3HMeuYAua+0aTJewVtpFn7mmIyuzITfP8M7p
4TIcOQ9Gzl5G0CByQNaAP7l2ixz4ss0ME7aa03wtu7d+tiidP/BBUozeJTLhjxIhKu8TLUOMJK/L
pB1TDhhAHWMYlW2ABLH9+OEuPIRfycKt7/3DIpiZTpqnTebnOnXURgOxHspzICgH8gt4Jt42k9wk
6NV2g0FcYRL6zaDTnDhTVjUtDm3Vh/S78iU04cR8PI8/Od4hoU/oovN8Ru7tlbmtaLC3CbZARlj/
Qn8z7VPvjCa5x5sAjDFIJoF7Ht9GAtQOLHTYs0AM4pFYg/GqpnINQuMQq2/j3WI2Yx0GpvD8k9TC
nyMBiI5JcpWriyy8lKTOP5rdXg7HnjWa7qWS3RTROT9on5TPm/SGOOkudKUbj82evRRxgVBdqCDu
LBU9PCNBVQQlPvpNzftzir6Ccmyhlqh9odufB57p4H8wJrX2x0G5S6XUZ6TSPlvvDge37y6KjHRJ
MCkbwHuUc5Xxzlg7Mfn2XHrRAP52gntCaedhnjvCUO7b0HmoeeFq4jzjKIsV2ugpM6eSJDTkPwuE
EHMxCQZX1YI0NwiikVg5tJixF8lyq/Z2gtpvT6qrGOrXcZrCAMsdcK8d16qbAQCi4XCO643gKVdC
UCF7ooczZjWnJZiRFXbxZJMhGC/ncdATfW8vAMWWiYcOxyIV/LQ4EOnZrGBeuOSY/ANoyqfwUPjR
CKabGgt35pk9zUmd3tIg0ChYTo4kNDhsERYP3Xrk6+D0PRigQ8GvBwU1eayEkT8GirY94BxBbaFT
Tw2VWBbQoJmnjdU+icjtX7zkH3hZ0GiAt/89lUK04HKLxC73GGerzaND2iFw/rZxUD1A7HEvs/sZ
Fqs6I8nSp9eW2FWbXr6YGXIzzB1nzO/tHKuEm8mo1m+oc029iEepOAEyGzKMycOioRGyPdZC49AV
T1D+mL5tdT8h1NThERHffHKzYy3fAApIM3LTTzBcNyWJRyDudPfXmGjzxfaeLd5Nme1lQJkNwQnG
FKmbhoaRdjIuJyDzwTMUQzqgCGj2Obv+xtxw0XS4njtUR2Cj+n2wlbmB47Mju0voQoQVPki97d+/
MatOdnO5QI/nzBPgmgG/GLyyRQi4MbVw1siVWDNSEHa0uxY/3rnQZQxY+de/iWMdJxzwLWwaCHT8
8/yVUd8sIdF9r0aRYuteE3hr9QzDwU1AEhPu20r5DwG0F64mbYby07GncbCXAKUxayT7KO9HSxgf
8wL7j10esFmbpGH0zHksekMXsilr8fAwF58u+Ya6i6VIt4QyhUQngikUoUWv1SJiLHLIHabUVG19
TVXzctiyj9z8Ufkbu3666GAOwfghuqNKRIulN9XD7cMHBwMF14gCyg3FuRpnF3JqzYYL8iOthz2U
iQz+OuY0VPw4Ugq84uSYAXlBmpJLnhV/ll9uK52XoyM6Iy9Kz4L+5CmhvJmfE5+KkKYFqG4w2/BF
uMXqVFaf9NZ4Yo+ZD1Y38ueKO3J8s4MsWV+t/6PGHMzxW5O1KyFNGSIMAYQ/rAqjCPHW9/QHMtCd
SLLO7PXeSbOZfvLmpGA65DgwvgW+IKaVt8d60AHiFD4+U+J6XccoYptN+bNaPtEAFi/WSWv9pxdh
zO6YGe0quLZb96Y4wYXQUXcy2NRUaumPYU2NgRvxrsSHW6fAgKA1AWBYWQDfNvD9NWj0Uy/N6+lN
GgiAmBc/IQVAfn4F5SWNlR/UZdXD75SOGYxf3AnXwde0AOEOQDn8eIW8ciRWC2o/jVByQGkGtm7y
r14U8f8D+dNXn9Wb64Nur92xqCigBlBjGrOdYHbutxx43xXUI49GN8jKbkjlqzCPx+U/tfYJKMnG
7pCSeQoAD9BWthqEFBWyKhEFf+Oxs+z43k4OdCP/yVugr0YvDH3fE0ynN9ZvemNj4UvxnWwOj2/p
qkDhaxl9p6k+e2Tzjj72kLuEOsIwAvWX+V3qi+fy493SSURuGYJ3R30VlB+MZnTncsE+X8fTXCzk
CH9iL2oMTIQq+e38xrmNYX3M+whdO5UuyephZUpZcVMzd1jnO16RYGEPQcU57JMEMGBt+HIVsuCo
CSml/dW3IpPdPwsoVq2q1tGcyBSeNpgKBr8Ayez3aF3OUKkmJPalg2/e5ezUlG3tIVybtTFcRrWE
XxaNtXTYhnr+EIL4e4g6miSeC3Epek9rmOGOmCj3d1RopQPPZ2MJkmQMAL5IvysWUGvUgoNB1MFL
5b7DZzlvOlj2Ga4Wwk4to4QEgQKF+U06mxf1Jr+3dPdUVLNTJXJzqw4PrvctftOEIxCMbpxmLQ4g
a+jGa8q4xXbK2o/sZM2iAOwXBc60osVWzXfW9U8y/McATH379ezRd23dnsJi5x5qJdIywOqzo5ux
Cd6We2uaUMrbcDgL7eYzO7RzeUkO+7ay5XQpH8oh3qkeEQn7GDLiXf1hyolLdGliTi3DGRBU9y5o
tJENcV9jo95/IHlo5EWV07Wol3ZmGnCQiJXaY8bdifLFFL9127eZRH0USHhGLA5DJ5NDAJt/v9OD
xq/ftPeSeBYwOih+DcypwgX7B44c+JTtdniMgmFQXvlB+UVkRFPdTV34ZfYoyxG6yno4RghjLUf2
N+gLtcj+wuiPJHMYc733jAap2Gh6boesorfc51/6P0TQk0C64p54adqQm0CV7/93Ra3aMaSR0cw6
AVLTd7Kh1XEmKMmustysVqL8xTm8Q6nk8Nw1zJNkSEghonBM8iNXaOnEFK3YigpPNkZMjJqj69nO
gdfEW3jIAMMRVFaKyvt8L7Tn6rPERmCnkIan7oHAxEx7ETwwzwin9l+jdOsQqsZmKwHTn+LoALB/
AHsPHGjcrMe2Vw6uLLtRTkVywioauyrbzL0HVxAwz60TeXynTeQRoEFYckAcUWEWkE1waT7G+/9f
thMjPtAo04EXuRtK046Z3Ab/UOPpmpB10HiVy9Y13oB+Wi9zdUGJ2LbV/CMhiR2ehP6Smtiby/hS
ByqtSy1vOAVuPJ8ea4h0dTW42mgAH+RgcnFh7wQUQcNef8Yor5gSm2ljjSFgIeOaCM9HEh8PebYC
u93wnsZvp7cMaZTZprYLFSQ7mNVlWzEQaf3lzGrKnSuTHx2Sl6RYw6FtVwV+O5yx5fB4MVU74uIe
Bdc+E13xAkoU5LaR4DDU4zxia9ln4o1GA4FC53jnwDA5L4/gBZ5Q9bPiShOO1YffbD+1ZicyPrbT
5PvEPr36gSBXFuy33WmjEKjUajXHkvr3ioBthvrMcBSnVRMRvvlcoEJVgB9gaeG66xZ74CtoUFsg
+RnHET/yJ7TkYHPJ56YrygJbkXGuM5+KU1n4UBxJuDiH+WxCqyX3I22X4sqUzevQrZ/1J7m9TPWB
HF5bfjqsttmGfCAfIgGjhmiymMcED2e2izkH0d6blxApfW8LFggXrLmT9DAoMHmGsQzoaJAUYsXI
AsT+shiy2WH69cwntcGeN6TTHAsimXGSA4vrYN/e6OIbkGr+hk5NsVtK05WmNzxZft6y+GhNzg/Q
Rlf7Izk6LsKEyufaWTf6lWezZSRR7Dqhd/bj73JRJl/q6q8jIy8wktGMargDjEz9b8JKLmKRwhGX
W9HwlIziCgK0VNc2QkW4KSzJASEJDoY3l4el0R1+I7HqjNeZUWDfhSyz6H/tktJAbKWdt+lOiwBQ
gHHirwtp+IWYBOw4OGiJmgWxzDyjDzm0MGaFe84Ah+Ay/MPsZhiiNPjtJfg8NsBs8/KXa9C9OEQa
oh183KQbBSlIikfUHZjsC4gp2pW6rEenBxVjkmvpgY/cP/FJDLIpz9ssQPLj+NTIz2nx8Pr40YdA
Eldtq3EZZ29pW+U08e3OhndvGHqdDIakbqhVW2zTrwSEbinELQGDli3FKSwxaOFoNn2/SUzGe3/O
3svYiiLKJSMTNnmX8SnOGG40ZqjcrEXBKAaE+GJ2XfMjvdgtn6DM5PMrX/t2HejOtvlRZKoB1Pbm
pEkgB9Oz8/ctU9Jbf/aa9+fE8gifig1gxHdqSof/qs/DieBgtOkluOQB5MZLZ5/NIcvSxEqdTIJg
axIx77oHv3QDu04zeUTGNancZGTtC21zJIJEBBr9cAhkz7vGeGAOoGIBVYAfnNwgNVs3LRC8EMNn
xhqtgKdNNwdmFpq40xzxbpqTNMYG9JP65TyZrwVLMYtXYj/36dJNRWX+w+bom/VWsbNeb+aGEcs0
fMCjOcd60NyD5SWgMAmHXJc1md5KOEpiyvbPEu0GQTdSNcukcSbWx9dej14d1H4jwJ5pTCzHXRor
B8w24pjtoScboV9JSJelpceK/7jMNZFEGxxc64gWlFpG4SF8ksw7THXPbhUPDl3+kPsrTtYHWnOI
EGcvtKyHZfM/Vfjk4oyl65QmkjoKVir81f38NymSSX3FFtg4SNg2xP1pWc5zzE56q2Z87lafyOMf
CWfQgCNRUxztYQgJRurgJ+bcRZ08NugjNRp9OdI3xd9fpTzpkAQrgzrOma8ktjWj37w/6w+wQgwb
1JTwdIsIbo2ZZyJK+6TkzdIcPv32DNe0espfspVQD7SbqtH6+BIsIgse3sIOGogPj6PPkq6GmArM
vBnSAdB3nds8lsqYdqhWk4KnPpVY4H9iPWDOhRMD9WPoIpXCseEg23mS8IRWCMBdrt+XNFWwOpDP
crmtqilQUpVmAhn2vssJioE5g4S8mP3c/jcIG/HVrSA/6GqQpMJbFQuMD7BbRxdXEAZsIMrOyr+W
vGCeOfN+2pz0QU7lMJ0KMO3SHrY8c/QalmgVBp+MY3dq/kXxtNR8DJ5je8hMl58PeREINL3VD1w2
oHFPm4KgE5NfuNZHq7X0tOHrI5CmV1AT7qXByPV7upnTf4bsvKHrmHCN9P9iZVgdiud9dkTOrY2G
6oeuVuJzg0MEcsc7TjDJ6S4ZsZ+tJj87+ok+XwLRotItaaRpZoAVRfIWGyq9cQFW/Nod4C/iCmTH
K3lMQRUJUqWaxISsTtSCBfDKqyj4dJJ//BwbMeHcYw0cbiU9XNKwfKpUtPfiY0g4eG3mEa1XLjeW
UfzsAy9qu4NwIpSM+81qJgoxkLfEWFtBjL6MSzGM6ktGuO+kja33hLf6YbvIbD6DQNtdb2SSzfdo
MSsyziJGjdgPdwEumLHMxnBrgtDYk37ouyTv+neDSj1jKtnl/cw2n6Y9VAOX7R1njRXzdrMOj5zP
tk1yXoTdtOQQuvxISzsRk2Lcdoiy52j2TPwAsMS2aBoniTZ3KCwZ5uvKeQzy10zga4pnW4XzstLE
jDfB0U3zRcRSDP8/qLXBDVGdLauode6zZ9a2tlumvts9Ikb9ncUL8BhnBuwltM6fptPurXC0y5nG
6fFwhkdsCIq8ZHKSBXtrJqQPtuJOo5eyiWghEcZnWi2rnuOk85njXlmIB8Mc2nrywSZUdmWxQrKm
8PjUrK0ggoLZs0aNrTHBRLAYo/XTOsYxP/U3MfkhmeDrhCzOSG9Ef6RYse30sCZiSJtdwasNWoCW
3v0NMxX7YjhzicEtrM+US76wJFiXCG38RoelxkeeTqImhf4+Bl9BGQ3IstIU4XHEQs6Fp/1Iw2Yu
O6F+C7AfLgY8MFJSNNQd2hy/j88RRilgrE1TgGCSz8iU78FqfASJfitHRJ3FtHuM+lC6TVjqmAjq
l34Gyb5IdmMoWcoa44Y9XMylWpNyUVUXuNyxtXI+JgIC69H+/OhoqhITY228Do+M6dEeE/tr+rSs
4pVaKybn/LGhV14oZSdwXC9s2sXE2Tkn9ZRJ0wsH67LE1rdoiV2Vbwr93lqgjieXs0UQDPGzhugE
XSoTwxWJjLRSu6gTVVvx/bbMQtCI8BoeVX0U0NCj6qySZxrZ0PC4NtswILR7/8MBqZzJaf1lywH9
Fv3hhVxJsIlicN/oSPK6bV2XL+ZHf6SNVU5tzG2fBYQOQWb+RYFc77yHEcAyzcnXx7444mkpidHb
XxkU2FFAUSJXQH5TNALVZZuiGiwzJeYb/CuV5LuC+2EMsRY1+9u8TONRoGRgo9zqR+oibzX/ZA6V
xmudJBmvJZtIggVPUW/9A27WVje90st3Mz/P3u8cS+iQ6t7JGPX34dY8h/WHg+GjV/hT5WruKJwS
LxhvIz5CqM355q5RlbYy4FvK9cAIry1BdEesa7zMeb3Pjd8il3Z55ZVGVpfSxxrgMGPd+8Z80gSb
o/16RtsJao71jtATf3lFo5Oy3/wvXJnIcTp0s0TQhxXHq7k110OE9IW2E0DuPGVCk76H51h+dJX2
c5jTgm27wPfsZOuG7yqfLA8MNnBRlFOtSizfT9yNOvQ1gqFMuiPrY8qffogh2wKnSxraVJsrn2+7
g0QH7eAi+3hB03DbBwxPsNpTMwgAMDIHUHANKeGoIbvB5SprbBABripPhsfJgD8YM6kDRQ5vIU9P
gBxc1dKX/LByXEaBTAMqZS3wIiOgUKPZwffH4SxNRtzW7ZOTtZcgbELd80lbzAyXfl41MVPLsZYF
jfW+KQHMvHfxDq9yX71hqgh6G14oiY9QWFFgkjZfHI/YmznqgLFL17Ezctko07V+557XaegM01Nq
CysmOqiYIR35JA1UZL0Ss/IV7onM2xfuyqohqduHU+eN0ffvCuG71vNH13EGw+UT1YpXDbiP58K+
3OwUhN7KGKNakdkxjA1FDvmJDAAbuIysWrfgscezLwBfTJwmygiTOgOTGl2Hh86tYJGQ71EB225E
DD9opE8vYUzsDvGZ3jKDEHg7h8NxcVONh1LkJ+vsb3fUkww7312v6x5USSx96ardeTn/pdtq3MZc
gzRviHIvYJpBI4hu9K4K2KRQkVNtvJBIg71Q9warWoni5vNWVXp/pKabhgacoEctT10g4XbwPSDV
FjjRSSsN+nyy3n4AyZeFs+kUe90ufqxs/4XD55EytPkImAD7nLwHQXRfaQOl+6SyXux8NLnSZfxP
Tz0VJvDQq7uirq7FsuSE4a89n/s57sbD1ntPj9y892aFPYQvPQrl1jpxNlFqTHz3ZUccNVtvTH9Q
RxYPXgrBRYKi64cl3aWNRS8YaXEnWXM8eyzMeqzP04+/fPPrnr+wSf3NDVPhwUX4BXOfZJ4MwUjn
Hdhc9mRnsQ3G/VrbMDNflEqjN+IM5ax6Uuaf2QAkzZCoRg955/3nBfGvKmM67sXtYHbJKJI2V1/Y
SV/BG4rwfsoXf68sMvVYycSdqWFRpnfyclatsMrJmR1zxMFyzj2iYM744JP535JYuTpnKkRcEAw/
RIRMCFK7K2f/Xf2MtFNtTypacq3xoR+lWUujB/ArbjUiUmkBjj/z0JZfagoJhghA9bEHagjrZkBy
pnJec98n1o6lwbv1mSbFRedwm0kc4xmh9wIRcaAVwPslw4frQndaa9sIbJmrawCq1K+6z+FdbHxg
CfGzxmGWYsPatIxrxgMrMHgbw63KUhuuSJV4SnJIXdOZazNYTzkrDnU7N4lTPSrn9VeyrMkXhW7E
blaLpJg2RoCZl5GAy5q+kIvvy7VASCbvM4bMK7gl6VRTo1mBXAu32wE3RvLpDyU++/ik8xhxi44f
1p03ONOVzLXnROHnFFvDzBda/YzjncyMFHIB0BQv+BREcABI8z0itSXZuS/OKo0jqS2PqzTgycjq
osAVLHuZQJnKpNeHDW87QClOJ6LBDLLcu4zJC6rTzrOnz2KzhnhX9j3hdkYD3CnpDXO/Dvl/3v7R
m2oT40CrVBxUIo8tDEP63W2koJMpEeJuS3pNDSCSY/xHG4PzVkIXWkAYsyVLrGqi08NASTMy5ewU
+iHF1jOu4Te1lyxMF+x6Wc9Pti7y+JG9rNr+mYh4Ob8ITEubW6lCpRnQbC9heOzRPj6/yUt6FCvX
tbuhrOSZkoYCIfbBFFnEzM3ygeNTj60+pUJupsAhsouG4FOVLXh+zaUrzNAk8jHqX7F3w2x9I64J
FXe6tdo93rFBQKtl5WO/HgbAozRJYCqorC3b4Czl2uB9TWJapTknZGaJJgUcvSTnfeMlSOZqrdHJ
RBPpQ7vAn227XeBASvfY/8Hmn/ma2wkdKW9gbAIM2EB+wlrWWHWyjOlLCZfPFyLIvQYlsropIxHd
+iY1X91rvqbpN9TKSuAINTn7cQoVajzXtxEwj6tZwRDIvudDnsZdxTXQkz25z1Dnz6Q9/wEpkW+B
ej332zxBNVVSOdpx519FNywhadZGcTLFnOyKfe2mXVV4twCky/RNYVhU77PGNhGGXeqCVoc93HKT
DJFdLZgFT8sgP0cMi57Kq54X7An/TWa1SVlxqUAeDO81cIVBLnMVb+VIdRxWSXUcQ0Un20IR5rn6
VydRSXQGCRvlvXS4msewmCz/EjnPnRz0m3+AnripdkSVBBLnfe66cPz4ZMDQw5CDiH9Ey/ZJk+B/
LkHgm1xhjbWZPzENphlZSJ5DCSCPQPJSyo1HzKXYaR0lp6XO07bGPYNNQq/cl2ITZtlK86hmVvW+
vmOULP+h9Fob4J5kfZ5OV6xbSauj0vh/GLmuqQMSvqSa+tqZOxFo0X15ejQxQx1OU4G21H70LNfA
9+6AZwJNLEh5H5SCzmjfHwmlnQLvoZ1tvfgYF/2j84QCbjLwbGw2GsVP10NM67tNuo3p7UcZpvI8
dRuOr06XuzE2FMj2WrCZwTzV6RLpkbmBs4Jtjv1VyUpcLXACx/P0wLnl9lhiR029YLer6aPx12VE
G9Q326zDA0EsSA0GWeKzx703XW2UkD5gHjQB0fa8yuHJ1RY7SDrOV3Oeyu7gcNc8mcAmUpnVqtue
viZzrndmcmVulAcv9SbBf5mkOcsec5heTq4lOqqKkgHrgafG0fYANxL+dYkGv52uWECwB+GFzjGP
EYoZdRX7vg+USvu457ZRPBZ2Mrr3VnOl/Fb76n6+ct1lQLgZqhtRR96CSJXMWoR1t/oX06RHJ/Gg
XdZ+dDr8m20PZakzab9jUE7EIqkIvmSztRhqr8ANo9yWUeR2g1iX6Z3tFbBJROlHuHrEavlptICM
ft9+xWG2DI9Cq6cGStrBfXeDgdt3utHCizPQxwOD0mwWhnsQoF6rGZNo+IfjPcd42xWlYN02/qI9
01VIP7VtkpqNPuKq8/smFegwJgBB1IdPKrWRiSbslKM/eLNSiv83IHMr+c9pQi6rnWpvq1s5AC+q
Hyaifk3PB4kQ8O13eVpVL4csn6DPsQq1wvU+nC2v6ktUbp0apL+i4y44T/u8/zDRcTnnRjPqQxoD
ZzLs4PAckpUaezml//TTzItdio5cGkSC0DiCL++/c5CqFhZwA494DSLoG5IHCDDWJcpTtzGTJkFT
JlmbzGEPlHvIhyk4pVRkWJqnbDD+vtzvbazfzbc5G5u+vJbbk+PGBkjPBKgPaYnPubOEsao0o9YS
OWG0uSFVfjy9Qab+1EUjqfMaPNu7/c+tQF9oJO1m+phh4KjoPM8v/i4qLdx+nGy2dSNwnPTsyyff
uA7aB7mqGtHF7MDjXp+evUI46Khv8KUSYZ85ry14Lu/j8R73KiyXoy8brBaH5CXAeZ+iQOebTAYK
pi8u92z8g1dnSsNhBMtls8A0zCnCKlDz2If9kW8kz6KdMn4K23UaF7U2aeOsAiv+BWFDMIcUYmv7
MVG0LLc+wyRXhI9lo7bSKSYpbhKpznxRUon2Qplczira1EpocXhj5FOiOMQLwxI8V1/oIFJwRvcJ
QZQsQFqdg6TLocsFkCDxpttQS4m7FdYql18hZTfhnYlqXXInfGQoee13rhNqdH1CeVBXe4mPT3tD
PneOymeC/yS6cXbTDe/fQ08AmaCIdukD1+1cuNtS4pRGmcf9K4kZi/sfsTz+BD2dMbhZHjcU9C2a
ujINnYsVOQicEhkaKst6FiFPMwO/omwZ4M6xe7tpWV0VZudSEYkcpTvYQ4zMzm+z+2dEubz9q7Su
tODwSnPx50hAw0ns3YbElEt34Mg6Sb2MB8wBuEuzhv19azBkljhXdHLWpcSxXrEn7848hHz6V44M
S3i1FkDnEgzKP/GS8gCxiE8sHSudP2KZsXC4qWTlzSeoUfXg83esyAm7UVonZ9VHLZRZTnkF9OYH
8ZKoxku9OpwWqyCq2LZbRtYHHmhXaqKq7TkwqdLxxHS+qpv5TPQ8wn19sKGBnjhuGA7elZ0S21D0
92gfrH1RXpnmE9zfzJgxF9lp63JP45HpTI3S3Wy0DQ1pbE1soLiKluInF/KjVlG+x5PnDwudqPCS
9T0rSSfOccZB3D0pXSWlhNfwx5v1tlENYmJR13yca7LGolcJAZMnviyhNB1EyjSzDsgSJjjbjWX2
0a9AnqQxDfIAjkqpG2ritk0tljd0l+rwhSAam5FCtXeGoTO7D5mfo3uvSCU1ZG2o+FeRmM3P8b3U
v3JLim+xoTQ3tes1z8DwHgKryTLT9aFWL8GgKsa7BEYuaiHf9dmZXd4hCrf5I3d7O+a7oQ1jfsP8
9ai9zmOjymAMIIbsfa1HqvIuZnSQqaFOx2vxOguXefBXN9PZdbqpDKAs84ms46qjqS+Pad3F0tc5
iNRJFXE/CE6m2r7JMQjnyMEk34uKIpMf6PpMgh7CUav/FPx6Kpb9k2WoYUBDQnhuAEKN4/AUHIzZ
TQsl6iBFZ+PUq0NNPHMfacrMzmZFxbGLozxAvEtklYCXC8Xy9qcy2V/AyMxiseRAReYKZAvXZVSJ
RmIIKf7Ld4vxGam9FSlRYfUGWZDPFqoP7hHMOoVXoG5er0n19mFVq5dfy3zfzZIzxEWs9lQG5s4s
06Nry0SQNCghiJIYHIyhEHgW4MjSbVzfsfLsT0b+uobvUfNeE32ZEyOpSTDC3GRLVafO+u+2+nTL
yccEnQYFq15sYKUOptUumEPXptzq5jPu1WhameQq1wa7rVimFGWn+nVIGv7ZPT4RrQWDWgvfTXkI
yps8cTBIm9UQHJjUzJ1iGVoxJTUhb8s+gm+Dctd6Il9kng/H8bHozm5G1QWtgcsKyCcj471gdZ8x
h/tcGu0BNh492voNug1kq3A6HxkvGxXy8Pe8JojkioztuQsQB8Y68RhtEDGIUHUtYEPpK2XQWwyv
DfZIeAzXU95iA5+HwxFs8d1g0Hc9cnrZc4NCsucYGl7GXMF9T3EVqQ8wS6vRETpmczGPdUj9rnna
En9S5RWWiRqykMwpb5sujCT6HfekTWIrlWgK715o9oEx5wT11wLzvSOTA9qpB3HEqNvkPstiEHUX
l0M33W/H6dCjB22OocKe+8Ntkl0oMsViS/i5FvoXVwzje/g/WoXd4wxPSFCLa8H7txpkIiGHihtS
OM0VzxyCm3B70I2B/lae8ty1R6PX4WR44X+/Nx6pyB2YKGpjzx0WuFnFR9JMPY1fSTgyBAhBxVVc
qUrMPMTuAkX8kkRtkcOLVUibYnPP3x7vHtIdmawwH/kVbPD2gmbFSI7T44ao5CMoavNlGCaIhRs7
e50Py0+7u2wfhTJrReGn6J9dyglIti82cwQTpGtszYalwvnj8IWy2YL9SabN6dmsusBKvI4lCFcn
fTN17zYWJNbanTspZpue1FAZX71n8TuN/0/iTEHX5QR775Lg7+vnROMo0aTmf5wumNfRIfZNW7cf
rZnmF9/IwwiXzIP3igK2ZldUv46bJZqHX0HYzvrUFaUoZ4f6CY1Z+hlLrs+JR35tKMycMIOEqgDJ
t9v/3uBVG6Aaz+LX74ilQzVXGDaYOv7h/48WAmjLl7aRPagu8vDWCHrnYS1X8uJHXnwXXE5Ta0+l
ocxnDmjmXxpQKZO4YCNQzkFiIehFT5C1NZYZ0ozeU376p0jShsYmB6YLJUbDwYp5txTtcWvPMg/+
QB1Dr+WNNlq/E6OaOpkHyvZYnC64xRRFyznP4Ew6sNGv8Sz62/z8MYA97kzQU4MgJApZIRdP9Dnf
OgMUYHHfiz60i1eXxyV7i5LDOGKTUU7GlLKwYLdwgkDBdIFFdbG4ysiyf5aaGxXXHyp/KFHvIKbg
6dNCHMLIffYlfsKI9OGNcQsuZSxmUnjqdU+NDF1iMvywtHvPCGoM0JaN/gaf28Oo/8e7CmjxsBai
SRr4UsdzA5VitAKMJL6KcJGL+I50rvR6A9dHuMCKF2fwln88D9b+6h3g3AyEQOttYdb8ERq/s4fF
R8xeXFWR8K77bnzhMOl+BDpvYkQQGNUFsPcvrmfheNgFhL96ZDAie4V6uaAg2vejH1bos/sPQbcR
nSLgyWwU7Wi09AUY+un2Nu3A8EuxDtW4PezY7Df4JtBNEL3smcKlr/1N0jDmgIG0BcG4dcB5hQG0
nGGWYXwEcUYc/kjWHWhky1JJ8XqyaWltKAFUVJINi1EqTNJALQSUREPgwtNXXE/SlhWath1Ku6uI
rFYCqeK34vcXNBgnTQ3kc/YqC58egoKJqkln8WLvBt3VyUmuGwrwNrZSmTKVYa7JRW8GYi8hugHZ
6J+Vh9E4GLhKS9f2+7z6mZxPclRiKFWqyEGWvBmTF1cE9hcbjWr+vhAJdNvRUUtmDtOfjhMhvi+p
v3w8tt/7QfxIckX5QyIQiQ9OTRD1C9Te3qflW15EhHy2RSuN3c1Zmpgp+glWM0r0fTtLBlxnUE1H
TdlDyW4wlGOd69rpAj1/C43KVOZfpUN6L6IsajP6H56ohDPQW8KyhcIHmVt/QWC7iG5Mq4Mug8T4
llpt92IKxoKVP+1Ixdjx4KRuYM80Vz6hXTyRK5m9yo9Oj+GG+9V5/MMSC9EA2tOLUzD0HTEpditY
TPkW84Ja+/vyU3Q2j8z5mUvevrfMQOfq2h5Wlz/iYj+YO7FPFGM+u7QmzF7tlir7163eKy6urI6F
0VmAA5/m5vM6NHe+uL6wEYwuGptniaHsfp9Sw8/BVRtDGxfhSTu7WbnhMfLfSReNV2DH1Q6o7h9W
RlthEdXAb7IbzUjykw1Z+cBoZG3emQnkvMe8GQE8LGh5kHZbDdZvz0OHDY4xk8xFLaFY+Aen/zo2
fvh5cU2jX97m5s4iAAJgPEwVjDuZ+RGSi003AwxsfiMYnQEuwPJk38SUdtuRh7ki0Fx/lO7zSvyX
7IKucjTDFBZUcRgOG7hrmKy59h30y7A/jxd4lW5Hwspm4a086ttxmLHIGEn3wUfFAsl6FjJq3iaB
mkuIFnOjH2RneACtYiMUDGF5tRORFBQXscAj1yNQtITD3+FiJG9tru6hQu7uH/mar6eEULhRGUKs
T3n/FZOj/RAcOvyQuJtWxOxZuDP3Mokfdx4fidXjhidHp7F7CqY4KSeR/Md69OlxMuJtyf75B8Wa
DwnohX67aKMnxoxHP7LHNvnuHAUlr5xHqJLs/KsZ3+AHezls4T04RrLVj7tCR8AS7ulHevzBWRBD
pvBR//490Ng6zwolmcQxm603qHWf5hrXHG639Bc+hiqbdNLSfBhXVHwQ0hsMGbvtdV4EAp0eQLVO
9BbzIhy+mXtpEU+DNW0MLc8a0DDk/fMjkTa/Se912HQEs/M3tZIBcbBjoWrPTaJuVZ4P259k3bZL
9XobfMVo5/b1UVy2v8x1kZiBiKxtmtTzH34auI/DqpByirSIAnHVPQvnfBbJ8z9ot3bD7xfburEr
DzkUO8tZ6jraFs7bo1MkWleLwqKivhVBXblwp+YEc2gJ8ylbpvAFNnnSjjBUCyipRuG87wP7KR7y
LgKCwShd7DWS1VZRZCXp5KDaBjylTLKCr6su6+1zsBFlyux5qCBrqQwt7LxANb9nRY0/5ZdLw9IV
xPa74Ef/fEG1pSjRDAPZvos4LVq/1kTcN96Ugyri0++z98GoXqCXpZkhrx7gM52KVVSWhK1uH6Gv
OaSgIOSSxODEivq0a87644G1kzTbuYp3Han80DqoGGrLgMsO1opgN+qjYBDNN8/dPxXZtlnYjQSb
qqEnH7jsrruzXH5REAHwKpNOhCSIKluqbAQN+KyvxJQ+eHtNNaKXd9YdFJj8VH+ZplCzyBr3dZVA
lK9AyIShbO4ynvmRmsdFqLVg3H/3k4ytK7e9kspEuO1NIbB0ENCmeVT17OOForpkD4UaVkn4J5jl
WZDVTR2AfxE+msiGB5ZGpkmj1oa1aCw4pz8FNdnnETNfLKvzu2HtiaKRxocpbFlAII+d7d7IvT1f
rnQBRrFzC72SA0ooQukZs/VKNnuWFV2dIMMAI1dTHaB+Mau807/GMA+ZSVeXmsXIL7tq/ianz2ep
qkMGp5OBb4O6yE+Yfyd4wbzLkqH0BYUT8UhT7X1ZlMEjawu2x8w6brHGwgYVzA1630+svDS4gWUt
NygujYqe1VcfdrNOsHM8oCyQP8RwpejZYMNOmn/R83duX6RP5GTcIC5siOK7WIKALNP0rNT1I7eM
jrbWS2AmKBwp0hl/pKiYbvmvUsTH0HKMSsNLd5Bet+D+OOGNZ4zz0CSr6fFZ+MuacD8ViXusC6JT
EYa/A8qds9eVwDoa4SjumDMU54ovnfmLahKl5OerX9yWfL8oAXIfkhIWzy1lsqJ3Xi/RXxRAwL+3
BSPr5CGJDjU4tDmUjAAhCR7ryiTkq9LkhYarcVREjXTzC/+MDc3o/9M2GCUFL+ReuqzTwH3MrGBJ
YZkHQX6cxXTL6+lMqUL6ux5S3ECHIi1VH7BBzlICdAjRZocNbHKub+lN2g0EOyZwW+7Bb8K1wWxy
UNMtE5g47KEsD/3yh4u60DhCyNZ+NF8f6BCOGUrIT4C+bYApQhvKo+UwNsyhFT3EAP9H9rC5kceF
CPk5tV4m8Am5MJIc/Gx8yDZ9TKQSpwdjK2Y/FSTtyn5n3G+WJePQMtDdue31anpIuub1HUH9GedG
SCeUodL0QLdBSKzKhjo+bpaX9WD3pH6CIEoaasoNaEp/jWWbgcAJfUJhTNBi3qAnjcoJ1Uy71C8h
q9kCKOVED8ljRmAFuJIZbHO39Bea98e5LTMBknIKuR9/dvPesZREw/OkZVEbzAl4/ZvixDo73FUD
luYH6/pGMvG1c0zJqaC3+wTMhnTsesdlHcH+z9GP86JNhneKw+ZhN8fwAg497w6wmkPkxiWGCAlD
Q7x0Q+My7BAr0uNT4jfZcooG0WMI3dg4vJtFvgqdJz5GyRgFwT92fp4GbBYSBJ3dcxK3WOP8kGbD
Mn3BvLKF2Wj2xuC2selt9kxT1SViax10VBpAd9XqLA+GEjpE31VNsIaJH2oP7g9YyJW59rA1fL/z
F0YI3lawq1/3U+BUTlOE+336kKuCuBgRk+c6xy/xegpZ/BC1tM6pU15uBvP8Tx9lMtSfv6V98K93
ZUDjsxxzUrZjjmotcSNAQ/ykEtsJIkasHEtRIWMTdbnXKKxCKvsPMU3GDv4+FJ7CJxvJKhmtX25V
iE4I/1QAMBm2114Dn/gC/rHMqeI3O793yoGetlds3XQ+qyzFULckMJlJNizuXNcBlF+ZrxMZ4U5U
ySBwMFdXKI+yWKDBW6luf6O3dtElCIHFwG9QFsC9LpYKf0omn/6S6HewL/zjhoMBr4LxU2hIDeXu
o9Kww96Y5joLrbNZIxyiuqGutSp3tWy6bNq7Tzlfjftuz9kT7E8Y5P88m2F4XwAcRRr6Nlc/to5j
/mmdcnz8MeERbKqoyMjJU25ICPhRFAd4Xhu8muRW9tFSxDqMRCIU8M0x+0E+pMQf18/TdV0RyHQs
jOewau6Khu3c4b9+vQGY+PfJIyMWiLLKKWl/Hlt4Ujhi+xk9nzJg/aPPGmarZDF16jDYr0nSNSHf
4m1h3bplp0QfK73hshh7TwOIvazdXlelty69UPGsVCZEiUiSPz6U7WtHf+MmUxlucgsPS5knOJ4q
1qqnIhir1Sljt1YvGDfsDvn/NuSQof2+otmlI3kzXgWRzkKO70qePT5cFSu/5pq19M2dMBgGAiSR
Jbx1WUCnbpgOJEpAn9csDOLkABT30qA2C05X6DfLzefv3OU/1QayLV6Yji3FOqdvXH1BPDV+GB79
P+JPd4eJ+kYqM17r70MSJO+M8bgSKvmJbacMYTKOraXTHGmz975AFxbSRInu9aBvK6ZC5dckG6g7
1XKS6shMyaDFuGFaPF63WOsX89/boyaCPaGXBC24u0UwXV+pHEKM8v7doGdKy4JaF10vvb1Go4dJ
IW3jJGyPcRLGNk2MzSDf5ZdFS3FS1LcnTHZfFgyGqnLeevfzWyykqqkNV2Jv7c/o5ApB4wuMZn53
s9wxfEPm5t+Ghnbi+MVp3/yWFzlMij/rHa2AEserSsaEPZ2t8BsEOBV1JrNo30V2qm4BMXR+rMt9
pvsFrqccn5lMq/2v/mk1PzRFERoTxT3hSi+S6J/jGRHA2S1B2Vl6dMaWeu9FzAaSS3WMAkNJi0cI
LLnxDO8cu1z0ZbrXmLmUMCzM2LVW6PigXgl6Ea7p6Il8stc+pXWp9gvZricvmKbWGjyWCxXElyo+
5owumstGfxK15uwVXuXl63HJlQ0KkiZ9cU5/leDZCfIkB7LhlhUZKzMmEGvk9ynCYQNq3o7nN87A
xFUis42dQ3e+eOXiiApxjZwKe7Pa8TQW1eMMTJNOqtM5O78qOEXB2DPh5y/+2Od8l0IOh8zPX7HF
PSm5PEp3vA80AbP6z3jnAD0Eec9OECigBGnj3iAUkAQSKda/Xmh3YAX/GS5noV8kQ2CnOl7Cvp/R
Tr3V+LRVGgTzmR6sdlhZoNYXm4dYlZy422lVUbg/rH7+03Be328aWCbGGNC1N6fYUuR8geBVLmCQ
M2ANS+ua0fL0rOTxBGBGOUygx9jb7a/1+MS8YxkWtFy5P+dEFgjJqvsGT3S71AQJ3IcJSnlNHs80
whI/6acf1vwYDrTWkcA5Bw4JU3jGhBtSX6f/EHYRtfnf7ykA63aMSfjy+tIiMQCX2MhIPV51Rpl9
LiG+GOrOrGwmTWRrVKrRdgYZ8Np2Zd316mKY5pcWX971FfXaJlz9YkAP4aYaEOyLtRc8sqq4hV90
QCBLyucHb5uijxRJCIctNMkKOY17tt+T9raQeCjK6Dl//OjsY3ak+QmwmONR1U6MzKL6Z9sp+/gF
fcXBagqRNPpwWg9rjPfr/hinuOki8fkZ/ZAPckrwGcU9yr9fLoAkzJeB6T+3+jtIk8pryWQeAEDG
g8NCVltQPmDMncDPYvpVdoj6wP8uWbAN4gqdyJ7wlxA/lmQxwSf5evAcWr7wAE2mwDS8VGt+5PlF
ZGxmTbjjpsmIk/XjZ9fET1fTzArTYzSFE/1QA3i2JC9Nho5V0HEEzt4nBlSRxBlm+zg0VTTBxnZ6
ljp2MqCjHkqbcQs1OV4Ce/WkKI7sQO2OecWg1W+ID0E1zmsoaSuN1o0Tqf8hRvcAt6vUPnAoS4qN
fOVu/9GYZjHsAjdLVC/FO8OdCkG+PyKgs6l4u8GMnA17ttASoIevJfFsw/tZb2R6J9wu/jkjM30T
TJHvNHymBLDLiQsTz4bXs7kfk8Opr7qCMZy6c2npAG+BTti/xbcAKr+Yloq+2ZmFQSZylTlfMejd
u/e0JakXHh8RI18m/tcTU65FJyOZ+Eif03rfHXBACy0I3OMpFtx4fHYdXXkJUBpA3DAQOO2693dS
KqB55kV4v//8PjmrVwreJ7pV6hQ7qI1Eqt0MoODw/ig+uM/6WTTswCjf+9i4d68C95w1Gl7zxLIa
gIw0c1VAZnmAIPmQK+U01fiRbWxK0GRlRnDtOdLMeeM6Dv4lF6RInPinzLzy69nWCJMm8mV2cAmH
BK39wmnOnvStE4k/gFup3zDfSZ7C/NbI7WwlEP8sWiOWZfTRAmFbNp3A27BpXKfqT9vnu7NxqXGa
PIf6pMGguILK+hMAkzWdjafpkRisI51aQYkZ9OYzaCFuLY60PBEpDcTUIdyCw67H3QelTMW67eDE
FwExlPktjjtsOqMPWMt6gX8+FcsP+AYd8Vxm+5NXJ16c1UjM9QPEFnRt/MkMUlFFcYZLNdlNK0UQ
App7nl0DTuNHSsjHA+BTvL624J4j/0MFi166iDNkLNKEN4dBTuhVH+N/YJ1g+rU+k7yw8hKxjltH
itZ5gKurK0HdTUaEPkDkLY776nZz0864Dj/IVBpZ5nCA2l8HFvP0uNOnl/0bT1vitDNjjgqoQXRA
6pxTnX/zOX+ReDzzIRs/8fZ+ShSR/itFfgSURDFsy6GLnGE25AEy3F05TC4Dc6moOWm4S/TN7dM/
G763jwg+9H9lCEnjfDWjf6VmU1hF7jiQffoAfA20DysbDqcEGHzO9KsTQxoJVtX5/iYoxRlVhL1A
oTePRlBuqjAeZjmQN92J2NT54WegntFx3HaMQt82UmppTF0J8jz9fAwtufikpzHwGmYkouGrNs0e
hdeKFrgMsIIGY2ufJ3bY2N4pA3QCskkDgUMvRI9JV3cPw1ul455Mu1CUb0uoWR88h6+YoJSjnvX6
ULj6xnWL/8jO1/Jm0XE39hRdglpmE5VBK/1gWPfULM+36c7CLLkfsAyio7MqYqvE+TacmkjQrlPw
7hxaYepM5pjJhekft3cjB+Cfm34J8eeCoXoaSpL2wogAzniMT19JB4oHU/bfXhfztqpbp29fllUq
xKVIqBExjTRiC/J8nXmYjeABW3D4SJQzS9JIou1xorB+YCORsBRXMKU7BOZwKXqvjpmjhHtoupZu
84YbbOPqypFP5RyTS5Ay1rWoM6NsnvtAhNRUAj32/YQa/xex4iqP7q5beY1thxXgXpJUIDJUEDwp
kHy3Xcv51U9WMgBOX99/3JxVx1oiKvFaTWj5bZSlWe52M9LfQ49nZGw8+dgAiOLKMGDGT7Bbctq7
ivgrur7PXSoOmTypmilybIpLriD8WZkvl2P5ppJCeAVnD4RXnqwTBV9cG0mzE1JXDg9tg/2L9XNI
0C1Q9qv8MbT/2lmp8JhLK7D8aqzqD1uHfrG/jFDRw+zXK2os/R3OfVI5c5j+x2K39WPX62Kx1ee6
q9QdL3ghIbte+vr0Bq0JpwuyZGfdluOAbzXrWRa5wOzohi5yRZGkmu0fEORzMfmfhPd3IVEwpoJl
yrpfYQKNguyGd7cSdwN4SZnH/GtRgVXHjugWnnbD+gmVSpDVp98l0qhzQkul1lfWIIWwYimn5qkW
jt29Fwbrny72UZjrzxBux1W5p0JtHUQP0vZT90oAbjeT/WUf/7USDcBfjItE0sogEDKjAXNUVej1
JhS8fYWj3Zt4lmwmAZ1W+etSJP+HGHPTvZ0BDBXSDXT8pUkY0h4XvHD8UWXHK5enOugsZxIQn8nv
KBQWOPyfuSMSbhvbmAX/jbm9mWUj0sd72J2kyGbPMWXbixOsYSPCSCl3E7aVNs3SWX7Eaxq9xKPv
X6X16IHpEhj3j9PwyQygvkzzNYhdxLJlid2A/oJfYIGxVf9i5dfIgtLh80H/lGYrk4iqT7w4VqZn
WrXs0K6OOZrU22zkE6UN+gMtU+IVDidtYlp8z1LxsYWSOOcK0rGZp/044b+0S2EoDdbrGngzNzrT
lligz+kWNzC64kvddRrt53UvFZ1LQpnRTuz0zqnbeXuicpi/2QIXCr5R22kILQP7jKvoqvHSxiyK
246ZuSkVvvCVDt/6vU6X9PEr9gkEN1lNwTOuypV/NLHAWYa3RfB6j5H3EechBEWRM+5Q62L+d/Kw
DlLUrjsKrapSGBZBgLeMRTCL4ilqlzEa6x5KAsYMsDnlyaqeTuy6F0LFEH1CFstclVBX8OJ/+yDO
Ws5W2aurs9Or2xnmtBNfZYjGp8LoJTjq/EaQUav0hIWt8ELTUmViV3YUZB3JhSlUXsd304kq+lOd
AscQXqRUdzGKj4ofokGtvOIr4hj7aSpN6S6CrW2daGYC7HAfi/MpALSicLrFNXog1yAfhXEIH8w0
rPLbqbHVmzQ08usc+oTTmSe4+Jo5GDmDq3tN9yKo7AIDEFXqRtPGDYr/2sQ81go2gzqVUmMfGvxW
rNJ1h3YwcOb6pVpAH33Jq/MC1PWWXAww77J277Bq/WbMbWhkWoU9a/W7Q7KQHG4nNCOCObOJblMi
ajqy85WbR2aNfFlS14c6L1KE/30/TcPqPntFZUyDnVGCyk7gB70fu9TLYRmftylV5CJw9EWmFd4B
AkXk2g5kv1OUlqTYSWe1QRwP+dVNsxQk2Ds0VrO1AhEgyl8lMn5CLol/SPDzIKaGjyIm1jcUUma+
odVekPTt/4juBJyQ6xdGHD9oQYX8RvvV94nZ1rx0Q6ajOoKUtSFXh3lXwty9AObzDeFZAIhOEFiM
PN01sj6Mtr9FT7W9CL87CkjAE0EuBHyMiWasStfo8SYlBuZ8VtGxySwBGN+nWh0lE1GxqCAvgVxc
JCXfJ8tKOiQaQzACmRahyv+YP8LfUIWrG9+gpIudOPISOAslxAlDQ+7yzulzAqqMOY9RVULP1UBu
Sm8I4yop/8zm38bZlVRnaWRWa1ssA59sYP5XqRi2/UNDqyftMAB1eYB4EJHuBI/ly00jr1aRSnDZ
aJvBlj1bRVkJ8/sxfNFIJ78Qg9gTNgf4DIvm7bJot0W/+Cn4AclxOo+dkoOQj96+CbyTO/ScLsA5
FyOmiwIPI83ck3qckeYuY356ueANtUzeyu52yTBAct+YkUHDP8QWB5fzLCi8kNWAWdlKAEEwh7vI
ALEo6UNB1KSe1YkMcP7H+NDvffuiq5zS3dLVsPiDMCLEexZFuXuHQfKMIfsy1nmxqojl+fZJw90R
iM+InUHByzHMvOJufFOw+SQWgt5Alktb3AHOPxF88rYHqpxayOv3MPEWDq6+M17Q1RY8qJaRfht5
9uCK+Tk08F9+wFeXS+PKOWyYY/7UKuHGmv27itHMBg/MHb5ZyrXCCrRdG+Lwpydumn9X+nGDkpoT
fxytX8+xzqSmJ+g=
`pragma protect end_protected
