// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:35:25 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
GuhlDIADd9kTXDp5bwKYIXGsXmMtsRHyG42WBdRlBrOwuv7YTzyIkuLqyvjQSkTm
6AlzRVNIlsS9BqnHsVCkDy6GR4XkP+/m3NlOVB5D3wWnAkZuk2Xkc0ZOCVwlNZkj
XMmjLnSzXlIv41RmQAMpRh18pzdLBC3eJ4F3ggtfIM8=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 9600)
+498GgdgOtfEiRrJJ0ClNWkfj42EprZ5i7LIPa5RiyCzE3oZYgUaXftwgIOe498u
BEtg6nbYZWCjhJ8IQ58EmjybdCBxS4edWZbHorvWkrbaH8TYmi9DWUtYx1x356rS
Uhny1+oYTxFDYKn8X1XYM/Fe5BULIRtVRROSocZBWVA9h32Cm032FIKpcSVtd02X
pePi8lQ67be4r51OmcFq/l5qwfsSGaNs/o9VxrvPWwk+/X/TFMPHkD37w+53YbEo
f76LJeA0eShUNU39be1UU9h3K2GSm8gina6Hqox1P62FLn3Z8d3DD+TL4t1PdL1I
Cu5do9fDNLOoDmAJ/4+b11loTDsQ832pZe9i+FED7qnDbkIkBTNWBRNxowqlCm2m
yE78Ia2MqfAptcYRRDerWuwAs+mwjl+Coxl5q7oxEPzxyvORoJkX4KcKcATswznS
oyIa+UhskyN5uuTx4wV+XDjzCbRlKFbE/PhEyEcFXrvRRPjfkEN6uqS9dF1UWpSd
6S8NkMT+7hfty0vyuUpnNHTAEt2hJtxWRtOCfp7gHwDRXsE7CC8r6cgQ5u1xakLm
KeQm+ojgMXOgM4aZVn22+pCY+dJroF1pEG6zF0DKhivnc3Bvynx41ivey9J+et+k
vOAiw8c8IXOkzfpBiDucnuS/xBRerDL7H8+EHEXu2W4Nqopq9dBXQWAnnA0pXG89
JFdOlB6lM0g2QSOMaLxQcRYIlUAbbUm9psxjrWvB87k/FKnNpcYXK9VPR6uyq9fG
X+hsljSf6wnx4dHvYCroGnRumGA0G6JI3Pzou7CgtVVJJZK8daejy31jh0UQj4X0
zGT7/Mda9/kvXzIBHhO2sz+i4Mv8lcB9jvSVfs9Oxj1DQ2QeD8qH4cvNvnHFpuf7
W2V0Ol+btFlHZh01OPys3HaxpAHyBb4E2+8OkAlze5WucxF97CEKkSo81Glltcdd
SIe5H8MpN5LXQtLlCyewIrmwTTzbMBHLXPir3ZDIyL5FUQD89KXYmFnABUe1xwH1
rVu56WhR3DziEGIPqHieLNFgUjfHrFnCxKwOMMgHqItB0+6K5NZ8s1o1hQdt3SzO
JOpGOOK+llJS2iEvBH7zmjS5nFlvXcFIfwY6P+01SEIGnrE3NoHbuNrMAxZqCjWr
2Tyw8tVJ03F6S0qZewLXPcR3gsBf0lyOZg2XbfN/HTUc7KJnpyj6rS/i79xc6Es3
cAXTI2bUvGexWa0lAev1RfGK/KzAnkTbFEOALFQ5rRg3sxZAgqy45kGoyyKRTbo1
jzSyTBr77aU9RWs6NqsQB+m9UbcHY1U6XQszIvIqIOBKeaankWHcK0oHhpbpedDo
cfOeeVoWpCL1wgXIMbgV+jk2LjRdEBgPUt/JQl7763s6r35u9RIMOTzfgjvvZ32z
9UoHTxCJAnOdwHiWDjH0cwlCOyQ5M0sL0LC+BrpwMT0OGGNbNxDaHOGXc3lQcUJI
8HF9baAVg5Pe9H+DCFUerCzcQD0qXJmIFva3ErOIGXW2DkJnzOo3kBRAqat6pzfG
1hEab7LV3kbphqu9LPPCeRjRqSEPCxKxdy5OvA1s42R+q0dxDlvVWi2OBlXSIO6R
tMk7hsj1nH6ABUA7appPpIZEhpQwXNb08gKnh/kp8knmw6Eot6OW89SaXKti7t0E
PEBvKGORxkhoiQs3eIFHTJE4r/1fAQDqPuPSsiOjB8rFGzm2XowQ/3F3Cl7Iv6gJ
6zNxu2HBcTi+edl1FAm0YglhuElONeREP9g5tn5GdlkIukkeitnBuTTpufA7v0T0
9gxlNb/9p3IPOf9s+Qw/dZ1xSy056ZH/+55bHU5YZrdVzGkLSp9tTB5Lm5S8vG31
L9iX4JSsHqVidhMABuiKZeJWAtamgFZEtY3jc3UEKI12ktyRYOFcbPB9Bfo4bPo+
US8FJu68MWzjBy8uM2veRtIZ2waKpn9KB4TVZddLYtYvUW0TDn6Yr7spI4UDhASC
QF3KU/E6uibVxYVvomu2qUNW/XISGfO2mCQnh60U1BeDDMRJ+j5a8ZHEHYzjJj38
VyWS3oN9k4hkz8hs8KmGAxQ9JB5H1ae35yU6aHy8h/GG1BSi04YDsI25yIGqqDce
xFyOv8FS4EnUnxleLH5S58pE5JaO5bFduINIgBR9OAyPyJHuXAOqbYbVO6CFXrT1
TcBWGqmcm+AVtqa0Hgu8J6BTXzl64j5EXFOx+aIaQL+VKqwj1ns9PAuPbFs/Jceo
czh+V4eqmKm8Y1ez7qoVLKN7eyhzoXyqR54R1rG2hv+hc3XzAwnOthJfzjIJi+S1
5YUBhCMIXnA2ZI9fVY8pVc5hebT4umVom9Y1GQkrE69GbtfTSzo/38jDauYnJ/Kv
oDY3y4oAj9dVGaui7mKNeJ8p6FC6xdTStJFyvqPL/7aKkb5ho/+Xxcw9h2d7cwyS
y7DovQBhUT1nhxKcZ0owcK2PuqRxFunLb9DgCuPx/eYFU3NCls4ogir+/sSTxuSa
WqfSz1L3OoogHuCmIxrNpVU8tV39gAfZeDAe+ECD2CP8zPg4ANRvWhi4JWIDgOAP
GmPQgE87QGy/s3eDBuUN+7io5knWGle9v+G1F1LpER+oDKuav386YhFGFT/xLRNK
N5UNMXAmoNFi3s9gkDxyblQaVy/xWXjgmtNIjQ2jeTzZmK09k5QKQqXJ1VS/8E1W
BTXc267pxyl2fOUfzKJ8gXsAh+GOI3D7iRbchsU+KhwVrquHBkgXojYOc1nYfZpI
DrkKoyqGsV7/IKR+G68kcSrc1Z0qJRwSwKLwQCgl041bg8k+IOdiVQrhPf9W4Dtq
+fGScDBg7BLtWzaME34AnOxWGRdcB89ee9ecszWqdOdjEPK3rDjDKjPP7MaLrtLZ
DjTTm4q3FPyx9VXCtwtySRrwiyGeFrgE4Ph9wvV3ZBp8Rm6UdoBmqjy82NSJzTPR
EVHbOcHKk5gmqAu5QeyIseldFpT873fjuTD8/A9Xp8M/IJXf66zlFnAMWUFO2b0C
AKtwjAFfZDr2AVi/Cvt6j9+dleDwgPADYMuPVZITsrMGWeYKnENnSI1w5f1OonWl
Bjo+CsSzPkmFPwsRgLqSh/wU9TmbbY6L/CIu/uOuqdMC6gEaZi1H1wov/zXAJUKb
MZ75VtDgsWslCCNCxSoc+Ptx2TiKS/cc0HIbZaadKbswqAYEOW06oxbUROYRI3hZ
MXuiIDE9YrgsCrPa1+NI4gWWUKy5ZGxNaJjO8LLtkv9XT8WCkrhRE2r4u3Q54IJK
eAjp+FYgymFCbD/fj7Plvpp5mXkX+UV+0lbdU5cZjfEq5f4cDNcRvzkN+ZhtM1/Q
JKxiuDFDqSW8/VP+ZqvPe/UKjBhLW+cVEPDowiPAztYBPYpot+a+wW9v6fIOJWUG
Ir2hW5jwkhyHT5gZQV+DFKzUreQQaSzgRXsrNe7X1ivzkKpw5xA2WBORqHvBHyJ3
5f94TM6UV7jSbh2AN3fT5htxgrp4c6RCDo8w3mE+7NoshAZkzu+AIihrNmbnEZtF
JKy9pCIbSOFrYjQ7x6zYQ2/Yd/OU+OxJrfhwGVziSwijvHfTTVFq3txvNIqRh60c
4XI78mpIVZHW1WCCmFWp/RuoFQ80xFdXr6nWbcAFEVKctvkUsU7ujyr8FjBscXe4
B7JxoiwXnVC6HKgcF1KA2JGGjuWFysoibdRIDATdDyztQXl1FqjTaP/AhNZlNE+E
jNw0/JrJ5lxbSH6NfNOtzJdnl7Wma/+LQvcX+7p5T7//NyQPSd6/VhtTWffn0xta
eXyZW4U4e0eVPVwx1C0CcceY3n1rcqoqPz4M7BOxRtINDK4JMeL2SzEHzqqB+kSI
wH2KyNuHzt6H+fuAb9QQb44wHM2yDaT797j1X4FS7NNiv/ABzqXzFIJBYnUUXLxi
MvRlquV0HnykroobaPFk+VttWJNAp28eqVxTEG4Azc1xOedOXhnPmi1xM4CkcJs0
3tNd6ziKhc6HPAxYnVZx2Nftqwli51hkgvumDzb/KQ7fgFjgTIndyH6hRXE0BmY9
pZMqHW3UHxc3TWYOh168LtVYXMLEhOJo4zv3XINRqsjcKUhu923U+qJFqvU7lJPF
SXo/yHvMbCMJojtOpHa2Nj5zKEludO86hEfj1WgT55sjnukz/tsMYmwq27Ny97vX
bioNuD70petA0CT7VpNUtvjTrT3MyvcCt4GTboxIJJO2tUVVfrTxjK1ohpmWHr9J
ypoIZxMlMfqMmO4QMIHIu5+4E4ePBJknuIDB8WMaAVt6p2FjLoCZTVr5Nnxm93Dd
zWtVtyOw1ktR0Ho/goQgImVXB5Qcy+A7qT7/5IaLyAsJRHqwFYfhqs4Ho4xl3e2G
I407ajMMAMnS6XjTf9r2BudqdJkkh62MrcO/84bE8P1O5DL/WRQnR8STN2m+3oqp
oj/jvDLLwOXcneJRNideISqwk450KVKeMahKt5N8d1mYrzcB62y/lE7KmVNnBLqi
/ok22+F+3neILrtH54UvN9N6v1r2xhPg8I5/ZDLRbwMb06cBlRvJFuLNI6gz6HXB
KGzYuDPkPh3uoxo/pDybjMnOxhQayxJRyHpqG7FD7zQ3khqhtCkWu3QBKtm64DS3
tyvnbnji6uN0qniOK7isVQxsR0QmrYQMl6UsIBMNz690VzvIyYYfv9crhIF+7leo
iZnpSjsD640fMZz4xX2/iY8DDppbfQZBTJHoKc6tgJKOToWLS1SQ5M3GH6vV2Osn
ouS5d70IO4n8n1zHzn15ZX4vgcGfx96pXdb27nKkFTR9AhGQxVRvjEVxNq2dg3eF
fG7z38x99mdqsgI67bxfNm/E1uZC173/m8nLUkUUVLPpXLwa3uIQRtLJX9CaeDHC
Js9Aeh0VhIxM4nzOQY+ChZommdveqnHiuj4SFvCtRX9UOW3NFbZywORKKJ7TITVJ
k/CSv4KIBJd7qJd7bMKRNJL6e48yWM+Lp6Sb/crEBm5wOoDsLvvR0CG3+62vpWO7
OXj0/3DKutPvL74T/USiW0W3S4BycyO9KycY+Px9u4/e2rgRW6hcx7cPluJzFKbg
TXx082HT0c9DmmBD16czwyyYqfkPzKa9j588CjH8jsWciOugctktQAZdU75+iUf8
y5p9N0+Vu8zANv8HkslQ8ZUSuzFmyM54khBAPzsyDMGcl2ONY/9/iK59NPdzvcGJ
NeUbHiptcDIs71ymc/eC7eg5dXvnA+b65zMp5BEULVqo4xrMNyZzK1riVkYCgNgM
b2MDqzjTM2PkdkTFRoYqaFWgaU9uS4yiOw+PyOXGCkd0dgPrdxyqziBwbFC5Fa/C
n2q1fPc995LxwGrCgbR1xqD/tz5NfiDpddUXjVUo5C/UIvCd9eDW+C6nTsA/gl1v
0yzzxA1ba6BWqu/y9gSwQhOLTYMd2Exq0XAehGSlarHGRzNCtonhbOjdhsEuVurR
M0dt+qITnzOYMxvCgm+elKhofQFUxd3+Rd5oCX1xPv4PUMFiepw4OWmP5Bu2JUvi
Xfvg3P6nomR/m92bf4bNQJKlqmHVgBxJrFVMAirbvRjstbwbefD98mwb2BflwcAo
yn/69vywL+lPqdgXzgjWtdsyd6UFfDMCfnTpBNK/jxiPOoonkYN1nYat6Gf72FXg
yWoujN90aqwrbECs5YzxulseF2EwV8zHfzs5X0VaAi5ahb6v+CI5+bchAuEesgia
cDBU/VfHP8a7FlTzRwFbiYL5NoEft+aYuGblitQRsCQiu2L4KOcreUrzJbP1H+sc
a/1H2MXC6CULCBhcQOFkOOVOKaqNKlIr9TeKX5QbD7Oaq541Db6Y5ZnREc5xJno7
F6+tuVtkcDOZdPAGWbAQU4d/V+CcUcWHyTNIm4XiuKl+Iq5EjCbuhPgDkzYsbRU7
keXwOP9qMfFOhIXSNkeBnbagwYJ/roEJ24tq/nsswLumtTbCeLewwVUZ/jAnhbXI
0d3iMjBt9st8Zi9rHkmhhqg5ldJGrO/1ZAXxt28sLzXR3tloe8f+c1bAAP0DQw4O
OIje8xI/EW9mqgCGvJ4MaK8drcMZKpm8aAghrq6MNTxuWllBGwIuXzXwCyhUbwMv
pUNS32dVTNf6P4X9WYLIjPjn68lYsLQTgI2Nj1Ywex2KlvuA1tjADp5v8/pC3Kr/
Z/DmA58NFWn6nLNSeWsPonUhj7MmepOfcRWbB7zax86Fkb+UAHPow+eK49GKIs99
9yfLDmWAxzLrlA8GPtcZs7PZ0hiiWKzyzi3nY09GReSz1+rG1VAN8zk1x2m5xdpg
z+O5Yg09UfkbBHM1mKIf6uN60pECvIdcqs4NKorudc5dhNPKMpfhM3/4dx7yI7lV
VeRt+bhDimox/uOK2gT4usPTa8eemli7r9E1rjvKRfAqtGgixNRmENwzWx+XAJhR
MzabRTPnViTeK4uzobQ033Nl94XLvZp6D0+4F3c7t5EPSd6HEAdnHSjEuz9k1+d/
46+6qRHrcJwXz76P9h7LAmAly3jQ+76DQ3TNuYUjrhLkDbQthStgXFX70WtICQzq
2Am4iq5+G2gGT7NzcS3GRQ2WdyxnInxSlpEM3NnC/reanMeBpmXhyP68Yu/WFsZ7
/kv+YPK/csxSI/0YNkN8BxCp/m1NAFUstkeoa1ULmgwdff4YLhRigFbAeUJp/zIa
y0pQuSdIc145CdttjP8Mgv8/rtlBccE21A311L50BeiOYA5/hZ90j6aIxaXwYZGf
yHgRs1hDk+zX0Ebq5UiYMrLCsbTuQrzzORa+Vo2jr4WOE2P1af2AYcFVL2NOF0W2
x8NYacLDmAUoKwrEsmko+h2KZF6BjweJVfEUE114Hl2j10IgUxgUduphV6gkQtDt
Gf9cranVIIeI7OxjCvOlw8/fPwCnS6wUsdjaWhuzQhW+WPniomLbxvxclkrHbnou
tG+UyqjFWbMelTUqq/Z1pVnGVrBPhF8x9nt/fRAJTdQoIwxnOSpnPDWzUKo9Z6qP
JXgc8fcrpyvmNyprBfoc0yQflc1qbWmXFkd1vABLakWYvgLrIEXEFV7IRYhnl4ZN
6z4pu3SZ4UwdggcNjaQ/ymsK5WYTGOjzjBuDW7RgdAQTK5dL/kc7+Jvubq+mJ/RI
8txWGLK5SFbvjdH/sWP5KFBNT+jqBgPgzsmfH83Qr5HDRRzqFv1BybSilKgpWxeP
Dr0YqgjgdaO0YiuReEaVoB0yxYz+RTe2N8JZZPRgxACcwS+5OJFomI/w49s9Xp+W
54Gkl4IuZsJcIsvUA8WZyg1jQ3d15IzFWL5UvaGdgx6nsLjwi/UlfU1k0Z24G8+T
Z27xF+uvGY6y01Q4ROxW8CprJp+qZQmNKSRGpLRK16v2IcEDGxxPTJ6mq/n8mPZj
IgwtSNRsihP6g1S2zHwvHVzN+2z9enfTu95PZGQKxZsRW15k3dUQfXvdY9zY8uQy
Ho3ykQObsj8js647J2Si9bfpOSETwj3FMd9qq/rT2qYvoCRma4bfk3ZETa1LvFpu
6uAiyqtilZC7NFhX2f4/d6LyXiXsmXcjZlpMtpuWZj0A0pdOGhKq9OHUP4HKwxtR
Er13p2svKDSsAJI82pasAXbF+6wFTtgROgtHQ25rT0mvK7VwWnx7W8SDZEkGJ0ni
Ox/sp9NMItUiGik/biGLWaAboiq/KMP6/OrDFCcCvVjnttuwh0zV9Z23wE8Sro71
uBS07OyX5sZnMc7NyvQuz2uxd9bNiNrUZ+ZizCWUeHM7pPuZaij0YO/3JO/POp/+
q6WvdtkZ4VtugMsrVQ0VLl2Ptr7RBsTkyi3ODHXP/tOR2wV2rorpLs1gJHCLJ6GN
LG+8qMs7iWP9u7RJjtHBZ8rMXMhGws9D6J2oQvw+mVD+38tnPhpIVBO1mcNXGbef
T54lRqNW+ZjzS0ShUi30kQhMidorxwB2ynf0cgltmps5d8QCqgBWcMh3r3jp92QR
9aq7rsfadCdk6v/QF6M1voiS0PH99tdBVLuAx+EuOcdZ6YougDojyOVVyaxvXKCV
Cp193+kfTjvE4jzwvvPue3a8CDJ3tqs8Szv2o8loDtpATBAb90F+aQqy7bbecpNa
Z2/cZse5PxNFtV5pidbCuv440fU8fRR+NYM19sowmIiavjmLUu1/fWERY4nw8SRt
TYA3guCmei1yMyuUhJGfNd2CYZT9npa0gdI1N21wWmZxwMQ4s9QycThLurxrDVvj
oL+UhnzzF5oQCCa++CGZpCl1+dhpQ9bvu6rCoq7mwFOxnWwK9UBNI/dwViMHSfCM
8g3XdtfwPZItP2NlPc9WAbpVvdRhnv6SJxZpmf0VSYm9aoDg21mkxVshAc6zXMjj
FK5yAAx1cisFlndgw/9R76SUvqnNtYQv2YAui0bOxbNGZJSLK6PJ6TY+1c4otXfL
p8ZT04vFJxHzXQZ9cvjyV0etJTW9Yfjgy3I17G8IdCJvW+41OroHLEB/bigQCYNW
+gqMrJ9uYztU3F9ipWiGVhhceGcBXxWVYmVnFDLZYUbAGq8LxKCAe+U9e6m6lVBX
w+WVEuXtc3OKp59HBRzJ99hYlcGn8Y86CzXrcx3JfqYAeNCEzYoaN9hYcrv+0eTU
9z0rLUlf9tWvmYSVPCt9hMGg8gY2nMA/lRLDkNSS98DcE14/rxaxNDwIzrfhZdBz
DD08j6g0nmRM0GP7P8fyZzxsosJE5QguqhHHG1vuMZ9RwReUNazrEi447cQu4I6q
d2eOxPPQh1IkqEqhNFiSRa6ShKWsxtU5Rmb4H6U65cOK54VYxZ1l7NL+RfYX+z6b
sUEy8m6ozakhKwHO/7DjVSDGRNMcvMJfGRnD0Qn6jKDr4brdDtxJkVXLNCmN+Vgp
UP2yKhSILBTZ21HMy1639tjDKgFVDZA6J41SljH0uSxV5fzblVhItUBUm2BgBze1
7hOKuam35ONycP5g+GvoXy0q9IZNKnGUtiAMMpYsiAFLbK9aEcxRx7z8mYZqyt9b
uLZ0nH5xMn65AA5pGNWryKn+65r1koy3nE+nQI9t4I8nlx27awqCvc9NVkDgDbF+
x+Gr0z6e1hga5UlBgOrdM9d576GKff1LPE7+W4wBFt78JSNLLsCs/wsXPQxBcPZS
arfriceAoZ4WhkAW3KJQ+ACnNwQksGA248+6tahwvWb6ICd13G8B7LYldlFK7jfB
D1XAsEiqlC+t6FC/DiOqqRdcpJqTGMBhvYOk6kUQLBfqup6XPIMq78PT+SEDPXPQ
8DqAX2SCKKliJoygpf34LiD8z/ZmurPezDoorbiVcl3jgHsLrVe9iIaV8NHNaSnt
WSzi582hdntcDaEagLRtDdwVSJ14O7xzMicBUL/XdU1b31pWlAHUEOECuRprHNG9
yz7GKRSrFQ6eQPV/eejVKSSH3vJT+Xnz9X/LrXcpmRK4OHBjb8WdGLxVCCSFYFuv
ul4wbZZvq5GLoda+7mOrnEHw90r/iox8cESetHUmw6gpJCYFvKx2H6pqo5pRE8AW
akJ9OMBXaii+ERAryeA+3SRnCAiZqu4ZN675f9nI/o4TNAB9p4azLZ9KfMaqWrG+
uQMVQ3T/lLIt+7PXlsALywxaa/57lMt3PlmnSaNTrVkOs63lJI0q+BLeQ+Iphu8x
71uPyWLqLIm3bWQxnSOv1CBRtiNvADLGUI03n4tvt5fn+bPM7oHEoPzD4IWNvbzZ
1iHjRSFulzf2fVc/zPI0daCU1aehJqwL0ck000bx+3exmlosc0R+kdRsXnR+iVT8
F4agox19SciLr9/+ACiKXSNL8TZleOYZfPUnPupZbyN0bEsD87DKa1SGuc0E5UD7
K+9zkEgE1ogmfn/FajQwSiNKQorEs4MAcURR9Zp5yxeiWXCkOdaAnUrEMlwwrPb7
7u6SUWBeoEYSr2HFBQAZtIiboEzcJm+eZ+9at3CBJETCXWsTA10VyigOgitvyhLR
r/aA4Huc5kPxW4ZxHhwaZEBrlDYte4f+O3U2C35EaGf2EBAx2MlS08h6BiokIeOg
EwrhJ7LLJo4Sz6AO9FF2H4weaV3Ts2XLchb2TdPryaBJGc4/HCkUM0WAM7DH6D/V
hqQt0+VVSyZ8x7uxuN+6FL3C2LCMhWZU82eDJg3DhBr3SuhJHtgg20j/GjZx7fLc
XmfKBbz/0G1WiQv6fPoQ6dUFd7xGzSUqGB8P+k23bruDZ+QpP0DhwmSSCBUdC3/s
i7IigYlzQuBkv+qVu+vcshai1b5UfWT0VgZL9nO9AMUSNA2POHuEVqDVV4hBZdMt
QR9uOKMO3fD+z+Fkl/8y+O4BsoFGUveJGJq8p//ekyGuNCUPZbeymXKudUK8iVzf
VHfolCnyE5HUhUhDOZC+7AWARanv5/JMgf8MWu+vgu+X0v44ZLPkR89VDVspOY4j
ehe1XtIuJm7wT6jyT63re0SPOsNJYA5EFXCh6bmKD4oKBwK39/s2zbAw2Z70RZzZ
eWdSyOjIYHYSai2+GCQcOa6V1OGNcfIQiJQFeEq6Yh/Bg6mnItZFC89FOGH+Rjys
CQIofjoXcV7X/1MUHmMh7/ALFT0FyVrf0oA8Ee+VuZan3bh9sex7dqHs8xhTix0R
EIS8PlJuS9fQhlKHshNyBt1Ieuo7NXddUM86eXHvpeOCAJZ0y7bE3pYS1dtKs0Wp
HcjBiOT+GPkjWinbDc2CyCEloJHxqSh5lZ0KxPFlYoXiZmiA0PcG8wlxkD3AnE99
W6cxFdQ38iuOznklPHzZGsldWBORtSFMN6N9XeN3bi8+Gdgnb8o6DePBC5VSx8VQ
TpLNS2bGaAJMSnBenxprMorF/hkTUnrw6aryiqDo7vO19Vdscy4f09h6I2W+s2fy
IBa7RHjVczP8YPNTO7VtX9BPZakzEM1bq/nuMfFxeIQiOy+vJeAwZFuFVmNC/0l5
TfjYmfyYK/ddo42bzfLsqFt2Fc2D74ZTKVyRiDL/s5ALxlnYKopTELZ/jIwFxXA6
jvdFypCdl80Wv/E1FW8w6zZilnqHmvk1aOQq1AtnBbG5lj5h4YrVLGrXZAzT3ncS
Ph3yY1I5CSFIMVJXXlhaA1L6/A3LLCQnhI2NK+9pvNhwUKZjAb3LUWm9kFtbO/NO
QTtfFP+eja6rIr7aBdakQpO5VWBSVX6YabCbxfwJmVkxwelHjaI5BPst+qJk4TN8
qhVFBUevtsTuZpa0re+mbjgSAZMLdUdbgDSeO6N5LrDPyJLFoFVXyRFsQs3c0mqm
kTxc7oD1KFaQO1rFSpDvhyL8oQiHiCZ6FrKoHHX0n+asTQYo6cWCOAcDhEFggpuT
cw2Wf5ggKa4CyOGNiCpuj2bRIAWMS7fj22TITYXANU4H5KIZahvCOh8Irs5qlDmm
S/iCB6Qgt0fuyZ88MZrJjgo9MBXvxfjOp4NAywhwjN8Ut/edRUYAap/KLxK/kUdJ
2dTfZX0Qbv4m6zDmyNGjuiESW72/uQGz0tVYBbVPl64Me3TJ7FrpbZFQbkxEPReP
NnpNvcioNbq2+D9xhRwiYns6elwwyKk/PUzqVlPtP0pDFHHmyfgOPlwLKjI6Nnjq
xl9bAxHzAlkYni4cJo6HS33FtkLpCMaWm+5szb0HHqcAdtF7VSJxncTapJVSTrzY
foc1PrCPZvFsdeukb1uV+J/rgPuDmbkZIkaLpS6DRU3Bu1cGdzR1jODE2MlK4c0z
7u758hd6FVPkaZHZIlwsgcE7FAW1wsLIZFYSLXZ/JlMaVCsglKRaOFxDH2jx3tIa
3NKuyULUg8ISJq8JiVxLSW60oJCSYWvwenMqX1SUs/611RJ5IoS9qwirOf7cs3WS
CpMt59rFnpMoRKPPjczF5h9j1NHa2yR376s1iniSEsRBuv18f/KWtQOEt+BIKA1e
+fZM1Q2HXKqiiOmUVvQehQ+Cgyq9tqWfRDQuUeH8OmlcAjBaRtZSkHWsJE+omWGE
Q2UDFgTQUn8MOkY9kLqneDkVkQ1BNRRH420/KdCVWTuW51dc+e4lJFFpNDqY9ndp
+CC4veBs18cKSs5AKRWyHvBcupKW0Fk02PsJkZzMbWRJO4uPFcu9UJ9jQjNam7mp
Zg4Z0MaElDuEB7Rdm9TopjApfsL2d9mYf2ULogkipWYlC77qrp9/cNfJebch+fFL
88nDACeUHCjcT8N+7bA2qrPP5GAyMVCQQQoLESw0ZqWjvkzlHnsE/wOD922qU0dE
X6WfY1hOwUb7KMXnUFsDIGkhm6f9SDgBIPFMMFx1KMuzGHDtY8fNoifasj02O45o
1JZsynBekAQ6AYQZ+ftjKY+T0plWWVTOHSvWNysLaelhDIQAN/Eul7p9CskF/u8Y
Cm0xwa5/e/02/AJNE6pQbRTNQrBhv7ijBZjKqWNncdlFALkG24CfiL5EYUdOHnrl
AsHbMWmqRQCfj0IxEgikRbMSipLU7TScn1+gECZVMpQzi2XMxgufjI8JnNYDoUGN
ShOIm3QINc/0OeMi48ue8eXD8F5CK/Gddkkg2ZdW1Omkx3hEtPM42kZYS3sbsdyz
lcLPlbkCe2/nP4C+b3LBgpuZsGl2+fvRlkhQ9SQGqaS+dMnaDBM7v4bRGsT6w4fP
2n6eAEJvHCbGJ74IPyog9GluWVIUhCMq8kgoePYz44WDD0Y11nacgfOjz8uEf463
0zeES/xIM2OXJQ96vqRzRzBs9kA4w4bNqlegJNblJfNXGiXBVzRKMka6MEfARLLu
yDES+ywWxgmFmjlRTj+f6+lPYjFgpbSG4dZBs//1B3GMOiDcq3XQfGcuOlt0pPnF
yQfyX5lEv0eRkPjfvgCVV5giAqXweOkUEa61LslGgiVILQ9xkDhHcWf7abYiQBtA
`pragma protect end_protected
