// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
YZKlCG+bpheNYl3ZUE9uQghb9hQAgp6xtAa45MSDXfGCoYQNFyJ/9dgjNDpYZdS232LchPbxUeL5
/B0qj5aus7cAoOqxFhjoQM7CD7p2qrmylE9ut1YmWgoJwhVbTPSmIOBpDuCLwKSyXoSLBjwAxZM6
408izEnVacrDSJ7xY7UsGNn4YnU8yCx/7wlWArTFVFFaox0J+tGinBw997PoUMDoRT1jVS1yncmc
knS+4qzis0GRHKbfbSoQCzWv9aDTKrLpiJT9RStaKvToEumtJbC8f1lkb0yh6MyZrUdVy4BJZKcw
DTkD2oEMDZQK38Bj8ZSEu77YRzV5svkOHoH4VA==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
yTnbWGBS9U7heo/CJEirPs7Oo4UuvFWl0iqciAFVruFpV87SrkdCQr9F3gxs0UwxN0lnjl5h6PBF
Ei+WKvdT7cQGVqeTKh1112XeZCvVUqweasRA+R+upSmd2qC1fOY7CGI+GmzlSVMfKHTNrdgCGU7+
qqI9QJ5Wj96ckQ9chSWDhz58F6xqnK+G0WpQK3suIypaW461IT5p8rV7BQirH8hB3swxDEjxpodt
UcjgupgRchbe3YD1BHes352LX6lV/BwKxf9BPiM7rtE2KrofFQ0CtRW5tGpdtqGNZH86OeeE/Fe+
P1ABv5V4k9t9OPM0YmdAGIhtanTYvmqKLVh1zdRjByV0kNhq5ufD4CYrPzH24ymWkxhkqK/IrQVZ
dZDB0yX7yhM7dhHzV3Gfu9+osbn+aPstEz6UdnOUVF/6NblKoeHcoicgX1EN/Vtv1KXQIyR7tN3F
mrz8yXily0ziYKGoQ11Vi+Mez05wR5WaQrtq++xhzIB8k6ZRBaCdvwU8RjWsyBAY/QM0JiNr6BSX
9Na/DZBLoGW9mPbpcvgJSOgbCmsvbTF1d5jpMv+satscaX4FQtqWyRDG8p68BPVvPsBPX7vgvY4U
8F5izkd+PugxuGNnubwjfw3yAfCQyHb1QGYDY92I9Vd8qJrcbVkEABgJhOMGaXUlLZDMowlY4YiH
45OSdnZNE0qc7lWXJMs9+b4TRwvAS78wuT4mXTdCPKCFM66BpIh88FV/KGx5DX4QH0siug7/GRKO
rtt36AzFgeil+O0XKGQwAtpliyWq1eJG9OnyMchNAMCQzli11BKk1SEWhUcdulmjy+EQ6oYqBqZ6
Ec9NKDiJqhHD9SVKX7F0HXTjnynsUaEFc47fasUzDnjngX275Eiaqdugj4dGvrJK1S21sAIgT7Ut
rO1yeysuTWWutY2X+NDxahw8ciCuHvPsE3oERCK3wSfE7aPntKzemG/kpdpGdGSjGhUwCtT24E/3
vanzIKiYZEiGqDxAyK3cu1Lca1m64tmBGvqIkYg+xk6FfCKYDjSxZOKJzf3Q8RThGHOcVgLElpxT
9aZny6a186XUruYnuF4pcXV8o6wtHHOtYyKETWqLUS4faNpY6ndtE6NCQOaGbi8PGZl5Dg922UhO
iQ0qTQSOYaQDz+CgRhmV3kHDFjItQdz2JuKH6ZuAPRJKcIY1Blml0alDjwQRZJKPBapgUot8PyKB
jeX/LaJmJJ/O9TSW2+2F+sxKxzOgNZFCS3FaDBpQFnwNgbhHBxF7i8tL+HMkIJ4T0WqYQiQs3Yhb
ad2JvUdMyy+dz64g85qMm6C87u/pjpc4CH2VTM45GzbgxTyCtQQMW1Csu49ABJwgQ6kAigjQBdWk
bzPqCMw0cI4wGJ+eRY/tqcJFZoL/RDpXJ76AjAgafj7rIxTUy30314utkWVh6AGKfOcqVDcU40pw
0rmIB5DoW2gZXONJS0rANeMEP56tKWkr+txSF6YTUt/wWukds2StOqIe41G5Cliw0i+QD2l0os08
wojNAPhoxV34r7EQwexdPW+gghTNUk9Eql2SsVZhV4qoH4P/x0bTOni8sRsbPcv7UpKeJoi7IL9/
2YEDTf2V+poDUW2kmvek2h+0lFSyowvYZYIgEfc0O5lsAH0mQm4CiSMY+sprmUuPDB98Gdal4kY+
SC+uDfI4hD2Qu1lHG6/Zx+TswiSchc88fidzjILGp1WVJjcI9x0jChTk/T67+mQaGN6lXXFC0Xlq
IGC4umKzruaXhJcWE8ibsHfkygc4LjiFbDb0Wp3sv7KH+6eb8SUYmRjrQBXwRXbAIjibyuYjQjiA
kQKf+GlbrlxTQGppZF6FTofLz4PhnaMwPKx+IOOctrreZcVxcHXCP/tQfZavEHrfCWhC15kP84fS
TgLb9v1UDhCgnrD/wvQoF6ETqo5S99ljh7x9QI7uNwyy+Z9TuSXhnPqAzRL3PPbKiGylojw2YaT6
m8A9QSrEuWClCAHwgEwtUbnNyubT0G/LDqrXCiMyBT31EUUp0QmbHzDR2s45br6FQh/jRucufB36
gbwB385j3i1oaymWmftIvH46SskCyzOiLSv9RlRS2Yk9ZJOxSefK3LuEHLWB029UlLPPTF31lJud
laA7/Q9Izd/lTxqzfVjOnAdIGRXJM1/o3LP/L9fiCzhlJqVSN8x52Ay8gcOMxySWHfKP2jvFRa2N
8Y1Vbfu8Bzi9rJIytXPQlE+j/ninVN+zaxHHg/FIj2NRZDhnRk/+FnZkxq5xlK8ei+ykcazKTEpy
O2D2eSyEv6Fu1EGImk321FV8Cur09vcoP2MEG96An/2UP9SGpcalicwz1Dfbr7klmEPPdRhAFink
5jfnSR/f/fWO4iHIII9yzU4TvN6SRPonMqQW6duZYzLKxrpVODDdKffCEVS1vZtwzNKrJ4ozssdG
o2SuwGnEj1lQByjCzwzwSbW0cSS0XicGV0EGZk17dgflZvYZnTyTAT1k2J4P1bPE52pWmQ8Y70Qp
xtDNMp6xZbYy0tKaRBYxGwifScLc47YjTdcCrTZtZByOsgneUb6Uxqmcgpr0u07aV31/mwRpCfYv
k86qmBYOrqbRB2z1HZlb8aAE8caxudiM8Wu/XixbQ2cgi6OVCc70CvmTIkwFv7BYE1iP72n90XI0
Su43E27vM4UAmh0415sNKqhbtJAQ2UWMRSUYXRsIHP1d4nTyAj1trOCN5Hm42HM97PF3TDtaC9jm
gT155HLYVU+fiHPtemBwkkMgdYbI3p4SHLrQz2BYzpBTC6A2yxBOeEDgoSFiQ7V1E859cTCcgrLq
YajLT0YCz/Ib0a2X4yHEFITN5pXdn/MOtsuig5sFHZV5Fjd5phVHYR0ttIp+ubqsAZYTpWLnV8hf
k3gFSqOo2eK7TYfSuBWdY94dDHKn6Ka1BEmdO+KTashMbcoXYyRySx5BeWx8o279bCRbUSCixMNy
CpUKvKllbeT2VezEFaHyFUpjM0kj3Vli3lRcHEFChLArk9tsNTNUxjdwUY/867BMHOZa9DqZ6njZ
3QyZugfvvr/aK8tVykGh5F+4bOI0JhqtTE47/U9lGwpBdq5ON21CqS3F73YIGoEUdszVZmJywWAZ
gh4/S3AcPsfwjBtGW43OCgrf4qpldXcVPQK7hL+5ZZ9kjWeKFC5QzAlep1waI7qS7O9+zTTD7o9N
+HUTwCnP/DhFdgo88IRcW6GT2E0TdX912eLYahkw2ELbtPE/57VH4E3O8S+LZFAdeiqBiAYy9s4o
rMBoSRmkPFWtGgKvv4vePviHEacLgS3r5+HNU9xnmsThBDFXoAZKHDhMALYxTJeuw8WVZ0ntLojy
jeYU1GB4TS+jkQbZ/RLiUkEE8oY0aGVoQlp6snWJdYZEl2ukB+TMcL8fM8eHeD979zpHD/ICHwWK
NFN9Um/ME7y+QWcG8YeL8NrVa7QIDgyTzUZp1kzS96FMxKQky92aHK/GrlX17WfJrj+/Pey33RAP
6SCPpyA2qx7vTGuNINs5UtpANWnzqYnBEn9/wbJkx2y9rm0v2ckQIMRzLBtomPULiEb0u9MH09ZJ
VFr4YpcYCzNNGveS4M0pGWIddF1sqEfAY3fohCC3fsbNIqLHZ7QoEsZ0jMCe11osG5uosjjNhUgz
UHN3nucs92vfkoldza6xgyvSalK+2AZifW3W7HMeXI/jPFSTFLY1uXCqe+0T+Q0isXFNpjZWu/Xd
ixGSAW8Um23e+6475Is8Kzz444VXBGhHm9Ulue64fNOefkBTOnuAXDjJFhcFrGcq7GznXENyEorg
kp4kMfCUB008glLf5L79FhLVJM7oxojLmexbQDHAEfqFm7RVs7ak+Vzl3/B5zuNp2T5h7IUFvrlm
w3Wbyc3/cizQi/5IUsvBX+MS4MobCyf+0cdkTmvqutnPtC+mNRTg2HFcarWre1BwKFN+hV7iM2TR
/GgqskCehQ6mckKhPRIhZ2IkVoay94luKjJPMaCzrNMVN+5C4rie7rZJvmRk5LV4Skwh8e+d9gtc
b/QjjyuS8r7RitV3KxqEhKj2w5uqWkjgsbSbzHKPJFfqLrgVSHQQB2cSa4tiTQLJd0orhmaEVIer
9VN4DWWVqX2UzQekS0nupsAZXG9oZG74puSYx8lbx7ftOsg/XhbE8AWpQeMmtt89Xny0Al9DQziu
rN9gZO/kU7R2v/e+BMNsi2s8IwfmDKHRzEGUCDzu/0H95yWwfbtbf+McrCbb0u9MabHt2C1c7Z/p
fKTFfUgazfdTIW9L2te+dG/deOFMZqH5Mr161OIwyUiWWUJrJT5vt6njwEfHwhwx5l4Qs+BkeYM9
J/oadiSEk4qQlXo4tSsqQeF8gBFAUaTfTQIjWSrD1Bc3yxgpemOlYdVgmf5GvaeruszBB/CLn98Z
w6SmDGrZaRSS84m/qIeaddVGRXPrxx3yE7L3SbNfEsObPAbyGb/bXt/G++xA5053GfL0i+/mCM4p
fWEFbCB4rIQW3cMidrH5DuN1tvTDvVqHMkL2brokQC0zku4jUpHcbI8hbBm9uRC1SHXYdxomVMvf
WBgszJtAsvqDeu6OnFDXIkLRsyusgvTWmJtH8abmZ1fcG2ufEqFadLKXlaaoL6bi5AXrbRm37YW/
LbTXqYLPI2gcN75XQwPi9ZqJo4TXSn94STsJX6Va2pMnrFcLQq69OGDMHDbcA6hXX8dKKsdDLqhG
4nq+RcZ3eGmcnsRQPSyGIAePRZDSBB7GAl2/an8Z88eylQWiaDwzxCT2IrfrF5bP3rbdM2s37AG3
RKS9VpVSLZ6FdXqtp9iWVeDotW5O/SuJcBSNGD0peYgvjHYLQVEc5dxzJ11F1TJXd7Vu9RSTpT8/
9+8Q/HnaMaoJFTopeK8YVLeOeh77Cgb1Dvi11SDTFgyji6sMCLeEn1tHS9WC1luV2VOVxjPrmNfJ
XkQhr05sBp20XYmUMIpcUN/ensLDYns6qcbVZNwhtziliSQDCvfrKa3FpZLQfTO9FIIrP9E/niLS
V2qc1EC6TehIqTzmp8Z89ChKF0lRKSGYtkFNMdkCPPIT/INjg0x+HD7924RvDRtosFlF73LGc7xe
2TMfS2wDDI1dJ6BM2H2TxbHnfl0DVW8rxr1EHusnQpC+5tjnAIAAGG2pohzug88xPjWU2ARN2P33
38qQ0qi1FbV3YNkm755HhMNh0fZ/3cKP3K9xtX8FZbTK7iT1hPHKzPv+HYviz7XYa7kcJuGYKZ8l
ods+a9xvG+8eQVRBa6qMY7ZBMw42WeTy0OpPK8cxCgQ+00ZtioLNFP1kFHP0W4dwo3xno8YT40LA
eomwoo7dCXq04CB8yvRRdVAIGNcAY8iyxYs8lwRfXHMNIwHraII3XRx8lpOoGCObnQriN/6LE0Pu
qhweev4j7ylwK0bJMlKZq3yd7Q5LkWi1VKfryTFi34+7BJSIM61lZoDAfGhSujsK9cf3BE2GlHof
ZSWjRL52pskcDBqlUVc1he1Ys7MAjjpnUCl3JC0PlRV3pm6p/EHUqP5Z/0nrpTpvbqB6Py37n3+z
vBFfhH++Z1Gm9CAdRhEmxky6yBArGShAQ2unRH4rRB161e8JOsmuvlgLZSQDhlBWen25umCADnm6
9IF6OilZ8i5sdhGZJb8kBuZLaNI2wTatdL/omPKGZJlnhwwZG5TDkAKPe8ZDDFQ8TMbPnjg690Xt
b8rlU1XVX82uMjs4+JTWrJyup+MsaIRLETTt3VIzu7e7aRYt0MVDeriGW5fT6nhWQImpToWnE9uM
jNrDLeNcQUZYQp5OzZns1LfgL2ojz8tHQs2Ccoh1YnRhI2yoedsvX10LZrLVT+zXsNas4GUFOZ4p
I0erZQRpoJFMbtCixff9Zlv1JEi2x/2qahaKjOxgEkLuXGY8UwotiJDOcegYpeTAFdvUowd0aYVA
I7VLzfHCeAQrb0OA9Ajb+Pbi3D6T3ZkxuUQBbPJNpfl42BtGaHjBPyr9qR0NZCPKe7aymxoEYr7g
Joj05CSdrHyWPoTY6j2YLwWH4I4DdDylctQDblyxauCgu/JGfIOTw/QbfZQGeSzjU2ZrAyNH5Bxc
xvqsQ6u3zhjIFBB71mALIUEZeGmUmOFgTbZbdWDXeNR8sXHIhW8WtfJBUydNlu6cqYdNYmFeZKQR
FRCK2NTO37LPPuXQPcRq3+MKVWee5uO5C+DbFpzm5G7MQW1oPXwa+npVVXImeJnx0oRi7fPTCAx3
M3/YPV8SxsJDUXc9lT+XmtKshL/L0ZCOoBhtDnCC5s3w3rqDEyL8YSSJHZQP5Y0dq6b5OoaZ4YI9
ouSlnW6ngtjlvj0Esr42X4d4FNE/ApYA/Fjpn3BPVALLs2o7lO1xfrUk/qr6nQPWENZkmlGiRiKs
RtWCKBxjoKFcytVzyZ8UD/1iMrFJ6lCu3piPEPHWNI3nIGWPuFGSpyLUTLVmluuvpL/JAE0MF1p+
JJQn2m5mjkneI5OaMpJDwfow+Yr6Vn129JQ5nQN7kkty8KY+1e/mpCWVUcPj7h80aFFnGh4D8Tyy
RNg4obQxGyOVH9FzSE5IvLBdv0A8QEdE74NVJ1+unBxiOBh5oKU7uQ12uqN4EPxYEhNG8Ot1HUJF
41D6NAd+RHnn4Ro57viT8fZHZfARX5N3iF5R9WhHOFSSXMVX0D4T80oBKI4HzUODJvA4x5gNJmrT
E0GLkAIPw/VMQejsuOef5h7PJyrqWFlH60EtOHkiCpkBpQLguxehEDgfkxqEzzP9ohS+g4gv11vU
mAXcw39Cwy4s/nJY2ZQ/AGp4xvgOPj5AZDrqeHHkew0VUm90sln74Wa7mOiUARbdexZeXCbJQMfN
3/o0o9kO4EJBojECpxFy3aFxFVKCGYmCsQSwRsuj09eTds3BYFbk0yZE92k20BNrUqiVSgs7aMrf
o06KRZCs5BXyyr1eGWgBc0oZoyUAYlO3u5rx8d/DWqf7qMG70u2/5Hb5/oNnrxOIRyg30KHzvgnd
30fiJVZ+UaWDSFbkXack8p8CHMQUJjbDoT8UGV8mKb/3sDHaAy4F50rVGNK3+eEArTi6U2tD3Kis
bF1NGgNe0VU5sJRcr6YPkAS+WyGsEjhp/LMoRY0lV0pV5XNdeF6Mft4WydlE3Jukf3/FjLautQT2
TEn20a8cNYQAWPKytuMbpGZWkaHoalPpS7Z1gv+S7rGp/Bfn29w8XE/9OrEwrIVt87fMks/eZRSN
uBuCYbbMEiF6CJ5AZhkCY/cGmU/ICCTbk0TUsSIxnfGQ7iObpRGPeExcJzY7EVkP0cs7qE6NzSus
btXEl+t1dWC9hYMjIYD+TIA+lIReUbdG7f4a3WqlfrrXAwWtthv2s7bKN22OCgXiCnvraakMBERf
dxufLG0RrX+KZRN1wGuslvswfxHWsAln/HkoGmIqrwOWwQsDvZMOVWEUKUaBalKzcoAozA1pTYT+
LDzoaEpwDn2Bh/ZI6lqexJLXyoL+HAYsRflkdJo9YZTFhS5bR4dFyl1SAcFT4ABSc6kq8FnNoqfs
c/JORPOWVjGXiMxugG+X8q9/99L64ayWSKtBXpbci6L/0xxoZSIAuGiR0S8XNDfewwf9CwZFGBf7
okgE1tInXvzpFbRHfZsuMtltmm5haRgg+c8cTAdtpcqBED9fcZVioUkSvb3wL4iJ9xJ6eXWIa+wD
CdYC0szG+xKFtHX2ZWjmDGM+MP/RnNb89Y3585PUi6moiNxGPIRA8MwIEzflGgiW+UENiXWdrjxT
aE8yHEqlKtHTIbCfL0Qggqv/QeATk2D0hjVy3BuDnrwVsRTpcThImYBBqq4dTFNkpewJTuDKnd0U
DF+/gtVxT1LnvoICk1v6g3YBQlSly6LoZyvWP8rr5a/bXAl0WWyEbnWTHNRDJBvEqWNBKalDs04R
yHBhsm8HBR39l25Jyg19jnW7BgEPIklsKhwUh06RkSSIf1ssP6DykEsr6+JLfh5KVstXAKcP45T0
OaJEjHnfHWdDOqakck/T2iYPqxcCpa8ECeyfTR8mefTBGXyKNWmEJEsDAFjCP1REnqaWHIpxP1qF
HmnxW8JMOyjXg3+8tVJKWKUUxqCK1xsHoRL4Cfj5BGKhMM0LRYn6WqRElAQXuMI/QRjt7vGDhICm
lBU4AYOltyMfeY+ir7O6eaP3gFfXmiDuKyHtuGpIXwEZIcvDoqjvMfdZNiq10jfgfs28m2w+cYnJ
7DoL96qHZ0ksUOoCKFwMIQufUqjWKourCfWqvjruf3uRj1UZXDVWzXuHUN+aldb8zbDhijIPryQa
9TzWHYkI2LwDRBU7HZ3jWRHOQyi2lMvGvPiIDwblwdOUW1UxyGgvVo9JYOXjGxNI4zMF/GrlFY8L
q7H6A0cHwGdmUtTJa7lu47CmPK104UKupk0POA16PWfrB54kkwv+/pKmW9NyrQ9l6956Sw1A8Uwm
6O73um80kdQdWQXBUZUeVYFlp7JbOM21zm0gSSC++fYjJhDxTVTdw1/VwP/QQjv3Dh4VUOp8tn+O
TMUawx49oEsIvmflPzbOEtj5fvIvXqK9oUubQfxe3IYmPmlaauX029EIh+nTxBEcy9ye56qirkEP
6WNkB3qNS2w7Av8yiwvqbnbhjiCHo8kKS64+nfjLFLVdmv59CDHq9jYaintE3TuAvLc52bMuuXd1
n6Waj8BkEPNYYR3lZcsjIN8dkljy/pEO546pHFJYa0kcdJruy1OD8lkPnqIaya9tGTJX1g93aFd7
JUKf1l9FCGM8UFSUIHN49k030yJm0WMxogf5EHtAuH8QbnZichc05lHuR0PF5OYXasGw3Shxc/h7
lvKRzHf3lUOeOAHKxJp/V0jsuaRUrFT/KA6AwNUie5V57/UXwzElXLrtb7svHuKR2RIl4M6BH9fk
ytSprsjn9k35bRIhK4/o7CsZoQ+Q+fxZwgm+Zz2EYtZcLA+JWuTcofe3GA5cVGlXs6OVWEiVkoH5
Ut3KXPP/CapIel+MjQwDQmTwbRatBAnz+C/lmIscSBZ2T+xVbIkSCCsEARX7/L7RsVNTlOhsRjHk
ubTUhX4KcZzucuja0x6H5L2OSZk+HgoWybzoGCsLuhiqvM5dyqUj4+cQxZDaBAus6sAyp/SjcnHz
bskTB3N6uYKV7T04QTe0XARONPNVkreqV/c02vPvkx3ZJh89AwC9mtwtfLhzAUDmsgFBl6Yj69wx
9k/f1GuGJjhwsWgex7Iwu7S4QlufgJwKAcH7+hUAjPIL55i1FPes6c79Oh3G2zxsYjkNqarNRaEO
2q2yyfZaw5eKD3j1KRUgM53/KNQN1q4nTu2SEg97lJtv64S9j5BHjoGPdo/D13ihaw4I+hsh0jVD
9vW02aOLQDrIsejchdfIY8yHCROItkrLnbRUL/JyWqJt7IgsBkiQRJ205ZI2K/RUPY0FBQD2uXcw
IIIJbvY82HKrDOJdqFp6gYkMy9sXyNNfdtIyZZQ0z0a0NkRoeSQYfsJc0h1MQKsQK3p7PfNREUVa
PFEcbDC7YqRDtXOJrYMOJoAJh3UimMwcZshR2vSP41jRYPUQu9rTIN4HBcaWa7Wl1IBT+2YUNTlT
Z6U/qt1GrVpZFIlHz3zH4w5MHurU+YkClOJEzoa9ZMfgs585+wYylAcj8/gEvxPPWOotPh+xKuQx
l0AEVyqW5uXW9Zm855RZ4fFusqduFVzV5sL1MgSdwlQ1g1AeFn0vVyVTCA5X1B77j5ree2vcLjaz
NSInvJN67GOjn8AhHBGhko1QMrIFTqkniPPe7kcbosupgKvT1bl6baznQBgbWFNSHlO6q9FbEWuG
PYQwt2DCpk790LRJUPKXeaszWW9haC3DeAee+na9JORXqpsyL2dzitpp9wtJHdLmsIVLRfyRRLeJ
MLkfOO/yJB3Wm5W6szNIKA2/bqn2d8ZoIQfm8scGcK8YkQwx8iQPithUJr7CLEPRH/ucyX/wkL0Z
EOmrob/jy4mDXNFcXj4r34B4pWrGbf+MHpFhdqzW+iei4HMusPWlC4PE2urAXjQWTwKTZQdt0wbt
WTwCdMr9qM/jHu5zbZXL6lLxaXV+fAwdb5GbhCCxipN7/Twx1yARRG4IQrh1o8KRWEWaPrgDge64
0WNg07t50BU7xqUqDpXNAMcpgv+0phlFWLbPKxz+c8vCxj0YjZZZuaLQRS+XNkeeKY51itUY0foM
855Lw0wf0o20u8Ky+eZJ8h7INsXJzMbcJP4D6P5xwQ5vqvgde4gqZzs48U0Fd38eKDYkImpcmAuh
oHJt1ydNElz7esTOCv1n37YGjgyCwMIslSONzQxnzarRYt9xMorHWAwjXrHhlNeCgyRsh9e+Dxc6
22q7TG935Btx8eAv1WfN/cmKOq9igZ2kjLj3y1LrRjJ0F9sdodz+Qvzio8VEaQ3x8IrL4U5/vL3A
s4hjAio6IB+13LIIv6Ea/P4B7zsgPtljFW25ddYtLQiJ76XQmPOyzQs30bwgZ0lZ2I00NJLea+f/
k/6r4bajP/0ONQzSfIMxVN+9rRMHJFQ/vqEo00VqcvXGaYpZboYPAo0nTJ5gy/NwUjw4ywcCD2FG
OtwDmZrYuSOnvg2ihNJ9fjHO5XNGAtMlYJJJme9FTTS80sppIwSbR4bWddoJ0hPSvMlH/WuruNKO
Xxz6fqws2Wwca4Cw2TiD1DHD5Xzj1Tnmpht0iPFz8XN4mLB9ZLICd1AMrK4e1bm4uX3/TgoRQojQ
gBAz/cY+oo3+0L/ECnoOySChowuE8yN8p+SpGDmUhWhswcYrUilVvjcy65bMQT8osKlbXFKYpYSf
8lggbD8uf5DgyGUBpJxb4AMR6P6Qb1v1tIVZQ3yzGh3mMK7v3EOC8cTyW9PN4KcHjOShg/4gNvF/
G0pMBv9mm8LJG12uQGp9vuyF/k7XrQZ6H9h+QZzRvY8NmRTYy+4YlrQGyIBvKtT5IhDqFEcTUpjs
oAfWonJ6i+90BmygL8JnQ4Ij4ajTLNHwhUGNBR+pOFBFq2isudlIfcjo/r8EW7504JY9xNKnvYbb
DMowVTM6PFX/VqGtV7YdLC5JYkmKjYSjwyZCWURP3pGgBpyWE6Jwcqzmhn+WVqIAMhFbEXv6wqsl
VWxx3FzxkHn7QfJ09A6XkqlslEOydHoGmkE3H2KW1vxbxyuaRdPv0yIkN4sJduGhQsg2DjvdFi0U
4G304VYIT0gV18O59uqC07+I/+BFc0vUhzqh51sZ16MjS0nh6OUVumNHygFCaGvvnhQW3nGxC5Ng
ZNupOJFzf3W4+VzuC56ltGtGdf13GKHhCXSubXVpcXFcwQkpi5MhS8RGOZ+bWQtXK27wJnF0m2T6
zj6FLqgRyLcQAVNW8fpe+rON0GjfMpV8fnxE8CVtc/P6GaaXL3fLXBrJJ7CXMjpG8faV+doTHz/x
Y0JPdUsHSH3MbQJskIL8vQWpA0yscgD89k1wbG63EOKCuhjq0FN6xTEam1/kHbvQN0gWZA2xY5/q
MnWTQbSpNwO54W+ComRQF8zzlhNRP0ewzcp5eUBxefRL1WnPJugAo4fOe/fH2im5vqC9j8tz3MYe
TgeJuNvmhYzLMOqgjaUoG/kt39LZxyd9GrI30v/Ny3nacUGyoOEqmrJgzqce44BJxnUwJJQi/En9
gwTosiK/yxp6H65lm8E1RifeUGZmp3oTdAJOH1CelzW+zUVgm1frWfzHlZM06vWKtBnpbaKBkeH+
EMyApBVs
`pragma protect end_protected
