// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:35:36 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
c8nxaNAwAYA1GZ0+d/NsJZntKUPHKKh32a3PgCY0O+S2trUk4Sa0pM6ssI/1aPXh
kRtV7vH//+NTcgpfjj3ab7h5fWGtFwex9+d/aUxQcVf7b03Xe2GEqCGV+N0ksH8L
YdXxp0A+x9EbCxfBDzF/nH+4dGaruoz9hL6M5AAmTzk=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 7344)
s6TRKEBKp1OwZb2yyheUBh0I0QrIwI9OLL0PkH0RGeGDf4ZxDEqm8PNGhPU65tFb
cSZDtFrgo0AnWl8NCHQuFGXoQUbbd3y3n1RRpgRicbL3Fahxrm3ZWyE3uEny4j2M
+BZy58+vLO0Xi3Iyff51iPb0eAw2F1KNmNc0t91RnmsvRKG3KxnHMdPYQPWyOrAs
KRFzgGwntVYjwa36epkbHIw+ljmf1FktYuKy2Fj5xXTy4ry5O0utrYST83mEzADD
ddMuZFtoZknG8bQyFk/y1LRiO8OW6sCFW4Kt+Y5woy1z2HInjRcKRqkSplecVbM/
/O3oj1hHfhzqoF3yXaclYacTny+ZHjDH7+HsW7FnZQsZYkZMMjfRUoxsvpqS+Fl3
tkFf8rpUxPGzSvOcll+JoT1zp7AQilTWImO007Z/Ln81j4Y0jvk6ujLxd1aB5QaE
y+Eioh2RFaWMwxy+zN7CJ4OW0+lX9QHD8iLMpoA8g0qWWdBCEPrOBwKHX4qjajtA
9Q/SPA5vrgDinRzkfQSgivwIACF6Ncj4aQ9oa8EWSuFsDFxHJbLSE7CdkXpUNmkP
CwV+G08MY8aJdVQW+fEwJGXB3to3cta5aiRLpdFOKGVfAecjo5qEE5hloGHJQN3w
1oLlCME45j5YGV+NJ4SpuVPOYQI/b/kVjUHrFtw6vP5tuYuBTCl94qi+bc5BS5xG
m12IySU5ED4a9jwIdi+X0IMrXzFZmsgvTICEUhFLdhS4jXN1JAiHDTGYBcPCaNrt
58xpOB0efzKhPgVsZOBRqcOmreLU8hMv4Jnh1pZ1+1G53kaOQh3GuqtUOk3RTNI5
0TMljcv8GnQvOUmYafthfF0vS7GhIDqosVM9HH2lNOcTO94zU9WP/P5MXP0lBlR8
kr34AFg7Ia0jDw6UpyL2Kw6SMt11eqPjbEHoYlpro7lpWxGNKhj2Vp6JyBYl3Aeu
773x9hnd7w+ROoJpRMRLk547xSlL2s6QwVPhCo4w5HzfHER9tvEqT+lfG8rd2BSn
EM+0Ibmu7jip8AjW4TVlzfj1Ovxz7OfVt8fUdIo/sPIqSPt9WB9vrGaCR1NgeC36
6WUGMf3jnz1fxkcSYUjNVx8F8yNW7b9JiimdYTXHBK+P6TF5WPPm1zGutrCwGNkM
QW8Qf0OOwoOOVO7PZmmbVbw/9Y1NAbS5raVOWDLVgpco5htWmiE2IEvNJBBSULxU
hmfdAMQ1l+ZphGSrnqzcsbc7nmg//HfvyJXC/HLl3+uF+5pcbgkchwXStExYL3Af
VANUjvlWRMLL03S0hB27OiFYYHrSgF0VPMgl1KPJ8xnzfXFD9q2hq2E+ptWR3CqT
KoskL8cHuQCe6lMDNU1kyTdChAv9pkmbG9AfHwqLHr2hAQDEUFUULD7oooLr7qAi
UiGgaSaqv9WojDQdYNtSHyYsAz7FREeN1Gp2XkQYphWaLMQ8bvAvyNVXF8eyJXWA
kyKU6NfKMB64/JCdPdRkaM1vNAkOfXfSncrPrcNZpKi1v44xxsuQC//KybNymn40
wbPKn5BIGb1uKGD/nrFCG3Nx+vK+Hb2b2dPlU93FE7zHcDzUugXqvwVPZZCnevgI
/H09Fo+Wn5sohRm0zZL0nrgCkS7UqAAfVlFjG7vkLGH+QT+dgXAHPKXGV1voyRf5
azmAK+TF4Ger3572K5dHsVlAfnO8T301blOaYQp1CWE0wyV6pjx0+ZOVFw0SvTLs
yRzxi72W4kJxe5cHnkwM//acTNGn6b78DAyuHixZuo3Sc2oO34SxZd3JyoF1/02w
q09G22lq7p1CzUlHxspMMEia9WIaCkLnQyTKw6TJ5Z+oDpSQ6GW+Qgp4QfqXMIen
dQrS7gkSGtI268w6ncx2Q4CU404Ek1I5w6LHxYftwdQYddNcnNyM3wQIMSYDBwwt
oJQBZsbxGp2KPwBTUq9hwDN/AZdf0mQU19IoLxkntWc9hSJb8EfcgtDdW6liqtyk
w7rZoVZDtIswXu9Dz99qimi1ZCpiLGP5UVv0WjMgaogF7Fq3EumK1GifBOgSkrJ+
+418GiCDukNgsh1lnH2y2HfeD5Dk6fOTe+fPzkL9Irrj7QuR4vx2Q/6NBFahzfVh
W6F4Rjw/dQPJqcmxjXBPMbqh6pKrPKjH2pmHPYXeYhi5ImcDbb5/kD2q/F6r+Cdl
qSUI5QVfSUHaiVs7durbj4UFY7SZWJQqiqQVQSbl4eE+QXdWiHVLLCWF0PbodcpJ
DK2I8C+86aMsAGpR74N1GGo6HGfCx3eFRbM1k6aRIqbm0y6Wg+d8qs280TwQtBNP
15Q68Hdh262kqYInY63TfYpM3noNEzlP49zw6EiafhQEYGkyDTK1jlPbujZ2K87X
bMgqkxXj7do6cxo8rMclOAFDCGVhKLjrGXI+qSLpuC4P9moJZc3dY6n8csDlEN4r
rFxJAVa6j/ZoH6+006XEazikViv0jAVD/3fwJsvymD4HVvjaB+U7QO8U2m7zaPo6
0A2AabZ0CJGqcHrQ6cdNbc9rCGjj4+pj/EXYdqdNpOz7gMQfz4rh3hygfW76eeoW
K3JyKE3ylzJsE2gltan70ahxqdMKSju9sYNRG20nlsqc22rlpBqCCzEmpz9ldo46
dheVSqiSa16dTQNwkIBIv5WbfVCzxKEFsvrcJ8E5epYcCiZ+SYIDN5D+xaMTVG5r
D9E+PRPOzrt4rXTV/QM33kzd8u74TPpuhEwKLEz3ASu0C1dNhxpdjwXQpLxRZJrZ
UybEGBFWFaR4I+nA1jLN2izmUG1P0G2fPK/5dTvEGEguXmvn4ZeuAddfTAwQs5AF
8LzyLE+3JaKvDl2cX/sjM652pB1ZHdyMOjQAWS6vVlw/qKMsUVAQQ0rh1jKj7evg
hb9nlqncWj7HRoQA/frMk425I22cXWE0ZtOpFAPzuBJBXpS4ujH/EQpEhu3DbTXo
PYv7WoLAeR3GHb3rFN6JWPRH58LMs9Ak+x1pKe/Jhbyt38TZ6xr1fatY4JD7u+P1
2d17qBMNGNRSlFgqnxNTBUO32t75bPKSu/uU4D9LTA2/Gfq6MMzh5yAFPB4vuTAX
OPcbe36HD+Xc0c8yoQ1PdWXxi4AH5SONIcP+iV60WS5VPusrol+OA8p/dLOOPBUs
Ier1BLtHV2rDzhdwTxa0NJhyPUlQohIc5zvdngAYy9q6hP2BJ5BW/I5S8ek8PZkM
NPQL5bCABVO0xrrUrf5bbYtUZ9JXI8rJO+cOuy2PnoIRYBzND1OUL9D9q4BxpDGa
KXTyfX7I4t4RypNKM5LnxRt0iS2njPXMTW89LIMMrfDRW5YTZdxXR8leBDLfS2LV
hq4CuF3nRt535rheF8F49ngQpyPdP0Xp/9XD0QiRxX+bgOqyAiNpOENCJA8hyDUQ
j1tRwZtjbj/aIEv9Ezd4wcHFv8i/SmpKP1dYpeb8TLwXt6+Zj1aGA7GuWim8zTrZ
7wUDUWRWe/WQsSxxM4yob9N8VOKrzWqjPcDLuXYG+Usr9HRYKkF7CT7f0VxLogcI
RXjU9l20vddO1ZMeT8/+658Ov5FTEGRR/YqPwNfnQfJQnyboPrV9UD5aSutr1nBq
yHHnlKkAQnuxnVNpNN70sAj/ZEZWcUhrihHG3oK3o5Ef2lKk9PGHfLdyXKV2jNfF
4P0weY1EKa8BP48WooW8hrzyDHHOd6RqUxvGtDqC9y7pWw+8c23i+2TTSUoBLdtg
ckGjk437ldpYF9WZe6cLaTpjoW8aQCxgrJJrRVxmip2f0o/wKKnc/v1dXovO3uME
Tu5IM/+6PfhB7F0tSCHSvxO2HXfw1Snxm2/NVzEAMoMAGNT56rWEHBKizp1Zah6v
3WXjRMgnuVvxSLzA5VKswrESstua1BGtWjrx1G8W09KlO8FIxw1nh0D70wp/hJqH
B2bopvYADJv1VYiv2QYelYt0ww0OFWGmlPiRvEoTVuBjynpNVz5YnJN6RO8afc5e
5EXB1lU2QUrpwthUUy1mBRQVrZTnxcHmzSYA9OK+zISX6Jj1FBUYr6gMbTi3naYP
n3yPQXUDXX+Z1xNyLUNJwZyToX7//CUJMXXxufhsD9fOincui6IhXwR7lH9zZkgO
wSi0J7dHNU7/yEulLffrJlQSGw69+spupD5/RtRd0LQnhJa/6TMZH+XjPGPGSLPe
H2iNAHYhblg7ZBpI7qRNninDqfFDboGD0WgactgpzjPS8Sie8Cpj8bhlqGcQ6zcd
FxKFh+hhOOfgiygC6h6C5gAo4mjUi2QXxtiUImAtoYFY7/R4OWMWWKZZKyXLsXyg
4qUEB04oz5YjXHv9hJ0WlyfTwXmXjdrGK7WyVQONJuruJmwRCraLd53Ll7YtZYt4
JZjMQD38avtvwi8izOwrMW2UVeGpOML4xQGlodVOHNQe6phSWLnJdg885AdJryTF
nb2Njq+3TAy/YtmHtvVOCYXDuNe0uiUtK4MwG8ScD207L4mKrl+YsLT+ztVMV8jE
KqTuyAj5PLmuFFl/r8yoHElJOteHCdPBSTElG0JLOz7XxDCEdiWgFW1aGKbwLcT5
IzEJ24wgPA5f0Fn2lWcRRawtoWs2i0HkgqRL+9Y2T0TXCYhu0E/m89/ZNsx5aefI
Bw9q9sceUEFi7nw2lImyxDSFQUfWjqNcjaQwAZngbH4GUSicHTDNE+6Dh85X8Uud
u+A14tth/gjsZztFF7r+quMy5D1TjdGgtMsT3AQRZF+5JSfCsZZ8AdTa7XZI1ryG
nnCupOg70JijAm7MMyMXQfDBI1dIb68yzem/4EXPla55JXEHFw+3k2Qa0IkSdT6k
BsF1mXnXyowgMtvQmWxKYfANkRuy/1+oNUZ3t/ZhETFJn5Tim9KffP2NJ8Ubm79r
tamEgIL2uCM0yczgcXRxmP/L3qmrm7UhaESsuF8jebc/+I+gpCIc4cSQr9uwPIDV
JCisxGJtzt1oANRV1t5vQb2YsnUjCqKnDx4vyWbErtxp8PuWM3ud42PV60vUm9Vp
PMSvPygDbZlQyTIEhe8lly+PH2kBqRGGr8xJwC/NmLpQuMmmulbqUT81AW/UEaKA
lQkEbqRMEaG6njuTCuxYZaX1xOif138R18zLcME//ahNIUw9kDAerxH09QJAopNX
/6CCAskoQ9kEYtiTylL/EASa9kJQCMrFkeygNAJJwypm2/HkQqs1eJv0Wnpcuay1
SQSbuimPPl5xyYW1njGIaw++8UNMda7scw/6/uvsE9HPIWYx81ftnoN9E5XsLxd9
GRT8cdEJb+fNJPmAwiDgWvA4TWNarLUMqL0FBO2fQBD0lcCKtrNwy+9i8j2LkTM2
LufngD1DUzmWy3rPa0ob6WIbw65rFohbTwUd+jJGo1IiuZa4FkKrSyMyCpgJyGFy
3tN+YsBkbGzIU/Iz1lzW0XR8fDwOd1KbEzX00yQzaBLqlHozIFca0qzg2I6L0RCn
HDthw6kVEtcU0VKIT8gKRo5xD8Leknt8QVSu/StFzxQuWkWo6mzMn8gWtSElxysk
cFKNjuP69xIht1cbAYHcXi8RrQb8eQaOwrwhOaOJy5r0IOKW0uhKaD9IzvOrr1E1
ec9CvVzHNaUDzb7kZDtli1hs0lvCN11ZmRZYWrMnQ75sekIGgrkElg3uNl2eqkuu
g3tGwYlvU6ar3Rfm7oB1sOIRHJYN3cW49sWFGELhzgPIdjHk+kRM+iTGca2Qx0GC
Jz8HTwwFbYoM9wLCJCK65gXpMfl4ETCSJMWyCzslEiVuEEnIpvrl40F7u56nlKnx
paVPxRiYiGmPzIZ8lCf8ksaaBiHC8gu8OJ3kO8jrnooOisJCMb1Tb4kXqRpxM4gr
zSOWXgfSNLbeiHhA0CCu2UcXmAweR2xjHH1ew4dLsmD2eMlx3myl3DAfTlJfvgUw
cYcln7xBPyvVAHGjIzRS5j5csk5/1bcE5e1WDw3W+Wkbp6TOZev/T+woGv2/Ct4N
OVALNe4pgMKgbV1hTZUoITklAXaFuXQahvWzVYcZcrlgtnb6dt16YptZFn/8fwTU
j9bRFdS1GwsMF8aJiUcADaX53iShKOvpXT/1DOH0feaTe4d1wFRVxvuOSUIlfyA+
zCjNvuIsA+kKgYH96K60KrqA3ZD7xmUCMP11ZjyOUNdDYOExqZ1ZsQ0YFo6+iW2o
rSEOmCk43TJIn/myREZ4nPRULWCuHZOhaEW2qhxs+USpessSra43mEI572gUJlHV
FZz7RjKnP/W8W5/HJOvs/6P4vWGHJOmLAf8msClM7fKWSPWaBGdUdgAKYUHOS5XQ
onnsbCpjxVlOMh8zS2nBdrRQfoAnyKjcbMuTGGxe6oDbWiSCOjWlpryowVMCXBGG
X0W6cERP3su1eD4lFhjARWSCfjn+MI2vJHKnIVER3ao1g7MPLdh52T+H+uA/brtG
5FmvR1K8iQ7y7e8s54DEd52zBfxyDq4guD1zKaRlpTlOrmXqb8ioia0OWlBHtetJ
vkXUlAq4wl58n/J69dv6VU+XOzhu8g0KofYBCUAezKbckv2QYI70/u/HlAtJGx3F
+/jHhYC7ThZ4rcmssEi2pYcPdH0i+YDqCZNKfycDesvG8PiLeLbKRRCc92sDrxXf
+K/gyCX4qQVcLQQ+Bge+1l1fD0GLPK12bgNEa3oKpakF9BqxDfMhNaeijRRxCQnW
T+Yrciyg6aQv+t8bbD0U858KHif7zDLP4C+3wRjYELRvNqV2cIanD6FtMgK9ybdF
zjQZRWCGzlF7WdUtnW95Sx3vYvSIyCJyIwdR8hZrtFNUO27Jod3dnSJX6SbdPKO/
d/xOdJHe+9R+I47vxywVZ2obNqoSnHt/5bJeOC3+aAsPuntMp/xYuwyGZ49QVvw/
VukKl1TfOAsVN1umIKHEMQ9kn3PpbNNP7GccGez0Byb8a4i8R6fBspTET/qOEKTV
nsl00VS0voFI+jQu9IwwKI9gbC0VgzCt78Neiq5UFsRYrQk7F3bTB5CVQHQLTP3h
ITAfgwIFhmFY3qxqZJdd/XICwjF/nL8TE0kpHBHYmhJkT/XKlhENwzAQvX3OW+rC
evssXPxcnBQPtkDiL9Hz7ASyiPlyJm/DTvCcTsT4/x6p8NfCZuWGK3yjkJ9S3ntx
UxNN/rPKc0JHTkpIbbtaSMPy6uaSBB/Ozk6/OeFY4coN4I42bgff39wqiuOj+3tW
xdTNbC6Od/b+BZ2i2nK1+GIIevQbAXC9ElBOk1S/aWPq4q32BnjRXAbKl4TB+4pO
zkdMNmMO0vJlLLPhKiKfeXZNfDz9PxZcTzPAzfvGIFhJyiFRZxxrJ0smjT1GzUwq
q5YzCzsi3kl6JfQB513nYU+om8i98XwDw66jyg1DRgx6k6Cx3AcDzuzVtWIC0UYb
Cf3yO2wX8iIwHmMbMTiFaigvrAp3WmakZBq/Fwt9JAQ//f/vP9ZHldy+Ijvk+dW4
9wBImvBRH2ZyMWq80mxKmUdfwU/O9Gv/VWRyAa12WMtwI57/VJ1R1SpPkBfIo8nk
RkPMJoKNQuLQQpE1Ui9a6ZXJxsHto/AtwyQeLLfWOd7xU9UT2la7uV+WvR4gZXWD
qp94ptCnwp4BSsWjDe4I8QmFSeV96eQ+FQzMHUDAMsfdQ18yiiEEdcv0d0VK0dP7
zHgeoteydE95lJPqr/eLQ6R8QO0/t31XP21Vazxw/fKQXjHM06TmYbW47hCrzVgz
ZsDlX5ik4H0pu2EWu+EWcOeqJXftIAgTvlNM2Q5lldZk8x8bwqpwqquvTfKeHoHA
WFE5m4AK1RmuYLRUCj7BawberGjENYBqKcpt+WchrTl8tMOAYyrx6fS4KwAfVSP4
1WhbWxUtvLgIcFSnlbo6PD2BHrjQqJ5WUyZ0OJ93JuoSfy8SCr772YWTzYvbkefE
TMD6iFXkMgbLOFZfj2q7odm+dBaxoYnCxrNtWCMeM7g620Xayuogp2MTLH+PEgJC
Og8yLYFkavbHhBzvJ5FDlw0mBhnuFbhjVi5AUdC7NJXqnnVmhiAjQqa/gxVP+FAV
PrlAe0nuEyL8vuBArJXV79y4FVJCVMwhtnh8wUZyHetp682Hd2KQWxbB7STQ+hYW
aB+zD3s6X6Lil5nZcTvD9Sav5fkiub2dH28aCXjP0imH4F9DYhUgCM2+CrCt7EVW
Wq8v2GqIbIS9ZQ2tlV7R/0A5dcqA6rPPSTghoY/+SBISUa+NAPaMet/TMwaFO2TP
jODDdjrdCywMbkx5uReGdYlkfl8iMuRmwdQ2pzS+wuGE6Zi9/pB4EnspbbJ292tL
ix/f+N/dD4tzpw1BMz5TVRYR6hLGaEYbw3S23o2Ji3ISZGtMKSeblYFtB9GOThj0
JIcWpbGCRqg3vH7pE1jubRkTqZzK9e2jYdyXYvram0/otTqmU7kBRXwtdejVde0O
x8EI6ZtR6C6DjwI0wav44MW0kDpWM8hopmdai9bUQCPdsQU5ItjMrscs3IzHBwGT
h5wViIHVxkrF6J3hm145kJmIXmuYZs9sTrH7qkKD+6hGqqKgAkUBE5a2HEQHoZ++
QavNO9Fqzn9JFbL4cTi88Sc8FpaJBjcivX95pV5eRRAskawjv+M12XMOGPoO2Gzi
WLrtdAGK7oQYmnu322Mijzi2WV4m9mvn/nYntvTABJXBGwToZ4CzkRAbqFxXoNoT
nBCALq/Lc1ZTiTJFetG64nVkeleRQc4YlZqdE2IPmfPnGgqSuQR/pugUNov8ZAsu
9z1Xth+tvx1OZh83J23oCsFiJxnTptEPe8EWFNC5ILF891hDJVX0AeBrK2Swr1oS
EAOno9QAe8A3J8Md7FmB+F2dQzj184/Nfj100W7MDF3kR2E2pGEzy7+8ooDg4QUT
OLexxo5X2wGo1xDCiAZfciSqGoje4sPFkDq/mTwY5KeBPhDelR+B//U/SUOW2sX6
J6DH18FOPpXstN5JoouSntftbSJQKhZPbazxtzTtIUnFBM+4T/6yryW5ybBKQgNT
sqX3FX0SUT0XZDVmbhA7wKAnq6KB3guo2u1CIJ4Ii/MaCDPF2X2P7Vy1BfM2ojj1
908jWvX6JmF9xG9AaezqvhGMUNkmg5eS0nVz1k65Nf2Zo+UkfV5cm8d60xmePUPw
IVuOcHnyQNJhPg8ZAAp6nZkj6/SQXCBMnqs9NxtWczQUCX986esiVKu9sP1dTkWF
a7/0PjMCqc1QX+B0ubh08VUGUk2yDQk6SP2Vd6XDn3qw5NxOM4Ez+S0RSUiaaBtJ
JfC9jSegPooXAs9uEnuahLzzAnuKODlRz/42L7ukcHFTDxngKV3qSH30Om+5uvYD
ArgtOpKdUZtrf3bI5Pmssf50L40n9xO0/pwyoomAAczhL03KTgeShWd+Uu2lsPzF
cwdmFExYBxNlvGTTLskS9AHAPIYhQ4ikUXNZR/neRBw7Reu+oHewWHeInobnW8rF
975tcsveWZgN/+FQuH3EhSuE4ndw1MKkcCezVmmKIpcP07jf38JTCrx/2+P92VIw
SvpdTTu5BpuewSzkYt7Z9GCnMsnnnIYEEIw6ZjVESnajLT5vxvrVViZCk9cVd99I
1Lb7Wn7z1aQud9pSOmy2KmOg/3ADNjeHDDdXmApHOt50+WvU3K4kOl3o47AUo3k7
cSfI7H3mYAqhG3iHIZZghIqj8qFu2QjKc06P2VRIVDB3hky7c/T818v+uNl2sjxQ
PA9FCJZFuEShqdB1skxQthpDglDVDhjc2KWPgqiBBARn+AgA0uIkZxu9B/92OCRt
++JmrjKErzOTI1gv6XrNQF6/y/zfby/tjEX6XBhCLAbfLWk1yi6MD97QrKqyqrgX
`pragma protect end_protected
