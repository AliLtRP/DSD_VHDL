// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:35:38 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
FpQcgJK4d9haTbM8i0+m2TfGFyaYXCqTfEkIkGpt5UMl+WYidJiyvgSmSmTgTOim
HrdZvSt0qqouzNI0BGDIIvOCS3jkw3ZA/CWEtUl06TTXNMeH7XN0FLrlMVz2pGf8
cvUO51U9w9n/LYojwzq6VjsPGaxTJCzyk79qasnE6rc=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 11056)
Kaj/GwOg4CFGXkgtxFOfZnCycxamPeGh55cWYk7QErN9+f755QyogCK/fPDJcSlW
1QPSnpDCa379+RU1smNq7kI08fxOPO8Ig3V5VTxADIMWY41DtpuUH7WJxh9JZtki
M2Ig/XTEvHXQF/aCQBkhM755Iu1Jrr2DHEKQG5+zMIdgiQqbuJ8t3ARA3LrlKBlE
+a6j5Q/0nJxY7+3V14HLgb4DJrbW+16fbj0DTyInVuVjbXg/KNFP7sb4kBZCnpq1
gwezu9IVXHdomzHqWbJEuEBwRlBRkkNHkdP+IHds39CNqKVOE8Z9BLDi1m8ZWj2L
Ym9uxQMYE9MAjtnRSPhPB1mJMRizjYBab/jaM/t7m0Nw11pMxeShaTpLG4K1oBs6
FmqskFUJpWEISP3GmLQBtOF94hFqRpnIH31DJdW9a1dX+O6gFm/Gnelr2R572GoB
Z0OJKaUT5WsKsCpaLFayUR0EUYKoiGYdp8ONpiyxSX8xVoIEXoq+q7SPjsUGZSSk
LhM+Uvtrf+HjPxjXMJ2jd1v1DS2upnCXj6fbdTxzmnn1Rc+hqpfrNgHFJA65Vpfj
TE+2JM1MP8gLJTe7jIgOG3xDzV+w5+eqBDi8rqmddneSkI4sE7B9hNyQRb9ErQhb
0zxUDkXggXRsuVhCduqENEUP5+orncCTcf2Jk5Qtdj3Wn+xVX0IEOjYqOr8poOmf
7oyEdqOBF6YYC0f4YQa4gfc+V8jVZ1wwV+LyGm/roRRmhml+GkEClZBsdg9eaGRe
RMevL0kJ0XXtjFX3HPf4sqoprRMGTUTkg06tycwRLbs6A1R+wXrjbZADt/IwR/9N
6ZaqZHPd+mdgcxO8386B3I5TLkIf8Wgs0YrT+MsKDqB9t4O34Eju9tOhF1jJDGn8
xBNSX6yUcbfCcLvs7zFIn0TqZCP2j6cNh94LeSisi+jG4BtQkVVyxKUhBK6Zn8mU
oTlwcs8LqhbOkHEux8WJmeGvZ3giywu9KxIo9WRchXzcsAiQrNwcO+HxxXtzHKqW
kA1AYOt9IvQJkNafIVSmD5cV9o/pjhBZZB/nkHFaXykSlztR6SZxbzUVC6eL188U
MSLX47q0/RkxK5JkrZfiJusmllxId2CeUIrGqxsDssfuflOkgEM+WX94fa2/eyId
Evp09nqR/U85gXKzEo3+OTYEkHQbgBvI/FxgDWoGAaXBZlwXD0l8ZNmJtRpfElCH
rLpdffSuRsgJ+SYbx7RSgtaCSvGtd/BVR81bwhxQ5W1B6vWiuENJhwdekc+IC3LP
lLYAtxkxfNBIwF13rcdkKY9T0UcBFAY1hPGdiD1LWtQ0WjR3vzn9evPciqgUSVVL
XPBl7G7yViZflxaJc3V+wBE9YtClXlOlTDghE1s7/3a1qBkl8LdF7ew8nM71QqbG
+jn9dQV0BsCKx7xEeBiMPLTCM0yVhB9duWxJQ/vFQXLuzPn/KdfBmh80z5siIIYN
2SjxTm50OseNzghMoKKuX2484bexz/X2/8zjcYBgKUC61AwDBzRlopA5R+3gf3BJ
Km1tA7oOj5kxh9YZ6n7oDFzBE9H6xR6gHnZW2wpZnFUTqbi2y47LXcwWBp7+5OHT
f9lOXVWTuPCtTBbNZry7/83iW6Eob5GI1aVoBhnFVHk11k55E4//QyI/WFjUrElq
7s5Vb2d3gIfdlVjtVdxM2kJ2S5Rt9iXOE7Kn7oTCLOP/ZX4ldDKyKC0od6Z/SVly
FAPkpl82koPdGs8+HPS+8fzZ5NS6EFKONew3D5AGImi7xPOQ7wfa3PVmgyMtub0l
pWwX40jKblOYIGT1+8NaaV05HDRU8XuE8mofdXdFiDNEOAG7JmHyFCaiSYNWemmp
GT1B4VYVHw0cIo5Qe6kjbvt2hS3GFpEL4ewkJbv4vGbZv2PjBPa/G0efgbpmVXYM
MeK8AmR3NS3HbOcOzfm2k/1pV2drP8MsufLNGz9vF3FpsB7KOd/9INsSIBqlAhC0
llH4o0pf5K05Sa8JARgfPWdYqRvq7RvgnHeWsD5+pnEDIJ24BPeA4BjH9dhSzC0r
y7lw2OMYViibjX5p8fQdl0LcmqQmgUifJUzVJQtrdZ6E93zFg9Mui42Q3KB8jPtn
fR/beC+bTUOcRX/SuhLn3gtq3CTXd1Jh3h0spal2sO+nSMpkGW2GmNEhFpjptBxs
q1tJ+5a69D+mvAopsj94+M8bbIyIOm4TZ4/WXIjoQg3m5Nw1sYYlV+jLgmjZ+rAF
aGLVDqJs9ltMaeTIsY269SaghEpLhC6PVvl9yGxXUgOJRsFQJafuJ+Zgjfxwdzv8
jhZ7o7ppcRt0tGeJO3N3Vym9co3704IWG1maqfUHlunh+KyemrMvnC1FV3kG+aVh
Q1iccBISc2yTNCyG1aTue3ddJLmBFAz/9wjST3lZvvd/tgBGBulceuCR4LMHEbZj
lKB2O38dHXatgTJm6APuUxaFrW4Wyk5mACKyjLLA1rbxvaELj1/+k/YJnJEE6tFN
03DcyCOdJLtehLuDpFHja0wmfSbjojeZLDXjNK/2kS6l+54mUsf8/v9wXi9Cu24+
54UTn/j6MggpypdowLGmvQBOAuQ0jc0GwkIPJlsp6O2CQx6IIA69ovBbPQmFuBgO
LwxB4f2CZE8DRMbVWHWqkHFSI//XNjxBYK6ibXGD5+O6s0zSZJXyJGCIFKBPQgar
f0tmRWXNP4oFtPBNqMf8JKGoufAFDCZXxxz0pDtFLZFuG8mlS6rGgj2qad4ZNkvv
HDEXuWiyY1wEruK9tdLiIkPiqLilcAYdMluUkMEdQsK73SUVlfjWSVa6f8GgBHMP
0K5fkroUZ+G/d9AngKk3zHv33w8ZNP/BvCmgjsNX5AZ6K0TLTCDk+0eYaAoKZzZH
Ng2LT8eESEMUyu8ZMyltf4Fh8BJoHhh+Uq1e7txDuqzwZw0GDXkelH6VPmSmMHF/
Q0ZhDjZ24QeWFvr0krbXbOn2yXsap7v7CmP7I50CrfCLyB9axY8qJ9V2psuwvYyi
opQgDoWJwAnkEEIPMO1cdZCZRBwyckFIrrvYdbFuH5ebzD9laS9wNxcMzR08VI+6
P3Kq5/lKFkc2uCrDp18EcBldhJCg23dczEcFbDK/cKzpqiDSC7SoTAQ+yeTwNe6Q
OBrTbVfD3Xv0QDo2UqQ52B6Ev/8321X2mNWyx9JD+nX7LZiMTCUASW+15AGMvp9t
U3q49p0zqX9gcwXM2HsgJyP/Un2QVYPcb9r826l520jYnMZPvEXAjsSrk2TUYTs4
IsRj6j1S1wQJ/rkfHSMbXuWEoq8a7xqqMwdlXiKdkB6QYvri+XKXAYHk64cFqAlD
RX9yxv97ULId4zRh1ANWcSs3QW1VBxFGSNCITjgnG8CuzSHsZhe5hVqb7/iDNPvg
6kq82baZb9pqzwGcIcD2MVitUvgt87Xk4Ez4XByJHYc6gX3KqqGxwv8TTJMg4rQJ
qiA1qkSkJLSoDY+eMbw1N92CfGWSiyE3uraMsf8XV+WVYEJeSZbbuRVM73HCxTs2
lI75ouG12ZfBobu6TXTno9sj3Qf58BJdl0jVGP8oXDVHTSsEbPstVmpuA2iHtKk0
Kwm911OxyON69KmF7Uf5TedV+J4kQwYX+K9Kerly6HFTnVvQL07kg59uWVCLpB8b
RhuVHszz/deNgB3aROFDxXqyuyGpfZgVIXtfcKQC+fXs+jES1kL7qlzD0c/UtDWE
moKX0w0XoFZNQkFcT1My9dluiQGJzjBH3HWVvN7Iiw//NxBCzo4lpkGv+l9Jcdok
JgB1sWHnQGoYNq1Ti3AyNUoAw1AaPutrMqG245RPYXFAWIHyyMi9+k1lL/JAXmqT
8SYl1W34auLOzQbyRXRigTdz+1bL2deC7r+jkK/xp824OyGU3dTG402P/qcGwyd/
UlIGHYr+OEi46fP2ON0++orL3qB78pxTut2bKrMxcfA8nXBiIsWaKfLWANulmWit
cMf+VQeV+y2lIaJmchyPo8oFbgJ1aLq9V0NgEYKexCP3PTxDDFPJRojd6CQFJlvY
rdt4xNLY2JdBy275MoFwA2NCiLkWmbOSWWrU0R8vfC7i+BbZNf6WREvECiKzBoMG
MbD12Scq31ZhNBNJ9qhU6qwzQi7sNrmSSxxldQv48U/Y95wDMXH2Tf+XnnVz9a1H
/S1sVCTPUmIr04xyZeUIhkdYcQNrn8EcRPzlxh883t+ze1P6WTCU/o0m/OnZNZzC
lVwO6zXyMLB0LrRywaXBa3wRj37EtrL4bdrzYlGIehBvLd8H6l6L8dnqWENeT6Sr
l04lyY0DgXP2n1lLeYnLZu2e4WhB/el4GJkKMGcQePYQ1h/cjqnlp8qlaDtMQRUV
nUe7CEAIW/I99cSC9X7QCzYVmcx/6VkEZdNgyTd8RsmIU6qlSzjjqFfy/BDsv6IK
50aHiZ4YtWiwYQF/jaEUv9N3B4SOC77+fhu0Sxp7fvUXBv2PMuPCc4bIImknJib2
OTQYrfGCObLEb2AfyEWfhjPoLWPgrXpkGanAM9jm4RTpYy6yeNBDwTMAvMGPVUpX
YZt+G3FNe1lk5UZ/kARrf8AuxoPBo3evkRS3dnGSy1Ss9M8p0hFZG5V2YWfCTEIe
lua41Ix5UDz8Y2jY6eXA69I9vgTierUv0XVPME2oZeCF2OYidovXyx10Cc6oiNRM
y6PdcAlVLyfszl+ePQoKId8YZjD0CSu5o1bdILYy+llytFZX0zWUp3bUgeirB6ZT
aIp5oQxfVdjgihRzxjvwGc0AcbKktU2FzVUIRhepiM9/5Uzz8XPyEjczSmwCEjb8
p9b/KnfN3COaugq8Y1ImXtp+loMGo2kMtqSowBwflTLRvd3z2R3R7MA5+HvORJ6E
jITseIuVRGXw+sialL34rXk+Q3FHcThmdktteGvws69MYoYl+XEwCM4oQ84XUUyz
gYjhL05TFdm0JiYf+n1/i/jawD7M8UYpEnLJVzs8xd2FSMWdYMm0mkFM0N/OcD50
AX9patR+QEPV3iCbIXdgJ8zRsk69tg45AHOzSgLNCQzOgFXC/ldJCgO4g6DH9EQE
zUyzp5bngkPTZW3AEu1FOwR0Gu9VvMButZSudkm8nf/vd4VfeQ8m3INqWFlvSLht
zWYnRqmTlLdxMNqdOqhSclvt/u8fPKySfXs/HbQm6SU+O31t2SbD2QL7KqNBj6Z6
Sgi4UrrXlfMHYNtQVRToT7yyGzPaIX0ilYuKrwece+W+DRtgbVzGi1OKep+D8tHF
OiKO9C+w5rVYGZwi0IksiQmBD2SHcRcOJqAUApbA6dZKXRVWC3mkUWkQ4bQ9MIU7
w/ugAdQuPt+hJZd2uTuHgOakXxA7vB2ZFRNAzdsBV9u6LtP1Wi5Ykik8rCgxc6nO
0XhlXRIRf9MbBr59UxI7sWWf60XlPhGJMCjdNfTHVyKf15r68dJa75xWXoDEsum9
tMLVJ1K5fhg5O57F/uyug91WxaFVPHDndWLTiVgznzXwUyZfE/lGl+X5DkYKGqbP
OshiACe6Iw1lO1og63alOIrfS5RwBboCXzFRKMf7Jdea0vwf5REOeWiyQ2yXkDUi
mERFjw5zrkU2RCShgZd0HRg9NH31dxhXll1IJ0eYeHQmeY4otfP+T7cLlXm7PTrf
brij+78Q4IdShitonuSqk3G9S1PAwxOgP+TvX7znC9tVWINEH3yRs5Jkju/0QC3J
zrpSMRvLzUr67HxPdfeTl+D4tSKZDwv9PXw2vSSYSm8jD7SBzRsmds7CNLYDFiUu
M8o+MitPxSsZiViQGGuNrYFmqmifEYMixSjdwb4eFhVO6lgdpMcV8P3v1d6xCNX5
eMmOMIyy+7GW2v7F9WtCil8Dd1ZJnuNjl/gCEKp3Jqkl7dX1i5t3tKe3RBXeyVU7
vCyGcpsj7z3r8zS2dt5LN/ncTn+Q/8oZ0YaiXhuxc06zPD3OeXxhqCylVXIoRqkh
EyauM01dM9XUQQ7N7mPsvq2V3xccfBPTrvJ43KMBPzGJESE05VD7CxadsmcAL/vg
8IWw7kIehFauUMMhss127+azshKE3KHCaVoT+B1tcR+Nb9c/clEfJVm7gYPn/uqS
RxLHJf9m3oQAIMbDxikX8ijTl4QhPnY7yHM1SIlmoU67v1SPFwhKfQU1EyHASKGk
R/AyegAl+EoSOx+ohT0C4RHNGwx+oC/zPshCFMgHaA1heU4ojtsMuQf1BFNpxyFo
eGnSS4/sdOmPY1ndTPZumsRcMKNiHgdwIHm78ibl3UgN4UVYFvShtLTNJe8pzZdT
kRzo6a18Is21jRpeew+ibzRFyzhhIGfMRpIbVhGvdc5hAqM9lPQ8XjH8IzruYxSd
iLxubuR3HbNr4r0klpJUHP/ZtGhvt+GHUcgrxSdfo3AJC/B4Hp2gGWxdEXuz17CY
vhi3tXJ/jFMJ1YMiBs1By/Mtc8+yTf5A8ZWa+NANrqqYzUaTMG5DbCd5w0ULmTxa
ly9AEh21pybmMPFD6XKLg4iLLOdk+3TxR38tcE2+Cg3zzkv5J5ouUPPFBWffQ+Hd
864VMzs78Hn80hIomo37N1SWhutlKF9f8wlC7dj/V0tEUfvlsJs79fSjdzX395eG
pjd97P5uLtc49XVvddbnYA4u5qPANXdTNuCmDMMBRYflaoTr52wvsKOdT/d286p7
gQG/p4ty6OQcUed/k5vWcphdo4n+SSlTII68DHkdudC4y0Ufg+DaM8z1aqhUEDkr
UuLYqOxu0dn6I+IPZv1xJvpzHM9hO5hDUh2ivslScP64t9IGDEushviUxxO4L+3q
ChJJE40adrnk1kUAofyJysl7VmIwGpBoTx2coutvBw72ZQYlwhKjzkikHiLdkyMH
OFqSw5Vd7MOCXdAXDB361bTKrFMcWz7Kqa0l7n6qUTTX9YVVt0AU5T9gh7gD6AKV
jBQ4x10VBn1sIwmHo23RDEAI23oG17eGQ4N4mP0R5OOJDpm78UQOYNhYvUTk/ool
Ip6LG7Edzcesvug3mKkLj1/mM8XSCPCcqQLmVgfhLdVVrChx3UlC1QYB7mgGTL3C
++vo9d3SY4d5kdXqjsl4WzS5/AaInDk8iIuADiTZPIq+iqPPihv+xGSjKeeMHAHL
TP9nGl5FsHH/VzXNYPWFYw588Xm8b9wv6j1QkF7+6u2/1yJnFNOKmcBFF4fjHLAi
nn9iQJX2/DAmOjjsKgGQvP4A9aAIRgOIFWI+4triRO6Tcml3tDyASiumUduw8oM9
Z9d5HzifSx2BK4D7+51RDOrK3B5Zx2As/oMYv0v+h7I1iSuLtczQflMtrcAFLgiZ
G6/pEqZIu/TqH7k2ztQ9dUvaWyh+gJeEIK84aaF9RZbOQ6A1C2SIp0rEizWynObz
z+3iGBHgBDErHjnUvU/QC/e9OdZnA22Y8RJpbzoPkKOfNp43C8WxO4o69gGIevwa
b0OXpMtffc/cHwjutdeVdShqKwH36BvP1mA7AxM4L1C890POOMmfYJHgSaiCKPg+
9twmPXHgRd5KugZYmB4oMNJH3eq+uiFQIxfD3nld0dJReLwPIOZImNKp51g/cY3E
hp7i5OhiEDqN3REUT28oSWogVJFUcDFUSYfnr7Wxsf8bBqFjxcgDROmNFEzaxGnP
Ojr2s4MAzEa7SUjF55B8Z3rW/SHFvFsxPmVH14vjrM47pG2Mg/hg+guPE1eOw6B9
ntwG8Cp2hJIOVGIHBX+i3LdrrXLXLHw+2IgnlifByA+F7BQDQ8Fn/0A1Hva9bffA
h5JyMFUTeW32nPRvDk9pHjQVfW98lc8IQ0oFfTK8BdDwAn1BWMWGWNCJrmMFkmHw
YOw5dbDU0aSVvxWJzUNCaX3Gqc9rY36L+IwtPrLsP+7U3QX5myqQQQrGbf5IrAWs
SfqG87ZaGhV8PGEgliDHaEZlMxS/xPVMAj/pL34PBSsn42dM7iJ1C7MNvFk7mv6/
6P+vCT8JTeUZjTuUGFfGqfOxtfJGSqcoUBB3dZLNREMBWGsQSU3Bq0oFbi54Bkhl
kvx8MNf9vYLGYiIT/u0e9fxERLdp++AtCvgAy/trlqRkljD713FRh2xEuFrUutLK
kHA7/F5XXVAUIpPo3JHo+44Du7l6c5pMp4ONhx7UCgDpLr3d0MrJZeDngLt3UJUC
NQm/VO+ZhjZoBbeM/akQCTefTL9LKLf5orTVlx2VI65bCP2BoYgfAngA0LcQ37ib
35cMuBc1d0wAxEjEmtb+FgVO41Q5iGl0KfZY4MT20MHDDcvtu5/69t2lf1nzRwXC
JNexlVUocBIPQoxk6H674Gv7z4t1OkG2QHCSItuSr704QyeM99LVkcZxxXuRVT+3
EwsQ2to+vQbEpnXKroy+igrzcKw7OOiS7p+MDNBV5LNjJKUB5CBKnCDnN0IOJcMa
7Y9i/x24aQ/9+f1HvM8+jxaa9LRrazy5IG0zazUN4N2kVa81zbvxbCw/C38R4M1b
sxjLWSqTPtIGuHH44gP9IKn2oxlGaZtTlEnlDmEfco7+gO0bOdFV88NAL7wGp5BA
qVb6OiGimlM3cbHWc9V/xB2Gg67VJ+bslB2t0JhfFQjnVy6P3Lq/3FaB6BjRPLmP
VanEN+DoQYA4W7bN48ssbcD+2/b5NQoN/MHiHgmJ2uBh2M/goinypdPsoocrrMyS
kf8k7cVOmZBzxs4CngnfwsXSHFEnzq8/lA0mU+YhjDADeEAYcaLvvi/RMo1bbYOc
w2tz05WbAFTXAr/9Nl6g6aV81UpKbynQfWEhZXBzWWs2bc2TAR6kIkRbPKi6UIm1
uhdC6sDuNANNHsCV55Qx1xG7ww95P0GTtrhEjGPBJ3fCQazJI59FDrAxo4cwFqSj
mWJk5S17h5gMOHL1BSoU6FYvMi3owo8WJt1UcD6N6dbj40fdQyV7fdydhLi8kcqB
qDqKtMg3zbq3o2azkAva/QjtycRfs8kPE4eSb5o29bBP/EYpLGCsw2lUfgx3Y+xd
VOHuMHRcZcJt5DPdekcN4aeVb7SSue46GcaH/7JCdaNOiedvpF8CVcD8e1LRurni
0qU+v14kPl3EeXjY7Dhw7kNHyelvm/9d+42otlR0RmiFPNQvL8W05lHlT5ndQ3vv
5R0DSSxe3c0V+Jetm2vXvZcJemyzy4JbM1lDueIeiGkp8u3TzWvc7Zd7LdJ6R7Fo
2sEzlMwqId0pFQHQg6V4hXzlcUiCiv42y0PtP8nYRg6dDJKc6e62zsHgUZGX2zwX
2xiu9gfYfQFiDu/gu/Lu2WN3nRjKjNJskBkIHBY2lR7r3/DnSfw2NzgszsQyqHj6
J40ayD/1O7y3oscFDW+roeiPnQNXHgm598SLEzHFHTvWqTK6K7aOcBeNBm08GA1S
NrE9qznKPIAmzSG4T7E8FywpTE4qnQ+RUmTfChc46CGm+RpmyIrA6M9e9vH5tqxp
ljPn0sJL4a1y+EfU/grxqAUdzCS92P5oLosjCzxVa5pXMjZPIoGbKPRzO1t9o1T3
EUAH8eqYLdK8iZjBcRcJAnGDXxuQtht1CISRxId9tADcaxZGrEdRJqh6Mlx8vMVQ
/RMH3hDCvV/dW1l+t249mr3gSG5Ow+BSnn9FaA88fntxiPkJYZ/aHUArEvZzDaQw
WI3lmSQKyRN1C8opYMyrINti+hOHqZKbHazIwe3Gj8frGC4nQA22o84LyEY4RyVb
dbE2WL2T+9sZ8BE0FKe/ggJ7FGduxvlvbj8JTeT2L1peayyyknlRCFZj04vgU/2I
0j8fSnGh1ygY/Ix1rEcBcmplaDf4K6qxG2UMORzpX1vbZ4f5Y0AfoXPH+DaYF5uB
ehzZeybd1l+yLOZGrkBEMqiTc8stO5KHXXK9mQVAGh+Oucd2eZpbXhvGFX6EnuBy
Y1hL9ONVMdOeYNuUgg4O9LMc3ylqn0ZpTckeXvpxOvTi5+KJl8R5a5z7JOgV1UCF
PNPPcjNgaXsUFLDFiG1mrBcDoTdaTVx06ruU8Qxv7svINj3/3Nyz2GlLHdRpX4T3
+EXti8DIiVFMnWqF9felRUQ3zBrOdkNzA2vbGkGe343R5Ge5rMAb2pjx8SY7L91G
rF43927NKFzaXMLa36HazbDBLIzV0p7IPMtJ+pY0flXtcPYLPu+kcTwoFO6WegJR
okbJ2NFfiXwYrUVGVUgzv5QYFtU40Q67HG1XJaHXG1Lu7SAudHvtob+EDIetEeo7
CP9ZockK/NVuuRTN0IBnFDifeUh3mZE+Luv/R3xyzaO5Ol4mGdEZAoewZoIFIiw5
cnrxbsIezJDGNouIGxoj/UFW09juG+BO8ghSVeq9PfR4nnY16K7g4lZb/hthlBge
A3jKzXN5OH44bUMnje888EXlUZ0a/DcVh4Tr3a1uU7+mXhDVjBpbnROdhm79Amhq
t3/E618+X6pz4LVGpbcmk3T1WIcVp16utIqE/V2YwNVaiIs+Rr8Q1r5HGDkfmllC
rlnTv0qqAxfAjTHxOqwdkQiob2oEWKIobimPBvN0N0IA8aH4v0g+gqEzf52J/uSk
ZbQziAOBxTHTuNQpDOifrMTRp2sbHTc5lvdzE18ExHf2nCo75b3JDmXv21BV7ZYy
M9RW2X0fgTw5LqeUx0nbh32VXjYyOE7J9vFpkJLJZskW4iZbEaQybF7IBrkrQjSY
y8vL21k5pej2Hm1mIkMfql0zXac9pm5XzYOH/24TnW98W9MrE2ntHOHFd+04qySC
rE7ufOmKvOALVgoxmws0Kc5Cex3tN398eFjYgWLvObnQk6ZiDOLi39/WU2OoSKsZ
o8jQUBEbhm0i2JbAQzAKQ3kTz/offHIpfju2LtAL6CdAe2KoIPl1VCGKgEWn2v2J
fLxVuzh46oYFDIJwyRjAtIMsieRW63AU0riGTMsobSFPO2Qii6NFRQv7X5n6z2mX
j79ztjieluC7TPpduWcFlcVml7cmeNijH4IihcWK6p7Mo7W/Z8SqR+TXZL8V7+ls
cnJfbc16Q5gZwWGV6XKIKxpiywWg/T4Hi074gXkY9jte5oCPZp35aFswLUQAfE3y
+vvjNOugpPqTsO/N89xDu8AJyE5MmZbnWt1cDT+vAzdxN3xSEYVbc3TtTR0VP7I0
a/ty++ah/PJHNeyLbUCENEKru5ysSEiLf+akzUBuuIAXcaehkkEhYw/de4mv6MCG
CY9XrNwe1PVgLfSDZDF09GA2yMR8SgzRGurWMQXPm15jdgFSiiSIqy3mc6hRxWZv
BCczB193MH1c8KHV7NDCignSYYuhO4+ndh+YwAfsk7ARg6J4tgZYyzfXAm1aJkOj
vXG6qsEQnAB2pfBf72m7HxyAIVVVXx9G2QEyq+ZaNMI2uTbHsw7/zbJ8elB5q/yy
ETLgpy1+P/ZKf/sW+osITyI/VzvKZn9RurRanIWDk+qtA16qMVE26s1/i73iyJtA
+f04L6Dvya5yI1iqlmz80zLewOm3OkAnlS8Vj4+Fybc2PaaClXtuOh+1hE1HQ3qs
l6qc70zhuNpZMK7qGrM0Ig223oOEujrG+cQWHsSl8Cx5trisZfnAQf670vb+dP2+
DCoQjTLLBHeucIZ0buAZq7iY6nnahKG15Kw1gcpM7NBpg5keiNOJwF/1xJ5E8gsi
SQg5lhriIu/NAJ5LY8Ik4S/FucAJM2Oxy8rSzgy2UJGK/BWjXGCDRTNjmT2EbUHO
1aR/wO/a3AONWPs9JlIS6ipHse0KNOzNt9AExTIsKzWkySvZHN8TONbaRCRmu4x9
ulsM6HaW2eUdtmIypq2c76cwJL8QNzyUeW/tyoONKRQuW61AaaTZSj+C4+aiuZVb
GzqdQByGvpF3a/dTGrfqp+WhZNTJIipyxneciF5QXEJlv2xVMh9XVuC4cNe8Ggv3
IjqnguqIKLgrPOnkW8MpcrVfiermhue36RcLGMWYHRTvLo+L2eamYyepXndGSm6+
whXux1EEtaPhLhWP418MMRbk63PnUTa///lZ+dw+jq5UHJN+mnU33tgmX/8LhExp
zEidyJMInU2kz+3XalQF8TE5CxjfkIos/YkztcNEc4ubItIPXig6lS0rR4gWMecw
ZOWutzp6gCCSr4wrSBgwq+1a9GGcqGOIikszJIen0kLmeAsJrwUI4JOcrbfFe4jD
sXW2bCjlSV4JuP8gcghMkUnuP6pqNWHHpgOFutaepqkUofIAWV0vm8K9IeU8uuds
basfjvV5Svw+HtVLJUWAuKR0ZMvTB5MIwBxv/VL1nOSXNDPkPzTn4tb9zZGidc2D
vl7Bb16GJl+/fn2mPPvTIiegc8Hp0jw0HzkZEWYTSdh6ebr5zQONhMpnjHsXnmGB
hGEUWoQifOpjbYkdt51HBjrVj+ycJDH8fTyeMIyHVYfHb0+wltXqypMPTjuwVqh8
b82L3BCTDYIEHjIZghz3WOfuvShqZsJ/Y/z8qb0nQOjg651qoRbZjmAhApvGB6j2
UXnLOerBTDObzpGxvOpZCghRp41fvKWyi/dh19aBAZJ+GfjJy3H2ZdxibBw+K1Ps
5WvEC23vnqBBypy9hwfT3+uEF3VwhguRiqreJi0II/EXYX65DSgG2oFB4WwVJOub
WSH/BW2YGDOBja8VzX4NChK2DFSR2/d+2cf0Tsjr2kyRQw2V91PAHj2tTzp2sQRO
VPcDWEFCJFXxDhg5geM2j6+32ZlGBuBN4IS7OQg0iO0rlZq3tDVPvmqvq8LLXfNE
gdCfQ/OzKTVVQnzudFlja8/MjbV3o4g6BlDNxQTtK/2SlOzQLr39BP1hOzddYMrQ
P/PHHCoXUDzU5KQiH3rA2FZZtrKIjSpSzKrMySJ5xkzm4upNmBtWIsnKmZJ7DKC3
kYIJgxJPKAtxAOso0OnbCULTX4o7457zHC+EQ9KC+E58lYYdtx+9Wn4JxgiFAj1m
ct/UW+ICJjt7//Bdj8pZwk67doRGRveXMeHIfHWzGTIgbWsF5miBi+uximyuxtAq
yxFOLZEwuIl2RXdIecYMPatS0xULOV4AiPlDfN7hnBUeoe7nOKHdsEYYEMQLtmIC
lXSmhYfjCgSComdqjMeB6ZIsUOxK/zIWR9d0JQ+spnuCzILfiMIbQfejf+xOu8EQ
nQlna0rUjDQ+wa6wdeNtCfrWWKySVsnKhNg09bBg4dc46e4lSH6vNvJ+JMJC57Y9
tWiSgVOyPzNAp/kN/s5ed7klyd32+k0rXMzGM7G5EhPDASWoSCL7pzvpe1lm2u3a
ERV1iIwGdHmTku5Eux8sKU6bKgV1sTlKTp/FDYjFhZcH3U39YzoE4L+0LRMiqyoM
x2B2wed1X6CYHCh1DpLCGZoKXSe5ItNRKffzVoy5U44DycwjRuShMRIQvRWmwW+A
T0XhNvmB27LGjzkD+N0uW8ectvLejkcb/bI3Zyc3NYb4Wu4Z76ovhp9kAFC/7yE4
G/4xpmH0qeAei+PcUR6AfmNYpdknwRFWlaTBjtMR/J3t1TK+zqbDsJr3AZT7JOIu
ktXGY+9eZJQg/9PUeDNTz24NUICtFbedhnHVpXWkpuKxrjowLtTXAZI1az5n12j1
ZTuQkKVkDn//rE9MGu90q3BPN9cH53MuqhHVAo6nFLPXv7yREa9F1OsKZpkpvKfL
/GdtzavvsE4OZD3bw/h/tWf7kBElW7tXtkPTVhNwvUyKCHuXN2SB5xXtggVl5wtl
FLSnXMQyYGq6O4ynp4E2qme4BBDEmpKz5vhNYq1uxh3DwUWVHVPjXlMZBxuzHq2h
QuWfzp2idWAFOV/zco+chhLl6y8sKKzSFsf7VP6mhzMpEEz7agqKg+kXvDove+lA
w+mlEsatqBbaYZQqybwYBuWn3yAlRUawsEIkl/dti94FG7RV57rBA4cL3zBwpeiH
WVLlZ3/jNUoh81AZrQbl+jbYegex60ZFWZe9Kn5a/lDU7Yz5o6kb8tkItZmyRasl
OpTv4CyJzhvKzy44BJdB0K93ONiR30243/wXf0aI6/cDh3zm8kl9Lo8R/KzH7p9J
MsPtLTDEEPRkPCx9+lV7cI7H/R1HntEu0sKtLS4KiJZ5KlD0eLtQ5DGkGTqDhh7D
WG4SFqgnz/YA/EvGy1NOFc3EMCaZk6PrihHsI+fOKjxCIgtJcAhisdKFsLwBo3/W
QBX6tqWF8gYecfM9w7G0a4Efz3iFU8WI2lMy5pVWtmMIPjAAQFb5ZJGCjnMptta6
xIMrKGCemn+GqJuP7LXZoRZAH2dxtHuaajKiSGlZZphH0bSitg1/rBlLAkGnLBU/
PB2uTbXjPj4mgsPfbGjjIrQM+T9IZlSey2guQsjldQYovdeRtoTRi0pl7skbdNin
3u8SCSVS1ueZe4/crI9m0ty70xtjx29TNPOEAfW0lAINJaVPe1UrnB7P4IPgyA6l
1AAal83jeqfurp8Zp0Df1jAWZi36AxHTulZOYELVuFC9aXutPCCwpYeCU2nCRdhf
xJVIOJKcAzjSvA3XW7b9Q73vbuKtHFpR4ebny1OeR4e9SlOCgGP7mYuOr9xBTpgh
s2kwEVOBtxWymNFr92erEg6952N/7wVYX4owV5mC8rGmCWnApyxH0cQ9nN7VGAbL
AmcILyH4yXlLOY3zu7aSufrTF/RmYXVNIR8phJyB8+XWdnwedJECnOYk10sL/5yQ
Cd6h7qOez6rc4xZICoXAGY5JKN2pS6AJi5e9qCoA+1FgliMoTuN02HbTFuA9dSkG
4NQ4pwJ7B1l7SeGmC+W7uyWibVhrfXDiW329mg6RO8iVyEY9WvFgpW8wiEOyAUPo
A/dGrbn7lCo/tYghjyYHMw==
`pragma protect end_protected
