library verilog;
use verilog.vl_types.all;
entity and_3 is
    port(
        x               : in     vl_logic_vector(2 downto 0);
        z               : out    vl_logic
    );
end and_3;
