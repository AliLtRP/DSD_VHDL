// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:35:47 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
LxV7MK995WmS6YBV3NkBw4teBr4NEIpNuHXU2Xo2ZrxDhzH2AgxWpQ5NbndjR0tg
+D4O1fIaVLsQcTKhb8SCYM2XaD3QCzXrfABXfwFxXwqTHE4zenCfGmfcYsTWpV8J
RWUrZanW9n638skRDyyFc0qKAcRxu8USHrMYvCv2dLg=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 2448)
S6fHnOVyfZusE8LopGuwYN9bjIXJtuHVKqoMaln5XNYWp7s2RFwnPeo8DSuBS0gB
agH7RCyYBwE7RqjvUKF1irkFoQSOAKgSsYe6au38p9MMk4wS1Rub7tRJ/mEpsDdY
DpawZXsUxDSP0IesSPEALtiQRHm/S62k1jmCeS+kSc+gj/1u22fw1ZbO078MdNQZ
hH4hGtggHUYoxu3Q4S0fZE0n1jldVTQcvgAQC4lfTisyjaKI7bwGt6HuMrnzmUGW
Gt3sX3z9s1f015pfuzUTnqAc9kpRGBo6bVdw4n4/5HrgnZpZbuRJYMvE2K5q4RmT
MbcHt9wA5gJch0hxjm+xJqsU3C2JbZSzW1AExodeUzxx1SaV5g8DITqfaxeLb3Yg
VpsqJFQpTtYjfFDGF4ZhGcnimBwA+Vi0sUAvwlnFWKd+tow23hN9oWxyZ1V0K9SC
NMrGRIoRaniovVxYT0WjGDsqo01q8exLkPM6TPBvrsBDuhbBPgKXsZFK8UV7bEgm
tHtp+T0sAN8x3SbIynGv5nomSgUNZpRjRer5ZzZHH6ntp3kmlENaAwAcAO/934a3
jmNmuV/PpK/SG1Nd9VxJT56sUw5AF08pJ+qqnpqV1Yt7E3/3zZCaKy5sATRgS0h4
nbetC4Gp59oVYHGFvBzLb4y9iFe3qoYQYwcXrl/B0E35i0KnzO8Ll5btlBrrskn6
lsSCK4NoJzxnWJm+H0+4kx/l5vhD0WIvDKhEIWHJ51nhsZEl3dijKvxoMBtDNJQR
u3imvSE5f9sdcNOhPkVZLr4s45vxKcv3WsY3g8XQ3xPK2NVomQzCY7T9HUAWQqBD
2X369j3tmZEnwR4V4CETKKmmJyMrbMqlFLC59Ttbtph12Qz5YPHwz5KWyYAoxL3p
1t9TU/eZDcHOwAUcV0Y57Xzle/aBM92bu6I1HC+YGi05iMWxzJ6UtP+ZySv1JpWo
TjQ+dGmTkmoFvQHhfBPpWOKWaF2gkbbGcSqIBklYnDwNgW2dP9VB4XsfbQOtbPV2
cFfe7roSFKc/GdnKgFV3RJO31leaAQyRYTy4eLVCYFOWZIggW5DjQGNW8OI+mGb1
oJ7VqmCLcDciJvtZBGy9ukZhXEqspWqm2YkXmrgqKetvOX2KycwTfcQK9Gbpil7F
Nv018tUijmCDF0nWds7V19a+ThQoG04YuYFm1XggsHz+sMi2kFDawCA3viTzSOv/
InpiWPyc7hPabnwgzHJnQDPb8PvWRLQW5yeAExRvXdqJe70RVZbv2coKAx3HFpji
zmSpbFbSGlviz4fNhUAYV5qEgXdjyTlz/n29FBIKNbTOSSWJktKeaOU5tXPvd+Rl
BBPlf3MDbzflfn2YfZpianz1VHVC/dDKjD/z4uYglmzNcwjOsSyLeU4CoKTkuodS
I7yIySEc+Z5N+VPRCK49y4ajOSyRJbehEveaN1/ZHzFxf4yFvykAjMGGZBKMKH/l
9w3PrDrBWPNhj4FGRjlkNGY9ru1c5EOu1BFflEJURwHcNXKhsQT36KVrdtDjxc6E
pj4Af5wTbaFwnsaTIunzfkLDwQNVidPsKbSh1w/rJhxDmbJVutr89LlT/vf6+ctE
dy9/FUmZ8cZ4JH1oYGlTgYOrBj4D1YzTz2Afd+RVQOHP6yUsJcyM2qiKjtI8xqRN
rGBlvCq0JFkSF13PQoYHeGLQvJfqAaKgmiD6F4AxAK+bw7WJ95jGePOaeriKwTOp
eLOLwtxQMoBX5LgLaze4nkvmo+0iyiQ2b949M/6XjL1X8VjnvPY7oM/RQcPY1Iz2
nnrK+v8xZl7EGjakahXR2dQkCorxtmLp0hrYUcRtYqIrz2OAjf/23WHTkdlYcQVn
QV1bvMr42lGZcyYIqrc38UivqdIEKxC32KM9eGNtnIlAncGxA1+Z8QFwA4duhEup
lDYR+yMzU+l6ZiW5rHZ0ng+7RnEUYxTeGMLk8XfGBSv5SOoPaM3o7wbCfoXl5Tk0
1fXXEiXdIm9tOJO8z+RQCBCBcPqLJCM6LyFmHsYwkBjCRpwR++/KvDTJJSdVneM5
UCwHQyzrfF3laIJwl+5Sqxex4Q6fmyB+MCDfEIrflSuenT5pJyMJ0EwUvfGrkH/+
MBPpdCbBaRTilT69hyLOz2iXVBKKLkeRNGEnRv4N5i7I4Rae66svBASmJkDs9klq
Vn5X+SG1oIgJMo3x3x4GYOs6XBExFl1P336ssz5LggypkeIJbm2+tlOXsq6f2Cjj
x7DUiaKClb5wAKGTpYdViyg5gIvYwwmz9w6f79mfR0gaIOMXwHoeG9Kuuemv9fmb
5Aznn0EzyASLEXV7GUP5lem90NnsN6li4ow29SuPmu+wH4ZPWs3dfQwx4VQ/JBvn
DTvSld0lKNwt8+FKl/v6UZ2fUTMy6FuWaCDCkgIMIjQuuVmyVdFX2FcdcfJZm9rD
ket+FefQrxdhVdF2aVxKNSY6LfoJynQ7ZTyT4JpoU+y+7OQL4tO91uE6MtqfXrVO
YaUSRYMosvNY0GQYHTo0r6RzAXl6LQKoALae14BBu422ThdTrttFMT7wKfUOcg7z
7iK/giOs27N1s20PIWe3HaXOaw7seXh01tMHEAcMPFJmSbgpIe8wZ45gdYoEau9D
lOdgtSt2hKWfTgCqBYvn/0/43gm0aq7llLICF4v09/K6/xtg7zt2dq+WaeNqWnMX
2taGdOgN78GM+lFqYGj1CDiyXqiFzw6G55roj4gy8ZB5yMeJxTdbS0W/jEbRsrHj
p13SOUfn5I186oeq06Y6L4GkiFCUA3U3r3zIPNPA7Y6D0BVLpkscHpsdk3A5gv4K
fFwgLsfdn+FK9uFv0b44djvgGbTiKhRiZyt8l7dR6r8YIVNFPfMDt0xrSr1k6Rc+
cBy1AUmE4n/j6iFTS+DnSRkUZ2oUJPBv0FoEk2X/SLu56UmEX066OWH3mFOZYkqC
G4LqCGtuqGncbRZIjT2XLZHFa7510WWsVfoz2Nw/CTQ0gtDCtqqXfgPWq16Q1WN8
caOQ0XyDhUOxg/UdyFNcBC8Iyiw3eK4mOn6GlbFOeppFK1I2rt/AWNo42aPD9QQD
iVifDV4q6mavcI+STGb3ohjL/99tuNvu3cmIsxGqw5pR7gonz7aMWe7XIyAl/aRb
XvJONDDIx3CCGf8eY09bC5oXYukED4ZeC40orvMbyRSIl3qa+pBj5zjQz8Vr5205
03D/5xqovoza6cbGysuL8C5D05ziGUoTy0afZVyM1v/I7uZVafNc5U/9jUTN9X9h
`pragma protect end_protected
