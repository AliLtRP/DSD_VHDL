// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
tlyreKZPZiTIEyklKHLQgPShVGphLlIJuP9NltlkNWb2mk8NT3V+vDSBHGlYEZPyNI08jfL5reI9
ovXNvzXxBZ+Yuk4emGD4+MVZvMC+CHEwFmhHxe0cimey3CxCFEgc4pVaAnjVd4SAikoIB7dJ6eP+
erN9Hi5dTDsZhiJD8cH+sznRca39ZlAWrYgxqmT0KIVN0r7NF3q3De06+dYADB/TC3rGkuEgrjqS
KVZCT1Tc2+o5FqrMhPr5IBy8cpmYfk7aMsjigk++kNuZWPLw21mJN/RCSX5RSXogInMt/MmQlh1J
fovQQ9TGgXD6CA9UhdnargNYoBx8bgF5u5y27Q==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
YP0hnFtYYScHp95g1b41ixrKHs4lOHNnvjn1jPBVgOe86jWs+P+9nS7UnJ4qz34jIzvOmi7kj+BD
yP08yQLLPwHkK1/MHEzFLD8+UHBOBHEmfMIq5CjGfrWMPkQxQ4izGXdhqf7o+EX1B2Zl0D7duw5y
iu9KLdBGVuC6h9EjiFBxOfIiPZkk2SXIKEGR9A//+Ad1D94jEoyD0CWhLcOb9fNu4csJzSC3Meqp
Eb1DOZ0dg7x7hWf1ZLpQRzDkMBOu+yk7qGYGwfMRoPIz/2xDPcEf9i2/RTXiZUF5d9BCF2aw5Dko
3igIOBYc3iaToDnB3MEysE/nOgVs9YbIL2/VQ4paj6UyOXeRXt/W8+2nEXFd5uy09+Qh3tyKlAjz
hhnAn5mxfIGWEk4GMYf7HNHNhqnT1OLUqXcj+ZafpDloLAz78IqA5VGHesJWGbN5l5MTRWyLuwwY
dbUiUjm9ge8F5BwQPbxm9QvLI3AZZiuNfdEsf5wjLhwCEtG2t2NkY6nSchm+9V6PhVFR2EdXhbBD
pWVMI++0ZZ2qm3fVvx0+lko57vnJ3fXRwQYOA83ncf5ONqagehd4AdFxxNRmv5Z96Cd5Z60g+Mfl
bSFW9zwAxc0K6wxUnM6+v9QcuniOob3UQQ1Nk1hZyk0NqTNw7Xudy2HhFv2yEfrf5+sY/m4gd9Yh
AGJgtZtTbOqafrmiyUIPlgALJLsnQYpLxm3FOjmyXG0gKSePa2wd3fsQYREi3tTkjFcoMZ6srejc
gpXVGAUinWr93FshiVIpJePclTI7JkCVyFsqIM/sBTbaXnfj6CRZOMowaaImhYLhxuyqLyWfRUZe
XHpw4g0qRrHgpsZuPeaLqerL+cHtLiIaSFjQpyt9kV5VvK1CNnLGQRxPACaL1DfbSnABAhnLLgXR
BXj4AOa58qwOraR35mfgTvPbycHQrkBzjL+w/fmv+g9SySTrnKTEuIp1m4664fRpsxEsutJ2bEbU
vtyAb+jN90+TMpTDeg7R7MPC/RQSHfVS1LCnqTkOztvZlnD4d7WGKYOV/z9/1wUbV5WvsE7Yq2Uv
zQWeHhjS5oKiRCxbphn6ABnohtVMx6qgtipjAxCTAvXpoeFvvHxrL2yTk3kOd1FJ91314GrAh1zR
c33uOiO2E4dNiv3Wo+iP5lk4ssezfAQw51JzghFZH1F0nXVULFCHyiOwPFN2b6YShux7joLXI2Ft
Miayxj5lFzt5EapaYrRaaZUVCyxcpPeCgnkyiBQ1u9WGs6vj5AcROqH9c10cjNZtg+TSPxoE6sxH
BgmOXiENoxzyiCfDXJiBefKqJ3oKaBYORPuMR/9iJEYamhHR2qz2MdgfJtJK4ZkiMpoy5GvqhAX5
kitq3Rv4tdC0PXg2BdT6dKXLnHsVCrGJg6I0UwPgikP2aIYpQK7485hcbqn5oEcOrz0GKrOcqELK
9U7TsUA9VmdV4wOu+hAwCjAyv9D/BnG/FvAEURqci1UUKP0vWd4FqRKnbXgWAsnA9lTZWevW8tr9
prg5VELavd+IqxZwdYzjvKAUoosL2A2aAtYWzjsNATLT8WITuMNDuLbYQcWNpowcKTlximE3+yoi
IdrDqXzT2n2AvOBLcpn7F+ppI6c9gowW9ewVzmQzul4r+YAeRU6LsLmIFfrQRc4v+nMwRqyz7qTg
+/Wi2aHk2x7JUFJmDFz+YTIWspm7mi6Cehj7O3fLVIRNGiPBSZMrbxsX0/kX2yqZ6eyLHTzpoI0H
WZxQAKCEoQorGuotAwqE3wWo04aWSjez9jvZbyBeybSdpVGqTbUtcGAMUiIQP6AZYUiPVpcJ+wrq
RcahjbigdDQS7eYbunkNi1VNtzWG+usHr7AZHRUjwroAiEWafLtBr2KffKE79wpZsYjnL82/Hk2k
fFygkXi7nE8vIMrrT4gpsxU+jQgRKocT3fAvsnZWl+r/NijG7etHRLvkzdsNhwQV0o/5FyaiQmc0
5/zkQQLmPfId0PGDRxIQt9SiM3fSLvq8aSyg6yTQmYAAGp06F2yCa0XuGG7cDASRn9qjc3OkCz3s
EZMOqTHVQlOjnKMXsxbOBZa1K1kyUuF4cJsIQNhNXjSGLejOER0nsa8VZdtHi3xx8D5ZMbL44b6t
7mW+PlKR+rgxTZOqgBkZ96y9u8vhkhZyzX5XgAIXBvR6ZtufzI+zZo7ygzawrUf1lB5HRItQj3Yf
9ZtCU4x34oFZqouqX5LUt1ta49n0FM2SgrnvCB16XL2I32ux/G7uYgWXBXpmvh9XC31qdi+I0qtz
u4TiLYnrbz335KipHZIOpq+by3I/ydIQDt8SsmNUSrPtOKArRk+PSP0f1xjxPSHFstbPOMyp2AZr
F4Ehw8rnMYvT9poZqykvO19BPTPieQLiunAP/CPUXWJ7WS5HilPyQtTs37jVWg/M+d3sN+2FqQZv
KQ8sjSJWjrpbvlR6LjzdGJOtynSb119WvYCwwBHkp5ZU4htnEI3IRpKKYN4NU3Vv3urZzu0AwDbb
4IQWuXMA8VJQw3ljhoh8RxlFAoRnkewoFh1DYK/ldGe2ONamaD8nHSmD2e0lAWVOc6fD0Rsp3eFr
8B4mA75QTnXUj4K8YxHiKxJtLEEBscuVv1Qkd17JJBodOE18UTZX1Z3hmXNV3lD4qFnIPlEXSNdp
CCFSWfdCCP6YpXA05zvfsUoPTWSjMeMpOkJ6v7pvSTBhSMtg2J49HryeuH9X8hiqC7685YWDcma4
5yHjpi2sHnW8HEu1uBs9SvP0jopw/hNGSvtZ3HmtZvYYTTiib6DiSz29REU0yvGdAPN6wkN5kyEj
VppAT3DLMQdXYVYli2oc/vOoCvKl6Wv9FCMWwacZgQgCw4UEZJHXcOYVrkjMF+m0hSTjIZRNnGZS
ZxF6rtyoAXmq+5NiJApMvSdcASNEej8mALRdWWNPdwcPMM1MO2A3KaIXkD1Wuk78n2egPqhYLw30
T5S6hsOoroVR2oaHBwOgIM30FmkHaIvS2QB/grUFez1GZDQ8Zig4gc6GdTR8cd7W5ES/agg3VUdP
ztE2/vjnilDy1i5DnF3SDSd8nVyJvcOjhxHmtdZSeiVZhfaPKphrTBR3oECu5LONd/IbQctEGKU+
dsR2vr33UNey1W4FEG0YLO6un1x45RoMigi54CqYv+qBwgA7BvUNJCpvWB7c58hjuIqzZGH0ZEHt
sdtYEgsno33jpIVv8as/sHm1TDCsGLQSw+Snhi8dP9XIzzWCug5UUXZPNGWYi1o0KnwrQWrjYvF2
2kY75c3nErnh3Ty2zsALOijAxT4MH/2ltIXNSOM/btgW93wg3FrIc/q8Op/4qUb0304IZe4Coj1v
pJdcA7PWzrj7eX2KcN4yCswUsvfpcQ79liaXjhiarI1cXnZg9gcNl3iN9fyy2MmicD7CG5UrGJ8g
6c72p9Aesr9CZ8j0kxd0VZQ0OqifyJLwrOjVQYqiMp1KNxfyptaRkBuLN3JIRh4/EGe46kkvrsnp
Wl4H0qvh+g4soj08PUuvXdHlOkI+3PtDoQNjBzIBuI2/r2NhUk0+NWfafZMCjfX8ODCaqB+TWdWp
5rn4FlB9LpJbMo+WpyBpibrFJ4+1r0NYhOlw7PdgyuSaJ3GqB27O/gdUU7v3fiaL3lisMhz7gnHh
1dnjtlIg9rD0WVFMHcb3bkZJFbRVJvzTOanh8CJRVKHe6O4wjweEUWcY5QVbdHRvc4RG8gz7kpgr
zjduUiawjLPLvu9x3vhKVxhbSO7dpuS1zFhhXEiK37neC5wbtJP2lCp8plEmkdl98eoJAgCfJgNB
tkUcwN4p+VbxjYoiXxaZjezqoe7RQ5iFMhJozyGlkh5Mq0n9x5wO2MIqsX64j35Zs+M7dTlprF4M
3Ua8vKpXMfHAo+vwQ16x+LrxdxwZCqkPinSF4/tUEm0hEimRURKRvaNVEXW45EXP2OWTe4J7UkoD
Cxt1JqsftUmPU+kwIEdt4vJmOO6EnQrWWkZYWRRFd8F6daEwchRRgveTDu1gQ34RaPAeG5052wfX
vF+l6QrrwRSyBIk5bVkkIjEzz70yCWZHGsDRz8nJMSbELJsuOGP/by6F3JINfUFZf4/u+Eqg3r5f
KuckgNQIbKeeNOcMmGUQgads0oA2oxqcgRG/78Ie80EoqpjPsEbuBibcwCXtCMyBlhGuBIDDhj9E
R0+oHCg+1r7NUF0jXbo3c7HB0V7fa0jZJ3PGMydpeREoJTLVBdH7VMJFc9dOEkefUhSLNULXz0J3
TLar+ZUfCE5uEUmNMQCh+wwK208Z2yHe5w0tHFN5cADST/zpADsl4kU9sAGPCKOBa1mBK8dk0uMJ
iwMBTPRmgn01ZMyc4oh/7/6osnZNBgUXBv8eJeoXJj0b557AyOExdxp03kR+zafr+DQHvosCI3UF
FLcGKvTl3H3WIphT1O2cdnWhcQI/k6D1IxQk+SbHfrqHc3SE0Vjvru2ynrmf2kmtwH7q+ROBwMNG
z8uL51GStw3GK9mqXGMnVxwIU1Kex/c4JzLxAHOB9A0HAArkqm9centvc0ftaS3+2WfDMJnHEEoV
B4e8cWrBTbj38a6YWFLuZBxZlilfO2dCjcXEInfOyLH8e8X4TMRpHkLu+y4AmbBEi0cp1EO5yT4F
jPx1w9XXav0FSuwqNkPc40yp9xoedv/qEBQhACTWNdVNcz6Luriha5HmWOGZRX2tuOFGoUdSCQUQ
9Xtlk0Ipwe3M4y1rDmrAh4z8FJF9KgY9UZpxB81RvlXMYTeeNrnqctvoyVvsh5wt3qdHWg7l2a6O
0jkh1MPFMjN/eNbV9QhN49CNLwMQcYDBpJnBffcPRuDL20BYwcZZDxdMMC/XP6k5CD1yeE/sNcs3
aTt/JQ6wVdLMZkydFIhs/HrXh6Hv6oiXSi2Z/OckocZzG9Ss5gw2quSk5+PsKMYtqOcBzKQ4dFur
3AJTmvd8vDJBZRH3TMWE24v87zasDfxTyj//LXzof2ogMI3rDhEJiRuINSLYDnFoGTUjPnW+5mSL
AlRKhAmMKOyvgrUj1B8knJbaMpTKcyzmsvATEuJ/MDbafMjIRi3pM06kAeJeutJyqTqJDBfNb6ci
P+dEKxXLYKTI3xDCJ/LynE4nZHNp+UP1fisIscXElyF/crs4dlzKEtAWvBLZlKfqLjW3OlxPZGND
UKD8MBRxsWCWA+nH/2H+933kPKMRfWK6kQJPVsNEf9kyACALaj/5GEitMggSpUVucQbgr1hnO4FI
EFZGHiCmJwLX6Vx7Zq68ApLWAJFNI27K7j3OffpjSqFjzC5y5ya9wbM8DzbhJNB7PnNEWUqGY5/Z
DsPJFLXS9Ty2wgUUwQoTSsPvGnYvIJl2uHpqIuuBeJTBswuKh/JpExDoTUUj+4m3+/bNgC/ObFmW
nXa2F7K0w+gKkQ0h19tvgFvNcuUjI9OaBAMLD1tzwZyDTku2y7WDAzNzVBVkPfqK54FZ46zsWz9Z
HrmEmueD9pBJ/uOvUAjDKv+xUUDFaIqcOFCvmMtojN9fcPB6a4c/Z7SerIoD8lTbf2khX0cOz/u7
Y0YjEds2BCdr+JysvDvxe14lLxikocTYI2noAeFV3dQ1z0t+VYYs7f2PC92BXLT6VF0HGsc36Kcc
0pO2hStXGUhlxaoIdXSE4l0BiTLRdaBJdxU9r+ceFG03H9jNJgf1ol36Hw0gbJTev57na/AXAE5j
sPOIBfZh0vEetAQwoh8RYdC5sXcEDxnr4Z1Mge4avFFFqDy316dzg1oH/hwbPFGuFvGttjgblJgk
IjbQ1oXosC5x4X10c5U6KZrfApP7AhTWWn3bAIE5GzGEh9sVcu73KFmHRoWqeIcWjmQJur2pMQ/Y
6BknPapxZ8qQPiGxLrhs55CR3bIT05ZkyqplG9PH8KAx/y7dRbICk8NQHYZJeDYQVw45YTgwW0iE
l5k+m3ZPkjVXlgLHIgeDAMvz5mxWPQY62ZtLuThXExmBaAp8Rxtf4Cso02AOWAKFOT74SZ78Epsg
hnGXsLLONsmGvdjqop7biIIiUxvzhifnX2et4+TatJfSxIv1KMPE2im8GAkDNIYBbiSSzLN8zEhA
h1ys5Z8wu606Cky7fCS8WRFxd4jMbP5OIAi5JZ4IBLlKBNDutokuHkObrE/D1ErTzORI5pC29/4z
9DwUuhvjvCFHZEtZmFWjbq+754MWwVSyLcOOmyYPvtbdQrX6/h7uZzRO+5sOH4TKec5fV+U0McoV
6MH6PQp9yxEPMz8U9fb3ogdtjzLq2ig4MxCR0/hGQiGlzI2ErzFKTgtNN8Kh++shKql8kG9LqxmB
rKVuJTmirbCPsc2eDzztHz/0a8qUaFvlX91vK2tUjWq/UxjoEuKMANuIdEpySJXQaSGnD7a2oSxz
D2vCyE0V/02Lt/++r8E63qVYYES5jxg6ZTQbz6trMrpkJbJD5LRLAFrrtx+cI7LM5B6c72icAivV
3FDRBsYH177jL6oFtBITXcARJWHIgxd1GebZsjWh2R8PoZxpMcJ0mZQjD9wG9STA+GqYvN6mI0IX
PmeMETXSb22HyBYYjNxgUJAenf7scn7ip0THWFhPDWIvye19IPMmXMGmMdep/U67R3wwq/rG7hmZ
g+eTGxgYlYpGn9EvDx01lV9MrMm6KaYMC7WEOorNmrKoA0HY60oZRH70HxEpi7I2vZ1K+OB1Jfy/
hWnw3Qutim01/Kv/M2zyTVm58gvZyg8Mke91K2M6oL5sOwH7TrHZRN+/OLgcmlLZOPBGYeLGsSUp
pUTKGWQBEVS8qxJBgbTksIvOuF56EuU2JDFw67O/BSx6zeMxi4QszBymbcxQXUKq21L0cGHoNoAR
sikukTsrTQQS9tQygkkFd4fqQ6C/XqbqMNFS1TKkXTr1jr2zpqt3Ne1vE33KvzfUgdM+vqsnW2Mj
HtpUjp5ajQG4uQkofHfCWr/kIzBu6jJwu1UPIDNPTwjJVrwiYBhaWvIdwE+QhcUFOoLJFHnRv9pp
2EeHA74XjSyt9g6IMekIsoZ4hsUFKj865dz5OxTYZztS6GypEnfvuNg4nhYKm20tFiOXheWb5bvj
HGzIM96Q+HRjPzx31RhQIx1M2FRCo85NFtGcosgxB/Y5McgtVV91zgwheyFUcuuIYOI9GbwBQF1q
lKmvmn8GEh1EeuDlxsqYFpmwkMdYU6jqnRNWCM0D/Apu2zu5YVged6mzcrMCXU1sbQ5hXN5LRjAw
OoiHuRKb+m83NJ/OrPspRX0mVJxuSHfBbXmoRxrs2h4EpLRdNVTsu2PedH8KaSO4pmW6ekYf1oKJ
ANnELBX4wJic/JsU9CVqPt48OBFSJgAtvPiO2a0v0aFl+wuNmB4gAQFsVP3icsnBs1OL8Y/nPeAe
0xKMyIZaoAyYBjy1RrGquUr6D26g4oyqRfMISj5Q82ZIZmUJzu7r1CzXfe7VqhQtj3Za/yWOekNr
+3j7LEbvKFi4PJ5DTdMfCTbwEuuKSsg/TZPnx5Ebnj2Bf51UaTx87+RZ/t3HQOFrkEaoWxfCKl1q
oVNFrKawN/EspU++kVYY2ZDiWrd1//Hxv9eSZvfEKM4XlA0MtbHGubUl0WISxK7hcsHvScy9oMKY
7Cw8XBU5+FSsv96/ZBTUtAVk7urSPTx8aQlcgaw6NI2b5cpAmWc8kDjM4lf4A5cdEAbBf6e0Ck/m
qB38zMKV2XtJBwySESfoY3QqSEHWL/bI+fZD1oNVjfCE35Qzwnv0/2c0JPWM0PPfZmhfuE28XS9F
e6EjNSxpq8/yfUUVxes3DxImUAGFLOIguVs0RgbQ/QVmhx7GiBruG4oaks2xIIpCS+vjJg9p3O+w
1Lz0duzOJg2LtrG9I0AJ/a1AHOzrw34pmIxG0mnPMOOxNAyZujZ8obuSAEgnSUFZSlIEd6mTIvsp
xXX7jKl96OqQ/ovxoQroG7+Kl2TtqVYETd1ua7sl/fn3MnhWA6FWx9vyf/p1IePRKqisUE2JBwX8
6TEFSLSale5JUTMQQWiciaKmpt3MHztl2gtrLajh7shXYPjJxUCQSCHn+OFH7qPJAKtm9fmiNyXN
soFOLG7D9yBEWc0Xgmq3NplNdI6O7VifOOJ0Kq/Ua0qXd95T6Hua33yi+fmtD7HHHL1L71Y8gA2x
UPQtpUjbbtMmDA3dJXXIIUvxVwmHIF1B0abRYHUcZE24DJMOcIlGxKZHDgCh/sG84oRozHoKn2tW
c3BhawL7BVGBrVmEF2Jak4abaiTs2aukO+3z3yhRc+aJPyBn5G7AB2sBkmRchKpYNcaLbcyVFfXX
kxjZcXfNmqvSQMW0dAwbvKMSMwGxKo62rtofoDQmS+0hGjxyR6BIHgqTk0kSk/YyaXgCbJpUuGqv
MxzqAmn8UNFLb99aYRMj71bjumdTKwb/4phdlRqySviw4YPNEOcCCkk3IBALT4z79z7w7UqZS9KB
VDGXAflXOkNa/XschcRibNPgWTqwvfMnOwg8bv4A/LYCJ6mu/kRgr52DRRmEVS+nGf7xtdkD4+DQ
5BOfGTtHvh2dAaGf6IFHC+XYwfjyL2hlm5C6Eqk6v4zP2ifdb61U7DzAS6Id2kQX20RANWjphb6y
dU6UxJ6691Oz+bFpSvcmDPIo0WWTPZnO2A+WokYGdHBfg6jiqEP4Fvi5931bRsrr941uXCPTEHWF
p+IWzJBJOxlwE+EaaEKRsFaa6AJbumqJp5WRorPqGKLgLO11vZTVoofEeki1F2Df0KY1ifL8ktl0
zQdREtkDjXa//mZBUEywbw4Mbj8/y8Eh1PdrN3yBkkHpNECES4X7EofXkuDDEyS6J7a4k07IJerS
qlqAvhad7eNSi4C8yhHMv/Lw+x12U0CtSryIbRyzk86ZdjubmmVs+Ua3W9TQLpLTWrup4fXy73+H
v8W/r/xqjDQEVpOBAs+McPLyuFJ/c2TQWjqUZMozGO0BeZTu4JqXjVh4oUBiIzyQMPh1dEC/fFUZ
6U1zHigYJLe2lGhfqKaRpBZ6MAMfmlqJkN0QrgxzJOLrrmFzFpObDJjHp+cZ0XufDfs2cnXia4Im
3mYpFyhCTesdna9/rmPtlqcrrc9omxKPlTwC0zFId8jhxzLZ9TRdoomCHFCb/hx5Bjfy6wyb8kb9
BmymSfEdYX3nXScEhZ2c635CEx5onruZoEm9jIhWuT6wXgSeL39o2Xu1uvyl6prgKJaKGXf5IFFJ
R/CzOu7XdyabsZQM+QJ/JKjl4ovEod2Mi9tyLslLrEcJfa4UInVlpJBsNcDzIGA1KykHZgAHiRe9
jJuLy+/foMfgNKnhfzUpmCtIU8gofwlRk9Lm1TnIhcnrQmy2afKjk8M+HdwBmfTOHFDWF0HdkSDa
fhs+KGIoExgmb1U1ycMIrr55Hw2aKs/06y0zcNkNNL+2cn76Fct6JiI4kvF3G7MatFHI1K9JSQJj
nidzJ+PtMhvMSK8v6CTerne1iGPfAhayUVcq6JIDiqHmVnBrHUOzaFQW5vjKxGbV+D1CPeiEUiCi
QqMjIvuIlQU9JSa2AMkyOc2/JxeUJraps8douFxFmNqnDo3Cdwggq7LSGdPaYvh2MgdAWHNamgFN
bkNklNKkDLSetvBI2FP28cBRMysZrpsVLD7ACbuLffjnyou+FU8/Si1C4MAsjGRp+5Kctgv9qrVM
xTHj0cIr6ITQRRl0PMogd05BUg5NtRKYFIfZsnv2Vm+8DkWuP2Ai4jFPu+qrOPJ9a3EYzz22EIeO
zArvIjVuFrtsd8wgkBMXtOePpVE7ScNVF+e9DWr95Un2oj7Af+zaosr+dY/evasCGAgTdlu9aGjp
ZrS2dgVXWumpKEX+Oazz1EZBmHakRxQpAO1uVR1tVJ3XwweFCN7KipLLKT1TkzMJkpvRTUP3ZhCZ
ZfHPNMPRZMZ48Ol5SPkhICXS32cbv76HVWFrTWZsiLX5eD3PsKPr34RdsvvkYnkF18lvQ/hQ9U65
vouZLGHyrxvHfh0J7NZju4PQFgidb9m8qZzkY4X1ZWjzk+c02W5UlyEPsugivRkXG2FRec/IIUZK
GY3imn4OhlBi8EP+Wg6kXuKZQYnImNbPEjkOk4+ClS1M/CoUNfGRZP7Zc+AFrYL62IZvqZ8g0IuD
DHk7Q/DrLnglndKsh1R3ImlT1OuH4yfWvWSxkJVMd73+TMIspOyFfUMJlEmfjo2NWlrCF+BaZRjr
Uonmc/59Foa91H59ncLog3FyegfH4QjwXtLBzK6EQksSJNNS9NuyNlq4pt3d2YlnCBdxS22JrXGP
4SDQMvPrHQez1R5KpwoqFQWtdSB8NgRTDj8dq+wu7Z4M4Fc/UTHVyMlgINnQ30vFya9cjPrIIoOk
B0KpS55K1gwFXT14R7UCWHncaRZqCJeujHcZhKWWbxNk2PqMZSpmBaKj5yYH/JW86F0H1D3xjIZB
kMYAksBIQjH5KZibhDde/oR2zz2ydNheYYsn2ecTMIEUVWkCsOe+gg6skmV0iNnpKuuEUs4+XDUV
J0fM9mVSA4vNuPAMHtWVpsja7OPVWQNBzU0y/2VU3YJtqUJy1eSMvmSOA/gC1BwF7jaZkUojR1Vx
fjH5yC1HqcLrG/e5ZqcCCaxk9RUoAmkLd5qz+fMd57Co95VgRdmzI9HYXXivczcda6I3h/2eoFqf
tRIzfM6TZcSb72QDdXh7HsKgoF608k/HbdByWww9zEjdh135YpLg+HwssZADbEoRJ2z/Te0sBKiC
bk/MyPo6PTcl24RyeZzg1H6ZA4LI1uvn+EZ4qCJicB2YpLo5jlkKQul8LW7B5gLuKZn1zt0orZGX
6UDjvMHIKU9Zp3zj79qVBwqIH46nPmnAFYNKQoklxuI/Q7jkMM4Rqmp+LOTA59LzVrxZsPgAkfvX
NS2pxKCdkwLXDpkL/lV1zPf3vL5XwKii9h7YnQaQG8CJhaGrSIc3bs0mHjJLgtXpJ8OSP/X2EL2t
SezkkAuYVLn4Xe+fs13iZKN8SPLMhx20ZKA6UebP/hUUIu4iIS0J6bowkTmF7VvahJi3Q9ZgW41F
hGQQO9eaBBluQ1q0xRMv/Szqc0m9cLH2hxhl85PnKPbgfDL5V3g0M+ces2bbbnBRRdPRsiUSDI+3
D7cjRaZVjEIGqYpd5mroatcT8vW8wDO5Nbux5LaUaS4u/99udDluUpuyf7FOuy6j++ZLJ71tQY6c
0xsZuI8fCMxWvKB/KYnyBUMM9SFYnUf6k1VJE/XI89uCxz5+9AdMBmZ0ANQfUwLqYYZNNUkn6Cwc
OTpIGlMQYVgJG7kO5t5vp4J2rrvd2oV7V8cMjsKMeKN6sTWwrGaxqYMVxr0RKuVsy6RgZWGenJPM
IgU95MAuj4K4nSggrJk6N1SDjD6h5coFkwTS0lMhiCiREtBFj0ovz5oPEeJuTW7sA7aReFor3SG/
RI8kLuwBQxi5TEmAypesyRrin7+yVd9sR+xfLY2gEJ4m88/sWWb3qZQ7Nk7s7MRVaRJx13m0Xk2L
Y/b7PreLfpfYVSeeKe9PREwYe70ixZrmTKvw4IO/KgYby93t/1AtHIXvabNHwepttSgJQOWtR+V6
4D8iwAsoEzsBt+cDz+3+QqMpxAz60dUFdJBNIfN+Y9qHwFpMPyG9aSBFEoPGCyGi7VmmTF2JWDYS
rocB2JjYfh56uDI7B2p+1vn/q0l01bt78djs1Z4B2p7B8xoss0OidGfJRRTW8+d1bSoh0VelN7Lq
gZC6+0AjXyPS+t1+/+vVAZy92nsJQwmg3y091vNlu8DtWIufd21JQJth5jbyQyQlQ0iSRLA4b8Aj
g6wMh8MQxLcryceLoSBQbX2Z+cYUGs6Fog9EljrokoKvMVCduYohwPC2+gorJrAicTtmVlU5VaNg
iZ+cuIXn0chtMe4BdRS0ufM+kgaC6g9QjJ615AyJtoDttx06YiENTmq0uvvm+b4Rh8K7L9s5Jsxs
j2epcvZCbOauB8J6s7NLtFHYt9uZMELpZu64S+KnZZyI7cZ6+YLSQIw6OtSwyUl6bYUUXtLlWYK9
FTUWsUq9aP5a6iq8vMhrPAq2aZlre2Up6tMQO1WrUixG26ELYxygm1Dr1M9OGC6yMT2+cqaerw1Q
nF9hKNqWygiGX03WUSg4yYnvichPssqysEIFASsAVu5axVcCAKEmQcqwWOkOJ1yUYGjR1r48u7qE
6Posb1sidqB/a1cc/FdVQkQn2/AVqTLxfHbzQA/I9N3yR6SJhr6wVUMaFp6aqyDNXoaOpwAEMqVI
cM/7f0TweD31qzPwmaelCu98hoGvvjv4PAnHObB4yTi6f0h+ei4I48mgNajvWJNE9OGmtJKS3GwK
Ii7ZlqAmn/uw758oaHszkHBqfKfqUH31r5Y3L5DzG7tqj1sFXPAEkDpy0RVXzuJ+fW6b/j3V+Pny
SJsuhy1wyHaToPD0OOQEWA6IpyHO/8Y0e6oDcIPq/8ge88q4KI4u+01BcdkoK2NlmpFmbZ8z94UN
ct05bb5t2KFPWcZWNCDPKiL8v/PwNQaxTf48Ax/lvPZ8DbfxWj5J/95la9STxEovjhRz9EXrptDr
/orZL1VSqQmVUS6jZBCIdBLubaX5QDMumDMWGkjvv/zmq4O0uZH61vn+izNtLgkekJsDJ3Z9h7hY
j8ZsaomAKZ3eV7qVStvRnhCPWyg33bWmxwWQQlQlw+Aaz9f4qFxfFWbpzzyGFlROwVvcaJe1FphY
ov9jXodJWCJ8rz9RIbJzs6jfuvSqV9wwkwQoJI/PUSAAI448+6xvhuglU2oMh7ApmYYova9RDZ2p
d3Lp6vDRKmV3A7b8JYOxhUkzKcPQOb2tZtwBaifWJ+vFen0WjJxz2LBYtRhfInstLn0lM9ElHPbf
PN9DAaZUDEds0fsEm0kngmRMw+/fizX4wM5QM+9AfC8/2u/r132N/I5ZMAPsD7HCGOmMjeY562KM
QXfz0dG1E7KiuSS6UGulXWv7bTRO1W+fg3p3Qc7SliO3YDHKdESBCrn5tAEqOQbZC54JiwoXLGaq
7H0+WcQnXxGCTrx+s7HeqBZv2oAQQswouGI7Qk+YgnHoZIwrCeQ0xFM2nPRNXSBVcXXnWIjmYvM1
1LoS8FXt44vqk1EO9sW8+cahamP5ry5zDkeE0Hj29mek3KVo7frc7lP2DfFl3AnqaEt1KkRnZ69w
H/Ner1RnmSQF7H+3ETCYjoecMaZd320cATFxOOtpSDblY1YKvVRD4saGb4QAyhPGMOHUy/gZRelR
RcD3D5wznsavWv2K0UMcWehItCfSp6fygvhYi5N9rwCyshPeIuN/twit5IDlanA5SsLNRo0gW1+7
J9oTDzevUOEIDfss2OMrrw4AzGy0fQejDxTAkepzw/Y+RKvSkZ8rX0ICsGSssByFdaCVQd7vAXEd
s3n+vbiNWUfqWnybkIABOmt5GnHYzbMioN8sOZRCDbqHvvUqe5cj4Ep6zMojjp+4VYj1Wo9Hh2qO
jSLn36NI3PFRkLD0HlyiH7eoaqQ81l32NjBewDCCcj2xeE3Z0Y4hfEx+Ovbi3mG3Yi/e7vfzGSGr
TikkRXJ3SLHMsAS80qiS8tKfj8NMNbeTKOtPSJupswF+FrVzr/ovIBnREx4JUuOWmq2un7HNQ3O2
PEdZFJx4Tu6TJaswR4n53qvQh2gUv/u/i+ITrTpgAAbhDi7+nUBvESm3pzB65yMwj2TISfv4Z3IY
RJZgMEHXYyZe+zUdigiU8nuAmvX2N3c/GEZjRzLoUaEVWL0I+dArFCJEuZNFA2qBIFcMvo3nEMsF
qdZbejTByDG+eLEbJxESJrrz3SGb6K99tisnGyomidpLaaS+eKGFiarD6wgF+dIrfkB2eEq/G3LA
bcgNTDkAhMw/lPz0syT+F8q0rdvdxMNvhaXZln49fuZ8Xdl7j4PdD9cbx+8rKve8+1CpDglqSHDn
3AIP2KyIcwZiUBzQEBtyQxRSAI8JcVwwCbLqR7V6iW/T6Z5XGaVSzdoKo8w2rUSMOdnJsPR+nCvH
Jq5XxHFuWD4NRNkFLnL4bZtLL5o75sau7H1qQkRSlK48a0JyqQWFfWcu6m6PylAFcQRqpKETNaMx
USnqHmforTIr8dpsfRMADPSVvTj79COJCbyoZhaWpgcLGEZvaruh2gOqLQJucYFgYM8wVc4/+8K9
RWprmD1e4wGiWjlrJJs523uMOlgK5ShiVIHQOXLnOoBdxmGBmV+j1swWak1xUNel5n/3I625BwoB
u/tJPlR1XIL3kDHYYdULPj2IoDtJQ8zrFGw3sSlFbtzVvI/blhNFahHFeHNHvz8p+KY0NPuDwl48
0aSuwo2NwxbGSOw5CFZka6Q3vbcaJXlACmTSYfFzvLTtWZEc4gbcndKo/rXmd1/Mbr6Thfiu/OoT
nBTBmebSfVAlqUAO9oBzTmuy99tbr7aCGs2r1vQZRZAcQ/mvqUw+q72oATDKXVo53ztFvSbDtUEe
UnN1AF/97W9S+o6DkK5spAvJ8AYQu2KqrTIZYsLIpp3T//Qj+To25sLrxhxvrupr/U6gxui71FT6
kGHJuEthzmz6zp0F5fMUbawd2BhpJO2iGzH7e7Z7ewSWWKoYloG3vZeR3DVBs3Wb840g2saxNLbw
T1rfss0Nh00JIIvtpy0yWrpwUaJgz0MYgpmqQ0lycT8jL0umLCC5m7ow15SCeLSf5L2JUxfS6w5G
3Dd3m0GvoqpzXYeGbIcYY/QBfVWLDzH5bbUhovxNSLSDqBV4z5ilgyFURo11HizFEd2wbBpVHdtj
PuMln0eJILq5HA8XI5G+N68XbJaV4vZQBkfi+0YUwUSWjQ4fGRGlLH1rKFXR2abTxxeFaM987B7L
bmGZW3hfzqT72Ndm2+lM3VNMOwqlSvMyl3I5UQ7SHJW05UvtoxjZlxC7/W1NPR/ulrKPh9GheRDj
aigHd1tvtXhwuSf6UgVxgVklubmg9u7AAE13IbVWWMMW9iHMIr3m1u3LH1q+VO4L/NttajvH7Vaw
QVwL4uCtcuu+11AK6AW1RtwdV5aWcrne+VD8FDpNTsIlJpTHSDgewvzJb7DaMDt6+4CtLbIwZoU0
YKTOysp5iLrwtsgpP6pXmuDv3phXNU1OrTmwPW8ofS74IuI/lfYiP8Q3Jrd3P6GACVYdAMcqrRns
9/oef+2pKi9qtBZTOg/q4kFtifZuA0EUH0VbLowKhrYobyfKzIUSfGkSsLOeW0cUuvM8sk9l9QSD
crG6rREPUnNqurfBVXqeKGTfqeGh1zBdqRGIzcw9kGZ009EYmJOQ58uEjG3Z88kgyFbzcUxiwGFN
SEadMpIdd5yOWLWTuspY9gctAAtR7ZQsG4WARXi5u+5eFoqwmhuBJvxwj1g3fuee6aucFPdr2H68
ic55LrHeyyoONA2TzYXCBrlUw/TxptZctoScEM1IRhj+CjKhNyYmgfE/t29uDQYaT11owfidUz8v
/WPW6RQJ0fdlZMHE1gLraVylx00hRDno2Yf2M5OAaK5oB/TTjoWcXAAgGT5LLr3dWCxM4ur/7K0O
EC5KctnEzRQgb7I3NN2C/O22n4WYelopugGY64A4qEn3Jrv6f6isIEi2h3IP1WVKwuGd61bEwsQ3
MJsd7+EeKgPjRGN3GqQ2mYrd2YJIPI7tHyWsJhxh8nLvdPNx7S5nl2aJSGxhL5a1zuOfUC3xlSdR
SKOiJ2T58OID7cIiGib79rYODUW7uWT/4WHXTpRj1uZDb2RQBfbPXOiuVQx6VROn9ZrxdF5B+7vI
cor1tJBpBRAYlEe5EW/uRUFAMOXrOPdcCVJ9KbRkSGL40bhFO15Rns9qHqTfmy+cI+IBEIMgiYBb
O3kvzy9ABNETQyVMw4AqebTIlQOQndXytyAd5vfhYV5CKKno/pCeD7JotOla79sKsnAavaWN52A4
Hmnr9KsnFaDsGSmyRr/nFUsA8yp34y2xk1jz3rfcZG7aLI05TBoKPT1MOJfbuTA0eVCT0VhF5D8l
L+YXgKrGSup760l8A/fy9R/yDGucAvgxHfGPE1c0gmFA6vXcXPyiTbK5Jlx4NXq3LimCo3zc1dYt
gejhLuQr2EOP7+9u9bucuLzTo801IZdpSUn9tIYEtOvZ6cQlNz2MMU3N+H5WDn2wPCc89kRBty/5
iUfG9X9usuZZZlKM87hfxlDgHg6J7XHcU0WNuSKVDPQGLjWD9UF3mGgH7Andclsg06mWqPpRWydG
/rGSYZsL1A6ReXrQHtVGbLKZElBwWeMBHRnjoY1zRxo+Cuwm2pniPR3KqK5hcIoRaafzWxwNk9ej
Zulx5lkmzKbxalR0FkXPQ5Sei74+Hk7k2wmo/oE71XU/Mo8HLQIUaVFnnk9gIx5rxy2W5XOkv0uO
8wrvGpEIXVhEVDxn+WqIQJoAg6DtibQvsn4xsKAGVZxgZfyGNS/0FpZVNF+eBQTZsJU09sGIQsLW
GAs5aq3FltM9JEp+rrXBrC0Naoa6rB6tsMvHBnY/2M5U/WEvmDp0+i/IAS/hw07GpX6N3pxMNaDO
8CCOq2dvjKCi/Y4yC/ItggiEm3AzgHXnJk+xBqWYjnW4cOrGny40MSYy+U/M+KAcBK4MdmhKwfBh
U0m8GNS0mNGwiQeYMxpcDPfJiVdSjn10IpXlAU5Tv9Cw3huluTd9URkPlRGSUC3NH6zj9XvRbBLX
A5ni5Bm4z0efOQFomEddNidRyAkF6cG9o1t+c8uqJDLoMrc9eApU2Dua/l2Y2DmBVYXucm1y/2aI
RSnMO2Dj3BjcD5mAFT8smh47OSrUKU+P2Msx8fAV+Vv58H7UyxWLMKWl+KcM70TMzYtHnL1J+p5H
5HTXv3I6xwVFiIUiNxWe5yxCS0dQODV467h+h7JlC5g/o3KQHeGV/t7FTs/+PJD59a3z9Zb5banh
wzJfSb/KKgJYdIGOGpwI4FKeiqEnv7ypLFdLGmLVnQ/XnVLGu+9xAw2NieALy/WOS6AfOCvxstNs
mlZhbdDJBKMDzrBm+ztaH7sy0ti1hy4KjAGbqUTmsODIHOHjvfvF/wAiDLXsJ1Y39d8VGqeNUINa
33bRh2JBVZO0fWxEbqk2ChwQNuJl793iPb6KXvVEv0dcCK9PEKXUxsrjHEKV8JpgjoGwFO4a4TW6
42lah1EBCKbPfcl9DqJdLrI1S5jBZDyqfBMKso4zS4fPulMZDZwWc/mcpZLJBYjVMkKd+Bc9JfWV
8t+lrBmCaNSaZY0ZuzDFpv2oBOaLrfkpepr/jcbQq7gCal4XUTpbvlOWJrU3ne7ZzFn4BJOYfXMJ
+GSrUvgQsqeQ+y9J1qNbRIaNIbR62bnSL+YxNrO3nxW7opHzfOgOLoZ7YdJwhJlbeP+VfCJhT/xm
zjaPdcE6nCRfN745SPRd+eVgP7XnCS/CAjKX/tdwI929tKoYdbWY0NqHEbk1/eqGP7X/UxYnJY/S
B+bF5Azu4lgYZP1QLtJO08ISTWAjxnssHOrl3X1WMVOPXGA1Ys5pRm51zcwMz1l5/6tVgF9v47oT
orgrBHJdOl4HSO+IEq2UxU9WLW0VV1BWxAsC5v5lNF8Oq9Z3eX+KcgSMlMYMuJFjt+J6n3gHSOlR
NGNe+bWWxqEP1jw+Rxhuc4HadxnJ9tYNR4wei9ll89mfVS9beZ70160WLAwfgtAXURePkynnkW+2
pqaiHvcqX20DjPjnX/Zf6ZcVlxMF42NfdwG3p+vpwZ+fatWORrsHoJESoFGtsdQF3m93hjVoTgxL
OzD6ueynMfhdFi8CHwWXUWzkJdHz84UgKZ+y7z6X+3nI36mfKbwKqPQG2v+NYI/ZW0kZgkzTBXvF
UC/KJDzs7qTCh1Q+cpb7FJsJ5QuQxVrXrkS26nnW7j0lInWHBVl6DikTYBIKs2FYvuw/yOi8ogBB
mBt8JNoy1Q/hrOqX5DBg5hWx3TSN9EYFL1570eDrhfkIfAOR1YJNYYFDtBsHrsg/ntDR3gWfZvSq
btKx3lbbD996a/djs4wkLZ+sa2EzzuGEJmWYn09c7NIDHTHq/oXtpZSdXqneu0+GF5dc6fvyPrg/
0ZFHvMyxCruvvdHjEq1U+1VCrdbAZwh9RWP7p4fCrpur+abFjhTp+C7uWfqZKfPuCzohafXJrDTh
R14a4P17rJLnwsBZ0TTv2VdyUbaf0esKsAV4DC+Dc/YlF+myFsDDs0ITROtJTGwgtHv9sNDqchgN
QZk1AQ5wkDTKIvNAHCuYKL02QqxpnCbibwYK5vzAX8kPcUXnTTm92Ueqh7cXLQUFf+EoZMzEzm6p
WtF5Q1VqtAHS3Nx6/rYP8j/F155iCVX3aEilutbEtlPF1OyaLgiDTJ/eEvYQGrfnCQngWUZkJIMM
hjy2G0WmA29hP5XtU3QMyZV3oOYC1+Vgkz1gJcPad7uYpxfVJz6f4ZWZAljGVSX68dX9r5OJL5gC
I38Is3BVEJT52Z0j7nZiEUG0LCzLK846KmB9eIe3OLvyMndqrN4I8REYIosX+vpgJMl47kfFrcYa
0IBuin2Zobk+Yw6EzaT6kz4w0tso3KXIinpiBnonzVRa+0FWn1AvgDSuO25ekh2AYBX00IpE7u71
nqC/kVQ0L8g1geJxL7O930U3YVmrDCcoleFoamhLMGMGYjoewH76Yct7SJyXDal4rhjUiKfcwhC7
mUXizcrveIFDbwYHGJ/iw2iAdAh0ZxxIZqy9ZMed5fyFNkZ8AHQ2oSxrF0sUU77C1Z67v0YYDbrf
iwQTXgcOGiax+VulKAMKvTIZzmngyTvzxl/qgTrtMC7TVJov/kMXev3fzSeAcZJwyMkZ2m/bGYm+
p30xlYQkDnoriesDXl4fSjy1T1OzhSwaN1N2drCJX7a2u8xd918oRIKCRIdBeLAbhFprO4ab4cvA
tMk0aO3mC8j2l6E25MYrYgcyzqQy/cC4TPMlNYK93o0ZzHWhjzZv6votRfC4Rhd+ehKm5cPR97s3
YQvprCaqj7tYLM0kG5vc2EK88f0DzNZpMo9at3w7JxLpI8UmRzj0bGFiPTNRQ1rZK/MKr892/1hO
BkriXn5BA58yqJb+vZp9+YUX33Bdw5sCXIsm6z4XL54UcHEbzc4j4nXOHciVduaEHP/NKNTK0dsp
8ivqt3DwFXNUk6atWBWdsGl8fC6+6UHdSCJ2rLUwodPw2igh8f2EpKGgGlAvyaZnJ/N0MkPHaeiU
i0X14+mBNZ5atjvWZwLsj3T5wqMKOVg1r+rw5W4O55kemZhDNkVXKKKG4FOst4IJPVhUr6aBUru+
xAN6kVuu+R2qGF23zDU+Gc+vXJKSHRv/tOY6jC6QDMdsPLJw86yobTj6zpmHISXXZ9FCCbR1GJ2M
5LZWCQaNTd4eKoJ6AaMYIIYkBDX8Txh2/4lj+PP2pbB6AQlO4t53+lf51Yo/0pTxCtJR8D16LteY
l7LESA9/UFUgw405KdUskwxVMQVarNanwBq7Xgd/1GAp27ZLFk9ALWu4/dfPLT6x19e1mzx/mu1e
QtnfGcmNrTN4q56pcgOI9YcVEdlorv9sAT5kzXpDUQpigqiytM+TRXaH1zzTmof8/RybWKHVuh7c
17b7lTyoUAiMWVRldQf8EjmzneMsUaCjYrW0IYODBDJe6HQFUeCHH7v8W9yhCRGP5wKrKwk+mSSy
VM2v8ru+ONZFcY+KUYwK7xt3eRCJqyfucaIdH0HBiSOCR/5oQp+8UDDuoftrMqQTIsG5i8nEK8d8
wrPJPTHSSiqar1FnVlazzpFk5xmva0fiue4NQl8mIlUAmwJWEyH0e+DSRRrOZYPeN727QKo1rSXi
2syNaSuiUhZ2vDPwN/HSL7wqSu1bFBpKXxbW2Kp8Ud3kJ+bBilU99w9dvvph3j+Cq6XXIw7mOlDt
wtARtguBlVlizI1rRayPD4Fzs0YvXJMiy1seChknxGjnqKpnYSDpq9u7rGVEcqLunLZIXU9k+Wer
5YZqTkadEltDpzRW5JhdPTPI6QYqyKfZPPiK5Lzcs8mhSgAUeVama3ETJ6iOo/mwVuJVksP/q2Jx
dK8VGbtQB5pwRuHLpG7e3aNH5ci3c3uoMG/LvYzyPIGWVDLScYllrqT5nhMtZ40GLya1gbtqH05l
WHwZn+LPaSiiXFOLC12yl7BTz0lybn+RcGX18jUyumvLwUjpuf/pa/MZVusqgFkGZuSIJveWSx1g
KIOEEEsaSy8tconVYUGwUtMXrMWa7pe/djJDHfUbUQoRk2ipZopbvzordgMx2f/0Nr69VqXPMOw4
nC1n24b0gaIwEa+28H8yrBP7aTIPhxysjh8G3Fgjx36eWTbYjiF1d0FSC/W5S2TtmuALQFsKXKlD
p+du5uu/DwyfyqP8g0W6rbrMWI10NkqdvYWXpX1MzQZ8vlxuHgzSljylVSb8EVNFDOCgzZJcHJfF
ssQiG8kMeK2sANaubFZs/aKxJs70YaD9mHnJNVJ4tNVNW17f8j6b+0XIKEeDiNS+Vl6k50xrUtCE
NPl+tyiU0Wswi/3lTqo45nkkmuWMsnSdDaGLsuQAy1YrU4+4HrqCRyXFq8FTAeG1TFLYdUET7e4L
qJTp5FjR0IaXfvmWBJmaXWUDX2RqYfkhnmBssSRBLIXCglYjKUVcFV914aGY8SJfuc03Py+vm1pe
GohWQ0mYlv64l8GBIhCawJIf1H1taCW3R5T2JT+OPHLXcLXEbKfpDci/dPJ3VAQKKVFP5B72ibNx
rYJAXxo8OrIwm0KDLqrLzTWM/HN8wIQMVOaHryMlKKQtozpZl+N9jC/KL2ao6v5C4fvQnztUqMuk
GTtGJiAz7uEhSHpjo0RjMMsMX+V2nRunuX+kkGQsqavAOWMZvlEj9ZbuEjOhhybVO5oowsYPHiEn
8vFM+O7UKrKk+n8K4HewUr3Hd/tsD/UOqOlznHq3ylVzEhpEFsETdsiMY3qbPLVEevMV7+a3zoc4
HtdTYBPJe86FNcB3B93i+OhKAMCIt3DmG0HNFXSzSBW6ixQbIRNug5pQuStbItOtHNvgxDkiqq1a
cr0pfWIkC0Vf4BFmN4+lzNk7rr7aXsANyE/tXmnY8r3+i+q7KSeBXXQpSEcOFvgl0bH8e3WovUdr
kbDNBETae9lj9TAugX/RT6J6+KPf9Z8k+wbqCXZRSGj6cGgOSjlUe8kn+nXY2ENobxofl97FJZOC
2GwIwFmASRNsa5iLmW6+fMaZecfYegBGrou6fm1di3cKkTF8oNUOzyatk8NRZrMrdZ0gc8VmWtj4
+lEJbYpP2/O33juHRU2zPa1qDVMmlAsQihT2Xc4tydIn+Y6bBH5jKA3iJ3/Fgqb236ZOEtzuQP1d
Y1gdmWfnX3FlmVOVyGglv9KtVPLxQdLnCZRbXi9R0JCUtfu2FrGCi2WaKNLz1WED+tVkooK4H88r
aah9zMniIePsRxnBXfxKrH8c5VLvgfREWI0TxzJNyJW+hb+2gSh5KKyQBNNHdXC1DPZ2sscvhPqV
/VmWtCf+ADO5JKBZPAeQZvNTqXzYTMKTb/KwDwX7VGCeo4gVwvmGwDYHSwKKrYhVvGJypgjjSKO0
7Yky20d48yywQKbb4ILlQdfBI1teAoC5xsCkQDp12ITBE26YOT4Pxvj86j0UoOTX5X1Ztpy2BwuE
LghRkuRX185EKdMvpE5Gp2tyui/utIeAb0DtPHsO7oE3X+vczoocxnA2LLlFW6ZqlnFK5R8YtKwp
ehn1dxYun64sXbNl+YXHWCs99CnmMO0k0ndvwlhFsYQX4Eos4jIfRZpnf8Qg+0ehdofyif0cuSie
IK7Lj0odrdczgthvfbtEzvRpfLfKEzab69XzHjncGz4jQIam5E0gymFIYmAhHK8yVWk1PJ6DY6bd
Zt55bgl6sYkgreqgWL3chz5Tti/Ct9cFP2gnDfBBFvG4twDGPLtFqH0a3CXGk1sIjPUwcgJz0oGI
KUnjEgwpiYWAaVdmflzzEbmD91u8cIvZq1rugwa9AiH8lpSjDEHuytMuiI5G3JUiUJksbNoFs3Th
OOMpssS5EuSrIqQ3vdtQMaq9+A2ScbeHTkt4pqPikK1ppuBInPgIzdc/ug5Cs6zTV+7AJYbmRRzI
Tch4zvQDgKGBGUevx54ORGd5EZTcUC4vzRxTMopCvYcNbBG1PeyfK7Uhc/+GmR+TNYttbBNAInB7
9T0Y2picoOo/iyNChn+WDc0u0AXBBaCgy8uYWQQPNTjJirLm2dNTpzeQnUYPegxlsZE/RXivkFfO
0u+6DjWI4jJIVTOhfoTIgMMR1Tgn5WtqGJcSBL3wH8YBVZzfzFVO1KH7OfdtGZTs2WuV6tmN/4tY
3AS5lcJNiM6n5DNiskfqzXbeF/eR33W2wBzZ938L7ndDymDPKI7WQGP1MFGe6lQBhHb5q/TZa4UU
xeN6niTzGsvXSWrN9L/ngdW57fn9rGDQJSdgnGp8foMqVJ8wuoRwZPUxkzmQ8yf4Q/bw+aWP9hMS
Km6ZXqC8Uqe1E425ugpD6VEPMuWcI+KQ7ZETUJJNievTxaE1RGErtpgSvnsRqoA8E/aKpr5o8OGa
8NUne4fivBkrt23M2GmRMheRflbxV4KWMF994lJFpDz5r3kTmABx/LewFbG9megpwUv9z7oPlbr0
QSx4wJ9I4CXeKUv1Xk8jEdfwU7/ZrMj80efRmev+kPmqPiZv9toSylFy8+wht7pYBozL2tUrp2Rr
s54BFKFKgSsJtAuqhKYW5Kb7iCmiFPX7yvcwFIDIvPK8tBqFE2ufCAY/jb48BwrMIljIDZKQNzGx
+gh2upqKzXNQOTDjlDNZKklAV85DiwTEmtbVcBglKU4nyaSY/k4s0wBf5LOIaheWr3E4DTIU2Swx
kWtfY1FxweEzUD7dk4F9XvGQiQz7ogjz4AaV+TOaAT2O6CzNAxgzfGDyBISPUDu6b8fqRnSmJZ9i
wd/h7c2J3uVaAdPx8/y+WKAMc2lJG2MLn3ThlcGgB8P5/g4304YAsSaW7bEIgxkxQHtCbtWuPwkU
D6e1tFrysuNw5vDmFsyKYWyttDCE6F7DVq2VXw+38tvXBdb/OovSp11ZPorYz9uxd6Y3AHSJtb0s
6SqHy3qaxLVuXzG9QPqyOh6yrFN28vDKBYAhkbIqXf8GvZ4biQsBYhfLh2CmnEvDeRs6atHFtp3w
JhAc0wL6Hv7n14jscUJg4z0Y57Oxkyg5qJF2SNbhV+ILIXX2yVk+mVnZSO75a7fkiB3/UjW0qBHB
Vj9AbxG878ifL4acElMHiK5xnnRWmQhibQ9Id8uZa80WqnvmkZ1UzGMrJqC+dtGbNQ74ZQIs2jTy
vEstp3Rqp9ZZ/K3EvsBetdLixPnxIgLT9sMOK01I61lg+/1vmjwk8bIkyHG+TKQGTdKL2X30Jhpk
7+o5DJinf5VrC/2a7cJAGttynrIomNjaA/OsNvLG2Mowl1/Q7SKe8DPKoSI4BFNrsZt0huJ2FXpt
4YYMaf/VwZbE5Rks2OCmA8c0sLAO+tMEuHvr3sZumAorPZoaZNOVxWppyvoM/xUSeX4HLL+pMSBK
wRKxhIOSHLzIuslFjtNpXDzUAS+dNcJj6UO8Eh5QXQQFiG3a3lWtc7ykXxJ+P1Vp2P5VsXA6XsWa
jh3vdWc9ujRLSayEKdxj0sWGnZnyoWQw33KEdqEMkTtCyASWIp9mTVHzw8bCW25u1BkE7xDm8ma1
rnQQG7ka3x/1nwqqv9/iCfViH4sRKqvKF2iwM1X65WZhqCjE0bpisu9ZQh6i7KTvlh7DQrqDtDyY
Xg1DkheBAUmuZoZrRNyoMKzbZA0nS7gx26jZgq5ywZvuTfqpTz9JEOWbfoJJC4+lUIECQXNz0xXi
CQWzr0Vy5NI1YwcEl1FtemMNYOThxbHRqBH4UPLpQowz9rsKP+w2JjGwAp0WUkZ79mbaxlEvDJiz
x83SmYGuWIx/oD4OHJ5U0bbqyTxp9YC521SjjUHC9+ta/zj1N/4BtM39rQeJh/g+vHM8O6lawtmg
JcuHXOtiybYS9YsPcSG2LA83DH5pHvld6idPY0Qpjbm0jm4WoLtFpXAVtbd5+zbRM1GPsDmT0cRn
saOhhZNtE/ZlkfcbLKgV1XmCbbuBZfycld2hfjyYRnjYe4XZVPbKmiiy+y8qzDam9LBSzTMI2JKG
y/i4w+oE1wkxFj7K/YkvMOSiqIzUCgRh59Ew+WwTj5hPnXBtitLRuJfNSuYd6n7Uu3dpOE3YWAMK
7DpMCceVSolb52MBYluvArmkEVv03gyV539OX28QVJ8i6wTkROiK8dWLOLwMc/2KrWgjaD/YgRrr
u2VyYzO13zgySZW/fZZGJG3Bwn/KP2e3KniGrL8FOzQdBDGRzvaT9iMoCTqaVu/GqibJhhaUji5b
XYXTZLlib5CKjSZ7kuKCGo/9Vl63y3BF3fXHgYtZWiKKqqKnrdvREbNrXy0XuCloTSqs8ocM4JMi
Xt62uMJKp4EPYBMTN7vLDqk6ot3PWpyJwYozn22+eG6oyNSca0A2Z7MOdwiWj5g6s7K8dhCELNRm
9XQfRGLQd6kUcxF81IOJ5LEy0bo3f+2q28zbLeMdN/X6XeqFHW4vz2p6Qq8jO2+6pVZS8Y4XfEl7
cfcwivIk/EaH/FYH3i77qVG/tp4vOV2sFxnnK57tydA/+nwMVJ1JNL8hUMOtRAu92/3BDIW2A7iQ
ciwDtvRUxWaT9guLsaA7O3g7xKrIfM9NbXAiEYW1pHaijeYJHkCaXuY6q0/Kdiw/SrQgHlNoeZcN
+TzzzqEzoL00Xywsp95917VnuQer8jKO4N0TSW6sM2Qh/zoI+LvGtDp5Gwbl45T7S1Q9UzUzYvzD
vtZ+OtGZXwVZzjQc10Qr5LK42sZ1lvopBhO+XmRsmzQvCPfPjAqgzE++NCFXqPsXipVnM/Hvq1mV
h0vXldmY9gWv9/AgN0r0E26leK2me032n83qcGtJ/J1P6ixijIN2LhR2DjjUcjLM+HqScYd57PCB
WNMq8NzNpA/xhitSXbilMfKhU50Ii7YLakR0pWOa2Ol6PGFkIBmtqj74UO06MkMV3nQ2pxPz8yig
Jsq66SVbfR3SjMKu6sY39rOOmMfj3zWR5oiCoy5KBIoBibRt8K2MJ7MSphEZ96+2CSvJOe3Ygg4D
nMDRepGnRAX49DqJ82scyw4UaYcgdqPzib9Bv5SE5M/FfebgujNiaaWurk5aC6LL+so3AIAzMv3K
iOyi8fGNUTQOPn1dqFUYXdSbJQnHc7+ezqKnwfAPpympyJR46prCdjpAaN6Z9GFxL8XYte5EjwRD
rNt6TZmDQD7B9g4bwTsKB2+F9oKk1UyADtK/ptu32MEn0Lc17iR8yQCEq1PJSggOw412N+Egh8Rh
tACZupnK7XGwlqvtpme6RFuLt3qlVHw+6LdgNTA0N+48ooM/OA0RkoYaIGOD1NHDpWaappIBZ+W3
0pqybwv669O++6lvk8S6Rw2/rXUYW6BeLJQ9Z9w0Cqn8cKsFW0LhSQmrGWKVkwGd7fXTqTOYm1ny
RAGA0sQTduGf0UBlMKeXAok4DCk1Fbqt6nqsF2oZKhPvbAYJKI8Y5s54Px7nrRV9kMqqHjHavHQ4
j/sac+4l37aRAW1CviYnDdmxMOpELQYIvBcxwwB3d6eJoQeQhcB+3fuvYfW68yrButMS3fiSjEx1
kiOr/r5HuzMjznyG6tZAxYuIdwggxhH6JMxmHB8+Ng1uY02ac2jIi8OJ5MQRnCm51WLVFGOZz9be
1qrMj2iEEWKN38ayCLB4vpiLHaVm4dmWk1N5E6CGNOLaE+G8uJyT3gPMJJOfg7O3M6CfkcDKdTlZ
nKSVJWCoiMnl79R9rVQr0S3wrM8LR5jIVEAJujierBz8hUnEGD26wpi41UJyKC4kxUlFguzifdEr
mLH0tsV0cvujB/RhOqsUV+5gGO9WKS/Tk12xPjO4AgpZVYJHSo/CKbLQAHfjI5TcfeAJr7i+OhL7
3L04HbIme6DK9Y/wVW8sDIM68/7Gss+S5GRihL4jD+9B/1h7fOLqoLU5CK7DMDrTPz5i2HHkLIdl
7XSjWPToaSE2WkGUSFvm+9BZMZtewZrEIVDFqTy4wgth/Ea14K/RvpefHbWSU5ra/a8LL9t6VN0u
LpVjEO1c3c1dQCXjGY/RuEX6XqyCFgzx6uYnAk3/rVx0VbovZ7R8nFynUQ7xzGr72XkNlmY/rEnL
YyvY8Csye8v7Lj6PdWKOIIse/u/27EP+UvtH3Jip2bfbCi833B3/7cVF6OzWq+tebW1ECU5XVL2r
uQOQANVeQEVQBvpFJR/ZiosapYhv5ZTNqoELXuUpYKt5Gnky0sEcZlZ5XW10pY33qFRHwK3TYJBz
QEqCuUAkTjQH9+ghr6BhyAEob7TTRmMLAU88tZF5x2GD4uGN9oksCd66OhUArWkES1SDb0a8dxM5
meHBfO0qldP8F8ijzvnRT0utwMHzt24YaTMRspIPVZO/JCxy7XY6c+6i7PwgnHyVRU36LmZ2iS0x
1WJpZZ1+XvPJESmE3h7WNUwgEUQrvGAQVsoAnKeLgkiFrNvOlZdDU+JnzZ60p48Ylo+BqwJ6zhbg
VALXMuFgmp99bZUldf62NBgE2PLLB/fA1QafXe/40omdFEM9bN08NtsFTRWLDGzRnCnHhNmWVcMR
hJI7DfGrA/FBwNKZIkGAnj8AnJyLelWw0PqchQ0S4zVHKY62gC6ENH6p+rsLkv/AZVDMSfDyd6Yb
8X8EUs9fBSaMFGdDgnNywruxpceJkHJQdr+MQjh1UG94ruuzgD6b/taQnHc42/vpzFOn68fH99nP
wvgVGyxcwZugeILEjZFgrskuOZRofxuc18gne7ZjE6HagFk10N2hBeyLsL6Jw5srEFyvwjZP9kN3
TrMzveR7gZdz++dvBcPv0dz7ffAgW4yQW/RpeEH974WWxQqPLTY61ZhIA25SX45c0gL/1xcCrCh8
dL1/u0sn67Ko7C6+3ZIewEEqiyPH+vXtfA9c8paRgxuuRX+86fBFhgNOl5oATNps0uLbWmQr+1tv
xHhU+9l74HhdunplC1bwnEqVDqtRDzWXq4vqXT8pY9CVFD0+v13Jq03t0NMKCB0kedx+k02a2JPm
VJV7CqqiGoz+76D27z2F6BXkrwyN3AkzEx5IKu6qwUfPuuJ+lJFvdAcS0V4lPhEIST6N45Yvm7yP
s5g9r044jC44ia56C/hBiJ0di8Exb0p7Z458lbJZ8nIcDYUJUv7Fy80TXMUzFAHO2P8+qp+Kh68F
fWWb9ivZRsC16VegjxYXoR2riirrMjPdrb8M/E2+FG5f1M0f6I44tv//812hrTFgDG3dPAz1LUuN
pJq1acDF2Sm38Q5kExN9FLtrJXzfl/NRSo26BeAvrExCBKHMm6RKxsoNVr84gpJ+RWXhASVYYysp
ErGlKHwygvakTBB/dpYTvR+5rnc6E/A2QDRLeffPIL6AX6w48jMP73/DDxZif/1woiklXeGnTmeh
agmLGOPg5/UedDXcndglygG+sPr8vUL9oNhYoCwITaC2QIqG/gYzXEGpTUySTRBpT+nAju/18yHR
/0XXEK6oCeHs4ZF8cWL6wa1RVhlkEHjt65QzoKNPNKumK3pM6Zpb5ETqRZ8R9e13ur8BOegHNdq8
ZVb1m/D7iuP/KHFUe5c31c9oMBec81ois7i0gf6on0saim/xg6Wkc5RjdFjiLvQan+sNd6vWNKyT
a5JiB3JSGEHnjdPS4uf5AGgH5ewre4ytHCo6CWnzX1ZDX9Wo7uWCe8HzQWT761T8V2w/ksmVViSk
zWNGufHX4dugCol788b9JA0eWZRdPCZe7zg0/57rdz4mhX4UAhPPGHOubNje5TwS+EIyk7W5kNOd
zSu4xV8DIrE85tj3duZ3TC5C+yH584IoyaZ09SEuf96tB3ARlPAKtf89VFpSTVXVfMvBhNiRXA62
7xOguJzklzl+T+8qGfjjioXDeqPCT/uxC2DjzCMfXZ5VI922ClPkzd52GFcKnwmpvvGYwsHaEP5y
BxV7N0OIdV3SMjk7MuP7jSd3s+HRiPbjRVk7C0i6Yeh0TDUqmyR2W8rthBWvX9fWK1Y/fDcCjYLY
om5xm43Lnpi6cEvYgFgiS+jj/cS9a2jKXyviJgKYEgHY62Qh0F1/AnZ8NAXa9NY0y+ktFYZwjWHn
q+et3f1/oSfipA/RKL58Iihinyi8M0zAFzneYk8DbeTF0zt22NT9gBSg8fbE2G/dqnL7FtVklCqw
oNcKsGq/2mtr80bdcjHcpHvEqdgVmlEgsmOz64HukbftzN5VJ1IWs+PHphHx9dHA+8BfrMV7h6LW
REQLVaDZJFFbVhUZx/K+5aL2BrT5R0bfCB7WGAaNfXZ4TtG8TPPXwmynU5JSfHZqfk377momDOML
y/Dl5LvL0PtPm2hc0kBs8OCOhbL2B5ituXUBef6gqnLxjAjhH6LiJTv/I9yFOQsabbC05Pmm+IIl
KlrfJLat/yz/L6EVzy3AG1yS7enIVpg/gwRQipWHHYXGC5jLW0Gfq4hQN/mqngjO9WSiH/DwlfSv
XeBdBJJTP5tGR3ShDJ1vnYIxfzwfEd+FJP95E/QTGVjwalTf6m8voU8tVieRs/8U6clGCCjzkNiB
LWavr0bvNr78RdAIzLtIeMwtulG/4/pZ9Ls6crq7LhXRVZs6VNQQp02Rp/HKS6dtzeKHWgUXHkRb
G/8AEOMa/7OJmGheOvzmWo/+inPCx+4Z0J87aynO4mwnK7PQBS+zabmU74szGdR9VM2+b4D2nKAB
2BjNJtNhD9tN8EPBE7jgwfS5co9kWDt1WOIYXbFuFIMcj/5oKffm9F3C0AMD+RUTZplhERimXVHS
w8jcmEjuE/uTTYlShdneJoKPvZ5GX1NzjroaM0Klj4MoY2sKMKJugA8Ha42gJ6HnsvT46s3oI9Ww
bHujsO/4HEIH5M8fkmF+aDfofXvLGYInu1KpBwDdnJ+reiynEcen0JVDxskOBGqguZmmgUQTnVkK
h9P91+2O1KjtRlvZ5key0LsT5ZIErOCMpd6HbS1eywmnVj6OFMoeItLRXUnfMeeaS5/eHwtrRawA
QhHeiuJmrL6RMXlX5TvSPPVntD6VR/iT0BV0Rr+ALa1d537qYXgpqOmr3PazTmNntopAMMdySMWy
WQrwcu2KrOCp5c0CiQWMe0xga6USQfSnTiUjSX84Ji3UTyPP5F9oEgExNvmZfP/k0+B/kCilNQCr
U6CJa+QJDZCvixLYepsBFoxXIQocPrqOVBiTaQ1DywDNZ1S3xmYReh4DOQMt+ZezHw2eIsluosM6
zru2FyaHGADG2T9A3QLeUjzOr/prB1rAVzDavHEfpg9P5Pd/VchrEVBaoSzxWEsgL0N0c1gnIB8Z
P+EcKDrMEBLqzDrWWbpss8DBXc1zJhCGWOpOYFEEYQz7K+99uvczFx76AWw98TgBfVCLU3QfNSou
RIS8btQ3YwoY8DE662QYvoTtL9b/iqJKrZ43Mhqm+0h2geVnmPYF8Gli/WuuJcFux+/052nRu0Au
fMJ7tYcl70DAxHdytbhy6fU04SKGzq+A1Cz0y3+nvjBm9omwY5AQnifAejTD8ScTLxfxj5wU+CBi
a7P4nUbqQSti5h7uPiLoTsJcVqkfT1FY8jJjqo2nvd38gJUMO8TDaF4p4uziNqYXbdjy24V7RaKo
7h6Q8tm38+J/SEW2iL9+4qVgHXF4fwQMmjfXwp+NgeathsQO8Q/673sr93PQqRSNiDyZve2v2CSF
jZ5phPl3fJRH6VZ9NYjqJusefBgeQEOsp+LoAudvg5uf1QMQ6tLqytemSCwiVCjOpxaOoCcW3aD8
YpddB3rNVv8dywBprEGkYvLKj3cjN5h0LwL9vQp2AD00eAacuh0LEmkHoAYi9FCrcEzRiJoguhP7
OjGkwjYpLxqWuu2DlTimfMV5X9dd9ytObVrS41cm80WXfZJlflsxi1v3JxJOEhRjvvu0loIltA6B
DHmYV29O6bbSBNJY4hDwFh4Kele9WUNfp2TwKGQGMKBRavsWh1rmEYVroIafWCRAxJZ4d5MJPXlp
OnVo6iP9NbyCILkxmv6WqlBz5wGkQK6p5C3NmC4VNDaW+5lNBbRyxbRIffx7nsRUyo0YJ96aDpkl
sMARsaAX6GqYAUymHICFlFtX897ZKAX0s5cmwv4f/7BilOJPz+iuQsTki9fiktaKL/TfKkzhbWv6
4dtI7y0MhOXDcY8m2vYsl86ig4OdtpWIWtP6ZWe2g8rCDWRERWYE+2BPnv7NIaScvEdhlRYVlF8I
QKJtV+V2DJjCVbMSudbNRzOuB8yHCEH57iYoq2h5b4OKAXz2GOEeTwFZmIXbdQPd8V+XVhvYezds
kMMY0nZrfIGtRj8Nt5OqV3ht0onD7eNxd6Y5aiA8+J0rfzbI/C2fGYk5XqDsTjgCydkQGZnWN8Zv
W0l/3MbjG4gwctBCW9S6/RPNIjcr+o0zOvLws+4rhvr6yyjju5lsHbP9Cyy8yQS5cWid9ob4gumI
Sw+9fhizY2YnT9Zx6b5iFX43P2bXeZRI38Yztqf8pv9njr+PMTcsp3SShv5ZhnIjg5OvWBnKu1Ln
STQ5OXUSO6VGiPYDPbjSFkVOX+weF8QuLxiLweVIvlC82I6DbLGWpquVlLQUCuaBxTY6cypVs0hz
6BzPQZY2hHa/RmpYc/2bt3PkCiQgn8pKxYWIViQT6bV81IcyfV1OH7ABfqFfsAJBZfR0X8jeCXYT
cJ2avoWxNTO2R6rP8C0mcXiEwBvmU62zdyfYeI9yhJV8eUS+Jm/fOQbueUsa7kruNNc1mIocZBmH
uI8/xXIZNLXuDGHJkMigR/CzXRHLJbNn6wrFGK42/Pc4Un+GADthCsvbvvjPVtmyomppW1gPBkqm
zrDeKHTxQMWQss0Qxzs+DVMabWTruj+7A+ARCPFafrVfBv6KbxdBfYmMC/HDYoj8nwilRgOVPSix
Z3BD9cbRohcJ/H458uC/KQ/aFV2Sg6N6WEHQKrRtjXcOD+f54ZtNlqy96vDitYMw+terb5LBmorZ
XHLu0o7N/ykAfFhiYoe6V+I0bp6YbsKT+HjNaMVUBx6GE/4/lRbFTD7fjWHZzvA39WpDcTREC/Y8
hJdHD600SWUa683bq0s81z551dMhRixZyxEIQdRwqZviq9wuO2sqO55jetaLADQCTjaW9D+YS7y5
5po17yNaoPBDb4GwXaaYaVqrwcTye+Eva34zYYJjqM7EmxEalrTlsVohr2pEgffe2pfP0MZq2Sen
UD8B1fLeNUUjkQhgMuQh+T7XKyud+mls0D+7EDJEXGEKBo3SP93WQWmbzdHxcXtTpy/6t9bebLK7
SySiksnhaIav6mB1dX7CL+xHlisjjVWXC1jR7hVdak0y/pLa+LVSKYu0ns7Qhy2bh5c6ZI2h0/xk
1Vtw/+3rVZlEXkSa2CpP9y27W8oM+KaFKZjbq237mnLkh7gZ7zbusUp+gB5q2sQBFZtF/fSkUM90
wrYtXtIjyNUfWP6kHKtzzq2V7/twoeWqpT2Pp95IWPzT/uRwAMjN3VkYkMslOoJMseygWYFbrYJ/
rhh41F/aedoEGlp0jQRx6E6If3fYruIXbZk1RumRJZRIgufJe2xKJ0T6CnGVTrctIm5iIu0kc0aQ
ephMIm0HHditog1yrCwXWOumvKyInj5xu77RON3ZS+5aR6oHs9Bue2zYtESsKVmAHe5NGWlVpucm
OeoJEYHDn9Je0V1wKGvZUvkyzYAuTRsEe9xJNJgDcgu1lC4RstJEHFRilDOhMWpfX0/spnaz1fxr
M+zu41f+3OgqdFLPUyAODrR3KFoJr4h2Ap0t6dNwhX0NNJOH5qWChMypCwV2wo30bLN4Q+KgZdQq
d2uqC03fAECxvvQ8QDzc/EHMIJhP17+Ojcvnqf3vyA/jZTcnkPRiQwb1QxJA6O2mEwW+VNxWbKJh
6IiIEszHl7CusZ7WIXkD12BNmeqzYAEYafq+WYv+V6bLPZy22hP59eXBCJFlhVyTgKYAVwHMRLw2
iU5ahk0aSBaXTwrEwYX8vpzRH4xqbZ1oeJl031pp3Ui0+vo0HffySV50oToC00aqLlKqFU7pzDdK
iC2qdtiIj/eUoiZRI5c5vaxd0avoWG80uO+xxsmbNFeM1pvXlXbsN5aoBQsHOAKjpWTGLKsyaleu
fLtBAU2HI9gGJFskVg7Z6BdzzhB5QiFAte12jQ5N6kMYK4rvx/6KM03VGrkrn1vPRSw2uZxFbcjy
CsfcYotWDSLvProggQthbSJBdOSqk8oKZd0LpZlf//qRgU34JkpnWV2TQECx7Zi8HoMiWS46toSo
l37YmOYAdCPSRduWAjT+RAbGqd1UJyZbwybOgDmy+8J62v+DHoQfTVw1+fUgEgZFsMZpe47QYw5r
71PgI3Qb6GI3coBZFYw/OE3BTd8iT9+sxokbFOkJbuPgCg8YMu/uKj7YekEF0yaHzsqoSwux9Nz1
t1eaVopKZ5JKDkatMbwybZBBLOXbiFKLNehGoOOjm3Ojj2mV5nlxBaZbP4ZJq8HDU1MqHS4Yt1+N
Xll7G9RyLuw7zPhb31GNFSaLGbw9LN8CQyJ/IKlibNPIwWFqXaMpU5GBGrh4aVm+LFTqwE20edsV
SocJM3T7Gm2wdd8TKy4hzJhF9sP7ohqKChGz1ug2f+Lo+CVSBto/+U1DvCPshmzHomf+07LoVBgZ
gtxe1ydVbNT8KkG4WI8/QaPqHzK3xCgUqiNAtxKElOvfPdGHFX1vydra1d/x6Tw2UaBAHSuyY0Ak
uQ2/YKnv77jbhwL188drevVuyfs6Iy7z20I/iDL/lED24YbropzrhiDBF8JEpmWyl2AjXGXQ/2ej
L1YB3yWMWRALvbD1F6bkzM+e91MLBm+WjeeuvpSZU6gI5WDMXXLTxBIAbsHAJ0MPaDFiJtJhxpsp
6IySY0Fl8QXbBK4rwjTQhRmzHUONAGaEY4fkPtexrCVlZmOCODInT7JI5MOwTYsca0asyovBbrXl
3oSarh/gUPaBleVN0uJF5aRk+jn0n0el/7a2+XP0Lp9z4iCMFOpYCbibk069FSL07NRHUHnzneDk
q2BZ1Sq+PYBMNOdrlMw/pPmpZjVL4deq+xFhGoHpWXKO04P16091oAFewGWKaNNaYHNBqKPUZTEB
1zFg/WK6hfXD7V7Snwy2AzGYHLlJ54iijacXicWVEVl3oldErFw8KQeS3ck=
`pragma protect end_protected
