// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:44 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
JoquZONtc3qDzw04Qb+2oleMN1KcJ3wfVNndYScmsGKMjVkcsDzX82907uGq2uwn
Wpoa2c0MWVzoBjygLurHM9/Nn4Rtx1bukXUBnli0VJ6BaYk0PcSKaEg0lI5NvPvi
qLK2Iwb2wmqg0H1phMK8R9ooZMIbR1h1k8qkorWpNOs=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 2848)
z8lkqRPl5X7F7wq8tLnlAOe4Bf6qpr0g+MVRANLjI+MBbAP6oiaxZDgZTBotA4O1
6vE8zBpWbnR77/OmOY4q4F4jEa/ND8zujOa+/dNI/a1zIeql3HEUDrHOsLa6h6YE
XaWhlX5U69hr5BzEH38g1WR6XgO3ZaC3Y8tkqk+Vns7gfLqRjL00suQ+hH470jWm
PuZdnxdEnFVX7UR3bU7BUFrU6sxGE9GEs1Y5MTpZvx0N5HGiLGwTrhwOaCvmEgbC
5C6lHsjYY/WFzch1JTwsb+yHCGOyeWIGXUbsJ0Jbyk+xCpCWjvFEzHnJtbLe9/lA
yLMXxRG01qRc3GMqG2tEnrN2/ACAlW0fyHX0wdhXjJSVbgsMNAp9CQs5wkJueHSY
AcWTR8U7SQS8tJ7nid15NL8QQSQJpnz82IB76lMp+b+XvxPM4GD7VIV5FOkEpj/N
r5OgfvPhJHKsBtFlVEGKAdTrE65FCzattvcgiebFJyF5ytT31aGeyt3lPyBpgzi+
Jy60BwrsfFt7m+ejswbpACB9qApqBbWzUz2WT5knGde1Q0DGxjUaGDdspR0tZKgW
dI+/BmZ2ptV+F6LgUG29nAMA4XCkuIIAI+tTY6saJBzDhaBdypwRd+SkQ2rqclU4
VkJx78mAgzWsMT9Mx2M91fCnpmEtuo33B9Es8bHp5pSqURksSeYdB/MYQQP2Fc0T
wGE8p9yGEK3S190bUO3gcmAzRq4MKMtXH499HCrIKUkg2gzXXQPwWFBDi9JSBeVu
rPGgJM7lnc/rnSocGPFqXmYD/LPcsOMnjZ7NYgonl+n/oVRlxEh6RDpGKg3fEn73
lQB/7AtbXMrZB+99W6n0kwpyQ7YeFOlVAu4ljpCd5p/0My9zlav336dLktN/iKjM
cDQ3HrS+7IHiZJ1zkpTI2kgl2IIq+Pj4KVCf7apyuftRM8tv9JGxKzdj8V/ahkKW
KnPA1qnicvVKQLgbXhnCR8/JourWWUkPltwOYoy+4EAeltxtwpVRv4/iPKpxOPbO
lvNBJyQo89uFFFplJJFdMVM3b0jNh5YiIHzPic4pYbLyjHQaNm/YqmIcUZzjq17f
qHVj3vESpEmAU6n3D0OJE+LmViGVUQmFjT9L9T7Ef5kiT9XB3NVsJBkb4mk6fNY6
IxPDsWgoqNLfYeLjeZgK/2gJe8LcONjAYDriin8g7P02GCEQx3h6WnzFUFzHKGAF
J41UfiaJyFHRiRJzCwt9X1CrjNIF6pwsM6xoVBXlDlbsLq/Xs2BM2tiRXmDm8ODn
ECeieRjvGvTon0x/txn7Fx10N1pwXQcAgowRNqGGhp5Il2E3Q8hweXdtVhfP674X
RlwiErX0rR0swT+iMdikIq7I7+nqxzgKonHKC+XbTqWIMYsfyKr2R9CBbWXLP2CX
r04o0XaXggOddTVDzpiVJtJpIollZ2kGvaT7Q27Jw5iSYTzmS25v8OJtjkXyWxmo
dTSfFAPwJrBatEZ+1c+3zFzSo+hZGOnLJcyLdXt9s1Pg/Bsx/zkzQwc8xqjXT09X
d9t7j1wsgQQOK/RHzLIfsDZKXGGiXz1KrBmKtnJ77/1APVGtdWH2QRwfc558MXvT
o214zWitIIxvSF/3aVyHV/guckwU9Jjtd6DEWdFLe9JW73E02U48cK6z5wh/3D2Y
obmgUDwlmzx1jrbdJkqfjtOb97GGoxwCGnuE8REWJ6HPs0msxsjRgzqeMlkriUsM
Whj5SKM5X4eno+Z9TwsIDtTsYVSBwlfCG8MN2kUoE/DnAoP9l65zJPkQ1Ir5Lvd5
ADkkplqJnjNuyhjTK0jwXbRGDD3eJOxuRQURPxP4H/8gGlmGpmF1B0OFJrCTVnCT
VsbRelm5Hu+2/Hukx07RVrJ+0IOACnaBBytGj2VSy3ja7DvfSXkQoKCzmcvTNAwO
H2yl0hd6UYziChF+4Xnq98FNlb/mNh7KOCWPVnP1ZqTye68Iy2znr8ytqQ9ModAW
wxCbJtcG79J5YPJloS+1kXooMWHPAqmGNwQYDzuRsiY6M5WjRzBZztSiI46O7HZZ
Anx49cYaABLzkLwvforkppdjTAsUr1bF1WS0DPqBQpaqj4hzQpmv0G6pxfruX17y
epZovoPhEXIERLvnuKKKdtOZ7tphgucTf4S2WQY4b5FH9lBH7xYqACAUYsWa8cx2
+Ec6hXpKFyNpDnSVaXJ7bOBWwCmGy5d+AWJf7nVe+7d7X9nGaJ88LOjDBN4/b8Rs
A3AD8rL5EUTRVkrg/CGA/lyZubEoHrbi9XqG4NQJ/xIwD/camoPl6lF2+aUAls5i
bpysUJOWkZximB6nx4Gj2DhW3tZxmCH7aMPiUtEaoNqaxmJup+V6FesjkpQEE0B7
wB0SzbAyFn7br5vnD1+1bACjWv/o1WSAbA1cRuSMvjFEec5M2Dn1pyBdoUk7ue/M
RKq0cEfXpEdsaNG3W2gCvIlnWFiaGNP2kYXFO+repU+EhWkXhIDXmbRcVl+Pp6dk
LhJfj3Xc0Aob4okWON1B/ceKupxS3jtrlZfyE1mVBLkzgLvw/8y59q3BYo+/IV9v
KH5JDqjgM6pKP7e3cL8aRwOAVuaMnpcJfan7yKIxiZi3DfQXapOw8GuoBzEoJik6
nqa9GcOKUWElbEHS2jAaCtcIyJoiC0R0qHT4L0Ze9VkfvxWkP3MKydb/faF2jKaA
XfZdDm5ymyBW22iupvr/B1CiR0G0yhZX8e7X+uZHjvtAs6wd+2us/xPNto98O8Ep
HYzDGLe+HO28GPR4vVUQ+AEujZ3EYdfZtPg88ncf6ON/Je1NyJcuIz5ZR2Rw9YXl
TMFmQLkItelKpmdyRtOwVOwVXE4uCsevcKSOrJa2GUJvkajNhL4jyYDP0fpQjkIu
1PlKA3B2tDONNMFQTHK2/keIqmZUTHQ7RzNQ23T65gd68hXNjwZGYZtNk9sqaclc
c6uyp45BV1GI/MZa5TmA0VbQEQhWwlhC5UiyVgA8b5djTbyBtcBeQen2P9d3wvXq
b6x44eAN31cxotJh7BhpEWjgpYyS/bLwjRmle73sTa6nFhfqavUcAC1iLwQhuAPb
3UtLJcpOYm97fn9mA0Vfhljwjea9ssYdz/iraV3P/tjySdcaCFlBiHJiX5V+6YAN
3KZ4myKIkRVwpFecbpabJ02JO9cBZsQoHKmrlhbCvRvqKiQd9AHXR/EruzPRbSuz
piA4tFm2yHPOZgIcZS68XtgWoLLNX+6ez73xZKKSTSP08FO2yYHWtDM8Jf9QvPI8
w216Vo5bb+6IjqNxJK19bhAj4DYc/xMRxsk7HT/OQEVaVd4mIBPRnh4yfgcK362L
L4dH+SAsl1j2f9+O9FnxKV4IrL1B3JnYmFjJ4KuEyWkEuPlMtCuUC4zNYZtJy+Wh
0nVQA17PJT8ITA2b57EIbguUiy54B6ZXX2vB8+1CMI00Yiny7GZbAImqX4eGPNG9
k+gUu6LhoH/wE+QjpgXiHhfFt0WBwBYXDgKN0lsxxIukExZRMMLSKcaZG70TkuiO
CVra/IarsLc0P17fOx6o5qSxIpzaEyh4Ne1RBOAD/RTqvlMqaSk2v6Yyp0m+LiqY
GEyol0olPfLm5cSmgdb8zmfd+GzBhhQW2TB9zep38VRRc9O6nbXr3P1SWJgbYoRC
ublp5CbvvJD6SXSos51ix6NotkvKeUWh5IXHaUBQMXhDwx86TVhkSCEmDA17gvxq
2IUTyPYl1sjwFoXyvkduCjhLp2pB7pRnHsxlEeqiZVOjBPg/klF76MGBn1nzB7+5
9pBekbCy8Zx5xyWPLnzoUA==
`pragma protect end_protected
