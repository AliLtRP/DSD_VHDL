// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
NF/lQmL0MZMYxrPBsW3KhK8WgfVx5dX29lrSMAo+Ir6afq0G495ANrcF3LinQdmE6lXnodVB8JdP
Lfcr1/bfa702rb7JHRBGh5nDrkap6WmaQHL9174i40UAUFCB1/MlKekTNq/1EzDXWuegBB5S7SBM
cxXPLmYX9CdHd0huykVyAynQxR++fs/c+8+PIjHNiqs7/prNYaXF+HjyMQp1qNUZzKKpQMLYNQ29
7qjLBU+8UJUcgVJYzXC/uAgggabpp8ehNAHAC6jy27f+BtexJj40/xRJZoD2gBQmJ3IC6uRpdl7t
mQlFWSj+G8xCAwwBs84cOvP0eHTbprEefVWL5g==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
Hpo5Ck3nGph5EOYE4xBEMJs2OfIY4vP59gCbtgmQTAnei82RI5OGN+Gqi/kotofbEZ2owsOW5yft
jRxqxUsWOIl2pSYatXEcjja32Y4AfzQyZohPxvrh9xMOESGuG1ztW8VeTOrAA3tbGa4Fv2E/6X7z
boMtD8IWP/stKKPyYIJlVKcaM29fG8/hVR0nA3ScvrJNOTIxUaxZFs9bviBA5Rz02nipnoWPugxW
XWRc8cx9JCfCo7AWz4x6MWq1RUha5GAo6kL6pSO7c8WlrYpwuwnd4YBBxixJKQJJpvUpmcY4dBiR
sCfMjjFd4MuHgNcUi0/XrGMm1OCokvOD1yc1QPk0kUoTQAKWAke5UhDKIhPdcI352UeDfurkZ/Yu
Ac1dxaCd0GRreupkpNLPig8KbcvvLsCSS9Ln0pY75spMVTkkI/upd1oPQSCn4+e0sUQtVvhMtDcc
4SgerDYJCzHELjX9GAXEBk71d5hJl8KoEBcNQjoh5fPW09jVsfbjTxPK01CAbCOHVzrkOo8SMomH
IoC1UzXinyUrC6V/GOf4Zs3uumfkMEyMGnivIp2+YV6q2eQZOmu9kdzJP7QlSBIVe6hUrWU1jVDl
LUpWmqULlILRrEK55rPlzYONFa9TiEXyd5TEjIwnCScpHSEXmQychUK+eq1NPv6SpgBPVlMPL5hD
966BDN1ErUgWOiXhi0ZugdeUzZOEwuuh6idr5fcZfKs4Vdgvkj5adsrUxfvwAWu1YmvX7PyO+JHS
MDbbK/46ucDrfS8DAOCayHNNIC8Rm89iwMwBXYydT+VrkDVQ8uWh2eqPfU9G8vXxc/quU0hKWzQ/
CKJiX4lWF5GXuL7uJZZdTzHhqx4qXb307ygyA8B+pDzYPKunzhDQGQSEzWDOVoIRiXq2dnP3V/So
bwSYWcdZLi/75A8gTW0BKjhjw/4HMzomH6ejCSF8hVKYT0I628Z96tnj8KHCzfB/rMTZaXziIifE
SdJQRjETouDOt3hKEbf14nvRo2KMF4vAPZGm+f63OANKaRMklcSfMrCF5hQhOkj7VFUR80/vJ+hD
uYsk0L80QI0GJRiw4P3ESdlk+qyjdvkXEkfic/TlanKvWJ9aCtzDGS1R2pbsJCU4zb1XYje7WRVb
6M2kdjQo3u6O5CKDPpr203awSbIU25684f99YZDaO0yIrIeV7EbrMbs5Ml3VfyA66Wh31NfdZtir
vwMkaKQXXU/pfB69gXg6kIZGE8KrvDKsomXMuIhsH1q6nCegUddf1XbN2FVoRvSpn+CbxLLoQmOP
iyYrtvjaWvYz95Bo3VlgIBH3BcNgr7jUv/oLv9QvegKB66IQqz1TL/X/SImPR7B9fsEAs7HmwdUE
uTdh0Z2nJ5tIF9qTN12eHf7ppJhIEtLbh77A2x8EGOX0u5OjciTtViYCTtELbG8GHHxSoaI05Uq5
VDcU/TINqDslPPQb5JFJKKyWtALRIpjt4wTs33pU8mv22mKQAHQmbk9Fs2lYxp0X+TjXNCdaqZC9
Y1UOfa3g1uUrr1h7px8BDzFJJQvPtmHA5DeMFmiF15VnPW8Ux943dcuPuZg+emHpGkr+tOCYG7rf
QqwEbVRZyD0ITGBva0VmYJ6NCGdSgQvzDcEicuNAZiE+KcD8FaNbvOVs0H87lVzmq2rEGHqIDWbx
nNjg1w37uGCBW0bvQ8KkN5GtgnjGLavFZM6KoV2SMBC3WtfliPerHsyvR8+n0nyHfVlIPRbYgP9r
c66qp+maBHF4N6ZYHMOGnS/y7XW6S+vz6MdGU2ikx25WO+xpqVt4BGwsUYYbBUKIG+Fo1AYO8623
1ThLlzcMafFScmidEl5sqXH5uO5CZ+zc8AaKewnn/tS1wsksmqjHa1JneYtsIQp1FiDGI4leE2UG
IBzJhSEuSdfjs821JzajMezgrH2mQHg/uONIRqoDDYcZH/yPoPeO46pvrcDXi1UjtlqoHye0Gh4C
59wmxUmi9/SS7kEAFpexL6/bVA4gvcIr60KY2TOqxvXw6kCSDSt7QGpKpLRnyUp0pL9lVed06C31
GArPRDi2Efm0ZgbRxODXaPCL9FBTIEcIR/LD9WRpUDXFJdQG9woXRqSsb5zQ2JmHnfNis4FbLmpt
fABL7jq4lQ88v+Rn6zBINC3KYvN+xrfT/+uj2PdocOLDr59S2duFjUbfwBLwMqPw50ScBv87Gvpp
TrcydgC8PURrCLf0yCkbiJHIk1svj3Knsth5Pjwu0h4iu3ShGP8uilP6x3tDJACiSIJf1VO/Z4Ll
lSOpAIRIZ9ZjMxO7Dgh6I7IJmhUypete52sUm+wWUqnQMGJt0YzpbBEaZ1nPrgzbrZN2c06iZY71
fTR96Fn7FQodN6qdVtYfBZW4jUyLeYOWjVPaWg2FrldTb+JUqA8KNxW/DwQqpShuKASwG+0sAQW/
wgixkM9PhDmFmCeO9BvF4Op/Q7HUZLmH9VTj2R2Ki4TDxjNsofcKcQfqDR+RtAC8GIUwhomyRsxG
xZ6Ud0udO+aD/jHB3fbBiPTjJ6I5Z7169iqhPeuendRVKKH4KW2/2uw+xTN6KaQmzzmkn85j20tQ
wUrf9NYxgJkBWc6uX/XK/HMOTubQrrafosYe9oS8mSuVu2TTm8vRryvvDR58HPrBh/gwFxG8GkLH
zFTifZIAEa0oThWc1JpRysfUKHuOgtHj/wCz6th4hDpuwJwNtPw69txrOEaUjFHz6afpPg8pH5SX
LH9gbzkoN86zWEfEUkhdeci5pdv9XcQaOeP7TbQvKLXJGnNPLlbSBfAtSY6GvzphLqGEgJUOLD4e
m7CtfNvXIQG/GF2jih5h/74HKcmiofpDtm02wJIFVFtgqx4He/JZZBz5sFf3XlNcyNYZ6sELbArY
v40hTy1QUV0aTneYmNUtQuJPD3iRRPVzSZCdETJM1ZKRGiBJjNDXe0IPuGf0ySZtmbnGboovx0b7
s3vzS37dN8SNZcrPOg4RleYNaE95mZ6iOyJzde/jGVqh/4ZepyY9wJ3H5pzev2i44wsmCfqGyGPj
JimxIW65UBQBOwSYrJc5dWgSAeW1XOVMuziv8auKcep6JDp6l6XwYMbukF0W3BJ+wkHMDnYpF35t
1bHdNudnxzgoctgF1yVKeyYf8mQk18fuLmn9VFh/CRIIpZEa9hQNmqYhIoXFutYHddKwzv72KFJ7
AmvzXUdrLgotKN6lMtSKleOWH9XMFU9bXmsKIpJRoDSzmV/R8sPv9I/vBvYzq4rz/fUqvpwsRKW0
7mJeYQGvJJalAyExabJeir20I/inFytvb2w553E2imbeyHoKLPda45llxVnJZ2sYHhd26/MqpjzN
vLzQ0KYaSFNNiBBOQuwvn9aJxEVZnshReFvbD6QUdvvodHJFfArM2DHEfYMC0EX7XZLgaNBksW38
FjnfKHZ29oZEXv1T52QLhlxk9yYD88gGKNlB+2SCov96dLCXUjoElbhKrwbSeHlt6rSHRuKPGVDN
Yxs/CfQvzRMZ3fH3mwBpaUB6mGetSTKO81Q5OOAzC+HfgJ6ij075BA6voOXFkbGR7Weh+eSi3dPW
9mhC1ztHrBGQGvJIw9RxtLWmvd/FEDKUiN4I82t6GljcgOAd/KLf16FOFt7G2wff3mptCng1paTl
NKAQpZ7OUOoEfPFhU5yuGEOn89YiiqEWsoqQmtOCA5+XinrxYJDbcWCS6D6fXjKKY7dwyvqXl/rh
gk43IJNOTH9JPbKhwIaXvCOkizS3sVnWfy/eRy9pvWQMIwPLIq96Gio83KEui0yfoIac1qdinVFv
LcdpbSZUV0SjQAw0lYYEp/tfjLdSALCr6Z+LJqbz/3MzkwXepbZTzNQl288l5oRMXnCch2af1PkT
Q3NdtLkJORhc48Wqd65r5Rzw6iwiF1+6xvJzh+1Q9iAuHPOaYrSQs1fo7SBOj/gLR+JGEZzFb3eV
SqQcZlg72j/IHGAiUn+SWlcpFH4CwE0XMQqE4g5I5ugFyJ9DSTx2i4FjzTruJZFy0G422FmTFdyA
RTCZ7KPq4YSWzEyEpUdI90WEruGYU1NYrW9OzDQMuOR6in1CuPREb38KhELpPOBByg2+6g7mHTrO
ycT6EvjV+7beaeutQnoBPJ4rJvTWel/nr2lAzFE1SDBlgTBUReS1FMMjnLW4rG37LpRXiUMdhSqd
5+1kEy3VVNUgdZv+5UBz6vwo6Q5QopstMOKt4D8rOsYQ2FgA+YHEM4b6hV4QXIPRzBQDrc0MwSt2
U+Imz1cWnXMFq77uazzm7ZLq0AJ95Yk7DNWI308Pqeaa47EYwQXfucMOh3+TbPEXZL/R8iusUuIJ
pzuAUfrWdz+H+Fm+Jx6BnxuhQCdUb9NVJLj3TshN9jsz7OuBE2EHg5d+3UNctRcrvkgBnQMjlAKC
kPrhQ+VJje4AaONst0UuMrNyJ6H31YnxElbnF68IGHj0HENtg/VcKH1Uam7f7vBakz9di93woNak
LKjb5OrcDQKanAHhMR4NF/p2VcWGae1YSDoC259x404wNGpwaj4BRpvc68gKtLG3LoGaS+SDi3Op
9UXKaRWKMcCF57bl7TP3k5vARg2JAFgiYFs8RsRpXmXoDIEFISuseCGabpIEemMmKbXB4NEOBECq
yUe42jWxHedIL23igyeQ75P5c+lPooWJCTNqSQO/1MSlriMC36BeS437TykCFn/gjJOMvLIT9mqv
YUKSzq3TiSUtmhMb5mdmaPgUOYd7vCIvV/bIwRP2wGnbr8yVxMpU3zuDNs/CkPw7rXZrbOddN0bi
K6e+fuN4pKVN1gyKbh2spj7kntJn//8+xP+/1qbncB5INfwP176s5Q/QtHlj5gGcxM8mVBPCQGbu
cK3E3IqK1TXNBpG/lGBbZIFMhixRs5gRJH5BDZO/4cgIXUugedK7nzqdq5A/BS1AMXzZ1m8vMWjE
m4t6jejDB8aEIXBVpGzG5iffvcltgJYE8V9Hj1DGNL7GorBltbYaJwpjoqfKAAAoLmzK0TViH1CI
gtGk0emLabfD+zpONu5wBFF9WiqySVjxBaoK594NY8rmsHr0esbpUrEuszG4KVZYfbrbq0yTjQPi
Oj3Lh3jIzePx/AlWjoIVO9V1i3WgKwpLc29B4bU1uaenlwU/xzBiUZTQp9pMx1iG6QjjbzfoGBxo
NAb/H0gn46MoGDrVh1j1Q0uIcwf95bFdxcUE2LusuP9w/bw1W+OEiis0JnMOGdAFyibm3jDgic3I
rve3wPCyOxh6mf8LbCda1EpOwO7lDCbmBGidgzJDpjfFe9IENhTZQHPWr+ONbDSuUOURaWrgd3Vi
ywWTHlZ8krTyvA1/Br4XC5/R7r1EoVLirKYGJRtWAI8suIfoPEGDl+eeL9G7RO2yWJvFaHLYkETn
fLQOjuqssrQV6zb8GWj45hEYfDsimr5mQlqR/znDmjJEXkh9jvVIzEPdtPXqQmivRY9Raffc7B8Y
wf19m9u+YD1yDlipYoy1vhRDE3OMEzxpdxGgR48KL2vsLhvekzmn/zjCs7GgH/JzE08QRF0kqlJK
ndJiOs7DmDlUU7lhpLBWW/XnQfOMIoFQwuTuShtCQ7QH5+Mhph2546qKsn/4NCicc5WjShQVTfDS
MzoQIfPwCurYqJTAYT+Dj24VOBbRFATyZ4ob4alProCqNlxhxWgosC9KvSwC5H819Kd+ZL0bU9qc
SE6wW7ZPGmdO5OqAKkXXH+/z++eLwg2S8Y6EHL8yXzvuXXqArGJo7gAwcs3lX9w4Cw9GddRf0JPF
5IZ8wzHAN3LUbw8lYGtA0KiBVXe3YzUlqZAcaOG0PqCuw1PeJ/+pKlkEgMQv+MwoEr0y0nmWwEDA
VJ8I0+3KzUmqPmz+W3beS10w4c0U63vXRyp2QUas5qsfTZzZX9I9hPIhF/dfkhmxTRjX+CbTsf7L
UOguzLqn/DQRExE+Pgvij1LmE5DXLOgHd94K6ATU77ppHlzbqSZ4jfdjsIRXXaRcIR6df2YAzMv+
f2y+m/OZSIdeytv0lAl3Q175Cr2YPa5pfs1NXUDfy09P6duCdlPl9tvUx07q3M6xr56vPmTjuVJy
uZtCLeuFOcLoe21GaD+kRzGuk6925rp0Pp0w0ZpJn4vZjNco7jsyFY+1bCZ9NE8s/UM3EXUjmXYm
kv/PR3j3zymWCiuWJMMZq5dK7VMd5JQqyfDMZrXsyqggi7vVaS1Y+zO5AoFlYYhUUw/aH0TfY2EO
mVo73PkB6Qwd93+KkJYyqo+MZopeAXaj9eJ3vOTuohBSCyNAGZgni6xR7veh8Nxi/Ap5hFi412jN
DsyE2gc1F8Wp1rPpDiAwx1GtKFMKlcPE5N2S6yYF3mVZxNxms6JnL2o2DyWSsYGbnKoVyyohJGuf
2MQelqeRpaNBeGIz4crtpEaFpGsHqNYLYPAwdwMkJyJUjNyNeQ+fd9QFVpYeHM5NUPbWr8rEepwS
s1ZuQwhX5zlYlojjVvFvlTjNo7M20hpEaalhv7dkvCGaHbP8EGs9XkdiLjpERwcCtxeeJjB8vJyy
8Mtla+nkpmtiWUsoHtxs9g3HDDHxj3+3vg12Ntkvx4pzi2US5PlKimmQNvanl3ykBjRBQqu5+QaY
vOP5m/3EkcfOAy4aYyO+N4XJHlMoe9kLZSYQejwKXoURbYDXfppWv2hALTfRaxYktN8ZLGuKaghS
fb9R9KNWU20hsOLMOX0YOulVCjfAVkStDvLKK0RVjZ/HdJa06LCZT9ax5potDE4ypVhoJm7rRib1
XMZY+ag9+l5APrc0YYqqgaG8bt6ZDmveitTfcxqsQFkI9mybKv220yCNHnyomyqUoSN+2uKlq5ac
z8zkWmXAovK0Q4qF7BZFqSNOi0WI68zD8P4wNs+ibJeVTRajwUFC+K55NWg9g6O/jUMO341exiaA
GvxgT4GJ7eh+BEeXIxUFHW6d9f3pHW7xrKUTRjYf2FN+/I/YYHPyN+K+iucTteTbCq+MAxcHHn6z
5GsFnFJlHP+xlewl8+BKBwU+s7xcJg75WBQyIvx/B3qO0uk/7Ftkf2ovF1Of13v/wM/FMNQ2g5Ou
z2USxNc1TosggjEZLuOzXrOqWZYfKGQmRzHX2f+w0RFsKlxrCSz3QRdioiYLkFyGm08cVnSB7iWk
3nONzactok9XKwMKJc0GPcgTzwDZiWTI/ukKMTJCC4XdMq9ni5aDfmICcP+j/ldD0OmWbOdav5sr
OHYfnAL795hI1+X77a1cdFwUb+jNCnTg1Q06Lls6xCVdiOfl/U6bkfnmzrfuE109Ky9xQhqtJQ7d
RXwYxNi3NYYYApEAA1TOb4BeBVOr0OaReoTrzb3pvdwxPO0rW/zR99esMIJNe8BU01g6qGgTpJ40
irfEN4BCM+4ep4QXGbNNfhnSICMv/55usc5zmMkU1UOMfXoz4n4IAHLif4h6RGtEKTMoZRsuclOj
ILq0KfoxD7fgZBG/L05WBfr17TCCKlIZmLBErFtdD75tS3i+/LwJlGLsBjPikayvK0kOVGfZS9ce
QcSLJCaffgYqFRoinqnFanr6xzkCBnrFG/w5q+i2eISFPoenECn2lcum+EM9d3XVnMA1vXJtP7AV
KEp3TBRTzMr0vRpUOCV+GshJoTD98Zh/wWeUf2gOJFdFXUIeyWShWBuLzZf0VVt9qfilsh5Ccur7
mBOtJYX/5/p14FBXdzL7Ru7aJzRu9UaFp1Yg/as1IvqMlSSwKhGH0OdV8ZG7XTsAOCc4LA+W8F0Y
/Vi/Kbu4Tv9o59OrZkAK5JVFdkbFuD6JiKzq9Ozz5ljwxA9uCX0sLpw76flsRdL9xIKo0PZY3AKX
acCAXLI5tQ9dX9E3g65P6qb8tB7QA9QfEQ2C7uLVK/WSk3nzTuEJ+8b5PKaDgCzV+pekWWJHWi4S
WyKqeWq9xhySaU6PgM8reSP9uOx1bMy1VL1dZDRxmvSqWGYPE/YiHIzZarkudJ1wvd6Qzo7cdfKX
jQfEKbeqLprQMeJdnLdK+wS0ffqK6e8F+9rEK45lhvCJmbn100w4k6+fJxN43jjCFpM79IzJMnxY
nvfwaCLnpje4EzKs1/nK04dOl5GFXdVoAqpI9+fv66/Oe//uyTESBFiekR/TO7yg5sF7JFhvlh6q
uhqHRwDY7Z0I+6gWYvRMH7Tx4LMjCvOEjLNddF3axHTWiHPkYTzHa7Htlg68TK5tDmr2a8xkpfAH
RzpR0pUZfjyKHWJjhJ4A+5ccLxh4ryXSRWYN5dYUN3hq3p+9XTQa+A+SoOTNgdLld4sJikbCrDEH
8/7njK0ZPSCr85PHdC0E5GEM+7xuTLEFe5UxLTmhlQBUbpRRkS1SiQezsfwk1plXxFGrf8eLBAII
9y7YGf2j/3L2tV3702gDtZyqWj9MlryJNFuXPD6T59cJEOC/rHZtZSy/HyIHQ5F9Ul2H5eje0CVR
OJXkI7qA1/E1NHldDYcNQkcZFgLIgH4tKzFrtVoT/nZDTqbFPRzJmi32HTeNiM9VSjm67SUxbMX/
eT62KLd1sl3hV5nFp+gahDYWMvtIlQ9DRwyb6DPbqLHKkTOoMY8AJtOgrY+Ea00Hepzt0ZEQG2Kk
/wpUhsxPyOBx2dyQlqvGQ928/U6g3J5rQjg1iCWgdw/3NPSiZ26u0YbyD1Gwa8Ptq5PjUe+tNvel
C0v9FzASI5YQAWPS2dC202Pd3m7bGFj0kCS9WlaD2NUQZfB6oV4SQ4csgIkswZI+yKpihaB+JloN
ARNvS5PL8M8u129cuk6cm1KvY6a2HDgkI9S5ybzhEp13pd6fnLfvOPvYiotfeuRwUwArBlj8D4RZ
EMWhqiz8wgQyy1+5wVXCc0MGGMT9WDUy1ZtW48HQbHLLjgLS19AFruOTPy6oSUzPbE6H+EXibxwp
adAFvlKSFFFNbUqQq6uLDpmTQ2aMZ+/SzdLTmhULrBSrRSOJIZUWmc4so1ypKN1vadOghxYrAQe9
7PVnkIpi0o9K3ynMYEXGoaYYOMxJWpWeBUbbOqmpionGbcGMCjTFh/i25zOJyi9sek2SwO+zW2R8
QiQnRIHK6431Is3NabOZBLXmhcPRA0gwmy3wdQJrFkzNSd2ypcSmD//eeLhFG4iKhfJ11oyHhRSP
WKPjDezp5dWtPRY2vM9w/SGrYmG+owHmUjdbZBJ0kzSG7/60mQXMOx00+2t55yVLpMp81cbxakyl
5VJSTiBgYvekC2E11CJ3uj/r6sdhsoKB6MlksBzNGOCGA7k9vn33M7F0O6fX3wPH9TMpbwnNBWUX
9c9vXwhLiJC15xRh2Pyw/Lb5YcDpSk09qn7HPP7038PpA2mQgvxTj0mdzuoJWTDy9k4OPcpS0oo1
GBYNYx7A9M4LNAKVeHnUvGuo35qjX3QmvFyh20m2xu3rEpHlVcNbrtUoTc9SVZxG0IUdSjN6oUDH
Qk4A29zZK1XG3lUslPKS+iho9zWpn9Wqw4O4hz/dXTKF4YNqmte/K3Mr1PS3k5L61cD6MHPNZXiF
FUoI1rJFSToX0JF5Holvd4UVgqSJ+K/SQJLixHo6vnKb8i2yHRdFXcNOC9x2kEvjgomrDUM115+j
ykigundh8k1O/sTnMbDY34CHh/Wm+KLb6DLtmCVgKAVYEfm8r4rkLytxqiE7sqrvSdRa6axq5jwA
dvOymN7QQdhzCOeKx6SOciNW8Ageujo90Z3Z3UvW9/W+fVGvywhfogIl0Z1Rs2OSudxsOYS3vDko
0E5ZGQNRdIv+d/717pxRYPwUlkvcbrF4v48sQZexKaIJrRzmJPwfMipxYWAXEPyGD8y9Dh8yPDDU
7u16Ud8aQs99UhKe2wJr3BAJPkhbS0NmTcUxgrbBK4fy50DWyYGRh2y7aFDoBmSDKSa72bShlhVx
7omoqU4noIiMr5JmTJYixoKfRZ2Y1m47ZWKpXcOo3axYUUw4XfYDTPogNMo0DP7VE4HqwyW07xnZ
/Jx2YFHkyHcFVfjM9ElFjBAVteSKS42E+Ph+MwFt56cKROlNQJFnDvuBBBaO7RWjiRLDUse1MSE0
HLsY5jxO5bqCDS3PtvM+S9AHmN65TChpuq/pmRv53Rr99eIuwGqcl/sWMZmamN6hueET3ZKPdaq/
5K0X/yzm7WGYHcEzl93DLNCVzKZnC3guToQsfhYm6sNvtG7KQx/g3fneYWjVCeFtjLO+KoTcrAE1
DoVY6MoVLXwW2nZwPHHPAXdpdxU2LmTUMvdsCJFhy05HmHeu4lUFkM70AmbRnOkR1bc7geADe9E9
uEEewcyTwJsnjrTIHOPQYkHo03gzb9DahpP+lSNSisVeWHDEprqmgtjS7/F5rVNqjIpgr+pNXm/V
+hcZ1eyI+iz5DZu/d2GTqovkSiUnOXlzw90gi0Bol0+pyaXFmf30SBpW7jtSsWsIfjCLZaB/C1hH
1EiTL8F4hIoOqhzskREB5x9lHcJuYAk1XG9/xcN0FzsDlgtnfaw91WyNVzEm3jbizZu01Yu92wom
Sp+Gs7AcUZTkdzDRCu6ZFwqQm8tTY3K/DxGSh7352/0N3bvcAvv8KIIRDWeBdmICnIUQ85fhB3lA
D2zbr0EtEtBr8+p606tJ7FVzWSaXCBmDRRar/tqYlCAi4OPG1suAkyVrKN/rF3a3VU2K8VGjL1zU
LZyxBQDoqIuzPNLbGfezjAzbbx0EkP0WDKhIa0sStZ5jxZU+nmYAkxd05or+KwnJYmNUul09WHsK
sriHWHkJQE44qql0jPLvxNAgAg0YjY82GRLdYT+72YHRYhvjxck9k5Gy6AD8NUNL0zvnjHUJXOsB
WrehX81vK+3rK1yjBEVGRVPIe2QsvlnaMJRJx+GSplM/x/3c+UQ5Nij1w1hUtibsNWSOtY18GkLb
0vDrsnC70yt7zfc6Mze7pkcjdlnKMUpTwZdIyHIqV0vPRQoYsDXBuUWFTptz8R91RpLuSke22ebR
P2G6mkH3AU3rM0vGTyQ3KI1F7Y0F7Pho5sGZ8rLt1ijuVuFtcz4mQbh5q8bCNWAWmB6UG0hsw6Sz
g02s4SBcfTB4F6lnr7svW/ihPf/A4W6uaREgpHTB2RtUa/jE49Kj9TJhJkAY44s/voEqCxtn/V9v
PbbRIXqPr4mKp1PDT58Kpv0kTURcX9lqYld4QkT1OYqWGl7+fihMct/7O5/Dd7TWYw7yNPaSdxNc
43mWKqTsbbJyd1e2xL/e1zhN/XEOB8K/VM3NekVH8zwyZNLo4Ho6ekrsH+3mgHxESJrGRM/QqT3z
N2mwbBbdDjntaA7iPopvInlFO6K9sPTAxWtQZ+AE7sOrz9gHEmp/7EHMJsHr81ctqWFil6nn0PcM
212uwSE1UzQw2125CYIelfLr0JqtqTjX2/oY3nnf50O46OtYYPQfogxwgF4LzpXMcrZIoHyBDfZn
uAfOPBD2+YYduusRD7TkLo94kl9mSFfKes7ZO4mOqeuNXep/o24fjlLM2X+U3JSaND607J6gbBAd
SdPdN6iZerD5m35nH7Fv8Tu8Y1XdiDTght2CHUeNuUlqjL/mcugIVN5jgvn1u7qJuct2gNrATQyF
+31ZAquOpW1zmNRN4SBLi3xYPJY7Z0sLZlbvNThUOtBGehXcckPsb+fqPd/xtqAwDimTCZ1dH4yP
2hXPdEyCvay5W+vbU7A1lgwHgBSMZ1VYig498aPoJKrDwN/XxTRBRbrUmk1A+lpIDah3F8riZY22
HSiFpznK/YF2Qg5BqC5YRWo+mtAQ9PK/xzyGedh74FRwchZdRW519LV7+2bRzlfyzlg8afS7tyct
Nrq2ulZsAfYI/xkUqDdKPvaAq75gVsxrcPTPqZDNBJnyhW+pKU7yeYO78lOCqlWHIpvzmfqRdJW5
wE8AeZF+cM0fUyCBYfDjgr2EwAl6wLVp96Enmhxid2IMCA849rUoZbA8mLkw4CzVESne5ipkn+e6
df68XsfuhpxEiPrha/wUaUw14txjJd3t2hENSKV/UOS1p4IA4bfKcXnGIqdZkVA/aKQ8+Bg3Tz+I
AsE1+5irZtIh1n4urzkgQWR7XZad8rnlXvi+v5YTUsNcfQhSGubtCd9TJroxqviaV60RScvdEUZT
e+MCLd3xwvaB7RcZb7ItHy6MUvhrq6CqKWJ35nTNZWv6yeFnvPw0r0O62gXzpWP09/AtUexsz9w6
nPvakcc9FJhO7vT/7pE24t77H4FKgRiFwsphM77F9ttY+5zvPpN7gxi2Vy6nFmi0/FDdryKQvUhf
q/6+sme6SDUZHXO+aRIEQUQMXaRdQ9jATijKOuP3h8TyRBui0BQfDuEq7QIwXnwIsbrvGLBfRAG/
1ZFXPr0lHXcmRPrjto2PxpkcfPjjNeyKlMtuJayF4uKw4w5oH+CkzEVt76asKn+de8Q06pi+w+Nd
F8CdrjkEZT145d77ztMuM1FLVTwZAiBzUXSQH1uCYT33tXxTzc48DGWAJaH/yRIV3rWFnwg4BnHn
jA/RmYmG5CeTTVB7GoWjZKZHre2p8tfe8igdxXb4tSI47AVI8zhsUWHGpx6kkbcLl5Bo8CSgbYDD
K7WaCWzLA5bhVmBNmD2qnRZaRZ3z+wtJU2agQwvDTeiy42Pi9CWIuDbvKbzxpmn6SKCjB2Mp1q7Y
gN9NoRXP5Pgg6FCNc/WAAXjfWxN8aCDbwMtVmsBTL+W4/JT7YhlTqW65zi484+46Z7RrF/ahMs0N
/Akty5f6KtvOWyLc7/kj7Ep5Lw7uff0fACXrtyNK/9RrTTiXz0fWBNatIoCoQFtzFFo9MPs1r6IS
t93QAO9KIEftoIRoFMPRh+EhybnMW2lKiEdqBg7og03REz7JHCHGIrERDwFpGGnYw6L/fDKL6pka
tB0gTCgJCxfTnbpnwZ+1zRTInYospLSqFzxWa7BskJf9QisBy6zQ0yLDW47ZQOuo9DhlAsPWpwOV
PZF2LFtZGUJwHsVZSs4167WwDmsjLET/sBUMgi6WC42Uima8RgwXrlGUb87mPAOI4ghtg61BBeTP
etgeygSO0NUUCRV1I4tigFXRQ37LyzjGpXb2E72yA/VnjtagGXaeTZ092eYU1mbA+7R630ywEofo
+RAhpjXaPaVPLaEtwRUmuR7UqVWvZNkVIkP2aEMin0jRcb7T5QchVjfA++aSBrH0PYwmI9xozRpc
pnKyZbiMdeExVQPXQ2vpd30rE4opRGjvzMHZk3ZLClPaN10aXdii/XeJ6xYLSK3SWvCURHTmc2bI
a1jnXqgiQY74ZIuu0fFredcH3CPMfZR7Gw3MM4PAPDvUOrdMQm8irUG+y+/NZqGY3TGRmaC0kVCT
mCYaukED6S/P9Kat3XvdPu/5qY72ruhnKTO4XcZaPwwug0bPEFv6NmgKRlfty1BhVHgMjPQU99Fr
tLpfRoT8GL8AQ8Q6Vm+/HDXiuZCd6h8lAFuxsCHJjYMkwsrLPHgq7SCylop8p8tGLA/kswTjNWd9
S49QvbtMOLLVhXZh3Ut/aQnP5lLWCyPgvORmjcVPT+MiQ+FMrSE8hP8mVfsUuRLKfJOQ82mRYZ3z
2enuHYtg5lwQkXLBjnSTcS4HLOYRPEFk6scaV2n5rmpY2IlHb2CoWmqc7RwOIeiY916bzRLYLDhj
E93g+7TsnY4LhuJsaam5ohZ9jCmLIE5LVdfbq5N6iM7wIjnTXBWBl/78XXuW7Z1wyBl/Q5GV+qGY
HpX+GDHlqsyaYZt6wGFPDBnwiE/fRCKOnGXlwaTmB5SBcioFAKL3XetwVnimLpF8yt4g+ll4O/zw
GmYua2Temb30QqhXdaBF5Bmyf+ABY69Exm1IAWP4PDd3iEZ7cWsFe5Knbxx2Rrx3vtdbsQseVXCC
ZRLW7tbdKIcU+pUPa5mLppXyMjFYa2ZzZxTzW+73gVuTX3GzY7E/YJqc/5WYoaxUBPlqIWkxao0f
HITmVkutnOeUiz/WaCf8YWtI4HGWDN3rjxDrNM7AXv0Ch1fr1/xPWl/mYJW8Y9QmokKSUfo2goL7
InKxPa8QdHEIReWqzsYFyWflgAe27mDQuO9GJsNpotGq/owrOAvHTnSvkN+kcdaz1fhZ1fQ6y5YN
VEeLFmIjBGhfbsTx5wk87ALgcP5mC+eMc+vU8I3b8CT2GA+nthkqOYS63IPiVyNMf4O2q/Z+5u74
ALm2KY7gBZsja0btw8XWxx2BkqaFNbtposTNnhYmWCPwDrUmnkTSHBZOjEHSS5QfzCO+NXzYnvzr
VWCnln09REl/+eUeuLnnxU6eAfBW9QdbnNbzegCmpR+uAFF7s1DnNyaliwtqfq7y7IAxs30l7I06
kcUbRtJWUMaJInm8EfG/EpDc8N58sJAgSwsdGrfKR4qA/IJtUzIVtVjA/N4f6r1Rlm17h+r1fGOX
6zo/ISgwR+W+oxf7hUaq6y6UP0LrAvgw5uAItOr7lfixsVyIkyfMVvaJgeIldQw+62V/QfzEIwqx
SEZi7bITA71ExvPqw/ppwYvON5Ju0lOlhm65eQt6ARr3ou2lpM7f7FYDrED1GQs/wIyQK45gCG8M
XNRuzypS6r+o+N7h2+2gpP4S7dalNutGSz7Sj3gNVyh2HUM+kqGGfImBuC21RmqXTPqWN8E1cX7Z
W3hapqNQTKpt0niGWt+p6lpkWJxuHP93HjTulJBqotnBXRqsUyDb6cwmPPcuCEInvkDOL6PMWAJ2
b4xGsOas2FjaDoaKSa3Oj12Ry0JYt17kvhakQN9Xg5j2mqkcWnGqKJLfbnpVaIlGe1yZR8pLOuy3
x2v3Db+5/6Bb7I6BFblvrH9Z/9VSrLqVyKg+vvFSKj6z5i1Qx6hlKQkysng98Pupjsur9qErTBh7
0Ft5bvg2auRvkj9Ror2Rw15gfinbESs+YiE+PNJhgoI4PzXt9zXeHUws0QpMPQOEKYkHIO4vlNcq
Y7IYUnX6snLrKmW0fd1Bfq4NG1BmY6c/KJOnejETjZexOlzFDRmJeC2o+RNWVaRJzsIdJYKQrTLp
YMqJDKRIGkauuQ0i0JQp2YKxbPJylPbXuCHr+WynlWkdxCUrNlLgDUF8ZsOU4Nh/XVVP9JiCS6d3
NtOLwPgPedfQ/p/9gUx5TALm58d5qRBulxg5b//QEkN/hAyrhcou7FbIkamFNr6RNlIwX+pHbQu+
z7e1OgidSC+kxZzOhHnZnBjOzKMsqSjRXC4U6IUzioMjVvWcw1pDkH7w/d3FIkXKgCOIcngxa8fI
BSJgf2j26v9D+aaY6O1XJvOVLVVU3Dmz+jfsybS09TJ2W0iKQg8V07ZRwXn6PfiYGYsjWT76p3mf
wLiQ7rdzq7+T56NwHGRUb5iinsRWKF7R6+Ef1Yjpx0C006JNACpsVQrel2XPFc4Mq9lVe1YJlB/J
rjMJDnDsEbH3b1Qt56lguILT17V2NZo3zfzPRRRwnRBEClY3rMSD8SCKmNGIS2jegtNeuCG81m57
rGYBC6+CktvevM/veKUL/xipDLUF+tZw8ANxHSUNfsDKCfa4SUBoEoAaIo0j+rab1hAU+R1FkSZq
z18BW3JR2tlB10Qj31TGwbTz+QoxW+rV/8nXVnzwAR8LXGMURNQJuhdD3pIVbM39J6tC+9xGeZmg
LZnt6pV/nfx8okwOt4faxfRLG8P4HhK5jmYkHrDWbHZDclXU1NbR5fj4Y1JaZqV8mkUBv2v+7U38
hRh3xPJJj+D9OStQ750Q8qAZTXChoCcec+gPK2estQp2s4ev96PIfC1buMvrWR+09ebpM2QVysG3
UOmm3SjmpPU52lFLyja+uXsLPx75gTzHEOUY2iUOao1h8W+Zy2UcUvIuil0161tnS7WvlquDjtJE
O7x+iVKh9tH8iGbYQQCJPyWxssu94mI87Djj7brswTvRevnY20q3Z0y95KtPYkfHRW/D3tXrZzOK
MDc4CPms3y1/PbXlrEkQwjKnMAgGlqWPqvjLRHACpEfvT33kvDwR2cZo2VqVzGtwnRe/0mzLdWvP
UXkIDB43hciqIABH4zUwSlfKhdG1JFhyihCt04X1aylg5CUFKse7ZzmWVaQr8WHi9cWiadSg2sXV
FGpzM7XucZloX9uVXFMLtO8spXWg/zUQ+B6J9onRPDRNMAbECN32YGCqXkK1gOgXrBDPrBJVQ8CR
fW995fzDTp/3P8ZmvtfmrLOWHXxq4rf8la0UgaM1kctNezRO2VUaGZjS+zpwGHZ0IaanFYhdWiEF
MIlGle+yYH3OkkArPVQzA7awfLwr/RpGLWrEEa5PuRyYPUZGxaDQnQy6JlP7YZvKRjl6i84YmlaT
YUU0L+pc57mg1Q/LsAksN2aWgVtX1boWaesOA/kaL1EBL5a0e6v1E/vI5kT9AwM/NDua3+GjrnbS
ZCMZK0bCjOy7x8HRLRSKZOmegrbzrH/oslgUbaIjd3ToYYg1okS/cX4xcAPIssK9he9TaRtJmKCA
PpFZwa/LBv4t/NORe6RRbR405D90Rh5WlNGTf9KwMZoW82JpQSSlIXdgxct/Dxf62Vh9JkYacq8+
16EG/bIPAifvXGAhKjrsTaIXshW3A4imNN6dHEpMwFafy+X+V4iS32LWX+FpBZGi2ebjO6+uNp9A
9NT9O+FWyYbGx2GKCm6jN16UGrI773fkxhKyUu7mJOSsK4lUPnh1aWPUnbKBjAWd+JZT9Y9DErPn
/fgEtjgjkBMDubWnRBtpCNZXjND6yHJZ+ywmga6W6uIyw7oAYC+pmPvXuIpBVI9Nv1AtITPm1mLL
2MOWws6smqvgmUWfJiO1OTy0CMSdiLsUCilN0xhqIm/3xtN2QSMJeydbSgvnAXi+PK1T3GLQtxWc
klxO35Th4Zucm0C95EjNnz4RU/s2fUPzylgovq/2XRWX9MtrKlR7yhDaVR2ZDrcL8ubkgL4i1+le
ifiyn9wcaQA/SG3OQa84e0fm29bGlr91TqgY8RqFQ0LhN2lk5czwQ/F8sNq2l8rjKWfa/R3Qygru
2uxuRLHMZ/iInr+mFInF3rL8aQW3yEIN2u92oMFPYkHBNwo0HwEITP22GM5sA/hQjQSv8fETHKQS
OrTR/ZlA3GNqIMbTy2t8m58Vi+BFGcWAaw4sFhfIA/ITDbvG86Mg9vVaxPafqHegH/SMARPetNgg
DA41/aducrZFRJo1OBrlV+OmCfU/hTAtSbaVFfMBsqVFMiUmbrTPKRyXqS5t1QGx94JVipip9UcG
zDsXCooJ/wqTNo8VnmqzLQFWO3UIyyBaiYFhQJ+M518x4fCyxJKhiE2UNPqV5ANnDtkj2J6SQe4C
djXxXg9GgXvczqfSpwbxaU4XyUJsCv5bqdxlvn6uzHJSXaOfQVcRhcvnLIEk464q+R0zTMHjWUF2
j/O8ExiYrbfHofElyrYQVT9OxDYISnCokGom/QnqIq/Qs32rvYCsw9cX7Y/ceeWKhLqcqWg7XbU+
UkHSEqJASqIzwUxJTKSnqzcDGqXWxgYe88k8U27KcJM6DPRdfZjPFf1RgcM1FW8tXF9/7B3rJ5BR
O5aSpzavNfd6CqEfFGIdgdV1fw347NZrZhR/2IDG4GjywthbOb9hLHETVrIYKP71qjhBQZ6pLZWD
yMwX8w86x5/z8P01zlqhzCxwHzWMcxfe7rsuv6oWNuwrudO1bqxLRr1erOVhwWmiyw+m7iMeK5P7
xXMT7jGhLII2hu9Ol5JOeixsOMKINlhsO9O7lf+icZcaconncW6Jv9bAdVDfrGYY9OQpQl0ROyg4
Cg2VSsTsK/aynKCPCzflq9RYjCMzz40fA91dPTvN749dR1XkghSw2hoB6fO1M4isj5JkQZ/4pvE4
QDujObgxb4z7d74Vom9MiwZVCKHWl2rlBmt1Sns1NCMPQ7Sh0p/g0No3o9rXoMVqNjs4Q08BcGYV
WNlf53kZ87YxPZeiSvCd7ImL/BlVO2xYhPk3sZBb3N+PN49QMxPHYWl4lno3uD7MKvG6vGG3jkra
C9wKwdj3Hx9BMdTu6DWLN5FrmDJm8BWoDMOidBHTu7cZ7LS7SYMBIAcmqO9ZdAjS/zIbckznHDEC
XltcF74UPxI4EYau6ZhuyFQFGuWgFHaUuL3CZQJ+vnLnq4/hluJUIjVx3wtU8qi84PzjcaHObdm5
QeysvWjlNGaPPBWpsO+wg/+CrckCzLLtEk9UVs+cWetsiXsl+9bK9iECJP6EWa0z8BHrS6csWiDW
goEDSCJjfdo8b9N6Qm/IakN/LFmiBNVamXexjUBBnCNCYmB+Yj2MfY5Hkh7JgtvXFMeVwSjFfUw4
uKl3evAJLsL7qeHtWQmz8VVraIXvVNNzr+wajuVYbS8TixxBfzj3QnqdXQupSoYXV4aJLzuy/M8E
rHEyfw9HvPdO1Ju4hAaG2IlQ8PMbb7h6Fw0ozGAGHzovc1nDqWaJ9oVFC1RUhPcNI3EIYwcvk6RP
y+0g31g5cv8K7+WYxGqUKzw4B+58n4zS+cryeivK++LHVljuPItDtHp3HU9Lmguu0r1oSzOPPLPQ
FjQqJ0dbqs+OsDart38BmUvXjxsEZsRLUFtu+DplPdzn+5gTEyDmpwqV+9wghtxG3nH8NlwR2cK4
u3Vk/GYKCCM+w3c7p3ZJD5rsvbafn2cgIAZnx2MZ8ZMK8Wn9qFBk0jHKYq49Y9luWj9nZOPAMh33
4ZW5F4loDurxpvNCY65E2yDNfxrJSW2CTM5TuCE5Gaq3j95kCBVz183SfMaGs51+bb9p6afPbAqU
jpUISK7hXMq8DLTSWV/R9YmAznhNetKM5VUs8aa99VMKou8Hz2HwWbc6wtM3SXZEbW8tsEXHSU95
ZhbtmvkUVfkGp2pcdc8SEBZR+DYwlOT/YcCQ9L7W5OqnEbv2LRPPgWHZTCWbcQHxfb39D7MRA2fm
giOOnsD0omInJqYoLdeb08ii37YxrzT7p6pljBEnr8Z2qraORIJju4SVFz59KI0UPynzHmxzSll4
9AFyBLLXUcGFaUJCctyGnqT2FBtwNE8N1ZpJaoaFGKVObNBUE60/PsuKkow71Wxry4t6Si4w8AKV
fynjM9iVIZlBWhF1SSRsQWDBVQFQimTEdOsyuYrBOGYgjgzfTE+Uo+rMkcagiTcXcCnD8G+OqOcU
a8ZY2zOueY6jLsHzu9Zw4X9FTkD0ZBspoizRqJTxZTYD/nupisze8Td/claymAigvd6mdVA3xeFU
Sf+pa038hlGm6+JOCPRRL6D4mzBoQ5SVT6Qeeyj4aoodKVndL2OnLlMjCjmq9GEk0Kw5VDhtAV1h
xWxxtn4b8TpZzWlaLejvOGray+ErhVyyU6eH/8+79qWIKNKYQfvQBHKoEP+qi6oGAdMgBXPeoKwS
RXtvRIrVfAyrIVqLhbEyRwgLdbqYYQVL1aFVv6tIhw6edO3zocW8wF5Cm64d819I5OCFWOiRGcU4
Fm/FPw97U0IQjrGfMo4PB70DDOKWp/wR1HOJ5lMsGGjdEugWBTgH5fH6hJPD+AK9dhQTaBpeS60i
81xxvzx44zV4LsprJRKvmLQYomh2d0Sww2RG+i9A+MV0bDT+cZoLtYtbGNH/dvuQwhTTMwfsfpGT
UYVXswJzqkvgjFNkSm2hDSBdyX6j/cheZCyerFwbuBrT0w+IAYvbQ4HW2OQmkT7XZprqtnqE+djV
z2+gjLS5KWv8/YG81yKaD2qwg4p7EC+ontszFDQIElLAPV5Ifg2Lts02hzHnEaMjQEGuQ9AS5M3l
4W7N2NEZCwh6LX4PPn09E8ND6pMkZk4P6VC8y0o/jo9k0sqFtrcxc04PngaGieRtElSZ5ok1WYjC
tWgrZ+u5Pyk6pfCkkZwfMBAoA0N2/o0EAcB84GDNiJsXAkeRu9yrgEAiG1GAqBwcE4t0FcWMdB2q
opv4P1FRU8iGmmatXHqRSNc2Xk7CO5GJvePpUSDK89BDDeWpNkhfDziUPMJpWCsQD84YnY0L96fQ
F0oSIcq6j5rV96zYlok1b/cqrzl2H0jxSjDZlMKyAeJiIFRb6q6bCpIMzulzHMF6sLwHoMajvIBe
fTnJQ4mNNpLD3j4l/aHzuk2NyNaMXrTzwnTc9gFQCdyEGHKjpy63hvGANXq64/9XMGsvDLoyxGC6
0/zk4inroLYzUT9740w46K0KXC33nrWKv4deIHdcV9hKsrPMrlHFOeQDOPMHcepbGw1wm1/KddR5
E2AWE3AbJxLk5+WQ8qayrE7ftttSdLfy8GNWdtZxLr+Y6nQcvn8tFg50yRMJjabqlvamGN0pkSzK
T226G2/MZwKQ29rrvTrHQkPzku656lNAik9wS1A62ypa+1wSRf9HzNHgZVQRlCCQs7Oy73MitQpA
mU7cOK58CI4Ucb/31mNK67AFTzzcXKFFtfJGykcnosCGOGE/1ASR8vHyQm7v0HEp8iSZ62wfttC+
36ppwE3Xp8w8058wcZvrakcsgTyfWkb9Ujsjqvcln/2O51XlNshfQx2q4Veo8qk1QbGue/PB8pZk
WKfGf3JtsI0LHn5cD9u8QIVfRyxCnp8vxPe07NCuzx/V4oTJBBdX/Oj0e6ak2Wyg9dIV3gFScfBC
sB3PQQxj4ku952y8qY51niazVRZZI5TRfPvUw19qZIRg7cUIvCu+GIB6v2B3QcnsukaRP/eY5GQz
6MqkXZziZd07Z06lIv8vewry+v3zfUkGr5I+wdW0F2/8j4nkFc0yk5nhtccf9Ktz0vpC5p1DGHIj
JCavURQvYIkGmDaMO3HLYVCxxE6ftW3ncvnHVWac+t59ebQkdePud6LKmapLigpHq41uHINuiozs
+VnWjgAMK0Jo7zRBK1lQpt55VjkiW7OsDWVT2fGnU0Ov6k+DfhGDuHTDrZWRMUNXdlSQxmubDy32
cJHNzsOgmkPCsdoh96cPg/Ja7TIM3rNiOpLfxT1Na+/xUUUZJ3rS2FwU2cDC1jNDS68gWFgzv8xB
7ykllewdZjFEWEsI2o8Cg62yyFi+ARJiQoztACEm5yQPf2i+HrF0BtMgHwH4//eJMKj9q2YoF7NA
BOLm0jhqpfG9qA5UYB0JcnUm/m71l1V/auTUclbM+965KvpVsdpXraeA1GaCC944zeatXrjKYTXf
8Z1CNpoh6MNbDA/nWw31iUpjmCR52cVxVLRcRkFtRNv7GMdagjWJYz7dKLtyWgNTrOlVg+ri95Ad
JzVwL3w3BsChp1OIwZQyuvnWqlcRD3mcEClUJoaeRRTQOva3LXCGuSoAWkJuSv2/CRKKvGSthVIb
x/9X0H8rBnC8IOQUEQMSOuSciq+hkeS/nkZH8JD/CRqNxxaQyo+r4JDkTlJFGhCrTI1O4X8fVfiH
v3CurosRzzg27E7MWbqPbURpSJlPYHfHvSWATqDsw3JSjZ8Gjzq/MUVSrNP2D6RcdslClfVy8bVz
ii+ZBXfo9oyRrHh3/Ez8kLoh7lgNPMHgNKbdCjFWoBdXG+LqPCHZ4ins6QGibs3NJ08KsIvfZMqj
6VLH8D9me/3Kv61g0II8VvPhyw/IL5ljv73RxCMIKROXoXOJ4BU+uQolP+Y4qRHQ+K1CMflr7L7e
1bGo/VlsGhDwGZXdgDtODWte0ygP++wsQlytY9fL9f207hfQ0hpQM0+7q1qQz8A67yAPOHAX8NTA
l9nU9RlWuHE/rRdZvle2ewX2paiRX2ng0n08wePnqes0FVYVJsLczOxut4MSs9SMvQNxgmSK362A
Y4twH0EuGvxlzKpjfMoLnaC87hBxdJyZixDBw540Ys/htRiMhPZxRnq/hRYAJhGkDSQSmXe07buH
mNgs7cROXgvVSZ9tuvwySUWMQp/FAKnl7LVDdSsVLtKcLdAaU7IfD+QH8V9xRTKgk9BTuE1ua7ga
Vvuc0sRFUDZ9VV4j+9v4F5IzRtUWTPAG3a8x8C23ckgST5s5LHyh72qMUFKDwG8RNAfkxp6xEYzk
IoCR1h8p5/hvCVcqhutYbIWwB3v4/qvdpw0aQjL6V371D6vUXn57+e9Q3KinqpV26Z6si2swVnSy
+Gs+DAKwmhZ9i5bthMIM7SHBZMYWno8pLvawgPJdtGi0VZqoqSYikkH6f1k3OsnoWQOYRx/nLpWD
RMT/HM5Me0S3kwuOfqHGPPwNodLjRN8gSsKJsDpByTz3BO9Klf/3rM9QAa5U2vgy/S84mntY3WWn
DzYmZS7pFgz1t399oUpK8F1YGKf2d//+ec05m7h1HHmFPBI8i8OmuzoDPUAP9VNd22Ro4s1vlq4t
+KF+dwGIfOqrB7/dxWB3cBA2yBayjwU6ZX1SvsqiBNnrcjDWY/uEXPVdOvmlX+4FTz6uWrAqPN33
0BtSFXpRiIa+y6CmFQw94NygzlU/rTV9P4Kj/lBYMSuYDB183ohchDzQwGdK4H5H89FK0K42zWrY
aeXU5sTTwQ4mwU1B9kJNeeoGekyd9p/uu32cJ7sfrt1+dwXfnhe4Zk/g9AwZRsG0/+fA90J8jOQE
OPvpHlENcVTJT5KEDRZ9Xi9dH4yD2UyP5bFwrIw7RfGEuZo2YmxMpPt8uZUJZ9l9s9nnN8ry/t8Q
CXb9jFXgmJCSwxYUxXbgFViXKlLPP0fJohmeWqP5EvtQG5lw9fykw1G1RNAQRhHjJ1baXIe5bU9w
CE1E5uw3AVGN8B8cemHiRwjyWGTBq4SC1SwKhHmeQ6Ki9e+OhBX0fSAOEsm866fU3n+EoGUpHu8U
B8bB/ylm29jctRemBuh8XrBBXJBrxHl8wUpAV+0TYZGbtAzjBXdhmcgYH6alfsOhgk4Yc3F9yDIV
eSHuLihgFL4Lpv+OBdBVVC4SU/hevuJ/ORlzs1njBl2p3og6m9FmtpVds7XHiYBi3wGhVt7mmdBl
TvE0pvz5HQ00HaXtuoEp5jedc4jPh9k2AACVl99aj8ORwHivp/9QQfNTB79Hje3VfdGT7fVge0PU
k7MY2gB3Humdj6UWFu78a059KTaaqWSd5Ios06Rlm7JxK/ufH3NvcvHCsMvkSE3xXH340CuBbu97
UyGkrZqH1sUAk6CS/eyGy12KS4fGHKJyKl4uOjlkrzzB/PmyvNXi1JlJfsQ2lcQK37zO6AYVlGq6
KmQ/cOEEZPj8cuY2OvNvYe6v4GRn+zAl/hnVFlVfe8Tf6V6qdE+R04hBqfo+3irKpsd0Lqayw3GO
l1OD+/SIfl589xPN68ujDGBRVNJw5JVf++X330wepG21079+bK/HvSUXsgmU2nrPNlf8Fm+YiaR8
cFf6pq03v5CGlHh9cQoLryXcvUpoKX7FBh+x6D5GM2sRyrle6KUS0DD6quAiEdYrVmxOTKTn/uxf
B+irbsgINg3TpiWd6TiEXfOQlWsbvJXD9GER+mPdJhz2AoaPRFxvTBqul3ToDhTzdCsxPxneG6PT
ztUolnGmKxBfyACHrzbKz5XHIivRzBCRP1wcuOUedv2hoO4cZOa7XGyY6M6WLSaEu9GUnY25cCe3
d9TPz4nLqLIQO7YN6mPl5qZQtFa74JTUl0n/PLnQkv8CplUhNcKsfpSaKGGum/4hpECkK42L263d
r2qfiGfADff50uqC/IFOV0y5ypXJcdYSqcVrjNMkRds9wWaT0TlJuO5h26OCJRPZ2EKvpXevZzKx
7ITw5wsK3HeZMiZJbFpdmK6FaekzRkrBvK0jJdC1V9CX0ox2NZz4SRr8Raz1/ubxZY8+V/gH0JHA
x+2S0pDJVu1KSo+AxZKLKob762UocoB8zGwWZr5bcUSQshRczLQ1H49GhUmXgwC6D8KYJHFtC9Y3
7Qdg4nkJ+V+q7Kw2TPkIUNmy0JJLg/CN0vdwk1jsIJgjLJ7wi5FbSBFpvAqroAINxfkRldhRCcyF
lCTFCoX4atkhoF900CQ4AFItWURllD3uOk473wniJjiqKL6oJHq3zVXNZrsaquTajaKvBgdTyU0J
uRjnJGLHTk9GmPJP+XN5E8GQDToA06yeqCVKJScyo7FkvLz81Un564BQkhwk/AqVzvlmL6L7MPt/
uUxw6enAA8wby+WmuV6PEtSu7FATHy28Wd8yZjn/QkOMgHy6oquNdIeJ1ql3dePhQBVhkc56+dcv
uBPUKL5dQn3NLRk0UFPzFtGEJZvm8hmT7WIDbrEcaj2rD2smEe89uChRhsJjXMk+NW3XxFt4QQQ1
CWSTaCDQ3/+iRCCZt/6WewHe+eRG7sGgeKZZCtG7txEPccp5fa6jYQPerIKW8/i9Q5ay7NRQDezM
lGc1LQ5A+XnWxsWyB/134BFesDPrUkeSayIEQDqx/3DOZ7jDBqnxYLtsQu1HT9VXeJOenIv8ySnW
55dJ68EFoxcSpssXzxo/gBSznE0b2uEh2T1KheWI+tJl0Iurf18GlwRdusDai4IAjCcpZ6MLuIcL
9kR55+hFFnmbGRCJNzHJ2uhGOvE30/8sStRO1gqwkJ1T3ZklSkDpomI69OAfr9aRxnOa2DDLF+/c
qky/6hnvA7NgP2/2MhHeZbMKd95qJQuOosPnd69GTwRfTCybKeuX6mRTRUTmrr4h95j7+SuHtKcX
kjH04gPSQzcZbQJjl07pQduhvIB/yxY35agTobUe
`pragma protect end_protected
