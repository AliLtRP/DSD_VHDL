// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:34 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
fIwt+SDasQ8CHIHQIIbKkxP3iH0O26o30un8ehHN4bVDPYziPhsjoiupRHgA6jxS
t0AG51/5TE3jmVghQOKwlMLByipUTzuL8BZHyF87lS5GJAxgrFyHe1Ywafut+11I
1inELwQ4W3RMKcTDSC0XHI+O+9aVxjIL9s/wu0r7L4o=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 19056)
WkfM4doKg/WuK4rfQjtVCaO1RN5kiPrNto7MFtoeZIOM9pamA/a/qvV9QZT/2kXF
64lK0APq5YaAYdRSEwXxai8DvGEWJdBWo7wUtUvzA/0Wum33WqCgvdKFykjD1bEs
MDZ4BlXg2CyO9XbcVwBBLIYV8Uc7obQOAz9No2x1qslKbX3nh2+9R56ipEycFTDZ
lhBPS39pEy/aT/LsjmRlLN/y/edPM0uJqdC+QdysrLB1zOhjWV1+fngqffkkRRzk
s9FHSghvHmTJCqiq2lE61etPES0LjbAhQX6uNvkZOC/mC5yCHOaJ0cxSlQ973QJg
cgdqnngHQFdJpVl/vhZkP4ze89Rvse05in+vVdsKAZPnC8InT1Q4clYgpTzu3mwn
lljTxbNHUJzHrY6AZxpMPRD1sfnu5h0JeBJZKBKWZKbwVLUj+j4WkwxCrugI6udo
z6l3Xs5RLNJw7WPLXsau1D8HYmITlcRFQWopX5gf1t5M2Q1OtUHqZ4/jCzpNJTee
XgRNMCDiurk4GpcHP4VTybpFsOB/F4wnQtXuetPyO3ce+KRrQrzXvLNBbx1Mc6yr
1XKAY80gvpld64sb5ccNdO+v1F3DxAzfScPVvdNLqOUch+vyY4PuOFWUxOCEpT4b
fetojDENN1zUeBmLfeXFst8j0SgzoQZ+RMQrU2WWa8w3MeGMewzU4OSeQUfEvM1Z
1kys6pj35mgkDBQOy/bOjTJhSBarhVtIVLVI1SoQy/nbz+Ca5WaAW4SiP7R8/R54
xOmVclAObWfBtL75rUBPR0ebXudaPhQdoir+WipqQSeo4Dd4um/bqLoi7s3os6l/
S6tZ0/SFxs6mjHIcPBPkIBKt4nhHowx/sszm0cuu3Xn8C+QPukkkPvQvrvXFMUJm
+KTqLDEkNp/2xgel3P0lW8FSTNA56FHOI//oGr6NfFsK6BYixh3trc6xJteJJEO4
AFisKTXk4oUy5Yzrr4YNiOSf/MFVvPs+8MqdmoMDC2pelj4NWOCIYFdOHts0G1kr
RhyvLiaL44tqdMmUVKNefPQKpSlfWrm1v6/bGWc2thmhQgSWdzDgogelq/JTkd4O
iuX+tcuUyQSjprbNKFBIFYaG9e7eSlqFFMZjrFUZMqupY9lVi8RmB0awUHKQ/kj+
2wvGFE2H9u9aLRymT4dfn0PziduZM9ZLvCZJRK7BxjfjJrVXpbBeGKlCtU6LAEtH
DrmXjOgDT7aMbbW+t9Q9aLs9PmvdYFhJL2OlCjwiZb3JkTd/H39Z+EC74/4VDpjw
j7lFFlJTEzYkC7sWKAhEyG4knyZVg/M7XDmCOEOF5lQuKq3lM3kjATvr4HGexZY9
ryotm2Re07Jm+0bPwdWPwRuHSmuDKuKawpx7KjyLSv62EPpRA293yzwfgaAioCKn
rd0kAFakG9S51hqW0CTSRyRSZJXdRoWUljZWEUaauY5qY1eON0jaKDj8jULUhv0k
lzXMaiyX9AQ6vAs31OCVm2SNHr2G1Cgz/lbYzH0FEFJ14kETHaTVLl6eFRTXAeip
26vrjDAqEfaR3gIcQXMIemJMqE8ohtLlmJofXc/wo4JoUFH7x6DwI34eUt+j6XBz
yDyH5T8DkqrIWtcPJiffyGLgZ/CODDexw3OI20JcehEXvdTBU+Q0MZ+JZexurUmz
qKDjsBCQNOQQdQu5+NxSrwEB619X0CuArhkPb4O+PXxkaVPQwradtky4zO/+IiOc
+mKNKedj6pa6/sUmMAzwQxh03Gqi8QWPYfp8Fk1586dibGUwhZQWQzS0kxxQ8Elo
NjlkdvqOtqPBmqWUaVZRmoENlWx7ZGywxK3ASelg6jApLLe03Gc9vYv3TeCvwdOK
rcQY7COd+TluAuZ/Y6XgUzsRAo7wzbeS1uVywmO4Iz8AU7zMPvG0m9w6k2MoEL1A
xcTcjstdODiecvISMONrerYR5DKtQzyMUk0kZJBIdlmNbIbT93Fevs3ffRNhST5/
rOz0AnMJ8nWHjf0cAloPfrhdNVXspSRB9yBGtbOMkscA+w+e1af70vkrWoG9xKNP
EV17hoUMgRBLH46A6kXpVjgqLETmhl35pMOZhiivLGFFQJpXNYNmZ9v5nMSkcaue
ryBkdxSchpb77gKLYCXN1lt3dtolAk9apZfV09OUCpcEv7VCkO9Gy3P6vEimES9m
ezjmoNVhbbbN9uVNeHvAXxQCqYQixytGt/n08mbqVWxz4JJlaWo8stdDLmNOBdyC
8nkBcM9hwJEpgUy7GiJ1dkI3BzSUogG/YlxYMxvr0hEQRNmpVyE9ATCuXG/g1tNx
zYYXFZ4tlm6F8FMdKMGV8XXXJMuLk80kpt/bHJuj7bniznK69u7VpO5E5a4Etu5V
y94VKtapeOxfcHbZqsgU3NIAPJjzqI0kWl7DVddn3gJUiSmtkamfsoY8OW8Bqvua
+RBWUAXiJRdy1KZeEgvwVTkjqC3Zr8p0wA+8SpPeqAGDP7Vfp2jfssdFflyjYvfo
XFpKnjnLXOALRJcgomRObnfMgoTnt8SdPHFCVKDCAb16ax1TfE9PL/36QWMigYw0
aqL6bnzFdp9+tVnUKS+GYfqOehWcVwNl+PDwQoMloM14lKFjFEGud0Yisoza2m2n
4vnQyZ+HBDxWA0hp5OiIPN7jQys0VvDah1NPhiiSt52rTsDQUNt7EKfCHKVNqAu2
rVbdiIE4vy/PQa7EWKBjskPpyAt4R9PJiq++/xHdpKIVya2j9I5K1eT5aYW5QnIw
PCSUMM4ezHid96+2qPEk0eWk49HuHgiyioOLTpIaz/8vHl39/MDu8B0nRWJRQzWz
fumSJ0LUk/BAuLV0m6ndxpQ8A9qrSQO24uArKRNBD4qGzNOdrwxxUWePSJV2gBR3
xwHgpYd7u25z0jlmCvH2PoYVdk32wzC19ujurEaOQyKgsHYc+Le4h6kP8sdUw3RV
oNDtghi5FO3wgHkEOStwQEIuA8EBzq7FBWMAgYgjWtaaQzFwuZB/4xeEj15RoNw3
i88AVeIeuvL4Udh8PZA9g5lvdsknM7f7yw3ZO1hxu4pOorh27VztORsKFvYah2gU
Eu4PKRcsFeeWEMpXJOXQjr2SygyIivmo52YDOZjHY5kbBP3C9oxrttRnaffczVir
d/8CaSLG2uAeSIMG/YUVYDzSpMpN6tfAZeFcn4/H17yjWeQN2r4+MaB4fbvb7ept
6kC2pXZDPLjkb3lj0hbHyCwSiCN34sLDlMzJTdJEvoaM3i4W05Jylma++mFTrcPj
9TeYEKLDItpIjYmcpY2Q+omLSJS0hc57S3NSwe6ReQWGjbU59lnHYNbfei90eu1W
6dSGfkqhTDqT2Ha5RTxssbpz0Dyl94e7Ex3fLwucTAXezZCDQ+RTBXtIyFVjKHSi
Z31GgVjKgTORaEmB9gF+RNTP70aRA7cZF97+z8AuVakKawTDuOqpzlWzq49VPfOC
8W4HOirmweObnR7I2ngHPFmQnE4Mq+e8MejduB/z4NK9PBfbat5y7emoNhIb8XkP
X1h2Xa+5yacOhvQ/auXx+nouJ4RdkSsBDhlIm9PEaqyLSH7/PabLpdfmXil4P4yz
XZikJQHiazte52EpGBmNnxEHYnSL7qfwr6/gfqUWTUNUIFOtu0pBXJuMJLcXpFQO
d3D07WN6bVrNSW07RM0rsVwJYtwQod/qy9IH4aOEaK0bzaWQFi6GovGLSx+5G6nH
M5E5eB4wJFxt9DZwq1qDOBepn/hXSdCDIz972xmj+x464IRxOH2t9xBGrhUnXDXU
t9TlydMHoTYTd+nZ62KNk2K1F8vmSkMKIkjlGK8fTLYG2KeK6c1B1YjgHNbXA1Qv
qWkBkOgER+JdzQNa6nxf2eRWnUWbXSa0gZxNoClibqG28YOwkKTNLIUb+ixweKNm
HdVbOi1wnxwrpevUFfchlUwaIxOhoe9Zkh3H5kEEqfHuq+H4MKvCkNgZ2xTIOAKY
zVuWJLLSE5i07QCKL5ke82qSoCUjxQBr/3qKoFSt59+gLOB9AF+JAusB3VP74gER
xB4x4qA7p7fVH2RsrMQMiZ/66sqViF/VIBys76f/eY09qfmUi5u+8FbguBGGSmye
eFlZQ05haBAYSTgDv78S3385FbVFHPKqxpSXHC85UAvF9wBTuc49nfVGJ5WxSwpd
ft8N+6SlLIZ6INlClN0F436y2wMXPTBurt3ZQfCq76avjUTU9yZ3Prh+hbUXVUTK
femmSWvGFx+N0AA/h+5I9qllfmOL66tVxz063EO4hAYO/JO2crfcEfNBefrlllll
OL8j0TiBnlUkiJve5bN/J+rnWT0B/sb7qv3Za0RdFLTBW3mnnXUVSYAFlyDHMNSX
Ix1+jfqDPiJGRT6SpYvPe/iYS9W/fO5lvA31bSRdZgYCoWvB5pbdj2FzLz/XmESn
bfnO4Iz0oPqylR0enH4YmdoLd4gwHF4yKKcDn8FEe29LwRXl7N9rpoaePm+gX9+Z
qkTMVCnAIIkcIS/f0eAqZVfT5A3i0D3vtaQ9RTd0EEMFuHaWBvzyVvdN/FLtsHF+
gf0NqiOn0fZLYsUsLWLqjh3GZ/cmZ48/5GKSmAxJgkoW9zkPP7Bn5oVAFtVPZaml
j/KTfSZotT4PepxBDcN/Jz7JSvIuBS3RYEMb5eSKqYaxq93K59/CBZXSN3j8N5+8
fES/OEvSouZ+NF1ZB+DDb80G72fdblWiLXUXSh0MkMzG4mmX2qVjXQbI9jsSJK0a
ruYMwLuS8xU1m2If3jS8cqevbhHfug4UwCN01bgsHTeWzW/QmC2GkoUZKLpJSLko
ctmF8xxELAC3OvN8gZkvVTVxSC222UMi2g5bVCwer45AB900olpfZyPSVHNx4pzX
i699TTC9MApWg3R1Ev2Nz/NXJuuT18Jpyzb3uwrcv1oZg+KF42rmpRpZfzRi5+83
WD6oG5qs9neQv81Wo0MYjhpP+QXe3QbfW7tI6piFbefFzLYcziwh1fUTjXd5Wezy
cdqKa1NyFZcDE/wa54gQJ6uqkvPgWx6qfkhEZZbFS0TsFg0qnFLjamHwq6YWs188
FrLTEER/F2VymKyiKW21l25AhQ9yi177cDjmu89nlXYH9vk/ylTmsfE3witSH9zk
8YqVfoJ2JIpnvlxxahZieaZZqaBQciEPVpW5B8cy/7WQ1Ai/jy+3xd1rGSvAz5Ak
S+3fME0v0pLC/dJBrj2EWrrzldj5ialVuAmQB0xb1jWdobCLsNaAjaHRsc8QMIb6
Lk9wYLdsirAr0C4+bAOsv38Dtfth1/J9JvnnEuc8UKB2UW9CmKqDEbB7uuBJ6KHx
UlruGsQhY7p2jzvD0dHEdQNkIQg4Pf+asAR8pu5NzjdJqonR7uoAA/AENI5KxsDG
lrf5KfcTnwmEv41roI4/ur8WCdm1HDodXrvnH+ZVwy57ZhRnjVIA/nw9oI4Eu+hg
G7t3nZRkpCK2fmKv8gsLYYQBJ2z4rqJqCLdXp3hTFuMAQ4K5qmb9AyDS2x54dpH7
Iui3/bM0OIr/kT3j/IULj6bUTLq1YoVJ9bR14GPxs3D7Fyuat/au77hDLjZuW5Li
RggDllgUor1J5ej00Eu6/UpNHqmgAQgBWqbVu+ssvwU5sWYV0UJz9HDedKdtRPPR
4ktDL4xqxCGKJRe9VnHq4Z4QEoR/UEA+Ygma/w2ml2QYiomw8cQYr5kJhb8JTi/X
Tk2EGQn7462X7nc7uQr5lWozaqJBX38UBeHl/abUvKhbTpGdamaHqlMFssMoQek8
d74h64H60CmcEQ4mBOOrTXUjdJC415HLSx9cA8XyRRZTLhyPKLPAb4cS1mnqtQwh
ioQ8j3CwOPVGIlncd4ogPMUwVhAlwG+mwBSwGuGOKKHi99YnWClQjYRaJ/Xkh+I6
/STCyoVBmlg+CknbcZAJFHWAeRPdAa1eRoQA4EIikfDEErjrPbZAhy8+Hw4NX3hW
E4PcopXogLDjzyPVXh/dC/MlVwzkK72Lfckj9sKyXejRfIqpEWY3m8pmTNHrwYUF
HN+2XQdpnJtoYZdXvYbnCZj2qlsQ6awTKjib2oDcD3hZXQuXT/mJfkcTYifQmXJF
cmehmmZb4LvIdarFyu/APksDShuvrYxUsax9lBqD3GpRL7jfVIEqp5nEGAjOl3xq
Wr6rWdSz2KoMRA5xFedFO75iR2qL0nVLJpoaCManY1onZNxqV0Tm7JmTecw+8rSa
mh8ap7r4i5GCgBlAAOvOyrO8J/g+QbD2tA2XXZsmaqfz7VLgWDlsFuZV7BtkLKnY
p8EwJb7lCEV8yPsiqp8DMzy/5ArC9LeQU2KzVidK727msYLPYkFN/Y8vaEqJcRdn
usAoYkn1c51Gj/UgNzkzMLpmR1mUL/zWmj/m3p7LMt4TL4A8pD/nlOO1Taq3oSZM
5Es1SDRDEwb6J5dZddCL3YOKWBKOOLXRkwLnspbLKBOUHRX2h0tSgsOhQ8PBDkmd
UwZXF4vLtAAxwchdYIZUlb1Obz3Q13z8+1+7RwOXom6ftBIgqNGQg1wqnB+VFLdY
21uEdNAaOiwpQuO9GjA3Whd6mBnQB+laZwKaudguCJCPJosb6UxHeDEVEb17qbll
5ywABCmInhcGYdH85bBsOo+ERjIOlbqWQk8cKazDYKRlRlfl4MVTLD43QLadZtjo
ko1382QZiPTt1I0ECX/1UWAkOAzcahDcCB1PVCGbOnuhUhLTNgV8TrjxBibU1npp
M18GBaFHYZCETyazgICnVPXTKibneeBAlB2xb6wW7IKRy9+GkbzgcaywW44i72NA
V1Wt0s5U0T8Jy+FJtJxSlVvM0ZB5hAhEFEAD8Zr+oVgTexQ4v5u2DhI3/YBGHuzF
BH7NtT03ab0GkWMLQZ5n2/yRq2IwfruSjYpYoAKuxBqi0/rOSQElN/+nfHZGHOKd
TX5wKdQjOvfSK1tlofI+JGgwKd1C9wSOO0fDDPGElJtjPNopUAX1oC624qm7b4Ke
83JxwnaPSzco+LDrzYpK29hCSiZU0+s0LjDMjQmTyA9pNXTRFVSDlNeFJrSEXWnR
l0SSe5j/oDuc9NqkQcOsjfSIdIr5iWxgHSCstJjr/gVPLVG6njdS0wH6ZFVabsDc
0tAlSVM78XPYY51S1vidhwOX4zaujkfNW5BCSm8Il5IN/pMZbv+0CKjasLMI10Gu
jWh3pp3Yc0E9F4yiQiWZdK52R7aWhW9vRB1l9Eu05FztzMMoxvfqJZgvwRyZrYLc
3XsNF7X+9bna5SwXjc+cllQ+I1g2xwvG/E6lf4lQT1bUrMGOokIhJZuKeKMl5MAa
urG1KqB3vocDIXshblJT4SmGnAW00O75/hDkzbwO4Uofy+dWa0/M4GcGeo+0lk+H
fjjwEhKK4hTHxcbEEgpJXGmIyeIi02k1/WN/ht/IaeGMu3wK5PpE5nqip3oKrDLD
ZUhk1cJtwSDJv3VbvMxmPT2mOEdkAEjnJAhTftDgElz2QCnhx36hMibW7dPu0zon
X8ZxFhI95LpruvOoosBAYTFMmDcd2gNkiCMp/m/kPw2o9g6UqB+ijuAenddp5R3D
W1qeZKffV0f/7NBHeyF4zh+ny1SOxH4Xfx81UzBr9WNwswmp4K0MBpPWm6pasDVD
HQ7HRB6iDazaRYD95RFxvM4Vc2Y6lgJ8VvoZikzLAM+vLnqRTVMg8rwBovtkmozP
BWIZQJDxkfFZ8PGVkG2WrI3DztHxJU2sZSZJmwSNcvEsh+zi3pd1V9bg5OaA9nyf
7/5nALhaz14CkDIpKmsi6zgJ8VwxuZ5/brWGTwRvp017IVTMno4fRz/aeVG/z2mQ
w4zlvqSdAF15gSY632SMeS1NW+b/s89mW2KJLSYwxNOGZ17QpbNXVSjdlZgEelS+
wYHpemRisANizz6B5FzW3qzlamgZUDfEDq+sA0Qcsv+x59aSdBMT3L7WAbX3aWbx
qhQVBQZ6eU7VBoiuk7xuur/FluaZWBlLH17qpy4Wl9qavVp4F15N1jOegv7bcuvA
gLo1EInQ3uGX2k7AIX3puRPGgPLgOGctb+bmhUPSMZOYl2BMYYBUqx+h7MCY7u7E
YzWuxk/LTiCbR/9Rs2gPLB8o86BmCHBeNeRdAkKLKRJ1H8eb2ZTK7JLsmrkcEklC
WCLD3uR7mW7H9pvZSb+Z2uvN8ccaa/e7PqHoSsbDFXvazUsSDt2/mzfD5BLg9Q6B
RFgebYbogqD5tELOdhHczd5rqVPciqSOlMIqDNCHw4M/OIXwWMvycU5ypbHKWgRh
z1MjDsI+A9iJ4m/4+bqUfmfRp76svCrNSIJVlb8PHIOG19ldcoZc1bkQpsCFBKUJ
S+FZiQbZ02cdvfT6Xaf5RLXd0T68TgiwB5AI+L4Lz96oJYR893DRVVxnVSWhbb3u
Tpp1gBLbDwD/KBEDCwxRmAriCFvqfXqkmEgrFStnGhaApxPgylOsc7hA5E2KuJ/M
rsC617AuebKWWQDvv0eskCMGjbHNsaWoyUnEx3TSPQ0CDEA1lshCwDpCX5DTaI/q
II+b5RkKMdNZuqzsZunSF5Cc8ljzS/d7vXWAZZVB4JJExtwsBIY+59+XXtz60k63
a6WByE5pmTI2f/HaCGH/fslVWFPh4gZKC1o1w6lg28d0urZhQ1dtSQjuPXc/r0B8
KHvv1t061HHUECZZ3PKmzHQZjn+5MNWdX4L5zHJEOW0iTf7gvp8ijCnStiW55M/v
jdmjPC484dKjXU2Rt/+yzgexLi1uFFYehC1WS9jwTzbZCK6y2Ogk2ia+xhMgPZGc
iP//IpP2OBX0h0s6+tojrN3pvt3GxcZd7yqfM5oJ2mccCS19P95KD6rzRzIpp3eM
QShG3R0h9Iaacenyba6AtAK09P+NNRJUrDMT5GkiWJs2cTeXtlsRbKJPHURYQjxO
1pQJaHPhaK4KMIkeL0V1AtWMNrKCPH50sGqKoPKtnv6n6IP044DUzQV4ZjodhZ98
XZCrj3h/XJqLJBd8crAYUlzQUoQr38q2cIBriWZQXH8F9BfNQ14Wug4QoHZ4Vq1q
An1fPwM8BUWciZmcWg+JOo43tc2Fvsv3qBBxX+PS16h4AXuLbk8eh3I3OpN+z3w1
FK2b1Q4NRUEt5QuWyR/3sUF6+5wGaZWavr9q2C7Os1GB8eK9snrMvPyitx59DYUR
EtSxySjIdnOUUzQx8Nk0dYjt5Dbw7N8mpXQ8tpvmD9rsovOzkbZ9GC6mm8j5aMbV
nNQshGrJEF363TjqpoFad/0GRqHVIR9G8xGhmKnEusizS9RolWImTJTBDloFo908
eyz1vT+X7gPy5jBxqkeUFujjNhvIVtvVK725sjgeGQa1f/X9vbnzk7qfDsF3LWc2
hiF3/G6FmxYiYQYTXp6qLM4NK0WubGueCOajEnhAHVFoHbIdf0lvNqfVuzTO2Bje
erodIrblIjfd1XFoXw5/4IkMyA4jNIrcwx6XBtYaooq+ZYzOTBj491pKBCn1yOmJ
DQBt4KI/q5mkTME7/UTRUsprkb4R1WFk8WpB4j9zWOLsYKBMtZq21qYIA4b45/nl
grXvzixcXYp2kuI31d3ZficT58KmnpIl6UanLOSLU14OjtY8lAEye/gzj1Rppmni
rMra7NBMz4o+sLmUXTZN2fA9TTqZ/tRH/lfyQFtW/8SYEHgnYXXnoXF2IYWWNwFO
uKhQ/EFtomEJwL6sjPQcxWIi1toRVcaJ4C2cWwkax/N5yTAe196WrGgMiD0cYnYx
5NuGRFVURFUl3EWwlLIUW3rMWrN0dF5EU+WtZx39exDu44QwlQl8EoiHRCfqhR3K
6Xys7LXP4FmRaJ561HjJiNXGMvd/154/uK0bL8dohPsJGzlbMkUvJV/OBWlggzoX
kehzVsBdUzUNtxND4NhKSnvS79C2hgmP1XA7TBESca31Q2szRU4xhvAft4UwDZGn
JpAEPUkPdpUBDtrRUQDpSqaQsEC1M6++HYk4yX5ylK+k7+X8dWuPBxJyF4R5Js3j
45368QJtkt0c9unoJU9H2jhWS867NQh/hauDExd5vaTplHeKCzV8S0hyYepL3IiX
OyYp66qxy9i3oSn3AYO5HJiqkfMyPz1cTOJa3BKAlk8Z18VToJK/UQyqDGhE67/5
yinu9kxN/vo7ZK9K9c/FRCOP1eLfQXeB8BSfnL9UrLRwmRL8LWPhJUBPzhkvlZnc
LkqFKKTbREyx1wW0g9uClnCOdBryPNEgLgK1his9iNgr5Fyei79DG/z1ccXlaXRT
53aR08BFnsLh1atHjUIewd3aMqNFORzk2WrU0JEibXmPHHpATVxUizMgVaAe59eL
A//RMbv6fWxGYWyxNoGe6d93WUKgDJEY18wbFJvQB6zyIOs5ytZCnyRroQQhtZcF
jPnlQ6svw1WyV652XyMQUMKk1YlFBT3bQqPTCpz0/5hiZIKras2SlIiETzitVaNx
0IXjyJ9/v38MhHmwjnGJfUhcVN1E87H+GVfGwxc93sUk64tIIu1CSaaGmkT4FM+Q
q+WrpAOMqrwK7eev8aBidWABWEcwKygoBdVEKe/45NJmmxejSdKOSJXrRF2PEbsD
XIb//58bpeGmpfrnMqKzYlipioHYK1R63liHSpqZZHrwoqDQ3NILdW4CUgOsIyZo
Dvayksb68DrqUEwt4feI7b0349nuRQMyP7YlyOhpbwytzQkylyPuYsuhFfTP9I3+
CezL+8dVZ7mHudBOBoYz2D/fqnCguoM4+qQH1XoHO1cVSVMr3MCmhAXsYYf/lmUI
Hd7c/XjY+f0reUxY6XVrARfpSRH0kx98ZZ/yqY6NHoOYcnnsze21HIstPmf4+hKJ
73ZxPhSi3hbSSGFqi/vPqTK4DzN8fd4LpzNCwOhZM7+uCgnQkyeDMzyTJ30IbZex
fFeY5LxKIBrT2o4dZadaqMrgQg0SKJZEEA+96lufWWIn+9q6wB6pwpT/xeC/I0m6
iFTdUpuU6Kq4ttk7BhNSz4e7AyRHCI4UKwvk/XtFAD1zdrvLTn+HIN32Lfc7jSIB
9jI8gLbIJ3lix+HMVwFO6orEKtGffIFvn6E85hiPj/+38auOW50U8lCt3caP9D9C
Yey1pR8bTcJWmwt35uY+uWmBO0YYBSljhsypv/FFCBWdAn2YsXWvQiUOQB7ESi40
1RwNvrND2AG0JTFWXWrJGXdgXIwXFoXjkVcngr5asyPT9HcQrV5rzzcyYkWOLjHO
1x1T+1uFir5OG4ZZF88s01JOX9dlWkSY1xaSAzJpJHnkMO/RmRVzrdZWevW5D+zE
Y801mypLylBA0sEVf0pfJERLyYzu9q16QOCek6MoGxeRaehNc0eF6+iR7AQ1HEDo
bOS5WWHjsNeu1vMXknQLX54PKpIjSd+kwy5Ymd/9w3uN9VuOHNR9Xp6xJKCt5rI7
ZpUv46hWD4ovelQCDOLM1PkQ9ljen3I54EEKxRZa0khMOMyrufdetsmkgQGy96gk
Y+Rfk9OiXNJk/KGWFcRvdPivd2KEKxXwQSCGX6KciAgiAcrnspAS4Xlf0+/VHULD
GPos3hf9sUBm+foJiolzpVjD3Zyc47j8GJ3WLzsLPSNUCPgy2O0b6qU6jqFIZO+P
eFR4nQE62ygLeXDmBrDzY10JxlZ5D80sPvdtR/eyT6NXZ5oG/8N49fzavFKoQgbn
ipBn7uocB4OwRyt+bnb+r8T9vrwQPhCt00bMKpfMq6wBy3MCC9jAqrnm9BNhBWm4
iuKYgWcrHm/blJ5ty56G4lTc3bJkig5ea4SXH6l8rm/NOavQDXCA+U3y08a4Qlyb
HkzrzeEl34udffHKqsUyybshvkKR3InormoLOt+YRb4CrfjILMoBlHVd69/pPnyE
duZgjrgUiuOVgcr0Hu1OXTIw4uf0kytTpDlhhKEKZw8sBkpv8TmwhaiQU/iY5aku
R3nWUk0SDYWpLApGX6tbhieB2GjoXHdGa0XWpsFFLkxWcXDihN4sprHRlqAD6yML
V/bvWtPWgolrGS6A2HKM2h7Tw4pTc3bV8eq30DS9yibVFPi4/43ZqWTaI4ViB3bT
I/f4aMb3bGcqCEK++jFllGMTY54GwW+I3lrxO/89nNH8Y4TQrhhAga108VFPPp8k
exFb8AlMmb0HNTK+pZD1WvIUrFpxJ6ZSrShKYlbLmxS8CgAzMWVu7UvjtybS+DPL
ABb0ZgKM8wfcCLvtALoZGS68UB8PB//VSHTyiRpEMiv8iIAHnyXZLOZvNE9mYJpE
yK972BKMWSRb4taD4AtLM6/kC/pDSZKM85VkeCCHYi5O5RDZgnUKbGEkOgZK4/S4
cAgYQ4M2F/yg2Pg/OWLv7I3L/CET7gjiCXP1rfJ52j3Igxmlz4EVHIwL+mbtKK1t
AqUwjkwsN3+0IuC6uXnTIKGvSIKfnL5EeJ0ZQrW7bYtnVqu6J7+lMjnNW9u5xRM2
nRHvbMFTwc+5WgiWyAOX9abF9JJSbbaj+3ClSikWDmTQd9TLSbiRRDvYjgwgwISH
4YzNjiyb5Tql9CA5MRdx3TZPTFnVp9HWe2/NFO7EDg3GjLoWuaVeMC3vRO0RO+vV
G++yzOmv6hha2ZsA0xY+fJjfN50E/q2v+36cHnM7aB4+BOWnXqs1XEu6BCzc+4By
TJUyWOQA3OezHlBt2rhxdjoU0Es/CxFDJq3HrcJYGNZc/OtqjuRGQbCqMjOEGKqx
D9URWwFqmJX1D10lJa+0ZJSo+tnxvhR6PgHpRRHXmOfkavWzNExIilCq2s4ZLI9H
e40oVJSEqq/ugXN0ZxPcCLh5Nf2UYQIJ3Btq7sRJpbBZSaYXFeHKPJkV0W+ba6Ho
JzK8obSbyicxCNNVHfky0AhkQnbPCDyLsEiqvaJmmkZNnAGLhixsEahYtjFA7UE6
PFr+IP9XyjrNEVWJF1IrMyTBzeVU2LNAHRfIp2rg579HNWI+g4HEx33yWzNlNoCP
8LyafjqYBEqoTODVsIQYNaUg5RaOydkj19WNe9sWsRTxQ0nXkzryf8+MF0zBfDIN
h4dlcJugMjoK9LI6NCedkQNmLp1up5mhfsEzeJYUx4TWRJq9HnUMxrP8mvjCkeBz
njoBPUbvu8HboiwhbVxPbeFXXLPjPB5JIEoUEX1vzJAddSST36Xzveb/d8dNRs+9
flVdm9S90jwF7lY91XHmqTpoS8+adkDbxTn3P1XlcPrw7OoN8QHG6wsFn8qXrRgg
z4ZhsF7eHX0JPdSIlcKWFQg140s6qtLkJnr8Zbj4tGo3zLcc0BQ5YTRKHVMhhpKG
qAp0iF/qZchqe/SVdFXT+bzzCEK5ZH/1FFXxnSWx4WK6FDVap1VztV+yN6x9NiTF
KH/7Jh2erVkl9XnnqWbzhCRdwGH33uqJRqp2iGQso7G9XZMchEnf2Zb7q3iiOfWq
Lhme+pkOjXUsFduEbeJTylqVWaaaSmoW1etszGU2+DQh5/uItsPSkgM4+BIHy7sc
xCXIkn45sqc8NOZIgX3D/0LhteEYNJBq3nqZVTm6sRZL/+Arfls4I6C+9YSYVh8J
LguVAg3rV8u2Jb7OCFozwNMgZicbIoK1dvVgW7aLZneAhBtRSfjm7yp8ArK1lOW2
MlMEnT6fZNrd+F8ijDGTPbq0r3bg3x8G8xH4JSGuvZdsLR6r4Hk7q7wA5EqGKzwa
sbAKq0rbQSaKNKzLxn6xF8qQaA8joqvbG7NNXnCn7QASceUuk0/f8Owb8GW3vebC
s9ZUDo13T/60KaEipJzMvrV9buKLSn4Ki3NfaW3Jd3dT14fFKiIqqtUf4cgE9f5B
AecLJo9lSN7pRSEugGjqFy7R8j42FN/PomHJPK+ihKAPuktNrHdxhwnr6mA8Vye1
ASmMlKHAcUdEg3v2diIjBz+hA1LeaLIb+i0IZ1+3MRvvmCnRzYGygWJLR5V5ugVv
iCN282mpGUM/fvm10JuIJGD/o36KykI6IyBmqPOpORccpP45ROWUZaixC1GkDhhc
uXUKpMmW30wP6n3ZYOq9dSU99PjcyGFukzf5eVIJxik4QPzpk21s317oj0+4U8Mp
LMOBVfEO5mu+/AzoceuASBQjo0M5HvtpwfNUfNHvfnlnCYi1bpxd41sOTe5QhTXY
7bceh6/ZwecyAwe8C0v8qQUXXL0EGHunDyH9uJuTPlIX1n1D6Hv2zoo8E8m+DXf+
d8UlyJNPKbpuVkE3BOI9AUCnAZ58ft4K9ugeVR/MH4ti7sPVXK5k7IVWP3RQVUjL
7ZiSQ2sd26Ilt3UOdIRN+IthIRkmRYihK4IX3DZOs4ml/W+PcN3Ogct+oNiXD6/R
6HWBoDDih3KdujgsdADaLAjyAG7mDjtb1Uzhjswb2GbEXPkkCvMmV3SEx8ssE6QN
BTtuGLXOwcqw/718Tu+KvGdhyqkyeWgExaJhcXu9ZKPEO3VGQ6eD7wYYlZOoffeV
5JfjmuJqgQSusoSADYg6w8bMZ3eHAB4ITHua7LhS53gwdIEDbP86jgYs7ssSrlHQ
XsapA1/lCK3fQVLVmaR5qzH+m3VAZdcuMRrlwf8WWNnpcfdnUhGpPKxMbECRko5d
xyNUHuSgk7yI5qnPgHxuwjA1gyuyyRprJ/9rxBuCNb0bkK7nwAiE6zkopvE4oMn8
AIB+UsM8TeBk5udJKro4rcsPgwKoSAtMRLjuXQMx5SABQUOUlV0J/pNt7a5fDmTS
mTzR5iqQvf6QYYl+S/nECVSKwFUJBzFyXFw3LcLQHmtqLJi5lo2rTPgAw0SL/1MO
YGtHS7LgdvmOcHJNx+zpzhkF0VlWx/A5fL7LJuTj8lit/HaLcc6uJItr5xPib6nO
PkxFRDF3J89KL1E/sJ8wbi9PRpy3UzDyMHjf5SBVTmZg/XmnJE0yxuIVhJ78W26m
EIxDgE0cfXkhjYuzf43nxWEZNNDUt3uLEzBt5Xbf4N+1IyN5aZDdWnYCAjkZ7g+Z
g6QLAYi3Dg9edEq0EoRtxldG+FwY0+LVFiy+Brz48JTQtxrxzoKA1F56sKSYZAHA
t+eZ6/3vtjP8UuO4G4GRsDHFPYhWjqKfk5pmck8rk1wg2p0oypl4pFmBC7XumDs6
iPFiAgbI3l8vdHGWI+JkLNti9N0n0DTiOf6uOfxKlhYWNE5irm4iSpgaRo3a7oov
qeQkD0Budnff3Ve462oN1AYR0fEl2VQ8oHkKGXR/huFRftqvbvToVp5DiK+2/Tob
HjYOnpLv9f0ckgvdUlg8vWvpf/+kffnxTI7wSXkt4Eodxdwl8/VPCgcilkI5KoAW
cv0auJ0mTr3Bw69iLtgoFnjm8XgDYSwiLAT6lIEOfAsKiR5vwnA12LAzZ9A9VGPn
nO9uKtIabsdjqzZxGl2G931sg9y0AQQoIJ8W2uJWth0c4+HQY6jCxlsuwSgHO3z0
PJDLsUR5IRHbtQ/fYV6dAYH4IZnEs/nrxtsZXMzjXXhJSEhqx5Yn4RsgRnN5l+cm
xjcjZlI+2BjSDyOfaKwVf18svmeJOfYbTy7lsHAt8RGkptBqrq2yZHplNspAVBWC
vWxzFF+3jiaZP/7KgszNqz2cC5kekr3Kvqx5lbZLTX9ht1HSez0bUlA10SKnsoqW
tatYCAE2LBVt2uSe452joXvujamerTKkeanM43og73IkABo8UFpubpEgl5JuogKz
MrjVhTUOtSv8Xoajvg9kFURP1YJFs9N7FriX9bdq6LuYZCWKdBg3f92WCkOmaLY/
m0aJdwG35gmkWF8swowqHnF+o9OyhnOdfcCTna1AfTopOLxA9Nv+lfRKWBp88jnb
bZh9teo0OigyRWXuOEldGEdU0UVI/lVFRPHA8HNXTImUW0iLwZm+rwfAB/NqR3lQ
As3G27W0Oxu1WT0WUpw1uWLtlcbMfQENQpyhp0Etd1aNbjojqf+Cy4PjrrBvySP3
RKn0U5uVbuVys2o1KhcRpbAV40v/hs05V1KSACxeLUn6AOaD98YB2QvdwN2IlhEL
Z9rzisOarTjhjf7BMq7V/YJ4zR/GBZHn8wvpZoTjsyJYIPeiW9SdpxlpL6JU2dih
QJaVUmqYdsO9wYNGZ0RiTsNJcoszy0V2+es2YtksogeppHDsmvgvW0U7wqHgKAu5
LhpMjgSBq3oN34PNy4znTAru/HLP4lbahXGw1zwMHDZYRBH7e3tLJv0b/wDsuF4o
ZkZnWw8RYC64vIOnSRPGZVwkzjyM51/6VwSlWp12qkxf46YV3At4jcwFtFIBF1/N
CAbTTLBwxK5lU4CA1pqTb26dUKIIOrjPiH1v4Cbk9obXJeg0TIyDvdIw7K75dm7I
Nxip43CXnZeC3rbnpId5i4HuKiY44015QB+o+smwRLoa6ChFKBJa9fC+P7ALjT3h
S9dX46pxmvA/5ZP4VsRNXAsyPvDvKLXVnriruJ3ii6Sm2ob0EH1Ch9PHZI4t62Mh
y9CBY/TquijeFMMhpO+jxlrx4pnwGm+BaQ8dlzqWfjRr2tv1rnzJXq8t84l4BroT
2Rl7vG2WRturRv7APbCQkgkRqEBHpPPTK/OGL7Nc32Me3cRYjKsrYPNj1o8RXDtw
iUp7uxro0v3M+somwTEy3Gih+avbj8WIj5/yqCbEV1WwtvcIu3/NJIevK0jivrNJ
x3EfduRsHXVK17dtIVdKXew9jlSyfCfyXgpBN5xVsmJITPiOE4/30TAzynaAT9DS
a1UOzES1PH6YTZTJDfXxgG9ziqT331YEh+uVbFEr0cby4F2tRtdKSj+GMa/lbR8l
WH7lYGefHmSASSC3AxYObw8VDb8ac7iI/E4mXMaEMTn6JTiID7e+Xbgce9ZV4E8S
q4tiOKPsuPWZSjy/sWU9UBNn4CdMIoP6MeEkKMrnM+FghX/SFljTZbAa3oejK/e4
JzNTdRA7Z4TooQZKGhi1014b657LoEgpDVXNOwO9RfWBhC0epJfTK8n3TOAfpVZC
Z2kapTgpWHiCAjbPDCF3ArivGzl5uZy+sjq/KGxNcO/aDB8y4xQBpohkgWqVkBAf
Lt4Hsn2mAmScIfeOWblIn+/CJUmLPaw4l9plTxwxDMR3psuXXrGtfSBaBe2e2bk8
HdMxi0bcJ0UkCg2aPc8e7sfUtvEXWSbfCgp+NvU0tv9lxhpKZtjwhYUJuRn4z/Qa
6W5XS3C8IAP7YBkqYaGGWf+hdWTNDbCf9+i0bHbzKdIWKP1Okng/8jTKdoWTfU6j
yXOS98Q1dK/g5WQFt8t6tja1j5+iKsUfy44NYgxL1c0zy/six48hO8I4mk4Nu4S3
jaHs4urRfoPZY3lWOlU38Ow9EeDRRmwf/kHWANqJ5qhdbH698s6K1gtowmqMXflh
amnfaGeya/U7Cq+E4ob3rgLjSQ5Y4ftvRqObdqNsreehsozmskg8aTLrS6SYQFcw
+5C8V6m4qCshk1q2Tu5gNbqy8Ehm9w4y+ncMEH/yEwnpb3oN6DDKTGSvtlQ3VZIt
l73APnWSk4mHGnxbVFuT7sncKCGF9onn8pIGb/VjBmibUt9dFSU/Px3fCdKhyoEg
Y1HxJl34RLaBprGyf0dEABpzyPdM4hE6nYdwHXGgE1UCbqxmJsxMLkhyB16S3/uS
CtdzK11P3IEEfYlLfSluzetrWg1p/ckHeibitWy5SX3qr3iBCUxytlQIrR4mQRsV
40ofc+NV6JszNxDUaAY7cWAmheeiy8DsZ9kEGoETWCbPBgSA6pn9Mn4ulINlqTpN
U2JMuId4eHi620xB8ajyuzQtiO5Y0xE/M+cyuceEwjxgkf1h8us9TQajemMCNlmq
cyE0kcGWfZUkqcQH6ZmDxPr7x5z9Ol7YWHtXZzd4qSidoKqyi6UFWVCbdstzxRLi
IQ8DgHgIs08vQ/tEd/Q2+tzglT5a4hUXAQv4MqETmiYpHiWvn+YsKDRQ8zk3EeDd
CJ3Sd4DdlHfC/bGUNH0sxHf7O0iRaFtQb4FxXXvR/rLADWDkr0lGC167HXDZSGVl
p8p+e+RwbFYyDAaRXjYtXssgBzoR2r5HUlc/gCShUP+xwBG7fTseoK/JQtc/L10h
jxBBH+QTLKyJOQoCwaaiZ9yA2NuWqGsgKugeJXKsJEk0ICq7GnJbPwvBhcEA24jQ
WZHzGVKZqS0ykvmXDa3npm6A4nkCd4LNu1o0Ync2RfDPnJho8xmFf0NEokMh8mk8
sZVOSadz1LfPgJw4RJJTTphFmxRhWCCzz+XMJ0Rraqk18o9ttKfvgs0aJ4i9NzL4
K6tlqnMk3zEb1+Oib7DPB0+0B7ktmYRLTYI9h2ap3Dk+XgOiFtpHwllY4YCB3aPY
KPMgo5T7y5RgiP51bxOzzpr7BnPsoxiNI4QOS0XO3SSZ5QTJPvZojqHqvRsSWCt4
n3jfqO+RDc1Mq2gW+Ykj5rjhw5482oZgkeUDyXYw8J3eo0z8I8iW4DQiiyCZcylL
LWX7I0+FqOZW7C+adaSOaqEaunGxY9B7HK0lFWPR6nNSkI8rW/zqzjbVL4JIoceN
msk2fypbU/B0i1fyvMvzLvdxZGTrEFPmF1wpw/vwwpl/yRxuXFTOI7CUhhkXgTmL
tw0ZwgFewTf+8eaeIqhP3miWe3eWPWgYl4k1n2hf9lH8WN7tNTeMipM6Q2B6CT9a
hCCNBYQAZs30KpZ30528K0M0J9NDSLyLMfoxW4yzs/NIKT9knTxjkP+pWg06kxtF
LV6dbpyWl2cIV5nKzvQVCoICZu0YgTEiF3f8YEo3K6rPXsvGT0gFdsp2RDQBg9HB
ME750b00KzAicUk00JllJ+0bGACz/+JrxCSG7xc/GqWrm20KcM2d3p/0kA7MgggN
/2N3HrTeHES4CgLE7SmCFigLccxcZ69x23S/4iewAGYONH+B8KzBBEMgeOpiQiBU
uZf+W9saS4kEwNpYZzrHusBctie7ntShuO/wkr27q/wyaftCskb6QWaWWn3EAAsq
s2hILNejz8cMO5QNtMBggyEk4wCWxnBB2DfsZf12fFsasuT7v/ND57pFiWKrphG9
lnjPPYE7ahm9WDKhUifuA66ScAaCGloZanaHQ4rRTiHQAif4V373UGGHu/GF6sBT
67Cvq83Vj+7hpYR4TdvWd4LC8MIl2dL29HxDW6R+PeApAuW5a2okKoUwjY9Tj/Fw
LY8x1Kwtu+0q/MixNBQs0TTqIZnyqRDkF4mbPdmwx0kVvaDS+R2oZOu7GJMl+2LO
IKK/1Ur5onZl4M0Sn5LQwkl+eqDsUuYimsq/bN9qzZpqG7c9AvQaDohiCaKpumMV
X/gfcF6SWeicQG8hRAp5DHH3jT64c2mMWxqTp8MEPrl5GTrZ3fDRfsCX9zSsssK4
Ds8rUq6gNVyo7aMk34USMWOw9p0eSBJP9od1IBFsbKJImypoC9J1nM7l003PIUrL
KEfbeWmdcHBWI7DS6JUzz/OorEAcR9Q05HG4vB8ZbTxSlRjDsNzAseVD2qJpohnD
YAzHsu2ztiXKekcqiQ1xZaIPZhtkotkEW4RaxwUKtvdoRw8dces7MDHPYjyNf/m7
fmz/tcDxx9t7JmK6LcpqLL/GznH5OXuxy6+HRQsucu5qucnvknkTxcO8K/1RUyoi
bUhWDAx0dwJ2O3x0eifAea+fl6+YmZkj4MUPk+3iiCA+nsiXEY1iHObCi2OGFAMr
hHBXEnKE+jAADFjqVwspBN4/SWTIvuvdxSo6wxYRnbvcMOd5cyevybLtE4dUNSfV
tI3V2MrLvyoP6tEAnQdBt0RReZr63gOxUCznIOt6iOdiHDY0jD0ZDyzo+5IkBDuu
SdVBSP718AM9ED7mM66s503hqPaLE9G4WI5ZGMH+vXmhCtSq0ZzYA9vNjN9iuqvF
gfHnIRkjUvUs2fBgmhFxFst4nt9qDgiNfHTJkCimdlUgG3s/WiiR0M9q9ltiUmbp
BTF8Lldqno2QHRT2T+YMAmh7ARtzsF+1y+5l0Q+NGV4S1NGyEywWgCvN9t5YW6Jw
hZN3D/EZHzrvLftLCWMT8V8toU4f6yYa+ZeCMNMXqvUAhHnfBIzz7Ob0+1/0bQhJ
Lhl22+ecZEdPEJB0m2LkgYJ0nF/dnCV16rTeWHktb+aFzCp0rId+2GEH9zx0QRjU
6F6VAGHkh2HWEOLGrgoW7SoUmkCVvC9pHI+AqjzJV3DdGflMCoBbIS8Sm4UQPHc+
SFlPk6iEjSNIK4qJ/Xxo8H5Em9zgNMuQo+xNSbbQWFJQuY6uXdCeKhpxaAKoDdHg
6SS3xwlBIU5zO6AOZCWNT5rXKNCHwFLHJvreBfXh7B4cSzPiGzIi+WiDBbvDJzTL
r/2UjiSC3n1cnsFXqOd0R1NhKzgyXm231E6khiB7kUowU5HPs8sl0tktDzBnr0Ll
uaA7ro2aquPf+Jn65zYGuvkK/R8oMxvLnZzWqt2iLPCBjQ84uB+lurFvurYKPSWm
llfL+nt+OK8bvNHaux5GnbtPXFlIUHVzmY4Ng1eradhMBas3nx6chR7CrS0BCY5Y
lRNV+8CgRgHihPwOIrLq52vXyTd8rspB6IopctnAzcDdSeoqrd4QqvyQSjKRRcgV
8MieK5CcEnTDuH+sUB+kcaOvzcbaBhYyYZFjl/Agj2Udkx6f9/NBFMatpyRSL7V8
KPRD66u7jj0QAgUEPpC7lQ5D6OV/FpErRob/JTEVoIQK+wi5AUWeawePTP+pHNIs
S1RK7pT/5Iga0Pgf1TC8MKQwSE+uJWHEqYhRmG1PzfjIG6AbDpbd73ASXdguzc+/
Ghwm1YD4Kwjds4AKCQdF4HdmzRy2NCE8+aQeXI3Nu9kZLj3cVXmtHCM1Or4Dt8Ba
5WqewiX18xX/1T07dT4yN9lFvFr3aV0t39ua2OxykaihuYHoWiku4/IekXK52dRL
Zpq7NL+TTAouN4gQ5k5+GYiJSTAO1l912MhHvFxA4f4LDnikdlsrrL5STvgvBZSi
EHI7ZuxhRRvfGApIwFkQC1c67y4kPn4HzPxjzF71yF6780pjYsiaQ2fBCgJNB35t
FlIo35hTgMouk1X1cZaL5LgbyIfEEKCfxL0fJrajd8LmRZdLcXeqtLRZN9hqZopX
Trs8oAbM9cwSnWXaCcmNq/jlPzkd74bvZMA+ShbEsjZDB6wrQxbMtePUVDg8qPrn
9lVOiN9tFAtEGgWkKkwc0nn5OrGT8aU/juQcg4J2rVdx2plyJKYE6i9KnQ66Csnu
99ErwzdqBz+7Us6MoRx1pP7DS5dbuN1GD7YpMcptY6wo1r2k7fdwPPBwoGtjFGOY
DqRBH0r/HS6Wwra08xL+v1Kb8SXbWpPV66p7d8AReerkhtoJ11pLOdHYkOO4urnW
FdyUfK3o3zrxPcMcaA6WaCk5emSgcGiiIyOHY0OgNjF3eBshsnRlnMMPj5QmSHFy
2NLashw4Ta6MVQkhzLJCwMs/pi1T15J52L/LYNZd/XcLbO3YTLRnCbXUlVXTNBQV
zw+o+h1debPoW8vuTir0EyxJccMHivKz/TqjVIp+2flGEIV+SeSYLkSt4TEYZKrn
lN5F8L2O/q4XdgGORNOWq42uS1ztoHdC4UjifSSWWqTuHMq7ZDAyYEi3ZJ3/kWuu
IRmBmr+GGQeiNIvpX1Ibm1Ih5M3Jvs44QJ36827V6A0jiXacB/HCp86l9FWCDPur
bxjeyOMHZlRHWhTKxMan8sPkYi5tLcPWD64LzAi8KXjGuLacnzEi8ckQil1AvSQP
YORC8Gu6JBveXy6JocgKOkBP700+865Rso4+Hd5xQ5shKCWeoPfU5BRu2YrGmflq
FU6wAoYjcbeol1yIDvDBA4/9tkPTKChmuv/059WL7Nb/y1r43hwYdKx2hZDELbfZ
8dpayuAyBJg2tK8iyj/tWi/23ypXOzAehhFyrSRAZHDZoARJqdY0ZyTbqqYdB0ky
kuJ6W9zaexd17oYD/dNDrop5O4tEZmN636ENwWrhvhhqtn8B9Fxcq5nbEISsJ/Dr
TNRabC5Lw6JNO7tCxMalC0iFGNmaYrXn/r4SFfgBoKpmUSaaDLq4h+4bmJJv0nFw
4A24NKCg600bfIIi6dE49scONsmoMtCp3tR+XTfGigls2u0GtZ9GheGI6fdf/e2r
kB6x1Dnn00mOrFbfjuMaTBNJwCmFwhAe5kQOV95xzgxuitTtYjo9jZjrWPVh/ayp
NoWPVYEUBMNqC3dWuTKIWZB0655DuTxdquLhE1NlndhxMCjQmWAay7cycWAx4qON
onLfIzecAMT2S7CCW49OHx/WnlVPe+cA+heHuB/uqeeNYA6jkHtDtADSVYd5nMTZ
slqy0wP5kJbsvUYt19nRrkuIJBRWnV3SNMEgy8Zp0dgWNCeebesRVdHGGrCfC5qe
gxQgYI7JytLbqjzFE1OZoLydRA05VNS0g32CN/eDEJ5whMR3vAUeREVdb5mWcZll
v4R5y5Da3I6IStpWituNndhPC5kJykKiyuD2PcIH5sQ6xLbJA8IREH0/RhXIYP9N
D21sqnP+3KAvSg1qLGJnJ2RjRsKx4obOAy/Y2cnM488if1EkxBQtpAB57RM7GJ7g
3XPlDF+CTNKOtJjbs3MkUvzDhpXFvcVLvpaJ0R7ybh2KiBSQj3pxKNJaCmoF9Kau
Bo9ugHsVQmkHaBzooglC+caYAhuYdt6dhmjwxvJEizZZWH2mIzmK3UU5GLFdGcks
SAaIEONl/QvRSxmfr5qKHBcLBytV8yvL3+arOiSKrmVStK66TM96e/bFCi49BINT
gCstvK1CQr5SIMKkkkp7k+IfyroMg1i6zjU7OdeMiZ90nnkZjviM9wJ8PwBQ0c/Z
NaGK9RbvbDRoD6w4VnPWvwxD0fSup2teKV+yYGbNpBkY89XTZ9SjXqTZmRW5Bsm5
q1XF+xPUn7PDmtrTWArDJknrCEFAA1DSYFGGX5rSItC8wN4rf1HX/UqOSV+cLuKg
LMTuO+byv5+WLiqFyvQXOR/yhxKXU1ViSBPfFF7mNAn/QMBPqaTQ4peqS19kpjGU
YHJCyF+P2zdIvstfODu8Rhl/hCpD0FcLn50h5PaQaPgV0ZszP0EHJVfH31eRUl9h
QjvUVXalfKsdzSchqpGQAaTbNhS08AC+azf0x+WWElPcxlwyJVuZDx2pPVst/SZp
yp3/U+Xylu44O/sUKbWo+lhNwpuMYYoooxKv9qsvfQcC+0GgO4yej+yyhUju4vPA
cDK2d1dYPcvZgqdZOuk/w+w9nQ3diIKSUR85z1Z+zzhNdRlvHAZsYJ+ePvXW9Oc3
u0cxhpNgGq6d8O5pmgFKcV2FMnT/5ZdlT53cfUbH2ASSlLZQzgTR6cow7FcmSuzn
K8G0luP49K8lpkXXTtsBTz/R6n40eE4bcEP17dS9TeN29npvlEq3GoEWaf2eU0VW
98xg7jgdaY+57AAt6VA44zo/j1aOF3OikPagxJrnjrcQqrfXVZ4dNP6uYaaOj+kj
BGfB4weZeNmk3oS20rZj3HJYOKNucJ2TFMKqRl+lhtT3Pq0mxC7bOMDM8lYmXspw
6cWH7VzOoK0aqOI6EVPrT4JTPCa4nH8LVmNJlSy7DNV+KYgTPjEcEXJ8hUeJNRJe
99yFmK3nWJSB4ql2LsiI/cDPQpUTUaePqWTemOTnY+upgaQ389HREDHpCPsi3N/q
aNpjexHHDq7wgqHmN8DfmomFYquJ99kOsf5oaGT/zvnH3zuh5D0sHTxdOwdk7440
YUWPRXGtqpMeRdhV3q9JTz2cCeCbnkWJ6pKGzBSJYSCA35xYrhU0BZIdwOunTgTH
7HSE8Fv8g+7ERVPzxMsZ0KzfQkFh7MlU4Z68hs/A9pXFTugwpyly7O4wS/E3an8T
03yCvHu+LhnQar8cA4KeTyDFe/7dHZCq9zs03AQ2vvmREG6i4FGYSA7QsFA0pFcK
gVCvfISmZpb7TsJ5p2bIz4tq5eKC9OFUeyPhnRTcz71akPds051s/zMuAPVQ7vS0
Pu6QtujPQCgz4YB5BOVfcWKm0+VkpaMxGeXmnVm88bQOmoRKGVAyf+DmhU4uM78+
OFYjYnkgHBbG7H/Gj7RPHHo+mGC5p9AhVaMcV5VKUGNHldY8s2PO9yxEgZ+lvbYW
65OJh+9tShD/sSNh+7M/yWfYwk/j4sgk6o5d3vJwvXaPXgbdnXnOi20EWAkGYorN
YZ/pODjo7+A8OlYVE/YVflXhibDS9+u/OL6BvyEdabdmsxY8TGGRJBh5ApVuavyO
Y+1ziJVXph7Lf64VChOd84+wEHAbK9Qk7UuRXZYSsUFJLk7G03zs/Du90xZhBmvy
2QgZUDA12N2otOaEjLLXDpVNQ/IhFBH3suIPkNigfoeq9LsgUvKMTBZRtzkjCn3+
CwE63xy807KKV4zdRwfp0tKmbsaioACxuE0n5l/SL2aGMLodORWkqqm8YHJdqV9N
KCzmDOv3IJ0cwMFEMiadJNtYXYZ52M441Xgz+hFb3QfPuR+7nE/O5p9qfm3CDs1Y
kEXmsPPyeCj4APrZCkwrd/cPHdw0cTqEwbIAmLzOqU2OH5QrCfJ1fzqnTo+E3RS2
Jscn2WmMWOYf7z0SBOeDcBiXyQPsFQI4HZaAn/M9R2EA2mNpGw0MdUz08E5imrep
GV4UghGLvDsQobaxS6h/eghulc4RIdZ9QLIc1vJ4hQFJNnZcLUWV/ZnMAgNrgscr
FTixUWYl3uwoPDuTs9TB0SYxSR/xK9ojZ+/Z9nWtWbBNg1kgiqcesk2MZLjAc7EL
yEVjxYefbwiPvre6P5op/UuDDCrZB797R5lxZttxh4dk/RSVGiTYrjWpInyOldFK
1NcIS0VQfXpUF1q/pSYRDJS0CUDX8KzyDwvBRjASBmEdlmkWJy8jJwe1LvOcdn3z
VR4rY1XbB4pdXz04/kRTf9ZAtqXKMpn2HtktjI6LyPjDAXYUpv8RLr5AloKPcgQG
1gSI4Yw1DQcwPlh/LY+EmZhZ07jZ0aebXi6yrzjC4ikWdzpj4RcJPzVxfCdznRUE
dZz4J8ZA9HIU642OGNId5txUyxg6+p2kwU70FpZsmsW7XzVcthTiMbxvIDVYL6Oo
YCuIpz/wfYsnU+GN0ORyakQhcyKBNfqVQ6rIQBxJEwdZDx0MYMtdVvwUsfpmWZqG
nHx6osnsJAiFEgvNiQYOkEizQSgKrP7mUbilC0874hhseJ4X3QoLnq0grzng7yQK
RFlHNDk+mrUi+yIyxYcIWBh9OSf7O7tSQisi+X4DYadjAtfCIm5Ry+LYQ1SJGJSr
d7bAdrR+ywHpGo5IE1UMSmqGjTL+ZqxNohjk71iiwpFmW6/N9ahrplYlvcHNC5DR
AYVAa4qjVEgX9fEFdju/fwCCE5LzV+PSkDmbJJbkKgfn1EPWiLkYf7CLtVvTh9CF
6OqGAsnNAlkdW8nXRU09bdz5NW0EKKfj7imR4IekotB/8W3ZfwKQ/FcAJqXI0zgK
DA3lylxpQqfal+Ce/5yq7o+7ulGzeeSf6ynhHRbog08sUm6ZCegXfBQU2cx6LVvG
`pragma protect end_protected
