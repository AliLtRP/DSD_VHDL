// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:19 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
kU8lr0d1jbDZPuwmEa/llsjuEyQYzIeR68ASp5GNabryljGGuyrccn3raBvGMxo0
bckDi3Ihngrb7hBedVD4IpCNZeGjiBWIjbtpEMvr9Zx42Ul5qyWF3sfRtKPPJSCz
mbE3+Ioi2UjvWPnkTVIBpqnw8fn8ec9BvELLXfjYF14=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 22736)
zBBIQ9zwvSQmJpEN2YkOYrLuxWhVlbH2L79FjKR9xFJ8xMDrDhjnHGd35RqBfmBn
V/3N40A4E9eAO3h3ztUARi7QyqL9utKj08Lwu/To8kV6nonl5jKpBJ95O8dn03Lg
0vnklfYqI8pz+81brYrvtckphxEJIHaiXN8fGBvKNj98U6myfc4bBb5KGi14oZXD
EjYEaKG2NyID+zUBN+/WUKyyTlOO2ZXvK8by15qt8/0tM51/NUPaLwqIq6ChAvSs
+V2Xff5ia6Jvs/Z/wWNXp0VuZwgSGdswfKD0wzt2pVEIcf7A46DWYzCH6JiqFGdE
JOHFbQG2Vnem4CPgt7lVGwYxI1/EkmiQSFr0WzY6tCSS58Y4FhQcSOGM26p1CS2e
B2L7zHtFBYXiDhsYdH5v69yo1eQiNrOKSKXCQEEjfd+aM/4bHefLJCzS0QNVl4DL
mzdV+1CLJMbVvMJPeQ3SpEsRO1Ju9mg7EU2HFHFfOhHo0DRUZudLzRo2uMLyPBBm
amxBive8vAKtPnQtvcOXFZAqMzCjItlVLFhqKaFILffDro5cJpfRl/nxqiQYZhex
EOs+3zsLJlDZJXaLxDSkMSezFfDxlImLqLAozIRUfrsh7GurF2v5l/RUYZ9/pyJ6
M9BJN6qZkEHWy698GdmUV89vS+K5SjjS8GTFaYZZr4CsaZHsEM2riZwIaF3Nh0Ci
0v3EF074yRubFI0nmAdtG1KHP2KJzcoR7IcSPaFFGxh9I0+vKILuntVBHLkK5Mgr
rPe/59azX/EX989WFw58SJWI8zBl2vShLPnHffx2T7T9f/xYljCdMDM1YE6Mo9e6
LFYvExFPqwDRD7XGVQZRlQnZ0hEE3YVP5jlx3G2sVsbA8hxcop/l1peY091n0lBp
VtpZx17qoVLbzvwVeoiwU4BzBVkZDbjIaTF/36IbE0767VJ+7ANdAI7nmTqkAJud
yj0zyeRmw9xLU1ymlKIb/jyINedIn7oxFrd25jSaKppq0i/zSa3PDVKtWTOERXET
c1VpUwQgOS7iOnNiT2Vif9GQLhn8+UWZYG6vuRHQbNBRmi0j595FMttynIDpdG7n
SgSn3/G/iD8WeqvG0Bp0R4FXLjmxKbBOzJ05W/wDBgWmsD4sjYEX/dW6fk8NP4E/
HMFvsnw5lCurd++OZXr4jRz8+QSfGa8PE76VreWAYMp09/eWp7UGoLpo49fXylYF
JCB61/3pDHyDB4xTqsfKB1lO4u4tmBVAieo+wLVvT5csoZy3PlCse6JuwjUFXGG6
6oZIzqNtP9jIkTJ3kvjceE34weoudX3RgD1vJMu+gdYcgBojWTYdkGG/WRatcW+k
t80TDqqRHYMawpCMQtdyIF38lZaaSSQVhpQz3tVIspwGKCJBIlO+GcXL3RAT/ftd
8ozqluk7EsZZRv8tZG2EuDQi5u48PR71PNgaIuj2qnT/+95eIY+DswPHzn37zWlw
l+KQlqNBwKMXWXn0T2IgVGL8xpkXE7/id2G2TUILzgMBM1e7MWD+B8xkz3q4KrSY
vGbxu9LKFLbMwkk9IAB1/V5chThecukBy8EdTpiMuknfxeR3ZkR3szyz/cRGJGE4
IWEjsAhznbaKmfW9emluBUZuTvBdZxoZqUpOw3iHSGEAEEISrR7FVZQRfkhoPb1+
L4RGLTykuAM9Vr6u6c08hIQt/6cqrd1kvTaUFxwHbOi7gYdIjDTzpVRMo42Fohgo
CDe3ydGA63yU+y3McWln8KyrNFsvIbGUv0cJ+vfOEPKcMZnRQl4yF9bPkZFK51ik
CBWySTVQN5dP3JimF/t295lvkcpuQU9vGHY/z978FxRDvOfFxgET/ys/ZG1wTyRQ
tBfenw9Hy8GTr5ncWcR8Y5gtWmmKs9oWqAGn009CEq1tIIko+WCO6Fedn1xV52Lb
dGCrc5Y/JOeIwTQRgxUfpfNReJXzfeEthX4QEqLd3avFebNjnaNPhCr+vJyHpTvQ
dx6zFvhF7C4P1eDJhT/0oGowjz7lJLOIvYbjTSuhzK4nKYoMt8iGysXrT+dIXKIv
6dBC5FYeOicO45tgGoEfYYitJYNjLoP08GaChuRScSduvaNMY8qwXirA94YdRg8L
wf4Rx3Yfqf6SkOno71CGFH9qxxajDQ2mZ4cSdg51fjpov0A3D7WyPAke/ulPQvz9
MdPzPq84NHrhLL6PB3Qp2yvr83XXD+nzd/lmQymhg8u5W65pc2VocDFE1AfeDXTX
XD8zn3JIdovjZdRLHQCCSnyz9Z/YkzAlkTGikumfB2AQ8FzwYT4+vT1j8I01JQx+
MM1Iiam/VYBkSOm03XzNNlDm+6q+fv9cuig09sKAsSrpKEHAYKnm1G33ehqa1ivm
H8wKioC83IF9OjgSRzZIesF1pLxiorW7ni/XsqiqUTeaqWnC/+M7rx5o3CHDRcI8
H3AWBaV+0QL1sqt7zuppRA6aCsf/m7hYIDMgbmcYWvIw/kSuEEfjPKg5tVcWQzX5
WTWH2i0h6XYo/tQO4Wb6KzpnA1cnzGdQIUHGnEKRSIfxsQEmmKNKQxKffX3z5xT2
FRDyJnHhpNgn6l7wcqdhTzRyENZarEcDI75TMJirMEbuy7eu+MlHdjuCflHhosAD
osyd1SkE3+oITCom0A3rfH2FdBolSr3NN0QFEAuwG8KmOWnD/IX7GiKXnHDyZJwr
VjaAfSAhCx9YYOAQDDI9TK9T1HIaGDvQGRa1FC3RED0psdPJkfm6PW4DsIMVMOVI
e6aL26S/2m5BK3LPiU63oGuDLheq8zoTf+7n72p/JEGF4INdcTWbYl+WPj+0ixAt
AYqtRLHtjmmFRu3XUNyqm5Zf59VvYrnGJC+98Nn+629AhdI//2ErOBpHpS2+OUvW
6LLKBq1ybacnKdy7dvF7z8oTtHD/Wmc0zE9Q5mc1Qy0m542QOm6DQ+j94kzGJ4F1
0w1ax0qI60fB4F+2thL1eFHXHYbdKzxT5lQ6r2/Zr4DyYMfBTAdtojc/qqgA1ogc
4wQqMfIuGabh/iJN4aN4wTAGPI4D5ru2OL2BMJcdwjDOscpVviZEj9CHB2lP6lvL
Fnrl0NnZKpni56uOVZYPIE9qYqbfJ5ISwfyaZGK+cQaal/3uebMHtQpHeB6hFDbM
ZncelYT34IvZTbdXWD8CMrya1vPjv4DL91U4/8qVwm/l0Vicg9qpO9+HbhpLf/t2
WrjHdNqRaR2/1wGssKpaYYemC4zWopIbdeYFUbCthU8P1SuRKsjvH6NdkI/wks01
ZrO1gp6DpL1jDQ/7i4JbS1CeEZOOiHFSWn55+sePRmaF67SG+hbMOj90mPvGRErT
6nJYbx/B5Bjleea3N1TsgmPmy7Wr3EJemP9ZHaU/0Fdv3xCtMDaZUPXYuBptMLaG
J4loekktoRuQ2OVhN6WNA3+bb4ITrRu5EKMaqCGudKWGvQPwYVmaV0vuXWHch1Qn
i5GOdCYL9VWPZiVdoMPPB43+Hs47ESRUHl3/FCu4+w84ro/OXwWUA5NMfryOPygX
GYnUmUlNkJ7slczha7jdGKBa+u2C/LK2LJh/TnQ4HlWMmQOwySpx3Zqe23Psh3Uc
CqJSrK2UREie7o2uVp/TasnxDN/Wj+adctgw5kcZAvvi09PslcRfZKLhaxojT5py
7do7CL1LV7GkWaFdu2GQnd3VuCyc36taeB0yB67pgDdCqUjZeZq2ZApKBgko9Q9V
VpX74yEJ87wm0Z3E1ecpfh0DmsnsGLViWg/EMsCowuOqTYIwr5TobbZvUjfelZsb
4T/pFY22QxlO6pz1xHilmuoOaU3/gQ8JZWM6rI2SbbntwnBvUvxjQwrz1TEeNMGu
2PGgGpxIWi19CtRUejgQ2Ry9Xrj2eOeWoj+k3VKSE/O6NhQPplUGFrXEIUl4dHeP
mSWqQzV2s5tNbSUmmZXhXt47pJkpFF0hVatZOWIoIR56xx9sbPQbbg4t6IabzrST
mq5C85Rxzgj+sSlpHPo1RSKaRsriocL9AtoOun7YHnfdsKSVAjPBy0q8Rhnm7w1l
/Oru3XJ38IUTRd+xriRxPmYsUaHq9Lt9UZ0aj1jKo/yAl5WFGLGqI397t2phbYw9
BcxIouTIaFVIUuviYPq7igEswYZit7XTyDCXBGgC0cKnsQqIKxy03IszgbwcEiQK
/+PJ3bWRLgAy3fsN2dKMFc+dx+7L0iTo/oIwAxCP1K/8SRl0vT5W8Phlty1nZiOg
wgPNsrbeU7MCC/MfFiEP1KB6cGlSI3/DwxrM+F1J2GkbzYRNJjmXEYNuoOil4hZ6
15KAhWWxFnJ14D2L+YdE24v3HXpe/ziWX1C+i1/T0snYQfqVwp9422kpsaNzt9qq
BRgADwSqxAc0vsE3o+TbHiv5wUiRjMHWGUu1nO1N2DWZ20OQ0ZvFvX62kJ4M5qzv
a3wBCRJT2+i+fxIWRQpA+jwxlQhKcNqnB0M5gl6be97V5hjLS0dsejP+TpjycXoR
2g/D4jHNemHly589AFGnAjdjJSaVcoWAWkCvmUxDj3g5crgCxUuNn/tEPAwQGUIl
UikLPn822oYwU8NJXr8TpQvNZpPH0+1Ng0y5rdXcgxuC34wIOhxDPA4tXJVnq87k
6NTX1NEwlcTN64xJDzEe0uUCokG+7iQ/Dn2nyKo71w6RLitQMCVaf3pwoqV46zpl
maWqOS85OD055Bn7rETYdrvdsKg7ZMQAJy3n4wapIeWGz4r7i19uOvDuo1L3m4FL
mvw7KJiif8S+jQ07yFOMe+VVVpZ0c1iZz9pxIFTNiDeBtl5bB3LCYpgNQCsOURKa
lfXId+3W0bl+Qc9c8wvJpljyClL4d8KmKOnlLI32+UCCebnoLb4SIuxtT0CcgmPx
2BAMMfpxdkn9/5+s8TSbmlqhNJpPNJCbgzxQCANFNG8vpFk7Krd9lHAKzImaFHVh
YTgknzIkNguaWuRceU7/BLPbV+t+eaanJMf17pO/AIrhgHThFn5pJcr73hmNDnAv
x4qsLQeVWON72pf3T9SjPXPTPSzb9wI/mIecwRWR2KkBuSbAbzu5gmofOUL1tL4l
I6Ee9zl6foh6pM6/MNRuBOAld1L4Ss/Mp69CvZdUW99KBTu5ReXva+gSRnQ0/JHF
PAPeo8ji+pgGRIwRsF3eNp4nNNGERfNYY9GdoLlvzxFBTuylqMf0OitWgQUBZsdI
nmPJ/BgWW9+XLW1P2wqSXOVkHa+R0rumjplJCeLfUik4iSZLMnBeWdr4N+C0y15v
Ykk3yggwtUQYv37HY2fJ8NdEpm5mKbZS71Aeei1TfZAD4Mu9q05lpBc7NG8WUHZ+
/CC4OmZdfcaIMYDNxshZr8e5TbiRLjhC+EKkXL2zGIwc/qw3d/1jxs1FDO6w5YSu
L4UtT3S7Tu8U4LOl6jp7/du0+MX7TJLZCz1LQo8+x8OzQi3upuIF+OuRVVRLjG+O
ti7Bq9OTuTZmkJWPkQ9nVaYAtQe27Z76a3c2hM64U3vuSsSx6tUh5cnFCe0JgAYd
Z5zFJktPJePovpPoPD5f9gZggwaICuc77nk8g2HVRbECxU6D0q4Lg9BIXodqyIhx
ofwZGHlB/x1wrPleDWzklpFM0zK6XHTMjNOvqmhacbtcKG+xNiWuHgTvzRtvGVrj
wlEgk8OKeFQY42qRVVlBt3LyU3Xre1BOm1BW0U9oSO/SFlgw3VLA7uqKRJLCNYf9
BBv4wIktlmbflW8fCp386pcYDMhIPOute7s+gq9/yqLHgEfmvKJiynQpVP0phXn/
CL0sxdkSMl19uYJJb+M9jN3mu8KyRxu5sOJ/nhDvkHSqUJPuw+YU+UJAi4zisoRb
cLKQK0nxtMgF6dX7UcQkqEfkh9HSIAp7PBX+a4T9Frk1qHJ8NH1AFBPDlvzobOVb
f1KoYU15oBlULikwLeav2Nwj4xnsaJ9fbd+DYrb+yfETY2JDKod1HkvPb2lcqoPL
ZqQYZxsUHGODOlcjVrkKhEleTFLYAx0PNInV4VB9PjVD03U3lX3koiv7BNiryenj
dr9QTtj3kMWySvKa6/tFXyIEub9afkLdoHxA3JvWM4Hz5PTPe+KyrGx4lEe328KX
+gMtQcJeEq93YTITz+o8i4i1wH1A701PKkNgiLpyOzpLyOe+ZOi64nj5gR13vTqJ
4r4LAmul6NEMWkJOi4ppB7L9RFObQ3+UQ1cp0GCBhK6Aw64DHT4IngII6XB6GXbL
GKIUneM38nj5SVwMXl+36GI6HsD4817Yiz0VmeyHSFL5Hu2sSeonWzBVjS/N+3Oj
lujDX/WHuVxjKHpw09evxlBWG/GfjlVFf9npuYea/87MPW6DfigxBK0693YUTfcZ
Gdb2Re6NiXpYIRZRJI19vUSahyGav+ht+BCAAlkGiFodiPY2+8xVGDqxh25Kt+r9
9K0npawUBd0DwvE0kLXYKCQLTH2oFggPtSyEJMRX+O9Pj2BgNcrW2tmbKd+CI9wZ
WAPhTjOUXo/8dLTMFAnTLEJVJkTXLf46B6nPADg+g5mfcpFysV+UJ9eVEnxsBMWf
R7aX+k5u4AYmdj2+1+d8fYKVbs8XMkXECWwroWtCsES9JBqoZ8c/yNiWj9SHtI6u
aHkUUg0v4f1eIaRxkXy0azR7skeFaXIbMMjI8yNHhy4yyaQwB0SQhzMPSOC03o6C
YQMSqfSldbpeeyGICaNyc4GsWBzd1nYWcSkKZjipO+lTmHDWfdkWkOVfWUPB3j6w
iLgpFOqo9BKAkN7LGfqQ6biqYHVrjzVDZhS3/Yx5xV2diyFhKPoiraLzAG+N7nf6
HF7+KurA3TBDcDHk4B2c1NFNySNwc/f/3aihPgwjwXxiBY7b1yx48FIA2BKJFk/K
IS0ALXI8bYUqEMyjGmke9cuhJKILB6m1ut64miwBuYK9YxirnoI19v5hHWJzi2UK
pAUjTbQNHDmc3Cfi0T7C4qSkr5Fiz160lqxpw+I+81NzLVuiBWIzGQ26Sf01G+hI
Ybr3LkxiY3gHBCEfk3ehUzRFQo5GzIIhMEfaOvH1Kyt9dl/NGOHR0OvroVqHFgU5
FVMUkUeWRyb1GKMvcNzVLJ2pPg2AP941KyJxLv1JfHZaPY4hSAyZ0fW/qP6RXXpW
sLfbcSXAyrvRHmH7fSxymb2S2/VpgtSvMfv7VqhlvVe3Cs7Z2U4lqvYmPkFJqajL
tKwDS5oOFqQWF+w8FqjxKWgTGN/hyzYDDcWZ0//8WDN5AY1fhUAS9a7a3/WRwq5j
WsWIzLXF9MW8ORZ4vudvJ18QYqAMRIQzXIxyF84NQBqhdlHstHzHQNRWHYZo5s7/
Irwr7pHPUQ7Pa9SCiTYx30wFjFM3Cfqljo7qF94OgpRMAMlKlUOjn43VwwkZyfIG
r4jMX0XYe5fg/8j33NoQz2HpKmO9dVNhRX4IptDlJB6DBwWiy77EjGsXIzNO6sMF
ZSHM2ndO4HYGn6lm+4GW1H4Yq4Wd9T4zYpGg6gQhAOwfzhQunZPlL4gEMK7pbC8o
TL8CP8Vc41cXCZ87ouyoe5xtmivNw94pPNab4+dCxOSHV0W8NCvIPOo7HXJhgrr3
u7+RkGHMu4mgJWyKMyLngcs2jR8dPJ3RSy+8NIs9OFUmJDrAaPJ5Pc1z56TR4uqJ
4nReCM0y4rksDyjnM5qE2I3CZ74pcImaSWwYP4ZyJ56xiko8wc6NLen8csscXER2
oU546udXBUBtbqZ9XeFWq6AyZ9RkEnOtmThfsrRTDszirZiK6H2WpcwnllLTfvuw
ye9PtVsr2DJVSnH/FKgjBRyrvq2Q3hy+8oYuxGiElSsxNdFroCsLsXJ0zEajTcvb
Cx+N3lj/5toMRPe7EO8cs2Z8jUVP8NZHUuGvzOLMOQMPsijVNTFzGvgyFRzvqPsd
vx8mUxFtvvoM+nnHtN7/18ULDOujJsiAhi0jXgj/We9XP/bPLOyptyjO1Ez3YoUF
P6nHlCYvbWYx8HRvTE8v6vEn467OFaIFHOXqDsb/C+BDnHU+5XfoMA+6O/Nfx9Yz
k2ScGqOCtMDm8qMBItGVrOrqedc7ylUa2UpzteZF1LuUfcFXIQ8mQYbhl0Pe3nY+
13JrPdnhaUa3RJ3qmtSY9tqsjjOIinfqyrdlAP2BlEu9wRxOsy6LeK18IqHP0OEw
KS06MMtd8Ing4RR5jhdyyk/lqa2UNfzSxcOQuGXMxK+7DuZtByZxs74cSFeq1CNQ
f/ozZEDAX09dLt3+Ayi7YKjv2o/c3m75xoOr3ZA6HVLAMbNF9jzxGjamG5jPkNRv
/w3c2g4H/mYFZWGs476KoxnKGaipQB24QB3Sqoqm9wugpMc1bTM5s7Wd544yxp8r
xUZHurKFHvHYZbzX/dnqwxegAlL+IaXQj4G9XJXMUohfmrk2Qm8VrHg2qpc2l8g+
8nDW5WVWWG+gh+3JMDtOkgjN7wDUm99rarRH5zuiLpll8YTZq001Vy2EBZjmDuum
UKn7XSHI8qSB+b+Jtdx5BBJAYhcVqECWhkVKLW0UQNPIRzVU0zNvPT4JTtlk9eW0
fQPc9n0Tw8+Hm1QnTEpEMepMHkiYRG9b2kYG8ybIC/ngSFfQCgL4vcdBRNMhD1j4
hF9Y/FQNDjlgLroCno+KgcG+EC4LPxB63KnH6FVjlXiaXwQdgnIGSlNsI4j5bCuu
JPOSTkMT2zl+tl9+104A5UEDsYdaiXg0jdKfjTBdgXKlO5tOhGR4ufpAklR6TvRZ
1FwE8AGOJHKjfBGCI8f4PW+vWiHrqrOLhD+UJmrlGKWmy+E8A0dz0zJ5+Dv79hci
tjcumExLEHPTCqzZP1u6QKkBA9tZ16P+D6773zmFER8A2z7u5lqlkvUdF0o+jPZx
z7x+2QhhqiK3rT1QvRzjvl9eYfKzEd9Pe9zKSymAXTP+3RaZ37Dg8N1lJoJ69OWr
yE4y1QhAXKi+np7VFJ3RwTkjtH938QsTIwBNK+rzWM13vtpkso7ng73XiHDUptDw
TqIlNzlWhVmgs74p+g+KhDLRU3qkoQ5GK4F9WIgeGvNmrdIZMP+i4P9Q05U6w13b
iZVG9kE9el12Iupq/HRoE85yLU/vFKAVzwkyn8C5sEEwh7GiqGZfZITn6MqDslKh
P2jH127+QAkpBABynOlNQqcVqpr3J/RObd/ASWeldwvw8+iMJdIOryONDwUYL0Ez
0bgm4fwR+8JD+fMJSIkylTfi8Ox58HX5KUnd9PN9RmLWZMSQ23Q7ZPEqX4qu7/zF
yAKlfct0VUXRXYBLHJdA9BxLiLstsUrnBNSqfZa4J5X+cSXHF/QG+HkWxZHt0ZtP
OGn6HOXZMxjBMXbPiiYyDE+aZi6cRJS6i46/PjNCBQYOiYhnuOzRb22QmZb0NlaL
PrRmSbDi8fMlVVYfBlFXjudn9mBW9U1hOLJw0V+AqZB+M6wklpon3SV1TgAyiUAP
Qz8m9znDcypHNaRjLoj2mjr4Sm/CehO86Y10pRkcB/IlEH2EvTEb4nRMkeYCZ/Qx
GDiERLQV71G8NdDQ5z7jt4em8719Pw5W50Qgrgeq3W/CsvknDY+nf5YgR3XxGQwq
fGgPmii3tfeZ2rCxnL6QwFSy89H+cayXu1f38jI1LCgyfcXsesD8I404/QEvzz6C
gwMqg0jb8QhErtaYNkKd+pB3SfYX/ovZawQggG83Whg+k+FAZlTqbsu373jz2KF+
nTnsF3733tXa50M7tHWD49e1rH4vayF6QRgkCMsf9jvjc4QOsZ582nSMK3Pe5M+B
rKGDkONnM2WowLyTNG6kFQDZpo2+UH+wMDEeDEikGCP1GKE+y7FCrIsPt/9gZred
diQA1I8tQW53WMFBcTeoxugdDF7HQuodjTwGaelkPsXtifw+xYdhYaPRujqZXAWd
GyQ3jhiPsllQviUbORjuwWd6oSKHYkC3kPrGtGfiLIipAjsJsDPEVy6kJN7UhFDj
eT5g0A7fUlrkc/i+m+21B9wOu2RUl+TB//0m+yicMCOIMnGXAdqSSdvALhVaYZV/
jkQAq3VS0BaW4qm5OsyFRB4Y6dsmTxT4x4r6n/lraIZx7VySk5crIHIzzcb0LYx3
EAuIGwgDtEhdkPGbvj6Gb5kxAfWjbgYewZng29LVNOkKKtBQ3L4x1uwbe4xV1VFN
wStU5mEV5pu0B3g+43D99jhqAdZfA4jLT88DcNxrl6vJLm6DRU1bdb2zg1qtRDZv
Nw7BnIVGD7M5NMIdpbRdB6nc/txsk0VeHZIUCB6gv3v5qqg0A/aNsr77XYt3Xmi+
RmgfN6Bkp/5SHBVaYKBZYBoW9/ua+N0nqJntRqmHo4e+e3kiGZTJmDlCGtH1j2OH
TWfM9f3MIU9kFQ8RwMgG8vMxkA5No3vFxrMHBs+5W5haUTBciaYEY4M0KI6KY3Yn
V5XVgbUcSjfZ5zpXsBuZYjIPF69OCDehUM7OSvYSLLLxrQ9tUQUWpW/l2lDrW4xH
qsXqzJA+NPOV5D8v7ojzMNRyCChLk3l5ETr4IVl6MxmuOd0Q0Vxck5i/amcLRsCJ
48J0YLr9DGwveHI0ykgvW24yE20mStTiVGs02da0fzFfkiYPkB4GGK7Oy2hwpkSN
C5fSNP8KQ4RuGqn52H56eOiEfA0Vgt0ONEc2YnnHWGWLxWYCWaIpuXU/PE7m0MTU
OrCUpIb+GYWEsrYse/6pRtLum6JuEzJ1wItYefnHjbg+iC3ecZAW2nTqQSVxW7Wl
z9ij76i3C8PI9Jbnln+k4gDWBW9K2BzLbXLXiCtDsiuMGURq+FRd9d0j3Lg8mzGw
UeVQiBh9/gmfh5is9YNRMtljbDe9T0M02YA6kCRra6viNSDFNgBh6CYIxtA6xUG/
S4GQsC4UvL7JRSBaxF6DKFuBrvUhx6LbmwdAscGM2CgqtIkpChXop8JPGivQ/FqO
v6IZhRCumd6rS3aBoHwuLi2XHhAgbu9kRcgWhDTPiPoEzvtxvr3vuWpWkUiT6bZo
ql4RN17Rd3wpUYN0yL6F2w+yiWsGXvW8Gw83vJzfUd9R/TK63HiHkgBVa9tpxz2e
4scUIQlwrH9HyD4vcWR+l6hyapq0dLcsiM2sSPawgi3PpBXqMG3EVmTb52MzyVo0
0u7QChFOv7ZUJxV5IPVo6HfvyeL8jghuz4mS2Nq8JQyjmCNiEh+LXCMPFdMdcpck
Ncv6x2/N8hJV2VJtCqDtCWe7ZDPasArV5Y/LqiRLaizIln8P0sf7xIJAfLUDBun3
1Aa6RO0riaXpg5YWGMUna6NnOxiYBMeh4f3DfSTIgAZ4dpm7rzncd51UPDc16Nty
MV83Zsqg8/GRXAeRvGOtClhQH/UT6Dj0o0fZL3pgVtFyDuV36suiUzSiLg3J4OSk
9lvS+7/lBQYQicjPAvIFgnxKbg5cT6LJW+ReYm64+TwStnB+nGTLR7kp1KoczFhs
4Q7OhIPxHYeE79ABP6SX88qAMKhlRY32Y5JUZCi47WLtF5tiAHRPwd7nsLqV2vU6
WSnC0WNQW9INvyKzdNAaBBwLKrpHwYVn7FVfPp5lsmWyBriF4opOz4GM2hrE5pIo
vM8JfWmQSP2x9dSeY1zW0LvGr+ho2S9ECOQYVHC0aTK9BXNtl9dRjfWVfTbjyBc5
M3aQrbC5HeoqS/yUMYQv1bHhkC5647ZV91/VfIveE4V8EKrpfS4MlStzbFC/1Lhr
Y0iW7MriaUT2ResP4L6gX1oME8Y7ish2E2r9uLj3Cr1YH9InPZYVNoszK4obd8R+
W4RIRIZY6O8gS2dyB6t4Ipt4q5zlkXaR2TZeW9pHYdPMOiRUgp8T5/LtrQlubB6P
7IweRUiRLSswWnB2CkY+qeTT+CdYkqmCVoc1s/bXVbwuONcMwzaCUHQl7YVozzHL
62Y1Un8Umrk5IGhW23MAGIqWfBU+j7T2CLxI23mg1NBDoQMQXDKoxauBq9P/eFFp
3+ZrqSPelz9H+5vByYP07y0WVhlysH3OX4OoIkK1LuG3tEdzir8hEu4DCOhO+q7x
me4pHxbwYrZzQg3bazcZYRtzA1ElCvAr2YXf7kqtJY27GYRi9mDhj5bL4pd84rxg
8xgnbqYq0EoUmePGLex8meJH0J/tKUlCcVGpXHQIyEpQclpzdZHebkTiFTEEEHDH
JOfFGlodl3skEkbxfr+FHWIae/RTVnNLBi8pnQmPNjyuvvKE/gXakPbXzLMz4T3C
gV1NGmhvOpRP7M6FxzE3NHSjM7gNSL1I4NmnJlHr4cIi+UM/KdEJ88wRUREsPF+9
JrIfPvdo7R2oH5W++FD5SjamyJgK7Sm+pyfELLUnIjvUM8PO9oY3OC9XiMyC/HCJ
XHcm8/wUm9cXvwaHrG3MGglUJmlXlERnn4tTD+GgE4Bacy+wlZ0jtOdH+OikgV00
vJVi4dfD1KtD+rT+FvbBkhf/pz3QodVlMAfGhuuoNqvKLv2hKgZHd9MAmRWzco2c
5YyF0dexGDkN2Rf/ki6mRL+MRN1UldVMHWP/3i/NDZqVLKCPTkytgfW6bN3y5wmk
NJjhHIfnbU67sd7CPNj59q3xeLTSXwgJoTeTau6z/CaP7XMM42z031C2BcWOAxy1
gkVe9n1AmsE9wXjGS/NmZtliS+8DTU10OBagdJJdDP+5JB+r9RuiiKSFZFfhonHb
xNjjBeCI7xwSTq8eKqqoWjZLPVtGjwdwzyDfTIaD0sQishFAnCQGU/lf/dmwwIFk
+3H3o4FZJFXS1bLSf7b2uvkIxCES5p2IaQIXeyPKYprWAVKkv6pa/XpTKYmdS0Xl
0yNxJSRtoaQzGVI5d++apJ5IaAobUOKG2lBxiZU9RW0zABw7GK7SGRCy+b7EV6Nz
dpHsz4wJmP/gv3s5PQNBnkQ8UnSkZvgxyZmQ7TT78RS/laAyZsb/K4mYxUuxgY6X
AeO6T3dnZhOJj5t5RfWFFgb8qXkAjkXLLxeQkMTYYzDhZeiSnl3h7id/U8ptrZn8
dHf1VU9IbQP/U5EVkJXtTrZQ8JorriEJo9jn4oSEM90z5BbinTgQOEqoNjeR8xWj
o7XL39FfbkK0PgNDAGKI3dUREX/ebvwP8foBkF1OAwgMx9TEKLmtA4qcznKP56oR
NWx4IkXdW0y3EeLFJHtc8gQ1YufgbAvO8QE9dWaBDz8ZybQOSFLiIDdBCClGfccE
zB8i5Q2JntoIFYJ8p9+iBYiLDN7YTOIaQn4UfYDkRWYo4TAxr8ol1qebcxmeOW6B
uXnafsdKvu6fnxhKq3F9RtlKl5lnYVsW2ogvGASXbKTYAgpwzDhDkKSB7Qp8Cc2o
aoyD9kSjBv2p3RM3lvabJcmHDK9hPSRDPsEfJwDO7+rdcFkUdiClap+pP4FguHkI
Nl1qGCt6QlZDbFDfWc/BjFy3cx3nq6wFG0Yh2c6+W0BU9NH+AZ/qDBZbEP3oQvyE
oQjj9yyORtLQrbh3oqc4Tr8b5cHfnHbcYYecirtys4p+BqFeDZdVRePjuYvm9wfX
Q/nSBWihd2qpPe9sEn8NJh5mv3dlxsLnseSDl1Rb57s7h4R6RAAdMe39CKb0QEtx
z94k+KtgOGCPvBxki/oz3QjcH5pBevghWTcRp4xAIZLXho250QES4C5vPbmhHsZW
D62HhEIDKlmVbxV1ixamq6/r8dOIKg8kLDL6Bpz+YjEDtmUWeNQa0FTEzO8eEqGJ
2aUwx0dPKJuRo9zrXxX+fOfoIGv+UO/t5AE5xstmmBQ4YdO8Ty5Khn84QrFGu+1+
/0AAPCbYk78scjWz+20v53C4y0y1yeh4Z2rThZ1pL174kuDrG/9rrXeZiDuSQ/gx
wPSM0zt1ZgZAXiyRsXGkUFFgjcWSLuW6LvRpBr2kM3npF9CBmg71V6nUS3Uz+1dN
Vp0+gnhHnvVl72RYIHRlRRh1iFV6DTtWTlKUL2qEm9ZMvb+O9os1roPH2Sa6LH0K
3EU/NdwV4amGmdp+f9zokGs6L5zvKYX13Ium7Iv1xuE4qvu/t4Q/PwoHCyktqqAP
vILRQ1ZxD5uBrmR4mBxsq0ixoD1twviPGZDr9gh0ygg39teZERyGTP4dnRNW8dDF
oEIV9Dn9RhdYt51kwINA1MkPmGE8BsvZHM5dcHTk6WffE4WbJYhLDBLJvsNx9iZh
q02smLh0WM6jTDfvpiivC5gp78dCxV+HWxrN5g2f6ZHylcoK2lXs86inibhIFwZd
ifJ9Ggk2aw3k1fBV3S2JC11yXqipmmrMq30/U4189iYJGHo0IFT0hiL4tjItJBoI
DOSTqPOOVk/TAlOQyH+yy4f1NZ4p8fb70t62Q8XdtgOhqY8tO8u42oqBsHGJUW/8
C31vITjMc69He8SCYaeFeymvCCdEzkG1mFyuqnmTFRIDSRMK59AGY7lnwkzkB1CU
uZ2LsXjsRGsw8QSx1P38gfi2JSFJx4i41wskycvApnBK7SH5iEMQHDEbLchzu/aj
TjEmHXX+Jbf5koWZ1G1+5izot8r/t0iQJOC4N74HQY56lUQ6/Dmzylw+LoiX78vN
950SeZC3T3ba+qRRefa8WDLGs7v698o86UXEWarDxbruS77A4Wfzpz1sK1XZ2t0B
LtFK4hIFFuiQoXu6JVJTmJrs4xZOv35wHRJ778Fjsd8L0Mu2wZhKxQuQ7TEoAyJx
8ZvDWXKx3BYDKFZa4/YSkhMWoD5YcwhL5R7pik927SclPWAPNlbKYU2PRhEUt2Ft
h6FLWI0wSXbRMUB27zsNd/9Q2kzoOI+G3oLBuUC6xsV59JTc/T6y9k9wpfRzR4FM
JpCH2xPey8PmK2VFoj1wROlBN/hQ+miTSN1F/BAo8PXtBQejK7wSV4IA5YP+FXlz
ocpU7CsbS/1+YmwbanvomtJCmklBU/QC8QV8J59QFqWTLewWH8vQf4gpPycLMxU3
P6OaBgL9W6ZF9DtMsCJjAxYT8/Hju+5uYBZRFyDMDADJkhKeEz5Xpz5v1RGTUCPt
ok4mn/gIHtXP9cgvcuEz1q5TAMwTlywqnRUfGO0RxRcBBfkEjdIeH+ewzEQNxlDR
YGdiK6QLpWib/3i3FKn81fPaJrBWwP5YX7JA3+1ov9tKi9e8x43Ki0XV10xl1V+K
gNd83Y8D2jIEPtnzy+gGq+swj1IYcWuQRsDWDkCiQPk2C7lCzS631Y3Ef0hEWaq1
SXxoiNPJ9oKZmirX4BkhszWrUPmPiMuFqdaxxXRRBL2cT48UksPj1EJiL1mxgb54
iuP/mPc+9/KXkUaXPrVbHwlo3T+rfOZd4TGc3w6vHv2Akr9ELzaxD2kXAX98O7Cs
foeGS91vyuwAtCyDtHIK7uxmre+HlpQ/liLY7gcGA9J63EbiMwIaCBPk4l57B/Du
SHc8FRbl+vVP41Sp5Yoy4he5uBox6+IOdYKq9GLewZm7+PF2I0CIWfoUqIo/SxR8
WoG6qJA+BpnfsACLXq0RzkhOw+eOZ5MfBDvyoeteuUVRw9DrO1xgzufzlVNPYBNE
KKhxVZUImCSoo0Zbll/lNK18P7DOw6dU7z6hf0e8OjseMDh6G9LNi5qERRuKdlAx
isgOf1izZlUnE0UUyCkbcxlLmrqocqr6QSKaKQU0Y9cV0zHtMecS1wwpdsw0Rw2S
q9zjzCnf0qYRjwg8532m75b/2mG9+YjHdpirZicc7pwED2mZ3CzOoVTyOVssjS0D
4ld1FSA4b8XAwc/jClU4AVcKWvHsKQQyC/1WshTTF/elYYY0tM3SNNfqewMRZ3F+
lkXnBBTc4D3rZni3Jz232gMZPvaeybaD38a5YnSBi9JBKD2tKITeRITItNRewCGG
IsaEnMAVPx2iZZ4OINDDz5TW7er6W8bJDxGpCwC5TiWJCUM/wRC3Rq5fQkZhZett
g8pVhzlRwupLaUJiBWrQIK6/TrWPc7xaBZJeNLNESxo+Xjx4I3+lKG+Z4+6NrWLB
mPMI8q5exoChDVSlICeJKaFPGbU9Ke4tBK+cPBeCVjdV/uniNJRfYgxARoAOEsRr
1q27pYqgNn7rsdXLVc9/aA/WmhX/gBy7JML21Fzgx6OerXnMRKLOMK4K73EjgMd2
cgFeBnIzPMF+ntaJnz5/8khKUsqMzDLKEcv1yyg9vQbmauZbxzrjQOSTO9ux7raT
cn05gDsiQ8BfGS81wiTiNwepiNdYLmrA6OM6CAxSc8PbrpmZLjgLX/tMmMkLBT89
/c1tDe+/XzR/njud8lLhlvd7NN1i09hjCcKQALmOr8LR1bgEGK0PMVxKnlfgae7e
BZL22I2Es/0C21xw/kW4LR5tLIGF3GLZEjLEJJZ8yshVYhcn1RiJh+BQnShHrmhe
Xcz2egTatbjMaRIUR5UMlUKA5Zzqoy27P7cNNlozi7+hYCuNoFErpEd6shBbpOFy
YOtVF04Zn7zQfCvQzDgJ1ZSfQZy/7HgWJr3CuGbdsNRtMhueVDu1AybSEQMHBDpb
4kqJX83/nScgHiKffTZTa+CW6anzFtZq4OnICu702RhRtGzrFVGAU2dfRadPqT7p
XxFwwrQ5dtr/cPcRORw4BkbkxTiLjO+eQTkqL38qdNh+y5glLi16RaUDDnxF9zlN
ArJoCex9s21cd0iqL4yZ1ba5kshWDhqUYQI0sv3fixzBnAvrVo//OzrdKxfkYkWK
i7hX3Zcm3Pk6PLhsIiIE1zD6rAV8kdfch7IEq6xlEnkiqcg3iRjlnZb6GI601V01
aXbKDMCmNof5ycdL60Ij06AfYoE4XSSUXn+JNIyGG6LNFLj11YYE6Ki2N9W3T57J
wpnHWr8I0NfxsVMckRJm5SX08j0gbtwzZV6+e6yJEQGfp53Vk8jIsh0LmJ3JZrjm
FhpSzawIQlCBQ/6nwZxmImT5Myz/2BhI3qz40wT//abaR8tJjdEZBi0vT5BgAeAy
RMb8edbG63rcihAPgSgRe4K5avWhhcO+9AQDS9ubfq369BSP/rZmV++UXetOOYLA
6At8C4XekeH8ox6yPB2dEqtkQ+u/bj/ojn+ukLQFAh8hLF0NXhx/3mEEhtXCK+NR
73OPYUOPwW7mFgPQqmJjnRF0WEZzMz+elbTgegRk02TH2yHZVf7Wcaiyt4MAEscB
0wZkMzGWriuqs2QKkBiuWnKtCoh1SpsRfxBL/4pBhiDSCbvtPbf/kDrS82IsykPb
pKROEaoTT3OMbcLqGcPvymM+l23tC6PZc/4QfswYXI/wd42InoTIPteMFzRGJ8SL
Igdgiqoi8SLW9E/0ZdgWztlNEog9SzI/u+eO4cjcdFRS/4wNip7xJ0MCvfUpnuqr
Rv5cuXGzJCnq/uFWA0TG15hdxJQ+4HgfUNhXSDFr0KwGvI1TXuz9zhPAl9BjWg0a
7WHrz1zEXzGzeX+ZWDdqlcG306yIfrgreYGKqa2VLJgpwAhzxu30TUrfr10EWHsG
tWbrjsrXD8D7PatfEBaqT1jZJbybrxRgDWyh1Mfa1UuC3Dq4SEY/XdNCMvBpVxkJ
z6HQn1sgYt1/cCNdaTx23+S6j+L2Q+wXlHN7C6Oqaycc9mSDYnLfGf2VIHQTaOJm
0enBsCwwIVqhol7uHxadca1ztkPw0OztwYGeBzs+6NZz/jLyfok7QIJ70qTCW2Rt
W6BcPzjj8/0+0EI1wxzYLd2nXkhO+BpK4EVuJtPX0hSegkkyANbzGm4mfmACKCJP
rTBrSeQY4cXBu+th+fSJjpZhkVUVn8jQ9U+aI2antDoRfe4c0gFHjEvk+SYw5DZM
jgfxlCeVexT6/l8PRcVH+Rt/18vNHfke2Bd4NKufo+/gAIHnWudqK4uHU3Hz199s
Jsk1Ssj45bkKLd9amE+mmCYVT4bP+KTlGh8UkffvyxStxjOJV+ZGomHh6cBaTliP
+05uXw93F7OJaAoVla2J2UMAC97faS6qjYyF4ZszZRfnf+BF7cE9X1p06u0SNp6t
Ui72Vgtb7zqUcFRnfeyGUpMQMR5ZZIvHsJGiGI6MXomY7Wlod+UJy3IlKJ/iVWXg
i4vY4CVElhhKqvSnu3mXGFcjGjx2tKOIMQosUteMXmzNIAUjBaELKYQtYN3bZjsb
J4k4K1rO5aWp2+yjYdCzuMZx546dilQdyNmNrGfeYfpD9/fu9Wov6K5CInUXvJu/
fRisXmd7f7ztmwRwvAIYHmsJZn8wiSEFkydTfnxQeeIhB9q9T5e5NEm2FQx5Q/tw
G0jACbSR8oB37b+/0iC4OWXhK32rdNQfT0dg8CdfToQYaRMTVD8SVDrv9NyG/Xql
QDbhD8zt9keI/Iys5g3ouW6qmEROb4osl4/CFAyKl+C1YV5rnk4YKQSGkRy1fAbh
7U1TzgqwFHIVar4FaleEoU6+4HVdy8pfQv46UNzn79SKzrWi5NBMwc4x7i8/2vhY
eoz5HqxJ3zD5/z7jIJiniFMgPK/d7PG+mhfUMJvn70QwHJzMlRDfWYRAJ4fcRbgJ
yWsDq1wFj6DnIIMyyUmvDwainFCCewSG6ViycsfEKa/lDofs4gkYdSqFV4tta5Rg
0NuupjXNQzmuWeO7gMwZASKMxNMR0AoGuhSzMueZTpSTzdtXsK7O4RB8YaElfAxP
i9B5m3dEGg+wQH2qPxJUwF5S826XcloNBILZm+EZ5EhIuWYbMOPwYOTdZI3I6mzd
z2vID9AZmEAc+w2A2C/wI5VTXrh5tg0ZiApDp26NsCWgjsQINfvi76Z7pMSmWUc2
2Ai5A30X1rDUsJMssGl1Q8PuR/mf2jLYMyJpnHhjDJh7/RJ8s8KptKoyFAv7oJn1
Pk8Mph1w/Xe6rbeIKlwcMY0q15wj4TC7Yo+wYX2r40lvQFlqjbqvk23WjzpOHkYA
23Mx4VZ8b2c0rR+Ldc4NfuvIGropjeo/IhpAlF1sB/lfXMUPenvWBfRpIzI0XaXD
3CvoDz1lA1hcCJG1WidROJT9ogiiT2a+xQ603z+QO77qu1vi9GyKmyNZCJukG1So
dj4AJCDUkxtCk4ZHq6bURsq8g3csHeXhjCzFx7Qtcc4tFKnv2RpJG/843lsr6Jss
oQ55U43fqQQ96nF/T0qsgdYN5fqV+3zNa2EB4IrrXBjJW5pU9hjt9iTqsMatGe2B
96ymSGq1bdMMTfSOHyf6Bx4LTvz4dVWcp+10u+0TH2zc7oi7bTY/6gFGKXa9j9MW
GgZKMKWCvY/9fVnQ/tkqWrmPckZE/Sykp5B3qw73fU2g+wGvMaSa9cBzq9mgqz3m
OTFh7bGTyZ2nGBmiNXWdPryhT+qDnQzgh64sg78EHFISM93jpq4R1G3XuccjQ0yG
Yojn3VwfB9EpVooZYois+k2DKilUMOw6m0JkHBo6uNviBhCNuS1VZa4SMGt+XCZx
Fa8RBQStgNqUrmjTK1i8jWQ/ewcx1E4HNVsvdku2bTOSdv/U0i09osFe8QyxFkzC
TO5WzAk38ZvJgtqVEJUi4LpzbBgHy5MsJgsTOsG8or00tF9J1JaG5Zs7itwjVa6H
uSiL5LWn/ABcD8GCvVNazTBDXzkDT95TbsRtHNj5gPACEvnzklWLzvsH0Gyh5Tlx
c0kyweoegi/rpJY7Tfi5VzpM9N2icSZMvDkL55i6rX8Epd6Qe3ItSS4OjA9dswEM
5nk2z9iSd5JVixRfmAnhgZc1T7xtmSR5Er9kSq71ODDyv1+FNcYHAZutPcITNp0j
9Wul7g8e9UzAElf31F6aEKaW+BSCJgD/cwX3Up6SGzgMCBRTx5m2whU/fE5fb4VG
nWYLhsgPynx/I5WgGrA1eclP3Jc/HLiq1YDsuwXW2oM1iXLTmz0yr+Yh/AB8sA2U
UmseKnSPCv7wUOvTa24myucGpSBZ9TeKvIBB6Aus6RHI3NJvcOGMOWcQblFnBNHe
v7pcyALkuxfwkLCG7L0LdreM/kW0sxYAKG72q3PnU8Ezcqj6b4r5gua6rNq4jCa9
qJiA0ryzfQd2lgDASJbxxlLpeVrOyj6gWQYN77sYrWoWM/TuGWPiJgfl+/oAps+T
sDqAHq+10RgY0EzBhw6wCK8C+S436Z4aDy+K+BsiyuNGmQxStbFdQGkQ1g2FlHvH
JkcBJ6F/RygnFh1Si5vdDc9/1pOmNkXjV5EG+cKMC/dJE/wvkCug9vScIbwHNJTz
OLroRxroSw6ky7wqdSR2nSDqkRbxwA2ZppR3b8vdihOS4QydPjVk1Y2z4AupnXyF
7bi35uYQshsrkp8Hd9OC4wN0rlKxVzUDvPpt0zLK0iwi1FYSnP9UxSiV1ynsXxtM
uUXskRQk4K3+jFWZnjQPaJ/R8RYNaUsved8+Q1HPqjj9oD/CPBHDWBDFH0VFJG2t
JBZHJUrQ59sj3x2EIW3TDIbrg2lwERpIM6kE0tDloUzAVL04xSDKFyYvTpWRonbB
ULfoNBihzWg9P5MxhfvLe8ArxOSSkGHMTc4ity5SqkYPDvZsplN9rN6DPtWwbDxS
1529gK3kHoSyixQ3DCirHM/N1PzlGzU9os5BnfG2oSc1ikE6bT020vajTczykMwk
eypwBGeqFYUXW/PUaZWFaVM6Gs/jVJqI7GIWjn5me4Vsi4aZV3F48YQE49NlSTye
wkGObhnR9Q5kgneFT18vIuh4GFVFKx+R3gQWtiMwqWzfFabFd/lAEv6eDYW9FI9R
+PToJmEBE6wMDNFqXDPhHVtRCUUCBcQ2gvnrUjmi8mAS5B1H6jBjjlJWymE+PfjF
QPlvpzjDJpq4qEw0pDN8Y8u3U+nfYJZkcEPTBhroKWJkMwUAY3yHVvAk/V3wLZQZ
4vA9kSG5Mbq+swh7RGhIFnpBkcJWUKgl80ElLapmQkDUhGfNsJS6QzBS6DEwvKy6
59PQtGkrhtfdFp+4PMff/FHWM1akknKvf5/B6K76x09ibVDx6sFPELtnEOIoz8ys
muD/l/75ngbfKLdYrXehxiVSWKG2/5NiAPcBBiekm77Hwo8yD6Yj3qCstj4cAt0C
mEXJCiWJxmBHpS1qWgdqW9i/VV3XkCTMZ6SiJO4hHNdRfuVPZnBdiUXH/Ve+OZQ1
BfUXMM2QkiIzPBHh7US5WEi/CRStkOBx/WWbAzq5TyhfuEXTH1Yd8huv51kzYJCg
Rp/YWsTGungxM1YswN1FpXz2A+xjTeGWlntd08leA8XEKVtfDR2lE8SflMtGy40J
ugpAoKngrnMTh5Pk/E/1+ZMmMYTUdfDD0tQ1OdXodNdxXiA7bEl2vzRH0JeYWVS5
2++0YeZOGqeurkETY5mA6g0Qb6+yLfC5JUXekmc7iOlzrDwFyBCOSSSDIbw2QVAV
dKz4QZsUyCq3AP7YauLdTZo76WbuCZ+A+OZPtvJkG+Yo4V3+k85maI1OSQXEj06N
1BnQpOSzASxuNWeukPfWqXzi0fc33DRZ8yhttHneE/7gi/ptPsu2xADyCrVaI0fE
YQKlFrw6n9fs/aCyR8xZwfIyFGXDOf5BXbaSSXPH5HcozGgRRjFCPmkU1z2P5dPW
YpsPCsi5Svr+lrIsZWD0Jktx/qcZk8oRiH3CzJzmfp25NJLYZLPRM/CjM9v/V9Tv
w+vDhN6ViGugpi6S8ZaHuAx4G62Z5oQfqqsud5uuld/H+BWu0FXGd6IX25KvVXKn
Dz9NWwxtHujqakniudeL6xAbpu0e02Gu7tzsWjrbWH0wdQ9NdMk44ewu08diAcP9
pnVj3mbRxoThNu7YqPbaWQmoRsMO55m5y95mnQCJ4BoSeTj3hjZZWlqptOVFj5uK
A3SMeCsrNYBd0yDNsN8yS/xT0rwmmYduehfqxiRtANXxuxZPkDn1r5IyAxV+Tfmo
dYkBomwS6RSlc5SyMT6IitWjVwkmIJL2BEIdxhS+fYD5FThb9Lr4A/n7n+uEjZH+
uwvE9I8OpEhSxXs0n9ua1gwT+q7+a+vj3yjgb1xzNvSyF9DxhRS8t3/UGAC//zrM
XyE8wD8PEoi2pNzAQqNT1KNnEF9QI2OTWYgoS0A3abo2ZPCWvyHD4+rHfxBTS7xn
CfS5Lc9Up58MT1pkESx8DMeje5NbKhmq3sQ2ffJkgexINcLeHAmqMahwNyRENlO7
yaVXULP+pp6IdQVVlqq1h9Byj/Ak8OqKWr9cCm5dERhKB6zpg509xmMq5EKSuURM
Wv7BoTEwlYE6K4pNj/NbzWCHCAhfnzyIPfLYtTPbhs8ezlYQtEJ5+14F1YsTuvYO
YnapBhWHrlo/GnCWF8wgy3Aa5GSQZ5Gdn/BOuVraOaM27mK7brLNvmOrzUgGUHeC
PM0OOOSnyorubnN83NC/SM1ypU4mD47hiS6rIitbURQUbGoLtHM4+hNSN0K4kf/f
2kyGX+RxMu+MwEgesqbc3oopMZC2CYSBN0u4ghMgMxeYqCRv7tItS9+KlpEGEHBS
bQN5gD6Gb+CFot2TWOnaOEvkZusPduKJatrnyb+6ik/rWPR5ptS+4oDz7geTou0v
flTjaKkJCOYbpxFfCVqsiG2qJMXsm7ai3VRSRRgX7DJViYGm/4k0LsGMOdzvPkjQ
QNfao443ZvGIz3GiT+N51cDX0dUy3YaSkOPWmko2Fx6qyCYtWfAJdyVu/4VsoK4Z
CWKF9ujk7av9N6ZWQE1qZ1u4o50M48gaH8ti4D+9ItG6+nPvXWFnYcsWOy1imWoI
cKapKU+W18kDpI11MsK2diLhQGKzs+EvG8duipo6d2iEjKAFKVHvwXbFGSSjn9K7
zHbkeVYSeCQWkpGEvA4scfE4+BAW56jhoahKwla+uzWcFyAbUZnhyu5XFmX7WP4p
PgBuQ9GIDOICg8K2kk2F7sF0epBMoXB94HI5tUEQ9xac/gM+kn2zoXONCE5fPITQ
AGjjsfkiP0A6Iu1IOtnj5VY8vlnMvtAHVFWcfVXk3xnyzFfWSgeu3HDcgisfjfOC
jmJL1SWEBIYgG8KHrb6N6OvVjAyOJVYbLomQYyjbrLClyjQpm1s6a95RFsdkN3mH
TItluV3pRq1teDPHncZivELER1/Wy2Yq3hGVUG8xg+y9UQTOoeVMGOHW+279YW+n
CiFokpTXXQ+A+bq2ZfIuw1t4ciKX0B2g0mZM8tviAUc0jZvkrzss+USrQlsqi8pi
i+xR2vp+XnQrkw+ijUQzO1wHE9b3JHHrEL9F255/U9Jn+9FTJO6nccGnVoCxQH1E
Zh9RPK2L56bbnjKtjQ6/phRyTYfonRvYMn7pyO1+cNixm9hX9fC+j4QuP+mpoT1Q
/jmsHGLaZMKxBjIYY76e8+tb/7/y1uN0bkXKdw/M+81L/WvaQnc2+LaYnerOsn/S
Mi878E/PafMuP/j2UdtHkvO9qUuiJ5x2Yt5O7aEBJCr+wGJZwf7gccC02CdeDdXj
oziR7dR80Fz04iUKHHag0uyUDxn/3r3/IKYnQeMaN3kflhTsO1e6Km4x2CfdJ5GE
A/3jA38BswUiF06FeB39NHx5BDwkVo7DSkpG9/vHlq3KwXx3iCAXEn9H1r479LMY
oaB9RCSclrOPKVB5jxt3GLt8x2SgNaVLGtx4BU7/L2z1gsYzqyiPfGFJWQLxtHK+
6iV31TYI0MUyyeGOPev1yNQvNsvkZtrlhZkJ3IQR0MEoLfUWEpNldyxDeDYfW802
8ffAMKjvhj5jM6nP/nZZhjEuuyd/nSLwlt9MePolv0JXXNJK9YSH3bsC9MWJK5hQ
2gbaUNhRxZc2NW7iyBvn+uw+P6foZM+ERmk/K/NkM1C+NP+AYdO1cnMSKgpYY9Mj
FE4HxsAa1ojni2Me85otPegkb0MuU6xQYUqbm5vGhOzakjC8moxvyKlWFrTkHND6
YXJPNDrZ2buQ70A514vJE1UnR5FwfmUs09LdRiN+VJhtx9q5ySbySqn7T+ArTPlI
g1N4miR7+3kXABp74P3dAOgg4g/y3oo7xoeOdZ0ReNDUKKWkYeC9ioMUgLtRHzE6
IAzFM6ePvqgnhsDASmrn90QIo7bcj6AZaQnOANpBId1NuDFfeOEbxlmwDrTKS47t
/Js38NZtUkCnGlZBztJav65pMZIvXBqOLHbHhq5SC8leGqt8T/Ninr/W+o4WJRHv
QvUCXahFb52HJS1iQgvdknPChhIXipUUzg69KhLouQ+mz+JBck9Q0rxznqAPJRmN
h2VKlBqAFhoAygMsw0Hayb866zGybXAMLJaenhyLzpxaOg4GpHeYvAIj/vz9fP5A
x76PWhVidgN8+/kyTt7W5TSUrdX+SclBEMC5ABtRw46ZVFpQcFee8glqG5G248DN
3GzIfjNApUJ5cL8VoYacmHxnQ8i3r0fCZ3F1l5J9t1djnxA7YMjAOxJIaa8PO3Bd
6q5KsbWwoF5/64OJO16va/jzgjlmFnzojiVnpFlXo4mLFIJeKZUXWcrkvl31Sm57
XAHMofKMHDgoNCvcND4xMYiVBvhEO9J9g4t9QlYUjo0AIjkCGeDGGizPc3pB8Kxy
Y1HA4qIocVFpGpWiZCuytmJalwiTzwTQwpgGWTRtyC7aNrEIMZlLLDXJLbqK7qaZ
48L8+/3VgiJpv2JxV367pLEvIGr0/wZCZdeUlx1y/7TvBh2CpYgLPNVLq1fLSqhg
m2xWt9RHdd4uyTil2WbJAoiBe9YfJ2Zu0Ea5ufV6O5d3GaJjYLFo7Gnhlt7p/X5c
9cAu0Jwdycx1+A9EWomC8v0Xpsd/uV65aVcYXspRuL6Uo4fbwNHWPEU1Y1jYhljc
WWh0GmKGHZwXW86TXBIQ+UiTRXC3upOKtT/RVRnogP0f5L/S53AlGCoUqgfNRGSX
977skd3H8Fn4mxPjLjWWgTcV0nfGUyAq/qZDQ2uwi/fRBNnTI35QVzY+qF+BTyTK
pv2nFdaK0NhOjjufmy/N3ncsYkKeiYBqHx2E3IPMltpaC+g8zM8z2caJe0Xlg1cA
ikJpUlE6FXsWNYrc1so71+8hlXHiQHWovI2HMhUiiVULvvAuTHwm8iExJB1yeHrM
mEfRhj90T2YG8cp4jDIMs0PbIrTuwdL1EwCOhcSmAkd0zgFqDC/Qtxif8Hzx7DBt
4cPlmX8rLcDRado54rWHP+m0+BmewEvedfo1sXh0L07VMvPD5z3azUiz9zCasTey
T0kWAyxocLvp9TP+zT+NzPSWZiiuku6FhyhIU8RPn2S5MDgbsHQ7/kvqz0BdZkYD
a47RpUHsGHkNcOfx/YqIeI4HaeISgnNO/dJJwUpKhqYup/VM2GeJCEZqYMBGZ5AF
INUuyOx9QQL4wbsPR6oyLj3blEy6W20I8NSv+UzhSPfMRvMIJe/4TaBNxuPGqzE6
JSr9xipQ9cXxeB6/v4kIEgUalywLtWfAL/cwGwGmwd8qpyjVdzcr4286k4dqsQs6
BWdOMrEj9a/B2NPpHM+Qp1aLJQqq6WHhi9My8TPMwwPGu8NA7wac+3QT7FhTAFWa
h86U5XbhWiGD+yUG/aiLpYopBLhyWWyAiVWSbTQ2qXrLVoE4vq+otBxvbtJkIYCk
Z9pPmTA+etetKn6D1O1frPWpznatYjZzVYWfWDtG+7X6uSfPHt+G0Ulvo1/7Vig3
uwtTVqghM/67EBayg+ecM8E2oApLj6uSemSMGWxsMSaML826UMDXAML7Q3hlnMNH
oEuxJ/Xts2tlwecDPZLzo1zyXkErH3PLS+rAZfpRSSaAEACogehj2nVKFAI457KQ
zt9BTNmAjhCeBnXIMFyIB6+9rJ2aB+wfBcGH+cmu2f7wSWjUOQcz2YdZpXVZ09/f
bkl/Ur7Ufsvr1HD77tK/sVIeAB1TWn+nzt0EzXzNNmnyfvSzzMvaJZCMWJC+TVA9
vjlCbrYW3G3fIXyNRqq0mPd39BxbYU1w4gCFOQdPhUCpCfyZl3nxzZf6UPscn/n+
m3tsYAJVTNJOv3gGhyTSNTiootFUleYQxVfZYkdNql1P7c+xIl4X42AFqc9V6EeK
SKeGzp7IZ9WBOzF2Ci38J+GXzzl4S2z2E0dxHnHTXNuWNMKeihIC4LNK52+7sBwu
3KuAJqVJHmK70SwnQZyD5uXcfjjcyGVPviI8Agiuk3NQltNwtCNr00eXconzwH8Y
+tKqHq0U4nHdOOOcHLllLejTI3XH8FgEUXQKh/TIAjKyHzh+oNymW29bek3bD1cv
0Lven6m3xmfhvyDqRGXjNSSpwn9MBuvHMmXeGZkB1jNJf7c1O5079gvWAuUW1a5q
+U9hQopyj7QeVmIIpaG5LYkTOCAei6EIocPGz7zn3j+g1oJ93FdISQNi89SuHlIC
CSV/Q9stN6Yyk+5J2w6/NpjkpIE+7J36IhmwgLCLyZpPjaKyCKgUUqf2mFsN9sYW
hOwOuKl7f1oh5jXyStwzGrVVuwh2q3RU0GIn2LcmMmEfKPrAW/dPJSfZO0cCO4+p
4h/kZAMj/6nvoKeun2+Awfs5bzukfJ5w4Lril91lGQok8cjxPNk3djTqgk62do+f
7+cG3eEY6hGQzcKYl/VbGfLz/3fML3KpOQKg37NNzBqtimBoWGzmsXwW0j2fGGk1
eUyDvwrWgFVNrKuOErI5byo+CcwWL67objyhsbQeYLlu/8AsM/kR14iPCDtB5eOw
7WQjPALXvEJVunae3Pfaw1HPjbJlhHSp1TG5dO2HfTTlL639emCzpcAThzrKqewu
P8zVXWy7veSTNEGBL4M/98tjUT+1dpcBevOXDAURoFdZy0PhmHGU8Ksw8RtDLTNy
G3bFqvoF+7RJ2Uc2dL5JtcUU2gOdcCmyTmPEsobK4zWyaLLPwhQZGzWeX8UiqQvS
vdcp5XHPVip1UbHLjtPxqjvD8lBE09w/GTHf0IhsjjtVwVNYD0xWcYZMkohAJiGM
pBMI/lK8oNGEqaNrCdvOwMh1tXS9Xne5QkqqodjzI2RzebZOd3gOj99t9Ws5x9dZ
i4dgcTDzSQxEX5YzqWw58aknsXvc+0kJgB3vB5iv2wOsKnMd+7WaGLkuNvlgNJ6G
EDqicSUfB3q0u5NWDZSv2pnyifruL6kzmmR3BmWJp8P2Q9xM8wNjVgHSaz+P6S3D
TcLwLTbF5Au15jpmcggtWc1rYsslHwow6OmofjOyKG48W5LaStRNKHcJIe9oZ7DT
lHw3QMnNk8ngVj08MNbvk1PaTQZTtBRe4kJkmK0hj1rYSApo1weCy9JEZBxTbJ37
4YCEpq/mtQ5e/mK3tZqJIHNhAmt9mCdcL+hI188+A4/ErfgrSDHRqqKBnOaTfqnR
kZEnbiiRoVxMretmchUBlPQvhaONCW1CgSHgN7P9luXVAuDzAkTPvEY+sLTzrBnW
0Yxt3fX6PP/sGJTsAK9HfmtVPyjMqnWPKxOLh32aKlk08fkRTO1Nw463hq032OER
zUHnMYG0ejuys3FbFXpBdd1/wIcH+/k0hkxW0Pi7g0G0BtmjgE7/nbotmjiMqqfg
Jsj4MEGNyyUqNZNQUytKwHKcSJNRmGi83/xcmZQ5DlG1YG6gi37OEJ0/Ibe0JJ9M
xqXl2F97ol2b96Exkio6Ww5nEqohlhDWYh7w+mxS+YQAn67gtbwm3mKVQZrfNmgC
oaEcSY9ijjevxjZGNG03pO/5ry/OCRpcOtzGGyS5nTuN0I19fJ7oNgbRoUbncCmx
XEDrXieifviIo6F2KYMHYQsqauj9DQWpmgRQmv/yDnH+0YfZFPtFwmGnP959wy3v
8nDzfs2SOnuASQ17D0q+KmfggJwDpZxxXD/MSOK5dmxykZPsf8enopNX8afuqzi1
5fg7Dp3xqiZJjaGtx6vjOwe2DcMTAr9OyDTBeSq9Eitm8KiXnt+ZrhuEsZktUOT3
cnPCnKArw1rsIRc6gLQW3UlTOzGoOGWfMQPaVxElxVRnoUQG7NOe9lWwhJzeETtu
F4HCav4GaHoWlBJ9e92nbhRe9VtX0H1XFlO7imb6fcSFll9nftcf9dC5XiFY9Fvd
AQlLamf63m86doWx8P5FdAP2IIqS8xem+xYng8XE8Mqu2VB9sDL4PdiutbBUQ21T
cRbUPK6xkMR2Nk/MqzzScbtf4hX+8CPCR3Iljv7vVSGxijRZnY0wiKVcF4uKAsnU
jEbJRBF57dmev3qko17iwBtOmAPk+ae9ra89rk5QTUbOHezLGjGfbtmWkJQ0yQGH
lvQphXzgIHhjgKycEoFLBiCQXsSwbiu9syZwGUBuWRvLIXkAK98j1LH9rdexj1xb
Kpj3aRzFYUt/NI9Qed6bhZMzO+PBVyveXJj342GJtjbQMWUoNtdWuMWXOuwlNsEQ
3K6Ppd6+MMyENbb3rOpwNze5LoSTcE5xtpLeRrN4/MZua2R7xMCW5CdY9iOIpMF3
HSDzg3PgisQyF5wvD1Jbo6E/23J/O76I+FZyAyE83zsy2NuVN7rBA2pp44+0vmro
GgeUEkwViR5QmCVuBK4JNylNg+07KFmf1Ti9d+fRyUKBxM74ggczWgwYmx4rL8Ph
9g20vVCvL7Z4d2rdvU3X0YJx9RvYggMGNecHpyoSAx6Ao0T7xRkj5yANn6OgRUc4
kvLweBvNfuv1UcmMi8Zl3E1T8lDF3R/tyLNeiMvhCZma6yqEagp9bv4s49nyVi5Y
W7gvIxoNeclPesrfuEHzmqYcnwiC2/QTkzAAh59c547iREcs4tPyP0AcVGXGeC97
4M7MLlDA/cOmIavUwJBsa0CQ0iRF3vNnc9u1iMxqGaKYxI9AhPj0dE5HC6norVQC
mYVMUcJEy8yWt+Ghe2bWi7aaHz3gB2G0TjtPXBR7zytIzqYi5J3W1V3vChnYWFxd
bZoTAN8SAZNyTxKE7iZBW+cZTS63WaekiWeMBsB2GBTmoO5/67zScsx+a7Ng3pG5
eIfLNwIyI/1tDGUUgke6K/+JnaGpAl06MUd4QVLjRX8WqlbW30LaWODp8r82qduE
pwTg3FiS0VRaTuav7fOH0+KQjGVvdo//ZyTWwCf5RpfdjY8eD46m0VuBVOWi+z5y
26N0UTB5Zu60PxS8MAzqfBdXaHjrfG9Qj/YMvmmRCw6AVN6oSoSFuXyVqlkEi+D/
Pw2LinV9qePvXZSPVzfQoLRVQ2YLyn/t4ILAypbRqFmOi8LP2mk/d05caF8a4Nzb
ERoHst5gGzpe6wrov/wPvnTPnZdnhRNakTCJbyiKoLa+WQhSXbJgQBwvqn32DgYH
yjIo0PRgyWwJGHmOuKjns3JbP3lvcbAAkzIXxdlW6K8NUm2k8BQHgGNJYXLUGPvp
jfQExRrSE4S98m0F+e0l8gX011gLAaQH1AIUiImEVv52j+AgpWxID6AjNchBKFRg
AYoHPAn57GQ/6bW4pAFC/M7T3MMA3TFExMQz7UkWG2QJpMaCQw5GRljWYWPTZS5L
R9iMs+u2CYtuCTasA918k+MlqlSteFHEfNJdlIssaCNZ8nRt1gj99Dx5aeFVC92Y
csX58kaqx46FZ065fUz4ikwCmNyI6aSlRCQa/FBm0Ejhyq9AKoec/zxqdPqQldBj
RnqhkO/cB3sZDHCRlAEuV2jVKkkrgeGytYBK0ZyNjHTAO4wVcnEAbvUvh+y6aUMH
EPKmlMB6dM1NzE7UugS2N+6zFk4CV9mOeRWBCJkMLJdG9q7bfvETbNaeP/2BKCji
uTIDSGsPahpDieBCLNh4/xLtluNAZpv/b2VuCZUjM3o0cQIse4QkAglxB9cvQlqf
T98uGV2olKHwusE8AITNSawLzjmVo+J1popTic0kYPNwxZJCgszLPipqDmHHzC3I
zh2sRralEGfQ43ZiO5HB4DTXDum/IQLBScH5XjMCBrKalymAQD7lPwehxVG/x9ql
UOLBuZ7ZKA+hatePnUD3P6P4drRPeJTp8WOf/yd2xdxqipH5Ho+A4umgoEPsLZKb
BMS4pdbnMqN4i8pE6Zm8QDsuemFtewkN85enO1ZmMoi6GwC6IGxUi/Odkubpe9bq
nBTm5/nue/ImJ3TF5UQT88c5q8aW0cXrLEMD8ggutCMGDyBhoKV3yx103V5qGqh7
05hpL+GVTX+x8StuM3dBrcGNrtpiF6Z0s70QfA0Hkc5FaRJfdQp+NQHuKmY3dCd5
W9nALPtxxeqZG6xEJJwmlVsFJB97nOBEK+nwAuc9KwcSwFJ2SOVBif/BDKf5t0ay
5KokP2zpd8BkBLlWWcnrdT+lpOpLDsDDbMTneoA9n99WMNpAzxuUTrV1uoFq+ss2
BmviZKGbcN/Rblbjr/Hx61rvOHCL/jpZxmqxTzLFkBDKJXKsZC37ixPQbnAIDpmH
np+LMqZTDqtlb8lwLGFGi/aUE0fDm2ByQKKteq68zqRXSUV66UjTnmjTTci9UJUB
YYj9McmIlv/ASlFEeD5qq4rAur55nqZJAehyf1WFdYwNIClowwcBCJaO8NGnbT1h
SKS6HuI7lMa01+GWR9EbNzMt9gEiNAheCdrYHqjORVzGrpqANzVugkDdjOHPM5jZ
pvh7/U8v00hRIGn/a38kGuNDSvSeBw35tuc78fXyVHo=
`pragma protect end_protected
