// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:55 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
gCEaH8fCSDQA9Cc8s4p8qq8YSzOxf2JP/GaT9OoyKTa2s275hjl33GNrZPWxbM5z
AmcHMv95mXcE6R+gaLVdqcdM0uvJcR052jMYKZXoRHhmyk5fR8cfurb0BNmsrVB8
iuk6aylXcafE+VIjiU+lIqWOZhjZ5DmOVpla7Kf6ZMY=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 4768)
om8fx8ds7MYEApKhZcNnpl1q4SvkUuRlk8O+kGDb7rB3saCKIet5M9o6QmAY93D0
HoSPxOuB/Hyzkn9vltw0/NvVA4EuXQlUBsWC5fLYvPuLfq3qBXmDt9rwduywGkBZ
sNtKRlBWJYDkuguwGhHVPjW7/HI3i7hjAsu6Pdvk9stSeODJoGM4d47oyY8WdNEK
720GVb7rnckatcbe4WloF9MAHkXMCZp4ATPxBxOyVMpGXymolxmV/TjO0DQTgsLd
vON9hZG7YCa1tWTK49KOcRIdv5y+FQDUN8/MbJFYvMdqEJfjMOvPnT32TpLB352v
kSCWwCLPPYBXb2i66e++Xfil9Axx+8HCbPKa+Hwec72vlZu1fp/adCVeKDTgBPyS
fKEANU6zb0z4QR4fLKpsvV1m7RvdfEoxuuWaUEs3H0ShMiyDuY67DxaNFH4+l5jx
xEF7GVWEsP9lAAQL9aMbs5b9h6w13Xwi04jhLUl/JILKcu2wYEMl68B6i+9oKcbG
zQhAg8tYp5Ucy6oumrt4udnjesDpy44Q3zingJe2yEIR7gP5n4J1M7aTUlOib2IW
vcosEHoUhxKU3jpI/YWrL78AhNtOXfwRVlcObSLFByrI+gEw4fwfuV9QeVpTnNuD
7et2/hPEvo7SWew0qmzFjj2F4OZX/CCbj5SxtuA67fWa7OTqUBRR0tQ1QyRW2uUQ
I648aDTN8F/oddiGzYCbeFbBUHMv5snR76iBo7AVAPm8BjVpLOB/OlQLLyGxI9xv
DSCurPNO+5Q/lrG4T8TCtxpaxCYI2vUXI2qPrO52bqHN9bqzqJhs7+Qp08B5Gkii
P/MhCbVqpVY9tbd7a3rDXomaYvCdsireAkiod3Ggt+JrP/hfxdVKEl0JuvDClfnv
faUzzwrv8pSZOuuTm8hFnvc8UTscqi7jR3Cla8Bvk2qBMYwDXg16CCY69cTlIbxT
xsFCvThlNhU1xArAokBGEZfbc4kUPB43IPt7z6N/EjIWDS8F65anPF1DOoGXgejx
dcRKQxrmsWfVaizzRTzfk5hL1Vg2XMk4wdN2lVrmVNMGDZxEZIUfljXknHiyPCrw
GktLp2hqqaU9EGrRX5PWz3ar+g89CncKXYVcTOo3rBO9hLo+bixiiMAHEMzILadT
yoDpZnq78JSVDEetm0k7iC0OBN7wUOd0ivAl1pgK/eA9isRvUpemShyUwurBNj8X
yWdxPCGOuHHFzRu/apiLmJbMTwym2c/FRfngKu3eB735Cc0PbS8EFVTbkLzi/0np
8Cp8OahSPTWo+ueb3RdAGZrYIUbt0hZlJ7uVQ2UszWHZtKh6iqxDaUwubZ1zFxLP
ZaJwrOS/E25XcJdJnzEeauYvLA6ZGVTrP9UJttGNYLkBUFkdFj+xhYdGKYJtY47H
PuLCQKhslp7JX9eQLzsNsXv/hG/uLI/zbqjoBV4yDqigY/f92pY0wXa2YVKW0/JD
Ct3z6ULXu3a2vtEADMcAgTg1Krmr4jINzOfUcSrZ3Hc5S6SC8SQ4QAGI3ZJjBowS
Yzf10MVyd0/BecNFcmhC8y5h3N1bhyDnBLJZBKh41ulCpTFUz7EDtlDmBVleIRLp
iWSQuVOPmT53ncDi+07Bsz40jj/MLj0+2fkA7YNvIvv65EhC0ne7Zv8zwXNtfLi6
8zFIKJCHkogTVJvrszAtYKBvnAc+lM1pRo08aKUT9lj9e2VMiu5wgdHBTpdou7Jo
HG9xNTI+T3l3BtE+ptPDthiHiSGaB/VlmiBoKV0CHoXWaRLwB7oTTu+cD5/XBbxN
5IgdjeKL/EALBR3BHOb/Rmbw0DGTHuM7PmMuO2wAInA5vDzpLtqHjQWu6gy4kTWd
U8w7JSS5RRfdJiNteNEAqhQpbMcGHHf72eOTIT9eRlFs7NawiypzAHmYk6ufNGJJ
jHVeE5ZbIKlNHM40E6VD7u+YqlxYMECnYrMs+jjIjR6S+odtcNVAoqV8751BobnD
N0tEccSFGOPXs++q43xw4J8zEwRAu4ZDAHu4kYTFnt6hGRasPx84qE9K/QO0t1ka
/5xMAU6MNcAqyji+i+to3u7cp310eb4Y/EtmiUmlsugScmxHOptIzTOvFLsctrCf
eP4V107cprym4x8bpLg67rSkY7POapN0TRXXfc2ZY1bzVhsUpoVvnJSYjynYAr/2
nd18Cm6nviNwCkwLsyZ6NaqbCEFHNUdewPgAYocWc9nmXhHfXrRfI060pgki0P4c
zbnEl9q1gHvL86XL+D/SJaJ3viBdfMd27UHUBTjUurdAa7yiM2xONZ++8zsM2WbM
0dpITkhVLP0pCzZJT4sZr/Fae4UexvRaJrK3jcUiyMfZSzZNW+esqAstBsBeA7b3
99Z3ur/1KRmgCEvAHedmau6Qlcf3IUpAIxelIhzd1YrcwQOFupqe8WD7m0eDBVn9
t671S4YnRDcXmhSNWcNeGk2om7GNh8u3V4kt/q6tBaYvWdRePvZfOUGHic3XwNFL
rdyU/0M4ixy0khOUjzw9QVNc0ofdsLn66FIsWe2lhBqjtcXSXcO8QrPjSm+A8HDo
9tcokCd5XrrN+SFb2m3j/4oTd+MW6AbK6X4itYyJ0HpUheVNeTNRZ7EaybuuxWkX
5YXDc7l8r45LeoUjTx+hI+WytHeXBAUytqMGcV7sRS372WjtXvpcY4E2U71yNAOm
ryCDmUX9WIMAKIXliZiGQMFMi+dOvGu1mDi9LMduvoh7+wIfdjeO0kpHQHlfzIuU
9SqGYRNn2OKvprZeYqLtetuWI5gccEaO+gJAZY8bFOE0u/lo8vudMY8BTYznz7jK
WaO/lQ8ZPHGAvBPYJWxhDkDmhTxjCRygnsAkJlFY/Li68L2fBXbDnjT4zeQ32Pr7
MmwNW31bcABmD2G3cDL+74pVyQPA8bL7NiZ+AX4MPZYfxzc/nSAKAPeMnQB+w0xl
hnLt7+klMXhvpJa18ZmRiM5tZzMYVnrdC5oJ0kjk6tBxGvKJerCfz1c3D7znZTn4
2FQmp3XU22S2jy4FECGzIaIHGAMP276fI8UPuJtOaZjIqzv1LwcVZxN/J6pkWz03
lOxZrKXP4Cg89/Xz+NQ0ZT/o5htQAxdM84QgppLuYeQarxdwELOmhvWnO757Qy75
3ynW48NkoMFAEd6UnIxr7CE5EDW2TlTKfQRafCXRthQvneAT7U1sObvBKMa8s6Oc
lRZ6Xh5Ft9sE0Z6UEdLBqq5fttxyXeQ+jyfL16OR+mwbjEQTGLiyH+rRfnvmUOMh
zURx7hnYOu4xgqNCeiie1S5JMLD4e6NKqPJuN5egnYZcjgo6I5x4LEWCBAlh94tH
zRYwrrr4JQ4w7O/F8LCC//HAD+AKULj1eOAQ23L6unQPNlEiX3Wswi2zUzcFLSfi
FdkSn79oCeTn7KSj9PxFVgEkMe6g5aVxWz5C+lBKkkoPMEbcH9SfqVNF+pRjJjsB
gM9YxpzaCwTDYQ3iqMWMiCLLRFvo8HGN3R2WCEo9JGh9nH5vHSa9Go2qofeBbG+9
R7H+Js4Bwv+rDLfrfmCdk4lL6/sXAIQpDMlQSM/NgjAV5NT+AoSiBCezQiq1ffxo
8fGRHgfJnul8Kh5AYzGMEIva2zq3LdE51HipqwgF4yydWCOlR+lMp0vgLtvpHv9w
niq8wvaz60FnQ+doAWcwfcuzviIH98JctsKwX/sZSbjnvuFWBep6BPFldvreKtzQ
4BhvryBtfB0C67dnmgr505znK4qd8f5uutUQj1PHJ9Ol9wHRv39gRpkxoJdga87v
aFfG/LNITW7R7IjRqAVgdYYYsXJvkX2CXky42Ikls5SZo0uFRQ4HlofliprWxvgl
c5Jh2OqJygEeGhChlNYQbICmKSikoYF3FdC/0ZbTIOvygcT7xR9jbbtHJMF9eZ8p
2O/wL5KY/6TCHMfuXg0pDwX/5Nw+heAyYshZ2djcYpFN3gMpvKEU/sMlf4aSKxdN
/AjVkP8tqeKZkwdhAyPuLW+YJY6nr5hwUXchvptZa3y/d9obWOhXUzsaLHZJT2NM
xQ0btMXJWbknha895FX4/CNowS3kmGlaWS6ntGrhoj/mB2mIe/VivaScwOUehH4M
kSgONqJw4Qv2A9UXPRVo8H4zZ6F1eJ1HXM1VdmHphToBTVDI8AYp4gDnkXEMJwVK
eRVynW1l3utDuks+ggu7jnp84nCnOrGpx6X0QINFu1ilCNhebVPpuEyluYAPNWT5
Y7igJbODhLbV9/7Rg01tB4Bajoowerlky0vZS3VpSNkGdBoc9lJM1Gj5csow2vyv
VLlktgGMkF5XkaqhPwYOsiOkf8EMdlRtXP9eQY6+D1+5DzPNL/XhBznpVSlJPDNV
iLl3rUsNAnXZljuG5kY4Geo25Khuvnziuda8TY+gKMjBcDwhQvypFflTgichA0C7
eOPaYFxtqk5kMnt1o43ks6X+E+/9vRFDP3EEUoXFFsqqUnA9UBgakLIqokbJS0cO
o8pqrNmegu7VJxFWdyB9h5vmoFwQD9gDkgmF+Y6b71fMDEePYsSt+4yFWec5pWej
Fp2ZrPfZeQQX/fNp+bYNVVlGOZmsaTcxsQDkBR0NJ+l41qCKhYdYvOmBXYhc0DKS
gHGoDq6YDRclF6mzl+yXmbpkDwHsqKny4cq27Fl5mAu9M0J8avoYjrgXhwCYmO//
AZ3BIULReMzQoMVQs0ZqAKo5NVyBqqe2Jin5QQj5ncj0L0o2lgaUCdnxWEvJqHyk
1+a/0KJu+l/oydQIUX1M407Dz+KA6xp035BZvAr8IKUp+fLHePEliJUAV6AQ/as3
MqaHLTR4XuHp+cv9a6yJ1kC3ZnMau9optPGhhIa/Q8adHhQVEmZ91CweHi0y4RwU
zfPKgGGvazDRGKVXkEYbpyAchdxSTaNjs1BujFqbRNxsqZlY4WEusV4eT8qjCLHK
2Beal4yfSA7rZZM2Fa3xRSy26G0bqev0Apu3O5FfQEMnWnkDqfTRufsM7cm88JJ7
aJciipgzkydSszRohlN6nBbyivMU5ITqzzlPS9qu5tiwUM70F+uyYOaO/vaMZIv1
Dp1AtQ4xnRQREyDGpMDNNLiwf+rABIJS1EGiaWl8TVhUEmBj2AxW1FSilSaRfx7b
G4C8ZUl47Vb065V3JXsYFlNNeLLiCe0IVk8xu6lODLIJ1vbeiXvLksHo2uG6iBLe
vYa03Io/2eKHwBnz/H+M7hRJzVmkOOHBxUvCZlmy0GKeRIwIUKLuT70K/IluEiVy
f8FYeKZh70Z0lLkgAi6JVpzKfgMnIMxmSIlH5v9D1YfQb9MYzLpfZATKtuKTOosL
/I4hUJ5AFtTO9gehPukwW0WU/myDGw87X+aBqkAVEOHAGZIzXoeR1YxKGmDfGJ3T
GH5rnm0kVclrlcGTi/yIyqZQTRX2TWiJaDO7himPVU35G0Kngkd+eRi0kYByFKT4
qVlZlG0uE9CrXhoD9vmanhHUUzltNk7r3HUaDgMGEDhcezuoGxs6qYzXC7CK5Swy
pRtFPAv4rDRcJz5+BMwwhVh6oLG1w8QLverikYmt550B3x5t+bWxSHqTpWhSdmby
aatPhTsgc5dz/9zLt6v9vCztswoEhS4RjE/bMDCTATvXwniEIFFg9lfguOO68rHl
stcUwuQCH6xdqu0oVxxRdhbPZb4AQPj/m+cdm+/FoLxrGxTk7eLQGYn2ANwp4pZx
d2Wkr6D3IrEn22HxqWhQIKmAGZgNjvptK4xZgOnKsYUooVAeF8BmpOcCA5rnh7YD
jWl1DL0lYtbE87/Ch74KlKo1ejoMpQ8vf8ycDdQRgemTAkMkoiOi32i4WiZXk3x2
5j7Sdi36L2FLkl4R16HeJnlie7NB5QPdtTk3NAmRponEmMlNaW86slpcCeAhR/hN
TLkhLaT5/VlzpVogsS1RKGN5Ecq4Xyepc80ZLQpMtstVQabx2Mf19axC1JYhBQbo
OQcS587qiJca6MgKuCrfniQOy8rTbQZuZVr7V3nqzZffL2iiSHnmHEGY3p2GRDRz
5eNFOKgfDJIM709ukhRFPlOBxPcoKvGrDbYrAxNLdZxERTPc/WTGKSJUzIkO7WM7
qQ2xMe3sc4bhcdLG5LAslg9enGifeftgcluQ8Gf/aX2y4zSzQjwNlsnalUGa+OyJ
HAnEF181aIAhXvf/gNYNHAvMZV84o8eMYM8OtaTkCA42DlR/BXDFd7x8zXvX/bRC
ndEuRIMehbSARctLZBHmPIB+GJ5ph9i7E0mU+0WYaaxDAHq1HBnF9MGRzk1ZA7Vf
DkR9gmddv9P/ygthzjBWHr6gsmBM9n4+hNHyjZ0st/lPH3kG+vbHbMfj5E+wp/ng
SRhgdeBUmkWtpUSNFicCxQ==
`pragma protect end_protected
