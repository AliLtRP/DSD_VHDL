// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:35:32 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Ne3NItCs0QHVxNxn0ZmILUV3fKuasRrWNz9a3dAA9wIPIsLc9gsCOJqnzGYg/WO5
A0k5a+gJu2hqFqOodgeVva+fPDKXRPkDaKw5Z6eYoD7Nq/XIexztlVZJR84i439Q
pdOK4CmNx1+Nqn/loqo52BEMQOOOKLnnoS/0sP71WqM=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 6368)
7cWMPQSbzklkGmaTCoG/fWr2KQhGSklFg5UeMrkB+wOzfnp/LC7xawfGaEdFNOGt
Ip5SGN5n0dvy8tnS3L8MbUAtRE+A/H4cN2tjRzvIc713e0bwzlp31X7coYt6FXlz
Ydqi5gRrVpqNcnnMPRbkM4wdmLsufgTUsnMG7p9aYOG+QxxSktwtaGZseJD9ONzF
8SnE59iVIBkDTUlFhX30u0f/MAkzLw6OXt2Ba/jFCpomkUgd4LE1S1owxz7yVjp5
pwPpSskFykisTr5Taa893vF6mpTTymDX0QdyWcd34A0OBiXhKdbJ2LDsq4eLLmLi
jEBaIr+hcStPUtEOb+8bRG4Exmqb03K+LsIXSRQ+ZGDonqELmXRiyNxP6J5lKiFO
T6D2O6kXv3VrzBcyBlAsyRW7Lgd8Noc+JrTuHRy+nqlFoovjruA2UA2XWJ7gAKiG
YpBlNxBRetWOSHNo8XaHvm4JfJZ+HfaOyNDrIuMpOUofTrQltz/0Jhf7bigHb7h5
H/Ziw2+S/e8g1Jle9IUNkz6MELdjZY8U1OMaWCVYtwqZUQcbAd7/AIh47Vf9n/rP
vtodbPStWzAhyuyylWs2Hi82VKaBZZBXR+SGpsU7PXrp9ZCVtQSY9/4/pS8AEnmV
g/zUSglfYU1cra5f9WyjSiF9MURyebZqiBUiQcg1PoLY+YDM4VuSoVhwMvnYSnov
QrAvauNJzzMCWa2ND1MXRWXQ64LHkGvd3w6qkq93G8McljDOHmnbQihvE8Xb08iL
4kFIUC3nOZfawnQd++2iGobGUJ+B+S+jRh2BtNBl16MAW5ZGAWPLVSA6GyS0VUAs
m9OQmCoOurrxmtM0oguSQ/dsppN/l55Mgvz9j5zlcRvlq+zTExPWK5WINtUafhLu
pGvIkoS7ieT49owHLSrmN1TZgLuJsl52DO6eJwC5y7rDKaOIZpJyrPz1cnOMFlhn
U0ycStlZVvoKGEOJkSH/6FyFtN+YeoaXPpYsL1Aujm6fcgJP0jQl9pK5ZrQlSGkY
UzYBNDmNLapl+4JimBnNhMeKdMns10Kjs9giVWUpqTxPT0sEDd544Tc4/JOc6la6
g44cBC6pZYmONP5aIeMkHv6PMh4MLNE1fit9J80lMq2JvTlRLt9zoEszBdzNYPrG
Toqvtl4jVi3iBkJTEygdVKKzKs8XyfV+jMOgyEB8HPoZ7Ubg8lDXFvrRJXDec3kO
427+igcgf1md8AALuoBh4pgOzNSrK3Ig8xh1HQoHyZxHQM3E++nUaF7xBsXSnCfq
uF4NVzpSbg2SKFRNTNZRRWLEEUVUnlsMxqFViYpn188UUJ1M4OAymI81joRwN941
R80xxC5AlURHN4gj+4hug4yKzjwyI2BvKsUtQeZfnWnlAmi6uc1z7veDOhEqE7zp
Om8l+JqvXjGlIbEjJEJuQNplkYCVoiQKVjslChgIA4VEj+T68mJFDAuXuOfEtiuS
1gCzALFZZpkMWHVqwnGMvazx4/eBre7HVzxV+oSPzYtFL+wLBy13IrJf3IiCe4/i
DEGb7UWGf0yH2wGzNrG+Sgo+CiRXr5JgN6IcSxQgIH/dW1FBQxIEn4+7KvDZJwQT
ZdTc1fmH0StdIYu6O9Jo3Q4b8qC+TCqcCTfgIF41Ab9rQpo7YTl1oOVaRO4qu+c0
f3nmQ1b4FUqEoD9NF11X6EmEd+0Wa0YggP4zeo/NiMEeFfqoLOWCjfPzS9cTo4ZY
mJB9jhQ/GKWiWnEkez+y4ZbmM/JMdgPYaorcHF459UEnbJPgWbWdIo30CG79w/Ez
JI2UkDRda8elTco4kU7tfQp6q3jgyQh5n/gEHczfx+9i1Zz8HN+DU0RJOJSIFQma
Pfb6EqjE5WISjCCF5zFV1SkA+7HTuCe11ekqTw3xDHbzxRPa4VQuzpM99fxmQ1YV
a3FXaNf5zlRd8E9rfVnMw6SDfkFOHixF/mZj7md6GpKQKxInSWCy7mcOcz/3G5qk
KWA7gBB7yRDh2THPHGUu1qjNkWocAUkk+/9VxCRmFbFnQ+6CNUCMWZaKiAbyvU+t
P3Mj+elp5RCIkU1Rzkx1ccNws4jpV0RxOMqSHO4OG4iLTa+FNrTJC37jmHB5rfGZ
98XRwz3jL9I0IuJmp0L6IF4ClvAbfwzyD0wV9FQY86NWswT0miCwNjEZX4XuBTUO
9ZDRYrmCvrMrHnRCNN5jnKphLIOxPqt1ys4sN2nzZBaGCyXNcvaxSCcDtya9anGm
+PPlkHL/G5epAuVbg/cPeZuR9PxoJVwQuYaBOmXl/dwKjoeLNDx1rr3Av35e17i+
eXfOujhJSg/Cupzf1s8L7wu+MSypmu14NTgu+jbOW1L6e2YJOHe0vvCw3iu6Fp29
LHkUWnjJJxErT3fL0GpvTokq+HksjertYHd7PwbSvA51bx8KU4N4HTsmSym4i3wB
+Av5FIGf4NSJU43Y8fkXoI1tgdy4IdkpfjFYz6qlqj1nodApm/9yqUZGUBaqmFH4
55d31y3SQ30FQCjnsQ8oAoASWOerY9mMj6H9NHDpyN0L0DkUzFy4qsyHyl5NreFx
ajwUPkLDub2HTLedCW9+vpdCiZsCKq2108k1rjTjH/2Q4bRuwywTh20vVnkyfiig
4feGjd2wuDkmg5AUYUWNvgXounJJQJpb8MxjZnTVwrxXWONwiCaoEnN/DlnSxXSU
dNpq/jyCPJPZi80iuQUL5IrjSiVSFoAKQcPKjuQxj1wYrmF4M3svLjrS7jBhoQ69
xfrKV5y4A7Lb2E1dl8k47BOOqLnj2ogrlU4u46vpVd0o3Jy9dZAhdndDeO+wUody
LpaHiruAA09Kxi3496Qi7jI77KO1XZ36ARjTVHvr7EQj3o0XVVBe/R1iTs7JrW81
qv0+1ybdWw8S245M+4w8u4zDYjPn5ueptZvs9v5KqmBkiknAhjCAalM31/3Z2kjd
6CVwS2BKaimnyc9g5ogxXNfX1/QujDQnl5bg2jxU97BLS7ON4MOKE44dONgXtysH
6C4REqpMFrXmGWqiRm9Awx83lvUAP94Gz9MvG6zQXIJMHhMTq/1K3V9LC1kdGx4u
wBxMnjo0U5TpM6oVZdmco/dJeN2fVssnpb+890I7MenEqkJJBEKariq2EntIzxPt
X19zQGWJ/O0cQbpI9c8fHcJELirEkM3GxVzKVfzh2B9n8Jdz6nxUkedXNjXedYB9
5k1gFeu7pCCNMKdBxa2A/DUeodi+bcVI4rF+Kjw/HTD8briDdP1GX7PvhCZYqmb5
yPZoM2kq+4Mz1QIcxQrCvvHTjwgYJ+xafVi2+DVb2ddq5H8bN3WPfI8nKD3ofQbR
5l5UnIpWHEiYd6tOdvhuqlaQB7iTnoEjjbEDIIlrOF/xwqyCxjV7fJwvi+jmkjG4
24diVgztyAxzQBIE13wnIXDKjROjMlq+RM3Kq6zk42DrjTU+6p4RmhMhSiVTCUJ9
0BizlIK+1OFnbB1VTlub3+URiM703kG7yy9RQATugPxKRtWs9QiO+htds2UJs2Ry
SxOsDqyNmneJTu2+YqCx9pmSRUl0Azi/OEdiuWqgMGXaXLVQZf9LJXWgz+MwXYW+
bilOavSz7Mozk+wsVB0Wu2N/AZ1r/lN8Xh9kHHXuLz+qSIO1Q+4os0W8PA5lJBds
jl66FLk5DyPXehR22MEMjr3pHzM5+wxBvrLAmzRtzCHV0yZatfu2JKkLCloG9FA9
5f8bgTIKFMensgGmdoesdf2XWXJSZVFvrlyw0f0XE3QIcLhHcVUa/iZhoRUsTd5H
MkP4RNCzanW9KEXB1VGste8b2bpp2EhaSm80+Nj9HjEiozdEKa3CXCa6GBrp1bsn
CzqfXdTpsp+ZYY9gHcSe8ctGaj/mBX4ukWZ09jNGsvme2L7jPSs6s8BuVwiUlIwr
ZDlawQj8gsz2lwuixIl9GycpqC2X5dMV8gnNLXi0Yip/27ezburCmZmMgWlcY8lv
/rOweM0aHHKE57E+uShALNZ9v+MQiU3tbh+0MWMDmdU8HY20e3RJZZH/FzgIJ2Kr
1JhQR0CT/Z1m31Ap5MVp0+5oAoTWWziWZzJIqY/3QO8edtwPoEYwCX6Sa4oIj4Uf
/NmD8levShwV+UzN6ro/usA1xr2lNSPNTvw0uVfHi8o0e1YsC4LMiubzC0Q81YsO
/IdAsQqRspq09uc5T4ktVyFqr0vywYnx0wFjFpyhjOn1USt9uv3bE8eLfT5W2GPi
DDUU5vZmCygTm1+nuTQEiw2h+si4OJNGQOnRsltZdZxqDTGmyAfaAB8UyDv4OKe6
zjAuMPTpYBHqbisrLU3A71/X3kMx6qJN6Kzk2xbDJlgQj6bxSYdZuaC35gvGVo2q
qLSmS7DwLhderHXm+3+vssqqlT2I2dkLAJ1zGWQcE77i3WpQZs+9LyOtu0TLZ+QD
c7EEwXFdExd2T/Ew8RVJzMCVE7+35I2FUOdNrmrtpOHJDyhC3PJy6JZrSvl/dfZk
LaxTNO4kFXRFDeH02VLuniM7gE3fOXAsp0aXLLZLq/oO5Yp/rLWs2mL/K6f+KS7P
/TzJ69vFAwXXHGQshT/BOvm0OLOhtPKGhmNVwW3rGH1aC3OQ7qRp/XwDvIfZcPtl
Kh5lBvtUN2AiibKXS66KPjMskmzSW2DMfxgNt3ak3OdHt3DqPwSCiFd9Lxvk75id
muO+dRzwd6IzLGEe0PL+ujU/RUUWe1eAk1ZG3m/seVCal8BttN0wIo6JqACMnPzJ
tsssuNf5/B2RH+r/yVkU9IScEufT9lgb6cocpk+blRShezdsFu80eX5B0YvC1izP
/aGp/eo9rhoMFY1wL/TjYSb54z/PT3UT1fdlw8K+JDFeOBXDhBT37PKm1itcHH+y
kH6gC33ZB6wrRgGNrR8bDGZ2eHc5CJ8wBKY5Ffdn6vJDHddg7AcTKK7bL5l+/IWK
gsgmHwLAWIgTTy6EIf/isUCxK3YizlG/0ZNkpGgaj4IdUo5T/TbsCvj/rQivqcBQ
K+ZS+KCmaTS0c537us7RyzI1Tkd0wISzDVZzOEEGd6mmawKGZReEXUneYvzSd4wd
4czPm4c3Kof1Mzts0j+Quzfw3aQo8GTVI4Kh2nc2uWKr15IrzS8JUV3h1WzRmYA6
bo1xUX7q9UW1h/xdxS6xyDypQsJW21rjFMDGss/oYiUziyhpUhbnU4ByMpI7OAl0
Vg8hnhV/dLYKOZ7yS6C0TwbJtJiVFBk3XuUhsr+7hmy2BA8u58hedDdDGTdgp9hj
lDFp2KG9WAEc6ZJnq95E1vIvFl/DoPm2HayRYUJuzsOTeMNficJmb8FyRTOo2/FG
lywbR1PGtUTNRU/Cixhhum8Ql0VsTOhiAUZN0sSTgr9QbVNl3PUE7fBSFtaYDZiF
lzrRImBzA3BNGz3+bXCucVmjCP5SghOiA6ehbBKZyNJy76wiozafh0YMS6Dp9Cyw
gsMVUsPDcSqGymfUAljqcYBBNEzTkdKXRs5U8v+aH5UcAIzBZuHlylhprmWl1Mtb
Cjx+rKKAB5qB1inYRAE8ptwUMqytKYgaGFhKpMc3HdnrlOpD5FQsr+w6R/uVCPF5
gHMroyDGKAqusf08k2LrZCn8kFw96ZWiECEuujVn66UMnq01nwVW65MRcJOMh1kG
3uJiQhEyveUAt+EPPVfz4JRN5icaKtwJuvvNqCMwg//PcwrfP6ZAlmF+mRK6S0+g
e+DAQas2gP9MOeWZzZ5b79D2qB/NjpqNk3a/1yqaq9NdmGU1Lg502PWrBh7svj3c
CS5dQOZfkz0DplwwFkqYxwGqltmjPtAureN2PT9QKPAhfGcqBS0KbmBlXolMrtj6
IhXtBttbL8BDG+bwlvDY7wMMY1RwEbkgjVz90FUbAI0EfFMt1TwFyV9cKEivbfTH
kP7TxXSELshd9Gx5OYF+RW73tfIem3RVQkFu5jacEdi8hLEpD1mQTQHpheDHu70x
9Mq3bDJYxELS/2mt4JZGiU5ZbVcmNQf2CbYXqCmNimqUqp2UU1c6YTj5/ANfBMYj
XCeRkOJbRZoMTZ22I5pY+KArR8ViPMcBDRovFMgiSDHip+MOAMDxt7ouvX2lKw/n
sMdmKYUl0sZd+8gWWx8Z2JoFJ1uxcS8fU0tvs5F2WyHPuaKUpNwIwlygq3yVISFp
0hbB3uabf8v+FCmTWxyxyVX91gRiIDlk9rWHpKPXxLHk7mOUuDmAkNxI/97HR1dS
2wIt0HP9SCrVPB59J8GMDLb+3bGXvwOXpHqpeeXY5L7RF9DIM4+sD8VYB5kupUhx
lEDUZQJwRewcg6xRsKAGYPT7TuViLtNvun4MzFaab4VgTDb9Y0vtFKyagNVGcR5J
qZTBaaKnrUaMe8+b+oaM365Deh/25E8CQGGnZTOreiebhSIlG9p0pc0Q+3rIracU
GM7amnAmVuwSrdK2V8pUEflw0qFBBdMJjHTCr4JHMK6P5TSC9MwuE6bq0jK8zyXL
1c0FuOm+Ymv+9bP2GarZP1AsiealN2HxBfD0HxAGtvoN1U1BmLOq65CBwCEZ/PEg
AkqC5eOY+cOfD2DpjAVkVLTGZnJVbN8Aj46tddOtVzB6ofP5EgY3lahVCnoUN29c
nkve0N30l4pYDwW3sV6Y7TYD0km8uiJv2L9/YY7LHxFRXZe9/BRENU5bv7LjGqgX
d5VKGj4Qziu1zO5ZuKLZ6+NlwXjcwnFOu0mWj4XeLKAy6quma6mzUTgRjYzZfzCf
A+3A5J/yXrBS4I51jYNsa0KCCMtnpcEAf33fcEO81HI1HrWwpMw5zDQ4waWD/y7l
c/eS5Vm5002l2vFkl4wvSIUrq0LZNY0SdimOl75L3ooCu/vT7Z9yduXfNOVV7JHk
xHW7XK2cRdqAljmxWkjR8A2BcVT3tLYQs5ZJXzxaM6pzU+LVP6zCTXutnUOYnmh4
72mkTnTFdB7q2U0/Hfs9eHtPrFEnVbWH9clqYw/ymnzUU5bIUT9/XZpAN11vKjRJ
bgZklDJrr6++Un8f57WYCzRkag9gHYRAOL5d7GUKFJDcSYgE4nctMnzGm5si4R1t
OGBF4CxulM2KxJ5oFwYQkaOvcW4I4aSaInc9UT4ya8o3JoS3+NhERSvV1t0e/WLL
60eLkpuUG8t7R3a2WNuSd/laR89IepVZ1aNz++fxgCYLE9VC0gZme3t7ZiGUqiQG
v72eIOdudtNkL3OY1hzLFxBtEiKapT5O9d3jm4KeX83f2EPBHaRRP7oOZmOpZEEe
Wf2lodBaV2JIOgr9EkKgxZiK5yhpR+e6xjrwKzfndZwShQPUH4griwdR0FngoU05
o0rRPIUiqkwIP+eGh7r9xIeqs+NiKoTFbNGsubda5OOn5Gfm/bf2mpF0+ZaHTTiK
8JNG9WArHgoWi++h1lnsg2GIb+A++BGRFu5rDnxqfIcyrEybbrf0YittEMS08jVZ
X+LBMZKgDyxwuw8l6fJDaWRJM+H7t4z8JH66sxJNaAe8zj2V0HT9PRXdsSJQmWe6
EpNIUbvMuUN4ZKQ3Vhz1v5vED2AT3YflMeplZHCOnmAIBPJI0gTkkUSS9Ruu7UdZ
zbEQQ1U+IzNySANGKvc/iVELntfpylyRM0j98JK6cANc8/oEwzZm4Tb6Kl0MAP4B
TaOxU5cp+DxNc7DYop3mnSKUY0B8MCFmBdag4w1Nret088cCmggJiqazq3lBWPhE
PQFxEP3GW5SrgkLMrufOu09m7uF2hGQm4dO7uSot5S82mgKTBtvDjKwe6bY9oCHF
TYi9MdtaqalatpPOBVuG//Yk5VV7Xnt6Nuh4YT8ci1CmRJFKSaIHHV0UXyJ1eu4J
OtmW1SdlYPGVoaTWeNnJpzlrK5weciQ3XpkvUZlt3T42OSlMGVNkXqKAqVXKeenV
nglhWdsVO6RiXRuDPTTp0ao0JKOOrV5Wro40LPJQJ7zZn1boe0tU9GmJu1WV7BE1
Kv75zMKCYz/BSoagTv7ik4SAXJo2ABVf9HeF8wBObinBgU7Z/dZo2GmR7I8EZJri
mG/G5xGqbR+L9Suo5NfwBbFMfKwPmc2KT/YishC9LiJAmAzXr9OyG01doiCAxoGN
A/oMyd85ufUMOSuhAkRtdYInoNJH2tW49v6HgzKwkht/Fc1bxgW84ZDtsWPdxEEJ
PBn6niwUqvB5MKh68gjzUqP90yRcoRDczevxKDYQ26Mg8ZRWk1R0d8+kakDCG3Dj
Q3bWJC+o608qf/eCnTzB07h2z7RD/TxEnb55X6cNkDvEgIxH4ARxQczci8Aj3Otk
tXxt2yCcTWAXLoPD+Tof++C/ATLazRhSIMmjkbIMYJshN9oY0YJ3nQF7CCQzL81N
QL/xbMoc4vea5DoiS2LN1PYQa1ZmghFXrgXOhRUNZkCO14JsX1bdLqd6rMaAhZXz
3BMX8kTpHpz99XcoSZ++MY94mWlRzZd0Y+Hmg8IGHCTJ+fz+5qBYxHbUdx9r/da2
tLLZjKAuMc2lZFICGFoGTtso6+iGWj+zMS0MVtXc+7E=
`pragma protect end_protected
