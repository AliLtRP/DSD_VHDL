// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
Q4liaarX5FI7LqsvA5c3kPle7WWihGHw6236ldWldxfbO5deNSR8qlRbHz9qbhyPxBRWG601KiKV
XeeePzt9UPrkxl7wLcEPfR/BvQCdZ/HDo5Vm0MqcsJGpHYH4V4BMYgS0r9NxLXjT76ZoDSLSMbMy
fefgwu/MmcAowksSSYN7NEv7Zklw2mPTpL5DMvUSoQGgRUtZUvxuQBjkYtx+3LZRzjCkmiplf/2K
0mhyYHIvn8Qb5QYDHvVrjY+BM6DJlQ9Lr7BzQCQ90rmT1jOVOyL0zQNd/uoDXQIwmL0uQ9ZPhQ4D
LogHcQ6wZWzMwF2cjhJlb3o1M+xCmxebIvVNAA==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
txZJ88ckg0+ZZhE/BKdlX1k9Nk7I4yOS3tiw+Mf+j0yb4kanquOoYJiaV8PO65MyUq9IKEXA47/6
ftko6SE0g8r2kdB3yfaoJG1MdvrtpSxnRr41OaEtAgTwJb3GWGkDeaXDPKMD8I6NvKDDqft6oV0T
qjgvA1BeQPNIcR7AqoSCg5CoM7Tu2vCQmrIoUYECbjRZfWf29XKgukbHDvPJvISCWJf5LLM7ztQq
ssbJ68UeowhA51FJYFz0kmjUJCS9g502Ww1a72KcIkIAzAzxazRabFV+wvul/6YU7qoCW8yFkqwy
qW+oxgmdhiTqFTvuLs00uz8hjwbpvCeFQHXjLfpgWiQ5V7b8PI5Eky7Pnq/k/ebLJgsQMg1MElTB
uTPJFNpMzsIFZm+yD69XpgiFV0PV7BwepuoVJg+vg7ihx5uvMmH8gMjh2jD4fHT8nJBdXXMk9VFd
fD6IKNOSyVZaNRaA5qN8D33pYBHnfyr5leVyIqHBxQEHxAeRLeLQ1uKPsFUqNCOVJc7DWIsDZhrr
Xbh47DI3I3ErPKhi+s9DvRt774hJa5JuLlZE0bY9kA/9IYOnzHGcUcieR+GJTRZ0sbOOV6+dfpWU
0GezDJCzju21jC3KPID+vk6LqVznQyurXhPsv2p/P8si9x3SZvt+iyrnNHfq0j+bpJEsNMI0WpYp
ptRlnRy6SK8fWacirVQ5jMBomcUAr1x5i/x+YC/t2WRKl2pbZC17+9kbsm+5UdYsDIlxUMACXoRJ
xM8WDg+OmOVuwohb1IWrI4kxz/5RXZ3TdPyiRytqL2BSdxEeA3id6LrajUUTsG41CBfpr7x8mhtW
k2jC4VeBqgK147vYGd9vIW2xdv3dUI6Ecbji0hVedpR3p+goWnNfrrQ5WBVTQyruPbEM7VfO9W72
Fb6aGuamUdLhLPqT6PDJircY7oV22o4qL5NFWrELZ0n0FblMDun+cnnxFGhQiKltIJ0MDyXQnxsb
ZScDO6OVE45JjFsOWqizypzWZsFZ9QISfbOSO/zUJkcQ7ezPtz4iNP91zkQD0sQQFoPDY0v8O8vZ
7v1IFF0NZFg55duvFrwPms2eEizobCzVRJAyEWlXBK3Wa5E/C1gxb48sDMaImHSLhTDNJLhnP6+Y
K6AAsy1Q9DhPKu3HlUF+oa63zu8ic4YhfYfQmuZdZOkeLjpJ2D9x/9xyFwBYe8KhxRAbX33E6AEw
ONpGF+J3s80PlrYILvOrchor0SxL1nj9G+q8IvgS3w3IZWu5LyyUJx2Gkr9wzhp6WUcPZPMWKdpY
4EI4lgA9zyNbo8rFAqQIOXTu1kw2zBtybz9IDLJou9tcg+JMs1KEMg8QF/h96JsuEAb6rgFB76SR
qsiP5qx4TJzsHlsfQ3Wb1jqLi+Xwc18KS0JsYd8MlnM16UTHSPm1jd47hgZssM4xKGRQv2LTSz8B
49+O1yEqbNlaEr4BtM5aYn3Dg7NIYFevpK++j4cdzzJ+k508Y5ywfi1Mb6QVAxr2oPkdiHqh6T6m
WgnCrMfR1ZddT17p/XlIZmhbGHwfUG69iFRM3+oosCk/wMqnnWMQYgzHHfcGtsWv5eyHY1pLjUsv
+1oMmgeJxpHV6bgY9ygFCtUHgyM6ITrai3NB5rh1CNKFRuGJ7SuNMAXd09ks+c7R1wnnM7dQERho
FgfX+yjys4mJMYggpmsHptjYRiUZUeWqD7T0ymrH4DF5l9WeabVZamxukf2wIBuqikuc93xuNrcN
cv8TtGykVty2vVzEdEzsQh3EphxR+N7dMnmDhadpZW0wLh8mkKr5S0DXK9/vLWZSEK2l5VUIREmC
gedNmrsHnrh/d9wenZkuLSh8yMlSPqENG/B+QCwJOqWu3CPJ41FEfgcgJxjRGv17Stz3MMyw1PW3
0tishNv1XcW/d94RT0/F7TrL0odnrUVEwGW4o2QSLcOexDX4gaDxozcEIAAv7hu3vTzPOEITHBCg
+b0GysJ1pSvHHmn/Oy+vKgtxOsVXb7EobhPZPzGENOLfXtTznoljp+61POKtvcjcWE6dgwOLE06p
SE7zDkTLAGUhtHwMQRiOI9s60DVcJMsdQVWnBY7RhrMBrRLF7b86eg2/m65gyEjzJxdrgroUTwrR
JH3NpD4TVT7poV1rITPK67po+Dv2GdmFFrwLPwa7ib+i1YHQnIpkTQCtjmXjHJHXz8DaYJajDzmz
HoW5tzBwWo0jD256L2RNu6trvsN+0pXqOlOeEWeWFOpCJ0I6HZe0SK8qy1rkJFkS0xOowvUtsSIN
3bB22+IAkNgoqt9hVK4FNIMTYWYQdN/rPTde8/L8QCWEgxNRAn0UfgFdRvD9s8ng2GQ7j5xeMYAQ
yir2Tjcw1PSO8mN+WAlkelYSlMgAB5gEeu1ADvf4LDFt1q7s4IYouLQtRIH7DFzo/S1Z7v66hMw0
rmqU11EDpOjrZQk/MPTXdD/Ke7lvA4165nXdh+miGXBbrpIPDMK6f5SGmY+mReYuT2L/Xej7yPFd
nnHON4gfHRqp8FENAP3nAVJzUfEKPBa4RNQpE3VxM3zNYZsYb6PBsae7w0k+8CpOQptB5/9bXloV
2FTN94cK/ww6AkB0TdspnRbKaI8EjzCDLV5xx4TY/vhHAtpWxg6Yibol1cMZbldV3fN4g3jVaspc
0PZfRMOb+j2vs0x+1YiGgho+/AN0wP3iY21WlDDWQ08RtwCgqA89QjCajngagBRGe/UxGmU7PZY+
3tZN7PhrNHn0DhqbXNkYjIBeJtGg3vcQ1GwFqiMOqakPqpLIv+1BzR1599cisLC3o5e13eKFCHTA
sPys2Ds8N2/0el+dIT/UsPhsYEaLM6nLzM0FqywrPxbqFu3sIzsSrLijsxIldrWg/P6Lkt+8079J
bXx15WULDHjhViZM8Li8R7sorIE1cxrUfaJoEmx6Da567QY4TbMqtw6ql+Ol3UugG+kiDVU142Kz
rhLzMgu4AjtLwXnpzazS+8Wz7gsZ3bfoPLD2FpfJbsGb/IT9vAOo6H2WMvEb8TTGhsa9nWHsRkH/
ITUFGDVdps+oWFaDiP3hOfKjWzavTGGhsJZNo0ODTVxTKFKsgVw+pWVrjNX8ohbz82dXjXnWtHan
Kluu8OC9TPrp4VZTqHMT0muvSl1i0ivYBz5gtPYqTbr89wAQ/dHZjkd2FRaZpLGRblLk6DqhduA4
cgy/ME4I3CqZrmKAnM48EIkhtvj3xwEskc/eG1LFH9mSnGndWxZiwuSRk73kXTdP3aav3Sbs8I1I
V3y1bDCtFwujNi6EXBAh2FSskdc32SNHBRZ1gLeLeAaDC5ps7QSsYEoX4OqOvrxuN6pd4H6AbCwx
G1jQiK7fwh6OkmgmzgbYIkLDRoRdQRrhrhmI4eZx1g3YcMifFP6rvb7eDQsMLoxGRs+MRq4wQ28t
BJs6omrsoAWw6mtU8fK4Rpmh15EBTPanBsdGTO1dY5Iz2mz50W3QwYGyNkPJmEFY8s0l2DgVUHnh
8C6Smd88xvXUk84xUJPGvz4InzWagveONwTbeIfKBwtdTna/ug/RQcupESF4Mr0zk7LgEvNa001Q
M4JPjPPlbGwTuZe2+hnwyeOzG6TDHfRshvaAgCA3HA0rih8JfTma+poydmqJY3+xwqS/AlP5By36
q8blo4f6IKvtkvfyOPZAEL2tink46TF7JdJG+m5u0oFcIaLtDMi4fyXD+UGGbDpgJxTMprXgooX9
H3W+jryzx6cG+BPJsW+cWO1EOCafIdmFa26Jwe58z/nQEzlrMOYLbwoUtL4UlflynFpaUowyUuuz
k8YHrwcQqz7LyONN1r/WCl0aAYHmW5uYaTGVmOCed2ZBPMkTuMGc/ZGYf0jVUxScm5sVE5nuOvCi
l//usCKVAOwZ+JRuBmPwMy/wfLOca08hqW5gC/BlMP3d4mjsw7da0p2FLnLK89T5pRVsf8CjyRuq
7yEljs2W6SOi1vrE5t1Esiq1MRP9ldV6TZOlM3UqSsxsSuJDIyYG+wZbxmG6LC6ONVjJ+54jpQr1
9e45ku7DxDh67XA0PhFB6z6MXNtPdwPVLd/IlGx6pPzbH9cH6BPqtjLozn1XHx8L7IZswkdR1ajx
/nWKAOxNBh6oQRsiIfXMGPhHFYv1C+YdKTeQj7bUVUi/HjjNmpI71gySI9p0H3E/9CS3CNDIda7+
xrx0lcBofN1zh+ybFso8pgCtbBB2jwooSLqToS3DUxiCBELEMYnyVwp8FwR6ClqV3K1cr95XCXxo
09y2i3wTIDDFqUwJV+nhUgoMCKz7/+QqyBhYcJS5md1XnFPUgepH21I6+VV5+q1ujaDdad6Wqtm2
VGM9P8FzFEsc+9D7i6Oa/ARFIh4fFq79MPKAVYVdEyJmPtPvvCAn8AYAI78UwaB3JBALwXQLYxel
ZeNf/+PxS+cSMxEfMd7rQWwXdfa4RXUtdoquOBejoCxoObzSmM4KUAEOkjTpkTKBkMuVIEuvE2+I
Vq8LBrDYdDCRnxYGNQaiKu4V441qLaNQLw7UtSf3a0GdXHATWAAwU2nMf6W6os7YCVbJapGr/kUl
vBPRGUPegw/NRtEXPz35H9Xz7dHH4bYMvLkemyMNJ46VxgeoLn0loaI5bBj1129d7mMRBFUoJLn6
JggwicYPx6hj+pmZQUk13Am6U+9uvhd1X/ssl24UtNmzHFrEzrnkn8qj3NcP+tFWgPXGojXRLRJ0
zBmQ6ux4/zPvF0o3RbfJ0Kc9k1qneL3GlGk3CHLWdEaL9WwzAmSr3+gl8PJX5AKhkarXr4gyPzd2
2WtVEtQ/OUOcRSSNeXNiIq4bVUpaDOvnGKU0jaF+j1HohejmjseQ6IW3x2eWntjqTY+BBtpGKL0t
Wrtj6gfUZks6uKpiKM7GA3axC81V5uwhGshyyPUHff3oVkIgM79TpnW72KZpqA/jIQIutCtzKhiy
od7IaPvCe07KJ3jEPsXbCSCPH7cfv/BxnZiXSurZgbpb/zUpUUq+xmPxnRUqTPT3sutqyol2t0gl
ZcS4MAKXe6MMls1tBZmZ78+PgCS+yd9zyo9CJ924lF0DFmIYttqPwwjEOWmHzTvdwxruJ23uFCJc
7Vfs/20ntwI/spZWvZ6xpSwb7vfh1g8+NZMGkEuR08drfzYFHLEfeIoDzNW/iCDDE4YCcPeov2jL
0h6jlvXfxX8CPs5dI5c10wbX2wZnm3cVxaLqVc2m+giVwQw1+PR/W1YImA4LvxvSiuk16NTFqAy0
slMOk6Jg0DuosQmH2dKrTE06CdMDF2XECpcwE5ttrj45zqgN4PrjRP8c6H3OKrF2QZG0VqssGcFm
CU+SG20F1LbHbAu/4zac1hk5kuMkkxA35KksEwDI4obfRrAUHDBMhdlmNBOmMAyFG6wErhs9ROyH
Y+hqYE8ZqZbNyvoaej+oipr9IuVS8Bqf68aS/S/ldPg7/dS2DZOQGLFC7pG5i61PWYSv6I/Xgxtu
66yPbxTk6BCox94V33p32rXyp5f7m/SlcbRdFqIzrmL5EcwtYdxA9xJce7hirz0mV1MAtRqiUuXX
ygqtIZXfezxBDf+qcaeYhsJJs2UosEA2MFwFQO/valK6dOcFBVVCrvdi4dPQThvFNrrqFIFAzpfU
quKPxw+MKAgEZNxbN8nu3G5F47owHtJ1MoHDlipbI3PCgCglIpRLUu2YoKQTLOLoeLXw2HN8JuTM
p33Xiiy74zaUMrFcjDvkv+GZ3eEwPsbc0IXLaaxZVN4SmiTDVTTKaHuX5YLovPIQf49fRDN68rYG
EAu76RAByFeIB55UYOKJLMT3Aki3IkGM2fshi+xfRKSdUBJVBOHmzP3SbDHcTLaULOVTIdyz9zp/
u+KC0qWC1R3FLdOsS4og3XMCtmjaazWM/bCbLEOkxaf9L4QyF8thFWFt/J1EtHYTV3Px16ifgGKG
k8taOCVaphimuwy5PaDddMH6K34BI11SEh8OXjIbAP7xrwNK6y7r6h3lqQyv265PtLXNskO3zSvv
2H4cvJohbf4JY3GawgvK45Bu8cWG02QpaNQ9p3tb7YCjRzaAcfPNkGPMAKcfzNSg+lN1n2rjnDGs
Vp1Djxtmkj9Y45YXNjpDBMpzKgdRVZoRdY7temHbvraMWA9Y48bisXFIRwxFl8m+u90p78cgNg9q
HI8pDQ/1u1VW8/8MIG5UXkoPjGizl2UsWsFaLHHLzidqqoqNU9D97550IW7ff3/qIwcIikaMaD4H
w2v59NL7ZjIcofAUSFYAhBe4YM7q9yRHICncGn/jKyC67XKWN3MlxjFNN0rWmvcqFd+L6he7BtBf
ug1bouWWPId9n5tjuun8TprCulavznKxFL82EJIo09Wie/sC2iOhpdKEeReel2qlfqLimRCrBFIt
9CDA5wrl9YW4FUiGqHMxAqYekxr4X+67WHx7JSzWCbov0+x20xMX2qKEBck56e+mLrL6Gymvyj65
yoS5jr7ls14nj9q/fVUVSLaP7pKCczpu+V6x55w1McPv1L39ccNfaVHl0J9SFINwSHYi/aNkXeL8
YxqS3UWzWCOi3f4ycMnkFgpxWHRHILqSWpoqGIv0QZncrZiAGx14DVRTIUklK81efl9VTJKXyo9T
pLLabw5tMCWbnyG4+RZ9EneuW8W60Yv41dXbH5afHpNbACIsG7oSF40aUOdUedBpjOfUo6goXwZi
BlGn/ftmOEE7s65jtH5dX2yU1w537xsaL/k625KBkQWTJpk2mIylZQqHU47Yl3p16K6OP5e5UgR5
h7wU63Vij6ZgnpvkSL+WWM6X2WrCnXr/iEmp+hpyvSUYKZOntkAFb1yUWfY664Y8w6+JClebOYct
JkwW4jy/t7sqgw7qPY09cnPvxPCaxd1pD/gDQ2hx+AexGE18X61IOWHWSavnjp9WO2xSpzdNOObG
/N/XU9hFlQhJrlGO+45kKS3BV0hsuNd7uBg5RwP/ZZ5JCuTNzesuXFZeY+qrXJRp0u9xLF/FPZ5G
gY9DhVC4bYbdsjczpSJfU5Xuqn3aNZRlZfp9uUZQmK24mNCx9ZOZKv3x0eA/LTCMgIzGURsuI/j1
8EaqI6ydXDEy6wstKO+rJuPgujTDj+VgEyuKwIq+iFk0aw038ZY0Xh81TnybFCuIGsA8DfStEu+h
Rk9GtFVYe3AIsmvBdXSJ07XC3S4zZPNOsoeupTqkjAR+ibfUvmlTqM5Vc0jW9Ksym9kPSpD/st6x
mRxUPLAuyL8Bm/UaQ06EhaUKEC5+79H4Z8n7GLLv+XY8fWoClYVD9Jl3HOD71AM7joTz4BUpCMre
IIobKZJam2IyxI/OLCLBgVhz9cLC/eEhPRdnjT/+oTXFQp83DjcatgDEJ8o5EQWyga6G5EYCFq9H
6ijrSv2I+sbx8Z7MZpGDdCtumyGh6lveeIEYjY0DaaSvCuMcunjVMYRtYztYdr6T9SN/xEJ+Q+Q1
Wk5o/VntTftBWYAjpMO2RM/3n4SqOheI65BA9GOqYfrS8y7pRvTn04DNRJR5Z2AUEeaPmDuysEHX
zNFSJMN6cTMyiaSGF6aF5MlkIj2VxL+gdawCwEeSNbLFe9IIAWdHW9vhwQ3LzE0brryepe7ZxidG
g1aGlKzNUJw3kLKXKp1cMcbLqNriCTpPPVqSkTNc0/2sE8/aSC+ENo2YE97juwVjxIp48OyiC9us
zP4h3jUFN0u02TD93vUSdF/jcPuDOQVirSraFo3MuE7+qI0DhAEflx8DPFteahTiGUusiYjHqEId
5ZfIyDz4g4HHpdge7sXM3vEMcRqkC3okGriDFlz8ArYMMWly6e1xMu3SZ0ue9m/hRwFGv36Kx/aR
PdgpchLkvzTKH+bCoABtk2eo+lHksPWZWLS5Wr1h9gJ+HD4M1RGz8j6d534Z0ZbU0ENXHjuSCHRf
WOiy4s64K4htm8jR5Knvxxs4m5DC/5dFa05ccXaC2/rC6Wq0jlu7hLvHIk2mJbv/WpN9JKkLcfj3
XdhOOcWD7ZWv8kbW+LYdTXypqx1zBRS07lAaNRxOQCAbzc56pC7rkRuYsGiDFDGRzdnezjknulaX
2xydMJgYk5/GEKTRZqHKUH5PvgPAOpxpZkoopxEoFbUj2Mxqql8EYP/Q/h88tL3FYmYzJNFYBN73
jEJHf60L43sa0jnj8CGfXYMDVU0l38CoQZC3F/DjuTuswvfdJNHpAW0+Z9/egu4DF/2O6HGK7rXo
CpQ44s4EEMstC+Ie6Bw0Y5f+xzctz3tCON+6INwM6Y3l1HTaaUHLPa1Pyn9GXdeDA4G61fGukT31
B810lxMxV+/CgfIaqgXjr6YQkVTkfurLfJloOfLAA3ZNJ6Z3yNI1aE7wqJLimNm6F2RuNCxxpepN
fd48zMo1DoefrttoopeXE25MrgXGB2RwWF5FhXTEKvVzqbCda+F8Onu1372cGRNIEUvCWmU899Gg
81YqXEsx7UmGG68TkoaW/w1A5ZEF463voaxjtlpetiuwHoN2m4xjOA3UxygQeZ5ycpuiADRApdWg
e8nQlAWEi/u6VKIeEWrWQGjrRaBhbR+tn2iY6C4VTRJ35fI5/0D1KtjFTSfiw6q4EpkiJFL5NLfi
0M+TAO27lKZu4D+3FsK8qg8AvIku3nOfdSEt8gtknvRyNSl00uJ9VdVR8309pj3kB3PLbYb0H3wo
LmgmjQfHSlBYHn3fPsKkuGE5YluKfDblmpZkWfVuauQ5bm8D9X+D18fCVfigJTJen39SykkDMwFB
VowSokipnTq46oao4aTDU/1a/2oSU7S0G+Y9UlHPdMe8AStGeVDmmf2O1E7Czaq45xvSSSik3nRR
Njl19QmKcVSnpxSLws4OysRXEzcvqRXwyWiqrg==
`pragma protect end_protected
