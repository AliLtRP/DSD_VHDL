// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
U3z7/vee7jVl4apokayv1nUy/pwUev8mv3bqdn0Rzkw6fVuiZBRx9TQGpztfgFTsuQqjZemOY3BF
o8lQEa67IbFGUT8JQT3K7BVa0bYTH+JHomNjDJS5ABLCin+FoDovnJjCMTAvax1ctrzQL1rfslux
a8suw5LP+0g1p3XqZTKf81uaVenXVdo4A0NgfTWzKF9AOwvODATDoOYSPNpmbKzShgZPRc+OufLh
yTGFsS+qFbbxl1Q9kd5NaYcRoLPRNJcVdrJJLS/lAPJ04XcM8bHT4B/2F05Yhb74+IPgOy03OovR
rEYnYw3t6tEpSxeknU/UOQjuO2n3Agr8nnfLPg==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
vHOGADdrZbaI24gvi8GwdDC2b8W4kRe10ouhhsuTiDYVexuBPFzUhMZj6nDfXvEwncPvd88Bq3LX
lflAzRHtzmELHetRUZz1qQqlgszzI4DpR2kDbrFriih89XB/V1XJ5NdiltsMhhwRKW/56QzbX/+v
laEcuFIiBDWV3/x1k+EscpNQqDvdtG50mSwsEmKA6msv+S6MAQHl65KBht+F5e3Ugpy0Be3/sS/Z
5tOILCcI777U8OTBKpJFDwUg1VYCCSkeCzqQae7iUeCQ6mC87OMWRi0yrx+qabIruwsqojveSMTf
hHBCU6ySqlH7fYWtzEQmrk78DLxcLFCCTivM6rPqUjfJhqRtd1kXPdiFUWqxs+xPbIunAkdmQmgs
fYVEUqY+XYS3Y3tNoK+TyepGXsBdulhIGQ6AtbdS2uPZAqPf46TX/YNVul8d1KxVg3OT3DpaeMfc
OpfAkaZJF87RJ8Qp4u48psxzkeHrBrcuewc+R//55jSfque68fA0edNrjKycrksJIiksHDkhruG0
JP9FHoNwvzhoeq6z71a8xXt1aKjA9ssWYuWew8YLDYvkRv2YtoAOABz3N1vhCaV5GOKMQLf6b0Km
f39iJM2YIWSOqU7cDabSlOiqTCuOSm3ZB5LIRQNtRb7/5fTl7MkQgZp0B8rZnPUma1hgwOGV+3L+
0lgflAM/Jk3fm/lxVYsc7UjopX4QWno10uJxGMIrlMZLRyUFlIBpxd9yWLJKjoazg6XCnlVLweKG
cOVo//TYjCE09wJHu26II6JyX7vSCHscZxMHFjNhh14zxigoUlZUnEtVcG4mX3bygP34/VqbLvwd
JGSieJ9AFqwprxqupltUGTh2f23vo8rTtpO0MRebS1nZzBd7XuZs2KLB9902juEewosW2EUkT5S8
DnAEVcaeNQZdM7aeHeqEjDYAE3wMhqxOg5/JbKCqOevXgyH3H0YsbXiqkBXZzLTKnTC5gVE2OVVQ
4j4eViBAMyvr8284+mCIzE1cGtXrX9t5mGP/9MEsUCsdN3ktZiC3v3LwnuEK+eW7TRkzGZ7cht/h
i6iwRgP0SFGB2FrBdxdfazA+2qwFvGsL3XpDHL45j7tn+6RJmjU5zN9iRMTJKC6/uCcmZm5pWRXS
DTwzeinVKI9avEB2uzb5n5XreSjvRgOhX97qq3DDDM/alLcy53Hl+iBsFcgZVvyxE6Z7iZTXaPGV
nUayoyRoGRcBdji0ydsDciS0b5SLHaiSHgKqR4BoTVk8HmMrkvo/q0/4PD9CqmTvGoKA9nLWDw/n
EkzfZhAGl1K3BEgkhuXsKPFNQJuVGTbl9i4LQUSz0xQs53P6CEBgvfefOtjxArCL910DjZJvsY/z
y5dupuwzVlBk//ICsDzq3FaOQ7NTIUhy+XqmvBstkgz/LjQvFEf1BA4J6vFU1rCEtZw8uzpVNL5H
3/Y+YJQQ5SR7zS21bU5nM5fpErGFhMkj0m2SXhvieA0a2q+NE+WcCQ4b7PXPug7TNzZtH10HZVg1
YUsZpO8UPk+rdy0e+NYSrvX0KlFQg+FAbzO0iLiKJlp3oJkE5J+wdD9mq7+VTyk0Rc/dffs65yln
W9n0NZLu3nWbraSz5mJMfhlNrPNQRNjZVfJyctv0OB032H0ryx5dWPSwuHCIz8CEQSIJCBZWFKTC
8Gbdc0tqtU7EZBFRYHKxcy1o0VZxLuoReX/l+kVMkYf0DSNkl0ebsqGQ5IXHHL+ihOXr3+4gxqLv
RxipcunNJbjwWORI6N0tN3oHSNC2JzTvdQnqxz58quMeqiR7Ou0oiSTc+ajjrVimsYiBA2TPOI6Y
f+UEPV8hlzIpbAon39TTMywBU8OzC5qWpD4/9w30viGWKJk/l/bRLRMXjdw72kP7xOMl3K3mtfhz
/m403AC+T6+QVxAQIx2UCDNHUAzA3WidGYi2CCqnP/3MvycVH1RCfmwpKCdsf8wBNV6OkSj+wOET
XTdt6v/JKnNXVNvLUAsZ28sHxYt9ks8/YN+J9ed22NSLYeOtQfUwvP66WNDQzFjXpCXwXqoQ6sSN
g/Wgjeg6heYlVHkJLp6h1GQUqTs8bb9/b0akKcVMaKwozDvvWkjN+z5fEq+5vK4MlDb+bHd/lLnQ
bTIb+vWk30tH3G2TADTIabRgs65So/wY9xOdi3Na5xEHKPF+46LNgkcWqzVeqd7SCdsrn5j54tvh
73XJ1IqFUOIzCC0QY/eRzSB4Uj5xw+LPHdfIwv9lDQVnVvTLOu9Vp4f4DZp+imzLtGOqKtL/+RHQ
viyEIMgiiLNIpsJ4im3p6TTVdtZrhBfdCYPhGQUYorY1OiSANyc8LJpZ2iCDZAl2HAOTzwy6p8Fl
oEC1zNTk50n6ggP8oLNT7v2lU8pTFtCVNeNU88kOHACzMZZuPFOQsGs2DGdaxztqMjWYwCf4xOtv
dRn3KAMMq8+o/ZjR2+beX3RwCswxJuJ2EjOhaPdDoogn2OuAvPyEnPtbOlgNHTOnz4OdyrRa1KUF
Os/C30NMBao+lKTxht+tKCGJhD18U3juD4u9zh8muLb8ykZO6HSLdjoVYTPbNh2l2ZKw06NL70Z4
mcZB3eUEOrMgT4OyKxvZo80/3OW6a8pUoLpf7cnZT7uPWVGGlsPXgNMkEESf6JvjKOjVesHDuNco
noFu0uZJVTdXnmj5/JmlGV3kpVsSKcr0ymVYJfsY1JmoNjyrWS7o0P/pnfPhWzTeiNXU7K+rCcw/
p2RxwKotv3l3XXUjf2Sviu6xPpOaIVOrtNP2o064caH/lfO6rg3ruzadTToaDSlGMM/5TRYCQeHk
E3XWopb0QXYx4W3EdzLeoxULlpw4LcPEl9iTnYdD45RDEF7QPrrGNVm5wZLLtVKXQKMi+w/5rRSg
dh373mAuLRJIS9+ti/BTrhD7DZ2FRLG8MaMDX/ll8aiaI0VI6TUwoP496Pp3acLozt67JEmcxecW
FPrurEVqrPJKQzn4ITw0nviVCRAaxLxue9f6EU2TUgFsxswsZiHIUN0TjvbCvnOiERyT8JPVHgCl
vvbWvfPtaTYrxm1T98qyJ2M6KAHPnNX1hkJmjxR7zEbtSa57cMTEREFeMucv5kTwSQab7utuOY0p
UFUrYKK3/99WF3fIp52+5bw/SF1VWKXCza86f/3Cp0uk0b5rGtihqsQv+iz/32L47L+1M0lUPXAe
UJYzsLdZGV7oobY+4+QSnQzAyCETKpjgrz9uD3w6EF28Mm2aXfB0gXggBsaN0Guy7qrMFKsgUB1U
nsyS/q6Ud7JxcPF/OnnF59ld6L8VUg572RSvA1l22XLwIc38Jf7UTRw/JpaU8jQKuZNNLXuPd7G+
PBUHqkLAb8vtW6jfYF/s/RiJhfAQfo0E/HtDd/XzdXOyLf6T1iNhV2nwivhUjQv/gHmS4Mrjwmmi
E31QnQKabYiRwr0TUxq6lDWZ3Jc4TRFdNvxIdIux1Ll4zjQzb+9LcY1Qi/hqxEVQBdXzELKUVAO6
Qtjifa7I5Q7vlff27DoUiepgGR+eTK1jGSznpvql+bGTJGwaa+3vNa4qpkisSAH48Ruo4yUK4sdH
SvfUCmy0ilu9bb7/cX+hAEAf49jKgyn/Xm4mpOzloEnLEx11C8kalZV39JaoL/QBlSv9xo1bgISj
XAQkVamM9Jh0lBvnRYI8aRSEZUIXlevLSUKPhZXvqKC6TObJHTIBKxkIzkKGnqRFm9w2G2Cz6BGb
RvcSN26M+Ln/16laPt2R5BfG3XEaVsDhMZ6VCycMJKAD88azbK08OjNSD8Sb8MKRpaFranep8+YG
v/RFjGYtO9nDGwCo3l6KkCJzlTVMA74B1bgntaXvhEidjWdymF2kq3CE/WCuux2YewtFxbr1ga5Y
kvr0uXgDR6vDtTEu+XzGrvTtfkFzKKUF1iNwerWkVCLhiKV/r2qEyDuEGAeIGP3OhXmMdQE8cvM6
4mtZvlrfjTmfZ9jU4uv8l/7ttsubMWeN7Cd4hYxsDuCaljXUnj9Rb+EpNoaMbXFzo4oWElGFHdx2
IDsavN6SdtQMI6VXoO6yrERFBAlmRR9Zbf5LAVYIFpkzkys3DhBlGsZNmxQTLEg703m2Dp9h9Txf
hw3k70bGRx0RfQ7j5d7ABj9j1HIAkvO65+URGKSdkMB16uQ2KP7zYCKsnH6OUk2QG+uxUahbzLjQ
/sStYJZ3P566AaDNvDSoYNaKFJ4QL+CvEkMhddtGKOzh81MkAPHlBFbclPavpsRv0DdtqlFbjZC+
ktcIEsWAvwEfYA7izuunKurJ8rqRmdGg/W+Rv6ejKnX55NJ5SIOUXQ7IwgQ8SS0uQqjxXSU8XYg/
Sb8GFMqk99X/ZhH8sO/uiGVtqDu6EWXfto01DLmcuSUoRfavk+bl2RhMmDiemYqyYVpITnhSDfUD
rtkRIYi5hXCa/9QvdwprQ3PZNU5Co7gis2UFF0KSaSamSb57m2YgFY62Cq3SIOeNRTYTdTkDlbev
tgw7L2fjD3RN0GlyWKUTv7pngSvswQ0syuC4bj0M4vsSXfrdMFtLaO89lkye5J8+R5iAN5GADgoq
ItOnC+cK+GTdZLrOUvCoQ5L1CZ72pVXikDpFVlgSX63K6J/ZdO2SC6qcFkcaPPnx3C/ZwcP8m1kh
BRSLr6ueUWywiNkZVVhoM/5TyQ/9MnnRkaM35H0vAUf4xgyhWGugLzGgsRJCa/L6osi+x+LO4Nhc
TTC3zXqSRwvWdxT+vv3XFck3XWuGrk8DKo6qQhZP8w8an1k/VqjG3ds2RcqZXqrjDkcAFtbCu0Fx
kBxM/oBcl3LLEpq172SZ2XQRFUnBa3d3qlh14ttqV/aaml7Q0UvU7nzVJor6GOiJVjxPOv0oHOqO
9NzGUUKdOOc4HbAj+6qpmamxSxsyMSN8hlMzRD8+o4dXGOSQduJVfhq+bPTFs9aAhweqHiuhgc7a
m2cfBu4txuQ5qvVqlFT6q90uJ2xeJtTHntv2RFkNUxroQj763+AkZMieHLhCIg5UYRUHpwp+Ukkw
ZQxEwcH4i4yjDsvrmwVPK3tu/hAexhEZyN7b6j6KmsoL3qDpvH3sEngYzaLWlnGQsC0Ks2hUTkNK
OUUsbsBXZig2QabI1W5ew2Vyp46dFOf8LAE6YcBqwMOBoIWoNmqMLr3C1NbGTSCce14no8PnLX3n
vFxr9VKmaOY7ngc7lSrtn2uwSd2gDPfkvt1wTR0D4TwOD2Vvnf7cWq1YbrFTuVUG9/6t5eI0mPi1
T/S761zpRMwscK/D8IQ2FmjV8pzq9yHGaKTWXyXjnHG3HYeqt7UmpWL1JDtx4XCXrjmBEkY3ctWI
mWuQqCEfhDYIJD0C9/qAofnPWc1bJggPqjOHQpNzkjB7wehs8C8ur0FRkFmr/+fZveJq3+ESt8R/
okJZ2uWptQcNCauidKBpeqULcsI/md2Wlf4P5LUoXmjRfdZbdWGAJgLbcsnv0uS6KHkP7F1UnqLh
r0qkW9aYvaXpXgDDLkph9tf/9wc3hKWr4ECs1fgiwgIJROwO2n0FbSGQJB7MtiFtG8xnsHhfaxuQ
yCiAJnDwrB4BTHjcBcp7AKP1uUcDUljo7HiSkBmtgH/I6BD9uWt0yTlMrdTLUbxteFmXfkKoxart
JjrNtotMWUI3DRFxTkC6eGvvAJBAXFZshRK8i0AhZ6DzpLSFBzAxzW3fISeo3FgquojCeOPswZFF
16HxAUuLDxJungXe2DKojDqoffa9321PeEnC8XiHYxODgmH5T8dO50l4iXgxu9GmsN1vl5FuOVa7
JGs4OWs9g1/+rp8EoIj4aCBKPiTgqTqBy6BFagoxHWZAfa56klOeQwiBBFN2QJzPP8ccN/WJh6fw
NWZEhesx6HGZ1ASD8C7+UW0qt9aIEDR/7mt699zi3ip4mXnzAr7tJMQ3W+dETkaFScGkdZ3mcz1P
3mIW7XmtSsS5/flpRxZElQOQRa2uDk08RwfrnQO4x1p04LIWs4khfLgwAGWLftTF9PjTWIen47Pm
DDSZjY3Uy521Q7LFjwrKE+N9GpFVs/MsVCxU6PCpxmkM3oTqVyESftQqLppbHZugsz2sRAjM6JAe
kow0Wln0OBn5H/gx2GQmJc2KXI9snJFtKRPfdWwgp5VhM2XPlrKL9E9Zh+7NgedrYl0oVISs2llB
9BbbLX8rLAUJy7IGSq014ZxlNfDworGKrsPQ9aYErKWbXBLvUaibsL5Wu5SyXv1iwh9aw1hF4m62
GdJyp16UHJjt4AvO9p1SO/xc4kLXji5AV3n/GTISoc2aDC6emU1z3HFx7DdeZIBlO9zeszpIxY4R
Mzg06uDhrm73cbo/6wgMiSOyb7XcIj4/HS4iCo2t3W8Q4lBVIQgcn1gnJDDzxsYAF+HOHHcApSNK
0cHtZPOopVXH6L0NjO2hoEiUT89PN8YeLG+puEDQzqlc1YG7e/Oqkb6LgUcDTa2FvuWXENkGPwYV
55g1pPaU5p/lof5LTUYhBX50dSS/21m7uf2AlE65BrQtxW67Bl5BdrV3F47TTicLnsDSTfXwgSFb
+/SXkikJTZLKE69u2fDrAEcsTKduPqVKALPOtjEQHRS8Luu+jba1DgJy9dE1zU178ZnvBNZpxHu/
gI9VOORXGPENb6Tn40KIToM4rWKOWmqzPtTgHwDuhjMTyyWIW6joA+viS40TQ+ntPZtJ6HLxasoY
+BHKf2nkH1ft+KJi4vbCQuIvR92GB7csq8DnpBA4G/0LM6Jfjt0mOqn9RdDiAzpMBF8kh4W1/BO7
Bpflh4febI3suvkzOE7oHmlGTMDjHWe6ruxHnEc1G3TF/oe9VAQYCZH2kBfdaPE3uG0Gv0kpRfXB
innHA7312LtgD8Gg082+xTyGi+xGjK+85HGoAPf9px71MBXJ6/3QkKsUdFeNQEEEiXUxH3nTVw5Q
6IB/WePOCllzbgOsA0wNgdPcIWaGiXf6yeBVARYFqZmSISJIfZ/nL2MYY6trt+mBAVx6kqbQHUNd
HeqgYCkHIBCWUOuBqkT1BM087BXSmtipEJqBKJq/UZmHOnr22+JRRuukfisK0ktVFIKfhzaNnsQ5
mpkJ/M3E9STRALVR6dATBfeTZOiUa3QDHgYrO5pKLA5j5l1svXyDifxIfqp8z8NioUHzoPEZP/ZG
NIVyxU+MuEDNutbP2vAOhXTZPW87p+dX65CopiRY4gx8PEb5IwmAzgJtRXj6FAK/kqFW0p4XoIhG
1a3EFEGju99bWk+mTEPqqN2W4uQE12qrC82wynzGZLipf59/DKRhhlcAxIpq/TIKNAqji/M252Zm
dZIFeKgNJ/UYC82X0G635TrrfW6jhJtYLQFODfidy76ICzqGrZkm0Bw016gj8ro542qX5Sq0LG5Q
0toKaKIyj+gyxnhOK6ji4O30IvitL2YbiG8jkeT6G/j7GYjG4hV6jX43dr/4KuZJmXaVixRIWAxl
miSF99Cxs4NF0hJrwdAl8Q0xUP29pj0jKs4QEuPBMD1Jlu/kVkgblM7mHPtbjkMBI+uWjIpXVCh6
pxTnsShJOJZPwEv+wWNXJeE9YDyhgyEHbo7KfAxyFXd5QL7DxOxv24H8PQAecvlnZQzsYTgKsIyw
gzpNEVdmwSqHs634yAsD+0gybpSJNUpicZYWfN4oexZ7ztbBXkMzsi5E+9JObmYICvdhLMsoLttD
EE3laNTWlbjNLBo6Oj+6VBtdt80cRkPPfbliCLHyv6tBwzoR8cFYNBKdU67m0FZ7KRFMZiX1A1tp
DK0/7AVbmQpaMPcFuWCd9CwQYzCBfokq6C03Q9a9okmT8EUkme2pGVJy/IwC/AphqbLW47hUDtlj
JYPmVHj+RzyJFZkgqCXpZ/VlaZGhq+XZc6RWdEF9oMhfX0BaDOBeFwK35ucUrK6ftprtj3fQkj1N
MQ+nLhDsg17/mXdK05t5iBHcyNcZ0MTC9U1/UJQ9hOtwj6aoyFP+g0oVSJQLeE55AGv5cyWb4US0
bRBkH6PPUvlNHjFTtWPoCLzUqIYgfqh6B8hy63gCr/IBYpGPxRHq704omYNZMJhL57iNCwXgEG7N
cLpW2g4xPV8FgzBG7eZxFfDgQOuqq61Y2UQZ2/ziWaprFhbu/GuEbWPjOSmOea73r+elr8qupD63
FX6Prgkhq9yYOAf1LdUxCisczmB9E4H5DhkW0qFuDzTrsvtIJySrwp8a+l8kkGk62hp9/TkwHJlZ
ls3Tijc1fXQH47w+yHBZ3dYdzTe4PC6wsJWQoHoVfAGnMU8uH6xOA45iLBNayjqITvWNI4P5nSQc
zobz3mdmryeHfZXhS5nnBFmONoSUhEm/Beof6JpBqr1S7DVL5OWLm4Qmq/rAr+2bh8XlaKlwpwlN
A/HyddfHvQ789GaZURuK58AnqpFdZwYhzPTnjiihyrx21Ep3jxS8wkgTIm7rc/5TNw8hB8fRX2Zq
k1XClkXJZjPKL19tpTqeuZLaJX6QMOEiUDGH0YhYw0qmN51XaNZKyxse5kGo8g5b/sfLj29l92o1
ymWNX7XcIFIk4lK6TZYmmcg0j4S/JdGwtz7vrtibgoj01BEf2DUK8MzIte1fRZLiTz4y8TOE4+Mh
oj4LVGoDMEa2UUHra0t+wUMsfvHYywp7WOI+m2FEZw/8S2J3qegq/NNqSxY2hzXMb6WsYvp2EXVn
DSz300FhTpbRQQPKqnfhR6Uk4JJn8Nsr5TDqkzspilOuFXcwWzysc9+fo2hpjk+KjRlHyGznW5nF
M1UUmZV82Qq0LR5RrmPBX5krU+w1N+K3dghvsyUj2/d65hJ2ZQFJJoa9O7mUf1OcJa+jAgGel85y
X+aRNthzoStZxlNV2PBXJpvNGhFPbpBqflFAR9JGz4efVomJQw/9u7G6tPCYCre+d2nSMTz57zSI
q+g4iNFdoI7J364KGcrhWPELjxnetXJtjt9cSq2p13ze7wH0JnOpYfQvMr1TnBpx6qqOn3KV9yPR
sLtGLGOpmbhc/voBoVx5EjFSVeiDCKIvW6OEadFObfZqm3JzWR9SJNkFDaNQEi9X7DvkfmQ1/xmp
VvlvijDqcw1l/WZNEZW2M1zSHYYDt88AR11o1fmJFjaHgvuyRgBp1bFAKmnK2kSEs4NDKcSe4nyA
qnCgJiMJCCvqhByryABSQwwG/62isoeZLS2+ezl8GAOwKHWyrgDmJJBX0z0RkkMRCtM2PLyl5/vG
1nMS2VySDUx05j8ghLvLHnGgDcYyUg839ZI1YIMrWJGG4IvVcKRa6WeHPU7/P0fWto8+JAXEphHL
Svou/xE73/ri9zoV4JUIMo4SIgwFub2yYYHqCHLSSZOUErT7k9fmFWEXbVEnh+3Aim/9CVdM8/ze
c1W4tIcNzf/FMIRS6L0uo2GcayLnU59/GeWP+CCXBO/OwLKYnAcq484pLpCJzAsxLKUqUH2MrCgd
jmPT0mnysQbC5p1Zak/B/6qmdV+Gmb3kw5nT3x94rn2ERDi0dZ7Q7UJGNukvvogH3NJUHBwUtBq3
o7IeH23byVdt4Cvc2zEbsV6CG2hCdBM/B+ZGIrfThhtHm4PKelSgkHmDm60f09KWRxfpmmtpe6/I
UHkR+ddAZMeV1Bqk9bd71i9KArpJ0OAT4Bf9N5icBj+0VGQ2TPlYRPsdIHR/f3toOieUH3sJYqMT
IIcIyoy4BiDeOMjw7tTa6l3ddrDyrIruwI1BjCMn0o83pslNWwqG13/cbktQJQhiVuFIjqwGj5cH
Mqmy2Q9RI1RKg9ho1pqGwFQcF95uLr0XrM9zP4THORepy67+w8oqS/CBF1ZUORsm/qBfDHI3+z6E
5CJxZv3VLiia52rMos2LxO45GPqz7I/wPWj/FYR1Gr1lSmDz2hJ0wgz7cs5tnFx+ZF+GDJdJj9oM
yGSbNyPeL06ZThNS72fHuJ39z3DaJkDb3u/ikVEmKddvtVgYT1ck6SBl4f4+6HQ5PvGcdlKqB9k+
tZYOifDkBMvwseFt2K0V8NeGKlxpKbudywOfPfhnCcXBDYxsFZuJ0KMT1evAAvc2vmDW8U6sG9jE
36lO0HHOPyq4b8O5SgdMPlMnzCSTaDMsFFMSfIZIzuAICFvNKuOa27lV6aVbnKaGYLTcRTIZbXzo
h9ULb3gS4FuU2LhPBQ1JWLZvDpJ/Dz/5yOoWWCkOwi5qNBuKbAqwDl8GdEVaC9+bREU2pqsVjTLo
nj0yphuoRA0PFLnHkxDQyKMxU3dpAFmmATQb+btRCRmAAHjl8ix8sXBjUDHzH35BpBU0waUoyTbk
YbMTN9TO04kBvDDeg3r82X6U7DBNhaHuXCVmLCIPrsrZqqPeYGoomeq/bH1QuB3O7BRviAYYSXVP
hdxIaM3Caxv5SuGLTFNpmLNhX0qOqLFi9UWbleYaUcXfJqHKAzHNGCiWxPp/FG2tsqnLd7fvcIzV
Gn6A3Kt81hf1tj8MYNzUq0LqrJFhd+texetEiN+iEIi2AfD41ZYFCnnrGxDhgbFgjt7Pgpev2hf1
TafopJ1qjnqIidQPCPvcKQuB5doc2xeA5FT38ixczjYYvbFMOXPAbVkatMu170Vl35GMf8Z+BSqu
HJzxlx+14VezgnsBmi5PABBSe2lhLp6AT/ZafgGDWfzVwTuVkb7LsHpIrgmm2wtN5NkluwJ44oMy
sAGIg0wBpw9O+oLaekaDDNCDD0B72We1s1ALCRIoZnANsaJ8O1N85qo6ZVkakbiGlOR0EncwTzHu
TdKSJJ9FzNqv8VKaaV7qa9kGkj71ThoKN0/L6fy3hdTBwKmf/i/f7ckD1CHfLMfA2kPPQ7SLBX8l
KAucHJzCmMSh10VLVUsCfVlLM7fWBWeuB4MZNgv1LQcNakC8kHgreaEimdJspfCCxTKzdo7nmaLh
dpXSSpXhhHWWWShydpkl9m+wR10O/yrC24zd5RCvwFiQRjblToF/Cebyvay3PsIpbxjGxEctQfk2
WuwB3U+kxFkSqPyHOk/Y19enL5s95Xc0DU0rKEUg7zHNTX8HDmT83ly23svmdgol2fFioE/eYIt6
96+7TJ1MAY85Iq4iwKhxYvi4SJxW7RMw0gmQNg9tFVeUQY3ikpK7X+Wk+MQLQq1bwElVo9RF6sUl
Wt3lmd8rpN1+JpJcAZ5z2GWsLQ6MmWM/5JrScjHqMQfVNRbnU+AT3flYjaB7sIV0d7WNJrrXUzcl
HiG7h37VFlsoTZ7QnmXmHD/fCNg3/Lz5hAYN+TOeCoc3j4hwDYjCnxk76SP9r4RMqxAnD3Vj77vf
df6ZpF8uIIHmIUva2Qjqe5sb7t08dtBn7KDJrJaD8MXNs/sMJOe4mt9OV66QL7mH8mukSaS18xSU
5BScUQAzCEIajIdhx3bXYjARRe/i80Atxlya447v4FZsZsVPD8Vb7sC0oy9RTUH6L6uaDKJiksPJ
kP/8V6wYEGM7gL5T3ADPiFeGPeve+SOqco5Hdrfi/ymQg1Ba820CvEhFEDckjfelGh/pPR0riaE4
LCC/ioYgW69tFWeU7zvio5WsMcOQekP9yf40Xjwcmx3helI3lWwVsaTfQmzjxocFKKERGF/uWNjW
8sllNb0ZHaqvfeIkCKBH0cO+6gQudjwkoc9tFxv/XJyLp4kin6J4NHfb6puZGMj0WexHmiQy/Vxt
vMFlPRChSbJ0yUuUHXXovF+7vBhjcI+BXkzge4WcSowfg1arFqHoyIT74ctbmT/+BW+wSVfMgnRb
1jW2foPK0lFkqTe6J9Z2XAkYWMIGpp9ckUN2Jz1mHjK7q4cUAmxD2UxuiAYB7ftnGrftqmfeWV5M
sFBkBtTyUsF1iixLr/gYa1tuntGlTqe0bCMlol59y3Jt+Rp0zM3hbq+PzUA2Tj/9Pdq78uGz6RgY
+BmPg76FkfqkNRW5yEqANlVwssjSlCaTQA+SLuu+7+RpCIh8Dmx/NZooAPuWGpkdn7SkuN6FCsjD
pPolQosp1jPpITEwOMqsA4kxQG11Lro7NdknDXfLRyx3SZNId05Es/Vc2c+kIcdLGK4yrm4WUNIS
oLBnQjpM7HsSHWkMWa4lkFwa8GiRKn+gWlkA+A4Gr2VIQ7WjObKRIGnoxTRzxWavx5LtZwn48Z43
NNCcX6e4W70NhH9+d+MR6oC/JdHKtk00KHhvWwqZCyJZ6hhxW7HMttk1Reu2/MIZHXWxXY13m/hk
cfdzTMVbE+AL9oHBt6k7LWv4cOxvW2T4eTwXNXiWKgt7tLV6jWKbitB7auYcI+t2/jYzw1XB8Cs3
j+6AsYAXVxWd+M2Npqn0Zwtstyw2LPaCdBvMTsPGp5M5WGK5K3HRm/46o4jO+7QU4O/eOnxt1xum
GVPxLZA6TQkf0smh7pkQN5yDTF08QMzafX4fPsLIzhfNVmNrtG+v7vCnzDYGFr5R46HvHVSDSMkc
nJIC7RwcSd4gcUN7k7PlNOGad4n2NzlNO5d5u2Tn2qTo3bwjZc8xww9AhnLm8FUuO7iEyJEF5Br5
JzVXPMVooEZl4XB7L5SZvLybmCxXnUu9ccFFdgKoJytDXzvO1u4Ze7nlPgss0/WXpLYvzbVv81Ks
Df6l8DmLxA/AqcVUImbUQuKebl0TVfdFzO+tPJCiWCgFF2llgwwzxvTwZb/B6pOkwXWeOoa07eyA
sOzpCUVRBIDdvePLr86rdmjPsFfBnSeac8oGeSmlU8I/nRytESptSLh05lV+BoBsjgSL2eGXaqpj
VzfKID2+5EwjH9uTcmVdn+YqxdQ3v5mVRlR4p/wz99ai3tk4kZX+Dydylrb6CksQTi1qyCtqg3Oe
G9U1dN8ogyyq0Kaj9CjdpInrOzghT/++j+4K9Lw69tFOYPrTa6D0rLYgHuV3/UHhc9n66K8FIis2
oLSkZmRS6emAQbFH2ie8K2Ypl9RgRU1fyOVuS4lZqAcygdQtCA2xeFTFJ826dkw5SbeWsmILtkwg
ryPH2wbC3ycfZEpc6z0MpYRTmHRabZhG/jfGtMlrfaAxEGaUouSHIbsjMH1a1Kkv7vVn/fJRvXH+
/R1fnfkJV2F1x6wzNIvyOn54mTrfqgb/vw9gPTz+RDAydyLDoB86SiSffbdGumglDYuCa0A1XqkT
HizOS1IymUvD0/lO+82tV5GlRc8R1oDv9AfC+2MWhWisckVHXX/XZIgwoIjixBDMib45gP3w00TM
WQ5P0ltf7S+Vi3fH0hpLl639jT4KLKuj2e185DaDXS3e9s4ndoQEcTZBq0/JTkYEk+3vWsz4tHUx
jrI0kSvXe1wxNTuJ/HYBozGheZs/wQylKVY4kffR4H8JBO1QGtjztcrBkjCJuHKyOczKmkryfSkK
oWxBkbFNnB08d5OxQfcjiugBwXmg++pvd6Tp+WXZJmL/eg+G19p4RC1phgYfd5+umxiXWKPKCaLo
6sz1j1xAfcWG1M4hJHRSRoV7sTPas4ECp+jRsIC+YKwjQhqhFiD0rL1gOPk2LWR7JBwt0Vw9dqjT
Vi4IPDjMkEzl+IMVlQUZXYEYMkwMqmbmk3U132mgb2Wn8lQawTpIb8cssXpFuuApw43TYfAqaxEm
dS/0UfDzktH5ISm76snj4p9NTEbTLvoh0iMzKZRJrSkYJTE218NS65lwkuhbysJf6D5WEFnnxk9e
M+Lyd0CjlRxDtFUQpU3FMBGBmymB5SQYma73R+2n6US/BaWV5qto5Hmy9TAiIZJxbKtlgm8LieN2
3F5R4/icB2ikUR1zWcgfBwkPc4jsEdvZKUlXwHkRtIrOZjFuwCluqsBNcpJ0S4qmreE7BhMFjh62
l6Idic1EKjF54LGrddETLZihkAuYWKeIhXUjRXGObjQHjJI5l77SIGC9U4VkR7/41iJBw3puIu7U
kYEQIfOXUJ7YowJlTiLo7Iu3ifQ9hoi3S5ImH3mxb70v+wJl7+hx6fWLDK62Ej+Fp/fUIw3tGdwL
Zw/JQXHJ0Sc3D6TMbrntwdkX9jsHl1kxpEyfI7rNvati741/P3otugOEaX7Y8ZEqmO8phmdui/XL
wA2SGN0Pm5omqgub+BEhm9ahwK+0vb6REj8sk/+w5aMH5VXhbvvKiAydXXmdOMF5LrEWWyTSzgjV
9+/vIfMOPz3T8gwFQj5k9VGlDARS241xZN0hqz4Pha38POUrR++Y+8H+SGvNWurSPiPXLTLh9QiZ
9+xSl4qB3oaTVp8Kr6xj74mTuEG0BHqM3/4UAqEK1eoNO/t37U7TOx3RjYUVdzdIzXhMHuLzJik0
8AM8mlmXMWUAkhbqWTJJZIifCSVg/zjpvWlD/DossEci5A0kEQoLjrgvOLq1bDO+QYcbPK/UrSw4
pgJGxAkz3tdjUJOeuGpL1kB8jl3z2xrKGeTJ0YNNzEuRPO4kaMKkq++hEkT7KOEmDdmkIklS64mt
5M6w4/n3koCs/zRzBUqScNonmmDU8gvaaxZaMD9fu1TWfN/mJBEBGM++m9fKCtJulGKNhO5H1hw+
oFIaWDb55Akid7Mc5kCRT+vsAd94/57cocyaAwbVXQwpXuvK0TLx8V5grV1GDorhKxQi7WKqR4AK
YFCvwPaKbEJJ7UDm5F3vFW8G4r5k3KRNTro1AcMTTnp6UVK/OuL4X29xlCj6uCqAlWf099l/A2kz
zeCot5y7eodiyWMY4Q9hgteLGLDAbsLQ4h0vPtMWgCuUZEoEdk/n+L4vJFdhQvW9AOLs8fZyZ+/6
OhKnqs55W9HYFGtYETXJnbnP5EcqYOp7/oMSrdLfS3RjjATHQbg4rnUR+g9QQEAKupfPP3YET9So
bd1xhCbcCc1hCQJTKL5PW6u/EfV25GgZ5zB/1hWoE/OpfgCE2Hw5KHAbgqld3Y+jqxiuHHJysJZx
flk77Ji4xLGlce5Llev/pnA4EMZhOrw3HkJB5uq0MDkEk8QYrEohMv4/CX4a7GnrIhFgOR0t+UCi
jw6cTT0DsICbu6OxOulZhp2glEoVl8ebTa8a5JxvxiW+qFIfE77pYlzGCq/PdzermmmaM3CLFyEC
iAY46ZUzT7YWrP+2oopAAKJOnXg0Tlk3dVF2cctmCPoEDtQswZlgPDL/FKMLPrPLCm3oAyvwrn2I
GAxninToEc+MeGDzVuqM5RaBRsaoK8Nmp9csEMJ91bA9l+uf2WoUV0IYSfJNmtiYjhv6Y5EkvyLj
I7wAMX4O1bJkHyy1pCXjZj+vOuXXbox0d5wneiLBZ2xzxnfYAPP2cmPaTuAMhW/oKpqNDTSsA+el
m8fU64C0ICmKFBNU+mGqYvEqk/xJCIUcWSm/YnQEYtWOwlhzH4c00DucO6n15+IaXwg2aZR+7iGa
EsYS4Zzn1t1mBhgWZbrf09aypkGRB9gaEdiAEDCH8uIQfwAySRv6d3x+UWG4m/LKuEDBRp5a2CvE
nnz1gSZzQ4k0iFsyFPT9uN1QhL4HUnX72+nyUt/qky04FBS/LluowikVREhLwhEYbMVB+e5Ljkeh
9YMgo6odOWUtcmdzUnGRX/eUugTpsC2U7SpUK5y08vouXONFui8KNig3Lu0vnuOI0VnI66hmzThy
pKG8xBSr1A1jV8dvxvvel/lhUOsHi/x96l5X6q49NaNR+8GQH4KBDFJUP51VE91TEhRGjRkpVWgF
oFIrdlo/+7z5GZRlYEy/tWN2dNT6m30WbdnWMSxX+uZwPFiatVXsV0yKuuHROVmr5kkuPBBbdrlI
YerBYJG8odrcGnuYoTkDE1FQWH2jCAcWklbQsuIu6wjQa92NxopdBtpvaPf5Ab+oEUIBSSV3g08l
P5vg8LdvcxBpwJapjaI6ik+alVxciqv6j17hmadwMKQQGAx9ZE3TI+9vBq5wHgpCSEeEbiI7va8K
TMdHqJ7VoTE4RoOTyYmnH5NVWm/FY+BUWVA2idXbdvUcgEcVf5A+LqO7KokFIc/vWszLoc3K5zQ/
TiWghXMJCFGEYuEvf92fItygx4PDrpWZCbGRnyW+JOFWRFVEBN5yj0ZK0RW82QGrVF6vMPHy36KM
PbVmlMSErrwe2//DJl6UkOCT2xIvTYEGL6u4GJfgH2ZvQZnQIxc0Qreh9mndpZBpzXCbOjD5mV3z
kXEX6S8SvHZtxZ0h7jWfBf1hIqYcStabZswz56nYCFQsAPrYR5l8+smydW8OCk19oG4TmXZ+M/I4
fFvJfSWDfyT4z146OQogM79qRWkFGNEHq5vZepXFkm6FlkLAmahWArgvtPvX5py6FOPXr/fpx4ep
0WrAnkEm/+cPbygDsdyxSzbCVi0Y64bbhwRRPITreC+vKYdlfqfLsu6NlJVtO9MCxMxAYHsCl6xp
CD3dVKIsCPaK8fiYh6gO/5nHXBqHXP3DbEm5lHle9rcwOgcNvjy9SIfGeUCRrNgLfgKLSjqx/x9W
crSx5LngoJI3C11UyTAWkq1fzfYHB9fzU8mY/tQhsisrI9AiiAHpY6FJz6i406TQa/wEqOnr1FF9
aZMQVSIN1KOFx1jHokxi4dJOYOmhslcDKtaEyWFVqJR1qgxNDKqbXaevpmIigoaGfUiZqNOWJENy
OT0WinwxzhfNk0wjwIeQM9v8xGWRdNJjsRZbNONrhPbwOmG8yL8TwoS/mvvx18srPelUHDuk8jou
lZ9JmriZ/MK6lt93FNn5jAXKpptl0HNocVttbAOrp7VYWqOgbJHsLKXmE6e/ftkueELFO3+yVEEd
G7eGRYfX8wkHTbdYrRaz8k0ezPZDssu7YNXYsw9b459K3OiYDy/JC6yURlErg/4m9vlqhujpTng8
xTIukwQxOW6ToxNgqIy+bL1tPbeBtm17P//EMxM4NnhM0TLz8bMXhufamGIDll5/gbitOITchKk+
lgUbb8u/uXHML11GtoanuZT1YEpxGJRgq7zp8gPRiPW/nFNXvYyJeooHIOVMgk2UYHd3jZ8uOFUV
pMZ95jYvMdRoARkgI/cM0GHHh2kAGtGNSblnh3BHnGKlqSLWrmxsfzPuAgGqgFBW8iquq4d7uYVR
/Pu7lhg5Abr7NgONDeVteSlwKVKrTb/XIVoRyf9t//1ccF8p701vmFRVE/ViTgk7VG2EvPEpVLu+
eID0DXviBdkangskF8lyMyUNJAVjgkjgEFz8Zay7sc3vixLnCcrIRQfIjZXW9wS3DBTObxSejAyL
6rBsda6+1x7ZRVGLZtGHt+wORGId67W3ghh48lKpWy7ohLQoMkefLyClS626nUC0CssI8Qk1kNny
gAS3brvH5XV3T80DK+4bj718Ql9YFrQcrKe0yJVXP9qs31dGb2vlTCuuTsILYXndh1rwBWRGOQBc
q2X1w26bjs9YQDy2PiKemwqw5tsi7vHstpwGGK1J2rKO9vNoQoy5RSuDMRPxHYiqB+MbtJLcEEkb
iGduuWHCrJ0J6iGE8lTD2mgYIl3cxmCb1xxOPAvS1Aa6uKreq86KGuobhsOtbz3ZAz9iAtj1Hqx1
ow8OAKorrnf8JYr08SB52Syt1yOT+f9Ax8BUjw4e95ilF7P+nkw7MwlUxz7oqGs9Kx6IyrhkcJ2F
QWooGWEpAD7YqPjQ+iTaeKCjZ8QBi2ww3fuubHKUPj4y17VDnAAJmIgwssMiH4fnja9K/zJuE8lG
EKuyFd3Mz1f3DrljiFqBaac0tBL5uoX+nNLpu8EPv/PXYeB3+zENxxAi4UiOb/d9QhrIfKbEnQ35
ZbUSzM8KqurFR/KYHxxhZhzM+OpC1CB7cLUwBvOt6NmMWNMwJ7xrnQYO3cPh3pBLdat/Qd3oZk6t
PVgBGCHXOZKiJEfkp/y7QJnEoe5gR88l/AHLjeMov1bpRGSMYEhP5i3gfP1CFj9+nsM40tk0L7Ag
7I41YYjqNdmnbzASElc0iF5peNQHLGK3FsR/maMSQGhjRsKMuwWWCHpbwA6hsBBFFEnacxGgakNr
PIKDfgRoIzunSoda2H5k06WJnO1MEtUG0wKBq0Zx5IHbQ/aYgZm1cZupKCNVRiBsla84jGK6Txgs
fsC0AQwWpkBh5/bj2WwDkEnT/RVT8oc/0F3rkpY/euYq0CWF+iMuRezoz0PfSrnHgBBsHsimmjX9
VJJKF5N6n7pIRK0bBIebq3K5v92+FqGmWDemclDvkvrdLCnB8rHLc3XkLFJLMUgkXmJ9yqtyy3P9
xS3oCWAks8Xf55TYXr+fgw3uE7pnI6egPY3Ejp/PlLNDCQU+MlKqLizuHB25z5+vBWerxVJaO98j
g5rWyxs0Wpl/1Q8ZNPrTbOdqKhu+JfjLERMTIwyKmCjzcKYPF7XUMYvUKo1T5VDFMawvGIT89pu/
nHp0OJn0jr3VLT3n+dH9Ksbsh96JKNM8qiSndWepH+dg8J/I+Cvd37oA1XWQQRrb4KVNBcLbIh8P
TpHplO6MASPcvlBA8cV5Je4Vj7UvJzpv5WVUWCJ3dHXMw/j3jV8Vr1Akbkyzks3Bt8tKZgzIUsfQ
1vp2oohXMRwau+5trB95cCw1HTTM7oYftyP8/DntPbm8+EJySELxWFpZ91LeriDyxGKHCMAbhYqc
1IAYvqOKqvHgaQjVuP2FW7fMawChI3CO7Rx6FId0iQ3x06w65Cw3Vnqax4msu1r3rjs0czlm57mA
9agXWSEI8ysmjsaAumrzXlQSo0bwRwCLfW2C4k2V/ZhRLwZTI5X8cpEmtBkNvzyoQWm/Hh170sNJ
n0+/E3PKlezkg/rioWmUI8MT19ekCEQog+x8MZWrTaxJ7lhbCDwaBrg1ICUZ/6aOtf2n56zMnTVv
n5KBQkgq/HSoZijgDXSspGpqwgnBz9IkRfea67ygbBfNrURQ04Z3nFCUNnNuj+gHrJ5njnvQmx3k
yj8ItoQCs0ZpyfuUvISUVUuQ+TaySRNfKM9WMobSoomNLFuPVDk1a3sm3wX4QrAC1nPEjGZ45jDz
y34BWksKBeI727/xOJF1B4CScq7EdEMwMyC50tqMeZZW/G1l6fsLQY425pWjuDCiO9L1i7vaYrdb
eNri4BSq3XCfNM9lK/8pR/WDUWQC+hjdEivUcernvSXTduCbdypwWYwr0gSAsTarSui06Nr/1rIw
ViUlJYHEsLWhi6m/I7VszA/vJaeFAxp6RUCtVxalCiExEe4l4GcNY48jm35tWAvgLYW6klfVuTo9
52+EFhpzTjKsvuz7KAZahIUewhHfznir/eYPQm658ZQbK7AoNAqHTHLWijizw1vEEDZYlGeBqCxA
Igeb7XP5E3fPUsVhoARFIALkdrpbA7V4AjRAyZ5yk7N/S7xjDn1HFXCbnXqzb8GIm7OftNIF1DJA
vUaYDozijc+NqVWgMVIqeOUT47oHp4HOK/UdftbQuQ6AvDx9VpdTrWEd2H7ONL1/XbR1pZQ/XKkl
TBR1B81Sab2ZMZkUEzxEN9RC673eo+VNQ6SuE/PZvL2F90xjvguq2jikfGnDzkRtKam+cS9sH4S+
c85cOSlZ2vZc61XxQw7g7CXnAkccuci6Vs19HXLwVuyyXqMeTD36Fqbmi6mCbIXMG5k2f18A80L1
enqRm+nq4+/EyesMP7OHvIa6+QM7p3qTcX+eBWPF65o01JdlaskP3GR/qFWWCjxKozrrisp2/74c
ajw4xn92ZAoJ0Yi6lhQdmqlq7wiKrniUuIjru7U5EByplfz1A0XfZkyVNgJfP6fycJcsAdBPWFcl
xPfD1NQRS+V5rGQVJ4OJ34Sk4ti/ALI45KP+J03JUJoCEeHpwjgS566RaGnReDp4JWq3YOPNdFuQ
zVkGpbY8i9Zum8gPnM1jkyLIrYREvFnxUJCr9/uBp5uxfcXCe2SCRbNxy6pJOfqBBnHoe6C+xKb0
vYGdsHqZKMOH4tmLCw3fDXlR1U0TXXmo88ls9jwKBnMdK7GVCT1Z2WpnRZObRhtU2HaTTvYY87ac
3r/PsGxg3qoAb25et6XSMr8cSyciLJmuqQxtT7o76thzmmfdHmprDWsxEA4X9AAVJLcITIAA8F1r
qwJcHfl0iWSNordzYLT7IOFEsfwg36I0hDbCMGqZvUQYywNyqtaMpjaCdp9ybZhCmvGiUKNLK0sY
vqufPs/9GYL4os9XRSvbMDKvPa8Mm0X8JQK+R/M7OqBTXjn537FxdGF+hVJ/6++7bTAqW1ZlUVng
vZa44forJWbLnjQ3pqR2UxIeuPzSiCQVrVv/f+MgUGfd1oNgWOfTwMJ4D7rnNg+UHHDKswUS7CXE
WVQ0Fn+oJYGG4/+jK3uuV9GONqmV564+UNPyju8wWpuF99jROJUNnk9EvNmqm/+5HAf6JdzRcd8k
1bWm+Rp2f8ppSF3gre5gBwMiGTnLO99cXiUBkgR4yphYqsJxLdwncvs3bChTwA/yMM29X3veMiBx
nyuWr7rvuSjjbxJe4vsntHPeIGdcrZTIaij9EMIIGMXrNrGHOE3GIBPzofBKGhvAhN78LRPI8RxO
cs31/JlD12WZqi07PfcPO6hBUYMCxKNS3Dmm6jhMUL21NAwAdf8T4jbVtETxJQ0cXrEUww6YUPf1
54FOLjU7L1ggDDk+1c3b13xhgtY88D8qijtHoNApgqiEQIB9VglzNVSJOvmqoXZgLDrUCf2MZy+V
CPRZ11iBGtLJqSC8MloBjD35QQCCxBK+LDc0QfS2YvgebEJDJjq32tRJxZ69l39FDkMpcB87HDw3
O3u7cNtmNuHwoq6HykTVMsSW8kK3gGIqeCXnTeecriiaXCD5SvZawdW76Skd9NlOmc7BvI6dN/dd
+a7pO3kJjgFpQVtC2n4xUJs758yOf0SD6CjC9m5i6ZfBeRABNdvhtiBdTqFaDqkTpnQFZ7p3QKYT
VK4TkXZEx+N99GVxIr0fu13qAZqWcfjZCsWDE19VqU94oA6VvjOTgko1HUfNdb9hgvcxSbqv9TvR
2+D5U6hyRHQqU//vchGplR4gpbsCCX1Bc3rebzaJw6e3VnrcK7yffi2ngS6bAhCL+HDkphMOV4hG
oPUAhibTNE7sJZqkbiVsKy5rEwt/JAAM7lX4KRaou+DUnOIJjMgildEmWpGT8DAcGhBnYmYjQ64F
qUvUsP+DxEcZ/xpAHVslK14xF0hgYUD4i7UYIN/2Yh7VztgFyFGZ9MIUvVKo6gbJvLMWZ0Gv96U2
Z4D6BsswkegA86eH7r8Rw75fZVYCl/MhOynsls+moWcnQ0CtQsFc0FCmQNOSU7ezAXt7bLUEIs5P
PbHpeCpqX+sVOMni9izVz63smDc6PBipD8HrFoSSe8tNvR02ovVZqNQGiDw5coGZkO/h/9GMJGsb
pxAhk1Ib5lUSf0LBwWR0zJMzTUOLcPf067y+5YrlLus8JqJ5kT5HpTalIq0HiCU7ms42H0j7aDSJ
ow4THtA5R3X6pQkapEnCL238ZInM+pM4iq2ikucSEKZ+RHqPoCq5nHjhWuxx4lyF3udPBfKzJR2s
csPaUTAVfmgZHeL5rOzEMyRtWLFi6zLx2AJvOrywxREawGDHjUFxXucKEqnFg3RuBzKTJk1LE8F5
GYHCfr5cWpLG7oEbs52E/QtsbG9qLk0MtuLx4cMR+1yypEh//KEIajEl95Dh65lBm9tPYIzOQb1p
csjobf3pzLVXKK7VHbhKWtD/Ot+M5D+b2Ayu+fmB5LGXlvPJhzTXLrpBFCXVGB2PwMV/KTFWGmR1
p0u80ig6Qy62aw489G/sjeYvnL9X3z3C6brcW8Qggs9vY4uDAi8fWv7ABz4n0xa7JPUsg9fuc++0
iVryFTOE9uhZL2+98dhxMO5jO4tcADfMUAiVgKBZ16q366LpsYysdJgkEYC2/G61v7zXpyP9OyJN
aOb/vMitBkvQCis1m0DTtZ+QK+yM99H7LncEj/KJaZg8eshtN3/Qzu1GYt4vTpUkrI1FskPxm7Qg
GmUIySmIOOHDT1DHdO2eAtIun45kuO/+q8B6XotngazmSOM8x6Sffk9/Nz4cWgumYs6V400rcrk1
LwIjloBvA8V6QEtxk9RnTWTYhf77A9E/WqokoOkpTKCdDtDqY+l09fzi8fkM00Kl5oe6vH4hE/Sc
IFg44cNVhZvY/vEDUXRYPhXjcslgNJyA4FIxyrPVRJW5A48L0+8xBfxHnAzHmSSd6kgiUQgzDz7d
uUab6IxJJULL97Sy/APwLqZwzJDeY1PSmQBlfTc9fGI9mfY4eDiXYSHSS1toNrJLxLBqr/hae125
CbV0p9J0lwTCijpPuKHj8WimscUTxi0HOcySIW+d6s5KAjpBXqIpPZ8rOzfq0iXX7YNzh1Y+usEM
sGKCFNhzYyzB+Oj7xIdy9EZN1WtsGO/Wy/zpR/t6AhNT2u7l4ZV3EiQeY+eiQyWfUwtONGR82W/v
tgli2/1MUT6+mF6ENwB4F5+XKKf0sTVdbAIbyJF4eARQrSnLIZZNSPs/Xcs3DQVyIMehUXx+JKyq
x90MV6NJeBXtKtBHIRrSkGZ+/dX/+z4sKf7WG6r6B9r6EBgapD+D2G24Bw5U869bkEQJQUu+nzky
ESK4ijnizuL4DoYcQvHhSpxEvYAJLhnwjMxWvllED+SstQRUSrRRxpufFATz7PbNetJsF9uRO5K6
Dh/F+zYYiz+z/An7f5FBqQvT+E/jIn2x8/2kaQstF5oETulW3v+dZ/HFU+BH1xnL8YpTB0wx2O5o
nrKVCHdPNIBwYIfrHDTCdKGJ2N/puB1Cl14ILdzGSPrfd7jzaqUWDAMUjDxxtGrnL7P0EYmZchHJ
pKfk1Un+IisL/3woZP2Yq7LQCtx8qSo0y8sZTplo+WV1l5mRngSqM3QZKDqStozoIIJBcJBmNNUm
NIHyyGNOy5vDjyd7Oq8IgcVplqNfWFNnh25mrvI2WmrZGBZyOjr6rB+ykG58gcJqKZQn5k2qn4ed
zltpw4P8BUQvQcXfgu4iWW9KsjhmanMyQ/ryZ3vThDzYa5OTl5bXEo2Urq4SAnYcm6Jpto5hjn2j
XIY2fIHcNFlSrLhgsu1pDx00nkUoaRW9B8oOpPsYbShSGHKJwf9kD7LEIKusMnWhUHiTWDmrA9Et
yrGP/ZLfa91/CI6HrXKyzwrH4II9IoeLHNFlBnOkSVeDfmW1hNzXH7uP8kX/zIZ6/wpC9N5DRD5s
2kYjBFarffav1t+5tlf1+1w9upqZBjOJ5uolLkb21+tqrF+mpJ0Qb6LlcdjuFLi4AIkweAQhGGAO
+pPQySQ9aCrhkqI51hBQLwfwrkK6lHaJNk3B8CtCxxhS+LC6Y7EEqBeJvAJCpDCAsGGb0WEGxe7e
rR66CpwhF5p+iIToK6hHl5/As2L+D02n26WRd9fkaT0RBHeU/Z+LEMRsFgZnBph+BgPU0oLTV9Sv
/wMUv172lDo1EuTALuzHmgkqb3QKP7XkqpoiBM3sia+HKmbJn4jOUEAgOO34N6RBPIFicarQbh2o
DzFAjW8lPA/psoMx0pvR1AQq/faDfyZUC92+ZeEb8400R1whEDwq3C0r91ULOSpg4M7A4qat71h6
xcYCfAndLi+PcU/ZftIbtI0yC2XSlAyuD/K1w4CmDzfm7YDGdrmM6Us4DwZez6NEO4EaSG339/fE
LiuncQa1jleSA0ns8sZnd/AStAYGCT15SAmyHiP31Ghoo33Js+s0VNue4acAhjZ6oYSQjhGntXJT
tz145UDySbcte7mGj3o8f5KwWM/+gjZMSJPJiH/1m6CyhkZmgtLpxkNlY/ubRDG6UXyCzCymoCc0
FKBP4s7lgAoTs14Wg9fu/qF7SyKBk4FCu/5uOumAtbVTB+n8Y23TMEkxB1qIpEPsollb+cIzGlor
HwrIl+Wu3DO4hoaEiUCShGlQ8daXiK/eeRix0oz6ye2tW5jP6wIUazpjw5Bz9eKOUn3qkz2LBlYF
qwHzfWZwQ5iIy9hcUsQbU593OZu1VQUuSqPcWRziTe3lKQINKpaHVfrwiVIpLZkpImR6xqlzXUy2
Z4on56PcNOzv/ZVJQngm11MJKP0sTn3tE7C0fPsmP5bgvmXY0YnpVm68lmcMgykTSDqgFID8oVZ/
oTy5hSC5Q37vVw+3DDm0uKouCnLsKf5UVxPXzGFDb/R8NK/eOe02PD/djDsyNEWkR6gxRKgeBPoP
keVcm1JEg2zqhZ42XsNxQracdFyWHaJUytCRdDZ0p0ewiH5/ZobcmNaSG/FUfZf5MCsT3Xf1Qjht
in10q859PG2mj4TnlZIJIC5O4p55N/3kv0Lsl+i3wdlqELzo2TJaaDlUdrlpms8HTSPXKmOjTpt+
UEb74NFC6YcKcBzVT3QIl4pN4QgqGR1tb4jbaXibS1BqZPfXGxkVTnCa7YFjqzMbI4DVrdaMXBT7
heal3thma/VZqPzJa/GlLHOyEuZUbCJHBP4AHeBOMKXKpUHN9BdTpl3+eDcsL59FiHpoDkbWv5YO
y4vZR85Xg/iAgpgua8gfBU7X9giO34XSG9HaOluKRak5mx88d9n0hNWoXtnJZ3ENsjQskcQW4fAP
UhvFb6Pk1N1Tk9DxC0lYlhlTjtP19rQnv+jLdYHbOhhGZSjzPVOgvK0Jk+v+McDZrsy6uW2jHJJu
0hRAhskkSLNUVsNy69ywY8STqQsyG8S6kHZb8KLztsjakOHtNWrFOSYHF6JeNWf6JJf4Cbqm4c0L
45Cphw5QwXZi53kNhu7v0v8644yWyXBJRN5hWfpDteW7bdcyYTNQR8W3NJckk56J2tEz03ibhPCo
mxNiML5IEZxfdlbTaas2kQuGR69l+PI6nEid3cwUiyxHT0MwG6FOe0Mhs3VgDk29K+kawLXMzZ7P
E9WjqIGWd43VDfhDOiiQzlBwaYm/QBnNKB7qr5aGTJsrrRal8FlASK11CZ/1nz67DrWJhuv5fL7w
K4SyRdkLkVaD0zbWIrdchereyQE/fujlT93Rq91JOyHZFx2RKpGZe5MQz4LTBNh36l13mNdZo89U
v65ylWXpXz5rf/xRB8G5Hx8F+DbU0y8P7W5wTOxb2RBTy/5G2tWi5X+AhMN/EP3rZtO4Oq87beFS
ptqAa9ESWAWYISh+EZUTRCOTsdKwNZgOf43HL9342neazQkTZo4a9HCNo1V9rHYR4+hyC8v5ZWgA
DzFgTH4P/FQe0vX/S9Q4sB/a67ncEVjGbUaveHMmCeTLETFc1Nz6x7rk+vPMrVFZTH9A+xV0yibt
BoF14Iy3XkKsucecWjItNyaEiTnY6Y615cQ/l4UmLgJ1eD3vv8Dtt2z4DwYHBxdhHqZgUv8oJfhn
AfzhUKB/DP2q9+vXB5pz333A4UzBJUnlMojz+sP4I1QTF3swskVUbL6XctRj7rngegqMo0OS3lT+
pMwqv1vOFWDuolN9hEfhw0Pt8EcIuEaVoZ0qyNb25iKa7bNhIX/Lpi0qhpte1nbT23NLf0WSojfd
1QIOZ8YphROSEwcPEkrRpKlN4YJG66S59PGJduVa/j39ZbzFNtBuz3HvzXyzlAsQNrDWwv749kga
jQlJD+mw1z+5EmIdZxQnUsafEdVewJ8lQWi2BoKQBKOBWsppEF2XgXAWCpLrZ2HyAVFU63YxhOEW
z1Dylcol8jj2Gzg3gegWaSS6Pr8jli68HvcJcR+YvPMOTWHIIZuK1w6sR2jsDcnm3kBm0Hr7Fb3z
pteP4Mr7v9kZbgb9IBpuQ2FDntdkIjzW/QBRXbt76N7yYi0MRR2jFdKmZYzuNd2DYf1ZJlBupkm4
34WQbmF7kKbO8fax3ABOqdWQr6u9lp7LEbzkob5GAEarVFV1RYlxOPdW7AXq5fRF9TUL8tJeoZW4
8hdT7m6oEXxcTxEu3A9+GM93feiQWnmd8vnVQcFbL0yGNKZAA9eMiYaGuFXTJpu8z4HeMLbe+9dl
snpL9S7Dr+xWtAgKijOesddncmzhkElSudgFBBGSn3z2xdlicYMr1vNJY+mFMFpwKdJR/kYAODwp
EIbvzcntgDXU9UENr2KJe/h1mCMuU87014YvRg/bo5DkkrQMdKarBSUZZmBcqIRI/zsjmnOXWUYh
BHig7lvOKOBwu8q8NiAa1FSIKmyRo8HBDYG7GHHeRXPpXThCPMXVITOF/phLhAsyk2L5/3x4DOrE
uzsnw0WWnoF3PimCJRyhcbphDAmJSBT7lFrKdIXaCwEgU2UV7EZ2mkMobmE4P8OAEHgE5iC6sZE+
u9bOIzzyEEbXQeZSgr2QdZxeMiDzm2OfALhz/mG19wqYwk3lKzufIOhZKVN9nwFtG2hqXm36LQKO
XrRxucS/RYHBcgGxcLFCRy7qh0Zbqqae8yJmsNNVY5zOuP/P+2PKQQvqB3RDI2x/OC5wUWDJKlEW
NrSOHngyctKwGAlNNBYobt49NLkic9c7Rarv0OsRbFdvncJ3HCek55hkTyigIxIWbs76qK51/0rJ
U+bp2UOpoAk0WXDIRYXm/4kSk6/94fcKZKt08KZvhrqExHz/E9frHvjR5egHD7YxSKvN8J5u1gXU
JE6HozYJvLSMyl6e9zx7dKM8jApywcQPFNmrot9/z+knpmJECNy/zNMqnDlCaSZgJcOG/Zr/fJ9q
tZzl7FfW8OL/0/PVDATJ9EyD0BSkkztp+/AyUCQDei6jgIXlyLanX8S61Zh29ju1+V4FEf03Kwrh
mFp09H3I4V5d1jJfq22ohxdYFUT3nUJeE0R9uBcKi8w07r7H1vPMg/DkZPzdpC2fILDlb1FQEw9w
auNRMKA1i4hKyw7mkmAdK2wADeLr6494ntXlLcJbf6mI4FcursEaecHXaHzi3eSHg9SUXIgSmGCw
UXA+Q+2nGF+ofkcYMlo4KQBuWDoJmksA9Oe8HYvVxPGw6Rcq2tola7ac751nMOW+9FfUy+qV0h5q
LZT8LSeK88mWyCGk13eh+vU2M9Ysk+g2wgWfgTu/glia+yjyIgOpTgRfdbPwr3J37u1G2EkFqd2g
6mbWyGsrqsqowpbwfH3XBlem2yuJggRhCZSO8hCTVDOXDJr7yHGFaJIv5gIlWbKzA6OxT2G1PNAx
UoqQCvvAuSLSktXRjnBgPI7wVNUiUF7BlUQfkyePr0+ambCjNmFL3Pg+JEBWG0tpaTuHoihwOUSK
Ips5zlKtix1C9/+9YXjjlB+smgJg+ds6B6NbDDTm+UWbvC7O7whgtk0xskK3rrNPu24JWysh+Qua
7Xfo2Cngy6wk5Tcl+4IF3wnKoEKvIYJbuqrcccC3WcZ8lnkuJ9TtYExdN/ly+hRymgR+zp7lLRan
K4yot8/w3u2eXZ/AS5o05qS7yCSFccVfRaN7nWPvADEBjZ95ZutrtNiJaS7Grtx8/WGNKcJDW1ev
DhvGnsHUoHogHEtw7rPKd9KhQSyK/tDkM1nlsCnvmHVnwVyfZ5s3yMc1dVFJVbNc02u0mkjJD0+J
vWCHHCSNExTxjp7clnsXpaEQVqw6jZTvLhHqXEcnRimiZsLdQ1ibL26mBjbQ3CohSTu1/JcP9hp9
G39to0Iu1QaqFsyKrIkttQrqRcDr0guDvEMtv35ldMv39GXpi/72r3WjlnhpmATk2yWmKbJFDFIS
VWpl+GhImxfKzeJRHRHyhdk7mdA2W/Nl2fSywMEmftX/03QztIouDk6cXnqAKGAxDjo5Z9Pyknb4
90GSkEGMH7iatZKT+4LQpO/Iq+unnekNCORfgGKEZT+Jyrbk9xbm9/uas6Fq9heXfu+UGoIh/Udw
qiuYxVNffBp+cYiFJFlqSX/eOYKeE8mu0UX4EWLnJPFNZs3OhbLMqymNahCQFrB6loAZX+6I6h3i
22+RvUDT8yAb1JkGLjLmuEUfrgKkSZ8VF6KNbo9mWbHL7czmxFfoqy6ozEEuwVw3ktElE3YcUHYg
83beim4pepTeAP7D4p2bc1+I1Wm/ztiLGDLvlxbFqeZHlgEu6m2wSoKrGtCUxRCxW3lYZtCSX7nQ
QzFKiM1L4VxAyw50H/z5jVpdCNPnH01h+1igCOMQ4e2gsYwuLVYCPWIqQoIRCCJDb1uO1FeQJqRY
hGHxWtYIk1quvHAX4T/AvcA9akak1SrobCtitRWojoY2IZDtJci9KfLp7zkALezRoyL3SeeWI20V
Q2aPYMQkB7SFN+kly/4R7V7+siTNnGuXrhjVnFQgIKpXhliGfLuUqpZ85kTjXrIrvHbDfuN9KL6A
Hd4jYjAXoeuRnrG5zQekNFb/6ytjzE/cvD74g6/+riLYfJHsZWuPQzFOIEJgOMGDqSsi0J4LBbx0
fw/IhkmrIsgyG0dD4dS+xTdbk3ASJdcd0Wv7v3/uw8Hq1oMUnkYbDhWy19PlZBUaK/TsQJzAfJ4N
5Zy3zbYzwFFISIIsjzwx4Gi9u6+Kp8MNKRndtxp1Sr3vwtsvm2nOXeL7ZGcT+RuZTvqoXtgrLGhz
kRsY2LTDIQagElVQy8/j0kFAy+Rr7eZIEin4l7Ze45kpHWFx52WEgOj7VY4YGrZJMzuCnRTNzMvi
cNg9yv4grOBMIW7xhzEcMGjBzpVobfUEntEnFb0wdjf2XoyoArnfUbkuoLxKVvTuNTNDZBu855iZ
fy19M4QMlrRHmFkMsQOLgzb8nV4nRigi6VUksuVKh8XJMGkjVLQsbuVcF6MnHGtbs91t/u6TGL0F
Tq9Kd5lfUTfbPPTy/omUdymdQMUjVOxKqmg+nr3ZK3+T5QrgXjTpS00j9B1AHTEyUql7g/QG+xdK
w+1nBy53xPmIbN41A9UJ8lJD6664KCBI36xgurulpzL+9FjRrhwTCnqrXZ/6lnP7ezS6wOTrW/wF
tMt4wWjBO1YG+y0LUm/DJehEUQKWDBOn35yFaaS7u85Oc254JQHmmFKYO7TZQ8FyAhu0i7MYYpGb
nfd0bezqV8neHd6Yjtinxz4EGAdtO0M2tpw9Qz+deIUnDV/UK87AzXmLV5M0y/jt+gqxTuGEZCiX
rD3Xcs8/6ZgyIA6RZ7z+E1Kfd+mU9tNiFs9LaVVMTEvKjyyNXNx9riya766PpAauhOQmlUfyU0Qb
2UvqIu7wHnEwmnGRz5MyYY/L1XFqGjlloKaQzvmx38AfroZ4FyOsyZHWtvPag/rLs2Vt9fmAa+pr
rYZCZzmoG2woqtWmoQQSXHLG+Ml4s0eZ3ysc/LAF898ix8EpblExJX4TvrZEod+kbNXN+cGQ8rFI
Ff8klkIkYg7jeFMKr6EnltoBDqDvypuzJoPk3U71721lPk0wAiw9wveDmJCKxicv7VsKuSgcu+P8
FYo+sujF7cY3soBc3r3rUB0la0N/+Rkl2f0FtwJi9c6wG9LWgzfpQ0okA6oO/Qez73WvsqsXQcCQ
kkfF1lUh9dalo6K4F1p6JYi5J13H9d1pVeTgWCHiXXLpD+uUo17I/TXD/4+mwJLnv6nvcMl5XRDK
00w7UOlJGZGcWN03jt/g1oRT77Qm1IA0KU5UM2XTthfWqsKJM0Fx/ijeT4AP13LzlZeQF+NMjzBP
0ovahaQCwjqRHo2/Bk/IYuKbNP39s2slUaqvhCEcWmgFFYUwBqMfm08Kojdbjna7wOG90gGwmpx6
1nARxW6xULxBU6lpO2JtjpO7unK/S0RQnpen588TWQv1yuhXU+V5TR3HH1dYYgkAaObFKEhWqRev
ZDis6RxN7IEhRZyoam6NCYsYUaF096hxpwoT1imAH6FWQwHUTbUMRFU2gRR2mLoazVFDghKfEBA0
OLxPVtgk79/zz8GSJo7rjGXoOiVtkaJKOr+TAa48A1OQy0JfJUB9KmnoejF3sHvz2jd8vZ9zDI3I
xCh+dK4y8rtndXqcFBpEEzmDAKMPrJUpgz8uQeL2rnpuPnh1h74xOFDYz23uQ53jbL8fUhYbc4cL
2CPchzkuMWefiXcGWGkevgjy/e8QDeGK0Y/FJ2z3ENh6
`pragma protect end_protected
