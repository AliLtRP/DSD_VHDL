// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:37:35 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
BQE0H5RfM7OZ3UfoP/Qd8lL67gaK6YBne15E2ZBF7vEZOAT5dz9Z0JpkcY8K2zdY
gbvt8s2JfpMtAsrt4G+WAeGDR0zNKGUhtLcNyqywrTz70/13WuXj7gFY/HJI8Pl0
641pbK4uNEVXAqsu/ylBH+Ddfi5NnyPl2h5Ptwkn5F8=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 4864)
mu6yQOFvMMVJ9XT6VX7BMkuFPVLDIb2QBdTwLGwoRQpGFk7Dj1Rx7pveGvgKp9bo
bMz1Eqwvgsv0OVtnGqPCKWeqfyWjQDIE5XtbEPY8w4lEuZAIXdC99x/GFoPW5B+p
743Vjt1nPznYXfnb5JoSgOpwqT/WCfkB7Ngqjwd6YuY00hWhI8BHDO8pdV2WjQdS
65yITEMedBhKCz2cJX1uDjVag9XWlTDn+ikDFGiXpDxz8GWmd/Loef8HG9FAiB5T
hE7DyLvwQeb+gQ+94yB040KgXqYtx1rE7J2lr+BJMSWweMGh9pbUXe41mvN5+NJk
lKxtbDQGx/1lDeJrhWEu1GifOaKOMBxIN37EzOH6jCD0qXHF+Bh/SdKJb515JQso
Je74tgIfp4xBA2PUj2J9bpZR3xWk9gztc9NycXa/dRDCEhGTUd8IMqZUkdT/5zDj
oBN9S6uiIB5kMcEBD6a4DAuwr4Eovi48rxjTNn7ryy+6oLrJj2rY+x/L5udQame7
LcxNruSo8hQKMSDP2qfkWiWjyhYgmq5K9J6l1pnMdICCrWHqX5MBLGKS8bjIITtg
4Pppo9OLYWiXMZz8RkwUh3EFOlKHKKZRdSO/zPNrMHIBhCP2szPM5qALga+5YL4N
COKEV/DPtPve0QesYYvR9wlCoBsJmCLfflovr1Zbkx2QGi5Y41IIjymAxjCa5DWW
H/W0HIZuWc9dsNnfmeTjMOVipRzqKbKBfDkxCTLzeifkC6PkO0PpgbBkaBoejl29
V3uCWa3v+3yZSbNnlACpgerVUW0+fT++f0eVqyrA4SMC9CE/5krJqafdN29Qu0Wn
379KE9fasmJqg8DdBJdW0+hkcPBkDky3f1GmrjF/FjwdkF8KaODwigdytOAgPb7t
T9p93Ae/HAePWbzQfp6d4HtzGM+GORo0Q84lIdCzxJIzB8DA4z3hMSt0//XBQ5r9
3GzcYqsjD3LlLZwe2kqJ26aK5CztF2bGRKuPS8b76DiTfRN6xhP5lGxIt0IBS8/+
AJQD/Ff8isFkCki6qdVLPGGCKXoGMoEd2sbF3AiVNnhyNDlLi15g6KxorBr4s7FF
gZo1hAIMt4qsYFRCKoOOUV5RU0J3RfEfShQowy+/MNwqcRNvEZvxa5Spu7I2UKXy
Kgom5XsXPBhzr0YjyAVdqEut2dJPnTKwYtSaIiaCEmzMSIuEelsc7nQQPuLXr2Wm
8xCecWgOk/r0bpKLkl0B2CWbiLwa4msOQYQNY9zZfp8tqv4eeP4Uynl1D7nHBNFS
8EikLybgxMF5zLmhGlJHakcXv81CLJ1fwPbmqkXRF/XoBmxIJfzE7hntWJ5qIIeB
1BqSVoO6Ym9fYfzHxeMOKqWZdfGD3v6hv+h9fhvTj/CGO65qA47SvmfrVfNkAsxs
QL9vujwGnCTZWMPjQjlFof9iEd1GhLUXCUWkvP7XUgz7gQLlhlmQukINatKa6QVg
Pvb2OMF7DDjqBauewITQqvP1T94t9hkbICnl9J1H6OtF4ZseH01FAiZ8QGIP6tt5
6mextuu7QlRjE2dmy4LIGtGztHfTKtoigYsxj8Pa+WQluiawYMRUCtyd30JlFe3Z
YE63m7D6RcpwFDt4H63La/eJT610u43GWlWGUFaZ8cDKY/DQ6+H8wp5gsqI8uyok
gxQrHRVB6n3neV28VrVJAdKfcBUGdfZs2QU3qFuE1ouDu1EHkPjMOgIYSmg8CUOO
gvnERKxtyyyhLx1vTyXPtV3loivbTEEiTMp+5Ey+V/yQBpoA39suakxNelE6hG4N
ehb5EUiNirPCTl/pUuHVDZKdzSEzZXLqUITyqEwshxwzNdd86CrM7E3b/VnC5LRm
NAhdTeixMVuFM6s42x2sAYhPzXWekP3kz4nT9y3pt6EkoxU8Q1nY9SHLUkOL984Z
crElmVWkBZ5zETPyKv+C1oeVlQPDmxyYbIrMODMDwh5stTZZb6wzx2eQZN3AFMhR
QTutf5x2Q22Fqx4k4Z82GLwJU8XfJhnQs5Mw6sBaKzfj8J8VP8ES3NfRv/ys64up
oZ/4I1Qr57aLgIKy9JYhZzXGZyE+Wlo6bMC58Y0OIOoG9sMZyRRRl312zRyqFqxU
tndwFtp6v8t7POF1boo0alg0vuDlMqQMfbUeazHE7cbY5lo1SStHkMfNbWNVp/bn
T/dAS0/vNu+WOQgMZItV2ZvTBZJPBjts9TvpWuan6DfyRtGQVmZViKyDGMiD9cN1
945NomkaqGOwZZ3kXcGmHuGfVQ/1MIWQkZ/n/tfMtizkvsrpGb76PRRWg6Ff4G/w
Vr8/2eBKy9kguVbBK/uufv6QhpsLjN6YQTcZ5SqkfUfAr7MpXxmJu6FE2siI7w3i
aKtJYTobloRrAak96rULd3xInDmzmsKCehVpZcZXHcmkg5KKWnd/1C1SdqH9SDvl
3/LVEuUNI1Ra5o2DAKvgL7cirYnjEqdnpB+L12AFHtMysbIb+VlSplmd5mb2tqXd
jMds8NPDIspQJHfve2TjKK2Zk2PIuJHWPR0+0Bq4u7YKOSJCcDQWymNabeCZpusY
NohVD3ARY5ENpj/g058XZezz/GWt/zWMZPhPJ89s10F0EKwm/svNHcYJ+xum3wEW
1ZWM6dPi3YA08kDQHEoVGYE1gMda741O7H+7iTmwfz6HzWmEMHdkhne9zu7n4eB0
dX0kNW7bHTmkQW1dHKYwsCmSNlj0gTFONS1GGDDnX8bqaGAxKmrXJdVXvf4bvwlc
Zh8vENLN6v3ukGd4W2/tE3Jm4TFJlTVa5P1Wk+dE+ueBpgUsyaYoNwOISNPzhLqD
1sj4+wDgLubGZmN3Rn8GRlmEjruOK15YeORehD+dOqvs2gtQkqRlKeuXIdMLPKpQ
xSnvkYOjRLFY3Qk7lZbxLM5QmA+jyiDb/32Yaj1ExkI6U3u6UMadjRZEExFRn0Mn
9qpzW4s49+em1rnx6zkijruY9omgp0rZ9aw9Q8WlM6xQLTm6urQWZBd17soGlx1V
sAnigIWcZXCkvkyfjYsSQrf8O3bET9YETt688Wf5Gh8oWlculIXqvXTL8iJdVVjq
KFgPG/MO2ilM2whPZV7uafTJKDrAqilciDzJBFIkb56qGVLX/Tz9zdOtvdwCfx0p
eaRUz+AXGytbuIr658gLT0A3FF9x19o0p4SF6pDNT6qVDLrYyYYgdKDxvbYYl/0h
ep6C4Amnsrle3B0wDmK2hyYkgBokQrjW+WxYClUqT/SLc+UQ1Iut3NCwgduOu3tu
fFgGNt/Z0UlbhP9apmIT9IpiPBnSweIwQQrQse9Lh2Jy6FXJtaBBBfWS1rzwnqJP
u9Rpn9ELIgyEg6Dp1/65ddYcfn0YKIFEgsWeM5Z0KnFZHFjQ8DJCxcCrdfNzq2cS
Fz0O/FUG3OZ9xdtybyMgFo6X8/cZJ3YE2bXeJ66Jsj3CL9Fpmgt1FHZkhiZpzZcF
liQDOOXYCqbWTy+rlH9KtxlM+KhUUQnyezQfMbDpALV04EyPsqd5hcyfwhocmHsZ
sYFNskoK9BFxxouspxAhb+w1iCKq5hUdW4g56GkVNejPvaZBuf4oD1mN2N+y01q5
OivImXuMyJ5+l/R7jwdsN9+awh2X0WUKsjMjmczenzCEIgkQJUTpwOByBKxHOVpA
wWlXTGzzlFpB7IFDzAvm2GAk0m+S69ba/UX327oaCX5wVhNoUk7o8+Yw1uDmS9L+
BuskSZNR8GwhX3nL2Naf3RyNLJliksejTwVrYNQquLsU0EPM5ECsoP/xWre64VN3
f8HAqSj/nf4LTJHhVdeifHDika5aEn+4GlUNnGAYJRgf8txn13QaX8YZ2PE5vGPF
aUQZgfshleVq0nBM6nL02CIBLI95sRQlz6+fKGtLZR4u3bm9Xg7AaaLeaL7l/KrA
nh3UAdyscckaGcyWXnlQfiu21P5vQ/GlLP5zP3TBFE8SxgPwdC7vt0tR4ImU9OrU
WCMIePkUhATEyhtlRoopriAgUNj3Qe1be0FkqApFmSLrf3bLH344SbCVYIt6kqWt
3Hclvek/sKzVEwFIZlaGP1PR4fSxnW5VNZDuhYDaKdiX2AqVyURR2gdWmZ857clN
cUA9Zz/Zf9Rh78+IQ+LNOAPr6A0sJFTrgydRZ9A9D4cW/LzJD5a3K/4Qg1Fod5HZ
zoDF8zuIj281CIm3aHJLc168xx3vMS5Z73mTKxSlmaaboToy9V5vlkIJdLGMExCC
X3U7svbsB9qrUCUcIViOx1iAcb/jZqx99aQix1koub/kWi7CYnelCIFJ9tbfV6rB
gPENM2dRkzmeJ8Mq072xQ7vin9crAed8ETAKBVF7eLjyd9FTpSuyjtujWoGxRB8U
YzXlR9ZlQfcUb/iFC/h7heNzGbYlIpq7Z/U4j/eMeGESsws/r9qWDkXxNsOx5+iW
DaymcwgXW4nQXRlfZdFF7BPynxGyCAC32e/Zni+3SlmzUlKhEqZY6du5efGO6sI9
RlJg2GhvwHb1vGM95dLk/gXiQOJUUsj3Bmv0fzxD0LAL1dt5uM2/YBNIA/0Dm1pU
UhCcjPPD/lkOs15YQ5TYNzxNEHwXSXZLMWoAMEe9Kw9OFCPdAPjAimMx0G8YqS9g
Sy7IwbRfiDfVPN2EpsO8kF7XoL/GAAmAfn1u7uMgOCArOWedTnobt/6+75aSqEOT
5IsFogqY63UMqEEASgHXsH0WU/HZEvfp5uqPh3qd9URVm/cLzBMgo6BwRE3STx7Y
K+H5uJ9w4kL1aA2nD0zuHbInFI8lh5bhXHtKN/aAGw4LcnUp8bq53yPNEZnh+vYe
x+goWXtZ3/cJ5/+fnAQPkCRJ8uH5jjzPx7aiVNqbluwp6uLGFiM2/pBoesDoLNtm
d7iwTFDvEH586ekrZ0e+E5yaUlYVK9k39ocJoDc0awim7mxtRVeERL5KlZEhCvCV
L41HPv/gVkSCiPgk5IonB4v4QA6K9ra+H4Pp2oNqkU2AYmOaT5nwcseVYLB5EDMu
nYYeeNvDsxLA4Q9GetlWRJPjp+txat3+GrG4W8zd7WvidyWkj9+Q78S+Cqg5vUlJ
/SYnSVlxQR/aU2RPx8zDSOClKAGkuZ5DtN4d6fBFNygJYXg4/gMNbJtMl52a+mgi
CgwINhmXJFRIKsYtVp1eO625S6opBszEE5T9JkF8Am1YVEPsO9zNZrJEg5LpaQUW
kkrdJfK+J7zyBCtAii1zhn58yknQwko30yiptGH/95rawvxdXyToRNch5yy0blSr
UHWDZvUGaZqoWZC3Ti+o2Tk/s6F9HiSyqdxt4KGW3lA0u/Ed15yKc6ld99V49qxp
shV4F/hMXaMhG/XlzIdaWlalEDvxsrFHrc1899BscbPFIOm+1B/Rkp4dA6WRl6Pb
6YoUpcDmhWgcrfYPN0DlOve1zXB2a4Ae5/jGOuWckohEmZlp0ayIJO/t1RdTCtSS
kIh7RRtcwdZwssE8+Brxrr6pWQVzdgdez5pcvuGU9+pFf8iT45a0xgd9g9NMO//j
aOpGRR7EujNqWBsq15/90eyYy37hbS6eOsViM4aAgn0/emuW2gTKSSLrkJkVcOzi
TmFko2pgVv2eGsYiDxDHQ6VYpgG39oZeRrQBq8wD/8b7XuhYeu3hAKQUr128yvnP
bg48dUnuR6tDwqpIOWfMJpyDXCzw42sKHZHElGAVfOgXFoFoFjJJ0vHUDBWYqBnM
PwsQ678885JiJgCCVUHjvkrEFISAJKiqtslWzaVkwUfR6y7YX5HcEM2r0TIgHicz
zEvpDPAqNKiB0eTTsfJ9r/RCaOflNgORclEOjAUoah97UYfE0k2WP8F74+pWRV+O
OTFDtFFUVufzbI5tJzlkQiad5yQ0SsZcb0zH/vJPEMJgfmUGVX8ixtgQekE14W6p
uP6pKUiONdN9ivbotFMNQsBTMbkxDdLb0sEeDpTXT5IJp6pSOssEVmXOVWZM6KJq
30ps8BH/9LBuH+nfDejZ8Eyv7iKjsNpJ/FHLFgQ0HRpBLAJp1DLyMsGHTkFqsbr0
b40UPRNdwypTmU7i/faWCxPdHWJ9oN/tbvXtl3ycCOBEztJxlmVnpAKkRuyqKwB6
L4luuOPXV3MDfX5K6R/kEdq10S84hYtIZUPGzM2I6g6E6sj7AYIsdmhQU+KnqfmH
p+rCEbKFY8G4Jd+m+GcagZTn0TsuKvdcNIfRHVPp+OCYMnb/IGNIvbMFrrV/LG+q
a5kIXajbSgBYYsauFansbW4KcTE6qWPNxLU0HB+MqcK21dFzSUPGGjDeeAtG7a1D
WUtinqdckdFYcgacpfBKHzBh8B2FD/xYKxcU/wJSvRqzjna8Aql9JkE7yyzcKNz2
89Sh3a11mSQoOeL4OkoNPNKipOIjMyG7Ooygz3gDcrlYx5QhPgxrw5CgzbhWNkZ5
ao2An2x2ntBEy79lWKxQu35jBinnJ7W5ZhLndb61e1ed7h4fr91fk1Pa/+YZ/fO/
HMAGddeVlnMw+qXXbjihPA==
`pragma protect end_protected
