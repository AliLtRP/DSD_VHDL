// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:35:40 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
dZpv96DhaQNy3vLCqCvRRXoF7KqYJ02nadWyoKW5rgbJ4pElOHZD2Iqj7O+KD4uF
Yq/yXMRChrGLSKLq7EJx7BOtyKOqnsRmICHRADAQ2sE+k3R8mE1NczqbUjhYjCwG
ekAtdAFeajuZRtOPj5WdAJ5QGX44JDj0yLdaxtg42y8=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 7280)
kuMHno1/4LCEDss0ev3LfDRD5lNlGgntTNrku4JRf0Yd+AwG8vSBN5ntrhW8n8ko
y3unyhuZwa67d07YfGhDEH8MR7jPIY7wLmCwd/ShqoBGr2CuGyGmLNPeDr7qglXj
01Elmkxe7S+MYsbRB6+VQTJBNCeUwh1TzbdT9j24JxIP6lmWF/4X0ad1Ht+wpnz6
K/rW9MSBe7zO69eYomv2AhDoAyY4/zsJIhKJx/NL1Ejy2h1JOY+PfpwS9GWD0oGc
x2i4H64duB+U+IeZs9Ofe3qyCzDGd5JrI71tZpcr2dw5d/emid9v+R/egNgTljAI
TBkOXEsHYw6xh34Naax6VOMpGVKh1i+Juqz+FNr1znoyqAOlVT22ymcR5hqjsVtt
VFfEvE0c5GhKzMTGYwDCJz+IcqOMyyHIQibUdIp1Kwg6uXW7ZZBhM7h7niSlYBdX
dgZ0mQMmjSXY1gOGgjSoElEwOb1LzveLi4a/Y7wkZSP6wHUtztZzceuTZfmqNNcC
2c9JrIKAJyUhQO9mT0mdUblH2iyiA4wuOcQ9+gb+ix8RYi3sf9RtPamK4prgz9CP
l3Np+1cVBfGWK1fAI2mEAcU1Tq1DtgNoLZzPZaKAllVUrQPNF4ru/clGtmf5QwXn
DD7j90I2jl27jfo0M/Qh3OLyLwSqlJKiIH5ou6bQTegihW9aF/8k4GUbaOnGtYa+
lJxnkd2prXTBY/w1VP5dE8qtVn6gB/CldEi6dxWXW6sHfEdGXIF/3EzUUAkNKlKU
rGrWUFGva4eFpMAhi2hvPH7bfswz5nnWEYQMKCWEqCNPiidJ0rHlOyYNilNUDGWO
mfwB+Ng1MluKObtnriUNh3c/OYtQO3lu6w5g1zl+1+ckQ4rsAraq0RQx5WLtVlx1
Rc4YCjtfjkTE4S5E7F6+DHMfK3kBNlR3qk5RJww0Xa2OikdOQDpMkk+LCGgrYq1M
PwzWdLCbLAq14MlVL/yrU+E2M7kFy5YC/JfQmYUUB/Ger/toTXPk2/DjexSLsl4W
yAFGgy6RkiW5jQhxFAMqNWi4ZZ8BYNYJf5oirbPdompc6vYE25OvEjg2CryVo2kP
Nt0ggi+hssPjd5I3JjEbdMgiJCFj/+LquRXJ/2u/CuZ9ej/j+DqDHEYhV1LHZbwN
61GaVyhCvx/VvVbAlm5JzJeT1df9h3zEabYrqgiHEFHKADdQ/oIwB8CxVFyZ3Mxh
JX8KeoakFxHNvwKdJm3WniFciaeHZA/ggRPsu7rsoYUb4AOUPm9iPV7qBSeu7+SI
7uGGHPooR/bSU4z22hxizwd+0z11SB7fJmRSGdIP00TPEpqWga+ZWhQQO/azszor
5lz8wAET0M0rd3H0uSSSEHbWkT9PjfrbEXqWaoMVKAm9sYKL8R1c1ihLluGuUbl/
QwiPTBfhfb2jPS9UYSBy/frWV3APvv+IRG9p8TQmKMJvCHpvUxPkAd9aq2B2QS6f
CJamWBlm7F7u3njUZ2cXUgsIjjaLOh+yE/LSyBPK+3Zvbxr925eGTvEQiFIa93gW
NgjKE+cwMIpUkJiultIh5RQ8HN7i51kuosr6uVxJIMX+kg6Smb1JNeapGtRDCTyx
22mMFnO1o1nOkeFMU7G5DelL9ubvYZi8I4jLZNQF6DURsMt450qLpKs75gnT/plN
NWhlneJs/mWzYJeoj79Qkvhj69ngz0ioFgfSePiwi5UDcjQQRZ/2wMlqFQpIVdRp
kmt8pUMsWD1V10CbYwAHIh3GKHdBr38Vs1s4d3FzYO2RvlYVAXHJQZ0RrFjqQQBU
7fZBf31myjeY0uKU/3fZnxjfsQyeXZdlo5C2NpxSiAR8brdCKk8RfGsaYXwfF85N
KVm8nuSziIjs/Qh12rnRu5dUVVaAMmPra0e2jJgljoMXU++nCgOgMGzbXNKUQS+G
Epx1cYg0TuYbIApkhyVaYBtYDOoTJvbsvDvd2f8KBuJXMj7tcXQM+rEghOpqp+lD
GPoc29fitJ24pX8TYYycqwumKgXxj3vLx1VqNsfP965UyIfD1ZBITpoMqECOnH82
s8gJ9iJ9bRQHCERwgqFqUh6SrksFyPJ+Tg+gjEhg+jLgwEQm7MndhLZ0YWYIweXZ
FARS9/e0hth8lk/R4WRdu3kVnM2WgL/XIWwLE9Y3gXjjpN1HNpecgWiwyy1yYYwC
DY077WPwmY+nRtRuCDVtoeKD8zPkeofy2vu+1xcWTs2DXZBeeXFtZnONiegzlpu2
Zx5WIYPkfCMlEfYJDE0cj7oeZ7YxXwB4vFy/uLb7CuH6vFLBa3PJzxKgzFk4zS18
QaGs2Ekof5hxOH/j0URU0KtjNSeWy3bzM0+gW11Ttn5QoOXMDgJNWLhwYvjoX0tl
Lzi9sD9679ifbCbkAu2V91uaY4RazRqOdHYgVwnQ/fPev058IezXzJk0vILM3Z0z
fMHNs6WOGVUcwB6HqgQd8CxBnHtkErYbztP6HOTen/O7WyE2Yv8TLJqW6F3Q8GNd
y38vA4BTiihEs7Qb7xlkWchSWGboINo0jy48y6NF8NxN0TUPW12FUnuWCMXyl/2L
l1vL4MsOCMp2ItAq3xSShzViXR6MCRBqXkCVt2nQ877UKl+85zFTSqBin0sryLzV
P61bZjveAb7brI7nycCyKW1ixxi6jDo4HMcLJWS7KnaAbegv959ooM4VZQnMKT7O
O8mvnouPiRLhagpOxwtH/lQ1BRzAn/KhVgdIcWaHVzzEFqpkTajEBZC3F1uxtUAD
6V1ZpEtz2Ze5quYr86GaIpjMfkr5QuNzVHfpfP8mw6xQJ7mQVW9kYFK3Fax7gKbE
GT0svC0RX+jJJHukY7kR2maR6UTSZQga56/r2iQw2XfbPbc8aL0YMhDy/V+ePJc3
F8PVePeemktYVxPAv37Dt7rNBn8nmjck3ze8MvpFKevRD6+QdpQWWlIWIG0jNr25
Gx6YJzMVpzx2x5XhLyWaeKjpy7Snx2WToWeTA6+o/H/SqkQb1ptQAPXspU+Gy63C
hPSd5Iu8WbWdRp3ONbvaZZ9ppZCdMKqEg4l5hAUPxtHGyJVQAHYRMjjiqSaHedl8
g14H+Uf4l5qPTCsC3NQIkyjPd7SqDcf16vUgfgRelvLQIVOmbNlK7qAMZDFwD7Xb
fhZufhQVV4i4DysN5k1UgsJzsQAu6tK4u0B21zg4I91FL8K5c6yokMNk6jw0dYTN
6DswPsS8GmoAw6PFODCb6xm72PdnWg5610kOqLniAHxBU60BSDQ0ggIjVgnvdBor
rJK9XZK/OeC2bleG9GFJHkw2GhDGK69IX6Eg+q+Vb4Gh6mY5kR+fHsASsCrK6aZF
AVTAUgKtdkbH3gTwNmoJkN7ws5PuK2PCuGgvZ+CTIwTINuoKdgH721Fosrlf32+J
356yqGjb4K7BDgie6JxbZ3+QfYSD3pP6UdBzSTOXGBWFVBe+1PHR3eLimP8SrGkl
0TTuWIp9GME1zCCIiSQ0jaxFmKJAaNW0T4piV2vGzMoJ/ZfJvX9d9Pm6/1Q31rdb
URokTe/yLas+MY0F5ojVDpnW5GvdhlCnNbpduMk5ODK6OO4X3GoFMTJF5Ei4uS/W
SW29iu3swBUU3hDY1JgGNoP3ue0G1r3QYB5ZOVEKatXhKf6bjjKZVQORw02IHXkf
c5IwM4250/HCf1IgKwf+oLunB6UNRGUofKCrJuGN0jwIQAqoVyZNwQTppSnsQsR3
7lWCdXnCLi40xPAqKGB+KqupI7nrJcQrDsKaYH/vfinipsOIhPB01bDGUQKOlfJa
+wiOg5Q7AQC1IDHvV+WkRgc6wWzYJqD05eGXY2DxalQi/G+68H60vrWOWH1328Hn
+rect2TzGgaJXDZ3b77lO5NormOEFI9aJpeCvr44Zc+fjeSqVGgWA5qz6/2TCQGm
H6h2AZaTVtzGijTAJ+hRFdQAouiq0gmJUzYu9ECptRVcCwKnhdBUSeFexvKzQHB1
jfTyyzncrxZ5NrhW+s2qWIXU4yiMFkIC/NXM1sunqoLC0Zh0Ycpd/M1ueEAf8Ot2
Yx36xORdfIvmapK6OOXdIN/Gmt4AgX9yAKRKE11L0V7JiRpCsl68zlXoQt195s8o
kQMkz1mqpjW5HYu9hCaLRlYXAYcpQvdl/snSrNWMCgOK1q+JdEHiLi/pWaliOkoN
P8hByGTbNnoTxsfF+kC/Bxidfqoi9m/A39jazHdBt8NZXllTBR9fZkF2X48tQ+Gt
dDI1/M5y7S48gim3KKBqZHuZ79+G/OV6h1NIyloDtkLo8d9d7UK1ARgihAdomARK
JZxZpzppRjek+8Mx7ekJNbfutmD2mnxSU6ULsuhDiFdabNG26ZJzbLDs5d/A3gme
GbrAvhLFCpMsYDpzxN/CtbgHffcs1xhW3xP06rWNgrjsXGhFlPFwpohY6Zp04uSt
F79ioWhQe0wWd4ekEXzcRgFsz7xLqna7rlrkVbc/5Ae9PT205hUPtsPVGSHEHvLu
pxyFGlYatU6UaAxGbKDeH39iFsQjRBOzwjqR1f5JKvRT+fU49rqyA/nCVBCn99q+
qaHykNKfLASEI3mfDIAQzSEfOSsl8IA2I0Scnw4z5JUz7qmuOzfImI7VcjhWiZmG
4KbU+3HHadrejmvdZFkxYfu3KOnWmxM1aTq6slIjfTat4iBhYPWMYrbkI4eJM/nl
VMtGS3Pj9kyz81kFk9M+mMqBkbThXSIhl4D619Mh5pyVdfHA/pOk3LuiPOvg9gDg
HQcF0Lut6cObnr5YBvJe/jHDtP26d36HvGwj5t/DA+4kFWX1tsIy/B92ySimSN9j
cv3LLiVjrOU/QehyfUTgyCmh0c4QkNsmf+NB+olec3etH6VgEzjbrlOANuHcxD67
dPRvHPILX4cdWJ42SVPU8b/EUQuOgPUfpjwD5G/wC+KOHzTY57sNRJaPZ1ff60UO
NCKWGAbD+vA5HwuxvAj2AIChtJLC6R1VGAq8jAgA8Mkhaxhxk+YRfPd/h08ocywJ
AWwC/myHAQYQB8rl6O81kT9svYFkhXCTP8z3Wzbo8lAG13w7DTIL/TpzKgeAE/Bq
FonU+Vv/Y+yYJA6fhtOV7gAoaV8VPH25GhV+2q2GePqaNn18ZGhhrgs0FqFgw3ml
jlF6qPl6c2wL9zKan1ZOzZlgXSOzcVRwwhNUd/mv2tAyfDNmN/i4sdm60rRQ8R13
u36xGIGfVjTZFinYRUrE2cjC9winIDtR/HC/0qe4xHgMrvqx3mJtjDC8LLM+HcSz
fVajihu7A3NF+YFA5P/wyPXTVIHgCwzdzUwIZ5jKIyYpsdVUEcAqqawDn9fMXmn5
kX6OU5E+gn1Egtb4IRw3M9fZSH551xtPB4Vm1FSPxc603WevpowCq0vzgs/51UY0
7LJ1Hx+Ngrc9supDKJ8pP/9IuHLAiRm91R9DFw+YqKvUpQo4St9sMQ/IHrbdM3dq
6LaDLMAvjxVEP5zbRLi6hhWeainfGWNHwQ7NVkLSiP6pyHftzR/2dxQg6N+lfp0g
gHozT7V92QCVGQNZFNIfWQuSeL11C0g75pbD9idvkwfQ8aaACljBZM9GUEGMYEmI
eq++jSo/i4AI8tV6rO8z1xQjn5xvtAfeASGVC/omEFNYgr/XM+si5vlbQm9ecFN0
h5QbXGC86dIxXlGO7+cPllxF/hL7raUcbRs2y4OskrSUlJUQ5CoNQ7yWcTzsstf2
bld0RxtxKKhBjci/RSq6P+4u9pyVc6fJNqTGk/YGBTZ76jIxO7LvB3/ZXKxB6+io
JQYsAUB3R1DXa0Epgz7T3J/xcrbpn2PZ5p+KhJlVL2K84q0iUELUUCN2X4mcHaVs
/K9JZEj5ZXsDUbn8CxlG21wItDJtgI0bKJ8bEPOppZAXWR64wCNK5M2TIIvp8PR2
osgQDCNXy4ux77t0469554iwieiSzXofvAiqeQ3pGLq3JVAq+8WsOX5S+gpDtcgl
QggxwFbjB3/EK7W+w34s84wQQel/li8s9wK+UFQKXfRhMPA32HNlS6On4v0Iah8J
ZzUtsOjEvOUEEpFprmZ1qFRoFQZEeeda1EpBhDM25QHYcLvP/Kvg51hNlDvKgxOa
Q3VJ5v4d+jniF4jl4884V5lYcWVMudseCAlHu23wBS03rA45ruX3E9YLwXfnTRJY
KLyoyHKlIlvLdNi3ApcrCWcrmboxWFHKIgK+ytj2xg7uNjoJuCBGGatjzaDMjaXX
8FRr29d7O3LCvXhEsJ8791xZEAa9hVGgPTW3IIyZh4JieK5KjJVrmwacNY+QZrkK
RVC/MWytiKJQWjm6jLGZ5p+asg5yQcS3pffNN0rIk8jKbzDp0X7/oKaZVApsXrp3
hFbg6zf4a1lajm4ihq6GIgfYVQQu+qYggs6pP8rG2+DlBTBrwTKWybXJdA7BjIeI
jiWfzmXd1EvvEi0cvjCQ/vIVFNaTbDo3MHihQAAl8pbhWs0D5Pq+4wFi+rozn6Xc
yLsMoBEzW8qJVbd+yGX/kheI0TbRz1JF1WXm1a893LZtxYQnGLosFkKsUCgKuEF8
lDelXFxsxYWhFyZyFCN+hGYHDXbakhRSvMatVRJp8uuV81ZXzaGjTbkg293+8ktv
47PgZp7R0yIztwgXi+02yguhw21zWjPmJH2f7mULW/G4eTCpK478RDzd99+gpOrK
dXDK3VBWI5RuKAFVOJwpRmpVIkTkWkoBZuHK3NTSEeYzr8aGCMXUbO4An7VxNW97
VolPoo6CrfZS+cWS21YeAvGgECaL1ZqiXfKpaZJ8ChSUKG3YuZkmue1wXV/a6zzZ
cgP0WAU49Tb04ZTjnOnBcRHKb3smSPZk06Z5QLx4n4s9YWStXNRJZD55Pl6AdwIA
seeZNbI3mzFokDS88LzueKZ9ncoh+fE4UgrzVgz51WGAYPtO0JMur9NyLmMmQVhu
7U8/jsWJ/zfkVRUi/gwdHKR4Q9lb/zhq6Fe+7pswUvyWfgZOsHGOwIy7SDMqppHY
ryWyogndK5YmXq44SKOgqGwVtW4n1qr1vVbqJ4sIPSNiDS0G3r0Q1jw3nac09oDw
7F/zGgbo2avH3h+ET105oop1gNSqkj58fTMUATP7bVUEUA6aE37vDLbfj7QZPN+H
67h2JS9pr3w58cnubJMTdzchX6e0FABKW9uwm6jaSIVsivmKhu/JikzOs2TIRBoL
GE2hTXULPRcRgWw3e8+N6EjZJQiiOSaLhITd5Bd1hDd6n3OdMIzzSAlX0krkJkHG
ptXNlmJVLDRp84Iv1TP+wGc0deSEqwOQQR3MJRHb8LV//HivEyJKU3hK68Wez84k
zNQGbMKYYUL5aWsICgRSO6ncnFt7XWN+tVGAjuV0gSec5uwG0vWO+mRqBQWLKS6i
MAtWANWm1f3zfjaKn+8ethOgsy2URolycE3V1TdAPvgB99h9b5vRfznlgdZNgAwG
bI4fAmSC8tUeLJ938jpoHbifuCzYLtVoVxxhQGdN6bgbNAlrPKVRT+2ngd54w/+O
lOH7oEh27iEtDizhHsnIH0oa9S7SWpEpwoljbIDEiTTgpsZAxda0vmb1xVRWQQJj
nChoJEqWi0q5WG2IKwKJbT1YyI5J6pPTFawD+jQ0KZVO837JdfCsKZYn7OjqkY+D
h/Vdujh7Su4EhYs9ItEJNCpB4DOPPbc9C862j2ASnCWI8A7oZqHyk5qsSTZJVxRu
sRjZdi9YZ2zZJ7g1HZqWBE3S0C+Oc11z+B/LArXBNX5bEdcefGxjs7A8yArWdZQX
4lk2VIWktVwU55MPUmA+i8LGkLwod1bsiu4WX1D/GYbsDlM08s/FDWyR7pa2BY2U
lE+VZXGYwi3yIsQIbwwzwx42dih2x+KHuSj2Rkv2wzcAFctM37cE8qTG9OYnsxPc
RIXg7utYmFFCnaC8/2B/2tkwh8+VfKXiJ5O4G4ymn9BrA557qGQPPrhYQcOFznlu
jrHrXx3opo5+WW7rOuDPLG8hr5LaO6Ij0cv9JT8Ch7t2Zg7m4cH1VeXdVT7mCoqf
Nr16PGOerc6fwd2i4oWuiUBM2LuLCQhyZH4wEtFyNe/wadWb4jGwfw2A1Bcazg1H
eEJvdJE5B9VHhTqRywuh/CFfYpvWZXyPRxVK9MK36EzVzhmDqXLBM+dfa294AxYp
WJhV9QDr5k13JhbbrOx+l7flDPHGN/R73yu0V7ZQcyKw5f1fVMhyfwIvklEBD54E
iO1DcJ3VYqVEit3ltSUGQzambDlUab8RHTVJ/JZiRpmbkIhwh88YOCnZsiCadwLC
kuZPJCh1F3AhV3T2yQDcI5vcZwZjBWz/xwJpXjbB6kMxJCtm2cOlR5SwpBLQJvJK
XBteTpKhkV84yIWctfGgRsiVgFU48LJYiVl1EYUAe8LukG5ED2lzqlMbu9dgU2Q3
H6BPlsi71oGRfZ/PabHaJjcpYWxcSeC+ngzm7zCw6m6T7O3ulb7X6+YaZIUT4h9s
DbAZyxhz9kN2doOjZJa48iIYUNWhOMWRoOn1JspEjBHh1PCO/dQP1tWt9eTPUOmc
xCYryedVcVUVMIqRrDlE+95qihdI2zS9wARHgWAEA3WENQq7grhua4AkA0QVX5I5
FQ6WhPWr5UzZNh1ifZqFNN3BE92UvRo86Eqls3sStSxBIURxHDuMx4asMug7c3DQ
AoNAmrprdLEHj1HSRiW7cqu6NBHDIDzDvYaY+PyE3QNKaWMkQWfyYisWvdP1xKUm
OLClDZo3guJKxonjRdG3a7uGVWyzScP66bb0FWW32BEjFfkZ3R8K6odW6FDcXYmT
ZoV5Q1kljD7y3nyBJE7aHRH7HpyP5rBCCSDIyFW/x8HXZtwFjanK6lIk7TP1GFKr
J24cjxBUFi58hiytMpb7ks3MWSa9hydTJlZcTzpBp1uA3H4k6xeYe1jG/y2UkyBj
LCkSyhRk5ck1TCAvqezqUbRT26NaJZu2mP7kApBZxTmuKuXufIDsMd/oNScYYfSp
llR+/H1kQw1LzWTxx4MjZd1fht+Xn149GpsND8vADTHBqWMKFeAdixX+GP9O2+ey
e/v3OoGZMrdGClHhz5eFDt+TLGj5BWoBrZ2I/aBHzCELnX7tfEXsdVX2kUCrvgU8
VcsV20Ih3o2r4h2SYcrez/MrOTqh2D9iVCWeaWrd7MZAJChhp77cAxdslAMcDSUz
QFL+q5DekEoGalle4sEJHyAtlWCxH/TSuyONSV/3SB5skEpU+sXbs4MFBhoo6WUt
98VfO8UL4+IzK1gDf0+J5j7UP5cG2oJG3Qs7xc6y7IkUbMRD9+nQzxRW9dOmVNRh
k5sQp/AMAasQ2tz/zQpa2ijdvyWsLQrL4/WC5aVRMHfi3vsN57eZLezVgMvRLJE8
PWcTzK7Ng/pQY6r5ojlkTQEjevjnU+UgkNq4o7M3VjnPzdJqh2Job17A+7SOvONX
ANk4NsnyAWeZcz2ItS26HaJYs8rlSnozYSkN+K5gdIjSV92rNSbtWQLJU2Pv/nmH
Cpk8N66DKOWA+NK7b43B4JENGaUY6TJNBmu5YzLLvs7aNsZSu8W5h2JQqvM604Fc
M5FqHZNbls+D8W4tbVx7y9dCpcOpCO7LrPszZzH7ypS6ngssmQ/rTsaqBxrJEIxe
4BR918/ZmEziEY2F0iqHgnio1k0ffhRVXUJYDmhxVOuVIGq6gJPiNDRK4ImuoGWT
FxG/MqOr3DvrZ8laOB2R/UtaPhppTvGvzRFxVnouxRY=
`pragma protect end_protected
