// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:20 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
s+7fisKXk/PqCtAcFN05lPWtjvi1iuXM+XT62wZMD8I01lA1W381xu3lBLCZhoMd
jPsZEDLLLJVfGkbtnPfNkvgIrS40GbrS6rruGhYrzH6sSyASVWcdtwa/794WeI+S
OUCHxMZ6jsEHZF+2fHEpStliQSWg4o+Sa7UCTURR3Bg=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 18128)
0dHGCshcCUtuEr/q7h/jKT+4gk1a3e/ubeMRhen69KjHpBzpLgb5khLobQwn4tfK
umQK9I2fNm2h6fDUUwuQ2gTSIZdtQV9HV43wXEb3ItTfHdZA38Fu0z55aR3yJB7d
WAzwmmmTw+L17ZNhKROPpt4XlOeXCgKgya8ppYO9Spzl7AAzFPkCcn9hI2XvdJ4e
sqjTGAChU3Qcmwsp5kih3+ige1i4KTWUK38X/IkfOn+0+AP2elKEJz2xHghsqp04
UQALLCFvv88+4V9NffWbnI18Pfz63LfkGjgng/x6zd6e/vzWxX11d+cJLzTCJkb/
Xh3lEjfOXk6gRLK5Uq2nAeMOyrOnUrvgzWmlxXG2XYdwYRmiKCT55YKQQmrhb9Sk
/rICHUkIcwvZT7wDLgo6ZyhohH/ozXqh0vBObXEBLks8EnzTbvJAlNU2Hh9Q/Vh3
wUjfDNHEoxFmFgP90v5MvVhApM2C/bS/mDarOOYfSOCqJAyFHBjn26TbsRGrlHRn
go6YI+Vu1MPvz5gFsCNMs/oWNGSuAIx0m/qjN5uRlVCjj/ido+ovfxJeYFpC2Sqb
gV3u1KF4/RmVNh/Pl4y1YjIYHADQTQ+pPEZLU5Af54S5BT26kDpC8hZlQlqqoGF6
QEoa9lQbnAT1rHw16tCWFo7zmGfDjblPf5HMa1P4vNEbgaDZaluYnkThxTmiyl93
PS+gtnQE0n5oIwvkzZ7iR3Qj02kJnb7GyOSCEYLqE084o/q2yK7esCIXc09LrF8a
UYG9nd8C0V5irGFIn5jzXIAamFA41KSaQC9/7iM0LlVZYl2FRmvUl01gnkCOBm/H
J3NvSauTzCqEoOv+MYQ0dBj9fyZIIu2P7afUz3ghOrqlVm1pThyTmMcbw8LKmC81
+kD0tuN60JzG3/kjnNQE0c3lGaSJZio7YZ1BL3qhfXNFbC+YZskTp6r10sAbghXd
9T+deo90M/2wrPceWGzPVfDNrenKxDt/6mS3XFTyriU7H7tASX4AabD+pNY0jk90
A6SDIFEdH4gizTbU+6VdddSjSOvYjaJuJtFJwpPjJeVW+2pmilW9gn5N+WtNWLHx
QyOqSUiJ6LqJR+3Hn1JJ0prlyD9wV+46OJqdGTM5xMlCpqOnK6p55m9RJxqmW8dS
vzhHej7wIglbfgVpvQ9tq3A2ovdW/hi9Nkt8GcOonLZKxdZTSKWzQCbYAIcqo16u
0q3AuBpIBfRIaSfXxo0R6vOhAEe2tkDYrEyoqKMwEC9KqeJB5j88c3dKoGKNokq3
bg61Qy7JNLz3rEeTM7gVAKwxdiZ/58vQSXAEq+YLdOV/910MIPy0Q0UaYpE7Df4q
h28jeqYETufGjMXTWRoH2vsK465YZx4WK/zHO8FoFb/jXk8l9MVnPcDpB6iPlofA
b0qdRV4Hufi5Wb8QQE5Wmz6OfKI5IdgOohmXBWzbnVu8mV3xuWrQBjVX0O6j233Z
WwT2S9gpKIEWx6eRQp3qg/6uXsjE/wHBJuAvcTys0cEn0aWN9upr85wVXjR+mU/B
mTEPWmi1Y1PEAFJXLxGvY6Lm7OdRDzwaBYFnGMERF1CkyOEx90zgCFufXYLkr4Rm
uaPtqzw3GIL7tnmYGdOpZczBKdTwNcn090/Bs4Z7Xb0WKDMyQ7T4yAoO7/1A5m8X
Kr+9mqD+pu2WKsrzPlb6wNLMBzbpMxEDk29aLX1hZA2A1mesEQzR16fFIJOb4maM
NXau6e0F8Hkfg/OH5nFwIJITg85G4RGSHEeU8kQyt04FIwRCJZmwwQKMywtNzRiB
4e8SUPgwc/MZU6GrCbP3EpJwMyjdRa5z8aFX8OE5VGCbq409yxX/dvIRKeYK00Cz
N4ZfTsPDxxJekc6e8I+NnJRBAyfiSA0FaHGFTfx14e1ZuZRrIrQ3Az6TDYeuyEFi
OoRLR8SKJuapXGneFTgubTYGyND70PXUsEyxSPy8fBYr3IV+xAXgp8w9ogRXIsZ3
2hLdn/OMKgPU98AYcAlfv2bH+W6eK9OgFx/yc8BkGal2CBbu4w9zcg2Ll/1+iV59
jtqDYV6FRvqFabinnNbm1TAxaOXtFSdQ+WmIElC97kbYIvEz18kuTdVgyAhjyotK
CNHf4mL0SN+h2qOvV1vADTgowMKBkkxs5NVl+zztWyEokEBxg4RGGP3VLrrlIkj1
w7GFzAwwFuWqgMH/sIsPXorhBV3w4u4hQObsMxMlCDfpZKC7PUUAtIob/ujhScO/
46uFG+a7NWD1AQ/PWVlt/1swPQUcHxAKEfST+uUYyP4gmN65L/e4Nlh5AQ4VaGfr
uCgmMYAnQ6T6lH4M9Uwz/qmFdd1YOHJ1w2qwApHSn4uTUnx7t8SCkLHKFPDZczPf
yW698lasQFRCLnLWEB/HYaHw7Xc2sq59NC6kRakFHWst/J75/3ur/6jBTtJr79ku
qHwJzHWmfUHmoIMG/5uKLIGY8/Jl+bICTxti7Fvn5dmSUL2DURkD1YLU2bTPsHPj
mMoVhS6pG/xN7OpVPkWUGMopGOA/SyFOA+EN9HTiA+XXpfV7UBgETPSP7bSmp0ss
zyzvZDIXNrmZrqYO5TreRb+1ubtfB2MycRnbbvVWGu5Ik4yFw4N7gqtWWJgEAGcm
bWRtDFgHQHudwqlFhD/fa3OeuOlmBHn1tnkZ3/rbG7HsHT//utpTr5aDznp6dAio
E934gYc6Y290MyLMpH54UsL1UDuYm7GgExW7uTShqFlSN9c76Cgt3uPUHHjBMqAI
t97JnugWeVx6r/otI9rUeU7v5cix9QzCt45IsVL8Hwpj4vPnqxmiSlmbaxLtpwWw
E9zDdaukrLjuuYhvrAzBGU6mYU8WW4kZS6G5q8d81lxEzldYeZh9QC1VVtxRz8z9
hRhzWepjNLqyZes6b0kso7dxc98Cl0M7Ff+/ugncxQ/Z2Qjyv5mlvFC7sWxsZ5EK
o9b+DzSO/dx8EHCQ9tD2sul6uzdo0fI9CTIXG2T7ti9U3BXRv1h5AxP2/arKb25e
MaUBRh25sMtgtjmaBMHSR8Ni04pjvd2CfwAU1EPSW08IPBPCYdlrP9TPF5GPqGOw
AQLrUl4msa8fGBVryyWo7EH15pcWjSc8wCD8aOQ4lkz3xXRr4+LcqVamng8iUTw6
qU5EHZl6VByltnNq7I/eK37sDacC+v5oLyv8lcyTfHXtfV9EMoXjWWuplkQMPSV8
LzqRsJElX7n3iqQviPea3AAFQ2qB8JT3T1X1tdty32R3XeTP2ZWNsvR/Duhtn8na
PkCN3Z9mRmZBpP8c7vy/90YslFwnYzgWlPdDqVW0QC/tYEzUkxJzpUuYBrwVtj4U
6hQjc5KJg5wQp4XKUxl6l6wGLygFLVJQLAhbDWnQs90WJxWHg57ykT7vXUe7jaxb
5Mz4IHxskPMxuhchfRX58OVMxFpTG9gW3qT2a5T39D9w2n5ech9j+HvFv5F9QEWJ
08bOktJK5P1PQ20n4I21Ecdzr8NPg1b57gY2YN9vyARFvZ+B7lqy5+h2f6PnEZ91
SYfoSyGi4wpTpEoEOqjTaFXqCOD1hHQmaGLplh6QeGrTOcl/YgXsju/oY1yT5sRW
gtyB3nHdqBCvgomnYJBoX6z6dn6L7btBXwOTHTCUy0JuprwyeepsehxII50pvs/W
GLXlHjNxJyD2J/7eB3p7yqINxfVkLA6LICndTPR4baFHU2NPHJtA38hvjTzkxl0s
kFCeRol+wGbj/XUAKGEsa45DWDba54OoZT6R1jZjONxVG6QHwtYiDiExkKY8t13f
vmlZiUnfjAdvQO0sf1m6Zz9hgjJD5ruDYexiei+hqgf22GctCVh4ocw9QoQQp1+t
2kB+cK9MG8shQ9OCDggkMUKxeRr6mvvvMExXX8SVv9ii/ePO3CL46JAM/AAGxZZO
+Toy9vW+1nfYiPR0Y1uubcVauwPI/pWmxgagyO5I9qhrvBFfPsroWNSuMDhc8TjR
7MLXvM41JCNjS0oIs9o5RXGTqeit5dHxZ20PD0ATIghgOku497htL+LhzkegRIpb
G3qWsd2zt3knr/625gjWT4JdEM2vfEccBEiny5nDig8Ir0C+hWX277I9HS/M9rI+
97NTAjLuXqkj9rWFaX7nsFZCwYdld4UUPUMnQPEQF71AVLn0g8hKYuYFhOtMkB1C
KNjsUrIFdKu80D/SvhqHbUuSYEHeRKhvYnn+VD2iO+EuBK1UnbXvu4SD8+79bPTv
2EZNuNgYowISA9djkgCwwIOvhc7lex6sRSBBpWSwBFf7wG28FAyl4gzE4+1b3Gcu
KwV4k9JGvnw3Ppi2IvI1//2bM0E4p5XagyxXEX/kpJI9bOXpxHojKNFtvfqx5nAK
W8ToHrSMA1qsJ20oicXcnWKEt2mOCr6eXwyt1+n2Z068ovloagJlni+8ISPstaOy
T4N/v3GqKxvMt1hatQIAKNqWPp08QQ/ZFlMNMjAJ+lf3pBOJIFZxlyDj8XCaFBIf
XqTR63ECLkYjXuAvPtwcLI2FRE4zQ2jUVzfqKlvUvqAKP0beVPMuEkGv2/Sinc7b
CoYJeCXdSGgKn1gWfHcWnasjMwM338LkIbWC4rOQa3h3JeLyDTGAk+ySQzP2zeHp
Owb7rLYQ4ULg6vq+8Ip7YyonvJHu359/0oSRHiLa1UJ1/Zl24pcEEH6O9D94aX1V
5monT4J6/zNN6+lNOivkhj2uRhx6uXdX044ePbJja83Ddsc/rb8Eu7QvjoXVnYlE
vSP4Wg+UbxAQSEqFI4j5H3SqhRc1hs2MjPYJZ/tYrAqxi4dvzG9/2nIQj40ewP3Z
mmF9PPaNOIJ/zEFwAgTWi0uvXP/PEKkw1fTGiP3e/wojaw6/Lo1Z6kvgxZ7KHHmr
33duplzFluxoo5rwGKMuQ6sZQ371zpfvm201IzgrntfW0l8pknfiw6Zy+JmhcErg
aFBgpI3ENOZPTmELHjTLAsHFEuXZ5Po6lEgnib7oFDqHwx4T1FPOyVixEBxWsA/u
xRnno3spZ75lWiY+0SYCfeouHfNMmClT1q/GRV4UpgEzB6YS32xu/8NYrqgzuBvA
65LF7vzUZxuV/q5Ks3fTOkdu4fTgN90JyWoZUrHtgTxI9D0qRjy3hrqwByu5d4oy
pas7CU0NP0wHHwyEl+mDgggHPlmlDlAFQwgSEDloPd30q2bG2QG7h72JPbTBavl5
P9nKpIap908Whw6vg5qpLbjGt3iIi1VX1/TiRXS9Fj92xz0TTsskZ2yuJgbJ0KkF
5IvbfkSLXGfzSX8geFT07B2oaWfk8/0kXrZBuoNiZ2UYkDtGT37cvgJ6sjbMqTKP
T8ZlUoAPCA7agUts9vISIy8UJugkF9sOnGuW/jq3k8i4g73xzzv3jNTRLQzhttDg
J30IjQORUxefP6ozqmrEsx6keAj/3vtmc9RXrYTvGhEBpSfkjxPphDYOPp1PN134
ISS5fQJNy+3Tb7zucnUp5iEx//BKoGKQItWJWo3w4JZ74L2Hlm9yidH6EdcGpI/i
VyL5pT/lsG0NHHgcQ33n7GginSaJkXrDsCEySOZ50G3PIRGJg2hVCZo0Owk1ZgbZ
Q13VjFpDEUe7ErlJk1EezphMLXDmXukT2NUZemQDqUKWOUgIsytE8bH2AasFLpE2
Oh21euJawJHh1XYdSRcW4czI/8j7TdgmipELgt3FJ42LH1TR++YZdXnlPlHDhCna
pwX3dfVyHDpGIhBFoVz5J/LXvP5pl7U6FkdSurTePqbTR4zRywCfC1zmh7QfHgmK
LvOvtOAR+dZC2uCL/IO0T6yvftMy8CBYCydP7JfwbLh2Ph5qT4lOeL/cBKNtj/Ms
DbjU4XM0MvttsXeF3xYXotB6xKpQHA11C+eFAQDu5AqIObrNOI6mXi2IDZOftbMu
uxDva2pND0dzHEzzvG2yCIZA3BVSyKPsaB+hpkyAN0iiZ2YVomilUQddhwGyERb6
80FaNClnxYyFszSzuJAL3LcDI3FiSOB7YuYDNPAy2wQZ/Rs+L1TEp/8stz+5uvpM
2JHrAGxzfqcKx8ccnKH1j32+skt7Nlkaq+ye3DPj5vpfgMOzfyDydzlRUyPSBDpf
nymvWA7+Oggu1oILOXLVRaL2y+ezpDLeo6qb2m/dZ4J29DM4S2h0V2NM/6r7/TRS
Ru7d2PH48nAEnY/6Zth5vu21rptb9/oEs63Nkjeb8127ySM0rL2f1najH9FyU5+y
ddXjexv7rfF/4MdIm6tATcYppenyNzNDQloBWBVGrHbkp+Kl9L2uxAAtd7T1sF9n
+mPijviY56/qmxcOhd9osB/K9FhWNtNr8urCcYxwFKNjVVd6ko2U3ETfYVoCYwiJ
V3EpGbSyh8qYcImFmNL7efuCxnCEfhWCpuVxbp42Zjg9pPPZhHONeABWat5fcPEF
Fiv0Chjqb6GMRLcNsmt7CrQwHFLxqoQyk1epRX/tytu9FV8F3poy22c/qsZl/AlK
BfLgSG0SLbHTiC12X6Ts8NgqhkVoxTkovQNPr7DtCQnrnF2MGez3YR5KPFg59DxV
Qjrn6CZCq4/Qfyvb43JlDYKvHXrzdfYUU29qF4nxi8kv8Ev18/Opsee5SGzCvzip
q1CsE1nHcB+xzfIXrRUPxj5ZIIWco/xGyyiV9MHZ0HelUfVd1XOcW6+N6WsKcVfK
YvPzOINN7YWv36I7ubHOifddM20EhZGfEDgM53QL6TQq1vYMDq+rFCGvw/18TU9u
eRZQK/q3qV25KktpnVG8aYspDgkGUWeu8CEz4qSX6lCPOTG3a6U4lXI5thptIBzP
rOK9qEwNzhC5rzt0ZhZnPtNTC9KmAx5eCb0xJbmXZ/Ul1sfP1LVUN5exUyCR+iKe
SX25iHNCaxal1jgXix4bs/+WB0GL1PqDUWD/s8FcJogbDhywfX+p5qyB2B1v2bp6
VwoZnkee+JZ5SvUnq/9Wwg81RGDfGEdvw+NQQwCEKTmVcJJ8rBo32C4TasirMyeC
aCGtC99Op+LooA2ACGepCK8MkDa0SlbZzw+B8KgpmudvsxfOKTkMSl455OwygznT
fimZiggvLaj/n1mU4BqWGhNFfqEpAAprto99fPDI+SxXG5OZlWQlj0xsDdiAzEQN
88ZZ9nHZyw9/smEqU7L+2c12e3Hv1XRlEQJG/13dQxHTNDxCF1NhZ1vWZnuitI3V
ddRF087kxk1t23VWy0xyDWiFLovWcS0RQvhHaPARhQufKeYR1oDnfYOiYY/uOpzM
QCwr3ETri483iZckjb0eVTdRBJOzyeTlvK5ehDFo1OAjleEvSEidQUwSrWPivN09
/zImtVYvgHUXLzNRYdaXS0mH0TDLz7DIHWrN4oOtJ68g5XtP3Cb71rPoC2+M45g5
24njoK5dbad1ABQ5U5ErU0oPPzkOnrN/h4qFlrBKy2CxLfK4dKblqmiPNmuSd6ds
VsiGgBh8ABIDYVyUICrlTjuoFXCcIxmKzaKDdGGR6Iy7+77aNOiIbxNxB/JzqGbB
dKXMRPxoCyj7QlLRhZd6nvGuQEHRZHEl9XivTaJGbO3i9LQyulEeJ3K3VfnF9IEs
CZHECcqG7bfPf3AzNsfVs82l35cY5sFVjOvfQ9NIOnV5giB7yB++7JocPWmTdU1x
9eLled5epMnU4qOm5nmoPUxuHzlUJ/dGdX2bwDVyvVn6okP3cCqjsAWwHsfvz+ah
hQ5sGwjJ63LeaW9yaTtx4Klck1XKBLSvbBau8wg0WivYrlZU6dhJvRkUVBu+Ssao
OsaLbeVACklONqHadXa8UYQ8iGF55owfpg4xo0T1dyy8NV2QLmy/HZe8TVZYsjrT
tdOnsbMvFKg9gzFA6mRWQ1wNl70H1Jw8U0ntwaf4+38B2onSDP4tkZ8E44rAyIFI
Udw0NrRATMhrbS8tBYOacF7qVFdhnkj3Ih/bBNiBgAKbS6X79+7a/g2dIG9TqYLh
mzW2f3PWlFDHe4vO5lUBwR3ljBd8YYvlGW2mJOQrLEqdA9ldzKydCM1YLKSi+EVS
s1fbALM/7jyTtlIts0zCGUwd8WlVLtAWifeRfADZUWdDxfgft0bOCL0A5o96cxBD
wjOGGEodZ4EoqYCpY7E0Zb3oCTGeI16Hi1p+sJgeBy2e2qg/25qOJlXVUFE0Qi6I
5LQMS7uvBiJ2ZSxtOgFHK0Mj8v2ikAK9DAU+/L8GVK4asdDTehZw7P48q6MFHId6
3R36MUm38JlTZczO2HZogh9cEaXaKG+sf4KjqfOcwHuo9BaRLNhlDvq2mqtkdLP5
Z/SIYGQRbFLGBtMIhaxHz1hJGRFbNXLsToQwhcpckkrJD/sFxt80YA0BfCLMwViI
0RgV1/8aXL92RE8eeEgxgZ79c8F5XCvik0Ez/8O/aKDXjfyvBicfvdBExSl327GQ
lHIA/pstiX+jrYDnEv8XYo35rII2XBj7i+QQ52Fmho4Cf4bP/uYnBsOuAT0aPGEN
VilNPcgcXYMwIGOop+mFhaObi90FAQjZa2KONObw4OltHHzUy8e7u+I/fDy7YgIn
CxseSa8in8Ax0Rcf0wKuzoTJeyrQMqHOtD+wj3lQBL2GSgSl6JxLH8HWanggzGnp
h9aaoDH5mBuzh77i/IpzEbzvYAgllogjOR6FtntMa8BYQPoLhI+aBCXLmDYIY76j
gWMhUSiHvX0P3iowZAi+k0ysEOd6smx5VI2KSd88Sxksr7N/+vmbA8PsjNF/i+et
tUNG2vlpumb5ypehi64R1IGNJpyJVNSY44Qtl/6BCSTPksKLAhyBz/dhxyFJFySs
A4iJKLPvPBiOsScJOEYuZAWD1ekOVTp3RfZMlnLyDJ8oOEAA6PHwF2IYeY9s5DuS
knMkDv91Ptj44IsJJR4djeeBV5L7IdgyrkVvKYmTvHihwdCoRAcDOmQOzLPjfHP8
Z33qtcp9rkwN12ZYvd0mN9Nk2JQFlLcbN0OH0jqCGzFbRS8NTnseg4ZcLs9reTxK
DUXAV/gxXeP99izXRfH44S6CknEeWPhy1+HoJinmWqTxj4JZDoXH0iP4X6rJMj3G
C34wguZCKS5KBsIDjRT3Uo4/XzfEkgTCHQxF+pGOllz0jupOHXpQ9/po6hMziujj
qsR3Nmc7ehIgKESXUZKtLxh3koBfev39PTKASCU+tjFwEREtjW6l+XoFgyVjcNY9
1wRJm0+eYZU/++H4zzYieoVK2pJhDzT/T2KIIFCtCPkPPV34H2JmZXDS8Og5ZDy0
lD6ktTR6300Gata8A0KIJFp4t9xdygCvYNAuYGi1TYY7lOBYab4LsEA7f8+DNLW9
2DC+qzbg3urLIFN15IY0MMzqYWUCICy1Wyp+7dggzhRdHECdBML1LIg8ESCsevEU
7m+bHJFsoHPutPqi0qQUUg5qFJVaSj+MHxf+082zDbgUAkQJGTvJjE3WC77tmQKm
uGY1BmZelu6W2haO8GGQIV2XXjGRHg2CPmiFOY6L+YlB0fQmeHC3VmIpv1/n9qeW
pvF8FQrS00kDJ2jYDNIiLUl1303oL4OqIGDsohDuO44HC3DYaIO7tvAY6+u32gtO
qWSoMUWFet06qJuFlQsSlZe6aumjyvRUbfLV/F2KjKdrAGtG11TMhjO7oFKfnyD3
ZxghaK9rm30tpDNA6W3nMQQeuACTVJuktgo9sts+nQQrJvSz8gobGzuL0b5SIlGY
Qd/WQtzCjYSIGwtnSDBQRRoD/oXeV5tZlZOEy4w9sZFLBAwiXCvwLgmWOuVv36X0
6eWwyyw5YMsxJvHYrQa2hykZEIDyIxuZ8o0HsgC8QAn7HsLaEDdqSp+CMWgBT6WA
D5DIqT8ZDRCxreYlMn1dh59rSeIm94LMjmIxuV6LlucoxXxrl5moEHhweO2AjY+S
dg6wmSmHZHW1RXhRXwN3XS7mRiVznktiNXUtGyY10zuQcDiUyZmq33OtT5p66D0B
CbUPDKMPP5xeD1qVVCM2ZqJPQX/rdR/2FyHoPR6eVHSwpYvOIFnST5u3flBSGPbe
EEj6yIHU8XSfoXTdgzAx8bg3mD22b5k0wgtjw6qRTLuiOlrKJZG2NjyNxAngYeRw
IoTyGcLEROKLIjoLp5ddRLEMjQUUBhHeusNps5taQpWrVc+mjOlRTYhyxVJqWMUJ
k4W1SMqQ8A7xur40AIMOziCKiOVYkVDOm/v7cxnsJKFX0cCw9l5mUpWLjcaR1pBp
8BFLYMJ5wV+NHq6tCGfXh+NhJ6dcbrYKOGnOhgVS9hQnk4l/sw3G/8wIwyWhw6/+
Y9plD2gRzX53jd7uJXMToyO8Gbx+PtthzItdpB1lEG3aYzC9OQ/nygYZmZUR9y82
193yOYFDnbtsVonhiddIsgPjxy9wiloIH1CbguUyz7wzXf6MWFjWf3FpjYcnDEck
Jga67x1CYA4TH9L+waSGrLRnOqAeFVgBvzsSF++TAkVrylfmwh4/8lcYPEvJnODw
yDRilFsotjh4QEbkPYJbAQ1G2bn80rn3Td31bn9a7s9iJTP/cceaUEMj6iQHtuO+
j0O1dvCiZgNxopXGkWD7+DQFCu2rnpDCBOtX/3jOiAJ4u5B5G8wPaxwcgRF46SDI
2/GlVKlXDoWcbN2hxXyn4kTLYmLZhtNc0WTTRVoZvtOVo8ngUN3dA3i3RiEwhaT8
bWNLX9x7yoo0IUsdfkP/ZeIKqDnbaGunE9Ufo+tcJkao8hGj2aeTk09oI/00A/zD
NVwzV5Bf1jkbc7VEwX6/JwoA1piXI9mM4PmlmNSGrLemv/SiYtpc21ztoOKFzJfM
CRvAXZTe7MFRUBZmzxjKh+926TUvhnEAR4HrdHSyDjLwKcdXnJIkqFsBegQCiuA0
KAJOprMR3QPI70cUk4OLeSMu+E7BsTpMQJsI7QJuSVijhOL+ziA78SD+1Umt1Naa
7jZ/J2vwhKPB6uZPSaeBYBvtd5VgSN2gRQD2t8S7xXDwHtXB8gl2Bfx2NQsY4q5A
my3M76e9I1TWfmYfvgTVi+ukydGUQXDbRMsziUR4joWRDYP338sZMeeAqG4bHhIP
6SCyP+1Ltt/6LTyTCMWOhdMQiarTlkRJSK9D6Xj4bhs4K9Y7wNixHNx8s70XbhVv
KSId1KOZXLIqYl9TvzXiAqk6qDa6RPCzktUA8FDIwPqgLH3mKGgbq7xy/RiDbk/F
hLcTiDqadtWLjXWHRGGIumDecnysCEP76PN6rJNd/GkzDM8J1osNZiW6X/Y72t6D
s8HdOdwZ9dffdRf/0ECy475pmtHfW2zMKEPcFM2XMAkpCgkNx10+GjAxsOse3TDK
nu1HivSr2XrzRI0HHpoM7eyai9qPSduzPv+99Rip2hUjwsrn74PkV+nkUtFp35um
XPO2ZK2aHlxq7ENSW5ZHJqdk9V7rhUbSnSNcyTEVGbqy0a5yQ6HgXqmoYE7fp0Oi
UiwQHXgUbC5pP1L9ojtuALBIZuNdo7iV7Ka0nOelQOYmFTxhpcltgHMd/wBdFlnV
jqI2TqMaMT2itVpQDdHkBIaUYD34OZwtBkm4NgtTG1x6V0Zc5MdnWNiLdlh6HHRJ
xmYXTvihl9+8TbNdaqiU5DC7vwTOawc0l8gZIGh/CVQ9iGG7lcUO76pCk/yorG+m
D3P9iL4P3whjL65ReCtfSWgZ8VkTxJ6eT3121wkJQSwyBRziODZah9fKyqlELoik
HvereImEx0QU5US9P8XyIYaf2Jij1fpQrf2K7NV07XnNRyS+ETeI6Pma/pTdo0Zz
HYOVSkOlIuE5MKqk/bPFPUcZEHwme1Jomjz+d/H/nSYfnysER2Ej5oDBVmJulyht
9dSig4wkUdXzO5czp5e4xNbNCy0zpLarpu77Vk6SXxCN0ldwYTUhv5qSGQv+E55U
X8FEx8lVpvasffbWJWMXzBqAJgmigp50mrA6lwkDRk0MjimEPrhth5qpaMGYh+gD
TnansGjd480xbJYahdS+u1fsl10PhtYo1CUXPKMkJhkDt2vpo46HaSpQVVPD5jDk
FbjSlQ9d6EVMp8oSP/1r4B3rah2HnPTTSRtTchoe17nrfvgee+KARjAof2U11nv2
ShFLetr8QN3dl1e/FT0u0lwOmMJkhdaBj+3yzKlicaYQ1yrQvF/bOvfWSujZBVyN
ssqK/jOiH1hnM0NM7KzMcossqbPjRBmaXbBryCPnxNMKATeLzV8IPUr7DenuY45a
NqSgMZjLH2wcNnciKitlfQ8JDokWviAqHrkBYvogzGHxLskG2XMa4YsgDRfJ0v3E
NHXnTEopbfuw/v0NLwmH/Nu9HZnTImj0EZMl0ws0eb60Cerv+sv8ifVg6jH6azg9
GpgUUOMVy9borszkS5TYBie1s3pFBqsdcPUFMek9xWB+zNeBY2++PzJkn5ogNr9g
8zBf+v7Nn4IAodmzCkcn5cpZ5r3czHxuteQ2uszw8hjjBa7miI7bWPZhyDcNgYPY
/pXOcRyexqr9RXBl0Ew61+XSk33WflO/gZrQkw9KWEZWwEKVGxuW6wOqc4pXpoml
FZQPpjYwYYX58UTzZip52B0NoU5Q3Or7gSvbw72R0lXzbLhXC2q43CxkUUWtx1fK
t4YKp02gZuNYZ/m5K6QM5B/aBmy7JnTw12amXP2g/lA6CVrX5Wd4twEE8MXZBv6u
FZ/NvmOWhMrhJpbvq3F/qpjubGEhbB4JmWwjdroRxOpmp2Ysz3DeDsVhg8WTpwG+
QhebPeKEDGveT8YLO7yflmICs3EhkGO3d5m0wXFoerEo/ZiIIu0zxHhBIgFknx7p
tZhzWHK+s7xqLdDyTQVZWVdDP5V8TN9hGjXrxpbY3gGcE5VveFv/xL6iHejCLJ6T
Q0C3qs/WVVch70oHhZ+WlpY6ZiF7f+J63NNN2X7B0ZbTDQof1op0HiqWU8CBzQ7e
pcY3GkhsTfNoXn8BrwYYzPQfRAfp8AHB6MBsGbJ2jY3JF82n2QuX798eoTyC7b4s
129WzLF0uD6EyFmLg6RFqb5oKDdSgG8gHohYhZPfSaEoTdx9rSadouwkAR/O4MP3
wkuix/u8+K/V/dLkQ+Dt9htJIz1Uwf1xTQd2vBgqjCriti12o0pG+S8bXIJaOO5Z
cYv0eDUcQ/9D65DpPU3opCbTd46NlaMKwBicQc5+5OaqfC0JrLzvtpVURLk/rrAJ
6s9akZHW0oVnku9kEHesFB24lG054egzS2Fm/LFFhWCYA1guXXDtM6Tq8YCZF7Vm
KWtUI4KkWTJGOXbch/GSYOTwCVXAV2l69TKkUvYLHFmgISNdY08VwEdT5gxTTExN
TJwBruDuWbfCf689Z9EfMyG8i4NTWJL/g0HPcfEd1NZhnKIyNfvf5sv9tvR2g7F0
rIqnXVX43k726u0h6XkhTT2IlesGgx/fJ+rmVH5luKFOQZWf3hK+iXUh/YczxLV6
Y4krhqCvMiZaw0neNKYNdjCW0mGlnCWXSjJcdWsXwGpRntkJhKrBWoOyts17inKK
eZR8k+yfmM7p8Xmj1Z0k1zXQ+9ByjdyKNs0fZhXWEPPfjiouGzEDaTXOPLhwjb/+
otwmIXGfHS7Dcw8ihJUhHYmvMZz3irn8dFcTla53tEtiF9aBk+73P1tQzdvxfO9Q
2bj5pghSetthuG26vN4rTKrp3AgflwjOtX1eysdYzlAOmBd/2x8/TZ9WyqAPjH61
kTEzeL9xq/MEZ/Belvl3uixQo8WoEfxUNckCYLOASaibCPItLwDV1UgX8v8Gdtv5
BgT/3B8PDrdI28WRo1dtNqSxWtLR9/ijOjrGdI8gupmK7Zfkprfyio5UweCnUstH
Uzs8QjLS+MBc/1BfRxq8hzo1U2b+Lh3NuQLlRL/yGPtNeJEO6z7+DE5K4sDqaWWa
oe61PtGjAjK5zcnbs/Q6o5e5UP8v2tL6NrEAsInn21OilMUHavUm9XZf0wICf4Dr
1h2do0ehWDJNypnTSvDoJ8qh4R3mdQpuEY6vW1xhqEhelnUSwPBo6Usbl4nZM3bA
xrGRnoz9i3+fO2Y5yj3JLJYlTFgBz915u/Cltr+m/2TwvuASYi3EYkB8wdmZO4EL
6rA4DKMXF+BtmFyGKT8TRWq3Tdo3ON03WfK3VY4SO+59GLrZ3zigk2zWhM0mx9lu
VPr0ZheUoq5uJ0Px9T+gdIZhJgh4FXDKyPrKg67XJjkQTiex/uwoqKIL6IP/4u6W
iKZmzE08Duz7XUqvyqfCTU/hCSWSbh9SPBn5PAco/r8iV5E3nfgif5N0XARx45HF
68BX5GzQwPm7MGXgEhNk9CKLWHTNui6g/XYLDOyhbg9KOieuy80HVsli/qws5AlX
IGijHmLt+qza6W0IE05LF7pu2ufaohKvirKl2fL8ayXl3O4I1+TyUyi8gPWaE3Ff
QNJb326wE6axXstsfkgFuWy/0lwGfAsu9ggl5hSXCxiOt+U+f6blGUhVZO5DwjGr
HPbyS+C+byPZVpCg0ehkHFRhYFUQ8fxOS7lPAIk3jfCv9Hj78f7Mp/mW33eI74nd
T9xMBTt9JLEHFxKvXnI07FwL9Z2rHReZlXn/IAynWIiHNU+DrWQu3xxWzH0eEU4L
Lr1I8+uJElyR5F3OkZUXk3MubihonZAesOp5hW+uQjMDrhkw1pkBneO0PA9+K/jp
3YeMZ2+F3xjBdz8FRI+l94hE2ZKpApndvczIArhBykuFdhuBnnBrL6UwD1eY6rsj
PzDNDbX5eSVpLsXf2miqCedNaBVYolpU+xZ+rQt4rGnSGwe53BIHPgdvVLXt2eCA
p1s+ePsNJw3U2ZdL9XRMkaknZwZxYR1W/+csiegVKFItgDyv0L2ueh2hHpi47yBO
RaDpY+fGFOtVtuh3xxwueRMQfKXt37YpbF73M7I1EsPgDWMZp2N5gRtlJjb8CNnA
5vIHvPazXaTO2TYqy/IlJ/55wSKWlvECGjllT/vRrAm4wCUFMvoEpBsGjxNUjlNZ
VREA33c5AxzrAO0vhl6eRP31jcc8p+Dr7NfO4HO3a42Z44DBvIhZuCNKqoPCJHig
rGB/IzNSVsQBRwFwnGd5NhLhm34Af903yq1uW/8G5kWoLQNzfzE7KCoVQgVe0OoT
d865uogev0d7kmkKP1MYATFXnsBFW2uGEwngQzYdjrlM49PAjRVNeWSMxkw+Qg5I
DEd9KrFR2fQeFH5dngFAmsME4jbHGpfgXRk3tTniDtncx2o7C+uJv6jpQoW+WVMp
im2sfcZ+VgfgypscY9lIdaiL7sK3X3oUvmNU2RnR4PpMmzq0mYOhnf5SyI+XJ6/b
47RURvaX9tkTlnd1pO9vzmf6mDLnV3fkDPU9rWAF4lCbuQZGSIgflW5+xchECOVF
ndGOwrHP/UbOggSOo8/F9H1c3ig3+cXSIxXfC/FTN4hZcJAfT/uEOhhUKJAshS7o
6yGRpMCSoeSx4vyc9sbsRLKJXJ36Kf5wfWZcxY8/8VA3pYf7Ec4ITBOiZ2uyz1LI
yA6psdTyWVqaTA4y945PI0qIJY0c2dSVzbXE8klN3DhslvnXYJM4TRD5bkhCyS6Z
/DSIDELhjVe5sxscg/AFhPvwO4GzF2hElO/8Vh5PvzGPjwUgaf4JDZCyNg0E6v3h
aTJH9Xb1Rge/crliJGMSx2PX3h4osXzXjIk+RgEIAijYtpj8YJV3/eS+Zl+XEk6P
icINTZGg0e0cqsAiTL4Xb9idqtSSrJh+FhcZRNLPANDCBTKPJdv1wmMm+vQN6iHr
Mf5kY+ouqfmVRayZcsuXgEmvn1yg9qOvWn1sG41wnh53lYdbf6eYPhJ0fvBZnnQ/
++/soGCM77mOS4fgFw4hUxEq5dJAbMzsDvepbV43es6dirLH1qIvYeoqvfqEVXLs
ZVzpAqICgJuugDbZ5CBdu+KC5hRQ8QkR40301emqqZGg6jL/RgqZhwg8SefAjN2A
gLzjyMC17R3VDNiEcsDOuXMe5UfjF1Qh2KdVb4ydU0IMdDalsgPo0BOsJ1t2pPdn
wt14JTcvvb/HpNT5VpKd0WbxN4c95521bRvQga7OZmtcQOKbsfgk/gEWKzA7I4Np
6pkT1escxlkolJZTdfaClUd1oW8wkfkodX1ngNFk7T3YXfkV2qkHnG5t8aaJliGJ
RcwjjBdob/PWq01zpX+LA4eK5Mt7+gRNMOL+Vo6cV+JKuY75d4/jiR4J+A6tfoI4
tY8LQ4l/o46VYll7HLoADIzDCNGW6lHZCo6PP9jrR1Gev+6gNA/lewGvure4kxdj
2x4bcfpDnLijmMYbSdvRBZBRep7NBfK9s2vSZcScB2TR6bU9Jucp54YbYZIwePPm
xkKHaEHsvgIpzO4xysMBHUs8/x8NsdyugRoPozW3Gd/N4D5NpYGYRE+1RDebjFIr
mC8QkZS4MkbT+pH9ZG1S26b0GJuuifB6u1wYFEBdQsBZO9I9wc4KLHHCHkX2Ip3o
baOnLYVWjA6XAsh1jpd9fsMe4ms5IHwJWMBrULAXsNibiZpMrSQiTwJUNHPc6DVY
7/P82BLvOJN0LMW5IAT+kdV6me3m4nWB8MHJ/DcW6MIXaAAlYhnJynQGKiMB6NYX
KWku1EkR1YsdjTg20zn7bxaHWGkXNaDEh2K+LrSEr4T2bLtkNPB+vKHdQrGUKb/4
yNSlyd94xYMUJzjUh79U0/833+4+PBgbnf7+a9AVA3NpbKu4WX8gurfzHu7QE38g
stuiOM7P5Sc6/U1TbcY1BCFHruaYtKpZxbC020TKvy11AT1/Xv+OaRJ5YzCKF12g
Y8QmF4ZYcdglOSixO09I6YJ4URN57cLXHaanFWeh6E90PLSwLxBvFYeS5B1hJlC7
1VbXRlK9TGeu2w8yZGGDOR7NMUJ3lZ0FQDsXvSsI6nZTMB+eWMvHtrN5WzvlHhN3
f/xYf6cF5NYF4XAI7PlxDrhSqBKEidPsUoirslZpR7Py32A3jgpXpUzJ6dO8kKdU
eUAOm+Nedvsc6ZkxwrLcYs3rJUbWI1teWiikuAbazfstNf1dOUMl5vRyhkNg5JPE
MsxFzTNCP06m46zVwfPQf74KBJqssy+IGy19N2oyay6wfs3/aQE0A+e7bQ/PEGiI
UDmEgghpX9uZxIbYts3Gvcks20Hkrf6YRnF2BItLFyQY8rvzNP8sov3BPSn4rle8
6HwEBDkm/FY+BGru7ONE93g2RA48f+2N+ogGIZImkY8ceXgDQLtVUEgCIBDaCU4M
f/E8083eleyl9U/JUp8RUgSJCUetM+TfHmrkBelS+yO12vZuh2h+A/bhidkn40EG
SRuCNIzjrCObhQQd3uxMZIzXJAXwgjuiQmyyoiEaTh4ujl+0fhxb0JKC9cxKd/xc
Gw/DGDeo1P43BvpRnldkqT18OISGanQaNkmEn1+755uNUciW9Pe22wrrLuwbFWsu
cYP+Zisq9LFwg69BRP2aQssCS+SNXoj2eVGy5zYiXVy2lZsMTqbnLxmzYZ54N8tW
VIWwFE8M8HEQ1cvLlzDBkzVZ+M2z7cy7Ovb13s1yCuP07pWQr3s4sAx9MIfsvTDj
M6LmDQh4RDO3dufmwi/+QsaPhKFuP1H6MipvyuaSzgHUWlI31VVKC7q/fi6cghPe
NFDUDw8KT7VkxV1a5wIiEbXPCJqBTbDqHcJBI0tFudMC2pPbYsvurTPc/4qzTJi6
5GXu3Fymx4j2Pv6m0FiWkRaQp3oIsF8Q8cDKBtSIYpwdOmrqfmSpikEWnE5wT2rY
akY+zhD/2RHgoBunlmyhpZ05FLPhciiiamPqtO8UUHEIyYpZ/p3TbIEWVjQ+2TgI
VWK3QxNw1hmZZAyLMebENPyD++5i1jggniFE3NuI8ZGaW/dNHqqZca3cYIQJCPs+
yiqYC+Pee/7n3Wd5vMwpPCI1ptX+JM+INmJ+4+4utJzUKPB7t4/Ng6r9hkhFhACV
uKZXjwL213YjDndiRvCwm9RA0sTD5gpiJYs24WTRryvuZuCxSwUCeVo5qFH2RAKZ
DwvluPZd4syQwPz3/dBbkahyY5Du2ohrLjaKZ3t8Ya5OjPKJXRsPMVGehPIuvFcA
p2oF6IKk4sd/EBknf+YZiZTixEPcPog72MhhLD57kO8A2dEcA5SpCD9tcRijVOaO
esq7otabbMAjdhpcq3mZEVLOweWecPvvfYNU39eHrvTirQMamocFvNbhShD5F4sH
z2nf4ppkQrj/aJszRvr0MxtIUBRQnhWSyyxrQ6xvkJDAjGjNG4pgv6iqJ1kpxtMa
qe94DLcycSNYHJ9GVxJc/NNW1QNUdYssIgNzfZ24Om5LPQSgiYFifCgzGBVm6gbd
xBe8XRrV9MXCuZErou2nFW/7EfKiFnCYstuc1sF+3/47hNKwMUuTu+OJiWXaHMcc
hFAPHgLaMPePXLErd5BlSG2XkZbMUyJ+gnkkFeCJmsAW2KAua0PxhXk1EW77Fnhf
Wk7fctWi9RbOvSjT4uBIEj6HxCfmbUhPSRhjrnS2UtlEOujqvC5dhZs6OZvCTfl/
YjvB3phqQtsbGVzKHJBDsCQoRDQgYDszCTjOg3DbUjUyfEPH2gYEOK73Lg/dCsoK
kelSRMjYaqLKIVt3xWmDRxy8Lv3Q5bNydN/wIjA2JV+fA/xTx09XPQlYAnN4wv49
K8eEnI6ig+L9SW9YPyoH1558T3eG2D23rwFjJm2apA3tLm8oOuU44aUbUuhyUgOB
2Pphl2q6SmupkB705I/uxJSigPtFjXC8HvN/caDbo01dqXNNcd4yVE1XY71FMAK/
8CY6d9dqUVnOCDyFsIXN1EDI85YXfBnJ8AB4Kx1vQGg30b6tM5395+jjLq8prQ6k
hUnLTK/x0XfokUOkBGS39apn5ctn/ESsIoxFh8dVaVth562HiyuVuocCGkxIKLAf
c/SBAogjQK53guHhB7BQHt+iZDIII+/oM8NF8PFkgOEcQ7+ysYF1KEKGd2ZN0u/L
Fiu0WC8b9gN5HxNgo0jxWxOw++2ouZ/lupFKK4NKmqVfYf5HCTPtrc8xRC2WXwWD
NXMj8DLvl2JTIp7mYwDoZogCXQcZm78hreWiKC+y2dLcpQ71JtCuoWppMytUltMg
IIj06Jlab+l/llRD61a3PQOnw0eVXhFCOK/HS93jdRbBZ46FLO/PL87a7upTKH2m
ZuqiPwBYRjDVOHbkdL+IIuAssI0aCXl5XY1e2hPh7Cxd2sT0KEvBIJ7IL7JJNgdd
XzIJuohsW510ftPRYWsbF0vmNDmFoZU17Fo/tsXIgMc7BH6s1/WW6++zzOSERbT1
N1iHmxpGAdUEF75RdUdeuA/mdWV2AopXUZBy0GRWV9D+H4I2FN2gcpijojwL8H8t
vJEx/UYp+hcv0XkAQ2sOcpXqkYdZNSejC/86XS03XYB6neBKbjHKBIJlUzHUzMto
qkgnpN3QbANasBVLM0eNHCYcJNF3Rc0vuEijDF7kllv+FLb/FXXfzzlckocmteWv
jOLWQUsevWSdGJioBN+d9McnWOSa+Mp86joWzGG0qE1GEUT5niTJYCwbYL1TFjyf
Ek1mJgOI1C3UlsF1SWh1684d3fAaXhTtDvI+9nuuSZkYkkvLXNxVr1hv6SlihjLo
x4bQtTOpRlle64Dav/g48ZplaAXFwEpI6/Xm2FfVsSL7bVIzYykyqCwB097MRXoF
dNBBOzYgeBq82wyuhwgG4SySTIGNXeKsWsRhsh1E3XoGVnPGI9ywKoZ6th2vjdAw
tX+KxBa+zNNY8MqtuUu+pA/WIoQ738c9qtrDvKIrWZH1myD+UccrjeKkyjDmznGu
A4ater50axVJ6grKjrEUkgfnzVEygjBKi9myvm70t0G/ZrjVcApzsdBkPuR0PaXH
R4nlMf8+/oSZ9g8iN7S/mF7m4rjz+0Si4qz9P7zPb6ByDK2qIXMdEUq9KL96smwj
6DvS7mv9XwIV7qp6VgaO2s7FKYfP86Ob/SMA5bHFBZILH5Zg5yL7WUdKTB2VsV2l
GALvrMkaIe2PMwuO5wN9d6kNTwXGK9bkubtDBma/GhM/fkDnaQMb9IQa7AxzRhe9
XjWwbFafBNpnQRXPDy5DevXuvs0xogzu8OJlmqhYfoQw4x2hn/rbohAeFKHf6wFR
4/djy+umH5+qOx5YezEwVWkkDp8T61X+uAXnT4GhnownQenlm6td4IYwuj7Pmw3c
rP7Gvwc0iz8e3WxlU8636Uug9+qObMkfcSgNbvzwyApNJxnFhCpl6vcHWpk2+1x+
fAINURKI6KPBTC4rQLV6r++ht98pH2XnKE/Ng99dnho3hYSgVhUrDTMtAzhMHkao
qMbtUvntMBoA9TrH0yTFlxPSHPjkRHOpBGMkHS7gE3HP2eofXFoyXrEI2LwkZDPi
VliNw2oRPxC/1PRRPUp9MGFamhi9ufcZA2ivCK/P5NqtcaBhOqZduJhHO71bScUv
QBjmKsB/02lnpLx4mGBR3b5rpJreSgNhXQZrDAB9nNnGOn5K4Urb17xwaY/OEAaR
eLvGlcGYxyhpidRgdrTtbzZsJBlck7ClAH5PXbC1dA8vuSM1ICmJThy901ajR6fp
cKvlMe00dfK5SfrpjmUcfp2q/+bz+6GYK9CYQIvpQiOIgy5Fyk7YfS4pFajyz6wt
DvNvGnB53jzQJXqHEGsJEbXL+Z0K1OMCiNi2y9BRECuREKYlcS2uvkoTQa8X+9kp
OWYgNwV1aJAgpO8PCf3LcXzKElsdy8knmkAx1obi061SYkakQF55ZETPcycJlv8c
aY+qs5ibemFh6sWmYCgnik+grJN2bo9TShq2Q8Ey9jnwrPX/Yeq/2Ui83X1OZRN9
nUW/1xaloqIUi+ybhS4uGqrt57V4g4lj8cZpehVqc9r1abkvv+fuFecXY3/hnrRx
M8Pb0BquAee5Wei9LzeayjlnVT1MZvYdQnXjCMzqjgJ570bhST1rNWFjQoUQdADi
OsyV05t0y9w6JKuMXJZiK0HFqo13Uqx8hbqFulBS29yfMLfJ8pMWgK2Kbf3tZIGv
zWSX3iaF7OZydIJZxQcj5T1EmQVR2Z9DJqLP6Pa0HHN8SjbpqqH/R7tm27t/+q/S
1PpNW0llNAc0xY5AduEGgEsLhu2+iZXARgLhUBiienCaN3OYHwMhed3BDdwMUz03
vyE0ePvs89HMt+zIv9p7pG2QqSxBh6ND/5Sm+aOg4n311HYH287c7UmV3uMDIkag
gwX/nCmgEvIowOzk1eRE5c6N4uf/dDKsGvfzm3ZIjLh+K7rrF0ECqdp0LgLgY6La
tyKCudR7sNF1VfZLqbZchXV0Q2M5Ed1jEzbCm+uJMNadGnDdzwSZWhRYDkhKaqeJ
Rcqe4HbAIDpw+8lNW0b8+vaPuCGdJL6ZPYd0fkkoGeotBo+nDKbzD0WEKw4kVZe7
ZIll1w10bCZAW5dS6YqT276VPyIHFR4X1BrrY75nwJWm4gTwafblj1dOPKZpAGFe
WEQfKtCLZh2oayD1S6I83jae+9W3ZhWXS938qXj12XIzI2n0xPKi17pf4fXaPo5W
+kw6vTLtHl72mV9rcJ9OPNWzXqKjSEq2RT11U5st19fJmzkA0ysqH483Y8imOtxC
en84hC3UCXUJbcCnieKLr3v/9Q3aLssM4ExJatIabQyuJpP1EwbDiUmqk75JN8OL
w62Zk39DH6kqXkgc7lhaLeNeTy5xMHPdTG+NqnfJVl7j7Fcjl2DvcY/KMlR2etaL
szUO8RrrwahOntUISA+xLogxo/cdIA5elmDSz2dN3GYj+zjpso+2MRZmE74zJ8dq
Q7NEcO8Z3Vv+CQf2oIo6jV/ih8s7RAx/u7Tg5FM3YZhxAR53nD9B/Lnc7V7kDCtG
JSh22aV7uIT+9MozgRJ0deR7fLeg0qqpLas5qzTPovOtSYzyeJ/DoRexfoJ3JFlR
XmDlSYFH18VqOjZ5IvgyJSrXq44c47ErXigZAO7N+qAR2Do3kmOVAmv/RSdF6kCs
CUd4w0i6jiICie4STtd4B3thDEqy5oI4v3AjOtNFsyNiI+OO+6q2eJEB9ztaV79e
q//y4tEH9E8uZVS+5qLuQrszl1AXoUxS+MYmJvgeQSC/8pfQ9Ut6odPGLPxyEekq
iyiif1d3iuflnZFgjB/qHORp8dGnsyWwZIavIc95ckRgagDcXo3K9M03O5r0HEFC
MqaWoyP6cLohxp7ckzeZdh5aLciNiVrOmMRBLppYEhkHZz768aT4O300tWuH8EzT
i3SUy2F0U3RYKEZVwSMcQvbKdTZMMBm0u/X29ekFU447MY9etbNJZsA9ItO3g/II
f+lz0kYJwS0Azvp11+85bWxFGRw5JxDa/rnLLmZ0QcsaX4+p5t+1DW9keybimpmT
c0qVV9Xe340aSmxrd/GVYxZEDWwcXiY2eHNcekzj9zmG3z/5kdkRSaZCJhjataRb
AfJMBFH7pUDubsB7rJmUQcPkAJlVLAmywB8o4ngWpbawI5caxxX7tLZ739o0EVnW
EX7/DBrhc2mDCAk4lskrzAWqqx1suxyg8SWzteYPimUu/icJrKuaxkSHL8I7w29P
JFREu8lTXzxF1yECQBhd8Mg+NOpDoYdxFASDIKXzuqKRCeFQRgC3dBV/4JGlRtUd
+0kb+Nr1fhNLmi1LfqTt5+e1rW1bAhqEoj7mtL0SK+2K4G2EoPwjMOZAfaACYl21
xpnlzv802C2LYv7Fr8++8LMLV5IHDJMQj+fr17BewF6MvJ/CEHdWvW0AKrOmED/z
gW3QnUT7Om5aBtLjBSjqQh6o6gmQ6YRht+8OuDfVWmCdzJ9VI82sHZqw25fsxWne
cGkWylwKFhLxZqV1rBvg399w0JYeBl3SSXrG+TV3vgoqK9OIhzXQf+CjNGnGo6/5
oEizlppIz5HdK7JaU2lZEoT+mUk1O38zz3F6bnRungzfyyfOh6mNM04zz4rcja77
//7xA+ejnUX38HWtX6JLdslb8jZ+9NC5b0f44qcyKaMd9vHrN8m91F7lSs2eP5iR
TaM81L3t3YQYJ07jKnFYWVvrxZ8E6P+rhFJIA0cDCoxi1QIJAx5flG6O6lnxG7QX
sJt7IRX1mXs6/zK/u6Q8T18QHik7hwg9DY5aBC1nHPGiLgZ0yhd+Fqb/88ljSW5L
jMPtDq4n3O0zrEWK4g2N8YgRIQ5/1JKDEBfnZktoKAA5AyV5smGXU+T9U/o810BI
kDH2+NM+xX/liAtP5YjjwKg/m4BkCVVdvrUdokS2cO6Vdk0jivWmFKHa0ouRypxL
jGiFG3BvKKaru5rU6GOmnoYlml1QYp6fdFIii09+CK3SJ41GogwztHIyjyxaPM9e
7PQMshHpl8IcNyxnfvEgrVP/nZNnXqFPd82FRGdjQp8SNotV36o875fdChwucWIt
knMKKLlaRKBm0kL1IkpEHWv0+EsB08b0JTHJtHafnhUe3aAbeFMdzBxgwQPb2qxE
mQUOu5EHQi7zjML9EEQM10GaFMLF/DpLEbnljYuT6SvOqGntwrYS45+NQ+sLCLZZ
nGKDBodzYSxPiNiEBirpA7D7sJgtM06+klOQDk8FGh6DVYk1n0XBEkfwYGGlv8F0
gNoMsjvUrlAlLFgHzUtYYN/0uHGKeoDsU+JQcYT/OCGNS9b6Dca88pUyIMRjDph2
HNdxH/6tnVIaRBGhcT2aiZ8mQ8Ic6nJfZQepiV+ReuU2+2FLgmGCOCafDci0Xx8S
wsjQEnxcpqzoV2KWFqS8Kd12DznIIQNUmcHuOe/vYeP8auDKqC2SOil0BDy02FSG
AjaavyAMSwW46H8Za2WnmOXkIEtcczTmXNWUjfoZWQG0CWJVazMUW+68zYwJdoKl
9y7tcON9jJ4feTC91NKHNnwQGo6moG8HiyzHCAuQjkJf0OxGpQbJgWiWN2ksWmBr
PT8aO8lQ1wxekyI1907qbhMpv8MEtssnK+pI++EYxI+hsjcGc+grthkROX8i/BV8
JOItjEBe+9QpLYvn5mhYhEwqbUFfYC79gCSXm7jsZdt5dFPYgziE3CSYi+MDMboD
UJGDziH454iqGRertgueyOoBR4sXGo624gJkdv3sYyQ9VoA0OtFWAd0vO62cAdEd
YzjvF0rXJ2WbO1wpX9D4R6bkAfkGAgwaibhcJkuLuV+qQk1YCTOQw80kAbBrV2fv
rVoYCtQKryLPUEViUE7RhLAsHecLeoJWROyI28J2Y72FNHpYxPO5UwWuuDL2O5rM
OGbU15ON8Nu06rg7ntXsykCEVGIxNgeE3pNBGuN1ZEw=
`pragma protect end_protected
