// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:33:36 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
tC2hM2e2K6rcfBVwLbsMlSOWyNa91BTw4+2lssSUPVkGyLRKgpfcpnXOj+qTLxTw
Pc01zLE3W9IXBZsHlk0fc/tqVoUFZaTiO3yhS+39cZd+E6rbvZdzG8Fq+1hIexHo
BzxltGz2WTGw9LxsAdlLWSLEL7OKjfD9pOF0nuMCMcw=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 26736)
Pl1a6Os5IvOkbp/Dw27uYgG1a6LjAlRsWBMJ/3z3Mu8USofbmIPTqubg0VrCbtYG
Zt9Qbi/BP2vTglc3uwOX4rwRa4BapWwA5aORRdLju7WB+O/4RUJ3VUwoFbeLc9CQ
RS618aUsmz9TNyj7KzscWcEoYP1Sv7A5O6Vo5lZTunILgb0jfDjgCpSUgMC0cRkF
6QEGxpiEIm5jouvWtpH+67xCpJ/lltjHzXZBnbRfPkOvbXxPmK4BbvRmOrZkpsHC
gU1ysvQumfz1/cPW5Jfxt/rgv0koVjtrLcX7pA2HvvU/SxIDqUndw2OpyZVD2/OL
Wm7kki33wALC81yfrnPPgxUqgLk0RAompHSx9wthfRwAlegWoBb36pg/dNhDDaTu
Y6Eeax3zOPqKXw9nCO9PpYxLJ6ts9CWzK9I2hllV+/Pi4zNV0BoSM3upE62Ktwln
sJo0uUhQxJoTcR8XHuzEHTc+f/c6IRbruzT3MDRvAhUlAUPdczlPyLa2Vh/K8Fnb
dVmCxhC4TzcrkZiz59NFX6MVUpf9QHqL8VlGNJ0Wq6y+qBuEFAMlwdMRX+P5HQ+V
EQhtDdenY2r1G8qPeLG635pLS8lvT8XrJI7ZjWQ6/UFETtGSwmynT0J2GVdDpWwM
ZL33HEI6F/TcZoQ33SKm7m1LKSDwqfcaYhP1OwObOyUo6uE4DNChJezF8ZWZ73m+
8hqDreSjwp/bNeN/O8MnLrK5vIKzSwkoe5H7VFMJRfM9Sp7eOi9zJa9AXQVY1I92
EITgA2yx1B1bTMjLdj2WOxEgqGoUUyBLduFcYyDBfBqVwqn+8HBGNbelCRk5z4Cg
goghPd3ujyci7wL+k86YqUTaT4Kw7ldfT9Hq1XvrhNWHjwfb49/xg/RqfDltFk+m
b6XaglJngRzuRsbbNZcnRW3bXxUftlhIDAM+GaqcSzWbTdieBsnCVhrYqkj3SWNG
MPOb+7967AS1mozfg4jegITbX1f5DjUv86OtI/tw6jFzOjeIOS7luBsJceh4f5jg
goATNsmaSkICl+aYIoZVyIQ7+HmwIxXbC+v9wA0tmyljzMelpaHEKZYISrHdu0xh
a6U5ePAINcc21wr7NuodDndmtmT1OT21vk/sdTY1W0KHU7FnOnApb1SoTEOOgSt3
6jsGIQCJ7wIL2LMrrzoyxxQCp8mgO6Ahx5wJ5QWzYVe3bJH6vYfx8OSI6wzWOoKL
xk92ALiIdsBRcBH4cRTARMOeJoxk53BqCzeutXKsFUFZ4yQEgsZLANlntmG62lht
2PTShulwIBDcZZhbIiFZUuoRW81LIcornf0+CdovuDmTKmv3UzYAKPg8/vof/Ugl
PJab2CKYBdbgNY+9H3aFcJ0pb/B1O0z9sRn3aTrSThrQa5DlLH9hJw94fF7iJoof
thvTz35sx5CvtRUILphsXR2rYopOhcp0BS+URmxvJF9RD6D3QrSyG+9LyiupEwgK
ilriDmQbfEDX8lZswC6OFzEdzJoteYKTyLafJVFA9VUyskADIDoYXgL7uIWg+Jdz
3xbGTUaD2batv1cWEfHZIUYyP2ndpa8k/Ym6erNo3ZojFRhwwsF9ZeoiHo38P//K
z2F5D6nTjtEeBRsaXnbOjyuCHhWkNeYsL+7VEpsAVkiRgt0si8vqzQWn2YUvDmQt
O7t89zeZU8knsAFIpo5zJyC8noP7JZ5xRbqUmiLn0x6VIzWyEZJfyDT6A3fbn65y
Yg0A8aXuxaNf6WyxgPpmo1Of5PAw0QoMRRGNY2M2n9UQ3UgPd6cvlGRk0vV2/Qgh
dLFxcNjzgn37+HK6HR4JEcyLe2QOeg+JOxGX+c3qkBPta0ZgtlOfJC9AP6jU1Xtg
Ej572G5DpH1exIxwZCg8loUqw9hfAe8NcZ9TTfaOHrJdXz23pnM4rxcu0VGKOimX
zuofX9tHYV5JR3jL7UG91HK68abVAVK1corbTjVWYL9FIgFletffVIuuVDi+8nY0
Lf536FpdeiNUEkz6qFrKnXvuKYR6w/H11j4t7aTfvXD3zeIbCWzCvnn1WWOX6l5j
WEf4JSpCiydHzHSjY4HyACtmnMu7ZyQjwe4bBhTG68FOT0M/3k2ISNp1Bv8HLJNc
9kiTUOv6Cg5eh4qChw1ZA+hDT3xWW05xRWRYI+bifEMSk+SujuIYzdmlhcj5XvNp
M/BVJetbQ0u6waGAj5wlL48msLR6zY2JI8hzsXiplTIb9AX9a8YzWe5JAfIaAiCO
ZGnmRZu43CMpmy137vnxCMtYftcP9bHV5uezt/iBAox7+hQd0+UIZqJDZzC7vbEi
oo1pHqvX1a/+7MDN6/B8eRBKJjZnxoF6TWYnhpPsX7utWrLbtYJBCL0e136bZLqI
SqYsM48as81evmUDoEmHXnSFd+cQ/vWZUskWzOsSwrX6CP9BzcRX9EVhiGig1ZLf
mQ+7nds5rRYiXA7t8hieGaPeM340rnD1zR5qPfrpgJ7Bu7ZzvwWFOyZMNVzQe5xH
WyBP/3cjygrDv72Z5tGaw2vIMgVwLF18ZsToSk1ndpl6bWcl+F5wgnCyivCcEEJt
9y5TsYvdI6twnmHfY3cCd5idHMGo/FIri3RmTYz45EQzIdv77ftPICnGk08yCCAS
IJvrQlu+HMCEzAykeTY0RTqWcuqpqK9BXFfPRSOG9qTIN3Vng8XfMnFF+KJmYEP3
P8uT3PfoCSt4qyQTlQXZaDGfLiVY0p4Mgv4dP9mIGv1w3l8x3F9bAfXNPeaBFa9u
wWWhSaLQqSdzn6ItNa91y4xRQc6U+ADhjv0saXWk0Z69PaTk0v5eoT+kc1RngQmb
AO+2orZwcLBCc9nhMishl94TFe4/QzXFpnC45oRQJIn3oISCapoVQhB2yt3DQlkJ
ehisM9+fn5Ri/dkcUZJAacfHqtR5ljw9U8mP24d/uAxZ+9o1vPxzhVi7np81ZFjI
wKF3HdVdktpcteepxLzCqSAvUadC8hyxrNMhgFt27V1+Cyg6Cpb8XT+OEJ73nO+7
EeKH1h0f7iwZ+k6nnJVOilFkOIcQu8sXuwm69xBY1Y1XpJyuXBjHJZgPU1FwITt/
gAP0LEm8HpkD5WzAjlSq5nmu8piTL+D6UL6DrFK75C4otcY/ISNfhkMw4QK5lK6K
GRPXo449OzYvqRzcNqxXZBJNuMGIgqgteDy1w8JTZ9f+iS6jcE4433RcX/L8vwy+
8d96lBVrKh6atNwXoIolWjhcRwaegdfB6ff1MB7Nojdf109u5W4seprha6QiovZN
Pd2B61X1XQJ56cWpQG8xe13jMDzo6t3U6eTkKpLTzrL1TOsGAKAJW74PImXt/PK5
DwG3zSbaBlZROYoBmdUKdqzI91Q92GfDWcs0SzCSgqF3XB/m+sWq5sKgIX/1me2H
ivG0JGj791Op2PMbxZn9rfrpOYlpXe4Fh6trdpz7SvgjhYbNJ05mzVER3okoczVX
foz+mQz/5vw5PBYHs0CFZNZQEBundNJmUgBXt1hqMgNfKxP3g0iySuCraYswaDWB
1T/Sx1eiuXutViHiTZSrvoOi3lG0X4Hxs57N4Cdc7+5Cl+iHrHew7sTXkxHOw/uj
jMpEHU+BD952Og306xR5c4dcpP4PTEtPzyzBWxG54uAz9ugpXG56nNRXU7iqDVP3
fjVNuRx55UacXJe7h24eE5RXdpXVKn03iylXYnUzYzkU5rogGenAh/XowtF0Pjr3
Ekcp5ZoK/tCIa5mosdZ5S1I6eyIOQZ7wG01Y/v9bSRi3oRS+5uNPjbGZImz0Vr+A
WftzvpT+5yrmF+ppKpekNzYpDebSKJHdHnG6Iq37YJAiUdrLNytkK+WNSch1A1wK
SNcApkH8tH7Crv+g8xyxeYvSd5M2sDPXnMEoLUm0DIVItP8bO+uQJwOhBVxrzHPS
3uqqRIjQ93FUiI/MVzKeBKwZDzsw4eChk9j1aO9MRGSGzczl5BODsV/JjP8LKjqe
nhY6cH7K7tPllVkvnHbYWVBH6mlSlBJo+U2fugir/PLgsoFnj+hYYbSEalJ7JQH8
5VHLIC7R4zBBUpauI0/dvPd58/rfYptdvwp1bPLqzxPiqLI70q+vKBtqaXUsUOTf
e6DGxUij9Omrb1sGYmXW+Ri8/kyih5n8zNP3neLujnDGM6yQbSw9JFR9/5qhke3S
hWHVNnMxNPNOV/n+iPvrGRHw/r8ufMLkaxNMD3kZWVWYGl6hEIlmAAsbn8erHG6F
5irntC47QVffyHIzfw5DCrgmDkksgIMkBZAeUZ0Y68t7zygadwQlMYVEtRoUy1aw
2ox73CU4TX5M1bNedl6Oe1cK6PbPiox6WOgi4M9v9+rKJ4M5CDg8RDh1i4taqL1P
anUfDmKoXQgEs0nanXLlsrmMlcHzNtDKt5XRUl3xlI1K8y9uXTeAWlmyvbB6B3jL
6STtOJJ1ySWhxyVD80bM2BkyjldieDegm9JZzietQhPjOTy8Rvx7u+sYjp1rL1o7
LFSWE/RYojlAVu70FL/ZudhYYHgZCkDqtJ+f5D3YJLYvM3J1Dp2Pr34ZEn6fJZET
2sid7A1OY4GpJiMkDE+3WY4sk8WYZ3LiH2ymQ+AFl8Og5LW5PptcXEoJU7/SuAjh
rQ+V4FRkD5FnQVc4QgHg8lMBhqZ3RTTlre6RupSk2Aiyu0QFVNLhJDt5ky5625DG
4HLnL1dh40XCxXP0P40YwLqSv+zwLd5OgDmRDSrFgTgIqVpOgr2HIoymoR47hJhb
YozLCLiXX69x8EOCeCgNEQvR5o+wApKdaF7xNT0VrvsxFir/Qsl1axLaWUp1l2nw
R5dnlxcSXF/XhAoYdWgztvwT3LfaXP8XFPgiKg5WwnLRvT0yyUYDzxPhxRJTJPLP
Mu54Bfd/aIwBWfD0wk7CthnrF9fn6ucI5X8pHTiX1bDo9rQLwjVMFbKJE4inOCwJ
w/yWCF3xUxGJNifXxeoUjAN8b894pJDxubkD3KknhaqwH/LzXus1jf3OzKulYuiJ
UfGafPjWAB5FSUbGfZ0JldnIAiScvqgslU23YhR2KHli6kpWvRByZ6wHiqlLeXlr
k2OesLgcPcjzE1BHjqmFdCr9flg7IFzphfGTy4Gl2GwjwAXn4N/uUUJ6NmpmaYXU
5hLSRnaA05E0uO6Yu4dywriWkVgrRILNW6IRSG9m37xlRVv4MB48jD/6CQjcBoyh
23lxtQ1gAAByiymrCHCchgS9UGjApCha+RjANrCiJ0k+EJfgDQKq0v+fAf5V51To
ZGoCKMbStvMGIEpfdJRUIqu4kf7HDp4NcCtIfYeSe/+id2lEDufKy7DkzTuMO/Oa
9QIXTgoINT33zp9CEmwWPhQQz2enFi7PfeprBeUlngLt12GmWQ90pUPZv9lAxhEg
v6HFKXJofwLnfE3objY6unkmo7fJ1HEqN2QtpgqhEAvez79A4i92dNPPAkxtlKlz
bS3JhOxHNlXM2I7BRPpUDMqvUZsvcT66vWo5KTeYGMsVftSz3CRPc+GkYoAxJaB4
NG3Ston+0qP5GMETBGqy7UhChF3heZIvAg9GBWGBBnRzEilikQMrfZ3BK3XmseZu
elT9vT6kRmgvymLj7bvnIR8ozDOz903IoafLWcyl8c0KFrcdp3AMt/J6ih1cFlj2
+MWSD5PRHlfYM+1/O5PcBtgS56ktBKqiIW5Lws1F26Zq7ZiygCPoPknoeAVdg/ps
CpydV115ujynJVxI/FjLwqNOngsqEjFpofdr6NwqGh2Pquyt1suj2pHLY67mXuHV
nuxZlP3/wYwOxyFHm5weKMK1/rKQKOR0BNWcNaMorE3+0EIlOJnyOfRFEaSSLklk
H9oaACR5Reway+zh+wEESngOoVRM0QeUHrDmdE4ekHY6Mt95cb+0EquhpS1+jxG2
6Wl6EL9trDOI8CqH6Vinc0RnzZsM1Hd/v7xk03Gil31f0LCBwWX2ums2oW5aOhvC
iun53sk4ZOfxDzXM4OdSEUx40PBhfqbGL2E2pqa7wXLGhth6V7NQ1AJzK8cXSEii
WxC0apyjp0zcY36h6j3zb4nZHyo6nJlcJB70dlikBKZqfb3/CDc1uDat75OubDbp
mIsxIxUG/WlutByn1VUmR48XN9earDCHWb0S3kwLzRhLAQTjGe+6Agwj/x51uk7I
qwDQfCC3/PFUMxVs+y6iKGKQ7e0kea3nretPhFluK8BL/Vcm6T3+ccgQSEPKWBfF
6EoFNdGJ93rlL6vuq1jcid626MltyyD2xLTcRO5nbJXbqORVuFoQiS2tu6RuhRn6
+9bA/jTgL/70w7+ZeHsQff7BMc4Bt37eHUMHzja/WHos+0RhmYpSeN0P6yaFu2Ha
tOPXak2btkBvhWrM2FwCB1U6LeoGo8xPFSV1u9M09UGV+WX0iXK2XtyrUsyojPPi
Te64Th/aW9eUwGyNgmU1kTzSI5KjRAFsIrNloPZYN24scsokmxEMNUI4OeDsjmCO
4GR8RCq4v/KUTzDE8DRh6TbW6DwITW3qf0xXwLHPPCWyKZhM1Ai6c0AAmJQlyvCv
8kR6F4+7L5DQuSOTL6LMkcHRcm0P+TH22go6l7gGSp4WXxqEGUAqJw4vBmbLctYP
GgrVMD2107FKb3KkU/7IbED25QWrOEuuEPHWCOAPFaDxclG/rnIuwCSW6LD5+0P9
6fjvuh0WX1vvowo3tUAlcglydbAtik/X9GDDxrem9/+gumUrerGfFKj+zf/5Ioye
8r0ELPqY3l61uKBUszLVTrZ+lF6qv0WDSN46ecuvXIS5KErlyjVi0UGDqLdr444J
PCk9nvtwnkSFwco3TrglntCbgBjDyCovEz82hu1pl9Nd6c7oNHja5DWytNYx7hTi
JCRI9tpRzVDo8omhsqD9D5LHZFCNtXTLjhEcOqdr0dRBFBQQ68B/49AjEN9WJhZL
BdZkvlt9tVQDSknw1/2vscfU46/oV+8WqPRsEQpBogNInIQ3M1SBOkMADuvnC5oD
f1ioH4r2depSBKayIhGdhRLeXX1jAVpKViGPCEUsi6/9E2cAVzdwY8jMOWxzUWk7
PRdDfX3wVAF3UdZ+ckL+bqmJR2RIEbLPZBYkDAeC/x8l0j39c0pZB/ivRLdqSnif
ULCmQrJLjFHd17GkoSIkyMyodORyGmaWmqj3zF0Gr9G0oyeL6B8+76LDjnBm2G+Q
vRxVMBOMWa3AhXpjV72m75YZvUFPjUtybD6/GW9vkt4D73wkBZbYpqp3fRk2ha5o
/O0m42qyfQgEXEUoFrJE5TIXKbQSJHw+FqxMiCjunigfBS/eLnzmu9M5mFSgI37T
qYl1rWUr6vwZeIklXnr87YHK4HLzjV8XDP0eMnmj8idu32ymjrqB0VEjMs/h0LsZ
mcaAvaMK49TbT1oI1u1sgDssoRDX+CyUUUjzFQftNdCIR7ns6WoB3KdxL1Bhq3dU
zlmm/zfAjKyy/aGinD+ewGB25M+pFqLKhZgoIzHYHcj7bvkSb26S52bjYlFm3s+y
HEP+yS8masXtHxC3XP/aafu4261VyC3EMYUutcNEoh8iqPwY79GOYsBUdSXjYdqU
PM8GKbp4nGtzIFWL1Fkglmak30RbNXhF09N3httbNzjU3OC69L4YMPPNf20T5bUC
CBZB6kcDjwF/aouyTGTnEMYrNMvwSJQMZ7czeBz65wk5Hs01UsyFVcipSAehT0jp
gu5+hDlwL+cVzHq85B5IHMF0Oh8pdnQ4oo9yf75/OcHA2p9aBfL+F5DZmMLFXlBD
UqtntY3N7bZo/qWEWV941CfrgHtXq0UKCPOvTd/I3vljvKW/qDmlAkJWigSZeUIV
7LHwvmlVKY0d3+UlWsSVQT1wGMgypMfqEpEOT3J9pZ7ltG859rEaVuD1tf4L3qbr
DpDNOhKjGlAm4qxFhSQZuYoLXjTsaAqVQwsVB8RqfRcQ2TYCuLo6xuHEIZFJsN4l
u1A/5EDMgHPzMSDjlbPsVxeI8j3GuoXRYI+FqI78FQAcDMP7gy7ej4mdgoOHuXNh
GtkeWfrDajm5bXKVH8Cm+qZoE/KyrUKIJGgxPrZ2yvVGgdFl5Mksua/0BbJ68gL/
kx/Q0b3ghlzTyR/9Fo44EFXawYQapb7S6P9wBqgL8BtQoTccBSq9wih0StKTRJLF
6Hn3oYguLK+acAWCS/dMBV8fhQ+C4c8srF0HdWcXvpOd25Vq7veSyfRvL/pekFdH
nCbQ7+UfNxzl7L9rZNaHmYq9Gb5I1bC6SoSfKVwapvLcU7U/e1pTzdErzxIDPAZA
6pXBdm1U5lF7t6DcF2mJNUzVALXsNYntviRhZYVdcCw3YVfM/ftVzz7LrYImBDUz
PDqT0V8F3FzEkKMMmQTuIYN9HE+qIBIh2bZnL360X2ehzi0hL39OdYfSOVTRVrzQ
HIw888IcnU4Q/8pzHWqWfqKXKvt7WSLhsddA4+iPYtnUjln9jLNrG3961sk6KaUQ
FminQtpYROByZz6vFqKldLgdDZ5oLPV1buOivLA8Mr+uqO2ufRRs5pIvWLw5k0lM
yquGQU2fQwVu1bn65U7fxKuyn/WQ55Z+13RLec1c5SNK+N3WI6NPvUzBycUvAKsF
oWoMPTMFgwYOz1Fvc7vAIJ8Ia3nrFO1yO/4lwE/ljwPLjOw7CDrfHwrsJ1bjZ66l
A470IFlXgKE6lThknhId7X5IlB9BKD1865ufHa03vavK10iQlUB/exE58DCpm2qM
ZC7jN17T3WR6XZJrJeip3T5VtJyO1nT+OhpjF0r8bPn8lYv07+unFyq8KPox47sk
4bIewtMA7tsZPCWWMLut8+dbCK1zRWYlKiSVPGDmKEfVWCqMdmjnxItJSf3iEeUD
YeRhctr2bYQXRNCJfA1QC+/mdfISoW9O5w5sEd82cAERkne2obMJZJXCSG0OQTNM
qzN4mBxcn0GcLHcxygaTD6tfNnQFM+daBGuJWI5c8bgeMLb3u1NmXdT+gWnwPMal
ddFyVRB+TtbAQjIJxzPFF4KONv77P//1lZR4Th3+GF2PBstqFBLLQWn12J74EEQb
ZeNPRprF8SI4eTiRBJ+9Ip1HnYZcGjcGxHFrqv/x8/o0Nmrsw9dVxAZ1FqzJXr3B
qW8Y1/iyr7My8T7aJzNvoz+XO9Az4wQDmSuTsSBb0GVD5ZKXMZOnaywF5FL9aMDj
svO012BQm4WrBvq1T+bDbpQqCfQM0DbOuhGAA1hrz81IXJjSue+Fb396bkD4CS5w
UVKKttuJpaEHe8zFh8iHwyS1tcfk8vUzArWrbPXrpwQp+S5Pko3g2RjTSHCI38Mw
AnfnV8pImFXwXSJUB81mw3D8VgK3f6iuoplsfuly2XJgVgLZ+s2amuxwHVFsAcgA
jGEN3VOGGYCCf+uf0TnLNUt8IOxO8avgbpA1M5LlIhkGEIhfQzUSgz/DpOJkjNA8
KQmm2zVNckaVJyfKVkM9/ov27z5ewEzebQFOXXDQMnyOUogLrNNP/5pwEr+MgvxS
74PKF8HsYMVYmYjx6wxfFvb3OGtffzKGitK/YPjiVuoxnDD680adAkTO+YqG7Fgb
91fvNThdzLsk3ezX+wSx454S8KZwZGP6TS/dXj9KZ3+lQOsxF8G7zxnIV+9GNov5
SixCwMd+H+OqJDlq7qxNEy7hLMcRw78Ii10L5orjJyD8x5keHU+rKMT4iPguIp8b
1tudqtfxO/4ZjWaZWhirobGNZZ3FUTn1E06bHU/0NIVEWc6IDvQBfNHfhNRI7eja
FWg+pBgRcMnKvoT9tqDiEJAyjB5CTB1r97VflDfNWcZ7ap4s21QC8y1c7TJ86eCA
lVhu3KMm1MIyFaj6ts6tnmasCZRSqQjBQsQtTalmctIYQF0FGgWWW1hHjZBMh2S0
thUAFGQvoFMF4Dkl3kuUSZA02uF1s07GcWAkBEjFm7R7VZVQwrintVgLE0cQ5IEy
kD1ryU8nm0w2SLGQU9out61iSDtRWImtg45etG2VG2u15i9h3dYyj3DD74pZaP9F
1A065znlD8UDuP+NaB+O5nzl8GuqlFkTId6OLhGBb+soP47U0kl1IzuHaF0WXiks
fwSxkYD2KLL5/Tuynz5AuoIvdSIlTIArG1ITDRrwGyv/zgSJtqyXrjhWDavEnW0W
P6cSoqK2ga9WddyIdJK9BzX0WEO5Gk7TiIn/yugZB6NQEvC1QA/qOB5pb8joShSq
urPw2cXUsQXUvwvZULPAFdpHKksMi60t1hgO7J/QZnVJ6AFYFhL50fe5saXAWx3T
8t9NN6d9E8nSqM4LSshw2im8UpWMDGImaYp5mKEDJ3Qo2+hYpVrBzSb3HnAWgxjs
o0MOCVe8XsaBh/ZKTH2BUArKTGOdiiB+8bJQkxbUZKjCU0R03jS9Wk476XPXTmPU
vaZGG9aP9rXP5Yzz4+ktWV57N4zmj10LGG4FL1otosLpliwAMq6CDgKzcbHpi97u
pViNef+hCh2W4s4PgtExr+sCbZIuto4mlp0K5QsdWHV0kufh8EP7jP2XbRPVWNFI
6lFEHqUPSmM88imL1FDDNADZf4YSzOX0ThfJI0sBjR3QyKW7ZzTLCW0T1Zz9jy8i
CMliSiFLiUfLO/IFwjd7CPJDcwEHMI/znMYKYHhEpW04XIqJzNbXWi8LJphdgiQ2
QgQvEwoKLfjmqJe2+cc7opUYqLqCbM5SzXNHmW8gl2REU8ADsSEJ48BHomlBzLsT
AST4qPjA7HqhbxX/0SWOVyWBXiLTS7iTX75mic8CSQW9P3M2YJRTogptE67Nr+Yk
K8M/TcrXUWrtRjtuOw79ciJXRKCBFVXiuTx32yFzjkhRTSeruqfmRFdAYnX0AOOR
fS0zS3N2KzMM0pj/4fwe0Xh5Vpqhdrz2amsJJr9QFqjUgKIRPOxBFDqPW62W8/nN
agVjf+U265fR8C6M4VJLYKUTkgRMxbx4XMHGHWlCx5ItxCmdB8NgVOgW97+tGZj1
YBNSHL2DJR06wuVX7whM6DsWNOh0PThx1zL/DTq/AYhTkJAULU1H4v9+MmaMSYrw
dZWcAFwqPDXYwoBRC07iPvO7i4j7hWolYRvOp6nlpeIu98FxLewqLQh04Yyhy1Y4
MTlnYW+tH9VrbnHZ4nga5BJlihCxzxt4XRByF43oBupfN/Z6Ji1h+nOuazhHSFmI
ErYynM36TE1FBGjnMWu98JilWl8jLCR/DZncTvuMGGaadZVtq0cLEMvppmHzJkeF
VINyyfEStT9WhyCYbebuXXcscF6Tm/+Ajy6qs5cuCcx4PCHzrPoYgLcNDcCIVc6I
3yxB9EYejcqjznVaeW9MGFDGC8/LoeLmhQl/w7m0Nu4Rl0cPrF8Z2aJcqkMnABhu
GJLWC3qJk8z1drgh8TB2WBAxBECY4B2JreOuOpLnWomJv3wdE2V1ULiXF42JtqaE
/QGpBvpMI5sCuE+iZGvPpu6Cs6k3HQ+wQ5FrLgI8VMlIxFDSJMZplPI8VTyfX0LQ
fzdfhEzx/U2tsE93kfNzCEMDEE8USDQLaMtSKAvu2MRcQR9uk/7WKeVDzhDNWoZ8
tSsMfLiPdqqJUH2itycAT6RFWbiHZi539iwlKxxi2NU4T9/szEYz4zSJYLQ4oH/w
WGZb2vsc4L1EzNHRQimX88MkUv54DsbwghH5f41JxT4LVhHCSp9qsUY/LrDU/zD/
9VDlnEepjWVcHkrDJvq8kRkDduo5FrK1cFE3DbnCjwQBwQHDD7U7Mo3Mi3wDOn4D
pOOkVM71Ts2PhMAEQjaYeDrSGmD9vPP1kUR616LYQ0y3CL77GAQYN0IBqETizvEv
sdEImQTYNXoYZorf2wCy78SdNmc4u8RSVGogBsY2mU1rNCBB8hWY2p2+z4XnFPog
AMP2Xd1wxHhtbCBVNESqPmldQVrBOJ6D+reXev1cplg+vlO/3DzK7jKNplKx5Zg+
aqHctlh0GIckyGYbRinoVSskfxGbmZuXbR6jOEuUO3Ely+kKJwVi0o2jh3ARtVS6
EDrRS07tH65nj6Npr09l89gI78tH7hwKi6A/cnm7rKYJdhN4dF17foOCaibqqaGB
V4ShHbqMp3gWwbE090PRNA7ZtP9MIonaEaqSCUTIqbiTEZog70hvNjmYbTuk6NqG
qZDK11U5cQ0DVkA3JBGuKN+WOAG4lkeR54WLP0sQJMu32o2nHsQvn36pUMro0FfM
QR7uDDFDjg5aIcPvF30k7XnGAhFGS9Bx+N1o6TfyV7e4G13bth3c2XHswOACSiy9
YezAyNtyq/1Tq8HkFmNSNXaNVuKwgEugU+JhCC5e3/ZEjg9sgb0P0yLMKUdSk53y
vd8Em2dWNy/xtFuoeEA4qjSpDyqPMR1xFBGhKR+gP6y9UMNPTP188iIuGiDy3xSs
CmRpjK1iqAy91cioVqzr1ZUUiWZnhAhM65m41PKIE00DnleBjFaDPAzppvri/A5i
qCR/+KZNiSUaskCJM7Wcum7XKzx1E8SfGKeu448PA/MrL8YUFef6+NNSJIw5Co0E
IiqOMilmEOJAXSwvPEg8lGJs4QVRO7ntueK0g4nmz5UIGTkPrlxooPtecB6+F2bY
E46e4Tuwhinnh/OrBYO+bhlLGByvxaZplzs+EiQvkvcr+80BD1jVYb4XCVLURCsm
VWFrObtkqZfbtyzHhnwSTtGqNW0WtZpwCNCZVYNkuGE18FgVFGfiKQ38l/c0ezEQ
+RZT7m9BceP/MGB3Kv1KJSE1hJkZKdJQTjO9bPAaS7FPpiHV6Sf8fc1TF5i4rQD/
hjR7p2EJQUIufYVoiK3vC4ncR6B82I0Ay2DKlCA/oeAiEjN0Su8G2fBV6gTXJ+4J
rCib5HcFe9rWgeMrz3tlsJFsZtqYngiM5WQmjffzpY6GbPzyBZ7EunbNJMYqo7SQ
LWoF3+0MWkPK7K8lcrf+jNpDCVtDly/RtRTDi0w/y4pBOb7bUX4oC/0dqoR5b4I6
IsNaoRwz6oUzLPiy+Vz4fHnXKhrcbJsYPoJgQg+Wfp3Q9sNMw59luAhv7e5EpO9k
mv7S6bVx7BA86IZ+OrEAxzbPBNI4ZuBGLWTfXmgN+Q60exyAqDUizMMIN5pjxUoK
2RQJdKdqz7I37Th36ER76/gStjnoVwn/SmumgXx3MnB3FT7kelIuzUatnQOPS5w/
fW2Cucikdq/OPYd4GwJTxQXKXZe6L/LWzBkRQjWapE4uvPNF7zM7mnrYm66IPZJG
w56mH/GY0Zk0qM9cyTfAyLJVnnQHzfizXXkpPTHnquGbXYLmfrqggpLLxmcu+dkV
2/h9Z/jDSA/6OSJtmJx/gpWzDbm5fp80tqLE+QrCme5IMxZgIr5U5KYACJvkzePb
fLJOjiygaIVtGrszf5DslHbfTZj5yPLtB69c79EFMXmBOa391Nc2MX7GNPe+8Ku6
4smoPR3wMp4K0e8YxXFa5RcDdU/U5G3gFljQ8hhNB9IjsJm27yNlgMWIxbzkxBZO
wxaXWvbYs4J2HeuKnA2E83x0GarqrttWcffbNbtkN5M3BptNowq0GBy0eIYn7B7i
7NePw1PwkPjvX1Mzj3q0Qvbkgy479/joFy8CNe2i+4FuvAaarObeaKP3yurnBE9A
0xczgU0+O3E0MxrhSDz9lxQqkv/PW3j9qKnsYLpNy/VE7l24dCU4J5HzILKPnRwJ
UeRlZ37K+3jXiVh7DNjw2boHS/9SMIzkbWI1RVbgoTBX6gXm9Ls+Trb2NC9BtG2P
Xl81wjoYSQ3QEth7eFtp68m/MDCrwjOX1ejQAPBTEtzfDgwphUbIWpTZfRap74Av
52QRQjfK/Kqzw/oaFIeF5Hfkd9SvBgKpmyCHMW2VLMYo+AO+ryDg8WY8jXJC4XT4
BQ0h8s75SoWrTw9gdEEXcHmM0KJ/C0x0ExsGQ7vYgRIFoOMZ6cjc2vMr0drBPzu8
+YjL7s0Bhm+OddG2kWHrWIFXellbFgGFNyy32hH1u9f7m/JU+U42In3NHWe0VkuZ
VJ3uUqeKE1AB2+MFDU48wwYVuLJ3S7L6zallgBJ9heMati6P5S3xXu9strAcEgVz
9fLRgWVvEM8k9FytdT1Izb50IiOdVbKtmy5Xm6HqxiTeyBAAk5rLhvYGyoPrzPaT
WfLGj1cwyoU4ELoxoWp2JhuXfkppd/wWsiEzMJUbCdkB4KGkLiRyqpXsKkre0dGF
qVSpOM+YZ1b12PEVSesWKVunNmj3JjxMtJyoN+ZJxLlh/C5z/RICAnu3LmnzFsL+
QO+K09+3Zwm9Hlgu10a4dYMjWcbH2w4QEK8HFw/aCLjEDz/bUwwWY1LRHyo+Li4z
i4ifvjFwdBIuOmNA9qJcMi7BWeU8YbmiGlS0jimLMUSucrMN5beSACikpv+MIEdj
2upOKDcgQGRyWIub9c/fT6ryTIzCI+lBSXo+/LPbEuv4FuMqB8BCD4lf5vwLTWq1
GLZz8tssuIfOCdrI8wvTsIn6ZjnJnBBY3rx2Yx2g/rqHo9D0WxB+n//2vMWwjS8q
qm1zPoazvJmhf6E8LYWoz58xwap31YFO6sNAWziRxoHo3n/c9Mydlko4rG4n8SI4
FWiyRR6+RWYegcrVXjTuyQUyvSo3JjyJZf51Tjt9CweU1UL+RbuL6clOcUl4ekDQ
uq/9JORYYYNL6dHal035o6txXY1240BDEXzi+HkxVy4C9ZeJMPs9S4IcC/Y6VEFp
BE31of7D+NXUZ89zhB9BAKMF9hxPWbnxTZsCXOuhNmYxymJQNhZmTt827pEn/KPP
z3QMM+2fjtqNvr36wdPbNiaGIcpNNeAO+kxJIOJIq8SNAdurZYYUSCyYRy1M5KU7
yMvtR7Ihgyy8d7t9w0VeHkNgyIi4K3rtP36QvKeDEcpBIgwB8sVbtYhI7ne7SJl4
zbexoW/rQ6CRQXD92UHb66UongbsbEy2M/CmKBtct+ji6ZqHiHjEQZekoCJvOIHl
a4IZZMxzq+CVc6YEH3isD1lTfJX5Wh+xtMDcrxFgcnF9WnvmQedTZVXVpknEvg4p
bZzZRbUTmqfAT0QkH5hcL8FHeB4tlSXzoKqnM9JkAO07Bs5keHQZuWlz2lnqxOj/
1vLNCpq/D67y/c40vaBuqCkIYSnENDGh4Dc7qDcQ9NYv0+uXvaZFn6h8IUQVc/UJ
nQj2u3t0X6A6pP0sfVYjHBCFqPTpzZm1I81gLjGP/l/Kge3Zy7LnBrhGy3MvUcZi
A/879lXGa6+wKK3rrPDgC2GxeJLxW/TRDudhKjDnS3wSKoA+KFQNRuYh7hXLV2Fb
bs9uE+2mvu/T2LqLCkuJkzKYclirczworfMJIut+OMwlqFbok3mOCyVVDX2ByFnJ
Xo+L6xPUF5qAvjhF5qP+Kw4g6gpycPyCQ7W32qBHNFVC2eXk30fPUOsp7Ta1UtLs
xsOQ37Ho9CThxlYStNRqF/dMFETCQHnSlRHq+Wxsumt7mR0TozQJNSFu2AFu0dzk
9pwjcfNrp7ZUQA9Tz+yBj4jp1f0hECuQNUYAUNtNZRTgTgGmmZCioBTjAHx1k+AO
a73s/hXTQ0qTaA4CS6RW2cbQ/PuYdie+Pcdv8RNbDShvRY9mtM8FISyGIFVFlna5
7IJa3oFtaoPpRM7pV3CqW9pxVSAUZRpGyf6sAbYM6RXemHB6GZHzZnMCZ0VgVGE5
2jEqTUryXRlMpRPkVTVE8ZfWFzuVhN3YVfMy4lOBet+lR1ugFcNyMwJooAJY5Cbj
7yfW//S2zJKboBZs2dOD/0+UvHgjkr/BI2p9BiXGQ6bRlB9YkMtjXJkDN3EzSkSa
mGdGlLv7QFJw3jp/WVzjQSrVdgZ58b1eDihd/Nbt+DCPDLVBWB7wOsMefVTmy4tx
1VdaM1t/loL1p2z0QwIMVVdF0d1o3iB32pXQVkMgKqn6yWRuvFlMva5MhvEDUQUd
4U15NYq1cqXWxREgm8M8OUUB8KQQFCvaI3lYGEry/l2FokjGGiFWtqwmADYxD3wQ
6sVB7eFbtsDDKHCiYOL7BJK2bVxtdS06iTXpQuCmj2lx+p04405J4v7tXBznP/jQ
thH4Qg4mf4oo47tTg7hmOBcdeFmZDB7I/cQQmVoVNkG1SqP9Yq9g3n+WzUfUERS8
GIMKqoPDP1BgdiNrVKlgc45SrrW1Tndk2OwMHhtgid3TpEA53Hx1JXIoD1BYQzaD
xK1ilq5R9sFFAXmPl7U1repm3elEK/J9ALserzVfDP0kjJw1M+ol47Va6up/a9Pe
0LTCEyL8YVnLJ7h1q9JSeusfZxlSXFFvHPSvKIKmHPE1m1uNFubxPOJ3f8G07W/A
Xdrq2h+6QCff0xg+eLZqmHzjzBGznuvpOh+3Dip6cL0mXymCB5bSWauLTjxtWP1y
7rzGd0OcT3cjrQP43CWvT07kMo2Pjp52xYBN14KaEYhZLBP6BuhZdTIf/ofpZ9Dp
T4ERFapCoLAO9zjY4XzLzu8TT31A22foE1VxAJWhr3miuD1WeOYOMB1ceE5zyt4q
5ls0bstUoMReQyKbXLw4HKDKBzYpNSRpjidV3oMcTIxQNRYHdpWPAL13sBPlFuKQ
b5quyULK4RMSagzVDKAV/zj9D4Xtvw1DLF3MpasIh6a+AJdYlbwxI1CRFA964MQM
xQOenKwx1BWBAOCgsLavGmqgiOvgRnjK/0ZCw0QJ/jYl7JQe+Uluaa1gdtH3fBU2
W5zw7Mu5IumynUTkRQeilQ2FRAxDUVItbxkPulikryoZ/bdFnnzF7R67OBcexxno
Zv2TlfCJomurCfE0keuT/Zm6GfT85XCpkJvtGgAJiGpkSc9OlgjTdW63I+wRAVDR
xqoWI1O3/d7DeVUg0N50ryOXi+PQw5IMgJzikmfVzxWMxLLpU9u2MxeeRFbBMZZg
24kD4eHu4j744EnLolVBvbZ1Zfc8QIyvM95/+NDxCThSkZb4Mce2DEdeXCtsp0Kr
9Ek6zsG2nFpMHsP6UDKfWdMmwMHBqrBA5dDvQprh5tLYbR5Dcme7CUIcJZvIrAuY
POU3QTTJRwIMjghMkBjWXVzeKQAHuEonDu5MY4hL0kJPeCsy+FHj7rUmIN3yfB8F
mKXMtGHpsGsCCerdpjt+pQpT8xzAXldcBpZr5pPBNgmVWSu0x3z9OBpLKv/ihnd6
sMTCcE3z7dFG8dl5JBuEJllF9rFkBIia68jkshg3dK+iTtSbo773Ni+ov+9LHhxc
qkCiOIoQOSe52ZD1mbvwG0clqYWrdI/znj4jFfonp+PrRF6ieALB3xVDTPXnTUiG
lQGgEb27e1Xp8Egxvw9zy6V17EGQ9Otmgp6CDcgYyIkqdrS7WR4CIF4GskkIEcxA
mlnvjmspDGAXR9qg4ZqvLBVlU7vgNKCTvB1tpkOCMKK4Bl2r0kzTgtegdm9wnQiN
E+BX/SV5X6uBZBbhUmTYCFtUng5fEEZ1IEnHrK1ZPy1AsC+PQfQtQHdwL1+hVt/Z
rx1EtLu7lLJQFXCvVVbX3sHBHPUWLWU/W2yAV4qZwCujVVQq0G4pHCodInNj5YD6
nHmRovihAenvL8aSXerBbEwudXUQXwbcb5o/nMGJZNS83P16kwe2jRyouKSST3Zy
h2JHETKB079+k5JPxFXNhd4c9edRe2660XaoqNWCodzjn92Xrgp64s4Di7O21/g6
Kx6nFRnaQtb2QGak7tBLme8yJg7jHH2zoeXJDwIjG7BE1qSa84ITeZDHUFAGfcW8
mVfU+sjnpXLH7x1rhF79qDdp6PXeonCCI/02EIIcPAUIlsluDMB1T1AWmdiZu9uI
v6lVcFXOTwLDJG9/PnkxBAVpEWCMkWzef6L+wrEqwOrGQiT0f/x8fvdQEKhYSrfz
MOsNf8cwfVwEWQ/I58Fo4nkvFbGwtCYdqD9yHoPpGcFbZ35cE6BPGWxEQwaW+GQN
/sNoufxTIpv/5+MYlFeCbhavCr+HjmygeX4O2lFxb6UgJ/nzPbElgiBdUDftIqAi
eu2OFfXGw4aOKNUfUnEEpkehCabworEKCoypKFW/bnBhSmgqZTSAmUcMvFYbwkIx
9SSe0YGgO7aHaFBEl9xgTxRvLexApUJkpDnBvHROnQnFXQxx9TzVO6XwwZSPxt0O
vjlKmx0B3JAPgOtRgLZjz4NcLX2gXQpOkj1Kwm6vEvo3we14WdTdtqGzatDHDgwo
UlI0FAYSbldoXGcIzVfSNPXxb/STnCowEPiw8EE3rf8f+3LqH12q3YkF0VwO3sV0
imT230aemaZd+hDGKDlO3EWXA644Vi+kRoZnrLzNHEynb5YvYERtlVDHpeHuUezn
2cvc7ut02jpq3OJNAJps3pn5h1du5hajuHBn6pZTBPOXr3U9vgJqtqVnFeNxBVZU
wlEKQHMOZAwHdIlZJ+xXb1Qc9lFoLsxqfYe+rQ6OWqC0PV8nJKtvHcd9NxALJJeS
zAbg4bzt9ELfDsQmY6mRpgM6XalgqItgQKoA1v+vCN24rMWDs3DhCdIn5F6ZxcUA
33tlGH3PWIhYmcEKDRa9vWr6Fahv4qefuYTfq5XGYCOflsGrYJ25sSjQYEnSAWgZ
1G7j6GUJHGn2VdnRYUQVqfB28CsoFsXuvJWfqyxNQj2oXwqm5HU7O8lTVQbyjLZF
M5McxO2cbNbRir8aV8SMNkO88qF0moc4UrcwfFS6pYIA3MCe/cYZPza+XtEP1cev
1VxAD4vhPjSkZTCrcLX7cDMhjsCbW4iDlYVzdxV72RcNMR3vw0hrrbGIXkDUlhY7
FU4IL/qGmtqwQnGKXSv1ywgxdqOHV2/9ZlQKpczpBd9KmCSGZWEHCv6dYM06gcRH
GdAXrSmQ6K5fxYTxPNCraVW/tzFXApKhmpISArPKlEskQq8M2Kcq3SVzpgS64STr
CG4MJXYIJ8L30cCVCkKt57LT3GHBHMA2db9r62h2uukYbgjQRcc4V7mP96+yHA5m
VeOvlao72sA/tHV16HhMrsoaJDbJbGGHf1wqQiHNrb2BJuYfoR9jSk88j753AaYa
kl8bzlV4QsLxITX2bz/9uCvAMMN6fTRRpMcX98iFffWuWAvCtj3zClz80zXMwKJJ
nQmkVz+Zgq5zBrXu+ABbfc3kp37GJMIl1ktphq0CPKEoKQR8f2s4gcdiTgFtzvHw
SpbValAaiHHXgpReyMy4B0mcv1mKWTZuau6hylaLIq/7wfcLmF9bn+fsc8IvEVEB
Z+koS4ycgs3fPjYX1nETfxkkoB/aG0LZwRM2m+rW+kh2f3c3qEYWXXrE+vrBOq3a
MhGF66+OKe2lgljTYdZWIcJlBQLV59hrBSThJ/vbjPpRVaS1AcYbTytMLMMzQ7jI
iHGXloEBKqn5J/+tAR4SGZuQRGtp5yn6omnc7uzD+BSjlD46OnUlMGd5i65RhtE+
62xJHoun0M+PdxWXeHQu1Zs+l2QQzzfMZYN02ik6R+PYjwqJaz3YT1UCPa1uHDjZ
TTfmXffLi46Y+sKv9hXhz5pMC0p6onqYNVBjPHF2X1VZsBzmASgowfas1LqE3doY
YyAa7YxwzyZzowwe936o/5uQJNBXgPdOR8SrvSMCNKKa/PuO2ReUgI+XAgDzanhs
EjQsh0zwXBY9zwjidoemtgI+fgchKHZZ7CBP0xIhnMNXKo5ld4OASK70QT+Y/Qwb
7tGw1lgZnoYSA9Iksx2GlKx5aQrc9C/u6xqKv+yd7TdF/znYWmj8d0+PKDEqEII5
Bh2n6xnMMieNk9T9FJ1p4SDVQLnGiogemc6qSyR6B9PkCB0fYMIdaPTmKe3cwE/C
70JePwCciD/hFN0puE5ucDgcVLd8TXLfML+82yt2uP/BxsJcYcykuJMsR6ISidMr
CtJGjXlfGvZimoyHjiIGDGnWNF0WW47JuB7ooOh5anMQmafsiL6TOJ7okKnM3L+l
rZ7iPW3Ij/dXZdMeOJ2PPJQPC+jyc9sqiS9LXGAn9vk8P33uB5iqIdldIekGmWLn
xthbqwzVeHuS+sXpw+CM+XiLgJD3f8ialHoWpEVjfajKch6DUe/L3PtaaeH1WXRz
D+pOuE6ImgqXLFcK1UlpLpMCErFsauCDQHhZwi0Rk7Vpy5dMMrk5Y6eRMc6jp3ia
1r5RQnkdyZNjZ0JJDCOJKLPhSxbGJ3gvA8dNlytGwUGbY0GOrGo1hQnQTnoPeqBz
k6dEz7k96UWzZXzEO4Ge6fqO7doHGs33SRkMDul7RvYovYXUNY45XI2fwxgDIzZy
C+AqAI2hNanLidYCnWwKlfjS56yCU0O8///ZYvQ4u94Ed6/7547CdUw7EEMfjHG+
9vX9O6JZ0eufO2hOD7VlGRAD57mpcp4IGRJiF3J8MtaVLrCl29A8aRLCa8FYBy1y
2tFJswqkP/XkMw2g2oHEOG0D/sgCcu54bYmJBo1N2+Ov1GTnvR//FZ87JmSujkdA
wVUO+eO22IxtOkSI0r2IL9GoAjfqB5/usswyL2UC3XkP0bYeovYfhESnoBWETU4k
XV2TdAlYdvkHVdFHDmpru+61ZxuyEreaK96z4B8I34+m3T3V5fkRTHkSBTAfGTXj
3XKFeVJ7QQYxbpS9xU9kj81TFPIVUUlgbzo5nSuC/CP0sH+I+w0qJHCqemMqfL/E
cxT05nnvWxqQJVqeLbjo8FLKziPwjYjYTgTdNZtCealGG1Zcu6X6AbKkP3jmrovn
I7rrXFGS3rUwuSx/TcBIc86dpGvmtQPC+yzgHWfISmeBUc0fGUARTFdY8hJlYg77
v9sL31eQaY7RFx3qStliRLYcS5KlNGVR4tc4hEsRb//FVM0uRzs1X4nvASozSPGN
rUSgTRM8kcxnRFYpVpjMbBz0bD5hYP/ty+mpdmWcNJSD3Pu2/vdqEslZsVNsx1FO
NKZtkH5zd1wcs9e+tqJerBv4kvpxCbzKcKUtpugZvaiNODOnr1KD6+XxYXMvwG2K
kKxRurqvxwyq/g3NqRGYC8ATZmkFTYO2DSZ68DpM9I+L9bXeoZcWZyjmDICFBWf2
AR92zvuJXF0MLt/asBAH55zsg3IbX1pR09Apv2G3E9U7lKQb01Uy11s/kutf3877
CPId2H6llPPr79FrSa+OOiBP7gUkl0XOq1dnZLrLxnQRXhHzq09Tgc7Grtn86zVd
vvpkYGKmEApdclZiX0pamq7DD1I1mgxbIFucqmRN5CGfBCQHnxEasPkByPVvn0R0
dqZ6N2sm7zDTgXr/HqTVIPGTuKJyMMK0K04Pi2CoXg0p7+vjxJHl4pxKBng5UXCL
QwJMPfQd54nxr6+EIyOH0QJL7guFSdaBUI98MDluKx0o1rfLZiACee2ZF/Ed+0js
mo/ZoeW1HpGNrC+aECw2RCwPrG4GIln++jQxqyyu8BQcG5BBWXx8wBkLymUDiU1G
Z77ZqZXgszR5um1Fet50g/qImOmFD/+RcO1U3E7QHpg8aNJksBFHlemdSrt0Rsmq
rZ45Iu5GRx9RLVJQsIF/F6cMa44mBAvYrgxOkr1vDvXmafsc2R2Sx6Bp25ISGHCx
1c9+nuedCn2ANB5dAT0ud+C+bAhyA4gI+6ChmRK2lygVCrmLxnH+pkOLHwUEOeas
LVMF9Kqd9oZFUUDt6pIRucKsV6YAaJIaIDDhPYJcnIrxOidyLF/RYOmTPLIy1fiJ
kSp57MdwGGIUD5C8+kmUxYQ4wsHk1DJs4QLL87k1DnhM/Q4sL7q8tAfW2mgsL55c
2TEG5zD8BydmKdHtX2VLFvIn8+A/b+r91hWdIlkWYcUaCrbGFYJ74ghdr/1Ub9k7
jYZO/ua+NmmRIkJdFRIZrbj1rmOcwoCTfdKiwJVNgw6pNhwgJPR+wtjBMgDEyJ/2
/YEWH3cxuZ3OjiTwE+phuKngcW4R6nzFZXat5w6q2IjfTSLFMhCQoO9318D9Eioa
09Rbu+t5bUEt8FuwidogB/oQDdUOjU2vVSddGA8Ql9nl3fRmi8FtK/G19VERIEWv
U0fvy+xIdNcwBaLJ198Zy98J+qvVb8uvsfvNBFGoA1kQ/8P4CRwFAUkAFcyY/ron
9lKygwfVxsyngJcQS+30Mmv+TN3UUlXN/XR98EoIunve+Kxfs7Rj4oZe5lU0StHM
YHThT4H1msn3z2DUqwmOUthlIbok7UxTaiugZLC3Sw5yizrB9JW3/mNOKoi2aeOi
OwOpDCiqz5rC8xxv6gYwelXDkLLgPuwa8z3fmgCxUAVc82Orq1aiS+3dU8NLS9fh
cLKW/EOQ5d8cb3JIQvUIQAfzzLKPWt58x6j4iyFQ7dX24i42T1GaQJw2jewHIayN
mhK6kRuP2U438eMJ+9N804kCOe1Lsxoc6x8DlVFHBZ4YbZORZlsGd/zQS2m79GQc
qYmyk53742W5e9rINtYUMxdMGBbQSI/nbsnrD8V541E54zGyruf8MzSC2I7w+MUy
fuCDDI9r8QXginQzt6Qzr2tMCA1irah0sZOnIS178FBKFhHg39P35g+zbyPGQxWY
dhPXNlQbzq3y7CXp2lLmkIOblsGxneYTGMptPB6yF9etV2SOihnLNqDyGkNB0NTv
F73pqbPDCFBSw2EwMQa9DKzSJdMePtTS7kLWOPjHIGVkpZbeaVWHwCXz0fIybive
ZC2Hp0MYODOP2BvWKk4cMsj++kP1FQJh5NS1xJ2qgUfahOHqgr5NGO8GCc1Y27vc
Q4HCmyAlHgHtY7DFHYdCZgIcGEC6guEbenaTKz4jyH762z03KLQIAxsZU9eo0IFj
JmxLIuXeZtErBMOtbsC7C6u2xDeKDNtDhOFRxFrz0RZIJ7DwdsmlLkH4zHUASNDg
AfiH5hdpHCTvDY3djr3C+CgE5iRIA4JtxOcA08joiW9B1jluOl2+48Y+7xHnMxxV
vYJVl28Ob/3PEyWwZhgy0hsTZzOOCvpXYkS6+NkjvKcVY+ug5Tqey6v/Z0t0tNoy
F+SF+bRKH+yUZUgXZPL6SPHZOxB5a/HNhNM5FuAE4DTHMVsVzCGOEVT+F/i11Z4N
6U4K7r9NDapfyaxZpxj08zYJzwHA/kNvaEPzIcWFTGfE4abkeo5NCYyh+Ih6NpzL
nADEXiDOjZDMLpFd5AdQA8jcJrj9adzJbxmKjARoiJ2/Ld6g9lPWwO3eglR3ZBc5
7cxNUZHpqDyNMxKsXdTkTejk7P5zeqjQwz35VFQ0BriOr+Z1Tc4/vvR1RzonH9mZ
A5/lL3s6FG+hlhw4uKhvHgPeT+n4aPOGvfPf8yR9WIl/ik7lbag5MPE9cCL5TIVR
cGLTPWwLDHilgBZY57sUKru9JSh3UTpduhbF5SYoyAFLUBj1PhjK2DaX5Tk7PL7y
El6bqUd8YHJbhngZgXFIUAux8p/gDa/UM7fLKUeJGFsRb6WfmeTZmfHF0t1fLSgF
Vdgw2dkocs/jJeXq/JEU0+9YNi+g9+W/MeStD9iPmMCh+O9dF69jI1U4N8wLYg/Q
JoiuCokHS5EXDOiTmMRCzvb0VDOe30lT6SYoK32zWn/5HXRTrd289++xWEqo5Nfa
cth896kI6JInABiRBKSnHkQ/BaX4ODP3xekxYPNb4rLKt/+7GVPUuvg6J8RqezDx
jal62DnG2t5S1L4JQqHzdIiVwFJQNXOpbr5s5Ers2YuiEWG0UOXODH9zdTQFrodd
QTWuOr50w/7WaRQDy3KoEla/wpZ7ZTlHTavViZ/UOPS7Meko2I+k61TUUjVtdU9C
EDEeBZwNTRcbh6boF0JnazOgR1cJY7ZVlbF5WovSKMTE6jMdk7HPW2+vq61QUxno
zZ/pNdHf9WvpqWNHI2OcZ+jJeK6RS1NZigYpReJSFcvmZTMTGRjPJpwA8gmp38zq
unEJU4jhcDai8fWPgIZvQF4+jgdGyUgeIBciCHE91qZYlzlNnGDXviUrukNn7rFr
z4NJhAPBRbOBl6fM5/HIT16pobHptWjKdFh5Zfn25ks1cwqqtS8RZJ44tQ4KUKww
Gk0uAEYchcAqQVgGGGGUBgo4+fYUx3rKqY5WjDZn4oKdbI9lYblXXlcbgglzcC8W
1cXNIXH1RdMLOui6p6ZopKKRCy6A/IXWay28OmZxTpIuWuZtC15GMIKm/x9x/1SH
EZLRM/G3LE1ODlQFcoKxHGI6wXhHBElvLrtOPmTR0h6OSzigCDHngrN9wtMXiu3Q
MB2guvucWe84an35biU5GP8WdI0vk6OjJcXto30xasgInzz/0aPoK39z8ducr17P
+ttmTlYA9lbv8nLTdyFHMqha2phIQHJpyjMzC88B3iqEaakzrcHnQPzOUfYZLf/u
WkbeWqv2bBxfdAbUGNDV9FqFPJr91OpytjqpmtEmUpXzuwOSfw+/983Ga5hhrNM8
o9uwwWPjtN1EzfMr0HU8EUQlluvzKcyuWgXj0tk1baL9u9ufP/rxG1Q8lAdBJrMG
FyZtVXU1HnIEaVzLf0QHKU9husnHne7JqW/SHfNPBARa98KwrRiswKIdmDphEmBi
mLYOESl1s55nt19jgTC0LtmMQiDxynO+6qz3c4GzyOHttqVlR0ISd88STUizGQTi
CCQ7uRaVUw4RW7pMNcICn4VhjZtJih63JsCmeB7M8dP/YIsnOxNgSnfWrkZMPcQs
enerpGlc3+ylA5+c7uqJn1ciiw/uhJ+OsAQXTREFbMjpbnJlH8WyhjNc4Tu6ZJvj
ivCOjbWLemzixOTnQ/GK/uFiBH9C2XO/g7W1hncXJNfY6dmnJCmgIjSBkF7/Cuwa
IFn2nRel3xkbAo9XL0P7/XD+r939SKANR1xgH7csXTBz/Ww05CT4601bT1oFZs2L
JZSTy/FApiEk8XB7biVTOmK3le1xSOr3RXuAmIwE+tfdWz7ZBPt4N++3s9X32RAc
bd3Ux9aUyoOHLs/3QUl98OvOVHGT1j35e+91EDPnyV1xTVMlya14pdJQTUHOYVli
uUxpMglH6mRCyhkgzmwgOzvEbdFv6G6o0FtMRDkFSrnBMM8J9Sag8Ww6nouZplHD
wEEaaAJSzQSCGH5bz+MKyhZmPZgsVD2y0+o1J2Vu/+QPLHxpcVX3VYMPPSJysTCc
xqJk4vzfFqipq84FvXx/G6Jb0O8q4ahl30OpNLfls8nQSOPAAzUF++C33WbRzMrn
QzbvB4wgLI/rULVtZX6q0WHIMlEUU1fEiG6NCdl6gn/K4d00dC0t6CYfG/KwNnFI
U8J+feXkFS0g5SMpFRklBBS6nQRxDMtu0GNt81TyXm6RUkeSLtzGC8LWmM/qHKEw
5EptDoWsGJr3u80ffzgviKls09DU8KHyiniVIVpwuzE5s/zYKOPF+K1YPTkOEFrZ
SX4FiyV9qVS7ol9FQdxJFFQF9U0nUxK3L2rS6ZCNcwvJrdIa/qkAiSl4QXIgeywq
TERxWWEpOwMen+JqW8AoDm5f55tU+A16Yk3LtOkcpvXdx747rxPkq/NxapPYTsxb
WnmHPU63ujlglGslL0d29RK0G3WQK2tmPHkotGtOiHZJoUP6qL01608e3BigDAbL
YZNUPlykKTUWBx9lkh1T9jvYk/g39F6f6zjXD67NdwdoRpIkAyic76tNyCyn4KQ0
5ckF8TKw+0jfj1TEMM27Yf4a1xO1wBh/aPzS2U4cWaSKylx4I51I9/Rq63Ywo/GT
j5jhIK6plQfPtNLPXF/IgxUkT482NSOvDuTGgniTswmglawS8Ugl9sz9Rf3GjhCW
77k9TY/usKzr1fkC7qLRp/2q6RKpAtmpzWVh1Sij33sX01akXnWl5DaZVfTR3xy6
zBmaQpTzYzwcMQvTtdEAXZYk1IyWfC66iGnfCb1sSoBja7grMxjvZH3W7Q6Y4ReI
/9Ld1mFTpmwd6tGWRDWbk6gn2ApfzAR0lN4siO6mCRZsjNVXapujbnCA0G3BMthd
5smYyTkM9XTmgIWd2cIOD4M0NMskdnhdzx7r8oOQRuXZ9A0SH8JirCLDiXgIyUtr
X6VRRbw/hXoanMOGX4Fb6ty9CQHwe+nQXkefIB2At//1GrdIZV7msCvxMimveg/a
cQteG2SGQvOY+P4LJAkNPLqtMaFKNxAK8p+WbD+U/QRkgZneEYbbGfyXiycVvwdD
xZV3J857GejJB1fursUqJfXXHGj7VUSJvg5vhK/yFsPUgy47dYcKCrKitz+jR2qs
mIBfSLxN2uRqrs/FNXfiFkO4GW5l6j4drdaf0jChFXt+3aviCQmyf+tSmYC/paTi
hxYXSsj8SYWZ2ESs2ZIW0ZAxADXjdbjYW6JYFNzih/GqEZFfvB74p9pWiXinejqy
fylZCVY5tHxMaiMGH5Qa0JRfi1zDmzinY5018Oj2ydVrhiStOLrl1u4bx1HtTwgX
fXlT+B1X6B7uWRaduoel96SfrFuwFOj0LbSHrQ07Y5Uj9N1YQUXmpwic0gqdHFFE
u8s6wOJU230O44iNEVJ5ayv8RC4WMPj18YGNH+5SocB2UF1sxOzr01T3jzut71ob
poTYEw3eKO+xSXeoqPyG3N4X0geh9rjKcrGLIRnPWO49AwrcSAgHgspcMAzhI8ah
B2inOjiM5FTz5SvTF4FS9uBzZc88karVd9ZvA7lRWAkdZ2QTkne4NqAAh7qWMaMF
GGDEnIJw2yn8FVO14GtXWbpZyhmTEuY6vqwpPEu7g7ReqxnYpGeMlONQFFBgzhrl
LOS+hq8ksSGM7R66CeEZv7B4kSs0nhis+lGwlns2odigT3Lt8n2GIO00sSNo5eyz
IBRRhKx7d6Dl1MxtEoa8rUJjY7YHD1uwxobSpI+5+3cFxk0HzADVmYOD+N2qQ18u
US1/TYlsbYi4ZN1S9AAFU8JUWBgaLywU2Xqp8JvqTt508qJk25KUfKFY8+8lJUIC
lTUUvcWWRi3BMs4hM/SqdmDtIw+BrruS7VKdQb9BcG4tklexyhHvGxt+A7CQDiix
FdpxzZScXyA79sD3btXVPX7Jl90bScSQcdjtCjcKGyy3gGd64qag6GgQk4KDJr65
/+OckOYxd5uRNa/Ue4mTLyRfwDB3YTcq5lnmelOBgPjdxmkFxJDQ6vXsfolpIBVa
Zm5Mqh01tiCMKpKcAVpjH/57hJLrYx5seolVv7eE3HDJ70nvNkWKT+A5Q9thsBkw
QOuIS//80T4//+JgXBeneotc7TOfCsxv20UtofjpuafIQmOIlC0CB2X23I4m165W
j9FwOmFFvAEB76LVUS5TrDzU+QT4nVxFmyKX1B0olHgvCUIZaJkLP2gYMqsnJ2QC
TbczysR3cqAX6ATIwcOf6wWGoIT72faaJtedaO1dFH5EzeedJE+AJ8ScHRCy7Yzd
Yuu0SAHdxe2Hq5tlaeB536OULU98tXQDgfLIUI3d6y99IKO0rDBo6LfT3Y/Wx+/g
0ZGMuKPuymlCJSqDJEBuiFLK2R6hZdOsWco/89Q2+bIlmrrZf+qXkh5iX/DQ45xo
siAhTK3WFeh6l2vqUSg+X+Knr2UZQaXiXtF7Ob8VhY3APzhbLtY7MuyHbLs5GcYp
rjXQaG88U5XcnbzWbi/pcg03LIiY9vkWcfN4xYuf4Oc5Xs/J5LgzB+HCsbO2TIel
nURmUhJ1R6gZ9CHzModxfPuIMY7P2exEVj039ZKte0SJL3lax315JEP5RRq6u1Uy
3npWIcgYdGqSydBa1p462A75Bn0C721zitpJyzlO7f80BVSrGIeFn+autLeF4UHO
jlrLkgs+YzJsjk9Q7SWTTAbkkdI+5Kmm2QdFuKmAAPh+7xQQYFPKiUs8+Hhy1DZL
SAvxOiU/4w2bDhr7Bp/M/ieuFEkJrsw8v7Dr9D8kwG/Y4FyzJZ78XJBSa+SqEXVL
SY016cRT0HXiT87/KXs6gunyyFXHV6JM5o0n5DiLvUnWqUW7vGa6/Jul/cRUZP6c
0LkWufCr6Z/S0SHfYzLEAZibOAOMUzXMmYgZc64pUGDi8g4H9fymphCv//ufrQoA
NyI4tmvRiiOLZEHHnc6RzYag8G+Ff2xZ9vqQ2VQQFO29WmJmC8myfMNgLpSRcNnL
jSBDrPdqEWo9TVGJmYaZtamTHcuwwImZ1/Ek+YnbXNGXiwAYlmV2tc4bLKYwWrho
n8QH+35I4CXlcFdGS9aFS/rtnJe52IXAMvjTrAZnZvklAQmEHDLmeRt47bK8rWiA
xpaOxzS6SK3AY5BINd7vzwJnsYfJtMuEyu5ryo5S5Y0Io2/rhNhlylS+Ru5PQeou
Edxo1PwDmNvubXircio8V2sHs6NPVijwvHtvkIRj9dd0yPIEoIVWx20B/DRIxxcn
sLLG5Lquorx36l0O7Te07dTcOdzN2HF5oA+/vmgjzlGY9DqAumjCD4vmTHqs5Ibo
4eSfCvziNrgTtjrLCT65Oi3WgstWyUgDgTvnu0EKC8bLU0ki/e/iKM5jPtZC/s7W
RDwXLuIKDeVRezpkBBokZ99E5I+BGPKvX7aSDVNtfYkR2yEBQq0u0nPcwM8sDcXG
LYZNZmXRsgAJkrapQYH8/Zbkcm2WedmCyz7cc6nhlk9j6hlOmJL6KaP/HF8s7Fdx
upzDCGoDOuplaXY5LQ+AbDDALvxC1xDi6Ene6XUs53+rH1twGt6t9OpGUBQUCPJh
hroENeoPins9cpcr4RrUoZOIh4mdtp3zPh4R41CQMpopRs6+6dZujOIMQ2Zj1moU
VxJIaGJ93ZroCo/Ba0SoXCwL7MnclbAxkSH/+kVv7E7vSfnYmGJqlhR8gAi9jjcr
iVo2StkJkxXZ2g4hz1tZchLIwLTdWJkNu+eMTHgkhiFE9QrApKYkNmoCT3batM/M
UIUgbybjeY+OFfSfPz+qAJ4p5j3x4RpWZT6IMsLhV1oBY7h4XJLthEq4qYbS7lAL
4RGNJrRt1JBVx1g52SGeG8XhbzSHect8uf3j7jPgBtN5J9Jpy5U4mXt8khLdUShi
sisVwksoq35qr21utIh2A2Y25vjfBh5ezqvNCTx8CjKgTqzgPLjde7WrFfojvm5x
URkHfnKb/hpiZMEbaD5OXea9sIcFuwUm31KFFD6sXppO/6HsI80I2jR3R2FsswcE
KgC6l45XxoZh6PZSpGGG6IAX0WJ47xwdMrZi7RtY9f5Zkhl+KZS3JPGOfgaQUU1h
G8hqlKvGP02JvNjiGQPY/7yK1eHmeC6MhQUOlJpmLd2yGJhUGu4nUHmFpFpBmgr0
tRj0SI1cgsXUlQ478oLg9EHzijE6zF4eQjtzgpp57vBv33Ahm4Av8LR31xkNiln+
cB4f6zBhNO+8/7vJL+9aKkTWldbcn0pjUtjpiuY+0c6XETzBlBZuPg8behPJ7eUh
gO+ELYtpcdSU1Jk2T62ey153aKOjILiSn0d2MAMJKxBsMW1MKxTTdx3E2QkVykg7
ovluLlvU44bFA0nY6lixn+FfLyKc46IKFzqzLu/Wd3Xo0Z9CNfb6ogVVfgf2XkFg
urE9+G0M/eLOD+QVEFKT5iBm5QhggC3rUbdRyuD4fBrYV6SLshcc1ZfngLMMKwVd
AZ1Sng4F+30L/6Sg5oh8IaQmDlhlu2svg5QAdNpV8h+5SsKYXJQcbN9jDJDKoOik
4asULvkF6FTfCZGbP8XBejrh0v5t+5OauyZzXQ1xAnloj8RXVIQCvnUVB1/320mQ
Cj0s7NQjBkutFMBNAwWvJ2gO8mRhyQfP0Tzx08Wvh4vf1cj6F0e66bPWFCWWOG62
mrXDcV3K5tt3z2O9XeVbVs5bm8MBF25Pmoh+388fvGg+aF6AOdYExT5FRXiZbR6b
YALVSgFozKUeICDfpBr6bsEaEIWCF40dlr9PKVS+kgM+9eTsnAWrRzzkv9rF2Jab
XCWZzrF+RDkfxPMLO9c5XmZGiqF3H3FMZgGNPWXK0nMfkCU9xa+Eqtg46I73PE4S
AbkberkkRZ137qUZKpnTVaQxxlB14tPQdCkkyAHooVneFjBtNBRg7oEvoSkc6kwt
VISw/xb6cooPArXDrHOwFijHWyvcqLWnYjxbs/E0mhUWUnPgGPfuPSASneTUZnD7
9x2txILakn5AzO569Xf0dcJ/TErgBmGcHn3rD5raMPJ4U+SU/fzxXDqFfah+koGh
8jiZVBnYmX4qCM5xdegoKow38I5vnN3ceTWKm3/LwD5uW6CoWQY9LrDToJDR98yH
H9NCQrTWChuIjAciRhMl1Upkr8nqyjAqOMiOwdfuB7E7oXH4ELaK/5WadSct2ahT
m9NMk9BCA7ECUXg7AcevvyuIbZO9zTCrcIS+0Icm3ejyKyVpOiyEaccANlHFKFAo
QuAe0A/gHeVujWOnMm/kXlv3qAl7rOZAbMSo7DaVzrXwUDnMf7i5t46uT2uNXl1i
J+FgI2l8i3BuekKALuI/lUK8wtJNTl5Pyg6dU9FJaGDN0h+NGzgWnBsoCR5vCZc2
tX3ZPIYXgxCI4A+/o1x0htD2Bo16YoSEhLIt3ly3tB3kHmir7vuHxBab9piQjY9g
e7vm0DUJ81Zd4pDPbhC/17fO0k1/KVJLutLA2zFCK5qRN2gYxpuw1mZrk2cNimKj
H/hFpoDDJoxc7zTjUb0n0up7SOlXdKOKq0Kx7HbWHIr094dRkWukXaBJVK1ovmdQ
kG0jZbOjxxUY3BM4TZTGDzKAfTV9C7heFP5GtwrLHlJZZywSJ/e6gAeXqgyHz5dl
2t/f5daK6118SJVUT4B2QTPGt+KrJNEqz5OV36INVqCW17KDDyOdTO++OOY0b2RB
k8ARCLfsU9Gg66wnD5FeJ7hJAjh0et5h59ZBbEX2dX0Ccvj3Y7NCCD3r5pXKKmF/
u+NMjrFry7Nl9OxtowAb9DD2eMBy2IfhCazb3ouMX8nuZ/XLPHi4fDLbtQbvffXN
j+4MF3jl4hlp+rKNfvWtwEdrZw0JNuf5jwd5FDzYZyPsLYFtdjgNpmrStd4pVDZx
SYERXE0Na9JrG9D8e4nj1LGeM8ODYlmFAtY0Bu1QqWpywfyjlGoXfgcEhbgWqYgb
4IQh9Vj3BdnrK/6tpsJIKtga9Kp+j2AarnZdwDcET59TiIwCrwh2uPlYZXgvX8EI
8Gw9Vd1P6rVSzkC01jgwMSvYCqJaJDr6eN2zJvERQ5CohIpUn4DkYdG9ScMpwXZ1
7q4C1SDnCvY1gVTRWQlRljTlYFNwt3kFuFTDMTLrSvtmxSuV65pd0rbmVU5Z+aWg
tqbFAKWDPhWgYGj61IrpP6uGUtNqFr8n7FdzkY+WGDsMItanLoySXLslzlgO5O4q
iulukV3W/pi4eijwircDmtMGJX9sUMM3+3s3irSqEADJ+gaqHyCaK8+mNwPiFzib
yBl4C5ocdqHAgzA8MX3PeI1X2wTPRGEqJ46OJX+n+UAr3m3beT6IGSDzAGYAr1Uc
sppkrPV/afjoR7Z38mkJ4Es6lomYcTHVyjFU4El7CFmJ7FRGVxXBUf3o+HtZrhIl
IoOGPQTi35PNTg3w9DynlIIzQhzBiNT0COSNTaCWFEFQmc46GJH3Cvq5XaA5T2Sm
9UmfjezgluMQTnX5S+T3svombrap1U2QOJmSf6Ps4CCMk9WcZYXkntMybvpLs7KY
IyXLc9vc5D2EQDzEnZ/IPLvIpJ14pFU7g4CWc6shFFK7KO4FbxxeZS++V7j0yWqY
wqzJ0Cm1Rn9NVUZtBCrw+3I5AkzmU4VJkjHxjJf5nvJtgCDMFcm+gVMNSZcR72gA
yAfhUPf7tMxkKYjwM5RSWxGMRpR5/5YxtgQHLhBocwu21Zl22b/yez9SH+azVwOp
spEbIGgw8yOtBXFh3TOTkAcYlWx8peHMjK8FXx0k592LM2pv2aaGXOcjBi5mOL/1
pvRCWHYKQBDqWCUm5wxMB0vh7Or0sJB7KNf1HLjjjJc8zZa5t5jMijLzGQ1rzN8F
MUxJawb0g+zbg8moY77TWHVFunIwDljNX5Xk45GGV5pwYlDAqfQ+R3dYkAH785ns
iHBm0WiQsRk8FnMyJYbnlrgS6m8T2VsS81DxgktsI8NPlB0zCH2tMRXK3Sy7AQke
lLXTDQqFEqy9iqbwoun8wQSgsVnyhAuwCkHQ7kT2SBaly0osCEABJkMkw9+qRR3C
GhL/M9PWW+lSyL0Lt3H6zDtVUXQrbUlERQMlejZvCMrPnyIsBLHpgnmybRcMcHnU
HIf9+JDhg570MiLTMSERSya6d3xhI4rQQMIlAGUuIIjNBEGR8aGefgfB3L8U7pr/
mely5HUmuBJkUTMoOX0gU9jblGMGR8clNcOkEWbz2FAHRsn9lFl3Jq8uzcOzO6uv
plvJm5IT1iyI0yij7JO8Q76zDFBwxkx7xo7YXcnG3Sijq9ZClPK352EdG0GmlHcn
0G37R761iIlJHi0zqDXOgHMoJUbtK8H/PleXTM2XEgC+XUir3hwa5HjpjQV1O14i
c7G3OuYc0x6KUB7sGmREdnB+nWJ2f5r4XDniLOO9wv5RTpH+lw/Kv9DDiJPOvZD8
XRwUnWG3u7sLrEdJn22z3UvmW3O1Rl9zCCHCcbDOcN7E8Yg13/9JK1yS4Y6yn76Q
radla3tf/oekE+3OgxUzToDblX4+or+VBJaWLCsXEXnY32yBTcSEV/nFqXddWprv
4z2YejwSOtlzlbzh847gOrlZXuKExlDcndbgB7k8Tlb51mh2havIq/rD05gnHha4
IPY89OG7prBSWvv2UxuMhlTP+Ib+jikCzN5117+s8DUf2CnJseQDusmC8A0krg0g
VoPg4qWXMDUKIQTBJuS7DGw5fON+KPQY9X+SgQ7xXCoXCMvT1QaGr7D2zZ90+ZWZ
Qhzpd7rDcoeL3qrxS+TIc85D5nPtJulE8+w6lySAlgzfoCiNeQjPOp73Fo6ABFMd
WfLEDLBh3/SVglzNCoSjnGMD4pt8VoeykP1DMv7fcdXdgEqUPU1ctbrl1DqiEU42
ERa71LKKfS7IF3m6g8XCMTrHIUaHJICz7mI3HWxtFoCd2QnROEJ8CSH+Qv+tdjWp
CSsziSVsd24k7mM+ADd5x7tNuEeRMu91ETPQh1Z+NG3oNpnxbqSh0B0ZTXM3QxUE
DoYviJd6ZDADRNGc1aa2do14q/RoodEg7weSGm3SmWJn4LS5YvOUtV+oY1H6ofhk
cZqlnyHMmxAVu4rAbWnJJc7mfrLY71lPPTQlCizBhEFpVMqw0p9r6Onoov8APB5I
jqz/nwU5i8ZIIkTXOk0sVuVhexyal1O3ZgJeNB7SJZMuxQN8SkW1FVm2rGAtpENT
PYTAIZZmNtmw3wovty40YCU+8jHYW/+GliizckQrSRF9TgvF6e3x+hPffEIrXlcN
XblPs03AS7pyYHvoNHjpJBYDMqLPoPhU0tHu36+CPJnaVYJ04/5VfRrYHRCA73WC
odAS6i9MrHWjf3Xp8nkAhS/0e0kMSK2lI+xFudxevfVMRnuCyM8wUbgMRh3fCwuC
ptrSNjWvYN0KtVVA7IQaHBcKqXKZCNHRhLVbsbrvqdscB1L97y27rDFn85Z+Nwkz
4EMMJQNrJRfh4OzPkrTqvBayRIWWOG+f9Qy9M4eQsmIaay706nPIfG3WuvkDDCBg
B7iGZvWt4hWIAMBLOqwiJjUrjqy2hrnCJgrY3ZDrjt0ZdheqxUkoORyken4MMqnk
P3sHzwhFUVr6psuZ+QVWpAue3Px8qeoM7VMlb6cL7qcbjK2sfyWZSv1m74Ju4/np
V7o969ESysAAnzVTVOgGkGSFN+ai7Z5rB94pztjmj1WybKz0CVb+HNmNbR6H45zE
265oCSqSQlKtcmbC18MWR53t+B+6CguRBN8Rs9BYUQ89G8oCmUfPLqKO9lGSxWNA
wNO/pzv6v4mNhd7cJltomlyNrHmJT8hmTPtM8MKBkIY3WJ06fY0EEr3n65vdxpUV
U2CBAyrsfcm7BfbNS5gxvL1vbqqjRp/R2PKiUNNcndG4K9q75K+gMScBs9iBFsxB
3Rrg79Ad2qX4TnOpgNpjVuV1onNheno02HcHv0gXkXTDV6i9DmzAUAPVk1zu7Uvm
6+2kL77pjaG5iOysTqglZkroZhXvNfgQfCYeWdnLCopQTcr/es2m4EbE1L74zVcp
2ebMpe/I5R3PSMindimZnKD8dmyEii3L2eNV7uYkrCERYois/IfcAVIDr8m8u6m+
njQXU4oEfma2wpO9Lo9yXKPqOC/dzxL82JAAMNKNUUOUcMQDB7FEqGm04hl8zS10
RweWQwpaA/2JCkWsEL/ZLNbBx5BP9/BYWj/yRY6Z5+o8+boCRY8WJ2Gw/4nad/DR
yMP9kOic6EX1ZrFmOJhiVnSKqvcyIsAdn0RqUCXQvNwvZ1ENDXz07TCsxyGJdll1
TWteTFd/9XcNDpbs2+Mm4VyBcpz0zPkWtOT6LP/UOelDRsqHUh1vR3hTHiyLzs7b
O8UIKmB2lOB8WoPY9Ea9lZOfTavQaZ+mb4xpmPju9T/2w1M+PNRdkE+wmOW7cZZr
Km8RrtVZNWvK3a4wFpAmGWP46Atz3aP56EG83d3jmGXwtFI2rW8+vVKKEkP416KP
wVyAP9xDRIZ8XVU9s0/y8BSmPx2P5Owb8DY94Sbs93eS0+pzzZ3AYdwStUlC4tJq
4mGGE+xKAMG1hUxhCevcsnu288fGklHAt4gVgRDF03XIT6ZAyaNonCR7AapX6PfH
me0lkL2NdUmoZGvj4MR/5keYqmleJsa1dG7XcniRl16/32HF6qzGkVWq6Y46W3i7
+eY9NPxjnEUKEItoTb34xcpXOgDvG3cEy3hqEsikiAuFAEjMksYkm94o7qED4f8j
iOO5bc4kMm3sGGsF6GxlF+OzdEEAJZ/Pwi7vlMmg5pCzIpD7eqhBFgclkbEHEyuO
NbebICGnfO2DFjCt2IT4GeYcba8Zft02KV9WkcrnfVXR64QMfzmUuXggRPmzciGt
2aUglnKNp1/R9Bhh1ZzaU9XC4PosrjqV/odaVoPd7DPJWR/7qwDG4pNAYz3xDwX+
8nitoE9RGr6snuMhvWrhCiE7oCarAWBRHsiswNH1Ya4FL2kU46OT10s+Byky6De3
YNJHDJKudo7QNxPD9dBxQsFTuxPKcaGHOjyrvDG+kfwlmTRTgvspDGHUgy/Gi1op
Msd/S7LpoK1LSoWSojS8vyBoanz+gA6gDWSJkAbgkFoWKYPHntvGRgxxeKQvhS4w
nUCea1YcsymGbnG2wEcqKXkVmrOC1G6nbBo+mOyyPjLNTjTYG9K3uuqGDuyISb8v
wp4UZgxzOsJ5YQDpiy038Zinm0ALWjv7498ki3JDy4kcNU/rpb+zhQGyrUi2BQSN
8k8s2Ge6tp0I4sd2CfflGB1tH4MrTpK0UZzz9RkIDTCwlk4k6Ws1XKvaMc32Vvd6
H0BXLTyjv6s8Ox0mLkL8qFSg+xeGIIvdk6WsdCZtFBMGAfnDGD/w2eBZoyM5Qea+
g+WNq0uDoOWqG14PKPCz2pz2tp2A1sG0BQhTN8fZAM9eDl7Tnf81uoqYpNOLo2L4
ZXJ5RtGAZHfLDNgn7dWjat4fzELOQMiTbrRnzMPPOaC2GCvW8iRG98HSSppm+4dV
3IGdkU67/Q6JRl6tyiJmozSlwd8Nr5xF89/YNWjl6sD+hvTXkIz5XH1y1YXb3mjL
TIHoNczKT4kNGf0XyiVkk3ssvkCohRSrPk64PgbxmULbXHfn0AFnvP9W3WDd3jre
asPUq5+BY1bELqLffkpRYSFwhxpUA5pllm2+7Nqj5BLnbxHWOKn5PDw1Ov5JYhmZ
Pnp5laXLa9LbnqyvsaMCTdJPAa4E21rWq6dC8WiedUa8OPQf3+OVoqbKmLQrLrmJ
`pragma protect end_protected
