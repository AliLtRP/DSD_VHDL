// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
g133MZLVGbkFtyp+RstN2GyKrr9T5tLjb0q/C/MZgXnJNUKTsgWN2+ZwiOhohYklpYNooiGXxD0g
op8IA4E2/5opsww60tQsngBUYUI0wo7XlewE3qCP2vNb8ocVV8o6cJcsOcKurjA0PttR80gYUFkj
IthE34yLRxFgwLIDE8Ljd81YzrRCLCWjZ6l4wT2C3wcYQIOy3wZrbbURBQIrYRsmQIicH7jnPGo+
1mxIG35vHJ26zLG2x7tjV8HrPCUD1XZyPQl0LJtIBOnhd9iECmh65uW3IKMI/O87sWD3B4tE3nea
SmIQ5B0bX3BNgOGhvcWdpoFN06I2yiRyGHTiCg==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
xln0pilprv9WDCebDBrqSu1mqDchXF7Cz1XQ+ScRHxzSIEoD26PBpbri6LwidGrSvjl4rYWX60bO
lX/UbudF/KF2Q76bTHgFmZuQnkaLyNKltj6YPNm39htVFJ89cwpfKJaKbX0P95fhhUCddjDGkjKu
/Muk5oaYKVReyLuIN4dWNTu657QsscLWMTJ/tjp+wYVpx31DBmFU2EyK1NnDfj6dfT50Fdpffvk8
RIrDiX7TOcJuQUwelnzg2jVqyakp6iRtlvbEi+HxxCy/82W8mpgJnk7qjrhjKtAicALiQqcVeR7C
j2h9GEUZtwa//+MD9lCtdVyzqwKA32gRqrqXMR7yz+hr5x11qZTAlZSzRpEjCtBoMlcHkgjtAmqk
yJwlkj/eriNKxaZ5rV4dxwTAS+3HoPAPZZ4+aUqpjvc3T86LSnuqKweaVfggpzTEW4smeP+S1MqJ
67WB9F9W2HbnRfUPI8BaBo3/Cz2IHShAO7Qbg9NGcjiLrT3FrBOsq6tjiJUqiBrw+H7dPWRJZ2hX
WoCaApwcjq0I1VCLY5QzLRaTHyXJR/tUKz1P+IQfycSOsn5nMMlc29SLpRcQ73iTHoPCtG6NBCXk
07txOyEngKVlRYab/naVWBfM3S7I8haaxkKFZj4w26gFRRXmsBJSelisGA+qwLH5EvJ38iu75+1C
8GwvcOrwf3EOR2hdWva4r8YTmIsjxBuYYn+fVaFVWY/43WyIO1P6lthVYq2VkfCX6m2VOQ1VErxu
Ir8VORkjwkWFyjnoVsRwGVJ4ToEMwRvIGQchFdgSWCl0VU7RAtvyvuTM1n/4QECGWQfngRlJ1d+m
L0TwM5RmGPj0zcTuVg9YpH6JN046Z46fmB/F2z8KAAvuexyxG65gc0yRcpcQLiOma1wIVd0FZeRm
CT7vGTuXp+6ozVH7CB+vf47ZrnzRhqnfhbH2YmC3MKd+QTb4EH9IcVc90tpMQl5PELSSHUMBMrlj
SXN5z0iuBM9c41GdLjLyc5A8FWtPKPCXAUhiynB2MXPyVUyJn6TEzyZjj73U0eosIJMm5hWMiPRq
gfz+T97z2WD1gj2931OuEsR/zBWliu+3SNH+5Y43Neg4Ppxy1MYoAXXeF+KByOJwsPTxz55td2lv
T+lw8IBKE1GeA9151vNlCshcdEawm6WVAjmRyf0xY3ugsmZe4o+iw3eIkjbPCklcuL40Fq/StqQ3
8x0h8oPEofaoRmgn09Yvz6ArBl6xtZIMe61l1id0LvdVML1zunF9Xkqha5Sy4y74dDKgNVoPvpy5
UpPutSWUWL0j8tijFOmd8XVIDd56ZzqXYTCck59FQ8qho0WqT6Ojtlxeo+TseB/asPXnedsVsA8o
UMqWyDkcrr4wvhoZZfnQIXKdhWPc8BFG9A1ikvUoD5LkXMOotctXPN6W0i9rKeRStKB7YLPY+gkz
6OlhjqoOQg44IVgZOhIA2XadvdRQH1qNLIKTedXW+tD8Seo2VU9SSGv2dd71a/6LpGSv2n9lpYzk
vuhjb7bQwttxuvex3PYaq0pRzTqa4wMr4tbQD4qkMSpcpfxrOZZWlOgIaMsUAuYZvJ8ciID7scgY
87UpmyhZUtt9Ce95uPanbqjx/RmCEqSxQlknCFdriP1aviQHwlJvzjyW5yuYadJ+1PryhpD7vAQV
pPkYTiZjGxgE457D2w9auP3O99q16QbOo191Qc7Y/9Y+tz4rTMsNxIjHjwaGtW7SCRgmLkwZFDaS
m6oLXdyMK3Ndkfxd/2XvUndg7rWf82j9U0wmMzO/LQHUH0D2jCSLY+rbfJsx0a4t4pLNd43vytXg
O/O7EP9vLynAbmHm7ZcDEerHMe7ih6oNEgEJqC3DwauTwm7nhu8YtVEX/3M0p99AOwKP3N95g4Y6
nB7TakeAvPSL/DdsphbTmv8MTNErQsBCk+s9/jVdxsdPqQeQiifioWdqUoHGXByEjCYj7vMRKgWO
wJ0gOqFvahGENJMBTEYSKNSgvzY90bA+mpC/guFPyINWkoTIDm+W9M3rWaOkpB5ePittPTI9pXby
35L9x7aA8cnBWsAyqPgfmUswH5X5NQ9Ov5naZNS7cKJ5HwcHC459fWZtJOBdoIr/3WXQVQ1AXB/f
kv0Rq7IHqFESn5osnhNzXqWfjYAGD5ZkbwTnbl3c79HGeVO+D9rIRI/XDsNJsuPectF0DRl6Gm1l
3rlmPMzJ7jOCiLQp7W+h2nu36a7Yv5dwlaI6B3f2AsOdo8LuF4nwcoEwLGs2OPH3myI/rjrcFGhN
RX/pI4vk+euc/vbDWwIOj5+hQc9YvAiKCbwTAE2BNfV6L5pcRk0czewEu51E/4Ray/IhT3wk0ZIq
DLx9XVdpROcRhFNCnEvm4I7AW8er0GTvmYi0/L9fiAOYHWthnXFlbRobY6sul4Sj9pQIwf7apX/J
mhc4MS6QS9GY+GoV4HWTQGH0EaI5w4O5mUZp4X1TSGylEnmsjZZR/IG7YjmbCZonvpm3PK3YbNDd
vAZlelquI+tflVXubaye1y4fWx9HQNMnFa+/f83ySq1ngZrpVIGSYP3TxrrrMqJeyv90nDo9NeW4
HNxssh1SBaQykiSVL/ZWKXycvRHVX1mMsGaYwwEK6freB1pVAeiDGrTCStcVLZCzRVmJCWrDr4OI
3sJoubHYGjGHoo8sYE3EQ6AOvA7qKvEkNAgDv6gTYflq+ajXVleSNpZBsWpGYRAiAXm69q0sfEF0
9pKDxs0DT1/T6cCBb54IPw2DSCP4E9ebSvzBxEkFEAE/fXZzdOSWQjWwCiKvh4K+o9B5/utbAW1F
du/psLa3ufhJgJqBvc1X7INOrHDBzjWMm/reQNVw3XMH39Dj7CJsw1kbEvkmkuyuXgjvjKrv+8sm
F7/GZtxSAJRxv1emljIsf8g/p4SUSDG36EJDPSzLTfEujRRFGW//4J+n7xDPqYYT3RWvu6isvEIv
91YVp9cE6h6lckznDyy3EOm4sxwp8AZCEfVLye7PUMBmRdexiCrHPebHNUUnUXR7tVGBzHkXP+Dn
7AAnSeROOU1MuU1e4EPOtiP+H58eZyWP5Xe2jxD1lI/AHUZdVNHmRtx5zJEWs/P0KVmO4N4FMZfO
g2gd6UZTD2cENvxiSKkNAHj9vjsvjMrqFI2SOrH6TUKFxjctkcxuTcXwwOyjVvyvBKTuzTZRvM8r
Pk6ky5EPQ6EqRxXZ2t7k4xwYkZRUMESs+JPFAwTjnrLbkJzbwk+1zHHmSb+KUyKulSGdNbbGMokf
Kcsj1u1IfiBqMKrHYvyZQ3uxiU4InwpQm1sYOAScyqhBJt7BOwv3zaO//LxDei7f2nKs34HG4UQL
rng/keH8o/4n361zbIgRmBlfpBY4htGe3cj+RixMHpMiC+tol4cqi7/hLoVj/QHjHzhfwKL+yrFN
CZrwV5fQYrvcXw/5n/yrB1vTCMTGOIOl5BAWrir9koQc/wU6M/i1tUzXQ719sCwlnz8TJfJUkPWY
DJ0JP3azZv9UqCV9H1fCsMYdFaBUw3ltV2zItDdvc2nk43W839wn2HAo47e4Du4L9WIDO0JNGwn4
koazlWddG6FApIOfsbxkqqQVaYhDJovMs9fODBaEjyT0ep2smvGnHllHlxaABALJAMGZ5/fy2kjX
uzNKJeA/CVQMsf6ATOJGangRRvRQ2w0ePbgmn17e3fDlwB3mAJ1vWBrENaGKddVWjHPhAoYY5h0F
irryWKVmaFL3p3SxSBwOe/hn94JyQZHqqPkd8h5fSzfDnfY5VvfwIEo2c9FYN7gCkY70TusvjTG+
clITMfOEd34WXiCVOym/g2Ys5/Pn+0zXtFTWg6SNa/L0dsLn/pTJmtRV0u/XzCaWalVZYmf56VDd
6p34+bk6FbJysLGGCwiYCmRVQ1bnwWTN6ZY46xN6I2YS0zfbHVpWb1AYA0ODSc9EAprI7kFDrqZ+
6jiomgBftIpqQ6SMf83nlodfIwa8C14TaYyBVEF6iu/YparNQN83xuEF5lpWtY15AGlVeiaTyx1P
XTXh9Se72ObVt+OWou7DVZhFc5wON4VHLYWrHZE1uzZ/6L/pJUoRdBbLg16HgnwJ6n5DzJ69reA8
Kei/h4bvAtWL6NLKSo9He28p4eNrIBl0pQyDfE6nagcj+bWRn+tkkDzvt276P1pUswY8Wm7N3wSg
BfR0S2/YmFGcxnMdWSPTEJS4tCD7gUPdsnQysb3QKWdIlfdDTMqzKfif4dnJB9yxdFmvoTBNba/V
UNQ+hGuxyTW2bf8CmjR9R5N4mX+hEhMvcQ4RETLGWsMb7kd8Pqjx4p44zfDEWYIdYbK+PQnpNgJ7
/i4UMaVotGZDfQpSMo20oFECvU063++so5RuiH0g6UpKTlnNRabZFAh3835V73p1N5h5jDOlzqyq
FWXPCSNZixj0uEHU2/HHVrRQ/c6d6ycp9OQKsA7BghVV1plgwq+0RgmMDYD6EFwAa95z4FIASmr2
vdbk5SwjD5COcBfi8aCRlbF2D8NxxgMJ6czK30z+5oBlJq1xEbAVsAuh23QJXdf9TNPqfwVxc3mA
3pqSI/4C6myUBVqm9I2hEOKZq/iQhlaOoJpx1Fiks6kLPsQhnDfNL6IEQuq1jMS+stFsGo8vxO3N
1U2aV63xfil7GtqJDxKD3Dr1MGS4PpJ9x6v6RuIrZl3tdvuxr+utL2/O1vm13pTYiKP9HDba12tC
zFox367PHC89YP23270cNgB/ClrOHIw81ybBq/lgBTFEBDmjOU0oJoLeBDPdCxJFl3qlmjCJqy1K
+FkEQW0xkHDZzJNN+LnAClmSwUvtwqlnUZIPp2AvIucri6cV8S27VBguX7rzBC7CNv2FgeVqp0mx
FEwTMUXyNiPj3ckHt79sTLamqjvm2r/lh0VYxjyS1Uu8q9iYKz75pKtDNxFcDMU0TIs6aC7YP90J
pw4VFpEjgftRnx1t+ywtrAwa7Z96swbFhJlZAToynR4D4d9UWfpsHhhPnM4K785WYrrzU+nAVfeJ
pB//1OvCYia2oMUcS6/0wzwlEmgY5ciNjlEVyxjyDDEub8IYmkhyu3y2fmYqLluBRBZlCx743HOt
h7DsFxzUOaFxB1nJfo4rf50BnXm8QH/VoYHlhsEfex2FSFNrrjgFI7E2/7/0PJpDvjATc343ieJx
Liyk4u1x/6Ijcg0Zqg37CWwDXL4QuhvXdWfOwrnXkO5/5S4rRMm5fgm5KeDHJgJtT5tqqospuFMR
8bQoEfoeQl3a45wUdZHzBZGYh9ylRyVa3z6iWKlU99DQslXglQFspnbAiQDKpUW2F56VzAuRKojB
wKfLKlVad+/ITzRLhj8X69X4ExFtSfhjYtsgc3jSGUK1aVyhDHLRVmZ9K9WHKB4YshgyIIGFBz26
Ngw6GxL0OHavG8Lm4aql325pUjCqYlRT/ziZpF2UjA58jKXUvBbE9a7mfzNUhZRWF5XZ4fCSRhDi
mibtxwGqc6zEAo3OlLEUk2DoqGsZ/st/yDSe0KaIjaes1X9D43NxIx6o6zfUBbrFxGddfsYlHzdC
VnCm1hC4onPhNB29WlP6hg/ET013adXW33RhslritWGbUptwkvtDqW2ibWUTgWEyVb8dli/Hj2oF
tbuXRNem5YR6giHsOqSueAphtca9e+D+g8JHx9FNOvdk/F64C7TqQDxFaQjeuzkYP6cPQUwjPhgM
SnQscleHSeP8TNmRDIbU8T9lalus5SAHiJz2Ml3A3aXWNpYhYjNAejbeeQo86rEQ80m/PnLprDF5
ZEbR2KsNtXCpsP0zYHoEO62bOZF13Q6bISjvlzHooSV3+fc2geVhIayMRyJgHDfwi1QQf4a8hUNR
tbmOX2x8z4g4wjcowNlc2gu7Mj9n7HqAoTVIfkN6/mtYqzkfTKQ82xud6o61vL4zNONRd57bBYTd
n0Tw6b34Hk5J6E16S0aJBWT9o45W/0TBdjRrOTx+oSKYAnbMPJkqsW61sGHanOBavIvlxjn1/wWx
ZI88+gWbF0JY5jP2c/dE2Yi122x0RifGMV5hxd6FPYBn+W2pp9RoTGefeFeONlXpVVa4loEZ4wGU
6MbV/mHtbvyT4ZkhUUZS/W/b3ASYuQ5M/QK/Pb5YP/LXtKRHWPXhqDOL9DTRDu8+XyH7WJ4sFAui
3fGSzMt1WCAiTXBS7ts0p99qYiYZZq2rTCJ5JaoYmhgwGwuRnt87V9mmADDiOamZyb4pwd4x0/KF
d8vEyQiF9w+HpDQJ232N5DeMexr65VkEn8hguiivzQzeUc4OSQNviURMRnkgmXxQ5RR8ayZb5SSq
U5/mNYiBdAP1VMsoPVjdQ0tGNhQRZHcE1oHxDDQc+16cDVcOthwwnOmga3lWnVRuIuQx8aiPAtUB
e7qUTgnSQwTIqrS2WmaKmwIEcbXjv4ZP+GXf+BsiSkloJMYfb8y1kEeGMQEDRNUPtI2x0bOSb+9P
vzjd0Q7ekIYQvqnQfpyZR1CDk+X6OJl4b51A4pZ/IhMqqjCW13liEny9aDDGdqSi3IJ8pSKogFOm
haLD2gl+klDBARxhN4CGu9h4nFQ6PizgnDhs4Zt1HGW4PtH2XzFRhPZb8pMNt4xt+IIJuRz7dHNx
uMGFp/VC8Y/z0jJ68sMt/JlmMYckwlTPIqymx3LKcmGmwQPFjDxEZxT9YQoldAKJChLtloF2JbcH
BugEYGpEEKgJDguv8Oz/uL8Pte84ojiLqBW5I1Od3UKQnja+v8X5QaA5DArxAOgcVStS5I9wMmmz
rbiGqLiMo1cktPbUoClroFW5jswsGnzeeVhz2+1pn6qt6HvDwcWOVz6DQUGu8jerCkFJAPCTQScH
Dsd+SxeHX7+Xwy7SDuzakUpv3G+95lrTxOK9EC8RLAMk3WgAaszAsLhLuDJs0YDRyyp0xbYK9ULX
C+0b6pFtY4XVuW+zl+jQYbBXgrW9QyvN5Rn+7ftiOJQ4548UE+xaC2z8Ce8hLcZdBoULBatpwb/A
GTFazRcGMgq0hm2hphQFZ5+DolUcN1D/7sxXPhejr2IJqY9CUNQZo5Zv6QGcdrFY1HLKNlqj5XlX
b9sZ8+wGLHr5CkDQtoCksqrAFGH8fVfAtjfOeI4dl9Vy42NPEYqIrdollQ184/vP8rL6Sr6N27t9
av5/zozgeubjJosSCVXiLKYWVt3bQnlAO7lh/+i7ECQRGzftX0sFPUOhcNN9JSAUrpHEQGvwXzDL
kiiqsh4Vn2VPyuHsmC2yjfJPdB5O+sXTpm5BhqToZ9cHWZQk7vnREF2uX85o7c9wG87HMrYKB1vS
+GsdJ2fQyMjgihKWYJMx+AaVHjNdbPinsGJmyJGOZajZoT9OL5KC8ISsiNxMretaHDjkBKJxssTY
st/7uGnJwckK7qZpLXVRUmCvQYjDZETUxHJPg4C/rQv+tykoXit3VPR4L7jfQF0Hgw8U9ueRR5g+
/P9IsWzvSmj/xudYQbbD0YAd9QSsJ5y1CypSyLaF7XXXn+i18dSDKbQcyy9uibofxdqvOcpnzEFb
l2qh74qF4OldpoELt3ef53qSgm+H/wjt2G1QiQl2zWsyzm9xffB4A3nKHV14f+UwbFu+FX4z7ZOh
V/Ps6h+1taj5ha3y3V7Q+t5B/Y4ocw7wU1Lx0XABBmFXxHuyukmKxfjVf9yaE21xFVVtoKsim1cs
8P1GaKetnUuvebKhcI1kMAbBilZot830wRODTZlhlgtOVE4ACwxBqexifU59bzC+o4I+4hhDK+hS
PICXLSiIZLkCXsFOE2DagZYhU4onth2q0u6YJApfrpDgco4BtyvZCt7Vcg3C/QvAJEcxVmEtfE9o
9cfjz/v1iGhaJPmOYhx8R/+3yrUVOBwxafW5BzMOTNBxRbDN5zRi+CjpF16tU6OIQXyPY+bJb5ED
qJzTD09w/MZgY0b4RjU9XbQawz1HHKvjaanqkurQNYHqsdhkWzaNyfKuF20fZRDDct7q4XcJWP0F
2vJIMdhDgG3phu78F3C3dtmzGo2tqajskIvtZNZN/GXtUP6QQf15gRVg3CO5zTdzU+muf5Zh94n9
9kAmw40iu7BtQSYPzEP68Oi4nsHulv6lQ8ImB+KG45elFO4qTQGoGVODmum74d/wie3wVOeOSDSI
BVVj7/WqVSPE6i+71ZXeL8VlN/SsV8W7Vxf+8/2YUxFoT04FBaboMTAaXIQy/3Ut7dqc2hln8BPm
UH2wckkEW+qqKrLTxC6aFspiGbIwkA6xHJYw2lUhWMSMf9r3jh/Xp1PjISknUtapFSXkMBDKrsE3
Wih1Y2Rk2XSy6IpIEIl+7e0I4FbLrFAD75YwH6tA3neVrblUaS56IhpS0yj6UPpKMWQG8JsWK0u8
9YTuEXoFoVuAWSRFmw4GGXnLeo6jEbFoc9K/JJEwgnrw5M/DlZoeSgd+dbstaQOBk3i6644yvq1O
yvaVCH2ukC8xe19TiYdcDaaH+oJl4/LcRwE7th7LQHyAepjo1RR8Gas6+diD7RCJdfLIq0z8bYuM
64gsTgIuKaA6kpkhbW14t/zuxHUuDelP2h5hRuBY6VDcBxiExNIcE2olWNKRM13UkGx0/YEVVPre
0Y/RjaBluGznfXyzTuNJJ24bzOeaZ/jIOZY42rNrLNBCE/PaS4GARFMMW6M8FWuuSxfb6len8zw+
UO6EFSRDHmaNIXWy3Q0orKJ+4ljm5c/48gt9nUaeTx+D6L6n0catVzPmFvr6uA4gl9f3PUx9u8d0
qFiOo/RpF7mG/3QR7Z26JoPCA7RymPFtLOKD36dV8F75ADYYpm6mjFlglwWuyDbYfdn41A3JcaIm
YxwhAOG5sKYlutQlvm/hhappV+AnMsbvUNbzaY8bKrnaJ3jlPoEt/kfKF0FZrghPD8ADR9eUEVeT
GxFTpHdmnDI7wRrGLzPpTWJkhVy9gSYDCQipbhU3HBM5hnMfPFMMaZUZS/PiQ2x9GFnXp13TLPcV
vqZv6GXe6ME9GT+JRTboiWxuFo9beWQ0gaRyjh63k9HKA0si9uuv0rzTPQGU7Qn3Jq5ECkRNhG8R
qKTXND7GjRQXSR6xMX2xzTLYs4oSHyARmec/IIsCtFmi+UoPpwA7m1nxZ7Mf5JUVj/WbEJ4h8WzI
shvTlJzgVGrD8DwHVbVFtE30SWEN1a57ga7R9DLrQZDlaN0JzDk0bP+f+yev/KZlGubgKfXDGWuY
hQaVzFbLfYzvvLY+xQn4qu7Y0B/KylsjPaMun2DM/PJHHzILS86E+yPn78mHef7dyRZAYDd8ac1S
N90qNf4nSFHghxnxzyBTJEiRPjU6JM08ok8pdbEBWcReqL+vqIyELHDxYJcQqGemb5Mc8MmE2zRZ
+0z+oJ2Uc1vsit0Ag3vqSH30IMWYIN2klIfXmE7BaAJn2K54vaBfHKeB/TliNnIYNvsh+YbBPrEr
Wd7dO/ltFOxHp5aVLyu/w06sui2Wvhx8Ql57Haj2p1WygSIz0gxklIgaf73Kuj3zD8dg62t3VLmW
AuazAoc/LhjOYh/3Oyaxlrfixopjm+jamX6hCGwSFjd6OjI2k5rAsK8e9kA/GyX+cigZDPfxdoyr
xWJtKAgaqVZOOO5ZFR3xLeSCQOb/prSfxrnWHUQ/G55I/f455qcQGh/QqwFTufhMRHB2CBJ/5YUg
sdOahwdUuo6SbLkZtCZ7+SyFSFqOTKo+smXNZeYFehETR+YcgBRotlSir4W4V5Lx3lShzFhI/eEc
zjeeuEdcfYFzvmM2odZChNENryKEoOD7cPb+zSAKSf83oQ+jokVw8GgUlLInNvHtma9xsJFouRno
wcZJK/1crpmkv8NlvUKQEYZPvTV8gKxJ86G80jlex40xOEuWFGdBhhkDeoKIHYl7It4hB2nhAMnY
0LVzl2MZbu9eU9140jDFc0EvHr/Jjgs5qpUQcThxYGDPFmicOiBOW1gXJalelFiNeqQ5aQ0Ie+u9
KZNdqI4eABvwRXcPuR3P1JvCmkiuDRn/hV5joMLBB1gcaGybb9B3uARqtAoblbb6ZS5hisV3YuHi
FDllWHI5z/KPTNHo/EoD4V+eDN9M3Q/KLnnkPu/inzs50IXpWMkFZrQzLXJjMtitGxptUEb7OSrr
w68txDTgfc3wl59KAqhD7sM99OqXsPcy4kxLm/x7egrFyUzneILot6ZoIe4lLlAV6hr8MDMomxig
UljSl9Ua38VxCDsiLtD7m4L3PeF/l953i7GwYQUx8rbsjsMSJYhfwQL+ldnQl9HadzrnqJ/zHa76
OigzHBuYRujq2Tanpjgom7LcMwvijQDqVCIea6HOoYSVwf6wxxb7hnYTL/uk6TBczT3Cqm07zidi
N1OCikJoe9206+L4eXEUq16+qBhun6QPtmkJzQzr6+RKPY5M5PUW6dD0yhf/9Y595tdWchvwtJX0
VQIHXZY/Ba13PpT4X4rC5AjcUiHF0w3OxAm6G+cK4ym+pA1F2JHCyrlB/VO/SiqDHgq/lA3pYiQw
xk/EujFCBcAASXuPsMNacN19TtSWhZnn4373oepsjn+n1mF311Dl69gpFuthk6ck1PmgPb4qK7I4
6R4QaNfr5HhaI2xcqraVDCIT4tIXPgt5hJT18Gmoxy0bfHFsx+hL3mKl5Ts1NG3Vndm7S5ctFyph
2zhZUm8p32TTNLlD6gLRL5eyNXnGXpnxa9+7Wq9SxTnFZOm2roEwDB+bUCviUn9enJhIE88U/ZPl
nz0ryYD+BZ4A+3aoWbe67amuJ266exM3XeQCkN0EYXcjTi3ehA+WyeI9paiTNCV4PEJ8AKGnIFgx
UT63NihB1BYkMh8Igoo5+t3xEOCZlLrfYSYje7gfULQgU1SAc9KyMNjN9T3I0ZQMhpV4YPEASAXd
/O3tQyoBjBX9ZQLRc1GF5iSqGKyCalBCRfAXQS/IWUfrvmQs7dROfOsOXYdm/bI62EXJG7KzCr6r
tEGZlvyWHVvWbeUWchiZKYBm2gQgJ+ho1Ha+7LboEWa3RWrLGRlJi759MdZUaXLCcEoyd0wFMbx1
/DsFZioYyms28IwF/6S5ZVbUfYp4vkEOiN2v/bhvzvYEjECmEW9w5H09umvNPpXulCKrnEuG2Y1l
J8///iGhPaBcJKKKdZLSG6HZYx6QhaV2R4l6KXElj2ynvFdO7tZGmTzJ2YbFDBuM9W3KfG/pOypd
TEpaIvWAgS1At9uhaxYs7Uml5Chx5/J5jzPO9n8VgO8kIz8InCabO8mYH2WoF/c8X/chu+/88bpK
e7VsNyXQVa0bAcUWAdlJtjRUgGsk7yEvSrra1yKvJRRHE5LKU1Wxqkawl7ANFjyc5K2T7kxvwreO
wPuFNQrK7DL0s6iW6Qch+rUJCEASkAGa886S4khJhnHT7r4+ylUtrkhjr4bCZqlbojakd8270D06
PRLqs5N8qTiscQvhi1m+lFyTIQiY3xDIc1bUtx4fLiOhdsEo7/ZFlTzcuSqnMe8qK8pEhIxKScY5
h+U9oTAgu8BOsvtS2Hnq64sfDgBgvlfRT7lgzH4adk/m2zbRa2yXeyygCAcS4TZZ2bXn/fjwBKlP
xp7GGN8KlVG8mbCsgiTcfi286SPolUvC4gA8l6+0PH4Y3uLYd1A5yRfC8ATswrQOCCUwVBfqL4JR
VQnAYjF8R7BI4YawFYYKUPRC8NFq/LJfi6I0d4KddAwFnA/LECL4zbO3abRTM9EIw79XnGqBnyrX
uIr0LEpOoRAgaxSrhLZA2fLvi7xfISlCs7pXu5ZjFVDGJknmqoQYd7zEW31ZXCW+AoLSVSovi83Z
atV9BaAXavNf5C27bkBm/3FR+zV6pJTd4iWbcmDLuT3fVht8WCdmsPvGlJWUN7/e6BK5ip+fzFUT
QsdL4veVO0snl4cltJZDoEkQPObg4dys/TtkMCmkp5B8RXdk0HEiIWtnRQZ/BB3WreYEAs2Fucsn
xWA9suGFQdwb9gpXoAagr9kPz4ZTWW1Ox5hUbkAE3yDWEj27hy8jfpBmXh6iLWdxz7nKAahxQEwC
dTD9X7Zf8LLeH3EdRZHoHLQy9Ql5a/auvi8loMoLAihxaD4cI187KxfThTuIt/N9x/Ka4BNRT8Nn
aN+XOThd209zmXYB8Nf81wdZ3/xEDxzPS1qO1V2GK5y4145Ix57PaffdbMaERCpVfzxM+77eBjoW
wYvTPubLHH9dHkIv+2BeT5b1W3KN14K85dr+rVKIbSzmsJiPpsxHlldIbAueny9oTHcdcCoTnL0Y
Ql2UZjv4tejGMT2nWz8v0KwvQsl86FZs26v5xymRMOatw7EuW//SvW9IZCABc7n5G+L0SyhxwbfP
tNREmT2Gm8t7FoJ6JY9C3UzQg3Xvejl4SfcxsLHMUXU51eA3ADd0PtBfuMB+bbOH/6id3rpAyLVw
dPrNh+eoIuv51fh5qmzYtlK5Z/PXatGD/FCCj5AySkS8yp9m3MQzxhrOcnBbfGlg5BkHy8Ae8Yh0
3kSyOzKHkFUwiK37Hj98vEhmOLu5dDwKibKklym4CniW88edjP1pxE8BvW1wG1e53VnX9uWiaJsh
DIvzFO+MkI3oFB5ad8Ybehlba8rzH2986LjrQB0piE/r5gBP62S8j3g78Eg1uhCZb3q8irBzwn6N
++XRTyNBohf2xW4qXhX0pJSeOBrIF4XiXvg8+HNmESP6v4o9lIfeSSg6ngxatNORIV1W2RtNnRBq
o2RyuARuowp9/gwNXyQbhn2/81qgt92qdq4DOO8rkHoqx6mN3+swKfTV7EkNS4pv5YYboVszE2j2
ceJt3YQ4mA32IcpcPwcBMS++eSdVm1QjOfR4YsnuZJ4Sy66J9nU84LFw3knr2P0hgMH6ThZWgSTd
hY4xJvYjoye5kTRz296L0okCxcyOC00F/X2kbncYzTaH3Wfvb25ugjmGNJYRD0PKK/HDPLNwCBY+
PAdX1o5EZ3JH7K0j5I3LsXNi2rZrtcf3cvIWzTaYWuxZQjrPNAmxYvcdLa21dd3tU/Tc+cdbX1ea
79hrDNgoNj/8tvhMJX7aX7PxJxA2ien7tu8QxASP3FtEZQTvbEFT0vxhYLv+DWLwSoxaIvF+ecwI
+nErO8DWZl8glaM6xeDlC0//0/o6wjPwWiUkP7cqK3FEvaAFMy3uZdAAbjVReTes3SjXWhtYM6Pl
Ap3jFRfrYPZ0Tk4Tjo+LIyQzPkMPL4aWHu3oLLwAAXzseRwwb6qOCIiel+pGg+KnOtVOygbKkIdF
R5hYs3XOBCAbsvxLeN5llusLsLttyAHcK1BJA/pKZMUKPHHEUu3BO24sycKZeXLEybqNapIs1kMf
LYw/NvYf/SaHcWJ2+UwShSMbeV+As8E0ld18vmUzF0RXarIkKxnKIQO5RUa1TW4y1zQBPv2JRDMo
dVA1ElLt/AeD9iLklSa7CbboxMKk11omxW6WE/k/A8h/rfjovfPtVVWX5DB5x7b7/mfZhydg3K3f
iFxmiloalNR0e32T22RQg5OQy/Na4Dnog5OZWhBXlZkW79aeYLR7d7tLTd3ETHowj1bZ3Wx/XKq3
5NgFkZLbA+v7eextWq8fqHPVchnr7Da63UDvVEwXkynFiLhf2AXu8UYNQNQMVyw/Zm7XayEkVuwe
nQHVYmu9ACSftBCPlG+Ohr4u66b2W7b3xdfsGw6hEaPElGI5xc72AY86yW2kzH0zaIqYRG66eu1X
0Suj6LIgEuh74euPO7vZMRfe4b5nvympvO3ClEnUf2mVxPRU2cdUNN5LcAmPzjCogJMH6yDP7Q8F
RKalpaDazXgHf2tL+B4d3ACl9tvL2VfO1D4eEekYPldE8rZMJLQu6C7Pc7/JrNn3hLWNb+SUoJbr
pTB0keS7pgeNQHxikAcXJqkpgsu8Z8NTLUs0FSS8OTe9LWWbWtxqSCltbbpN2tclnRptZNAI6esN
r3Plz0bfy1znKjw4V702jBLegjAVKNQgC1CEeNKa+4ThsB3S7xGUj9Z/yy5dMBdHKVC6OWg1qRnu
9Nu7WTDX2LgHo8B/9kw9wIvZE0x0ImniDILTmhFeiDvx8Jf39NrKNJbjeuUUrtJByVsc/er9pDlT
AJ147uYdNLr+IzcFHXLof8IZt0z2O7vBkMrrrZVWw4EfHXqB3Zv3LLR+VjxEWvLEGhdCp+qxxffY
9jkLUXFqxyiL8wypH3yvMGdO/PzrARvJCWCsWN+OXntx2aqJzFufVFMM4svR+WGw0lelmO+GLwU9
YY9ejYiHBI9XgP/CN46Rxvq4y3+3MGUGNxGT3Jr1JHp2MD6DVLmDOCpgdXX0pizKYe4/NLO15stj
FobJoLBDmClYTgljM0Mnzf5TJ8bwtqDpefmvjjUUipO3lKT/mqxiRD5PhqVZhDeFl6u5a79Smy5Z
roICwHY5RI6OcN4rzUvKNtL/qSan3k699WB8F2PzFCUsPXT4Po+aoo1KWaucN/EM/LzW2bcROrID
F92LPcyTy5vC+fdupDsiteISy8po/n+zKp7dsLiT/Tb/EbRRcWOBNFSdPw7U0Sx25xRDl/HHZqZY
Li23vTwRuAwusJaFI3BreJcdqgNs+3PbEM20lyYKc60bvssVUIMD+45HvxFcyQs6wq0bOAppISIR
LKTf5wZR27bT4xPmG3EQ7jKnWdyRS2UjpZ5pFRECaAT4A2ljvQw0P3HqMym37fq4BybU83BNcz+D
ihL4ywVeehFj4/hG7zfMoQV/AQF3jYW+OiYcxSuX0Ghg7Jr3QjcWm5XDIsqihHFDcBboQQ3YLQ==
`pragma protect end_protected
