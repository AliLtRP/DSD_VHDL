// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
oPSbrqtLzTlb78JG6MvBvinsmqAKm7k4DoKul+wRlg8CYfXSvaILNiZt9xT20iWi2hJzZU1nJo+l
HjKZmLsA8iEDZ2+c0AkzM8QTmXf9PPDjNyNvsU9We0cE/GgryvP71nzEbaeD6M9rD2q8LW5w2bMq
i3zD8HGkowlSabr71sseCDE+eobLuaF6UOrBDBbJQ1OkWRLR6vYcPZilCXyUvziFi22fZyj+h7cc
Wts4RMlOLxwWqbnQtmd4sUONR7KzWo0LDD+W3e4Qe7AZ7YjwTQIRc3z9dIM+YWnRHj+5m0lkpOte
4Gi2Etoa+u1p3cXjR0t2Le0D//r0XQlfx+pKXA==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
uWxZwxMoPbYnqwr8LsMxHxQUEMusfjCiI2IkbaaEArjJR1m5AIhFVMFFyfjVtaIncXju8ce/1Vso
ifBpjmzIF478kIZ/xDvENbPDREjn/gU0b8ra3yJ3APSOjqXuXCawPUKWqkirG7REEbbkSdJBeXuC
rznz1Z0dsXSxzDdjJTHX07qjr8SB0wJG8n8EwhEkOdNuv/raGy4c34BiYxNdaUGfQ6BMe4qU07Iq
9Ln4E9pSXxkfP1OVsrXcKFU/COQmDaJm6T7ZQZzZY4gaDrexrnPxzcz+3g8wpcTMI08ktLBcTnhy
OWoeZCKPdV/0xkeQcQ+d7G0WzmqXi6JXsJxZtB14ucFa7g5L6Xjo9dMdHebpG8sE4s5ZzLKBKBfQ
5DIB77ChQ30+igXHVTt+/XkheHYoRBsCI1r9VpPNgPwnm271g2xpFT5P/0/JWtEpSNwHoHW+2jL2
DoOF3KdTKugCWV8ytxUx3vq8AxYXB2zXvxnFKrzdOWa6aXcV30lz/aum4lmVzchgbl8tzqXesilU
6c8NAJyaCPsDIZknXALY9Maz3zKELJReOW4BA437L0H+EiNmOrL6jcwFU0hLtPkIZHOQZh+vR9Vp
lQGz5BAMdYbpPb56VM5dTh+pYZdEOYwSiBAbrCDBQtM8K6KofTwQEFJBj18KinsUFSRD+1bkSwUO
5IsABjaSnfWMxCMvsy0ICBFdarFu0WQ1wZ+96ZVaCWneeIdgw2G5oUz7JZMjqqeG6HW1LhETyqVj
sBc3kt6jHdWzLnhBkXH91EGqZ8MqGRqEJobH0JpmWLzUeIZt7wDVIFIEas9vDM+vCAJqdTEx839P
MlA1MB6eacdgk2hTBTaY1JPfVEFHcrmaBIC4GIov/tXAMVOeYL9V0q6pLEGLwYeaHpTKURfBTNWQ
9LxiZZ7OjbFq+kX2F+cdq8R4Axe6OmMnB2t7e9X4F5qYjSPwfbWZJv9seK/yjBvpiLoB0qajDhUX
C2lt05dFpyGLs6v0u852Zv44scjFDb4ApPH7uHezLLLQMK3/DcS5Dsoz4kMfRcs+mfEPphVnLuV6
9Z6kq7POVY2LT26R+XQOn2rTm0og8ZJctgMRxSphddMJRbKHtES0PyU6V/zsHu2MExr73JXuhalW
AzjiK8WZHeflkg5ymuhfZ1p+pQFEP7BJvAGSRBRCAgrddhiX80UIb5j0neqF94CpJzch9PutMNWq
EHlkp+nfMHQf7FVcSo2RtvG8jHL7ceyupEGsmgqkrgPJRHVLHEhvSi1Sr6BTQ0FhGFEVFfBX2fl5
1XCw6F215ZZyG/fFoq7k30QduGsQUi0EX1PW9jns6rTIVgmY+0rvmhfoA1pgm50p81ywQaxn+ttU
/tmYA07x+hCeO7tENGiihi8cGIpFvXCUAIYy9XAWGVyA4yExRsoSt+5TscWMzAI84TvGjXChdE8X
a17XW7KkIuy5e0XaY+xO3ZvaXnSPclsMmXixrXEoKz+FQKgToqxHshm8iLciRBddY3q6qOeLAquG
M4LNB75ChttVXx3sxgaEW4vkiaRnCobCnQH4lANGSNxC1mpWScIAkZW3T08i1OXs3nt9mHr+GC7o
+giNzAZs1Pk1juhU8s1zijWRco7UyjXgQSv4RKM3S7dwzSrodEEMK5/BuTRxTbIJBNLZdK6vPToi
R2jccdYQJa1Hi2vu6GsJQz5phy41+M0YAHT7FJJfTpOPd6KM7gBEs529ci5d0u0oUBXvh38yBMGb
y6Kh6YE2Eb73TW+sQuQsvTB9US8RIps1ZtTIk0BYlsFyGZoNmUSmWyUAGVX74XvX5esk/3peL3M4
NPjCR6i1wb4qYf/DsCrw1DTnPDph4bIqyZOqxXKd/iwKpcRcqcDWs73ttW9DrTNqBV3MlM3Ijoxz
Otlsw7uUFCk4SFzHm/i7fpfBfHUbGIiCp3TYMdA+ferymIFKplQokLFloSHwhBScgZ80k3/l1EPg
BG99nY+Zcd966BQLYaoR8VFbPWPVRJAvYEpmzAdg9yAxNN5qW4tK261fMJJSqHVDD6pY0sErRpGp
jLrBygeMRqlhmaBW5rRf20szZR7IXHchq5UoWpOA+bOlxGTCRLNf+UQh8qavprfChp28ucH7W9aD
4N/P6PX2PJrk2KEbAWLh3cHQqOiWuDl1CaidbNibT4JuAEM7WgUS0EDEfoi7N+7u2mFZVJGLhe8+
lka4VkXA3gbLzpp9jzQwl5by9nR3G1aWSNncP109Tu0BH9MCDVN4MkpjVAmCE6Ue1QBMm2lRccgq
IolLO1a/MBVQfuw4uznFmrWsCsTg3dM2f6Z0/ri2T9VBgGX8W8vLil6DWK3IHQt9rkcnZHUyebhI
K+eMVSKjxhwjPptr8+ytEnlQmakJgK95ZSvpFf1nbRDDyH9XvrDWvmAKiRGNwrwXIjW7+FP7lNfv
Qz/aseNcmIdZxUEkPTphQjsYwGEjqj538MyydvztrfkCD/6MBlppwFBLhacwVaPzdsQSvhspLBVS
2sJfUTlTnpzPM/GgX7aQFqZmACLiUZHCI7K3Tg4QP+obWGd9O8pvE10g2zapatbbNe8Kc2ECak3F
pdjpHBlQucM6f4CTdsms2t7wFXG8diOMOsgxprmm4vAxhcbfEMGcRSbq3J2LHEyu5ty7XgdsDeEK
PeytwMWn/lOi2sFddVOkroTZTYfDW8mPDONHdQXbelAddsSgg/QS2e0RgmXZSmavkQ70QWY3gMrw
KN8/QwGpv4y0rl4jJCfFgoyqwE9nuenDyT8MWzPvI2Qa8pkn5lFL0NJ/GLA5D1rJ+GFanxR1gNLS
YvFN3BUyIoI96pWhuAPHbX4eH992nu5E5/DnSCZXgjv53Rz19XPszmSuijwikHauxF6qs1YTusH4
ES/gwe27OTQCxBwn0y5trPv6j9PUR/PssC0uk3ujZBPI7ayLvrU74oAjAU+/O5QVihps2fOcJCQF
QDka78gUNW8UOra6ptCmMRXqgekZ6gp7VbWoqYl/0xC8zuq5dH5AC/5nr/63JCI3d5tCry/T0pKM
rLkuaE9Ep+QmC7zZQrkVYDUfh49x7aWNRL/bhKoXQcXA/bM/0BqEIOHB/MQEjdlRoP8p48jbVPAi
SvMzykGQ2W1oFqNBDr+lA3B84sxM+DDIUvbbs3eqY2MT/jHv6Qm4GyGp9sJi7ZNgySLG7AxJNq4g
GI2cHY3y9e94JN0jkn2FOIjCVTM4+Ts3viJfhrvSGvPWZ0jbIPUiSKk9X0pvCUpDlEYv+xiA5Efi
vUVeAG2Ab2ZfJyIft8J3eJEV/5eapai3eNCdMLssj8GnQmZQM9JXISoS2vqymmJZ0e9cQsk8RgKT
dO65vf5dxBJQAWbiBeaj+7cIwHvbVv/ILfnZvFxHr+rHgegU+WgQkvNkXtMCblQFW8kGLtRC1bGJ
hTvwlQw6qHo8qfS5namop2i6Wqq3dBLFlhuaLx0sdCuZaXmbO8skjIun7H/UtUcC3GamauUBkcMi
4phcnwzGcIQjHrhUtVeKugqg+49VF8WuwSJ92VoOniCx0YEVBxz1TUsYkU8LvRhh/4FsXIIkLZHn
GOG3vVVAHlh9yFCW3QDduWnAkbD5nkQO/9zG+KZ77OQyx4Od/GHh3VWk6lU0QsXU8mZNk3b1zTkO
wgtEnmaKXgh4RBp7qpT4jFSBdyO0fhuPi7gRACqv8z7gDlec0F8ewDSYPSfioxyKZ3gdcOExmc6A
fjNxU1r4NBz+/Th/kew9gIt4Kg5Ce4/iDsAkrO/fxSRlXJCrMfu+Y2XM39Q6m6EeX+Kfml9pUii4
NETaZTpLZg+TL0njNDRzorDAk/g34pmzQ2P11A+gE0b1M2evw1RMlYCk9IMJ8howhBuiIlaLSnIY
HepOKCta4AKBRypnAGYnTJM0VTPkcUNasAkkl8LQmhLka3r+qALtkuGdEbNvPbvSBLBd27OHyGmn
MK0MvclTZwGMd3c7uQaw5PPGqq9J2JA/CT7aggLmWfj4VPQ3nlI3z1wilvoNEOihWMJTBszZ8o/D
NJB4E1HM6TzKOYRLqZDf5eba3ZA2PcPwuRUwkMGP9prs8Myj4NbYm6wcMa4zbj2TgIULWy02JQ4l
IOpkzNCIbiH4oPCW0oM40zVTWG8WLFr/SiiDVTzJ01GqOpRb/uTmXGKqV/KRnwByBtyBIokcUe0W
12QDjJjBSGbadTyuiHYY6ccJ9fyyQKFdelHx/czsIP/xgk2QJTcAN8r8DBweZGqpwuoYBofup/mw
pcz1zIfYRWfXQ5Wnn/Zek8y/VnngUW0zZOmLo05XJkYIUXt0R6VPVHKgvqnUNIFf6NPRH7aMLZYp
kFSI1WKRUA0NMRpCfvjt6PWo2+wzQik1XJ6UR14PnXVf1SrTRPTeV8HKslrtnWt0LaFDtdvKgKYe
SjqOI9gxJhLRegEKZ7vR5xGm1T9cCTUfyWsmRpbkhgx62AS4ITPfnIfV+YVf2ALz8YjJq0xZzoU6
ipG+4NauC8fO3LFa2RhpYCi2igeB0RaHk5+POquPIu2YNBUany3ZFqHSDpZDM9USIOds3j45ku8+
sdRN/ejgchzMGKO5Un3V57TYtRMsxOs1JPyhv3pVjpiKEYZSFkI+IIP56byfGCBoay39fLz8+NJ7
4pf2VmaqBPD2VU28Up6rb2p+kBRImeu2skujeDyc0zeg5RnmOM80qLpBhG3IMazKe1CbCbEmPPou
PlfELhGkcZab8TKOC8HbHlpagOEbNan0wptamT4joVBsFOZn/Emjon4v7Q/C05IU5cpJ/aOMlZr1
nOboWmY9wYmehCuGFl1Do2Rc9Xtvb1Htw+k/bW76cvbqzdQkEe6QoOKaFoQDCmOsz8OiB7tNoQld
/Qtjhx3g+anwTPl+bKdbxURz/jLRniRvVAQgwMVEVa6xjGF88E9nMkMPy/yw952RbjR87TqLhDGx
YZrOE7h0BoTJ223E50XWS0Pu3ODpmYHcPDFPGQOQs2lFYkh3P6y78qSrYPqNIQ06b47UWL+iatYP
qN5c4Vjo/m+8hGK/YrNzQT5Z/xUahDPQqEhL5k0N8xAE0qd6sA9fnS5sZ0pVsR33TSswUseyAU8+
ah1YR/NWC5qxwlNShk5WSbGW8eJjHreW6YRN2E+bN31k3YkDIpMwH4ZcPmujH94OxN9R0SgrHxVT
bLl+kDD6hSSAXkdG9ekR61cXNqJMrw15kA1sVXja53NbsUzv/ySP7rIstKvJuz7DWraG2OhXtijM
pQ0ANBSNs3gMakPP/Z9VXzG0toEx7iiLfWqZWK04t3aqKbQ6m59F3KXc4/dhnHzJBQW+StVsUWb3
vpFmrwl/GjmaN7xcFbBhZLX/+bjLCJG4+jefqDKi2AQe0/EVIuOUDXLhuxdHhVHkXuXmtD3EFSmp
kD+T+PmVco8oJ66xmmVfC2JCMq6jpVwsvParL0/L30qqrjMj6Qd7wkj/5Q3ZivgO2U/joevFFiH2
OVuCs5FwwpT1WNT2w2SyXfgBS3JTiSZHkQuFshMdzcz5K37UVok9GHzeEZ4r6NWQWNSXl9KayC4F
6+Rd7wQ0Ys4pAGg0pcSuEJMWcYnb3AJ8jK7Hk2T9EwnsE0k8Ey/MH0wlWfCF1CSibv4znDbVQfP3
zANfaPFjdCn9uddJsmZnpW1aKRPHez3gIUpC2FdiUgJQjZM2wJeuVW5FKh3fitvpzgDXGDVg7v0m
r1KBrZ4O3yjhZ1n53Ow1e957VxeuVpPvND9iBW0rTI5XhkuCYM/JwdSvhLWqbhHdX5OxHIGepiZw
NMpBznVHc5BPcA5XqnsGufyR3SqF3Kw5BjUkETBIweMIBNvQKhqqIJT3raE7fx7iGrH8dXu8UiSS
T0LtgoJsDU7CMC2lc3DLZROvahn0EEJSUK1qzc8U/1H0CkY02NUSzuu0AVWLP8a2kJGoi6FB/l7Y
XuWXf5Km6kJ9ysSLS6WLGSvBVHkjZLQ8RINeYVIgUDTEH+6FWoBiSz9SsWL+6W+U6MQLkz1Tqn2s
eXOlZqHVy9mzZtphBHNFsH3V038TgUMJ36rIPMA6OtXy6LQsX1ZVnYsxsUEoHD3thwPW656qLUkx
SLSpdZUKotukwme4H+6yEQ6Bb+ZvlZPAdIoe5/UEHoVdor8OCUp4qU/TuXLFxNwK4aRObbH+tBbA
fRy6YvecgENNkECptITFeButpwTPadV+1x+FlIZs9T6M+yHg7ugaTFHm2sO3MrdIBdOiFIvh0r/1
KhKhskSxgxHiMihgaRPL/O/IvYBr193xpD1wghMhAC0RBdEnsPMp4J/pasbNSANrArJJWI5lpKAB
q7cITkRB6WyWinzg7+JkE5+RHYix32ha1CDSJzi2yhARZd/ovsijihCSkW2npcDp3hzNjNE1v+JX
whufWrsjDgz2l8d81B3iz9oAtxgJlLZGbtWUrBItohkouKminc0vb9PVlF9F//tflhNGXcz0K5SV
EZrARF0qLdtHZ6ya9r7B0Cijx40qLkysYv80jIs1AXuad3kXxDx3beUO2l5Ze1NdTFWuTlEHfCb3
9tcLZazGxNQnWXMqCk6xA2F5EmRhFc4mlMDL8EzWQNNLXOh3L1iu7P1zY9JX9vNdIoRCMZi9viVY
s05MmdApU3AH7dc8swjO1Lnjg8Lz2nbfWxgdjOD6Zv8arpHJMqfrGGNPMumx+Brc8A6aOsIcQPJp
V6E/QU32eeZnCZV86EyKLy7gD79leolzFESYbr/Bu49cTBloWsGRVjkVQLKn/fadkUEQ/wkzs16W
pzm8fnvK5j9Umq7UdyKEph+zFzqUtuFn4vYLtWPycmmzrtDg8nOIp5Qc2NchbLcl7pEXeXFfrBmg
ovz4b+rMHRZsWpcfIoxqUYGPuZpCD5tgDOcKSGmmNtGksiIcZ6TZrLx2mPy7AnaaPQEIMdNPu+Qt
/nsBblP0X9lKwGmQcKBMDuS3hS8ywXMDBiFutup25H4fTqBxD/stCKGwOQ+GyyKDuY9J/2eA29Lj
/cRNO44Fm9fhqyJVvfJZR1iyYFGg512dvHlutf2ytVUoVfsL4Y3IWPb1XixEMMDpg5ILFzMhx7af
VOfVRk004yX1PN8E9GE9gOJduly225liYDWq+3TPmsqQXzLz6BUZ+WaUeHePbrx/8pfhHDUPcz4p
leyInbxq6a4LTWxmln+D1rGQNV8NQ75UYctAg5mNcp9N3ydFmCDc54PrQ1r83G4ZaOLZFjbsCGRs
roXA+tTo90CRdtRnit8ddYLX6CeRo6GeOEWDZfqOYTFkMgULa5uE1GQEM3qvzsgD4Ul2B3by7+lo
9vEVpgMWnoL5FQyZkB1Y+Osoa57Weup4uj3U6sMouRQiCxTdZb3qLHimrF3tcdZP8E2ISaa5H5Jw
hsRm8WoMSF0YUYUE7JHf6oAx4O7cmh0d7zYMsKCdswO4A25bmxYMptFibSCCcgpMxuVoB7SPob2R
IL4nDwr428Mz+hsdaZ1/QX2WL11ETN0Fp5Mr5ckXOP0Cf3hLdBVTbFLPvHclDOkSrJ8b4GO5zsbq
GKfpC6fU8CFkUQ9N+Ao8FM588EzJFdMxeYFtMtqIIy9N18ObQI8IOvxHnWC/RuGolF02IVWtgXXt
y9Kxv5OM4xrD3LSbphULbPnWTl+bvNjZNxWG3PZWlfdGi9TyeCi5bXm+FvGGxA5T2YGnZNa+hXDG
jk7nckBVTcapYHwPix/S43WY1gAE8r8SQyy0ROwyEbB4Dn3nFDVwgRbUD9RmEw5zhQk1nuseVRbH
VQ2Y7GtBmOGz/Tv1I7eFJszrWu7tgyQYLhKtiDusECOUasjqf8Ti0sFf+YJkOTrM+gnvxJsNXMCD
TWZQoJXjvzTTGH07PqYesj2JpT3bO3SQ0iQ2/0o8MIYb2ClfcbKRuCMXwpf7nogco8UufbeD11v+
ZeWm2YycESVeOCaBtJI23jC2Q7kgUzpNP1DKPVdjvrm4/7KWxUhdYPndJdPAzmHboIpLQaX91v7J
Tq7HQb/j2wGKjutIf9bTMFJ1y6pIj3FE4OLouBxqeEh26ZIdwYO9QJ5kbYZMUue2Hh8wk0i0aW1/
nBmgFeYSOrIw0mgHW5xRTgKpETsSl61fv8yI0GhS2ptcoFpKytrCMiOlVA1bohw6pVNHagw5b2zw
ob7m1iAxvox29G8Uvml1uLg5wYpMhE4l3cVR0m8jaGHPa8qvvyJEFk2NdIVOfwX7ysgWfXKsJJcF
84NwJ4r7DZisaZbnOKWh5CJjGciRzyA9ywYHNJELsmlM2Zur0KmDGtcN49oG52NGJs7JGMgrUUpc
9eJ1RhFS29JuOez6p73nFyVoJoCOdH/7I5Yts2+/29JDY3QUJ850573vtk5nNPVPw0C7A1alUWJ0
brtZerTFAnJaCHt3fJ5JB8dfhjg98HBlPEF9Pcpp1xQB4slZk6q81ME4V1okZsy+WDuBVwpb0W0K
eQLpBlqWKlPSJ8Eho4iT/UlBd+etN4TwjHPZLv+pcFEs8NIUOTMIQNkIuSUcAZC11XnREm37C/S8
49SFgjHW78DvFiA2GMCaHoqd9l4VzD+iCdlsj30JemZKBW0gKlP8jAS3ju23L8UOQPG7upWCMYcV
tjo8YI9O3g8XTnm175yUL0bp6OQ/4wiMaHr+57ePSRlZkpD4LvdV/z8f6gr1jbO//YRAfvDtgn2q
TdhUBjdycv7I8T02NDSiyFPIwS6iteTzjmUp3RfU8GJqdxTo8f6pPo9s9ANvVtUU2bgi5NU8No+q
kIANtXrpgsIWzZCKMYwckNf89mGKZktUmzEcBlmpJPv1kLEpUcYc47v9tkfbIcGcP+M+UzuSgAY4
KLvFzEdeJOKdwH/NsBNFBS0uC+KZXJSpdp7JzlXtM+iqJBeNUGsYKIozVDseMECkJckYi97Xc5ij
x8wzFRNw/D/qKJNsMa/uSr4kKQVjFPOColo0eJn1YPyPSoWR40Oftnp+atpaLjD4T2muxD2O2UXJ
xBfCq1UYPIs0/1iWrEHdn0q0CsSXlhOqElhJ4fGMb2bsmSznIPFrV0f5u/z3mzuwy9ol4t815QXx
xZOf8p3lZp4oz55NOQJskDssZCoOtnMBnOj0nOzAllEzEF6hr8+qbo17QMqw/5mnLRQptjqUaZqT
cxRSpOkprEwuuCM3ynfdPcoTNgvVHb/LqoYVtQcyt5FcTpAZDd9gKherL7w5B7KvDHb+HmMNtPqe
x4QtLjMjhZcuTu7a8ruU4PIVtJLKOtY4+h6p+00VmNSA//Li2H9kkusjDSWklUsSwIr4lGOXIKrx
7eXSH0F3x09sCgvSeVKzHQ8fYYwbRXJC3nUZHV1LH0+Yv5XMArzu/5CJEjmlaYINAUgk/qytjoWq
f1wqMXPbytWdmVvs3FwXj9CkBMWVA8gNspAftqecL8cogcfRwoIEBx+sUhA1tIIAIhHsXVZgSxDV
l/i8iUl4WIm9crE2O9pEyXyWB7dcyE+6ThhjhpEuB6C6WQ/9F7W85z6or30R60H2JkfVSQQj2XL/
f+O6iE4pVHfH8yRFgC0I24gjNJ8L7wy6R5CItKDZjPizE6Z4ocwQs/i6AponXGeS+6ahGyOfdUVE
+i3M0vJbU5dGKtOfdkLWfoyb+O4fodqGBDBXFkZb3l7OiRhpo4dSBAW73pe2qmgYt3pEU7EMt5N7
RIcyALpwB3PJkKdtSK4Pd2EGLmH2BlAdzNbXhCDP13LTE3K76JB0cOOaHeLdpF9DdyvLEode9CRu
nFSPgo7dpbPDeIg9Nm7H9sfJcXpjfmRsc3PP4q10ePa7RHCdOI+MDMmIOChHgl0FBW2LWzWWEwpw
9YCjER1fmiI7Wp326HDnUvOKWaS0UFJq/9YMKv50Xv2m7VVEwu+tqoTCQm97eFI/3uwow7yA/KB6
zOiQuQ9plxhYjR9jGRtnBtrPVo1ZX8wEvKEY7U4BNjrk65Op362mhtSWZckZPjjF6n+S1nv5AWWW
VSfZQLzqzzQ6VhmMXsLKpoZh3gCfHC29opbIC6BpzXm6yuJ8ZGix3MkDuKdjpr91q/OlZR1erbT2
LvuVcVHfsDK19/HumW21RQb38/YO0AwF6AXIS8aKjQrg27CxQB5qKigMLYfqgOE2jGTopK/hxMx1
1+4kY2bzGMcWgEy4FBKGRxYF5noAkl2odFBmzfnrIhcpHw6jwT6W7a3E4Jk4Iev6ihh0Wl7KdE3S
T5TZeNrwwx+ujYlCBqLPbMgSuTK3tDWdZkbg31qw1Osj+vAZ7VRSosOk+bfWSfwOg31TZQVX8umf
FprO6p4N/rC0seUdn2JaGfPMPpM3rDAiDFqGKnPOSirNFkp4qWebXQQ9ioSB9QD1TFGqX65EcJhZ
j8YF8Ma4VK4/w+1kPgQ2i1ZooxaS9dzgeL3j8mo7X8Tvslz8X5v51GiLCuX+uWMSR6eg7XwXCZaN
fJ1sTts1KmsznmGqzpj+Uq+XpXHuiHeEFBXJFLKnDFrWacnbn2x4JGog/NDpYRKXbyoZ+Ay6Z9sW
bswMd3ok53bZ06jGOzUJjoWt2hALjtDlDH/wPubhk8MKbZScKfRDW/JqEXuMlNUKuOXxJl5Xaiiq
NugaHiI5m1gt6VoF8iGsXovfVcd5zwx9kjak3UeckdQBvstyALXIRKbPePcga/I/lfFL/eLJYOl2
IUPK0cfezAtfLCvn6E9Va2uTrvBvb9AJAvyrQLa1RXzeYFaYhe3OpTg94LCFjW8Gk7X+qP4v0vB1
WYZJlCxDzqwf6wVgdh8PJUMpcc2+/3wCdxe/YzbNuNDMb78AG5xLFjvY2cO835o8Rfo9ramFhBsv
+P58QZbv8VCaczDrb4j990A1dzNl84EtY6ARgFJ/UGWtXX3ZLZawfjQdGQ1dZxhlolYxdRTFJ3bv
sQQIaVMNWONF6FEnABg3dmHxm1dzl+QbeWLcxDeEm3FQu+F8a6KvE6ItZV9zXCtMDJj9lzCQ9VGP
LYYywRlmVUM4TpuPidC3vbLhYsBURiPr/HdaCUq9E1I4lW1Sn8SSgJxHOfCOB9zMJZn2KVa/fbSd
aheR6o1DWcOXb6WsWgCqqKHDVomGJZngoOx1oaVbA5IHl3iIpnRnBoq/ncAd9nL25DRbWwuXZf/0
i3CLmgQDzjNK8wplAmoM0N6rp3mh92z8ew6NMVivuYIambKeQGq+UUAE+QbOkoe/Xjg5R8xqBg9u
qq1jL6kMM9ATZfY2mXbmqv2UfeC9hNcfQv0yHWs9zcd5If+INzNGXS5geTtUlIcjOTo2/6L7vi55
uqt1h7LK3mnsD7cE9smEIg7LDD4HZu+R0d2xuaFJ+f9LpmCpWNlNPMOeoDNLwir26XtUBgsMJp/5
mehBeWWcXK7sghHcadiMFqwZvuaApnugIZMUIKp4nWI4MKsRZ037ziOYbQ/HRUK39N9vRgCfhlOG
bsZspClyKTf/3QoRgKfb8onLjQyM7muN8ZwIKe4AoyN7y5DGn1C79rQ9Y9Xludo0z7vb8xTo2teY
mrmTcod5xrdvVyeRegy4ii9KnYfSTsj4fMnDuw6YfzAkRY2JEbFkX5HQ5OGo8RiyXL7uP+LpMddj
Ew0UYH/r9egKO1rf+r8/On96bxacyy0GXHg1SUIt1yMOo5P1/nTaWhLJAS+QvDXbhvsupgQXMdLB
BeMC/+L7NtQ0x8iK6CbisY9GMuKp++ed2vRcW03w8jPXvQwY9kJnbcFnXkrQxBWKFuRCz7wD1zMX
8uGaojPu8EvedQoa2G7P9428rPbV6JFNO1qWPFtbrv2gPm5iXKb3AiHeaojXnrKGXg3Xwt1+R3ov
tX1qAF2YDV9G3KpKVeg1b/SppY58von4MtZHyGctADs23oURZVe9RwYgxEMcBIqJ2Y4wHh3CfR1A
L6CxCli5qngLo4Xf5tTlVCU66/mQHqmjDlJ85mssvWrmPGVBXa/5a1AnOzzDE7yIW9Y6OGVhgi62
ObHAVNPrifMXVjgXPq9q5AXZ1wca1zUS1JITxTVrLj7zJv4TTynJvWep1jRX6OtkQ67SS1CN/3uP
gq1qzIo6m5q9zjM2RdFqrR5ZRmJIY7bS+dDCNgNXsnxFt2hkyx22HxE5+3XS3aLtPQYMMe9opGw4
SrhZTmRK94m0zfirfEawDnrqM88ZpqqcaxQ0KW3PTMiRHvmJ+lCgtOrz9msERDjRLchTmVQ21YyR
fcQ4LYB/zmiNAX5gSV0ZvlCDX4fVw9rueYfTHRaBsoUhKMXzpGkyyQB0MWD0MmOUrv9PxjJMjHdU
QxtdA11WnUNbUdUaIft4uHCkMm+iZxToKpi8URru11C/826l/Yihxsxq/Kz4+v7UEt47U2jMxSq4
xLxlVe7JT62M6CoRVbHC9m3xB/7wuSHwS3jkQLeyzdBIv0ru5vkBPpKHElPUB/z4FjXZ6To6hoVx
jLLai/2KBx70J0taHKEQqBkI6QWF4M+pzVVqxwDFAe5tJ1iyKUDoT9ZyTQbvMHHxCPJzBCzhiGyD
QgYcBOixsqxeAeG8RtnSOZp9T2kOWe+AKrQcCNiYQCBPSQ8ngs3p4qzs6GQzy5ZjKatyTTUo1knN
nDfrjMEdL/660Avtqd9S1MQv35EIu6HfzONWFNkDYH7khV041Qb4POctTBoNwNDk4BfxP/2qS2Z4
qGVkVbdpxBYnca3leeRbO5agueooa/HaD0l9HGrmYLPr/SLqreQnd0KKhglOe8wf+zSOztLI958s
i87aMacfXbhD1lkiAIpkt6mVbl2yylz2N1iXGCLvdOZwJz12yn7DufmWwjAvIGd0ZOhyEZ0Iw6YR
AtznY4gi1nONScCfp0BpoJOfBLCxCeFAbUmaotV22ID8iYOjVvMYnZ6sTHcmRiqC03xn90zBl/hT
IzSQ/Esrr8dM4q0x198DDv9e3ooABUOv9XR12L8IpmcfsM3bh0UyFTwzG49t48vjopr3VkFcHf71
LEdLPvVO6LtY7XtiFZtkYUhZvFmdi2DSwX/iH5pvrO5H0XXxMQlDHmceecyGCWWtsd+NLWRG7afu
DPd8q29sEUb770gXIW8btFxDENqo+btBTCp1kI7vFf4Fng53mj+sIyaulFZZb9aNjVBBu7WJHcZ1
m/CxwY36ix2kf+lECPbDkaqWuMv/BkKGqglV3g4329Dl1VTr6XvSsjxw/0zb2sSSA2nDWV26qsOV
Arpca+bCjRONz5LGMqObS+rnDWNGFJ7Y8hAXmU5pspEoIsEGlpvi+TPGrFCjc3yG/g9Gl9X92psB
8DimZoCOHWCvbi1oZHmBv+xe5uG+hA05x9BHbJ2Op9vQgxVnGj7IRtKC6vJoMMxuxSvtxZ81SXCo
z+4fg+YS9VTtjm179W/IZnYwAwyaEXIN1sx7T++lbqQSAqKHRNmhg1mCGWjBa/Bieawqqca1k9Gg
PCaIka1H4/dR4qej95VxJQC8wFCgxVKy7Z9B1ms5OBMCJYYQ+CFywyPjwtzuXqHX5hMcsfmqVYM9
+V7IPCDCCxw1D5lCK7KrJNIsCCBvpLixao+cihRmC4c529VW1vht6Q3w1Dukx1o127ZhQijnQ1li
VpYafj4dY2gb+Rq9Adl3gwAKdNbyXrU5n8xgOPIa8OpEvHNvVt41/FzFns2I3+NcM68eGUyt7LWC
ZA4R5Tq7PDleSv2r5GnmDnPSQRsK9DrvSstj/KflKXAJ5iFijaXuJEAgWKKSusYoYv+KGrnGlpQk
UAMpspRSg2+14fG1LhaUxBneazie09eEySD4kvVtWHEjKNE7fvbKtzTzaoD6NZt1onOcIpsi/Rbz
FyWiQGiKyhUMBC4RmOXv9nNURtnWefXwZdVCldkBjjdz3aGs13Pl7lQlukGKqVopufSgTaZuBgLH
AF9hv7Xg9P3484tAF5rEG2NCxwF4H2Im2HogWxuezlsyqj41FmPWxOcVG8Iwkj4jiB5yQejEnoxs
Wp4iF5Pndp7k974/gY26+VMuSTyN+mHUqn3T+aPvtkA+TZLtTgnqCfoQu+nw5YzFBkXst6kBNflJ
qlfFMxSv0W+wBbsb4DoshjGR7JYAWBuehxI64r5aIDv/6wgKp6O9cwbWJOTmJU90J+PayvbkHqUc
JrH8iV1W20w7i0xjWLXQHoHd+IaPuZHBsENJrJVElpAKttVrFextOnOBmF6DUcMeHEEdj58qxUao
ogqtNHX/lrVQXINvtyl0y44087+5l2CF7RA3mRSX3AZPRZhlJW1voi6T9fmIV2Cy/ZxDMAwop0wn
VEAiw3tDDFFBOncqGp6jqtXBJgxT0gwiS4jAPyYxfyse+Ve15caBpB6lnOWdSpyGOEUOYz2EfFl7
jKCSnpC4aW/OWSPplRukp2xc97M5ve+ogCVStjbfs0oN5bJGW6pLzSSsolVV5VWT/vBLqgXxwIiQ
ZPahoICNuskFvm8M4mZnZMPE5bCkN46b4RAbx/4U2cCTBRuDCGS/2uLHynlv8qq7CX00EgTrOFsL
+bdbD/84JPmHjwAOoPzHtzAGTCUqlPPre2GFnkWwXUSMQBsuvw6ZBvSXI7+rE0aed9CwhMx7pxDW
Lcvs8fJ4cf8uFf2PTal9bV1WF6LfTTHJX3bx+s3ZkE2D2I5L5S96Ry1u4OtHX29bxFfvWCHdYVWR
TAJl04IliXwONPISsuplWT2mdiAQi/c1rrwf7smYVlYOmLCXbXkpatGQC2z6yaicgZSnsqwBgwK7
Z2Fu/SQnv1+xCMA1N2WSyyS1qfBSDC8M5Qr1puXYG9pl29DPsXKpIIDBrTKLyLwMPUL0F78FOKn7
X8O5+0H4PsX7o6szM2Tljs8ICDR1xTIo4F9z6P1qzD3aU4wPzT8/DfRhcn/qnyzHv6Ps8NzhG0yI
m+TVywl2Af8Jo+B/cgn8R1TMBnfkfP+YUjENSkRXjiO6Ex3EKaxxA/o46GPvQUsp7BIsADLUxtk0
T5ONMciQjo5oISMBqoO+/LhIHfVPU5z7d1LEvWfdLTfeDLaNTmMJ+Ws2fUeRgrkL1d4nfyWkP/5q
O4LAdbaJgUdNJzhlak7o0rYa5EZgNoO5fxKUlJPj+ZxM9iKy+0fc5TO0hUygd4omukHqIRf59Kn/
RzGsTcrln4s0VxSe4Mco8heLHk1IzFLnDPbH/PAk/gHW6NHHKx0/rD6eWTCpK+LaCUyr+w4bbYyM
mVbTINknhWYHaoK5EU06NALx+q8ma8oY+fu73QLGXAxk2RxgqGBYgjqFIxoBuErFG/9KFgXUcpdA
YQoG2rgUHpid97sJUAfn2rQtHz46Xxn2WFd46FzVQas31UzYb0nZi3VMiRS2qkkVLhyV3VKQ7FUu
O/9MwNXCCpz6+190Y65a67yqxoo6sShzoABzyh+zfekvmrVkUUN+NkUrgVxRtZtHkPoz6e/OyuOz
3M7RXU1NC0Ce7/J+YVhQ3LUt824x7qBrd2m8AGyTcUES+Ym/9mXEJAdAzm5Wuh0sfXwoTQ8sWxmm
GjSw8Z9kOXEiru0ZEwp9I7aNIK3x56qKrgJWZR9JZXOVFgMOjy8cafc4MQ4yHyq7Ww/BRGNfl1BR
aA4s98I0gAHpCpIlXO0gLVsDcy/AAmirf6rHhn0bBc5Jq7KWE1XNOpOr2mXgldMUyoQBXfH9xvUn
Q4KDx4QmTsVa24rRCh5JAb0Zx2fZnKJPgXs9nptSI9/rUo10uaWQ/sUYZyT4QZAjcQhZtFfmnBrK
vYg4uNEROXlCbRXOdoUihacur5D2nGnPK66N9j13Xr8Sht5IC0Rb6taEE+X7e6SsAEBCvGouxhVU
NzEsNo25qyD+WcCDZipQ50Y4HH20J7WGuzihJyOpaoiUi/zrfE6UgZk3sakg0eVextcv0roW3uH3
O8zipLzblAWukkddC6x34bZBl68MC4Cwxur6Bphx4LC9RfQk9le5Oq2a/ouOucVxPJS5633JYgTy
2DIqXoCW1jc90mvz8YWEGzKIWRoNKUZe/Q06trXFJH5srFzoNN8/HaIEARQRVDcCg8iAoaGdycXY
7zV1xcWwwClKHfREofRFpOWj0Z44bc69GB1yxfDslGG2XcaThwVg30uHOdwvGe5fpOgQItVzRhpo
7Yac62t+A7AySDr1SIQ5m1xE4svdNpUFvtZb9QHy4LG4ljDO77c6pWQ/zHJ3DNO7kHVFZcGcFxqK
evtrZg+aGVYb2ZCxZJkcngtz/W6LcJTY53RLncTmNGP8fHH07HS3Cb6osQFGANrdNQDPy3zCI4Pm
gH7+AdR8KH779GDfu94ByQDU1g8qzu0DIN8e7Z1OaosyopsdmW/DtwYHXa574jsVS95GEZBD+CTt
nuyTrCdR2OJjdNMlNXo4ATclqFeBjfMtUoMlVRL5NmDL/78KtYx42OL3Wkaovur5pikioiJ+C9fb
BGZWtXW+yqND3la9NjM4sLmyu/YX/4CMFRBeZQmoh/9g8ZMOTbq8wXXytytiW7pTINhxHuo2YM6u
GnuZxw8GhZxlmHUi7J7m97yKbf0PiXlmQQLaKx0OVY5F3GjW2WGe07xysHCAIkecYIeR1RCYpvlO
q//nzHMTpCwHIwoGbRFGtMDgDZcJr6ftFPGIubk41M3KVq7GooacRPxJf1khXB0emLmKJ03Yvx5b
phNTHQRfljhFSHnSbRvyVdWKldyxHRxve+vz8YakyXVK0EyfI/8oFhFhr1rr1TA85UqbgmIQ2uHz
359Bs+k8z3qScHIPThwvVE0w/X0B8k/QoVHg7bb70d5A+NR6+RIPPY6ANOShXXXZ3eZLHcCZ0KCU
VqUVufFdjoplHRyq61+yRHczPrmkGmkiP4ctu8S80U5f+SylFWwVYzRszJzZkmVJWtKEKA2teNg6
T8VK3kZNbtfS1W9nLxxryKEg8Ns4dHXd4ihlkZmlw4QN4dGm/FccWK1JigwH47xEnD6BMct/mt/j
qyaFe09vrCMusgLLVapNl1lztE87EXtk5FkTADZVX/3ifawYG9a1b7cWENBZKuNdqY1yoZghrXVm
n8lRnynWQsE+Ebiol2xErc6iJYH8j6TeC4Th8/QHqIH5hviJeu34gxe0UpsHBZCOgmxcJLReOYMV
MlmykpiaJXFwTRlVEUWNgkPlrBpbtxZMqN4dXtQaOPxrXhNR8k8fiqyy8yPAG57+WMLAupMPwwTA
Uy16d14GHhcw8VtaZIzC/jhktAQwuMJKF90G2L23usDKTz48NddyhfH7ac7+EZjbLayHWBRZn1/r
LldPBGOnT1ULVra6tCPkwaP03siCmBV+2PBmdYXXHQAlOYN8rizS4d9KmSzrj+wCWJUnJ/J4uf3d
CozQx4B+4GP2A5evAqS60EoaMdU9jLpLDvOSyL7x3jGMy8f98ArlNNZI6J4nWCsfrBVmOsTLUUSl
1qDJMDomhXPUTtf2jIUwqMw0wBdlc0NMVIAcve49Fscm/+UT3tzzZ9AcQedPn2TTWZq+61SwpC+y
bTqVTRm5p8IZiBZXi7jY6z3RLqpceBbVXuq+Hb0hYT2OrcAR4gJJLBEElbQgjHtQ4CzkBx9tCFPS
mOGywUrxvqvqemeaEuBVjcvWZvEJnKqu2G1yZdveyzDcn4ImL6meIx/8aCpjVGH7n4LO8YdNK/o7
f8PjkfeajEQmbJ++NkaBnZn+hOOPocyairNq62MK79qWCzQEj3qLxetqyxmXoVqm8tMSOaogUGnw
gXK6kw9ZC/Lyk7wv2H5lEIl8cWwqLru581rVGcy5PX1CFp/v0+rQ20FRULCEE+4FYefSVBG/yuER
IVQeQPXoL1E1qmAqYdrS+bbXl/M63Wcco25ZZo0+hwWnWeZLGxLmWGc+WZ0hvHnbKqYYnf79BQzI
C0wNaZLNSV7jdLUsqbvM28T/Qgz+MczqSrNsiFeTARj51ZNwGX3Qdf7jE0xQJz48Syiqsi2Rmn42
Znjiu8y1arNjmbXMUirgnwW2icx2G0KH2KWkbc5U1shB3sSH4gG2UlFby7CpF6fXFeozxNS5JYk6
b8oudj7dRgo+OIZGndIC5QgzaYzdGSgUojlzBAhgnli73MHjbTixw7xb6hUCkFY136KKtQhroP/a
Jcyno+CwrLcyjJeGYSxcZn3WaM/6jtPnWesxKt60nJ5v19lBcv8XONwCcQY83RfikAGezS/+K5tS
PzTjTWZNB7RsQ0qfs+5gD3i84DnAs/iroXO/SKDgDheVkljvbbOMrJXAj2j71It37TIORw2u1BMo
nGjoiwegGQxyG4ktOgU9S5b1KWFME/RGNOPN/JY0rkBEzp+BK8QOa27Y9iS01dYWFOu1vZfAwy2F
uGeptizOu5xkhJHZxYAS0klpUg8ZpVa6zdMw0cm5kmqP9WGu3MiS6EbPUJOLWa5MJeftoT7yCom1
IicPcFzXBqClkJDVU6irLw0gYUF03a9AaCtx8guicxRIDPxPPhZRArDnu4pJinsujzeqBKkZk6hE
+Nykw+pJyge/NAgna8gwTxK3yJKYUXoYa7/YU/2O4dTlCaVaXXGZa+rntNqhxjJoEV/7Qeb6WbQV
li0jWCSvJMP5aVpWOYFlUXEOMiAPipecMPMT4BYQLLCJoRlSTqlh8DlmOuVpo9nTfjAkgXnmxPbZ
0f3Hf9gZiQ3dPNGnvpptO7CIV15DGhlT1ZFz7SXG+OzK4vxRhEpmlpuittFApjiB7LUtii/Gzfr8
8ag4d6e+Y9jYa80Sb2eAjevPVeQXl/7Bvz27FQXBmRB3ECpw61NppLbL2MmGArnX59ZzraHTP0k9
LpxnoEFtU8klmiWm3TTkGMaxK77A56T5LKhJH0EP+1tDZpy6UblRiQjn6RSwB7k1r3/itKnhWKF/
kSiD2c6A5i95dObakzgkyTuDTgPQ6ez9b42yonoQhk/4ao0iJaE6Y3FgHn0wDcWW1uJRQGk0Xefw
LZClxMiDa38nGmlgGe07sF12FdE2259B1ucbNna1Kaz9X7pyH/rtHeyhCozRf9yBJrpNvxVGpNQH
kmRU6sqUOw8+wy0rCbTKxqZMH8WWy3XuSdW+xAa+5gPDPGFixWMClRJ6mYvMdEyDhn58ukTIh+1c
IccXOKuure17C98gg+A7kbHoHhq5yQjj6x6/PWIH48qMVLPm5UuKmGT9GEo24MDxhAZlD4G/jQ38
HkgYZwUead5+gx5vwSWR7RMT4dCBaW03uhyhv7rTv9PTZV/ajvBOLsq6IlxZ0WNBmbpQQh+9DJ6x
fyVL0VAFyW/0lbC3DdKXaPysDqopGUOCiMAr3bCK4NC9lNq/1++2sLPy6LRNC1Rph30gbtjnNJ5n
GC5l/YyGXROkN3JxNXLEbEt7fQZL5DHHaEi+5Z1k76dAvFtqVrgRLPy8agjxbvIl9TW+19jLYlR9
tPgHacLqPT2wWypb2oQ1KKS9QS7uFf7WAFNYck2T/0CQGjveiMSfq2JjkwAFPnGSU9uXjljAxZu/
3gS9DVi4idGWk2ff4SxAFUK2OsM842wIWiZA+mj72r4DfGDPHV7+Fh46x752FYM1smvWHJzZID8e
l11rcSSG16NlDsZ6TBQ8dVpaEOQYS00m2nURl3NTAZS5IZVj76qKiNEfOp90H5Nch7/mYZKEWSKW
x9U+cG6McVxSns1ynb3PDu3whMJvWlSaVoBDcLG0l6x6p5zvPM61oc6+j9O+j2YTsJaZrKZlk5Xg
jq+c83qMENuHpIMVRn/YzT8yVB1Fvc+2AoP7ZZtvKD1R6k9TJlxbnaYkAWyA41UguyURUIdma2f1
PdnY6jmOdAmENwyWNb96tCP4NJQI4yWJanS0IlLUSH2QS9usK2GhNCuHygkCMi0kMTYkRcgTJK0B
P3h/csobQmYQNd5pzLm7pgkDc2077MeJqJuQOrRz/I7wzRr4prY00U7hkl+mJwt73pcFqZFt7ynJ
PrqwNeHAnWNAwMXnSirJwonMzgCI4+Pfd75vSaPVMHJk18HrZoSIGAIRg74nLUMyz05bcvPEwsB0
GBh6wnabMPB/GWxP4rz7zVuIeovkPyvVwKve1cbkWgZYSa3Iq4NV7DkPA1wOaOX8BtYyIk6BOSuS
cC6HHFBj9duUcRwnLB4O9+Hgyo3ClnVWjBlQDM2cWBb1LsolNMrD0GmSAcTH4midZSoIsYJh+p73
atTW50NYwLstFzyv9wr2cdzZF2ai0F+Ef3zfst1AeJcTUcInH3H+uQRUD4L11idDhusNWmqZcuwJ
0MVH25EWKEbLGEGWlBrXw6Jr950VBru11XfNTUEwJHfNGqjdLxm+imn/FihowGgoO/PJemTn1YKr
bIWVRJZQXPzwie5Dxpp13Q3UBsN7+UWralNQhABpLAoBZlJr4oNWq/xaAvRCVlOHBszZc9Oe+tJ5
3pDyrgIcfoOD4JT9zJQNHMaEw0bOis2AZRDOw+vqJLqCvUqwxneviKeb0R1pIj7rKnIsYw9El/Q1
GCOTsQFHyGLDPxtGAiUdHthQdHFjuNTWQyf+xn1XCagnQKeXvevTaJJbTY4JYcEZ70uJURFmBw4D
krBGBwXTdeZdKzX82xVpSs3aa5wSL7Ow6OCAH+zp1p2cSlPihzl/jwcV98OYA/ohw/jV7He3C0Uj
YqkAvSFJmPFUT8h2nsHAWXGNEvkAre3Yse41teOS/lRgWki3R3CObcjJEGfZNkYQ2zQFTZtgKG5D
CY7JRsI3oLFXvUj1PNS8fnM7P+SwtE57IpRx/OW6AfAf3gIDCyGf9VyKiFy8Kt6jaJLcXmGlkmUT
e2EGmBBwI+ojWQZiTZ17SLtF+evizC6nXeoNE3kSPtbMEWGQ8GoLiZqwT/NWcTANXcWAhLOh7La+
gbpwmKLoomdnNroE1mc22+UPoXj7IU9/udzQjo27ryUNtLjhhclQ7IVUkI4CdFhoIt1AeVtMl4AM
GmSfrQeFh1h/XvCsMHhdCCb2yBzWWTjxdRW9+7TrBV7qxLoJBvzNfvVt7AnM/v9aOPsAM9FA5Bmt
OhK4AR9yjqg87q1sGWYo23XsgPPYiKaQOOPkiBzsAMJJpyt3OGBsCREy0+d0sqXMmsdIPq/tz7cA
8WnhPtfHd2qHzFvMFyWK2Vf4CMKnaikfZgBHu0pVGAhrVH6fhpG7VncK/YE4hUwL7oYkjq1Zim82
ig0AVktW2h/GrlNR20NuFu4cBmiHTCDE74tiCaaZQg+h8wRxtPmiC3uiWgIP2RwJCGdw+++DMWqI
alAIbPHXMEYCLiwsr/qck7mkcg2NtJuqs8QhVx6144j1hw6709RojUBZLswOuNPdeVTYWwtrO3Er
LmDRKhjLfDvjX713rBSf2RzVLM9xvXr3yOP46kNT6ev4fORkB03fpYL0CVIREDfOQuO1mtIWbbvF
V/7+Hoim6AejMomtXv1WtgQ4f3MBYDC2nuPj94m5JuW5ks03EjvQ9194xlTpgtpQyGmydRH9NgEB
3j7n2qLfJlzhLV+z4Y8HdSzWRnVB1Vp6YZbbImt1ZUaFyP9/K/ZZ6rSDAPfqtvZ2R9yRYSqsUxNe
Ju8wY752+1oHMUujafnrh9qBZdmYVOO+8JEyQGcx+wrfV69ET36JMjlfAJueXNk2nNWkUvpv//6q
s3pRFkiesn3V6KFrC/ux27AVvjbApJvkBwmlB5lyw1NGPllj4Hg2WXOBXvR69fMlXxTB/rk4ZcH3
vzaLVMqyrPw1kt9gWztwv8FxK7h8ymNuLLVsChDJVOY3Q9RoU/aqytwe1P5pGg3fTIrDaETVRwB/
Hp2yRIoawjm9mrRXFzfhRYoA40ac9ugG6mjw/k4HWt8i4Aa4IXgGnQ7TXT+cUxuqfXM9h8BIzWdo
VNyzF+X/DB4xE2AylasDiZNI4U6lC0oW98H/fqRsGD72yZtHfPgZfUcvyhdcL+2xD68qDIuKOkzs
uQcZ/CCSGfvvyxGOxfQtvAmZqOMA2eEGpuXC/jhhZ7NeeZqt367UPbuSfOYOCmCi/dFW7Fqcj3ZG
M/LnayBz3x5pSGmEwV1YgI0DzpXJwze0CzCZcIwN9OkzsFtS7AJbAtL1J8qI3RIa3CdN+bsuX7YX
/f5/kt22eGqXdj6x+HxE32uXoaGHc2S2aMhd9MjCiPHdhRJOaGciGbZGQXNdJpOvdLe1lqt6FGOa
x/1Fp91DtMIke13NYsb323DLfFlnJJemKtSlTiAcmhrLlHu3z+JIWPPoqDy0YQSUPOcGpRcfC2ij
sYzm+fs/tnS0MEn1iw3F9DsvoTMMwSSqGAhmZwfccj5jbqRG7u+D/OEVmPhbnMjNiisnTbTlR98f
0i+dcOwQ0yzb/oHTn8lMCTNvgQoksWwrT+5mOK1XedAEnprOsSM/d58Shz0fPrpihWNlxeGMnrVB
HrMkInaUqsfWJyDLdpu7VjZqhjIgHI/ITyA2A2CBlCmhmMhKTeqaQNJKvU7cEQmOPnONVSjGbev1
AWnT+BwiPPFDGBdr/aVqbFNeEK6CZ4cDUgAuUOANXgYR31SAQgW8Qew5BkCWbAgaNmuoAfCoWB5y
tXBc2VO6bSwtuK7+clGB9FYlkfwC1CoM4OM6ryzLLH9QP+dVj6gu+bYUROR7MkllmqTEyN81RpcO
GO5rynQr9hO4djtx1OznRne5zZmCwcqBXohGwnmr9XPN6bVoAeKxoeIbwFZhRED9/febQLWu3Wfv
kbj6VBeMr+dYgT36DJzti2o510xK8bRF2LM+fJwgSa9XwwI6nGPOVO2XPVNfgKLX5aZOsb8xnRUo
5g5DUrTm7PWFOUjzibuqn5C022z6ZFNACP9IsYAH0xgDew0vuDSxFLL+jeC44xG3WQ7TYckhujHd
yFV089mSZ2CPpyyXBj8uteaDCnd96N9yKnVIHbBXmoq0zrcXL1NG0uPqSvXvNGggMoJ7Ow5jI6Kf
U/8i8LKRXKwPvsWIqiS/O5/lOE5gbZaHZyzSekw/4SVfTsR/ojo2z5uLJwov8kLdgKkiaa5mOxko
7wLQFfnyHtuR8RptpeUaInBH/oKeMnebTpWu2nqzNOiLV8GUOmVKM4IxLpgNCMVrRoiTGw4tTSP/
INxAqsUmfk60mpzgldtqKz/rmszwR3ehVTPQvICUiW6amLymrJ7fOKUdSWcyad7R4WkXH7g1nZd9
lxvPde3vFJXQuC8trndmYWagGMGjwCU4YF0gH2UgdMKz1eNt9j/oUjXyeEbX7fzcabWw9baI6zSv
EzBMv/IGkF9qDj25nFDBznN54Yjsp4eZ+pxRXVKEuKEbihGA0BSuTKiTSlU9BbLGLriWrZ2VEar9
L+vCkqoZhhKPXrgh/9moK7WY0n/hhF8r4ImZAt8PZdfuITeLHc5v487fcA/azrCwSjrhBQ0HjxF8
2WK51Jxnqkm3oeZ02Hth7eoAAvUtj0JzILREtRxAfP5HzzGx+1GTNS4TC1nGm01N7K+M0vslJ853
Gk3D119QxY4uQ9EOdb+j93crqTN6Tk+lkQPQsveq/6Zq08YsrKStgDeUtHFLCTXTDBvBm3Lr6Aus
yUAbhOxaigq2XI6cCRiFHJCWNCVDqYnFODWY1+en1zwRxie2YSdOoQdxs/Rb03wJ+MHZEbxyrwC1
vrGWpcKIItmzlVSq1o+5UHHCOtxVWQMjZL5IpsPQIz61SZNhivsaRTpwY1GmF0BYy2qkvRNvExhb
IAYmrZ41AMxFLrTI8iU60CCjVSnTbiHylncGq1bgJyf9MT6gFlTga1Yh4YoCfPVdvvCFeS5oWGFS
+v0kIYb/vRoLZDHGzdyj2+MPsz5QFOK/Fiac3C0i5D2/mKXNLiiUk3q73XMQaUa1dGlMAIZT0C0d
PO5vyReUSkCTKCh18vEKGztepHz3diu2vveyH4cB0oKM7/eaC9aThB1E1FTr035vHE2IxBE5hE7y
EgLDQV76MLdkjV0eCTEOSD+V34s2Yq1A4cPCsWngGr7w9Lr+KPcCu+6k9Kzyitr7exu6r4KPj0EK
taH5RcUDHRVEtCCLa6UM7WIRFnZZxBe372l88s+Uy/QhgFJJIuomIcwJtcmUVqaQpfGmpgsW62xd
WGSbC+NpWKfX+beeMH1AvY+cpPy1y8NYdyTU6Zm11KzKzOcLE4IrTwn5kEf5F4+hCcGTxctFlftG
CSRbSnqx9vA+7sqCeSPoYFdxhvi/3s3AqMT6rHho5Jmc7w3Z+W4H9BVw53CO+YFWAp+JcQiyFGn6
nbocJRMTTcqfm4TbcXA70RSSaS0yCg3juIGjaNE3zuxLhg0myVXP2kuB6Hb5FUROnu7IiQVx0iBr
WWVhYtjp72aJkYUaAJ5aV3/xqZMpHRxq+QOXkmW9zDF9fQ1vMPcIFk9dgXaFeHQd8P86dDbCTBjE
fk6B7qlOPha6gvJR5yqxJS2o7QYwyYGyUE3/g/xgo0Ek0uajRsK6mAMT47AyB5GX9FEIJxcRCXV7
lsThlBftqltprxUlRoe9G2xyFz7nJgiWL5MjGuP28Tc2TWK2B71XK6LcfxPVZEDgQAEz4It2yzu7
tqEalY2Xi4lEvYEQUnUl/MtNIHPxUjgDt0or8sCvea0unOMoxlqp13hmDToO8W22nuXQ1MEwBzpv
pGX7q7pxmm13pi9ffvmSj/7c3oLTg2zmWlCIApZAPFFsTYsX+cqszwhUkMH1nTHgvwPDq0aBd2NZ
VEuiMYdHQABo9RnbqIxNCRbnuc3azh/Ccg0Q/Uw6tlXRPf1LO/xso+kUIQN87ehi9JlrgCNumUxN
DdX840iZ3pVGXKIXxQYkR41y1Bth+WNMYaPPea0vt9CqOsgtfM4qYNoo8Dn2sr/BsCWZ+wsZ5LnZ
io3sxohKbcCagWQwjqlffFyKw0QCy0sYpMEHJ61LnfGw1+/A498dLBOo8F/8rLrAJXojW0NckxiI
vaBmT1iQCOZj98JZarTdh3cuzziy6EPuii3xQdv5kM4fN2Kqv9Hrv5H6mnw52E1Axchac3UEBhZS
xjYxzVUdk7nCCrwfIIFUqalTlqoliiPZ5j5/yV79XA/Fzn/32ZYo9/URPpK97I8SB3FGyZDFcwAl
KjoNoh12YuR8LcN1aLzDS4mstUVkO9mFz3YOlDhYSdj0NGVlIg83Sp/GJK1zr6Y++E8sA7vtqQf2
EaXaLoExXFwa5NXFE9+HK+HzHEQhu08gZ6GPubz0IxJ6WN9sJYruxwRu3Jom6hLmYivH5NZz/4Mf
jy9LFXJGBz25ABhQ6gND2x1+NMFF1spR8BHvHFgJ8Z+1KfmxrohTb4LXCAyWHfsqB/jK/klYtKQC
EvsU+P03LsL4PWCL7R0Zw9/eihapH8t7mREDJwsY88m4QqFSavNwHKHCgkXCMiv53o/o4/WyrsSN
jDiCJvy1AmTydkUGaDS9kiPX9oXE2tZUd/NctpXMiF6BO3n10aDXeBCO4cs5md+NWfSuGYi2L1EG
iQsHxwrIzHhjvQAiLq1sfHXELTAscckdysMkWK66ai2fPEEcIz1Wd24rdc8bomjvKnso+kLYKDzK
tVzZVZoheIMoLcFAEc9olHRsFFy/BHqewzd9qZv26C3jgzd99BneSzWz3twRnFxDWDaoQf+PKpec
5UpG33ipcSHOH+w87IQzdiVDc42fTG0Uda29I+6xwsD7BFbiNswATRkQwRJqePkjOJlhGh2YM7Pv
wAAJJT9xdmtZbN99P38BuOXlk5EZh5i355Vl/bVjwYgrpuT7qB7PvZkoDnEECDItZRRsim7zqMXo
ZD7+cJjukzpnFwqt1RM+dGXapd8Vl/Di5C+hSemhR5N1/81E+snsADtKli56cEt/8GyLcy9rUHRt
MZxpInLbdwQOWJuG0mBX8iCOtHokwQUMbzYWmk6TlPiVkzhKMtVz5etIia+5QzWo9iqhd/0A94Xo
nqchAeBQFrXZCbVrhUwP4tkRFBFkKi8sF3HhENWa1/1ozqCAM3p3rPBINWs5ZGh4b3hHTLN1D3uf
YmeHa4s6/rbAp8Q7wyCC3Nul5F2m/l4pO+/A1R1BShWnq/nTW+q1xaz3hML7FJKEuVScvAHix9AI
TuQGTB5MEABukgGYFncbbf04RPgE5CILtgX+pGubTh4msVejUpHkQheb6H/h7SknDAC93Fv4//gL
8JKUExgg4dp9e6nUg2nNprllz7pqUQAdpGcm47+URWFnNXsvqxvTQ2wyuRSg0PNLHI96L6Dujc6f
fWxLSBmJfSkF9gXdanLc3L7qKDwqgQwCyJUOlu0qJrRO+8cMKmTj4SFsafEstvbQbjglKdO11Jq+
0RsVcbFTDhsmYlgGc/B/5aIrZjQoU3XOzMPEEv/IHcj/wL/e1YoC8PlNg9kIk+uvoVMMshEY3QkA
iTZK50IeQRFBHpEVOdgFZFchyWTPIO5kQrZt28YCgUCtJDrXhzoEQ4R7eleu/MgJjhf6g5mV1n6e
5CLfsy4Umg/NIFED7NW7VOVQOMDIC4KbXleq5w1to9VC0z1yF/U1y95SwNSap5q4wDm7XekgAGek
WjZicGo0q52h3Jt/Vhc8uitGhdy6dBWuEi9x2Qzzcykda7uo3t+MUNk5yPMQ0lnG2WgBYPZDXX5X
mmUxq+teiI5zKLsBjTbPGwVHckE/mMzIX6PepH55owPpJinY25C63W/ZbdxZ49eGUhpxDUm3Sjxc
TFTxJvsMzRYfnT2U6I1UNaQ6cjnVWnROYrsF0kt1TsN1dSXWttXySZCneMXzpYRiycAlxJHljrni
RuC50nHzae01GTzANPkmxWUH+U+amIARmUFIAFL0VVfBQzvr9SzNij8jjFYlywmWNDvVFwkI7Dj7
TtIXkQ/ScHYFL2hAKOdbFgVfq6vE31NjHyxEfzWw/YG6Uyph8kZSxmhlggo+FOUnwsiiVW8dKcvN
FWN8p21PGyE/T2FcEVVCfSNA0wl66zus12JmWCPxZK7pwRnJOklU3KYBq54eqzMTtVse51t/BlIm
iz9X2FcIW5sG9b2FK1uGJgt94Csm91rE3Kp9e+XsWjT2kx1vsoUnVBikDJ5z/CKGwAj3cCEP5mXC
eZsXB7Jkm97TLfZIgl6cxaaZWr69tj+crBHCJ6LhL6nN6EGPkRpcSac8J+TiRS2X4ZPPh3LiHh0P
w8lIsbeA+iGP1Fw1NQAjzQZVg0qS9x/3cSvsols8EfF9Hp/PKFEopC4vczlAJ+7kB0w8T8MQzvhE
6OcdM9kMomRYSrkcVhTHxg6bjzkYpqzVk9jGBs9ga1nCkjk3EPFfLZ4HgBfndbVSo6uP/feJJHTO
uTc7+NVxBPb0M6w8PYFYqamDTpQQizUV4U+St48vD++6ghrMEESOkIisMJhDEs/JobjHiZZw3D82
7wunPdB7bRuPT6G0dp5iQaHjVNOkHTqD6jIMvk4+3SMKXtxIzB7hX6AIVMtbDaXnQRNjI89dy7Jl
ekbog3m6FSkHlysDv0RX8o2l+fXX/NgGuLJOZP2l9zNNfhONgJNfFd4vf4rzD1JvrWf4P+xzKo2x
WPxdq08d5UwlFqD01nfJVk/xrWWc8Fiwso34TGuip6lxnppWJEaB/SMPdoawPf9HO0d5bjaqKnJ7
eZmUaU0ti0GWDuDKi37FQy+VQmcV8lv0bxDuGfddJXUTGjJmOn6Q8f4I9aXcdQU12hpZHJA4HnRO
b+Kd8cPA0wd9QWeHrgy5v9jitY7kJbxOOMbHfq+ZGvMmXUbUMF8Ofzb5WugkStQ5eAtO18ejCoKs
jo9k0RA0NnChrxHw7cx1deS0FD/EsOqkFS1Ivl+2tcegJZWdIE/FwBFedpHAdLILy3G8sWiFoWJf
zB1E+UUZThwKAa4lq7HfnEFKj12U7jOAitv9xnbNAATo7DnK4Lf2FhP0Q6R9dofma42CUU/Tgd4g
wWpkyAzhAk1HvwnZCt9pVsZWUzUXHW9R1CGMG5EPVP9Wi1GVx/7/wgxBVEhiXnmrcj5d0Yutvv13
2zywUa1LyAujZanOmJ5aFAYh1xMbskp3bBT7XpguS5c0EzuHAHTHjzwAEP/gWqBauyTVjkVgpz5o
I1pJ10c6AO/93ZpW0sctwmbHvQuD34q4QpqLepuUodBIzLz+2ivNJ+6E/rWdmjIVD2fCXh7G3r8V
9Se53CAqlJxK/iffeXdFaJ8wy1FIoif0BzBp3UUXbt1wUEnf9A6o788BIKP1qcOPw/B0MwRcpPAR
EXZQXdiP59mZWRDAxc1oZStcf5Xj7/y+rUJMyCurEx+o+QJlzfLWZ6EKYA4VqXXPSEyvu6OrUoti
aj0jcVnxxuuOL61BPIGw8W4vJY74jzvryvljwCCSR/FZJ+mjZXhURTmXgEFbSxWSFLxVOAGziI9n
M1r5SHa9iwQE9XPN8Oc6AlS8GZ+rA1BN8+e6v6hIUHWkse9JJM78fdusvhEVl0/EOWHuhEtAIPCK
gOXPpD5kY2sQ/MoLI/dIFu9CUlJ9oTJa9AOooC/ve/L0ntUtkwnQBmSMqmjtiImyKFed/LYx5vv2
t4fb9m23SDoNfnvqBt5dlO+wQh5QeUJkEQ0Qs97t1HrqD2RtilwjPO99hLB6lAfm66wPs6Dl+cid
RG7fYlXjkq9NvqhiIEIshXnr9d4W8dMYGA2o5giJyN3DXP4A7giCaXwfKqW+TM/89RWGLPnhuvfZ
OwzsVbkFprud90r6eiudNCJ09tNqluofpSKKP+3rewBG3rhBiKy55t9QWguIeNFfa5of/SYFln7S
EemfTKrjeHx89cG61RbzciH7bEfCQFr3I0kqoSvpxHi01pxw7R6Pd7pfCFS3nu/9o3mHyKONSk1w
YGFu/Dy3eBZoUOfRnKItG+MPceHGUa6JNbLXC6ccgcNGBY4HXUjWC9V1mJDY9WGfOikCT51x7dBs
hFc+X/HA5aSQMRgiVL0mOopxjdowkscO2yzo563ku8WnVyzwwwQQsOQLhQ/D6ckIyK1EObkMqqfO
eOVo46eeae3YbwR1buM8+B1tEGS+kCWtV3QQWOzvOSoSxmwKI5ceHkRzbdknmerrdgpmbewnJijV
CyXmHIf+eYtn51/M/eJOkETTuuBhauH/Quwq8Ei5n96kstr5f2BlD8yh/QjwzErEyAoKeDxc9261
JYoJT9fxl8ri0iko97w2oGndugszI0IxXfUsMUZVB4zLugZXmZ3P1S77PMlZMgLvy8EMXN9n3ZbP
vrpX2Y+AnokLYsjxbioG6CMemfznbg0Grns/xVrLHwUA1TjYBrdzUoY7Blc+TQuk5Sho07Fgd1Yf
5WQZ6aWRBE4BamFhCqf8lx2oFOZggD26ChSr4TP/lWlDBS0MaQ0NxRbHQXfosg8WKDHDEMdk59GF
5EGmLVYj846ghG4geGp3B4wN2nYbsuYVKegw0nzK0AL06mUUKDODMQVZgXeNEHO5+UecGxQaNnPU
M07ssXH8JQjcMQLM2O709Kfm0Xr71/3ZirhnE9FsCy0w4mCaTEcqvhePNLNwQnbWan6qtAd06UG+
EU0LvXezQ4wSf4CyRwxVV7pDAhXXjMDrazEQa+i5JDaNENiHA0HR5p0ksBcpDut8FVR3A5mhlB4Z
GXcwcxfl/FWM72AYWBbcJVeHMMG4Wul3LN2Z/up90yvhuZBEAbrI7OJyGxlhrnGhQwTnHVaicuK6
K8f2x/DOs/M/eeS0N7adR8PtCZYq9ElO3g43Ja54nMzxVAEh9t93PdB8Yd0coOpiYxs5jsOmXKl5
+SZ01Uw+oa02xBFHQtckkO+tvxBzWd5cVRmBm1f9Is/xlOhKZhrY09qIccoO0aKo/llw2JfCexDJ
eNBMZaQGRO8oXN814dEibYz8m1eFfESQgt9sXEcJ6p+un4/akPDNtSHVtfwUidLp8lhdEhGz9281
3AZHbHdR4/4AooiGzLNukLUo3UXAJJ89qHLY/TamsYSqtKSFBFQGgAKPMpbguebizO98ugQlKhmI
EDg5UdkxVuxYkrmvF4GRuiWWOjViwAsvbN9Zpp8dMR3okPAxaBvBjvxDXDKboo6JATzNWxhdo1eB
9K6qcvkN17/Aus6p4iKDOfTbCbdoQWcWCEK9h/Ok7GXpGZDbMJ6pbXhh+JMts3JoT3zhrIn9lSid
Qx8NLJ2yVdB2dy7fWH7vrmsNRySgOPlkwXrYE8PbdqBOiYh1jy86wM3Z+xC83jsoO4/v4U8xhc+E
W6CIi+nPnIwogEoQffNRDE0xCwMb2tz60i4SE0B8PAA88AsHyZt0YkXM7YMKNuHK+2oTzl4oZ2hf
SqqN+gpsSghBqOJHEC3dUzWrwWfcrdphPLbAE+CX0aG/zBEX5gQPc77ucrQAsk3v+qjgf3XZkG1x
jS9dfguAvKc2jYjwIkM3nwof9Xbx21+yDJ3T7A27n6yiAeaLgkAVhiKQX4b/sCz6rK/CmgtxswY+
jYhZje6NSGvd7I9GmgbkuY8vzun1sBYcJ24/0zBiq3CH7xpLVh2aheyhcX2MwYbyjzafGzE451Qz
Bli7zgR0W2Ru5mkPUaeuj47yBWd3qD1MwNKaj7DnTj8gNd8KfZSKBdV9euUi6sk8lo527mZZ4AD3
2eoIn1z+WaWrNdwprUuMFDeOVPdCEi97lkWSJ+BBaTahLDh6YiwPHIr9nnBZ1iDXMjTNkAh0hekO
pYCcMywjiTWmCMWC1uhwKp+IzdMiSaITIQalo7c89Mqh78oKjoatsq4tjd5/E91iXIuxkBqIqAzs
U/RIzoP2kL/+SCiZZhOb7JUPdjViQRXLM5mTmvSUxAqV4/5Ic2/V5lhbqB3EXm74WpEC8KZjJRWm
OIeNJzVvcZsftA4f7JLchdVIhSaaHYQkY7SJk8sWcJDShC7/a/lZoPXiFF5tBz6i9b30e8IcWn+6
TcDi0QCEmIJJbRbQBoX0orrkQcchG76iXnyN/06YrN2jyeVldsbkMUiOYac4sEEQZgFWxa0UIAKA
9YBHC/DnDJ7m9p4fqbXXq1GHsAsEdgpknixaTYzpyTvVbJ+QohUPtQjuz4RcsnhAxiFkke694zY4
/wONFomZmQ7gZ2r0Fh/czTw+Q/Y616El1h5iwpAp7tQFZQ28FY/FcNSYuwsGUTB++2/6777U7U+/
cV3WaYW93vwjq6kD1fC+OAxyHlOgBZ3cEYr0fE7XMDp3AXNRoA5J0bwgGIE1ukvtZZhqfaR/43YJ
BTYuKgKwGOHV9bkl0ZV04A/Sf7mCRV55IJZOFAmDANT6++aFJe5o3lbadoM1AjpIIeVTMO3RIdUL
XbjqvujCr0rSbWKpVJ7WNOhbDgvlWie1n1jApre5YbshZVtuHFqhGMFW/dPyJ2/o9pBC2U/hAWQj
HaQPB3d4ZcEYjBdDFRmu5NXB7fhrbPHXHE34cQNRuIMcAAE7ae/N9W/GcvEtK3UjB/YxsNxXQLdv
J6HbIqsh+NSUrXns218uhAB/aYjoByYROWcKa0Lee5BXpqXTjTCgubuh8EO1ihTOOvnclQ1du4KI
VeS1Z1blp+yoKoDaJFrecCdX8CEmAxikcpJjYiIDpc3E50CTulcFJ7UdxJitqpb94PbDBaibvLtN
xsqrtoJ02f+ZqcXzFfGQ92DwfENywLXWxAg3IS1ykhCPvyptH6ofxE+C0HvCKB6owaNyjmK4ymHR
CUeCrNMu0umUuTGKWrV5A5u/ICwLav7NEF6DoPKEvF0pL4p0Qq6pmNk2FUWgRm8Tt3TWgvw877MZ
XZMgxHqqcTm9GOnRZL0hcbJBFR492VH7GbBNvBPmCIPHOf7OSAyZf8J/wGbAvPZIAi3yxjvS9nxE
I9x3B939gaDe3jkKTNQguCyH/X1utIicUr3t/ttljzkaob69ZfN0gH62bnBNnPP6xj4gEsoYmKr/
dhZqrN5yOQatD7Pl23ntaAAGmPsqx5oQoFFUL/R1/Kg8ciJAFEX7vm9U5L5RX61VeI7RI8xJvXE7
3E1qOXMDIrZO7E7LPYi6hO7ZWCTDv82F/a0+zhBRxo3dmD9vFZMqjUg3uf78lgG428nFhKqXOPlC
fMUANe+4vgHJsgrZGJpX8h92X3LotDpJgVcOuIfUpELuxNedLo5JO6zO1BP+ZzacOuz0lXAqwvqp
m/DKc8UAHDkcZHUtl1d0K+CkiBlmU+Y3uoMHZFxCq5DKTOvO42NTvnpCzxBgdw0pEfSt0PbJbJC8
QnbrJFsaQqpvQKWJumqLfWkw6IPPjgYYRRELoIDt8fFrmfRTFoZDdn2b1S68XhYm3dSXZl+/Pacr
BrHOCQzmxmXA5NYdo82pmIWqPLzAwT+/BRQdF8ecvpZmblbmC8TKI5L1fCX5f9j+jlNID/SMkEIs
Zxmb00IOI+Ym8DZ8Hx/CI/M9G6N/mQnlrWzW1cM3R86+LTaKaRs6nGGddjnwzwbQ8Q69jKz919tu
XTMWB6DRAcqmQIb2QuwnnvwU67DnzYQnufLFNgan8p4g7H+wbi8fDQw8ipAuKd55N7C72EKqfw2I
NbCuQkuh3d543MsUo8kajudc/1wEfQ+flxWDIlVuJm5IA6tUTH8Ti5BSg+ig2+2GM1xcJkWHLUCK
iBTNec+N3e4ypmAEvr5KJkA2d4PmAWLtgy4c2RDZ69Nd7q5YP+G2l/9ttrGK/BXXl0sw33DSsNa1
klvGd/6CNpOfYisXDx/b2M5Nig9HkE0zqGdXYpZmJeWFKDD5XkLbiMG+XPFBhjWIT6vWbTBJb5nT
x/j26Y6BnHEFlGZoDPzR2MsCxdi8antdpvauBXs7lcwXj0ky1FlfwlIpmME+OWEDyNYpr1PNcxJo
Rp93RnDVnMbHdOF5nRf1hZV0eCro4fVJyrHWaVaKAiU868An8R8+2VDg3baABx1xwNYoewqaA8fU
BrYBLlmT1eSUegO4IyKi/jad/1FrSN9Iu3joykMQVk/+hjzW2o01WtM1n1BazDrHzYRIgH9TIHCf
L2nXvsbLqm5vlgoPkrFxIkPR6ZfHsfM3BtW0xgB7xV51mEnBFmI4GlWgRzhNp3jqJ8lzT8qeWF/6
CfeRbxgHjBEFJxGOrzrqCuZw2iIo1JiNYh+/oCmVoo50BDrLYxRCmzsTYH7iJ8WTHo7rO5qYtaG1
ApiED5U2h8jsk62wQuLjmLWhIfUiPmRghAmKwXiA06d2KXlvilberDvHtxhDkYG5TZJHH/NYlJAR
Qfg4gKV0hL0SeHprCuh5IBW7rEgDOUr4GovtTUrDWAvNIR35ARc2Fr2PN94falAgIsiUDTk41kK7
9zcnQg+FZ/ntIZEYxKPV+ahwq3YawqdqKpwz6S9JrViLMOgkG1lXbD9346jdC3z0Is10XLu3rLuJ
KFQyxgxj++DcV7nHd80gtWOWlhofj7X7A8reOdNf/4GYsv6UpD35KbjVByz8vthJ6g7UXEMpFU2n
dR9+r0z29QisKfg7mKNUnddtc3klU4p4VPdJQOIU6+p7AXSWH0elSiqZyZr9l0BtUH/HOMbzmqQC
WRRC0Y8rXUTCbOJMHw/fyrRfVeE9AAEYn7FJAFMH/+UZa6s4US+/r0kfyu4fHoy2oor8UP99Hd6h
sp7pF62jaXdi+2tHfSKsHvH+oCxK3Nusz0krLGU8+ztMBjBPjmfmh4Spm0M2gdTd+NXDIY2ZlA8j
xalSgdMiXGqQT89y0DzR8h+QSPW8NuDlkOaWmgZZxrOrRbv2R0riV/XoeGI8/l4aeHGKH6t6p5vF
sztU7ied1IPI8EgURUodMUjr+auQz+fMTn/aJNMxlBIsqwXelhonKYk5W8a/pQwVQsA3BGRlzLVE
fPZ2l6oZ0leXhMxIrM0z3ioQLuduq4X8WArlEUzWr1TC3BdMFfWW2KFI6d8mjz6k2eMNL3pIer1b
ZyocCKefgEH7pE8jMPkXcUZOx/u2i1TgxTXKNDT+eRGBolwNG+XglmWOSMUjd8tr1/KAu3JXGxnd
dSYIfwqDQzpGt71K6UbHFyaHUWgOSsMLUw0fvLZmIM6y8GdQUwvLSC24t1xUhSrAIb2hiFbNQkPH
k0ywrzXl4AnOfgGuZL+Wn3KoFgqi1KdztqxzTTSURiK8HfGgSvhc7nZ2RSJgCOu7RyETHm4vGYaF
3oYNkWfJKv518Ri3jIeTR8wbNVbwXpgDdjtAPTGFIFklfaUNDt3e/AsD4QUZI7wzq+JvBaXt+9BC
fG2ICQRnQvxQy/bpyhBcXOtbbAH+HsNO9ZlJVd/i28liIHLM4ZhIgoVuifjqjlGGYUUpmTqf5l/M
TzVJau5gugsLt5urSOb3l68xccpnz4wmonQUXeKvOqXYTpD5JDVMz/yO3v2DCLJGmdNQzxh7NpgK
aB5zZ/reuxB4xH8iZ0TCIf2JdgQ2y+CCOQYZ6TxOqDxR7gfoZN9iAGk7oXIRFtgsfn1Dyf5b/T5G
lGCAxKdZrS1AXyx2wqfgtP3KgJo/q+pyuftLKJfkBUgUPYIHIU4Nd1vQEQakfXREp55Ga4TpukbI
QxYhrrnClpfkXDhSr8eFEw397ztmqnNeC7eJu3kl2/QPTzihSWBJC5p6T10esa8tTrr+cJFkcapU
9PHlk9tfOx5tfAKGnb+q/eh9xtsJ8H5x9AMG0kAUjZRMb0wsM1a1wzE2c+73fx2t+RsSCyq4DrPP
xXBgOzCIX3W5Jq5x/Wh8QmA1o/BLfdlpee0TivB4evPGNUqq3W/kOQkSkSjSFQ6e1y8fWO6DU76S
los/caYC2J/uObCQPKGYt/jqNEDQN0IiG103sdnB07JBACnFdWZIzNpBlNJdgSoujzK+s6o7aO9S
cHi7nvegVYkRiS/NepGXU1fXSR3i6B6qQh5nOs8Td4RkNbJKXMKgPu/Hg+ZM17wW53lpDHsG6TAN
saV8Jb1IOO5efVBJrDxbPkcK0KS3VSIL2Z2wSUd9OQHsNIOqTAcppPCMPwF45TzAKVpPxsbNvB7T
hFRxkgCBAHS1l19EL0ZLvh5wwAptGPNk4mdsQq8ul4/RbZKsmOAmjgI1jsYPbzRDV7MUXOaveolc
7Wa722zxHTK75Ya8CMAVb/lVh98B40MJM2bCsB9uhnaK69+sQqaq5FmzyCm+ihY2qlaoTVxvK2N+
uDLlHJBzBRIrIFzccDymUv1+y2QLV3yUHg+v3k127qX7tfZEXxlG3TeJ6vyyrvuTr7gSPT2cW+FN
Kizt16EyNO1tMJDT/fWmBUIsDhjQBAM3NQI/zHxFeuh6OLhlYHezwrivkB3euUX8UOXqjJ+aj5AB
uwXNJuUQY4mBgQS4wD2xdvAgtyVXN273Gh0/XxPfI/CcX8uFHDFunnANSkacD7MckUNwtYvOm3/W
MtKVkm0/kNss//mdoLtlqCcSFR+siG7yZkerNgATfMww4vCikokNXlWyuoXNECZnji1DL9N9NExW
hd7/VKIGSG8jccNEArZtf11JpfPGqp45h31yepU8G7iDtHo0LZGSye2+JU3e1PwGjzZ0+ENoKTts
SV1qDML0+JbjTJyQuq0gS/GOgFkhfnfB5dnHvNWQBXCYJ3wrbLILAZPm3LAuGtRGeSNwrFLj8h7B
gg7v3B2nZduAV0IFhmmOXys2rL0y02iucccO8arif0Z/+Edvcx8cagkFB0sST0xQFTqS1Is5clMH
YteDcRB8+ayHwjaSb9CcLlf6n3hgzSgvCC5BWfL5IjQnT4WOojpejKvaJz+0p8HEmSd4aSoaoW99
jxkoAxsLC/ao/a3iHcKUWC9Bi37a3ynQl/XrUWJ/iu/fTPRNKvlam2w/SJ2dIMwFCQuOIOri/gA5
8ko/AYX3QTIbGT5rYLCY3YK5F9VUrMNm1FI6DLKXfE54VbYLiAWFTuaesHHWVvnmx0vVFzRJh2Yl
SQiTcv2iAD3jbJ+WFehf48r5FenGLu31V8LdW4HnRCsLJqTk4+4/zaKIgWHt7c4m7Q8Z6wdE0Ap9
4W9ijwK13VoNtaRcomnHXHEn/04KClwPW3EhwT9hrYSSCHLdOO8EMPUB9MMudTqqJmpf/Ijo0HUx
M0fo1O0JT5OIQd76meck3Un05NIaUPdNI+0ZRdXwkutJnBB7WIDpcjOI8rUG4cQ6D9Qg/AtOoe/b
Nvf5u1iR4Hck7I0RcXrn7pnjYAex3qW9fQe/Z7yRp5FrDaOPB5CTf9YRCuWfl12P3/M3L3fRFhSu
9mB8ZsJwlzmkmLhTW+daoiUN8wDe8qwnJ/xRlR71GOx0a3TwiJqDxSQMN3AiSZW59Bj1eSLQlVsC
/HD6tlKLl1QDnnNq2hTbBEW5MITJLbCqdG+ZjhOMjATah9nbbbkj6CKXY52aDh8IiWJbxyVweSia
FpIZSZkCNHHBCGAqgkRKOpwpLeLDA0R3wWyCQdNHlIUAgmYbceuQhUkhA8flHW7xAxSXF8tr3fEE
hPrDw7s+rrE8wEXbS0RVRw77jpF1braMgofB8/b5z+c+PAWncQpRE6HY7qap8m7Zo6M6eRuSJplJ
8W2JtoE5zL4LqHernbWbiKuGJIia3FSseOJSqjZ6JsVLJMQ1D3Ab5bsWoflPXjzHYXxkjN8SvoNT
QiAMRDuJ46dPXrdc86P6NPEG/E/+4uhRIQU0wc3+2BpE2Y+K+jLu5H42SeNoIRyMDPRYhwj1hcrH
oNUMggE/TvCp3PhVN0Kw7lxGyG9g5TrjuP2YsNlNxL1+MZDorOFvITFPEgcUvPjd7dc8BTgZlPrZ
3pFEg0VhAzi2sAL1m09CoXs9n2iRA6LBpmh+cp5ki685T6SOLCOTRRViW/AwYfSn8qseZwMyU8Qe
fsPGtBdpwTlx5HcMoVb1eiyxGGAYgwdCakEzY6qbHY1CVSKxajus63Xjt+a9hO1v+vRf7BZMtsCc
6YiuxNDkyQu7+1QcB8JhOtv46OPZUwbbT65Zi14dGFQqDNO+Mqgyf/GDDLakvlcZqqmPKf2OaG1d
ZcREB+vKs2ONgbZBgPvVIX26NoS+cUw6X9JqPCEvcw0DcNMpbV5WpPvJZithY3gZ0bN7dRbZoOaF
/RTcLR9CDzaIWeAKReQ2oksI+alXURCoKlvYmtFftBvs3pyV33m3Y3FLy+YViuqVNeAYgptmVDLP
mkuxUb/Bc7DU317o5+uWJ/urlc+rV45q45gk8xquBmJxkyC9NLwvs+RJMwUT0e373DguR+62xPMr
Hp95IpQYIkdrXrp2t6qJlG1kJBL938gnykKsHNsy6norqa9I9KOBiD/Kejzoc0Az5qp1Mn6N5/fs
9RQdJQQ6Kj2/MofZkGrB6u74fHTtO4fm67SMYDrntJr1/8T1vOQifJYCMwqUaMXA4i8JkCwImlnR
8TQk5+kt/6jv6iEno801I5yjL1ikTvtaaImCITaWDPPiK008zG0YUSHH/bDKAviEdjpDbetPapM/
E9WWIqEBdHqXrmGPOZYZC5NvtBczF9FVEj7lN/R8YEVU5JUJIgZ/9Gp2SH59qPzaFd9SVKQiGecD
RekHJTfugymXWnPzdIBzOcYSF5zigucxEdykHZxQkESWXq/dT/rvvn8oiTTMTuPEOoJGlm+FTMS3
hmzdGsuNoBu6eAbc1gjI68eaBLfpOOSQTVrmCzJJmk9D3+mGFwCRbw74BOtG9nAvh9qIhmc6CF/U
cgX7o6dSp7aSpHH6IZHtImLdBFPE0GoTimmqM7qrE7x3+JzcNlJ49qW+xCFRnywhl7Z0U/m/r/xq
kCifhVszUUXbpfKW+GEAN70W+9/BkT/KNI0AYe7d+QJvB9PnP0n4VMouFTDy7DOhPFWDkVxlFykT
p9i7Rn6uFvbNVOjKVNYrRvhczzAp8khiPxz+EZzKn9xFDFp2hZfzpGi8XciokwDR6k+0eKcaIdj6
RadSw9NaMMaSW5Y9CHjDAbqjnx3uguGeIabHBGEi0MlVg74VFTohQh8DnUGxSw6LOIE5F4pdyCIy
xBTUuO1tdPRcTZXaf5El4nh0hJYLrHBRHCTa773ywjZyaIG4CDWZ7K4unJSbmHYswd5gwZZNWvN/
BMTtAlar6tw9RyyR6V27IXnFh2mNKQu3SnMgv1qLpyezzp0idvXBNk6cYJ5ThRCYSmell0SIJEMa
P44X5gq3nCk6Ki3OKqfd/0+87AnBRbjQ5NANaPQckftmKvZhWwi8LXyDivel9PM+vcv16a0pCzaj
AWK1PfcmaQfMOR9wdMlHyBX12obZ+cIZfXXX2T2O9P5I54nWgthJ4nZ2kjV1fqXdVqeJlfQixiu7
d70l/jfVxzO2hCoE9zzUBVphMxDjGYbc+2pCEw6+O4kkyJa3Y8Tc2zNtosV4udlXzRQhmHPN6eYL
sMQ4v51Ffu57BvwFBBuhTJ7UZPuU2JmXGp4kL4uGgjZsaN28BSNaWeWIfyvez4hEESyAMstiNLSM
61DO1A9wb/+2ERTxgxlXRiR+/PbOpx/rQLq/DhHHnvntCOzjDPUYiGg+VqAUtOJRCtbf6JcxqlCZ
ZamY/tj04QeOYHfKqTSGLh0zrhyZaeC2/uKPpni04o0CHO4+RKPwWs7i6DqkrernfTAxbyOdpBt4
E36MGPM0MxMJWWoxIzGrw2qLqtrw105buBH9S2nOr8NgWkLUPuQe6xNoIQxF9ingUSTOmWRqr3mI
t5j4ZK5osmo799EqPC3l7QpUxLlej/XkBOF32lhm6OcCJwpT9T13F/oDKbnIBu/FmKc2F0s3QjUd
UkStJwJppQgooUHOO6Ye4TTLHfmMXV9US2iH1Tu6NsKdQ4SmiIjyb2MPxEHe1IYEvC9rMzLC6pGy
hw+aJeLYMLaJ56pAJxyypSXMXGuVCodo1nI3vohV8rmd5x631BRetApbV2g/1Jiu2bCzXdv0Q8W8
YHS7/fc0CNEIS6cP41bwCJevZOsDwiNqB1WCiYMcfIphJbUfhmkytDAHASZXntfmqgsp6VlRFm2f
ZLYgIMIXCqfOAXxWB2ZJHzczjIE2ET+1w89KJ9EC0T3OgnqzasHmI1VPwcftHv8TwM0vOmI/+uxX
GbJ/4hSIAyf3ydl1biv1bNadtvaoaDWIslnr3meblSIoePBLzczhag/9xXg/W5iZiR48FEeYogo0
JQBxFUItvZdoTaJUWSv7ka6u+Y0ZFYq+V5Gb3hpuE0UEaARkKzxqjpVo/Wj6ZXobbjGKfZhVVbjh
+qQiYGGygvb5Wb/ofvsrzB3aUF6S3Hrzh5Je9SjmGbm2duvRr+JhAd+tG3mSBmCB0SAY/HteMG9A
un3mXoHDerPdfpuJ9YIBQbNPQg3MLpvVCRD4P+MuErTL6ua9G7+qtJ1MYfh8oHtSWlPkfPS22O91
callRJv0y6YlYaGpSvYf4qisMbzx01K8mOrtHrjRE2lHLidCHgZJEKwzr9o/1WJdTJmnwgPC31pi
41iAk4h8XltQwno9pnBZ2kHkLGGqJ+3mS53hKleFa+uAawjdD/VpWXdE/pRbQ2/NEXuTNoQ5P1Pl
SYuvvP/UUr9RLKoT/9zJP5vUV0nha+INvb2x4vzw6QrmwthnVHo+MXgfCZ6QiwmY4igHvhnk94TZ
JPMwNUihPAjX43nsGGy+nbTc6GRNfHmVWK4nU6S/Ku9grogQj5shPJ5PG2ScOWAMqiByn5Sa1amZ
41RYgXO8Sjw8c0gImVQf7JWkGiRVObjDnGpkxBRxLuh82KA7+LpG4t/oX6Jd8EVpY9S/olaHXDwc
XdN2tgMkmnOi0ZbvT+h3B/BLHhjnIl73ZB//9u385heSTUNRefsMtpc8z/BJElBu31JzCBQ5WEGX
FdHrM2n9W57ZRrYrrTAXyRHgf+xCPi8ubei8o3LL0TzUixKa1eQaqt1WJFuqnH7IzbDSacPOG94E
5KfFNsTYS7W226mjIzLTkevzm29qQpEe4opRZ9QxM3XxZkPPqAnPcUvvgtadtK4Bmx9qAJLcbvXj
Nj7kXRr2RXNsAzG42KAZwg+JlSL8l3pADh1j0DrPY66ApgjwYhaFVb0Y88W/NUl75vHpN8vJhb8H
x8oZlGB/zr8vWnIr4JW7o7r6/NF9I2wHOwwCZWwMcxPlOTFEaulfKgDzw0YBwaQBx8JA6ubmZWKA
nJQ7KRuEpDAApbPD2CL3T3cJQpwW7BsscOEZYEpj8Rq/18Sz9TJkJ7awCRaAPHBrnsWM0VK50GOf
JiQbYLBYvHcyR6I6Q5r7P/zkJlo9+yceAr9/e33aJfAW5TVvO28Jucf+0lsSRLSy/RQEHN1VBlTZ
cT3IvSC8YwtgGZND3wnlollqpkcEWxQFmuTsGt4e235u7t2w5h4qC34etTO8quylG2DAHUv7nVxM
assopH7RA0QYR6t1iMWYdZ7WK65ibnfKxe41niJYntrdsaiK54xl8JuKh49LV1j0oh92m8QbbpHE
QxCqBcxEdM/LxCEfyx0nPqV434ZBQTqdOjdVSTumHtWDDhbMD7avg6Qs6bVhF4tXlaUMpYgnBmtd
xfnAB/+pA8ANuU29dN5VjTFDjndda3p+iVhNq8ysOiSKgK7EVzyKs1+5CL+YeA09cxKRlJ+7sq0U
bJ6cVfWA+L7DMmZV0z7P+pznoLteAU9TXGqic5ghXI9ARjn878QqHhM9xO2/6iWxQWVijG4Q6RHz
sm2o3dNNkcWjEWhuBkdrnZmWwsZ29V3nQH1rHwnPtAeY9Z5GnH1kVCnEfbXQzfaAkRkkrcBZDagV
WF5+ybOBEZij1fXx0eLhRm4srxHt0stPzPUU8P5NQnUaWgF6/ba6ThkC2qjEsDYqPFuigMwE82Xr
41nB8cWpm51WVm6SiKgiAI//2AzsYhw2UmO6j/xsdtcnh+AuAwJeSIlZ3ugK8/mj+3WeleVt8Dgz
Dc4yQihijgWZqGG2ztTOF3BVRNjVcNLarXQIgHq+uKg+rdwvNIS4QUaPGm3EFZ8cftW/g6ZS3PGg
CVjQcnuScIHrt6JM7wncwywbFVf0OfpdutfyT8In06NaHhFrngymEoK/NzDsEvluvAE126Y99IOF
WZzgV1h6//Zaw6i2FRhxd6J+RvzBUHV/dGyeOsM/cHl7d7UdUp8dkJhGFU08WlNns3/PyO0xTxu3
cX1nJUkaF6Jdd6O9CbiVI7Ys3IbmxWgalaMsefG6WoqMgGSVNiFe7AEmlbUDCZCj2S/vKuRoTSYu
emlEceEWsZL50X7pJ5+TH6pnKCj2IIm4bDniu3nYSp9S4HAmuoWC7igRX9IdDMgodQ4M2ORqtBrL
nT/+G2qKlobVqylvVrY7fbHkP+FSZ/I2avuB7/bm8wQxPThqbWGnj5Ad4exCGRYc+aekzCeI6vUF
5hgSg8W1q7rkIG+4Bj5DyIxSY//6kSSY7RnsaX+WvYImLudGzjm1whp3AIZvgxpe1Qej6xdQ6ARD
GOFNJ9bHlxsP5DPvrynMgq8GU6HOzpmuvdvh57Vc4vLBeo2s2NpHIDWZ0helQbb6R2sa6WrWKiU3
gFbpKJaaNmckiUMe8iJcKzAvXb94F6Me8gRYtIGnBkmPjMg2aaXUEsNhR/47cPEVEivPaSNOzOzF
/Mm+CgxD9SkHNXYa+Qzt4OufVcUx/n/3LW5uvtz7PTB3GIzONjxcLcmqWQIBpkqTOsx+eVjwLc4C
r4yvmUMb03G8vydEl6VrqGjqxMR60NC3+IVuBPz2Q4MQ64U1b5YNuHVm9eXQfXbTWFeGoO4tY3sG
DxO7yOoXWSWuYkBjCmxgOe0n+n9gesX8lv61SYLoC9wjGl0ygWjTf+r18fMi0oPAwYJ4RJu8cvTT
wH26D7a422InJ3XhubcAfJSYFK2Yr3Grvd04H7HXLhk/8pjwdviIwEESZysRCIHqh3PG7poHMYNY
5ccQ6RxWbKWi6WwsqKCt9UMZbXA/befSRJ+DZSCR+R3Rp6+IQ92/uzKVopV5EldFh1mMlMwCEZqi
ENQNc5TBgK+s0U96PXIdzDtziFFicyqtgCKTTUacLwqVjrzUWD5Wj+PbXOUeDfUPvOljGp1Yd5zg
aou8S9An9cuR+aSJxuF5j2Syp2qz67nUyjsHPUhkx4FZFd+Tfh9vi9qwRzdaRVH4cw0xD/RvOs19
fwrlFQWwqOB64n/I1ovTsvXJf1KcONMEV3Fezh8E2pS/nM6y6+17KeS5O0uN/T0fSn3JRxXuq5T+
83cp4jFZ3/fmsGpMENmMJxsYjfFb+Eb13TwgnFt3GSuApTbKq9NOVR7ZjSha7FKGJ3KChhcZOjJf
YwT7VLiG16hEUPLUXOE1eCXeIzglFfSlsWK8GkcJPqgjmlIA1K1ZlQF3FFczMSumQhGyWHe8ZYsO
gyNV9Hv3vSGGfKaCqSroX/TA/n9x/sOKbWfl29dysMR6RSImPKY1O+LVrG1AwDW27Vz7NhNA0POM
hH9MLRkhvxpI9DGulhdH7Amm4IR4/bkFeHfM6Xt3OC5SzT6gR3A345JVzX/oSxIZUz8/ipZlkCXI
/og9dQdrohPSIbLuEaw7zMHIuPbTnMU34IO7Dhegp0linmjcK1niBJfeXOLYwLD/4DM5tah+bMaL
NrKjN45OakfugrvjglaTrY55lCvije5/lDOAoaC0n7uzl0VfjYPUwFZZozbTLv6YZ8ZyVyP1KShm
73VAnbzb3zXaO8E1WoKH7qA/W70xDBD3FhJtmOlUcq1o7yMc25cRtvRuKcfTWt05bTbubl4xXpIF
MYOxp/fNNdqcPtByRLPeFVU1idCac2sD2p3sXjYokpwsQl31ORu6peMzW7EKYLoUEnO7jLz6MTN5
mXVlKMblOveWSwDpw7yzomlMLilHTFxR16IOJ/YyYiAjyf+xVzvW/Do+4xtIvwgt/3HYgyEyBARn
BVYAZ6H/U0SSaTdZxPIihM3y+IGv/Y8YmP7/rP/xGpudgcJQzoaQOxWT/rDvTT1OBw55okaOH1Ok
ag3P6zuCLewPw6l4glETsxlab57APLrV683nvjJnobH/n//RE6pWOQM6x/puhfVpwK7XrPGuJP+3
2DS8U+Gitn3k9wOtRmV1UJnZr+tAptwhU45H8pesyCK/qgKMwR771olB7nT9cEGuvg7TSICyfB7D
cye8psexPHOgiLXHbyIpSgU5Pi1X0vlN+2OCIk3OPN+qmbEOvBu+BGhNGQc+LxwAasKcRWX8cF6Q
xY8GCKfGe86ZTzE2iyBSN5lqkaHFO6kcjbPPsMyEjkUWxLAPtMmiJ5E1g+CFgPeKqzy5JQu40yQu
sC3V/eUS9DdAD0k9+JJ+a5WROuj62vSrAYN7Vg3EOuGVNjelLQXDkQTWCJc5zcCdKMl9mhDKmTbg
p/O6muNU83WHOcqwwC8C+g2TuHnKz/Pl1bWUViU43/navh5GfqYDl5kFczChY/FPKuH9rjL0ewC6
9vm+mzjcr7JK+mrJnkNPMRuYA1XHK7zRS6MfMd3xef1nQ3JW08bcc3X6GcJJtVZFAgVHT1Jj8MhZ
njcX5OeG6ohfRU1tzR6lG05gN5k66dUt/pC4zrQD08Nr5aOtJ1c5CaPP7CQMddKSalkZhgm8B/qW
dS+AMyJPEZZydJKN210OCWY/suaINZk8jHl46LJqBdIs68xACD74F8xNFZQfPDgkqOPxTzhMjUBJ
9GUM4bTe3dYexiSEYIMUuxP1sbWX8mmpEdRlUL2MtN9XjoUugw18zPwd8OCtqrVaoEmxW/rrzlPh
JrMdh/kDpElWavgK9T9ch8mNTzW5OrGGm57WpMoxXeYTMr7G2DJKtNjz9G2uRmNY1AmRqmWSfMPI
vWxXwcXhYtCYrOFUOXXzD4xI9KkSUBTvDn3tMQaabUWgXmL+yJot1+PHv3+m8uYtTFTZu7aT/wHO
SqVMKUv53RAlsAm9eIQHb6EzNPFp1aWo/LfhZAmW1CXSoOL6XsjAn90ZjFyRTEgh2Fufyd8GGL4W
jK8Gd2HSxP3qqfC+zPhaw8DfmJWKSiJM6hzzUrXPXXJjJabzYxaiquUu5jCHKfY5hUv5Rwh2eHr5
dxwuTg7nLy9cNhj5am8sSQj4zwusvhfB4mHzA1Gk2jM4JL0fSjBea82KTvFXmdW83GUgNFEEQwBA
zK4Nq6O35HI+P4HfxdYghCfd/lN/4Ex7aXntWOJac10yPptUb7BxGCFJkF1oBjv0tnsDhIbaeWGx
2ITqSjODUfNLE5aHev48s7bSh4A+77DmOkEMeXtifsSn04DfrrxlzOdAYDPVP2hKlRRfuEoYFT0H
RTeg8R4ENyN7Vi/wfWqu3R7yR7V75YIQowup19EadAtzCXT8zLbqZ8NQjeMq6u7bW6mYBy5Zlb3j
IiNrQrvUTc6arFdE/wwi3WtWPla8ff0NIQzJuHj+KJHI8LLElFLNNM2Vo0MrDnM9RHHbGQRSSwmx
HnxRTZuljQ0KYCTiuwgqTRUkE+XmGBkyprHFKVKjVakcSLSiWzwK+U/UCdWrW3IUF6mrNwVOCqMs
vf8PNiWA4fPXEA5ETMyvCkOhv96quIrKh/o71LD0yc45iUP+LE4PwOMq3xbrxsMD+EaO+DN/WPdI
Fnkcb3hQCckyfzDUxG7CcoxPKcmpWo5C4DlxxwoF4AbQ3Pyms01pFenaoBGbB8CZA0RgXItameg4
lk3aVbi/VaY/WM3h80j0sHu89S/i+8DvNZU9Olty+OLr/Wyj++SJKGzeyXU+Zpghv9F1/z9aa6bI
bhpUO/Yl+YkdQzlEyExL7Y8v0333AJ1IDlU2n5qzUR2xd+fOkD01uulj9oThBhu5WoC91QENkj85
HMo33jSeZ5jj4qzyfDTQxn4cum3c+Oln44P+1Clg6tBTGu6hLjhIT7J4289Kd8IumMABs7Sbg4ok
03U/WvFRK/w2B2DPnIwMT6IFFpZZpYynrVZEnylR8NRfBqUfXFTj2Web8pxV9pbIx9OA/BiK/xlN
Eze5NWHAggfoCbY+7g912UNdE0xnPaRDB+0t80tIYFdKRJW3m1icEbQZh3sc00bBrnKBGrcvHRFH
leobtEp/mQuLuUz6bowHg55AhQF82dsYJP9DjGSG0LRwk+v16/DO7BtId9k6ClBULqOKmLuNeglu
8VwrL+xfffRaBLbXflqVMttmuOg8RbHvdgrlYPApiUX9zK/3ik6dojFiPvKW1OTQiE1QjmamJIVz
cyd8ND2Lz/v6afSvxHvdSdOSKWRtp8LbS1PvVWvD4EPGCbgv5IuGJ2OnDlF2e3gF0neD4ASPybZv
h+6Ubft3U3wf47lhkD0bvClAXUe9zXzfDS67K8cET0a9CBB0EfX8bgvGAenjqTNVlIGxx0K9ZgVB
NiPTWuVfAzGUFhDS9vbsvY484VKIXPxD5GxVpNJcNJcMMmnGnToIumB+xLqMGdjq73HIpKftFlDR
wCZwd9YgcXeQS8ieBB/yLK0g5YGdVB2+ZtwTgt2ia7Bvoeu1forp8+om6NNss1cO0bvmkPELsaMA
8ysrLBpZLQ4bI6bHfHnF61aBTO6V25UqXGDVJfcd5oKs3SI8vcKV1cFdvurUO50Kf2vy+ppiZcIw
mSZLvZusW3L13L9SZjiGtgwP0HhS35G2BI7VHUelYJQGQ/LfgwT3QMsvQgTPJWX3l1q1L3bq01Yc
60WWCPTxgiKMzE6/9zVyq7Pg8IXBXv/nwBrxVJQgrxSmgcXZGAIwLPTsvpF6xWCob5xczSvnwdH/
j1dHmrrWcYDjHODr+aS/XXjxTVXV2tjSFabiwo9VI1E3pZUqflQB83fpb2lfT3goCT3jjbs7pNrk
BXkvRjytz3t5062TthCGFXEwRz2x0/ipqQaIavwKErQZ+zDBiN8+KYVLYLsGRywIR++KPuUEKbRP
/oxFwjq6uucGrX4bsMbjOeQlXUnuwVD5RGyc++yeU+WY0GW6UC3cj0hAjLSOWXYDlQMvOQ71plqW
Chq5RFYtdUmoQ/Pq7sKVIbdghZJy+m+O901ReZpRbK77I3FFHESTw8H1oYxNpS1/wawlOmZ2KvzB
ImOKKI6/CsQ4+wcf34nkgB7R7o1J1efQdamQDKYdAXdyvqeOaIZlHBt1xOl3oHqBQfiYXDVwSz6e
au8GrxrhSIGBUmSisaRlCxxfqsjtUWFDNpdhI9JvJ8/QGZLp8JE0SqrGLTV2WxoGFUm/1CYIzVhY
lVpEfdcO3//6kWXcBs7csTH7eQOEs/pFxRgMQt578TLtXFdNlyQ1+hSydQhEHEeNQXJ/qVPiSINh
u4UqBCYRykCEnAxtfCojMv450T4P6XZEER5HmXrmeha+tZBS9Y9DQCPRsucuti4P32WWO3fuHE4P
yf5FPjmAFcEKhNXEppeHYQG3/NV8usEmBwIU+hTLrPYKnAgn4dvJ1fep/mKw0DhWTCg4htk9MDNM
GBvVshz3Hwy8XsVI6w5lYoqzGN0Nf646ENid4HwEj5drVNpsAba95xxs5bHK9ux4SHzalvcvpoPG
1PpX3Y0sY6zwukeYodXyUlvoaKbnnC5GhiTDRVcuK8y4+rfA+OUvi/82lJo3Z7M/n3le05LA3rmK
EPbGrYIe7b9HpwHC1i8Ymv5Hypch/vLOXdu5uvf82t6qBOHZrZcpnj1iJbR0pDrs1QkFeLpdeNQw
zCtF99guyA2FXMcBVc2WR8f7jm02zLshfyHRrFIUMA6CVO/FHtYyV61cFlF0Nuklg3VYZd0lefeA
yF2ikPnT2MHP21nRye/5xH+FxbifrDE2jWxXX0vQSZFMzVrD2XDg4N7dqV5nBW7yozLf+10DCaFv
nWaTGEOmtxfCKv9hiw6TisgDP9vDkIAFubgXjUQwaiednzVlDJMtYrVXUmcC53rGPOyFH1Ud5Y6t
G/bdYHsJSnx1OPlUvLI+Pdgc81Bnwrr5FmtE1DBBRN/Tn/zpAhITgMjxYT3qr60qmgYXvJ9uXzTu
wZCyu81lMOVlwCslCKq6bKLlV6qndRMhPwiDy7tMinZHS4zLxvefXrZqkSm6nnt6T8nL/XWAWYVO
KeKafW74WLpOwA3Tq/56aMDHcv+jExqOXdI8X6yrV+dI19bTpyynPuZ/SK3mwn6ZRiFDXHHNCpTT
AeY7xQAxf8kpoo86L8eKGvHmo1PYUO7busOJ/7+iJj82bsPjPGuMCeS6n1Hz1SXurliOvj3RLN3L
4I6I25m2B+4mSo/9C6f2owyeTcXygvgCSW1QwYvxw+MmAOyywOd1NyiA8svkKfc0+iz74003XuoN
KmK6/uSmqYhKsCSnuXhJrOx1KpLRQIkSlhTT1gQKXCoAndZOgwISFhOOnmn83ZRhaqIRYZVyQSEb
Zs6SSrpVJw3IR1pxs+92BnKaeG2SOeyD/hi14+uPPDtuOqtjOun0IvTkNiYt7DMdAR/MNhTSDX8S
unxt1vWd+s2IJ2c3ZeIbTKW9rliWXzOqQN8XAIfbmKev2hXydzf78zbgLZukNbmUKDIfkoP7zXNh
Cv9HEmLW8oBipyU+gHbmsbzhxo+xOjpXQ6n8G699SK6X0LPhOTEZNkbRFPe4N4Z4A7iItUriqTSp
dsiqHz3/1ER6DWnOEEfs/qcPB10AKxOQuh9ZETFb94qpxtqGpYBNZ6kQcOIpCbCPVDaTWT6DaowX
rnsx++zCWA3pZ9lMq/Dzhv+1hrQacRy4OBimpbxewS5pkI3kcWhCGWIs1DM+1iTM4w/nnOrvLFqz
OhOF8Q1gB1QEocI9nwaUBabfpcd6CtRclx1I5rVeyH7tZ2X/I1oToyRt051hjGzdjCZkiemNwlAC
cQxV81GpM5NCgYqpDkJD5yHUuvsvCQaK/xBEwXMur+SwtRuqbPzpe9VSDonC2g7N6NSldM4nGnTN
C7w8hQ87GqPm9PqEyV+SmQPtKZiOCT5OWp95+ZCsBeN++9lhy8x7ZaIsgrjROg85O5F9kVQroxT2
2DhtXAwmtdvPzO+ivT4AZfOYPCEr4xNW8TPUWtO/LDNjS0S46M/Z+XAKxh4OLdbKhBqNamVLbeFU
sNrjmKqxQBCGKG1PTHFvlvxqWNAt9SCFgdEGdgkw1K4nXZt5Pbtml8pW2LvAZ2WPiVuBuF2qC7j+
0TxyOG3J4VufuUYuf2ZgdhFDf2K0bWSgB8gDJXFUMZqkJih7QQlaS69eSKJqX7QW8iS83JxBkICh
VhOBcMZjJdWuWUd+QsALRCSPoksRnHIbBMvtyQ4f23fLCkTNJJsOkyCo0zVdtZtDNWBoayJO66Mx
d/thOHc3uWh2/CWn1A536ABRnbJculP85TCzfg8T2F5yFh5hm8hbgUgxbqnOZ3HDpbph9czIaLwa
I7plDSuSBrwrtJNn07nzDXnytfVVdvvMtRdOLz9uH34pNCni0e6CjmfulgQ/6WT96O49z5Fjb1n5
E/3FMUbjSnsfKONy5tiLj+rltDqfw7gpnUgosaPm0W7PgSSWYOHAOxrsU5WrjWe1vC/i/HMdVXCC
2hSCUuOYP39NpDvPw9+MzXO0RIQNkJHX371/lkqfMUgJUvqjhu2I2AqdCk2cMH74nZEb54UjYoyi
GcVmjHL5GI1pFnTsXGryNYZg73hvqILbmcvdB38AmjpOlmvpUBiX77KNdI4/TfOtd+R39VjMVNi+
ce2KPGQhRYsaJlQ9RzHezDnmcGOY235BQyHqjsfVcXPBNS5/UW2oTuKrHKDmpwKJjQmIDsI6cDD+
w0kmtJul9gVKxqAaViXORmGZxhVWdRY32yJdLc5yy86R+Bk1MvTAVA5sXni7K9PWBwsy76cQfO9w
+zzGimY0BERHzTESyUnaVyU0rJHGowq7Z7C0kdQnvZektqCD5PTaJsDoHIaXWznFwKn0yk9XgkgI
x0axv5dFw5N+I9VPSYKF6ewvVC+Lg5pSR/XR5EGpVq3ynX4W+EV+Grp6WcZlhCfe32S8IvqZYYA1
3Jz4kZU0oTNtjduJbR4a9TOxQ2/8VAJInchxD2bK24CLDK+7teUzGucv7VaBLhK+9QnSjuJD56KX
UYiUK3Db0ATi6wtYNH/4dtQz4Etm8uVm9N/F9oJ1srG+zoOOY9XWYSZFVlrulOi8fagKGy9TllBm
WcSLAAg+z2O6BdPgrumPm+JWq1NKwZ3octtgj3L2KEPDieTStqMNQ2p3JGDTOQ6D20sJEYKpK+6K
bu4rGnMGEuhjLtW0No3GWwlDvDJhR2rXlbfS80KuNIavDdwx+9Xu5Mv6ZOpnmn8a5PdV1sv5/r/h
OQOddjAcaO3DrWc01tSoIqROZQ6Qye3/47p/xKl3m7Borw1k4w/YY6tbQlQZLD+/6DU5lBjfFPp6
eYW7aitSx0CIswl1nw5R6ULy8via+1UGNs/uUst/p+c/tR4POixL44fM96cenfcfUevpppmJ2OFL
3RgsM7w46p1W1qP9+0lMZutNbPjYP/EYAdrOW6AnrnpJBKgiH8gkxKLb2JueWrLX3z5S2wGzpP0a
jwIUnFv5m4XjepcfzQJcJJOrfLL29fvXFdkYAgImfOoZBt0RGExvs3l0YP9oxYPm5HpHHKQhkPaM
rvmcHLCyrd7nLTyTx6MVUOBIrmQooh6crtMWzOpvsAzxSd/q8ojSvobN0nMqPtvcvPe9uIZ0uVpw
1EhSnUycBaOlGHmji05N4QYuKeaOcPD3AElSjRWIxGfVNrrNEq+9YVU+MyvE0MVhP/+1dd3THArr
aU4bTIdhs785kUXFUPvlWyBVtjTsmrDdOsGvRlBSb/vfdkfxDsWFB+zy5c5pTBiCoN1wU/1C0Sjl
hTVL2aWYM2O8+wyPccQqQtXbzLDyrkDYAL/9wbidV/r1ChrDFA2nUgpU57kFu6DlM3hzb9ox9pNN
wAK/bSxsHJJpuxKYRnyCBw2pCQeEp2nUtOiwO2FtW4JyCFjE5eMYR2Id7b8rWcPx0HCGdK88Y/tc
z2/oc1x4IMIJKLyFDzX3h0D7aabhGaljFKW97EWblAcDstsZvRRcP9adasUzph/L6W6aBkpHnla1
yHyMjmxDg/wxWauqMiDUOOwZa0upDSDwp2xaIht6ppU7kPs021TZGfb6FtAIMdlr6nCNER0LqPOW
+r31QhlNjPgG6Hs8fiquw92IhZ0HeWUAuP20eyoTpYOTc/6CIT3U4bP66Pj5tYSLRWuIRGuiG5wd
i1KxYeEYJpA7aNEpcUXgRURVpdYG0sgV+SkXRPvpVJCtEoaZuPZjq66vqBduY6arZo33mDg3Iz+j
QYePpAS79jxcNbjncSmaQg11H77PaMZUYJMr62XvCPotM4PjjNfg/6XH5b96Q23fwec7v5JjRZpD
KzEuXiSd9Csw2jwu6ELUki+CLilPCDE+ekSBJgZqymSoGJifSsg2cs54z7//mUmo6n4ELkone7dY
5HH/EWLqJjmqGaKqDazvIFaZGkcwZ/okh+dlKpbiaP45DpJ+OxZtYZK0rFAJ4GDH+6YHjHYt0ZE/
eWvnNuKw8cxhs6X6jFQ/KfVzXA/UrZKR4yOKmsh1vPVSPhFFQEHJWufiTD1WQS84rhc5y3XGvtZY
mIHFnAA1WaST77IoU3x1vOF8/aSlL/IFpck5aA+2Pksbm7CiJsX5865fv4bX6zFe08kigPleIyII
JXsYZQ6zFxgHRG1OnCja8KEN00EXddXbxbdprtdbHlKPy8FLpDJX4RRoLb1PzsYwCc31L6M8rn1V
50Zgpa6wCMYNOv3iCTXh3OzE5RGlES+2NVwh70fWZ63BmgZS+FvSgQzolZAlvq8ys9PMQgo/rnmJ
669MiOEHI2tQikD0d/VH7eQcdRJZ73ks2orIaSVGBhyVIF0vSbI2zhvOPFKEqorK9KGCLBtDNGa+
AbMdVtg2idYuKdk0iyQbJlRZ1iVZsqne/rqnGY4D6btLB6j0mxQaEf4LmLwb0g78UtMP83tgWd2T
rr8ERKwSgzmpHJYeMyRHaDU9JYhPUrzdeu+6l0MVfU/fYCof/rTi6L+7poi4kLIG76V40xXMF082
3PVs2a/YEGzR4CuE8gRWCdyHBXuWGbNEKpfTikPgTI+9UsTXxQ0MyIfdghHcbXwi5X35O6pRqA+u
Rq51jw/8qo3lezJIGX53pfz0U1cogIqpXjPK2aOae1VB0xQ/lQU7nxTwZCkFbb8urRBUd4mKRv7a
ec6XZPVq2FCr1QwWWJy2DQqaqMpBXx0FJ81zTBpDjFz5xcKqrRC8ubL5ux9fTgifJmrA0x103qRN
3Fild8cGZHiWQuIMTzptRO7T9WSJHttsPCGId81AzBmgEz8gSDOLiVYqkf5kvVP54X/dmciXSDlG
gBPIxEVgX9NgOmNlzaLtPkX4iO8FJkBn1wg3Q8iSw103Ag0/eGVgMgX3bgZrVrUesjAfrJftzCA3
06XLS8JsLrLd37h4Y5XfLpT2VisHGl7uGV4rhZ09grtNkawfTeWCgn2XaT9DmVgUWkaKAsKF32Rk
GoeXIH++Q6UGa6EyBj4Bi6NHpeQQTSLd8pPnAffYWUXunGLgubwEG5IbzmXuiqnM69Ks3iwXnnBY
xOxBZIYo0Gx238ybvbNv8G+YZC7rGnnrwXqObyG4idNXukQgRJ/s4yilI4zwcPrth4blMzRsZM59
1db3D43+TjYKSn+sAv545IL9AhzO0Evogk9Fy28ou0fOe2k1yWmFdkTu4FLPlbXP2dpQKozeNFlk
HMPzuCp5cVoddyP4mZZ1HstRgtmvE4QFCoC0zp4iKdUumWrJjIsIPz0UlKoI5uxla+7ps8ZwbD2X
0E5z0Q0WCUG+GAchXyvIoMkMrOadBlNaFgOLjY6lRSkqj8yHXTEUacFLiMtY07yS9ph4wcbnJqFz
Qg4IjV+liXHm1uLJoDiSaqDYDReTBnFovh0cUgaMbLYAsxF5kPsSqVqT7trtKRUz4lekSRmMGP0A
AJr8lQLTB5Qn/8qIKolqN7c//QtgwVBr32UlFL7IO1W1Sp7fEU5dqeRcnJhtK9JZFB2dl1MLwenU
zIjjqAYhO6LO32QMRCzd1JnvklrNo16CGg9T+EyFy/8eamEndYSIkJ3G4UJjByf2VHnlkbRJNh4A
rFvPuP041WnSLMepcAbdGSt3KTNb9BC01skUyohfbYQWJsY/iRG29LSMqIaJLjkZJoARRzCriXQz
2h7Yr33FaBbDoejnXvWwKCWhHsj8pUueHSBkOOxWOM2WFfwz0MulnVY7fjzTHo0asMeLD7kTCvkG
7ru2znSx4wucjMuqz8aSjc9VKf0x5Lw4zxUc3IVg2N9AEpIb22yWseFjHyjdWzlaZwyfOsgEPQQe
VOEE2MxMTgBVhuPYGSd+chjWwYtHMMi2AipAwadyEcprBnYroMuzutfYc9BbOk5aIQBzk5o5u2DA
zuX51PxKDluZOFfKUrMklmRnv1ITuDedlEwZIPijudun2x9+KBE7rXtSifFlFG38IefASiFJB5xe
48dWqPu7JOhP3nPeClWJz+4QjOqPyp/CEiQZGs7obw17JkEPMDoFCKjCH/XOVjqrDSFxluku9dPG
a0hrcDHwTCa/d/x6lNOxUz/d+qXjV48FrSaalS6e7kL75zbZtqE8vUV9aG4a82S7mK3yCDeMzA1k
seqVt4ZewOtfagZASvY50pJmhlkxjVPdLckfkT8bhmGvifg2eyeWtwFoho3faBqc3IXO+msVqTch
9Bn93D9ClszCzwTi08j2rCNllFg0rulKTpvi/tzZbRrCziLCF0ecb8QQQ3f1uh17+H5ndDJRhI0h
eaNNK4Q+TG++HUE4bA7fb1/U+VPnriD58yU5v1s6WXm8hsFMqBozqoCm1hJxQTIjZbysIiFmfgBI
xcNfeeveCbVXIcAgM3tH1ZgY8Dcm7EyHRvcitGi9bU/UvidfS5mqoJhsV3k0zTNbJRPTZtht14n5
315PLSgyRwJIPizkKsSrOfLy/VvXn4v599m8/TmA4jqJ5sIao6UDXy8kERs0lpRcw72QfWRLvQX1
M85H/SOv3I4YM6O6gB94K7XF/dbaj0gclgTkKWvozcvyM797ldRe/ljs6d5q7jNCKKkPs5fzx3Cn
vRtnsVlfoMhZW5Q4clV94ZPxsOf27X8yEyZr6yVPT8uxA28Soe0aIuVfAcEgcdpffEoHJJUdOPLg
3zhYv7UAjFNgci4nKL1oeEMY9QxQ3TN2d76enF06VYj05QalbjLIAvFOpL7e/CXBjqFS9Rjs6Axh
Y3Ne5odyiD8ZI5wtNeUT4Lq1UERIhZ34aS446gDwJr+37ayPqVDSrKYQuOyY2qeFL9wqXEprhOt8
K+6uXxziaW5fyKBJc2/8+UR0gq6xvRPp//1R2eEVCNvIuEWE307Z1LRnIItR1+4TIxs60ixvuTW8
/mgQ5rBnvQSQr5A/1bZ+GiEFQBrLhOgkHu9brwGxqCpYpMFhueySr6zEylaoFJsX8VRk/DGPIAYR
9Fx3Po5pHmiI/fR3FJxDnl7KeOgFcHkByq2Qe7QEqBOnQMbLdGWq3XGafH5kx7SPJsjvhpNfcDfa
l6OqKJ6fhLgYxN3sF0QCyLn3W0gzejIrpHy/On/pL981MhLwG39N1MqC1agI5VjvErGqu/MVmZCe
oHeRk37HhVndavEamyfH4hUes79u1fcfKnxGebrJ3VAZVhCU2ocC97dbqmjQ7KkJePzaUw5Yxt7K
TMxfwgBPs5/WyWfxTz+E2hb/OecnJP7Bz9LGk9t9qq8fn7jaPtADY+eWCwjZrPHnPLOtv2aB75Up
WDuEnyQEF/UD/BduTvxyeTv1J+HHoeb/xQWXxiTx+GRDDeZEIRBp5Pl3x2esvhtznYFGWPTAv59x
89nzxBQ1EAFF/Yr0eJcAC1NQhyYNhyenZjg4IxeDfE5SGaj7OHDnwrlc62I7Eu9H6gJ127Qd/bX2
7OKQPNzsUSsBe4B2eNCBzFlkrs355T0vVMS+n8byW92+Aex3V5VR9g9oX9C9RWOXp1H7q3EYfwxO
uT1A/slBRrNKdpZ49/Gt2YoRSJMRHASsCk3mmUJs/AMI9OdclHY7fK1U7ycc3SKetrkVFAKbycaj
oAQm7ImpwMIekGaIYlAnBO8EXKaSTt3bHO/eDLhd1E68cvhKV2ry3B4OWXYxWKXbnV4SIJT3WJDt
kyEXEv5WGvsqg7Orwd98oa7vows0Wkp7AbfjVhu2wb2KxKAYVNUAjSu5idYK6lNWHhGTEDXHEkz2
tgb9a4/Sw4/ai1KKEEpw+588Wgp9bkx2mL2BuF2O0+gq+G5ZcmThDs+Bb17SlCrIwF/0SXJ5Irut
UgSSAQMmPGN2DwD2HT0xoBR50SU6n+9yp/wC0H4fubq+DSqL5L6WrLwwt5qR1mUnLboiH7EwBxs4
1D5siMPeLlHECxeDP27Ns4zs+ovDjTJ9Zorq3+79x3L7SFLKwNez8VTicnkK+bSfZprqPoezhSFG
yrJrFskYuAUaNGBFDbxJQJjzK6GIEADkWH/JIenl2pvQ3YzTLSGvl+SgFMiORrjN68diTPw59WLV
NtfyRw5GdTL3Oh+Vw2XXs5IjbV0ei3mbEgiQH7GLuevSo0jcb/Jhv5WrFIqqfq8UvEeIU9v5kpnd
3NH9o1wRdg5j0nuUuKmZICVaPB/gMgkpXt68RTLVk/WsKdY4Mnh3vuEWpD9RUO5CYE6reubwr/Ab
bpTZPp7kl6wkGxpNjstE3ISvYU4M/EDhw5/rGr/tpzVT8dn4cLIPuyWCodjeznFAC0nE0R83Xc9B
VqlMyMFmIRkmwAK32k3OyG8uFIsOQshMz4lGNc9GXTrBoKU4D/22g+EplODJrmKi05wAT1ay265a
thz6KWb+gRpbWCHxyhJRv1niMde4sxGA/16rBQ9RrJJNO7pzVLknI21aZW7NipJBYDAu7uUTgKKt
v0s30z9P/wPKadatL1ZP5XK6yBoCvcX1s7vRRniQuM+I9sqXogG9dpb6rxFf1PHkcsjNhDb/s2gX
OPiIqSz0nmJlp+cW71GWOGQNIAQf5oQgnDf7+7CE4Tv3Xile+Nzl/ee+aBxXRLAZGAj6lL6H0MCx
15CobmocKJlIYjGORdDuTzQtzaZwZ1OZXSHNUgzMzw3jkKNASYjE6w5v4Pt9otdTSHTAbcQfAL2d
29CadZnamCIAlGqxXBD8Oax96cm2qz8GPz4dPxssxJT+hK3fhLRZ5UfRnqYPe2LfJ/2wXXIllgDt
D2TytER9PG5WQQoFqrwFsmqqMAhRlguhYacfSYT/5KBWkB/2dl/xoMLjg0ZxM5dazA0o9krzyHJi
B/vK8eGqzm1CMXGTOPvOulplrnZKEtXkwO6qENMdg8+gZXpdaAU/yC0uIqUq7RJndxxAwzXiqUzh
Vf+MHxiXkAP3ggovG6AasbwqIpWBcgyYV+tv/o1h4hfMzSf0c9OiWZUGYCOyd39mWvs4t2NXTkHw
CmSkwPjinJaignNp0Pfz5ke9b80MOC5lMraF5NqYjhCLxJ4+w/6e8M8BeSTx4Mh+8iJopX9FiE8l
i9S1jZX9uqJ6NfWOG3pk/pe+zfCtv/hwJeYbdPxrGDJ+QXaiVSywS1TuGuZDYbHJkwyhcu9PrLma
+dfqYKw1rUk87wOvpTG+AaRM8oAmnovhWdLJWMcfgNUNdiJEBI0KKLDGtbXBZ8Q8/u8Lze+CQx3g
wwIgohJNumx+zaYnplfRsjhTVx2H6AoTcLW2siAJJUTqAM8/SDc9SVOMk89bXULkRVbOfgKLjS6c
o5WzCdBbDxnTu9woDulpPrFR7Kq4NZ9oOM4YCXr/A6TJ/cRd07X31XCSTyQdZNZkaaZIBs98z6G0
amOvgobpVgknZ/UvOhr7OuVk3wYz3gPPNUdNasBKv1bK9Q+N5/+x9ZhypOWpf+z9RKOJJey/DXbq
JNfVssGIvMQ88NOqHGNrWGOOrRF05GAWtnBpQR7RwNvsEAhj7cw+FtELJRdu9E28Ib0xXNC1rXvj
D8E/sgafcHLnouSC/oHWQ3FuvPnz6nTSTvlKEy1xq+HkZf5sBi/Ci/Brq7QI6jziuxgMH0jtue2J
V563tbkVLYoSc+VSWNCvngUwU8L17cbm7ka26JsBhfwKq4G7qJ3buKuEm8+/oNDj5pWy2c6UE7fx
WUrD4TPrBXScuKQY2UK4CG2N7lApepiGfUz6hy3vROzPWV38xg/PKUV/2YPnWKh3HcXDfBQBDuiO
jBN3NxH6mu0+Z0yTyKQAu5nv+ibAx5S5uqwm6QzgyLOXqjFh/sLrnVTmM9RUWYzkiR4RLlfhp8C2
LQTvi7hgvwCLPQDCxWl2IEKPPO6yHarcn9i035EdyWoNU0ud/ue4vKeIgFhCJH/PpYroKjZTOry7
6Y8OYnCV8QH9tCcvxfNmTlarp7hVxvxTLlOEy3gYVVF1RulWmsjzJM2OC4EFtnvU4pP9M9adeoC+
TguI4JjyvwDn5QsyTYNlURejZ/D5h9kdNsPRF3ZYFy3Im+t9ron5RILmShGLslMsFX8OgpH5cHPS
7eeFEiC1WPi3VtkwxrG7/ezKePrwoCPOJ0uCsbeseOBkXB2rDEUqAHSlSk8QzJWZzqeG6S1nwsOE
ojU11iFYk0chVBItKJpdwGz5zgnVLj74qZzzo7peVkYJuk+AK7SpnjTX+wlGOnTx48USvweUDNmV
Ha7Z4nihO0jHvBecJjybMedzzMSKRWW/+RWrsJRKDwbtyg/BsZQ8BTERMlT7UkE1MAVe4OybtSGW
I/5xbb3xymEqAUsAwWe69bwzJNcOPfrEckk8OA8eoCAIytoMCYCbBoPjdMQfH5rxWQkacjMq8EKA
1+K71Qf1IVTvR5dJSBPohcJaqb/CnRM42+CTu02DcFxJpeSxKNtk4Kh5cxTtkzUSB0EdoB0jIT5f
ZMJn90XTqnesYZY+pjI+l0ZGHzYGhPIIsWn/UO3Tkg3gJ6Rx0+URILhxrYgkK2pYkAdm4+VbbPaL
KCMS1lYgy2ypknu9Cz8Pt06NbHUFYC02PC3ZdSYH/yoRFbqCA2bb8Y3ettvTNfQM9fNzAjPpLOxm
QxXSFzgtaYvzz72lcflbg8LXysyoAnXSYJSp7em6Zxml9g3GADEszNJqho8nh4Cq/KUq3W2TEnma
wgAk3wKIXP2e9xwUzzlgZUEkpvZQ0d5osfEZHuLBUzT2RaMZR/iHTjR7FXMLumP2bSpGRPW74nLF
wI80r3iT09Oyb91zez0Lejz4ovRLDLqj+RbsEmDzxEIiS7XJA4W9KlfRh/piR+h5TNJo7sQumziz
8STKNdlEl7//vmn8GC6r3lzg4tW9L5v2n7PCtXSbHilcw614hDBuj3DBxkI1SiwdIHutVyQjFxzZ
vno4u80oYqKarY5LtrjeU7u2uNK6KbzfZiWzSO1q9FkVQEF1nJSE/b0NbzRVbGvzcLH6NW4qfrgN
8JKYwVvpzCOeKIsonv6wfIoM2Tbj3uAjYLpZR9uzaWqa+ITtA0sbM9LRqbAUisAAgs/YKeerMiWy
ergzgPCq16E8IBguEGAmp+2+DTr0G0gCHB0QwLTsrQwGOjCpqoc/bz8kWJ4C+X3L2unpxam7jdlo
1jooWUAEu5/z9utz5O32/dpApM+Ez0gG2UTd8bGutDlAL6tfvgaIWpOFVrASgesM+uUf10Q+bhe2
MSoyb7C6wrDo7B4pkrccXzlHS09iayLeokUQSbUwkkMTQDJBIpi9pG8za2a2OLwlNY7VuITTqa6c
Ax77T/GYb7MdORhjjsXgBZa6poDqw/D5qboKkvwxd9r+KOLtVgbpkYFVui5D7zRerWnrAU8B0Zx7
7apsA7aIBfnMsThgZjkkkun0+Rw4dwq3SMoWpLsP/6c/fFbakU7pPgxC1LNluWEs6869kEURq7tR
PidvvvoWNyNbvsW5EJdZY11t4zri4XQqLQwKC2rUo517tZahmtvxJ3KVLtA8cZKKqYazlur9/JKf
dw+E2quS8tUG/7PNAPXI7Z27cQ4zcXjGQLoz3bo/xpkd9LqD/dz+tdNAEOLa8XFvAsycy3idcH+k
CZ9ggZpSQ6W6f5rgvtsQCWw2gxRFWGTalJj36wrwYS/xzY4f76X7YNQh9OA6VjKmLOJptIV144HR
VhyhhxMr40wzCCYpirudiDgqN1J5zUd/n9zVzqfacAFZwP8m58QkICOxg0ju2ayHx3NQfYY7qCb1
SbcKnQF1IHwle8fqgKRrIJ6oxnfjkPRlE2TGmsZ/+eEAhqmcvfX3qkLEU9nsZVKPdO2y7pjj/4cs
Oiw+4whBUvldTyFJt5n2FPNvm1VqkbFmY/S2ARXcLFvUNzUEjlLHbGgiLkMKwCuttYpLZ400I2DU
OmAk90NZumlSXoa3DYf7G/pH0meR9iJKSs9q7CFkggQTjl6sdaqcA8Us6u7ymDrhvgRUWoFPNhd4
2yoFUxHKnly3jnJ1FONzmc8eWC1xA5cz+2TZqX/TNm2BBY40fRXsf7l5I6hnAH+Pa7hVtJyorm39
D+KcC1kqDMJxE+r3UaS4BjQtqh7vyJLrpsRazsJJtmErqotKROAl4NlO9GiQQqAxlADJNIt11cuY
r4mCxf+h6jr5cy15Mkz7fgDbGG3egrF1lbQCLTrpis3bF+qxb0vWALcwv6EjPQ7JQpxjtT5sPIbt
++LLczXEky+YNzSL4hDu4fNGP8NX4KhvXATVxkxAjraI807IppRnKmVn1gNJcM3dqeeh28JRaHnN
yeWfvHDm6geazJOd7dptb4X/SnG1zGIh5+Ek5KrmbBcC6nqNIO88SSJQXFm83PBJckDQ240PC9t4
dwijHguIb+6SZ7WsPWXVQEGiZbVKco/3ht4sXIEa6tGnrTv9XU6LjwP/6lNz6mZnWqy/wnV2iS8l
5pGLPa8z5q12QNEVwq0Db7vYDO3DG6IEky2BQiyZt4pxz8kBS3DcX5PtflIOyr0+dN3uVFRjQ6WP
ECJHkNS80KeEEiHdIj57j5xZtrxBCXHxbFfxa5E+EgMSTCUNQk/f/Em0CkSEJYDmY0U8tqSozdHL
usrZEWzCh+3P1jAKjIzTUg6wkiQR0AcFubx9Rli4ez+NNtYOq+wLlVZH0+XA/prpGY8my0aIlnkh
KV9l6KHPdSgqMC1wYfeY22SNT3ArZxNjXq7s1wGACjxtrqiKcf2/sPFFUMxrGuSJgU4FIcoKXjfO
m2PrzFXgPQbJuGRbVupIz/YNym4xmVLjK2VE6iQOqaq62PbF264n3xF/OkYvSxnAJbGW2zzYCM/r
QsWdEHaHw4giEDnHXYG6HJ/tu9P5gQpWIC4r+5A721KxnaIPjDOVL8bnjKGdM0rY9Aabn7fwIxt/
WRxbyQ15GYusnPC+XZiELky3qC6H2nBg46fY/YA+MDOP/rUhc1KniaIw2Zy90M/377qC23MOH7Hd
1JoU8CZrW63XZ/Yoht12Rbau1jhMkKSIH2RvievWbwfIqJ/G18YFXxUkfHACRUs/QLnA3Yejoc5x
Q70wXx8fJQ09/bgTH9bVPkQNpstOx/IJ49AWA9tU17DAFzVr0gjsp5wVuhTfHCWORG+Gt7Prcrji
ofC9ahri/xMoPPpxKEXlQlQNy9IGyvqAkOl9k/G9adZDzY3Pi4jFyJ1nZXP13oV02sf7Rq6Q7HBp
xNWF+iWIO0lIXb8J3vRQDduGP4UzShvJrBPHyVXzzIlRatTizncqO6EIjRracYT25bklsHGqYyMp
oQWBepVSrjbRgIAw8fHpGDz/MY2aBfiZiv4sn7euuRj2a1pnm/S82Z72O69kgSFDG4ceddZe2Svi
O6BOW90mLwgv9jnLdRnD8PclQ4fHmzVs7nPtOimbqm6l76nP3LrQkMb3RdTXLwpRsXyeZjnXlQ0a
pln5UbCEgrche/4jnps5ndQSSbhfQEmLyuvg9xgt0QW9vFXhQEdvtnQV40xpgxdv4izeIpBe/5pD
bDsq/RvELlHSmm74ypuGxgBJcBc0iq4B64GXW5z2G6wm1xRxMkZBv06NXnr9Aks8CdRdvAz6PSFK
NjMkTRwiihx0mLnWQUx09ACXREoz860x5itudLw1CGQBtO2RSlNXOWYe4ORbK6jA2pcs2Iufc5BK
T0xeQY/o4uB9s44TXgmf+/5Z1Q2yHuG1yVGmtykjpVMFpdmn/gQJMWqRbejbyk80R7KH8cdivstR
LAyZPXggm6DTpkDOH6VSzlvDDypezqRv3RKG+AORz4x/fhK/FbpJ0EEJFJ1x+tsFkB3edmm8LGXY
LW4fuiLfuhzgBb1CwJckmzec8vZnKhszhi/Lfftbqw/n+LRiWtNDNXH77fYpXHkdKsEGEp7IK7Fc
bHFD7kB9EKYv+/iEbfCqQgDVxNN53vOV9GjfuaiplAOPmgaXrfUO+OCODqyz1J6bHhRJO8k4UbYk
sUZdRe/C0trJEbCfLzk0d2zukgHKT5cbg655wDD+PULlHKAFkac2f6HV7dJhdBs6JgLI2OeZ+bOB
MhiCszVrfqsZTYBP4Cf9HK096LLnbZqmMjVWn1Owtkv+iVM25+a9PfTVTuYmPVCBmocY7Y0tsw/S
NZ9SO3/C7abclskNDkfP6rHqdV+Y3zixsLpGRJBFJJUDVNJVmQn1DyuAaBsT9l0dhh7MnkQNqZu1
8UI5OC9VtkQ8AcrmqvrHdNkWQlQyFM9cthCOvc5SjwGFtmQLP1iq6PAWahxrxGwjb9ayby6Z1tUL
OE9lHdcLiLe5WtVI0KzeLiGMQYYAMyzXJqZPVoJ078Rf7sBgVD85lAkEyVA+ylGIEIiCDRc9X/yb
sa5ikx05s/0OM34GieT3BcTkY2jDiQPxzZiDT+/f579ARMV250zHco/X9GwR+E/fGKr+sSzg+oxB
5eKgf2awmHarnE3b3iva4yzRrcdKKV8zIj514XLxsTq+eO/Kgi2btdfjNCWzZ2JPR4U0aV9N4wfm
NeXEMZtH05UW7A8M9WqmNZ9UglbPWoSVDPYijY/8wwkYIuXhrF8T9bgpT/HMZKRlqOwTVbeIliOq
FsP4faHWTB8FE/GFMd9MqoZEhrMZrfUe8sYSxCSx7QQr3ElEcyBYKbkSi9x5Cjss3Ci+ZMhCS9Yt
e9wAVRazdgTDEI43eBz1SyDOdqqM6vmLo8XrZW+yVnZGa/LuR+qui2k8sdUQrs4/Tl2qH51BE7fZ
wF/nwiV7D1z3a/G9Rfr2AHxkj+jVX8cvGeBLe4ZYVJl9dwzek8Ib60LVdrrrONyN9Zxefey/UuzL
cy/jHyRiwwPKXy6F/CZ9cDKh2K6+0447OHohuIrKo94ekJCo6az63uQDc8V670DcmrlWOCnMSVPW
gJ8VzD2HfzJB5j03vByzAG231Vw20lhiQwDiwbvtbHNW+pMpuwAXI7KDN0EdL0wXHdkD130nWgxe
ZrXZ48Egs+1wRgUxcsH23PoygHP98SjbpuChr86aNWLExBrfB6oEtRB80+IwAozJ3iRtHypkRbSp
M56rgCrwfpuXnVNJditFs4YQgcAyK06kSWlJ2k6T97WdF93g68x6/KpkC8QNvNnvt2T+pJZJ/LCf
jJErpg2fQ606kSE6e8VNytnLiRzbfgXsDmmKOByznaHCN5Dehl3kBXA27v/Pi1tq0p4oK3I6aXwJ
7Zx67o0wAt5dEiJQI02fs7JFHBj39PcRjmFKv4tJKLxYgwPSnYTMUENrfA0rs5KF/KDp1CCFyfge
+Q6FucPKlIeduXMuIkek/JvuD25naiE7yC8nUXlo//BQBqhb3dZFD9/Kad7aG7LX0zbtk36w60ZO
1+wBWsfcpahia3ckSmTaSfrWt1pXGGPiYmFXplZh9fL4bMQlUGSBYD1diJFUdKoIf/SfK7Z1cIW8
fSQs4d5dLYPVvSU78RDlRlZ9Qs2mW3QJXQfaS3i8yzGkp6AV9UIu03rGRaQN2MUucx0QTmJyChJg
NYriiLYeSGJs3Mbo6aqxpByE69LSDzJjD4izrxJ+MFnZH4sx+pn5I8SeXMDWcAGVK1Tj3vzCUo3b
B2vljIEkDl3Sshii7Z/QYicJUYJbw+DSPFcswQ2g2LpxrLYIIq5eyM14dresfGa5oLeiUtq6AtfN
W1BG1TxTsenrv0N8F7MOPuyh6IHVChHFhCrCuI20naznj8y44XZF/O+IQwUzlLrRd1srIQrmBFQD
ymTDZt/AY0mL4dRbwGk0WqtxM4jt2UF/fGPTraWZyy5Hwg8oPWiuaLQFLJh6R+4URx0lGeNF0li7
KL/kbsZndIvYFjzAht9BEa8k1cKnNHeCRG91qcXO6a1wiSYN2fwK/Kzp6B2RxhimynRZH5WcmWo0
xHglAXGVTRoHqLfFnQ4WEJAZbpq6W4yJXqzLnkCu8BCZqFU/+w07Cs/X4BGyrJpk9GZOs9R6pM5y
DQK0fnFA4JpJEaV06OzUiwT/wdGy6q72ffj5BxmT7+XQsv+uG1KkfTzWbAtInuOFzZ/9/q5ZzRgv
jUHIwmlXDj8zi49zw6lkfX0mGiQKZC9gR+Tr0r5z+chuPHU0P2RHzk49pdfAuaXDU9fLn0cS4vi4
zVBAVnUeOWY9tLUEqTcm3RTqT3tU71Az5mOMU+G3dEh1L+C3ZUmlV/+rP/Lq9UclFrlaa1xCTLVO
y7Bc/BnyU7xljtDMGMFX7285OrvBJ8vGfH99lZTWxIHb7wexguxdj+RyrLPzG7ZUug57v6JeHpJo
lwAr1igfwJykCUAUuKTrxlJ3RDsHH7L2YGqD7wxO4j38aplh+AEggNf4V75s5jdrqSaZTEj3hyiL
ZGq2gnKkWL3Uk9En7f0kmDENgDSUOXJG+PQi8UgJpLsJ79lT3+TSwiWTEs+J4Uh1fOCBM2UtSLMU
wy9OoX6DAvwdKz34543FDrEhqi2LT4ZW3m5l3HKjDfI4lXuACQjKK5abOKtbk9RRcMP7INDjyBeH
1MU4EzTOxVh3ghesp5/iCm6G9O3jigQdFmeZyLdtnaZB4uvX98LaGA5zkzlelOhSho3EVFG9cg3W
wiS4Ah2eyZYkoxG4gript/4vvzqlb8RYAGq2QlyPcSk3DVfszjnh5dK/enmgKFPqdc3mYtNBLxIQ
SYUFzpw3kNjvaMfS4zNZkeCyZHm308b9uJ4qjc/yzw6D1xpl/ItB+nJ3oNmS8I31R10yckpIQEZf
xAymTXfIUSvtP0wP44oOTJUX9ZYJ263P3X4Pkz1/1VPGQGB/DEhyrj2bGPSvsG0ZsVGFT0PSY5a5
qoXoyvi7hSrVVTHazH+/R8dh2TBDahR8ii7f9nz0E1Ti/AH9dGkJ8MCHdB8kwSOnp9rXObeeslym
K7oNMhejT4sgmjJaLdlqvWGyHUjtyYcF6c6iCcRQMdyVvlIL2siFP/5pSlizcUifF3Cr3/UQvBWx
zzsE9J1klOvyOWySNhHZC7tSCvJWSTgER5Nfc/WAWXx5prr7mVGxOsKxie7zqWaDWW825c+pIqQ/
Ag31wCl9jCVSGVi5EbpkBV8NiY2syNwqT1LfTxhLQ19Oq5pyYeOdcvKDxiZbZM9YNeaaQpmpm+3f
4Z74grhzvyfgZwgmJxcXNSPxPznR2btptc/hTIicol+768AwZ+xZg4xhtb2pKwYTqcGkis9pzx4c
FjA0TsdyAA4ZotV7ji0D+ACddqDBxcxR/eHbzjoTbC95mdZ0wekNSgHGpoT5M4SDwud2Jt+MOd95
qX81A6nGmDBIvVseVQSzwSYDy5qvWUF53uMKmMw9UF2Ohc+EoL0/1xGxY7r45Ms8pQp2XYpizg1T
7kyqLGRAOijVLNFdaLG8k5DnhJIA51c92nEYQ9GiivdSYdMaNZYHTE/eQE5BS7ijhLnXuCo63sbi
NrCAozNfqiEQoTQDgFqg9EhQz7oHvqGhloMZhYJe1Xum1wJhLjyqbgFeKMTlSD4OJJ+lN0FhWjO9
kYj/M1B5mu5uVcgCV8A1wPXzMWJbNZpCvL1vq1kU+d2Iw30rFyKQnXwQLQdN/t7+8Y7oZVIRvFoe
isDTUNgzl+7niNWIlSw3kxE2r+ssoPZmJhYYOzgUU/4WMVBekVvmv77v5gRjEbY6nMonAaLHaDA+
Gke4u1fRxFnSXFFOkMZf0qPu19uqrEPMKpoG5wTepcTyRvoX4otY23OwN/sSkCWY2u302ZuGussD
fUzgefKQtmY1g9tgTdXK5xwCUQ/btFwTUavqOad2NerLqRyOwV3UDm9UOeviLcEiKCjGhizDkTg2
f6BEQYABZ5QIZI5Ne3FxtFYzzNc0D+Rw3bV0zEZsp+tj1HV7Gg75Lv7lfqt3YCSlxfEGShy815BD
3sOg8Qu7XEje8QJd3+XZAozeV/3fnrreVBzfOGhyrE3o+dQnjGHaCXddQhgHFxORDM5QIip1HdQh
WbcpMXeC55N61sk2r9/gYuzqxkulCqi1Ky536tmRDNtAVxZPUDKgAL7Qd6ectRbDQmrOlG6xBFR4
HfRABMIGoZrA6twuYAOLPyLhTyGL4N3Vgz2kfx9AHrtMwI16QcNcizbXjcDxd9DbT3EduZp/8QRN
be8Ra/QTBoMLVru0JmYO/fiu2tCox2/XgBWO7Lp/e688l+jtO9KiYKzJ3g0VJ8n2rE6av/fr6ePp
gY57aM/NvyOFatgnBVoDV1ULhGgU1dUW1xcUhi28gpSHduavOXmiymf6mnRr0KuA5HiyEVmhR4ax
NcUxmgucxFAHaKgdTLr8ZmJNwnpl4Ipf8ohdrx0D5NRaGrcrFDd3V7+H2jYzMmfTYsu/oa4QyHXX
EEKiGYJ+a546HAc/XPEM+FQOZWxA9qaKejv6kEfti7TwVDcbYJyEcDmBB6Fp8UZTflffjugF9pHZ
3+ey6ThdM54h1/EkpPMiwim6xUpXIVzVdqIT2FJJq+NoM/giTWSZzrNmQhNhVFaOmvi+OP3Wfafy
UeyWEPkifKCCYe9+V2XRYJKHgofToi3/YNSVE+c3cwqcZ1QUpucUhx3MFwPHi2tXBJAeKnxj18Yv
iGInYtDF2G+kDeOd/NaGKSmifN/WejYaXaU6o/DkN0HKZ6kdZH4t4OM3AMX85CEXQY5/t/3rTFqc
n5uMjkupkitHuWYZLN8A73MbxcKwdrsldlihx86/ncRkAufGVGF3AzEVug8FDyd0yt9Kc8DQ3+U2
qJJvzcCh53fnNUe3dWSPJbYQiYvImZYhpAVCSe5/ALn8ugBnEfBfBb2LYArTErzTK9rDFQJ6Hdv0
a3Os2tK60g/wPqfNwF8D/mlbCbM5CK2LYogj0L07RkoHGeFcgAHlIAst8GaXheqbhBCWgCqe3qIa
ovhoXHUHKLh0+b32hk5qyk4Dtxu51//dk0gfM9VsVsIm3+7K30s8y9FVil6xhBGldSxOsMzH1K7I
RXmmsJFlUlS0o+XOZxcz2QhO1tWIrQqeUz0Z/51LAOmZ7Oy8zFaYUdg/1qQtNqg//EXikCA8ZOqa
ub8O5gA4dEWQH/9WlDXpG79juRyUahTTPBvF4VMEMer9tdVHNE7Bd28R/Kn8+q2Eb/vtyHuC60+/
S56IaE4425xhW9hh32b5nQesGMODPnr3eN6DPJ0sFD2FXdz0fmgguNZKxoNJT/zsF2MrtO7iE4pp
mUTuMXYjdp9FMx5cTRJ9X+Rk2umw3wLT4jDH75AvhFag4nyD1zHilXi23Xg+37B/5a9nagfsOn0L
hnf5k2aNWmJc2mgNV5c8oGt5yFwGpvJCQH/+Y1Oi8Sgb9daAfKMPHDklsFMokTusZfkiDA+CO3ua
GJAUqzx5zKbfLSKtgVmi/e2Bh90KLhYl3pBg7VNAhSDm5UioxRrty6ANgojV5oBbwHMddYDfrBL8
P5EMzChrUZ6Hy0XZTU0j8UuZ6z2TxQyIgXdilQBAXN1ISsVuiyD3rRvCoqEkUq3Ka9yKSroV7M5A
K2eoMQcDCQi+6SLHDjq5BKWJAnhpAdoLz3wayUK86lSMiO7iTAYhDEzK8cvNSKQWwAemnEB01T1G
INoSXVrvPT56bDUD6xcK1S7nStYKRhx1UwIe/yhiy9Lm0tchgTKojbJnav+yNZjpEvb2ODTih107
HPq+eOqxS4zrW3IR2wUhikN+jROr5i1mhnpaIvi5hPuqEIyiFNaOcSZFX22+G+g/dn0Pu5NBsyJ+
XNG7luGQQ3ibszH/ml2HhzBcTZ6d/XSYt63lSmfS3l6Lgpirt7q2zIkFrLinRArgMFDkBdcGZfrL
oq9TA7a7tdGr2z1ZWMoTsInM1kJCrIggCtbpIltw+VsLQJqrSzGLCDXRdF9WIROsc3eOSFepZYll
KyktGG5ZTgSqdAwSUQPxYiUfgf0W4MYgnxlrpeJVdO/U7ReKVm667RGOIKVZiLbHq4voe74CaOxQ
DV0YLpDQI6uITVv0E1MUxeJpkBgHNIZS12H/dhKHrmeYUwb1IfRUwKuBDooKHQDkk8IrRxzsV0Kc
5fySXeTOQtAe9z/DjNkbP/nb4FoGpYBCctdQ6/kXvivTno/Anfo0E7sof4OgEBTiMlf1RS5xtwdV
zmJ2CryS5hk3vVX8vfaYKYP9RBf4SPrKIbxtTq66XNdmqAmzGbX5PD0EtO/XpPeyM7qcKRQK6IXe
WJNUAwUor6rotDN1mujbgJzc8nccvW70kfs6DBmovjiVGWkmvvaYYicU7fRgnC8Q3rzKPW7Y59ar
gNbfWpujtZ/EYWgipYXUWoUu/M+6mzepBQ/uMJJO3+xxLZ0JHh/oF7jyDZyC+rL9Et0GMq4yFA40
wOE7EZZBnzg1UEt2JM123f1Bfh7ABPXS7h9S7DN0H7ywyrOeh+42GL4CWfjXJg9X9xkylhb2xxmC
tqSAT8LXM/gZMTk/9HmrqNUSxV6OCzXKiXZmYnICe66kIqgSzyjGcmZSolkrZy0XlYeTT/2LiQ1a
IFabT3Y1xqOyTcqxlL47ptZU3gPC3LiXMAr/thF566wns2yPPYab2wljI3quXIReKBLLsS/dtkGa
ZFk9wJofTr3GeGWRrNxrpbuu1Z3KcHfTx6l7c3O5gBBedzhL+m0IkdAdJXLKHEnndC1fxG6sP8Z2
ltXqw8RhKuLoQbyTI3wwBtNd/ljo+mZh0nfemNFUBLYctQWGlvc8hRUWdrqpkpvB30B3uqbKRmn3
YM5L8rCZyYBwI5f1TD7WlAEcOi/2tmt516aWvehNOB6wOSYZpF1fIDG4AewU/hQ2p+5axMDAHfTE
VUl88dWiSlUb328G/dOZRCPvf9W4gr80noSKcMZ9vdzdic8Fgm0CZ41HvNSMor2Qr/8ii7bhPiqE
8XdpCP6eoJFKiQVYWMH/u3kp56CSfT5hQJGGWer3MYRzGS3V0FjNUQMj00gjogESkJ5yEVEeWZBW
zW0Tnp9y9db33oPtZ55jkkOStQ4qE8KWkWTs92GFyYITNskmTnBJVuHo+MReHRhuR5pffWNnFNnN
PgaYWfgrZRuZwAMFSik/qBeF4Kqw1nVvlyFddJM33gBK8hJJvmbsQV+5OTYr/IwC8WtmaMKBwHiv
uYYggXoJ6Jm4+VkbNDTYL1NIpq4H8K0ekC6svyTFUP60X1Gc4SyOVbkzqJ/s7FqM9j1RwJCOozEt
NbzYLGNGMx52fYz+rVROkNuMO0FuFAdaaRLiCm9ZeFY5A9gCebL0rL3GnlhLfh40d3OAhzwoMnxi
QhLfZS+H/9VnsQms7Bk4OPpipYCzK5JT7akqDHNh8NoIyll8KRQddNDhtYpqiWj2PyAT9WNXwska
Jmg3/jtXVBpiieTjWGH5zFnfVqIrWPhOia033wQDHkTBI7W93w2mPEdT17xcA7azEVJbIZtJ/lEy
SKWARP842ZjM2nLa29rXMagQA7GI6QtVkvIovvQcrvSRIiP7ybYS82wWFILiPZ61UPD0SY7cHFmC
6uZveTdzfGHTCs+GeNE68TB0OfR5rpc50rdQIbhMTv+RLXJPjP5WizPp21kt1widfr/OQi5AAsHn
tICm75x1qEXFAtO3J4xe4uX1dOhF4f3v0sLSSTXMi4ag8rvk+zgWEfzmO9dz+UF1yGJk8aYN2uIt
sKq3sQH+p5ihRwA8iECptdx64yjtWCpy/BZh4qhVMPVkwf2Cf9oeunFBkMaxr9kS2gx2ujhbJBxK
z7sFeOp/tA28O88t/a4G2zyCftsR/StqgztXga3UJJ4zH6CHOgvDStKusk/+ZYOvKPNlcn6Rdb3x
p1kDJeV8Eh/7Z0arwIUHfbXeTrRHQyNvwyTxr/THx1rMxT78HgbZxGQu3wOey7P07gAjJJsKPcNX
QwNAPYIGJiqLJ4WRDQ34PHrWheNMXCnV0c8TdB3Sq7El982Wa4lwgToFNnh1ZbeCCpqHsFuhf50y
THBnwgWlqi7GiUvMWaj3LV+BqYu4VOVsHpkEkjVn28O+ShYHnuDBoeo1gPymXzFJM9BvcLGypCYC
4dU4qTFatidzUjZFXlgqTN/9stsiDaTj9SLq7Ft5FUBQkaUxJAslJYnGJhpOWDNsGDU9Foool/2C
rMduBHRd1ygcd4hFfsa8lwUTmFzl/DkqpXbS3iTh3Rz5BBVXdbZiaQs6O8ZnlATWRpSUawKPw8nq
cxuNmqZGgnkK39vGw1PPmqTRWmUsfUHXomNkgIJ6esOYAAxd/0oCBUf6higiyg7fZmvbKLB4wslB
2exUcvMcs8v7bvWtLUUE11PqmubRLDoyrx/DeSj+0sXHC/8pcCksFX06FkJ6FmAC1Z8uIc2wc7uX
uXgt0sENBWoXqMSIGuj0ThQj6Eb9xK1sf3vc0YlQKJX7kTSXkKUGoPBu9xekLrmSfzJEn2bad6X3
4mE1in9awDx1NwuabAZIPa2/vGZXaWhcB2X8tvMRJT4g9qjMR0LGOSvUJQp0rgyFbKCGBY8Ok6SB
UKj1AIV+inVU0vnLdRMZg0l4H7nLBSYKf1xze/j1HOX9trJv/kKDfKnfJc0M/z2jPMVQ3xwbDUb9
KALa9rnilyG/o97R1RibFApjqwSdt35BHQJz6izaS2vQ8aJ3ZOjz8U8x6bnXIabXyENJENIygTBd
ixDYZakO2P0oUta32idu/vM3+Aoz8nn77PAW7ZUI8EJp/YyQyM6pyTzcg9gt42ZKfFOaIok7PCl7
K+zH2Xw4maDoEiR+l15D8CasgiJok4F9zmm8GEZ3AP55yCzuC7q+XyInpIpn4/3uq1mRsnld2ftW
J9/u99XIl1RqhQeNNqZcOsoR/K0ZcfC6NIo1NfznKGx0GI0+ex4tw/TdJqsx0ZpiS7Jwzcd8kzu1
JWddMg6zpQ21JvjdKrnaw3SYAmrHc91Zqb3bAqlT09i7XkhkK4Oz3womWZngOGwjweYQiXOlBKpC
xCauMfZdJDb7lI7XjHTzrZkJ4uPegVEWjKiHygoJQDirYSA9Rgy/cTJ5NZ88hRoVFjaS4LzP1AES
2yqCGDVggeYscWLDt5dps9ZGLVYiqB4wDSo1FOOXs2qf+G68n/oVYOSKtQiW2Lm2fRLy7VyNy32T
M/RQ+gDxMLUzjdvB2Ot1m3Ik8D3uUUmAcR9+tTQ/g0Uj8H5l412tkS4EUWuRc/tGrN6+GN0xKaqH
F1ySr9wr8BFCcidEK4PYGG7pGEOlt6QkFEBgT7a7V5IyGPstrP5U2a/1d9vOJkUMPDUfMWTyLFww
YZpTQFQYkT1uewJ39+H2XnLNPOPR9CXqTIzMSONLifq4IPX8HoUJmkUuT3+oG1OMeHlT4sokrSLs
Zr4gqj6sE2oLYE6L0KEs3gHjRD62V73uwXCo+QBXZBhoyCJacvjRgWY6uxsErqwPa3dd4piXUcIW
LfJ00GYpuskcgrzTaAuoLcltPF8i6jhkDfR7mclTx73rkr4AUyyezyY2z4eiJEIkYyYm/cWDBCb3
LqSVKDZfuA9GcawsAj3p3CbB3lyPHg+P8IAJ4FwRrwlo2+wMGlXnY6vdziB7CmI4FwfdbSayKwcN
aG0spoQFp/YZfg5VgHuqoP2wF4Kpo8b+bEJ6I5Ss4NkworSMYKBvd6h7mysRFklpplC/TfRiBJ1b
cd9Nvwz7970ZfgnXTMATkrmnSBmbSajqj/2SJRpC9GqzjbbeVTk9SAc6yC1ZlKNoB/z/A6R8vSFQ
FjIt1Foe2SrKdsVJmA/lKjjrifekGuL+EcPR5VwVl9TKk80mAm89DDSlToaesgxWrC5780pRZhX3
WUwrTVAEgvngLp/P5d/gj6pG740WZ74hBLDHd7JbEtsZSsdsmODh5ByWs0I+++50aZO+gnwPq89r
XCnm+8rs+5GAYtYoflBrri4X5a1xJfOI+09Coqx7O3yYsCABInQIAx41IHNHq4d8cJHLgFsQgfkd
PSDcxTTlp5+Ln9JYC6KLk+vpFXzvuqG/nhK1266lQW+ic6+vwFrQXn2oljbDkrfiVFhjafq7Mc2E
Wu0PYrK/cpagS50ClB/M9O/OyX+sCXyVzMyI9YRb0bS0Pf6jc7CyW1w++iLhA7gu3uYZJLl/8+Jn
PcW39L3rg9fHgsLQhAHI7DeelcieQzGaZaB//Ah4Nh1SU58cmhPAFrlGuc2xWJeaECNCCT2cxBxP
nm8BoTt2DO8x6BkQ68R7OB87VXxAwhPfu8IOhjf5aGGBxVBqo++CNjSvZPnYr5PuqSTbIVLuRNMj
hXXoJge3MmjJd0667Pbw4UN0gt/t7V4T//D2mLAIn86MvGdPGF1ziqU1xLVw7BPivv6tBoaBiuts
VDJhd4uBcebxUnmConVvIshw8AWYZvieVEoDT0VKvkpaKUU/a0z9kXjPJh3RqC2NqKibBH1uZHQV
JRUw5mlzWZhv4ixA+y4kiqT7o9uYIBh0W7UtuCk1yws33AToYk1Y84v5Md0hzOy1Rw+Ty9xzsMyw
ypafHuyzVi/MrdyB8y3NoDNhQrct0b9hAj21yp8umP+7ZJuendKlGakN9FCQacehQdnet+07TZ0y
ygmgnn7ztSSc+tulJBoPmtG8wrYsO0K1ZKGRxYAuk6XqzAM/uE6+qEsSBq5lSZQ4rHhopwLf9maU
AMliR/ghNG7t2H0VRS5wXovo1oZL9oaw1EXLpz/MEF48TpcZ+0/F2U+Pgq6TBE47qX+4xupnPxml
/+t93xY4ZQzypi/gtOzuWQIp7s54T1f/b/S/rsx5S4z0lJb48XCsKiz5G6/+PBlnbfdItrPdJVsS
hj3I5Uyo+aK4IpdpqKHmfTod/O9akolDXaE/3myJ+v4xqA25QDpe/yVvULRC714Wbjtu9DB2jfpj
64lwgFUOMFU3wjLwHlpj/BwqVn7XSJUln78NogRf6lnShq0CQ4yOWpKbBiMguQB0uScmvNiYoZC9
alDg1oz2+9T+3PbgNiBZBz0NShOompYmI/wDcndX48NyopeKP/V9OltbjyjJwASoeLyy+CSnCB/o
/ksy/bhxuaoyFCJreKL9W9BgLYYifDIAR6JrlFpNUF+XlTEPVQcWHnhX0oD7tci6IIgUR7QUfUCY
zcD6D98rK44d5fstmPBanqYDjpdnuhGaVtMZa+CEJpbW3RcImyn+4Ea6/Kc4ZS+zSrsgVg+uWmGW
+8RAZAl2hVw4O6lSti/CYNmZ12qTBI69/6Zi2e3HZWcRY4WtxmdSkUj8qRVN5OfKLa6dQRBfjyEU
RG6O3aTjIOlfWpIYuYgRhuDVk7YyY7EIi9+VoY8v9acYJ8F7ir37xjzMR5gTjd+qHdezu7S6E9uk
Jp1v5v78dVpdxOy/0r9RfuoOeT3brUY8X1QptDVLwmBydBgg3J1quJQJNcE8NjiU76gY6AqUI5kz
UxKom2ZJJ3X0BsOh3IhTe7poFiyuqJmPRiMY63Hnm8ddAhLcZ+EkpCM+okRBhYx8yx5iMmrJ96nt
+MZtuBdFYf/F7Dzm8ikOV+5EAz8SuwYiRFNWKU2D0BzHiIZ6leWksZouMwL11wa3wgvabeblgOSC
YHJqGEpR/zM2CJDw2OjiZXxAr+apV2P12MXwZLDk7Jxsp7IjW569DlzauenBW81t8hZqqabJUH98
UvxCEJ/rUdxJg0pNvFCn6MP/WuCa1LT7tQ2m+fL38IQZXbaqvFz2OYWQv/OT4yq56HtaXw9uPpQ8
pCjE3LPjhFsw93wzZ1uOxfubN/6D0EIHhkKzywHBg5O3Fl97nFHQ1RajJUsIoqleGQj8qcAS3XTz
UMnM1ZOdrMG9c4DYQgkp92EYew37V4eiTHEiDkZ55uHUydcb4CBFsLEB1Vi+5+03sEw+7KWiwSaB
xW1HQK51aREkhFEQXUsbxcgVyVN+ErHmGyWSUARaynM+YF08ge5yYZTQ9Sl6pg30+iS61gK2U3p1
sibS135Aa63J/rovUFmnP3g15QK4eurM/BBwyVVoiKJCLeDqtMudL/CMoMXW3fSdE3JoE9CK5ZQ1
4e1gSGVy9a5l4iUbeqDD6Kwrwi4Edvb7aNC5MizYAtO8NUvd6HmfcKdSfVWba6ky7+An2CMz0Wy/
cRq1A4MTpMnW1nfINCm3CB36FVCYs1n4vpxwiXw15yhSqGOCIhrfc6QBiD7rgCCmdp1F7wxg0Xux
QxCwLTHrnogjH/KTTa+Ngzd4yrZbe+XDEJS5oW6mL1+bLRIlY6sQg1DwsxyASiQBj+vfvgqBqKZO
2a7GyNDyrRC3v/JzJBUp0qIfdAeNhmFE2oRTU1Qg+l870Cau19+Q1TvcAV6+S7H/glwjbmkyw+UT
Y5PzuYNGamRrJ0mWbGJTBQUDsBaLLyPf6CVcYp2IiB/gpAt3h/8TBhfTG9KcsRRgaGoIwPuHmXya
vvkn0ctC4J0wJKmyX0c+wyfXio3Bjaya1Cta9UhuslCRcnAu2BsXYDtU5+rmJkp+OcmiVaGddIC3
pgSYVPCKQOw1YXqs7USnTF3QoUP8umkX4mk7dT0ARY29cotjP8sadVtIkNpig+pfFREdvhQIEnbu
gTBRPe5+Ev42HmrsZ4CyJD3BGPUoV0xyQjtJUiK4J8uCjbK3nt7HWS0l9hXwrevqqUvnQ5lDUJSF
e7iyAr+KZR7AMy/jCAdWVz1zzHIChTbJTYtpZCz/X/QQtHh3kK7DbDGUto6ykhCRqu2U9I1X/P3s
1kvV6ru1opGWT9MC19GkGsmGgMeWzGWsXGRNgMxQJQGITLAh4tAiKGGptInXAwW0XXWPYYZk9qOf
8rhslfVar5cHJQV4/SdqKVeLFNEKzkfr4pi4dSgrEFn316A3t2lBJzWn4lrEjmxpJrzrWrptl9CN
sB6Ovup+liLUIs4mFYYALPHwR5Ym+36IS00KdrWrpnf/h8wF9tHSv+Whp1cuITd51XONp/27cp99
z2Cn7vr6QPHueJnYXDGEe1CxcS00OJj9iDNS6g40U/TXUSGKkDqxdT+/PY/kARPxL9tdAnydx0Em
tO0sgZiP66SPy0rtYLEEDuNhXkCMDgyVngU2jWve74xN3p7iNHebkdHTXVYVyUlhEjRsmEIVMGay
EceDlD/oTbJxCBlMNalu8CyGeXpNqxSatFq0UzIlk+HyHNZpQVIuwPWT+mFXkWVG6JC6A1IXO4y1
FqUkMUIeTBQPFenSba05oDx7hdgcqS8fvJmbehF1tyTzR9gcYwAoamterdKNvmjrneDXSsdMG7GB
apdgmeKpo7KwBBoZWd3Gwgjkgjfvo9UHyNptPWfG6xnPLYq1QocnzF73KM3aVqEVS1t/RX9QCMdI
RMjd1i+87mcztQT1EN6BME7NkXOsl1lMMUGzk3Xc2di53HCTtAiD7GiNEvNhfEbwk0IpeReaaWt3
Azow8UyjLFNOksALHjBMn9NqY8vjt8fHO3QwCPbwHzfZ3x/1ogHJqT83h6xbYrddJ/9W7Kegkaxz
9iEW+lLDkSm1bWc1p1nAbFyJNgGxsb2+wBYy11fPt3pVsG0kAi/4EahPI/Am64oFCTsa9nR1cFqR
uoYWxebK5ZfphnYbFuFE837je4nZJmi4He/pneKNuriAnXoJ086cNm8TU9+3c9JA7wJe9jq/m3OY
bNpY9RNjU2YajmSQXSEuLBGbBF5HpWfjtfJi57I/HYoxyy4YgukzJt4JN4Vkf71r8kkcZlhT35Kb
byuErh0nCAcm5m6UGc/JGUvcekO+9Pqt+Zy019+DeoTrB/Nl8SgRRJI7ekYwR68jyma8/vaDywK6
I57jyvksFrvap4BY4XcxE6u/hq8Wr1CGI3J5qVPZ4ml2ulACPLMs9/39NcrccUAb41MWpjXzYnX1
t9izLvn39JzOfiNCUt+mkUKUQhfgUCOpM0KtFrTrK8tHiFOzUDaZH706l9Nd1oSZvkpgOej1d5Xc
BmZIHa3X18ltW0dyZMDDCHDe/FvG+2Aa7MioquUyPXgtyFAjxN9ZnSKcT+BO9Bw79rtF4TuHH34R
tGO2wHXY9CKhQb0bOYa9FI3nQqTCWGgp2Ivcp6dd35qlnjrcLneCwQXPG0WVJBjL59duR5rjByB2
BmJTvsNmjKdb403tBR/zgEqzVATMEVvwcjbO7a91wF/ojmHGsdi/iUVGefyUyxUeLHi5Rkuz/Pup
42f/CwFYpqe/L300PQzu1UVLmzYC3XMCPWLBtAda5NR5A7E6XMDIpUJIdraHkgfaUVDk3fe0c1Sn
cex0Ro+dIohg9QTRIVTazyQlN4Ytxd6v3vYj37oUAEXpHEBxPVgc2/rn9GQ2M0yI/kVF6N7i/Wl0
xngC38rFbnoz0bPXGORfZknfpnicXDgkO2SkLgoy1ZVtllmH6Ka47EIHIcPsrZoWMVx6DtkOeHOm
9a+RWC51YEhrLBmCI69eh+y3mjKlq57X+oNoPuYv4tlW6Q/hAB0XtByVnh23hpBppg3B6Udg9ZPZ
EUseV24dHxAyuptle1BXgFZ9V7t1qcSonoPWzywSEZzeASrYQHajJ4afc+R6pdElct7XxHeJfCS4
0KTB5MSbxId7aakpnQSt1mdknxLfqffcuLkLWKjXgXfPDqD3RqlvJ0Sgy4wtAvHPQ6d2RoP+Sko2
0K0dm9lkXk+ymnrMfFCA8sqk0oV3AWVywa42XqklOGmtgz+5xKU2gKs7Ie1yfn9mO6dBW9oxN7RA
lZtkzNXPYyOtdvtuQnP9WHwT1M6aDKYbB6rccczzXAyBX0bjZdTTrKBoc9oK3UV3V6yuh3kj3EIr
AnJkJzVGHlDs+1iiaegOL0inYDQY1Eiw1t3WufsWw9ykvBGZmM5c1S1ZDvf6G//zljSmVb09bNEM
/V5Eu3qOyXApDkA51yqk+xwXrxFRp8UZ7n+WDJJvbadXehl3iKj5umTr/WtiA3r+hYNqoc3Ykk/A
aY8mty5OtoeWAeTqojd+2azok0zVFDbIM+CryOQ6oMSnzU3VlvpLCpinEJFCf+EH75/j2TweauUP
CvSGKUtVvYmT+aKvtIrdbRVLR9Nk94vUvc2Lca2HYTAZZMJB6QEPaUtFpWq1D51Z+O8nNBmrXc4P
rJeLC/VXwMGvBFcubeqCZnJVDLOYY4XA3HV5F6rcnCjFfO/l8ycd3TBTz2Zy/JxBRnvf9FYybQT3
QenJWAwcqxeRFTIsxfSoVWaAOv4tzPVIoI7VrKUAKvCKleSJ04kdw8Nze1QFJZcfUJQHfxQzTPSd
Tm7yJH+NHgFLnviAI6erYt1Iqt7DwR4WtTfRB27rjUAcVwU7FMrWmPy9aayfBcUYQ/s71S9u2XTX
nnnm+/42wO5t1w21ZiP+IyaV0d0oREK6i5zJFdAT9aAkWoPbPAiQ/eoM1L0DGhVAK6S6Tiyxj3g6
gvupIFaQ4ksAfFIrtsH/kSNrlJzJUyFkFqx3zADp2zfxamKadLMO666WDtJNHXIuOQlGK8EQhyIB
irnVhTeM8vbSUupNHZ08Go3jODEakBhaqKQAcy0mjByMspTmfACwZtkUgwSgiyKTdHmS7QqYF442
oZpxQnpuTEnOEwDBagqR57g4Z5h55iijHXsz1MlvjNnzoGNI78mDs8pGZ6g1wgM0nNxxGtL30Uyu
ITzcTiYYzk/OsB3bY3mwQqy+RtCpxv6GiPVc+BVhluAtsvZye/bmtdjUvdY1dMdRYM12bkI4cVPC
TKMJ2PuJS9H/qlLoAw5XyCrW4LoNvkCgeDPZdIuTbbSNL+SKmOJANuNVAgvPsR+AsrctqsHmfqmQ
GNGS8/GkIcQ1D5EhtRStA+BWBAp6xTqsMi4fDucaZWev0DwQ79A2kQCNVxnR9oup60Pdk/fWRNJn
1h42vTymMOAEWnQqXOHyP0vG/0N65MshB+02TOXJ8AsLx/WQVWd4MzHvyaGrRw5O+9rXZtRKYmmh
iR2BzhZxBaof/u5Z9IZOp5Z2vC4LKnvdXvR9s1uca+492u1YsydF0yQyRniQUhaD+NzFtN6Ph0hw
t8UlvoJYOeCIgxOH4bUzw1tNZIzL/0nSpxpXaKtKrUqlmJa8ONZzZP2PnM2Cc0Gp+FxJDy0HIQAx
OIC5BtJacH10yt9akT9xqYzKQlTYsfNr7P3aoR1OPl5Ttn+6Nmcewho3G8j3edEaJ3h9uYslrmdP
1iA2a8NybCG9F5DivlDVogex9GOaxGha9WqoTBObeis8iv9p41spUTgKN5oXdTUCTxkEftbvQjhx
gfpDt+ljV9/Tzs49+qiRb6Ls509Nl3H9O8tPmrBUvHU88DDIrtkTLQKkRBHRO5A2x820iLcI3w/F
taIQ6vc4bO7g3MJ9odpq3iYjrsSmBrRFnI3AaaGGtkloqo8DN8/81EPl7o6EWoUb8gvAeP1/G9Zc
NGo8Jd9N6VvidSSecs8xIXmR6o+XUNVmSE2PYRkFOZbh3jYsho2pIVKMGk/+Jnsfm3VdUjvVKsSJ
6wHgy7POVJqZkUs7pFjoX6WztqQLSnCCv8+iOcJOuufZZXNj6Tq4u0s3jCrsGmNdTlO17Yjq2NhO
14WKymH2Gh5GwCQ4GRhNseN9Rcnw104MxgSXHXrpQcjPZkGYS1bnEXzWOk8YRIRj3TdvsMbUV2sO
q29KssjcWbZRJBRpsK13Wksldpj/c11KYVTePctC860z5YQkGTyVO9pS4n+aKxQBasvnEZAtSALM
yxXxbJzK4QE8SbzOC97LtDCI/1OnhSGJc+4BH5Vi3WsvkAo6MJAZr/cMOUZx+CGmzieuso82xg6T
j/g5o6E8yIOxi/zaduibmUr+8uYmQWS4VoDy9vAEsU6kMt5DttFB5j0qBfxpnQdDhSVHyJDP0KAu
2B+bCvIyfln0+Kpv7xCEoBFkbSM4TzU6YjJPqNhUkQ/i+Hirb3bwVbPnQt+58GwOmSLROJw8EtN5
IhuG7vcLaAzXC99r5CI0bjvEWDl8dKnEUoVVfYifXKx5Egr3sKpIKKjYWuKf5AtGeNHo9k9GHijN
tDraUsVG91zy2fVC6xBF4YCd8Ui+mbUZgRYQmWjF0ArK9u4UCB278B3m1e5wBO+lA5aFVoeL8YdT
mMYwKK27Y5zpo9xOJF3NjmZFJG+pwbPEiA/JVTepg/SgO0X40W4rdCt0YO9RHTy9lRFpDUZz2EAS
kYAHJlsBF4ZnKw7TNlYwx7eQhu2y3Hb1X83S3r0t5fNqdC6+CramivZm2GsI18yoyamnW0nGgYMW
VTCK3Pu70MLiGv3UHLa/E/nFRwHckA+FDH0sbf5wHowlk7zDZfW0pGilGnW0EVAemWCIO3ZBU/gR
/uSXQEn2EgQqD+jpATLRg/iHAlCehMGEwdJkXZOeCO9nIeh2xvEKVONSk9dmD26dEZHTXxGf1B85
o2mWRynTb6ueCqKr/7LRYp3tE86CQqW6B71KWI/Q5u6A9po64l1Zk04phLiMTO6+5udMMd0FUgS/
76g5+B/p689Ufbw/CeOYFpfjXgPb85AFGcGbtOKE/RvTDtsqsxRvJNDuvJJU4lfS+dli/E9seOL4
K5/b3ml911goyaTvRfGomWPWgza3JUu+UX7XQoT3muiDGY43HNMt3BQEXjDS8Apayuhd4rHrbYZw
wHNVyRqDVhwhdg2H12JRgF7/L/HKYjHKvhsx9Ah12MSlTflFJaF2NrZP6ULkCk0C67v/u+wUrrC2
vdrzI/ByL6FRrPtevJb8y7/ePTg3pITwcI+2GMmV3d5MnYOP7ZpRFEXTRKNYlEe5Jl2ea/ymPuLz
6MUQYZFa1rRhM3p9Yrzw55ylcpxxfKqth3Iqa+zY/ep+KQYSOqQjEZhnhbbfSvQW6FQztAG51E3C
DDoPNGe+GJMjJAjR3iMsE5hqbUFq7wqUiNXhWGn21le2CVqbiE9SXfTIbyOcDUKJllnxTP0hQ4GR
z9M0aFnWeOwGRL7IRwPhsPWVb8oFkrKiuddjd1kNUcGuBLunnAmKUVlemeqEIFiVG0FCtvCMPxy+
BLKm8Dh3fgIGXCV+hNVKNj5n/WynMMGYPRo43xjXht9yIim8nefaFWe1KkkseonEEUik9c9a0CdR
7TJ92QmKAw2KR3rcpSu+E+0TUnsnhAN8CitVdXbnxQi1mfq8kLkemXpiJHgjS8sh+I83seYLD9lA
hOObR6KkQls3inUDoRPGRf+SBfqMMTFlrQo3ho4jd8L6Kx2LwhtibBASOUZkxrmjlr+cWkRVvj3M
AMvbQFMNXVRfaxMNMWLEzi4r08dT9FaypCRgnjFZSGQLOk7f4jvWvhlvrQczriLDNWHOy2kVgVaF
J9kIT8MjHGhdfKAf/b8GZR9k3HHb1XFIxbZqBJgfKHHHhKYpXqFdU4U4MHqTEroinKQsoQ81pAJn
ucjCxm4jweuDAabQ4ELCSRx81ijGxxz9xDqBRw+89dK0xo5jPlsvaBz6vds/R0AlgfjigAN3+Cqu
R9wxxRMWqKQEVWliMoeSE/4O25muZVrhFD10ZvkCJ5BAzmH8+kmYD3qmJn0bphv8H7g9n7qe46j8
WZ0dUr0Y1BkD/6iedHDJYlnzCjje7ooPCydfb5cnoAKjXQsAzzZ+2sGOUJXHlTriDYEjTeR5md+P
OMyO+2ATgt3MwdRIx564Z5JI0fMjbm31y3p35+aEf+x2crK+3iRgF20k09/pwWjh7Teaf4zpmb3z
xQlvYzIVVPO8xMvgGcP/Qq5o3pWRHKShImtTUkOGl+Ccre6YZ44JEFYvwZBLhaScfCf+JVZ5IGW5
LY6YryQYZqQ4sFfhrsIPoPkN6Atv5g0gu4ArMzYLNKNRCbb+5SGqcpCEb+2/83F+dz8soTo0tfwx
mPBDs2akPI65ecNZpfJ0RLc+wGQFerSe3qx4ghi8YNWoHNLig3nxKWik57ILKyvqSALYhVjc4MzW
y4YMRHjDsSSidYowE4m0NiUBOPKN57O4TiMuEq48xTdZF7VkUx1pow97RYdEXCTrLruXzJAQuq6P
qZPb0lEDTYgFDJ2hReaUL+LqoIjal9JL3auxZ+xElCbiV2AnIFBZc5cXGAQ6sD90nkqP8zvrl6QL
628mN9EL3QFwK4qK/rvyaRkjBilcv7wY2WfgA4lJtOsFfR8x05ov7ciu9B0bdvUGIW58wF+viCGt
j0fQsBczhYseHAylIjcp+jU2VZr1wgphYgMZ5hix+DR0YR29GfqBXJmzALOIdNF4LJAfA3cg95BS
ppQtFdsdkTPfFnXdu7TBB6/nAxkRyZ/WQ3OHanX+NFiVrC5vMHf6iwH597dHlgLdxlabKaQPcVl/
K2kPGBDLksnJjpv0pG3tt6NGY66E8qzyvgTaZw+0pkDP8i5PBpQcAGXJqR/ztm7GuKtYD1OyxA==
`pragma protect end_protected
