// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:26 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Q4wIRndQN1eSmaZ6vOXYI7uuQKaH2/CTec5gDLAt30GZ8dbbEz9ezltJnBsX96OM
wsE9zXA+fHm6EvLLG2fTNFVJrcSZzdJusECDQlQOXEAfhY6W3EyZVXqKBP+MSf2J
cfWBIYNjOeXA1TlJ+HZ5Yq6U1wPAsJjAaK3ynnI8g1w=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 8432)
TJCoGm60SVotxkgwNvby9g8l6JJl3tSrgvgEPX0vFMw1IpZ6FERqgaxPuDZs+1Bo
ljhGxqd7Ix+yPzwv6hDjsxe+gTcraZrzIu/ihiHqG4YefxIeGTIxXyGbQMazXGeu
QKJtsQoOhPVT4QrVk+gFOC4uuv7or2X7wR3I9CRszgBJYi6DwF//rEAfRBPCckUT
Wme47pfh+UlTsnGMgi82Jj3uLS0n/nJW5rRofeEuG/xxyz4xW1dE6f4E1yQMNdvG
GfmiSS4cqHHwFifYI3/v7x1p6b5S20mYZU8ZC7NcDhlR+Tb6wczxUHL1pbC0gn65
lPFxcgwBgQx7WMuxHx0kwoQrNMv/VenBS/f9KP41jJuEl4bt6QuEWVHabnIPInjJ
LFDEBiXV60KRDibrHTLsdaZxPBr5IdJRVC24TyMKT53CBHQwff2mfhneOkR019ZM
KHbOouwNll/McD8/sKGZWuSu2gjG97guVDNhBqmpG4WfiKebzrRtEbwpZMh5kz5l
gtvxbRiF3Albd0IVzQPgWFxIfB+JDRA1SaTPj2rddnKc/SmcZmymGj81lMpZjPWw
uuxWpV58rTbfOXGnBaqnVq4HpO62mKH+fpP+tvO2/EEPAxlWuAxozEh0cQ+0lY5c
aOfrfoAbp47gTXubcSXz0vax9FSLt6wLk/8dzQDYGT5cxt3BUCUIWqXJ4fTOFNDN
EP6+sRFR+yZyspWD0U2KWhUCrtLSmUlqH0842VgLPQI0AMhmZaZVtw8VGg/JHFBP
/PbVJLBG2VIhsHVKcx0R6DFbusWTYRmNYO63U/4jwPRHVYGPUhtyErlyo23MvnFT
xmyb7pKCmsk6aSPzLj8REpvQvozToTJMeyLUnyq/8dWyhjGPM2/SG4cxkILH5xt8
CjxKJNN14m6m32bGwTJ+cJ3KV0xSmqvGAKsa5tgDdMax/+7gXL4gXyF1CyDwXLp3
bePLXGX6C9Q2+NmiEp0nPv52h6pM5vtG3NOBsbEK0C/bcE2Npklds/FdkNDFmstQ
dpWkGrvoGjScyUYaMJeUObdau3D4vHz8uUMXO1vnyDReZkIFcp3WQU+C2Mvq/f8e
jXMB0dcHlsjip2wr4aW7sZdeEOl6Yt4zOq0nlKvlmBaPmnZR/9h813u9q7yPQW+S
ONnAosPGjB8hSgfqHkKLl4/zzlqpVmPnbus0WKnpWS9/tToydnC9AoLD/oQP/muB
ngPVNGABcLkF/UOjvUKeuoXJvDnHYJt7YJMIfcmOAtruVxUh3fjGpy+AXj7GUVe8
GqwY+H8dhPzBXlHqAQ+Boo30zJyWsySVAFLJhxTHkaonZIOo4jMsz8P69mW2hybv
/Zp4HYEYm5xg0Qb2MT0WxxjMPkc5JgbXCz6IbsLgpPJuNyZwQqtcFPgJOSpFj//b
i+Pv4kAECbIL55oWTzUp0cP/+qspBlFAGt5I/owWJuLC8JU8cY/Dadwbi/Xer++P
8mLA0YeqV9KclggoBkrpmKnNvAN3roE5yIAcNQbRKGXg1gwwHsjqVvddiu6q1DV7
aDP79tlgHEiYacOqzBo0dPbPxPIY7KWO3FrCgJ8JmUHgM+6POzhFvENnBPmFElsl
gR6jr33sv3Bni264zhVWw1hz9ZLZ1f2zhxsK72ncGrJlYiVm4cm1bxPhHgB2Ffh7
1y+ibr1k2/s+9ULLqZKYUCR39L4hipNoNh3yM9qGuEZiGsByyVGGPzN2L/wacxVu
WNydxqM1GblHRAXC4JrsPXhoOyswjBqVRIOmo+ZWQ3qw2oxPfjag0w8yn54xSisG
xNFer1W2n1YEmmcoAup4JI60tXpjzSvskav4gT7EitmiaqpiuqEe+Qs8QyCvG6fX
dzP7//O4yAM+wozZxWIuqUMBhKU/UQhMNDTRHBPrTJkDrnkxX/DdXY26n5RN2uxq
o4pZMUSyXJUHhW7/koCJ0onhHDpDLxvPy/izsf4ISQIgi9UFWfVhYCRi89flhSn+
UDqfdNW+pybHgBUJmDrN8lL3EG3433w+i+UHVUhk/r0+WAxg3f9wj0gz3gHy0D+L
JjAQASef9xV2/uZO83Hhs0zDIsXVxvEWgZdEeq4Td5UvIVzW+QQDoXHPxpgNW/Ud
P+ilN6cLpkgNfaOrhz1Kb7qMZKZd4D6QusFjbfLunqJXEQo9LBfkNviLiQTuSder
fha9BdcwRPNuKSYT5n9mwqk9vKj8Xnoq8zA+AFYW78mXzZ/9UHv7PfQotcIDTuOw
VSCEAeFj4At1n6ozmPpoyI3jJv2GQYv6erU3iO+Aln5dyTV3uvJ3EfwgEZWQYrue
ASIGtJfOYRnvj7Mu8nzxFTfUjP36iJ3ZqcE6FZe52AXjOZGkR17tAODV9pvng8ay
8eIQQ7GOxHvUqiv97ralXFfnn4wBd7t8c8cIs+iLxfXnC6aC+BRaFP7DlZ8gP0zu
fHuWwCPf2293syE1lKO2NOCXwB4nVOQGLcKjHerHXcwsW0jBOVDWfMQL9hQ19tSu
ZE63hS5WzLqM6fP1YrqG3VkSiSPkBeTu/Dlzk/0iIFfCqjieZds/xhLD2/0TVdpO
rYYZBPTG7z/eLd1teUtlyaUjAnSYLscq+AHlNZZkqoJ5TtEL+557/VRljfkVoEhQ
bhHq7M8OClEk/a/f/GjVt8unvBGxTG6cpE9F27PGaKv2d69ErU8yMbBpYBwdh5qE
fJYpDm9JqfRtVTwdwlGUTrcqD1/KDLGCm7FsfuVIhKT37sD4WcAnEht1jqmh0IFV
83xIeOXdZamN+8Zj7UxkS3aqXijDiyFyk98sK5LEB78JmKPxIbaRKDDQ5smQFl18
7F8T8xLv/1tfH4NoxntyrhU+wVB+Sp6wL5qF4gS7xQbbjMg2k51x8KaRpXWRdu9q
ltpHgW3YolA3x+cPp4d5l7YyVfsoGcqhf5QzJyI/GI1gtBMhqe3O7BVjo4v4hq41
0ulfu9Ird5Crr7WUEPfieLW+10I9Wsefma9ntRsXjuxnp+IzlifRNl30eBnL2TPb
/1eL9dCZA8ZX4civlZoGBSgl+oD9dyTKVbRA+nZFCTEx3PGfpcN/68yu1CU5tjUQ
5NuIRTv0k/wOaemX7JT62cKJNqsJ8kvJEUkpXwAvGbLTvwgcmLH2DTmX1PNgKZmb
4k5AypMDeSRPQ0uSaBv0zu81rkObWdeYsg7fP4UbWGKFlrwO2l2XDQljU4rKn7Ls
v0QDLDzLVJ7HCubGuqzw4tef+Jh93uHz+/TQtStgms5L+C8+/3lKhwyD9UX0smkF
4BSh+Ql4Fgr+baW3tZuITsPZ3osR8C1A0Gnrey+YhqmOzeqG223sDba76Ndag+Tb
cG0JG/yJTv7SDD1VtWtv41NlSdAiT1EDaTZdkdm5xdsk3pYN3DmyDSsDjOJPgkQF
qLKxN0rCObynCMGnQuNdKsU+aE23lemU/h+cEpxQCD3LnMa71DnyBCe5LmXHFFX4
5q7NqWYrupYwep18WJFOz0Y51nvXz1kMkJnhcOIAnHPHS1KP0TKAV/AzoI7WY22g
WB6bgMftjdirpFvJcLugfVOiYjfVTzyAQGkQJiUEylO07qZ5Yw8n4UNqFg1aRmt5
SV0XvrhtNG5De6CndguX+P8eLlv/5ycEOUfRFIDpE7Pj2fK1qhJAB0vSbYral0t6
fDEvkpKdZuuj1fTOW/ZxDH86eFBtlRVJnV0k4DtWRh2Pg3We5ZEUnqWRw2fr2S+u
JBq1WVN3XzRfnRxrG2JBfMp+4HOhxL8MkAOyV68/jkBWzIWYYpP8HsS+k71ybUrA
yng+ErKEOohZfVX1J6qaCeFuI1I3pyYJN4BUnVpQ+4dLK7Zwp1Cue7C8CuUpI74P
ul6IC0qcG8xxTez73c8OamlxmcSA+xcyR36S6QVlH1FfDKBHQuj2394d6MGRoEMf
KE/nsfvCeJkvjBfsCMugLVAxx/kuDQdkIAShPr/yr0JpdTr+Fc76WP3lIGcKo3/Y
SC1iB7MhcLzxZ71RWtu4DhR8fcoqmmWZtN9bQr00aKf6MmL+N/g7i4b2Ys2rwg7S
WoHmjCyIyWaIA63Zy3uMpGxw6zRl2EsfOgayjozbSfYYQZrgd/gjTNHa5unXNCOE
wzG+rqUCBsbuCONp8JS6fmZohNTHLo0HbQvlJfIROyr1LYqepTg1L84Wz7oH58Vf
NQsXkLr74aTfc3XDVQQmqLx4DK8uCQC0hwPz47pQdgMwbbzG4NAWotQs/hC94BeR
pp+VCspDN7wJrVIB+WXxXmoDFjVqvplgwYs+CVkqK3IvQm2nVpvE5tWN14KZgxMy
rkqT2otzlHoFuoUOA6f3rl28FpKUsl2hJayTRMPPa2MZ+YPXPGf+oiHxknJX6+rz
STaJfK7rTsLFGH9wWyYuf+YWlbjubnRcai7qMi1ydW/KvlLQ0ixDSuH3CZSlkL7A
vJm90x+YKajXregwJqpoNsrDEOR3KHCfKkrqlnLNVasNlWFieNhACCXpegPRdcFj
R1SyIRFdnFiDr8vG0aPF0hmqJXZ/Q/vfJ/Ky5mioZEpxgdRKRJafBYJT5dm8j43D
iO95NN5PlwL4qNkwxoBMeMKC+54GXU5nlj13iSFg16wsSxhRURomYm29zWtY2ZBG
AsrHKhPBOkmvCeWffSeV6yRePpea0VKzd7fDQcux1J7ZSG9/TAvwx3ejnQIgOyHX
etLTgEm8QZzbtmnkWN7ip7NUn2f5UkS2eh6xHgnhufhgYfhax6Jr74IMtISJ8lX9
N2a80dc2Ec8OBs3Ln4bmtradG1n28SGzS9oRSFFVWnlb6TQ//I5y+ObUhxUNKYU/
MPijv6gGvHoHGBlRPrZ7/H8wRGU5z2MEzwz8mdAGi/M9KUAP0Vzt8+8TTaZIaxQw
+Soj6Ul0pDpAskkNmTLibvN9U2jvMydi0sBkjtSY34+yM6MJC0ZgBuhlOebXFQrv
EuTkch2DRm0TPwkin2lYzYzsSQKvK5D8cmYMXAhYgwdzKLkcD45PWqEdXEMgYSLh
czygkMD3J3SrSOBvNfrysFEp71d92c2uTpdUhbqq4UnFqxxmR2yD/K5l3WBrngCo
95SWcsEhRG19PRxtVSTZAPX+91WtPtr5UD9ElRDjQYKLtRTFEtpGo0LJDzXSuVpr
uDi36X9OjoW6aVIDkI0+0cVBvBbGwytXwWseIrNaPfmnCr4iQhiuXn8aAyT9RyGQ
+MiQSrmvX5NZgFEbhcJqTTCjXokz28kORBqcl4vi/PMDavBsfBT82cnIsf502GUm
ktf7De5H8YhdRKDgUyeCdFP+2LBfWWFrci1IOz1BEFcHpngSc5DB3fzSSPkcguri
ZL8Fd3Qog5j/RRP8KgmSoqJOTkdf5VL7WTd47pkLR2XCV6terdBsRdtFkvuifEq5
Q35/eqrU47G2skHFXpn1JRzF7pISQq1g8tiZ/rVTqC3XjancJsn5w7P5ydBII015
/6QseDy/eLuxu+dqGfWvHsPIOyqHnTU4KxaAD+m0J8NHD83dZI87kOhi+LF+vpZb
3yMEGaCq3NyeQWtQS4GARAEnNWVyBcKRRGMJ7Q+YWY8qCDzoDEX200sC3REdkV2o
sCF4CA43o6Wea67nGCzFzSRHPtYYOn3EKSprZMF1Cxneg22b/LIOrSAcNJ4fx5vd
m00tRzoy/tcNzoVkbTq8xIqBkcxaebdgsHT4LyGUzaT+TCZ5TBNJsJBKoBa/tCuK
AHU71Wl/p7Z4sSKa9T/APAB6f0GpJqdwgkCjTrqLwpbQSriBdvemGCmtoT/3gGBS
8IxsDyOFGiyzoZqpL4Q3VCiDuWKbN+TIDaTT+Hj89JXqSsyRbmKC+FTp+gaWUQhH
a1sgrdCoP0bS96ydNM+OFeLa+Gt7ZX3SJ8ef5xCJONJS0SQ6dxr8rRjjnaDmgbti
znpmSUfseCvpEr6zANTs1gAaC2Oog5shZmTS6k/2y9uP+toq5vqF60odE5GiEhP/
O5jXVL7KlWkK1Er/BOU0nqfRF4qbP5I4yvlguBYDmfhHv726mYw0SkkC1GYt5ja2
30n8LULJUbPrLPVqqYLmzlLP2IaqykBnbVBxqCMziyV20x23vhLvy5vzi7YUaF+X
aO03kJu1ZyqlT4Tmt/JIYZosXQp/qZqBkKhTTb5b0zz8DGhi7aLWxI4S6tThL37G
k3Ao/SMnuWJ5yvYD2g+kz1wu9iH85Tp4qbrqrudrQb52/MUu1318gR4AE5TcZa1q
hirV9+I5PdGQbh0a34PqgxtOYiqGRv/SumCJSmsNL+8UG6cbBBhd6581qf9biXD4
3WPxHDMaC2+yXrp5OYP7u5HdEEUgpu2gw1l6ZzqCZ2i00FdWAfom6zU399t49Rvv
I6UbopZ6HrMmENDEW96CL4MdjC1SKNS8ncOE73Bg3B/cNPASgNuyqIKsW2cbqvLL
O9aBRRhjGOkU4WP4k2QSxVluIUkwoVKs8RuHLaTVkeKhknW5qt11GcKHcZk82ZRp
ggnVDs9rHSb9qroQAFiPv6gKKRplAl/Tz/NvRgVq1zjN6iqG5F14B2kE/2y5pzZS
09H0sxfXBtSOe+DZRI5D6Zr4Nm25/vdteu8cYZgWcq6+ZqnK+MoTSgRkfE+ntUjv
Fh/JLp/ZxjruanHYm6kpUHQG9oNQS8Ya+l1zXFQbO1WwgGofgU4wuJrSK1N7pefd
iS0y5QYjLBIrKp07bbMJpXEBAbgZd9q9+teXyoPEOVAon0KAuLLPqMLF1d1dGuhr
t9cxUvl+3vaaK/vL6ABmhgzfJ98MXGXhVSg/+hPebpYW5SU0vrfYqVxY9BmdsJsX
aSVeS+SzAcoPeNg6PyQQfQ/xi/XaARDLDQy4a1NzIgpXrLRI/xYsnvCR/QpBPBoq
JSf46SHvqtursouxtDCaE4s7NZP1Aok9tWeiwn/wpDDxUE7I089DLrzNfYY+uHLW
qrQ06y2gQC7GcudO9fZdzwdZ06wCwctxONwijraN4w4fPFpxYM1Hv+vs5O3ipGSx
kvKLErr5P9zltrw9dUfRu3L8PQyXgCQE9qTpaNGR8IUNnzcn0hHKOlxtsY9nyVJd
BYXHxCrkrMAQe++EiD5GLKiRH4dMDAp281iFqkPKBzmTJ9PlWp8qXU3+UjulwLJC
HlKo7kAkEMwSylI8XZDuv/Iq9Q7NcdgcTaNeAR6UKc09LspN7xhs8U3/wntlx/CJ
dDdfVs22lrQPcwCUYEjBAzuxafMzlrz8Rxc6EDLcOOunBzG1Zez9RUsowFz/kXiG
6bXuKi7HJ1MSCmoif6+tr8hXT84/jlHYNwF+cSrkDty0oMXH1jARrgfsZFaFChYL
v2st6kZKYS+y4Vm6GJQ8H6H1C5I9LVdmHwJ657ewlghh8Ck8ylZe+cAceHb8vetq
ZSZxAfSJLfE9oKFwGsPZjfebkLArX959y5tmgDCC/wX87HPQ5FLCw2qPUCJ9cy1E
Ip51gb1pvbOBF1G31yjg4pDlwoVtb+zfZLnvzebskjSdGuOZIQjRwae3hlQVFGJH
AZAAQ/No2WOM/1HLGxfD+TJuxS4L2HXrtL/Y+/C67Xp/8fXaXXeBUDh8ST91LEFl
Dt2TApU5nhmDFpc+1/TJPQzTneBhhLEMeCgi3gz/Ly39Kw8wpRqDJuZxTjibdRxn
OhUaeyFs7ID7iSKu+Ez+MkbX+6yGOh6NSVfh3t/XAMxDqwEMiHFSbHlq1AcUYPqS
kkEhJrQEm64nceFBSnKDjiyGvMp2oXH3kl5LFz0vM6HhSC6WUWdbONm1H/K9Neqx
FR/ybWns2jkk9RLpkRi6W4Zl2yERzs+mLRYO4uQc2l9+eNlJsRXjtRw4g6zz0BYf
jsYVvj+pV3u06ZHilwihJMF+LNQX0kqcoCKTqFSeqWVTaH9r1H174c7Q47zvORoY
/ir7NDRxuyITldJwHaJZ7w78OJmDfExGsV98wsddxImuT1UFc6scNhW5h0K0oRmS
tlKk993piHxAW1j0Fh7XdAiOOPggHi3jpn0c7HChSSSRF/xwfnqgoaErYD+YpnxJ
m1ot5ot7b7e6wn3tZpQjMLTyag0kQ7SyRUgzzSENuLYgIbhf7DrSae3xlHlPpSP4
jRt+LVebLVNx2UgBAgwtR1+d9pW/3EFKPO+v4FBGQ0d0miywx24tY0jG0ZWj5wDr
ob83jagpFF6cfRIozQfX864k7Q3iD1birBDZnCRtd0r3d+WRLqFm4npn+/eFspEu
rl+cOP/1YLHYUfmlBZBnx3B1NIPS6R1Qx53sCG+D1X+hlDFdG/XkwHSHcxXQYPvI
NSshOR+ca/3EBr0NM+GruRJaD3fLjtzv/TaERRT+VpETaKGZBkRlwbF1Zp5AvYbX
giQjQGbLRris3OLb/VwabVD/qM0Z/rper2hJeNFcIBwxlmoKoU61WgAuV3Bwfx0i
FRVAJB2DIxviF7T40qqM957GQlvwbQNqzGfmlbnTDxgvaYl2M/SOzwNnE/nVjdD6
RqX4M7Mfzmushzv27SN49QCbkPa1hpPs8jaSO+eZRNzalAAvP/d7spWxML5GOCXt
boorHVHILljWzVC1OGSl6TdGInv15u5svetDAcdumlcfSxS0f1ge4CfHkyFmfaP+
Z6fToUYyy16wSi5GlWZK/PPtzpNlxj6CpNgPe9rdOSt5FFRSINoU811WajXatpPp
uCq8r+IA/1CUNvfVtO0prr2zRSLdKz61du8iPgGN2zKlp9T4V8jsADWv5P+shrAK
fEXcMLkxTOFryHYm3fovKgpk3XBDC086623qqymj6mxez2VDyFPymGyOYbw8fEfg
50eCE+OxpqYsQF8cXkxauHz9nAkT08aOxevmMleB8Y921teDw1Ltm1LFj2plagUK
J0SX/AKzfWc4f3Eev9gK2UBRzUadEsiucA788GFvZxYwv1E7vBUPyGnz3cs2H/Jx
KVyCw/rfZY9bZkUrM4XSv+muGl+/Lo+BvE2gTW9d3RBd62zabmFm6B3nPxbcIvk2
wcy/0UUuvKDqhR5oU9e10/u4YhqsUxUdcHCXESwqn4Fkkli/NowpMIhfW9hcTZJk
1V2h3OZP8LfDf9sfQwVj4Z5FxxcvXqpY8FHeckS7sfTWTDn6gPgYmL81jjN84k4J
M+H7nIrJzbaq85WFVr8z4QegOtc+vX2TnggFu2yHpSBAsIpqkBGwiSOBR7EKHAtj
RHnpfQcDQ+9Sg3BaBJltxjL7gb8q1O4WRaIjN+a5TJPYRm22kZCga7gY80lqFBmW
XPdgXwjR7UcAnOeIuzMeFpy1K4hu1pge0OWhCRnYTYRdIK4/MxTPF2Wg2ix1ZllY
INmumAv/jPAfXXtdhBubEbMtvQ14gC+RXUXaIikYBpgPDjT3mJdvQIrxk0DIx2Ps
vcDUBH5As9Q3lU6/OjFAH/KjY8eGYlEz1PbopaVQNQHrpt9W5H8y7rBsCGFTI7H3
DjJTPt3zbSoWpy+fF5iiag1Bd6caCtsSSabyt2cuybkQWByP8FnCtHiSEdH+vpOH
89wrupHb9lb9r38mqK1qHO/So9lUS1NGl2VrY+HgTv18sMbR5TSArExhUjB8I62e
zcyKo3l+5SWlCQ9PwpFu36izNif21046IMsj8HrCmd4c5nehc4+/oI4gp4y35krV
xOD3FCUf1uXYLgBtxdxmfMR3tjXo2HqU8400nwKpqwaeYTOsOvQvRGce+45L4Ak1
RLxYHF/McBg0rZBvP5gS7nym2rb8bHGnzdSwAO5TcryZl0CVl04TanJSrLYee13l
vPbLCxklT9T/RrjAgc9WyEg9SbGJ2ZCzPjqLigoPCBbZze+Srz5Py5KVwghyO8S3
fmzLpKA+tjx2+fjYAKAA6in6X2WwBcspUXG/lPNXJCJYqTRHvD6qd1rPUNJ1OVpR
FdsJYGLTOJWA41Pz9WmJ4vz69iHy11E96YGG7tRPE1oQkM83NK66Nu2i8FfYrt5E
Nj/OHWSMm83gWMRcAL6CMEgX9r4rwbgwTGeacY8aQFaUnx6BAZ3NJ/Zpr7jbwlPD
lo0AIHa+9CGRUf0CMqSQ5eRP64ks9zxcEdmV2rTdMFJXuQP+h1arM2vcCOrWrmAZ
1YQxUIbqm8U2yVtiNEsdc1V5zcRBgccMe+gmdmy/m4jcIEy82K8mzFms/UcJIhGu
MO3GVKMOpQymnqBC5h3jlQUAfiiVfgl3uQICFOGLPM4PePcWhcbPBPOfz7VWUrT+
BIT8RMu/zggxAlJgxf+1oBBVTHRph3ylG3+WGg81z8BDySGo6lejk5cWmXTZnEl7
APTpVQu56vPVeHA1ey70pOuoR4OBfKc3Aoz1QjP7OakG/1ks/VprTDUDN3l4zbcR
7xDmSUjob6P+W5xJyKpcaqHilB8+wjJzJL3rtgY6+k/bodQVWvggcrAt0+NjmB8z
EHq+8CVHs9TmAh7KMUdKpBIF632l7it1SpkY745/yV+Bd/6781fAMxVv0Vjka82r
suleEzHaQyuykNci/b+qd08aw0VO9XcrcZv5ZzmnfI6+TfMbc/jNvmb81WyVYr8Y
jRKCuIGjynRZD4q7BmxsyhdBetChWMDoKOvpdh05XlC5y2XGxQf52aYu9jDhT4Z+
TpmozoOUqDA9bGkh3yv0ux+OqAC/4aT4tQkoEih9QyFPTDRLRgyeUl1UDZDhAK6p
ki1uDyhXNRznFcSmQLlovnMtFENzbqAlWteDazm94bnxgZMMNQKisn2Wj1MWW8KF
d/IoDWf5gBQszZ0NYuvTexmAhlCw5yxlqD3ZLP6tx0ZRXkmqc7pxE7EPup5RzJIQ
j1N2l8BTeFgKyv2koqQMZT9V7xUKhOpl9C7JUh/WasTh93XeHZLhF2ClLgLHp9Y3
1hKM4n6V/Tkdk62iCAqBu+0LzUoEaJbpWepRasFeU0WS9V1j7GSX9E6SNVBgemzn
I4ALWUo8z/zUSf0g5WF6+qQPt06yMbmLTh13lPP6zaU547usN1NmZQBX0qXoyS4g
XaOsYQc6sWBOQAShqSFFGSMKhHExGxrj07uG+9lFNugkTpUWahhseAUxD8COeVIu
idaFHLza+8uhjs5avoYO9yGL+NfAaYHzToI3xKIpMonrdLazeKEMTv9vbi3T3qxx
Oh6mPKFfpGXh/0VWAYGkjhbnw5WRwZ4ERpJ++Pw/xLtf563mGdM62OODX8mnz4rj
XRRqG7Dy6Kbx6/VGLemi5hdcf3A9wEqpNkFNKJwWSMwTT6uo3i1DVqHay4A1BGX/
y/kzYTb/Vx/GWHxNLoJM4bMw1JFIGfZyF7wiZWv/iJs=
`pragma protect end_protected
