// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:35:58 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
PmKQSGaoDBB5xrM0I/mdTLt3QNvTlgRblN5OXS1+bv6xf6FcrGCUBwpR6KkK602c
pCztCn7GFwF8AFpoT5jehkKkRPSTPaGahjRfifrAhtdhg1MbfryPuBjcIUqgl2Vy
Mq0zzv7q/2RHngceI41h+bJfidZNB1HUhlyZMR8uGw4=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5184)
CnZpU4/5gPc3F/dAtwtG4ts6lyqdDS3KG/o/Fwt6aFLfPsYOoTm/Lfk0QMCkypOz
Jxxs6Qw5tbglyAVIAFY1Vz+G5r5EJtxfNelSgxlxTD5N75EDnCCfvVmKXF7uZKNi
pEC2emUP90QW6UTMOGTBiYwCRbH0lwR+WmEPJu/Q1C3Pvc9twwpaMociU8Ejx12f
O2RwHx9Czt7uGOkdwtQLlOn9wvXCFPhp9KicxYgB6yVU9Dg1B2JEU5dU9BW980yE
6nF6YgtarAw18T29ZiGfdw+YCzZ/LjaQVF5BWkGj6sbqr3LOE/fGMcG3PBnVicFm
2aUOtyrd/n0EFNnBo9Z6E5nwbTL/IXU4ygKBaVq1KfSIREhCGG00ZdAPWZa5Sx9y
VJKFs4tqMT2QcrbTFNN6in4cM1Yq++LS/m7uVxzkPQnAQwjfAMUyoOLZgjcvmEF7
oxB/uFJyhoZKTKQIutjYcwTyrw45F+j8xQmQF/OmSj9ggEFSooxSkO0LKZ1H1DWp
3KS9w1qSJWXAtS0Qw3pnwcY4gKwatYP1D6pqxUglBwOEXmZMdwLarT3inZfsPVSJ
yQVJeLsGsYjLYK+0E4MNC65XtarzkOlljp8v8Gu8aOmj+8X0O4maLywOaBJVa1X7
V4Y43fBPGG+H1ImY4r3gsvvv+gZAaJrh2A9NzMvFiAfZuRb8RzValRstcwHZFGPx
1GehbVcWMqb0Ck6KJktWoAV9xWqc+16S1SElDqdaDgjum5R4aqsBUkMh6X9ukQoA
G0wT4e2zLKQlwyb83VzrehG87Av5KCx+lnRIOBjZlZKYrCFurB6T1uca/HLkOv+K
ZU/iD9u5FaLCG4ckwT4zqObBzA7FnNRIgfj5yHHZyLMsoXaPm36TYa0MEX+hOo+s
o/8I8jxTyIuOuGlYfbUNQdxsY+/7/0KEwYpiTRrK3iFzZZlNWNbjmuF4Pmlqz5Xo
LNJ6LyvhDwEh3zCQbTniXl7LHl1xPEppYk53ek0ZGWv6oUIys5i35Hj7CJNg/8e/
faY8zXE3hdnLM8DIdzkS12YJl3t8u0h7rqhJvjDeHkdv9MmIb75pOczPcnEJa3OB
T0KfKqo+8BpgiRfAk9ZRG2HkJv63Iixp1UEjCU52sdBdAtZdB8ejZ/xAlOQ9wUyw
nLYxWQ4dWLNlbgaduKUKBn/bDFdU/XiU1Bqfp7mtLyy5y58cL9xEueWCabLLFXK7
LowIKXw0E6OuE5fgmvXpZzTOumHvkM/Znq2A7KGKAvdBotIj4KJ5P2DPJyGHIFFF
/umJ8SVRfe/V1ZH4DybFwy3rH2hd2Zm/TLGnbEWwkAC1oX7hLn8mMdadG7r/ZpCe
RkCzggQcR1Ts150HDlWJi/RA5yLvKKND2CqOp69fXSOaL1uJGWxSLPHYWr13HWE6
VJ9ps7hcTS3UKdQ9dwk3NJq+Iz7NRGfO6mRjpCi+wKgx6Z0Qu+CqXixTiUQneqe0
yissWC75bYCZbapd1jPsPN1cNMB/oAGMlJ+easbJKc4njYrXAjgjnNmUkmH/unKh
QkdTMmJxftmAKTAOP9olrBc7Tf7tfYT7WsemYJWRi9hK+wt8DpqoAUf56PBgX/3r
C6Iw6UY0X5+4tw0Iv9kSEpQ2yQXAztFHXAL9pgYtZkgpa1KNcrUtqX6j2gTTym60
0SWgDuqGbOwZhom9gRUHpdm8ahBLZ8rvkBBFIY2SPXnNHjc6OUGOFw9oh2LggRXB
UguGASXWeTD5kt2ty1yzrCYEBp5HWoClnllQ8NJkp+KgGeebD625JIQNVBW9lv9f
EYox3/KLybNlLIqeZLtECHzseVgD7k1n8ai5/GqZ4A8uo0RcyfOoN7rg8kTPef0q
ybmWulOnxJLrseyQnsvA9urZ0lMfltq4gcilmHRgboJLELVXDoqrWs4Qw8+lhKzM
setPoX9tN6yBNNCsXOz6DV095MUbYi6p67B4R9LmjtU5Qc95bBoadSBpy0L5vIel
X48k7+WDciWOtdFRUspu/pJS63S4ZCKCWGKUDbwomb1esx+ADo8CEjB2nnNEtT5T
sbtCk1nP/osX6IwZn33dgZwDuf9zQvvWHtocrNnrTVSxeOwvUSMELO2SptUxENcH
6fD9wGgcaNg3P8PcBgR03hMEPRsth8/nojOBYtgLZ/iEd0m/JyLPI/F41CQNdbyv
9b9eXpyVTgwRSzNm4tqS5x4/COHshSQebIRh0MYAtaFZfT7ds3wZeqG2u2Qhi9Xl
sfvf0ggIVgPPG3MYSa+JnMd7MBI88jrjHUhY1W8Z3GcqD8MgnzmciMxi6XdHtxXd
PZs7i8Satx2rnWgt59i+8MjAGlAwMxB0S5ZAKPJI+U5HTSBvC7+sR+H70d7n8NK2
LzTVdT7eYDGzJKgsRcc6JcrHSk2bj9/MeD+ir+bxlg3rdkyCW6YsTFF6P34hrtB9
G1N52y81L1iCseT+rJlv8dlfVmXcPFGoR1bnLRwp02vM8rITbZ76i2H9CvIm2LwI
eMOgLpPUv1ujOvV/aI/FAfMSh0yCVvqkVzdBKEqFQaLDrVLhIQs+I9pnHri0p/dV
4lDYAv8HkoWAwxmVgG9O66qiFdj+RiO5f/xi+cqd0c76aDt5okUHBu54fMYoXJC3
H51mGx2G2Cg99v0UTGfOtw1e29Ac0IX/DoPdN3RiHWaE/JwHPr+ZQEwJd3dO2ZrY
C+P4PA3GltYX/UVZ3/a8CRDKpK1O5pY+Do6W+dTSLZuXbqozWAzSHzCQzJpfS74D
6uS7e1HVqnWABQ7iP1mUujFeQDlsnCQWxyqumVpd2A9eQ8esKqOrLVBnmOCmylb7
YD1xSVcSCcdLf3LZPPIID1XSiMMxj9NjrTRQiBKNPI9+1jEw6yfiiYTLL81R55Pc
SMRKo/niXwzdZrHhDxgKprR6eWJ+gSIkL7LvgTd2hSaXrVOPSreT6mBPEmdFwUuS
IUQ6f/N+qIw/AdncgmZ9IRnvD+GJNxP4M+wPg2YcbbeL7Rodchx7BkDyX8bzCIje
uGORSHOb2ctg+DA9n/ed1NUgzXLWT/pK/MPzA5rHBN/U10jhNd7zZP3yb2acXiFa
9d6laOxhPuDzNCw97XisEowc7PFj0aZJo1VEu1ycaFLUELDuV8XvohwHUWhzVAIB
aA43oS1CZfJhHWUAff6Rbxvw8D7oVxeIIFvC74QNgre82XkYs8hEKl1TdTQ94FZ/
sNxnYtEc7upQP8+9d/At+fdjikL8IGHO8FooPBnN0NXJjEryuE5JhdXDkJ97Derj
qahEysVFm/eFLAfoSjDwhMuD/U4LYZFcFopRwMEX/IfUqUizIOS7fmpedS/KBYip
E5sHALhpkSFYWni8HyJL9udnjEkuVmGeS9OvpD41oNHkhkIBfhsJwFzH/4MHwCOb
UPmiZ+WHyI/LODrlwR2a5xfGqPlahT8vXNIvGeQZxJ52Cz5INvRuGO/i8HEwYEEM
Srvxb55tQGTLmKkMSaOLlkiuSYcOjacjR8HopXcUZeQok9XuhnkApwC83v0Y4qG7
O5YgfZHsD9WxLjP1Fe6lpxsv2d0Y/UDrEFKnBJgcUT7EU97bphPpdqiKaTTKzzh1
sBmB/EuYbXgbs6pAzL5diJMUFxuGYHvNVHy4scP/R1FJcEQVfMqLyvzz9pnZng5H
9DxztaMAY7Z18tP53GJL65q8UAZhNy53iRGhcG/A8/xjVWMzYsoVdeuyAHXW27iV
GPFE7sqU4F81R78tqPYa7K4LNtUlhLgyygFoxI6g/cXjF6Vg+M8S2qGpqXAC9DaH
FpmBLPfAdeKoHRVbWYph0aCaMTsTgKPnP4LboKweYH/GFAZ2+chIQsePBU3m9vr/
b6mjf6SsO+LsoIbv98K510B00lY/YRnR72XQO6Z5giJTAkuq5Rb5zgNcJfz1rbf2
6t1t/PON9z9UVT2OxvZkubw6uAb9qkkhl7pMQysHG6N3kMtVMlMNvziPYYuQrVz0
des9v+ryLeGQq8qA+zPgaemhmqHxdfFUgohcYFwBU2uQcXB3gioGM+O4cQHRBXZ6
M3m2CTGiaACe6lSBUp550KuLbsit6rxzkcfd25akJ4oe326GtyIfpkdCmnM6UzxZ
LvWCv++o4tfUcIekTxtpQhFn8NFb8WiAYDgQGvaE/r7+MGyiDbcq/TpfAlzDRiiC
GrgwRaFWcTM/Kb68+FKaUVd9gjkSTQa2Pz7ay+fOZnYBk7Mwj8jku+GiU1J9yU9k
Pu4HZNpQKC7yjarAcE7DSCLWCIuCpmoaGcgmTv3DwPSOOUKv13l6kO0Yo/aTh9uk
XNhRs/3HdnUbxxuqe/3NEYOP8ao8D26yD3ecZq5xyNfRKrNaGE0aeRL+kIr2qafH
tvqCERC4rhli+2bS0i3FoOtZSRuKPXXNbQ+wGjldcvg3exCKKF8DvuEBhaeLie0m
UUGFqxj9KbrlXy6plujV7LjAMi8ap0ai38yoE7mldvAsI0XuRrAXtz38U5v2hw/t
dQsEchEU8iDQGI+FzuRh79oWXbCNteiLxhC8R6ceX63Pecz6TbdLACtT6sDG5Nn9
I0EoXQjI9ADuFH6yU0UHOcs3kMHdKniJwxUXjsANigGxKmXQtdshGx5sBBVEmn5z
yaToTqexVa3uQWE7RS9IXDa3YxdC/2Aq6urG1GLSlVsU+232m+5EQvKjjDONumHP
cXFsQtQNf71/xVYP43doQdP4QEfYUCCpFjW9qLN2U+6PFcCGOgCncIg/kArYSaas
e8nUC9R9rxtrQ09YG2cPOAYW3TDgxCg6Sgwwh06lPI21Oz5k1l47z7wbwd4K4vQJ
UrhRPP62T/1PlH1mfXwU3s7eMDaJd7OI2WeiYRJ8HrQ/hPwr2aRpTDCaXPh1D29O
CHdlAGEZ8XEsYX/x/wfPL3XMVV9mzwNwUi2tUMZixEwRNCzZC2uawsWjJTIbANup
M34yzTGMZxKa3n9buyONBiNdkhKeXlO+d86WLeagS+vrIkF+FbTsFMocYcaHNr+2
QrZL5cMFvRgxpjDrbgF+NB07GLIXBBoBSSuFV7wDSs+BmJNXLnCcxyedKXJRRAsq
guok8FcaJqQcsxuwZkl9OkXZh4hmqxedPjGnlKhm1hff9ay/33yJhCXp2I9ANRxa
yqUgYf+CuF4Y1yap4WJLMYt8ErIFG5fRWJh5HIayqtRcbE7soevvMK3uBuB6H0KY
eGvygH2eZtlpblkyoHotm2egdMz3kFSmkIXhgN04J/vgHa0bdbsU580KMWuD6l2f
pNim2JypTR+cn97tZ9SaB01AdNQ6mYlGVjn/hGgBx1+cnGk0X+TFpa2NnTIi+hQv
s/6NftE2n1k5SU7fNaYvAf2mL6dHXJlI9wiNsahmDwB/qm/ip6b+Q63U+d9A1+YK
QC9ALezMF95Ww8X3LMB68pejql7M9K3kLzEJZiAjH3fh9LVpbV1iZAKUdPG+cfGf
F/unsAStfAiSz8lEvWUhKY1RkiGl0nJATyrt5Cp0XTJfoLDuWeqpyIkmVP4LZurK
lDPnyOtqFzLrzo1dBFW5GB+4Srk5wrvgMDyqilTe5WRKz54JXxT5K06lM+EnoeDe
oHgL99VKeXBSC+jPL2g1Ovocu7BcGHypd5d4XnKDd4fAP3s24ZCcXO89blk5Obak
OqO0blThA1CUXP8E7K9gI7a86XCYQn1t9/cftYW4qVRKOj6qgNk5r1uSJWjZj0T9
Lev3brtqtm0bJG+n/tGSIXRVYTt+vZsCqxuFyHQaiHjxya6y9tWlPk09npHkEzDg
oviDLTbVeGelTk0FgkZW1BTPXUO0c+9knAyEak03fBEEYEOhkI08GcNLxeGDg8QI
mrJV6cYwK3TlIiykzSo79qOakdhhwfksddAj1UhpBGDQps+0frGOJpWUfn+Xkt7X
AaR4q1K3uLmbxE4uSip0xyQHNAiB3WnpiAe22kiL9Z0kFDgLIMa0yIqHyoZ22DDc
uAE2MfPksq80YSKK7o/H/7F62ukPCufb4eTpTrgrOGATk/ENPlVr8yaGNh6JHy/B
EMfSRoIMH36HlYc3UbeZ/CmrGCEoGYuZp1JSJA2o/0jHhV8zMPdkV0ZAZ/uCZM10
CL68M0Wbj1QrhYB2awdDGFMH1cJtiKtwEzMnI0Za419xMRdkXEL9JfL+ronicZLI
lgoQ7eKzg6vCB+LCQd9PrFYNREfKqGLqvFIO2D3Kr9KZNADcChcPAlONEUEOYYpT
AEjC2Hf4L+yxjWSrNx/tleYw8ukdOD+3oWPIImjSDvcXR7O/TAWZaof2wRcQqfKM
Qpio3yE/n+URpDh8DupvOCvEFKldcJe/yNdNDTwXwe7Hjds/zU9lgxVAWzLPYE4S
m6ZxxiXulR6tHzNTdFkubJGrWX8kvpv2ug056GuPZazYMyP0rTDc9eiXGJM8aXYi
vDNIHB4d51NgeNB4tR6LyeIc5rxVYq8YceyXkWGUHiXF4JU6ehmGEaj9VNsx0PiF
IW6ZzYOfBuo8r9cbyU5bowz5SHr4JZjeqJZARkLgI+moVpsV9fQPjB9mfsIWEq5U
W8USz1xzRvi7TdafMvlq05KhIyW6dHj02IDnt6KVrz2VHbxtrJb+dbLCcW2C/AT2
RKyS/vyu7CjFQwb7wIvyPUH8VSisLI31p3rvpmnd1kc936YCiDsJCPVxpRjBc3o4
e/YfvVAyeWD9sG9cIpgGNG1BJbCNog+rvsf3lqnaA6CCBpTAwjq0F+BoDFlQxpdV
WuqvhXRDWzd5Gx/RDek79dgsQlskrwtD+t8EyFvHuUbqVUaImr5QCdm8TJgdofyI
/gPyjp/KUHITxLBTnmLmOWvKXXK9VuBO93pZE/A0lH53B5lkEl+YGSoHkwXtN5oM
Z/yBaVs5LR/REMvyL3Hnf8jwIGKcGpWR/oYQM818B2f4/2tE7WEojaavP4YLi1Qg
`pragma protect end_protected
