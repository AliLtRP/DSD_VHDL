// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
OX335OaQ1o+5yzgiROJfr5Dnz2ZEyATngtROj1GqOBYhJ0jMe8sLRh9zdqPRjbOsF7Mi7EULb+xi
vctJTzJOBjxwZnbG3qteQ04KSof7hCqAU2IPO3LEOH0FColPp18sPO69ANHAtY3hrPntqVv3FBFl
cx+BzAKT+AXM5pZGeJtvRdjvzF79mCIXLOhqvHib5zJCC9NaQkm4yyjleU5ovAkQ0jwmSErbdZxN
IXGoAxtu1CTrCwgN3IhA01OS5SF2u88lI5rAWAEN3ONZr49HKa9UzPP+q6dbdwes3M/HE8D2aZhB
juxZ4rj/XCJt+UswZjIy/Z5Zl6ahu/PUkXamxA==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
RI0jrLM94rDAg4tKd/48H5zLsIsOXC3S10Y8q1odml+AbO861/fCOlyfFuCODD7EkEL+GsjrRP4h
Hvivkl2UGlXNtPZr0LPpZqstVY2pNsBkdbA2e4jiFaoNl+zjv7GMR392KOCbDxMbo6lyrL7hwZ5p
ijqEvrk+Bfi0ewAiUyU4fQVfBn6SMGOBOt+4ohNEaceVIHuycvyJyAwN4mlP6IEoKeqsF4ZaOKQq
HRSALV+kLniw5x4Fz20zx09Nv5hayWRXTVU3EGrQTAjVD9lhfUhTb9Urz/GL9mg7ahp4K+1Dnvth
kXSVVjPfGFiyl7wEQPn+XR7Gr2sISJ9TO1Ci9dWhT9acXDS6Os9mS3wtnsMIjHHQ0RpMT1ifKJ11
xW3D6K440OV+5pP8u05nUuhCopM8rptUjjNRmg8OAeztQPptm/gk6Nq1S4H5FfqN29YRO0cIolen
Xujlkzfunxgy9v4I3gB8jYHlmWadwS97E6f4PnYK8gVnKP5THev98qQK+KvRXxJYaEBt6CiQMpqg
O/HsLB8499EeYFAnBZLntYNxGdUPBLobUNLDxtVlMdnfcXO38YopY77+WyXh936mhWbto890l9Ww
8lMIy3rF7Qr30M5ikhTfno+GSirhEA+HmrRAMLOBVY7eUBvaWEZtGT8ht8AN/xU0b8QHY+TioxK9
csjvMUhFk/QIlkE48LVAZn6or111nRLgMMmvK3LmY6zhHEs7L30mHyIDx4S36gMrnyPiriIYklRS
+KfnknO1qLCGJrzFuCbWd6RbPvJgN5KTSZq+Cke0gAp1JJVask+ltyZ72/TXwViB4w9U8Of4sGEs
jpBCu/fgT44zuT31QHHNdzVquTb2Z71j6NuTWE1NqRGXcy2ac6IOxifaUM75aM+sOXZDKN/xVcZR
IeKMp224ldlzQsKAlifzokXnG5SliIsSLUKCIqhcwwb15Q8Zo3fS/sJgft6PHMlWH+p5gAJsrzkQ
JknqospJG80AclZouwzwqIm3LscjhSfrGTHkiPMhYdUceeqeUSJ5/RSb6hZk95OPBs3pKWQKSTAZ
f++dEu7GFn9YOpbQeEALehlOCv03ZdeTJHhyHRnKpDFevX0LekfzvjqQNb0dauYqgBQ6CLFp9p+P
frj7jvm/k1sL1CaWGigbTS+MGpGPtC7GPK7UbYzzZA4XB1LErwr6rMZtl2x+jgCWJCcfhTp63v/0
XsJCyHWobydeMZRTy3sqpI5f8KPGOr8b3isEtQs0PQDj+fLaWXjJJWZ/OWJ7thkqoc9n1WEnukA9
6uhHYb0e5sXD4dc3VD2y7suS+vre51b0TipW7Feym+5aAvdd86b6vup/qm1BkYRliwcMEJ7oxlWW
dbUHrcMpQkkT0qbMTfl0M9D/A1piAGOnDY+xh61y2aubSbiU7/elus++GxnXoGXoC3mxzwBc+rql
JFnDG4brZluuO6E0hFSKQV1mVpgXcLbfBQX8srIVOH8SQ34XGvxyd9LpHJHMFLDAp7mwm88gFAb5
Fk70li7MnBMbJC9A0qnPwoIdxDIS6NUOE2twzcd/t6dwR9CIzsBVYWhh6SvlSo3kml6HPzjiHJuh
1KP+YpHeuZZ52AFC7SsdSHKBfUuWa0CKUPMHxir4zO+tSGoWLpiWbmsAM6tGw22pCr/+GD16NxwM
GYywgExoGH5TrgS5db5EMWjZWgsAgVF5js4H1Ut6wkDqNBon5pSF/+b5CkXfoMgAcJkWPAVcmzuu
dxSF/BhZRD32LOG2rvNTqlkAwmJkfPRgqkgJ2tlLixC/7sPA7MpcKrl8wuHzyM4ev5RljxT/Uleh
Ias9fhknKadA0SP8946t6QZKR1xt4KPR45OOD02Z/C9GU9rIK0tB7gnqRXWVHZi4q0hrfNH2RHtW
tNINKWwytL3f6P4unv243ri3/YrnI+pUOWzN1gzTXVcpBjbL7lyQdMHJpmRxlzYp6pvBAidBrSEH
atZe8fcmYVVQNEgWdenqhsHDoKFguLObzQ/l1imCylhx4AIpAnhqz8et0oS1rZzb0di2h1K3UMBU
WO+wiEjP2ncUHc10SELVdq5oyaCBGT4YqAQWqrb2Dfxf5HaWMk5oT6W58ciuimwNQC/oB35XqzGp
ER3kxC0UXavIPaFyMXlSL4/UzGtAjbwb9BcEPb5ppEgnuUFdK+939/itBXuG+77jRQoPdLXiHiGG
7OkOY4rn0KE16oNyo3IW8/GXRfH0PX6uvK6Iz9USns6zX9bwvYM2i4+7Q6c5Eqs+X72SOIR2U6LT
dJP599zfNiVDD6w5rtTm6nvLmEiF6k/LXZRZisRVkToLvckeWQS+ZcAS/TKP3AtdAmqAtMFzfrxM
3GDOt8tRaQip49/EtoIjCebXIosP6AdgSKnopC7WQVUy6+f2I0HdJf2UFS26VsoTpjKD8znDJ0BV
BsVPB4Cs5GUzrYmUqQTbLD4Bx+arZ42Thl8drvuJGnhNPkfoPYTwSM1BoOzJyIhSPWgNpCd/pYrR
YqXHfUY7dGpn2EL12Fz9LeheRQQ9fYyuGaYFufSsYwU8CWJZWIBZ4vYLlQhHz5ny2HFO2apaMiG4
LVhZSyXTREisDLpPp0ojhB7ndZGCFycsXIGhNq0RTCXrUz6AHfgk1oEuhF7sWluT+rNuPQKbyaMG
ki0s2j7E3LvHV2LcVtaMIZkfDX3NDpmf3WKtCvAcmdGKUGe9Fxk8FkB8jj2nHNRmh2j3OqSI0pYe
CrXCyO1rWUnyBYXlBzL3Wdx7DDU/2yPHfdQQRrUy2ME3MviapXYGlF8hETF8nNl3qL0Szgs+2jRN
KPcvQbcdVD6et0xUBFcFltC6Lb1K6qeLZdWbjrxmnOu7jGj8FrwoIrT74PWQLF38FordJcMzvcWr
TkATTV/a2ILvyX9+Y9XlxV2oGlOStsO/CicFLklsbC8iWb0x1PFx7aONVc8P/NqpyI0Ab1CZZHlU
NKZrmdzXfeBwxjqc3BAQ63atximwc04K/kyvb9eT2kqmDnPYVbYUJrBVmJvZfR/3lkUQ8muDFNz3
QHqRz6Ndjc0R3eMmkOJf8BZnnrIVgVcruWdVqERk5E15zwO6jyOeU26cFVbpkMydyn72E/0fm7s3
JKY8dTEMwrpRhmzaFMHgIH2mFuO8Byn7WWWD94JRn1xoJgDVVI/VfJWv/7GtioffXMyzJhQiWwoE
d/hQXs2ny9AeOdATrAwh3GjL6I/rcXuxAlleSFnhqjmH1E55/RnvCNOh5NruWy6VbGGc2z6NHU7u
20rGgiDfb0TQl1P7I/VYzEn+MPTZLdl57BxY1q55s1UbZ5RgmWGevMuSnl7fii3ConHFU7h7SddB
jxHie1MGw/V/OOHvlSScvatGBFtai8coneQVLkNDndw8MH/GSP+317ReklCNB2IIx4eW65diSivD
GxOKZvIck5MmI3ucpSW4p9IKtM3lsfKGQOrip05owu3Lr6eny0OM57+XSyNAKK9UDouGwwq51s75
8klcAlK9QyKxJBLYz4FA4trx7/qYHUe7KwF7Qd3sDu/gQfv95mSL/Sk41g+at2NYpF8+8uCKFjFV
sEbyUywpwN+XudolztGxb9W5GEkdQLObFgjooSrsT7gUMy+fF7svPKtE8W6fr1V9vblJ1MNHY9fz
mSF/147LNzbmtBqAxghMbm/gpLTnRm73jYNZOSla8sRa6ECcXuG/hP/1sWtu6n4DQZ0HNTXj2nGC
sbhAxwEd8kZIYphWu3FJTcEWU+9Mfjf7oBpEwX0gAj/6PI4pGIpV+TaKLWOxifRdnDHFSkYZOazb
cHspLPAsHkNb3VAUaiCogC3EtEcuR/SZGZO8YV/vloEGH+wICbf5vL72EJCOf0gQTc3pacU7vnEE
mn8LiA/BcsHUSEdEqWbPhEayuExuNMPkChxHbX3CZ6jppslbQyeCqjwvNl+IXaDiQwoXFraj+juX
//0Y6A+9hmE40ntEXCdgh9rzL/A7uLTSu5wk5OQhVPwBm96oQbk7FsSUTLSC7Nm9h8XVrW0Kz7Sk
I03GRZJCbPDHJLoqT5HodTQ9lwO3RdWPaAfDmzq6uso0P2RNlkKCm8ZTTw2bqJPPkMoNQHxHbOtY
/su8UQtu51qJr9IQqqivoGjuoCJr10mpvluupzTy3TYeER/zijYMrQsEMW8JUQWHmdT/fwowWyjJ
0owKSyNixX3eGQunixvqfTQSJ3UWaMMp/6GaZTILEeTAqnsDR7omaSRhc/7lx6/2sw8s4PVTX8RA
O9zjlvZQenF+jRStvlkPYsmmUWpjq4/fKxc2T1dpYE4ui+8JRIKg86CH9YA5KPmiDmHxi92Hsfhv
TApPGLBWTg6jqkfzbpw5ub5SFAlTsxitv/rT4Okla+cSqJKeOFfKBD/TqeVjWnhYIWHF4njU7Wsz
J04N92vNnfiwtzGDrY/GxZzn6HjNqagIGmKSaILw/PgZqv7mGXmkniUxdAlYmyFqrnmUtgJbIyy5
Zjal/bZRyZmCv9XLRs84CZ4mpYsrogr9U9M5KXSqRjU77spyXRnjdARgbFknqfcpUua1Bb1DBkUM
u1e6zI7XWeDCr4Bd1DjwXNXvAbRditt3x6Pc5FnGWQAPEVU7e3sQbdV6SXtfXQaLoST14+sBCSPu
a4VQ7wll9adHyVLNEFR+Z2nKLV+ciYCdFhvX+C+iQjXe5aRjgsmNmSqE3wjTteK8kDynjDCA8WJG
jAfGvD0k43/bzMkOUnwgRe51Tf4AGjRltLNchomXJiPxyzdJUn+G7/nii2zsfmpD5dui5gdUGKWB
f9Dx70ioqYAn3EAQoAzis9ZzA4eITYMYQ2f6w4SChxuKV9M3hEBrjY8zPI0RPhvK8+M3ysb8sUWZ
2YsqZ7tjfbFf1xT3CoesBiqaUur1vJofXYVxBQ+6foQDEYSy4jRRYhcAn41Wl9TfocpFDJYFGmet
eKlx90i2JsOVu3AzJkP8bZyYRY00TjzQ2nV3uldMrAGYM4XZExhKjPY2sm16fBczcGWHGY83SRtE
FUUwXxXvXhXb1X3TntVCHJz6M5eB9BYC00dUbBi5zeGJdIe2PpfVCE/DSWU146otkWRT4lsWcrzm
Fab9DDPZmbcXTzFcTun9EdGRwFx01z+gyayirTKYWH0iREPjAtXzLL1Y8tyDc7eIZzjHGMjLpP9f
2z7VnxIH8GDMPEerClqy37OGX1PzUhMH1yr9FyJOq+KTALSDIS9lxK2YlG/4Vrelv+DhtLQ18P/k
Us9+FolB6VMjfh1Go1oehOMx63GHHXcghQKN+VNerOhCSF/+0hQ3RUKSr4Y3VNE2u4JIubKYcDUK
pApxU4KspLlK/gQWWz+uzBa//IAvSMMgQWDCweA9rh2Df5b9FNyFiaiEOMLPGkwVrdcHPnvPX+a6
mMoEzyE9qvCtC0tjH88cDt4m8TDC8IC3m5HA9+wn96AzawZnaQtxqX94mMP8Y8VVniFqcyJh4sid
+3CbNwHgekb0GtFfrZtuxQkSfv5d2XDpqoJ9SjQPaErHbUukWTyrr0lIpCqWBD8Fqm61D1YTLaWX
Ul/wk9A/TEA7dh+T4rXQlAoWbMbtM0Bzds8O7vbVeEGmvzrDMt/g76gGbOZGF6JLELL2uEXcbOPR
XAJWiJ8ECruSwYHmpWhpeiUx/roGnMy1Bl5v8YCPypC0X5RPgqZZUXFDzeNUEe4Ij8ImjqFFKuG6
7VU+JqfPlndnbNjeVlgde3tk2XTaP1mORqVNt1hY3fwjctvEUm8byOo0RTDDZaS96izw4HuPtLBL
lZhqN4mdnvY012VSKvPgj4920Z3OcU3rZSrT3RcU/dGNwkMm0YgMYQN63dYjAbXBIBY7WLJIZpGx
WZFE+1nKDS8Ve1UxL2A+xJv/p8N/jq5s3O1I9J8a4zWwxWPPytCbo+k0WQ/uKsCrT+ipRKUkaufe
RLYHF0g52S3e1gf5jXXN3bNS+RL2KOBXJg4oYEEwgmijNLOUh6hahlulhgW5CfiPS9quB66/yJre
LAgEHNflyqqPLR5XU5rnVy8kLbn9rhbZhxCkaUnkO4G+nsyjvGnhWRw2/nbTdaqfwfVnBq/DmWlQ
6RfbXrsXLvV8/6lQNsB33q3Ze4FZigNeM5BE9ji/OUPn04w8KmYhqqLL59hCbut7gEpIXs0FaEn7
bLPaRawPN35y0uj6SRU0YtAqTSxzeao/SRaRuwQugfseDaFjk5AWLuB4N3Ed4Kwu9bNwcMijUIW/
oJPd0bZge79W+GtsqKf9LJIfBTcnDTnxtsE47uqQKMhxPQcnxSf4QggNGiCtLr88d/n+bh0+GPKz
FMj4nWumMm/fbYJx7fUHXU9Z4DQGRMfUIMTAfNY9SAnvtxXBFqnNbpCQoU6qFVy6xuggLegJgOyV
GNvMpSNGl0UK1O7miTM2vznxrpsxVAt7mMxe8SmX3v3kS8Ng6g2fT1en1HCZCSEQT3+A1C2CxuSt
3mQka8OgYjZOIBoX5uquqQSYi+VCMceiG9pftBQEwqW1xHs2xnajotDSUThfGUURKdMn9lKRfx2Z
hOfnel1ab1VUaO1Dcga6qeMwR/3BaFVBlOlIv0P78gprH0RXAdvHAoKwCp4u8yHooP9nWYT46V3T
2x1ejBT7Q25LA6yguqiFgkoHlI4OWZUHVVKHL+pD6YYj72O9bB2p+r/Ikjr5b2IvdA/+4veOOoK2
prgFUjDfcqXiQFQImxasn5q4rk9IqvWaPOV0O7+FcEEZT/ZpwurrEdZFuoqxFdCQyH0yMqnVdeG0
ZQzjgCxQ9uhST+UShgy5OeScS3f3YAmAWsr64m7HE6H/4kDwl+hMXmLdjI0BaAZYWYUSWvhA5WhA
+F5uByLwD22+1COuFKCCEsp/W+wh7wT5yw/ngpnfCMy6YHGiCACUJB0Szi2xYebZrTTtK8VbUTFC
5U4/lXi2WXkRhIhKMWOwzowa0a9B33y6PzPGoRkD72lk+rAW4FVui053KsV6TEC7GV9caKETMrsm
Y3PvtgO2XEzrSE8bbK8tjqalIHiBvsvpF5SKUCHPevk4W/JetG17avex+kn9BcieCmhsHrmG1x3A
FjZg3h2V3v7KavNfPxjojyN04+rc0kDO6HOuI2iSj1OxO/R2cO0So7nwKt0k8t9JksKQZcNH+Xko
FEnK9lxCGf4/WR0xcCu9kQa47mZlyYngNgVgMnBRSRghLj7h7hzbz0OOCuWQf2+5PPfD8c4YXuYD
RAZv72Td2SVlvp6uyMnulNQAbc2DHPIp8lLxU/jgt5mu+++nnKB1IYdjYQ1GVCxVvrbw8P2ndKOK
KTHdgw+qtkOXHZ2nJliOB2fkg93PN53BsOSNiG1lkYqoYMRLlI2AgcYF8Onh29cHBr010ypA2x0+
MI5H7QXGbUCj7IjLsFEy+asw9Jj2e1r6XrIu9yY4RotMLx7H10f+fN8hiJv0OyW5d5vXszh/MNqM
cX/9eR0LIHx1t3nJWBei8N1/F069IAQufhxWM67peX8YlHFanQh85ZqVKv4+6whcaU/PvM6IheFM
7skFWx6gviC/W7YiREv6J1CmmauGqjKpcCse+LcEk1UzCDbv9nMFfDCAdHLlesL9r8GQIkBWK3Nl
GnAIbxs0+7ax3xxAxiIyz37Hfi2h4beaMFAhjkt9F66uPsFXglOvSDoITcB0pL5tVs+Q7zqhSiN+
ot2C31rbLXpdqy6KzPLK87BFFTw6U1/mGlpofByaeA/TtkWsp0RohuhLG8Bu5SRvLbdJSGwj7CFz
/gkvR3/GSdc3uKsSiQTl+4mZLGgXwfqA3mvNJ4TES//ViF9hWLH17B+RBS+7yzV294WZPTUMlIYa
wV5nrUk/RG1z/hqNNm6/opEGFIyWi4vGxdPhPcTtnzDpw8daBIn1a6/rkQ1HqTJk/Hf29aL05SNk
rAE2dHtswHoMSYepPlRR8P3OCinAWhST5jTh6kFqKBBiRkh/pevuGsbaInWFuspU1hsUM9RWha0P
mimrbx6Pb4Rza205EU6fNKRstE2JXr+E24wI3r5foYTpJPeUT0hwnJoTzP3a10bGw3iEJE7cq2Yv
j5jWCZvstOvQeRnhSffd8vjNGeNpUlHgA5AgtWP0hKVqfYC4laLNpx1ylPEIGVEC9t76U1nLlWPB
bY47jaRvziHTvuQJRyw5VkNI++DRwtEhdQBXuyqY63MjsRiTGKlomA3dmdrJlhBvZbznp5FuYmh1
rHRtTIBWVHGVAAZHrcoNdoZ1N6SPRVsZvdd3oQzvBOkiDIopNS82TgjlgOkK/oXHkfH9Y6sea5QC
sSpbRPplzunXvl/o/KVhpKO5RrVzhkZKgtd2roSgNGTK3MwJy1Bfhdn3K5Gl63lv0sh/bhb4E6d3
rZqCQv4xmg8cSM5KyT+oKfrZWQfKO3Hqy1hFzjYRUU+iM5GL3QiBmtNlBXpFjmA6F+m9sI9i4R0r
BQsBM2jr8gfr4sAGjzfvzS9usdTDbzyx/dt7/NNukzy1qLfGjtkmRin319KONgcAlywva5jtnjFG
dQzxxDGO4VeoMfUtYqzwulKokwmOku4mV5CuX0+1qioNcSRIeD08mJSB8riIabuIUeMkydy8i3jG
/u0XP6UFku+buY07tR4DuaFb+SDSzvHfzfhIfD8buLlSCdyEa8O8AalPkmbQIDSBmu7Pszbl7R4i
gcWVEbbOozOOHkkxivjmyU2MUdTN77/Pr2lr+tIXtXWS9aOgXTIgNGuIklEMuvTUJ6eb0ISkdSQj
ocUCXI61THHsuKsW8L/jL1nrdL82KwFm10AILMQofrt4o+QcFfgIlI4QfQVYcAgeWEbHq+4vp4Nt
sAfA6xyI3WzmaSDZQ8OBVDmGmJmY5O8nAyPmPHBNluX8J4rzJikbcM7C4ldlZVC2xoD9EytTnLFK
VNjpoYvSlIxlfI/UsDadbZuEQurN+8lfxEbxgiasAOcSjYEIjnDC6Wzdgq45eRJB9pm0yX+3DRTk
bpUvRR2JRiLx3qEvnXgkdcjv5Koz4hgD5CKuYGwQ0W30TDcxxTyvAtX/XFmYWRt+avMy4kSYENZt
rSb74Api6nBkvSdMdIB6xIqMpS9AcGOW8YZI7NYEfxIbMvX3UaahkjIBZ4CowS4daL6TcUQ5T/nW
nPnmab2aNH1a6XwzwmP5qFKWCI9sum1KRf/NmY/K+29lp0cUSVD9OiSLcB1PHAHPhZi58q5XKsHX
lV1UQ8c96aKMpuY4SVbEPn1BkVnROCKId3kMHOqEn8YYiVCCYeQuRnE4S9qbzMi1RqM1sxRzEHmj
85EvUGrtUVWwUWq96E4F6Zc5pGJ3HkNivZZDlBnVlxWjuUayC4lTu6yk0GMUAoMWuYd8qt4bwsRe
jQPylnmUTB0238b3LjNateQfOHn/wV0Aeromtsr/E3coR/p4eZ7whsG1e/UHIPaDmC+HW4dRLdfc
zav6rVnIgHRMp3YndgaPuiGZ3xxR8n8tCxE6skNJy8av+2nsfdQZsaR5GfNrUwArWUBDAgZd9xRm
tCY3UA0pdWRghBeul4dW6EZjjCnvgKqDgoVSQlTWbhultzaVup8oprGaEfmGd+vH3+RRcmYYr2Hf
Js0JJT326X2NR0CPs81+VN//FNoB2forZh+HVLb5idstyd55ZbJ6zOCMhMf1e3c7qXggLcY6qZOG
LI6vrwAbX6BpeEHPpNSzo5UrOMSlXLF4Ef2+r9KU2wQUDN9lgWpiM7/wzXr8hXgUVR6w4ePxFT37
vOTMnVeieRfU35K1ZQrLfNFT+kBKK6ASRqX7zomFT9HYO6b0CYyd5L8bcQfGWPFKU9wibFd/+Sp3
5gRxGxsONl6dPtc4S+I4/120gPfJqxVAqAsXIZWI+1UBhpTKAuqISgvvMitRmDG6k+GjDmiFNan6
aFZ3BElcO4h5uP6nSzhPCU6K3rqAcfsvwotPtcfDChVj1zaWf/zILrsEDgN3QUUhIOZWL+BhB9DZ
97WFn9cUAXEkpLyyTF1R5PIBkq7LcIz586X1OL3htFJaNc1fEfT2sOUBHOqLZNKmR1Mkf5suryct
INilIvjJNiQvQBWGfFyIEunoRMQFNkvLNWQPfBtxCICsj7DXLKDELdF0kOO4kzlWUz9auNj6ddKE
Mzltapv+3R9Kk5hPG0pO4xuX8CN6k/NBY1mi7CYmtlwpeuesPqxoHkwHYsoeylEcv2UdOSvkyY+A
FtqPHgr6j4zBL8zVhn48FTSOvYc9DcG5SwW8Y9qkb1tINpJDj/BviGBcZBcZGvF29Fr0xbKhGPCE
LC0WiuRVJcig8Q2AlCbCEouxWZdnzMLSG4Z5hHGwgm1ZDccrLOus/RF5VElHGTTGfQ7Kck7038wB
G/cqyGUU/53o5mxlNPVYpfFG0sgfvGje/a7K9rcvmCL4sB68ZdEVdwUUyWdb09m8+orrtTWapfbV
evJEI6BuVNnkm7wANhKgUPZVqeqp/s6rgAXZhA/islHk9O0Gb/NYLEVrKGta5MKDjEFz61+gz57A
OEAJQHVOq2kUu7yY2SIiwjujgLP0c/b5ZzvHmCF9y66qm1wRnUpVuKqV3WV8fZnUJAwzFS7B62sJ
SWjEZDPpGIX0vvcu5SwQGMuqsg4qqisPdHq/NOnQlHz0ik6ftYhduHrDeevz5hNV7fX5z6dEzYNK
1Bcaf0rP7ZIAHxOfwbRBIj56KVeMfFstqZrWnV5kjqoND5k/+93oLKKHWF5H1ydkebYTAOjgEwP8
isBjoIA//l3TCzqkGz4OHi3LRsAm17tCnqT5IcY7SK5jIrQGomXuXofqMadvtA9r6fSC4uJwQWaH
fp/eraDlBuCXPHKOVKfeKZrl5yuubGoHXOFgwkAaTwqnQA5sXRKcqbT32687YcZzuG8jaGDXCtxk
SYGRscb4vqgM/8rVaakjaBixtc0UHAq1RzZ9zvr134bTa6N6D5FibAkfs5Dt9Og/lZictLljoqPP
BJl8X1pBL68+LwTom/u5B49voSSF8Wqaw8yGT2EsGWmHzI9VcpKK2IfpchCOq8WiHcFuLjj5Ivwy
NmSI4VjhhibaoRT7w+y237NTEjinlgqgQbUrHLIfPcNErAwOP0KJpnM+DpZ4P+iaZqzU05ulcCZp
uz9WX4BgDQ7AQizEGu5oVNT0smYj5AfUnY4uCvAQGSUPrjNdn58GGE7Z71+4lBCpisMKYcUqLwUh
dD31Kwc3QXXyaeNXn5xtUZXDPWb111tUxkP4NWP0/yMcZ3VpD7ZXYSKFUfc2WjLgzZH+IIY50XPe
+M9LiIbOFhwcXK4NUhdKft4ooPyo9D10pyaWRftS7auXwCTQH1lb90iA6lEu5rOFpQnKjSxD6Fmb
VHG5S//x3YlpVyojKteGX8sbqTauwvJpskIRhpGnJlZFgbRhWeknE4P40YTtmiHD0j2mUaSc/QxM
0qvcTri8iJ+/Wv2wYn5O/rsryBm+CJd4zp9OYfKcnN3z/bCRIAe/9ysyEoU3NTNj2UmPiEtk+MJL
zMJ5PnLmAhe99zt0vYc9Mv7Mjkh7e6xP4AQo1R+KRszQBAO4/tt+fFRz7otKTn/YdLZcyYxacQSY
2/U/L8sgh9L8hG8ye8+kFHJCX8D8aXc7F4+IYwNO3SUZfby5n1TvehXoT6wsA7eejGQDg7ZDhBG+
iM1J1yileZXSkDRAQOQfvMXten1eFq3d2nnkH9jUeqch5xwsdd6cL9bHZfEYfrp3h/fsRYmB9RXQ
dqpqc9Dnge9tinFJUhyfqnFa3ihccTYQobHyeleUEwXXHtpGauOL+2yAhR8ZeTuvZIOSC5nyaqHZ
kpR5OqUMlM/N2KMlvRPud1kcg4v9xSFFh610WLSYgFO3Sf997BuwYq0dPEG8LTBIkMrqTdy7O697
b2QdBi/qn3akzFzIKu6pXLbn5R63b1kURgwrbiPFSC0hJIk66nWyCAFwPFGQNqBdMR3pfDJhKupq
CDBRj27fJObEidI5jWWVHphIcwy6hP725VNU2GKeTVvL7em9esx8UcG5VmkYh4buGlDTmCOk05Aq
z5/Awe5Fv1I1bwzeEdvtqCIccVEFejTTyGXOp9WuCirWdC6rTrtDiKQkVTx4gxw4rct/h8elHk5f
H158o4xHf4/hRSrZqMMweovBA2MDVy40vfJ7c8zLkEV04qWtxU/nAN5EGIX6IxhKgd887MEOr/5Y
r6AvXmv12LxWhjzyn3x2Hf9+JyT0IrQ4qsTicbEG3PoSbf/v+Gf1gcNln4Y3i8kYQCJuuTl4DCJ0
BhpS6PiiN15daYVXm+QGqTqPEq7FUu5lyPZGHoDHta/tDAft6TGPcvjJQFaA9bH8+npu5AIfIyyy
vJ7sDpJyseQmSDS94jag3EP7FJv/60YSXeW/v8eg5slmLAo7V1RY7hrcqN5CcDGMeMkHQnp7oGTO
HTDvPctVo2pQFi6UvVp0A7OluD4S0Un6CWjx0snkw0zx2r3iihB6WvylfZ5QbDsI0jrk2+NZP85d
Mk0X77V1qJ2ZjsAPcOYizjA2XZu1NVGL/Ka/l3JSWcrWwMWx8ijkZgjTAnN/bnf7d9P5mKR2nj2G
jbmsIS21KJW4248HbLhb4aBMR72n6KYqu0jZ1njeuONr/d+uWGMdlYw/j+tu4tYt4SMPBZZmqaO7
MtimkoefF+fS2UyfZq+rYi7a7xUnA+zbBE5r30BCdFjfiXwR4RXKC0v9JT81qIP4igDvpode9b9T
RzKiKCZ8I5uDrF9sws+CwUjMYoT3q5Nd0eee5NfoGtqUghuyPgxeDkMgF1LN1DqeCRoRCIYPIbLQ
as3/mlBzdr5HZH5LzCPlP0WSz5lXZZC/b7oPN17VzOFNrPSTj/Ae//KFjUa4BEuB6zn/C5Iamddf
mBG2UXm23fxY3SE66vGBqXogY0VL2+UcTayQ+uBgcBYMNDvFBJVmOOxdj5a09AeHVcfL+d0qNpRW
AnmPm80KZPF8milSEYxEmi9qWYVkKI9p+c4srqh7+sFuG5WkJB5Ay7mCvqSEFGyiBWQfE8KB2iCs
MBhUGA83IywIg6cxv5aeqqKY8gEz4UGST4iURnOvGwNN6u34Bqy2FkOFBcnxlrjo6dMyznDJtfUn
lWmLlLio2vriB2bUyqEJbluY5u2mO7nFvipKFsu315FwHyAif0VCEpTGL1kgwCmMFHx4jPog9RzW
MMJA0dQNWF4tDXQCXhrL8qA4f78W1rWtUjati6L8KkZfvZCHkccEE0viD4gQXqo6m13KZdcsCQU6
2sqDR4PsH/r6fIGgfais93vVQSzDXjSD5Otc/+qqAXK3tGIk9iXnT6uE5yKkPzh2R5KQxZzguhnO
+zMoE2WLm+d1SOR4xg1Uz6s/Lje3yqyFl5phSL54cDWOIiudQdE1yypOidNNBAga4c3wxnR+MLL3
Fgiidon0ZIj9NsxEiW1qDBr65CYbVdUS+Yu7XFPwXdmxFs10Z56kGQxp8gV54y8troZWHZpbfpeK
MwgZ2wEpbyF/9g389wVkmb0sOxHmCoV50HKTdx0ZnDSpk8Pr5uHNjcGQArAH6J9aVbXJunqxwHXz
0DgxrSCxfz5jS4t3RLYsPlMWh+Yv2/hW9LNyamXZyZKHoeUDLIsPtLp6U/phs2dP+8VUCVTwcbB+
9Wpap7dVkGwULTwLtAHDHN40eBp7QqxjUyiEsja7OvcKGubkXstiievz/kw99nvX+xom0ygBmNAy
JWcEpqj1ceIQNJHWUNU0sKG/o9gJ74RjpFUMycqw5+1UqZ1IYTURlWLGuUwGoUwK/xtsg9zjpzVV
Noup6S5z4FcAx7JRpH8t0gcAU/55GFai90d4UF+fE+vndt7lDhytjX6jHEjwro2LIyVaN3x9rAjK
RkJt9QdA5AHz0nK6IIEWtuaunUwoMR8EDZWUxGOir1JjcMTvd0puU179MmBG+B41cC6LOiyt0VAa
SwMEBHPjWTLCI70LEc5tHqg0SBSQxcuwylc2zOSACLW3IS+oCf4WSp0VCtrOGGu0KT1feCNN1z7+
SitCr0DEBL4BCZFF1F7sxZMRUcAtyhcq8Oq2PyZ2hjg5L/x8R8r0XdAMJV5xPkFOVO/Ug8TN4rn2
43BphAWIx+TPeSSH/rBSc5mXrgJTyKdRbQTWUV+NI/gpOY7fLAXlZa4tbk8gfzHG56csNParVOEY
CBfQOtKGo3e7bP+HGbs3mE316z3ur/rPk/egRMc8QTD5pJ5Di6qIoXoaIiXx1XjTHCJ3kEzfU12x
Av4KviJ9/yTgg9LsejCTrHeJOowOoIuSH0+NpumxJNijAqyna7rozVc4nnlETuaOBOm1GEeAE3+4
773fgDafasiCXxQ3h9NGKL+061p/laB871HBwXTA6gvKcfbKeW1vMMyaB3NbNXP7zuAUg+dDPJ5c
ZpsA6pRoTlYn44cVjScn4g2ZJ0TtKJoAw1Q4K18ZhWLznfHeLeyWmx/QeFezNjDVD3EGWgzRY5Gt
3tIMPrV+HnTqb3m1ZAIgTs819jS3KDthMt/T7nLHN7v/V5vqO8X7MfQapF8zZ9HtJPnFen0pwFEm
VCluhSSdsSCxy9qMjC3dSPUYOqIKSR0CnN/LZD0hfxgZ8G7ujgejZYK1waDGLDK+bgxN/VW4dliL
4G9eQ8DOMlxnI0aBcYFZ4P8nwgBEw/cppqIXwT+BNu7W5kYEn8+sBksoblGNEgrmV4VaDS42d5sN
+G0DyLhFnErasEhDvBmH7fTjL0jEhYy3BgHzbOUB0Fz0UEGxcvLVPHHv5McqevO4iVGdHt48ROWV
+jJZafLTJPjuFRXvpqZa1gNM+KcIeAg98BU5vk0tT3bQ7mmnHFCy1mYA2ztgahC7I2MzgKVQ/EAw
SGuplpgsa2f1pA0DBFr6eJzrribuz053B/WgDK0UoBim354aumJuDHLolJZwRv1SSV/JdP5ylU4N
P0zoUCjs+LuxA+v1awxgL5BxExk7cVqGLMiXMTNRXnQs9It9lEX5X+JDR2AydtXGonytco/LWU4H
obl/LT+r/1E9Wpp1+FXTu1NDAsEexyIfdX6WXFUlREADNEHIykAFbSXMMecGII7iMjBvM1wZAwik
uMXRgrQpkCXJFo2Qx6ewN8Wm1vUE+sEe+bIGpYOVt6PcTyPB+XgZJM46istVVbjO+F4T1SrJUGBE
aMLvEJTo99uS1SDG2GJOEsdvpWHS/Xqogwk8aHr2DgKPunwyUvGB3twKmEmuY8rkZHdJc5ETrg0+
Ou47jy3S7r2lTFuoimDeDd14xz+rC41mGSprpcpkYgiIINDEUhiL2xa2F4e4Qj1affueaL8dmL9c
jr3LnlUQip2DxxyI1qxaU0hGXnGUH8vvqmrh03G0bDc8DEDuVcKa0hgGV4RS7/bq7coJnQGVcN8g
LcEfHwPh0m+b2MLp8TueaZXTwR76ISrsvXeYGX76svDOSs6W7g/0Nx5XwqjTHVuTURP7Oelge+n9
enWovFmvPQ9dbfDrxCj9fhKkJ55Jt/vW9y3dMVTlkeSjBqkGugPaAMmxkLVD9USFsHS1d8uokaXJ
+mf1deajszzcK9hoeb+VTxB+age+RclYQCrqgQSCGl79xEL0a+gw6u28RKaG6eBWttkqMMWXDj2n
kLo+jBh5CyXuyKt/qbgQitwMJgh78QTF6HP4saOfkRUg4bhiJrNnmE9CyX6wVywvgJEVDZG6FhQl
qTZq6wF+z/tB8NQ8VYN/VRbgE3sN5rxKIuQJTXY2Z6Fi7lW8f5fHHu3nqm6biXyZfVd2Gb4l6PRc
1BgV/qkVOoneKtyR+WkFB2ELB3uU/WgMufc/prm4K3HG7HU+oiQii8sV+FlA9SRgnBsMaUYPL6/P
4fDuOVTYK6NZQcoZxXA4H7gKl5JlPS/g2d9W4Z30znTkWwQNwPMiHaVJ5zO3lKe8mwOS6GLlxsxd
K+2Nfp/YFrb54IP/Tzl/fA5wApbPJPMF1PA5MC5aiDotNbo6LRNANwqDX7JDKn+RseNx3v5oJGc4
k1iRLKjag5HDTwvETi7fsP082DEQoYzJiJs1RYA5s1cFVIVlhgvhhaIMUJa2c3ej+gC5+AWapGzI
yqKkYdtTm/znPDHScAzvw8pNp90ZY1NG4SKMCGzgP1IykZmH3wgNkKgCItYvMAIBN9vs6eYru95D
pWBTgvPAJZCkLBuBSVSy/qTEZNSjB+LMiDMWjD8P8Z6rLuNt26VF2Ol0wJx/EgBIG3C+YtuWkiJU
U6TwerdWlQNiHVtZlw7GfTlrnOFFnGkHydqwyJbahAbhaq5XixHmBEk4q/6jEVouMEjrJXJl8xlu
E8kMpnOpuCphXjCMjmLdR9z69+QYBQe6MlIRUJVt1SSKlyxNoPW5G4VWP2hsLi6XJCcMsw409DVw
wHgZPMtS/YBVFzwq+nxzRRLGt+oUlqYVvKEZWXKd6M68hwrCQ+G3IXaNfj39icCKNq+DuGhxq5rE
JiUnxh97T1qUbFvH4XSXH7aw24zRCzw0J1Ri0XRoZ593zaibTORgAYQsRtMabtWnpwe/0Vq+ybUV
1wm4g6e05OOt9hlG6C4uhxmEF36SPFR2wVKwRbJjGcYMTXUp34oX6g/vYF5qj5npYe2LHsofgSOR
e1uIbIwvOB0My0SViE1PB7vELHxYXvKqKgChzocqIyLWVzy8npr1wI1xQjwvATaCoN5G3wO1SI8o
65b4031/OzsoR+kN/XVxxY7gMFM4AlJ2E4EnVNG0XuSatwIwlrn0XStR/tiKDox6WtHrPaMqZ0t3
UPqr4iO7TivcfuEQThg0icO7RVDTCxhrtejcu+LwqC9VDvfzlyZ2WUlbsR5dyPCHK6/nXotK00uO
OwtoBdifGGhU6Ht1yswfu5U9ytxeuuN2pwoZ4TvdqoJCrYw5I8RIlMIope10rxlrCRWMRvCW6Fft
7hoo4hAy0hF9ZxnmsH/QW8WbtV7MoKcynXt4KrKACyV3GInbOx/Thx4RLMtcPrb7TCUhC9mbZQYd
MTRSDLmE5bS5OM3ZQJREecYq70Zo1hpFYZVCw2xS0kji33QpcQoYUu3YQs7IVUP4UxNiBMzuTGdf
Yw2aq2+JQCFGl/rE89C6sF3l0hZKcj8WwkunyVnCRUgSJS9GgTJLJ+EBtzOocbK2i7SAZlLKf7mj
2Fud230hMsouEgyzEQ/sOaXfcgXjKxe3KCFd/VStEWOKFRVqadYwwwftsinBfXbclz944oP7t6V/
xMu+F8WbkLcqUjA2JsdHPQ18Ho4L8qBQms1jk2XcBVGZo66TOLLmEG3kDHHkEr26HBwYelc3dfei
VzC2Tl476VaQfKUNfxjbvZoo6td8FRXUvbEzZs7IVDroqWrC65KfHHW1amVhSQWCjS6MRKPzIJ2+
nvbHdJ2wsqIaQOMOiS9BxEQo3+xqrUIOchroMidQw8xZ3niiTNWng8SCXJCKfbo1gZ1NldQgqtAp
jke6LTATQbPcSM3TsEwzgHLWSJVkH3Pk5jxmbEuG3YZNLYOEH0dA5bsMdBjpCCPGZ7T2qZU9SL4p
xljdPJqIU1F3g0EnO5vg1Ntu4hqyMWCjIYqXYsgRM4AziVAKHM+Mf3WOsV7+oaf2rIZfedaSLKCG
gkvvtM61/l6UVS6heMa9KsoVevjSngjriMj9H/+KwqUMSXMnb+ikp2CaCmwup0CLAQ6B5lmVszqi
4OkvfuN21zheOd99UlVb8iHNG5tYqxvZ3DqC4/KntmaVFrg22FVoHGFip9bHZgWzVsZTtzuNGuYY
OPuBWdtPAPVx09bigNr8H3wmX/bDHf7BnAJrL5TqioF3VRbxUh0I4S7ro1QB5xeUa8DG90e89RBW
4NfSMOmjrvkXEV4mQKuPDVxnKqdds+dgDUkgxWt8d+UXQs1QjUcAdVtUE6dMy0SKRIu0erstTMYZ
kGw6dsy6bx1gfoUdP/MP4BhFad0pj65UrUGVdstttFgkVNMAOL/WLBKyWLP9gZNUpd67OJoZD1wd
JdD8pBXpBDB8+D6lYfqB1AWa1L0XdeMUpnV6iH81He7UK6kYZdNuMOJU+rr8hsH51tzoEeeMfmFK
fbbIAoY5nXrEJmA+/D386/Y4hcXnv4//mz3NqLqyPMiXh6rTWJF5ov8/GbpiG/k/UMfeGPACkXb7
P/jiQiPATmYSLAQd0ZLrq2yiPc82nZYdDB3xMhWR2ZJ3JLMxL0NyHJVD4KinmooCb2SNW1xLw6LR
l27Zd53cAGWG33m8dNCZ0fMb9IKh90OKwf2l088MrXMGDQya8nflEmGsYlJXbYXkyXpbrBxvJorb
AWWe4bYuxglZwahRdMJ7LGcCJC+vo2IWz2J+c8n9y+HazRPrbn6bceUgyOS6lvDzS1ju+bFk7Xoa
P9suyvv65QLGFkvzjE6EJLeu3DWD5LpX6oc7bLok5vi3bVihFKG+IgKkLuUYeq+rZjiVc4rzh9Nl
O2SaWrecjtMKtEnmMa4Tey6BZZb+z1CmPfqRYaeFLMP+7GWq7UIDGEeuPtIB4onE6zxW6yVnydpb
hQ4E0GgVGuOqLvVnb/x8F1dnz8LCLSI72X1jgmEUfVXwQ6nj0TLmMte+ekkM8Xh5NnnoKUjjujx2
+xMgxcJqzfj2WvMXX0vzbB4rgI46eQCwGyVo86eLtiVZ+EA9IuZVsHCScCQJ2dozPcdmay5oUQEp
AXV2y1Zg0oUohRoJZH6aVfVZvWNUAY52TCeb5k+jdCSu6hT3OPASjyRFK7QFJAzHKeFmFpD4wF1A
kEtuFwAJgcerPnHRKjZmFjuwi2vPBw/+LLkzSmE7ztjdUifGPg0opgkktBs79H7LogORv1br3rjQ
nQ1t4ICQ1yiNG4IN2Pyh92RQpukBPPRKIYA20fjabEL2Pw5ltSDzmVaWEkGusH4XGdVruTIrtC8W
Gxl2egehm3B/CY3AXpmz55JgmZYt0eXPDJVZ6nm6uvrOdHZPJD2VgzJX76+tO6bqbHj6E0d9yikJ
CNTbOCRXAxzLd6wDerwQ4ta1hReqcIen3t12WLOoEpJWf2/WJ4d8ah8FGpmfpf3ZdwMXZN9aH6ry
Sgi+yzwm/9rfXEwPRv+2hbzICB+y75dkaWQhgr5uQwoSt9iz4lXpziMJZP2rBpM1OvIlyMCPJRPa
ZwiAbJhp2CKSbvNXdJg6G+q8JICWSOl432LCi1cGmUZ+4V9ExO0ouXwxfhjIWC25XYjjyvYd5IMQ
ZZciEiQ3FvfclqHCVhuvaNG5IMd3mZxVSC9kclmRMwu5amNl9iG6GyHdJ+6XqUABd0X9u9SfR71M
YASx3MYvwcObUlKVifMLIGa9/SrPACYhzUqZGxhpMTkAXTVg2fept70bPUZgp0Clsv0AFSFfvApf
SztjQ9r+n8LYk/nmAqneVdw0wQYaYGcEaPtZVk6El2M9ZuPgwr4/mh1A7A5QCH9XYK4yoJJIoiwr
uL6OLzKyHqmPzsTewPA2+VKkPgxNKivLviW60A3dpDcO/k01orYWQ6K8yBrTFJiimegpZCtOKId3
oVQ4a8hyLKtKInENvnXEeCmsC1HD/WJMmxmZlSCoamAfBLT1TOyxcChI+N7K8sGEu4I0WgJluAJE
AazRKXIhU2REU48fnqfBiFUVev4JCg47tqyl1Q4qdO2rPneGZkb/TBoJcArhQRed33kbPIaFmAPg
RfJIMhAeUAdCjqAKhB98M8wNc2M54geq//NqVBsXdMlF/mXDHltzqyaRYoRAoGl5gOzhPbeeS8BU
nRnevTRpyQFG8U5mdNR0bVkMhsLz+FL9WQTH1fTVUmVYICTu9JrRn8w2eMwnaBcs6iT6Q00V/Vni
6cVyRrZ0Pa0Je/gsD5fXSq/vXHhRzdlZHx1dIt3euM/L9AO7gE2WW++CIf9YW1g3GVBwsEAARbQw
A8iJoeOHXlJ0/BwgpSsWdoNNnAuhxBA5mfwN7qdc11m6IMEtpYx9myVE9U6csNaVM34CyHJacDTK
gvUZpy/0f1VoOXe5vCTS0z9cmlyBXgK9Z43ZEb0dKXSVIgRAfe0+wKTX2su7b8DH9+hwo3PP2V69
W5vU9OoqWHAHy98pZ255cjjrZHNXx89IcOXXbMM7psADtzlWL0r9ikzo896gyOeMtvvpKHm+lK4G
ajicMHKuUdc+WhZ/UJ0XvZl08pNOD5/p/aUftj47CQ+XzpPWm+6389O7sNOfo8brZ3g6GDr9Isuj
9ZZJ9r9JXoldzxpKJ64Ml/joDWHnZEAhQ6mo63ZxpAF8B+xUd10fW1KmjELfAo8Z7BUgI+s6MEc8
WpC0D8qFNvgtqbWPIAHTglGolg6SZ/6MYbDSOzLCRBL4UFP41M+XIskenZBpFscvvLg8plU9WyOy
k/k90fFg06S1JzIANJSqT3sv90ecfpu9vMJ1tzmD0DILeDca+E4irVDrN263/qokq9l7EPMIhG2h
bhZrqYHiNMSw6Ne+1Vqkr8SVWFvPIAkG6hwBXTiX0huIj4/aYz+OK7W7z9IJTeDzeKD+ntdDk3JC
cPIntrGVrYTYdx9La4G2dDqXgz8m8jRkVW/t+NxkHajXl7dyoiqIyRPl0D7ci9VT9Ss5E0nMO03D
w+reflQm2uoPKImnDehlYbKpPZ5Z0NuSD+HrnJTWNGtfkKc3Z3uNZ+M9lfZHqKjJu6QuKsZ41b3/
YIZhC6IjFvVILTCCjFc7uA/eABEbjkarYWNDw9JNn08tJbzxjZOYqcAf5DFi6uNqLf93B0+vVGLF
fOrWNeI4Gia/mu16HWrPxD2PF3ehjIjhlfnTEBx5tdmkGGBRl+b7vBFXnn11EV9DnI5MlDxYSKXV
Xt2fq88P3IZ5QqRyYcqxBYl0FGamgl/GQbG13s1wt7cbgY4Fu11vsFQ0CuOmh21Uu0YJxuUEX3fO
KsF+EErUdrpJG9h173u+JOk1XyE7MfX7LWMNJJ4qlmC+p2OH5P0u39B2oF3DuDYpMOYdO1u4uwWs
Etss08wY+JZVNsEODbHB0IHid2oB5/GnkDgvA7qx85DYv2sFzH2kMut5VBs90/RwyX01tQKHE8cR
6xhLRUUcAYexk5Nd/DcWTz7aKAM6lVJZO0fqFdBQW32L0J7IHUiAnwl0lRYqrU7hC+1BMn7GjxmC
cLKKvamxNS+hAU2bxTP+x4SYkfko6X2vbLDyUNuiUx5pjv7DVXVNKK4+IUv7DWZpGQym7BShDzqI
iyxSL5Iy5M598EZa8q/arCE5ETJzgJPXCWkgfrMulX2kIAWUwpcdwXcxLe1PnNa77iFMana72bWZ
BXnFjPB9wenp9+3Fe3/IsYOAkZw8NeKRgsWHtDgFBCKrlji8/zT7ReNDLx4q7Mn+dOUO4M7qvLbk
qbP0GWFqeNj7jwVsSFOlJlcGzwDis2PTJ1NDo9O3zrBC+zduOcWgCrt+9HamfIv/SYT/obSDstdt
PevJjVljmwX8GaJYddm6mhb3rlPJn6ohcaZiepIpLdUy3HjXH1yr7QmXishQ6oDbv/nCfZzGZTHo
p1X7aSb7Kbnneee/0OXmIFHnWfvc61XuizG/y/N75Z5uUo7IO8cXrRVW3b6dpkb3W8x3+5eNO8Kk
tKYzlAw2ITaAsOacqHd2rQmFf2taV7qTt4qrhEd6d6sSBOatYPeaDmWARACqq2XF8zlbxqXNLF/2
kAUo17J9soV2s0aWvyvEaH+jEEL62KZ8bNejktTO/UPkX5QotnPz0KL7P986mIOe48MYIE28lzLs
JkLEkJK4k6uHzNSyUGSUjOE2Kbz4RAKWejtZecvVpkfEUG3UfhNNma0sCCNaQPR7lj1ucWcaqvuP
EPDco5lWcwsJ/1s4Idm/W7hsT6twihffqbitvd1SVUUV2nMqyTkBUWVIq/Fk5la0aK6ZQLNaXkHc
F+kzzVLapzpKDOFX7buclY3Yg/gNjjg3XXFdaxiDLlUSK7A2TteqtbMJIXX+2jctDovHM3ALq0YJ
/yiSbllKG/icm/AICKJHSOs2+GToScxCh2GZliL5BYONbhS5RnV/vXtX8XvPczreV+A5cWzCKC1g
x83LzdLY1hNQn1KEZ4KWC5NBO3obkOKkFUtXrUNi3XDsLib5KV7gXncsdCKqnCQt1ipT/bQWEFi1
zZ4DTj9lUO671ptcEVJ7SbRPCcfZQ/qjFTt/LREz/xG3pCrd/NC0gq3S+fZdDyR61QunShwMHrzY
w8cPso5YHn3qwyzc5QhmvhwdHUPlZso+HkS46DKSkKA2kMWnlw7oSSRmw9+UBivUtZlhhtpXgLgT
INjyAf4wCTrikXgn+o1FVwarU5eRrzijL0xtUThNO8yuVTVJ3DgjavfqAurQfaBZj1109rAwXDf5
lyV71QiNvpHqFc6L2mY99/xtntumfxt+prJf9jtVGvAh66R2XQ2h0bSgPUxMGqKndN6us8VZ4wUI
HWYiZUxj5QQyorGYAAlwY++trrJK6qbFJNqPi36/9bGpHs+cOll5ZKLUkx+dWcz4DD3kFBpbanVN
usCwZlVO4wkkjjiud8NnEv5tXkITwA32vbpAAs9LyrvQVQshGchjvyKqfquwKAP/KOZwzW8CCKMW
bOCjNumrG3F1DH8Vspvu/3xtVfKlZn9s5lwqUYruucoDktPJ5D7oherOdeNlk10goZ7GHujONKv6
SczCn2Yy/ModKefVFpSTVsGczr/Jc5FmGQU86dZVxHIelcPlu1IHUbO77diOjU0lSAB69doRhcql
mQPpb6/FW+HiHwoyXAvtFtlEp35/JJ4QZ80i9+sYp1hXN0PN/xw4D5+wDNe19lpnvfYvmmMl8211
2Bw8WJ6WV7NlnJcdc7906j8zhDA0vId0tTf8zAdZk8cV/kCeCYxtI+c5WE5F/7q8HRdi9aEv+7a9
RV1VvdWVp3i14hrtkbwPtAYqHziWxPpSisk004IENFu39KY3C3m8syazd9WgJMEVT9GLBrWTAtM+
8wQ1xYjFbS4pwA+Wje29L5d6FaklncXl8KikGDF8tqjOO3cRR4HB8UjErjImJzXvaRrLKApx/QNU
V4RJlI18IafrRe29mkWV4F9y5LhwClKkX/+WetWMTGGnnWOQsWH58YX4xEMwi4iTTCFQkDH9uWnA
ldf1S0LR+NCFRZ8YtOZy4I2IjroJW4gk80atA9gyP/b4wvMBUeQ5PYTzNn81d8DPqLostuNMhnb8
C5d+pf4BUcSgfT+YPW/38BR8eYg4Crgjsrnhs8w2wr4Os3kD7jK3OQU9cDBZDpavChrWqdrGk4l1
vq4DFBcnEQzFhECa31ThsO9YB984OBFBMRXtck/3cyGyKQ0Z3qox/WhPJYPXjpZLVWDVM6p65GJL
h6ozqtfwR8eSxzIl5pjylQ8rV4QWRTnTcsSmpwlSQNffCKh56vdLDybDwiBkDyv+buiOAM1eJgg3
HQBqA/VYACFit6A8CpyxL6zvSgouhIcFvutl+bZxALeYXrZyCb0noSSn3CC1nRgJeEaFEXd0FyFs
wsfTwtMLGivzrgw8kRGzNHkqVZ3L8tWSU6WzuDvtT+QfMOJ4QE8CLpWeL35d/Ptzw+kvivuHDfKa
bd3r/dVAVymyU7FC1xN28XoGq1zpoPIm2QF91hCjPlwKmd0LQYx1w5ZlRszA/YcQVzkbOGcb6Qf8
kO72uurQ7Ph31TjKQJ6pavcFSpH329lw99Qg1g4LCuggS9E2Xw9+tz+Jc/j2TMNJ0KNAUkJi7BuC
ONuEiM8bPMeAlQJIeWF3TVS1rqHd8Vs1JyfUml4ovL7m4cyMQC7DMjQmTdhxmIg1WGHvIwPbmcDQ
RmyrSrwq2dVwxuPLRpRakaqCkEUZ8yuuxoxDdj2K3mDN/OlMy8TESA==
`pragma protect end_protected
