// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:31:40 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
qVgwhgH2IPufV81xR9h/tEpmJCsFqkoOLjk49r1QSymmbsdF21fIZwC6QQFlCGaP
C/ieUYsw0YF7VAtpl1EyGxhb0Zai6ykxEkW+YnjyI0ZTxlI7ZU/kIv8OMZjXXfcW
WnzJO9N9MsnqK6UxT34vGVfw0X+0+32Mgtb46cVo4bk=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 26368)
2NN0/MAPzfzl8ygAsp5IvjVoegibHqWaJlvRiRVcxxwRDjELH8rGGltJiRRhWs2Y
ZJmLOSEJGPF0dnv/alDDLFu7JvxMeGWCjHILaZG8esfRJpJZWagxkP00uqPielq9
0drneaPGiIgrWPChUQ4mtXxSMJEXY2/i7L2okYmr/Pgltxlo7FXhfbSJfNrxqFmd
zKf+aNzl+hX17pF2g8HS9cABc9bUkhnjPm96TpAaeGqxzzcm1UPmNlVFvneUr6pk
fiU8g1gsLXAUvCe9K/xndH5DenMo2MILX8nL26xbktA0Y9caDtWAT6KZQFVwhJGB
fMNTCCd+uuiRmFXHZBko5yC+rf9CqkwXFQKg+8hVjL/bVM3nVSVi5eWcLIaYS0xg
lG9hWGm7EQfRMe8Z4YdwCLD3TZeCYbp6jB1qafFWWyLZqp0mMYlgIWLnAUy0/7Y5
NICXKsxo0p2z4SJbwrO79Nh/8g+IVC5gpLg6tR1xz9Xa6si+8nMujwgvuHPliObX
pYy8l40DJ6dhbqe1ycWhr8R/eylboMnznrkH/2YChLs0eqynNAz2uwMTj70mkRCI
Skks22fFk06/L6V9IOyFiR1pvu/0dwmg8LTpWNYKS4aAqvAS/jedPDUiepU5+7l5
YNHlivghuqSysI/IhFPX2t8JZ8SQzXEcrM/FSolJfUoFHmWtX7+Cv8nP98IQu4fN
yF0NmJzrb6VwywAKlIeOjzOwr1sdnD2+ct2nQQ/XPYm5oy1Tadt0xHF+ujhYt785
uh2/Nw1AR+NyFQwt798Y7QF+rliOl/RvkdXX5zD3oXKd3k2vRB0xT7+o1UDKyecH
wocaF7kJFFkkZfJNsuL35T9bkcMELl1t46S8CLcVRLxCn9gOr7fyvYmBy18EHYZH
xvF5XqT1+u0Ymm/Ec6LABWTGdsK9cDm8RqqknVbEA4AZmKq5Z0rceB3tQiB9K4mP
CghD9fN+BLgic79xszC3EIlzYurw7JUitlPThNrtmU8cNs5bhNUr73uwE7m7XZaF
jXUSIs23FVk+aTJv4NJRXwxl56OlsYNnQVEWj0J/i10VZPZJKCpaUZ2MiHT8+AcG
y+xuEXUW2lgX/ahKzRxabBVNVCIsgiWbFDNND6Jx9EmXgbB1OqsuO57MK7frugrc
EWr0/D7ihe74rFf7aMG0lW+y8K1pH6oV4JYFWd0NrloCrsmVfn8fcYzgwrC8Q7wv
j1gYCIqDaQbVCksQA3e/atVShHm2nl/J8o7fnWPKwbeEJ3hKKeCaiqyEOWGPHlMK
zVhXq6xfVsBPG7c+xKNfSI4PTbBWMGDGEjokm1wE4fK5BlVSp1XJvnxkhWuf3zOo
XY7C/DN6SVNcpiarcBo7XSm4GNryDqJGVOatsTd2Qn1qfVJsGzUeE171xLoZ1H4D
FFKxNZdjP7dihAd6jGeL4W/yPTk17bzd7KblbMAOQxQ34vkXxWcVI+oAzmcOMGOs
KvXzmpnu6hvA0lMuDaDayvBk0dBUoXaJptqeZAfmYXsbKjS8DIgnIKfnSoDpX1Ur
b5NXLD3uzugZP6FScnPx8hPfDhhnvkiJgt3h6Q8MfuypSomDKHoSrs+bDpMBWFlW
UrYhdftCUM0iiMrYpfRLFi3zmi3x05PNVjy5t3/oiPgiRJidifsOMaB9fa9V8E5W
Dx8S+BS7qMkY6PeWnqVz5cy70HDhnnJVpDMuJLUiZbbR6srnFYV5vq+qPbMvuMgr
hGxFcoG6JNZw+YWwQ0cC2Y6dMVzoqdcx6bKSapEUg/QS2rGiH0qH4egWBuDZ0eRg
odAYZCtARNj2I7MnrDq0JCPFBlWnWufmVHCDif+6ZcA6FKHw/vAq0ZpPJDvJV4Nl
ATUTzswR7FPsZmeKyU+GcYcfDz4GrYEg4Kt0a1iEGnDFot1LUR7vP+5xhiTTaJm6
9AioFUjSxprLQs2PFCZtCgx8RMvkFlwdFesHpYHzXHJupgY3TMgIXFYaK78UC/Yz
zsYQW875UaFuJE0FI1cQ0G8z3+W9eGDbaO7fpL0cLuU1cMbAXOQr0cE9F/T73ecQ
Jo2taFhqjGVcDfyzJWL7VvLV0LtIM2MfHkvl2CEJ/wxJm0lJH/hlNQV0koVOfEVc
jrpwGJuEWtp7A7YDhZzoZvus8gfvmup9TN3nAAmThE8ulk9XE+Ktc98K/u+9jDU9
Opu/dv0eb0/Lpl9lwJg92WnCChJs9EGIxg74wrpmUzJJ06Tyrr00TEbJKXwapt75
4rCNtE+WzQ1cwpQv2Z+0DJNcuTidyPIkSLQrDIKY6F5OhIMpBhiJxx8BS7pl9GyS
Y9hnYBuqwgv8bwxvxWj/s2kpLOclPFMC4DqeNz3PNwSoZ8wkInwpV8/QPHqYeKka
/eDSqFFBaC2j2YEtqTzJM5mwr3O6JLcXI2SRRJcEKLq/39Qm/jkIe+tb8yBQ5fyz
yBPLSnv5I6kOAnhaTY4zYBacUQ7uJ3Dv3Y1bjogj5qyfkZ5/tr4ufPmPDiFFL55p
wEOKYR54kIKaIyguwO2CYg0ljbrY7ZpF+AIzNjjZ27EgqKVWfGvqTS1K61jIm65Q
MSwGUBuchSBrWE1X6/PfLahASQZWYbFxT0zNKmOjA2kAIcvn/BiPhBINKP7x6GfY
WoOPCdcUXdYKl6wgY6Bg5ue69j+5/abz9GOAlE5vHDH76JZ+AA/3A83LBqwRt4VQ
U3jj3q8norhwfm1hDvwMUFAAIstA1YLw1VsngNEwDgRZs7Zc1jZBSK4doj4Bh0jt
NajZwjT0FMUounPIleJ3/zk1myfE/5p0RFWgEIx6GIn/4j6v/JrCyEm6JOiQtNsQ
kj4+if2vOD3V+F3T+lHXKJAl0lpvM8WKgH1H8L25AOsJPLtu5+A0olm3u8lGOqh/
pvdxdtLBcLrzs/XucPXrWhvftEEckdmoTTtqtf+aRVXSwB2FwOo8AgHTu1JjFQsu
CbS1QjhFSTqkKi+LykWR/2SH6ZQpBfUZYde7OE/SH60K73tK2v6Typ+d9JijkspG
pRmrFg9hcpMniCIKOFiV7QlJsSOo9USLWSLLqvZgH9Ii8W/3Oxwuz7VY5akG1uyj
FG9nqeQKoyyAzICMeWZJlBZfN1UKJQc71e9mk4fCinKV0yS8GX3wo5VWR0rna33k
pg1ce0SNCSxoCXJTZlSpSEXYmfJqg7q4ca/uWGBCbnoe6xfDJtfygV2G5Ze/HORK
KTNMQJryVFS3vIOR3jMhMivCxYgnZo64sXsPTmdYUiaMmlB5vkUJLVPuqA1nKjaj
s4Vrmv84a/XV+M6PCpLP6mtWNgQwLTcRMuH0dIkFTTCkdrv9QAMKdnANI3F/FccE
oOJMflEiC0JHmASRJ6Ppxf7KMmrT+BQjq/5T1TOyDloNOw3Jmtf6DKycoETtx+rI
R2gNOUun3zkQqxrLesCevRbgOTsGV6h2WNhiOhLps3U1Da1InnjXpagxglIUm6Yh
kZc7aK34sadUvJVAK6WHR9sMPNANX0ww/ixV5mq5dtdvDDtaCgdm21HAATMStZ+X
Yiq3SYShx+I+7yz21XVXRKXCAjGCPYBukor73xDsO3wYJKLah4ySV+RzMG4q+Y7Z
cewlM+G6/4fAMzqtmf9s96O5thzViaxOfkaTo3E1suJC23AteT6LnHvqWwMGm4d5
kksfGiLtXmosFud1trbbdzAdezqKQmIjUWASYa6Y58DZ10H31pTxDrKQGSszdToQ
Iux5Qtp5xvPcFlPHQbTZR6O2H7w8h/vfAxSNS2tYyYHhPXQef+/DuOjTiG47l/O9
X2Dh55uI3Dj2qeG02FuUmEdQlboJtnFgwhZgyI7ixd/x7J+0S+8ZEwQpwNypTAWM
oWdrcBB6wxN0DeWHEv/t4nfiE1JtIlZPfIi+lvqXVTvsymMBf9lOGEmLEdIQnpO8
leIRZxXoabttRVFF+JgFNReb3++13El9z7gj7+asZ3prw7x/zTAvU5cZxtyHxSfC
eRl8z3IbRpytkkaAett353LmsRhJ2zQS3iraX+dUQtHTKzQqsiiM49kKwZxq/+jK
b2EjG97Pt+g605edwXRj9/MsH6rdq/wt00/vqU4jF5BaNYgLHquNeqhc/6ZrP98/
cJe/AwWie2C3315awS/D5lM9bWttImCSFZB3PclmmAVCbFVYXhrlngRwKq7XG0ak
C5tYhCuglvKwXM9elPe/qGJpbjmlZJqVxM/vvja+SJJlTdINqa4DDriOxzequ3NF
RSCtWXyCmQ5wQ4IQVvLbbBQ4ehLeWxGoFjACWdObWfYC/Z+OOeeCZajX3HyPvzyA
TXep3rM9rtnmuNi6+DwYLYQx7nIOAMSRi5rI+oVk8HoD21YdIMVM6N8FUee/39Uj
eFxN5YM+SwhjzUQfGL9UEezTRBo2A38b+8aGBrkMmmZ22BQ7XDBptqSBS67KI5Md
JflgqnbW/Asc7A/W0rXw5sz5lsgYfPnvSiCJK9Ohq+LQqc6u/KfAr1EXc6817K4n
nTkO6Z6cTPAXModzfHC5NBe2WeNGE5Gfz9J7wm3zvzjoJYpBOLiNsab7XeB8pP8/
uzgp2+Fc0NbDFF3Hkmr4FUPhj1l4Ybbh673+zbM28KtWKifQhKkh0H/+htn5uy3T
GCnfI9P644ncrgh34zSDgOzA+mgQkmZ5mHNRa1xWN4AY63XC4APiUCDI6hp3QgSu
+RkMmAopRm69W4MvcvutAvusLFZs4vh6/xW8c5kqzxwgHRvZWWXpdMIeCxHJRFan
eulnOZkvsc8bM8D45i0OTF91mWoMKoaoHKdNOIine1J6crS6yZCaXIoD2NftQ6gQ
VbChoJw7lYY4+bOKDlLQFHNY6bKsYT4UcbwtZUD/fTZZdziakDVUYNhslbSGkGDt
/qLrX072z4s8mwx/Yr0Ss0OgiXrrSb9JsjSgtuEaDAxUSLofe4FoMVoYihrwjULi
btN/X+87Yj2zJjbF8HNkQzFURCCUxWeyaNWUqTlc4+z2OQQU3wBLJN46+ap6OQfC
0YkbyOLh27P+smJGv0LM4sbpjma8SkX7zWpmW0i3DFzlNU1KanCbeGukHxPkflrB
7biJIBPCYJBKbeUFAJ0vI9zR/lmcboBqQyblNzIQQM5rZt5zh2cD91eL+JZqTyHm
520ohM1avhwF3YSRUv5Pej6xU+O9tEiP5dZDQBCqEy1PBwic4f4qEZ3UyKzyXAT2
ZrHNdoLuf75ogIQs853Z14hoQX7nTybuH6EiC1/yPFx/YJ6YG//0ksGQZ6/F00Uh
OWw9J2ZiRGSyfIMAM+pYQShgi3+RTzSTyOOme97br92+s+bIpacRaCW1ohKOhjV6
T0gq6nWBU2RD0ofPxNT4g9y9UMebGC8S+l0/+kfATzr3HtTNYvty/DGSeefvfiWe
dG2bVDcJtyY4XpWTu5jSZmV6hWDtJNm5q3dTNA+VaYUbSYT5qfw8zviiwPHDmkR9
qx5H1NxTPmwYWKbFAQWWzbG/ilxbwSc8iVK2+cXwCbvOFv0fBpXbjmqnAch8tQCK
ereiZnwi+6Ci3CT+ruf2mbSxYrNQndUiuUAlZAtNAoZ1TGml5oa2TstOsxJbhF2U
eMZxlTHFqodDVGB1c6EzzwU7//SYwzSsPw3yVb+PHsE7bdKQjuo2j/goyKNEOCIh
FBQX67nACDeR8+dee9YMKXpUPyrACurP4w7FM4DGTrrX5yaixvHmXnFYUa7Z/ew4
4duNxH2z7M7Vbvpmn+I5OwQ1/l8l5x+d0aU9lHunfABgrQPQXvPEabhULxqe5XdS
Z/4QkxoHOzkb2JESJXC7LUlJC0eGh+CSxqDf9J0SUm7vAtqjdZEPgjh+46E5seG9
fh98TTbaKdbU4r6VsQ0/kVBKJZXBQSEicVQYPp2cQ7Wm9b3vK/xjDHVEaKTH23t4
wZ7NQqWec4yAPB82/mwJL+FtqdjC1weVX/RnCKflMR71nVnrJxMsO6prR3N+vl66
lr4Ic2dfzMigoLMoEmReSFJKsBXQvITTP91g9EwrSjqlAbgVvVe/RJ/Bvzur9Eqd
oyEtXEtE92jcYXvk8c2CLwJi+sbLkr4Ewc5HGaoKiTh0/k76EUrA4WQCuNOyDsyE
D4JdJg9ZtSjm0HONR5RqxeSSSyONbmDis4Bg/6eBUYIZTD0kLjyN4hdVtSi6iIPv
EkN5qFQiL5ZpxV86yRuQex7RhNrUyV4WEaoOwHEHyJ+FJbYqb1j9D2xzGf9b15q3
7p9EMV3fp8/DX4YMOLDpQwDLK5qEQ55op5844e4pUgvbDmWHjWBoWD0DLUzMBSR6
0qcO5QaYAN6LQbBtLBuM0muzdvnj8lOhN4Y6encfJnkRlKKQwRgf1hIdFkLpmS3K
KKp2Ew35gkFZlPtuu4kka8I5Wz/013SAFOIuag3xaRPuJwI0aD/vLjsVxUGGCUkz
Dq3w5dZBVrmiqhwG4a+U6/qmFc3bjxtCLTJmSng4D4AIBkizRHBgQE/Zd3cEwKxn
iiASjVJzqCJa8aid2B3ZYSREP19Bt1hCPafuwHciGshVjV4m6Ot+cM3y0r/58/4K
/zYZYnOO16KwL1GGVzFDVCRkcxuBJMnRdIn9MQ4JjURakYUiPrlX28loOBQVqdHb
miCakLKxL6lZDptQpp9N94wCiGI3aHZ3al3gd5SEQjHBNlPTDnka5Bko0hl9pNM5
gUAK15/YrXYepKfnxXeBmWJFvKOiR8sS6VE+0SK0wnjlaOvbRbPAXLfxiQrKJSlA
8XSeISzd/8ywWSHVe55RmM7vEs48/u+xpDJOwaPxwlgnPRUegh/HJ8osH1vbZxcL
OLOKuMacuDPGe6H0S3I5wRrpfIyzACeQyqpeBz/dB4gdMOKIiSQiUxOJTWxoDgj1
j0zCwxSsP8OyQ25Wrt1i/IF6k9esV3+QuqtbvPBk159OJtNtdXcBaJCFkQB4/3D+
B2tGVew8JhlScpIwmDuWtGl/eT5d3SAxL+lFaYKYyK9oHi5kdOhV18h0TvQF//cA
RDwk+8YtyO7YrBF+NHF5l5wkMzYOf0WAZ0mfLF92uN0MYg6GjqsY49Vm54hbstGk
E81BunWQH7io/oJXuyM8a9CjkuSSZSOZ1hyQ8z/iDF0F4rTKEzB+GAGN+q95FPD/
U8d7mBUju0g+5ZEfrivTzB7T2CPAm6VSZk0oXOc2AKovsKW7/Kz6hOAzmvD97vGV
DV1l2C378Wb7DI5/PoH2FSADbPKw2fTP+0iGgjvATW13pvP2BWAyAfwTqUMXD7gx
pB4LbM/j0qSXzWKhxOOxwLHrYFjxgbiixXHwdE9Pv2/4XH3nqmrELOGhOvAkqOzJ
Km41lgIWSx42Fsl2MuckzFLEhAmViO3YxGokSKgskXAe26KSTysj41IKY3YRT2h/
kDzS2cNwnYixdIsUSDBugH1hPvzZNU6k+y2qwhJQ+VA/gFBDpDBC6Q+0rY/R5KWw
CVlD7ldDsATj6yfVE7fLzphLLvMXt62wA2r1kDq4yL2ow+fk78gBhjEZUjv3x7mE
DLukh31ywhViuvTrQZOyrz5u/pYqJwaohlKoOy35ktAUVIkxMZdO8OugYXShI8Ne
Nb7gRLf04QlY96Jj4o4ELbVKSLxqi2fLyKFbA06TnSH4FQE9BBZMhvr3d68XeEFz
osYEbcq/wsedBJEFFsgPzAMfcE4GojeEr2CuGjnPD2st+dk1H9B5vDkERPur8C3+
H7m7Xr6N7PlZr2d2US8Y5R+QZusq/s+xXc188pMQwhB7a5jL+TETFferu+19o4Xs
kebqSyLBgVgblXDJURHNaJ0QgLRKescGIV8xLHZlT79HS55UqkZtwF1YvvseUKET
HoAVJKg4RscfSHbldSRYJH9HR9clCjCRqnl2FR79eDoTpFZueMk4i6+cG8y0+srw
fwLkJ+m1xU4r+FuTd+hnSDLOtkX9lg5aVZTWeB+NqR2lRMc6cAfL/OzLKPmk4y7g
wcceN22NvqNT7pz3YYSE1vOCElTgijJK+X9KE2l6nTf4aNq30/64XdksB4ecoNtD
igTpaRq4LtcmjNCff1/pAoR8ZEWTQJqk6BECGf8dHDbnRLivjnqLqXxG7rLAwq6A
xIyMMdbsiGxTqg2xMX+tODPn5ATSiKHgXuPNDhKeEEGhZt2smNihyZDxI7ZzkP+u
mMoDpJolECbaW3ZWGQbFsfg6ahtKjRUzyKsgsIsaCuTxcM1DJKrf9swhAsJU1NXi
mSJKaRY/1xa27K1YCbHsEXfgWJ1ahBLEIYOEN/Mns5rKo9nt4e86/Es9LytPHhx5
+xs8L9vgUF8FSVEDS4z8/XozU6fjz9wl3at3jmR3bHywx1basoUxewBv4VrQRUgI
MZECNDer6bL4p/DkFaZBOeia8/aJQErqN63V4u31k+obRYy5wofLsNUnNOyrkyIZ
Y9dyNScWD+ImPvWHo+sxSW7llHsXJiUFOIQEqLIVDT2VMHytM0qB300Co0GDl5ug
nsxdklnFYZjRndibVoIzJgN+mObBaFVMgImicliWbGq75TC9PGEUhvYz9Or7X5w0
UP6L4t+n47BFQ/XvU49PyAdB2fZTQOVLcii1MB6e+IqGfgOMLEwIhYHMzAJOpcuT
VSbhZ4haDDMoi1oqk4mW3IE8nCyu+2H4/zbw4ByQ1Xtx9fuawFnngZI9p/dEMUw3
GVqh0OWBrh/YmlMfUGy6ptOPiNceirOR0q69Hetvjyu9h4smEbq0SRutCxOQ67Y/
xtEpq3l7rCa4Lx1ACOp9YJwsBaBNFakTiy/2UUOIqKSICjmuzH5a7mFfgO7kUIrx
ddpLB9RV7w1MaSPepeGnUGmW5EXpYuf+0RfM2qXmv7MIHKFXvmxRvEEBpgqpENqF
l+moAFqM4OxTSj/d9V+a+YHRJSRd6CBIk3Pg5n8vxa1eGz9MwGn0XE8Uc3/hWMnu
DBRy5azmN9APwGFPoNgepJa2ad+HvuH3pg+BN/l9FNERHDwwsXlMcPJTzY0dld4t
X9Xt4n0fhc7MMYhhzMOmJlSux3H3jZ55VekEbr8004xC3ZLoEGLD7goQZ4FxE4Z0
rk+BBC8XQcJbmMLqf6cpT9byjslm6QYvnwAppUmwih1tghS2ykQ/c99D7sbiPhRg
N7QH8YYpiquzGhCEFUKF9UtEHstBykfwcs53K0s10n6XbWqRNxb+jjG2HHeirMh4
+eglIlv85/UQC2H+zFgiWhpaFVDNWeC/xtB+raLWZUZ992MJyA9u5Sndbpm5sjFN
NZi4lbSybOaLny5++hY7yzphjVAOfUBvpvb/1WNnkx36j9eCphgM9fpbl01p7AJt
KrNbHQDZwDjtSCwZcG8/zdcf7cp+JRmq+9CkhCiVeoM26WWs1vwvdbr06QdTlzqT
Y+vgrfrRfW05gGTag7FRSOAhLsQ7vb61xo4rD1Q0e9TfK9UhorScojG4hrkXQblH
utp7IqaKPAssjch1CaYvvlZkv5zYmaOoRBXLbhgkoJjNDGwIS3s1JtSxZUAQWUn4
pFh1EpkMEtdKoEtVUybGMvwkUZ7ZKuKGce6a16ycKr1VFqhgYpP7LeuOqIVWr9yP
COjRB7VWl+0HY/siuL7P2dkA69FTR8Ko9N8BEnL+2Jvku78td2HbTednJA4iyzGT
q1jTd4M2ftytxsrzD8gL9YtaSIWv4hfV3b9wGW/x9nUF/hTquOSzfTcGKRSvyzAK
Fc0Mju0SCIiB7GMVhnMxzDFkhRPZzBCKf05Z1C/DDFpSoi250zALbIKJ0tS6LxKR
jHtI/KYrWSy1MjIc9gEuDyOw9O/ZnWhfmB7a/XC6fwcC1/6oMhNyqfvrF8xNRmHb
V/Blp+aWzBM4mT3xbxvN+drtMdOAlwMc/t+K6W+cUmh8Wr18zxb9GOhDc40OkSyg
A2VRXyTpjI0rSWVp/ro+dzZWjjACGx55zK5va/N1RUjLrDkUsMFQEP5ahjHlcA9p
rR26AwYpUy5ox/CSN8m3h6NZeEfuyTsQclxxoYVL4ecix9Vr2sfXLXCYnIFjfRNS
esVf69QJ0DDgFaBX30es5/vsYNrNTSm8huWxRTB1DBrIQhYT1djI4CrmPdSgUW26
xbB0IsZNWzMhBNUtXUp5u4jSa8DCorRlpk2UmF6zuIot90rOm3ykHO764gLBceYx
xmuD6pHYrfuWc42OMywdp3HFHjKc6GLIAlnI5nGOTNepKx96J11jOfZnleP2VEb6
7hHAvs6ue8NX8c2RkonsZ7U7G6inDG4z6q7lgvG68N1fdCAw2eukYpfUVfdGEQ2B
lVIhHDYGx3pNVHr5GO2hWLQ1+2sUUIymmFT85X25B/ecFzXbOEJ4rv6gwS+S/nB1
ag40QPiz8kp4om4+ol9cccU/6QwKLlRyfoQEp3QJXw3DR/hPN72rG/kp9B1rGjq+
5XnFo3xHyR44fIeIj6DahZQQEeKxZTig7cCH0IT/Adnf57awiWe32JdlUjUglWks
sLc2oVQkQgFre3um2Ic81RtMl7haBEpc4EeDsJSsFa46rQ4zE8Xt2/55tyIaaXlW
lXh4N9fgRQ2iXI9w9h5qQ/RNnagd0V9vAyTB4P7ca21TGgARmZoMqer+SzEWwPr1
26sYRLCZuq23HBp/Mk78csFP4ENZP2kdmWigxzxftuRmzEfSzwarf/FUgPormTys
W8QOPqxnzLpQL6A00kYCZaZ6rvlU5Xil0PpR8tlfLIzUj8JnGFNRy8dzcrpgGEHU
kpgIwk1MvOK14379MSYI6hDYRRCCziMI8ppIQZpIuOAjoeA++N5DLRTXanPI2GQm
AL2s7Ys8zw09pwx587K+nBDOpLu/1Y0Z+gqO9/WiZe2/gp3uXgxI3iaCp/WXyWPj
ciSjRL8O8LTJoDTCjIbfVA96n5DaQVf3FdJVIVr8VoCfgEkbMETri/LJpq7D0NFh
9lKeoI+PuJ8CGYv/d27BGAbtITMpiptSAo9v+/u8JBF672b+TYDgi/olD35jUtF5
1PsI7ponlopt4mHH9wejQT/S6A653WYQ0wztztD1nypPFjl3mVPtY2eaJ+1h862a
CxTm5+h08caZPkiIKCrjXbXj3GVVeT4JWPcLBexLDFq4FqZLiHY7/rP8MxDgd0lT
wW1uGSYaqD/i+PWDBNP/Gi3Gnl8irXenUcN5zVop9SJkXGk597ADdbXJSaqJ4yZD
b7NV4qXlkTMVuk1D/DJvzjNHmpsZDNExsmzveXeyqf4Nhgv3RljUh8h7TmWSXM2z
zOMwkXLnckghgXdI+msAG0M+HQ+P+PdcHAD9Ah5M67iMyDaMxLAwq8z2IrE0F7gJ
nMy1veDMvYWidmWPbhg2TfrejicLzW9CZ4pG3JklM9000FAb4CHkpXCxNV1Kuar8
v1PVl76SQceelAb8AiDBaz0EOvLGtC5002eTpWXaVg7safphwI2TsEr8CDibbUuI
tNr5txZuo/uTSGRt9AhkSK6s4vuQ3XB0kH0u9V5yoq8O6l5WmSpeZX0A+tUSXMSn
6XWSZdKwIV5a9F6AWGH34DqjDgVdgsqUQwWMvCQsgYfirErMWw4h+yNG4iFADjnY
1HN4tiw99bSbMTb1HGW9DAM8bu8gyaRL4B4lUhOh0TFIxyIK2r84Zm7CePMp3lfo
+UFSvR8jhZsjhWPdkwq3tdlWSi6y2V1fB2U2QPYJ32SRt3XFv7tVD/v7R9Z/SoAI
Aaf805dvvoVjd4qCyi+wH8IGcxu9sY3NqTWIs9jrgGETMAcd4AN2rbxQ1a63g1Sd
g45Sin2RaLkAfyz1Yla0uH72H8+GVrZV7mFLcQF4jasdkzswAFardZI4/yUm5r4P
4AnY/wPrA6TU3CxILHKLNh7TZpa6i2Vha/7yZDvH9pfpsLAMBcuGS8BSVbltZ3B6
9lKFyMo6njSC9bF+D990zzIb2HOPNeDDE3u8fDQ4a+sOctq8mqAHwDYZJQWS4yh+
qufekPAMSckOx1Ax3dyWRU7rdUYWSHVN9Kqz7wiWbmR8wsjC3CTPIoDm285loYvX
9u2/10wO2ZUXWeeVsvRdrcVAxgc1ecDDogqQbMzxcKrPRdZHLGfLtVdI++zzaQa3
LLPDI2ww7Y1xjtGw5w3qPhg4yA+q0HlxroB1aEpsxSEMNS5ox7aDKMnEEjp3we9x
x9aXpIABuQyiUyxzMBd2Ukp3fOs67oz/EKt234czjwqq4Eysxg1+aTq7ibAN9e1D
VSZe8+02QVkr4Rru8qriefdrHIqC8eDAHIY5qK1lLoS8Z0lBszC+azLAhKqrwn4d
2En6Coxt3MCKmOzy4nboUNWRip6P6h3ifzUlrcJNtBGxBJqqWtf40YbjaGLL2N5L
xSpzakkve2DbuVtsprTzvgSwoAP7lqV5mQkdFq734gOwcuYsPv3Lsy7mDNsHyizl
P3Ui9nN/B+KY3hv7RCJ6/ez27bLbPA0r9j0IVV3YYTw4uJEODuvyZohuiaK6THt5
fcGd39/9oV9dzCcSaP7Lh0PWlu6dzGELT3MRaytt+L/OkiggduY8Lw01hcLptugx
R/dByILRjKsmde6pWlaZB3B1AqklofkSOzF77QtFy26lRvwXXjO0WuikP7Md/pZ3
hCcojXo5tsFU0cNBX4vrYtxnzUpW0OSZhkzQtNZdIlVtbzu/uZZ5lSegXa3+HF4K
i/Ci8fGqFLYwFDiqKo15a5Mfl7e5f2jsw1vv2Ko76/hHJCodnLvt2+EXRfvhjt1f
KxHjqpi2rIK85sBixB/9r/1sE9PiWV2JxGe9eksx5ok6zdrEGOE9pzH+OorE+9ig
B/DLXU6LSfJgrijBgSOPFJT9LJmyL9A333oI+7Vn2ygFGRyv1OnliYP+Is75sSqn
Mo6549a21HEcoA0L/dtN8CsXzx0CKlf6GrzICDQvZQUJo7JUQ2fIkdqrA0Lc0Q4y
amg8Cc9kQnG/+v6aVG0CPw1ulynjED8KQvMCssmkZnh4OzT90yF+j0zbntV/K/d5
S+aNp2ZrKEdTpnJ8bnLLizh4QI/CesFakt0Q0okiTUE1wh0a1s0EKLSauxe6vfy8
30xP4izwS+H+f+vSLbqrVwBL7wSYkBPSoNlN5Kq3EEoYabM62cz8QjAoJfAayr/l
JaWU4qjxFgl4wBl+lV7B5n0SpQkN0jYmGkXUoyz6G/XLg1kb0gSL6HSxpzyEbmST
YTSJEcHDIfSeHhm3xAedSF8SjsEOU72i2Dy6EEVH4/5PpzzX+jZhSd+tW3DHvC0m
aE9zCKxnS9ll7E0swSXQaYh2QymDJslQE1qod//pXyx8QN3g2eivzKKFxzYqiwo2
8Lqrp15I1YgyIDY6RU/FIZoG7j3OgiM24ztenH7ndJhuap+CNOOTAMEKwxuGPwT9
hV7UJ/xzl16o1BIgTFcebgRneBEHVsF8xGsyLyrp7EHJypMjd8Bm2+lIJlgGNTOX
/aXft5q3j+KGk0bRQEtMZ2jl0mpcOfp186Y3Vd6/WAbTFkEQE8blL1Qcc7UqgaQU
dTKB4dBiRpURc/+flW80KZQ3jmqNWUD+xQ3w3g+3+cACCxvUHzt8lcztXE3GAdFO
g3y3GkNOW5cD0TREgR0UqoTgKPy8qG+DhQInXJW02Vv8aB+zS3cIFUJyQHKmG3Qq
a73Bzmb+MS26rncmV/EwG3EJHrHLIrJs3YLdoGKPzjg5mA2BaMUSbfzVspAm6EXD
Xi2o1Q1WSfpvTFRDdqAL74OALilPK2w65gyLJbGWYe3LJSrj01pSn9742c2rLlkA
BMoN/E7fwWF7SLleOOZXoiOOSzqYviuB47y/bNPyWGpmegDgQ3a+i29td3UJc8Ys
9XcwfEvV5zzjL1+LstFV509VTDC/rn1bjASlg0cG+YJVRrEelolP3buXYCsL0VQ5
sPnJBmMqQW2JXyiJfdyOdW1t3zhCQmvxkRwVjUdkfWvhfQFmHUFuMhWCxMALXT1i
CHQ4JL7USFtOG3S8qMCZmFinXii4Q211jcQTsk/qq31NxWHTRUQHcy/qCkIaTIpO
nExHtuIzwz6naJCICYI1fC/nNAvKcx0JAZEXcinFLidmT6QlW2HHyZnihuhlocTx
bXHVmTrwv8Y3R4ev39nGoFEn6lw8c4LEjsAWUXiu7//Zclr2TZXgtR9fQpqYVPUO
o+pY/BnfDkILXf5oMhnPqS6tt0BFJOxrG3xAo/uTwYqK3vieAmi0pI7IQR1SjzT5
vHsYh3drH17Q8u8ELryRZOdp7Xqww1r+qNHxJuJeID8B1rN6cyArRcd/1OG/zkEz
KZ/Nq5dHvcLC322oR2IBgLt+BbaXm9ooajTiB7e60YjLWStaCpWHrd31PmthnybH
7Z3h1lpDutLwjwgZKCyLhlmG1EhwOpGu8kRi4LDSPWdaQYSq9GzxXS1kp8ZrMc6g
v7Ya/AEjBe6xcs4Xdzy9H4eWjz5AmvRyP6U5BXXjYX+IjgTzonxuUL3ujNxmUEzV
uE2EjFlpYaehdrXLZ9tV9Z1310pwwRYd1+odFSSJj9/Q2K0vHw7ZuXMLhoJ0QQa+
VYT2xeIAxH9iKK761bMJAcxa1tT73vKRhBWLEa92wrOz7PTgAzj90WrXSXDlxSGf
V5BlpXpbidVDdiB3khoNZWpFKK2HxDgRi6CuHxcw1602Ci8UG/TwVkngUPJW78qw
UxpkEFJv5rJ1fLN8vr+jQ2ztN2GVDjoAxuAzoxcusqswNZYqdaR2Bpuw3yOyG/+b
hdb51WIrUC+hld+9MpE6jkkDUfNolHZex+1mLtQ8m95hcODy+hwOfbxTPa5z++GD
Njs1evQFWpwwDmGe5DI1nR2b5nI0l1WWQMH+pvcJHaYCdUhoT68chu3ip3XV/jy4
LUzi4qiLeiO1FCOnxE9C2MWRC08fCIizQNll26pExTWbpAnmvq4OwWwvK4q+vEx5
Op5Dq20SYKb2WdMPBBLVjzRkTuUzgmjiTDrfXE6kMJa9hjb3miePUv2w4luWnM5+
C0fJ36T7P2dReM754GErMY6BHcTFfBHTL3db2IN/kYjbuWL8jsY+U/qefnjuLMGL
dDnZwmVIc+pvmxtzKTtRivyWBKbddCME5yUpCulKOQkIWvD1Sf47adpsb9HG4qW7
6FNPV1v5wWirCIPUooJL4UvCO8FCaEuUkd1Igf8wCPLd6wOE+HW6NHHBQmOIbCnC
DFNfOWSwP7eJdsqDf874tCm2e2DHXtKcDyVLonKO03TTUcfUsIpSDxa54ZSwYozr
ukqgnrxomVtZVzUM9E6D053fmO7Cqm8227VZa4HWcPcDlJcKK+WZm8Gv0eq3mq1Z
Vix+pLNFzeJZwLqXmSW0X8TXSqXcTMLmUrmzmyUP+TVH4ylpBzLGs/JLGbQyMOks
DVTHAfXvx2LMqD/DX2ubsZrPlQVWJB3ra+iFs2c1hWnef1ola/TT0JYcC5/vnquP
yaQNk43AsHp3vIkUd2rMRDsRvZcVkFz6I75PaHjLhxT4EqSKdxP7CsV4V7wpBVJA
RUk11NYk2lgrfYF7VcYL7qqGax0WdEzWVs7SDFOjVZv8NzhNe0T4Al0I9evGRohp
TIdt8n36mix45Hzw6wNnSeI1HTpUQFHSf21fBeRwF16Ss+n8dGd1rfgJ0C9bfSPq
JMp+zPwUhn7BPknw17Ilxq41uvL4RTid6rHUyVvbd5oanm3xmtq6SKhAlVy5eKQa
ndyhouiXJgm+3aLKvNtMz1JcfA/V3gDTqg0qJkav9pZjiWfrkXNc/0DLiOtRneh0
M4R7tLaVAmTqrY9tFvw6RK3w1uNrbFF0RiTjW5E6P49Oc7bn0om5sNxnG4rkRLpF
UJ6jz+mzAH2y/1cb3pzZZXSRKEMATXI0KGXhxa97U2JnHRFebytRU9n2vgd81jc3
gItFJ5zJ9HHBC+tYSaoUrYElJuwzaAYysMk8sLo5uirGnj1pzm3xwtPBVky04Cy4
8BKiGaQKxF1KXCp9S1Vs7RdoKhtPZZS+degJyncW/ezv5p9nuM1qbbWXlxL8R9sM
dNbdAneK1hxoYe+vMQv26KBK79EVRQHcekOMRQT10FbhiZKoY+8s7tM/9aGFvEUS
nCcdOMIC/CgdSwV7crcpvLiXy4Mu1usSngK/O+mG8yQMhq8F+Yk+0pRgckc+jQEL
6E3SU+jyk6EqbZnBqTVOqfDd4xFksEnRPSq2Z5RqttJyEpKhj3m2rmmC+8cb4x7U
oNtTijO4+0/ha7RoeA/RasuyEqcP87akICAaDg5OB1VywUxF2cKgG8IENoPGGHd8
eUwfyQUFqWvGCAMDzeZ9jkrQPe26qYH4hrnSyu1QFp9xVUWeOW2Pe0SWUEG1HKsU
1m5n4X/i3aY6AIC7yRAUXVN4nU7r3j53kqIi0qRgqlgopruKYAVuXziKTb1jKc+1
7E00H9DwCxFjsyLwlWLMVWmxs7QqBhDNh5NsVAC45C21hiMXMdd7z7XMA0Oj9Tkn
fwmlKjw0YwFavMXjTL2SA3MgGGY/omPIA3nPu7Dlvjkaw4u5ZYHzqtaLCgeDqrSE
jkRMGYVOVZRBtxE1X1Hh9nssU4oLAzqXaqOqyNgSguan93pQmEVesoaLKy/kAUmj
DLpmloWIon0MQ8570yMDp7SljSW3T5ZL9xe/UCD9k2fCIFD1gXuwoemGJyXINyXr
qm0P8muSdd47H/M18iJt0XGN4QU3807K5kpc6SCvtEghhRTGdaULHVrUtYyr0I6J
Wyo8SyTPm2ESRVMLaT3h8Vl2EsMzdFT71WTDTSSWyvaAeEEXRrSYDe1cGMciLgvw
w4Pl5/FGR/k91/VkT0X6RCJztEo2DL24LxEt6DVUhN0fCm3/cEZDcitkZipBBBQL
G94DB76EUKriA343fu5UhRGy1i9nwlr1ikfM9TmLipjx2p+QgLYC2bNAZ3Jv8oVC
SfohXTE4PMZy8K4jm4cjcydGqwfAx92AWWjQb+M5vHxzwP/p8pceX9FxhPgFD5qw
1B5L/Egxmmg4OEgIM2vjg9POSiFh52v7bsmXdbo9Z4cecr4ZUdsmq8yyxHZaHW0P
l3RfUQBi9Y5Yc2ZtDzHsiIkoF8wpRq4wLw+lljr+7yTm7BTU6jfqsh4n2vaY0QEY
Mq/LjBfOMRcQf6ljBwI83ekassWspw9nOEk17yaWS0B1LREWm+A5bAUSWNMVr7i9
WQanm+O0ZBck+uO6Wv5wO2EdQ64jOHD9DYztIj7C5ZD3JnHCzYCucqjaXrCnYXfu
EFG+juxlw+hXGMWxYD7H8OeFeL5hmP+Khj3GdnZI86ft18JU+YUFfR8kldsDnDfn
2iQKFpn1mKvy4lRHUGfCY40HOloUN3I2p8mBn63LkfqDaurgh+6N+ullJGEzyihr
8egeMhPckZUOzDeQ3acVr4MnsUQCedypuTlyrrwzoFlA5mwSB6Yt03AzvjA8GhVY
9Of0P0PppeJ5nPykNN4v01i5sQd9bKx/YG/ZiRiflHaYrOHuPM5gaSiJdKkEtPhg
iRpwVTYl9XDYVQDEGTjQY6nXNrtE4T8c03cHg06UfqXCN+SMJDsBXtbBWw4++YzG
WzLPt/nq155ZJi5CbqM+EXAs2dPawaqKNPIBP7g2VWPFfcmtXXASCRX+aSw4r7g1
bZexGX2iauaEU/l6Qzzhk45nB+eKdYy1qMnlF5K7zGidtK30PsJKnuwcmqXPGSny
8W/PClFOQP/UQLRGOdSraG3O/YpK9FXMZ196z9n3Wid3UiYpwd3GFM9n1RwKr+4U
CVLb81dAcuONM/OUF00P72UuiddxxoSnOEUihhkzx/9PDl/bcrTtUil/wWHiDZNP
Vi1YxEdmp696FnaQUbDVZ7jskxaX5aVslisasRkWYMYdEFxF+ZpHp0ttgqQb0SnD
IOwFvw6ZCjF0KRMY1MEGTfpmOnAC/hIS0T1U7Et/SewZlsEGPnHRm+vbzExrrGJZ
ePBTVdlCj/Y3ShKi/EMD6oGnm2EARqEzAY9ZsAp3AciKTgyfsd0ABOzeIOqh0O57
qyS3pzcZyoTDAjEikc1Of1yQZIYQJPf60dYscI3qG6cQB4WBkpb7S+dKInAbc2Bt
hUCjAnQEWguNkMLIeKHAZXZ77rO9EMIPALw4PocFbr4gd/wtOxCFnlVEvV2B/Px6
MSIERYaS7AbPu22lsx3dDFsrSm9ZT8L4STtHw9fg3+fjGtjk1kxYI9uD2EF10UrY
Qce79jn710H9h5rU2wypzbNRNIo4eB95//rFn0ZS0k7TkLzedl4ByckYT3LyxTfs
A3Df20JaOpbnaT0UxPFQG6Ql30hgGHubHeKarQMSyTICeF7VQ9mwgZQkf8ySMuy/
qsj+Q8Iip2Mdp7RrBlNfq3XKOFvb5yCNFykOxsktxghKMtBFQdr2R9DaI14AFPID
7ibeP9gGLAKJePBe5O2nySzxqJD2TdkiJWF6BmgpEtPmcR+PtrjJfLwpK/fau4Jr
/2TSgmW5x2PzdJKvhJLLOAzW8RICxKL8GBt2J2ek6HV/Dh8/Ap8VdmZ2Zfo6aDBt
h3IPnL3gg7RmlVVtbWxulvBmj3Nkca/PQ/PWanz3Ihni0u416ddwcBFPqsfK1urS
0/XoCnLFLhc3SfBUK4Slw2sHLWat99huWulT97bs09pNC8KjFhItLuY51FaKuGLY
4R+xsDkErOU9M5JLWWkZf+HO4XtUg/F69LRIADfxpWRxUyNcpjpPdB86jfkbkJoO
hE8GZImRxUT1L2wsK6nH8Fwi/hk7z0JNEHPjB+Ei23nu7OPSlYb+iSQhWxGyMElL
rPc/bhj9os+E0gYg+8g43vJWxMvDSGG3nZpT3k94ti2mPJnJbgMw3C7rNYFvqpl/
xclQHwJOiIv7ANcF7HkpkLiPQVaNBvF62f224m6l+79rzuRt46sIeSYbbf34xoA0
G0axCADXJRlA/UGMMvB/ZL8TQ7f295rjODkqnnQImZYaJJtSdIYwgNTGIxkeL5tL
MUeMPfSVFDexp+udegfcEQP4lFkpjppTqHZj+5MpmtqgG4DlvvyFq5XfqPVy7lS7
d1x1BbE7NMrGzk8WiDGup/Qmr11T5D0K5tQnsaecY8td7+U/C+jhP6je6XIPZn9H
VFVoMqiyhytvbgaV6DkKmUFiYK7E/GRew+8q2pPIIpK/iQTwsk5XBqJJnAHCoZeU
s2HFkSeuFAtQFKtU4tePOgIbBGLWfnKVqM4a0TTeaB+w9fQ7jSkAY2mHrRtoYPqr
j/hVsUSmKuvgBfAA2s6NoGm3IKMLc0N0i7aK1Ek3Ew6M54L/DEWgNQL8uM2T0qja
sf1ZUYbTYEmWSUVePiGytcr2mzYCqtFMBespfgrlQBtLAhpbXAP+1ONiqj5/psl6
oR2C2BhAGvO8+FpJpPZFDnv+b1dY2J71dcDXUHJBcboLDVUbdBCBrLogTJvilOXE
e5Ty83yJEtZ3UtcPiflf8NB44JWD8P2k4bN5T73lLDzGiDBszSRXdH0YkP/O9I4f
VCIm+zcD6Jl836J5eX9q1v7+X/KJl7TMCM3+iX7mzy8fnnap2uB/7wnwmYp37FoS
ZJ/2GQzbCwBXmsMKp/0X2eHhVVXHfGa5w/iA6tjt6yZOzReqHIBeGI7ECR2a9RZh
RNoW8BgQI7gzGNpXXXPDny+r+9lJDOjbXprRu72V5luSiOkhMmjERvxgpyanBKXz
jXzk2EuCs6g5I/Z1mWDnDPTjG2Tr2lHFcGMnJdhcefm2ZfChFbhcEpaXkLJ3gsN3
y4/Fh7ieJu50+SIYQteSS6T0uWv5o82zyK9wyOA0AvidQi7r0QZKIvelb31CaqvJ
NW+hSWcZRpCL6te5teGfUHsdNFDjV21gfYEIU+lBHHsIFPa8O9KAxDevyKsapKJW
AlWnaS+HI2XeY0eU35WIfiIyEyn1aQW6iCiGfQjq8e/mTzofhaX48ICTLj24quTs
/iD05k55f8I0gfdFLjXMxKs3frHwYYkn42nbR2sRSAQrgY/hZWo5gJUytYPZ40PJ
wnOSFkObltXFZK0EAC0QvW738oMesawHAhRSpAVDftIeV0qHHauA0pHmb5HYzH7y
Ek/ISkvu+Llh2jlJyGo/5W42wjvnzxaUb0mbbze8hCZmDMqhki2dt7W5Xws8EozS
Bz93PBVEeHQAOHjHxmYbX3ABcnOjGbHi6lM0fZEConbhzsSsSyrBzIWt4O9yXZ7l
Wk3eW+fgw3O1oCLIUCD/nqjPeeBeapARkO/ayB0YobShc1d0Ptk7V00s7zhboru+
nnWXZqq2ArxBzBhw+lMJrbaLuYe0L9nXpbI7vhikg3smoeIMq25szdgWKYeyMk9j
Is4wB9oYAi8zmHpqCgxNvSWxkl0wr77dB4owJ9rkcAxZYkbWxi0eNpnODU2H79AO
ZZ4OlO7cs2OB3+/GPIz48nCqnZPvddqjHKM8lrooSZ6s1tcnjo8GIHNGUWhS6xi/
F0h0qZc9+PKug6eyB3w4hJXMdJyUQycbkYE7Sz4PEuxUewsJjCNpsR1hur+NaWyT
cjuLG//mXFqpDja5YqnCbpwUs7Gwc0kefbq8mlApMgSWETx9YaR0W39+uvIJdeup
d4YXgruWLzWeAWhUVkO2UInYe6H9934sM+FCH/RDGj2SFnRG/sGJjWsERisE5tK3
aE/H33Lg60d34y320gHtt9Hq1e0OPin+sIek6wfA5iKP8FGkD+upx8MXMHl1CO2C
p8n6z4HaXTo8yZebFxXTA2X9DsRzupkeP1nO5ljpjTKtfKrxzcr61BUHFxNgx1ZD
+2NU4VhDw9GXIgDGe4ZBECMfMLEKHKdALdu8k66xQ9dMvSK2/J7lUiCCUL9fth6Z
zSUkxQexW0BfzUHnJkjs1qVlmxTAvze6UP/QaHFcnB5NghRYMA6uF/QDFju/WHyY
h5aBJ0xqjy5HJPIADUz0A7hXIRu2v7CG4SglkBAKshbmQFczhXmE0MmS5fK2FwsL
sOqsh2pKDsDR7mds/aajmEfHvrKGIqySJa4b4hC9ksS03dXn/J1uqKneOO17sQM3
2VbfxhjmnJjYPd1oIiQQI5xPhXkXVGfEHn5IXbYrW3fCZq8XS2PyxG5nh1LFrrPA
68viy5kOd7koVEAVIl+T+nugfrce9yvR4dJGQc6YlOqSuuaRi1Kkj8Dm3Zf4yvEH
LgWvYbI3yx5p28rt0YBomosvrD/ijkKwm4oHcG7MXMMsKd/K6Y/eBo21Y8u9nIKo
Gw/wbXXqp0TRqcNRYA7vg2d5imVj9TVeaXD4kO4UVwcqSWz0go/TNTHBUFPcfs67
251dQkUlCFda2APEJ4FuY3yuqwehrmPewhT225r7EWcnLOKHMUuY+S1h5ud7iq1G
IbpJgSv8Hn3tphHikoy2h4uo2x8bsHE6lr0WqkJ/zxz+ShAF6KFWL8T1nmkTH6bJ
Hl+TKYiMFNLKEk20j60q8rEPGe9xHkLjIy9JOIDzguZp6OS7wuSAGKRS7CtJk0oq
tZrCfFuaokWfIy5DrkLNcdjBMoC1EoZBW3WmzmudxzMoD6W6I1mOT70DuzvJpFT7
g2sZpQsYDyeKnzamFNBfmTF61aLnerlVUe9Be7Q5p+pJfb5ii0oyDsJSkBC3NpNE
FcfQebbZcAvEkmODSRjN/f/+AjouhGO0sfryZnXYnQOPL5WXtu0JK2VsjpbTWcxV
gntiGv84yKqwPuzftMDh6jcU9F5XJ+yqnnBKulBNGnHMqpwIz4B/m72bb3J89NGq
uPa0I8YH410HR5Gp+zFEcqG2fqmO7PVmKS8mYsj6PjNP81YAswybTMTgC9igG/F8
oH8CEZ+RvkikW0ysleXiQzajVBJ3D4cGHPCTtjPfv6gU5KC38ktfvpwkfxZKtGL9
40CoXJlnOFvu8J0MijMz3jM8wHgxV7FNGoyY/EW0TxRREkFcEQYJaUcmL5k+vkWB
vFLbdK3T4ak4AiOMBs8y0AG2wd9N44SDvTMsTAjYrSZHOcY4XmfG2ssxJWqNGVvN
wA8VAH083x5vSWtQN37IcnJLXgBBgUCtr6u4StKiRWRnxQOz1mqu3+UCwUIP+GUq
XbkYprCGsSX7BcEuOdv9pleXmEWOAHSl8N46AsN7HJbK5KZFeHJl4YC6hGgcuVCY
YWA3tKVDcuUJIl9Yy9OeIukE+hjjolYrwknFqIPlHC9m7/my7bzCKKWTJQSmGT4/
OpCb5bwDVoPVbgkZnc5eI28FhZtWeSvniZLn4PjEY9CfXDiXJplaxrj14sqVqPrm
ELjzbQJn3Q6uFQ0uPInmZkfT+O9LB1FwUrb/cP6L1r/+aZfgkgpc3zB2+S3Az9Y/
CneOJftUW+W1USbXAhWY84bUe+k1qYgvVkxpt9qoDiifQRYzszXiOWlH9o/KdGGv
lbaOtkQnPmkhClDyMOL4pef7sWXeLTIKh7jiPWlCuXrqQ0rdNo5F07MSJm0dvMQr
X4VTNJFddyQV5hLYKYhIcNT0ZeYa6cp/+siTuZhB4LLYTXZ51RLHOBD9hF60Da3p
0dPoUbEIgh8765PrHa2gFLtBgybwi7VPXvhlQfz7DbzTPAcBVWqbGmsGfyC8670A
dRVyqE1IMOWUaFaMawKtOeGidSWV1Iy67A091WMYaqF8vs6cCH4YEktHal25pwAq
NmicI+gKUDAJD3F8kJ4vqFObTXAOFt232NBVGAeJRE2Gud9JMz9Y/Fi5GMofSqNM
Q5SIvvqSPddVhrupI2bIP1YBGdyBD1xnl5tFW/3OZGSi1uDVAbZuUCJ+BUOiWBoy
nt3lv0AIej8tDfx0MlQKzH9lu6swmUYh7nagjtJ1JTuwBsJ33jJFhTx3c1kBKu3j
txOu9EHmOycsa5cfUQY7Nn32eS6UdHDp/YXG39VKsw24dRhx1XO/bRuRV/qAwS2D
M5fupZjzKALVc2/HuV/9bduqAr0aT8JPX5CYulkdOve3yQSKoXs6tCTdEJYgxuKJ
S+v/BiSLMgE8UwjYX77TvKlEpLtDrztFRE+6aDSSVqpMd3kW0VfeK5rBY4w6uTEB
yQdKRZH3C2y8lM3fZZkXdtCAku9RwdrpiVMn69pr9c2T3KDKwBPUwBanq9rHUYpc
OgalzY/1LHAE4/CBzJi/mXMjy+KD7V/sWGKMtf6aj2cRDzHV14mlYudrHvkk1EnZ
JeuPuvZdHWjrIsI9CxKs8wRSgfPm1zHJE+rUxolUWVDIJCelJYA8QiTd87WE1L4/
EEjhyksYuiLFHIDJSwJ6KmnGBXZ2lTk2ZbrGERuTJF9vZ+MCnUZrJEPlvzJXVHfh
TrAgBSlVtAwu6GlPDCOFJdyWXXwCIl3CVOeuC/JjMqZOdxrOmArE1F7dBUoIQrqq
JHM3y6Ob0eDmtEmN/PwXoSj+mRL7neuYdHfJiZOo/vDFpglP3HhuqStrXbDzFec6
aBxi2oZSojPY1WlnURbuFnXEKlx3OdSf9M5xIgq/bWpHW8CJuLVUXgIIDu1Mx8Vl
7G/D87FNM8QyzUYRHBqj5/uykK80SR9BUwZX9/T6emR0s92VTNwttHIE44N/88dX
LNQM7OQKxedY4ecINPQ9RCuh4P7WCda3pXew9GX9zxmRt3qGh5Gyl0Z4Whf9KwPY
jh81MxSnWqGTwt24geTjUWTcY2maneRTa++D3hj7r9A/aSDzdScnDQ8OAngxC7IL
6mjObIYIospQ3h5d6anecUEO0nKYNV+ta/UejrS4k/GIN74LsalppawvSGincKFC
5ArlRCbR/+c9AVe1OSUE2tDP1PHeL5GmJmak2qLEutkgM2i1e7451vGeqEedYgsi
rkRj33IlSl5ujjSgdQnOS26vigEcu9sD9VVHf+SzBR0yA6BrTM07bzwgnvQbgbxj
N2mjsaeDvOqQBOjwdWjaPLK7eNHO9ZA9Xj6tJEj+fvj4Da9zU4oqVT7oG5pi3iVx
QJkQBu9PdVso4/sQn7SEU7YugbxnV/buPjSYawSyfG0O0+kktuP702Xpe1fdaL71
NjurLP1kDEpTUZZHcNkgCWhpvsf7M3Y8ioeGLkSa2UPlW5xEbhkA6SucKE+JYmyy
cTn+HNyuMVeDJVFr7BgRxxoJ3z3ihIxMN3QwMUUWLGccYPVMgBMjxaCXQxNmL7K/
zsh3b/hxK2Py/M4haJw861Ix4qtCelIjsitqxlor4CQa50ODewp1XBiB8yccFiYI
e0v36oew245cKTs9txiBaQGvndnujCGE8CdvfzH2sWGRX+hnrm1/6YWCWREEGi2l
fZDXA7f1SQPW9WAHkxNhCASVzQ313yVePjZZVQmdnys4lgsGLqL9NdhQuoxvmBUo
GsjJXh8+vco0jWY6FR8VD97u+m/f2UfQ0vTq15bEREUGck+z3CjAjDDrns4+aPdb
cEUp4QJJjPx1d0HxJpazUYtjRUzGjk5e2UdELDHaXbMcp2iWZeqOvyHkn+hu3Y2Y
5CsyyGhiFUuef5qOJQ1U0/MKLdz2wPhN/Ad95cb54TY9B64hJSlqENnDV5To7zyx
DPMzo2UGs2ENyLuSf/Q/ndWXMsJoGEqZ/higvkK1gCWowWMF0AAZrYIlbod009k4
pZWRExW+CheNbSgT2CmoxG28I5L2N7Q4vF/QCTnRMND68wpV33iiLwDAonpwWIE6
qlt2eKYxr7pguFkmDOORHl3mUBGdvyXVoWJjKXxActnBTrpNFIxf+RG9epd3Q3IC
GJ0HXUWsxv0jN8Eu8xzy7q80j2naB3hZx1Slb+qRpJ0VW3NpaugSNCJv+eLh1sCW
sUvgl1oz7hABjxCq5Zg4hEJ+/MZJbCIh3h+1CNwsJ9lIXrjnbXsSJ/pGfjCjWPax
11c4Zjj2Sm+5unAQxRbb2mm0hye18Tt2qvtKnqjSBxy/b8Snyw0BY9ZirQTC0tff
HUORz3TyNrhAhmBHCR5k5JhdubA2uCa9tF+Vb+tw2+fqPdiQOVFKo/wcIGdLsBeP
c97TEtpNnkt/6jQGyujl48DPT3Kbmq5yvWop41SpGepHk77EXH+Nj7zGVB1Og6X3
QaKZRmVmw5zyi26/n0Ro79YwcBF+7Q6bnLK1bEc+dfr0oFaoxx2JFxVGBWp5dUiI
Lv9ElBiR86ck9Yi/r0V7X21EhYntrGbgAu8Wc9by1aHkaPBcZERCbvRWVdl8pUOh
oJW35m6sAC3wkLfyNAhLW1mw7D6ybBxkxvOaEyQpVtCPc+FQsNDlM6iiBn21NjyY
EHYVqBgHV3rKKEoTS3YcBLokAubtuH125WVe5uJFxYchaJknF0ZWmV29FGdG2GM7
AZoBhIHKaMRmYe7HthtRHFvUlQi6jJhuqX1o0PjNMch6quWY+Rs9bvlJQxGmWSgT
gpcNFWDvIXafXqzneatCE2Zk6XWxjp23sy58l7Ii7bAt4xhaZ0/72mJcBrTU8Tjh
xtrDo400z0/mCEDQ6MHVkOtsoSVjVc6eXeZD5JRDl+Qlc1vOIqLMS9/sSR98KwTu
2L4hs2R4jfvUg3ZaENjumxtziWR7erqt/7fqrmLIyOLaXSBE+tFhV8r12Cy8r5ly
tuEqVmND6DHCI3qJfhZUWhNc/XgTJ4+ZwYYOQORN1m/11IoBTb63S9SjdYylwKa5
5MS01hWh14Y2XKKap0cZJL5xynUiTcHiQZCuuaJpzdrWe/Msp00SLGzXPufvV4JK
N5dZ5wP2vFA42ybqXa9ixEPhloZOhilqpZ0+fAAFfsPIVYGFR+sfHVd5TJxXpyS7
sgZs/lD/sT7jiurgYYkxGdCxuC73VTw7vF75utQX/VINveqZrA7ev2G+RP2pWYfe
0GQ05wACttJ/k3pxFWj5DBvpTCxXkEcdoNDNRaxauzMRhewSnyt7yf2qeJaO+xuB
C4VMKKShcaBfOj1m5GPIEqn1TjGEWKaCu/BUOyJ0RGOFeQ8UomG14IrlYMyBxrPH
eGpK/7U33h8MnsBV2TPXcIyiKnZcSiCPjKBmRdUk0Wsy5rVeisXjAa2DpSp6yDFM
xeqDXf2fhKSlgNU7bLKJ+cMvloNbkxCMy7zjJzG6pHRX74jgSf3WUOEIyCnsEpUF
4YfHZmKIorEJmi8flj5kQu6GgSM0IEYAjFmRJmOdbPPehngz9jTJtwFcsumlgsd4
tIXt74dNIijBuF+yhnTFTdnsJvIgEcJGuCEd/VmEXL6lt9gXVpQl9K6aLIYnclgn
ukDWnsVlEBDtABG2ElFYtlIkJLvj2LxOCae2pTuaN/0hq1SYiGpiDl0QIPLgi96W
wPbhfkuaeYwIMJkCuxbe9LVKyC2CvF0zXND7pDHkCD7LOXNsywB8w1as6rN6G9hK
JiMs4x+7fv7BKG/fe6cE0CfryB8/mzb3fX18aUi51C2H20qRfJjQvnNk1dc1395o
mfBm81xqG+QmejjDPD+C3ycJ9/+FGockc+PqZOx873OgthaH2A+xMjzBcg+lj2ix
cB2hudociS8y65osIyGkNkhVsKAh46wXM8ZgL25aOIRYByDMpz8WpPqR2BmupVD/
D4v1UoqAhbIsRSaxV+QRPDJ/h77FIhaEGk9Ye2xlUoVLadvrvkn0RkhE0ib6c6Ck
m9l7QlWMpkArrPY2Kvc3apP7bMSUl541PX+CBOrfGniXBxnGDzEtbS4dlpPJQzLj
NFQ1LdBeRRQlkD1/FXCc4N+nb0Q3JZpsYRMzuA43Ky1F/i27plSSM8pe08QBinsI
QvoPPkacA4K3t+C++Cm6E5CyIzDOu7LFsJ+qD3TAPRgn5NQftFL11rFn0jMrn8xH
W9LtZ/CVI972LxUGc/Y3MkKjqapBj6hzwHNUr48Bn9h+CaWnuKvOMGjaow4wegvT
xxz8Fuha55v7QWGet1eksnz6HWJXDpvCeERQA7RYmmQgU3lNdl99E0bVE5zj4et8
Qu8YPS+iFZyS5eVpnYfZXG3jfF/Fa96MelOm0pe5MuzKFBoFKhq6M9YArsjkOwtl
3xr1w52Lgj3dBf+JIwWiJFBid2PsR5oVI+SlFdJevzJnWglb26UmW+qgDwgbkmb4
4ecQmOmbOR4jgdZUfYZOHuTNz3F7tKoILvIiG4Tj5XkfK1caiv6GdPejXkXmh4eU
pLGX6+9NXMU09fMGUfymars04GLhYRJIDiGt6fQvQRrJb5uGtBH6mLvhXJn4PILi
qLimgRJFPVSAq6MK7ah5Dw6zsSS9jI/DTTs+YrjF3ruYAN6qvUfOhR95Bun3+Xau
MLnxCbxZdEJ4AsPGMKYp3p4X61EwR41dOjU+5CtjrobKfe317FI/Iy+f2TA63e9z
UVCY7qiMttteYxq4sUy+5RYd/uN/ksuOwj0yOLnzFb+7AlHHXutyENM51lAdsGwJ
ORlUWkW/00vlTV1T+eIfcl2fWa8BHQIdQ76KrqB9gqQ8NwpIqH3CAJMq7VgAVm4X
mKooBm3bp5s5x5Jkzph5ITTGMEhL7wCFrfSyl0cGvwvCZ5vycO5AIuq4tXZ67tjy
vXgGTMFX0XPh13rIwWIQnA6LjDWle05NFHordW1MXrPK7tv5Q6NpeNlXlC8RuRX+
8FijDONn4gpPNx4k+RT/6nMISmsfS+aIwKYggSdSXlQsrj5sOqLf/U1heL+wDYdo
rNZMSRFcBWc/+h0exyD4zw8CZxf9z9IDuWtAu10T0X+vJ3xFatwZaC/RR79ePHn3
LLZPmT5k55mHnAH1AyJ59bmZ1M9EQH41BwaJA9QMRiSBPMxc13YXkcjSFWuptRE9
bRAU5urH/86YANypPMWb64+nY0Hb7dgIcskZQ69XPUtOuGccyLnALKsuim1Qy8tJ
LUjhGPoqNgKWdwzvUqIua8aLPAa+/j/gbtiESCFTWUFJ7+hTadK8A8UISIVoeLEK
hXjeaX7c5YlygLqH1LzhFddwsqSTVW7VBocNIaxShsHjj84Wot0czoIQOPTNTBiz
LNrLCHSYvjKmrPx5rN6XIMll2IKdXMbw/w8p1Gsr9gLxXKA6m8slSFusj9RcEUEO
IVR4jcSaoIiCOywmhxbB9Mn1d3w1nv1B8SA8DO0v/L7L3acCRKiMZ+bEQc5HC9zZ
uw93n+0rdAUf9P2MpQq4cVRJi7E4O3qX0I7AjB86yhM7gPKv9wbKzTtQSGcibuR5
f9yxNiYyPpFgdIJW7+wK9qt358hOkTvBjI5MP8jBqztD48/wWlolbfNcShr9sIVx
QFlToP07Tzag665+r/rSIZcoP6/G+k6uXNhGgQR0fGeP0Qidnh4AFusyoR1BGxnO
qx1HUidoTvC8fje0Cw0zRs4RreWH5zpOK9Bthr8D8q8PR6IfoQO8kvlsK8U0GF9V
WO5Er4vW95frYlgdjNEP4LwtG1bGZ7flKaAqICK8v1+Gq9s7G9DOhuK/2tuWCFg1
ZS9rqrrAPzha1si7P0hqDJXckXyPGp6tLtEt2TesxngycCUq5Tv7Q1YawSv6FhWX
wKxzNkb//etMInY5NB0jUDC7OnfmmF7xebQBdZL3mKQUO4zrgO8qYIGrYLiixCqs
s+2pIDuJObm3dZyvI2nnfULVsN858S7eONO/htA7S0z2Em1LSETPR64lzJ/qMqsk
VRXBXJPhfyT/8qFtzmfMFyg44lCF6G/2m51IwIPe5afb+Rm9m6XgdIWN4T6QvsL/
eiSHlKar+lo9iV1ZpqTP2BTYbOKDJxJFLtTkNT15JFG+E/zjo+vIV0m1+KvDfH7Q
cChIB2VAz7+wELclOwtO/1VW+hhzRFWiUsKLxczIYElgirnYo13ToeA9cnx3Fv68
EiJCgXPND1kLhPPo+rf/4pYGQm9WHtKEJ4ISI8h38gdHTEfiHfLyCQ0p0VrQScTa
ERlSbFNmpO/dxdEVKUTnMVsm38H26vDrHfxW2gIHVLy2kujMNEiaaZiEo8cr3imn
FL0R+8my1XpQ2AuD4CTXoBeqCoFjjJTy3qHKOfsooBReuz1gkUvu+Z+8xhW0uoh9
HRtM02/eG1qcuXW+bJuSSKA5m2c3f2nlUvQhoBABkkylueoNtkkEq7HG2YHz4fJB
pf5JpbP1ox7M48iNYuQ6vPOaMB6iuiaO4Ncy4DQ5Rv3gPG1LPotFuNM5hDLus1VV
Hxqb1eyHeNB+0y8vKjqP4T7g4HimzMkqVTzPjMROAapN38UdPolJxcotF3iZQvBq
mR7GxFipu/tKxLQMpU8DFAhTIVxSwYhQLqV+A5o4UTXm9oqIKgmzqdOm0mg7OUst
f4O0Lk50M6PF7K8vncVt7YS5qvr3C6Kh8XGebthh4Z//Cil2vg/Ms1opzwAo5Qla
A3M6kebNllvuMaC9+ZWAdIXBNh7aQJ2Qn+qVVFGf0n0mKJCaI1wps8D3oUUocEkK
sg1esOX3ca0GFYHZFgzMGhgMn/fyaMBzRUSdVfjR/ExZ6C+cnWsxzM4PVG6xBDoU
nUuMG1PGLbUnTx1tv6StOEPPpNBc9FZC6RgaYcrD1hxYNsR77bf6nZertxafpnwL
d8EBI86ceGFDCW5B8+sMfYVZeO3pG+F4QlmMZvUtBqnAnM0KAtChCtOF6CvfTPS6
SnQNhlI0l90lnN7RLnfSB6ePPxkuDnW/5OELBAIz16gW5Dovh2TB0KTlE4D/C8h+
BLWyWgm87Mk/Nn4kuxvwluDsisy6JQ3OgoHidgMy1EYmEFTCV6pxxLiWv5S2dShv
VBPw+SPYKJBnbdxyXruXbhTt4f6OsXdcnyyOTicUzg39yqr8bSbfIQpUj0GMap35
oCgK8BGrG3K8TFGpryEMF+v115A3qWKT5OzLn9PcKuv8bkUb1N8wo0c3y5HKfrHJ
+/etIbFJKoe5a6ZNdkB4/nWNtGpdPgEpZVKu78mUmiFXJFPsM3n+qLMHhp7pB936
noi7pq/vZWuKxeFRqGGn9tGjATrcoeE3lm2jztvcOiqc5yO3e6itQCfj05YYY8Bq
AichXNKbDLOc6q0o7BNxD38ihISaPd6Vu2h18TJHEbWWShowlt2Wfd+mTiui6D6G
F4QYTJ0Vt/Ha9HU1dHD/Ie9kSal16libhzI4MlJv16cpiOjy8ZVAByW1VxSpNpCo
p+JiNfS6ENODatJaaR2bExLmXQ6RNYzjisyjns+tp1NSa7Ib3C+hD8TqJO++3Uyi
QHUvix1GQwNH/ZpwVAQKGEP1Cp8T9nSjGT8Ovup3NQfkZl/ybNtuBKb8lCnO9+0w
YAIpq9SCAnbelGJ2d/sSmxZIqQZEFBPqRNlM3ETfbg/lfcbpzw0obEADnaMbuufl
hrcPOPtxBI+8vrBf+r7tgbNuPcmyleoytdC97GKt4NLytNsSUDn7OWm6hNpqWfTl
Yh1jpQee7e9zbBseGdYcO6acTRHcLujQIEAE8OBgAjC96HGUxashOREKx1sifVvN
S0oNlAyHYCPEgTlGiZcFnk//mwB/DmjdEdjvQS62OkkVlm3aIU8nwHqunI36Oy+Y
IWqqXKSLwXh1RPMzsh14qqLZVD26jNfqSBaj2HuPjnizDLrg++1pwPvzi7OO3htq
vQmy80MYExgS0G64iMy9D1+0LAy9psi9g3e2wM8yW4Og3leykYugAMoG1REC7Xxg
XKdPblmlBe9JbiyASu2sj5TjnU13EWd1qVLHd4z7qL9UNEmNy50cmOp26P1IBOsF
O6O0L33dj78txrI0D9eqOTduyytciXmXw2xxDFbc8WBOj9e/3/yaz/LFKbU/kiuu
UcwOZJBIQ/7d3+cVTnKlmi5UY0+JCDXaI4KRXqX4sDQJeId2bOpi1JZPFo0qTWcn
WZXXG4IgUjAJ/Z2ScDRlajp5fp7+Kk5drUhlwmmAQdEtkxhVNK8p5cLrDwdQaGZT
y00ZGqOFnzdhE1oOvM1iqaQz6v+IBNU5zKaHHHhhzKUwfHImp+krglefyQ81bsJh
hANkg8gzZNqwP+hin8o+qHH2F4hVOBLgLI+t71Jyk+x0Z3YzX834BvIqSIBpR2VK
tXPhV6l8oQow2DTWMC6dfB4FGA1camLY/FVMFX5IMhHMRkXMtpu43KCtBZDn3E3V
0OiCcRB5OTEOfgk9nxM9GKA5/iq2zBfk28Ua9R89ZxJSCDA55TlO9TKtd2ED7PYG
84+M3hpqndmuE79DSInAiiPqbnZQ8yMCUU4li5dvY3vRiFc0TqgmDEBWsd/9bEOf
bqlBlHrPkg+DKvPRys/zrymFVz5Fy+jcxm/w2u/fyfHQ1K2PR+dLy90iSmWx0g0I
viZcMjHuoNZHnzgpdgYBmd+UcicAaR1VdXFLFy5UJH2RJBhH744/OByISW6tlfzT
6DUapxOLG0bRugmGjL/j7HotByMLUfzdCVoKLyfuZB9Z+J0AAqtyOXqpnZmhec6a
v8l4HGWUSLMO5OtQu0mQD791GakLZW6o49sGABSdk6MJAdZosIXn7Rh/pF/YiXce
cKYCeNJGlgvp7xKSbvXgmwyf/iskuOmAXux+K4Cy/TYYEvCJQMMHbE9vgfpQCu88
8k6fM3LBZ3jvBqig3S9aYhINo/9BaiyRHNBGgZLINZtLJnKYObrNbID6uvaPMXTv
EuLs/cI9YjgVF/PU2V8s9in/vdEYFvoS1h0oB17vT6KpWvujuJxV0iGL4fZnEunE
cMDVzwJL5iZdTmsn/pJWM2g61TLGqXloppKaNy469c4VDWipFn+PjES2vHWCKdHX
PWq78AHIM8DaiwuS3j0+4z68M6Yd4SNg/iGtK2LcKEh3jopAAY/6+H115UECKTYe
FCZyXsQO61IbiNYxI82GevosAsdH+dPatOYm1yliWKfNEw5g/vyz1DRse5BVkUNm
WwJN65Cf/GxgPVTvI2Wccw/Vg8NXzs7LYx6IaphJHq1bnARZFAZCZgVWbBxBnMza
PIHkOe4nyWYjS+aCSW339xueeomf39xwhNdTt1W53VaLxMrQKCS7ynTuODzDv9zF
cKU37n6y9BSdg4j+efi113/48kIe83bXdE4uGUJBynpnCv0HcfjBdPTo5cb/z/50
OeF9W01DqSEdRe8lEkmV10KDiaSJprrja4T95agWOTeGiJHoRXnctDcavhW3t5WI
9YV6w6R8C9WUFyw3WAunwVvWY7QkqOj9zmMDxFL8FD5onLUT4/03U8KPgekR4hSr
Il01Q3N6EQLDmoL/CNvnECZ81s9Jju/VeB5gkWhbZdR57nVe2bxYeNm+EupXw4A9
ux1F1yo10m/LzUpVAgVsDXRZ3ndLvGV3VMUUcApUSGeC60RSkcsuCMm9xG2UUsuk
Slx+rL3eMrgbde1zaGMoukKMD41xtBMJSe/DeKVkYRHLCRbhhwASnEW/kIAUHAyo
53YTLs+bgBO+KnDqkKxdl0kpm0bF1vb0h88kztR8nVRN+IQqKyTfEyJEm+Qfv5iY
HpmtUlzfCYAgjbgu2dlDOg+kj8EnPWqvzuhlPtQSdsqwsagagB6GEiXUDyZImKJa
D81W5ha6Nl7clDDKSQKR4jyQ+L7zE+CFIJkvAvNsEGdETRn/ENyJITf5LzuNLekh
QtlDOJeAg1G+Ydf2eJemSa/2BajS+R7Uno0uDfRe/0S6ganqTKGBpuge5q2tHVY6
OD0QEJUQcsgA3nltMEYCXehjcsUzzeBSdMMcc68dZtq5dMRjOUI361wd4k0BweMV
h12oK75iurwcZoamQd09WtlBipY27K0WqcQsTldVJ6aE5pVe3mV+FgxvhHFsGVpu
zlOyaH4YwHv8YckIavIoWHXt85wVejDjJqtwBxX62SIJkkmIpZyPkovN09EBpdZj
XL8BDcgP97jwDnz+M32ubgj1/ixC+ydUVEmg4vcPv9PkOR/Ndcvaq6HpLZ7Pphb3
3KQ3eziA1T1Ct/X1wcuxcnu+q/N3nyuGlLkOUfitt+kZlA9Eb421hJsd+pEUXe8h
uyTmTUEaylcd/We8nwH62GVm8LqKPiJlirG+hGVMnzuN9m+t1fVn0cS79Belfw80
rO1LMmvOJDPEa27mTeytAatlYvUOqF7XJMotA+SHay49dJ1F4g5Pnb9hghZjz87z
9weLgBS6X5abDqBOPB+jsRWBxlZ/Nvtzuf6E1zbk61V9jMtxRV26tkMXMyPVGtod
a1xj5TiwvewiVhJAAEwsH3IT2Ykp6i4Eer5raug3XH464d9o5orDgEk9jHLrBUTF
PjQyqoycRMgnR2Yvuab4AOVwbVxmh/UrsrxrguUnZwCPwmWoaPT9LyBq9pZK0AIX
Z4CLD74Iknf1EDH8wvmyOfI6EYmX6Lur7OO2Zf46FzCZI5a/+kFjXYVeZxBBsit0
YKMcR9avga0hdrZD7arm89kgV6JuBS6MBRCqPAMSLQ8JpORyY0hbbmIjX3V1Ktv6
VbmTwl2ML5/GPzLtk3tg8WVi7H5Le+pfrDAJo6iaSmcMlvir5b6Vq3IAcRbW0qPM
HWvH/J8K8GdSjUTYLD1sBMc1bDxN+Cu2YsCMxc5SVznuSjFV89U/JS3a+m+ikOhC
EOusgJR8Q/yMPoE8gthDD3SyUGbM6/xpt0GIYlDqQ93pWxkKvFPzj4GPW3UYGJ3q
v/Y9Z/+ylk6VGrQtb32nVd5lr2SI6GNUjOLLX4pNUMHZ4jkL0DH1ClvXq3E80pTM
wJXmI+7wfLIQqLp2FDKt4di2ca+IxfF0RcouyiWzwF+wdSoYkSDg5s0YhodUlCZo
EqbYRuOOc1TmImLM9nzFf7UJhx5xzJ9bajgT+dM1VHyaqsLt1cDMxYvUVm4AUCAP
2iZe7OipueOpqQN++EZf95WPoaWVGLltJhKjwEIoDttti8lGxzhULtIuYsn3HWTc
FbiluNdIW0InaLsDm+7sU96GXiuZ/uR2DjTnjA3esZ/X0RK9f/daUK0tW1qayRin
ZH59huALC5uDjFN7URvhZSkCuzARt9/Gu5mXYZSyyDRIgpW/rTb6zOP/bWKI1Ovj
zdSqVQYA+gV/SKRjnYkwumI7IjtuJ8kogBpyv9Zn1KexHAGIvPfuFic51b5QkN5D
D2e70hC6AcPK+4NbcI9j3eWdGEuovoIQ4uXm4qAfxMJSXD4qWRzm4RKMoQ4oPlrZ
wuZGDGj0bW6L3d6wRGzEbblv/6eEZl/gNSlh51hcTD5lxtdlK3QPgreLRAecxqC/
BOgK6Q7D0TyiC/w0TumkBZxd0jhKD6Rb2Szzvuo+/SF5hqVQnVM5gwaMkHnPIPHM
MqQN4yj+8xDQzuBXaAzg4C1Cxr3vCril3p+57zBawaPAa8xh+0loJ1DTI/k1HUg5
lNYA5iFHfGy+8BjPIqMPl19Ul5bKRsVkKgeC4U8SnUPDfBEtgl4MH+1uIWGYsot1
6sM1r4MaWRJZqvPPx2RFY3iS2g0Hl1+bxBAwzG62E7tCQ+vVpkyw8LZ0Q1WfxZzX
P0bMrKBpgObmJPVCsTEpaHT8FTDCunGwjEwUz2SuQzLJGXrakFMMW5gKrWPuQLlk
f3RwkcA6K6uQXJuRqjcfdRKiF78tTaiD1eQDWfwYXd/O3Bx9/CUt1qk9aofqWDKy
zbwK5mPwHAHNNFJk5onBLsxGbcE53HWQ5ciZOZz8tovljeiWxLrDPCt8B4bL0RID
bN6hs8zfMNIIAzmb6S3bwn2DlJDjvrs+sSl0N0ONxgmpVefW4+umNwIIMg1YHbsj
33FiXNTzXWk02cAFJ3u3XurSCTHNzz5jMFcQxt4JLvdiroBSJLxoh7afoBLD6ArT
BdVhv9K8qA1fZwNIykHLS0DISuOg8vS+kgW/tt4Q0M1jrq5ZsgTl3utmv5qodcuA
BZ1daF/fmshEQpD7rCOatdb5WGdp+yZOuldxHFC7jli5qzAyTv1AO4UstvrXBs16
2YQaYMSIrw1TpNPaVCDif0mWY2Xew09NM9zoK/0Qudz5FZOtXoA+6gXXxngkJZPR
ms0dKMRGWYLqX5cz6TLlDg3ER16BccEKGuaQUhpSYgeS2hWW5xmXj8KKQnc/47rg
AgudWvzQRld3aqCWpPO5IZ7RRHZ2eAzptRtA3pgidq7WbQcjxCRuZeGtR3RUfcFE
OHEHdV3a+JJpFapOlq7uYidV9aD+7ItPqeBR2qyHCeZeomQKWZBrc3ELr7G6Byq0
EzJBnfJKSwQPO3BpduxF4N7BFp00/jqc1AF60UFEMbkUOUCyWtsORa3fUC94MN2W
LEDbARUXDsE+UyC9NECdYjN85W+PPEqNrPaBuwo7vJ8/hs8+kFy9+TYMPlkkoZo3
Y/poqQBYVctOtFD6T6jCjOHuKi1B2SC1QJBRQ6Pwt9dJlx/MzsRTu2ziHDbbqZHt
bkUn6moVoi/zuJC3ZbylMue4RmtUkMEZdtuA1z+giZshc09LxvK7hrYOETjEdWz6
eijoBy6qOSDaUiqf6m2N5Q==
`pragma protect end_protected
