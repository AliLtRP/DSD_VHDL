// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:47 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
GqDU+V0YFatSp+kMYWOHBZNrvFQEatphg9PwCSVX+GtAxKGOl4O/eXOdpoEkyOOV
At6Z4xVVaH4haYlmI5e98vQRT9E4b6EaFUJTzx/DpMsgiwm6aiyUmCLamc+9DFbD
MBDSD6LMO8ZWxcTq+MD/hr3Zhuz4wACZiaKLhCZibm4=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 22368)
8kLX0yqtAsLIUfy+fSWtSfGqt9Y9jn0OPyUQFhmzX5ZfK7ilsl2XYRtR8p/gy+wh
2I8855Bo0ID8HSnBgzuTKhlZEHQsrOe7NGkV8QuEuMCpkXVvTi0JpltrHESCYdlb
eeWmmAHENOwzCkxz9G5Ccf9bh13cUycYXr+dVcB9GKKX91P0SA7885BKlE2ohR1E
m1NPvW43GL7rKafHOTnwJBgrfFU+nz6S+tBbYn4CZ4RV7KdWKph2fAbd+L3eBv4F
RJPRfSPGcM87t9Rl03yBEJUVUlaSCB+92E/l1OhLz7Dzj5evljB0o6z6jCInPkag
Pb4NQrZjXTaSsd6kB5MxYwVRmS7+bZXcOgko5k7/QMPE/XTj8OrSGMWD1TrzdTuY
Ysu2JC5S40iSIOPlzordHSGPIlx1jVKoHxRWD8d6u2cFxatOhMn/Ir0rGA7GysiA
mGapcoTqvvZVPGbsATILMTdvqx55JGjcWS/T4yO1o3425IVqUuQscoUQi8vcogz9
CHcfGMHw45yisBCjYg94H8vkkpMr9y4HBfcxAZhRj29aCC3eGJ7zlzOtWdGkecT2
pZ96ZvDLhRhgAKgHTBkv15ew1j821vX3/VzDAlShL+XnoXKcFzY0DZqvWuOykxIg
8F+/vH7SWhEGZ8PpBVEQgMoPgwW2krg71v6oTkfnk5zFjZYdwHSKo8wtfOMZ8nyS
fKB1l+SzykTOLMx5PF4vNmLN31DlsoYcoYYTycXmiw1X5VUbdRJYqdtxUjhjdnjB
TU/nXYONWUCuhlsjR4YowwfooxHFQUvtPiMA8Ldl3A1FWLnI3b6mRzPkRSOJvHVz
Dt9Ay1RRch+n1E9PcHX5yADSbMWBLWCrvYkmxbc08O4Hm82eTE/J63pmEqV8pIdB
iMmWKvQCPLqvRkFizRd0Nd6UgDk2WpdhXl+H5oHcpsJscdm9d8+DUfnCXwqZv9YH
y9SSC0JPda/jKWonIovxJftf8Lnna5bEypRK5K9NJQkAdrfBJ/eagTwvzJqFol6G
oWCm4EK6P0C3l0mQ8lgDNrH+fdPS8qH8w1DYPzvXgPAGSAOxN61Gy/vMywoSiFqO
ZnY/Og4g5kK4CsKsM31hJtJrY/O8U5TdTmSWRAw4+O8NZUHhDvwevMd4cXLUGOTB
PWGlEWj7oKaf2fkjcGaRdkYTOn/tQBlJadCjwFcku/PRF/y1MMCtfgWQ0Buk1Upw
nLm8zokQrZ/Ca/IhkU18oKO3qdu+LrFpb9su9KPJ84fd4dVQR9fxOdsYxQUXjX3X
HqAVV2Odf15OFip5/AE8xWY8xfMBv1DuA/GQ7N6Jbv4iCizxDsJNJL6C9nnAixWN
LhuxcSrXUIzdg+kfQzPm6k3UgjAA1OteR3XPlUyyaBDGtdFrXYEjkk1UO1Mc8zTN
BCiirlAf7RmCiQSvqJDNI48K0l8/7At8HTrDCdrcFhnfyvAmvm1RfISm5NzeEG9V
dXTP+wWBUowKEE4zvDKBhYfIWiKoR+7pRx7nSuYwkOwGB1sNMCGxcaXkjkJQcSXF
gf3GNxvFTBA4vZq7F022fJ2pgxmV2Y4erYaqCZ7MwQE2v54+E8GFAPxdxiYwUzkX
w1kW8gNipXmulqxlqzcw2q/EEsj5U4/tQEKxtL5G0lLA3T1x5c14xvpM4tEb4/Rh
cJzq0lqXFGtPULQcATN/mYppjBxQ5dmj4WKm+9WaOSqgxkH0XMJh9qQBTn0OzOvG
4bECLXgmhQA833VUf8HLGCkwBiwvF+s+N2keYbdGwULwGNUKAPAHQp6JttLJxJlB
cWbBlLZDj0/uauq3e9KZnkZeC0Qlqjz+6h10oX92kCWJvfzNyLith2tcNPWUD8Gn
ot1VpWMU6RTg15CmNCn3BQgqEqEBvjWNFHFMcU3VagZLSuwhBcT6H15Mp/Qiicfs
nIpo50LaiVetrEK4lI/sYjH4RKYYE+T/3tj5M02ohERVCJwo+0CmlpL7Eeh2n7Uv
iHSL7Xg3tqAEktO+rKq4bb9kibl/mEeN+h+k2ItWKY+CzfXTcltoQdYYxETWimoM
e45Z6dBjHHAn7HwvgB5vh5gd0wOfInEPa4laqDRjd8f9f3SyosrR9FTTTYIGyIce
whqwifvp1MHe01nAZRUZ1Cf+cUAVNdzczcSfwRbABhW5yUK9yEplJ/NRE3rF5tmA
s2Au9UjZm0qyjPeUJ36zD2NKTO8/cj5PCaElI1NagFMqeosurDigFbu3d7+dxlJz
Q3cw3ZajbWpu0s9LDrqY5NpgzI8xFllSWbI7emnz/gQcWu3cr7MvRwP9dhW7vxVd
8fYnYFn0I4vTtcwVehgxKH45VglH7boVYoHAHKnFZL2Jt0+YxC/oMjFkGNB9/bAr
e0aFgjXVbuaISl6JI4L+0/eloxVaK8YJecJ+aBLpqctgNdXbUF5r9H3KNsAgp2Il
3G7xWmRj7akXPvH7jS+ZaNFJ1f4N72Kp3JesxuMKZYxce5e2M+r20drsb3C6jyfa
AZ/De8yV4V4ZA2otoHekTgMvpBVd0dXi5boxBFWz8/Ka8KDbvB+SOpEOj8rQWqoH
Fa+BRGvPB+SvdOD5STOLgtlxRpExq76Ix9pqq0vKfl5d1Ri0IGxoauw5Md/FkRhi
u9HhcutaCO4UgVKkLhE03GTOkL7Q8b+Dw86ri9kzhkNKewVt9SAjfetkSMylWdTa
yKFNjUb24ShkEIsBHKyBqM1AbMYM3w4egJsDPcFKH208VVrVqgDuBu/+xgegE8Y/
TiACZIIScJMOZQwhFYjrepV5927RwrHCkZMDFaKehgufptBKsSAdz1sCwg25qcXy
o7bFySeKp+5A77rUqw+CzxjC9f0HMblipMbmDX7mG4VKbVDFsk5oSty8y8IqOYC+
CVnI8+YU0I8xca7U69QIlUDfa0f7nLqdId/5od8jHfXZPy7lqKtqetFEldUUDz/W
UExTgGAAGTtKXEuAMYyTYBNfIAYHM5slV0otO6I+YuVlLGkJaDMdNVfVpQX7dK+7
hG46vJH4YGR37JX7GM29n+alp2kZoulJEaKFffsiWoE/87TNh80BijsU6Ti7/fY6
s/okqOijTR2ycLtA0gUPTAC6XY4laWdr9+wd6nXjJ2i4N149VmAb3Yz8rdLIjKw9
e7KDSomgc6dlnNtnFOE6hvq6DVfSCPiySY8FOYmISX2xhfONSb3edxUBzbLU7WTI
CrbwqkrJq7THmdHvj5/T78aKa33C2yG5VyUuoyEeOgo2TAOMXc0CVP5gn4xhJgRP
bMLllK9kNHZV/3LoTvmWiZWUtwecFwcN9cD0JaGxCDK8x6TbDiJTYM66O28XDYAA
XYEjy5GhqM7wTSVOVBAiPqbX2bUMpZ/eWVN1P+VoEy6+1OTLbiZiqzg68Qp4yvct
ivteRlampoTupHckO4sitAhFQbk6KH4D1rjRwLA5tR4qDK5mmKAk7XS94GXj6OHZ
PI94e3ATChg5ZyspB3YvpHyn9qg3vgL25Tvuk638JbEanmmYyC7yNrCakLsovHjX
Nqk0kXKxApYQVq0T/XCDfy3I2e2U76BlNLsAmTIk1fQ8IiU4HGzGiGSCniOdzxwe
TwCs99MougJT/Ap0qpqtBMPefeZwgHKCpAI8WvylZJUwfLFo8vdTCVclZ31fDVF4
tvanktA7IOSpp2RoUYa5zVqQe04no5EksoZt3cJyMbqZ8WLYLW1ER8RaLSDu6SfT
d9KZVmVtqE+EOc8BD8BQPDgYwfFApxb2NLBOeI/UP/pbKLpyk4JPK5aOd4VmUqWW
93JqZgrks7kJh79DQmUkfbTXEL57ibTrEnCt1C75y3alz9UkMSvhi+FDPfZx2R0B
pPgzGzzgx4rnSN3leSvSWMXF/Jg9LiRPKwNh4j5E+UIc8dX+BiidNu3KErgZ053p
VBXg6xGEDBohlE6C/EoNyAl8v/yWobRV81Av022fdS08B08K3u/kk77r/iMP/E0z
pdbMkXUa4YQBK3adohVM77GhMBJ2awofyWnYo3zMhFW5UYQBT7Lk8JtE5+e5nJ2b
nOxAZUYTBN380NfaZ/7Hh3qi3Ivs0vf7gfKkYaA43cU584Y7eHot7hK1jJquAjgy
Qxh2pi0sshBkX90AVFo/G5cGKLw2gQe+sOMM8B4EcMzDG0dmcpdgDIhmI2ONrTMj
iKPfVoRdW80ZKWmOSiwOk0ijCrLwtiDY+9ty46rOqvGwou7E0OJpKMAZD50AcDcu
urvQCpJcjGKK2AnsLpfBBXubG0vm5bWlhgu4LNIkpCO244k/dS1qEUThGsUkuvWn
UGSjdWqXUPQo9W4fFqAQC3fBlXnil4XzoX1i5XBm8ZeaL7RLRxekHilHuaNDyxOs
aM4h3hevA4LfqW6udy6+G8KmmLbmH0U7MI8urHfcgKNB6VrDv1M93LufRrLtO5uN
RBDuzRERIV/ZQUaD+yggOzXwq+0rnLcB1yD5dlfjGysqRY4tio8oOygMKaak3DqM
9XbXtoyrXWwI+V5kv327Ul0dUKh0Cav4d2wVy3d5Q/mG1VRg9bUTzy1253ssu7+j
6Y6Jd8fBY7dU28c+E+l/1T6yZdeeSpBV30WyMNnML+hmrMs9gnA4dQEW72G14/HH
mUxC7cB4dL1uNZ+2t/QltRJKeTrg0p0q6zGseXfm5JxOx+OMZjCKBpy0K2pHvqSp
FA1LpBOapFE6GtHp80VFXRzhZ8axWig3WU+oGBalrWY0PRN7+qBR+5r0IRj9ouuy
GDCUWq54SNPDGZ0ZHF16tsxuVwmlPyE/tZ84JINK3Uo036Oo2MQwNmzVI0v16pgi
x0Ne7znbryse+cAdvlclPpoascYC2uGAg3Jbamg8yZ65C+DDMnGC5oya6y1wVmyU
eXTR1fcgsjT3KruZKDl3ofevxNBuF9myMvphWCrwcQh6Xw1axy2NR4GgTvmQh+iB
TprlyVO4AAat/5mSJuQgvlm3CJhuyJ0VZyY78cnyc6acMH29IaIxVhyMaXbqh4hK
YBHqnEt86PAsH/W9MzUGKYmx5k22rQl9FLKfwIZ0LaEwOKe8hJ9FCiL6IitTmdgb
a1lRFPLzC/L3QOeSjc5HC8FrShdrs1nb8mXc/+Ma0VeHfrBayECcrsae+H7EeTwa
8KZODCA4LYjL54VZWXDdVIxYr05gSmvCGl8X/GNFE0DJMX+i1TziSv5zJF+6tW0a
P9fSKN3u3TXx5+MNBXqj4dsEdS6lebaiW2pGAPDr8Bih+pJ0DAZmdn5YxQtwtVS4
JJw9v4CEEOoTO51stGvXYZnGGBpuV2U809Yt5CzApsEaQm0DYQrKFq6vhyuETiT3
IGYLczkm2d4pCY+wrNcuSJoBS8ZR9ui2YejAvacAAp+Pqnn5BBSrEo2+7+vA86Ve
tzNFjdolFeX+wjlCn9UyU53bCEK9v0l/VQpmQDoD2otpLSiSNB2NmKGwsji1BjRB
wc3MaDQbmaO8DOPvG+9FuVHoPsL3/cfqpfU+49rZ9DVT4NeWYJFOsEehkgk7wm2j
cauQGoKPUDKHY/vX6W8iAUQytbYihtNcL5yhkeGMTUeTsZNh2JiS0xW0zx9jd7jG
Z++6qFK25eGJiYZAEVgX2tLvAivf3ldM0X7JjqegUDPMIt/K2k/UVgxF3iocHQNe
7jSzVAbOMN+bVRv1INpq8dyP7NOqwqW0O4SLu4rrYNCNCmiyCE5LioGmAlR03cLC
HVAS1HSSzxe4nhrT1u6FIPN3up8sBBVLF8fXuCxHuTKYSxRseAeB9z4qHueS5TVH
jYzkydqZHhSx+hfBP+XhPKt0ULo8UwN4XhGusZulnjdvx3vSCMjNWHPV6o+I8goA
cFaBkeN6YT9RdVQkvcSaRGFFUqISqq+04tfZlBOccZeb4lv/DDeyncJA5+1Io0xD
+ZR0tp8WDIsg/t0rnMT6Coc5douy4HvMQLUsnVSgXixECigVviv1u80W9zIz6Qkv
K4HdgNyzmKq6MnfBTQ5vVkgBN20ciULbWn5agrjdDNCWFEyBCJ01uX3qE+u6Zm1g
TqYYaz5BRqhP0Ab4YNNVyMGmYCwQcudS31Wb/ZwdzgSi3pKQ19U/m2YBixNY6MHJ
CXwmkDKdzjOnzwAImB5PxDZuZvCnMDr2ujenHkVvg4vEyYK7KVQ881Lu2sopCEdP
FltPQofKTdh7IXC92+ZP8/LEkzEQqdTlaKirAVeu9/qtSh/MkTLhDoJCMRFSsfoa
RRnRtly44u/IwSOTonNdpB9jMWKyYOZQEzmI/e6wLGuUzrfFGpWVYiZpmYZsw5ac
1HQNGRc1Gs7Ed9R/zRa9gdnl21K4s5L134b1AzLr9zqBLXC6NGKjiTFNOJ5odaKT
LMcA64kSIqKVzIptai1Pfw0zZW52A3o9FOYmuQfLm02Imte8U/Gx5LJj1Hz9l6uI
0mqWQCDgLNl/KIxOM4Ch/Uip3AwhMCfdc+4+IDdBlW2b2rjxIbwgiQVkIcsexN0S
gX0u+s+gBywX52u4eiE/SljuTs4Yx7bk/UPh8yQ2Daqlo9TDOZFBSgKDCOWiFG+d
QUYCLqxC3CXN6DCEhLlVmuDRYeyczGOScXeaeaYmX7TWllhQdwGsshAOHnKFZgez
ZsdL8gCgP3o3l4J/TDh3hgSEUIbr3anoDSlBzgIdJ2BN1iNEn0uumnwHc3ThnIt0
NbJJZpMUiMVmXBys4+sio3rozaCcEY/W0W0VcUBww8io+J7bb8FC2f64PXEkLGHq
OfYkRrgW311eteyjhd/bP2kU23hqJWapzSZ3xk2sJNsPdbQHwz1os+nJMOx9Ixd8
XUKzRS0e/UQ/WtEFW+A8Hap+mJywLZwA2UR6v06aBHMfncZBhbSBbXsr1CDftCF4
UHFLGQkZyBhPrny/L63TXnU/Em0yG++tjlm9gIJRjVyoWum0L/EJmEKE8oo2tcPa
0yTws28Vd3wi+LnH6PSjpYv0eIAU6DXpCSN5ZowPrEoF4SqsSL/s/qFkSL8JOnMU
Qsi/U3AMSemHojDmQLcMh44NfwLHep7L/qFPcvrclDPAum1OarmZEKznPKybZSCy
o9L/yjHxwafP7IOBKJ042rVn192N2wvZLCKFsyPsZF8IpwGDLlbadgHsoG43cZOi
pGYYB58zpNWGxfjhGZgQCO+x6CrZwGtq406QtlYsbcIa26e2tV7gPOHjSnjdMDiC
p0m0/XeZwQoz/lvH3rW7T34mpiiR+2RjKNMHNi06fiGBam96wphdtMv57DclPpVv
S3XBXNemnFXQS+2fyg1hht92pyxzSThrW5lXQX2ztKcUqV63HrI2tPCI6ImEhU5i
UD9Sb2trF6hN9D0/HWI8ooFZ8Y5i2uemcF3KoLVznyP9qMQqNLI4etddyNGgJQOG
gCjsinHdHjmI0BE/SPdRsSWvNd/wpmxVW8ELcBM1PimLK2UzKqF0sCKNk8p3WkPA
ZNSTYgp2rU46mG7evxr1CkMZR/lbHR8zUQL637uNNDripyI/t3tG8qXYfazUVQKL
Hiz5XyqnZso54Qmy+E6xGV/ys/q8v62PBPCUnpjb61DLXxs8p1SyciLaeDmSz8jk
etuTYn5UKRQ58YOOsPk+t8/qjbVJOv5iPY8nbv06nH3pb2TRSfoFN3klq/obU/rw
bSQFhGYds2znyVGhweIJQ2I/7He9pQUt4qXxdNhbpc11f5FMKdxCs6YcoHlG9pkK
wWgd0J5S+T35sbJKMKpuLlayG6b2J/xM82Hee0eBCiEyES8n5VbgjYZsL5wo+qlj
tflVFT4k5qMHaqSqNrCBd01CzTqNLjeeHNbdNi2Yzrt+DRN+VKTt92xk9eprX/OH
fFsixL0ddds0TFOpFP3zulMhJ/Sn9r2r0XgWoEp8UGzirZ6bYpZ0+JB+A4jehzsi
56obolyHmu+453QhvEH94vEX6BogEIKNa9SCArlqEKF77NPsomVR77pzFLUyIF3J
EWVAxuiJoU2ONYwCrBEJ7JwOyZ+4U3KQu1diHafLplrarKgHl71UVGRGpN1LMzTM
oTCTfDJkrnChM/24a7YE6QZnNVCKoCkFMrl0FKWyAjgasBiRdVMX9+6a1/WAUAIY
2lWxU/WrPHcxTYTnXFwzCJgn1v2nXljhp6hReQjjtzboAM0QpVDmdF90MNs0J/6S
pDYrqR4Nz8cbmaHLME4CZ1yvgXYHDLaglyr9fExyUl8mnxKdHwmBrZB/qv30oSiP
lfgO2cUZEdakqTwZ05wx17+SMVZE3cP+wRBz7ku3ppGuMaUNDWv3fzRR8C5ISzOS
mub98Y7dWlWgUpiiD3G4yQpp2GDmj002c75xrFSOu8+CJDz+sjgerrBuQ6wlT3CP
ClOKpDvoso8jK2wJ0gyLxfIB0A1cfwBD3tRLpUVef9uTkRXcp2R8rsUW+xEZzodX
GC/YOgh9OGF15RiaXC9ZpGiEW7ir/5C94VTClpfCOZCdp2OgtEZsUj8WiNgOn0rU
wN+iCo19OU0UU83L17NCc1DRhd4Kf2JcIuASL5QRkpSlLgQkR8RXFbUrT/SasX+L
v/no4HjwJcHt5s+EFbIC7H6717lVH5LImI3f8kzFJUv4i8hHrAR6QnO3A5rDYzjn
75In2bEZ3+BjHUIoCCVqFWSyHTjmGfAaNY957ysduSdIwaUuPB3iXplW7kng5vM/
tlyT2U2huZGEY1KCvstRX7Yys1QjxSAochF3MBF8Hph62QM1BM0/hoFzaqnsYd9g
t/LbL2mViyUaPftIEhON/g66CAXIMbwHWdRfZVg8Vtr/ZUAcXvp90BnlGpijtOHz
XUvTU/tRDrevfC6NSFYzitz0oM4Ofpatb4ZhPUX+r/M8oYwt3mncuiltEZ223Jv2
+aQmY8jP/o2xA4/SDPk7nMw8uOYs+XradTvQ2OBXgi7neRX14l69RFg4SRgxvD6v
dV/BvHXffdD/iT/lD5mYruG6UakOARktYiXIOx05XWdTQPcWgZehTeLGgKDi091E
rJp9OM21ozqvI2Vxp9c/qxVkCQVBCZp/j2L0AX5wmX5aS3nMR74Sh8gSr51A1u1k
yrv0DEAN08vAs6vhn8b62l5vYyvJqp0XLOGK7En/U8aAJPzKumO5o9bPnnsM+xPA
VsDgOO0ZOXCFM0FDVDwHsU89iFMkna62QZPaIZgzZezQ16wMA8bM9ZAMi9YTzjdc
MZVPNdQHOJ5SrP6gtkktoG8Bk18ZVB7x3BBN7gPIxc1/5E+2ik3lp1u16pRDd+T3
U8zHYtBiA8KFI66h+YPncZKLL/Ys6eJyIvis4oZeOi8s9o6jePJ2RU0IxF7zt0Yz
BrEjLJlb4WaXux79jCOPwOTXKteVmmXBC7lCr7cbzm2NbgVmF0JdzdfuoYFJuCs3
H/pTdP/VqjlyocaI+WlLgb//ubtWE4s9PLEDZz2KYaOoSgbzpoRCFuwNbZb5f0BO
8nLOSbI4PUVDw4Ua3G/6NnOcOH3Fw1W17OKkrFWdye/U73qDYbKGoiy04GiswLAo
wV5YDmO4Jz3ep4YSpwocmnWxy/r1DtpmfYka71cAqAEFhLso+X1Ena8MTVeUNIw1
F2/cae5Oll4NFzJDCbMC24U+EAnwuKANXiCbSuwtjB+BQAlYXKLgv8pbw5Xh5KP5
sWKMpvYJD9KGT0o8z4az5K2rNRep+6Wv4dBl7P8SVTNTZnlK0n+hzWWgeXKeMzOh
aTvpXJAhxl2iJ7eXWXyUJHEjA1mexk/wRgUuRpPPsl10lOpMPlDYcvZuZlSMnn9u
4xsKmilJqpS9lVGJGvZ5OW7jp8i33LarhMWFRC20V+3HoRjKBAGDV8ioSt24JBLC
xL9QavU9COAJZygPACSwjAWKdqYvu/XaVhgMberqr03Cdr+vbIQZG/pyMX1TYIOy
hiinl5XGPp72jDbVvmdYGJFMkRqPt8LPIfzR/9h+G2AKaefLtofotQL1MrCGYLPs
ioeW8KqTpKWHPMINEXiKGg/o/s5cO/BOuBnG/XSIE8FYNzD9ptAi1asRiUFRcNqK
hd/b7ZPSL9wrqGeApnPxAgET0oJd3laJgtv3jtgBms390dArLVrJPl196xI7Wn3S
N1hiydg+hHBYh4C7+1or7CeWTE4XREgLjyU3NsWoJ9WYumXOhiZ9MenHbAsxOgvl
AQuDVySQ73Jk3e/5uX4voaMGKoBW2js1KuWG1o63VnQtUBogDLFK9qlN4Xp1EdyY
Rbmz/Ap1gRKMRRg8zf7nN1k7hqQjnbxTBrkjLWdr8sE6sEqpBk/KY4YMFGqcqRC1
JIz4USVYvXUOT2XiFX2+/tWiVo/JVmt8ENDf5iaqOiEhm3go5IMI8OzsfChjmYVv
T131f5ot/03oEMu2k9NJXcNPYIswt/E7V58reQlbwIMAYeBQLuh8jHVzVeD3Up6H
faf4dSL2oNEUNHJ8PYRYeFgRQ08Zx7+QgWW5yPgZ1x7TSNMQDjGJ7QTm7xB2sHwX
7JVkPOpx8AmVQCUbf74ZsdidyCv/IwW+d42yZh6Q9Cvalv/q2V37B3Y4AD4pFYqw
Oto+oF3bl8uWPMre651IusMgAXzaybIbVkJKDu7VIndndC/WF2oOQwYGpoCd0ZCN
qwrmsFV9pUbuD5fSeMiOc6lBDcToEZYNatNzyoO5eX7VHCDqfjWNCEdMpmVQFJi8
Sxyfr2z8kPDtvAiGQ2HPuR4FENYcA+fT9VvfciLxsuQ1KBxmVeiKSuRATyvMuhOu
aK/2ShXkQDJmzWs6b/tu+uGHIFehDfZsne+9CSf5xdnYW8JgcuqMr2QeePpqtx+7
t09s+fpT7oo+Ymjo+goSoHp29EHjkmlEWy+UAHOwf7Sd6cwMxCKnFp2awxXlqG8+
yzuq5qmB/OnJqp6WGeGoCMnReT3SaomBLyXmStgRZaCDCjVTfd6FyiqGKR5uaS7r
YBE17WLFowstklgZ5FWtuskrUuEDWfDxMyIGi1GD6+bdaGf5eg6JppnKCh3EWdWA
RLArEMvCrT4EDTk1aj1zBbYkYG5shdp4kh0rdLFZ9d8QxgeQDnGh4cawGa1VTBUh
e8DCTyT3fiWeq4EQK6GYIHzKA47q4btOQgHEuDvCKqy/bgFdwEsOJbkXTEevgMr6
H4v5K2ozp/Gi0pFOKpoDr4syzPiN8lFQzgMNLJ1SigOh69Pr0vSe04O+iXu8atX9
/xIsCLVkNZSwtQjOZnjvgZ8R71KZsHWcCa0dZBPkHfuYXNFdbgaLNHnLF6EGAWNp
nTf+1WpKlYoSHGkW9MQ7i2LU/yxxjTO+asaXwByEV+A398bWgBgq/bHtEXDAi+BM
u1ABNU3leEcmqkmjBn9AZFZiTR4bclN/qDgSZwThHaVKxw8D2mIv85bZBxs53tRN
/bKLj/a0pWYou+RJAeuAM1BUn36/TQjym2xxeG3ZC2DIAFKFQV7mT46eJsSf5xaE
SnPo1xAamqSLrtx83rvnl6pkE9/LkSYvElDT07RXdZE6E0l+c5Q36am3Dqv1L6s1
1/o9asmE7cXa3ydK6Rp9aHYDmXOj2y/lp8B8BG2owWqqA377ZvXcHpwl5+/VqRqW
bhvBMV26ilfjPEIfGQAsArxk2N6z0JJ4/rkFg/+C3tRb3QFqjiyJbvcbCZWChtjB
W4VBx384befAWQRHcd+gE/894TuRZAicNiAKuDmO7qZO8y6Fquh8a52EEzwuZ8Pb
sT0I9XcDyPCYF+YA2bqrkrJWgy9ZGiLUhakC3QOhVG8qVTxrpLG4wJ+LT5sxRC8N
n0nyBrrw/vLvUEJBwCw11tyRVVvvcsTqsKEe1dLqKHqPNf7ogEIUwKxiBL0zDybe
2dM7OQftZgVTas0Ok6fPrBtm/qasahA3x+7FnYWd/R32HvxLAE5x8D76VRPqrVeZ
HzLjmaozB4ahcAYYN0CM/5vA/g3cuX2FAtqcYoTbCqUIN8rzLJIWHbupBlhYf5jk
MnZVUSEhmwr/MiFc7aFqYPZ9wmTHqvFd6u2b25czEmLncmtNT5O82NrA0X2k3wUc
wll+SP6HADHq2EG73BKnro5eGsczAhWPn/LRBLY2BdSqzk8TH4Z3AlHnYIokPUTO
JKabl+oiBBDNOS5EbqDliWweJvUN08XG9xgfAk6hRvhbAa8+g3IodkCa6lHcl+fJ
cC+39uZhdBJwGRfEJ7xXd4ZfDmyP+JTrjcfE7AWvjxUFTWUZCvaErRRx6hvvB7dt
k9U+dliiY4uk41ER6CeSZ1CdejfEkNwKxs02N5jNaGlY9HWG6ok1DASvma5/Xacm
RZzfIMtnSAkmUOVWTepe+ySa6hs+OjWyT/MHMzLZfu+UuI0mHD6/sJUG13wqFvMy
+U2HcpBTKQ8hn3GaENaMjvb4DROWtw15lhlU1Dwah5fp0Xacufsgb3/8Xj4Fh1Gb
LW53Q0HNCPwXImNUI1YgGdIXsLK+BsuR6tJjvsximYWKl8Dy6QNNkOuHKSxzuFdV
awVBc9Gc5rGelVJHTWPY6Zyi+/Kmw7oJRyl0EPWcKp10VvaxN8Bk3lM+eeKVXGBc
UTiOXx8TgrlZc/+kfvJSVrTQlf2raoMtnv5ulvQTVtojHZGYn5CSBp3SaSwE2Q9H
FI3Ig5bBi0Na8akslHnq/MpUoi3thySBV3AZDiUrHULLSLoY/CT7/JDcoAHJCHz/
HPTiyOz4a/uorHb2+vhlY+s+R5WxoJY3RQOoAqVfzic8qQJKtci7zrxCMJznhcfy
Ip0yDjGAH7F9H4HWhCTVMX96DAfQPPtkjGzKDRspSQjoGp5gEh5jiW4S03ylhdtD
n3TOKUreulm4DTJ9LpuwqY/VlzqazofAMfjK4MjkhnQ5QPVSCEiA2ZLgTGOiGvGo
NI4sm8zNOVrIIOipMxBT9H2SmVEyyKAOrmMHU5E4VFGZ3bCeWB+4UV5j393Ww7VU
dB0ASV+bX1udY1PiyUZWZdvCytCYslWM1+jDoLZfZ+3G/5PaiTEybODXcX0xTaiV
9tNKNqhwNm9oq00+sPCZ/9KWrkIg0nJCAPjKwgZWRoUHRcge8/4P6KOltGaYfYH4
mI2iefyo+y49BvT/V99Lu2Nyo86SxZ7n9Uv1WKQ2G0UB+HLQ4SlqQ1OY9gVNZT9P
bWP3wQo6oM8gzn5yfnl9bVzItqSFfjpU+erbp2ftiDpdKGRX9+Q0Vo7wEAM4Zz+P
/GdHrefOiwQZBaKc8WULiQ0WaaJHmGcOQlGUqt4sRV4/PyGb2BzeHF4/wAQj6KoB
sSn4EVrKnv9Voq4Lwa5v76UrNyXi1C7vBO0mKx0yITKvgs3B2876Zpo1puZHj31b
b7Crhdj4iIN0/RDWvwBlvwrM9zj8YB6j6YRxFO7069CiGAqpoCEbU7OXOnxK2G1o
PusAgl0bqTvf1d/a/2c4U2LPv8o8B/OtbtpiPzdjDZCfnD63ryHm6UndVMtm1TMC
fImCtGof4MXdbe6TIPTgi77y8dlJF/SF1pSZerSx36fR8XNMFhvwi9o4e3J6LZA6
HG6B7IyxZ18ooNHbP32j5WP0C3nxBBHMzuCi/37FLQD0Mffv5NUZj+guQqtvIGZE
5/q91KqThX5IsKAcYYsJAqBCYeAe/eyZG1xYxrz9i+AXFQ+R+u/ebbEHi1c6JQlF
wduyD+wHIRFT2upscgy/qNDSmeYmpl8hE6dTbOh4yZnMLy9rJUT0NQPDL9zHvhit
faLLdr3jZd0TAB4sIj93xHEHRH+tq3ae+2S+TlB36jDxptzuXmY53gvK2Jp2Fs+Y
p+LE/eHGmPpSPGK/My3SXHci2FKeEN/LZ2oLYPLpup7ruyWqZJC1VwcK6b0V8tR/
jeZpeDMbxMxF48lukVO+5v3NYWBxY57Qy8zo737OyWsJEi78sRf9Rus5dko2IXyi
0G5fFa6Vu95A+JJ7alvg0P0fVO6P8yHPaPf2woIwvBCzRCTKBl7TOFBKK+XhYz7c
KezUwE94/xN93TKWJbAdvQBfTPIUue2ydDAmJ+7jVXqBpzIwqr8ytTY8U8eUf3V+
7rKPvVb8seyl8/301guuJAFcvgyCtiZBonjp0reM3rb2XmG6uZYBpAvBxVfzokT3
0HYPz9I1MbHDMUAcm/RaxNoQbCnElCi9tYhVjLq0ya7S9w5hMxJN0HqTG3e1zbVr
x2wsVmEEOB609PEDut/MuShPuHBzoV6ZnGCG9Qw3r+6IfnCHRWxju+nujr2t5P53
jjSkvizl+IOcgRLkK65yZgMCpay7xQ2ybGDqgeci07keDbnWn6EtAn11lvzLv21V
15IefhmTQQorvN6ARNRhZkF3cuMPY1Cb5xE3MKOb305nQaWAu6I6azzrCu2tSE8p
ou1RomstpUc1JIO1Tb/hmVv7qOjAzNDPfjlHT9R1AR+JWBoGN5hHMdBPXa1zim/Z
k9UlyCx5skKWHEdqooTZoinEIHBrApBA6rifgXTPp5V/pINu+qeikTKzGKs49tNp
f5dUPF5iv922Qj1vEyIIQtd8AZTDjTYYQtZHChlfEplXgnaTzHgAwJ5R9X8EZ//M
kkpN8c7INgIFsdMmdqd/8KHHqegDEBt6zo0YrWk61RQ+YU2xg7iKgnQyYSXp7hOl
yNspQuCBKB5Nm/Gvw4+LQ4yoCwwomElkQ+JHoWaMtLrQDKirWsrfNzDhy/xkzUe4
RyLTEIgxcdxP/gRgl0pCFtLlQ3nPU/+CoiO+c7oK+oKxOFo0TbmkoKzZdgiGoKhx
1uGWZplA52uUuTeBHGG58xWzerFiUrR9Sj0dt8AZUqjro1xaWxWHAiDhnUUWzlA9
nbIy0q4Z4InleRQvqUCstThUI73uvA+he8Y07niO07sdVTKU0ukQ/OdQJyXbFH8t
J4X+LrvW2Xbfp1WKWB2WL0thy0lLgFZQP52gV6PkAPZlxxg39EJkBVjDkI3JeqQP
NUd0HjUb/Cx/WfxsjJbKLntpx2hrTJIPEfyjqSLNEIrIXJP6RpXaCfk6ku6s0Q5h
C9Th2EN7hAmK6aPPf8969g8rFlIjgPw9DrCEsYzJg9TBPW6KS9Yzn22zNr2tJu+o
rGtqUIWuiciT2dJxMnofMjlddBR3+JnbffYXs3S5QjjaeDvROyNCd536pu86kGW3
hhoqI2ZUjKS4eZasA94xRaCvFR+CrQKUC48T7JjimFtzmxcmJWdsHSPHmdNfB0P3
zUhkbyicGcgLFEcK/E40fzAYtL4+Al0pEjgPJj/G6G8oG0WxNPoCdwv67UOlOdn/
xUT4FCpPiwlDdhliHWkWWn6F68C2eVWdEQdPjCTMU4TEiC7V5I0siAOm18//IJa8
asnCpo7lc4dVdPf0/9+6DPWHKQbldvFnpoKDRhdtLAnGfUgjZJUt7W/x5Ix1Cwpb
zd2gx+YPFWYVyS0gNILWmi0EA0aiBLnpF4nlH+j7RK3eIS5IOvGD1whyho4CUZz0
OJUe+Vt3MY/Lts6ILwF1YJcTsrVwWaAWuGHBmkTAw+EkdwMf/sigQVxWw4gvjjte
ie18F6hjf5QBlL+TUCmvOnOM6QLy952A7C3YnTdxep/iw+iKG/Y90sYp2++yhHlv
Izu3tdBhF9sCf4o9l/dS3GpHIuoDs9XLE/LERu375qybcEbDnzMGqDQdC3wNe+Pb
hYIdQpQYQzrVkrjjKU9J5RtvLRKvDAAi/lN54CuLURVl9Gn7cxROAYJ7Jg9yFD9o
WoYZ5nmdPmrmKg4nU1JgR4CV/ACy0TdWq+uaJidy47G1lGgrBUcxjS8AauTHO5Vo
xJWEG8ri71Mf8xa41aP1XLgih/ycBEq42+VG7Eq9YSr4Jkx3PM8j9z2oj/90HAyN
kvMLHHSmEiWAxJ/tEWJYfPaI2U2r0m5s9/bJFchVGtxXgb0SJLoyiPL25Y5Uf/mb
u6qQ7RWh62AWpLJoDn2q31OledobvbCAZeKOAeIgjPZDh2MoWMbYHlrVYic/Q6o4
qS3coipIxB7F3JzQ/Li0aKKah94wfa9JIwFy06vtTxygV2+hE7uf7SoXbQot6Iu5
ELiFRLkmSF4BEr8xddZ1tFbVkCcPQH/GbSlk7BJuruK9PLAAVZzF9u4FOW7mE/7M
IN9ZhAkkDoVAge+bTo8iff/j5l7qvB03wJfzpmMMbeYHcnYmgAMBwFVmBvL0u1ZE
RR90wctOP0IWCxQpPWgZpOeQTBAYrv1peDbeYoxQaRGlz+Xelzk9rgnQrhOpbOcl
FTI36XcvzKWPGZKRTrb+AEbR/JgFZpEkYSKgLy1hVi7b2NRQ5YXVABH+e3QIz3z9
+gtWucDmUqAsnXQiFvGwnGQ/r9AiYkXhNECMSZsyfZPbi+69VVKvqfsU07In1pbt
VzUU3la4axxINfCVUB1u3PkCvMZeZ9P2h5O2VxzkSyUjjpswJBRCJr5K44xzmcTi
NC6eFf99jyqbIL846ec4pXcS1NGTPABE2yPfQl1rVVM7auHqWZwc07V7edMueB58
FdIq5v2NXvAXzk/5fPvXw8VMOTc4FqloAnN42TjpaZPfn+DijjUdLZh9cK3O3XMo
Z3hzeZ5roGF1kCg4ziYaEGkCe0TFFJhb/ixhcbe8lUxBga4mPGmkR7KPx0mAsJua
G/DTqMHits4rPh+/qCWND+KnhVbQXObpCRX8VL+H9re8O4AMWaJYgGDjz3lfmPoP
uHdJHzYJ8/MB9nJ1wnJtHXm8jxZdHEshP6Omr9dKSpP9+bgwHs+y3kTbsqQUe9iR
L4F++PaKL68xrc+iKAFfU4atd6xM8O1EJhcvv7VxX8RJygA/R1GPXhE2OB2LIWfY
3NYQRpdIcUsmpzb6tdBtobLEnQDy0yYGU/kgHxbD1eeiKMHY4QBz/XwC3xhZkTfD
nOQ8d1iMlAnhdw2mXNLtLJ4WRZnGArSLICCl5T1iOVhEjQgC+7KW6MOcLyESfx0+
7yBd7OjOujV13PMvujSKJ+NIpum1C2P+/HrIItc0aNnXgnM8bxWY9z7A58gWHe65
XDW5l29KvzpBPvwGHbKzQOoXgiEMDSKRgdSmDmimLr+ssLL4Ue0c34NvEJvBXSV8
K4mqtr9vHPYnyC/c4nkQG+2iLqAr4MYoLqo1ZJZXPpsJsRAnhN9dJh3fxAIINcD9
SxyYmxqXflCozk21M06LUAUmjGSgQJUe3Q9nPN3wtxFNsnMLcchndw77V5vwAanf
k4R5F4ne5HFwyaFeRQCzqbQUwbFIPFTkiHkg5/TitZVfoG+KJYEsSRtCKsMdeoF9
IjU1qVI84Wk1W9EAtXp7UH3SBBTj5wTg898B03+pBsNIXDoEXLTfM2cVYCn6I2xC
jdSgRQfMFkFxJGco8ZGndjLRuRGsBd1biLzXb3Ilg7uXWFs5pSiiXy1PA5LlXZH6
Jalfj19vl5pG7wUg5+gwOHnYVkEQlZirVytTs8yLAuPR8vQeRtcGRObm36dGRuVo
+R6rm/1UmFFFBaPFZiV4toH4PHF+F/5bdKvvtrgadpWqpyKXJFXz1zIfJim0n3rk
ET/akS18wpfcZowcMbkwa9rRRMlOTGdne4lVi/7guHs+BFhpnUlamO+6YD1XjYSq
+CrG4UEh3sHL03hA+W9rEik9czw4whyjSijEm+G65/r2pz//KLRdUqw9zsA+zM2o
KQGjy89YHkGMHpzHQZybUx85030Smo69sr6+xmjKmjgJiMOA3i3eWWgCGmqkgNHR
5h0rC1rOdZOgIFUDaV6biO9lSSFEzrbmFkuPSi5ro43cy2EwyaTQJu2qEl2FaLwp
P0I5WucsduOg8x6kpv4n3IcKIwX/uGUAIsyp2Fl6/hXgagCrxl+JeWRwl2vbOFKU
gHDZF3HxpifbCZZHQW8OwC3oFmLocKgn35cp3nx1YpxNa6xkslXtp+I20GrSi8H4
VYRu8nwdlngZoPQeKmVpic9bIxIFrzFkR2RVNGJ8iFfiLENdcz1Sug4Sux08/k6u
W4yMaCnzeMGhjk2eRN52GLhZSspCKXOXjoulFPdh5lXNVQLMQ2EMSPsDjtuQExYC
3pmpadTnhvKhAXPbO/PNAdBTWebswOHwfqJ/5Nuyg+52PeRE6I44RctI7ladcZNS
wN/urpzYQRQEd6j2iIZfagumYs9ZcqGR1UASoYtCOCkR2jf1TS/vGhV/27RKE2vE
3Q2C/PMOBOEp/mmBqI2Qf1mUujledx7AF17v2ipISzuOqRx2KHYKp+/nv0z//BQ1
ONGdRssV1TDS3ZeJoLbUzLE5OPxCvVO1AQWiXFmUDtF4ijcZowJyDpBb1I52uchd
7H6lcJ5AWntNFpkNEbdyH2keveR/NC/wIzwdmOPGPaX0iVilys/MPVEexy+GJtJx
5gbz0c+LPci3aoD7AIGn60JOo//vf4J13u4Sbsu46rjlc7f8EFEls2IJmb8+6HPL
OKBye+tcTHdIOqqkbew7PXFMA23DZr7fZBF9sGyzWxlwFN89OGCfWSjb7prBkxEj
LYNLZHNvkQWwwrtvYDu4Bs7PoxO9QZJDa67ZbBuFxKrCWqzinc0o7BOGK/b4YL97
0BIiNidatB6es2nPNW/Q4Ypq0kS2HsBDg/n4zgzrI0j9FG6lwlNr//cSZfnX8fiT
MDHRLNklnOoU92sDSukM8oI5iXjgnXpGuWrbAxHY0RZvkruBJdlx7kvl7dct6xcF
LRVRyC2NE13h4NOj4EyPaY4zdEsdtdWCqGiULXKyeDa4mM0NDoBQA/BZac8G7dtz
W9bmRbd+jmIqynEETggittjkQsMdWltyrshnjwQAtZo0Ru7OxI4w/gF96GwPSPa2
KK5EZE0GajebLRjX7mSM62krX+7BivLx8v0cPO768oQ1T/Sm6R49pPKysNlEMj3q
MpBd45n8GNtYI5MkGIHIqyPJ9nVXiARewck1xf/ii1DLgHlpcFwAn1D8BjdlqDuH
2kkvmSCHOdDhT3FeClYqNX/xtEEM2CmGnmOmCCm+krNLQwDkVCBlfBp7A3a0Iv0X
REzaaVQ72NjLIuzye798Ow1/cSPzvphk87L22ld+1fYV4EWLYI+MEpmSG6QxAl/O
+UcQKK1fTauEsE1Utylf/m4s8Phwsrg1G5E5gEO8uwOtGnnfYaMryi4OOrcuEJ5N
RwkshqSrpd97U9E/uqWkmj2ke6T14H2QWBcq0DOzL7FjS/rLk5mXEG5ZDtQIbSCi
319ORkrhFAP9vL+bBqTeJFZxCOqUnVH8gNwCXsSXpmHkxUGRqcG8IyIEjO063mfo
NqSS740h0zAezjH0lHv4N/30+vD/lEZMCiHmtUurxtEn5QHT8q1CPVOe7JXaW//X
k6o5kQO5d044eA6tEA2Etzu1M4XlaPJMMNO1AEjCtObPLtH68hJTzPIeU0uOYU1m
9f0SSec2srHkncHQSKOhCf8R10sq3ivm8y8Py4MFD15gEXTbD1Vq+uI7sS4DY06z
syo2YyhQoqSSaW/7cdHhvdx/eXsWyCW06Hs8ly3C1USCIu3D6rYAQMrGDKZANlAQ
Z69vCYXvJdRPGDoLRvjDzZH8XEYeSe/CfB1FyNfHrM0Ymw5IoaSvWeu0SuNyeRVP
960FQnrOT3caILPzWft2zhvuJ5WxWB9POji1deoGyQN/0jAs7VJ1YDxHgi5XC2fn
FRBEL6SlAbh5fWbCG/U+nwkOju1jiggMxt8URn4l8unJdrSSVHq3StL0qmny+58i
nyoMmUGrNoYrtOX8HDWsDSoDMJf9Sx6Pxro945v6APJ98HtJkG+SoKUPVdRTOkrw
9wg+Fk31pqz4YXm3sBRjtdm/DqQO2ffSSEgYV6FQm9raCf7n0+S/mwcSQK923bXR
YA38DwmNRHvayOplo0vBZovCqB6aQ85Fq/+L+7kefXSt0/wCukDpUg8bUbtCB1v1
o17G61NVr8QB+dScIabc/JhWv2NzLHPaycQWWVxkSxAywUjuEE1qs/KQ21F4dm8l
zbK1QLAWsnlhUKZYg9sRcmoWo1yUhZ3UFyoqs2+N+J+0BP3SssXNWV79DscoRfko
i/e3RfECislytvcUEez3TyXh7lErWVeElmjE8hm00KfKM2Y0ok5qY5pu8HKvVhTc
WCwwLRkuDamSO6G1vB7UCaRammgBNnhxjuygJ6yO7ESjRRYuEvWl0TRQPs2owlIU
B9Ir/dPm5YV6z3tuaWT95GWdc1SGl2Q6baD8lCmYWVMehbwX4gc6IFpZH6ZNT4o7
gW8Nvgyp49lrVGYiAeQw9mBy9QKs4uw2KtEJIiAtX5NXgaqJDUAzBKzAw14bE9Wh
p2OuAnd5zWYEeMqQOMd7WZXoFi8nO2zNouEZnxrb9DAFLr9PEKl/X0ONLmA2/9Pr
zmqGZbTuW6/hsdpkKWuOPk91uGSCxSH8V3dCUYifMIOBy8HKyYJqao/765bLwSqR
UkLpk0RQL0gItKGT7V6mNVRj26t1xVcuA01aoGmB1NvY2yYSno9uLUHtbfMfzraU
aBK/zVNE+ErNG2Bb7n7I5HZoJ2FdBi2rbk92Caz8yww1873TXGrRRg6csTWtxxbv
R+1IG4f++WW4CH0Fm5L/95ltJUbFTKM6VFgeHnX4KzCPGPvqNoua2g1pE9V3wA+Q
JRd9UMnrZZZ0ZJXlgSUCVARPOkgwuMwBh0Hy171BcKA4vSSu9SbS35z0qICXqEOj
cMgeE5UMzhFNyeV+aXEuArFKeRABEDRWokrWNHVK4FKoA8FWa/LTJ6gTVm+kTzj0
36LaOaIl/40D7SgQSxRugLTpUf+TiXV6Hk+521yl1ffNhmABhy1wNv5CmHKK7/DY
IRNCrTBZ1FPhtzrx3v/4rrWUWRUyM7TvFhVrpB6hVFE0+eF7J9vfLca/gZ+SrTDH
ysONVVKsFPk+XOkQ5/vm48N7gNQ7HTt6Cg3pawsBPlmG7BRwaiTVgaqtL+anrbCf
V2JBSqUXX/FxW0nNTEhI/piGU4zNThxojztibrKteNl5nuNGnJZ64Cilq1BKjL40
3U8NI2oVbyiVc2tLTPcZnB5Sv3goFdNNO7t3Ttqi9vUiA4MyunH3vkjnQzhbvIce
Wi+W+4i/27ku8jkQHyfj/UWPpkfcs8aJvXe9IerF1zFLDCQSeu6QRWVVmGxRn0O/
uqg8K10KzDIqYl8PQtqQgbk9Z7fw8SyY0mDH1AbkwESGLvCg6dSlusc4dFnxWqCo
68lUn4p5BzNzpIztIwsqLQakAOdJwSmd2PA6WquolmY+/jnj6nubNh59tExPe2rS
iop1rMIF/Hd9bbjfL10s2E58Hyox0IGh8dZvB9Jq3ylHeNMybAi/WzRpR/LGr/98
tkd0YCH2uSvei5XHHTx9TqP2C1//zMyuKIK+8vlxe9v+AUv1oYEyM3PRrwnSh3b2
7MJ3qjZbnBUmQ2vrnE9jLcOfw+Ar3r5+oVBW45N12mxV9M1pVxko1iUMlkCyJVrR
gxeJstak5qaJL9Hpylgs4W0vXOxeeZPPgt4cLzsWzJ4HhcFXFqmUsHJ3CYfZZTZ3
03gcYHrn8SrtRkYJ7J7upp/0+cjrymlZqrE+khe8m19P2Na3USoqJZFGTAgpdOE0
dfEtLyATt6J8IyUKuFpi+MBc2gTfOwegOYAs8EHh9EMSR0kJs3yTmwbjIIcfoCHC
rz9Kbz/9xe8s95vGhAjXO8ht0Olt/cOXBWEGnGDgLj5jwDA3C5HSSK64zHsoDYUt
zaELDzgu1xS00BJGElgfrbxOf2KqrvXVAmvdYsviik4D6UmKPBfq3MLQEbTtjlh6
IC2PbPkz6EwAqPgxVlNJtFz2e2y1ORbp7C+HU/t1BYaaupIpZk3WZZkxxIa+4tv2
ttj+51tKkpkgrJnbCQnQSaB/ompWtDFBGdtziK6c/bK2AESOQEmEPAeaqtUJOQOS
noJGG55uoRboQHS36oMw80vWQU7czP0dGnRYG7rsNhN+LdzocpIFuMZfSrsa+mks
OWbqJjdi32AyC6FHA+DRABpUr8kFAfMvhFQqNkIKl5y7Klb6BNccFPldb9kglw7q
z6AvPS9SwvBpg3uLYh/y83HoM04KYXoXPii3+FpmOa9T/gFaGcj+HblalSveRBWC
q04Ij3EkNEPwXvHh+msIRiI5gZFmp8PegwSoHdH/h1URg/xOSmq9RESHtl9XKMq2
lStpTdFlFpT8t1FDBKdYg9PWmH2t/hCvgtOxASMk0197826lbJLdAB61z4VhC8eu
Qxbh3YQQsErd0Ba58rL2rd0ysgKqTl3+MdBqzeRWM00K3TprkhqcTq5CQaOMz4CF
VnSdhrCb4z4XxG5vYdHnBaOW16M5L5iyrwi7mTSi4FZ8LwvMmcEJbRoMCnLZ/OBP
HZaJzTowhxx7GVjajnNvhxBVFpjXDNlv2j5Y2QIhihTRSdc2ppEs4Gu7yKMAkRRJ
15m1VxKNIhzV11V/8um9kWt8ImOGMIAlvkFfSgogdob1oUxuOn2XyGsdtUbVZlWw
OMxBAq2/uO45l+8omc5hnD252lBioiK4JYwcsPaqdAwXG6OjWFknJteQGoJ/TOf4
MZeP2tDXECobOzZDZPcK1E6jZIRgK8m6hj92A+xcJs0OXdlpvgI+7sZEe6Mbem2b
m6+Ud5o+d77gFfeas7lMhfG5dL7+NqvkDV35OUl1wpcB0k2gbOaoR3jTVsm1xRZc
H8VHdtNnQF6a4RaLkuRaypGv/cyT6hdHUW4o29p98PKQoVl/BD48s3CVsmB2uSjd
jYngcuf/LhX9G4CQt13Af5Yu1CpZsCxaOLm9IIIFl9cTM/hTOI7W/MB4GL5mcyJq
a54brKKYqZKayZp84aqrdN9/99CvSN9+54x4W3Ixs6Idm9h0ld2hZ2dxxivnhgdi
7JitmY9Q16lSk3gBQpkYsc9yFjXhY7SSFFqEDPsV8KKU7E4cEJ8EpYzUXfAcrisZ
HUHQMyXCjIv9hfSLRm2knbMZ5UpyKfOiGocRM+iH4a/S1tbLnHhRQGJyN+YPT/EO
3XDTC9wjqF1ByJNzAtR78Txdr3toSX32ejiDj9MdmTxbBNcsr+0N9Jf7I87aNOfN
Nn1m+8pPgRsBDRQg+trfabjzngez+NjbNhFQSPLM81YwROJu+eNJEBAtpv1M+RrR
TYfVGIQo62DDg+HFVTNcIXcK7Adr8ZtGcpc5cDKJRuwHdFWX0JhxyOkmG+B4nS7u
Njym8w+m7Gb3Y/HEKaB9WbUu/qnp3sx5GvfjRnWyjwnbU7pwfFCc9JIqUN3UoMO9
X6owwJ9lFAzVqmUx/O09x8j4ZUxMvb4YDjnES7tiXC+rQ1Uv5/xnebp6jL2Rt01p
fTQAKItCcswd+Nn4ztWFebA5O8eHepwN5T5zgLtlP06VACrg42JKSoQ8ZZO2KhaD
HL9EJpoBoH4p5KswF5UIypIaKsrhnZ4s3DtKqce3VSgFqJ28WkUCcB09ywAAJCrI
tMjaAjp36bblcCsX0PtCSaiL4+WxKt8k7+WewA3TiFHTRj47393THQeHSA8ePpRk
HpeTQ6XiJxhoWAFhM1qBE+62R82XvvZRmcePZ83HtZ6PHM4LIPTsOSwcwp/+4dn9
NxXG2NKIjqwbd0wRP0TReApjHOnKQaejdNsZDPxXyGsr/NDuYdbRS+vlpa0FOVlc
8INXP7RUN9omkbHQLvtylnkoy4rF8LDvPTK5v6bGPl8O/2seVGMd7eHxVQ9w+Nd1
V/GxSFCXDAKCxliXjlT0YaEN1x3i+DCZBhsFzu2hxdAZn6RXgR0hkPn5bewQHtAm
PgaYnxGR54Ps9HGpwm64GMuPwRsi7dGDpJnH9HhjQFqR95+LZQ/temjnoKJlxZ/6
mG/9DZOPMs6WzV0s/aB/9le7ZwSgEZ8fOWHInwiCvBFMexbGOzNvvaGr+1y2YpEv
U2kZheJaodZUu9J9xr8pfEjJY5zvj4aqObV9tJJN1S+axD7cT0ze5SuBSgiwGDGO
x0OMamj5ZBLUbwE07s8HDBBEBamC7aK2jH6i4M/1ZXQsVmfMvBiM2lmSFZ0Jqith
jCM7PLquGx+egiFBNkbO6M9Eq21QuOuMVJgqKvdGC1VsPA9/Ll1RMkIV4gcIIbPn
LLcFlfg7QkhOwa/tKrxy/1IK31T9oC1RLOgEIe47umhoBAzUdIRYB6VMpKaeyCaW
VNqhyHnF2isH1pWYdKuuwo3+beP0R9Wi1itc4Exyp25g3ysCV2iQUBys+BP+EF5n
LB4uDvhupvu+OVbiZRpdKdFSS2DpAQMwvjre+okELOLqk4hAeP8v9d4PJrKopXYG
gHdLiiTocL89OZJ60qM654w2eFjb4aRLVXstIDn9pd66Ynr+YtK/ju/MpUl6DLp1
LGoTDhJRyf9jYTEr+hpneO2S7YUz63pVCeRAsTDHINwZYBkSfawiEiVyG/Jb18UZ
UpDUpXdz2UJn163dIlyqMlBdcVq6e/VEEgBmA3inmaPZw7BZnZelTXL1nkmYZP5a
mB2/BAirnvu8VKzeFV61mjwuxVw7KgtW0wNbCIY1u6J+Fu0WJuu6OSE+1UMgPDk+
mAB/tWInib27lB9rm1brgfT2aHC2xr8Rqe3nlLEHou9w8mPFDJJK9fB//AqfNJvu
G5JQRsfb5rSBrw+dKLS6Ggx2Tmv/xW3fRcoD5pKFz1m8nzQhHkmQM50MB0E5BBnx
c2qna0xLaoS5CMWlzlsTY0hWKRNxeFaWPIE66MM9OcMfk2r2j174pqEetvg9p2az
nYz2nZ1lKQ5BzpBGV03H4dxiWtYFVb9YQ/JvfOTcGlc4EA2CClccbwaZmHBtwBND
YtUy9gIg6f+F0BliWfaXzO9mKG995FnJPPZD0VdPdLwhrKFUHYr4yPbJ5IoCvIqq
ehEQ3fcfgTWeLczsSMN1wp35GnSy5Ikax1o9mSs67eFkSSIJOynXNd7rRZlXpH48
At0hg7SI8Kwitk2fw9zEpjdvzhAQPR3e750zd7Gs2OSaGGMd0VoQofGhDoUAGYfD
NGoMp5E4fOlApArcBAHuGxXWzDEZvNtL0bsDfBx2NRBfMXQWXz01l6/2R5IAjP4m
AJW7u88fbZ1e6QK0eDrJMPGGt+mJ2IqmCwfXahYY3T8JgAcyIgJJ9vVFeG5pQ6FI
wgjjIIqFpMx++TXQZiMLf4mkbf/j094wxN8rZBRvKttVS7V/sx99etrnM2jLDIdZ
TSYeLHqNtYdubl9iUO/5bf7dv2i3NV9CHDCOMPVQqw3j8MNxhfCOUxX7sJct2d36
iM9fM6y0fGdIWoH+cODXqmhYH2h+rkm+bHDvjOviqldRO7euYoGr0x240ygkYjFr
zlIJyO+iRT/i5qHRMtbGpn2XXYQkyfc1wOfv0J8RItu7BzK+1Gbs+x/9/DoGIN3n
db9xdYE2IM3MYWMBy6NvXn4wxQLohbFVVonE35Hhv65XsRPfrtSTiZKWDIxnW8/3
XirqCbbi2faHWlMspAJx9DOoxqnXTIxDxApmG+aLJZyZdNhCLtyEEzSZXsl8Kt3Z
0nvf2W7JaJ9onCV4lEH1Vq8cYuiKDBSsNF79Rq1WuxrxzLTqi4tPHsJyS01ve1VD
wUCYYRhl5O2sWJXUqWhHIZS0FokEM3wkpG2dUFfzYPdOwXUj54ELWrwIm+7+jRqO
NsAZs9971nYMcGKTdGYU/Jl2MdYViwud8P8M0urGIf2+VmFXrH6PNeWZBz/u+hY4
eotRL/XhDp+uRcwckvQ8S+a9kspoIez1Yt2wwh2nlOHfhQQXfrm0/5ILTepU6ZDJ
y7QayKfwLpF8n7PmOCtOlmc9S3qZz1H4dNaBWGHlgVgnNy1Z2GzvLpvsI5H9ZDAr
OZFTBbO7loUum8tx+yhuDkxedSh7RIvNgOR1FaOlGKKajI6czvRjAgFjIfhpA/OT
U4AuzthR5nPnsoV6grxf7mQF4AouHuRVkkAq+14L2WKKe2JhvXi98t7u9zfqNNXQ
bIe0tsLD5NiOinrLY2n85DpVGHVMFwNKS6yxq2tCLwGORuCbcq3Ccrrd+PrnERDw
OEKf1FryFizTWS/7wGKKg1tnZH7UJUUdtAuR3M361+6aMtS8BNTQGJHMwfUu+hs/
8dLZWVUGUNnGVRqrfbXbwMTAKiIRsq0zQ65N8FyzcX9kcx2yXtEmLAYeH7oNnSTt
/nRnW1i2btkZeVS8QWOqS1WtNn7wB+O4kYIJDLO+u8/lovjks62tl43wzDleyLkJ
synjgmgwmVcDd25LZfxBUXwPzqymGahr+I2AptapTZexa0D/FdAXZRezlhI7tYoL
JYYqOiLR7k9J1VsR1JFDW+sx+lQWR10Qgqm63+AgUOdJW6OQG8tbetIpbAD0Hvi2
2k3dQ2a132zmw0+sFKbAfdv1IxfBeRyVeYtIEd0LZLEAjAqF9Z0901dURP6PgXn8
xOBERaA0igQgq0NzCzAqJH2KciBuYHNx/jYmstHXFHYDHgG/YJ9PpivjlsPYbLex
Ch7u9Fu4Hy4YylzY3JmTdn37BFRs6ypcAoSsObNB01XlozfJ+ct4lPjRBWt9fI60
+UhZxrDJwqeHnVQGApm2v952vQRv5kODjuqo6jq+g162idpt4K11DgFe+n0uPyg6
mD9B72hElMJuaE90RHnJsDNhnDdLSceZTa5+AjeMImZbKNRA3o/Dx/5EhO2sXI0a
O4R2k/hlSZXzgRV1q3uVjXRZbfsFMQiL6N5u1onCUMzk62bqcfCCeaFqVLTEbFNw
QlrXU2oyngvrepwpBa3Z1lDX8mfisQLQf+pAWUMQ6Cx9qbYtLe++PrBxLjX/vBC8
mFVUZL4wEtu3XidvWTwzRhisXm4kG7czMZ5cV+TPucjg9RmVZlE0wgmJxi3+5M26
QaUg/WPy4thYhlKvbEK9fuenNiV1tSRK94/9gAUxeGt0IK+zN39LPjb65DYumtxX
AIdAyF5S03v72MHTo7NNTmviXjkKrjvnJfR0nO+YwWX3FHVoi7P/qCJ93eCeCEal
HEeyRkp38D5OlIufB4GQcv7UKDmwLuEl7q4Ilxjg4YifD7gkIgPXqk1hPiLS4PIB
aI9tDu3WbHpJLB8RE0Q8TgHBqEJG8ateM3v98B1Slf9JnQuU6ht39jV3fwPSmk5v
RK2FDVSv4pcZbVAbp5BOTerhDg1cdZy/9xBcmAk7RUVFAYMl4K0RlBkVYqA5DfK1
98z4LI6iSDSRzSOx5LIdBzHVqKAzwWd9dCZdWZKv0b9o68VuI/AP33IX4UkrVfG+
sT2M4dwnyoH4aJnbM6Mv5ZpNXckTof/18HVJqEHrR5olP4v2JtJjhTAdYpykSYtK
fye57xfO/MqY//cOE67pN3aBH4oMihFRo/3Ut6OBoEUTa30DaXAyHF6yHAzFbU8y
eD+o+VEPx6HTQVjCvUJiDyqpZK/ZMcDTYGBab6ddNDMI0j6ga+i6lRdgNMnsXD/2
oMzJGjcuD1Zqfgk4Yk8yffc9XsNmE5ORm8v+XKoliQ0bxntVcckV1ZciSoJAE+lY
tW3xj3mY8Y3rWWrrRwthPaUJYwJS3tZ1w206MxaFxNjinjBRiNm5tzyRAUWqpTwc
iuBPCdMAomG6vCa7z4DvgR7MAvWF019KNfyQWw2EQWwHISfNSfP7TSJ8SJIHFYgK
jije3Ek8VggK+5aA1orDmePGN+QZLosWcuSchYRrmmVa7Ov5c8vmJRTRrZBrFfOe
vvQ+3tenqnmdfGhroHzW/ZeETjoxtJgm7Tvs2h3XLmiaNNPUQ+V8RlMdLww3z/XE
fODzJUFEVwbb/0/AikO3vpHd6iRzfYcEG2VecY5a+zaDyL9J8BP1XdIXYPeWIuE+
1ioHhYwJMmvPVmmEOLf+7suW+BkPiEUyWGgjok0+dai2GuHF1NfoqBXHew+Cp9gH
Nh5Q2+mln6/6VPe99v//+GLr8MFN2KC0MznXwbz6aofIkn0sGdyn4WXJ5PQu5uOr
ZazEgbAp/SUiGXbLUUkXdrM+7hmAkbKqzokp+07p6iyc22N9wbPT8IW+4hHM2je+
k5tevrCz78njIoL7RJ3f0yGfQdmRUEiVqJkiwwGJAIPYLRb/S2uXSXHfpA+h3Kyn
RYQkgLksuAhQsFpaRlktrujQXU/J6wIGjGZaDqa3pkd+eaX6Mpy06hBrbKXo1gEJ
XgTXJoj3dh8MKI88RlLV4qBGlJledBArROyu+1eUeuJVMv6hXEXXwHPEcGHdNVoH
WdR4bdLyvMnoGxhWd2nw1kZE9vvgeUnrMwcx/LdhPginEnAD3P4+7TVsTne/cWJY
dzTHqODMx1RygJf1rOEkxd907PAwBpPFj6YflnFUYS9e/OrPHAkJtexCcJUL4ebv
itgUGw411OAUd7RM/5R7QJwHM1lGI4GuBAtYDSzYveB1DrCbSbMeox9x/diUxmjf
RiCqrk72PUg+3kGzIwSsN6wtQCmyWxhc0wZxIEe9EuTJhcCuzPgdGbom7Ip5mzEi
JoDEC687Ku6/b6q9sBHtbH/oCglZEWgaJ4EUjDqtP0MJ/8aYh/VnDljhToKGh4tS
Q9Rz/CtDsumpLaDnuquK9Q04KPIt3iUT/uOy5oflaEv0vrQiynX+9MN6jDd36cL8
KmNUeaiTFNm5cCdK7A99eJ2fLTRtE2HqOislnBJF4q6Dj+fKWExpmBdmVZFqOwNE
ZPBKvUu5cO+/t4NY5I89lU60HHq2UAk5qAtqRCrCj9qtf8Lulmwxw/WUIQO4ouWx
k5KbeL5lwSIeuIVjicIT0OEjgO9mK3GSMsIWVdbgFYgkPyY68YmU9E2w5XAoumen
9TotbHKuoJ18bKvS1E2VNF/0+Ej0VjnDL5h3B6nSLUjSym8J1NLCYeVq8gd64bMI
7av3mAxATRlEAbnjXaPJpKcsdoTtjkL9uphskTeN8lUXYoYu4Zm1kQmSv5T0fcIg
x4uHl9gdaEeQblTNg+U0VcioYZNREEZF7LjJ0F+VOSNpdujHSRfXnA3OiAqx5GZh
wIUB/1p14V7Ol5iICfTrKhls6EV4R/eMz58ag8ZCpbTP+Jkq9UYf70Gpry3siO+D
ETL3aIxE+srWzE+dXNR4wUJx8UFevehaVlzbFxjhJZAj0+gl+08YR7XGpQV8NIMw
SdbNNrx8Iykq2z/4U144bVrSfCKyVGL8sq5vAG6U972cNhBvCzAjmMbGhbun9t9D
Po6UF3OlT1MsrHypjLDzGmplTeTyqg5NoqdyBRCwt1n2y+tyAT9EfM+hvezDd5TY
CQJ+DskzZfi1EiOuIQRrXn4cNkG3RzcsPPckOBpfTC49IeGDuTc3cOte6+urUPtZ
+efN4TfLCwYr6FRbMc8cZSEcKw9llsZzuAucDYoBDxTrD6aptRqBMXxNee3aV4Mg
Ch28whghirYIBwCJrpjrIvBvkdLHJunDYPamR15JHXdrjrRMgf+yLAdAgMuocVYg
4P5NLD+nuSSyoC+JO96GtOS1qv503LMLmzjQoMBI/mW4tp6zA65Otv9NpycztbtH
S2oo3wQB+VURlLneKGIC3z/LgUN4Q1xYtoMRqgjwgstH+SweZ1xTtG+p491esXzQ
07JY15rDk+XnuiAT9HaQGXT8iYvCKLvZBRvFSzOKnco7pnQ7HdrNBG032tb6yqu7
UlUut8bBBAVFcwi6xew9ZHalQO9fjaMwBdPfwJbTlaFZHX5VvkjZalsnPg23Phil
PZTJpPI5os4cSvv+vou1kM1o5NU+T5EMwjR5vE/ocPR4zcNYZCPJ2CjUG4m2Y6fy
WSrIK9qqDy4hcY5KX+0KuexAZ/OGK6W+DvY+4HLDafvluII1lzsz3bBj+Uic5zkg
0/OgC9bVqS38/dJqM7w05cxILAXyV38jQTThnZd0t37Xc0Rf3xm0aE0zYqJDdJwZ
uzBuTrhCL9G0YgcvYmUWUIj2CgZW9s3OU3V1shvUDvFQbobWD51NKt/Y8kJA59Jx
6tO6Biwbeuy4nVfaQEAGiAmcuwJLQChIYSaclROuFH+/lyHEaxOm9IJxSJsgpiif
`pragma protect end_protected
