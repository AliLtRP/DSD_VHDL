// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:35:57 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
osflYyXoPK9fa4dMnnQM2GbLm6xK4UWDsBPYCiDJeUS4hCfxuYiHxNxJpbNRXtVO
wRy3Xc7So6rWTPCu541GDlpdrAHbHf0MNKvFcoFABB3HMqxd90JhjwIAdBWtsvZo
6jKpf53wKSqBoeuX9wkRq0MHGymapU5EHg2nLlUJe1M=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 37920)
Xd3FVOFEDzSewJV/rGnyxHBSMMRvHq7CskBMbGdRX9pwLzSpNdQMl+MRQJguBBwJ
YXjJz2e48v8bNwU8L58QFOoma1UW6SMo8aJugFTGSP7pXawcEuo65raoTbMZaVyz
15Ay/4I33Pc3Fsqk6A02CmZT9n/6J/WniuOZdthy+WDdNsoJofcbXiiUxGwxNvwk
Z3hYrP0xk2ExMTRY9eQk7IJDiTLeHBuqUTZe8qM33pg21mW4sFj51KI10Y0/RS1O
DuEyvJCUBl/TsYlxjBqJmj/GavH2lvyeQZej4EX1trRftKRMbTRXj7dKiAvaJA69
sZVUHjcERTmJaoTtCEBMn6wIL8NRsQ956gGXaVC8LdlCKUrR8vXERDGHVEM6brHw
PWlQnz0vZMFHBeSZXv6Rsa6W5HgqOxoA0Jifr1T7F7LM+FGRaHkY6EYVKTbiKH4y
oYXS9C9rDf3wGOX6ptyL6M/7P9AiWluO+GOND5GMTU3QFhazbfSL/mw26II+HqYH
qRTVtVr/JWQ9hBDgcE918cg+cOEl/ZySvQyHhPgsD7brXGvx++HTv/Wps+eSPA86
NbUL9gENrJQ9ksg0DtPqnPxvQk1pZeA4y8aZ2faWplClCL6FwmgAI/5dO8JtDNLA
2HGy5zwps2q97VKNQyZKNKo0Fm9KrGG9pJjPspRCSmTQg67tNLR4xNtEBC1hrhU8
MgcUzyctVPFfeUOWxNcWQvgZ/ry9EeS0abDi2jAKHtmwmAD9Lkeq6hXwHSHjf9IJ
CtCUBraAtBeQlmLgL5O2u7wRqi0ynYnXHaTY50BzD5xA0MqskfRCP9qbT59OK3t/
hC4pDw5dnoF3SgzfK53BHO84U+Zr4lku6VOsXp+vxFnnP9X4mBknJgTJKb1WF97x
oXIvBMrKYPreLweiD88fBEumjG2LiXni6/ikiXTY9vLdmCqC2ocPxXv8Oebb1Mrm
bcUKUJbE9rYw4XoFkYameL5iKg4GgCZvVuIhImeOtjSpoyLWOy/N5bIX5R0pge5c
UUD1rKwTHEa+xCvqB+VKLrqT4nDrfgaS5kX5ztlDd7qk+r4VImKUM2S+YxHzMl+7
YbdQDxhCQfvOdbAmglMqQCq9Er8RTAHdOVKT+KtFD239yONE2TaM8t4ozuzV3cdF
qnqhHN5pBzqTafHetDLvcfuk7kUx9I/KP/SNta4zWpc09wCBRjxNGtGvSH5/vHHT
czOUjvzTQq7QkIjbSBFTI+1Da1DLt7en7eM3jQxaq/fSPAlWp+Y2giV15ggLg+jk
hZrZ04smUWNuLlbmyeWH457jXBCYvy/RQerf+cw+lkni1eAHscNAV7o+qXcGXqL8
rXDsVIIhMjmt0KQw2bnxKYZsP9E/v3ppsGxyC4oKYnW30fONH2iTL1G9ezAoAWgp
3YNpYESjpcptjx1LNw3mL0Q7YBUycNt6SHDF5DFJy7IfJ400tUlbr83okYZL/K+i
KLFRMZaBahk/3OyMfM1tSiQj6VE92tzDArXSVPPe15dew8CjcqB+LuscZo7xSKdm
RMz83mlYzF9sVbQHWgADz7SQI56MQG9YgKeNk7X+nOCB1M+Z/a0XXxwa0zAmm0Zl
qsZk6sVYczHTx/5mMttDldpQoNfLcHBV9d4V7TGarXa5/xUhfjzwxOLQENbjYnSO
o/DR9o//klGfVMoNH1bOP5DK9oZNtjjZJPInK7x29ALG3/9VAdAdAPjVRYrMzIgv
KM7PYfiQA4NfyLYyIBecfeaKn/+CkOa5kbZwBR0PYbBssiJokntBOkWbk0xOh6FW
FhTzX19WAbZjy/ZJwtmBWmw8MuxbalYmhZJlUz4m4aC5GNH66a156KpPT2oO3+Vj
hzN/cUN6t/ZaKftovaFFjn+OmwOkeJwP16yH5VLEIc0lD7lwOqG0Fy2yt1GcU8W6
fRbTNOnEyu5t9OnIC/BJag69s6Fg/+U9euHaxCZ+MGtF0iP2zgP/UGJfSm092kQx
/Gk6vpSHjc52CcCSyAcQhTmiIlXhhfYj4xq3rDWLz2a6FG/CM3TYIm8yVCtWeePP
9CVtKEvf/mngB9UR+gm4wpeCagEyBDHDoJihAnEkQYD9MHlTBepd2tAjbbDL6A8Y
zLqkJSwBdIIVxcsVHUGYV2YvM70GEhecO4En+FIKuWjGpP74pwmFE82Cb4zmLHh4
v7yrD/99AaFdIU5LREhJatLH+/YAmi9OeyHPGyw2hpXhN97rw2gqXgH6ghiy3eyp
Z7MuLBvgbtu1SemzcXEMDWlrr+ShPhMne+iUHHuQx8H+MuCRqe7IVj1oNenWj+c7
dF2+dERe3/tqIYLTvpMeoUIRsh2qqNfEl3imGdnkCBrfq7OQ3aOTe3yW/OY5Cemq
FYbxyHqBpDxVnMY6DdfKXEQHPnrojLPRqvTKvOl0finrnH6vAxpGmNrp7mZKSzkY
PbPrUWy2uxvi9w7xxp5hMLWKeM859APUiPoJBXXKE+vBk60MUGgozj6UTH29NbZL
nHIQdXZYJpShrXzRqC1cN0lcw/poFbnlMqiehIs1LEwsYIqBv9Isx2QarHhxGNbA
pl4zj1Kr1uepp8TIwWu5vhukO3/SRWZasMMu4QVgL8rDrqtzy0Nd+5Kw13ZbAizI
j+X91q1yVnQT6fZoZoYSBRnCuCArM6bACA8Vkji9oHLe9dfMZtgj9PlwlBLEWYFl
pdcl/uRghKWcj938I2J8vSUgYBqa3ygcFuehBKd3MZeM6nUnKx0ZvAOHZk6PLRIh
nKuWowhv0L5hKkxss65oSYCHISkK+02jNsjSkxC7PREW2FFNiyFikI/9ruvP2xmr
Y1j4p50+CEUkR+FPsoVamgRiSS/0zjYW75ZjFieMz3+xEji/PSx1ZkjO3CNYQliy
drpr71eDEnl1oOUdfTVIdqk7yT7aDvvuH19B7S5/pFyRWkX37B70+wlE0Ik+u7NK
yC8WITe1BPvsx4bVV0b3Es6rjW9kXWcUSpa5dccbh9IaILILE0eTNWfY9MqPbSh/
qItzqiV9jvv9gnFq/t/H2WMU0d9ZEIhu9Cl9sDH73GjDbppJkXpojIBYrK1m/58z
KzZMZlWykw0oZav6bHs2crPY5w6oqUaSNiVtHEzFFC07uJDfC77rPDEpWRI9iR9T
5G14DvwW3ul8UiOwYSGKPVWhqPKLNHinKKbX8aJ+kBDM19yYtjQtCBYTEH+D0bcq
4vbWq80tQuds7rycDMc8x5L9EcYc6O8RjOgyoea6Xwp7o77hLsg8ch4aFhUMfyZ4
B0k2AxgnHFcqNF4eRHqe45UPEQtqtmd0UGhgAwKhA5O/g1vMnuG9P2lUf2Ct1+75
PklGk6u9CsB0iVz3ryomOAmAzE9P4Ogk7kGXL23rFYpUbkE7N/CIB/Ud+vIqH4Ey
QOg6F3wlLXOPjPg1zYatMSWsULNtVPf3dVacTzLtZZQsNEJzhFvCVjE2edf90R9e
45yC3vSwC1y/V0AHHTTicMsIE9nA1AqOCedG8sCyyr1a0z8XPMHiDOk8o7v59Vu5
x8hj5zNEAR3dRJ/uvhU5K42zyyyiUuhHpCWbdA0n/I6eYdUHXlSezpPhS0CShCc7
IJmmj1wEIbGjlPQkOUD81oD+4YDcTkEcXOiAYFFO9hg6n4UmofcjKDz6aF0B4hiE
y7AkTios/V375h+HylyKjZjeBp8QuVInYISAulBxKl+Ai8IdxIYrbhD8RCmLJiWv
gnqtw9iIqvfkZA4WhAKll0XWzfULO/DF3NF/PyQBBeFe0RABcBqnuQMqLq3kMdPy
jiQzEAvaonhQdWfN1BW1L6IGvnoDjXWjG/dB6xQetkW8ntDvFhSPh15OqQ9Qge+J
MsJ5KfiSBex/UVMCQCXHlO8rN6HpeslcC7pqRrhy+SPL3Uy1PMChy7Rq8B9K/nsb
fOPtSKMFLGZ3vXXswAQ1fkDJN4F1+TfXqDUwEnfiabObRV0/0360dHvAZmpXnc8i
aA7OFW448kQC3LGSjMLHy+L+IYFZCJv5ZkR1CtVXmmepOpWsGotH0S2k9mPbD8lX
YgJohL3OWM6qaBxzmUwh9AViqWgYKxop9w6JRPkF8NHQ2dE+4NNAnF/qgqsaZDrf
ijskObCmh9toJd94cHyL+ei3ZpkDjXauv0bND//7yHr6Id5n82+NmYW75BwPsoGK
GIQj24uZuCNMyOBZqKDH+5EZR2NUD6yj4wZr1x/zxusIDmwt271S8jUOPRaYeBXu
3Yx1MvBRrOJDyir3fzaAPf5ShgfWWEDGAztZpUGy9qtnSB69es2Afl5HvOHRxluZ
/khVeijZXEnFQjwH+mZOkh5mSY6U6GxB1DmdkOt7Xxqmvi0MudBnq/ScsJFDx4+w
/VWs0DMGN03GjHvShFRajpYSqSUTVwk9PwDINre86pZ1CBQXMMDUVRfixxR4W7CM
T1o/giRkz2eV1j6MGkFS6CRzSkjpYO1z4wRtO6hfLr7Jvn1gjoBGQdP9UFMmnCja
iacirPuPAJrGagX6nG6m4oriTljjmOMgCgHbfc8F05jl90UHFw2RL1dWd/SiJCWY
z+P9pvn+isLSsIGhnmOWLNJGPjxSKxil2X97b1X1ZpVCcABLYIMzrWKGdJ+yKhJr
F547ppkWAFajgsWAqSIRMa1GXG8nknjD6oxximmrCHSZUSF4t80pxKHSiv7C6vRs
7uKZGFSyn5Op/nSr3Fwc+EnXhM67vOtzyGtHFQ0HpACA853XH0jgnaMCkCl+IAhH
t7xUYjG1lvr6fliiBTZgWgniQ/cbMyi+jMQ0hy5EI8R9F9HGpZJbwxzPB3Zrr2w9
lOO2bKgYtqTlR4/JoyvznovooTsvM0c0xwiLwCKz76t26arR3p2MIRRHIO6Q0WRp
t8tQJX+LtYQTnd0ajesFiH7ywRUkLqusH60NPtjGUCcyt5THDewOuiptL7yejV5a
1q7XheRbDqc60qNw9RYGV17TltWWLMLJ7MbjnsLvu2FfF3OWtAKhw5RLZKzqnYpc
piZ5E2lxGY7D/4yBqnhiD0UbSm12IK7Ei5ISCIG09QiwO69shgnO6/U56fbBEBO1
mKUrsPx751/kqxLStQNCvSSG5yrsJzegjocG5EnzL6QFQXjJVitNpNutYEOazDlJ
OhseHEu3+NS4BMTOGnFM5ljebqTWPdharNSIV4um5SDM8Qap6MeVHPXzuLQ39ZqT
qG6796KRHZfF808VwqGL8opFFCKXfApIsoNLRdNCH6DiXx6QDQufsOHB+kbtB806
DZSJdsPB/k9zhyCW7oxMKtmQHmmIh3E4KBzWkS+HAK2lQHaT+T6CAi6FLIt7BtUL
NrJijsbOU9ytXvnjlAq66i79eLw2PLvAySwVyN7I0vimvk+tsAHqIBpYmr4F1TUM
GFp/GDfTnvjMJD0QotdoJoQxyJEVE5JLjyL7jEbsWSXd+7tH4agWdiRmc32wcw5u
bi22SpJnf2BTPJI0AkkrGoQF46Il9VUCqj/NExl+gGD8/RaxBpjMg2suMlubx+Ea
8Gq0qqDevGt8OmberOAgKPNLWlw6+V5atYu1zhjrs6wvFwhb4w9LJHNlRaFpz3G1
WKvvhQD9I6gg1FIIjkBMYN6W6aPfvP4KENzs541Qtdux4oU0TF1wZIDHw3+dU12A
MxUxtnv7RYuUArw6iu3VCroBACyMyVhSan6fG5/9toWLzbTgKgE7P7fPRNeM/I7f
UG07dPJz1qWfTI0HiifelgGPIUqdMQY5YPpZED1WJ+Amvr5vcUfWybqBHsreQvw3
jpMslY39PwszI+ObS1wOsoevXU9OFckPOGvm6s9VlCZm+vT3T+60myjIdOIEAPXx
7gFuUtzty6WkT7lXrPPWugCc+/ZSM51hMWqzH/7guDigJvObchru2SLe2SbGEKOC
GLXU2O6W1v1sw9oaizjjbCFKMlR8eOwAwAA6vs93+bgR8ISHKPhYD4GeVdxXulLb
WBoNyZ1Jyvjh7TTs/iDiFOXTiOosTCI0PzgHsQi0vQT7Y0lX81rqKsVF2GGex4RB
uX8r/RYGvPpdoXWnF7//v0Mtn9SToxlxcu67Xwd+QyZnGYiLnkD6tI8T5QxVmFJq
bIrnygw+B4MjiOxnzmdmnG//lhV10A7LygaixTKEGXdc7Geo4IbDpE1UyuoN2zOG
7Fro/oXq/Zn+5gn6RPb6KndKMMHiuwfRBbjscpOPzu1HPnNoM8J+1RtBOn3RqlYK
0QnEPuA2FUbCUnxcSBChLTOA3DXmWHp6fwOE3AxN3fCXUYV8pdS41dO/a1og++7p
8SKXcx2Q0NMPvR/8uwVddlmsjlJsG2oISqIc39A2xtR4Qd320s9aF13l/ZjqpMbI
/PjmApgEDjiZELjXOp6ylUQ06MmCHr+SjU+CAL6L1lPqkvfK3VeZoa0m9CctQq3v
b8Y0f2a3R5CZvJ6LNvK5/CH4R1Srlv9FAPPWvL2AKFpdaimXuYUV9Zfpw+YuakYD
VliKIZ+TTQsi3I1/a7AzEVILI3OCGT5iOXLqjSgz/yriuejw6DeJJcYv1fNszN1F
sIv55RDbNDOklvfyTxr6Ss/r18waJRZxRTZn6J7BEKl5D5SGN2V2elM4gWlLR0aW
Q5BYxLzSD4aYAle/btbISIxF6VcLXdH7RIClrpYe0o9cJF77AbCe4aOZIm8fAQpi
WnDJS8imiEbc/m4kGGErsp4AfAyTeTZvVxsiUCVlpk23DoP6h1w9Sg96RjgXi/JY
MNg0JVxXMMsAz13J1OxaWXN2VNGibL6IDMRYKyb7t/CFdrMPq6IxplOl8fA5MfiT
CydYIm8QTORa7yCVDL8nUIKiQLo8A4yJy3WsliGyfV30ScJsbIJ3Ob7lieVgmhTJ
N43FlEwJ5/VbvBsYBgb931pL0uQmXiiOFhAKyCAqCfcCTCgdX97d8PVV6k/qYFBg
cZkcEyWrdgt5d4hzFiG/FKTDryfWneuGcllglkulUCFsNQmqgudwLFBJqvWHtuIm
au4PFWBPnGpJjbl9Yp0dh8LhRmFtMK0tGMSuKdfsP1XPpMb+RsUsxpo+0x6zIDg9
wD7JQ0IrYej6tlEPKXMI/bbm3a7XEWXHeytaTDDDvmGSiYTkhIoRxx39gvhXTsh1
a9GdItVmcTSXTYrH/aW89lHRFWIbCr+KBlcDArIbrv8Xjcq8oph7xvK1zqxN7aRm
p9Pkn9XGvV6neRGr/bwC9cBChZ+rl/1jF0UNU/pf5BGXpieHmOAC1UcaBP9D65WF
AplmH6rPLV7Cs8RTTd2MtvCYUzfHSuBpe1LIFsjjcpCt9bxPPnex8T1D2mHKCo1w
EbTROzN+SbWyEFgDVRdZmxfXi0Pr9F/BqRe4WyndVHkI4awTXizewwlnSKWZU8mV
1FsNhZAvwtHPhEwSwMY84lTLdYcCgL08gaWdxVxdv64mTlwP32n+B5U8EHGcK/47
XTwvn/FfMgHF1cGZbAenpw4n3jVxDLjibDPRawIMhL7bK54OwfR6zdPoD2APk+ez
lS+Lswk5K6jKy3nqMF9yUpSZLZOMWbh+3Zpz7MPFmIyDKEX7zNRDRD8s8wTe/4LB
EbsJUR6ZFmbccXfmUFhCg9oBynJOBA+LhCmlqyc0+Hqdw7IRK4jp7dMNflilVHMb
namkFyfcgK6ToCmXlO1SRrgN+DSVYp8lvPaXkNS74sq1yLPAKLhJyFg2GuyovtPa
20laUZ4p4T185B/YlSiRfI0XK+OGqjY6afIsLRdimrNvY6jp3JA1IQEjsjtrtr2P
gwB+MVdBOTICIY0rhjM/IBixpcn7zyi/jBM1VXNHwWUIAc79hBVh2e2+Xwd2TKlm
vOL/zGqCEu9ILIomAyQUp3OredKqi+u31mAgBys7xyfZwLdVgpWxUbrQXl/pMRWY
m+U0dS9B9WJ2Po/7RXXzI3yStIREfM3ghDztIrSD2go0GWCfjM7dgzhTJWGWU2fd
3YX2KZVJPjTScnH6Fqt/QRT5hMYfSwOXqNeybZLcISJ4JUAGkwBChuQtNfUdr9kj
WaTREzpEruKa6ocgrg7SS7d6xHMARFs0Ry4xK9zAI31gMdrPT+6t22Lrt8mjte9D
6oYve1BAcgXpt1Z/5MkAKa7llKu6uPx/Opkit/PDXtTRiqiIaAQmAnWnCKdgGZKQ
cidJc1kV7we0g4YV0SoCGLy8gCoX1HsUSL5A+krPXX03tNwJNjzQ1cIlMTflcra3
4YiQR6oojngJbaTvB73PPS00Zyw5Y5VS737vghKRop3EN5xC6EJL+cAcn46BBzxp
uX15qvNvZCDfbVWSe167mfjfi/mM4xZsZkggofpEbLMwNYYZ/QxzvzBWq9m7qIpE
oghHr9Z0W8ySL1d9pK/rIvVBE4RzRNByiNK9B/jItDHY+a8/KbBrsNxpobEMdXtT
3blkC9lM+4N5GkIRwJUjT/Ae72Rj+QLAgga4u5Z728+TrlzH+XFaHIR/W5RtgOxJ
QEVeNbSNTqCQRDmhp0lSOzkDDSoVkZnJVkIUJHSoE7fkSzvTZ7yZ3kytDQkRdPnK
g3rwWNBRk+4Pb9sGaeqz+3EI/q46rRwWPM+6lNgwdOy/KbglxM2UfhdU+deX71Cu
VG43cU0I0spL9OCwFfl9GxGIYeNu2eyKZrNg+Ol2tx93zYgpTkZ2LZQ+hZ6NiP0u
IWv9+lTI3rqMiN/S2OUmICJvBnyAW4Tx3dp//Zb6+YqZVzZZuQjSgY9PzwPqqlMm
hewpqhetPHWlfZ/PPiyevxGXka0yaZn2T1OqnRvevUq9WfshcD95lo4PLp01zqkm
/9nxs9ktQcmxGJ2EayEvegk2ivClv8803ZdyyrlrVxQEv5UpqwwjLCHViTOFkMoj
Xl8tf/QARVQv9b6cUWgWeCwV2DUlTPDlHTlggmXbl5RPvM0UfDTqGHmkqzhd7Lzn
q1FwE8d4cYZaDzTTLHjEw+ul7VWqCtMB3p2hvv0JvZhvYGASIFjNCmvwcF+F8JuH
KWElfPY3bhsFTXShvVZX3+1hj341ivMzeEplChisM5tnTe7K176upbYmCvrTXcRV
cg72WpZ3AuMp4bTixQrawyXDRQL3DCFsWW+SsP0Uu1ABxNX4PRb2ONtVYUxkH/+3
53EBysA8iWIfDIqX6109XsqYQMyHQQZNtC/ZA9DfJu7QxiyKWZzt2bwDTil2SvKv
5EvYMoeI7fe+wutH78SjdC4uXWuWOUlRMmx3VUs7qFOBOhdZTkihCGT2gWEAJgGw
Aev6S8ClDdytKTL9wa4OE+LGSUKa1zVZ6xpckpD1nlgO40l9NGr9jdhDBi3Kbp/D
b9xIhU1pzNiS1It0gBC8aE+BJs1gD8VRn8GzSS28N42+b68EotUj/a53oamdZ72k
6Fjl3FxZC/gL0GacCfygMe0A5zMIXBc8CvBW7CfCwQwr6ow0pGd2qskXcEU06S+c
n5Cb6TOdvSVgDqdEI+sfDr+v2MzWd0cpNOZGlJF1dYZiO0dlK/uAz8jYxaDRTEVs
p/ANnGu/YXn3f+7rE0T0eToBXIu0PFIt0EKp8jj6RazYTsjRZVwCzIjGjZiicbTp
3c+u446c4pNwpzkep7FfUGMICy017ZJDUyvbkS88keWENthFiZonr0QaW+aINZVb
dYpwhZWAEfxWaVznxJTOOp8eZP60fNq51b33xZbQpu4uzHAgW+CxgtYPCdc2xqEW
Ko/u+XdWBZaMu8fjUuO0RZu3xXVOF2jFseczn9PXw/cEPS5Agan0XCCBc/Fqwn1h
NhGBt7MwYFdmKicLHHpMKFJ5hgFoZttbPShZPeXknTFMj89V4HCXw1urak9Stb7O
RWL778tKtllpkT8wCQ8tPqsnMPujikKjZoWFeVZXKdnAp+6l4QaUUcBUDAhxuUFE
2V+GEMmOTQ/aryOk8yr+zx/6Z9WxKhQ8gTHE4u3gAWooNFNgrKTW0jcqrewLmpHL
o7EjfuvhAhQKIO3der6hHfzKufbRjBUpT4qqFLDwrzp/5cwfDDRAloScSxw2PbS1
GM/aWYJnMuuF643k5iFtWR1n64IKbdW9q60X1+1NBiMz3KYdugMhnYV3hFolMRug
4kengGxnmvT4YK1ZfhHPOwWbqpFisOwvbXl8QUNMC5RFeupHEm7qYn8UUbs9ijYx
xCQUCsfX6MBgcDKKIerD0ejb7OEWbPKHELQ9lemO2AmKRnstDgCek8YcOXXftbQ/
ECJjw1VJTvd9jaFNHSoVGKLgjuCylMsvqMINIS4MVZDMii3YGTBeGSSzIuCVOhDt
Jn+nNfiFlKBOcUnsTCKMlm/EpdnWS/i7yDu2gTApw8iDUx7z8nKsSs2badks1Y20
OTfeXS7OkDmOQocWtlASvzV7HProxq5RpQOsov7BlwbfZmjBRq2yEmh7LiwXfDrO
pgg7yEv1IEQxUFgdynl0O24M+aFEK/MdIgk06TaUOrwGudvG0Db/+gksy9jjFwu9
dnca+oTThCOb/hYvWAfToOVNqxqWVuQ3QEBlsYw0zXGWxf+G2a6eU2vjwGHZkWPA
szHSvqcbgHVNZSAGGoMfYu662txai5b7YChTjW2sLswutYD/5iHrEq83sm3XW9o5
p5daEWKxcyClKcFYJq3sthAh5JemSeguUOX0U/CvG9LeMOXHFi6/qvQBVGo4IMJT
MsWuydvCv3E5a3W1bx7aKy0qYCkaqOikzhrRdmYUhJkLjikITSJ5dSvJkfQMSi35
2FNZvoDMvKNQhTamSFmy3HcxBx6OdvoK1AGRXZUWrZb9ucU6PY+NhPF4zKbcJE44
ouywivnCakBIsEbrww7oYyLUHRRBUEuCPxFQ4LOPdSCDZJ3x6Zcn3E0bsJ3WNRJ1
j2bV9/E6s81z06eukp9h3t8aQIns74uhBLkU+qbpacv4q+CWk5ROzvOibU8uJF4B
vZrMBqFXcPOqTPaODsnTstA9kY3wgXFo2mi5Q3oFSgZjuOQZ5JocHQ+RGy8+Ul23
stWK6j33MywE/8BpiJyGtGJBXsZKFoEGmOUP6ubV8jaaNwVAj8FrlefasUbKiQmA
/lJRobSfAXmHkSN8h5rw91kR0gjWss2nWiAxSAmSsUzLFvSFcAarfqgVJxCF7RyU
cTfyc04ST5yKl9h0dyFgeQGSHcbjjSzOKYG+cVi3Pic0On2oSjT8G0bdyVddQU6k
fGh21W1bxXRfXkVS7gwEPZvwU1RkjoAoh7ccTRBiPAK7opx/DPr/ALm4kbN6VlDX
zL/xFmWP3N8wZJe8l3S2OIO2elLhrLeBw6Dz73m7TxLhpIeZrvxY+5zwogOAaTe8
h6Osn9+1zTyBsRW6WWVjmZSWTpu6SCdjAVnWrnmfGDJTSYo1TmVDqUQIhzySRQpO
558+WLwrpy4eKGcBcMxSVpTYWN+tM1TFLL5F+bX7zfc23Dunqb3xriBwiofb0fXF
9LRN31XgqWZz+SWXHtK4NIeE2RD9q8gRkoTQTyGsr/MTBeg0ZrrXgs3odMOQwrGL
ZQCk5Va6stdJJYoMk/eK2W4MxErcvtDB8lAU8hhcviKNTLE3k6hYsIaJVhdeLmLq
amV+q6awdzLiXbP1fqZ73ew09eSx5mybBnQ37GMLH4IpEUZ0J6kgZbe/JOIb2ukj
rFQ29dul7a9wmSClJYRHmj+LUB07UsIUdNFkTxPSX9vaeaCrmxbNQ+Tf+QX4kGBD
yMv7ixdLjrR8oe7rg19dPTv8dqPo2wtIPBS61fB6pv7SDSHycnMGJG0t3wWCoPjb
scEL6kSusaHHlwzuBPiRFsTJfMLfaxWesE66/MSZPEoFfpF9175X1xiDu+hLBDN9
VEcHPncDjBETVnNGH+w/hYnazApX+QH2TTHALKIza9Hp5/Ljaqx03D8A8iMmDrKR
gChCvB9Hq6l0sKdop0i/pnx4EREM328UUcite5naGHt5GFduxq/OVHMy3QTRn/Lj
MVE+ZCR0X+bX/NGhKZMxgBkEONM3f2cxOqaMlt2iKqTi2iyov0jQQQV8uNbVI4th
/4fnJ9/i+5SvVQo9sbvuQDjPioYlxyuo6QGwaRyY4It7BIDu5SPIkJdJAMESdI4Y
LZWUzKL9lMEOqnebtG8ywVUtRpx+jzNO8wFOOkWiv0k9t/ACfg4iWI0uFuosLKy1
4COzRfgYiOxAnHd5Lz6TwRpv9T4vPZdsYMUSGXUS7y2qo7C5zloO4dHytGZeRHZ9
fBbrasUsmbfhlZFsn9F7BQ7q7LF/awwVkjxRBxK8viB7kqUsS9Obiwj6vkl9jHBz
04uJW1JsaY/RSd7sUFloMapVnfaA/jH9OOQLFsffNyF8bWm/25on0D7H7hGfMyUP
pjRBFfwVz5EGS8qqynQSmC9HY6hoFGR64OaH4fTBD1ofBnoV4JgBNuMjaHWwTLoX
il1N9tWViqP4wnWax+e+mv0Yw3GJZFDQEyQgb9Xd/y+ynaEsVz1bI0xcmCUVg7rB
1zN7dLgDjdUbdOGUMDDC3HaHyMcRNmWCkQBORcCu4++13fLq27JxEz69ly5442Rh
N5EWgK4WAgajaQKaQma2uaGUurQW19evJBT5jhBfy/wN62BV+YGjHfrjOMliKnmp
53KiGB/A1P9aGs58mVI4vX86FJXFo5rKRkp7n1hPDoMUBr0/EPtu07q7GPc5GfrB
he6toYcZld7ehTDBnTP4ZhguvvuuC/3RxGsxDhQXlqjEzQdDdhOTRyQBDvvE/Lun
vlfzJ5UQl9t2ULboyenNnaKMzUgdYxA/WKycM5OZ5gNmyGk0BW/+6U2riEji9KwQ
HvQV4Hlz4ScpW3EZdBP6W9+PLhXHq3SyJA55AFZEkN5qJt/QVY3aE4DEvaXUHzCu
hOVsNtPJlZsZeXmO20O52BR4WRIjni4CbbiOvn/9ZJLurS0QVxor2uFbj/+1efoo
AmomN0peAQ9lw2M6d8MAWO/u1UI3vDBOVfGmWbnK1IAV92IKbVhJ45py0iMv7H1o
zRPWHVNLyMi+XU0gF3zFIn1+7E66e/XYAy+4wffmWJsNNYcTMtegU6OXHCwXUlmq
QXHVN5XVPon8TPJPLr1F0vO+TYW/VrvlTrHeZiqYElzy2gGnVrLRmhvUveentMJx
N3O7VH2z2ieq4DdzV3Sx+rEux+Eg71XUKJXQThVdZuxDMOhOXZVFv81l951O8wKu
tKLCzW4WZpKFme5UbCbuu7o/8B2F17RWhIUAXh8O9BXYe2f6dmAGgaeqYLErOcUB
NIygFUQLMmziIdrCfNO/HPz2uWkSV6K/4QIL593S8wZvd6zBAoXWsG20I2883DCK
ZoMBaKygEHwM63kYp8jUTBCaIYpMcuURReeDSWK3wqouE3Oz9hwTKh7l39Cj4c4P
nqltc2Dq+7qslvTsqMi0/a9JQ2/j5b6W1FTnmVtOVFMWr2POfXTTE2E9GOBe6SID
uZUsxD7oxjxuqkufCAsEZ88ldexivyRn5xOcL78PICnUrtLxs3qPANtpGW0XP53m
M/ZPQowPNGJrhN2iTRrueJILq/dHfqmSw56ndFZIzhxfLM3pMrr5/ciAr4g8kvWb
c7hbJG7/fpBL3xR1GwXCUrI21lkB6wkYvH4MrZE/4YPt6i4bLPl99VS2sEhnVUu7
j63RPr8tTOggYspHEekooPwuTlhPzPK3oYoeTomg3alFTnrJBDKrSTK9V4pmyM6f
Vvdn/B9HHvr4xQ1gbw67t7UJ8h2d+LqsDqowMvUFBq60PhtRMVBn89d9JmOdDpKQ
EW+dWLPv3057C24xS2Uaq9JPjrgXjSVupC9WyqxSlbg3koBtxY1Xgf8rAQXY8O3C
xHkOmAqKhp8+k+y8tmNs4TXM07R7ChQQdwj3oNtpAXqbU1BPsYEyt56DPFGgmDjm
vsJLnOAtkVAoe2ekwpYbWql4RnVTeg5diwaiVFUe9LxktSrE23bNApvaMlLWekEO
j/XDN2HgtU2zmvyZZQF1v1o/tmpTHI+UltDla7xEj/znoAbZtUBCK/5rwa6bHJ2M
COjh68JaIpV/Alfqm6QYA0kayMAZvBFE72gGXkk7npcnOQPppkIY3ePx1DlNoEYu
Td9pK1mqB8J/Psfqxoifqj4+h0AhrIw3r4WAbdEW3eHJGiq+UE93qXKYG/K2SrdH
u+bExUF6tGmj3Ylc0EeNOfuAsdNAo7yZFegE5AlBMNRf/oI4uInKUH0yUXgVtTcA
bQDX2b4iSL4yrMdKqEPYt90ovZOeny5nH+rTyvu6TXOUxVcVooCCACczlMUqpem7
46DrJDXjlNejz6/HFijFHAReaYC8kxjz/UdqwgK0U37YRbvaBF+sw/e2dOhbMVa6
h3zoFvkgIesEnh9aqussZ79CrqDomYuBH2HbJmzMnHfYRVvaEa38kX7CYJ2jvpnf
iWo4TVuShoyyi8yR+c9t4WZ6jMYzU0wjoctl6KcQjUKPRNCEIfuhwTaF8Nc+9nVs
kTXW6DpGQJLcdKIb8Kuqog6ke+a9qq1lBkW/Q5u9fBSKUTCW1dSA/b3HGe8N42JQ
/o8igLlUlkq+IJtm0QI1IBNDcN4vuj1+Ni9U6hLs4gc1nAjJo6hKGnNHdiUdnlva
+t0TSNVQ+WSURreMJCOVEoTRKgXyIfj9dKEZaMcvB6v25EVHDipz4ta0vA7KDYj/
56siq9eGd1vAFip5pWPVLbuiYukmo9P3Bj6HyDDls5KN14CQxnoHUxNNYHHkB5wg
TfZwG46lMiJtWyjwIRt4o+9dU+bCQG9vorU1iSumewnHmkgYltSwBJBrg7wGdwHZ
Ad5WuccO0qUoZaf8dgBLZQW3MmOQvqEQTpuXU0OqKdLWS6KIyoT5HkeYyhtdbQQR
3acsWatCxb0TjZZHG/8WH8IIn0WvQ83WIYgjPVg8va7soAkGBguo+rQCU5CBuH0+
U7Sqoa+b40HEHEFfegU3jBTjhXDLxRb0Ofz3KShRjL97M1OWQnZFkh1cFaKijNX3
+Iogxo55a9KDJ5t1pGi+qhuQbiUCNSLJ1bbbsUr4SLpywxBTocLFguxvstKhi4Uu
swoVguQE4sBVF4Jg2Ky0PbhDUaryY6pzszk7xOupSY+Nl7vRUxETLnUgyo53di9v
SvsU4DTwEI862lKmQDUCZAf3AiooM2jXuV4h6zBW5YLI4Ofg9li0y84I5xYZD1vh
85hh8/JTQ0ntrE7x3I91jkInLJMiwm5IfvkJSXrk0XVpfjzBrME281sS3ldY+u4v
elq2af+upuGc00/QnCIXBa84B/3fQofrYpmhaSN5fEMQ8HwEdUBTZS6Hkm4eaDLs
XxLmyey6SRPjHA290Q6dDcz/+vdl6w3lamOEmWhzogYTbZ/es/+iKsk63HGyCkTv
qZXERJjaQ17OP9e8u8CvViy0RVWwGUbEmXZSF8B9d80uzCdRRMSffwj0V4pHPwyv
oB6RujjXVAy4NnOVza7G8B1QA1GPLBfPXoiW6ErC9XidDLju7MeSfsURJ4a8bcAI
HssUOpQbFI6AEzYY6jnkte6hObblzIgCILLjKBg0SO+EV9aQSi8Sj7rkNx422o9S
o6UdLSwzC+TeWBdKvTXreLJqGp/QTR2xtu62/SELLyLR3bVtyk3LJQ+q53s4Dxc9
oG58l7uaL3TRxP8e+sgXfcW1lWAv5FAc+HKhf2/Mg3tbtR9yeI/36ZYyl+K8NyqI
87q3SLseRFPqZ7vaFAEqfA3VUAc/M519mdhaUjlv3cl4/DKP71zvrwlSjNLS/1Pj
C8dYPSjiauaUW8J9Q0K3zio9YZHFJ/7nC0ft1nZC2e8XWZHAuvZBUUsSv0ErTy52
AM4jj9tooUXhPHLrIorbJFmjKS24FIcwpsTMooLvs384SZI5jorsMV6kKGbR9b9W
tdrDntalUcBEX5Sy4EWolnoysp1YAe34USQyvYAQei1IUsGjHbrPSfHBrp+MM83+
0CHGoprjwmbJ6FWNP5+jdQ7dJAq12kprjiU74L3pYumoBlFvgmMYVWRXtzV40Kgx
Be9TfhDTmnuc688ZB0UqYJKDT2A7zfpTymmtEPkFdphky3iBJyt03qugaCP5X3tP
3sGs7hBev7FCaAgcqh6fpKlp+UrbFsj3SN/7Sg7Cu6r5staYRoQrX0etAplBcHV8
VFhB/K08M9V3n5F1y2ipeuPZXgZGam8/0Nw9VN0TwRXqabbQiWNmqXsDpuiMYfyj
2rR8l7m83GzA1DsN8trx6/wRoxnndljS5t0K+M9L9DcD6R0+1+Tvd2UcZ0XNdAoP
Rz0npgcFKgLPC1+GAd3eTB3AoeEV+ZtM8aPVTQRmmzvHcncIjmbz3TVeOKBwmdOz
sTcSAWICERFNNX2yIOr/xGc3zlw1KMV9S7n3nIuGdNCR2DaKjri1XW1qI69MozBT
t3r2siwvNXqofuvxO3zMB1qGHc0z4/an9S2bTTw1ZKY6dNoOR6L1Uoz8MqEWO4GR
3PVghq0oNZNgfwgEoCzdfv7D0CfE2YACznsw4v6IMoCWGvLUT6+rGyYvSOCK4OGp
6aWhgfRB2WwUlMknhTE0J5yPWMmAX1SZ9yFRpzQ+HQF8eSldeQNIo44DsOdY0G1d
N75GarOkqDLnISOne2WKXlrzbwjCjvR32GgpIDGPkGMzYvW0X1AOHCxYM+xwCpCI
BCMTrKSPX1w1AdiIB2WHbLOPoWXoLAKyCKvHCtgKvDHauglliZPTx1kZ05xG2NDd
7F40rUEWSfabV9ETktj7JzLiAEfN6oTvR1BUa4igcRrzl6cBuuK5TEzBJnr8jX6N
nM5D65DU1Z2BkoFCMNUgz+RaK1HooIb1I1CeMm5MzbaC9Nm55BgKxs+in6U+921X
k/c2FmlGLsVIRMM7JQW1xNtNTUnYTSrcBa6lY+nGZxobH3RUZqapn0vHNAzjJ+5h
Wwp1MW1ElaiGtP0ylRZx/54I6G+8nuN6rOJD7pkpKGmhyJk/UXUVBBu2Y60uEa+q
4Uci/HKwKpVp56FAWWzZdQ0MrVp4Ls1c3eZ4+jVcWIqXU1iz+QlYi/FrwCRIw3Cj
vJEZYgAZdlan5OXCjZKWUWMcMFNyx95BenTUDRpHVGQis4jt2a5oBp2SFYWdLqHN
UXWN8HKA7yo1aBRRPtNNj/TLkjhiEeQXcFSZ8uNfvkP66/KSxy9Dz0wbRBoiklji
ya/6zdbCqoRmAUlif87FOHQ6MoQmNI8VHfE2C4S6DRImDXFKRtHU1IZHLN2dpV+X
ZXFRT21JrOKXHjf4wJUYJbmxxQtLpxcu9JeIxEIil2JKlzYPOzFuWXB6X5nKuzGK
ZAuG74voewLkSYctF8TdXSrdy8k7aLpsQx0nGCefEbfYoZopsTTIfo7nEmuc31+n
6wnY7T7B0nUGgMlgswugpChn93XankSD6nsev5OtMWNN2B6HjON77Ibtf/GcFewr
r7McPUzDJhRLlCy0TUYwYV/Lcg5R7Dl0n7nGuqJCVNpWNMLa8C8hkAVTOvh2kBLW
1sIxapPNb3wZ10hMKl69fyPBuasEJ54vlJBLpy/vhUf7eq8zVVXHmXw5y+l0nJbE
o325A6idAUWBcgOfSx6IpCTVISvviZySOA0WUdPQA2Gb7v7heENz1LpjoyTG14TV
zC6aGhIlSKlJE6rmpnYOe6r5KLWQL0nJV0ikIwUF69YrIYJIKPfljnMoBg2ZPOBq
zf3YW/E0yK7UBdhNMPvmQAkJdyrNs/4hzztQRHN4IU+wU4KVFWtUFoJXwa7d/B/n
2LxK1/c5ZoUcmniyFzQbjOnQ82X2SJWrYwmlpo1kQK7UBrHY/iSRcHDS9g0FoSfn
mpVXhGv0+gVurXmpqWgAnKg6GM5Ed0rW2vpjtucXlRpRS0MjvIwtdJ/hrXGeHaru
pEA0ufRaSyXoNAhp5aBYp7xmEO6kvZxrJMiUVuv3KkYKkzsm+1uGacFgAzBzSloD
Xp1U/SW9DtrFgt+7oOBSCjWse/H5QnJuZF1WrTdItP//jVkH7ojO5dTAvhjOBCC1
FwoHVnW9lcfU8SO+uSj+XK1kLPTG2Yn6le3FNOUZ3NhvIdT1i5DQxRQjJ4UM/8Ba
2gB4KY4A/39NymBG+qshRiq2ImlCAn/8mbcsEKh3SnwNYUrKi/Qkoe68f8fRl0Ta
6Of1YSpavNZVr8wNOQaEZYsaqFN/F9D6X9N7XrJGhdwcuZsyHHsS58N1LQY1lfxi
NxFtlhu6odN4Hca1M9GcVeoaOJxbF3L9AOBCWp36Rl5EgP/iAQ+7ZQPxQWssNUTd
bAL4rQusmdMVf5EDsm06rwNOHEM/wB/E7449lniyEMD1cQS4Fnsaf6O1Yh1rdiSz
DRmrA5WmJzj5npAIpWv+hcHIJem977x6SQeDCWe/WsOb9E7L7E7MiFuMchaEMdBs
BSJIZgkRBLPdiRiUGUKCi/tj5zV8PCotgxQTkTnkguBQwjSX71rXlHBcRoBSi+Q9
KDUgTxAeBwLAyHq9/YRooCsiHXFjfMHW9Z0GVsku7b31sfDl5hWnBOShap6IgU0I
utocY3SQ/utJrE7fZ1xzSUzuSDdvyxAt69Y272hplZB2PEJLDdGkFCtO4J8nzneE
fLndpcbQ37DuKyuJCcKBUmYnDbMGA+zD1k8eGP9xn/8qntK/VFvj8c19+fSKqAsX
LArgT8gqnADdIqdKxAZ4U9Ijm/VEPc1CsujswvZhkl7rGeLL4Fc6S0RII6xcRnea
p2MB7/0XeYKCw6B/9fL4XESuEYifSingzWrNLlBLYwfNcjT3pEpstyYuqagCfqFv
fdUfTJTiaudVzh//3tDHHj6gRaGTuNGuDdfZkT2Mu2U8SNdZ9ll/6cd36MVf9rC1
3muDMLGfsnaUCW8hLWrbSNS0/mVU5vHogfiptxIcLRo6Zaf3lw63fX/AsJUdY9Pk
hatABJ96dfHafWGeUj+qEG9VoSDS/0wu3Nj+ZUEdTLvS7pafr1FK+bNfEw08GrEo
zHxVJITKsGSZDsZRoA5BRUGwsyi7jnZiYFF1zJcZmV/OvQzHdpyTon1fpTQhid5c
Vbf8K8qiwNm6A3WbmzFg814iBuuygjufjr6gl9ajG3ad4T53oK6AgnDOn7HOe2Be
Yzrjy+rOkM+waENc//XYwc6rv5xtY2Qa4UiMh0csBzEY2aFuVH+83li/V4tuH5a3
TGypZ9v8E0ga8xwdPhg5GRI0f5unMAgsd07KR/V4Xn8LXZTuGFfY6sZ8ZkSHC/1G
bqLI96HeqLmyi+9AEWMbKXyEbsCRnLpIRMgOH0L9IPB0Dqn7Y8ys/SxBEPhieB8x
LBhr9ImYQtQwcjALrx6WG5/9nNsD32qdde1PEm2mZ1lJBudddaYPsS9fK5QCa+sy
IQqou7vcrW6mrZdbNEtN+yFNyC5fT8IhfwrJYtQoXoawdArZUeBT9enLlfAM6vO+
gbJ41n4KkkDz6x1SW1blHV6itdQPb82tOCZ9VFRUPKHD90T3Zhf3zOBGhlLirhVY
N5acRoRQ3Mt05Yo+Eg2kSmUem8BqLEEnw/POizrHCbFuKxg+VJ4UmOHMYXtjXZyY
ye+PV/3ngg5vHPGaNfR5uiDj+0LbsJCY0hLeW24la7ecoJbxXT7uJ3rTb2AROUro
K3DUU1e9yvJqos1NzrodPnTaCsN8mbKoSCXC0fKh61KgqNwW7pPI93sIjODCRm8q
TYR7R4l/Y53jMGRCb1xsCBk1aHi34dx+xncFgE+tSVY/5bL6eUIEfI/t6u6cy9Cc
WrX5TbT//z6jmYNM2arL8ARRoUJIweNpcuySfvZiGi8S38YkUSIz9XKcy7Zs800v
22WKKnpxW78oNe8OY4Jn6tqXpjt2+KLOaG20U3jEVbo4Wsfv8nx5LLupKnFqaGi1
sf1lzhN5JXOS75IYbfzlGX5FpTq2U00m8BwzMSPPkFIbADGqGislddN4xr73gwwV
f/0kf4MUMFPM8xGbO455XUQGFt6c7b9Fn0zpjpW+lmwCxEScMPIq55EiyQqqX9uD
+YL2yh6+bR85AFWAGxGzNX7WBelW4lnVppctKWs1oN3JaSTHqZvAcsdUXApR3LNn
Hw9u4xkJg4hO5yTuSb5NAXfk4/N7G2QTwzwXTOKkyvfpx7lo6gpW69Yhy//PoaaW
svFTxSEzQqGS/nM46yKhm2wCYZDUj7x51VcLWjPaZeiV2WWp0IA2Jlde47+4E16H
VU3r2kP7QobxWjR2H/pGTelrKmZ6fTq0XIlUt3iVhjrKFlZGymQA5SONV2bi1TlH
g63wA15uxbLA+bVvtw88+Xfb4gfsTEhq5/MckTy9tl85oDQTz1TpPy3fN4FSaprB
DNQePuA06ezoEtyCSbbCJzCNHm1yiOTqk2GY8StkleH/Pjdm9L39hr/QvREkXvCR
pWirBcGh6eT+1SUEOUBaGADiW5UobH7kbFBSgRad8fyfz65tfjhXD1fVIw4Yxacn
wCvikp7zrzh0wJRUXo8b7MfRn0WSg0A8hMaqt0FKJPaViQwrHtRTwLxkPgLETNEP
bFD7yUcINIcva78PywcKn2XpLPy9qTZSXyNZc0gcXb7VEqEoiSaSVQW0SC+4bGg4
xg+g2oLTksBj0P0qYPjxjscfVHRXi+O88HelJWJ5hMw/MpGqBI1sahTFRlAum11q
HZzlSNw6QwvSCOIY+deg5b5dgsFtmsXZRmkgZhACxrt5WXsZRqpoU2mIf+n5TAKR
VIMtp+OUOLylBIsqesMWQHpyzvTePoQ07TSBB55vlZY/BHVOb2184efiY3by3DcE
feuPoUoOyi9lczfOGe/zwXo51leD0sHeF8irnDAfs0ck+Cb62oTjlbxbbJyqKJjG
zHVQf3arX8iwUByUCoDUOpGPu3pFkYUw8qKCA7mgBCEejwX0TY/QCJpFKekXVxAB
hP0gw09TPqEJTIIOPyjxGQ3J1YCcF3dcAhiiEvIg0MreRiu0W+6lZb+hIh0bc0aJ
mDZs8FHXvFQgy5cCx6mgzRUJvSca3EimE71C0uwXmQ24zYO5zH3sNsLy4f1kDlk6
t1Z0BQZ063u/RnM9B0+aBa+guawYMKYvyrM8EyYT4rxzcOAAXlxFbbo6yYjccdNM
5i2wXbw55ctO/L4WMvobGnHlXgJr3R1QRCQ0WWeD3YAGvJCuFoBI8I/TeScKayOf
tG7+JGOLJd6cYmJFiUUKWqivJASojVhA5TnJtWKqCbCDD57rp5wNzChQBbMQ8trc
WRYrnA3+YLcnjxJkDD8Rk828cww7EyZZPQWAA4vl/bHULxMXlqoNB+ChCf7kTWdU
jHXhaOLopqiKjiPHPCjfmNIM8osam6GmOGH+rZRJysE/izZreLk+QfSToKDgcwas
b9fNVlpIj5zL38U6VzOxC2ZrptR3I3LQcHgWDFNLJNtSWmzkb0+h1+kYIMPbv4oz
tfcTOPNb+PZ8+ZsAuuPICSiOAjgFtc671HE9zD6IhBe12M2uDoM9Swwx/NKdQ/21
cGdHXM+ZJGwcA5cL2I9ln+2mciqUVc4hKeCdU0O9CJqoL9CzulA9bYTGdmy/y952
QcsdVvkuUDdJy/1t40KBpVL+8gGDqielgqsfjEAxBZvjTKHXdPDV+RIDoXHDeFto
ddCJpx2kwnh+KFuoOopy2PuLfuUSxd3h8ZM01MnfceAuBXzgBpQg7tzz36aAWhAk
DEQq+RJdHzHiexcO65dqZSj0qXJD5dCZ0QELcgkK8sL4+3LZHyNGqtinauqGviE/
hgVXMJAmIrQeXhR5yJggtzX2qmKY3Cg701cILQqF5urbuy18Qu0hXKd7M/JxEK61
l74OpDsxyslkuazTgRqFq+M6rW7ISClTjhkVdhAKFINDlzoQjqbDpFwWUlYXgnnh
LOXkdYo2XE/fjkyfV/e5PY9PM9ljxbw7NF2s3sI84HZgDh31RrD5xYVL1Nf87Nh9
sxKMgDPhhSpcBqJ9yydldeTWR7pFXSSXNPk4AuSs1BrsJKNa+ctdI/VoTMDuKbq6
ZY6O1acmiquQ32RYwq2PFM1Y01+GQKJlj6+udQDWanoIGeUL59OJXonv6blKruga
stOETyEgY1vDXFI2QRNklpfnQ7O+eQ6SN9PsZG6M0emn92qQVBl+1Wa8Xrw9RZDY
ONgruXDfZN8dBME8PqgZtPdPyQZ4ERxidbnLbrQenkCmQg8m8qWFysaPp5lpho5V
gFXp8jaIevVe7VcBQQReeS4VPCZ6Hy1JDGHkmdZYxMdjknX7XmApNMTNOWz4bpAl
7w+MD9738xEWF0swFbbU3Xm2Ja4HqsOaIEUo4QFRH+UxG5Jky1oZzccbsf3JVFKo
hrTlRb5mYRRP+yNeyLKPj6HrLkCBlWaIhKnv95TrjfWYw/qJ6DQF1/IKgFKhvFs3
EenqOiZ9WwyBkSmEhcoZrAeqyKp5980C/0hBB/Maj3QMnVpche5CzynHAiUFQPfE
lNIKcuQvHP8mlbexM3wEPKkGGwqT6JgR8AhPdv7G5Zvd6bUg9jLB146J9NYi1dne
328dsdyJKg18EDLRTkWhJtHvYo+xjPLGatt71naS0//qV2dEvp9qE/dhgy3K7MOJ
jGX+jhpTm18Awng4YkLSNhy39mIAD5zeFlZRBJCX0d5ndoWVDKWsjfBsJ9nh6QPO
oI5pRfm+D8q+dcBxJaeWx4DwwRHAFUix1bxJb7V0kfsTgAlSzzLQwcg5Sl2nyw5Q
tCOC0mHLOwjlw2P30199/gUK4PesOe7Tm3BUbw46YrCdPpx8+eNrqzm0Z2ff7z9G
j4Kf6+a4jKCTFaeC7OemjQZO2dHHa2JxQMeYOISWIEqnb+AkZ2qI2aDkvMMrwUaX
CpOXL7WE8MKw31vZGzUlcS//v15oSbr5GlGwI3z+Xo+jBuJ2eQSlWPT1Gc18XpVO
3QaKzNYyirUw0Gr/G5fDPUDJ7o0ultrSlswlaeAJU4hp3+oTZwugR41nnmsHyb46
ZqkmhVQeVxsCVkB0hx3B/83HKXJHvZaogvwM3GYEi3sOFkehC8LnVO/mvDysihcA
NG5/mwx3czvbE07tOjftz3zAxbpu7ALqBZIV3YRwiLuK3ajARSCag9r+ILl2gn7n
TjS6yE4/gTdPPNiqwlwrMAGlvW4zNsZiXPUjgcrIFYDmiKoCMVRQwFmcPMfEkg4x
jUTzEciwyheBpE9QIfv4eg1BkoQu/J6kLPSMbX/rbln4bO1KQ/BsvjZYXOfv/ouU
+4NBZXXWrl+PTSE/Ka377GbS/fpBXqDZkLnlSiuVQOLEeRaD0XEAIssZgJc8E1rr
SmnEDOSEIhQz2HxV3ZTyD7iEJ5e2MD8uItXx8y99y/jkQEeNIZAstg79PEpd1T06
gox1eT59vDaQ6gGP8x4duOoesPFYy2c8qUk//DzMcHoPhCkXzzwzF6gnOxYZx6l/
DR7c8pBu332yIKITd4tmGCpvp26MBJ1iIhYnByt6jR/ejZovrHw69Sh0wbf2hhh8
stFz5dtvRMoLIRmPptBVPqSYuO8TGe8mHr9fn+TW1q9wdCQGXTmA9zjpC/RKLY+3
vrQgsIKS/82ytP2N/5+3x43f1muLQ68SoT3aTnjmA8eebWsj+BPVn2P9af4G2CfL
c5Mz5YWki50uU3MKM364CwrIGeSbA3tBfyFc57ErTW1lPLTP6bq/mbLh2vO15GGL
B+XJ3NoNyIHf0IflHq0Z5Y7RlVWLFS/3K6WzrBGRwcLIbVO7kbiAdZLXw63tEdGT
0z3ZocUyEhzfP5YjePrvHjdv8+kgdgwPuwq99KZdfTGIkS0TCQwvDizPEGkYUjvj
VZECWphNs4tXhnXhgC518Oaugs5d9j/5bzP2xJML9k23lUvxoWk5aywS2qTikGCj
fL7bcwCJfRfOIAMMNjer6JVuVJHiNvFIa4Dzhy21lnHjrB3sQZuLwZvxm1/Q4UlW
9JNpKBNYLKFsDQ+iut/27z4g+w5u4DhDbr32aBj+LNk9CsXG2GjlPmxoub4mQ0ix
BzFm22rdC8XpHH2mF+npNIMbuozkDbbOpRyeV9Or/6RUKg2THT+7xXbiBgJQQecp
yQ8Fe9BOkMDY73rObTioqwN1FIO6vIn4J5QePYUyqwDs9/ApVZ9JstiJiE+/MnZn
NLutDQLzH8nO9V+WxdlVgXpmQ8yHiv9yuAxUdt6V/DfiHJ0X3njPm+wl6VuuHQtg
zFR3DcR+NfGQ2bZFDFRQ5QR/kEdXtrSjPks/gwKB5cz88f4Aauu9qwbZ/rRRBlX/
FFIDDN8cNOjb38EVuwLd0WmRK69bd+gb+LvAp+XFVryOt2ykM0qZKBtIqOgwRXfS
kgWY4H2QizqIc5/yS99hgZUHRaWyBW3DFhJOc59SJyR3sSd+LkTVPFxQTLKzkmzZ
jaRuvWnHsopFZK4s8c/fXPgwvQ8Y5F82h3rcjTM+rjbAS6BXW94Afvm1p2aAKA2r
QOP7jALsxwirWFgaAX9ahnE+OahUNxuR2ygw19iszZyfDVPlTh6RrgXL0BD2/U31
8BnAcKP7WqOpikyDCspkU9KiLLxurKy/Sfx69jHysq+hBKgYdBTfN89Sj2HX+mrV
8xAbRK7yWbwdy6cUf0QV+SOG7u8t/L2a7AHmvFBX/8xxL5Tk8DZFuzgCZZsstjCi
l/vn9QYhp1nYqHFIWMSwTh9Y77394wOUEBUavaQjAehJeQD8VIC4Kb+9nmHeFbz+
mwU4eo94OabB9zqIiUWz5CctcjTEcWEr8nvJrz40pQyoHT07mHHp40vehmeoSjKG
4ith82R+6goU7/wCRr4Xr4/fXQj9vQKX/XxinFyEAbQqk0rpEuDvgCHz/6Wdh/8l
RtEH7nrWHVI6oKkXHBAhaSu8sYpcY566FQFpluhfblvpLp+l9SrIiBAZ08cKqqwm
W3fN2CpxZvJrrF1L2CFI7JYLDokerDa4X6h1npoMcfP8H4DDcIsLesJhKpDlFnJo
DSWATRh98pI06bH2oam06Ltl/80z4iDmpyDrRmuCXSD/LcL3ocdYpMVMn4OB55/1
xby7vO2EX2y4TtfPBwJG1m9G9xs7gG3ZT5lQjpwitcITMiH2d/l2zNjaLnhkxq0o
ypuoIQ7VH0f58HdWGLyg2+DitqB3ZSFBCO87egxJUbhQUXRO1Cyugsi0/NYhcbf2
i+2Q8fMVYE4Xj3ZuSINesAo5W4C00jANxiepPSVb99G+glbm5xOTG/xZZibp4d5Q
8//p724EnLGpOm38NDq29i17Fab9/fw7crfXqHGfBPVfQx2jlfzecyYc+0mokN86
cwJrEDqmv5UdeS4e3Ym6l7pfl/LgjnnBCLVzth/xcTGDc7jA85pvFWXQdsLw5FR/
2oNsMj1p3UHIBuH8sFUeAsPMVpsO/J0uIL+DDV2yM0vLaVGc0pAkBxAZ27crP8vX
UPYQKx+gzO9ueM/kVESz3+0BbBx0Q424Hgqj63gj3DfRY/tIqt9XXxd2mF4dtf5z
d1fYNaUMSZky9fP9BxNmiZCRBxZzDn7fU4Vf+NKPAzmEhOL2E50vLq5VR6qJSfFa
61brqXNlSElWBRkz0CQM3lKsY/xGr/aGkqyxj8hyj7cSvUh7RYLAtDrmOsPDvAXG
/BdWWEsRO9kkVv9P8NoWIUQe7uIT8TrtwlLm4tfJIwMBiWBqPspjnUBhK9FWW0e4
wi4ugYpMS81vUpMjJGzznUu4LWnzAwyk2zq8oc8fV931thNLSHwBXEs+nR0/UyjE
B6VzSgRz5/zFqwapvn95wkr4y5QZu66jlAEIxXYtk66BM4SJTxhvO/aK4Ok/1IQ4
Q3xBqXzvLYCkex41SNsvWFi+1PS1iiyhv2AcLPhqDckGPDObChY2SD3Dv+uAkste
5TlEtq/60WQC9zDknVQqZM/TG2RlfCT7nXQ81TmDl7hh/mSr+HBNPeZOLPnTnARD
OuALsrgpzlIPIX4BombRXily1JVP0vu6jA2jZluxYN+sQNPHePMPW6lYtFHoscUL
XjcaEABLKTtHhK02ZE3+X9AxYRe1OTxGNC3Jc2teGAkqK84J88AF6YKFhCPhfCNR
2n9NebtloEJT55xITx3lJayKD+ZQojG28hu1lmKN50HcWJzCcNVArWL+SO69uly/
N7QoW58CMWwT+b7PWzKxZA+qlRu2Kf2Pg1uyIH+FUpXpp/bjr6Y1bE5ppYjcsc/J
6cDAKpDnMplVxkaSS3r7o6MHE0NsPsD2FGQcCH++cXCRmMHxr7OTr7IGBWGOWiK4
qVck8dnOQjxLxBOnrqRQlhGJsmepdh7EapqNWsUSTdNISEDuSSG27/2rMAWU+EWH
upOWNz+nFnyxo3otFzvMNSzYJPyjz1SMnX7ymvtbgiAa6ye8zeLHYBjbsGqJUpPS
2UWTftNYA8bQSbETsSniHCnup6v/MXVzFkXdj2HEH9TOagioBPDTlJ/+glwor0Be
ekE5EqxH3rvBrDBedRQtJqDb4hrxj05Ui/JoU4Asj0uo/Q7XAb4TqJFCKo6VnLDM
b036lfCaUjPLP18dbIW1IU7YQ4yURJngDK/aHjY+WknQRiD54WWA1l4AUBNKJCsQ
vi2BRPzei+EgMKhkXAiYbM9LCoJtn4jpcps0a+d49ow2yj3jLEv+iV3DhR0YwUos
NuVe1morqPgAx5XUwnzbqoR0VNrnT5eJsqIu1QRO/LpMwpkSqAXGBCZWZwF7V02k
v+pHsei92W/L05+xHxbP5OkXwQ76HxcVdx4oIExVcMkH8Bv5w5nwk9Th7ZMrTBeC
jJtC2h9J41FEZSHK8fXVlXhQ8F4USRDUgM6PPCmJjZ26Pmf/AMZA6aep1BD4rxS1
wXd/1yHqhiFj3yBZZ7gdLvEsfsmukuuXo22hcVmVifAW9l1VDirXDSygfgU6keYw
PWxIgAod2RZaXMH+LyJMWVDmotkz/IbMlo2xvMEJDOSY2kmTAHJecCBTBArADc1Q
ky8/7dCml+31iNojhOmBzd/MjDi67cG1sbVoBMkTCC04cYrdVznpjCZltYeJsAy8
lb3ZIWaVKQmLgD+7ExLSG8Uf4ZrVpXsOjwqqN3ya8za/eoCds5Mk1k1/dt+MEopP
E4O8pFA7ITlVCKziAlDcShLj1JtexCQleY6dAmHqAn23RaohFcZ48gZQrls9TwV4
tikMi/yJjpdUXJ6rwZc94AjZdia1xlpIznAFhrnEwHOb5O3PUIIY+KIqNRhoIlVZ
D9pJpDFXxSW4f2GtAehzpEQazvipRXnwyGXGSJBBq2OOLpqtuap2EvUU4DU4QG/w
SMG/P1tAJXdjl4RSAJGGHD4pCHaG8hGeVjnU6/uS02QgjGSHEGsMaCurVPklnTUN
zT8GZWMAgf7MJt9fJuZpkbKfHwEgs2fn5S8lRA2tG8BVj5BL/nKO5FqvnhdXi5zc
gLGFlY0UMKMtMo13WFVAOnOnDX1IOYp8SSZgVp2Eahm19H9y2lBLYdI4fZBzdkgP
9pdT3nfV/7nQ3mIWBtLFmj3CYkn16RpK9yWDNIuvSh2lzicxsWGD1/DwA4gfQE+H
z2Ss67DOBDdZ4o7TZ0ghO24m5s8Qe1ecfqFvQ7Y1kVbPEdVqxln1V/NJcJVhRBIf
mDDM73kF8MnzrwuRvtPvPxSRikuTRVcxFQmgMHLGMYm+0+L8wxBdbkLPxYN+4ZzG
WhCwaIrEXsn4QNX1hvbUef17WEzdQdjZGSCVkCPIJSLymnrr/4OeYCUgUFUbo/pV
8CwDTaAZPaez+MGQxYQLUBetgkKqJJa486G1tX2wv33T9CFPwXrVAvmxS37L5etf
A/xNkvUBPCfICZKsrcJcIQ1nl3Q18mdBwXGfDJzy7pMFCbEoUymIF6qyXfT/CpZH
p+ce2xVu9UF88fv6lL50YytoFYcb4KgWrLtfqaHOjNHyCiI4b+XlA/P3GdkRyApu
+GipFfwjCojqg+ct1BtNUcw2A+ATG5GFW+nXFBPV7qjr/whMztEdhi98neKVnh0X
p7nBgvYQybNH6//FEhRzPIOmiPf7PnLe84RuDgGPQo2AAKIwR0rFuGvHQNcGQzG/
Z56/buoMibaxsJoCHJBBODxmAgJQVN6snt8Kh+5ZWzEVa0tI7T3W0XhHqOlzFXLH
OvFD5mB7SNE8+hJwSEQbrGVDcfDY59vsA49dRlAM3rGl1hGituo8eLMKOQzgJqtk
hIV+63urVvkmjponwbSf1Rx6m1VDIFP8+7jpQ3ZI6FvW58DjFScur+R4OzW7DY8h
apfF3R3SA0PIhDccyHdf2/rROb4xYAuqS2+tDDVnkFWa9CDtN9XtHoUiBWP5HAxJ
5YPWod/kIPDwoezaGEVB3hGWlXGd/LppT+KCRGKFXATaoz4FzT+MdNqUghqIfd72
mc/p+pmXYwHwwAxl+s8L7uLMc+DxiU6iWRW4bBKhylRlJ8A0FYOuaJWOoBZVB6xc
qgraLvMITC6WKA38srPY6BJKHlyF4Ouxms7APiNKrNce6xmepcYlusmj6jieFgiS
QaG5CzE74iXnQt3PgXvW8qV5moE7iohk+O19DbNK+iIU+ph/Fh8LbF/ZCqu2Kkwq
V88qUR7skURt5Div1711Kyz18xmN3Q7vvqRQX7rdxybXtdk263Cp90FWNzlDSKWh
KWkg9LlcW/vHHvFhhEIf2UzanzlGW7hlorcU1ArPAFkJuWfbQHuND51smiF4i0en
GHgVGMPRb6hDbiMaswJGljpwEXVzXx+akY/C/JkiqkcanmwPhmWKIQAxyn4G3v9X
eoEZNomiStMkWOlL1WbvhsWslp+aWxMGG5jMCYbWzVuHjtyMKJDqZ8CyRDaFDvRC
RKe65GVGxtqTBZ0YNRQEM3A/NXkdFmsrbWvQQqGzp74s/B01brHMqXaIUbumSFeq
LO97tcCTI0SxQHio/Z9JP7xIolB6n8d7/sDFbvDHe3gYhy/irv/t5ShXgAdN2aS8
F75fFYffRk4+dl94J9qf2sMbGsXXIuvlrqy4XnFOskV2NtnMqshTqm67AVlMuhuv
hsaid48ze5hXa47VKpP7lTwz2/U7IZ19hqXVn+kih/XLLju0KYRuDqbu22+uHoA9
6lL3GGxlDgs90MbqoBSikJNfOf3W21W9W8Zxzkg4IxL1r6tuWKtAp6KZzd3ZCm6u
kXB2VB47hUYusecswfNM+BHfkJIn4bSPrhhBBD2gB4GOUWVAtmedR2/BXTdRCHhc
x3v29d6B/Ofjj11AJTTsTIZlB7Uj6/1NibEWtD31yAmtXWunyrTjCKeWxiCIBxVi
q2rlW1I8/qaSNjX7/g8BO+2MtSXtn6Go3sdUW1cFTfMWxMxRnwSu0yu/5ZQA7dSk
3arG4+ic3NEFEV7p13UTWTs0pXxzPUWOQWCgpB6fvZWpWgJrwpTnm6gEEh2au0Xw
S87E2+3EZrWqb8kI7Yz2TIW2ZNozcPUxCvgnweQNos0ODFkXp2+8Rs1l/hKHVmjI
FPuyP1Tjmt0GHU9QXCHM7Qhd2+/ubCKrvHrS6b41u03EflyO4fQSqabDVYoSfY2D
sFftY1aD+sCmBvECAMx+fBh+0udRFUw6WryuPJrJcIKBSkWfIiFuMMfUjTT6MI/f
wFnr2eRcj459e+s+EZQs4B5UkeRunGlu7NL/wWu+Wonf3E16fdcHjmcE/qY/24EJ
hYps8HLcc9mvJuT0tO3RgGpgZpVVAXSH3efmJZUGqoUB5XZP2Lt+3PrOvc+5GntM
/8U7XXsUziUxvjhYmBo3f0PIDGk2RhSEtZHW4oMMTXxqVBTwfsPSdpXB9onE8OKV
B4Rlnorb3FUI00byjJFlfgrAvQgMnNUBJBIn6fKpwbbJSAC/d3XtU8Ph9ULpjF9e
4r+7TMZwreR/MSW86MOantc+q8YHkYttt8DN+Pd12a/VLeHJN8VOvbb0KA/djva/
W/rmZYUJaXeGjEpX4fQQYw0zYdq11nduyZc1XKH+AXu7bEvxTbBsSjy42hCkH4mS
wCnofag16VKr7UIa/4dqhDocVJ26ZNt4Nk4dBnn4F2aYoX1RDUBRNMkJogOVcAL5
Y3FWGDT24NsS6XGZEc1ihGXF81Oewh2A2JZL3EA19r0TdVLxyv/WgvKyqOD+RWBL
8shuoH7XD9x3nRm0ynDaFRk7rYLxBAoe+U0U/DyCvQlS1YasMg+jWqR8uQrUdzQP
mz5OoGxc2YoJZgiGb1j5eC2QSVuXR5QUnnYPSPIZA4luhKCIpTkjXJpcCiitteCf
+SM9lT3FB1A38YZwibKrdAefyZQWEEpro7J8uZgqONp1v84R+ePbLjAzZhoInLDw
VpdDc2R9WI4fJu9303vKDuGm12K4185rvWkLu7MRYzI00pc1OdkJ5h4TGNOZ5nUx
UfQ43Mp7KRsZ1tXNrNs9T3NTmT4GU8olI8tYvmb4k/00MOzT0O60nF9JOuSmal+I
5kxGNCz+WratMa8n92+riCInI3d0IYRu5OSsS4ifxeurz1gTQaXoGpGB/NFOBUJB
VFFj2LfPyi6Q7RfV15n1Bgks1aNsrUI9ciaXjRFxBSb0fq8bVBApIJ5gyLisPgYq
NhAhIckBNRokS69pBSHLd2XGuGJe3A6zneYubzAtb5V7NvAm7pO65echYm3qEbVF
1lxwvqMSFrw7IqcheWhn3cDXF7aijWkFdtBO9zim5c+GkognInqgoCCCjCtDg9h+
ipL0dZSR/RGsfsaiRwvmeRBwQyuXtUbNFTW74bu4ifGnXG0MRcG3MJbGXH5bBzeY
Xk42pIB1EJZH8CuO7hjKEMytK26TwjgO0SQsd1x9jdefMNUD4veQTNwxJa6Y5AH3
G+fRsW9ZqEAg8rEnyW8BuTY345t63pSJLp10b2Mf7bmcaySc/4cFgFW3SBzMro5N
iXr0/kU4ctrtWy20h7I4ToSH0UYYWtG4UEx4yCUB5kRnUWoV/ux8YthGETPcs5+d
H23BPU3ZdXDbgQdJ2j89J/HoJc6sOqboVdOoOGUEl89rLelPQgFyKjhvNp9B9lTD
Jyo5//CnyPNtYfqUMnVrAmbCzp2yy9pGBit7cinRp8hGkce0gNUwa8BoTqfUVCa+
y3eLsce1k5fOQmcxRavG15uuGfXXNWXFt+7jYe6ibNwzZKXaDD29LRLAKfw68uxc
b0Ky7hAQphiYHMocsCD158nNJUrodXY/LsPWo2C5QrUODmWfHqzKCQp56e8uP4zo
s/mT/j9d/HQpXlKgaa5Koa5Fafo+mV70IN9l3xyh/kOtToXe1Atb8/VDkGIJBZhw
NyHhLECH5yLaO3nk40eNpup+kFhDrSbTw0jxA7PqvYfp7lSNwxOL7qwS43vIze1W
nUPpRilFFjhmOZw0bDiS06OQjlXnKy3E1XqMmrBu/AS4pvAvk2sfQhI23vdwCVqd
ZnXTuQYs8IYQe7M/kdlZ2Q24JaDLHEZRTBh5ass28H3G379lDcE/llm/SWAr0p9m
jMQOu4+uZhlYSXCs0J8bEOzN2tqsg0aFQuaRIIJpR/JIuGHoOS/gQKusWwe6wDgQ
e3tgq5xxtVVBav3vHFXTjVIxmbkfkzQoAyG2ldvy9ZoptG0HEADIjFxY643kFBu+
mtXStRBW0AuOhES55AZqEKGfcEPYF/bfNSkGhHMRalaynEGS3FQpIDLC8CpgjaPX
bTTlHJKfSrlMWyEOrCKQutQ7W79zSywJLiU5vrEWr/vuxe+VKrD99V1ztOTraw9A
j0kJwaLE5dC7FPlOZw2vb5KiYG49crr6gDSZGK7noKzRMCdf9lrlZmMUly3cryfl
+TiPYD/0EYJUFdE7jOuq8ZezkQPkjdphH0DMV/vqw6O1CbwIdmAdqF8kb3yfdA7M
FrJthhhoL/b7oahtOYfsgogLWwH8GTvomZsH6H2d3cmMFOn8EfQjmnSsOf2FmxEz
2b45n2Yp0r7AvNnSWUvFgWAxUhIvF4NY03fJq7wdIbuCh2cLB5p1u4N8Bgp7sRJA
CJ3IDA6TnVLUkhWL8ryW/wR9i/5clWULBD8NQWul+tVEudWun8Sdg7yE7tSK/WGp
V8sf3vrZ1zoK5kVaQjFfkIxImttqVdmODsUL0CjJL3K3EkWmwaII6ze1ozbJGtoB
btHz4HMRUBkLglMfCtXq85f5uLFg3lTd/ZaHGX/yXrNoCh0+WcaDdfB7BrLQVMta
dJ9NLd+zgR20iiEnngO4PDFxU59IEcv0x0mliMtG1pM5mDiSvgaJQJNPJLkiHpQI
flVGkWZ80GIzQlEv4Wef8X/WRLW4QBJozdIqRnrqo9N7LI6slArL0bCYYim6o2M4
JVE9sepkCjdkBdajrDkfEYWvvXkOx76pCYKE/b3qhrSo3X7iwMF4R+5pXRYtj1Qm
/no3lXajteFWz3fkX8PH+cck0o4Z4dG4aVVufNjKrpNu40yG4QNlHSbw5ztyIFzE
keZQ6dzS42jCfjouOaDhZL0fmal4qGzO995Yq54QMS1Yz3QY8TSkul4NSasmxDrr
jxtSkNv0ke8n0mDXGrlB76RK7JoxsEF/Smd11+jtUeNL/A9m7GLwpAMdKARq4JxN
1wofYA70JHqvgC7UO39zOBWhgF/gSjYee33YN72UK/8JwCx2vyI4g0Jt1VyJbuyd
xlGGPel/eb1dbxRKLxRKCjMFHszhrdHqLvnH11Q9ePDf8usoQMdkLOrzO8xh6xzx
MbEQc/bzSzptFiaYjWIb4jmAdANLtADl66i1SUhm9BO1UQK3XH46Pz8UimDxVsfI
FiVXzt7W2KrzH4QxvezWAg8i0OkPtNu+7CODRHpAUS2eVu1wYs+ULm/J5r6qtlBz
213gKgIcq5kmY7VXJmtTeI92nBVhu4yyBnHonCqKqgiFwiKYzcSgcNG92cazrgzP
z16z2B+RZ7xkyTmzPPlj5XpCuJk4W46RXRzqBa5WYQP4wBOLJ4/ryeMHLpENMp2U
TMsI3WIz55NBau5RI0LPjkNuRMpNLie7K0eq0k1OsiSEkPstDrlm/rw6ihmgfoZ1
79wPzdfWOhUVibeUl3bCF9KyH+i0+mcZ/0Kvs9nY9UmGUNlRXbilZHHc3c9xaT0r
t5XtzgLc9Q+eL8kekhqJcACKZpSzelkJZm+rCySTjVJtZx+9jnLh1YydfEkde5d5
55H7d6gGj9lsxR6pPaauAyx+i851tkPoAvMEROfdARibcS067iyP8HtChAPw/Ii+
KgJ61wkfwmm5xtDoAMw+y6Et9APhKNtg4xCW/wqVPuJn+a/kweqZYis8w1kWuYuh
xmREjJJmJRbYUrYNd0WyEDigjX1uA86tPSA5ZMkd2jbVa6xz4LY9DNcC77TrBwJ9
LZmsLXil6kshHnpecBICcENsDIkdaVhXu71vIWGC04dR+kCMz7Aeb61IMIPbcNCw
tDxfTWzqgJL1aOvVp9JhBYe7seX7KXmPlXx/m3LtEdvllV0j5gAgjA57Vq/EJvT7
W6/RQdjVztsVDtc0eMi+0t8N2ACoCZEz+9SVkAg3N4ATRUCJOnU+GJwkMbJBiUfu
dD3c4siJr5dGXwfUndWsSCTlzyUClFaJzs4VC1O3WBI/PqdVBUfJZMXgY8EvFMs0
svFtC2MrobQ7n7VT9QEwBKnhwuYg4xe4QpVPkMR4hCbZitE6kOkty2tBrAPssW6p
YWPgBP8GwTQIqDYOZlC5UW2dwiOpSqx5diKNgKRSRTxtN8MlZlvvrj6MScPAapQK
Aw45W00XCZv9qOQ3pXS3GPDjRSygjatBQu/yR4wPD+Lwz+R7yy1trD1X0KDRsAWL
CT9CAKTDqvahQCSPgLSKtZetxZjs++H73Ao3oLFcJM9Xs4q8+dRIE3u2rVP1jTZY
+61SDR5VccmXB9dnxibF0yn0z2fV/PAzkyueqdCcp89fPJYumhLjqWJIi846ea1I
Cvua96NGYWOfJY6dFL3HIVSC9P2XN2xqRsWa2QgdInr+0ZH8wvOV5lFk0ntps6pZ
Pd7oykzwxZ4RUF4iwb54K/BD9NegAttHj4sIuR7cAalalxYttNZZsdx0GXGXN++3
LtkZayORl/q7t6wnnXN6+W6VXSJGjh+MWH1YkygYRFxVQcRG62SxMTQ7J2d9R8qG
SWZJX1b3Z1myIA3gd0kK6KUV4wGnpzJaJQIkScq38j/XpYrag4dke3jZUdY1kgqT
jPOW/1tiSkKJ8U7uG7zBX0FZvkfiLZFMLwyzd8k5kTbSbrRRWaDzIBkSvgn0z8lp
p/OK5SLgVdljwKz+MZf4e2wvPLHHXy6fvQybZ71s9jYTYS6ajsYLJjYLLkzK0J/A
ftnqHuzh0yuUCAs+NwGD8c8wgWWZFxTzgrWE/dq+6lMWxTCkEYjsEQY2Am2LiloQ
hY7/3s8kT/KmXbHogrUMycb4V/bencS9zJgC+xPpaRkBYEM+XvptuyPKh/RaoD33
pUe8TNBymGN/F+aa+txg6yuevZDU9Rr2ViD2OockKOAuLA7SIVujAgsweLaSU7V3
rXrC2rsLwv9aEqR5vx6JZHtnLOEYPvYQObeZ5sxNfFar9nECvmxjGghshusbHclY
IBxrDcnZvpBbH/wUAeNBbaQnOgp+o0qKcEK2zDf8VqG9iLYXXsBT3z269k8SQsC9
97vyxON983o+PV4l6JHKbHDnIaIptuCtZknmmPwtNm4MMBLUXSy6Hr3C0FFhn8iq
bnVjzbX1NNhAn3Glm7NJqf2cbTI45wQy1y1WOURpUgS7PoU0ZQM0dn7zg/1qvjbY
bbG3PHxpP5I1X17TZsgotnMv5j1dKXfl4JBLm7+wrsSVPBCQpmkPDOnJwvcLvZNK
jPkQ9CVKW4CQUoMxlfWHMOhAk25/5t24an1K8uECBgylFby9r83lXnzBCsfLXNpe
U+wvCis8TtDbXjzoaai9Z4ASygOlEcnRdo9+8f+TSBdQlozm63n3E/0QReDK0p0a
C2Ly+c+uqQK0/BfZ4C6h4xsaRbTDD/GqlliqpNcHF9abP9YlL7JeX8SZzCbZomsa
T/Epew5+Xbda4cLxNg857eoum/61WFgxYxuducV6MN69Sr9dkqe/hRM43x8l7CKF
KaCdJfJOCEXtICy8T3QO75nPhL7iMtBgsnllJkBFT+VcqSOqgP8Om/z6YFOu6uPx
9mcUjo91AwWdCBE7ifuiaPxoiS99iUQaZ+8o50R5ndZd55t51ZkpESleEusG27gU
xSNCFEpSRLb89M/suklKz1jDYy+wILRFE/Vy3H28HO3WC+sc7D1+Ep+XSzQrjZ8c
Rf26fUtdtljLyQzTj8e5lZ4lNMkEbmagUlAnPYEui3vggiv0A3R2OJpn2/UgnoZ1
d/Z4r6L0vV/Er84nwXY5MVsXaG9FYy+nLxAla6go9nilZTkOqBIrm3xYNacebZMj
JVsMZTTZ48jaiCWrb9wLcNOu/+UkuvqzNgLDG1TnzomZJ8Alw9JB998lprPYf/mn
Daz4YPl0NN1VCFK82E2FdweFxkx3dg+cJzEx30pakVeQ2hK4JwQEZddU85p0Mqzx
2M13DPToDTc06awuFtL4CbyBd33gQJF9fugIoOQw1kS/A/wwJpE+tnwBYBvZD8Ql
Va0BhxcPaKf6834HVqtNlqbW+LqDpEpWQNuq4yW+s/In+5Fhft/a5w5L0he0Ift4
+ix61MXu3dxxajRpwKTG5L7LGEInqIEamWuvpWt+IO+VgxzSsy7xZdzJB2RBFUnY
uDOJfO49VuPURnv0FUqoBGYrfDsmnil/5y/T8a/2ZUNR3VCTTceZvQ2DqUJA8ctc
NiKk56jsAIZ0MlAJc1s65OoUuZFIYbHeoR1IwdlhxSOkwqAdCYLkeXFOJ4jHEKQF
zZLpszTp0h+4xGvif/2oCcByxlCV3Yc/lz5g8l3hhaWUgdBDwRQatsqi/IdZIzKb
6ZTC4ThzEyK40/cBB/FNtmZfpexgtgmEBVsubHSzUkX8J5dzPc44i2XUG5VV/Ol6
oMCYduTdRnkPTiiPqLPBrrEs8QniOLLGkxS/4GItg82LTBAlu6iZJCo9gUBNAjCa
28Li1wtcZs9/HP6CdClS+OILCQoF5ugtfEpW7Sk1GXa4G4RsAMRSqqBXi9hnemLz
c7339nVObN0pj5Akqk7zplArwDXZvRc8urMHUu80DYhIYq5L8LnRvXWFY/eRlVml
s+qSa8kXNah6fApNARnT2IbWPpx/f70Jcvm5k/LJtPljjN72CihxFR8O95eUjdzT
5Iv3Y+zX4T80fW5dCM8+lr52HAfguL2i7m0DFBuco7jPTxCa5OqlezkoGe/m8w6Q
fP9WH5ObIGu2IMdH5PcveP21NhIrFtV2SOKq6FlQe3gOy8utnbAQqrF02lhIaYH8
YDn4w959ZTESoVKkYh5dgbwfPM6rTRHvReo4bHV5SVyZJS54HRrycxd7MkO04wYW
EZJAn6TEYxyWMC+/XB0QSRxHZHKPACZidwzT6PaHCxe2HVMIqCx8KuJ6RGYqYOrz
5TJMldwdgenO50ljsSkHphqXJnCJKX+OZE05QoIczwJjv95E5KhXxE+Tl75fsvaw
x2FfMyLuS7U2OOvd6vdkpuoLgOCdZ2FQ7yvKo1pYncXZcW05S1Nh+HBXMZfxEfcF
jAhc/WM0sdRQfL4YX9ohyNS7d9BADUi3qkq8tNN8OtQxFy/4l0/Ayz8hfVWJde22
KuG49oliATPWfiQE9FTjlSDaB0YyVghIjLdLC+MAWPg9WGSQv4YeahnXnjTffIWT
qNUXfEYrvO0gv+BTmvfHnB0bdS8jEBSypal6LTNetxSVYV4JjGVtujyZhI1Q/gYP
cJR/Fz7g4mn7fm9hI1aTdzQWTbcIqYZuuUHPuBcsru5DmKb66V5ZTXvti1I9Jk2/
/L3ThGZstaQQC8eUPI3JQXPYl8slHQ+nNqQUJFBMHp7WqO8+zfdr0aw+mSqODsqe
YU5P16g65arhC/kbbaiXx2Q6omKhwyNtasZB8GEOTavA/FixGu0d/xv1h35t3ahY
jLA3P3S2x6hQOsPSJbR/PJhmv1ZMiKNFtdWp5uxR8Kelm6+PaQK7dQbWTC8zMERD
RK35HjYuGK9Tp75PkHc2gESDndb8ylLLbzoaKPXfZBAYOVn2UVdUaMLrnIMaavLd
p3gGxCUUvNUpN3WELQcxYbx1jm5Dm48xY4LzTYJjAfeSS7ztcBYbHQXlepCyeU+4
jNzr9DFfs17pDMKG1K+Zgg4A2NsV9tuLlXumGBhc+YBdYXnLu5pRwaEBB4RH+UPJ
gwdVIUlFEajK4f6lN54zkWOV81TQBcHKRqR3xUrRhdrQPw4CIUOWy1fAuxAFJGDh
JiBtrxDHVkxfEzqJ57bhvALq34+0vMEjM7gzRpK8gDglZafL9F3L8eJ3B8XQze2s
bifdu32FLdehrq8F8M9Bbxja719BIzgD5ZGj76zULYSEUAfaQj1Y2MHfEUUBZFiq
y3Ot08BDFb1eqvNzChW6g+B5DvgdsT+YgzFeKbS0sxuNu844fVVSxJ5Obld5oyC/
kQ7YiX/uzhuui6Tl8fcDtLO0+vkC5jiWxJroD1qu+6um4b2M23QsMz2FFBMlxaov
QGkyVDaPdWB6JORWQbXoXQa8J0lxKBeGjfaPT7xTd0mF46E2SA8T+knVus1FpEth
dFTO/cpawQGWD3tIx6WhQZiZvYR4dMoVf+/9DGDbMHvwoT6fss4e4etJ7yyPP3pm
zbjR4YgTe0Rv+3NZNh8kakQq9OjZhPqpP3XcRvCn8Gq1RHKG1vz8suWDMjK08Vwt
eVysKHVta2qScRnCDAUfjEIXQzF8gO4eMSNww1cO4UL0nuWEtb8LHKPn2X3bERNb
grNT7Crki7+oIAEFAcw/Fi6ykAcMH0WQs+sbfMqIXou7GZ+zzPOqbiptVqqsX84y
5zVXYUj5AWsJEYVqAxlxKhmCQcHYVC5egLFIagzCeaqIYXuxlu0B2cCBeASX6UVl
xtvG0HRSVDinVxIsvwakeAr6es+9WWoR33wDvF1wS9coMMxClYDuG8wMdfzim+xJ
cTnJf3vlNOI5Wp43p2IVdqGaxOSHuNrgwEbgAPgbWQ2TDcq+NrOGuMv2urVkk9lK
iOJwCo2fdfSMt3aCC5KT+eTrJn0pno5ORQI9oKiueSs1yqaiXrS7DkFoqDeB463x
LZtuHWxSBGg9FT0q+8AopMMySzAcjGG2sxg65Lgg6IANfHtNpmPpAPoGopcEyVGm
/GNPX7MiGk8XX1miTVT+iu7VNxjXYzFz2InmpcI7wfMOcOi0Q7PEKnnMUUHaFc6p
fJ6Noy6IWBWmdhpDIFoQ83iFqASBn49F+QP7qJQmtghpaVrJSOjEYIdoSAnOFBqz
IZ2chOYrDnu0Akku7A32qmlQ/MnMDsuLefW9JjcikyLh572bhWVTSsqs6S1P1BoS
zvJCCX0Z+E2HbwfyKhUeM5Rld77ZBZm6L8+KpcbkmiD7NqBjQal5TaPa0/0gqw1Q
2mD2aky0mGEaMv+SP5VyCbAYBSHPCKtOnELDSOLTxVsPwayjoYuHdvhAC70rah9x
k/mpGdn7rM1fhPkzaBWXKaLggW2w0FhGr9jvVzJjB1p/7Kbtiv0jcumjMAul+OJL
YRGoi7bGBSl/aeUN2IMsVAOb/t+UHcCZjv186o4T9JMz0WHXvL7typwp126sUCvD
33pRJVtTHe0vL8OnoxboeovwJ2+BjFrJOwUf/YvXDz66ox6iQBHmjCUZq8RVfvcu
SwVb7z7Sa/66xa0/VDsiPkgynaK/3Rw4Gr8GJuRuxTTsT5paPADYbY1XrStFzd66
6sDI+gwGBSrZrvud6KMxx4jEm9dMjl+50UVg1Nd5s6OyLMN0OVjBGpjQGg+jN5OZ
ldKHXg2S21pnXGZyd9Yp8HWrnzXb6cLjUwvHbtWaKtG43BypMKfUGa8yyZvi/3LQ
JBhnM9vd4HesuHogivraCkjC7JOThXZxov46NERLDu9mqihrZad47Ud3Wacy4rgG
QzOKXSSp/79Beb8/3R/DU9f1Mqby2WCh6Wrcge8O1x6UcKxpklB3n/YVnnLWFtSw
8+g0oW65vyxNFTrzh3cX34EQ4+rx9z7nR5lYpR2mCW4Jw7OXAxD7eSpRilCSyUsO
8/xCOE+gUUsGaD9Vqxen8HP6zrymnKn7chq8x74BBWKnpHqpuFFYiNTOVz/XXd8N
niLmM5I6jQdHHfxu2Spj8+zbTbuM/hQvH5ZZorw1GEL0NKwRh8UB44vDd7lqhetW
MQE5ThRt258u/euI1cjjAZPPTuE/3Tw98dk6lLswC1IrYAP5UbItSrP/Nkh0NctG
0ov2I3X78i+HZiOsvLpCysfQK8RxQ31b4dUFndwCAIIBr8/VlUbgwDLFxAj40Zx8
ahaebsuQUbJ26mfJshSJZrgsNmP+EqprWi/+8bLx5S89yOIQS4kYma8/ZRyviFFk
O6uK8WLpup2NZ5QRYyNXaBTIf4+naZmjBU3tUJMQEv+O0klYNa0Vp9eTmE2GNMFl
zvncIaO0qdUnteKK3RAY7BB529P/OhIy/D3PK4rYaxUYiX8vN+W1PjJoa94qCwrY
0fNjh1LiDP/gMxbWzzwSdkWncOwv37mklZiSi9qKSj52NFifW3fM1zknHR9dSFv0
vrsbRF65W4p1bU39y2eCOjP3LdsFpC/w22yfqdVqDhmMOOJ3eUl1ylszBdAk6S4v
XMePW09mlSCZc90chaFTAWbrNeFbLX49UxztnCCA8bfFKiZHyj7Yy8vAT9bZJWvw
hDO2NrfwQ5bIWKg6kkXmevDDHiFpwjJve1w8lrLG9uS9U0JoBGaicyoOYuS4qdAE
O46PRvBCNCZXwFkAmxNGLzx+1cgJUVqGnW1UsYbRacuIMA53I8Zjaka/W/bZuMBj
oaek4SPAj/lA8RX5c8GhALaVv/b16SoznsFhnTLznR9n+pCeT0duNUjPP/5PlKoW
f+dDcyhYSgiATMghEALk1faeFs+hfGto1aGWiUOSRWe5wbyAE20YETlP6lpAc4Pr
0troXrT41/s8DJQQuIJ99k8+/TBcesOVQBd5/95pejTEGyNdsv4Zzk6RYluMKAaE
BVDoe6+nAsET6a4uOfLtDCUQ61lUZKCP9phhBGOmeA7e3dw0YqGrQ4rVR330wrGV
Kz1SsBjN/vjqSp8LREye3AT1Jmd3dbQNCctuqunRlEb/Pcn0jg9PH2dWev7jwPdx
U1t1zCvzd3Rtr26Mu6RQjgAYffadrZjKLHRQeab/GKy7ipDvcuPIJleB/wkP3wB2
zHS4M+dZDL8z/UZsNqhXNZIff8OwnDTk/HIypBYzukXlaEplX/JCG5rxXIr8/qCK
Xxz0KzawVKYbiLT3KGnoMSyvAuOgpZJ/tt4ugC4Vz27lcq6A6A43X3TYrto2tCTh
GW7L83A0qRxpZHG0YzTNFSPSv1/81C6ItfmqjKff1xwe0OMIG1jRpNM45aleYC+i
gO5yc5pKXqe2h/zrOBnU0ISOhEb3O6BbkxUz0LKaYMdQYyYpVkI8P9MtNBzuFScC
PJQ/7iWFGd9G7JLRpV8ANEQ9kfAUUZe2LYnl5p6j7MXMJ4yRrczaKyI6ou/oipcV
yx+vm/Mx9h/P+eSVH+ZMriGHrZV29KsJecGs+G/gJo4p//1oOHEdA728w583F3vg
JwujwaIoYCzQX/nOS6cOXaf/3V9kBrm3rEFGwX02MoSFbf+h+meX3lZbNA3ktriU
ZWIgzqiApw+IX/FpnoswMdCxYbR9LTS2LEP9qSRJ+1/15ckX38WCC28BbJqTOqaW
YuIAnuAdSTArXtn1ObX/WP/YvCJ+k70LDxcCmUBxH/NKhPj3BVa8Sd0tyuMNg/q+
hMAzyrcHsYwq9725TLXfVrkobqAz/PiqVircENyPqZqcn1wWmLNwB33J4yioUqcf
pqZTN/qh4Vtksvv4mb4fj8/Fnk6RnRZHlCWIQfx47PEDYM8QbAkdEDCc9fkzHK6/
LwZkWylVCj8qSnJWH6FrQihpllVfVxVt2cKrQJKMeKk71aa+Scc1iWRJOF6EKUjT
/iUVZn6anuEE5N1P4BCQ8979XDxVDSJN/v5LdVbOWwf2gufM+fs4welt2lvRSmqP
i/5Ih5W8NpTLyvD3EYsLwDS7xS4CD3J6ZQjxReQ2+KYdGgm+CyRoNrnAbz6g3wnd
D+fgOfeCdGWXK2sfuGiiUGD9n9XstNTAITi6N2xE0IPiiJq5nSgRIkZGxWdmE41L
YBTKWjqGcLI1+9yB0INiwyN1DQITxZWb+oJWEhoEhIzhkvUyIYjOevEBHcaU43aU
2hhDyWwtbHxNKjGSc1eYHSEkvLTkXOllzrPtuG+RbX54eSw8ysgFmyFeRarhnRG1
T2dIo4rUJzVYjWJs0Sn9L6lS67ht5IotIJZY5KkxySCdvMnlp9WDF6hqzVXgC94h
DMcrLWPV2DFu/y5lsLYDnhGhZTHQdlW9N3W514Z5Pk9W2h8/I5bYNcMK6wWjOSK8
PR/4EjJvF+5JvEEXugyvn7PLsfihBA/AhARrnlzrOuHOJZ26EA/uUpD4RzU27v0j
amSOJqoK27EteY6lu6FX2UC2hwLE8GSoDMlR2k/K545bnL33usC6BWAgzWXPxJ5s
+A00NMOlckL5+Am1WpSkfKk/C5kyHiiYqWtrolKkEo67XoiRLf9+RBE4WjbZw+/T
5Zfw66lnuFyJz03ZXvvhugdnWkJ14yb/nY+gZOH+Ti1r2+Oh7/BdKKfNQB+E3dH+
G9wXzoWslj2T3oOU87CBjMqZ1yiI5ZzD6pk7vFfYbzFlhRlXSz1JMBtpkLyUVToo
JNmkW1p+vKyamSuY5U9BWH4vP4v+VXRWylR3yvRED6Cca6rzNq78HNrm8McCXpm+
CbBBOIc5iAkJCsEw1xUuTm9Lxx8P1LUma5gb1jH+JYZL0HMAu+qVsbf684W5NWiW
WiWrgnSc44q4Y3if/MVnQMKKwRPcXpd3bMU0pXIY9fYLTfYjtNHcl0LPKnaHEIxd
YP5TrsDrDyOYMNvbmliKfLRzj7YBMMTUSMs62TCfmfpHezLQBodfzH1M51DAzJry
PTK0CuyFADhmYKYifmDnJfx3+KnsJUqz3/wi3D9QPtgf91BJ+lEfG7QsN/l49vUl
zCA3bX2kPX6UwFGGih505SMknISXCFu8175F1CXROb7KCX890IpvLN6uaRLwEg95
TQD9C8Cd6ERUOZ3yOiOwB4xzyjt/5zTvFjXT6FI9aFeAYf1+V+oSGS7HTO22cOP1
Yb0gw1J5kO7YH9Fp8C9DouFy3Me1a0uDfe3vCtUDVAvDn4B7PvP9j3V0OfBUyLx2
XLxQGwtY60+ih/ChWBSfYEDKkUPz52DwrBYq/hXdG5uA3fAFi2HrN9bqyVsI8mSk
Q968x7OenCOxLt+hDpgzGBIqJtsPyqeDy0RSZYKd61TvcFC8binOsUxqLZriRQWe
vd5ifw1Jb53VrM7XjbwT2Ru1sWQtKF39eAsNQhmFmccbiU0TEGT3r9Ux1qRt3Jhk
4+nMcEY4zky74taXK8VJmb/U6kPHbXTRQbDGqT+zJfVDsbOZJ0vCYaFvZ19vmVT3
nxNkd5U6Ua3KSTSQ5oZwvEVwQdoTbDwr08Ml+GDwH1N2lazWo23/2CegFTGeQSIh
nimFYjC5U59ghaYMWyLEoKc/FdVBVUWWQDMdeir30lqdl8LQBB+BdwAt3kNSSmAP
GbSn40bJ1bLLEy/MOKgD9CJ1ecY47b/8IKAPgVYhxQEFeJT0aVet1AcisHQkXER4
WcFBnHqPlbsjOsNvi0ckdT8cHawWfA+KCHAx9Agl0/rQ1SFyiRsGhsfleXy0IFuc
u0t2JZhSp1Jg2cykAsW/D4DMN/3XP9ubCCU1YPQJp7YwRRSs7QwsDZp1Cex+HAD2
hhi3tsh0Sh7bKxZm8EM2LZTh2MlHwZfw9T/xA5lI3cUzLu2lOpu+Xnrq97U9myRk
0le0+RA11aKlgqxgNEGO8XpzDFNzksvimIKckwLn2/nFhbiLLYyt4UKwE6+9+4uL
vEVvbukcymimMmXG0YkLMPfQQQ/RaV0JmKG2Ne8vDoZYlRxR4XnNIhDV8u/K+GEN
lNH/XrMd81kfgxF+iZQsFpD4SUZESp39B64l0rk97Dd0DKm6bQc+un1wxRRPF5dw
qpIuyrjQ2EJZqqQCyl3FXmctMhNiEUdvXegZ5bCY+tIxOp4PyTCfI93FYiIKWORr
dpz7t9+yJyhStdQjObaI+un9hRgcDjQO3sdogn6vJdOoyy1p9dmp/MFpwIos0ocp
R+EBS3oRfdpbdUuUDN7oMCGgnHGtkjQMKoyaEIfC6gtrwm4SqBxANrNiIohCvibN
bQgGTNnQ8FK0ItFhU8X4pN3ZjXOXIl1gagJ6rs8T1A7OOuEyrbHbl6g1UAz+oQYN
UOtwlCfHykTe8htJcQ6GjVR4wwnlgVfY8A8CFDS0C4pSR8QNF2+yAu/gbs3HDgNU
Z3DFMQJPNyS7N1pYxqPpqAvXfEKL/LT3/NzoSEWEHikgAvWzxbDc5o1wlsq1rium
/hqYnrSicEQhh3cY1h1MOIDtiqtu6nYYcoPM+4b+TF079fcs8/+rmDqioRxsTIpg
ii+c4Lma5/1pGNRwVD8oLbpmcUfH/pwuDdOR1cnlOyvJK7nL1Wj9dmbdRvNxzB1Z
O8xb294jUjAYnZgIZxTtDX7pX1L5fYhxIMc6yRXZPdkcgFA+1unOCSNmwU38Fedl
bDnkX3rlq+sUi9lYSa9usJBVAB2SMY7+SEqQ8y2dDQA2Pklleuh3tQ4LiL+KVjlB
niMA6q8QTTX91BtgD9BP67hhp0juCvd1cXW/frQIm/M8uak4nXUAKYByoRxFVTaV
yzTkAQuZGpwvB5I99XBCyomjfziLa/rwod05Xf4khKuzpjZT5XuaU1IvoDNG9SSj
2GgkJPkMOx33IQHVxqz7hQQ45XbSsRKPLB7bDf1Z4uWIfzp2ph6sNuw/CdrDlpKQ
pJTDQ6ax1QcDrsaKESVzWhBoQRwfjcmZdvGVw9ZfZoZm1bj8wJu3M6MYTMQ6muCW
LC14qtJ+7xGk/FXc96PkE3pPsH8SJmrwWQJgm24LPj/XTSXhHqUKoTJTD0tPVk4B
hc497CHx6rTw+e4Wx/iyquKYI48etDJzH2//sdIF6VNt19iHZ41Q8eTvtuXtckUq
mCczMuITz5q1i3PUhqnTqyGhRHJjs1UsVdJdYlsUVbT7x9YjXyMIUAtPiYgHQb+f
uLUe9GPjYZoIJ3c+KE+u5Ovk/XJmllcC1rlFIvCRkgnHRqELci4EyzkGKezAbrKe
UJZXZOglZw3LEInFUOz/F8WKiT9ZSXupqYEggbGRS65UJi73bWW3hx78zo3eU6OV
BdYg5ya/ZbGirh0n9V9h2+1tPDfmUyB0Kyd76q0u0fNHTWG2ef5oAo1y2ssh9ZnE
WXh2nDBv6B7XnZrPsqspCy9sK4PVJ6p7sbGj9V6EJG8hIOIHIkqu7mHDyyFO/nKR
AYUiwMz4B4VeYC/lSqbw7/tPWekTRMtXNJpxcBo6QNVeZO8ZA5Exr1tLFN/UUAUC
j9vYrvLha1jYMnwyyqDH/HhiQ4VjLDPMBYS/bPQutdkzgvm7B8K4O/g45/aiinOx
FVTXbI4V4IZrZW5kgA0dK3xW/D2Cnxe7sLvVXPfvmqKQX3obsAUdx7TrzT/fLD7b
yrXBC/VrZ7fWZ+6e5AQU+s9kKRpabqlYeP5dS5xpgNynf4sK8Nc89OktEv1bXlv0
gLuCF9WoK4aMRA21osseOgf6gI0t9DXtRz32eOEtG2DDxXpV6w31GdcKaOUpPx8o
hHM9JMeO0mSd1DHwpFcVAMbL89Oh5zaVFz/iuZgZ+UadPWWmxc03GGXq/opuplMJ
iJOjDCuyEVLX5LgRBStp9C4oDpqiVHG72q59I1LI4xX39+Ryx1dvYb9zXCYJj+N3
YCS3NDVWAr5f9TpCvuy7pEXcPj5bFua3mOq9iqJ6DRcth1j2U1QJ7McRbfC3zYNW
qCNrOMFWrLyYt8lpgpov93xYj/Ptcxkpc/ernszFgRs5pBq6SOg8cGZdHrTSnyYc
/4dwe5afq2M+AMdGJ6uhI9kbYRRcUC0uP0UAqueWV1pxCHV4tgBsjkGqjlBWQF9Q
M7VaFQxey9bawjSPzX0XoieFn8iGCH5D5a/B/s42/dLOnv5mBpwcq7S8eyf3jCi/
fl/CkEDOeb94z30WIq77PYGSYHxKeKQ1CJHsSllMaquDJ45yHfKOz/dXevQdrwBb
9IfoSXbG5JUZmbBmRvfCixUio83shwECtBhqsCTiWFwdCQpqHLyBKalcuGQZ8Dvm
MRBW7mN0fmR9h/cRwI21PxSOKUE0YyMSzF7lO6YymLcH5KDpXUVgQrcmr8dt5G1y
A534Okw3qRwGDB3/nYswtw7PKw8WpLnBy9lIPU9ax7VpH82lAGaKbFwzeJzC20kT
KY40zwpjAk1JoIjzN0FLZ5XwCfKI3Ryw9d/c666aTFT9XmTSA/EAgYIyJ5AbuIq0
1sQWfAkRyLOpQbGdObCP79+6h5/5t1U/GZwhezl0p9rdwPtGKn3Ov4pE1MFbbprz
6URFddOfdHAxdzHDvf50N45LQkzEXJAQ4hRa/eWYGov2VVW9FVMF9ArUH62cfR7w
7KkanvPIo6JAcyrllrJbnLohvHNI9HMzD5FBUBvUIXpbeYCaWmZUz0hvqoJ4N/6E
dzYY0Wpr29NwUf+MKD4u9wELUrT9xvQ5W4NZcPrNTXoDfx3ZThwwWkYS3OEE+lu3
Qvxou+YpN71GBp0ybFUJSLXpPr1RgzP1xXe88z7A4ebJV1rQfe9BCiq7MXdW/xbU
R4aGYmHcjM00s2xYHQiGKfKCbDtdQwPCqMz3DSngdxIyJnawPdcmJYXvTPfZwZY6
k3SWXMirPcyjrZTAMumGyHuWmqNo8ipCeuER6x513aqLkFqu3LA4PKNgSp/MhNhA
MQQ+XwPjRzMaSRYFIMV4W2XVyVRktCVNAHdB5NZD9tNl0g67jf6fr2wpKdDe1cTA
RgDCKfjWRtCYIajxVFyG5Rlnl79Symt3eYIxrf7m062BpK1Elogkf4tvdDagjs9r
PsrDAojOJ9v6rnPDVBwxD3P18caVW+kAMIO1jd97q14brGPc57qSOT8COT6YVSc/
d4osX8LEBKdqMEXslIbDWGIiwbhbX976Mg9h+ZsiuuZp0TJcZd5nXukrpszLN5UK
FrVLMIJbwdsOXF4iJFfJTdl21Gb5j63+Ao2/k81EnTUD6oTHKgqt5NgyiUyWub1H
NNweDpd6tkyXCPMWN6j3uTXgrtekFSNHfBGeyX6zjLQjXFWHD7IRYCf5YSpnNU75
kCPUwpyDj4vj4uW4qN6XlyOAgXKYXYwtOh83NegXASOvG/G4AsqoaI10vddQIdMQ
iOYrh/qNTSyJshpqdybDSknrCviuS7UDknhJg9o5ULS7nQMQajV1OFwPvfNSSa9D
DuOKZpKSNDfIKxpVgu3DgKxXYSbzCdZZmTXRoH80rYPN+sW4P3maHueh1XnR/GgN
uM8FEsEDAEpaRRjxBquM406Lc0jIjuNM9TTVRiup8W+HOYdBPGNC03zqO2uxSDtZ
FkxRZCW6+44qmGjez0Dw2X8M8uOnGdO8nRDjJeTjJ6tUAEsdO2ie7ANpRy4XP2OZ
tpZHp1Jzun/tsKhNGMat/GSLNcGya1A47g4nVxBB8WWHounUjeTKTNZbiMPFw0an
uGZ0KHlEk9ul6Y2wU9xTUMrmRRpnh/nsm5ZDrzBX0VsXeoZjiqLCCyxingxckXlW
TajkvxCfXeNpe2I/cUqEV3AJ5ZfxkIevUwuLytJvtv/bMoEvS+ryCCEkpqV2chWG
X9L+d/ypBBBmlULw9Yp1ehs8ldHpZ0bimcjXd0iSru0GlTaopvdO/oy21ccRSyXR
ChB0hYDVwJwQBMBHywhv9OnK3T3rWrsq+V34Az2vpocN84BgQym+gHgW8XaGpmCz
zKVosN3OzcbIMN8I1WNfdvYYd93EtY0nm6bXm9Pl//W1Q3Sy0Eslts4mg8uA7MRo
o1iK9qNfDvFVxhyvdDBRPbHCzW+c2jLGK5ZwV6sRHmhi3HK5RwgTqGicvXmvVCw/
xi6JRfaetaMneWsQoZW8VtW2fEZEctAEbzJU3lV5H/Mk9OjtThKw53gF2qZOnui3
leWMaMylf+TVs7HWfojEMA5cXYoq9mzaUOr50aGvCMiIi2VyJ6Aj3nqiGuueU1ky
HzgnVZ0kHgK2+OMiDotIuTKqhfpO9G6R9Pk7e22IE6pA/44CJeLGXrHSFe5Erxlk
eViQH/7VK7OcKaRy3gkfWTLpen7nk+qKxteX7Csa6oNmpkBvlnn7cKF9xQs+1sEE
gtYbV90r5dWMBYaumDdoqhSHRTm3U9//hI+4+S8wH+J6WGN/tRZ46c/LJD0Ge6Zm
KAywhGEvTZ8jselueOgPL/iIKWd/9mJ17xCFp2Jj8/IS1WqDBa7eQYFYceIO1kbb
gWjR3GMqG1atArQKKLXubffforc35b1SfKHWvriXzq45Mpe7CtqPatfiojndy5BU
0VymVKC6BkYM2RPXQtm2LZy2EnkccmZ0d8VUnXtgtzNFgG8jltczUcWIM/5ZWsAI
ELVnVGX+Nm8mJ5N00932sUjn/URL3saEvQpS3bh2mftvtemf8gzb2DWPu5Yr9mXC
BK7o67a3kBjKXzdnBpg4OZCY+TFwN+2sF1lOigE5wC/ycMFGxCzlN2d1ECiq0w3B
lebVn0VxRkXquEk93EAjwh+HHtgHptDHHIn+3EH77jGkjDLx2Hdf0bhiRo1JfiU2
Q3tesB5CU1giq5g6qU8ETCd4SWT+aR8kQxFKFCu5+dyb6SsKnV68EPIEANOkZSRi
kndnCuBLuY36alXqxz1PzsvHPNLP6DyxeX4vpzXBzhZUp3Roq8PchQQGbt9N9anU
FLdaHC4RHv8JYBPODbNe028KRlZ0d2vI+cmSwuONQUarzFbmN7fGC3ESL5aNTEQU
BDeCzkxnf3JzUdhfXsXZ2d31eBuSdC04HUPl1q03TkYAyJcasXgZ/UdNDyCHbjmJ
fi/a+yyUL+onC2Bv4NtvU1qB4ZEkm8C8+AQHM86StwkLnfMfh1NSIP5IYTUzYdc6
ou5t9wTFauG+ndvDOfNfUemzoMwSXITdMKykADHuF1KlqQyNIm+L/otZsIL/N8QN
xb9/QdqSNW8Raaj4bJUmbEOb5yUrsX3M1XbYtzJXSZa3XmzDuFH1eOWyOpoyjVVj
4F/YJgZo1zLpKR1b4z8OmoRN/QZN+O4t3HreNcn6ZbteLf3TSR4kaOBUdgodzyQY
WWcOO1bNNh0PczJ0A54KHvLxXHQlbyeOwhr8v0hPrWRIESj7E+aRH1OVqb9WWOev
C2SxngEfHhSsJqLTIuHf5UXCYxo3kxaDvXeN3zbTKO+zwtJRCt51HTk5EOmj2mwA
QIat9++AiN9nC1WB8modiRvK64sOxc819EK1KqvhBdoN09L3mJdiH+L8sh3umUWQ
SvvKgARcJ5Fj5QvOfaDXqxTHJh7+7DtuG2aK/jF+OM6W1Y8HW1q1Xac5LL+T3jHJ
O9KBSIAnh+1UGsvoLTL4VW5Zw+7xNvL/3Oc0X6OMyXiyE3F3pROkdg1p3HnvPnC1
xiQJ8QSOAiTb/RvXJe8T1rTiYJDKEiH/CR7u26ofPfzJUAy4Txyee9UpcQh7F8H2
MvsSIAkUdZslRMyPmEfx/tbZVWsYSGiib7LIB5nlk+QSsUvXqYTIGSE67hQNeCMn
Cwg1vv7jSFdIrW28E0NyGwEvzwF4bIaXxi61l12LopPDNAeEvdnm+6XjlKI2icH6
wNrgFg3f5OxRDHZkhh9g2aNopTTln+vdDqOX3U7auvy9hpvUcQsMW+0mYJSSbm1m
k0vs4Hf2VOH/7aSPN72QQbG0VXCZTKl7PMuUYVdKUOKd7HnJkidL1ebTn/UEl68Y
s1lIMojCvv3fNiNhggeOTAsp5aOyxPWc/BpmtwJFKCYY08vI9sgmrUw/2ZbyHD4T
NyeNVRdn0gU47klatbfWSG6CrHj5gAdMqaixGN7kTmFEeORQ/Q+cRPJvccoge1sB
RAWZ47C+2HKa1QDcEn0MnI4xhFJhdrFxDwZAUBZ2FskIx1kJyMWjjJtmHP/O+FFX
11CYV9uBh8VnO6QSEc+P495+tSrzN+Ecywk7CAjA/7kKfGY0e/N5nogLXUc2pukP
A6h39rMQsKca81tMH2TAlNu6zyZH8bOFbCanddQnc76AHlh+6upbrFG7XhBDmZyJ
Tx0oN/RBR9ve7ODG6dMkzh4KhPhMXca4JCvCGChWwFyeaYEnnc7DUCUj62qSMu1C
bN2GH3exu/LMooxG761UXERgW2lmxeKUOLBFXKtsKAutZwMfyCUDDPBM0u5Cvy+l
t6D9OKstfIFMdrbVO8lgRCjkHMdV0swPECysaDkXbyT2q8s3jrhB4smLbER8dxCM
IkTI7niWJrSBvrZlg24M1cbljtD9bTNttjwGC+P3D2DZXnFURIim/FPcjFi8TlVA
JudxZ+hl+liYDgj/DeL+ghYuu8cq/Rpn9tPHJ2HjKYCgIWEzAGgQJPhAs9+VYCey
IfLehMGYobQJMS2H8FA3/7VZnwA9VJ6ydin/SxKb4se1QTRl4c2xKt54t0fr8K4D
B/5WyuMEO4PHi1QBMBgCHHD703LaWnYTVcUV51dZizoTqQRdDk75uUxzLl+IYtA/
es8BaS9zVp9PUUSUUEu+Xvyuo2auz7kJtRUtIoc5ybMeQi7MT3LTviwRnof9jLUR
qAfJegg6sfAOAxfwRKChnM/CYZI4gTVYd1B7iQW3HTnu9VgdjRKfsSYPSBoJr8rb
XY5UV8SMYBMDgtJpZymgJvgzUXqTwcLTzdzxPns67jfgACd9CM8EpAsE4fv8Ej6+
10WsPuyq2IZM9dDOJkNfZdGpjhHB3FJ+oOwIw186Vdgjg1UCWaZZWlK7lUNVHJ8o
ZSPLPlmvRBI0JMpdxvzzLpyg4lHYX9V5arB25yeJYBghYLaV93q1sqVaEssaMjw8
1/Vj24e7WJn0BZvmfYVCYlNmsqFfA4V5BNoxboWKGaREOsgo2mRSTKUuplVQjEdX
SksZM1b08DKK80VU3a/Dm+dB8BWd1csYKgpJA9I0v4aEW+UvdZKTD2VpJKcUALo5
TrI5iWtB3ExO9wrXCONjtFB+l+VksX/GHZVxMN5il1DyM2NL+/ntueaN4l0+DRdv
N9KdayFMMShCwPry4IHGfR/07Ha0cA0zUL8ZEqbZKwuRdz63dkLP3HJAPNK4b4Lm
8niczb9E8uZWzoj6mD+aHrVLcLgCvd0exktIzDNMmzYQ/aJ3fj1OjOgKdCKiKj/8
TkVT5RLtG0BCbUoK9dgl0LQVbP/xHgzn8c7r002EJb6yfav2CPqS5mdfScxOFSJ3
/u0zCdf/pUfG8nmwmo4+3MVsiHpnp2lyXMhzpPMBqDxeRoEhC+A1J+zYzjJY7i0t
gOcz2Gf1+rQ2qL5bvto9m4maQBK1jGmqhaE3sdCcCzVkeHNuh2IVTrXkW65OWuxP
5b6YN+XUpkCczoqi01zvOKXkdys1bYfqEimxJQ7/FHfAwTHTzcvyw0bdQpHfwzJT
X1uTGfveaKGHgPtCs5Nn8lWi5VIqSCH2a6ku7ZfdTjTfnm2PA+1yNKJZRgzCyAJJ
giAOmzZrl65naRTnGX79C5OjUOh5Y62lC8pwI6Bs7VxcvzanV4hr/rjxdDXGjuWM
`pragma protect end_protected
