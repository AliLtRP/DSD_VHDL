// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:40 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Vu01SuqGjGbCPuiB0a1LS6JXgLPyA5wpAFD36fPkBLTIrQjz0g6aNaz8ueEj0CK/
fNZFXSYj2MnFwDqd0gZRfddEG4pjT+v2Bnv+u/OtXPk0pt3JoyPpoaZYhiJ10YET
LncehCSVtsRH/5vNqUluBBL+vXKNDmXv2FoVfpyd4pU=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 11296)
MgaRNfBS0cmo99RW5/v4joyHUGPKBFt+NeO+AMgFNZ2a9hmdaF8xQOCnMAKQXSng
jBnkebVZyp3Ev3VxkFcwr30gzLb7vve7GEvvNhWVnL3tBoG0K/hCurBUdvxv1xbC
a0dSnBka5TuvgtuyuVzWGUxeDUK6XKOyvvcayYLhayHNXpTUw7ivKzuZF91TB9hb
MA/8avbeKKv4adxhDZEElB939aYFOhppZT61igsE2DtSq+XdwPxHk78mF/aQ9Psu
KthTt+4c8bjRNJJdbAxeQ5lsVGY93f9PZ/UveERcBS7m7PbEGRmtl5ed2gWfK3fQ
DqU5L7l4F41Bbs0ZTi/8wEZ9MGtzD248bnEGFKu2psv+59e56o5vC1buUMou2vub
cS0ifHUtxgYQEq6VbDNiEbyg/cpF60CKOMFrYhJa1GBfDDpisWe3X9wDKwlK3Yzr
LKYemXiJbUx8Y77l8dV7nq99Tr3XQLWGMh6F5h6q+LxvkIFRPMTwz62omll0Fx4G
GljZNpgGSx+BcXf7HRD5B3AXEN+CNkAfOZsSfhucdkfuWkORNWyBvi4UDuSAZzwT
6hKbWG16q6kfxxeSDpsj5xYoe+I8It8cSaKoWo2OUVhsmkN646A2q7K8o9HqqvZG
sLZix8mS4515+Xm2J7IqSlF4NZs9viIY0Yop0oRy+QuyuurBMnavCATj9h3qlW9n
5gAIEeQrI2Gec+XeUkvdyr2QO/Z5u6MF/fUuqDVN5hb0AR6uFPPw0QKrPAQu0DlE
wJLqWtY4KyhBKV9kcH+U9lJJp3/qgcuPE+vk6RDb/PkgUyJ6e3n1kDjGPiVNbNBM
63YCHcO9Z0pT09yulZqOZ9JqvYRqI1RJX04cnWCOv8M7LIVqXzZb2oghp0e0iM0L
b3KJZnqqhn2azVaUJIZAPB2KVA6vF5NFqhoye0N4md8AJ857wgt1VmQdWcH1bRky
4C1y+mjzYBzRUYMCrZmxl4c7rRsNknNccPEsdyQtrV3kh/E63fUZz5+NzhuHadju
UbmVElUVdjEVCupLc/MxoAVYHhFcD2Rleo4jhIDvbZo0wZZo4jDEPL+J9k5zx2kq
PWEFKMtf478xNwqZt4DqPkWBPEyHtHbFJgP3rn4DQZ4z+GHVd1Hn7VN+sQGfwGaw
OSvRt/dK+AjGTrH+tOXie+dgiigTM+ZNO+ha6NO423G8Z8K6QAPIP+0vUEiaJoiZ
n47Cegb0F6zatUkcxPEfkqK7jojLXm7gV33bJhkOsLrKBrY82WmWVtBgObWKuX+p
T6YrgPrYsdmgn8EBRRbfZf8p396xHRUevsCNKWU4InJlZ0FeU44UqVsUGCwu+FLo
MivuglezZX9yoHcFNAmQGe4oz6JLBpI3efzA0DSI7xfYAdxrXGhBQgKxZ+/VIEup
dapLUX39E9BDPCZQSXAJWEypUs8djOemVcpmV0S5E8zurEHIaVBERdV6eYaBRWfF
3PC3ANBEEnVx5z6rxaDjgLVMdtfMV2MGSf349WaIVJO+5nqF+FAmCSUg0r/4IhH/
LarOZ1ozk6+TDoPZfdwRijOy57uLO5MrShPGNRk3zsfKsTpyvhfylfdZAIAelQTW
8DyD8EOcQ3+LRc5gSLHHKssn8bFl3J75PibU40qhnbKKQkNt+F7QTXpNDnka+8UW
jdnyRImP1VBxY87TSOCXbrZ+E66MUcQoE3ZL3Z4ucaZC/Y0caZN7GxVzHnhb2Qva
J4oTMu3ovVAoDPmlSj8Nc+HKx97BGufVPp49CIFQR7o6CDRg/BL8qBoNnmiizqSJ
jRInpjSeBU82aIqZ9R/sFtu+Oy2oRskOtW4ERUd6/JPejYdf6VFylSGzmDEnblO5
Mr7UuC1dDUWGQ3OerVcEVbKCEVUGaMgyxn1++0G3fQ/EyQC405yJg60ZXzH/bxca
bM3y0D871xeOwFPw9FkgTQbiHBPu2ukwXQYRIcS3CqLPJAkELI9YFXVVjGukFMdf
59OsAUZ42uQrJfbLgOHTS8NkY+zO4uYX9trYuwKYIwp3u9EvT9HHIV3fF74BbSW7
rp0O8TXGQU3b1+6TYAqvi+LI/6YsUY9f130x+3E9mQh4kD/EKs7bZr+YaCwqOLrf
tmvtBNcEdoQQKpx5CQu505AkYiYMYD9U/8bZtxs7zTCooPEOAendKJTM3QDOOPH4
KprTziuyVKy2wwjIWYaTgHKt/AKdnnublZRjpt3mmWz55NJRuSmuwEEkeqsoQuHN
lio+4fB3L3TXvQZ9nUJbmPK/hc5gS7U8221RjrtBsTLisT3suw7pX6rNn6jqJVcL
HiazdWNs9hwUdLyEp2BxaU3Sx3eLuYwitewsrueQZb56OtAcZF7FqQo6IfIxuCDQ
6Wb+0ntB+0RyEQqqdJuaLhbpXqC0n6kbtsMZkt9dGvaYUzkzSI2xGvyaM26NVKIg
/X48gCVn3c3DUrCqx0FtZ2GwgGdKsGasNz7B814LT73VCwoiYesnlLiyd8HF+bc0
tfBn3p22PeCMJejL/JX9sFyaZV/EwwJxcRBZV+SJoFBKBapLuQ+UXqU6cN87TfRx
dLSPAvKbeOdqZS/be9bKnHf2Mwyy6wjG3vr3a8opy5ricHcL0LYGsOU7PghgCzSb
NvhKhrzSLi7CVblzOf6ysfFhoXlpalpTw6HQtK/sZ+ybmpjI3ulMeVZ/orbJNTQ+
IsB88Cg5BAv/eVNyhFErNx07cZP9QVkeUYQ/UOvEbbH39eIvAnylhI0j/KCrINNw
212SD1Vz8AZW5UfOzfGX9O5rBl8qvpv+HeIfPbdsd383KOdY2paEHPAR9qSBaNLq
QVez70Gv29bdEutt5tcl/seWJ6L8pIwjTsvmjc732HdvsyNfuhfOurAKxDTWVg5v
6lcjdzLGtYn25QopNGWx+pXlxP28jSKBqH5ZIPxcxP0/7FxtqiMh1Tej1N0tPkm0
UnaZ6x8mJMQ/eAH+XME6XUMoAYHgiPc6nO7TNe9hX2aU98UEvs29X6WvLVwM1KFK
/sIu1pdcxnmVtx/zFQ2n4sHmYeZOLPb0VP+ayFnsvj2Th1YV7dpKpKR5bE0J6H2T
COfTjvaQTBOBNFvV07b9I66cdibE6+WZU0u7YNP/U0/6yPhRW1Q0kndnbdAuB4tl
+rJxSXJrP82Qi31b+d1H74YVUJ0elwX4BDodoJoldhKzQvP5lBEPPeN/YZepgAWz
XX7OOmhllzXD4cDitCzykf51ZrT7exHhdAWriJQnkDgtLrkO9SpG7WXWMnRqA8xZ
dxlGRpB2lBo33KqmBRm5ZT+BJAzAwHEaZGluXrIoDQdhTJvOjWsAdGUNnINvuM9x
RL2XQudOqYNEBlgV0yRq3TTvF/P6WUCf6MHy1F/itJtA9tqDqayk55S1vuzrJ3gy
9d6GX2380ZihetbQD6hpzQwyk4wWPTQwYhBIvGBGs7TVGK/chrSS2o5Va+KNrEWq
JBk14lZV1BIbVJtPj/daS8Zh0U05Dff4B7skf3ybkZBLYNFW3cckajRFETwd6uGx
fd+AUI/wCN2xC3Ol8utkKHhrKYdEInAhI0FIJ21oMs510o9opF7d6jTmFUeathmB
qYudm9ap/nx6rCu67qcftZMcvaI5/m8n5Fr+dHBiCYB5aP2UT+CMLidm+QFEfe/p
AptBu1mg9A3dEBiapd7ZMJyNlz6TzflkOQVD1ssffpesBMdh/BmWSa1H6xfeH72z
rOazedkvG6wyvi+9M/xVQwleuyqPLt8jtt5vicnBSusjvD5eNJnNi9jeClhpxchA
SSjgjfF9KoelZVPdB3hJeU2kBw+CfIOfrRbo1k6YxCTincZW6E3wMYTAys/SsaOx
cOs31LgWXRYACUZaRI/gUIEBi2bgG+XvfQsem30fBIiTkLk/XlMi9ZYTuGI4q9Jt
r43rBukgYOXNs2g+TAqxqYopfkuR970VkSUgpkLHrOZIXPm2Ch/KyoohmHVk4GnB
lQIE6BeXCf/zAvB0RMIW7Say7RXNOo2I1dm/KEbUSUDNW+TZFvBbqMH7pJ3SaL8h
lrVJx7iTQlamhCfD6bwzgsr6s0+7YHYvMXVD3h+8SwTvLT94HGQMf5Jo+SKl3U25
KQoh6MFt2d414aRSKCqS7iuFv0TzsUt5Ala1v7pITRtmgymqoX9jfc3zHlTJ2U+Z
srdU+kTfzg5nFYrvI1FHsUoNC46ofNSC/LWIIe52gCWy+vx/g8/uBFT0P4yS0fgt
B+iDiRSWBvD63QpRaQXZVW0dgRO+oIzwH1VK9drpUNAjtZJpXlDcYzzVecU/1LvY
gwDc7Qsjje0it2tCYAY11WOYQVguGYAoWPouPF906qzHGsryOxKCZFDU4JPfT0ZB
K5HkuUZdeWAfna9ExcN07eGd0RxhkFsvqt07VDZNdwiC6CahG5kDloJU4hs5TrqU
ta6JJo1U6kOFQsGQC1D51x5bRwiAXDNviXYtWOcgu/uVUdodZLE22mioLcO+dfmz
J94W4I7MYOKxsWg8kRyLKT6A+HDiREnh5B8n0edE7pS7OoJIlB2L2CQSwiABdllZ
T9aQ6HYUIopKidZKYswfZr1U/x9IG55JjK1X7X40qbMSi48oaNI53BRgeE6pwipT
TdRR/Nbn+1yYeuCEM4AS57yMtmQas0DgqDjxdWJNOx2EVSgn0GZIz16oaBAI1gx0
9IjLdjPCt6Sss3CPf99Ug05vesXvCYHONIHaCFBadS7MhIO+yFvML+3TL05waziq
L6syl5wvR0xkO3h9AFU3R4TeLccRuHJ0kK6tMUizdKeSSqO32FjqEkVMlRxkbLqd
yrqBGqANeCFV5Fguz5PK1fRF08wLna99BvgXaE7noDjISLIsMnECIHzJUXHa0tuZ
bc+0BfW2WrSm4X2Pkpo7lbiFLqHlbzcZI+qQvQwws56XMuIHyfIutXAmn8RG9+4/
kkcvFqst814mnxBm9IU1kluGpzIubKHT38SSVkOO225rBJUziCYjzTSrpoJ6ULPq
lPQU0y+a/5E6dJhAurnmuvYbCuhuQEZ2g4D1b+wn6xNkS48wcxBuaQLzLOTTtzfz
cSXjBQRMI/Pk+KL12JCid2pOJgXuI0P5ec86HDRIcXTX8skeGaBH5qF4lPnaoBHG
egRsgKrWTVE5YmujMIiH4fiR3BskeO19dAmm5B0PWCjsCvQdSJLNVGXB0YxgxydC
d25+nWoneeq8YI086CRGEmF6IUh5O6dap5OyT9gjug0FTbYEPJ+N22rquGyCovmb
gHDguorimknI2sQSJPGP8eQm6+LCCkS9/z7f8/4mUtILoY2JF4XuiivWRV+s9EUw
qOKxf7B5dCDRw73OM6ShU5386rtZzG3gxBaW6MeGxs7KyZ1Lvo55yNDEOQ/05yvY
ZnegaPF063fkWCoHyfSN5ZH/UCkrhg0y5ZkhHD2JcesdMVMvYwo8UhJ5m6JIWefz
0CWzujQmJu78jduMRItLMvXNqEDfE9jm31PJz93saurNHQqvDij5GeHiOzuHv5VV
09rfRNHG1Z7RkmoD8HXHSC+8bSiuhCGwtKQibw5iFXkfs/I6TcWqBhueBdr/9o56
OLQLwS+7Sk/dbhBHxd9BCW2kEMGSEqIRRE8OnU8lZWu1mS1UkhtolS3Hcce8MWIl
7FDf0HIJzfLrHZwI7v5TXjyUUs5W/uSV24F2SyNPq0m1I4ZlJgEkMlgIJB6DyfE4
9BWd3lBBNmWffRy23r0G6GY5uBrdktO15poAEol5tT+WNRwb62JtBxkf0Lm3pAcZ
bZ6OI0kRk3uSHmoZi6CyWz+3mqbQ0TTJo4sUFT8JtsSYUAJSbdIBlN1naSmiNxtb
4ltR+FdkbfhGuv3HDKtDnQCXgXcsoU9lUkD1YvCU2z3UabB+S8ssZSYnBB77bOeR
gM2tHVKMAcQ/8fUinFclYzAAZm6J3UMkAgOttvfgnTjGEbmwAR10f9rIq1vKTB76
DMyiPd26dcSmfQQFp3//BiJJsueBhxSZrZV2rjdt8YLwTEra5JMSP3mI6evqLxnK
H+mt0P5tCyp/2+wBq0zUMgkMbvZtITEM2cv1MVkkFPh1c9TGCuuJbDSWAU4NJpQB
gVYxa0fW1JxNTsnrM5T+pV9y262tET2fJIYMqjF+mYp3Im/pov/wSrh6YgdbXcVD
r7qI8AAi0pZ43Clv5+NgzPkFzXmPvUcd3lq2iACmq/O0uTcKfBPquu/jglpLCfpX
Q0myMsfZhBpYdNgPslPS0K8H2VONOIXCWw2BzOW4Okvg+gHrJbrVLGAaxALYyVGS
lCfftcQ6sQ4gA8B7yPpUJn8XIIHCE4zDOVhg3VXSJK3nV956nOrTcBBZOuId0d0/
q7LE15Tc61l4qnbu7HQYn4fkMbUZQEhbtr3BQmA9rfmF6WxicJMMn2WdqhgTRx4r
8qDlqyJah4rvQsJbiglQ3GoSIvNWrNLUgkO7zUYbAX8NWimLtud4usGmkRZDdnpp
0QY13eeSOZ/qMk6upygrQQCf7f1LzUP+o5gtev8yZ9jBmwNB7AenGFzqD3wWmip5
PcEc7ABMSaLPk+qr87N036KYYXUWZgI3hOl+SV80ZgCxbR016ZcVv97xhV/KPlE5
Usar0RcggWRHJpx35Q8Bx8yQoWKZok7UdAeHuqMqV09waLnt/zhVGSkXTukxV+pT
5B49S6L5CPGmdxNDQpaVeYmtbch5UH3K+OGDXYJv5HVRTdKNZ9A9DCGfGccdGk6E
/G/BYrJysZBOpss6VEDtMjUUjFoQRQZckD2BMZhITkD3iavRNBq/bW6XUWIaODb5
kwOz5vTAiP43ejoJS1UJGFNOSpHw8Do5X3do8uuWpAcsGyZncBsgzg/jVGaIJI2a
wFm9skE2xzA7a+SZm+OjKv2iLN+qtE5SIxMtKAL5EHSxeLkxsexnoVmqN6wD+ZYM
P8YdaK+aBQFqioiqgnmXr7ntD65ChNCy99MBNDU85pnjeXJaEYvn9EAkjFpmnRfv
MhnNnFzDmXTpY3/GQBAoLfR7hpgMoq/OQ50yx/eJiFXREyExzgxhOspTgUmAlBcA
LIIepFbLPIqmeOynwFWikwNyBlZwwGJIo2kCzFvERYg8CzlTV0eXJpidXOZ5IGC6
Ocr4ULIOz54vER0TvoeTS4OIVRjJiQ969bm2xc5E7hlz5ReLfnz9W71tDuiWazwi
0rSzHASOSWHQG8PZEGbc/VelPgcklqS6HHC4hNz+EPNawjZxeT3cim90jT0ka0vI
c3iod47lVC0NUht+uM0U42R+KhlIE+si1Nq4rqDTJpuNIj3rSZ+HXJb9B1rYs45O
5sP9qpJA07W4424twBMa5nbT86n69LtB1RmU4XuxZeMY7IuX7A+Z1ZSvawihqixx
a6VGC+O0Yq9JcwygTkwrocfy722lpTCd5AaYDtOxyrEdJuZq+dvR4IFQ7/dHcntf
tBYWlcJFgsWTAO4/pEPz3JNEHcM9Lh1ARVTBPh4KkvW/ZyrCiY1iBirZsmxdnokn
v7LzFh38bw/VvgGoIKY/yr+mSVUFl7NScKcwoDBh1vQwayBJmnq85gX3Hf2IHVxq
ZHPKSh+1TeZ0J5YaLAj+dP/GBSyt/IJ8uzBRDWOB8twfmk3kF/MHiTmDTUV4YIxS
qmTjSOZNN0VFVDqOlm/7izI1Ftprp2ujmGg/3x8VOZ4a6lif2pJKClp4t9cwyvNy
duauCirO91SdNs8o7t7mQa9KDXVTY7yOVn1AbM0aoUrBBlrkwNR+aff86mkz1abN
8V86zgGZXOquaBboFR0jZWlFfI/olGe5OP+Lg5QcBu5ZHgyu4odbdae6nTmZqAZ1
yXnGXCVYqaAe/j5wAT3Dzsv58HvlFV2MTH7WHTRW2zYlss77dqDkmztCuuO2OSTF
8T8opsJE6/HKgh+0Ep40/Qp6PLsbaTGHZ5WkjMQgE2KUYnmZCYk7RutNVO5M1pkM
vVDS7HSNJqv4Ns9ZvjX0lxHK+C4tbubDnxCRKX7U2K62xGlceZ3BOFXrd0QlnRnK
Lq+jhIxTBwNn5+/g4ZRNNtCN0WOA5DF4I/amMdrWZkraA6kEGmEzjFrfVBqIvycx
6DvP78Gf5l5WrNioRA0r+M4yG6jfQPGeQqGqM7+HDQIe64NcNRvcYXRoz02Ftuva
IMOlzOS6GKfUV4GAq2Od2rCvKZyzj4u7fFvabuYJN3nrfjGpaH11nWuJ0/C4J9Qz
mfo3ZdpTWytRhRp6rGMIr9BPScWWsTP8/xOUbratvQWMa8bGpTkbIcdkvXljROFa
lcuhgMz82ge423a1EvhzF5bzDjkHcs3nwLYPIhoQ2RteyRwpNtGvDBoaT4pAtYjQ
bkNcli/hGbQk9A1oiwJaoicy/emH6ONlDXQs4RRKLYUX3n9QcFyGVu1eg7ZX4JjI
mZOi1HB6dxeimEPgdy2oLluKJccQ2NqZWIp0Rx/zzFiGrL7SeE4zKrjRuDxlj+QF
NXrvbmpnzuU3iQ4K3Ch7ybvB+zZ4aAOBu6W8JSayDoyJ/RAcHwZCZpxHeGmNo93o
wFKkQbov8pFiCb7Fvc3q1j+Bt1M4BJwGouv5srurCvHqp4TyXkx+cQEDzYKPIyLi
gVMXFODJb3YCItqv9fZZ3xw16jruA3JGkZCNg9pNnSHlpMgNPALQR0RmlnnNlkEA
e8F6NRoRy+/cau/QQXqxNBQEGhqznqnw8+cwSmpJvrT+pjQW3LfgXtwzPKMP80Ta
e83Mo2m1x9dZHrhkcAkssvKDZjy9g7/q/6gJ6t5KtepjgwC3qIIESkFAM7BPlZ1W
47Q0B6An3uNa+6HkKiaSmHVFBj9a9taykvR3AJTb8cbEPH6fHJdfPKmtmXxKsi5t
qqq+GHgqvzFp5HKLb5lBbojYcVlm9boQq0yUtmPgEaXd5waqPuDt1/Bx+pqB6AwS
CNknEWBbh/GfaombDQ6kUCYH1Sbu8qRNanHwUrmEB4UxSt61R+1H4ddQpJBQhYap
P1J4KO7Td1cZ6HaUc3jd++cnOW9VhWN3sGUX1zoFigFP2tXKEkc13hqZj5seo3O+
6S2pT90ngOquV3qxKS4lhldlV+0OmzF9Gr3stnmoBYQF8QD/f+aI6kmBCc9zzvsA
yfhwp1gd7lCJxS5biOPFKb2VpbWhSpGrQvJs7MkPI+vIT1HWKgjlEGD5S3Wx4T9T
UTLiGfMxIAk3eZ06YsE4r6TfUSK0kjwsOIfp0KUG6dVCOca6Zs+VjTvEKyHUgFVy
0gv9X2qm8Eyn0uQeBls78Kg8VdWcLWk0g0Asz3TsXns0Va+VteokXO0wizfeIm3W
pbPJo6vZ1DaHP1QmPQOAgjDhqK++cPle3q4qNB8b3mHHn2GNZiSF7hnmaN1iQC30
xQ+01MfUs9sIoElSUQfATtfSjjzrLBrE5+fKrJw2nINhLbjhRNtGkfBxyYLrN8wQ
u2MHBqQFmAXjiY7Oqm0X9YX/sXuDRsLCFVCOurryuJPs6d+3S/GnaoWZ3ALXVLoM
FmMO9Y0XLRKN/crW/WeiGwMlR0CrtVB4w98g45idmwpAWaCQrQh0WKPKqB8ZVxpT
bomDqr9cXRXhhUpPJzJJ8NEDMHtrdlUEN3du7fdCzDl/jcC1VmhiXzGa9neGOaG7
AFGu/lsxL032lQ8ITS74R8JIxm59AFdbAOe4CfwuVpMhmIN7JkhWaehHg54cBr8h
znxP2kgbzqAUtp2X8oW0zbn6+7J+SQKElctjrVRGeU9U2I/BPCyx/5cnM8bi8OZR
HllfkAWcw6L8lEX5ZPQx3tcffnuPMfRKASpICwkjVYZrRJc4BTmmrLWvPJbGWemS
3HLfzlDGmi7zikW6H5LUmJg+lxH3DOg5SfCeXheRG2CDYJgP5pwKxs/E5wcDTiYk
2Blx3gOz7LgfVulT8DxGDNds6ylbBu1UhwwlDI6D5F7pz8Ka0X4/iTdCvDCQgYeg
20+Nu2hPS1QnDUMiAl85TjGSmAxgj5wlvw5y6i/hzUxGsXloDGmU/LpMPIgmbLOD
AXt9uJ4jawVjasEJwXPosLtmBlBJBYIw1UcSU+QTMDtKPIvUrFk76wTu/CvXT2p3
rDYFCduvnn5IDHt+S4TeAj/ADEjx3DUSupnul9ASKJUmgJYczp248dhvnniJVC6W
yUD5mCBOLtRVCSdIv7b6K1Tu4/MxpskuShLTvjlji6yZZW4S3v//RJ1Lq3flh0I1
4IMfb2Vd5PVCfFoFhtoyJF9PxQm+5UEJPe36di9prvTDp8TI/UBQdRHbPYp6cMbB
qa6CODMEF/+o0ToyMNgQ/gEWIEtECjwSA+Ay3/FB0SVoDswJS1kq8TBjtpUzQbBf
klRIRimfKe5KfUbwqsKcp9EEOaBGwREsLmNjYUxWaqgf2WUXXko38YLCcyonRsan
6Z4rUN+mL1iZoXFG16YD25HNrk2gxqvvPTPjJSPzqtDARM4ZVhNqB/BnUytfKmue
CvRIBtSIe147ag1vtbFQeeqbLFrzBkZn1jTfLNm6oDi4KA+b/7XPM6On+W86ONp9
3YRkY2AUtEXJ61D4127WpN7+TCTZavIFdZ9CJEDNy0iGlIlDwVGSpmFYwcC7j0U7
kzRFSN+GxZ7LBa3WLDvVo+wnAof0Ol0dA/QV30hjC3s/GRBLilfRpub+U0foiWB1
bJUq7OuARBcm2UJnIHXZ6FpZ2WVs09Cd1pXdQXigu1ecvChTHvJS4I01Ec2lD6g6
wrykZZWLqQWG3JnEDRHXrSqghP7dmuwrib9kADn0wVK6RTwo5qc3DXoeLYAcSPOR
mycaZC9yoo5Ts9Sc1BaCuJYnhAg27+2/H4u+Vs1JqCgHXNPo3Az+o5EdDKmOuuqe
tsASl34y4PjhM7zIqto7anfRDlko8s5gzMo/i4Cf3a7zEV+dqMyOdCSG4529XxKu
wAlZ+S5ahq7jwD5lcPr6UQaEuzxz5TCI+rO3D4MlPbh9C/UsHBhMGwF1jRQCiEEY
4a8mpfJIwUYUO4q9jmG9FMvvniWRZw3ywxAuxTq8s8PASNWYsnrq2QxKp7dlL8KX
t+WAupLV3VPXXV7nOO0Y5SlLE06Sr84shSEzhn6DWAL0EEmuVPH5DMHFS2CJd82f
xLv6mz1RP+VdflSp92etlXyesTUmTpcmQMMKeOa8YS2eC6MDLv9V3r7fl4l5dIBu
Df0ZpWRA4kmWSiMVtHw1JlB0LU5I/dYSYVXI5SPTjGdO1Jy8qbS6USmQy40/UdtA
VU1LiK9Fvoh3L73aGNS12qsgySIxw25k1BL2DP5mKiZkPsG1S3zsCFqAer3bewTj
puJcWD53MUQxutdm0sIQS7r/veJEXlgHAisD6jqjtCUVuAaDqEbdfdF2aL3gAgYk
Y0MFvEwwQufdx6cgsdjqqIGZHPOudIQmRRo12Cv/T1cvMS1XhQA9nEYhg/eTbDpP
5LQpBbATdQBJWD3MzfuJJ2QWLIyXxE2xzIdo2CoN9zJOEVw6xcrwGllQhcIVtyV/
zqoIFvqR7YKWmLDeuNsvqoHy1f/U85TEGDwmh4bm0riHYL0Q7K3Ig+KKKA9vGGjM
wWi/AhG4glKVqjCU+HNXH+XxTAdpGNrIvc6wC0ooCVj1WvZ9EbZzt4qeXZHziXrE
rurCT9PkdNQ/hj9ArJPEfrMexg0sbt+P0q8NZcaUrqgxWHLGCcgudoudw7rPIB+B
hBxHTqz519NW3Hh4HIMvByHDVbFgEr5jvA9FMDUeD/fe69LoGiQEsTSYKt27nWrs
HH3Taj3eHe0kO9cMNJ09Io0bwHKEegxU285ZC9Kb6TdvhF58yFHMqCFJQM/VEhd4
25L3DeJJUqtlMt2UkWmpzBaUyrsv0yLyh+lZ9z3UKPzke8KXbq27dYVuVoKpMwrR
L6QEON90wmQ0c8HcNSOTtSWuXH6vOZpcXSHDi1wxYQwOmY43X570XxHYiomntEv2
gGsG3Z1e2r4NQUb8Ll0qeiSA3OLJ/mfo5LGdqN43rHztQBOi9RFYPNGbV9tsUzDv
cBVwItu6gFPB7yez1VI7GrP7nOrGwMfcUJktfCdRLc9fxWCQSDFwwji7MTc2T2rH
xcGfvXUSNIeGKXZCI1iwwX7TFFRaQCaWWJ8GYMdEF1L2j6XdqkmdQlkVOvWqdgqc
JDSSZ5KB1T6tfz5jHNqLV/sKQNXhWK2Ksb8HIlrrjYxlHahO4Jx00KIAE1LZt+cQ
JZZ1I7nWb6BkQ7DThiD3AYs4qpggox3oeWhkFGwaFX78sEZqLisRSpK7tl8G3o+S
1hexI5+n2PIwoTZpoxtK73xEWi32qqShQyKfL8VzTWLRiVdeeCMvHc6S8w1/1PE7
UTLb6wSv9TTOas1Cq6kyxjMIrZE0Esk3/GAPrg3rfZzUr4FuRZItTJBL1ZOyf6oM
qKQnrY34mltUQ9USTJx94sBPOfloSnF9jY2p5KM6BrFq4+J+XWuaFrC65wxzZ1xC
+lT94f0TicdmCoZcX31iI8xoVH+Bx22oZNhXgIcieMWiK+V/w8iKt1CLOYkL+TL/
5YOEXmMRjLekcd+jVEF1JTzH3fNJdzBvel5etlP2yNNBU344qIVW3JfhvG7ZAaOz
6MwbJOJbdv6H1rfrynR/BG0K4vITwtWoLc4uxcuiQABY5kr196D0G/iOvm7vaGT9
oDdJEWb4Czk6SO94bDCck9s+clfSxBGV3xa58imyEqDa4hs7ZZUQZvNzxy6l81Mi
1Z48W/X1oGSfhsFZZsf/lv9PFiA0TvBuE7RNWs2aeb8E2h+Ld9F4XD53oIp78TDE
1TIlJgqMAnVfy9nlzxcxlJ9UYNF0HwpmD6MGBxtOtspNl26+Ps64TEG7wEhzJqKe
svBTYDauq1VYlDixHdc75aGjHc6aUJtexaLtp3yMUphV0KXIlNJOyeamycex3ZL3
gaKL6GLZTQXh8+mpgLx5jnnstRzhuhr+jvwDGo8ZB0gDkf+79LDBSm5erQZrk5CU
/Rx4T0Mth02gYFGd55/eWz8zwF72+2l7z86V/qk1WHMhxtwz2imMpaDglOAjbeFt
XobbtZjs+DLhyoN1WmXZhZLsc6JLUGSKy/Ph8XVMFd3WvJsTZkbHm90BP2HxFYF/
Q2t8t+fjSRCuxTwB7Tbf3M1rpM1kvEgZ2fNN1AcrncB703Pk9MkDrX8sfzYuUshA
F43lCGSZ3ysusWn6UTWF8hRZggpe+3SjoXHIPI2KE6N7TlEQ8bEJRLZmQDUtjPRU
mKC/QLv7B1Ig3qDTIZOKingssuaORWuYhZiTwXvD2is/olPXDnxVMNyzuBNfODRC
RzMYZrladm/a36QRhdV8i/Tb6NHB/0hXdcFUMuR63Hz9/53F48NNNv9lCAvlFJQA
g5Kk+NA35GnWMg6fO0n4zpwc05BZ93PI1zZXk0WqRzXiOhrbt4T7Yr4fK6br+C15
Pz4k8IxkFUVckAz96303CXcHppX5K1aXpE+C/a3R0n6YBLIv4F1d5/WSQKW8lg9q
6wsb/bn4E29/hVQ3nYskWAoN+uOUdwF8d1OVBiVlc3Sk1BxcbgGCw7lI9JVHlWSd
f8KuTvu4rIHiUiW3hhFacstut6b2s42W67fWfKHgACtVJYoQvSnfOXIhFma+IoI8
R+h+o7Znuq0F4F6DcGMIIZFqJsQnMRxVJbdb4Z01LD6hx2TGvnVWXYjIjUNC8e+9
+5wPnr6hFFMy+hA+LJHSMKTBGGhrRdLVXDIyWSgTECLtDtw53jBB5wMH994QTWGP
LJbn8piczZx0ws4EJEqc4wH00l9cNmRfQJjseW4reLOSDTAs+tlQ0P8jqulis5EU
Ztltb3jUaaB+fvyM+Hn14sUbNao+Zhq2OstIsbMfcRfRWUQQ4gCzJkgdiJPWXm7E
0wODkE/NF3Rs9eVKgyzIZqjY9pbAGdYBjmJCyIzLb5LpATLkLPm6SKly068GFuOo
0S8mMTFhS0YbaJZV15uRz9N42dbp/HLsmRAcagy/JMgJiZsLLrVOnuv76kvTe2r8
mqCzAsnQPHtDXJWvVOtZUfVyC0o/a5FvmW6Vdm2/OZc8u5uPoY30I12w7V8Esw5R
SjtHQeXuRyl57InPILEXhl5hvCzHYFHCoj2sOnLUHippwKD9gLUXg0vtKXEB3SGm
A9HneA4/q+0bMsBgLE2pm1+sl4dEfnKPDD2nPgg3N0S7imunNdJnN45c/gcFQUAQ
XPM/tvkwYPgV8/6A7a1ovX4NBxeuO8WdSKwSTWSD13zGfCsIomrNnNyNhNxYidhb
0r7v9aH8EIvMI+B1IAHmXI4lRVzK1MnINzHGlfjUWSDSqVJPBE31qIvc3U1yvcG2
APOtR3q5r41FKTPGrueb/wqHt2SxZhW9v9+KB0S0rHTEa3bmJR/5hsxpv3JxKx7d
Zk/cYay/rBQ+nqr8iXsb+BCJiO+GHVhZPa71WOp/ARNVBO6dhQPofgEH1iqg9GPD
H7ZP1ib+QzU4eNKp2an1YcSXJAOMrfGWNDm2N7lNE9ZmUYOqi9FmplSrEJC8kMA7
cBYFWpFxmdPk9uOZ/Kx70yySCiY254Dxh3eJkgBgAx/E9VU0RP+wxt4+IcZGyLeV
t0ikVY3UdD78jZGd5estFZsnCekrxxje6O5Z+ZJehtdX/2iI0lryFgahn7PLaXf/
qB469PAmnV7maR2oh1t1kAgH898jz9GXwe1HFivdlE5BHY4juC+f2AY2yXJZORVl
uDK5pvJnNDf12JugDOg6nyD+5gIX3O08W9TRv0g+ZW1hk+Cn2x1TRM7uJYmSPTBy
F6hIGWkSPSx3SyhxkhrbXssq8iZgDEy3NyezIascH3KPcEzwcEMEovas/a5q7SjO
r2v1oEL+wXB8IS8AzFgeO3BuFusG4nzUeK5k0X5LpfWhiRmUHaM1CXjqb7QCh6Wl
AKG6mE+NNkIo3ViWWhhn9Gq0ZQyG4IO8XaDioeaGne2G4BuvCqxxka/t9fm9ICN7
RtG8OYQfkzVEmdSKulORWUVqJ/YaH5dYT8KXBkGYwl/8ep0r08+NF8l5yTogWUZR
5GVCoeKw3gDKOXbZnVmm3BdYESjVZn5H2lUDjqsBFUGoXsZ5SkCU1PF/DpUzeBqo
xwdn7AvIA4F+8652YFSURw==
`pragma protect end_protected
