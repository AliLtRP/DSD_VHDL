// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:31:57 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
XLy+6MVWPIvOrzAjfTUhwKv5VKl++AQwRHKZp7CmmnKFz46pCnRm0vYwiZlWZJpt
ULEv+yltLLzHSKvHunK+1W3yn3mF3QWJ2949gdEB040ov56OhE23qEaZrF/Phps2
vcrvV9PaXaCHeg+NIiRuARnDlwIMq56P/svZ1cnKOiM=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 15008)
bCKKLnUPxKDryrXarxhnprRCKcNbGULHr0GFtOJWRmEoj74GDI0uZp6V7gaKySkJ
P/C0Oep2Hpp/nnRw+D/QOEFUB3N3n7Bg8vWwZ/YIvZtOfc9WS6BT3QSkFYyyHJL3
es3MUcJxulhQkmYZ5TkJD8fyUvLh83TYWgBZdMvwFYi9JH/IB4ocbpSvBzkDu4+M
A/BgsecxZAxmgWVjP3Qe3rvwGiiMPCXfbFqL7xg+tOKwH3Jhq/cJtgcGQVyWqZO3
hkYtd3sqIeYLCAK6TwhfYoXstLigY1+RD+WtW+bUXg4Mu3Ry58SmwXNZS4iejfpC
/s3Ix8zZwNYpsjCiDHoB4pme8Vgc7N6x9VegmflO2/EeZpBlVsiEcR8Ne35Gb9Lk
2GK/ExidGD+zg8b1nBq5JKl0s0yyXfJsro/3jxGSAu7H6mg68j/8+QPBA4noehTx
u7NmLUIYnEwcSDiUqrrVe9QGX581bIqCsukJxQkTAbN4NxkxcueEqVoBUaYZODns
Y7shcJfkUQtruXAeZIaRjwdqOemWTgOq2nZtAumhvlhF0mqqJEMENHbrKPpenMzZ
UwFC1dJK+bw/+cUghFGs/wIB6RMeVt4plz3k1RuDFmwo2Tj3+CXUiHOlBwxpNoIx
h8xzTecB0bIzNj7VMDwOxxkBDLEZLf249eFahuw2fWwrSgE+xaU6b2Pd3XtTx6QE
g+GQ4ONjiAm1dtvvQ8OOcJ1rLD6Ga2SBaO4b2FhZYqhku+c8QrbZxKvkpYpf1Dbn
LraSIf1jyVtM9xgeg0QCyp9uRCdIoJ2i1a9OOXaCYdBSrDE3LzzN5JjGw8JAqQMK
7qawDPEgnoX18xsUZXSdeHl8jUqExafj+GV2Z9ffuu6K3JXSX4T0yHVzpNpiJdKP
o31ZiUooDtNBmCPTrdakYhgMNJv6986ggPRDxIIxBLOIBeSJFU/LNs/e4qWvNeWO
qkFcQFn/woeERFvJEHrg78xR07NOP/A6eqpHf52Ce46VEv1W4H7lo7cR4Qrp3zi3
r4YGwUQEVrkjtiVUEw2QyxINuXbneSTfJDNjA6c/oeFpbmkK20Vj79ZXjTNHOVXb
LsPAN8QBcRT6X6/6tE5Dw1SrhSO+Hra4hXHNoky2mgMEeDjQoS0JiuahE36IDocG
bD1FuFGqoov6Nws/2iX5v4evQwQeR2sybzYa9Mg86cGgH9x8qV3iEdwRBIm0FzyE
tOr88DY5Cli6W9VhzTdNfCMioH/ElI9ZT715RCP+AS4zbeWECNln8qqNFbtNeME0
YPt1PTi6nk0TYU0kqpWUetNsNgOlsdj0/ecLTdheeqIg8B2WPZUce3l3Hw5SRmS/
ShsfNgFuzLaTXBmLX3t+zcb3KONJTxCNMKe4G+PBVe+nlNVq+ifUOVKq7cSc2kmZ
hCvst7H9FpZqUErf6RY0N8zO1UF+4hmN0zEK3+cLdMGsx2qOG2o5BeQx5Z1laGeH
jPzQBt/4Yw6OFLe1yk0VHFMbbrlDIDxIZOOxV9RDNmlahrC6Lq1Ir16XLfNAe6gh
BvIPZ89zJFDiLjCcw7JTkZF+4God/B42A6dVPuMvxu8Dy9mrXsNziMuVTyl12V/B
hUfraUpExO/Ktg9+SPTb/YwfZzNf8ThCbLphpGzXNaQXzaAXbGGswXlFwiRBs0vP
FITQbmqWvwSNRyMo6AwCirhNCngYJaWIkg9WCIDvn4KTQ2npHXhrNA2iRX3G4d6y
rgkltaO16ct+7icYXjzTPxD5a74yJtGeClE7zBxpkzlvm7zc9AFYeYxNS8FeRtZe
YGdKXTkYLaczjeapFOxLopJHeSAqAK0gV6YCYmyQxviK2kVFIq9fe135yztosJnk
qWnT+d7/Fn1aWRjUjMQnfD9aO9Xn/7Ho0m4Lcx7A+7bESOdb2cxMbELNgg/4ALPY
3zpmObEt3dQzWliGN47fNUiG/EQsALaOudSc5gG/AxTgZojoM1G8Bi3181TpwW0w
NnQS/xZe8saK8R4Yj2PHru7DlqVnyTwnm5vGztE4u3TMmQpfqBQcYHLxJGM7gvjv
Xqfj2KMcN5mrcW5vbxpb+W4vmJneag4ZVuGr6qpEPya36nH/nHurED+aPLKQu3Jz
AoRPRPccWlt6zERLW1es2viiYV+4/BeXf808gjOeQyf3AUoNNoUfSD2f6QR1N15G
UO78HO68WX8fdGL9JX1Hcvr7jBCw6FQmYpyY+OtbmlN32gYUrhUNC2uV0uXBbAiK
lkeGWiytCM1S2yRIJJ/TPA4GjL4zwhGXkGUitSiJwnaIQ71tpEEe28ZFL+hxNUhA
FsJlawmLCcT/44gchIS06JaUt8AyrqEmGlJhiG8PC3sSEypyEFoyjAuXv0VMgeDM
nA7kWs7PB3l8Zua9OAVT909vFcsIP/VJzcMRnnSuWcaATi2IHSe+BtIi02HDv4W7
CeI0K1CsyvXd3S2R/xWHT3zD7GEfHyK/h+JuNT92JFv0NUKbfYDzHnhCGiOHmZJp
5ppj5O3MLWNPdaSOsBQ3nHCbiz19h30E5kt9fhdAjwyoFYDghuPxIO6U2kW1B2Ti
rlZnlSKjsbS4BSMrkfA4pXQ71WHqSz6GMuBtLi5DLBJwHCYm+osO0arO2kXv6fCb
4ibgqW6SsD0hSaYDW8zFGcuJdkwbQ19tvU0h6YYXnC0rJUq6+joDM9gMgEkoWooa
abpz2IXacH3KAqu7+ta99eS2AMASs2lyFgNXVmIxYGcjdScEMpBzFlEkHwy6dzKw
RMG3ULVKqF1fjX+aIFF+k/nPA9C8WnfzB2By6dHGtDo5z/B7kHE5v+JzKvUuwdmM
O/n5UqhyC3qlTmGlc1coOciqJNdp/2ouHnG+Tr0ob9u+n79/2Ww0izDIwiGMlZRL
jRcjQst7Fjs8fd9xQN3IdApRt1E4scadlcA3Xi+CMSEMsIzWc37vLYpDDdUPH17p
cSfGr3VWAmCBtDVDpTIK3+ccr2BvLBClPi97Rm/DGesfUGHdWQvhdcP0WRPBILpb
rzfbtX8TC5ZQfnCrwshbweNniXwi07s6boBe2z4NDhoaA4VSSfuMKLG1PgTc1bkO
eFH65fOI1jA9Br7SSurs9i3+ZT/mvWSIy0BcB9fn8lJ7r3mCMDZ7UYlm4xdORn46
TC8s5uKRdtecoOBNzQXSfiFFKpWFGweWjXbjZpFlyB3Uo7EsBvirAWdRXrmnULv/
5aig43lEcuqD/yjTUrY/7blbv+sEjcnd7eLcB1LFQmEnxBvXiaqrGhdCBz/GC9i7
KB77bH/6kqjf13EJ7TQMoKeV/2B3HOD+iGq9aL9BcgdKcxFo8dyQKSnwVXfSG1q8
VYMeXiV+t6gooLTjdepRDqwT/MOW9TKH+UBEmymKw3eRvdfNMAK6c/hKCRz8QSKX
S1oNX5HLGXvsFNssSvhX9T2Uhw0rIrhSEbvIi2uax/quuZQs+2IdOqdJhgQ9R14/
sPPeyUWlnWjdVhFdxvfmz0+9iWE5MzgTVcL/E4IFTTW89rLSsoTqjpuZZwE/5UFw
SHV/S8QFFP8VOiffzxpi1oJvSOtSsxuyUXxA6GmqrzVEscUobgPj2oJ0FzlnsGEz
g28G0vOPdapfgMVZmWjws0drGBrWWadlQqQL0EO35SiOUvhbauiYcBTnW+1F54v9
KoVOp7MtfBu4VpIL1sdh7YY9/EwEP0WALySDDTvBLf9Qk9x38L46j2ZqhOALI1Qn
wNlAGtL3WH2r0Mp1Z53Y7BZuXSslOtIrFwoIVq8uibhzMAZEUE6BseaRjpmMPHY0
pj1tPTfYmesS5S1iddJw2KnHpIoazXGZXfdZ9xZRKgrtHmj/3sfDNyN+Bu31o7G2
cg5EWxGknlqGRuqdbUyoWB7D33nEogjfMDRJO8u0YOpamJ9wg3mAQ2xNHkZf+ZN8
VFt+XOfh39rc42omPhJrSJVJzW+qdDt+yHkRS45bD2lFn6qKMBW5iY0C1y8ZSClA
hXR6pq1DxvBTzZPH6n+n3VmFGK6daBzIoffdsYnB23pUIB5Ap+3OGdj+RBaVJBuI
a2eHkZFnYBXVEOk+MpPRdrjjH3VfKUKzK7sCqXMbl5hjcxR6XoKeZ/l/LGWFcqdM
oLTJKDYve/57pv6B3xl/6Cg51NVtUqCcUy2Llr07tP73QJkN8PLZVorAbDd9/apU
f89afB+noJ211xkO3wMBrRZjXBPZmgxUO4190aZuthRxKz+OL6qUML6zHCP1YYVR
5cHFdS2djzB8KkOc4Ctfcq7fVl3JOfFq4jFweij3WuEfQIvOJSE7CVS2xs930Jxx
m4SaqnGKsyIry12z94RvS55CkKEQkZUg7ZfkratHuD8qQxYZN2ECqesnPWfKqyeU
N60zg88A1y8NDnK0OM11BEJRzVIU+DLjhOtduuMOn1Knd7N0JIdSzKWy9QESZlDF
uzt2HWf4FednX7nPdIcK8KlCtmqbn4YjkO6GwgvnkscP9yPAnITK7ht8JseIOLUc
cU7t6Nwbv/DvRKjcllwrwI7ZouwdiE0Q29R9JmbpeavOxd0LaG4wG6EhafoFrjua
Ztqva8KKhJKU96aqeWXU0qQD6M+gHmddsq5DDbrzNVQcaFgS2xu8+RlTGMW8D7aY
NmmBMi+D781aMH6wnpC0AInPMB13ALTwNz08wTXOOP5CgIF5yiFEP8CQghBm8nLb
v//NpMfSDYT69xmrENefNrB5Pzn4uzQjbkvz0WBOZbuHj1KoRXRc55IK7YWuokjI
4eR3369NJ8zavxYu+RRBEdVShVKhQRfrVew7uLySY3FCjILwd30vapg+AoNsSYTp
Qk9mYj5pS2rABX5lhJqdqz4Xiu/a3uy1Aw5JYvYV2Nf23F7mI//6eSDfnbZDFAoW
4bIeCl12f5u3cOFEvi2cXAgSnPIqyjAYaw7z699TTi6T0KyEfGiOH71dQWjAbfRq
yzGipU/B3fBX6t/T+E2miA5Ed1pY4Hem5O1VReJabVEK/rbGr9qe5j0AfxmtR+kl
vMFzHb6nEt5BGAH+cvlvfueDizbWTD+QQYj9HikObtO9zb0MeXk25xvmgxpikTWD
xeEeXDe1+wGUZrxdLLK7wbfNePJKfU3NBtc1mwvNbnzsBS0E33U7YkGPUsMarUSI
6w6ZPHrIJd9fWmsFGNihACnAuMB26aYBsQrSUyqaskiwhbX8OsAEG5W0F+5achi0
aJinMMC8CH5kgiJzNz3Vgsl1zasFpj5Y8QmAx569PiurMLZR6uc5kpG+ryYLatHa
LWaRZ0/MBOZeJO+v+RwrzqIplw20IxiuE5KiYCkeu3STzS181IAzgEUkFmTClVcc
M/fBfUOuuh6lRS/gGBA/yLy/NLvVKn/O861+EQZkaO+CMJdu1wl45yxyQUCbA1+j
C8yYVhwQzSAyTgqgi5CyatnjxHGM1hc1OTY7LMGYnTQ2DnT/8TSjTLHinRjWJcoc
d+SboVJR/TIQf3oJHVlNaBWxUDz01aaphQNMQB9MowxgUcmvSVS1hchGj2PBwXu6
LMzofoJCSHR6sGZDSREBdGwXjCSN2k7k9bgGBE8yhHm6Qi2BfzimyLl+4+E+xMvy
sA6aYYiAAlUZcmDMuTwZt4A9Gvyd1TaZHlXlNo7bHy8zJpvGhODhULQCCNUFbL4a
14pgHZLwZ9ptvMvoWb4TS9zwLgNTeVNYn7iVPKiTOxCIR1ZJgq2OcqwysxlXfMeH
YXkOnNxndBFB0QSlWjbTBmnEJxQYG+hJURCjRBQgXj5EumtBMFB3RbB1KvYM4/Ai
33/oRVjSwOKANLm0ftXdvsBSo4N+Wf47nhywbsVyG09aSvjGMdLVJXqDl7X0p0Z2
uGABmV+z8+bB+ZeyuI4fOGlhvgfpLegmPUNUHloqrPIV0pVVJesN2k6OGGeDP7qm
pE0HC3hHa9m/5q6JK3vuuOmXfDXrdzwKQ+ovqXQ2O+ykGmk2izWWALJ8IRnX9QoG
Uz5gFQ4a5rMsoygjuJHylhQOdwyC269oRpK5/eVQ8SZ9K6vliTfkO3YEDbSB41SX
F+P0tonLGSI2xnNhr+4tHxklWH4vjR5RTH3C7oFY0WmVrNyr4GzzVN+7uKCwK8ls
FoJYMyEj4IQz0cHwIXofQfqa040jGBloolZrImwlH5uMSrLi6S2tmTJl73i63xvg
EpydWAIGI1gNzD9k0+eH5CS2DRJVxGCgZye1NcLEQV8bwfE7wKNqWbu++r6vmV7h
+Tmq/4tmJEWevUV6vsYliQIkg/VsiQqWOjIwy/CvrMAURzKDKu+Hfz7bo9NLJiyt
tfbJ4ShPt3vFf9qZ7E8YlACKy+p7YvhAG4FP9W0FZATTsp4VunCEoNv7XrH/F5l1
5zKiiGRuULW/p/B2Gs+rNqaJ2SvxaVYWauYmai7O5lv2iuz4tGvIEpd+4yVdsbHi
uzlBvwVH80EE61GEJV6yRZgXnFs3NKitwNMfO9+X4uMbYzPLVBiI6rQMKE/dZkjH
W2MGutREaqBir5uggukulNm+PG6f79VbPRNSIadmQT1on7/TvZOGwgzftlMnlk/2
hiujQVqNoA4M8M7QY2J5IglARgAB/BVsvAQIbBiHrv+lvTjdIpFGLKgnsGgMUCqx
zJPtbbq/GjRpejxU3GP0QHX273tYShEsMn8Njsl4kUWIKbPTY5YCm4iqzy1VOcRE
RsohxOyNjwCI/r/0dxPu232DOLehnc4cf+ivV029is61YajWq0UXmojjRKN+0u+Q
zvEa/7KLZrmYcJ+/7u11IQ97DesZG/lZcQYLGou6hYXNlR4yoeyKFwcr6Wj9ejQb
kGL7nIMXfM8Oh4APVEvljncav0sIVVPpvMAUOAfG3xMvoqu29oNQl1dnCFBgbSl8
QvUy7p5WO+1emUUqhSBoQdB8pRLLGlSC8+uSTTn5fYij6l3+4N5z9w+dGciPvoyh
+wRTn0XtZwSuYwymJ24iF1ZMufnBSCtC3u8DWteykgBvQyGHuZI+3mRtYRBMRQfm
DxvWs9cityi4t3kA13Vlj53DO9/4etmJLChnfdpjGN62UQ5elTMQJu9LAYm2WTsV
eyYyLb1NAe4e7ySO+XbzPdNILE/Z7KoPAJRlo39Bwg4C+4bj07fAewkJLzWf/Pzq
hxCScAyWvPqDK1NPY6ZvzsnR7/OBsFg4krpFt5ecYXyOUAmhDCkZ1YHFPMoqA7PH
r62dwO/REv+2kD0HWUrIPafLlkx82fb2bcpKZrSFbaMcahNNLaYdD908wNfZmHh0
rRr1OwCRD0GJqGf0S3s+7st7/r96q0KuxhmCeGGxL83nlqmU8CsmFSyb8ZQCnDoQ
twCcEpt6grOpHppegdY1JAG+mFCkBmJ5kCT7j6YoSWUqfIGyxTCfgNJteTjqPcZ4
rC9gBIJnaN2Xrt5CXd8/Vsc+RZVofjWioghp3Bp9iEl+Z1ztmy/WZ1cDKV+Swzmu
tfMkqwzzXfaybusXWC9azEJfj+90HMyayByOSN5ZNH5ECz/G0Z09ww/zqA5bCR6k
7us+6E1MiGOiIin3UxaIjF79cfXg/32b42MajusDq0o6socfqC1mkN1Ms4E/cOMM
QVgcibDQpJ4PHfzORXx4Fg9ZsGIY3DZ894m0Pdg4hnixAzuAruuIHET8S8+PJWm+
NGpCI8gMat5GAAGBJlc3d+otFiXCtVaSNJIf+F/D9QOMsiCBw6wRCSVv/sCwnl6N
kxu2DmfdxwJbq1IUKR8FC92KGQaplTaWW1oLmZmCZiuK9ujVql17PXi6mrSIg88/
mozkM8NaJ3LAtAnQvgbCGqHBT8L1SjNlQ6ey1qMmZGH9/poQKRmwT6eH3bE21+BI
0sPKvvEm249zY9WX8rjwrqq55xNkeEUBI1UCpNmeoZqXcj/qSjW2+Q2QHSF5dgEt
VBq7xY3fqt/1+9cMzo+qA0vV65g5M6ktt16Yb4rKenuyrYn/YZlrtvr7WrLVEaDN
/XUE3sWbe+5KPpVmuegtKHW5ULnz4pxzdOts4c3X96j7GlKmr6cZbVh3cMAWQx7v
pkX5P60S3cNAXKSEV/yANmrQsXRsWbSpG1kstHMkRiJMkcWyhyVoRK4aPDYTFJeC
z2Cc/K4H30K6O1Oulz7Nw4cMbuqLNwT0Ur5IQD6bUV/JyawjOyhx8LfPQZz7LXf1
DjpHsjBbM02/vBsLA7YCiJvegBTwm1wji7msCfT8wAT1R6oX+mGD96mi5shOdVU4
TpZAsygJq892wI8thPpExBh3RzNd0Yr2dAMuCi/xGBw5EtZRXc4dM5IulEFctsqs
BuYyU1X9GS3Tm9CyqkJbd+pRgarkMwdaNpneLZzJlgWEvaRfszEir0EP4LmUwSty
OsRYEzB6W6wcblespp1R4ZREsAkERwWQqOfGtZt6sT6AUScd9icprA1O9jhMx+3f
OfvrWwvvzB+rg0wBT12IXWaGqZQ2A/KvsVPJkwbbFJepDNi0C6YqjNQchDsIdQac
C2x3TlsxwzwoxZ4YuxGf9MEA3qTQEHNj3SW75PKUbJ1UAU15qx4qlIFPreOx6r/s
x8QiLoEfYVpuxbERA/SdWR2osRFTKQ1Gy38g8QSeqQY8JSZHEwxSQJDCSTRuPPMF
lHoE1Jog1M4r0UOqMcnli62eEgsmbF1SJi+ZK1bmDVwNuy1zYGnr7D/+mFz3m8sy
hGRq92MdlcxbdlwiR/Ycu50iIlMrNWS//ADDYB1FKk01SjRkQlFmGe4qso/32ZJV
TnD0KFnW5NAh09VxbcZdu0KDeY2QXHxT/wUo1gKMJj50+3bvXXjU0zaDKdia15hx
qy4HnM92DbQUB/0e0sv7TvW/nmwIsMzbEfKTi9XqFbKhWoc6MP+QXrYCyjgdQCj5
xJoDgCt5OMHoe79OCnXKI5YV3PJ/4QG84b7z03AiZb7fxoTsZmqvVdZK2O9VPWS0
s5Rq6bZxNcIYPgiDu7OvBEhxC4lEwgvZHR/y6r0jm/Qatn9wqtzsNwW9Mtihvhab
S9t0lDZ6LPm8S72YXRw2+zGE/vv/WaN/IN4fWiuLjfLXfdcan5lXEVZHAyICP/oN
3gSk9jJBC5K2JFNIbFCyGf4wOOYeHo5fyE37u8ie+ZQh61J8d05gzvZ9anGiz+mW
tBVtR8xxl/6B6nwjQViiJJFYYqQs7AKJkIy/+cK/fwvhMsHxmz/GX0UQ1/bKyRQ1
7M85tb+neKcP/VSnkl7dif6A+VdzqHjFcDqkXnObp9kI/t+oPi6Kh8WmagA9jDvd
KouaFyz3vHi1Q17/UfBW0d+SkVOUP9KKSUDo97f9TdqE8+sncenfnhLpOsoKQ602
8guNj7sN8lnj7xPFHMDE2iyNQVlc6F++N+RlmpjKNhcahk/l/XmSpm4nVY472Qyt
HfTvuJP5ppvullKHHVz8BYx5OII/YYYToDWXEFZHwuJxlaJbky7iwrcsxKWudTGv
iE5zjdJ16osH+33nxzlxw2XV4ldgpiKJCCXieveGPHc+WL+fVEJlq6XmlTJwG/rI
cSkxZOlQOs31CB7ecwVqxNWL7V1khZ0WYoGNm9SaqJaIlW6dktmwtCDwq2UH3bGF
xgb2byBqqnIqYiq3Dp19gRoBirbyuMT0RIr4vdqLdXJWqrHF9jrt/w+NF/42TGsw
psie8MmyjYZeqp4cLbg0Ne3WqaYDboh9EpNaAWllPqFiBxCs782NyDeYn7K1AMOu
V+GNNxb/oN4A25MlbRWfMFkb87/KIRYXOei9VWRhgQ2CdELOuh7KL2WEVaDPMK+G
88ascy2dew3jHd7LB8zVxSqdncWfYtA0oy5A7NA3iJkJ93wjz2Hov0REv/2braxH
1l8DlRTuKgaak+QqMCKwy1At6zbuXUHWAJUSC3a64Qn/q8s1sQw6WNEY0seJYsDR
qQJ6vVa1YqvtNRoHtV73vlJEGX1cNxBejBh46sXuJQ+C0iHtXUSldjhhK9hYxBvR
t7iJH+3DWByCsu+YF2IEELI4L5mJccJJt1XaYyrz+2NX9A2gFKjxRcqQH8jAtOOz
6v/e4y8UDCGZ6RRyDIOVsa+wtfRwZB5PKGV/pALTpeNPtaEcYYPoNxV/B4LSTOGt
lwXjXBi2/sGY29Dm/baLqjdreTPlwlN3lGEodrzPwjpetedMYBGALoB5Hh72DZam
P/Eg0DNgM+KwiFghlIVjoH22dK2TEup5m8OAQHIFDfUIzBJ362daxS7QZnIvlhv6
rJpm6qMTQCC3a5DKEysCnb5tWZuQieUBMj8NsuWaMlgd6Fh/GJoDkjWcA3uHb7Wd
Oe5n/jNZV1HWtc2v/jLW7cBNy3g8ozIFU+3lM+Wsq3oANu/Qn5hrDIwE71t5f56v
sqXDK9IeZvoZVl3HPz1c+UBGrNESiJ86yNSmyDuz3IBbNMGdMybThjske0/+c/K0
zi9YA8SfOj/HfVMtEVXQ9W4Zs4c3R8W5PA0dZcgJNISfRP9vUWReyyfpWuH98Qs7
XQ97sBgYfI5FNy4ekQUqHTvLLhykd/otoRGsEmsSmf3EtKxD5H5M+YvmKezXB0PQ
i8QCbgh3JZ4RzKvzvQRmnEuPYWNni8QGn4JtpAwAyKd753ShfDV/UJsUpvJN9E/r
PXhyTl/TNRJ9pgXFK9MdGJy+TuCBUm3o4rCG+jnlNOgosGK2hYy55bUxPcC/qGC0
tCu92sD2HjrvQjl2wWWopXBRcYUgSKF2d05/0CQFe8YNrfSY4v490VkSIXq67fd9
Ca1LPZ9Zc9jxv899HyBfQeqW1uwSnW/VQRbGXrIvYpHJeW22VtYACX/RERojwK5M
OmzlTZJQIhIMR62rOOB1C4RW0TZds5uK3t3FZLLCX6ToPsyPEWZcsCQiVmpXxdKM
RoV4FUVPXlsoLDtCrMlBulDy+IAlm59lTWIglPCdvuxzXh0PYZoE4kaLyPyTqZGR
ISJI5rASd2Hkn1P7Egl14YwxP80bfcXO9omKVh9D81xwtIFSDgOQ5bU6qc+8Dl1k
cIhNYy8RgerPnn/wMcMRWdpNU/39z9TLMoQZsqktxipjl7whgMFKZ0/QRaok5xxw
eS5L5vZOkUbcJ6Q1O/pNhbUGBLM45bhmiAlsNCa0V5h5X6zFZXx4CjXu34o6HKo3
N4U7IBiF6LUzoE4NajqjdzPxq5zkrvhhp8xKE5T0FPSaI70rA5KTH0RNUoVTC3cL
C6HiN7NRYq8nNZBcHifDnXd7Bmz6y3hfZnyRcV5/nfWbHiJA6VItJMtdnEFT0Spl
l9WbComKAitPiU3iSxe6nm9DWi/XvRm8BugCnsm30VGMkalpsv2M+PHzv8PKY49c
jo6/V6ZgODKD1yrWG1n6hAbC+Xva5l3zGCu9OYLC7j5i1tt5qZUJEvn4PPusLH7y
2h3SJ95Hjqr47ZA7GYAGeiG5+KZgLLkm8SO1Ywt1CK2GOXMISFvk3bEPSuzbiwdV
mQ7BAikxE17UToQ1pek8/x5Uyb88r0dgsTtXFECgxuSVIxNYrAjA76Dx7aXw/d2Z
tjqVo+1XKoqnDhOTQMqVhAFxUuGDFqklp3emNN+34DXXYdpJl+lT91I22433D90I
hQ96D/8B4SHHElCR+3gbkyEuDOmNRu7qlmSGy7+VZizGZRBw/JMTy5lRGvogStm9
TN6xQ183QOF1Pd+1dGA1DNGhZ9ix2dWvAw1mLtMSiPl0eS+uOS1HmCIIwCBKTgDH
7UXFs7kQrB9yU4h4imAF37USgnkpJeSyg2xZEKqMeRVsHahx+g6DgsgQ9OkvEsxh
YsKQjGEfM1bQCTwOsR4AHiOd5GszhB3FAnvXllaNFN10KcoKioColwVVfI/H86PR
5n+maVxgEeS6lbMVDh1gf6+AtJYtMfccZIUS4lcZ7aA7Tp0/kr99o6pJPY0+BIhN
pCkFyN1utqOXiCydjJrQBSMT/Lkzf+Xz1bwp/nUbdjAyGa0FVZBaYs9qOMH9vzhn
gC/pHUHXJ89liqD1MuGmXZHE9xcV1X+N8lk+RLcagFbhnzSMAieGMdShat6qFOKG
8ULPkiLiY/g8MFjs1TGaNgwBnG7gHdnA9RknX+Mu7jO9kNUALeqbGFcJfgIj5Tpk
Bgxg9QS+4UY91zCLsIghKjb/s6SLS4UMGkMDxKheFO9ev61/srBep7lcI+KNIkm9
v6YaVUFPBUZ72TTbR+Ij8duA490vEnYCkUwO5CgDcrL6365WzJHpspAVjB3db3a9
tMj4o9szBwEHhmjK2Zy6LVZpg9QRnQGm7y3/1BiiNKyigSyyYLbKs3KCVcXIYctq
W6CTIiIR/3GdUw+L3noOTGaMJZt1jzB/b6zdKUhVMBhdE2+ZWdOgolhyau/MwQ1S
3YWdXrNe/hitE4MnYXc7Ly1ePHeNi85+fqIMZDbMCDrczPgnrFQQjJIBbkfHVKxq
65qw3NjEFMYHCdo2opHSiNCTUAzDZgVtMqBs8NQFamuwg2KhFoGE0Y/M+QLCF4Wj
/wO+rsFDZ/ywdT1nBGn9Ypt6VpWbI7EDDFUymqvADSTjclcM74i+aMwNezx/yRHx
hxNl9SqsLY1PVJvgWpUwCNMRBpjeqvKIOXrolHwU2An086m7UF3I2OzbPm/zBaLq
2ZxIofWRrG/+zSEE+H2y/oy1JuPxcSHhapZC/ddK41lKVP/Z0t8GaOvWBQM7tt3E
29mPgavqNwK4Tryys5FcfVE7FjVI9+rWDX3QFoRzUY6z6/gCFQRL87+QNOFk1hko
HkoYgvPLlkGmbY9AZ/8UWSPuKDDDmbBgAXY2nnwpgcKOFMtqDrRzQDy4RlqjxXU8
2JFWIIOfG24DvcUEZ1oUP7ik9QqBdU/nabolIqv0vDQyrJlKhzEYriJcYaFU8RTO
5trzhNa5/LahUUp2mUsfD36RWg+p2Sk17ul95yP+yiKjRR+Ewa9Ez5JORgTb0wUV
/3Q9fZpQTXQwnVejKfV8ZdEpV9nmP7CEQa60C+VKeVGGJ4a2M8HPOnW1aKkGZXKl
jCyD26jws+Nt18netSr4VTSDzxJG/RNTgf4hox7RWgOkEQnec4QMx6uT0UKCsmyK
flHdFJ6c5ZF5hvohXCybuN6HJZ22adqju8zY/GnmYf4mU5ynUHIWjeKwdxCk7VyU
PDEJOZDix1BgbQh/C7Jj7Oc40uA8MBc+uMiwy7bVs23ycIFtNVfHPtftsNXweXdJ
SchkfUZ3a8GZTBqLPS6TsK/FilQQXHGg4U3lliq9YPEcVF4OjEKzJLTM5GdRCFn+
ugXQzMdqfnr3rUCbqvYRCbeSIwibqyJJ5v19kJi3KTlfM62aH77dZASqqxi/wLQ/
BMy0jaVcL0N5V7oDEsURmjS9QdDEDlpDEFK6pOfTpK62nnOjgsAth4nL/p5lNH/g
sZQDBls07wt47Q9stpYsjkI3Oef5VNZOl5V6+SSasN/6lfe3Tqri7QeLNpk9TCpU
lViB7i6/qlOtOnXHl1szwfEz19OgHhv8Y37pmubdImIakJ1X47+6M2AkT2ZVND5K
vZV7HoVlokd6PZp4QZSh3sXjs1lrXe4Fh3eptQfvV4zHgnI++gMgP52UVzJKDBKV
Y20SHQkCqIeTo3CDwN6FmMpQVtD5N8bu4qSY9e55N1DALYJZClBxGjnEbqk+Bouc
3QuyaZWalX5xi+LpJ9ddbEjdYKedTBQ5UNcEjla8ZhM+8GDWrkrvvyYZOkdUNGJE
ORuNgGHKGmlNW3EJq0hKnlADFTo4p5JKnLjP5mcOCoAvwoh2wFq8xH6xYAtFh/xC
SGjrQ72PVEoMJup0WXUMkRInRdNmGQNg2iS78+imyEAHnjeroW2eok7UOFEQW7dv
keW/o+OmPpl5fREykaqs1olDoz0QujJsx/QQ1WwLUaYpC6veMK4Nfqmw2USH3chA
fA80YdtrSWlaXYXSwSaD4Lu+uf4KUAFl5vNg9Y01B+veD6bOETYOydbJbcrMTasB
gRYEfwsuR+RBTXqayWJYReOHvVlmhiIv9wh13gSGw2XUWrcDkvvpdpdWJfYq/egY
I7eFrLf7HI80pqwOYzM26djUAGYDRfGiPVRy/M8Jk5KEGfniCTa4Uv58vTeGepbJ
JYQXpooQEOStdg17Xo5z7Yda+LZ1Lj7CmBiGyAmFq2vI/tunKB877P2laP5IUGWd
7spZ38jBSAr1LGmktEqYw/TMKtYAEsysa7QdK9pBpZSB6eKW8MLS4QD5E2E3qgUS
BDj9D0M+Vho28QbRo8XevwYq+Ug2y7PLgVd8Hxc1qgkePTuYrRnnQ0e2W3i1u0EV
0BuKXF1IVVADaT0FL+ZmkmZ/pWQuF+jtrGgtUN8/k6j+QngSt8+8IcCVKr9Cz8v7
wL3CiB8JlV21EVMt2mv18IOQGjt2IM+3hKWkrJnOsaatmw2jn3au1XGpCfT09evS
2zyYqmv24OvN6htYlWxzTt9Z8NpR3GUzeRt6B1QdZgD2Cj0sScswEaWeO6Ogx5FP
tnTBqlOffkXKx3zgKeS21UzdWRz3p0uB0VHRjwL7DOhhyHYBuUP7ZeV5sdNTXpji
Kg9bGbkron+Ev5dQBR7Fq6p8juR9fjtgscS8+VS3w22NuvhSnA2THo2FHyTOaLhF
qQALqHj/iu3nZT3NJWVcS0YNP/K+2Uq1/THAaF7JUl1X0KdQN/BGLPvtY4jusrfn
GxIRLOnwvv6xdQQkq7S+7n0sbZ17m5J9wWoUvVWJADIvm9e4pxnOZbzIwIEc9CyH
IFreD8g/YxrG7OiS/1SUVYttHg5KflDOxOUvr1gEv1K8HpPjUOfjZjK96JdWqdfO
Xdkj0s4gkkhV30U5SN+XP/EK/BwtPgf0/jt+aLvhlHdduDRsZkmbtSn9PXolia8G
FXbdW89fsQcnvziOGJtsi+FeKNURqn+H32Ug/XMc5rolzq2EF50ap4nGe9Z/2PC7
7xaGBLJuI+VbvXrQZo9JJi0FtZDX+Ri4qXzKapXWgUavuMuJO8cNmRiNit66W8IF
l/ArmLLqmt6ncIMhyCJzuK9FGdB0vhY5LvC1zkWR0NS+veOeo/67UyRB4W7DPziN
Xphep9PMWSksB61ffu8UlK7s9kjNTj8+y3dvd7D6stNHtq5JHaB8f+kB/DFGLCSF
1O01GZB+PQBd9oY3KQL0vIrrD8aFpGZYXe0j8vbeSNyf0X2gg5m2uKm2JQpHj4OF
MRpePuZjim75gKdvVP8LQ6p/Zl3xHZZylnA0Wwv/2WS1OU+5sPGlIc3iQcIm1Y29
uttexjGeBiNug+kIH+ZgzDux39hJwdndbzB0tMmfOUoofXemEm3g9JBxcblY45eE
+sauw9f/fYY7KACn9Q9jZbjZFadpZO2NDnB51dyeg1RraHfG/DIjBrwhVer0NU34
rZFNCx+kbBg/hj4ac26zeyo253iAG0AILpEs4lzGLFTClsqkW0KrK4p6NQa+iewL
mEUHEFPaWLRtoP72pPDRcVM5mt5JqiAHEd1zX9FWMrkM296Bzo+pE97YLpMGwyE+
KqmOfmI3bn9ezc2nExAzGnbIq+mxWrTckk2qVgWy7C8m/owTRQ/efnRZWhAKfCH2
PNSVJ3I03c7qOLPuraPzCVcvBa1DxBmda7KgHKBG0/tQT3Vu18CEAGKbFHwAQuDe
KvLKlqttql3DThyCJ18pHM0PhGQAZ1W7VvNbWmVBGAnEi7HMvdNCswb4g+xnUprP
1dU5dQTN1oXNf8AuedeMjrtug5vKycX/2eSo6sdkAH7J0ErWHIrK0W9S0He3SoBH
Jv+BnL7ebIhBABJVtWUKroBOiXSs1FOtKG5XZ6oyRCXidFZsOrqofU0ZNQMMyQwP
Z0PGAp5i6hBkysMcjcAIy9+Dr6hP+hltzXwUZdmbNWBW3nNcSQBcjETZOq+FNnbc
RT6rH2gOBnNT0z5/oTF1ky5oho1aKP8DWnaw8GORh1NbFgH0jh+E4eZbwsN1Z0ZB
zqem5TWnZ1bruEGiWhHN2JrnY8vJRPqnl6xo5Sk3mXdTDVNw49f9xYTCIdt8SOAR
OdvAHxKatSoSbinH3kTgce/BiUEg+tSMjge1/jsJ/6BEZ4X2cVTB8pF+LLqLM7jK
6QeP8UFaAK9QTtJg/o29BpnIXMaCTLPwNtgqX7cfzoicfvXfv994l9gd/VnwK34c
4L0zgpq8o7ABwmPw+f6igKdu9Nuxzs7N3Nzm1RhgleDMvOXDCGsgyX1Bv9cYt7S3
8nLn6+/v8C76oxga5F4s7nCvh1SiIq1ASniRIwthpIJCdecuDQ65it2bTiQdlfRS
APanZN48gNY4uz2BuFx17iMZIQQf7T1np4NkMB4bTZyOPTCFRHrAzT0fogUI0BcU
vWWPEFicrKhT+YqO+y7+dPu9wLW0CT2ELlo7WK7zOFgrFhg35Dthdl721MajiCzF
pIH4uudHnwLrvHcpMmfsaSwbagIr/DxCoLSV7LxaKDt01NgfU67oqYuLoyQD7kCR
iwXnn37PzLGZ1KdwGv9LbyJJv7FrDP1QdLUTMsn5eQ4xiy+3y8FbN2EPH0d5ryH8
oQsx81EzP6ELhO9HQbfi9aUvOOgaE6z0+5H6D320iAD9B268h6cpZ1ErzlqkIPjx
L3Szhae//92Qe51xfTINTKXGVTd8cZX3kRWVxMcc/OIzdUse6/NQq5byuKlBPotE
7kk6SyL5KSOHrwUaLC1uPRcJ1O71tBarZdNLpiquCSX6BYeY+GY/7KNou7n7X627
N4iNAH2+y1ThyHdV9Ji1ku8C5XJmUzhTtQGKWPjHM4xbNBWhUPni6x6HcbK3D/H1
yviwbAH1G7N8o6O+BFRUCkS+HtUTsWZ7FsAsnxEhc1lo07G5uovMOvPawsnQ0skB
tfMHucbx6ozQqtfIsN1PX357F458GR4M2928qayPxL0+YS5U5X3nzoSB4si6tmxk
HzS7XgoHkfZDMyyucPNq43DvPBfLuPBFHCEpX4mPJOIdOpbgj/Vepeuo4yl1lRgT
lpmNWlwQ6b09fvKLWY+en8kqLLaPOhKVyU3EI54pl/Q1s/9d2cPQDxm1CZGo3Wlr
/9+zbQdSbCVW1hkOB6z5AqtlZFo/k3NO9g1PbPz3MUI3fgtVHOd86K7bpT6qyDaU
B3aMUA4X4Y/Nl6GWjsdr670PaRgxxfSwY6beunWfqkaatVtUW5KroM4xm8xkg02G
r7e2CMbKNrl3K9V5BibSwLvIuKjbzCvhtg/J232ZxiDLNamtTu2wYAqP1S+7Has5
Ur4liM90+DzSHx1yHk3F1oPrzBwytB+kWOYnkU9jG5hjG0KmoUdWptiXmO5A/1f2
mmnAXIGlfipyZQcFPphZIcawfnDdX6D7AtsKEjF1ekp8ZAn42Rz4FCEvdn5rak31
aJHY6HlU/dahgaNKDSXm6kR0CrxKWSTWNKHI3PQBSkRw2qoz2Z5wC1HlcGiVJ2Gd
2Iri/ZTMqoMIpn6FceT3VNUPkHshEvorJ842tE1FbxSuqDCAMNpC+BuKGn7Mb4jL
cEakx7iAtWDYE/NGXb5Cgdsqin4s0tv0tQLa6WWQaiRoIbeBPpsPYx5Kx15JLc3K
2az5ZA3+rHJrdwEt9gyZij/KcdCpxrD4ZngWA5VhmnWyfReLiUEKDNrmM0KPDD09
cfXpeWqDyl6LBffwTpsuhge8ObOv7vqQ1nvzwR/t/cCbHCBp6xJZr594y2YspOU7
0/fOGwCG9VhvvI6euI4qboBXHN7bIRSyhWvC2Qtrmpav3zMpwxDjS0FDxtsJVekS
0pTH4GRGKv7egww4DsDyKgxUB9Uq/+zDHU0awiG2kXCoSaT9wVz9IoeMLnAYYXOR
OvI2wmqL4rqYKV0DgRpxLcauotdRQT3k5wrOsbudsTIgJnMzvyDymwh0sYAbXQne
vShaAj9Cuk7RmFQz/ICzI/xwxWmR3Hvya3ErMgCmQugWyBSYTZlNl7cJohe/b5Dx
OpXw4sMLlh3yA0ZbsQnqMEQmf9OdnUh9PkJkXB4QhzpJos9NfSQ9gtYGc/NzjbVp
H2u2bgbp05zU9PUeXn8zH0v3ReAiSSydIeLBa9RDiw6t2sh5kMmPfoD6L0R4sTdd
a/vwbMADN+haKIxBtz/BNKJCQ0udmY9kIWRksjdz580oZnpmMVxZTzAZY1umSjHd
woU9pJ3GKW8XoNdtnxmws2YieAYcgC8LP5vIPmI1dqGjbAs87zgqPMVug/pJIKVx
qA8+IIPTv7zn+5IbDdrV+CG0glsG/uwXRZuTjFxhPxRrDs1SQGYSYN0vzW9P/bZH
rxyM9AHct2OlfhOn5KPrAFGTKyZpMQQC6m9B25FP5vFLpgcWulrTGV7Ffh/Y46mf
4KYp6U10Cs7mtNjl+WR0E2SqtsoJg8ZIdiZqXOCKpW3jNhmqWvR9Av+Dh1SkfmUf
3X1xsXnWVvKuboR1j7m9I8fQDpDE4a2lvOJ5XMAFuEb0Fez+YK1zlB34Scqqyl7C
hUPKUgbv8K65gCHM6l+NCADVxtGyQNPG+5jsW4ZosyL1YXQ2TjoQxa2aT6iWzV+K
aW64nP10duW/U0p7BHPTCD5PBbDo5cDLceBx9n3mBy7Wo1SiQ71N965E0d4KkdHx
e1Pul+GFEmc4M9OmPXxoOtvQ02L5Ze3LzfZmOAyG10VYeDi0cw6W3sXbM9KZTF4R
we7WAe5sPXHRAnxWKrURh0GHwFf/Sjoq2U6CnxpNv4XYVIPPq9FTJAIzfpMznkqM
gHaeOPFPpB5iEJPMTnONTFy1R5J4tTUVIz3e0uczWn1gl7l5fq6Mz3WWidM0+Cb9
/nQvCXreD421RJ+gYNpJIP78qW66+rez6ipLyacPkjMxrMg6Cd0uz/zeJazjGyKX
F7X15E9nPdF8mHc7vVy5qOsVtcA6036a0JKo9fewOJOVck/cqLbUMNN4f1jwIq1T
YufiDp5tnje+3NxPXh3JgQTNOsZ1VHYPUk/1p9Bfw8s0VkljhCWP/xUOjVChRyxR
KfFXEScqQ+Gn88U0RAl+enb7NHumbEEmknXDSR2ljlQHwz32igfmr376Ylmqwt6s
g4ui8SNBotBUUJvVrfui6uKo9oEHAXv53DtMq0UaFhVbbqSLbWfDzg0mozJOmEda
Ca3ZQbBp4nRjqw7wbYqLc5NjYi7UaBe2ey+l/zxA6kl5klsLDo2E6oIWwpBfCSMQ
6mQsAg7mdKTnFf4oYby7YRXMzX5vZZNzvthV0rLWG6ndBEj1J5/nOqE+TTIVVVRL
5Pw1AY8pgIoAgK/GBgi+m7O2zjN8VarInP4tm3ouvItb3zdiEqK69z8aUKy58zy8
lk6sG80e5HFic51Cks6ATwblCdJXgb/7axcVT/XM46UP38rD30bOTzoVrgNDf5b9
VGK8nVZG9TjNXiqXZu5+9zGXYlYRnPkQlPw5qJnAK0ynmY6rZogVI1gBjaHE6FRq
3AJrbmGxb9VZSiBcinnozDk/7Sl7rgb/KriHFOUpzotZiblDwl1i7XPP9g+gLXKz
5N02ZD2jfhFIKogeEiER5QLQMtthOXU6lGdQew7aSQv58XVsyq7VQ7UTDgidVVVx
QqOZS50HMku9o9FFnwPwgDUOLmFaMXb4nOPNVLtM+J2pJfBKR2468OcuhVxW5jzp
bCYDxCTknDW/a9mqlqCtvejBH85bKJoTMqakfdDKYhunryvkJKhwQw2c7HIhEALy
+T49TJrP9aa68EA7FkQF/oT+8wC8LaPM7ihbR4V2kuYyXLx96KWPW+x0/IDF3wH4
dzR+VxixyoDleuT3lPxzhccHe+lLcvqHKRsJwmnioJxhF9E5gmBpxIXi57iuRHq2
yug6oN0q+pqjRZD6TsFTtYgVl05MXQhopPWWulptIBjtUpCh9xByDP7GRmBOB2/H
6QmhvO9qK5Zgy7RCKkqpXrF/yHsdBZ2yWaQcPkJ7Vr9B1/INhGDo4J57poDId83i
yDEZbZwX+vHHmUBL40k1oeG7LKjPBWNBQbVqJQ03+3yuiR+1MAd3CXYzuYyK4Uav
PLLmYv4KY/TB3C7k38+Zi4bUx7xMlWS8V2geYrFMnmSzGBWvFhUEC5Yhs77Dz8CZ
3xyIXmgYR0MN02IPGoSGt94DrwNDnub5mAkwhkbB5ns=
`pragma protect end_protected
