// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
JsjEWWZe5zLNJmHGaMme7whD0aRwvcCGbg0XzhmkghcZLMa9TG3E6o2JHLvcfQistTVr2h7JS5Ov
fDVGDCMqu579NCABPDpVu92/10ksCkn1qqUQS/7b51Fhp6weNF0yFZQ55wIKHd6pe28rcUkFEFKJ
pQUfDZXw99qjpYS2vq+W2zdS0zlQCpiDYE/T0dB4qPRInlcLhuEteYCovX2oKKB7z1UOUeSsK9GM
gjWK78jS1n8KsLEuSvrnOXVkvlC9cYy6gze6I/uJtRRVDzh6x3a4r0ucVHRUoStsJy8aBUVOtIuw
wBOFadwHfTSyyNrNAPBGCtvYBXVQICeTu+VWYg==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
N7+cxh6U9lIbyK37fYZoYUoj45o3d2nrWMlRJ4Caftbng7mU6yv73/wzYSDnDn0p9pTAfbZobGP2
3VV0tdTGHtej3QOxA5ehsydI/Y7df3IOv9zDxsfun1L553hjalnrBEB5sQp4T8D+MBSFDHCpPdE1
CjqFDjKmBZXe9Tm1s++6Kxk97FgGdEUIqq5rZA8oGWe17bJ2N+mchwgIW3+hJC7F1/CqwOTloag5
bOUPDH3+OLrF29B09kXpv7evvUD9lqu4gvJlXniuFMgXpqEcDf/22mBjIQZZz1ycCtltZR6bcyz7
2S40vYKdXyxm5Mt0rGtxeJIiMSdrsuBIOPnh+IgqZYyAFN4EYzbF/rYocZldqUhBCPpIEVNE3oYT
yQUKTCdGeARkdkDJVsDV/vOQYg+ztyt0uDuhxEEpmup8/YOeRwKZLNM5D8Is0yk7ySylxsL94sR5
WmTWM1mVS2QB90b715lc7yEZ8l1gD4cUgMAFhMEOde+DpPrCXpOxwCTlGzfMflRfFKOZrfH5lwt8
lwqQ4GmW8tXQbQSRRcnng/K1wb576v/jqZ1mD7Xr8E925oKzF64D6PkmxrBUCTVvkew0Upxiv4Nz
ibSsRXwYOjPRO1FICArKcqfOcjfnGwOc11z7ySW7sf6BlocqvogXeUDIVXxfjcPtU+h6jxjLwbON
QuK/3C4j65dYgJEIrBOLMPSWF0OGdUf/j0Xqf5mjYJ+LlU01WwN7q/EZMDiV2lQh+y0Daw1dORjB
+F0zHBreHiBkruSpboXeFNIpkBAK8SkUj8moeJ5GsiyGMpAz5ekOxbKXEMHHZYUWwsXJP/EWa/bY
ZgbPwbvtNn9TMAmTQUk+elCAhIluZf7bAhFpAoO9P/t+Cf06lZ91e2QbwddSe9yBK5/tycWvQIEE
xhX0BJnQUebdwJmr4FLHWwZVcLCDImmuyIsXyiRCB7D6TkPaJ9u8GE9QyXd5xIoaQ7snw10G0kjU
4rrxhUh4vca4BaTBp9QSoSjG7adjfTRM5otTxekX3rhQEZE+wyRFsQhfvtTKfpbulhm2RJDu22yd
aPGkSRLLtiucrHZq8ntRccQEnKWB7qrOiU9rnGS0hKO+lxMmbn6eMT3ipNoljXov05QPv5oG/YlC
Ap8UWvv0H3Ntnez9JblvjB9nedII2Akc6eN11NAbucpQ22lKPe82l7Qukm9tc9R8b95fM1QS9idE
CATSLQAU4VMXsejatn6KN53Z36p8tAg6HnwI/LjrKPk+owarlVLvUr1t+B+lFRRqvo8KbMnUJx8d
VArWdeLSwpXp7OBzt4IWkh3JmJbkifTuLHSNm7THGCVfinSwwfpYgOeTJKAQDQpe07aCJT7nsetn
10CLYnHBLNDLe5Jp31K0GgHGK2b14aks5iLkMg//jGtKlH9Et8LhIxsXVUkALtPjmbyTuRi0Qjz/
k/2K8mDK8178DhR35/Eq5POsn2rEhOST2BOqSwY0kT93uty7NZlEM0SYg0W1XqpNqM8BCczUD+uH
iO7GctLbWAewYHsASTYMHqmo2sEu36yL6C+ioOwbqeIl/hoPN+qnNQTX6D7oCO5dm5996+5pJI8H
B6NaJwwS6P7CHPJcw3xtBcNjcUWIoFBNdma8UpJz13dmbGdq4IDRjCZDQwQirpIZJieqOfKnTQV5
FdIR9iu5cg5LMdemKpxlfd6Y/Zmlc21xJ+kWVoZR2TiajtfAmpThMpMqMb8YK2JkK3fEM+NV+q/g
uqhroEorKIFOmnecx6IuwYgDpzHECQNxCsuxKOt96Y8L05kTodOmu8MVaZs0izb9uw48UoasxI1M
KT3I1dbrzD8xnmg0YaBhGdOvHWAZ8LrKeih77mCHBofKjctHzHXUUF0V27DhGlLj5kIE0JuRZlz+
b1vV5/mbhPzvtGk0nvDddpP2OB35LS+4A2Kfr7idEC/EwrF4XhPuWou+2xQu/VvL3uY10TFigSZR
uSAMxR/7ONnTCyYa1/RqtFDYeCdT9oZR1HDb18ZbAh57VMLlsFz+V0dJfTdUxveuV+ULUkBcTd4E
Bh39s1psqOMTvhxnVaEOgavgLyWzqPCCeuxngnptdGf6pqGOGPf1IosRT2kIZRdgh5bD7Ub6NKAY
qmkg7lKC8mAsMfCsZUsiIftf9K3n6WF+HKRj0igbIPDPi80587d+NzMDYnAx+DE/AkEnsOu9VUgp
lste5/X+E0NoPwNyObkB0MPNP29pbzQ8AVTJhYRhJvEYri3hOcYnbpObx0V3lNbNIJneA6K8AkRh
z117wN4Hi7oE1KChllzJssCKLj+z+nzORnjCjZF9jqu8+/KwJ/3OWm06Xzh6SGZI9GODTGLJhnRS
sxb0y7+ppos9cbtoI9UZeGGJ5ZqjmiDwLjGvjmUckaMXAUsTrhaDcWd7eN7uw/f7sueTwZUtkRhw
PGn0I38yalLG+IeKP7dX2JASph2SsJ5WrTLwIn5WLvMj9D7c/v8VT9SEMqhJyPGfdwZ7I2ihcJXu
Ylg7cYKHuDRXD1rXsZFcb3cYVVh3F8mIAFyFpULMpWMP7VXrnYFbUXGvtlLZ5vdjoxgywB+TFIK5
fdbLOPb9zzL5KPH86F1wrme8MnaagxZRe0NY/BPDMVegcyKkHIq3ax78GUP3i6TiuTr1ixZX8eSq
EdeRToQ66iVa6eSjRUo6vBGC0bf3nMvaMar7NtLkL4/wng3UfkSsedNmPDvVy8GY5WJyrQY5uE11
sAIh8J+5Ynno8ymsJLij8q3RAmfkd+bSJt7u0ELXOa9aFgSqRJh3mKQB7Bjmq+4WPgzlOcfUbJ23
uWp/4g+ly68Ol9ZKQJc5pAn1eQ0X83E2Ich/z0Hh8e8/DbG8BU7Dz7RG36WEMCdUL8t/QJz4CRVj
HRHqW/COBaqeo4NcoH9HX+uVB/N3elrEjf8ltwcUsFvofwY4EffpnfKiWQrTAMZfTh/uivWsNcRl
JJ2S+Vnq4MKXgv9K6CSSbno0KHnwju4Qx+taeImJYPA5m9V08aBg6TYaFpPOxkIsWzoWV13SCcff
ZEhRi8P/ZTFosOBghrYvQ5/u4r4M5ubs5kxw6k6+vyspkerIDiyo6pC4TQCZJFYhPRvpamivdvFI
RkMpblQz3XLn2WU6AzxkncsbpdwZ3pOqyoC+3C1Fkc72vH/xcGlOFzb0aKywmQA3f9tQVHz56gQ7
MttJgU3Sz57WYcBi+CZwjYuBS+F9CvmjEeH4S+QXoq/gX+L7VvkfG07khKBDHU90dMVtR9kplIZK
gNn1kU/ot4u/jqDZ5SL1cJ1JB95oKJilr0MJDzWBAkkZ9fKm5k9aIKxRvu5lqlT594NCLXsJpdZq
tai3PA1IvgBbMaYx8zjHCuesCjWs0ddSTPiWxFeICDrMDsjGCCaeH6mFpFLKYh48dSC4h0Vir4ya
yj2qXgWc4H5Oqp6+oG0hyakr+HIsDt57IzGru89W2TixDi0Vkx2lY8XG1E7TLpH5USuoXo9VFOfg
+oxU7X2jXwyZnC2n25wIovFNC0ISgwwdu1qRLwCkDA+ptxUlSMa860Mr0HKDQxr8Vji8ohTDfQhD
PaYFy8SeU6NqVi1xAaGjpUAJu0W6Y/+xqwvdVg4BmGsZJmkd5CQED4YY0Qbd4kauycnbLwCxzw7l
WfDaMcQyx3T5yKN7WVHyCInBof2iqN3/2l36T/LIEStAvoCzsh+5InN1ldEwAfKkmCRkyEolQVwP
vL+ou2f8eMaDIssF9NH1T4QzXPisaFNX15MBNVcI1NVEhuYo5ZJ0oACCSGnBgXqQc8eyBQBABvv9
5a1czjt8pcDF2PJ1Hy26srFcMMZSrUAAown0vCo7ofV9zBsEkb87YSHit4yzhESm4fsYsQyJC7qe
Qx5oaC2/gkBT9Hc2JbX9VXgXAcZ5HMHxPOhEt3Lm6XBgQFOC+uKW0dg0vm7PMdQKP07fSaJjXZ9G
0c2GAn6NM3ud384VPMgZVMW+WawtrxjiEPU4w7oorCUOJyWNjAF127EzsHBkcAvtTUZ02pQN6Gpf
/yiP8Q8uoytx1BrVb6s0h012KPJiGhEMgpI1XhHf0yfaaxTptaQIfVwAaLVggQbOs3P/ED8XrFdj
XjwLEb0BRj+VL7IMC0Zi6e4MDtiwjmcKv+NTKlQ43VdVUJcOtqv2UmorHU9xjU5BlX29JhjSoWbq
bCAdl4eegzqoNRTM8AQUgqefrw/qeF3ucZTvFtjv/Mv9axsac0grRQf00AIBAiNw/Zz+N4iC+KSz
Oe3raWte3YfBS54Vikyh0Nk/ZKQwVUfYLWcORdNNaPqdzZce69Rs7IMxH08NhyCL3cH7tngub+nJ
Xsok+OuNaYDlsHtCXVzjqHAHLKuDpMGlyuX6vtF4X5jHYThxgJbC9ElgZW8IYchSgVbosjvwMM5y
xtfRQxKel8aP3c3ZbQLSDaNxlxik5DNOPeCBY5u729YoR4F+SeVDCJTDn57n3N5sWDC3AxSpUeuc
MgKaetQa3nWMVt9CqvEUnaKDnlqi6kYtljz0QbVjvlh6lRpOpxZ5L89xlBFT6ybRKM0esj/i3jCs
0bRaHcAfPZaDAjKJ7LE68cuNzbp8H2eFFfyf0Ou9nlFrdDxGu35lWUulzhAiFMjV36+ztXMBvfd9
MUqB6b/nUD6xJuNUoxMhiSpXF1tXmH9aJSpqpP71TSgQKwDcgtdE7Ya/4DhucxZ8yKikWY37YG8n
gZ/OwiVJOmw0VzqiRmqnhre2D5JvAmuwyufDKq3d52v5GwQ4F3+KGqfdVAhpgEVwSwWe1VFmyjR3
ux/nzOz3iVgglwkvUXdj7iqNCG9ZuVejHLxc/+oFVdMz3gW9mHZR+RGKUFfBRhVhXeneVNetl0an
tI5UpcOH0yd0R5xDWByBizrxgfT87u/SPByWddTBG5kE+SpyNkR26XyQ+vtxcX+gsRTrza80el/3
QWfn8270tRGeo0KT9fuSWaAJ2nfMCsTcLNScH17l4Et7i0W648pDW15VIV4yeRhFBag0nLTfSt7P
SpYoWY/XoTYGq0cZLR4u1xLIrCYwtlZ5qlzh1wfG6E3cxmX4WRKICK3qp1P0+6UR6s2own5OiZh9
N8GbahzoO6t2ngMBC83jNSLCnV8I5ACimkh8yMt/w+JewcgyzlYuEVodFo4tw/ldFIiWAxtMrjT8
x4Av1RkrkzzUIrLlrDWkf1+4ZnTmw7W7h09fmGtyUtEpo5mikgLOe4iUKYnXSLNCbmj4vmwzjxdx
eBBh4tswAhaRAvZDnJrDrrBg8WJlLzwlGiHi1PKetHgs8YCcw+i/xsyDwtAvoC+bL1jIu0JeMkPP
hrq2km0PLoGHxbrq6cEvqIAJZZjLAgebcjeWFJjmleXoy7h/9jx5rJpcH4Ls5qzuauYclZIO96AM
I4sYORu/8rIcsR394SOWWnkAQ6sABLuBU7Zpk0Xf5vX4r4TvhPRUDoz991MJNGDWjInHGzU9kD6e
reUXk0u3Xks+p/nsxFdKyq9VUYQnQfH7OE5YS9YnxmFuEFYsrozH5A4DAXLSdRUdW7gE+b1m7y0g
37E3G1tS418vGJ+0SHS4xgkosUCKmNGcvou7tnPF22ucJF7cN/jPp5hxRdXCO3Vm/s+Rjh/L/m3e
Gn9nidHhFvNAdrJbIZV+86mz3SbXdpXwFh88io1RWFJP5S2g2j1PytF7Ack+MZzMkbCJlYdmEZRC
K//xh5HTicUYOTxaCEgRw/ncF+8rXrq6VQWht5iE96W9yzDOr74f72BUGr/gsIKrGYzmHUv9vFmA
ZdNnT6pWYjNarn7iYWLN54eKRm0sZqzSnJH2OJerrrVLsAo1+5vbFbfkIQV/uDXUY783Af2ExdBS
EjIZVpHRHRNqCSc/jyPk0RtOwq8q5NvJxhuQjSvZz5aINmYdU1s8vicrpH5eV/YmbdHv594yvBpH
Fq9PDsr1GWd4IE3gBz8p2NvvbHzlU9E0/hi7G0Av6BIGkEoY+svQYMx+le3br8RlE7b0Eln4emVd
ItB1RIXB1n8BTy0KjqVid3qQM5Ie6CEDDuk6x+3Ru/2oxf1CftPUL68v28HwS4jf5oQaEa/a9N0L
7sewGFNptXkN4ARvjiKroa+ZPbJLRhXbM5cddRehuzNkm1hl7LCJCRbR0bVQHSAa72mDWRsfZXs+
HTU0kg5u+jl87Y61IuhUFzz54wKEOJrQULNLiq/lhLtYpH9plk4NRNWN9uXUOxxvdJFwbYVDMgd9
vdjAKBTzEQk84+nkZTACxzs99ZZL92Exn66Tk0m+ySlnjqSzclCVmIXWJiFO+B1rMEHHn9yPdasJ
Xv6bIoOk5/VITnxsC0YX90I0iPBzgMP5Nevzz3NrgeC3/6pogE4jyPu1muQ725LRa0GKrj7qk93g
3b00LZgPQgt6tgj8jga2xUvrGFOEaJ7FINEj0NdEM5vPNl939xJrjqs99SVro9iBMoGEq7LOPbzu
0aXVKuqUnmQ4gK2KYe3eAx7+Zz3wRmpq8vz8j2adyu39ry1/aOOPtemgheIj+pbHidph5c6pkwMj
QEn4jzxjh95QPKdgKL5xtFCkpk3jWPZ0w1rZD06AJ7Wx1FDbr7Yey6cq9CjkIA6qdQJjQzlDbO8X
zf4TpEa3H9yHmaTdQ6//RZF1N7aAJp+ZtV27vl0YIrNtdClGayYwvWdfRpoNg5g2u21ikawg6oow
56TEon4lENJS4exLMpL+6wUPPndxftl4KPMiccM0oiSDOui5ocrdCKTC4FbvzWISf29cSVdgw6Qp
Q2UEGmaq7qel/KFqPbtUjWUTC6hvtvk2LTGziN/PjQYBnQ021bk3d/OzE7172PGumxpI4s4gYbu3
N91kV3CBwL5McOpDd92oI64ZsnKmtOf4BlegRHloclGdoGFDmbj0gBzf7hThkVgQKk0jvqSaC5M9
+QfPinIg3ksY8P1oeKf4MAiHt3wsUQOlaIPJhuN8d3QBEVTgHSigPL9nN6gcNKOzoWuoetvXv/hn
tMc9cwamSHQbY3iVFoTdsOUbcvfRy+HqCqWXwA9KETA2BG/bqfzjoxlD2D4aFzJgLBEti/n/YAOI
24Z49iMxSsACrit9pHoc5OxqQ+C16h+ZfByz3Qc1NZkwFGGEMSLSCAMudylwBoILzc6E4H5xnZCo
Lp24Pq7vV4dcPbMv+GMc0ySALicstHzRQ3EjYqtf+sQX/mpUySsgKPyKMg/5nIr9T8Ed3lFCj0S7
0cWUopeKl8U7ZzqhVaZo2WQE3gvc1/m2Z3jzThDqHLekT+6ZVfmXK3pZCrdYDTDADF42288yr4FQ
ioA67NKtUWsnc7wdhrfmAQjGcEpPScx738eatMH4hbEaB0+2Fz2TWP+zr0uChuO/cFeGTKyml9N0
rbtJH1vqbCzlvmSGRi169Bdg7V0q1oh+m6V4FD4EYfrbJ6U8Dcu5pAoRZ59il5rWiQsOYrgmqG/2
7MeYjTr9s8oP5pOph90Guup6g6g3yi7UEDTRgta6yvhDwz8nbshpaI52QdKq7ZMgpL69SCT+IePT
D7Js+CiEAedF5mkQyCa3PwdHDDpPEu+ePDtLHMqeTZj7sM758WYNbrdjq8r6YrA7xibwr7iItcZf
r7vFqHHBTB48csPGEqfsvmxWaX0KpnBBsDsVpRtm0j3QKKYO6tau4xjEQV3gwnkjiLWgW2hKExsi
TsonznHf05xyvWhEVvtKJAh7EnphZZkxA+tt+FprCNZkXIRsYLn37XTssyEedU2+vaq3FKgpHuXq
b5CSLdD0mZ5Ii9uL1mnOOAufRXfeQtvhfll41lR44otFG/B3R5gUsopbbnbfRlotkJC0nfctRlrw
87IuTyc/p/h+mip2NF/IfTA7cSNo6Q/IXgU6WEeidHcvyM51KWn5zwGxUrMG4zma/2378AiTf7x3
qxW9S3MUSPrVbVq7Av6G6AlGISZZ+W1kt0wcLi9zD/+9WBkOsgGOJBC7ouEVEJ7NRuvW3eg/jyT6
fUMjENMb5HhalY3KDjlAr3ZhC3Lb9MUr+mjmKfTsmvh0Ype3wx6hVX8df2QO/bkNlhNnLs3ekEqH
pWzo9x/eeKYSrEP7S3mJBvin8GSFABaFOtwTdyJWjOtCsN1SkZ2dsKVVrLr0yGZHAOXaCxeR4a7B
e7a52Agyyf2M5YEqT20MXM9TkYbaLtc9MWEyFbVj3wRvGCp61e3uq654iLXre20+xpCskDi6wXM5
cRWqjLjftksPOY878IRZe5Mvu1yuO0ek9SL1y8IC5GPdxqy7blgln3vGH8rFUUJiCN8GQuwNAmee
KDx4aOKu7uqkBYDy+gtnYxYFOhxKS51CHJKnm8rHwY0Rkehn9Roi7+X3XGU+MC5AtpcmneG8yXtq
PwmizwQLgCOJn7q1qKJLvbDBhJXMB+S8udubyO0NwDY69a31w9u/0BBI8XVLGBfYHfvUrD5P7wQC
cXJGFcVXtAnfGAWpPRZOY7OZ8Knj0OVAwR2cUobLMAJpYs1AapG4w+r4tDPQ5ukd3ghpcm/DiyIq
//e7NdopL4uLfCndb/LNNPZ+9oP7ZW0v2c0z4xutVLQz+5MlPxmfrAX1nN9/MfxjwMy6ClV6th9u
BGXabNB2fWqDus6BQqSLLs/GBzF58+Ldy0vS4WCZcHzTL/VEX5L3FX56hTlLCaXiZTS4mwBjFk5A
7CrkDvIUC5Nlvms8ox2Omu6bnwQoRvdtGhY0MqTituu5KsQZx6HH6R5QbD94X0Xdhrjer7UntngY
mO9PSLgFW8iMCCdg9XpC6uHSbbK6lyTyx6t6H9/+UTaAMsZ2gt0Q7FsSWB4stTLz34D9OSKTxZJF
I562SzO5To0yEEr2iIVgy3TjrOsGXeh1lwc/F6TIhf0iharro30w70A0WZgoYrvkr2piNb4omNjH
YloYHhk1KyWQnjpXfCQK3HPIRebxujpBVi2cgBS+925tt2u5CHy6auAcwXKFuejcuuB0J1M0Z1/g
/C32sjItUK1uj8td54qDg1gR/Vi9IOWxXPjeEMZ2UtlQ8lOQJFFQGA4LSxtuATQSx90DHJG+Rqoj
sgfW13RiTk8V+4AonRoW11UnKhejx44j2N5HnwOAMgncAygtjb5T7S//iklz7tgmLQS4F745EoKM
uFS6l36yfTj0avSmeMI8XGndLn8VdNCNmD9mKHOGHb4Ctfnj/14Ru7MDD1qYu0zoZstd8Rs/m8KF
0GbaIn/Qss8phiEbkMlvfDhPOtgsF0qYC2TWC0s5d+LmsjEzLjPwmW2Dqngebv09Gp3vMfJSfKMg
u/25P9t+elpghGtV8p5JvGbOyPHAvI4ZX83QnYbLPnf2YzGrbs2b+GU7E31CMwOW1eHLVKPUsWkk
ULXeWMP6qu7P2VbwZ4JGJwiRpV0MYGppqfNtFtHjMbRiUh/9FQArMQXtWvT9xsjuL1MYXDjVWT7r
cmqyupJ1jRZfNLLALmUZp19tuKHnWed706d3yexv7P4pT9lSriK83gjUP2FcmYH18ld1jzNHGcdI
OZlM/2U3FparcMighqobV/Q/Y2bxl64d7TBjnBH4hvvOfvaMtSLgkyxfHbQvdK9Zj5nIPBMrwPOg
lL90XR7LfDnKpxIcBAQGdzPT0x0oXicdid0py1bTr5/6FDsRnHM2pdpRpXtsZiQ6HxplT/BupMKp
BQ2oTwXaSBoEdqT4w7jGMcWbD6J/Qhnlcel0gQ7UJF9rP05b3rag4F0UIvPwliKSNS475fxJ5+WZ
bbpqjAzLIUa6LvRASMkUxpmxbJwQX18cIWvrncANyglDSKgt4qUVw5RqRcN/MI/3cvzyg1jktJSP
Wp6cmkZkekHZwVxtBjnKVWj9ER4jaT7s7uG28/kRUxkPXrNzlLChAD90ZImjyHCafW1ih87gG45A
na8ofqg9+YBFzHBCmQQUsRopIR6sjzFdFItpNoAnGrgEo7X2upgBa+R0WTN5op5mx2qSBOJ4ArGU
On+Ckc278xmYsc9B5VliU2X6/DT2jr6mVNj2vF9OgwMqjJH1ObQxzTddchtr/2OJjeZpm+Fa0Snf
9iKJC3ov4mgvAD6+wnI9+PnH+0BI8Mgpu6E6K15d1u6hOIkemepf79oUxVxdmcY/Ok8vopgoz0bl
rdEux1+z3C49Hn5lf0zNGCyuaehYz+M9BuUkT7AEof9ERCiyty+PexY9zlyZ6qg/geGE95R1+H7t
spLZrtzd9gseQ/igWYSy4+dRX523GZNiOrBi6UB2wgqS5T1wp+0j/5mxzzwQ//PzUYQW+uCgsggw
5H7rE73prAKx2LVae+l4KwBQ7JzGW/EWzZv+HDWom67kp35W/5xAlhqXixlEu1wJvP8OECBrGBam
BFi9CHzYVHXtt7RdRMy64L1E+VsBM1h3Llc3ueQXsFBVQkHrq+7BTf6Al8tsVTmn3TYIYIwYYaT2
sEpg5g/zeUL+Y2GfY9vsFk42qTcgedCIDXzyJ0RotGjoi1qEuOJE/z5wxsWtsPN1Nlxe4lPz4dAI
K1QBknQEaJxsethmZgwLqkoSTbGS41K4Ai3vJhDHR2fZbAafgpOUSzJAJaVfNLKADraxcM4JuIUL
2LlPbAsL5tg0uRJwrgk3F8LK7DTFq1Sje7UEh2U=
`pragma protect end_protected
