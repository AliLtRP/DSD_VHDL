// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:39:13 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
SQ6WsgiLBiVUG7QqBI4fMERXX+FgHPvt23pn30zkMaSXpc1BcR9lkRE7Q0jDqpt9
dEQO+ZRG2DXMOfGi2ZtUkLy7CDITEzOaC9f/njpMeYebXYOXemSZYArWyD1Vaie0
RqUupTOazor+Tcthc7b7tS65zTmiaxQ1ZSoKnXtl+O0=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 25664)
7G9X9VDmGzDYYCwPU6rGDhI/fHvv/Vtfbbo65y8FDFaDCA6cnWj/G3XmNtqxE9+a
OLXBt00Ziz2SMSO1cUtaiZrps/PDSXZpOGs5pgNqz37OfE3l8OJlf13qZUikMlDK
8osxF5P/aFM15Errj3mOrs5QfJZF8XfdJmCDogu5uBiqOP+PtMdG8PKOsM6a6+mT
wmOr3d/S3R5i+rystJgzDQeDCF07qHo5Xb9qeOeMEbubNz/BymNxHqJtYhoVpZj0
VqKIwHxEwkXkFsqA+DzZkctSEKf+cIcBLeb7mHZ+cjQY1R9nJzPYZz9hsmB8EII+
87otQiRlarvmwg4ecgbp21DZ/HZhT7p+45bndI7A/Lryg8I4qqUnQ329T+i1Jsfy
0xgUjrqraQacXs91Rq5Y+0ysrs1F2O5vFosSCTIcM3yEDqap1bGez4yD7X50DNEf
8TjHvrUA1pZ/XhDFuKY/zigd/0KJAn1Lm4emH0pOY2BiEw6VakAtew5Kcoff9Tch
9UpvbgOJbnF9axuL4I3ZCI0cJoAQRXqUUHc32WCLf220szX4JW7ne+wGW4SKrQqE
DPPkwfMBWK6kiYWSS65tZaE0IUNVdHlqovS35ws9DFUUhRcFXTr9qfp58bgHi7Z9
9c8z/PP4qxvqPoLeJ9/z1U1uv5dR6SK4E1BpKIJgCTXmuXIT4ORhkI6695tWlaDK
CXD8hMhzItqjtPq5wccCz1q6988928eN0fC8ql2JbF1ij0q2I/hxydaG6ZrQsAmP
DYzrKFC15x892jGDqAOvvNjRpyrQcpcb30EZcOYD4Fnc6xtNTFftURGafF2Jkxvr
wY6bMKWljs8ZXU/O77Czw9Z9Z147oLCLZ20vZEYWg5ur019ds+e2fD7nj0mav/vW
DXsKj9t9/L2BjIBtqnLrIfwum1ja9nUJNnRYrHV3Y3ZfhYuyE3R3RoLg9isfHnKO
vGjo9It5N025v+NtrvlL60gS5Rr8K744zTUww/hwW/t2jQIbH+QwlahhLRrpRFw4
wQzBOan36DUREdU2SjfAlgVWFYf4/dcuAewNEOPPoh+RGlOCgyS8dhAKPIEeZDm0
oKK9MxfvO497LQ36Je19vTlIza4dECIk8Pi+LJz9njoRnLJf+S6Kdlff9s1kUM7W
dKBWH/y4vw7PQv4mc0varHEv3OnbBSChr0FIrn5Mke+G0tMVO+rnVjsZujMEG27i
pP/dZqwnoEGGgs1ZCwUx0FyG54CdtQBhJejrzRpYhXTsbxox+79xHJINnLRCx5sR
9Jpq4ftvwfJUPP5boX4ZuE68gnkFTpFO6WEK2buOa2DPMzuftLwZ5ogmE3pEa82c
iOT3HRcfPlVP+PsDake93KhtjnbiEtd3enmPudniNGAurBvCuSI/caiztgbTmBvr
UQT8oAxnt0UfaRPYr+eH/UpyyM9Isb+GOXkY9Ru2QxdGtnLoqo9FyXPUWkRczP45
GOy1vONkn1UUfXQCQJW/h8/GNl0T3kboa4UMpz+6i4iemyPo8Mb/tEz+eJGGp455
7vBAqi1JKxMvzzGNaqBRoBz3Stgd6iaAz4HaptJeo2taGCeka00X78BkyNL3LXcv
VD0xTkE9dTmO9ZDRRrbcXLzMSjVLgxXbhYrY3gotTAat+lvqDKs0aIxlkcTHwHIk
KNjI8lzB5maP3Npv6a0P61OAG97xtCom6Rm6vyM7i0lMNf7UfsIT4iluY8EUMp4p
75SKQuTzgq64jDWf//jlqugjnN1B7FGzvo0/vXhhqu8IJjVXPnMSLfZ0bysue+5X
fqsbAPU19xRbHbOEoS3RpkGZb2mFr4YUHDIlt6vb1+RVrKqdUhpvI/OD1EHnnoB2
nzyWMvCAlSDYSNmvgrAyZ5TFa7DP+Jnqo62I1BgtvFAmDxDGiEO7YHunRhsCqZby
GouNDFamD2XCAEpZbqhph4MkbzX1oCBjVkOgE6bsxEX+9LLUbeZcq1Lvj2H4jMaN
20MEdHnxDRkulr6m1HCkHNMXTsbh9GVDFzjEhmp/QtiZNnG2PNejFGy+OgvupFPx
+Hy/1ABY2nW2jsOESVjJhAOmeXjemIovwZUEtzAEsoeJVIAUnKyKUQQoGflVPBiT
Gtinp9NjwJPo3kkO62+exmzpS6BSYCj77oQws8nTk9MeusPdXyCiFHmYYAL19QgW
ekt3pVecbmFzTeMU9Ait8Pv55FG1mpK/StMAapft1AFfy1Qc0ik4X+3hGBnbMwij
TdUTPSsGT3NZdGTQxQtfviwzjQiS9aEstlWy7vLH64MYUcUXdQshT4FPKrxCBTjc
ykfPvUiTgxOqXb79tfccmHXaNkDQoHhFlRA33CSBsS8WE850M9eyQvt6+C5onudr
TIxrC4Q6WBk86VymDvil7Ct09nN488l6JnM5ZCX3uLYvO1K9OzefQ/phyeT0UxUV
JkuAULyEGgEvNLgz87o538TfWaxey9NuD6Ux5xtsZqTfhgdDnMyflfgnhOG3bKmf
WaIY9DJwe0W0SzXwrx4EbHbkirItWBoPIFZm6Knz4MfwQqSg9RlzERo98mXmATOG
06VRlDGBWvfD27qnMqLdC7XOtVkb4QcWHGtfuaCKPpmeGeQ5NWC51JA3c0m89Ygc
DKsJYkzngt5F97ewWCmvQWBMuwte3rxmfoJCHg5iAU02yK5QMmcAgALtkmZJaibq
gLBbk/209xGl770Z3YagMdZKrqJPrkJh1KyFKR51u66AkgY/WgrPzAIgw9C+Vdpu
IEcXR5gmqxG+ZOujHdfD+BY4zTkTnadIUXPuOP7wuaxRnjlJZZJDKrYFD1nF0ntK
ZA+Mgf0Z+I1trsgNXRWjERRPfUATRFsYA0p8HnXmyQqZb8DbhRYy255olN3qVvJx
r7J1MZYdh8NMu2LSO3czut9QKcTMcEHkDpqLqIiLRGLkW0ZSqsbPO7C4scVQzk6Z
RtnRJXmbwh3ixvEbWgck+Njvr95G32jT/zsoz0V2XW1ZNIo6Cap+806a6CZCQhWa
3X5txQ/0cD9n+Iet9jYdABSIIEaZCBZAgLUNUKZgxx78GVVoj+JK31yI67l/Rv8F
1GUVimPvVaEYxaVBdatv5h7CNKw43DiZcG9xDCAF3AZmx8wpNq3JUvrC/042gkfs
qWi7HmgLn+jc54LwjN0teHrcFBjX6aVIJGKfROWPfVrRrz+ZyuggCK9qFODyCYP3
WCzAAIETcp84Ce47VDsgs+uQEEoKSSeTwLnMLZWw1ImZpimJTX0qme+fu3M/zvdg
eDPGDSiMo6zUEW2CV4yA74mlzXYKudRJvjDwJfVIBvO8qah2+eZEEA+BGWaOMljm
677klaX6KCiTimbmAeFPKbkNwNW1IgyQiVSdOZzZSm5GSL3KqGjB5IDahZv8Lj7M
UcXopj5dj1lGRY385vE+ckziYvdRK/C05R31H26Vgv3UVDnGZIEagUssIRPF3XL3
kBWUP25x+5FvqYih/XSsrd9c9qVQq3y6no6C55Nq8foxOb56BzcMpff/qkt9vAwL
ehvoyR7mMyEPk6FWl4lhh0MrwB/blWLdLFyowiy0Oj1rAnn7NtquSC9wv3lubsq0
eRTP8arFJ+XWRP8ONCJHxhzvEJ3Cwcq0FHnUGNW6S7EvZljIil1qcTw29Gc32pgF
vtUYOs4UZweB7gcGdVZzzEJRluU88MWXnUOkX8zawenTucDen5RBKEEVjoUEh3GK
5Dz6t3yj+mzB43sL7idQpXoQyCdLlAtDgQx/5XOUJY+nhui2uJT0uChut2lzvl1N
/a1JRZLBtROMnHsicJWhL6vbwbyRlUQ6iv6F58kaMdXAs5jhqq3UlmsE3nu4QiaG
r9oAOV3Z4CkhMcRCZhWGeQIvPNsTTdKERDy+iqXMLTYaRbnjiRQuSRTAkMdhWpRq
WtW0cQHmVUXH5pYBl+3S48ymKvy4Q88u0/OdDJjdLI6YU57kfKXgPrH0Q9lxoxZW
rLHLdguupIMce82lxsFvjQoJFPYcJC4WyeZSD6dRYVTo1P8rDF6ZJ6DLMZm+wSpD
/LL4gLyMOI4x9Re67WGLvodWklZpMbJEV5b6MiknrSgbszcwxCewWlZykDpCKMDR
Z8xv5b16tCh0gWfoEh8wycXnXRBAWULEUOVPu/m7IuPYn8JN7esB/2rKoxHhdK4r
FmtQWsyTDEHkj7qorq7Ds8Q1YC6z1ppmBWgF4A+1E6THqk3UJDFk7F+Y84mjRdBL
vwm01cP8ce53de2pIs7RKuLMBXfbQgJvid9pCsH+bXknq/ac9is+tCTOUwEC4Lrb
ODxgytmoIUDKHaxaj2zmbIEHMnrQduhATqof76SwTCXZPvQzrIZZV3VJ9FW69eh6
FSUW0aPy/XCrTSuJjQICkRAxkk/Pjjvm6x69bQHZgdofz4uxqyudcaYHMeZYjb/d
VwtdonuH286HMYfd8HGllOvOKe1tZ9Ke4cTTZEjAnpl0jrdmZ5jFdyCAUiKdrz9N
fyQHePhjV25ePhU9KqYorlYU2lPiy5eg3+CNiTN9lQ81jU6E6pADQNg5/09V4g8e
ptvLiVjLNtLFL0v1Fvgl4k0DciAQgsSz+7H/4XLQAVjW1kRXTnBVybn7dj1mWFOz
n8i+bBxrElkdhogVLomVFPaTOLhzDvLuPt7A0nadhFnAstSyjeE6TgvSCj6/kq2s
exo+NM7wfob4JQoLbEUzHwiA53NATUgcWhsYrNXCCn61TBqn7BJHtKo+XjTxsohU
e3KCaNeKPLO9ZlVRRNF831W6fRNFt/otP+M0JaWgpwnKzKaJmtVAw4l5zubNKQcB
bjnt9gtXxyktzAV0JA3FkEJcVa+nd5MXTDlvze17y/b+/LLMSb17D3CXp3CcRi5+
0KZrL1t9h3Fecpxp+nj23joJa8NmShD7LSo9BhAvt5iWz8ZMCEt6A9yztgjc5h4n
p5TauH+6fAR4abXx3hhneLo69a6iipukPDZdA6FFd+IM8K3EbeGvVPrRRsB+oN5I
taz0om6VaGR9FYflgzOp3tMHvLK7FwqmTfwOg/WPhFmV4WxD7DthJR8Ywj4ywyBq
dy/ugp9mJ8v7LT2CPBsHpE6L7hhPwqnNrDPdJGxFrLEEMEAsfvmjbHjQq6whOVa5
xOul0/dGjnQL5A9NAeZWA8JaP1jinLW973N2oqWJR5x7M52wFbu7xMwIOO///VaZ
IG4GUr4FGnQDJJDDogHl/VLPXOPxNoXNu5YiFZFbTzVbKX5u2PtM8Z9bak9ck9RX
SkMUxsVeI3jqPipIXpJmPMR6Idmv2UZexwMtb4PhTiqe0lKkhBQ4N6Ql+9K/Poe+
p72WaJ07t8gX+4W/tyqDuPcwqdP3TPfKsu48U+ZB1qGyHbaLgbN36iSzJC0b2wmd
L9gDdldlPjRJEhj6AqCE6AUi6E50cq8XLRkJCb1U4V4A0cznhFelCjV9uSisK7r7
A7eDXzA44sh9VMEIJA4/p+bJP/tzftr76r+A4G9AuWvnM8ePTgUHzHcaMkTJfgE3
OF7RBj5PBdqvMPrk/1Uef9O5flP5KVXwBtJXtedmWY2EoM4VPxG60yMNSS8shB3W
8JFwiYQn2jd89QRY4woGzuCu5heO3sgq7G4eAiVehCQSkW3V96rTQ8Q/Kc+4EvHU
6BfDrnZc3PLglsgqFAWNTZjblcpokTUs4Hpjtifdxs6oJQ+voPJJDjN1tz4lGdbK
6JtxDAsMXsMAPZUaQMr4D9SADt1bYL/ADBVsydiI0Lv0grIYxR1G1aUtLcnf2GLZ
Ldfwnd9WjHSIrwKinOx0+ICMNvkymOBXnv73qxhmJ2w+v9RDSn7kn64CmAvvNl/u
BdpXIKvdywWkZHZ61TrWv+U//xWNau4wGYIBlwREh2ql7pyMjSqOJ4Hzk12a49Wv
HYSeMq8Ki4bzmO2BKgs35iVlLT5cwEkdTObuUkWVMzHDx26z8wpCN43G+RJt45CI
MsQR4+F6pJwYVlG6EmMIBJN9FqN8CaEkTZEiqYX3Xm7XW/AKo8EKJQGAn4qfrlux
lAvWFf0ueB5DFa7q8rMS5QMr/oLKcR1JT4GAKX+SxwCQI0JrOpenUWSt9Szkpv9U
fxQaJXvVeXWlreK5jnhFyhU0sfT11v9nOOtkM0CQcDV6BSIjEzSeZaLSLDmbk8mu
QiG6q2DSxIEh/Do6+R1AzxYwmZhYxpbuzB16F09qvRKvg16MkZgh52P8BCLmllQf
ulTFUNLXYJJXDI1lDRgC8odrt1URTvaFAnfsC8SpVB6eImNrVjNJp0kt1HGfyBNH
/A47rHCbsoxZ8//Y1A36OhqKoFAWN0ybLq3PqR79G2x+MmNY+st8EpibcHSnXZ6S
6nPExBfWjVYM+GDf7tTXruarpGTn8OK4WhUPJorIDoIk+8ygE+wU3CMh+uaGTVuL
CzI1n+0M3hZl/yY56EgSvdICWdNIFNEXlKKxAGRyhMA7atNIC8R8P/nN52k9304v
1aUKuPz6/gbzw8utkrCpnBbxDBLUjgirqk4UmAQ7Z0YKT1NufZQnpXpVdz55rdcv
fFwD3Fwd/zZkYdykDn8qSPD9xJtKBWWkw+XLIoaSJuRNEuaqPPJrAHtSFdqZBvyO
zLCVu5p0Nih/iy8wTLd9GklBwvteX7vHepUrbnKHCRO4q0mIJQkLN4QkW1+sOsdo
9NPdgHQfa0M5Xng9HyPi3nMrmtaAqqA4QnoEkv0GFGvfAE7UI3O1gfa7hmlr2Skt
FU6x9VMFhIhTymnuQM/Bv9dSe7xSRfx55OS6gNpaMuJzdn0O8qMz/01hjPZVush1
SYpmSwXIQbHi27OK/V0QMmt+uwQzOV4rFm1aQPckkV2+wsk+YcNZyFXlU6qpd5Lp
VjT/C0BZZleoFk+PPiHaosyKpJg6oSfkp3Pfec0oYAkAm2OBoCEnFIZgu9Bi82SE
MOfoSXwToKvpmmEdmDPBi33/BG9QoHQJgSQmQtvfsqYMEm9hwlMSrO4OtJCotspJ
Nb9p7NZLtndT4DmrVTjFhbpMwjPISVmStYV+DB37pbqjYRFc3CjIwZsbOM+8auzY
aOfAMCdLOpbr0yK0RTOijvpHBX3CDFfBq4/kZB/aD7yQrx6wu0j/o+5os1EZPd7a
k/SCbFn+4Wb39AqxmtdyTZXKbifmqVHhfbTvAkM6UxOac5IEkXO9vDIpu7vqRyF4
dg9JkqRMNj7E3KrdrlsFqbkgfCxifgmeWTfF/v4NMK0zxKvdF8/0Uw2UUpXoBrlN
tB7wobRUi/aC0srzNoMQFy8QvWtvFSjXOo3Rt1OQlUrUIfukvGf/1M88IwnfBsiY
bWGGpD8CNFlRlz6pSvaCTZnFd0tUstGjm9xDwbhhC73rqVsa8+PKYwu013eRhlPF
PZfocSVaREoULx+ypNVH9GF7BSNRS50TOW7Egr5uAUdB4/60lUypHt31dArqEoIB
hmR351pgT70d2dll2FHnSlde8ueRQpNseNSgrIZlEBxhCp60EgisGCe7Q62IKHwr
RjaHvw8HjtpCA/mgDzGYu666Ba1h/U0i9IokKzisstnrdGYPDJJ02QYTd5KeOR6q
5F6vvuvDYPEdRuzUvWOHh2xaxTsmKS1eGgkQU0OlVqGtuyfcqf5+AJLdKMPWPFqo
F0CtwoAVpF6HwENnrvIhfuRI1mbuh5MWnKsAb7y+ieqp3RFf5Y1edqJG6zDSpSIS
j5LE+f2fZOJjxzB0nVLiFc0DA1PeL95HDQu/dVF5AMcqBtb8u4ThJgtOiTK1S4Ap
jf4hl1rbiPpRhCMVZci9HIjEtlmQnR23Uey/wc4g/yhZ2/143GedPENQYz780lpK
hK+wAdn3JKEjAQho2Ki/4ms4aY2o4s0GwJETFAW3e+QR/iW/4zNMBjXoFKm7DDYV
7Fan9NNg7+kdNszrbcK15joHVZx+vTHBM8V+Cm0+sCI7H8uWNrPtK6Ny6gT7t26k
CjYgCPCay/HnVdsGsTqepmU2Q+igWhSoGCyR2+JSsA5DrrXa9Abiw30meDY4efwX
D0x9rfmbP2ihUTdTCt+OJk1m13gr8NnBvbhDnUCNBgsQPH406853l9tIsuVnjNv9
xnz33rOI8VrZshnCu9XLOTFmZmZaZz4x0BpLoiVbRaMXmZ0j1Dv5u2DPVZ6RCaJr
ahfC7T+P0hayTDAkezq/hwtMqvnmR9GDp1ItaEP4LWpigX6LyNDiKQrT2kfG9lKL
fuJXANJs5hbwNuofuyF4tBRpHlUZCm7R/X4SA3nEv58Zb5xy+VBeJWd7fqLVkShi
n/LPYEWkFI8gkTmSRyACu7zr+oTuWfogGz0VGiW15ZeoXrkStQCY5idAD0UdLV4C
c6AjgowghfJlVCgDXfpcJBEhVojHgRMi4xnBkGJPXB3/mtCa1RX42kvsq7FgBPhM
+eB4Qww4MBz5f8MglAjRtlS5E2N4FRsjERtHRbCCAcgTN5+8QTS0AjtocKBsztq1
+V8O2NlEndHKJeox6bF7znRpzZA+hHq1XAxwBR1T/dG3D1udmwUcjBV6+37qA4CI
hHRDYCZp+EkwZVmrk4xfdgX5DgQX70KTwkdl63XdJCc5CVrjApWJdrLGmvzAXY6E
vjhpTWoQ6ik4RqZ2BPu+4mRyCf1LSnvYNhHcku5aNmzoc9bQEeEh6+7sJ7D/f7GS
VyQI36+RtJdRAwnouDiPPHGEWt5YLECncAb8gxaRJUHjcc4asxV+kzYH9IoGxmsk
7mCTVKIGe5mGWFFvUkKKdZV0k+OlvkTmgRtw6s94ALYdC9KjLeO4GgfOG3QgSJvF
/ak2lTErbOAmvf+mdd6fbF70MweadijaJyotnXDhiKOjl4k/nQ5BXD9AqkMLUAeX
hfxbnWM5iyYWwh1ksQXVY+ukpbMVEse4IhwWP9iIr1yhYvK8Ixqx/nAylc1FoJ3P
9VErB9JP0qUAjVU7B5oagsO/9v50fpec2AzOq7yZNfZBaF9P28P4bfFv30+hZKKM
OmmRhoIQ0qyk9DMUVJQzZPtM+1Ee1E0UdWKwB4cfFVU1jOWrxqKJWowpwO396JAt
zGbtcFWSG+CzInfhAlDU9OriXDyAbjsqTCi0FkTU+78WLnX1j+pqF5Th0za/6FEq
ClAA65jefwBeVH3/2hXUxp7axIrQHusykGpJfDyXHKFaRPuexJ3acQ2nQTR1XVpo
PPzISsjZMzlla3fqveHh4tSZS3i2rpm+KEN37NxyHZUUdWwJUnolvDf5QM28O0MR
j5CdKshi7oEaaHUo63eLL94JNvoF7mk60GZdtGc+LeZq+5Km4Ao7thMT28mM9Bqi
A8HifOC6OZ5IwHkw/WkYevXlsrEjbvz4QkkgH2qWDNHNjjFYEuqrjw7LKRGrbgI3
Yd5ZZUY9hUDEedmEyo226pyZ4C9RPF26LHXQFTi0vtowNlfkgbV5gotaH9N/LFH5
BUa1p5juhBRh75aItep5JEmo7psvzVj5ImxDm9o1IGJTQGh8RcW7eBNz3MZIWN/b
oKp4y+37/C252gQ6FvYiJgeJEfC5FNMZE+tlhd9Je9Gh7BsQ0+NvJ58izIwGON9I
9tZ1QnAHEhyyd1WMO4Ml6oPci2t2Jv35X01KlLEXj1uMo42dqWZweDME/s9vxLy7
lZpcVVNiVyWayyH7/oual5TRqY8XxGGIJ97VhJpdlqyaLVoIOI42Q9B6DStHpQHJ
YPH3l51J3HEvjCHf2Trmey4+2barf5BJMiCP2ub2gvCG3knlVxhMicat11l8Gngb
djxTunQpn+HWdfEUW0BJo5tw2RCeq/QmSDiyymA48gr8gbuEcdqlqvyYzs+arZAS
PDCdQBPs87gkNj9nXvOpcU1wEpjz6+LpND4HhPXYyhQ7o5xIImByEBJIBhy/2XdM
U3Ak7JQc8wCi0FBxpD+SrzUUV+l+LnyZCFTl3KeEw5LfeSoEDSeMhKZpyk3W2iPG
54oAZNMa2I5UFAemdoH7BTcZAAGE91Nx0Apn2xEIxeFcG6N4xhdgpF4HAe62KpL8
0wgljCJRzfteq4ASNwJt6loia9R3Lxx0SPdCFVtfVDw/Swikgiwc4PlBCkzCQEVX
Hu3eajttmENVXNnGrrW2O6eDWTrqGAclbAdxe/TayklUUkuop7tah2nmlV8BMu6J
wLzFviYVTcJYb596zNK4XPi4XqzY3ntLAQzXvXLqWlo4VNo2ooE5sq+0M6j6godC
0WiEZeKDx69UEzDFWXn0B/ppoIKj/YkWjgV14mUImy0mHQkCi2GdKxSNfWW4tWt5
MIsvaJ7rqeY91SlfpplcUw+rIdSmcqNXFglZcyCgbX+qRHZ27EHezk3n6txNjj+g
jHQhMdWG0CWzq1uTE3IQTHTyp+ucZteVxPgmLzFhMab9Vza/EfLxR6oUOPPm/1nH
7VbvpGnk9DFHBz0f/Ponwdejb5N899DuwPnOvlUtXnRqHg4y2GwkgG0w8iZR7CvX
ORLAQoje7ZnZl/9BGUiRRu+4oMtHUpAxTSeiQySNWaPp09YDLkkeUcoH9R9I4Zvn
NZ+q1/sajI/5JMXKPe9FHw6Q7L3lay9AgW1QPPbRCKlK+x7uuWfrcb+L7JUsIaYp
EATDKufjqlOLmlTO0teQ3eRkmV6bT51ZTHat3xxH+yxLkf0OUDEQD5e9noM8whS/
VTmnF3wF+4esa6Zx4xiAfyMt9rbmX/97ppvPT/NgZToNn+OZwyLfFuAucVI36d2c
a3e3OcMpzhfqYzNkKTJQKXILC2pTs5DSO6yEsjdqG6w3SPWV7SPen/sKS+f3uUIn
WTSkDChc4s5p8GHeHZKUFZdjuuIKdPgefrndD3k09Zo7xUu7HDffdPYptse6k05t
95E3Kh1Bt01OAm/rD/a0SjwhU11VAoZlaK0LtfE46VC2X0JvczqxnoIxlvbxSF1O
+RlTPm0ys/urjtP7VuC7mhR1T3esrTrVchICkO9wJgO+Ocdv7SRCjFSYKy/rdwpG
Ya+6y3bLAE406PrNxuSSofKizjk5oxrPyjmWUh2la3xyS7/s4myw+a7dDNC+Xwc9
wT6MCI57iQA/7G52SP3U9/NHp8AM7vujsi8xfyKmGVS9JA6w/IWXSiAXJumU1dDs
1RNWX/0GmmdrccGAdN+rDO7I8tJNUeSIXCshk3lXT7x6pnoBMA3JDfFOEp4OPi8/
evNJ/L3HiiTbFXOhF4nUzqi7GzZDXGZ5DPXeGZQUKJpDzE+sTlOSdyMqJTylXnLC
edBgPOKy3+oBFtTROLTrG+qVLbWTF9zxWha075ABLEakpFKytVVMqCXnddVwG65Y
gECFWWtmRLiy+lwXTWEk7KRqV+iY+BZGOHXds4DzccyUqnkivt449+UcuFCTvKfB
pGu6j/Op2VALLaCMEzqXLcOEB9z2ewJyDl+ORqmhCUx2ttjIEpJBepRe6jQxpjCs
z/wJdh8sVuIYhT7KdfUIHL5UWMJ6I9sC3OrjmFnKFvMivO6uojI1NT/uVRRQN2+T
Be0313L4HLU84all08GwdQH1tO1Npp1M3pgE3zEpdn7b3Kjd55ApAqNs9RbKd8sZ
608vRwaYT/zCpOPv4wk7ljc6aK8/KceWcovxKn7T28oqt985lyrZj+M/v386eo6V
uScOrqAxQo+inXTzGMvwkaxwneoaHtXt6LHUhroqBiJEvMmz294AVFjrkwolve2F
LZkz3xzz8J60JfGa+3EOOzRqm8hnY+JzyE+MF99bKbvLgorrjDWiRwRB/jCoe42y
LExIJXl9wPMAQSQFTJvFkTa1Gn+vq3dnPz5T03w7K3RzT7BFoJ8i8HuCByA5Q1Vc
sHZU4vmrCz71ydvBsBC+s5RvnoFBwGoWtM2vXY5P+Inhljlh8qjrWVQNauOs0w3N
GJZJru+sq52luJ9c13hVDFSwZ2J4ziVCEoyZATlEoTIY+sBSoDRLoAvREhti6veM
8LU13qOn8Q1G22q0EkxBV4zJGUD6x6/mkpJ+2zTRK7mu1OiANnOyjyq6e3mVezSv
60gDx6bG82ZOfo61u0ion4TX5B2Sw07e77aD/+Mr/wiWo8219qD0M/nWYWnYUHP6
VqcHWYmaZZmjrysA1TbkN9X/n1Q5rRLyU+KYPUyi9dFRnmP5TCpCJXBSq8WR8KKl
ifN7qyHZtpN3ryI7n/BjtzahgS7Hm4HhmmncQoVM0/6OV52aD7OKrAq4LvsHxo2E
U4H0eQVldLc7Owyj0XA2m2PkQ2AX4xTBaDRVaQRuR6SK/qPh/DnjJ0A4QN6P6rUS
bYAvyauFSC37PG52q3GH5RY94SbWKHAExSqmM+sf1nH46FLyT4NDwMicuEJ6bGXJ
DtXekr8o6YhpXgrTSvb96qkPajcMiAaj43hrk79i0xBMINwx0GbH931atTJSvpRU
kgCAEkMHDIthRGA4ZmNKePhDjXCNAd/ExrLa1DKv+O2Q8yDvDJNMr/OEwE71yf28
FPOKq5v8LqqaFi47n+9PsbEgU64HSR8W2SMEVBaQRO3PEsDP0aUx5o+iM97TnIDz
Nyx6yphl/vCqG9L7iHqLuiosXAc3PupFBWchWKbkEK2QE3nzo7E19qccfifCdj8g
QEmFSNuZajilhPbvE6I8FtRSyjemJEbeMhXNGKjQSgxEZ7+QI4bTJ1vhFEQycqUC
v/T5ov+vXTvpDRAtjDfpeIjJDbvFuAYTaYO1DKmNluCJIqZzt01uedDbfaHRiLu/
BcFgW/fqHnRtjU437ATw1OQp4Dyg9DNCOHrF6HLT9PTic8JqhZwvVAvIgZjlQK8s
ugDPaW2ujrr4Bps48p6J2V+lKb65owXlRz6LB3iEORpQYV5wubEX5jmoyq+fEdvf
Rujisrbo6rI3jUX7Hj4EbKTGYZNorzlzEhHjNJcgFKHD/ZZKS5vOkl0dP4//GE3N
ydz1jDXWCJVBHBjt+uSexFYCD4zM/uSQWwWiZ2/Bp4VbKeY66J6gvAM2dmeUQV4P
P+tKuAlSFLJ3rcZYgEjAkuzlTwW6iLFJMVNCA/Y9EgmZZhcKEIFSM1FOEPj6nRCW
BmQk5XSMqHsfkiHqY/NW/whWlVtgvfZiXWu9KyNx866dfmHhy/lZnEfAKj3Hv2/u
H6EbOVe02HLXHJ5jg6Q3ulTSGkrkjOUmGu0HfOF1a04ey7yThBFGvOuWzNHrxDZA
l6P0o/biLZcAytxEuprFvreG6qNxT+YHNCTqHTM0Tov+lce79wkHQNGJunikbPbf
aCseFxLhXZmQ6sqgiGCwYnvYEjy0jMfCZqIfdWd85OMOSTXPPHbVqN/bjtCGh7DB
obEcLJ8nF4GLpDETu7mJQaEqpB/uz0altVzAEbokI5L02srqn9bK1bADxN+cYNPT
6PyzruhmHa/j0SM8VUebMZTLG2G4VDLz5Pk1F4vpZ1vEdsKC8eH6KAkIbRm06Elk
WLBVgsmOv9TEOOBkJ+sOAYUMFulKU0sGq7ZOj5TUSjM4alIS6zJxVsltRd8Wmqs7
FzasB8FgSdk61oWasFzL793GVyFto045ZF6b5GaBSW8N6kqRdwqSccC64QdUmM+v
s/dQGd+ur1ygdPD5Co7HOs5YDOnef3MJeuKUoWeoo0rZM2yqBi/UjVfrU+d4aTdv
Vx9UtJ2d4VdLlV/eLlR3NaPOFSTAVysEfUsdho9FWkciKgmiAYpPhvYOy2DUWwgs
MAe+tMAejQ5RBE17qYwMish5FsEKKaZa662M1ywcFLvLpuskkjMLbZpVKVMKeu9k
I2PcVkWVtci7p6dthpHSHKkifS00dtBIKAabIosKQQfwygqoFq71omtP6yha7sYx
Dly+xndxAdk1mep63SJXezFm0WXeBlxjSMN+Rts5glStZtkW04gVk8wQbIVARy8e
ZUn+mNgo/A4Vo/LCNHKXArcDuvpQXkAnOzR8QysdzoYFC1DnSbzW2nMcI/wceTT7
I+qBKFU73Wy4vBQgqmFa+mvU7bjmzHEXc1MUh9p9wVjQTCaBD4RmUO/dztawqYmK
tV5zA8uPm8V8T5nkS65RqfmCZAvo9U2W/fP0CiMqYgh3qr2dXNQfw072k68+XaaN
PvPKKS26iVxR2DuUeq1qbTK0N0ltP9w2raxGaoE/h24Ga6aCTvkkT37tzRpmzh/Y
EXbwJ38AxrcWdNGR7c1uhrp0WuGIW2DCLowiuG/T6J7vHkedvZ08JmWkhJZzs6Nr
Me4jBgOU2AclKReacuBsKNIiNTze3/sr3eKJaryeE4OKYE+HTmQ89C3ckjV0TdOU
NPHubgpBXnaEGdoScNxbmU/npGRXGnEexjiL/LKOUaYjyVVTZgtwfvpVz5HwgyGs
vjF86CgpRh4kVswgXLwosnjI/fxCL+EaFM0pNJSJiC9q34G9nLPgOKM2LWGXtkGd
suVo5ge4l3yKigesFn9imdqrilzJu1DnnW2oQmcDUJnMgSWOjEl0+Nku4pxKJfAB
cTHOMs8Wvc/RXCof1M2xFs8nivyCogSXhF6sR/goiFcyoxvj186NjqbssYPL4zgS
7lQOXr7guApNrhCKBx2qbJQdfVRE90o7TVql8LfjMkSSSdAvwvkK2WNSjPOmIeij
OBY9U2olEaEuoOXIm929uUAkXRdigmLvtnRDuci/VBLwrHQ8TnktUSQhMBHwVXGo
dmpkuFegNuNu2BDrcgl54K92NBj4ohFUWrP8QlyKHjZavv8wGrNtnvLvjjXOmHAv
WX6Onr84z/oAmdsvmTNWA7H5fiD0eZy5ua7e6tVRlHQOcUP7A5Lu1h0GozY0sxfl
T1/Gpm2BD4xGp1Kl6T4h8vm5bnBgL+RXggBHbhQRjcNL1NTkjEjprjJc4hHgIL8K
fsJVEFZaxEBQfdGK2aFVRyGS1aD7o2D0goAehQFfFxT43EYjPpQTZDcBDuMfYcU9
zH1xfSJHFdkx3miCnAucapOuSo6S9j8Q//tOb293DepK2M6weT8cHOBwIBtENpH1
wpTWAMRAiKpjZGWMxYbyT9DUJZpUaq0zIH4aaMfurAOBAk2wriBdr/MmFu6VBxVV
vWtxmedeJcojdDVnudlDBA4LQevWj5Hc+mldIqiOoEZLofk0IH5pHPdQg5emXIeM
1ZYh03zndWO5zjTCZGnanB6imBwG5OmatcB8vVMOzp1mB6gn9ww2bp1CRM+pKDE8
Hnk8yBe+w/UtrrBIPXicA47DSzXH6oJSmMiQ6fC6RakimTg+tu2IvhfnCfR/uP0m
57qdA4+bXsUEGLsCz/fPoVZU/rpWH86zez/L1GtsSKm2+uRMCwahN5CIuPARKcU0
t5dKz07op+t/Z6egGNI6DrepHkkbZ3ascGVBm8RvDoAmd8ze25P3KP0DqETQDJqy
FE9zLW0eK3QAHo5WE4KM7rQDFhhAfDQ8kV6YqogZEu+PgITJ8HYI8RUx6Ftrlyel
BXaLYutBLBAuDtWxlaGju2n4xQ9hpNxU0pIde3k8jUNOqJPeF5sy0nBT7KHHaSkm
3rVJSN4N8ZsYoTzkqYKI//wGPX5If3mE+QuHzcpU8xeZLF0pZNWqP9ssivN+Gerw
DQfMK5swAkqgrnrzU4+GNrGqC3+/T4HAvkr0Jc/rpdns+uqn07KbhC6hgzF0Zlpz
5AqVxcLfbAPmhrTnbBqJSt4MbINEBm1yK+seFzUCGDFyM/3KjzPX4kizxIDfu3BK
f1mQAwmDEzDp9Whs8NtqPZDGw7wIppwffGhS1OHcc5h61oyWm/DruNVIHxgP7b5c
xzm6U2MXbA6Upq9JwMyGE9hQMPjiDPH9q2ysUAs1zp5JmRjigN190P/4R9gWxEwZ
3Jpdu04EsSXJulXPX6baK3HAqvLIymAH/4dfkZkd+9iEQaPCh+Ux/jrXC5r2X8UN
7PG7wai41GZaTnmunwe9v/7+r9h2+VZO00iGp1u0hNiLk17HJpvSNUNm1af4JVuw
hIgjk1/IfLT8G+2oCJsuhQfLVQ96Sj/FtMox4R/IzzdUW/i38H3LMH0hICgSdZX7
Dfv6jdVqpkDtAcoBJd1ke9IQJkpUNqr1HDaDluCCxWNbq058JDP+xqYFI+6126zD
6OzWboWohJ3Lj8eRgMGo4DWRJk54UcEO2U6QjNd7Yv9G9V3wwsz52hYuSBWQwM7o
GtaPHxPBz3i+FjYElBBCmhNqsEkMtxqaIlRX2MvSIDaVvDxn2g28imh8qDKGJ6y8
ZpG6bjji4UlwfSEGyiGAZMz46HHWPPx1Z/yOqrTupIypeYoCzn8fdtAzFmJl/VE2
l2UjK2NW58aoVNwLTBlUblKunkbiFAugIMoh68tIsw2ocBhejuOEZYgloZXzaa3x
h864oCT9/f6Lcun1n+4jfOclBnBXyVNSQEPv1d1LgX42cswHrNT98fZskihPP1Hu
qQOkFxG0L5NqhE6Emuz9SFj2/R/4deaTlMutArtFIFLEC4IFWvKs0J9m0KahKFnt
mm3ISRkVE4QfdjlpYgW1j7iCqzrQfjHqc6MJ1r5/F0JLYOfLJdgeI3bPUa7KWSE9
BVzl13esY7/I+LvidVV8kWOdaLh7jputY4J6sz/zoEuGlPCeCJBS1R/w8kH+umgv
T67ms0+Y25af6MqGNPxTZqOiHcqj7LkrZTjNs4SX48K0P6we23znhAj5Zppt9E0G
5+KtZNJEvvIObevvgrMJunFZrk/gxfV5RrRkD7whl1wd9b85ISEcukCN7eYpKgIo
NWCPkiSmn2ygU2TsNO0R4meeA3xrrn0wJ7etac1ziUxhuiLNlng2daREtFLrFJNd
8ekj4s0c6AIRPZfzY+DKjaAv3wYoU3uFWsYTY9XcCqN+cEKFGYepPjr0VeqsiGBQ
2ibhjB8yxnJGR3eFdeveOUkUdoHwHpCi2+QJqFmLmzk86iKxqr8nzh5bwL88H6S+
9qhv8QsDok0Zw7DXkxY1HI3eHqqOYr6lUTP2dJVNgzOLqCVer04gucuxETMyCDZN
yrni8/o8b332ug+zME6vxOt+6lf8C2SxmtPFBqoi6Li2k8k36zoXJ+LAG5rPil0c
ivQ6N/hiql5Vp6gG7eZpSRXIzilqxeEult0aUrrge798nKrDg4MlQtw38RCJXLUx
HZh77YRhPBWrMzm5zs5CYiShSlsdE2Xjk4F+3rs/X7RDq2Zn1DKok+ERKWieRX0Y
TcVWH8xLHRAUpsJ4EYo6srr8ZHA71v9w2bJXT29kEzVj6n5G0jZZZWSU/ubSMM6o
uyUVepnTf8EW+iMS5nG/Fbdq0SYbzvbDxIHkTx/IZGtPIgpp2KjlkNfKH5Q58G5N
N0RaIPrisULxiqtSIqX+zP4nzm66OYKc8acumxvHPW/7YCm183MBB4UYjN6GDbro
e0H240ycuk6QyfJS7zPJpkY2LKU89+BdfLliM7bFJWgVBvVjfLYLkn2yOKoc9TtN
vWdCEC54Gj0eHPfzU9akB95v4SwgfWbetNIFqp19vKiTRa1onvWLUJ06PKdrPsaH
PhI+sQlLEBUbIoy24O168TWlurkcAQgh/Z0BxJFJZ3v+PcdeTA9YV9Sg1uO8JVFx
b13LP8powfDklvkSXLrXckn7/JjOaLJEsW6WW2fY0IY29kcA8pDYt13yFeGuLGCC
UDRH+QijAs0f8OWIRMrM3rObaX4Bj1QcYDsG669vGEP7uOtObhnWo7y4rNd2XdeI
eTiuLW5VKTpjgpjZc1q8OCnIc0cflkIpTOi7ZfLgLwVvD6jsUffo/nJ6zwIA5NyG
0pLjvhmUk0/Q0CWBZXB4X5LPUsBFraL0KQ4zHL8PDh7rozMr09szbr0Iw9BHfznG
mfK3vneMfBA8pxThoP6p6IhCfpjkiuwpORlrfjRQtOokUfebbVXo3KZEBsUOAnz5
+FqF3i5QLr/g+NMXPEQsJiO2vqVRgEGq/BvOJgcXdqRJqhatJbZi3+/HNWoLFOLm
ittLVotyyDzHdQg9LZ7jnREu7G38m/XmuWvYIUNDeXoWAUCIlXvyU7zOSKMjqNZa
CJu2tfGSJX8eh8aWRtJaQuWg83kX1kTkfFJdQS3dsA5S/5FmMmoO5YJXdijBebcd
UEf2ZgXXsnxXAxMZ9Gc6PaARJCipOWCcwnRGk48xlkmp0ky0rXqYqm6wIAvz+s6Q
1lMOE1fSSLIE0wqKAGcnwfZQOT8qJO4od+UkDEyI4vI5XW6NICDtTboQ5XIciKaK
pXg8XW90sUwacC9SHp7yQYt+qepKzXNfTFg9pCgsW6FXAF9mIEcGrQyPrGqmu7vE
1bCewFFVzIQTSL41qL/RytLnA58iCGTkNw62UZPWPqk2XDYBpQQillEXoHSp6GAr
48/hFJ/8OSN7sq74Gw5lRxLxwrUNB8HytkUGNqqRNujbd/jiSeyOL6ri4C2XxYGP
T4DS/0751gfPH1IaohMaJQs/+afPWWIkoE8LxfM3FzOq26ZFiJrTh4bJ+OGVtsts
TSJD3uoZgE59X9F3Ja7WFH374KFtqCm2WTcUkRT7uYLPjiJbaZIGzYL7peZQOI25
MZ84XgS2/zSYpUNDdo5v1N0VSZWOCOmvnynF40PbWvGL/qQbemlLT4h5DRuud2+A
aAHW1IGFM8tp59ywDfnk4uiu+u2aWaP2MbQ/T5VCWkxyQydFiXcDLpPEUPm9P26W
FiSklpZvQPMW2vBlazL+da7IazrHheazWh6QJNyH162Rc3jcyG4njvmaVYMjI7F6
Jbfe3EYAXtYZR9XT/y4C0nA4sV8Q9eyPTLIsqTRX7QsPiyPjWPrqaFYhi2tEV5ya
yAZsP3tjRm8cqN770LyDtJWxGgNx4P9ARlR2suSbndGS9TZhM3Gxu2INceQx+6HI
IwYKJXRNi2KkgOfzQSZV3ifuPjTsQuyKMuW/cHpkv/2CJ2R+A2X4ziaaWuXqcjf4
uSQRw4RSnFGqiPwJVoTGQe+0qWbph+8Ns1HDcxF+jR8VxYHN0dt81+UYKN0ltGZw
h85c5rJJm6KVehN2UkcYLoI074UHEp2LSI01OIn8VUmw3gC3090YEMCAZoCmYw5N
TqmG7+Q3qtzXVC8uQuDtgENC+faMXNE4fQxAuqqmG/0Nz4j45VRoL57O+hvHOa2s
r1pGwmPf1yQe8HKzWv9PWZSleqIcgnmClbAk/kWMDdBoTAv0kumMD3d0avgxiGPa
nie/c6ucd/xeI6XEKiOrjcQFKfrOFBu6OGYFeBeTkqBdT2shd524lYCCFP+aaFH7
WAm07Fp2ERgtUD9CwwZHv+4d6NFFUFCU8Cc7wCK/WXycJGJyydw3RIowTUj6cjfw
LZa4B7XU1g4nra1o9jMMd9tgeHq/oG1YBfPtsEkc/BsydPYjrAZ61KSKj8O3BHB/
tTKsIMyXpsgQO61LFqBNt5+XhiaqykFXiv99d2gvw3RPFhLo2D1OveBqyOa5It+c
O2W3zrfMDdceh10D3nhj1D6DX7+nROk5Fj+vvZd6MzMlfIE6R53yr1lo7pVcwqLv
idebjekPFM1TRe1mK5B009f+m8S7Pzi+9H6EU3TBs6lj/hAsw9heq2PgtyiZ2t+s
MAzigJmipuxSwk/CTEw+uZ1OkAbnYSvoAAFa1EpTDV3upfrTDgR+TcsgO+fmlJk8
/UTr0StZF7/icfqAApz90wcSfXkp8D6Ywxj4Fa/1z5uBcgxcHyBFFKOSHOQCCNc2
D1rs7dihEP+uJyat9bFKnWpHovrXdKcM5+0l3S8as0ztO4mvtYh8YuDj4jKdjdF1
MQS7O6sV5yQmmGDjET2g3lLEOcxn6xdCh9BQ7/BE1u/iL7I9JTSRZDubhfr8w0vi
SSiL/Nry2yxVLQoyAOFFkad9EDKd0G9nMY5OIRBChDYTGs0xFEQq97xgUUBRA7b8
5eEOxFepBbpt9Xvnnxmt4JW3kEcWQ+wLaIz3/tbuGjb4NdYvJqY6RKLeezWntXdy
JIzi1izBKwZVIb17pxde0lC/amMYIAqB4sZxUw1oM0k2QVIGSTuAaDR51/DE5Emu
aEQno1XBM2s42mIme49Q11CZf0xVrcHhf+HSAfKxdomKnrItxeqgA4zmzR31VJxN
lxxtUmqa1GLp/hiLbGCltGeXcGZusDLWqqyAa6amJteYEP5qX/Tn2C8PQmraD6hV
ppC0DMmSdn2VTI1xp8UJt9rUzXMgRztsZewTtkwBXA3XG5A9KruLBEtD0fwPIc8G
rK1Ct/ybQlvIwppdCKKJ2lmDRi2H80evSfjt2MjmQQkTKk4N0HGlwugSk0AiVQBU
CU1Zn8e5ysc7KrZHHe2QVrto+rKfJypHcslCKRofOMtKn4a/b0u2o7qaFA50f5hH
7vdCZb35fsdWhHI+1rMxrhVKuEXMYbeJOmhjNildpYXnNr0labwD2siKDp02CVeL
gDADMxfor9ZIYLgvuRiPMJomtit22ioP+gHI22X9oNUkSbg5ml6g81c+FB1h7vdS
PiLaVN8jMkARFavmlNol7WhiLG3u4QqBJWNaqjk6shcI8WlhH5gU5P5jl1kUwoSU
gRHkcVAWokRE6DvARbC6cppb7bRxy7GNGz6w2Tddwk2D/JUm2LSCn0WjCAa9k8G4
y55g14bVx+GRZEoG8gbfHo1wRY/A9BI0cnBm92athXTiW3kkCll0bcOENr85bDgn
fPEknywMcgFZJ9qJHqMQwewfNCObVeaW8Rh1hAAkJRwzrq5pQ0jDpHV9ehejGMah
xT3ZsKWgAYzPjHKg7RRIGTR3Bd3wdCZeaH5Ln3ivmtheV0HdPF0cpPYykKskm4VS
xfrqwpGcDhzhXY750o+8ZhjZmmtUJUBASZdeURloH2J/Uk71ZEp85cknLL9U6V3c
rKI2nyOkV2hir74+xqc3PXOEdQ6uGy6gXFP9xKbjK3GmYrh1GmFpp1d6r+4IJJvu
TWu3IfQg+EHcBkzk+fEgGoCk3Poq3xq6afhffAe83eHuDZF3mvVMtcFXnWQhZplE
1JBs6JXaDg2XKj92MpQ/dP5QkDJe6uRLiG54mtdLo3J8Ablw5dYfYTV4/XMNOVL5
qu2K6Wmy0r5wl3SBLFfKFy4yYtf9vg4ig+7fazZLXI7c2PMuo3hs3kT/LtzZmLhp
0nXgRsF/CEV9nkaZ6LTaUPqFvaQRkwc32KpQAUQxyZjVJVRI2OQ9TVVswhC39Sml
eCXTl0pltyeLO9rZ1ZuWo6fEVNXvTEJp322XEqpkSfLupQQqEEc/4H/LuT3WOH0H
S/5Pusm5sYhLkehKDWvd3eLYdLfgM3QIbaXVJjjvwKe6IS14mv+rVXNV+C9OMEPC
wuxHGemek7VEQNk+gllufzTfTRhK3y4TyBQ6olQOYrpmCbRBCcW/8DCJSjaghyWl
7ZimhI0+Wxyt0eMI0TMjeCgT+i1hHxX6oH0KXCZ3d9mPUX5DYVqQunNFsXQsRSYM
5UVW6YxQmGHbpmA+smSR0Gp0Lvvv1q9dBGhiIhgDIMiId9+VOZ8eXFM3rH+bmY3/
CGhYoNATCtBz3q1FaULU3msDYWoGC+x4VjoCZd8dIZGECO30OSSvwBvJA+3iKAuz
QXwc7Ta3+NQR/+x8mcv4xb124Ql3YzlcWVPejJbPGtnRj1P4xtJCFyQNapUeNLBL
f+B69ONNxLPk8bGfmqQd1jSQMcAdEiIlgcSeKKMCVlo+ombYCvuXRilgTMMBh3Ff
NeV68FtYB+1824Mm3Ps0Eo0VRz9aXlvjxcrJaD4SjgE5V4pnClgh3U8TuAMiykHI
Db2H2RYD8sJbC7//O5eCwUkaW8oZpPM4U9mwsJc3F0a7bDSV5uwJq6lOp+TkO7+7
5xJLpajNCctLlEled20nrUp7hRtNp0SoIglQyGS5szPYft6wni2sxRfmKKSPHUfr
tuuZd5llogeJt3t6hBJFrOwVEAA0A2otQVlB5CJwX/2UKpJHeaZ0lM8f+VbF91dU
E7YWLOQS4X5CBjm2EczCMmz8fAaBHVItrT8O0p6WefeDZFnBLRUDwV9KxTmKtvOT
MJovC+B7/q3rQSUNkjdLU/Q8LePcDPenJ1B7Vv3aStZHgShEft7mKDNC6fGfTeLQ
5vI8PAoLJvYKgDFjHRmGhMDrIaGeAN84oh1IoPkpbBTaP+U9ET//e0Bf6Bw7kTvF
7Dy31K1J8CVQzzUhHSuujVHsNb1IwqHeCgQa6LOLcXJ14nOgq95eu+G6ejoVQGoc
SoK7k6vivzL01LrathBr43U8aoQu65b30ocg1kqCfg5vnTPHLlYSgRjUEZATWiIe
5td/XZnTmQ7zuQonTjF4zd+NP3sFO0zZKyhdhONgeb4up0sbozrnfS4rRC7ISZqu
9DZj0pe3aKuNbYCOP/PF9vuu0QVNDFKvZiDujdMHBfHUH8kSEKOIBi+D9Cyh1k2V
S+B9e8DM4szs/7la8FVnpT1Y8bKiGxwcAeQbQkSkc3HYHFlnTiWSsGm1cxnsLEc9
9lbLzAWMHhv7mfQezfuLRkNTCFgSGEFLm1UjUIKJVuthgr2EslL+o4hmJt5k0yIT
ae4xKNqX7HEvLhEPmWkjmInHsZDbDiK9d4l92nf5hBSC7c5YXD2/ANC7A1Lq54qx
MuzQ0IYQDRChJMD3K6nLSHsa9Wn+Kck6bS14Ne+m7FGqOe5XF5QRbQxc+HJuBQOH
W+phFoUV45tNH9gYmB4NqmnrOoPVG0IhD0lAfXew2G+im4NFrO6lzijy4Izu3JSc
MdaKzJDEIYTq5ok+nPT6fK7p5zVv4yzjHTg3NIHk/2TsYDhn927xiJ0PfjHVN+l1
4edssqaEUQMEFr+otjNYHtdSn9td8ppC+lrg4lczOn5Tti1SmFThT2/J1AGjW1QU
VIQUAlIQRfIn0rnx/DvHt2yKy9elX+B3FBbxBUgQzKK+3jCVMIu2h9BV5MLud+Au
nrGQD5Xs+m4TIkZrkpFjx2UOoQ6NyROofm54IoJbTtrFQ3+H2zN8qpTm3vcXH+Qc
MMk8LTMATU834BGMYLLWvzzAdqK6RvLUfqYLZFH11O6vbdHDTp7BECuFwMuRFinw
N1m1Sqe6vRDf01Yip5d1kZt+xw1bjVzLSeulNcU/MIqKJe5mVg92a1Eqd7OxYeMg
5HmE45ADQb1pJ0vlZO/dTVbYtPk2zMV+PTamlYfgtzX/eyhe7D01G3I/ywTm5kHl
WiG1orvVnZEyW6Aj23ArQuHN/FK+baKj4EGiiD1dbxz5aDLNMJfZFCuxvDTzkQBu
lg96g9hoTh2fZzRgaNQTPwdflESDOV4XVr1dupzLLX+vmwIuYSVHrKzmyLWVpHsC
sbKJSG0B7VKFyu1oNNlC6FNrnsNnj0RwLLCzK9GSIz+r6Bq6GJgtx8/HHFdjJgwB
BDTeYIeV+W+ekWO82UV8UB9JYH4PWKJpsfS2Klwl77Tk9tpEkDNyjVsGym2klNO0
/eSM/kqYuR+eRrSgkDQdLKYgy4jjdl2PEdrImBHHXy3yy90MeWUXJ0DuLKlqCM7R
eGiNzyhHbU6w1T+aOlWgfc5kcLQrgi4K/PYGK87JdlqBOgjccTswa3KEfna5mdnh
JDV44MYSEA8Q1ZmFjFlwURUSKP726krUpplv9hkdumaChi01AsFuEqKWOiihyj5W
MgO/DYRFDL3Ls8KJnhWhMhw5t/63FfSlnwEkWwmkrnQvvIdxaqSHCM/BVFfRV6ZB
3W+pQc38DyO71p0EmYmygI/D6N0ztDjGm029FnpPjGlZElWnRQrHrNjPhoekzV9W
STJcc0wdTxdvHMl7ogGBZkrWqPmKvaSpVToWLRjHDzt6/9IQnPi5sUQrhQwTL8Po
3r17kjdeExWcEha8ooJeLaahDseTm5k1q7jJcNa2eUfsMmI/bGL/2jdIw/aaQsul
az+foPSaL+CRstMDvoJCZSdHCfr9MRBNhe3XdiMEer+Tb6BswIeR7jgxlPAIjCq3
PHKG+L3e798WD8OFBJx24J3Hl1HS+tmn8t8FjZhSc8eexXb115Ejo4+GKXADXlmK
9rE6hm0VyJNMgKzAmAezPDRGqwvzB3OFHCKKxK3QL7cn9VzutjEfRB/X4S3Yk3fX
Ev+PeDuRLaCT+by3u1sZKhuqr+Hb044eMvy49yDlRUNv4PEJENu7ttzvSKvJ84BU
SuASzLU5mWDhm0FcgYXS3agPnT8tWyXPvJmOLxDMjaZoVAXwVi72z7Ml99iRHDg/
OJLcQxLfRw+Mrksw+nB8Uen8iLxWI9RpQHSbKIxN98jXskMtg0Rmu5kGbGPwfD3Y
9w/gC3AHFGommQKXxUOtfeUrUIl0OcbukVnIyxpxmSlVEFfz8gapBzBB31VQxxBs
6SktbA30EmgURzdnSVwwvBJLo/y6Xp9LjKXOJ5fCaP+9Tr4QsnLPa9MOLUv9SIRH
bU0pLfzDmfJ656z0CiaPgTNJ2+SpPpk0pKkKaCNPgy9t3S85jeYrVg/MKX+Prhk3
dFNpV7L/QS9LVs8X4uaxhxEcZrNeHgja4QF2jTukS3Pdp2cAe89GzR/y2eidsQ4N
jlzj1T320J6+s0IOBI90Jlas8pRpmorEmFDR/DgyqpusVZKOdYAhHTw6ZQeQMDct
jfslDGPiov8t7JUZMERKh4boBFRZO75IvaQUpuuyaKKzEmrx2T+MR37Xkf7E3tsk
XjgivceLhNGnxfd8byhzoZzcYqkVfZJymYk2tReKUcRgDzWTec0WyGwhE2RbuiFz
MLODXgabKnzsfwSKWx0bjKBJy8MU9HLOsQ4x+CSX+V+yI3j9ar4GljLZdtNhDWAW
pfRiMd2dkQ99VnQ7QnOjClX1qJ3Q4dIkUNVYa2Mf15OmrGC44jlJB2wLJ8ywgJXr
ncRx0Dt/gtE0QjwYmYcO08p3t/S5l0hvUXe9IB9EQXeb1mcCkY+4301OaukJLMa3
yg+K65wXoAkjQhHVvWPwT9ZyjGY4ljd5XdA3RIpZDpEMpCztgrmkPwEEOnSPRYiy
QHqwm1HRuREM4CGFee1Hm+UgYrmzvdcVyjXCGDma5qTi6D0JCkaLbSxVXjTi8atH
thhwQ1jyUh1kr9OqP2cVSn+mAv/UHCXQ9WIOOkpyF6qJXxIjwym2r+9ZYPLYZHSR
3x5OpBzOv3oPBrI5p96LpwINeNt7DKxspYo1HorYLE1oC1a9qmWd5UH+7GrJqlF9
KUiCbJ2bgQt6fZK09RtHROYmguZEW/LUv1jxDBrmlgEOGJ0aGZ7y9HYYKQmtQkRl
1lRfdJkygdVHRbFp676m5KvZszoo/27xbRt8uqjtmh9yxSM9c6yJqT4Gsg4j9eWA
qHz90VwWbixiF3K5/NVdc5pwvDi9vhPw9HPkTjR2jjonBZn9rUSQMfTaExfpAX/0
9nsD4BrsjO6jAqqve+JZPTcOjN6IGhNEsALwRDe2SoiZMEGmFMidckvAaE3KGjzk
42XIfvZoND58OMT4/Il5iIu4qFAK+PH0f2ixbZfXYcnt19QeRs27E27gJvrrODIv
7DZDn4Lt62GFtbSahFnG7GIu0GChF7Rz1+Z5eGDciZ0M0EvQtp5ANrcmWAaTyGKj
/VcCKVd61mKtQO9r+gHv1YScvX+OPzAxQwsN5LV8VmGe7X4HZPmIoufvZW1fLP41
OdfocaJkm+PYqQBkfEhDa9fwHR7nn/tlCZSXf/bESBeSDvD0zGQ6DJgcdOO7hwOU
1h8lrWuzR26iqS7IQOyiBpn1Vpc7xc5GcgQqpKDwNq+nnl0WiEZgvdWFjMwMuvhp
OmR03AddHVYk1bPFdSh2h6JyY8KMWSI7Kxk8H9uqzF3AAO2EHJjnTf4XPNIB8RP/
WhOHUNf5YYRL1NCy8uJMXod7cUmF5Oyw4eakUCVFdp6XMAQW3gIDGS5VMWumgeM+
ZJeIcJ+GNckYC3e1tL/DgPbl9rekvrvEHwsyuiizYvAhxiNrQ6SZT0LkBv5lReFv
6K1xsn0rh7xM9OlqhMJpjSrUPvkzITpUSotVrLqo7rISg9LudtStWGH5cs+OqOJX
6P2vRxcY8NywMo6z05UUr0cjg2YjssJzqR5KV0BDtGChrbWxTFqnI5bvaZ8A4ti8
Vs7F7Y7iV+BrX1BrG/twa1hckE8dbbG40ZRbguqxYxgIZAmW6niFcevogwLS3pnH
Pl+w9f+lL2OE8TsJsd6pBxhRBkHiEMMrnhbVxSmncWDZ8ED0yLA+GyLos9PuObj6
K6aaab0mpBNEEA4BnSnWfSrPDCIiTjsuBlnsueM8/D0J8Ifm308GVQiihCAR8y6T
X2GcrGyeqXCBIHwHJEilHv7HoqTcB7L7mDPrvx/B8HQ2kp+0c/mPI7imcPfADjru
BweXsDtLeKDjQG8nNp2O/mfxWdxVREYEQG9tauGUxdezajr2K3jfyqXW2ALLic7s
PfPR+2oQnZ7XzwtRKWCNe839HwgrB61rGObi0879Aap0yLNjGjmjzps0dJYSbbOp
hnfXRuUMINg/9XSUDbJcG1qPHzxdd6OggkmoC2c2NCzsEsgUwpOc0R17EpXGoDi9
uRqB9AYX6H6so/Djjw5C5zcstw+Tavfk2my00/dlMjJLep7qbo9kyWudExEqvmxz
RxAGYUy6Eb4IdMHK+5xEk2J0gt+Mklh0BY55LIG9w1Mj+LvTETncQckwhMylbRLY
c0D6GtoDFsdwrvtGq7z0J5hPnreQnoN/FC8vs8uF2dDEbygo7w97dHYyntE6MeEp
tLWC4KKOldTLkjDUGSJDEUxQqcd7eUFugTSyV6mOLQn98CccRCpkcwswdKWVW80V
8Bn9hXGNDpp8ejUlDzc5mtXSS02SUw8Hxca2OluSaXpmlcEeaE5hlIFAwu6Qal7A
E9KBX2bY4ThxPdJPggNyPDAB0Ro0C2vkvcw8BY0ZZgtH2c/4Eyffp4S08ZoHhX8D
XI736QV3pEnQvchh9peA/hoawbEcS067ALQcj/7CjYfENbLuX5fPapvXrsne6BYo
9IHMyZsFY0IOEm0Hhghj9/SSSXPN7oPT6DS3S6oem0XkWyL79BtghY/Og4DmY9qm
8oWw4UQnheRJZP6LAhcPZTr8SFMvC3hs35bH0R/tyq1g9/aMMaUGFTlcj3lN50fy
1RMpUcYQ3csLVAmSfTN+6B/6FhgJWJ2bNzf2bCSMita2VxQZ0x7ouD2SjUXqN8+s
OnKTFFN/3Liu0j6FytrktFso0UtUsp8fNooZmfPE8Tmch1D5DHVnx+FHiD+AJFSU
kCdpyEJ0HCGo4Q9xImW3SKgvmylKUhsof5zwe+4dxsvSP1grBhYThX6DzqxK50I6
TATIUo0VEQ3twa/sRpya1uW5DrYR94aHh5ARB/F2C2Pj3x0JZZBKxW6q0hH75Yz5
cue50XndVhEcQMD9rYImT2LXg6oiBROvcD6j8u3OzT2yqNM0A9nk2YARVc1FRMs1
yQX+Yl973/x2fJI1gMY+UTlW5uV1539I5AcxvGAF3oJcXzHGyzSdwKL2yiaHamG+
Y9VTT6Dh2zeSLW0zicEns6h8qxVSLCiC38PwKd1CawjflZOHcxj61vaswILGXweC
aNpznW8m8BbiG+vuuNu0INxePeE175x6tpApjoQDyMSupFGbCv5iHU4ba09Yu7cw
6NV+grg+EdUbwgklIhjgm81yqqkjS1G3LSC577+xw5cGVEKNAa3iDevYwSpc6Nwb
Lezw5TsgIQOcP61as/cHIrKALVKKQvdluUNYoOr/Ljzgi1qnOWGHYTZ1xCdDwUXc
b/Skvy6WClHxCBxvlOuCFPdftBXnUzul/r/NhI8yoaCPhgqTIQWcDO7Dgco595xt
Kitf/qBD6I8VojU9/lPERNS6TBToTCb1wnDwpVvQjk1FriiI2U0lTjjalNxejmAa
VkQgGjtMk0ZM3tg8166b7ZLBx39zpw4fKe2Bw0ulKSrkwAHOAlLIrJ1hD0rAGotp
GGEktKSeBq17dRFaoLp+7rptn1v8O0xWbCfdMO8cPLDBlS3XEL3sZgc9o5pdWkZP
A4tawLHF48c8TYZND8Q5mNgDvEuOvcEd5xMGdZFjUtCpxQLRnrHHjW8vfZpOSLJQ
KfpdrM7ZcOdSjK+JOSZbAcsJcz7ySdX3U1awED6C6joynDTDra1Yxn/rzI2/4zbV
9fEXn8bOFWOn5gsjp5awPmxd39KeOvTQayj4OtIWRTjguv2BAG6lqcc4rMH96Wm3
d0EZo9+9C9e1/zlmeWVAF6oH2Ws+2KTadRNPh7FuR/9NJOM46lRZRnulKIQl5NJ/
A/gQucO+9PK9yeK1p8BL+6mJjnZEG2HawSB+VfCZFpFa7/8x65HMoLYvAsGjDlCr
gIWRLzl+RocwOX8qDTEZp4Ty6NKswbxSMHU5UVOvr3mLHkfYMT22cH3BbpzNDdU/
T5ABi2UOJkRatdX4zrcyyU9WvAW3PaR30Q3nnulUZTg4FQNPIjUJ1l05HFWBasGh
bntwOG1n3eLTA0M0jNtb9fGdM19vX2GSQiW2eNMwCLOb4bnVHtJPfvga3m+WGqZ0
t7ShtTiGddyl/mH+czOhFGh74QMKBEM83Pk75pK3BHzClp+QU3UfN/NuVB39Y9Tv
jMorFMKupLQdvI8uaPnx+4Au5cwsEEZpY00q/dlO5Ts92iCrY88kEjXIENfj6NFC
uq+9cg/gaqSXcCXy0G5dQzAc9RzcZpnMbasmnO/fprAdnSEOEF2wEvtC0+vMa0UX
ahtzS3tr076ExurkYknVuHCENjFZdTpVzXxhOZhX85R1ztKEQOGn0V3m/XD/wqIC
4jFh4pm/O3A0Gt9MM8CUMq9nwKb9rwWFOpsjZcAfoVkuAYbUAWQJ/2MgiAZ3Pzvi
o/IRL2GRI7XqLOslFIC/PIx5HCjKlxM2P2wRkj7fvSzDWI/nBrQ0gcPMZHyXKGhL
wlhOM0Qz7cts4zvRu+vtFD6osQjxwTvronSiLWKwQ/eoFnB7fSubMQKM0yZzhKVC
oKMqWT/H0DWycu9oFFrS01CdS2qsokZN1njgwsvcvQbPjNlcYuoKqckjQSov9Z28
/7mqrAAvfZ+09ARKSlqREFKpt8Leu1YWRjdjnn/wgl12hXBT86PcMBbJ9fU6pLCB
9AuXoiiaUzxOL59d+SththZSPwzqeEijhTWrEdhfPYPTkp0/NAxsMInoy6ILUuTI
WflPYv61nG8rbwvImZOaNH6sJorSCuQmLZqT3u5LGa0OToEfdu0fMeZq3cLjdRdQ
qugVl9QXxCg8Euasl5yHOyQKhryPsmyCBB8mI0cLTEoSZgzfvC8pOAE1aR0F9AiX
P8XVNCzCd6tTs9OPTZsI1h+7sqVkwX8VFHXd7xwkZCZarNSXONa6ghxN+HYCpFOH
PK44ugy7vED62mg1aRJKtUTq98aYtMKNOR3mXFdtP+m2p8GNlw5v/YzEkloKuIj7
2F3AGEOW0MQoWNjZkznElkCVITyst+wrTEhQI0pCn++SWSSWiqz5kTSlOtNSUlcW
8XdZijccqFEZ2bbpz9cRKxWGCMm48HmH9ihnj+eOA9CXuNi1TmioW/PEVIwEXfHm
mDKQJxzU+351wtwNTho0C4czIgDXW+PnBZHA4UvZpzJDO1SmF6E18e5SQW927alv
uSvLpqYUSc0igqjSy4v3ACUmx4ld6sOAdlw1XjwK/DXHYKAng0LWlzwYfMOuUfVO
fk952nOR1etcq6Qytn6ILZ/Jxg4cV9UOGAUCjmvrW5WzAyE357/QN9p6QzI4LNu4
bd5pLGY0HSOqY6gR3XYUaZwe42m1RGV+YQKgZwrP50atQIH0QEQwY+upNxToO8X/
12Z2ZnlC0N8teHBBOEnp/jWibfoV+I2etoO3N1WKPGel5ltKmRngtpp+ZzEx7C8q
sFcGgWvIJIwm3PTHYAM8Rc9a2NSrrAI+kbLy919RoTvZYlIR/SjGxWwT1uJ7H3Xi
PbIbZOqoaL3Q0VF5skdhj1RA/jIRwk76jWOOxT7NtCN2yyHthRcceFXlJmgYCWVL
Eqjt9+yqbpzUTq2ByQpBxX29fH8C3khDfklOPJk6CCZ+u49UC5Q3ZFB+5EPgq4mE
518USDqTm0EzESW0H6gM6TabppvAk8JKXrbrLBigG/LQ8/sDz2rVMwuyuPAeJN/6
qBRd9Tud8VwrgcPk4PQoQRBtTTptRjgtpMiutHWSk+oj0SuwJapX7T9gUoApnHwU
ndIVKYbcXZRFakJ+whHJCC7L8GAPq7NzbEmFML0PooCz1pvg9Y2A2kNVFpKSpC+O
T22zkBFR0NW1k/ay374t/hUYjRWQWPU4MguKf3lAulwGwdQNyhcwMMCAo5NYdo25
TXypr9SFHSOrguJsT2vM6tFK6Of4SSTdMoec91e00o7AHivHEa26iuX3L+GeEgqW
LMITbsjesXZCibJiQK4c4x0XGmkA2iYnZgDnORjcsH784MuhdaRxbF6odR8zs9nG
yKWoGAu1aiSBDn9ZGX/LH3P0Yr453S0S4umWd5VnRMUYvmgAl53XKTAw0glRJtYw
xm+oLAQaytDry5WHw4R7pcYhk/jSRvocIUTvKacmE3x0ZjXrIL6bMpCOd7ucasaf
IaefZP3ociv+dTSzi+t6egx2xT4QhnVnRZVKNrSWJ0KfxtpkcJjoxIb1GdsBsvNR
OuH1hfvqsdwdLwr6jNkznv7ZtcAJhiE4cZ//dTh0LCDJ72axpVL/z1CSzCIjZ7Sc
A+zd3/Gwho0SgoGmvtdKgjVPyGlfdlvsiSRpqV81SkdJFgtJnf/96gYupaJzHBSP
NILrDGK7qWmZDhzLeyHKs06Tsqnzj1lzmzCavf0I/WopiiYJOH5BRb7oocCQwYyc
mWEXTdkiWUd4ofioHcsT9Fwoxt9I/lD62EQH6WgkN5xYvQnZWUrINnXhZ3QLqJ2u
Rf0EWgv2Avb4v0uPowGCYO/p9/IavRyntoIaGc+AXRfdaaL1+zm3MJkA7P83JEIi
+r6t8Jh5hDjNVgMrm+tdOARb6fftGggU1iDt1HaXUtX4+Vr1ghpN4xLloARyAiMQ
c1s6F/f6lCSHpiG1vObKWcu6Lq5dmynydR+jPcgVza7kLhOvz5AfR80y5IBi0gfN
rl0yptPqpWHpBxgr21At92qT6DlyRVCmcspwG4IiqDaRrv/UM7kU5o4DKXmglHpo
E9io5grDLXgPfEyAIwELQnpAmn2fA/9oaQxdGqXNkwi8I2JlnbBQBO7I0zl7xEjs
KOBTVzWFNmOU3kmiG1xIvFeShN7E6BlT0oyNaGDKqR3WVGx4I7oqmmS0RqyoXg/M
YnmYdv8opY/JoGKLQqjCoMGO8wJF/kQPhzjSRLENI/5fyVKhv2q5AZMssSu2wSmF
0ciCYOaC0UZ+rjrkqyBTH7Q2sm5ZyDfmiqlbtKjFz0YmFcNdaAEWKimvzK94tJ9D
7T39btqF1AssdU/Ufb3R3/0D4IzTynpE9oAllfXO1Mit/JNY8FZCG/Fef1+upWCX
XJf9xZaJYaI7ZZXgDEdT71ckCD3wkchTnQHjVAOb0NqxvBNehHf4jSLHfywKO6jl
9BAB8Tt6dYV1nruTMZMlguXYRha85DY5Ulsc6hEaP1NkdCmKHaxorN6Ecvqp9sSt
vIuI8Ntdc535Bh5/DSLTuWikwCdDMtffOUIDdr22gzNfMRqra1pOL36BiMYYEZ+F
PohOjelnaz5bVIKDJ/sh2ni7CIZoOK2SlzR9VeDwpUOym8yGqtfFbdzC21xjgCce
UqFB+0y+KuWPaB+wIFJeWINEGgnycS3Bf3Ukll+JlB30BNk3WP497uYsU0XQxc9h
1TWG5QF6C99QlljbIfJSXQt8NDybe3YM3oUvONQmlzQX/PWZXAWo6SATRo576OAd
SF4AOIkDLr7fHB/d7sE4+fbr/FbaTslezaME0S6gCDBlIa1wLFoeEnXIXX3JSBPc
cHByZtZACaY5ZSJCo6o68WywX+9e17ZYsCkF+IRc7ap5iwNOgvq0JL4GKe7zoGf1
RUzvIJpGYXnU4eRNZWo5liO+v397KT/uiLWmPi1iM/YWzch5EKt9P48d+vQvNhNh
YuMV5lbMWc/jJuqsMK+UGfLojWRZ3V5SNgHd71yoblrLfjf7+ZE/Amthxr7eOCTc
EbBOZhHcUm/jZd/Lhv3IOnxVGpvbovYG6v0nbxXhRnxSPjHFATyX/5c5UUNeh+qY
p8dVC2sIB536eNiTpAOXdxQMUk4g21rHCMs6ejV4EFy6YccoutMBoprIDQpt0Xue
rTLLgOCRuaWzdAdLa8AX2d6OMzuiiAB1OraQpuugwHZ5yGxg5t8F+mMSu9tJbgQi
VVIBgcYJICQExjqLRv+0p8ToDxB4DTw+0yI/hFZxoZH7JJ89NAlfeFj/SPzy1D9X
G6jhHDlEMvjx284hbNBp+Gv/G9F7roPF3PVGGya+nqrPGR6zoKe+MKVHwwNBkdcF
T2vgfGpRQstiv+P7wu5vQPuLugfhJG0vVF+RKAmhzI8+BHRnmR+2sgVupG5dJwhg
1lir+ob2hN4sZZDe6Xb+E13U8QW8z815ZZvpGXIGplFQHOrA0WTaUL2rv/mBB2yH
vZjocvVgmON6vDPFLBs8I12p/qp6ZTcyUjJDdxHRQ26hPXhhYRXatNIeLyBfDjrf
u9pYQPL64WuU3OwSkKkpKHUm1g5XKkYPaiyfAh1m5cWMxwW/XK1gLvzoCnaWZib+
boL8jugtvpwBRaA+luAu6aI9L67OjhNh+zMJChH1NFxJNbR0NIMZz8q7eH6Hb4D2
IlF5ibizHmbBEZ2Vc+PImKJNhiJJfYz8CfupqdJCBM6e4QzFtqcJcYXytFRCCd4K
8CyuIhMB5OsrIHl3JSCiWONJtxn0F/Y9u0p/ow7/D72H8D81hO2CWr3rQE9GP4fi
8n+ED1ZAwAJRmdLtXp/1lHlZ/QfDX42mYQIWZ5mc2tUvknYaaVNVLk6UUBxi4xHy
QpkDffKSvJhfwnseYAmprLpJg6Rf8CCXHI8iPiyFt6NZuxQdmG6KhXfoCX0ubmNL
LFDvOWjDVo0Klf8w+4pY6BZuCWVKa4cwf7woSRUa5IJs7Z8RynlxbX4CjqHXpU1B
YhqAIq3LdfGf6QIcvmtOoZ1hBHmWjN7I3SGXX6lhiLAFzmbwZGdaCiIpDzYrIxyB
ATvVZ7TewhfDL3PPW3TX35pOGQYFPXz4qTZRuG4XkBLa4qVchhYCbbHw6ezqbGb+
0DXhYoecO4FjmyTFfxdAy4RDhh5hvbcBqzebj6ZZSYipj86CZ/8FqeD9itlx5BW4
ixGzMWV3XKGfJnFl8Tl5SKINVQ1r/WoUzb3yoFQVvYLyIExmqN4WZuGSKeFqH4Tv
NWDKS3EMTwI1ouF56nlPAYi18zQaZupiZe4Kd2Ld9S6+dsbjmMAwX2LqcYmDyElo
BBagLy+PMN3HnrgbuJ1rcBEKOHTtXkuHV+1zcdTnWxBTt51uNEunXpA7/FCQFMnT
FlzBfaCh65PUMTB0xrx71JzPdI8BGKSAKcNBhkVDLuyCljxl6M5BTzjB2HzHScUm
YIzeclXE5j4qcEBRhDVFrLzM9gnXkhr7lhBUXQhRxJfxAp5l2fXTzlRJunVTusVw
BaZVpLv/0vdJagsMml/eox+2P7qYCFniV6CVoRoHjI/QKWUTySueWYxNNjR32h5W
Rv0eMf4h1Ju4vD1RMUsplPVvCgbEG0eXRQyLys0RGI5e3R3oXje70F+ZeIhyJZV9
YllKAv9N3rXYPfAydt6N0F5k3UvpoaFSz6I8b7q7Z1s4KHJ0ha0QNfmKAzj7bGxN
AvBJ72h9gpMkhXegfq83u7/BwrlIZKGorxEPbhd5anWaFyAT7DeNRWknq6FGkzLA
jpajahhVa0AhejkMFIrSm+IKwKcwo+FEcuDmy/t0NRGDIjGbObhB4vCP1AHIm1mv
FmCMHWLtTWu9O/hMERRKDJ0EI/0KMluDGJI1bphIITwvbsy2gTufzCjGTN7Mf2Pd
clW6TRY7YGZJIzzQrrM1uYvHRu/9UCm1SF2hMzyfiMA4yTnYy0K8xh9I3xLmaB3V
aBd/bD5f6frza7OD1HJwTL2PRH9M7+Pd5JJHSGXP0hkS3R//Lp+9nHQKec8/BWsG
AvczdUTM5RudhKZNAn1ogcG+bOQvQMHtTHr1mPg5x5/tfqfCb34ICXpTCUjJqkTc
ntHnxNXvfqssL9RWbvWbuz3ePPInxALfiKsOihyVU8S+JP68Rn6JtNwBqL/gie8N
JIpJ5FU4NUfau5iNmWo2cfT6LPGELZTr8MGOqhlcFOFOp6ofzGQXDFH7k6BdrT27
KW5NdPDxvwsKbUED51edYhJ1/oC+fD99uu3+4ZRZrnPImYiSzz6wS358JY+fUzGE
dak7Hb8UtTbghXiOPndXsKatR1Tzvpyz8+Mzz5OYK/c=
`pragma protect end_protected
