// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:39:16 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
oqlTr5eg2TKXEhjn1h98a/eWG3U6ijI1RRVtl+yY/ZPKASyCC9T7EFlWCyRtRAj2
np5QJId7/1/pqyRfysumvYc88tnfEgv2S0lSNqjW53iRl9ycz6Ob6OupYZ+bWbv0
NbNhI8iRjOC4DaRhJT97h/SrzhK7IWBX/vjTVToXuxM=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 70112)
fwrN9/Tc6qiMTPb/Ite9UEl8PobSw1PYBgDH55EX0iAdVcFTmSb547EBU7sofXf9
hXMqOQApg5ZNFHr8MRk2+YqiHvehNcMc/4lO6bHuaiNKUGVrvGfsYg6A43OBa4by
HXDuTJEtAiPVbC7YEYxGIhBkI+ZEM3e0hQrsfqjyTUVV0AJvyFTlV08NUwaqueTT
+jTenubG746onm0Nk3crxP67BPnLLPkOfWS997asHsNsRuKH3o9AtUukSr+mg+zH
lMxw+pPlDDYVRDMWYQqJ5Wu5G/Ry373egCgcOoOtWU2s7N5Qhd6uPTqJPZcfMJ0j
A+mD6tvsfIJD2kvD+fvH5looSXGqFaWNm0e5Yhqsmsq5s1zMIWB+ORh5NZrG2A3s
MzyFmbaFQQRFJjJ3NUdqfaKWhc9wtypeXTgpy3L2Am0UjdY60r0DXNqoerKW41UW
AMfWzY1emcn+7Q1HJVBoAec837ndbTcQsQ9gBdjtPbOEnFFm82n5vMN5MymoNFAj
G1n+C34fCaJA6mjSYvKPJMfkOhDW5daCk1Es0+cXBvgYp0yQket20WcLNzzQZ9vQ
sexICtSt2YYp7zkWUwUCv6+fvQ5FMakUVncc97N50tY4hkXNmPOIFM2/gJy6SiE+
qqOEJWfTf7i95LjLqTG/Qaj7pXaQI5GWSMwcIgna8y2S3LXKd/bgbFNmRiUmlOJH
XDYP0FpQT+bttdEYPt1pY+dNHD8oMV5AB+e8tcQXNe0Zgkq8bicSaEjznDEoqlvK
BAWZvu8mQWJ6NS5qVCMr+pVKAh4Gi0PLyk8BcGgC3LZLykXVQ0t5JXgdeyKjQnbJ
zHApfk023oGM7nPKmqSGG/I4QkDcMNjhLJ+lrJwaklajRtyu3o/+E0OZ9Yt6PRFl
tOTDkpRZfi+dnyIyRWs0N252nSSm4UznoTvKIp/H1mtugyQcsPA2Qxa2J/l+z89X
WG9zjnGWD9ZMGMFHqYvWk0ddX6Jlnh7sHCw4LoMpJphfqp67LeCgc9he6kJzPymu
trzDSUa2iUSCeZzS77L+uOnqI1+OyG/5CKT7wrh9pYj5gjEmE7UAc68FriLmxK1L
aqzAQh0N9gznUytA90kuPonKvsoi0gfauBmHDbObelY0NZw7Rl7oH6i5RV/TJ2Wb
w6jjMq9XZBDBBEQliSgVK9Qp3bxUa1m+sag59H5rdbZwPu4UsjOb/yBLpBPwdugu
fy5yjwN7Yhg7IHeXbpeincacasJsyPEcoAWL1tJHHFOaf2eEp2p1y6y8iyOKdLwO
0nzmh4bNcpfJTXuze7fysIvgiXdIxdUuPFmnFn56JWtZpPqu6m+1RptCLB9bK4oz
teGA95WM8xA0heqJ5GfmGkEQCmfV5YsNjNKyxtOFDUKAi5WI2jOPDEUNZjVOYg6h
AjoC2awYjN7b5LL5K+XVDKIs2S5Ek3GdO0r6wmXEAjfWwWeyRPjmthUGTng79gMx
QC3CIiJqPEaLNzWM00emgVRfY4Qv0NANlkpa/QAl/Ikm0awXl0KeL3GOeAAZ8trM
1uSjOHHEntkKdhccFqnDFmNdAMrfKoxKaUGFm1j2CvYfSmicQPy5SgkVLyyxUfNA
oHHbSUsykcepOFRW8TrTeeWTf+C2VB++sQRMAcL9Ff1RY1TmbMA8gXHOtP9+ZIP9
Poc4ARpEvzgGf42Ul31fMdg7SirNDBBwHYLgf8V8aFi7aeJRL6yc6ha+XnWgshv5
mxziREXHnKXAFTsXIKZVw35bIqzSHVM0gS13yIjt7neua9ltnFhqkpUu/6FTBiTY
1V1OaoxNiLdbu03yNjrXVPXNWAMhvUqzklRr0MkbIm+GznNBCIkju55X+YlQkeKt
IIgko6ZkIwMgvArZyiSHypO4nC8r4NgTONGw8rG1ZWid1fwtEV/MSbsvRVb5oI1u
R0KpN3t94bza/RjKuvIIL6zxK902653T+j/N5xuZmqIMPG67gqZ/g+Oes2q8wbzz
aX0UKCYWOiC80zCMMtnHWUZrG6K42sWC+xaii1FsHCdevhR0QLPDCd2IMPNAt50H
QXOo1ng9vBZrSB6MfqQwKpIboVWllqzajaZUoG+CScl32+tLNgBaAWP06uMNCmc/
65kv0b5NUNwVtKdoEbyZF5zHtvA03uo58LLJIKqZMRMiNq7Ch9qd2FNJ4SFH2mWZ
aKKum3iVg4GpRpDjfgTA9uAG0FtJRxnIFzLi7Dw3vbfhcqhIV8xbBFpkklZCZJ9A
aTS9Nd5E7qmZMFEZ7K8LKqj3DNUNTmYEluJIffrZxEjL2K14wHSvGdMIS1RZDr9c
QPVHhzI4xsaNvZ+w4byBsIhXvDc360LCaanktLi2OgOAF8OuHR0bjz/Tn0E/jNSK
IYITbe3u6/jDtz+HU9mJOyEnJS4lrGphgMCNvEqjo/sPkm24ckQeoPysUtuo3WF9
x8astH3kgRca44zeIG57WFCaegbiLAJd5tfvNUmur3jziJ4QDdLiJTfr7ThL8+7v
8C37iU2/8uXf4JbW/SL+L6NzieLxAaEYhZOtNQ+jbAwCaRw4rB0JyWWOPEq0Ic/S
Dwr4Eb75lu49t+eWZhyCQFDsU/G2IR3PMyonGmXyfhJHFTikwDQNp+sfuX/ngUBG
hjIl9cb3MTGQiS01upB8z0Po5tnPIKwcPRCjDz0R4Vwp2k+psIWrhl/kgQyvHu/o
m/i/ahfQyXcjAFYUUPR187Qf2FZyTsHVZQ6tw989jfxAxs62AbK1x75htxc1xDCO
r/EKCOPVpKQ29BUKklToG1J/6K5l4BlM5ID6SjHaqW1r+vEfbg9ydZI4Itf6QAp4
w8X0SU6E2S72pNWJ5taaIWDpqc2BPMEOINcvkOE5H7DeKW02qQqcblDg09/jsDmM
fpAwZZZQKwJLg8zUNpIOUMrJimlEqqAFvt+qqvwRpHOsnH69lsRXVRUeXWf+bI5k
YdcIu7hjgmq7xNpeYSkTp8TwtgihsD+zxA5fBIOxGbZGw6fmXd5JHKdQytrDFDxL
4W95rPERoFctOZYZ0/b7+gVIrrFlKzaoPjKqM1qXlpkqLWoM2j5V47U/YQ2DYHtt
TfQ+lqC4WZcFWt6MAG9epW3hvwF1BI6JzOqlIl/8vzHiwh+vFdCt6K5dsWye87pb
gqzBjhHBZap4l5f2k/x1LOsFNMmbkQ9uZ0uArnpa7tGXV/acW2lrfxESqSomDDg0
xEEl+bZNjK0/vDEXcu3qKt8H9pksth9xlu7FOydI17hqeyU2atMtiL9ZIqbiOg3T
P0YO729OXtIPjfOqUpgO0N50o8/xlUEdUbVoMBbPBggKIUcLq+TVRKZMZ3eWUhdE
BDWfb2za4Op2RW0BB5ptqVEIhHW3BFK726g7TUmnRYyhNmChoWLRNLE15ItsXnnz
yiVOgVKCV4OHniQsFhA6qhhI78sICpUWaHsdkXM6vGS3ojEVHXZCj+5qC0zhi5mQ
IG7gkn0WV53xTF3/sJl8mHlbLKt0KwOykeDOAFtYSn5lvCYsgeI40SSXYKrTddKl
oPSXa2RVRCAvdkX1BKLTuRtGya1pcB6Fnd6ASgxqzyR+YMJQ4rhpGxfK1JL+GG+R
eJLzG79zw9d2knZNPQjMhqdQR1a55igEVheNuo3aeOzP2bAES4V8lskGheNt/huf
LhWHjaAgo8uOD1o3trDNNf5M8yaQ3JS/Lzsc36UfYVnIaVbmYWheIGk6ItpbAjmR
ZW+2K4s5Uio2RBtmmo4MHSn2qetB0uFDIYtwALJtv0XHGjwHX0tUquiubBUa5Cjr
BtgUkJaqBg9zn5eXPulme6xNNlnCwfp13GvasVf2gQVl0UwuVVHO7ruXdJR1IADc
xMsQUsq4IRp3MwtL2au14t5Po5TXWD5gfXh4M2kJs8rBec0TKjtj7j3r6N7qI/RI
hD4/1SQQl6R3S0+kDtviMCxw+pYvOqo0u181Pi/E55Lk8gDZkOUKWq8bDbw3dIeJ
v+CD6lJBiCYhpFoPCZwnr8erc9J2F80WpBD+CCP694tUQHBo15OXjnMzNV1HC/Wx
FRujzpTbWg49q1R5B+l11Hc6eGiDkIURS3XSZ8v0Ej0pMdUodgHQzT5dm/MtyIrd
iMz0FDztV6fgP2ASQoZ7jZJ+4ozKZtznWhvDZuUGwRhgK3AvU7re6YwkDO+nOtwj
0KSr+JJOesq5+UnJ+qSzCc3last5gfxuX/Iz5BCkxDU0dMlzkOPrHnsjPKGUV1PM
ih99goX6mzcFmd0w0jL3UaXfSuI8dXID8718UTO3Jj3RdcpuOq50MD0UQcERdx3t
WulK4FBB+kxxzCFhjHnMmbqOb2S4PiMTx7UG2VhKMo1F9b2Ki3N7V/ruXgmjUAfj
Yn55xqIQhQmEpk8SV6Hmrwi2QW7169LO1VEtYTm5RIuBeo7Xq5GLi4J8n6CMk2No
YSIuxHta+SDpCKxjEdBd7s9OfgNNDFLiKdq+qLVlCdJiFhJ39kIThcqrtJU4ClUa
yo2r2iE70KQQR4gJ1WHlIhVQvMDWbitGCP+9VFkp0SMR5D+YoorcnIILmLig3XEt
rRV+pFPHMDGl6sCPeVogVJhvSjjBl87SIAFpmCOg0jodMK+aEvurOVCpPzkPWkzM
2ZchQ1uEF8F4TeT/zUR50yc8PSKzx+5RuWvPvzqUdGkrJ8qo82LPuIhp0+1TLzPY
p2prLntm1nejyEK060TYro993jU8EVdayMRcLZsgNf/a8mo0RLSKp7I3PXigWtUK
tH1GuzVMapYRILaKbJzD1jXSjjb5uL7aRVMIUZ3cm0Qj6cr3Fv8RQ1qIMoOEKVjm
MOpggv7Q8pKEvB8+98XWKjuHbkVVRia9t5KSq0VFQ/CmjYDdHVcBiJbfiRy44cjG
UrkL/3slJ3klOsG50QiJTN6jy2qJGvoCbRVWC3/7lIaJ5YmM/SUQGrDV8jwE7/bj
+kYL7i250YWMVmiw77Ce6wGt+dmlVn7VLs145m/aDqMmcQcPjwBNXn4MJXA89sIT
Fm5ZYBi9DlgDjfaKMkR1jLuII9jtDKi+GVQVQxwOKOZYnBxIzPzVt8/akSdAcIS+
JjwiYXGqF8SHGPyzFdLD3T1ax57NnjygFaB5aMd0k7AauVY+GGM/3qSyPEu0hqUe
9HpnVtE3giHQmt0c8y6gCcBxkGVMsL/f7YXk1AxxjaihhuFBLtlNfBTm7cwj0rX2
Kn1J/0lt/+bKV4zkicNEi5yDPpkabFwOZ8ohM5MZd1N4gYOKPxzKdOHBxyvB7ebb
uQJn51T9xpM93GEx4PFjG8xYBoTcOqLo3E79UFpM9SX2COnqXs5/2dmcGOSem88l
FIfiYG3RfFA5SoiHPHja61RjO+EsX7x/+xTJK2Q//SS3QDYkpMvAsm4vdi1lWtXx
SV7TUnOshCVV9oK4MPp637EmPo7gULyy5fl9YAnzik8DaGc1BUDzT4JnCPTquFDP
h7hb+7gmHHYmfjBTZgpVXCKaJSHiI4XlOuEtu9CIRLT1sAPOl5a4XgNRY7wd11Kz
SZJms2p2Xws7zMXtBzcrreQxXe+c9GP9AT/y7wjvTvY2WMG75nsu9QlEUcu1ViB1
uhSY3Ezge8onpKRXq2NuAWmrS+z3uXG+YNeURe/LbEKstvQkCEH9Jcb8iFHr7LW1
8wlmowZIt/9mC3uHeoIPq1wTykwD2Y7AzjDylhAF3Any5riR4h6jzxf+C4ixlg9E
U3BWNXfEaXM6sjTsIYBhjp+bmkYkHPjaKhah5dL5l6XkegwrYyVayLTHxM+jojmT
MpxXByYw4JkqmiEGOam0DS3+9T4e7Orv4PmSmQgDrqKMekNNwHloqyPQfcFxRXtv
yDcJXlFQDFKWhKcKrmf/VHlLHeKAunQrpmNAdoqlkM2TDi3xCia53AzMTGvJrlU7
cAZNQ4BqNb3mV3O5GfaHw6GZKpjHqRYGD5aDB2J20iTtkQwBXVYoWRgwNEhFECHV
v1dFenO+FceQDvdJJiijyw1chf3V2uHBlL6XohqcikinGdFIsCstVZP2ja3v6fZW
bbinO8wIrrChrSjwy/qfmMm+J57dQb+S2N8wB0Rl5mlwS5G6hRgonrEctGqZ+QnB
A9cQAAfFbRMb6KD9ejXQ9fMMWwF3c7AU0EON9MLToLsiP3HQqQSGIDkaSHHSeeTA
LbFLVEnjztuI3mOxVuRGNbMiqU/urdO5/ZQfY5vhtz/PTBrZHJrUSIavrEC4Zz7A
s6JDGQ3Ylw7Y2RJJjf1AnKdnk/qEB2qSDqX+TvBLAg8xkWTPgRLEHIo1SZji1sds
6D1uA/BDuRV0EfTjqVPu9njG0dyw/MNKMZu0rNhTj0emLIht2bAnMWc35c1zqkaS
s8dMYfCawroAnaca7Px+chihbZsYTWE9zWP72TboWJINkr/Or5seVCHHd2fGAcO0
COdpx7CCBrCMoeuuVWjWKzXtoWcSLdAdaR0s+JXg0vgBBe0+P/QgiXkVnFEWnma/
aOW0gKX4d2zsH44YOyOq2ZFLNdmRwmV5hAo5gsTJnYUmVs5Yzl5w3niFIK+2OOQ5
zd+K8235RNJKQY0FVtArTASL7twSx0trNIaj+gFrJHsf5ZjevgaIaPgh4H2KIOma
9uSUSUVH8dnxsck3OM8bu1dKe3RipB/0bWqwyOgEsGBRebP0sQgcz17EghOGDyLc
JcviOsO6Hbd2prh+oa4bqQpJnV8HqVwpf1LT46GxZjLgjlAJ4YQ92Edkmag9h5Pq
Tm/NqFTpRX8ZdeSxdqji6Pf/uNFgx/nmF1c6m/wTTSd273ogPcCxuTa60ulnwJV6
sccAr4Q8fEeT05fWrKzmDfFPlKKTIkRQUJAjew02qgY9gobS9EIceg7Lb31SJup4
5gh/0iV8VIBndT/dSMHHPJSZv1efCE3FUhVaiRT58KlfQmnG2boxwrZHthR+NUII
MpuS9ATjl5sp30CMMcI0vtE161gRGB8aqT1r2Ss5yW6D4AiV5gCbVKxjzllG5Oe6
7q6ZaVzInCcVqv5phToqoBBYjWS98AIPCZsPqlDkC3Evg5+95LUPzc70wgTzOkGu
YVc1pFfZINIgr7ectmKHsFeGCR//19Sjfaqc+ULw7gbvm0SAJ5JzZnB/Igf1t82w
u/U8VXhBiFNSrmlU6lLgjZQkGdEvbKEzLxS0lw59KMJUorA8XInoajX/ZhfezWTf
o7stFPUTYogctP3zGcXL9Ckw/S2q3PV7kXRCrwrhsBZjx5qqbvDbRkuAYMMuTbK6
0gaCz1VOgkifl6OW8k0TD9VaCJ78sNTJpGJGBNRlJiSr3JEhMERbYDElfaj3Y6jk
D91wARplrzjTrb2zcU1fA8z9L0GGhWl0gMtqzT69lTCJbA6DuF7g5sO5jHekqo/C
qrTxZMMalhwfCnHMnhsECR6DLJNatp9A5UgIlad+NmmMLijLa+oFrHjdQz/b1fvS
+sfubClA5RACY1DgwVsereJzKwG+fhYiLbSUKXYi8KqCfif9DpdDnRk3unghx++r
WaNoSMQM65mmiu9YQXPCHBHRHU24gn8XzIK39XXhzgx4YiTvAsqulz7xXBccFYxd
eM/Yb2YIdoyHOoXihP7cq0GJKjS5qS2gxRi1vnsFibfq+6WUyBNTZRTcMEqCSETZ
H59HwrVZuYqst0DFiKI9/ih0ji6E1EMas1F1hRrkHJzXcMOL4kkVSCxl0yvaoYiB
m0eb2Hr8F0CnkbUePWZA5mJgdOZVdHIoYVeVUTje4BjiutFw2LulwmL0sBaOyVqW
9vlb3WZirE8YW1gcEC1omYUKloFJZBx7Qty1y+lysqjlBUSEK6n3Rr6JYfgJ1v7U
ycqbgX5+22L11WmmtBwdo8pTHzYIT7TCYRaYx/Cx6zu6uf/8ImUBH2Fs5+8ExV73
uC1UUzgZvbrvfQzwO7v2lA1iYNUohQ1HK1QiZU94dxGQX9IhRh6XqXbQLnKYiWYr
vsD/s9d6wxccsliYLNQUGcSW9DeeuuVXOvKMidvy13oMHPR3UsghyE3nnNXHt247
QboMa9cID9mAZrYSkTBGKsoWaNleT8mOmJH4DfCAMFetuI8K7YS1Sp2CRRncbP51
XWHNc5SxFRfaHr9hGNIceOYvErGGjaaIvZ8Eom4oPJvg7az/RIGlt8giv9RtGWu0
lRmB7OXKYQxVI0HBCq3oiFR2BAGGZmnYipGv2stFaLlzmM1Rx4CVidAkCb1KngJb
2kEldWmy9ODouPoEREyfRek3dUmGfKei+6pxbE0dIjq3FNH6mk9KuxAFXWw/o8I9
V1f6KqSR+psOje3l0l00LtZAVhbmWzuIB7LiyAW4kY4VTejaRXWsPTv1ro7RhqL2
rASV1PJwqPELGLsZ4BvNAwZyiObZ2sE5uA73buhYvKBXChEwvNeNK597GRhZX0Nh
9Vh8ZhZlKcxwCEbCmuqsS7hwmBq0FNOZaMG6x0XyldYpQk1n/olwCAbAC2Tym4Fl
Bj33pPX0UZUcUyQBfB7wAAtXock3VEuQlroiTtnbgLgyNSRTYDIp/QSN/MMwUYK8
QRxeGhFjpZ0QyyZorm2CzjfrQu+gFMeguM/WOosuufThyqpDG28s2kVFu6YE4+4M
O+++0UX5M2I3MxHWB7rfffPqt2A2ogY0urwz5aFnHBZsNUKnJ6nViqMGD4wZegvq
/NwWDaiPjhQqISyH34LhOgEwjUdX+P2smZagHScCVwoIzenQyBRY68pb0JAliTgY
fpphQi8HuPtdyMx518qjs6qI8h+iVPOTBR8mmhVJiGY1GSIMs+o8jjxoFEJ6YpbF
DPXA1BIXFx2g+xnJnFOZ510M8z0EywLk64/o+Q6Aeu5/CxOG8J4FKHuksI94wAl5
5DiAzk1VlU7mxGIei2PqcCZsGzsLxzh+V7TCqSan1+rb9RO0a74Vd4xm3U4S3jVj
0cOvFrL3h/y0L7DwabmLCgNPLZh9E9wv+SoDaj03JZV/o2f3Jcxq+16T+eJfVe3Q
tbjiBYPj19WrExAns9maT6znCvhsXoXH4XL0oRdFgBzWehhWuSAH0ir06DpyhCFI
lXi7gvTE5SZtA5ahLTALD5wRPxrkGCLf3jVmTuk/3UulAoh6WL/eGGA3HBbe77c7
Mi2/PNuVwo9lJ3ASCMoh5ghvVM2pq2J9v6S1y13Bf62wCzxAkiuK9phH8ErSzoV8
2A7ex6xTEBGsLSIwn5uIfYAVhgTN9XX7xh55nRkPJfycfujD1kNVQae3YCNfHPj7
tBbLIDuDdt8iEbj9bTY0w23xCCUNJ9FreZn2hpOGDLLLHt40KOp757T2//o8wBPX
RQEf2ELZnwSOZoG+L5lVaPU9UySrwa17BrWYw8qUJjoNOTcPVKUlSM7Ri5Z0eI6E
+6hQpitt5tV11e3MXL5M5xjAuokxqJV1NLo16izMhwpGhSvW05UgiD8WE2IrUCki
3FrYvdPXYFrdz+kHnzqQfKryDwn7cz2L5b23++s2TWy/FjTrnph5TaZ70nB/e7iD
irLLYTyjlTyRzXFa/fx3g2Latem/BqZGuo1DjwIc7xbt2LMvIEbjRDC+5KeZG5Il
18kuDahCldqZbsWJSGW9GeqRe6YwcuKqHCjYq8jG1bzssJHCc2z2uHu04W3wLvOH
PFi9RGhlx6aNAecd0tzyDI0xWLjQixVtcLIWuH/DfEcv9WEnntrVmbDeST2lCuqN
4AutwzfaaZEVMoEY3fLVu/27UWCR2og88dnIDxYCkBOVDRGzlRqrEnTzMrxkDozI
bqQJdrWtuCbVbrzfrORx8tGLLtq76Snd7KedJtWgRT5g+mizqgAlcDcZytepZRkJ
pFbxougAwQfoMilfeTsZlEQZVVarEYsC4EF1djNkDB0P7t9lV5ZceWUJmkirWkkU
OTbKdfJtJUUCNU5FexSVrUi1wPiEitSxytblioaH8JTSr/CqXn8JA+BOMRdtUwqd
5wJco6Ja5mZndG/VsmWudw4WGNdjbXmxqTIFLn2U/V9+OPdwf51WpOCjI2ahvq02
4W/KaB1Z+4hILv6Dy+MCrgfwfG/WsV7Zc1Jaix/uLpjY5LrR9y9gFoiPF9VyYiu7
Kl5AKCVEAeqzhCB2vCKTLyuSYOR2dnFoxGdTIGqhLuYyU40ZdkncYrLJoJHzMQDN
jWyjC/n+jKA/mtNOX2d07jleoDyF5twt+la1XtV3log/5qKbuGjmI7e5m/b9Ct0Y
g5kak7BNO5VApq66GOd0G3QDpBNWWN0N/DWdcICyBjEU4Fa/aujyrwCybnbQ8gI4
yqtjLpI9y+2uq/SwPVYF42BCwUgycOd6zNC+bndMBc576J+bLPZdaLC0H2ifY2Ny
ZQIgP1j3u/yEOU+YjIBX1kaol4hJYXqaB4l802HcdjzTDlO/t3SB18iOcsdvSrAJ
bRc04LoQ5YZbEz9PxCvrmzUkpZ6m7swyrgZajl+y/svC7LYE5ZitqVnndGsJ+DRU
Fc/d3hGR/ZTZwXgSW2sNeRexfDRomG29SPM9U2k761/tiOTP/mtOn+sa66wu46qN
aC88Lh0p086/6oI0YghaUCdk/ChGh3pdKOpIAg7gt9ST2f+0hxUR2tC6BgZqNyWk
P0OGEAWxK+VopGQe49/0vup04j6HInxW8L69tEsaNCljWgKUyVDlMNoO7+2WQIHu
BTXiBualFlfHZkmP9cz8Dn5VSTlUb/GE9+dYLMMVny8l7CuusQMdp2S2yEeQPexm
ZR1BKgW0TiWCyzeI5NRwSLy3k0KFz0Lcff/oabkbI1/TTlljXlQkoGSf8uF4lCyx
joc6hrsHKgMPzZoDdSnHafB3lEjjv32fomy2ZT2Nd69NmLYIPX7Ckv35mGlxis/d
CXrTZCKbeo8nUeGaNcf5aFg++H8GuI4o4aivEKq6xZLrZLWQ3DMx/Ro09DJ1Szod
N2NyxJKwKwpXzDHQ2ZrR14jl5MlDiJuQ0BbWsfX9l575pkmhtvItkqpCPTABT55x
c+M1zXLQkKcTAZEM0rbtJmjBYQyGplZOk49UlFTPepdU82lBmpYyOEzQCKjDNC01
p/UXBLfAxjCjl+kQVSBwiHfMZJ+TzEEkyTzkI9Lqa+Kk3WZnmZn1+i1ErAaLN8HN
e1HKWshanlNycmkYCDS/czMDaxy9vEPtdGkkDwweCq2mB5/UUsol2pwNnkd9Qvr4
WP2TqvE1T22ssxYxcmIXXtMA5pz9bFvu2lYDGQdSxN4x59p0YK1IaGYERz39aWUC
Wx8CVNIlrZDllTg3zWPoVFnl31j4cu4T+Xsec4+p2y6odV6oy8y5kOXEeRrcTAqZ
Qkd7aboAG6QjiHyfFaE8chEIG5LjA/DsRBHLQt1d8p9fYg0U9cgGoJMQ++M2nqs6
GYQe7TgIuLaAZwTnsqAMLHC9qioZfHVgX6ZAfMAios6GBBEgNns4Wqx4R4GX0B0v
KIzz/dztEgBHgOKnXv25wQzBUaqPHoQlp4EJF4ZCAQZDZ8oDn+7D70LG+DXOO8G4
u85UKWU7mY9f7UFhcA7k6+NnmH4LZCshJcb5CLT2gblH9ZFr63Ye9ucJ1WDCy1pd
xb3yKq015yFqCNVy+IRKgFCmHiNPDygzdoMURGV0+lE/+Wj7byQHpxwZQedCd2xg
l/OfOc2kHuFa9EYXIPbq3vVSfXt3TaCCVVVU/kYRsMc1rkfpjhUJGPPfO+fJ45sq
3tXd3rz5xXpPT9uocC+ek1Tr5moX6sdDta8nJvBdOrgkb0q1N0Bh/3keeBYZioiN
2n+QBMcfRqgq8k156Vwj4xcGy/+TyN2ZPxUKKwJkte8bPR+LYHc6q3zwtP+Sglt0
vbYw528DlzQzXr8vLiifIpqEaj9iQEd8qJCzG6nfKmWnvy55u8h6EywHEQ9ZtmcS
6TPd54CoeeOzZUH4FrXVmqPhX1bNdpPuFyA0+O1JccHzObKIq9K1o0/nVihY6fa/
lIlmlJJscCZggiUs+lKEYjWm3t4lhoQG3IiHTQmoiluwn5F8SMSQIoW/8wo+knnX
LIc449I+Kla1NJsqAqV1JQGllxsMtvnYgxxB3nmmRjHYPLWWnfUSsKJdRPiyD0jz
k5qRhxdV+szIwd36vR5w+m2A4rzPnqmOmA4xzOq24auOTMPjgwz4I/oIAdIRecXA
33ngYVGLQBbLMMmgcAHffC0G4yZCh4GtYBgfU5FHLMRIihD+Oodn5U7wqGaONS4D
Msgr9wAt29RpT4CFuSHb81LlnvbfpghtRqzbIgoIHdMSGDcS8BR8XTYQhhIDayqT
l7NqrslwYxtOBtqwn4hSeZIj9AcBDY5sPE21ruUQ4yuvlkHV4ob+Xjd2xyCGikKx
vU3mumKK4h1TB3TLMiCoKXk0aV4kNbPhBoNARWW/F+csO0slERiq+nbT92tbmwlf
Tvr7L1h/sz95QRG69GnGvnfD6AMZGwfVyEp0e3qDXSI6EWiiXZgbBmI/rI/o7Jpw
Fbvyhuz4ozOyYk0XkH23TLEivJiyxeHHrn910zPqBcHjdwHIaZyDX4mhyJp0Hg/S
Ija2E2YtWiSfzpJNSWbAajNPcUhyjDNJ8DuhX7dxCuhSkJjBDMlkMJPMT93Ynxlm
L/lU8JGOKackd+9hCBcpEL2saaXO/Ul6p6R7QbXcc+lbm9fDrgVgbWObzBcHLtk/
Oke0HwBqblWNQ6bzST9NNRgFDFHfQPtw/BbN39H3newwOc0LBL7Ex/02KU9qVRU1
af/rzPjgHsB4QEhTrJcTa06m0/1viT10yEGKLd+5WXMtC/qIBC+c5QkissXx7y9X
lzXc+mXjTUS3vU8GlsUPm4MyhYuxw5uXSBYGWIqIqWgTQWyUZr6EFZYUAe0SZ3Fu
fCYzUwI4uyIub3TtFFPS1ni3ALBj6eK0/LmTlMyQqQXdfnNdOZrTlKtWdW1t3DTH
IBDvSSRCwFmRRmqsMoqAeW1l4Ln5w/uSSmfbbZhqpjfAqH+tEdUkAvEgWik4dxt1
g5oCnxJUQFGbuJ1KaytQ2dmE//3hsnGUhbqlUs/B1mVmi1vE4JhSRaj3WrE7yTL+
95za4zXXiM0ogweSTjKwZ5BBNc21E5xojdtbD1oAcdcbz2FlAdxyoqtHO5c/U2cI
SeiZofirUddnto/8pxGLRIeUGJ5KdzTEpb/r1Omf2QueuARb/Up5kpMDAXeti+Mw
XxUsn0R4DUuV/K4Xh2/TTWF9k1ZGmeMtOkVbMbCwRmn/bOb3qSwUC+xUSwiNWEWo
8UdahYrxwRurcf8qZyC/2f2V7AIhKySDKLGi/5O4iofmAJ5NhiDN7+SgnzfhHqlO
RHX5P4H8O8y1a2ZxZhOt3hk5tFt+bk3lSpsKY/tWU5lzxXQ1G04aDPBFb7qUvqPu
fQB5dL1nbIbphB/zbSDzKtmAXLhhzPX2d8WusgbclPORHYEl35wvttTqOY+9iQHz
iL7vXI695SLK/xOqhYXyKEKYph1Xk970cxayvuRoWXq9QIXdX6jtQag+MqCaFJFY
kvoWEQ2XNWWX4U3m0o8DGtX9TRO8tBwLOxp70Ah/zOaqcAUNQLMvCdxL5IIYv3o1
bu5OOuaabvE0w6v8lBk9yQMx8ymK/DlnLpUIKD5yKCz21M7YOUjQEu3L/iihATAd
S2Ie0EtgnI99ra2T8212YOYZKamHSYEpBXe5SDfH2N4o0+0BZmQXprVNiKSWgrz/
PTQIwoBovBp1V+xScK7AVMBRDOnWqW+MqkYjBLePCB7+/Nql4UqnaRjxwfl8kEu7
uTKo2v4NPFaBu1CNxfOpHHt6MvBogJDNYdTgMu6mDFfp/wCY3vvq46F3uc8RR3G7
71w2piwta1QDVGokfW8sFU3tekpMo/7whupSEryDcP0HsfzSjMMcWg6vK7Z6cCYg
dfnDW2bH4F8Q2tttvp5CwLzR2U7mMPTTtieP9TOWyKg7A23YjzvxKBiIb2IDsq5A
wR6zghmKeTP/I7BEvtopK0bVVTGnkkEVWEeM31iWnT0CUxDNvDQXyCLGZxWevJ4K
T2Vwo7cMflfbAHExGpVNscp1/dwYR7vVVb2TTMv765rcw763mlREE+Kx9A+E47FX
+p3ja75nuBAseGAoim+KZ7uW6CuzK6qG/wEKLtVsPVuLc6TJZ5X71No4LncBPnQy
nLLlFUmRW2ObuXwiffuCWm3eDYEoKFHPbCC5yz0nF3qL4WaWF/TrOKKs/x/ZoDHy
b4mynvSDCp+3NK49pePX3p/e97Zd2KwjVOKQfCuD2E/2cYllO1TDHgACT5tKr7H5
BY4YliMNgGLiwy7kHA1odek2YCgHOOF/xQS3yizsmt3jpWSnhAOaxlARxngFT4ZT
Q/tFVrH5nPfmvuP510w9vQNl08BYuTWWTkCa5AphG5tPpq0KlqfXZgul5+gioHwo
/S2D+3WGMlxrtKdWZkJw68iGQ6smpyNqgtNYkUvMKMRv2sN0dkzT7cRYG4wmA73l
yCUdqNoRyvdpUc5CjHlR8izGIDhNY1jCfBFHjStTXl4xpm0QNPjBRhXcs+c2Ibg4
pGLv5v/gkmTuGFLXzCGXIKvzX1y/U3FDHmeSo8AUY11uzGsYXn8qvVc8eLkjtsyL
FlzYJVjRbItaly0x63SxPCDbOfHgxauveWKabXHsX/LA4HKStfuhpeHadFVhpVvm
idWW3lC7fiqSMTLDxbhbq8Q6kPSX6eoJh6PQafHi/gG5Fkcryqpzsg2pPuJmZapd
MLByTIg7z+zAnkeNRnBhheh118AMz+pHI/2I9E8qsrBrtdZKHqAD3HsWi3Fjtt2p
gS3oCHTS0BpDx6WYDhPAyTnT9HGPHbspmy1DCIZSpCQQuliZEPUmaPKw+2iSgYdg
soeBF/S9JSBcvcc1VfEWyVK9oUJkPG91XYAV29eUZsw+7KfpalWVyegk2TmUFrrh
d2y6Jo6QK+qWlZXiIo8RcZjRsSnZ248F7AZHLaYchYMG+LfEIPCjRg+JT2GC1RyC
n1XgHM/lDgcQ3Xa5TGRR9g1tvo9EkCcbINlrAGhFn4VTs5Tmqq9E0R7aHLbxmUg5
Ft69a9c+ZOHMf3sgcEB9XCAZJrZ7+Nkh8PttQzvBMtBnz3DB8wIYJ2UOuARQsHHO
gm1YfrJUhNaSDsuZgzitmiX6Jj9ocfOET/MqQjw9cOildC4ZUmNcLWJCMGbcwik/
gY314tNXcnQwwI6l5u1BJakdNyEttZu8Lmm3uJsJEmvr3slitFR3WugNBuS4oapz
2w6jiw3fRLjng7uBI8+1CO+Yucwhg1LMK2f+cNuKhspxrM67uUoBUKTs+Jer9/O1
7H3Edcjd7rOGu9PG9Cp4IGfqw9jlQPHftmD/akmyquUYUmu6KVTlzVMXcW65bI4c
0jMfyWsxbQc8iBigsK1jwR2Ls4gWh/GI5LVqdOQVVcSLT1k4O+P7kyqgFgDt/+ab
WFg8HiGFT3h46hzyggRHLpkWh5M2UyW1KQtGceAyAgwSYdqAMhnuRSCsI6OeHsgx
G9nUiZHHLFPajJgJhb6sDBwikMBaVmj4s6KbuKYW4hnTAJb0vhgVIVBOsCLxu47h
mnqw6L1dFpyUeNCaPXTZTzO3fe1gDTss1fl7MtYWDQcd1JoQZKFY/iWo4DVfoN82
9GAtY3vD1VWBuo82GInKmBhxbPqTzM4pUqQw8KN029vZOXL29L7VbPJUKayW1ueN
7x7jr5OjA4yWSPPVQniKEuIlNGGcYxugn3F7xN7divt2pLTYQC7gYL+8p48CdBIL
iTrZWPS1OdRThQLzmHsYgVn3Kd9mPA6t481Y1zeeKuK6xfmlDEr1uvXB0o18zM4Z
7Q1ZMSAsq54s6q8ffijYMXZVt7vIidP2VkKrVF9QomUq8wnKDF97Fzk6QyPeuT+Y
evGAeg6abDAVcV+eVa0nfNRYFYlLlaC/TV41cZ4XKk82Evb3WCsyf5fj5QIgPvUi
UpkMFeMiTNOrKugX2XbU2+l/Rvn9BEvJrXzJmzSmwWtFpIeGGYncq0V7ybabICjv
rjpgWM8Wd0R0yEUUWvdHO3jmlbwGXI2Qun6mOtsCMCA38IGpkUk4AxWo/U6O/3Mi
xx926jA5r/HfnFG31O7Da5Xi/KUV7nU6pRANAnHkyu4HUePjCGkWUdizqmg6cbx0
dQNCI40UDNA7JNvdUGg/rR5otRLNHPvH15l7Xgvwy0kkV51msPUj54h++1+AyyHg
n2kwQElnJyBJuUbB3G/Tt9lI9jrd+OZGmlDgcgNsVUkyk8L2i4/7nelgE0GhGTcz
Na3GZRd6I4Ey02TJqS7srrdipOju2BF9vPZrGrPt5lxkBcYKAd2ffJQkduWl8IOo
EE5HqwvQgX/tlRkYs8TSQdDSO9lrSxPqygSnWz6U1GJg0gTl0Gx2g2+V9G2iSm9c
1hPH84kfJR5H6X54X6dj1u7Fwk5dLI9NGMtDi8s6eCmCbYG72Ty/AJibzV18FLeU
ld28zOuU9rmORGOQGFa9SjPGvHzgYRv5yuZwDfBTQ4hBE/RA611ssyAj41hd9CM9
Uifj5kC1DGOJ4vA2wxnrmF9qIzTsIy+1ImpNjLmhlagFNLAp01fXNgpYSBaVli4G
Mz5fiJ81QwGLeSRGpQo+inlJr9wYWinXjikx5qjdpl9mI94z/hUihxtsCIptIxG6
iKJZvb5FdPTQUWVRmpZGQ3VBbaCveaUheEfVNB4QMIx60jdebnSMlep9MRdpTEXG
jRxNo/QkBQAwSfEgY6v/YruQ2x61d7RQybX2DxTGBI/1Mwc6zutskAn21jdUIcwr
HXHkRaWHpID+0x8PMSUtPpI0x415IpgTbd9xKb0gXU673paiTbn6awD9KNEMa4Aw
eG+ceR5AsvipFDcm7MJDeHYozVSpRKcCjQGtRafuX4R9Be2uJEQFFKCGaIhijC3f
GEt3BK1JL/J6ZLgdBjf0+2CLY59go9+Zfu2XPL+aODiP11i4BlHZIfJAzr/+NFjA
7TuHXY1aMGaFjFng9J0Wjqfq29dW61xHySKZYaHO3txQN/ZLhjrIaCyJNrUV/iLE
GcUw53MEKjnErQdhH1YK29Z5qQ2aUKl3cpbhCgAqIEMAXD0D9ULmdDsadcpkTcE8
UII47Ky0SzvddTYbm/MgzOHA0bLiQxXy40/7r/hsDbiYxKlwxTABxISy2s0HnobC
cCl3+jQ9Cfw8qhySKDycVBjMKWyUoUbfxLsgHB8iXoJEI9J8oVfm7hOG5KybtZ0I
pDqPm/Wuvhvy6Wz1Ud49iyHQ5omBDm7EruqxSfSe1kZ2V13JGrTgE8b0b6wLG2JJ
QotlFXp4o80TVtYu9gXsZaPbQEzofwoO2vr5XJYPma9QwT9B26haIOUrZ2hZr80q
tfbcFT+QZqs/8mnWgPbQCpIKnqRjBoQGqR/IdU5wXgVnPRMlcXIi0OvXvVylIZQx
Id1gXCgy/LKQDCFJpBbRxBktMpYrnzGnRIcZAhwIIy6cRwpOeIhVdFEWRtR92+MV
NX7kFTRNUI/LIUSU2+ga/++VakE2a4qScE7AdB5DDMzroYnIEi9U9NlqC//r5lUr
7BXKohk5j9j+/3T2BZXsVY7cdqnXufzKB1Wi+rqhEYpimOIp9fotMRvvb5IxDbK0
q5U3zKHM9OoazrwBTi7yGpZqBldI7BVlFTLsWiq7s4NWY+V/PKC+jiyHhQu+YNxG
153Prd7U7vlp5qapCYqmVer+0JVV4j1ovdPkz6hgT1qlELZlGhMzR8y4ipCDO5x1
ux71e0S16KredrGhIadmDSSsmtTkYNoYpeIcZMeiuZL/e08EW7tLo4Ujq1JkMMrQ
RywC+LHCxdvSpnD3Pxkb+L+Cc9Hpmzr0bzur1khodZ3Ol0ETchthgGVJzL/SHdsu
CimKxcEgjZm9LIiw8plrlY0gWyG5a0eUKblK29hJmw7pJQwq75ujKOAybPTrYOXZ
VSFR34FWNqJ+CINu+FooUhtKxcDOhqyh9gY5WRoLYci50AcR7Rne5K8kUx+SMxqw
GXLkpdR6ML90aXmhMrNOCktD8UfXt9WHOborBOJO5yeScFwtGtgpPYPWR/1HkgHR
SeDNTaEx48OIhcH0RPHLp89sIA2inRuC31/5MyrOaIYsrWvcLktBvQVHPCsj5V/q
PTNXF7EG/CVciPdYa5PXsVLJLEQMdJDqBg5TnCbQs586SMT8vYJNDwtdC7aa9cdf
VZ/SwWyYWhF6gaZEckipzxDGd4M8T9tPGhCILqlEVgFuanvD4O7eL9iLaaWm/9+O
jjfSWzhufqu7u6ZESvYqXOkgRxNJBZbv2MxL2GM/F/9wvC5xmRDyW5HgTZ1eKHMZ
obJD7vkgXeCyZl6fZPktuChQcrlLjbO7UAnmfUf7T2c7UMVlGqoI0CSdfy5KsYpm
BkH7/GOJYoVSP4Ffb1a5a6GhmD5dK1IHf81zkudQhKY5ilq+XufBfQfMEBmnrYby
MtO11qm3WBIGTcyj8K/jzMDKLbNFxrBrd2Lvv94KnHPbvjqnN2N9ZP8CfGDyKxZq
oJ44EZQY6uNuKd5keVHdmhaHmxpWIFB2kHDqRa9V+KV0BqVTCO+Bdj3mt5RGokuB
OaHaW7Kzz7TaJbm3OGEeXUMjFihEF3yfJz8lory/MBc8UTaCPKPkn3H917ThZL1Q
F1ouNDNkzem/0A3373xOTmmIvX4n1c1+fz0Az56zvm+sMkfMPVa6Q5lbapD7ptfU
aT/FsQjbhLs7Y7kemUQa5cg8pel0KAiQno5FP45LWPRPyxDDZC9ipxPTVRyEsIvj
o4AvAnnbOVQgWumdshrItneyKaAFC38T2WoF42+Z4k0WDSc9tCEmL0ycBR8nLw1f
Ptc594RRvR5cjL/TeeGrkKVpBsHYiv3Pj1YuypYUTICFmceMdeZYycdnpPM3/51R
u6OPLS7PlR3x8SQFU8iNPCSlRzQfNonXb+qyN+cdQGeeuCU4g2qzIDVX9JFx7c/V
xJMn1hVQg55XeUb1oQo5feSZtMZI5WqAzo6wxPwBEc+ma7IsThKGNRqMfJOpSU/y
7kRGHQdzQdEhXyHA3jUZzlC0EZGVFkQt/hv2gzOYZlcJZWmRimdtGA71JAyAfA2y
t0Qs47p8J1AezYXxU3CCJqtoIalvFJlDZxArD4aZw96780LY0y02Y+iRXpar0EzA
WUZEJcljeJMRx2YhnC61jw8I2vxkfZ/B462iGiAzDpBA3JeWB53esGf/nOPHe6PA
1GjJV3OlWE/gwQ8XiMIBaOSQzF8wBKN0+VC3aRcuPuQDNVXtGfAr7QX+rVmwpMFe
7CyYze8BGh0gDuKAdlcoaoekvQ3zwV8Vrp8K42d1JWYDi4LFOih2vx2Kq4h66d2R
dl/Hr8cm+bWBFXgrG/17jTak6yTbus3wpXFp1RTdf9GUW3+tK4DD+2o/mWvyhpLO
xvOECEm8jbuVBpRB6MN8sHJcqsLcoEdUCfZYutIfZuKIiMSWP24zHT7nBRwO8MK3
j3deGuofkjCYd0uCw0l8NAnSUVQ+y2qyTLphyyssubY1ePbmvC9pWKAd/UFkU/Sd
clbssBhHulRBVK0JCCKIrata3f23tFwuCC724PJY5dJHMHSHIt9GUM+GLlAw7Stb
oZ+16Vr9HyMQsdLtn5WeurCM0aASZ0aJ3LswgxZbVhWmok3xvibPle9vNTcsg6MG
mQUFxDdtH+FS6m28c6L0Q+A45rUZu0eZ/jAeWzsACH0tphhjP23IbcrG26/VETHX
BvgjnLDjnqAdyAEv57L2KlPZq1AhMlPN1cYopVXWzRYAV3yob/bXxLFP0MJtFdpk
7oIKJkM0/zTBP4Slorunt08sIRMX2p0jZ+1YRjewdFU7L2Dt+K/v55yoJKcDvWRy
FDt3bKpQUPDJTvueAaR1pBl3OHRT4uB4wReRYy9ms3EHN7VZvKmW+N1R9cgPPCla
4bYkRqd0ykf8B16yjp6qP5N4pcCZ6MX63T6Mnkd2nRjOgbOZhnpz8gfhwS7l+e0V
sy//hiNFWY9HZ0BRKFOFBxdMUb3cbDzv2iUx2Rb/VfQYrQm7NFQxqycSnIEKIb/H
OG1GF0N0ydJp6IjRXJCMIPgAKtWCsh3SM7eyCH5D3jFuucVmsoKYt1g8Fu21QEM+
3IC+JiI6VlGFK3mYQ3Zg0YxunYwBoaxvfGT5pDMdz+qPtDV0Ka4Nzlg0X4NBIJNW
cVXk29c2ElWu19/RTquNhKNAnmJ06kLk3/VwS1/oGI4yAJjLMY9urQw4GoE+IEV4
MP9N2lGf4HMSkrCEyLyN+vZU/DYbkKXSFLnM53qyrfyhSa/RrYEJydV56CpdWsKR
gH6u9qoldSqvo1NGxZlSFknXYle/znG9zMqF9yuBKFFBBK5WrE6ielYTDK8BlA3r
9x1tY5eq9P681LcdKBZcHw2LaakKBcluOMUnoQxDSSQb162AJQ5pnQHhp8xne00n
jErkKIMRHn4V97jfvaMLjmmKd8w46NgEs/zC4/gd24cF5o7C0rtqV9EJfvLtUBqp
B2L7PFf8+6zx/dk1Id5PLWDDsMOOL1aDpyuw13f7D+yRzv6kCE+VxoKNB8HbUaha
oGvd/L7j8CW3uurScn28T2qNP6/gh3ZZBc4ZkwAJjbYFIScayd8nVnM7Z1KLj667
tVXY8C2Q87vFtKBIsEUa9qrw60/vguq3atbCMy6fkgo1vPmwJHiISJ+2+SrGc4SD
m/tJAfaRazfnsYQAkv87xu3d9oIqj6p5m5hzUKrpxp7B+t6vycu1HEA27TJ8hbmz
fHXLzxB1TXoa7+p76KI2AsSwAph/gS5hlx4ZBQRLKCXUFL+8+4W3inL4ErfTgk9l
Qsb7IVIeUNW+9AUxvLo3kZJB9kTrLhLnXDGkEsHPwzZninm7+1pqbnPTkvnPD9Ak
AGrI2GecV2a0ESbAABtfF/CFgUeqU0jS+Aae7ALuAw+KB/KFxzD6+8Vbt+m2Xu7k
6Mhm+ug4yGTMkVfelKzXgkFocYT869w9UaSwJJvMxsTofOK5r9eyoK1XamYyyoTf
I9kf52CkVlOz6xagUziOYjAUHFgx/FThmE1FxzJV/U+++8Gz/K/VdRmrZ/IUMt/y
cOUCyxZOkRk8RkjD5271RpBEcgAWpMMCE7cmIhI16gDiPG6WSWoq1xml3N2XGE1n
woRUo7xe+4XGUvU7AwX94ZUur7IAOZytGOjIeabCRTud0qdn3PXIOHpQOKW2crk4
LUMVy1tpy8v4+x/r1RnW6L69K2pIp/GKBCau4IgYUc8ZQV0kSEh4VvUdayHTT2SQ
poyIm462pHEzFaqU58d7bgKFgSQAi+CoxjmuSfu1zoBLyukMKOpWbXBUwvuXm00v
KxZGvRnvSfJayUmT1DPUergbjMKp7qQb0SdpRGdloeTAkAgbOEULPFB94TNORSV9
KxPAh0x1q/FaBjk+6LrXMJ0/qjIBOE4Yjulxix5P1bZ+EZObxRBcLBf5iGuxNUAV
UY3z4+XSCqsl+WO87wNfYDMOBjYgShF5ldGkIe48xhHO2bOW0Iqt9FuUX9otgefL
PNYCSAWjMZ4JBdakuMZkDQir0ufRKdM8QGokb3vHdLG8t2kL/IfpS96Y5bdMt6PV
3teKc30GoDBnfhtc7jVIDRnTChLU45b3V/yM+J50AOA1nLn7qJQfgQwmZKyXfxYt
K6sOB9ZIOnZ3CCn2wmvjJIAQS63n661b0iRD8A/x6SNlUgCZBWx4w2pXOsxDMr9x
ycxVUKVUmjG7ZKGZJOEpGOTa4MjVGbIoavIeAw3hAnVW1RiinsQM27pysDdNmqkb
UqtpF9naGLmf4rQ02FGybl/a1vqt+zFkiUwe8DBFMASoTSJiN5Yxs5Yg+SqezHjC
gMy1FrCk0TcTMsKyR+aSevMfq/Odo95kcQMR5YoMdikxybw+hABHDtQAfZR/t15x
XSScdKaLQJgZ+mZ9jDXhzpGv9kUIu2BQQnpyPIn0NQJA2qIRq5n6vAbmM5uQzAff
0BVtJTC+kWRcc9Jt9E9bMi3TNlOJJCLxJbU403sfE0bJbI69MyvDdiH81MiQfY23
oMp8IKwWdc2eCmCDfofym9brk9T3xkktS8/s8XKgiP5Jnv7yQ+5lMFkS5fgKM9jH
QWFl2L+YrpkpK8ueU2pnNPIrWzmYScg7A/eA7wWukOIEeRjfSt5qCFzhEIV6Z5nc
FERq8nt+q3zgrWBwAHxKt9uR+QDvuckXAgvnohUE/2wMi7ayWu8moFD6PpsgN9wM
xzppm6Sxs1xquhPehZ62oNyv3w17wAQaCB5AjiSOXiQXS1em04RfaymIgY3nP+UI
t7H2BGciAsvN0DI9zdDgsLQsgrELqteLd08t/u5+4s9wDL+slS8FU8cFQ4OR2AO4
uoIVHYecVIGom/q9i08ZKqRJ4vZWy4HYMehbWQAUfD+GlCytPudmMsEhyUjsL9Sb
vOZQTT1xZYNoV728zG8/dW/UCIwS5LmuUd39Bb/ppmNcNVm2zkphUlSMWcMNX2gb
pMFF7DEBGD6FcZaXn+uXP7g3W7ksT98bkPn7sP+xHZZbaq+kTUCdEQpJDdOsZx/P
qUWvqIGt/zQ9l6JM1e1DeXrPXpywGavCLv3bjUKgnGKae6vu/5Q5RrIYOPs7Mt5M
aZ+2wJgokabxfWU339yRdZ3/8ZiRhpAqiLkqgdOJuoMCS7j52WBurQIywmSEM0pE
FB+AwhIcGm2DG7yvUuunpT9kwPZTSTmarZ9yjk4SvSv4mXwhGAwxBGWIL7WkuVth
oebX7VPNjqcbc3bBI1ZLudB/0WuXPA5FCHWwFhIXxF2wkRbpwJj1GjW099HTT9Fu
aTEPH8s0ZjhvLVS7Mhhh+XfxKy99I9EoyxoHL6lIbuKW6tkdGuRQZiYXONu0VoqS
Lq2Cm3mph9YXortes+n8qSXa0sQUfTjEPET5VR2Kbx9Kv03kGM0ABCkEPw8darJV
CzmQGDRPiYNJyLE9OB7PU7Hcm71tf2Uy3NrqpXzgztNFQqQahNuZ3VqbqiwqU1eB
mHQe/UyIBZQz1ZEfD01BzNq3tJQmr0DKRfD28eDSBnyLFG7zYaPZeS0AKfuIzRii
w0Z/ZSrBFDWkiGSdr/eb7Hkb1bq81VVXlgs7Yv3EvVhmtj+hxj5dmdq495my+A7Z
XjWBo9B6YFWAFKLw/ue1XfmS9RS2T4syRxUGtjTO+KFq32PqjzkbWR5UqqRv5vRW
HvQHFLRJJrq4/8YIsW9x38Uxddsp3tk6ZGzaYA7vomVxIZKQl8NCoeMMS50D/GnG
3FyEwGqSltDb59gELXDp4RE7Zu8tSG5UiO6b5alNoS6Be5xww/n/sruXXjHqJH+a
Bscj0pwTUUHCEYDE8d/qg6uDFOn9Zc63STbREwjx+KIRDm6vlwBvTaSBoZyBqmVv
oBELsckUwj6VirnZmNsMW3HCfXQBOPsohCRJkTLJZbEQVC3IYveMk97kyhyx1+8+
OKuIBh0lOqvqGnyoAPvxHH4oebcR/vCipS4q+NOxkICyorlbNsyvaWnAKoBiU7Ag
MkQGVfy7IpIKeZJ2rCUQLKPMseroTo7bwRf5ivCBJI5CWl/GOZoMl/fhji2id2KZ
emv4e4lQGLg0fmxN+j/caLRFdTYBBnjMihF9wIpA/LMRSD+5TONCZQZPWaWg1BF/
1r8gTKm23rTS4eMZTc4wnKum6KTw61lChOPqD1klIqxXM7o0JGEvgpogp9mcE8oV
IV7UWh+PsMs0pcHHEQkLazIhKMyjjEG5aKiDlBJ4fl8WSnZVI8X48vxRv61IOfxG
Zd9h8nCzcNSa7saVEFywJrb1sG2kRPKxOzLC+3rkf6zUg8XROb0vXrl1Xf/m8JaB
W1DIfxCjnf0K7muJXqFluydHU6LSFYwRMBcu8URHOB57qSI+gq1IPQSQ1QmhOVU0
B/ZUJrrnUbBzCdYAhurQEmtQPSfjSK1lPZvjo3rHl9snVgXnAdk0m0d8sQDVI1pT
ph6hvV9ZLazoKNRRUygQCH81maHQ8ZwBSh9qe9lUEzrBn6/BTo2AQJAWYZ7YbazJ
3fiUlVxOcokAHwXo5WW9bljM3UiOykFxvL8fa8PPgBLTVRnVWavYH623SpULbJIL
eeglA2i2sRh3qrX7JUD8ixkY1eD8Cxy0MR/Ymd2dnBn3LGoo2J3KlaRcpAwyn4Dp
0vozbAzZt54BHGkvlmlaMQe8SQOoAoBC1wGbOX+3y79lH7cKMgvgkRmJelWSI8AZ
a0x7iHXsz17TFwutfZhimAaxNH3ZfG5dgR8BivWWTPw1s34d/9DlfhW2xbB5Tuqv
LMwPfVye+6bKI/EhYLdQH7hQ3rT/Fny5wYyu8KHtV07HyuwRuyRPYHwMFAvVb+HW
F9FXIBuQ+GGDoBMWFGk3psRGitOw4qHCEJjARdkK5f57Uu9Na+MS925laUWf5jsL
O2cqziMG5nWODZ1Jw/+wxJsKd/HBFO712b4ESINmkKjMgu6pIin80SOefwLbuoLt
XL5ea5GRnwwS604s7hU17EKtg6u8RdUrOnqdJRrSqNtNQ/yuL/IPf19I/CDiR6cR
G95QVyqpbeZvV4paLHcU0wIjlbjMNrsmnqHG1yAv6xcOUh1zwRBh9mXzd7k5VQM7
BCEkeEHb0+S3c5/Ll0jud/BFAfsN1HAm4tV+hFzGteH2PUTmGFH8EzL00JgCdvdv
8slmMGI38NQEAZ03aY9fV+cfCqOTZHn44pXuv0prWQ3Igu2ezlDHjt4EURkd98jT
uS4DHgBmEHw/gOXILiPVOjjywasOazkMCC5Ip/a96/yyCoL6LJB7YriWjUkThwNy
Zm7fKV4kG2VgoebzqBNw+W79MyI3s4g8c1SohEySqIo8X1ZlnxWF8ravtprvjXTP
a4bZqQlPuc9VpD05KSsj0+xtvpvyTnVxsfVbSrUnAUkmK75xtDOYnPBH+Wt0cx5U
vPCJ/oafciADBeuft74ssUrsJ86B9yqgAqOrP7Pj1o0ntoHB5mJuwWegMRTrhC+f
jz3YOUbGpd8zV0Ey/OoOtQYfJXUJcYMLokHcPQGnscRxqfviuY14tHuin3U9zRvU
hwaGp/kZ8IWOpPt5fScgZqdrhgxNO8PrEFkDQ80M9LaSEvHiQumAqR1Oxxd6VjfD
Kae0DAII1HTvj3yOsutMOskq+qHkb1QK8ZYQMK9FNI1kS7eDqelv6bJzOiQosXWc
wR1pvmx8JXNPF0bdtPbvKc20Ep6/TwTAa/z/yVWPksMNpVjPmKI+stM03GmGwH3p
FjVkcdBUOoeOnoAHoMWr35UzOm0wmYZuY/7u6hr+Sy8DDSUG/WYUp7tnU9Emn0Xt
d3D/i56D+r78SZEm54o9zwOrsqQQjnXiDu3LbG2Q6SkRLTcDDcsghmczNr8bA8Na
xx3jjb5eukN470hF3x//NVPag8ShdNEu9NSWU+7EJuLmDwg03/KGg68cj5e7X09l
k43Wzbm9zhSWaCaaAeV5I1Ohhgr0SSpJeUUnu0U0/cMK2VyMLMTR3O2T+Q3S6T7Q
17AjPCFWtZkicL7Jo9zzuIdlMu1k1fL5twnsCQyyEnYHiMHXhE2QjVsT7YF9pvVG
cmSEKHCMCi/jMc2M7EE9l2YcfjPC9H6i2dk1u+5oTvbXcPT9OveXHdExK7VsqanM
Im4wx1fWmPAcrHLtiV9kD5gOu1VPpnGnjVDFuyM81NmEqa8SXpQkZi+3cLM+gp2X
N60ofpqlHwUcQetnOfc86uIz1ZSZ0A6aTGXnqJMNIGOOR2Dph6pB/f3KDtbbj1J8
tIUKQyP0jadRBAwcbJLRIu8jGa1X81XXalMYYVKsyflWrH11SC5rkroQ4K+gHVda
ymNdRQudoFiOVEIoe5cIIwhJOlGD4RTRZIv+S0sKBtXyX5AJeUdh5F4RA+C7yntY
9FczkVOkJUeahjG0O68RVdmm9M/xnOQJYO/2djJ0+xD7kVm1sb1RtA30yECCxD0w
br2DlzcbF3c1Cxs4d3YUvNX5Scm9LoupH0c/7DA1Rcy4ovYFu27iaHWjrwdKZZIK
LgnFZ01S0ASz4YbcZSLl7R6uWIkg2Hi26FTL4ug4hzzh/EEW2F6ljN8gEggPFew4
pd3cAX9kKo5jMeh76cUQDAE3ROeOXDOsRzGe7eUyCo3e5iMRvCztyRjPZYACJj35
WRXc+jU7oOcYOKBq1wOcW0roCROHXWeQk5cR0QmHj82ucsx8nFbqn7vS98Py33Zj
HB6Skoi6kIpUJ7JlO8Owt/F3SFu0ZKL2zBOOPGCPYKwASiLubeEbNPhhP+VzQYtf
EVggpRKADxD01WPw/mxnROr3nnq/h1ZFX7YT4Y9mkl+pEX0aDZz5rr4TEyiLcS1e
rqNHp+JDgMKQ73DgVBDToM3zXl5lxER4K3JD6XKvMVaNHZvkHiWT6qVab4H9L/gi
SRZ6AYJMNPK5PiRzo8ccPhcetHonA5nhS5kvUbxFGHxpIIY2o6LDbO844Pes8Y6Y
MvwCvuy62jKzfgoVVu2UYi+yCQQ7eF/+5CCF04KfRGiMObD8oOzq/DkoDHaqmnMD
G1bHeQ9j7vZukWJoeLC7+Gh9iRFRGzVM3puiN2jKz5hClB4C72h8sYW2JP5QQy+9
waNGNm5MUdJ3AUnOfYbIHGnh3MtqGX95TEQQ6lF4HFWlhaTtKulJSBXVNPSbYzlS
0PIV24QRqXCmzQfSJcqGLC6n91HwLzBRVEkdkGRgIQ8zXfzMPaCgVu61tEAzvHpV
XJ9Icbtsk9bGkRmzq8k0o22ADXYiL/B8LoTMrtZp+rAg7FVr37LxjTAGXAZMkNgA
NBRFelKjNlq4KIbrvLtBmXSkq5Tniue9cMaEpl4EuMDggUjZPUJclmOAV89h14NO
Rqde/d9OKUE2HbVtwEnvgJ7XBbE88XLs5XrIfj44TU/FnI3NiEHth2G5vJG9Mvee
334oXb82w5N3MRntYQUhPeDPsKX1WOXaUJFhcMsAtV4mjGIiqRuIK+rscagUKurR
6kQ0oSmsJ16h/G9LG3fuFxvtVB7RD/NNFFIXgWtfRa4ybSFvpcTQOLqNWB1VEfWG
6oA/RUNsbWEJmWGNbBhpHJbsi9K+1+brcDs9LfSkp+30EJo/L/4ZgFZAQPO7GAUt
vp3QanKHq2mj/gIhBaLzAnYawEqLc4oBj0tS6YCA2ovFFBhrkDhBza1BuxML6bsX
4H8OU23ST3kHM0S9qu+qsGljiRitWB8QYPGXq8zGid08ihvQ74aWjeH7rQNezoaP
nCqDs1VRF+Q4HZtuETXx2/ZBBlEwLCDgBShsrMcq07kaInTI9EULCKFV9xagGmxR
gdK6mnicfEoXtECWwt638kgOThhrwPU6pSLgY7GBAdeN9zzBrLWwKfK0E4x3qBxI
/hCKer4Cjx+AKk1DbR2zVVwqqc124skcbhTOex+oKdV+USSc9PUn/KokqQ0TzS6G
mloBq26VlzXxQzoajoYikdt1Op7jCYg84GIl6WXjO9P03Rx+zyMJj0079NIL2Qf/
7lIRXa5TCCO/DUTshwRoQ2JXe1ziEl2UrYFYVqo59G0PDGSnUDq1t01iNoto2vIu
vZZpEZAEQSAtpjOAgKXKzjmV8kkLmF/5g/6J57tYldUqcN0s1oHre1g1yTnE3J2k
0A1ZDtJflVD6wcdnZKQK5BwwMZFlwAQqZtfCBod8/mkEP2QTN6Aw0Z0qp6JekV+E
YFjjbL/8+WePbGp3htpVi/jiUcJQqdmYFJMMPRnSAr96Mm7lu9wjiB8CMJPnlLdE
MOMb/3ok8PAagz9Vi4QKP0oNZGhp10ZzEGZXKw5saDrqtM/Qgfs18XKgckjPAjes
jqKkexTAMJFyrh3F5NBG9gthD3GlGT6iOisG/8wIID49oKxyZ+c2eEkv1cs5munS
SxhiH9Cjo4F7qofyUcb/lOPZHX+G2QHDl5zzbYLF3gWN6eTE/fr1qD83359NEbv5
e6R/NoclQoqiFSvo6i1WSz8HRluypEWIiltTholFf0VfUAkp9bPUWBuFeUnrcjeH
hBw+ajXuVGnH4ORMycANkY79TzJbgCVovN9zofBvV5QY15Ei99zDDP8LksrEu1PK
y/xeG+I85qDlgRmgPE+8LEi8mKKtkDRKAII9tbrK8N2yaO2l89fdq3D3viK12m3V
xbnG/ZdEZ09lDj9QtLVOP8ZnUTOWZgZ9j5KlVeN0yKAFA7G6zBujDVyfWSKX+jkp
z9mnLTQD3Ei1uQwcxzvflepNCXV7a2lLdvxgUMmJLg2m696rIe28RrL8qfV4MZT0
3wXQqKjpOYOzMBkIK/3SpxdLpAu63PjscUOYVvM9GMYasbmweymZdDKG2BMTLvDX
Dl4oa3w6BkEk2v8qv8entJgpwqsjQTz4D0Rhe0SqeJ5mh0Kn+GEbPkkSJIiQ1hWp
gSwCZ/qfz5lZ+bLL6mvjxsq4pa+9UhVfX2TFKtq6ZU2ki1Os7cSfpRmz505wn/YR
cvHA4i3TTfRqsG+H/+ssqlwqklauS54VDKjUkWx3/qZdXCUt6YwpFl66iRdZR6Cf
DecUeRYxBu71mUscaOcH99z3vMlHMaqqAjowpPK6Cj1sUi+Y883s1pmk8powFwc5
/R2Y86URUh4geDIT5ZvTtm52TllG3yoQhVXt4BAYA9x3rKoCN/5oz9dOykISjGKE
PuuOjcIPP10rliExuLTE7FXE75N5vlyyE7P7Ks6t6pgPaXtBUsE5LVrqW2j9CKEi
DRAng3mHIwmXRDkPjvVU+kfCCbYE2K548TQSsqlv/0vMRwBZAo1A3aJq0dlBSnDF
bZ+A9OsFau25ByVj5iIxZ1AOXts7yFlqfN9ulx3+SbINzrBAwJO7H3QEpZF9SvxC
R00uxGesQB+ulzWZRC9GGiRmXf4VieYcZeJlXJuZRTh6IfzyqmoNAoYAbSl8+qFi
FXFdDnza8d9MNF0CAdg3YrcSk0ctSLcqxAi06cegfEcZjTrSecV2zaHXfiPawmKG
cPaLEyHp1YzEgG0H99usgC6oxuLIkHRn/4DroONzCPqO3DAcNfyl/p+hClnh6ska
2GztQl7HDCpol4lQbMuRgHmP1afvMbP8zBiqhsY59y65Xpj6f7Q8F0dud6GXMiBW
0VwyUiMl0I9ltB62B9RGGzz0eHd8bjtwcf3oNrQsell/emOb6gKmCAdleCAcJBjl
OByvsk1EjuBtUikbyio6h/E7daN8a/Foq5TCwe9cbe+8GIQA0n6opRSkH9wxSDS/
jiBXjELkzn6gBVIOfPotvPLDkv/XL6xzWuKvPi9UUy+qmj+8gfB3ss4p+BjX9tnZ
pYf0TKHDtZjjRYFUgfQJ5zVIZwLllctukie83bgiPg5LWGhrJXpSv9Np4Zl8MBH1
invrDJdygbo5j/5gBXKopQnusPUDC+uGsEy+zuSGDZ7pNqHSUvS7iWgjWIwam8Hq
cjeuUOOSrWhEXl7q/boT+piJw8CxV03cBccjnd3cbb1M69OTTIfLg3xEJ1m2eYZv
8OVVk5NMmhl2vcsWf+muIkrP36v2Uxm2Il89hmBbnmaH7YjqFNTEUexUYNypvhoR
Jc0W5NONr82Tx1AAwB+UkpIy11Sgbc3ybG4Qpy/FmOqBM9Y+LgnpmuOAxsMwvVdv
BHNibLL/dylZ5qoJD+cmEJ5G9Cuu+FjAMNu0NmX+sMClv3fUbjxnTmyLRIJlgm7x
QOQ3HObkEeU4ibu+7G2lJfw6t7SM9kU11JrI3trXNNm6Yn4wBAOqyxh3rS8VHVWT
hhTAzAbseCvabphM74uQ5wPrC/cfE3FM1MEWiBeGp+1naP1xX8gakP34FbYS5p1G
S6r6nwIMu18ipYLySCPWqy56gGtnjF0J0I8mDZKWI89v+mLs9YZPwiQUCNdyHmRm
qiEetiwvTbgP89o9QOzj2qV4rC9/YjK/E4OAQ3uick/qTB7/0I4fCK/KKO0SpZME
0tg+z3hv+fo7YWDLxCurmkqegQPbP1b1FG4m2nD4wHD6ETVjZs4fGY3zoiaTBWB4
vW0gfC5AjXTDWlJBsSKCI4+SkPGwPiwMojsWXG70iwSq46yJmojfXtK5ICOKfxkc
5Upv5Kjc+wWOjZUR0TgBuc1b2A7v4T6figQWj2o4RghcYfdOIl+ne1lQE8vr3110
PPPTp/2B3IS7/7d0IXJEyZXYIYJ6nKf2OE5KeHAtxDaw0VHtBfqXtq57q2P3Zv9N
tJJlOckV+65agVXM2iK+4V5AaRhmDEGDhiWL+RqlutYYwT/s6a5MFmHnZ3Oo8Zi+
ZE/FbnWTHuthaGQTbZ/A/zEe0VZ+nvQcZIADJkfJeAxVxsonwGyyNPv4cADCQGFP
S+u6J788UDACJG2fOor2sDqrrx4vpgViu8ZIX4saL9nyYu8cpyW6PbtmnENiKLJh
svdQyksLH1SMeY4SYB6QTwzNVRWF1ZE35EP5mk4VM2a2tdDrwwENMFNknzqyrOOJ
fUsn/blu7Lb/Vp3+mEl77I086esQGPeqHTGKBVtnBThe8o8coPremkUxqW2iS7OH
FwFHprLgF4Ksnp/rsIqnPwdHj7I6tfRE/8gLwHdYwIy2ohWzkWhab8XakkrCWv3T
2nCtk6wJxya7NnCR86y4toxTQr4ou7Z/o3hwxm63GjBuq+8C/jLe43dnbMEyFj26
2LeD3+caU0QGNtliO2ZalLC/Xh99QQ+klpyUur+JO2E8A0FSz5bkOSmku6hDY93p
7KyfNbFWEhmoQp9zzAXuo+Q3dwLSgxBKRTc1uoPDhPDPtnVNchSCaPmFxkWsG6WV
I4OFmU+uZY4Ui6BSMxGeppUE/QwhalihoW5QvTNOKLgBCJw42WZuBhHy47E2GZkI
g1meyAplmVGy0ZVZ2piDN3UG3sG8T8luftMndbw9tae+TdSin+Hrr8htfKyIFiCb
iT0cwHvoZfN11rTeZM2Z9l/j5FKshLzb5XQ+xPEHS3ia1mlO9xEA+7JVZWzwB4TQ
P11NjP2bUPG/86ega/9emzmwgKNkBCUvAo7MlurmhOPZgyiWO5jWeN0pTxkIB8zL
AJngGK1x9ZcOFb87MDU6JFL3TjLocjO9vs8kv4/05Ds3FTWBMEz0F51J1GhkEaz1
RzPmdwjoEc/HRvZhF0pi7cJkADu1/54X8OPMwdQxJc6kDyPZVs4jPt7/MgMxHGOU
Vh4Qwae3mNdOv6Yx279+nDQHUa7JIPKatE/+R4K8d/igJO9w4WDcCfxbcNobDHan
SlSl7EsnW28Fiz31wcghQNvxM4SU531ZgHWj8c/hdAkDGpNHTyQncQuHn1KebhIX
r91sxh/ASrkpyxbxBXab9ndDgdzyg9oyM5iPqg5F9oVh5OPfP9xBm3r76N7SxT0t
XR/fN5whYaFjwnDd/bUoEpAkvGaGGr0XS3EYNsmyOiI9OqWjulVhzllVRmoZ4GvD
usT+iCJrRih1hAACI28pDRqzMtunHwHsdObK0EZUK1MJAdzpp30orth6J4ebXvBy
wgHvLfnWnT4BbNtS/4sQQN2Dxw2q1LkgduL6BpvxpWsaXGxYX+bJuNb2e3/kp2V7
TMKlww/SS8hQ4mfICP7TYPrA622V7tRF5gI/41bLUM56ECSEvYgXHr2iwQRhRWRK
XP5KXBHKVkoUBGnwzOzwkKmwxkCWNrUkbtJZ12QhwgL1HD35ngaKp6thROWv7vzb
bwImbEKYOpATFHymG5SVf9Db64MW6ig1TMUvywonWP3hhTnX9RPBedtbMU5Q0X+c
E5DyIHuJTFSMqWx541U2CIvc7fFVouZAVRihe7M+aS3vSQ0h3O5p7ENNvgo6++rV
kav2juoHDA/q9tL78t8i51BIW14sk85YYOtv4ID9KwdCCL8vbAp5/YbbM+7OWEEB
eVt5UTH3rALdxtd/nliANjJbqfCC0wHMCagHDked3pRGlUdZ9w5kLZwWM/KaSpA4
fJ/zvca1dFI2UD4qtiKMwgaAJ4qSHXWl5sdIWlcJdBjtV1I/PTGtyobPpN0J3F3j
oaZQfhB11C9uRe0wnJUsfioRFNr+QhMmKJUjKQD2yHyqAebenaofaKGtSqnabjwj
/xlMm/iK6zssrFCezR8sPXT0nxDSFtqLAk3gnRDXXZvkQ6MaGCdzbhn5yXuZ6JBD
gdLs0TZkHAkYxnfiQe7Frm8wkIeABSo7H7PjL9xmMXLrpjRbB+q1NxHPyG8WIrwK
jw2xuehRi3my68jpgX9Aj3zXmXYPOkT5VnK+LvadqtL1g3pXg2zBzpop1IerKjot
228ChJM3OH5YRIQIRjklfLxSAFntOFDtC3qvLjsi3G/PwDCs1wvEBXI2EH7TQLhm
mw7D+sOSBSmZwPPhT7o6Rw0OOCkSQVKSlUj0XPDwpuZQbp/VnLjnss+14UKhMdQR
rtJhbOqSlkoUdti0krzCHgcy8I0ZePd+rsPG8dAe44k3K/lWDGHD/Hs2vIKBlZgJ
woE2eUyOjnvN6omD/cvu/W3DFvmW03VrENnoIfwNlK1YJGtrTIOQEnVrbMvmti+s
b9LIw1VUZMR/kqH06TNJN6cVDJjU9MwhzViouC113NEmtbdWOFXhaKwgR0xqojdR
o3BQ/U62NKdIKZrAfcLUPswQRnneR1p+K9yN64FAPPojUuz2hBeiiIqwL80JnkNp
t6GE06RrArVCQ0DaJpuJCaHCb7vJC1u///SJBWCXlJ1TVI5bAfSuDS6HpeDwzjGR
gOJmcJL3YC964I5uUU+4Ol/ZTcGsMRbcGZSoKraLaXDo710E/5B0PXPLyp0Bw+c9
+raCXj6OYdCVCc4MWnVxYB9d/Y7jG/ngnAmWhi6O+lKmNsoEdh+YPHTV4tSiej1y
VCYzdsAYofPbA54QEtDeVC2HPxYALdOkHCOe7moQu7nOJ0r1eR+tePHVIZ+G8+bX
vcZfN5vkyqZu7uO3hb8ui3dHrqVJ+FIFFAxIlYNs086nVKW79eSaWFLXiBac7hv5
GMuQca/TfOhfaCXL0fBI92GD8iL1bwW++ySK/CiITHkGw1iBXf5IjvzGlZeM0dvE
v/UkKuG3BzQwBtoK3hKLBXKqI8TPLuUcSi1BCTBvZA/4ARXwtPyjs07NZ1A5nFmc
HrgCPoqT2PY4SdTj35HQVnSe2jy92YndZ5WQOAxl/j0OY+CDzvPHTae1FMmyd/ah
raQG6wTInyohs9P8Z6cXs1ReL9YvQosBgPQgwGRcA0ZKT+HNFuVB7cCVrCVisxwe
VVTPgg5poI0WpQykmGw9vxE+ThZgB6CR9rm9C+/qr2gMGNrNY/ELpULDgrloINp0
b7fbOvgGMOAWCDawCVJgpJzH9Z5yngL9scYjYsgF4rybkJwMyxmwAgOsadhNJg5r
1C6SGmy8SqmBRNfM4KH8KCumYQMpsa5qvJYbDdt0GvfJlV2elsNWUkF6drW8YBL3
l18OCkxM0wLaEFF64YOJihsI8XvVQnWMtM0nBijMrZnUfAHM/aHBvbYSNbf6iSoY
XudM16zoAf34mZoUP9YWgGIe6e0vCGmIg/OZ2dC89tcNtvjbrHpEsBXBmDrYbi+Y
qnioj4Q5Irw3N8y+WlctIEf1g74MxxYnOtb1CbGSbChloo3b1K65dpPf6xbTXKDQ
5UtzOYPvgiM066wdQgB/ttp0qNok1Lm6V49JjPHZf2Ij1RzBsAZ7LQt4iNP0iuSA
qUQmc7JkfCpODFax0lj6ZexK7NkLcZtEGfdsko2+IlnXVj5xjL2WzetkPLixzVwX
puLIBCYbm1ivbJQ94HymXm9WMnBDT4dh1S9KlouDhLemn6eSzSmPYfRHxfKQmFhc
4BHnVLd7bfMKrJpJSSVg7J2OZjs4GdDb1F68jM5m+Co2uiHwjwqQpqKsnGFfpuyT
P2vY6n0NzRGyeTCM/NfHzqUTvZO1Cw5Ybwaj468YgeOMGHJZgDx+/2WWV7s/ITzB
/tPG2BpsaEqfRcyvWRHQaZmYcjRpdE7Nrj5/rZ3geOwYUhH31zQuVjB03EhhiRsL
xt+9g6iF3QQQ9WQHDSsXYx/o9JJrFWwa3WrkgGZFtvfB6bwK9Gd8kdoc+UNttyeH
yJPa9F1JsD9iHosRaFXos57cglADTwDZihsAcvSa+L/Zi93DEQW8A4IDgbueXcqV
VOnCSiFPykjRJLqW82M79276U8P3FLpcZufvvJaTEx4dFzyQnZt0GI2xfMA3ELAT
P5SAg83N/VDZoR4yAggGR22c+8me/tkOgFhrpUP78OXB3qI8BPEPSBLhWDYgKs1Q
sueRv+RbyCI1MuKBf3Mr3oAuv6SNbOoAK6ov4gBv4djzx9tJb6oyjenjxBVj8B5x
cqMOu+bKihceAFtLTI6fO5OBcYZ9yNvgCfxWT94z/r9PkQkht62l/o+dKQC9m9sS
lklvDUusbkd/DE5M7fLoE2S6l12d/uEQGmaUl7Oz4kWGUc/dfGFpdauM7I5IUUSJ
Bd6XMWzaTMibSB38UAjg7YdHD/ihEdYHPv3EuVgN8+mqQLqWT1hcgr24R7BnnLHR
2ZuoxnvjpqiYix9Q6p8Mt+uxaa3O+40haDl+Eknv/8okj2A6ZJgLmnG6BmSSDa+Q
ZR10ZUmQVgF1tZ9YblbiGgnsW2gUyvUMUIRJcxt9EP44rTq16hOIWOUFHe+kGMLo
ZXhxHlD+RR+2S2Pl5ZyTfvvvQ5BVRb4n6MbgmApH0H9+LTPT63Puj/ibEU72AHId
LF6EsyuZ3aHvfmQAYxaqF/iDg5vlMoJjqwTuNJH9mwWzkT07HXylA8XjvhWvoPLy
gUlVY2NnwT5CKn2GAjTREhrPe3M2Br/X7FwA6JFyDDPQQ7crY2HyVobYYVG4B8F3
wj8LswzmQw3c5DCUgaEst4L/Eom1Tvf9SWy7GllznA9SneRhOMFOTLBUWhXKxk5l
ooCAwEbX1EG9XCtR4kYZ9/wcR9ZubZymiu1E7XWF5B7BDquUfLJXNaQ9E3o8RTSH
UmGzyfjo2pozfQwpIdNfasXDQ2GLF81v0h0KUkSDceCCHepkgVK6Km4PZWVZMM7I
6gK7swzLAZD7a6RYx9IP1O0X8ZsYlza6D9YA7u0tzMUpDAElXxPQsbrJwEZSFkH+
mJOhXFM+oTr9e2ILGapFsI+5GcQsorJKyf+rxmQriC7VJ+cIclH2tC/eAGNvBWme
dN+W938U03C8eWckiSSS4njRq7qAEu/6o0zCgx384fDUJWhe30+HB2xRz3xJaxnq
bKm5b54gI/711J1ZVOTfg8QS5CbtOyhnx54rt+qBGb3JtBrsOfvcOc6dbBBTcIXq
l7wT/Bu6pMtLTKre3/CJHz2KtPIGHU5yKlpTH1F7P6ZHidJDmPPb07ettFsXdxra
SrnlGhJ1SkzzcsXLxymTaavB/hLbNjsUF/e0F3OJd39ajP7aSYK2lyWqwdHcRQSd
Iqaxj8H+pj/lrhom0kECJG45IzO0AhmJ9TV9yydaHHu5U0hKzme+5Ce+0Lpk5nVH
b1IezwXCKBngXfVkkG31wEZIBNIZw4fN4FzkRRErTcwF0bgIS0QWc5Ohd7PUHWre
Cz06ldp7Wrh+APlH6DOgUUmsPikN2iBAGUzophZGS+k+t+MABFIZRhyO2CC/kIVb
dxwnlrkufQdroFdqKaQ+7iGxtiKhk3LJ4RqTSvwXMH72YCXppCsrz4ZpYIqbAvSN
VWxi+QvwEyx8Xg1Ee2pEZGxBA+3PuyD5LDO/HxK1cNxgjaTV9Cu7wXOXPbYsGaZz
DeZssnXPr2YyqTNLIJVWvwRQfNMzUxad+VQja8E3Ezoq7NA665W+djhdJDOP4Nnn
uau6AKfaE+xXLHFUxex9qMobC6hLV4tgq8hzZyZWKqNE1mQblL0v+HpeWNiJT/4K
rcHhqgpAfrg+czgVWgcA08kKgB4CBYF4XVkL3esh+l1xqe54TDWYAv5pKjHLgeCb
Mv/g2b0AYz+JQSFhfy7OgBRJv9g6tl+GXXpbIVJJ3ba6FrGV+utcioXpGJM1RQve
9xHVsBjeGucqgN1GCYW5lGus8su6aF9SDKxpylq4+tNmCpo2D+n+NVBHi3mSRP5+
xMt2FCfUTSrX0RZ6Sj9FBcXkEkt5kPrrf8XVk7v4gzBB8hVcBRZKZ4uT/WMjCam3
GD2X4bsipnToQVyPVHrfu/k8uRBQIzv4g3q1vhud2HPYYeLZnVGFTvLLEwYoE2fD
EGYzWR+HeLaDlbmKkWjj2FdJZzhGAOwqn0AdyhGH4YH7bRwJGbvtbyNXDwLLV+ML
VIViDvCmBbkx0LyvIyOM3ICoE6qno7rWmHAfxZotZ4qS5ROF5jFZafbMcMhJLLmH
fQnADQxUr/aJWsA0nRDRiHzHMrJFVxYV5VB9wddL99tG3Z0P4OXzrTOCzmMcMB+E
WLH4RnqY5OGsXWlePJw6VMlh0ly/0TZ1u0S7V4yVnVOKIivzyB3elG85kBjt7RhZ
Fib8RmuV9Jey+kIu1vucwL05yth926n6FDRq2qluHrUuZXn2H5Fc/c0qPkEGpqAp
Hq9o2CSLSQ1srDNLgOyFZn5b1fpKpdQ/G9Jyd0Db232+71ZsWGPCcTgBzI0Z4OzK
4LZx5vXw79XeMrTQisMFM0u50IDOuMdnoC69Q0lZhWXD91joELe/IRjUpeF2DB23
Xp2dHiw3b25cmsymVZ5+wlSFr2NaFPZ/9lASCWVo++wGQaDqqxZnNoSs/en1747P
85DrscaL122tS+EDqd0hF0N7BIupCLSsbvOXngDyJSvnLveith5ai4QfIK3zZ/ve
+I1b/m3ziY771g9iVtz4zrGEJf/1aT7I9M5NsYCj6/zQWzkkMpeITv3Nb4DTD+8u
njr/Zw4xh/tuzE3p0NBzycteRhQkSlQ3EZAFclVieHn1TYX2f0K8rkgd430HZh7t
UAWyBh7RXjqIoNfapcD34nhLH+06i150wMw6mHchC4pL0dDwqr32y0QfGtG92Aa0
eJfPurw7XI/x0+QG3UWynTe6V7UHjsJ9WiHj8nTl8f5XT3UqxOBFn01S5M8pgRK3
CkkznobHD+i2UbPSEyGlh8fgmjd0CXI5u6FhEjcoVq1ciij3DnO/pRUMEVSH71FO
UmHIm5o1YsEGN/M7xoUycrB+fDhVG65qlZfHX4pg29yAwIVwZa+UDACtjJLf9Ugk
kFQ+fZydu9K4/oSlzJHlOUTgjfFUHzBVmVrVywlevjfqcc/yxAK1r4VwhLKE0P56
xir96X0wYpnvQuEZF6sOtXncTF0G+55cW/W81wpeMtsp+jxeX3FBRDYeo38KNcEW
CqngXbBMSpLpja39oozt1Y2Y6jO9YuJtGnPKJU1wR/ZnQ7coIqccv86yXKkLdzeA
nPU3YAy+xCgpTCAmLOJYxACPj0PMmPZarkMtOh///1tCkUKYB5jWHFJHMNNEIIJe
Mm4WBwQO7/ZZG6gQbLX8D1ZRYx3u+by26h49O1G9bRMwrfYrFDrJOG5DsB3wug2I
ydZ4RSpWm/nu91vnSNV873n7QZ64vJHzRdjLu3VawekV4ZnwyFIFv2r+PBV5EUjR
ZYVpB/Aglf456+380dR2dxYZvqqraQPmChCDow2xzxnZeiORl2DOV3CxoEzmZv7o
IToMjLZhCDTMmd7+sbimf4KlwlVPRPLOAlzNBkFlSgB1kJlezpxn/A1+2ZI4dqn/
vXcuSRcxNnXU1p9nGIMmFukafTz6y2FCNc3r/WsEiBx49gO68ttV9VjLEOiCigJi
akDEEa/tW0ONAkPiaSiMIcWRlRkgr5h2fl6DxotxsyCvk+yodGrUi/ibgnnqvYfw
NJI56DnFAODjX3VEvaCbLcauu3J3wQqGTNG5ToJXLSD83kTCTfsX5pnUTCennSen
/YUac0T62LLQGQL80SMV0IUImkoWt47hWB9iELAKA2i0qrZF30CutKzLvv8tmKg+
jo9qx8XU/87Yt7Yd+P2KI/YrPpq0y/StkdhWF5yqkA/NhiWNO3M4O49++orOTtYh
EEQND7gr0jAP8OfOo1jseDvt5jXHS2NIP4wRaxlN1IuZpHK/kvZ3k6PP/IjCSCPF
BbHbzPEGpgBfvmHZLaMKmP0CojXddmupqBb/1lcf3tz9ctMTgjld89GafDYEpD1K
h5shTiv21c2/rRXB44zoSLtLNWKC/E70Qqxq81/R40YKJZAJnwhWHmqEZc0AAB1s
GSDH13M5r4mW0S+dNS7zApCQRQ2emDLPupdK+MZZ+F02qQBREJqvwwRpYeNo2dko
Q0rS8d9tQNxTRoH75Mxao6MiiepgydzkNqgmp0TxCgM2r4VnbBUnCZmJXmObG+RL
rhUl5Ch1MBThjZkM0r6whaqdPapNK7f7GviC3a1yVFdZlIiPA9MWw218OzCFuCW4
dTR1oNZv5WuHUU+o8Ax6VsDLdn4/VAxthNBTnFIY1NHbGkS6NitdgSW2dplZAiOc
cwntBxftcTTJFE056H6hxY4zPOEiU83eVffA9u4I+R1DyMg5mFnI7TEcs1UszSf2
X9VruQNAEqWBrzXD83r9016Wjt4wL+/D7DQk1efm3FB3kwxkgzeXxTgwGzH3K7+a
qQQYbgHSCDHApIlId5f6J0/4FRX4uZU68XWyCwk2y5l63IGMphZkoQ09ICTtYpXk
VNZvfcerhAyrPwZPA3IEoFisniM8/QlJB4/NWQ93aatbMZF+ahLFIqxLOFfyrcIP
QPD3FKZllGHTJwZaR6MtpdShfwIFJI6n0QI8zOU8iEqp+ybvpluLXeE1TkgPUtHF
aRKt9XmcrnKpJYQN3Z6rShgzKurevOtFy16KSPCdefjTjfpmr52FdruKh0Mi9HhK
JOiXGQbpvqhdM2qRtVAcITIa4kO3VB4FtywwTHvNMbjSTuz/OtpQR2jSRvhyDjcW
MCHSoPfrcagMPVhcaYeU7eUTxLDMEEj/2i4T9/tYvld7ltSZ7359Rt/nyCZ73cbK
x+/UHCReI9eupV8EklNF4Vg3YQZErMIVhjwfsuJZpJSQDzUqMD/q1HwSHr9FS6c8
msHcL3TqD5w9FTqYsaHU1tnl+qiiHuX4qMxpNG+szrMBsw89X98ONjodJqXqt5hF
b+EAbhohhFux2lMG/bb/QnaQiSOua8YYLywAPTG4Bdv+GC0aV093/+H4GmR7ymoB
GVcEJ6QNuvMm3PRYw9LFXEto32Ss99dMk8EvHwT1bGna2hp3g1xIaTVsX0r004QO
xQrF7URLETMUw5/gxqSYy+nvBpLZjXwOVsnK6FWWEZLRapol9lbnPbKTdhrU9dOe
8f3dvTKXskfUfEL9uWK+OhAM8HTwsuHo3m5YNXZWOV4uOCnUL6jSCNG03I3di8Id
+jdSGruuJtnOIVrToD7qxHRSyZp3ICEq3Vc2WQSFp9KDk48FEsN3U+ADRx1eF5VT
9W4fsf+umYpc4TRVl+nBuuaV+v4FuBqlIwMz4nCpsyW5nTwcRCqX5GLdFmHEUgRQ
Az/YOz5TzvQJCb2i3hnzY9b5x3k6cSa0VTpgOpc0F2pxisyM2OAxzjOftVeiOHfR
JA0SY2zXZNbg5X6bAQtpG5Cm2Spd+AWeN3hg87hxR0KEE1ozQFGuIxycZlFgqnpF
RwaWvBvDB3RXefVOoQ7nEBba8PzwI2u80swpvFCzFP3zOhfRIPNYLiHtE6x/oMLz
MBEfOg3wwxwt3UIe7zPzONvI2cbq/5sxQ3EzaMUheCKOKouw3rdodp2PNkcZ3Kap
ca83BtHoCdepnt80IGIZzANHAojMzpPOc57874NUsNLM2fLuVsb/DNnUCjkH3K3f
5zgPBTH0A2oGh0kzeqX6gs33Ej9y6ftOMxU+yXf93DIeTJC2AYPL130+4SaS/bKc
mr8BzbmpQeM7TwV2Db378/7A6sYAc83POWLD1LyqW0pZBFwFeyP6QuoZ17r3bUtK
SW6cnItn1M5zCRKq3ZQ7RXOs1QhyDl7EyWJgdmfC+ehkbF0tfJN05Lie2zOt1d+f
fefdajYkR8nBn2M7plY0kQKWL8EYCa9JmHi9qnCiGaQGzY6ZoFbbzJEpk8vomBpe
u0JspF51ek303CUaytXtLvoFFFnRb660Lnr8nH+uu/MvChSTiVBJHZsQ/bggABIP
TzqWmwhP4xuqquu3dg69xfVze5TY8X7TDaAdfCpFXQicv6WFzTNCNST8o9YGUlop
scEgobROj+XoTqxR3P3zM1b3bB+Uc/1T1Ab2UoeIihc3qRmy4b2YwUxTpfC6Tsr6
a/c5h2XSZah6gMd4XdKmo06j0f6jhegL4nhKj74JxBDoPKZg6ga09eN3okMBEI0V
MIG9XHsyvB+1vYp8980J2EHl557ZL9aMHWBdEXkeRQyZIHq+uclXoXB4rFC4V9rZ
y37QQHhS1jXB0CO/PQx6dIYoofFUB01D3S0faPDrRIqYmHyfyVQ64jp+YNMjW+/c
+pVrLt6lH6ib+JbNR3Fk57tY+zCozFB0X1NA10ImTmTz1JGMoZHt/T1Jq31roxRA
u6pwqfu/vCbHbztcs5240uUcIpbAziXfCfblQz2obdnsMCUrTKfdsDorHW/gJCJp
TzGdKjxBlCcCjHLHZBMnY/kPsu3rw0JLMt9CqR3l2SJGwX3oZxR1HeFWSd0zdGT6
t2EHQ9Ij5FvFQhRr7rOxJlYXgfgYVavx8ntfIp+qoTKa5hqCkQUdGUI9FzBv+gDz
1ebz5ny6qznBmFdTrp0IZOL280LuxPr6rjgdC6cKmWDTHpfZaJ/fXWZzyLq2s5JV
aVE1VApr2q5Q4yfDphcTzheiRhydybn27N2nBiezRYbMznWOhGVgr2Rsak0FNv8X
xun7C0Hl1EUouapsL5A2CzUS6R+bz+b50QCPim7QAhfL44ygn9j2bL3k35x+4Mqj
hvrGZK+PSYX5xyz+PoE/EVwhwPDihwosdBQ4JziSeBFy07yjcrU55bl45yxe3EG0
djB8B7qKRGCNNhRhxRVpr49JZxccSNqm1jclrftzBhqBhi2omJbmchDn3s4w0Eu/
41ktkyq4PZsAHNkF5rnS67iqoWdd74t1fkfOpJ6Xf504/Jwq27SiwqOTLRNv4Rkr
w6nxJP8UhJOzwXehPJLt5ioKMZipCiamFYVA/kCts6njR87o4gsd6DnJmtmMqTpt
G0UqFllw6f7cmgpCSeqTI/cBQqEtY6uRQz2V4Ezz1rQ3efhkpdhE7aqsFEySQ7HZ
DhkVPG+G5PSfRmxNfNgo4VyPvp1PBtPHgZ9x8KQA0uw+6QJie4vY2ZLD78tjgzSq
P6bvOCzTyjX1kYaFlIt+9D6F00CpI11Xft9ZsNtSFUNTWPgMmkfNdQi0pxtgKi+b
da86D72ie1NIKVfFxRCjrHt3rfRupZf4qd+k0GPNSCmJlDIGKtyBHv0w/vHli9bP
Thuxpjt0tC4iIg1y6O5fV9uzh2YjczTVX2yUDbbFUkQKdgPZopleHDkA+/HF7Jzr
l28ywZahEL4ByPdW/7tw0mJG/U9F0KR5Rs3k3zyqdGkOqeMEIAeeteqzfttpSVhL
YnYyK6Or2vG9CusIM0+0fXEOFU2qXNlGcWiat4XEzOzbenL4byQGgcIyw/4Ti/P5
EvkAej93WOV70btzeD9SZ7NujmWrKCX6J1XtlblEbiQTTEqCmuMnKbRfra7qjmkB
+e0rb4mcoWeLgNn+aWqXwe6W8SQn9ltlkqMrCCahL57+VGPr62DDX5k7PIvsAn9e
hi02a3FKEWivFcA+lkzt78oQ+RtVl+SPxfRdDZO7NIGmfNpK0rtlHyopPrOFIhh3
Q9+Oay9dA+BYMrEfvebAHSx8796lZhoi/Y4xlzBPpX2KDUIvOjMhLf5/ckcMahVT
jd3aSEO+99sfOBx/djNO+deTbBgD5YdBQi5T3PidnBxliOuk2NuYrdHDvIev1yCe
j79TgR5P/3pbuYr6TYm8q1Amddb+IoT7nmZ/zL1VrJNSg+AznCcyBkD3rHqBIKKN
pYqFNAlV74gd18/dkB/fZVeS6DTR8SRs2Z3YVrgTsK4IP6ZVxGOnnVXhR9uAz2Cw
sijXC8abVacvOA9TSY0g+XldSN3kkbq7j4ftD4Jenrzh3MnAGPgkfHcQQHSQ3eu9
VP07lBng2/ChfLn2HbhPUPeryPx00SBVXumr3vpss0tQLhwKamFQ2KREYwmBJGBD
E698YDyYkdXTUer4DJbY0bs/15NsmSSEMoZP9P7oC2gRuSh9DrDgXlF0NoUAk8HY
nEiFSAIs0gEO2SHR2WTe+LPzj0wh7A8K3LUQ+tYr0cf3y2wsZAsxeLaM1txKjb1F
57n7QK3jXXw0PMmt4dJWO2+AFM7bch+zcnW+Mji9nT6bmN6ajO4ajM9Ac+/9s/0s
OjmscpkLUBs5MNh6SrAljbnCwNihFuAWxm5gifkclf6hYXoMC/An2aawqmdPu0KA
pOBGPIZTcSlxoGfvymjPTJZJhhrWytNf8lZ7TICOEfYZLz+8HEPpQed+C62r/IBJ
kWvCE8m5Fg7n622i6ST4l8kvjqL40wD3lWH5N5TtNsU2G1+lRHuom//6lAUwhxSt
+FzNVcZXlyCtsOW4VAsM3uxQ2K+60QcQka4mpRaB49cgJjJz3LquDbia2S1FFK1L
2fiNvfJpkKzIyPYHlf/zXP8HdALHIEwdidnUeMB7fsXWMezlfr0Zszy1dqGGCLYu
JY7Zp+QR4jSY4oIBoQH4VsBYybHlTjLR8qHtofd4yv+NMH9RMSlQWy3mjS1ixMX0
mpnKe5PIr+LL2n7rI5zuZrWfVKgzHkSNdyNQRvveRzNgFCV+ueKO5sAB/J0SDsde
6ifdqO7wX2lReQ2AMvIo0PvaqdqakcYXIBAhbJHIVty5WSoD6Al7hs6yCSu03uCq
nna2yexvi3Ld/Wdww8HimE7kkxm+l4omQnHQR8n6Ul/1cOoIRckVrrAjZsz5fxPT
h49fKS1HJ1aVJWeYyfU7NzUpfA0B+W6SakgOxu34eGJ12CiFW9tE0AqqA+TBQLPt
bIsn12BDAfoij9v/wwLTXnT/MEwWZp3JDrR8PeYtdFbdk6tAnAor6dUs66Hif5e6
CmZ/nSmbsAPMLCgE3d0DEzLbf4c7znpnxmFdeO/yelzsfALkEFL9Adyb6lu6zGYT
TGZhd2q+L9EYDdMKjFOZvz4KQGSf7l9+eycuspH9zXzcDm5UYeX1Antcd2Bi1bsn
1g6qztnwR4C7oCAGyOTXzQ9GtNc+MB0hm6nu2fgZMtMG/OcWzLgtv1F5YS1wWySj
TPbVD/LlfgZAI1H1+/LdpmFGx9XoKbYXmu/jLv054JUdCR6Xzh3NCiZDZdvCHwQC
h8l7WIpr+/l5hMNDZN7e2NkpFFkwDlva7rR8zGaDzhy56toWOgqy+ozeOLiSpNWt
HI7LykK4NmdsDLl6OHQQN9lHEU6NbGMOxV8S6BIlUSr2YUNLeC3NLpLYVLTJg344
ZOzYgKKHTaWHkjOcWayecWNlmQ3Lah/V2zcAnuVG1KJWwf1TTRapGaFOiMVKCR22
kQhCOFpOky7166oS4Kg55lahBT6RSuOJTL5iMnNaanl8cnFFdjpcCWpcdY+n6grp
by2296/2eOJIvDi2GU2lW40q6vd1JGaUJmzAKdP7hENlSe992pE/xuk5RzbdjC5m
5KLaC6TgOakkDFLNP/U9lKoVRjM2xDt17YlgebkwTa2vyXmsBfCoqzzGtQ/UFGk6
NElXQDtpR9b15zyP6BjK56AGAjrCeI1IDW164PanScpYSo6mfDd8f1pLsFnryBaQ
f/Kwl/ap1LtJsGmYlBj+WbEl8aUfdFomgBsbYFab6hMxuJSMgzG1mhG0DsnJyIZB
89sOoXf7b+TiCE78NIKHwn2hFkQrtT6KrQEZ0XDILQU1+4xd5TdJ4v6iWGhJNNKZ
vU0jEQg6Ual06uuTs2AymlDFofKDLtpuO7fGPRbCi7Wa/ptotl6GoUagFTGX3qcU
bnnbiINYkEZ329gFhOk8uIweZFNf5C1CIj0UZao2l/qVk91+FxCrRLuGi1PoRfQc
Bg0seWcTyMEQrY9HEsu+cv7hl2rJxsNPuJ3fJfRrDUsapS4Lqeh1jkolUPXHDCD8
ram/5+9sQIDbJn2UiAb/8oTfwvtrgr/QxhmsvttfA2JTvA8KkFmcT3C3/fV8sfFA
B//qMKm7KjtKcbygpxRw1DTOHAbHgAJOxjvSdif2QUOI1wZTG7MSoRIgzBVwlrQl
V8uducacKwJB2wr3TTwit/9OtlI1GEo0O2p1Mxy5ZFTH/TjNp49pbVTgpa/C2s6H
CLFwwwiq1kiymqGDgJUSK2trYLMs8UqcOPXcGbzTD7G9HBuHoQuvWR3V8oNkxYZ9
fVIdkUftUUPH7L7lslWXEfXrECF4e3TyZlaFwW86YBQKBvohQ3iLpn1wySFZssRM
7TUIiDscPD11oitJqm92apZyA6EGSIwweNi+8EMfVNXqCd4WeDVmV+GXLsmXrLlJ
PoYPJ3sEwqNzesbQ06GONjV8+yZcZ6RkADdMywGO92IkR7SjlI20IsQ0mS95tOe2
9d1YAzullE3FEzVrpAaWTYjvB0wQDl9FXreuVYg6TQ6OWkHCuSLmgZ3Ild5XlHOJ
xR7G8sbMYImoT89YTPUVMQ/s1HNiy/BKTDQMMeyDuUFL2QvyHx4Z5P0+qaHT2DaI
gqtyHD9WjVEcZU/dDJGfhR0Xb4VVbPTPKCH4sZTKDqhJkb8SCzBdquywJfGjMbTj
dhHpfN4OvIT1k0CoyBNM99MN/6RhWuGI3HiV5iwOSiDg8QD1nq4NzpvaojUbHv+R
V9Gy08HdvmvtqX+BQTRAoXp7WfyD/Z88T4TySws+UYvJwnZAiSgxyfNzmbZHeKgG
7AekxZJaLlowymkbmwPnrdIPFHKeVXNcYPDSI9INXARmINjLKjN1kDeB/qTEhxO1
Yz1smgc9GlSouLSoxvLmU2MHjcs/mhiVPxP+QYSmCj9cRL7Zjd7v4bLskTB+iiSY
B4xLH9NyPPKeKA5AnUOTiDmv8Eo0yC0v2+ijWthx9qwKVM9dDIWItpWbLKDDQWOl
uLrHeH/ZvsS8U6JUKbyPRDgJgE1DjSwUk3/2/RSQ3V6jL6CNkDMHJ2DqkkNuG6gd
KTdvdNd+3Z1dn1wMylNfMm/g91zr+FU6Sy2rrjFyjusqZRoZrIIBIJ3PHzOpZYIH
yvOZP0XxAzXRmv1Ghm/d3wMCwWfMIyGKPDOInmpIZ96CaRvwv8lggvJsUppBUiY5
1pyAJFFS5IvpptYb0T2sl2xP0HXROKFyM8IiiyTgq1o2lPqnU7ti+w1YeKD0x2EM
AhMDEtHt6Ug1q90jlFrpU7ERDOllSfkL5AshsOf09eVszg630a1v1pRdhHvrmthZ
GuptdXlVpHvdKQRHo3XkSZihIdCp/zrxj+7G8/LU9+IjqVMRMiGzXX0HCezk3kZ3
kw8/+fKSXGDj2njCEwSJll78deORT5mb8NH88Aat298IX7Z9cDPM5OYDVlC4zS5i
nnbEvVf40KmQanQsoJSVj45ZE2ka0dVgyhbKCOOlzzuguGsK9SeezZTflkvToOwk
+VD6NL2zTO2V5OdHRjDrSL8O+0uSuXAxov5ZWojSEZUS5eshQlQ4AOTCqhB8W1Ak
eZvw+2CLEju89qK2P46+jqeHzdTVEmYpVT9D1xoQOoduQZ0nrjjYLRbDkiK4e4YI
VvGG1jzqdljUHfYBnSBedVI5H3tDyvboW6+iUS8LnLcFUuMiQilYer4pUywc/XvX
NOkhzmdf1PtJiMHpP1upSBOTSODb5vP/Nji82TS5tw3jS37uJAnTNTZ2CkPfGs3Z
7dgMOB2HkwYY+2cMmFdqBrX5faXAa1z2CCZP6IJZL8efYcGiyhZ7WBre9oZEeC5c
Kx9ZNzdCyGoNmvf2B+7ECcvJ+J/xmOKgqJCcMErzj8igkOrXzLqLfIfkhSzrheFg
zbGmgD5CkpVLKdD+L947KZGH3+YA+4fAqm6qcQ7BMJynN3tzNImTrWfKCBaJ0wI7
Nwy9BpEo2qS5WRDkorChQ8SJoFrwuOhYSPhKfVG+7I7bMN20Sx5AH2A6Yi+FqJu/
ULK5C+nXAbo/r0/J6wDBzjJYPVxw0Vy8Q8aTNl7fmoPADomr7NDnpnSSymn2BorK
ACMxObBbV2dlRraXbFwd0KtqgLlFkwr1U/tKJFDaSur2bGA7Z5DoVEknkEAexWqP
4e5PV5B5iak7OCL6U2tEPLYcqVH2kM/TyHTYJihzUuFfjQj3jtdEONNgTSJvyV8k
jK5Rl3f0GyUSb6EP74T30wnzPi9M6OnOmxH/TFFY9LBvhgql2J3rf1kUkg4R6qu4
vlKP898x/ujdaCtOpRnqx8r2byGch9MfTxt7ZEOriO9fhg7YNkvsGj5s2gHofdjB
dvzwWAvnt5iZQJNN5tYzojfRzigKTTD4ZJ8w45rz41Wl5CVw6LeVIL/61jRBmt/2
GYkr/mSsGI17Y9g0Gr46TKRM1yp81dTtnSahBCiTGkY3eNYGy3NFTLK5k8yG4Y9q
Md5HZpd0dlUBsbv5/7ZU3mJZHDL+V9n5CyJlJjg3UpVanIgNBYBXbETRYNmbyzeb
jsB4eHpMV3KEyY6psZHWiuWn8LeFFwhA9UhBykHUMkO1kEqoNhRsLFy/swRyJj63
7q5jbB1/8RNUMiEBfyhEzJzFeocycol2YC5YzvRGS5CYlTL7a7Cwz2Kcexj0sUEG
pSdxySWL6BKhEYfO+uxDIIFeTPZPeRghRCDwD3oPivtuOKsNnIpFzRbXH3HQ3pcs
YDPZoL8WNCtLswVBETGy0rwEv7JAQcu9Ca72ImgF+bebTEFV6j3lT0P3Wa5p0JKW
uB9klpi79tQ3c3TJdp9PmW9cWsvPkPTJ4N46bEJwuQzsYLrStsjbUlZCGN4qIQ1g
ICzYvrgEpRUCkySiFmey8BsFtkc70fKGzheQb15BNV6aFb39u9t6MJ0q+oX5khY8
0vv0uB8g36CQ8W3TwvuQZIw54A/sDweKQUDUOJ8BnpCqCnhRGfDIKaQmGRTIgDFN
EjoptS9iE00xyInoNwfnkg9mlIPpy1rOP1c5o/Ewv6oR3XWOEv3wkz6z5bwyGwuO
NpRcsky0art6FfHvyHpVlE8ykBQF+DyOm4oDipDYRtwhzinlHCzF1b027LmLRN0G
8oufQ3z9eRWQ04ddKSMhqDK2PUCBxzfP1p+V3W9Msr9Z3hL3GoYaEoO3Mmo1b3kC
+f7Jq7JnIb703r7I71XaLGJ02Ro4CDxzjxq0jBZYNdy2b6Kc571+sZLEVYtZDoXF
T/4NPiJPorE05nsnY+UHQDevRtLhUVH4SyK6QLQMvtV5R7dxvq54bg/C7uN+aLn5
i9/1+b2Wi0cBo/c7Wsw8res2VaXndbOcfsole9x1YSOcUq9GyovoyAdx2GBZvv6W
qFjXmskBrlaFQa1lDzFmwayH/6pL4EATyJYecvZcifA3HAaPwso5HgrsL7lwvU/n
ppSVBP70clEAg3Qc2LMMpc/tHi8hscF11tpjkhTa9n6XfebKJLT3nI6ZMQnQ8dlp
vRdSJvse0VLuh+LCa1OZDkkq2vHWAAaH4BVc274ULKLstMBs1v4oLObWtyAe9CRQ
mGh1xIiDTuQK4aOTZ89HnCQL33LD3kxrcLXiE68QN2FHle66SNAiIjQestPJi7Yp
z27a1aSOPhmTWDZKwOe1CVcQkvdvEgQansCfVsxe+0pATkB+P0QdIP+skMByNyoy
1EXwrTJVfQquh0XP54Fm/N4BtJ1duJT+YwByPb2LnYBagOTw8FrpegLSJ8ffCiFB
HrlPWOKidM7pazKHdtdc44VNDxUXiCm8Xw3HEr2X4jE/4NfH0ejy6QaZnMUfQmoa
+Okuvkc/mjD2xoUQwoZyzUzI00icFQeodPC5RR2QkuqV0Z+ttl05+1CPObiEqKv6
oOAnp/s9i95bQxxS1WlYu2TsHQfCtoi+KaUxvDaGVf3TOso4LjMjctvzmWN54nvP
qctPwGoMMgb+oVIT4E0UH3vOrlncMUsTF0rD4zmBAkIPplVJBzs5ICq7oPmk/o3N
NfrvSfaP6tuD3N4ciCpbuwBD5erWuDIkr8CO4137rIZ6UoXWZd8vXFs2waJXeA6M
uDoNOG0GBdSFonFsl0Lil/ZXSoh41d/H34ZGJLVsRvJLDzki/GyvSY3jf5HPGTKN
0R1DC+sOV3ZBKZ+e8KxaswtVsjKQYcqNKd4ogqDVOiNlsqyZRCiN8iliee9Ip7JQ
EdM50QkBInVyhXnDfnil0AnC8+kNoDdbhGomzh6ge1tZL611BIxTMffcJ0lcJ6VZ
PzRPCSNNQS2Oiou1JaUQ/bTyNQinHEYIJDYE8f/vC5+EZljq4vsaFOo08Ivs/X4t
IVtabfjLgFhWlhd8PBu7WCqITjeYfjY2wKUUQiDQ/U4TLKw1eWAN9cl+4HVxP1d/
ARzq6CFr8CRzvqdJArsWl/yTjCw5QM2ve97LwAcprl7Lwq9/0/nHxUgU5KjY3a/g
Dx1ynGcApjcMau5XLslZWLoe3nF1G2Pu7gewwP4Bq7vcsQLpg/WM+EbM0ne3hBQC
iizak4Q9MhYqNcjdbLoStEJ/7d3HRwRMQF5Z7mDNsdJ3TwvxlioM/nFRARhYypmK
d/SwhhQRnzTCYrq6OWbt4Rtj0DHnoslo5l8l0cQoaxuNmEdHxfl9lq3JmN3pgrEk
amsR4K5zKFzrOr5koc32ahROqSJh/BguWpPkfP1gEc2jAzhE7ts5kDlpQ4DW76KO
vPr98wc0pP4unebuOFLZvnHf7BdclyJEbTC5k8HBEU4MyvRb3Aedj+U8S9OgaBsK
WbUkROkJwtQFmeYsK2ze58ct0pm5r1vIf1dMzOl/4MROPBGF89Qnj8tydpNFwdYQ
QScC/aI9ap6e6Mn+0gYQtsaXkHeyvWRzaL4v/QdHpMwiSV6Jw7w4SLAn7hwPC4cd
oEvgup66lz26spv9PD/ngzCgkBmsMaTkgGsdI33fe8A41WjQzGXw+HTJmSyzxQhr
UCEAOATnkQaMWEiUvjXoC07THFsRSIcXzbVWq7s406x9SjuQQBGJ8GNNWDWmDsGA
4rM22YKtFDDiU3nQZ5eKZ0eb3kGtANWVPF8lQrUqGXW9By9teuShSEOY7+8kX1QF
GV2TyUh9KLdxctTqFomgCCOZWLBCqFYgULVVNXmovQtflmPqt4JbKulZfxRj+ZbQ
AGGyCTDa6sR0aA0CaZv9TrRwfwdJiDVgDYh2n+xNTPzG2gszSa89ZkX7VHC5tfVN
W+ckLJiTJ4wC+fBMOHPgmvhUSw67cHuhCl64q+JsjURKHG9r05nJgxBffJu571XU
Y4OWcQ1BNoG9f9jwD+SYVIa9DWMDsw9uwbI+h/Wc2Dsg9xtZ/qewgu/HhP3206Ms
h2Z/bwjYF0tRY+qCPSguY7/XByDmVRL2xKxu+6nYMjN7nJzsMbW++Db/otloXvA6
W0WxfvxyHY1z29oguL9SR8BDzluxxTjslT4wDej+5mOZZgPV692SVVsbARCNXgVk
5M52/lkOilaPqyXb1CVdjZnC+et+oQKbNrcvj5EKpwGpGREJk1EeiZuVBrmOtuC3
WlHiAmPxsSBK+asKfnUYnEIFptOOAd+WlO8p7H5AZV97gJSyDuCLVVGCzd2SFLau
/7wwDExM5kQlDTpVtXQotysUC9hW45l83ov+VKf3yvzgBxc3PO+KcXvMmZ7Q992e
MYctRvBaVWMh4+NytYwKUhW23P4MnQ5kmNSmCNMgfmx8Lev1bLAzdp/JlkE+/ZSP
HgZU8OBoEVHKH/kZe3y/V2lojI639M6nwZuEj5j+cSN+6XVSplqWGqaKVJv1Z3W0
W1WNcbS8cCBSJUs2rbvDVR8qrtS52CffSu9OrPVp7/eOMsGNkQXOCzFJuG3YJ17y
qjpYHjcEBxBfBTn6/GmS/2HknVBW2QU/9HQ5Z9N7vp3zgFR6IehwDn7FgR5Y5Fi9
qgzDEC0qUckcYatOKtjEJBNfjR5HZl9IzVtHtXaex6n0LIPi8idl/ZBTL+lGhzNp
N79RFs50+9ru/6ErDTGbkqoPgJ2w7YvYiwJifwKWqysQmMt+81JUrSBYeZaGh5+V
vFaf/ElJmr+AGqXaO2jjbiwapD1eVy1Fbafg5mP2+efo4S+9vL/wZZo8SgcGALA9
lwyXzMGcZNqByBKl9Hoi6Fcgx9MVi+4IN1+CGrToFfrEmc2+60kzeLksQXUG+5U6
CwfLcPMRmSFW0nq0mZz+iaQHaJZ1Ktcwfty4MvIDR1SAlAf1o0a2xcG956kwOYeC
rsObv6nAre6jwqIlo40RITEE0MVGXLxMST5WzQ08dmGZiVeCw9KDAS3uC49Ez6JW
MZearae8XN7LQngiv2u3cpEvWIN3OYnY2R7VnNLYXT9BIovttZ6MVmvLe2HuGhd7
6Gt9GLX6j/KZ4zA1JYibNycxwkz44aPWKzvbjzOCMVcZ1Jjqv/mVxAe+eZkjUwQ7
cdulZEorQ+feO+/rKRbWkpeWrBfG5JFNolnqgHg9Uw0sYpJua7TKO4N8PYzTdcgP
gTgnuAs54KCLT9rEbyZ02AWgA+Uj57/XU1eKlMpqLC/mkjfQ6ftHe4o7VaS9LtVc
0nQEq5D7poBUcWnicrc8NrZRzj/HltUgLpRrACb74RA4tI+GZRIvO0CGp5lpeCF+
TaZ1iJH6lHgmFU9qQvltu1IfSc8fm5b3IfSTuxJ/KhrtPFkzDWd8kP1wTJzcwbGo
fTTxo2KLr8kNC2Iyu8JQEwQjuCH/t/XU8sGk++2J2wKavBPpM4FHOs26mQVYwDhw
/CtOipJ9sU/FR9sAb6QTIgJyCfducMR//V+fKKqpX52abxJ3k1FTov8JLQZAQFJH
nUYYfCSPHoK5J1qOFn6WCX5wAKMzpvWK1oAVoRkkqOB5lyfqkOsnxmUlHcU4k3OT
KrNmMxbdpLeSwGhERKFGudqf/BW/GL0m9imJQzmw1WPqPH/lq9oR/4jCQ4ICeM73
NuXI5NRHNKUGHWdwyvfdqDMuzaQiP4kY4f99kS0xjSdGx+X3Lmxe85IgkGMm/aBc
Eri0q4Iktb7jGqlNKvraR1W+3W7iMBKKwJvDiX3z2l1Caloscqs4ZUZdwxC9jTBV
PiObaRFxvcxE6gUOmvGeEGBcNRFtQgdUh70xa7Q31rsAgkTGY/HQIQMAua1flGKb
xoCFd68lCEIycvMDW9Tqu32MSvmwD55OBjPgZ1IUC0tn/MwP1Eu+aNRFirRoVA/j
s5zXZfP/mo9ibVs4Sn/Ypo3qdYP/YT4SpbkZlYQ8bXUBz9A+rsViNncYoNs68xsz
vn2RaW+YIUQo2kjFOw0GW9FXplq/6zWYjxMV8hyawnS63a1O1X5XItKvOAdqa1n8
htrblcUTsiWUA2rcByC6mbURgvn3tMB4TEdn21w8FbwF/7c87o/yh0O9qhGlHZTC
Bgqoc1eNmJzmKAqo/sdWIwB7au8163GBjdO8cfCMGhyQ/WYErlNZvZzwcISnplwX
Ma9V7dTZi/7e9UQ71AzubxeXLfOj7RKHp93ytvqGsWCjg0iMCnychGia/AQZjYI6
Ssuu3vcEmYG7UUdN2bsxKLD21xd4DeP2uf8PfAuJSEzpVEihvKqE07lVhZvH6yyH
zki4a5Nx/ioOT3dAwS5o9r3B03HvSBEwbUDW2F1BY/l6G3zITAEaxx72PpalsYij
q9f0p453Emu/l+nmcCH0mJJSDSruK5blw30puBs46aN1rbAaUD2JlS0+pVbPRP55
I73cdA2PubtFdyjoMiQpUtsQSndSMGUsBbmriDt1IXzagbPQBkDMfYW8CAWypH8r
//XtA7yQ81CUQ7+BkwdLZV+dHLD6Fvjfz4ljOuCDVqU3dg+oG/974hutwcnDDnw9
R7+YkXJsLVKj1q801XYKaUnbOflX5gHh/lAvjTBvo3uObJj7gxA9TE4YHeuj64ts
U/Uqu1GQCRp0EneRcQZTLlwhFCEhAguUHyAUMyawJj7r1qXZFyplQvbEMsIwInjr
eX80yeV1qEaLQy/5EcgjEKE05N5Kw2gXX+gA2tOk8+gHlfsv+RZM5cOEnm1EBhRE
n6swL2kZubbbt4rpAy4xFZLStWv24I25V4zW0YS70R1K2m+ZUybZEimQsSaV9EDP
5TnkioKcJzo4iz/6+ZFBHCQe+2BDDwS4A9o5zXql/2DHbsPFuAZVgjDC9VHDXGNt
MtyIg2IGn+ydU3N7YhuI4v17EnMknSTC48+GvdSrZxrfnDgyq5s4AQdfM8gGg9Bt
ssY60Kk6DemRgiohH32GF+erJ+qN8kcHrLFlkqHo3uB7ibq/H8s9AUdKkb3h3Ykx
3l7Zpz6eACOl9/SloSvVgFVkynlgPAl9hFdSySmWu8J6ut6+gZZLq5HBr55uH0+g
XZ4XL/ujYhLfWbXm4pn+yrvQMWotRzZRAwpNKjs+aD/pOEjcrdQze+7AGC1Vlh5D
xcnDBPtduL+aVkcB+muSDcuwzBRJHazJCFH1ugZWticmw+5wO6Hb1r5/rVV4UPKr
78Yrw4BGWitD+ToMhsqqkCFLLPKO6pfdThIKnBoQRvl3EOUbZ3d7fqlJfwfBF0tI
OpDMsyNPW7ZJW1wiUErvVoUJsQHcflsFGum3l3ktZx20D0/n2jBAO+8vVM0AweNJ
KFlO3DzEuJEru2GyaSBcXcYh80P7LcaL8fRF7dXPXzP7qKTlMgz3QDUPe6d4hoDy
o08xDrK9ecF1qKR+mWXABEihbhulKMM0Vvdje748Kf/XYIElETsM26EXpgbCx51n
4HBBVrWIITsQp0n33+hqC4fzUfOiWNhMkRUhl83gGgSzIbKHjmEmRfpmauN0Vri1
qXfoGkn8dR+Dn/OD4w8u8CULbbr+z3FYLq9DrkceuImHdqNJGVZd0FrpJ7cddY3y
hJNoiFgOBiGXq+Q7RFMyx1Vw2Mg0xjQ1Yed5UCwFCe3Wh30r3Wu+XqKu71gDWG0o
4CSZlaf+8/CENE/Ly6pucvJqP1rwUk7Z/uA1ndxBZvwz+rzfvYprP/oAFH3r491I
ZbQTRFMjvt1/SghWHniIJVuEeSXPRmEMnzee6ZNG+XgWTgr6R+qQYpQ6JBnwypt8
ZXR12BATvgCvJoGmwTi4pO6T7XB9ruFIIJl91knHzOw8cXpXx1GFDq++tiVXjuiX
CglHr3UHzX+rrvq/1/ecuDcJWgNEU7a+jtSBxgdLapVc08UmB+BBYm5y5tLLA4jc
smvcxXfQYslGXHYCEAdyFK+Bpba+DJesw2GirsKRF4CfWVB2hujtkw2jNiWPEtIu
7tHv2Gcp5uVwOAl5LvJA4EtAcD+kOltGpX8zVGDEv5L0bed4a6nuDJrVMn80K7f6
jEvFE4ucOYiROKEkwrV4j/L3oDKIT0aKEnR7TNsCuqEXB94M5b1UOGC+FHBdt/42
0B8/DO1iZJKZtXHgp94MZJ8zeoLfCJ93okYNnFQh99Pj+//jRpeUxYu33T3iZpDq
Z3C6ZQhE70tloXz+dJ1bTpju75ArqEZBQIZtMMb0QI5n4QKHAYXSVTKvy/eZNokV
dT6kT5CEVlnxKmLad4XG9GzPg+ASr0GKgkJsWoRSopF89rCo20R6msD1z8esZ1tH
VFywsO0krBqGdpTJxCFp4SPluPbcM5QWiirY5E+JYWCq+sIKQfn9CBn2nmv3U4y6
ELTS5WMAYW0LcSpHYCm8WUQ3zPt/j5rvDa/07lal02Qtx5Y33Qo4hAa+47G8xdRw
l2H0sl7cMdu9aSQJDKVxuHxvnPBQ3y1sh1qj8FmrAM1lyxd5Ow5xV2/gYaeEXGEP
c74gcfmNavq5km3Ma3YSLnHYlnvqezCllc0/uAvmL7+jTVsIEDI4X+itdcTAzqke
yxnqXpfI/QB4pnyfipDFLtIHRo1yO+W8wlJVjPVtWWFXZHdhr+SjuaW0uSoDwbb+
TXJRyscyWA5SzA57AKaqacwNjCxjskq75hiXPomiL6ZsIHpr3qOFaTcq14GPAFJ8
RW5KWll43/QJNoOmaOQdIvHY3Vg1qscPP7/Y3MtG8rX3Zr/ey5g5Ke//x6ijg480
HrL2J7v38VaC/dWuSXHpFZrysmaMTwPCYK+zqvxE+YUTVqvCO4EMouXkf+clxcuF
fH9cUEo0+GU8u+sQOvmtnPweb4lVIwEPS0DqKoI6YLyKzjnG4VoRvZeAMAvmQkUY
YemfTIPEcGEBY0WWr6jUYFB3AQXOwiBaj7Bze9W1GfizX+xtwGpn7SWkrQXuSNyF
oBmd/c25DPwKz+AGRZ8SvTF3Djz14rX7BCeLqgJvx2OR0HZwKNvwALo3E0jwXtDW
5A3OmSFrhmXHSA2ocaTcXO/wyv/R0bECsZ4axfR489hiyxPVgOgAKKAvqjPTFfzu
yWpHM8MIeQ0/g7O7tgv9Hj+3XxofHvZfg57odoDnf3y2IgK3OrC6GiOWfwrq1HAu
HFgBWth2pRhdPu3kj+OkyPcY3/RgzYjmWlMcnIw7A6TJ8HY6KoKJzsfxamFGdlSe
Lg+54U8+zJy4TVmFzMYs1XR3tqmRURKvEnXHJ3j7Wij3uIAUaC9a4P6tSGNbmCWJ
/0lUJSS/DxfLm2wrmKD888W66EwBM/jbuTdQUolk+U242je8lwCUlqFTmLJ4EK3F
byHj8HcLUHZoytND2L67Pi2Fvm+uWL4K9WuUUuYck9d/dgLTgvt0iT0R0URXUZ1z
V6Fg/kYTlmSdjGedW0anned4M+3zrmPs+6fZuD2SLULSEupoHysmL8D4iJmDQVVT
dGnd9jHgTjSG+bzoT6Z55hexVYuZ3fTnO04yRV4ke3Qzin4BrIRC67LnQQKEb02c
Y9xZrdfIoJch8mFUfq1813LjlP4lJQVmcRO9CzW84JiTdhdb1bZl2mvPd++RRwtQ
In1WVUAvok0EJFf5peqDAOVH13BBqL2GSDxHAayuF7vnpnjb+2qO5bwOdAP9M8s9
Km1uTVgsKRrG1Dv4l7F++YP9cYOUNfSSe66pb1RsAO71iGXog3xy7IIFuXV1jp5y
TnpXJlzRz+Na18gQrG7aw70i2kanmpjorPQvQpX+8TmHppHttdYcl9xhtFAlNUMz
qbgaFJJFta3ISqJdn7IxQOyCqyR/p37nN9qvMt72ryxj+h8bnWB0Sfe+ESwG8D0n
2e01B9v+Z3Nlq6aIL5RRDU/yxrDj5t1K8NbVlUrYPvrD9xg2emWWygDf4mN5h//a
ftn5uxnjfKqW8Cn/e4wcuqr3GBnQyneYoZ6S5DzyL7ZL61ovVuFH71OIF3Y+ApQk
WCn4/jSOAbwaygYivNMnQDl2wSzvHQMC8wuGC4fteIPf82HqnOwGbLR4fw+33RkY
7DrfgSRQrQKcj7ZHHAZbkai6WeBBRV5jSGuVcyuMULwiJhdg2PBMHkb6p3gCW3TQ
3EOH3gx37vaoRM+LkWC2lqMN6ViJen8qUk3ef0yll1ELR33zaSDEsu0w2EcChexu
chaeUORYKFD2aOMmG9zciJGyPv7orNA+xkOTfB9ab+Y1Z+PjSlV5H+JTBTT8QKJX
YaOcA1aI+CXdzasjtoHpQds3Pkp1AVA+P8Do+/cxy94Sx1dLts5CUPBA3wCGyJpf
iDhgeJ8WHWQSxYF8Gi240F+cIOnVDkvmSj2gHDfwhsv4UwjtoyY706tEM3mA5TAs
blM0Rv4kYw6P2DMlDSFNNShEp2BIhUfp7PTH+mE1vbRIshjomU8iDib0tH3aZqv0
T55je9TZ6YtZUmfTIQ29QXTP7+7tM7TjxPXHOrW2z4peCX3fWfBZg5uBn1OHKCP4
1aEc1qD5hRXmF+KPwMbFVGyrN76jbPdFsbSpldNOUcjio7WXefp1uU7sC9FWHzSc
9Hpqpgc4yrmUVRUwIACbi2XNQoLIF6XmFGsu1Z7yVFHIU9LkXKouMXpNF62y9Kap
1AUHQ/xYBS/wdChE9RoEHRhZwqc73GQpOwC5+NrNac2jjL/lNng8QXnjJodb0FRx
XFn9sSwn2shke7NbgOO6x9bsSbeppuh7htv/D8GDoW6a30QhF6LFlKicY6472/L9
0cssJU4e7y06fQ5o69NwbYM9+KUEyP+AKz0B+AEZjBM9SVpMbzU4B9JdVweLTbIJ
06ozkKidA7b91R+AgRE3oXM7ktwg7BQe9rTozPKBap6jsSyccCXnpt5JSWy7pKwN
07z73tTkgF4mxy7sFoqNwIz9/HDiwEIzpSNdbtg6I3yayhljWi4K7DpMKlk8p0pG
UgT3TkDd/kPV6Z5TBI/X2Gf+8HqGYGCd+r58DMVLZzTLQR3ia2xBr7ApqU+o2oiy
qPu5U7qSG150t+ltc14OCE5iX65UldlYWPniYZjtiMns3mFnButntWalxmGGUmSI
2aONTJCAyXoCzZqZdhp4569hSRTmlF9a6z3yDDYUTuT2fah05jF2wLirqKvzik7j
McJPCRAgxAv0rJOTuB1SQ+Ph3jqzOhsjUiwAOIccmkmMadIKbaC2xz2Rj5WmkNfO
+6RTnkTzYgPGNUwEqnrKij/J3jGgIQGtMtwhbfrr/+V4mYHqtXHx57W3rNA6y2R1
WwHT5OOLnZKzysvESUvyakJAExlY0GD/mqI0Y0xA0XYRuuffvTgsD+KlyrKokyW5
Q9vLYbKab/+xEnpXV+NMvGptStY+fk5HwoPK4NQTDpHk70Fu2MSn5anU2hbHmv8F
UcFaV7xrTWw33+cw7CKzTcENZ3n4DnfbyP58UJMYJ4HV2e+BMHbIo7LbgU2Eksb9
cC8saT7JBqVziKaMzOzDdOJbtzCd8dZrPnQW0abUc6AMUzWwiVY4woP/Hpkuro8N
Ji+vFvHRTJFQfjlZl341pbnl+7MNEFbaT1066a9TmK027HEx4KSNZyesp5xuYTDU
y1Ok0g4d9qXEtNTThG4RFaAjm0ScJl4VYAFA9k3bvIfTEsZFu58aYB3QgS8IdlZv
u9YgQHALlu+TqLtSLMy3tCPjeTiJLAU8sgrRrvxVnu5kPnjMuoG+VyoMALDvZTzQ
F/PWDB6LYI4w9kR+elysgMJLJ3llfe27Te45No6KRM8HFs3KEEpiGsbio4rpnam2
nOZ8113GTFv7LvGTTG0Swk7PSZ/Rt1QGCTsm/lyJ9UjwrAzEGk1AjZw40yBbkiAK
Ns88pzxa1xpQj45GWqbLwseLQu7Pov9MLRFnyfVPnuok7DxtgbCkZtLrSpmcNbsh
2cMB+zVhQDe0SxjQbyicdpRZN10dFE+jyE8WblPcqRJ/AmJ3SmX5rQvpvhJgWOpa
4UaHbmqUomZ74nfiDkKI3R32TqS1Um54gnlfjYjyL5L4gP7YXhYnKHtyBUD5/55+
pZQJ6wvcwEXQAJ3s2ZI1jYZ9Lgf0gVq/G3yz9YRb5j6UUpGhylgJPCCfNiXFSwAY
Op8FRJ8LI1T9V6aiLN0Zvq7vj6cZLoD/q/zvpzmBNy+ADzhyuOMGa1q4Bx69JSQu
KCUKJJjFx3APFUqCIBt+B5EdUFNwSVEA/C/5aKu2WmTblTve9pzwPVo0+ZwAtWEH
MGQdkGhRX5a2MSTXoMquHzKv+Ffr8bAiNo5y63/JWPXB0qKhPDNRnLPXVchq9P0R
IAPPcIg663DtwOsrI4GIHkzDeLU2SkZvgs/G/o5iN5T7hV8IOb3OFalqb8ud+kFC
yun3daIhkaR/ti391qXFukEx6hYvB8ebnzshP8zBccjkRj/FYgfbVAFHCnX4xPZ9
g2vzGB/FhMsT7yTgLjT+RvBpWrhwR2osE3V9qBEo2G7DNCMXVcf0ycyqswk8d0XF
a1sEsb9KWdgD0+SUZxlHln8+MNpEW33wNQQoxLRS3Ns3pabxM9yJ4CxWFDe1b94h
ML/d/2/N4ILOPQEcfq+MgXxflVivWeveFGt8QPNJq2i7f2Sh/DLqbAc0WqzG5/AZ
qtg2CBKWYc8bRLw9v67hCXhYoCHAg9bwEFyq7miE3t35Cq909RLbICgYz5UyqsAS
h1q4zxm1evCLM2Det3MI5x0K2NTWD+ER07ISDo/oEU1UqGJhllJR6gL/olNeG0LD
P+QhMLmgSWds+DlE5B4u9YmJZywfELjMrU1R03acZbtaeVuwSL/COQP7Ziynr2Qr
y32v4LrL7Gd6fmoHM27oOQLwa7ZmQuMQ/TNjln/ugJZysrDm4OyKRHbge1sQb8Ol
FzOY+GQHVOUnX/Z6xaU9KFARsNA3d9e/AoBIgQJEqgb/ckXG4dIhmYPzIKN+zTj3
1s/8L6SCfM56Fj0iKh1eVDP5AWNTDPjwPQLxyL4HOwfNcxXScLBpQaEuq99J+agi
m4o+71DF1qYayYF/LA8elS5WKbbYyxn1Bo0kJl8AOAKLb+lxPx+0PbeHAde6A5qJ
XbKkqtOs15ZDhOnkpUVpw5Hor8TW2NMdHaMvWV+frkI2TTt8WRIFGr93DNKkmQb9
ZFSIUdlXqBxyICY3N5Y9UcXohPj7nkHT3nJ+m490mTIWTXSNM3zSc53LpFwK0CFu
w7cnfF48JpuTJYnMeWhtQkrdhXcakU+bL5M1Fwx/gYvvgwBFlpeq3nVqKvzmGZzQ
XblSR5oiy2glYA2RA33Txv29M49SzUE/67c/ZMF12KP66QgxA1F5sqLPpwUcqyBB
0uQeU2G1z8fajwY5j0BO0k7IA930dMmM0+mus9AK4MOT0GCcjsj1E/E7ipLbbwKt
EIKeorFVat3og/VU3tnlKFSePvI18RYoLtZ40OsMxAoOhVvx5WVX13b+0YBLRI8r
g1dBWf3nMr7+BRJ5lm29NTKpYFEi429Zuxi9OU5Z1o0kBpjlDWKSqKgYndpMm7qq
iZWTcYFPdrbHjp7dFa+n9niQUmxuJk4IWuz65kksS9m2s0J2wMd/EEMwPlnWeNc2
U+I4CufSM5nTqR1ZDov2AZORI5se8xwAXqoMuIz6ffafuG04L5VJEKA2q7YHbktA
Y3iPpDrxukBc5QBjnCt4Fw6cuaO6TnSd9Oj29VjWnNWYKv6q0T6xU1CW+gq3L//Q
5R4n7HGc5bhWEKwz0RE+GQA6JxRBGxKlds+xZlbHYYPaed2RM/F+zueMINGTOR2y
KnW0TerrFU/yfn1XpbsVa8P7j58LYYcTSY/UBbqbhSwT+AMe6HPh5iX4eAWqh/Qe
z2rBoC9AuNmUZCL/YK40VkfVcPBwoGHyKIbpXbqSv18kLa0hPyGgI3fImsWmSlb2
sSWnW5/pCHHVhKfdJnMA9NOg2PMa+ctZfGyjyLdoVA1mm27DsKsuxzb0xuLquQ6W
4gozWP+rjjm9uXhOxgulnSM1A6XPzWWwHki6SgfIP5OJj0tu1Z7NI+3Tta9dOJsz
YiuiW5qunG6pxvOzetzkkye9AIXFshOX0eDiqYyjDb3psbLyjtPZoc2hlwEPfbkX
KFnpjsUTrKQ/mEy9uMvsf2yp+EuKxhnKfVErcltfZUtWo564AO8X8iDjw/QqBfhl
A9HT4+6PWhuJopFBtDqhDOBArldfia+QcRtzKIATX40FBhAmufVswvZ2dqxMaguB
qlSB/9gTWeYo1S6dbq0MqKOWU7v56cMdC+6ebOlxSctg2fi+xrQGjmi+JDEVTzKt
yFajYxRfCiWIRuWr2vJbuoX6HcdTbsF9MuzGwnTHSzk3HFCSEhmZFrAz7v4DqPfU
cbQZaNkqiCiqlEZN0lyxTuboiBP+LiS6ygOwr4XI9CUV8UD1g7NXr49lOCellV0F
ZKOPUbP9TKzOBJ7QMeLP7SfAAuRllXRwa0Pc+/gkcSZIATseF8DNqLxcg7D5F2a2
0vSyehj17T654VmSIZCCwdaYtxID2WrEqj+8U1JDffTft2L+Xu05bO3NV21bWmcN
bsYefEu+tVsNBVH+tF+yNiiM/w8gkf+mSNTsrfwoh+4+03TwG8MrpDSohixbPizM
Xv8cR1tnGlW5YT09WBwijwEbykF6QBKDkpI24MyOraQF6yJGt3RzgcNovL/QL8DY
1duM3V2IyOV2tjqp5U8HYwj1lmA+TA+eyjDGuZxVIfI+QOfO6sebhzNqY4HKVi6p
I9xgBjgLJyrDlIgh7zyq6/Fxd3u9qKrqZju1tUDhu7dHCPlP6ATwa8GfX6dJd3AV
WeYhJolnEwr7wG6dOBRmuN+zurkk/odTxI0Y2ezikkekjnuhEm8KrBzzMxXHKEGD
TxyOKD6v9nGck5INyA2KDsok8fXPzjVTjHCtQdWjrK7SIK4cpSWXlTnXmNYOef9n
WzkZzXqR9EXqz1F5WCJfoTkHxR+cDvhR0FVjj66TOOlMG+Pgk9/vJ6nQsh+HCwCM
9SK6crpETJGTIAlY6IExwCLK1uQlKaRIsv65AjSrxGMJUyQ+g1AofpPMKPseAcju
6GHjRSHhBbsFd2lrJXhm1gesiLTA8z8lV+JlYMlxIbYnfLUrayJjqZoCfcH0Ik2F
QZx7vuTnqgF3JhF12HKG/Gs9nZxuog2rlLgcHGss8ocgLqpLY3e3yIUHyI0Yfowx
l93akjhXnKzv0cfEd+ydorQQ6kVxXeNBqgAJ6/EzIl0xV+K01/0nSDUSFbP5rPsF
tSdwnBJ7/71pfcwXVBE7FeR385OKBJ17JEub1hQWAhKP81fQB1+x4VLh507Zw+AO
2zQS944qzTNPCmQ/ZnBFXJttUmuqfNxpOBxIktQXlLXHMRxeglOQQZGo7nvKP6CO
H+w+YPS/qwneVUqvruEJxUU4y7/5M76Fr/wxsfPdiLkH5UCCmeYVojkzjLnySBI8
L6M35OIscoyWJ3zfd2yZUhHJSA0d9jUsEPPSrs6MrIXrlLilS5J/MpF7qpUvW3+o
kh/S58uclaCnWD6RwGVSmyBJEz1EpyzP2HgduMc3ua+SPezS83JoSeu6nUquklEt
NeWZ9g4oOtu6ymO5v2+w/fFxm3zCUIbaMSBlfD0SG8sOYJxScLRVSSbzHXAtxDoJ
7c5CT5FKloNFvIIdrLzbcBQ6dBrJ/cQYQ+2jHuUnEGFb/Gs2O41a7XtPP61drgHa
JWQOAdAtxavaSna+7dMvB/C9zf8JiDpISC9yxYDiIGVRpbT8IfO22GSePtbIy/7W
a732RMFiazr61uHyV7jXxN0G0/UOZigDtgamHDD7MZrHg8HjSlURsdZ0PpaEaKEq
Lb2iyop5ANPVzVQGESh2iZFhwaqczEMr3yeLATHE2w3qxBFpfb4aFxVDCDCINroP
AWRdktiawYCHFEcT8E5nJSR8ouCcl7U/3aoNgKvHcJvhjG8NceMfWPZiHspCCWDp
sUzkZMjlxqJ+tu1OCFfr45XXwrGhWSopbqK6K0m0q3q3j9zxNfHPqJWByagMNkZ8
eewwmRZQNOIkf6fYkBWrsZ9mcc3nQhF3zlout8fieq7kx4JBIs02W2x0/rRadl8E
tv2nIUUznZq096/UC+xCQFjkElqdnLD28/tXYi8s2znO0t/3zsusDPoXvRPimVey
NDryGQvRc/atvTnOsrm7e2np2Xp2VMoUZ/9G0jEjANFA3OZZ5C+NZ1vrWaZBuZR8
rtisCgh/ju0vxXWDKFwELp2godL2JF+zlsHrsWBY775yGtujKuqWZZFuUMOzzqn2
85zewysWIX2l9ZpphSL7AmHmGCx5wufe5vRwdCgFc1mE6GZuA+gKIkLYdCj77wZN
sb7od4i6mrjOgXpNzDsLkyXonkIaQptjLwAzv67wbftL/0PZ9ZSBVkCkqEVYjlT+
9XtqPBy7KFB1NHvWX7NTUCfieRANAiHb6Q02topXp4IhJ8IKU4mk09nTJq1CM9Zi
nzVtX74WJEf7c54kBBNZD39ZgHInIBH8cHtL8RF1GP+QF2X88HXal2kOZjIP0T5v
ABMaXiX5O+/ZHWXqvTTTtYIbdiLbzzjJiI99EvVDRuHR/mzHTWgQCfnQt6m99+8b
l9Eo4jLzMhxfj88ESRuLvXpT55uVn6YDY0yyPlDQGdRqhdPw/ExIwVtj/af9PVeD
8+kmGDABIN1rVXPlSNdSvf/9eSsvAMF6ljqUzFR/p1pVs+K8VecF3l+T/gYYI32A
EZU/urDqSF7O+N5tliJ9oxIbTAT0DNw0xDA+Bi1rwzj03iA55goc0uKioyCUiE6e
m9cAD1uUOf5XWFap0fUTezdQJhZZy0Ye5+hLzZ5KuRx5XjqtLBXFY97eLaMvE2fC
Teemf7AzPHXXkLHI5lJOG5jLiG45jeI5yGMhzeisSW6dVh6HbPukr+4WkzCWj/h+
rpeMc0Yc7sHR6xPW70FHgwCbGV/e+rrNRoiF1OHk5kBJr9nMY3M25BeHlzgah1OA
Lh9rFSdJboCqUs78/ceOQYq6YaonmCKpBEz1o9xI2kDuACIZme1jui5hVry8Q/6s
DOJf97Fti0/moJzV3gYPEy7U8fihDwQ5z2CJLTQPRDsyBgXinv6sjXsTqgR0b1fx
gJOKOF2gUeizWTil989XoKafMfM/MbjIcZ7LUFT9JORDL+sFLA5tZncydnEwtcGx
VLkNb9wPNskpepEkSaW8C0nf8xyEhgWa1xnk0RHqm3zN33qqVEvxeec7Zafs6oN3
mxT8EgYYCrfdFzKETT8keT+KJiUzdLC88SD4NMkHsrNw+qCXuAk9bdCBPluZikpI
FiA0C+SOmbXAKGc7VFv6V2H8jU2HVpWR0wLa+rwSBgnj0EWKe0TG9E/kUl6ZDFOM
MpHoutUe1UqBrorJtLYeFNm17k2T1cahF8aRGhBfefsp+Xrz5iKW8mi5m6rF2yJW
meA/LJDpna9oEXeXEC9b7e9BHQgUQbfimXsUELnHy8j/WMYfX9dVAXjqdndgc1U3
GE6F/UEXKDerlPY1rXJNUkn8HjfqoDx42K6yXZyvdnZN+uxcd3PbWuU/cHqbqyXh
1EClUyV/TvNYMRRyTMX2FTA2JkIwctYfhwd8FodJw3Euq7TCfMniMrq8rvc7rf0F
Lyt2MpSYyyNmwFXU0bf0CXkM2d1/6V45A/JxhBTzTOOSQr+8nR+Qh+WBpeoJSeVv
PMxip1/byrkwDa8DUY0RfgC5M2Avi85R5VwrUyPBz+CUxfDoH1RtwnukJ+C2ZXSR
CHCUjV8/gJuiHLfZB8CyYBUAr4E/UbAWQqlN5ppkPm0futmGekVq6mO0kERqTzwV
EmoMttEf5ZVpvyYwQUySNBcZVAdWLLofYQWhUFLLTXYtnTRHS0R8/7OmAVrcsyuJ
LY20hpklf+5wVF5y4hgaPCZLfHb/v63KUlvn+04hZnApn81dEfsJ3OSDIpRsrTwx
ZoZtYeX8zX+jMsaDPUrNWLXBhR8DVAfGaCMdbPI+ZbbXjNhUjR37ox+LmfhJ6Vkz
Fzw/HcW+313iei9gnTCRBKXp4F4WYD+T6ADnqJPsBU1KZbdvdYzIGfibKLzlpUwr
xqIvml+a4oAr0qVVQOs1w6jLqIcaQDIIDbKa59hXH/XCz8dyPts59TVSLegpT1sQ
EtKLHGRXevA7RmSUXtqWmeBysKS2+SAzXAIpZG5AYd312oY4V5Ahf3UAtCJCRzoI
fvQ9pvyCwheHfxjlNFa5n2BWuGNdC6CtX24ICO18EXP9MaLSkc5YQWoDNzcrWDz3
i7COwcf28sazCVobQB+cEnKTLb7FW0IlRdBbNyHDMDNIV3mUJjIAxQ448KPCriyS
ZbKx6vqEiVYKa15a51BxCDlRQAJTvAzyIpS82mvgqpisq3t0BfC7uTYqvIZi/bYq
SHzsMnEXjMz5u94A9zLi81p7lzSMqgFB3nDiSNkiaSO9xYkRUaC+q2+c+gm9rtmY
oRfyedlpYPLc5rhYVishOl/krHVyMPOheVGlztfre+DOGh7SeHyabydbfR78FkxJ
MBa+gRMj6zqdIlnnUTDouLpVtQh70oXmCT1S8ZKxWO78lulNn3hVM/2TF5kJn7Na
WwJfN/PSboXbuc0TGwdKLSwZxLNtoFw6+2hbRwJ+Sr2qveXe2cGAWUI5Qhjnuk1I
lBjdMdHzJ2Xy95LQQHxX96LiQHaiUUNDzES+XhrAgi19b22nLmhJDECd3vw2h0aK
hPBLM4AP8iJ2oqd03/Jyj+trIMAQ0hcnTZluVk/eQpfqz0RaqIR875Ezc5EJ2iHL
N1otnCDoO7U6yEMiXQR7f/Up9Su/8OR/sAvBPJHkUCi7BMYmCnWDJsVkqR3EgU/2
EVlNaFlUj98tFjk/at9hcUtEWGDpfSWCrefQabRc8I1YIB/lL3WQ6bu8CquZ8bYt
zRrPdWT+mvTkAbbbUHpmP7GfOOKEozc8SB3CPzRAku6xDWWWR/1ddRCpb4c3Lmmd
VewJh/w69zGHTLDtvWiYeynrI7EqCmu/VH1brZIb+Ftcq16AjMhtY0q3yLbLVB0B
1fPGW3/+mHLn7WXH9MVGkR3dcJqq6V/JFCJ1mF213MwuFk16FeWpzA90imYZvFlh
tomcFLafugLsr+G2ChmxTRaZIwY2mcCdh3IgNqlm2dtnAldAUQ5HQHvfDFl5HyWc
b0wOI1lvFXYN5QvtZQIIPJa80cU1BcbDhjarZ2b5jtaBo1RLHlKGw55HuGILXpM1
wsrbQkcv4B1Y/zzuHHHbMoCm2Kgc+JO7Rf5ywGfO8wpzVKU5GzJh/TwFAH+6Jo2g
hDkY1uvTah68pNehkOFFyXwKyr5i/lsvCT86XjSq4dbo/OQ1GbfnH76k5G26llaS
OP+TSb7UF2Q3C61Sq+hcf3x+rObukBeE9bNJMettVpOxYCSg4YIx4loZNDSwbdRc
bnMEciVjdCI1ZRvPPNvv2TH8xWrvfNYao8VlDK+X6z0/RSkzSgWMhhekkyAsedSW
LfM06jpp8wqZ81NUGjxnXqbxbtw10VER3YZDUWYy1ybpwLBtUOWXuqx3uM6TNxVU
wudYju59NyCATAEgXzMx7jklPCDNwGIPY6xbvzuk1jcuTA5ErWhIYdf/KDIqny5R
85MqiR8w6CkhOVHVtVBiIA4fsGi1x6RmFLGqgcDKIGwMyhyMzAaRJGeaI38cQhn+
5wopIeLu7t7iZf6AMe44TGkWvKbDnaeNoLPQNi16UOOy/DFj29hr2YuRBknZhrEo
9cLXmrmjotDvi4XvFzP9BoCvtM3fvkJIvExgPv2SC3vFlscQq72IpbXojU7fAUUb
nSssUSe+KhLRaKh6t39TfTB2sqLexGhTwUPcjOzcRCnuMGkTboke8Tz/TZxfBsWq
BV1leHnDsJc9eMkP2tIin/gRYR/VndxIS6BuAzM/NoIHSIMXiVxgO6qpG0xBPo9X
X7ZG1HcWNQORoC4/SSrBNkescoN0q2KzLFWZezhu4Zg+H8K/OR0OGFoBiNx13YQV
L21VrBz3Wg4SKTZKPBK17Gr691RXZtS6RlRokxkgNNPxqXBFuWAM6g/iXEAA/XnJ
qLlveQJWTwtoKslGTwfcPzdbxFcQVK49qhw4WNS5N2DKQeKmh2LW08AetkSRg+94
Z69VBP5antqoJkrp12EiL3W4RmGZ4ue3n+PApSLohxgV4OFVJQw67hocJ8BRKsGI
oxemKeEMjBFynBxl3JXF51VScyJq3Yt5xO+nY44wJxIJQfTLqcvxGVqlWp+MukU9
SAC0Di6CO1yRb4Qkm5B/ytBIyWQadfEnDwnrQbalhfc9Hx0CZmKjgGUcDoYINfly
p5RabIHMYyj7GnIyuG9zcVJRBS3HHlkQGKzVsQ9ral2xwK3/Ov68PNlj/GfgprSx
CJcCiM3iC5GacuHDhfZLcqHttqjakbqrRw7scUW8xFsgPjdvFfZsvFO989Js13EH
OKqWFavxMi/cnn9jMGhT39NUDiHQUVeICfw7XdUpKvaqQ0KAuSkX6829eWrxfGQY
xhj4FSa4Sto57/IxnEzEvqy1zqla+C8IdEQVs9U3iUilUDaPSmvp5xCNO9+2+L7g
bw4zXMuRLE9YR3KN3opy0FeTE+3/2gwJ7oesloh8eQQ6iYv94aDuNrS6S3CZb2dl
mXOJhs8uX/Pd7a662gZJfT1B9QwRPLR70viWY8H09EiRYmSBeugcHmIm8PBAvKsT
iljzAMpQriUxRF9wIl0PqjHqj1oPwVLFrBf2YO7c9Rh4x4E0/LSx/FLTCmXS47bc
mRF8CP/aGkaHT2C+IGAhDHQmRNK4H9BaKn4Eq5tMUEm8Yw5qAxJKHP/tnJUx+LA9
0hO+0DrLVShVppL0CHqfSFkOmO2tfAJCbZWHWaCsP8d3wVSyB5Vwn2hG1UaUT6AX
DQietuoFo8kVGfSinz2LwPlNnkPu3YHhOMq9/Y65aNCgsVjD5h62Ppko44fmITGY
Wivfq8z40HjCaDqGCYt+i7uv1OdM4ECoWuoZ07WzO7HJS9bTjCisyr5NFgr/0uns
6dqvtAgVqTqJ8S6vC8MSv4U/rVAkPKsGYDVrCK15MbuMOdlf3XZ8mWbW9Tzq/3K2
gazXXtOZpnkc90uJ6W6h+IAiEpofgezVNl9J4askgEK0opIbPvZWxd/im9IKOAA7
PczG4KcgSikz+Tf7EAa562A9nFbnUhM1oMTC1hj+lCQksNWUP0dTSIhvPCMKweIy
abcSj3PAx1k30wm207b4Bxi48I1w/qRdeojNkK2yo8tPLpYIomy8r+GDt22cF4wM
5C32a4p7PclZdnPXBtEJ54XPlrgiOGKMJBLkZZfPQXXYik3XJIE62OUGELiY3QlM
6smCQoFz2qbs+uUCmWv69IOJJ6e4SfD7Wq2Kk+HX2IEq8QXbxE1wuNAhLkCzXMx1
ciribD+DUbZaM7bnlkd5kCYJXQLdpuHpKPnff3CeWE4gVQf7g4t8vghkJ1LEscx3
qbcA7crtKzgrfx7GmcgdSDwJal7Dlwn6U7T5Mbg267NnnRXSW22xjyG0mDCbaegg
lQzWrfsModXo/h346IWhcoG8Yy02zvumdgS2FJ7xJHOtC2OWlT/9pH/t3qzv38QQ
bXyTdwo/dienADM4iaxJukrWJJomAXWTfzDI//bFTBZaFWDf1p0UTuOecwJHbXgu
pxKM9u+EqwF66BhUubipR2j1bYAqZIQIaIL3hmYQA8yeZylcF21/u+aF33tAXcSH
mfcYqKT3WcIkvxArO3WxCxKAfRFQ+Q/yzqPWBDQU8p7sUIejH1PoINArendxydEj
kC4wcH8XWLWq6XhxOqCtwAszMs4BuNQn/t0foXmDWsHSUx209/ARt6WV+VUXuPYl
NuTOiWaGww8ijN6bMtMb7Si5vHbzeNb7WZ2AdkD3x2DIF9AimNbM8QGpjcBuxMse
tcNUjY9pKjTmwqS4bz/tRUfu7i2dOuPnEMnX7MaXjZVsOwLP/4QZilnb39Y79vke
Gzg4qSfoAiD/gh1ehdOTJYZcFrvdx0JLvL+je9qXIGEUjGKl9e7JSXDHD0S1euWB
MCMgqnGDVrcS5uJM3cajqtTuLvMGYc91KgVyMV600ljLRINU65h7it18rc5OJ/gV
EcMM44+HKjcBNJwPeMITzj1QQX0XpKuEEIp+elyTefjiJR1Sm94LgMYyHgIudDSe
UhbKsm42a0i8geSJrhQAjGYiMezKupFxvLWMRa0l9Hx6qua9YN4ZkXL3zQbTR4PU
B7Ic0PtS+ErSggLEyN9BVKIApwuFMqHx9MFcmdNuJukZt35cV9G1pFrrDFG8TiVA
62qNO88z79qhGKrhdW501srCF8WMlXfTMC+PzBS9BKK93klE4AgbDYJO5ocfVRVv
bjwOhaR8snPhd/VPy2NwM1/+b9bsorWwJoKSXaLK1zaDbOiQabE86tr2zst/e0Yi
A6zudxk/RFMKB0kcDxAQl/1RjiiJt/KhW0z47o7vhTsh3FGhmV0L+prpu7/5hhBB
umNIsWhgoHL6KpEFLV9F1b/i7OX+Xhi8P4aKL5iVXTFwJeoGXRJVwlT4n20YNF29
G7HCVETKRyaJqWpxcIssK0Zhfz7GFX1NS/wSQpmLN5IxA/6piKcH6NqETXpvvQC2
jKKLWqLwYZwvfz5c/eXX3k0wy3GzOdF2EKcQp2hu8C/grILqfWWKxTIxg9dCSzmS
2gODD/JP3oV9ukU2PGljsj/tCkO04ynCFLN2gKIHquSvrQzPgFZn7025vF136tSt
wb6Z+PEOupvfGzyvM/jCXE3gLer2+jT+QIflHcjbH0jJ68UxcekZfnbt0rd7gFbJ
Zoz7VmYYnOk4Bj5ovbFR/+P9bTXdxzTas5OKShxwcXjQgHO6GFPVPSxGf3/+Z3Oq
nePJNvcdUU6IUOZSv+ASZoo6s3nWPW4xez3ME5yk3jBgLB9RfVEphEypY7ICPVwP
Lahw3CREbW6b2C7gTkP8c+XPbwMPOXIc+ghQqJe0oo3bg9zeZRwtncdFq/vC10qe
Y/JlS7x2CHVhaaAZdTiituVGKcyI3AXhSiG65V6qUkxmJMtr2fRZXSCB6YRpfZWR
hT92MIGl0saUPXDKw3ZxZL4rIY34gcR97KBG2CH9uqRiM6IWp7xhV6iBhrgfBTQ8
gGz77qspW88O0xzjJ8SbxRIyCXydmU3S10hJY/05fI4244OfOvGlth6BwKYbaUpA
DlMVCbGbaKlGSSR3SoIcnVqabW8/LAANKYmI99MA8f9Ly7qWgM/SoJeEurk7UivX
hIXXOdOS5mwemQl/CaVogDlcbkcSqx2NPi14i9ThZ06Nckria+tz6Amv+zoj0QwJ
cGRl4z9PO9sNIbKWzfSqtdWK//mM3lgfjx9jshZz+KWTp2jVG8ThKt1pbAJxOhli
UJsZbaGlYSC7HamRKyJs6cgAuKf9zO0j21UYtBJAQ2Rk/9iTv1/C5rREA+6fTtTH
IDxsJt3Qxo5qI+BAxdOnOeCsYQwFkzPyASMNytGq/Z73pBVnbLZ04iY+fVNrgOxp
3BH4L4XymSoOXEQUdk/RY+1uEYRAZVyiacOowHarDhEKYhmcMkhYZRcRrh54D3v0
B23K9EuH8YmMRG5coQzQcSd7s1H0SJWYwQn+khkvF7sYwf1pDTDNIOfXO0UShqTT
vHTnPTGFoBZA5rrbkxtkoN0QV7v0dlf6zxoo+aIIELJ5CSKO1RlqhwQEdb7ASEVs
e2zoHKc0YxhIKkA/2FhXKkvD3IsJQhJgBfhtf0nvHolF2z9DFBTCK/TpgJwrxPNi
WAK/1CwqXpmgnuJPLfVFQMbEDrtf8vGvU+Vkt20VFneyvRWvt+vnvlpLtNxQ3PqK
DHjsN9NLhxZpCbUMwxZxXpHGiEcuCrlTtnqfVEQCmNtsunVuIOARAFILzl3FOmPW
b3ap2wS80izT6YmGNXdM7vFWVljJwASRKmyKUE2iGnxVDO21RhlFjBjVc2BwDXw9
m75UTqaljvjChSUZ5BwNLLgvoHqUbJy4Clu4w41u5mRUnLpkkloRCGv5PcsqYjhC
fdqbDrM4EyBQuWOtGlDkZQXHGNSxw+atPZ+rNg9e1BGDTaojAaN9pW9QdPX4MAD7
Bqpgr6lercMUx0+sVQqcH4my0lQaGRszv3wk8dOwCZGqhWO4Iug2Wgu5meWIal2h
mYgpwpdITy27PWMOtdEoT7SiUOrs4AhuF7XZuAS+so1PB2W7c8e+3trSaELvVDWZ
r9MCWVrmWM4opt/z/VxYcTd1jrQ4QjKXoPq7jQhiks2/RUuTPGTRCSKLHLzpux/i
UaaMQX+gowcXa17Gjw65iNV72elPEr1drBSt5Gok5fUTx+75gZxfJD20vUUehF5J
tVGtlJoUriPVCzOjZ0PUVtgHuWlkgxhkzVgcozzzzRZlA9b2fLFSK59YNc9rPFMh
SOppqKkXxqR+dHV27p3n3U28Lqui10NTe2WkLQBCxgJsT6BMX+FK1i/5M/kWP9AL
eoPa0fK2NDUUyB+zdrevsn18PHdWre1inr3uZSljOi2uWqOMBqQBWXB0sxIM+Dfs
MeUNlhyuISitBF2V4KmCFPJMuttonDAicqFUZJk3304tvMUG8LY62I8p1+gB5wh6
SuFwJMTCDPO2aGbOOLMhar1xjdjAhcveOf4h14P1YfLvf2ZPzO8nbupd50Ca0+mM
28OCvvOs3g3+Anzw0pFwMqs1yUnm30Bjs3CvqGiyKAL0+PxPY0r0HlQj7OWwOKBq
xBgq7WC+HFtCBJoanAbNdLFgpCQFgwfldd1CRIDeb4OuU8+TgJyxAAMFgy6gQFKK
9vBQzj+11W3GMHYHdnLnBVzr3M/2RufpFqy1qccM08hsvd95tWBdAcOf1Wih49kA
KpuN4lGLraR1o7DzLFSRd3+iTOfD5MgnLkFlMegO5QJT0sQ0YnBZrv2E4xpVD8xX
KgvQL4lCsh7lZ7aNwA8IlAD96mRagyDsPFwpeUulAFXCWn9qFyJMYHHb1Zh5YGxV
v/qfaqpnSVHnYVxnFZUUJJRr+NHyPpOzrd5JBhRXipe7dUSgcJ538k7/WhsR7mjC
Dt7ez/AZ4WgCjeXMdM7D/2pvYZeN+iNkSjtnUIY7BY2jNnIQxImIHtQu1mpoAb41
Vwd9aonW9KKKqwFofHYYDD2IRZAR9GnJfGssXUkt1PTyAmDs3Jzljlzu0VAGR/Nx
NBbl4I+gjiPpCWsyA0DwPzz6xyLYshTKIM1pCoj4+0O9x8q1KlKeknz+Zau0wfEX
debzdeIS4ukr+P2wSkfBvKLl2NLPi8AVbRhEECqIazdWaWCyN2hJTI21T8Q0iv2G
PKCoATJSjLFq5g4I4eRCYGPe8dWhOi1YTKCGcPAcxQsM3YQg0mHb8E9ayxjwV3aS
+9E/4p6cvA7DE0mwTQxVe0YKRh/cBvnGfCVO2beeWll7bB814JYwo+7tBcuglz/E
HBiSCPOYXxPAtl8ST5Ibv7aePyRyvhkIEbMvtByt8Ntds62HOvP9KbIZ61yfRa7b
NDVQ7yXUJ/1FVac2uP8MVAsnQCVSmuaOR/qYMGWqyNly1KBA6BMJ89JOkQXGRe77
PNPJdoDvF9KluRgps3xABfyMQ2DMLP9zS+n5gesFekrR1+m71JolYp3TQNH4tZZP
/PhJZTe+jx+WwWx9lMeaRQh2um23Jt/kqCbQrmtwSbznKDOVXAZuXDxp1VWu8gLX
YSIwgIguJEVrFIDkwSVGDyQeTh7nSyF0jrDobpcR2DBvElXBCHHOH4qir1/qn35q
y7uqVV4oxz94AxNDnvKY4XBS4j04TieKpF6FKAj8MNUujB9SYiz3BnrDtW5TVLOx
/H59kWgIbgRfOYVguUApDNre+tF0hIcnCO4+JbNIGxT1DkUJO5mAgUGqEfDzhCRR
JypMp08hDbS+IB5wTMtM19Gub6l8mv7oP1lkzF2gb1733LNT3/f8INQA77vKljZ9
cuyrgfgiC58EmSupqcNoSYwDU9zHmXc9rJ3KEE0+w2EBTP8OdYzINMTlEsidYr9R
eW97NIoO/26R9vJXa5VuCxzeXLzQQ+3WSAJd2WMcIsC1oqKRb2f9uLpFXfmNYt9U
yVKy0oSQJboxoMjffZNHA95lus/uIOf96zp+/guJOw3KV2fgvE4Q8Rm4A5sEjGa0
7Tuj0I+g1KBgfycYVe9mdu6UryGlE0dEoBUutFljqzewZt4N6HjhEyiqZRDvuC71
RjI1BSXLwymtjn4q57VluJ4rTLsdpWIRNH/kfGoGxvb/RFNTsNWZeTStpBv9Xq9j
0tb7wi216GLMoa/QHfPQO6NcNMbqaLSlI/vtvuN9uDNmLevZzL7FWY+a0gthDPaw
gtj6NogigX75uez3bGVXUaVBf2gAnK7ARw1y47dTCG8B+Re+Ej4LSRLiDEVi+DWp
gl/eCvF2MoV32apdyRuo1naDzbhxxuyBrZACSB/U3E23iB6qgagP3nwBwB2tYC9f
1bO9DXMovkCbX1uaQK6ASHLEa010hRdGTWTocq0BPRGKOH2FG0fdHhq4TjzCD7J+
1ldb8fxuLaajA3teRYyOGqDkFEYpL1L2Tvq+Ogml35Kekn9qOt5683R3tWf3WJPg
hIu5tQrZ6IVNNFmuE1XlbHI+SjRXWKPVfG2tYXx/pIytrbYxgBGUUYhot2GFI2xH
JnGVrZVlbUVqIAVz0OsG+GnwkeLeD9QpEoO9xO8RLqjiUSoeSFXTO1mznmBVjXfP
lDss+8JO6AzFhB16/FYula1cBXHZmugAxH+r+xjaIBPhk+N6OyfUyJ2kjNLjm6jA
YnXTjdHakXvSgyucurOXhqpDpRCukLI4JlVMb0r7IdTICEV47VSsIWockXQBafIx
f0mafrSSmfaESxQ0IC9QPKNzSrf7idzWDINAFTea06N7iRnRaBBqHBIYaF3jaVkR
KcgAs/bAH4VUavZT1rVxE4EanSoxWtegoj0pgqs82JQruPevU88qaU7t+QP8vvXa
gNR3/4K/ja/Wb1jjDdDDaDwqYoVwpb8qzpPbs7KmV7Uceg0vHIkJ23zYSEAuXX7r
x78TVSD4TxIaaQDr74taKkg3nRp9ruc4QC90uwC/7COFn5wZmRCsPOKFzuY3JbVr
luVPowT9qavqUT1vectyRcMJWqzF6zlVKtGPlxeGJAB5x7q8P00YvjypbzJBQ+rr
k1Ao1w0eHBvuyd/IJTlKdJGZVAAHHueXReaBJsVzZvL7TS9Cm9B7e7ViR1oprpiv
Jpyi7tjNXP45xf6nRrU2MrQkAfGKYsnZ5w+T77uz/9+jfysRCpOJMfJiiUnOcQsa
XakfmyLpwrH0iiDn1UdPMq9H0xNHiQ/58Ggr5lHpNlbCOrDKreGmM7BwFxYUL+oq
c2C/F7lKgnyAcZ/DHOXrd57ohjPjIvUwSZtxOxODlbGl6gzdf2fIyqtA1NOR/8tq
8y1wCHcBThViWQgZVHNbz2J2EWLHtr6P0uzoinpke5pb3TjDbQnWt5XRaHM2LQSi
Ud/q8BO32Z5Ihc8LOj3YHjWzbDe3ahHFa7mqmcnAGJ2RN8jwNygDqDVZ7JZZU9KX
h4agK4vzaFUJXj3EbugunlBx2PxDCXchhxC0VYQVJ/+WfqO3wky3AkJWjCDMGkOk
vEJjnsu4J2Rb06FC8SgYER7e9MDEEQpUGWJlvzlUKj1wHloPF62SUfJywfPlxerJ
mI7FVyTIjpuuSNke/a++yI8nHzk16UULXmabD0qGB2yb4d1XZEfV2TGir/T57U5v
v30uMeYt0OlgJIg0r9iXH1z3ApbwIOjbE8I/BIkpgdMcmcpbbuMp6i9YkHupF7uu
p6bu2QjYBrFLJH1A/WB1wZV6uIYmFwD8U602ougWZ/nByEQAeF/IbqTGcM7e+utp
1htVjmwARhU0NuNtg5f3vuYpwbUfUzNVwqotgU8MdKS3deRVqqpo7Oj9TjuODyYq
YF1jIAimQn4cdSMLT8WkLH8Aoc7oIXWOnt3G0rMJNqEWT+inHCW0dCR1ccAUWuKQ
W4h++lvancPPvA0nAwuuTVhamcbKBYkT/7t45VM1EXi7fTjZADKtz1MAIHKiar5t
Q+8UbruAY4i0TFk1SGVRi6IJ18kcYkYRs9PHuLgA9eOu9iw92JizLEpFGYNrPyhK
BDVGmrV9VgGfNBjDILpTlVPd5RSb1m7I4BYAM1ES/IOmqsPTqr2p+c7Bjg80379r
CXy5JQxXl4yckcq9lY1MWjk+2qHdjFQyx6mutmGkpOKB9379fYK0qkrVutumOlXu
S5/CXEZYcGBCRuEas/KGUvjmBB9mAP1UVkIA/K1cp3SD+qInNMTAH3jlZnY1tnL0
yI46ih2pw/IJeT8IipCxZZgsj1hT/4ArnLBF6l5g9itBuuhocYvDDN32B9hD26BG
dBkGtsiPFenjBdk5tKSHbsfl5vzCL8NdOrVe5Ikv437y0VmwSF3WCpVCQwcTRpqm
IXaGYJG4kGxxnWZ0Fi9qiFwgIFn0zBfqjbLxNk7SzNyxDSfRjMro1dBEHMvWBzUo
lB4cpse8OIC+aHay51IXJ6s0SBCbYUEaxp/SnjFC2gVhQdIg03gJLniQuTeRel13
GUVIh3IGSATx3xUbW/8QYdjGBiWERrMjf8OSgNeFfxfeUuSvk1W7HqejSG93YUsp
lM3MtJBpyFDr57+I1P8yIV3xMXbGaN91r7mNhdmrYbBznrX6rE1Cv3eJjyMZ/fXB
90Xi2Kh7I/VtK0ZjadtfUZbDzlgTUr+uXwPQr6a0wnCEcjpqgv5QOHJWX8WyntDQ
vmZ9EaWswaJPU3jeOYdYpt6gLJOzpRHuZihWHfwGpvhIPe9Xg1AX31PnGUDJAgwa
6YuldM/jf7Sppv7kZQBgGkCOlfZVCy8h5TY4u2UkfjZPbvT8K90Z2Q10Iei2idf/
9NFXkNljIaZcj1ANhAD3t+eIlQL9+DMpYDJqLWaLPwomVX9YPMb9VJucCvbww2wl
j993ILAgGwo48QREfQ3a8GiQ3h+P9kjCH7++FRdn+OhweVzb8gHk+AG7Irnr7nYW
2GCDrdvYYGYgRYCi109N7aZL/IRm9n7TE5nAsUd27BIYkSWe/741CLp3CLdEJTHP
RgxBFAersjP/CNtTGnL4nO5JCg1DuD/iwtPzQDHg9DfR+Gn1GL7IpWnjS6hieH/k
I+RF+dTX8R/8trMY2lxLr9R9+5tS9624VgDqzJ84uhb2hulKnZHzikcMSOZpGYxw
v0ZpW8VdJ25MlNOKTWStPYi1tisfRC8cnH9g6/UDakB3tN//A7KrM7ivVUOXdAz/
j+7CTVTaQYtTiupzNFlviOpdeN1t5b9bM77qUPeqgIm5bJxviDC7Y3iZ6pvFSdRl
eUAmGyn4mI7UvJvCEJIFL60oj59E+vfzu9Lt0epaYpsRmvxMazZJjuvxjhJFKsgG
Y/phZ5nGyuux+ppRjt9xbmGc8cCg07gU0n/wC1dQDL+6lk7frsHhe0MP5Fr/V0aT
uMtgZ57EN2a+/Mz/A/gxUCVzjy2mxo+E1rNz59eY98V0sb9wmIDvbMTAdJ5ZdPKs
lkslv40Iw/tIa8G5ySXqac2n6ro1F5tED2p6nsVY1g25yQjxMc/Z4adOEDg4nGDh
FZ4lCKdarzSCKWp6wRgeXXDB/pBqa+1RFJX+/E6YDJw1JlMWdofKseaAP1QAyJt+
zUwa1o404DD18UagRKKgisRVYcCYQyBUlVbuhpvItBYsKoXVLndn6i3PeC+zp3PP
KQ6Yl/EGEGWocuHt6QgDtkPelVv5kuolbYJ1GXrkJo2+M4jk+t1bG8SUqEw2C+Q1
CmsG9c95oNQp3KWOudy3goOrq7ALt1IZVohgUfqh04Nq9Ukr1C+zIh8Erz6w2oQl
rl5eNG0QSRu03wyaSbb2evSOvrhqFT+8iLKO9CvR21wcbhOlSQsUiV0xYE91Ykk6
kWeuldGLf/m35DT7HlO8H724DI040GmLQDbDXmlN/IdLhAMv72Y8R1Kps2GWIAmr
5qbmOqHjehz0sIOphd7pu6MfzGzGicY6oi9Ikg1wgyFn+oEGQruc7jGtT8vMWc10
iYLY7K5KiVah2K0XRRGBjSWP6TDoreyf5rDIUhbVL+GhznQhupSs8d5EiBbOUQuY
EOsXTVLS/SSFB9Xt30kkbmbqsV6yKFXYXceiwgyaU3z4sJkf1uqYIVJtrm21YC0Z
1q0WNJdxAA36cBGAvS9141O93CmXhaK10fbb5C4n14C7DnKQ56KRCR8rnMgkuBDS
pzdppOEOVg766iaZqWjH6OCiprK4UCbZJtcP+EJiFQ11Gqneyk6nR9FXrXf/xK7U
f7eNb5PiXNayixKeKKss88U7AV45vqaaYGKwHJEMQhubVNlgT4WDANBjQoqrBt12
M/6eexge/TecBCFBckWnT5ytUqrSst0c/HZJ0/7eaHfg2lfg3EjWYc4o7tcXX+Cl
Yey9dKH2as5b+Lj2Ljy77Uw9s8aXQj0D/YQiB+F9KAmkjm+Gl9D08bBaWaGczgJ+
Ai6t8llfXqpVb0QeU2SjbF5j39L9AtYSPG1GpaUK2V0gT0OGLHInyp+V8/q+wCrK
FIpCfz0WtzRcQl3QaNQ2Ql8f2c1mRRQr/f3yqrg+GbNWAIUW1SV4u0ds0Bd8To6t
EIG74CNWTskE/YaHyDKSn2uy0380+1wcE3g5KBSPwg2uFQUExouZ2V05hw60fKlI
qmnsea8mZNSk/h/BFVKAeblAL0aIZH41sakZ5kj+YQ4mstW0RXnbyjFGB/hXsJd/
q2FasYHsGUq0teXow9y8OM8AU2ZcC8nmAgeOEzZOZCu8DOTqMOaQoF2Bm0p/nmYj
33b+vfEZe+bWDXV1yO05i8EFynQWhyjRDWpM51t8V38qrKNPVJIQehX5PQwP2+cc
Lyjc0mRlJDyCYW5NQJLlVmSXREsk+MCcLTNa5Wb5JZD28Xr8XWSldaPGVjGfGrbB
LsZpYeCfz6YSLDcJxsH4ZZaDqFypmFAsggqLaUq+sa03euXEEClrAwSM2CREx8w2
byRcN04p7ju+BSc9LTlGdB8Ns9AuAu+w9sidpYhsejQ50A1yqvFpFCuLkA9SHq7R
zagFvzAwsa0rEC1d9iWJ8fe27OqXgzMB4UkMWFKt6/rYrfxZlj4M497vzkG+dtCs
CpwmCFpi/awSe9eeBn/LtkfwXJL+pVj52v5KGjE6nn7WDuoXU9pFf8yEiof5e2Df
jOYJfq9sk6VPH0aW0nNuj3gmaFPuHqrfKWbU8h69uWVj9JJksBGnlJ8ixSStuAiO
fRSOrQM4ni+9rvVaI6Aql7PfN4rq4X4fqWXvLdipnqAaf243lF5AvkZ0Ey5NDwib
2VDfsl9R2upvrtZb9mSPtDhZi75OUK+bEaPhmAOcrG70UF1QE6AFVgVQAp+6emhx
lBtzEoD0TbvrOvcxXKs/SWjsLtabpJiSOaTzh2rUTCUc915QhfSvylBqCxBy6PxR
25RWvJo3irz69GtI2rvWTKH1Fc4bLN96c/pMr5EGiIijcWNn2DoraMn6kMLYSEPg
U+8is1saxsfbNMPrnTGTljvylIkRP04eSdQgTSEMu8a1F1ArFKJGqLijHo1wKR5l
Qbx6dXBUX5hTEkGEmsJI9rePDupNbG9grkD7oZ2VDZHVMF3TLtcfP1QYS+5Va10k
acq2mbVsNTGhO9HXmI66qUSZFC4prTO9y1Y6yPP27hF2R9kG5pH0dyogG/tLuxDa
WW3qmQLFU/yngGInMN9heFj4+GtZlf4MqtwqwUtSnd17DuaoTb3hOUEBwPb91IjD
fJDJlHaeX2G8uA2QZlhl6z2YL7phcY5GLvBCBDli03oYB0rltIAtA//hVBAiGgnA
KaT6ZajZoWx73mp5g74SP0rzzWpZVK86qKSx4eLie3ewaBomfqJsUZD/CZOFbCkx
5/1cJT/J+UAo3bLe8XhMe1r50dVCTjInPf7xvAVhDzL2HVMtzjqqXsB4HctymdmD
ISDtZOdu/nI8+S2rOUymZSS44Fn2aT89dltaozUGABYlFqdeDFm+OH5alIB7bXjh
83n3ANqMuYB3tDNNt2CaQyIwsxrZ/ZHf7LiRKn4DdmGRtuh2hbgPvz3mdrB+7A73
Li1v43znImQkNyVZFxtz7ZEDBWiEDYZTPfbfZlqALHqkTvqfE4LQHRgF30ktRrvP
HAvZ0l395h7DyugYLZz37p8VbVOYNFeYOFRBAmDKoqO1NTwhAhHI19Rh6xjIYqcW
JtYhic3s4XG8pXroK1vJ3mS6YNu9X1fcXAY4TNRopXOmK5QWujzj6p7H9aYazdiC
tamE3fqCj0wbfPaBeXh5y8jsU3BR3SUS91kIIAXh7fK7mrx6PBm4zxyv6Le6hhMT
cODfjhHIw3UNIXcg5ZYmDC+cUlbXozhiIJ5qZPEMLPzBMZWIBE4QAWNyrAfJbplq
eojbPqgNUy25srzFJASuAkZV0SpLM8yfljPHpNV9aNIr7RHjoA5psiPVJ5cgbzQG
Wc08hcDxPmgUCGIMQd0Yo+x1loUIzY2V5gno5DMAEXjFulnuchgw/NS8pXZwH8xw
19dfhkRtKTpdljjoDCtV7aeJTKfL5k/deFvyb13HtpIKJ7AS/8Iw3dvsNWYAxKuO
UVN2WkTZXQ/WtMij5+SFQ16Bzhr2vVMrRklYXcqoUOPbBPRB2VhbzQX5q5A+P1MU
JlqOGi8MR9y2plKuBPkpWBdYvKLz3lPzlmc5zuO2y27/WK5cZEucoLJKeCv2AJkL
qioy9v0aPxzSHHHY2cfUB9bblJ8As5IwftXpTDuxtf0TF0s441jh1XeFVfqHzr+C
Dsc0iD/HTNLCt9ILzXfuLT/DfhhLscQZMQ5GMrfQYz6A2gLhfUJS6oZgbSwNEBIn
8u6DtrpDTwc/fpm1CnXWefw58LUdpU9U93w9LXcfa6mAUo3Qoyqh8d78gqf9vzVu
14VCA8BpVQCmVGq3lAL2ZrwM5VnULmwk4SwutbFEUrYfnKvIOow1LsLQuvzQ8VpQ
IoTqlrtU+QJgl5ReFSQObBIGCdKb173Oaxz86T2btIfxn6lPdcHv8m3YZ3BATpve
RpLVGVcrVzq283UokWSfjUxi3/s5ODlISkzGK8vvRfw4CV6NX8puelDJMGNJclKG
5UQwgI7/pajKEzuStrWmPdQBsuONjPCVgK6P7llLQKvZf6dBEjsRhTxy8wHhyfIv
18T+ufvIrf2uIKLXaILsN7UQVaRu4zEls2dP74EI4SrGPLTqENXRX5QkZgzOzHFs
w29iCu0WWCkz9Ia5MQeLb6OmRHT2fjmhe7/zhcJiWKj2YzTrrM5/ktGHcTXXj5eV
a8HPOT0T3nvcPMvk0lNMRtUFticXOE3ypeAYAn3htRpaPfwhomyItTjuz33/HTlp
cXRjMgKGZ9QumduBRk+i1KEyy0Us6Zy+VgNDryZE491FjVY7vbVblA+jvEUaICCL
PM5GVUB8VP8UFkcYqLtpcgJJUFzQbo21u0yI2jrFwRu2PzSehHvrxXs+pSOgA2ig
fJD1ruIS6WoK5kKV5ZhJxPUptU4GT5AWzSi137E0WMdFLt7i+G4fBoE2E77dj4an
A5+sGQ5Dm0QLH6UnxcLhNq8aL8E/VVXFWks2Gv+b66SU1+p9f8VrkPMOK1mVwqFF
129Y+Wh82ScYnPAhvZEOuenHwyuUuJpYaWn1LUEg1BCY8uQbaI51cDAtId9xAiR+
LqbRFRPU9V+LiyEWtp3iEiAKLnRHnHHWNmAU3E6S/qlG+SGm09A9ToqoVARYqdJb
Bq3fkaGLf7YhLpuvdsLJa6fW1Po3Up2pkqJcr+MgonOCu2HCImf6wPKmySEHnkSE
i9sOP7u2CAzpM/eXA9rki5rGXURm7gq9AUIsezL43hbLv0eSitIntG4r+QDnRUb9
0FgsNQxV/xtY3219M412SKzBg7cgBMaWVI31+EJBzdaE3wXBQYyevLkPN2tAkZCi
4TBneqso5ZC8kPOlwDbSEeVCRCasK9jgOOpwHZh1iTHA46sY/Tsofs9fhoG7TnLm
w83bQylwgd7pHYNU1gm8wZmNVzgQHLv8ZuL50VwTM6ufSgw3gUY/EDaFeIO4e76U
3ra3jOybH7laK2h/Op7pz/U09OxNv+tTbqKM/D6Wz7t2Aij685z9XQpPGVxUZGlW
4Pwrt5LyHuiDWKDUUITnIKchy7LQ5uR3tDk2NkFWUkkiU5+gagsGpeSmaHbERwEX
sfY1l9p7rtKjvzctyNk4bKP+5oI8s3KnbVANvAM5KOADtXixWkfNVqGwHrz3Vy1l
8nZURA0ojq/24EuwM3OABQA/FDJzYrJnpEvcBQdbV6L0k/Va5c4773QnGaXpIZiu
eeDU3KOVKeOm5K9NL2nSD0wpAXIbkogxOhb6CXAff26zY4vLmcyk/oVFN0QAJ1A2
WfVzhbIvll4PY5T8KMnClKx0y6GXstBBBtqfSm7M3RPFxD2hhBAZ8g7pqAsnFpXz
PS6PN4stRqyLngPKBWvvuOmerbCCfLkZra4VTKRTSs4S0BLfjBMQp0yCbN1x1LAg
hGh4RzKdiHPofASRgfWMBUdklIjQEMEqhY4WS88/90EFygzHfbbq3xhfGVAI8dRI
MqZWc3ivBFoXeDmbvhtlGA1b3qAvqu7dFBuOb2LGyTffowBfurc729hJlq1KOZTB
FpczIgMtNHICxHHjXcHyVoUIsltajsWYHH/P/kiWpik57r6WPu4DYz3ruDxmVmBg
DzO2JC3WgNOrLPIc7nhH0/l+TF+IWw3q3j9bQ99wINA/FrL2270U7Lz2FnpKVz1H
Vp+GVZzZ9D1I4+zsuAH6+Puko3bKIKTfoXV0n3f3ev7kfjIDcVLtpNRIwDQjwjSe
d4F4LM7KYoHkkE31WlZhpjFWJGMU3hICgNRg0TO4msweSIdZ/3X9PMaGVIe3O79X
hsQl+qcLVrmR6860byqTxfradvnB6kOiRwEhqvtyFe+dVZWLXY5SXBY9y01PSqUs
1E9iIjfxFM1YOVk8eVgIuu8h53IxwafmZfcRg1oTiHBpm5Raedvev6d4Arv/7lFG
M40Wk765wUbXKcTleNxB24o4fPUiDHtd2skNZrbmpoVYNqswBfrCFm5blf1K8I3m
JDgDbPYmoJuFMw42YmLXDtG1S8cVtTwKISMFGPfNJfTxCuhZBQi1tzb42oA58tml
N7i02N4qOZ99G7/qH4qMUiKeeFcIQDQQm49J3phlCbB2+/8c8zjg+BnBI2/Iq2jn
E/SFdbBneXkdtl8FVQbl6DWecPXN/dDaON+SJnTpWx2fOLZb2OyFuUln4zVM1zBQ
m4onUegZiHGzZEexkNXfj+ugyTBYAPeJ7NIX7+0m4QHGKjc9d8O7Ys3fitzYGLeW
eXgrQiliM2DW+4dZDTmzp7nM1NoAEi2Jgho+VTvNmnuVd0jON+TjDzY8228IiHaR
VDDpghbHef6po8sroi7MpHRva5k0Ac7XGico6JZJXId06IYE35//b58JwQqTOe0h
mv7M4s7M91ut8ziRi0paDlznMmESY3xoIEF09qLOUNDALYja53ePMz+45bTK89Xm
E9hOTT7UOxn1eKiQalmgns5MtWVHDkcNBbA6tc/HbKDgt1hxkrNNr+exAkGFOXAy
m5nt6n28xnPd9Y8BKg2ZVeVOp8CFB3Ez/ir04HMEPw8Mt9wBaoYRK5gwhTT/uX+B
aW9arrIpYfuqhc6PdUCSfwi35782UIZl6vH8rEScj1OV0rnhwAmtkw44AlCmKqe/
sUScmjSSyj6gAyd01iw/taD478CV50RIf7bvtsz69LSubqtWogmUwCOr31L3O54z
RIl1tgVBNCXcYexgCo2HsoAOHeAE8dBeOdu+wB98px/+f4Mx6+57C9JneThPwqa+
M8RXbXw6DzjGTUMVpPAgfgjvYB5cfUYBU2Vp22GicbLjU+3t5MvQ1lPse0PZAEnf
3GsQ2QWk0mRh1bK8VF/NbzdWtifBk2NS7bhgUsWkzsH4AuQmIeK/R1mfV6QKi7bL
he6sx90pF8zbXXRbbmjhFzsN/cKHxyh6PvdSOpRVdF2jjOpSSh/msOeJa/1ebjs6
v+NrEeKwaRDFt1dVx6AZkT0TG4O1i1r5CT3YroLLYiG3KO0pZbRJopR244GtoWnK
q5wbMaICVuHQMxqYbM7LbgHJZRy0CVWf0yWqhTD2rhWJYvR+tHqkG5J4m+53Wm2E
lSthqDnW55iwJ3A/H7XG4fZRNc5fiZi7WXqiefK+ByS/hH68aOis1w6FzY+pgpHV
z8uLL+IQZ2Ser3fJSDU6eBR0cv3WwZfTjUpNCIxex5UfSFAbTkIB9V4OSzvSw7Al
b6sdC5VRT6x6Dm9Kog1nO0VQAl1LUO5mFXwV9TycMCQnKRfWjTQOBh/Ckt0VzKDZ
rXTe0WM3rj2UAJIYKJz45xckeZeC+7Ns72bL5keVVkELkAE6jDeDARyng5FpZL1z
mC9+TK77SsdAC8XCGKu7qrIQYEGBMLGPoVeIfIQGY3ZPncaTJi6/VSv9yA7M2HCh
O3dqry3AEcKTm3nzztdw1ypbUC+zM3DSmKAZMEnNBqDBWyHVQeVqtQoVbzbj1Pe/
2rcdRNkvg8+ZK4iDMpvgam+2JChV1P5CHGmj3kCM2g3KmTOOjx+FGSmmfxCBp4SO
SW57Afk8lZx1uSTEQkKV8rGiIGd09WBBwgh7p83gkeiGHs8TZOCH849VDvswPUiv
40udyW+PO8CljDvxhCTAK7VmlXgRFpmMD3tuw3RIsTReDnZ2gyx0TA0Hs++kLMdz
bYKPerGiM28ir5W5+UURKJH5OuWswKAvAem2LRvXcKMpdkv+Tm3udZDAdlYLmhd3
6qVBQGy6saECuCjO3g1j29bWwAn+iRApmD/kHkn6dA2pZTEsQiA4zasQ4Q/IqAk5
lxu68B1d/O5ENqBXnVGmRZXCU47fmCMK6rrSwRJG7hUbPELBangMRiO6Q44VhR2u
qaK8v19081m23kn4wW5kgy7m36ZezaN2XPve4n7kVFwIhEUPqk5AwrRrmrOQmLIL
0OmHAibOCt+sTtxQMPt9AzRl54xyD3E4gWTMdQdxwn334ci8rZGVFRP7Br91Moht
GUfINRrwookg+7loMR2iJwup0AGWcPZuHaLwembzE/eDIO97CtaDZszx+kEu8Oe8
JMk7PvaKCA423dI5gSgUNPLrfLa6Dc8eD3XNBIv4xBnqQamu2mluvwaw5lmwvpIK
AG5wHxuGt9dqlVautGe+qwIxmqPhgvP0p0p8/fJqbaAWf5+XPnw/JJ1R5Tfg7oxy
8O6y6HJ7pr9njBRyfN+tAtARkmE3CGgzB2Gf6SNgOdtScgaawOg4JKnJCQCpWzvK
2nI3jepprRNbPSThLqNCST6+UtPGtMROGTLYlTGavVb7AirT2nTGQXQZAOSwAV8q
zyXcw3NzqamuYdZ2pMSbzEndeRCz3Iu0mO3I4LonZzpgITMX/PEJQgTmzI3JZYGG
A3KhINRBYJG9RlXGMAo4w4eaIlqBn7bBD3zUsTcd+7SqLDTbdFZ/aopopLTDTLkx
UTrPvV6aJfPOxG0Qke7hAQiJiDaQTZfCuM6lblTbf0+yBfinlh6fipMeeRuSwl9R
nAI91BdftVCQVU4tHHWgKURUMPUiEUuE7+NV7BwF+wiO0hVLRL3AMbA/gfbL4doF
GBHxSsJY4txN1KUoOKURUciM0nv2WgBmFR5Bd4iI7TY7aOd7O1uc5yy+/vIO9gKV
C4Nezoc1p4Fj2fsdwsAhzeCpMy/qFzi4W+B6LKFiTyBioFFtAIS4Zyz8lhXZPW64
1p6XxSMq8pzaGfS8ZQXW+JCQeDcvj7INd8UglMcPZ+IwvddeDd2fz2o4mvZ3fFAM
dyUni9FAuc9FlcoXiSbl8vyOzov/a5Qe35ZgWlvGKqy76uaA1kF30ROhem8zDK+2
gjTI2hv3a3Zvm4xTZK8oxGOZewTwgxG4UYo0NE1NFTx3Ip0xV6Hr4DRZdy6RR0M6
svSIu8Q4U4RHTChfH2PeMD88QMQNL/hSu/SByiB0vZ95AsLyP6ZUJt8PtfULjRJs
1CTlCeRKHl9lx7zC03lScshughL6WhPGpsHR2d/s1/ex5BWM0D1SxZskeAZGZRiC
jruiCJlFBzLZPujGLeKzG0FBZ+AI9l0F177wtNynh7eTW/zgc6feduLMLawoq5Ln
zUcDzbk2Dl5zFSGnnnpl8iIaRkE4IYAKc9nQg5AuKMm+UQM55FsQ8jd9gmPCh3qK
6N9JWUJCJGlfC16Q6h0iD0j5OGZMpmwrA7bSTqxj/PposD3BP4pY5t3IA1X4YG2z
yvYhJjT91Q06BhNN2ZfUwbc2lXioL8dbJ+YWVErnF+JfbwKaLHJ3bbaLjCUDUDNG
BkjA6BVqzJqOO3uBONRIP4pYQk++XGEqMGBQbQT1ayrC3C2DTGR90a+3kVryg1qN
irM/pLzh9SFMEZsTjyOmfPO04nxfS1WZhKb3yTWVewVcZJ4getWnuFkXLm6IXUMg
qh1jNCQLh53OKEkJsOFl4WdYX/NO95iu9nvQBHzvxntOXpr5XfqRg9/qdIWDnZlA
DQs2cL8ta7FEjgKZ1WsQvALXJ35BBZm9/xLtE6JT7eqVxFJ9BvLXY7wavs5kZf+D
GjifDCri7mplIRS2Ed4chmDwmKSRuwJvuppOUJjkzNy0O0Bl1uFBQl6GxMZn5gBZ
VLPZsku0QZ44RhNn+ddyOgcieCM+243rOWeS0EipGoh0lHOIAzYya/Y7zEe1yAXw
btLy2I7/qmOyKbDWWqV12jAFc5t57EjfSnn5IBDLmi6jRhNDNSIYTWGJp0NEfMHJ
jsbmDAv9rDyRwCfrFxzKPWRuDysGzHZUDj4CUPAlz7PuWQaPMN2GMuKjEdodYLyz
6dj3V6qnxHyMhp9Vu5gzwso1UhGq0xhmWAKyTRJ0V+f8ZRVGbkuBVRN2LT7IVB+D
PFMCvrudhpv9ri3AFWj/9OrCJy9YpjDRktDlhRb3doaoDTRRytPCv3XgKgrUuluV
4llXv5YbC4hte3zQyZ1mP7pTmQ8jQbs1D42Qlo2iULVxCL862GcWatgi65WubvRR
p26OhUf2LVRHl7r1IfhAY1CAWIh3EFD6Y8Iz1+h0vIB999PcXu3aJqN4y4E56Oru
aeSuXkaFd3HOpqpW1TAysDElq5WvkSFic02zI3SjIKvE4iey1vsJ9vH2V/UwChfW
bxHuWlTSqItGNZAnsD1cOOHl2iAyb0sTQLdpOIN1zc7b3z/KurrDNFV9M96+IlwM
isIGVyMf79O4Fj2/1ltQbbHFTD7miL8LeqONqfKZUdI4HsSOowANuF46EkQSe5iH
86rOiWxWwQZ6UupXnhpYuKrLzUktXXN5VvreG2sZQ01CD8F4vBuEc/I81nr9w8tX
Km+/5ua9xA3d9YErEeyZdW53uCzTtUulAbDDnIhowEAAzO041nLCf4uaV2mQdHRU
vDlc/X0Lv0HqjonTpN/IvDSsnMMYjqZWh11aA0CTFBr0QsK74XWqi1eQdcV3zawe
RDkRObFWoeb7btLaMZVHJF1xobOoBtrD+7h2XO42NvQiaQv7qftsiIu3WMAYyZ3b
cxiCH/16KB++0zaNGBMTshuLqm62N71PPxYCwDSnHwg9M5TCUt+jS1B+0vFIBY/2
loz/eEjYOT77Xn1H/Z6+iRIxrUVKqjwAjaid70koXQLGCoy86lyrRlTEYfXyUhnl
UAdxmbHhukCjyCiXoMiShtU+exS3xv2fzE1YKPyhx6FdwA0WTsZisR2qWmCTDfOj
w/1DMb00NKCnc3IYp1F5V9AjYWbE9RjJXluXm67bhlqzNKrMZYNZ41zWO+iaaO6s
zWyDlSNOZEfQ1ucqK+vefauXjeAZoU9r2N4/phnSDUjuItjZVEbL7th5Ftcx8Vw8
PrJ0tEOLstuzUXgarXthUcf3IB6Ojk2XiiFtJhV3qhu31DvhKiIlIRGmGZx/S8hh
YK7kThuorrn1Z4akvMmAuNo7Aa9uuMOLsM8EbUZ0+81AUX8QbwgRqT0YkHxW7Jy1
6c4fErNnk1u8Krvac3xZHGp/kbHn/Sg/ZhfUDSwDIpj9JNJfEjYpIfi5CsPr3LMx
2tbiI7IUAQEXl24HnBLRIIM3DsDSnZZ+OLc1YSG9LuOBAcJ/ZxMQzovYZZbfHf6f
ngjP7f7mIzynj0gT/1ZyOoPTSIb9OiA6FWmX1aoyqblyyGwzlJ94WbwLN1KFDRox
E3LdIzsmX4zEWtq8oZWip1Uqll5t/yGgN3cEhTLOE3eZ/b+SG8HETq448cJdUct3
aSlQ5ogudJYR1+i8j1YnrNo0xOJUCCS4eRrZECHX31wUh5D2rXME9VHsQ0PMvzwm
MYrEf5TYSGYcbFew+X0TwdKbbbbyy2LXSpglHRGtj6l4CA6qhPE7Z61chYRC4njV
F9k41cemjv1awPyjq9FO7WadT1H6vmfUM8ztd8UsNPtDAgtHq2wtO16ySUyIuzQy
5Ou1XJXKxHgPVg3Cal3Z7qXnYys5zXmwuToKFc2OokbE1Z5Og58P6/8yxpEm8UhM
atAOTn7LS3oyhosi6IID3sbmGxD5sxWnWEB4C/a4YoPdOBtJlKY6HMzQolnzdZgE
2Knc5PznkwjW3G63Mu4a2606jpllcTTlyoq/WSja1cogH3/6j4klmppiLvgDBzlx
b5dR/S0oZ1cF/ItJPTzPNWkGmraDC6qFqcEZ9nVyEbOL9H5Oi3MqfWXfbARZcitH
oyrQ8rd4uh4AJsfRQQd4wCUgHpK/DjupOf9cKubfC5wWl/HbvRHj7tKuDAgMqKEL
l44Zn3R+8+SWvzszs8c4zWMKtnXtEDfh0fCyTAqxrSoEnxAJP+Falz3kp5DzPQ5F
4P5qEJWuaT9DDCo4k5CSkKvZwXYVD1p0IK5Fa3oRy6GQOA5DkTY6j6xCgeqUbKvQ
UZRKrfPf/z8fBLkPQP6r6OG5vYFbe6qeUp19pMESfcsAo5RYXJnQahEyj91HbBxV
YH/Z30OWM64FY+HBbonSE3pcY30OcsR/SwTWWxGYce2Us9gICpiuvnXKlF9RKnp+
aT1yoEOarUwFCHUadFqDw7a3n5F1y+Q0ZK5BuT4/R9+7699vqqXg21smXwBXmpwb
kAwRyMX70YCN/fYsFEND7t6BozKECu2pjaAmI4/QKKQKe76tN9srAmSxfjgbgFLg
JRE+1WIe7E0VNa4Wkmkse9OTHGHW3giHbvbZCMPvcvTjIXXIsjg6W05m/aInmqdG
bjDGR1jQL4SQTGzgYSnPvyrJxhnKyamplTBD5EuVAH7g7HOiNFurYAv6joDHRzrA
IFztmzavPJ3PQnfEN/2eV0/hvOhFC6P8I6qhRCRjzk4QJWOconglcGTi7GvheaE3
5JqSSMTFLKlzmG/fmu7u032dOqBE4QGiF2FcXO55GBiBu6619Y0pvQ+Dq8+V20nH
Ge4UOofpak7V/IrMeukFcIwnw/w2VfsEFG2Np8NXct4SdxCATN2+NcFH45JIcVPm
L+V8rwx+bLxuDxVmQRJtFxiwkDrko5gW+YkZflF/ddvn8Db5TbHrhnqHBJ4d22vw
4QBsqTEnQdTaf4XIN4i/dJasMcXZLB4ObPkJIcmBZ4fy/3LPUjeqR4DcM/BM4heT
wbVI26tArBdCBr+GTnF8sRHAZHD1zMqLIkmMrbdNnGjVjxAX56p1qbwOxLScVG0l
7LOxfPfihPcpsIUNuv7wp1cRlRXd95HYaZOJrpZcriQJARtI9vNzZo/BfOZYsk9t
uaQyseZ1Fl2pjfryBaupwpT8Vwa0MbcfIy8WS9aBYRrSh6o60wqlWQL8Z0BT22zs
xQ7MaaF/hZosj8myQ88mfXd6Z7b3izlR9dDrpE8D6TBUMMrwLU9udP5qlZjJTUNv
frO71t7vKw+s4YSC8mDZs9yIsgCoFlUZ6DKmchT4kRQGQp2A2GeymnatpJvWL08X
0//5Ompu2kwsb7wqaP7oAJ+wAMOkTXkKSnEi9kZKkqj/LYU1/s4By64mePWs6G/g
uhyTPcQ5X4vcR5r5pu4h20kL3/BNZ+fPwrty1N3wFJICwzgIC369z27Xa4M7aasy
kpKT58SjzIVliKwKmZ+hRxqYInreILIOac6KRycTdy0D4weF1j8RpJiWC0arohJA
3GMOZnsRpGYK77VLwpXiy+aEEaeIcoVQMRFycyZUcdlY5KxHnMQtgfdmTk2RoHhh
bdNDTq21vWVAI9veNh0gf57iY+sM6DUB23oShlJGytrEfYvRISRJgqDnWXwJu4OC
nxAa1Nssug3lwMEtZBXIankENw5bAAVozzSCNdRMJASCJlTPd1MP9FAvuniJs6Mu
SzYRJ+D+GXtVoSUMCCJ3h4GFVYseMnsQPuNbTGVbdjgYAeWxBqptLZA4cKLdfkQb
4/xUFSO2QctZiYwaXxb5vzHcHFuIpm+3zA6jF6qDKy2aXs9MaH0GbBcS7EYKtSRr
A/uOM/gBP9K8ZA6545hRgE5gtCzIE27o0c0boI42yKyYpwLOtLXRde2lwOKdAVwS
XAsE+WpqsccJW9SPOXj+MJApY62hYggodyRr5RHgs3gz9C7GCxevdmCKJjTIPSBG
LjNbD7FOBzHyWALzI+AsdKazzdNZZb1BcZsVOCj0zk0NnNSWUC179FDp5FNr4mvI
6SMnvMb2Pnn6CY3hZtMTSshauw7uSImKtV3bwcARE6KkIKDvnhOmnbaHmNVI7r6o
lXyS/VcdSFBHnBqGb5qfe/R5YmpkhI9FmCumjE3e6C40M78GD0IU3GylS2WOoMHk
vyKMHXhSlSOaWw2mb8yrLUIBDccUhe+w7WQ/4yZRzunZygfGAKrjGXPlIrbf9xqR
x5u9U7EbneHccBD5DIGer573Vm/7w1hwmQEII9TMLkHAtdvwz78BEc33xteIvh11
I913Y6cSFeh2Ip3+tWgF/TRAHrRIO8IbiHA0t66AripquhgjnkaBMROKiUr8Mpi/
mAoBWeL7xofP7A2P1dHcUoNgLdLCeU/WbmkfiaSsZHIdHKu/W4w1cJIRkT8xZhKd
AiJh3As5csSDyYl73Kwdfv3CEr5rlctOhKqrIrJDDE97iLmVBP6SCyRLM4SuoWy1
b5YqMcWes2UzdDIr5PJ9H4r+hN3J9fmLFOIghX8MG98daPDRFq+cHzNxB8sK+bZM
hxYV/TEzTdXTAxIZTG0jDCPQ7tSo9ht+Gt90Tx4RrNVnjjnnCxssOSgQmFmnZUu0
G+S6EO1iDT27DDB6eV3zy6L6E/yxrp13gn9r7/pO5oR+PiQOdyazpT25Vm0MZndy
NmTg1NeT8AQoFOT9r2ts8raFVf5tH4H6TkLmS9JEJliRIsRM7EGs+8JJRPP8hflk
ncoez/T1dOkOgND6dPmP8cUrgL/440zz9SoLKy7Pn9mjmlirL0vudOPlKWVx9XcN
dpxsLBTqNUPYaUL58+Afiv+rnb8BkyOtBPEBi+285tNgLysh1JAkVdPD6Uyme8zd
EcgRJPM1v8thJInJPIQ/zJRilYXtAniYoLgMCcQDKrQ7YlP+TZgL3HZFglZPkn5W
PzGtx1CM/rNJ9Zl6JSisgUX9TZPWuZmfKbIbPSiSIrbAAW+gkccyQuoiSutImy5Z
/WZDfriPWxkqfpUoXqdi7uhfyKMaPJDI5ExqAtY7g5EhrySR0VXbQuTI3/QL5Mcb
oIf+vYEwty/FRECE5ohgcdgn9uTrW3htk5Z3KUmPiydWMtA7A10TZxBQwmMEDqRz
LIpKXr6PIT2Cs3YYzLXQRdza84SEdy0d262Ui7GXIymOz29Q+GEAaBdG6xnjmBYw
wkn/Rt+8ZdAhbervFRljOOD9tOYmUAtLkVPxfVMuhJCyRCIuBtfLjzesmT/I5MW4
8rBkvleD8sF+u4YGb9Xq7U9yHBHduCeUWcJRnR1lsvsJpuYF8NmBET7HbDB4ohFW
AUfQ9OvBQcojkVzZ8nCBLr1QT9ZNdXx984aYSPgk41GV4yFvY7FhHI9sKKHBv36t
Ov6ydOsLEtzS8gWuRLVBAv+V7+xpxbR1zmi8DApdFZZqHpFk7j01Abmn8p7MHfvG
tqpkYZgr48rIVmcNcRaHI/GQ0Zkh16QFi7ORaQapnSdFIrYi+lAa1eGEqRVJljcO
lROhnbdm/HyN8wKFmkQhEDhsNwkPjvOFrENT5xr3D8BUo0WwMv9tA1B/gtcY2KeE
kRvhQxhO2kmO5Dfckfo3dj7Y3wQuCoypy3NiKBsZH5tmtammRCiDmFwoXjQPzSp7
9baVR3aA7qw3Aw+s8bW9AuIf7P8uu6P2eWhUAkAxYvSTjBDvAqYk7mfAo6wycalm
UM7qXpS4oIBBSsjG+4iZubvPXydffUd0KwmXQEIEchZjT/fXN/IfHMxII0Ry6WGl
G7lQfHEAmBOONHWUKNm4mvm4LFZggifduyi/UrPrS2V/PRR/I719yNfgtFj3w6vn
Noi20T54I+3WkfrgbBbloncEjwFwvTajc82w8DMXG9g4YspLjosk8PmDZEcutJQS
w5GZce4y9cEXjVwnUOOIV2YmlzBguchxh14LoQJ3XaUCeslOwl7bngF45p3oTd02
C6IgVgHsrHpmYakDtHw1HXTiNzK1xnVGHQol32y7Vdh5yvlXZzHfXeRmB2Z/2lQP
uOPRTsYUIVvoJUgW1f1Yw8lXMpA0UeUIGf37J4Klzg12HA7iGkTuKzqrssOuAWsV
Zjo8fHCusJOC6oxks9Wms5IGwJWcgsrKAAp7l09tt62XRnT8lucK9UwUfwLSRjEf
4PfxFEQQM05RT6TMoPKMUrhdTbR91LEcgMMiJG3VCfiu0OKYh7hHQtp1ZLYd3lcu
IW8W3/7zwd+NfkTM1U+Asx1HOdUjFav53fqzmcDqx9g/MiMV1Z63TgoVOHtrFnPg
JI8WqpfpP6xhqrHpnKhTw5HEUY3XDAbY5nAcUQ5avS1cIoz28tnP1t0qGtdBN7dG
FFaQ7yKg0PCAYBkNdv1Y2K3OCsbi+pyE4Jr+xQRvSKtkvHxKJIgv4lkqe6fZ97a/
jX/OuCXGQ2EdiqFKsW3NzlskkDiiV7f3e3tZEZrYMoPbKGv4c0AyN1o24+XPP0WW
xs1rv8nHsu6psimneC94JYZ2wtXIfzCyFlqcxCI7fcH45lvAqHz/syhLHV4Vwa9M
vb9ozba7hNzdX3Xh4OjhEtbhenNtFp+zUpIPVkUvkniNIqp/wBZWJFPosjp3QnS2
OQ5pq+mXHbqF5ohQw1NSxiAn/zmBb1PtrAB7L856ma/gc0UMAVukzeaOmbRn9m64
tbCNFNimVVxWhaRBDsoJXyQuN4lPqnzefx1L8cEFNEhLxyuEwIHu3Kwkn5361T85
tjxsL4NzA4Mb2CgXuWFe2rQxlN0poZqQlpfG/InMAdjG0aVdMhmU6xuNY607BNjc
+mqCvUpZ74svr+jh3PVI6R0UreGQ6HLmHAAIKicrphYm/kxI9m3MeQ6kBy/K/GMG
36ESEwU1z04spefv56PWX2tE31wHwngF3tqpevUmxFmIx8nq1E13ErNpKlF3vI50
tm7209meYwEtUd2iVrGQLLYBkK93tXEx7DHkrcvYG9NnXOnyEqcCMWv9EAbZffAy
OQT2sblKduOIiWZycZpe8MIqGVBjminOKpWTAJdPVDIt5Noj0H957lhhyEv6hLgP
KJJtCVWxblj4iLMRn0hvfhIPGm+FEmV+elU7r/4SrQ9hlLRwy1zg/R2XeFz51f7x
LPbuU7RCbJcGriAjb/xzqeAdqPGRTxsgkO0FYQSAqqfemC30whLmFEh0B4plBsx/
50AwpGQWS7bPZadGIkYVVT8K1bD60qJhME/M1FNNkxjIzQybtRghNRSz2crNP19p
4XtZhaD7TPTkmulwAYkxw4f+s5sV0gXyhk3ATi/SQyg50YXo6ymxigPTIrypbPUT
xNOTgwJ3y26yZgonRjehXK2ttXsxs/RVfwzUZnM8nESPOnnxGnbkVPMIE+yB0rKU
IDOWj0UZ9WUX53/kFdGhpL58ix0Bc6H/O3yTvtmJWaJbtZJaGAJ1THD7E6yBuBjb
4WwyZ3nJe1wKa6lj/iB/yzLM63LKnx+tHAtcLTMRvAJkk0N2K3cpCZdUJM+RjQx7
ZL9VQ0T49Lnfs3HLG9RKdngh3kr+kNZR028bR1d04rHU0S7SvlTlA74xwfYBP2Ww
4H+/4HjFxvR9sR54K939qsWGHEQoMZUz3KpTHTFFbZwvUhvzgdkDcaZTcuMiHuET
7RQ4qwKm5n29WQoSfT28peuJnSBItcjQPL2OTypqXWQEPQAHg5iaiU0ZeR8UzhDr
AIDmJaLMiET2yztehnZVP6U65cJBxr9m4ydUzfGE/M/VK9FoUX7BLgJQv4bjgzPd
Lc1VMWuUoCpzC+ca+F+ncBhLsz9IxVd7pz7bV1Vn8VSIQ6vwSAqe40nWkqEH6cKJ
KHtyMcgThq44e0iFrHskrtVC3ugWc0PeLekZ0NfUnw8tj3x26PcvnJp3GiR8D7Bm
w9ere0EDQLaK90j+VPcxbm2/87Bh4w+ApUQXMrdxA9cC4xFOKh6Ljvk8IRmJVcul
UCLQubIay1SO+++4SfzbgmzfQp0KJEa/VwbHprBuMBTKZxcFLgGjTDqNGCqKkW6O
YSB7t6W9UAJCCe5pI3Fg8lrutyCycADOMuKGCj7jrZgCGsLsc+Mm/KKpRBcPo/Gc
2PkFbf7oDMpaX9BIe5oF0A6uWyrKo/woF05J5niiYfsOuPltenuKundUauYtRGoc
WLTl3Mqhe4o4ed/hDor8iz5CF8nnY6Mbhm1nkyJUByyFUoP79k3I5S0FVL/CfiSD
Co+VUsXAvd6lmN3R5YJcy0sOoJEfugAT7qoKkPgKoX9K1bkf4ckOrH5uHJ5VXdGj
upRS9+fuMBP5zCHc0122ZTA/EmIrzQIHYkpbkY44b2LFa2T+IJhJz7ggzhDJmkzM
E0fyM9EOONridpBpFCd9bmMNrzmDRMjgS5IpcSsPCw9HQ67MaYNTbSbBuExE9aRV
s3Z12ILkaKg+tme2oNt8Nsn54sxDwURPP2B7GbIhqaBI+qrYVSon0AUJmcw3ylJJ
g6NwJFGxD5d9vpCcawmL9uREp30CzhzCX8r7gDVtByzR+sZ/DzudzvRGsDLSS8Am
RYhhGnBxExEW/UDeyLdQ5A/BR6FaAqeEMrQ2OTqVN6K9+8SCuDABDP6oh9Mhn6/n
59ab2aheB77jutWL/cdJp+SE9Y2hc/dby4Pjd5YbJPTl+MGGyDEWAT+p1O14gzcD
2C8F6MMsbwzwzShl7rRllFnbpckqwulb+RRmvqNTW2zq/IBF3fKTzbuaz0Pvnko8
fDvrGopp09mYTlBlbYuVNvt+wJpBAb76fbwM1Pp5QDI5gPg6V7PPXdLk5N7BRlUU
zA9nW62x++UAarK24hB2wXj+wnytalEOfucLVpfL8i96DbkKEbnlzClhl3Uv6QtG
YfsMPdcsSTd9k1v2ys6L8DljHbPJr47Db1/YrDOW/Oz+OpMSUbkFktIQhCkHaQKr
mweVNHE0g+aX2yppjFkxYeRiUKDC370JVonJpPRFjZwio2p9VAgPiFHPKlEc2Kqh
QyyMy2pgnQ2nALhLcSFg3lFomwhA58SCONppWydUfejQ2ZZOQWwyUfHnnTNWEpEt
DyqoBTQZ7CZXpOPYASf1ewBhyCzK3q5wh/nUE7Y9pDbZLtyWq9m4qbEnorlOltDz
j5L8YEvgVLfFu719wuR8DE8eh1iRGl4TAobpsvB7Eh7367mxQbyUnVuAUs6MYB/2
IC/djTZbDjvOqRWm3W16jbMvfuoVix3zBPcWIwRZrSEXAzGJioRXo9Z1ZibXCQxy
8vuUtHw/izYSvXPK+Acp0xI+npF/flOiJWEjokz+gZXyAA5atGl+AqEOzIuFQJdi
j7qLCWXm0bFRHbfSFbzW1OSt/qfw7dLQe1hZL0TDporDN54WPKShxe5xyMdb/u7o
8F9lyMpZ0SaMpmKAwFP1zAbaCGQlkO8gGL9pEBnBiBYoLS/GhB9nefEHeMJF6B3F
G0Q9G3XR+Fnsw5cGDSZmHvWHg2xq4vgQlK2eTuBETrO27lKqS05GrwUpxrE55j9l
eqaebwtAwTx0XrsmbED5KmXDfiLfJdTOi2A96uLa3EhwJ2AUb+foGEjBTXoq9A4M
UqrBPhy6lnKDqxgYmumATa7go5D75Ay1rkvRXT4FVbUYLhS3e4tBG5SS3fz1Jo40
dS22wPQBo8xrU9Ty0sbUxKziBT9QCxwOOKlQjDrjvSMSk/434uGpv3yxexo3bvrU
QKLgBFfsiNZy7i+V+zdUT5M/JfjU2DXpyTN9eLt/veTN//7uG5RONNGYgWOZAIru
fEBUMIr6UBNeoev/HTJ4p4XtNicA5OBEVDTB6WGPjHE=
`pragma protect end_protected
