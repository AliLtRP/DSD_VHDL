// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:35:25 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
VWQDDtYYPrq4eiAqj0J3+5eGqSUowhgxJkKkvn5VTPnWwoT8Ze4jUHAv+4ZUj9qx
ePmSYtQL4H1JxCkx6oTgWu8CFt22MpcnJWism+8pT+OXayXpIajURCK3IZVqGDqM
Mq8hObrMeIGuCJXVG9O1N3uzsz7tpEwJG8H4VKwDdk4=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 13264)
3gZhY9Vm2KHhrFMsYQOajguTrOhloUtq1nq7lHYHusBJZYC4GIe4reDzeTkeSCmV
gF+GcoHT+e1aOBN086JLroR1ydTuu2JdpZpwB6Cqw/EPz/YQuAE8jJ2LAZBrCsFx
n45XIgt7IdeOffljca1EsZDKvZcvF0WTN4oF2HDe+KnYOMS5S4rA/QNW6tV2zjEz
8jFM9T6NO/AyhdtKOCS5KRdkaA2NaAXOtlaVJLMLso+Lnbs71dUOCUnNEjaLVM+V
7UbPyBuJDxVdTlBhqed/XkasbgPHUOcDh2QTB3uj7iSiIsg94FsA58sL/vkTax92
xzGB9L7F3FjBSZTFUylZiwaj2eBE6YSRax7Y2mqwWiYGiJF4I9etXqxRZsEAfmVN
XgtMEK9A+BXg0FXvqaVmwL/6KCSH7q9EwA4ua6szi6umCVocHU2GfRUaSeVhnl8u
w/FacEJfrc8Cu648B/LuJq7F7y8kLtWWE4lRQXt8iRbd6zc1Ja1z1LE8N0a0Kc4Z
kPBD/0LEw1P+GZ2z5x2tJ++BWLrUdyDaU8b/ChL0ZTAc5+ZufHCMX6lmq0F2Y/cc
uY25nZVm1973qba2saVfBwqVQ2oWtRbCKR5S175hPohSVIlPLXfHtLBNsCa6Ac8U
LaNWhZOiKlgnKW4KIgPEyyvD7Aa+E36++5z2t49Vwwm36ujfHkveMrit4t5M43QQ
LavAzWf0cWBnyaFK/Ecm3DBYoaP/rAgp6OiXloa2Abs0C5fjNR96IhWWsN9ZvCMP
0x9WVZK3u5LpcDRcRVHUfgF25EmdTB8ND21i0ySRZUY0L2ZWA+mjVY4BsSUcnIKP
dE2R0SqaOkquyrOnNMI8dpCCwWqPiVWHxUKWNgn72nFL7LcecUXqHQag9iU4cKlx
szgkf2WeL6JKKaoOalucjHB28GGoSzox+fmKUzfqLMQ/qUeDyqScAHn38VSFxNbY
TfZQgM3WhH/8lly3XetQtWH4FYoikcJMQ31z3VD2j4lRLM5LoJGs794q8pWPf37m
fQWb2FDjnMj9myAwkIbYJIvUnp2f6lU8ajQewqkxh78sTfCvxyXpzWQUIIrC+9Cj
1uLpmRmYWYnGu+abiqgpf14gg4Frt3KeVrUC9HCn2GTlK2RF3H6yIzHoh3Z99rZ1
Cohq9gERhQCRxgpegH7FqOWIqSVFxHWZCsxcOGnI3lslSnPE7HPWeAarQpxrUqwe
RO2Tzm/0OpLOTqmLiDJWOMQKUgq5Yd4oeey4vAWxcVPllIaGiKuZBP+6R3zBhcD3
SyoZj8IChGh9JMJH7Bf6yxIzCmeESOBxWhKwZnXNt6Emoqy7lPw8QDwOko/9QM0b
DRMJ1Rl+9i7IrZtO1QTw77nSSG2lmAQyMyvn6g8+oPUXPw88Hb2VUSiiXGnYKHcI
vqbBkWOES+lObu6Kx8MJNxwePFql4vo2ucxfzsUn3YYzYWA4nMhgQb36bX1YiMSv
GrCynhmObZYhCM9B1NUEPTjJTJNULhvyP8ZOYi8KXGwjiouM+4LebDwQ7s45+dao
6P0aG2a/TtBWfASoOZBdFYtGyfzedeN3cye/2yDpWEkl7HVwUweiOfdvjC+Uw3lK
Haf7wmojfswhUqMZMaJkdrPuAbVtxBEOJ0s3DVR+VIWV9/1xFeN4XZWhBf5g6ENl
2CH9CcfokP11WmqaIqQXGA/xPhCGMoJUJeBczQ4kWzXG49U1gU65f28mvj7DHoi4
pUNcOAID46bzCkqoz3JeYeITkDTYj94bt60/AHy6GqeTC5GCXbzTdK9M3+ibEcHb
o5C5hsb4GmK7+7UZRVPuFRr48kLFxGsT8HU7Uyp5860wyGC+xdpvMzK6pCI5osfB
RJPfLmNcBt386LRg+HRh1ZCWPYDgf6IlZ42CkH81w/7EgtVq8Kz0QXaD8rJwWUAa
x3hqSfzmWbiXJqoTcp1F/hQ+18fg20k4DCwjEgJhBFrTuU81FksUJ+cfOiG81iIV
TsbyPT9VOskA8sQGl+U7865LaI68Y3SYHu3/VHckkGn8N9mcdjy1aVCSN0P6az4z
d15UZXjXQmPXybXxCA9qQWWptGKD12E5/yN9gohkeGr79VneUSFC7dcaK2qKFcc9
Wdby1//YMz5sDYbyylWZVOG/AoeAb6j6a9v8qJJLN8Lizyq3ib+m1SFTtJX3ajXx
3alreAGxPhNUMipm+y2zUCfLW6Cc4XaHoKYy2XyiSZW+Jm6c3+cmueBPm8eOOfhY
pPRBcGbQgxFE0ZidmPvuQ3+Y+CBwHBSMeq1KOjcXlKH+fCrgt0I+nCGOOPpQIxx9
JTE9U7FX3EXwUcuQAS07lruU5+6wOOKVJD6ARv4u263bdzeSChZI4Tty6HzmFe2k
/yTHySTdos4D/Cz9m0vs9+lC/cY/c+iM1LIUUh1tBFSw9ez/tofmeDmZDO0KIJXx
cMlum9/a+RkJdawveQqgtziZPzgkRP81grn81VDx4Kd0OGgI9OOFuo1Sf5+3o1Ic
nQGR8E+iXgCbiedyo9nufL4JqH/b4GmULIMd3nxL/m7IhNaeu+904FSMbwv2WvqJ
1684tcgrVNYK7JbQv4fgAiqQsoG4v45B0F6TcZjdUMjUpHaZZlRMcqGz/nCZrFwC
ooD5dxbqKSi4vwoNZ24D+acw8XrioINRhcsXSCyHDoV4SWl6s/jBQoOCTRs51VGB
N/pkJ6zowLslVThrxrWlFm3hZoz85gJD4Y1UBmOhAlSGefytQCc0wHOdPutT4t1r
5Ojh5+Hf73uXJdxR1941mm+5bs5zrhXpHytb2lzooVEyxlHDrH/yb0LTkg1Z2Bml
4W/txG2PcXJ2MwDfRNeeq+HAzKZKCnD4VJTtoY36VHXETGGWfcmrQhjWARu+yC3W
D0gBuOiLFGEcPED6EE8ZyuSupf5ZO/9tSK3UMx8gmW5tHp6CQNOZMhgBp5ZjBhQA
tYiVGxXsBIpnI9ytffWpxOLrax5p47VD+Zqw2zLUR/8agvux60vvpkYZRcskk3m2
nYvETS80OhmG3NSlS65z9dXdtIPGm2XCmwbQqSWUL4QVTW0Df+823NjKYAdfZca7
9uY/bU6rHHxJ9mGzwEx5p93rapD85pq9OrZNhjaeWrqvHNeFHL1WfyEXSh1cLnT5
GWj2JAAwEEtG/nK8pa2GV+9lZh50EaDc5wDyXIQsmoLkjtFyWg6hW1+g8fDf6Rbt
XJCj3JHMZabS/lee0UVQctwyQwyUuhgEjG7tHkSON8ESyM1OWjDJlsIvUNB76jdv
+XZvV60Qgo8AiALfGEHxh8CJg5AfpVJze0g4ETqWc4NeQtvTXo7giZHTVmCLUCLE
9JDdjH0XQVYxT6bepg+t5B7juOuCK2dbWrqTl3IEgGH5GTdA0Pti1jebRdjktz1/
i6Kln5Of6oK/u7x6XtYTshJJFkQDd/e/qpbLCmz9Zck9ZWcqGx5OLOz7hWWNXUV4
Eea9tOu733hgLIOVXWQzo/D5QL6awtXV79xZNmZxc/t2Pzvh4rrX4ouQTZ16kfjn
FVOIvM5sxrXfpqAe7DucqIaYrrZj/9nmpG2IBGALN+UcKItBYybxK/+Ar0o/aLvS
ZKAE5Wsn2q/J8KBpG1CMBlzzRJ43bMcM6UUfk34uYSBO/5hjzDZLOjI9/OjxmRh1
6JmdbzYoFh4BRbmqpusf7noaJOLzHw8vSdoqD0d+BiXXtiesliRzp5cJITgeBZ6Z
z95D+YZvL57xpUnwPO8Y4uUdxrc7HfL+vHY+xD6p5gxMNxPX89lUVUM9L+0wpvcp
defiXGIURwVUQRMQoSD12h2GpWrUfwyi7wo5SYiF7F44U/trWcGLv8r1W9WjQt+c
LYuJvXy3CF1WqQi98kvsf6Hx/jaGOMA3K/9eAtg5avWOuPiiwbE4LWIeMEajJxYL
qNx33z1zJULfxmFNiYfmcrSftzyMnze5whEZ3LWsS6D0WX47Xn5LMVtNSqfFeR8i
lRPMS76K1OzaJFFJZ+beVDIOI5v4Mkr1Bgzr6JiuP2phhZdSUBIhGb7SAhnItG89
uqUmLadULQG7W5K1do5zCv4TRtzcTkYX7pVzAcD8GDXWm2n+/OCO498gIfxOCJOR
q1AU7T8qoCdzC6QsBZHxgx8dHLvLfufPR4dQQQYacD/xUFGkiMk2KcdYlQ4WvKMr
9BitgAdAk93LwwQYBunrLmd+scNc+W4LsdRG2Bpv8nnTqeuZfRSJRLMuNhe28nof
q7aA8AcnVi4Txi0L/AD8pRXT23WoLeJCg9DFZta6uBb3bM+c+U5ewG+SgKAedSvn
oLrufezg1N6/xObO1yZc3GVpMFJKlpXhPS9Jv4IB6zCpApLO2KCbrMuIkA23vl7n
N09QqWTT08UQ0pA9tlnrHEaSHruJxF0DcfJ1HYlUzzOt3Dz9Rs3oHm/VBOpB28Vw
R+i8uslSM5mU0yT538h3dpNNFZIQPmEXZl3mYwI5nuSam870c7qbUlZwV+pz9x6n
U6+tfcn6v1PIIzG9kHJMfoCPvb55U75TFo0QELBNJH/pGIfe9W+u/626tc8s726c
DoG5OO3Z0fQvL9z2aBj3AWvx67uB1izezifTXVi+zVvdqqzZLCpgPB3USFyWPrcg
plOsJz3VYD9wMVnYBiRf76L283SKA0wJtupT2J9xxT8nQzouwgaA653cLp+1YY/s
ngel6ZVS2F4qIPKe2wrM13whVMHj3epJv+HuGp6EBNIE60rl6CJdb00GANjvH1Z6
YvGCsZC4njn5gTLQDOn6ajPooWJj1hU7aDcLx1VTSuIY5zs2RPex7ncmfNdkvtFh
YkRRIEe7rQIMhAWry4rkvZP+xrtPw2sGJ7DQQxP9hpdF1UyJdSlhxJtEq2C/5Y6w
1BaPZzplRzenyF2kFSwrF2DJgaiAwxUQ1FJYTzRvc1aJOFoWc9P/Cvj1Odcp628R
Ve5lCX401BR61plVXKZPb46Hh5n7xE0R+LLvJ5Z/qnX3gXmk1CZH1JPvRMUhUk0u
Crqr9jgdbU0LSjD5HUOZODh0EUSYKr/VUm2HA5AoG7HdASKyIj5PwXgw/Npt4EEW
hHkydiQdkBqcD2bcVT6DtM01dpyRzRtYJzdrQ2HhrYAIwfHyn/VDwZqNbiRBFE5J
41fstYDcQuna8Zdm4tEt6+vaRft2XkQvNbdm9J4TZuol79OwgAPTTy86cfQCbWsn
WwIlorDL0e+XbreeWGbQ72oyl17WD0+62v00X0k3v6iAskY3z959JxaOnDLV00Kh
pqhRGHdS8DSEMgZGvZmYQ6p2b7E+dq42c3jJXbnXZEA2x9DTP2aRWb4oVGdhhvUY
mn/HqkEFxeNWp3FyP4e96hnED/duMDInn+p2XzOzx6yMEGOkEZsgyc7jWbtdSMAf
UGbOk7NlrEOt1aI4CSwsM/BLuQ3QE++8Y5JrV6yt/OU6Nyjb2ZdliZnoudOW8dz7
eSv8dl9073q31IameoPP29PbK7Fw0bDEHJFKkE/ufKvqAvgpp+jLASdY0f/ZGTct
GoiwE/3Bqftv+ees1eH5MtDYEctnndWdhomAPD1NJg9guyFP/pq3JiQwXRdTe08T
tAGBn6Qv/FXly31t5yQsccsoclHbGEYVJOu0iKztd3vZ40/xeh1LaDu5QZIOR20i
RM0D0Wo4OvfS0r6Z/2fjgvSlT4aguFDt+dcpy4vk5ZI0SSpOW38WDm8cyIYgN4Ms
UJW/SLT+ztzFUAdYHsnCjzm/TXVJRL6dwdI+qUaswr0DD5CHFJ0v7kMtniM/MYg8
sT+SBcFyAju37cwJTg6ykgvEo+Z6Jv8rkULMpg53UzBoA20Uor1sZ+LzhtgCK5If
KfdWyr10uhlrjMVC7Ec09feyfpZPoxrMkIZ7q6Fv38zKUd4Yb6Vu73Qe7F6ymOFJ
k/062hOcRr9xLDVoOo8TgSo8kKRa/llsBKQZJyml1fnfF19+al4WCu8glBWBcfUm
nJMotc0UkAqhOpdngncyUD7Mi7/aKWDZG7PXwPbzhxcxiPywvHuM0Wc2VArauSfb
sy0Kpm9/+omyN+R7njIbhcdieWbQ/7mHnOfSYYhRY/KBE/q8u9NVj35QlZ5gWz2h
1co/j++xSyZxjxX07X7/o4Vc7na95FW6Rsp6NLxYPfggh0TeSgujdTVH1fO/qcXz
/QsI7N3lPXiueMk9pmZObdiYTmX746Ox1fTd9nByrIf7nLL5yyeuRYuxlJAqmQH2
DfZ3PtNKj5IkdXCEgmJfiUX7fPeo2svHZFxIkumjHTN5fDKuWjdL83LrpaAdSPcR
krB2Jswkpa3TAcxycRYtm6Rf0D3PkTtdncv+TyncJoQGRcqeOfNBJEFJAjgVAlPQ
E7LXjeBieJiOXsK/6G4pZbZ8MkGm63ozOyduaUoLJoZ1RRQ95O2kmE879aXKUL7V
JFy7+DY7fdR9mT1rSc+pjR3VgGV9Ess8N6suYhtHwmdsbxNdYSLWyamdcQiVmhN4
nlVBl5Qi2V/bxZzTWow1DeyuPjXauFZEP/Ms5iIptqrEA0zhv7joWs3/8vqEjqOk
1geeLzQ/SRuXQj5n00ugFzlCFc8rfO8h3aXwXbGXTJzKlRPIPmtfnzApSwyaXw/0
6iuQcV9z+RadU9T8hC62fw5Hf669fyrZuT0uOJMI/H6QvdymcwIqN4LNB8W77SQh
lYnuoY9+ofUm49plhweFupdoOF749HvZ+5yDDZV9+e2ueAwaWDL2sqK28+kYiyrn
Cie3slBkrLtmpQQ0ErOayV0n3BHhZpmHMA80+O7QQxykEQGKkj9hV5z06bdQE23v
p7VMyE5WZGIXnrqOdfMPKa6X1KirKGoJPmHc64Lg7nA5+qlqsLqfltmYKrdH5+hX
HuiC0xI8oZCRED997JXrbP0X7y/vZOnv2cHWIed+NdU+fivWjnrdTTInevs7uAOB
FJ3i+tCH+bajJf3Q4nKW6TfJUct/AewpOjvuzp+gimSAylGQfHTflggQyCMpdSmp
UeTK7GWV7foNxvb7H25bZlPJLcTy7gBGIOJBlKUKzibdcC7WRebm5IJv0Ic6Y0fa
9gAZV8rA5g2LItQohJb+qF562CCd170uWDPtqpqu6Ne3/EzczBLNglYKZ+LUU0iI
nh5PixvtdAsSpUyZsI8CCRrt4hAFi6rbnRMLyS4TbhkYB8DqFRW/XaGtg0rY98KA
NFYzs4leAFvrJ8DppbNvgBUVJqTUANEJzWhKkY7927uJak9qlBu6yhzDto8f9cmX
tBxNdUBmBannFBOw5UBMhzhWLRaTa22e3ppPZgPUUCLOnkDUKtzMjyQadu1o0VpO
xFVa0iLak2fKbq0lD8OoUreP9v6HcbyNLjRV2/tjn4eymMIDCcXMT9YtzCW125CE
0Z+SN9LFmmb1WZsnts28b1rS79FoMgT5LEijX8UazHV1Vz8fxNjliyRSrD+R+6bX
QMKxN43rlsLrnFd3G9SzRtXVPzW39ydFUaa83fmipUTk3gFVmJ3XqsrruAaHbEXj
9cciM3mfhecnop7QYgxUxHKG5idFi5oefrg+lUaPiiIoK7OZ1SkoC3vIs102MPtn
yfEFodD+enrO4PR4h2DbWoD8CUsHkqFICHzse8o1i2D9/J89XRBabHePGO6dN8Z8
AF+QBfiR0/YbEvAGzPtTaXfOJykxY7REWtIOkHCvXCTgsBx6LTNe2pXyP0j7ggUd
g9RK/pOZ0wQp2gXKJeTO1Uueg6Ae+iMo6u68qPT6N1UUCK6ME2645s/ampnsfLOn
Mg0L00qDP0F0GZLs8+4PdPEz7cGzximajrSbU4yy+Hd2e//DnbzWqrXo7HB701Zo
yxg08DuWBhhtshIdNU+oC75fSWS5OKgH+ErvqLnCigIHbIQpBm6UThp7qxoIoh4s
lKrKKIa4Yqbt5+uVbDY0TEddfyIOLrFtZiMZT2Xj/jovJU75ixViXBSLqSSeH2qt
V4YK/xnWX3C4VxUHzAWT3RPUPatH1FNx0vPcFfOBYzuYf7Cd9Iv8x9hwER4CK1zR
AuCzHB+RpNuDQqsu9I90wvA0m+8w8B9ZeuM06nEU4zA4+YpH/jcl9xnXXVHEwqaK
126JRigQdUfiQWWMqVXai4xENEHpHgyNA6m08pSNfByhoP/wLGwjSlyEbY2AVyLF
/5QrKV+Fec3Ybq5cESiS+zsqsBeAtZQsHKiCw7E1LdOBKQOoGNeGIfAw33Afyguc
ZGOu6T1QI7YgYOXd9DV52cN0hefvWS4ULnoRhp/Nx2NaoCu1VbaZTLj2gUtdayJs
iWz4z8GrUCbO/X12B3kGBm/LcJ415Q5cRWXudSOcltoDcmk0oLO8dIwHol9pQzLW
GwGRkJfhwZ6C8718NBbXdAUya9dtsHst00JIoTCtx3S1NL8E1PEVXNrkUY3/Vitd
UibZ8L90i/b8k+E3AO936uA74Jb4IvdImdAtg5Ike4H5jXNXQ6LFRTKhGJLnVPiv
Vk1XPF4haomppw1DEVo5G3+SQghpsow0Nv37XEsdW9btx8Tovcqm1oO3LN7QBFZG
mLcOm2bSa6bhp7PVxubD5SkbNalAnOtIWMYbp25HKQlCFdPVC2cXJfPl+zshZQAJ
ve/jyViPgm/erQrUyhE+bOzMiQX50acxQm4hdbzcjh7RhljuoSSQbuQxmPVLwRv4
3+wgiL4lmQ8Y7AbH/kX5wl1Xt9H6s+gK18rXIFOlsxc+VAOqdxjFJ/t3ZHUHgcWu
8Z4TEeh8w96LDcwH4R0oU4SxK+cacQy/KHs2TkuUAE9Y8h4FDyYhhRdF6llROjM5
RWvqcHPi0aZHmbSBO8Qfom5v9JaWO7oIhLANhYrGfT3ztYroKgBhdqqWYC2q4BVs
vaYxQ3ge0D/dnj/wYIhmh9O5LYfNBYwelNoX8stGh//vCxQYYfP1BCbAY1DszJW1
ye0U5ejM8BwPWIl8nFfBSHwZrYaq2fGMd7DG0X/ndk6kdxlKKdtvmqKbxxnfDGch
EfkJxHl/O3WHE3AjvgDEgmbhieJ8keKAo99pONs/jAVARypjn7LTiLAoYjmDRuYc
IX7eGsW7tAw+MPXejiy5YnaoLmWHFAKXpO/b31Y/Y8c/4RN9NmUemiRdVO4WVgEt
6H6NG/IkrPVdlNoZGmr/JM4fbStJSRwhOVUwQs2CkqwXvtXOmsJvj7fabHY78zeS
0wGlTvQ0p9xilVk5SBqyzmp5oncck4lQS+5wf+g95JeyGbSkDTAnZh7+pOZIm5o1
YF3KL95y+N5MUndftn8sFUv1QPulBt0n4rqrrHFzS0lLs5EMAWLhRQtUQHVw9V8F
JyFdwV04Mypd4cof55RwqFRt2SiQIeEp3JdtrWKc2RXLDF/hWu9gX52Qx0cIOurW
hWWGXIcnufLQSVHEI0HLPssbh/N5CU7/FVI53uQha795mYvcyafmGPiGuVSfVMsk
N5VTIMU9BnpF3W4Vm80CrTaKXjLDKG2mZyALa0IlD7vUxtBxPzSNPYL8zCRdbwyU
ssblKhqKL6jDxT1IGvdCuZN9DfOzU4e2WfUMmQJN/rVu90zzeH8xFw8nlur946TP
7+S3w/+0H83YtfCQ0e5I/2AJjx2matExClIJwWVBohHGGUBRg3aXhLz45wou93yX
lXcCJUchNavYP1JQN53fgsH9YnIkuTOzbMnelVyfC2xvmuSjzaOgb+gbwnOwZmnP
CHxWLuP/YQIw7QexM0L3/VROCWTXIwaccpKBkStUgQopuLaEWrGKgqFFNttLK3a/
LnywD5XFyiXU+mdV8pFfFm4SBGYfBcDjf0lkGpeCv+4mEPQOZtYFvFuD8SjWK1ft
/hRO2FHNbTB921o2SEeXcWhoDPFrI2lF197AXimU5RtyZmOB2Bqm4lWnHe4+pj/D
bugciBvLKESkTHF5wsZLMewqzau4QB3U+7y1kqlmp3HB5+kEaWb9qBV+m5CWrhQH
Mh9EDcnvsQWZgm83fbim2gCo/EKFGBtSSOoMA/6Qk5NOq7YvZy/BvbkX8F1jcC1P
dDnmZP8T4BWv+Qxh21+HWCnnFllQOn7b0Dug/Js6R2CMxu1Y0XC3ixoQvPcHEaJv
6D/p6eJc8/FISrFJ0EsJL6ftnq6MCptfLjyu6WIPkEifqns/I4eMGEiRUTOW0jDC
BUDOb5gC7AuVetEudBjYm4oZ4JkFP5bSjcmdxM/T1bE1BFgsOaRKvgBzLhLrnU5B
Y53XlJhueS+DQL/w/02LwW/RsD5qCrJTo7geTkaWzU2bAxN/6IOIaxZWpSVAa4YT
gkzZ18FHXGoq+YhTLb2uWzOHGiSWBzkjRsJU1UIeVt1RL3f9pYbMfxSpycLJW/CO
j9qLAzVJnQhYJNCnqSTDwSIZykViSh+t+GUChoYTzC29PHXCE6b92gCz8nyOmasT
ufr8aabohWxkTnWJrSiDiTS8aE2633z8ghYxKOEYl6gBPrPtAjOlKRIhDDLjpSVv
qMvGI29LFU0fjdBDVTbggq8nnIfw6un8ZAXkdxmp0vXBE+rvK/WXb7IdSxwKiMFm
mB8ROt7M5xrRhtuZfQlWPKcYmaTCgAitxk465ZF/kl4TCGbDkDFqswkfXlMJ8mUZ
jiMPdZ0y/IzCQLdCb++f3GxS8X+oor12swmWSgqdMTpG1Fa7So0mvJMCFs76fO1g
CANesGYS3iPMwczM4xQ/6PtVMILMqyIQ5zdLWHtLfU1O+Y6vOMRdwLCbxTVBScBw
gI3VwTp4Zh6y5sy1CoZCHppfQ0JeJ1kdSj9nLNAbmIseGeFOHIw8dy8iMnIu8dFL
Ecd0lq0WqgJWeUzAQFnwcJxZFoc+NZncIj9H7JmCU6w5HH8XXH14kTuj33WA91HV
L8lhFBfuO1jVnXxJjkZehCuEqJU+eWNNhYXV0Qo2Z9TGfALAaeYnZXLiXxLuW1xH
uY8UypwEVXmGVpcXA3/MlMoB6QAtoOo58VaIyyXJPKImukIKiu7j9Y3AJ6aaru3z
Olm8BpRsqdMihVANYpgtwGDbWk7l2/68vwvuKIa4pDkqzwDv1rcDwZGGV2WHyxyz
gLG6pe2imptgJyJRiHBxqke4YXco44gVq/Up2HD7WJZrFRwZZIPDTJK73NhU1aSS
t9At47mYmXN7FRNPqRw/8iGfD6YNGlUX7mBcU0uOA22rGOsrCKyYT4Y47LSiw9w6
F+NefKhBw4i6eR33vmKdjTm3LEXrz5LDr09ITNIfhphnGiNyI92PaUBBejIx9XXR
rci72oRdpduWMag38W5KQm/qHyWxzwURIgLlR4QUrX/3Rsl5q5IYu6BylCmTGI6B
7rtQIQGLG5DxCwLjkO1Q9lIAMuhU5CZQuHPC3GChj8yqOby12qnGYp0AOHgCMCAU
JS4UtTLwXQbicPdYkYOSHqfJFbsytcHOkG+W+SjdpwhX/xkk7GBwCCh0W+XV6RRA
8I+KmG/YGUAaepz9lBAZnMZakzqkzVImwMNGhX/yuKIFiIPz3VTvNSLXVhwgaMv8
2/Nm9afTvatEk62RPTqdxe3nrH1ntINluj4LReP/jceslyUGID1ud1e+rZZfnM71
N/QYOb3goyxeC/LFw/x8EIBUc1Sghl6DWQ70BEGyzPew+r2kqCRfG1FJL35EgVvR
ro4gU4PlytCqvqGfbWc+1NdwagA6GGClo7E84RPp7MmujWe+dmEGgYvVMpTnWdDK
CiivRGxE9CvbAQKWXoLVP+N8NOSsB2hiOiBJYM4YVnm/pz1/53DVojkecaKiT6sy
l+19ERz7eva/qSedsJ8fSwUg9CZpSQ5G2+Lej0aoog54aI2AhpAXsG0mAf1Bl/VC
iQpd2KAHUqOIFoylc7Q124JFXeCqEPRcKcl+oR9Eiojf0gW1hveP579oTx7FZPeE
f1GX38Qee3O60CaQhqmxq1O0snbqQYimReQFou3e+9yN+TZ6xALYzl5FfOy1xaNF
grWiSYB9QbnhTaBsChYqU/5NrYF/VqqYsbrtVHaI1nEZwMtuoEv0Y3/ebmqgJ3BM
c+PMy1GUD3v3jzeXO6VbnRlD4IjfEPwJ0IDc5Ut0RT8xDg2XxNKvs1rmntX6n/wP
m7/IupPwLXudx/f0T4cSOb1hXfA9F1dtghfOYWa1o3IMLoqioWmpsXEuknD7XfWo
qVfOuvR4IJ84GQrhjWZiz14wv+zzE2jCUu9y1CjoEVhY9mizmFVI7HbOKnjl+H2b
B3f1ZTRqrKgVcuedrWiX3XLL+qLy2Krx/adZC30c89AKbzzHk2FC0oDHONk94jnl
TPhiVuNT2ZAkM4fyMkcuQEpMsMmy/b/XO7rOioEToBzEKBrB/r+az0zHW7kytE1o
BTTNeJSPR4VdM4z9493O6x/N53ZIxrn8EkoyZE3TqGcmabQj8qXgs6HkJVLofZ0d
LSR9afEoiMQTkuLTzsHDCGKe3fRiB3eWmO/jNP1eA6zC28ShbrrHGX0iSIJCeW8N
Rth9hAbWpal9/F3btE4Iypnx5TFZul1izOP0tHfo4qC0kpTShM1vXVWRiU6+XDCx
sq8cdwwzBkY562i4ntB/ryCQfu4CKknm4keEZX3MLC8TErLxNFmhhmjnMZ2AYfKc
b2CF2Bb+rcGpL4uvrFPo9illEdlQd5OEGqXa15oMToQBtA21LTvpWT0mwLNkkd5/
h6jvNZL79j0/G8oiCX2AFUjoVwwsoa3Ry5uZaevJtdQTMeW+9KoSoIesCR1CL1gG
5nbNkcLV5oyhVLjFJHxB/2SbdFnUnHH+FRMKuNo2il6hB7BLnAmxrlAeZxyxV2d8
nhC2PBzhKtID9/m9oa4p1GODwR/3Wjj6AcyaLyryZeXyJMThc6RzaqC00UG++jhl
jCMN/q8BXW0lXJ4Fj/aiOKSF/MMe9RYeRf2b78KTJlAoNUlUkZwWuQqzE8ihMRyL
07lb16FjLhopWukMITZlnWRaPYsAMQ/7Gn0kdToDPr9uQLhDgZfc2HNeIUd1kcCn
RJNcx/HM61IjKS3VDXgaS9hQvwRALVaSMOYXr89G+G2EnWNTFTTENryZijS1d9U0
CCnhLhA/K6Vt00VSEOHHN6qwzGTLLj5GRIs8FV2THYv2Ny13DgpBEBAT4ETe47mN
6WvJ70pnerXwS5f2fJmXzNXvQeHXQiomYPNF2MTY4dJNwC0GNz+QiRpV4Gr5pBTj
3lITWJYU6GMwTXhH+vAF4aQQftcQ81xe58as49Lu5EmujG6b3rzE8Qp4Fq+7v2qT
Y2/C7p547bPIw4VfnxPxwzR3LkoQxsfb37Jh8Jz7qIH36YSpLzFFk8YQEWlqeWp4
t5F/rC1G9QHSBV3SkEW24b7xDKi2X6RLQgQH8qRgaTRRtzvHatZXsYavzw7VdQSd
jZXuxj7mdf7SBw/K1YkiUsg4PxhqMpgU/lNiftET9wNpO30vyfEk+WA+ymKHcKYo
0K6upXvN74zljZ2kR2CCZq5Z+qvODMwWo95mgwlTAndgC4mY0neXgapdENAoliNV
f9w/y7Dwx+5dkPVozwxABLEunzb9FyNUQwWuHrWmzwyRzVqNHaJXJasWmFlDDVSA
cOLZJ8mvvulqnQyJ7uZom0DzwFrNunaWExcLeW6mZxQTChYXTA3G5bMiwQTtohYw
oOlpoJEjIYTFPcvtkHjnDXux0m1io9UIA1yNubdSWa4i2jESRvMYMew8dvEKonjF
voG35YGDWp7kHDYxhyqFqMwUjNyPHJFXfdnhLiTHOlj1B7KZuLOGeDf0M9rvFrco
Ze/YAkH2fD1lzfqHtvqT05gd3HKDn6zDUuuK97pWQ/hgMy/t9KF/7upK9uil34CF
kvpWO/VKvHbfLqvwEEPe7DG8kOMcRFTCJ/b00OrSmXR6+aqOY/Omh5BbDPQte42v
+utZkeujEmq9QAcfd77yjMGe5ZyGXspkPzKqEQ6xyMKFXJe1K50/0noMw35hDrao
UX0aqMmGB9DILVciH8ARTdz3Z6pnsaBQF7wBqvwg/f7wbDJBJGnX/9k3R9HuyAGE
dwpdoSG57nHuBz0D5k6yPU3VLsfGJAoNL3NUxmR6bDD4e9KpvLAppxJ/dt7RfDCi
2fJE3CqjTNqFTrl0whFFqPaCya+Ea4+Iw58WXHn8uwZXVBqacGq2NID9IsDsHuq7
5fRIyJwbFVdn8rjc8Oa04C7UnnLF2X+G3ODFSueChqoDCa5364kSJhixEIQUrWrJ
D3WUHMifavpIk39xR5N1+7txD14qtBfP1N52c/2WZ2yFmeHf+SbZt/RxLRAd89l/
zfX/xHBBelYE862Vdkfb4I0pUqZDMXb45066028KpZ0++Bps7ZsFe6tw+5o30SiL
mtxS7BVz0ZhuxEphzTXmbz2Liy7e7A27M24RyNjySl6h/4bM6OT1D21aHkPS5g7t
ihS7NVtpjifD4SXJ/YA1DUTJm6F0h/dBPR7xPhC2fJRYGDUPyGDmlnxaGhwoIkMg
8NpdP4oRKZ/RXQg2fj13qu37l4rbkm5L/L+Y+F8UU5rruhkzvksevtoR3aPQ2Hxn
s5U106Zkt3NvbpkkKvHJF0Wj94iNj04dzEQ/ILBxCDBuU7JbnOMl5oo1B5jO8npV
eFKLQE5as720RVmwFjze+8xfBbIcLvvH2NhpXe/uciw24ZMzrap8G00trj+8QQAC
8mesoQWl95euFTauOcjfykv1qj17OV+W3jWXlmxzASIBUfpYpookzzd9QUMSa3K7
ovmjM9+N1zDWRtdS+EW7tWG8f5PF5zuSZCk5xgiP+08Jj5JmlyVtq4S8/NjRRYEs
2rPqalYWtLsdeN/pgr/tPLeppKEXHPjuFgaAFdoXE8+r0yIraSeSNr31YibNjG7o
OOvW5RQHTU6UbYu9H5iTbJNRf7Kl3Q+LfhtAODt6+KPJW6tgiiKVSlIVu7cVIa4f
yeYaXwOy6hrM/U3j4DCEkm5iN7RFHlNrZ52lofCKt1VSmUlZ2B1XmLUABwumOeHI
AL6xr2Sk+99F0ULNa3bMqaY10h1KFTA4ejt3yQia0K+FDHKEM/X+KzPZSw4DN5a8
cLAMW26YRGWyfRthrLYT0WJWSwYtHyuDrzZu/ZqIXJXc6+oCLoI8dpZgOwZ8OBDv
0iAKrLwWOv4dAbYgrIaG8iwCTh6HngSN1rKJJip2ooCHkcsuKc70l0x8rhEc4YC+
D3sacp7YxNmsKbg12s7v3i5G8rKoYzNh+6FARoTyL3KeWA9j6bCDkSHSFxE3qTFB
2Zw/6f6VSw6tfUgVykYMR7BLNEGeVOXM2dYXLSjoQGLhYBHAAC7F+ZKhiNtU2PZt
E4/ZJB4EeN2XlpO9OJHChHfwkN9sIluQEzgagKNxb5WjJylnsUwc1Dt22b99iBwm
X1s3iGein8mHqdbX/KCR+DJbw4dAUTLT5UXV6Bfc21XgeKaEPxIn+SYW4ZeDPr50
EOVNmLiwEO0/tozMlZFKL/lzR/vusOLuQiEMoiAJpAr75rr0tGskGJZ+/WJM7cBO
WiOZKBYbWL9BjtiHe6MnP57UEpCYippbLuBmwLAhyn/1Pthln/qTGvK4mvwcH9XO
boUjPABJk6FqliZeN+HZOxqeUcOJB6kkqZmKtXdgoDa0rk9+bOk50B4lpCHC8tmG
L7U7bWR785b6EoRRY5hoN5x30RhUI0XVd4//w58kGY8wYJvenJ2TTbnpTo03CLfF
Iym5p2S8yk5rU7oluPNTM/TpbgkDn/Rla9J1ToAP1Dba6pb29nk0HBasKI5VcFFw
sPihDQA82YkTqYHb4m6bFw7a9sOIbZoFUt51nWPoXCeW5YvL5bRw1QiyxeznbZl+
o1fBbQUmovsYpP75Jfp87+UAnqbglyAxfe8rdQeaALjzDbM0z2PdGVUbEVTB89tl
Hs3WfRz/FHQtkMs0/jH+TB+pXu7P539BUobJ7RsofXMyt2xd8Kaeb96HxH6BE1nH
NRKqzhP7k3mpBFeUXrG5zLvF9DBkIrcto652hVvB0l0u2E0P5KvNpYbdEaG84ghJ
BhMUXbWVBUjivTtEf4bKxCg4la5zkXWkjjI+6y9HiecMPJ562qwNqSao0cPQTVIp
X0/IeNZUyBWnCYjJLYtcfujdfN6QIzfH23+uPXUCJY8QaXJ63oJKEI06X7g4wHoA
7z+4fU8EDwt5JENUR/FzFMojo17ExSAw3rO9mpPO6vmDnbhRcsUm1xFFpKIwvNVB
2+SJc4r8lmS6C+8+zACfb3ol6ISI81k39t0JtDm/7Jiwjz4ZeyO++z/4CDmIJ9LZ
UxyJe5BD6P6xbmfnWyQ85gIYX1Gb4rYKaQqCrM65d1B5gXrsf9Kxxil0wP1d4kTB
Xk8XCgaRYdTZXMYgE5s+7IiuH8zMgZ6Hs2QctnoKiFdesrQqjLlhd7aAvz3xbkEQ
Ks7MKSCXtlF+CXJ5NJm/PA76Ug07qI5OQEEOJCMBH8G6f8UvxTNQxMvX7S2PfWcJ
5hZM7nUDz2HaCm+YTcLCIUlPg6Awe5CZXPjO9/ZFi7Z41nIN4sMsb9eHv5I3Ggz9
X7bzDKA9FSiCfqaUawAksce0CJaPflsK09Ojp+nT0b81n4KkpXDJz31FLBL8IlbK
+JXt0X22GDnf9g8qrsqGkpHl/1xLLVnDshNtUzDA0hp4bbs0QvmR0ErtPzb5wcJV
tHeTivg4sQf+BAg4NS0MYhlBiNA2Mk3Vqa2VIC3xCkZxmvbo1vP2OitLMSPuHrts
4brIvcDRc9TIH+4i5fDWfBdibDP5U+PMlUDK8thcGDHBIR77LgtWtw9BsVnmFjDk
qxEnPSDMr7/Mzq/bgQM0ZbgpjPwRYl9MTN7mShlVR79CR9/avj9UfbUCDVPGzA1i
0LwD536rAp6wc9kiCWGGUgiaNbonejGn/dibTi9kz9vFLd2Nus1CSvFIa0x99jr8
3K/yg+aQyECjYnEUwK7hIlN/PGAdWRrzP6tRPYIz6v4CFYmzV2lhMQ5ec4i/Ynw2
GBE183p0k+fviPpRqJLgnrQIbq7plr8B/gFkbV2jhnk2l/+P+bxgiRC8vDbdHlvs
2Jyk/tuDp0dQlW6xDuTkLw7L/Zhmgiv2nqvD/rGMYwx2QhkFAxw3lQiexIEeD3AU
u6K2DPPYtSRWn8pOs0KqcqOq1aDdboAabXMB4IZTL8M8ueSb+taVDp/hUuGCow3s
x6RtWLWP3AER8nVagwPfGhioEcjq+InVKo+laDtCy1L9TTmj1tYuZr4BeT/MIpMZ
8Qkno5Ekygb7IiHsYvxZGNWil5zoS/C7ce1wWCaKKKET/14AmwgUn94Mt8E/NYbb
vGifGE7ZP3843yEFdbTnhIOQuKmBCtpDbp0b8xt8jCUVfQGf1ELD7mStPiuypCRc
Fz024JRCJhurggP/wFQw4o3LMceddl6YKVg66OgYDsjUIzPxlkv6/aMFJboQY5kp
NoooCjVyNVqPyBOVp6uzc2XZGIddlEh2Dli26Adk1rIHby5WcI5max/+ux4rA/Cv
jUSHnflHunvoxxKj/GFJsJF29436NAfm72/MgqhrLWwFwlu9G4s5AaWpGUKBzjWk
KCKDAct89Gc+TaBdhMp5H5dKOzE+my5HODNadjvBL95+1vk1tTdTspjIjvL0oSlQ
yDrUZzdK3TS22ULndVqxlqj/K2kh+1aawsuQmNP1pQ9VgCl5QrY9Hl7tqpPPgwDF
xfmnwBcYhzbleFGIImESX9LT9MKTXP0GWQXgh8sm5YWt+3JO7/Un0ocRpeqV2/5n
DCP5k9G30B1ab5jcywSeBw==
`pragma protect end_protected
