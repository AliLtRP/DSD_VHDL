// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:39:00 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
P3yt38c1oL1Le8/+BMfgzBM696qZsDLpnNX1X8kFT7Z2lkRxbv8H4Usscq+eK/L8
rg09vs41/LOPq0BVaRGMN0geEAht7EBXL+2zrp8N/Mh6au/iJDn0pvLBTmyu3ujI
v0ZkR24UcAcGY2u3Cyd+zHqpSdLkGjgqnwCzv71rC4g=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 19152)
tTLK+9gVScZXNK0x+ydZz7rEe7ttvkY3cMFow38r/UZHQPYDki24TDkmhS4Wl1LP
C0indpNNtqgwyWxWVf4Wb1bR2rOAjpnKOe5US7/6cNJT+wvPyLFuUU0FxrdNarVu
DiUyjlo6CIYlmztvfw8cKHSdq41A+TcYdxgqKcLhh5ywMJpr2xadJk7NiTw19DvN
iW3h3YetftAIwpLouqKRW6F0ptQ3nVgzLi61zRxZKkj8vfoAlceJLBAK8Q2GAWVM
1v/fzkL1wh8qgFWLnG37wb2nQajTrWDuTgPwQqX8ENSncmTXgn7ZjMsWu/OK0FqR
KIcQ4r3CeBbaQGeHvMzAPHmjqrSRkhCG7A++YtGUIjs9Bo1LlXG+N2KR9zEk5Lms
y3+fb9pxj+yxdfTNzSRpxtf/Dt2565DMDIsrfbmrLCRAf3nANCs5xCnMfL94WniO
RT6DWn8Wz3LAYch83Gr3UnsNhWurCsr6poZDWojQItghwMn46f/F1QvoXRwCLIhY
wXioBAbBBhW/bg8mhELqCGM8k/FFIYBXgV2izZ/E2Abr+TAJyLIzdNO/2iESpKki
kc+ficxuByfEAFpFPHwW4WGS8uwhU/S94nN3vAPlxRLLku1+R3NITj1EBJxR4Amk
nNkjpV5fSt35G5uZrATpY7H54Dw3BPwAcnTqw7EPH2IYAuztQKnmDHFGN8+AYDsg
0aohPuFEPDE3704owSrNwcHWsS3ZF8B9enB8CKgAL+ZVVKv7I95bqOSi9PDDj6Xn
1LQvLuH5HuKQCkEFdUEA88ozXsNvtpgG+kfJGN58nM3MBWFiry6nVup9IBnQiRHC
Ux9oqyMB1T1YMYPbKiE80brZnFmeTikf7iuDfZkzLxBWf68gewAZDNek28L9h8/8
MLjlsx4o9Qv/xpw6IWokT+ueDno4LcrL7Lq3X4xYOWONKnE9a0NvsKxlqut05ZaH
3Txr5ASSDabcFJEFrWawB/jj3BIdZcza6Cp3zbed6ylfH5uOVsGMmaZYDAJ+w5xq
yaLTan60S7UW+qS25qyy6IXokhFdF5bqmYsabCLWFd9Fb4VHS3lTc0+MkjifX4sR
OuQKpOdYA9RMTEJvXVqUnwsCQ9bg2pBtfZBOgXGIiBE6MvCAW6an8+AuS2Km5DK4
+Rqf8YrgfQPO1PDWIw2sNB1tjYLxAsVhu+ccX6wQjK//zdB2PvNyFZ5p/UMAST5W
I3zHuSWD89+LxARuzyWX6+hPjR42Fhq6b/dkGTs8WTSVAaIszodrRatu3j9b1Qh7
YhPDHO1dETsL1dykcAF2s7fJ+KAUSyWsLGobx4rqMVRH296wFD+4ju+quc4k6wgT
b4jLRVwQlD881icvodw7MfG2cCDyusBXEybr99o7p9OjOFnz8FshxdnTHwlyYsN/
8Hnsi0PDQbIwneeCCNRFZ9UlPlsTi8AeISSbbhkjOcydFTh+R2HcECTWPa0u24s2
65wsowl70qwWsniI/+n+kdQW0BLComiYiru1UwecTLhpx44jl8EQmUeblcJcmnJZ
9NiVp0NYlyc6gaXzs0VO6yQjmcDRQPl4BbqCNUSSZoNtt5hGraO+UkalbbjptSsc
6qz7RymzuSQo828qf8oGK3xniL04Vj5jyre9IXt/AGRcX3QPNBRFM5f+reeUgwIf
w3KXucZ1Qq1YjFu0TJYrgTxfwJuizV8wVLB686iX/qiEdiA0tdnP4eiV/IQ0eb5Q
+e/k0ZgbTqzg0Y0iaBpG6O6t/Kfok/pZOQObdDQ17jpONAvhnW2Yf8TRGDMItMeC
IWbYUDlL+ei3sXoqMQF+7er/X9bqrqIJ663XvVa1mwOapjgJJMez6BPM0pVfVi7K
xuhO4X6Zd9da5BKpahpnfdE6rP2Lf6H/dKzg+ochkdqKGNhDOPIGEQtLGVmPDHly
kxZ8LQy0WqEd+oAw9T6l8pG2mk8QqnbdtMFylQooYCqiwQnE4MlTSKdhkxmysafB
1AuTN92B0nt9w4nCFIZs1AzwN3GraUuu0d50Yz8cMk3cPPsfmuM/UZxTzBOtg5g5
cziKC0tGgfkjNFMN+CK0Uo1ahXPSUJGxcfiLb4dWDu7zEqa59pxdA4LLkmheXffB
RbU2Rt3z/06I3eE3z6LO5+9i6a8gGXV2/O1oF9GPNnS296dLRuGxZ05aDwCkhNmC
TTBghSoDmu1ymFavHtCBnYvIGbmVm3WgY5jYzWVb01RAkTwkrGlzBZA+c52gU9g8
wij8lr1xPtMuaztK3Tg0dimjcTAodg+x/3zKScDCo4yMplTSR8PNcR8yxk0L5NHT
ID5NLPp4ouz6ez8G9/D0Qo4H8tZARg2JIZ9gaEMW5tTD9BY9zzpI4H/yG3FnPjHN
WGXJAAbXb+e1KDrhXOMKsbdzhn+xF02Y9vn+q4WF/hocTEelZWc1UBTvQMH++1Em
bkKL3mBjE4b+khuJvA/1r6e9zLrmUlhqamlF8/bn3T4EqyA4D3D3STo2DaIjhLYo
qyNmwB0n2qujS6LQ/7lIvIWjJYDuU7Eaob68XZ/UWQ1NWSPkuqb05oUgvr/OVasp
PV+LQz57jv9yPymQ03hXb9+jU8EBlLHT+qxUEsrp0dUwBMmadKtzCDO2VG2/8+vM
dTl5d+T2b7QFg4fiYsZJ6hH3eDfFkSiiNGlkWnBRTWBhOsWheHXwtW3w5L9ozQlg
MK15KRKcLIt1nn+ro/EGHG71g7Nm4YIyzRBPQR95Krtzk3jflYDCwQm/1LuG9ywq
lMZTJrJmKDmkB+PwoUZd/vgjOy/PPedWpSJtYeZ3k3F+iYm7yibdx1XgLUfzFs5+
RgrKVt4WnlKB4ltR6IkwIDP3ZYnY1f8d7k6kyXYmYUjR2lONtrgvKpgWVBwL/if2
kzI9ksxgXhwqMQxIxcgoruTWXcKb5EyjRVu6tC60UzXkskmCZhoA0a176wfRoZ4J
9MZ3lK+JVHT4vsWqdME4l2d60tZM59Yhmaym3mtQYJcd9qfyP7bvDzO7Cfh6CRcZ
sgoel+AwBH5QZWw6/lep/Y63k3rutF2Ah1L0oYymVgnagPonuUi1cDpCKVp5qAwj
aXbCPA6nXjp7f6bEd1MFasMKo04Y0ocyG934cXj7p9SCm4k8l94GYtN0A3Yr6MlB
xzRwkcHQ/3J1eNZU6a0rwS6cwqYg2/pRA+hpH0MCKMWfEz1k7U09VV/YkrlG4XRp
EDE+p8m3SbDFhF3lylOLDk2LRc8dglCrdds5LCm3IrHs0GOOMWQtAmHqc1QlIIRk
cxXqXYoBnVflz+nyhllBp3mHq63j0bzwoqzqjiBN+MEKXrekBXrbLF7EDbmOcvmo
u5FR6i33knqPW3IRHav090vWOQp0jP+XRbgqbpGFabMG4Xb6H0SzaXkzdFToaFzu
vlsmzXyiULm1sBdD36Whn8Jhmf22qd0EZw7T1pja4O6DFP0PowHIuS/zSFrox/aD
yWHDVmRZKOWcsN65w2/Y9s4VcrZeFvEbOFc94JU0t6/0lv5tB5Cx3M247UXh7lOI
2BzMyYwWvnMSfxEyB2INmHYyQVRBDVyLYzKR84/HNBnGqLQFV1QVw7lc5dahIs+5
+5rZkIgaFZBlmTBmQ36wi6c2MD3jBSRHJrz2QmQG+EalaHyHcVjl7k+RAlHizhe+
l7Ja0LSMWG1wAfKyVu2bcR35eF/i6HNW6xmsbJFwaqS2yo8AChhmVVU8IBWSCXOJ
BjxPCqBZIYiaEP1urv1GZtzv9CDA84HqOw7hZVNbukIL0agk2FNLvBHl87V/NGXE
InRrTIOxXcn9BCkxb5xP7OIcz/q9tEERMxbJ6NoXbLgH0N5H2INLa/eYO8BhBhL3
H5oYNWs4I7JsPe2EnmDcPVNPimSh5hBDm/bClm4Em7NULRknkzw/W1M42dgiWylo
TX2hpSmbjuOlPrClNRIThvjM5woODAmOlobUrVHzWSbz2myyJUZxJiG+FiVCKn1o
jc+8XTQv9fgGmcs6heNDq/cwXYPiitahMnwseS2uuhg+MSrSRJ3ebN6N3GoCJy21
BE5XhH1wP/XoO9hxlsxxYjK1WrRZHdQN1r+HEPfGgI/l1sMgyoWaW/7YZzYVkjGk
6liSG9JCX6b1kskrInxJ9544eUKRp2h4bCq9K/ZiY4wi7LELP/9cw1WHhfCG1GcU
u88xGbq1dXRAIRn8lbDMTblT3NubAn5O1/5VmJEBcmp/bOCpzMTsTtCI4BDG9rYm
McKJMwMLSMFqEYPoQP0SK+ffTCs1Q8bQ58bCVNNJXrayxVxUiGCrOWTH8hj93Ao1
Jkl2xjJhjD/DLGcr3ptNwCKAoTGGLvpQ/Be00z9vqjxbyNXR5L/NkU5rXm+KOOhX
AmqRIECVgbfJk9ecFuurgAN+JiEDgdrrPLilti11NoKspfjobsak6ElZbynWL6JL
DV/1kguL5qgY3HbMRr933l8lk2FBKUSfI3apIdJ4wJIa5osRB5/zDr1TpSSfvvl4
DBPoNyU2R2ygXmtUVUKZM+sm+av7pIUJjFqklIhNGx5oHRlQ3hrYBe+cBURYUkLB
8HS6cDxsV1MzjCZ4y7dk7VvNA5Jj9pq6DpRTMCZyGKnZf3EshM18MKs4onxBadmF
B4BpYtS8BYYg0FZI1/nzmQ4A0lURI1bYC07Z7qbbsKJ0kFW4TrvLlku31ngszsX7
e3agipuwDWheUVyFD/jsAbT13rqdOK9lIlkddztV5HHBW1mZf6D5GhFtPTiTzw0s
mopZ2+U+q9N//UkR4WwRst66GWvs+e1KYpJ1ghceyW1fkCXANzGg6eGLt/RD2gDB
va8x28LPkXsF05QzfFoxC33DfJ1fWO/3E4ayYhA/MSHukJQF/YZQPygi7/2rp6uS
eEFv3En0eksVDlEII+/6fZV++PZdAs2nAef6hDQX0h9ntrJQIiHrkOrzJThhdhjB
4FfFzZB1X8iJ1LCEhtqqugjz9FBSCEJfoXSw6WkJyTsIph6+yYFyeBboTYNaGUqG
kz1zbF9VsgOzA3Fd/Y+aeO2QJWsycu8Modj8QocpS/SygV0clnbbI/kZ2SDf/zxg
x2k3PkdWWjvJsFDck32CABOqhPo99O8kThvAXwllpake3fRYJZ6xnkOGxgY23tg2
mHP8x8uQGaD0eCiFGWCVTY81ZIGJJ1Ijslg9lYOvoiVxA/clX5vK0b5R5AbpO6eR
40D+KkpuICoqUlCTiA3n51CB0BGQc47QyYSKJSitj8S/A6KcuZzfoyrgNxAIAOJx
Dg0ksk2iJ/zhPBGmQs+2iRIDsKMU+fUwQ1D1T4grz6fCfSfAN913ANdSoIzkFOnU
3/HWIwfuLLIw503y7aiAIbAzhDZ7gEyox+wHiGLJ/cSbV/UVZdJM6V6MC9G5+MrQ
ZkDBKnRJq3K3r9GdBE8bWJDhZ5yOit69YHWhJ+kAa0wl6MU0yFpxjRJwRgBCDn+g
OkAluFOLe6fk2kA8zqk3gfJNd8bPtCsCs2Bzz3+beOhNXBuVSnpgpYMrZgwTPiwE
OyYauPmLqBWXQTvt0k7desV5RvUD+G8b1SnOM1+YfOTZzzQuwKVe/DhDTm5KwU89
0u5/kja6ASdlBNmfJ66wUNQzoW6vD9zgL/FSuY6X9ulGKPukpL7nxxhNfpKWXB5b
iOXmBQjBZise4z4tgW8xn3edkLmaAPcSbR7svh4Cb8rFYu1grhhMxog9C3DODUYH
AbELaC+9SA/nuj4n8ecPN7WzvMAXvJcvieX5SjtD0rGb9dvZOctC1UB+ZKyYF0xz
0bfmaWXHkPjdewILJ81lRq65ROebUB19MXgIIvXLR5CB8vFnt9nJVaumBkf+CeF8
I3QYB7V1T9boPwfKnOf6c2byHR13FCIStV+oLSSyaf/9LhsCch/cF/2cbVzufE1b
TtfqfiuNgMEpzMvynwTSxiBFlZVQFAx1U/yRFxMQGMlzuizuDG07qBnGnyIanRRT
3ZFnqrbdRbeDvLSSKei/LrB6c23+TWgmpi9gOLb1IYm/adrt4glNneitA8jzeGom
lrBD+G9/026gp+B2P1SFfBB+IWDKjdGIkrB8ga5dLioDjRgAWTKK1baQxzUq7Xe2
IPrisLuOsAxxbP9WGzXrNf9hXr5NKrc6baTe9Y7Rjhp0jwnyzrkbXIKIz/Wq9MvK
fkYnNMlMg8/FYtYayNmM+n9b3e7V7kuxib0M6rurDJEXM3K6yU9jGp1oxhE2YFxa
ldoALfsBCzt3prGtZLwk9keTwXnARZSwG4NA+WAbHIMEe2TA8u3VrwxGRQaPLGi2
2SHx5VIqjCHeMTsS6Y2pAgFwU0Z/wt/TJEBjo7sf49LH4U31pLIe6CD68lx0QiGa
D3TFfj2eBdImTwo/tY5N31hdHQCUYhZlrkbjrHGhiuOhftx89bW50Z0B5bc2rmyL
Cbgfhtp4XkRbFhQyfvzzSMkyAjBcOOW/6DXMm+Bqm7lxaD3VzyJgOOZ5c6OsZ54+
ihgQDIdOxXmBrO36zS6ALwKNWqSIgZk/QP+A8oVayyfq7d64mDy79FyzI1A9wPsr
tW2RLM5CX2bCRl7YQLbFBuvr4VLgFdszZYqyys+opxb7+Mp8mjaxFDn/7waxl6tz
5uvZ9Ve1VKJujW0c9GWDbue1WL9Om0c3UIxmg/mtNvlkO789PheSlYslA/HibQFB
jd1Gvdws9svi0UKDzsUO+N7nmL8A+3qVC8mgpBvtE2oN0UEXAoOsxld4yrlkJ/GT
8Lc5fDaElywtS2dxCGMXAGoY6heb0o9umry6gtRNTfTxSQkC4ywmoiIotTSoRgoR
fzWFKy3ddxspYG0dl9w8wwMsFBvErPEqV8VTtVKZJ+Gzy7m2nTzohihIRsS3wZVr
dccungEWXWli5Xha4oYgODEXy8dS/eo2qnWCUYPqrJVIQ4lhfpTa3NQpzht05203
qIwb8PVeRJp+CAgV1CZJlAeePirE0gtu5iiQMamRqUlwb00Fo4TdVB6bxYkhiKHy
I7YQgEXxvNU6B0WIn/6VGnhiBWrKWLoZwntcpE4Iu/JYhv+5MOMX+0aSvUAziSrp
AyzeMpIlowRKjNfra5z1+w9Q7wvE80Y0JHiiafM0Q1+xoGZhA70VoJTQH2NjsuM4
OzSC1f+qx917qY0lXyKRShCHBKtrxHayqOEa/qEvdjqn2g3Hk2KZrun4R9jhXpgY
tDNSboe7HpukjvQO73DLZqKz28bvPLLoGeCn1XZXlkrqyLpg1nxQhbIIsOmF/45o
2NVi8qH+sbD3igF0AKFYuyx9CgPJSVvtHP3I2Oxxr4WCr/obWj+5LwJaKak00gcj
nsoZxjAxf0wqVtE3VMPqnWNCN2xtJBb4X5bfyEjGWyXVNy1LrKSD2Un+wXDEzEfL
fhmeWu/RZFQ6jOWHwgHk0HKxowLpKegQxr+PT4fhZyxFIEwng8XxAR0rXBpxn9dc
S0Q61v31NeDT/yR09cMhO70i2+dsYhv6DGaXRUWrZwbQPUvVeDXTP0WDDogMmDl2
Y0BGck7bExM/BvCGTNGa5tt6AcYAEGSLUl2RYmwjA6XmoQOw17RefY9PoJAAkWgN
keuhBKlqtneqjjs0v3Mgq8pKPUFA+PTRCjk5Kh2k4BUbFNGtw0eJnFVla2b5gKNj
NkBP18RbaI5llMk0Hmb6tB+V3WzG5uirtGtepfxcTMvBnR7vza9NWnMQf4smxdNM
6tKctNibtKCzBcMgRib2+kwthjUOyG4+Lb56u6OjOJmKLsKnKHinn88EqR8GJg8a
S+od/RzRwYO+ZQjxvamZhnoc4yQVUhbfft52qnVkDnHV2JIiezp3+J4rcoHx2zDl
Cb2Ezu6SvDrN3zhGQq4ITuhwIzDozz5uSycHil7Rs3EcUBIaf5BvQyQ6N3oobdFr
iq/GTDCWGdXWQ78ZSvgdmXAlEjt5xJmtXfU8IejH2+xu5Lv8R9d4EL8PdaecIEsD
ShMt7yLUaBRv4pSYJKgvFTuQ5cHzY2vwapUkNl2D3Sg/1dLZJbu8hnhU7bXmfJtn
yZp5BRLrMnX5Lg07FCAdNwbG5061tMOysGTnTniaLVVFgq//8q7D74sqpuyxfGQw
nBBnwlX88tkI4lYv+MedeOoSSWIZNrXBEAll0LlnLHKPVJKlLMswa7v6Riig3cRJ
AlkDfgzp0mZXvslzxyN3SBT7ken0VU2vhd6BFDLyX7ocr2azFyefU7LqQ9XAsN6Q
j9isP6loUzIqKKSSBvwpGohPUmZIE34Yz9UH8y2isPK4zVRIz/KgN0SelJlUWST3
c4gADpDXq1qbLmXI86iWUXqMYOhHussW0IThQgAi+Fy4Urewob7K6BoLucqzjgKq
j1SE9S1pii3xJm6fB7shBd7eFrRNcWy1ILR4EDMiMyENZP0mgSEX3IG/NbOGMpa4
aRkIKUEqfgDaWLlLhg5e1GYCLbQK96MbFaN3wbdZyp6BmaDeCzXVM1gLMTX8DkNE
Q+7uHjc9viwElfzyNuJH6qgHQoJuBmAzbD2BelcKq98I0cZoo3t10noK+l8/Z+gN
hDVfDHI1gWfGYk2hx4CY9iSFS6IXdGvQUzhCxuMjto2on+qeAr+llIbBvmO4aPDn
xVCQ3RbCNYcSoGwBmBDqvP2GvlShM6Mysh7w8xjOftNndnOi4/X9vKH3fN5HCjJG
ZZzOZAC4vnEiD2D/jj+z3R7FCkdpa1SUPsMW9i26ldlCf2jhyVtBCEKigjxndgR6
qj2//R9Hb2h05SY4h/2vFu16NgikmpOk8qDsBHQO0hrjIcvpGy0UlqocHNha4xtV
Pyql+CUC8tNhA2EOrIL/7z6rsvdfcp93jJWaUlZ5226nimqof4nymNUm+2u8xOPQ
t0hok9rgBck8lia8pRkOW0iHXnaVWR+UHlKJ8iw7dh08GsB3mNS9orpn4JLBgbdA
SILT16J6xYse7Ec7TOfnGbbzyQ1GG6Kgc2pWORpqFUt1TApksEb9Jpt+2W70BrH5
TojMuLgYN17zKO9kaNHWJbWoPrnA60cp7uKLuHvFM6s4Js8cbdKa1jaOIlItjNHl
dr/bP+N1cFs5DbDiBH40I3CuLLDN/AB02cDtyEduor54lRP0QyXdmQJ4XmFp5lks
9wmQeXsEhUNP14HIM7pCAefEYHls4LJgg4N363lxs4JzZ7b3tP3+mH6WTUTJCLTb
k1Alu9JAC/Lh/as4jfBKvDQ8xTCRJCBijfJnmlzxIdO0hn7bUrabUnT7jPrVvSAB
G66j/ogzFoLsANjNRGi64y8tJFOIWyLwWdEFDVsBvYsrarcoKKnmjkQXvNBUaOoh
qA/aS3a9g+9zRHwC1NMu/Brt1FV/+hIyqXiG5XBABcQyRzQWVI5QjETTP/vdWiR+
NpxHIr7AnPMqDXXUZC/zzTcbShyWqfaN8+QQejNBtRBR9vmkdss0WUNztgT+JKWd
kbvFCOXcD4EF/uF7iWBI+CrDdlDrZBw8s4nmME3wGuUN3vrwQ5bTlQnv+UKnjYc0
8o9wue6F9lMHNkyz01mJuEdiu68E26F7rwj8nTlEMgcgeIkWrg1+K9sKSgipNmvN
LnD9lQe2ZaOfxBQigGOwKK+pghOxK2Cbts8j3+Jz+/7g1VEI/o4cmgMx9WoGIF7c
UCmIvjMQ4IgZjl7UBOx+WiO+peRLdNsWal+2hoGHrIGEjiOIU0GlaYcH/uzFbXjf
gMcJcXXMmXfYBKN1ZiBJqzG8s6dQbl/h1ekIeDtDBA9AGldH4HIQde/2tMjlPOIS
T4gU4hvCWoYBbPtcZtw5XbkonwsMb81qRUwpDSwp5IA4KSejZoQOdTJlwYm0y8vW
n4O4MldikmjlyFbjZqGjnwItOcgc3a8tLKJ0oxH1PWH6pf+lNm4VYtcOVUU9HmAB
2asJF9yIcG4K88RTsB2TkvCNELKjIaIMl5/ZMGl/zczNDkj2vnepyJKpa5quXaNo
Txc22PYOhDX79Mzh1vXPgFSD6oiuxJgy3+B8HtPwkOjnbqn/TxkJ6oB4egL9lVdP
5Pyt+xlyf7vYldoZJMdTkhffhjKe6EgYHnBe3u3Dov5EIV+S1S6AISCKMt/tR9GK
cwL5HuGiheExUv03rliPl+YdWh/9wu8Jz3o02PoSMBeRpE3GjFAbWmhCGCXxodG/
Lj1crjcMnYKCHCOue+E4UzJZ4HzLnlhMeVuqIdeYK45FIvx5PGgi/IuOR6pc/P3Q
DGGdsFBqMcit3v4gwjlJ7PIrL8RCoxGQ/DnmYteiPPD5ZjeyvlFrDZehCmJ4K6Qy
Gf0keHFLayKuFkW2xlP8eb1NEOD2AD40tCpnNx3LeVU22uwAegzGQskYOhzuni8A
I9BC4EinMw4SdTpIIpqXBndnWiv7p1XzkYWIo6j1M8DmPIaWGhUhsAvgCeo7grvx
/0GVEjOfMIPGhgBdEQrqA77EXhev0R+H+rhHep0HF0jSLiJmcsaXYj9glPGpoDaI
8Ko/m6M8t9CxkhYcV+Hv5QVyr+JIjPGBMr6CTUtaDJwO6dHV+ocAE1RqHr0Oui5N
WOSyfwnBQzjmkJ0IfyGydUEqzWarbQW4jFZ9loPhKh5vp5lzy/8uAQr/vEIobfSP
oZ53XyrMb/rAPRe5vrc97yoDavbFAQ9gzK7fqVT1ZCq9qfwdgPlcK2ruOoEp/r2D
bGitlsHf0rSTAOqeu3PWSwRoMsFlCrO2PnSO/qKnN0vbmsdqmtZYU1xOGEKWOSNk
bLVeB6uYUFW3hJPZFT47r5RM4BHFSEDnF2BCkt9MWAd0lezxdm8LAD8m+zkRyQHu
pNl5E8ZRa8jfZo18AY52+aCzdyko/EzpsjHvmo3xAIx0It7kV6CSbejxRWq18ErN
b8RbAXcjXJO6B5gkZkZt0+q8HkNFy+Sbm38rvS//ZTl5W1qRbRfySsqpA3hbJZp+
GSfxNrZU44AGNGvhazEADN/zsHCT+0zIfpF03eTmUiHDHBpTqUyKGyYSO68JxQI8
Q+2tOBAk+xB5SSa158IXWC1VJjjr+RHH+ny6GlxQNhne9QQGXoskcKcHa4UYK0Za
Pg0Nw17UvwTs29r6r5mXX/0rRFBa/vqO6X153Zxi00WtbkDThKHkQ2cVJfjuOLsi
khrwaAWI3kQG+ZRrXUu9GPt5mAjjXb/tpVLqFYDth98Red7e+xjVfIszpk+yLh/+
g2vOhzVh4UZqjrMptWchfWpE+ZulRno4S77czfPIb4jaGwYnAXYGD5nTB0+3Ktpm
dAjZyUpxkNxaU8wueaFXQgd3JZ27+gC8wFpVVQBc8QA4RUP4nxOoioBLKMEEqHxg
9x5IqYJHSFC6CZHwHnaSXmXk0rmQhBgCHleOERBciba2mdcZ/RyUc4F0st8gNQIM
3l79HjSH4qszho2agFRAsVC8mh04QCMF1pwBJKP2lYe22tfe+boMRzzdtr/TFCE8
L7kiXS0n7xTzSeCFIt0SbdsT3hDPzchQ7azrcnQFMwF4JgD8Htu6Pks645sOmDt+
xb2co44uJIWUwJ09lm2fQYwuLmnBp3wjhOezFvkSffZqhiLDjKxdMUQ9cCVZ5sYR
F09kyjE14vhHZZrX7KHeqZWn3Ezgqbv4ji2B/xOMxsaWNnTV25870KCIpfYozk8G
FQiqJq5q1fo+dqfc2vc/iunYLucE2k1OJvcAY5VI1MRAcqa9wR4Y3MfX90AHK2jt
JFdxT/HyI9sZDbZXfOdSaYWy/j1efX34QK3AzJrUfUDoaPmK7A1g4tnfx4fF762D
edfP0khTKSfJ54BZckqQ/4D30AF2LlAhnLZK/uCTZxdN1AOikJFt19UY+rNm+zZC
lXvVNyo67Rx+FGcxzPbHpCnj5ALR/5l1HCfwjspspovSr8wd1A2nW1gIzTVN9252
Ug9cRJZY5PKFJhOw28XHo3Sy9rKToQ3JTbvfbVmMf3qGXMdtl/otSuK6J/6tKSK3
e5Xz+D7X1lbiAkfen5IfikhLigFCVTg4PLYJb45kmZt8SqO+0Ey4UBojDl/cQC7d
JJA3izS0HoY5oI9a7r+lzNd02GjqSFvryQ7s01zpjyxkhkutiytLvFjXWghxw1Eq
4wt6E01ZjdchOiQ9Oek8ffE5jjAiQoZLR6JGmtvIbm4mrGw/i3zXWCE44MUspbU0
uJhaEx9UQgYGmNvVw+HyKBeR5x3DgtQL5tYuTezXZzcyIF//QNc997bTHgR2tC8q
ugrXHqru6Y4/LsKaWCsBCMrdfucbV8zQVhDUD20AjVl+ECkz+CfhAjP5Sx02ZcC/
rmiWwLu4whALFiivsaTlhSFeTVroWNFaygToTqClbcfdv8vS2PcLgA6AY9Hyhv1c
j7OPQ95neRSgaS5t8rN4DQWVxLi33Oj3JEMiXSLuPVGa8daNI9x2wRM1DhWNXvCM
9kIvGQM048T9CghWKERoqw8VcInE82vW7lLqoHQdl4KTeEzrjmIw07IHH/0K3JeC
cjmM+fAMtMuTj1jkpKWbBaxTpUTwfhXLL5LMMpjj3F9quYBh7ZD2eKcIXSCquqdy
HKQz9KCJCsnkNciEv8a6dHu2xjEitssaGfXLHtp5RhPAYyWPSIfowAzts6VNi8Cu
4FCFE2rbmD9Bx1VRRkaYkh8kyJiV/YbjKZkXUgyBKkMkQXCdEv2f+OxEEF3Tph24
X4qP0of9hoV9p8FFe7DWKguNCrV7CLvnwoTi31JQ4/ALuL6xyyn+0QYyU1oRFhdT
MGbp2aOVquLrE2KC7+Px0AP+wvb7C0L1yjAMSC/jrpO5JgJGt2xKkQ8rDSfxt0sh
KMBltgFGSxrzxF2AmLZBKD2KzOII6qDoidJf1LE0XaqnYE3yMd4k/K1rcvz0qXQ5
fENCmQkEV7Hp0p5iWzsywsBrmmSGTEq2AxFNkQY64bt+VKmuTOS4tRC684vFSEwj
z8YWUWNVufAECpGmLrJHiCjlVfy47ucR8piQx/NP3n8Pk/eQLHwkNR7NfhsJCPPB
ETM8h5qdwZNTjG/W3zMSmLH6kGEjvV4PlK6twrgGZhdBZTefrf/ZGVFp6MYq86lv
YddOvppoxtkuYfeyFhM6qlGGrCKrJGGO3c6SyFmmWVXWbWzS9EXC9VqWffkmA5EW
EdUkfaBCPItYV349cWjHmbnRbi1QU7jKJWLHPrF9i1YxV1qJlzS8K0pC7yZysLoS
VVlHZ2vwWfcvsMdH+ulw3+pMm4MbazfKSAhnmDvzJeP75C/0njK5SiYsGtuy44ax
LQVQUT2JGVsbOEM2QA8UG24MPnx1/sVha3vQyKvgzHzj91uwaqvuxYWQotBUHxdn
ZLHn9Qx5qlAa3oAIIlThue3lx6jRRrW5BplfW5rV5nWUIGR36EZJuRe5Q72mFknI
AvzoDJs4FValKwyVmFzQKePCxD9PbAuRbh0IGhwmyMIIKHNhefjdKOoKiMceBfTC
N8zLDg6kAnXLPUK7D8g2fxwI8tuvKk5pa+CYD57C+/hO7u+ksodFoiTex06vC+tk
8ZA5dHfC7VVoK+GRiof4aUwCTE8nlMrLTz8jw9Uhyny3yqnVOg2NpqjptcaIDgeL
Xoku0u9F9WVZH86xWJbQba6OR2/NPT4lqWWOng9pTGMS6dSqZafiBJdfLF4BGq8A
QRV7MYj0JqINgPw5oGXjnCT4dGjLPFjRz106g/OuQEVGv/zsUFeYAxew3g5BfoDS
9f9qJdl5yXDnITk/j5o49oGIxD+z0MH5Qcie/CWQZTXNMClZZSrc287vZo88KTdt
wNpYGJtVAr61zbKqrThKbuXIorefDm27Abj5RNspkdApupQ2sSzlxtuRv2WIXpG7
O9BCvcJQsk2FbEGqguyhTTdntCIeS04iZDfn8D+9RFCQemyfUjCjNfPDN5TrHvcx
2yk1Gq87EgVvJQduCYIExe8qptcoYESm3cHH1/0kMc5fRGQbSsQJ762NJLIvzuJ0
YgbcfODVsj2gf5OPoRyoLkGljOJwUBrFVeMjvyu9/5FnsGGJ4ZVUc66VRZA5B0gL
Fs7KzcBWv8IOFLJzZ50Pv2eiNrnodQPF5gN8LYM8qXkPY0DYAxRZ71CwAgqeFiuS
vC376NPxenlOUZYSRAGAXQuzIQ/U5nBEePYZvHE7G8ZRf+QtwfEfzY9qT4EshMzS
9gcyoSLCcXm17+OQu64Nczzm6lmzhdkQNNOGU6Srul7e6rw2e7vh+I00B6JXUAbz
oOiRzeKNGVGTzUjPighVgVA8v5H9IhV2K2/t0TnwrfB4RMY0xpVQRlwEVgyg/f0T
E4sK8R2PYf0aYLheQgTYpdOeqbqHLmn9LFz+C+IUOHkKBpaKifjQmz0PQN365j0S
w8D8+AO8YK0kOUOneeDJkq6EiCrFbdGUzPg/kXaz/PCxVM0Xjhkk2jyBXMqDlFrs
9YXdR/Sr+C06cRKj0/x0Poui3nWXz1xuQN+glMkM1RHN+pxm9zs/maZ7dkPUiZAE
BvnmbPIMKdjOgPQbiW+nx/u86SfIhz5rJoG+ABz/db1DDiN2jg095tFMlNAv87R7
2E8n7eORUEIXtIe6jdYx+Eo2rHfEOrEUGlT/QD+DR6YlkK9bMZHMyrow/b5R3dXh
Z8D01YoTaaTiW2rYBzZlt6ckJnHuaYhmAcCpWEEWkEfYdKofgGDCt0mpjRd6qHFB
GXUE/vEdo4XxNTUqeoXwZNe0gVVbSiKm0tU3Rn1YsbgWVmkb8M+8nWGWsXiAAsFO
VGtXZOKorYA/aNVfESDaSAoGSEO2uYcwTdyoi5A7b0y8l/d0nTkksQ82Vvsa9LOV
rex6Fyx0JNB9r/hvwLNy9LmG4FYOudtb2M4OG3t0lVb4+ZPTaSdkyAYwyB3chC3Y
ZoXKfyuJNYSyfpm+9k+ERe8Fl0RMPUstKzwtUvVesH5QkTmkK0MQy6Z7/uGw8hZQ
KaJEgNZJZh87eQj6XJyOjEu/gBIDL01fjniu76cIz4rlAQwGHbp3dEFXOm4uraib
nPF5on8Wb0Uee7TLZM1184y53HEPuI7mXK/ZUxIBAl3fjdJ3gvrG8dr9I92U/4bz
PNkWt8mg59x7jPIAIce9aV8BTojiyMcbnLmLyHoQPkD06pBQ8Xb0y2T8Bh1qkjKl
0411k4VqCUmlSUcXRFnU+yOcQuo+lelRBIE1pi/DJ3TxgAKTbbCznRKbwpuLQ6JX
vraVr4hVZw4WFi9+monoY0Vt8vO3KucCpieFcbz3fJ8vnqT56xS7oUqaUF788dbJ
UzQOY5MNwpSEgE5v5kjJqrZ9v4oga3KFNNy3h3fxkSAiB0H8srMvsIkwevjX821d
7tK5RqQR/OOUdQ1nci7fh7IVs224szryuvxmvIu8Ou/ZsoX5jChMKNCABwhmdyRT
etNXu2bS+6IFS7//vutR5qq4v5ngjz+TGc27W+1eD0ATkX5m9f4W9qyO2gcE8hpZ
EFK4r8zxyBRBXP+3n1I9nMLptutIaV0w8+b05T1DAvvniFbTHTfG9WV9jHHYYGCl
XB8bbivIuh0NRAVDYy38CvBs54XYm82pdgrtr5Q6RHrWeYO3W7m/V3QRIJ1XXJNN
K2OLiUGCYMGU0dbKRXEUGaQHrdkyuuPZnMKVDLd1nlVDN1daOApaq41RijAcXyja
r902MhPSRC+o6LhBJCgB+EW5+ffmzdCEWMK8zACqVUtFECtrCABTpoNvZWYwbbEA
8VpYoZxTo7AyVQh63Gm6b8ovWZw2mCDinAkI/ULrJhg9USn1P+Vcwq34esttYOCs
AXKzovl6X1pYIWUAdfm6Y2PaH0pA6Y4rp1vBz0WDvEUyr8GJ8wX1dNrNEfgy7xdB
IRacb9Hzl4QctdLvH1Rn2ZB1i1Vydy94oQGsOAnbgZiK67odeXthJJ1YRK9JPZPc
a31o0ZeUjkITiD0b2/xBQ+25Ob1xJ3sOlWmkupSwCu8Uo/OvhF1uSaWJykMSTI2i
K7dqcUIByeiUzekRZ9NtIpbLQ3/YT9IEZLJB3rd3F5thxTNaTHQgkWhRvdstp6c6
SNICg0CqA3Gxxl/bp+K5amMeBhd/xMox5aJwmX5zGPgXSWR0cFh5oq5YfKDaM2AV
ctYr5DQ/ZqP9BT16xm8n2XAYfaNrjFN28DDfgnTq+yZTVj7b0lRj+yqmQqiB+ZWc
7TWjiA8fbIp7ytbFHsDAeiM6gTZr4GsDeHeWBHBtGFZXVRSmLA+zd1queK/jaUuC
UaWGZaEkQQK6OJGbvd82I0TcQEzhhClURt2tdttsq7nZwwW0R2l48rlwnkZCZsRF
d9STFtSEMA/up4lbxDTi8Wbhjk49CXpuxBTNqM9K+FAqLWF7GLdkQbbqrAf6bF7/
rh7Fsdqgrl6b1+Fesl15b2e+3lM2ZVPFSHIZShN8AZlirphbmHVGVEEtECCqyKqK
cWHk7pcn373FPHwW0YxcFs8A8xPmg7bA+YY3djSz9zsZYwoizeJs0nZZ9OtwhB4/
8zzmXpKEOuUxjwraI/5HYFkhrtrcq7K4T5iDKhOfZqZCdjEnUO/WbiK5eKJgSk+C
btNMbI4n+YZiR1rRYXXJjSn2W8Rh6z4NEiC4mPlSetdZmpXTjrLKqSILEXs9oQXS
kbOGwQZHvzh1FgOLBLIUnSAfZIRXStkvJzaobacshQqBwn+DPNR2TJC36yNywrK0
oPgsvM3FSl9duIkt8TuqK/LN4IXcmoZmGvlpqxMtSoVJDgiNtK79fdHm+dz64pVC
uVl2duS5vHLRN2Zdgmh5DLCGW94d5zRm2U+kGjl+4d+5y2gSmbp6TKuQynU6V7Zl
h8QwDVqTy3IcRXiw0OfrHKdcQrCqe2Yh91vzQ3QOQndlui9CC9uVk8MqCIxULfFq
WTt27q4DtnEQganLBaNshrBa/3o9B2o6v1ULjgjqoPk0zAWioOumAFWvMH7w+Ztx
WjUQZQX+KrPWNUByj05wubm6xuMg4xwabD1eZXhrLV/yBhvJ0Z+tHyxFjWzmWw0k
8I2ko8Ja1eXHa1VcKhI8HT65vSz57GwntXu5MqnW7Ma5BrBEUG7vrFvuo/K+6tZ3
N7BT33KiGSZJe6mL6Z3Kw6fFTSGqzKtPmIKQTznscRW6njiKCdEkmhUk93WsyWv+
eSjgq5EoOAvS2PN/3oMCwFcAGbrh3QpgvDti6km71BN/vAkCknVPIiJrpeBTGZ4x
XBFPvdrKV/6T7VjKNBrdbv11k4GhnAaY61EZL/EzseidrKA/MpURPD5+nc2U7yuH
TZyozJgaRbYQ9LJm3qpniLykIJ8xQpLA4RnuRWrIwL6eGWS0eM9aTaf1Wt1hsluE
YYzm3FPPUlu3mtdKFV7/DhSbssSyoRUTUOzkxDuq9BGdfkTMPkw2TgeFOe0X7d/5
hKEM88K1R8I6NpFSwh3y5YUxy+Ps8WFSLg5xSppy4rEigR+n5kNZWjz6GEqrR50Z
s16jsTbImudLYSxXYeda2Px1B8dKXV3yu9yqQdQH0xKLUdNk9DPxJ0aBokH6toQd
xVJ0/M/ODnb93pG/F6r5DtKEq+D/JQDcCV16WYjnHuAAn8deS44UpVzlqvXp1yDb
A5q6hho6MFWB290RQf7OEKnF9EDNcDHv3pEPW85FCgPkry9OB5tJWEvxsQOSEd75
VUNS5+B2PPBJ1thcpootXQep7zfDCuU+1Dym2Scm3sh9RgNf8A+77G5IDqnnmd5N
kTk8gfIlMoPCNCZtB5Y5W7SwVskeDq8aWsgHKhEyVPfou6xgHOj3WN0ndu+ugkLX
k+qJhGb8jvrhu5Jvbl+wQOjpHSvQCTvUar+kUdPEQbdleB1+2jW+qvc6JJ+sGMYU
nAgjENlBzpcRHWD3uFRGrbFTje35QnGH9HPc1xhWxBb00PvTO+om/5RVm1tG4DKn
VBW5ETZI6xMV739PVn//pgv3Cn6SFfWSmUI+BUuoxN1UdQZ7rRiM5whLrm2TC0bk
plrtpFARDfKnBwdnt/S7Bx4ry2SZn9R4rjNhdDawPBzWCbWGPRdFi1aixZ4O6BjG
yNni7lfykEqQtsZke/M8HnR2h6o86rogtKnlhCKSyWnRqvL1X/yo1jTAv6sHWvMA
SsAlmIiAPiGRL99vtWRlSDVIwYd/OPIUTDDawMTYTju1+lv1ur8IABrga8oiNdGQ
f5G0KnPqPDTfH1c9EFwID9wbnDzBYbffbY62D9VPKlLiyMonbuyVZ5/lmxkc9Is6
bP48MVFFSK2uzsfo8ogQ9g6WelcHr1u4SeTg6M4sQJA0WKu7Lanr18Rcm0SpBMmA
K6QuJmsP+oZpD+0Lqi3BH1bgU1xVcywtC1o1Z4i71Xv87MSwy9Jy3LpZlFA6sgrg
+s4dXgRZ3/LlvjdTP1lGQvg2WMLZ1P/YQT3kzChY4eInRazxEuoWoJ3KzmFvFfLh
4HY3QlHz+thPH7n4gXxPdX3ALmIeiR2rvnE/EmxzgBAe6Svs8xgssbjLXauEdtw5
zTXVW0BiVhj/CYSfgpzH/fcZ8tTHI6VBs7z8X1YCZUz8W0WeDAEkMgEAfp2mplqt
Mtp1+GL6iWMTlIYWZgBr0lKo+3MQO29ieWcP69DPpDVJ78ldfISJLQowrBesAs5T
ca9A0uKCvtUazpuZBNeDSQaX48XZCMYc/MrQ93dvIXKNxt+dgPUQXVd+g9Juv5c/
a0DkmUHPJUEiQlEMe95N74uxNyOmBbmBSeSWnxjw5mz20cuZpFQ5zrz/fp2K4FDI
pXPsw7u3u+Cv8RmqyfmVNPll2Jzianwxz9wn7Fa8xresj2rut+XcpRwbsWEfvJGK
CeGZwzM00mIfaFAw4wj5v1RM2+tBM0ujyzUgBEEkvojLMCrGYmOi5dzBl4fTe+2v
S97noQtWw+aznLMnv9KGSy/NEdylmGCt8m72OpQjE3+Yrr4Zuc7rDUgFYfWRuKLd
XBuwYJyg02rBiFz8GyPmFYEcv2R9xgoFz/25obGxhB4T2X5gJZ6yTmbs9v12PT6I
MAzD7lRAxe8ZJDYM6m6Qb+Qnd/hPMmcHaR8dSDQEbVWLMqfu0OGBqq2anMoe31Sm
GNkYwAUQwA12yAvth2qK1XWktarg11hDavRWE63AwlQ70ql+M7gjHhWJ7GJwU4ft
aXyU6SBIF3/H0LePlTnRbGHcMzU6b2/S8YNWSWaRJ093bynKqABfq6hR/ltPDmuN
3u7g4Wb++Tif4/ZdTpPiKPZJF9KMqY937+uD8/zkgsQANurZLYV3pbvNRMnobLO9
XStopofhUwfJ56qYXfN8Hj+xDjCl6Ps2lutJaEfODGAWXrAnH6WX38eRWvOZkEb6
q7pdhWeUhpB8hnMFa57kAYUFZSY8eEK6PWuj+5cjvKxQfyw4VF+gZR3EOx9B871g
qdngdQfxiVaepKd9iHdosaj6CvNoG1yxfVRkBcedejET0cYtX/MQm+MwUyGqz1WX
IOcmKrFZeQxtYe70KPoYc/1RqlMHV4CFUwsid8g3S7OQbYchvK9PuLXFS5/YGsAj
FQCVFsoRzrUndz3ngpxjgY/941ONhIdXHrtwraF7zdUwwgSJ/fK1TqQwSHteOLX5
LIEFYl2KjZPK902a/B5h1mWhAU5N9g/qqT7tBNQ2IywjxoVzYn9auqzgs2IzOiQm
5CLh5g96HVTzerOwyYDfew94gxWyctdVKeZ3oM1sQ50U/LCr9F0WE8RIQ7BCVXcS
IUQIb/U0Iq++uBnEDqAlxRVSAid9oo0G9FI8sElvhlRIoWntb+HFl4PPiNoKSufe
qTv94q2z+G9y5Ripb126ATqmUlLKYBJlbTG1kxiKMJviW7cndfYPq/BWa8fnEJnz
21hyfusYlMvBS8z5qJyOfmtZy19BVcFdbqHpUanroceVfEcj8Tg0WrvGeL5j5+L7
paiYxqRotZGA9wST3nFFG1scmSIK24U2uT8phqzesSjVzBUupghJ3vk0Yw0nQ0LB
AF+LKdTInZKJL/5qCQarjSqqVeE7gkWZuQ4+vML/AfO0P5XUwFoesmsE2oLTvfQl
EZQxXqfCvFEnJOUxjNoGjz8nOI39NlbnaA1MVMNG4rHzWSubmpOdTAH3nyYwzRjR
YSQZI3DstbdtdLZqUAmmhY0Fjez4t2oEidhsZDAZHWqpwF0Itwm/vVS0uQ80JdDx
WgmAt800AcFVrQ5cOpEr8cd/0WyUK0PIEpU6ggf+wiIQyXIKMdJi4h0674/RPzVK
/XU7T/+nFsbJTVZDz7HsccHe+V0vq8XB6oR1yLMrCs2N058WiLHH0W9ncTOpArSp
chCUZanjpDFh91xGI71B45+77JXR2jfy3BXQOSWnImB0ZIqMLsDP6o0Rx1xwKRm2
XvlvvJmJu77LnKzJ8AfBL7QBuhTi80zy9Ya1y2hFVcdq5mkRNvooMqZluW0/YExz
BWIxqB/nI8NSUku7fmgA3DASzfkq7MNjCUtjO7vyXGy14boh3m9oPKTnGI5WMyXW
IeBP/Mx3IJYxIq1Sq/4d82x82w9my24BU8aARATkH39733ng4605Qp3sjoHJas3m
WIUCjVKBy6DOE+Ua63QtaV5hVGpe3Maa0n5+T7W8GwECIRTY/91JDhGg3sI9ASOZ
xTxo4SwOdIEmX1E9eJKP4K7aREhc1AeC89h9vbcPfO3lNhwmPTyqgBqH8toYOhih
XqMmO95eJR7OLyJhqTvr4fBkEWdYjZTxv0UqSMa1xDRNC7KPzGEmNVx0oPi9j/1G
E8J1Whb6NFmxBSSJvo6G8D+uVlB5dLPE8NfE/P6iAmqmv8f6m+bfGkLVHFJmq1QJ
5mAk/AVcY45RSuE4XZkLr4RXTm1dxmwt9LSkAnkSnAOyzVRtK2o2uIRZ3AglNDUm
20ZoMSiOO8kMDBwPvl53f8CHJMibJnTL20P0p3xkSzjqeJTbOM3fEBZh1ycNvqip
eHJeejesD8vPKLFoi4PhzbJO3/Zlk3hMCq6qpOqSAxffsP0guJEkyoBIlz+GbQNf
GfNSJq9UYyi/0rTMklIkV7ozzdu9U86dFoINSLDVTSUse7YiwSdATdmLPvSeUuC6
2FG47fdQiOZqC8K+IuVJcjsxeeSzTj+nSk9aDQd62KgTAAK8aghOhXbEKvGKLE+H
seTq3nqdZwnWyUBjwHcZ0Z0xrXBpn6rMHk+avIPoDV97m5vf4h2sxhKImnsReXjS
3bs7ODVLp3BOB21DGl/PbnYLjZiRXCxLjvaEeEW029fVJXotjM4NSo+qZ4sKyOXj
YB+Ck4VOWGf9oZ/glhUu11kWykBlEQwEZlcGg/PXH4OITyF1ePBFVdgBpOIdkkf+
Fq5ItX/J6OFVn/U0yM65KVN0SUUrGFDNOgHVLKx50xKuVRpaCKB554grm3tYWCfh
M6OzsTF8+RrLH+wpnwjV5KekZ0cfQKA08Pscr4OzSDRXnP2mUyagkxiUxDSFA5iN
85l9GQaidKKNuRpTQt3SUHimi5Ck4TYZBBuVEHlRFIqSvjMTIyWSGu6lsJqh4pX0
ohXSPyDyFyVidsXVTG7PQPqBNwJABwz+sSy02NvsR34S5/e1iW/NiBjMHFaBWhsp
Dm+lKpjzaxqslxILbM/7C/vOX/5wjhLtE2I07faQButDEKmy4wtkIzCkDRHx3U/e
fzMNAgpaoGzAq01J76gHdBTzOrPwyiwIyD7DS9Svf7VxRJVWvDARnHRhy4dvuDOx
8sVIOPnuPLqtWxWOGZlJFCeOw1yuerVAVOw5rlM0ZjsUqYNEnvz8HHnKEUu0jLc4
dDX/zXuJYi36jLB4jzzTykalkFJ63ICX47HzXMK6089t3IDNBj3VA223WXYjIGnv
nXQIc+vCVeJz7eT2RKvO5qX1cqbXuytc0+GDvrTb4NJ/UorCtLglWaLEHbllGggC
jiLDgn+QdL4DijFTewtAtCr+EhiFFnviqQOJ+1TplkqoRudK+NFx4M5slsR1s5jL
tbycBglDMMcn0ir+4yT0y66j4duTZv2dIpMscVJ+oOghejV9sQLBx2iNkyy5m7FC
KXiylU28/q3an2W2i0ukcHHtSthNEfbg5oOr7MNOAL6y8COu0ftxXy1ojKdHX+RL
R+VQywJU3klwhoJysNT7Ur0+awmIMihwNLoOJRvt+XLKHMEOl/9KICZ20acFTIYV
WY1+vC8UgjBjPTYhbqp5NC9Q0q6uO+/+rtD5RHt/wuUU9568QN4kxgyyZnyfu7kQ
YMeM91FJoRjkyT2D2PdC3Lo1ktqmUGdVYvoxKwq/lFXLRAAGjwoFKmlX8ncwHgNK
HV0p5WHvmJseTlPUh1Wsam7F9Mi0Dm5X1XnA4CFpaGe993MYYgPZPReHQc8LdUXH
zZdpUtax+CWLzIb4MGIuZ/Cg1qqzSZu0s6bc5cqogloAta5d6AeNspUeBz0z/iRm
jz/UzkiDYZYNM9hSFrjX51zUdQ5qz0UEmGZwLp+LBhpZg+CD4TR4jHDsLnfFCtUY
6jQOmeRRBZum+bGeg8omAmzzb53oSCKNKZRHWlsrMTyK9HOxbwHo9arWTV2n9AlH
L6J0Pa6vuKwHzoxZ+p9JpCVCsC5lInSeUxOKrVKnZPgoIXFdS8Jgec2/WniK1v5s
sWzVmoTHeyZmWP94Cg+618Ot4lqhjYAUkSe1lCR2xNWyrvfFIh9Q7wnn96bgbUMF
GQaplIkNwoo0CueFoezvlRIqXkbcJJxe+30lVvLGmQjczoHsQ2fkIfTAHl/kkbe4
vhr7ntrJGD6p/fJT0nn5EHGH4aLhdELSfrjJh9L6fmSW8pVSfTAxyqBLt2uWnGiA
fBBfQB5uE6F7GWMnc7FfNF6W4h4rnmHPP5xBGDtame+4xPvkUtYUvB50WcPWbva6
YG5+gOLy/MxCv2C16QW3LphS7fb5TbTAt95pQMgAJ/KQ3QTQzkoRIsyO3+GBRNlV
4a89GtD+fXSaJht5MjOozRJ8T1Xm0ErmmF1gNmBCoqc8VIEzT/2LOUI689gGGG3b
ZwwUOmm05WpF4ozx0CfYGt0TboLEOMdrQS1kgFb/XwzNJ9pdt8ICBq0ZfQxA4ORc
gwYl+RiuTcEYjUe2Fk3vlZyRi643G3skVzQCOx/MQNga8BnC7RDNvRaPdV1sa52D
voLZEKuZsSpmdj6L2zsLTYeiWhXAYIFlquknJb+c2ZXQU5m19T2gzpDfIMr8fJlN
PjmEfkKkwcJapZy0jKb/x40whW5vFaO8GsckJFZoMLDezEWLG9dVzJuhQCUhdT06
KMHWWOAv9JsyJguUek1vC5cDKcu/pq4WOpKdC51iGk4VmTTZXOYR4LWclzY3Jjq9
adPGwuqYpiF8XxnxA5hmarY92AcG3qrR+uTARTJd3ANvdHOG/GYZ+x6VPziaFeHC
jEfFXCm+LR85HhYDzzAIL55tBMPvJb+u8+FKjfKIklU3A+93mxq9Afoieb85wxEw
GAoOIw1zx7wSmakbuv0i7vMTu21jAoyLPy7nDLBS6wHg7fEOYAf24W8TTYHExrAN
jU38eWfp2n28XJJywcVH1fu+T8QyBWfTlHjJsvjy5hA2cB8OSEvIA2yttcLr9FB2
5JFe6YbtXh2z2Cfwy/TSjVhPJXU0e7jwfTu6PcklRJLy5qYbtmhAnuIMROsJMUbj
HeAkHY2Xp5k2RlZ10ZEZnpJ2FNUH8UIP4pIMs3033VpD2s/CtOTPmGnurYTGmyYQ
1NZg7LenVBW1Q9Ea9UUoK9LmbwyQ5jmRXXeBVhGROHUq1j42i1wqHc8JvWLBerPZ
mwZEVdE7GUHEt4NY06ufovr6gZw66OykLAQcFz8KDiaEtT/F+D6OzoCeMpSrkXcO
8WW5RpPbufJ7Q0+1xnCKpx2xJUoDPQhWyEshJUefjsLvY+n6MMbgqaGvNO7iiAmA
x9DqCsYpkzXOT2UoiD54uK+QmJdv1XK+dKp+1dh3Jpj8Nc2UJp9ZtoUQZqAfCKj5
vsZFD1n86U/oviV0LFooAQil3p6P/6zc75d2akqX0/JBnNvZqnaitI1FSfWqJrIg
2pVwflTKexdxSkQY0FKcv92MSCehCQY4XIxM3jJ8EcKOEPZkbT2jzOBsFHRhmue/
iEDN5sEBUpqqVqh1vnIq1Ymr1unpNIIVkCpR7qoWABpw3fQXTxc0sc6WAEvlxquZ
LoqLurBmTJM9uaJ9ydiQEfuFM3s8isFHcr3tbdOy/4DGwMOpE/QPLD6M6GHHH86R
AmkvCWFHi7nDsYVcGAzpn/GWQretBwr/1FIPTSKdjn/LCOksKERi5rYuvhKx2w/3
JIjkikXCGIqkctOsn9R5T/9Z4jVrGqQS43ulMZiDLOWhVsNvkmxvbRp80TbklgWA
GETs+wPMa+j4wKBVWLYZTpGE+EiKycjIXAISi08sGJwoUcODrUtx6jzVVaSJ3BGA
gzdDlqwcU9+sjGp516N1nHv4v8IRwy6FWb8yChakuk4W25U9J+0uGHCmahbcEkJZ
KirvQYU31joQzlh/9WL/Xb1Dny3FEO+rgKF3FYZoJbLO0SD2RpUbOsnTOuYdxUoA
bbUb9z2YhIq3wxvoDZjpaQ2qzRCfPAo5iBWZsckNKYv0+l+iNewbPL0wP0zEuKsr
OQxdyxgjKxF2Xn1y0mfB5w5P3oJMnrw+uc+31/Y0X0pcYSnk36TdZefK9JdA8hZ2
HduQvpLYvC82B9pCjxoGjqEMWNHIzaMo2SMRmVpEi3SO6BIOvP4M/4hWpRzuszhB
JkDLg4mzC2JPmwZZQ6Dhd6Y7Ot13kaBf28dyL5rz/nIQ8/aJsBG7tQG6SA0VpOZw
GtrPXUDnwZ+IjYNtl9YORP9ELHmQuaAYTQkT0pTJ9uB6XCC0jfxlPBJRa2TJM2Te
Nsh0DwernXXhAreOhcDqm0Q6GtI7Sb6bhfzTjkP1CA5qsZbfsBg9zgHpKwEx+Jt9
NF6Ly0A117dXA1+wPyUwI8HfNYIPLcbNprHZrJxRc8YUUbxIaN4a8AuVRGLwTWyk
aSGij/Y7HCS2iIhKjoPU2rsLGGBZP1Pz6GLj53UZZYNvznie1RiALD+rTkGFB/2M
qGlmeVtJtB5aNOtfebSAwC0c2ggWuLpQy/UV7WZiLrGo6REr4j04Hn8zTu5If2MT
DZIKxz/Ap+Ry/NONzdaUgwvzDmQCn8xFjshdLQf6mHvMJ2POyqbLeOKym6cmw9JJ
j762b/e8aQTFKqBJ9qexq+gEEPvMthflPI+gHC289gKBSvj59f3JnGSLVknlPTAQ
i/dVmMkIa+fH0D+0D+l2ZKj4tITnqhdDhsuHA+wfLrB5y6bg5MIZ8OYXnAjNK9Mp
a+pQ3wOsI/79+k6IEJ1/cgirS/JIgtOq8O7uniwPFxvRhp/xj+SwOA5IHQT27c4v
zsfIk2cDF1sJUWP7Vvbr8JxId+je8xZVrzZ2qsHOsRh5G6HHSDJPCdvULFMyXjSW
iepTwhvjR6LtFBYtOnX3cPewRzoI2X5zomQwP3eHo6ithOMAldD4Gz5erHDmUuM0
Ap6k7XrYui882mgknxb086RzClE3EanSDqG2V/PpxY18IlF+ZpchrOY063WIVoV5
hkC4UbUFuJRVgsNYT6pTUQYn7wdyU+2ELutrBwwX1SkCZQU3sU9l2Rxw73Ht58ny
81UtEUwi25zkuu3Hnzq7LaOZRIJakN3Z3zM0ik9mLaGflQcZiJpdYbRtsCmfvByG
`pragma protect end_protected
