// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:37:34 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
RDJ9gDa9XTJ+VkUW9zU//HZnXACnCsWHORs1+YHjfg8yIu60tpDEdMyp0q5GwfXC
NIUJ+12xQqQBdbMX75AQmScLk5yUmWoS8XRkmTq2f3hIL6r6unIifHlX+tQ9kyD6
v/QMDGSWtRhQSu7cq8NpOrIaLAhBGnrSTT5QD0FRAOs=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 25216)
0YtDo2vnZwnD6YynM3VpM5E7vDYqmYNUj3LA7L7LpiznML0Qex5T7bVI7Zt/9c/P
2BQdfxvkNoOKkeAt1fLgdqe8teDtdbD7z3CS6QTigqRlFiBWChTfrEY/k0GLzCG1
CsUyQ5nNCjd+sOxUMuVXhUIflAjNZME6HS7XWCpZ5OcJcRfVihuRTYhNJd592nca
hpFaM8LIEGj65VkRLEauv8lYrmYfM5lCcp4zVBjNURdNLLTIP1LnVj9d3Q0mD9ak
PT9C9fox0Mi180pasm3n6RaaW0pWmlCWJxIDW5Nace4aT1F83ZevSMwKC+T4Pjw3
Y5pcDOVksRp8+iX+OMaxACmOGPHIKr6fJ/aEZg1fphiCplcBTDu8vnM+K1CyhoPe
Hi08Pq0BKIVOc02VguedlN55cUa9JygrahSwQUlxivNS+U+4FgVDqaXEbVHeFR3c
Bjy5Wd4TSS3G9GVrXu5B+khYMVdeSSy0+ARhEevmj6H20lvM8QSoYWoxUqFbfzbD
i8sdXpp2zPUBcpqZcg6wmuCZi9lJ26a74PgKtMFm0yMXb05ZltXNwdXFCpQM/y6u
eJeeVaPVHw/PzoLhhfhgnNS9Yda0AKVJFtLCNZ3PChUuz1WHmJ6JRKzoan/LzG3i
O3iOo4U/3mKACeVSZcpvIuf8FIZwZ+Rc1HVO4Y4BJU7QUbpupXnNFvkSAtaezSSx
UG6MuVAeejoaa8lafof01ziIt//FmGB84HDOMfPDjfykHn7HAL6UXk89D/gIBxPQ
fIrDG20LjNq6Z+7aA3hAb1kCKqi7BVTiJe++PWAbROSuJIxSack0wlVe7iO1zl6h
yb4blg0ZtqdZqk0rLkXmxKr8c38uiBkWpYyOXaZArETbJfMbsnBnJqF18u2xOLQJ
dAfOlAOH1wtO/9AY/0RLM5aINmgPrRzmqAHQXDC2/afKtfadrwTV9q5eTsUAzvyK
nRpMHmW1Sa9vUa4TyJ6tgJ0d7pIiJMVQ9mlF9K7R4CAguE1GhNuKi7Wn5PGeeMHZ
sIXZ5/IR7HTt8EswZUnQXYqtmyLxGdifziDmGzoF9jcoFmwvZXE2FTMaPaMzji+d
xVP4RIf4Hvpeki5hgFGgWT1oORBFu6OhOoXX8QjiYLlpibS5rrZLT8wIBrfLKBEU
2tmyRfki0Cf6x/spzuy5BIvp9Vr2rYmJF/VeycYQV+cYwsNBE43oeUD3YWbEQ4Vd
Bn0WMOfwT6x6l1xA9OcWV9mu+lDNwFc/GaUSMdX3J5mu04tnbSFCX9UGTKK/W+tc
RIvx4cEHF0eONX80EwmphkICtql9TJw7hOv9chDNzxW/Dh004YT6O8DiO4tOmhQV
y1A3QQstVISyeZTFGiPsSYjFIfCvTeRfArlOg9nTjZ3I7x2FZPuvFevMPj6wMzLM
Pef9O7R5T+r7sHYfP0jGEeuVbFdegJLi6QG+6MGAsum969Pr/kgBZAHFRcNSt2dh
EQ9CEUe4hZRZOqmEhdwyj3L5i1Npv6l56ShDBTY4BXBa17/9KxuS5nkErNcM15JD
dubaplSzLF1JNOHsQkObiIxnc1KKvq+TMv7Or3c76HA8+8CnySrcxD6NX3taJT91
AXkwWAlhrwSUuyAFoG0Gi8293WjTbmflhWF1OsKGLxLFhSS6VLzhoKz4R4hcgct+
TGJFuhlp/yXcnRi8IqtQGWQtQM62/0MkW/ye/dpPrLlsN/ll3NXcudI2v3Dodpet
1lO92UhYWEwQj8f1PISD+9+7fL4dxab6wR99xT0TlaLxdFrMFB63B/a9LPFRrOpF
97gmuYgYYkEV5Dxg5MGJpp8xUkRTOp1KB54wBB1rGwHJE6jRmcmF13kbtJsHz/Uc
pB9y6h2YyXiInHxer83DarwMiuDO8UePR/2SaYxl4kfVqDGqOkSFTpjm8a2ncO5U
fuWe9+vVt/Q4++3lMt4e1/F0h+mHd7y9pr+ZlRB+r93ZEVcA5HU9lv7pjtASZksD
IXXWMyirkkBfFcszvv+7hs2FB7YU5YjDz5aAJlZMQoUlqvH4EDWwZV0+Y4CU8+9b
31W39PbONy3vQ43f7tgK2TfFAMPCJd7v+VKLZQveLQRsHIPNUekusC+ViAXwu8GT
jN4Rb0MjWZstbhTWCAgU5CbxvZg4d0nJt8ofqKuPEPhf1YmlWltj1KclgJ2Hec3G
ku3jeWqyDdQ92WJHjCPcCGQtZodgWkDRPRKdVjPAnZrZqp6sGM3MnGhAjeN7nGly
44Hsks3z7dZfHqMLOXR0A+hlsTukX4175mazh3BcUkM3193HDgRHqOwzF2C+wWFr
In5qJa2N0PPFXdEaRmM/naKHhVSG+VqTQyM0b0OirQ4hqcRm1AUjWCupHjdWyqXS
lO+pHTWRC0phCCw6VSC/TLGpIrtBD5F17XsRypZpzP4qv1DuBsUDihHP0OS4lPDj
TjUb0LVpLWSSV/KIeH1qAKZj9rXAaz3ykf1stK8dEhj33mmHOc+uBSIC9DlclrfK
cxxrOGVxE7kHIrqlY/6U4b3TFb+9McrmKinsCrH80xxvj5f/3UUvtbCH+2Vcu4IY
QgdZ0CuS4UQvhIYpio8O1iyC7N5+O0TifpIyQQ56EacZrUk14uEw1KFBqWqbtRFy
j6AWcTZAi6rxk35DkNtYVy2mcsVNd0YoEWRh+yrVPsJHAmQsgsgsQBvfCpnliHnS
8rnypT9yrzSinN/gu9QrjvY6hYchXp1u8YTuZelsAB2puROACvtxrSBXpWOeVW8g
bphcmwrPGJQNjSL25GwcLYuZVEmjZTjXhs063wWRgKRkWYSTNEIuDdxJcLmi4V7O
xAyQ7ss6BNAAC+Ja1q0yrEXxSaeejKfEiv4Nm5g7RVu24HThu7g0909YlRrXv+4g
bPVqj6KdfaptBossoW6wTv846pTQna5OZR6N7q8TXII3x6eEpLrzJTjaN89l4Eag
/0CxDzwbxwZMfPgnAFTZAPV4JoMpybGSZP9GGo7OgSuefoJJ0Fms3BOa3Pwv+Zbu
spsDAp1tQvgT69Yz6eiY8uagxX3j5/dIs4GxrhP7hgbzR3VLQNm0lBT/o5V8+YwY
1CY3IAtx3ANy8+z5Xhga4gFteCIEPe6SV4X90pAs9ltHy+TwTM0GnQkDh3933sTM
Yinz/1Dzgns68ngDUGELyycwR+rlXZLJhUx9OmPb5Z7qx0B2PTsKCaFiESwqg1dM
Ijb5QV1NAcsImqV0oS+tHdDXfBUV87R8rRD4pBpFkTXPFHInTSAMRCfdvH3e8C0d
4B6qTmEFWwD12xgchkiTYtYVqj+yiozsxfg1b93Td0uJdWWQ7DsUOnfV+pMsO8r7
i0LK+zPkoMT1gx8+f38+Hc+J18u0VFZBHh+zbYBy96yU2YwYoPRyvt16O8KI15P2
3qfB4VR0RhydTH0C2VbOYVfzfii4hpZ7ufOU96DKIaHzYlD/jmBPe6murFqO9Vl4
35cm8Z35kH9s1UWe0ZA7UbWx9lWV1vKjbez6jPqtwwK4JiqAX0R6Jlbkwl0PEWEy
hwYBZ5/6Qd9hGSkKbMhop6wBlPldLi5juca1jFuD1hL0yhOEs7Y8HskdvGEAj5M4
jHUy2oqc6aVPeTM1MTLpg+uCHy+ZAi3htlnZjms+pn3a92/vP+CEii9hjk9Jqvd1
bNB/FsSGY4z/jSIDdM5ZvVz8sShM/N+XN8Zzfe/OyB75Nk6FOOKWXB90DerlUUoT
mS3vhMc25SybP1DyVQSAtETSp/ZdNinEAGqH153WSYgBWKGohdUr8O1CPMLJ4oPW
UxZuxLPWsDXAOBMlnKcrEWTkwYuMdqTSuGzVu0F+/wNp+CiYlnLkN00yWHDOWwyQ
3j2axt+QGJOi06uqIeIx2171U7xyI4QptxCg/Ufn8nP3SB61n1PRn/pJLbxKgy55
CtB/iIuWB6hVWeLJDfJnDH2i2fcC498kmWZ+ewZC4STURbYMeNROq0mVWh5yebE/
phhjzQhQG1Eyc8XUGRLCp2jckEnVhCE3CWHDCWPIv4riCEbZ9UvII8ZYFL/WZvBK
Dukh4eeVI9BA/5dva7gLUXn/eD1SOGrgZMT1rVbDFYW/6LRMe58QRHvqCc0eEK6N
yGE54qsho/q+jOuahj1Wm7B2taX6rR5yDpHqZjJEm7iNU2X3pe3/a0M/YVGskMNX
OY+ghtk/lAw79hcor60k99HynTfYdjFZafD8KNeOzYhy2krKleFmm8qBv4oTIJnH
XUn75g41YpmJuNZw9M3Z05Q2XnGCfeWIUOruYQVfwZcOGbJ7tVKAq8KjUVvZJ99/
rv4fsRsxFnBqoRVDSYyz+vcyM6SzwxOj64oPjJX7wK75AkI2wlcEUr8jqnNpAu+p
K7oa88JcjkMXaz4u3M9QhBYhhaXzagGrdDgl2tsfcwgOzYlN6BhWK5+2HogS9VGZ
wCgJlFEXltouaTlfBBiYIaBrP43uQ0AvuJIwp1enAx8Bo2FcinvUwEXKLn6ASdxN
nttaoDkk2kiMT43drEltbT9woNw+KT+Vg/c8o2ezY+DtPk8ygjW7qz0wfGe78AXC
ouetA/c7K9nCuSZRHlO2houPPtEbaVx+lEktHbNwBzw0e+A4YsJ7KcJXmKNHGA/C
y14TPtIpvej6qrCrIgveVKNGCwPUHKnHEda3NOAn9xIsT8ZOBkSyw9/JiT8X5wJ/
gz9NEWef6CunejUBItTeyfLGCA3Nynlkjnyc6KBUDe26efK2QzJrh2CT8p2Oggxu
mHEvpBmYDesJIDt8SmkA2huJGWMt18DVCMqsJ9fg/yK2qmnrj3hxr9EcAYEywWWZ
gVU9Hgs/FFj/oCaCmvniPPh+S4qWy7CRn4HvZq6viOiJabYAkp8dXyYC/kNBz5OA
QFvY0lxesS1vjITVIlvXEq17Lg3Zk/xHkq7kB5Y+1FIAvDWPmNhImToHSrBzrLjG
+bW9yxjRa93XzNIvFZL78Kh8Fl1AuvPaHE+/MdJQa4hqoJxvPvGrggWLFP/G/6+c
n10B2WTcIkIQMRT4WYY54I+CSoCZ7T9vo8Oa5KvJjkK8UT+3d8PAwDz0FFo5xLhN
LSBOB77upZXuPYmyl8YJhGYDgMKnKQT8cuoQaaZ4YNwjchUsg6QAnuyPab1QfeYJ
0XhP//spzOMug7NuNkSiLZaGKaQBKpZmcO1Eek/rIQaCr7elDZpwYiTFKPnRKvxI
lfBhZYoTraAAuGZNhS/580oQQ4wG0kXRvO/biNgaf6ixk9yUgju6qADAJGe9vjM1
1dBczKWmsHXMFofYeEZ8J1QUzANaa42U48r1ggOMwXKnUmHORDeXhKPzbX9DEOz1
Ho2vQ35hKqdPzrjbHdK5lzbo76XvHDtgnyskQHmWTepUtljxOGSGmYJ2RWYIx8p8
Sw4mprqMPGIwvcEV/D8uq1V31qOCSaCJGjKdco1IsEYWXFpQ8HzZ8+Lq2XbE3U9P
0dJFoUxX/XD//piFnLDXWVluNSFbNJl13iXgSlJvw0/vBLsRVjl0Alq0v4YH8Sev
cl4n+fIvFLNzI4xw8PQGETtZQJlP2GajLy+u1jSpTcCW5hqRNz7+Ix1WhKT8vBpg
rOwJHT7nxlsIsxvItIaXSTMvsmj7qc/oBKio9SOZKwoP4aZkWEHHzCLkxPq/zt9a
38KJZaW82qXA6594lKaQ9qiGCd/6/0iAT/3uA1VvMq1EmlJ/fc7Y8jfd0IOi5pF0
RaUSbeJ6Dt2KXQEikctvaIt+iZq4dr7ZPP+pCEkOXwKdc88McLYj32vDifUy1+o4
RaJ4V62GGbjE94mdVFocc/oEIx6/ks+/eP/zPO0cQylz5DtnpEEa4rmDEtvNM7z4
VWoM72A7SOYouWkkRNaEvfrqOxiL/d/gAqi5g3qnoqiYxF6zswHRGvI4JPyccWGZ
0fNAs+Gjiym0n6GpJ5lmwoImNwS5Zm1/k+6b417peLBb+NcNyGwS5NfmDUI/NM2U
q0pc2ibhmhpxQvkH+HKy/JxJ6ssxNAq+2HXHBL02oTMWnBGJ962Kkff9R3ACyzdU
RKQ/lWw2PVFZA2ibuVJP8UA5emUNfQNep8gSeL2JIKvw3bInqKGtInz6ApXG/Cwi
f7RoCkp5qnzzda71Agf4DQ8OQq/YF3OfhpWKXY1VK3wtTzHPB8AbZLmeqrhlBLtj
BW4Y/lK0x1qlA0RXmBFmHZ1/LG4nYF5mA42+aRsuyGTii21Z4Nou1Iz3Xnmmfu4x
FWedQDfirSwL0WUqBxKk8R6xUJt4jOJ3UI16wukHhlEBJFJwnMyDdHCQbSY/Mbdg
J52hwB1SLSPGfVYE9xZOnhWyLaddGy2t1/pu7xU5R0xfD0PHFstXUhl1dEHrh3GT
0iAplhUzaM/wtWg+bVqKPxGmgCFkN1XvPpj5YjiR3sgCWBziUF4Z+ZK9FgPjcOxV
rLsLqf6bWs1pJeRdyy7DNJaiM1rm+lyRrqX+WpKWsYXU7J2NVPAYTmRFEhEgt2xY
WmbVV6x+PPrthWsr/NXC+t1cV9LL+x94+Z/vLYnQ+Ac0nZqChR5bFc7n8VEHfnMx
g8vS1+ofEdLUxm7IxUSlKU858Hue+L/xi0RZbfLqRxZzRppj8CNTjFymNm2xjzVl
Vu/YJmLPZvY5NUlPJ2hXTTcTnoXiIuRTkMtiA5qdA3jLQA1GKPExzyHMikizHMx2
iEfhSau2vcC//U6L6Fl9mxHmqYMpDQsfFvp9H0TZala1ZfUptAtNT3GkIfDVtkYN
gZuAzU1trDgyJ7N+APJJyCjgbfunws5Gv0IKwddbk8Rg7GIpmiBP54kQptO+6+oU
QnZs/yDsrtBctj4DkRs81V+DSuLAzvDTdj/KWYsugxjkyXwg2VJ0eaz8AICk47Kc
Vh70VqQV+hnZJOJJeqduUq0YiVVNYFtCslP37kXMZQEL8zW5qS2xDrJsFrFHqFMO
XwccRO4RugtxCVl6xv+9ZjgMAlLml9yZqWtvPcBTR0C4VjtYcX1bprNuXQBeEBDi
kYXxtNh+YAsMUD/FfAq89UDfjqwf8TkUj3QaCtI8jf/j5ZgwSNOwd/66u+iCYqqI
aPS9UcGeR6VIcTzOXUERuFQzxnXWTWQ3ql2jbieIvcs4eXvF6tieMxfbqKcWi+sP
wNREaky+IIY7f2J3SCkvh63Ti6i8eBaFQ1T3VgrfQwtVVg8zHovHVR2D09vo2d/o
o5qQQGZq4ZF4nmcUI7NEnVaPBOhiLxiflCRxjb9UfttfUjq9Vicslv5ENM3gs3CC
paiLfGTdO567lhJwaSudkwj8gHGRP/IiKU2//eh7ZLN4ln2vbxrrujIHJa/Kh40r
Ql7vRiEauZM1fKrDQnyx+BaWr1weH4rCGlWC+XvPPKf7nJqptdriQpgFoWdEjWei
v9ciS+2WwGDzzxDxpZ2mqcIK9nnwbocsf4xdeMAEiDuB77WQaZIAzSjnZwd3Gz61
I9vFqIdaIk2PgDEGaLyl6TpNb9+GM77X8hgD8uYwn1je3cgdX9NOFRNaPORPmXov
Z4Hun4CxqkVSmUASrgydXshuWWwsT9AO0SHpknWurnl1ynNeGwl3X00Dz7lE8y6H
6Vhf1uoK+7hym3ctK+R2PxHas3hbvM3DNG9q27dbUCWibA1f5+5zZn9fzw8IqnV5
EWrNFH+DnR0g2mTih8OfFur2TSr4Nh9JSVtsQPUdIangRqDT3wM4B5G7uHJJeKo0
nbC8qeQKwoUEYPXNnudSBrhtVNgkiYBTpgcz4TgpMPEvbE/4GlGv69nBCLJB/Kzo
D8m/Hbzw2pQ9UsXfcUWwKgTLInXWYTKGRdX3+6lPaoBSjlJkJiUbdhBGBUCcdFBB
K0bm4L5jHS7Jz/wclRSAwgtJ/bXFidAkLdY5LNeGPMJBY/EkvhtAtD3Q0lqaZqHo
OkpaTvgf7+KNElCSCM1WI+c92AnspUuOVCVCSPVE74VoKTHxUH+hD7Wg5ECvTylf
aH52v4V49uJ66LfVeUIUSCJg52RDVE3nZOSZVILAmEckiXhet/VrET+rlcVR2CH0
9gyezaepJa8qXS7ACRVjzy65G1b1KTU1cR/k5RmtYTpzC4eis6DjdgOY038zqvy6
suejtG106gHxvmi164MDjfWKpJw8nMC7oVkW1BHoU+m3G4tcyeVU1gSgq48cyH0/
TpDsgb+qDmRTnG5C8niHM+wIibx4BTQqRHL+FwH9T2aX3LfMB0D10VI6suUPtlOx
2k6u6FMX5nDmMQs+a3QXuXxF0DSm1ntYZhXuOc07TbCpBkiIhqKZRJRC1ArKVa7f
CiX9XYGmk0tsVV1dA/Sm+17orwehzxUXVcF2lJwLYIpA3PNnRSgJ8Ic+lEMrRwKZ
PPKBYYe7ytbP14HN1Cc1eDrMEd81zcXoO69FJr9Duy+/XVLvHwhOrVePVqkh5BAO
3TVRWqrGSxkqC9f4pg8gwHuOZtvX4fEAGdq4uoopOPCBYLrdQka8Ipt31r61p7Tf
vuUqeEPKrK4B5c5Vhn8UT1CJNc8INoIjIOq8VUY9MT6v249q12P2WqBkn9IB6qyb
mxzvvrC3P6o715jiE8BvQbJ/cbtu8cssXCUv0rM8uVJIxtwFrzJRSnOrzcwC0jsP
PwMh6hk3laIKRDoeNDThog3T8BRXqeazHm9RpigZI25fEG+tbbciPUjZ4PAPPrf1
iAAHnGsldj5+bKGscOr0EWPFGksjnIIUyy1mnjL3M4qZtvyXRZt4vZ+q3e/sfx+s
W48/Ln4a7DJOuhTntBeuJdwp1QSFn/+fKWOG7X0HwSJOYCJG7zKpDoMdViyp9zRR
ttGQ+yzlYMXb8OlEB0Cd57U+9rY39+5IuMeSb0EavXNhSpSvUNM4yNkBcyWAGTnu
B+eeb5SQE5ZTANMyf3EFA1XFTN4686DMQdocuittUeWdhOEuM5g1sD+9TbiGhu2/
9PVApjorspn5MtyO5OvXEyTsIwS7sAJgIa3qjkj/y0Q5uSYuEUmBuw2xQFzKbUIU
TPSyqyfAD26fOISwKHF9ql9bYhHrbt/Eq1lmUfmXOqGXmP82gHK96iHupVkbluWU
on9VB5lbz+lpn6w85MUXoe2fSzNZDCWZJzcO9MZgSsG3t7jTmVG/WTmvRChGQBUa
eWSpWCmyBF1rT2dHkWzFDWDW60rZp5OujNZj1IUZsd1IBph0PwLkaRQLvopxSFL9
sAF8oXZO2jiYnq+om8NaE17bShlSwbo7KwSS5etdhh1QtZfc4ZIspEVavW7pZbZf
MoSq8k4Mjct3H3nn7e1LDRce04vA8DU09q3HgNZeOT3GLJhQvoVPjBiKmhID3BCT
yr6Zwhj+FI94gDXt95J9EkhgE4xbR6d37Q1HxvQoS51w8KaNFjtoiJ14SiOoRppL
tA3sASj7S8mRdcFuQzz0QjJZtwcLSY3dTM/brh+LhmvtBzYqvBjJgN8sZ0bYb+02
Q+aVkCpRW4HeLWBQ8iFDoY/WMF47tE2DtNe9cjeKCza+ZXrfao/VF+72J9A12bMS
ouewd7CBE2/oKyKh8Mxyk+UKnDgVQXG5+YJRdXGt59r+Ixnrs1q2WbU0dGp3U4W5
zj00ZrAI1LjR8GOix2KXCObbUi0hWQ+INEpVySzKQWjXslznzQLz2SXRfxY0spGL
hAqFchlhAFTtI7+zgt3fSxv+sdgjhb7235jISL+PJ9+ou4V3ZTrp++3eyHWgA8uR
oOnjRoRVUFhRlGzs6uhTl1kbR0kEa1dFloZyi6Q4m5dx8bmrKKNFl8mXPqutQ7bh
WQlv7+c9dgMpr5vmJ1JI6kJxa2JF1uEbAizF1aeBi0OtEXbYT1rU/7hWOy2kTBpZ
RYFoveK2bQx0WIRTtz9r8Ml3jTKOcKM7b0PdvBSFiVb9UZEYCwvjyXg+ddY8LHZs
Di0LKfXw8ZK6I4pmeIogdHL6hPcNNuYceU1zAvG4S1UttjueOLsNQL4LynhOmv4e
Saas0/fE6VklJziHtvj1uJgkSTOmDc51kqL5aVs4td5u3MB6deW3ApDrRWBXIDJh
I6C3gJPRf4DW3+rizQqemoh5Bm7u1y8AGqtDL5IEI6mvronVRA4FSCQMAhgYZf8k
a5OO0vGuxH9o4FS8U2VRjF7DlBwPptXZvm2MHnWS7x2iiayykHD2EzrlMX+wFORC
eEe4aVkUuuEssDRcCEHQYKG+9e6/Q+MunUFRLOJGCaWz5ntpX4QHqXAQZ3avSrOA
dF+zA8+uXw+ECmvmxURh2tzd4UIO5eqMqtO9XNbupJKryFKO2J7MRV0TALzy2Yy9
uDmiE8KiP8z7WiCA+jqRRN398e1ZEDnMXx5bQzOyVXgAmyRlaiishubr2BDLdQf/
0kCZ+EbbmCK9ojH2glqRRrkxOnB6T2nZOiuqHbee5usv3ZKfJMow+Gt7ktKywSJr
Armyb/eOiRhKo4PRBdSmlhKNNZqD2ZjSbqT1v4/3BETxl2mzgBfAm0yAQsEULqsI
tcThYurEIS8SqhMXbe4kAEEFfOenWSJE95IlzI4rn8dGbdJGJNFXXaLbeBs+INtC
M+1yBY8y9J66WCQNges3dx084Abf/Z103Tsg2cDYTZqYW1K7KWDw7rWW2Fe9vpFt
+55ujzO3dTPEu4+ptdDGtZimR/wpoaLXZxShQ/66b/CGfrDVf0pzcuDCr8dvM1UA
q2bmxY4Kg1ir7jISizmf6yvhKgEIGtpqe3aGTx5/Jo3HvXqOrQKg4K7R1CRmWQjJ
UKTz/akWRZVRcpKzlvmtndjC8GLMXlctIckHB31Nv6gQ5Jmhf9T9oi2SKB2DPOuK
dSEy9ySbSERYW55PO9bPoSffB7v+OaV676vraxAylxocUjRHnuoWpHCAsq77RCZt
yEO4xi+ERPHsYEbSpqBhVNf25xz3d/lWaRn/oHsr67lp5DJK4Vrx2tqbmkq+OoeY
7Q982r4xxR31OFhJGuWOjnqv3jMo4bDIu6r+xExCNh3cFiVFYObEikhCi+ARDo11
LE7We1AhysJppShjrbu6O7IoKTnJt8EAaXl68sDb5RAu/6Bh1T29vI6xHc+rUjxz
cJHzsVtNhVJii5cdQE7KUKBhmsO/yNOICbhg246GiEokr/5ud3GajPPyJl6j6M6R
V02L9kqZLyuVGHlNnkFmNxMivvrY0EIOatarcSv82nLw3tPFLs7A5rzB8iw3lSJT
YpplU39aTpk23TthTORcDPv+dAicYvzNmdkh44dwNJU032IlQfc5hPqk82ql4XPA
XHHYtHFU3hTYTdVgNEF56k2eFPLXDZ3pqkeGnrUw8/Q7Onz9XXi/0lV4BLaENJLu
nRENsmLaqkHxrmueOcMfarzAp5cdgLl/nUZ44tb6Fk0SaODCLbQ4LssgU69u/qzm
gsG2D4tmCWEAJjwje6UUxO27JFeYYMNxLL+Dp3Bqk9cSVWtdCTepc+P/naaiJNi0
cCamxM3NCM7VfY/d3q+d7Qe2cgsqXwBV6NlxCiRA/OEfROTj8WSPqNQi9GjPfcUo
9ulqxhGJ32kOkD5UF0mgxg8OiAIIvFhsGUYhrMIXNKNdGp1OH6kyD1TI/eVvtLuY
Oz7iZFQN8KzUN7MSeqCX/TGUUIFLe5laJegvciBqV2BUyau4BleQdO5COIJV4w4C
KBK+vcUJZqxaelCPDzm/LgsV5bVDRAXuyNWDG7i/Ho4sDJy1irOT9SiQA67rk1YF
FYl4lRyO9GmLlq9YTa55S45NsjOlVDxw6E6GKSMVmSRKGCoSzyCatNdr0Az+kftl
NhlY4WKDopOwHV07xuajwDWN/jxdITEoSMaOh6mWnzDd6AbUqL8cjtxKcU8CjFmb
lc3ypsmvrT/fg8AuYogL7kvYJQUl14xsC/iZolKjbs9CvHDIM7Bu/8dLeE2cDOcO
kyv66NExfZjsuFhrgrOV1iO0sySDIv6vOo82zBfXbw3zWnFUZTG5jkJnax4KixFq
7U9J9hwlA8Dvx7QywWRd8ywKG4lAljcgESApuF98ZBoGWSumhAt96pFacqg2ED1I
MzCjmewqGCfljDRX7fl8kH/ziS2g8d2sx5uPjQ4/j+r8vzmBWZlILj9IqVemiZCO
0NibrZgnNPS74nbDgCVcXb119tSU3vUmSStUndHp6ZflPCkV2ltzq4JLdq52peVh
jcOWMBlnyTjzEY8W8RFadAi+CeSu00od+10ExEZZudbWdQNWILf8gR8mL/dk/YnQ
6gLDMdJrf5fc/lvEx0RyVK8ZICz55cfBoqdVteZcDQjkVx4huyYHGWOK7GmaP7CO
4nbTalzZFWDEBOX81SKmFcTmHUG1A9qdUqeKdo7mnnZFdSFQI4QJluaUxMBv0IBD
yO/AVUS6hoNjsBizhdJOFvIHG609kkV6lH8Ng3CKwwG0vs76O1xgpqTRHiI+cfGH
29ejUVw/NAn0YJ5fOmRwgIcvMRyqDQ4VDhg9m3BUA9ekslXDXJRqEa381Fy2t474
69JtQK+lP/3rjnXsaaqngMwTBL/pRQ1RjMGXBlfAY0i1xsF8u1jMxVL5/jWdFjgD
JoKSHALAIP3uQscbtdWwcYu9E/4ksRFyLDNY48G2K+XrvqJrbeH+CHqxftIqUl/2
LskrIkOqeFHuzr1BKIPgnhVZNCGRmOhIZp3umsMWpgx7DlMDKEJQv3eJOECVxLcx
qOnW0wqvPglvE6TBX4wshAe63dxgdSl66yYYxdru7iMK7jrBrhF6Z5Efv6yw62ST
JAHvD2Q9ewy5DXSy1omM2JttCGWtbBWrKXZ/XOuLnTSmw/jm+ETdwf5VWqCfDdJR
6tBQXCFblk1xNlP6GRTWS5XDB8hDb3KdWXubeZFDL5WaY3g+MWXzfWsOh4LHkiNT
W5P47hKIY1xdM0MYEBcpMvx6wRdupeQ3YGIsuyIeK7S9UHGQBgF6axV0/X5Dz4GN
rkjnuR+dElC6hN2O0g4BAV0d5045BJSbM2RgvjfMa/a/hxKygpzrXoWqEPEaqCX1
4yQKlW5+F6qqhwQpRXgFqLMcMQMIiMscy1sIM1fRgLjxlyLoLwyD8SJdBbSHWCFT
Z9nMJS0gHpV7I3Su1jKJV0CglOBGBBXrwrAi1Q7aIaXuJtQllldVlJrtsyq/5KBr
rUUnEcEgITPX+if+aACgaw65HUvpq24l1nn9DWU0uRflJzcbXxl877Wi1o6D+f4a
AmWBJcV0Ob+B4odEPEyYHV56n4bFXBmxw//Go+WrSMIsLDaKiZZ/81bRMmyRuWxv
1ugWvYC+OslrjXioM0n0yPqhbgF4HsrkXVqHvWHhvXxuIPLCKyyso7IQIlN3D7LV
U/U8V0J80tfOJJ0Kt3knhwr0DwrA9+QfidhBfdgq+tlawdN/6NXeRcRhllZWiiLN
bjRycMG4V/rYLsw5APHJzEveNClIftdmmXNlYYRfgY7uEOVRiPQXYcSevjEZVka/
gozW9BxCBIknadAtBwoy4xr8kUry5cfAHvHYQxIw2lupDU0hav/CY9Nzz7ftOhxX
LDlI9LxSgc2Oi+F9Aj3iaKG5MS298bAbhQYa8UGprXpQarENG9EXhJxzsXzPiW8O
jNV57SD4OmDytI5cl6lFhDj7HLkYW7NplJs3UnPTbFAUvjPlYgESRrI8EJ8F3+8/
LeDpBMzbaUaeSrCUcUAEWMKAVgCYhsKnSR8yDHaE1VYlV/ZqrrkU473H4w82sW2F
JPcb4vECUHlOwp7YpAdt9KOWN3V5+EWSCpw3XVlOs3z8PHY0AT+T3VfFSwxgLvYB
UZYaz/saa+mdKo7uqkaky2DtL4vfqFslocryk1PWl7TXiEXdZuAtqLyVf2tpIsqS
Tc5cFvUYQUtKxqzmTJX/Wgmgq546j/AAXUFS0PqsPKJW5YTjqq3f2YbIaqKXBRXD
dLt2fCmSHZBgy7uHCTvGz9Vn7rfiPl3mikPDBTrl8LcyG1gLvet6kfyWvTNHqv2o
Kb1CgR8iRjIMwxdIIF82G8RboepLhiEC/ah/75vDd+eIXNGQ+519DkExU5g+mPNa
ND0RXxJAVjhHtVZSIn1f8g3CmgKYrb2IC42QudutQkkDpdx6+PE/bSlPwuOCYo7s
yVVeHDFnyQv+RU/0Uluy8zRgH7FvWWoYO91Fk9IYUdQZNIfiFgMwtRh5w42O6sYk
GFYFm+mw0iQMRCDn6ytrq6k3PUl72Xgts3t412Llyitu75RXcKJ6SOlWLAdGtomJ
sIUhsau5FcPApb39xVlfidEeOGa0hyVp7pY3KXoGCjbz8wDH+6t2hKCfYb62/7e1
hy+pn6muz6DoV6/zZA9l7SEhfJ9CTV6QdqA5CBYrpScMrHUtzLyOrV0s8mpqNWGq
OiB5tFGufEQrXnMyGO2eBWwXV3AMdhSIUOvHt2Re82pCPjV4K/qKS09wx68i1ijs
ICFqB9UfenJnA/G8D/BfBqyhT9GjQTXLpe+fHS8qXDetvtznpbOwe3Bve1+zgcOi
/d4UJNtATOrmzn/TRMvdja5UPCXr0AJhxTefYOoF3bB2FADd2UyTNPE6BQOXXfYE
K5qmTjkL7Msz7klxzTy6qvsH69Vf11F33PZbJbJ5KXjIldY6gTtZ5Fcg/VCsleQB
/9/tGTPgX7gVyOkIeP7tm8+2OZ73R59aYS4wa5kNcZLVDkaGUjP1Q3/XevVDruLz
BSzFAdKV3whgxw9jYLwN1gJgNJkEsTUCvQQLDKadbUsjMWsto0qO2XISA66Rg00y
Yp0QSCkY+o1qLZ6UExSXqZhtLiJlgcHlPDw1Uec3iZCU5FpGpjKF4tmUZP2Uy3Br
xKPuM2Ojd2liFKZV90+dn8VcFktjvp7ANKu3HpgST6UBvlGgeMhmN59MdW6Na9X/
VxGlFZMXmwz4SXCgUhLvy7JPLH+P1gsgHQqrlsa5qUPgXoQ60pAWiHFmW57O2Dfp
w5AbyS9WERa3ind32XgRE9IdcvYgtkUybc0AKiBzHt6eF+Mi60zGj+j8VYmynEyJ
lOTw+dK0IH78TttKJidhzgYed5EXuYXNlVldo1vr1UVsHU8q/zbrxCiyu210KTOd
ea1qT74rW3OJz+qFshDBtLWzq6/LXCUgH1iHirOPn20hsAzCb4ao+22F9X1W1QGc
2sbMoYGzpYu9kFlhPIHlwuPV1gq8LCxHHm0eDyVDqk2RLckZG+Y/y8VoPoH8Y82f
qYjtpgGzXRZ+KqOY+IQgyHQ3ad9RquuPzbhNohNDZGg79eusB5fR+xkNGXK398DQ
od2lmqju8z/PXxWEcDMOYKj2A7fs/bUDSE8JeNFXsHYH5qIKLscrXvHgFE/bFfYn
B+LrROm6AIzqgATqIRdBDLlj7S22IThSjxq9oM9nItKD/q6uGH095VWvtI2y5Zx8
YcYf5je7lo+PUVRcd27ImApNVJxhLl+O6cHJvcYsWvVZVPZNqw6Q61x7K3xX/+9t
VKAIxOI+k0M8lEYuLyhyR+iAVzIR+VKATaKhbHFbzZzv2WoorWAG/LbJK8e7os9o
jXRVrNG3tUEijXvjBHpMsO/MxlvI9FH6xXs6FvCXGPyn/2QXZi7IRyvUztDesU16
sorVHFtDLvy9dFt9ze1MYizJeWmQqcYmQmw+hhsEuyeDRV+YMDIjtBZ8INL+Gi2r
Kt9P6gASZ2l9Oldb0lZ08Ts6zNikkYrnY4+cfm++W+ZvC8KYYgl4CQrg5QCudypm
6w8bi1JMqFUDxqR34d669c3DFUEkXQOPPFsG7v1IqLD121AYEaAghp8HbbfaZJzj
EB7T/99UcBi4wJ3rMas+TXHO5JGE8BtD1OzwJz9z77iYTRh9ByL/49MMczV4+/Hz
2EitCym86HKm3rV/4sA2TZ/P+tdbOvMY0uHRp+hqdvOEivXGXkZUSK4T/YuwDdfj
IP4HvdLh4s+WglTVVmTiz4dPoPrDNBCC2RHpH3OQJqheb1iISObcrhP88kAvsk8I
4ejYDoSMXgBmHTT7igF5S8COHlEF8RkIeBaXzkEXWkvX5Ch2BTYMoa5qxzlPolNH
K8AbBuukIuADRDiG2f7FeiOHPzi7Jl+cazyDeTV2+N7I5tEo9NLVSxaBYZGR31D3
JcAfq6gqhd43mvZBfoZSV1zElLvH3R+lr5Mrw2HfyRrAxxISBZAxdj8dpaEDCv6X
vWjua7WITmQmeEt/7+pFfL4Sko0wPptSuU448tRWGrhECEgtVCiLQ/7zD837gfDi
RKjX4Stlilgubw6vn8O6kQ9zf6SQr+nbAH4XIhgZqS+e6oUFLFaNG/NgweYRdlmV
BsgjnesUo0Giav7ow7+mwnF83E1SzCaL8ckYlNx5HyQ/MEhYNzOJpcp3ixO5ciER
Tu1LF8r6XyyaQ60ztrVfFFO5XeU4ZeGZWzcYk3DFwxgSOsSweId5iHDuWPKXqw2f
RhDobHSo6Vq2w0BAx9IBTgaIK0AzqnaOhqzOC30N5YNpuk7kvsHize+uQKN/nYRj
KyumL27USsqBPnSpXIhVqyf6972k6VA5mkr5IpaZO0xvnqZKpg9UE56aLzeJ4tpk
v1Jg+wb5yaQPZVr2idWrWROoPNvRMDwrDq2r9aRz7DngTE2CHslGBBqsTaXfLH5M
Fw2BOh2Onqv/QobMoe1mWitObqHZ8NQfU08R75jCg4mCoTCLR57q5+KJq6evZx5X
S4ojxYAJmfXnEAbEmHHzbp5YEJweWpAgImd41Dim1qyUnUqKPhiXUKo3DiG9kLWu
JxbV0FhZUuNWmVyuJAIawXonDIDxYL+zSPWV/VTAl6DwsaaYnHRW1Z4ztmB2sNsT
QP/H5szdrDGzLiahcyXTzPe6Q+xKTUFIeyWJ2PRGYE44dR+bdR84vdJM2rlP93gl
RLm/7U5Myn+KxpjKwVtVOpfPvO7jVUTVw3datkkhU35wOK0KZ6U7VRIwZNuOGoYW
bq+WoLZNgkhfQbgUGlLq3e2il+B2ql8mB1EIdGhZqevxcElYFeGEn8WWQTHuY560
sogfe8jv0ipfXYxprwj8ti2qry1YHbN5ufx3jTOoUWsI/idAkXMZZpc+WJ2DfdnG
WTO1b2jC36kGLXAslnOKZ9cHP8hZNiFtIxVpW3k66Wy6Fz0xWo709ySkkTpHS9ZN
R6UgJgim27vJVcDZFZg/TVjyPShZ2OmGE3Y5go+XjNgEFV7RSLVcPi0bWdYoNcTA
Zlw7mRh9wVSVpqAS7pYLiJoaUGqsouk2g4pkV+C6mJKLVVniDzuLM6hVLAH4tIoj
exNHjoNzadwwafIgXKu79ZSj78c3gkEJWuCw7i4C/c7V36AphlU0kDzHrN9AwsgI
q7M2kNJ/vTCYGkWmIacFnOrerG3LMpVfyBw9bySITRu8iJeGfnXYwjpJ6/g5KWip
i4gEj6AIicDl6roativkuXkxtI1p66pZn/jq+4cDJAyP/eTt/XMrztc3Kmm5KNBj
lf5iGjQtUxQbUqugnVOkTjqHwb8yR3N3UovqfCmEpI8GD3Lhs74l9oFDIEK3N9yz
FQdg5XChSliZhQWD0tIJDb5Zxl633IvMPFGVby5QM6j69b5iIa+pmc6iNKXSSexR
8hmbpQG8yNnU51/WMIY1WhzjsrWyVKGJmdw2MYPPG3OP7h6gNGR3UjlXReho4Adl
wqTyqkg9ebEn1exoU5KGTdlI/1CY50EYXLcnJg6CrgEVH7Vy87L5C3aMHuF67afG
My0vBsx9rq+ww/NboJAz3H8OGgYqn0ryzi0ieuxfx+E9xZHEGZrHuBzKZ87KsEVN
Dye90QPT92qfRwPHk/PyNfUekKOqLzZ1CVLuIom2kxB2nT47n7TEXfB+IH7ZE8OH
1Vs+FBh1H4j1knamx5I05VxcrkafBhylaZEBOWz5Kr2ZXunjNjUu+4BvZVg0+uWc
ypL5gfeiHDIUiwFeFrSYLkqMz4SapgwNtuoCZAEhbFjXXdX6vZEJpx5mf5i/IzMH
EZH09hVDGvVq7mK3DhC1MNMOi7ihNGsrbU0jAI3Ctz181pGJkUR2MpnP6Imp3uDu
bZNDyCxaxuJskjW0p1MzLoJ3OxGj1ZASONMuKO1X1vrTdWeeUPqxm17VlKzm/AHE
InfoK9674+RtOR6nffUYH8uTVa6+pEdKummxnCXY/5y6WXGpBzoPQ4HvedugN7IY
cJiW9NA8q68/meIJTTNAZQHRd7/UHtsbkixzta8ljht9dHxJwNUL1OL3c4Nb3va0
cpfORrv5AKGqot4J/1oULh8o436vl6NUGtA5QAszPQ/jxIB/+bLmDOhBbRa5Hpsa
7tqrTtDojBYaVcLxWYU3fWFo7S4Dk00lMMAGFFxijPKjcaNgkOQDobWVeoRAop84
BTkmS2AZkW2F8A6vcfGoudYPR0VrEF5Udsro+g0fCAh6ZclWPMdWdd3rQMvVJxJ1
nyoMa0UYm+MDtzor2Kqo9cBBgKQUyri21oddOGvBOBhaRqlLKqmj6bYEetSMzwi1
ABxmrSMFcStI07ZDRTm7Dc9MfWLlY4pcou+/NvfHuvPyy5oJAn1D4zEftoqRmyj8
fSqgIMDmDD0+rSHqPxwD2F49+NZ6q4Ksod7u0m38xhsedCecCvcOdXQKUPvWBy0R
3Lx5LkoGzJQn1u5DagqNz95av0FG0b31GzvKJfGRfk840dyXwirhtHnAFIf2wrol
fq0+5Ik0y5tRaprJuJM4I+aKJVJmd7BCf6Ad3QrRTn4POTOZbaM4jbjzL46nWqxD
BUxFD8nHVhOdfJI/IREKzwUH22srBv+ZFuETjD1eFbT1gf1K6j0cRGwPzoGfV1iX
3vE/qLhoFPu64OnEadtP0GeIHgBN0+ROTlCwuXbYycRJiBD24ohhQFbG0Vzx+GoR
N2FRxVmMGunAFzcmskdOqE17nGeXR/UN5Mfp3h3uVnHgzJB10tr40VTSLTzg9Dua
SZlYBSaiScPJ7tfk3aVKcjtWFhuMHxJDvAJaZiSL3gaKl1ZA1g5GI2DuZvBOIpG0
R5NyR26pun+f4U048FOzLpRGuno1bgLlLKn2DdjRojVfU3ISonHeMiOfwMED4XSD
V0qZI5IVxHkfYefnaTQ88N8SMnlX/lByj/HA2aIuYSN0NgQX/eMK/FaQRVnzFQEU
0i7IxHdJsuvdCzIZIa9x3f2zqKT9GjVF2jJKQ66TP7o3bDYknvPgkED9MXNt370v
ygGpbhMCQ0tdW3cOcVfolkEL4qsjLYb/mlFMMdjGIyuMXVyMzZBZ8lZzdNgvGWCG
gLDdgs/ENpkWrxF28l3AeHKvQl+Vr21I846p32NFSn2fCj3Rx0Vkskdf+bbdvptN
xbAWTR7G2Io7WqhxUVhCHYJyOAHLTmogF7JDUnlMBAtIB5ejR2xU7Sl2HHe3UExP
YrNi6O3mR6959QkKJPipfh4dJi5MPtRU9rK9yaGV2/+BPBjOhGEgfFgxnIhXAwYR
6TIQwz9dpb8njYknALBoSUDVAsrPbFhHs6/a+cDHB5wrTuIKr/W3QcTnGNfns+uD
tozaykwY28jot4GgfU9twaqarisgcN618Z3UmHd6BOQM8BVlSRcnU1fdwwnmTuq/
TZGkhlho7VTWnazyssUWgY4I0DLmUmdvmvCosrMixq1d0Nmj07jpxk3+Z8x+cZ4s
/hMPZ3ug3EevYuzMJfWkynFgiPIJnd2ROp0ASDtdjr8FdVhlYNxWHRerhl/W+1x8
R+ySnwyPfcs/Iqv3zqNnWNHgGKWudjMCYQAEhCk07man441DSkojIo/RJ3N4+jBA
SpP6/Pxy9bn8PIETUcNQouFp+C2EhIDxMDWNmbgQVfp0ULLOctzXqwndfl8vQwAL
BsX5SclCsYV82sdjQ9265VkPSsssW/QtMzWYtQOEr2CTVizC8TTjW8dd2hyrEORm
GJeSbFdeWD7ek3R3eDGtBD/Tu2Rz3NL6jPwATINTnt5FyCOsqhxyIY+WVzaaDtO9
3JWZEMJXj6PMt5yN9GDRDDF3Q1HcJaoJJ+mJ4BDIMRBXjrC6SV2G9VCNmXGsympe
ZdZhpY9CC9/LmSjjip5dOVuCmrmnQcrjanRnQMRaI7oQnrMQvCnK33AVE+hduqxr
mCcTZV9h7mO+VV4GoP7saCcd1pq3HIqkqH3ExRWx4uJe5ngGTRoSj+ubiAcyrM3n
u+GyeOqB7QRpBRDJhYXt1BfYvzhn5IP9SB5nK+dXu1jyAZlCkXHeH2iaSb7Fwj0a
KzC4KyQA2GVD/F4LtuBw3n9RmEVAWeRku/QjrVLPG3ZMrKmsHnObJ6Y6JaRwPVx5
rZnDOQxTW3sdFizqX64syCRurkH60sIhsnCWJxsIpDFJl7N7LUnseJ1Jj/I82Tmz
azeUG50QuzS7z4/EmzlmhQCfsCnghCCvw4g2Ji2+7xOmTYzgYHHFU0Zmau3WObXW
X1fhZiMCUQ2n6rN6szYOWOtRC1fIPWoe5qFhgXUDbnIXGGcmcnzAyqEs9Sph/zrb
QaA3SMkqiO7LjRjkKAumFpEO8FOGO+rzaMSXjhg9rZ1PyiE+S8DZYve/Ccha+qWe
/neCH7fKin8QN//T8RLgomqgscTyy5KHTEMz/139ytDEnRM/ig22UcmlYNCULNqC
cUU6gjcFWgQDTYEv9RAXYKxwY2IOExE5MNa8VhRMYNzjrF3RfyKaHVbkAYfJ+aJ8
NEqBKFnf7WtVVKIU4UhP07uK/UsqjI8BuEukaBF4G8mHvAvTx8SmHKzYlXSA56mu
Okhs1uUAS3xs/FMqZQI3aaqDSKxs+ynEVk1rVKTCTN/WnLeh9dLoiAGxlc+T1Ao6
mXYeTPTbNkBqLXGMsXXfRJQv6blp4kgsNyZ6OUxXpFgS2xnwfw5y9Im070mYmv9x
lOyJMlJTAyd5tye501zVG4DO7GdwktgzJNcEWMomXJSzWNP0mgo4lE+J92bIdqiy
tmpXEWKYywU90CtubwQU2Vu3+hANFpNIY84kaVsspckVZd7dmoupLQFjZ78fJf64
kZmuhTacM5pDF85Gw8HyKoU7wb9Dmu+FOwcS9YbpNvpH8PppS1Mg0csozmAyf1SY
nPQt9mFk6g0dJxr6qnTfUDmSiiS46SpHwMLNfeGcjWkRQTA9r4cc25QxxhOqjOvf
h6Oi4hz+PiCjRrd71wCOmx7tZv3LMzBSwwuSrzANJlnVibh5fS844iIjb5q3W5Za
wN2CFC7Vih18xBlRIXh8XllALYUCiflmx9b11P1pFXTxLizNwhNtMYkjogur2E3j
xmQ9PZINOP/+3DE5AgvaX8hZwlJ//NkivLs3cRPVTq6YNvOXOVIi82heSPRHSTu2
OLUQHp4bN9emL3Jbv9hmHMYCVwbcVtDCiOb3AgnwpWzSWX6nKbExbxmsZAJSLuei
LmqOgmxCYcvDTMkjTZsin5x3tpgIPLfMIZUiStSMLxwXn7eKWJ2sPhBgmtNlDek7
jx9W26cMx9ofzy4cpvrjtc2rRCLRFvNFcb9qNAuldhb3HPCl25zudf0K9OoNQChd
RsRc+UDRvlV0x2M1n+c4LHNCbco5/Ts+2gWSM7JHK2MUqImieDF0rzn54Tnnhb0c
iyZUL1p3GLESWPcm4flOmc8ruPNa/pNtd9COOxc+4rbtoRHG4HVbAUFElIB+sQgC
5erGLQegSj8nUWJ0FcuQmycWN/TCq3yZF3rU09UNfDCBRPJIz8zn0JxhiYGOrOr+
zKlkoDpWJiEOQQq/YuzOBGiOsr8SjeLL1H4vEYkn2G6dNtW+altCeTxyFp4Y1fGf
4M9kmmiguv0K2GmaJO8JebTZ8aMdv3JgM6gePfkRWUZJPiy10cdOw8D1vgKcph2H
jmvf5oEpWGAMVeHkEx20Ma+4SGHCUnYaGQ/7jzUsYZbRPf6o9DAxzTpf6IzikDjV
UnXJ5TzYNnEu2aRvdS2aB0ZdZicS1FG11nEkc6FlC3mRlHA7H8d7lw7hE/WIYnwG
sjxDthZU9F5lcwWjvmtzdoVkUVz61PXNy2Npn8DKff5h1pwQ7nfAmZpJbMEgkcbM
3vDuTXCxkHr70tbhZlqjE1jw7bb68YH6Sdy1ChVtTEWzOOaP1najYgZFig3WBa7R
gVMLuZH5dJxiMkbPVaRJ67xnEA+iz9m0r4BiscNt5RhYnnIM0f596LU+6QmBN3OO
ngbK8+i54KcFZKf1NrMgRkfHEMu2QP57tOKQsvTlnWmgtp1u+rVsCg4apWF9ysLU
qh0EzpsuTjQVQW+27Ae3AhbVYg2cK+1qdzNnRHkyFco1QMwiFNXKvJf0/JR4SXtL
qg4xnXZrax4STI+TIJco6cIiv3MTGFgKXukhhkWTWUiSAT97ZfH3mrbZDk8C3ADb
yTSyQM9wSFWb4zIE5qEeH5elRGo+L7F5y+UvekxSO3ggV/VYxUsn0bayV7TxwOVo
sZ7CODf2101z+GetsvDu1fhqTa8f9VBEjKuKd6Qz5ol5XHxG82GcmEfixVksjUuv
Ka6sXvJpodoz4vhi0w6I3OAyuLqdTAa7rl5W91y/Jtbyd5O/QfPgqnTBwzv2mNXP
JbTRP4GSp0Gn00MsKKylMdk7iTaH1sJMYkLYzpDGajoD5ov6y7Hoxq0uX8YplwRJ
CHXDuHyG3cm366Af3KKukJxTSQPVnXbaMbE8cXqy0eihaMT8b5NfaU99283yhLzK
sM+mh8/YwpUEMWOtmS3ohrp049nLmyj08br1w5TuDVOVdjm6z16GIl76F58jdc+n
GwotJehKQ/qNDC33calSYm4fXU6Hi3svM6xxrqzYcSjfG9q4HUHvbsg9iUU/+KzQ
zZBK7hBKcDDBAY8ItjJAScuSRwt9ffE0nyCSEHy/pgy+VmpUhMdBNLxy/U3Gi9fA
DQwN5ngQM79+ZzUe+l7pWPHiAXkDyrRX3sV5vdHyk6/dRpswmn0ijqR4TlnpuNc4
YDQnGPIyXsIYlzTh1AEsnKOdRwmsGiWsXn9YYQ6BBE/iQ6+VCcJAVPVKUoRLdv/c
OopTOBIru9/w9IKofnNU/nQULQJbFYKCwJGNrWAeKKU8g04Bve6rgKri0eX+4RrB
MleOY1rCdhtQ8rH/CRnVqhJ8YRJ8BisIsfNi16hiwIjOk000PAuEW8iePzTlP6kP
9jDL7C76m1hYbTkrSOc1Z/A1yHKjkwyoGHGShuqHPCIGDS2ZjhzO6mZ/3QOR9FlA
uNuFxOwtEYdg4wa8Rz/4dY2ZXQ7mKP9aZF5seuj9lF3ZLxn5OUHnf/W26Ealvvx6
uoasWaXc0lSMbIzIMs9hYnl0f9ESRKJlLpWYVZeWB9CChwM1kueM+pYf6eC1gd4y
4q9HxTY8msrKjNpfkzA+DDUsfw2/MpFCbMBJhbbfEWWN1Z9bzbcCTcjfMSK76bcU
lHawKz1aEcXr1MsCthpHc4qT9UYxWZR8u6ikiN60261SsppdeQEahVVCJdyXnwhi
YYKDYiNz45vdfajFdD8aFBbhHOJIJZjU9gwp0+GyzpFElk3EfcmnRT0vLLnwXPs9
lelFHrm72Ex+UqROtD4w7cd6wapcSPWJ/LICKLJxostQ30ogzHBV8qLTOSx18X2B
BC2edYckyX8qaGJekqDJmcKXhJzDgvTN2sB6e/KfCMg5bjjvjy+j4Aj68Q4gMF8v
U71F6fAfsVfGKJ0OXKEPNwrXzObSVpGq38VEPlAiQfflGpjx8oFqZ5ZSNoX28LGj
EVrZkucL0d5U2UnBCVPIvqMXJ/TvMkGdtM1P/dIocqIPF+HDP0unIeqhrm40TsQE
a7j7kYrdiLClzlIUU/Ry5j7/IO+irS+/H5suODqChGNVhvyaBt3akPBRbnuCQO1i
9SEDdCeRTEvfRE1jQ8mu9F463AtTN1izptyO0ujcCPOEkySZOJhelqHTaI7WaodN
eG1k5ulEgJ/UT5ZNF2e91X4Dajx5aqv9ZUBEZPw54AqAU+KKx2/OyAplEcsnnJg6
BU7m9OgDdjto3iEUEyw4Z0ZsPruAng6tpJN8/Rmzka8QNXWrmZe/XdWOe+C0hrSm
ggYpQU9LJR8bVTNa6g45fUu62OXqJD4C+Byg1O03RirHL7TCtBKIjbpcqnxZLbp+
RcDmFnk5OFQipHBe889SVNNVPgYS1WQhMb/wDKnU/L/qIPQYdOyS7OPXkpFF3xzU
miEZ/AYuT2g1E0eBjHclvT6ga8GzEcDJA+YZFUzM10BDiFz1pJfTMi6fwY/qyww7
uI4qYGSjs2K84HRqZV82MkhWrn4T2StnryOStUOKrk1/nLFpAeDTk8j/t/O/FeWt
juZa2jgmjkWeGc35u6FcqYuzV1dolLXGVvYQnKe8JLioJXXTjp8OwrIt0uaijXHW
AcL/YJlTVNiL9ARWpmm5M1WJOTeFlk41mFp2hkXYG5AI4niJ+bqqyArg6ieFJW1T
bKeiZuy8AwbgM6l2iyg4iegGpgruO8KayTCRzbKfhNaNREvRM5qZYd49mVYnFUbB
k/UxxNC6H6tGY2y3zgSjDn2CXjnMvY1Wi/RFm06AFlVtzMg9EbRjbTokQEvDccIr
T4mdeq/aqF1eW5CtpKtvhtq8RC0lGq/YX1bfGaoewzsOATTV7Sv5McYrp0K4Adyy
Rw4hzUS8Z1UDEH39DZH/+5Dg5Gv3QELn9D6iy47tQxg5OG5qyD2t7O+GetAO2x7/
RuSUAdZP4Vm46j4XnapAL50wAO2tF3fz9OGyYT/nJyxJO1SP1+te/d9G8omnzz2q
cFMaaSRzslYIni1Fy0E2m+TN/n+YRArmC/JHZ7o3tiS4s+oucoKDz9OALWyHus7d
yk5mDchyAjSlhuw3kqkCmw2yYR4/S5RmhlSxUt3fvmKVwiThiP5+FBQMDwRA8k+F
lgiDcjQKv0z7AVal0YLgplSDXdAOSE29OpbqGJT8PFlx2UvAp7rp7ZWIQcoAYlik
bkroDO7xZN+MT1G1ulVfXQw4lM8JhmbhHFrZ0rFHF525/ZZtpjIA6eWI+pnojX3h
sg6HEHn8boEm8kNPOEWazhzogSn6NSv8tloitpwWECgDiQhXMkpcXuxmSEU9Uav5
ZjIZUl6T6ZjioNHN+NhQ/XicZA4zadiMcZyYj6xaTf4bN/XH56sG+4CgwwUGKTCm
K25SDy9NcWdRJpVltfRcXnt7cMmYYSbUuWKJvXrXNwbk5nBYTTaAoPEGHtxnAi+c
ogiLp/OdFuR+BNfyrcHYqQpUCTxPTHH2MM+N2vO4OWyYnuR7kzDBr5clOgAmyASb
HeRAinT80IIpL7cDADvHEN2Z7ciJJ3sZ2FvZ0pHCb3YSbQ2zY082fkdxpTfDoZlX
dKLhgJpri2xnoycD4vXY/cwJ2hs2md0rrQHGDO8YMYCjbwgN0SKEgh40DTt8eWLV
v1t7vs5NgOOV80e+U8XTzCVLsEm12iv7xbPPtc+VFGIUdRe+NNV1wAjEO5+DUwyw
7qoKYw2PE8boMO2OpbeFdizmA4zxCWPYhNySFqm9i5XhExMIlz2977WBGZ8d9Kae
qOGLoQlLIFMKnlECk1jBChh2zgmMOCikGsy9CqlcufNihjf1rteVZoKl6gA3xsqk
+Algw7IR5CGriwS36cuF61FN/nMS7y02PsVW3z+9OVe8DTOXE+37+5EZ+ov6z0JA
Bz3cgCrxWFbkk+VNpL6YeMuOaqBPsoDAfaiyrDMAHXkPthlRPW484MqGWdo+EYSJ
HOGSWqeNnpfxL0vrZosxjym0poGsn+VdTy+iu/TZ+iY2FUXbMZshv75PvfSltRv3
zncfKgWkHfmILbUkoVIinUWeuJBOxscYJYaBXBavAtM6Tvn0ESq2pvAe9kotIiBk
ulKxjhVxfJHDkUa2wZNY4THhpmIif/huJ205BjhZweV9+ziOXlFc9GWdPiEMFJm7
Sdsyr7ZhKyDAPmu5haV15wW7yemGdgNBWKUHmJ6SIOlF1nbepFcpljVmiqadXQRQ
ClATXCj+TPXdDqu430vXBZL/n6Cqq+Z/qxWGoj8f2JYV67vJniDywGulTPLKTHtg
kzPks2qu/3SqzgYSI2mMnD7Lpv3QDlkopHH01JUmfepiCQK5GK42rNm9k333cHhE
mfyzLWTrIksPrkSv3ZWwDSc4SUJBKZJOTp8VlJHeh2demLSXWWKRV+Pq79bClbq+
3NLPOaHTU75VX8+iem1cjrUpaNkgo1y37vdp6P0I+3/xiwr+kbrO1U1VvPCzlIxs
/JM5tb2K+at8UZi+4FRRVxG5dVV48dXNG6yWB+EQ+jjxz4CnCiBjgrvcMgcpie1h
YkWPoqHjShhe/JACyxy8X3FxYXy+5SOSG+bqpHUUhZ4k8bOMdHPEvELH47LQpbnl
3LhcL/51frztj+s8uAuL8AXgqD3GQceBIRhWR9npPQMVaOVsUNjSMFRsf7hFDF/H
XanVC/rS894vCBYg5mPVP/I+Ax75xNZEgW2RVvJSZXSdo8en+n+g0qpOoLTJWh1P
xFIJHxGNOtdZDI52janez02jmayO+WQz0+yTcsF3mrxokvneazvFO3HeMX7ZBMdu
hD42A1P35iR5dERESm0hnqci3Y5EEPiNFQnrDPWh/jfzBYCo+VtMi0TvBRfxbRde
/pCyY/t8JwOksDt6xpWasjv07Jl6cB+UArIAreUGjKn1hwwYWYDnsNe2MfWHDx7d
I0gak2u6ieLIkB+tn7UpkXw1Zb2xHBwlN2oRZSZeoaS8VpIxpYxjOff4SP2BE+eW
iilXS5861Nnf6JS37b6ZWbM6eP1Gqt2kzUqvRPtAmqKTm0ADPKBgT9UF5NCcTRpv
xodHaxIgst1Eur7SJ3V+HLCFztj/+WDxL6Hah4292BX5auzzXCoB0C1J2qlFL1Gw
Y6oU0jIIDXcIOPG8a+pgZ18x58ci2MsjOTLFTtcxW2lsCfeTVeFxMucF9PS+F210
b85hrAaCkXTFP9sk9WG3sOqNCJ7UO2/8yvCfqX5vf9dswczDs0Tn5fwCbHIM3AE3
jkNkP/ZIq1z0JOlPXw9H0UrNaiQHbBXVETp2IU4nzzKqI7Df0t0SoIqywPNeJB9V
M/tTaPnXjODZ7FNZwg2j/zRGmNK71bnIrKB+cjMN06uERVarWaK4OZWpncZR9sRL
D6kg3d4ABxt0vFKRxTOTB+SZnyAve6lrlVfaq5a22jDL2888W5HueNAtbITLJPBa
YbaH8lRg//GN2TXy+i6a145RYnuHiEHlPqH28dOteVb9IP9JeNhrFURPmEdJhIZ7
Ys+3oQkdgvpE0wkaFs73Mc343vq8c4k1ii28aYFh0Cmfj5QPri52gxZkTlI9u+4T
B7u0styBBhJrOfyEc3wHNOIxOr3Vp2Kz+OlJeK6lR4xwzsO4qcF06d4Aq1hCqYAy
MXE857SZty2zfv/KKlzyrQWrUPohGheh+DRYxuHVMsLt1EWE6Vo+21scfDpkeJhI
z/SwXo4LpNM+YiNWItsMQJKFLDwli3/97dGTXTJs652PCzlYuhEZ1IQmQV6OQyDh
IXZzk02HfepeoraGo3cpalrsguEeUOAZIiNnwv/qlUa8+YvB6abTLuqcQEQB8oW/
y1VjsWEF0EdLJidFYf037JBIBNI/d3d2McsHdXGq49uK9PHmuAXeHFXdPfYeLylO
Naemu1pw6o/8ASBLba8Vj6uigWvbzln9jOi5Jil+TJt+vuWF296o51fWXPilkduv
ejtX7QHyFH7PqZLPogJomC3KZCKhYrR0S8NsNZcui0idCziybbH8wU3NhWNRjqoV
78BhwCKj/q1tOtLmibPXwTRMusOuOmHImBbH+KXVlgO5iqZHCuKdlNzALYOFpbMg
362isAkmhS2ccB1wh3WAM8eH50emfLm+gCSUbtmSLiXQewACM+R4YIZDkRzDMixu
X7Ins6dzRAq6SSzdzzHUViDaxp01DztWq3/dW8WqNT0xj38SSkMyuIQ4b16vc5tM
wuWxqQHhUGDAivp148RNNC+yRkHv4ZjcVO4hMrO5rfySF8pdc+jLqqEqWBZvdwHA
9iyXXaJyIBuOH6/PS8cDoTrXcS6dmDVzNor+JDhkqRQaxpMjfs3TkHRHaZhTAm9d
3/4kzRuVTV0wFXt7NiQqPZtIHC83wnLAQVgiwGLX+hmc1gfTOemhlt9IsYLu5Unn
JdQ2VK9b31R6B+xZrjke9fq/Us94sECTE5p344A96rQTpblxS8zDyktCmusDjPZv
k7QYkmmcefb6Wns+DYQ3NTYGOGNk4pqSVvKRciHYdWaAGAXltll7Sr+n73673ly8
aLYY7tQEUNG+xCb7poJhs2G8sLSDojVrA6uyyf3a9HULoQ7vsz2dZWTAgLTYPZce
iuWNcz1ozQwSebxBRv2ORMvCqJieO7465ZqnnJGUNAmqZsnFJSCyzxC5XHsk9vcT
qtHq+itqSo5Zm2Bck0ZBBEbAZ/SYYm7bSvd5utvz94c6TfKZcbGjaEz9l99HKjjf
ByV4IzFr3heq9s3T6ok7axgn7t398kCRV/3BchB/Vyzakio2NcLy6cwUzkejQ29I
t0q0Aw5keqEC6I4Rpbmk9JAUFdHtw8DbkaMmUfy+DhugLEQgAJfFJzh7v0w5GDof
NZxJ+9qpIFtTkNlVXE4XxXdJBc0iv0iQXS84Pw+NuygbvXvsFkjWRZB/XMQTOEl1
dpoi+uIIVcrZBk2axUcumGpym10kX+0r+yjmUWkiVWacHLy9mNl81xBoWvPIJoSo
CiFU4TOgtot97jS66mEXcI+roVJ/w+NQ1c7sz2RaUQ/ABGyySJLsHhXLU66ZInOf
EjzqvlmYRq29fUucptClvYJ50UF8PblKrfBWk35bmobTlqiZuK++9immDPHBcV+c
32/rv+mcv3CSfZx8941Icbv8bTK2WVaZdOQihbEdb9yvv3e3+Z3D60Y81Zv/Poow
5SSG0fWDGOILmWGxu4ed2DrtCoNCLJZomJ6z81mrHWvwo1ChLLEPuecbAl1pL0oA
eb1SqDNJzeIWc6R1iagltQqB7cpvVVyBJ7x0f15SheryfHLk3eRSDT/7oytiLPNs
PLHHIhg6g0oCiBNsMsMGL2ZH5jyAbose9xTmNzmGRG44HpU1N7OLe6gv5T2exWc9
GW+roLaGkJYrSV5Du4kotyV55E5poWYW4BuO2h5VeEFkeUzylZkEc25RBOHE57yW
+6zV030lqOabrVLh0JFO40QAOjqmWDZ+my1soW1cdhZ+qy5hCLCzjZbPywVlbcCS
KUDkXKH/WCgyq1e8rEtvw6c0fSghuvqhdMDYKTYZ1gSdvWtZr794f+klry+i5v4Q
2LwNc9SDqfJuag7/863FxQapOnPA/nJaJgUnDuscyomIxSDeyZgjZ5mdKyc84fza
lh4i0MpKhjWpze87ViMLPsYF3TNs1teWWsy5TYJ2bSCu7AZ9OKzxoKLyx1jqn5+p
rYzke0x7NHoWKOpTiNFqNBmQrlP/ADDOq6T8XsphAMY+ob+jw+8K2bb98TpIietw
sg5NJXpXllhLXZvuYKM8L1kTkgNkhyB8tF/H2AlCOBuv9jrN7vvNZNhgJ+Sm5UXl
2kHWNkJy8vydcrrfGzKMWPxQXu7TICgGyfMaMTnbyelSQ3TEKZ+byB/NOMw6z9Ay
TARzw6wdG89GQ+ylKEzJDOxUH4+39WGQeoUCcaycWblHA+Hw6zatWLc9kAyp6mSN
+W6wpQNqdZQqgBJsUfPNUQPcO990oEyw+zzNnL7wlZy+DTVYPGIuYsNwdaD7Km8f
fHvvHdu8Ge5lS6IMgtKzLQY1JEUHnwt7Q6ao7n/WIOchsxUuLCyCUP4rAk64s3EZ
eQb5ASI80pSQX4KaCGj6WWGhH60Yxd4rqPFS1P/3uDrZOnPwFm15WBvibEQz9dzy
PtHwgIuRdx6WOwDmpEaHnInFYvbSlIcblj/Vn/aeMfNHiOgZSHOWAeRL8j5ttOYM
HBxSCA4+Etx4pR7bA0FUzNe1r1FQdjPdrKmAiBmuNk62WMFUWcpaDTZOzWiOwyjT
RKllazXkGUQg8OXOz6Ogtr0bKPDUkEq8Bs+LKsRjBYgiBSWQokm09h9OqZn2VX9O
jcSVEPmY2kOkqddtl5bb4yw5m2W1bcM0+18d11YFR0yVtZc2DSXwHlRCKvaaR/XI
0R51El/pESXaAWbPra732SwWlv3e0nL/jsTF8Xw5N20EBrmbmSBObPsGsYLZ6gJz
XSvBu3l9hi1hNHWK/Y4j/kw6dHkcLTNWJXa0j6ETsSg1olUt3gfiblRTWBAHxXfs
tU69K6dWVmv/Ux9Fy5ZPUEkIweywUY0ZLuYMIJIm5/Q2aF7sFh1iojfzzAfgpIlt
9860K/ius1PtSMlUrnRMOWeEb7OopIgmp8ei/zZG42evzaryG1J7hgiKp5bJZhK/
LGihXoyO1ddDq8pRLatkZT8nRhenX9b1aeOtliqkySu5df+mQr6DILVVt9QQSBLl
jraJMkcBNcalrSWB3hLKyke1KBkzO4+G/vR+cEwGArbbrQcRIQh8Ymxzo71Xe1QA
gsj7EB4y1b1fVr2FcAa1qn+EasUd8RQZgZiySWiHDCLFVyAzsWOHlsF3EeHd1vKy
k6uBXm24T6e3to31rVZ2j4IG75lLXCMmN2zPi27pFTqpZ3YofDwD+H63lI6rWxz3
DsuctYBeSBTMx07h6QmsAwP7j99+pslgo0U72ILcP8C5HGdarJCtS1IiuwUTZRhi
OzpdzLqhJrQT8a7REONPVV5Q6p72pGFKNFd6D6ssKMYKmr909TjS4+13O1by6z4Z
7dZtdKRjgMvO1gK7b+m37W7L0XU/01xZW2U/qTyUOoMXGkbbTSJT8pmddnHkZxyA
iKEm+LdU2HviGylRQEGVvmNHf0OYOYMw1VvfJqlow0UnGaq+DZ8wNKYQPUGzOEW+
PBeETuErMWVtAAtVkGsaWXXn6V5Ov6+eQhUlxIFigAYvyocA/TRPRhGzNXtvx/l4
SZCXNqHYjmc3rhpRENRhUvvQjPN3LprnyksLD5o2psJIHuGH0So44o1ApmjzPhM4
H1p9NLK0Yq5zJrKMxK+l/l59XcaWmBc9FdaydiJ1Znq2lS86an6xd9CyQ3JEZMNX
xA9RYw4/sYfap5pT4Ar6VMtjwe0wUFxP/AsNlPA6fqcMeaxRfALJp+MadiorPDA1
qdHaoNi1Xk6nxI+Y9U9lqP67JyaCBx+32pVVP4vN2rXCgAEM0MrXmSdlk6bq3lPf
xzsj6vXYOskJW1Gq9DzYim0kd/JThpyDJ3rqnnsdJTMX+H90N8n/ZGS2+gxpn1ST
eGRvzTLWMJmAJP02sN0k6ySFqfl2w0L30sHNrBf0cpMFFBy9ghDSN9NeBV9SV4fw
Xcf/gOR7auX5QoWx3QzH2Q7dwPvUemIRJE8g6+Fu3h0A2LHqjzV6wOv+jOJqRkH5
n2h3V3pVQUrzcqzxqsD/bDLOAQweLtxWgnKtBmT5+BBXTcN0HRcDN5+hlNmH94qy
pWJ87wyLrXNTz0i1kNyiRxflLNxho2KpzcvsnZ8jOpFU1hTZLoDES9cKI7U7UqFh
JQWwFZ6MZVE+w6LcdzkBdoypn3JAIk0zJOHzSeKkttgPTXl87Ms7i0k1SMZ0natZ
73cuO/72pYswH3JOI41huqI0ywzCy0+EFiXIt5yNV26012BpEwOVgSeyT/S4b15p
UNfxdfQbf75+AsCciH8rw8E7nMWAeBR96sZzOM1cZMZ7bMWA3IAFF+W4d6fSua1r
snEitnxf3nGmITMZpD/2/r3SfApZaj5yhsMiur1DqaJ5TUPS3gsby/946PTjNBIr
R3E2/rAws1K49Rksx4Ik9wP8LhZ+Uo/eCrM2BvPG/84nfAzXW8YbKmL5/3xAkAEz
GbgKE3k1f2TiymdRN1EKJJcuuh5hw0hLpk1os9hz67oJuUGbS26MAw9FvfM9mhCV
KlKoFC/gi/Rm3aoI5LLsgov3NkL2jJuRjRDUCUTzziflnxEX5pVKPxKiDbbDxR/M
k3c4KWGa2G4gNZJ+RMb+DieTJU4gjnZye6U93I/1k5iHD/EcM55ct4oLggNE+DlZ
aHnQrq/mO2YE5Drxw/H2A9VTaAZyibDEf7nNONY/Jfg9KAiuqlx8+yKD0VV9B6eL
/N2XgJrKPqJmzhU0m49K3f0HAgJA00cm/vkbeTbIIfEZtRHrVVo0C5PLCPCT7+9q
f9hBP9GmyQ4wmmzrg4x9yIg3IB5B+IpNfOB9BxnWRLuAlgv+zm7RrzH6+WxLdnVD
43McModcYMXWbbjneHDpm3NZ5v8ABs/vAyRzhBrCfTBBmJZc9cl25X+s1mtabikO
PUh3k1YAQRzAl2ojBboGgI2pVMsVQaXFtt0SL1/2H3eyQ8VfsqPMInxZnyiPuSDh
4PubdKCqNR6kV5Y4V/8i8y760htoGVremPpas7v9lKB/UFKLeGRYhA8Kfn/OuSH2
rwILrzbI/uGQMOrAmFf5MMcaaEBFfM7MMPCFGJbNIXzYE/eHFzpfhxmi2I0uOVwk
goHuC3kZ8nL+HrAyshuJsQBJiY6JUVnNrSUW9FkhmAarl0OdJOr0RLDhm2l1D3Mv
ON/MIdfIwb15uH5jgbAFNFkrQ++ymcayJHWIK9O0u15Io0DKrEbvDRNAI+ysrFQ0
miewkUa59JL74YFoPOv26D6Jfv3ze2IneaaMToZ+Paig42w8GEjmZJ211149tKlR
TdFjzD+sGZX9ekGsf0KTEUO3S8QBmGolA3vIHLuZ59KvBPvboLeAH1mcB3s1hU1a
5Eljpdq9TplTcxwHbvqInAe26dI+GSGa2vW0Ikizld0/jJ+r/hGGDZ/6+xFyAwJj
JPRwkkAGpRSpAfDSyA1aZMdvBqUHOHDruOYhCSYJCHAvKh7LHW2CSGG2BTv9s+Hr
YfRsWOfB1NkgJOg+y6A2oBjaw8yunIt++xNcBpaLAxc96jYgJGKSgJNkVECJ5wlM
6Njs91wK3SZz55YPRn1DDyTFpOU/Q1KXLCeORjDBuLtrcoW4Mc/aVEZ1EZ74AZWh
CSjxZp6xN0fnP0RGSknWQQHOf99RyQdT0SmuiaVeuhpkhyhOHL7aZ2XjkjO4zp4R
jz8w8WckS56I8r3IlDKv8xlJspHL2bIQKm2Tzljt/VPH3JivAiPZ9Wmn376JsIjK
pmtfzj/uG2akyB596ieQiyLdikJty6a5rsZ30dRwMt/i9LiCnXE+fNSrl36E5p8L
0l0LnZd3OD67FHS4n+76KiZiIoEqjNC9w/CpHQG/qLtikokFU0QSS09MimgOVtsJ
omAfeSaA8rLqHcorWxNIpILifY3T0IKzIMrgZkgVzdMYJ4/xU8mkxF908eT41IkP
xwRzuGI+4SZRNBXVIIDwqIMNsLexWQTKwDm7bEFsRgvtNp7zpk+Tux+dXR9sj+R/
h9YlaI7cOMLupdzWmH+j0u6rmBbk99HxLKr2cuyW2+fxMzHLuutecgnamwigsxjd
GXLTkWK2DWT/V6eA5FchsG5Gh2Vo7YU9XKu/BiyUjJp661ZqUEtR31iJBshCUBci
WNth+/0HmyIlPMX5QopZ/GhRi4LeOsAO/zZuHU6eTQSuvr4W+6c1ftyfiDpIF0yu
9RGOS2oI3gh2iMS4GWN5hTMst+ytkq0zhJI8M+2hnUaZps0aXPK3ipZyasDf+El+
8bvJ5Ra7QLTBAjRVspCweV/jaHfpmpibzKxOgUQjrHobyuSEy7Gds9F4/hO7xJs7
rGkOJxBv7vGwA7QQ3uC3E4Y3pY1FFNnpck7aXzBvjoXVzS2f4kdnofQYdxVkvG4H
9tt8uBtfwG4fKwizJHx+MQ==
`pragma protect end_protected
