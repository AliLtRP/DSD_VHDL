// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:11 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
bt9wgtK8nVQlDvXIwatHhyFNMmxlpgFmja5x0Qr8j44GFd/6YCtrwyryr4nzUF0S
7hBdR7sB8UZxz7FjxZFaXqH/dG4Ecdk9VC2otZ4U1aPcwyDoS2l+H3puyPWnNuQF
96Chj8dz1foZAkIl8VGygmnXpga34DChIUvfMs0cUGM=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 23280)
7dUzYQRDmBEU35/lWZJBVA93aN1SSXbe2w40xAN3TJMQTfyDw7bom+H0bvKYnczG
6oxm7wVTEoI+RgIaV5Ri9bONGO49XUCZxMobiPyXrSXsXgine6wEV2b4CAxe59q7
VbB6iQWwImoBDkckIw1Pz77jtj/BWBUfCiBKwchWLXewQSdV435sg9dIe7DUIoHr
KRZoTPpT8Qyvkb0++OutWo5h/D0zCXxlJxA7HAWtGhAJ4mRHyj8jaRtp4Kc3/Hth
e0NRlI5A7e6TURQU5CwUVubm+q/cqV9xBleWIwSYTJJ/grBzYTsSaIGWV3WLlN04
4Y7fj78F+JvBIWaM95OeOHsdexWqzeZPmJuK8Tr72IYJM9Okq7CabCE8R2Ywk2PA
0ZLu8bcOdR36eUqqVYt+7JPmCDiYMz/yqYvsvTIpBGluwoKOy6qsX5dlskzkLE21
lk4gGHrEdyJe5h1jCGTJE60btrmP9Wusqrxu1AbCuITuw0sH3xAfimU1da+Ol1Wm
y0tGd3EFLCvUIgr+2+F8+ZuiX5P7IEVmZVwukt9OwyginMP3FeKKKA7UCccNLeyH
3hDDhfn/KbFHLGLodmY1epeY5XnFK2wZexV6xKaVds5pudiCp1GAfLSEkPH3X9F/
DDLqaBE2tHvWkBIRg8hysgr/TJ6/CzB4ahhHXCvQ9XH0sinOne8qyToHIbtMRxF1
E0cBZMZsw+3FnxrK0TbDaJTC9ldXfSaq+LrcKxF/b8FW2jPAIY4o7TgaB6py0OKq
gQFAw+SCg1gxe1pFrYIsDO+/9R3VyKslUgwhkQ+3y9GNpHsI/udQ9fap4DEdj4Sf
pD3aC9DihqVFlsRA2CbolKuvz0Ukvfb6ZzjlA8KDRtrjzG5QtKTIyVEDaz24Ce+w
/YpohsKt8uKP43MG2W9x5RFPdfQkkIXrHBJNPRywEkmyUmkDOodeYOIuKSE3VE4R
uTkEIXx+bxiYW8lSEJ+n+ZX7Flz9Owoj80zs+WoSZl+UtNcUIo/3fWtHPmwVGPPX
yiSUsT2dYOalEoRvrv2T+GoFXhC3iZ4elBsZI017pnGUv1MbCSEzCvUfFub1aL/S
R2sP+KtpaKbFz/vRJpHhYElYP3dy3ncEzLVcXl1fJJm9eP+ofGqIt5iXcVXDNu+g
0BlnEPznzzuaTGg1vPH42MT1JuqsN/5lFjuel+kKd9vGwrOCY2f14xbRXoKKbswP
fD+U20mclgD1Dc5zm8jQ6dW3lr93ZD63Zh0GPLpjZdLdJbuDqtT8uKmB++b5vZ9R
yF/Gb2oGggmY84DC9iEcCljCUzs4uKUM6YcqElmAj1BM//QB2r5gOaO1Lzt+TTpJ
SKuNeFs+wyJU1fVA7iqnbHoRXvFBw/QmRHwZhjyU+0hyX+4PZGJ7syXaC7DQXW1j
WzjaHsMckY0rLQLhG4MdNZYpPQUESFYENTKEKeXks4VcdrMYDddWIxyeiCro+Jko
A4jNX9SIw6cb9IXNIl5pNrdNCAu1drVoszl2tri7T3poanYeFUci1q4fQGkKpDmQ
ttE3r9lpjlZztk0axsg+EkS6jiUg2wVVgc0W8LzO69DycaIWIlnXNagj30dMEIxe
Dw4YbvZ5HqXna56uTvWWlSWzxZRb025alhhizPJ1BM9qFaRqo9gcwGwFoOWwymd9
+oXC+XWWgLIOS+2LDH9kjl6obfUw1sEqi8S9ywbfIznEZ68Ip4r7nH8qu95bL4i0
r4m/KP8JwD+b+Le9GC78xVnrQ+0irDc8/NFp8ZQADDZDLqeX9NZW9g0jwPNcVw5J
/bRIYDGFSgFwUzUjFr2CtkLwsaVmoUpOo+sJRAeDZwKxtFQQXpwlr8VsQ65QfPFd
S3BvcpryqgXgL1Q4ZKmIsuRXmfW0F3GXyMfczDHz6o8VOgywiAHCtMXGJy6fMX7m
Hkdx2FtfSYlGGZNmnpnKmsP7eBP4B0JvYEEZ7Yitu9xKmAFdWB+PtJW0anNGrqU5
ERF3aWOFylNOz/1EmjTcLR/GDAZiEN7MyjS6lZKPZSFHDYYkmxfCeez3+R2ElTRn
TYqARsEXfjYcawRcA013aeaNO1VX1FNlUs8vax0aXoE6b/2GnbzFqdB5rObBb9n3
nGBimGAwxkyuXTzQ/VxLFjVRIcJ+/W+vSLW2XeT212cVzIVZPpdU6lXLkDSmO+SP
Oj+FvuI4qm9EmDW5b6b4j02MWXeSzrYncq35O/9KkjTIAqKcjh7qGaRGyy/oqsn0
X2qZW5Dup/jfEq2ruotrfxFh83/H8sgZDLMTzHYzCNtjl5d9BPJXUEzEeX9nbED0
baZIcMDt6QQAhHGO0IlEvPYrBINfmB78T7iJP7n+A1xmsA1Q3JQwOtY9Is/payy9
CZ71vjfjlJyjKvSoYdpZp+/RVSjUJ4BoKAQfbqH0sLdckYYvv8hS2qPpUEjuz5fq
uWBpYjYOAZ/G0vX4hX9XCzR1HHx6uF94Im/8pAEWj5GnP7aIrMCAC4ncypefEE+h
t26byv/WgBuTrnXyHa9Yoh7mY/KahyZdWprDK63R8g0IkAr5OrgwvyZd4+/gmg42
vhwAguod/uwnsdrVK2KrmIBqnNo2w4f3xscTOahTi/JFrKvfHvadbNA1EyFeFSVf
c4atsdNBN37hyAa18WmvK+zDl5cMHfmMn2DMgeZy2eNlAYH/GnMlpcUyPMXbPJ3S
LS7FcwIWOpsScyerKq2VcVcPnroeGeJyO+d5PY4ek99+3JXsLLOSmZ4t1VySXOs9
4ezvEmtUTpCDO1BOw8lSLprZa5OHdlBGfTX2b8P8aR604OwEO0208qRI+MwOOTMP
+URg5wfA8AVP7EJ9E/y6LxPuGT3NlY1+NpvEjRIYhFakj1TrY9h0DGdstfqvfud/
x/3AdXjrpmU+iv2jzFatfwYBh/Bq/ZREGVrcP06IzJk5Y/lnrO4LLuCEi8XzLPqn
DA3+8PZA8Y3hOqBRQVO8nDRF3x0IQh/sOL009+JP5ctNkaAZRxesJwWwkG29Tbbn
vXdEwOnhzB0uTE27Z8uh1EBa0K9mlI7FdjT/jymWegewtk9A6NKulvfaoA0QRROm
+3lgOImOtIKxngWDEoyeB4gCh741J1r40qvDZjt+Qapj2YXFxx1MS417COfXp9wc
Nnl5NkDeeV/jQUS8tmaXsBZy3dD6BriTWqxadNmWKVS7frHaLuLTs9RohP+5OPYq
Wgz3/Klf5d51632eqdUO+G/34RbLMd4vswkkmjpWWRX3ZOyWJPis/NLJ8+l8zXZu
ndDi88DByPsCk4ZE5Vz6bUhm0wkCiQkcaYHTgMpt6B4WDdJjhIc3Ytjf4mtPQy0H
njG2AbxYgh76efK7C+4NBeOe6ZqQJAk73rYOd0hITWJQXv9Llk9+uPEmbipxwTQS
xIx4FU4igo01G/xyffK/niduYq/dWpiClK+2HlB8motlH7INSmV2CSXTO7q3BRyj
5eVLezsLXd8ZV6Ko9FHtVJmjC2IojdaYP677tqAdkogI6tWED5KVDVOBbOpmTHTK
5eWj18WULQYYepaRxtO8GdxdTI08Arb0UCebiwTsl8sr7OtOWAChoASdnVZbGQeJ
q6poXzOF6BP7d6RiLN8UDFSLIslaSoOTrGMn3upmbw+ZkaL4RLAvh6eS5Dpn4nwG
1JLNbixNu55eK4r9cLaRAizWoYPl+dDN/w9EU8J3S7R0397IikJtxCq0twMFbelJ
Gzgw7kTK4VahCZLl32a6XSv9ebNi1hUzpkF8XtxV3WNXtI9uyVuwRKp/p1IqYQYc
ZaKhncVfXsSz8obPHyEdMNZ7B+D3Zns4yEV2jP9icAx/2tCDuEwROM5QdvCFgOUf
1ZqklcWGey0OQCMAhkdeysQB4SzvzUqK7Ib5l8WWFF2rWPB3hFjjYUO1C0xXUBK3
i2EHpNhRu7jlAWhQeitx122Qk6mmfbiDqHNUXNL/QzG7d0iucyN0v+GwNvDw15+M
WAaR4lvZ90kU1ZO449NPSumMzbz1lTfJLdhJuNAHdZiHfH6EyEqGJIeeFdqq3nIk
4eOmcYT6cg+vHaLeylOraj8JGQnpl05lsoVGc5vRbaEZKLFl4rc6jqCGrUR941Hx
iIP035+uN3QGaEjK1TKJvfoRjYBbJj+KHR9F/lYDJbQTcQbfVlHNu7i+yHzbJilo
htHkcELXBEZHNyEmBNVdVkVUjpjvSiFBr/qrOah57LqRuAQWzbaDp6384DwEVdaa
ScMTyfkGr2w1YoPKRV3n1R07IgS8zVMLYwNuxuwyRMPYUO9dTbHS9htP8Hv77E5I
ZP56obiWmjnwamfE4EvSHg4AJDz1Y5oTla9kqaIIqqf2W8Cz1RGlSRTNVYohf9i8
39b9zRXzmthdJJ5ZfagGb/9tuWAT1Wy8gZ8JeXjksgdr8IVIo1orj5Ej/D+3TWkT
fSKrJoy2DvjrYPJfHkGjElLySX1jSdVvDoZzO2RT/V5r/ZMRTEoNBv2HFC5xO0pg
PcnE5HZocrrWyAtxhNYZ/OM5AIxtBfbp+Yz2OJsRmOss7nhD3hkK2SnNFNHwtRvA
POxfNJa32nIZTK+kko3jhlijkST0wkEaLwWwkwejmNi3Hg0Tj8FGKgaqF5xeAbCp
U72TzuwWPprmRJtssEDmc7/8N24ywoCu+QZ/8z0YDFuGr0w5BrJ20407Q6slyGkx
9n8gyesCBYBE4ASHKyzckqGro/eKx83WY+fs6inWFPga1gPUeutIq7f/NP5U7zrQ
XfeAMWyqgGZXX7eTE4Nuul0ABUQKo9LmOeUq6pojMrAuYYE9uddJhZLJLHnuFhR7
4cTtocAEvbyR4mdH0ibNFpiL6b6SrXPCbM5+FjlxDfhOHmGVE6/tSviXLddW5Ue9
Ys0251sYgLpjIrHQ0vJUww3OdknGgOKrFoumDWdK20cQ3y1wFivdvFw8XGsop8hc
INAS6UG5opWE2UDj5hDKYgY3y1DXwKp4ZMByayZAwGvov3c2Y+I4Q6WamquwOKN6
Lz4KzEXGrbUeLfDUe3Hm4S+iQCSzIss81UM7kKsYCRabpy/7wAZwF7YMB10K3/1V
pa8uWDruJ+IvUYAgQJOMPMg5IwbecK8zgRrFDM7S+JMsK1cb3hnxeZD/3JAisA+y
tLdICIOQVskHH9wlaqX+3tbqOCpUYTLl941BiJzIx62+Qabkg8+2VFbawlxze1JG
O/PbaUjngCZWsn0kccr5l1ACIJYzJ7K6ns7Z5jRr9OUrKUjDea1x6UaqvuLE72KM
lheWAr+JdCfwpSX95TPojcUBER31A3sDvWU/bqVLyo+Lczq0JyS2byjLJmR151gv
OGi4k2aO+dCf1c+8RoyFTQxUAMKEdigC0ok4enCdLx1vgvdJ5vkzIOYDRTGkCQno
Qfg6Z8M2uL+g6eCI+Yi1q1rT5Mkdu2lcsPZngEAVZWQCxjpoLIySUoiusNZwiQQZ
KPZASlL1waQpmF7X+g5RJkz2lsqFkUREforragE/HhhP+jeMU+ysJKyPkasU48/6
8FUNNOt9gC/2B08y688nuFFeHnn9vmyLdOBV8qC7h+l2UK1bIGi++qQT87P62cMj
siAzYnBuLxmVLW2OErOqdjYad/AGwpd4nibe0ZScklh8yd0hlaZ3MVh3j6qIqMBG
rVvxqMm9uuKTyWmuacpE9YymSkcEhhgb6ZkKwmvl3p9DbCc5r4yKmq57R5XEggK/
8sJDmiT7DaBDfgH+Uqilm79wGo/FoxAOewdWggdHUeyr29lgeLsNURF9TX3ZMuk5
pGlK9SqDxxHHrmiDa/0dzDsB9iKAErGtSDo4otkOjyQSbUrAlL2WM1BVy4ey5PGU
3qMi1L8D60NgsR4fiUvKY4mm4eQRYmqbrnLWQnUsVvQLYgDgfsTQ6hrgaC7gDs3/
LW6AdpRjOoOAqcJh8wb2VCDZpCfyGFw7VrZtoL6cntn9gZrzTj2N50YqePQER0WT
zDQJDA6A84IYgoNRRiFTb8yRO8LyTKI3DvBbqALwr5qST6idx4tWOx+Rghc7q59L
4XtJgvsWbkZMbQgG4pjxWkFqhx0ZzOJmVl5v5h3zsMoxgFP40/EeebAqtZLoPUDe
wDSF0jadcrm+bKxi46zaToKHToi/8blo2nlGrqYMhzdp/loyBMWoLxWIJHgvOE06
UwD5uAYFkWEi3ZBT9Jm1i4cXvPwBDfdSdNOPuLqU3tifGakwhZ5g/NWNgT+Gw73N
zXiSvDM5Ot6AZUeJ1Ky080FvgEcA3GDnAFU794uYapKH4g9mIGkHMvfKCjYkdoi1
BzN7+sJhYTDix0qOsvaKds+e/5xGYi0EG0yPMeYiOj4BFwmal5CU+M6vpInlbpMx
aJtkaArphlE3NrOWVfVOjsPAS9AcalyNLmozfORdFbkVuU3cO47hCoOjUej+cXVa
pRhfzqjbW67yr937vfYl1M4VlEbB9TtPMEDTNZVt1Ud+ySYNUCBjAVV9lYPisRWl
7H9XnYz7dUNy0vz59R7cwvdm4DxB3pJd/0JvA5qwJg8IRtk3YbfHj6dMEiaAhNdt
Z1M3yvurgg7SUxnUSCTb3Ygy47Tgm57EPWHxfIf2saUbhI9fdAI4Dy7sXRbBKkE+
3nyLIAgxvz5Xu3fyhi7EOcmT90ZFr13mllMJ30BjmY2dKJgIX0H2VGNJ4cyyCl3O
enlWwxrtMry0qmVb6PoPhUqw5lbyZjlRVuom8xgdIAYeI7jXDrSqHy5d1GbAF1ht
gpMae8UlxAuvvHCWoti7GEXlWgB0Ox2fgVcJ5N/c33hEF0qgWo5/sTdpQ3lTDTN0
8TLrQ8DnOA7WlV4CwIg3KgxGbgK8Z+ZBBV14ztYcHyWhprezWiFbKD+Ribmj8xT0
TAgFt+y12J0b7QvPJJ1xwDfCa9CTjnHor4Z0Lsag0YHVQQGzlAE9NIgVyocr1d4Q
BsE5MY4eSpnaj8zAS9dDSxrtWyEriQdNctH3szvvIb4FN8qq3UfEhfEkEFvIN6Ft
ZO++ZI82eFjtvOhpS/7nBTVS8kp7v+KJA8eWmMTDSxunMlErMUaYLep05jPSQgaw
rd6L5ovSZ6ebM82suXMm68Xc/m/sjfxh5cWmVd4Nn9RnB8MDQ+U7P3lLAiaLyIJW
W+o/20MvnZlaMAMDAx41ZyP4SuS1TTGaZk/DD5R1Gs7BWON1pARJ/OOKUmYW6wne
G39DrvRZuK0iW+QzosYe41z5DQIK+9r3rtTP10K/tCSqY2bEVAgfCezyKBbxr1vd
CJ2uFJrD3WGGxW1R6mTCtymoCfjHVWCBqasfwfU1OjvkoFUBJd7l/Kx0skdonyo/
8gfyABUyhsK66NocGWf/PffbssP0ddtaAmL2VDzFSRA6G6OHBOdtnQUaPFDw3DXX
Q42NuhLijZ/FjMhx4hPfBlLynqWLYl/f01QwXCKQykcff5kqUA6JtFoulNySycg8
chUsfKRa8PONgxgkuXlv5cUvPLRKlwadFM22gNGRgSgperLrvLpIA4/Q2KKQqdr0
YsD0r8f7ctOUk/e+knRyacdVcsnL+LFdS5V643fpWOy3PJlp8OUYyXsJizikFD1y
sWvVxt5kY+KkJ78KrsvrupoRJEjtL+apTeSRSe0WYUUAU7Qub2/NtvI1gvkrpij7
Px3Z9Hwj7Xgq70F+QRZzQNHcM7CP4r9ZCZbJtg+Qc4GWDlEFIaGr7KJR2iBW0GTJ
maL546tjd3PE4KQLh8MiQiPT6wPjS+WHQzFZcxtwPa2dE6KE3RPhXclwp1zztc5z
UsqGKoyQJ/6k8oR7jBUBgjX5McJrxITLQ0T89alIl4jQv5ZMfe0Cd93wZyDj/SxR
V2V1cTlIjvuuJDhsRhjoOi7M9DNqw7jfSlFWRVyQ3qAe1ty6ZMqumBbDAWKV/RQy
a9XxyKt0KGKl4arshLI/35Ii47BQZHdHNYlPL+g9lgQ9vkzbtyMByT4WclpLvLmg
Nco8qQgSEtlYWTB5MFc/pQ2SzlnPqqfNHQeK043lzDnrhdClfLixQA92UacxxXim
x/R/t/BVTdsCDWzGps2yewOvjqbOfr9dq0Ev1EoGIZky2jj3vl7twDs8oR3xljVU
bdHN18RG4yJ1s3Fb9somRmBHj4qy5xVD1vi0xhgtn1QOOYBxKtBYdc5yQKqSS4m4
GlHsDAMSup5xsb+3QZ4aw6iKQ7N4gAOHQqd4yixLN2C+6ci0xhlw3NEHIn+G0jC6
a5njEJTroBNehKnwfgrLj1ptlSB0nd8yDbi10EqKTV8g8wx2QwhU6TMjNnlQ/sX/
aejeKDDXqeyPmovQ0yeGj7KhgUeb2ycdDfRKrBxFmriTYmvaloWWUfWHx1FKmJIP
oziytCE9/qXfO5HeX2CeEXsRMTkJTxO7P8FI6aQfH6ixOYIlnUSsM2DA1MtDF9nH
/lYCSWyXHHxZCiubldDeytYhulpZS8axpT2dCANdM4kegh2IPDeKvfc56Y5JdDYe
i3dE2BBty0EU0tC3Qn8nTPCsl/vPn98W6ex2f+Pd0hSlifeeUHu4CLpM4qlaHduS
ljrbMdIB/843xic+Nnjw5Wkzp8ur4UBYcc429VOVXXTElAu9ZbZX543q83DyDvfv
7hVmndmAyu5yrtUgngGpX8GJDRfJ4arXyxphCWWVwOXsz6iCBx48YqfgqzOmXU41
cBNwFuTwV1zPAnGsOKNIFERLM0Tk/JRbpeK2wA/lGheXx9AA+n5muAFEANiUYvzz
q8g6Vk/AgH+Y2Pg1tsmGUKHuGFuAeUYfXH5YvGzxHcXP5Kb/qTMzW4vn48oNSAwx
7/T6nFvTsZ6AbI1YG+nHyh47eFd1/TIf7NWk4m3/bFykR9rfJsAZ6GOHfl044Swg
wQN5fDIqwVDgFMNfILITFQ0o6cdqvZ0paUBUlxX6JTIDbrXG3J9+pk+81X0kwnbE
Mn9pMr/lt5XYZvHZf7gkCOswgRhixhVaz7a8R6AlnnmB819kRGWJqFxGfnjrHUeb
iHr1unbFay38FCHyz1Hg2YBg2VaI9R++SAcTtKQu1VJD729mssbqj3l9be1SK3BL
Q+gGAMrLzQxoNmgIrCGSj/ITOfrFfgJSrhws12kFCi5gcg1xWBVAUF3FE4vynZ5V
SK5P1aIslNNeTVcv0BJKHBAXyHHpRO71nCvIzqk0Xv932+Otc71O/AIORW/m72yt
jblmfS8Md0iF/1c3X1zkiKZ0HpU58wB8D3Gm2ekk3Fp+dDwqU2cw137YZfYrYB/p
cxh84hi6g/3Gcntuod+b6LOMwhF1mhvQwEpLyqqVZa0g/TYWFd6xLnRaXyYlQceD
NhmBNJ35sRoTZfFNWDq7yWmLtQPYzXOcCkWGkqs2sPHKm5B9oDazozziAKiIPoSv
YpC9yNDkRpnKPvkCUj3x0DKDB9pWQ8hMFXVZ0XtfvuzOrnMYJHKsjIud3pF/m/sC
XPx7VjVg3LBoUcvhcDRdUaFGgg7hadVDHsHhPGOfwH3ZhtnCev5YGEFSAP6/WuL2
+FGTiEJtDyFEUoOkYun8A+HWJjtJGCewEtHmLIMjzICC/SIgfx6VyIUpsdcwhvag
XE7zXNIbzth2zpjSpIkJKfICn8TD3438+9t2B14NBRawGsX2nL5sFPoygzy1O23r
BbYKY4ELdOpBMw1yrmbGGtAI28ynWtcs/jMW3lz1P+gE7JLe2IuuPz1v51ODz+kD
tvOzXotRP+HHaZOSfn8+Zk+TBsfKu5gJCURbpK19b4/b2ZWZTT5q4afwXk1iNqE1
AE/ZUcLeJd4yjMHTPj/1hKvUHRHb9jA+SYzAHkth7RXN3yJ1/vlGG2L9fGSALb8b
CO958O0RLsIGa4STmHyr6Am3V938lZnG5JKPP1pJ/7hpP0Ml8kqLiLOalbOQJ0GR
2hFnvHeIQkqk0G7TsYWvrT26lR0QcsoNDQ5Xh56E+V7TpusyvyTnXp5ZpYnNMwAL
ctP/oFQciPdSGQ+9n2Gs+LLrkJlhgqpjTdFTtib88yiMqBqFczI5Zee2kLha5+QS
rCZW4ajUaIoV/OLxUxkF5AI3238zCg2haxcGtjfSNY8ze9Dhe4sypEpp4Zx/+eEX
zZ7jrDNx5MU4tBj59Wg7WnDpRjDeYFegY/L+xKHyu8ncyqgm4l/4ifjmQzaI07cO
azqCoVXfl0zWCKNP7lERO6S1Y7z+qZWZajXlN6tjlZCV65uVjwVNm0iUJsBUMd4i
moe1XXTNRdcWCIK0/YvMwK7wz559Jbjtx5/J2AAZLQ0g2CWSpOKYMtbBfkpNlFAq
of6TKWkdm51PgS2HRL4308N+qz8DaDxVZ15Kz/S2gkhCUNXUoVon7c2aXlNwfg1z
z1XpNlEZB+qA1/S1kvKCAv2+6C6MudcmYirmYBClQ8/JEkUrghJRYQelTw6VtW4f
GGGW1UtnWLR56zfKeUsXmZZrQJKzvb8vJll5eNCK7BWyB8rK23dzdYVz/9xhWhrt
OAU+tChErWY1k0vnpP9LpQxFsC+3jebhgyfy5laLqkVgCMXDhtEhWnPH5IWRgzTM
F0EhBTAFB/bUR999syKZT0Eg6r8UZN9XHMLVbjWbTsEHGazYfnMUjjfz9ZbVvVjM
CRi/TJx/APtzCP4lBySDBjB4lWy3TSbm4anrhg+o57wO9LPObMbJxzUKIWLV9Lze
bk+ukATFZyTDShZISDygIVr/HDKPDbLTmkzvI7OBkYpAH8O1Ax5CwudD+3CBZ/+h
4WDhm5niCyCvmo368CU2vBcGnvGKubQ1orc/4+0/mlkKv8GGHxKjAT8TvR2SZOqN
6RSqD5imrH3BNCrYVjY0RBxPvQ5tcqP5VhEmOBA8ELsAcO56Bk8zzIR0KazywsE3
pyVZu1v/HzFlEtByFMyKYANviYBxgQNRjqCnezg1e3TcXBKajRjIwmwgwT6a/TYs
LL2QPtS7GUNc3wB0F5dQOCc8eYB/fQRDbdNODXVzs2h4S//7n5j3QMSt5atyLdUP
c/ac/wFGX3F19nPhzWf8xKvO9za2Tu573yGNBc0xNaSzxlIp/bvKwDJaOGLOE0mg
fBd9msxItbcSfgZ8ee32e1h6YMPz7uC2oZMaCa+4NdWA+AwlPG3kZbTrHK/sDNNo
oi46IG5JcQRm9TAXtO8A2RoH3NBDktQ5kGPHTZfVIk0XgJQzgkNjn6xFNhGvF6Gg
VI7MZhzO1gKjMCWcwXR4sPepv3bWroLIvdhNx4LkgooFHHe4RyFQdbaevMatvGKn
tpln5R3YQp1LKRXg47x70zk9vFCEYxVBvv7WDzZZISkFkzgdex/SGYCNZzB1wiuq
Xn2p1+fmGQRNEWfjIZ1wMB98/G0STCJph0DP03JsLX0LOf7LQ7XUa+Oy7qLtoxnC
yXOAi0azHg47tUzaQ5b4yTzhBPKIgFsFmkBH6t/T/Adrl7wG6Y6npVIRuoEb8s9T
6IdOAdNT9xS5hENl4WjDtsFg16HPwPGRM6+cuP8338zbiTNqelHEGvzuOVXEWYC4
BYEHR9q0QGmwjvJcQg/uxLsNPBFlYgvZU6v0A8c+oU/GwkVgi1gHCSuSmLHmw/se
EcR4zS6411I8TLepMGxip8P4qYBvwD7N29cDWcg7AjHzOlay2ofXxvFtbOT2qDUq
9cg8ve2ePGte2d+hSgRBWdv6yWE38KwRwoUARlki9DikUTTLOGbxFZGNbCEU2xym
CStlw9xhAGYscW0g4ZZiq8anEXpTI6ArGy6IZBORCVeeqsWBVGpX2zCsKC180ege
aZ+qAHxt+n6mBsN2QOTreEiO9zkNS6O9ysSCLVJ9i75caYPufqLXSMoHc+I50Iu0
M69nnv88Z6RvD5jjUJmC/qMc4QD+uAUBs3Y309YgyeN528+MJs8XXkR3cxAeDmmo
rBeFPxEVKsWJGml3ZBJJMxio4aAN/nIpe1i+ifogfJ16chUPtkVxC/Me+ocpj3k1
9f/QH+wOLDpJvZaYYeosW0qpJS8O3+U4FaiWwnl/tkC0hjt1SeUd6v5CsWm5OaTR
QaYlGdAArYelzw2X5KBs0ME26dnU/PRZ5UqVcK1nhNAjs5X0VSCLZCD8Jn/bcN04
eKA/ZLGsdZgpnlUyNvH6RiU4wW/f/L9CWOQ6dNRu8cOLCOKSoCh3j1QLccyxNeUr
C6rD1XMCHJwGiuDyclqDyCgVNAlqjACbc80Ecn7t/F1iH/KOFWHOWa1ApRSyM2Ou
Ko+NKpe5ZijOrn1So8IRRC9dF5cXrZEPAArz/W8Ay0F3glgU3puN2Bh7pmj1GBh1
8FOgDLhGyq0FryrQdavvnqhbAd+cVhzm8S1NquvQpRkOKwKJTFKv2vKgrCQuNm8r
hPGo4JM/HNzKIJLO7rrFJrxhcyCapXElgdLZ8T5e5wIPK+qprnXjGvCW7QuIlBfB
cH7FuG0gjio7YwIeocOOccUOGHyWGu/IK6j0rsXzQXgbyKvT6zrAotYI56P53BdJ
5hY8YJAZC+p0Jiys3HQIq/NrOltKVMcKfgRmLx3uGVOo6mNJ0yTT68f2OUYjrsC7
ObL8NNg6x6YKEiR+Q0IRf9R7YWkt1oZh3VW2RSK2GnC0k5XHb6FjEZIenlJ2iu0I
35myHyjwzZdYHYJQIwSzi3Qsj6cBMEJJEVDMZH3FgMweyR4LW4Z9owyZNR4RZ78n
f0eYxt7jQAuHtCR+WEC2KNV17GhsIe7tVbmjvriXFUGNfjShjvLnHnMwE4fAH1ch
iVQ9Cn0BW7dux09FR4WQrnTmHkBoTuY+NFkAIcIvZ0ywnt0DCjlKId4UDx/loD/8
RSQKF3PHBjG6pnTV9F/SF3uetFJj7J3UjP7yyOtxKhSMb+VWAYiJeqRWmcAO04Xe
lZs2BOYwObRNR44hvswoX+x6AULhYk0Z/vtazSi4PWyU5My+qJ9rCR2K2y/1J5Ny
lKLXWl3bDWM3gmullE6iNnkBP9/auYxcCjZP5GocsyTCmvsDPri94QLkXnf7nPo0
DaTSf9EmCWfN937L1KxpfO6mcHlHGLgNhBboM5Mp7MLuvSg14PzF7CD+/8J4f3Cv
r4ydkzEzDs1qpCOwvg4hJB1RnPVEBpAVASjQTLrEo0JtikwhdYDCIfrA0iC2W6Kt
9WhsDPkRz/xxndWXX6+RuRY/X9h4s3Uls5rZMfaXpWaF3kLGfs+YAjAUH9EyeiD9
qPoT+tU0Gbs29sJT4udkmkPxFuGi4sCEMIEBvJ76PS/fbpu6+15EVQXGyPbwDdcn
v4zNCT+O4+uuSfkQJtbTxag87l5MsHMULpaDYcglAofS5OadMjx3rHSh9q18ILgc
nUu8XOHvbfQnNyR3oT3GenDtU8glhbVjs9MVr/m9WUUGfKEyhe/4401rAAKx/XtT
lFY04M0uJMspQjBkrupXSN/+FAjDYmwY4h2dV71pE6nP4IM2qs3xYYi4U+HpeRMR
Z9fhthl68kvFM95dR/2Rsc1st26zPeXUmePFghwJl7OaH+685DTy2YYecSt1mxdI
doi678g1pnN1HNoJ90ZYAQnjXD6j+S3i0z81s+5YDDswwbeYL2kGTQBf48Ptn5BE
8WoNi6XdtplEXqPPMUULojKctBPpNUVL8PWXl97bqxkG23MJ4PGJbaEwu+c7361m
yTQVAPWYsw6+aA23k1pc+8WFEHzLAY7772/ZSstzSED4e2EyzJXWWDimrUtJitjN
dkDA67YskicuxfVfuDdKj1qph9pWQEUKxOJm6UIeA60Mu3DHmRbxvFo9N0oQ/OCa
nBNDAkudkWD5zxyAw8OL+YGEqP8mpKyaUtfhoAqTz9+hVtCJIkTrOUiYEau3p28T
ZFH5aeuA7RVbvZVUsaI2zlqsonZ1neQl2HHA6ZPtJFYT2EbgZ2hRsGBYGzsWNrub
1KK2gyaC2xbO6IqAfZsU7g8P7A+Cg+AzjtwhbpNlhYF8CnRdhzuSu++wG527Z1YU
rfIPPG6tWJgXMaFgaL7bbtPYjcSsL+mzXXuLUMUuBA+ZBbwBKt7EQbT51HkaPPgR
vKwCOGbYJMnEekkFkYOt5XQQ8i7/B1Ix5jLERf9hymUloCNPdvWnjEV8+tEkAsRW
8DjdPE9eluqNJve17g/txw2IarSqPWxQSI+Is/aSb2uA7CUe0sE4gOTaCCzl1ior
ma75cGzCPUNa1NLEqp81d+Dd8c4QKX8OuZpoK7nAXPYo0bEoHr2LDpf8A+7Gu7VI
U2g4mnuYtTKGML87SLgpkojk33i689z+IeynppWGc24Cep98gmFa4x3gFh/rnutL
ewtbdTISriNfT8aS/p/mx9dHG2YzHwQ/5S/twHFe2wV16JB7KgRNwpvTwHDaXJEP
mb99lQ24Ng9pMIatFYQoWrsKZ0E39aPLNRVvxzRqNJi1EmZekn6eySB1JZ/U8yxA
aVfYSV7jF7tqm9jPHfaIPwygkPWUeSttktlLpqBs3BuuQejuTMR73CxWcIV+mvIM
5DWg2q2SqsDAeoZUs8uXg+aRoEIOG5TU0gUnI6pTEUOurV9VMFzYfCmLt5nU0mqr
zNdj8UuDUFoEFmS2xY8O2Uqg7MdXHXdgbeORCdyqS+kq2KwJx8HRMasZdw+zhiya
wAy1f2nLqxLmAAk+TcpAfYFwRNJn1OOxCNGrd6LO8d8f0CqRx9h303HkSmupm8ep
td3gcUL81CIfcYk6DIXFzVp0qFHPnvJAc1pRWzmMMNL3V7ci4Qz/Hj8DtLYeHq/5
QJsLyvI6Y1wjWfSoEsalyI/u5BYWTk+d6chvIAdpLiGOdfFK6AeA56uy3FCUvcTM
6DP04P04/y5HvvEnWxXXi2xXL3kGP5YXS5ARSzrG/UyyFANCgDBSGiB+crYHp7WU
XaiOKFauGd69ZtOMSbOGn1b707JygZPtgQsL9tEy1z/+dmAErHkvG/IfOioMjP5k
DUhVWjV4Yv9xnBA+WD9BCVysDpfUTe5Um8blFrgPljy0WOsd/w58ZKbkEjpxRx51
qxl1NW6UFMG3yL4oHIDweeQFJCETmvOxItPApZuJjbJJ7rk2fkqrYhDDq8B7k7Ts
RB2R58nRYDkm9VWpXj9pWpqdJnMCqKlf6fn2kOge6ADPL2N639iIxrFcfPjBrkJR
YPioN9zr5W85OncwQAZ/L0PmPdU33gKiuSpT6uoyelkYjb1BzCTspXpFCcmMuOnX
YmKL6VoQtEV4PcrbSC5OlNlbOx3h/YhNFghZcYIAIK9GmOYp/0CQ3SCSRzpAitiH
TD5SwoutcQFBQbrFhezRIOtOKZraH9G1rt4bncwbYXodJnirAt5KP+OnNSAP05fM
zVIQBrP9XBIUtAYT4m6utzEBxlPiCc94r8qRmxZoDrduU1Y4+sz1wqNejydBmWT+
IqGv0iHuDZ/2yC026DnvKcntOczffqztV3OS/ZUHsAkniNjQsAl5fjkrrwEWjdD9
FhJKYLZAeo+gzL5JEdpmuvxOIqeGI3apLt1zKEuLdxy7CKsYYHzO6P1TdRzI/cwd
+4RMkN1XxtYhggP1umO7Tc+yH4I2yRCh0AwUZ3Dp6BbXj9Zeed3WPqgx5fl6+TYE
z3mVnnIC+fzXdu60xiFZgVnyaFypvwXM3N06TTsQ3ee8vt5jrvk592OCSo2TytwI
PdBlkv7Q5ThCntXMj+3JK9w7vE+896q8cvaA95GrOLRzcRGA8/ViZSmJxiTls8qf
SZKhfnHYW4dYRVT1PvvgS1TuQ3a4ntCV8EZKWs4YmcdxCnM9aXiMOwjnmXRotffs
1loxFsd+wh/2/K+V4KZgl3kzQHt3lE+Jm1567Bwuf3X89rIYh2aMLgbV57W8FCPo
Un3SOPucyQSMooaOxAUMX+qzRneSTx2T8IdFzgjfyw6lBTVCZBsjuG8TZzAGm6Iq
TxDTmMPFoP6D2CF72tkeimUcYbcIiKaG03HxUasYA2OfHZoVnj24h9EkCefXIyO8
m3CytiJSABMTgTQwrUUUWHoWJ28i+4NJEkrpM4oV+w2m8LAc8DYNOKv+xgQxXuB2
XYnYjHbrmYc7d8UlOctHOykXtcgJQUEakXOYMVBciGelLZTL/ZSnld4eW2pL36qR
Feb+MrGRn+zaRkozjfYsLflbY7h40F+AK9mfWJ50IJmjgd784NJXLp+sp6FOtD+X
iAOngRxy9ZUegaTL9ga3A5I+C/H4ULekAl8srVx/mmxhFGN/GpLvbukKXC+cXIm3
6am5N17DQLcCbrZt+HFtwMmbm8Yv0ENs/Jp7VAkaylwNtnrZDw7+zkvaVuqw+zIq
rYzeu2WdT8sOxj2P9ytOTyz5duaRYFEM+sYgDeUqqvqIg4ubirEa+W58hjXkunYO
IY4rLXEp0qBM9XVKYOEZrNGaqhnWQfQfBX/71oNoY6qEG2uk0Mnr+FcpwB/5RlWt
nF/jq4GVtLnwz4ntXRYkIo7fLlCmOtb480KgDzCGi56HYVccO4Bo0p/KpTKhBAwu
Fwf3LddPKWuHEo2ol719SuqNOltWO0y5gi8pzqFNMqqoIaF7Z5KAP9NUQF6tFu7z
0W7jXEjYHuh9wc9KlMKKbh/aHClYR+HHtubDJFFATu601stxvq+4lNOEYSEt+zAU
+Rhccdzk0Y+MKbDuixv27kCxB2k3UIvDtmo8EbaYC5NN6v7quspK0zdMa8IGb/gG
RwQw1s6rOCmMS8sD32qjpUUUw+AGestJBT0jI29K1aAtZ8vWzLDDPfCwNfXCFsZY
6CFJ44CU/X+xR/bzhWHds30DXj4itNsuRSnGhPvqz/2g87w4PcTl52zhBn8td/Q0
9KnH/Q1vrKiBpdji4AsPn009nA9GBSmcwoDXVokfnxitwgDY0TSSQ3qpepDxdo78
ZHwSWED6rmctp0k3DwCUmGo8Dd3EEzgKBLpkvb8q3Zk/yfbdK59GNNUZ60ALKt81
wKqVlXAi6Szd2VyYYF1DLBDM4S1bW7MIshRtVgusWA9YdMpqjgQ7cyxMeVlOuhZm
k7YVb2MmTv599QOcVAn1yTXX6zGYBDJFt45YLvcEfivFutjhEd85EaoxV2KO6/od
coUu9DtaHBQqruakim6UPr3ppLM72W7Fd4QALYpXPlL1n5UlbpZiqGFilTJE9wNT
7nfHxSJWVX7MW1kyrrFPsiDkKK8jDPcENAkeiftxtzsCMQZXTIlrs8TToaPr3isw
XgwgmI539et7q6qqkRcr9a8Jxy1YX3/swhywm+arZqRaQYw8bIWYaLfC5dpjsbJE
0QXE4M8dUDRd3xOCKims7SOcca7RN0rlxuZVQqmQ309jPpfVceanQLMTC8v4Zk+7
UGd0+rWy9jzxFpUFySVRhPfKeSf4/tZVpKVNteSqqP/JN/gmzVfXZAyzytd1axY+
5KSsUg5ZMDL/XKo5MywK72W8cKsz9LARf7FmwHZFQWrO1fGyuL8IoRr9jXxn3oxS
yJ9g9PSovUcIaGSVvjJ3aXymttVCYZLv1t+uFbyr+ym3v5Jou2/SSHPaPtnZDPUc
Xrpw9h3OxCUhcd2E/Uucjb5a27LAzgINY5ao5f8iIcraA5KHFEuFLCdYnMdaKZJn
rt6SmsvoUCDveooRtVoJjyPgqFKxnsLXziQcmtP+BjiP2ePH/Bw4od75fOFJ/dEI
zgUi8cq5GHv+c5rSurY+mPhKW1MISI5rkRtyFxdUZDy9B9NJOFyGU9yRm2IjSIFf
LzjDU986CQkVajtmvM4RBEbLSaf6slXv8C5Fz/TejAwxKhFDFERcox3lPO77tLSa
CCzZ2DQ+Yy9gjBIllGCBE94tECqc7dLOKu9QeUIbO5Gy0h+etpRl2PEyc6VvHXp8
OHqlzPWLoPDQFoISiJH/k5IDvwZGfv64oQbatM4aopTwDrS/9oWkJs6a8wuCyL1I
XH+X/qhck1e/bwK0t/lIf04rOrpzfNxfG91pImjQiKKlnwc+hM0C/j5DVtmetuG0
3gQuGcUhB+3JIWBe0xt0iQIiYsHx1QTq/MpiOPCddBZ/jHYRKDzdjPt3e7SyrwI7
BwjBPvSQwF0csJXL8M3BRpYp/hhFcvswg9XxvNaje2oY2OGkSP4cgnl9DG5jo5jL
MQ0inS0+hdHPWLNb4dAGSdXhE75Gm8C9kD+d6yV/oaXjK2toLO+dhuTgQXHUfdyb
U97z50ueiwSj3OUguO0MoLNin74RQp05+bAkoAkUDk4iYb5SIyv63BR/0SfA382U
RoAwR2vAPATOFHpGcGUrosy5s4j055OkGeZ6TzLp5mSaorjKdK8PfULP2EDTC6I/
id2jXXUutQkCyd+pF28akBVlfMgTZOSxC70PGx/+OWIo+jYGTLKzklJy+FFh/p5A
7Pm6RyC8XYxOCzGBHdebZc+QBay1GUdmeWANtVlPhHt1rykDa1jccMdQGsAqWbk/
AUv8MLR2Abk6XvX4lzI09E/4uFtXmrgDZZayXW8wYbcQ3s/bVRHj10MtAVxmq5jC
yjfElosSqUjNXSlclErfbCrXSv5A0eoRu4Lo6S8eIj49IrSKxrFJcfZDTXbniCmY
aC/uQYFqKiOYoH5nll5dvu1cX6neOn2RiyiV0uEXMmYX9ko5ax4ZCkFFe8+f/bdi
BoMFVWV80TZO/BqHzXvWpuH1h3JYOULyc9AAVueQUXNOEl36OWKgbOEDHcpL09Da
4j7Gf20M+UAjEhNNNKzf25uQbbP9MklB3zc+R/X/DyNDfmC1JdgQwm6iQLnu+aF1
vfyHoKptajH3hwHTsu5xuBaHl+88TVIdr9/LPYGghUa6mNb5knyi1kU31dH2Zng3
aF5xkV3gIXF5a2duVW3e1vYRRHy4tAGe0FPrNigSr4szQ1Dd8+T3YYIEdxbk+Ojo
y0IAWdzUZxAgYOvwA9DdrgGM0CzGuVdoNsSbk6eMsfb/HfSABWlRuCEmHSS1qHPv
/r39JRC9Zs77MCqJSl/OtOFpXUFvX6PD018D9kYyt+gXU4vQHxO/DMhR2MaWLGKv
xYmy8mWqsGKU3oXV5OFW/gUwJ33dMisecGEdr6LtnXCMRtY9I2tULXrkXiBSA2tM
CO5dZIayKHB0Ea3kh5C6UeXpDd83hYzKp779vXDw6jOjDzO0kTC4VZyPq5qApIT0
NjWtgjtMS94cifn4i5QfZNQ/YidEXEuHNFw0n1GbkIS2by6BkMpOUxCvBUejPSXc
Ch49PsgMPdQ/kj1yLv+PTNJQxdQuo08RJR9bkpKMGntoSMTb8kxnYjr6Zla95Mos
VKJhK7hk432w8ZApreAutjmKQLbzv1zOdm698zwfj07AeQAYGj5R9YUbVomNBnkk
15xH/EzCOrj7SeBIZbDByM+/kxNDLZb0q7gHvwnmZTu1sV4jZHQsn7ughz2yWS1j
6w9CuQpWNXAYR5W8w/2zQPPWGTwobALx8dxzHff6gqnthbosNPb5W9cVw4TjSR2W
IvH1+ronxaJQETR1If0l8CLIdZhvvoYOcTIWUE8aTfjLTXIbUvxG8uxmJSb6s0M2
+qJDq2JgTR61JOlkqCprf1p3Jom5dBT+pRZx0but8VHKZ5beH7pcZ8xZvvIWIuCw
4Au8eWdbTOw/kBpzR/E7Ft9DmSzG25GTY8c11o1BwyJdtH2nt6m+IvPKe/6S73Ie
E5RcLtXcTrzuUPoqqxvGENyzRqUbE5F6ArtNG8Yt7FIxQw/srZ6aO3xomtlVbvTn
AnTv+dHQRtUP2oxnIueOHsC9ji1ybLNdWmTCXTPCJtTWsqEv2vgY3yQ+BaZhPAbO
htb3CHNFy3eaKQ4LnZULa88cjRgU+nP7KFWCE5x6tDcJzgq3woav2zk23QzYclKy
c1IX5v7wLejD8ebo+1SKjMtOWKC1t9KPpx2EaARqwpsfLaoDEm6TtcX1WOE3FB2s
8tyspN3s9AhhE/1liDy7Z2WFsoOo3HEQ1deSmjn472d8rrQbA8wktGXbXOcbIIz9
3jif9U82FLQ0bZSLgNV/+Mp1t8FJlYHH6TS8KLfOoZ+pqN3HqPCyo7ENKT80SSrn
zXBziZ22ry7Js7yuLWO2piWaWESm1AQ5nKaaSYYgzammCVog6IO0NGzzWo8rQRAI
l/WpIc7V4dJjahm6Smcsin1CJfnZF1U9rrxs0lrtjbD1XJUbB5O53L4EUzZAfUYB
7NL95SKnTAEDydbV/hh02yw4Fb2HWHwUW1pGGxo/ZbsYuHXtWhSThFJw9FuSUBtE
PCUvO1z3Rh7vnSitJkxdSukW1HaXC9aXSzGxY3o7c33P58sHmqGyjz8D8ffHplYW
GqmtoCKxc4vUBFc4XdKaEYux9pkAnbUtkKfiFb6AY/j4hZTZf0roMj5TLmg05rDD
OdBORYu3IJe5Kq4/aKdTCU4MqxvhMg430cRMoB58b0JtGnJpye4tZCuYcZFCH/93
dduCXoAoGyn49Z3mtnPKfDcfMnpkMiwTWHs4oxjD+xPF04yayex/R1F7B42GhbE/
uDWkJ+UF/DY4unq4Vr2eni2lK4dbqEiLPNMRtC7oKZcE3DNdS8+n9779dn2kVaeY
iENOrna8njfoyJ0wzhC/uzmrZMJ7Bv9d9zQYY5H6zaMCbpIUZxcIgqMr7F9w81Id
EBOw2FLiIQY2/mxWOvG4ED6XqbWI4cYDMhifmhypeBA/HQEfGM88IA7QIv5ymydE
DU7iCREsxylOeBUiB72ZyLaaS+Cpr62u7WOqdejQ8HL7kEy3JHKawgUaESvBf9u2
IIJUFJdBKAa5B+jGJmp0PsixymBeOOqpiC1n13/C+8fzBE2wQeOKSmzqqEW0rEO0
8eMqeq56W1OWxp05Z9RNuJkcgKpCZ0wNlhZWFREAEPmfsXwKBdz2pkpAgT0aIFxg
mmc9mg8Hl3pyw3u6qY5LWc48WP5aQ7I1c8uTVZM3U8lrmOeVhW6XegdgF5nMq/Ki
phPsqIHC0lWqSlFnx0/7PvdTTuBDF4Oa3FNCKCAAxTLu6gXxv1n1z6zVLBn8ePyJ
Zywg9F568T7vodNWbDIefF2+Yo2CTsUzdTlg94LWuUaX8RKaGL6YMxZtGMWLct0X
cTNsOeFai8L5g80zQsGJgg7HQsz3iQoTJzWWLw2/esqHHr5Jyz4nAtFJcmik0d2L
72+1H/7vS6wP/ZyCVMqDXyR7C6XnTAQvfuWhyvsXkc7s6m3pW065wwURu5I3D6Xi
DwLJKFGb3zCeuGLhn3RSH0HHTGZbgO1yo13zShr5KWsi+EWBQKQBefxmE5UAqvIJ
R7u+9lXLEYBfRDRev5q42/JIOOgA2s/fedFGnKhBzilv3GTVF0yEBuhZ/kxwT7RG
17QVqEakC4G2p0g96Yk/AFNWYM1hXbPsedpLML3bpeHmqlR6PZ00iNcpT8R86Qcl
iyt1FmatiJBCjFfYOZN4xbjd4h014ZZDnrssXTqOVKZ4xMjwmQrOTUEUwBrN2r5m
di8VIBq2L9twV1bDBzxUhtZiwabHsSW8i9hh1IkOB0DeiK6EfMf3Zbr7cPZEb1tz
lA8zPdQLi6CD2+0BAQImh3iLDRiU4o6YZHGjQDtkgz4dchOoBuox1xZB8ThZCpO6
KqXhib3sHWYV3Hb9f5MCAQXyba4T+C59xXvRe0U39mnvykojN8PBVs0TTUmP/r1x
5p7PQShrvQCuLq/pK0S1u20Np8bHodO8TX513JHwgYbeqzKrEeXJKeGe2XBlm4ln
5Ck5TBxTIGpC7eKNTl+XK67p35C0QtF3xoUsHvkQ0QhzZcwlB6jE1+3my+0+1ekE
V25233BSPO7GLyJT1L+mQOu7LO/gfrxaBa6j+Bn4Bf2qX2I/y3T9MntIIUSvgu0D
LERmGPX69har01T86mNnlalYmRFNdPg9AS8/Alg6HUKwuhtFiRGxOeHVUenHX6Iy
IJXYaI1wDmXXsl5X3nZxVpUXVGoVk15JHwLxSQ9auZcahm79iiq7aWT6w5/2MqVr
srbH96AjcKvWsZvVruwOk3oN2gbrcDgzXz7FEx8Ki7o3adYOZ/GBI14JqxjxGaUI
OuG/2qipNVEpcU01ID+H1SA1MOetcR2RSw2AAvPueRayps8gBk9rY8xgTZFov1XS
SwUgsuLYyQsFOe1J5QrEJ3CAmva/dXNkOAKylb1jjvwuSqNHO1IbuSMimMZvP1fd
TBLEC5dn2898wzwj0ILid+PY8adJcnpykSi7Af6ww+Ee3ka1gQokgjRu8Zr8FAV3
sExUZI09GRA1gJhJVoz2GFOyxB/yJc8ckSqnzeppFUEF+JzKaI70O/vD0E5lQJeo
FRSrRmPwUgBJ5NShcYUhQC/6RxvvMJ+8oXhR05KZqDetcMoYjuTsOAnXfeco3Y18
/iL7QlWbdxp+BgOxtwM4lIiw2khUFOOPCkKL9e0t1zvSAedatxN69bMnCbFeR0Uw
yHQBBkzWXQVgWJSbB2vitUBqOtwN0IMgW0Len3Jdk1WMQKUHbA6vq71yQqNER99R
vRjgpjFKv3kRoQInAjN09HywyhmsuPOtuAP02dQqt2EfcFl98xyDHle5W4tViU4a
riB461D6N2KtVAx6GpOZyzE3SjI4UxWLsko+y9rofrELr7zWopUOu+sSesfvrMY4
mnB+OBBUGEQ+EWiEBOBH0MAUcj839FD6d/mgohI1/QXgZbYHNBmYVRLIyL7rBzav
VVG8dFIPk3/q2G5gjAQTe0zwrLilw+mjvqKOKB213Z3S54r42zedR5KDLoVx6HzY
YGELF62Ga/YKTL8VY9At0rp1RAe4n8lL9Od26saRjB5L9f/bFz64WN063ZYdFMGy
0JOQV1tqpXLg5qrjV1t1iFriPpEoAmz6oaSEAarL8N2TXG2qlN7phnfR39M1GWi6
GyKx0wxiMxQexCcq/yYqfpFycTjHBs+koozPiIIPwd9Wzr8YjOMfrRUguJ8VCKag
8C696EROnBrW3Q6PmFB6A1vrfCHk4oHlTTljiKrWOG7XiUxZSQpIXv9W50SlxN+v
C5If1f1OBBEO/MrP3Y5M9vrj2hMm9ioFYPGe84sofmDPy3bwysYIc1Yn1oNbLToV
KGMzEwPfVAr4caawGI45AnMJZG+G7m1VLzjE9/HfQTnNOnrBPBa+VlP/48b0W0e9
hZTn1uDLa18L1zKJTQF8YBpp+bX/XwnlRpaJVsFuxts94oS0aelOlCbqSkej0ykX
mqd+Grc5EmYWCs5oGREIE6zXVZsQWzk+4TxzGu+mnGCnn/CuSpuzPJbU2cQ2QSt5
Sv04ZWtj2RQG6/NsxUCzypySHFuhCo7L+QRzi4Gk8c5O5nR1V4sDNgCN7WgVdsB/
7Hy1qNPaI13cD4GrhCXtovubvPBB65KwNJhfaQMHmBFXTI/OPDwLa8GTsQr5yKlW
vw3e2PeEZLlAVZszTayqqCzKaVjPJ38rkKEb21GriBWKyTv86FdbL8lxMhhWpQNJ
KvOEwxDFeLkbfHlYzxgyjIk5eDs8JpJMhKDJYLNEXUsyaBV8AjZ7WDe36cOR+lPe
RQAinQQCBowdjt+zqiEtfllSJwvEKFXQA+xNMkmAbnUlwgxxuWry8X0LOIvQFI1p
SnfTi9ZFNpQLNC1do6UBicX4aFUT+htNE+CDVA1ZTthoQP4zB5Q7gEZJ1exdhgNR
DPXgOP1+N7GWRk2cFu07ZzhmaDrL8GMTfXn234MAOUKZ0JFXf+85Ta3lRJBW2nnc
20VKafYEMtO5Pisk49HlMZPgerT7y3pDi0xNLvzHa4eHYeTmJExEJEgfbherGEFP
3rr3QZdN6hAR76NqpUND9qE1o/qBjDzO3nCYWQL92w8c0orhZK3o95NU67gz5iyJ
TuIxiOTBrwr1MZLbCCq+9Dk+/C1I4y3syA2j99tcDZkxH+qR8qdIPap9EpB3wf1Q
hfNcFYuFlhYdp/dEun7bS6ViqnFLN9pXIEHgfSt0+idoeL8UD9CZYs2+vy27+RBM
Z5Ke5h6oAQP2h/Nj8eiTdcFfoEBheRqw0Hh4/YXheU5WMKIdxPRK9GODtSb3IZqz
6Nj9NMZyS3H1j0l5aPx98HhJ0BsyNszzSaiKlkK4QX04t+9xxo6FNth1Wqyx+1pL
mDrjnuEztSrOGCy/UBiwpWh+9q98cemCm+ELvV+m/lDPJO34Gu3aSWxlyILj+iIP
oyuXLAI8+bZLTsf/h4pjapqiqs7nMnJ+PZ5CDO9UT1dt0AJjQeTdpip1Bn+wX7x3
HRChGckRzMHHkykpDpo1By2MFaiicIH7RsDhDbmPr8FC9ZpHJyJ3+rLhRkKfWKwG
5Eei9lebHXabjgPo3R7MSuHHaqAVKw+BAumxJ8XXIYGyHX1c1QQ+Ec60WZZLqwc6
OyQV0Qj3Vhc4Qg4eiqFdDHVlEsYylWNaSD4Mfvjcg1tpgPlwOwm3nv5e1FChvAA4
47xrNcv6wrWlNeh3+xKhSLHsCRQ/GWkSl2YFHENzFjVbMyKsacsCWJADyRnWZiit
JshyuGzkm9iC9OBxckf0joChk1iSsrZm5RC1NzeEMxZLSC31QdXveNPltc67yf2V
eo7FYGKQoOZEmSZ8mjUXe8IUxj0VHX+qLOlAjWMgmsj8D7cj0Y9/uZ5+uMYRdWLn
Gp0mbnBHutgl30EXWhrOAcp/8kw2UM7FO2jRshvo0aX4Rh+UlurY0bAwN/1v3Hj3
GTBVsST/XGFEYmGawkzXtasVVQFHLn1sZt5UvzsB86K+wV4hKxakFSXVTlIv8msU
mI7YhGuDMH9S6M1uzCzmJfF9hIUjcSBqe5vxV+KlGWFJ5WmyvCBq+YgFZGrsr2Mg
zy7UmVjtwyelmRMp09Rrf9lTNHUKMTMIBhJQX4KGswoq/Gd3VFZF/qGiqvaJpsnE
yEigx+ZGPi2tGucu6JZ9k/60HlcbRv7fHWH2Zn+6cRAODIDjoAExVv9cQBTNtyrl
Z51Jzo4JVL/ehCHQ07jRdaszMcOXefqxWAj+nAPxUGLU0UFSA6l4tRBr6U3eRWmf
eRfjf1/Zo1JOgYaxo/vFZXx8dseXRnxgiyoogIY8wM/2vtTgnISEkX50ysTCv28a
WrsBmz8/zqZyjpdkAIjWY6IyKYptmV6PcE56z5KpDjKC5r2+XLiKgLeORtBNEm0H
/t3YJ39fJz0NrQdumCidMjr1MUHwTaDmwnNsXaiSwDENzhdDWmle7BaKen2hpmFL
JEX8lQZikU38MCUupWmiu2Xn8iKHPeY59XyXV6uGE89u8VusCv7hZo4tYUjJ8jgb
xphLWw9ZFBkXf3jUPG3MjemRi7yJhcZhjpp7YEQm1Ibd0myA+P5AfrGfTVo4dxib
nNO1jfgvGY2Ar+hpAcHrFsvQtuhs4UJSLbwKTvNJ8ObW3cn1IWWNQTWKwJ9aUXu2
Wei0xJQfiumG3Oe8GlNs8wxH2FhAQSk4XW4Eb2TXWi9odqWG6+ftCG/6aiFHFfV0
59i1387W434II0fom9JFF540jd4v7WcAuO2JDlD802MqR6+aMbwu5zbUAy01JRdX
ygC8xcg29cDLLa1ftd6nFicD1uy+TpahMrAmK8IV/gYXUuBX9ZgmKZdQkZKi6gNT
dL7bRW9aQKAOZrcEbDWHL8g3IhseFKyZG14sg7P3B/TgtaOqNJXb/g1sMT0n0wnW
PeAc0E0BCbuRZ9xPnnxbLlwf6UNIAwTIxgJahg8fhTwwEZjHXhUDyehj20NUUbUa
vGSAFYGYZeuzPF1uuk+zWG53kKNyNsznQv0ef4ALW0epBSju/tY9SKsJ2eOiDn3A
RQFDAl4N14rQ6mlYWnyzXkrsSdcAeXNymoA74tGXMloo/jZYZSfBdiUZm3n4PGBT
rWfbx7lFEaQQ0AaLJLvcuOwN8Wvp4CrWDwT4PnYHk+ar0hTGQP4RHY0gowFn1Tvl
3Xh/+f87uACv0+O6Q+cGYVmASxWFeNyyOqUqZJqdXR0xfYN9BM7H1/Z/zYPAL9c7
Y/o5biOtx9phWzQ3diAx6KRjRJn2ipX8pzmAQENnwN8Stn+RXlW1+TExhLeCIolI
cp859xRiBxN7TA/Oy6SQkSYNyaQo4Hk0NqniYk3OESar1nsgemKfJej634NU+f1Q
/f+8KOVUUJOlg3dWPb+5WzJE2E5W4tuMozGh6YXYPdl7qVJ2Torsn3KZHk8SBf1C
ZIfbXt7PJeBHq4eIhZaGXV647FyCS8Rwgu44GsERl1fct0gz5Vigtps6DhZjKI2l
1RJxLPd2Ir+wk2JRauYtFL3lNLDxyMFzDavkF5CJ8LA2WrQ4tVtFZw0jtMJZNEDx
NoJ2pmwgSOdhli19Q7QkaQdXCRN4mxYjlsZJA05joxu4UgfXww8tQBx2oncbZrDO
+15o7NSNowiE3vYKRMRd8l/OV30kpIWMJu3ohvvvE9boPABLJ4lL0zGwrBGkt4bd
9LUbKOMt9MbvhUZRsdDr88GnFyHVpp2mWYc7GvlWtt1LuQi/sB9w4DTCp0eMdOht
B1Xe9XZReP2v6Bt4EpVILTC3Dv1gp6LYqhJvMnAR3mp5lxwdSuXNpYRrdUnPT7LE
F45FkKAejVnEwWsge3pVDizk36NtSmOBgKd5EQXO8CSdYjTWNZ/VlXC0nqHe+3Gl
zzOhHgfluBtnCf20Ux8LdwAvXKnJ3a37t3zK0ZeGYv7GG6D5WipU8lnX2zsTySg3
fUGzxKm/znbmE2KzHr39wyd9K8HwGfldBLjnc9BZ6zuht01WlW1usPFiQzhu79l9
1TjCmPqgAWlH7a9LKDRZ1PFAnPKuuCHNpHusK83zG026DvrRjc4sdMt8ezUFMR+1
Msb1Crn+8WpVlimazHHY0AA3zxySNsq9/SaetSsCAh+DWqkjU+9i6lqfNtW4ZtHq
j51GKznvSQyYHSXALZq7FsYo/EUGApVk00WW15sqF0XRfl/BAzJ/EhOLAs00KS6+
5pcJD8MAgc0pTlSgkphISfQZMn+NPsfC2JWWqXvRr/S6LRIAbx59yF9EDDw+tkLI
PVUXN6T2oJk3YSVzW+KvK4tQLhEYspcm4rnbjN2KBnkHeFzEvXX7D37a5ugW6HXb
zxk4aXmYrFn7rpidzW6/sWTGN2GEWtlczjXTEgNHMCetfMEsyREPLt3PTKXmaZWq
VzgJL7OwimIdrHhrh46buq8kY1I3GcOxJ3AW4lAu9tuTfHc6xacnaZZu7PuFHefR
BfIOR2B9E6JFNbP4g2bxWsP40ZFI0d2gZ0BB+bIhhXr9Vh3Jktu0dTEm3Php7t86
lZmOXEPyi4hg24jiiNF1yDDCgs7c92bvus8QYycKR5q4ywxGbar703A2VoRJzYrp
AOib3JoLJS50cuHT/VdkCvaRlPVp0nZeGJQVKKVzDevx2buoFxe9ZqfBnF7Z8aC1
cQjEcU53JoDBTcjlaA0Dshw60LqgYPjBu1oELroPmrU+86bOyHQVUTNRnuv2oSrf
po4ahqmx54/WBgeKSO5D7BV2vdDW5FDoO8UV1K3iySSqU7kgVqB0NvIftB/SFHJi
oF7JIDNVOia+TXpcIEv0cwkwfRxB4HaykZqNg61ew2skGTxnt/QOZa/UL2cDDLPS
3LdBUP/MJg09VhHbOEfeKcgjov10jsVJ7owZsm2wdNURNQzwsnv15XVzPLdlWxxw
AfKFSLPVdgBG7QXBFWTf2LRoyxlmdb4RnsKvOPjRWuTXLeAlqgGNqTSf2SevZO1t
D5bKJ0kpqZCwGYyraYvEuxxfVSHNxwqcsyM4Rz91B66YuKqPYTjS590lohbZpAai
YyxXB5w7xTbM/5SN1tOymBIzjS+g1Qreq94j4ixjKDMNUKevDKnzWc5BtOo18wPn
iC5lrGzCUzDHQChvCLmvbeGnbCUfbUXHn1mCId5PqLka+ou5mT2z+SP1Jtux8Pzv
OUCIh23IRH04RgASg+A+TEOtP38v+oYUeJVO3uZAQkhinxcfdVS5f/sv9SFfOe6K
zFB2cmLim4Nk5a/wnEJueuNVebC5YZcLs9Pp602+hRV28skGebQ8wM5yhgZMNrzq
xyiPLXHTm5VC0KK5nMmRPeFagikyQ0yijEEVMlXJc6zXoUbM7t5uCEJY5Aig2BKF
zfruD4XC4jgJ22G+M03nuYaeR/md8XRQqe0q05Px8v1EcosSEiAJJozAAtXbSZDj
ueWwqelal6aWvofbM/LiIGHfxFFr1FPUj3jD1U1/doLy/tLffRdu/mR0WfCbbjkZ
1MbmlzfjVs7wYGzKC8h23t/3Jfc0LbF5c1tb+2ozeU9k6b2qRWgD2dReycnqAxzq
/Fp154o3X+B3hAMg7Cv9EKjcFNev9NDnaB7EF/o8XmA9Wn2qh5iexcFkXgq+rtx0
/1EtHYieMGahmecWOijGdQOsUiOUzKdQXeiaZlEmQ68OccCZr1Blzx5zsQIyM3+P
rJ3g8nFlQwpVvSdGS1fnSO6Mdd/dX8IhuJ1q4NUicpNcPinsAZ6xXa1xu/yx0ttH
59nxj3kJtwQXXN2GN1I1LbS/EeP8HtRyRf1Uucw7ec73ofrm02EbjZXzrdmS1WRH
5T3Lj51z3EXzpQVE1RUV4l8zmn83VqSemIT02RhYWW3I0/TCWx76xy/7oJihb4HM
imeWdkk9nRylIx2txtW/y7AVwl9meypJylRkO5ROxpgH/qFl94XITUhJcKHpkcjz
jwtKAwMENmXSxqX73S5oalrZpjmA7T3GVB9u/ivwfa4Boaj0kbdbAFH34vWUZV9D
F3jvM50sBwwQY00ye/2bxPu+4SUzAIpBQTY+Ogxq2WpXQxdGcmEZmmRGba5fRxxP
mqKXpS4WHdib2JmijeZkJ1D5Ke/UDdRD1SYgJcloGMYuM5TrYdknSjqw60ZWaHXP
mBaBa5Af9k333t0AsTtNGZUD4EvHaCER9h1JkseIMvnQoOohSeoJQiUCYZZuzGAG
qAMVAPfJ/sdMWAjuWAcs0a8hBgwWaKwy8GCaUhlBCdFl/oD+bo0kbhILLCLl2V43
eSdEA3ruVU+gbs3SPXTV8nKgw1yZkElYHrsK3Vevw5bqtUQ7TlNnyojWsFNY+CvR
f/Veqg4tE/BjZSMk3ZoKb1QrZVv8Pv6c+Ldf2TtFrvplCwB2lC/jVkzmGd3MpMq5
0aHGN12g5+4U1+PptLbGrTYG6dCDucRC5/qYYMlmActkY1y4gkekWIps7MGA3kAe
gPubpC0yEIJWBflJJLF10LELe23bBNhzqkEn8B+jmSRvVS54NGUDSkk4f7vvW7IR
sMrm+Nf5r6NA3TnyOeSQ+238lHJntTtnrh8wq41E1mWpkg8gPSmRb1vev6qjloIN
3TydE1sMEr3QRpVLOPrg026C6Lfk3nNHaFKfaKfe+4w+Qj+Gc+nZbNxw41gMJ6wj
gt35uXJqbcUV0ovW++tJV+nc/uSIQBANpS2+jEafVA0LxTd38mPBHaXGL5YwPMNw
gVRM1QVGw3DcOi6VTdQNytCcCGF0NiXTRfkq1IuAeBAng86tu3zWMYUeJSqKuVlS
qGCNJJDrIxB1P6Sg6VtDqm0xQMPTE237s4nNVksHELBCbbhci2pf/Y+A0u/L584g
dHLwJWMGTxzR3BVDjg6jB1qEiQrCb5rkr5kMoZ+ohFkGN41eEljxIpK6kbUUlCqd
jzXfc0FIORMdpEGoQPIHllbav05b/tHDCF4HTRdpl8iSVdCLxq1dOP4xkIr9gBb/
3x1OyDEUFTp79/UkgHBq+13xD8UAnkEhANWTHpnHkFO/3SLKBNpuky1nTc6xKbZh
TSEW6OSDwy8N64sjx4L8OyXp3KWcuVslQR1yligopIdIMqNLZJUNHJ70fxG2S2o9
VouekwoNT9KvFAImwHpD95QBAbG20ZDtAI8M8eNt7nQHC4B1A6cb3V95izHJYYLQ
3U9ZMNvdoiH1ter2c/8/XawqAu7dd/vbOqnJcRCiwBaEnUGxufMCAaF2oolCeIaK
2VQCPRdLlCA3Hal8fKhwywSpoaRVA8bGQ4OFfxkjy+Du3g8F/pJTrh2PDa9lY2qR
0zgR2Q9ja0Ne7p6X7cDqyB12dGhMZNM7U01c4cPI37cyqRpV6SQTCvYXUrAMtRDX
43nA2JOQcBSmCzqV7zMiAj9t2mtt2dhJfW81u99vCRkycPvL9029OHD9i6f8KxMa
fW3/VrUEKh0JgEUJkD+K6WG3K7G21gvjUrypJaA7Pe7awL1JM5L249pqd6VsR0S4
ilvSh5Hzg0LuTlikk3qv19y+ywX9qoADZ/vY1dafht7smWnTVTxVFOseMJ7McwJN
tHot/vcah4eEfwIjwYsEORcJhwLeUrHsNhGsvoqJZy7NRJgxMAcep2Wrw0E/38Pf
HeSFaqSSo+q+fi4pGD+XMt8RDsANoLs9R3xjMvgzcJnIXJP+yE236aM/BlKdao7i
eWPDA3n6GC3/JPS/ReKFqcal3pmDmSHeq/YpsD7sIc95ZbO/LVEKB/B6c2Io9DBY
NwzvIeKegpttnCQcyEoUM60vpAgCAV7O5G+Uohh2fNFAPeRZ5R2+S1/ub1HIAFzR
IaDDp6KQzyeGAnQwD7tjj64Z1xUUq4jabExzY3+dV5aK61DQ2Nr8RcfV5/rrJspe
E0/uag52ktpOwcQU2FLVYhlMp7jtOAqClzFcU7wGGEe5wQlWsQ2UZTl+Naw2JIF5
kk03lg7XRTxolEU0jqemVizL7GGHkKQvRzS0/G8HDcf/NHCFvVpK5MOeO0lI8FJD
SChWab67E5cOI9FJ0XGoQyutVf2D5/QX7a8ah0ctCSKqugnDRa4vEzww3kxs/lXd
xGNovRe4u5R6fS0smaOTyJqfHAKyt6dLLgTgfdEa1u0SRPM9VeB6zuSVN9B/SZ21
qiFN7VgEIpp4f8cjPrQktGx3HfTJHGdM8nwVb09NHcPX9oA2Ggxyo+73KY1lYwyK
wGwOH/UtGSFcDgjQTlrtt7BQ0hsPblQV9MUoHjs6FQQhOjvkI19Hu0qV5Yzl3uJ5
js+0rUmt/aZFwmY3qhTiPS/g9FDrROns23/o90oGV2y8bqzU0bS7g7u6z33MMbG0
pGru0NoUEMdflH12b8HlERPJnV+nlPR0X7d2UEMW/2KzE0Tl/cYBj7cslRB/JcGv
vowG8KO0zsJaAQnhp7FsUU/fEDc8qEnUPCJFpsE5bc+qpvqrFrG7R3TfFZihY5/h
0kGV2dLtCAC6RMKSzesJU9MOJi8BhH8szFAlK/EiqZ0ZFJBmO+8uUBtJwp+UM9jb
`pragma protect end_protected
