// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:31:44 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
LPgkaVhq4kz5DcRk/bR7k2hZ7sf5iArhICqJoWNUtKXWj5vcjP0zm+JhIaTbG5j9
7+pEfQFbP/+TCV6Am2fNzHyCCh+kkZoz3+H33jxFxt3z3UaVRZ2NmMTmpg10NtcL
YtxpoWlg1BCj6fjCxh55EUjCU4g/8TO5qBAnNeN/TQk=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5344)
c3bpsaE0CFPcyhj7XHRbsXHuUBUAKUGoPg9lUuojC3+G4Ub12hNh57EUHOY/tYl+
iQ5q/blOy9lF4Llt6Qw3JtMjJqpwdjGBXAp4/Vg8nE1IiSp14wuXbW8o6baRSQIJ
rSbpIcc/4RJT1FFh5imG6ZFUupcDIkfIgPTgBlImN84WBb5cCNUUgzkSOjN2OCSV
ZikzyYr8EegXvZoUAYbfslXg+eRD0ydQRIXR6Bdeiiye10b/83qhCjPPwwBE98Vz
wVaI0B8CAGDipejkVpVaNqf+KsK1zJ1LYPwlLYNIFhMJS+JYBcY+9pkFaSZQkEM3
kdtGtn2CgQv2MtCe/AhZjkXKvUoqo6R4PkCim0330Zhs/qpslO3RhgxuFj3ji/yd
qcuO2kYlh7uVi4zR38eQH12m0ov9CzKxDoUHrl0K76rU8Jchzj+wK5nx10inLVNQ
UebST28T73xw3t1C5+59ywrpZnEt/LKJCWQz7rYeebdcMZlxUCY1zlzYoUHZ8beH
c+L0PDBpvDaKmBHlFOWIduycVu2rgTSHzmImUfGjJgqaah3ZE1TViZ99OUVNX4O1
mvuV87DDuhM6wNc2q9WyiNcZNH9T7kuP4rC00Z+qtNT0oH7W1ki+3AWZ9W1Z9kYc
TZfuu2R2erHWtXdKb3iddcwcY6cGEQeWR1iGrdoy44lrCq0OkYOMMqESVlnqxeut
nJqRGwL8MFsvfPt6EyJJ1/lbc3HsbL/AFfiphUIma/LNy+rExT5jpaGtcJX7mAsr
+RzrhOFi8f57ozGHhO6E8Jrt2JjmaEspZAPZZ7Nq++CYxgNMmA3eq04IhG7Zy49z
VMtI51tojDIc5CUQP7GVoYGnmITZ/olw3rFwegNjeSCwms/erz4lc9QGzrW6CIRF
rhc8hmE4oAMqZSeg2WtbtbOcwlG1oYUCVp+M0vIoqq9OQHiZH281gjK7mZ0i3504
1ONDarIaFkD7sR+5ThzeFvEvW/858OCYIHvZ7S6UfVsUrCYP0XW/05IQcfug9Iyu
UeL7OeJqtF/Nlfdtf6DB5OzLNksXyQFy3rakk90Ukbz2doM4/kU3kJ/gsbJV0c49
zNGJgysP4qu78392LFVD7TD8UG8N4qLJyhdaLCPOLa6/KqmvUTkkY2Y3A1rog7fv
py1FC75dLTJ5w8hfx9b1YRL4adpM8r7CFlYvmQpuBWm6ZOmp29CeP/7P4Xfladi8
2/5GA4CVm0yWNHqzqoJXYqG4qz/F+ZqA9jZ5KSrFNtP6CQj+tB+OK04O3YnIF2IA
PCOLQK9NUh7RqyhWJOybrk68PZwzB7E5nCQxuYJpPB8xlliQUPAZEH1hUoknXuxE
kJEHzcJJ/5JR7Jxz+EtY2jPJji+utLDb9Nl2tOtRSMZ8gOrIlpnBBZ8UgcWPMC6r
aQRBwVOPpZW6fw/jznGT2+t6nqjSIqo7nMJ3XB0WH4yV9sBSn7XaTdACuqqS4ngf
zKm9ciPuZpijtYYcgTNtXhwrzYflSXvoRpPam3e772won2shWXj0W0MEZZGqb7BA
7M+hdHmF8exdzzEWEhpb8DIlJi1NWU2a2c3UrFCM+octwUEjAoZjGsrWzKCXTdcN
Ex6GzGyTmPia5g7bz+lG259K4TFTa0hf4MD7Np2l1632HFA1J+cdMAN+puLUbTtB
JTvGag49VRXonEZ3XroijStpSj8VnQR0HT/7UkVeccWihI8OCinhQVUOiOemxdCv
aa3wF6AEJ8NYKu6fcxz16eoCypPoPYl9DMpCG59fK+CseL8hnCy2r8+EM6w17UfX
yvmyffgZmSOmRl1JOJqwwsUO+Z620evN3DtFAcTB4gS5pfPTnDFzut7VvY+WWt2n
AFYL736n5JxKBRx2JxzKKXK2o6qSS/20ki0ohVNnGSCyXo0d5irZSAC83zYNyIqK
tjCfd6R5AoyrWxpIznuaO49VmRKBgvP6cp3fo+VWvOTDs2/akSfcN8glFM2X7fGh
XDBm0gE1u+gad1TPAlEMBSfeDQfExRXtuo+mQxdqaYmOrU0qK5MZx7Dweqy09Eww
UPSegPS/qT6Mq1Gd0RlEckQZ7MnkbswlNuR4zcz7VM6u1TSLlUlQy2XUGY87mtEY
csjwCw8YNkSjg9H1Bfs5MuVE7czndmb15ByyiRJXg2X8ir5dECzwHuapOSF3V6RO
nBv0L8EslDCeOxeErDzK7Co/HczR4KmhMkoxIYHCFo467lEJYBo/eN+pLD6wIzLP
TyDv/nUJFX1hlvQf8fWkQYFXp6BlBiIVnRxjlRMOndN8CblwgY0pSu0RjyQHYx9W
4KhePufWl9yE8WtaktCWWcVrtz2+MP/Pr77N2qyj/n+oi86V0ZGbBH3dgGkhX2BN
pfqSfxq2bxy5N5lCj/HYCrMMU8Q3YXQqhdRjRDx+10J2aDJ/3LEmFtDhACKR9EeS
yoZcNuvWHE4q6F1Dl0oWDabTgQIT7ASwXvK8pv4sFQ2XDD/shCUCna7lkhlCSEsI
EX+VBQHlZiXJz1CIXwEixnfcLiDjtG40O4HgYftBhTzq3IxNx4Iyi4EHJ1gaAs88
KOudvsf6CXSp0evFMn7ot1PgoXWP4rQkXtJinzrWxuehXJqio0a0O3LnH5w0DnuR
hOz/16xfavljBMy2K8kVNJeubQZL7LDONUKU475IeTZWS4N7WOYsjqwCW1y2bpUp
M/SXj50i4ndH/BnWIkA+1+nEsWPwwsIveOI6p/l1T5an9wkh1FVPEAsYmrGOtd8/
IWuDFTYiOE6ZfetGfJEBnITexYUYN0SElZNGJpaI42P/T5GXnYcoXqyOedal5WmD
ghHN/bpStrqV+sdmhdvsXC5SiOXfKJsiuMb1KU/YX1cPWXAQzVw0LzpCMLbnxUYh
0SFNW5QTA8lwl/ItYLXKRRBEAGms/fd9md0jTEaMZyRGp5avlw6299Ay7j8zXa1E
ZrbOIIwRGdLpjVH0V6xz713B8TGX8m8kDlNNGimDqBHEXCmMzE4OoNNjX0JSvcXO
f39KkHOV62qNCZ0iHdG8O3rrH4odeNmR5q3A6YNno10qvnIpRNxB0Z2xsZ2igeD4
ybXMboTc7g5S2tkJ5nDphNuM5Yy3TgF2bite7YC8fP8hYRCRckrLWPIdIC3DW363
ayTWnDawa1z7j5ZEEP7PmaH8U5axtEQZkmnNpA+4RkaZlhT2dHbfnhXmr2TchmHO
7FmW0Azb0epJi5NLO8KX2BCEUc+7kW3Js7DfUOoSvFqpzUUgFR4AhUKCK1uWo/ER
kCGCIYTFOFxCg/vA1vFPdaZo0fLu9eIX+bzzx6hT3gIvyGx12I09GNpXg9mfe2Hk
TP91vZmRTEtRe5lfQqtNwENg1boZq7ct935nnKNVlNM15XlGqRJjRfNu3nDxXmpI
Kq0PL011uZOzdQHe9XS68yt8V8RbUZCUxSLK9JOZHULNrYnIiARNouB4PURqHEAf
kTjA0L/kNNCeQsVmxbDAlyKKou5hXDxx1D+g2+pJKpxMpjOqFmItbaEBXtZeiPhY
OZBVKl3syR+6I533ehIutin9UcCZib5H25CEynHT8Gv1tVCh8VISEXq/4bce8Vsx
DYRV9RmA1FugR2AU2GcIWH2oiqgxkHi7z+Ku/znYnmLnD9D5lLilfr5Z4doUgaKh
60LfuvWd3ZN5ExuUyudVyJ0rYzftV/HteHS+ufrvA3m37wJaUo/F8EPxoJQJn89C
vBofx84wcH6/nMu1dyalCJDZK35AN7UA9rVTAtB1LWuVgYJ5gJg1NJ28cc+Pq+M8
wrSXSGFN7QbLWFhhN843j/E7V3ulUsKG+Hiu/ahYOPC7m8nzR4/DB1e1r5drmxr1
MQ0ad6cAnC32lblTzwo+rXDZu271rtLXC7ego3itjvJnHTV+tMavQJnUxIsrCHtP
muG37C9TNnusLg+vtt0U5M41DDL4W7n/N6OAI2cn6t9zivitnUnA/Y+Eb8KhgRhe
c9gXPlTNXPAsuGfNrvFRm0TfFtggHp1reBTUsYRPVgR6LIoihhYtvKQTSUd4q9LS
1U+M9IPhUbFRj/5fNFOAUwClI98iVlldsJXr/cc4f5HhVvBR4K52Fg+MfYyn/oFD
dXZvzE5D6LEDdIeXjaKdk3pLY29PUgFRXzQMumonFAAjUckJKZlbDAerhST3Tkk0
unkSn6/A9pppu/miRgGVyvpEpXRZBoPu8Zf7qg2Sbor2JXZXyeNa/ZdeyrM5lB2D
CoSYRyzpRrBE4ogtdXAiMjgzO1yecmqvlH6VuckgJoxDIJ+ZjXHc3tapMwBOjQaZ
0en46r/ZCWOZb4dmcPZLsQyKSwocu6kB9YI/a6YsLMkD0ShOSg4M2Ah/2qDc9rO+
PWB0Ly0M/omXcb8s41Ql+Lju+AysAfFoY6kpebZCDmjpkFHee4a5v9arkULdWLBy
HElrh36jOgeAVUu3NLzWgI3GBKVCWvyR1XjI8AaO2i8TQUSezn5afZxzx2bbcbF3
TysaaXz+RpYjrWEah+kPKkdUQs8BWYTylSyF4pickEMPo4jg43o762+64fo2fR1N
8zobyNYun1sP6dQ203udSa0CocBxTmP1W+DbX9QL2X8NPoRr07d3OqlMsvY9ktHu
HR2Pe8FrxPWCaWyjIMiwT9oHHrJABq+EhPIsecbInRCakcwZN9WgcxOLFJuuozA8
NArXdaCbdoxaCuMomq9Z6nGjPuQoWmvdOSnZRdzoxIbseBIIa7WCtkTqHcruBIfj
7K/u3eMjlA0hlYgtLadBUb6M4CTvh4/sSO3poTPI0Z9cIFF0HI4xSkGXKCM9p6IZ
zH9AKMpAvr2/yzhfh1Gb3zMnl+16LDRSr7qnzj7e8EgP8kFp10CLuz/e/hgQ+RaO
1NkBwH3ny9HrwtvyKT7p9x/cffOMuGNONrK54xefv+MVVjTrJLtqJ3zG5wRCCZ55
aynMh67ttO6bYy9Ot3RDpv5XZJlDdjlC5tpnjq/7+K4pJrdEHZZwf6vpwon7RoYu
QIB9ZRXZ+aWYvqbDh1Dmde4+LFFRPFVemZcOgMXoG0mklLM+kEh8IP9FugpnxExD
NMhOmFLLDJHFuYAVrJYojxrWSr6v1IGk+ThMoodr4I7r7ZOzrvibSqt0fxluIwr7
pgKniaaMqs52p8mFyglgBSgZtRicgTNh9h5FYw+lvIGSbyIcWSrOFgLh9bEAITwA
REuJFoCogm3wcfvVY31s1XwI8kaAPA/W7iPL6yo/IURKjK9gAkSt4spV6WAmeSca
2P4Kbey+gw22I7jvg0/2xomFLh66l7hl9EX8WZaPElURySOpl6kDPs6hYVkg6/Vn
AmSBhm4f/6rd6J9mzMssEtut83OtsVTxbC/IPIVTj5rPQCkxKarefipdlPEoJskn
MUWjMOHfjN9PiRPA02H2HbbaTF/15PEbsaWYlgB1YVpLtZLmuCNqrLbr+DYf+Oyw
tYrrTFAXcTxNakKPHiFwzV1TIDiRfquNamr6DOSe5sMmQLx6jB5SRMZ3/4OEMueh
zCHyEcvjweYv8dtBeJ7M62IuUtukKojwpPU8xY7btD7parTdFkF85Bu0ZqGpGs6n
oN4tgmfCI87ie/AOgWA5ZGPA8etmMi02XDzvVAaMa9bk5sra5XaXQeCCXTbtI356
uXapd2CTGNRnZbqdgknLnH6eOlg0TZUYeiDOnS7xxNUNERdNa0VF0AYfqX1rLYpk
IykSN/xBNVAJO8WfAQPPW+jNwZkTwR/F3NR1274e3UI9SdFdCnTyPqVOlxIGkNfe
dQssTbQ8nMDgjUJtDkxr/QGYW3Twtgz7Ao7qeWVOemonC2mk7o7Vpc+7SApIecp+
GKsQZG1+4tGkTH70B8Og3huOyX4oitWkcl4vIe1+NCwMM4GR2M/X0eT7I1Q8FqxU
EyxmraGtCiX/89XVjFBuYJ8VPpJyLQ7zv+R1Jznn/NDUK2BCaDSN7lmOXmXMHX/s
9IcsaIWR0KN9NsziN0SOZu7sui+5nFloj1Cl2jh5TksMbrwV3qJWhqPHCIGmscI8
idoPX26l/SgJW2L/D4rqeHnnHBBZpbNbqiu4YGiL25WwfjJ3C/NN8mCdl4e6M0kY
+2gyByAecHuVaEiNJD8RivkGsvtROjyNtu5aZt66licSrtT0fpH5+HSP56x6xWCP
XzYNI3B7cNw+0sUf1y/z0E+rHW1Il8laAkxd68FxfwAemwh0gw3z4NsgEaQd3gQs
3Dpy0cuh70fOUX1rUEVRJyL5abz2HyeRKcbTv92ko2LrQACdzyW/zlltj2Yhe9+r
/vHY1SDx0VFRsvHWVSWZXXS9dWbH19PlafezK6gN16NQk0WTFFcHfX/O9Sec8xZW
0GTwvcuDm30iiIAwjZZIInA2UEJZZJBgf8z4jDlVCUXljoI2dn0q3uFspVmOdDbd
TmiYDfbORONTxDZBh+pREf0cJlMmckz2JwVf7tcxex8MpvUxst/EUXSdu/OhJJUt
ts4mor0LApbrasaiyErusGTipP2TixPAHIxCSu5zAR6YBQc0+Ehz6/NRPXxaB2vp
46gaMdfoj/bzibHhco27Sj8auQLEpNuPcyPpLpEq42aJXyFHdmjlEuIk+WzVqSiT
D5sfonWYPt17Ckq1u8a0VSCITSjQqFN5XbwbuVlLgaQBsej7wNElXvoBy3cg5LDc
yFyYs6IJDBassVx51a4R9NPjCEA/11jbr60W76U0rn4wQc6g6+saYTzOXdLdu9wQ
Nt7vsY4zkjRatkIkOXRqJ9T17LPEj+OXT9w4mSx8TX6MG/+Rap46s/es1bV93fUs
Ag6YlrUnEf09Q7cdx9KJgIkoPyhyeWazRjBEiJa3rbPGuao0FrmCEeK13D0cpzao
iTnmzz4CvibqCvHC+Ktm/+RK5opjaHHao+hl2KJUNgcdn5Dq+3V0g5gowjivR59Z
CXhBKMoZdbtWCqvLrD1YCgzadLHMm0+SURyTyPYFo9zCQxa1yucCVx/U7AdyUgen
FW/C4PAuxgPFvZODFy4QaDLaqw9bBQb8jRP1ytdM+HMnqtXjvZxpWx/vxEaxLB7U
IwXZx+qbiYuu9RGB3Lgo+OQUdnC8nB41Pg2FNU7p+OEIQLWQ+xAMkb2lWtWcuyly
yB6BS+XeDvXDfCi405U1Zw==
`pragma protect end_protected
