// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:37:16 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
HEcX4g+kTvpow/82972qKCjV0jSB+KataxhyuquSf2MEJHR7E07+nSVIxklEdFGv
bPU+OtJaf2uEiKuzu0qjar91HNhaXkYJOoAHEnvV4TFM7pmc36sTAG3Vfim9mOMW
BvFsnm1V7JIfXnunIp5UqeYXmUqu/dtrBmr/FvAtrpg=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 6672)
1SdSleMsWXVx+PU1HWfiB8subXh1Igkc+iI84bipHts6tb3MhBTHvm44rbg0Ul1s
QX8jEd3V4+eFR55aZ83e1rRfr78USY3z6KkCUNTrtSVefadHOOBMlRsQPjdTTIQO
5E2S60PoVysVks+u7mB8F1tqZR03yJJ/DHVbWzxkzfgwoc67JBPvKzBiZdf/Gvsn
8ASmmMTYcoRtNF+81VRDtdgphsUJnaWXzZuoK7QSZCL9aqJGZq7WIdkNlXJKEOfn
scWWM+Ct4uEQITAlH7kKIAWJTbz5dNBEOXq9WWr51tRBbEGrC9JBXgHG7agn3gnz
rprag60XwgFu7UuaZ4nnBYapB21QCJz//eIf8nlfh3xy+2IUnTTWFjFPz7rEz05s
9QvsAERJdRvKHz/CgALanJatvdZN8MJN4G/NIsuOO/AVFWuRy4ebkY7hjeTaQVM/
dpxSpUyaIRqL4g9kzfoicR6sI4bClmBgkQN9+wl079+mHFlwo9mAPWCUVMxLu7eL
y7+au9+6P2053RpGrXZwEGeNtj+R+vcjZiFwrYOojoXSOLgtztc7sAbrr/CbWpfW
SSPqrDCvauInqp2t1R3TyiaJpHYTHpzuAlMFZnmqGDaD19ykzMNRiF0QK96mBFhk
y8/MtpcGmXli9yTpgd49W9fbNd7VJroNlnEZMU8LYibfZEPPmhV3vAqgtwPD5Qc0
pb1ss/1r9fsKsef4wa7+0Pf1KoxqGUuWw8US0KY7rLTl7cTEUgSvLi1ECjzZTEuC
+gA3Oz/3xvPvLRHtosp4B01y+a38pPT/Adfv4sJuptBqbhxLRehIy/RIrb8G1v49
FbEEuy8OzWNdLSVrjyLiPztsUwyxOAM35BDhS5n9/2u2PuTd3wagyLZ+phwYlOkR
WQm26bTVI0kULjoUgVOb93KwJaGe33qIKWeMAba359SXe0+QTdM8nvJx2fieW5Rz
9Tgr1X9imPBBtrxpW61Qn0rF0QOVjAR7RFjHou33vydyjrBlxuzUOsPnpj9tDxwN
XR9vOvPvRDDl39ZWh8HCL1+GvcDvr2okV70K8ZSc7pRNK7fZsPcq+y9DPxn7DV5Y
J6KVXPlkkc16oqV8QqCyQekt55PcbF0IGOGxpSqMe0NeQinffc+FSpCHfCDREQ39
CDQ5cJloppLiLUenj3pTD40HFlOkHYMi6L+Sn7ZkRJFJI9RTn6szzK0Oqab6xS8/
YbE5S5mL3WnvhKNpX85tgL0MvNUh4dY2e8Ml4ksOIYYrQJ1BUUc1mTdp2/ZFTgg2
fSx5CpiluGZU8CpElwBtsKg0UFrKTLeG3hkoL8H4cTr7ZCUqQLmhLzf8nNvAvLAA
WQcb3i3O4GhXbsgTsKRAxRFG6DZKcpVVO/Ei0YgrpZ4Hy6trxA34or9srrrW8WS5
LJiGXisS9os+8epne8SxvlA49Jlc0e4EZYlphGVfkkZlNf3qndGRTzPZDamg9ykK
OkRkXYYtYQFYHwN8Z98Dkug8cj5uB/xySFr2giVWAqg0y1m2rSpC0/6dH3K6xX4t
Tfmcj19yINptTL/CsR+DZota3ZLOAwUtB+6WSrIDi+emOT2poUYyHheXSUPHXA2s
FB7JC4CH3n7G9bu06FVk5Wu5tic0VJLN8O/x6UXD9GVewUIwbU7nG3Z6wsi/Z47Q
q6VnzdSFkodhH0LJDsgvMvRlZV6ezHILO5govq0RAfrkGh0ablVRdyo6YA9injWM
LA0j0yhWG8mbwAggcYel+UlXNZWfYcl4CQcPVw3KxJBRXv8fXsks23NTwUcsdbmk
UKGmPGi+AWuF8McvyPQBnKNKV7GlxAxZgsVU9s5uZtJDFVJtg9/ebZXrYhkINkYP
lC8I1yCF0km+U6aUU2g45RgHFBsv+mFP/7A5bpL5Mox9F7681wVX+r0GZYf5QQOV
GqbiqTtsMeVjxnqHs1utYLs7hAsFxhg1rHLtg1sYQC+ot35A3Pz/nWFn1kDw5dTE
NuCevL5tJH02Wfr9oEgM9hJyNodADCCsi1Et2y6BxxWHm9Dwfy2p6DQL/V7plvoA
WuEVbGVTcQBk/BhcUXU5tNxvdrpd+uiBi5byQ9h2CvMOcQRJepNEBptDf/dgxf2y
f6mZVcvr1plLHBeyaKk8HZWikZn8MtP8R33rUekbblh8rg1HVsAySGgHxrZwPCqs
Je8F86P7Zm9VOjAnwKsRlPzxFhZ3/n8zaI3zTfha+gkwwA/QLZ3YVRZwdLLfp7BV
foI4fwvioE+sNt/nv4GQjfHH1cjjyeDr2SAeP1KBICgr8am2LfHU7oi/5LpkNd4j
rdA0psck87984sZ/pdbTFa47TkB9vvBgv0Tb60cg5OXdIyTa9nobHJTZpVizQoLT
vP8v0FKnpbCdvstZDKug25IWKrf1W0MHion/sfD+37lW9NRXHg3Bog27iQacyirr
gSubOOgap3qbobrysAIFwwryaCKMXhF8AFgFQIsGnEg7ME4EwMVjYAEf2DRNSzqr
PHhmd75AJdjvRKrHW47BO/9bfwAfo/EZq5MPhciZZv8jQxaetOFZC1x/kboQNJcA
UmUe6BXDCoivP56YO6CF/g4AfjgRcaUnFCtVrnyq421QR5/C2EG6BKfv8+bmBQuc
FzwolGJYvRlJ1QDMsLrMcRFa402Uq5JJNPSFfF/hgiCTVdlJhgQDXNktAgEnjW7s
KclsazLa1Nw5FxV4JDIvs1R8Ci0ITGfXeldlQyxQBSf3ygZXWOYbDNCGJEpslDWD
zHWMB+4CWa3ofz1zMjd+rYUhBwOiJKPrQzZL9Jdi/rKOuLIRnd3nu5cKxEqdK5zn
jiDeD9hWDAzCiLowxJV4N7d1SFkzMLZrXnovPtC0QgWcb7CtZXx4rMUoxfrrwTff
LjwEjTKjVBEOw9c7fg8CiqPF7aZezlNwyoYaftCoImVZ8L49JyA25WEomP4hHnmu
T4eLk1uPBSwNeY4YScDVd4d6/VvLWgjJb0dENa8ZXBZ/9UcT8nogpwT1LFLCA2yw
n5qy1MRxdK81ncD7yWcUt6o3hxu28WgnVOlDLaHHstxW8Ycm22mzwfEuQ7iwjDvZ
tPS4vab8C6Ga/E4w49IzD98qcWXWrOG1zX74CKfiqvHZdETjEav9ZclakLt+hPJv
YvL3sPhch+Mlkn6TKNb/nXG7y+nlKeFUC+SpbnoIkSiOUO+04OyE0fUFAjKP/tWH
y6IR9atTXTIk50TBymXFe8sN42lLk8MLPjdBWYaKJ9xcepOaqrUJqNsUoIs4K6qf
PWmLkamO5PUr6nvYa3TqnUv6OkSHDz1//FOA2FK9Zn1BDVzsLa8nJ9NQmXyO/xxx
xptVDeoI50yFovGS3t4fToz0feBSI+CK9L6amyPaxdT5hL73NLG5+c++m5mCeHIt
qZLNizpYRK0nozCkNvyQtGCbMAFGAySHq7T5OekWk88mipv4XlptNIv6E0H6BZhf
od05wQrzZIaXnTmgiRXmeIs1K21eke1ML8celOG5XV2wWTHwnK+3TVtKnm4DaTPd
tZpXcy4PIGJ4qXkgWBVtgK27k9pfcOOrhAjHOgf3IPUCllDT2JazZhI+G6WWCMAN
voXdRzVDduri4NIsa2AkbOgwLK/1fPxUrnYnadG+FSYJk15xRKPUvHkwRa7J0rQj
BpIoMRAIIDiTGXS2ohsyYOfuI2bLqRx4deAahOSZNBDIA26PXLmfcgLPDQVnf09M
GAVYUYQRbagTGmC5OKxfFAAm2JuokuyxpV4fNDl3786ufogr12e0ckuhjQYsLvkK
pmlbyWpcGMuzEDf/lT92F4FRXjaUeVwHjZFyPDjiXeoQFfLveBjDtvK7rO4DnH3H
o8o3qm0OaCFt1RoaAOyyvhcDOw22cUX4nt1H6DJYk5DJ2BkwzJp9GH/wCuOgd8G7
WCWmgFFbA0uDIMyBVhFhg6TT8SNSEgQl5aQxntS2gg1L6/xYks4fMiV60A4CHtof
r20bh2VFZG7iLYz4dkOZ7pc1SEKO28zfK7+8CjLdPK1DZY4Bn43ZpvzGdKF+fNOA
kvTFZ9hDkAr6vunxIcTIDZkuMnlofCr3obmmaZWEkh8sCAmI3aThid8WLj8ZcjmS
aKo58VgPhKM2l8d3B0Qau2p85D2Y7QyHiUuyblEtTIt8rzBG+dz7E0Jpv//Z5jVp
OQT5eP5UgzS4UPXMexyS7zu1cdBQAA56FvrL0SqVqnn3aRV/D9jj69ZcWHRlUVwm
DPhxcp6ZwUMNvzPd5pmzWuwvjnAmBHZQ4/MJUPKI/EELRJBEk1nVVxYRSoGcf7kl
0fJC9EDCSwxSz4guEnD2Izm29KPIg22Gc5PK3kHrY7ijG+UKDnkl7K9PqEQ703ce
6pFBTpy6TfA1mGIc3Fo8YnNPb+7JA0zQMkDYyPTXFHtROcy9ertCYI0gFy/TCaT1
Vr2w4YhrP4XASLTjHvHtZ3DF39WiYXLjr+8RmCHSBXBxX625XI8dXcPv92kIbX4v
d4KhfM33knxbV10ZFMFvsxrUXpNzJCv4/XjWAzOz+cmcQwyd7lYmrmifTTeln+f9
EaherfIuI0YJraSBBRRYe5wPB6MfGucROw2JbfO78/nc98jyH7sXUKvbquko+3GM
SwvlKZ9aK40kVqNTDbcBVL7gcVT/LRYBd1yP0cb/EcE5EdWbO12tfk8XP+6cA4kc
h4pbxdJmhgo8UsZRceqqh3pVDJQWBw3JKRQX1K4d9q6KKJS0cELcp+qX+JLcdAKB
zIxc60fFhl+Pr7KtphvZzvZllbWwVZTwRYbtjgDEpHEDjIlZTk0oRlZ+/Ap8zQ1p
4Q41aGkjh/WWkNRXh10vDehBGCLyzUPZ/4ikfIv4ZIzJHoEZMBodv4Cr7ctY+PM7
LGfIPUv35EUdGGWqFyU+It2a/IZA4iU4mx3nqrH6iiEaxtPa2QVgmNRIT2iYkrSq
pRNcohXiT/7en2SCxpPf4N6ALmi5RVFihMTISdSGGV5ZoNaInTyjGbUVekPMWfzR
BZ1c6JxV3j+0PLbDvIkY2YIyyF3t+vkIOonBWQ5weYvh44yw7Xgc0AHl7Mb2k9YB
VuVUq7ATsl2YxmWMXgK/hZ/eKDFt5b1xewiRdKAtQm38XgXBy84sZ4vfBmUlrDCh
s1EpcZzNWqCrKQ//ePA/+WD9tVwDwtxM+CvP8tvo0sjJWbTwrBcNEkqNly64YRc5
MGw0Q5OMDWoIo86nYwIV82HB9vz3z9sltjWpbyvyM3xGXwHHkCe9QRMskU+uSxNf
ZITt9tPyLVxtj6HIbZDNCo1XYXOPW00zRb5crKWsajpPZ3Sl0RUX4tDo0KtuDn0a
8hLiNRnIy2B+acjmgDVR8/k2zxGoYrH0q6W4YUdu5BPQwd4wv9YuGe1T/zVtQAJ7
zJFNtB1zcyEtNxHAYonRddGiZa5guOLKi3KZusaHNTgOpZ2HyB8l3IE/wBwAkFZL
tVzpA/GV8IN8N13mZ6RIsbsSkol1y2Aybnl7beso0oIUruYPBdGSViuVrh2hA2OQ
EXNkTsQskvrCkx4Z61pnOYMxNi6Ar/dhv3koQf5MqhHrzE1nCjFEnO2zrZ3/Ku84
anXipaAg9DWyThmgGkk9jYDiufO9NxKUwFayIKUltOTlnCsn3u8U0N+qy2e9feGd
f8IeU631PC6k/RN2daUPhQAvrjgoBHdNPoOgCBipIxy6gF1e4iS2w3nd5kNcBDoc
AdxB9iQJIqsMtijH+wB3cSoJOyR7w8eVflFOzYXofa8nUwtJ1Oc8KO35ERAl0+m+
W5KPA/LUyYAAH5kb6D+p9GUBKG1Xp17MGNi+4bZI8xJwdERyweJkz3zYnazucwIk
4Dvp3Q1VPF1Ij0zf4cwnhQmDrwDQpPRR9umhw/Mw2hTTF38j7uk+ctT4L9PUIyMm
7n7t6qT8eW+jlGD3d0KiLDdsrwcpE7N4g5oeaBPhnVxVy6vE95HNxtGjhJvoegel
7tHcWabpWhTg/UB1Uo513riksl/OmkFAAetvLuBFMLev1+JgD/BWABXTSueZUN4G
YEpM09D+xxFjFWXedblTxGDyThly1Ydtzce+cAAgIbwNo14uDaoSCJ8wFaNZoHwW
aYwNypDc7mjuBndSPpED7aX0dl80jN2lqw/QJxavtTwiW08ys7+HgxXryyIimI5w
LTS+7u3mvokctAGVhzcdl9o/273BQUMqNabMKs9LkJYeRTnORIe9r4QJfhU9tNA+
f0j3bh89V/g1NLiJRrzU0c+oGr0+BTnjXBlA9k48hpV5KdU3RyIbDK4h2e1wTK9D
ejAt2+FcTc9fiYfZyDDj851JJuezZJD8ZICv65BkYEtazK8pLJrwkM5vWM+d3Ubx
QRmIwlXRgDPCrmBgBCF8vcYadB5V7OAEAWUdQbM8/OJWEy3p54KF9rrS3PX83Khj
O9M/hTOtZYCjb2Cd/jLsTT3Lb6UQcxvaTaHbLFizhsAPPa4Hvf3PsLLBEKSNbL4X
qppyxwu8454NjS3pjGGfbKDOqZIRLFueMlQXUtfM/GYQvRXb+fDSdj7QqENuW3q7
fqOvaR7V4K9uS2nFM7NfLWyZS77JEnTawuDKpd0qX4x3reRPfIlJ1hdWUJSj9OId
n63rTLbgx1YCyK5Yew/5nROyMUO4Pr9WH38lc3zuCaqDwfkFSJ66qNfX064sE19l
xtpMaz6iXiAzov3RUbkhuqiO9X5WyGbejaRvT7Rjh16MsydPF2pg+xea68zO2Rai
TRUTk2apC0YJLp0+r/OyfhlyGPqa6QwFBow+A6JO3PuNW48xoM/F1Olp+TFSi+OJ
0w2QcJEDeXpgdl8XQ+7yTIciTED3fBwKhSR7edKnlvew3PgZd8JVfv3pu6TlqV62
Esuo/Wzln30DioIcNSUkCbeJgHppjSYTWZDWznLMRkIya9X/OBjx2mS6DabxKARq
ezZg1AiZu3TgHTYIuAd5dSBU6edm5CmdtU86rVAzGcvv8+WeKAk8JjgXKwuuHEDu
kx/Zez8hQXNaExOPBB6Bgw6FCVoCTad1yxkd/uYxisjIVB8rUjty87GmPdXw6an5
eyUPJ3N0bPCmekWKlNy9Xkw8uoGrTbw83BNwZwUp8bVG/YV4y6vGnJ3xIYqajcGx
SaXGR56FuUHXFr7Qs99dUIQ2JFC0Ol+snoUa1X5fn79ZIAmQ9X5AbQ8NnQapvdV1
/g6WoyzwOEVSpQX/wAwjU4g6++m3QE73kiJSCzcZXqRemPiGckqB+xP1agzzLEBi
7pepXUgdMbh84cekl7wO8KPOj9cAdh7GOlhZQ3QaIidhqEk+CAjQ/VSzx8Pz9G8h
dyNISAQPy4NJS43MaItToUCRqrNOHPS+lXXmwxGNm+69GMpK4I4KMIAdb+S34uYr
uC/QOVBZBiig4gHWdDtFvjzZgSSQ9larLemotvzd6/2GBLa5LoVH7/4h8AmetEpD
8DRiGI+bSI5aqweWVMunCQhyhNvOUpnojkEzXtiPFgfsd8gB2OGqYgB7LznCYwdx
ZQ3Gd4z8UwMNK4hGg549EwL0LYjj70XM70RlLld6rAesCW76ftewRl1+Q95ez0iT
eH3ts0vyOf4iR6NBtKq0+J9RHnXySeU/O9hUoNKU0YYfNiUuQDphxK1wPD9MEJ2k
Op1synhaYGvFnKBRIlBQ3WIzWnQ/DA1JtlX+aerSZodWneEubtw/ieXpNIlJ8S9B
aSaqypxjRKPzTqd8PExZTqflRrjfKKFV0a3SEhJIfKOZ+PQ2PPMg0duN/Lhrgwfm
OzqgIOMwehhkjqBQv8SxIfQNs4d42aMGf4oQuvukIotIDDUtG0KqG0fuOBNyX9//
3g4pfHbysjrLLRC+dFHmL2miUAtVVNJ18MhKq3dErgYvACFfjMxRjriVLApJiU9r
isbTX5d/9pElO3AzPwaGjmlesctJrweEyFmIgVd2i9MfzQvnkWxP5fSAW/D8fg10
4P+sBSE3WAcNiAs9jybt2MpOCE7Qaf1n6qOJGKlW0WGN/rwy2IsGGtGa5Q5xtVrr
WQGQtOziNOICfB8DTP6G1pJSBpTZBbEof7QYh/cWNRIp3W/OoVKFj8ONzeQ3nC8C
sfN0o8Pr06/oWhbcV16u6rMcelA9DC7tzSnHnRaVBBs9XZhkKJ/Eogd890qTFcOz
nQJ2xvI703cIKsCCViN5dU0UNpKyDHMzTx9fL4RvsvXvFKu8oguR+TrP0mxvtKW+
r7Bu6LjExdl5r/8lN79W6yr2Py5bg/NW61KVYTzRZH69rXJp56LEyvDToyNlukiO
KzPbV0IRoUvy5x0gsxsgKs9ijC/QYrdUiXVgg+huRSha6T96NFmINU7kDDTOsubp
hMNNcYpa/3w2SpYUIz85AASE27lC7vPF0CAxR0id0PoIQLrPQKaQvuD/P1eX1/qY
pZK9yjUx1czAyQUmILDqVINUf4OgBouesaxaEoFIkA7hJrlZHJ2XIet9x6+frbW/
bJTa8xr4La5NPTaghnRiraKtLeuoJcbr+xXre3KSbuRdUYDWn/Mg6XUHG9GZNxZA
ZmGi0BIrv4L080MqvjORqd7zpmZn5lH0IrKwPPgXI0jTyN3zZINxt3qYvm7eRle/
5YuZqOe+5HS9dEmQ4Q+mvTg/frsKEFVLgQI/fi/LTa+X9e39gXs628590Mtdn1DW
7UZHyLXj0aag072LpP49gDpIuKI4TaWRryGevIFYi+7DIw1KnaHEdUqsdYyccxEK
VjI5VtqZbaIrtGg7xKimzo+6QEi4UUD5xiDV02pKzy515cQv7mno2IvUcvWmJS1p
2Ot2ftzoLHU7oXkUQdquOhNAwrOvZZCMRt6iWwKainBhZbEQ0/6fwJr684GGEglF
W0rTi3MM6a6/rh+uirrnZxoebptVh4k59NUdmZeINjxBmBZe4piXpnWQj/8T5gZ0
`pragma protect end_protected
