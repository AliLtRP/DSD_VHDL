// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:49 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
IqHrlzjnt20JU8BucdQ0JxBrHtZWkdvHfAxT6xUL9dmVNjgaX1REcR40w6tDqsmf
UhEK98EA5bdsTXdcEIbamPndkBZF8uOtupo7Dxz3dsXS0y3s3NfIi5oZ1NzlEwoF
BFF5CdtYg1eJQ+7xDsC94b1CQosTiRn4qbeTvxmH+Jw=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 9168)
ReI2m9zPHggdtwTvjBjmX5Eh0nMltDWG5+XxLAtpu3GV2VxNNcs9/HlfCKV8VGxK
ydfr5OBxDWeEJEL+3/ywnlK4veF+WjRFF92iL0bGSTXEch6uH/IulxWHDG99Cbew
p0CwT9o4E65zx8bQ2dTPRV06WeRwEfHwc/NZsJXnm4Ik9kVYB13W6GKpwBmIe3Vd
krZTWnvCsKJSI18vYWPsyzlVRqwj+2gGxpyJTulUIA1d4amhcOfzgNhUkk7Cskgy
YasKvx6Zlgm68vGI5TrnZx4VBwOU/kZp7WRD6qXBtqDxiYWRhzgXzJoKjjYll97P
mcz3ho0Nh7z9y+bt4B99co4emvjf8KxlRaVGsyzKgd62ZJvUZVm35WSeN1pxf311
g1QmawxBW0eLkudc1rQ8Wp5DmRgnMELhSiYGHuHk9GafQwKVm0kb1I3ieQvGVbeX
TNChaJgI86226BzWR6rMT1CwFduhy4CppIEh6Ix37WVHG+mUkJIPmtcIUyeNu1eV
rediDGcgs3f758+1OYKiyzp/XkrVB/EKbHAfdFTO1P9jlyKvh1xndm34Sn8lXsCB
O5VUGr/Ok/Dy9eGAI0tXBjM3CGn+ZwohVHruxRE9kDmEYOFKKgTRNWVeqyD0lmSR
zqgKMeL+mB9/g+R6LT4FTMVUaIapubWvTW5VVAyx7V5TEs44fSGUY9SYZJR0J0hW
UlrG5Gqn1IoVO9ZiXTOWndVdqBX4HaO1cMKLp0cgzwZCFUPsN3e8TuSUrSSzMySq
Mqp9to8m1cEiZLLagU1OoDZ8RpbLl41duFCJ6p21cCfFotAB8dFoobcrWWDZv+pp
SRrMBlxcSwXoG4r1Goy46Tr2Oap40ZqbqS4I0ZU8ML8rlDLlGLIuviTgQMJ4HvIA
TTmqEHekywPP5+G+/3WCJpYgVf57RtPEgar4ySNFFRCzD1eCvssC0Bsdehjn0rP5
b/S+3HFGI9PwrR5LkYrN0mkaHUFD5/vKiLqVmKwJWIc2sZDIuoJKaOH72FVrpur3
3f9RHxaUSkvyitklCC5PahVUlbfmJ5yeo1HzB3UFDVOjnXn9CHgQ6FmUD2TGCN4t
c+QAdn3d4QnjVJv9zXxLN11DpjqsqVieAx4N3KdAVRY2tWmrwprvGYwyCd0Y5ltJ
fQTMf+ojCiiFVlK7pIOFxSzL4kzJyWcj9dWskz/3Hyr7gu1BQhJkN1yLBzGYSdtQ
XEYVSig9IfSEVqbQT9iS4h590JY0GjUz1xdoAZlDa7xFKmGMie2PVrYVITuUk41X
1Qmok8CUmQkqBoAvZMitlSfezdkZfeWy7TVP46j0p1VTCecIxXQZRg/3gdUtU/Ck
KFSqDlAz35hLqqACbNSFVM1ukB3Je77KjytBigztYE1sJlFQj/QMecuMK6MJM0p1
yRBdHZv+7QNW20JdqNLT6oKUL+UFALW1lK1Q/JziW8WymZXmefNpwEF5azK+ARTO
gLaPZXb+PqPo6SsndIYXQ0phigiSyMjxqP9RWI2+UtjVO9g/lEahf763ZjQQlpAX
K6EMH1XW+IovECEDtDrPkLGA15k5ev2pKVlHHUMg4gETWIjdRDpcsowt+enPpeRv
PvV5RKnuiCbvwoaoTnfgq+IMM3oY3P5iOxSRMoLK4uathPlC7WmQMxek7awhCUX+
n7t3mrSAFmM2CGEYPR0m6lSs+fdtqtgEoy1UYrLTiRGvXMSW8/2eYmVCNiq3JjOD
qllXYXHXiJoFGxhmswKKmuKXkTvD+yuAMtKxvJ8Xx3DZK/5upDPuaiUNhpfX/7bd
GiwtwuNT7TZ42kzdOJKrvzUOnoggyZ0WgY9CnlSlhw0yPZOn1Bvrw/66Pao+WoUp
xx5k3KmEfpLOjaxSZ91RYsvZy0G5x5gwVTZmf+MwI+vA7cAaKKITgf8Z9lGzC7ke
qUxFvkYsO8kN7Y3BfwtUfTJLvewe7M3zQIw9iVEoFKrSR2I5yy8vr4T/pEl8NS1r
EvnM+F3nzpe12Vk27mKbipqBp7B1mb8Htg0ki7p1P4eq6ZEjX7aTzBo3d+33rU1W
HNiYthf1gRinbDC4S7hXxxRihNqgKybdtqTZOlqpw03Ygp2fuqn9iM0zP6nc6zW+
pZn8tbDf5wNdxvYWgf/kQg894twnwc9Jw3vEvoahTd7oJET/cUTw/8RGL7gW/l3w
mZj8ycwamaOKLm9vGANhqxY1iniEWRZ6S4Wo9q6dARa6Ryvo8EMx4xg7wLv/+IIh
//8/Rz6pINhfktW/MbTgOqctQelSP8ZQy6/uzuk11M0RJmhmd4Tn4Wyec+MnkL07
fSVDzQbdQKHr9Xc0DDk+v6loqDk+dKPkAOuNDN/Vpr2uG09sWNcxCwU6DGK1+TMs
c1ODydOfly7+C08IkVL6ZrOqtRjWtWJG80oenM/KiXid0La/oIXPaeBwG0Xtv8O6
0ev56ARUoEWl6SjQzFUtlFvOSxLE28fcOuOfjVpNN4DalNJpSgk6xF4OkL7oF3TG
E9+CH8DY/NqahavGiR71hSYWXgFsTijMrn/IR7E6S1dWJbEROzdn5ioibMUI7Gu0
6D1zsbuCE8nDpp41r7XVNtYeRaxV3RchvngnuO39RvYmWTW8NgBWCm/aEW1SAMCQ
OxyRipXfFefuivJYDK18Bzh7pmdzWsOrw6HGAmOLVaCyjDw5BIYYc4LJVZEk4l9D
AGLxWb6Pq9v9ZHCrY9v/iQ9MJ+pTefRbe7LUrDhY637N145vmfXtZczIb4SRFEy0
O5HFjeCSpxZZikvmNN31ww2+u5+Vn4rfUbOV8qCcXT0CeUabnhEUjsgqvnNE0FRd
vOJp061TVYY+RP4r5PaQ7PVbsLP2Jlv4yblDi5Q41J+OfeMN1hYuDeNMbuKF91TE
BddnZO98tu6WaT9i8r4zShhqOmJyQJGOpfYWvDmrkPCO9XKqtfmtlvfO/jfHxnXT
cBS9NO5x/qFeL1mY8JZSyat1tyWFRKTWwQb9IHEmuoy0ygfLIog7fTu9oDDbxarJ
EkIz6Rfqk8OyyLBVAf4/rsZvwtoiCbfFsKKnq38kFQ6MjymBoPDsgKoQq8GlM0mi
5TnA7gMDYuE7aUaae9MRulOe3ONRkGC1ueddI/2/aIZgr47+L47XGkZ4Kw420gzK
TDCVX12qbBSMPR0AOzj7zCBMjKvqF15QDnLIna9MhQwV4inYjCB0aLzG5K6m6GZG
QBqyGt714VDlYhz9NJqIUed0AK+OQgz0E59Fp/5c5Fr4PHmjGAllo3vriINOUwB1
yFN07Yn6c+9kezM7fl9RO5juTnxCHQAQwmfH4L8hihL4Pf8ljvmufDvHZKjIEh50
NqUzR/idfB/23/uJkDLvLa8SH1BR/xvp5Q1ARYmUNN39fH+13ScbFOkOTWwSWRcF
r3GxzpVcELAp26fFcjFFQ6hwSbl6jSXTD7dDjZ192ngKVlfQ4qCxncaiVtlxWrCx
cnrk7SptrFGKfiBNG7XP1GKc9FgATDz+9EMJ8Cflp5xPFZOPmZyhpHlZbwhrqX6X
qSuPl3amf7AkcIYR4i+dLG4eUa3gyFE8pfQ9PELsOkB2dfepjZCkvK2LCDvjICIw
/jTMocMMwzJPqipqSg4KPFmSJLlgT4I+6+/dgwtAGjgWhpaLezI+NBGWe6vQZD6X
ez///3vMUzO+O2gQREiulSsERQEi3BMw+Mv3W/lTL97Ok6YnD6Txmg9TtO4V7J8D
SKURhTnreHxT8tvXxiUnPtKqK2wG8V0p7zA71Oz8DgtusSowBW9P/1Tvof+/sMq8
4FrvwsH9vFb8TJ3oZ05edw28AXqA0G9CqKYlzMUwxAixwOenh4Bta4jZr2MxevC1
a5X9GBPAmTiuGqQP2YHiqGDukwgZFd5EeM0Qqmh9/uEHNGYAV7raVQ2JgkB+h2YA
QL50od29bo8RmAd8Lm6kQXlj6qRzMW87FX23zQZPJ0gQSs4mBXWfpMlb5/xR9NxU
71daCNTxKh/nNXOJ/eMQlwzKGqwLHmMr8zTYzh71TcrvkPebQ+vyKGjjt1C4lQPW
7uNByI3HHhvTrtTyUzPHNrY5+OXYvw3Nf9Gv5AP4XRVJp9pxg6BDDoOlPaeVMF4l
QT0SOW1p6GTWL1lIS7izO19yACt95ybNA8PrSTd0O73H/PIHRMq2gP4sC+ffvpuG
5NcmyKQAoamoCTzJyQWyadT+xbayKIZtcBjhj1hTIRBIBhAJ5+nXJJaXN5eLnE5u
L6VZcl6qOGW058qCFa8wkJimasgUfUF4hKy95oSpNoeupk7ug7lWqGpTbmdVxG+J
e0LTNQD/GfFigQVadfaC87JPWmOYKtTvuEf66qBOTN5mqf4sHYlOMoX9CQIdyAFq
1/VujwYA6zzfHitwI1B7d0btfBTSB44HQqoK6YfYStLN1h0otfrXL3D7i+8IH3tt
JTqTMJeFBVz868sElqCaaodVaC+gD3kZjm/dIivM84SMtKLcUUnC08auR/EpVSzH
R245WmglbS2PPCX8ZCwCyCC/BBHA+nfi1U+hU5gXeAgApvWohjlH6cNhZWzdmX25
/LAbymCLMrKGGXqIs4RnE/eQg7kMspyzdIsc5ZMFkOLpEr3m+CCiE/St2qKMgV2H
H2gzmcQktnU8j6xlCy+SSQTBKIG3kw5TdQrPCCDsEIeP78IviACUis+2bmtthUPM
BtQX3PqBrvmz/2kHO5qivOZukS0mO28iVWk5gZkdzcuFN0huCCRqetkK1LBmyiwB
NClqGQFgGtyAzzgxWUfb71MJ71oMp7aEcBL+SH47j2t0UH+3l1Q6kix+uvlPUhfH
OIRY9C6hqSW483Df//6gd7Sr0tN7hpTLexqgg+ji4BCWHigZKKGch2Rr/IpoIRxU
dJpLmxmJOVx0LBFua4lwhcfjYuDflZdQmyt1aghdeW1e0NUQrPPkTtXjiS+PMDAx
Kq2ODrY6FG5N4koPSz3ejrnv46bWl71LFWrB70Z0DkPCMqLTpelOU0G17Q2NlSas
ngzYlzG6JOmRRKigbp1QZDAyKFsD/OQXcNvRmAgf3lnXTuLr6lX8DfOm7II3Yakb
Gx6wOmIkeyC8Y5mClX48+0QIZVVOwcCWE0fj5+1kfxZpO0Gvg2/JmVvjwBObfuvI
WeU2kEDxK+Tl+PpTERKUG1i53NVvglwYc/ATqOFGksLnHJ/GmjC1bWmAbnCCvLA6
AcgZmyvaSbcwSUhjKCFIjHYLNN1M9EdZDzrjz/U1cyY5w2y5PU5miMzs3Zi4rrRi
6bsDUlOkwrEMcv4gqLXXPJWc0kZT7dhY/11t4cw44m9UYkrWgDWhqWzUld/kDSB7
R8CtheKS+OD34krmTSYHrW6xQjsAq4IXEhARo99ifC8pQc6pz6YF25k/Oxc/SHP1
n37HWCacuLNA1JM9n9YXmJdIJ2aE4y2GTVYN49uoC2fHDPeM32qrAPJi0TglllTS
OUoUnOWRN1dNVB80hv8/dXyDLf3G8jSOvihK9schdTjo1P8ipoVru2XLf5lZ8Mfj
cwSdk4Q6jI3x/0y9zwtqDb3+KwpFCEdjQaIFk6BP0mwj6GqKBh2z4sSEUbhsiuoS
PsebTBnGMJ8Q1SFG3XqB29JxHlNNkN1+bEjMFGhEq+gB8xQf5UbS92XkGpArS0yX
rVD0ijtjU4TGICF8DTzp/L43/hJl9N0oPEvgO6yOiJVreipl6RnZPWYEqanmA+HK
YmoIxi9tFtuBuVQiUN4v/f5RGtgxwB+27zxJUDXb9ENe42eegJ+G2jkbRDFr0txX
zmvSD5/m9W6OgfpecaJAM9MLEjuioWulEmvYOMTMj68gPNDVhRT/vMhCV8UIwK/l
nQMAOE+kOzYojzfHbYz4icpSpPCAmuPEM0KrsO2LdgzK9OA5G9IiwJ1/47JaRcMv
6O4VZnzLoMWhKvV0WIpqf/JQkmA9OraslgC4v0ex3bPisvIfA1VkgbSOfmiALQr9
tf2ltqZJFBW/T5SNF0rTWzyYluhIsjJayB55C2idXC6m/BY9CYPSI6AFW9ocw6L1
VquUKQVcPnubJ3rD+SjE4BjI5whWUPEs5JUFbSOJUYLKl2qVGes9Nmqt9p/h/uJC
XByhvImxSO/zvExRKkaIzeL5rcqBlIv1HDSZeWEgrOvkAg0NkrnUFitLRuC8CwJX
sPivZzMfua6dRVLXwLO9k/8IRFT1VTHJSSZIacNRLI3/qyFGZdOCOHgqP187UKWo
vHXqeA2hFTKvoI9aWWJfhU7KDzcJANZOPHNVS/JiBRf2OiQOZRkDkI/WByGOkDF6
PZ3lUBi27gZPzmwozgEBpZGggawCyaP1NIfgMHAVwkfh5QYAxzunT90+qP+9MSO9
Bi8AMsLzOmbKq1vYlXuRZIzD13TKMtOWBkZlXEwfIaNaRYAA/y8YGG+a3pE5uanG
4XFSydsVdovkayeXTZzHu1Ygt6hr0onGS5md7vYPBj11hxWu98omjTwfStBY8hwK
SyDuYGdijtkq6llXQfUWTVuUKiPKy45Jiow+q283vNBe6DCQWrGOdXz0GeNcCJIC
OPPsJzXc80uFlf8yG+wdb1HrTWeuZZPOYAfyEpkdJVu1srUhGfU3CltNuMhcGRck
Ypj3aMz1hx7/Bb5pvTB/fcH7Zw5oPXBCs/qZdJz+nRDgNUMGkUKcsXtcn+3f7O6g
XkUSuMI16A4XXKDPI6R3uIf49p+7eDRPq66wD31+/wpLu+VTMPE0FUlJ/kwDAe9e
7vnD4RyFPf1N9EKD4v21XGPtlWKH8B4Y/VPsh08rohsJjT1hrZIm2GZsi309PQzo
TJe1JUpc81+xqQ1gBEqeFkfaG4VcNfD4jY4/Fbz7ksXvFO03EUwBa8yoEyeDk4Vm
+qNHrwoRcXu4c45DXh8cN/vXltdgwSx18NUNXaZRdtv9yq/Qeng5q+PXyi9vHlnq
4e/aqxdRlBwHPXgrPQKq1GwmGR9FlrxWdwNTnOMMwPH1Sfl+5z2p4JjMH43AMMd0
jimisYCp5IjVj61HN9FUaEjXGgjp4dyjWqe6C9UeH5wu+ZIRoHvSDX4fjfPPCSOg
CXcmXNNMYm3DTwYi6OFPJ8JMEW2HfOYn6lYgOrRFo5HHAfTWvdlCBcBkUINgM+ld
20MsPN4aHmZm4AksmEwi7tQ3K1GSf4Qiq58eUvzBXSmlkMAIrNR50uNMCRp2I2wO
Y97BLuy7HlLcUL+KWoUnR5IxXL64IkpqciKll3ZgrFyx0h7dHZZe6xf495cskD5T
Lk0vYCjUcLASDRSdrcOL3cdbokIfQ9ZgqNVP78oxcnRk1ENlSHTbb9T+S4YYcSe1
ysEB/E8l6IdiNYtMQyx8NCqn9Kic5LccbvHG/SY6S50/ju6zc4LDNtn0eCGkeVt5
fcxwUQzyqSdHTF8pBl1KtqzBlQuJ/VIDEkQ/o35D7xuov22DBS3hbKannYFrB7Ed
JJOEojMuogqXV5ufDtVfcMA0KHS7uZYJfHJlC5fDiNfkWErDEW0HJR+wxD8aeZTC
hb+DmOZi7gEenY/aJbkwo69/d/VI76B/v67JCtlZUKosXfjvd75GIcL3jZcyIBnp
alPxQJqtXPYHnx7qYKC7zUH5nu6lVbx2/sX82mlrdqRl2xV7rbDamIkbbNWjhMus
wBmeNzwGJDXv4f0Vf+IlnwBvyWYk1qLSQEObzShA4nUttNO7E60y4WLTrN7NeZxx
pqoooMhTHEKL8xieOe2gapS+6Lxgo+GzSBDSHEtnO4ddJKY+tkFuVgBqAk0yvg52
v3YoH+tmT7/MS644/r+XT8UjNFGGgKj+FRogBi+38b0EF1sivAndgXZKwYl2xSmx
OaNclhwUXlGveB/MfEYWCMWJyTViutvXRkYq1Mv1ntUhpOOP12p1YBA+v9K4j0vh
F52Ztlb1big8MZTq7Jo+KANxnOs31WbenmH2T7aNZigKFsFyT1a5aTYTn60SUogi
hHsHgTgfYyWhbv+fHbQ23JoZO4JQgDeOlQuDEd+GyWChQIOdy5X0EV9rAhHkPxWo
PWuD21LaHUdxbphotVcn2k3UMWTiuUR2qCFLkrJ+OizcvOb3k2zi0lmUWACPpyHD
tKZODLsoqqe20O8medUTyMVVwR4XBLUKOYS6mrk88zWqyvXbQg+9ljRIgEoY4RwD
T6FPH/JRtELFEFA6fSUzw5xcnXPWLypzKFjl+s0l78/bI2KpvgLnt8EEHTkP4uz9
phQ0zegKt4ckaiJkq0l9Gd6hUs+e1Yb+HIrVb3GIuGUUDEFbCeek6jcMa/JmlgXf
GXYxFlo6GEKitqt0Y+Z047aKRlIHEdFxT4KROv6PnkEgorj0NrRdQwYKQesM92jz
hjuFk69MQK3f5h6aelfg4joGNduw5DnHApshKkvnClcKXHi2J+M6+hl+zwqP8LAy
GUM8KXMpgoN/uC6VAVNatTWH2ZafmcXB+YS7N8UzF5Juf85HFu6h/vp9gEhZAdLH
mZ/9tn45kyV2lFNuL2jg2TunHGw/lIJEV+v/6Vq+CP0dcYC3QLi6fKQGpReeLB6Q
zQVkZu8foCVhhhCdktweQ8s3t1OA2WVhwob2EBTpqwhj+1w5PupmRY4eufubTMTP
fRG6sDXjNlImtYWTY2Y0OcNJpyBLWOxd1ivit07jTRvYIkPVgfUHQ2/zU5iyr/ds
fl+VLqQFpSBNWX1pw2XeMtTrU4fbCKNW5aGnVX1Ti0VHjxF0wFr0jMYxIF3z/wHY
wI0aipM8TUogNEyWjo0nKskw2N59ZpYqQ90bgXy6HU8nkcYmZU+ycCs5+FgyDq2B
K4rFarw7zH1iPCCCDnRh/TFbZdrbGYotQFh/U+QzOLkxUTnmOFgEqq10fgEPpKE4
ZpZPnhFh9yXl+QPMaqlHdwK88ZfaPsl47TA6pBSTxZQaXXI1zEUsXAbbSn2Ef8/r
lpklvsH7tK+qoIqf7mfjulT3B+cvSlK6jpTdm3gEb5M/2JhL6p90hgG3FoH1qjPL
fdknhYj0g+aM1lQ9E+zBO8qZJdEKwGhkncGPZmSPbIrqv384UqPVA2eB57F127+8
zpp+00jn4VPQ+uZKfYg+IZhj6DKAV2MkN2U6Zu5zZZiW0O4Elq+EJFsfwKpx+Y6M
65RKXAUJtFIzj+sSqIeTk/azIL/DtBpzVaRTvIQcymAPoMqAm7xfURZaRiFGKs21
2SxxExn30UoElpRD+xinbwdd8a+XJ7HCvF9wVJQ1VCz6yN1qS9OdyawQ0M4A/MdC
5w0Iel/LqnGoUaOaBxflY+m4GjcvfWiLAwbE1mViVdgnmT4vW38VhNuMX7vsatYh
oidDAInL21ku+V+UQEi/EyNAjJmuiRxXRiJkyPn6UgKQsHSP8HnlUGUyMJpdqT7g
eCBnSAFXhLqfd6EeXf+oyU6Ss/yhb7P4Op8xt2rbEL3inF2jjLkjDbF7XKKz+ZYy
2kYHIP+5rIIZDiZ8GtlJeJYxnfCSxqyqyJ6dKX+Ab0B7eZGQIeRGyd2uyt6h6MFB
f4bGIOL9KSONR/eEI9vwRNv9CGqPtK9C32Vp9aLGOQAEqeBg5Dg70ntzflqDRypR
MfZgxwRcIQ0YSOa7s/vhYITdLcPgoYc4E0l7Wp1+xJoZZCp7Rd+tkGgp9V3HrkSt
CC3tGEIsP9dky4xCiTEzd94rakaAR1TE6a2qQ5hXC556hmSzvfudUy1ZahycBxBK
reMWQrhrxMCbo9WtqUKKxBoXYlglNlQl4IeglDe/OeQuobMmRntHqx4N8zlI8Uho
VaVHuGFiPbms8YS8JHTviqQr+uF05/UgdRIp8bzMaoFs+C2Xsjyh0vlhPUcFSR8V
wntiEcMyevJqY6sNSkCJjX91bys8zM2geLZaar9f1GQHhB/n/Oeq93nhl3mftImL
+LNSylTBqD3dmzWIVDrbSD7AYJNh4bpOAOLLu4meY0V9HpdEs5r+W6uA9tEXRiu5
GlSG2Ea9WgSbhFSepSSm71AfqtJiKpHWSZh1wco4KrsNZ3o1o44KJY/AGOC6zmXA
J+lg41xl5FfNWiAj0TpIBo682QcnXpTbefLpGjLwOrskmGNVkXgumX+ghtRHPhMu
41QwE2GeWP+aiSWKQZI55CiQSZrcN4ArtwbGc5Q3omZGtpBhqlkJj6SgKs6gEbD9
23bCDSZeodxbQu0rWA4Cq6HxQre4J4E8/2JXzXjntL995Zdd6rcdFetqNZv1VWRB
H4PJcx8AH/FseiF43Da8KhRlx4zfa7zYjgWHTxGnACayjhuFBg3+zHjdQy5E2jB4
GrupzboJ9kNzCHc9DlHotqPzlA3nk/0gLXlPQocDo/j02zFubJQu5pLNHdqzH7mR
kPV3tS47d2A/oO6Iz6e6r3E4bkA4b1fNTVQHKlmy45Wj2zCihbQfHek25xZHMQad
cDOwPOCc/Frn83BuA3Mk6er/rk7AplGipNqHGeYQNFnnPwWDYuF30hkglIyrWX5a
uCfN6CDG1451DnkGIzAVGDwp0RnSn30JP34/+ax7ptIk51nbkIwWfaElyQdQ8jtg
1biaMpdzx4c/taFaG2xUy+Z0XQKQ0d8DgTe6+O4JqTpdbVw/RTUOQWH9dKxBB7OE
+VjQXWEM0UmZ5nJfUXKQAphfGrq26OwEU4rh0J266rAovx2FT6cAD2ih613MdteL
e49vC4LD3jJwFflKesBaK+5bdz82MW1/rDO5Q26BlFNDLYvyyEYo8cebvvLSll36
UBK0JwBLVKNefzWPUQOpF8AXKV7yLaOgwPEmkGVvwC5ON8cVeyfpv2ezIAh9H/F2
YkVWOkbSDX3epzbnTmI3r0EI6c3hSaRKTTtLB5AdTj8GZX46KhBo9y0t8dx3FQT3
zcBchxgb1K+uCZMmyuCIs9GWPMYtF9FSCjhdZD/abqKYEWRcyOpOjylmHMVgyogV
LZ2tMkx2kllyr9YOQkU+PuyzWoEMEEGCAWv/RAVGynkcq7TmkVvzqw/KzEz/X6dh
xy6VSSsfvmvuBok8p2sSBkifYAUSx6SVfAqfBkym1/fQ4IldBXpqGot4lqgOU0bd
8KVmNIR9EGv5ea6NkixRHB0VKVBjSBWmV1x42xJr7hobgBB7kyHsan8J4AmyuUNS
KC0PU0wl7478WlCliBmnrBqPKe7gMdniztzy+Vlhh9lNPQSxG2Ldz4xb/DdNYvAI
6OXk2MvkR3ocNCTABrMwc9Bhgan3FjAveYORRggTjb9gVPImoCjIpUM3GXtpQw6D
j6xYxSSYSXV0ZyFn+AKipzZsH/dQKC98UOtyHko/MDTT2tMOMMOmR9cgr7bwIWP4
aIpjUpJIthhsKmkraElIqrpDxVEHFDQEbStbEEFF13wjrE7xwUG1/n0LmWlbmtvy
o5s3t7QZ/BqOsO1eo/Ro8bqYvTnf0KJdGszZLXfyxYeR/ChKZluNrc4VUpl4lDMA
8oh7AuX2MuTfMzDM5LryzumgJWMnqjTjq49thq0PNQofsL/0U7dgAFPZUjh1B9Rp
AbTxVnEPUqLZ6oA2nUICsujNeSDg1X0r8dpzvT0HRTCo+qwEu0b7npjislz2EpbN
Eq94VBtKLU6QWQQk9VqoBRBMxbPLXgsMs+gToyapKxVu3owDVcANZHT1t++0yxOu
JFkyLMiAfD6ET9w+CoKMo7nI9NijvCOT4JdEuCIhE1x47oOv/srs57A+T55ytoCB
LTtOQLSgwaYvp3yhTimTpEI2bAJt3B+TkcUC8NCJYerwikfnj6/15JPCFrZmO9FL
oxCA48o2pTml18x7HCrWT+dk571SXhxZdU0eVpH2Od1ZOqxgPaMMkABUymkRQslK
zvaTYimonwyE233sXM276J/Js01o81cY92JNFxwVX4KL0jsik2rntwd+hPiRxgWs
lW7ZmH0A8wrDff8gou26eepn4CtVwlS7GSxTT+XV/E8gFju4Dpz92uBOb80YyLre
d7mC5OwfyWSEf0qrtSVvewxpeEqQAfp3yiYTsC3fYINNN8qcU7QsGdPY8KDI1chJ
53ZdtnTQ9q7dvhbzMQHKhpkZDmwiDs3t54vXuTzhPwfxpyLPWjvlpl25NVSsF8As
uZ/UUCUZntouQjPBI9C63kkzqftRYxlAMSQnZF1lw4bo+ZbQAK5c4T8O7E9S1wom
JOMV3YBJzY8TwPv+VMRrbWKSk9m0KqTItj2rG3xSgSASduoGCHuBpstQBvZ+yie1
xkI1VMd/VRkLlVbcIxtMpB7WEz6iFoqzxWd+XqJdNFiGpVVG1BzD9bUD8+9CQN/o
`pragma protect end_protected
