// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:35:49 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Y8kcITo705uDZmRn3W11Wp3KHPdTS2ddQwABAsK3krVWLJ2ev+pBiqPTckvqN8wE
KCOCIkWcPyGr/ykbb1fi4fok0Gb2iDWS64XWDj5Yaab1sG0kek/x4kluw8ZbLCed
HJ74JVnRMvr9gt68mVQShvh8rlNf/JY610Qj4pA4LAA=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 3280)
ZaG361DBbXIJAdbsUhHeysn41W3oOAZBjX+Ceb9inYGptIW6bzEnINHuB2gZ8S0V
abIfgO82VSj8U/W2SfGHd/dtcWVW8PKSYW/yBZCXEZOXLrflII8L0P5VYsz34Vj0
Suz/wNo2mjojk7xGM8gbjrwmnCXE3ckwPo758BPEUbLISrF+q6m41UnHnY4k9hd0
122fRHI+QcGNhuVsQYn3ZVK2Ywt2/HtVmt6V2BIIhkO6iCYBvrUUCYerahfCuBQS
DtZHO0Y7XZ0U5EqurunijvYeS1p83z7HhPWFEG0TE/YYAi8gg2bfNc2kVWakTtKK
M7kDoAiG50VDL84YxBJIQBJYVG1IuOmGkPVBETRUn7+iz7sPzbm3lkDsT4LGDgD7
CY8fgJSWw9Ity6HgRPn32NG7J1i11j0eoAL+EQaHkRAsdhFF2jy9la+Q81itVIDF
P9Pj2ar3MN/ZIV8sVyrTRZ1/XFx3USvEObc2H0APK+Tct0hYnLTu1TgvrD25ZxJ8
KCQS7BOsrftLDhf2ET/8v3yqvbfj4U32LOUfz9bW1RsboqS6Zh5QOAM96Kg40IjN
QNfZ36m+wuW4LrFE+zbfsEJ4fSREiSJ9ENYNNqk44gk2gD42sA/7SfM5sWOmuuWe
5WowcOb4yFT6Rv+zXQxKXgcvZt0aQEy1Hj6c9jbem8G4qdiI8n1Te+dNIpdcbaw8
5niZH/U/THITm542csOVmjSCILe6GxkiNC5Vu5nMh3aQYaB2UhYPS8mStqgjCbFv
ROC30p0yeHeWC71kdwDa14b+cgrZBgkmkDgrLienDZ9H+6BJIxau9GTi/FjSRa+H
ZQilxKv58Xn0x06ION/VzTBdaenmz/dm59lpFq5uwNq4YbgF5OqVniTPrxn2Ze+N
rWgEMwQHqV2CKHgcDj/1JXRsRH3Xbm99UpgrqyhRrkTf9tmN7LYjAipcZut7bTyD
cL4poDq7479S15Br+qPCBNvSrznmQyPFHj90Ab8YxVV5H/C1woOFUltn5jM+UUZW
IR/DlF5QKnyXPirePO+p+2MJW9LVRjWKdOle/xw+VgqYNxzpsuffrIqjDUCQV+dx
yHT/23BpxyQjTddmvxHekOX1H5bbbhZJKehxpcs9euuNywPX1RjhDRk6vzCG0OZm
lFNTn9MamaY4l26NwiniIMwkX+A0gPgFj7myypxGHHZilyZsogglsPITNgxe5/4I
9ry8owvuAD/5t94NpiXERPTed55RJWyETABucHhOj+wtHcn2jfwpk+B5kTTBl5vP
rsTfCkqMOKisnrjeZRqcMkCsxmAHYtVyn/9DwFk/UMEUjxU4Tdh1MIFDtQKz9Rpp
lPtuGi/2JaQ3zTyaOCQCaydsF1mthJjjG3sNVMcfFxxGjqMNVPs/lDRZUMLfManf
XqUG1Qq1yUwuq2pBeZIEZM+K5T/+00DMe3syiKHc6o8VEHchH+xAkia1z+ZXswDh
V/uy7A3iT0+NEvlN6r5INp6DNnzMKLCmjKkebZC2VbVmZYczPDrY3NUkaDzHxNeU
f9bV76wgst0aCKpxQYc8JrqdGNP2TRgerlEVwAmOMP4vvXGXaHWuq60t58wibCZF
wCd5LSSuy2t8+D0n/okCY0QazBBJs2Ltvnvx8GsrUMdk4WINpMn6FK1eEChFvCW+
r3n6rR2LiRYKh0UNvOBg27/mrbhABQaJVfvjPeuCj13oCEyXUaksBuuGRriBEc03
DX7NWp4WSWJD/wWM4zLWVpM0x0H5moALX7eXpH3Wmua997eaAqTu2sDwc5clInYj
W2JlH6JjTVNAOnFDmvnLBHFccDiVD7p/jeQ9RZ+othoWlO3Bai6Lcgqr3OR1xa2y
p4oPmM2GzkIBaBqcHimp0fLd1jEo7/IFhDLNresBd3S0wP52ski77eHhbYz0eifp
J34CjisPuQGJQ/AtMKHYO/6YcbXxwlVrQiP/g85G9qD0QIVNMRLb0tfjKkt2uQmm
ZdGC5qbZjOW1SCzmfE9n7F84JAthVr4vcAzdzh0SZA2R/Q5n0uIWdfLU/f950Wx1
mZ4hyYjVA+y2IkGNnG4z9G/9txtqDPApFw6xdIOVFfWlHBaZ1jsd3W6sJoJLWa8v
zQtmFb2Cl/0eOzws8o6jK1vqWSq3+FsNmvE4ch9p7ftT75Ya7kiGsM59BbqoGHRg
TrVPGPk4u4GHp8dlFLCe8RQB77e1sIPIyhUdyU3LbfOKC/NwVMENaEiLAIraIy95
rplYw491KNZJTKGAS1o0hVhJRmiFvmnbHIKBaX5iQqkderSPaN/Ja5WXv6Tw01J9
eUQu5L15PavBDwoAcHEpBrjOIGOnmmqgT+CzQywog5JD//Li1216O8RJ8Ka8LzhV
DirnJnZWJvTGxOFtGF2vnWgDVj4C+TGhCvE6Kpaysj0z0KXp78mXpcPPAxs9fXJW
iaCMbG3T5mreg+kGT2tqcm7MFv6TYhJ3Po4BfsMEEywlBN1XBSiKMVvxE/sDv1Rv
xWjrWv8O7d4NHD7uS3LyYr3h+B2AkDxO3Qif+Dj0MddsFLuUpm7LEHLIBBP/etQH
WjUVX7QG4TozLV1ILQ7QUsnqskBvwCJnJEdIpAMYvXPpMtKqX2lxx/EdD9gFRkUK
GueYv6uF+CB4DysxCPSOGVC192596bfZt6r0Umq0EMH5inMZa8iZSfSVsxVxtkjU
KhLC5f4dMPaMfvbWkl93ARCYM5Z1Y0eZz5ZcrJ6T7eJaSQYJEeC3hklIW1Kcvygc
LvLezwwks+y0PCcRq+WM68+suYAiiSWysTZpiEdnS3DLTguFvkvBKMDeLhjvCHIf
JbkiW+DBRkS5CHC73GwpRJK+Jprlu8PEmmobCA2QH4EKSWK17RfWRhLC5+yJZzTd
bXXPJyxZg8PsiAxhLe6cokRmetAcuWoifzNZEUpcAyUsijmLaVZGdAVN/NrWGZ6X
PlNDrChRyVFswstsUGo0AJAKJRFoMLefhX3o6r+OhIRuAD94DNxdIrmXeAnLKYvb
s0uC3Ub/aan1J8wX8a1src7FgCewmeFDBL3aAk/MONo86W09SqibU6CSQvn83x2h
CR+dDlJhKUwQFm0k5qZaR5LBptuqjWdAJqqdHwMualnQJ7WvRqxu2cX+qFWyqKPa
z0OlOpcYe9HR0Bx2SZ8uwVnI8Xgm3PWpFRwKViB+WhyKzyq98fYSnZA/RKGPHaiK
rTtj6+0PujAw+qEkiuMIipIVK6Io5kQLN9t5G8ViSNGZSXLRQSOQY2/AUO+Fk+V9
jsa2o3gRhmIssB3k55oAmflJcqJz4vOvl0K3NBv4lBiBQCGqLilBgvF7B8xjiPs2
BvV/MxhH/zNEVBmnkmFq0FqOQpHW/H2HRaJPWdG/dHC7xE0rN7/oCV7A26uc98Xj
g96QFuhyf6SZYajuCbR2nRHjTxAfCmw+oMX2vynNJV1tSLlioLadbVXi9mKCNMUB
XXU6JSzo/o3QwGklOe7oWz8NPO7VrJRTJ5aIyE3VIoP8PkrTC7VrXthuoY2LHiWd
Zxha9dulCuHaZxZ78cynxpeYnj9Eb2dX43vnTPd4FqwdZg2og3TSoXthCbOlZsdw
22OPRp3fU5X2/YNZEwvij6OcFJNHe47VNlPhL9y2B+rQugjg4hmEw+btX9h4/0ao
BFqkmAb95UlEe4loqIZ+ULAHrUM1wPuBukdLh3dHT6dbtJAmh8jLekuqhvhzMqIv
Wsv0xX/EkymNcBuVspQj1WTATWkMOgdoDxfPccFDqtvCVWQjTvkwd21qmuQlwBTz
Tv5N9zk12kRJnULRXx2ykQtM8CjX4QrZKUpImAYJywMwaEeaYr0DgzReHxqnURQ4
O4fNMKPiyPFCLhaX6rKuipQjZVs5zr0nbHtVVL+uQk44O0D+1ZMOwzmKofGlccWm
ZiONZRkKsNOhQKe6y4HO+eN/wByK55tj4oZhKpjpT5y5kNrQMrCWIY4Nzh1OOF5u
7rAlFZ41MnWs5ozC0gzQThlqsBpjglnr3SMJtIB2Cs3ComLrD5iC+4cjPswVwOhs
vxhKo2sFjUkaFGfFLe9BkJFs1MhX1Vq1Zj7/HY69QHiSTzI8ocOHzmtLKyac4H79
ZjdJnkH83BLpWyC+cURfOgB8vWOI9VY+6cBKAS1OMab2UrMSY9bF0U96qyEJar4r
jN0VOJTOT7VgPwxzRpzaiSumGXwGK4zHo1+yw/NCmyYiLuk4b5K3RF32hOK6pArG
6HeK+0126yd+vcGJfpIx0BUJrnE1zmkm5PJgG/GvV2xsYYPxVOGQMvlfKAFe6ftg
+kr2HZKjA/PGohs8emwseYFDO2P6VHj8SfmQwAd5ikcToPUn2dnQ+b/2f/YIo9+L
gFHjyOHCF4truXXJm0HxXQ==
`pragma protect end_protected
