// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:39:16 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
UbVPNFlLlTTohBhQ6natykHFwXhuzg0G8pOkjlIy3f35OjzuEm9BhmGVlRgsHvhB
OWdDyNHEikXCyKHPjej38/3V6yXlFwuKbjkfrMIDYuuydNK3lt3t1b8NeDfF5Uq0
bK3zoVd7NFHxqCLkEpqM5UCCZ3YaZoSzZUJFobTqq10=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 17040)
ykmFqtvP/ISMiAoexwWR0D0RoZGRYyAjDqFBGZkL4k0TuQYjH6BfgDvzMo4zmLDh
U2a1MssG6ABYy7403h5MKdtYazFXE2S3Ex/+RpTsbhAXSatOk8SgOCRDInesJ21O
Bl0UFnOToHbZoQgES0UT/OdBnIeSwRlCM2nSGy9Tqkun52TrrlV96lK9NLTCVNE0
tBjTQg79btjKWC/dVh67RhcZAYC7loJamuiI8fq9gL2P3Mw8TyFNU6L2o7kclwl9
Wsks2e5ORwSL0ojzz8GPI945wBz/9YCyES7bvaPCe/Ys0z1FZly9PD6V+dJLjGmV
E/S3Z60VOWz+V1JkH9fnGV09d7tplH/veMvznzn+gFb3n6Y3bH3SCTjyDZ4o1sD5
Y8AsbCMacHMM2GCWFTFDebrcCTC54+PhFLrS3gQB+u06fB95WE/3z+OrzEA2UXeU
RTwzzRI8omdBfchhTzu+tAS+J9jeX7iMDz7RtpnCU7CEzfBa3gJzH1nJ4q/cmY1t
ZGVvMGphZEIzh/mAiv8uz0q8sLMIisDKNBsbYCRrf6n6LW2pDGWUDYif2YUi2gUJ
za/ouqCqad06QzfSZUkzrkvAqel4ERGsi0JEG2+xu3Dnlht0q5myfWaLGRyGtqan
3PaNUuRDV7tvMIum60nOHgTtsaJQZiTjl6wUqoDIc43/teQj7mPe9ZU0IOJNEtPQ
xob5NBVIZEAIBA3uvKBxSK6iOifJanBk2shbx6O38EI0DKULLx0Z1DLF9UJMKdAI
n+0ktflfr66cf0nUkfHxhQK+FLsjvuLoOd6ILyXx88JWYXnw6BuAqTXE8LGcuFay
Dd/WJUhQnxl6upNtr6QLQOvvi3BiiDHmLH0R7xckwig2/LTI5SzN6o8btOrFrlrp
f1Q4tJr0OSQFfDa8I0pMoLVe8+LJpy3ahXxT1cjxSTVhd+UfJjmQeQBr706CNcPr
QC6jMK1gnVcuMEhqYIdWfGq9e7zbxkzXPjzgpqxDgberONn1XUqCNjqeqxqWDR2t
Add0Zf1gcqQvNopwuLRp2sb/mBg0pKZ1236t3DAhSosstE5L5/b3Pq07nMw9Ttkq
Gxr6LGcT056pwU9qf5JqWJFY30NutEmT48yoxP/O/dAcOcAvKgkNCbE4se1Luo8M
jeI1MDb08k7FUuzP9AJAtfSiHIt6W2lDriT/bCeYYNVywHOvDh3cgWNJgB5imhhE
K5hbxLnhrwKHBc9lkTRuXRXIy1S/bICv+6frvjX4sBpcFeHHiEBAT7SBwtFkksIV
evHAYMfDqevg6q73+n3spZjaIAgEvnOSC0kdahTkLXORDuXWu9ezDjPFngseMoia
Pr2NfnDhg2Oy0QBlEEwojaLC74/jDt4q6XX9/frLbRCUsUFkIu1fL46zhUOXOTOr
sL9FwtAL9JF0fPNEPCFn5aNis2VJXAcmkW5aLO/1lyoSs4iUzT0Vaw6YxcnHwiLw
i9pRPweyyGyH658GWemxE3GCPbA7Z99aMkfk8skpVgNfa0e8cW4tor4pEbNeRald
eqEs+FrF+i1CrktSkfwClDPp0bdi8/xlxtHa64wvqbb1nD19JWhuR2wX4BnDG7cp
qe4NfXzJ5jeolmZ5U57osUgx4xNB2s+fWPOpb6L4BQdGxgWlPX5akOKKS4qsWQg/
rpzUipU171W9goQEgXIRsGJpf/xA5NqWR4tfuy24PogMZSMjensicP6POToeYGxK
BKrrz/gKK++qvOIEXp7rs2gfn31a/LWp/IFVrTgtUhZPXI4aF694n2qH6Jzd++0h
wm3pCAg3cX5ogWr8vxrg2MxtUrS4/uihSOaYyP8R60JIpZaw/IGl8xutl/eFipKL
ZuSBcuCw+u+rXcsbz6ZsYCia4lL8nFRRMT8zDK4RnCy5ysL/ReK2wL6VfYFc3CSH
MNRmgaWtgGvYlRACphRSlxBXuooX6uOjsCTTS2YBMlp4Dnt8tgIlB9zLr97GzkRR
S2kH73wJroWEqrgakC54qoekqNarMqxOAOFPUafdCUeZvRB2Q/H/DGNhZQKF40K+
c2KewZlvdKsn1oqQ0/428CAxYHU4Y1HxTcDzQQku/Ls+yKnF5gP4HoMbdqT/T3hP
wU/WpP/uNW/WFMTsu5bYBehOL2Rssh1zjX15zaukisRCbyLa6fYnjQYfqx6KcT62
FAd/WBe32tyzY5OZAwG1jzigTyw7BEbjvXhpwaOeicppbhx1CmrEZEFEXkif/Ayb
O/iVgw64AcTHHjilNBYSwrHqdC2eFKpJmKrYAF55CCodK/c6NERQY4wVS9+AMlPP
a24bGQVp9KDd6VHk0QX6EKtoYjQbHegYFOTR+PZ53JS6zpG9Mt489UpwQdmIadr4
gPQFHp73a16zXJuDzAkRyppty7tJDHQBvuA0+e36gGjyWJb5HOROFkgg2DZbGgh3
c8hYeXZ5d5XcBg3sjiZWDZYbVBOn+jvF0AuD+Gd6I1P7U5VGPxoTU8LX2B1RPRRJ
sF0MWnsh32Fuvsxtaxok4d17v0ekXLFvvwSyVckc941ZtHU7jWcdAJmS0YnCB6B0
WQMIP/L7nS82Bx0E+Hr6JLee70dCL74tX9AClLMicIppy4omQw1mwEfOhgfLKxZu
XJHjCcMWHw3Bs02ai1owXBjiCoxkoSW7c2QzNfzopRZnPzuj14n/t93tQvVF4evm
BQt8hVc23Nsq4ffeBLAUrmzfXAce5EXxXRMAOV2KJqjkfmgyx66KBNNr4gC59rFg
ErsbKS+eumUA/8EOoHxxpaXNLE9yvApVb2/6QdbTIjwZbbHxyMbo8XFmfFaRtWji
Cr3BRPVXlWsb5GnYSs5X6v4p+77nHRwz9DJhiE5gZfukdn/KFB5Kr/UJ1eAE3fHF
IDWGoqgVK9VmRHhlYAC0FWjQSsB5JwGIn84FHalUPaMiJ1Wwp24cImh0O814EFHp
83jFXgxCEuS2UUl1Fe4u3jQSNxdjHc4eS3JwkDTnjxkv5awmZyLB5Zk6GvY65BAY
gUUjCgN33awVIm23tXLNvIR+o/QVzTuedFZzN5ktuJ5Y4GKWRXMTsV6YXm8o1Wjj
Wlh34ovPzlQAbYe7F2872Iq9uIoFe6wcKsmhFVfe5gtsHHg3YMpsO/QgRvXbqW2p
poDKoSpAu6FlssqbN9wr6ERzkk6CM5kaGHW1CSp+yCqKWMxwVPit2+BwwwXngrFV
cbuPzAQTq7COPSk1IOvW1/isU2MuBL8olmN7j8rpimrWkM9zhxqSIoHlj8RjnCez
jntS//2qVu/upiAk9YUp9fRTPDoQmC/yktQg72a2iI0+hvYvvH3me/S5yPf3tFly
Zhtzo6DJ0sC2mAktrm+pd+Qg9H8SMe1/MgEl2Cu+aQQix07XZ9tielEo/yeLgMj2
8vNqvKFINCj1KrTGc64yeE5Fvbn4ygsg8VFS7nIZ0YVZdgZtm8lExDUn/kcUg5wA
X9E5sSiiUaySpiJZbVDk5b2ph59JW8taHbyOo1V0k86uf+v7y326gcPRmZQSUEgd
53e4OH3TEKqb82D4vGRDEFnF6EQSBelYJ3jFvs9oOEotswgkZDUD9CpPD+Q8gk5S
TXOIwXAR71yogsy2VkrJ6gEx+ngf4Ac9Gtmax7Z+sR46zNR0WS++mpxd1X3VrGnD
NcrbVgw3Z2EWb50LdIfkMBo8Nn3UBVj5s90kb36EIPVIE6qI91BtsIbAFgRLGqk2
ms8C4smi39ROTQ0YVGKd9KIH4qLJ7KdDLNWncC9QRSwcuswpZ/IELZTqfZNu6F92
Vpe9K5WttMw8AHcgZqzx0G4k/xKjBbasjRHLl/pcickABMynccLuIPn8C+AlQGTp
p4+qJFhgjIdODbwsqOthWjIHUzVhJrZpV0FRss94//c6hsebK4B09VWkvHhBaxxy
oJcm5EXSIAaZLY+fRjFxnxwN1BbgRKD1+WKBp9e5tZPzok4PtV5re5ckXSuVoHq9
QsTstTn8n0Z3EmmiRZSnb6r00c/Hx4RIBty6CaJwm7AX+B97+FeWGeezcIBx08yf
f3U4pD4Z975D14SF/SQAKA4DE38PJ2q3AoQdCT8EuSIbru+VHTkFvKM+SW1J0P7E
dI9AqxfENd+cMmwmuivBONds6o5cycs6KdFuQG/0ePfjfuvRskDkd1f8fsGy2MDt
NQCFpbU7Iyb2DYdmUAsDqep+Y2iIWafeRgIvol+mqJsQ6iF92LkNlQzKpo1Puw5/
5DbKjfzi4CY+W8+Jtjgc4KIE0rERVOEFbGKPDHJvHGeAWjj002WYewi3NKHicFKt
mP+CjIA4/wHcyqZSYZZjI8LCOY1A0bG/zVx6cM1SFhIvssjgE4B0RiblH+CN7fXl
0XRdWLk000nkOAAIzH6QmU6J/boFzxiQzuE7m66Z3VxkDvxzuHWAgmmAuX81xJgk
2bYi8KvQetB6DrgJZiEdr//lM441o9hNPYn00iLol+eK7Gf4Izv2w8mxJi8x/SmL
wZatD8UWOHFianUqbZdO7FQEpMnCeaxtYHR0fsvV8yCONOaU7VNk1iXS3WWnt9Aa
CVKnGLaSEOgC+ORXoBTR4GIbpxdFRto/HvAwddvojRz1LegrNhWutHhtP8Tx/2wJ
dBPoRGd2gyaIBq7QrH610Tx98jPONTnWfjwTzVHboZxU2ONDway+Hgx/8PJLcWGk
iVhVli27dw3aOSL0lhPE8FdFQ66iqzT3kzssjyVVP3Wca+KCljLbmF/Blrn1v1aS
1u9aR656Q3yQoY3DtYUv2zi/HJH8R0fW46LOGUvyOxL1svqtY9ZVZXo2DNT9KfgD
t5gLMDNcjzIBDF/vvmrIhHpntC3yHrHapSb+P5eABGFpKdxMikGP3KV08ymDbIwZ
znOSFN96VFISf+KEz90It0/0fyrlnVXASUEwKEwRekZClMH24orCy6ouuTno9/74
tBoT+S0vrZx7/CiGjCoeC3PeWfwO0QXQjLHjOTXq6N+WC1LriSBMiJVwsXwG1rYl
wif7kU8it9Ga8ExeCxlqB128cHmdT3M3Dh4+En8hW5zjbFvnvrQ2S5akzWBshYII
IOT8OgH6SZTRYwiy1Xd+DontPAI/7RLsa8Q3Ha9Xj9SulZjJocuHhUDW3iedIKnf
eBtS/6752osS0+hxj1lk7d2gKov20dHkUArQuffgaYrCzd9CL/HicZGS1PTwvRvt
09ZyQAnoPZXLNGUnna1wSPiMZWV/93p/8LNM1LZbApT5UqVFscmP+1M3Pd+M/5eN
Pk/1XnwVWIN8CwuJ5bMv4/zX4lKjzQUkuWSiki9kUPOkLzmn/wqK4ocsHMyo4nuv
CTVHGldtZY0s3SeV3xoQNnL+pG/EpK9HcYxLsKHICBBYwx3MnAjS+6wR7isKesUf
F0ValaLyDxVMOQuLVVReCpMUp7G5Lt3DkvU2ip+zmQBjq+eZB3dC/mGlFIuxScpq
zz0x1H3WU+lQrUMyw4cEC6dGCKEAxmc60OFHJn2HCalrL0zqyCqtbBx9TwDcDLaG
c96ZwxiINbMWjx3dSA1U87/1hOANHg/WV5rGZ0cO3pDz1U1q0cuztULlsu6cc3Bi
GADeX+5oNVZKT1y9Xm/oPhWYUTDgo3uMOoE2RbuwxgIw+duUTytb6pex04IXveXL
g9LSl3aZTJxEkxDgr96w/PsVBuJfebgOUtel1yIoIZH9ssCz41TdoSE/McFhaLc8
9sdkPd0XT0l2df+gBa3NLD8JBVwfkEjR4SBe8y0/j4G5GMO7eefRbAuI5XzaLtBe
PjAsLw6pjBjzQ9afQQrU6KUmUU15xr71TDBPaCIfj7BLm5XeKOzLF1opKcvcCN8v
87XptbAOM3MuCL9/bA0zMyKcRbNcPeR9hQW0W1WVyU5xROXAAVsrgSdJbShXfI9o
BjxgGBoIZBbNUFZ+3UsTqqg+XluaCYflGjX5nHigl6vfo9Tap/Bi9vxx8/x71sDu
hCOQacnksvkWSXH9gth3DcIHOi3nlaEouTSDcabbkbpX/2QkmLxgpKwsSfuCfZgF
GQ0SV7+PrbQaYEtkJYvH5kNcJq7BAe8uycVFxc7hY11B5UEZxxE613gkwKytZ8L+
TgeWi+7VuoXc3fQhG9ZJjZqOL3bUjM6R6U+fpxsiLhIRqB5UwERuOt4YYHibW4AV
GYanDKzZUWYg/PnDFHC61CUBSOR0u3cxq081mLK0STuwDAoUiE/L0kipEo62hqCn
hYtcrheHBwXEhRf3ipgMQlAWiuW6B3SNRMulENQgsj76jEmvHwKQ96/dya0Gkp/J
wL1lL8QPtYcVZlos2kzulZLJTRj0eBXctyTk9U7pm7PNk0yuy9j3F0Oaf5/G5Yl/
z5pIGrwVgQf5MG64qpGs/T2OnHYHsQX5cQJH2tYpPdZRaUZumneBUArWclMv+VOB
wreccAlneSzg5smC9Zxb+I+xDqIG4bw/2enRVbMtqcEuxPvY1TLy10PCY3KFhI24
H1uqT+jl2BLJinuWpm7d7cw0J1sh5ReZvsjDhDnTnhsOYwsZLRcu0nbRJFY0ZERW
rVJzQEIJp2E5+E6Oj8yodrSCpPpjdCWhbLHCzHEGfI6Qzs3ng9wL3QuvuqkeieUv
98aI/vJs7dN3ol/q1kvFq0ixTDsJ0nxjtwz0dlMtrEQhysPTM3u3nwLxc1M7muee
Cf3djfqdLVLcj24HNus82op+FvUP82ub3QClsjV5nz1GUGFjeeWVTa2GiOHyEW/E
OfGXyOA2N3h3E6lS7aCtWP6AIu0eWB2T2z1xRgZn7fLuKXxG4+hbCaYfoNdfUPQo
6fNKGBC+QaLeeKy2ZRo6F0t9AFlHNNk0LxDzTN75w+m76Y4//u1c6dQvK9rOT3AB
JYbSVNEQzMm+wjoC2K7G3jvgGbe8pN3HhsMCv1REnuft4PzZlWC5sBCR6KJoFj6e
qfTNJHTE8Ugex/S7G6bo6AL9BTJ26l5BqDmbe5Ub31vBpa1c1etTGC7Vq0KPWK2s
02YUEzIW3rgLNHd+F7QdGI7AP8ZZ0EDx6bMleecQSbgN15HvK6Daiqc1w3CzLesK
xnH4t/Uhgnfb/IZPkWAVj5cxmzugI2EHGbn0wmlwho//kfcPN3R41BELWdPKRjB2
rglAfqtqoCfBHyQqtZxQNoaHkRO8iSzmWSeQzYzhtdQMBmhpLwICmXuHSmd5j178
PX5AcXc79LOE4RDyzeIeZWFUsErEpZ9X3JkjegfBbCIdmYSAzqI2u64BtiDf9Hys
9kT95RJK8QLagsj4wnfvyb1cA5enSb2yBB1fElDX1HyIkTF0txSrq6cp0FYJaIgB
+rDdDdeWOu4uuw7sqNDJ58mnWL2uM5sUNsaz90WQt9hbGalZoTLN8vFwKjpFDNDF
Qc/VHBf8sDto3/Z8Hh8sVNOqwDgNOGqnCZazKPApV4EiJ9t2hIDM+mjAkLG6zAUU
RW1WM5wncbYZeMynaRXkGXzMqg2zt08IZBptzBOTnR5cXq9iX99dycdRXrjt6V8Y
3HhmtbnfgsQ43uyDUtKt2H2RzpYxaI+bRTSVVwXMyKIiD/NkDNu2vlZIV1+xWTOR
W56R5E6oQKw/7iewXSaUuAZgEgjfGVG4R+XfNRK9FgFP0ACOeRgpPC42/yQXHNFY
36KNizygS7elD3w7Qpz33gxA2VHPq5/R3pEYVY7TMRQpbcQMl4YDS9v/9iPrfB9j
R7tQ1qmqKUIyIxPHjmH/BAJvKTEPatAxiiBmwYmO4Z9sVK5xhS3o3Lv6bznLLJeQ
oTiiUY+ufJIHafZQimvt4K4nHkUQ0FUz4EZBUbrLw0OPB/DmtqYCXf+GdIBVNvfC
fu9tClZBKZto2nkyYNuY7JXdBlhzcMHDPXe9sJRishJoT20cnLFvM6BdyQaBVxHh
zXByvvNfzrvcVAUjPufAzGKJRm6a1c2scUsn9MqvGL2bhnlMm0KIAlwrDv7kiwSi
Nh13g1b0KLatDoIeywcnQ3y7x4DXMkJI/jbbY4LkL8SSqdNZ2QEGRm1XlxrdoQkp
tTn/frB1c4iCapOU2/LB3khDUWxuXHjVGV1gniQ1uAujwp8mpLWj0tO9UkUUMIT8
zpDfL3uDYxgDFkODEPe+p6J9iBflnS5ogX9QMyed1ubH5r1+EHP1Pi+NVT/AbPKD
KYOAkOb06IduOJDkOlrB0RRh5bfgDVEXeLgFSHo610q4Ub9GkA2dbxHfFJi2kFWh
xrtA/ELGe8NjnBUieQ5Y7L82pOZeQo193JtfePhNHkS1m9D7a+vdd8Qo5dcq2Kyv
YNPntf724AMLQPULwgFdM+uUFJrDiPO/boGkOMiDVjPXZ03gWXV4gWQ+7C1CAFvf
4sFEO570WtecOCjKVOokMYLxBhDJkXS5Ph9LoeKEUqCIEFdhq7W/FS+EeYFPemAR
KX1adrWG0es27bTx76unDGQ6l5JMrmDn2Zze4Ahl6orNI7yIJJT21Vta0Fhg6Hiy
HgiKI3XKHwXoR6YujfeZ2DrYgraNlhZPbaGj9/msb9RqH9GCEb2KbwMLehuGiPR2
16ZM8IZLdkhbNGUe5W4aa/Z0CL5yCUXGx83/skOS+fKbcdpJA6XrXOo+1kbmxY+q
WVjP1uYo3CjyiuuwVjdIWdhK36elMXT1PmW0IpBUa6hkQ04r9YzBnv9ux5XNebmM
btY5PfCmBW1kagET+DwngNJJ/tIeYhRbB1JbGysfO71b/ZPfgREgo7NgHSM814Wh
FvASYN9MKBxSqIosAxZqZdFpnZqZdOR7gRni1U+QXnwiDoM09doxsIsMqowXua1a
iyGqh2svL66QFTv3mJ9HY65Uy7TgB0OfqOpCrA3jkaIPPnYKwgSs0IE5ODdah6ma
OJAM23AYSUrY+TNi5bamGKRu5QLAZTOAiYIfRIK0BRgEvwjNyOAWvAbp5VNnsYtU
fTfNILKOVBsA75mPkRopG/IK2xA4djs6s1/qKbY4I2KuhHMVpl9WgENHDklMQdS4
oZ5k2gx1s8voUaCZujs86uJ0R/HbcFOSEs+EvuwJTb0d3lAPag5K2uVsI5w/C4z9
cfRwCOc6+Xh1rJ25Ckz4EMZgFtj6JjBpXLXzDuT4zB7No08Nx13Btiy8PhcukbGm
aW5JfyFqLv/IfoTAL0zDZSsJ5g4YRtwqKfU7KwYZzhsnvgOSv4iIW6mT095oYxVM
JEC1P3nPY8FPDh9d5LD0fvRr+nLXlRra+d83bKT0AZ7BGTSHnN3fGKkX+mJXVeuz
+gcOx2uTo8JlJOcuJvTyTfgUbP3wXQqIcDybGr7FACQ0H6eARURwGI2WdhZlo06X
TEorN+QoLqzozh/6DrKKMR+NpitS/h58cRN++XvJvXG0M1DWxgXPKdhSUeKhXM/j
F4+Z7xN0sqEcelc3kzeOW4/ipIdD1tnDFJq65UxDoVD4LOLnQSMpN7RSs5jyg9Ck
8eFNG4Y31Tn6A9lYalUn/STkzuns3JtmQoKEtu2hj+iX4zHoZVZlZNoHmfbIGglp
UutLnAc7MGJkcXDYE3ESEN62GwkvOm2od6FiB6HdeuUd1A4TaxuO2qMZAo+jEY2o
Lbe+Ba5Xt1PNtqsfN5l4Ebl5BXtO1PIo0akUjE3RkYxUlp6gtezSEnlPwcw6upfR
TIrPVpc2CBGFzLhpPQxjsVGNi2GNFvo/Ygra8952MgpSfAUdt88iyGRFl7zX41sq
yg/tsIiy5nmYfxgs3118MnHF+GwLgDsHlhxJJIoQzoDHrW+f8hbu3njgR19H1RN4
BrP/vqHuj8/Y3LD4L4SCcOh1V+SgLnRLcJcczJN58FsZDVV0S8Th7wO61xnMEbgI
pZrVoB4cABy8ufJvju7pe+NRSFZurcb0a8QCNwQ7PVtslvu3vwMngxlqBKW5bdDW
hA80SaQScMYD121uw1Bb2IgPUxWIkaRj01JpT56xpo8AvEsL1nL9bfGiOcOIQqhn
0L3WDS2dhLF2Xl+zrTglXexObd7A1Qzp/xNacT77E76ttTwZy535gpfcJNgTt4la
J+hhF51BZ4ltAV/QkihVwLPJ/0wjnYeRfh4jI0tm6YwbFeLnZkwhr6xiuXWGSYKu
ogXr8JQ47Uv+PXtatX0351H3WPpm/iwa7XoQjq9mym8Pr/s+2e/HiSiNAAD1kSLI
JLlM1IUJIfqEj/0j1WThlYfH2H5SsyzyG2JguUcw8WFO72LOe2yVI6ZVMOdgmWlX
PSdFHuXKUACSJGoTg1tDuzS926x8SlPTeNb974mZHtFWFmhAbv1JyNm4kDb3dvA6
x/gJorNwbkAzwkmFZOIkByGzaa3vGA+1cceEl0qaFi7iu2PfCVscvqtwb3nLXit8
cmAxjbCi36ZkVwfigdOs/e2Qu5t8HQ4MCT9hYVUVsQxxHhbbZ1L9zmk+3OVnnPTx
xb/rUJWfWwG4wxobI7zUXpglAYpGsf26R2KqzmMy+8a7AGl6yq/hpThYWha9IYfC
j+To19MjTtKWc6+AeBui5gy0kOtu+MTzf8UdlERWFxkgooZgN2m2XBleJgIbyBDP
i6nY6yxQj9fFv1hQZx63KJbSunGqwHpD0LEcTPTmo9ACo60Gh7AHlxyWo/eSZlSZ
WMPl5GyNSCt2g1I6Tz5zduvo+DAUSl1aOFIcjqPAZJvNmOO52G7nbnZTmTbZm0RE
2OjvfNhmW30NDJe+UW1pMXGeo3jYc8akbCNdRvO5z9T9u+FUPu2lbO9mwIAjbEVE
90WjLtRsPMxSOfxA/g9ZsBav/dja0kjnisLowF18WKgdS4BJ/F8UP9qkKldDyRWl
fJ61j7bFcLI40373FpjylSG4GMY9uIZ48Y+xlWsKUnZLrg8vQUXLGpOKI5ROKg0U
VE9PhmZN44g0hGTaapickTRwJxKXGL+DnFXWiQVI1XT+xNB3iYRURr3B3EveYsPl
HZSiNZm4/RikI/FFS31loT5KKF0xdPGftsmjXs1pCZk3TDdc/Z716tHmw2UP/ClG
nY8QCQ5EiL17T+nHzgkgo8vxfdH6KcVv/GF6BjZ0Oj7dJeXxHy76NmHLPEbxMUuc
9VK3x2IomnT+FScd3M39w+FZVlGmd3vKmd8xIl+YQyv63VgIARxS+/oyWXlFlmed
DYa5QlBPDPIm7BdHSifU2dsx57sxZesvJJV5dtLYM6W16+Amrj0hwzBuvH7tpi9Z
sSkMCX37xpIl4UyWHgW9vZbBIuS1AXDjB8b/26vqEE98lrBRp+pqD0s0zO7fuSj8
YUndvCNyw1uevHV9cGuu1wLcQyHBb1sWYh6J/Jz9M4B7kOxZZw/gHkRoiJp1utlM
Qf+AOgzihC5FDmfantlJtZ0cdmlPHN3wACToNLXs5K9SdM1Gc0LUwiyqyYIkeh5j
R7nspyGzajYZd1VGYNakaU3ppPILDuKfyXmCYAdcZD5XTcuz8YOiAm4Lk6c9tWH2
YLBqNniAiAcT4OGJxcXMpyBOz4XuEZSndCieNjNaamSVHPyc731GKnutBv5DUYJQ
vqoJoR34JP/JnXFL1paHJlCPTbsXvA7k/MKHjx0y2UY/+d0Dve40DTq41iUBJlD0
Gc8DTvqZw3fyMmYd4fIgwRCSDZ1eD13vLU9HjVLHqWTpxfE+kgxJ7oQ+JXhomBjV
3xxlJzijewbHKHrhkQgi+FMu+R8yupelmdVhYsQOiojKB01JeCOfC/4O8LUuwTPm
lKrwqYyRoE90mwI2JH8cMrkKDBRMUPh8JVYJvhQJb//jab8SAva7VNVP2xB4eTqS
+9HyHzKxrbmuTqcV0uVCi2gj8SI5VQ7zz9qiiMWwl4VV5du8+/Frtr5vwf72DeI5
xRCbDrY8P5T8fMRJRiGlTbWod5aw1SSG/KtjN9dMYrH8w95VSclzgOXASf8Qmsq4
Nza4q5ET3ZsYbGyY8O0nko8Os3DapDTevizqsGLRO1O1WEQuwurgthHCnagB6o/y
Za7XuuY5xz1RKLqo+y2QChw2MVfCxKuYNPpikokC2U9vKPxkvLy8OiDc0rhYrUsL
VlesWj4CqdwwV/dPSWe1wIkmC3kdpKGxmCkhMxljzf2E6qyXvvJinPnVkWX7TbOH
50tMjpQQKSyiRlfmFLMvLiETUiU+DOyQm0VF6SiDnG7ookLrx/h6VZGGVZ8vLBQI
xwfGwY932hVB3JSvyeovr8gM6i+5Y2SGc2b/YGLEhxj8OnM9Pu4lC6o5hg/e8Isy
qescWbyTaQKG+hOaHbVtZVUJdib4GFLlFOAua8JJLv230HbzDv5XDEkjMFh/UL1Y
Mvm8EP0qjA3Ujt4Rb6zMkatJytfmgAZCe9zrR8lIvWkjQYz4gE4Z8fBj4Wx0hNFV
9RBYlpZOOz2EDS/HchJ7YLb2IH/ukwULgSM9pICAUJO2nEijiaEC4wy9+hMzABuZ
KpUFZvNyT/RLF/25cRVLGk32/Ryazm1pHUsoZN6z1cNZVDVRp2IkHf/ooVjgNkfN
w0Pynm4SgcIB9CTTyS3V3y2dP0rPMQwVwLI20JUiXvv//P4OD/ett88Uv6V8v+Ey
BSbAdXZBRcm+4QrRD9ttCQSejyNGrRK6QJBaUWRaQ3hpHW4LyI5VedHYLP2qnEBm
PPWtOSkPkDccs8baEdjt0PArMnwMNu93vlLDIiRDyWNCtE4p2i7IAYB6WVPFzqxJ
lXHjOQ6rMrbgEGVrOzT7EDyqbzF/ZaDOWY1h6PFM3XO8ROgo88LrB9TOopttobmo
Tw8iZff2tCHBOBTicmtv7LIMX0AXUolqy1qnRWP3TTmJd+jFoSsnJO7LFvr5SIw+
a595k7jM2jDFFK5rF8h5wQJxFZqpQyHZHAzP7PD4PgAlg+GKxTDef9C/vt0AlDCs
3oooPMfldUnyIPcwyqo6RBQWeGb09lYhvEhfxSSts9liKKtiOY4wGFRwtM4OIAUW
Yrw/hKQLLQej7E5QpFR6rJG/YaSB308OxhKvxwtIlIOREICwtQ5CZAMWtgCquwY/
7kGR0Ktj618trMgNPj9Je3ydQw8bCBN0bY1l/7D8oN3Hb+e2AOvOkjpuVv6ihDfw
AyeESBA87+PWdsC8+i3RnQPjV+Lr7fycRJMQ5ZoTlViOw6AKgB68xNQCLPbhveNL
8YcwGXmg7r5kwHihwz6weB2TGIbNZd4Oen9BiRN0Ik55oVuNtVl1mkT/EO20o3bs
a8o8MonU+6+SF+KCjiXsMCmlSViw+KL3BqxjitqTV5vrGnL8QTQXHU8uHy0ytLbq
vS8iNjH1A389LZSwgVYIEzpp1aHIl2d/jN+HbXyzd0imqTf6T7mMqxaPB5zPpfze
Ct2l7RLvVGYgUT1FJHsQMPRp2w6NAbX+eG2AdEKJtGp9NVdbrDIxcS3dOZr3614N
6qiqf7rab9Y0qCCrLOtY2loNJy/HhStbWJgqFPojolqpDizc1zFbG+9vPUymTRMg
ITzk3Qe5rkxEGOuXCMwJlvkqbUyFpTpSmVKyM38Fg89V8h9+m1GgYZeTny4Zl2FE
6U5ICP2JiHDKPkEQ/i0NRc6SGPNbQM9mvQRGIyZ6ZY23SKoBs9l2+9fZfuHa4LGs
Y1DYFP2sCJF91rpIVUrhAqBm5pKOKL9vihDTYBKnC9q6NtrEu0fjr6BLD6z+F6Ni
EUypzERM4T5VNtPfZnT9yg79ayJgN42oD4Ble13HSjh/JZ80QWrvrDeBifAqHfg4
awp9m/Gcrp+uoznxoReWkimMWXxHhIT3VyV4eit4QuW8s+V9C0NLitkt1QciC2Ut
z3JtMuFBvwUyh/hn3jCTt4B8QcRyZQu7QpyBl9Y442Izg5Ms/F9GPuz7G6XE0Zax
b2kJ64sHxUfebmWHY05Sopn1Tb8Z75/dO0fdAsjipa6WUp8SzSJYlgifnH0nx3Gg
QW8TsfVaE4oHA6U5jnJeAQiH9D4y7PZqJvc4aSdUn5bUbBydgi8fTkTHtuZwKxNu
Vht6jBNrWWtyIwTiKg+OR2xfXd6LHqIR1H/Fe1Ak1CnfOKTr8nlxHm7euCJClgVm
f8aa7A4EYBHxgaYBcp+DY/x5zLsXHrJHjvHnuCKgfv7EK6BXlw97WWFJDiT+2FNU
JzWZe97IoGVWNacpnR9xc22wh8XJUCqJz0bQKojJaB1g0OJS+ZB0+uVK57uF3wck
Pg6ISjkKikLUtVVdOUzu2x2YFU07MN9rh5iskuncW0c4cRcgFFjAKhXtCBRpnSJb
CTXWZUxo0K+/zoWhd2hldYJEgW+28Aabam8jXt6mnc763e81WfQbtWuRhUWDVqPo
xjlMLznb8kb614qTITuaoRclKds6sP4/RNb81QeGGck4gm1NuXHaELRfjjI+55uN
EBMuc9wuTfrTrmXv25i3wqRTf7kI8CmYVACcYbkdcISX2qz2qV4pIgcyuX3EFz5p
YrMr05+gxSPb4gMf9nYlA2wwItbdS9Yq3p/WpGwV5s5n62g+6umKCJNXCYSRjuGr
8msWf/BWliXz+jkblJH3Ttbeued5iFycqV3/ZxCy0RiVK4ER2HUeDBfQFHrYaejL
AIzhU2H29VODoiZLWlRZpDsi2cyIXLuMjqzAhRJiX689AHHELGe9MhpPFQfrgxlm
sCk+aqL2IQBxP/QQizzbmEjopTkToPJbZ9aCLaipLt9rbdprX9UCCv2JBrJ4Y2G6
5TOqRXHtp8NSxbrl85dXCN13KMkVhUbz0Mr6MNCgMbWbCire+99ljqB7nPypj9DU
RfoJdvKkVXfi569jL0vpDABaaEqEC5AKcwVjffgnIlACDeDeLc1ZxFo1MbQjukst
JePXCvpP/ui68u/eMVpkbNu9cjyAYZmcvBxd7zafxsXd7k7338dsRFq4+m/lzGLX
1e70886r9Z7CGfY4xBlXdivUW1N2RosSDU/fj36oJAOXvA4kR5hJTCJ9505BUw1H
m3h4tsANp/ZNATGt+MJBfi9wBNsqPB+JxJkJoYafY+zjKbywb7R/K5FZ4+1aJZux
FRbnbrVpYT8EEutkKQPAXrhjZzLiOcR9VuMQQOWhgGTzwZ7tbbpH5ym5mkpfDRzd
+AfN8UEfn/bvUPyHCSfNsI4elM+i0sQD+NZVnsN39lE8tkcYI6FjFoAXCiM8yApi
IXfKtgUeeaVN0H47+qu/wbSKZLPAWSlXgPbfthLHTM3tkahZbOOla2WCed0ruzze
LqzDyAW7ddoen7uQQ5Vb8klSP/vfkEfonvy//twy9eFwLV1KePfFuEJyS13yVbZA
/Jr5y8Y39BXzGfE4IYo7J6Gl/vkfYqBvKRDKYMrkP2hihzR8mHMhFY/58xTum98B
ZqH4HNaDtcP2CUMwUPe4FxWrWph8inGGyQ1uGqyY8yv3Z3KaKToSwiUkwjuuo6nE
XEYu1szG2A8li4WKArFMoie/IIx2J0aAfFZX95V+rIhw9dXZF7ij/36rYUfAkb3/
UNN4qvI/koVRJ7kFezPWsSacbimXPeRbl5xxGTzpP2J6tIKTxWzVV7QP0OMLyqDF
qQwJEC3Sf6LhV0dYg49TJ822HknM/jNQHyz1djVVaUOotiHDcPWpzVhLPjkRYuM8
clu0joH30xZDFMH8eb46WrSIoNutp8hKDfeNm5IqS23tFh3SKfPCGsLejm8FlHNu
EKNTc4s5thBmxK0V/eDNtHpguPyqnkTrD9MLRGlOxthFMwBjP93ilAR/pY3XY5Jl
pLSspu0zxsJGe9XrvHqB0iy4JnD9zmNftiLjbZQmfqK2kVuhYol8AuBAP4EasM80
vH7KzmzEvQwWUwmlv0sQZcjlqHTWk3g+RooRYZQagDoLuPyjDOiE3RFUqdN8r0rK
pFdlo/FkZaemnGHpBQ1BwnMnZF4oGbnlktQS08DokjyUjwgczuJb/CYb1/6r+Cpv
6iO59qAC1Apm2qMbzL3QOJiWRx2DpBAIGgJ5/HSMWlw9iYeTJ90Fh/Vo0SoaQixG
QtHsWXPaYwQoQSgIcGTzp9cW7Jlc68UPdYeDDeKaH52pOTPeelj2RHU6BjF5Sqr8
85Cvvjo/XaTWqCdNGd/BzXLNm7yuWaRi+4nnbQ4xSLAnEd6bcpCeGdePUzH+4Shp
LlzhJ6NS+lb1RLvuXia/7BiA+Yms6eeAPVoA4CtgfxBO/1Cxt2khKTcEW9Xxd1ej
HYkXvYz3ayXs/L7MIAn5mM/Cx/Z/jXRnrHwHdSllA5sutOtr/cJ9vwOeATv9jkDD
gxuatZIufP+GHvc+cZLkAJt+tiS2Y9vP8IC2k7auFUcqZvgzSpa2NTCkJMPjhGvU
9XAwqvITuIHbWbMLyDW+PUtnVxhq6D6gogzSivUXx746ljtEbAbl2h4mCrhvvBas
Oiem0OlO8M2PoKvrjWGqLrTsNSZzqRxiIBBuV5IsWHkoIKE8UniNV3qDWfGbLiKu
EcHSwUCkEb+SnoTHTnN8yNO9qq9JiQ3xY2jIRnPKDuf2J9ybbhCOG4u2OZvEBZcY
dRO4VmDKL/BJRYr29AVzHpliAz5roldF8Uqu7o3Zfco26xR4WH7ZI+3MRI5e/I2g
WdXpOalCYw9ECTf/OJ5uFqG1vIA8JA/2au+9CqgbCaUYB6TD0/ARHSZ0sYS+/0PR
bx0GPswLxOQEqqxJ5e+Id2xYoKUtUdpNHAVQT5DeeU1E47trqd9m4x6oqzmhuWVT
j7C6n29lLGBypBjasqyVsDIV07nyeijcvFt9Xm4WPcS1cy9MxoIuu00Js2lt9lcD
2X18xWQvcZDm4RuOX18FEQUkjsqVm9/shsYMu/qylBqhqETbuASlUoZ3hrtqvryG
6XiZ77smTsCDbrUYDOWtdiIOul0zNt459gFipoP5SV1LNiUO0/7EKG5Nh7dLU3gy
SXkWXSHtt4FnOVK6XW5iqUT6H4wG+m9PkIzJTGCQom4Ae2/FI0pBCc46gELtFyZx
PAtYKhMEqXejH25e0Xvj4IZafpElpkAph21hko/1pXSsjZiz2BTuRhEFYl30le+f
eZMh79XJpUa6epzmT8IdeV9V7UD1htevDoi7Dd8NunOghDPnF/Yt4F9pmsVV7y9v
bFqDBzSkNA5WsJFdTWh/xqKTogPgJHyXp3/x5SNhMGa5tDRKFw8/yfL/QO9YkaJ8
/RXppaShsBJeDSdM0Y14/4L9zC3IF0tIygknaSAsGgIYO/tq0PGP9iMAmjmYAwI7
wA2X1/NLXm44hqrDSi4+qRYhP26UxVUAAqTNcnqBx8djD8JADGgBPamQ0mXNOgi+
jYBFs5473pujjqrxtGxzl6M3P2EC2GGK5T5QDqoxT0NDrrFPL9MyDFIEejfTrYwr
TS2dRWQdQ521ooXf9bCTvkHKLCpjS7Kyusa3TtimfdpSFWDEebgYUfnP26P8TVkY
7PYdK+R2VneTZx8Lkiup5phIv74e+paQuEdpGCuTzPPekTEEbJdTST4klp2rw3Sg
vCSwThf+/jVua+CFV3FnEL1G9xo7H2/0aaO6IFXlXO8i/TVzZyrfhEsIURhqikIV
CQ1KdqUKViKsZgM/PYVuVQRbiUBzVtbfXMxTRv1z84pTI1LECzMsey0YDfKaf+9H
fG+aFBiVL5m5gtezQ55whvi9vfBUWbZJDdvEMScIKyhFCuOP5KGGWnlhknM+/P4i
TQe/NEte+3t9pnnuBGCCnQ+IImccErza1sNS5PXL+GgbrBOrqrF0im7TfJv2dcTL
tM6dncHPFJpi3VMurrk0ki8vJffrLXQ3ccAlSfYQV++QDgu5eDU2NC0mM3VtTWpo
sgrlqjXMQnROngvfkREJPkChMW8QoS8IOFLhEGNBop2I7XPB+7Z/J14U6OB6DURj
bt+d2Uit1/dzArE3mPrZr0KOAKKRgqtoXhWp+sRXESkT2qMx0+Qi/mSKm47KL1qs
O8AdNo+OOz6a1w0rvG+LyNcmatQBM/eNZP4Kw1MNLm9oUFELR7ua+yxoR2ulvDpb
iZytT4vq8+HP6O+dI1iDeIYi1cQt6f3q0VmrcI7nmBiYedSdmGr7qtUMhstkrQFz
zQ9JqvywiOh+DM264wCyIdA/xs9pJRT40h8i9a4SDtMZCxmYQwW5/gXOykWfK6Mq
zexWS1LxjurWsgMSPJhMrT5WjKId/AbN9WeMUcK8gnwHoefOXaLapEJzvOcsE6Pa
6YTpXl56cipkMKwsUaAkbwnK7jNG/CCscUS9Dvo2B9ztyTa0Y/AVx+mngPv85Z1U
mb0oEpglXSfoqTV2kqinShM0sXkytkbHGkNaZN9i3NvPJydgNBiXAgbf96Vfk7MX
KBp3BR7KVX4W/wesZbxiRSmpez5JZR58w1TccJWzCs2UUjRVb+xoHp+G/PUdcXJR
NXv/Jx+ASuZ10XqGpBqvyQLcGFO3SDN11/HLBY8pDoWOtMu7TO9Lh7baT55C0g7I
9sNlKHDj0+c6gahkiFqY+NhlAYS0wWMmt9mHgarYL5wnrkNg/sQpllBx4F6bKMtM
tMRiQyaahflx5/K55ZAf1bjCKtxdPOULAx63I7WpmeHvbQTeqIpxQaioRPYDQYzT
lZXfRHMp0hYsq5lDDmmgGgJi3b3EglKL629/VPc2wXOH0RKKFhMLN/MMqsiXfm+6
39z5nahbWy6wcKQP4IeNB+cDvEeruQt2uylWdO9yEqTKmJxMmISCneNPuWd63VvW
EaLfVKS50QBlG5nZIT0HbSio12/d8vwQIJ7q7YzbN54ZLzHPNNhaxmJnM6m+tSfj
plVjr6YrRPgO8ZFi9EzsP3McVTcGuZTel4JBW0xbWdfb8Grbft6qhmEE2InGJupo
Rl6KwqiLGATS48CCK4zyKAOTwSnfvGsGJBniZVMcvxNULK/I4EEfGMKaby3Ug05I
a/N4E24lxzJMW0hyre/OvT1yJjGvtGCNAf8OYdLlqSaj6nUpr/OjuMJrLXQ3SSZN
jb0/pP7kn+BVNjqd26YfTd0znnloKmWAAgEOlpvL98YIxp1DJjJ+dfqzfTYLLt09
hocroogotf6aXNt9vEv1kT/R1s32xSWxBATZbPTZNZ7qeBFs69tsyV5kNOVGrSqJ
ZstCuCjDMBne3YmSBaWAFZQQcvPJOP+R3U6DWoyaFGqqc/YoyYlRwzc/JKGk2oXi
lr3pIscwt35DvjEsmpZRHxQLrsptuMYP6+7PTpTUo4j7oEtDBSFQ2v2Ud9wtahKb
APZLZrlGHz/wIWCiaz8W3sAOUsS/Gv58mEwYO8GOnGUiq1bxBv6nkCHgkUFK/6/+
D+Xf/KjfY3PgZcThFSoHRtdMNUMGowyHUYIGlzPusyx2rzbbodjpfonAAgCTKQY+
TZLC1oPlV+IN0TUbUKABniPnIAuoRY0wl8MCPx6AOKatDDY5XSEVDNqfnl1DUp9x
inXMikj2H2DLoEm6OOwBMtpSWL59wnB6gzXVZesrbdyELBb+mdGDzaSdK7MFpjCb
ZsV4Ldp4IjzSt02FghPr469MHwuYh3qwgMhZPE5SfmHfstnUvf0Gpg7gvBEJHLio
sY10GfTE5EqXCf8fbWLgcnRXS9LbN+TABI39He/YuzLaABlvqs1k5DWmT2ZytlVT
F9YolhqIYXI3jMveN/iCnge+AFrsP9pilLU/ilR8i2Kikbd9KGj5/1ZxvaqEWTRA
QhKtMETRHeQ1pczKyAQeBTukNAjCn7hXos4apjnYVpLshtoK6K841VQl1qAT80mS
aBFaJmtkXThn2EwBv0WJkcAO/xfiRLLl6FFpM1f1O/N27IoiS4rD4yfdm460/SHL
fzZ7COqyB0W0H7MQKb9JF2lDfIeuUO8c8JZRkH46JFVAd1D+M3Z/I3n/sOXMns5M
WutiG7nDkkb+3f/ffTiZkyIufCebu3hQdiMKcUgCMv2k1wdeNvAeV2Fe0y2i4O5A
idkm+veP8MCTwM7nuVEiN7Un0qDv+MMjVz4x4JW6oqmagKxSltS4SlzyLzRvBSSn
7fMpVEPNLtK5OlIRiajPirR9hy9gqSdg1RA7tJVObgfautdQexYvKXIWSmwQcJj1
N/f4RCRVXZfSKep7E2jJLOCHuiWEQB+YJPPxPMCMfcCxdU+6zpSRC3vRC/CmtfUT
FT3Qu/0XNw2vtJ4NV2gG9ivHN8Bxv2S32lZq/rE/cnFNjBB+51eS8Gk8WBXaSmMR
4w4kjJ9QTSvjz3TCU8k19ByuRgRpLBO3JSicN2m2+qMGqHmLYoXSMKyj2fnOIIpC
XVvq032FdA62K3i1gAV0KR+mB0FM1pSNPV2eDQHL6i0EDzfBmoM1RDVdTzwuzFxW
WN91Jm2rU3QiZVDCSUecAGghFsXzt+1eJgzgyKH4uzmPFlv5E7GRBnpeZ97+u2dJ
M6EoK2DHH1fjfp57VIrGBfic3CyTCx5gYNIBIIe8HwBYYJJSuF0Zi5o8OpWhuy6I
IHvukCe5oD8hPEtFnDQGy8ykg2fDQRPqiPRN21K0gzJckNyMmtWbTjj7UhnGMXTm
vYc7/6je0xpikiyKCL3MMt/7TC5Nto/P6nVfEiTIZVq7Db8HnpaTAjjHT75RvbYX
qeyIw6t5suYgLNp9SbpVptXF1UTbasgFmqcGaMrixtVJaH1M0yfCe/UfJUzaYewh
GyOYobU8PXpdajVrLspkU+j+YRuib/fX81uMpHLMhMiUexITJRGacgA/dsexXot/
fIBdp0FR4/QyEVuOPlkzVLfoAHBM8yM4ozgo/ur9WAjJeoUyXPDKssN0vXBqCXPH
y7FVRhIYXqdMPDRdHmbItU/AnYeUQYENn/O1zIJzWlh8c1o3mZOt/X5wFVGdohG/
QKZen1Ziv/zf9+RwSZG4E+OIwkBlCA5w6FyxN1SWIfaeTFndepGM48xmCrqEYN9b
dNgKXmNpRf/QwRYl8maJ4o+6YGSgq71dQWnAVRpjk7mK9x6oXOAkRGmn3qE9PLM/
spQi7bdY63xC5OzA0rS+4471sVURVCKUHeXnC65WQrq0YCzGRgTx+b46goFBCTOM
QMrSlpNjOEu3MUCGV7kk75JYB8h158y4OcL0Ka7/OjKm1qzWACc5COyRmO0d4+D0
T9Fp/P73BOJnFqcw4kfHSROa7p81WbkN/YXxUzrycoC9DzlZ2hxxK3V08fVH9k2n
Xo5nAIspPNfQpIQeFuaaRncaLyCZ471AUR/DNlf0U7Iv3C5bXuiENJVxwMqXrXw6
PGyyFNfJZYGXrMp0MPLtRmc6sycbR8onXZSxIiSvUXpFr81l2HwaVNbR7xscubTa
KYWoL4zxHxTA/MqcYtbKCcnspqoiucg1aaA0eDph3/4Zjbs4+PNoL90oFd15JOve
A6BAA83yAHMiddDTolpPw4vyZeWPhOBblZcfhkl3XBHXTI1xAfqMfByvdJye5MSj
L8wiimyR3XjxRrQqhSYY44lRwrzii5iNVUVAv7cGceZCpiR1HpdWHHZO+pfA+WV+
rfJBtV23QrNDMwUkwhqq26HJuYij0ZFquIrXa64Jb9IUaAQgOCkEmUd9obkrk0+z
8PsaoXQuQNw3X85Y43FzAOJoLS7729a2GfGGNC1evS0oqILFbwOdAElbE2ryC1LK
EcRDzeSs1C0c2j2drmwGlebnXu+K+hNhZ5sl9IFP98kceg0VbIkAMCGjBUzRJvXN
pxpMdsSGWFGLYVTbeo/jjxr7nHLCqyRQz0vNSPyllqTI6NS9FPX/D/9C+vngbbHU
fr1tNnukgVFYp9vWl8yB769IoSBOAC5RzY6JVwa8TEIxUoif9SFnAgZx+C6oFoTx
JkaHCgJKxDQxwdOmb4bhw817qMsc4Scfwc7/GX2dc5znC6x+B2tAlBrbGGz+v5nl
rA2inp5Q3Fdl2XQTvFYMlnaFZl4zhZYBOauVGaKJqwIx7nuQofpr02PrWZ5hwe4/
+wEUtVYDueUnpMm8GutkgCttloPidbeUuFlkPGN6dPE9YC7v4fZr27QtxC7iv+2t
BdtbmNG5tp6Gf7BWs0/ykrXSsetqVHGQjMAbvhmfp67/OeMY3M/VzQWZM37vnpiC
cd0yLUxyNUjIUhcY019vgcaO8r1ZiswcDDcOpO3ImE6veIPQXbe2wGIN2SWtu54c
OUoT3BL7RawCGGhFx5WK+t6QcuVkDC7NKWtJieTcQRR2IlGoasSC/4eyuU6If0Eu
HLhxgfi4469l2OAe0Ia9WD7GwAng6hnkGAUfm2MYTtMyzMQooJdss/xbA6OTcwjZ
PgtIwD2qmT+GnRuuQBM3fNbYxaz5VutWN64WAoJjzrECUJ5kPvNOw8sTrtBdXCFo
gQdYmR+N5kxcBE834ENZt5OfV5QXOAxcVb5pI5c8vt5qtdaxeqvr+1Y5E9Jm0DtO
ugkaF7knDqDFtQFNOuPAuJa/+SEftYJFQt6xcgmOBpspeyvsmNGbzeLHDzJncPxd
jck9aEYTmg69PdUTIC2jPPW++oqy0pWeM/i/58mZRzYCNiNhNL8wJLvz9Mmyvxcq
4Y6m/84T/pHPi+8OiKlvP3EZ285thTkN4pAniKsTTWxO14ZLrcTyIAzg1VlemOX2
YLC82aagAZrRJfkFPO8d5jZkgP8c7N2/v701gndX5Rx7DZGITXPDwQ5AcpONQdfl
ejQXDWocU5eyIgXPDBgN36P9YD1LBwtfEcee5ngQ56oBqq0MvH16UOLsbAu17U3K
E6TFtV2mA+IZTVt126A3uEyCUrVhXOiQpQRgUZWeMxMoDRe9xBWOAK4ACRJmvuSK
Qv588BnCPM2TScNzYBsQKFGBtGwv2G0U3nCVFut5L86/ubnAHPlmAxECDe6TVXec
eVvs7/TQBM8cS/jUU/EyQ717X+R8yV3PAmz8ctOKdCqZ7tkX1HC1GXjvROnFEgLB
`pragma protect end_protected
