// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:37:16 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
IJpwJF4TDqP/7aPfcN2c5iku2BeboEJ7u2N4nceGtiCRvLLPxpjBQcnMrA4TTCB1
vy7DkubVfbX2Ed7A6yrDTZTw1aBm7USaV3uP3XQRCjkqaedPJF5U0amLOQRsWV1B
aTRYGQTgeL/wo8mMJUJju1xXq90ArRziYu4FGE+WROs=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 4752)
3VKEO6/OVMn+FMUfr3pcjnfgnRS5WJPNxOdaPi5dLgZSxQosM8G8sJ0X/nwH1DbJ
QajHSO2voob/PhGNd04dnvbsy3OVV/xETygFBLnEJhf/RSjuvanFfkXMl/yNJxeG
lvoldgw+x6j/kmVPVo+srg628W4lVyA/woO/qEk4JSWiBocoJvvpBcg1/6Gd1mPb
rPbXNC0RwjuJihxaU56q0CtGwFL4eh/5O/U42NPi0LH9oTFygnpC6mrkGMUTs67l
kRNoEftnd8BTQ6az7j987Tasvt1qrzF+ov4b3qLZh7iknuQ5rxsUkfrWC9L8l8D+
eV0ogJ/g8i15XCzoR5vfM/dH5UvllDu6I+xTzSWK05p1aBhv7Dwb3tnIVHtXN0LQ
RuBBcXNTD3mqR+rllI7uKxMBlP624+EZMTw1FWdoQ/Gh/+oa6SrrWh3Azkd5XPQM
l9es9SFEiw0Jxi04VypTw+4rhazXEIvv0GjjShgsmYwCDZYCHnztrEjhCg4oejGT
KqjJpvPXemCA4hDceZjsGT+2GbWE9mPionSYR1yzz36uv/9efXAA8N2gH1rZTJoI
r0PVCaHiTJ35LQfOYjbsvfPmJK4jCgoFx3Ba/NSLl/+FNm1jWWYHdN/cEC2vMMtC
/+3P5bSo0NsPOy14FYR2/H4SZ50pPqMMNKZulkzXvxdj3Ug8sE9CkouMTRc8vWvy
ak+H8dO5zgNisjq5Aolf2YyCRjb7DOxo64Cg1qFO2g5GwjgM311h4tMJEDgnfPc8
ALZzjKfF56xLC7h4v91t1xj/whOWlWkX99pZvKLmDcDJXI+iB/XmLkEmeeXtp2gM
Je67u5kbBzl6ib92A9glWLc6Sv/x9xQihpSjoEFoHbnBudCiKMsstK+SsNQbGW5r
DUeEoRCDHAtN2+XM/RfETVLGLEDTSuO7hxiLTD+JBCY6S5NLoLmZrX3DI8Fp9O8k
s+nIo5L0Mfxbnp8qCKDkYDXb/KiYhjBnIrbTxYp73ssAsbsnNrg7vhnDGCMprRqg
xY2t2ss+FDE2KiVD7d6qnh5uy0PwC+t5xtmb8qYqCzQT0tbMNiKWt2kgdDmsX+FX
BZRGSTtPdg3wBlvQdhvVb8+ZtZy12KVGrrt6QhnlXzycCi2eNiuLgzaqGv0ZJnq0
81gHOGrl8Xxxd/2gOmZfhDo1cUaMrIuxDYKrAFeucYwGg1aajWrsqR8X8M09ir+M
ECAuIeWYCitkR90n/J5WrJmmjHLJ0vfktUscPsbUsp1AlbJziDvJPtvv2eeMy22H
tC4Hr9xzaF9vNZkacjj1yzcUIhfEPAVN16PWfvMXJDZQmja8VblrHlGmT7tGpXLS
kLq/2HYAE+EE4C8a/krF69pug5/zU0WSva/+nO8W9KvM4K3xzb3Z8PXXHDf+eLiE
JHkm9cIdWKYl1EaePYsLIEl9xF7CG3hctrOfNfLJgUf7lav6capepR/9ablafhRY
90NDs19F9R8sv/h2t89WbOMfGcAYft9cap9Wt1FZoqWNw3BaYJzX+Pf07dx4Q4qz
/aHZS68qw/uH2ihwxhcgwomTsX5kN2dc/XPB3MDgBg2EGbrbNesA3Q1f8Fr77WBf
N+W0QUg5VNswRPqII3vvN3Dppxn8BtZs322ULdvcn7/61M9FeThiv2LC/mqvKXy+
l9zESVjFEmOm3tNyW16BESnSgz32yby6RPv7PVV/bGBI4Sb/7sJYDXZKYgjk/EJt
0xbgtPHRgUfUItQmoFq1plmAyahEvuPdoqxg1TbVgsoaFd6F7KIkcfZGBfO+IsQ+
C1g676Q+pAMXYExZJTv5Vca8Vs0lp/28MA8ckshHv/kMOGCXYbnuWT0zunoDmHLH
Zi4i6EQriMljz4MiuVLuBpeyGsvW8p+PgCC5iVnnOU7H2x1vZh0IGE9ZSSGDS0OT
islaVK6YIFW+kn6tmxUNXAX9GTMcJ+jFlOacx0ProQgwog547gbYlvh0g6GlWab+
cO+MdA7U8TXPAUkmnYaZ2RXOLscz9watQcteHCseDlQiukmCkyo6KmUDy4Wd69XZ
Ifr99qtcS/P5TIdu1j6Eb6WvGyEGki1TuKri4jI27rMYKoymiFnouYI8NBW+Twhb
COz9nQ8E1smScRRErsR1ai2Uq7E02R5guy5LQPexGfPgEc/mgEF9dgdXiJPjEsy/
UZD6rjYHB+LppgD/Jn9Dh65IrmAJtOZ+WMqNxQNsw/e/SGeZtwrR1Pf8xaxCurQ7
p0jUFMDCCoZZiUtgOvgu31km6lBpwNPI8h1EJjGv2ckFbBLhIbtUf/AjxAFD13HN
Xx8j6QW5ub3mIlmnB8DGdINPOtvj+skXvKt23OwkpTxyGHcSa0wKfs89cvsqaBF3
dv6PKbtQKooB9odSVHZZ7P2Hbc0OErIXA8U86bcPyrWIlOCACTbkVzEM39tyOQfl
NhUcGlsFHWCL+5jNScJeJhQPj8LlwYPTqRA9CfcCEb6Ith0EZLyFQqjXTFgfHXNn
D86WuC30SevPxmOPzSKuwudG2+XxmFI4F138sRV8f8YKppNnoGjfkFPkPAxNqXif
TtNPecN18j+r/Alxh75gZVFyyLdmT37XLZz8qTGgG0xB1WtZwrc+DDHeeH4aY4jn
AvoGmVukuT5iHt2z0FA0UpOV5+EKwxiU+gqvS9IT81cRGIX4XfhtOCuAV6nLjbhf
vcTbQRpANKe12hvQWAa6zQiDFJ/5QuAyDR//pBdvcM+mc3EWN/yhUwGGHLM1uqBp
NTFSkZjJYEGnb1JJHYf7OGjsoXxzRdd+Ano8ixCaqRBXZczFyGUIWS1xOPYnRlCK
nqUfRtmf3pBCRXoamCapT+o7lQpknyr0JU/H9tiHihTcpjsKhvH1Jk4ejVADu1Cx
ASPH2EsNFAHrlO9Z2aJQZk8XnAlzKtPKU77tFhZsA7BiAM0zEfrNqzbbeP0hTOXm
J1C8rz5I37JT5vqkJcrw7Tw3boKMRLTjGt5E7ZH9CzaFAK23HmD5luWmGN/R40s/
4HNqz1/K9zDhDRa13kgTEVbwzPyI7Rtjtd7vJeuTyDQc7o6ndn3bA7SLaMfaOWRJ
feYi/tXZOQlf52iX7GAjuALqRD3ScDeQhrCKzBmyR3oAA07MLj9aT365aqjLW3rN
vvmOTsthFcU9+mrqf5MXQPtvSJpd6S7dDmXmtBvR7rWcjCpSd03sx5E+CeXKTu9C
ModVjg6MimzakMxbwdPwRvQ208V/Z+xbm5YWgS0j13iZOcAlw85QMDPdYDOlLWFp
4Sru3GNJ0sl6/1ooe64iPL+bCYzwE55a2jBQsUOj3RFvjoRYs7BRo0tukh8apCnT
N2Mk/RqP/hF4KOvAMf1VwEd/mEO4Xw40OXterGm/W8UaKkoeuFGH22GWvebeVmLJ
N4st3bCQTK2cgOKpWY+8FkVMN+bgCPRVEG7D4HBW91uQ+jsCRcFY1ncro/+NKHd+
ovQOJSo8qk7pO4gkqvlicgh6FkRM/UyjNUO+Mlv0jo20OP5cb+Gwf+j9OZL+mBNY
fg/2DF8fyrqX8jypnubzthCAIgzTvcY8llg882fdI6tLlEzuHinrn3CkTdTxl+df
/X0RHLoge4s/+AJGVvUgWs3fOqN3O3OFLbP3tmGZf4Ih2w28lGHk69/JlWCEEJCv
FlG+cMw6+aEE5DW3+bkQGbUB/LzeG88O008ss61Pe9UIUzoWC6Bs+187MIvCxH+a
dH12NlQdfkFHzppTh5v9EmjIhUdl0dzIaN1r4DVUnV7cWzZtq5yJ+yuKtyzEft4Z
80tqHlxNQkOze9Fmrs+CHn4sWumbYMGcdvBYXN6bu0jn6slRComPr9t5xgAfWURH
QAZoavHKl8+cfPDoGMxKIqBuEWn1Ra1TYZ+gBi2YYGDtkKAjEEJ9XF2Vb6fo/GCp
i69v0dJ4uM4JWZRD4K6pe/4G0gb0GGCydtnx8LccRdpqzdp9bFLar8+hdWTz3jb1
8BoRczSH2bjKl58p7cu3lPls0JrUYUVpH9p+eAWH2aS5e23FBn47dKm6JJJUt3FF
Dc8qnpp4wGqVvEFE+0DfT246rawcgF+K2HsEQtj4Zia5coiDImmAhS8WZRkldLLr
5/RhZzXQqW2GaD6fzeJUoqpx1AK5wWkRd6iOIds+yAoOzLOK/M93zCzKQtYuIVvy
jyFqhLlWWUPBYotsv+RZRY1ogXRjozYJHLwkf7ZQaCxzx+RYGeVojPhRDYarccrh
OGeVphqaUAdmV3dsl5l/dNsc33M5MTWURktjgMo4B/LA4DSCjf8vxOi/vbOzcCc0
oJJG1l7c5XiXPqA7HKkRmST1utTAv6h/PiNnW6tW1jXV0P+NBcd6fiYc7lAKyhcV
xJZnRsMuI2p011Vi5YaO0nW6symw7+8c4eK52SRG0Sl3itP1G6JTMuXyCpKZczNT
5RwxxIVL8QapIVRjew3041JHMHJZAoG4sGEAmPBoaX06C0zxgD0ph3tXn/ZLHuCr
r4FZdaNBjn2NHG1bdOcYlEK8Wcswi7Ip0up9TSpS8cbRYvJu09DCR/LCD4H50yUa
e6yj7SrP8bpRnrhc3ohbXTVPJBb3X6Uf/nvjgTocCFtYF8QmjfakLaHv+Cm1/oJn
9Pb4za+DdSCNqo2aMtlUsXVHl3OsqpBr87SB+elsYH1wx6xYMg1nefJht4FpdRaT
aKh1RkQ+FGFqB7fQqlT9D+8HVvc+OrumvXlpVTQ5oz2FkkEBkNOfLL2gK0oWwtSt
sWFsH+jkmaK4wy9QEmBiYtTsVorw62N09mi9119VCg7C0gCvqzVwiEcjfVREtHGd
XZLzA/rPsqMRubVFcfkuMmTQx5FDBLT2Zn64z5WyXbyGf3+TleOeJEXBJ1bjnTAS
dI6f4wFzxu3olI1b25cb07vE8N3+Y9a8eNkSy7f2DVQX2aM8amqf4LakzCbzz0Sw
XgrNkbiiuJuLsOlx1IZA7y7pcIMFkY0bOlFlHfP36NCGIb73+No2mwvh1Qp9pwFO
XHSwmJlKa6UnoCnuRa+owiT94uLCtrKVa9Q8KDaI5jjX5kv7YFqeBTblBCwQcwOr
913e32GXU2NPduR/ymgnQiKT/tsrmCml2oDx9UYlIYafrM2rLaf0m3irdoK0s5KM
NlUuHD7YHiw4J/10yf4mHEAkeZqVKVDd4NTP6Dop18aZQlQqYMDBnuVak5Jik4xK
/IiF1ZDE07Odw1LR/VAVnIovaiBKVe4/NRUKkJrr3rh6MvV0wgRWJv6uk+pVbBut
miuymyzTM0LSg/QZHnI3udGbBoUIW1AvS2OZHLDWgUHt2y4DA2vCQAtSAc/hNyUv
xifS0wPjvFsp6ZmWKq9jv1/kt03agdJD35CVcI/Ur/zTb3bZnyQwQK398vXgzbNQ
g5lBKuO/BaeqhxOx6BdONZ1gfZls8nOtLQG1OdZ9uA8AF2n25FFPUj6PVXc52Gdl
oOQ0/aEIvRWwAeOOK3SdtDuI8w43y19X6c91JOpCv6ln3mnNFqJCSJrh2P4UhX6T
jvRIO+CFcQWWXO+4I4uv4RQtfofUBRQpEdGOnFQXd8CfD4tRDX3KR5jrrBqAGwyF
kItbJRxhiF4wKd1BPRSJwZH83uzKB5eJNP1WJNYNK5gzfJlcyyb7xAMqctuFVtPt
+j2O6EwO+8pU/2MqAThd77shBNkOdziy0P3NOWRePjrIVhIAa0FScXfF12yf9mu4
cQrvrVrlK8MhXQVFWWilxSGJ0Hm6Fa+HRZVLvd+8UZ1sgTR8iCYz2zohiSA1ZXFO
utnsaa7cllT/5i+QdFQGBaXJ/INyQQyAXkpt3wgz423YE5WuCdCHcUZsY9OVVeuS
U3VLAMAWd81Y64TnCRP205Y6GTAQa27BuPPxNnqeOiSYkljwMHh0W5Ryt3uqC2M8
BTK313o/RzrmcNvwHEgoC90kMfvlrsOZqufVwjuJA7xK7Lzz9RWhvnEQRpDHT8dB
uqVZaQ9b3gbIL6Q43rpSlAEcE3NsETzNj24FLPGfaQJUrYtvrQOTnaVmYB2zJz5f
2YWMNkqBg5yftuTdute3zk/slk0O/AiShE2DYkOh0+OMLEwjnMuzjiiHWFdBbeWs
V4gct39/JVtIqPzU0apK+6QB+pvjUO8CvlQBIb0CyQHNmX1oFgYOgY0qFHejWXvT
1zZYQvd3P8LIBeDPM8NZ+6piGFR4AxPjXykKWsENTtdTOMpOmf4CYedQNG4GRhQF
AoWk+zJaCx6DRDTV1ztAaZcj4AE2cuUniQ4sWtG/5sXoA2k+b+S3Rfatik4wBY9M
wakF9hD1Ch59kl6/DRznkvUFKp2huZljC9a2WO0uYE98HgCmMrJ1M6NhJ3elRl/H
`pragma protect end_protected
