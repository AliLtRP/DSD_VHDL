// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:33 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
SctBAOFr1EsL1bv9381bPM2JFai+umro+BmkWoJ3wDo3vVWugSLs+8C2CB7x30VB
UIa9o05yaD4f3k30mLVwvD8tazi3qwdV9GZw1ztFRjHv9gTYzCEyupxZGaAbfKIN
ThwCZeMrpgPC1/RI3wemBsfXkihKYqwyjFfS79Nrvak=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 7216)
26D1BrNlflE1V9sj0/uyBf5IYP2KNRwDQnfPSc4QqbH/4F5Oct2rb8rOjk8BKqTh
vSOax+Is7/aqtGw8pQQfFOGt980+LR2HYCKdHXafw0BfXEjP+YasOcjHWcaJ8ZSu
IFb8tupiPr0jWg0gP5HNj2Pbi7brbYb6YYx2FyFh4CCpQTzZQYjuIaODaa1ae74r
Cu/nHdG69gHP02LD3e2yj229h5Anx8gy2VyNjESe3l/f44BsdSbCICpp9SFXsCG0
ub+dAzuDPgQprs6FZp6I9i4itCCZfDp1Doc9+Zm/S/Xr2i9od4f2nFeMCjUTfjSy
CBkNaynKD3IMzkIdkbN3/aTY9xZS4jrXjQvnzpkaAqcNzdjrfUO07Zdrwi0nPe0z
X6MCmR3jJpjR16GD7MEZwKcqvDcjyJaFsBjFqKZev8/4+3TPEjD01gpZeLBAPvYm
F/k73iCAFhov8W8nSx71gZq8+Z80rk2TBr5ns55W5/sMJln1bqw71lb92X5/CGB+
1RtRQvE8LiY09nc7FvB7MvsA6siv7zX0YYun5GX4yv+w32tG9I3C0ZAqyryWWcfO
I9gXzNYhOOcDj7HrnW3otRahOjxSoO2st6FRDpkGfhZc2zIVbw4MuMxAYC0pW1Ga
ZWb6wxpkaW/9GfobIZRN/j44aev74XMtDB+1693yDa8GkAflDTwwcGBJVcJw2pcY
QP1fcJ87LajR9zmog1EitKJgmuiqdJVEUs+a4DTdzecCdrNk9jqZbhgZYnjMsgnG
IZLCISx/hEZ3oJ7frL+VRR6N452AaRWUo07DvIv41J5UpO8PcI4lvUCMzy0mU7jw
MWkr6iDRoIc/d37rIPnm5MLV08QKT50YYkQlrpB0Ewbc3TLdiY3Tk5d9MhLuh+Ce
3IgwTnkJxh8m4DlYZv7o+CQVMLm0fIi70gonf6i+6CPTiNDbyKQkOCsLumN4R4pS
KUqXV1eCWKHrI7dR8CPZSDOYHwdW7dJbQxt9Ze8IQ2hsJHnwjFo/VA25Nw6rJLWG
Qe9FO2fXwTmqoXSoIyIhB0y5mx4rtPV8ZSzclnx0AK6z0H/mYlqyHi+yVj5TqyYl
tYiufmqHBtGNcMtuxJY+W4LN28F/9m5q3lHI7cIzqlfAvWSQn1L9JLZDOzYM44Iw
yjE9tgEHNjGQHh9IBZvXdqjUxeoUSYUw/jrI2rddNzHFxkqDbACZif/Jizb/DAkI
60V4HCNh2O1Udy4ebUfep7hDpoccxN1UOj7FEMjvTls6NpoPSZ7GZGlitxtRISdQ
Uveyn43kPb6i+Jk4cdlr1pZIJPTgoqCpPl6DIaKASGSdQKVLZFdyhNf12V+DjBkB
b2+ICKJocveyXOEpSwdoAethf9U48bhFGscoK+v7+PU/Zo5LClwKRpTQi9JrxYrq
9hce4fL+F+O9Xn34yQxEKA7hNYNg+XoCU9T77fa474LDbK4yh80y8RpVWqvTelyF
IWU4DbVMjerXJhdLhS6KqT7sbVP8VgkCWN0Jv73zWOcS9AxWFeeO57I1SqZsCtIh
BTZSiI39py11bxh2B8o071qa5d+JnuB1Rm/w8G3mPqgSOc8sXWkJWcDybhmH8Udt
jeYXXm9lHHTue5/KvQeRuBLQ6S5fHz/SaUYm3hOx4CFnC2LA6SGO9PIPZx3tGRU0
KgyYjUaAdBDXMsF+CAgQHbO7WwwKPbkZTMEzA8H4ZiGan0Q4HfrcJwg70s+mnQ73
oxuiujixm2/V/ZrvG4RWPztrpb+tEUTe+z8dbc+/ZRUMptrMjLalD+P+RJZptS0N
hpY+X5UnOiGyyyEfUym2PEV19LuDamRRvD7JygoPBS5PZuXty6ZZq4yYp7gkE7kJ
A1roLh0GGun2dW07L5a6+uqWSeuSLiTJ0xO2L0VI3dJ1cxOXEa5XREMTWPuutfOB
PNxp7fVRnb1nOOClfRNPquoFgUhnpWJ/hTwY6aOSNAKukTBlmoHHILFsVMTwIwzO
KzEgfKlo5DCMIDjOhSZpWzuB0+BMOjM9Gi19Xo4ze90oIYcXMbk41Bi0vHp8witd
J92LxpY3kitgJ2JQyVdQ33xMuYFnrk+lB/camUft6O0FmQty/VT6nt1XnI275YXA
BfjVrLH3I55tqtg5X3hwHbLmcjq/nsA+8PWe6RNmu+f/rqp32BGd1ieUGFgINL4F
lyqdPRemguV0ukLupQy8QXAnWEZWcpAjXaWLkOSdRk6/FmN3i6Gi3VioxLZAY4tt
DXISHLKkk2y6AJ0W06YQWlxCwaBOn/TqAlZbJpMoaKwxW3DEgWaAqPcpoBxfV5gZ
Qwoqk8CJQ4g5yIPTP1wScp4Y7rHVwT6JIN7b6cJg84cejYVxkT+2LCRqpsaMk0Rc
rEi+0c6Z2H+DJnKFPUCm4cIUWc/dGUspbFNgDE99MwRQ9KMXADkZPpYHLhD3hVb7
RF6P8IHVDY5jEIskSeAnhMNxid/LusEfCJvlruB/eGnthKpXn3H/ZCJyuC1+5orM
wj/8GMzMs0yGKdmqfwmRjdRbfvjs1e/EmLD+wK3/XHYKOQww6aVww8SfjTtf/XB8
zHJ3jlU7Bt1HCDle0aOY0PMCuDboSz4iphCgW66/9wnAiPRrcl4m1dfYzbEwG86M
kbVrdSsh01o+eZvfC8duCGTQPZRTYobEMP+bTP80yv8fIYkPymWA8okpGi+V2ni4
PK8QI8y1T3DClHpcfFNXXbuZS5hk/58dvJLFvDD0/iQAPZ5S7Xvq7W0iw3PISr6/
unFVD5LaONL0UjEuACk68f69pHBnSlrfjsGd9EygoZiLxjgN78BhaEdefLToKILV
MvcX7CYLNtjE0qDdj1tLX+vakp009I7ZIcDU/o4hqan7F41d0Dh23t4R7F0P9NnI
cGKM2/Fir2skKhL7pbC3Smw/F/rGBghCrnG3s4+dhu4IgtDqBRvqPvGjdqJOxDjD
lA8pZR6uOuqi5cWDAa76MeGUU1QRGivDJF7k4GaK53Ttvg8YBj3hur6/C/AIgOyk
1TUNTSnxNON3T+Kls/3R8bQToBLxc9rmSdqjpCV1++WFJk+aoGCTKgL+WR7CxSOO
UR1vLq7mlm59TdvsP14SwD/OTD/xgvuUX3FUpdaC1zAjbuIudVYIaYDMv/dYpWSa
ztz80qwMJ3c7d3P0TPEZVOR5pOE5WQjokpQIKewSTYp3eRcECodR9EO9BfSNRYE8
D1ECLBQR/sXYRA2YKS/wzLiA/OolZFMxkO5pdL3UGtQhe9KqC9nE91CW8cUpD+tA
ZN6DWTZoWFka4c7q3YPMAvIj1jTZlx1mpZtnZr5URAexhEUchY8kxNBrwKcVBeSO
EouLMPfYIcvTsOiRvJ6Tkg2k+EQ1ccQgF9CXEh/2ttYJPfVFY7PXSuPJ3MTPcdrZ
yaH3IthCVM2HDLUSWB/GvbxoGRvyzr2581PDmedx5073q4Y4Fa8uFguAmJOMxX0z
4R6XpSPPDriKo1t0aFulfZx8Q4kovfrtwcuskeXP/tK2qQ7uxScD3HQ+asVbmWFB
knHy933PHxqkvZCphBWOnAJOhbNEql8g7SucDb2cpzvxJulH5hoth8o7Nq39QMFc
6W6vr65Yq8mDv+tSKZl2Mmxat331OtPFDOHqjxNjClWDyhA7hjXhJLRhvLpjCLoN
gdAJl42Nb3ce/JuMoE2xqla1yxzoJ6oZOTKIiOe8O530UtAo69GUZDi2R0+1G1co
iGycY4Sa/xTW/WMgkR4HojOJmeDp3jQdC3iCGY9pVfDAbB+HbgHrsEZYS04uxYNN
3UTMYJfyq37AXybMx86UBF2khTisD2VCMNX7J6UWIaPI+Tdp8i8PEJTHGAfV+hg1
F0AjotP9VQZDwnjrEdFRjpt4VIPbZL1T4w4U2cryDMs+JT8Qa0vPrT93RW0bTln4
0J5fPaH66IBT0YI87F1niKVdF1O8EV6tTvgEIz34EESBnSZOrdcLrm+KN+Kju+K6
ejlwKXbfMzzMzUdALgYGVTJmtq7aNNEgughOEdq+CpaHArGnZYg2Q+QoAhcLlZu3
XRcDdXm87IsDeQ7x3d9A+VTnYYYfvE/0HKE5xxx3W55HnMH379H6BM0NdBKdELEk
WIn8b0ZyZmZwk5TES35sxnXBmz+xO9Bb/sr4iKqE+NGDIqhQW4sxyrJFUEAnqfRV
ds3VYHcE3eeHutZssSMxbuHrJnVLSHR54GIr0VqGkGKiuTLQeHdBsT/nAZkEMK3j
fv+xEt0eXpEzRgDSawwLX4f4qSmocivIbejZ7HmnJrK9La9U7afeFRSg73AtLbom
1AsBfKWMHGPoy7LMSF1QbNg9Cm+e7L0E5iIqrdAr5UXQwXdBbx3HIrCAdb5rjF/f
IvTh+yOc9zQFAuAW9gaPwSZMPPhVwBmCzGbWyc1NRPtRDGViLeOk6Nb8O2xQBDct
VozAVBGpdvKeUwKNIB9tLCXk78Gh8WxNQIHGWLf3zveHY7NfkrRwSm75Jci9QJqn
EuT12f8su0ieSKXMxtl+z6wxw06Bd3cC6F9C3OOwAkrCRi4Sn8/BfCsg4Z1uJVSN
Pt023AVQjIP+pRqpvRUUNyoV4l5kj+3jZS0yLzp+S+A6ObmwHfSKLdO1UOtJqBYE
v51U65apiCEbWlioU2fwrFlWt087Se+hWC8KLgqp6g/S4Zja/cKGzAyiH5cmzJDh
jasA6ioV5ZMJf8GbNBNQI3M2OjrP0esaPDW/CgbHBhbktsIfVLoLzNXZlO6NUpW3
zYffS+ngBueXuryjTZnyCl2BrlTbQgsSp9LUkwTgc40/hSJz2XTREUilMAuvEQln
Wmsj+UbRGwHjztC/wclprZrvtsAXjNlajub6ogFWrUjp8i3c/BXmPv4fngelbJBh
g26koesqKbSzJ4qDiipamm/Z+ByweOaBcpzlsAsa1ybQnTxzqe8bGAfD8/5VhYAl
x1z4Fdxc+/9g0BVQDq4hS81nK9zvCT3O4fOW3eEPJTRTsdv93Gpk0K7WLzVYyWSs
Mly4Ffg5y4FDdmuyoYkLkvdw6TfYMq525nUZFL1/0eZsf4FaojSmRvhKKmjN9+RL
83TRLl+bEebapgO3VMHNzOiKJ8EMT0jHv8+EnlUdEPRla1lwDDCwNZGwWPDsWC4u
of77u4F25sMUFo0oSrLrwDCyHuYHetQ9uVjC+e1xvMYnovJcAtZFLJ8gp61crU6x
n+iDQv5LLyqHyA0Ut/C2dwlCbewwIYa2ujemO9DP4aFRpzvXwUF+ujSV6aEA1R81
wnTd7vF6p3EfMKuDVMRz5hn0Gf+FUTCEde4862mz8LCAValsOgSQzyAVk9UkcZ3B
o8bzwRqgV/ve8cjAiLifHM3j/vaR2ncdGv2s4Tb29mkrhsIcbD9Ba+ZT4k81P4RA
j4yHEGPMVMa9Nvrwcv8uM3pgOWwG0v0t3W807u/lcZ0+vvEcOqcoHUi+uwf7Uvnm
bmsMO2afeqbk6W0IuwMn47Ec4ockdcdesdDaNTMldJ1QFY4xRWlQIWgp1NjXLDxm
0dF4Mmb9vAV2Ox/msOgmkXts7WYBfglg735g4l/0zDN2j77W8dmuTEqYTsX3Smov
VeqB5f3jF2YXtPSlbwiqarrsVK7itcCgNqsDuj0skudBVh8ouc9dYW2ULv0IndpN
rfTp0uEBRq/J6qLEtICh7VIFOKMzfNITmMnSf7kQdyzrKLEwI22TDuM2pnDm0uzH
0Vq+AVolCpvev7Q4E7NYevcv2w3IDMSILHB8jkrMigYVpueYuviG19MQL1BQASEu
2LZZUVHk4zpFaDUrkSWTBzQhxW2obPhqGCkPJoSU9jNY5yppvwiO9Ks4xxDeH24y
PYQYYHtScwS7XCz9hs7dvl+qy4Aag5ivsHsK/1T2k3HN8FWeXm4LSqpJ9UdiNbG8
F/6491BVxG5xNpq34XuVemjDJihgsgRLgXR25g5QUOD+jQmVNxvC51ZK1RUICBp3
1/ufI0+Q8vCw9lq9CU07nhsyrpqQ8mBd/c+D/kn/vjg90vU+io7kQ5Mxwi6Rfpai
vt3+eYUcte8vJPQKckbjlvc14uXHLClAJuy6HRqeLA/Lc4yUoQCyD6MZsa/kqeJw
hvW7BRJzaxGUdd1DLdZcHeCRXgI9JB7IG/WbTLRqxYjnNoRMSoZmIHEYI47iKbGI
w3usr//lcLdmPIJTRn28QulQ1u9eMDZYoudqE6w9pfOvLhq6EfXpk9q9QhaV0i6B
U32aCnjUh/r85ZHncgbAxQ7VR9n3SzXnztlS5/+kQ/CsBoKrGpEHHrdbqdl4JnMD
9z3A3R77nEWoyr+l5KcWinVw9ewspr6bJ3nyjrmk1oSERvmBd8SE/i3gS05mkCJ8
vugpwnvzkbw3qlsjTEYUW9UrBJzBIeFhPpOi4TDtIhZH+A2uUWtcvPw4tkip0WHl
4j3wWYxcMO8JmKaiFzSGhkfaJ135rpxfFrHLj+YHVdcd9rjbRQSPpKabGWntMRl8
XzM/YhdGexbT97yf5gCOJVOI8kAbQbFFzUdyc/B8GLQTSoSh4XZxZg7Z0v+hrG24
+UJFShEkepbyAFtKelWXOG/ia/7pJFNoXibHJ2XMwq2i1W8J8GyNFKu0RynwovzX
8lxXG44HhzhndrK5sAKn4Zj99d7gcZ0RozDV6DIGMnbFdpnsfKBn93BIv3jv4U6Q
k7C0m2y+im7nNGmlj3f1KDGoms5c1aL+/NWoDPjMhLZteQGzfzGhHvuXOdxBGiGQ
jON5UbVqQ4+m5Xj9HnlXsb2OfOZjazpoy6RYnNetZVTczzh3t9EMOVgnwFv247Mg
a2nSYj5lbrqsmiIR1c7CIrFYJ/8sC/OPSKaoyWE/iT3B4UBRcMOVArR08NgDx9Mk
e/tS5WyQNwnN09/DSRxg1Q2z12WWD43z8XGH0zi5NJW/Wy9HWP2LbOKLsqiaZXAW
XArIuIDOQxD0Tydu5G8ZYvvKFHwKkRGdfSo9uanwX0Dl/w79SY7zFOXbCWiIW0np
FhjvBtxYBOFp245qTyo/2hN8E9xxMNtU/tNuuE4JmaN2+F6XAJQCpzV361qEFbTS
IAnnRvDxgQXW7WcbUYUijsbrMmDRJa/XMuuYaYvP8rOON6o2BqDDgckcXM4brNbD
jILX+6N+Ttppz+WtWnKvUuQ+P/n0DBvOysXjcpkhz/6DVY1Nt83CV4W4idVyEEJp
JAEAUaaINYXH2DYDHMgBXLRX2ASXsqf6EC57E1WU7/b9Sgd0JKItJ1GQ8zsvU9Cp
wJIMDTpUn3c3/7d/Qu6a7mTu/4DMZEv25C7KKjhYIvZwajz8Bu9wfgxdYji0an9K
64Fb9pqCYUyb2zWjTsTv6AJU4IFwf087SAp0OXDJHq3/ktpdi5xoFuGWdNGXgjLi
BQlnnf9+cmG3byZrZxPTkPAklS2Od3PGkkSKdLGszDx3B8XxTblPouAcb47CuQg6
QedMNwFZk1xFLrx1IjePTLnfLWZ8Hv64e5qH/HcoNbIc9LfBD0emc9K6qCZKEcNW
7l5KUPke6x5LabmTTjbPyKZ3U9BUhfDQmzfbOKKafCs+Yhk6Fy+rMJrxpJEuAmSO
QHbFmVDwszChpcYRv2FyCIG0wAECtAYJIdf60WxIg3k5B7hbxW7Dn56j1sJGfCZ+
9Ve42sQqAJlrsyUlA0CP0Ymw+H9YAicBap5JCaxq+yXjlOofQjzg6zAerRwiASfb
zUcc+qsTDGQkRC/ySWHQpNKF/1kZPQjdcZHJwm/QDUaTqn9QM8MgDcBycz7HTfvw
BceF94FrVeyCgoROBJ46DAIWTgwdGJzY6XHpXaBGrAyNHaoQsHWBLit/rxLXuL70
3AKSSOema8AE6usKjIG24oaqil2yyaT8KMi/YHBEddlwSPd2geB3U9CvaqLX270g
FwNC3IoLc965SqYYV5Bl16NcHzZOILFO2Jwqtiec6wKogE8kepOOQel16xYxmdk6
BnH0v3CEc9jP/Ueq/S1JUVCVxejljULHsfYZh4X93cg0Lp+J5Ajs5mzxHc1K2aX3
J5Cd/J8G/l37uqj7mq5y/4sVlvwilFE8ub8dwEkM1ysTj4VePncVj9Bj4RhM4pW7
LgF9rxU6VvOyZRpzacb/DQHDNix7xA8Yydt1QafSXBu0tfAw/gHr/AcJ1et7iHPH
V0eq22fJZZhhNlYvqxXcVoXQIvCmlV8UWwzIX7SP0nQUCCFeGoYbj8uT8rFXGo6I
N3HLBEtYQ3kksj2eVkF6GRKWwzDhbNr7c2pah+u3Y24EXM+W8CTDhhssagJKZon8
yNaei1TeHYfTRSpkYgF0TEetCOhtEvZKyTUNwa1pMzknnFqG/eSjmbOeHlPe0eec
VVamIKnLDo582Y9HaIjikz1KMfhDZGR+rdvWhyVy/j3uDhj9pLm2RpxtXF2I8I+D
+yYVhLGCNcKBtnnedngQxhFu4owXUpG6aq8b3H/bMWUkxkguohNzx3Nk/j49/WYT
3NwA1y6kyfwEbOmYrytZOC9LpLLQWr7XH0K70RB3JP5qkzF/TBQepKokiQbAqRmh
cdapu5Hhm6Ax2rHaTLqY+iQE+N/hPnO+s6EefY6iVzRxOyoeYFMGnXuwMd30AeaP
CeDjj5uAcgGAv+I5gis86QklESYjywA79O9+79F66TO+HvdwW/75+M855AFCOr0f
JRa5WqGWj5Fexz3OFAek7+1TskiQMMdSwVoBUI5jvlf7LYr6Lv9jmlDhC3cXiwgc
5m54wMcFXSMzvLBcl9APCnFrHwJVAEL/knQJJNx1YTzrfTUWpyVnskvyfcDrtNWu
R7A9w+xGMW5PngeXpuaYsOsT6C8XTem7Bskh4aeBxuxhF6QPE2zD2fnf43MEQ87a
sASFU4rQxY4KZv09Y4ogrNemO8TdM6yCe06km2APDjwHu0zNWc7rYjSjsVd+VKLu
je5e/fLI6JHdrmkVecqHn//Gm+/U3rlU1FEcw5w3/t17A1VCZQQnqF2LxLjZZuGn
C7NuMk/7hgTtzKoYd/wS6E3ZAwFsYh4ybBQGkG/8cEDHNmlClmt8hzH4W3GrQaBJ
aq9LlIDAhUYC8fmYO1rpl708ZjcJSUgiaLr2H0kl7MIZSRMmmryK89iCCNSVpBUa
S3McQ7lZj1EM1VNgOvfNt+AtggJP9ULWAtMxUU6Z2PDhpzzGKWubMYj+/Taj+6u9
s7FZEvauJGMiEg73vVhUvAGvD0//5nOiDO3ojrb934NEjq/gZS2jnNdSS4KKRWzi
aazat/mWlfx7YKqTgCSWweayt0tsyGAbUV/lzLo/5MoWw9ghpRgcPU9ASCtBCflI
TbVtYbdiDKq/9gaHkYEglnptCIb0um5EE2y+4efVwk11oAS3Ew2OaAx0HfJoSg61
ZqR81Y39Drz0feVkQc+uK3eTVNkvLQonm9L2CV1KHAPV2kzSxoEutJnbi8rft+Cd
8FEdY3jzcyTDae0l/COtuf50F63xUJqCXbVpGVuGKDsfvLaoajrOw3EZc5wOgX6R
2+Nj068NkRdbq3/QwB+LqXb7sw0KK0tWE4mBkKSQDIudIA0cBpfy7nR+t1jSUV6H
og1eqOk1iXixa0BCSYuCH7GHd4V4QMKIO77JnbQsu41IxgrMR4TbWp41lN51pxFb
NokoXwYWoUT4zCURiG+0ow==
`pragma protect end_protected
