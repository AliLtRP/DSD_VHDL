// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:45 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
pavjFT+dN2vJD+ev62J+c8OZ29WBdYugtTmSgNrAcx/IqxGF0JkqbNi5oYPEXvpn
zZbor9rBY0UbYlO+SJgwQDZ8o+NMiwjRXIHZ9nUI1itcxrHuQQK/J/MSm7VOzNcR
jk3dIIJENVhrkJGoi9+sdIuF5Vd3w43dUkbKeR9Mn6U=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 6784)
ar8j5AWxYIwLvNReN36sPrfR5szq5Po/GTcdtV9zAjKnbHP0XgfSH74h85XlLNmP
N7hb/2/LdJvcHyQJc/dpn23dPEfGMqTbXRVl7DXRIV9j+GxNOBNCeN8vJcihfxh3
9W0n6Bo0sJ/WtMNTg6dp+1X99V/BK512aaEsBsf95J6HjuFcbRgk/9R17l0TIhG1
MnF+as8Yln6dn9RWho8jF/XBgnCia+dlgKQoP+i8SRSI5ptRfbhTEiqOpHAIbvUi
T33SLXEfVMaXUxWfKkwrj5vYrKX3gY+lNLS1jibcScLLd5x/W4nyQKYydNl0CkoX
c6eStEWqqy7f0W+I9hVBJpsi/h3ScD9jwFLNb424QpZtp0X94yAhRzKzF044h+IH
vHIi0zDEevhNhZ9E9A7JuVnkVobKINOCMsIT5vW7avIH8by85uSQKodnv5JMyF/5
g/5WErCxeXd3x4yNIOEYYfYY3kzME8psD4izdpcTKIGrrBTChjB6U6jH6jHWT4+K
VOnBco2TnpkiwoBa7DkJ7qNlKbLRwN6v7imq61fglgqPSeV7b6J1dj7GPmalcEgQ
izdwLTgv3rIDuXPr2iYDr9EbO077a+XdHaI5zzgNTCYwbM5V5TPf7RaHeG227vIi
3MpDoiP9GgoQyxKOLA2AcXKUzU5da9lxfzY+wSOP9I9YJigTF3nlh4CqxDwiAl3A
2EvwOCRyYm9GcDUCxJV5FlfgCoN3cFJFYwD+n0LhJQs5+qIXauBm2yBCYQZ+Im0A
c7Rkeg2lUriCp6RCDoi7bc/RDCQYgb8voYeTLrd1r7fvCf7TS+uTc/4IJyeXE259
Ro8guck9tpZ7cAvd7ooCFlCCLr2y+CDsIy+S3Sr3zITBWTeHtCKw6xotWbTY1IiA
WFXD7JPMcTtAOh/9Vp7DvobOMAcICHmVuo2NEUku7PFBkgoXzUPAIMzEh3qm0lqK
kll+3N5Rqjm+sRWwKN8BOKU6gua9ytDFyq5cBc+VuPW5HvDeU4M5o8DfHVwV/dsm
AR4lDg17TrYPWs8hJGFjPiw0ZpdvfnNotCB/pY7vnIhGvldZ3rbzob6Nh+LTXe5v
Z5aBSclx8qj5jJb1CvM5JhtkbfxNHNny0ZUYCGINRbmS6ML8myOl4psDuagbfImB
8EMVZu14Ez0n2+leTq+GFnAgGT28JRJJZ6MmEcJgwgNYCSVS8zw0fqOvGnjitpED
zqWQXVmtc4KGlOIZ8yuISMk2MTK6QpsZnta8ssW7x1u8tKldS98AW4P6cMYAPrhz
inZii3a8s5BwFFsmTDfCax/IMjgoPSEbtPsrokZtCKDvlHTh3vZ+3cAzPioMY/WV
SLe3LZ4ZODXHLgMDrsy0tYAkC6tJ4lB2F+WRlsc4ICooQ+mhUVhvIz2vwaBQR01c
0vQdcYwYrcqS6Vo4a/LikqHIlyZ36/i6YJWUs0DuKUwWmkk0bJpYN43EWNl3BNaR
esRPM/bUt+82hs6ZEOHMSKt6Rs4Zxua2h9jolMnRWJQsTsu+0TVlpuckjtHh0/wX
3hgQ3KCkPHP2yAXkaeyDmfEipfANxvKuI9LnYOxhrfgJcIkz+LyBGr6KzAIHXQRZ
NnUuUQa1l0r9SXHBT+AiDRqgeSb0fOoyMPc4ZOq5sYIli70JLiCmnLvvF87Cc3iJ
xc0V908BbpMKdI6m/5mA8oJtLz7G/x2WIalSwEv1faWx6Y3V2Sr+bWA2N2BNKFPX
J8vtU0RUtByzRxYojG83t6GdN2GAdLqmuC8f9eqyZHDU1D6P3I9imUMvvB9Qfo4R
63896qtz6NSMB+zfuH0w872dE6Pj3y6GtdRrWLeR/62n0XKAjnznDTDznX1JhQHr
BGejK0ramQpa38yYUEgQ1MRsDzwM5wzAtwy+QTjE146bL/1hs/GwlgLTdeinFctb
aanXztIaopGfF1PZtPasUg+N/IFci+hrmr4hkfG7JNvRybFVBS6l6bWXMH9wx9Mh
Z2uhP+IW3PY6dmaEz9OM5aLzhUoSGdULlcIT8OeIoF2dV/R4Sj4DWlw+FrKikRO1
R+2yyCkVYATmtyucLEF3rDnaXBZhIpfPhjSj6VPfEMrTgntvu4LpRo3CmusSDJyX
CS8bvvumjR3z3kSX40yDMBzVNIgcHcCS25JQ3awIfLdYaXJ6vRdaxiNG5UByTSWl
rLMhe2SqazWVYOBTl60HFLfr/gboyagD45/gqqlI1WjIVhy8IxQriEfKvixQV7BP
RcOSTO3MRLRZOZLRB6DjtSsh638KCR3kTCl+Jw6gNAYx6pPrBBeksAP9V9egHb9o
xh6iKaEuz5I+EfRC2GGr2dpvVKgkPoK2ro1qJQZE+pChTy1oEG66u/R3DNtMlMDW
NmEW7tz5DhFgliHVV8VuIIwwbTsT61aigHHF9FnkWyqRRwlhgAnRFBKARfy10SmW
sIZO2QdfMLLHt+yNfyr61KQlFEDn2eX8jaqqXaarK9y7FqPv76rA7DMzhS7kKcn4
KPZrli1X6vo32fd1zOYxJH2KOS5dlHDNHN+r+sHLIEBad5b8l1ykS1/p/nMFzHbz
MTTu8KKUC8HopQOHyFi8NBnx8++9h23RBu1VRpcBUs/2MXpPBv9SuJdeqIKFB8tW
iaa/0VhxlwNrBU/UF85UnxdKQlk96/WCFsRTsWILn0GnXHto6OiFKa13ctmhzCPe
5whH4w+9qVxm3swwHizWFTJrf/jii7LDWoEPWxDNSS1Q4XCmVi1k7Llzibdu/S0j
2Q0wAvFLHoDoAh75jjIgF4d9fc1IlKgeyH/yy+knQgzG8xUuKZ8Z0OHhE0+1txA5
5WTgtajA8HuBHqbbdUAy9v4h7vNJMh5HU6ePOnf2yJoM74BhoDoSxXFemktcYEQr
F4RsNYv3tZnl41ckxsiocPs8XDh+c69KIRuqpILi9mgQ+cYTvZ36F0lZbB1tVvKZ
Lyrv543b5Qkr2rUZ41Ni0N9qPR7gkbGEiqGREg9WSbp3xInvzZOCQmGUfn8I5baB
zMdYmrUStPGjRzPvIyXab1UB3TrkHGTASkXU/js4OZOAwo2ma/P1FTkLmO7xIrLo
E5uFxlUV5eROicuY+1Gh5FpmtwDNacVnQ8wRzDAPMu+f1ZAq60DvbozA+9mFxXYs
yYUOaI3h4IPJzTKA5oqhYu1lxMaEDGIQ4xGFsEhiJgd88mbILHQG9qhAgPkiMAlr
mYiRQcf5OZYFXQDPcveJUxFRUp0f99wXrbTaejvC2+nSZ4+o6mKS/0y3MRgjap4v
VTkA8Hu4xAFYcklItJ2pZnc5dI3yAuOugMP2x8Pu7DN9hqXgs5lM99cRsuPVfhAu
pGaJwedCKIItbsURauyT5oxZg7vUD0fMcneZuGvbiqcgkICHT9UbJJF+nK5KcGHZ
rY0BNCtbD8dghBbFYMK3I571KBrUP1kSHuPs579iinm+Gf+969btDD73honYf7IT
SZdvUPezbT89rlEzg3HtRsptzprul04ltO9yre5x+aksgDbusg+D6NOFywoPACyo
d4CyAHrLm2e+JMSxJsE+VSfaaYvn1JmzxNbb8Olvs14ZC6b0+rSEk14npRM2VFbB
8367hP3GAGn1zv87MdQlgPYv3JKYQZlhATbjXvd63FniGtqSoGjsoETyXRLtTA/t
Ko6Pvgo97vJUBkzQetaAN/+5yscDXlgbELwfag9v67DeetStbYOTrs2JrCsBiIFA
3j6or/HGvyIaVJOT6miZhycxl/2p8/pDpAjAmSUqBgwZlRsDu8/gRsRd5Uj+54+o
QAgoq8CKcMmanmrI6cAcOhlB2GT+kuIKemL4tybyWSvIDe3yn44KdtxaYvJIAsMf
6PUir0AIdZA3AFeprZC4apG3UhFOp44oF+hjsn2oI+oE2Z35a4DdG7KUUZ5mmDyS
jkgQ6jizoxrTCaRx6zKpmx7dGJNZEInlZVqQArEzuMdtw5/VnS3/96e+yBrMWjea
ZcbBFuhNjDrFta+gQZXxoshKQ3QlsTKlnUfVjEdFJb0GOzdGIywD/O39PfPSo9PC
aoKnvtsmkO+k4Dka1gZcoxXvUwIOVUKw2RW79/oqAY+zd6ln5IeErGyzXLSgM5GI
VcBE0ApvlSbNrCROnRdDi9uqLjhaIlMrRb0DLuk2N17tQ5s5Ux6ERqDA6vc4MwpU
gwChnV/0+zrt1byl74M7TMmpudnNrn6PRMJRmjsJvnf7p/5UAiEhHpKuV+0z3z2A
GunSchECLDXzkHnVgPzLxYeyMbHf/O1eP3l2WWsXQgo9DCYDyROytqGGLfdoRpj+
aS//zA/EJpkVpfXWI7n9FGuzohZ1FUxAgw+ErWIplqAnM+go+030ol/Ch62+qcA9
niYdE04pTFx1A6tn+I/nAsZQ+kvpMWHmmXSDjEFb3m7afud+OcgEIqJA5pW5eKrc
jwoMs0+2q47xJoJuppF7ckSNeMgDyKxKkIsW7TKfz+q3gm80wvF3rjMl9jt/DsFq
vKNMFVNeLITK6wM47AV5Hk4VL7XqBYFlw4Ddc2CKYMG3mZm5ygPdYljAsGErwK1/
BSET1ypIpmeJFiy8AjQI5GLOzA6dlb0Gem7fs+uk09Hpi96NyoZdaY4ComvWvlMv
sybkQJq3kvhJHlmDryv/QrUHBT+18WM0Eu7Pv8kl6AGLjBlCHhXMaPOHVVajKw3P
dxWCcfT5h2dmJT1uWWLGOvBz1WcTbre2SdqiGDw2AkD4YU+W19LFhCTALQPjIXXK
cX0y5Jh9xN3RUPFawzylFUGqzG4CUmYULlf/UDxzWTARkO4OUvO5hZrqtEWYfgnm
7ziuLvrnxoDqhYLc2k0Qvvigma5XRmw9422HXm6GSybjjPBVeneobtYe7cVgmtvT
RTj0wia4h+1YDs/JQqFizZIxRHk4s4z/sbOquxtATJVi9ek9XSJ3prXO1hqywJVL
PAwyMa5k20pXXtEIPZXQeecbJWfp/pVhgIbdW+B9CCDNmkFLSOQh+/gNFpBj0n4x
fqOWOV7auFgMPG7FblEtLCj3EBt/homZRdVgfBrzQrNJrt1L3vjdspoENlYXkUm+
HpOYceXIg/XpbpmK0KOUjcYs4i4IfJKJJFo6IujVjFtL7hklSQNKHqC2FcWvhAUU
1DSOuOkpGescJchQMs5C82d7YWirTctJx6W0tFyyzlUSElFT9W01bgqDRj6kHGwf
sCJ69cZ95j7g80vLWy3wkDB43miIktS29kAZjZa+57ROmm2sLjLaN3ffUGPE0L/M
RNjPntommGyucvzoZ45OHrH9DgHP8T3sOKKgCbW7pVzhCnfj2HbJV7XuMCLY+8Ht
iNiZgq4vVDMFr+PPIjxkvDcavqbEhnuM9284TvZHlCAdQliMYYGsyg1rtneXbgGg
zNPSlHFH+Gu9QA/Eo8XAx771m1GkiAH5M/eW+BlrwrPoG9KFo1iGiFjMMGDBVvKJ
/w7Ji+jgMcLPp5SyQzyRJzP2SqRb4GGH8zqBE8qIV706QTs1IrJu5ZdnuF3tkPIB
X4k124c1CnNhCOOToOOQELZWWVzca377qtdtnxd5GEmb1qCGWR9bzAXiEa4ZOywG
UYswrn9CUKIev2JMTjNZK7G0hkFTS3voq/bXtvb5VdBiOGgHy2RAzsYRsJe/iOco
0qoUYwYGRF3fNuGpgxfYH2mwtzLs6ulbGjjgGQZpgBd9nf6fQYewbo+UiSCNCwPP
dWRnbQ8igUVrMF2sD8ZI0xB16Dz5ju3PN0mXXVYR6oNMOxI3OfouGbL94r69Hyu+
2bY2mNUUf11n4vlIcFLEinuPsx0cAPES/5J5FvBtJMRpR2Tex840OVU3mypFPwFK
7JEUXEy94gXCFoeSuigTBAlHvn6h1yhTl+DAerWj8tvX6ARnCi6sDtgxjyfzERG7
hDLdH7Uxv3ILJGvM3ueY1071Nbtm97mu3mShj5b9DvGZyxIjJMzj3vyeYdhpnWpS
NrlDXc0gckU7Dtcy9QcWj7zfyBiihCJivtC4hxxJbCa7Ap+kWYj8OHPt/mS2x5XS
+/Ope0b5ELG4EU9QPLywcKy+7UZaeH0LcyMJHMsJ9ym1rl5kYTVz3mhjziwV/s0i
J8FOsI6amJI5+PbjHweMpN5UKpfUTBzhdUZTSGUJ+NnClOU494R6C0jeslfePdce
oEjBvim+h2FpB8A/RQb8Kl9QBW65Xzmm9jawvLGAxKkqkvIDFb0haBbq45WXCiPX
4OVlTPJtjUQ5kAJFCrgz0AHWVOU1AKDtySG/z9bPlLriS+Qs1xa/4ZRasnlxGqZD
jitObnPx/2BYctrFIPcQn/pPbG8AHDbF1zD8uzC0cIXC81gBUTpWPgdr1UmM35Ap
E/oeCpWlgRPe5dZmsYM6m38EsYDW7sCcDZ3tC0p7jVo2jwftGQsvpjhW6KmORtjE
qs6AHm76hn+tdy+d+TWsaHgGxIUYxn7D8RVp5+39ulP90a3PIFni84/XlxpjEuEs
OJaLWCT/r27as5KNxDxRq9nCLphHOt09EkWacxPCVcjplv/CEAVT6PH/WHLq+7HI
GPDE8xx9kDq8j59eQh9M0PYs0k+2BFaWlsE4HWroID4Irnv22HLx1ap+8yC5HY9Z
GLkfFoyfnjVCiME/JRnqjl0n6gHgcytGMRiXhMGsymYo9MNTY+iUYoiZSszzWa6p
Pbsgq536FkUocKwQgiEchhL3IiQxbpfyoocMjrsXkNujUPi10HZ4wD6lBBYW7n6B
jmO1vnHKUEL21WvEZ/OP/Icd8K28tMrv96eDuF9finUfXryTtM5ou+GHF3tNAV3H
bTSw5YTeCfF7J/TIFkjuNIHINS09QAD0ndHc6jLHJEkqQPlAFanahfbQenyfaXwA
Cr/99NAnwL4ulpybxd6rc++d197mH3/NRiC5nozOQ64bsxRolYkOBLkBp6nv2V2V
XZIEtFK4xSO+2lXmF2q0uyfpbmIiFomuRr4vVvBLllqfo8blIWNdYCF3HS4RD6pz
7r2QjLhsIk5mJ7AfQwp8euHn9hiuINKDHXifOlX85Es6uHTlSXK9L4SQc6hxbRQb
iQ69l8el1whpO1m41FvqBLcUIzutQ4RiO8FgvlUT+qz4ZA84+DX+VXlHNA+EDxk7
mcIl5gqRWxcYTK8j+3tIy6sLN1WdCkcKXpxpMcYS8iOPwuHuNRLsQtVkQPeCxuHt
0bX6Gpdt78MWv2Bzr4d57kFcEJvU2UkLuBcRMjP5f4hwm6Yao5glOYJ/rJ5MVUIr
6ue4Gkorqi0f5rUHAhYjTgLrAM1v1Hlyf9UxYHRB3NheR1Stt5XmEVWsd2RI6BJF
tudnp8uMjQy8C4RbZnBGb5HdSi0r/FmX45FJCZaHh7jJfcEXM2VuHqfTGxRk7YT6
AoFW5X6gIPKEXlEZkJz/qmgQYiPhgYbF40iyqlqrRhM/lDOXatNxhqZNWpmErJxC
Xpjr/8IvgTFi2njyv4lQmVPaYHwi2RQrB4Z3h6zXdhyB+3ybT/sOw/0uamMubbup
jZYBLaeaQbhi6aCfXx/4etxxiPURIQOOhkAi8bH2YC1k3Zn4GOqDCNbACbhU+j33
TNdV3leZQyQ2rvl9qP8TpIyNsZ7/d/lktBq6pCOdTPVMI6a1m3QXzdrm1oT9mpuc
aO/hAkFSS6ATN7RdNCxeB0/uJeVRPYqxnUIDQttGM7dIO5GlouRlRdx0WAFumvdW
ENJL3eGOmTdQVTaojwLjp73DvkL5tNPKV7Zw252NRUZ7/LQHXg/wnAoaRi68h6oT
7Vn2dJcWFbX49lrpL2l6h/UVA3PH4S+ZGZ2dQFWlL/qV7LKlnrK3rxbF/Oq6jqLl
mKVIrlf2wq72ZxH02OgQ2HS7uNkldfKm8hIXTWs2iIGUYhz+fZEa8500bhErfWoo
wOESRaAKK9fNPSYXZC2ZEeg6keAiip95fusc/QU6nebU92z+/wHu7n1tNPrv4cFB
BrdvTV20vKEcweF+nHwd6h5BKqOS/jhtbWwVTRv4194tPenVrNP6JXKYcuBT6hCb
4MwX5UJmbIdxGGy9FY60bpMHDeyTevz0hzEumuFayO9+GnsAi8jP2zMCG88nnXBA
/4Ph5OtO/JwUAnMZu+j7OL0+WbmsZObfEg48sX+7MkuL7Gso3nm7CIu2koQfD6If
zrRykanuaGSGlVWM7l9MZ0KaRqleGqxsaIWxGeda5G1eWorzHLnpDHeArJCDEvZb
UfxYy3p0WaHnXOr+hdfXza7DUZU6JYgGRCR6MkQAS6dFa5rawk3CV3MWWhEdlXvb
dCyXpOysKQjlIFdYL9NeuNbRXb6jMVE8crWzwIk/GsnE7i7Tj+Jp8eAKAPEmclPa
JR3rjDipDimnNK90CFdxfJzhG/zUJMK3Qy3hq/FqI9Px5EJMBAZDpjQHnspThdSp
2MLdqu76kcancS9AKoCZtwurUuxbGa3xPvLqoQJgu/SOSp4ZZW98rQhgYw8toNZ+
JaLGViWCrU14SF0GCFtTU9bt09CUqC/7GYKfRVhGe4iz+of+9k3LJXI7aFtejTjd
dmeTKawGSj74no/vmBbclKYugX8trW/3cKchWfYeg15h4K3E+4CfvJzcymy/54eQ
Ss9n3yShAG6mgWRhB12eBjyIDrr3wiFp9KN5lzBBHeusrGrWeByljCR+B+C0xQRN
PQ6buguBTvBgUrczAXKc4PY0aJChHfcb9M+qgrHoMtcOAu0iw8XPPVr0W4BwCXQx
f3S83ZELD0gZ9f/oMaperIQsMLMHdbfBl/SS29a4hRU9ffoIWxU6i7aDBO4hi12X
TOR9T9M7tz+CaC62d7smRBGRWrrt2sRo5U6jIc14SfL+5pl0rFQt1Zp7gdLFnHDU
CDDNNx1LNsJ9IrcqjUDVdssrK++A6Amjmphc4lfR/uYC01IEP0YjcmevVISSM+k9
Qi8izRaw1HfORvlry5HdBWW9QQ8tEiaG5vc1oIeUyYb6Q37yii+8MNWvV4OuYDOa
Yj5sSKjeBl2iGrYatw8p+54siSdm3CBgl31KzXt5pPylVAjTyDa13LdUMiY2kRKx
he3Quoh4pnDh+iuP3OgJZg==
`pragma protect end_protected
