// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
L7JLiczspFSoUMxqYyCbrAE5m7a15FIHK5hizo3zVlX3RPdi4IaZ8h55UJMhaQaE2r5B1732LARo
+WPxDW9xYOGNa78lWj23Z1ubu9JF43KjRXDTAw3qoBgNP7+KXklo0gpaqi+hQs1BGzFjL8t4fEh4
uf+OYjbPoZI4seSmlXnQ4ek+y+cLLCVCjlup6v9zsQXokA4kLWcQj+81qqiHvnRYzB7KAH9P6OJs
VV7nYpyJUz/TrM4yUD9smZPnEpz+TVVS+tpVFMnVF1B8dnO2/7gBXGNJG85Bf8jp003SMibmVyy6
taZls2OWiywPnTIOsVip19oT5pyktUJQSa04+Q==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
PGF6fgxvrCH6GfUDrRhVnF40E4OrzjjCBOvvJEKdrH/uxzLyu6oaAAh/95GUg4u5hqZ9bHyOLNXN
FYuLc7cZIHJwBHyzizXQhoae8grPLqvYMbZL5NkCUrYfcP8IiVEzPYqSk+w8OCiiG8peZfnfoAv7
LGd5Ks5mv3lf7TYDiTTHQxTdh86fQaYucfaJfNOM6yMy07Mhu5km5BxC4ylge0jOYSnZgsW7sMSb
r2mOcuLQM581OWqEmbsDNmsacIQ82FYPFnaKldoecoW88+WF4z8YvSqnlK2nFYhwuuzFHMQ2HaYj
og/P1KyyUM846T/G7HJBUXM0BxZ4hCyHxrVot2kbQL9e6s4+TRlhM8ljnRO1bAnfco+AUKcFLR6V
f53Eu04MGOqsdNX5JHR/hLhKbs0Exwf8295em+RSMTYKF72OrQkwNaVGkGcJ8a7tdMWCD42/CfWx
T4FJTi286AREN+ez3nJd0Yl1jmxbnneXebrCC5+xzrZZ7pizjFEAeCFKlnzY3MO+OVRtYAvSxmpC
7I5H10TS9xzaLCdkLx9M6uTK4h7hYlnAR4ieQMUBgMLC6HuqlNPCjwSVLxP7pHdvl7HeSkUvq5Hx
fCmGq003wZaachrHsSbt8kCupHnHGGg0XUtta37Bi2qghAcZfTlYZNxGGI8Mr9GQZRGhU5kuPKB+
5vIADmrDKp1SCzjWJOF9kJ/TMBMUTTg8opcdNLY5EtFH+U0T9AxjRtTkfrjcfU0mjX2hlZkZXL+A
u5a5/dyn/lcnsBHeaCG1si1tLUezGEc1W/A6GN2dzoYBEqvzHzmI0n4f6/heUJZDkCshOwHKq74U
3l8Um4KlOjsNxsx/Tn9KX4vu+pvU/+LolURaplRb/+GSoEVpFr+OnDuFGHisKzY6tdBWprrgZ3n8
W0jYjY91VkURc9T56mOn0xBUrnoCUP9A7a7uD4TP0VBjejzrKcu9g3gHv3WWFachtq/XbVvuJAAO
hCwMu3HZQSEv6XfxQjKLResD7Ipfv4RvnHdkQLjvzCOV0Dkg2gJYnmIlSsDr5kxunt/oyqnak6J9
3/LZGM674fHnHXn2T9/fvliQ+aKocAKGOQglfEs46X9wvRJD7m/s7U+9UHY7xeirzg3K1lv8KMrF
G+oj0YNNM2FK5hNdyL5A8syR4KRpVyYn9nzIFRZvbNcNDfLbdxvuAa8ajREQh0rHs0BNt2DEFIyB
TXJgDf0SHOrOhNMPXQNBfdkadULDVGK0ptpq3zwCwm33cSX34M1sVVJ47HsSefrN/JQECs2mOL7J
U2zn2TaAvqgj5ZhYOhL6OZ7sx7DGM3xZ2F1TPy5T8pHfoRs9MQftB4Bd3vhD9ax1jAjRPfTAvMUu
q93EjwdwHOD9xFGxrimDIVPPlG1kDTHMOGX2A/lo4Rhev5TgahGNajUcsGpmzoUE2Z7X0glRidT3
jR81v2RJWC2xVB96oCFNm6JAfn7h5Z4yzjPylQs3kwTvQREeE00NHUadNREdJIu17hQCnxCZPkWJ
9MkzstqlR/RvGiS2XuJlIFgzNr8oxdf3EokGX7E8YH48W9+rxNGrjVfwg8ptCzn8zs6/EguHi3Sg
V9SFgILmygoOLlzrnneUKPjhJjAoHDS0R6RIbyWiEuaTyNDqdNfBgq1p2e6BBvGF2T7AMF0LoYtb
dacL9AyTYfAdRevX36rLVdCd0ajxOYDDWLtQqryp/Q6ZXJG7wGTYMV0Gxpog4xZx6aRQiofpicrR
OtY4R2etDSOoAcVHTlNDEWP/6l73JuK3I2TzPTUlEDLbaPxTO/u5b3ENpyblVwJRdBwqYpyyNSbY
tUCcHl/foq0JCkoXy1qcCTqk0UsrBhmYEiSukV4bhWuqN/y89rea25b3jhTb2iBdExR88btRRGXn
QjDxmltOYhbkKk7x5gz8ImmZLjuowkqnjgFtarGXVh24bLCRw8OytRoTf22W9iBDAWioKeU6wmy0
ZsrO4oj4ovZuNrNCVDQwocICsRWpTW4tDjJhRVMXyr7JYhcPjjvQN6nUHUvOOnY8HDs5GOUNwthn
+lWhxJ2v79DEOk62hnzT8FbjzKHXUJ/eVPE4yPZDowhIT1ZnCUUoeQYihPTRt1Mg22/CKW8DawdS
WU0ursZ7hPWN720+EKgxz40ztpzBySW/Gs3eBlF0PuAh2ieFidd7FuhvP6WDlWLl25B2xtWS/Tzv
vycPVCl1wmQEm1fYleI8tG3/mtlyW+ylYneSbmMVqv9KcfIWgNIVphXUIrJ42R2CVwXvtIb5hIXD
5k8EjDXH0MT3HncQz10cR7h7SgQuD6V0mt1DYX+BD34dbj972rP1Gi1eNbnMuvf/lEIYiwzY9EX/
XQJRmKmge6dRL1X9o5x7qyKFU8PMkCHPXBPVAtv0AOfu88fFpcjWgA/2dkXftIfvGFNmqOI5gs59
Cei/okz6BPC290+zxg1BAvGdAPt/0hASJ/kfqN9E9K1jMQJEeapLwhB6diOcm8FScd5039N+PjaJ
AcEqw7aEDgavfcwLsvji/fYOo+nWeTj5HORZ0S3u+i6ZGoI458tSg0JkUMRGN9nfJQfw4ULULjVJ
6bJbOgRUzlXP4s9ReEVHc9V1xAWYJfQr0jFTJ0PVaVStu31viTMWgH2PxdTjuNsHQiOB6AEkmllA
zvBd8by0ji1TJbmPqvpZP2sMkYqJpb8RplXX4daC+70Uj1wxKyAv7g2AjEE+iUipon5MZjiOV6aS
lWF1IfXVO5LRuxsA4Kj+7MDPPq7U4b11QwaIVLf1u7TJgEBrdHqd3Dc6Mqnoc9AsKfxTIf8k6eSo
Fq/rNpZGgf5q8dgxGBqfgUSPKjARVNMQb3JmT4Q6eXOasso5nq/IGA+j8mmJG3o5APwVTklT/scr
CuXpyeZidID+VaVpWqZs9Fs5svHxdslOjN8vgDcjq8LbSwonkPm3ohV8QjsjIwxx0vX2TYFp/9zq
Fb5VgrDPI2vZQPWdQY5fCkoMFqgtwZ8HUCEzQPT7b0SL9HNc0Mq6nz83nz8stNSXeMhqtZLOvd8A
DnV7hLmvyG4X9TdWS/Z88K7Rw24IgCI0O/wOwATSTFdSe0QofKLl5zo+GUpDK4jifeZ1WfhF4FM9
0W8LV9bVcrVHBoU4v1J275ok3HUuaxpxsihOhe8b005VyBHll5KAmEEDe0YbMwTrMtQ2youcchdn
hlz7IuIPy0VHYEJKW2HSvCsXstczxqr26l96FplAY3YJEqMkg1AglKgzMDdWi5UTEi0S9+iNFZFH
uxTF9169RAApIj7KvMUAItaF8RssSWJJy9xubQpCPh7KfCEgf3R4Ylq9W8Zj30fPHlGOCbhT0QNj
BzCZ0O0Wx7Ek+rM1S5ROQCBuzu5x8PxUA1P127j+Gi5PyeLHHqsHPS6nw8+KaQU/TAxM7S+HZpxx
sCR7hSNTrKQol4DgaZq6tDJtD05rJ4ihan2sIKiONm2Ur9YIb7aciYzEWqI7JOLPyBHqbdypNCgo
DGjF2fh4HnFPAMWZPOo0VKCSMAqsfot2h2IY2Xwd051Zx+drRNUCNRbHKxGpeWBOipOD2eRi4NCy
sG0GT2CT4g3URqJmyv4wUmC3yU3ESYVdvFOW5kpRZDt9fzEMppHNPgaHFzwC4/F8prLti5rWTGAj
OPDNdGKeu+jKK8+L5QCHZJCIXAxs0jRqIeQH7+S3vIW/z+nZB7sLOoVgBw8HmQfhQURpSf2Nryke
aw8FWSQIH1fF8WXKVENvcyw2Tg09j1PeofjyBxXzBjCxumNjF5YeSF0GRwk4R7ariDU7Icq6XwMo
GLXaxUmVjAi2CZUeorD9YvtjAmYSwDd83zoLP1aOdiwdYMbj9AA9kva96dqi8jJMDIu+IFD1E/q/
LP0IZwTh35j/Mb80t+pKGJaQLKkMVewBXJaICUW2HKsJ3uHcc1C55C9FMUbKnns2BiWPAKZVb+F7
zl04ZvkgohvYXSneY7vQcjesJIloQzorAU51+ZUsVFPVSfYIJ3c/ge4T3y4cyS2W1CQdPTezervU
YVHlsbCTGKvRMxSb/5G3XG+xkZU8nSrK/x/C2/ELDNxa+tQVspxDj1wfSjgCjzkK4obEGM+f/hjh
Q6ad2G9tOMM4Mt6ta2d13kYFgm+lopbEcQn63cA23BJwbETcXMziKvDGWzvhoITSgkORXooawURv
dAgscG+CX8a+3i4yRmAsnXenccOTAtrF4GMlmufaTVupR4lJmMVG1+Qrj6SkhDJp0/y2Q37bSVSi
8lanbpcUGEvqC23pw++9kzc/FRgPN1UBiYcQkf5EcbQrHXG15URySCrU9B6/6djxO+NN4wa8syOA
G/lwJe4hw0wo1eIPXIC+DASqv5l12cfwu0fZpNCaEQamk9MpbKI8rMpFztESW653nWYqZpx9e+YE
0HxFBGwI9YzPk3C4ITU597iu5t7Y+9uHTT944W45Kn2T5RV0iqUuSVccJglopJ0Z1+XpJ25KT6+Z
6oWVoc2VsRm/T5wo+iPJoJU2YJoMGCxfV5YFwz2iUp1znt9oG32rGwMzeLWkxv46Jh5ZJd9GrZ03
/eg5AFCLLPrtL0UaewHaLa4ykE54U6XhaKTY/7eEHuufhv2j5HbjLXgjNoYOND2nMELpru435fbt
R97gPNk2bs6JKlhAkLrvc5GgurB8BG5xJ5a9h5d38jf4YV6rXJg8KF5Aeiy8BPJfKNUd690D6cW2
CFhHv6H/jS8W1vVZ0txICJoAOk0O5zP1rdeytUoWKhWcDecZbdXwHFdwfoaF/cZgsUXVG3quQ4sd
+Z055142NUYbo4J45V5I0EM/o3+Fe7keC9TZ3d5z4tEBAWfg2CchZh2VvDJJKx6Xaq7rgkDLkH2g
NPrDfzYy6O2pkpVjaJefFOlp+Z5KSdaB1ITY8na3eF5y9wtxjlFEV9OU8+7hKh++PIIB6zqgrdy2
kQV0nf4SD0XkVaTY3DWvQHCVs1sLoKnMPdB3gNbic2MKP1PVYNGXPMCQsP5i9yNxZ9JabMVOULAv
1b5GEJsaA0gz097DsdjHhrUj5EGRfHSYN2xPsVrIi8Y5dLw0jY8jAAVFw8yhjHN40/2069Fzyzyj
iShAIZH9aThkWM6nIq47XDsDZAHVARIx1CoUXZ90LKMTq/kiTF3iYO3zEv3lyVT4R0PIJJAf+9UH
WmeAhGYvqc6m3R9F/XExZOGmfTW9hvkE9pgR/HeIsEFhIYrtVp6nATswkW7g86voOe5LyQaVVmpS
5tTygLiIp21IhCRUiUzLG+WE/xD6yR/pFaogs3281AQRbicxlS7c3UQaYGI8MbKrq4066o4zah4w
zTTMfI6GK2555G1H5v0fui4lDqFE3uwXdA5+d3D4yvnaSzUZi6MgZCuV73Fe+oIvTBfPgif+WxkS
wYLjWLZ7X0nx7dvOhLmBodwm6UtM5yuwuFvOH1WyGoGeHvngySE5/3jOdodoKtIxZjbZUGBDd1vH
SugLiliGNd+hzaPf+XCY9MJXXKtvbFNJdcD9FIdkZzPnWBFHyLacBA2m18LtsewETWlnjfkyYCQc
iTLjrRZUcau5qv3WLaFtlzvA6h/sQLMcwtPu1NeSdNXPT+sv+osxhkz6NuQDTYfIfMacxLf1Eno6
JwNU3jRkqPKpPDruLCD9uUkBqryZPx+/h8NmzLqE3cNzTlBmy74ISdMbwbaTfNq8HiEInhWvCX6J
AVLrb9IcYtjHwjJBxnDlQrjRg2Fk0Rl7d2pV20nNgGSOrd4Eecz6ycQjIOqusS3LqjE4o1DNKjfn
LSJasx2bdoQe68uaJEUqvLnC08rvvuGEtqzqI+0MPU0mZ6wFeam0QHLhNGqcgdrNMLUHWeDRW9dF
ONVIbMW7TG+2d4L1i0GuhHlKF7l+nEwNl9nTU3tdkqa9V3nZoiIYDOkXv3I05hUlApZoMtN40qC5
SkoMilxJ2NTwDsWucRK7JTt7bkf0OVx6fUssNv7xwHMG7vlCbKS5//ZLVcl25uGdvQvMS6MpW4/b
DaIvYmIxIDx75GOQ76+dYLjd5MHmRiEo8VvHFALHW4wJN6emrpT6fwgxgZva6QoOz1aQ0c67qsvb
BAJprvCxzo9yarHYPPwdQIkIowPgRdkojTVLNwG65f+euYdnk+PF/BWNgx8TL+8Dw4i4WajksjVY
xom2O1HXVCpbncA+fGKKaHKWdOh0S0QziasS0IQFS1f9tV6OYYKRA6diHLQvQUm3cBtZrgRpdatF
0tcG95QlKmgNkideF0dQRprBkxkaZlqdyb8ye/TqTKJyJCuQmPJwGCyoU1vpco/L4s5lrzbirAIY
bPNkc6yEeE4WLKO8nN+EFSsz9pwZMaGKy5WGFMMgmgsA7Y10+IXa3s6Xt9raP72ptffnZmYq2pvS
7M5KQxg5IAIJeN4FlWciPM8D4BZW51XzAemwkAsfbBvZVcEYkAHGpy5guMSqKOvPX7TVGjYnkKGh
iPC41nT6fws+qGNp+Nzq/xFEuzr0Hc5CqBSMsseVQSH2GDq6hbnYQv5nKi2xhqNArtCDD0TfMARZ
jl7L5zgMdN9+24wxzR0+eXh3GC5vd/TTKMX7jL2PuGsOijsLfvwoeznYzOz/WPjWsOmcykmjfuWk
9p54i8AT/pybPZlRXp7sUWk6doBoPtbXBRsESpNSrYl8eXSOveTnActb//TCM0oG7XE+3sF7rf80
/pZat2oKARfH2PBa58Se8SG1BpRzTeMzG76Cwh/ZCy0tEWz/omFKIGCC3gDCo+HUJaacAc2rmMRQ
3ELU0ktP9TFpzbBR7y/soFlpCvV8KP5lo6XyoeQKqwPuVzCsf76tOeR2EPi3Ma3r3IZN73Rzk/Vr
2bTLkMVZg53Qeps+PiujLtJt4OYzmkO30ySopUGzQZ2ZnI9ZmoE9W7qt71wZ4LTAu0tUdw9D6KAX
qLyZ8y9kV4ErWaOJE1iibLorTEMloZnNIWmg448LBWO9SatJiTWG2P++jyX9lhacg2GPd6Vmbrpe
4c83htvGGIRrbJng8iPpU7wtFeDxW+d3VFe5S2WH+CBSStI4DFU71JKscgpr0XpNWfzNOEcqFSqG
VGnbcp0dZk6g3e6P+VNZ6IFx8wJlHYtqrKxbyWbmIr1YXoQFFZCX+tZ/SgW+9krrRgbA4DWgqoao
G6ssYBKWsycBscK6SmYIMVUTYoF3u+vyxhwOjn4lpfCU2dr/mWHlgph6lRUztwXImmhi7WUheQPF
fIqRgs+VqPPZZcOgrrKVS5aHsEKaqkRKJxhz8hNZKAlCXhKBTfOF7AWCDF5re4uKZtPkePXHTkwh
Im6MX8fJMZ1HLb8i7igCGAS8vsrODbmm3h9Jdz03HFUNH7tg0lHybcA2INGqdjHDXc/u9j/ACfLB
A8h0g/YPl+GaGPseNLkkWw0u5xtdkY1na3jnVNCofQOQCdYJ4uSp4sjUsWy68JJ+qRsXqLY458Ff
wpwFwXiGYNi0USCb8/VjnCtl5UJsRJJyFAiZOmBV4JqNKcixuayTr7+zFOFQQBDJX29TS6NNT45B
KsqbrDqvMQKoaHonIff4JiWqxlxbZCNcz/4IepqV5lLmkco3c+Rvslpw66ywnsCX+irXfR8VBgBH
6Yu9/oeeTiindYFxsF/bEMd8WgahHjeOhtNqGQ2OIgM0j0DFcR8eWPsz9A5WqeEmA8x4PXCZK0im
k9z6nNNiI59ocHU0uAa3i3Bb4p2xFsY+URPybrsuLh09GpJzWZVIPKZz6VtbPlIvIXF3qxfNniDj
OKxo4vWrRkxQA7a6dG9CaCyZkPY5fV18Fcg3xaZt/TnF7qq088KYlE9jEGkOubaZ/GYQgGLJck/c
ryEWLi87h7Ci8Ggu8wv+UlXy4wJiwhBY3/Bfz9zGDPwWjuKjXp0/jfFR498Z/v5ecW0tWxISun45
b6UxiCcoRQA5H3RZobhyphmfq5JtYEFOyflzKgg2ZnkMd9mZg/PI+D7+q1dwO+oz+JhMo2HU9yQW
Vit4ivNKeJBre8OgVn8C025B1OPpwKWSZ4pXRHNlJhudUTI4699uzIKhEWTqYIpF7f0sRrw+9Qk5
oh57hrPc4fRE2VxesZ2FumIjpuA8dr3kyw1MNTZD7tUJvDbYiDJe0Vt3uqVp+wYtmv1xj5m86FOR
3Z/EfzpzomTMZ/h8h7QPhdoGM5stRBH/6EgGCDmLC0oasIlU+WanscnizKdNQsHV1wdv/DOmihto
9wjkw4zFUD4FMNaxFOfVec291oa94nTlFGjx9DzHXnxAfkt/i3e8nhsoflDNZTFklg6zgJ6n/Rmx
sSJSOGdVqIqaSVJYdxFRw8xh6lx+LryCciDLiZ7P4VER3y2M3mNGzXyanG41FXQ3mypQhNfvHUIy
Eonepci0G9yRmE0BS5dHUvB/5tVDjmCOpmTjoIdSG/1ZZkv5mQdxPWiuu/hNkIqmq9TKA4dBz2Na
mhQyigSLHDB1XsQUtjT63G+x90VsQsGbvsX4Um93jGKk/tg9vllf0hMy4Jejyx+s+KFCmuA59817
97K2VhzOZmr9O72XtEJeH62R6GQCAqTtSbKxriusYe7/9sd5zbicOF3fzq5AB4U48zY23y+vO8UE
rhEPUXrphAKqWw/Jd4PCtO55em7Jbd+pFQAS9h0N9J3bfxG1ZZWiS5silJPHmFq0wIfn9DhIv1Ry
yue5FnJvWKhLpMMRo8BuHQ/UEdFmU5xBvl9HMoEtZpRA27JUjqyikZtTNqj0Csd9eLIM7pm6IDn7
LPi4xopFlIz6dN8rlON8e2T2Et61G+FnZN+klkCMH9NdDgEt4UDVEb2mg9E4BScUz/dtKtQjnxV1
c4kgqsNMZ2a24ljDa+tntlrNOAw8m7hZCTk0HOwVC+tv4DcFrnxRcMf2urF5YoMr9LJLePahvgB/
1HIMBs2YIERAW8gT6uM+29HEM5/pXqcU/v798t7u6Xo64ajaVjc0oCcXkQs7sQ2+E2CLomRTpd2e
wDzDafizEonejiXdh+fnVTK00HKIiAh67XqKtVqYS7/nMjLQzGxXW+ZAywI4/0TUglFExcDo+r7j
ScwAdG/BknrZ5XKM2XbHGbEGaddU4iu6RXrjKSEDwcIDP4L9lwkEoSnlsYtnh5kE6/mgUmOltPb9
Axhj3pU3Khgqnk/ZWFSh1oTnmSa52EW74oBK+jflADBmUBKUk8SEVjWpgHt/A+MWkT6MjSlBSe6A
yBEHtFAHUA9zldSQunQmUjAdUGPvkKDf2TK0yhgTgVm8C3uyUoMStfmtkZ0kqHBipMEpzn49ZJB0
Xi7XG7OeQqNccQ2fjhjH5qjwho1O9WTEWDRzPVUyR9nPI004/EPYYCI4PkWbRriZmyzECs8tK5p+
fAxLewMPqLXDfuCRpdFkUmcM6qeTjK95/k/jIu47WhsiJJh1tc1dfejPYBmUMenz3xd9f+h63dIW
3R1uRSpvShB4cIcJwbwQnhanZOEaQxTaTTlhgQfAmkpqkjqpw79PPNSLHCYm8smiXLTQR18LT/mf
qv8qa0dMiJ3bpnpyjnDSjoFxieq2WsJlkJkNGhv0xHgtB7hk6wV+dlqZdNyOucl3Y+2qdy3l4UtY
FmTGmLTvkkkK8RrtLakRFRAQawSalaVehEuE504IZzAluZeS9AlzNVW5A9UExWwiBuP+1c8zWf1t
cOXGcPn+9u+j2KDMbfw1+9F9ppeo2KYrli7t3FmI9MJMFUwrQRaR0cqK29HNQBcazcFCwYQNMMhF
r7sinASzi4bCsnHLZNDHwE1H6Ht8qm4LP5+Zg/5pvp4AEoYYNXMyTMoELIelBXtg0eQW9/4LI9As
9Kty2krW217sjDS1nbXJkPsdHz7EjpsAFsbJXpYENksZM45LsCZ6gOSJNxCWzV1lhq159JaFZzbN
iJPLlQOnLgQ5zXACh36v3YJwi+3xrhYAA+XvuTBokRPFB9Ov+eAEDcicSoDP9gXt3Qo6bzBoPpCl
o6wAN3GWPMymEX/ScrQIUH4ivXkVzDFtGKiafBVrckJtXI3t0woDs07lN7YkPrPjliB6HrjkB+fc
mCKXk91NL6P+tRGIiNSu9dizvoc0WU6+hFbZBQVgZID1OU80/BYkjmbXJs3lJ81Cpaebd1LxP7cl
OlYs5+r0SPwllb50WD0yI1pTsvJx7wOt5dTE1+QRWQ8dmgqTLJn8+J0uftxUPJBCBriV4e/Sa1vN
RWL1g49XHK9PbhqfuwAYa/4GVeFhkvduFPXUHhQO9velsdj2j9en+1PQkKxaq/CcgEt9/XQD3IkV
f+LuO1n3VmMHviqZKjb4Ygx3187p3cBqb8rm/7pLVKYydWo3kuOq3rLv0mtmrPmOMXZRc3N0hM1m
SXfALfWoJVB6aoBdnh0w2f1aBcnDG42xhLUoM/acvGaeaw9iqcZByIdsiHgNvTce0pjlEEFM5pvO
ppx3jlfBnVyP0V6xlDtvODjk2MhtjnRf77+mERNqb1C1WMx0Ub+aSWcLYjKaDqRbw+9GoxUupXiH
aJSyyXu1DTEaH0CU7lR9mdhsRugZLaUKZcjmlZ8bEtTatLv0pBWU4rPZZ+6XGHpW5u2QyQNRB0wd
z5f7PaYSxuC8sEz4YUWj8Np9kMP2yyLfVtLkacwXBjXcw/S4qHmZIcnVhDjQv4PVZZCNHi0wu9Iq
ZMin3gAi/SQrYB5aR+qylFldXI42Wah7QD1KZYIMN41mFQ0elhO/uvAFAEJC2mrqznULAKTlsO+9
fYsSM6GTXqOHw2VRu7K7Ss+vx5WVlbKXkxqX+ciug9p+S90fQ7tjAoJ/0UcQllnIQqF9Dc0ReggX
RwJZdxQDnoCZJrWadgkbBL0I4VAl2XYb1ByJCEkTTKJ3C3c8zlVVNsNilQPf/FZwzk++6zGHe9gi
Ij7J5FvC1AwFsP45aNuMBzsejqnyxqmaGZQwpSzg+vqEch/24pi3bEdyGCH2ztP66Fn6buHPebWo
KrbB/66OKXnjsrVae8HWq5fSzeiWgJNNfLLE4jGNTxTs76xIFGft7AptW5+6COzSbtPVDbDlV4EO
FoGZf5Zl21KzIuPQCH+4B1Bft6997rYGCkzF/QjnE68ICnL5XR/T5v4o8RxGk+BfkbWtLg7Eb1N0
tMjaYm8jpgslNLDizxGhGxcwNnDDhgcyjeHfZWVR6Lwy5qpdyBdrKZ8BgK9f4XLrnvs6fkPdWK4X
08+vGnraf7tZo2rkZeu/c2E9+rd7PUgmKZ7zkyMzkbInvFwbomVCvOsOYx+hBWR1HUCxg9Dxrhaq
AfYhreY5NFyQE1984j6zZ3JpVDIC64KnXr9M3P7+Vzpy/GRSl5BaSUexlN89D92M3SuNJKC+9bEC
QpRykA+FKZLSo+HiZ6v8dkhb8pSm07Dxakqg/AtyHTAuC9+xwGPGQm3sC7ij2sbMJ8KKSIMEgq0Y
zlOor0bS0SGLeWAmwE9aNKjLxb4SMdBfOI9g4sThcjhgxcjBcoWw3IMfTZTJIa8vFeSWy3akDOMS
qaLwNXQU4sbMKOcIy40I2VZRP2iPARcriRpOFy4LAuOdPsRKF1O/uw98Kia6Lulk3ZpeGmjtJxiQ
iLnqmTlmy+ULIXbt63B6fwxQPWJZgej6E3XYW9w6Vce975uyIdWN07s7RMz/KPzuvnFxMp6l0TAT
eotpIi/5cW7/vc12pWlsk+DSikXaWAi+8flhKcyS0+pfQXvRuoVCMWEL0XJ6Tps9ZIOqJsIWDVqn
DkVmMPsHLNma6uQpU+Fa4F6Ulnw6KOkiag4IEa8fQ6AnlQfQuCXUstLmwA09PUg6HvYd/3xCzuge
/bbFyavjATvspuhxjaJor/Z++4+5yy7D8sJrOauCDYE7JbiGmZJKrFrrTuiR9QyBKetFwsNBioDF
TtqcdCfgKOKFhEw3lTy24uyc1IRuOAR7+hWydp9hL0JIVehT9E1hwr50cuJzZVXakbkeyqbUahYy
Hef1YtljZ+K7vNog3hzkxzpCzNhDcDlJIxZgnb7ILoAkQLhHqIbdCxADoZ/GDOhC5p+jlGOMuWh4
xv53IygkE9Rx8SJAO5w5MqbpzlV3uYptGU0l7bJxkwg+ErnrejUnCQ0cydFDmpDmbrV8VDnMhfla
BAASsJquru+1SkrTkbhdJLuZmIzK8S7PCFm7izGQspZ8teE0cX39ITq6Bc6On0izxn3yIQTbQ3sM
y+CsS1eoyr2RRVU2E9sk0xLItb3Zw4Aoz1DtDlUb6f9iVsC1Tov81Iev1kB/Ca3Uc/rlGo5hJRN6
2ey+y1Vs+FWeFK+9BhODogseP2YAWjfaIjH0kKuf0mATz8ej4DmIlLBU3CihFVqAEUKGTSMO/Y5f
5Kqxkm0DPIphPNtGfuwAw25XcHLm/uoQIJ6LshdPPWa0+lv1c/04HEGn1RjKddUoArV7bU+4OHqG
k44qjtu8lmbJp0iELRUVgjRfwrOW7J8AsUr3xStfUueYHmS3aBgztZovelQJqmVQ9wiJ5eXtroxd
xP9AmsSL52sD5X6sl6vsqumdrIFxDnfI72KD3GHZeDyT1YA00fdFIbu4LatIS6jNB9KZXj6R/HR2
OiF25DZgCwKCgR1AX+wWcNFLa/PltmzH2lvM2Ui0TD/wAUbXtz4cRUgm4xOPTNQ5Gs85EvwE8ZIz
gFgIv1Zy+uDNoSgQc2mcWE77QBmb+uIEH5JsD4E7BCgV7vr+CAlaIggR6QGa1EVwsQiIYMZ94zp6
yvJYsnXN0hSpYuU7LjPUORjEcPCzK678I9K0Ay0WI3AlUtAhmAsS8ONf6hMqUl68SsMC5PkBJohq
3fC5QvjwKkEyVA7jSXSxTxsNuhpbx9HMjyDQnuVS+ZTo+PbpAH99lE91IoZPI78JDKp3PoQhu3cw
hWw7i7av79eSaUUcMj/qeVEVh6ciT6S/cGrMTlBlmahKPSh2U/2xeKEkvblELhbdKve8ivx5tiMm
NR9Wemhfjv4zthEWDlxl9hU8XslI8sXvZf9F3HfsR5LrJMfBXS4bIBl33+rcmMOHweoPWMz3WPE8
YXlF7VLJ7m1JeADK0dlSe/ScoLN+8IIJyrPfEYFuMmvHo/qibftmeS0C8UXjZzNWBCkGM9hOfgAi
YugRhV8pPwEgo9fFTCgOhNbUi1qmiHOTlaEgEnjeO3QOeVKBYryiRQjW4KB12+jdLgFy5XX61V0y
0LtXxr3qqOYmjDZ6suPEH+Rlao4mTOMHNndRdq+p1sEp4RnKfeqIk2MAJofpjYZUfcAVPFmTgpdH
JwaczEP3xYr3v8NMRf5c4r0tNwkIASJA0qPNz0jjLo7tAayJQD+GZm/E2g4+cmCEb88IDo3kSkIv
JZyOgB2evejJwYN8zmQaf7D0TBfIYTSttqRAKVKAOy57/GjrtHiOopVcKbwlHhuIqt5sJEbU3Gja
rz5d8f3wsLrQQJtaOh8in4ECW2w10QYYNjZ+9Al7DNwlLpjZC++TWeNcNSorQeaZthVp6svjxgLu
MV4szrLrjUjcWylWhrdNAuEOeMvfrFAXSW2o8vRnOYZ5aXwG67VqInM44nm0QsTaxrsHvXvXEk74
sXIRnXwrxfYuGqb+KXpdncAzsVXsTw4HqlPROB2hwQPiy/2lIZeSM8uow8/pBt9xmuluF9U7xoY7
PhvmhUVYnFo5qy7GUb19jmJ8LHKQRg1ICgAOHRZuDcrecHUe2AcgUTEF1rOkbxq+eScihHx96Az7
AoFe2ztFaCSq/PiHkI0SQhdoP0ACwj2lZBWE7YrY5RZ5WPikX4/aJRYga2zyvbuteHkSgM/NEiHq
WPRLUGNerooXZCh3EDdn7lnwv++7VhhYEMKG3Wc0AvgRbh8YqkCjnsrbKfT9Nhri6pQLfveKwdpT
z4jtYcHnEjd/157Tu2zewpsouaUHGNP9SmIAeM/Qo1nCVG16bqhjFmqKIsjdXiGEILIc8ZnifGB7
jGvcyenyoiA/tWibnZ2FdaOQ0t2pyj8jvpd8AUrpHlUy9TJ8vLQ0qtUjgEmTawawmB1XYqzmBZBu
4+L0L9JznrWtsxHdjDnd2Wfn3AFynT+APjI8TwdzN3B4btP24EkPtyyT8M2eERZ1wr644h00U1h7
xkHK5mK5Abz6qp5oV9AMGrVUUpPppNDrwY4fwsw/cEik7oh7RrtLewhka1Ua98UoJpJV66GzQGq0
CWRtssI3R7HUSh72x3wDUWVe2qWNB8gx018oGbOVaMdcQGrhmVryGzdhFP3ZOW6y7zsRqwuoZwuO
JBQkjuGAa48RQjqUfWicfjqBrNoecIihLrhGPsRppX4bt7+sJjrie3EXT1NWvlX8EZ7X+jda1Z45
aWg+jhLxj4pBVgn2Uj40cgRNqBTneRMdGRdnhjE2RYrajR9OmF6wWoYwVGbXaKr8oMlRCSfVI3v5
xbMmCTFuZS8udEdWF23T1LTLgJ3OUg273XL8D7BODIwtVUDze75/9o38glKA6BLDhB7q4pYeXs5S
RyGLqvKbEnMH+isECaIyGLtr5o/cefdA9QWY/eML2sXJMSpzSRTKld5lpcRpiluEEymLSSnezeH9
sScYEW6mlQQxj0owlW/jxHcnkwlVj5VoZPEzwRJEU8Rhu23oZ4nMR2ca6N4y4drhIboVB/nhOZb1
v2uJHTUDqDacrHT8gZQ/6z6TdiJmHi0/0ikQ3sVGAmRopb+SRPDGq9ROouwRUtsffxSJxKqZXFwp
E7yL7Sho22Dg2Zx/5cPGvNtU7t/QmISjnxlvXnK029czCqNMg05mpKbXh91Sm8Lc8iehrD1lbPSo
ok9rqzoyqeWW2spEGHkh6w0Cu0CQly0vw03zvjt9BSaJp0Vwj+9cFDTdm5K7eTKv2zN2xIwjAP04
9WFTrh0KHxIdEOBvzSSyUF+DY6S1Jp6O1Z3WkXQ2TmmSphq0jJRFlxbwqKbvnWIBvwVfoLvqOhv8
iHPVmU+0Bq4RhwmiSoO8c+NuD+Zax0Ku3PE7Dx6SGlKUiqOXz7eNTyktRC+jfY8XbOyULxdLnCdk
PLBsNw4K9qQ1DocQhl2PqSnF8eE7QQRqIDHL1ERsJZ/1E0KHM6JcTq6PjaMv1leW6Pfu2UM/TS5+
IFX4M4ogUwldTQVfGdUjFcyvoHPDlNXBLL0HReP2fUuBTSyEJpCVE58EW/illGXEA5CqBtttf5M1
6t5a1vtkDqG4ntiZdYjw7aZwQZlW+4H4TlIWiF2rcEE4vI1/umVACAUGRVNJ+azn+Q6b1uauiRWu
OL0qlC02xhAwgo2p28Tt2Zy1pfnwQUBkIf7bBfgAX+36VWQhgdNLaF/dgd0ly/brkqX/qdDRwsLS
Va96pBigrtT6wHVrRWzTj9Cbd7sLcEGB0yFOspdFTkPmAPD4qW4kbx3ckMmKwT3+qTSJTT8/aEg5
3AuZI9bAnDVeTgSev6iyvecJ4a/C5ON7MaaThe4h+nZclIkvsaKgDviySTCFGrf8ZWouwn4BFk0N
5DUqI02bXjqqsbNBtU7RHWAEV74tPma+vMJfqGtGlFIRAqM82j1zRjcDu03gPbKjVRnKai1+EB/4
qLmRpQXQGoluoGYzAVkYNR+3MRIuXWoGt6U1kjc8jETbVCfo/CnaQEsmvOnmDOk69yzRXgOT6hnu
GLFe6lMZ5WdBpM3ioEFUjCMyQ+ixF+P64kk/jJPBAkhxDPkwEDpEw/yDbrwr3j9+tSOr0MO5LWCS
L+8Tn7h+S1+Pwcbfij1CojCoMJhsSZztmzjyVOd0ph05Pa1AKJQUZgK7RcDNSGK4zMzR4Y8RGqwJ
4ZkxvQevHdG3mwwKnleeKa8RqtESXxpt+SOT61VXRDI6y40cy4IP+GFchdD24c6RFwQyCSosClfG
G+A1dPh6IJqrArXWAMJyjn2QDG53lfH1ClyNgFbhKJLESGjnt9EyqFhd92qeuEZFRjnji7P9UwCF
h3w67+THB6o2YUuMmgj7t5M0Wi/n1I5gHmv7ZwLM4+d8l1qPhcFHZB1sERZV9AQ8i9MXVejLbhkU
niFDlG4oYYQd6iSWCJfjdkK8qocPTnfDu1Ntj8yCAlf8xMNUdrpsGyQQS6tGb3jY1q8zW9NSa84N
1bz3lg05W+kn+hqZZ54YGheqwvxtvE76KMnkVhkM1a+rkDkOIMq4s75ZPSlDpps0MTNNhXm17/Dz
IyJNtxE+joQuU+2fNwmLlYKI3jBNw8kUbCROeW0YcUsVb8KezmLPssyeDkjYB5+9uC0xCZDGz19S
tyH8ejZGWYZjEoP8ZSQV2YD91/df/Oc+8ZcHsFQsnTNNtqU2jb4eZwdg7ToRGMrpiWrt5tdycDX5
Ug9uS478hR4MW5GfV2b1N2msnPd2vZ/DFt+WFng8iE5hThSPZsO7Tg65S+RaVlpI1jmfZbXD4ygT
cpj9uWNSdwD3rl78PUP/Euz2WmRVwwO+Lod+LG6US7hGcLE91iNpb837jmeNZHRq/csjf+HNIIPY
A7X9nHk4jU/4oerDRRTBuA9L2Vj/xvLkqKIqsESbjQWQOpUtw+X5ELbIx30c9sf+LNb6w7N8cCgK
uYKyXIwsxahveyuo7bM2BMnILRsUZHYsdm1xFIbkH8efRvGnNhxAtKzmt+DA9K0HAVvK98fjl5yO
T1r6L1/KiwmTeUACtulFz/Xh8v/78eHikHtM1gAENb056KtVZlX4Y5D1mba75TD1rI3TVfPSBKSP
D8FvjH3d4+yMRkI4BRlQDonwaAM4oZgLDoTPhp9hKbnYn0FUFqhMJoSOflBo2g5OHQSUAz4CMAZK
1i3dkgw0+HxptG6OE5UQcSs1t4RrDs2sLrpbXr+mknZoarJ1vgOs+Ng7+iUwrlZPhhna2IdTm2IY
Sjqeex7l4Np/9lLxOc2nMkOIkCNcWeUpS2YNnqt7Pn9WFjqIPt7+fnLnPqPG2rOVqAr2cGmXAG/8
caOM3sF+T15k3FUdcCtedv3o/w0zyow4oSWdiJjLZ5hA/2AGeJC4g0kS0LXxRA72SnEknYBxkeh4
bCAhAVvS2gOTCX8nFcPJMlVSbgOEHGYjNTzFbVYXuuYn7h5sDObEFaBmtnOpU3QDa+aDvWXBHdou
NotRZG075TmCD4DWgdPkY3nb3z+S3FmOum5JUiKK7SvOz0dJ8XsxZjdgXRMrM37N79USh13abIEK
FESDPuplD55kCS68o9QRQgExM6mqrcrD1jlr55y6AM+7yVHL3fuPxSy6wvZhC7oNXth3drQzP1Qc
fGFT1Ht7mPAsHk3PXDoOWsiBHxRUes9NyYOOJDwphT0Y7w+4/1QzjLhamFlF3+DP3P7eXNAQkV93
DxGisH3loHifsMiiXJ9YgVA/rZx7+I6ssBsn7AIVbXVSZ9jW92gYBf/ief4pYhpfBua5e4eT4ox2
bIerzOLXT+SKK1d2q3Ag8IVaqYDDcM+uNDXlH0mlaRVwbg9HmEfixD2uvTindnB+UsieoCZQibPB
cFqt3x0HmDWCvctL24LOG3EAlIC2zQ810lYQHlyjq69CJdjo1tWiBqlzmtovZT43Q+q4OZslm6w7
yAHSFJzNGUNb7FTD5fGRvGrV6HVdOoOH71p+3v+Wb3MBpjuJ338QFVNu1NdxciQiHYtxTBM5A4Nx
59zSIob7MdC4j+W95QAdYwjGB09qSEjoxTjwBNsjU9YF24qtxlYII4t4BWWTqQ4YyOlus1azccDV
rW0w7ccDQ3atQDWcY3KEDmjiSBoTY7feLfPOo5VBmJrliMsvLwFzBz+2dIwprZt9eXd3rdEe9G1C
ozqxrT2Ei2LhZrV3he5aLLpu5XkvRa5Dps9e2mv4jkkMl9f33N0S/zz5Ed79nuqY4Qg9oEik7cWG
ykzW4GeBTwlAV4liy9LHdQsoeyl+F0VErH7Sg59eDBB40LF+7N42I1A4Hr57ejsus4oYsNypnK0P
k3YSq5yfHmZF/OI3bqQRekC7UpjWCa54sTw7k13j4ylv4LB2JScmoONS8QinTwT9aehJA/6X0AiS
GdnPKen96D+GnNhn3qaGIWeyhdXEYEoOi7qjDtiQFYZlUybQZdwVfxJWFUSMpBitWQdIyfJrUCzI
ZNYPUAMG1wFcTnXF6UPvw2o0J3USUA3hwJaaHL/ofzopHxR0OdFLbIOI1sKskHzlGvk/MNk9GMvq
2sh+RiW5KASy+YHSHwtXC05RQef/MgSzYvCU0a+/Chs+hgOlrpl5Z9EftvnJDHECJRwX5uhiQRo9
H/X04Ctl3VXG/TOX5nSXiEpdrot8hw6lxa1bihi8NOxDRXH6gCQVpK7tvQddSipasT/BsQoKo1wV
eP93JYMYWAZUI3zagLswowDRQrd9rvx9ZCtdnkY1WNr2gmqJrvOidy1wWrsZBSnKi8pkpmjSXA/R
lkZKSRTmSiQARiHWWLH5fOXagxIpR0i/QkgWAWAM97N0/Yi1r9LW5gdKBdeMHdiIgrn7+1RhJiM9
y1oyGMyVRk0XUXgwwTCmN6RkQuAT8pK2/sORLqCOhNNOhTXDdRYX8h3cOAg01RezScje9rwbtyB1
VKUpnRGj/7aHjEkK5tjw4XytmIDQ91IzJtavHrYYFWI+qKPA2t3PuI9QeHBoCJ1mUFg2N0aC8I+x
8vPn5ZWmutN0+QmRd3v9FrqGP44lpqAlQu3MhTZY2Lt5MfM60/Xq4762gLPbV6ZcPxThfC60qJ9n
mnfZxKnYIraHLz5fabYBOQMOxdufmuoQk8SsgOe6hY/q9JImEBCalZaNT0QWvBulp5YGCoqH7vaE
8p2w3mF8omAo35aEmSmpF5fqrLZ47Y9zziou4qlmD/SsJS0pfY8HDlMYE2TdNvieKY4FAK7aNCJK
Cj6MC5o/B808+Jl20FJyjE83sdT8Pe1egFXmbuIAcBH8xlIDs2wo2rDBZHtwOtLxUt2OWyeTlhfA
u378aycs2bx6VE35foy1Byr77igji/s3l32WaxUe+SjG3khcx8sskxYBxnf2NkPjl0YqjpC8QzxR
h/Xl1tNMkA9bJYgaAgvQE6g5IjUDBAJFwRWoNb/oHJyXulZ4zxc8gCT4i1+NpNIcRQ1InDMTZhQD
fv62vJaEg9qwSvPSnjgtoQkR1FfmYWBtrhVrV6sQ3cfjMepCvdQXrKozlHAfGfjlwnMAb+yNT4nC
iE3bYxyGVmqFCVA7kupkEPhfwW0cZ97P0rB8DuTFniAumirMmHcfqVoky05noUYnTDlXKRClpsB4
jDMFtCG5xjB4sIPCBbdCcATQgr+MDERrBEaVq3q45hIxHi6JRN457Lk07LKbBw1MAllaJZvECtWm
BqIkjDSIC6ZT9pgs12V3FGfsm4F2VJo3Pw7h+qvUfV0iWW6qS4BDHfiMl66YpGxrnSy9yNlClFVw
rmT47u7WSDf9ufyaanUU+1gbcwLzdMFoPNRWTMQYz+tHydw52aj983NffJY6wOeTgwWDV3WbVK8K
64FIGe1pgo4PU4k1ze7SsfgGi63XbV2ZA3VzCmzH9YhYolEsYy/1vc30/AbD1Jyt5riGIfvTwqGO
QXEjeSpEQke7Ur6LX7bOva0VGqcbIr3UlD5kWAgsKreSDrlGb5Mw6o1V684oAMf+LEkdxSsYr7YN
Rty/mLX2qH8mkbo1onO9LuXh/o8QNfT1hXJxMw/5L57RZ6NKUyiN8RylQ0IKTpMXZ6cP8EVslEfX
qZmxNfQHhdbZ9pgbLNwMaKrRifBfJj4oFjG9gDNo2eWtEFUvcQZtlPFi/39i/WMD5XwVF17/RdtO
9cYrtpdmk7siXvfavXe1FY2UhBt0YPfReWtUQ6QZ+k1VQXl8NorK7LU8mSEGYxJdFDph1uyg250T
dbK5ZECGCwEqVyzzbD0ynbEFQp5OcMHMs1x211mG92M/LCs28haAqF85dLImuI+Fp6JsnIXniBZi
z4iFdzQ16XYH3kx0uTimPEGiEuEN+FpfoNFB7nD76VqImeZbE9Ek8U8rGhZUfFkY5iqGZh/7bNQr
TO++1inGiXh26PQjrWXp+o5KQYpvTNIKrLvXvRH1NASGuccWK00iLiI5Uq9PgNa7WmRBTtylGokr
fmVG/FuyJQWO2qfR1ZvRgi5Z83kjyGBfud/7RmlcHMGeIZMRuE3qD8YVPUCCBJ2D+2wVE8nsXFes
YDX+QXT4RI5bofJqM6TM3fMYqLFrbSIGQU4Cd6XjarAbAAmHsTj6HqYgT/bB2DYSaU9vf5eji43U
RsBByMR1PVbhh8YWcXp/ZuOgZvIUxIk2v83BDm63QbfltUonIxuqSEHgmPSrYvguAvxvMaIswE5C
EveyZkN4tCFL9i/1es16TVQqcJxXbMH+Rs0KcXVgdTW1j7PJrERJ0sqW+xHKeivOMsSxTTCmIQxH
5x9QdRmlh/iogJzaMsTC/kyLKRIGiMs9MeR2ybCTtLD8xL9I6RWHdb20be1+jL28+/8c9ldefYSG
tUbSjCzxZqU+uORWpfF3JOl6VKGF4OyJvbuX9ux1MpYROyj5rXBn3ep5+qIA4CjRNMWfsssr/R9A
gQfBRry+JihQWFYkF/TsG+LwVt6VrEglNwR8KFufyAdohLwtF/l8HcDA01r2oeWsdtQJidkdwlkw
Fa4KW0e9AgLp8TA/POYdQU6oKdHXg5AvAahWq52Z9SbYFtT4aiykVuQ+ZneYA0n6KL3FSyxcDy6G
SHmq9RXo+o9yPzLxX7fO9g0msHsvF6fJvcgZryvol+Xzekg1cDNkveYsMFfTCDckN6BvqyD2Y7or
btIFDVoX0gEg7bvAs3jyKz5rvdW/uMbes/cgZ7r1a/0jHL/SNfS4he8yIMlx3pDbPYSF9fre4fKU
6WQckvmAiMphQg3R0/d3bSf9u6PkOvNPAltBlKTYckmQZ1j43IBIK+S27vlXQZGBKiauMsENAl0o
bJSIP63JkYpiLTUUkCDButI9PBYtDmm06YJv6lVXhcP0h3mWgasPdSsafoLOoRAH0OnozBx2oxnT
IqleMGY1Y2uXPVSreQa3lbldHFBWkK+WtoITYD1VyHAeXWvl+Gfk2uBNCBxp8+DtCcmU0vqgleuf
EoBGydpkK9ut5rZCivNmeFXe+H7qH51d9MZ1ygCqqa/wUQ1JqbuqekLKWClUoj73gOXlpYGrNq90
O5xKVY5olt9eyieRX7metw/av8mTIL6jfoqLNTJtjnfi62r9SCcQzxLk1lebyw56IQ8AwBgZjOIQ
LfIKA7j+B4NReg0RbljbUe/wel4RMYUGxDPoF72sfAWZ8nb+Vm87ol+c3UitPvWqtRhkFEf6TbnY
t8JZXWN/P2X7/GAPlNHeZtheEMyg7nz0LML+b9giGTXqv7QHu6s75+IryB4S+PW11U/lSMdaE2ZR
UkqFkSnIY+OFPWBjMZd6Y1cvuZoOD4Qeq7UFP8fsd2U9e4Rx2ESvYwibsx6y7u96yQUvv1Dg+cfn
Lhl/XyyYBTJLKKcURpSN+/EtoRLj4tIxJjLhzUyrYNVtGIlFNVulnAAAhLGRd860o2Ba9vbuiIzQ
5JOoVoBWhS5ym75LBpKerSez6EyoCZ6zRvxSGksyIJYOAb9bZS/220E8CMawIf9qcnG4+tO91JFl
qZ7xng+hMeqvL7+jsJoOwKMKYQ7S/iS3qQODfCS4lwpHfJuR01+ckKrKEzsJE98+EkyeYmV4auBM
ONd8qpWpxQAWNt4Kj5q0KFgFxU5xPMChooS+l95eYnAoDT2/Ri9PsNWAnD9v8jRHmJNQvoJ6B1Tn
WboM/DSEXxQKujkiEttFGjb8PbVgnXt/TYVBZ3fvcjtJyueE+RfFqPn0aPlOO8WEZut1HbfNtZgc
EaYk7nZJSuU8nvF8DexuR9BQP86UJBuJYWMdE2t1uZ+Yne8e0nkucnBmtgDwuxHFdP1Gp7ntq0t+
qOZZXQBtB1gOe1oREjlGyVSVHJzmIyUnsnvApxOAPUo0egliJcZnz4cwgFUYpfKzI7rFd6hKzz+P
pnJfHMtgrWOX9kgmuorqHN0c0JCSbkvvkTjI9fBKVjgb3HPMDsB8dg6WIM0AiAIA/jus/12GZLcB
NCfC9y/snhAypx4k9bWsCV1vJHu5tm68Y+SFpybcOBruhfAqkYNyCwy12xMps74PQk9vQZB3yzbm
f/PXdm5hx30w1jCyGI1ErNMa4dectenPIaGYLmCAeCcqm4bvB/vONOHXydNmQ9dMJG5Td50q3KKy
kQxexwr0mKQOik/TPOOOeU49nLIOomyNi8bD/vF6+P/aV53sTMFzBBwnbv3HGu5HoFU8viCKgnGt
NXiT95mFg9BVcP24UdMmc7R8+4XjuM/cWbYGnESK9u5rRb3yoA38BycFnG4uupMjSCgjd5KZXAqj
Y333SeCmg+8VKzAN2h0/q1Q1b+ezjrsHqimmNOhjP0ENRnUJteBviXhgV29D83XS4yHyLiDjWsjJ
8LRgXWjNv8Sv3RLJvdpt2WRoh2WTHyUmRqpOYeKFzJ0QRcFXA8wMQ1IpYsSfgrrTuNWNjLo8U+s8
kz4xwMYiSVb425w2t7+3NRKsxJEVK7EOEC7EKVi52DenHo9UJ0YFHtBFlBCnYQOtOuwij8Npk+H1
gadHrwzT6mxTYWwQgsFJzzs+07wx+yQslExwyUEICY58BLr0U3uVwq2t1LS1e6hFd85VZ2Ir/v4u
HTzIvGkesLoGYo9R1HlV6ATqvILxEjZ9XbNjQJ7GDNIOxZJylKmBPCDKT3pnPS4KpMPPgz4PHgvB
ZQ2JEcJMs5TkJwgcJyrkZxhv7fuy55kAWsm/DYmldd0/K/GL+HZajX/7x0ozUNHvqQF/WE7+Z4Gq
sXr4aCoG6gBg3xtaPSMpbgWqj/4BJijl5Axmg+sq5Y95BrCQyxWtvfbZQ1e5bHtUIdgCkTt2LoI7
MEGGL+7WJWnEEqYdxw2c3YhjRE3A9pj2WZNaOjCP1Mz5YeBpDddGRymdkQZWys8jrNWEjQ05emqj
smuM7f+0TTElCRV9RSh9q2aNhWRJX4ZztVV6qt0OPAXCuk7J7BQq+ujoMLXnbIIPCo1qqhMsuWyw
UompLjphAc1G/DfGZdB4Uucx9Bd4E0S/Klok6gTy2q2rQbuahPsJV1xDS3iG9JWfMjyCkwHscDKQ
4B5CGcixa7cewuqiGbLOgsColbCLL5nc0kj/MJgzFte11+FXaYjbBdN6WnXEEk3FG0iOsMX0I9lI
3eAQrouVx+BBhTsAI/V0NAxFO6KsfBCH3UVjGBXz1Fgbnz7rGEHSJmAyF9TY9h1aCBK49OcbAq98
liIJ5lLqNeLEpSqfBAWjcNuzIuZPobGLPtjChqp46DbJseb9l50Mo0uKQ7PoGRF6VUIlVij84wrM
0mHXRlXzsA5U/FHLhP2A2tEPh5TZK/hQRdiTRoQCZA/SBsqI4KoVqZm3uX1SSapn/okFE+Lw2I5R
qDWVIUOzINxG4n9fYlA9RSfCsQjh29QbKWL5fVkLKiRB1dmeO1K/BYJYElqJ1aKyqW8rXChAX+fh
K7nLhyHq5hN0NTRqxMZMiGscNvVgoObmRitzqZwK1qWpVNa+crDK20UH+eH5pOMeAGzPIhvkdZa+
/okX1Ii1IYwRdGusc3T/YIoc9+Vs3GM2Hv4q22SIpnLWE0+pAdLlwlOkFn2VnQds8ZuYYsgZL1of
ReR8LAaDMZ0Z4yrauqvpRiy33JUGIDPGQOu2RGDjBRC15L6Ibccy7eo1vnHznPbc9KuVE4ssjdGb
PMdWAMJ7TzdOzhl5kJrnz2GLAK1RuxptZt9/2jkUKDBYq1Epzw9t8qD/IGLfVlrrf+ERuV/t7A8C
BKYE9Viaba+bSJ4ekzO+kU3M4nfREIfQ5cwV97EoMRHPLf6KjgjPECMlpolGyOUiPYgKLhd2QI61
erA89uv0BMy0NywubSHBFNlgwbx8vahDEH1P+lj4GgwWwM0shG+XP2mqYr93Q95TYgCThs0S1Pk/
2+MDZW+amaIHPzvbB05YpVQhX+ZfQvV8A0+igImsjovOrhCla2kEwyxfC8uk6EMfh4p8WW6Ot1aP
rm6A92nkHFxEp8v0im3SNFlWXoe4lpPvhS8GTSlvsnjUqNF7QaOaaYcWljlb37w52i2pbrUU/Cqj
+1F5rrTnZFPkDZQIvkz9qaboAu6VU3AGuKK17GVjkElPs6fc6naxGiTwD4w9zKXDbtYYFUHzOMdj
ayyTBfMwGS3prnYnw4nik67TDhj97FrHiMvloyTP8I81Ani49gU7DXYozRk6MvStXdiA4i4jnWWD
LTwVH/VDqjbJA8xPdfm3L83/IYowbPzt+fmTw/ijp4tbqvhemjHJ34ENq+E6vb4Bs7tYoh9r1ZzR
vS6tEZKQ6C3IGCxg4F+KdjxtZx2TecG6jgrf8P5WbyJFbF3ZTfgiXkjDTx+2A8h3TaFar7UylXMm
3+kKrZ7PXwjnXb/2dQol5QGd8hdsczds7D4h2yR/ycNISURoZE8v+CtvEEHVyaNfHyEcpZFEkNvr
fnZTvqjc2YtRMq6zi4lKXw7ZY8mhYPgEFiqyU0Kz/1jWKSrxeWyy/VAyPJZ8roQlQ3Ny3qCBHMM/
TUsmoKdzYVXaDVDUWNfMMMYlH/Ygdeq6Q3nUz+VR30CN19oMLDy4djKo6z8FAipPLpKd8VT2LZoj
/2oW+0JQK7VpP0RiChvL0xqDQ8692I+/pt9rmlrfjd1jEQC3Y2XuFTQ2HbnniD6tW9hM37JBEUMZ
29cZM1hx2UoZPypVoApRAs+c5g0qL5zjffodu2f4KV0Iy9n/SjkVMiNva6/Ib4FRd9as9blVk1h9
3nWymK2QrQqamCXqdv3zuJqcZIFsCYvt/YwEhxJneyGQuiEgpHl7DRePzskmhALnf4bwsIhboqTA
KT3BzEJKdh1i1BCGl/4Phwt2WKScebYpAjHkwe9BHrXafBYf0iq8xEVN2Prcd1n5Kc+qD5EPrnH0
YTqFzvPVlphlRppSDY4Rgiq9O11QZfNSZvkhJRfRcwfCT5chCmVxnFkzjKKm4w/sohts81tUrgNz
Sep9zNR2LbAmm8iSZFBpOyq1IC9v1RFYu0SKTM1WGR9zVKj7rWvAEQmoJgCHTZiLE4SWG5Jhag30
MOFTuiOLMC8LdhnlDLbHJ7LJx2ldND/rSZJVupxSIFwdLhWqDa81wqGrMvdbaWethabHAbLGBHHH
ZaxESCq2+XJbdPQdFyQjIjJ9EmiWqS5e0cNg/3v+IENLHkKZ1B6bmh9mxAfqXQXPpLiFUv//uK43
AI4GjP6IQDgzGsb83n/aHPwDPP/fDhihM4HYwntT6XnWJKxl9Jb5X0wGhG6x0CpGgDiiC21X1EUP
f2WwqoTkfx2tw0tJIvLX65z4euXO7d0AYozSO06OSKPaMO1MiMDB3cVmI/tdNeMiOeGPjoOH2CE3
RlVfU591pp1TBsdHQKKT8+izlsFEjjfuat2HnqEjAZi8hwSqZppA3WsdjoOc5ukXWv3BuWannt4M
GGyASwkw6nxtem9VhMATWUjM6w33C859VgoT4mfGfQs2EwQbjaEE7tyL166dYtGyNhoodnF6tHYY
gkLRi9KeUKSFKqwUfUg1+vfB0IKfjWB4Ewji/Z2lVB9W6IzG6FwIm9AI+CywTA5hOQgbbEK+o+2c
gg2Qhw+5t2GMd7qx4tEZhd9kZgDwurAI2ABy/Sy0Pk2VUsKwZGXRAWEV+Zk2sRnttNaTmgTfUoqF
hQP5gRHc8sjeInYVmsbqWvuz+Zx1TSnlJ2ep4pOVPFhc/oNeBCkAW32mzyT3B1ITtJ9BheXORAmO
Nsz3QhjLHrBVLDdV2lQW9OmtauJeNxm1/nGuU6UwlKDlhxzVFWXuCIeR35kz+VgrsHePjieoEzNL
UvJ3wTPAAHPe86GR/W4sSk1yjhfBwdUKt4AZbZF5j3cUQGiU/WGD+6GFDx947I+yVbZ/Vy8FO0fq
Ax+KDiw9BKKvhsW7jWEF6OUUPsmY0Tbf1+8YYyV7SyIeeJiCAmbqpSFCk5y96w+gm+FYZpSwtcnT
TKwR7QDHedqpTnT8JRgSXcZrYE2QlwFuH8MMJnMn5R7eUaeneCEPlHpB6zTI6Py/YuIchzFwUtgQ
SkyX/8Mu3IEEif5+iCRWtocqxzCT1hf0uw0eimte4tpIBrPratDoerinxhSHqqQQwgUTjCE0uEAd
ePhKu6H8ZZF3veqhIIenuHG5rrGyd+M4LlDgsJtEbChKVXiCO9lriXhhk/Pa6+Yqs8PwAwiQVTlo
JJdRWR1FC3NjReAML6ir4lGT5GolVuGwb+tc/+sPcxy8+TlJOQZR74i/soplLbnOYTJIASRaxu5W
T4BRDCDRVxXW3YU/xhKmBKBKWURBcXbU0xcOnqyFhnT1K95f7+BNZ7CtQRWPHjWrgaJ3nJ4Spewz
J+PC73pzNaizwBj/dgqmFeUIVWnEsh1hzYpClz51CBiVxLXpStoslrS35mOrpWMtbHVDpHkVnwHp
DeOEk4gL5yPM5iy/iZ9cg1bH4TDwkjqLd+jVj0y/+MIpqkDZ49mbPLEXHf1xCmybO4vC2cZaEqy+
s1TZ9CbeJsRO5aDzKPZGel+49c/Wy6YHBwYFyp+I13Ej69gQoRuCPWkWslfogtjeXEF7iM9TOAWI
oXtNHkBYoF05mADRWciCtZC50Q/+R5k9LU5Dhvxnqr7ftrZoOT+hNgauFHuo8OxULnALJsF5o9aQ
0wNqDt2g8EDIDWRz0AIDsJRqYvBi3msEeaTnSNaZyVU49/jIawhwd8W16LvwOEWRphvSm9K0B6VY
EUMOvaxQY9GIzfzy7Z8jCUxDPqciE5fnZog01I6ERhGdEYiUBp+jfIDrm/2OkaZnqwXHzJ8PuNLr
nCVo1JG/Xx4gA91HFNC3i26+2a+jtgqiMR5Cf8XDjR/82sPkHKCeo1S4Gu6/OH2M7/OV0VBNN1wB
zjQ5gXNEzfL+HjUwm0ZTXQm4WFQWnvEpuBcliP7QHFvMuX72dD8adcut0MsfWkqUjbC/IjES2w/E
xXiRS/2wgAI6gXUCmT1PGSAydvyeOujVly5S9bnh8VuqeMW4xZ90PEWmB1yDG7O1TOeKUG5dimNi
PUl1YgKR6S8lbY3H7eOsMd8j46izZ0bPp6ajuNWxQFvKrfGR2PPngez9kQcVjdQzIxAaNuAXQN/h
o3p2AVEKHuJC9R/zdSOZ1SJqsK8iruBeYbl7MwoPpg/w6tAHZhHKswxNyCfZOoqmML4zCf2GWs5s
YN9HTcjw4tOZhxwBf1G1MEcsen7sHmBLwxp8Adwm/EAi6yen/lDIR4P2adsgOpdC/f1J5f7hHtYL
UKRgd5k1rPmcppRkE/cDqJ3YW5ElUHn9AGqzAX1SKWBgXASpNClA/4Ci0VydZcur5LaCP+gb6O9E
yp0VryMSAyBDAxwhpRgDzEaAsfei0ByhZGV09T665aCG3oFB7JhlXEJf1jvnWjuRxVrGXQZYpCGD
g4Z1GioxpO2IjyA/3izuQeEcHgOSyvue70NCccdDoiZbbjFqw5RPgR+5VqLmxmXoBVsUDdvTLbnp
NDGYMP/Vhj2Bf8Q1D/3aPpDKGp0qUrVaCogwm8xmiqdnhDY7517Bhj1tEdsuuqtFAZn5XCcv4fgA
BPavkO1lyNoKLTSE/8C98/ZBJQ5H8W4MIcpVQ7ahpxpxongo4XS9DSnIXwjjGbV/SpdeOsFDQBme
F//IR5sNZcGL3wuWRneAVtkVGNaGScb+mkVasjoDG9DS/nKaRKEsQSmAz49tyFdmaWeqsyHK++G7
/wPDO7QQEAEASwrOYHgjZyRq+l+eE6X3WhFHjdoJijlEy3n97Qq0/moTtJ6NF5m/JgaIaV4qVitE
9rzO7Ji0p+1mrZfDegqKxtEKdIvvO26rMksPTbseOSRVXRQ9WHvN7FBqWzHPnt1qfWFc5inoBp8x
nWzIiwOpiLtCW7oKPzB1bPhGG6YoPz1Cl4LFgSBn4CYKeA+foNlTJCit4yz4FI9yiB4GBGhAKNYP
Kh42kEgiBJb+Xy93fB6uAlomMqlF287symLza8V1xEOBhqyOBw+9oVq6GRPOczqTAhW+W8wsbSqS
/ET/9gu3FXpBi+veW0foGc7HiD2/UF5t5VlobAb9a4fhZe3kU1u193HjNaqVQ32p8lfJh+s6dbhE
jKK1f35Kgn9tRhPwMVkd7UG12YKfxEDIPYX4pYaOMAD28YdDS9T/1+HQu7yI5+l1M3pXTgAA4ZWU
JEPjPmmfpnwl5VHGeH4yK3QJMARcHgCWyey91LRWp6FvvAVNqfaGyivFwtXIGJoXVpdmS0GAcn5p
3K1Sxj4Q5Z48RH7/jdgt+3+Dw0Le6X2x789mdDQQH0n+WYMB2cj7EJfelTmapV0Pj095qVm/IaN1
w2QfaVx/VHD+gtVqPdW6LbMgyFwDF1vCVYfomo7AbQpF6VHL6ZCmuDJRj+zjSORTHwAX8gUQhGqb
fYqosgnt2TG64Mk4s0hP4+iUDAuxi2YoC0+s8r23RRgN13ZCidjJjNPXdt4cMaQVOHGQnCASmWER
MkSdlsVnRXUagkH0GuXMEEnITQ0q4a+steRx0OrSO6emnkATr+hTdjqJL46YWKVMxwI3kcCRHhNM
bB9+J+KulV5RKEHKglfnJk+zm/RsAvtab1df48Q1jDeY0xY9/vD00B4BZDoSw6ZBNUGCJV6fJfrK
s155J3Ft5A7gixRVLfk1m8EuRmXja1P3PJtYWrSW6S0VMzTpYBBrebC/guOKqL+92iA0ckwH+XAZ
RZW7IfSjCaoxW4dx8qU0jkN/IqYT4ZW8+0af/DHEfSXmQQYBkForxbxFxGcySEUwLmrQXcbSvOBw
SL8WYFseQoP6MczVIlVdXmWVoEslQ/jdIlHZTivhyThIh/LI7VTcV4H6u/scAlGwq9LSheD21UPe
7vCplUgyYv1u6lgCcKBkDCIhlOZK66Nd16VlYZeOe9lLcAFmPmkOXUn6ptSXGfOKv5PEKKIrHdaT
fCEWUcU0O6Ppnn9TLeOayNuqOEwtAXscFkB8lJ1siwo8SQiOjSXCSFkcW15SOdp904Qp7Fr+JspT
gXc5gQdAxExPK7UVX9nZ8HV6puAINW1vgdTPRPjn5IsiNLIOjXPLsQOL6a8IqxOwI4SldzHx3fQ2
nr4Bs0ffRPaze4ZKUBG5ryXJhBeJ9/AD4uiZoDQ6QMe/utPHsyIvVeEVPWM2DJ8pXyeu7Tih66Ha
8d82QUoHWwAIeLxp4/+UdC1/hrF4GVlCcihkJuEbPzYpL9SoMahD9hvOJF1JZsRjl0B2o7awZ5eT
5z/9nNXvTXmEsjMG5pVzjFA+vsuQQiYwKpaXcH6VtZZ4vVGgJpVYbKx5RKo0al6bbacqsQRNqxhN
Dt9pdjp7GDf1qqLAts5j4cHKLyel/unmBtGPQy9UIueGBWM2mE2oIKzadasrqWGiG2hWL8mc0B67
mIb1vnX+Mzq6rPxZB225kYWUPlQSR5D6K9VG37C7SJ7PWuLyKe5EqCuprEXZQ+EeYkUShMGXwEQ7
fw5H8v6a2JaFQMcZGb230Vo5uI4MqQTu1za5fK1tLiY4Pp0ZqqXDJHRqosW+whZRbGd9UcCET6Cc
+sbz/DLAtdZY5+7AugfmLNy2+r+PoiYtZrNfXnmSmcXBMQfxwxJt6hyh51VZkn+MvvKcCX3CTCUK
x1L75EHiIR5lq1CBm677ReEP3iXOrBtQOhX8OonROmh0ASB9zizVV+vSF3awcYP/GEeKBKWnImVh
4iABJbuUKWo44wigYR3DQCKo31WR6Aop2c4AVAvfa1W/kitIsNKgEowtvLnxqXusZ8VivHJSTyWX
0DxCP0vl9RabDz6+shKnf74FhLbwSGvTz1GcrgMcaCUhzLWr50y69tE34S7GLAwdYb9r85ceIb9K
k0JcvR+u8pgdoL3o6FlUm5PWRZ2Z71b0iUUkw2LRwusdOAUo7Zku31h6KCr4OBkPuIGWaj1SBWW1
wyfqywZzxXUnTghgzJpNVbL0H4HvQWNkwymR1RNn6soRmWnoc9igmV7o4LtNSFA6j3RZpEGZ2lIG
gxhikWlPt6FKFFFUpEuyZdaaNqKVTzp+9YOBPWnCuEJbr5sNFiXg1sDpUR74CjYPMdRdgs38ZGDE
ddNAoCrvlxuWIX3B28SUAFzogomSXDXKKoKqSrGEHGcIaxigTjYxbH1Rh1FjeeA0+8o52Sv4G4Hx
figYdG8m9DsleTSt/uABfBwDhEqB1YJE4/QLgzSyT++DK+kbHYQAPdlPgkwW5Pmh2NoFvWpGq3uT
8N1h8SsAY05DQFHIkmwX6r/Cbugx5YLlTpOB2PFN4z0ByD3AptIzkMk/F6BdaFQ+QE6k68doHHhx
gG6Pm2oO3/ycCbP8Tso7F+eb2zZn5zbmQKCN0MnNZQMOqW/UeSQOYmmk6xDsj5nTeJk4bOfgLNpB
tUHK1aTq0/7v65sbVT2pqiWYbscho4RlqG8OQqBGKYXk7f/6O0waG3Jf4L2C7OsEutKC4ah919tv
NMeveCxse/apPGD3+/wCsC1QPRyqds1LxZYzBqtilpAWsk0Dd3ZF4eQyXsf8MIBXUJTBlk71NRtD
j4RXlFsx1Y8vXxXdP8zOj442iwE7yB8mNNrX8xrhfH+BySGu9ulOhkjeb3YuDdQuMSvC44HfY3vN
qgcQBfBhygeKrGHwpOUKU4BB/xMUqchuwm1O24E89YQae3nOrzdUa/TItWN+NpC0rWRUe4/JmsEA
UMB5UR4yJdoZCNMomOQJxDmlSAcXOdkySZiVzJxtKacpbk6SdXbij93iKs7YK8FhqZjFsOilgnuO
muK2MqfTHZECGd1MHn75Cys5jg+HjAlMiRZlqTaaklcZAOCUXNsz9eLBpj2GiOuBZiA+os0r3yfT
NYqmqUJTsBvCLGB8mOjvrt2ewY+nf3mNl1s9raxQa6N8A+oz7KjJuIQ8U2DmOtZhBeM5Wm2XJg+2
5U03spEtbfr83xbzV4vyCEIhu63MBru/r+UG7qjf+FfusdNuWeggqYBJA82sTqncJLU+9ubVV+7c
FlssKPsupWt+Bm7lfyQyNeZlMnqaFRRf4J90YQoW/CVKwA+ypNFkL/WuLri9nGiHc7aEEYc6pMWz
6Ok0giH6yJL3jlJEpaVIqNJ++dX28VQlxzTrfzCbzVNZ/HyamjprirFnD/IgMWvzI6BhX+PJW6nj
D4lnLUK2HqhgCrKtKljEyoyG5sypqPedj196wmc/ApehtcehUjTG8ktfUMYsk6EuPv5oi+vk9Xzt
ccJ3zuDkAMgy3KdtwDbs2DfwppXLxyiwDOZ4t5OyhA/HYaaXb6HPxY84/BXkhthDMvLkiU18GDkh
1F0HGtSvderMcermUId9gyfVGDGAkA1EiURAs1Z96SebWYIw1fblJ0sjUq+gjtVBC457486RHXD1
uX47u3xL3msij+/t4i3jVYeNEq8IULJpn3/dmytgacJKwm4+b2wKG6mwHHcXPY9pyFtticIhenII
FjtZyFsASINkxwWFGhDCC7abBjxJreBlbZ0sZ3cQF+oZbiK2FrrwUoisgaGvkLOERr0Lmmj2kbev
5ttsX8+Ob6CjbfadqHy1WmxinfVy5+UYwC/pBwUZl5bP2ZNpxeBb559Z12GWp6NPTAMO2TKHxf2m
FDX8KKjsEU7qCH0ktdeEd7M1oqfebcVTcNQr8jGzlVin/F/63geZVT8xcrPGKT3yKTElofxA5gNv
skRwO0DtXbkJ9WZX4OFhDYRDMS4ZutCramRGs+qSPBbpMd+j7S9467WPJhGqi5pXybaCWbplWPh3
PpuqxUfemxYz2b9Lp0Y8k6ALC/e1cLpdjvGyBEgVwCNLLh31H7Yk41NmxMuFYKy3KXUNeiUW3yh/
uLhfw80zAud0KFcXcGOue/dUi+nG+7Tn5MI3rXR0PjmJKTPc2UVnp0xW82WBkmfeOI8Srs25pmBE
04v3xQD+nN2mtkoJAUfdzbMzecxczfcRx5wyk9xoudjvV3vui6zKal+nKRM3G2Qkj528AS906mZq
vIuqEp/zE494j9ja+21W0jYCQFpSKrZ6XPVaupclBgT7RTvsKi5xHxjF4A28kjcJx3vVkFqf7JGg
2LObL0jNpfxj5dnaTY4o1Gpf1f1x0MQ7ClEg+/tpjbSQEnP9qKIVXs/BE7Su5W+9OdU841igRhqs
VWkwls0NyG0Ux+oRO/R+yyQP3gHBSbByN06TyyRGtAmoy+j3De2ep5a7Zyr0UsFb/JmVtj/iYO2p
xxJ1JMVs1Q1LY/Y2MlixvHBuI5ONxYJQ57/NeqkLqodgJQk68GgcUuecv3pK2F5D1hH6gWloe3es
hpmvcVurRKJRj/3EMrkJCi2xzQ92p0L7BCcwH4z2V+A1CiJM4c1u5lH5mqOFCtQo4ZDwS8JO6pxX
DzzTy5y3rfaU1eABnxzlJ3YG7yuWiTM9sYUd5BNh1LudLycjhMnke+oUteWBiwytihRQWYBLu+hY
fUdjOKmU/mCCLzIMXg2ozG1LiKJT94AGd6ovjJdCpb+fb+r6aMLxTCYDXzrUpslbgTk8CsgAQ5gU
DQCpQOLF9/l6RaVT+xH9uZdJbgqSBwZkV6rj691AP8DhVPKScwh0Pie24RSgv16QLeyFOadqDc0Z
f6D4/qAZe8GmI9xdJP/VDBxkP3PqMfiIqybDRcF65FKd9q+xCfa/3m0IR5u5rdNmpMSoqKbbYEvE
SY3XbWXuJJK5+bdfMdjBk271jPn/IvG85hM/lymuu00jIkwx+fmnC1ehHAsHNJt1AihiowIizTmc
x7zC8Yi1UYuwJkyhPsYRMdEeryygCs1ugVHsv/n0JmGPw2bBlT45zha/g6FUVXe66GRVs02tQpby
6gQYmRWbitsq3WM0swXCNZmuYvewnM6huR4u6pBubf+Ii8JHOX09He7KL3XJB6BLsBspH8YBYTl6
yRyLUfmo2sqz+T8ch1O/SnCTUCHV15P9hTt7ylhc11H4tobKT4CWnHPCKe94vgfglGV1kXNqI5FX
QD00g/lBQi/Rn9GnBFuAMGnPVFyvWk4QftBNVYTkaQhjhTPKYfypPAnbX9uA/+cHhMzVoRP50uzu
AYdH7l4KNUPphV8yQqruWpUOR5T53wtBfx/M1zP25VTqBqKAM0KYusBy17qKEhcODWCZLdU0Jouj
ccWWXYfxavXFrr/kFEFYNxU4UvAazlce+eEige8ZbUtWqlTxp/kPFadicN8rQtV99763AoKpUqFb
kekda8oQ9hQQR2wCGYLcNMsslrT/c5giSAnm/Ze9IgSDUe2DLne3J+jD4YHrJ5G1APtL0aKOaoza
z9Xfaelh7D+6xdbS4EagkyS/gh0Uo8DKec8eNLNeca+v8WDEjhSWtmJronKMGrlFyn5NJY4faxv+
Q1ZoVlvlrLACNLmoOCAUFtF8r5xzPQRawi3GNDFAYyccDFeosSY5jgxzwmGGdKOp8ttQyfJk4DGU
wY7U+OWQnW3Tn5SS2DKFk1dPI7lHGRRo0w48rGJEAsBz31d4VfnLCbwumYTnTbGycQQQmLdb1QBG
1zSNtTgxw3kAQTOAW3uc95aa+I5YgCukpTB55Dbov/xuozmAq9TL1pn9OI56JXRpty7QfOk68DaH
uzBRHOeUHUg7Yg6Q1Q9FO9ycB089+4viMU2MoqxM+jbZyinFodSgBOw9tWVO2WDo2lkhKyKUH25I
Y/luAArFOKRR+6JKNK+Ne2/rOFvpjyCPT1hE83EbOM6HhBg3NszrXa1LHhzHfaKvZz+W0RrSjEkv
nQsNRhPJp2BsNbARvJ1ikIHbOQNrPqIKAb8sRHVZXkpR3kbmgJNtpxwUWJXju56/utChPnc2Pt8y
G/8SCeU/6zDF5fOdHqYOI+nG7N6qNUk3y/EkUmo85kaIfvA6V7F903DX26KrqacEGFShrUdNqxmT
71Z5cnsP0SYkX9JjuRZGPqmQWf/PJ2ifm2TLDI7MqhbS8AF7qawXd2e9ID63D9rsMB20DkQ+PBVH
6ok1QHDTOvhXQU+lmbcHdmSMQ8CZ2h1+tY6dL+tfTMdlHK7x8EtvIZaMzDO0BWhnxvrB/A6dPCox
vUNupHdcmJ9T7cVhCUNL3qu+qqhuHvWqZ+M4PTQSbuSG2KyvL+s22zTbqNYEl1cHkpDdGoQTKFU7
U+xT0BYQQYT2rCM4EvvEc0i5yI8r4egThXFMvDFdFOjAz+4uK4mCsnB0gZb9AWbUzT6cbnCcNf1/
xRiQONdRWTMGH0cxhVgIqDbFLEd7oTbr446QSyyJKrQj07h6TQgFsXl99EKaDYNlwefkO7LtMBvm
C6kaEngdgcipPa3S5fpT5qJZFo2pbJhQG4IBhLvqbucjtspHdiOpCkQBDQ3JCyBBU/ZLa0MiBbaZ
suCS5dI0IcZ4ZrYF8+Kwxk7DGA8S8jL280/Th4+W+eVnV4YwfI1p7D8S2Xdz8qPEzGCPSIPU0Oak
H5uEALMkMiuKuw0Q2WCfS64SSjXRSPUt/GKbVQiRZwqsUNxgMExFusFPjD7RPABLByOvHD0IEmBk
+Ho0bdnL6NHGnqdetwRVCpIu0uQxwA9zach9zkUmhSOggRgQuoMwQYkk7+QQzH82W8TD2nfQyOIM
VWERloJP/3yREv0d3iYPA2ndj2Irm3vh5YrMnolz+/4qo42Vkn8ACg+JnwskpxZn7YEAErLb3v+v
f74C/Xu5ymJdRN8bawDwQCn05Jdo5qga/Q05BSp2ijtAMMWbDQHxkH0VS0ZvkMGNq4AAXxyhWjY/
ldayOYSQSJ2uUXRqUD8OP94IHDyxCSgXOrq2lpiXPInMvExoeMso25obwKJ8j7zmwEQtNKr2jY12
7eyTHQrlqRIvZsrevG9lKeG/NxZFsAprlzP68NtAl+V1Dd82GrHChppaj5m8fswzFUO1+9ZyA/au
cyFK+PwIReWVY0vRbYVWqapS4zlZTL6xFxaCZs3QROZVFKLGZTkJETsPZPB8r5tvCGcX0Y0ZEqIe
50hvgiDUEBg8uQIYX4k8h3f/MOcfs5DViXeq8WowYNJjOGj1m48FMrx1HCgyU1h0INmHzQPsFtEx
0Y1boDh284d9POYSI9QdtZaSBBYNopXz2EhQNMjQOkNPNIo4+LVgj8NWpN2NvtNtjjYPf58pMxEA
/Ocq19RM6IYEar1HilkH3u2LubVozCMxhTpjLVbwIKsL+q2Zeb8L609UyICdlZNlvGmaRdR/AlOd
GdAKKTn2lsYdnLAHvERqS+N43jJsLLkRYJGrgaXvPotmhwnt4LtFA2F6XWpdR/1/a7hHY4NGYD+V
yO5CnB3B2A7RhnXIyr59yXi32Rnv5/XAawm/qsclMYDCVyGADsQtMZJop7veyEaSbuZjD0rV8vJN
6mme7T1FAvUy/5X9QzK+SiPsdYWIAH8S8bTkFqm/E7mPUzCrQ8GrbqHKf3TMHNy9iqiV+SZ+dKcr
o1FTCYc+4YNRi8OTDynVe3LN3Kx1V+XTlZSlruXyjFiPWRfulSF7AGeTJJ/ZXYj2sGNOVx6MTEqy
j1c0As9HAUIUk9MTVcgpZ3ZON9UHBFwmAA12P/gw061u2TfzcV6YzxXanV2t0h3DgPlKvQGqXat0
JYq9GRRr6jspskusbf1kPrewGajZz4EEuIZb97K4O6BpD3xTelKV6rfOFLbBXO/tpBZcoQkTBWHe
HzXWmf1+h86aDFn/PAIrONnWGglZ1XWuFAlg02vaPgDgZsFi+CVzIrORn4e4lyH6GXTIMZ/KyJFh
4hH5+UrJTq69nk/LCx2RTrcOyZTelpOS2JU0ni4EYs8vzMmZ2j2FgDbVHrex/nX+1TS0c8woR041
uf1XMoH22W1aFf9+orDwCBjUbarXI8ZJG6yKtW571A+IaVl0HWJC3nnvMvjYZT36WAHEoGY/QtY/
N0G7R1+Gpy3J5nRABMldjwKIRCdaXKsMrAGl89kak/Q0aVYEAIDdxsYtxKA1yqMHIBTJ+kanjaFh
+jxCgq3ZTc1fkT6Rb2KQAZQyhWP7OuBoPTzrhfEcDUpOx/16y293Y7jTjBMIWJA8pOjlE2DB5mf+
dJ1TenWoP+YA2zfAjXJZmq3cGcfjVlPbIaLtD69ItRKcn+lKP7CDDV/bhAcADM7rX9tQ7sdOuHmk
wwJ16Rm6ReKseSdlo6koNxUUYOMWDUIRcFxxxnb/5eX/pQsBv7ksX28/0NXiCNvHm8Y3AysRevhu
oKGI5u3JtwFL2zklYci0YUNLtmA8QbdtANni1IXtfTbdB+s1w6KmgbzRJ2VyIa1nq2WFLKInyWnS
sho3sfQgrh1XpzM7uKjMAqeIAXuv0AVjceHfs/buTIS8gZY98lw5VEg3dxLvtiTFm+zdmTZ7InnM
YbvZJeWvWWeo/gVzdQYCHP1rgK+J2hJEuVy5+0HeGVbqYLoGFss9IWiwpbprJupns+bzpXOJPOpf
5i0SM74VBh3+QyAuvaffe+dpfgjBjVTGHcB2hkCJ2ZMVVStCmRgo1AzRIPcrz09ZVsIpAxBXdRxt
OSQxvxFdhBlO1+8fHR36BXYaHZ/+yNLTp4EIyd74CdNgwXmJ++EARD5vw/ibqYYL1z2jD3CRK2lH
4T7gWpnVKvEQ3FtRR6rny1Cq+qIAEr7IQVne2VcbqT4CoNKZsO9Ze9MnRWRwv1ZiVoKLzMKLuXOi
t6to7uCc9pSPqSz8u/Yi0X4q4ahNsVbsBMO2SsyZz5HyDKIEIqjphTSMUvEfvDsRth62xQTOqyPJ
pVEZYpepgC93YKHgPGvWZUZQAo0sQcbo8QZWyTHlAtzGEyyFcsl+FUDd197dn1m5wxAVESyuSeTC
ehMMOBu+Fc6wM1kxUrZ+TuziK0A/BQ1l7ateAGAaPj7MdF9PNk2u7jehVrHUqM0mtotKxSuRNPRC
L5Pa63Xq7chefuVNV7TqJDh7+M98Y44UGOoXb2LjSs4rAV6Q2m0otY88vfnFmnV+11k6YOVdP8f9
UldV7kkCAoVkn91OCyeQNmztK8KK3XT9kxyBKVEY7i7f+0g3yuxjAQFC+GQoEb5nq/Wo0zG+LTli
9zIxKXgkenO4uA==
`pragma protect end_protected
