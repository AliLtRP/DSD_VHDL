// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
mWVOMHWUX6TBtGc8ACAe4w2LivriyCeBzl2EECcvx5SGO3TjXXm8bT+UXDGlM1E/Uhk/s0h0YHj/
V92jg1ugUcv81a8SntQSbom1JvS1rISyl+iqEgPH7lj5ZCpLtPCqRc5m5tt6Y1vQyygX7U5ONvbW
q98X9lt42CimA4xENYF+2cZ3BZLkp+ntuoKb5OnRPhfznc/EhcNQGxOqD4EodYHsMOGqRfhkpnjt
dyVw//WHUfSOAs9G+WcKwNVPvIEd1OYCYk1BSEL5duJ8awBMhU3DqQp68rZ5fS9BJ+xacA+yY6dA
c48h5gsYCdXF+e4r0eq75I0WaYnuDq2LG80YYw==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
BMH7LebBtBqT6og0KFbDRJzojwVOr1W6DOuw/ApU8DOzP0TugbgGKkvN7Aj1IBxW3nEFE3uYWE7F
9fcWrlu2X54E3lTFHTijMtA9Hz7pOFt8prkF+MTSNtKewj684ba7ezYV82lh2S82DXEVGCrc+MWA
AxJFQV0sL3yUA6Jqz2WEmWeE3K9Zcn3324yiUvxLMHDhWCLTIGI4rYKnIIZEW9rJk8mfe/bmTPQw
28WPBVmHdoBAc70XDaQmDNZFDlz39k2xHlXhHANkw5+k4HjA3+4LZD+HhCWjVhy1ctEk1J+dA4tb
rO9D4OoEsmGYRwqLSt0GXe1rRJO+WxAqdj/kKSqZASC5oTwabZBHT9w5BF3v/qCqEIvbpjxLH+4w
Z8wFzKjvi8eA+ybeLjiGxhTpP6Z3HHLxZGpg0cIn7jMNOMjRdjx0p6nvzzGw5zf9CMK15eXsj8p/
Tvhx+m0emIv6sh7QzdIzhX59Sj0mcGYfMSomechJo5+CItOtRrJZmrE6L0SpBx90chnFpmNbyL5a
LWK5nZFarH7xR6mJRuk1bbM088eie0oOzLOTZyS0QSGZZEnnLO9RNi66Rhsv/2EJTNxWgog4lG1V
Sn7kIlwKK7g3IsSKVSYwuxcmf+JIYrEjCVTamBrSLcNpefmO2WFXWSmcIu79zshD9eKGFi70Dg5Z
ZQAryx/mNiQNdJnk5QARSyI6A2zsOPO33pqqw8LSHdHQ5rqhzWt8TTHR/yVeWHRp0nc3FXquyGQ5
eaeZySgtCjs/38tPWcIX5p6hkR3jIGm3ieob+lTELdt4bFTH28fjeQgbNTOfNouc5k5ga3s12w6q
wUJbIigcHosbLt8RoatcCMhBiEOfl6eiYi5R8WnESVfiJ9t0uSGeX1IqPxTNXqVFrSetEesQjpWP
tHyc0czy39CH8xG9S2nodpJVFEfpi+7pAVGk7OmGgKroUqQ7C9JUNgG035YR7BC8JQ/2JI8Nt4Il
8s+yItYUNIdHN6+sf3+pir8jaaAB3TmfMc4SD4irg3cJlyHoMx7FbqJr0cxClNCQm2w75mJKyG/2
+NbF6y6h8iE9Xc2cpciZlKLt+4NnnFXTf0qUvp0WLvA8xCOMHpOsOYKFAHFFG1rUKbdH6bG2eLJ8
8FY3Gah1CEc3Gl1XCavHujGsPzetgJD9WG1CPz2EFhxWYu9w7LxLfLgYjxa1RURW3AnYGvztzYb9
JY5OM6ET/5Gxlpyp/OdFIbBrpB8mZt3AVawCavZIMweWXnP1pbaj+WUP84QFFTjZoyGaM1+mQcrO
XQDvO7oK6yTdy4/10W3ja8NNT0RatmHQ2HDuNtI9EyyGZ86wYEGu+dD7kxTIFsQTsMrlEStOGj/K
HiKpsrGMeFZQKvJ3306AC5LbzUiHjlJMM4MVNFUH1IWKO4Bg0Uk61QWOiH8ELkyR7F6JNPHxvwXH
qm2YXDO+vVb/FDAzuHpvY6rfkmEDQTuPD7jRCn+N3PPrYphq2pejGdC5mJo1cgEwaDnaLIRqd5EG
1edfQ+TORbwtUrnlM5RO7xZiH5hoUTmUDUnn0Z8u4EMsycFQPEgm1g5+zJDxKKpLFJwsVl6I7XKY
Nsqq8pCLfjdJTH8rOBLRAsrVPWHIUOE6QSHWeeVuM2z8q6RMRuisVPgHjvhIMXif1CUqr/f/ok0I
oEcCenwHrS1LwbsTSn82xMg8nhQA91gAB4yp+kk3itdg6Ao25tb2ZzQI1gwdjn2/GmyyQiKz2qYf
PNiAiyN8faIpGuSbzgtKvm6zDDr7nAebXyS/6wyNjBeJ8TBBpTtparHIOSiEgnin1HDS8R34Hzs3
cWZSuQvoFedv+bwk7snykb+ZDKFdqpx8PSgkOSIC+FHo5fHEUTznJrpwjjdcU5rkwHDN8TNGQEq1
69GSKINGnIOVZzPIoljtDPrKjfLcVPVVzLHMxMRH1we6pe3S8s+D0jxz/IrOvai1JXN1w5O//7by
cn+ezq3B/SADKn8V2a0EMU7BOpCgp130+lfMqsujTlNwnYXCj1lGMCa8yI6W7O3EqoX+U6fRBBqY
Q+8PHmTotT81mcByB1B+qf0YVvXhBLZ9WCLctfRKzeh680lYQ83FkHIdU9zIEkvdePa5BN6S2p+6
lvgG1YROpolO41eUYQeoI1Gt2ebP7X0ZjWZ8eO2b75h7nPdedrDt+9sd9aX3cvOJZCDYFpjmVa4R
KXakVhpc99Sn5IA5FE94fQcQUKQNZ0R1fACr6wlGjYLxV9Agr8N4SR3vxQEQn0mKCkhpHrcMot05
vwqP8qbdLbPNptmz8TPE0erdHZndsMJ+9sjStw61dUzLlYsJSdy382W+iP3ScFWXqCLzAFkjFkFH
7T2eIX+HI6Oua39Y8UKn+FQgdeUEgwi4j1oaCoG+A3fCNQMQXoIuSpEy783Vh+00iIVEBmy6VJzo
4FTh270CE2D+YPRrsHViWylo3+IyBKlWecM1lFafIctLIdjf7wuxZL7MRnU1yQyL9grF9TgbgrSI
QZi4GCW3vXo/9Tu2hhipqDKKcQ/bOKnEQbtUUPcE4n31ovvIsNM1Pd0GVV//SNBktnzFT4a6GROz
iOCS/uUH1h3R+OH2PBiMVlFTuLU3x28C+1z6XPh8OP0/oEd4hySe/kbYrUlOODE0dtMStjsZ0o0c
97avOwr0kTQPgFfZch0gDHeGGBbUsnTrfwQP7wDHMNXeQvi1xgRGwU2wSjlrmeyOcwWTIQHaQ0ft
bgCRtlgOKV2uxnch+JntG6XvPxyQjzF9l7HLdXLSVVbQxfftvDXv9MCvr5ha85u6ANueVfB+EzQL
Si8ZxFjeO6C1+Mp/BtAPNQAlSfALTVZxX5yX2n9XUyH4iAnenJenEW8+EdyBrTnWLYObqJ4qgHRU
ihdjFvG0UGuOwfoL0lnhQ2af0A9wKULGGFKefl/o+N9WhIWtTunRhddrUJYZFkLs8xlX+Hbo5BrO
Gg4YgKEC136Od+OCNk4f3tblq+J+7WUIHpZoKeBCPDHovxbFJhw6wW6QTssfXTj8wUptUaOlyxBC
XlvYClw7eAVWPUgpRGrVoSIo7LlMR9EUAYI8N83ljZ7PgynwlWSEFzpvBo7NlyWD7Hes/BHlSZjy
EmPrUg/Pd4oUy1WxkbN6OE3ssxFsvol4VY1VH127+egL3fM0kqnzgmTl2BbOqqd+mTfLX6KprvwE
1TbbDyLCVnmSMERx09H2SUccgmfNwIIcJgg+PPxAEmGhDt3CZMtc4DKFLnTtKnuNvWce9I+84a3u
oPOc0Gh3Ae3B1f41KulE8qqQGdJzJlFL7rIM/yuOiOVMeqtEeyNv4JsUULXgQQy585DRWl5q5FnG
lgjE/gvIPGxd8bWa6o+zr8cnZDG6GY9sVfHEttEaf0cfaXvI5LfhP1O3l1t/dfOSbcUMtxAtxzaJ
PwNhs7bSSAYCRYOpjwbHaF4zUQYg6TT6m8kelpfLy6tXsvSES952jeTxfexrOhoOwAfMB3UBY9xd
kQDO74hVaYuro7GZSq9Ik52gfxK9MP84D4cBFFr8+YkQzhb5t6mT43Us/RBgzcshcVRXONzNuRZL
jLcRV77yxgvQeZKVK4aOMVtR3E5qB74SWD73JbHb6aXteT1/pEcUkvWR5YJ5FBvw5VpZQchNtDQR
vg3bNyelajdE7hi7kUopj8siHZSFqC7G5C3vOk4SE7NyHlhi4J1p4K5xie54AdFKcw+20m0FXw6i
vZCH3IKHeGn3yP/0j9/YbhBKWJHKR84GctuEgIVLR6D0yLuuXGU/kEv2XXKVAC/0XHLaQONLs8DA
9665a7VaRdIiiNK8tL0q0PUq/VQg2qrdxcefbAQBAcPtA5Ykbe0MtiLdzOT9vcUQ9SVUykgcAzha
fconeyKGxwdTgacQa7rE2SBcL1VwrM/mM98hCY+U5+G1nkhXZPOOyE/+Uvo7wzpo3f1zG100F+A+
WglCFw7W+qJC1O8qVZThFEfbwyiYfORuDG/+i3MITqyFnRcri6v5GpTf+lZ/uEoCO046NYNGTmgg
Zj7BMX1jx0WNHQzenNIRrXd3no1UVUGMpynskpoNu3UQR3+vOQz2hZ7NN8pGBnE9oGNQltU3cbec
nQ/RPRVlWkRrL6yVVWMkD3N5w/EhgAecxtySaEju+8kG9w2Dg8yLV++6Lv/Lm2KVA0opMXbG09Q9
TfKBuuMOULK8Gk+rW95cu1SemCLwiXsydRfCwzP6eD67jRSfO9MApusi+oGODynUzSdx2pztPz++
P/r7NWArSWu1rXn7DN5Rejrcwct2wltB4PGMFHYsDYs2xDQfZQTJEdp1pUcPG+4Hed8vdBvIhhhU
TXqEn6J7ZiyTQJWj/a9DElgmXrZKLe+X7yXpDWOSBPsxjWY3Txv6iYHQIrOoV+drpRWt7WowLdfN
wRWbCVwg5+Yb8CC4BZM9OyXj1nbGHRR1iIVH22UNEJJ8U+Mym9iytkDJ/IZi6o1d0nzlBWQ69Trg
8E+53H4SWpXSTaAgGsrpQ7jyDHPgi83qcODDySJLMf6NqZuGiwlWnGWhCKauC/a6DHhpTBaZVhEb
9uCM/hrG5lUPI8U270bDnL58A/FYAHm2i/m3sza8pLlkMIClj7KkAdxCGvQ17vgByP4chA8hoeX2
6DMUDG0g2/REdadkFg+WaVxc+QebZeI7V/HNE4yW2l8TLZoK4qF3vQrTFu7/30T4uJtjgbP2zi4e
jBUeE+7gx795SSXxygKm708MtUqEKRIzOK+8fw4QrJxYXFBMlizD1wWKdBK4YB8G8fD5ndr9GQYf
VJYhLNY+kxSZjd3Pc9BPf2rK5jZwhX3DnabRMgvXSKqEClBhdAURboV8Lh0+2qAlZALuJvYPJ1jY
DYzqRazC4CeSeOizHIyzVycm/2csWbxygq5oCJ02dSnRgXwJP0wcwWMD78uDx5m21a35JEcN5CTH
cnvblMKFyJDmQNMfJrXkKOV/LaN5FJvQN20Ys2Ih2XbCAdkdlvuWiDtd3ZAsBlyiygq0bDiMhOB/
qRGKoAG2q5gleaw1O67Pre+TxK/vTusagfxejJWFVffYwv9Q0zAuPBSQO7wck5FO0HlCIEOFQFFx
fCdoMAFi3b5cPdOvKfDkJb2I+AlNERiZOc/yVl5mBZCgFm706t8wBlqxXzU+IJ+USlDEfn1xx7QO
ylzR4UG2mJSUu1HaBhoCpPLK/tBBtN2FfmqFtTKrUjRyLaCI3KtHNMwyjzxpe08ivGVeyH6PZ60r
jpBuawnx2XrKHcqrMfYu/ICe8Zzne1e2QKZ7QQTgjIVPbGTsTB0O3rguC5Kv2It+GZ++KnAgW4jz
4Qaz8QxvJdlT0Aa5iH9rKKrBj9oHtaeEYztfbZi0RQmj9TRde6xB+5d5nU6V/NplXIZEIHAcfmY8
9AOMuF07+LJfJela2y3rFc8+J3ochYj4ZOi9O4tO1RTpFr5i8t5fYpGuErVY1sP7b41iT4NqAul2
64dOZG58U5txlK9RCLAzSJebxLYdsMcyfrpHHXZZ0wqCfgAv3+jcHIVn0Bq7hSZHAGRrlqFcZRXN
Guxupce20BiPL3/b5ZZ3BpgbAGqRJLKKS4/iHieu9U0Uv8D2U0XvlNi9luBJI+/clnMdhBd/ia5R
YHDJAc3+RCjeHrYMoCCMe8X1wmPPM7spetGIyiwgiydyeM+u/YNydK+skBu5uAeZ/KvmY0vCyOdq
s/rLfqMaTM/zhTGUIc2SYkc3DGiKJD8ha9IgiYOmW9okDSKJVdJ8E3qNN6S7PDovXbuOX/px9Hl2
vC1T+L6MbVmdepyp06qHfQWI3xMlblJ+8Djokc47tZilOQzHwd4ROal9JmaBlve75OZfCQlu+vAk
JnUz26HNssyoUAzopaAkli5GPc7zRnaoASv65ZLOzOo9EdhkxzcrSIj7o5OTQ6AJYZ5DFs0dz8IR
O5II4iBPXxN6A3AvMF3Hff97YdTuIQvszQO5j/RpU1W+kZZNeW/NQi5cEvwP+C9MCBok8O9j8VIE
y97wWo5wTcTms7Z4oNJ8Bj5hb3wNcyb5b0mzr3cRKOvlTg/QAWoRQeLu5mj4HHgd5u7tjFvmTS28
8/jjn6MplFWzxcaGtdXKlAke49+w5TL1wdZTL6EYSkorDEQyNXF5EnYPbDEs3UveqpdCvyQmhkCO
WuMfKC9vyhn7533x9MniUZidEVyVBAdpdRbHeribJj1OWVmwVYChHR2L+QOpHgVU4H5jTlfI1SZW
CciqMbbNA5P2xltYzDfPoraPZ5iQBjaBYyNxnwosN84ONwRMe/fwF0l95CV4WFrzEGp24hv/2/NK
YjR67AZuGAO5PCZMB23vFValCRrmSko0MXxjtE7ylAh3r7eeB3x/CWsAmKtYm6sVdoczwT+5r+aM
tfCffRApRYmKDXiiFiT+4zaj779xF56EkIgzVAhgglOdcutpjfEaK52RfUAQj7Jp7Ym7REs5mOk9
3AaFljZrWmaXHOnNWPN3djlgK83etkGMAO9p3haVgAB0mxoyrzxBnsmVurkGno8MPcCgaXAhivdF
g+r1fgQVsRdCvURcKCqhvVpunAOnEwqI+CRLlTZ4zKfLMyA3Tzh5vMLmNd6m5S47WhSVBx0oGz9i
KXQbWquda5Hcw1OBu0x3D/eJ8KcH0JJii+mrfdJa+KoIo6ISb7ifwqY578T9AhnRuEhqXlHAJDSB
POe1yzXSkevUmtyn0r7K5vtsvMSUjp/c1FOwBR1AlnJiPvbp0lUM9sD+Qg4OPhfE52Yg3HI0Osvy
JHQ0BmrEXeBtODmlbDz3/fjybDaCACKN9sZP8ysvdRn5Ai7DPMHbJqfm5ebrNBkomTdDKemUQPVP
j+vh7SY1ST35vlt/XvR0RDgpVax3vfF89WE75sXJjki9ZZ4GVQzKPDp973shuaOuPOLPw/4uaS4Q
bTY+QResBaquPuinfqQWaIGyvYX7FkAWnd8tinageoLfDfBf8i61lsKEl5C57+qnYJu3HcphaAaT
2prG+4TDA6rD7/OOKtt0WhTF8nayD8GRAoEB/yWmnMW1DBUKh4Feks5xhW5amx9WoEJSt2MDyWiR
5X6O50fZ1YLr9fLWJrP4ldjBlGFqKJy9O8t2zWBJsvDjy/ooXD9WLMB6vPhqe8fPUDUNX5QsdtgY
4Gb8MGpoz+WPVAezsDoY8kSJK4b/LJzMwAMhU5bZQsKfKhjgXjG0NzBuH9iRvIjDocXzTBSKxI2U
SlKHgE1agQ2LR2GAuNmXulkW8jPuXOZ53xNiFLgcDmq1dURwcnD8HCTSyfl0ZkdVoSwp5mNI7uB1
SDvffokLRg4BBIi2RTcDUavxofflUEPkaw9dUrOiVKLWybX3e9Q2XtYl4vc406xmm9iVakrQYOae
V2+bq78tgHeuldinzd+FzHyVzv5BOh/0khvcR7/ZoydQj20TJ4Ih4X4z500XBW7SeqatjUQ92BFb
0Dcj06EBk8UimNJevkXkutqBTqIlysG5hIEevFAXcP/H4okCSK67ZNZynAUlMz479FUB1LVsEOJ1
lMeOgcchPaioHu7EgBmXdOfFDlfdyyDzQHvZZGeUQDr/ggrch+yTC8WVh2zEeSYGAU5EyqtOlIFi
/jw7UTmMpgb0IE6ctKzzZMUFnWE7SSXJjNcCzSMDDhLAcRRi0RDpVaM0nQFsjr6kJxzgzhzVsk9B
d2fmw1RepLOn875IujBJ+Szi0pqoYnl1S2T4EarZVdmz6sZDObYxvCwWILGxK3qN5BLP6Kg3aJro
q1+W6ubkFNTsHA7MfnbxQU2cfhZNeMYgkkj31qkT5Yex6M/lqBjKiuiws89LQ1tBvFHisDqU+VfF
p88XvBT0nbzwLiKBcFGoAEWUHtAZBPsR1KfxORvIC2hyKfniVYgUMBWByf2CBRZCG2dRqoM2zqta
l94u2EOju+M1ODhz47Gm/n48h1wpLzfKzASDgbxmnkdpUeFRBQ7oZXK5FD4zTuX7vManFefe/Y75
KmGKiv9dijuC2mjLy4JUwaTkpUL8kodJbSLQlEa5crwf6MMmIQTc+mmxAtM5gyBaYjdVZYsWRDwU
OkOEfFK6661dHHUNOm0tdpHWdF+uDBxx7C0LG3HwJunKgNgMhjU12Z+2eRtP/69ZOPbmiVgB7RQm
meyj4fmabbs5pvdlWHVGFHvMCc5HS5/Npt6r29jJye8ptlA4qY9E99ivKp0SNSneqLvYQx75gYdL
wVjB7elOZ1kyef+KFF+0rueFFAUZ1ti55Xc2ZzADkwg44JgrtJ2Zuh+Egcemml5hllJkQCyy2rmD
7bMpk3XxVFJNtVcbCcO8PUYaydxTa9PlibwT7KlmJNmw6L149EKqb2m6friTZ7JJdncVsKmb35kw
VvSHv7ibuHI6DT4wv4Jsp6SO6ppbgmi56IPWaafd9s2h+juSMoBASctjhJno4m0RuxbKBB+GnoAr
g9qoPp5KoT0XuTVvNCIqNivyOFpVkv9C51HbmP4LOJKFMAbEsOENY5uPC4W16Yl9yR39AqSguhAh
+f8Q+P1qYzUcDoRmGanQjpRilXs7rdaK25Jr1P36+J34zULGKO9qmadaI3IjCL1rL7jWGiPYWlbX
C9VpebCdnoBe/sKM1oSScpVzt6SgEcY/DEOSwl5KZZTDQghlzmvHytlwefJ1/OKBrpN8DLKVyjXM
UoEchODqFwjEbSlQXGKMn8zABvWjOXNY3FOEW9XbulDpsm5oJ2J01PbadMVggC9of6UhwTIQx9EC
jUt82oxpLSLAipzkU7jJQfTObKuC2Oi+t9s7YQ5753DaVNoLvNyk7OWsBPXwUQgVl616GWnUkNsG
Yw8nUjh7wxCV8YJoOEeeAlLTgZfZZVQ3/UJ1ZKTruRdbAHq/ge5GrsJ+YzDHchX1hAfB71w7JLSq
NuOrEnLhmFATCcwl3Lv5gXXAvy2DefaJyetcNLmjOCuivF/v3ud2mD6qeBHkg6pHYFRKrJXkzeTL
ZE4g0X8+tUtZqjmauy4VXVQpbEqWxixHjNGqzz5Qn69stpvp62ZfEvFf7AStPeisFphF0imLtlTK
P4uRh4BHR19EbvJdv/XJCQiWi/UDgpCxWf7wFWNQPw4yy56I7tw1uLoFBdtpqQYxSuFhgwdYvC3Z
RrohgPEhdoJIUeaev9SC/SbxYlqjtY+Id1TBjFhc4NDYD13WgNPdpn4ZSMr6eLbXNzmX2gZjENHs
IINHYgCPAZ3JilPKHhWwx2X4J4xDinq0XgQtinM4hlboouMSqphKH6oPXqozgd3RcwpeIVKXxerK
wCe+/YF0B3aEv1UXbJZrNlku60Bu0II2UnlAZNTu2sbfgggbbnwZKzVD/1pnjQWGTdOMdPCDMaW3
BN5qhifo7EFBEXNr6gctmfZiU54IWLvNY/YfHAzyD8o+rokL/yQYddrPnC/MT2D4p9zb9al7pjdB
dUScqgThaOOuLMXrrZf2CHSI1XbPqOWntKiGaOZzu5lhPjRO7RLAC09gxafxIgafbS/Lg0T3IkdI
6Nx8EPy8/Go2gAiMwbVnEzobY+wser3D5jBCREi4MLnE0aqPwgdrmzYapErzhj3sAIHxGr6RFnl/
X3JoFXEgbDgTg0gItkGDcBaCOUer9PPpxo+Gue8FgCbObx+wWbhvr8VimjCBj5wtv8MG/pZj2fNe
QPKzIwsIWY+lVy8+a+izZXwSCZS8tl5nMDAbwAK1mnmjC97GM72iAyfSyfMRGKh7u+ktaejjKZzX
30IQWzBGeIKbtXS6lql96ABQBMfORQNPR9ZMqv55VBeNiQ6GeXd9QENk2JDpn6wuzqJFXmnQYWjZ
AXeZssdqP1oFUETRGl1OdS/FNN0b0RMryixQPr/nUsqhEkEUdBZushit+rZ0XrQCqoMnI2ZOw1Ie
566k5BSy5yEtIA/tVwZ5SsN1tGrFUGMBTH8CitGAoP8nKi0RCZfaOByZpNqnLGFAb5vsKYeuetao
dmbf6qfno26qMrA0mv8wkPhLwSJjr/GcaOzrj9ZUshdu10HmZIp/EPrGW80lyMPX6/9H+7GRfQ8C
JRKk2yWQ0MItqx6Zuh30IwYCPRRar5RAcp7nblD0H3Whemu/pvu6VRtIOy9I7hkAVhXFgn3qxj2t
mzuNH+7QMaqOMoElFsoIycCbNadnipCMeNFOvuFNib+mdzSlw8FOiqjuB9fc7A/lcqpL2aoNN3e3
cNXDSg6qfFrpulmmOef0FiylXga0EbDZ9CAXNCenULwpytFlBWSJINtUTHjQILHICXyJVE21ANeZ
740PmDe5N4bxq0+1MCpIL05sU5Csjf9utK0v1U3WOrh3PN38FfuO/IGFBIcP3N1JJnQmiEMZesPi
pxHG07gk8CpTVATuiFct7k4rhdW4qgPqzJJ7jjLGs/bRzCI8Q92K56YP+Fe7gJ1DZ4gyjS/NGyAQ
LAmP8kbfX9FdWjon2BxllJ4hl3p2QzcKueamuYibMzjTTokvGxx8b7s3ssbg4OWfK5EKAWb0ClgZ
uRCUz8tqUN/I9Ds+j439fYGGk+mRBYJsSJXRw703gLBgnzamMkufPVw/b6XIQphv5vjot9LzaSbv
cdfm2fBMd8t1vJ5wYZhRejPDUghQReuOavR/jrBWMVQY1lgswzHx9lC/8gsUepuphem4x6CiM0ot
3dh9htP/sySjiCLDByvxXUIcsab90kFnUQcv5FP46A+aDbgejbIKm4o+GDAxw2oh0P5J/Zcd81Ka
igi6B1zBqZ1Bz6NJnWjLI04TGDfJ6jmlQ3uh+Te6VlCb0OsZJDWERipBOKq0Ci95cT4Pg4ooxFHP
OrCHyOBmR3FUB47cuR/Sf0leYD0arLk2s+XqnS/IjOt6aCJvbgzfXGejPfTUiI7KexDv3QYONNJE
E1/INsG1brauLqbnbvW4j6AdcVPeOY7wFFFemGbfqg7bKLzMqs+nYnq1X9I3m1Z1GUHoWZi799wO
YdiUOe/G4NZ6avRHd2F4FrKE3Uylsc+JNfo10DgQc3oNgKlNmXo4F2cYAVOpIp0TlOdeeL7IfG4g
upE0BgtBfMR1G9uz1TNoNPK6+6PX2SXsc17xn0bJWorINxgDPtbjYomdRTswwjFXTmkmK7VSBFSJ
NgdReK8JYh/45+nLMx3N31YCaPowfLB7LstLbzzFYKHT76mXEcTs9ohWVTqtSBuUwOnx3ifQSki7
WPxW3guFxEZjfYefxBYC8uVJnf7kHaQ6R9CatTIWNTcwv0DlYGfqEeT18RZhxR3wWneZA8GjueZF
wvnxCq4ZqIVwFKKNysqz38NWio/s6Lgb9nbi4o2/Fz8zzTiILwfTI04p1nmt+gn0qTe5Z86KkQcC
pxDDakEczeGBXUDwCJK+CLajtsCFkDLBfp/fPWlFkxiPGxhAZVwh0j9j4nf1IpedZPNSinbTHGJS
n9um6GVBZ0szTX3pr8MTR4A5MiOS90/9oozDbuykAjaXHXaLzKCnW8Yg63Ex+Iv8ytQkDJ67UZ9r
FZQYvGiezCPpnkYcfQWvIHCCCOkW3XvHuSN7fdx2Fx+BH/cCMmqbegwymhZ8HT/jTUUdA5a6JF8H
x6YybzXDcbjXrnOK/yhPcD67T5SG+1USOeCtC72qTXz5Gh246tvfh17rP6dVHF0SEb0tqqKFaCPl
zNGIEzqLtNRldBxGWThcl94GhOT1tc9RPovFhI7VB8GorSlyyx8G5zvcG3iOwDlUzKxEVVuu0nEx
gUkG186/0tHF6uarlsfTuEysF5o1zHuDRFyvpAYOAcSFWGr5OzkmV7K0lDNbPRIioEFf13YnbrFc
yn6ehJvyzFw1WoI5DO3CYXW267U7XK1OaDyG1pBByIJQRZf8gIL1uAEEsqL5xIN5ztPRVofeMYQI
5/o8BnzhtWJCDdD9aoidxpKpmhvshKcMqjX4njG+tiAXqCqB7qbTWEzjt0hJ7R9JplZOwqfQvzgu
n2cRTHP9YoUgmDjEedS7x99C0SGvT8rqqb/zJX+QzNFh3jGgzwThsCENLEscvXdQqFIizQd8R7bb
DwkAcUtJMg1qCL1IUdEZBTEqyxM4y5ty362inW3Hk6CjHgXCa/V0iEN16BOR/EfxShvOo6uc0EW2
byJoZ67Ib9O3K4Q6jVterFxiIfixfCPZD1bjZ+mFyJK/u2620GcW7UBLJvtkchUzjTZqdYPLXbA1
lf+bGx82N9056taSQ9e3OKfgQMMYw6RRVFA+7lMnfzUdy+2ABPXYQU14oht1sT6Xn2YDRu1hMtYC
H3YXsTs6aHWK+lEdNteZzTjyz2EjWlIX86BLcM/LNoV3RVjMNtkXQII//ZOU1dzCXklobftblHQ5
yqirZPEH7G0muBwQxYwMWoNY6gXk/sqoOQrVJ6FKWDYo1VDXHnoYPDEI5p2OcGBl3/Vbsjs/vDjS
RmVvQd/l8On6M8sQ/AO4JgW5DFfIACN0SDJL+jPFBuSWE79vm9E9RvObefVx2rUdTADj/jwMqbFn
lDxWz0OfkB/i3EHMV1w4/keelx8gxODk3xo/A2eDI9Y0ifwb8ODR/CQCdkLaF2I/PQSvkRjhitSW
1wleRXrCj9R87fw+OBKcH/Ck3Vz2V7TMm2ov9vwB67wHwNoDNIkx59p27iGXSbx6Jq/v3jf+sTNb
vak1Amw9CACuaWih+Lp+DDJcakIaI3tHtLsFEnZKA/oNr6bfgCjp06vnAs6YVAskheOg//+HsY1Z
TWYu3ZWD7s8Su8ICVX1qwJhRABGzjO2jTbMAEJ6a1S2FW4L3gYfir425QxHTaHD49UH3tIlFlQ3j
kxfA/Z8oZN2TWsm5mgOKTqI9wBW0Sa4f6+/0xHOMAWnzkjT7sMuY+N5f2zA48qsFH670roLAYUXz
uyhshkp5g1d8DT+9UdKauLdO3eMtueync1KxI0MbnHJd09tHbX4OEWRG6B6cDfJ+OOGIiJi+7XFI
RfVjD0Cg/o3yhYDONzElaAtElGz4IWQmmw1YaKAdOxTw2b+nYzb6kFhXIZRk0emjMR07Be9GMKLZ
8Re2A0s7H4PYyqFcYKTwQGSJO+it0snHSAXrGdjLefOpWvHtabb2iPsTY3KtkOC5mUr1M0l6Ln5q
J4pH1R3twurgDd0mjWjZkhlCNDem63YF3joyttFYoWqNb+6vPp6o3KfHtXu6W+MtiWHfWRkPU3Qw
+3RCLyVVCcktUE6KLf9Ei6h1bU3wzCi7CGTdeJEDS7gOEXUkrTdEHiOIPSmETF566B8nUFfUNSWy
tyQdECn2rRRMe2P6UPTuss2D2toIYznPn5qz+peIjb2l8Y5Vi4STVNTg6SHCfx7BuBqSxCgQJ4pr
NKZao13iMj+62GjS2ozTAgw4vU1zsmHGPKgpaGO4lynAZrq+RW4XhLHz4iJGiU7Mi6ZApe5sJPuo
8867ZMq5b6oYFmOlzDzctyWv5hNwztGFrXmgqp5puZLmlkGBHbuaiUh7FGlqYjAucIXxT/+JVzwK
2qwBVzWnYqD7hZqX/q8YX6ct0DCEoNg68+zoP21f59Tf0CFrwzp4DfNuRPMTINWUhmUvOP8+Q0He
Kt+SJzfzdHK6ubr4afjWQfOGqp7STdyhy/v2FQqTkFgUdhpYADdtQuMd7RUMgHydBpFu7SS0dwMr
qaq/MmBxxCJ7hnd3UftAS7LFS67/NivNZjXQ4ys0yKJdOOjVrx2FjMNzuqCWopPQF56ZoDgWfd8F
YUxDl7JYzYL00kWEMhrXKpHhipmpa4+2Q0m4P4iSRaBrFI50JGd/zHSRh9gCvK7J2PjUHOK6e4pA
dnA8cVlE5n3Nv7quXeUXgMB/zDWujoL+MiRF6yiSsLyvBlmEE/SYBOCi/qoQa/O8XqlxdU7wj8/S
/rwxYjGC5jCGaf0PAW9XPQbJyETdIdkMltevSuXsb7b0vdUE08GiNJLq2x82lOyLEyqtSmxAcj77
s24gcl4JCU2IqvJCA/ELUWVLrAqdmXhSk5bl6GZTDg0tsnu1Ye2UtyCOmrG/djQQiSdXb27qyvAq
9Ihy+e9d73sPebQkno+7yHBU3CwJOZyQ3++fBmR0sieCT4bxivSUocV6JkL/8jrC4Ldnzvsgbmyd
I5DGpnNXl7yWhux4eIncWj58bqgF/XHIFgHoe/QcQoDAEbFbDtxYVjVLk/N2pv7kaE6QdcHCQlnh
qQdxfDgmk4zXZjR+YMssCej05+5vBpYakp2wfRvNNXbdSRRwpkYv9zrfpsNEVovQ1zk681PWC4/H
DO/k5jFSB2iDO3CjyvdKCcvkiQEiC+2wGA/7f8H1hi2QlegQ9wkdzpwz6CziFe6RTpy5fj6n8JHd
MhfSVCwxwpHUgEmLl5/I2ZwEWQFXp8ahTENxvIxssMiTqK6kibKCyaXgzkNPqwRpVBUU2J28a3Gn
TeYhk5ysbINtFGQtjH2NHLKWN8utrvHm9n3F7rNDHG8FsnTJMjiBHiY/81AXilRXh8kHgvn3PNM5
89i7SYAkcQiiVSa7e2t90mMSrxJ+NQYYKqxRlQ0sKL+4YrTP/9/SW95F4ksATQRdvJ/+07RYN9V3
vOPI3cXY6t3Uw7uQKSyAfRvTAdKiKnAeiNy7klN504iGb6rFrfzF6ShnqIqdnlhygC1UKrfc25qS
W4A4jMvz66IlhH2ij5SVjXkmb/OCHwwwF+vGilhR8K2lZsWEHquK6YuTOSxROGSOR/plT/vRYlZx
cUCHQOV2AuS/2BHgPz3OeCT/+6x8Xk/70v/0XCfyp697Mo10x9RRyyn3hFV23IDkpTgjSviljVzd
F050z/11ZJ+m2MhJyiFWi+CwM3PdayHfoDANbiZX5Bbn8iSsX5d8nckzg8MAN+OpOQuslWR3TC8I
jhboJWQ5DbmWKPgzd1LrQieEN0rAPgi+9xqlUVZVuh+u77erATc45Yon6hnAQYGAMTbX9Q+g/tkL
M8p6leAyxPZs6FrZVbn1rK12Boovx0sUNRhcDhBesAmIbRpN+KWIUKevrdAIWMwTJ7AR16KbnF2X
PsqiVeqKbroJYVXw4q5on4LJHMMTaahtM/VwLtwqEIT3QC+MrhJfy/0uep6cVxIJ3o5tMQPxWMtE
XbLs17rpf0NVSxFlt3mv4w0ohtwo6bBuEERhTjgMNkFJYug+Xe/jJ76SsEUiRlDjgF8w02JykP2+
gz2bxJ9lgx8yYR4rgQ9faiZtaLyNt0qvOAMJ0M3xqug8B9lPlL+wtrMNuznxzn/vnzw9W1zRlapA
q8qzHwuv5H1feo1npPYkRaAOz4HWU8h3jn114wedK/hwmwgDvhFp0JMD0qt+V2CLkz8QmjzDgXT0
tavIUI0Pffo8ogq07pZyQcGKPH2jDZ4ZQyhV9QeD+R/QnbyKTSM4LN3OEHOlBXWVQ5DLxnISHk2/
pjITvGjoRjHZu+EMOolWCN3IpknVzkcEUoCQi9jpvKEaEaxGk01GM6nvf7L3JAObZIX3i7PxALh4
3dbbJFpiO3J3Wwnhpf1hXoVXNjVr7/TaYs8vw5Fqw/R7wWFtNntukvhI1FG43qsxcdEXHeZLBHAN
HcImCmsXFAZGsFsMsCrAsdFrCjjQsea69L8Q2j4FVX5Y5qwnivNRydxC4BLhp9S7Z7EVnU4B2QAK
IJbkvLT+BzRKj+8+Q+tOFDVBb4eV6ra6IK202C7YxDDYj0VlPQJB8Aqwm9Kj6kGkqOqqvcO063wA
bCYE9Id1cJ3j9Ouhlq0YbaX7Lv3Rgu3ODC45byiAVsS5S98ocsDg+dINVyW1fsnv+IFajLnPOL+w
mBiF154FJUnEsWhTIvuz8r4DlPL6E8Hl1PMUl+ErGRw6JbF8lFPLeaCv2pC2S6t/uoyobDeaLxKx
K0AIEYcDzSOCnrqPWrki3NCXWiofuRaq5G6v1PHZx5Z7A6PiV9L/b5JwtXZTib8hD/lcAX1lmQtp
tmppXeAE0oyWYOqtMqOriGMpTQfx2kVrQ5KitCcyF/TwvLJy9OV+U+fpZdvIBXPedgmWzcFNVOL7
wzfEAQx6HK2skMcu/NdnHK7ui3pcJxIAxFXHD/wKurlCt898RvXsV5SrnZ+49erX6wMQwCjViwpB
gjPjvlJOVSBhMhFcdaqULfXhRp30Gs4DvoMXv1qM8VK63JLK4/EDl4Kn5JCTCeAKMzLtKkEweJfi
TErkOiBPzUkodeAiJyuHvIKL/wuUeDuGTAchvZ8EdP5FrQgr4rH0ilZda73G53BDlx+3U2tS8ib2
59xQVAIK2rHcosgqfZqBgiHtsp7sgxRZW33YYJXVbBsNvTZ8/FgCqck2PnArBr9TfaQAaahEDo7/
fl/NOEO/LZepZIKC0nD5LDOFxhRT/Z/ADEQSG0yOpgnXMhElX37JMwn3w1dAfggDVAiWCfrqZ+DS
HqDVdDQaDJGTAwyfyGP9YBNR1AKg69dKCcqw6zKy1kUlapVmKBbk/quXQfX9KQmmfcu0CEdCupO5
W67dwd1eOjA9arfSrVzUc7ScNOZLoF80a6MkQvBsYKTztOXnnH1bDt6YdsblegylPUuHUgbGAWfT
V4FppftukYc6yZeK7U3HskgklXPcpMzPO+HMvVFWlR76Aj8lX1lO8VdmY6ymg4fBDBfgO1KkbFxz
eO6T7Bzf35Y2llXK0/DthU7SNhNi1NMFj5fusJBYVgVwJAWDcTigvykEYU5afklH+a0ghBg46R7V
u/QCeZnxJkpfZRBevHVxjKHJdwvAKNq2PQbksfl80rOiElMFojmpXilYwA90dmDmpZCnL42XjFcV
vPeS3aiFUY9PCRpo7i1WNdQ8yeGpg8HyuGxJn7t8VtGrACT4mayTqbnMkJJMOd2kaN9EBdoX0Auo
5K22Aac008UmHEPcDb/JC9AYOTSxt2fCiuRgVkUcDEyGtS3BdL2efqgrEEUWhOR/HwAi8kVofVZC
vXb1rAa9+8amgu7qihMBThkD6BllIrOUcZXutg+bgPAmKyNb86DQuUsoPU25U2+OulC4qTl/0dwq
X/N0QJGMBJ4Er8SlfZLx9Z+/O37t6MQhcuMshOytBl+/WKESKQ0B5ubFbiaMZLekMzPrgx5MibLC
WP1sVpInNa0HQNdTSNQqQoIfGa3Qm+erCx/Z+d1YgdHGcfwjqDXz57vTGmt9SeO2HGiszYQJmeiw
30KyXFyiYKYz7x6kjCpUZrbkP4qhfK6YBPfikwzYeCeibTDP7wiyjGD//4qfaSSwpSMAqyce9eJz
uGZfjGUvS3jtuU18qmIgjp16240tyP4tBcd2sx8VXmZGCHKdH/dn6bjUyB0FKSHzYw3EwohDN+Ap
ik6Y3WVFltp12DC6r4vtVK6t4He14sC1QXmqfFNt9m215kEdy2Y6KzLtdKgfr62Yo3DJgDEHm6QF
0ew/nuv6/n+XeKyjddWvhp86GHRn+gTVrg6CFRhf/IEnW6PCtVPI0jQNWGMMcrSxghV256ekOrj3
SUzwxW4Ty7oct6OVXjt962Oe10mpMpm1RYFUh6VH0NdISo2IUSImaKQVjhnrON8AH7C6ywcb7YuN
ecBX6luLexbyfBiyq0DfqCsNY9U7mEggO+ZzZbmRMvqDd9OQqgc19GO8PhfPMiqDmDhaOqEGgURF
h16h/AUAwV9bCDXFk4tzLbSSsOrVjsjI6LEepx//obwt0aiq4HTwcQb6WewwoP8STXkJkckgz1pX
384Ks4DufO12XF64pv8ue9HShG8rPpo2CUkX9PR3VsoVpciJ5xsdKdR2zdCqhO7EOKTq1GNypKY5
7GR+5D0KmjEZSK7rDRemsesvG+i3IpU6LIkhYL1MjDlb6N5mbK2rymMWMzcldUBJ3csey7R0P9lG
+onp85ucbaBhvrAbbYaoszt27imcu/eA+1EE9b7jlgswdP3GgZr/0s7BySpDVvbsGu0bUmhIcDp5
6LuqdafNdjtEHqs57fzMjWoHJ4NWpTGJedfu+rCsxy9ch0xSMoX/jjz4eK0RtmVa3ZyBi/USKcmb
hpSQSB1xfXfJTiTsZFTDoU6Izm0VIZWdiEFmv8dd0Us/QZrVxYs3we5Zz5gBtRBlsXSmpT8FJCjr
enzM6dEkJvVjJdpbdONzh051kvIQCZP+lUCV5Al9umw8apSpL7opMXrez6wZqU8KmhnDWz1eB2Zc
nIKeY/+IhVAynSaTqbkEPtwi88Wi3ZtNUy/Dkb6ModKDpLNsDKJtuVWMfD1M3Mk1XrsDcyYn2sb7
bBxhgA+vpZ1GfFcbJa49YuGbwV51sf650GMD90LgFZ/dAflRPyBAn5IJjSKxYyG1Gj3PRqSLKhPx
hntkc/XJX2i3VLbBXsU4327vPFej/TlU/WqO5q8k7jSouFudlETPc0yliVh0rE6Q/BgZYyzn11/a
8oWcbtqzAls0kXNCBsI84epXMrbpTmSu0hb6IMvrn5wvvgtLEIMAldBCbxD8gbLvj/RPuA/0EM0n
9TliYbDncTFbdTOFA4KsHmKx4P+EBPEjDxTOeS5JsMSR5xnItUF4okeuZS2TrHrqBd4RmQy2nnpD
T9Ex2ahQPiKWb/NqCFywEVvSS4mXkEQ7pW3JwESfWniFwreNnfZ8zqT2igrfSDfif/xB0SfOEY8t
MSJJsrcfKBLyOll+0u/mVLwO2lWI+1pUTh8EXSOBE+c62yPDZ1LgNqa8e3I8NNBX7Jusm887Muhj
k1lJ67dR84eultaaSD1FY5yjffDE5V0zY8gn0PGJuSeQk4jw+jHy+LlyfeGIondVFjUByW3t2xBs
CPaiKR2V//T985ryOIOlU/uGpfZ0ADpLiu3ly4KF03XKNcSWBQmcWACa9w39iPV00XvjGeMwxq0g
1jGMHeOAhovshJy+LTt3zGpjHbSa7sLFb07GXCcgPooIs+y71kyoULRzGp/yhN6TEYJ0MryZVlv4
q3RwwK0iFCS4KS2W2jo8CA4H6msIdLNfM9kj1zWvx6qNvv30EW1ya2qcasn15le+UmQmJknu7YJj
hV4QstCpj/YRgPswUcpZ+6QHJHWbvwm15XZQsCJosjpw1ay/DZlvGJ20jHkPBPs9ZHgiRJX0ifMh
G3DBu1F8kqWYC9YBt2pYh9qSO6sj5uSqDAHMWyvuE17vHdabXGaJ9LFnHVYv8OWRxZ22Uu6ocD4w
KiO4ygaNEUs+ZCYxzVKa9TQA1dnl6wwW3yCN6o60d1ubtfkLQ/BMaMMV59qU/0eyr4evxotOFYMN
b7Ma2ncWuHOM7/c4gTNk4kOxjByQ7gbWxwrXFKbs0QV+/H4drF+BhOU2+J0k3rUWNWuyrREJjwuC
6XAih1TX0daTaCp2aPIelVQhjaaDcsgWDyzAKFL0CqZ440QPxOVjQDHszizB7L8Y+2VrVN6yRrgK
fEYF3XcnnJU/xpHX1ccfoXdeixvgjL/KHVwcyMqbaFiu1+Y39kJ5UiQPydyVwVC5d1OYZU+zoHKf
o+XpVK+H4GcG5nZ7Iqlr9j9Qg2Ds00YnHdhhPl6c74IoM7ebKzyP+9LZRQZ2vpPgvh0q4H1v2XXq
7rSGIdsurv04Kg7g7xKxNnNY54Loxac1WLPn8oruc5onwnaqYN72Uh/7GQew/bEUFHoC1ofVm9TY
U83Kn9rZBS19NIKrK1gl+VmZreENkyaB03l2vfLAVDZmAlrtpc/OYATpSDuvkSPoz6ikOr26q1+M
ahKdAd39ynHecBw8MEPqOkX2KuZJ+4cSnk/MIz0Af1IKw/iJo/4iBr2LwiGk7T/FyOrMjAX3c422
HbvKrzRj2pAGfOz58sVyqhSIH1K0e4mLPrAmCnd3rmvZ/kwtDOUzb16f0TFJh4UpCduMksXC1v33
j5t1J4yhKe8tFWjmB7ShvDV87qtOJfYX7qNeCxX9c814R1SJTaPuPLpURc/6cpHZqbmiwha6hhdL
c19f0hBiXuzQ66tCGbtF4bJV5gcaKXZMf1RX3DE3b8JuUBFcF5T2vycrg+I+f5H/LrSTbNx2R/Zj
J2a7aqszxoa4gmxk1IzuSw9eVf9hv6mRTDB/YrYvuLXZrqj02MJooBKvs/reVAtFXQxrEDzTCBHM
JQ0DbupcGK9LoxRBhNYegKsJPU3uSM+4cTJeVaFBM9qGvCtszUNslsNROi9nseNQjhB6rbeIQMbN
JeeZXIhp0oEC1eV9u+dq/OJUxXFRpUc9LbjRH5+dxOxMV6O3eoQZX4Jl7dxsK46Onhr3HqpPiVcs
nExv9DWEDOAUv6+dTgzCMkfPl17+6wjL9lq4CiUiiyTkaAKqi8W574ke3zlCg95UwBrWueO+bD6G
SM40k13Sehx1gVDToe9WGWqLHFfeDUG0YSPac9omBgSvky6yNDukd9sV/2ftM2cWXtuM82hxe8aI
40sJLg0Wax0lLC+1uTYhtYvFM3SrOTzJLc7QpU18g643WWCjrHgDOMvwaWW7WB3K5orwuVJZ4IbW
VliX7I2EZu5I04oWrPCeu7QAbvN4ROFcgm7y52WNN2grtMpfJ718IX4cEx3L+Ebi2ViuUxMAR6G6
er/GVi36asDpyi2IXfXz6bsfl+1wrqcL6qs3dmN9XqlgybQNtnjOdkvSAep7dZww7z8E56UniCRU
eBI7RRVqQxYTcpany9KfWhzIT5vahCDz2wxwkKCx9y8b3CWONP6kRkupH8fUzAJ6tRy9OQK7wYdg
9u7okkcqfXQaioB6KvxvjF3MLPYrhs+sPvSHMpTmA3FzugSzi5opod4LjsFde/f25jsbMnrsyPEl
7vVOqbk23bNVA2qDojdxdJlOxBqeXVZP2eZaeeFpH4aIBmaijLSLnd1x3nBxQzQbiWNHLFIvceIq
ZT0zvEAsi22a0hjIMSAH23OsoXUSbZib+8tDiIqVTa4SgEf7qPdxOWlO3mF8LlPdUWiMzBy43sC6
s1MNu63Hr5asQENvMcBYbs6KGgEhxGyxjZ8n98IJZVcND2rgAKsQsihP3hjm+wvrXII+WS0Gi6S9
J7YDqkQneVnU8I4z+7Hr7E/x3LS67TU9DyGbZLFcta4tXqpCIT/O5fjyHCAkPFKm8MJMILAtEWNd
k4UDm7iWEF22SkD81KA3moYlS8h3eKAM90dxbEJOTEggbd95qp55f9+azQQajgO2kpcQeHQU99g5
Tcj/FfXi1CLHV740csmLjguXMMC+USdyJWPXMykQBWF+6k+GmTtMWR9nop8Gg3ge+dlJcYDmYPIT
XIlMN2LJO9+wNA6dlN0y6WzajbH60lSj0GdXQMjACSq0LmqAKArG4y83DqnNbRe+5PHudiRDqCH0
UJQuuQ/bbab5h9fI0vX/TN4A0Yp3D02rLTqOsCMyBziJ9y6mbMROPyQHhOoVqRbUO4JukJGI/pvg
q1JErizdSNeH9Pa+7d+86etiEGlgzoApWPZiTfOegHZo9DsHpdq5tw6OJynGewcL6YvvfYYRz+/W
RQ44o1j3xTwJNzqyqQ6l0R4qJ4PHs/RDRPYaty+9RXdGCVQJ3ehtyilSt6KwdHyGkrGynkEx6Nfn
WQdYe2IIcevjJ3B9Vc0durkY48Da4DJO2LrI2egH7094fG4/6LtRazbHzTueMZ0GapOF/wR3OeZD
aMfZBghTpsFM91Gqw1a3qS8w/40exU4rveNUBg/aKMp+RpLRny/QppGPZtU6XW9e1TxUu17StGxf
dSLhW4xjKqacuflfeKyRb/T2X25sltwaz2xn3dRQcnMApDdlkrUdhPglHub8tw6ud4lQx6RpFCcO
D7ULBXrV7jxosp0LX+fXg+RQdEMtcwI0NPV6PjV2H+YkxaVFNYYeHgpPATpf1nH3yUkxDNi2PrIA
yAaaUpJrnKuXJLm/HtuzoYHYaOIAfhJ2GmDBwfJMdCO3ji/NDVsteB+1NCKPQhlDjDBVHL91WlMw
jhv66Y7BI6KeGUlavlbxC52KhlbJHibGDn4pigi1shBB12RqFcJKVtfoH8zmFjn0iHgYX7+xaxVq
C7vRhaiGhJQS4oasb+nLHF1qEmZRYCVFwp6XNETao4Tk64MnDZ4Qxn//csMUyQADnQ4hhreGhhnL
fGSGZ9VCBH7q1zQjIuUhGI3vlSEy+Tpt0I9VvD13TwK2S6naOEtk3S00NjbNqQ9y7gFxw/WntHka
25M577OmOEg1dkTklmjJ9Zpm7kzJekBk8XcoIaHdL1CEzkLXus8PVPc06Dbha8qTHcEwsRmFw1QM
xF20Z1NO5zJ9Mkk343cPiXETSahgfroceTTyphYKj02/UBel4LXdzg7VjQe5SJ3ezygsDoLq4izO
44aLfVuD8kW/szXdYQwzEJhHW0yTwAmtLJc8SAkBOAXnTyTVy2ttXZuKaPfGX+2W6GcsXKJ1tDuT
NPc9qNUEV5flGSocnxs1cqVdyo8wd/uOp+8bmoyMt1HgNRchSod7yIWBlyYdgUvOwvnzKWxxNZXH
mE37G+g07EaUe+ASHUEh3tgWIULEauvwQi6PRY1g0hNLDKtKp8hLY+ICT9AKJ+Rr/GjChBhseihc
+oYqm+VfO9TfJqrBV7Kr/etP4hwoL5FOlVShzYDcqFyCXB3axvuAGGPG55MKqyCoZor1bwPuv4wM
phQ/W18/Uyn7qSonRZLBhJD2dCnONuxwObEQ7eX39yrVB7neKIbVsJfJ3hjuAeTvPUpFwz+Xvv7m
Hg6IPySiNl1cH96hywhptPyEPcpRqMZ0soOeT4hzMMPdhACcN1VR3cub77AHQShsDaulI7HF7mmf
uqrXC4H6kQPD6sYhfHCeRJUX1f8W3L7b+Kj8k0x8ljnQWjNwJhR3uIXro1S6RyovhQmcil3B4I6t
0R+pqRMSfEIeqFQ/9YmFcJXgiP9YT8rS8Xs+wR1hIkDflDp4FaOwK9Ibp0VoYXexA8sPkoUpdtem
o316f8AOGnFiZbRJaX+Y4mYpSM6KweySqtb4+3vLab7a2UTEJOsmKiFdLqqTlGwNLaD3OBvtmsZD
tE4/d/zkHDzlCEh2NLNIOzMAXrAx3SVF7zwxxuhZLhX4wlBP54KFsLcBH7SQWiiTGG4w5+RRZixk
SNYJfs2iPNItp2OMAFnryWyimAc2Hi54MQ5FQEx/HGWvVZN2nXDtS74GnAT98sb60Q3+dFN7rFN6
7yUxAJj0BgzpSWa8wQiSZASn8oAZRE3I8CbLk2QTZNdAoTs05xvAW8QRBEEHZ7pWqUa2YDLdUzhW
dHQFWYiOwERwV6I3Yfg7WeaexpfBGCVWLSOT+4ibYbsPCjVAs26jrLeakC+vOlNY2espTWrrJWSe
tGcfl4TDejAWTsGlXTWCgHXk7v0fkebPdL64jjhKIA377RCOHrLsUX8vvn3Rqs3lLKwuTydVZ80q
USsU7XvzpimwKn7LO7Wpp2SwG/DztvCStp7WFyJhcQg+zjlo/puI8qJJR6fiYOpNRgjx0AURxCmp
/e6VjO9wUCtTFj/sCLainP7F/T37L7hc6GHXiiXIBNeKvQMspC6nnchlLEMy6+E9KQ9cfZTBNTrH
vTuUy2vWXLOwoXDL8WUmt/dsYaeySGuVtAOxp4npEYq41vzPjLunUX/h0pqEUCAVZAnt0P/bJFg0
sEzYS5O7vkzRtsIAs+dnNL7FpcNwuoHD/Qftpvm+dSm03xbQdiZzyfHhsC/o0fSjfZpMFnple8WS
om3hDK4W0VbjjtYr6ySKmXvGeD+pxZQlOURPskSnE+M8s3FfmMxLxfTD58D2yhQQ3eiz002+wXPS
ngKWPeVWybPdmy4fko/lYIkq8rV8Egu7l6n7C1lzPrAcZfy9XMrNgIA9eXcbTbL+dwPrivu2KoSw
9cRMdBWJ1qfe0OcwXh7tEyj8bgCtGXFvujebhjYeLpUmuCkWBKzC4GQQ3NaNvOJYOBWj0/8zvrpF
+GflQHs+TRi/+tM+p5fo6tYa7WhaW4f4hdPBiAH8epen7eKO86ATkmTs/8MTSl/m4xlsdfIeZUc4
vKZVpxgy/jhUGwVIpTuS2hihXxslFMk3Rk586sWf2nMPHOh429ojAr+Pf8w5Xh6cvM4h6L51pFZ5
y7v4lVSr9ybQ9DIfzuEfe7d5SjinDBQwXITdSsYC/pBe9u50TBnkxNvSMuS6LRYNlIai3x+2627P
hDeJhYUf45QB1BUNmGFcAY9mUJVsbTBnlaPlVKl09dveAz3ar41WvA1Qu/5+EV5T71dNquGzUlaS
dDLk5OZElBEtB6BxK1Dg52wYve2RlRdhhZjWOkZPQ01Z7vYQtbmuyMrgJ9Ihujv9iPm8tyt4OmOJ
PacVJTD8ybedkPutvgeKCfca6JniEqYNF6K9imLbf6U6OLa1bzUI7HYwD9PZCDOG0Fr/JFtM0hpD
xl9JkaspxrhiYQ2jXUZuwgGl8pCUwD4v0MLPASszomZXgNsa6fFDgsObjjvNLZo0ikA1iwWZvNho
910bwjLnfZx2qDtaSWrlyVOfG2E9VczVSFCHzRWJpQdlQjmlGfTcO3HC7c3URwz8zuP3tTuJhQMW
qSP/WZ1qGEDYXTcFQc1lLNA9JWzBz5guBgR9/9dQS2u1H8CBhGa+4GL0KUgdhsn1kWsK22TejtHT
PZqwrxI1K29uHu0eBb0ClhVqveDVKH9VdbP8qN0eLf5fO2CQKO3WHrJthFhgGI65OcTSPW5OV4Ve
LoBqXXyy8yOa54r2OlnAjcaOebemMTKLaNSeFrqEsNCNis5m0bqvdcK53lYmQVZEBi6t0r//iibC
HGIy+hhxMqH5lBn+mi4bQgrrxTkdvhowndqZ52HbSTJzVFwkI4SkDlBhQM+ILBjt+RMbEvVmrByI
b9V2qA+o9gd/cYKuh/2ngdl8w/KKG7Fm8J0lCDZ1tY/kSYuCXcI0S3UnO7KEF6OQFyk0NpbanvGJ
OiExsqJf1IiJ0Mn/nDvFyW8BPaFSepjkDMThBARkhmFkwgfNDvRQSXev0iwolCbk9YcLI/aSwGBp
ggv0zh0X1xypcoqDZ7lfqpwTv0gFtQ3bghovmfwQCHpUS/9RqlAO8fAlPjRwSIZvBGFuVeA1EqfN
KCUodVLXLYdJ5u1gKkB2nehyG/j4akao7BXpnphJBotOerFVI+OX5AIOAq5CCgPoUTDQE2dEgPev
5460rofIlwXsqqz4036vPoSynNICkwzJFEw0p0GOjmB29MtjEH8Sq2ub71I92Papy/FmEcttxtCR
tVoPomeX6FiaZcj1rIrc6PpdkyUHisYJ+3F2Irvy/EKjF8QBqHyJAF9DaqSNztqfGk251jsSLdSC
YFtenTl5PFOQuRot9NUXNfSSpCxlBlCqaj1j/S+w+N5RaDQTO0NEgJ/ygj8sCJx9i5Meplb2c2Kd
Ag/dYinTyz95JF+u6L8T/vmHXjpnbc6PDYFUY+Ml3IT3ObsONDwEEvfru/NdIs85Wuq+Ls4+3vTG
nU/HeSa51FkomK0hFS6I8ViyabLLIZHQtMbIkpxbobu0Dv7bYxyz2X6Oy71rCsV1QGdIbUPnZv9O
D7ZlHYo2ZuN0qu5/shrXVsliPo2xg6295FPnT3WerEq3pL7VfhFs6yULVKIXbfE4AfmuIu+YpSGI
oUIJC9he8sOy6485k5bGmWOBCwFv3pkuMzup0fx6zyqLDKtMUIuWdbaRkzKLsqXZz5kCxIgwC0F5
wz1NJVwh7UclW6l2YKut4X4lb5LekgBnPRi7SDMO4XqU4UMqj5Uu9rQnauRXLzu7bNoVhUfCdBl4
YlvyEVQMopEZ+Y7Ud8CgLx2YaFftEflUbVwW4zdhS2rnUdUK37NVjsnRIuP4KFZlzHuB1a5kvQdK
QYF2Jvk6yFgZHWIXWGYxp9/E3LFnEoSEfmrsvz91JpMn8bQRnR2ZkRBeY4Xj4ktZaoc6yGj2L/BW
lv0cujwLLIpq6ANMk+N/tV1dICvBNk+FJOWofk99sXw36xev5Y12Vll0OrWNFZPOBABcRIiLSLD5
qLkIWYI5+qLKk45n9drdOn5Shv01Jb0uxrvndZ4gYO1U00Fiu5KJUryQNP77gsYjdwde+5uoZdEs
j+DrwZoAb/qvSzuSmHx2DMLLPx8HyZBWLnP+0QF90x8WgW3kmo2K05cNMrZWozjG4cM4xdqd6hbF
0khNJNCS4CDji3+I0mK5MozNjLl3glTwh0DLXxygPS7KlmeMYxCoZwJwgtmwqPF+h+aiaI7sidJT
iKKqkk+10VTps+UaX5hnsj1omOqrP2lRozPJC7q6MM/eHU3MZhgNVKhnHzLaeZav6iVI2r4dXI6o
jVYnN7JSRWpKQ+5ojtdsSK+arsbrn2iQ3fapMDiRJyQOgWgmrmYSGlzxsiqxVxGEISXVf4E7vLfU
FKhue/HMkuZMjvHCzteoFjF4Es+QXG03UivanrY1PdywKfEJjlGMTh5hu6TD67uYIX1UPPj4iCDS
oyts5xBEoZNc2QAvGg4PHHCCWmxjcn4fAtEEaP7UoMB1yKhGobhXcOSs74Q2djLX+zT7+Pesbvk6
OpQtLvnCczrvfUJy8WRx4qWSvbf1kjPgsFySrzBO5U4jDRU6Gx5MrFlZwBX6Q+9N8D535A/J4l7u
kLNQnDLJ4ZE1T3NcjTPR22tovzgqxI4XQDM5s8VOTgr66r12bozCMqag4IhfPIQgHBgzusPxTOb1
ix6MadkNBDg4RUSBIanKQRSJJyB+0/wJ9naN2o/uj6TTO72LULBkZbsV9e7WsDVo51zWZlAoJRAl
ms8YBVXu/TQjVuavVGvKdQfrBHyyq/bikiaCb1m9o5wkcQcAOeZ15kU30EHzmyoaCz0Ey5kr3Xqe
Kcz8YM+cGgRmorq+6yII1oHeHufMz0Jf0atfSVdI0E1NRi6PPm/fQEHr5/qYxjkbEinAOD3HPBDz
49PPNaSHf64TGcgAmXp9JFJAGg7jsukBQwanD68Ttt1BMBWhf82Zy6+61QTZsS88zMo7P3vKjwvh
57/nPg3LmswsigNgi9c+aAAvN/dcLvx7TOyMUVkAHa9XfmqtE+16MsiQ3llespbXW4iYZuF8jXNL
G9krnsL+1hbfH/4fBIaxSRcXmVyz4OtsHHwLWJAT5qJooOoM3lOij9X748f/c8Lh1b2SQz1rVhS0
iPGLb3FLDXfIdWkht8crm25wM31dbSQSiPwWKSqPT7gbMNuAmPwa2QbUqa1UIxscSIguMn+Z8tJv
fv8fJUJ4c3ft6ZGLSNe1Xfxu+wPJBdrUcKgk4zSXKg4S6eT9ngGH1fqcn35igqs0Rf2DX20SDJe9
OFcQELiJ4ZQkLGmMSNpg9zE6I3U2o9g5jDIfajh7o9CO6S++JqUKy/kSxilQp3lFLnGblGI8lRq3
im9SBcT4WWqatjksl2+JqHD33oxgzOFp0M7bEbm+3mKugVbFu5/1RrUSOOFOJeMGBUzcLWiC0zB3
iC+79M6XbjgA6CkaOQDl7ByFVwO4xvZJFSjmc1pKBE5NmFuIWQSri+RRN1mYPl85OFrVO8XHQuOs
2TJAvq8Ark869Oq0kZxp3PQva9sK9GAWPWHm9rZ5GUVXaAu1AXFtgV5WCIRgLw48Jd46XtjJLyPY
rU8o6XJZaHTWid6Y8eq4MnAEDT/AexhinRXWSMDgbADpJfoKdvcGLI2OXuj0IYX0ZxH+vvmmb/b7
LUNOzvOFOi212ZZX2Gz50BdfSxqhIiC81+G31TbmtTKrym/30el6mjDPK/TCcX+1/xf6DoFhQQgn
hIkpX2HB+vAbIOO2IV8LjJ3Rog/3EnGgcgKmR43CZzitBKJ1dO+7qqj3pg42GisazQu4gaYPs9j7
WQ7smHvvwsRVBhEWai76OYlZSVEPZwUKCfTGZnSMndUdpgXigcNZkFV7EdEO5hwkMaqF4xi1G+eg
+h94JFvV/zJ0xdtAhojpux71rQc1R4RdPBn06FPV1jP43vStWFX6uUsojEau6uV2QrgKMUwUfRAW
66t/Bilh8nYXq4MHG1xcJvWk9gndKl+WXsrDC0dvEOsmKkKU+790lwWZfGIdjA7INEJgVOpHTLr6
EUZuBHGVSrEgX5khLoQ7q38B/J53g/fMSsLItIqMGv0E8EUHy2XC0K0R/jN8rEwmjJvKjZHglNHx
4g1TvnworQ6FiwSDBYPkG2GSh+SabTek3MWBWXp0ppff3nPKeyWWOVsOB2Z67ov+jlqsSU8805QY
CRZZ6EMZERDhV50weVLmzLsClqC9sNWLie+v62quqGP2Jp3vfUGqGTmXThPV/y6A5Sbk+0gimGw0
0ys5MINKfhm+KOfd2tFHNTBpfkeComjz01s9Vg9xxJUtVxD96MX7S9Pk266pfIrc11Q5jE8MtASD
9Z2XYQvBIQumtix50Vj9kh76yAwG4EM0YvKyQpKs/dvswCz9bRXWP8ltMfynhhG/z+rdtNE/KwjG
ADDbSfcWk2NPTMHv1T/GYNEma815R/MV3DDIuPz6r+g9u5wbdr42bufTD7nLXOXVVeqTqQuqK42n
jHuk8mqjfBpxWTfQQauOj6gXQRzXgcarlmupCc5mk67pGm7RyRpvajW5uwAd6XBT6Ol3Zstf6OSw
2l2qgkmUvFSlXLIL7Sn8etMFgnkYtznMO0gLILKW6aL5MsDk4eaggZFOmFpbI7FneZgJBNbQlhN1
/jrSv8z+qaI1pL+NQrtXC30M6KaQOyQofu+Jmhq9ByV5H2dTlb++Jyq6mkJVug8i6HC/YKq+7KNi
zvWGf/Cx8osP3Fw3NyRY99IsSfdl1NTIaN75SyN+uEW9O/FR3n0FtUKJQNAISpoF7P6nU3DvLvqT
9WGrYgi3WNDPX80aL4WwX8wz5peQwV5PbYveWnGVvXBj3+Q9QlEky3URg+OMOmNG4A0KK9p1Ihup
Xw0sUlP2eYt8I/Arrxx511v2UoV6KFpdhjeAd9irlCBkrZtZZslY0eTdMSUllikG9XssANv7T8jW
GaQ+c1ilA+UkR3/py0kNk6oZb9TPiYp6oEh/Slg+2JfpRARBnE0gdV97LtawuYJ8qDHwpnW8F1Op
3o+hBVLXqWhlsPCtYaezNe/h5azfsDofVz5fRCLtDfGfrhpOaryCsXa2t+EVIIAsj3Eq2DSrFLN/
IKjTihFG5urJ9t91GgrzHIEvnS8Y6s6bIzxWZxz98SGGB9VLzP2MNKIoZJwgBycG84fC05BqAysk
caF6W+de2uJayJmKvhT5Rkja3EwO9zbpc8MulWCKhatnzRXAyAPfBlMfcNAV7QiyXBQ0Gv63RWFd
A7QcS+dYPjHCIq9vyEh3SK7puIdiY1xA7EdIgKBcxffPXXbTFeoKIKiU4U4M2vQgu+ttrd6f7D/Y
wQcD8NlaPXfI2oC4/24fQVB7buVXxDdCXdjrZcyIVKse2PvBSrK52zCHN7zYuQu3yi7w+fHnfc9J
LfgyuOJYChUU3/g2WydZrPpMosLyBRgKZFf86AHLPt/z4wPQ2YUF8bVh8V7xnoUwVMqWJIVwvp8c
xc+PtVBrnFRWlSF/uEUwpDVd6EDadPloulCKAmbE0p/sNKNVA4zbWetAQV2MJsccAQBAtrDxYhdS
ihQqn+1UmnkX4PxGP0mn7vGWBUQ4vHLJilT8qPu31g+Hv+LyyxHiz5TZZC+ehmSghRPCiFeDW7S3
olixFkw8MN2NSbLbZ+3QoxbdvdrGB8v8QFTfnaf5aWqU1QAJTwCSN5uyKGimePXhENN/7WlDtCkO
w++XZhoeXpJ/9YoM0TLcJIB7kILAR16ljvrP3S6pKzBWAhuDitLppHvjMnmJCKufOgQoKfvxJHHW
41ybqIHmrDm2PkWWxF/wmg/hDCSPJg1vYd06EXWWBVsxrTdwMyUHs03NQK5a4a3BT/Y4501Ykphg
U9ehLMeOBSywtGDMmpWQvNsBgCu/0ZxtOmO981d+Z4kg1OlqBn4wXYtnHv1dq42TAv+6yE0gJ1W9
axiNsokpLBJ4W4FF28OUscP9iJv2US0v9LSGHucrED6bvW9OL0njwD1QXHLMjJI+befIJi+rpUxC
/Tqm7eCH3mo6j6nWUD/xmJI04Fn0RoGWtJjUcv2LQXQwGtNmXGDYl0LD9J/ugF9+owqoUGTgth9a
8J8hstpveLBV/sUHY+mrs9VFgaqcaTYlT8P5o/0rgL4vYxh5A4XyO6/A7PWfA2Xz7C7I5E1Lhkn/
XnB0ACr0TJ9m6f0s+26S1qqfRw0flf7tBh9W6RMio5YyRmhpOi3ZNQPT/RrmecJ8WEzrhigVO+Nb
uaAUWDdqMJZsykxsfDtBXZxqkTKfOTxBMwe5vNitv1JcA77RjydAggf6x2Tzt+MLf5vOXwUKjFfW
wFggUBebTPxiKrmiA0/tqsokcg6uQ6d9xT/y2ITyWn6wOcIQF18dxAvpANa3dtWlEYHljccckYGi
1sTxR7oVxP3k5GkUnPGm5HdTvdOW8KzbagLarz4181fSXl+xtYabWkze40i8rOSqmZaj/NUGXYXs
S7y0qY1fEzRnAYXzQ7smF+LukL58R6PpeneBaRso2gutBVJjBDdtbuesNBRZWiwuSeNc8aWNQy80
ofO7oM2+VpTjM8B8cljeW8qyhxLNL8STZ695D6H9hCWpf6FR0/uUpW8tvA35sqEgneDB3XIwHkfK
CsRlSZzSOG0vWyy97jkJ3Go4rgZk+c1CaYMSeip9KCYV2fb+WMRn+EFTTdmwRukaknvDctdOTNHE
SdhY0p0obrD2nVPaSZW3mSLbetJygoImfjbY9WwqvgAuEH8cKDTVrUHrXnvjNmvsMSQfeB98jPBP
nny7Yz2cH6CPLJqovfGTPnEYwXbRWmGiG4qwwbtB4IkfNe/qoYSVmCYuHN/ZH8Os92kGsHJ8UiAS
5Wb5dnJMwRP+vCvYizhu02o1wqLM5MqYCLvBFF3EFLYKDHKZSW/20uzV78KdMdmucOYor2cVXxWA
WxhKih1VFPHCHWWGW30bjQLVWtG60ve0ouKkztmWdABsxoPU8bnCkvfSCFMpbWuLKCrc99XXhv+z
VJZjOQpOOTbQ6GGW+l9AJtjnCFuYPYsG+GPnAT28HgmqoXXXbe9IXLRpAajDUUA/ur2y1ibja3/4
BqwmTeoSUQGco3H2IJ3hc4AINwwQaiS9cMQJfhQEJsRV22B7pFNAz9oPletJbN3+Aoj+52gPh4Ld
TcLQHqW3wRr7HGZZLrrdEige8brPquO4GMoAuUpZLff2AxYRBDVJ1PkRRP4cU6eC9r4N9BLqoswg
cL+0xCnCQalc1GwXkPfbfmvx4dNuoaO24y2/E7rdB/3CAal6CI/Z86IFlQYkIz2COX0t0zQ1O9yP
SR6Jeh1m4RO5YHOvx64WulEpPpurhFcU543iLpzMYs2L/xSHZDSWwHqzPScNLq/e0zi/I/KxVlzI
0rQRWJnxF857x1aO4m8jo02TFA0Whn0IWptr937qGD+RhBMpmZKN26SkMIHssnHW5wdUoQdNYqdI
b8Mm0twdJjjh07fDxYeASNGaUHOS0iMoswHdlzmsP7sg0Y5m7PjyyDH2CSTYtjysu94BAVelmYuN
YSvhg0zUU1IxKKUaTkrTOxeJJHa1e+pld26Mq4Aeuf3TMELn4xfe4NgN2BaIbNMs8vny75jWw7Zy
Xfbbx1sPVbECZo7icqFtZ3+L
`pragma protect end_protected
