// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:35:44 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
FqDPGFfZtqdWYC/Bc932d8w7QVzpSj4NoYrqZWL15BHP+CrRgHxOarivlLgu1jT4
ShLcVwB0s7J2yjjEDLdFkk+OvLMBlzs2cJo7Rxp6BEGujNshD2qv2HsYCFxegCP2
43RipwjuUKivXnJpxsmZ1quOqUyO+3zBx880nsyPCTc=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 4160)
Hm6GTQ60gWmHN0ylAdyTHBWsie9KCIMDF6aTqhgfH7VW+kjojWZFff2dutoSaQ8n
5MxmpSVKJdmdVOwFRD5g0pSkGJR7jWsltzkeIeDzppaLLASWFHbzcPVcth6asRyI
Ln23/nFyDtaPrrlPM0Xm7jDb9AxCcTZBMCAe89ta8Scm4set5FmkzvUoTjf1XRhj
ESNJGDbR96cQe5NNtqgyo/wGlvEKUSA73s15DvH1hbTAQ43a6fJadjJrlMUnO2yd
4Dz7BHPVwL05DdKsOav/uJZ3Mno7aDKfcNsyXerr515O5LFR9n/fPt+rXMMdZd4A
y+z/iNXkuG32ldpSPbltsGSSrY/phYixaypIRsdwIMzXQqO+K9/MTgvTlxRTnwWy
YOYoxzgwr/EhcrF87C48ksWySB/77e6rp1+V6SVuZvEmxNYz4qKIQcIYBNgel1fP
GNkXeBin9CaWJykLuAtyC5OYvQAIXq/rbSvO/+mxakSnjjKJn2R/gkSLOwL4cZI1
NQJckOAybG2KjiZoCkoYFjdnLlkaHmWdo2CnIz1AqOk/sYFsyQq9P8vYaGI3p7fY
wsCr4VIQ+QfDOik17J2oENfoxf8DSv1mALHV+qM2OzfHh9tJetUoqjNteqvHYvmv
qev9kMMl92Tv/vmYXLRfk+wuQDQoQkCaOtgZq94ZyXYe0vWct8XAVJ7V/jbVGcF6
YHV006R+OfCOc5nwHvGC6p5mD2hCWbVuX52P+fZJ2Jj61Rx12rhWZEJLb73tqZrT
CzcKWmAA8mFP80dcyIKlfY8JK83shG/ZcgCz52Q6lIsC2xGKASnaHFuyNI51Ebzx
pFB/8gJ6iT8BkIUrMQuTbYJ1GNZmLR2VhHm61S3SjMHxUh+IucGnb4CsGqIxnfvS
/VHH4invA8f75qKDfeAZ4bfDlOXnsExEKaREj8Bvre/Snurxbbqmefxyhka8B69i
GD8H+ozoIfSvxa59/g4Vu6Ti62d+Qc4uNLT7WtbQ0IdnqYpo8Cn2m6ndYf+6CvD2
hrKkiDlnmwupZ5uPlrcwYFuVREsVvKZoZ77B+PgskChyIktCLjXt2nt3/h2IGh1D
c1m8nmeHW6ufqHTuZ30uewKCIo9hiExZQXeJvDeJkHJDE+43pONoLYqGe5SW8wlZ
H6ENuBOU4Q4X5Ean7q1T1ro5mhwjO2grzmdxTm3FKJlwPcc9meNDamdgsc9YRXnV
lLgEWqugXkMG/CJCJLD/SKRT6FbRzmptPhEpVlQL31Ljn5DPpp+PiONvjzFvBCoP
4sKL9aGad6tqNNtBWv+DsJsWRnYXi8Flnm8BDAn42sRCmVvFrJ20ABBVRJrj03lO
jerBe+TVuJMzuIZFZSujuB2M7mLAsb5MhBFDXS8qJV4sHH3EePc/w5/r5aq4F0VE
Bw4F120zvvUrwbqME186+8mwQ1tqf1jAXd/s9pylHOepvARwnBrxxLj6kU3sgfVk
7xRoUgr0wiBWldsYBsxSSDlKo7KXp66WD6gjUwPmUplsf/U+tIutvKm+zZwwT3BD
2kF5ArEhu1UzLC4ezCvxmq+o5EaI6NfB6PCXe3El32dh8ERMTWuljEnWvNbOEX3E
LSVCv9HSuae8gm7EAFbIGW6FBvnbR92q+iv/RW09tDQscPFtXCQTFCerty6i42NI
DP0pnxqcGlQSo+l89t53rTvrebQU05xDW23e8ysMl/Jdtd1gtrK8qUMg6/7OEFWv
SjRmk6HRRNu7IUYcGwIdNh1EsKrbVdyYm+m9Q0vsLK7ZKLCDBbBP1dXtSBzlY9Zt
a3NBmQcpXE6b9LAoJ9FjByVyMjyQ/fYeFsHWAaw1lzNQbgzK7hYHMMIc28mWJT/8
H3QD+fTE8WrLY7nXNFGJJAbvXKd6g2pyQL7yviN1hTiaxm4wZzIPhy0kjEfmYCl/
hXH479uSMwrELVxVBnDOZCRfx+IJ8IxhiikjqeTPwzXn2NZVgtzI9Gn40FC5omJy
vEOegs9gixjq+EJooWleug2fjDBJqCqfw57oj6Hix8Bc+FRJQbd57lX5bBtK8/D9
szPVzJ1y+2l7HSTId66svFEXsnlZnqqfFAB9sYOgw0ak05R2WC0+GTVdqkSpA38j
t0HH4TeFfQZUy49nDrdD5OnZkXqCBZaO1oTHgbBWS/eKvy5ymVaZOL6xyzaaBoqO
2BLfbdeltrfWy32yd1Mf1QWlcqZ8LNNlckBd5L+ExKxCVpBTkgn9uIzYQiG/PKPG
tjYiLPXLV+MFBycm2Q5DaON2HGWAnzlHhAoO9q/coN0u4WhyyTVGygZytpmKYERb
w+dFvyj9+JRpW1pcMceSSsv9DzBHCECv+LUQ1s+GPGPeDXI+pHfZSAQYoLriwOcW
8Lw8ulBHbH4SEufHKy3S6z9bne9rWKLs2ZKkmxs3q8C59GCodOzVvFpooVUXJugi
72EqAWGau2SVr7KYdFD+X9D+E5JR0NWT5XBHWD/t9YiMQYhwbzAqQyZ2OTeYQrcT
yqGA9EkydYcABWnYk0RuzcYjeTz1tXAyvSdAbdOgkGqSXGwkubzd+f4JW5+sjElC
wHK4T7dud2x2zMKlvt0lrPJm4kBdAyCIPQlkcE4yRcAHe5E1TD6S69NZHp2WZ4B9
ff/++WtRvUvEUBt+YfM8VdnvrzV6wDJrRSc3NHBaWE507iMR3XPTb4QkkiygrfRV
TuRcKqq26UNFOkVjjnMlqLLmoF/Na997vtkVU4K4BjoL4ALxbNzi+aA6z7uZ0ArX
BQPjCyPXv3rvOezcQJtEcQ/m5y9wiFKi2js1CSaEnHQLcRgr0Ej/GiDaKMnGzrKg
DujT6U1DWndqkV1mVx4D53Nc7tygMxfBAufOCOMIh1CfCHcDcO8yc23E1zP0iirt
Gq1EPC0+2Mbv0pEJrlq4nOBBHSCcxZUPu07s6ZmFJHrrXnL6VU28SCgBp+o3ceQ0
9tkJfdlsFNQ4kMQLjdjllP+Iu6qI4u5usvtPM5qA2bwjZTgeOHKsXdUgEnPcugqw
qlz2kDsDW+CNu3Eg675GCQ286q+YJWReRW6LjTj0FwXhh6F4yLFL4j+F2dT1+fk9
RodRsy2rybnNZ8SyOmqdlwzbqdc95z4r/YFw4QFWuEDKO0qfLiFCftXA0U4vT69y
/8PIkAwzDvB9H8yD+COpkLGXqYPI6Ocm3SuI66yycVKvXUU6mhgOYzeAM66xE54U
Tf7Yn5Q7hCSmI56rjH2h4X1MiY2cpvDlNM/bh/44/LfUelGbfrFVdD8RMKbSIrTX
yi3KkMmSjNEEH7kwYigARETqGPvNi3Qi7ZIy7wr4wY9DGQvujXz2Pp3vXs6niIhF
A/JIjUFa9p+dbZM3cfQ6Wi3a27OwfV2jTofoHdhhFDk9B0fQrGO4kIC6G2k/TdK+
AukeHEIidEA5UXaq8yMWpjK6lSDY+rwxBpfVRyy3ALvvGlUu3Z90JPk05XeRdNiQ
QZHgmnGXWxlwYZxaLWkB8pKQ9m3CHXy+unuvMKyZUdCXfUIlZbb0Ehz46YD/pBEU
zieqPphRdkWKOJiF6do6M9dRJwsqc8ZG8Zrk32BMIjm+kJLfV93i300DT5upf40D
rFyo7oDxILXFN1XtnM09Df6Nn7m5DP0a1ea6tgcm1Xj9oZ+r7TtepJ13TVLZgvbW
GzlXtgUlKgtp1cY+LTFm3NJr20Lx/ube1eQtONEFwmhzy30uHN6TZh9qafeM6UCh
1MCRtd9HwyyZe1YYihqm2EBn1WMzAtU77l/fFDddSSj5cShAYrCOUI9Ar8xVQStB
PQkAQw172KJKj4aRFy4ennqGBoeTl4Czsha89WOb00FZm9KlBg2J2aocdw4Y2RzS
Q0VOgvsiBQL/gRFk6d+pZ+Qf1gRx9wzwMluhFxV50+wGTYHUK0JXZesx1T3Hn4HT
kXPFF2lkQPwNdMt1mYb7nmOGtFp3PKdUu59la7ME4h+LS17gIZJMqFMfr00vlm5/
ZjRoj7bcT+YMO2vy+mw2eLljuMB+UYp2jxPUkGkGlxRNYNZvAKNBWhuWFW9Yw9fL
g97Fs6egDdeKmlDpuMHAB0LFRVtPRUXAOYIiZ4j07WcAFG6aVV0jFZ9Tjz/ZFBT3
RUnkYMHciRmhjKxYtg0pNTIjEom7TRmUhrNtTCo5eO2Q4W4NseDaYINtFqtol5f/
SgtJhmdDGI3W6Q8wdXEqfltbHPCzAImPIs9vbITKbc0SKWJXqFGnfkXwrpXhywyS
X7YCGOHiceNYoXLwrRftZdVsNQByPGD2xAfYDDhVxP6usuGpEaiSCqDP9OJpBSj8
/G++B0Wzg4ALEoi6qJgzGFDDXl6hfrYV6WlUDvl7mm5qGjO+k1rUzvoPfMTiAMoY
DvPi4woq8CuZ8i4j6nebs/xmC7tXHfjIApYVN50cRa8ssuHYJMic0TmTlWxrL/wk
tM5uKlUUnFaRDrhQVX4a1D3ihBFMvYMJiXbHtSxOcSUqOdySp6k3Hd19jAEHPm8L
cxdFEGUZtLzXrnQOCY1Ck/P+Yj63szmJeQIt43/04BZv4gQVdyL4fGGSpa/Km9oT
+BONuvJunUudki3TqjiLF16DNYepQZ9hZYHDrgpX5BNdAQ+YIi20K8o7bM8D8Bqh
mdBuGqg6bYgdYjXhnzXjeUdDxhHDe9htibEqQ1ryPgkho1hzyBfDtBINnmBdrK65
wyeOGiyWLPHS2p/QTTMd0RJ9897UX3zI/JhCUjdZOIO6DJOVWquS57iIsfXFfbC8
69hfhSM/iGLk0nxt+jXjndQB34UNgo7t/Km/QS/F+lWzUhK7iftbvBOnEP2phLU9
R7MADv9uDSHl4g3nYwmRqF1Wv/6R7i7lRxc/Al8vE98j7Y3CY1YhmKPyshe7u6Sb
V5h+P1LTjHqtiV2pFBm2FtFvlJLR5uBFimz72GqB1g9PJ0VOqdH6ysj3cRX7mSJa
daO0wYxa5283/DVk9fXxGtMIhqOrJbqMS7KxPGCnJRjAy1iGSe5jxcd1hNzNCqnG
lphd78CN7T7f4mKrA4TnGTXucm46ZYBv8u8/20/JbmDK97fb97dO1Rl+TZEqO+cx
vXf1VgBl0H0DmeucoWZ4susS1J9AdPiuWZ+vh4UpxW32hO6Uvc8Q3EeRKHXcpBVo
Zwgffb4Veru5tQPZME/92S628frfbD7bRMdPgEQt8Gr1783QPrqF+B6tct3XDJiW
vL1Wt0KuHtT8RBWYd79KhOBJHooJTPLiWdEQ5etdj8rdqxBrM1mdeV0w1RROgkfT
kMgN7xRIDaLMrHDabGebBCByH7b3R8G7ySytaPMmAhq15u6pm8fUXfiouBEhAKb5
mJGUUd6pNu+ldaW94cw7XJfL0ckDyBRjct+e9KBJyjKBiFaHfMWzUx1kl7CS7o2X
KZqf+Is2F3WRPpsq1vljyAFJ75bKIMMBUmijRx7oVaggu+yAdkmRdtzRe5z/pMW1
rif5pXP1UHwCDjfkHnXeQ+sFYJLsv6zfWKhBVxOaBBN/rii/CNo36ctDkWJr+HRw
CEWMLqjznP1A2gxl4rsKprStDfe5UuecKhUKFU6q660=
`pragma protect end_protected
