// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:36 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
ZFq4GsmQJOZMWWBTtrI5yr8V7wQOwCr5Fg1Q3pXuBMaGuDvO49753JcNJGewAdyG
c3LmxnS55qxC1bj6sfkuXd/v9tesM188Ief3rkKxRdi5tSjssxXP/XYVh/mSBSGZ
2SlWR5ORPFvwknQJguPk5T2qKz9+DwLzYkaGzkNm6lA=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 7504)
R1syXKAVtuL01hzK6PRyVlJRE7f8pBDxqYHbGaMbKTCTz4Fld4hhJNvP/hYGa0W2
z69Rxfxb22AX6yt/MQguphUKieE7Lk3K+xsz6X+gIT8RlpWMl8SbNePMsiSaGgSf
sG1JAm44ekUiWAw5n/n6KWa+8dGHgpmULes6es74biMsv1LdeBGJEsXpHddcW3qP
2citUpdvSL6237p5NMwyoFFqTYLCXIfTBqdES5+/VZE1dBfHb1lq4zLI44ksjxaH
TIl4szbx6Ky1E8Ibdbc03PqQhyRA22HRsHKu5gMyJAHdWPhUlpM4l/MKlSp6GnhF
Tlbi0vsTVOD7ycVMPt8vCII9xr/fsyVQo0L+Q9ZBML0pqRi4zOy7Yhb9TlVb9kod
wNLLmCp1PNBTrSVeoF2JyDsm10gCvQjfHBpDp7GHP9e6qj/gI30ZOI9ZjRP/OCIg
QkznXRPZQombIRgRvEdBYe0j7Ii4n90p2n2TXzfEjgXeRBU5jJpaOFwG2XOENUUi
jH3ExUgRg/TZuZioHpiWaJ4X4RwZvdbDYrTwlGIExIVqNkqiKZLT4smU4t9fH7xz
yiTNebwA/hDrIXV8qyCANVNj0aVv9rY7riS5BGAgsM3e/Ujw0DmwhIXGXzpmZC1c
T45Kf0j3GHTVbSy3o0UkQxxoY/+olDLzYQhvH0dwo6H62QJNJXc2aEm5YFCqD+Q5
5KclwkPpNVy1eoAH0liz9j0PZYOxsdsTcsDfViPRvFa+F5Xz5B+LAK5/4jHTy989
O9FZXaNEI85EqGYDAwqItwiAwfz2R+suIAWP/G5BqYfGkGls+4rj+JvXf/2uRjvO
58TOvHw1lrHx8xcEDLxk1N58LSa2HE8CbPDEzE4anJpsxfGe6pC0SkOe/A94qh5w
FyVJJv64RJcEUd1GKNBJT2zKL+d4NsZ6T0Zs/EdwYUJdFfK86vCZSDIHyRxgxmZF
vUElgmsFR8X0L59JKqcE/7y5J6utScCK8r0VkznBKY2WI9YoF+RlCANkbUuGTHzd
tLDiIotFLoZ0y9XTgdV0CfhJewyT33jsimyHOxsWRfYwwWpupQ0FJf5IM99jMzAY
85h/0QZZhHH1szY5OJ04qdBSyWgfDEHr7HqI1IxM8AUQoVaLWALoQPLJLAhZ7k1i
Rs7TqETtPQDV0ecR49+QIPnJ7niZB0yxQjSMjuUpiat06ISOpYVymFhGVVJPp+if
zb9HedYp3UtUz6fgzF6RJiD7qCnzMrpkUe2IHR8jeYGNQd179OGq3wx8RCrcF1IN
EYE8dtyBkLEBpAmq/oWz0Gc0G8nbvVNXuLv/s/kC7L1uveYU1IOlsLKbfr1ugsjZ
G30uvjpn14K3rE3+enhRu17OEH2hG3+INqupv5uAuowNGynljbGhC8zFkHjKX17y
AJTlYGQxa/s8tCafK/kVT8gu8wOLNCEBSW6L5SE/cgtB11gSYbl7VlKmmvXrGU7y
VeE8Qx3RwTqEv5zKhmGQW97QmXcrgXzB7JntuYUWy6qlypDAg+MmevqTem79JaPN
wUE3qdmwww6rU1gXIEfvbyP8tpZMcgtNhkdjqRpP5q7bfrtJwVw5PuVvIf+RJjrb
ejrfTHYpZDhqlO3eWOf7mn8h5rMl8WQRZ9ov0HQUWHAws1t9B2MTZ1yjrH7BwYiz
Av2cXIrHiuhwq6LhJ9BtMbec/UrgmGxcyx9QP0Z9s4/t16Aaaodv43hHyALJP7Ro
DxKhhzP8K9wAPrM//v2MuHXliv9jd6cyqHAtvk0fq2YTofQuU1c8hLz5E68vVQDl
ZXzsOCJWIlo7vifP74Eq771lXh7Loi+usdLu72Xee1DWA1TawYyKZK4xDNdGkn12
x1Lkv9IDLys+PxlyLoFDSQPONPB4N2JbdhdgK54w7cRrHLwNQ1icRnasYBVhkLbm
gGicdyJibK4+mxS/NqC6YZotASToGjh5UEV12NVimfvmVXDs+zcPugElxLBOVsRt
aERBX9shWoTXI7TYkXWbQd8uZC5j4slJcapIbkpgBzERUkJ5fo9ac5K+5z6uGoqT
Iu6ncw8QXAIUMF846B3bRMkrw2WGzDHG6KEn4K34o49iiWspvuNFOY2ZmXLitVuG
pPN3h1Q6+B3z/O2pSC6z/1nio331QaNBT/OJ6Ke54cndp4upos9IbVTdnB5RLBT8
GaQL/Y/NXa7nAd2AAdXk81RyfCzeJjmHcaJNE3KUE97LyQyuOwknuXvvfv2wsKXZ
70wSTLp8wPZNNFt5V+4gDK+vgdmBQBFij4PzwuVRSEtQ8WweETjj8wSV8CdpoPyv
CYvdfkNPmEF9vxnsnYJobMLBFX0qvc6ftcZj14FaGawg0uI1Og05WY/2F5V2gZPA
IjGm75YKyyBH3lBuacujkUzW6532Z0qEt899cC4wqLsO6F3HnzEsAp2BpE8VVLx/
eaekOrQYBOpNrJjULdEQ0EzkiKReYxejVsT3Qdzx2l8RufwIcdyDO79Tc9u80ARG
thD+XvmYeSoSzdnw7jgiTaJS0RPQkZOmUt9qhVGcEgKs/Sd5/Mm/pnn+yib8udtq
sZx3MyxDMJVcpRA2csoXEEWGE4WXQGBoAQuSRGodMpilvEOAryCib/SNp7mMqj2g
m7jn/BZT7KZC8RoEW7EEVH96XmD4JTdxolOptUzrVH5S9zQjDdbTwlFKeI/KkND7
HkJgB+DC6yy3hiWA5Ykp35CCoAYHKQ2btwrXmZGiXUYrylTvP47CJnHKqPLqGXE6
OiqNXbFWw68fZ1CAasJ7Xb9B7G9wwVcQ8ZjBJMtQMRD6uiPe+4vZIZL+ttk9Xwzc
s6yq5TRCik5WVL5IOhgfNppk16ePJOjijCXD+VWVxNuNeB2oqrrcAS8ai71Gl3co
56yzGSiKwe9PWFEnk7UwLdkzdcWLUIBuJisxFML+PoqK6xHtK+8DWyJQqM4Gzrm7
vgvrIxbVFZXiM3BYKyeSlBgGYcwWoZx5ptBzi9DcAY6l7OebZPSUue4fHCmP/eMn
k0+UszGFM2Bct5AHVBTT3KgOeitqJBVp9YKBui7rWDBYhNwOqh2l5pSJaiFQMEG0
kCtfZnV0iZ9es3c+YA51gCxpg0UMxR1ykAMr24+ur7owXWaai2EhEwnFs5NErNZr
4mhfgHgqmJfujZx9njgQem5uObAPrgrgUE9bXET8WK4qAs1RfNIzpnq1BFLyeFKx
squtrdQI6lv4zCe2ILKjWhIe2sYvIlNLsVZ6kVwKHIOcT5nKHJLjzAV3PMfpntTE
5blgakJ8GIhUsKwebkzQfkvceQPxV6Jw+17JnlGHtNMQgyidVTSg/ahJUFHy9Jw+
hub/sGs3z6cBcMG6O34fEbVV+DILxSRftYMHbCPYlLDJvPJMqtjuG9CSjxgiDVlC
OpvIQmy42LOiCQzVdI3ur40AgJGP0/ZDP5JYd/oO6zjMN9qnAjvVqgn91stAya9o
DXiATKaOo9qqXMFoK2UGp7VQ0n1Kk+NFlpDbJQe197rEA4eupGbEF38see4E1UoR
ucOd2xVSs2m+qvEnyeS1asNscF5BTGZtqPOrZ1PAiCsus/zrfcBP2FLapQo+Pdwz
4G9/pIbcO/ljOIZ4XGsBSR4XSyCP2KV+bm2pb2PUcq1Wh33MRdyXswHSImPsF3PE
66g/EOyGd6PD5qzhCvdrozQtbbRa5LJL4kDhN/+vt5DmiU2h4N5biVSGBVj8c0tH
tEuxFoFCQL5MJEkCCDrYxysWWpX6zzD9MXnzYT1YDt8u/rz+4jXiV29bjQ7iiZVX
HI4cBtX1qAtEkpEXtK57Rhb88x4h/DXe1FzUjQaA3rZjJROcMc56GjefuUINpDd1
yNbQWPh7q3ojIpm5LK6N0m9I9I84q2BqNWrIDWk5EHHNwgelMniTxZ2ztUld6DmR
i4DlygiszwlKCdr+q0LSMJ/Pb+EQqxPlalIu3WrPk7Wh18sPtWzNhWGlEWHWBlNZ
Za+L8bqERQUhk0MGxwHhYAUf8m4B0V6ktRkawrD8Lt3FS2kFNfoIKrbDRMtkJWgV
BeOtFO1Pmc/jKvXYnv8d2y8oUZOgWN7q+JpP+QLbua0guNdQ3DBSgQLk1XPghTsO
oxjDwCSkFJmqSU8B4kcA0KVQd1w9r0E7VmyptHI/eETYIucwmYzeAzsIqWsEN9g5
YSy6j7GOWnqzQgr6gOgBM3oZofOm0038/M6Vtt7K+bhey2oABzW7PHISR9tzwzFL
iTvLVl54tPDM8omIiqUerz+TFBO5f4o2tssI6eom6u3FLMf42k5+iF5nlTVFyJXa
A9qbIp5hgR9ONQUJkO9UQveTfjDS0qTZTjylfz+XJ4Djbzv16e3bQE+IkbexiPHg
IuRV+rZp44XLdvaFZAMi49CsfpK5BdMxaf68ucwVkFiklc6bKTFtnDwboo0UTl3K
Jl/71+5Z+yAY1iG2A0Kh6lbeH5HJizEIJi4HKAOcmJ6+oYv7i6PRgOjfnRlkGGXK
VyPNj1F6lr4qdjQD3xVMjNVRsr0GI6w4lLlz4XMXP7vZrICdxgFKFK2FWFSMTAhN
NP+R5VoNdvCLLqdevdXGGCWoG/CEs64gwJWWLDucupDs1/eAamsSQsy/kt4zBMvl
Ctwn1vpLDHPQOe5kKOnYCyiLWlR3EDuPt8+CpUvkulpFLR9WEe1Zs/ysxSVIoqfL
Fq3K4jQ13jaXdrLUxBsgg1JzPKVGzYDC6AODX9Pp1O6/m/HMka5ltHrJKL+HZO/R
hX0jdZDn6B57A6bW/CF03rzdiYFhnkXqOoio8srE8d9e123mSXtoi1UgJCDiRsNw
91a1VrrJWS+YMAt1AD8/ixo+n6g0Qq9gQMYhz7fpgnSxZmLifpnY7/OdFl3uHJAB
iEa7wyD84FXP0p57uNz8yUXtUqNvYr3odEJmpd+U6Kce1ir2aNW8wZph3D/lzWmL
J32MIfB/s0HnDjdB+A+6kd8w4q2/GRiIPtofXeZ4etP8LmQGDksxnwNAa3ue4HvN
TkD0++e8+ITrLZ0euBXQY0pAN6VFRyEaXoie9mx5ErN9abNC1VAeltDmL2SG+Rnx
sOFQOt7r7hHW8cWmvuVcfkzk+ZE94x78SrwEbl8TZR4/YQGLQRIZalgrcwIqjxWM
e/CpiG8yf7G2qKcZDF4iupwDqmEpagFKhAG++FKX6ylc+0yo3TBatC+zIvKsBJg2
xTlkG5kv/UzIrPBC0/z75quUb9qprQga/heS2VS4M2RmMf4Aqwslg9ncZayoMLW4
FzsA1h/9OXaSG/Dmo9B/1Vl+LYP0Npft3UCS0hTJuhIGF3uNxdRzYl1RlKCeTCgC
HMu1fcl+bnuGZzPyWcxLSI1uh7xWQdf/q8acDVYohY6+jfn5c5Bvt6300LZvCT44
j9lRtwcEjjlX5Uv0/fhhjNS5B9JH8KyQUMSmIa3wo6FveIAiukYnHi5s/qxS30vE
/9/Lklw9kL6d0UI6/BoVLh++qq6zytuP4Zzd1zxVKm1UnCnMRtAuG/RU7QTad6xW
nmr/UlzEq5UzhvxzC8Ezowu7I4vas3lryUyQqfASk/aQFiqctK1CuOKVDuHfnpw/
GlXNqqgnNmykeu27gM2i/ad1FRkthfAZSV/PwC0qq9ESnL4D+He7XBQ0Ms28sXl8
0GW9h1s3b3+pC72dLeswTDs/ue0DIG7kwMeLnAocpeZez91GJgnVhwvYW4lQP0pv
6tLq1oTxSa876tZRJ3szY3h2HW9Ib2N8ZDMgWfEUk+eWq9LGHAEZq7tLdwp5zG1v
kqm2223sGsB78BKMTbVF9hLrt70JnFr0PYPdBtNAXC3+UEh0AV0PuDhlewGQx4eO
/OHtfhbhNlHgiLUHfuVT3ucWNf30nOPC16aIsjXyKfGY/M/UDEIkuUz7tAW3GJgg
XHeLJrvscHNQ3+omhnFI1lbYbpkKxcYIlp3oUf6HV8epjdo4snAOE3n1MsWZFphn
eInd6Wkx6iszv1lTHVhzc72Vak1MQsHhASwDJgrxXK+KJjvU/xGUVCrXIu+gnijA
v/vkYoMt3GWlAWhc0F/LvI0gkE9iIvDhLcRR0XfOIaSsiOPk405uf0XDMBEIZuQO
0z+ATDyNOa74UiiD4CvPU6OkLUlpOcWMBG5sFIHkPN1n3iieYFo9P366/E6iRcVc
nkoMfPcxsmtBO+adefZLdxsCBDnfsMJ9LoMAaU8DU+MomOZkWR1oIpww6yT4zme+
0UdtfZfTHKigoC8VSM6Q0fOY9mtHee7mXFX5IH4CNlW5OhHSZjwNjIPj0UQNAPQh
yxaA8Nj/8ubLQU4Jat/K/KQFwzwPE4Edf/Rx3cO3UgiuSvkxwcIX05hZg33xz631
5mT08ijH8r1nOKo0Eq+xyGMpNzZRt5eSRf58tgljGMiOWsighVrA/UwXmt12kh8e
mNgQxDJmcbyLeRqsYgoETr33b4D9DAIFE8wsic2vx8DQ5rj824olGPQtSVWuhPkM
kvoS6K7DqGxjtiI2XPYuL1TKSe1WevJC+yCdSDNFcw5AwmZ1KcUjoSG+H5PE5NxZ
irWWw0cFwM2AaxQY16uXLytTr4auQDSwrvNjMsX773cgQP61hD2ewaaOrTAopTCt
PTQ5EIMBr+68YledipUK6Ml5bxt3tK0IcWt7lnrh/H7ueqaszQepyc7P86nS0eYq
0aqpiOvUgF/nuKadTUKotrLApPtMZzik5cK8fQHwLG8vMWrT2enjd6RuQoOeYBsJ
YKTKAdDsK+YGeMswHaJw6p+hrOHPkeW3ZTp7FPlc3QrBYewCTCMU8/7r5pFlBZTD
KIlB/BuF2n2y1/vOKCLmVIx9H2iGf2ZbVRcf9YkoTJ71lTK4EKC4GPTaYL+GxhHE
uFzt1iV//21anFtTSDtDLbZhIMMaB+75FRsBfWXOrL9DLV0JohdCA8sh+YKwF33B
rIO9KtCKp3MUl4YbP/k0mmsqnaRuLgKcPPbzDmge08oAxmRAvy/f69zDJs/V7+Xb
12VYz+HvrgwUDGVza80+Tg9RWPooMgSYOxY1P1NCh/iHaQR+u3WM/F5JIwyOkAUS
bQHZd3U62Qo8AWuKlG4YSNcxHtdPpDqt6lhiKMfm4C0qZcs5w+VPQwE971dIi2Kp
JbQOP1uMd4rKPja5m3n3tLL6C5yJazllegfCgLYm7GbHcdiqHEMPCIxSNqhtdDym
FHiZDhU0WccVS1UdxEM40rH7TXxMsbXGOZkleyUrYGpAfLzj1EqfLQlgYHP/Wuno
RZKVi935QFB7WM7zHUONli7leQu/oKiedY1ZasOzFwXmxYvD2Y0Kn3uYni397+fm
UHPI0LmZZiESiHGNsVodOEaTNeyzB/50xZvTKFzjB+t2xUmelZEIgkTuI0NgQMo+
vubgNTKuOYNh27Nr/UtczaKQ1Mp0SC+tpU5jeMzCNzEwQBjX2EYUi08YUf+KxQ3C
xlndFAm5qTvME7tqj2bwApswJSrdgE42L0ZB5QkoLG8pHxQoD4bi3q7KPOgQlcHZ
VpxGZ3ZwQtveZ7si98JYVrbDXuwQg0l60gewhJJlgNqq5M95198BToamXS+4UoBi
GBpAQuWtppo4wtkfJmXm4S0TlOzWZR1l1ugUkIVH6SId0Jhs1Boltf1Sy/6dNU/8
xV+wtg5UOQz4uv94Z4SqC5SfCrl316PEis2AeZSVySLIxOhwJuPoPuYZYxP5Z2V4
1zT7GiTPeHmqcu9kb4Svo1xHHIJQnMlrXAd/yHfMMp6NL2oDU/uKuLDT+MirqItD
bWw6WZc1mtpet80B6o5AG7HrEHeInVjX55bzuStTJ5BzijmZ430oQT9fVT+/s0Mr
fmkSAdwLkudsrvt7mSlCg31pJeZLNzHapnDVjslFBl/9ML7uCG1F1Hi35R4mWQvC
SvdMDpQRHhwA2dROulnhkUP4M4iV4gI6nAI9s1qyiDef+HsNzo5bD0CNsCmwm5At
jbP0/lt9WSKjl1ZP2kxpvAVIukmKFgWhNe/bCto/Q1Q60RLeiozQKrqq9o6baNQo
ePVVtRUBkaykwTBK243ZyUe9s7dLluvexlNutBzsn6YeO5c9u/pdSjxfa4L9uEn9
kvG9dzH8+J3CNFxuPJ3Orb+RonVUrQ7xflZz6wGDY+BaheIIzkadGTbSV3oF60fg
C9IP3bA6SnrIgaDpDNfHgLALjOM6G+J8Qh2QSGu9mOGJkcAhpiTeyzM1BkhsRSPi
9uaIF2VLdN6kximDZK/mM5MoEusBNHCX4ygMvDcUR5I8boFeHvk+mB36LtaIWCrs
/cWyYMMis4b+wPBPUbW3i0viAnKP+HWYJs5aYcuQPkaHOj3NgJM9msAFGByBGTK/
bgnVdbxnibVRMkITfod18O+b/MKK2RyWBQZysTB4eb2tfRBWOz5W1bJS1LyT6k67
bLPrkeNWPaTQkE8bbdUyHmdNzqVnP0oC9qENHCanxZB5RB36XmCAZ7DN2Sk4qecj
FiSHm4qhXTUA3i+1uPGiN9kF0AysgKQuq6tPw9uPUsWOSg4CC8X7JDEHW67mz/E3
ERh4giwpJoC/gJk3yMfGVav2qOqUyTwiNESZ2mlG97qnj6FZBPuB9ulKEuqAvxKT
yZh5IQlhWRjwML4gesEsv+H0+EdDafpSNMwwwv5odBbmIUUJQidU/xwhE25p+oi9
eo44joF9685HRuJWqMdw5+ma6pN+06daMNhNb0/8IzscZMlQ7WM5MehKko7SRnLq
FjIGUS9q/hVx2BxHdX4uXtFXk+FawHW+Q3nI8H/mZB2dhlb/Gfb06aXqxdg5w3Y2
bO2JpyE+EoHxsZ4IPjciQnlEWOLK9QnTz84aIvQ8fo6F+Soe96IKWzBlQVX1Jvx+
OxZ5ETTs3OZn73agowbvaMtdJX7zd/T2G3Kjw4nmhg1li7QgR0iJIgSwjk3LqAfx
fHjZiCEod+J3Obj3Slu0wPnP2ouLb5w246Exs1dPTcX67MEqkosSwBnkHBw7ZrvI
C6QbGa/0SRzwhUpg3W3fs4hQqXTvKjuvhmHeElyRQVIIK7Me8QyKkYJx836qB8wE
m0+ONhba/NesEnpkFuPncoUEBCph/6gUbvumGFRoS3Vk1OEB8xjaKJpsc4eOdIPV
vslNgLjnLcVrAOprCkfHWFdyXpWj69Nk8cxIOlxYBobmlxuA9+AgH8b+Z2V9bgbA
SIJTEL0RkSfwRSuXzvf547Ei/FJ33hhWlNjA7qM8lv3Nj8zDiDfXwQO3lA5pGudn
jzIJZ9Gkirw69LODf02FyvFKuWEesOxbMjrAbKq+sgI8VexpNHhccgLQIVWwcoTZ
pyDaRfBaabhhPhIZqUqlwv7mIhJeqWLqwuDvpqECjJOIKANSwSj624zPi0i39rLZ
Sfpqb/PbMujj+a4DEwtuTrUHTiT4iB7KYDKFV0KYm/waYCmNdQA9PUJcZmVMOOVy
SMovOynsmRZK6KCEoJi/oNM+DDpzM+zM0oWmX2qeh2tsuj4xUBj/CBB5QFyABBug
fAmOA2KdTRgSqYFyp4s+0aZpa1lDyXJpZmegMmFqJbh27ouFHijsEbsbiuPHgjau
SMPTC0DTDRI0aUJJG9ngfQyPsb7cDsaHFJoKy7+IRlG/oMIa6ltza+H2KCM5+LcJ
pn6gne+GR0o7u4D9MLfzG9FNfO5CG/gAztkvLonepNzO5jybvBVxO/3TGU2GNgdu
XWLj75G34dWdL2S1XOZM8KWcqGsK2DP3W67TTkxZUITcSGUpZwzwg1EirYguYsqL
nNK2QfS0xV9//KvCQ0rGznERd0bB9yKCNc5RqaiDJ/de6jsmHJXG70lPmyQbqUJA
qG93RsEo2LDZPcJFORbmiQq1YvLhrIWEIOuFXxB8I2FG9A45JhXG56NnCi+8FYR2
kNNBnNbi0iYadycSZ3uJjvU+lEUG+2Esve6j5Sem+sIAo1MsD3In7+Q2KIDQ6X1T
Skw84i4Q4L9QU2EYrF/TwN0wLc9RvKYJNjzH6pnL2lWh7+5vGuDRQXmQNHCf381D
kt+i3Rg0QvyAkSc79YIRxw==
`pragma protect end_protected
