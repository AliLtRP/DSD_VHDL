// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:39 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
RHhivzMMs0KvH1AlOhJJmr3d/2YziOmbXFQwYwSp6liEM1YZrojdO5rvlNj7ox/b
WTxZjNCue/3m4+m6t4DfGjnfIYvyxUDTbfVrhsrnO5NB2ldDjRachgSmbyKxNr4n
xmFyTadk6PP2wqnKCgK3Mqdmli9ZzgMccaTI8gGHVoY=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 30560)
/gmIK+fRRzn5fNL+vvTwsrOv1BqJIdg5mHxaZtVN7Mu0Gc2AXZSq/WWXaKte5tT+
fbtEYbSNTp8bHM94u5ePMOt1QG8Ri953ymr9eTb5LF7BxpAYEzWYacRLHfVkW+h5
z6m7wRmOf78XnrY/R7QO7RStX7FyOr81/ZGhCNuAB7M9By7wpERzwYAPyKF2Mukn
4ySuOmAUXDjf6EJ14Mo9ababbkkHWvLwupzIGT0zSJovc0Al+FY53+tuiqh6CtFQ
81sOEFTzGoFD/qduZqUA/0ya3hdRY6su0bT8dImLG3iRYyhrVFEQvmdIslzqY0fC
mbyE1f82sR+V35tSS8tvRKTbEzz0k6Wu5kOVYZb4P/KOuBRVr2DS5N53WYN6kzxx
9l1UJkMABD8A4Lq6k6QPyYvLkBePj8xO6HzFP/hJKRqljk2BF7PPJIfFMNrU+6Ya
+JYoS3zNceOmxrmIt1gGxy/PJRkOso/qwqbhC1CJIFmPQtkvNQTpBfA4J029AwfM
er2NJv/pYCdB9bxnZrGLRxMn7FR/IXxf3KdIEUl7zYJTllPJIRduK/dJAuM8OVCV
V8Wt/rpTRKLMGUybZQ31AjXR9xWxDb5XZcTSynNd2pVno6RIPK+4L/v4hXb/UujH
ponImg2tjdNHXibM83rs3Owc9vjjBaRVB8MF87mApHfZcnCwgNNnWsdmmdJqx2bq
+t5qXVgYyyvkK/2zb2ogrVWLZT3AyerCguS+rTi6GqfdyMft+MW+Lanzc+Sx5gFI
GAIfuYFBKIwIadtJcmpEUdJc67nYso5wgy4dU71XQ4aGNulA6Pix4GiKa9+MpJ71
+WiBpj8aGAomzaXvhjRuGGOfzeLzIqgupgFFAMegD6tJmoV88exFoHnp9bYWCl1B
52R4BWRVGvbvYoLsNLzZU4XdVijy5NdvANBBEfX8D64gMU2p1jcXa5eY5olPcl7/
T/rNQRkpSmaFUVUF74OVg63taF8oSHF9BXTljEv3+TK5A25Lu7Qem2J5y/nXT4ei
UZW1+XYKU4TDG6t7zPgwB3d+6Hfp/U+cPyq8A4EevkROGyMYKVt6emR8errBjr7x
JAlaXkLaib7y2TyWjsaEuKxToY9XMG8pUhrEulMmAC2lkYNe5ii/we/gQUOEVT1B
jStw4UwKG9pHVPu5D/B44AvBHq8NREnddT+VTGRyraRfTgU4Z3R3Ju9pVU7xtypu
ubkozH2kqrCRiNNQLOpDdf5DU1OdfpXJqRtHpVc5vgFwn6CLobC9tgOx0WqCytA5
Bu6IxFtsUVk51fYcacpm9bd1v0u+ubJrSDhXedcBd8TfSgcSwSzQFWb8f3qTyiby
Rc257Rk1OEqc+sc1jpGl7jV9qyqj2d5ZgUEl0sDmVrlc1+HPaF0gZ2D8m2p8g/yg
RmQq1dhisJBh/RD9ggMRjn+XYHHJZP/DmYplsDHpJbYxBzr+4kAf+CFSf9gdmuSk
jU5VNmTqDaOKtxizlOo+0ILSSRobcMFZ2OD7o6HOrSY6+6OnMoDnWPkpB9ii1BEs
t+neiQRc0KZ/AkVcm+SmlJ3OM58iD75ZE4LPZwyVbC+FeslNk4L0oqVRvCqxaU28
+KOc2NDo+Q13Pvqjai4clJr0/AS6UZpPLcwjo7+Ae2n/IgtiXu8OG16LaWA/hlLk
LOWDE2zl4MouQI/2XF/hAsKqq7+F0G0Y25UwP4Eua4WfzGyhkD+GFNMBFqnJyWpB
/3EKEB1+lPzgSeaSPIF1nPKCRYpb2wzXCmZMm7PWnGcwlY8Rhi/j0Dqm2yLgntWN
JnwWEwuMq8YigcYMYgVuPUDJ/NPjeU63KrLsPEOeZE2BtMw0K4OipQA6YAZGi+ji
exRWCs76S3WaaijJ/1sL7969PFUWnXO6ANcIIcZUlWMiGuZY+j6Xh7Eow1XZAUJa
r5BUDKHCt9e0wXJaPiS4EWNaezNDCcwb+D1DcpupXoBiHoHEEj19PeL7fZfuWm3Q
6lZTGyfKhZoMVfe6XKK/z6B+i+swEA+5l5xezLuSlYhyt9TeqD2LaKsloZbpWGRD
H8mzWgr2hgV1ibpk3v8rsk8Vuhq5AweYhcdovp+1RauctlmrJUPZQpmNqcUi+7Lc
L1ZjHAaPKtZlhG5fPJfnnuCP47+8ErDdEohs59sSvYiUAapUAOzUIEGqTSOHevl5
7mGAvNzLd4R3hxfImbKnJYdULLoofq2BB4iHhQvsIvUrbc+lnig9v85mYstlPwsN
PtkImWBIV7copbTs+5LRzJWdOSyZ+g7SWvPIPlPu1A1tV1O4lugNQY/3KrifuwAl
A9kjpNod1jcQGGtQs5a+LYgz1jZgX0rC6x6YyfLxsOdA1gzMDXM4P6tc1BGQyMX7
yxbRlbVVPImTFJ0HYR5qlZM1sff6M73aFDcEaBCsapDb9UKI/M27PBcMCmCYWShy
53cyJUPRVK7IAzM8wsHr3Kvh3Mjf7VMGJPTasfjttqdKg3jHak6g2OjXfKGoafA0
S99pRT/CvF+PxYZ6ukZlNgmJm9s6Zg4VcU7sjHPTHwsAoG/gAyQHeOo8WISyo71I
lbiob5c0cWcS3Hrozl3JztHJSKcOJmP8yLBpSMAiFRgaoAPZR+WOdNdmP0V/GNAv
jYiPOce++xUx2g5hwacei4mKbZL2yzBwWiG4IMQI4KjxciAxGFXZ7ZJvZeDYORTj
I5S+gViPTGNWkT0ytFO1MROtNxySiiVP7iP1DcUfGwhb+Qu+y6L4V5lj4KCSB3x1
F6hUqJgcXhnRgfn3t99PD+M1dKPFUBPZ0RmOca0LdHAUoSRzDQDHOHk2p7j1XezP
7OnnQTDmO3muYwmDfKVflWuMXNRGI9AlDdu+PvlrLR7ABbLT596UXQutJMnt5+rt
XHLnRXAe2d9+llo1VEOWVIyqoQxJBpW3QbRFAr7uPhxQQd+FgMNW31AA+iQPYsfv
6f/x+3W2DJAsfFhJnEYdLqMmC57sOH2Gqnjs4N8Ilwyjx1MrmjJnTqF8UAR+D3XQ
LUYckMF3k86WHv4VQY8eWqkg2HMkJ2cJrp9da5nDQ3HwL34eSol3UKe5twZlpRKv
9mByl79zHf8x5r+FFjOdk6r62bbsMt2aR18QC8qChIPprpnSnm0yihKka9YxKzWG
TMIt5SzQvlbYFzkrD5+1rTMgY58n6bC2/CJVdntnjaLSgxCDsyaSbRZCHuWA9FmY
fthm+8Mq7Bw1rT7J33Gq4SjTj7XBPtoh2iN5HVj4H/HQK4dqflV60ZaKkTyzW8Cu
TO11haGQen9QyVcaZgn/khOB19c+PwOM7qwwJ4ILTQbpGAU7599J2uMPeSSfDJMF
Ii8QGwXmy1kpXEl4R8OxKa+iMYa3wfcveS8USZRowf4/PwD3k9CaxEPqXooa3uV2
DjkaOtzpXuqszXe9rGpOIf2BGYbmgiSHvySm+45TsvAduIENKz3TLwPqIpMfWxer
wh4JKEmDnl+P8HCs//eC6qeD3l8+dxgYRdQPqGofnw/dJDUa6LNCcVq3moTAD0Dx
2vkzzoeFp1Rc9/HQuZlGYXQpIozGWprexxtdOBm3O6lLqeXUOe7BCOLCHDZwkXk8
J+CYwqzBE/8TfkZQQ0BuIbBylTRPWohESAluztavby+fzRXvr9FgpxRVGC8gdHaL
hCe9Wa8d5b10DByOR3JKSuXJzpOUgBA3Sr74gQ9GINSmtPo5FgwybOqyEF7eul3G
fH00cdR7/M7l3jcqdaRpBmLwRrpD1PFupgyy5kIj7sF2oibkA6bjnY5Eq5+WnJiw
sd3uIJc/936QfVgB1Z8P3rPjSQx3mhyG33NwaJxDVhR5GBUKm6Ter9pd75aP+mez
H62rzpu6vD++iPIbkSwoc1mki2N3hg0mtAvk+9cArLhMGz3rtgFlMUYyfJoLrCyo
dH2b9jzUH6uFDbJuamb4HJNl9a7DVE+f7QbMBYoR9AnDzO4V19m8RTVZgPCDPInU
UWTCUAp7AejA8crOtxGD2k4MoW0AiCBhy3oOwXOnX+OiNt6cWuksnN70qIxge6Vs
EJRdfQOaWaxbTlbP6UDAhfeE6bySonJyki5nWzph2nKOtb51qAcyIQ8Gj5kZXI7O
VA76BtjHfzHUhFq+vXtf9eqhFEer6dgTnuDl6txpd0Q97S0UI/JvN9iWiL6iiZZW
DGGLDzW0Zu1SbmQw2NreV+t2DfSWkP6lODGZLZ+PYWlYG9TrOk6YJ+nakNonj0jV
uUy7+Bn9EMGAEPnmg4pQxunMDJHm+QaDRLfo035FhJCyFQu2IynvySlgC8hVPzXq
5wyW1AeArAiysqNB4/P1CMng6rBoWNu1zptqhCxJ19dEPrmDuBZKfybgHN8ND3C4
bjGbfHBkYiVkjUsyCZOqmRIxQc/ZuSC/ptzeXEidQarIQ71F0MfAFdqu6439bNop
KCmcC6bJ96VPsSlc4G5kEsN3k6QT9zH8KF1nd/qkc+UJQawWx+ZoDht7PJQIxnW4
MqoyhsoXNdSJBeXZM4giZdojKeS2HIpd+voyUhBjrsIWI5AVVlwrxTsimJ6EaNsE
Q+f8Eb/6+oxI6LtbLPKxZGdBvNiVtZww2VYLNpKqv0xMZXYJduIYrZfIeVjCACJV
EGN1RdyKFyrpcCT1T1uIjn02DiVHJWn4aqNUgqGTUwMZ+1dNRzfw8rh7hGDDnt7+
yVsyupy+mtyqL4PT0+wO8l6yVfDzrTODJMtL2AXdsyP938xx8AaX5YVRLHD4IfSh
onNt4Q9eY7ZhsXhZZEfT00whaIlYMEzcOpmGc9kCP2P+q9XF34I+0JFcmVyd27fp
ilMTvOm9T175fF5DCNpepVEyg1zFe+va2C/Evxby4Iox9Lrex/7KQwZezV7Phoax
YESrkI6z4XdqOtKgqEvTuCH5eHGExPZXObH+39pCK8surOZtMbqSl6TqI+3tBO3F
SlS9qSMVpu9NxWqknHv67m6Aw/hDoVBHltnWU4miN37CnEg1AcIPlA08YnB/yx9z
jvip67ph5m/iGZHc4F3DbWPB/hTEq826F7vocbxlfkSooUB20sUKxdB/GzLiuFAb
P7zxArq9dF7mUW6Idzja6hpuyhUIsNFo9lCa2J32D1CViwkzZ6ssgZufmwKInXhq
hDoRdEkTIlb7kKxamxSd6fuQ0MWNhUrp8Xu1ivBhZfdLc+CjIVBsJZh+s8XUcf5d
TA+W3xwrzf/rf92BcO9Zju5YIEbFeW6Q6vOw3H0dmGDZ1/Dox1Y30PmgbnEY+2jM
/Dr2Lh3nGGGvEupYY/ubhKtFche+jjU3JyynZQrdtapgDsiINPXaimk0ZXJo1ueO
LZE24WEXjA/+DCez75s+m/J2oFCMDb17frzWmJUNrtNk1mguWuTscb/454zAh7kI
Fl7WwmLiN4XbqzsFu78VVoYKRCu7AdiR3ErC/GY2U3ZLdjiu2u6xa/PgUfjBQyje
4WwcEmwrnkJQ/lUa17p7IDia4n0W/efeJeebbc1mmPPr6BqPuRJoMFR9Pek57t2A
Yzb2mvT2jmrtLhe19gJogfqVgDiMIAb/DGEXiHYCNDCcUHSeSgQQdIg0Fo0ixd3P
0NfzsMxU9ZY7mX5XaLeV0eACkA3JuXwqa5HJbx4B07xi/JWWJF/OQEK+I3dy5XtK
UT0HxlKeJr9TAf+0WLbi0nyJKSfJO0fUClN3qJPtE9Z+cJodJJ0k0VuZ/Ouddd/7
DOpxAKX5yPVB4lVff3XmW4RBbhGa5bNDBiwkvddGZjw3fdnTg7Twtd/szhvye5Xe
TcQe3xZ9gl42obB5luO0mWgJXf56OjEz36uliLe/mWSpvwEQ1K6tsN/x37tPPfDw
vvgNa4P8hD9DUkVr9lHZM3G/8x1y3aHhODygWcFr7oyQPgTOQdwsV/+YlCW5QxTD
dkp4texSY9ocDZkS0MrvSVoItFgE9fSfwFMh7o+86NDGYoW/UKqzHiVlsKcb/4HJ
UB3+PRV9GocNuGYVnzHpamzpX55yJSCAkrlWV5hM6UMS2mv5J2WvhMEJMz+gfpAb
jfkp5LZ6tco3FAG1tw5HAWMuNzJuact5tKUGljH3BHN0HSS5ybrJNhQHvoMu0/Ie
K7fNjJCmWAhDAz41e+Z2i/4ebvW10I3Nr6slS5bT7tN0HtvO17gFUN0SOxLOBRBT
vKjRSH+qZAGJpYeyTDXdZVfWPvNjgfHtMnayNinDLKGSoE2ewzw/qREAQ8yNumFN
fkdzkSSZrx4FWFzLVGIzYfd3v/ym4BAt9AsmgmieeVQnSdpVfM5mH/4XOppd/7DH
GQaV0EKrqq+jiPBi0bi/dJmXjRQGPaVep5UJgmnCU2YHVodonZM5SmEaQ/aVXCFl
Hc9Juz+jv13dVimlu+/hQnEc2z0skrni9JxxmUef+1uygbc/uzEIzUGnWxc9ArC1
o3zjodjEbPe+rl4Hhrn4Xd1IlXbXsJoYwqH8JG4wNoxJcazJj5sMRXJVpgU9cL5I
zIBXscCNX7+HCTKhp4Dz+7ueJZOBfisbqKbx33j+9zyw/lU6fGjAY4R1Y9Xnf/Wl
foVI5+L510artonB053oshvlOHWl2V0tbcg3SYx6+ujMMwK2TKRuhp1JsxOPjy3i
k5JrUMezmH8qViBMMqMQdgw5XbS/3FYbrTPABREB+SOELcBwTQ85H8Og9mm3BRoS
82PdeoME9i10VwTxIda7KSteQJ41RQbqWg6cji153SwJhAKHTi3ybgu4fCeC7hFe
VNF/2Ig2tdporbdVHLcgs3x79EuAuY1PnJ/HZoCNileW4bglMEtslSt5ycBjj6W0
uupBb4qRhh+gDPjPVt3eIzw7W8GfjvDhGoNTpPaow28s9czR0uCvVaVOGpJRD5dR
Fm9XhnQ9qN6Ckpytn5hNOywJ3wAh1dtTDEgyAgGYfd5XB3SSK/wqASsmSOS1lgUT
V1lOszsb2Ah7oKShSFhxFkBK26pRixTeyhwUdE7MGo01DcxnBAeGgRPPfpPYmUF/
amCmJX2w4gHueyq6c7HCNk4y/lwVKBchx8Kw1TD4JgLmtS5jHjA8CrCu6Zipf8K8
ayMW2BX65rUM2sLWOmFZG2YdLS07+tbcgNvVtFEvZQFwcRhN4TjgG6/44Kmdv+e9
8mEacnYLpPqCBLuUwP9U9Fc5DdGEUx4v1XwxWatNYf4MG/Noo8FjQjhCvcq2s1/R
/eYgBIOjPNQ+KuDDpAl+ABqBX/yfk5ic+ZDiUB2zCJXC/Tb60co6d8Br7JHaj6AU
3pARM2mqV9bOJUF3ZQNjuHzr6w9KzPfMooKnqjWQ7Xl3S8t79eR/6hlQVKm6wzZJ
8V5dOxgC7rWE67U3xY+4Ew4TZxBGlhMqkNBxjJnjTtT5E0Wkfa9snQVkA2PoKb60
xPgjPYB0iE97HyobNlzCZCZBwuz3ARHxbGUk22OXYTG+FLU9sIYs2eCfTd1DWpCc
7jYO0JpCCY+Eic+fr20WjefzST/4eqPmdiA2b55+qYgdhvzs6IF7vTLT/2FEvV8F
RwCM6Ey8Fb9j5jR5HjSPjw2C8ioWapAvxO8rSo69UEikGZ6/FEUBqqwGngIgg6NN
1SS/3qcgut1U7P9gZEQVY79k4A9yi3KPlvz17VH2LdJUSj+UJvXhgJtaZc5EgTz9
Gfo4EtWtYHMPyNhQ5mkn2h0J4RoYPAykYFr7X8IJBw0Y6M04qAy0hv1mAnBgonvd
5Fenlb3S+FEXTPR7AJ/aRPi/T5Vjd+r60NVeHu1sWRHskE70VoXQ7w5RrHNKyj7A
XmVHBJvoFPgbQ74IxhkpFDXHkcb4GGkKZJtgxrNPolncb2e8S0YrtOABjobRDHSY
TVJWy4tS5gvxKORLjNsUVzbFoQ1Zv7T4z7tR4Qp5Xuehx6tKTywcbbf1VNNYvwGj
7/tXxCc6hkeFRyqGcjGhvlKLCDKU6EIxmRruXIAn3HHSAsUQORrVJpophmesxxCs
/yh8t5M3XHFByiQV8Shr4PX0lsD2VzA5XZKZOKFjvvqV3ICuu9eUNn/CaYjE1M/y
kcmjaJISvURxZCfsMIYBdzZPFocExEUuhaGClJKCqHE1G7uM7HzBJww5D/bnhvF2
nO1IDHw/W5ekdchBsv5wdpUTwbe1FfnD0Tc4msqIDxTznzNVNPwJRgaHvLKh34tm
OFCwvZrxZPtyykOtzHgBkhE2PMsp7hSzlOvXpM8dgW76ncvBZoBxzm49gAE2pO43
AotRHJFByXRC1Mqg61ScLJSU4L4EbxwS9znsSBfmdIBxLX9mS/WLnCHCEOYG2jwP
OJrkXijcpEBW8V3zoBDdFOjNnXf/hf+uMKysM5GTqG1gnLGQCDrL5EWzFjGJyADg
G1OHGwXn+Jsr8wy08kk0CrMB88rWjxzkctixFGBw5XS4X6LG/N1r5i9eqRq1uXER
Dj7PX+g4dmsLywNvhOTvncIf6uzGLR69y8U2M0ZG7eqLMLr4vaCuNVOG8dnTkoeY
OK93KqoSE4EaNR1udq8l8TSewhhSV3/vjQk0RNFf/tlTCZTx0FOby7wKY8Q4PL8q
kDjGqwcwnh6fNCS0jSYTobY6yP3lUdXCj3SlCneya5aOk+DnGRzpcDVtEqKaDED/
mw7lw4SMJQL81eHA5Yjo5cHvwp1NOj1tVbOSP+hRUFJIadVH8KJFVN6HUT36XceC
DiVX4qDK3UI2qID+5TtBn9D+M7XBgFk17+L73jw7p0n+1my8pJd65D8x9lZWPm3q
9rrL9G3VlB+6y86VI3a6Uww2WVaUk+mtORMMN7wJThQMWpSnZ7Ec0YlPNob203bw
FkRmXv8f9x6spsCIZwXv4ZKnqEtBcNo1/xuHXQNjEjPCCurZsG9gXEogEaz63hYW
2gOWJz9klIcuI5EvL6ecErBfsKKsxDD9f9IZUpdptiBcL7QfBBxX/41zW7mlWr/n
C5oHqU+9o5W8bFbhTHxJe3uYwklQT6dNx4WGDGNMBYFkmQZY9TVMGgvWRx+1IhpW
nFa8l37o3sJ09fX19akWB4x+hUBSrxVZ00j4j6OMAssxvlsbgdT0jie5uIcUZWtf
OG1v7LhVZJG06Z2Ot7+KdUE9uu4etm0+wz3QDhtYJE6vj8ZXCGtesT/TGboRFNiH
t3bbJBt76RWKUixkJBPrhMqBqA+1/AsEZcWrMW+fzk1072OSVa2g5pOtjd9Q/iDx
8Hnkpts6T6bnanaFfVRHr747feA8DeRxLSpHKLIbUcdaYzmBAAWZqSWeUHo4yoMd
Qqj9f6S/yaMCegVuzsoetHX/x6bQuMz7KJMPb0ndMfvbgi+vNuK6LtmVpDr5SJIu
HKnBnmMixF64Qnt0IUIURhoze1KXceXAmt3jvDdnISv5xrj4fdbGMfI81Ran5Cc8
3wlGaVwdOHBKmVZ2xpcKaT1pBV2/ynOe8LTbBonke62PM5Z21R7EV0PeSOZoeunC
vBxOVMHllAYcx6Aac6etWFkgntQrb55u6hy8My2mamcZUgBZs5Gl41pLsW1wNJpv
dZ1bQCMxSgEuUNq0NpWxI4iya4/iOlRzvW7haUEXqno0PSpmWBd3SVC0+xV4tSTp
o9jxf7lC0A5RX76WM2qtEsafzOnM07MbsiymRwnVgJXKXm1/PD3fQIbQPbNyZQ4x
nyQe9YJz+rZzCDmtQcUon3x/lfmVYeahAnfoG6A//9yiXAKbew1ji333K63BYDZx
Z5YcM8NFpGqcZhcr/FACkeg/XDrWq4Zf/YUF8VkdD2qybBJjcPeKRJDvtvTPaGBp
x8XVP8pJby/IYPdQHff9/SOg7keHxMlnL4uMhLJUkLMWU3+sqzKMDGT42lDoPMBw
6QO8fzTQGzBFHQ6qaKPv4Ephcq3LRtqh77zjwa65ViBvPgcH2nCUjNu1QqFR6xLV
nfGiIQVXzrlODSjhtquFn0r4EmDoipQphmj5GmoEnOZllYo2fNqxPJVSJcoLMavR
2R3khRMXCvkvI5ClVxAcaxGiZb+r+IBClZ0jEuMRXPPMKVQ35/fmhYdXkUU1GVez
dPLEDZ2wcec1zDqAoVrD0G+ZbR+i4qvSrYxixwFedBbDeTQLUZY4V462lHyMXVZc
XS9yF0cL4arkp21oGDmV4CLFhdJTBSbqAOu6WmtJ67HT8dEJH3cT8r/6Z5Dkpobl
ZzgGlg+EB7nbdMW4stpDzNSTIW2N6yCJ+a6kK0KQVUSCkyovd6KFMl4a8331iU3u
fqZNf/fjq8Oaq2mqd56WIDTj9A4d6cDmBljFQTQxvqznZTyVA9X2HVgZy0+c7pSQ
FXMqOcVARL5kyz6985zUG0/OEYfT0+wgunRG/QuQLajN0gVmxrp/MSw87gBhiLBQ
AYuaa/Y1nqOACP5icMrQBaVULZH7v2F5jFzGMXL2t/tNj3I3GTW6Sj5zXOv3UhDf
Rfh0quxnSTAXuR2k2hq/FPuwIX/xLSFKz9Mri9SsU0YddpTLF3lnz01OHfmgXf90
sjB4iIDHyLm6PX6tFdP4D6+okUWDOF5dz6c9uzwNShtM4YMWKx+a8sSsP4dEHmza
LaZBZgkEAi+WoIyz9j3eiUc83+YDB6yJ3t7Qwh+DpMuD8oLA+hsnl+4xBLOSyPZG
H1bArEJbxX+8p1ToMrr5T5XbdH2y13CJpg1QwDXclBDrkF4o0OIBeUYfC8Bg3pAp
AeDOujzE/6C8ftslny8rb3nueu4XmgOWY7j88el0fEbOHaLqwosF4fGNiIMuE9Tr
TWitq6tNyYckqDqSuOWwhS25NI5jpmYZbMIdhHkwYn3wHuIbqgIyGXpknVFqfPD3
+Hwu1/JejSwWazuWPHpqd5pK9/HOL3x25VAZ1ItzwDcISIMoXiO7H2mvou/da/C+
bQ2qBey5ywWGYcg2LxIqxwnC7g2nQh2ELrSj2lpcd4ISNMGW/IqeZB0SM/+Hm31J
N2s/Xwzg7o4TJ4fVqgvpVo6yYQ1lpOwJ8dVHbmY7nmQOIYzd6YyjU7ou9iJa33k/
7xC6KpHwrX9dcEJJenEhMP/eZc0Eo6OkwXp+Q5cCorhbHf6WVTOaisA+aD3R/iem
el5Khir+ZHbCYuakBc3F875xqBQ2IZlQKEsAcYA53+7d9S/nHCuYnCUeXeVfqxtm
bRTiDnbUoT2aHb77xc1cdlqoOp+m2mZeMKt0UsBuCXS6Ceo6lIEqJ8nW2kuXi8FN
/boGS7YjjaXbTEmpqLRzzR0TJO3LoxDIOG+CQ1l8A3r+fj02CdW7zoLtTDEStiP+
t0xWA75Xu3zMuNOpw8T/ZHCXOYmE3W5X6yGEUa+ZnWG9Gss07rAJ9BWAO7aFkRgT
eo9BAmgDrGMiFRCPLR+sUM++7iZ0JMEBdkviduggZzNNQ4f614WvF6jx+epVnQml
E5bE2W/POz21F50Vr0aQRwqE06HCjatriK0F8fPVyAXxdazhWt/z/tLxcTsFu9cs
YSFg7gg5P/5/MSedmt0Dfu/s6zTqjgMFJESEaNCkA84EmJ6SMnWNH9WeBaBKCfax
9JBQ/4J9KDeip5uqulEMEyMksDodLKLn5Kx04bw/5vKdb4Ew/QPZADuuCyTzWF1C
Gy8wv1GDEnyaAhs0VgkHG/oCG7Xicmg6uS6DzVgYKOjLuf9G74l4FJhqotXDCigb
22Fl8dPljo4yghsiYSxHGRSI3QUxXdgi2ThRUmifR/r/SyEtqficQZOsOp4thxYh
sQvTppQz0LahZGiv6oh0d4F3u6JZ4liKhmzjD+XCAJvApwyANqfZ226277CMdr1V
qQwc8MPTFj5KGzGr52AcfQi5sA5iVa1j9zEOMy3cvOscgDzyR/KGbiCHHdsd/M6X
kp0G4r8H0bhbgkLfi8WcuiGpHAF9gDQ+q/HWdiw9bPc1+2VCUdQ1T8XlwbOl+vZe
o5iSFPCVVYRG1M1Ul4Z1JSPECv6+IzUA9khJumsQ+2nuJxQywqhpmafEyEt6cML8
Exkrp/h5kx0OgTBhMjOk9NOOK1ivg1sPl+pUtJQjHfqt4mgn7YXpZNbNckG5Y4KV
OElISPbQIurt7umLXfO5b4SYEJsviBK9MtgCoz3tfXVrO+rvaHFvcFzGnieCC2We
aFYeiLMBytRvgbFAtiWWTaRO9tVBi5vDjD1mtPoilHYOGcZ3/V1+y/jp08qMBx+f
BzQKOk2aAYYAVFadZ1r+Cfn1H4E6ZtmgiWP7msCnOxwW/16U6KQW0ATL6ACn7pfU
PAr1hpeIGzpZsQZJaoSWQuoxraK7j6MB6uSN+H9OCArkyfkJ+4kyLCTSU0Dzd0ld
GKKyiQdHMS1y4nQ8N5/4S2d6gdXCE6dHvfxD7Zwp6ae+MN38JEoJFF5Yg2WM29i3
T59eh/Dpuop1KxUl+i8Zm8EIu5Vr4xZApImIy5Z2yR1ghRg2Rh4CuzRgtRaqVE7g
rbbDDvG26JtCYs5/5WDuHMmM1eA4ZmbpGrEUgx2Jwe7y01z4tCslXEEdOZgq9o5z
KEM6umatZYgsxLCrSsiH0FP/FWLbgovB0/DYql7PtpXxQl+q1g4k28u1rcPKhpgt
sqRGquknkuda4lIJgFXsb1go7Qxy8hHd/xonw1rKhuN0p+vpbKQSpR0MFoz6kgdw
vDKxMYHm5rEAPZKiRzn/d6yJDcLkeExTgTtbirUeLunPuVGDcxavHFhGPWBHEdsu
2N/8e9EPCV4y4hT96Be+bQm0jgSY/iHl/JDNZ0FaCvd88vd7RwyxB+OCsXkGbNU0
QY84j+lz4JDph/JiOfV8pNb42wf5FrmZaKw/JXODE8De1NmPdcE8drCNh76xZoRB
z9FG4LM703Xg8CBulmdQl4F/Dg49RjCL0G/VIxCzr7D2X2A7fKQPvbDkIaYcpFsi
vts97X0LPH2MfK9hpf2wCBSTpB5TC9ZGrjg187qjHrFjuXxe+Hy1THvJW+1NuRNG
Oz46eF8AMmL/3uxiqf/E2q3wKN1VbVNo2+DZPaU2ZqGyPIFGUYI4HGaXPUFI8XbZ
oYklfhFF3j89Dp4h/y9N/w/xHNGhI98nL9ZeGlKUdXaTEoxR87n296DlNyz0UGgJ
U2pXAhvHrCR75JALiDOOqZppmxuTkzmUkkmdomb33CUy749ztlSPA8FRi1cMY3ut
tSr0bQWSuCA8NP4TqPOJGIV8Z4gql1ZXIRl1/2hgmaVYhaXFFIGHmTodfF9EkwnG
9oBauTLJp9W0i/D2NB6vKP70Vas3KmLPcZ819x6oYxxKjpOLHONEVJT+3RiVIyPY
Fi+gFk1Ie8lDPjD5YJEJu5lstGae2soYR9L4jhkoJBLh+ogIhtXCDecs9Q7JPKHn
Q9cG3zWmcdrqBETTfvRUqn1ASrvsBphP/UI51GMbWbCTIxazNsW/RJ0JuTMv7jI4
xEOGO0YHQjbT71DcZ5Askx/I+ijRge0ZGCAiw9SRIOWXieHgnxcDk1aToTkOpZ0D
txWCCxMphhjejarAfCtoPda2PpvM9fiHI5BAVRu2Fi4RU9aRU2E0UEOmka09ZNjQ
icHV2kMHrNBh9dqg78t6O6uQ4Gz9t1nE8kbWs7QcdTc0UgoAsJPhNw0VH33I9UXK
2/BSS4GmIz2H67mEvmBZu+NuZLDNj1G0wqkdWrw/blcUKh70591HUFaS2tA0YK4k
0YTYTvIBiwCPi0FxwdHJO1s5s0w2zk24VPGpiUIvqI2FFDq8Vky+Mc+AX3wuro/I
gdofleW+m0McInFYkw89oYd5HGUd4Ua/vWRrOK5VMPu/w3Ifm1OtrQ5j/Ygni+i0
r1Fjdw8hZUkWgzXnt9BYTsyo1PT+vYpOd+KyW7cWSO2k7Jmu4uBeI1uBe9RBTkbm
/AHv7yOFgj2ucCGYvxkVLAXAeus6lvb7jcp+3q7D6zcaTeiwoYDDVzrZVvlg2hzD
k78CF8XOv3fBipRC/GD2dhBqPGikmyYKXoup3wyF2woQ6XpYn2vozDsilH6hufZY
GMUCSWm3uCYl/i2/zqjZC3Xn+qZ2oAA0D45SqXrg1AnlDrN42bzuoepbi2syHFgL
9yXoeDEF+bDwtKJ5bYr1qHE7uA/qIQF9JedUJxrwBcY2r+nYMokfYzuqG6RDzJBu
R4RwyRtzt+taBTonO9DzqqQktZJchla2YUa+kRSAnX9HRgw5L0U6o1GOB5fatXYi
Q4L+eb0jkra9eGMXvKI3K441a2KTvFkmNF8lRLhe3XYaxBycfd1FQ6yKEhYedqMP
0eiyJ5jToU5jqmE4k1CuocKkbXUt2Bw5DLVSSTKRLDXkncLJGPb8w7yGKpgT9AS8
TbnsOTZwdPB0sT6oQisXf1H0x1OjTzpuIDOlLSzdrTGhmjQozRp/TqNWohkH+Y0v
MHZheLymJ8JhvliwFQtPXyQjJksNkif11eeZeBwSow336JBAoZymc6lLmyka5iJ1
hhXDCFTc0kuPkwqIKFuzJXdvOlP7cpg6fZC5vObNUm+Y9zYAZptLvZvGBv0h/YrO
BW84JWp0XO9jWKRGnmq8rnTTd3pvbk67RCzVfOHCyKdA6DGc6bsnGSo+SScv3m+N
F6EeumweUBBBjUV7KnhOKbahu+hklFOCru4AWK+00oRLU+DeVYggIHVctFvmcrPT
Lj2JGFsr98njN7ioicwhlfYRersGS0J2eAJdtaJj/vHYQZpW7Y9d+EcDOJMF7Wb2
tpfP++pEuSjDUFLPki3DmX7K0xuPXo4w4jTOniMmxdnjeo03/ySP/aXlnJ+Zgo7Y
a0etN9KIG1ddQeRjRzwLk16jUau/bO6qNMOV6Ms7LdUxEzgUAv7IC0GFemJ0Djru
tomFRJjHL8be8nxmeBm/Jo2z5jkM+hCkCsoOAJ2s/iRD8dbw/Lu5NrDETvQxZIEH
Q6lD+y+giiGyD/KoBwKZPKp8lDNcydDlEvIIInxCJRQreoG5Lg/0JUdCMub68rwF
jwU4/0tllspC9UPeMomzOC9+2a2CJb+mmZ0BXvPI45iDqtTIW2apudDOedDzilcc
NAiYGwBpUzJeNBY/Fgo6eQgfLjCY8GHD750HF5IMUDU+RFW8WlCaR6DSskLpliQI
hQ/A/MRZXIaPD7wwosTSGz+DhpNUXBlGlJx4LLWBLTF1oO5+7VspweEGxxnWGVmQ
b1buPfUP+4aoELQhuTT95vjz8RLiqkHOB5kH5Yp2U0xBJ8WMcX8ZiyqWOJUTgdCn
VH8UPVPzU2KauIOmefZmReYdZpQnDEKRAQg63879mkycmtBFGcgfAuamsxoPjUOs
VajJ3uprr6htGLfHmei9SszBuKsQeLJh24OeKqACNA6yQ9gc32M8KEDI2rVcssUz
Qxhoen2jIfGcK9rH8ZvTP5NIvUdEuoPDPwyQpw6Zrh13+It/MpymjOuI0YPekgra
oweQ5IfOJfW1XlKz2Ao4MTChbXVKBGvdNys2et6x0oX210oPTpOTfcAU3ruh5+aL
OyTzbUPNrm7SHdw99GzoH/ky4xtzmYqVp7p0zbAc4aMf+xqCX7yLW4Gg/HT4F3cP
ungm/csq9XDHsXx3Pi3zEROj0aDRsONRChHxCBNOKfc3OsatP11y1ccIRLB+4Fcx
S4tm5/TtYrBg5MEOMb7crVbN4M1IpBEeBA9kGSb/uH96ipjh5KYBfkb065LX1yWF
7Wvzg07TDq3ONp80lsj4pnuMY+v5NtsUw4/rU0EYjFh1H2lcOWx6uzGKX9pixuGk
4ncd+l5CTtWmaVCe444zWtjJ+kgUzVGxbKgwtUsSrIiTFmKn3t12bY8VCLWt6LPe
aLX0pFaXNpPCbO215zcq2XWRthNVp3qXNVT72ufeJapiAZ/2k+nJKWotRk3aijNv
e15ZgY3MPh90LiCjT9hbkX7fg3K4K8FOtjCd7UIBTiCsm7E+XtW874FowwaVKCDM
SWGYc1vVqW2Vu1i0CPvrZNRHiP1jun3qFTkhv1puzPPcyV44zL8B6+KmAcAdCZI9
sTUl7cyW9edP2JeF610e/k2pyGkj70AQAc/MmpYBsLpea0eF9bGf98xI9dG6bp4y
nOV5z8AOzxuwKOtiWaBcTqVOxOWra0J93S1I0a40dYR4FbYGW+S6putDzHbtyoIx
0dCaZRXfOjykFvAxg3QhzKeZiQdbnKAaCHEQtXXt2vpFq06b91fOwyUFIQEL6iCk
OWswJiG6WEQSnUS14TP4Bl+aqW1yeYYqnkrKIVgQEUJcpIJ5a9uF4uqUOTzG1xW4
QnsUXFTR3mIkSxl704Ghz3qHxd1r8EnwPUovkgmFuf/V57sUVr00vUBdijhNqOw0
l95q2y4qtjKD8hfuiRO6yf6YG0CxNwVoJP5ZJSTiMEW7LLt/mi4o1cOt3lVftVKn
MjvDC+WU/V7gmywgmDVIzwfMKFipdaIjEbgqw4F77inbhBqRKW/X37vox0gXbasq
RtOvS7XPdVAyLVmFWr6LLST7617lDWOSyxMZ/BQdRTx/0zfqatFzyRK8q6QOmB9O
hoYEN83AFI1/cHX+QPoBKjLA0JgLYp8n5wiYk6SL9FzHtAtdyfeFnTpPJAwyEexW
uiUdD7zNPRHGOVJyE4qsjT97MdAjdfHBIqhMMAcZ302xTXyDkx0wo3ApZljDHsIi
cyGwC8Gh/SuU2XmmrkdVUTVB91ZoOvRAPWWHV0+yowDEpIFXQH0HbDGCR+Gnflg6
6xHoyVAgeJStADj0boSMC+BlkF5Xz/PsDAEkVUiVLxFC96OmqDylPtgpWWOua26K
NLGzILt+z8wry+yHz+evIUJZNMKA2aVefY6eh39E33XYvBf5w6Fi0IBVIthochG7
M1culX05lTHkEDu92SJfZQB9OdumDirX9rywbn2BJlYruUNx6uNk7EMF6WRizPI/
dQMrXQXR4oYp2Y3UequmGx8R81+0IjzyPt5jI0n+SoD1Ag3mKX8/TOM/9rFs28m4
WpPH1O+CKzjWAcuoWNi7dp/J6zbn00vZtFXsChONyR3T8rs0qR2wzBEMWBYvTBYc
fpVE1zpjp3jJMgkCAVcq7CnHSTRxnx0WCookUiCVMHgKjraE32YwJUTsxdZobkZJ
Tq7a1e+IBpSFtLvp2Js5NSOKj5a4An5R/2+fkirLmQ63Sw7PFWM+2Iq88HTKCTsN
7GX1vPyLMOoD8ZKOdI9j+isZOgpLEDHVH95IkJqVSideIW/mmWVm9JJs5KzKErxi
fdaKhu1oJ9n4q/XAbc3cmP1+R90k58CW2HVAeAx5mf6kfRwQEDADPjvO6oPHAio3
Y3DJ/Zqc4N6hej3KCpg1aDSSqYrUPAI0Lz3kzI8iUrSHkj5Gq3we27ihcBbvAYkP
iZWv8odQKLp4qPNugizk08yRZGzTGOYiK2fKRUcw1TZuUkiXJCuIPc+jjvoD/BSJ
JTrasYAfB6ipkvfwYvwIGaI8IEWY9KrP+5haIO4O68RomTEHl9Vo5OghQfMDkF85
8MhKHWvIt06rRmfkd0ITW4AFnkmX9CPi/+GXgHzpmdPHBpzbp4OGx3Av1ud9x7xH
Vx2i4U1ycEDYTMgYNNTi2IR3hmrrusNon2fy62XY0tE9l+IBruHuUSUhIWxX+5+f
e8lxx3SMY8el+5F62PCxl/yXuvApoSc/RiinmGxGJsL/2krDzLf4pIVU6bVgKIyg
LlwArX9kXkyJmopeDu1JFHFCD4WYF+XnSkPLYDpMCqj9oQlHxM8YiFpb0WmVtxEr
WOupwHrg+d5kuJz58yteZt1b7fBDhq5vW36lu2DDmimrNl8QL0APpl/O5jMenllP
yZpu7tmnuabtmBB9MkTCXzw5ZWKF8mtMeWKaUhceEnpRRHEPERizKsRrprJcswZr
F29RipBhqU7n0ULfvh9lzUkuVLp8nycN2TFLuakLbGuPvKKBoChjMlsqZvogFEMW
JWRNIjZi76FR2bPqHuk63D6sKaW7q4Vrh85r5CHV6M+Ij0nKBIrScwP/UIwfaa3+
gnFtd0vNTonseW0m2HpI6UW23d+HbNHeBfhVSusB0a4yyKepWAzZfsDVf0T5ThpT
PKcW7lHc86jqW7WlbaKa8hk0JJPpPgDjcN+LMfErpMOzY8BqROAquYQ9xoc988Zg
28G5KZMHU7KzOcO3aw1glrizPm0/3zOJT+Mnv8KZjmVKTS3ZnVk65NqDqPeYOdVy
5exQUieeOutdEM9xmrToDv539mcklWq0upsX0JVqXtLhlnIeCF1CmELgvNyu7CI6
7qlVpHyFhTFx27sC+NYgEfWJomHlQ/Ln7QQKBT4Jdmb4DtZN0Bz/D4txbB5ZNKJC
PYgnyIToyBIhqJZTZebDgIitrLbBx2QbwJjL1XUPYPZDs8Uk4OctfXEMHniHnlMs
o8lBv2d8+XJ6DoNY1WIGhWYUqr8zZwlFXPoTNOJBjD6v5juelHocYz5lTeQRAs2E
TGpwBa5IIYc2ux8o3z+3m+5y3XoKT3naCB5CyXcvAePN3Q3sFN2bNJZYt5+KE3UH
3rCx0TMk08i40AfTWtTZ2xypLBvZ4xb6yA77RbJoeuUcyYgqorbBEhBwRWgz38fT
TbG4y9YiwjcTwx2XB+E0j66QA7EDeanoUKu5fnPTWobqg0UHEXohrIhq299mYBvE
B0JVMMfhaPKSDwU2kYGdFl+TY8NH8PonfPazAeeRI4okueuN4U3c9UBXj0rn7RcS
aAQLOl1ii+XHjfudtB37Y9dIlx2DAAKk6J8GgI6pZbVzhVxQAkAh5t4Ejde6pTxG
P88/EeCzEWNiEIG0rkqqUYq/yW3wjDYgPFDf7+10E0aP8lb1sGg0oDBARhh7Gjhy
mEfy72Y/IHpo51X7Znoh2CMBqtaCLVeZIvTO69E76EBXfrZsnbsVdtUqQ98cFCdj
na+DJZ65+0VKE78zMUplPaDkfoW3FddiNo30B1v7GUn9BRhYBQ6CO/vNt3MMp1h7
JQHNBu1og7c6vYGjG7v+MhGIEyoARWAU1gEms/JWNhhxKSbf5K7e2LTHypqvkPxt
nHWrM9wlQOC5gt8jdJKBBnN+yVt2yi9iWsgsbZBmpwfLt1Oxc0L5WvYQwPLxdKii
u5CEkdEqNJ2CqpUEIZriyOplzCcSGSRITddnrbEIoyp48zV0lJBlkjVILpEXfgEX
o7QqSYK2V1jIrakIK770i45QdhmgO2Gwy7ngokLJkDz6sRw7+dkmRxKWgQI7Eesk
SSLrv3WWzib30vu9DObWcflZjKYOPRK+LAXLTTzg2hgIGaifNvoXlcCpAiDHgq9h
jIoR/z2oPk8+WhSXsCmY13aa5K66cetZd1CSpziD6ftzxigs4rTDr2YuUQ2SUEoV
WiADw1JCsufzMJHdcpOL2KeocatdwE+P2vRu4ki6tci0xlefvudGYOMUxhhAFeao
ARkcOKsYPxIIGhiAl7oH+3mLcP1b8LJq3KZYeSHzN/JCz/CgNWjnLBldXJqTwOUg
19wYpRWLDc7QTgGjLJ5BMdvVMgkzI+/XbckrPnMagnOSnvXBgpnbECsVxpVBI1MM
/NJNRB52HObxlVo6uOlbN9haykTGAR3x2D1Bvz4412pcY5t6501NuOjJMof3gvOW
e3e4WP/Z2Ss9VU5bJON7Y/AwUB/iIWhqHQGOXDLRGaLTv6+WCeGVaaCz2TteylMR
COCk4XtITKn+PRYScCevq8E314OsovohpttrwreICjEKnXZ34ghiNawkJMLg4pfy
3xmuNA84fP8bySpBEP8+41xtgzpu0lX0Jw43sKPwZTPkj9Li1Seu+i77SMYJzFhh
zQqrapStGVWrHphzGGaFnipaPS/i/xa5y8jnakYr1ov9LcCHfgeJgNLsnadHsrlG
eR7UwV85Owxm2kRd2+9Ou/JJVw50kFzAnX1lZMNxvBjA0whgaDfb6bNBOlqGWRQY
MyXSV0X/cYZLGqtLh7swq+s9tGfPxc0WAdbCKkQrvncb4K1sz5UkueGLLal/ZaFM
cU17chcToK55I6iOnQHVB40XKdhx/jsvt9C3TGcfPyqdyVyn+jC35Gk+GcrnFHpZ
u/S7MQMmQOUgDJT3dYKgHV0OvnWEx4oL3RfX6jWrlkB1xD+OVT3chWwNORfUgBJ1
4dbjO6FzqjKZhb9/Yn6Y550lpgKBXW5ph3Rf/W7AsRc0Ubo2AIFqw+nk3L2m/941
2g0++neYQgT9WXWjrKDiPocuInhnPlHfA92J11hvQq07g0Hr4XK/1TokBuCMr6la
eAhl5bVzGuL4MGq9hczkTtiPBtAy6caEeEhfimOXrU3Ctj9VnAjk9KBocWBg2kN3
Pj/r2vs598TlwRMgdyeE8JQ09QAdtYPpEGAlGRluJwO8sac7mMunpF1L3Q0jsYgO
FhcGmFevWlmt49IpzuxRCoBxxcTWmWeQgqJly4fNSr/Hs01vQ008/Qa3CLZkKpSb
0zQDE2AEVbULp7fs0qguHDk68d/74EwdQpJ6oC5LNSa1rBK5ZFMdt4eMagUHcowY
m8YEWKhUkC292HLLz4Bj2pD1KhTh285lE6+EBPyCHlh44VfIWO0sBxmcEq95rETH
Hhzc77fMn6jjRCoc81O3E0A4aTXiPuDWPMm+IL6rBoT9QkfX7PHHD33udO65BW+4
4AGqBZIGdykjnZryjs5k6YPnacmeNDm05nrYf262kQN8SVB33WKHVzL7Cyhv9iYz
hjfwVrQ/Ek5YLWBJYN5zBII2DY1apriYW0AgGgqt8GUGjXM+zaWHbD+TsN1BbSpZ
t2rKuvyEqe7+iQCmWmFUjMwWMGPD8Z8NsWkc0pyFMGXHbccqzmUvSmODP5IbpPf4
1cdkACpPD2EOWwnKpG9Yxb06SSnKKFF166bl5IWKSmARDA4u0YaSxtcvfwQ6q7zE
alLHhWkW76jwdX0pnquOyBi0C0Y3E0d/Fv0+TcsUOjRqZtUIaVO60xkaMjnDO0An
zqzWAoK8ixYhOTZnQ+1Ip+MY9prSpbf+phb3QkBo5mi4JfXdS5d8vXO2FH91f/uN
2oEh/EvsCKq8v4Z8r3FBfSLtN5BDL7zhGpyHuGhneoWTrOI/lxbvEyjrsGmPOsN3
Okv5hel9T7CKTqbphg8HSnGPDg6O5oWxitCGXz2wOup951hfqhuuEdcqMjfJkbpp
rjvuH5ZEf4v8VApbcqIQUkE/SVBcsc58D+MT33nMEQLQlQ0/3aBpL3GA8LKuJ2Jj
a1V+szLy6/pb1A/7ULKVhMmblOYiXmwhFZDcPX8PvfzV4UXwVAY4kk71RAATTWkS
StAElK1VVDq1oO9qDuRQuXKyaTXbw4BNzDoi42DRiKvOE3euy2TMSbxyQdt/Mrpi
Q3MQUwfJGi1is7SdI67mHCDZ5v/onMmuU6fcjbUcXMyiO7lHKqgLSDhniT7resMr
8AkFZ+L+s5iz/2+e9ZBITzrPW6DyFUXTCgxr0CZD1CLcIDSzEsbvSxLHVpZVR7I5
WbxEdI8WZRzZ7eGQJBkofCmT+61TQZkImXGAve8IYHELP0AUaRoffNQ71tE2gKeO
xlfQlwovZcazvLpUJIwCtpNX7dBviPLN/Rs6VCoM2oG0rXsfVFqOnjuYNrcX2/+B
l0RgnN+8VUY5HFa1/PnlN0N/11KS0Euj/oC5SNvZI4ro6zfDcEb5pWXBCZLLKYq9
Wge5laSsNpagb091BztBOBonVAY7FROjMPupC3YRUnwShysYYFfWtASXXKKR9B05
EpBu/AnC2co8Px/dZybYEZPqY7kK7pPLIOCn7kJwQRHDemGwCm7E1Rb/oLMBmS4X
icrGRgRSAKnlSHBypCZpZDVqP/2J889UimCVLXbRJabMnZe1gbqUMP7Cx3QKG+EH
k6puFffXvkxuP4qfkqkVaiF7Vrjv8aufymttXwE9TZdqojHEM/58m49qSL6e7wNM
2H5O69MGMKHP5fHVQVKz/qZUJ51StERf7AD+70UhZWjrfkwpLFgEyyGnPZarBpKj
qhNAkKbXFjZfaVdiew+b2ubTTztPOmOPL3ByHhF565qgrwhUKSXoJPcvajC5U92o
H1n7BGwOFxV8lEC9TSi3Rsurx4wZhIgPkRS9wb/+16rUqfKfGEseDZ8b3vAQSEw9
iXumZGAqggBioynVngRsHgOwupo78l4yPbf0ie7qf3zwYIIme5DaxKbeZUTWwWCi
RELV+UStk4s+CP/99XGFiBmVKo9wHCnbYHol3AM+Ac0XbO8nMhepBAjFAhlChuRM
+AGS5ttpo1K/ADIFdlQDHBr58tPo6oUMbvoxBicuABITsKgtt2n7+NcYtWinKMWF
QhC2QlDqTQFmfsZ0XAWjUYR7hPKLQQfxoB3SBQPj0rKZi3b5vv3MfkpZnmnjxo5m
KXCM5kK6QNKRHHY0OrAZi4+E5CfDhJa6plIWaE8O1Blly/GAIC9dcHyCO7NcH4Da
DvVcuX0vqOqbE1MkngsF3TGPLeQrVVY6VFJxINvS67KrDLflEt7c14HJAL8SucYT
Cpp5YbYrNFYTkf9+ZeweMeWKP2U0Nw+XmI6Ga/7oNxo3RPCNxiLRqFcupFR6WVXs
KkZ7FNevDXdH5NPZ5wf1T//R7+N7LR+8/3Obf/cjp5IBZpkYG1e8PF/yIiJV4Vac
ncqLBoeesJxYWocomkXv/+dZSoMHJlyuyMmd/LhJf9i0HjoGXcmKQLOizGQDTE7n
e+A0cggmeuUCjlsY3ahs7kSzGLF+o5qZZs6o/wOI+Pza6k67pVZLh+e5fgDelnnU
Gga2gtMGm8DXQJHCQOC0nYoFEUiIm5qeDSgwNer0nO+rCfOBKYAqPfAGkqlUFt7L
LcL4ZY/CFkB/hT71o7vQadSMg9XK40H68sQdSUwbgmso6xkznCmUkxW9WO2HjlUx
5/+YBzAYFm+Qdw3ZS1OIEY25OzuedvOxd2rfPOYtAF9soN6T+JmpbJpQinRDPGzK
KmLRDetFyaJvbqqgLFvJOg5oChC1WQ98s0oITQ04IQ9K0punKsZM4Yx1eiyLxEAL
eIjl+2oNieK3Nhsik6YV0nhpesw09y92bAIWI+d9eLUmzjEWW0O07Yr4JIm1H85I
njqEzvFezwF/qec0tylsM2I/WYR0e8yc4Lx6UZPRMUJZOLtaJR9VhosGPFTtExuV
59Irbl5DgZgMXpVd7ZKech5MmfuvmQHe2tPeM1ISWXl5snsvPHFqOv7QUBZ42F3F
4GB8rA5gZIJKs3U7Yzjii5HKG2dEMQQ5JRsvP04RKN4GZTDZtCI7CFs+EFIqvPxL
EG3SgQF9dhxdj/QAdzG/dTQzcU48BNxyjD/mKT1iCUwY6Xn6L2OIDTsosu5eeLrK
m7spzma1AYKrTpT9wgkQMNCTGxolHJIBdt2oLejuQgK5Bx/vRJti1L0xn24OFcsd
hatFtqIdrZddDYRcvDlmm9sneqZzkAVrtztr1K23SXTqCEbvntzsM72VXcNqo3CQ
38RBBNGQsW17PJBDMBdQr2GPbE4YaSQ0sbB5GhpbYl3gA7pPo5HtDrtGMWFzlQ+M
YCZleKIuTcj0LQQ5NffzHOkO3azhK5NBUsW55IY6hMFm+iJApN6xMki1dfjJFDBt
OJyIL9T/v1WgBtMfZnZSZN3z8qnaO0SqN7kVj2FR4Jl1YHGZKUbT5q3pJccOXnuy
pu7xlL9j/FTttRzsQTWcxIw9eSxcPKfjEEW8Uq9Esjf7jGdvClt3v7z098zToYGs
LQlvUXTtrcuoCjqG4DaDwIdYt6dgNM0qwmZnIOeI/lQNQ32qNA0zmFnfA3e+aXh6
kF6J2YdmJ39jf9raNmBugG7iM9eXFLtXzm4HpDCNwnrcxxxkXeURt7ZN6cIQYud8
44lwXGfE5qUNkbSr6QnIF/9Q+TZOAdmzIjBiE9Ob3Dw5crZEUfGDMzuqm+6tNHGL
JJdeckT8CJ6f1gDVAesC5UlCW+ZJndqvMu7RpyCMpGsqoVDHEHTSDDiH5j8LNpCq
PbG/py99RCuQs02V7dlVayKH1Ion4biqFqpDQyL1XnPDsOkOKGfojAf1sqbLGYF+
IDmw3JruGSG2jQayf245ukX685N2+LBWWb6ZOQJX7mVSFpO6mU1ST6C9xjyv/+s+
Xaj16nOBr2cs42JFTiD54NMfuon1L5kdl4ZBmx0QA0cNpf8RHAskbYbfGnpgUIDK
f2XlboSuyuBZZNU+eqqhhsImkOqEIEyaDvKFRHU/XlzDL4quiLEYFaMJFGeBfYvv
2sTGht7QgN5GO9kYxSJeFqLD0VWvFDVQDlPlGujb60+ImXHNlAOLZOnqqL9B4C0g
zSG+xrkxHz3Q8G6fLWoydtY6JBPErT15EYclyc+dWHR/ZbQ3k/OtnPo1aZywVnJ7
RzdT3jCZbgnpDmlIC3ZbeZP/5GBM7cactSlTICHUdKJJP9DDmXpn6siEiYkQ1aI7
zkwBGnN/qim9cme1gIy4yRc4Kpq1kEtgsOmqWeNmRZaVR8qKIYrjxJqAANWfO+Y6
rbsh93kEC5QGaR9jJ8h7W2cFCUeyP3QgUftLqRiNOu0deVSxGoha0OkDKlmj4APa
48eVU3pR5OktJUmTeLiucMsqJyS6Xm8amvfaql8KfH0mLH5UgD0SCjntFm/2A0Ek
PGufRyJbtfPumi5CVTForWBbtQIHCgErEHmzn+d9CpohxivZfp36PgcwXqwcafIW
a7w76LHdwInqf0qGv9/BYTFRCSyieRXN/AojbjT1gCGNW/PZeg4ls1+HarFAeCQ7
prVR8J8mqM6Or9IWn8mK62xZ4tNbyvqBlMpFKWRwNCRUtest4EYp+pV44vXq3d9a
RlsCREgo9rIYwzGHYQzcNzEuogXW4GG20oMPKpjXURDKHQq6Edfoja+1pn1oiyDz
xlBY2NFmzGE3FivWZzFd57TXJEd9+gYFwhpI4Ly8+UZqHVh0yvSQexG3UhJqcg2p
lkXQ9f8XTRBAeY+xecQPcEBiGSWjZB03RoGkPgbljHwEkiNpET72I1drmyCSD3ol
cB8XdFSK/QXg6ccH2JRN5R7w+2MBSNSwgBR1dZNtjFq4RqwD9sVPrMrSCmeoxfGd
ZhZvGkxByTMg9i4/sSk81nSof1crt7+6Dk93EnFZ+NnrQ4WqI1+BAwVlBX0p0OTJ
x351UyQ2TK6pGeyk0WRbx3w+Bt+gWyc0CAQXhA9oKk2hbeSvZExTjHF7lKjIp12y
9qZNGExO0dpQqQ162ZI54v9Rc9IFxXxhk8U6SJPv+MhfElTgx7Gcafh54ibjqf+R
xOxDL3WWdpaRAwDXH7WRxfr0YwakiIiH0uM5qgWFgNgtJkD2rlS3YLFK44FgFC5C
k9vKqp9lCOd4cozCqfBtZA1NTPyQC8qSerpWVkH+/XAlBB0r6oh7YB7hncZfaEb6
zS4ChulSzyCq/UBgNiZ9zlkSfjHxsd7R0jpZebKPoW+Dhin9/RoWs1eURUA2pLOX
Kqe0YQLV9iE0N2KZ4OQj4zYgpl4kY0cGFX9qby0wY7wfOLQOgExReoFsYw9MPu/A
4QbYNwidrC67jHXfc3ki6GixW5Xamucn1vOYOep8xbqY70znc2Ow5jN7SDhq3ZSA
RDQPfuJsQam1StfijQQWjY186hVvbyZYjJN8jpHPnTSXC1bIzLMIoW3T5H8LdFI7
Zp07bNhDxFAUJHQ4Ra+r1kamsfWQnkbUPZGRF+aFPhnV6/rmAJQHtBh4YqA+Ed0J
XFygJy/mRt5hYoPImnoQ348OFC1ebnFK2ZgQRULTReceL8XkouNRx7O8GkDJTF87
aKSSod/ueE5M9y93a1VOi7L6Eh4qUjOwIVFFnrscoa0dS7svWW98eXTGMNjFYI8/
bgrB5QY7VK49kiU7b8OCbefb8J4h0/gAGP2o9QXrPSgkeV/uHRgnwOPMxmxSh+Vb
SWJoVPbv/QCojdq1pS0WzbOZ2hTXur0Hl2jZcm65BAjg1/q/Oj5p1U/lgfECrDFU
SpKygIpEF8RzJVOh740QkHLtplGnKZzTbHDKO614fAnMa4e1TGkPJEFeD7W8NlaS
+JSfqeKk53i4kZKvo4otsznVL7n74b8eUovGgOPyQGJlq9olRkcAG9og1454RQ5h
mJ2Dew7CDZF3QmlQKUkl/OXT4DwEDhdpQ1y4UlIDuYBwjeqTW/DC12CT0hFHvW+E
NDRzmDKfeLz8XOMs/vU2PvuEW5OSmGu2c2taNpEvhtaCePCxUI0XOm0Z1EA7BEZ/
rzXA7xDIzboJOt5u45wjMVoSvquC9jZOt2GdWB63XABKiG1TZkpGGDQR8iQKBdFn
jEhJtzFptGceKY4wwpb1C96WfxUGXHZs8ffLOzcpti4RCQbtXYDxClRqeG/oGqgN
0hX2L2HDijyIM3mJZYA8TUmGtKxtUtcihEVJW/b0W0Z3hDcNGA67upkOXCqPv2V5
piMVtwDPUdSog5V4eViWQ5Ee7QvSO69S3X26hmjOLogA2rsSCTfxe+waA64ku8D1
aSF11w+Wo2GXfSKKQh2EcEes7VF5eTedNRZMQX5pcpn3D8RZ7dNxJHpAEuUm7e5t
6TyAbUs7lC/lVzugO6wsnK8dnLE4E/aIjSa8VL96Hx9Kh8DlYT/RcyWmHpjigT/g
22sB61o1rUAZ7x123PfnoZwDdow8C06uRrcr6jRPCKqThCBUcRWMaM+hK4uzcUvx
4eZCAVWnyPEAmdbTcl7Fo0Bk52HVWJdvU4kpjOqG/SeEVosd3Lo5wrwJPXBVhljn
GX1bNDxkRGlFCSboAVr/PNhJoPu/41j0aPzF8Gvhz5dfKE4qrqyF+ts6Yr6GILTX
72k0rYG85o7gt0xF/cxuaJM7l/D2pEEucfnYRJkxnHx0GVZMETzgcTzpMHKekBTF
xGOpKMQOgRsdYhZjHP8I4Zu3KeRXSW2OOVC46FGTji2p00riRmTW8pp6vRbEXNQZ
d98xk0WSjnVw7zCmD1kQiBdzoIWI1nrVaiaCUrRdZiA9SActJ68EIcXMuUTArZs1
UMm72QufMDUpHlg5fiACAwQidJSpHhl/GGFIYz+XPk6SpqotqcbtYb577CJKyTO+
AiEjoq3T+e/kV52F/iHXA5dqLNimSciWuGea89O4V1BFQXcmjWvYswIytEnzX9Ux
HBaBgF7YFNhp2kovHsMEQr3iaOdqMoxRiDPGKqiOIJR8K0u2gPbTJFfWGKKkGL+q
rwLzbVHcPF+5W5oFZWNcLqNu2D384B/yUn7jvlwD9GPktSxbRE24KmoNvKcJTOO3
6qkXIauBcNIVuRfDaitt07ok7H3oToWytrO5kUl9/sxpyqndzbX0H4UPhuT+XHVR
K79Pt7naW8NJdCze7jBl/awsg0djKzq6GEuIeEWF08rDCWhFkN/V6wSt3f3oml4t
rLlGBvgBQhicCtyGqTh9H3p7CO5d2CYcgB/hhQ5+XW72ZCnolbPVNt4gdkVFTs0d
7PeZQA9HFNixJbDl42mtgPlnN7rgUPCAFHvyneW5QLLX94qb5gOH6v8W/3XP9wWV
XKiFxgXvCx57uBHZ3VwfqGDRLswP22Gc5opXN/VIs/cZye637J/ZPLqk+IsFb3qk
6mEC6Y9Zb5oJP9hcjBqjiOnnmsA6JpnIeCBVNetvnoqIJzmKClDfsmaR08cUui6M
XbMQ5FxSieNLIFDXfdyw8xoHyMYcFp0dtCn35vFRqbU/vRWJ9LEq+pkqkGSF/ud1
rrZtFth97r6GCGKC3aTPdV2HBhgIYR8CEzUvau9rUi5cOH3ZdWrphE5SMClmzgW/
bCi2IZVcXiLxC2w5ApWrygZbj6JGOM3wzg+gzyy1D0aO7COb/8jHHdqKf2YlFNgV
zcVAz+vYpstMFSP6VfCHgGysbmq49YC8FWReUppPnkZd8Jd4uGVCmuvtbW1CbHth
hqIHKjzgyIjOgkut3KH18u2Q/5WAZPOg9SptOxR12UU7DsgmYHnI4J2t6yAv2acX
dTO2vrcXGxEi0C02WCvtn9mfOAmOuhBAJWW6aaI+vLAZuxASvGwBV/L3E2foLLh7
lG911X1rcRs+Ew3KyuKuKhIOpu9KFT7LxEf+aOX9doUOZ8NEc77zcCJYsVgDGOyD
XU7OmK1C7ndIRgPkL3InjjDHwl5+VY57aki21RgdC9c5QQgog03nWLjjyXKb8WAU
3ApVmmL7Dqu+LF0JzHjrPOrW7iyWjzDs6wqzieNz3WIVJ7cpGEbQuowZjwS/mn1P
8CPmlnFELHyjSW2Pc/sOtxAF9XqS++c/vxSz3/b5kGXGZUKv0KP9vGvLluhXS5LW
vDOigzoA3halZntNcWfUfSjJnPkoMMN7PHzT25i7lQw8kcmzTTt9YNt9oT2SUZW/
jlM/V73iLPeuzsaUMLYVUYHD/DuWEDDTtSn0Ezz+MG/9h34cdQT6fFxj3uYlbUF9
sQjXF96PdvTFQNoVKFWMTJxm9m/DrC8IIe0uvkKPXZ2LJxvElRRfGl9pnVR0o5AJ
279o3AFznq6ZjwjmR+AFT7/Z+9e4K3Q9XMEvyCW0I2/EwTze8pQ0QtIcnNkYfNwf
LIHUCQTbAhBkpZLtdDQgTH9g2oDjUxlM2HuE2zqmTFtpxBJFNvhaQf0CV/JEoFYA
qD5RtYHwbxjvD5sdSJM069tBMw+bOKp4kCZ0OspGQcLXJrRTN7NsVn/ZR61EAo5Q
METIM9eI/ObOwM4zSpLKRwGEyWgmV46IjtaLOl6l32ujnnE4kwt3+PDuaCmkfYeB
bVpXj0M8oAP0Lj8XU7jeprBVPEuKksSTYh7fjEavW6k8QwaIFJnurbuhkdT1Pb4A
ZI1eePpjpIs7e3QANntk3r28HO8cml28iBbj3nK7bmLLtM08oAqSxok7cbHmjmE7
0a+XRAiIivTxeoZpYykrCDAC3B0bgCdFzXxr0ytC/6TS2LLeRoL/rmTY7qHu+H2f
hKqDIR/Z3REgirbZMmj8IcjPE+KrfHovWPxm0WZO0Unr1/ADC8abUUMUWNNaH1i2
GcrimSR1D7gZoq8rZuHUX4RPpbynfIgLWJtOx1NkATP+yi3tT3tpKdtj2u+2sbF1
Tv+3XcnaiBzpCoaxAw2vzvllDEC2WEGBztwo8KfO4K9AJs87vRRp17I75xlByaQZ
4j0kXodpDSgckbgPfy8K8RIsx0gSATYDe/fW88ofgXyXhf1BdchB5bIbRgl4Q+w3
rVT6Q8kTfFtJCCBxiDl8jQ+2nQftqvs0H3F+jWrh9PCSDbkatq7hyjeOCALMQX6J
wnto63fAkLT/9DkqR3Fsau6vsUvegHndThKGcCJNEXY3eSqj4s4OWusB9dOUUWwv
jDCj9X7hXtHLj6SdEp9SPqG40dsgipJBgClSvCh05mayyk1m5PcwPRxEZ4LkG8sR
zFkzij1C5QhE7FI37ZF81g5EuuE0EZtjtI259l4i/9BfUq9LQrpAxcFyZd5gLDwY
E5C099/8Ld3hlpIWLjFuw34grpZY3E7N4oPpuN4qEPSSrxl7BDURHWJPxGgtUY9u
zKlC8MHajcobMKlXhaOrZcFiTMWiYw11QOju4+CilsD9XlcYhAAvZtjmcN1xy+1p
EUUyNsadu6nOBUdd3RE4DJUP5tkV1Q7gIYI6H1+8ivdJffrqCLV9PRwswnq3VC+n
pxDwCeSvTQ0wB2+r4+8qWa1MuqyiiEpLnug8noiIktr2JGY9NZ37ayewhHrXoBY2
mg3rmmyqs4QCylg0vuJ32zTt9pxpEcTfHdf9PpDOIliTevR61AnvqJJqmGDVhH8a
+QN9vhM8zc9919gY9R0a9MeV58x3Jm9eDsqf1eSBGHxrEQDWJ8sezeZssCTn6Ad9
ltVhwvdCL6n37tbJ1u5nehdc2mpnAmK/eqoiAa9iXAdiMYJSPfpdJu9Ztf4ic5R8
rR8rnbMTstnTEfkvERoyh39Gor9Cd+JfRjecSZP5Z89NUbYp7MEEOE0aftEv7IZb
Ls4ihc6V97qFzMSP6or97ExJQwEHssg0vYE3o/+/vPAsb6alQgZIW1cwdofinOuE
93IcE9OBi0nT7a/rqNTAs20HtqTMjKuLjyZp0Js8tsIZ16z8XeAdwpSqYYP71fRc
qu12pEi/pT/X97f3YcPBoOL1oSVJiajlgZX5wF3SffDank9MymISifQwJtvSI/4x
48JzmBLLKPCuJELPBVKzBOxKUINoDEJ1o1zIpFOLS/1Paxy/CJGsssU3WDVi0oB7
T+dZbxZEGZbfRiwgJMKYTj0LI4viAqAZPhw/RKR8k3fGs886MPWmbxbJEc+opn0C
3t91FxWCOJJnhC4EPkFb90FAA7+pLQJbxW2NmVKP7yk1atBwCzQJnekedmYmjvYX
mwCLIeqJr5ZddOe13ZfWmMgnpAcnEKqZlai5QuNzwUv0FtiEE+yZ5GEC3B23+NBD
Dkp0kBE06i6ejaOcHJzzFuMkBnxfq6uLdHg30tnnm+MbMgJBDG3kpfwpXiQ+51f4
AXZxt2t8sLOlNR4rQM8SfEQRGvBz5ZWRP2OdmmGi0qORNDZ0C6ODsSBZoBu3jg51
ZV+LDmJ6XT3BlHHmEdBvRUcbDk/yvD+JkHWOLCtCHbbzlcQB1IGeGuxPGUqRM8kE
ntF56bRmMwHvQ7yYXgZkNm/4Zc6KfdB02t/upz98ixKTGDIKHxJIHzRxtwttxLjU
RMTLDo7WKL0drnOlmV/dVDBwqzEGCTKAuBJaRvzGEQ2PJHJCLkG1XhTj+UVx2kok
Mbl5XegPCsvef8Hs24CtRtPPtwbCmA2kYJEFU3mQMLVWX8dt+qeXWDIzpcRnTk0+
RH/rSRUHeB7joCduk4krLNuYTqf+6k4ETZvzuA/l9gjNSADh8yqqOvfZeOuOxc1G
zlJulrhet/UOp5yAPw0SskOZHMCtTbaRBeIYpghjQwX4aliPBq5WNv6lKuTsPJPV
7uPfvO7SfW5RqYUPx07fzDAs4bQDmnXu8WwNRsXgbTXVfC1mxharAkPACU3YvNfE
jXWRRSdZJnykL0qCA5Xtt0sgRJ/QBcKj51V00PwQk/16FwWNtYz5CD7Kzko9LhxJ
IhqONuMWJhRzEIFNyV+0hT7MPYLL2bJWMI9yPRUDBpuhxWKenz8wPOR/8mwLICFm
2cZA6Nz1Lgf2yXdOc/39CGIXHUATQtDSKFL20vKm5WNWo5QYHn5EHf9clkfIU+zs
8B5W9M57DYhNSEoJuSUJQwvmUT57AvMi8Hd8L4IsN59Mudv0AW2jp2KhDPt25FUC
MlOV0LuiDRa7qFQF97B9qdUNezUCQbTq33l7qXrl4Yq15Vp1b4fJwA9DRXhal/TB
BYTOVLMtfnlzc7/kkAFaW72WZ2cMEcUnef4wzpLMXncpnek7aLwvO7ebSyQG/qhN
JpZ2h54/Kt4rhOmy95tZDlcLubvzDd8aKT+6GDvlKL8vQduh8aeAvGkR+aG+D+zj
hNcBo1dfNbaA6AiV337m/fCJMfJbRz6+es4T6LeLRCLt6sBwQ9VRO07xeNbadmf8
2JG4qGvKGkG6NXqVcQtaTy0hexiHV+mgCgexB+1TpiP76XcbgsbQuTvbcxkt9H51
V8EtLqs9rKtvi4GqrXY7+CRILIux2ogpvwieyTGsa/++r2TUaQGK9MFMs93Nkm0N
UyfXSagZoCP6/b7okpz1jhyooOZDShWRCU8qwVCMGt54nOCPXyUiLb29NDkGvzjj
f4Of3JfApHhV+/1me5CTgdlVbrPMCjXxId8dKy+qcDCDYECtbHIBTJlMQCjFlKZ0
CVgs4OsnNGtj2nZd1CDgxqSeVnG2Kq3fGvKPnNcExPUOwaP4+3N75my3XwnRg5HG
yu+kZ1DUPL17LxCrUn54RsWAq7TiFvD5QpGSy1rwvW3RacIjK4XJoak0SI7pUuTG
h9k06Cgd2ju6EdRLwIeLDnachBDbB0vbm347Oto7zDlANKnQQ978dej099MkmdqZ
tN4lYXQy2imkulqVLPvzjxPgH6RtxEhH/mcQv0rjmRmN1qF+d8Z92rHcteN+WcNY
O2BRSvbumZNDju7gMD3ilVo8xDpdUORWZQivbJRdZD6UOGJ1WEEISIIttgDUi6+M
G8FyPYGlr8I+l8zOvUuOw57tKoSStJX8e+aiYbujmrNjKvWVyr9rQ1yUR1/yJxfT
cUUOLKYAUhydGV8iG5iACH7SvP8j0RCj2XQldOC6kpGNWXKis3k1VkCFyhuj7KA6
FJsZrjNq87FJ7IOq0iSbVABQgpZVIUTKYlJZ4/AknsK1OK0Isg5Vo93MhLeCQuLJ
ztEEADohyqzavGkYRbDN22ieVtXxkjNNHG5u7Kwi4Hsn1g6FdUenOpUjDdwnN2Vc
Bzq5peoSlH0nOJEr7ZwDos7Qgfbq71plnl7Obe0wHhzxaC0Z2eKQByCJ2sCLVmgC
VvMqYSpkhOGDkinaXNH0SjepuYXYdiTH1u5uwC2E7IdNQdDImXp0vlB5BKgSE7qO
maeMU0wVLJi5hZx6bUEKt57MjS19Yiu1IUAxMEaOm0oG3V0oq13LJ+FYjVwNdkqq
GJKv0Xqz9tr1UGSLvbyT8JAunetX2NoUumQ6yw48znv3T5/YjLrXc8fL9t7VwFIa
FxvorM02PwcuANfPAzf+G2N48AEJA9Qph0pPo7nTImJc6VFLhZj0eThyj42ktR4R
0kvwD9qnZo40/YSRlDUeuSBWYec9rSLMoYxKeCAegWE0tE5FLRczJ84F/kT5JVWK
K2CTo1gK0aFAezYXSOEKe5U7dJ/cBaqnCPZpF1yqwKmtWReEbh4If1ho/IBJro5l
ZIti0PFrB+/t+TKNm0WDCiXx9rGljFqsnS8Vw/kWVYiqAeQu4TtP/PIaZQmWl+eG
+Cs1pj5lUfS7nchSEsrDReTJ0/j6Zasr/BCXghfvByU6SfXL9R4UGEch1i4KyQwQ
LQB2AU/oWUbyfzKbORE0a/EBb2uXBBmj/h82HscKIsHDYCg5Jt5613Lubrj66wPm
+v112MlxREeuu8ydJgUL5tn2k7uZErevvC31EajE9lsA7TsAcZ6XtaQ+RaypOMsO
hME9UerzDiuwRUAdiXRyG69lG9mxb4wA+b3sEBGuSaENFtdhvu3Ge9hgnBleMo/T
nG/vzScgI5pnGw7pDaNdYTbn2svS9523v84j16VIAyJgPKDRvQxkiIhagKxHRv2d
rgz/mQ+WqmlAWTjxq5axssqY2ecV3kWBFzRXEfe2UmqiJ3NNHYRdu1j4zOrjbtxN
qxaYDtZA7tsP+15tEhG+tt60qcnxfdepb46FvMumxMBbB1vDgaj1Cu8XwIKdsyep
WjtrueCIKc4RF/963ydM2WCkWof9WoYZRfK7utCC7LJAz0YxwnmI6nefV4RZalE0
6Z8dLqMHakCfJ2iiLg1nMunLwCZ3PMugGh+JdwlyeRbOQ2Uhkk1cQG6UryJ7WVbo
dnLb/R6h+uecK71odu16gU7jkSp95HZ2dbtweFybFlNGWXPhRhTDu2QIPfPgo1Rq
HOnu0gB2FeVJpZv5p6qyXRMlDCI/o5Ey2Ug6CMowhV/wwD1XbOuQzeLz6ZIFiKoP
VVULP6LguYv0UDUdZiusNNoa9tSwaVMpC+l0gEmyxhCpxcTqkNLQQirla57EY0l6
6ZxvoWIfz21rIBX7sx5GkpNza7t7d4oMQqana1HGMruooUHzB2RcjhE9tFcHkl9r
rGX7IuD3Wde1MEdzFEWTgg3fBKkMDePDr/DIJ4ww4mD7i3KsQzQD/zThIFah9rpW
pfjpSr3UEmECPP48nW03W38MxCeSGHhZVE1zfap7m9wYsHnSzH2UVnDR6xbLSfKd
4A5KMVMiZglaKPlqDjYm0Q10ZATiC2isYSL4L+TzvJotanE1kleonp+GA/M2FHex
rpLqK+AqOXX9P33LQVJslAHQ6NPqOzf2ghqbBX0KVhNOZE3Fk8N5pyetlOZgsK1m
tDh6mixRqKEUvZDXjsL3QWSRvWYuVxeLq+MNEw3+qBQYwvi+82CEAe8Lcac+Mn0B
nucDRMPEUzJYoILF62IVRduS3rPg5SYSdtye5JOiy0YsgP9i1f0oJkJ3cM1/QwJv
NGHIpbbCvd/wR5u1xshh7NNCrJ5uDXUfiPrKa1gFUhjWs5R231wAUO/crvsqXwgI
VwNDLSBuUw1aSOdic6YRlqssFiRGkmyOMSgqWe6mpFsof/tnbZ57OYivgVuuwbzE
q/FywWNPVpORY+tg1R+x42UzyxfYkibycD0K58P0YJSFfl/uuWkNXe+26numGwsm
hkk04gBp5K2DwUQU7LNN3GpRhvIii8QObITXQdlvIbb2vM76CQUz9iA3n47B0yU2
2AUtmWpOmSF4won6e50sv7/y3VHtKCtOi/3Kz9/A2c2V4Jr/vbGzdiysy7FMH6Be
y6oebEN5sm6bAUOxk1oooiSh+f9hEkder07SZHAg7kVNT4h3JdNC7hlZ7edTKa7y
NiiPvPEE0nar19eqhABCs2fb0TTsRHO8C6RZGRPcNzTdiK8rkbFchFtnjl/+IFo9
qFXvy9rkYXfgX5bLUIxtgoKyr6NsvKIQa0KBcO2Er/ZiHfJf9pRB5yJdZ1FqeOEh
VMRcaEzgvEiZ8yGLNiDM8gupAiMEtBnCYnhIwcnkjyki0YbZv81LepB+cPwrqdXI
XAWYWSgqIYMLZ5/HqPyX/8arDEwGLlR6zX2k+FE9We+NkSNbXK6fL78GsQHx3/eW
FQnohEHCY/a+bKfbB8CMOpumXUNiaFNV0gyLv2H4RlzFYpLjevJPmS5m30TcVeUI
8RclxpL+HIGt45tRP97wZxa1nqZuvB+ntDxlOvJ9+5/5/o9groPT8j2SUShC5JxW
xqOA3VVTCkUABSMgINoydlsM4bixKwzllipQMn3o8mfIIQjHvldfrFFqjVa+3x4S
1nOdtfy0SalVuRpMnxJ6DKiPMgLcgUURCKmGsL7A3PmkzRnnxEuDmzjArdmZksZt
5R/Gi7g0jhDAY+uUZ/a3hGAh0c2OzZDe7Tn4UDzkGP88pnZbrtcbj/tOlSwYDa+3
ISN8kzCflBbVTaMV2eJrKxnOn2Mnk+CQ6TB/yPy9JSbAUSuqQx7GInCYUEnYbCh1
9WHdRNdiqH9mUHzRCI/yCBi6Fa1BP7k+rif165TxiKUBu4Ym9Ge6ANglXun592JA
1LjEzGSUFMvgEiieFzgC+6qX1GIdK4gLaCVrOt+Yet8lDEk4RO04XpwuqjQnox/5
Uw+PZbaTHFxgjWT6oic8J23Jg40jCdjI5fAhoaIy22vldrHqyNvy0yBIDlXe5RnH
OzM51oveuVdxYUk9ubwHuZzIWsibYUpeyVWdzHYp14CsMhss0SRQq08Az2BzzgYK
LugTQ5/CuIaVvTsHonUyuYxMlht8s6I0ejVgBp6ccBvKoD7pKKIKRHVJr5dLkk0c
aWzD4+SLQ6AEOeV07FRfvOh8D1Li5+7pOFA2etNZ6ZmcvBK1eTsA+i7YasYkmuCk
CS0vV4fL9K0ZpF6KJZHnto+JIXBOwC7GTk94qnOsa7PDj9xIHeNeQdrwd1kWbwYZ
gf+rKcC79kX/dYWIcTmdzUwdeBOi2wh01Wq6NwywzmW6ORJh1ZcVdOYFpnZbqTM1
/rjfXk74wruKDu4lJ1gp5Hyu76uHdpmCHrDlh15UwFuX8nq9YWbVhdCKZCW9kdy7
zBAyH3T5VB5vPvXjP/bYZHi8ZDutChSHrQomf/wcivL6atTCnd+YN07u4YZWTSTn
4cGN5rVy1e4rl1X/ja5CE8q14sVIByVvNcuLU6W0s3veHVPhxWGJHTu6w6HCo/Y9
G5K1CFDkIQU+a0Y4E4JC2OpaJ/rntnx0cgLpa8GbX3ap6i5pGAtBb/HgJwlWz9o/
f0RVDL6Nc1RJt0A12HRSsufjC4XPZ4Pp4SlpTsiZkwq/eSJUTAOFMbeG6RWcR7hX
uCirpTtEZ7CN7YMN4AbQSdib1eiU+UN/eoOW9CrAJ1Gf0Ng0tfepXuHQ4E7rhrf0
YALZd8b8R8Xx/rItYnIoc4W08VXir5S0J4cIdfxlorQBvP9N+a3dbqndB6KoSbju
QYSSaoOtHMrlKT28rz0kB++NNNpYWK/kBsOU3WStZsbSAo2OEGfep0lacYJGvbVT
lM+RTbA7C3Q/UEebP34i4C5fz2jgBpOVic96VGmN/kkJlsZqkCN9JiTy0Ft4UtBM
6631vlwZaPr6CxE4SAlJxCUX2t73RP9/GUR1RGluhd27FRtKZj7aHV/Mq9Tb/8Xo
YUkVpEYBc688OrT7zVnM8laPWM1N6F1fTd1bpFqc2Pe8cFv1IH/KLojD0/EMbiix
jXKsMP/gMQRGYQGrdzZanTXAzUs1oWgEJ5b5g4eoqvzZVAHRkC+L+Iz/VGArBmrC
F1lnccWyqGozCXx5QFY+JagEMsSY5UG0elp9HBNSnG1Hqh4xSodrQDkq53uCPf1R
ZJLb2bzYhjitUlhtzPeYD4lNYnxR01ik77hWPdWJNIaRp5UvM1vbIBoU/GSMEHAT
1Ft+CmsgXxJAmcJuRgLhGQDm1iSBESnqenx5o2eT196JYRwIGOy4Dx8sndeJe8Kj
3VqKBdeQ56nN2B+LB/y1dfBiiibIG2shOLKsQgra5g+5VP3gWhbORRf13+fpXoGZ
bZaS9w9XbI2RYC0dgcIzwlvSnOAoJs65WiceHbWMYKjdoa3j1sBjGO3yQ7vw+oDC
yx+kXSoVZDH34DXJId9Gg4tIgbx3rpTbu8K/q9EK3QaMD9PL9SoOUgD9OfijMk27
YUBo1BiUbeMDK7lvj4dKNAilqSxKfcKG+PgwAwwE3dfu3LdUMGZXDyU0kexH5D+9
DZjc3rJ/biyXHoZ04RuUJIOKlEzKYNn0UQ17sZnYSv3l3loKUg8cWHEUqy0Wdd9L
Sjl6IotckoTZ2LhwGvokGbMNSuVJw/Yd9ra5BPKkaM4/CzINIcUxi+d+29YXkGBO
G345sg6MgIs1OEq7BtGl2gq2yVk/9NPR6pMo59Y6Q3QheDPqrJIo8KNPCRJ1ddR8
RtCuje5aSgTIcduDAS8iqeoUGGGwvdfoPEgFYLFIrjhCF/yf7sf5WcIInw+K+kv5
8005SbGXC9H14XS1ZRfQFVFnOEPlHQd1Ooec3LRZlDewHKxcf1O3ZASsL4E9Io1v
kvqqXpGfymNZVE1sK+lpvOc29zpwNd2JtIxItpgFXloaOZgxaqJxolUNY0WlJfkd
hQRlbdJxUsdj/IoXfH8zHmTQJLfOWLqOvJzl7Zf46L5o9Fgyuas6+nAH4KxwevG2
UbvFkMrrtHoiSKLsf4S4tRRdrt0qKyX4KVM1cAWQ4NXN9m3TeAHVwZ4ntrX+13Fs
oDGKtO5jRBROJ8zIPaWXNfgseL9/RDdo+KKiqb3gC/e1fs4yrPwqORlsG9dzf1PF
+UrKjvwXqkxwj+Bs40gTlDYPNEZBGMmNZF4IL7CKpjFR6duaqRQqi/npiuV1SD9l
wPWkqZKGX9EaCAHSG/kQsS6h69ifry+66A32kcJVuoZmEf64QvGH7tW8nokMdEOB
oy9UxTqKWTkR4DNz2MTXZSKLnnPQRqDo9qnjEal39hO72lTFqByaJ5PNDhgI8+fy
MD75GXa30LD8sV9g+edgZo81PWkubEKD9/sN2UqSjf9qwjlDNwrWfNxJWYE7mROQ
9ng5SFzdoUd8aO8mNg5+8JzOyelcKPr7d5DyXAU/UVovSQqIwz4e1cm5pSPQ/GwF
fnD5n9ksCP58nkf1o4XAjdE2EHdNfBlWzeYRgvfqo8XKMUQVxgBz+FyYTG4lBP5Z
WDPOqSfOQlaYLWHVYczkC2cryxf8EJ17VUSnE3xGyK1pApoPPe31wMnMHcylnYSO
VoEfus53gzlv6VTVBwuj3pSn3GdUyv4eniy0a0oTotI9hAH73QrQGUHEYfsmpkGO
iEMtShUrO3pgiUQw23Y8teTGIilscHMuSMb6kR+k5hL17EGMsSZJjLpLwkTayFqJ
QG5qDAMx8fEB/s/+Tbyhb15KmW7s9XEM0jy8m+hpAFY7B/UHSB3cdXG8l+yT5kAg
beuVKbtMtp62VsJhaQPfixOPA2qdfYNKB69cK1QjuZf/KCekixFAg/wHcfs2uRkW
ZipRHdfsn/RFedRsdNnUtiHiIW86DUQNsZEbH9E0E4WIPFD/+IDlmXEJKyHaGSsl
C6TwEjFhqV1yP3oS9sJ5zr8e4URB2HWLC+xqvrneG0EKMvuaoBvIPMtGJ76aeq33
uMdLMzd0a60/Zc/QkRbtGrNm3WqR+LP/Utu1mX8I0k/wfIXYKCeZHV/vhwAIUEoI
y4vzkOyw4GZ3ecMTnMt5UpNAdvMv9lb2+/755EdS5S16d96i3HlCcYC7QWSkalyn
i7+LPasKUtHers+20Ax2MeR6lTzDiyor0t1WRY+FeOjjfGAFvnJMvRwos2jIwFBU
s10+RJdpnanKYcRf/DJYz9OGfwHMrF1tNOq4A5fI7HN2pcFUi+WM4OBwfwzOYCAf
ejs2zZUr48SzixKeEk5MpH1PVYRD6Ebrh+DcmPMP3T6lwmlxMmInH9CDrsF3Siha
b1RHkVOag0TyJFGXDaKIva0B1aUL9RWoCiQTFZrDt/9yYsAazC86nHqjQA2qOGB2
DapL8RSEmp9GKFOylVV+tdbT5mhxlxLvgWN1II/GLcB6FMQgXy7G1Bp8RvxEW4NO
cgG+nglN24tArRNtm2GpkxpEEL/yXjWDL2dLdoxxPGDzg+sOSm39HReTo0sSqaim
XM8ASWuIVlJGiq8oYbUx/6q3ypeFgOeRXmRThaBRjpepkiBmLC0CnejtPTmCoydB
X2U/zWyGOe5fiz9qLJDsjTcnIBzrzulAnrN3K2PBiQybxOVkScrxFeFgImQnA0ul
iSDf42vcb4RMeY88qc0b6MTEHk1/UAjdEganltjHoneXN6nx4OluTgIIpWjoYFmS
UjUlkL3S9++iB3+MIHIyT9RxDMbIq52Lk1eLvYjgqsRM4OwI0EY3+LriDHvwGlKw
/BhiUIeJsxqlddIHmfFkdAUsqTd7GTXOXDM2zNbzexDB91fCpbaOprYOb52Hf7qc
d1SVmS4uXKc+Ndc3QSjm2K1XgVC6zpFiD8wsDFP6ZGrR57Tuq2hOedzHZJRRMMIs
cHr0cB4v02vtEwxNYn9/MHdU/aqagLWk82xoAWKV0jP12SrGvElB6HdJ9OiZ1COE
zXY/iYn//36EKS+SQn5zh/RedvYF/imweklsMeQQHEgwNl/onuU9+jpru5RRCRyq
FwuRB0Cno+D2fmp1YFe3IXP158MIxEEY2pocO1qJFi5B2aaiEiTxbOWjvwDfvMP6
ZMxUcYmho7FiYQ54Uc5LUemJorrOupxOHYZ0Xqny9hVDtLoHeND6ReXprV+uBg+8
bkmg/xbUDQay8v7h2pn56Jc78z9rGYs/po5uTW7wLPvEvk0gH2QFGMfvRl2CpLil
DLqA7SrR24tfFtPpp3CIjEPug2fg+0binXLo47INvnp555sKhq+qyJNaf3PY0KfE
J/2fOfM9JuLnp4nTdOl3BXnJsU4wQ/9TNDZd/DnElguFC99BLw88H9j2uUEVtLuY
tNP4r2EZqxte8cjt/cX6/bd0WAirUc/4e/ackUyKIaAvkC88K3WkKrSx+3Ce3JUe
j+d8yByYi7nVHrbtiyUbK4lmINhF8neVy2vVdqOMJ0Abra45qlLHELoQjKeeKa7h
+epxbLZJHyHU9J2P178fkl23gxoARqoEHMPUPTCAJ7YHMJhCiWdCj44BMb44L8A5
/Vfdq+I633zylbmTdshRbhpUccKgb2XeS7kdgF9pp19oIs8g8rsc+Gtgp59kcVMS
EFib8mnIwADSTYd1fx4nWGvYHWZBGksOFwICKQRhwQS7wuzubfeq9IE26HYskLlX
9KUuiU78Osk4prezJw0U3MlU7ta2bjLRnsAAhQHo2Vzf40FSGxApslltlWV+DQIy
xRAjuFoG16iSlWpwg2RkKuYgdDfV+Be3DrA0clXCD2sqsTL04f73aiYUVNQnooKq
58Kr5TLOyORKhs81C4q9WHbQvYsKEtCXrRDJMlHDVTKNRuOaLLmRL/KGuoNbfzn6
ShzLr+2EpFcFFXyfuEx5ez+wSHMCDc20DoFSOiGVRJ/YeJTQSlQGV38FJNzh66Jv
1kc9CBsL10ru/NqQJdsuFIYV59bF2G2qFwZqKk+KrBf+SHr7cRiayyy34oIh+ta0
FaYpbAtdSpKectc74q3uhDeryQAgLBsnmBBr/39dRj6lTVy+iJjViEyUXzbZsQnb
qrNuD4C8S7hn5tGd9wcfK3/JPcPft9og9cBfP9Ms1gdn05luyTll1POTFQoqyEsT
mbRWt+sceOA3di4LLKcyx8emEaUgNQoJOMvuJ/L/FCLlhwRwMAqibLPNzWLhMfvv
gN4qqbxf2TMF7QFZeW2WH93zxmmcmUg01Z8ZAjPDcce40ysXkhrc5wNz5RxcmyCv
LPLAMCTrWec5EzE3WNmtiyVN5M3IlocIZP1vDffIPcWMK+FNCd11Umf/uakEJT8h
qJrXMRipGPuvXqAcrY1cD8nphxuBFBOZQmS+QrE/1r/AYUhDnYmlYQ5V7ahFZosb
1a7iw1yFVyj4OjNZ0eco1VgKaoQezhzdqeNIPPxjuNFkBHH1XC+xprxuw8S/n2QJ
oMP+T6LOZq72RseRG0EVnraBT6xqzDuHE/W2dNwBd1VFEk4MnvokucT3Q2Pejtcw
646uyHuFq3+ey/5dOPnv90l4LhGy2YX73RCnUugBifzmRmKj33aJ6RFv99ae1RG3
UAWokA2dGTXcBQrD+7xAWzoQse6Ynw2pmXshh8susOIjloTGV7LxrEB3NuQbkNhn
68SpoSl5TnPwb/zGC4zVJoVq8JL2WNY4PdcSMk93XVud2AWRyDkfY4I92/avtDc6
g2uXCWd4QHamLMgOmP6v3f0UcrXHZFjwtyTjSJQJNa8=
`pragma protect end_protected
