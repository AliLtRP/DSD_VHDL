// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:31:31 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
FKBChaghIOsBxMo2fKV5vRv4xsZfDGn/Oq9lbctnJ2vMSqamILtEXfvXGhvAAZA9
R+42cKUarj39muavpUB34EnaATKWth8wtkC1dobOOoXCPMtO2ys1URJ55Ww2B7es
bialyNUajNoXM20Dp4yUzec2KRvfQEaYYo9O4kcunCA=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 38576)
1Ph/Y/kiUXESSrhOEZiuhbZVu7vUcKV19y9mPPzYLPJ7i9N/BlqJc3NHmLDV++Jr
f3lwadUExHBecUDPpfVUIeHlWR5cqigN8YHy9HQams5FH81EhaQwzjD9PbUFgeyM
0VbhyY8ftgUlPzNbvUBARgq8MRIsllJcZqVp58o4d8G6FpgpSlFQalR6vUN3LFtF
i4JU4AGWQA84k/UDKQ0HJESXZIqK2nqcAF82HugRPLHAVsj4yQDNBGL8K+SPO6Jq
j92uYU2uB83enxjCJ/LI5FQBASQBZKwKAct3w3CP+f5qlHpJQdHN60NrBwB/ep6y
aRqJeUv1ApzVGEXbC/B0daU541c5Jm+ylrM07ML9u6b38GtuRlAndUxHT2lH7cIK
Wp4AqgRsugzkdfj4meOY30fzbqfZwc7kZGe1ZE33nswk6S28kwoMKHeNUgoJr9Ti
Fkyk4YeKW74E4PNhVNQP58e9t8SidT4d0W0uIcxGSO7F1m8l8gYy3IkCldU9dwNu
qQk0yYEoG14tihgTK3pFyAXqOqcAeBJdHsRwGQeKUAiP3xQqYsf2C/S9ZekovMzz
lGp+0+pWFHyA6Y6XgLXj7PXhKzS1Uj8HuGalavIH1Ni/wgh97AvNtdelLlD3xo0W
AyXuxrWyO7QbF20EdnnjEEguc3/hxkdF1S/dNITsWfeb+GJpyZlknyLReHC0iQSu
E/7ZpBAkYnscGyRC0fjcqRVe8cOj3VhexOwOkS8hnmIZXGuwpfnKZfcHW4OYR3ro
39vnvn7UzP46Q6yt6Tdma0mqrkaJ2NPzNL/KPzgtTGWX584LczL6swQcjMstyN5p
alRkMj7AdVcDQCYPOE+vbdKHsmnrCQZuEBOiyD44gqkBgyF6GJJLyXljQOA4sTxq
8URnHwQEWoqK3xb4gfs63iM+cP6w1WOWpOAemD+4TmJNKIVvCiVtHOm3mYfrVxd+
P/014yEYLFLOvwx++2bLQyJaMWGWJ695DRCn9xlQQYUMfGRYL2eckVNHrTj3WWqI
lZIPP/9D4nusbQhL5ZP+eonOGK7vQJbmdbX9x72fTg59nLproDU2bG8t8ThmTLLP
u2p5rcIHT1mbXS724GMafikCr+2IxF+Vkb8+Rwd+YqLrucagBnczT/uG12GslXGR
BroYKx2do21g5ZBCL5tzxeCsnAj3f4FwxvwqC07cJlHPE32UTCGi3yp3y3RsRX1U
GRYifAxC1ZBGBJr5v5hP3lyo5t7rCKZOe3jbTed/IItOXxKrz2r58bHFKQOLaig2
TqCUfpdNCPu+0jnE+OtVTVCeE1t0rMAJYABLWNh+a4X188Bz9uhDaMfuGTM48bjA
sCdm9MVUjiFl8c2FV4Xj/ZKTXpjJLDJjOXiVuUL5OFymwILDoC01fobdwr56jdt7
cpvLi0gHFPJNqeQmCIbXJTOU+mur6NmQj/8YQ8OWeGq3C0CG5gOphkZIXLxROnuI
IVVzxqhYhEdR2ZF1bueUfCiKxle0pShWwH9yPHsRpc0uT9+UCsCQGMVSq3wjw9jj
VI7sc/qlEOPc70jJPN4gZAdC8HbH7+eKG2Ldimpx54H8hSHC08t86CXALcC1ayrG
tMV83MfXS+rlRKDh/feN70ADrUzEulTOsetY42sR9WQJEA6WklUe2EC8+v2I+vNw
0x+WR6gSMqjIP0vOr3z62Uj/p4EirRdpUlLkOsaRmr5KZmG/j7bDjiFmdfAbewTh
UHSG7LSlNSn3xC2daJOGAcxaXmXODk+7EO10qvWQ0TrVBwBVxWxz2tng2gThQ+Pz
ZG01bbfZXIaY5as4M4bhNYNTWUXcTPj4Gu4AIOA4gXgyEu0p4vP3ZLXbQJNE6CNq
LjVtY4u9iwcmNZhqMfwoj29a7Zj/Tl/182Qu9EkIw01IU4jB9MLLFabZ1hpftJx+
0/jfq9BCrV1WpymMxe/WLHyixlhK33RhZda4ATyEfAX+y9mhVL9NgfPUNzQVgZFE
fxUTjAjr2rSOzVnWGbc2yZfAGxd9NNYU2oDQPSXpOJlDcbQBgR18ImsNbOHKznXU
Pn3znq35hnscjaSTGpmQ/s1evoMsbmBBjwQ6DYqhTS6iY2alPlYSc6y3XNzno49Z
SFdrCmWV0uobQ6qD2N/knHmckaPggJYZoZkSW63qZcLo4IFi6iWfoDuyFL3vrLX4
fj8yqDtXwVJiScoUd5aHptGuX97QAZFPvqop3p13MT8iafe8o5f2xBXMbedSpb/1
JyZxusu8Q6Q0TaUS3raiTis41orxp/8kPZBUgpvZHfyU3rkPOHn4gAp00NI6YrpQ
6Oj8orfM81aumchyxUAEg6EF4aL6q89xoCcFYTZy/4t/tlVyNVZMU+8ChJqXWWTC
JFiwnZerhR6UMOO8hyRYQkdEsLIDxjFIFrijzblZrh5/0n2Z6JNM6hOCk/DSBQPS
pucPawg2Z1A1Gmpa5O1/pz8AQEp6Nf3dNNfiDNvdtSum5Sz7ZXGmxmCNx5p1+DG+
eFIiwQm5ibw/fU0mOQnfYn0veZjH0xeluAo5rwy0ehmDUOtHG4QaXO8ZjWOsv7qQ
qB4sUFE7jLSa+nvHTMNvp2nSP2VmdxhFaaY3dKCi/ovFGzrsFCD8V2w+Gcb83+nW
UsivWVs6Bfhero3bh6A66keHkClr+3bWSPSL9ZPUS76D+IQRWUdr3UoV/Q2n2OSB
0j7kRCmnVVZbOf9qRazBfsMNDhnNITyosjBvjeF6I5mattn23TOUKJso8FmnDips
qGQlE4J3Nv3VKifJE63yw7Vu+ARUCjqi1SjSG4lQyhi7w0OQjKlhkSwjP0ylp2u/
XHQiUHWjb7MHeEjKd8BK2Gs5oRSp3N9HmEgfdm9n7xFMuaz+HSo+W5BcDm1A9lz4
mbIDzFA8iA5/bgVJqhKCaDcGcWURiOzAMgKKdUYCbOiZV7QFoNBVor/9Ee9G6S/U
hhJb25USa1Mvct1Xna2u2o7XMiQFsNeL8HLiSK0jGhNqz/DS56eYyp9YzCK8YuhK
PjDITMEb9/doi29VpfaqohLjZ4KNlxTfqDt3h5VSbr8teRXYfPXd4fjtQnGJhs82
hmw21gpZmzCvages6HCE+jh+8XiqOxe9NU6G+vX8Du7JB1qB13KhpE9TneytdQrd
5aZZiBonnSZBUo3/x1py5D3cM/ZdN2lOVAVxavTC+11nPspg/wIU3JAFJNJAUzZ7
VfnpSYhhqn4ETRIT5ng6Qplnedw7JOqxpBxbKAEn09anZM64S8uzm7PVGoD/i6q5
cpADAQXU4aPcbcILK3/x3mAsAJBJ9VqIWp27A7DLr64vtR4psA1ORhEi2ayLkTxb
E0PQgphmHFan+tIAmffiEmw2Nc0pWI5utFf+ufcEChrkHpDM+Ypm4cd6tcjg26xg
I9Dh+Ecyy2tjLTcmRqTHBH6iqQQYjRJrQboXsZVZc1XbtCuT7FyQtyREpmJfATEh
ufxDo6fhvgTiwe3UzPHCOWEJNaHf3wufkMEDE1pLjLEYG4GYoK9bN3UwuubFYsSs
vD/kUANN/i+Se+nkDhzj4R24+taPBVwoW0QsSXoHCU6XpOB6MQQg66Km/i11nZR1
wMfmGboXIYkIl7TaKeEobzXIC4QJ3DdOauR0t6xC9zbD31bilMsoQ0aQ+0Qsliba
A7yHNikEnj9eqjSDihvgjQ1qPZrDUPIozyptlVR6QtEtrrV5yncj3HY5iTPRvm/0
wZKnb6KMLDpaUYwSnnp/byH3xHD8Ng3QntpelFHAZC2s8qCn6aRp/J+uDscZ3wAE
6AbdmFKJj/vO6hJiGQLJFiKbWrU5bZ+U8Fc7q4BEnyODPhtya/0I0uEl+yO7/lMm
S+o8OBzVguSxH4RWrFMrO0g1jADGxF92fux/U4vMytK7qXcg2K4gwFGUL+8qptay
MmbI9DrusP19oLSXRveuzY0HF0NcQH/YraXA1qqcF3otEI3r/I4uRxe5o+89I8en
D6reaCGSCrNeDk7T+a0iW8jsVk7eL7a+L4udrm4syS76mRzCAB1ptel5gt7PbuQ1
EGsEL36PQNmWA4oWxE8EjLWmy/rTy/Pk3lJz5VgF2/j13If3ThrOjLgyYTInPYxF
mexNpdIMBssEK36pqIcwAfSnSSOqzGfcREPzlm3/4OdDP0lbkYexjzd3/A0yeBAC
MmJ4xvD08msGDGkZPMwBDeFKm6/04wFoynYVsXO4yEQiESUHcGdHxd3qPAHgGfFL
w+1NYkQsJDL7O1pWt1f1+Kt5+xcuZ43WOtzDTXVcaJ8csHD9shnRametEDkX7niT
2ihzR1qxNF7QbOp/kED+5rKubz1uGf6cbhzlW51sXAQO2cNz07e1cosN9K0B2blB
ZAjVJoDTYnnKROvLa10NM7u70c0l3iMeU+rm6/NOh3WdY3DMjzzOhr4t9yjK4hFP
mlS4th0FZ9e36U+dlUzYalT7X01K40biYVzxI1kkFeJR/cGLeyqIq60Id1zKrec8
ZjLLwAxdC2mtNHtkyzdc/Q1+REd4aB6KMp0//RGWZnVi/ZC2jze+JIjNdIsq+eMQ
K1c2eAR597HkFjwnjS8/THtgaFNBxrBsA9FtozlE5a3pbEwaQp3JIvp7CMiWiXyh
Kxt5rIFtaOGGxkivboDbdxjaqvos2rLajOTmy2g65aPP1F3x+dzEEhlFV6PCTbT/
UlZF4//7GeI0J11fiyttsPwpUGWfG7XvED2AKkcsLgDpHgsx0XW7aaegMyEiPeED
Cp0uu+PutNmz8fhaH2Mf4tEEVIzd5xLG/3ZAT89XcFeh4t77BFG4YbPP0/K3Hvig
xuJwAyc65GGpUKGP/DiMp/KoXVxscY1linmYa/aCfCRlxGqAqSHxX9bsftFVbcHE
vVctcmEZ7UDJxVakhNzheOOiNaYBffJp5s3KTP+AjrKWLtFGf4pK3Po4mprO5DRR
v5H/oGKZOBwL+Txn+XlPZPLGF6ocR9K52OI/v99tKy5bsgJbgti69c8ZkMDuLg6/
wYX05dmOVmLBjlmF+ZV9XqrDnWFoeRFAmyIXmq6gF95X1GGKg2dkFhsocP4mcr2x
hZi+Ytz551o2ByuVrTwIWJSEUNSCAbwEV8oLiXaW4xKpU8p17qLjA9YzPoBKhjPi
W5sQ2UyeTyIQwUc2Su1urVfXDEi5SfhjgEEOvUwirUQrMuIn33paKPUy+G0eiAPD
4SVlUt8m+qJr5aeXYDSDIVUpoEPv+e8urfIMKixSaX9kMwkpwo6/EJBKif1zH3T9
jbWnpvRiEVTyecIkDiZxPYnOs+oGefrjBDXBaALW2d1rRBWUHknfnL+pE8mNBB/r
uGNGtljB+nEDqgON7LmJ3nzc9gt+t7TPb1C8nR1+PiBvUSZucbO71uSYb5mNj/N6
nv0ZELJX/hiBFohUKUFqy3DcVyxE9MCrq2YQH8LOsSRTuDNk82SGPkC6K9eEHrGF
2s0MchuREUGE692zf3fCU3gh7/Ui3pK854omp0oucgnQuXVJ9JhoR16YYscUMbkz
zcSg4yfJMwtrvhfOfo0FFKbnKp+BzM35v8GtKIbvKVfeHnT2MKXHVYv5W+FWdYdV
3ScQybG6ocR39qEAnEzmz7nTTH3lhACw/SKqURDGljnew5tuZg421UnwMO3z/LE9
EcIwT5Pav2dNfN3YI6P4I/vGyQpPUWX2ymYZdNBZD2i/oUdUnBPuHiLijiyepBD1
GtFmy0C+N3FDO2dePjrb2fhZ39c0/0sNd+91Ntuw2L3/JkEPl5pqaSAf8FlmDtPx
ZY59DNOnXq3PCz3r+1zguTIAbH3n04TZDYOO2+Gf8rVYVIjiekrJqq4Hm1IpzTnx
U5GGymesZd2wELCy3YK3T8/l9XN4I3gJSHUpid+BmGbB+Bil1g4pIQDIwKSH/Fao
H34ECrK8d1LDT4VgZS4eAPg7G18VZrvplmanIRlkML5jAGSExltP/7OTZkoeBELS
MpiOLFOSnyBvh/XG6BsbHIknXSoea3t5QMxcW0rA9PFpu9wuEH1TOm7CKdjnOJUq
m1albxE5kLV+HgZvJw1zsv/zWlwi7FQsWDVI9o8/I8XBfZOkvodXQCMM0+UNywF8
LKiJsoJkTlshj40FVQdawjWt+AjccpeEiR4gW8ZVcQhqcWqYuNOmKU+lkVVkXlnw
cgu17T9EGFEZcIi6r6n8GnP8lUa9qIWboIx6s8XuU7GbBcQ749d4Wl+eyiIQo78C
AoNER5rl37ukWRW74Gj5YLfh/6vOzmepT7mLtbu1Ns4EPs4EmLXbnhUvkp+5Iahy
Zkr2JebatFH6mRaOskJ1wQkHHKE8KNqtX7gY2L+pE01IQcoovHLxbWoxLyeHIFgu
R0fVG2tQHIVnoOqiMAFB5dvvDRe2mbslmcldZFJOhDxZkW2QXVeeY96vK6pWcnQ9
kUIDupEi42Ue5xkhswpzQQDfXuxGMNNym+2llmi5HtnErDG/9AL+7QW3UHKdEYdD
Nrzv6n+x5tjknsfmSongZKdHsOr4DAZ10i0qJsNkjtR8RMpRh01wvTRt+o4hzl+Y
yMRS3fExQUhcSP3mKAzne8ooKir+MJO97PqqFaRuEf9RWlwELtwN9vxmSgsb2eH+
h2KsbYI9pzrDv9KzqMV3J9QTuGKuJRA7AGvTB9YyNZIlpJuoPZwdHRGgPq/1Oyk2
he77T1mS/EZOxdSmva3kXD2Qa//HLlVJC8Dx/q5zAbPzCOPye1l5ncE71/uSHx04
Bu4sHUnWu2Thjy62aVTpnnJRgMREsgVXWqahprZDDOzfvnC6a9iDLRf4RnmtIl6f
FaySaa3T6Dcw+Z8zDCOjNygmUUV0vMsI0mrTGZAubp4Lj5uf5Wfp2skToXWzj5tT
Tz8hGYOWyvcInrvmaZR4Rf7BBz+lPFsJOGUkm9LywFDNu045MNzqIZKJICbjdodu
dHx9JrUoFHPEAZvWuWe59uy3LL4OUj4TVMfERHS5AybR7Z6ijhLpgf/9qdajiNX+
HFtRgFIpXE8B+3zSmdn+UKTCe8TpTw0YavnP6tzWAPn2aUsOsSYBIKj+xOsnBwaY
rr3SVSBBVvmU+n6FRazGd+YvZcyPaXSaBV9ODpD+pMuPOqlz2EEZ9OxlCK970uYv
QqqoEWEyoKinpK8/2lm/dC2bORnpb1R/Hqd+fGeH7CnNUyP+2l1yiMoRfHvVvfAM
SlEy4FJ1FaKQtr0oqwW/ZU9/9elfWcy5/BT3B+kdckqiLyYhoAGnYI8f5kTIqUYL
ncqkcEUz/yUMsqohyxrXXEeIp5XeG83GxniCN0gIm/tmbwU84QFwMj75zrkPklLX
MWfEDFs58lTYTn8/mkJSECr3sV6oM2urERlKX2/vUk7t07bgIOdEjYyDGRF8uzL6
Q4+qmuMia+E7ntxfipz161/nMF88m7YmlD6efW41BcJwbbvhQECxLRxwiZ0YYVIV
o7O1W8HsIscwM//cy0Jw+2yVd+ueQ0cl5rKJxampyfJca2EAQZilbVarL8Jt1rhT
Y+NRJuwtwuY+Y0ladO6M/4iEBDd4o40UeTWB4whrOhHrTsbN/B6dgEKdO8OTGo5f
8bKdxdDDVTTz+hV5Q53ai3QWHDaQue9F/Mqnk8NayXv1dX7vf7yfvycBWgk8dNbH
c4mhFiIZcH1LgQFWJL75qcRi47yhz0sKNKg7HgRCwGdVeScf0uyAoSKKYxoNpH6/
XpJPILdcVLDjWfk4e1qLkvs2qYIwvO9ixThDobtK5RFMkL3TI6604NaOi2XWEjTN
ex27i/iuh2Wfh9HAykCQsj+oKx9B25+C+ipP4jneSgTgGckOQIJFWZmqnmXRjeGH
Nxgdy65HfNw8H8tznKEXkH8T3DnkiaGxCd35lT331cDqtNaDFfvZ2DfeNxZSs3rU
TnXQTo//mChKozBebQVgXAWpl6e6WN27uWlOoVw2a4mQmNqkOoMonGvI2nZIJmHr
hzzgA1IMCaoPcjmIp9A446LaEoMnE6O+3m/H2RLPSovug+ntzBxtsiz9n4ItVYzP
drzxlW1mniS6ONtMP+bVrlJ40KdL/roiM113xvFpUQoyUR/F9hAO2DXIWhCGAWuE
Z9J1tN0IEqzJW5R21WT1Ia98pIxfECgJysbU0U1/VfaqoM7GmSoCG1PobM5h81Cg
cOrz6MejXFYgM6CNIUEAwrsAL4rrrLRDlIhKXGMuG23sgt5irLKTxSQbJO58hVM9
o7yQ9Xrjpj8XNeVCYIa23aCqry0bAIbCcGMAwPqrc5QZo7vXeM7mJUudW0fewST5
MCFa/Dnepd7g+kkiBMNMs78Pp+JKtYjDEdoy+F8nWEjcVnYjR01ViicRXXe+8eAt
kbp5UqT0YNedkObCFGg/prB5W0+8q7ykOwjLss+rSx/MeX9DmFc/H+OpsNpJ117c
89DTqWbDe9Xyi0pTMmDjBXZDwtWBG325IJJs827JwcSNqGUoaBJ3MpQSljc8FLya
Ul93tHjL1GQSKaubXxV5Vjab4q751O3JAom63/g/+2act74QJo959LnGe1yRHdeU
u7InZH9Y4Zxoz2b10yBV+4ZoCQgCetAuepSL6uXynryX+517+2xTHpBAi2TQOBhw
UbwKRUT1cbyw814b6ED6E0nvr6K+zRWxh2EEQpVH316kvLZYk9rCGAM9DZsmVnuY
vAvFz+13NgvMfCGK60Rx1mW2+rYQU6ll5s8y9JgRZb8Gib/m2VoqdMcIK4eM6EmZ
woVrIykZ0MK2WBlFR65BTGZf/1DDbWCmq8SPKz5gXZZ/Oe44O3E7JYEA6wyycuaR
ZiEk+SqkZADfdbOFGK9pUzb4k2X/LJTTPOudq35Sb0LvPDPEed4khWDlHo7AEr4+
mvZc8NQhUvtrr81KniCMZhter0V1eFSj+A+Zx1uB9LY4PQABJBOAVpE2odZfrd1J
s5fB3BNLLmW3E4Btczl99YMqgjYccSdHvIMpw9U/c4TrPFPR6S3RCFO/qw6VjaH0
zvg88XA1a3uBr+ubj+3TnaGL8b0AlmYVUpGOTtuVUOdu5AEnvyZ4uhB9aYJl78YY
4M5+yiXHift8roZ/8y3pVat6STsEMkySm6OHTVwUpOoEoOZDSz6vQSIDXPbTDHOU
nwVS39nTHmXE+8YGJf3VwnR8O+pUP/D8ozsNEhCxUillg+fpPfKUH8V4nER5B+3h
T7oOn/JSbgHcOTK5FEvZsrCp46pEe1P1/qble5cf/oWOP+IgE2/+Fh6gIxXjcHK0
eq8eG9VmJr79ZB7c88ZfB4kjq8bYMP/TgqzSfYJOxS8+vt5pi3Lj8aD0UdLX9ywW
QQ3cHxj4f7BTfaHaJSlKSgEQOsSmC3ze3aoM3MTm1Nmgnn/lqf4V+0IZVaGk7Rdy
RGNNUck6suQ+lFsS41Iw3puF4E1xqmrssnhDG5PtC36e4axIIhQaxjnqYkY3vyD6
ZcNHwGKUx/UGDDSBZxT8yV17kN405Mksy3dCuL/QncBfF5aqsZI4ZVqKYqWcF4n/
V1mpWtds9y5UGm9EVEDG4JBSMMkhVbj2HO1lClIjZEHQYZQRRT9BBsiCg4nNwhp9
SHSwzYVrBKpp6lPVF6CcAGk8/WpH0NSDzCm6o6iZhRGGq1JfNjG4zjped6I01qEB
rPVqty/AHeW8/0AsExwAA93r2CyOOlM1640yOQOctci0sT0/I4on5oQ0C8IQiq4q
4SK2Fl65c5eANStJYhetmTbCjtr5M/bTTcfM4+bbddHsN2+VF0NlV/YXqyqR+eFI
HUNklKz3nNdX/JgcBVu5QyyCM5LQGbkHDPsNdCd7qcdIpCsYtY6E7nOxYI0sTi6z
mH6LEXXTMEDGWrkuYFuDeDzXCJ571ro0gWB/oUWsJHB8NvZDdKW4EbnOV8toagMx
+6wYjdd9tacgo9uBC8CZ8GideTTR8F5N9mALOYw4fKUYwAtr6A2pjHkD7bzJdzEk
QCAhDNRjO2Ewsrtp2CyPGjIzzUqBtwUL6RlfKAFUx0nJ3A1fv57QBdOHVTY1RYjk
Q90p4RbEIQ+Du+FgRhZjACZIag7QXz4GSoAh1HO7s/2RDOKUgyajpmOJjD87ZyaD
hPqrE5OgQYbnGJX4bTiNkx8N+CUqL9Hgo3uygs0oKlSzBnN38vEchOeTf1yVYTCw
qIBSlAr+EiOEFnql6NRSSqdSfsQdPg8AV3UgbPZ3PO6Q3f+ZIih2eEY1O/4kUeC4
jBN98kCG/Azk4tyX4N77G9kepQLFYMglt5gyF4ZBwhpxhqknsTS5tm4mfDBGq8YE
41BBQtuFz8GFDZm8eHhCOVkLMm24spLOO3dMVkWz+qX9n0WLSPEOQewzkp4b5VRP
NmBRqAJH0s/1FEj1XD18X2wwH8wH972sHdNZ2b+CuHDSdkIz2kZVngLgM+LYVr61
oLZuZj+IbCVyGCIauOcQwEtFW9+lSRWwaMGGjAXa1kSBJoE551I0hNoxr084a3YV
VRBCQ0nrhSfYs642l6KwzzNB33g5/7SCgEzoweTj2oe4OMzCPG5pixFhxhR44wp4
BnEatdYHYhsd14LPtqUMARhLkIBqqHi6k9cWTHySshoCJDrBOzUl9ObNAPLAIrAv
a7FNgA1ZP/VOxtHt4OlzJ8Nn6aAZyhcb/iVPl5Pfq3jwLNw9m11+v9fmA0x9ezx4
NQiWL3mbabvSqUXxTd80ScV+oDJeywjacLVdYxfdIfI1onRkjEZg0Y6749l4NP3H
ThqarLGckY02idAsUlt3xq98PFknaz3rAoxn9IZFPJcRSotdIp4lnQVuyPbX081+
+GgxhrlCs8WWQN4UM3Fkx7i0o7mFZPe75RRHGCmIfnGxsln5GVNy45O8eLCARkFZ
PclMZequ7nZJe3kxkT3P0IWT84RgVzF2qsl9dD6sLEkaXR/gUvcWb48+XaAzP1xe
bA/dvg7PfzVgpaL2iT9v7p1miTzV2okvhxv/az7JrqVxy4KPAMZBaUfpeyKK2lch
9rDjHYn5aw7upOIMsxClJIt4HEqfkR2VG5+huUdnV19Pmg6cvO7H7b1uZf3jgOre
LB02JETSqkoUMF9yapubQQs2f98E0eNdFr2ktxHlBS/KmQNQTA9/Hpas8Z17edr/
U9pfEDo8XtLS2jn9ExiZAwYIJSEuaKWOJv+j4vwDjJbxKthjIBqm0UY/Wm0V9mE3
ApK7DDc8eMh883HnH8hDoD5CkriZEpqS4wD0g9cwAqnNhEGhUQhwuYG7PZvLTPj5
5oOCjnwueFkSgTtucwIH3dBpC0/gvNhY+MRE5dJ7C3LxLUSmafbXVV3rfxOzEmHf
UwEtBa1jNfH/pCW/JaNs13GdnWfFzN+ELW5jTptdugoPH/BIolVY11EjL8x/SJcW
mXFAQW+tICuqzPT9kWU8TRD4vTSEwe3d1v4KmBbZv/2A45rt2NgqqsHmX+ZTW7Wa
WfA5B2lJAvP9hHA4AIrEb9Bdjtx71GG1VkQBshdVaY3hf3wgehJnXMHjmLTN8kvR
SSD7YZhDP7vlJ9B/siiSRT4NqTw9DY9W4TKPrXQvLEq2ZHZIPapUl6W6XoXZt1jK
VAmLy7XrIGIraPDVL+WX6WQqhiOooZKcPSr7sfNT7ERPw/7ze1H7qafLPUehnqn5
thC0q9WZoskUt8z8L+KWf5DSwkMjOOwxMrxjf5pBs8cIPniRmFJfAf090yuHYyp/
dckgBZ6A8Eu/PN4hTMVVs3M3loAVjGr4ZfzZAzin0bhHxlNc+mnUD+lkMaP0oFrY
sI3nnFtgl3IELen1KpgrrioBrYKDun3XcU9r7R9o6Pca5ru9cdMj6XORAdWnS68m
uBvrMhUHzncDKxkZPb6SaQxTVEIppojOOd7H6KT/t13DkyJLseI9vaItqSJb60hQ
zYWlpof3j/BBeV4Aki/ewa6A2RmGBVX5U2Wid8YMR9Yz+nMKRhj/uEOJGR/jFtgV
R2tXwBD6cIEu9XnzLaZo5YTrff6YajsbdVVilvXbMrRuySTHdPpDfPyQI954rQL+
LPjUTmPbUYEZdIRpnRLGR1pFG1R2mW+S3MLY2aECdpt/f+bxCunStrymigUpZ7ku
bgWO0DPs3NlUddSdRy+LGav0K+c4pR0+pOOpxGDX9Kx2QMutLgVqlzGrsjfu03DC
CWsQiX5CwUxCNA5U7NUCoGn+9ypE8fMrI9/SPxJwiGJA157jxk3JgoBWgwdqzPHP
XOhIzi8QOaz7SmjJBG7i3Tw8m5R2XLkKYRkt7h4drlYn+3/PijRNxSxjQVgBB7tg
NCnpc2sggWyykXh+9y2qT7GIfHcHWpCNA9uaqo/e6IuW6CKZCIX0Dgo/Ebm7O94R
SY2dg3guS9YggKkEI9ipMb6ZIaNR8NbbX9WdlM1o4F/nJgEkDT/8bzkotTBFBkHj
XiT3JX3LWmw8h0jvCTNuC3OYRU4k33c/7y3AaydrXSksDp8eEkXHMf3vBFFF6CWA
zvA32SidkLn4DtPXVgzMPCd0fR25Wd7Ptou5w1j6cj4e7LnX8WBmEYZRBOGpWhob
L+dC8P3j7IVCMTfyTl9I4rCNQvQoTqJ3th7z+dNU41aX0iu6PxhdeAPcO+j+9LzB
JAKtBb2/82VRagYSa8o4TYZRUsPFsG3CywfjCy/DXptrlCn/r9AVSLF9uBH4xh6+
GEbVSR2uzmySa8BK00Nku/sz/JYKtRmO9rWGosYy5sQgxYZfPR/VkaDDYZuDvo8H
mfhukvNEGytN3llGIyShzhIx9S/7/83OjDYXB00ZzvCN5FlVr7Y6YA+0UWtk3wld
E6aeuN0waND5zWnfpgaiE3LWofKlzXvkfYok50njArtpekhhyRPZR3QfbynNu/3F
UpTSYeN1y03Gah9GbgxiUEM5m6R2mEoPYrimMt7c71MsWWGrizGWuz88kmLSIVWH
mRIRDxzIaWtyq71qUevhC71QE4EIkeNzJ+BogfmKADWl8P8jbWw6dh62Pzj5XUJp
HuwaPSeEiQEAf81wzBr98GKzWFF1AA4c2DCH4yl0WtLNakyRDn17AqPkfyid4sBA
M8O91KrlY7RpwBz011K2zUiJl6ttcNM+Ufl69o0/4bnJ0kjxr26ZUJlWrE7dJ/Px
isjWWAMkSsmCL6NQsKQz3Z/cS1r93Ni39lSACB+H60YZ4EUgPjEODtRDi/2XZtau
AybK0LAN3PxuZ8B6CuCxk70y5g1YXUnZ7pL4sSbyRDP9ila16zqT/aBdLssWdsHK
GArPsCEOhWUCLKGntCyeN724onpgIA39vvHmiNo6UwRFcFxhFPUndeyXu39FfzWF
ofmCmDdHaVuMj9BXcge5XhHX18/1JkjrYn2iZDR77BT2uC/zCl5sCMRhCKIREeAC
jaoIHbtrkWwGRm2Mo30ImBzR4Zc5FYMkEgjU8IIF5o7vHHbMnhnc4+nxELnMkduw
ifuq9/XlVDHl69NnzY8yw6C7ub5GAnzbPnvbvT55rAtT9HfA5A+A9v3ooC0Tyc0M
4jSTkE/FFCbV2UDLbfpuRffzG40CGFzR4r/808Rs5Gq06tB1xkvyC9BQf0l6IYR6
TDYQf7i7uLesHd0LFEIm51dKRYDBB8zmaK95/jRzL3GEBj0dsm/2TZ2ivee8TXKV
+0sxNjRkrze0Fwg/S15w+HO/csbfR0ZSeoOkLqKPsEadEtrpLOs4R/pQ/UyPmVrN
lBLFxdXRQl4IvFjDGy4JgupP9eUynCLfCF5xmt1BbNx4KoAqUciGESlILhtnX5Z0
ZLaAyno+fRUyERlx22taXPkqfeeyGti3rRfDNp2PdncC60dYmWqmIY4HzhBN9o0z
T68l2fcTedqk/kK/J2ZcrwbuyQXh9QoR733G2lZ+unxO2XHCXHL5E039Jf0JJgDA
kZWQQnbEwah5e8jiU1B2o1r+yoYOKgjLAS3f0ECmuKd/30PY57uMqYx2ginLxCVf
mujGipHMFfaXPlsok4lL+6h9KDx7XhZec0LKjgLDbbCCTWwrjfMahUoKd3JihMeB
50Kvm8EygxJ9EqorY4ErcUhjCTf8oDHYEItV6nnJYai+Iqf569YqKba1NgwkW3zW
4UMWywSoVJt9ifQgokh4iiEudm5o2yqPXY6swOniClKgsW6FMR0VnSvSSJof/Zxi
7WjzoC4XGR25Bx1jD7kAw2UtvlHNb+FRjDcDZIpYSo3lFsNpwA9McTh2eXxgp7Qy
aWRt784gT1KwhNRu7KjSnOZu0N9a3jIqwSNpuVkWTnqyQ3ZiLHoK88fn/WEvF3qO
BKoq4uQ0xRGD2qfHXslFU5wCBxLGaKSfyiNBD3UrC5vZfTS8W0JqCifoVrLUxH24
jt7QinQRXuiUxvFRAosYIv8e2aXpuZvvSHd30aKcuuYEmMyGTjYw12CsN8YpC6XV
5MdaIlXd3y+KyxDJ8nNNZYWvdheYKEk/vdfWNfTrr5cGvA1KORGJC3vmY520ba7Q
KX/ReR3B7tvsLkTWqvuiDstBaLAbeIEOR30dJ7AZM0tLRjwsWLy+rjqdJ7kihKBq
OmO1S1hpgqIWs4fInu+UzD77Oxm29WBObo9VJftcso6DbzbpbMBkr+peYF+zSrwu
Fl+VcRX/kZfAeHQejRcLX1ILQAmkP0yfxier8/OEcXwLPgDkA7F0GMs/ALR0eJnM
q2JI77GcQdDEqEgrZ0ji0Z5iwhApEVBCqccdCJh8jhMd7+v3n8VkVXOAWsq3huJ0
oAFjmGaW3BdAFwdVnQSskTgVKLv8PHHXfv1Ec5lcLwkM0Wpx920YtcICUpJR+d0w
/cYjpD9V/zmbc606ugR1tsZAaudpzgXxwmHjR0xEixlgI2BIZShf/ssWcQWudYbY
RV/pmKIGPoeMhvTw3QDIDzTESqXPlrNfQvqgYAMl5WKx4PM3/31AVQCYdAkJudSx
EhmcvlGX76Qg8UBz7zXD1x/pjLuO6smEYpxH1RxRLb+n7z6doihwGPTAYXIlXSYZ
8e3I5672kR6yRMkSldbQNsYsPEqBUJ57S4ac3rzdv8ryy7CAOQwNH5CbpmvgnOMU
C+rx699po7wZrNcoeQcz30wphUgjZk5Lxk0PMkMHswRYGsdTVdOTyR0Ln0kFpyVw
pD6c68Nb/G/8OOiUPAv3TCKlAG5FdhUltu/5cExoPuSleG00gbbEQefpEqvcAvEH
7GJ1fIIOknMvf+7ix1S3veSGs48Yfrfar+QsCCqFGzQafpndDZz0aMsy/bcFAEHL
012lijO30vfu2tKSo+FWpXqMwb9ZFK3/e4cZIuV0YfW01LlwsQIWyWL3oAF782ha
N7bnOfzXKWQp16EJuyFuPwEODhS+GtHOAq++HI1DAEADqkw8tuPlApPPvCQlrx33
/K3VZ94kG8un/7DjkStZWrk9fryrIRG4b8JLhwx8kPLc8JGOUkiheehxL+Tyw8Xn
C6HkSehuwzNc4QoIrhNognk1AEiXp6Gf7DA/YZ6AvwlHk0bgg7qSa5Tc1Fhcbcg4
vM0yVYm0FFJnolfGgQPEpjEjItmkGEI6HbG82ZweZDA0/4RP2fjOkOovRg8Q6NMf
MFadfNjw/dHO8P32ISPCUyGQXnagnxta1Oyt0pUgnrkg07p9t5KvJ7R2Ldc+bdaF
FreU/5k93RdD6zsViKJsPQAKTlP2SYKR6gi02Baoii3QKxJi5sEnOPfqdS0FlC4r
6KQiTrS7IZSYYs7Hc2Vle6ewtu51ZaXkr53BUreEdQlZz7MV1pgPtyVAI2laUp32
rklYZ3AvEkWfZ0f+6l3aQatksFs97WaCmwyMwJHOsqbLVlh6actvSZReq24G8luH
w6T6Ssl5JE/r1aqG0/2GsSF7xjQ62zlShay3ia03SyprsF+3YtK79OcmUEopyrwL
mfGG/SZrv2dqGtBfXJ9wANSTaedM5mpBdVOBvJy8i7eaIQeImE0NutRvs4LIb1Tr
TXTOHxyYf0acACMB8OaqGrCVwJjjsmDRcg/wdvzG95irsA4qBofGcBP9l9bJX4+Y
Uho0nAIwc8Q39/9Z+nWIxBE8Fh+eGqk03f2zikXu7HfIc0pZNWbuVRMGiB4A2MZ4
Cbyn8z572iSawXPjx0pf0iJLT0AFOQEkYRYP87fMnBz2m/5kMS4949GDd2UhPvJY
V2p1iFBqHZUq90YoY6CxZR6rHm42WUWDS82fjCklBDuIvfdYutKSgZB9rM7MJWHB
yOcI1w/j0k4aBqyCvTugfKurUXe9SWgt8+C0ROas6i3Gl+PAGThxbkcjp5i9OkaA
uYTQIPrx7mWrvA+RafhPKERiEGSEuxKdA042wbI7mVZQImy8Te8Z9zTa86JpqoNy
zia8TgxvELBDfL2I3EBSL2wbhXCo3nsvrF5HJEKluTtzwGsWFT4Hw4V94UE91a/l
XbfVlveCDDcmbFPilZDXnmscl/GqUFshjm2IGW49frWy5EKT0UQznnhjzvi0fV4A
2O1yH2ak3ClfpTASFsXM5S9L0/rZgq4JLL57vwtArAnErdcSzjb40421MMFmiwmd
MkrwdQaOgnfu5WzHaj3uThiv0l+iCh3WTd7OQBZWRMb1ITAXZrIVXJnzgP3HP29F
LJNZhVUoK2ahI59M/1/1tGp876xyz2OseZpUBraLzgHe0oQtzjn9oam1HiaXnecU
av6UUKMjw4JHwDflNmr5GHTmuSo7dHX08OCcpQ/MBu9YCYsgWOEwAI3v2VOyOQmt
XqsAZGt+UJ/brAHd910fyLJVE3SKzr7S+Q1DVXbS/AlKbHjiMLKHBJT4YWJ3ZtHV
CDbm63MLmBd2kQuQRGMJh1T8LuRTDzvuVrJSGMS5fR7oUCZOx7RlTsQUXAuM6WnO
uYHDyGjjf+yHfLnbh3jM2y+MWwjs/VK2fmmFIyThLZgKtWHE2Xt0eXQ+0QBIQ2To
2OcPMXdUOQQG70FRC4OPrs59XlwwssZeamaluMqST+mnZ6iBMRXzE9DEkiL9dU46
SmtYPwcIZPd5ec67oWg/RJP8Ce1kKbmheaiHY/pva0oUtgt3vfNcQJmCvDUxOG2k
qKZQHvtuRiSpkqpA8hxQMdvRs0264QqL90kT2pXQhpGJCm1FeTe6CXoQPNG/meDP
/85PJLwBrv2w2D6tDjlb5y8SWUUoCYL+77PmTWa4pCrV20xRlxhZJcZykoBag4So
3G1N8CGfGi5TgsoJNEToJckI+hGOsYhSww4WZ0iHem5Wbf6/43P/ZuXvCsewC8hY
uCw2vndxo/GxiFGCMqfubTVll2d9NxzOOl4KMzJhtahqWDoGW5InIqVxcI1cOYAF
vDddZkXRNEBLf2qtR4STJtm2Hmk5r0d9jJOTy1KI5nbBPzAcKs/aIQCoHVl2T5bh
b6sULu9fxruRyylCaaJfY+wP4TkMFxRyZoLlKWLYDMNLqX42UiBWcI8uS4movbtN
3kQ956cLd1Hkk8UaYXjZywMqVWbcB1l7AHaFVdxkje1vodCr4CkIGmFv11XECzGs
SNOKT0SRYdcHcbD0W050YsWuuDoSyZ7WoE4j7QEDiaYYY84FAyOVrzro3o2TyBBr
cXQ7MX8pdesD1ryGqZXXfN55O7vPM8B01oC6JZBpR8UZpt4ZULr4VtZ4bcmovpvD
YkUx9/lf6d8MZc1up5vJOJmWKw3i/px0cljslaFGYg+5TLGerEI6UiDqFWI6rmNC
C0vIq19snE2gCug4H356HMDhaJSk/Ri0cIJaaQPF6t/3Z5lMKI4elUUnnVKyQI7G
zlIhKBvcj4jQ4Fr1rygddCW4kRErD+Tvd9nBsRhLEdJzYnf1Sl8WVac6nVKi6v95
3UrLViufYP5/HCyGvjvXsi7vpxyv81a0zyu+FgkDiZ6seS5pszRs1b0uKgINyrVQ
GianQ1Irma1v/s995t9GOMxUhgrlhnF53Whce4Z0tdMxXFoSFJjBdrCRjyrOfRHi
645K+xZWCPLYu8HBSHzugieFMurGkNPmzIt/RCqSeHEOzsi/yCDDBAAaxJJLQmFX
n0dl5/ms5CWluYFx49ot3ukTx+cVkFwZZ5ydCd3T16lNki9733N+17uv4r2zKXwE
PYx2aONJHnwnxBLP9QjErFN+ySbncwoah/+tYnXXnr/xydlb0Tbae6EGHoJXBytp
xEH1dCRSgPUl89z3fxlE2L9YtjcfoxmxF4ilklv7eswx5aHmQDC6YjvdgtG6V7p9
6OpFM9VW5HSqLV8+aj9+/77anN3n4wYClH0nIiE+G54IoPw8AvSN9XWFK8WDflN2
ssCzgc4jS2NzBFAiM7ChjHfmeTIRZM2zQZEQHcP9NdNPeTXiubqbM2GNJraTegvu
VsnP4zvulpMADMNlnC8QmfjqS3O/58mPZgWZavb2hUwPW2QU9bAmnB/SdYFqDMyj
ryK33Z4YvoYquRPBVISn/4fcspezGwCNCmG2WZGA5JLmSygdzlyPII7cMepMcjWD
3slrYuwg7NFcON6Y1iEHLlXAlTD8a9lyxtmrW3GrOHHVdFu/b9saYs0D41y7vG+Y
f8PeDhWzAy7DmjKHc/0bDVfMb+R9NWkW4uXVr6E5mH8tSGEEPHOI6Fw2hzk90//Q
soC6X4KUwTV36r/z7z/md71N/3ojg40wxqXunZjwcKKUZePkLMCRA1m8Nvi1jW1U
gmCjDK3H8gHQati/2JJWUuE7kG9tFWSwyOEJHfa4F0ExGlTM8wpJzGLC4FEoBr4v
JeBBnqL6SbdDrH6sLc5tHCU6/N3ZjabmVTrnRySGnWup2ThatvI3x2kjtEJNk2eF
W5wbwuXyXXZuLj6y0tDVHTCgz4ojK+i/5PZvtOFwomQWywMkJtdDpBUTUNw65v5O
Vy9cE882s46zLPE2iIJMyx06O0A3ZBkZq+oDNIBNe6eqIdMd+keVI9GqPJ2g+wUH
wzlBaiS2EQKHA0i/NmReQssSxKXCox/qbhaotbFJudxKqH6E/qqbyVFH8RQybDQf
0ppv8DSnifagCpqkmAB4fzzuc5tkAukdM7zKOLp39t6+Nu2Z1eisdGORpjqSpO8m
IFnH4gd+JO4SAopH17KN9xlu3Nfc4H+1X7WdjgmEuWN06WbN9BC4CBQrnVqdIoo/
as0AbRQtDqdGpPjt3MwQxwATOV+iVKKrPcX6QkDND9Qn6rquxGzjdbE2cfx/7OhM
yf7zJvrUeKgmql63+cN8AosamkzBIzqe9Wp0I98OqPU/7BwTzDcweTI+ADilE0X7
wYoMgSQGlY/Yx4nVCm4QbqptzsdJH/fo0qjkUVM8/Q5DJpekY0zIL32LdjaqF0O3
0b4giFoJS23Jg1xQE5HLwf23QcE5uR/Bjz9h+TawsBqVRia7RgR2aI2JtATxkHQw
Vea3IC1FX4mXsQoOFv/TcmLV72oSB0t2uc3iNuzl10oapKIi4RJeohOJGmtcLp0H
sn8e5GzVnpiAz00GbCt5WE3QpyhDada/EDisKeqBr3dMCOGwvLG9mP61+nNJ0v/g
LjrqaKys9gOd9JkZlO+CSjtQBSIXs+AV3ubeIQcMzC/9YzTymKUnQbou2adlLY2I
WYAZZ4SKz5qqdyzU+g3Tr3xVbRYhaTG110Jel2QyYgRTwVyMLgr3VNwoop+ktcXy
1YJZFHM47TK8a8B9W8rzAjldt2o2fymaPmwhvcW97FhLCzMYetk3jTfYxNt5gtc4
fjiMfOh3tcQ5dLa8sm5KBczbWzvMZI/7RWUtQFGqdq0C6buMVT97/hryoVepNF3y
KOaHdH0OXrXkLivqudRJzj2GMmT7OG+QHAIGcmDZ/cwLL9H8tUTGvQMjZk9KOKk9
zAZn7lidCTafeMfneu7jKpprr32Z3a8B6MMR1RhGX2jnffgy9FDtrBTEKJkQoEUf
h9xCnP1I+RAYd+PqkI6UeHuwxFxGaig8j6BcHBi28YqYO9pL9dI1LhSFCP+i1rrq
YDl2u48xsv5R5hlrj8RJeMA/f3ZM63n70lf2Ml5oW4TUauLVZvRcZb0HGBvV6bzJ
++zRTp88vJzT+WlV2AX0ddtQ8XaebXyOV9NRPIy2RfZ3ETa95tyJt9VQRictQjeN
WAoClZiljCFmnSig4zlOuqe0ctor9gBOzye0wY7THcKvY+hhEzGJ5ibZ47R8wVaS
gecVvqY56hx9BsQe/8MiQd/K9lMLMNhZkmS/JCVNvBfkqK+uZglq9o25yni6a2IZ
p7+SDMehLzRbEpLgD2y3T9z/wnxAlSLXm3hFBJ/Itj2U8r0RI9L4ZqEi7jVNE0ri
i/vKDQZc9Ypxgr9aZu3/lhnrvrjjtk+5mdgxD7ttkWAJBwMBiddBsW1efn7TmDhV
ESO+yyqp8IgCMrulNqeAw3dYgByPnuIuRmHMroRpXV/y5WmwOjGk2UsDUjGQUzGL
dNvDOtuznEiJioV0Othg6nfkIAHu4jabMbKraoLtVFnnGxj5Jc2zrSpKapnzyy+u
T7FrXyEBPCtjeaEUA82VncJl4Q/Qj5C0eK2w29YR/cNiLwd4uFup1mIjEkSIz+Na
orym3PFYrqmv50MDsy6bfgJlqbs+6oeXyYb7MQztj8zydgXjp9FFdOffBmfkBEUW
n1gFzVcA9n3dNR95hnekp/OLNsubuci6QeF5AmbX2nIJ5RteD5sJwpdHo4kzVy/w
JPHx1Z/ILoYiOGJNbcJZ+R2v9qCPUFVVrj4X5X3F8D7T7Rkds8YYZXO5HP57O80V
8UdB5c0O91fEA79RPEKqpzf/YwzMxBH91Ootpd2SlDCVAK4Ea24rarW15kEC1ADG
BCwQxj/jWM6XZAtLX4UjGZE50OrCOWNBx7rZ+D9oPLDjQTRQVp234hu9KYx5Thin
E+ol+DfDR47s1L415uX25Ocm7xaEmSHvf2xMwa/MiIh92dgKXCinW/c88+8BUbaB
87N2cCzSVUs2/REf2HNaLGItlKoNzOAyVVe2yN0A0G4OGVCukENcu+1S6mbJgkpe
ucmx24H9Mv/s25Te3/66iKj6z1at1XLPHp0Slf6fSz7oKJ+Hius68wphwhBRHwSx
v5mjBA7FA9W6GgG5uzwadON/EHuivh4Qtck4W+1U6S2nQ2c4mH5OZT4x+eenzGMg
mTwTga6g7NySrC5fikbi2Mnga5oxobucvYhvMP5DGHW2Z+19UmyRRx0TsKV8m7CR
WXI3/WA1Oeg2q9wR7FBV1jge+ZdLbl0ojN/bawhKEN6t40p9Swn9XvKREsz7+TIf
l78VkH5KkGfmQn8rAnbrUhr/93yqUip+QmPrn5wUeg7uxvNaU0rgtWu3V0RaR2DA
3HCDtnChPhULLw6bq56+hOcKt2EYJznrIAgYsdhAnQo+g5yfKM+HLJngHkiufAqW
Ufpcuko7FGN3NUdNtJHvBhh0TiJ7OChCgLP1AeeQ1gDppVUf+y1tV1sO/yPt2ACE
f3Uj2oCr2cXlB8jcS2k+yd6sDB3EkvZ/eVGd9OrUFVzsmv5RlAJKyzaSAf0Bfeba
T6S7cYtpah+6FtjqttjWb1wOik/Db1r/18QlxOhF11VTfac7xml+IuikVfFFlBWH
4TW4wrVUesYplrm2ilkCSszT1C/XmcnsyZBBCBvrEdy7Nf/jpQ0M8hhO49yxgAkn
OWGSBL2V9ZdiC8ocRQjprUekCNL1Gr05blyAHANxaKi49MNpZKstKhx54LoAvbkm
bfl/65mftpr3tpn2N18r0wPwkxGg/EP6xKlys5KZd8jUTDEwFZvnQU4LxfuX8W5A
nOHAHDsoOjpZ0XaVoBZKW0/lpW/NgVw6HiUFaLZ83AkEuMQRZoQJj3Rm9z3X+d4g
I6v/XGf2sxeHqeOVtnl3aFpyUZdkeHv2/m/1jxJdcjn4+lHtVSH7yIfu9oIiXAbP
A9zPjBMRXuRKqfWyafvrhGtupaJWXnP1yjtk+EY8l0q8zOgyM7GyIqsRyU9Ylkdk
xVBW6CGvB0k+7JFZv3HsyNHZn7WWzOJVtr85hm+jio63uj6tSKepCMtdssLAhTXT
/M+4OkplD8TVCrSb7C6CVrO6t6j1hpgGPVmIdjyaAAp0foh4EkSht7mT3lc/Crhz
fGZzLWMJM0257+CDqgcVUNeWlS6hPUzL38cij8/wtfqvKDaSACTUpufKp7AVwOpY
i4u78rcM5hxGtnAejS1RJjCcoyNwgkzWdeiaTgmeZbQP2SAhvnPfVHS0fR9mDrIJ
N1TvVRG0wIgFUssnFG5p9N2Bt95aOBltgeB9A2BzAAy2dJI+RaThZC2qMxE8ndE6
xs3JNvhcIkT3XbYx2eS4gYQeK0s+Vntmm90u3UbZr6toZ7pDIrEc22vYK59GogJg
Frg7y6tcwMaorjAq7L3J791MQBSyFkV0FJSeT39Tm+JLeLz06UYLMp+TANADufPp
lEmBYeCYCtp97VWw1Iq9p2aSEH36d8teCc/HaeOwGsekEpCzeziyqVSQP92CJs2D
IF91kKsNndkUVnhGZ/VXowVTKzzMcuHQPki5RH+wZgb1Kburdi7S4MtDmgrzs/yB
eOYCexYVvipI8DHfDA+J6O6SFiLIxe22m29GWgXz3867rpBnXpNW4NdCvNciidEK
MgGRdreZYbjLcchdgEYjrp6fQxcjbMPu9v+CfAtO5sSDpIvc9+IWWYSo6w8RNniI
k/izLy+V+YAE+rR4bf0d6OZTFzLJxwRLNsp7yPdKVuCOHTaj69VIr31xXKUb0/G3
h6MA/zbm2WqV0R/PaDpBW1Di/vUAc/63yTNdWn92C6tXTfSPnKAlhBiGEeHag/Sz
lDADR4I+wLFFKpwBALTKvHpEDWfRWdwmTPs93ulKSSaS7jtlu/5Vk1jMoYJUZOeN
xSWc0qPicRw/Qw6X6C0JomNbsdOAfuCXQScV7wrIiXRGHMOw7U46fhEPPY53aNr5
eW9fNkQLm6KRsOhfIzopicWElu84bOLRPGg0HBbLCAfP4CVIF4ImjHdWc0rdA3eZ
jJ+y10P5u3xXjmdhr9oNE5yzw6aKsyVYBhs7ROj7lEwmTpYKn+01f/eHkqsliag9
2EEl4SFyMMbUNroYPOAXCFHn7kTr8AqGdBY0zzJL7OmS0sZzOtrQDOhoVMlIFW4V
2y5yc+tiepPv8qpHaPkElO7yCAJaagRjoxlm2gdXMjiO+E5/GPAcuqgRWUrvtLA/
m1bu3q2NOZX7bsoq3Ccr/UYtiXpNAw+FhB/R4xiDT8/eIe7RNASoZKEifC/o0idr
2vvi5yV85n9l8KOjQTbhGiJ0gEgJGBMOGpim+G89v+pLNK9ho/UVKomrvF9qMkWk
gFLlJIIik70EE056TahwkSRIva42cr/xsLXUPq/ZA1Iz5VXRymmsaYi1Q19GS5hW
c8M+mIO/8k3chTxodWdXvm6fZGJerwI9G9NrTzUuPcRt2j6EqiYSoC2tHgRYexbR
Rb8zFk6hXYXq9tEeLKDIvZIL+DBWGPr7BxDx/gOxdijtgIycX6qM4N5rMRQ1ci+D
Y3TXsgXwhOTqZKmRZqKC54IdMSkUC0ldakQewYANcRK6Yr/V1d0of8PaOAzKE+vN
bS9UViLrRtx9Pabh8ezSDH100o7QuDA6D3Blvp8lT+LTY07mOrlH75M8u7qfOVQ3
KKYKLVTMzWSYsbnnUexc2CulMNyVmWyrygmHk2Pes5OAtAYA5hYxhbFYRt7ieb1i
UxKX21qSDTjogIKWAB8ktpaLMEPTt2hxt5z1rTV/CH044hXFXiQSJNEObe0/lmuA
dm9LxaB6AzyncWfcZ8K6wCHQd2cD/iO3vEAqvP3eVgOOr6IxDOLLGlE6z9iDPPII
7OFNGdUUsyt9f3LUeY5ihaEcWHe+ip/MCDQxGArht6RPUjwkH7QgA28FS7pS3/PC
XzgrvQRuxFLA7nz1Ji8IvlPcSDgALCccrcjKJXYDYrM+HZAIbaD2lwX2bXyXStN9
7xvmEQnfhgGllaaSRUCzngFzuXMMrZ1wHYEYcTHGgdd//y0rzFtMoCInQh8w1HrV
VGNuDxxEDZ+TX8eihdTNg4zG6aY36zWNwZt1GOB7HA+HFUhmXxdozwWnpnSVvstC
E1ALoOz3LVnfEfcHbHX/oUEeULrqR9DlJIr+CkuvWeAGPDzr3PV/37FxdBkPQgE5
1TUvkKWubS/vaDfr/M3nZvOis+KngQ1vpuG6v/PY37R52O49v7t950GVAsMiYZpQ
0HEBLZzvmzSraXa8CfTLWUDvQH0uvFMrawE65JxHbdjo/tCOG5AIuRuxGhydWiqx
bq2C+UrcyUHKJ8lrO2BodwyB6a2uiLH7fODStab9+Hx4WNGkZm7Nn+pvTyNbu00Q
wRHiLvPtBaxzQJtPJSZUx8J3ScyTBXHiv8u9wEcgcHNJ6zGlz9VpnvNKQT2gUpHr
TtFifiaZOqTqSrLFfevxO0V9E1fDaKXCYrJaQCvfIsq5DfAlTmb1k9Kvdz24BK1B
73IwrIin6FmaFbrQlzz635QowgptZV+YdkkK7GltZAdE/aPgKZ6UR6kGF7++tGbp
cSIomiBHUvVlumkG3CIDSOez/gr832+cMI3fk/L6gjktR0tFsoFkKy3m8LQPaIAq
kJhAzMIRYOjaYcNd1Wb1FzAuG1OIwiv6Eaf+OfzlHvRg4QYoIQ4iO0tkhQdIb286
tWn1Kdy4RA62M2NYp43QWV2IFwI4cCszwseUWOB/npwEhO8Ufh5SGp7h5Tdle0Gr
M+O6FG2b8mhxuHLBJeBEXHDILO8jwoLJ1TnAcE7I3nls9c6/8rjPLYsX+rMWLTE0
WG8w7mk3Qj/KCGCER4oeu11SoY3A8rsTuYXCTOhgXThIJ8q+9l3+zwwbUiDlxYpR
ChvJSdjXL34SwSs6MlfrKV32cvmYJhSxPqBWK0x1Ueppama5r1YGckn8JqIoDp8F
+z+2dVW94VlDGfNBpchDxbIpIoLO1COaPa3NSUTOwKhWdLSqqNldkbQ6xoTfRVu+
yRAjCJ/tNM1nxHGaZLD2ysmh7cp0vS4KdwQVvkNstfAez6i2YK4vdY/uAO8JTV1L
xQUoLWDndV2Ab8G2VvPLWJuats/nccPYjpmCsMPeTdf46xL7Bx7MsdVO5uCba8cO
n/SQdeJNN48KIj66NeM3KnHXxE3YQaR3wgg6+BWAY2/CqzyiJI0OaVN5QPgP4pG7
tcvRUmGKj+i1PhlCIKKHrRe3W3ei6iN69o1f1l0S4ujiGEmI+cgz5HdCWsOKkYlo
F3K3gDwWp2Av3UcJrBRBTdtTxN/vGlkjeYjvgS0rEfoAMebeUbRav84Ikr5+BeRQ
iNUpZSlV7/hJvKhNboeGPjinvokuO5De5HuB+39vGXoCmlVeGKsgkwjCB1P4LmKX
iuzn1iZBA9A09FjS8rBnLe7sp06AaAE4Nu0bceIQfGdaclQjpgKB8SrJI6ENrjLy
0elDXR8f+kCSKtxFqZ3rvq6QUetKsqfxZP0kf+OXWvZdtsMoEoS8p7SAHgYVzjSB
eunGs0N4J/r8qWaiByT73Il/TX0hlwU4pncKn6X13HJ6TlaPczcDR8Hzl7jf8RGK
ywhhUYVrFZAfhY6Sl9wYgEzynzecqUkTJnZ9AGmZDt7QI9W9BYyG5hcWqV0avqOo
n1eaUr21PFTEf/tD4r7APpwD03tqIOoA4LxKzh6jhFFglae+b+C9BF8TMERZZyUl
ndbuKvXjVMXmKIArvw6IOLZ+9xUicYNrAhpUD9p1ky62YUEXipTdRIlpiXrLphwY
UVYh3qFIZIto+6IWTf4DQeUi9EBBC+Wu9x/RpmXksxGBYwyUVuTMWOQQXwOeviXz
HgNBvAap+oD00AmB/K+AHVOafteTYry7kOD2rMSQJkY8mELZgiOMioUN1CU8J863
uKQqaTvBq4vQZsHlAPS57xlf0g6GHzUb3/r2hb6DKgANsB0sieqFy9tPiCJU0tfG
LR9E8/jE5IQtD+zFy0J+4ndohGigtee4vZfv5/m4OgQ3SOsfR6BGxVhoZ18UOBjb
tfaDEQEGplLA3gYCA3gqqMXaLAJLP28NKlII5NAeu3L+hzhxsqFM50GH8GKed5c4
AITUB/mlvuOqUVZg76hBRR1T8kQ7EQfH8cYfFl7hs61Clum05E7T3gn1AJEX/dQM
PLs9PsweVYzAggsJzx3IeYr+il8VDyau3dz7seZ0D4g5KrKsfOOdAwRHC/5+dfcN
oJ4pvduod+YOWZfV+DC3hDO6qPqIlHwihK2RpcbT9buWM9tawnRJrsMsXqHr+DOa
V2Layp4euwSIjVy9wDHIAQjfFZiKAn3zOJAtdEw2UeRQHY9ecT7ZWknG5lUUjYnl
2RN/R4AfNCYAcI4gj2tdvEvFA/A6Ic9e5Co1uTveU7AphZnVOoY56R4uQcEDgsun
sBljYNUjrJV2n/gLCUbgkQ2bN75bw0IbIEYllY0p025ciHvMFnWXwcvFikgVqN7l
vF2Y2+CoQ06g2mHZ5ChfrCEkTBUIZwDaHn2GSusWubVpruLuM48Q875bHh6V4Y5y
fKOw1ZiVyiALOKUq56b79YlcAyZXvGo6xsVahobWPEQINcmKjLB6CmtmwtkEgPeI
ySGENChgqIhw5Ny0ycuVOqOb6St6jdCvYm/lC+7xClNLpbG71c4PvxvQiX283VNX
y8AFQtFaMIGpBbAXQmLoJOkab89ZObJaXHOOp7AE2Y+g8gksciCKm6OyY9wRC17a
Tl5Cwa5YDcintRwtqBtHmitafWyPY/i+Uw900msT3uM+k/LO8HKH5XioqjSF+IN1
ma6CWErBc45Y/Ce4S3Y4V/R4sYnTTcaiLneDIFxDcAVU+/Qbf+7lG9oijzDGMCti
hsUMsfvX1CdRM8lP9jYY0cHPAs7uyJoLdAIztfy+70T2oWIyTlpx5Tzecb2SZpDL
Zyw99GL5zl24CyPER4XZFk2SR3PEWC9W8yMHDfm50CO5Cfyn482fHxir1/7APMXw
Edy+R/bqiZDct5Kxdnc6GfiiBQHnDCgZ6U0NiHZFFGLahURyvAvTBr58SUBymrXo
jkksurQFDI3dg8DwmkmM4kGvBhDwKgHXQk0gL3IwHs547tehlvN3F5pyQj3GQSli
U3jClymfDYT1SVZ+PUk3Bpu4Q+r0FaPg6vAwHaM7tOGNtfqv5cITGJAQgH5CKclZ
TZzJypeEgHjKGRK6rp5ssc9YGO9wBIe5c3udI1FVck22xxGQ4lvLZV7zV9b+IY59
jAm3Qi8Wjl2zC4x1SrUN+nxlFnWyvFxth6hzhRMOeNmRH+WhzXfYByUN2+hyBGCF
2FNHoQCm+6i99rjESlNBhfusLTNVQonaggM0Q56c/LNyilSvtB5Mr9B8Rw5XMa7Z
9L30wmHayyuUhnZKUdtkgU8zphZBVMfbw7R1fjdwkHcIiA56E7yLRjxpDU6yx3eY
7mr2kG+IDUcdJWtQn1IcUSPt/br/pZMMMb5o9kD6UKkyQhefgn+vx2Ae30sK9tVI
tGqLlaEnA+UZg8L7BOX6jJPhdw1SJOzkjzOnSK2rMksg06VjL981jdSOWascOtpD
6wBwnRhCww9r6lyjOVUWXN6WX1nrzYzSc+PoXi+R1HCXxRv2YWGuYAS2A+Y/F82q
NJh3ElyZK1HihR4Ltd4VmRI038JqoXWMi7em9YIscf9479l3Tr13ZmjOAFke+vuc
f9WJXFdf0QlXWDHH4n83QQMhtevbSImB5SaVsnzAgXL5vIp08oksX8FH8Y+/3HS7
DPRuOzECDhTiJyCaNSQMEhAH86quIRDdLACUI+p0z5n16Sw0r+4w9RGAx0MHho4X
RIdN3mF4hjXKVE0mwR2CZnCHOtQi8TSQ2m1+zAA8Fg3ujKtVAQaks9zS+c9jWzjk
fYTT+CDkIuUvJcZkrKG+NoXOFmMyA+wOFWbsLkaWZWLdSQdb+TmXcDAlcUsLVbyD
vyyQ9k/QtCJf9iFhJo+hUI0hALwgymaIpQx6oL0luKqqZVKVF0KUnEg6PP3yiDh9
G7yEFmmfMI2XkFG5r8zHctcuN0uVh9t1FBezRTfKnyOeGs2T75IZ2BhWezrOxyQi
moEd45Bt9VMW7/PtoD7JiUh96T+NJj5vraPlLFdyPZxzRnFPMdeR3cQwQ5XjMlg1
UItoq/VOp4tnLsSv4MLVaqoToHKnk3lMoRrQ6r85W+a79scv6qHzWZTdOEqaxdEp
e2dkBXqtyzjzU4QyYSfph90HCFiQr64OtMbMd3awRMerVrz99cGXfO+TVz1ulnh5
s+6yZKVZsAmzqV1Owfn4NLhiQg+dZHgnwcY7u0L48vdJKxzNwr5wZtWk51I6lDiO
cON5JQfcyGI7SeKBY5oYMLduGs3RXbv2e3UuWvIqK920w21aaaLANTdkXDPg+z5k
slTueU0gvsprr5zmbI1njFigxwKAcJlPaRa9ga79NRmQxCK74byOJUMaHRyyeay6
njAOsVDQBLFSgBZ+EgSmumopSJpPswsnS5hpmH0feZ/9sZ/g4yATaTp5zy7p9Zsb
Bdbs6BxdDyi6YHChEsTGIy3hvTkCZQZLOk7C11RrfsLiMiVLzW+rqW6czW4U1OTg
PPNlEx2ipfwTb4hJUXxcp1X88KXW2i1SAHPgg9h45WhxUsNCLfaNjohoSJ04ROBq
oKBg7oQfZSSXR4QmSdVcqGeGwxe+0f6VYAuoTLiYkocDpJwRZsgOIcCVFsIBJUWk
1+7MVZzpYhVu1caSBFkfst6VMWjuQjuNoc76uQ4N5wpEhYD2wRJVwwJPMxd51HrK
re2TGUpQOGly9dqcQt4Bxkyp/YJHAFPkQor2SElkVtKEUXiyQ1QSmlh/nekpXvd8
oVLFhoViyF7x7VX8nIzlbO4rqTc9QujtIMwDAnCIBltWLSfX/Is9QI+aRfbkqG9N
GXslo//cECjviTUoQyLmNtQe65YcgFh/fN9p0jRB7/xgx48ut4vxFgaykJAiMlg+
wnYjhc3iCT2PhMZe/xuzWM8UvVr0VqRbpLIcqQ0NOwRQmL5VW/5ZqsGw7zRBrw3k
jTgLmhbBxpw7BpTfv5cmsyMbatCP5fk+q488ZkEPmUdULm3SSSc2lTQpoP1n8zoy
7wpkmZOypc1GCuoWBA1sqgt8rGDB3br/W86ukKJ4o1QznXuUYurVyPbwDhQKHsTU
zvgNDiEVk6Gr5qZoHk7eWr5vEriwKVp5rluVoNOY4Rp1BQ3w99Xiy4Rq3mQaXshF
7EKF8He82Bbl34hkAZXTeODnpWlG3nQA3aL62t6wDa38v7MrcLUMw89xWIgI4E7j
wfCTSsbrXnQ0D1gWNb4jLUX4qNoVutvdbLvt138E7sXAqyMPYpdUsSWad0nv4biO
LtSV7snuskq6R39y5D8rvzU4gENeQuhjRIftfKPUkIV+96bEkGAicepfKKslx8kZ
gbAv86IhlJ1bnKmmZ/i+QvuLmfQ8zU88Xxi/hqREECQT2LRMT9H6lapMW37tgXwp
LP4/c4NQJc6kFSQcglbEnuGU4091aiq5rUnZFd1kIVXGbrinzTBLbDZ1gFp+d2io
Aavq7KOwRN+vHDEXMZfppr7XL5DwHamIcvTOFlwtwBfqRc2aaRUmiIKEDXIZ4hIi
6n+LM2uq2a9Smp9+G5B1YrzvEFBG4hedJQXy7nSvZeWUnOtKppDL0KTF00HRFVEP
tR7i7PzssOz13uM2/ybKGzxRxPWvQ0sSa0P2TlTcyNtUyow1P9lxNdXqcacVVckZ
MVmKB51vduUphz7HnuAMtsZZlYzfCNuwJdtzGRxPO6snDxg8hm+oO+m/DVNLVqxY
QBnVDCN/t3oFlV2Wk9pug9C+5gDTqWvDQRkJXF9YqiULn/A0/JwXt+fdwCcAfUUy
67T7F1VlYKbMEJbSfNJsT5cvb5MneMnWcsl+x1xqgO+Hf9J6/wrBVN64ptexF2CA
M8cYhipPm9Gt/8FULAgUf/Ao0zzftBPcuyZGiGl24Y9r0FyfwhLqhHxLP88QaG1R
j+LVB2bNDuuDhzCHiXr0LfXqAai1Sq0lpdXva3nSeBZt0mCXw4HceFG3Pt4vc3oW
K+zyvT1dxJE2KTrBBgMKfwQW2nLMvRInTTlOeOrNy8HmaYFsANj7GMpp42ZFxOxq
ahsK7ADbK/S3VN2iSZazPcSCPAUPN7Pdsjw5Lb9K4xTTjaH1L13Tnd6cBcW7S3/v
jasKq3O8rA1cq8DtRayld+Jrkgo+a7rDMeJitjChHMSrDd+mJrK6acllDOL2FUlM
5gbDG+UGWHBjQ6Xc2MK2JeYZSt8z04BYbbXzebXIbJXqFlkmNTjYKrC8/xz8HlLl
v6M4luTersJEmYcD+k1aLjA1i/mGCND0pMe0KlE8onBtZCzJ3l/+eV159iXPhePN
CBLCJq+ce1gh3RjmVdf4upw74RLgeDV8ScbMW5OkiQ11V+w+23iGiUHrmPlyP7Lg
cHgIV+e9ecj10PBYokVyHQUuaxZtfLhc9U0LKad8DckUTHldqOARYaSmagSkZFtu
8AkjElm6z2ZYCEDkhmzwVQgrb5XfOBd1da7JfyDibpbXKxECrVEUHlL5IkY5ob6s
+VxhuZ9g+inbFQdoaLHm91GUdjIbtcIlKHc14iiAGFUajJr84e1W2zN/jzCvj0+a
dj5hDQv+NIu2DGhy2fpliuK6Xra4Fvn3wtM5HUFJz9CzicCgjedgHfS1dn6l2zlb
6K/0Id9eRXTbIpqPhvhU26bbUtQEeZgnUa675MZjt0cbboVBQRJ5v1Y7PDQFg1tn
SSi21iBj2zReaZWwM4KX5BdKgyuPdTpTs5rM37HlJQFSBnk+2geNsB37xiaehnUd
Qq6+ovUim2oHHjYBZFp694dtgBfNPYMML86FI1Jk40crs8P9G14edff0fsB/MVvA
HQaOIC3OLgFA1uZx9oGatMbt+rsVZqItWVtZqFJg+++4aOx38Jmqdc9cjuFJoGLm
bSkx1hEBTxGnVEb1Nj3hkD1gN0cxyYxXtogQWyygKMRnuDv8Bg84XNJ1xnsuP8iQ
kGN5Vbw/a02ykV7/aRU/zUgnsa3ryTHbZixG/QadcL2Ee5iH8gntUA2ShD38nPKq
Nvqv088GCQc37a4+ZF7JTuaNZNzMfbzOdxb6Xlvq/ZUzu39g1YKJt/JqkV5w9IHY
MGj31PvoUz2hfLHeVVqFHDB2Ifg6LahUiyWDfEHUxTxHIi7NkBaSajgMc+a8Hvxz
55svR8QaPzATsBIVEh2M45urbXAI519LinWfbihhzPm/8CLzQ3T7oqvMQWi36uw7
klYBwMgU2aneoAxpUgHhXerTXtl6hfgpbUn1wT86fvoko02TbLRhFGIj3gh6N0OP
FOSMAw3NrDveHu5VTigCEZmHUgTML6Ai78hWWHw7RwtKTXpPeu2mVYrVg/sr5a5W
cRybV1qnAlqYOTIku3tI9ScOPtVqjpgZBmXmadhC9XvYYIYunUzzHndlCnldFpjf
fejef2H1t0l+IpS2lavie5ENxRY4Bs4vXPcYC4/yA4ISZ0x22LrVh3S5ec1xFiC4
sVmlekpGa/rWpf93D9PXZfmQtRH40w5NmQ1d7A/0ltwI6bKzTZUcm8qEsKhJPIpS
v3y/q9BHI/Zra36wcKUWWKQBywGKcrnENSZ18TI25IUVYbYtelp/H54QGn6MpcFD
1nTt1jDuW0cghQU39IFcWvPaMgr0MtJ9ss0w96KKY4s4CZg5yH+6ibEEf+IFeLFB
PLz3wmyyKPiKvAdiEzBoGjb9cHzDs6XPuo8zL7TCGbz64USFgB/1IVuewCduxxol
Svo8T514Lm4tpJsW0oVdCYg4/SUK03lyG0zzQqFYmDiN5a67fmmMmP9RlWTQbsLV
CzgdFiHb2Hjbq2yCpu8MjwXcJObIiKsrkZo1KMcFgJQH0xVUFbRpv43HABY/4PO6
ycu7dX4kCn2oPBQdpC9GoHWzDaMsT77gHS0Ipdo2tQ9ZG+lHGNzHBoE+V+9YVDcM
kUgv5wdZN3beHS0fkZ6QL8oeZEpKOXQ1R6rvkbTC/HeGjSptqcs1pW07wcoaLvXR
RYh2N9K8M3w+/ifkgxKYuexWnEGnneWUlfmt+MVm9qknZV/hdauRUxl0x5GtKbbc
tlbJX2IJpchswHYsWre4mhr3R94EBtkcPBzWJLGqx3EKvOfHKbOC+XEcRfrpzumj
CuKaZM+IHf1Mn99wYhKAGfdJif67K1oaU4PsIZJfWln7oUErinDPNWciTYwyw1NB
LUFJvHq1yxjO69By3rDbcO6O0CFgzgUhy1hkmZpRZ3f/Qew6pHX1Lj/cIMMLrrc4
Zo0GwAqx6KzWBDVdVzffWuCulxW62U6eKGiZ170zrwrQekFUC3tDPB++bhGSbeMY
Q5ZDy6BwlxdaYueA2hOvxrI3FpxqHNmTbIggmvEEAlAa6UQIGDQbu00zaCYEwSJj
9CpRmcpr4u7X0PAHlk1YC7S4Opq9iYFNEDyy8xXZxKSEINYufS+o5sV9Chrh86/A
Cud9ZnnKM0cMpw6Vax/3xl8KQVJOdypXE+e15YZgunJhCc47KIrlDoRYXt0rETdr
sMUZE8+dOpKlKX8RB7XdSbEDsVbFBFPVLDQ5bjpzK4XSSYOPZXleo3VnZUtZNG64
jSqPrUzirZxhG1pdjXCXJq/cEmYHybNYsj1gh65Z7TtNUBUGVEdtzJUc3PaGvcGa
P303GheTm9v++DCTWD5FhslvjNWqPSS/00jJYWhJsH/4lfPvkPQdcg5sCgojjvI/
j5YQ6f+dSF5CEnF9gdzdcTYYgW17vEpKi89ENZZSP5PIWGf6tW8K+RfLnYFFE7Ld
kE8qi8St7zyuLibLfAYuKG+QQWqIql+u7nUjUvLNdlysNGMH+Qrd8QpVVx9d/S9z
1APmli1ZylY+yVqMiNstVZIvIN4UwAyWuCWxBMuocDfOSSrg+WNUMxB9JaJjBNeH
OH719P0y0/Ss/wWIWF86OUE0zj5/lG9G5dU0AMic+MNinnvhArSVGPID3f0j/2sL
sFF7kUY5OjI+BtuG1OeaRg1gXxWjOGCKtaew7d7XQYM+jEzxApDS/Ja0ZlFS6uPf
HlDz60OPhK+u62XLKICXiNFNv9j53cypnZPVU15GCnnvRvntwLngW6USe+waJvDx
vNeuZC1noCU1BgG59xwq2dDPEDsTZ+YIF4GwV8EvqxTrFmE0bc20jw9PE6hLEPuY
608LLORv8suy0dZSBCQYfW6lQome5162YsoFAUk9hdNNJqHYNZHPM3hPDr6qcYlN
AU6AXCj3HOb7vTh9ekhrSssj9p/pTw5FCYBe5cwIUGjW2pxiH52glqW9DNMIHspV
ObeDFdw9SyG/JP8FKodDvhnwpoOALrIZ4jg9A37Y1sAuMJyGdx+QyDnWwqgTNq3s
6T4gfjfPIF7XwJn8y0Tc0DJmHp5uWEObAI/aPWgHG8Op98RV+EMakMfofbA0N5MI
uuHXgMYnioMqBYdg4GR0dEvaT3wPmvgdCo6CbnLZxJ1mYCJpKKhXHkxj8UMbPwNU
tZchXf2qTv6Xrm6sCNATwHuXy4NwkAgJegzR/G3rAGSZuB1Gng/9xsuzJJDzuuQK
JidynZjgV+b/t/dz2LXQPuI1FBb51y0HH6WGndQAMev5aR8favCVG8YT3gJTs+Zo
k6Ck3jifY+yvTahJdXC5l5zmRh7apCa/WiCk5zs6ZvuVplN3ewP8yMpoSdvgwpa8
qzBLlsy9FdGM24okNKYiyVyN+KmKdUe2tfif7NDGa2MUk2CWuT7dONwI6V/1Rejf
fFhwXL9q3aH3OdS7/fH1nQLQ5wA20o7X/CYkqRDTRVX12C1kYPAt0MRnLLkr0F0H
JJNyK4U2cQaMo82rS0kvMGZ8O9ZeqBwpgfjols7uYEHF0RMnvodMWoiKUNftwEEo
19xAm+2GXBgm5Z+gaeHIEiET0VPU58L5Ml2IOujD7wm9huxwG7KgQtp3ir6y70ue
wgjYliGi1oOi/qRtY65lRE3fLEg9ye6ig9LGMp+zUkcSYoCofAKz3U5hLy3vB/Zb
ZP+bJ+jvI/gipMcnO7aOfk6fJOw71HXEuhexqLWNU0rtENBPvlykR1WmhN8UYysM
msDJGdvOMxDjMgIn96ppGW96y0/wdu1ICbqsRM7S7YJm0YxtDwG3SQN+6+8EetJT
BO0vqC4A4QMZOmoLojdYBW+bF2yNE8QBeQqzNQu54fZpTo3L2xQKexJFS05l8UxU
ValRXPs25RH9K98CBbPT14gI6UTZv8hCHJusn9ap6amKfPzSA1EMUMqhsYmc29Mp
C7GkNIj37lAfqf2APhw0qRUXEiuVkGHvXV8/TmJsiCH9dsgy0BjP5xHsWKgrt5t3
IBZIpw4mdh3guzhb2ztyFi/5QPS9SQdmQMNcawpgQ9NucwsYksjoBuy+00kctDKT
FBDKH2R30b72uqCqf04yIY6fYOgfEVN1WMcb5dxMCq9qVaomno6YwfWWL0xTo+ra
c5K6zjF551PfdpYVGb9KpEH3ZliYofCgmnCUXU5wK4G4/+8pyOvIFQGGbRxmgF//
CPVSjKYwXFb7R0UFNhg/v2FzbNYwY7Eyn36OkuoIy1Sig9JSYVBd54B34hB6cfI2
W3pbR+SCNht5PfUqDT5pM/ggUS8siWlzXp20bV7xF4sdyymBEQGgNVtPQG22Ojet
ugMPHUaaHfSlI9mU33IQpnZxeZpxOTeq8u6TuwfGvyiRBqrmiQBZIjQ9idUptBHV
3G8QDBW8Ka3ajP2Ktq9E1FTZcF4cAZZyUlPTehbfurxph91mXbRLT3mtXWZHePM+
JQcavogAaxCPL0xTZpIMAWoCFTh2K0nH1lacE67Vf5JSukOcKmmAifPE17DIFMVi
P2NIDsJZfJhApdeRBDBjm3OQY8nvdXL2HQIh2V+dEbzlEZrUoDqAkpXE5zwVBbuw
vQ+uDMrJqO2Zf+B6dts4igYXI+xqpso+hGn/Rc2qwdWmjPgOwYS764F90axy9Wju
56cmp/ftmLDTJkfN+5liYtWt1TgEAW1tlTWJjqHKyfJ8hdYpWQXQgBO/Rd8LodH3
1+UNM6cN3gRBvp3cYGddgqP8A6aMwfCRlxbPyxi2h7EnSnK8TtaexTC7gMzPSXmk
Y44Z7wa8jt1wg3CLgbI6NC9+u7b156doZqu1aXhpRRIX/un5Zl7JnL4y72yPq8n0
pMt3pufl/nsEOcCOprjzWmslVMd0GXOmQb4lILKnraTXVDYp5HuvBv8S4V/7Ufc5
XBumUn1oFBPK/OsNNjYPBSsfEhmvMTJFnpagPp/1uMCBIETuSmj1nOeOc3waceMU
USrvsengTRx5Zht9dfSRjzeUeQp9eELqeehg5ANJKl/47JvBwFuSoi6K49cKohon
vfD5v1bH2y1tZk1fdINcUpblJJhdFN8IHuXUxJkBUQ2954CkZEBzWbq84HUESaHj
1CpsJ6+4EKy5AE9V8VFRiEAo3nZbfHTMzhtTZ8x6idBF+7SZd3C9o8JqGIWFStte
xvapJzwAx0Y193H1FN2F96rDFg+Ds6ZDyjeiaOHSNxo6R++bsajw71CkWIRlSOEm
gv315SGnDV8WVnNYjv5ZZns6ftuliYM1GjxzjR7DISFh+WKlCwwlzUvXgOL1WExi
uzXshejlCeXCg4wiHz+k6tXFjIUOkWNKkkocvHrNROtpc+eBl3RYLUHtzDyzRZDt
+B2kcrd9Ty7ZyxJEf/Zgva2TXb9X1dqIJEX6D/wr3pz23lTOXSO9aQcZONlZURoj
wKSsr83u82B27USJDMSZN2SQQWxnybt5OStS43C0QtQ6rkp/WdfuOcdEkjfHHv7M
OGqrzm4e7kqVxYepkWHhKrLc3afJ9xY/axhz2VkPX7LUj5HroWKpMwqyJ1ueC1xO
Y8YS549xIi5Z+Gqr50PpZayJ5uJmb+c3DMxUSz4WCAPZeq8g0HS4AA69GY5brDTn
MWjoK+tip7upU71zR+UxvP+Ys4segO8loxvWdDA5eHwdG2zgLBL0/xzYG1nxo60M
eXtaKrAwVSNUhRTistszNbBMRYnaxAzTh2ZIq57khqguRT9rpWqwgainbPmZRSkv
Sxri+MkpnF040WuRPv0qPnR/6QlFbwSpaYq7PvTOxAmlw9eQ0JE7Xna/xNnA+3Oo
25VkeWKSBR+ueeAD6WvCzKeIp9bbED5SfiWXxnRVlQ5rJGg3n1AVuyUzsjAiS/02
5jJ+N7IB1NSiHUQlgDFtb1aJqI7KoLOicIB9RMGYIINsIwIp/trpAwDrAlUP0Uop
3kAL9VXk/xOQZdbUSnMA6r/T6QTjVaQUAv6LqNdA5r8eZNXJF9GZwWhKHBCBIfqx
DRN+Q1ZZCqeHQuYBfDclRFlDRX0OUGjBEELWDLv6FERZ9gF+n6V9UXxi5RXd3KHU
JNM3y95lS0gnUtXacwUvv8w647L2ivm/SD3SzdCa6h5XJ6Nz6TCRx/rcCI/jRd9I
hT623K6/Bs/Oj+EdnhXyhYPnfYLy5cxw2zfEEWX6l4mlmjIXWtLZjfcHIs6s2bQS
xavplaK7mDoR7sVf3j00MSAeFaOyxEArxniGC+wNO8zY2GgnPoRvH3qKs9qUE1zy
3ONDz/Kwf/jsIPNbvrHa93fpUEAdGVmA8KJr+gf8+5o5GM84frYErGc6Ek2UmIVQ
BSNy7iaCvSn2kKPlP4/X0FwORHjw1JFHWpb6kGuQzIrIij0c6/ZC7zE4pElAsqz4
/XOXhRljM/ibrMYFkd8zL67/IHJqLnDSJlzspr1GD8MivSBoDCvffo+zbqelaXjB
JV8SveP0+WWYx49VLMFv7ctLjyVV851PYFv85eH4WOwcnvrzEXKMKnOWJydy/PS6
tLI2AMwlpiu8DuAfx6C5x9BLYIm4nU36NgqZe7zyx7dLrXH7xDW7WvjT9KQKXLm3
H1I0LOOQ9VGjW0wNs7U6QivGyCt+38veokgglgkvM8Fs0mOJLRDDWdkafNyJ4rlP
ac0cUrm/ucEXJpeMHKquLtsMBRfyOWcs9i1C7gXfgDoHGiRLn9+ZRvKc1D15ZCeE
/fiv81khi17ccNaZNB2UAufGmFjZ0xvNUS9O3GVrQYeP/qRJoMrUJEnUSGvLT2LN
zTSpwSpbdnAyDo9hdMip9B2oYMub420Il4nFQlb5c/ZwPr77ziUD4AQOc/xVd2xc
eqXL2cDSJmjqN/ynxvLVR3+ArQhERacU8NasIo66fGnSSEq2d4W9z5HY3RRjC/OU
mom57zgIyKnGMAsctQhGTPldoS1azwkCQhEZKy8v7p/Ak4Dihqmb+xvS4Vx8kr8/
av/FijVpFst1R0ME2mfmL3V2y+nxFFswAB/Yl70Y8Ao3LOC9Jkdq/ZO3EhURi6EL
Xfuhsn4L+BC9Xgd62FBrLY/AhpxjHB7+h+JtGITcSe0xCqCbYJhXDsRmFdkflpmk
/BFLtfnR7Kdjyx5orx6FUt1B3GcVirWvdT41t50q7+6Nxj3YIq/LQP5G8MsY9nPE
VzFeL6omsd9TMKsi0zIWgQQiM6py5TwVm2ABUFdle9HwAc72y8yOfs7342ancEzb
G4PBVGiCXthSxCsUqeVGcXwElj39JMl3fT+Uq3nLy2f0awjx42YtWeVanL+G6yDY
+cTX3DfV8wQxUZ7bBjVYFhT8NSZW6gP6P6aI2Fevz6qO6uAUF2uv1kEjymygSkIL
e+dg3WkUrAWrhXJQkb1hKn0eoLN6NlKqj3b7H/oZHtFruFYptun0AYYh82+mjw++
YzND6yU5JQtHPwVv2sWvuVdQ2E4mtceadkXzU438r9H4GBL3/H82dzIMRmPXtURK
J+Z0EnSBVMcOVgZF0RhWJJwVwkoOAPKt74pEDzTMqNv5THCUJDMeOZgvU4Lo5kIs
bc9+SSHOnHyN21R9QZn6eWdFa+Z2C6U8CQEuti2FpaC1/s1cJ4q4X+oJMK08pYSW
p8EZaoST5oP+U9rMal+hC7qdDNpeFU9Ex68kbgVOv9fmBhn3qb2YkJ+aI76BuE+r
lRPWKb6EfJUHhXNvNQxjUMeSxBhgYvIr3qDd/RImNRaSGBQKgYum14ROGdlkPk3+
SiMGcM68JkbnJWOWkx/HCUfuoiy+rIMpm+rXl6FWnMHl/ZmggsLvArzvq0NrqESP
t3RUQnRg9ANmUSMCaDSJy1Ongx4EYftgals+2EWPYaykzJ7UALdAc93t1ZaM7MVP
4Q1qcF/xIg5uo2t0A6XI+dkCs4q07wwaHTrC5TJAMElXzn59ZHmg+Fy7JTf1H5Vf
63n4EO0vu27WPCZ8R7UR2uqd0mI/9trVWkJG0uakMSak87NAk1HhSRX4T8sgFJQb
88p/QsOSBtGXJWPmBx/86qat/fPeCu+kMjiEYhhD8DFm/Ai8q8iXWMeJSPdfCTlY
jbqFnQr0fQGvlKYW6bZEXkLW0AYYgDcZuDl28EDo8u14sKucuZd1Fbbq6W5a7NAQ
JYJtOXaTmo8/4b/VBuSR5bKgLldUSCHzzgKwalxnbKTJoM2r48Q0ISPVzNC7wrTX
+f2KeC5Crh9x3cUeakLzKUG/THg0xO2L15uRq5bL+7WIB+KlYkYagVp0+ZAG2fW6
xa+MsQbL3Qjta8jasTCuX4JLtcwqucKFRJTcZF/rR21AbQ2Sh3oazj/p+ag+e39k
7geivWQpp2hqhKU14kLLOtCQoStSPzA0nl82Zr+ca0maQxsro1dWOYngSYx5O78v
ZdgvcWEsYyv9BmBf+4Ytm0MC9aF62K0jbP7PPLbij7A9aX4FX1bMQgozv50+VI3X
iWblbB3lu3dMf2i8wbho5IkQmGfYBK17PXOQ6cCMPoN4gKsIo6DZzmry0k88nMDh
xeaMxW0Pix1ogEAJB8/B1chVuxaAgbh2ofUNzp6c7iIGEFAMMUJ+jbW1v8ztZyGz
g670UCXmp9fPP+yxy6TLcNpYxCJMajL39UDkM3Jm6cK9KL0Ge/PdJeMSglQ6Cn5C
+HK6A8FHDE4ct87vq38AY9IAyAtdXX+GpEmrGIFnxEQDaRYXxOAvITZbYmzcohI6
89bO+uoHjHihGkXHgxwLjuS088AxkVT7uBXKwm+g7pya8VbMTgmVtEqqfhBTW4tS
1+yAyQY3YfumpTXGDKgo5DQLPqcpUy6MESBGcQo4g2zoIokX10WMiZvTYZsy9RS3
EvXWshrgCi6NGdE58eu9UZWP9wOUy2vBWD3IsspRc1VwbnsxK4neamBYDkxwWYwW
Jri1jdcvcqhup6LnbAbf5yTF31pIZZ2Tgp9q8zkHcTcfiOK4VAtAqpk8CqE4qdk+
HtmxhYdMLoYlJtn1CuoX8J17AnDBet+ZtflNDJaMY+IaDYWcJsv1erHZKBOikp9B
RAEWpR0w7gSVsD6chfjz4h/IP0wQNovPVCn2OqWphEQNQPqiR2rwKpGoYnxRTkfM
a1Hk5QGWrGnXnhATWVY6JrZ7ZwC1Dqk3+X+w0PQDeN3CULNdOcWAnIwKfJ7EvaZC
kdq8CHze29xSHloP8FXTrdB7Aw3Nyblrmsq4TGjR15aNRZLrqrOE3VJ3dZ2Bec4t
lQyxIbiRCiZemW4/nYstneYvLHd5ce8zFL3Pe+gF4iRMrXQ/2MCtePDQLWseXmAd
TTSK8JvMb2BBMb+wG7dkFUsb5Yh6SOeGAJmgi/inOIAfPbuYB84WEMOl5vywohRu
RDmpz1WJivg4xvjsoH7Eu/gmC9Qrv64zi8QTDFKhm8Ui+K82JAV3WxP9peM7cz2h
PRjjxmqKwZHVcsp9TQdK6NmLkGi2badxAl2gblAo3OPz0ZBDVh9pUmQU8cELQivQ
dmXPXGLmBxpDV+GW9rFGBPyEGnx7VRrDh/GQmL4939xNyhPfS9UKrfomAs54c3Kn
uUTB7yxNSYqnJuQfFDUwhzJTgqocFbpEWZ/EPnDT1D4cyLjzEMSm0L08MmKPjS0c
RYcff5KQHoDrlx1j5TaeGu+1+t3MVPmyQAqkXHXJzMw93uRyH71hCy0PPXtMWo1V
AIK/pOWVm9mdSC4dbRbItcpJvfQTeG90He2zyw9k+fwP/CTq1SWV8SVCVpoOLzF4
VGNvAoTIWsYP6vWfjQ4UXlPJrnAaze9CB3e7CBB9RF1DzmYw6daldbWFPczzoVIk
T2ZEm6SDkhFku0cD1MJCDvBwIY2OEWYkGpUj10j1mKWbgj7/5oGFPJ0HBxunPIua
KgiScNkCOV/4/H2bKezgqXqkYx6JETLSslyo/ECorbEOypwciZ0dSf/05Oa+mxCr
aGE8YZ8DbOcG9DCLa5NIGn/i+lZNmih+j7+5fSE/XU1F6y+6rnUZwFBvN4oJoskd
+29QAtrJ62cnP4OZUN2IPQjHMzYPFULNDOzKC2n6N7WJFtbP0InIyJmlCP8zI9fM
aFZIrid5gvuVN/N7Yy437ku+dwOT+BdOgqm9DIlu8WGJJd2OzrsODXRHmgTj0hWA
p5BVgyMjZrH+NQZl5V4ra0ZRg7Z5l2mhSTIRAdu0CZgBP1f+SzAenAawAFQ/jnCE
gx/fJtulqUwy4ADL3gaU40bW2BMWV1eqmD59Lu+OeatL5+JXJJY3A80CMA5MoGXB
GF5F0zuJXOnd0iKyfkyE/uxoKQbmkllDFQN8niTF8XtbFm7lF1M1q2ma/MTAzJPd
6V/zWnGjf80ptZ0NUMBZsDWHdMFkKlFj21Yz9NLMxmX2zdYUT5VFUuYlYL+fQM2+
ZEsCOAmNoBaHN2VrAKuP+px3hSuGsXT5rMKFCjqYfXePsjgC+1MkYP5xxba0chwu
xJF6SJ4rptOM/qauPXlqfDs9br8u2k4lbIfNIwfPEugq32F6LbMnN12Ku8VPYuzs
FC30OI7nejia+Ux6Y07JJUiSl2JDYtcOoFMbsRYJBbvfGQzLvCQQk9TY1MJa82bo
SqZT/k2Yxkp9Mc0l85SXEkeV2VK2Z/rLu9rtRlSj5zRDpZBrNWh25IpUDok2J05/
fcGdP2LkaA/7pURHGkjECQphIcA1zGojhbqrrMI+jfs6m1PeYKoFhPOztafd+vLa
Tek3Y0G1+jaOICRJVvZTG4vA4/LxcbuKnRozH5e653LJOpmCb9x3V0VIor74uCU2
7R3XrqNaKx2KdcU2LohW4WTOZlmv133oCo/5+sR8YkODyCaT52eyOP8uCkN98cZ0
JfyRo70jfYiqD0zqxN8KNlmEolzldBdaZdlJzlren75jzI3LOQLj5Xvr4tCRJAHJ
QWckgZF97G7UTe/tBpULrdsEdKydatEuRVJwRE5qkS17JesTvA8eINTFcpSA5ctx
PNGwy8k9J3DyDHTA9PxylnCO+15M/gghaXx/CJdpgJZcEdvyEN9vwkiVcJXfnjQl
QdYdAmvoZK7JqWXpGjJaHDMjLcwpl5EBxtwY+VI3/98VKcon+O1irUsY5aKZDOKv
kZAHbJk3XlBoySHaDVqFySpi/Y0cPuwrMVX5WfZZcmDjZTrHpfEfb/dr1eoOqDzO
7xAaMCeshhO/9+aCBw3XMpMQGM4gETYQuQEfXS+DktdKCV4P3jv5fVKLzAehHqsl
ehji3KtzTziauzCDQD5JK7LXXFvc4SW/Sriize8YQcy3keZ0pw4v4GX1A7TSQTZk
xFqXMpg5gM3dDON/LsLmBtE/VPK0wLVeKa0qd+vv2PyXRhgnLW4pWIr82RZd4XLd
ZMX81eBcRQusvYqu7UjH4FRuWEmeAzv+VbzCiu7Fgr0TKa1rQYE1zcpZXQx4TMXW
NX8r6Qe27Rcbu/lWDh5t2XOKBcnGpz4ZL6ZtWeIPC1ROK8el1v9K8/74r0AWII2n
5VLFtXTNjbAyPfDUxOHzNI8T1KCcUuS/muX3n1JJ0yOQAoqj62uSCiZtOWdX2Gyb
M1BEAdBGj01ErozK9NgDEi2MobrXOxY2+8u4orAoaAyUpffHU6zb7RjZQWc5rVbB
v4nb2lsqjbVPE9EAb1867vMYjVk0izfYmjWvBzn5eyU9aTgI8NNVpcUAzru4voy6
gInBWTbRCG8NtTRkJM6XLQqBx9cQAOjFXpZyn7yTp3JSJQw7q+JKGzXGIoTIIxK8
GDppb6Sji3mzGhaI8TosNAM7TjH96R/Q/RgIcO/6moWCdDOJbCWU+zIuitsSIL41
nnczrfpjaHoAO2rGqOfmlKcrSW3mCHqnESJjD27VWOlezn0eRDLrDKuTwSOsfoje
uaaNfZPZid2yhOLEbxDpIamJq/E2WJIYRl/b3i8+DI8iGRoCyO+IBDHigo6smB3E
gUloKdmoAMS4XTc39qDinFry4ulJPVk/z8xWMarnmFoa2Yw9B8/IKHuGJwGaLagf
K1nH4BHB3VqL96nnJDrvlY5kNkhk2gWsc6gCV+drIG3QjNalcWujrqdb//nYABBQ
oK2PQUsVQKFqlFKnz6tvNKLe3BChLZqxvRJIO8pALr0R684u+dq6SFKcX1CqczH4
R59T014N7W8hQawtfHsUB0p1HiVJB6g1VMfmUbY5iAS1AvdbkT37S/DPTJokOpo1
xVHGv/wVR/ax7Mau22KhZSux34bsqqmEYf+Idw0uzv69KZvYsvvsGPzCiYiJONCY
51IFl03QNTIlvZplda0KvNaJVe/ngHZGLJK6cbyLHcCbi+uR+wGV+ux7RFUF81LR
7NwoHDpEvLMfphTdXhXKFg53YdHRvETTpDGJy+/LWwwfuRCUS696EDwShPsN8JQ7
AqwR9YMn6TCBidfzjlcvb0cGBDZWfhoGQb7pBp1zFakuTfdPexhvS695YPpIO0Xs
dmKGWVn+z2j9CHFbMsMQ8/3lEA4Gm8TkZCFyK0TY1ADB9Xk2NZ861W2Q8hkRNnbP
vIeLtXK+ZYclKgmUqijqsjk1D8p0znCk2VtVVLtjsSS2Pr7vVkZV82llHJ64D8TC
zde9h6aXoV99C5YTI/0s95B3yly1AbEmHKSMAS5lcLdVYY792UXSRUYIr/P4DP56
wzfJ6zfapGU4vPTyYjnTWAuxRjaTI2H4xjVBG5e36CbUxNCGYv5Yqwl/2sCFbw/Z
fcksLmUu5MJIExp7y3HG3hdd32O8WJrMBg5IVS1iaHaL871OTFvqshbH20O1lJd9
1/Y2ESvvuFXIji4+UlgE5FHF4LoRvGf+SLEbHAfJNu9U/I/wXdkvL3qhUTU47utK
fXjTf7UNegXJ0sC38WkP7Df4hWnhYTDwUe1zv8vV8rnUzPlz8M53ngT3KffpQHqU
akXGMbVVUVuBhPQlZH8fZFxxt7hwD60x/rbFzSsIqxZGWx9GN2owxiEAxkpfrkK9
0CMozAQ8Fb0Q9FWaYDxa2+S7hU2yj2XFS0BWnsyowjaIVANqfhUn39sNZkrqYC+A
4a1OZT4J62SFF+uXJfP8JQRvNXiFeOt3dpJKYzmHpRM+4dx5FuFNp+wfTOjYRT/z
Y2zdnGll7/pojUo2JC/wy7cO5tbaA2dSOunCb4kQ2fhHIxsrRhBsERQZE6CUVzSB
+9g7R/BmFbC3hfldC/ASTnpJggOQSd0KgKcTjVgZqmaYMSgx8mt6hT4kjmTyqj8w
BjElgjkvo3bQjVCYjf2E0wLKwtSMwjydS9jQtXYqqIKFCBAn1D2fJklatm2Tp5+P
Bl5W1MfvUr+prbqSgNiX1ADSrI6gkSReKLO8kf9ELqChJ/EaTsxdzaopXiuc4zDO
B3vijEwLm82M9rz5IapjGGjVyfx9PRT3SSHh6VreN1Q3heWfdOU1FUccoMda1KoD
0dtGUMwA2pmPrIafH7zeIuj1ckMgTSQ4/XmVvFOvj9nymHmNi1LX4s0WUkDKqWfN
7RhAp+hAwb8SR1Rm82TF300vr1p6klArXNFVgyr22kTEzNX8NzcaUILrWhcQ0CPo
9jmJzKd37BB8/IF3oWYgA6YM222x8vZhaFZRVvln+XRNZYsJFT2tB/Z/NulY5pl/
upy2FEC9MS7M/QaJ3w6YUep8E+5HHu8zmwAYb/56NPq+eAbxuaUq+iil/dOPbyOT
kRzwEKwnCXO5ae4HUTN064WJFMy2nz0Z2bzTVCvsWQPtPimRwpIASWAu+56O8OIj
hspywuulm7elUK3niMx95Ywol7cUHgSgW3U6ZGM23RZsV2HTl4ytl6D8GZUpFWOW
bktFadzzrsM0k80QuiXO1XuHVBOy8hx3xD2LUt9vep2q/kwtgK8ANB52WAZLNI8F
R7tdZwDDQAuMmMozRcWgu31OLx25xH+KBoL3zn1UZyqhG+JYenwVEABNcbZ4+gvy
f9IFV+HRQ9Fs6zLJyp3rSnQ2wK9a4fFrgf4BD5kUtmLTHKQUEmxyP1qHDf9IX86m
k9P5B4wCZT+GTxMBKUqzpfmJkV4fhQALMC+0jBP0LT6ymYlr/9W9S7VU+7gAcBGu
xqaiDmDdGSRBZDM1dHLq9VsIQc1YFvVG4KtOIrjE0lJTetFWP4CGbNStVa6r6aav
Lzfm/6gptIzXz0za12rI660jjUMdY5Ei3BtdkJNu5DQ2hJnZisfCZRLyHgTzp0yP
WPsN/M73m0wqqRZfCe/4bdMExmEyHef9A987iffCSWFzHgO3UY6D4f8uGAmXKe12
ucxiQRDh1ibWpIFmfuh5TDRi1bWOPAQEzeu4REKmnpsVp/a8VF6V4WfrrScXzSD4
Dmh8MBQtX/urJ+jdx5zH2dC2+1YIH+Fv4DWv00xIejpefHW7XKmopSJA/WadHLrL
6SYU094CEKBTEsY7xV7QHNXYjMe5awg2Fv/DkJUSJ2nEQZ1ncsXJRkrnyrg6x1YR
9H3LirrFSUE0u7dyyDVwORX7UWGYbTu24Y+BygxWpWG1yZD5wX4RLeVTSRAp9Ra+
wL+6rhELJLdXwfCq/oJK8UA1tzNSaHG0mCp6qSYTOMXst/YXft2m+oLTF1GNR4qL
o0P6mQ1IUR7gvBcbS2LAnu5msHGHvyAbSAhyIe30212KP/MFNclDhz94VCgrJAoc
3o3Xq6niFdR0UZTqsmTRqbsRns72mxUjFlOLGCI1nKdATu4f2Hr0Aff5XU2dkjaJ
HlGO+8Fr9hANgbfjAzWQOgavJmqK67EZm4pRLNhSAQXx2dzMeKXjqttOazny8yw8
YDJ7lsxKtqzKUJ/VgJYRaet3lrC8eS4nWRxPPF3y6uq7VloyZb+3/srgrMk1AHrG
R9R9kpOR1GAyw5DVxzRA2Remac9DtyYbBapEroRioYVrbsILINsa9szM1j3mlGHJ
tQ61PgyCLV8Gb38+1gS703V5gwW08NBvdHsy3K8H+bN9mzskpJG2UpNqiFexI2mN
F52N7o86koB8I4H9+uHVimvPPDt/PjYp4gBqfdWZAtrcWFJU3KDGzaxaxzHokUJh
NjxMz4yo5o3Q0gQymH2Cs/SfaAb1nsvsQbGoYGw/prUk/PjoX+u2gZrBk35F9d45
Qb+YGhMp9ByvlXeAhBoz3wCpgtU65NKoMIrikMCZvMfTE3BInilTYVUQwN01P8VI
1l0ZKROq9Lyh0i8NfX6tBqql8zkq7bXq7AV+L+f5JiNWr5KtDh2TrrTxcBbhFAzI
IT+6k1qZBKzYRwVA0UvaeE4lYtHFghf9hOpKrOO3QVIT80a9Zg/XwUBy5wYGvZSJ
X1xCnAnf50EZt97vx+AZ/LHc1a69Q/sE5v7VU2Xn19NKV/bP+I81v3RAVpntlZeL
CxYen9+28soyaFOOB+ZRrG/3K5+b9pbLqkE0XXrqRhkL2AEyyHgpSQnJUjwGMsiZ
APSR29Qquy50DvqWBP/xhCIWumeq+54VWEp7XrJbvrficxGxZHJdNrbiHU6b4dre
+N85hJKXDMlAliQ1N8IngGHwxhfNNdn1efG7irzyWGAhI3gwfY576XS9Upq0cx+k
iP0qds7HECY0Nt9k7yiJ2rM2Sk98UOtjXrIT2t87PpzG+3/xGxRzNufJZUjlZijO
I6jst0U8XuPscdxceDCNkwsqPtKVZfgvg4gD+yYRRieFRG6QQxfRvZvg+XXlabTI
4TFarOEazc8/fJiIntVgg5b7Y3j0vUKe0VYYZ0wNDuX3E6uCNE1FgnyywDCIbacR
Wva9Sbqbd3YnVi06ReL4I7SggN7Dx/wI2AnpU/FPmFR/ErHoGqQhBvvs3UgeZu0G
rjsreZQLiW0HngcSEbEIbQgL9YwEtaxB/R+QwSpEewKIK2nuthNr9ZAVOecIgKgN
jjLO0zI8tLp0vWywwJIW/S78d2pkvPv2zvcI1OGkicYy49OU9v87LoMhOAyKAcFg
G/ugtnfivptO9CEn0sxYC4lG+zxqX8XHGZdaePsCu3WN4CUerRMYUs5c8GRLJoP3
N0sKcqLP3xB8KikX9RiOUMyfwkz1QNAI6Zr5a5tN77ZpKbcRb2rKR0wNSVNaPQ3h
VYJvaTJW8gYPnc500O+GqVhazrWPBEp8WPIXnk3YNCuWW6Cswn0diVRTjEzn7SyL
9OcEb5JZqMhk+0cZeoiZP2CXRJQuSh0z3a7YzxV7jTe1dsGecSzRYPQBgebXbXjw
LNERYIoCBZHlqjlCJf2he6RcUswgdRi1pQjgSXts+U6pPOrUBGUA5/xLOSx3H0tY
S2Igp9b2W2u1GZ4ejkjnV9uMDLiO1b4viRO5wuiLEjeMouZAhc2wO7RjUAv5Xfy2
1Sp0FLaHgCo0+g+0kKE6EFH9LtXg3UUHkOGFT5zkC2Rhl9jG0NTVTuCvGrnMP4M9
Jbw0sioQQ1RvlfRYvlUghXeKyJlBE/3UBVpmQgf1I5J2uiTmBQEmybb5h2klW4IX
hP1WipfldU+ppZH6UL2GwArZuzlyzwTzGTs3zqjb+LQw8/wtcQWzwl4PIeY5n9T8
8xnt2hLh351S5xSfQ38ywswpLWh8IYJD2yJfXRsgW68dlRfhK7+lpb8fH2AwR4Kn
i7RiLHz1B+9V3C6HOjj+7dEYZZqacYc8y2WreJrVDTD186pcsFJeP7d2lD2gHZ1A
57+8eFD2DNxj2LqB2RaiyextUQoMRRcAZsHPahERaxfbp5XvwEZ0QUPqv2UfrBVk
6tH9BSToAJR0hkitcIvG5WlN6kyxCuuKXW//E/aBnV1CsQBngI9pim/dE6j1BEHT
QYh7f5Bz4UCGltIX/BNFhOMa2Rd5a+HTbN3Modd1HUR3n44ljXjN3flMBiFqcN7/
gMVcs5ZGQ79l8ViQlmFwwwDcgZOm8bEJUJvpluG/FtqB63lziwgImryUy2VAK7P8
S7GVa55IDDHdNX6JJgekvYK9/EX3djs3+ydFrcQ40l8H71L+42rG+uY4iEI5CSgO
I5HBJ3M6qpEbmKkSymPG3rJo+4zhY5R+8e4FUmRFyyO5jndhnX39Srd9564V2yJF
rlo1bqOvQ/+mBYShF+fuPhMGu+incNAgPHLEmU3IUqtr6GAi7t9ipeowwkOmLruW
gUqPd7i1wJiTQJ3enkBTUsqpcVyGffKYBifW4/VW0A++5Cp5ekpkcID6/RXMfP8K
xW5N+LGwAOI4IlwfD5qwpbx9o5V1Tj8USqozyqRxRjgAaL0g4M+Porr8fdgkYcGr
CaUrTVLg8Ye8wDzP4y/UbuQo73blZ2hIcy4YIGxdM4vLW6bOMRVMTOXenWunPLkA
y6+KxuzRBd+ASB993pz/SuNojtePpstmszT1qd6m/reWebo1KFA7gJkOqW0RLCVR
MWhtrIa0c4BzvsjRcysvdGZdMlzkCBtAUUwTFbuUsFh8GfcxFoVwveM3IiXOZKVD
FbxTS/o9/nsTdWyS73dwbqhWTc2J9GuZ+C6EkEmTjhirLGn6c2MI7wXsLstq0lDh
TBWDuik2xGkR5zhXfm47RaGWPr69MQ6dR0ZFM52gETh4wBrfWWaJd/fT8f5oqpww
8qqB8KGjskfHXRSzKAQIlRxtIVj0CmEW7XERnybNmJjkMxe4O0qvSq6NEH+R71mf
YGUR8e5wLgvIVkzh/Z1r/le2l6mex8jwzX36BRXUE8yhmO772V3wt57AgiWMpOFS
cUvusi50VbGWWMQmBdF82uBvSdk6UuW0ARXXTQ/YiyUNfAYi1519DvZBUnBE0nff
E6irqW3nwziCr7J4adZtkuO7dxSnC55PJ+A62swfCRauN630PJv2MLplzKdhpJtw
YF7c31uE6eoTyaB/sBZBSSRsxss/KXXcvnLGIrIKyVT4ad5EGti04At3pIeqbFpu
Gg0im303PSUTlB/oqg6GQGq2MjaRd7IFECPF769jPhMIwiOOtZy6vehPxnyupN1y
cZLZfHmlCmNLWd5W5h/IGBpvQO2p3UTGWuxtjO6UogbF+EhW64yoKvjBxoiyKWBC
6qu/awftKli/Fi3HYn4PgmQ6kgUPAKm81sMiEgvHQJct3v4A05o7ebJWkkDECwt4
3waFBBx2BEElu3se7sLUZQXHVIRCY53iU2eYR2c87+vskbykvVfiTX3qEeEqkH4R
5QOx56b2CeJ/Mfaznd3eGppuFCpuYzTz67If57HHy3WN7MFHjtvvGgX7jMjNmYEZ
S3ym68p5oAtJt1icRmegCgjMGLt+J/VVc+hw4+HUSefxu8N63gMYZ3zh3V1y2i53
vkcEDy6d3uSAyO8fvI89CULpaiYBETFZjHXa3z4bLdRnqV9M8No0W6lmpwdjgUTy
09r7U1/x5og9ymHIxc/D6/cbUBQ9ewrFujteRMKmZU3/DwSeXIbd38VYieVfMRky
oNwl2Ak63UP60srVJb5yt4jCDN/KZNJKXwXDAXBbKDqDhQhzUNyl+yaC6T6lb4a2
xe5MlyXOOpbEUu6O0uEy1nhnaQE8ElQJyzmkB/lPKBydLksDWGRGzGIGwDZT2A/J
gaaIFKRU3u5iLQ+ObowcNCVTG3WKsdlR0DNnfwGGzRaeQy7SlAsg0YAwZUfkt1AV
PPb2msWRos4bvHaVkawQrhisU1ElduKYb5SA0p10PfeK5BB6Vw+LLUliQLv07Scm
+LyOd+GYWRuSeY24RB82pZ9MpYFfCiKtmeFGZtFttwBWIWnQYg1sDOiZh93pbKLq
NBh43yyx+DVFhXywxZP7WkyZazOl3iMdQDGvKoq2kARz74bXpuJhgkY1vHKVk5O/
VajErRrsE5/rLDg8AWDUXv2YLXVCuyrVo8M/cluhthsDn9DkP2m7G7RoykC9/c8P
Z3iF8Dln/Ut5Nm6EUgUiCPzc/wQOFQ4eXRX/82o34moeoBreEgi9Dm7yxpwkuv7T
T96Oifgxy0NrctubLxiMhho9aRkn0tNuNir1LhHGEbOaYCgVCsdFZuSW6SdjGUVe
E9IKMtERqHXE122N6Zia2aaMoFXZgDOTZyFqo+aqCK1mufy+iCOE5EQ+/SPsBdjn
YlrX0DryH+ZCzv1/EufziOANN1Vv16/g+JCUY+TVTT858sLo1W1cEE54Hex0CsrL
g8CyCnjx4wsuzJvzjoD9CmSxKZfQ6Htuke4Mp6smu6NvpG2087tlo+XrqWHvcAfe
+xhSnNSrHpIln3AI3qltEwqcR7Q9WGI6/Sq1tY0XhJ8fRoAaZgwlmnCG3z5S0NLL
iLBkP1q9XJ/O0fH48RGyk/uVc6DjWHuSwgWwwvmZ7PT6tzPHr7qHhUbu+JOvA9aq
D4Qd1u7w+fb+3sFX5NF9hO1KGUX1cAikoQRntM92oOlm/hsXtO8lhX2ZVSDRDfqV
zZ5Ufb/R3+VxvQwrCAjXLzogtZ6N+MAV15ObSKAbAYSlMQ7vfXS+DrytFA9y+j9L
3En97o2e1WfXvV537aPQXmsfwolEKeeU8h1U31wwYID6azJ0RxPXZzvgauKDFVlY
Lb6PMcsf9ZUxcDyUf3V8sl4/ZwIpzhWImn3Aqy0h7bm3selGm+YhO26p/nHXdz9c
uVcDsjwgIaNux95ZNW4JPkbrfM6lSz4yoteiqaqBHyv7/LZWMupR34miw3kr0Wxc
V65Wh6ZrrUzyqhWqfwLbORW+wkTSpmI8CnoAub+cG4/WnRBvsrBNDhSRgkDTBDnu
kWV7btPdUPD4Arkwr92xWfTU0KRYxH/mVwjbTjXdxDgcK3ePAJilPkWRVJokmjLW
HBID5IM8sE1r/SVl2mrPu0WQJAsuGEcXlj8akWX+jHOqPTzBjVy1JxjBJRJGPyTD
/pIt/zVYd9QsnyDqA63iZ5Ft/hMAk6TW4ofWpV5h1erjd7mrWea3UyQKxUd5kHrB
hqIHeuDP6YSE+HxQbcoaFUPbsKqPTExW1ZfnkGBfDmb8Z58ymbyK42WzrCUgQjzw
F7H1wzMEwmpIuHhFvShow6vgTzfXltvsiQ2JSJ8WR1GetKdhDiC4XtsbKN+lG1xo
/TkM1bwj8V87E1Q4+etSef+XSsMRj26sghsUwn14rBVWltzew5ukZjn3HERz9RQ4
yzkDAPIc1890Ma9tYwJNw47VYiRUkq3wU1rq5UXWvwobWT7todrUEiJxcjaA8VgD
4ZpVm8FNRZB4sHCCvbzJ298EmGWlACe4RpNbpQen9mL9tWbckHWziWgtgr8HFbUe
/FgaJtZ4ShE83exziR6/Qdf78lQOJuV4IaNkzbvki5kP1KwCJLIwCb/0u+rWt68V
TzYVGgfnzpk6KQ0qami31C+gsQtqWCm17OXZBjrfaj41oj1z8BPK6bxTkvc7eu8A
0CAujWoML0SIsGHDK24tO2Txh7kk+uPC+rUivSm0UUFy+LCLcag0RtoCEybEOSa+
3rThFDjpVcnIjWZiFGzF724qgYOT9CVKSgOvn+ekxKfS5mlgOb6vePU+4sSlQf26
whTEOnYz4DtKZ5tNwu2kpqzOJIeNOmxV0D6/MnmEVU3mfL3Grgykm6WnnomeGyM5
Uqqsf5u5psNcNt0wthF93MMkBXczFaX+3gtXaXoII+dvT+Ex9GvMxh5jLDIGnYPc
p/zkv7Fq+0siV/2ADQSyKkRLHtMLrr6gZpvnLmGkab4XrSw2ziNGn1DivC2xWz+L
lL1CcUzOW/JQsSrlB575NIRREOnKRDSDpsR3yWOpBu7kbMnGlMly3f0+s73rBxWz
xA/BPb2EzvQmgZSGNJV0toW2bWqYVudYiIXNr3tdDTYQnIxUjo/FHWC3sPP0P2G4
FDq308q2CbKN/4oaD8Xwq9E4FNZhfFdNDaAjKLQbiA07VdwLJQnwBAI+8uhJZ6Rz
odEl22LFK2OZnfARj4d9HTZseFpcLtgstOi6qk5omKuWc3vX1TjJsBmlMmy3WAe6
QD8M96e65geCu7LvMPMRr4kqyOanyK6l7GJNy+wCF39M2GT5Ny8Uxs9iRMPYB9f6
Tv6tmSaWl3RxaKAEPgQK+clZHEIpZPQPLhdlGdxwt0NTPsvabHJNL4nGctNGELJk
nQ6g5Ntn1w0F1hEsj3L9bEH9GmZqRkP1WtcMYeziH5j6V3NxOMTOpHolXx+8g8sL
5r7kow9aE5pwFf5f/oowQPL0q+DRNmTV9XJOQGPa8KI4YGYdlJHgA0sm8NSDlIws
5j6czOwmeYCmDT2ClsXdrGRxC7w+fx2wxwDnQGkDAUrjioLm1hm0DBpEtdbCcZPm
GLu2t0I++I99BR/9EEnVRqRdDXUcKYqIu8Q/BNq/Xh6vNj9q9+U7h/CYHw4iC4GU
sP/gQp4Qrnd8JifJHasAH0t2NHpRt8cSYC3hkpRBZnMn7ogtfpxgh/ippbdOd+R+
ItiCiyx9LFIssUAPlFVK6hUkksJ3Z9XpNiSgnSGY9QA=
`pragma protect end_protected
