// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:35:31 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
YV6EmKO0HqdNO7mvogE5RTLa0RE0sLKsuckdUkv3LGVv0twLVzTuITiHskxcOi+U
3W8q54zQLMdpTVOnI2Tap/kBB4xnJhs0tkW1J0lfCTXePiiw92nZEQca2F5496a4
J+ZLrrFSPQwBr8wmTq5JGdzpe+/C1Bqw5gobM8gDrF4=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 6368)
F2ysd4cmrSC+oFjCQVTae2fsD5iK4cV4l4RyDuNzB60n2prRTmjFwb7TLB84Se/Q
JUt5CEuPbl8dzLFv58dbFW3w0o811S3WKyObXPzkc1uwG8G60Id9Ad+TEvJ473Xf
CtfO19Af7hECcOSfayZJWxYrtEf8PDPQqwSaU4C2cYv2Ih4lPDnXtIohYUQuPK7X
Ng8XKxTpDceIfXAEN6KlUffUGs8Sjs1fsPNBATJxgFKsjB15kDHKzrni/vaXcHrW
vI5Iav1N47B7uv4+VqW59Ute0Hg58DC1bpVZMxV85dt4ORqKElg86uB+qCa5es6E
efYwUrLSFkiQGbToGO5wG4WbACeZlCXzG4c1rUt3R9u8nmpt3aNBwv2tMjav5XwN
0MNrUqOgW6/dxfpU4uWsp24TADCbt4nq4KaV8TG8uRWOUwxVyFOhI/RCfFMNU62o
TCmho4A7FdMEaminuzc2PQmQ4sqx3zQ+//+QFyk28taKQXGb8RrqxBK5YdAYl+VI
3fuTXHOBvkQNGvItJnHMp49t1Xq99+0p9LoE7GnAXcRktpSqKh3E/he3fjTfztyw
zK3QYU/FyCjFwp5CCgCUHclQh5DJsw3cx6Ptjzr0IUWIbe2vd32iXPKlzLSe/l87
yOKe+lxibjeWVygKgIxhUwGr7qTIpuFNwvNi1+9gXWXDmyGZZ1safkocCOZqWJ9r
gW1bMCncuFwa2F9FwEpqJjOJme7+518mucazqjz0rNMDysbQyINW4e8YbrnEEW9l
cMxRpSzAzJmNLxN+Jn0lj2VsB90XYdZsPt2OYg2iIZ/QVUJ9Od9xOwVrV9bR1Ud/
RbTxm+mMoCEuwCDr702c6wCtLdsOCNrY+BwrypjohZeZ7JCIvAV7A/GrPHtxyp0v
f7zQZGJYluiR6eMvl76LNmRq9fsiJV/24A6iuPkIWB3PiFmHtJkLaMq+vVE0R2yJ
CN6Hc6O4r+4aDonUTrInvIKacYV9KiqLNON1e+PYsU+S5AbA/c9vYR6uVHwM9moW
igSF9FwfSp25QctyYahnZAARF7Wd0sIMzvjqy6ue4WpSukaLfNjVWd9vaix+OTbJ
Q+ki2eHfbX1Fy/7VN+tt/6nNUgn9EB9uNCQAIxakm+C6UeJSXINa0RCzGmDhFe9P
T8FsWSRLdqDLJPk7DG7MW+JvC1OQjacJYC0MOi1peIN6zRHAZavQfiNFjYX1/hdr
jkvanDHQWN2Q84b0HXKvgG8a62gob9QWo/de0WT670ojZtmZpf7jWh9vZa2nPiDD
DL3ncoa4ujaZ1EzBTX8aPh2fVtc+EV+g2g3a8GXATxqVpGV5Dv72TI+gZAZuZ6fU
Z8zy2ZGMG+LE71ar9rwEWEOMdu+1lFQ9o9IienFNAxMKgUWr++XypJGirefhgBbO
TSgj/8jhUXz3EfDKqD5LyGstOgMf3z17wGCQzTEAbTOAakj1/YjvQVUO58lnbJ2h
bmMHe0DBkPKzy/fho1IXPUrcyoFkyl3iDIIQJ7VpyERxMx5JcVyIEKmS+DgzCIWV
ZYVhaDJX9xVHo/EOJQkYiI7cTlyrlKbEaKJQ9WD/wuR5B72ZVU9c4QM0Bfqpxkej
TUePnPyaOPeoNc+COtUVvaqsAs6pkMb9zt8EKjnlvh81c107BTLeEZ0SY5rVCLnE
Sq7KC08QBKPaOj2UHNs0grvljy3Mw5kspGbb/00g982/ICLyCp9HetngsMmsqzdi
cvAxba1qt5SxcE/P1Q7q18S3nGxi41x0I8tDHQb5pP9d0prYaposYXvZG/EXSS1B
nzqVJ9cqyM9jwwy4cj0XUlIn8uBZcVKV8iAHvlcEj2hHNtsYfIdrIHtnC4yU4gv0
dSBnc+ZLQJWZsHw42kDv+ZP9DvG2iUjvT17fSsmQs+VPgjc6IShifB6DJ5nAwfL7
uTpkuaikTAlSJ4l5PMYS6DB3gI+9cOFddlQUDal1lqlanFz5yvh8gp7m9WPENh6p
sDka8fKHftn9VzrGPtFgtIPODSojZY77wFNzQQC8sszynHuJwYz4Hojz79YNTn1j
Niey9+zOYPX91DurRCeZgGKsMCMX9DcKc829adPsX2eeYHopuar9Qp2N/HKOwnDZ
u3DPsY24IcMqRkmNi7s8G5m4xOx2Zn0/E7/lVG6BWj2utjl8hB6osChTpLrUniao
wBi61a0sVQtpUctMN8waEc3oyGUepHE8EfFiFLMx/Dr+ewP9fuJ0/xzc9SB3nhAQ
KeK3MrZX0EPF1os7VMJEdSdIw99K/42aOELr0jkF5xhqR2QoRTUGpuUg5ZlTwHOe
cFvpLA7XNO6UuH0mWcRoO2/dPz5k2Vmmi0543Sk4YfIGE7WAPp1b7DxLCLbBf1Mx
+WXzjBnxLtmnAg9U/9kjQgvOWNDhlVe32Cg9mHNe9omTZPKBtFEpwqqX/rUrSOlM
K1qqv0EnB9viY8Ly/EEFMKcPORPy+FVaHUwtKFCcpRvrW1i5aO6IJvav2CKXg8nI
inafhPW2Ywr31gxKLhZFUEXoJhR9l7ZodX+m/pvOEXPW0n+8qN7BHO3OjF7L2w2/
ZFLWSEIxwhmw9iM+pG1tAzCPfqyBfD1DcwL2NRZ+4A74wKrnd+2NA7gbO6BcbZyt
EK7N2rC3Z4N7545t/K4p1vJS7KKYsAn241hji9d1SgLHx70di4PqRTDHQlOnydhX
pg1wR9pQDhCO/2c/bqfOW6wUuzru1i/XM3WAT5CFldiq/u1LSYvggX5Zr4FBNfK+
zJsKqrlXoUSQCXG7MSaAb8g1qsEcuG4paJHYm8SXA2mtod7a8N2943AQbHtgnRV1
VBh/gFBHs+y3Mco0fC7Pj0oN9Nm/8VGAzQ7GPeraYbwXZC4MSuMRrhLqQX5+ydDK
EWDDQsT//HGSVNQ2MLutOmHQohRD/VsKr8akYkU72iFoiTakidO9DhVmv9Fd22YR
nZeYYr5P1TtpbAc6lx98XlrWjD7kpvUVp67OMWVsHgPAQCRoY4pS9SYDOGFSNG87
Pyyc7RBSZ1/6PIEqbAne/RvuKqe8nWXtxbirmd5AHJy5OB9b3XQA8So9jDl+dTTs
nzIQ2YYOk2CcVs641vGbImzUpGbKxfzrmv+n/3dAa1r7oZXOpeWLiQRQYjqzRAP4
u8Q/KC08T1Q2xGChIuQ5lBBdsCxbnJysgTVLxWWh5rmgDIaOWLkYGZndVox7EhTS
LdmSqzugEDuQo8VRuJfyaRu0gwTTeGMYPbUtlT2yS642yyKAWjC2qS5pSqdwrVTT
GnkI8JBLvl+zCtJvxOLQaX/1MVciQuZEQR1teX0HO0/BOGUWlXIhi8cocKTKWdE/
pt6NUYm/cUSsBazPXTjnRzDExi1gsTYMI5q9tc3nSyN4RK5VdUJqMbXpn3vf1FgD
2YL9e7JsqNtSa4twkBFeUY+zFecsvyWoXtvtMGo8tGY+6cc/nyOqBlg2CcpRi1At
V6Sn2drUmIB2wgOsWqScTp6S66EUcB2LkMjVAcaKEuphDOqx5UDM7ToGv+bp0/GW
kriVOqEJv+lePjb3Lp0r3DC58SXWu1uMc7VzcbDaRVZR99icSvPL+G3BTRMCjciv
ma8GhRO9tfZm8VZeP52kcVH43xPMPZB8VMN5ceV9+2ennoj/ce6oinHAgNsxGoW7
MbQhR1cXIdqmohm3uha9onqzfXu3KSl30ko8GOhVtd5C52xR/KlzYOpP5Nc8mfQb
Ayf3s+6dcJzJjk6dHlRBDrR3euWcfpOZ0B95aSOanySw0NFivpekVFymI3fx5sy6
raq48pDUAGeL8BcRSb+mbgBD4L7cS7mpMRFUCIgT+WmPlj2OwZ9uaFOwojTFt6Vt
dZZcSVeKR5LoI7yPfITM81IdeNUaTQNLTncvBoJN2LIsOk937Ow6++M1D62gbBSA
bkaiTgpKWPdcPa3ZX3MGax0ZKAUZlFDOemj0lWviei3O65KtTrwu5sv19ddKmd/8
M/2WCWw5SW/p5hn/ul2bQFa2BLgaycKIu3Xy2S12uBBaDmqrYjqCj7SXO4pgAVvf
hq94DpdTM6MiKi+3vjbqgg1Wj0pzita4pbXgZt7NmyunlGUPL+Tk7DCcQf3KwArB
o7W4ckvB9Jr4jNDR6jdXsU5JZq8loyHwdmmkD5VYbBdvNmr7Q+unjUFbaHncI8nB
pk3OTFxgVEeBWNECSyzNOSPiyoN1KiH+rTe0l9E/pExHWmfIsWndYeAXjVbHz42g
hH31EayxyWFunQdEXzY0g7tfJ6o9+jOhK5Rts0lhn44jrusVMi6ZnZ5Ed74uVCOf
QgrMcyblraOeu9MNSAmRa8OvcNKqKoR+VDmL5DPcxHOQ12hhutaIYN3erxbQxkxZ
RMi3vr3hGBTWv7VGg1lPwrBfK7CoHmXZ8/uilV6xXdNu6FoRWDWQ9+VK8x3VxUYc
zvQ1iykP9FDKGpk6Vq+D6Lqry79T9C5BXucJ+IbOu2yZuwokpwkoWd7jigoCjRP1
krUCjz8C1TqzUuMID3IOhL3MteDkH1sqgxN0lEW7FffHWN/LT/gpMqUMpzteTG3r
b3dtMBSmgimikj3gG75Aexn0N4FRGHFuGqyhRCtkpSzHxN2d8SPjeBj1cj/TOw5w
L4M5TR1zX/uCJnhiH6fNc+GHixqc/qbMJH1irjSs56DPsFhdA5bSkbUOpOmETFKC
ctdX+hmwhVtSx2rlKDm4STFNRtkBP/wzLzN1qqZxJ9xCMPMzSdRzqOdcJYZLRMki
yDTWLSid605ctnf8xPpHrJvfPkuZtJgmlUUXJeO4+Xoys4+PMNRluejhO2qmeUy5
d98GjzbpuUVVAH9gjuYjnCahe05ehevlSjWkqb5Rn5Eyn2FLxSaoSF7ilDOjaOQM
fW9zBDLvAmbG9qyU3K86aheymrRI5G+NCgbrVVpG5mabE3aQjV4j8hlYxCU9HSCq
91PQyvW36ZgeKFqeC4xGPqfk1an2EOAnF71cD8ro8j3mHNa83mZ47oYUUDwz9u6w
ItprrkUubliTxyls048AmX+lskk6dt5IFG9gFliUurU7c4YYHYcvWpaSJgdwYzQd
jnu9jJWW6cv+c9oGQUhj4v8CnqIci+N7H86A0ilobdKYkeOJKaMoUojlpO3jj+pG
9p/Sy6sE2bowB1JrczDyKKHjd1f16hgXCZwLEkvofuakBavBNpx6Gno2SgEdwtTz
f6pqAmEjNIP3XJd4pgq0EpyPMXeca9tAxSWpAAtK0MS81Adh+TksUxTcDPJLidEp
RFZEFZcw3CY+7mDjHNqYlBUAqxnXq2jdpYgtZtpRTIls/67ZbqgkLOB/Mp5azZWO
JsLkDO1uuBtDKBTkrO4tvqpLgiRQHLxDi5BS8o3Er4avjJ1yv4MTkarMYKad8n+D
dF87fOyMvQHkeA7RrNH++yNWHinWYdDMl3nSXa2kea8JiKcv5fjZva9J8S7uL/Dy
9T4B9RtYl3FWF5grUKn8JxeRM9wip5kDdc2aqDe6ev3fdHGD8JqBU0qKvTD4gxF6
l7M5GBpv8YKChjaPmAyT915Ubmz2WKU2bDYdGfrgS3y4AGMMDDaYO+1MU35lmhWq
yxEVYXkgY4XalFosYUJsPXyNdoUxc4lYnQt6w0gS0QIftXmSaxyosamUwQ/8YbBu
9KMXqTqde4Qj6Posp+JTS/B3Mdl2eUvULD4G1VdJPkbJqb/Y07MkrJgGxpKqqxa/
FuTBNklClEXW2lOWyUXWy1860bP+my/op+wKgBYr3BXmFvpA3au1KRiJ5v/DvqC1
U/ZFu4XbwnUZ8ze5nAZbWSbYUmeipJqqEIEVxuct1Emus0BgEyU1ez7zqd0Flq4B
sf06+2s9reOk+Tc16A3pih8hQjv4u5qnsEQ8Qjd1ZHrDrr8R+bRuGmtr2mUdhzbq
8LrRlbMzok9T15IwjNQzmZrlIJteCOhHJyRJvN2bMqeyRdlzlIaBVTQTRKqw18CK
Q5TG+gTykuen3LBp1j+uMorQk0G2oRefprKwTDsBbQTLsrS+4zVVkeatnqFuHiLV
9fRr1gz31HCYzRy34kx6k9lU2+comH48Y+XTCAwDJ1/n6fYxLQif1sEzs+HP7kHs
ElLGNC4mFK38ezQWrJCfaQpApzZ0BaLvYM3c9YDO9L1cZN3nA38YUaNOGVXS2usF
cXFEet+0NILD7cY8REgAzBHv/9JjkEbi6coOGxBab8mD0uuAihnQ+RFdLfGX6WnX
86AuesIF2pXy6bniNSj85G/R76q0jiUGPuu+dkd9Uy78W/lX7NHAPPKuiwgihTj4
02uur3ekpj7KTXnAWiIScDM+KQ4tZ3PSucS33HS6xaGYsykV+CIfQJaJ0S8jR0W5
kQpnayfQKdrglW37dnGZzKVK8gQydFdf2J+r042Mbk2jz7jTE77iCmojcHRpVzr/
kIer/2E1d0rKlRHMK7J/qLdxeNN0rp2qoZ4tCRO0QgRHSi5wU8mp+zMLcOpBF/x6
SBJFymC71Nus580E3y0/TmbE5mDokFgantjfbpqPcjOwz7K0WHSp7oeJzoPyyE1i
TvrBQ1E4sQsCtFYnQGNRAr7mhaMLCZvSmfbmIwlBbtzIcRpO5a1MgeXaZaBM8e0V
MTWpIvBie5nlY/bwuDgP9wkKoWcv9aQoWyGuwzz42rHZ8D/aLMC4Ud8RWg9mWyFa
zySSOr2oqDNvy/4zQxQnFD8ycunP8U0W1ezBwS7IdVuQRqBenC4XvlX+r7qRyn98
MDCGjMCt1C7PE+b4SvUTFvHXVlswnVrkYaT3HCpRxTR7hoce2cej8/THuiWj20b0
2f4PobyluPc1NSrxr1UteWFfdDW7NMLuRDumWf29QcjcQmYp1k1qL3KTgXeqXoz2
4V0oQLPKIz0mzDBBUd2ZeDv7P6UXivcCAynrnfo3GofVDbqS2JAT8rx11EculwQr
dBoQ88tXkKjLx8Mb89D2r+U3fvQTTFkzT2SEwfhLTTAjwJAQo2iq/CBjRnGw9VK1
MO0xeGgSYbgZ4wcuXwEBjUsmefsIubH057aWsiVktx9rvSFDgZrn5MOL55mxYMee
WRrYeDsO4fWJS0Dxqo6g0xYKMh2YPQazca4f0qOP9lG/lJnRPxSb0nO25q6Z24vc
efDpeYfrkWv0N5sM0oJ4pZjZ+TOxc9/Uzl0MISph9F0MB/BnXXlPbujr6WSgxrBP
5xxBB5PH01K1PTO30E3Wrx5v1hWiyRKcrmRKgupCX0mu82EyrlnlEH1RbnG6PMpj
hXpt/Sb9olIpTsJ1jobj+JREZJMAQsLsw9NOyj8r9BcCe5+tNvSBaTqXdJQkCNtg
JcurWhthJJ2luLJ8j02CSBvq1mnls70MqsDUzKg2rInRGw1bT6vHL6roXD31tYer
8teGAf0wFUOaVtUepy062esDIqP1bF3Y+RXadGrQMJaU+55PlZwImYwALZpqE3on
sRcz2xZ2nege7NGBtBcsaBa8P0iunZus2O3Pc9RuGHZCUkp3bab+t2Sw67Kqnzlb
PRTNzx+Lg4mUicbWwWkhHDlfABrV405LzB2MyUfSY99Sgv1G4miZzehPE0Hh+iKS
suW5CtiSPUIXT0b8rh4gLWbS4EiKlqYe9sEEIvGVZbNZtxQvCrNWEuQa4Pb2nAIn
7SgZkTNDaoy1VqWW0E/eQ5bmlY54z8R15wsnXgRieCDa0OMfhgJK9mc9qGil7brv
Cw+6U75g/rsJjALfGDx44C+O5rWldBwJP9tvItKQEfR7J25fTNPczgkKBsNG4uLz
dB0PHQLO8r4JVS5iUt9v8FL/8BFgyLtm+hq1q1Ae6bOedgIVcayAHqXREbwMIsnf
L/z99UHlkNd9w3M6m/Z/TcwOjcmKVQmsn7ry9lgohrNCkSMHHUnSNugICzcCpw3Q
opPkAVXYpZychlmJWXeiK48ySiHOM5QlzPMo5hxvLg1fvJNs+Cw/RPSFxFy1/xC7
5Wjre9OSPVuTyZPL5kR8VRdUe2QYGmsGFn7ks/4BoxvBrC84S23iOXxi3hS1lE6r
v76356LCuifj2pYloqav/2uGRHhD3FD9pSaf0C+oLQ4yvAUlUhQ0tz6PL5L0Hzzs
hlWfu8+K4IO7rxMxCXQKr6Sr8mJTL93LEwItogrP1jIIK3JUSWah/7AKbNMSZFiQ
8iDbp0SIa2w+jyT4NhCx63627C+g/a5ercmlTCfsWIhdRG8viwvuww2eCqpfNweW
Dh3tKOEzaV9P1YluZLN1U+FXEN4YQrkBvoMF8wJeRstoferF8CmmwZzPz737xM5L
oUDy4tNPptVk0LMvs9ABdBF2HSZn7bucXuYXeQ1mjPlXbwdQYuhga29dYNtcZdgO
sLlQ/j44ezWokGzCkaXeHtukP4Rk4odIvfF8TEcqk1PYuN7aAPUysnOUqjT5eMYK
w8PgAYPXe5JoByQ2d6n9gB8OIk+CyVg6x7KbMecNlAnKIkULEqbXuhR3++xZufUu
b9Eif3jwfFxciKVR07pYT4KQDCza+3AaLsLDfZ1lN1Y=
`pragma protect end_protected
