// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:37:04 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
gzdwZV1dI37YO9QhM4pKHcPKC5uyJ3xB2iOMFPslBlHUoWeLsJrqjmCtfXuNJ20T
vqYvOrC4lksOjOvfq5oHU14xcX9qlcpDsyLZiVqNQxZMgikLp3QtFwPeGVmPLFUY
7EeB2J9FSBIbVD49eDGVD4gNUbwsf+wbsIdSm6ZdeRU=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 38352)
J/SAJPRSKiiGagXaHFYToe0kzKgijuQtjxhSJBXsvc50+C9RD7CYZy60xxOdiJnh
Y/RfFJA1SR779LS3yy46Y0bTjlACF61rj8Swdj1OvS7HlCOWuQ07fPsTlmemicmh
Wf1mqZge6pIZoAXDM4chrr4WGp2W5M5DU9F4ElurMkFbNnIq/Vx9TwkejXbCp5JJ
b+R1hhn1oxFdr7y60eVynawKcCaUIcipofJxkdl7E9ht2D+5G/uUg22CLT7GSEgt
R26J/OyRDi1cX3+CMgQQ62YIGO2bfk0B8uw1iVWuW6hyNmWHXOy4typ2zCjylxFp
pjvRsKAGDOmxYVKFbRhjCV3g+Cie5vPLwLVLyIgGjOqu8by6l+NohlK4+1Gua/Rh
1ZJOirQGsLAT1KpEAH3+INceB79+xb9oG/w9BWgD1cDgxLDj/01l0Ee0Abv547O5
XmuBjPSFOb4H/GIGcOzNOg8qUt2f2WQjBznAtI97IWoDf05BBh/h2o0LdPKuv7PN
IUP/dFJG06DZE98iJLJ9Eu8xx7UTXU2shyxVaYbu0kyWSJHvVmVhkp+4t2kUiKlP
cCB/bZi+7GoCcsNNruMSIGHERSQTbQaaIQsxl5IHnHiia89WF91Q82Cb6FlnINIH
DSzAAd4UGRmzHlkAGfY3kqy3gbM9g/9ZxEqgYBihmWSe0SxWPciiufH83hi7DDk2
cgxmJzs1D29WuI94dsVcdr6BTWhX2GYjDsGOuL7MseSMbafOCv875FHN4/yilLZk
K0fUgTZFoV0TZLcWAuPVdVloxmF6mVlsi+KMTNdDE4mFjQUrJ8cK60BjpMFhzlCw
6e1H3ohDSnU08K0Ys+6u9EoDcIkmFRg2+8S6z9c2WYPd0PxPYbobqVNq5pKxIJtz
zVZ7sdg69qkfjd9mYPuea7QZLi1lQSQCVZ7YpgsMJmHMdryGMEM69MC03+iDod9X
MwtTLdb3FPeMbmhyz/kO8j7FTA6aCL3G+HDDWVTaxx5CvMPG5zOgoArWufZUTTTQ
QsBt7nqOLPjtwlKK70tbqPbIaQneC+WH1EObfuY96cWFMhGyNye9tI24ppd2zdhQ
hk/9wvQvltwQFqwjFXNxLXMdYFblhJ9KCmmNN7OVicXO7ojS0Xna19q0L2WmsPm+
XHsWsmeGx9z78/N39XpKxnJjDrVlu2RRtCUKf/vCNyL+RQK4YWtVXfPXmSvACHaT
c9Rxsb+nyHCy7AUeBfHwh70i2LDlWKGimmxFCX8tSuQLw32nMfXikBSBwi3Z9C/n
Cl6J2z7vqxLBlg+YMssb7SH+eba92hzRWtPzu8JSaFp3W7kdmljdKsp13KvZFU7N
rHaFtM7OIXToHY7AV7SlC2F8qQBYa9H2vuUyBDRCHQntXcdlGQTjL7hdSeyIWLCt
bCvkmBGnHXOD23NMe8HOblJDlo6duc0uNpjV99TXwZAO8+PqsHwE1bSl3Cbn39Ly
HPiTxQnz0rsYSC28Dv4cY2zI02zJJSAqOdtJN6LlTwQ5HrIifroeb7IO3sq7KAPv
SzvsbpENzPvM8pkzBRoPIT0pQP9Fv5NS0vXvpSUQqKE7SbvpkKQ5hhbYO+KVqx53
g/ucpYmpY/ee/Sm+vVnNSVyovAI0kU59tGoIz9PfX+M+BVJ74A18G7SZfoVGkOeN
FY6ulUoCM7EjqC9/KFQBEcb7Ti7bkz/a/kfi5qQXhP5SrWTWTyHGIGdDqJ9AKHfK
+d5UEHGXkk0g4SkxP5VXMxZaXWzE8w3jf7ojZMJDsTvJkSU4LV5zfwz5758nSn5I
fCfQMHVriC8VhB8qnQgPHJSerYEVMI8c+oazBe+4fXEva+hQyURPUABGbSQDwQfD
Lxsvu73sD9GOhoyJMYpiL149aYSYvms4ygjJlCUAuh+Yh4tGc8ojQHaTGSyuLvGi
R902hm5896UMhwk/HNgDEBmqsEcJzaTd0Ry5qg208BGLNlYglyf/1eCStjy/owkB
HMHuYKzt1eHWCRcRcu7L7pL9a/Gl4tt9kNhG0mXZ/+g7XJZbYKvv5Nj9j0XqwXfI
/Db/Nfppozick0lgIrHThnQpV4HyYqbTNK6R+g0lAuSq5ad3F2a9ZDlL5pnJJ3R6
YSMp1xL+DgUX1fM9baNu9mn5PJQ3aCTQa5zbj2OIdahWAvOy9argNooO5nMpQM2W
tz48BDLNlF7a4mk4I2GYnW/+heLRDNYeCplgMF3JuZwUlwfFRE10peGrG1oeav2X
BborfbUx8Qp76m9RNSklk+nL7A/cD+mxg3rITB/CFzJ6DQ6ZCvtRNk/MK1YbbVDO
VaIRfsrZsgMarq8QO0dyltG6OIQ6CecgSXL3gXNR1O3akndAAUgSu6mdWElnI0ft
+iTdi1SThurYh2thcTx+jt+dx+oaOeveGvbfCujBy5meK9pd7rEle+SwU4lwmnET
ejNyvXB7ZWFUFtzD/v5kCFMMgsmggbJDjxt3/Md9yGnSwYIIM7WhynP1SZKoECQb
u+10q8ujHIX30SF0J7YAMrtTV6YvoFvR5duGrT47IwlNnSHTKci64bf7934yI1L+
XAZsFYILb5Gh8VUQAh6cOJkxuwHpcsIZgX16IT+eQWzBVefEE6edqrzFanM8OKq1
1plE6ZYIoCXvhAeF2jKvk/jpGZt1JehFSubYCC65thHuPSS5Lbow5ulCKYVaGwwl
YBOhwtWcuxJR5z9Y9Iwsx8p+Y9J2iHS+0aaM3/YmA51X8NxOI/uBFS9Smg3DHbAZ
UTcoQJzakyjmG83n7XzlnnOzwH2TbjnKl3bGWgJowkJUUHN9fUidZfWeyiia62Iu
5P5TDob4iEXxKPxksHVtW/p0pLrFdIyONcKbBvaI6OAcyAXTX8FV4HplN26Wv4S5
kl8T4hiwn+d0E1nzbtdOjC182EZh1Dr3vp6Yswfg3CIuA/akJbePqOASL3mEBJD1
lj4GCVV8oO23zQgscfIiA9qQCy9a7uzSXh85qZhc1Ml1EqjNgxAAp0T7Iplqb0TZ
s22ct/wIhgby74PhREPu/N/SmHTeQLCH2f3I6JI9hUfFlZil/KE47eqZgFq/CR52
/9h+6BmxS6bH9Hko3zolEiGozqTfRWXL9f5Et0ty6qTkY5B6VwYUz0roF6DO19JA
UdORTTxpA8jUxKIRJVaqwoDnx7Bkd/0yg0lu0wzjKgirFrl33Gsmr+SpxKsygxMM
nNiwTO6xWJ7szoKSqR9zlP6cExBA2YBlZQk54OOi+XFbSL9dGYSbZBg3snh7GFeD
xjzWX/R6qERA6kj5VuNZCUxZgK7Qte3vrV62UNZN1/Z9ydhJOlL5e7i7hR58dMT2
ZybZUORr4xvKZT2ApMKVfC3RNivI5YkJfkZLYHkO1RaAMLuMPBRfzhE24MXhd4ko
dXLOZEMY/ODF/+x6dmXnhkWxjRcFlGvDN3f16YxGm7WJzQBGtlLuVqvQJdZJYZ+J
Wod4uiD8c508MQZMDZTSYCs9ThqNnOe2SsW9EMTnygzhMvRjatt1bnviuGDgzcNr
XkIqN8lj+7WH78xZ5Oqg7sH3w2CQxGQeKJuDoMjS5XJ5SRNAL+MCmSLqovozQq8H
AKB8K+h6Qhv1a9gh01eh5pTg2QJDTetg/LadOtKH7RhqvXCk0zNLfcDtAw2zFIKZ
KLjMA4KhNfJiI8MMnCYtApKIXdJ0YU/0e593dyRhwnAxseUpjM9KV7iSIvFurL5W
qohXsDl155Tth7EDJci6EIzaP4CuN8qstTYylUx2cwzbUzvwSvNoUgOUGi3PgRjQ
021E4FYoXRRk5kNWbbykInkfOeZP07SdJF29PsvEt+4zhDT/IgvzHLaCjL+qhhyu
540iCIicbO6PswZZCxuevrc+ge6cOWtHE36nqX5tY759lr/fhLQirN+d2qafrTRH
iqw7oZK9ib0Dfquq8vFMp4MhyTiGjoO6d1wTmRcSWYo0GCh7AHtp9IESBbDEgqDZ
fhSai3d6wOvDyLXLJN57ahZTTl3MhUwHsApxBIEoHOnuPYhmE6i8VPfrSBAFZgpV
HpZm2aDmm3jGVnckUI24rg/A7iD8hhIOVZzd5//UIDnlQwOeEaoBL9DsvpAan4QT
GLOCwK1LFc0bcCNNPWzVuRKslYpcmJ3tf9SyW8ve/Ee4/X7P4ZUXL30FBEpia+bo
+WMTMFUzVT01Eg8CclJEcN1OZoyt9MfFVWgppVQVNJpB8agcjH++2JBLIAPZIsF/
2iuA9wngEIEH0NzUmWELRjHcC6zhA83iyHcbTGCiW3jQwl7kfSUI3YHUhY+XNpOE
9Zu6Be0QcITJoDe9JMYUmb/RP+px/GUvoN3/fqVCIJ7S2JdRepkjBgLvXwOMbOXY
bjsxhVUIA/WUdMFa/jW248bhDp3IDQ/7Cf2oEAWCJTXUiMizIoRjZlNHNYkK728c
b773e5IdYWat6FmJTDvtmLZareRVGJ2Hg1cay4eyfj0dt7vjg+7vPLdnb9P6VYCd
v3urpdBYxN8uAFbxsnAkNJfg5oCOlqVJ1sgO+YKPy77be80OGgNoRTMcaPevmnuU
0sIInUEukexdSwnT5PG8k/vKzZgCcPxVmrVjdHPR3+bi2gBXk7IoZxrfrGMAFcTd
Uhy/aL3k4v6/AajVD8Fpky97xg2J9330ArnDyda5epkEa+FyHNrSHegjBLw87b7m
GOXEJnOR+QMsgjWZ+SgnPiMpdHR/onalLmQvh6EhJaHAdouEGwCXqhoWKVurBfff
R7OAufjc7NUFh8w/bs3Bj/lX/IuvzJpRgIZ165OUZNcG/9OtP1h1VX181tLfwq8Q
sQhrFuBZWhpoxQ14ADu9VuK2ql2jbG/0H/ATnVqWsiGWbYDvdrmJO+4g1FkMmjC9
0iM2BHGQxdxkaZOA3axYveG6+Q4BAgmsfoTyAvt5PR5Fm6ijiKBPPmSPMtAyX/KC
VkixY9BNuPe6IvW2yB6lKCMlo4+WkkktgITjut2smKYCA5cBO3YPzUTJf1aNx0V+
bXSWjvL2iJvBGyY2HBBqJ4b0FEiXFzBJfxkEF/Nenrq8wiCIAyIgA4j+37AdRtqE
eQ355vLEn88YtEuri2vA6bQ+7nwcdVylPgd+webQ5i0ePOqKlFYbwfP2uPPJTWtn
U2F3/zFGIOmlOMBspt0Ls+Av/DE4CsOOAv6kUPhRSJoAFhwo7eabnxFOkI6R+7l7
FTD53SYQChskf6nMjhQCDJ0vDfseIRUtiYQw4Svyu4Pjye0lC/37g0jqR9lDV1mC
97DtK/X7y//Buvo4fwtiyk55H/Wtf70tvMFSfJJcp+3ntl1geNpj3f47/ta98W6z
fSGyDoCGbz3I/ThKb7bvrv8l3Y7G2kpWvcrPT2nBOs2XuTG4fMuY7g8HD+Vwufgn
DLz7p8R8nmrl1RLqySyiCNU2B0HC1+gsWQbPa15Im3GO32Zbe/z2hmEqtdep3n3y
Asofh6T+QEPCnSxC4IVlS+ACbpuEVNDofTD8o2seJnyt5O6NYkOyLBSICx+Qpy2z
8lMhU1cRqKEjr9mbZ/arIGPYh2A+3LdmUVMIdenJH0ntmwV53Jxx+DDzNdjakxme
CCYIsYjupGmpOyF/rBopuozYnnDPtDIA2pU995ZoFjK8uwIj82eson5rPDAdN1Ir
vG1oTbcilqUSg5930o9nHIBdzrAfTMWkId6+/6Yiyk+56aJkrl/WL1Jx2sQhC76/
xNs7fujY5pm0PeshaXA1jddgdadTCq5sd/f+O7tBtdtfYRA1paHkFop3o1yfXtpx
OKMnOVhqUWAwI77KMYXU/JeCdt8HH6Xa5l2a9PNg9eTB942PQnGa7SeqG6j4OIT8
uFKtsLQuuCnJpblPB0RCLS79/S1Svyv4+yC9hS1B7i4toSmFhUTVC9G0BDN6VU2J
ZcQgP0rzUd22X6fZvlUJIiQuZ8gYZoASWn8/JPzuJwdj0FQPicmCi3xIgoAYgWpc
0Xd5rgjtAQoFVRwpeuTqLOPs4wUJcEaic7A+GN96IBq78TlEyJ1t/Yk8N1388PN6
/eGeBiXIlrhALOlQMMPLVgJ2J846zswHwoQwEoKTb/+cU7q/Zf9XAzE6V2OMDJG/
S22XR7E4DmUtVhxvdpR+ykvWeePxiXccdNvxJL+uxPR/n1IRJzRTtqklpNjkxs+Z
54+2B+yL1j44KtrZtczrdm4dxtIj/q4RyLSEKRJc6uQf9pRSXtXzb6/FvcSmjk7B
nIilLohd9Po1+R/OxX6a+negwqLCSk2M6BpGieLuQIoi1pmWQRamhukVfo44qds0
9maKd24KwtGqwzAK+1QKB2V6G5uTBZfSW3COFyjIMEXEQ2lszyg/R8R7T8W6shrF
0lHdphklZCXG+8FqD3V0gx4BtgXP7vmDdQkvpI5ubc4A3OJzR6/ch5o27HwQivSP
L6XrkYGR3pI8dn7Vs4PvNxZDu91bxvfwdWz+4dswo4s0yssBuoVNZWRZd9nllUHl
lyDiIMjfrHp9GiILeXBrGCX1J6G3PBSp9fA6G/IzCOrHXX7dJx0Dz8R67TNeDMh5
S+zCWGhZL/yojV/o/Wj5sbiRJ+R0HQF+F0B+Z4dZSHS7fV6qjYEQ6XIBGFoTWuiB
OnjvBXSjbdxTFJ+Z9UDC/Rz8aDXzAViwB/gZmJTvlBacdiHtsMm1WzTKDkyCtzTV
3x05nJyeImRn2WWOIZLiQkusiR4lhDunr7uU7fWbgWQbG81pnjuwZDgA+2mk2fPZ
TVtNbUU2lPJe2tiXtOoEjW0s344ykDGXdEi0LxtaJ0+Pk2Wqa2io/PBZWxOdO+7V
VJzJMjy6sROnwbTZk4MPw2OBjni6qwHUloQUAMjG6nYidmh05oBe/zXINHjP8a49
Wr/b3pGXWNJfjbsrs6iSPUwI17HX26gyD1Y0XFOjMFSfwJoR8TTEaws7Z8QnCTQz
RA1qvhtJK90Uem85S8YVnD36SDC8vJAAp/+0fVNxTf56rGQFSVw7WWtvVtwAXVO3
uByUidWmwY/wM+oF4Flx6vwRhqakKsuef/WBAEgy9TO6xs7oCgL7pdKJOBHXLAcK
iYUj/XL5DFaGmp+U/umJlSYWf4I2B8x9a/Ief2Lcd4aGd/uy3LomT5QsQ1VeAnXZ
gA0GC61sj+lgNdZB5Tncyz3Avg1scZ3avIKP+syaGZftUqYXupkpC1LR+2FeXFUU
2dlCU0x/q2vlpvWLk3xWTsw74oIDXKUPZ9+d9gEeL3R0b2Hc16AbfsWJTgwSQ7l9
FdZncenHL3DxxTi/9sbxzmzsGLSArSxdzY+cEtd9HdSnMf3ENlWIhYnZ4Llx4b6b
ak7bSbN83Ht0fE1i+oQ02a69fKH6LrSWmzNNTQLlMTfcl9kEpdyrwoSpk2wtE3ZJ
llwXr5xZF6IjvkHb4o2UXwHpsac5681LN/eN7vRRJUMEkzlMeG/uWAKDTVPIuAQw
bXg/DE+UtZB+jSeworsLqtKTIKLTbPy3puvqxi8tS/JwUIMnRLl45+XM8RPVXrVG
eQl4r7uENabqTCwgsr2xTxOqZxJjxcwXR1En0CZTa2PFeivuYoh+k57cfdRNFRWk
a8BVbW70WJKaEg7Bf/JZ4T19TTl110vVd/zu3u1I1lJYo4MktXq4AeWA0yAK3LxI
hrfrlFRgSrnSa8wXtDrx+ZgKKhnmtZcW2VQYywE12qBzF2sUA0d7ZKSbYOUuMgwu
FR/7mU7DP2aqZMvZGdGmfl+fSSK3N8rd1XYIcRYGp6VEvjGBtPteNQmznRdoQ4Ss
Tz66qwjGMyHB/sBE+jdZ4RUBA8RTPLOwctaQLvrbk9RvqJgAn7hKwWLLUH5MBSym
9iVyhQjn7IceHaXCsNUU5+dSvThlWBYPl0pLaF5l3R88EYkzje/txgX4jsxkUOcX
UvjIeHux3iHgQqVEwWSLG0UbEmMnQeLrihCaZ/OUYKzWGKGmUI2kzS7drMoLS7CM
LqNRK03mn09yofy30Z77poJy/UZJeyQHzi7jQPTO8r9r3ye3EwRzwdd6fCaOtpc1
DYIukb24sj7URuO2qDy58dCt9ywOMhklYqRgost7HIraIC8AlOdVLBXaP9TmiPu5
5/lCi/gJsdOx8vfUtevaiF/PUuGkjvJNrEKfh1LjIv6xActK3N6cjHB+yTK3o4tz
T8j7StMJgtb4LjgD/otGCTn8CPj+Mk6hPjBUOXd6aLjf4Gyiz+bJhJssE3UeJQeb
JzevH91PFXa7kpepCDgqQ2b7fBQm9NRg2eFQdDtITJjSmdz1eX8JsHxg0YKrcsYP
W2qp+ShW4AqR/q4jb7ZAHRhGJZcrPpF7HV8fJThd5RIPGMigqMKb+WY1kFPT0rac
HWmsM0Velmvtsh8VTcte/5ZGvZGvv8BdeqsM5bM35XXuwPb8mb0HE2l6YujLpsKX
idJIxZNHrd469kP0xncM5bII9n8TNFaaN3aZO+Qo6Gt6kwykyAoDBGPgMyajbLm3
TW6qBSzBSmRNxNNq/b2cVyHuVq3JqkxX8TMqeBnmlvAby8laTmPyZhbwKsT+MKSI
6NQN/UcQiZqjPsJU/kYi9BOX2gfN9PTpHQmz6OcF1xo+b3mUylWWbU+QEooWFP1a
2cujbPRvE7P3c7e6KCpa3Dp8sMtv23SvB/IKku1sFhlwJNjeIm3214xMP4q0zi0U
ECmdQJiKO4cw8VL+OWzgkgjktmhz8Mcgin8XWaOdw9chCFVcOw7qoAYdUWCR/4Zk
+K3QTq2aL2efWLbDYS63UokCQWtbLtxC/2UGyVS73mIQrzPH6vZFHRfUb1aduowv
tZZf3UhQ/FdFj39nb5sPAA3HhFpmGkKUNs1dVGNz19bh7MgApweq9eElddbkZuvq
XqAzhMvSuB8EconvxFMvepVRzMmbyO3rnEoTFvGIJyE64/EKXRJJIHeuAvAko1L5
1N1Kcp3t5+6K6S5r8GN8EiUnHsIqIiPpMb3ynHjACS4tn32N02lOvc1NXjK3tbQb
qRJk79PSqU5SSBxNj3x21uBOnqsg3lKB1lx31aHMySk+nHWmFz8yzMp/hey8vYPC
f15ZuE+aUiEY9op/KzNZMgOT9YNeDAnFCFeTuiKV1IQ9Sz7LAaJbvfJKVUHRAF4y
riAn5itkVhO2A0DB30NvI5Pxhbcatwoainsz8fhg95fLSMJv+ljf4maLKuA7qLmW
XeR1VPTOVvKvzLNQPoDNR4nuPolnzGNUuM+lKVGHf3JhXqKAbx/1M7xrwnCgZLWd
ApvNPqcVu6PD44g0r2hnHuaMc9mvi5WQ55lbCasnvUUMQLZWn7gnYQ0hUfhoFiab
xA+JpJjkKyL5nV9pfe1OxCtwCNJFqaWyaya75D3gcDeZ7fC91q+dt0uxq5rArWTe
KZeaTA3D/4mussVIoN3t5r8skKS8OpM7fwnh2pK4rKWiCPlCfHwucZr2Ny+OMxfG
pb1ajrXPiAqtczRaezzbP7+JJ+tBjDnDWHsb5m/hlMeW/c4RoTyBROuJnTyHnPh+
Zuavhl3gtXDWNXcFCKwnp1VPLJdkmAlYpJoMblX5c5+wu3M5UOy++P+YcBWeVd6v
ZGPzoD4DLvUto7RxhHlMVkJ42DwKp70NI8/6IkrYQr2IkePM894eDuuFtL6dbcK+
dbVT5elHKwCkKg2o4YQoYhmLg6D/zX1GQhOsBy4HnOzUMbW4o6Pyebwm4e4rTM1U
HtpcbteUYutG72YQeJ2g9mhxTvywurkN9elZJqD0a7ezguZWzeM6kAB6TX21okUQ
sLrje1Sg6zTTzcrpxj2+jY7ZKzox1soxSJwi7G0CmWTL+MiUDbqL6ZeqzoCYY/hJ
nb7K4PwIJUt+OxUDpvjNNggFzEWqxWjn4dMuXiF2dpx6EoVMpNxAidthRffX0Oph
VSjEKufgFztGm9XUPshanluUOxATKe+1B5y9nwnPVGc3ix821wrtNNw/q0M5bbEL
hXhwZ/MJbV+3QxVWxnioiB+xM5wmPGuJMAZfMrgzXV0fNhjpG7+KDIjNa/l0w2+q
8Y4UxadDQaYnr+/qMacuyc/qh4jaarPBpcxMvNl9L7edOLEgftFSk5uNrwWD3hSk
JFEInn3wbLoWOoR7pe2JrIKA031aLpEKLQRsOm7co92SuYQRU7RNyq98hE9y5+Sa
hL3thQUWO3Z12o/g8dAWLWzopDZY50zOVj5JYfUe4IvAegFwY3kAUGThK0t/xT8l
nwhkORmKBvTnEWIH7jdyMHcC2bOOS3KnW5ruqK5LRgFfuI2Laro0ZxKKeTr3cGZo
PYMJy8MADoD/3Hivg4nPURNDB/D4CrrG4yWk7CNu83U7Q5461gefF7PK1HCVoL7u
XWIGZXGbAS0nx7bkPonIM+riHFN6UVqnyjbjHb5Sn2oJsYuamN7umG/kEstXpLvn
RmVBRTx+zADW9ZgKdBigZlME+VVPVRMAX/EjUrK9oQ03EDNXzXYg07Jb8YF02mz8
IUc8zvpkE3MrWBx7uCJGDFak6dEScJidiZctO3+VQZWvgyHZGW3jxGo019CXlhXF
/11qlTy8k5kPrYJUYXl8HdnuVDvoMaqz52Znhkml2JUkuIROUM4NLqdb33QFWj43
eebkPnkRePirxQIRbEsCWEp5rBZHI+YHmIaQStT7Ih8DO5Q4ZaaurK2ESjhwXC+l
C0s0OA6N9Hxn8kh7IDnwJXGy0OPQ/GTx/Texca8De9nug3SyG2bXsH53GtXWaDmk
o311hLAA40TTboZ6YfSucEIltaR9bq3mregUWxEaaqu59tbOgGNrFDJ7Bg3WMfC3
4TApSt4jFOX6+zsXHvPho3s7PY1af/jZa71QNAWg9pdz9dz7lsbVeE6b4DyZKPnC
ayV5pShSHNt7x3IE3LX/V2JKPHIoBVS7B0AShv5DBoE6p/G1ngHgOtGecU1gZ6L4
Si+AOWdmWsDbwyeyb2ymgQ13g8zkX3mI1wtQFUhKYk3GahO5dXr7dh6eN9bIfI4Y
Jpw3pj5LAUm3jtt6Pgs4oopi0jXQn56AMMzUexI3bcE90dQu0jQ7DYi2ozv5Ecci
KFQGddpdzP244O1uHNArPcnQONs1vCMy06bXz+Fnu27nlOSAlxOum2WM7c2AW320
8egm/QoVKAjsXt35J21RZNiXHPEau3lsN8vA+H89xFcxEgnrSCb1Eaa1VPU6ezTO
2sqneQbkZoEDmpA636TFiEvSDZrIud0fg9CK9i6pSOhXtRIBZZLyNkJ9Wv2FzxtJ
iJOgE5rfzn056A2zqvS1MHH6wwvEYlFG6cQEmgV6ZYGKoPADNfwvU71QZfOlK7vQ
4Cpjan3Nr5h/Usbq/qenkV23vyvSFtBJ1QWDUQBjFyqcLfE5Rd1pfWu3IXk0Y7UW
d1h55fEwc1NPhNennTFd/YOLFcUTW/qouF7+rbxXUVYklQnQ/pAAtiqq4PGQAQ26
hcisUZDrwzaf6uRh6VIZRzgUbM1FZTQ4W9jMmfLuCVCdAweqKr4h8+JDWLCgvs77
9+6S+1YLpNvag+NfIHkY+OCiRJkJIPQFkiM5t+SYeS+DMXWNyooJJ7aXBBh+yqXp
h63xnNHqsxDcleT5EMn+iU7xXn95qsKEYnjwYfldovCUhwIKKJRjZPu2qHEZdx/B
3sborUz8EzQFk3Yi78VHdziKbV1xx7eOKO+yg+e1BPr20JWNA6RPMObOHTrrz1ak
aq0iWxcJ5fyJ2s2Gr1kAZwhvHYzDTzMr6LZbiC3/Pilxdmy3bGKjhHvOt4lIGKBD
ZitSKNkEtxn7wlB6ibJC73onIZxkb8FsDm/by4fPrTD9ORGMJ7IUu7/5daGFwrgX
Agv6UfIS0Liqt6uDZHTaZzd6ybs3pd2C9DmEcCJ3EOGyFHi+EOxXvmTJS7T3QZt+
HLHzbdc3nb1e2LDHs8j/OBOzu24suRX3nnBnN5Sh7Ihk8RxN0QM3M3d2pxgudjOw
kETezq5/TqdmdCcFXhkjHThJmZliOCt0LvzfrdJ7IdYFcAMw+uYj3thWyA54CatC
dQ6scCrr0ifLC4i1SdgPc5coYW4LOpgOSYREna7LGrAgY8I7TN+B6kzMBlFHsTB/
kvhcbFJu1u/AlPw3bhxzMM4uCiTGW5c20IS7G8qXTsw9QCds/qFFdY2CxpmCyIQg
hXO3Fd1pMWeXO1piOEi249yHIkSQ0JnRp3Lgmd/fa3eRCR+BOzBOpHveRlppc8nz
yu6a7jHyyFd8qxuRJwsfzhD1gEVVmguFeSEMjXYLCeCzo4oMpwCrpSqr+4Izrbup
8uhVxPFFc603ycyt76a6d6dn71vJkye7hdjTXVU5nauA+TMByEYRTGiBX8NGGlO7
xVCVtY+ICkhVxGDBTXMnOg0YyFTpec58Ex0QVKYdEUWa2Rrpx4TWmVNHDrR/BZmM
/IYUMVx2cHjIoYYxh9EWukFUKPoFyuS0izQ+RZgOqUagQ8ndAZrwJ2RD/wt5oXvS
kYHtp7SIKvcN4Tk9+sVjn9r9RmLaX4nPSEPg8Ir8ilD80upqvs4H0hEs5N7Xz7LS
CuYhT4ad21aCRFYc2worQvjkh+nxZP8LfSozmlC712Tkt51zwWeWuN8DwUM2a89Z
ThNqFWFtjjSglHyONPLEuOz4lBDAxBhkeLknvjn3wV6GjmUgmKvcLkxxCpU36Ugx
h1PGbpeh8PRn3V9zk78mViCqRCg65G9j442VMkGVdRe+hKzv5Mawenn2KxPddBif
QIP46A8cTdhbpbuAxX160r6hDh6ckFqXmDd4nPI5UtJAPUoT7Z6Fhy8fv1Q0z0dM
gShigwiAEjtAGzdlmq/s0XMuRTT/2UO64p4hBgxoBh8YrNZgkRx7oGwca4HfLWnc
GjWOw/Zb9tqyqpx3hOdzWK9wPyYcW9xaWFTeIHA9JUqdKWt70F7AYHlX8TNvr0wA
9svaf4tMEfPpAwlwkAW//Tn8qOsUx6NjuTKOTY8ruh5R4YakTTVJKygSFtlvQ1eq
W62WvDoYrhcF2X638d1Igz6XY/EoAj5tNToabXmF2LGY1iFmRRq4bLpvo8W4ud0O
nQCaeGef1tijYDVW24I3ZMNdf+0rOkQKIv616BMo+wbeRT6rwfr1JfDW4AveVUqU
AQu0nrJyNp/ZbMdCZGEFQHzAti+zbIpS8Z1+rUjshVZvCKsKLulJZWartInKa8KH
utX/3QtWn4Qa9C/iO8bKh9U7Q/z2e/ZU5rYCmGCWwR+M5/QfDAefcFKE8I5puHvG
/PufyhOK0Ct8CSBYSrjFmErfcwlcmxWUIHyrT/dgvYM7Ds0XXdpHIs977OvYGWLl
vZV9YBnZTgleWTErjvHwa4GDk1651KSsqZ84vGKNxVuN0xN12p7GOA1WmssOgbqn
O3bR2jHlT6qQB32+5i4vPKwcT2QJZJhDugD/w8/LsQiSU19w15f0dRFnL+K5ElSh
OtwzNUtfQ6X+OlOqJ+B10rbVQ41X4LwiZGdIaTldWbt1Tsk/YrDjFdWshrfeiuMC
+XTijFnRLAqBHMi6H3lD3c1vE0Pp2+S7E4pFVpvCfea7SdLrTPJmPJ9pGn3BFF0s
3HOTJEeeEo+/GY8ViljHbXBVdLLoTWgbNdFKOyfhNbLYQIRXmENW8dF1k7ZgA69Q
yCu+n3JS7fPni/83e3Wr1rOUQ1EGRoJl0LDL0yGUwNyjpA62aENmNNbXPc7Q5Ljg
p67CdyJMoRJ5u+MK0AtQafdK2dsQzjR/1zf5i7b2VQC1KyGPqebWijF+LMaGIWuW
vykOSO4hPpzTjSOjxADxmAYls19gkKzZQQ7M2471sigM4vLzId7ylhcYINsKAFlb
p1QOY9RDy5bZWorH6suIi088t5E2gIjzNqUSB9dO2J6EhlNYlQ067AG+9wY2fP3i
WslMKtE2ZqF+kRStwXczad38Rk5UJqApjYGxUwT0YKJft1T4cHE6uLm7yztkauGr
hR/uHQP8bQClUrIq+mRlivvVSBvB50oHpBco2QYR4Dt8XYHWGAgKu1Rm6dAQVAx1
JfwyvEhy5w518Tf6jNmKqIYn57eg2l6tCs+kT/0c3Ld/porR7/ivq+AAS9akxFJt
X9m83XOFosRd/cYlJGNPVKpelkW66w2euGfBNmAXMPkUxcWJgyfBs8bDGGrgk4Eu
fXnbprQPpL6p+dti1cl/FCICZyyVJUqf2kioIzBgJum5Psp6mLSuSVQvCtlujqXT
MumLkagiScT6kykWtY1aul/S1wTdCYf0MCEssPyYz88CXarRaiJGfp8f4G+RnaW0
VvMMHmJQqvMnYl4oImZDk31ydnR14LzuXOBciMc3KE4f7359TLd6XVrnCzJMhbC7
CpAPu3yZ4ZG2yD2u9DMC2xOKvcPrt5LDMuB7jsXNiNrbJ9+EUXKqKdTtc7YHj2Yx
u2pmA/f0YpJ6sxiNRn0PxW1bOtwhtewdUc6aSy6ITHNK5n+KThiz+qJBKON7M3UI
GBvBsblsVuyHaFuWW9hvTaJsAbhgesieYoDxS5rqp6IPLvPF7AkMGedIUm9LvzTy
W/B66OPQp3+Sb8wHm86PWIZc0JzNzUNSfYDDP4koJYo6/ipttTMnLcRY/rKrSwHp
MvU6WuHfLj/NF10qbxjWIpgp62COXmWEoS3IUAO2BolHUX5rEzdBTEya3eOnwhPL
MWpTk7xWiw8quU1YyHDkf3CXS6X1oW4BFnlAlz0aCGqK9K5SC9bwAnUpYiFFndkG
cDYxr9lsSAqXRFFtGnApKws0dn0kXDyf0MI1YRI1t3zpvt2O1zim6etdbsKU0nU2
1xZijErIvHyZWARvelQG/mrN9w55OoWIhh1zSW4UWK8hE9KUcRU4djGiA3vjslN9
/C4krW+9TM0dOdcq2Fiqq8d6bJXkTA63dcKdbgW77pvfTjZ4AakBlVum/NBXTHE8
04OS+hI8JBHSjyL5JLgSVjBf96ce7Vwg4CBYMtemVBccuRUC4vdVVcV5S3DJ+pUo
i0m6vmrquZYmgJpcm/9RlenL1jKala11gGdQFae4umUZgYUGcdp+Zi9C1ZaIymvD
9EYhqXWiL5r9ScQ7IlnZm359B0o5ncTibmO7QJAGwAmHZO1Lc2GQTWVREsCfmgmE
kM82Kq7MuVdF3Tv4gJg380yKrsyDgaptSlQVYtpOl0Tti6vE2s9Ar3ibaXwp32CN
818tuVMQyfTxvmScAx+N1F1KyasU/oB/GuXwYd6wI6Hk0MEKlR3hGU25proM2LOI
/8joKntXocG4p5NiEPoOgXfyqASyLgEtL7n/5YxEwUC4MR1cr5sNX2PSVEf4uMQG
NAJNfeiNd65ISppznSxLKDE+4DOY+QKloa8GVIca2mztmkS9sKbTEtiIr7Jq6/Tv
ahVu9l2FFKj/W3NNYQgyMAmMEETtlDfKN4L4Vs4ltE+2OPhHttGJBz70JHDiT/H6
j3mK//2fXS1LzO35cv4odlChu7ZXrA1Hk9EfDyst8ya6Fa5s1yvEDvGmaO5rLRtu
Dp58zWv3fxw9oGtFT0ehWnnuYPWot86HQ37y4oV8TLkfdF6si8yb4lTi5S/x3eXG
EIo5VQJh0j/lYquqUhHoK914nlkWBfeqMvIFC9gKg1gVxp2xct+P4g8pW2d1ZkAK
xhNOR/5MYOzyGAIzd/5XlYZ95EcFdZuMYPJYdIUzMkvldcR4hZDH4fR3U3V+wRza
D+2R7ZxrWHRUVEWMnO6KsUM9yogEClR/IIOlXvxREV2QHcI5k7K2ElfK/T2kVBlY
+S2FkspyuR+7NPxcTSWKq+ahOovLtYNEtvfDX+Wu5FLs5tdMurDQbPXhoNfBKv4K
blTHoXtS+rC6ZMbM1Vkn6BMfQZozgv3eEBTkTMaPpOqdRhcJq624NJJ/rrngu0Cc
wCenfxQcqvb6T9kv7O5uy1ZYw6hD3Z2FR/8HN6ZBZmwoUvVh+Mn3XA2sCMUXK1nD
2j1jSD9PVGqdnnm/ZMmZjwZyzjpza8QereKR7XVG1A5p5u5cNB00xX0EwdpeU/FV
IWF349IL2RKpMGWe3VQrs2pqw/6Cjh5o71WjPgCe1JUoVtIGBn7TPiLuEtk937Gf
K+Aue5Ml/SUC+tYV5iRPebE4nrSP8H/MpPs4ffOMLIuERctBrffqa0FIOIr+mapl
9mhZWbNMiBQUIj0RxKjTjN52kCaA9JtvIq3mAXqzpfM2F/0A2Cs99cL3Mn7fGJJY
B/wCgUYi2kv+XNnZ91vFGTHJzCsy4ZRqdPqhyS8p6PK1XkGVv4i0/AaH7bZN+2jn
7Qt+QRxMxFpMm3OrkIauY/8m/WBBiyE+OpPsEdqgzuOyyljgsCyay0I4hwG1EB1I
HKXvAUao0pgZQRZLyFj1RiSRaBw14I0zYa7xR61ve6Zr0A2ce6xkzowVafjzMUuw
EiqFlxs5WYPrK8x9JZmbXc3AZF9FvhbXLGFFPvD+UquWK2I5G1MzhVY3MofklOJA
lq9N0sERJDDcWt+OPSQDZnjmzNC4Q6C7R+ttWf76y/+K/UXP3MC/z0C43BPSO0lH
9ljUO2F2MRuwSOAU5OVIbTNIqqjUl6j85+mIDpe8MwGOZYCwf9EWG45IlX75HmTn
dqqU8YIWh3DlChN0gizhsllPCI8du954bUl5K1g5Z8Y7TY8RGBNyqZ2D4MOKTqLg
B535ZP2nFCPohGA8fyXNuLgjuVGJlVns5te1R6DbXRto5g7ZYzn8jAtRUXGJw7DC
hfcIl9qT1Q8o8YKyb3NQ/NOgkTxh1LEi5ckdvetAsKImQFpKiIJwt/L4ZHivI9aZ
AkjGrJM+EEszQgQmrXwxIGuFucEv2c+Csy7whT/A/M7kElA/+LACzdd6MDnJkzYc
EQ9yYr87HUPFH4P8nWEzMD0KRSOwLx2H+HLAtRTs5fcQE4YthkSxX9d+U9t/BxCI
tPEDOFhBB/3HlQK+zYsLiGPxJhNrjc2St9/2+sBYAZ0nbgD0S6n4IRm3bmQmSTX+
fsVcgwNjxD3/dcK+f9rGWmJQUpbPr+QIHKOQR1HAwopevWCPJrtuKUqfuO35hb/c
7UcSLdljIoecd2dCAlPQqSvrMxjN+A9lqGxE+TlwcK4LCGwOFS+3hR5bNmsuPota
lfScWG7vDsthca77yYgRePInlKN3sIBDp18N2c2JSC8UGNIGV3Yxrx4rc0PohMhj
mASSgafzjzf1cnWARmAK9GH3nA9TOcZWEEbOzZKwSF9CBjVOUdNaWcRSil2cQGkf
apLMMwIeUF8bX5S1hy3g7vg6pPIF1OfN604RWSwZT7irH1C6oGBB0xTnsTKFXazw
0JNgwMHdLiQewS+sgw4vfVP31GaGZmig8yc84gCVbKUMgPmMUYBY+xlFGbTZtQan
VTC2mY+zerATATEdN3mQYjg54We9Pg3bEAyofKQfjYLNtIdywYaSesVZkC/gvDFX
baQDDcwMtIW3q45m3QJcIOd0wRMO+dsFk4WKG+7m6xipj7MLwpCr4H474aYCbw0B
wPOPsuYmJ+oW4eNr1dTdXs8VBcNmbRdWAQrqmz0luEEdsUWhzJMa+9IRo+MeE0/h
vPblGFYtv6xCxAVrYSe6s7XyP/5JnFkdAqFCytCUbB7aezp+3NsaAc+x24CQjUqQ
mdutnXMu3brJtPw3tp8WESO62a+H0uqdk303GjgR/DQf7ubxBKsqK0U65AQdcBFb
VGpXSJ9c5opmDYEKOhkVP46jpy/no/2/5vgXz/C5LHQVFhOGN2O/v9x3re1CYnp3
AKTayctx1JW7UUCDrXgK4Py2WxQxhOD6qlGBy87go6KP2hPu7X0kSEnRua3Efl12
MsspLkOP1HFs0CbXLYhuUgl//WniS2cMvRKQLGc2vB3QyyQQOKbOIqRrVZToQsdO
nBb/ReFp02uhyQ+DUIQDWkG9u5o1WkY1iNH3PX2e6DoZRFuWadRRvVkGvGJrezE0
TZTM9j/KoH4mCSydD5pQzQCUNvP8ZCdpcc0hd0zTnkN7zuAuypnC/eDGeAeOpQjK
RFcK0JP0W7RKh6/14J3dSiDSj5nznhFS8WNTlWP+1s/UnD2ufDrXd0zfvqxRnwpC
PYwo3Sd+1lxpxlnzWT2LPM7bukiP8FJOvodpemTUE/Dw4sRPP46BU/25Rnfvl6pG
yf1KuNHaxtN0vqMC4jzUn0wPhq0bOYmL2F49GztLvem5I3k5sSOS0b+H2WTBFVnv
ha7FjcUayNteV76ubQO3PT0c180ZP+mNwPjTHWyih1rDoSg15tzet5aqEyCQ36Sd
nnn8mvCtIl7h8ElZkEIkOk+A7d/oiC/7jM2K7/PVrvKgrzZbpD6naRvnf1dDRRps
wu/ChV+KcI/bokVwwqJ2AHC98qwqep5QNVNEafGrhS0URSIasF3WjHNV39AThfFs
x3XK2myxTlBgzNbTyBivGJ/OntyApWAFpcXmrA04HxpmTwCswEin76PDxZCpPCNQ
WrML+VANLnVIx2esSzWAIg3MFdQb9/XSzhLBH2GwNYI9CNx98ndzb4Qq6A45uYrX
6paR7a7MJNcUrnvotyUgX4vJ7vM8CJ/lo6p1rOl75ViRRN9oodCKrkWm8mEG7Hp1
/47f1FC84lM3aizfgfWTo2r9YYkhGZxF3mreVxuO49BDyIuH2F0Uc0sPBxVWdBq/
48w7qgAqgPQmHLMSMDkFD5sIneLFiYefXOExzGhCQ5iXlVxOuHhgsn1WaBOmydBh
H+npRVqBux0ByoE36ofe63iruzE9K5AhLsBMV9Id4pUNLmqssa+Ual7zVAtD6VoQ
8z1Y2JK4h8ChXlg0hi8+HEObZaOyl6gklg5xGO3TJ5ipbYH9McAleQGeCwAMa9ZS
kBC6jrzdfYllrHd1hMj+YNLQ8Jl2iymrs7OwT4IHaxvDArQKpih7yUZH0VPjbc2S
TDU+501qa51Ya4mIFHVOa506TUe0sevGm0vIJCpCtyC4fBjTmXV/KJKH2oaG4CtB
UAa1zjrcpGGTRPVoiqDUZHTJbuOXw+jUpkKFAyC2Le+1XfJcYrHfJ3iqvXhVoxF7
Laksl2SS/XIRd5NggEH2O0W1qNgv/l2DGF8jRHHU43AfgpFP9x3cdTvDkCXvkxYX
GWexLyvBLcXQhZCb5SmMA9gGzr7d3HZ165mcN0ZGY1+s3IFOT4bECxbV9GDN+qaq
V1L8q14xPUnIg5RgMIn1i/jilevazQekpijIjtP6j+PYFMh8pI/3Q811wSnh/cNj
VsCUZks8EguLxoegD7EdriLKp3jQe2X4zpixtbW5JPtZ2MKxn3F8S2oYt9PcH64b
Z6vNhPl/1iyowGaFr/hfr3J4zDpvfOzG8Ox8kzqpzjRnHegwQ0+yIewHXDXewEQV
TcrRwq6j5gkezMc6rrrNo2d+4xlr48eaQk7EVmDnmjNMWc8VtHjcPvUO7A1uDdTd
ppFpB6KsHcrw43NZMQMQF6daprCRcJUTDgDZU2L51u4YDmfMMZzYYwFa1LMSl7ys
53MZGcEbRZDANMBB55hq2xGBOD4RgIFX5d3H4rjKZNEz5/snDI6/65XWllFha1T4
todewfSZxyK9x7wof0Cqd+G4wGFkyVKdr+MdjBonqU/wv3+GAUM4jFTRNE8BVPSt
J/vBsG5aW7zqAMc24/JQmmwxNVSdBYQMLu83tTtT0wjEDe1lh4mCB2alKy3zLDYm
mINhswtcFkemxXLvOSUikkdF8hl1phhjjsxKyC0XR/ktdobQqaaMM/VB6Z6uBZvG
YJKGWJUBcU2YxY+uopiU85uncKhcOnCqIkbJTN1SBcnszSsjZFJb89JxeQYudseE
kMdCifxu0qHFdJDAHnLAYBZ1euCNKZHEtmu7j/ikIdlkL+BCXjbjgGPydEp9XcSD
GmaHLzdnNAUmB143eJ61WSTazxYAKBLZ6YkQEBLccElJTvU37jwsG+jZOOb1wmgj
5Pp0eEmCl28IxW3PNWPiLuzS0wVxTxbw+h7y8ECYuQXN/itpz4LdXGOXSROdpcNX
cG/NHO/UY/uAF8SrNVnGUdOXc15BK259RpR2OXY91/3KUkO6koItmQUvI8pLxoST
sDruUPeDAkMtRLJz/Y97NCX4jJ7B24tMcgAKkDXQj/FPruPjKuLMvc80wmIlGoPQ
zKvlMUEJUMaBOJg7Kxi6YASNiYNBP9V24E0TVPJqRF1MxLs9p2pQrRMegE0G1sNW
1ACWh4TD0nmyut1tRE0eQ5RGnlcCciHBsjiw90zoimeGxxH4MsaHVqP701wcaLx0
tjY0x7IH6Y2pYkkeLrd9DUO3lAIdC/m9rgvy0rWK1xsZFR71WGnvLJIJw3vJ126n
9KPBkbfwjR13TLraazIzGssdjUvFEk3IeEfxGOE7lZp6dem7fCycI7nq+fRFB77X
SP69nBF5D9xVcrlFpqmykVoDGNHVTWCpti4rqZOVMrWuhzzHixVyc7+8DyAsHP56
EIgijUSCWbVMNSBW/nDz41gj96ut14I5RpVNCqkrpHa2yuQRgVqFUxLuCvVeJbk1
VMpPDme4TKzZkWR3yWlHvLSPWVGf3oKEsqxXNFCpntBZkZ4ST7t/jr4/irV/F84r
aQPhwt+oQA2+R3RQMFetdB9ecrQ5QrVgiAs8A9+ekymmYFPVy8KsikqPZGgAwr+i
3lsIHETIUKb7c+rA8geKoU0ruf8Fr13jX5jtM/j23LH2evE7lNOK/4uCpM9IuyGC
1Vg9l7T8f1dAcKXDOfP0ao/bAAxmA4WudeCj5QhIrGI9nWxM7XFdtoGMdlBn3rYE
1t8P4CGjVIu6raOvNGiKa0lM6hjfiuqQt38izJJQjhiqJ51n+xtonA/OXprFIQGy
Qc8+OdXsz5wJ6iwt/oxA4eo2llNpTYzoQCkzY+E8qEYtKlXm27XKsGbVDEt0fqJ6
IeVv8iDkDVSTsXkhL1c5Uqws8DIu88R88D9fJniaRZMwZCZd5Z/IPErOlBWgB/R8
G/IF6dtSQZ4CjsOgRQQ9BoSf5n2fJ/03kwpzzI4bK01RaRBw+RcgVC1rewSuQesS
dFtd58FeF9N8xexYc32Z0J3JpuuUO/10/WOrQcTw4pLSeOIQyzETlLED9yYQp02j
pVQkpfoVL/Me8tz7siiiRNytSXS67w7GCRsAY0iKN8+9Gx6CS9DUAz5w9y51hdC0
kQLD/X/7KqdATZtdCaGgF3jpc1PlgfLk1ZfNYf/UBbANScTvlatSSrTsADoTE2I6
/oI9z9rZEs1YvLdHunL82As+vn3vlleBwEzpEqo6pUoJBCxctCeC8/61jtjRk8ZC
ch80tWa6fK8iUigNIJLVALUN0EgNeYBuJ3tK68glCRfSdkdjvLPs74XkA14Umglv
04z23YKljXPv6jFFOGpxXXg1IqFZCU5eraszTbgHazbWwKmNnJny5tnECNrwDH2J
tQypgfnUMlo0Oyu9V+z6QyEYPJ1pegspd+M2EmBfScS1bVb0GgIYKqPnlpDxWaod
PBugKvVHGL/6TE1u1ca1gDZc7VJ2/kGqDzyZEMRYiu6UtpnYGYaaILeR/7UhxpOc
TfH5oI44pnC0Q/miLL3TiDMuXkbF63eOpP20Rd1mfvN+YyrqtcM19ADzzThKMIzA
7LqmM2Iamhw35oDVcoz7DhcuppEt1lkNvLBpQL64JOKBUjb9vFbzhT6IcwUXujjW
G/fGuo37VI7JrfVda+sj2nMlOwYrUd8MwcjvY9a0b5jj1PFQunT3VcCyXwUOBm3U
R8hIr27w/9pq+7JGvRfsIYhES/7xq2JMxujT4qfXaAsA5puoLb7k5BLsxf/u1YN+
CWlhPYuAqU0OKmYcYhkIYMn/kNbhVZOLbODa6CwOpEmQoxxS36L9MYh3gFaHApt9
WFsm0WH9kXdeOodS57cvlL7cEdHjT/HTSAulByF/3ir9Vk3mMrZ2lLkh6QOfVXj+
fDQd5L57Man2ZjsmMx2B+80hTQ85ddj3NIkhR7wzNfENDiVS1cEq4hWokQVuRl19
jZD3g1hnkysFiX4dYs+rbTXq7OIxtDs9omuhU6Qe4JOUHN/SMoQNZtzUQ0+p3v2h
T50wt02rhQ6OaFE9Rx3H9JH4o7NHC1RmDSBwAonc5g8iRjyWjj7dEFK0uUIB3vfQ
YRTVAaXwRlgkeaEgJFiVUIGQGtbk4pa8sFyBjQIsVmCO2VRKwn8SRWbVPnx4Wbql
FPlG/m3Gn7P1URXLUNlm2ojeHrXKydW6AUCmCLHubz+jDk1E3XNCtyFsPZR9TaSF
zB1/QpgOLukPlhZw+4hlF6FYWwIJwoQRV1GKP1yiD0S71wkrzXTnpREMycCNRuT0
ELDyZFazeoi1tZzKO7DBypnVUFrs+5GRSM9qmvYKqCOF8Kvb/3dCcaByhPhg2Th9
iOYzR3JKTu414AYLMtXxuUhsJA9Ay1FxAakLxk9PpWVPpyqQxioSB4wO7aU1uhqG
6CT7MnpweHmtKPXWDR+J12Kz0Dz26Kf+ctbp9SjAKA76CBv1IHJjjlZsO1eZypFq
DoXxRcZjFypIf1PXfnhxwsPZXdAuuG6aFIREL1es2GEZIy4VwWerYZgqRiC59San
o6GhY4xEUJofyMoo93tSd2FcP5N/oBzijWorFz1nWCrmdVBxF2UEFpc25LtSF0bD
3mSjZeUTKaVb5oFhTo7euS/ZKL+SVPwEAZuJLMPBKiW5aIQkzeHIatpwtGoStuuF
UvJNetn173MQAQxvEl9M4Z/qO4Ozq5grz0hhGzj0q/UJR6cQKAZ7wvzRj5Y0wzOg
tsIyd1jrZMc4VeXINiZy0t37u9im8IqHrRJI6XSCxL0FGymiygRPxNKLh+HSnnJ2
pr5f8Bacy5O1EbUgsITvRP46qkUldsyyqiYpZNAwu9FxcFKu0aGZbXNHDyYxYIn1
ZODcY5gzwI5HOmX8bhb39SiI18d/W71lMBfvfEL7D7GXllUgOZK9bMmdfGNhSwhH
IVmADHcj1mVXLgMQuERZ3djhDOhhRY7ZIn4S5fx1JlMEHw2pYQitZxRNcsJFclXC
83w4aA9Fvm12zwT0sokaSdor/pF4BDVbVIQE57aftDsvC5iTtE8s70hkJFxZ7Br/
3uANsGwtWNP1uiHcl2cukKkmWjEiN2kKWuBvA6/NA856ipgVuIQ2azVRjGSDriLz
gVu8tmKhy2dlAgoy1yelKk+Yh8SxRqKjJmVAjfMAt8M453VXP0dCBOA454/6oBDN
KQm9be7esKZgYJYKHQemQ5ZXUFNyO7lalHps2lTNOFnWYN5yXYr+lIRE+QI98q57
43ZUD1/lPaCPWIYnS4BRLbXJvgh/xw3bpPZzENoapaCqV/PTrmiQCwk1MbTsIXzE
nHnWXbFQ56L5oySLAsNod9x+GKOJ2DRDD47vdnC4pTHQFZBPJrjXwrrIPwb7QVAY
DZqGHY3glyTqgD5XQfH3pO99Y1YRbhtVkunARKa0bWMrt/nYjwFEqtXuDnQa7Awz
1mucFsDYlCO+RPjMSQ4ReWXK2ru12+Wh7nQKCMGrptGe5wOpGMT6/MH2OeKhdvfz
Lvv3Kv/2LT3tQw7Ee19UfoSq4zduCxlv9/AG3Y/8Konh+0XWVTCtYnABpeo5sNsY
Oj7kPHj7TpQkBhl+F1cHqrTKumV7A7o1lmhvYxavH6mVXxUZxq4+mspNsUig9wnJ
BpZC+XemFYpkuEzgVGtfRB6cjkUgUjM9/z2l2QtRlJ0zXeLC7K2tgjTwtqkmViIB
lCtXkDe9V9LeYh0NkYyM33QrW6HbapvLadqn3p199GAG2qn0QMOpFchgT2cFIPBr
dV3vnmBPRzEdficOroFn4meSqmNdoBipC6Dn2CEOU9MXverMhIzDMyWpGReYx2mn
jUnt38PkmOs3vBHZmjq7osIk7CFvHW5fCDPNSFRl4HsesPFXqHPmFhAVHGOLPYs1
4q0bLBSGoHHEat39s9Zoa5BB9n8MPf0DjGX22efARpHoknccUG78gJY+xl92TWIy
1bb35Mm+rpaBwmVYU17mbhjwHEpsGafr4OOPH5hujJW4JM7lqsZygd34sIiq8i9t
7JpaKqS49aGYhPUNZZzagDATpBjbzAGrlI99mGYyy0Vx0HPqqmwCuVSr5xCSQBwS
bM+32vYmvtjL/fyrDEobm4gtsYKujyAfAD3vXyhKIBuclavkBZ4xRUes1cmMC1YO
PNFtiy+rYucX6xCfI8f3qlxQpXjY6zcvInejJ5I0buCg9B6bgG12MPNeC3SwylwB
9E1YAMxnLJ9W7rIMZGyXL3WL+XaY7OnEVvU5mW4Ha0cqAu+nHp1QopPMyRxc3Hh6
2bIaB108zTeTqxCFHMASkSsLyi/bw7CgIhO8CQVTE2mFAdLeTh2JjOQQjk9HHMqq
MwCuzivn9uSk26iAh/OQRGC/3ZCOqM0U45ZQZw3MUw6SBe2cbSJ7AAlIxzkUEEIC
LZCQdlVqUbu+TkQ7oCbZMVx77COdrgZDeOWAXZEcRVHGPhMFxQwW0or7PaX0l5GU
VoJdEvYh0GYOcCjT2gxEK+rRFSGUxzGIOPpegpMKumI7HHtVViNprxyZIopdsasu
0iXUe8dp2ISFizKzNNDcbfdT0ETbu4OETADJAB2/A3NhTQpPoJZhVj/dCJQTL9zt
u3eOf1QAPbDFvMbGrHC63yQJwn2gNxxz7P8IsoHIe265xlfdmMk6BOBriaHc2pBY
7Px60JaH1EzsgGUQUQHq57g/4zEJ0pfioGjOnjTqwbGGyxHj3TkiHz64lGFCnMTq
JqKfDSXTg9Z2Dh6d/lfib7W9lwM/I6f8SFyl5igrUx7Tks+mOqbRWhN0Q99l+iHf
N+rYSIZAl91N+eIMyTLRYNmhMBuAwnImAKF1oxo9zPUyiGmUdLHjHHW5zJIwlf8V
+osxjZoOMZb4tsc1r8TsF5jWMsvipMKlQRidxpAo7NKl9x7okhGZEBzysEn4CNLl
3VOECiIb2ClQddtJy6X+nCgJtumbq9+gPraQxsV17K2pZmqYYVtMOmVkldAxU+ml
tanBU43AyUr9sD6g2KA8T7DTXOx+cNCQn1w8QMff/14zsncrzVacCDHGkTWkwkqH
B9f53Q7JlQ5bKgTTBsEkGPaxcqpZCIhyskCcD9oq65NdjhxnKdZMpoTYDPcloVpp
Nq+7k/my19BdcixPNyLW9hfQUsOjyJ/ApU80I1SwjVvyISU++vd8NS0SIdgPjn0I
a8/uISdWNUBdBknHE19sjD6L1errBKUqWsP17Za9wc5sd7oqaRx35HGuMJCmfR1t
KtmqO/iBCrz//WjfBPsVmRhZoWD34QsSTpXrLjuTSBhjCatZSyo5j04/WYWWYZAw
p5Gbj7PY7etRpM0166jrX1wHAq8dyv70QFz4Cx0igaNYhsGygY5DaUpDTJgV3N/f
Wh6ivCcDDFqY/90KNUzrJDModr2mIS14mt0FgUrnUWAkT1vbbRzIcGqxomK64tVK
4nwkJNfr+bEfKN3bMJsAQxtihorCnpjZ2IMFsLU3+97YN0AWx3gD6BgW+ht7/93k
HcSfLn4BBiGEHsKqlzdOaKmSFAP5JgMomXda1SzKVSPibjDrVaPl1Vw+twJp/ZRp
487kdh90yhFxywOuY1g6Eid6t2tGEQRjHmZnaPVUmQuI3LoOXprUseM4sKe4WzXH
g0V4+XK+NWOHROwfUb6WAxLiFfA7qxrCZxn/YeVlRDsKmojInxgHXcWf6MlRVreP
tbjKaQSjkfFKzypTGne6qC+uPTPyhCR47oQxUMsPphKjdnfaZdjD0+0gXduDcfEC
Tjfl0pe404qC657v51gxryAO0pLX0peZqJmHQQ08aQGi7/cWdwQqDz6GX2mGiOVq
TeiFP8iNf3b4t7vwK0ECt1OvbaBnXGabmU8m/TNGf8bHkellp0X24eiLlXHqvWx+
z/xR2XHmS+5wLB3rRO2tKk+vO63v+sk296guVlNE47zKnZ8uQ5xV6ERmxruO/9xU
enjw2hwam9V0cpNF6Q348Vd5n0ZaQWFj+yvzC6PXT3S/C6HcCPo2pucg8pjLVWLE
XyL1aQv/nh6vME5hanpRmL70yOcF4lHyHeG4ptJEiSoM6hITzpVUunKt1GgoJIa4
DGaPPIIu0m1RMHPLNvkX+jfGWrS0gkHG/ch2AUBSxP+W2AVGPZlzCv8ykUjfO8P7
8IwHC3xHmOz3hJcRWFnMB3SbPDzEDS9ldGKK0o8e3sUfFiaKHsOZmr1C+l6lASYL
lAzjYiUseWOX3MSSl4kCx3/ird3bOewMcbxUcUYH1Z5lcx9YDaevpake5hc7f7tp
kM9CJRTc2E0pULdwilCfp0HJ6dEkyadQuJ2TJbRxOInoVUhcwusTuEWExHqXRMGR
VdycWf38e92X89jQmnfSBeY5Rbg8gdSM2ckpxMSnEErN5sW5tyme/2dZ8dbgSwJT
3asbEdScZjWpk75a/Ky0wo4bC5GtikIaCecXLBSD/VCuL/L2OoonMLTNL/CC24cM
0C7ANsuTPNcnvcvWOdSp0uNedM59i+47MTa0Sj+tw9VN7NxNwpF71oCFWIhoXtjm
FjHceq+Yn0m6vy/Ns/F1SvW0efIk7/V99p26pUFtCR4hIJUoPbbqo7wI25BQQOYM
gawjDsZ/+qceczNEpCCbAzJVyzPPAqHLKrpHx/BDvwks4ycvFXvnQoMMAgauU/q5
y/vosOKxpJU/cSk0pkkj3NsPPE6QHjPpke+YZIJ9WIkbTCsbm7i8UcUP2v+vDuDm
zB4TS5wp+3W73LKZ3xYAyPRjS5IdjVVsLN+O3DD5C1kC0d++UeUZJd6iERHX0h43
U4EQQZZ2LuMDcibJZ93GPot121O+4xWxipIR1yvxCWItbp7++im88c92IyVQS73+
ub8q0S9HTr8B7iWTX5xXqmiuqtdIYKJ+0oMCuAFheUBivkwrbzq52Mv8uuWR+E4o
w4vII8fo65vjb6zUsNQ0qZ6wXv/TCrHJfVL3kb+kym/wxF29o1SPgRrZbNj9btGN
7H9OYbgtc1Pp0nffixWE3SCZOVVmixMCpMZQjAQqmksWZCnAThhtES0Qo23OqQOf
Riu19qRUy6zgnE6bK/rx0aO3NAnLPAjgQceOZq9znsv0omg1iN1uUr3L4nBUgF9f
7fe4nNbebWr4yAmOGVl/7WoIYKn+rLAACtvbqC7wlmmuZQjV50LGoIYXDxOJN/NV
uB9hS0ALGBagAxsVuZJbW9NglcXuCHxh4oyaYogE6BWS+Ty4W3bawDpmW0nv/Ctf
QtB5YXMuceO84q+XrWgSNFkYv76qLlUcuVVGJx52m9aYicLs8NDyEqm2TvaEIe/c
w7+rQbofP0WLy0Mle+bTCg1tnH1IXHlGGWMSfvFXqyc31D0/7XRMMDjlYZxUzuYt
apSBQBNZ05tm4PgEZBcG7ySxMDJ9hSxZQHv+/c6uf8bAL63kHqEYbdoGwRHj5C9R
dinnAyxprRomJu41owNZ3sOa+7pOLZ0s183fOJuXi6QEaq5S9XdDDq3G3FLd5a8N
n4+ggZBZViu+WiW4JyoTW6Pmekav6lSuoDYrvCF5qVAmVOsyU/PvE7RL+C77Baw2
vgOmDzMHtyrxP8YoZPxv+h+tczlwCYOrZtWttjxYK78ylV2ZFecDyH+Bs8nZ0DwP
MHidPTC1/7Ph42Mubgsw47KZaKHQBB+lJpsjRWIFMQpfFFVL8Bn56+tgFSIPeWy6
YUAnP9xOqKUeJX7bFWZN0coL0QI3vTxUcPUhuzdMwcqOcLCyyxicVm/cmSmjTFcF
h+8SMu0REi3uqXM6tMUNTV0nXm2/Tl5nLopduLVo3svn8YwzhfvEkPFOUitW7+ww
20Qwmx/wrgVuTaJVg8Ibgd6m8UYSBnAIJ0nKylLWlInfOE8r5I3RFDH0+3bG0Dg2
VQ7ODM3evC1X6EuwkPnDZOMah3cx0KeAu2IVHUnhLo1xtSMbMxlCGj2roHz/3clM
v5usSviGQ1htLYDBtcUziKniqv5C8YBkoOaQoobVog7SMbV9fb1QjzewtOMZD9QG
piyW6vEabpbl+XMdZtDxOIlwfNcm4RyJrPxac0bqXHyNuGVGycA/YIHUwkG/c3Ma
X9JNp3TSbupre17wASsFbsO3vGyR6khzeLyOMs3OTJd8jJ0l7eqoaSFecpc5scXr
OKcB/F1/nCL1KCC2d+EyXaSFqRRuHTGXjjsvUuBclgw7qJriMooXR7G0eHxMU3oD
XI1yvRH6Tf9kCOXL93b78pjfd+w9IO25JJmqbn+/zwcX2F9344z4S6RwEsmjTrQq
tr64tFFZyC/CRpLhhTiVtpPB/Dwt6xXuvBIoViSpZS8CsSRT6aaLMLqz9a3hM+1N
re9cYlYr0+is0t0F325BkJDbU2ao1catiS7p/mw3E0ktx4+RwIOhtB3di6nqa9vv
dPXzIgoaQLxS+HPqIgP4Ax2C4XKf+iXVXHT4MFUlC6QgG5/DQSexNAXY4C3PRVbM
Iqeeb7DtB2HTqYaADzi3TXib8WZRIdFLUKwTSD9ck2a6uDA+Bb+Oiy3m43lp6vTo
GtIaYKbtjpbdaTVG5ZRwKlIhFb/m2ad7kbGZpU5gNjvd6unyscsmhfI8+u8cd/rT
konTnVAQf9PJLL7yTwMfTSlSNm25WxYqrZ8Xmf83Gf3FnWmMv53rio+RW6AMiODf
2z4ReVng2Gz5TbpAfO0qhfFlZaDjfsazCvwDq9habrzZz5Od5XD0JYFBZBJ32UnS
uf2172kz+S/fXLypip9TYvOM1un4pOYk8CBpzFuUy5r2zAI1BB705oZdhCMmQy0b
09FE9Int1idjdgZ5hycWHmbUCmxF3OFiCXA2rG1RP9is6gXMd3Oa2ta6V7/pgzXZ
vwHMKC2XCPKMv7jEBdsT8blWlX8P3DvgL81J8nyFnVtTgHUkllA0JfdIeBHCGIgP
SZJNXMczhwP14NEOJIYlL7vdCvzfVnS6TR5X2OCqEC7TiFyPSkCTrO1h7ppA/8Tx
5LmZK3Pwvm4VYnukKDik+UJY8a/+uRowmrhgZT0fg6Qd7oWwWPrktTdv7Da4fQug
Hh4AZGRUyFzSdsS/cQUmPZWldpi8twsK/4uqVbjnMZEj47wkC05UqDijyHV2+fCW
6Xm/lg4aEOHr4Ce4rCu+Y4+VVXu0iLTgDHWf5PsiAqHZqk2lgPhYul5M8hqhMCPt
qohu+11ifvK0cL9VTCB3ibiBpA3VA0iJPd8rqecKvgU6EAx/EWLgmW6MWTcG+AI+
DJHMioouaMw1d7LZl5h+i24plNR8r6cOgeHj9/E77vhJIY563GXiXjiHo+fMRdoR
XWTvm/IOAmyfZz65K3RtRSzWL1rp0fnt0RP0+c1ylhauxSpiAP3Ni04j1owIFEIM
xFXhbb/6Mhgp4hLYdHHbC6UAnXGGeYjDaQOokwn+6gFXyl2M38gGSre9Vjx8TiyE
D5QRP6tcu/nfScHkKMzgghyEgQoeikaofyD0HbZuSNIj0MjahvX/GwSE0qDZVh1L
j/pGHIjchFspINYaJvFuljYslkpewKNGxb7MF3SyeCW2+QEzZqTiZ8pSxo6l4I4M
7Ba+61GAEZkSe+2ZaPhU+5IIZnLma8DQzIOKJ4M7QoS70I3CEJU0Jh+rvgE5oizW
0xlKowztfp8+DaK+b9WBnbyK0cfr9d8Z0Ek9evXCIK2SfECh+E8I1yvJ1mcZiEvZ
xFq7BkWaRWuc4vP+1YNbDUBZYdbZwATfk6h+cgCS3MrCrMxV7wiLxPmkdpzsMzOw
7+lgRXW/3vHAWMQW/w28+jM7aq+ziWtWgm3nyxEuEz2U1bpIPv7PYDvWR4Jpm+ko
ZluDY8ofGuukZVaT2dwF9xPj6RkOCmhDsfKnD5b6sPz0UxCo1X/qMoadJu6MCYS8
rUCJPLuPPERzBqskSXzI+1XIwpL21+Tj5PZh5o+MgQNto9O0DI+mKZpBN8/2hEin
p8WWObw5/84X679rWoJ1zYrSuZzfJROAnE3GBa+VBHddePrgb+WsV5l0hjDJniw5
LcD5w6OoKy2u2eW6ql8vuzPncV+xtb11KuIFPXI250vx6cPx9rEE9Kn3kDcDEt1Q
+kK4vvSvZ9lQRtcv7iP991sQq4m271OUH9Y18NgfpcPfH7L+5FCWG20eINP3AHon
kV6nR59HHMIIb6IVXpSFeiILpTUb49kXUK/kZGwMlMbpCKnooYWnOdzmUiXgHVXj
sc80FMKMkGwIjLbALkIh65RVpX7zOCLU2YojYYG74Wbl7DlnuVweaMHL+K4znxyr
zteN8ECq2ZUo6B92Hktv+SV6KPmzki5g2uKZ0+AMuSqKyMFVLN2efeGfl2xrbize
SINJqoY8fFmTylutEZi0Joi4H4yeaf/w/XME9OyzWsvCUu4l3jYfmAwsr+z0k/M0
t/M8R3aPbFJNfaZy4pkj1/Lz7CwZb4dmqsq3dtIpuXrgCpQo+PJMhNsOdZ5Jl97z
C+tsKLkPMkXkopbvVkKE//D3G1l7asOKApVgbwjaE/lYWxlBw5I83lOELlltc1Ij
RC1JXVH/T1+LY9aBDU/klQutQkxrYz4plyhvRMJTYjT6KWFBOjOSY+okE5CzYA/K
xnjsc8m4VbEJd+ccQbW1fNvEy36NLHVJquFUJLyhfsNKbY5fuWJhboSqa7SbUW83
H9wSrIvvnu8wkIUE771im8jhvwP1LIML7pV7ALrR8dHck5c1/nIZKIxSCwpNT3BO
/+CKdxNZ7RrewjEnNzH7ekQQAhf7qNSXdExDi2ShE3oMrEVvmQY54M2N7Tn7oMh9
dcSr+F1j63WzVV1gni1NkZghE4KoitWpJCHaRyvr/WhEFA2FxxOqfOrDoCvb18e9
3sE7YY3NN9ZXJkWeiwRzc4jtKUMW8ULbOSg2QDCqjpOcKm8zUS1bVz3ttrQtZMQm
LFOvk+p1yM3Mgkrw/5BiUP23buVCeIYTNvKVvm4VMaXC/37RW30DiW20x/roPjAZ
5AMYgs6cW+SaptwVH+5jiPaLXGXtryz9bTfnPSi+utFDVqCnSugilNul+YeG42uQ
cRGS32o5FPkJMExCwqrTSZ6jlFCRButnsTlsimDD1Y3A9DyxJ6y7inE8B9yYijSo
wFHSYJZzohwOqP0Yj0F1z3tv30vEsd79xNG2fOaQqzuvjbyoCOcdMDgmncUCi3TB
XYRKl2OKwux7/FoaQE4nOStJOrr5WQFmcOyjgH2bMFs5Bj7rN4lRcwF82I3oXvD4
6GQRm4JCc06P3N8nIdgdS0Mm9ZxPo+ZngehuGpSQ0jmQmdEoeYWrQv3qsC0lbE6T
LySdQuQ7+iyJrA+k91SeE3RzsuXdYKZc3kyIxunugt9JOAAZN9bdakdRY7Zy3dtd
SKOu85rKAS/7n1RImiN0AKWyXMg3wqny7zGza1KKtyvUl29bvceVdqf3t1EvaDCq
nUJesXTXGX7s8+mOZJspC0tcEPWSFbBgXjPJg/4zdUNQ7xtNhZ4eKQx6QEa6wpkb
nJlSjn5nVAQ4hWY/TmNsNhtTjupMoZ8SwZzf4/nrdFC8DTwJkkMKbO89skBH0qJP
KJK6dUrkm5+kPgJo1GhksTvZA3RDX89WZdjIN46XP0j5fMnr87ms1+GDajQ7QRlZ
YnL50rS9OIfRaIE7y/5vDGMLtNcIOSoE34c0vlVImxN21piFBp0pSkECn7o98ZLn
syj9ed6DrOBatVylUUZiJKst45aPjtRwMr5px1xNNGBnEbQtjfbLebSe6bDtdsyR
9hbny1LDzQBgrSNbw+4W2z6VEN6VGN98GPVEr5YhGhywhcv9SB8Ph8rdNJYvbxzJ
nOxgtirpQyx0AelPRpasDJLCg7lITu7VQSoFk9sGWa5EbPBhIwEdRnFW8YzL8VeR
pbN/KU1TYYIrCreJDiVxCUmPlNkhlxTfKWKjwGAzLpKWl2TBT+HulegeOWvTub1d
OFM+LdXSabAeVwkr0ri1RZVNOLRLFuKtlgNCCksN+DvNL/0e0ytRiwdLxjYpBEla
46ifZlmtEcF8IKb9UsWGL2eJj12Y9Vqm3lJKX9zrmHIljmkKtPAJl/S1isrKShSL
Gj5Eh6tsuCA7iENsjo/Y5fVsyrED0ERDneNqQ3Fx1Cqr+wISZmHUqcF4rKNTXp5c
ptzHRRkzY0kq4rXM6Eqf9cAFcQxT9AWTvllKUfa2A+9+VBsIVCRoR0ZvkW8FXU76
9pzIo6dIw+g2Kx3j+YWtQJKVLUFsShV5l2V4mFLS3Qp/SxLmQuHQh0lvSZSq0nRv
j5hjXTCGq23pU43mw/yt5Gu6ne4YcQUqKabJJztQoCjSuuFLfqcjYifN2ersP+qm
fUacErlAnylovD5Vc8CqmtP/zzfB/tQqPb7hWZxRYzy9DTZYeCBljEpBe4SpUepm
5lzpbLIK35PyB3sjFsAKrSyVsQY7UYgU8LRZmH51i1M23un0+xpyRpHUfTsP54+k
7H5bsaCZAaWs1cDjMEPcIaGQ7IXm8ZQnoXO0IxkQ9l12mbINsKz/VudMUbVIqVBj
XmDJ4blsdGcFbKYCA9MjkZlOGh8ARJqPVFY7vBYu5M24PSoSg9ZnsQgreinkUdTX
w+uD5rottd8z3QeSnemslRFkmkvCVF/+7Xl6N1r9xb4N4vsRBmdKc1GFlHEL22ok
dquBlaL11VdQ3prPXetfMCqvFBEJshbWkmjlLjmq1pO+yWozigLIvdFqmvT6yWxz
RoncUO1TTL8I+d/hCch3+QiqGV8b7ot0WgNerNS0T+Rq1GXNDPSNDFarQ2jGhmhO
hFu5wKtCIElk24g2m8cSvKCiVmL+gm6M3nBRvN/OlbJc6J+8DHmRI1hyhdhd7Bb6
UB5dpy5RRe+UlRfvjhCROjovDsMIdZvXSxmnMLcKhXehWOQ1sUTJnOJIjMV6Qgu2
2JuyKtsuXMSqoMsGxg/2+gEdZgAoiil8Scb7WvDQQ63zViSVd71lzNwx1XpehXeP
PuCUDVoXcTjxTjj6dY3oZ4tBaJ9SQcivY3zDXYr3PZHOWsjomZdM20zTP2HxdVpO
vL9a5hlvIiRl3T0eHTc0UPsbK3zyCTsqQa6rpZFVMvSWe6ghA2hetsItmBqdeeak
1/WqSqHgmEYXCJp64GOVKYc8cbCHCXf//kfbS4sehLyy4QoHiio/wFXRrYHqWP4J
AiScUgFs0j2XCmr8xvgU2ExBjBRLIqs9gyzSODdnGUwylwC/AjOuSLFClDcMO7t4
4uAnltHZtjpw8pWDiuAKe7+lk8QTJqVsArCqNgzqAjiczjMXyNGpC92ZHPuMUWj9
1jDFXUhGOIvNIZj4L1tMwrNTiAaD+kzlB0a8aBe210EjMAcMLXD+3xZHZeOUVpsi
0ikAbp+LtELCV3iI9RbCKIUcqT9uC923+IGEhhDp13s9FTvz3ZBQrnHYY/0muX5O
4zAyKMs/cEqGWadNBXNl5sqitwsVIihlFruDUP3NAjla4ULECoZ5x4CiRv1e8f0Z
bKKa3xCYUxWk/bgrV+cm1PlLRTTPyms/Cagp7GKRWyPiLUsGLS+e7DTn6fcAIcaH
4T3Ng/b4YfW2GujBp2lrJzAFjSwYKEpwMkM6TOd6O05hC0yM09p2sGsrcTr1gFbg
DWlDlm8YdzGe5wB+/bVtHFtW2NU+LM5vk5Gj9SgupCnUUmX2p8CgVHBl08qi4zWF
4OOu4IajE7M39TNLAPH2elzLXQCIDHHsqdg+X31yp+QBpiXBaAt1Is0sWx8Rvl6/
1wIkaJbltqYcvu7N+Ro6ZK3pWxkgReGLKwSTUYToYeVUD9+4Vw3j+Iz+KCaxC5SU
JuOt+eextOEYooFQE3Z/tVL/u/HzZu22IOSSKccHsebbRNQVEs4RqKDR3y6XRqbh
sitSYSSDaa2Df8h7MxW8Pwl+uuIXHdfEObPKMM/NEQk8QM3o71LDCdw+rkGfPWAW
F4a6naTXXD6Zy4lw2yK9NDAz+6suWsYZkGXiFGebeFyhFojdp22hEmt4LB9UT+LX
dXzjw2NSPJ1RVsVcWQMzHzhx+jvZpX8iBaH8pAEy/JxQqapJkOTpFiHS4xpBo+3w
rWe0VKPTdKelB+H6JpSd5Lt7iMkwRTsgmHCztl2PliFq6MAz4N5t48ZtFThWRQsr
tZTj3cQDnatJNnCIssr1NlJUlB7FtcHRtgts7/eeY0/sPxJXQmxr0xk7FouIyTsN
G0UzIeEvCjsJq7ItVuiFdib+O7QL/3TA3iOeTjsf+90j7DR+aSsddmQ4Y1J+KbCj
QxRVXBgYk6EPRO/8idkFvWsRjbRnXVCsfySmiWCx4M0Exg19uMDFpws/FnybNwJa
7eA4jpmEsK8lwF7T4bf3ZNJHaOJgKWiqzqLDaqQSP3YRokkFmYPfdNbDQ0PB2cwF
0JzGtW824ltfmoGyY0Cb2wbHgoalYhQpNT3xGsPEAXP7B7iy3sx1zaBsopbEhpzg
TpBNvYfQDM5fiizzX1SylCcuIjuXn+Q/aqdpo2MM3f19csWhnoqsgdhwJJXRsgzZ
+dsj9Xy+PccK2TKmpAEe62+ys0Xf9Jf3xxzkzPzGnukysXH9DkXNaGRuowT6ZQBU
TeJiB6AfGi9kSbjn9wCy/Y2+LPOmblTjJzYp/CtcvTDwdnT1Dcrd8D71Dl91r4I/
yUVuUxkS2oKENNJOXIC+Eu4+Wznf8bo128SyQ8vx2sS2ySpjSde1gi2nytzqxNKT
i4Mw+20t/In8rgEOndTaMKaYToEH448S8xQ7sK4lhdDl2c1dkEayTU44UaZoJsh3
iC029ONQEC5AopYW0YYq5UiukJbjdWDNSZpDBPAXgQ87f50Ig5klRzBGy2ZssLPm
sN+C9Ge0GQsbUCrgvhYSlh9c+Rq6Xjw8xJH5xQscQJIdjIueZYvjMFZfPYVMlBZD
5nyIxeQvrluheA923vKcjuppUaXyczl4+0bPW4SrVuInhdYhZ6zO0vRh0Oqrx88m
gwsnlblY31aofBjIar4OQ0ukGCnF+zIZMWBnIMu1xs/CC/NjAepNjLmAgwhEsWIn
Ugoqk3VuYW5+Nsi/JTrnDiQbPi0hFCvFAjzLsNeISscrl13wvKiwZLoqB8zINp1y
2i2zfwivB4CwbjxkuR+amcYWaXS0+ZUL9QfXGkMP6cY3ldMN7l32Kx6ZNNMy2xLB
eG/RGDPwJmWvjJobqmxt92clokWFn7kvzLOg+P8+k/gFXfrSe+WqukvlT8JLVMIJ
fmoM1CVbOsm2PXU/vrTPPyEYS7xez0j62tnFllWZyVFoybXbfTuijY4QHI9JwhtY
NgPeOwHXwLoiNUD1VOkPhbUqnDvDkYNOKuHf5Wii7+anxB89rSwnSXYfQ17SOqLr
WowdpMUEGcDpeWOAvXIUJekmKLOVnUQuAdi/8oIes0ZMxg9ZmT9bSNeQkehqiJ02
l3Rh3zTGVwk8MwvJOUDPER66jRvh+DlIFhx/dZi+Dpy/O9Vm8OU/dDxYfI+VDdft
9FyzDOh/fS1fcFzT0aOxIW9ieoB1b0BLjCVFSb7Yeze6sR6zfoEktTNTSXicBy41
xfJp7tCfIS50uMabko3cvq/eAsA8Ego9dO1p/wpdZCFXCebc2azuqx28+L6HSVqi
pGOTLMQbu29Rfp2qkwU7o0C6GtnWZJPR0XlqlUFUJgfnTYH0zLkojawtQlOy/hlk
66InHsHVVAjnSBorFMrf9tQbldIvZpn3gqe71cNt2igcequzV4ppze8SVwt5POIG
dcJhEF1pg3k1m8pRhZxeoaJhrFq6gTNd1KGlPOnaxIUzO21xIuHTnZ5hE5uSmeAb
8ix/jivryLs3+zLyhUtFbj+VEDDrVMsVIb1Vfq50owCaKMGjD5sRjbryxPDPUC7h
3LvymMPFIXqv3XkpF8xfWfxJJAe5exhd51BN4fW5n0C3S7DtUZ3q8Sgg7dd78GlI
33D41IbDxLdh8MZm0mMaupFUzhkMw1JjIHUYyKQaAFKPz2ld/cYSutbxYcQ+ALQ5
eKHdUDyBEKZ8Qycu5SXNeVfi1vPrLu4agPo3YHjksXpl0HYJfkm7ymAwUfJDPv1D
1ISYpGQm9L+1ww4au/ojQiSk4fbvKteJ2uUImRiNa7QtBdJgc3kpMIl2htNYQbke
Cy7WPwGP62i58PfjmTZZzHfhORGjqk8TpIKEhZceKpLAH6wshALD7AgWlkqt7xy/
0tmsnaUlhV7fjQOGNj6iseY0A0iWEBrKAbygpkXkAbeLJBlN8x62v0k1Zn5aPeuV
EZ2Gt1b9jhYF0DZVxO0a7SiipBONoT0JNKuLzTFSTNL4V6amxIkH/31iGvkzNGlX
mFV3iThXUwTJ7V2MO1GXDion6tSUq0pcsnPxYykb2qGGfSjWcwzr4O7KFaeEpIPR
54donJEAt4VhPJaVHpkNzFXvLAT2fuzoKnXhGitSigiMi4RUuI2XNzZjuJarDK8o
uTfjAmq2db4ve7muYCQPOc/T5M3rvlc7Vd57A/SXkpI2DRne/l00mtpwc80km3kG
tVUNeaxuwGaB2AujRe4sA1SOmrKi+sTC7tnuYkGs9yrVLP3zVkSwID342hwunSHo
KyfNw7fnV0okt4giOvSmljbFX0V8hkZyTdB+jWGCWiv+zGmPDafXjqyNJCyHuafp
N7w+q2RwdMYcDOFsQ19f1Xeva0CULGWWBWHyWLZ1ANpo0q172uc72HdXOvfhMHVo
Mi5OXdCceEw5gvDOw0yf/LqWS/8G1Gwc/bjz3QYATIrpTuta4RXblE+eW12uIEmg
PqoGdc9EOUgjJhrySMqUSJxs9XEHtmKRH5FysUCpbBXTboou/GEvmIytf87jWOsU
p2Qqd4vPS0VqtGyN7Y4wG4kNjEdjiGBQ0Q1iGL0dUcRxyGOYKdZrcB/0chCx/P74
/6PIUlCj0UEa6ofx5s4bcOoHh6XcsgCaGyKPCRTX7y7097VevxR+LG9EKtma9k/a
6IBVF7BhYwP0csCDRPhdHk68IjzpZakDU/x7YQ/qWA0WNuvzMvY5KL3cE/9dxx/C
CRXtO5Go8/GKvVSbwtuTX02a7KL+wWzjoJnKi7QvH7S0uMqTeFjQsA/fOVaT5nY6
B7bC+ijLmniC2h4rBxYuIylyEblNE+0WfhM5stscBUB3zyweHicL6PtBWDhUbTzR
umhhM9QaXK0iJysqG+ulZFNIF4hHTbhT9vpbf7WwFi2LgsNDDixreDRxU7pzFvLW
oc/veX+DIH630zpzSSANICAPIpOAV8fjqCnYCXJmWB3EdTHEu5duiw28Jqa5Fdna
ZOMV9CTiXSfIhLJatsb5u7THMjqH7W6dsyaGNHciLFJV5NZI2FqOaFyq0aZAY+0q
7jx3MdvZxkKiwrPayT1LlwhRKPNkcDYAX7/we6ZXpx4yd0DxszIY+tl9J/2v+fs9
TAcsj6Y796G9YrITz1eX3spyiyRD4E0jX92TGSw7MBRCOwEFzQJdPo4N/d/RZCmX
KCSI41CJdc7KSdpzSNfCvZzDceK+cYTjFexj/AXtTHvZiUbt+qsir61cmLuLSkAg
3/n7HK7r8xfA02Wi/CvDUwoxNslYVR3xWAwo0knMQbN1uWC+vgUMfrsyDDeNtrBk
gXf5Rcq7NsJk0l53ANSPCHTbRE4vkHSd0tETi6/6oYRT4t8HYZUu7Sp7WTGcKX8x
UiftM/pHAXtzpLGyh8lFNapymTMQ/LEJpIYvH1flk0y2sQy5Hg8sOJXXFEpCjHqG
s17HF5UQhTitt2cc3XGmgFcBZ97PdCWa7orZdqvg+yDtgcAXm/+Ws9xif9fZQ3WS
V4Z7gVLHIDwpdG9CqwxpWPoojiTHyTRl6qaQeDwycRTKcJEJK9ZQ8T+RMfFEj2nI
Oa6uBRdrM4x/ZwLL8Zx2LwnoTac6ZMChmSvqasXINPGifM+WiHgc+2i4gwTL6Fxb
pSnDg1c023tlkbG7R6N9UopdI6+BGOe8p6bt9+D7NFN0X5SLDfOkA3XRrrHMVKLA
6KrOuCO82h9nDUZntfxAaKq2+w8p0owuRt6W3sxKTFwdOMZSilPS3Ir1CWXIcf2w
EwCQmJP0JSZLvgBzgFVaLFZzpFHmU2tQeDMDdPyxjLMpXqNHAZZrrdPJCRPcbmKv
zOl9sowZNu/TfiiTAL78x3+6BAl0F5PNetQtiX1GM3wj8cCJvO+UOVGoTrX+Y/4G
FyGZpol12StGwYOGAXW8ovF6UfSHKIe81imlKuZkhp8MKj3/VhAeNcpdfVhYPUZc
ege47NUrm7qrzQnigrmVWp26sU+VTeRYkquSobSGHqnAWyBC0BCD9ueiw7EZGHmJ
1FmxIhCZB1Mi+sZ4pS5oyFNMojqFczn1yoq9uIa8NeFAwaGcSJHWTVgE3HtOat76
l2MIc7e8gQD7Zkw94VeBpyTxQdA0f5lN3QwInWwtpBnhjmvOIrGJpYY6HfD+WzWK
TBNBIAxravGWRJh5mDbACGLmiTEFVY6oln49O+WcLSMO0q7JISEtH8ELhGqZ9fXA
BaQvDD276EgN3+rkxUcJpxcPD4bHfQnoXKVHI8tfZBHycbscqbMcRdV2T1I7qF2K
1pdVa+P0bsIHtoqh3YclsOa9DclEAIJBBhhTvYhp7vEH26SqQYtIJNMx/H+263YE
dGp/w+C+KC4GupaoudDpOar2NQVLyV1V+kBuKzBvPszGbuY9OMSJ3VW6o5c5JAue
d1uRBAggeKxKV2i1Jfb0MBSIjZ2lWUizgT7erbgbBX2nP6smQbdWAgPE5hXGibkU
SivXzZ0DAkgq3HGermtCQRMnshgCHTlat5d0Ve7JjagCc3pV09swd3Y0dRDeC4SO
QcaGQmARS0gY55FVjCHA7fDV4yThv0+aIDXx6mgZ8JonW48HeoOkWjMZMzACGJuk
yiObH9X1vWfx3dr32wTjxA92vbjBJ0UPJ1PEE01makK26kzz5wGEuZz7j594OEfB
FqY4oJgfVKqL0IRzOwxsnyOV7Cw7gKvn4JjDxwnXIeMPivD2njYDaHDa4NqzQOed
LE12IkHEM8MARnhNVv9D2mk2IXp2hcqgPN5TZbEaFWIFVARoQGQeUMzNHv+Rx5Rv
dD0Gm30j1fIZdyZg6GvE2EURvP7scKZ4P2OxZBRyheANYQwp0bvVz7y9PnwJRELr
wpcg+aRRadgW24xIjTcJj4KJqUNJd0RwdI9UujUXDrOSSfzi6FUc99y3zcehcDkw
sT40xOWxQvxndROXlGyg3kvt319YP0mTmrkAGju8DCWeT41ol4dX/Tvd9lmT9fKy
TtgvKq9EqxJ8Dhj7D0JSkFRZVESVXSlWAEb1zMOpjoWH5zc56evb18nAsryHy2EU
9C2RCqSrUtiQDHErhsSChCgN0FH9XTvyusoAbmQUgsPQM+wQIXqEjKlbxRTpBGPC
ekaIKUgVYRTZdxg5vbQHjRB3jTeiiJqF0Hz9N05xq79Y5y2halSlCq9Pcru8NzlC
CW0LMfYIG/ORszu/9zmYoVnl+JQini4l4YC1rA+vyzLP7WYxrg19bB9Xwj3u8KWW
OcwXHDYC5n680nc4Xe5gOTCKUNEyTigZ/tbPKitKXdwVEoaCEi+BTbX64sw2Umj1
1igSER5mhneyzAiJimfxyRM/Nr5v7Vy/S6TocyEhqb333BDyzhT4YJlmvDwHC/tc
NqPgTBgi2KKZgXTOjJLrXP7WjHlACA9fwQIeLCALeSBgltx8PUQOyeuOfI+Jpu10
P4BOGI3wqQXllIdqqWyGHFV8vQiF8CsJM/SvBdFiV446iB00h0cyHGb2ydZudWj8
rn+JCTCwtOcgXu4bgrrbxbpekkhffs5b3UIrKbw8hslDw3FtXSwsKt/qWP96SQnw
0AyTvOqaEsNfQY8TE0RISwqbKLFduj9wxk27hYgeM5lUUjDiNthwOydF03u4+F65
uaZjTlFn8izc6UIab46STQmNYgdlRzJ9n2pRoPiEXvo9QdYAUsPPB95727E9Hf5V
1leUXk+X9edyP3/n1SnoAajUeOCsImaW33zwY6FkqAM1v6Da3bvxwF6ydUIpE5/h
RkjtsyvO1Kk/OYh5qMFk4O5fjFiaAQkn5+B0kGFZEVt8vnPognFWtoIHjDgW2Vw3
GYaJkCtBWAyYcWMpSJ4DmBiw5lzu+M+CRTetEpCDGH31ZxVpaHcSRp0BF3uHCnVF
A4WHaFgWuwUflDggEJ3V+uZfhN5eRRJf2L39tfXfo93UeehjnAfW8QMPNgZyn4JP
lu/Ec6PA86Ne8WhiefUcAUrJa6YGGK2UWlYsQxpK4KAuZDBXvPK+a9McPTUia2Mr
MTqy9czL7s68SMvnI0QL7k19UFVOARUIHI/xO1+phY6G5j9oqkhL24uTmkmZcbKW
iK3ul22iJ1YVVDubSnIZ5kWt6Nd5ZWxdjn1ti3nrpq0Pr1Q/UqvneL74pxXS+scR
l3m3YC7Lyzsx2nYR5xzIq5QehSaRIPBv9rGGFVli7lxtPdu+KtgDb+cmjF3MoHLo
ANOKU699FVI5QiwzFqKETwB7lR6aG/YU1vyEJw2DMR1x+5tbp20WckJZapc1siQu
rc/cCvFdLtU5+VyJT3BK8aswieptEiLHiNb4qfrlXNsyE7ISrhhFiyy3F3wa7G+0
Y4AwoWPyGlxCOSPDWZ3tevWikXsuSLO2IT3oS+Idz7/bvN2lfIloS4KhyG44I885
6nEoWJKLuC4aNpgoAZRfkU5o7Xf6xur77M/7OYWFMcR1pgnIwYdjgh8ywIwa65G2
nPlh3dszOPGy/Lr+wy7Vs1GsSIRxdZr1HxyZEsNL35frLvBl1rxOi7xMLgv9vKZt
y1kZVvDCTcAV9/aEuvMii5PHw4V866hEpCWG18jl7bQahA1cPuCtdtXqNN4ybhJX
PTzf3/F0C4enkka1V7mQ8Ai0oXQeRhIGDBn/K7gClaKS0VY30u2U5Rbdnn1czApA
/Pskh9P9dJhE9H1zlQrY7qsntPkM9lDDJvAzisBiTvCraEPP76yexebdz2+1yhtO
1tb45m8du9yxeiyj5vY0DIk3mP23dLKYI+crL7a3WoqdYEdZTpQHkHksWlZ+TzM9
Fo7HCr3ZNI6XFZrywaL1iWjTPENQJLfTORcs9sNfAn5JAOvP4FyHop7HSFu6WmIm
myyBrRZM24ikwQ47CBDWoJUZL1Xlut9dckyMG6fNZYRLiuBTtJnYCDS1XwF93K5n
yGQPrBSOVuKd+7gPshcrBbt2FOyx7HU6H+pHFWXiZVZ5ZbthXIPWyKfpcd/YEpg2
U0iFLehsuKdQGl6/MK+KcY5/QsdaB9LhtbqidcVPl4qAs2upPgvFzNki3PLmqIH0
ECnbDBVnd8jfoGxo8c0W8vujfePdq3xBAJCh+vI6sz4nSZUNrMGFy56w4h4C+Jno
0YJG2Nv7UdAxq/SwcTmn0iwJRkGPkEXcXgtGWrW2bRmms4N6NY9G9u1D+UFkHf4B
UsJwLAzZM8UoVyq1oltFfG3P8a7p92HFu7pxyN03A7NRigDwVEZN1W2erq2K9ahd
TIyCULV7xLHkJE+fQ+uyBBR+gVMSFdafOHOCk2LkYxC8V5aCRdJR+ZUc55dqE/Wt
Vu8BdYJijDZEuOMLNMDyulYydQCNtrvkQTuEELFFGeCHoxV3RIVoE2mdVqng9OtX
hqvE/X4Rq3fqdi7DXHxSOs2MYE4ghK6owNg2kXJdYYaAO7Jwc6ebLZ/GW081ZNlU
XEKqkzr4APYPY1JFuz8wbYdS1bKgfzqfIPrsRvatQdFZDvzRRN9dL/nOS9UIa2KP
etkwYfRBCZCOctanc2X+hwu5KIf+zJUH6Ot6VEQg8+zLVCCMtNLlKeByx6COsmd5
RKnjamO+tAiKoqkZMZPvzS3tCWxLWRwS+AvmNLMxN4H/lW3m4IBdHdYQyb/VJfQl
yYz7PMLX8vP2nC3FReybi0i1fEUSgAbM4CHQeRQYy4m7NcOuezsjOhqFt0na9HZ+
JszUVu2M+uO1kweVBUwSrWAhyRKZ7f5HNivWbt128aK2H9fsHOcbNSMTf6UGaayg
3YmpZeuD/xVNVkObOXkfxEetQrhN8hK8DzsyvQAoYBHnH2aAwXgmbKclarr/RuIA
4zpgYXuAKda+n6unug/4IG3dSwp+TrDSi2cRKANBjZyJ6nTQF807QuZzqTeLW/0S
edQYV6XYQN7VFXxun3tEDptBhgSvjCNqDkbrfjVGEf/URxwUo7KRFLlo0BPBZsiQ
TDNZ8ZKCXcIP8qhU7EBXYZrWlHUT2jHB0YJz7tFinsQ60/m7bZChQBM7QQU59gTY
TPRzguIJBkTK32vCRLtFht8wJh2p4/vjkTNaiNVNRNrVVEr4s7IDiBxQptxPXcVe
w5zWS7gGQtdmqbYSX5a3RNgGBUYlwOasVLlgtX1icY726iIJCVWp1NHG4GH9dECQ
pzPdIsKNodyGrtVKYbt5Egjmfg5Osjw0e+igLfx0egIXDTfbK84jZf5Pi6qIVxo3
zdgk7iB0Uu0xx1JvFLEhmIYx/Ji0vTn7boOuoXIYfM+1VfbXBS4hNXR2AdWu+EAx
riIFtfz39uwaqh0hqFHa81OZu4MyXlMl4NZDuJXFWz60OuRNXh+6glvkfkE2rGGM
LGHhCVfLkr/2Ib1HtPGTMSxZPnLurILPiOmJdQLI0Vv38+Mnd0ciokICVv+KFC3F
o1Ae541Jt6dPv/544gfHPpsu+h0pTJCGHk+ganWxxzM1l/4nl9RkSZD/YqY+aq6k
AS6MWrmMg6S+T/rvrptdUTFvX5npWc+/8yQ3qD2cP3GQgEDX6yrOPAULWUpgrdx7
irat6PhXGUZGn7Fm+Ma4FQqDvvGow0mdctz7Hj0sl+TMZ4mO0N9StjsQxz65dVAd
OGViClwULBqYBaIVj9ZR5wGhu00TCjUp5MWXSjmY7AF1UPPR0SV8zg7fgn9aVjU/
7NRSjYzLChsNXVkKIwiWBGSCwdIthO0TG+tfoxyx4XSb/eOeIJHsdhK/6YwnuVsW
ofnCIbhk+42lwX8jgsT+Q8fq5UWmCdXFvucpd57jYkFvm7ipE1PmAUgcXwH/Fcau
xD+OT3aaoa3nYI6kIXPpfLa44QWWLaKhA230N+Ru9ZJPqt0ByKgsKqfE4ftZHE/O
K7caFqXPOlQN1QMbUQXK+3KTTR0GvGyTLhNiXOQFi1SyD0r+p2h6GuL6wjO4US9C
o7fpp4tIvrDX9dvXfleBBgSRzfOm65xb095d0h/ohYKK+QJMQXAtdyZq8rtE7tqZ
bGA/H6FxaYx5f0e2+v9/9Dppzb41t9Xhr5bm7nbLxGt0Nl5KQhjGs0b66EbvS5ti
SUoIojHlUVythENufndFwRsWdRqHZpO/gEhjs2XKG5DcLauZqh+uxFhxp9ZKr8Cm
vAFMpeE+lxQUvQPiFhEPraoeeIJCDZaEFWL8CRkvU/zJ/3PrvRn1Omx5Z/zsE4rd
DFmHeTMU41JhmWVVGXCYep35BS8Jz74BEtm2jrNegIlspylDGg0MIKzv7hniHQTV
vmhPAuxnf6vZjQLCS8OZmyyWGy27V2vCUVHc5d09JUqu2pRg9mM2e2OcTvsc+P9Z
BSyoYEjS056gqGLHkuvroZZhApA/asuULwXsMLneOFtsrwjI+CteEmn70hq2W789
uBErm+0/NK3Opn3DHMTqTH9eXsJX0LXrBH75sBN90R4wmtwAZWQQl/nC5nI2FX/n
f7ro4M5159EDXX3vpnNbAnizKKS4LFZrM5GtawYkl8TVWwpgqumuGogelYdFvu3+
qoLXIIuTb0r0FdoHvnnxtZB5gPl0QO6wKs2po60TCrexZYbzJsfjrxG88mDIndwW
pBbEKvlGx+aghpalivbJE9W0fZhpGnGtXEaKi7+b8nPY3fMYFD9uWJcfnJTJw6vf
2W3UtAFL16xIf0Kc7lSjLnVH//3z6lJHHk+8XIL2ih+sROya5pXNga5R1J1BWNqS
cwT5PKdE+rqc/wBKYj2DFR3qhOo5kZa3kcJWiTex3Cn0UVPM72SfcQUKKjwY2uQA
Eo2S3NTvTji0CteMK+tWyYtffbfwWCZPRw49k5qWlcuZaKCSJGWyb2grusBdnR6K
xV62j5mT/6kQWODYLafBTn8P+eHijUw7oq/ujFdSC8uFNxdphGq+0WpLnJJGOfDv
GERFurigkHtc9G/0noEzeoncxhN5iaJC4tqN/p77NaL1mjSGV+wWWMsBRJQpxzh7
xR4ciIl9PmoYorWp1vKBny1JKzAGJloVvz1vkNrhUa2BnbkFkmxFW93rz1eMpiw1
zuwdJFN5YduMjYBi53zRnWbefC+nbDEnigMS0t1U2YPAVXjgPH9tOqklcCm3s55f
Du5QlRo+Zsqj/YwEswcG2tWZzRx4AeEiDlg8uS4XUYDfjlAZA0fBlDlcv5Q30bD1
qeRGaMjlTOqev4Jt8MIWNAbtYQ8effqkSp0On892PNLMPTlJia3CqQ5QI0KKKMiP
+E5gO9sgKPH0ycnnIgCKfG1jsQ+yKJNTUIGKxE9k1USqEIHp6dRaL/CIKfWU9PW7
ZbzW/UKO1wCgf55nZF8GZT8YnpooMun2Dr/0N7mb5s/TG7Y7cO99jA+wYWKJm1HB
OzzP9zPOOAqrshFs6J0txz0kX3HsHOUH2ucpl8k6pnBGaq8zby2KDMHx9defeeCV
l9sP7lJox1gwqc7UxwGpjQHYBTZjK3VI7wCmrrwk42Nil0A3T8wpEe2lMO69VYmr
xum9pkuFX+76u72rJZz5ilhsFO8eHsseXxgkk2Krcq1TpMswFm6FMajHMyWigpZo
V0hA35thpYPXzB3pga01vZC1FvpTeQanQtdYy8etotiSwhpYM3rz4uXfmoW0bS0w
G9CArKkYdgDJ1sJOfYv6JP0pCDRszMCk9j/lnyuL2bg4QTQ7SKMnUpAa95HCqnOj
xf2y9fUrNq39Z2EALicASEAZZGA00T2Vvuj8XRQgy+R2SOlifi5DnN6o+m6Qjm62
RySmBGE0SBDy25qd5RMM4wloBJAjMYBJ1iwMqyT4Rn6Ll3ceO9OciF+skjL6mfTJ
Lplasa/HtO36Y1u7KoXiGURg/0nBqcqCgIjYj7xmZvnIGu7fTgMyqipOokDCDTKL
4gwRi/hpUnn1WrSOwoG7VNIbunOuxQ80rw1fpPqBuOtNtnIJjMmMXwrAmNYIuc0b
f4aDh1pyyjqtGZ6lXbqOuox6j3pFytWXIeJMPezPS+qZWs4IWkcFKpq7oLRf4UtS
xnHo8G6gZNjWETSfaD1z/o3KUg9X74zsX2FZozTucnhgM6GV9vc7GaMqU0Jt4B2g
84YHjo5wQYCPbbXVTuD9Wr4+7elbnRu43BG5TPmzQqCgQNYvNwk8NiUdyifaEceL
9j9LA4Ra0/cbHaT+n1/CA1WMau6RMvbgGNdLCTnrXo2j/uUlv/cleK9qjwFQdFuq
PHRMvYHY6yqR+O5cren6FRlUALUXP6srBFObGaLJQbiGwytEcuFUUQzxCTIVZqAa
cdnLNxpVk6yFJRKPhyWh77aDaHp6EaP3KXJbqdBUaplCqgaEAxVVpLfxWXzx7Qv4
R+70kUIHb0niVRx+FF9u1OUlvUHqLqpt1V/cO8y9VdzTbaix7e9QHpCsaFX5S+Mg
AhiiFuCjAsqPWY3MJl7SQ6J3mq+orBxAzOXBCc9UK9l9ScrSG8ywDV/695+rRX7q
liON3wTel75fx77FgYsmHBCWa3KB+kvAoQZzTGlv5+yR1OpYqPaW/ECmazgs7bb/
7dOIzjxHPWQ58EUzEZEbASR74MrOXoNMxVsLy8JeEdfBAk4aFyMl205fEMoaBG0n
PahyTo0cUWovzMzIloQE87H+vfbII14wtPRic1pjZH+reSN7aUkr9+/rTGD0jSfd
0SV4YMgUe86hOZ4qmg+4mDP4i1cmpFHBkRPoZlSDNUcWkrpGxNTBpdLdnjjDhm0S
nhz02PCIlVOFVywGl7Bv+GmMNtnwWRT8w3yHKuTGHYdI9XjiL7qZPMCPyUqBqVR/
GHMxElFNi849JM3rb1bL4dLi0SoPxWRC9gR9TpB2liu1QiJN5Wy3NlwHZ5OG02JE
MHVZFySb/nyitLg5im+A8RjPCa2v5J3WGrFtDEo9BgPjtJ7pKVj6AVYtAZyMFLhs
Az5Kscxt/hY010XwqYV5qgjJcCdBlalz+Or3NHO0HwqNsWbk3hef2CNY2r2GbcFm
Ml1eMEh+vMieZsVifvt3DL2yjQNVZQh84jyMpjElvANrbAw8+U6n5kgbMvFWJiKH
3DoVOQNSdIakGXG2S4l06IELT6QsXBojW6GvDdkSmDXdQ04hrFASa7/adSw6JEAo
YdChnyiz1+eAN1Rm7qy9Y5kD7hi/t6ukuLWxQsbRpx+4YnBw325ALao08PxHBGzC
f9Z0DRH0prPyi5jKAR48xTgL1ZFJD5VBIXlmljOoXPzkIhGBDGP9uNRTwbHD1wD1
1L4sr0vZJh3wnlnvpT7Lq1/DCjlFVefxapgWTtLp5BQpIT13gsV1MYJPpE3CVCeN
aCKHxmvq/kNM5olobPzb9tXccHRqDy+aIJFpdc7tJw3GW7bXEbdf28vMtjhl04FQ
GfDYO1/EETYrkjMFxyxDfpdF3mE/WSLEtFt7rNgYrfa1lb+kWhcvomRCaO94KA3I
noFSKqgbIq5gfcY4wj1hG8GobchBENS0YR95FdOBOhrj1BqFIIVhSn75X+FEK/4V
3wmXkgCuhQVo4znNrtua3KEcFdhAAV0pdelq+eYZzpUEf1yYGg7+iEg6wW1lLPB4
UUAJmNYe6PYVLFVlXKBbAR3Dla84RdpXW6vROovjHCx2454v+8354OFJYTN4wfyU
vnJtKs7wM2xzoUyu1eT3u5JDDNjd0fYRhUmrJ2fW/N49k30J17H6cjtuyZDs2FU7
h+m6Ogn7K6CJzms5SSsseqnuNHgANK5k5GHkFOk63vai12faFwBBN0wgahjKm+r5
S4d10tqSSxt7mjE60asb8o3xHgVSqe4se7/VymGNR9zPHwd1hHZRG/sa5RELmYU4
0Lrwp0dViucbW1j+mF68JpMFzYD0Vo1nejx7UzfM9GZdlvcNEtSL9ghISYAUaRHR
vEEUjrHM0aKJ8upnMKEcMnH+iDHezofdlBT7VViNVqW2ufC+coAxhhTZNrSm6qOC
SZRXqmSHXzqF/+U+HLlW+CG7yC3Nq65nyiQSFmsvjT7Zj5wIrlPLFke4feDswqx1
s3b+IVWa8BP8kPHTcGyY0OpDt2h+FSNF7njy2i0BDj20A0/GRD52qGsXJCUM/Hdd
AV/Rbkl+rvvCRH35rdEHEVgQuOwZQuTbTeEtRqQaKC+u4pwjWoRKCiNoBqOniTQl
joRd0wIV4vvtB0N0LcvrvEyqzg/wBacRomcadjcWVf0wss0zVNXGRrAQe/dgwVF1
3rrr7ZwTqSduCPFsVFl73EhuR+jAVThWopm2ZosKlfk+a+6874bqoG4gjL3HYI8a
gMpR6u9kCtjJsEaqI5prmcgKb17lwhtXYCHGXooDnp/jnBc+ehLck8h1YW1eucu6
oPIbasknGZXmvNnuKAxrNevWVZL6hAYMbXWHra76ynkyVj2tbc14NhXmSqnv0Aj+
ISaWIiOjDsNo55MMYBRH5efu70I5KDGvoNaaMCwMBV9xcKCirNAOE7x+JzdzytXM
tCXXjDFgArAFLNkMGRh4GeHhRH2DBHHGf/21LfVKlqF9GxY3GUzQPOXRpX+rgnE5
D4COb+XFzriGYqL8rUlb1Le1S6jtGc4pNtGoWkH7sMkzZHJn87PKzzh+vLeRc79q
09QNQ/Jqf/dOaVzCojRCMSQRAGm/UMNP5MKxfh5UcSYcu+BF4tLAOCge7PcTAzmU
DdxWBoyHoJ88njkaprqAq1ROf+bhkkWmVvCi4M7pWcOTIxotSBCLtM8Fu5gStrE+
0jV1DNlAo3x8GpYFeVBQjLJVNbvpPkR+fl8m+FpxpvJ/uWUIQTQ6KpgLATNgOz13
l8P478z0wHF2XV7Du8ff2DOLcBfgvF4U0ZYu49OW00FM7ynSGj5MWe9i0l/DJ8WL
N/lo0INjnWCZvhapOTMROi3b5s91bgoH0QMiQjl0swVzpiBJBbr1yAe17RYklSh8
fCK8NNyzo0Z6qi+Znun6xZt3kf0+qEjkKfTENL8jtBOPuPkVQLvv6bv23LTxkHR1
DIpT6aR/DcSYpGFlece1T3PCr333VGhUXdoNru0geWTEXh9LLO8SkUOX/t+cP7Dc
zugI3Dd0Bg0BhNjLXofMJk4F763ng6NxDEmMZDRXoIC1zt/M7Z7VH5Hs8CCDnQGR
ouxawBqBFovYylgDnFkXDHHjf/IyE0PiepHkT1QKo05Dqn37BpfhDghfGF4oe9HA
5nrZzsFxudBHzLYuMUbIE/Qfz60XGltqK21KsY+vN8SiVDcHpKHgpoDLd/NxQmWC
I6a5umvTczjNJBDqRR+ns9eFdyFs5e9XLfSPQHiy8A3pga76NyqFBXfk/zpZ21kh
YfVYiNp4+0MCm/gwYx7MHogt9UmRf1MCkpZbukTS/3nVcj+h5XwITQTaiXY4tmgP
eTzrk6UaytPe/0lQdCcUJ3ubNN8kuoxJ+U1ksyfzZUcryyDRd/QbEHyz34UIc8Z/
SSdxbpRLA2lS3gNOP4KSr09JQdEri2kDvthGtjvAUOBWnZYkbuv1r8aleREVBovG
+/hLHhUM1LoT43Hb3R30EWribVox1pRkaUt+Dl5eRHBmQN8/BxQlcGFgsC6//cjt
TRKDXKZBD2mtOWPb6rK57k6jPmQmz9QZXZsSgyVAaW6NBanxbySynTGAkoCNnhKC
YJ1ZOhaf4BpDkJ1kFDpcd0mEGh5j6VSc3uw7xSVObv+pp5wpDBC1TEvKnUypHlQl
TyllOJ9xvMyX1ZGQlVeYedIXozqKGZkcIpcohjkC+fU1znc1Qd/CTB1nglTmW7s8
dbEgufzl8C5RKejZ3z5oHe/EuBQhWUxyh/i62uEI+hw9xNYuOeakzqfln07f2Nqz
H1kPQZyMB8SxJFbZ2QyNRm22FEyzc9u2JLh3ZPg7KbqaBCl+G+lc8MXMMaGHUnoY
C9fg6wc3qDrCVxWiuaG6mjWlAht2auVcHhNA+phf7OL1IGJodWlT8sa2SBTMJFPr
5Oylw+scvs0k7qKH4MfjmOVW2OPmf3fIO0UZ34r3rTLOen1fXIWVP4zHt6qs9xFX
mo9vhi4mQdf6GdtfRzpEFs3iv7IQp0SS244oTYzClAJolHkjqXeWtc+fP5fBXSqg
8o4/T4qhrwS4cAoCiEn1i8cUYP2dUOQgGfZQxHrlsGWZHAEpDA9aWjKdXDMJmHYZ
dIudHAGia02C8ilT/Ipyj3fgonH97u69lStP/VF5NrV4mU6ZhvRVtx3+LpiyYvwI
6FwKDe4elwmIIGedOZyr8OYUf4p6tdbb2buX9Jat0SVgNn3ZerrvteWxA2tj9LW6
FmGCPV84gsnGCFqOYPwhQIdTx2AtjfZ2wzGFFzTVwey/rBvT5+3tKiZvOmi678NW
NwgiHw30kwcYctO+RImaF1H5Gd/nxkfpFrQG8pgn3On4QO3Dlul5+qIDVOGK55DP
7PBP4qGVFjCxB4rxpStClvuPWS/gBEQJlzHqNPZ9XSUGRXs2F2t8YpJc3ot7oVz9
JUYjoZYj2gJdDdCCzYKoluXhW/O7VFFpm26gkK6DmjPGeZOTw54drzqkjCmo8Olx
cC5cOmXdVQabLEd3cuarI75njG81PoPudKQaRXxHlknIVsD6m8sYXWXxnnPx4lup
qnBvK9bcuFYOpwFOcDKaG1WYE5yTXDrVBMy1A9e429EY/FkXw8UxFbmUZ05epmxz
hNK2d6pqt1X6wjnjYltirRlEqzkauyWz02PLBfDNa9hIrCCqR+Bm/iN7dmVJDkCa
j2BGeVCSz0KYblo/rYQkS4AAHAlyD3LduU0moTdPByJw8piWWsJ1fhag8KzYqaSw
7dgrHZVkidOnLGhf8GRsIkBkSV3RLfHPmBMkND/IdP1Zu9t8PEf0+gWpGkktdOd4
G75fjj11o6Y/zSIFgmj74A8PeSsIuvxMB93/qWHZDkGxuOrB/9zWPE7eZ5xU3a7m
0d985tHjh2KQ/lD2/b3DnGL5u0sE+8EwdMWp7z6mSLVijkTf9ONb4WocXMSqvIPs
l+iPJ4biJxlAAOyIbFgjhAcEmAjHZg2oHexPkw2Zb0AN/PUOtxga/xqiB7nm9Kb2
rr7K6bGWMForTny+t5Z4P16+Kaq8AI/5tdhASlfClS8AhjHFAkt1yu5ORVUhA4bR
WuOqbQ5P24WjCran6W2rcmpNNTh12LA2mPert1WcOELbwsADSXFSDgagKHmh7x3r
WlYx5cyhp9abo8rG55f+8+8Us6mZ6ae6qeTgDJGxqv9eNkHSDCaGdclUD20DaGap
8r0qV5dyzmKTjt30yCL3puXznIdZkXKu0VTl0TZFM0/todRQy8qT4ZOTwTzkRCoe
W5xzUsKUqWWUGPB5hCKtowssbVAjajYnll9suRJJQcEVOka39e5s6mwQCnn1leO6
O4DjSy7q/kSiXtCPwXt08w0OWIEMKwauXY66eX3MvxkqbXEDfwIlDBPFaxXDILtE
p2SdMHTv0uZ8/Stzurwqp6wWrVhsBL3GGCWOkaA0xjDvk7JKtt9drK3Ylz9W3Tkk
Yx4wiX/lAzS3LqWgWgH20n019mvAjdI1MiNcUkklYcxzTzFjaBNadgOO+KNQnUSd
UaZZeU8EiZSw7Sjgb9gEKuURneQbPKoPReOoklT0x15Nzkg/6G9JABv9FsXPqPb2
5wbw3Ih3R4MBn8Qy4zVMouhW1LKst99ZKuGEFGZhHri+AFgsmcSgbCCSPLTU1EdL
kLFNnYJbGULiiMi82cuCxI01A3+PomMttBUq/axWLhpqJ1rBYf6UqJGOihHx2LpY
O/fcdwbqu7uhK9Itn/xAkIjqOocQ20/8I5in65eaxcDnXbF+ZQbIMM8z8WrtTC8R
l33arbkVI/Su1gNBFfMn+3KpP76za7hjwyu+PZtwWPCHoohbM5WMQBpZa+cLvlyD
SkltRtoRa6T/FNIIKWnNPavESMON7tmwyJ4+VqW/o+4iaSy9r/kt1Nawbya2ATxt
hEdjZl4QXR6Pzq0JjaHay6MYX2098Y7JPgou22YpHKmuzvg2P3E8BRBUXYoGODOO
Qs1YHAsqKBGe6eeBZuoCJPlBJz7WMGxH2NvECK3CxfN0qjaZpARh6p/vbqeowzu7
Gf20r/u0s0ELV6PRF+XvVDdvUaIqs7EYzZ+05QzZXXGK31hsZl4Pkq+sLVkWu9aZ
`pragma protect end_protected
