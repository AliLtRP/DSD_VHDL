// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:24 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
WKAtW9XvMtKJRKLfKfkEWzvC1Or2Sd2IJBwOtAzeREcqg5aHEpI8918KferDiymO
TZvvVXO5X8Hl494OITeGZrWlo+BMRRdXL6hP+mAmNodrEtCFyV6VdzXxgfC2rPdg
3OjrFi6HH4VVEzR9VgqSe6Fk618TSQtul4j7m8/JMQ0=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 7360)
lBNQgmucUoIo6rkn8A1mX+UFbjKAbGgnQ/mGJ7jjvJfQHhfgpfj8+TQeiYkdW2w2
ci4zIqPbY/Zq9O7drX0VbFO2ijfeJVWPFkfv877o34QtbSZXc8eEsFCCkQw9CtP0
A5hu8KJZze2109VN062A/WP9xFe0UHwVQX7WOKS0DjznSCASAk/qoF9SwXoyEUM8
zU2be0gAaDiQXReR0GgllwRanU3Ic8s0gTB5kYKU2nYWwjapRoKJWtdwzj0seBxz
zuyp+RTQXwLVvkLTBvORRqQJAQIJ4PXooL3CD40q2sy9kBWMQ95UTxTImoxvRzdf
6ZfB4G/TyqLxNiNavh4Y0LZcpl2YZUnKneRQr4wc5f9LgwBUPzpAyU/zrs1qy/gH
HfkMIuMj0BDbVz70Gw9yZ0g7GXSwD6nKLdCUGnAiHXW2Hz4GifGgcUTCp1UWsBsx
TpIuOiRbSxu6hGgnXMqp46DTDtZ+r/S7h965+ePJ7a7BG6mR78le2oJBZa5Gz7IQ
16PX3lvk2Asiz3n+Lbp/xA+rWiRcMosMfRKjXr9xOY1T2h5WUQ5UD4DwQ007qGb+
y6fM5K+SYSbKIQ9qgVKVvUcq5F2R4Alh32XMl0o7pmBeRWMeHR0Cyn2v3uFqkguL
ewviP1K35cViCtNWpu5BDB6YY36M5dwTcvvtZ7qzRXg48FBzTmF6BhP5pcLp6gvg
B4o6Jxwq20dnh8Gm6BLQve0awAZ6JOqAT5aYwwDmits7oWPgfnYv2fi/2tYxeL12
6etZJtmtqzE9Cl61HGT6fyJcgiUo2K9iHzoVm1LaTxcIsJiLl0ZMjC8sWiB4cH4W
Sa/SeVEnTnnThBzepj3knOuqlCB9y89jcPLfyXZcVuzHwIpaznQKFqFXmeFrtLiM
qeunpg4CkwHzK6FWK/nR9t/z2eS75Fx+uk+gmlolAc6TD9+PMVNNmlNLB7TWBA0F
HpmtXspZzL/gmN5R6+13BU4UJWO/m5Ki/CaEVUcMdv8UpaklhUvJBXe2HCZrbHBd
zn97HiWARPQphki7NbULhGWA4cHBDWvQzZaPiK7k+wXJ0w0vdSvSKx1Pcjifu9fl
bkvj3OsiH/Vj5dVadsyHS68xdWjvA1TjxDp2iWEFOH99XnF8cLMvlexZut0loiEQ
EhPk+X3EDgS85X7I+KPyshMGR9iLIAEr/qdSOHvVY2j2phUxEAf73f7enp9ne4iQ
tcIbrL4SSlcoNRkRY2zEAMgZ2EopUS1YvcG38yWzQWMiwHO9qOxp7i/9d8kbCiXT
KMtYUrGEGux5ZH6MCpIkwEq+4i686L598olpw188xoZjDZfvZU8pFiliToRRxk9b
Rx5sVg7cWdTwGtU8BdS2VjentAr3ZvtmtDtI5v2UaI0DDkaKLo5DEBjJmnOCjBlS
8nKT2pZCQUbWnqctW3E2lHSfRGPusBQwQKq8sfkqV8Ows1f0B2bb4l2xdi11o9fX
iM6F9FdJuYOMgSeIOBqAGvcEpOdKBQKwgoaTYrqvrlDpmNjwADW6pjkCK4a2S3TS
CfD0jCvrPJnF+37kUXNBQVOM5A4sEZSnXdPWFN+T/OKU2zFKqF2J4Nm+WBOad81f
BDuJYYHIsHYlv+GdmdAU4Q2HV0atLs/AifGU7w/ltdcCn5nBjHWlQQHpI8U1PggF
o4DnaGDIMgnW5tIOoDFG9qPSJ/7f8UZyI/I/SQ3HzU8g/m5ZsLPlcfmIj+m4XVUs
GqND4FSWdpfQkvYRjvDdtCL7dq9gvbf30TH2NKKTf/xzMWoohkJfE62yeKPxLJqa
4YiKA/ZgTdHQjjIta2aSXNQSFy/f4pb1qCT6CkhIIIglJQ4Ire2vhhrY/RTuHwAR
REOrzVU2ztWQBbkQ2CH7yExQ9A6kuaeqlp/OAWtyGSiQtHBl+WSRKCwvjCTf1Urr
W73DJgWtEv5so9JDLnYpI1s2qpiiLR9YPScrjm7W9umH6zCXHBI8ZsB3+gCtztD6
2e/vQlPQnu0lwW7LFn6SEX33/hyfKYm3GHQsgiQVfb0IdS6iR9ngw/H5lEUMG83v
P8uNI74n9tSq1p5Xzwqwb+iGDX6Oy605P+fqNxQAOlTpsrvAmrjUACKSfrna2yK1
aeJFNaueezrUkI88TNjbhYifnfyvgq5nrfOxU9nOXVKddt7XJVthn53JFYXqsAa4
fZ754SecMbDmAYoo38B1SkNVdDsziZjRbmQoI679+hYZIkyh+3pFB47aEWfAO/2G
B3MhgLiMl+H5bJbFjQlRvx2Pcm7uQZ2jhWkNjoBksJFecqauJxbaIvcY4AxRNZLM
GzJHjIycpj4cL1jBKsDs/H5yypSMbi4wql1etwVNIFBFCSO//ZMgefDKb5miKGC9
boa48H4HnEXYVDJfKYhe7hBdUTmizclHNRSqKdHWd/4BrR4bdmh1J8NSzv/F5Rau
487fFHCvTe/eNZISHLyq35DtNCnYRJLrKhBil5lC+ip9LxKERgmoN8qVQ13e+IkC
53RKgIdcTwrjgapJ/EX4N8tRXWZLAs7Q2Lx4UAsJ7Jt81l7Rj6wXdBsnfQd29vvC
EbESeFlwJ/l4Zz+wAuriiVF6v8XfVtzy/jSCfGtcUtc7GuVOZBucf8RDMusM0mpQ
l1DJQrQIvFPGhuiuwQjtDhTMy+3mXTVt8hCDdX6Tqu30+CFcj3sHLJB6HsjwgEb/
VSRu7osZJXP9+cWLTCKSXePqEkWJ4FmEooFbI8NEnH09QenKiDglxgO3+0LXecBY
Yn9bMsSrMtIhUTYVRvuJBhhXfeiAs2Kd/EzbVZh+f0VlJS6A4D7FM9t6lOfZVBT5
X/d29Bap9jyOFUalC9tniN4M1SaxXoRx1h9nTu3J69a/rmg1w2O8SnrO8+PETbNY
zXNSwXR5mAE6KOVF+UPVKfOaTHXjx1xFRcJOcmJ2ESg9O25sJFZ5DCRpooZQ1sQo
8i9/VRtktCXXKUqHpZdOECma2KtwotqFyaIAMhExwBQy6Ywnx6dv9Q+ZYMuDHVcQ
c5WM9fmPj8igKAZEvpCx45NByyev8iX9fRf4Jdsv4rzv4J6nuWEKtzb8YQ74MwoC
Xh1nKFpnqzLRA0LCTb011W5aWuVUA5Rga7Zq5aF1WWIQCIp/mYHdwc8fYunB/RNb
hNMnctvgkrP95RKaFm2qA/0QNMe0nOJlx8RJtyuzr5pwoXsTbp/tl/krxRS6jUWi
+3fwFJbH0gW8rasRVXhvHmdU53bkwcvf7u62ZZIQ0a7Qfbuvcq6OoStY5wxUA7oL
5jeIvXnP8wrn8635TYZxIF1A7Erjh8dnGsiquur6y/vJT0xosGZrTHuOz5UavAdm
mush8IY30SmKjXIoc7+l95Ztfv8XgjB9x6vNIgFoto/YflfNjzHd5GbyidZl8bpU
YgTnxwOA0oFORJT/q379CYeuZ/2ounsZSBHQ4JCCUvCY6ggabSuXSY4KMn+jmY4p
yYWzteDLRh6dDpJA5TToXD02RSR1J3Th9fz95Al0IzTjcd9JGGVO7R4nyCZJWI55
pVIBiChZ+EAaNBYZsH7528t6DbkPBxrIJh7wq3E/3k+EC3REGNYN8DeM6egflDtF
LaPy3TdmjIr0oNDk85pAKC+4eNdoBU9WWAUGcUhu692ZNtiMUlrHzRYWJOX+tHHX
ExTG3EHGqyWiAwZsbDw3Z8YHVC9kMXlNtY1AImT3zqYy2EnTPpMjEpv8R0pDpXL+
D46PsP/7Ms8D5AZcUjiMyTvh+68LgrxEu0dxUpsLDksWfw/dTXIjP0fM88chOUO8
wGOBbdotuNms99Jicf6lmrGtlECSnsjESx2xW75oMV+Fru6ay1M0uX/nw9ewb6Zu
WXEmKJaWoUAUpbSpMTSQH3r6KGTfglrnHnArabdBICXiivXzvJNCwC03xoTNBeEq
5/d3whYzyiBD3Y/kpYt7O6aWiJdZDcy1r+cTtqQdlCT1xhTFEvaLxyIpTbWcN8JA
v2Izu+umukew79hGfxiYEejzh4L5Uu/ysihS6IjF3ywbNT+G0XcouMrjP7p63ATr
0wh4lwowC/xKn/D4IYLIsiNW061sPEE+kkI7OztwvBXK8OA5fjvXg74yTc1FlnK/
umTf9j2+JVO0yMgTGIcvOHZu9XulmN0uHEZaKXYobyyQ7J3QFWLXAaW65LnRKIbe
cHQKeVAdsmaeZFGhotCzOEnUPFbopDRZpTRdZjw8l2eCm61FRdUY+YFvftRhj5g/
OTLnwPUP4D+CJPh3wTfjDEwCQ8ftJ8NHqC1rUhUI5Jj2f7OwiyNhK7maxDkeqRHj
VmkgO5E0zTWy5COJ5pjY+EntlTuQgPxqzWKBEr/pmhQ/w2tMBS3yqiENYYy1uOwL
WZwejVlwTzSVjFUKN5vw0R/8Ry/lY0uIeivyLs8xQFkZvnJeHpPUUp8Mb1F7IgAF
uGhyWQwPjhBaRDf9+578rTw93UAhlmrIzgafA3LIFazt6/oGHz64CzSu/8YqqIHy
7r0I/l10Cvvz48ooVs79Xrzq2ok3AvFCEFvXfIC2pLKB2xcHWhnjyumg2kRPYbHf
3yLJ18OZE9NxPGA38yd2m6Ipxx6+Eg9trY3QAYQF2cBJUekJgtHrIhVjadexFM+l
KysPgHSYsVDuPYdZWsf+7mJ7jyfeLLD4cNz9/IaIp1FupX9+D318c35aqI3+xNxo
lLZWbYw6YRC/Z4YN/IlX+j5MlomPN3X7WTwfCE9CwGK4cmpiY7d97joUPvTZyXsO
H6wCr5ZXNmOuLVVMoeRcoP/glUGGZ/p2Q94OI/33TAe8r8Ed1ppVrx3UhA0n7CxE
zLKLy8u64ZUogPePJDlR0f0fvBRgnIGHSL0sCMYtFdP2Hxu7jlkwimvEdydn1yy/
fuksa9lBQq0vcDzGDb+himS9OOxr6X1GUXP7u7aQlno4/9SrutCQlgJPUIdelxIz
72AgILOO9cuxsDu2cfNYGJFMVk8iiRoxPob+zCwAvPuLuaYX+Cu0xInvQTmvVerw
jhQtZUOcm68eYRF4GkU543/SxmOdTgw5xOAya1x0RpQPT29WQuSlxdYahbIHj3IC
n+8Ad56J1Ox9l9HRClmjOAHtkJmAs8QdXubKeX8ivbd0u7hnIlde5cIXLuGUCSbC
TzkGapy37uuOLbQ7y2t3I+gfjtOzxOD1LG/JY3XiVfnaeHF9ilS5oNF51JVS7Pbi
r2hebKVW388U43j4MTqackrBD+/uUVprHIOKDahfNvyW+BWbfX2BXh5AiUAtxeqZ
o4299w2YFCYFVIBKIar790RHJbhkgaAR6EjSFYSyLmetU+/wf+Y0T6a3h9YYdvcv
ajPur5CbVj/l9Bi9dzP7eryHO/4EI7fWMfdsXBiC5ISPq9bE1RTYZr5hq9Xl5vGb
8kpA4tfzI9AAFBSHGgLogzqnb8c659izqtHLFwr9dr6hols/foBLlebGV9+935WX
+S2o07PLBDQPF13/sgWsyJw9DyY4TgGdjdSAthF++giXv0lDjRch1Lx3h33xtgpF
qr3sVX+MNGaB1KiIMcdDUvzkf11siAbHi1TFhMOPz2B2LhObcZV3O4zVoGQCFfPI
YbGYtLzTkQQRU/09gQIgAixk5bHNnS6faGhGFqh/WCYaCGHMMMwOhpMTwtH3aaJ0
/vWTdHG0MvEh2NXV+DuO3vvS4ucxXPmADgHr/VujWex0Gt9gc2NS92NC+niVMYpm
xjuVbAesA1nqGOnWoV1/9zczVvEYGEZ27z+6J9OHSpcrg6kPWp3VxX1RTWxf+5tS
SNG3QnUiHgsCvhPlri2drKwF6DsByoqARFAufTn6/1OmnOdZJ2vq1gGAaqtLYNQ/
eYLIFwbkFGn5EsSUpvmTJxwa2PLdsuTXjwAe/i40vx1e5Gx29mHSh7vs1lQRvBnk
mEYAm2uciH8E5DjrkvCnc3sHv0B3cRMrMdlShdRy/+0AKyFeESsOo4/RRfMpGNlY
lgHmJSDhKmEh7jeleTxZASbyEl4Wx9Y3CU00tPZcDAlVX5kZpcuAxv8a3bLxGi7E
RvGnHZfCvw/uZ5y3zwIQv7hZp/979heD+vsNTLFyOfTsh0S2WRfiqbeh1HyMsu1W
L47EpLJDMlN7NdCj1TnCzkcn0vup3YLzR2WpDRr2az73ht4LbczgLdb//zjQ/8V0
02c2iKP2crvKnlL6uE4CpuSQ1nGWbzNSVlZveTld6qZVij1JsOq0day5wvn0tGtg
lHf/xZZWOE/Y3kOGu7xrAkqF61lz3jjQadnimEqX2DfsNwVnHM2fBBphclbmNKMq
LLaLbHh7likoIjF/gg28E7jyHB6FrkTN6Z7MUsCtvzRSoiRuQeJ4Sqxw6dgJmPkA
e6WOY1GQ7nqhU8Tri1AY5Pps1RIuE7zrClHPAunsmciuUglYmvBlxNHViCdf08c4
M0CuUZ5F62ML6iqE8h8xsllTOcDDYLdmS+/BV9FJzvoH7l6FpUZdBDSQ/MOQCHYQ
bXHyizTZ5wAn0ysR3C8NeM7vHBPe0XpVftmKhUPmgSsA9zZzXHHvoEMUG0CKBB5g
HSCgaV3LynPmD4igPZUOBXmoKdOHVR2cb4/WmJmWdkUrbQUtUrfQMDo1bUo09dqs
6kSOZTmhtWs4An5GJQ6/RAiwiSog3mbXBhc+TOIT9tx1HlkNWomIwSU226zjuOoa
UirfCAiOKFoj2lqGIlkEXmUmwGmiLef2sRvzHhGpPVltiYHWO70/MvDzY8zPtrFJ
Pq43Tf3dBsqVEmBroqFanaxeKZC7Fpe0Sf6GpUzhv6TVB78KozGhnf7BGI0nYE2W
JBeTs1xv23MX4lSs7TPA0IjS5kDy8QWB52IU4fIl6Sbl4GVi20subI8UcNzmW6wn
5J+7/JIH0W1+Jypa8JFhVdCuJwLrgs4U1+k7p32JNX8iRRoNp/TLZKTqETniWzWM
vLX+rgubunElt2xQOHvSWr2F8APU44wOOQ9UouQUs30uKZNBBSXVE3rOl1p8n6ph
/JX7WmC52nUaHlkSuGUTRZQ1yVdelllmv4KtS2qLnbDroWsUzLEfgeSYFbGqfT+n
PC9DJ6ll5FCRtlR4hOIFdjj95F8zRE3BbK9qA5N88ZsiLRAdv+BDVuwOxHxd3FIk
HdJpjOkEGu1NoTA7lJAcaOcG64KW9u9aMxwc4iZoEftJH1ofu0bxEcuxPxGg4MFJ
C3Aqczvcpp9mmnqLQO9ry+vwt132KjjoPrLGc2XqbP2FOKPxrmSKlFVt1xR6VC/v
EMCtWePAaJ1k0FwTafPTP0VjPc3ywCcAzrqMWtaOCNQZ2XyqUdUpAqjaj5vDDX3F
tk7VzZ4MCLHU434IClDn9txpR2cPfLsq2n6kfqR+b/zZgW1p+6E1PSiArpYoyxDm
isIPXK7sEikCKXCdKQ/JYK9bSGISNF1YYq99EPgVfeq77TFj9PN3ZDZJU0hnc5CN
WPFikCj70cul9wZCNF28X4QgpChQnXALl1hR44fQ58nG1Ifz2WAkF9yPU7GTaqNM
yNt5j14HhR0KJwYmmCDgCv0lrHOBK7QjPklDO4Jhtrtu2O+t6lb8Nxulf0tZzvq9
n7nkI8xu4EkFQllLOa3n/XJTdAVAwPl8W8bcgw7lG7C3hqpZOFgIvoTh/oOHarV2
/EJRi32jfvfFA6ct2Tq9RW6nXAjCUurKkzP4wjPPRixDso7yJwIuqM6touTbdGXj
7iBcwI/8Oj6FjsUpHX8DQKHXggB97HOU50kMWehKuab6qOu48VLHc+3Ztok6RaKa
Li5OUT3vT+TuE3XlPUwUACapJ00XL9h/3G42zLbV5Hlg4tucGn4/uNZhP4W0YyBu
TZTT/C3IqVoRzS7EM3JwmYt0UBlJldk/aZt0XQC7cHQWMHhwwDeBLWtW1gZLQ4HA
stA2cKvfGGqNKqLCiIOGXUPmzo1Q+NOVc1ieMvKQDlAVOTjxatBShnDD+LvO4nio
oUdJ8hYSzJ6S3nHsD/JWT9yTH06Do05YzZtT8BnOJqmS4rZYVElMfNrXXC0qUvN4
PIYRCvaSaF7dQyGrwbUlDFnYDFvxLS6UCqZGwBaD38MV+KDTVb4cKuG4PCM3RuJM
NfyjxOLmcbUOpRNq7ymT/HPYlzZISDzgfp09QTskq7Gl126FAyb74UWfdsBMYHFQ
4hGS+GE+8x1HNixSYwaZ0XwoGtG7u25AGqkwDNnm7wPe4rRyamJu606ZmjsIGwsY
me5fWp3G9DfhmatceVSeprJ+eHgeHxVORbsVPAKkaSLnyI4rumuaHfw4bZ27Hr3S
bHg645hlJQYvjUwVrnk/PZKBV81PMyldGhS0cfr57evUS0x5uqY88LHKqzpIkRax
+FQzJjnlATtGiDaMVxLYgp7+jZ9PEHJwSMfiVT8rn4zjrxp6pGUiAx9HalxSfjlX
LjNDoli8Dd5uw+VAGZw1fcCQ7MwUljrFgSFizuqJUW9IpNh8DwyqPwdeH5sZPYSi
urCtuhn+2zXDI/m3aJpvGHTXh7K8GYVlvCNoLz47Bhe3cE6nAzDPdxyjD3M7rVgN
9QyB7z9pV/IhTyFws+DGKyI1xV9oRa76rcK0cUthFwiG/fYBejK1w5LDBbOz5LBJ
GwLtZvGEG/K5fPe/TXreVA3DeQDbggKlb+OCLi5jMxOChxO3Z/dUZ9cyZQJEyXSo
5G7koAiZtMQZZeUxfmmBLzMLxT+AbNcYwctow3o3wcMNFOg+SVuaR8Nbh/XT3Pa7
fMvul6WP1AoezjWnntX830v/CiOvJquFWTC1tMLnUMnl30FVN9JBfRBK3PAnrMkg
QRwbeSP/mVbaTN5oZdpvJqT1qGGAnwkKNrP7XwyhTzBGGY0qttTRG4rPK6Rw1eVn
VtEkfehUM9GMdXkXQbqUD3mrUBVOHofTSgzzJzMeaqHcEsGa/nHXCNth784GStOY
Qd+s+7ZyiK29uZuxwbphXM2u79cE8qyO6Lv8RY0KNX/a3iqxkCvvGla8fOfxWcU2
W2Dlp3D6m6zJ8FPG3LEnIjstjRPw33a2NX6BB7QLbhp9bQAKW356wM0YOx1sORVD
JpKDpwCCIAspX1sRqU/Kw3Tar7t2TGVQR/Z21O2Xjhi3nICB5F0CQ/VEJqZlVMB+
0Q6T4h9XM6HHuQVUWMN2O3X8derSwps/LM/HW+zOiTfFYdBnDU4ZWSoIXucmh+XG
PqY4iGG4NNdPTzzVaB87IzFYPnlsy86gbcpAjySep0ycZDOcJgrX17hMnmLYanSM
/o533kDnGR4d+xf3TIja0LCvLvjdqM6yZl1SiNnrZCIQtZzshCDdv57/rLl8SU+i
h54pajvCI1d36eGhUdZ94DcLbYUh4qpc3bR4tBpqpz/WasbCb0curch1mhPHekGH
Z0zvl5fdN7hL4eY5ArpQksBn3kBga0BERaI7fAUBEtJPw89O3iGSB37oDy6J1BHc
wGR1f4N2CmM16CrN3/8vutytaejjxzcJXAr6Ve3upHgXe7s3gyL5pnKjOXXLzZKI
kfd5yz4AaE+WcHpan6GdQuextIKiyLr8pIjFixYzMSdWpZTGE36qwF9SbptZVOiv
Zk/7tgCApadkBc2e27PvR4m5GIi2HLQLaOyh14YMD1MlQdfbqAyn7cYDstGmiQ3W
ll5iY0BvPUmI5RSZ7pePNmnazvnLwzdsrlkmC59SwXaFjgsTwtgAhk5SOwaN1Jfu
uOKPwgvmdU/k+hyk/Y211qFu4pr0VXvdGLNSGY6SltoZ1xryLmKbz9GYArHnNkky
IKETQKie4dK/qtdDmK4n0uMifeLa3NgGgWsr+wV2uqMbsYn/8D9BDq7D5bGc8Mvr
KCRSsi2l5pP9VD/axfppvQ==
`pragma protect end_protected
