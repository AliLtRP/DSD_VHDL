// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
qy7MrqEYnwGJpM3DpKShJWpnxUwF4vn8hY1k4H8iy1YzCWDjftlHlOMRbmPx5K32fM0SBkis+kdk
pOARv0IVWT18SHKBYtpjlro8XYOaZGdRurz0j0u42N26pc8ZPSwxrR6fKWmE8+OE1CQKyKk0AXvh
3lrBEZkjWAyc3SMeWxvulSHbolp6IkzAMYlFXVq+q4IBBhvQw8yzELvlrCFjNpZVTR4BZ1y38C7u
/jxFoVxCJCDAp7CVQkgSytMqV/0UYOoiOyfv6zCz3uSFfyFXR0uyzwZeS+WOXL9zQyJTYvgejhHU
mDBa4kZMeosvAk3gTTcSoPdDozDVSGiBt4kW2Q==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
mwjlnWgxV8ZiPnWBUgxxtq3PJuAJqIBtT8T9Mk0gWhT3At33LQQ9xjx/tSMZwXqrCaJa2k76lRyz
7G/3Uu3tQoTr69iZxAL8QJWqaM3yjVodqXCIFC7U0p4DdbCfXbGYc/ysteOH5Ynq179udq8i88tA
MyfLVeHO7nCw3Y+xMQHC0Cd0WO1n3tVINV7Id4otN7JfxvdCS6acvDbcTNLA6EJZbOzc+SOArhu+
gExocu5xU2F4IlPCrh8YfHI3R888TtqOB3dk1xlz5w3iitA5jTQ7atOWZIi3kUsxgFcnWFE7qFsO
wN2X3Uq0sSYLeIC0yUzx0eJHc++LuUYgPcujnsW20lYTbMG3MQoIpNB7ZnzrW1PkgS8RIyXSQqL+
3lBStLVOSX8eHIMDJSFm3j7hsx+4qlkll4q6A0N3LL7wEb2KtFE7ht+ld5aEgHVCW7cR25qV3kxK
qCG3awN7FVdXHv9KtVajAmwEbP99jAjwM2rZwcmTdvZvbDHvyQX/19BhNXnOAjncL7ja/0eplNEF
2z47qPkbH+VmTTsLFcr0Mfrzy1wx2Gh3bd1fQSQGSyMc8XelQBpzSVzfA1r4SHOsRv+QgiQcxbIx
IjLTbDs18BIM/XRISeNwbMYHtWKQY6CTh6bvnIkielk4AkXjSDmXmGxpc20l4IN5VQm1EYuN9Xxb
7CcDFx2PdU4OW3PBrzzyFd/4tk8TKYyFp/rSPyirSbMIzqZwtN9b+eBHOEdu7bmNvXqM7otYot4S
eDn8ak4STGFmoZolqhbFlJ291L+qaSdLfJbdnVz+wAg2VGzD5R0bJ5+2o8jhRHpa114xvtha58Ot
Xt0mdMWOiCy1uEkO/phHNZXIlJWxeSV+IerAwtJ5y8WHYXPLwKtGnYZrnOgV+y2c4T76BI/QoduV
QKfPhb3g4XipC6qUEt4tur31DmzLJekq6qP0PjHhNvLYBeJsHfTHmUEFwv0SUFOpVqpUr8N3M12I
929lFXouj/mYcAuGDQIxD0u4oacSavto+yZPJPy2gU6DJnqXpJmy9wsLBdzZaGOv6+ON2bZL7J6Z
khSXq3rnJwiLQoQyckei2lhh7a850yIrvTNHYDcp+DLmbgq6TQBC9dWsfCPemUPVOARcSrc4XYKp
dlHvb8Xu8NIzT902CoeV7zPvWDdQd8W+nbnejutH58XGxHAOlPCMBESRtORITDVvR7qRVTchB4lQ
SvPNz/s4pEzc+DqJAxo4B3A9E8NTwm66SBBNszvxpT2bQaSq6Vw844MnchAHtOsS+iV/Wwb5/3Cn
NHoo5Dxc5cZbJ/Eq1nPFGAyTxnLQBDoD+WvjYxnFNIhjsmORgbKLhI3jz39uiAlWDMJzRYSa9gSZ
xnl91FoDltdC5fitEyOcxHDH88ZXFckiRVRM7kZgONnbpTRMjGEH6pA3sQVXjdI5jU/G3gIf17Z1
0MP7J5h/eKWQC3AJHxix72cb/gv4nuqZjuVc1TvZSxEeZ3MoZfpGFHeLJ4VqA7otHPo8XREu5yJ2
d0fsPExLLj+l3XmebDNA2RF7a91k+rngpEY5EFH1cqW4hgfuql4bFKeI2527Zw5dXzAljC9AbnZK
Ovp5HL/CLkd6b1IQR81NNcv5p3YaACTWfChhxRN2poQbWjhu8vhLOm/3IDx0ETAMoc5tQ0H1q6eO
cIo9xJ4bBdaUemO0hhH5eQkDKdrTH0m+opSO9VWqIJPkG/C40JI7qYrPppw/osIthjznQCMa+xH+
1a+bw6RfxVlUXn87qV4b7IANYnUQd5IIwGN8nXZ7F648X0nyYhs5N86LjfV008WpDT5fdgLjOgg3
1/ELB5zvG9KubjaKn1uNp1AyOIFkJs1tG/3e/yJI/yS2BJz25oGWWCd9pRbrQMTG972rd1bzdRIC
pzaCcqS48Bf8i+2ssKVSQrdNsCtjt1Em7fZ6c6ccf2a7gNTz/pyzlph0E7oJU9eZIJ9jxq/sMlZ0
H007tpmhdXU8CCtmzcG/jo8gieu3IPk4pU8be0mtnt2As0OZ9118++K1164tiULI7NlTEMa5EWLQ
u7A0i2GBkllknwnY3GdvhIWbCyLaDOZq/amlV7fLq3PJBxTswEABjJEmXbs4hqwQ8H1i/dG/yyhs
MWWhVB5q1FFTCCd5nydYoywN3PdL1GJ0cyiLesRlfq+KqZgrPSfSqpyQcdaiUaLXIvmEvmpdWnkQ
RK1XTncyNh3bw9QI7UExwSFhsKEPSyfgj712uKiPzUOS+HvfvTinZsYyK9pK/z5y5s+AkYWpLc5H
ObnnkxbgSeccebk4ncSSo8rta+daAhOnUfwl5/qxxK12TL15XzE9AvIua2GRp0aI3+TsPtHSgNPw
D1yQgGUBDYDo0wZ4I88qeAyeSB/pw4BpmpQXT4OdvVsZ9u8HE6EGV8z3ogZWC3iLkNOWtXBV1RlJ
txKADb08Oe0RXrquh/WzG8x2bTpHFXSxTrU37Vi9epslSaXugBvlJIxPC/UNlgb9BicOuiUWPqS+
9SQwtcZopeDxmIWatf4VbYBGh8LDEEBhrQ6hrLNVDCmxJrUsc56JMV6xC5yvpzvVIP+o4ZbvuG0T
KyTvMYcmOXYqudia0X19whSLIcrABwHw0vqZYbFUciv/V2oeDRh9RPC7gvZP1je2cPxInQ9lG9eI
gTv0J74ro4xyZubQUeDKsWbr9xCPFTZc/odi+ea3a+IjBgfpZHFHhCvXjymSHMN3BOidl8UkHnwh
UsH373wN/Umh3N9AeNG1V1HWlnXy9Y2o6xEYcN9b2CFB5EXg/IPj3/g8lr8zK8uEn2QloKDFMf3i
3pdUE226QypZr5revr70jRhp8/jTE3VgB72IeHYu9oy0m5e160s3FQyypFXe/U1z81Y/Prd8GbZJ
7XIWl3TrM9bCFM8QcmmBet57V6G4S2pwkCUIqDZILOg76j5/zLGj8RQncD0Smt4EQRcmD6Fw3yM0
7PqSIMEEC8mpWSacGupLigXJanIztH7aAcm40UYluLqKrKMNs+NtOgEXZDutDe1IDuJS+DhYyoXp
8z+UpIR8v/VX8BigqQu7TaQyCEbiiBkJ9viNKtCcC72vB1zC7XuoyWxbKbauo2k9tFKP3mxDxboW
hVmiDdER5F52mabP3C5VtNDWVBdhegBSk6H+bjUcVrwH579+8mEb9U+FoK+Oph8d73j+C0CtiN3k
c5orJq2Pe9uq3Ha+EMrf/vqAuYEefEtplL5Ad1ritAaX0ioVpL0e7tFoj1EAa5eMXMqY4v8yhHoC
jhPrf5RXAzXFwXf1GFCx7jwdOlbNeKM3zkd5mOljNXFS0MLK2uI3VoU4OpmZn6nYMHi5KIWzlDU6
pGHB3IWP6ax+4W3QWHBW6jeNOWm+qRhHe9uxEpqu13IykxX8eifIMI3D/d+1UCoYD2PvIdPGyPy2
qNhVBl2LXV3Z5wrZfNBvLP3yA9O+4Lt6bjVaJq0vSZC/jtRBqlNt+loaR2QkQTgg/uoZKWSj2A3f
+NPkGMxOUjk8qlv/rxqYXFOixSlbzgBgZ7+0aYtPwdw6StXhG6IRWVWc+0iyGNuzo3UBUUbBfc6z
5f7yoTiVQGdqn7IsN6hrW+n0QJOR9XOSnRr2aLEMLEoXasQ+Fq2y6uZJNfm9/CWEZGbU/e1rMeaH
ebtgG3YlTfVYZf39rH7zTHHa80ur369Sw7erfbP2dESfiZGv4Mhceq0OvkCPj24cqecgRjIfZTO5
4VaEKpZkkEcbRlMMQSoMQeZx2KsTvzoHfLENCz+TuOl2xYg5QfgTjwALHS4LXj16YbCKjEnHfsd+
hA6CMihtugNtke0OdsLI0gCtP9JzGGaEEnC/2SjNtRNhT2CPwSKMLZID1SfHuJLRYfoSxHnsGxQK
S8hChDmPXndZVFVsgp7twrDlCeTKSaY+wYgNDyY5c22iSSsr3lJfjC47gJfySsb0mjhK4D03N2se
1MuAZAzqWDz9U61yJuTZEaMpJdNfSisJkoMACNQ38LgwCZQZSxD30z6OPKJKeIj9aNbUP4UFRSGr
12rHCQDEemUjOtdbCynJT3Wp4A8mO53amhPa0FK/CeRuv/Gvrm55EZTHe+XH8K6PDkfl1j8Ptc/0
kqAylRPYeenBJ496KpRposR6OOV9zdCFon/7MEW+JkOnZUw+8wJcNyUpDy5yr+9wDAllNRgNLG/Q
5XyodRjWq5BdW1X9zHJa97Oqbs2fzpjrLNR+XjamJIrCieM0CNzKgahQSD9w3hNxuBceiLcmfF2O
UY24XBywcomTkONZb83G/bUlTs2vlJOBAweehXQT5lHhLyUFhmw7EA4JQA6QDBBdAhimPqgTiBeX
GO5JW3H2+J50ogRBuXV/A5QGJpsK6yoYbk2eSN5XazBDaLKgqqIHepH4b/CcCP25pa4ldZ3NUgmN
NkSzPCbX443TLRTWHgyOkENbrSHYQfZaM6boHrWUyG1yr83PMp9/shKxFVZrBEW1llPt/rJhviJ2
yMTKY4MGrKmA6D/j0vUAP1tsetAlC0RxPrDFgbT3vMZLI0JSRu/+BtdsAgaPV/mfni3w0T8oHIZ1
nIdpn9DMW0WvOqIc6RmDCvRtabuSovrBaJsMuJWmoZxKGcpDQVGoKpOp6LC5w3U4/Rvrjuf3T2NF
33hAc1aUZ4gya3VmOthxRq3C8YkUjxE+yNx6aQfxPkRklOZ31k3/8Kf4KGuiSTn+WruXeA3kcGKF
CLrpQ2UAf1Un5QHk+M+vHrO3w2GHcMAdH1+iiZUligDePGQj2zPubBsw4OF9CwvM7v03+b4ZqWl5
PM8ZYtc/yEXjK1poi94U3BVnyiwVTBPMA0n6rBPk+CcEhRYMt7f3Kbq4INN8Fw4F2+NOt5Z3BZYQ
OpPsp7gsxUxjEhZ9102fPGCnRculZYzC2NIJhsGNo4jUN91WOZu2nRxCaZFBX+xXVIK/3EnVVXZZ
KdejUK/zjkBZCKNwFrhROAZeoVJy6Sr1YGAcbp+7ktM4k/1UGTBPDswRaGC31QnpORu+voG11qVA
a1TH6FUmtKoemD8bKn6tgYlGLazsg8AsIrbkyrAkaZxQUXeFEz7EO2NXBP1iwRkTsqs2pRUKeIEQ
JtF0WkScDT3ETu9SQ77X+LACHwPj4+6jl92Am7f+4t72VD3MXBUFwaJgD2h/DPW3Yiy8zw7jde+Y
SOfLnyxdxpRLr6zvnzxto1GHHfWBZmzxS+biX9oWt8Rc+D8jmIayPaUP8QoFqI13fufNMksCqeaZ
dTnwka6c7PsF9Iji5i8dbXknjVHWg3haotjy13k/AGdVMYlc9FqQy119zh4wAHtHaE4r4YNOh3j7
XAptfporwx2ycM04Y1sjVZM8TBX3H5okIMCTFbXN7ewjK8Vtcqd4HvKb0opGpvvX/14vVd1j1YPk
veyEcTZKXm+RhK9Auj3KUh09okwxh42RxLWs8nrRFsZXTwueist+JwTHNEw8kBXgkylovk8n2Nlm
vFvS8KKvzur8tRR0KrzuwXk8RosnmgLd0lbyDCresd+tgLhcrrtnBf8h24AA3ujNpXCmwlBbo73j
UtyVTJuF3gzYIWtmltbI/yiYVnSWr2VaXQdV3RZooOlQI10IsuGChsoE94vn94vTP4GgTCv1YBu5
BYKoskK6Tjq+YGIGs0gztTgaIbGh80Yqcr+9Hcc97VF4RaX1JRksvMjdV/gk9ksK0sdf3VIBZfqK
txzDFmjoM8jb67u84jSwwkJmEMZuuYlJRxWudKcKtqpkygYmYq1gxfHrPYpui1f1famlwoaQJuKL
CjQnV/AClzoWs9hkL27hz6HZ823NEf2P6L60OQrGq7BO6BisYd7bZu5f2yQWTM5XwwRf030fAQ4I
nGPA/Dt9kJB2+pftguTABbbGGqQD3m0mDAPeLKCKo+M+us3NPTo829xCEE+9Y3w18COjAJb5sEjj
yFD3dCtoEWB6Gzkx3FRoOBVt+QPd255cK8g8W6mxKbXdeChIthcEQ+6mESAT3IF91vKHSP8u8DZu
gQ546+bLX2jOzy6ESH+rtPes7sj44ZuUIYCXsbmvHxt5rLdMbRbFK9LOq1nMqW6gA4EyGhRrhmMn
14Ck7xILgJB7k2/70R0sf9QY61aHcLXJ5OaQm6EEpXzqRMhDEegPf9YTdXF27UvF8D2L8gaVGKNX
ypBcPxswbU7U65Ng1uBNho7y2Age+kE5B9P27IUdAeiweb2S3QSOG5qVSJNqjjbsKS2Mx5TKXnkH
7y/XsIJcEENAQk9pJCx0Qr36nc8740ITnkeb/PMXdC6q4WYQSv4qhwGdP8ncd7POSVXYfZXotkAk
fSFuz+8Uu8IrikkbnZmI8hqmuYFhUxT2GvWSwmN4jbWGZeoWJxoecq2K7tyClK4suQBF/oNC2YYs
OnAfcDUjW4k+bK4mY1H+24jjW2ea5XRu/MplX76dU/4GkRC1QDCcX2CvUw4LbvQxLXkupkOAuqKP
CV2XlU8cDzfEXsZY9jlWdnQnnLGPA+01RtrXdURZkdXfnNpJooTbUsMtggBwVZQvrQCcsa5CLyeZ
2paZqrdenJC8V3jbS6tYxSMOL86XWoTuvADhCQjii0vcqUDTCHQeMK2kI4bYa1ugXtT+JknHt4pU
MfWecijR2WgzaeY1DnALS0KqHGB50X5qOsu+X2nsUiUxz6IM+92OtUb2EaejSegMuPwshIMlOT2o
XBfiT0ILrbIEaHVJKUQcAv8cA3Q5Rti0jmUS6djObvUL/FMel32/BDNW9Pz7pJadwBQ+k1CMtjBs
MQzKW1rU1EdMJ9MuIpVZYhYBgzinppZV18Er7bKfnsw5t6bGpvJxp/FbZU807SqzAJV0YmTyEkYM
lkAfNyW49IKlgX85/ka5CMwGdyZYWRgYORxMvAGOJMILNcs0PHGyOso/A9BiFe7rvwCF+VYsNr+2
iX3iqPgwJVn6jwlRwT4BTDtUK8aB4XOL23NZipkf3Rs5XmqOsWHMrT3u+jSLqjWkDwuQYQdfLjMC
msVCCZ+q0I5NteOLZLzr3Dm1/DoImNfMQOMlHBW9ExanQYkFdbFmj/AfSC3qFCZ39l6WGhXEwops
MpCq8bbldOS8JBqD1nPCU+M6YpbtwfIJiH6oLJq0b5V82DQUVGyRBFBTXvUEodCY0il57xnRr8Fk
d+OK59sJvFsgIPh/Sfzykg2Lz5XvsWOto8S/MutvQ88Z6oQK1VIYbAl60ftZB5RqjZV+xb6uOo9T
26i2JUpPUjb1GUHWkJF2q4ebnzkvZZ71BLH0wcxAIe1t6RAWEuxt8KcWy7WQcUfhZkX05DmJrVoS
sCcn5xljaHs1WRrQjpGHK4KoPR2mX/+Q+4BnidJB3I+aMHqmREIau1nZCFTXoV+oElMkIXLM579r
2Ywv8At4CdE/nckXPZkSXRcNw4THl57aIUT/OY3sEDMvs8ERnLKXvZlWa8oNYeLCL5KnVCosNKYN
uHrJaIRa8CeIx7TeDDjeCTLWyoKRJEAHiajdizq9FluK47B7GAzh78qe55uB4wT+bbLtMphZ2mKK
4S5/OBP2fdNgDF9OJF84o9wWUbdqeHlWWAICHCzYE2nITfyq/x56eM1Ch3OcBiiRucSVA24fj68p
2curDxkmSpu96EMYj30//ykwf2h/4iXtv4VcA61beyulSxL+mYqvQ9YYTowhNGcbm0MBIpARTJUS
bUTW2j0xppVO7087O9qnUo1v95GJa6NltP5yi8N2aXfFKOZyfxRLPzvGwUGEbn20Dr2POEAvPEUy
YQt9j48hviOyIb4t1HtUPQrt/NJIPN/KerjXrKHthWAH++xnRw8oe2rBx06cXzvUzz7n8JdtvFt+
4yN4z0yLmqboI0iSTR1ef8BKqdxiUsJfvimWdSbHl0WFHpqCHAen7AhP/EAbv5Xu7kJsmtb5kRvE
MyL+T1tV/66iDuefy45zQIUbQNnMgDk+unBy2WBixi0d2TmICLz2IEdej6EHHavOLaJExZMcOVAG
lXRLx8BKUlzm53/YVF8OCVULsNtY68OIC90EVNR4fC29RI2W6J2QTfkVwwHDuWRwsNm8+2pU44oI
XpXoBUMG2q/ZlrxndVrIn5Dv9JttPOjjZKIypPO8PzpAKTDAuLV3BwJzjEXCJ/kcM/CqBYURGdqE
TvFJnGXLzJksHYtXHCy2vWlhaGSH3Oc3NNuUiK1+DVplHfGJfvj8OBwZpl7kelvUSg4zEewqEL5e
NU99S6WqAzdq4fTzA2UaSQlJC+e3jZ6Weyt+5V9E9Qhlt7MY7tAGTTLvjGBSvteghCbFJvt2y0y2
Sn26fQKxyy6QUbBj2o8ZWF0En32fS8AVQdHA1AxxpIzaLStSppHIAtF3CixobMGseXqlmUSZQMAC
ZM5crtHDwKpzKl5PuAUJ+Z5KljybKc/aX901iBJqDY3v/6206Rqxt6X8X/hsIU9V3z5fUEOyjNbE
mI9NF+RGWDhAl0WwarA6FD4IdmdSkXIqS8ro/9zNLGjIg4n58qnpz1JJ71+Qsf6ykfgPILPogYD5
rdEZyuTwQm8a+rMABLGKrzZQxwYe5IDcl7HkrAYobKQNfuhS0Bqr+lSl5coAVYb0XcXQ/muHE/Dy
VgYPSZaNNmzjBwh3Grptshw10bixlUsMZAlpMOzn9chjEPz7aj3ZWmU79JpQBMN6v1RoxQemEV27
lSz52yyQ76qTH14PFMM//aFYMcohYYAQfTGK7NieOWh6TJDA4IBA3oc5YzJkQZ7ol9zpoD79h7sq
/jpIG7Df5zPRdMf+jWu7odsu+aefnVzQS4IExPUATXiVCYKLuaPN+nWs3x5v9sa/rxzCpewMm/EG
vEX7pHXDHtHKj9EEP8TUe1yCTUnOebC1Xt25qoGHVvM5D22zm+2H2U32Oq2/04CRBWDG4NcYukk4
FQkqB+1mh+/FI161xTgfNbPvaP7rX8uIwKx/yCWYB5qPtYJp9Vln4upWfqhaXypeoPmKnLguWmAm
vt5YGLLS0F/fZXu5UNckFidGL61wL7rmt2dP5GpYkrEWoeXk7zKegQ0sXY/eGDvaHFPATVZzb2N+
g69twOOvLl+18dyW+CDUlyyESyqgVMe6cF1N0rtdOh9fi85lILGhdpwjHzSpaYMd8psR0X+pbnv9
hhJk5KCkJlt1O+vb1zLA/kPa9QxVdf25fYcxXvJ2NQtB7a9bw/xpAGSBeqM+YTeA8vy9bljHGMy6
2vOk7Bg4LCKMuzusclrXt72O8E07TZbc1d7EiqifOpfyvhrWYfBxY8gGHAXEkpi+ayVWOUvUZYQg
QPWciEUkNpn2TtP1IsfIHC6EbfdEedOyBvUldsGQfZrPVxyWwK6afYAj/lV56oX/3ZHsB1Sez3Hb
ydXV3FTICNsHVIeLJJd8crmso/ub3DQhJq9JAD4gsLlsC9ouojYz+TylKfR515TAk6uaFlV5Kfuy
o5JuJEMsdTzU+cr62GxXo8bWAKrK5IkLYUd9Dc2BTsYz4PhXsjyM/YCr44txaMdFkh541rHmOLnn
pZmiExvzB/UlY69Gop33UQ9iOxGDB1PGyNIAp6jloyAbB73y3Us+uijqcp2yNE+L4Kc5iQC2+ho2
DF7nvZG5KbPehaH6vUF+jv30zjT5ZMAjbL6d+gFcM+iPJOoLbzhbYIEpqNemzT6JB6lklfZYDMWs
/hBVuNNQltc01iBhEdlqVGwfBA6qhhciHwpO9JSLcvVD+7UdlUMfwCtK8rjdDOpZl37Cvqow0MkL
mN1VsLEaMGd9tZrHtIgduZyLIm2YadWKLmFloHR2p1LTeyNZJ5Ro3bBrT3sB8cQVpCpRaO0Met92
ts1v6I2J80tDjKifRv732QSTrjYwv/jTEz/5AMswsv0U8SiYPdLobaiwoqLiJWURQGLbLLGok35E
UnzSXGiS1lCSe7Ntg4btVoUy6kzHPKtRh/uCwyIwXSq1fSWMt/T9kIUL126WZQdQ/IejAkQmORD3
VlsW/Wo8oYhAo5YbDzIFJ1hWrhnxn9ws2yXEL1gwnsOA1DetzJg2TwTnm9JO9B9+FrtN1PyRh14Z
O/i+WfhOAxGFYFNt8ageXmwsBfmhiTXJP7YyDr9qjhT9UmRR3emTKKRtDOFGNR2tx2rR8o8VCCQC
ztAfL9/4bx4BzuP1lRHD/SCk9GEn3CJnuPt35VMkgcRJxTdKsLI+00Q+OlbTEsp1RkOXhUSpEomP
a/IfLt5xtgUVs8nog4vtdZEMoSspBOp3T0ykMVlJt//aUiUgV8VpSOXJli0UzC+eJznGu4AEM7Cs
iBpp/Oa868A4M9OOBgeqYrXxPPre2o6ggOTktVxMytF562qOPPTQYMSjq6mxVyFE8WH/m3pJjHnm
x11Dq/bI60mwj4WOHqKde4rgV2JjjvsOcgYJdBcepmueVOb1Q+Kuf1gIGibGJFNkcR/SuVHOjj7z
QDMvtturOnXfWj1OhYvY+70PByLq6EHV17kpLvvp4JEIQyauUVOWBTJy51ZmuddtOEeVlGM+fuVN
XEiiK4QUTHvKDiCFxSOg7f7hkIi/4GtOBPGc1paDNE+AUvg+I9OaaP9pRN143vuR1a+sW4+wE6OQ
ge3xR4smFtP5y0DGtVCKeZ/2vHzG6J6yQjqj+T2dvMqWMmiXOk1KTQ7cxNEcJpdboRueO22ROymz
MD6RtN9J3ONHgIcUdtDV32EQIbCfapSCpVnsV4I/NIwYdppATmymRth64ilz7coTsjQfxjI3/kts
0vcXl2Y9lHUykWwmBmjZ0rKf3hRfpgR+ugK5+2A7ezZ6YzObEiwukIO9aR74oGRI5Y4Obtub0quO
owzxkmDJqlnTl6cdyh/v8HZ3eRjzCqUb6tc6F6HyHLHqskPVvbH3ER05OPqygznJTtMlhJ57x2E5
6MKb7iJ7tZYZhRe66uJUUMw6QNq9ju7HtyL6v6RMe84xMqATMCPmQhHJ+HQ3CwFe1q+VwYKACuGj
WDJPQbY9q6yMrDtIEynk13YGcL6QixxEkQrgGzivuO+9NSJ9QBl/HrcGwjR4OkCOyJDjn1nNIwbS
TBdhFFXX07KmOgtQ1Hkl3XX6z2uye2CLZ4Bn2LJJHPiVBiXF/ww3pCUv3+yRQPyVq6IEWEoQzYFT
5HGZvAdu/zM5pzb90FoLLO8lCNfhmI/57DIFBBIddB5niKWWLOAn+nI5OPi61SJT7yVBzZ8GH7nu
Pl2DscX0oittjcP/y1zNbwiIByCac1R+BxNdvFhzOstuA5zQksvXqfvv5BV59cW7GY+QXY6YSVCy
FrV172Tz5eEvcPEkiupyqIkHIRflNvmstBaEKiM4AU4g2PhkJvlrdBRV0hBzDsp5HzA5aHnA/Bg7
602VeW4ags7Az6NsOWreSmsfPnmnb6aPfOyzliKfluyA3ikT9yQwF0I2Lpmo+dXimTddNZSjTkWs
QtnxbOKe8nA7sd6bulgaldylIxYCAXm2MEpjwJ2rIXm4SZqn9OIAdZ4TBmKmo5cQ03QT5HVls899
s3htZlted6V33/EVMv0KKG21vj9Whi/JmWqjN9jlh7ih+dVSZyko0P1AdRVICwzyPeGkayw3aroi
fEvB5qG4zPPI6c+op8olZqYjAchGutxtJYLt010MtfsrpBuDvC+GpGaJyXYAdNHueheD2h+0bLXC
UnLwPn21JNv5eNEe+N13wLp9NVIMc2CnxEm+JyPfj3qnTh7siq5ZL3ddnmWkR4NuvLQmC5HxvZgz
7MRlLvpq0etwN5eAUEIg5aOGyfNhp6Ms3uaUd+CRtJ+/IYccTipYqVonyst/uJx+rcbT6V4kUqA3
nzVXMjB35uIe0OnbNC09gjoNKCWIqPjECwbv0M7cqvPd3p3b8I3NkvaJU9mNWMWzZJVey+U4VslU
C5ixcZQuUmw+/FVw6ktZuWTVAhgkuSngbWR/zSPMNMGQmpPD5FH7PI+GAMAwRyi7uuwIM27jDTMc
ZeSVGtnRwpOHVimek1MnSeXohRPzOUV+mT7wCg7QhXC8E9Gj8MqgSkHhpMyAR+0UaMPweSLhTkjl
PhjV4yJfsiMHS07ikY5e+NBC3pfjIkT7hmtENgoSBEISGFeFbj1QOq7O8sVIv2swRWCm9PcViOrd
mVfJ55GVEzn+gFeMNVXwA0PuDn2erVLKAcQKKdnfbZYsTuD6hRgdxgjrOw3L/RlGkK+KDVSK5KER
QwH8Rd00M+ejYcuocaVXHNwiSfD0NmbvmphulJ2fliAefYbHXjq4ADwJURpa9aYLtzFAjh7+ODyN
Z0TvIvSkqAVa/Znx4bsO7Xxh1LULIxKjT/JZofkpTXkmwcNSIWiaPTuQtHMaWvikcitlpEHoJvpW
ERCeTptNPdfbMY4x/sORpMZZ3hFmmY4vRYF5oOVPJsn44Z5yR8e47WvbZRVCrQdVzFeGS9iLCJiR
Pa4XL98wHF8Sx3+8F40oLuM3/FAvDSboBDYs9y+7d/XX+otoFbyf31nF8AonRW7WSAMaewOlhCzM
2jRbzn2ZmWtvaJE7ixFBcNDyQUbUUcw6kkxuGFsOdcNebzkwtSi2d87eclFPy8MDr1TNT6pHTROl
CR2aFUOJVelttmgXGTPlcIbE4nHdA6S8WeporAHZo/dli9yExHRYg2WHxMle71W9lKKYakp9GOr3
GMxqYr124mT6RIjF0TqvNgn28fexMxU1JkIwWTFVj4UxgxRiDgltIZ5+p+wr5kxhBWoKZYM0WOuS
HmHkrTIKjwZis5I/TMHfNhCKnhyIvixVMWXXgu2a32hx4roDIdiBw2tk/5x5+pORepA/hay/BMVu
x6roGVAZssPG6SHJMipPv1S68QFZX5pdJlAx93JMlxmzWu3F9dg8vM9o9rR57wAAKUvKQi6Sg6V3
Vr1VoXas7TBo8HG2iLy6I3tiuIiO3UMkaN+B0FXuMIRml2/nnXcZNcVT5vy4PjzKoeFssCh1BLlF
9EcuEbX2bmsqjFr2HJ3VPWdVgOeZFc9peS2qYJ2K1dk1MsxT5rIYXULRspHX+MID37/jpsctdmDl
A+QCwRru4dpDcFQr4tXk5NwzVS7jC0glrxWJigNdFP/aw1TgAhNYYXtCg17lgvg4DYsFK5L9176g
H6H0B5URXF4AeM5xtHtoqqLU83/mygB9Dxj56l0PP0ehiaICZTOI2qFL+UhPPTlxnNjvViJ6X4LC
RW6OsTkNIH0Y79+BtPPG1WVo1rT2caxZXIHftEKW+QvIoMx0U/OXfDaHsPwRa7PqgH/UcPqq5g5Q
aXT4SOgYa+pwzBeaXqkdSlTPIOmIwZkZ7XZYw5eM8q0CT/n/ZrmX2H3f2vik3XKILpbDoVLxxnEt
bh7wG85l+8iSfC7OJLde7JwH6sKmVuTrMraeZJw3ZM82GKQwRS/e82mFeym3AVz+wVA5kU/JQ3LM
i3hgY86PB56GZE3Xa4+f7RySpf408aSuiYcl15W8xn8XEjmHFpX0NlbyJVzMTMj+A7669NE3UTkx
Olxu6ymRKISt/cCmcZd4DF83nMvyeebjO65t11kYvhJgw++oA3PYV/GG3m3ppXsPp+wYmE8IBWSR
K9DlETk7QpPpUJTjXwhl5FjiGrDsabp9q3t0AWHR46bhIhiZ9kOERxSMnhwFCrGCMwMaRnKp1YUg
8dfBtvjTLJVIaOZrqednngqrV3LIrzOsaJRaseCs6mzlQR498ByQS+OOuAhaYfXZTbV3XfCIti2T
FmsZDF2gOPeoHiGISN2XtEt0A0MR72LWuQ1k5cS5KrNnAh+ioChjO7X4QhnGdt1icdRlfJZA0k94
V/alghJq8KrRQAP5ky3URKHDM7kwcqABmT4bT1uch7zR9B9kEPX12ypWyDIR0Giq8tgcqtOom6qz
Seq0OObcVr5I60mq6IOLqk2rBWcvWd4QYj8uomF10tGf8fWTZTlYl/Wa8OP8L9dRezdo8cyuBiAB
lpKoUuJ6UFyTVW47n3Pjc7J1K6lbbFPVXXNVGosv1NkY+m1pVLk2+tPAof9SRWwfNPx70AlNZzra
Bud1NGxIs0o8jsiJvwcZ8Neb7yzCTpdm4B+Ob39rX3v/zelwARKAlQczmKNHOFxhrmqmZEMztzP4
urSasZMiAD8jaqYX6+0Qp/FR2HBqsSlcsTsXDuMq/dtn4P6dnCM2SLvI6WffK+dvo5Hc+jorew/0
FXxdH7LCRwpgPter/2vgl207Dhq9AhxRpKNkoorQWseWNm+2+7ndVtUYMEY0UM5Ud2E3DOEjDRLq
M6Gi27RpB+ovKj2YBDHb49phbmLHFeDm/7dXZewf5FbThn9H+7oDephO++nvlFXSxrH2La3EOjDe
dZQom1ErEZDrVFchEsLy4HUMAHePFTQdF98o0th3eP9U6omydNum1D8ZL3LlgvhchfhyAa9Bo2K4
feZeeJjMLbm7g2YrM1U2gyYupvZN4CMOush5Fu0lIFKIrsoQRmNetWyaoc06CWplq8fPaKy91dEH
NQhmw+TbAmsn++NbnNFM/nMrTr4ko957rlR6ZlEN1vRwiLHsQ70z1yx0AHWYAo2VNRvACKH6RncF
JoWANhvPG0W9lDyTJwf8uEK2wO9w1WpyRqWUs6MbFksTDOI8Nut4908C6FeJ/YG2niBP1kLUEvHP
3HLYPvpvspF3gbc64CO8EV59YA5Hd8aVZekxRjhzDxLUvuP7EXIUrZwrMMTkRyd0tjP2761u7foa
e2FRMnzhl8ssWvZqX7WFDMosz0fEibJDKlTbA/qaqvxpE/px0YlP8/UHx9YhU7kHeCbza8pBnJCi
Xs5aJJYp8m4r6c74h3++tKAV5AkEXWULVGG0Dzv2BIrMtZpcs1lnb3qst74Rt+AJoH5dh7JX/ljL
B7RIIvlsqvtR5AgTd1YZ+W1zeM057X3XVDxZBH2YgMe+FNSsYg5ZVrvzlpTVEAap7YV5yCKRu8tQ
TruaLjCgbzTS+EVv2wUGUA96TN2fo42M6Y9Y/bMLkRsErH0BwPfDIBkEBP8t5u19oqbFXMGUXi9o
5O9SEiPNR42jS7/p2RcK9fMoBXPEirN9yAre/VNOXbwTLn3F1ummJx0OYzFx3zvZttsI+r9MlYWr
MMxFoVtpxglEAhZw6VRZUElL+NS8PS2fJ1dTQhHJZLKE0aEaIV7xbo10Ioz6/yNRaHod3DiWCPgg
Qbf1LRSHKT61r07DSD3B/pqsE0GLUvEm1ySv6XulzoY18mUguBGcKD4e7tppUFUB6WbU5WP7NA52
s6stZqnapIh9UtLzO8Q/hY6jVyreZZn6UapVislXOKOYLXttoDZyH6UTgwtNcyqCBScMyKm+9Kvq
a2An95QG7woJ2yYQwC/dxsjVvRUXZbcht8N4H5HsF8Wp1p5ECEVU73Nt4+Dxl6mk43BrLBjmD2BA
c9mfJUQExVxSPZD6ZhSuB3SY9UTj9/LbuvMUoOFJWPcskMdvciD/hCFG5Um1JEHp8F9u+Qub0pez
hazzX3ZCgdw80Vs1rIO+o3vr/wsw+YUUhPvNoKl8/3KJXQVbqETiRdsISrFcGeotiIlVJ1kPVFRW
bhk3m/IvJT0DV226v7kGIzix8fWvh54A92HZWlitpjj6nAWNI4ivqHOgSa6vqIW2uCgKWWBz5TBM
GJ/7iN3Q+zE4nOXGiHQG3qC4ithp/o4TosyQEx/mxWTjfwKOERx+oAdATn6aXQCvUGb8ot1Xercy
GyONGO/X+AFAjoGOhaRTTEgzTHQuKS7NKDSctt1veyjC3G0OHwjuiupKgz0Fjvm5Zyo76n+SH1qs
Vpk/YHxzr3gUiOuWzxDlLJ3NkVGhkjZjpcH4+i4FnCjTB7YZu6TpAZ2bYfP15cBi+On/u3fqPR+2
IniLPR3FTwKKtMQDtdUn3wl7MUI/463p6IGjC/zduEYkFodtpHqgK6NBbZPUbO+rnk1cDcLwUCsw
J1b8PvYjK0+bO1p2NzviDKleS/JV+vmNxnY6YYmFY0lANdPfNIa8DOi6ZbuMEOuNDCpQV9mMFinp
Ekk5Ep9PUK4f/GHCOyGVyik0/MYzL3Krc2jMX6vPHSU0dVZDEJQ6M77i6sQkymt+kqKus7DrN4Hg
vcjjaQ80hqupRsKVkupi7k+1tWj6Rzt0vkEAssx/oFpJGkYloe4Rsw4ESdEeixOsMaiNkuTddksz
TAvy190VhErLsCkz0BQpyj6KPfN6VDXNiXn1yRldBTJLe1olgkPy6vRrxSPXVOO8wwid3vEaJnQK
54rDWzKIf0fL1DfGBZjRvdN96RaMwjwyBkTOerJZ8hpBNQ1He3DKxJoaWFlzkcBf9aicZfxUc0Lz
6JiTE0hxbMhiovqQ0Q2LaCCvucmWr0o3kx/sliu9ln3baEWijFkwzx0FiLg49iIuVn4ZABqjqgwj
8WdXyX2CH8oBuXTMhTLViSL3W0fKe+5BUgRIuis7w9+wOyjDY+9r0JHBdZlfGGr2Wgq8i/hKoM8d
V3X7XiYpdKSY7f5AI3TGiemDy+64/WPiljcFMKtXxXnNhsQVX8HbWLxYmMNsxxccIWDBp8TnzrqB
R6jUO47MBkag2aQA0+P85Z9P0ltciftqI0ZOb3G3+dI6ZhmUQWfRjricDb0cgCgUqfbf9UVV8Yh9
e7cbmC2afuhElmx5zs7WSZNc+XVaFhyEamleKaghsGNY1NXP8ktc8CN3vE1MH5nKBDRYvAPrW2MI
eU+7NyDFKBCCejZuPKc28hSdz761EJyF1bKzZhP2xc02q6Cp8ZiJJUup9DJkrk+FDkMk7crfG/Km
RyirQmYpigVt06QEMHnw91uE8vXDedSuRrJzLkrOKLD+fsVg5QGD1hUxUSy2oHueWH7GA/4yZzUT
3fQS6+Va78cuyj8VvMYNEC6WGw/YSop/lRC8oF3re6Xv0GdNhhAsDU1JTANOzm/nw1HnLsZzmUXj
zMFjn6xbBqNOQtdeKfd1t2KrRqsrgwU77+/0ng2Y+ezTNRIw3DE09csTTF7Z6RlzPHb+W622wuWz
ne7AG8tDmuWkzK0NcYpakGT1XBg+kObcOVcjbbxlgCoQ078FBWdrYj6qJik1PI3Doo1QtKXzTOFN
D9shULQCkXAaTTuEoyCohUnikZ3Mqv2G7mpV9qEKmh7FzITKgjNQ9HDCKrdhvAB6VyXsVTFVwfkC
b85g9TB5QTp3iCwicUVAPsIX8HxOwdcoomW0N/oFw5JpdoEA6FDhcUPLiAfgyNEyCOCfIPQ+QmhB
FzjTzv6Jhz4yrzogaEXeTpknOjnLEy3q9epxOloac7UMyt0aKYcPU85U/tSCWXNq9W+F7cwo7l0L
2OHFS36YbL5vxaJU4EZMPrPVyskqymDy/v18HnhHjwdao8+4eS7cRdvtEa1wHcRheKUKEJt+ssMP
bZJiqPcqK+dC2JGXvjw1BZ3JoTPEQiko5kBqzfjzWC0vHtbe4DLBHvbKvtT0mC/2yBpPyU0X452F
yFqP4EZAzXJKCRFN7MV3KueIrGWlKLx9bzHzCad6sEorgwhsVHyJouJ0vkPyuwqvijFzrCFaqQGE
GLWIRQU7Q4iPEDv9MOO3OSg9zP/Jw6XO3poJSRJHlCy6MKZiS23RMq555XjEda2zqK/w/xm+7EaB
UvTvI0ynTCwNqO8y6lSOeRSBRlDQiYx8em9h9ADiOJ7/FC/GOV36iRGRmBSYwKrO7Csynbk3FaJ7
NGWqQ10rUOCjIo8MNCs6olNiDQl6Y5UdSgia6f1zQ3f5w3cvblkmyMBugYEtYNSe52o63RziJ8TX
NsuCJ8a0JnZPcN6ChJ1tWWCasz+TUnXmdEViUPxmd2ns1wjA6zdO6WFDN9ZUFisD7fdeTSPEomVE
JC39rGoMsLBFoHZrorTRyCG++FlpSP7jVD2ltIrmBXoTmJApp/MawqaDDtGRK9hZC7zVDCwGNA1r
ZXzUU2rZXL4QolfVL6wvEXAcrXLxl9okvEo1IwWYLpfuaij+I7WE3sBqoHE2fp2tc3IE8cc+/NKk
CYbrk+3NKsEczT2x+vIC+PloP5sy8pUQg04ulFVdPG3kYHDLb4Npq2gQHXicFNr2yhOnJtG7LAF3
RWv/OmCpOj8dKPczH4X2cZaIDLT2+3M6n2ybqj/Irpv/PaR2nd/UnSYnBKMBTSw5QEqdTpAnfTRd
WCaAsmoStAWF20sJxHx60mfI6XbOyja86DlVU+X1k1jLttfRzZ0aBPkly7UPL58DCL7JQxW9dw39
4ZTyPNIGMHtJVV83IfJgM8Cw1thTj31+nHvjpXlydduWbIkLkGLt3wcBN8ghxG/5KbUrT+Pdy2hw
Sj+2ZLo9Sb2cf8g2dHdoIWTHyBvMHaFzPfnh308cmdhicxB1fY8/APFpS8BmAWUCWa3S2lKrHfLO
yNjiPATdoYo0Am8tNt+xidpk2v2YCAxwt3G1ssvZyhwPQ52mVkl4kmr7MCttazccWQfNysgWRvMZ
J/WmfaXhPEUFKD6Q1aAHbmSZ5N264drHjctLpXdYJBMNpWyC4b96zvHYSo0yArsXN3Iqw9qiJVzC
/tDMDhqCi85KhJUHxqmXfYW3BXheq05DAgJDd5W8lic4I2SZSFV4gKZ75HuTKtU/msSLHGK26yTl
k2WoOdU5m7v7iIFCdorxOjXxYtvVby5LoczYX9iikuEDDoYLeZOLHLQoW40V9TmMoULZuystbthP
y+HfLqWTbNTSXK6wNYB3c8mpTrjt/yyAdTnA+allwTFfMsemJQ7+P17zO5nX58kNQIqp0JAwtVpc
AdmAY7hfDhWx1HPb7jAY5GZrmDbODvNveS/AztHB43hSk/HjhunTYsbVGj7u/DW1erBv5bjg/L0E
eC65BGazSWk/gXGrHkMWW/OM4M11SHeQWxvhrCoZ11aEDnvfyGZCx8QShbNdTObd35srUZxkKyEz
mKtJbDGX7ZBvi8yCpDaquHsLF3a8Lolu+TG/hQ4U+a6eYUh3vWcy6L5bEMMowIpEdNPlxTeUVz4Z
CYTS26MCNxiSVvaKiRfy5g7YBgrCkKfZyt2k1pnDiKf4miasqxtsPKiOzLvKJDELJKskVcSkZiC/
007hMQxE6pGp4WECpQrsSLIaJPzbY0caq1V7HnD1cHwYEIIpi+uvK9m6gynAEgc0febPT8VMv6bq
d8vuVH/gB8cSdfOJ/yQaEINehSnfD/rcXXgHT9gMctpis3WdjJFpNOk4Nl0WjuMBObc0AhO753d3
HxFRMK9PLubmJ1SwnH8khasH8QRwn1iJifUSeoEIr+Icc9auV06H20DjEOigJxfRLTX8h4TNgq/q
0W4UhsawMcLMdksTVsers2ayj4lGnvC4cGv5vHGnCIopBDX9y5DLfhzm8MyunqngBmxcQgp5+/zH
vTAAcXxa35S9oPZwZZOOCnAP2Oo2EKMTIk9eee2KWu9ipEgv9qco4uBRlrFQZVqD2EfAECm3t8XR
pqT2550iCYOgyjFzk7J6D8KgOiWfHXuK3N7Yv43TwVk1SI7XigeeJs56BDgsl6QhKrGOikwQsnsX
NupWDvnvvO8zVmXJcJ2e2RVN29/sndQqhxjlDVYFn7bzBqF4GlOHV/Q3y7IN6bJuUpou74EGHaOc
aE1k0DA0hDglUSIOS08h9vEEkf1gATTBUtoxWApEzEz+85WWdLIhq8LUmQi2fY3CAncm6ue0Zy0M
tUkYCdcD6IS00vS3CpAghUoIods1ky4XWb6OC9uYpTLHeSKdGlArqv/pbDllJj9bxie0pnKJby0o
djhzygaynHXWIyUjfwIKFNjylFpKZsQBhA024wuTdTDOgUnewnxFZgixMRwGGEoshwYQM0xNMM0G
iIZh/lGQS6JS4Di6vUCCPupQSbgrtBWM5hnP34E0sifofMcIzzh8rTAPh1/vPksM22vd6LsqW4eu
HJPSzhOWBaXIVnHRB7puMppRccPPugrlWaCk9j1zJ8AKkayfeVtIhsgoDNKPM2+rZ08WEVW6ewkO
W5PhLAac5vm400cCMZ0nnoTy5kldinjt2CogmKdjHRCA1GFbHJt4m/D4uRzlg1xE/Q2LqFAW6xYb
PkUXqQM1rN+M5rq1OZ22eg14q5wfmFlhob9Z4XlY8nf1g5Sg6EoyPgEKjeaZj5xxMdDzNfDucHhk
wqV7rhK01BRveCN3m2VfiFLeSMR5/01xVZXS3QV9aXS6ygDorLXBRPEJ8m4gwQdcdak7PBacO6VJ
1AcGDtPO5vtLih8MZDFGaqriyMUhyqoEYe9qijKT0zFqQzLW87tm8jQrpJVGm5geBYNpHePBJSc8
vObB05Skt4XLiHbgWKp7UuSZuunSBY+M7tNx+MY0PGev30Yp63NN0VgXr1VUqC4f3NqF+zHMBADk
WPl77cdMTOGcMouvUQ9miIIaRq7R2L8LKLb2z/u2+xDBQw+MgVoDD/2rn7Ot2eX5QGqOkgAfUmfc
I06Oxkb87hijoVANTBX5csiqlgYECzHhyPZIewczbTZach+Td86awgU2CbiUIyaaZNnOHqz1G0Bo
LD61rA2eo59To2lPSeMRIOrZxENvXj8xM/Z6JdE9HtXnF40Nit5UwgzYSZa8/5DOv5JgBGybjOp9
HCkDbTdNS+RWGYogQMv6RlRFpumOS6VZSN7zcILIT6mbw6weVP1EdeDBfT6V3THiOzJuxEMEf3Ok
6+0qCnZGcy9uQ4cvkUVBmPgjkoodyIeqUj1xrieOa7oQVuCzbfcF2zhP+SkXlut4y2C4uv517q9A
Aaxj5dgWqDygxqEb7jxTpUY4E82K3TSa18Z08wV2Cd9RvwaDVg0p+yjonzL953BwzQ72Tu3peHuc
GVSUtMVRjLEkqvlH9T54lKdLoXv6/MfKyxLG3r33XNC/IKVS0gRz50F2cAkWC7InZTrFHwBD+2XI
wHNAroa9/LuD4a7VXCZ4PcYC7/GSE3FENzyo7VmostwLrTivtEitL4yy8zgXZIVEmR3h7+C9jxGd
53ocwsJYOZztCf/pYYBhQONhEwiwY+ni5Tf/9WK4SPM4Eq0rcwgxwdqH4ul3ZDAEMCQliNe6siYo
GnuO5LL0xGTDOGAb81n5tBsaag0U6NAOLCizbbHAMQbhkFnrz3G51Z++YNVV5mimnN4B0e2EzBth
IowF1EaejQuJ5gYg2HVdUDdhkMBPdUcjFU+6UR61D4AHQ4/RA3IhviO9WOLM4qESDfEf3OYHpTRq
SeRWeyF0WBNEiC1qZXeBCgwYB/alcBHjfEAfsO7uaBXbOwT6HbpuqqBlxjL/sB3Tr9G6MS4NUWA0
JPXDkelFkN8DXzLEjpjp0ovfpKY/08amV20hmGYy9gUeDBC18jKlzdo1KRKNgHBhS9D/555lVR9k
1QNxnc1NqPJD89H2y9GuTBEmNo69HjWP5iClenWDPXI3yioOLlrSYxI7JLOopcj/dXHZWiPrRo25
gfnhss+mDC1v9gGGJSWjLLO7bJOUeOBP0hg0GiIBmiggPKM9mosXWLm7dttylN9I378yCS4ldM1u
DXtlwb5sbYkZjPz1h45gGcQuhooaXOROyvtZfIkRtOsirmGmZ9irNTwdjxZFdccJGAdoni/9dSkS
nVDzNbUeo/9ecW5szeaiHH2/MdUu0euQKrIo1Gd0qc2duotZ3jFlsqhJVW7x9U8yC7rPf9T/V7wO
EmCDoPgF+4Vky+TezOe3danP6fTOYWbSHJvS5oE1kV9WBqgpB+kmfxtXqL8xm1buzM/gtW7Gkz49
oNfq325CERER+l185k2HRoVrDvHGAp9rOwcIlbR0RMpu0KMraoTnaVJCaNHI2f78jNPRBhzechZr
kDBdCulHNEBFnwW7oloaJeZVTKr88PqowFn1ns6nRzxH34hyJMkREnxrRcbyYA6Yq2qDFeF22mVG
IKaeU7CMPMsclViD9IVui6ZR4ODPYJ3yiZkVHClJvztQfnyw+HRqZFSILeC+UonwEfWjj5gU6V9M
VpLirUPnUD0aQboBp4UmAneL+jUq1yWZ95ecEBk9NbFlKFnpdIsGXDcYfMp/6qRZjX1XtSLWporA
SunG2AUHUK7NtO8yu+yUVYx0sj9tqZLwNtLnzRYpd3UPk8fan5AKxyFWUstK0N3IRVTxyHLUzvfi
ygqdDiJ0tnb4faKS06SihtHJwG5DksgeIuh33Utr4hTU2tCR2By7pXTXj7KsUihSjE1nWB+kEvGl
zYQYEuwI433CNzDjeCJ4AvAyqgKZuG28Z3Hu1shXDuICc7iVOwQJr7aD48Cs1iP/tU7DLeOr0Rsr
ela63G2w5cWD8RU2stunVWFRb9rfEOEl0sWhRyQjdufGl70J8XCtlEdFT1Fc+V20QG/nyQpRvtck
HlsxZSZ1zs5UFzU4sZmP1NICIzKLxEomDteg4oGWpZwc1vHRIoH73RBhYdUdJnH4plq43aSM3rZM
8/v9oy7wVDMhp/+cbfXJzTz6r0oWrfbPWswXErkMVaAXF0WJA3FC6QoVWnPgQAH2ddlXEkKlFzqg
Lkg2ddQbQWfC92EVQofdNv0XcUZBGObzPI6XlV6/fln4L/0fwqXJaiS8T0xT3EVkz3MeYdbU9RKy
TZ45G72M/0DNXhUKZ5Qwq11qihblScWLXLADCMSknzrfgfnA+Tec327TytKmezUuEzQH6NwreEhy
ItZE7XEKAgi3GcKgSYUz0tbr3SGo3ZXhmORYe2RbdPr9BmhX47fwNHs0aZZ4Aroe+/+a4hLeEQlM
XxPEhdN2HiMHwIXXhAfoju3wt07Go/QwrWrGd0PHLv+rPw/vRrv6/zlZdNUEGZLyZUw34rXPqYbU
KmvmZzDBd91d0qrv9jMTICQXuEbz8LUjZovDK4/w9y1xnXCPk0HX7T+0w+kb4Z2hpgU/kt2yJn31
pUVRlOnOkzWcrS6MTC2Icnp8zUuOXPBw17x6BvD2unIgmYauJCZ+NGC3d35lIiCXujKDL/jvtdxw
KZOQzLIYOfCczrnDRuqttuhmz48I05GLLayqQOVJ0xZo3Nm/68LT+9FSHmunh9EecP99TVHy7OpM
3U9ERz5bhwsxd49IXaeKoO47UvoQLLr0H85eRsOiIjpMtq2oDZjvLiIX7sS0dObb5LuN7m/k0n6M
LiQBZGE0I5KTFS4tLk+2oWCpm/VEK6THMmOBRG5Wc2jco2BtMjgs5cnUNfTtoflFwsy0AHHzQqnn
PODruVHGV1R5SYiX0M+r5D6DeloVVeKhc0vHU7pLlBaFS0oEHgM3FQJataSoxe2nPOi8IpTiVq1r
o5WW4kdxyM1V646OXlsa2Dbv4fw21EYvGCwBYE2uKYugGsinNpsEvBUgBQ3T36Xvzpbp9WLg23+1
4PL7pIrNryFDvjU3ba9aZvNLU4w63H8Hh7SIEXGLXbu4qdm9AFwescQI7/2AjfcS/E1LFW4MC18j
6MEib7NLQAPz8rbvYsLkTIqDGYdxo+DP3cH46cT4l1ckUS/CrZzOQjdwR0QelKih6vOFMfQqpbSm
mdxZQ64fhQnYFSrEn9LVexIY3tTDuyh5hEcdacfyxNrCWo+nhKBrPsK+TkyJdiEr1WH1woXxdu0J
UUHUCTHqNGx4eUlvj7HeWmiwEJ7xr/Vn8LxqVVyiANHYh5NWWJslGK2qElzd4OCOI0PsjZiKyKR6
+meKxGV1dLXqrbrH6kJjthF5Yf8FtdlpZ9/NxN2YZ4Jmwg2qaBB+UCXNYiM6mJxANg+j/MBAW45C
0AMgntMp+kVnGQZUoEFNFW2YwTPCaRUDIN4hTHdW/ddJr1RFJQipDI6YmFlQ5//4StI/yA2APmlY
LS90hWPpuU8c0nbwti2QCUD2uVJLUHRHtPll9K0VmhhL0qqaVo2m6mjZLgJIjYXlTtJB/MPoYDPX
RU5EgZXr0BQbGpVC4WimhJpOMJjqKxu9s6SQMyam8dlRLuyGt9Jwsl5vAmQoAzAVLUhsS580uHL1
wVuk9PXIeLZY1QtOOWcHI2xCMziuUHc9gV9CEeQIM0C+rQqeG6CrtO+Ah2SYmE4C3tz7Juz/s5P4
YJmY0uX8uyDRDW8HkeZOeZwib06giNI45Pn+WHRqzxYMfRdC1yXrbb3WK4iEOqreNrYGVprOpVlu
qgftifIuUtCTUzKRoVD56wTfOJd+n9ftFP0nQ9zMKAHRtAN4guxFwAa++j4Ltz3IKqVv6BsefHi1
AY8JZ8YZwhinbOZ4SmEl+YFYkUws8EE2JDTn/d90zJkkKsVGxWb19aONejNUlaUm8qBPHwWFIx+7
3RE18OIqTKbI7RQtLfKVoD75FXMaWo/dEZI4QVjQoPFcBWzAYMKJOhLfjUsQs4JGlS6J3JwaCalq
SmWHp+UC9xnhtOtLv8eepxRc+Ugln5tPhOSiijjM0Y6OH5UCgADI9O+nZVzLEcy0yYJpJzux0q34
NscaezLxZVfPzq1xb9vr3/vBHSTRLKBzuJZXi8n+9v/Dg4XbHxkH62fHqW78PlrOQctKANNAeP4I
Z5ERvTG6g8roukqgkuCM1hZMcONKmUS1L+2DidEr0m2yPOQcI2fBY7eqklPKpXcRyxKVkrVzxBis
uCIeJ9hGBI9TDrsfcoBkROBjpQeZt3qB3wAqvDDb4RExCRE6TA0aYAL8c6Yae0vv+LjE7Ju1t7np
d82Qu2Qfc9/s1wRsJuzDdPdnlQnEE++JZS/zvXAOvOV97YMrOUghM1+lm6zxPrQAKK9wTvCm4L4N
Ee65JktaqouhMMYDhAPTofktWezvTWYDxVkjAT7JHkW41zLQ6zDIg3lijeLhLBvymnGharqzbMxd
/7JtNyNk9alMbWvWb5LJR0QOgW7tP+PUHX2nhrLhirzGJCxjJcJL1mup9ZqLKSGqRye/dWHixYAR
v8gK+drVI+8/FxSedQzZgxhtQmEhoo7oQUUD9c+guTQa7Zq1XcmSNZ1uCgfnhktKku2gy5BcKIB5
qPG0d0B1EqrMxxSd1N/IHBuMhfgiJ7hd+OpWhUj4o4UEbv5JIVojM24pQ28QUP1g+J6nOnwloAGz
qFmWmvBywVJ6LyCFYVDypnAoyGti3fOhjwosd65bsrwrRmdfnIt5mtC1K3C17skXsW0oUDFsmoDw
JYn3/hsnA3/m+ybQBaLG3Vm3NXTyDGUh8nDMo0NzqCJAIUa12t1ISPMu8Qi86yvV+c3VWc62TSTR
qvjOzz2ym2tWASJJpwWcLOpMHKZbO7k9o5wOp1otAWkkgZkXJoIdeNjs4kCo1PoevoIRIHrj93hp
vjIgyHbbmv+aoJ3wQBCC+pZkaNeUcxILs+zdKftRzaxkO45/9rliJcNPdORamGUt6v2NYjpjoP4a
qiELT3JC/LhJ+cqNtlfWypVwYew3vVUhbJK1api8N4TPry5sosrwf6J7Q9FvH5iW96fHuD7yxP0F
65uw02PrmIWXwxYx2Pd36cHMFYh7+Msl4NEb04bJKzknISYrQu28Q2r/k5ziQQcsCUSYrNnZkdQJ
8OHBf/xwzn40twadZdtL+UlitzjAfNErX/MvUr+JK4gajqa2R1sONr0gxGN3UY1H8pEuvr6qxyiv
oNze5Y04/SDVuhYcxj2c72MttfokwBREpPoV6QYV2Keg1Ww3g5I72DE6cpEXKTUOmT5pLO8+6bnt
FSL3PsLv3GHagqrzzAIlnb/oxbSE25ncMW5AmjNj7TrCoih02BKKeqMSlRIIeXeOT7SnlXurePBH
zvd1YPj7tupENGosj20ZcEMzYSLKmHV9Cy8bmlvnCNNGEYwu99UtzzX4YccRG6upY7hWIR87TGN3
QhKQLs4qpJJ1G6H1Y9CnWYQq/2qTukJ8WCG1JkYaNhSfWYD4sqGw3YCF5QBgKaz+ns3lzucBbG+J
WTeAOWeCW2muif9EG9Vj/i8cplAQM3RyFSyqQaSEfsiTaAzYuK9jx5ykn1g/AyJDnoKW/Fw1UL8T
lcHFHpKMp75dKmQgegEG/y/70KqHe/oykhyGI4Fj37txuwtrpcG9VGiEjNTP0rSNjJkS5adsQHmq
PUPyMuryDVWVLhUpZm4Sx01Q/dKd5umCrkTTPLSF7zxmS0zSb87pXkyL6WDKIm27QGh8fBi4vTZa
eHCRy1Daq68rIuGtOaZaMnD7JqgkWL/Gnu8IeJS5L4vH22dNqdOvVMNGhXJ0Q+XrA478mKCDCxcg
C140VHajCr5mxWzKMvanko1gM0sVf0ETSOmE1jYN/ugyblh3hLc+uOAEBAEy/uokl4Y39SMbBozJ
efjmvAtG45NYijHrsakZ6fpWzYTWtawC41idJovDlgAKJETKpmHTaj8UHTvze8jYW4EQI9a6Yx1V
J0S5b7bkV5qmWsKWy6lbVneoIm8V0vqjSkeJvJuHtVokNW7iyEYch2D/8Eie2EzfexwCtNHCfGS7
T3+w3Jg/ME4pfGjQI1LK2mnF4b+FQWn8ZoLTU11WU4yrhBVHgbBzWeV3owQffmpVRIE7vzOUeJZE
wy8Tw3EEOeASnR/Gi5VcGUvXu4+b/2OV3t47kNk8WG/YaLtQQkIbDvlbg2PeYTawfPnJmGzKHI8P
FNarNurGThzrFi0W37rqEhQ3xnnyf9+da0rBrpMbDgCZoB3jJtuNbwjVdy8+G0rC0KW+h3iDHwr+
ijMlKcGOLrsI4mH79ECiO0k0rD8E6i2/0toV50sEkAygBe/Id1UZCapWsqnujiTy4VtR6ucb9Lbt
aWIewIg+FrBGCOnLzSQFyLrHf1KdCep/ytg2Pxs7Dro7UZOtgF8XLoIIX8SoCCqLBm8ULWucywKM
TyJa6FA6wCHy7/uCOh63o0Aw6xZ4XPXTvyzT25jmghnIYIdr88Et3M+JKR1kBHUI3+5gQdoXLrBr
nE+ZotVE0Hc++aOlZFWnu/Ep0IulOWvr7ypLwxuv1EA4EZi70JPEfKO0cctDuqeWuEZirIgyNadD
0Q5loAO3D4LIRbXU8Zk/mfm1iqhG+8unMkJkBOiZN3nx8+LgPibZyhx2Kj5tQ4WRkYaxSUhacsgy
vXrcSTnfhwF/ZcyZkC8FQRRrd8v3Vk66bXGV2MvRRbtRugIBF4oZMuoy2Jd+5ppHoixwBI+ACuf0
1Hb9dA0A93nSsGHEY6gZ09fOcPFZsBSWixyZmrYOh75m9nHC8AMHz18zSN9SAFQth6gzpZgQrp2C
nl8WYD1RmI8rELDuXwAWtFQRQNyAcRzdz++JBbPesUkRGS/9n/Giq9r2D3oNAHJ+6eSm7ckYsylT
ch8oYdVkF/BUs9OKwygFzIBwZfIyyZi5+x465SbTFsf46uTTjOpXQyciNYEf1zSsKgJ+0xGmBQ/x
Rg+XsMysbmIp9Nh4Fmja0DOkM0eItsWTjHw2Sd+7c4rdm6vQ5LXovNmU5C+Jm15riSUlnRCsrJPs
7x4NZSTCl64SNvseox9RJp7GurAJjj8xtAOyxdnXEckKUaXuMKpHCDFZmYNXAjeIJsphYkjVxW+S
rwhgOv47dMnoPQDqqb9GKdck71HiTccSQ0yjQxFjFvZh7/4Ykf+UicK9xB+gDXYbVkljwEpnjKf2
b3dEKefEmr2e+SiBbEfGDCE2NMqRNZOVA4ZrOs1dnK6LwggvQTNJYi+ILVcA1DMzv5f1MSxEFlN3
PPLw+roccIE4awFu3LIJTzOkC1YVQzfbinHZXYmyYX0dFoxzD6EldC5U/v+EcLoXBdBCw3IAgeD6
sdo0nnB8agSx3JyQIAo8B32r4MFu7G1gSzt6MqE7I3SO1aPPOiN+dDZweIWiEcVdCDiJNEWKhw7i
dKuxmsLscHe+5KzNAKs15DUdro6Q1nR4iLU2VBBr1ZeMlkDtLdm6c2rKAk37IC9IVaibM7qpl95G
kSFVhDcNYJ1brXwVhShqNOIWTfiEvGyKV2QKqAr9K2mkV4pKsBJBR4kfreR+izIqf/fT34LmlEUO
d/UxXtfrKwjiegfaq+PMpyIDqzMUUG5WTSr2maBepuP35NUWmkZxHbt+pXXh1x+btfcUpXbjHTt7
bPKBA9qpLjKXzLR0AAr3bGMu6WPr6K5I0mpsHEYrgzJmFW5ewT60yMQ4S2l7UDOmDCLvehH0r/OR
vNG6YXHCbGM9nFPyLVF7u1wht0yol1xMKPYUDzeCcbaedIqVaYIYxfS/wC0tko+PzhJv2zMy/yjM
8K7gHlat3jJr8JDqDz1AyZci51aaosT/GpmOnbLPvck7JUOXLKNbRwr9RQBhh/i5I9rLBN0fj8y1
8SQA+/XM4UDXRMnaepLjlRQu6j8CKkMaVrTSuTR1xrlJigoe4MXjXiT3rNhEgYbcsEKJLIw61MqO
Pl2StjTQ1SEMlhi4UYm6M/D2wDzgvpVEpuERHm4vyXpcflodGwYzczKdji5zskTYEHapdUXn3xiV
/9+bGw40OH8oJpUIwZ11+wsFAu/FJBKVNVZ+6fgT940kLBZm3/YnBrVs/Iq7iD1RblQj6fHlcWg1
UyH/LYlxS9SrpKRaOg6Fg2/Sa02ZOEi6ev6dDjHjchgIkeXkb8s+9wsShWEfmjixdyByNp81OfSA
0IWIARxvmcFY39dGwp6AXRr89VY0QdwgCv90DvroC8nx7fpb+K8OMxiR3v1sMUB7fSrf+x9vl/3K
YtolspVRGJB54bUeRNOqYtfuOYCBQ3E46E7cTBgnJpma2B74+wnuhn8tV836GyAmUPeCXtMXXrHf
SIFFYEXyrf63I8hp3/lh1OhsEY16uT6ZMFphlef5/OJQVF8+0jhpIs9ylN2bjOAWdPlcWNckv+0o
S9JidDdv3ory5Z8Hjtqw6RNDyz5Xtu0RMQVkCaK0TzkuPy4gJZaO4oWpRKyTzMUU9K6M2dfwxdwx
yKM+yVyQPjC4mbwQ0DJrraHFaJzqT6dMskn3IdYnXsd5IfruyjVJFszXBNp5OUMcxrStmobKBAyB
iQ9UIdLdg5o7ZAe/SzrAU8S4xq88u1ozoEJrVG30ruLG2ndbvxD4PphRpUnTg1RMac/dRJ8pfQQc
DP5aBwpRAy/LVeJx8wmCApZyUVlZ7b5bVz5yIxIH6bEU2wBZEr9NOWYzDcMNQucf4tXe0h4bYkXn
SYlser2qzghyW6ILVxA55IUOpksUMqCvC4hCqledL4DZJA0RlEldOKQgv0SoFVaYKYy3zcKdiett
/XtwAY7uHFU+bab/cC/yr71yrfopY6CvaFiazA4biaQ32SBP+NV+w/u1Iwl8lAHEjk1AzRRFK/Jq
YcWjQ+vYEpe5aPtJWJdwJDQ7dlAUAzlCAYNSGu8GzuYb0BZ6JVHv0j79HtAv8VYnBtEmkrgPuWXS
+AjUJFPUuk1YzeFELrlCIRPLAdtwpXNHTU+pNmwO7h4u7HR4kiLISW0bD5vft7Sfa2KFri8b/VJe
/V6quewK58lyK5ZbfYRo+StAsCsg4+7u5BWzCCr3EO2BKGNXq+0djQHdFCDfFv1nZgjKpeKXRfe+
zw4V2ckpfrYBCOTe+5Sgs77YdMekFBclVT7AiFuMr4FlI5UzIIchxDALkc9zGoNgaLsRqcOl7rbm
vnzMIOEJoXte15zo7CsilsjuohfUV92zVkfNb0U4SLNqJlYsak6WN9v2oUY0tSkjj1D1LeB1q4mj
htCNKnuOv9jY8DQVLq6c6Cra/h8eR3GYHmvapeH3doXcJqWnDRsumo2sFi6znO6l2VwWeA4xwE2n
crQUxXcO3d38yRrahNWEchw50dBYEQ1QqRhF5bgbS3Jfq3EWGb+Hy22Z68oN0/lY4Rz4V1ECxGuH
3WiLFkfGHNRXUpb0bGh/551iSxPOEpUIn29wJ8gYwNvq7jcoQxHTc1l4pLZsiqC9nG9gHq1qVe8x
Izmt1pL6K+kpi8ScHzIVNGneOZF/L8RwX2KjbvvIOrYuE2hUuO7etMZYwRIvjPbIFP10nvN539i8
jUAfU3xFKUg5Rza04M7No1b3j7Kc5JUAvrDmy5UT8P9zizo7wt1fCERkaC3rdrbwomyBCwAADy06
pSx0M19RHW5za8/5u4ef7FTxRMEMuyEOh9GBe02q4n3E4wKauCzujtAiZdrSNpTr3denr1CbfJwI
9E7BnlaKQUovRpzOIneHAYeB67jjBk2KUjnXxrnOizFdEYdiAzDOshEtcL8LTKY05kUZ/RJo+K74
45hYH0D2Kjh1piYMIChT4WJ3DjnN+Hqz+ryfkE3Tkb3ICLRLXGN6kNSE0cconfjG019KQ4wrtp+0
CJemuFdiswvq8w28En1MVlyx/2ipjZKo1lwWkAunSwr9hX9ME/bEhDE27Yrp02zLMKCWPdufoN2/
E31DcQM6GoPgE/SPqAyaPauBxIU8/sDyhRPhAB/y+UgDz3rNsR0PSeL87g8oA8xqZd0do0LVRi25
EqK4sznNwAMljhj/IP0LurjMKn2/VuxXjnzmMVHQwFb6IK6eppYcz2mvRam+0RWwPr+FFF7CCtPV
Q6gvJUpt4iNeJNGaT5C7rCx9IqRuXtu4zG3Tttr30Fd7pK09ZxJuVDs6I/Von3kquP2fjeysnalG
gZEleYJcnJe7DitWLvqZW2LgLX5wPc6MG0hGT6WtSNHubFMTWmRDzDYn6JeRhs+SyMGS2SHmhVe5
ohDAFT6S9/QqvbKwzflClh69gVgmaJT8VCbBRizL6d2lCr+lEqm+njQTuQSeJPAsv2fuF+zMF3VF
uzyZ8JP1r4lel+2ytueklTLzYAINHu5PKI7QXqhA1sPMOGazAaKFQ9OydWvqymFZ4YC9P4X1Qr5g
eweuyBWBK8mVS1CNUmu4nj14egNecifYzySn3W76bMKVy2XcjqODUPTWfyZCZYC8qXZ4POfU5baZ
HMKcbGfgZwSbCXilBd/dVOZgycqee72NMRAk+GkjJh7wYnXGBdtHIWULNGuZUrDxOdUwKTkRj5z7
wl45P4f1LmObdabZzGE3ut505EKoG6P6VylW6Y8Th1Yq98Ejl9RpfHQJzZaEXHNu7Qu+WObXcOFo
eA0ZlSaUe52GwStSaWjDSEFHenw3rywQBqCeoeB8EOTir7MWC7uepcS5Da+3F8R6hSVxZ5AV4Sc0
dIC51LrsUQEM7doyYv54J7x7LdVsSghjfq3bxho3PHpgfKm5BITpJpSpylu2JpldLKeF0RZ9XXpb
3iCbvlegh8wxxdqLHeFmXG5dDjhIPHi0F6DJ7F9gLbspICO7t6nQaypbB+xHxF9vXxwlV090XSZC
vc6BsmqBMAEzPKquKC7I/JsJL6O6Mij2OOTjwkhcOC1z8H+Mz1luRsPgVVkFvKRs1NWyDm750ZOZ
dmpHzcgzQ+W7uZZJLRN1xOEzxEVz40JQkLNA/R979zLKPzbae0CVFTdBgBwAlaA6tepM6V7BwI/b
AqhKTNmXL3a8YV/dL6ttZb7M1gc4MLAI0tSWLMnrDbyIMVzqKl8Qr9efYmgx75RkKalGx7qF7DGw
omRDUuDcSg1Wn28ygBnb+wqJPyc/IsK9HLHoun1/14PDzQnVlf/JonohyAolfGPim7dPuaFdhHV9
wacrys9l0ND1n3QQm7iqU0npuWNKfJpgTgG+8NeULV5Mij47k7BT/tbejqr/cNK9umy3uvOo5iIe
erQw8dETfKCBRZ48vwgMDZL6akz+mO4aBW/XSjc7xMEqKVez2Ym0dGYlEcf6vCg5nuEkPo63x3c0
78RtfPDm2qu6pzIZZOdVMMbcFWQTxbXvcfd0CnrkyGq1q4o6sSw7ukozFG1t01isOmbn8GUMKXcS
0X9mp2x63ppOHb1FMhi1+Yny1ZJW8C1w0TNz5ThD96PSlcyo6OkgdFBqL8RCeCknXgZ+OeonYnLn
7PfHj1+DlvIztgic7zwAD2g4/GjnsyMtqhi09hbGovmk/0KvV0GO+/TF+d+FFvYnU1Jbn86a5/Ml
9mdVSRRqzkNsRcLCOUNOBCDf1noMFyh+Pe5KVnEHjiy3FzOowIOtjv0SiKi+foHBLBcmSIRaoA4p
7ayJ4AcsUeJRBZPhLvlCTnV30peChJDDkUhBVGrmhme/vdnXXN0+gaglKtcRlvm3nM/MQ6Lya8eC
ig7p3hxUETCJiBlGjiTRjs93AR4csyIrTZcem/cfXAFd8cwkpNqU1gdgOwcjNuHAYMVLR0z2kvuv
xgdefG3kYcVIa2BbYQ/ZeaIE7/vwcCPsFIxTz0AT12glOOYc7ruQXQVGN6GaCZKJd9PfMBi2Mb09
sHN6CUYp9rdmRtHjz9hhYjhAKxAVzo5Nbno/Ke4UGj8vhaqop+Kjsa9x/V8SVJpJ2KnK2kJSYYwG
/23rLUvLL+H3fMCVAYzFJsVJlLKgtMzoy/t66Dv4UZeSWa1u1Z5ALm6tJaridN713ikAJdCTrYv2
uslJ1ljpv/RKrs6iq4iJpSHTfCKwL+ObzGR9mqb4fB67Ho01ZxprYWBYDczNJLqsE2uH7/BrkeIv
ozr7xkWkFvk7jDPpvBVNYjt4ZptkGmq2WMgfEOvPBxIzEMtO4+gYiz9Cxj4Ht5fuPPNL9nPWroPd
YskIGAgDio3hwUJK8c9kYz1FQHMZ0Tz55Ai1wDVVnX+D+4Bfx45eFo618l3bZreSDV/jItq+uUJj
DN000ly+Qqp31o7p0UGr7bsjc5vYVzAfswxj4X5mPpwyt/iyP/iyggZOgwGOj2gsBe8ZQ8rMZgLc
RjokBpynuFggWZqFU5OilJcMc+t0Ia4nwMRMiaJcEgbAK59i2IUW6MkWs+N40m9PryfkZ/mcftlj
oemHJsyWejHiBwwFecZ5CGIK9hhkdXtJsGdQ/8YtPqkTWGqHfqojmdiIcN5iuAznwKZv+fe28yzQ
+EH2FKu6xqC+YARR4DStY9zc0a3YmbOEFIrevuDEmdTIKkQPy7sYtAFTebsNreG5dFoXbTaS3SNX
qOvMwsamruura6dweisJwm5rKCjkjt9IFb79ZGH35ITycrON19Nm3ZlZLadyTRS5DOtMETGMmH8/
Ryl3VSlcOuNU1c1wa+4MGsVIBK2ZKTHiUGSi2CBE1Y820ACkAlB3q34n1sYn1LsUyBp81A4BMS2A
mZyxfe3zNv4G0mGciOUjuf4dKxSewy1eqF0wOKyocdd90vFzvl73Kx71NaZ6437hZWcFB3hbxS0M
7NbEKX7FnmGSBo7Xbf/qkyGu+3v18vrOWsdX5vipcXZ0ygRyV1jkE0+bepQaNJUwg3I/xiTVkI5Y
ypP1noVYG53jHqeFbXahz9nXHpkVvkhMZ4LHdcl7FFKp/eSxXV1AoOD/64ppeekHfvsEPJ1gDi1U
pf9BQmoJoz2jAi28ObuvQIgWNHLr8nHUjB6VTDyY+EFyFc+g8LE8VxMDK95J6jmSxAWlENmsLPCM
NL8DEz39dasToL1vCSUsgICVpQfL0HXyyeKSHpF1amNirrzyBqLV92sOHVl/KemSNzkjwCsNS/oD
FeM4h2aoNUr2qWSdXC/+RmPnkL+LAp+6FiFrhRnWouglqFFsGBArOqCbjgv09bBSdXcvgBKudzc4
+O1Sqk/BjGQsFx/s/ELxRJuT8CmA3AV3FNurU3uMWVGW3fYCZTxg8pe3UGDvm8fwLqhfttuD5btG
aC8QP1SzweS1XezOeXgEO6qqVso+nIyB4wsckvqQLGj6/ZhZ3Cpwxh11qKUsqeceXBwyOyLFZNB9
SFPOedtP6AXiV+cUJZZMicOFVyK2CcBZFinAJ345/gCn0vmjqp/EHtmONjjWb7RGOCB5UdepHA0p
tEOronGhZ84mZJoMenYrh3f+20qeBrSL4VzHuOWk1ttRvqHnRC5PG1S2e1YnlJ9vO6h8zCPuy/lf
zTdLoDHg33e9xUui4Lx2Bau/2YSb49uN3CU/XDBm6TTJ8+kWsl+tI0P9NUDB559G4oYlL6/1N+oq
TYcJey2RW7WUniNv661jlpE67ZPlRc5SGPQX81H24wxhT5YzvjYofUDPjHhSvAPkGunJ5NP13aPN
yVlEfxHB2Qi2E0A4nBHXCU+NZlrAudX9xriM4lNvDEkAUpVZ1D7LhjKWeOsJiVOenDjA20nTB78N
pBOG7Cz36lpuQ8v4TlNyJBf/r1kIdkeOBx76wUxv4KGRl39c1lgR1trbNf/JJpgoVhfeA0p4y6E9
47T39dBGeMDnO8GOvxvDfkhQw+W4zOmzMnL0cZjlP9dwqzU2vLdOr/q4uTGbDECLK8P3OCF/8EOC
bFDVbEDs2LJMIjBu4VOMaM5ykfdbPpfiPV0V/sBvA7s9kcpcbb34jdYzn0+4U2TwXUTTMOuyF3sj
CiJFZTak63dXcwVEgGtNHrb7TOBUWaFZPpa13d2BTafuXkNY5kv0yFlCBW51qPrQYsvkyaw7db4m
p+Js+CjPVQlFVDM5f4KETKHI2dtejc952/Arm0o/2+o9nI2uMHk80TvF3nDWTGA3zwpYzHbryBse
+eT8AeFkou7IjDcmMUT5ZfpEQSBj/v83mXoEHmju/xoD/6JLOJIae/0421l/jzh5mbgHNa6nbbQr
A6NLS0gQU7/8JfJF4wSsdUM8yNRu7hG8rNnsn6xE1EQJmwjgvqyNOnmBDBLauAXOX3Sk8n1T4g9w
LasEFCWZrsLEvlws3pWrlo5BY5O6DR5WMZpP75TDTwXR0fBkCyGpY3anjxIZ7vX+M04F7QuG7gJw
YGqDLe5bbL8Lz87RqxTZDpv1sHYgVo6fJQ6bcTv8NVv2fLpYA8wHq5YSoV9q65J69PUMkVlnkM7Z
+4IR7bjFJa9ULu1Sze88UNOGlkMFqGXXw07vITVsFhds7cBIf+7t0nY16FWEjioDSBsPyp/TDq+u
PHAL7ovEYp7XQqI4LxRDIdFfl3fEPxA/Lh0zTRNt1BFRA/+YG1pwjUF7hDPtwgPfTtQ3TQHOmdIM
XCqWCaXv2ZxXhyPswr2KkZdiwg/4w6TW4kHb5osSlbDPWmjJvR4bHZogP5q6Kqt04eoKhQqUixSD
f9hEifZO6UYnDjkPPRltDOQgVNcRjoitWz2qxLKmbUwEn03PfyfHjI+yHWvFkbeku8eZv4zbXxyn
2i8VcODt9S7mlVbI0tpFAVDUqvAWQmT6pruUEbJ/JucIj785J62Sr4S+dcvUA5yoVG17wnovf5J/
3337AXqsU4VE728nJt92CMV/KGuxi0Xi3S2qU4w2FSYaatvbGNAlksn7XTZasWi3gCP5KajiYl4d
2p70lZ2qolxJ5t1HZRG7hsZCl6uywe2kSGGqW1vY5tnNYPHYiQ5Kpn2j7UJZf3j6bI9KKUxXaVgH
KyvaY5AJczUGnYYA2YfoGQUvCY7wCBqX85/qMnirORgOub+qL3wB7crkPUoIB7k9rpZc4Aa7L8T/
6/P6wnyXN/EoCCqmZ71RvhRXp6KIdv5vml0EksVTsK7sKgOhKgZjg5ntMyG8VC/JZh2zurqHO4qf
uhIIZ5uPXBz5tSHqNLVlEcYS7AczeYZLpyOrQk4N0Vcc/QEtHzE8dCB+ZUCGQxk+wgYPq42vCFHO
dUAnFeH5wMtg8r63XsRc1qkM5dDu1yfeTqdb8qm66cgNXaOxJfOTZZfTMG3RsjTR0Sz5Mj3z9V+p
ocnt4axMTDoV47MeEfJ+dQl4KUPQ4gMicnV8JYrz8Qdstr60dn1wUuogfCtwBYMQ5QrMCDlMKZ/x
JIPpkRWbLgGGpyAOcqL0tpoI/BFhTvSFQdVdIc4kMSlxlAoKNq7PXYJUYQpr/seTTWEM3O9ijczM
25ROyVn2+MC3UvnKmTeZZiXfsEdhwpYSYcn7DuE2AEMzy2iScQiAxOOFT6zqXmsjSOlQ/cX0DVCO
hpTQeBxz7ZA8tQebQv2JBjrhzg05wJq3tau+yKHC4jtE+jIA1ZW+KbD4VT4s/XECEPkM4DhQsLZs
Y2D3uW7S+CeDMP/R6qnhAGSi2hhSy3Q9caAJSz2Q/N51DS3kun6kzbFHoSdcSTBKJUdHIpFGgfp8
W/oEBZbEdseOogv9YEezS5/RDzcWstuuqcdQOvmN1IeAyMJMvTy+WbvTyU0kqcchEYoKRedUWxTQ
dVS4C0n9eBZg42CLsNdgo7H8C8s3s8C4Cu0ee/m2saifnLTG3c9iilzZYOEVf1qEnG755M+AwNah
/mjPlgnd583WsZ8LhPqL+/ay4PEvgFvqYxncsfYBK4q/dHUyv+bt32BP9jY2hcum4bVVYxdClHKX
69m3StyiE3TZPWpOH6PFhY9ux6dkS3qk7P9GrXP7HQo3IZaUyCMHfP/N64D+eMfnqG+0wHK4tzh4
5tHkCCIWDGGHTIi89lrp7EWAU6a8OvetKu9WBxQk5XNWN3oMPnBYDB/YbC/M6VsNtJUJmPpql/Fy
eyiE4jNVcH9GuEEXFZpdnJG6UTJWF3aRP3YtkwK74scb/anTliJWvyLD1TYxZ+3cUrX/bdHpoNNA
45VhmnBEpS/KLk1xc+cfUpznlu/2Yex5VUErwiuJJXIaslrym6b7Y0CDcZnvpAoTVNAJp0hRe9nY
ec7VAdIJy42Ww6a89jA/ZVxFTLZAlMyOGCVIjcQPnLiai7Yuy7oWeLcPpAK4bU3e/+niZ66qKMUW
YrpgHr9wVNVjsaxPMiHpTRYqNHbH2x6HvX/GInG1TGBjEZFpgYQCkLruodnD471ySx5FHPR1ihHd
UEk16f+bLHKUnQCh/k9S0+0C8sp2LfZb/a/OO2wgjq2hSQ3C8fwjZQFEx3DvxPaUracdLbvNHM/m
A7N5jtr8ieCB70o3tt1oL1xhsQ+k6aS4+S8U69P22OX/IlNf6jZzsBEIdd9LkdLIVWnmPZ+QdXix
XBWvKQKnLoKdoUzf4+WW+Dv1jJ2VEUExKn288eUmXklM6nJHmvvJrzS3ZyUkdGjiuO8DtwwVaIpw
OY0viXNhPpXjrm6PPgBwbZY+orLPD2UFnl7XVxfyLBxrfPkBU7XxbInPUKMiAIguUHF9MFTA7Cra
AB1TIYFjVzulW0vTho1+EWuSwP8s7oJY+Vlzh6Z6AUtCJ8SoKvE5eCkg5lQfPuFwwwbknZQWs2eI
aMF8Q3YgTeu59rxnPDp3q8Z59aIsTYpZq8I/58oa1Qjx0lv/JTjbXws/Hs8tNK0xS76N+z6Pav7F
6WiS/rXj3w0hXjrVhDe1nQ3MDIPTJOkZqXBce+cRf1TcbhjoRFR4g/kV1MqVFgrMkueQ8B6l77m6
RDGiQiBN51KLV2li5AHLm/7njERFuJ/2N7HJCvXciQqp38o83/feKRDmtm00hihNZx+hohPs60oz
GAvwOBIP+E9hXfU4vuD84O+NqrisdwM7SnFGNIqCOz8qQSxiiCeRuFTYewu4dsqyLEQPPTWtXVV7
9nOyhLIZFgQ+KbSIE2ZlvZ/f+QDDQvAaAUWU2KjAljHlgjSfwqTWtRWejyJdyYdbS6E0r2Dk9Ack
iUiI+hrY5HpCMyF9QHt1rKEaM6EXLunKL2m0TFQzPG+J8jsobraOcsVB5T2lPf9XvSlWDDTFnUE9
pirFJPfTRdrGZOe9xVVD/CxKoHrR45I8ScxvD2gFjBxyGT0SWlg2y+4uDooccnaChIQb/dFCsaIG
PM6yjv/nH/FUjazlza1OkqBEh2Kmm//HmzP83JHfxcZykelxFxe7TgPKM8iNtFfuPYoFAh9F+Wuw
tnZkln/PPM/t2ujI5Oaq2TYid7j1MUMvSS+hPC1jgwEi4ytk2cWo8EsGMBua82xwPCcc/R1vyaxr
YVXsStpdgj3HUv9Nq/tKJwNCtKp1tLbK20fT/F5ZmuuYVITcBE7RXHlvEKrA6f2j0UIdSIbkTRwY
tNBsBbr6QNACmQKS0KIBzsrtKTJ/qwA7OwJd3GEkjnREDZ1tIj3x+vw4iCyaCkBXmtcVGgThuAs3
0z75A+P1oHlV5MZD1T3XiTH+Qcm1aPiu1D9q7NUjj99NTX2LCt6U6JYyUQGh7kpUwMLIelUK5TUM
5sX9Y+RxWTbeztFsycZNaHD1yS8S4J9AOePgKNwJj1X87l1HrlcDmAw49U2yGfcxR22g4W/LRiqj
uE+jiSyKhwO7S/aAAET2QiMsDSF3X4w66BVmxaCP00mx4vzbSK6cyowOaJ8vB1tgY3sTxLREnjJm
F9kO2JFhQsceO9yC17+0gJK3kthM4sFTcB8Fl9DBnKK9cYD+zBR+1Uh35VbxG7Qld+NkVPH6WvvP
car0/4gIanhl+Rn2GAwcXBH4c5s/h08wHUmd8Tt6pzUGL+WFD0ZtZLc3fv5nnsDmF8ERqCnCaGwE
YsqaJ7Vh1uvwzkZ/MB7k5xJ51AkL4spmtwX8AyVZhxc9hyOCYi0r9WUXp7Y7rXmujA1HEBc2iS6K
H2g0PmdYSbROeppNKBMxsw2dzWu8a6HpRhmnBE2IflpVHf2IQWmOuU5zQS9NIbQwEdaVKjMiZYT4
4GSSgQlDhKoJfXV6TjoQkaQRxIesbTV4HfL1DjSD1n8wtoiiqxjHLu0o0miDue0MvAsVRcVcbO10
sYyZ7Dfyjfg4yffF+yU8BKsrRLpmfoLpLgojviPE/FytQl298vYI95nh6sKkgeNLkTAi13aB2hHQ
tgGt6xHDh9VVPD0ANNnCJLqFe70FnTt3ixVXyfbi1gfGSo5o/cxJ0r5oVd5BqF399nduMaQk51FO
+HN43Q3m+mJt72K5sIQPbAjrBT6710UCGXLMy8eQIiBSz/1XcLFK3I/i62mBkMWgLVWUyO7LzMhx
Wiy1J1trOvdC4wV0O335+5DfkPdBHhbZnSrF6aDEMo4/kAAZr1FscHWcwW+JMDyoCxFNx0yeI39a
Nkwq95i24UAwEZATI08+ND8AEEowc0RvJK2GY7JuTCb7JBB/2wLny4MRB8Y3f0qpG29qjUgngiD7
vFRoeD2RXT57KG/JPO3lAW5zZCtt37oaXP3ItI9DT8IKmvqZSOkO2g7ZUGg7V1S4sNr9u/Dm/uUz
V+lTe3+nGZUwvWVeaZFdAm4+PPuEIWWXxWeeSrrlth0Q3K7RbhAjCUL7x4YB8T5M1xF6b0882GG6
HleDZL/XrhC+ltU9jQ6C/Zil0izYo70OLDjlEbjorK5ZwdYQU0QO0Y+g+huTiOGglcvJ6nxGIFS7
HtF7cqYQephWB95ZawzUP3TWfcXxdowhlHg0nmXIOVenq9kaqa3w2H/9UMICMH7kMRS2NBDcJROV
gdXbFNn8QWgHG/LXcYXxIa1NqaqLPCrLxEE7esijbATJPcp0nCsWKdmJDLI4S7EVTbBYMwgkjdUr
VriGINv2TPlQj0Eh40nzV/URGs40PT6ZQCZTTgbVxav3cCv0NGWQ0ZW5wLlNYLJ4OjSBjPS+3dzE
Z+LpoVxK8XyQnYpGQJ41hHxJKiHIY+AmkRLmRHq+RjYVG6A8wmXVTZivjS4HGwEh8CpRXRqBV4DC
cWfUXoS52ap1WBqPxfj/Pnbh5GQjW2cK8ZU4RM5dy8thIUDpme9WMQmWQZ2tiJDyQ4cvrZKtizPH
l2HMr+e7/FUSgHdXfv3RZR/omrHO/HXxt4ujEa2RtNLZWxAyjeBLxOfIcjtbYhGgMn9V2z0O4O3z
aY1h91y8pkigZJEI5kFnldrkTELDQ7gPUdILLo7V0ZorP0qrjRKWX0MMd/8S6RjydGjz7G/POA6b
5v8B/Ox88/+4XFv6lZC/uZhAgbnzzSOeSGyU0wHgrE0R+yxQ+Sx57hnKE9j3VCl8VdUh1F/MZtRW
PDiI+fwrqLAbrPnlrDZCXFBwQUlIE0UwDfMgRsvE6L4X/zMQJwS4mD06gnPBb6QEtzJHx2Ehfs5U
V9KNuL9hfX5tSbMoNyZP5uJpm+F7xqfVeouK/6YEfAKn2TMXvyyheY+/v7vZFth1NCLUwMVIrruL
z9jDSVOPidXkZ80bYh0PO/TRyuox2+z7+xuibNBaZ9rGzAUC0WR7NiDCyUCut9OzoiwZY34ZIqka
xt6MahesjE5wI3/j9vLEjNm0qUogJyoP8Qo0jujcxwt+cOnqUU9tPOxXW3NeMCeuxmVO/gWKW8IB
rh87/rJCIVxhPeOS1SkBwxRzg6OUyDqX1mjDhl/TrUZqdz0MhslS1EZP9qta+m1wYV9reA7075vt
mpGksoZ5IOdF0sndQn14upVMrpatuDeyk7R6Tdf7Z4rfNhbdaaaZmN+zZhItHo3bA5X0a74K8DMu
PrBW89DSww9Ck9G4NT/9opYePH4EIWkhxf5mD3HnTgymTub+VrpL6XJCTnXwGpnPE3Rkp7fNvfgM
8/hG8xHgAIDTTKDOmHfVXgNelc8BeshwLacm798A9VbWjMKG7J1aYZAIk/wJJ1PEZhhSe01axGfo
14Rh8cd7dIJQvWj074QLTA3rMSpq1UHOvIQhaKo5yBDn/XlH+2jQfqrT/1CT+igFFJXGbs/K/QNJ
79oGt5wNbInSjpXmTVoQW8JVIfzfF8td2oykP4kg3iIzA5aITs1NBtKBTIm3NgC/mm8cQBCaGyfz
eX8DRIC2KNDCRmLqG+xWWKwzYQ9oivPpsrga5uxg8uGle8pgMgJs9Rb/pGfECm6iwnC7tfOf3TmQ
DT3fK/0ZvD6O8qHgqbLdr+jaFWaHt2lrkvUu6w4rR9LdujTJh0Yf3x07CAfCq0jGZyyHyEz6A65e
Dq6KW8ccpEF4SGMFil6YR4R4nljm4FROVB/QsWsH+DF9+7mBhGUZa4vzHXFQAk5/MZ7hbdxFzRLU
4VP6u2VsdzCm6ErFNVaxWZIlmjYVoNoZOYGo0qWLUtOOSIywRC5hA9Q80rUCdvHJnwtevRBgTzfH
3SEYPLCgaJAlSFr/1z/hq18FBhRD26v2XeSENkHf+xVRrLt96lQAjFIsktAX0b2IXidJ+vVgYwf1
el05Gz8bNWtRtQmrs5v8egfP989Z9CwmncpVRkNqyyy6eN5qOXjlNRNUA9XI4LNtlx/09ZSdaDtg
DVMw7yJy+ReGOZl4bQcuGCqhaQRo1BYHuaackuE0UQMqmpF6P7hugJb5+Ffdx6SICVNlo2l3jhN8
xmhgmN/9Aq1M5OCKipBRE7L9/Bgf/t+HMUiFRlVxlWyfKyU59sPM1HoSrow7ahX3hNepzYSD4izq
9wRqxL+PykaORv4ZasqJXm4ZXUeZiYQzlMNRH6H1RtRgez4PhzpEO7H7WGkr6klFrQjBR6G9n91I
FErAsb1TGqZl9l/1QSOogda1erKeoZd4crvrLDKCT5b88wpcwjPy3Yv7gArQ8oichEUdiRnvBbAs
v0FiKmzm5CZi/Az8Z/FK1exSzSyBxV752a5CSffENhRdSTVnoqCLCsxRk5m/tXgid3Wl0pTgenGT
Y8+xAtC8b5a93k4Q4lka5Bvi+ogECVoYYpOW1uvtDJUmDLik5zFgVItZbeRwarQ6IvOkjAssEfwA
XUjq4oLJRTeVZg6PQLBX4VROI3SQ88iQdStQEArYXl/PlFFvT+9a8q1yoKHM6v1nRgPgauy+x0ub
AmZpE+0AGXdQ4CTroVZgxzIFfFFkXVrpIuic8zvZ0Pxpi5X2yj4KHUxBUDU3CyhphztctBMzJDhW
YondpQe1pQOrAB0cECyDdb2JznghAFfZE5mheJL6nek/3s4SLjCoQyn02QmifAlMJTKM/D0rLGMv
l9Q3/Ys6iF/xhzdcE/fI897/XDkv0p9jKRtwdDsrbyFP87BFNGhmBSkTzENmvXgQRqdkpapXgWCj
IPcHF+DY0QBPMpMYXGjAazHQrVbmAnje8dP0W92rpnnvi3z8uQ/39aE4FFXQHf5uGbFNj31CUXQN
hRV41a86EezHYqPhWtqgw0icANG2fJBYelH0vIj0r+JtO9MNUmJt4AbjaC01gnX51EynO1oTTZoN
0c4ViWrcUMMgAXu8r8ihDxSCjTHgD7+MWzsLikXAu9hp7oxT13cMDvzcX4FOHczutSOCFZpZYrsT
GYBo2FFLQuNHm2/YVyCSuhYaYcBs4/xZdsN8KvNGbF334Ln80XQS/6YNcdk/yV6K5vc6RM9K4Eo5
PeT7cL5+lyKT49HYc5anYmxZTbvQnxX96gum3kO9AA6CDFzLSThui5tc5R9q4huPuqHM2dqFji7o
Pe8Yy9TJmHRuKKozZVYlcjIOK3GfaYiaao+/4qKee2od3K4U3kSi0B92ikyA9apNHzfXfDaqL/BK
KENGkd7f/DglNoWKWnOC5V0vSGMJuskCcRpVe/g+70+cvcQD4j/dA6w8yIKISGYN3lZsLb0gdP0p
l/qjHOj5PyYX6AhFVmO2czyrwiZu/iWGrUibvLyF/kr7E+yNeJ/vTC7KR7aiCdivfeyUEaeIEjON
NUpAOk7J0h6mQs8bk7lsLul8dY7BVVFkV455gDIe10PAFp1N7AjHEJqHFO3/f40ivIUnq+ibhEVY
U15s5rCboWt5ZXWf+sT0wsGrKfBCtW8CQWSmED44l7Eh0sE38uGpXA32/FVw1nw6wOwjjWOvutDj
FLiohe2mT054XfRnPo79SKhWbKv3YIffObCZOjOwViDIV+gywe8hs5BloeTeQVXVWXry6waqZv8B
1y3ZbPwr1h54Ajw5ad1kcScp9dY4F8V2ADxLJ5d2cw98TxVscPiS5nmqxmjgel16D/RdgTSv5Ces
aDMNodHbaJJQQJCFT2TZ5/crGEwWecfxEbURcZqVcOYiFyGVq7fltYPiDBUq16TZG1Y5BWPr7GtO
m0fojvL4zJ6perh0kStwF/fBMlL1t4JSLH4ziZQdAYh+BC+ylyHf9jcAhGN8ZUdXPa2xDDDn+0E+
mG6a1cdr/rPdIozjkIOiN5OFzD8frFIFpAuoLezacNu9/runuWLXApqMo8kw8iZl7IPgX5KQhVo/
LUt7uUuRgRXsBk13pe7HseXZ9LktBywNqPKY+aXdX6UH+JaN8Gm1G46SAVFQjfAez/nNvKhOPivC
zUFoSUczptcdUgnNM+GySmuGsjW1PBRJ5tp7L7MXIZ3GgZ69g9VU2IOZd0W5chutaGoba6vc59m2
GviRSu+cktjrOZuqL7ppSUld+KkJbgUr8NQf+wU+x+ZcYpU+4N94yl/Pf5kajD+nwtAUge+7j+MX
7KwwFUMIZwHs9Y7wlg5MhCC1/0yY89S4pn6UUIZ4dwNEInqxbAy2UqDi65IqgE8C2aGu52DxNipP
0iqWH7FRFOQ3Qve8HR/ZM8jYmpma598ySO2viY0c02uiv6DJhbP2hd6CTaYsIFse21GRDx8qa/Tc
lAdMtQCOpuQn5Hx+14UfobNRqv9qURvnK+2iaNx2IKOMH/NFbpH9xfrmZZEnsnBPSIa3bWrJbNCQ
jUOxuvt5nQFA9TVN9e5N5p1zt6Fzn+je7j7iO1H0KWVUMUpKMIWkQkjTmw+JYKNyS1YqQzwRNU9V
EmYy7etNCmoYKccSRtQpDeYsclVIvPC2vhDiNWgo6pxPe2ddyxrWWOyw779M8rRu7WYQ6Kw6HyGj
sLU1AsX2WCU9vCWtEt1uGi/Q64ZMm0G9jN9xRMmrWsSxt5oPg+qUFFoQUaJXkbvvYTX3QKUEms+L
BqY/noGmUCEZv3ENSfdaOlzzhtzde0HPHbakgQ4t4+Ew2CN75iJUunCmGeFS9aATCG+JNNBEtoFc
qNxYCFKOqYWh4iMdXgSp3LdmG/IFvWBIYRz2sN3u/76ss94KjMTArPasw3mLK49MR2t+M5Dk6ytX
LIBLpHpX4xxlKB4wrP1ZaUDp+u/Tgim7y6KJf+kdQ6PyDy8nEHNcxP1kAMcPOKmUDqllANJA4crs
wY85ffDxzmQszsao3smRonmcklRFNQKjUapkylhayx+Ozn9+BNDFI9RoqPXa6bdTYI4fQKyfyPmY
w6O+suYQdiXkdNe/CZjmvgJIXa9ekvxCRHDmgkYz+F2cZAtbYfmc0seXePti6/9iDCnEcEXYtSOX
ZQHnyHMC/j/K6qjiEdIuzaG537Kg2KQfutyKDAxavJfhaEapZqYYNpVhD8es8fahQJXquUwmaTwB
Y1Thv0CQ2GSch9fr1zSO7VnqE1+HsDC4t3NIc0GSGKbRsB6hIx8Vy592aeXS38lmm5WBtwbs3oin
kGGYsROCCiyW7ZwpCbH8XBxUhidsSU+HfjlWEDNzT7Lb8K1oKKFe0SRgwO+jWwLKcRC0Qiex/9BQ
AGRZQDGiBYp18pOTgVBPDHC2V9X9AlbRDwkCRnGf2pKTGnNJIpNOKmozWZJnIGz1HUiowvz0G/I+
rUUQufjSOFjb94RH+0/bhPHnjGO1C7iQ/MLy9jsthoMl43UETJKXDUvDYP/T1DOLIvkBfz2m4QSl
N6jlqRLxy4EKdfAve+FmjzFLgLQT2n6XB9GDCBxjeafDI8k7WV/PYYZq8yaD29eTAAkbUve269L7
xw1NJbd9SBsDpx/HSY3tPtMui5fPMW2HPWHRHqltf0CvizO61GmosMDPX/rr523FuX5U7tBwZz51
OU0OGoaStyX4BZbG84C6IYb3Cwg55wnaJahj699foeSpDpIqbSS3Jb5JnjhLPYR8aXE97UxaMyIS
GAvXsYiNTaGeZFCqm+OReOq51/z8alQrFpWOxEzm93cqlSP6oGs1MHwyvCD1UYj5WhdGGnNK3fvH
XYNAKV+UTXbPx+qIcCQoMAkmzvrM+NWYYmX5/+yITgMWSrFAaiA8zHSF8cHIprieSYlqxcM5tK6v
Cn4ahK+uc+BCnq83I2Tq4E9JaAHefsSA3n0c2kJkfEM7NDPQqMRRrb2HZB60mQkHVPVu6hy8j4af
PHIbsO5yO3EWMEwtORYH/FN73ale9HtLkKJNvdCx8QLOrFF/LdlYRcbJJutpVN1kz+ArlWaP7nsa
M3XLy+mf2rw8XELKun/tQKKKAeZyZly2A3QwY8OO815Cxe8AswFtXOhJgIhcPPeYxaqFD/bxNBOH
dc4sfNp9Etbhi9uOrxM+iOMl2NuFyKcdTP96rGi7BLwlAG8V5dtPI08PpP0+f/mAI5jiAOa0Ywbc
t+Vh5c+CK6ifnP4gOWt9Nd2znVRWs6UuscPy84hZ+lBCmXBMtgeE4iAbjZYyUrbK4RZVhQEkRGsr
pT52rVHNUcQjacfklXq/3YZJT+t3sI++NfcVTUNwO1QO+TnOSJ8kdgl/id2EAJND5e9xkHmXsdow
CMhMRBtDD77f4dXfwmRfT6NhDCi5qMXXE16yC/597gATvFC7XvuJz5iu4TEMrMZIm0lVA/THPbRi
ihtUBNEG/6smpKwm9hHSpM3OqWO8ydn+TR0ENCQjYXjFYIvTxp3wyJtAo8CLSmVf7yDrcti+m92x
XI8dvyYTejLJw1jLKYq4Yf8AVkwGotAgMnrVR0ymIjlwg/0vODzVU8dFVzxwxR3zzhU9lCd/ON1h
kstyUWRT9/EWdl4A7VwBzO/mEfFtt+mFL6TgB6eh/8MpDWQgqEdct8pTf1wA4PjytlPnQF4xItA0
gD/jS07/WHLivC5mDfs+Fc9KFX02s5AtLgymWur7JoVHnhkEdj4762eNogXwix1wY1aP/IyfXOs2
fV/BDFh7sC3d0pM1H9J0+Mifc7He4oUkwjdhapSHjk/RTN24egzJ8Plr/uL/3mKUmI/BhlTpXxXc
SDCSNR/uPqmALXja3WaSQfmzX0iZ3g580y9ZimqeatCskKklVGVMdA7mT8fcLFjb34J+FqZTF3+p
2y0PlpdJqKc8D3VLDoP8SSk5OLAKdYjP0xGcqr7OLI/WbGgSoRHS2xlp0RwyiU2h14AZWhtJuSd+
MggKZZIBGKd/JlKLTD75bk8Ta1gJtbttuLXgSvN6A4JCIBy9AqepFPi/5jdpUKEMlUfEF8847CP1
lohbl4qv9dbNXKGTtSkgrE/+LQ8YqIxtkIzFx7T9xFHpdZwx4WYmG8xhFQusrjPfm1sEioo4WY9V
yCO/kb6izy1xziQ5qeg56Sbfd+S9mS0lJ60BvxJYPAKBTIDIr4ZORi3HSrcdEqknDkhzH3dnhjHr
iNfxZw4DDP07vlRtlnuUWgAFPJUkdGY4ZMvhQeDngx3tudof0rNuUaU1Pfk15h4qRBRKmhWeLF/z
lUk0Cs8i7G0gYuLn3HxPAjRHsoaHv6jB/FgNac2X+95YKOe8FrinCZEOBqLLHT01Z7k7+OFcdWm8
72DRmnwC8H5BnXCZ3ukUr67hPrWnLqwwxpLztTQeFddhMG1npLbV0FgkgJqMSBs86cn2+2h+XLYF
pbAtoW/A3x6h7q4BbGXiLCH5ocg1CznB4RYaqouyzF9cEFnIio2acEVH9X+5PJcYKV1W/wngpARF
f+5Poj8vmr9x2xH7x5VEIS4Q3coIxa5O16MR9AJwND1aR5Y8ZuK5pzateIUHupN1cdBiE7Qzjrnz
J/KImCGYpPJyZPlC9S9UlC2lWZc8u7vNSWWbmBtoY9Euv9epRIK4j8P4YJ9WyjjIPe5VbYQ9Yrql
VhS4dv0YnfrfwZYsZffe/YDY5jPwB5OhLSFq7SbPLnzXneOUQSbfsol9jufZbawQSugRjUj64JNw
+zeIKWM8dvA2B4SYBo5jJzxhadoQX68bTwgO3G+75JrMcLpWl5uLti/B9wkAwf4c2ByRUpuq1+ll
N8oQJkIjGKeuTHFk+k/IMSTVCVZdwUsrja2oayJS1AsG4Br+/ppZfZUnpnIxT94MXrshWCmmVDnp
Zdc18Js3MkUtYQ/QIsz3IGy2QUCb0dgS1KZ8k4qqDkNc4CBLDb286N/waUouwDxcwt6ymn6nzdC/
ZUw+lAhLLTNtXr4zy+vmZoVRcJWbIyZmqOWmPhHgsY8VlGo4h5xY5+Ra4h0OwQTF22KxpIAFka8T
ZEOxXV+KXhwkpLoMtA7TYuQTNqLuSiTqfQr6zPkcHe93Nv8k+zPJXJVQtAb8QQLxLQybhVUX4y3I
1MOaI5JmYHF0NiyP6RnYLpjlr61WshAHo8U=
`pragma protect end_protected
