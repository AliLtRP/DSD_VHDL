library verilog;
use verilog.vl_types.all;
entity half_vlg_check_tst is
    port(
        c               : in     vl_logic;
        s               : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end half_vlg_check_tst;
