// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:35:40 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
JXRDXgHuRWQZpxpglMyp+JUciZlGqZTjyCICRpXzjQfhNBoCdWX0IncLY1niQqgP
C82xCIrAAALXVhPpVCz4Q1ykt1ZLBar8r+2GH/yg4YW8IdExsxEs3YPTzDPMG5Rq
SyKJpSz0IfsFH4nzYUoL45CyO3riuLGJNzhe39kguq0=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 3696)
RVlC17YA/q4CgoCkCs9YxkW7XEWuNMhI1k9zIM/jvH7JaCIV+0OQ40vpxjrumu83
5DwrQym7LzWESwVDPy2rojKOU4nHgNsKv3yZ9oWi/XUBYEdsITHFo1kZ2n5N8nYf
bwiWcxKY8vxN1TjQcy1j/mwEnDBn+pOgNaAAT7DDRMkNCdzw7o7GuajekANjABuB
HFMUk4NKmt6rdf0LohOLWKHN1zi8/84M2nmAMX7KbX5anTwxwLwSxAJWK+g+py9X
dgN5w5XbbCizziGdwEilpwyd79hEpeoJy4yshJ7H9rWJRReZoUqNCSitPU+b5per
jk/36RjA/DLjocWvXHNUnybMK6wzLApBYoE3mp2IzVOh+4WptIlc57LZb3Boii49
4D8Eh0l8CqVddVjk0C63vWP6P2Oo5qwh8VQfv9U9I3sWCfBcc0EkQJuPs2Yoy1jM
Ih4FBvSPKKPz1RDJ3ct9WQXNec1vMxDz9iMhM2Dmz0MlKBphBHc8H7gwifGDYHbe
FRoCHx87NwntA9M7gwOkmEZmo5mHIj9xqSy2D+dI4k5ZnRrCWTqzpPeWrWIKbpvF
HTR75E04J0MUwkSVK87FXASDEA92HWSXTnli2yictPUENXyI6+1XBs8OzE/4PcMb
QVtu3ZgVjzqVX6lvm7+knxeLPxU6uNWQTQc3SanWDNNJ7VuvnsxPhH8Ebc9gAVfg
fuOZ6a/+5wjfXEpyPTwSn2B9lvUxtqCtYRkmvZjE3JxbzUaA9f6OMoCkIjmzkMui
hUs7+sr4/h1C0Qow2Ae5eA30PfGLsxjEeDiyg5WuV3mRTL9FW/LNPAFgeYT/rsti
l1F4WGesvnxnrdMcq+MU5PJ5RVi62FEQ+eg+xNHZzYrxXICgC+ZKupwb17D5UM/k
TS1sUN9VUV43YPdKO5Jr+f4nwBira+35LmgP38QkSJBp3y81FuONiXvIOt/IvHf5
aM5EYUMW2WEfGlDD+JSOeySjaJJMMpRtYUhLFFifIrvzlTeTocu65rOCMRZZRIN+
ggNpftrJReYpZbmYxM1DH0T6D2HMrWHT9/nBwO/1q3uyy8nsosz9UwRA6pNnIotn
12G0qScxAaLoe2Kc1/L/vKLorpLAyZAc7VR40Z7rKZ8mQaCwZ3ofECWgBnUSRaUn
qUByvXjFOAHvLsoSbHZ7u5ugaIy5m5YSNwwYxrFZ19UBgkS0t7UZlQfdRTG2XMWs
k7ngydo3xJgTjGlRIJQonT4kEjKR/WwQn89OHLMvnwmUeLfj4zlAWBtDgoT4a7vc
b55MPfAVSkuko1MrTvHAhUj+mRL1oQ7F5amujdXcG3lKpecGzlXsK5izqL1snKUh
7kBPwLUHADbLhHvH07x5lpjIJiLHXX2BG0nFuBZZFOgRzpiPkGSJSYup3cFHKEQu
e4fxiGNBPG4UgCA/MtrVcLFs0017ZV0Zaif2geggSqk/JQRXm9iBn2r2jPAqyEL0
+Eg4bi8uydL/C7E6XZp7o9+h8yV5WLFF0lBLWjsA2vdecBwKU/Q6vtt0oMYOhLku
z1ytcPVY79bwfcwRauiQuVuvr2Ne+HkNaxSV17zIC27aoCBpGHfOCqbbkzf0hKXp
NeIrkoqlqZPeyJDNq19K3+n7bMrOCfRyu7BXdeU4T5UcIMGxpicnnmrCrXD9XNY1
kpUck734rWA+jnz5cu+Mu7i2IEJB7vdE0g4PSBJKiMFA2kwHpu7DuhJXOn6rGHi6
8lCoZAbim7P5fu8uDungj8WngPRyWEKeqCcyBeZM5hmnRi73HGlFRnwbpUrMdfYr
79jb6PIpEvm7V9R1qOvzvK9tavsrWzxFLmTXCbRNxBhvom67V/eJVPIk0ibrdVH7
ectgs/nrvPayY0Sg4PEbjMpBWwIH/OR29weCqJH4WEitqDka8Ilca0dN+zkPmCWp
/M4UG+LHwQS9HLuZjwXjIVy9nwaz5iuzBKU8IB5P3F6zVE3FrNwVYdZTb48Skqq0
OEILroGlhqmsBm/hMdpYaeqTKJajxbjMwHJGwGJj+E7KgAgeHY8BhxnIvlcU6z4n
/MMXf/4Dktpd2Mnyx8OrC8hIbLhQSRHIddlXnaKWze1rrcez6fABA1U/Dy92/jPf
rRQD6Hvdi202lk24tCZaWcCK8n9ALmrW53Mu4WcWK9TcSKEegCFPCxmw8ePFpp3j
xm+BHGazaqrCyFwOx8lYrUYR/xybcyo4Tcn/U9OWeXFZdn1ScPCY/Qwe4OHDL2vN
NkM9UJPUWkofB1j/rD/P//7iVFzoQCEEV9z010LpF66o7tnAqK1xfBIVWzP/undd
Fqb5tNY8nZ0FWmnk0n7gdcZHinwIembC6MjCIxdGoa/meGKxG7DAZWAs0xqmFKCp
WZUS/asmcOzkWP8YZ3TfMh8EawfTsrAjoxTLcNgSkuz87bL25YzPA6yz1fLHZ8EJ
oAazA6MsqHf/Gfhh0HUm4ZDD/js+PxK8cQ3O9iElMoh/ZJ74MXjh9QqxBIOMSRQ8
ElqOlZyyg/KHwZXF6eJ4X6uJojYLLUPWg1X0uUA6+rMyS32mW0aXyipVbNpuuNzK
OnelL+XULKZseZMLVTFb9hjbdslmDWnwQ5PuIIDmNx6lBPc0i/Nz+lsFUmi0SQd6
t6NeHBmLYKS33mVc9tszLaWHRu26gbpxFUC2eS/lmmIefAbUz6XccqdDyEE9ibnn
E8vsIp9geKt5hqXIP2atCUNwDteZnzWbYpAeASyrIues61j0Bixrqo9/T/aLTzO7
IISF9DS1qXRFu33Hp49b08OB+asTUWZkcrva6xdtsSA5h0g9msTFsP6wieyKGPBi
Z/FMr3v3QMSO7eu4i12Bdvh+50uz5DHSaiWyklNh0kT3l+d9EaNIVPH+kP0Thq3S
vvPcwtB2+4vvgJV9+1bSJS4JiiT9rseZvPUA0fl50pKO3pgNEmExDHnSztu5/87q
3bthQ9F2jgGK3uAslapc8/Jxggq0ju4bpGAtqeMMCOen1ASHbOpU8aRAPw07EuHf
YbjF4dHKl+KeQxe0sjcxdcIJdMQ/XQbkGURRrOlsKREK5vdU+EkbFlTceJRTv1Nn
jMNOqkPP2D/5hVgscHHwl5VeUZnLaaTU2NY/jX056YyMCvbF/oR+qk3FG4aVrjzO
iyIF1jKTfsoOo++zWS4h84C8lYnIRxJpuUgd5GP+Lxy58zs3Kh7MV0r1p1Tpu8K3
TJCwdCI9ffkRc6sIbHztS9QN5WCImcHyGg6WcJG1XagPbD7s2L1xRI/2WaTZcJmC
wuzlTJ85Bm/aqEqKh6JZSz/QRG095uTBK2MaR5d/5BGyR5oc928pl5irE90gs1Ex
vOvEd19BY1Hv9Q6IeVQC7OJPW4bsF2I3Z9I19aIP3oiXeNUl5xg59ZVGBF6Vutdv
r5t0XJ0Layh4BFpXbCAalslsbWMqnjZpdFDLm4cvWgdIC7iq2Qj62tKJCL4BLfrw
fp5aOQb4X/gqbj8Rc1Vq8aiWbVkccElBm9s7JUFUk7V3BQDLEeN5f41AoWX1mSK2
UOIyx7cmyROR8jRQ9Fyv65MjpQnOFR2t6/Y7hWUmBOgS8fp5dmP0Gzzp9W8MwHOd
aYRV93mkBhGpXdBPHXaTK3hqFHrQRfueyR92lL3hGWsLBDHW/L4dSUEjKLmhl18F
JA+MSOuqeg1mZQEmPHqkI+OhHQk2oa1Kg5hOnVOd4PoYDuDS7v3sdOr+mXforntr
5A1RXv+1U29sEi8I55xYn2b76M/BXzwzBKrBb2S8OFCrG2/NT2hXfjkg+6SPCjrR
cmfehy4oM+1iBH0mYktoudKwwRGpNqG/EZewzQuuOfqFEMjWy3GSZpHmvK6jFIFE
JXi1SCTBKmB1OTs0lqFX0h7VH/qWQlz46sqO7MuY/umlPRX41Dz0bOO924B4NFxv
jeiQ0AkE1L73VOA6f8lIL3in16rjyIdSfB/X6xcbg2AVelC8g0WiMklFXaLqe265
/FdKxxiSMwKbWYBSMbzrt3ER+3AN3eIpVQ9ESESu8e5IDl4M0/74AGIIKBgrX9vD
h1/ZCvE+XMrm92XKix4ZI7Qyvga/hVZRfAM4YyVZoAuAL/BdHcJJq4qwzTDLHoHL
kwijan7GOLzKHE6Fim3IbQp+Q/1OoQRhcVkcn8eOpVqfApPL8K8I56ry++T3LAVQ
w9vRwSGOCPY6vk+S5lRIg4xUxF2pX4meSuEfpv1Gw/b1A9FiP3G4U8AnuRegu5UF
rSF1maNsN/lQG56+0dMP9G7CEO52tGfRalLs/xKzAA3OpkV1lOw8VZLD+CDMS02X
B3XzvraXg313j5kD4gloomYrjwHPmem6j9nsbJBVF8nhr/57sfdfDH75vEyX9y3A
5DAs71NwzMg17Bg8bjl/GG95B0C7A1b8cPAViDLy5PLmrYB86QEFUnX4Dn/aWMuG
3Fhr+QQbWoVcaugVSP5FiiqfjRbnAUrkS0EWQRhEznCzkhFbd7CxBsvLGWAVY+Ym
f5KBP+a2IX3GDC1KAxOf91RViuqjDP7t7sxmMJSOqI06WJ/x0o1zocuw1KSw2z1C
3MXiEofKs2yGKVjnXazZpEVMunXMlRJqGDfpdSL3a097y0YL7c5SwxdICBM4A38U
HtaYCZ3FV2TCU/UkIUs3h4h0lqZ9y+u1LS4loH56jefiqi2ZeQY5VpNor70S4s2Q
uIVc+podPe1L50P8MdeIQ3u6eJ/1+sMjk1EXK5PTyVhUKAFzfkcPYEeGQF31i2rT
lSyaGHD33Px9aI1PYVdmHJeiL5UI9z7VxiJ1PYmI25CU6Au3QF3Oy7ZaGxvZuIBx
dJ8da6z5qD8TY+7RkPqqB9Xu/MyoPC0JU2AGjtMuxrE47B0fFB6M7c8+4Zlhp/sw
e6PIZYF4nm2KOd74cG/45hb+NnypjJcwsB6YRkm4xdkxa70hpuvi8dB48QI6+U8y
`pragma protect end_protected
