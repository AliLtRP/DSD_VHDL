// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:38 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
pvOZCzZSPtwgR2ohOo+HHb2IRB51a9x4p8z2IVgNz9c9NaEzy95Vd26vsUH6onb5
uhMy6E11O8XlXU3q9OW3//avqTuBFcza0U464H4ddQtDug3PDmeoCCHzu7ScnBsK
/2F7VFdlLUEuJbfyCl7UhhCuMc4yNWEsvmA5qWRvzpA=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 12304)
FlnqEYcwGq2NQtnNhRDmLkZv34HUa7ywlJ06GORaCCZVXN7OyDBbznDesVsEHdDf
Zxb5lhsWc9QcgUiRYECIG5s6ocmD+iNTJtqfqjoaHnzdo9Fw9Ho8N7rMsfbnME34
p0P+HK2noapVjdAOsR8LgJO3uf5r6RrTetWdDAplDEU3uPEbGv3tiyuEP6hh/0UC
PV7lOeKNNNoRQPKOtTjgfuxiEdZxqKb8QMotdZnLu42myG3kEqbIgiS+oH7Ez66f
F49OyqBImUusKZxlNeSdiqaiP2flX6Xj7Y84xd8Jh2+yxziRbfX4vtA3yx0vmJKA
UMtY6anXdTOFsKfWMZZJdf7ogoy0o/ynaHLOE0jH6nmsQiHa9Y+MQxiYWSRSZx2z
vlxO7yIowp4df9k3yvWO5behS78Vg4RLd/mIUZo5plW/+3q2rH/F5v+12hXlg5je
/szO7WlNoyAua2MBITUbDUQPNA9o34B/vh8cmncErG4fFPsU3a/6e9wbwLUlgWsd
falU40DvlSUlALkoAIQbEQo9JoQtOdZHYsxUh1ZT2O0DUh+NOBeeJHQdS0eNIY4z
GJ37cO3LRBbGgBab2c7YnyexuYE1DbYMICJal0W/M1iFgWI5t7euI+gnEZBXbJvT
XNVDdB7eXJNjLKySFmhpgHoyWwqgwyZVLRqKUnpnMGQEpZdPQOUSWqBzmKtwpCwP
vA2f8Q5J8N8I5Fo3rI/1L1iVYh/CHyEJ+HP76i35KykhlG2/PYKtLO8pBc1s7D7r
RIs2c+HtV6hoy5Irp1+DJgWhIv+mzYFAtMLwxtsowAwWuwtvlOIPq9MV1MT9dhzk
cXfNu/AduN28KNfYZkQuzs5Q2cyqvIicg1SoyeJ9qujGe1sdFh5L9oSircXyftyq
jqE3o13GTKGVpAgXAXsuT5ZYHxus+ey3V2PZHocuU/D3Vkr77a8HkdJjqrUwfNPP
QfWMAClkj2iVvwEQwS68cw01yh1pp8W4WNkyNepeGW2KYSz5AZHyTg+eg0l3o9pQ
XukSDCTjeoo+BFOIaJvWsHDA3ikT4rC+Wy2JDnkDwixsUfb3KlRxp16T7/iq5US1
8Em61XQfG4H36cSSnA6gUX4ySki/YfJC9G1cQHwVhOb2F0GWRQijMmYrironWV/d
XX6dqGNcjDFasvqEKfHMLdf57i5vyI5WjC2gAa6t7j/p+jpm+WsE7zP+VtInrJ3M
yU15ozSClpw6DSm0aeuwrqiEOjhMIvSlqzyB2X0FYxMKYOm5ZFyXE6uM//18KPl4
rkBD655VxJNusUuDG8KEh8KyIUdlMCNnDKewttnzCR5B+Itf7mm4mi/j4gyjeKjU
kLx9YgTyOSYxTsjfviyB0gPIYDwD/fdeUmFoiK6zaKghJ27LHSPBPS4S1s2RdaX4
4QY0p+e9A5vf274PXznCwoVFTuFeg7LuaC2Dw4thZ2L4k1JD55kQhCGz9EqIKmhG
E3FWA2iFelBcQJk9vYaH2hCe+y4zI5TX8ou6GFsTf7KSdJRgpcmS13WXOZhVYHYE
Tw8jhIex9yAKl61pbxE2QwwamQptRkRuKGai4EOAkPZkBUqcA0fhPzqM5L7C9Hfy
aaXglnjiouzXKToOCDKgUR2QlB/mapXpmD27+2FrjlqUWEJok8FNwjDz8dY0ZSjE
ksAQa6TpVhtZsrlp5maIcQTzAe7Ox/oBqIFyhjbBHwlS7vfvdqzylXXkEMjozT8x
aMrBHHGlMtCcm/LEL2WaE+WNTI5V/Z/7VJtrVTLT/q1dqIidNR/wS7eBekz182Fy
c7hPFozLOT6yFokREA/hRhk2siM1rtu0nO8ISW7oOiQUSZkRdpK2SuXZ669jr7Tv
L0hOT3c9eY4gp3tnqlPygNOGNQ7nG3OOVoepEXVP/dTeIiOcsF5ieJxgebPSAb2G
LZRlPyFhQ7wT+e6SRLe34jBp5l1jDRKYLHuoOCsJUFLTSWkBcvNJ2YEi/SJJefCz
QIncb2zggL7CIYCgPh/8uTSR68l5Y14uggzr+3VLMU//3jeevE1JM5MEUf7J7ZdX
NoarRk/tBesKNBYaYkfkcPgKbLKrEt3IEo28a/79kgu3Gripdh939vmuH8gBWb9N
1cGrskLp5fELvxbb/xSEB0ZwX+wmtsH4YJ/Zo53JTJNGlDOM9QUEyxHy7jBbkBpv
YmK3UKPg9e+LkBL6dkuyLAa/kYgROCXHKc2Q6BKWaPgEnv7Bg6KZuhT8mtbYJFJ+
3pMmq59h/0oZ3nhj58SiuqMdVbORM4BP1XawyRNbJWAUY6o7NhgyWE1kBRsdV3f6
kF2H8m4Q9uQRzoGgLbuTCFG0mvrMybKXPPsrhbkRf65sxM6vJPIwDMFPOqbyvcKY
bpyIzrYdoUHdcjIf+5lDZvl5wwrNKlpmwZDdUqbsiVC/nR6n70nu7coYKNvKIa1K
HxJ93PEba89Gx99gpfVDbRJZ7bvhduozHTjG/oAr52CwcAzT7rTUntLVrIxUq3JB
ZHMGV/85JxbaxlJqv0HN4SRAMBlWP5BeGboYaXRzTfJg9UCAsUZELqJJmul01UV8
IeAEVZ43s3Ztf3U3PZOlf7xz1GQZUVc9wbf2TEzUIHeZnmf1BJzLY61gaJHYvUv5
kN+SJ8MObaohtzKxj2vWuukHOIiodaPr0JYa04gyKuAmdCUE14gDdj05gZ1gFYyU
RHnEVNhiN/ioU6i2XSYrPucZz59BtMHNDGfbux4Y3FbS2cNls8qleikggHCtNVgJ
aQflqcLLFNKsXE9WEwnN72hNRkAlywnjCgW45/6hYXlfOHDBw8197x7lOxZyNcTe
NOBFJ84F0l2Lug7f8l6KxIpcBRpT5WWdmqOMT8GzVflom+iTJr8mLapQMpLBn6OQ
MVmAOzFJDYi4BOTPROZsIphHsvduhvUcA/W+a8i4asjTTl59o7+8VR8nB2XPBZR/
S9yx4JcQJHLAt5KAHnY8RCF2FwuYeqphQyFtWhK1Sagc9O26KBycAcEixoAVh7o3
OD8WlIfmsQcoKh9XC0psTd0HmQpuankkXYBWn+D1HZLfkwEkLCjchLoSyDhu5meR
Ml+Rvk1NkS3xykDzuYMFcVGmAE2IepbYwyYwt3JXqqUS5QIA8gSlCCOLov2Qxk83
K3uF1R+vyqN+ZLE3zm3kBeSxOszY/QFAxfNkjEnnf0vrn3DGvzjITIvGFkU7Nf8R
U14CJcpDVap7S50oaeOYR/gyLEaDnpp9eXeb1SE+NAJHBo2/MQp7mYHj8Ld6QeIj
wZ22zkKT3tIqLINmN4vGkwaV/GplkBz6RU6J4V2dbouAAF1mBYlx/J8UJX9C0DZt
t6S+w3fln7SCj7CQVG7aXfyTMkkZtFL7KkaeN2fqeU3I2GIDKn2Zs6AyPUSvcXZh
k6uD6a2Taw9N/6ocL5yMODtGPQXrtIc+LHyxaHq1q4+SCkZiCM7yOBc9bQ8l+K15
1ge+92LYnoIf7bnQKdOfSAdyk4mJJE6rWlNMgHOtg8zQI4gBJfvJ/ZLb3hxQCWXd
mYRC0xbU60tvfIgDIzL9co/IQdLgY0h0HzqDVfoNrveFLUEpQ+bkBMkCldntPaZ7
Yq2sipElOc2eRanm06/OpnzUGevjlaRf3fSzeeaAoJpuGOIKU+UpPxbQ7+dGsQsM
ULnypwP+rXfE4coPRJLJvkDZj1rAffnUIJskTKoLOqZ2L/ZD3yV/S0LclBKbmlSC
oEBQt99uu0+UIkUEUO25SSThPGyqFLooIF5rVdsRjmjy/amkUYcczW+pFs5EW9l5
qdmMUSXFuOwBNatpfSY8IDSQK2Sg9+pRCWda8N+6+VJsLMsJlZ+iP1DsFltdtJSy
ihl9NBzaJljbxDl+VnVop12t+qy+eFsWYxEuDhfuSlcEdDzs+y1XpbsiLvjaosqX
RYWOanZD5nQgV/oiAlQhZ42kMZwc+e2IKzYAMAKKGGfhoU5R/2HE2eKB3C7gwztT
2sXS7E0Wigydjf+yOFLXiCOfgypJCjkHFajpXDqKsPxTyZtPAcIHLGEcqPiGnyIc
1h20bDujZJqXuF/4PCnPzW3APpHKceBR4L9XLU0neT+oE4PBe5qCvImo9i+fqCwT
76rcblz0QOUZ2TWpZbuG3wZQgTpx8KIOjmbInoKyzaZALjBWPwgyQmIt3GOFH52Y
KMzIW+X1N1CzQ1OMlaxTf6qs0OaJ4EQbf8rtZ/iZZS68cLsMU39JrQyPaT1+BOEV
PVvFRNsh2JF9b5hmti5lBw9kIXfziFeQS33TUG1hOdNVhtNLBKYfmJKaPMl5pTGY
mF+ZP35X1XR2J1tDLlOxeMwHYExwKw0ONpJg7945TAE7xAh5UV+Xu/zAnGfSLNg2
jt+Ma+HT7Q65fl9M/TRQNrT8jhipHvGBs8JVc4wtlYxPqC5tvBRb+zTQiEeoxRMj
1mgb72bmcvJNzSfOXmJHAfckIPkCajXjQK7EK2Q/rQquDeY+T8CXhvpFH3rNmHUU
OqMn9Xn29265bFwsY0DZsbq2ncurfOnK74b3fUamwheeq/rIPTYsO7TPbxa6of0X
BXhilPwBuaZKebXNOdKa0OBlpA34BKJh3Qymc+aFiUCYV8IZeqQUrqLUd5NeauDw
hexp6ohpldMDYypXrMniFapxhDMGTMduOV0mIuAd/3VEYwAqlX5b6YBEbFTZcIQ7
tBew8tSOiuV7ywbBCTcY7JIDEqFfBBzIsnUYfGtWXuS2GNkLryOSRST16HS0P6QC
EWJ7k5M2Cfgd26X8PNUKpJxJfecHpKa033bdOqZc8KFdxLQqCFj2wvLAUzDf4B5b
7sR0eaMq49SgHlkiEOMb9j1OzV5drU+Y1mE8HRP9enK6uhnv8ZZlxJVy466VIV1u
Tg5zZ5PNY5CzuWe1xFr9sJxEf18cOLnKJCCf7cOUyLjUP86PbepeEIZ7mWvjl4mV
ZNdtNM/6HdGsJCfVU2qkkgnp80u9YS+38n1fkR2hjm+ppIuCXOZ09b1SxnJaI916
9OIhY0CqdOSE40MbUX2NkjY5efr4EDpRXRo6EQMb6U/al8Nu45xVDi+jH3DkTUlE
XgRM636kO/dTOljz+b2vTPuomDzt0vgoRN9xoyGN9wC77zafW1+a85Z7JhWQ+L1z
NySWB0ShFH3uTBodD10UeGK4gcG7x1rDnVQd/hOQTQS4O3Bhxon4gMLlFkoAc89H
TYMAXnNXkK9e/WVfGo3VzaEehKGr6Kv54TbmtXLUqPVHEF7og8xIoT1XVU5PsM65
Wol4S6Mlf93+KuCol1ACJzbZHBWEm+WBmxNhWjqELHmB7BinRo7iTE1fjC8L+JAK
VRqEDmVB+p+yTJsBdm04lRzydQjweignm5JC+voRWNerZMKnJ7hs7NHolq2be84Z
JaSs5o45RnkIiG8ylwrJConfnNM9FPwEhRM5uXLH1HYjoSNSJs6BuEBAR7TvhFEe
M6XqEy9qd8iT67DwahNCxUTVcQ9yGPC8zTkKZ50ob07heNyp3+EfzaMIlKRqREip
lu+450PYcY+n2F9W1UH//OtJdDLqUC5XkC/IadvWLQce9y5kWOI7LCUMC4YAKTLg
zAIZoBWBnr1FGSmIiXf9lB/kLt/p5V97SadvEg3FzINxQ7L/G5Vp1D5tcbzssuaB
Fly4Dy7Y5beJBZ2FlSWoQYeLtp1SH0XPaGZSvS8YoynMRJre3nbIcmEYA6pv6h55
lLw3m6n97lxXmvJ7KPjXLrAgwIGcKBXZPv2UsLg6O1JFNV5JxC/XcqNTR/WxC0jm
0ChvluRDhmB6Z+W4oOdMfVb9K16bCkF/MD8D+2PtajhUKIw/R/qITP3pxbo28tfC
M9GQoz4V530mh8rDGyarw1Ec1H3hjHTKZ8Od5sSKQygVlJYGS5rBlPh92+ZkkT0B
eCSzU3y9lrQSxS2EuX3VAY2AMm3kPUDGfHPCD7i78CTpjY1F32BESu0KqBgid4nn
htBZ0qW9HdniqQe8kRWpJT01V4Q5/GzsifT9e/KUVQZVgsKQmVJ1MVkDxjpG/CYV
EwuZKie7edPJj1GKFVi3KN7D/01D+s+9uZ2NHNdaHi7UFzHSfk/egfeTBmsM43QI
h8C/3iLWufiphRsT1BP9CrDMdt5Giouq3D6dafUjNEzbinvD67I/+1Jd1Qert431
EPPalt0mc2jYq3PlI6jFAo4Old1lzeYi23iUX97rFNjnsCFqg4jkDyiaKe2agx08
GL7rE+oyUawhnho43+w9V1QgVvEaLEP+ftig6ukmTmYGJY30mxTQMBxdZs402/nb
RBAxHAgFhrBquMblm32EzB7R+zEZMu3oK3+WemoqqwDrMXunSCyntSmi1UZ0CF3Y
og6m/RP7PyOQqsXIy00fMUsEfy1LCDrV8WEPBym1ExGXk3KGxiuMzbIrqHqA5Sne
YE79fR+//q59/koESTnyaHqcoxNv83WURVkVxQd0eN1cTZ9TlzOVzBrrOy+ydENu
ad1Sxmw2ARIBSTAuyWRKj5+CQukVH8mZj53c8XHrjoU/mEmfeLkqDHxNeGWYMceY
c4jVOysDjo1BF6jMEmW8Ia3w9AZIc7NiZrKV96PcNn2zZjqzpBxZaibACUgFWSev
4k/EAqWr6oWrvURvMvp+qwogHP8DKapwWWmFVwppBuk0vmXw0ehqqZikKZ3C4pm6
U/EHOIlkoima0/wE4IkLy64hYTyKHIf8ALroBwmBNMmIoUttIDAvSRDN4Mc61aPa
sjniFa2fApOYw2ULcKtRMIAQGm98j92FLVu+ThXcUnjMbVPBLrbafqznz36CNSs9
QflHFKLk3PxU6D/rR99diuYp+zEy5M5PBCCBfBTQCMD1GVxzsoQwnbQu4p7aOMXg
JeSqTs+88sKkUQ6ZwGEd/kWG+ppUcnD73julnFuDNcTCWq7IL4fe8rwdJGtnbl8I
zxzjYM9nV1QFi9mkjMrvzwPPLh2CTXosypPMdkQ/d1wiyXoMB7ez9/l5oQuTiku+
lkXePL1VNTJKeBjwYY8NmZ4DTTpY+KCemPhoKCf1fUEfVdQVlr8LLDRCuOxGKX5v
BLJSiEzAgpUQ+ICNSzSCCP9y+uXZis9UkvmmPgw+pvDTKmmxNSxNZekf80SRO6Hf
pZA7bHR4e188JyUmgaELhlyt5ZN+XfVp52KSdSDdzze7cA6CAmMER9DhmZG/lh3Z
mEAzeMrdXvPCkPHLpkq9YUxS6PVzRBbZYLYjRTdDHm1ZOIVtjYWMybhRCA6PHG/e
oe879KpMm9UXag2wALhZDbvZiqHC5Ra2BtGF1bA3TO9cKKyISEYoutlv+iGV+a2C
jaoIkpr40KOVkTQywwFLF9208lbSl/vmRIsZAjIC4vcDy/7ym9NLaZPEr4uknwtb
gJQek66JMROvVrESQwiddE1ood1k2A0dsN7dmVtQ9xOpLeLAbVwrib/9U53x5ONn
CggrWhikV3VXvdghzi01Iqzctj4T0QH4MywJ7RllAMku9YtH3fwWd3EYM3vHxxKA
QU/MDLoVDnt6KtNl6zTJY2sRJ954w37OGRym70CWsl6E+MKAQSYhcHFmfNgIH1yE
UhZK1omn6yoQyBcPjhed/KfyV864EaUmLH0oL6ekRtrGnhlxNy+aEgkZCx2gcG8H
jeoAK70KxR23eu4hsmmlNRyOPHxKptBzLkKrJbK0tpSABVnl77F1T4NfYNkUFhqO
oWjp5/TPL+WY64ixHRDVGVWtj+txRkK54FzGoUa+76FqG+nxnf00Ni9uUuOlPZqr
EZLpQcSG5IUgyX0x+ATJHCRhCq8BzTeA/n0mG0l9UNAHIynRrbsZ8mVibD1Wgdx0
gOYXJI1l0D630zVcRL/zMi9069YCAyXRmobTkKyz1M0646NnGV50T2E7nJXvczN/
9QhV+gA9ibGPacP5zE907ZR2BfpTfZutYYSaw1hkR6rJB7l6zsyAZ/NKTd16kX2Y
uHhcMFKyZnX4dDM0B8H/pB23IrFWffpmO+FGa/aVROkWygdswdKzwGMjKv20vPN/
arciqTLUGvc90M80ZmqALxQlxMldbn+14I1hzM7r5MXZHmjsBauEs7NuLc334+GU
A/RHOUXxUKmVHQ8Z5YLudyfqs0oaMKQbi11b05+z5DGtoS+gPz54Vt4u8yq+bk6P
S2vfPS3MrzZNt+Ge1P79kNWxu9VxUQny8bewudzwotroSGEMiC7Xr7fbOJHsOgDO
78MJ5lQl/Y/cEwEmd4htzleC1ckhscpPKZvSzyksvVmBdslM1aVkfkVovWve0zeA
mwDHiZ6x5j3mbEKzMB9v7URw8maI/Rva3pdI7u5jQWDYth+W67XipSr7unMOsjxq
wHeouvF2rW35E6rO8ZvDwTozSCdaGQRRb7lV+NsyJ/pgSkIj27/YsBQH2FpeVQ3G
UeAu5SwU8xvJVez3NuFl/vSMdRa4I38ONNt0X3WZ0xBXk0N2huB7A6IfZNzC/VYI
fiafvDNpJgWJCyqJDwriPHjjdLTO0nfbptDu3H7WgrTLK2MDOtvqDRSt2HxJh6UP
B7TAN4gZd8WOKvwfwRioHsLn8uTTD9PlQQWqXus6YZn5PNtSObz/9CeH018fAM+8
WTojUDvLFWahoBDns/8VwIPBraBbbxtc++S9zvuOCgvIlH0BWxFmosRw1iSIo7AA
Ec3/zKHFfIHVWaD545cWle8tMU7kM/gL3Ifmhv2n3CV2T5aAG156QMCB6MZep3zQ
8J3H6ZI2AizuQC25Ibad7LKZZQyIv0cHEusT8XfpJY4lBPWCqEwFoygI13exlsu/
N9b115A1zSD2EDS9nX1K0Rg2k704voeJq1FnTGzcrELGSxyHr/hC4F3iNxKVFS99
WTwqA9poAJEXHbUfAFPPKuejNJUoJfSiWeQsh/+7yIjDjjtWUxg9pQM+xWdcV0zT
MtkDmLU6QbazqmhvW/cZZn4hOHE+OgKn2lIbJOS+KvJ3FV8+huDPNDi0v/YZG5cm
TDsNJv1b5QQDBtKT3kPhMveZh8HZN9h2jXSfeiBGrhMm9Te4yqs574SU10g43GFa
X9EJeyW+FXgJHsRRqnwAQ0v/iin4Wa4CirRQZ9+buvP/1vShMrHgdjxVr2/QUo4r
KdILYraxf78/+hPcJLDgNxw++JqkjS5gRN+kLDIFOb1tkeCXAWBAcR7PN4fex+im
oDzIsxRRhnfIMW8R0LAtnLrtYlQvoVme4O2GvsP1fzZytkDhF9x7Hhe5SiX4nDmS
m3PCG7gO05gPC/QsGAFiIpsTT8NFFe/aLpyRdFf0TCCEI/wduQ4eJdHxkH1GpFBq
/9MRln0/PZ5B+TGKVa2r/izTKA+KAGYv/YHhpovzsU+FgeLEM9Fv9sH6g/N4JGJy
j192usnUPwl1w/Xx4jB9RMidxZaigoHkJe6A1fNXQROeaGGPN6MOMQTO+qpwWi8y
qOXnQVPyPPik6lFmXKYCrI1wr1pa6cdRgV6mjHvtZzVJn3KBM2b/g/QCDDMOMqjO
pTsZ1cPDPSBqhArwoB+B6blUSSL/iidzwbBJWIUrDyYrIvq0R1SpvlfS2ruQEzd/
29QqN3GlUakalBCth0gKZsEWy5bwfkUUznmKkVeEJ/l2BQSA0MtDn3K24MEUzsXY
xscRPZ4PpcQ19W887vPr8WNrynEnkWgj/SAHNkggGvMIkXL+R441fcvMb+rTjTCI
3x91avh57dodEZlabkJDGXtajy9DTanPYRqwvCXXPI//858euS78MOF0SDnjw8KG
Oa8Z1mA1kzVKH8NFFvwR56NsL7M7Fz0e9I5jXc78Pf0GWLGExGaABygxYEu+Z3wq
2FAv+1UTFd2I5gsKu6oecrbq7vbwBslkXwHIFCEDacYWwPdghqihL1j+7XYygF4H
JgHtWresHaaQK48eKkQaOnHoYOjWrFyoKimi+8VtnCmTOgTwr5+i13F0riqnCOGD
CqMyg1yKDzQc8iPODUJoPq5gYqcKPdYIu6SDhva1BbtV51uMQcLT7BZU0kvtExPj
PCRaZvVhnQ1xpqX82ooh06Lxg4HKJ9nv8a/WYV3n1hErydnm66ApEMIuO58F0I9g
1559xWY/e8BtbbS+sxu49wgRhLYNOLUPfZu28tml1v7u/lqp+24JfPZ97KZCH5CT
4onjfOAFI5pv/CB4wHF87SYVTSIr9DM8cR8ZEhqa+6DRE253uiL2+1O25FD+PZAp
ZZB2XmapY6rpRgop80AgM9PMndB9K0U6ezuX9NjKPwyzaTw3qYVUyZLRR1d8qflt
uA1WxNMhw8AHEF6IYl9u+z4R34i/nTbCHWqnd2852a3d7DTx44RfVGCufQtuY2JA
/AAzPWBiAT98cGS/Q3x6wW1AW1GfuGXYWMUMN6baeZ2Eap3xKG4fluae7bFKJGJi
J/cztTAYSYGT6wtvE9uPIX2pycf2NCxKvMikL3AAPtHuHpLswOyWeil7aMLhjKRv
gtUtUvKS2yAAbd3DrryZaM/EdvvRg96u24uRdY9m2x1TiU6LQBw1uHc6fA/95uGw
ZLQNRF0hdV+9JkODXF4Fb5P7988sw/h/HmFQMJa383W9N/SjBZsSsCDuu63MO2IA
16jdiIkRjlJ63yWV5+27rMuV///HOk6vE0fA3ZL1unKWIU0A+D+qTppA7vavdaZe
uPi3UZjbjdz8XOeKd6pZ7Nj3nfXHedZ73l7JkXeLcqSL80/kupgi5LNICTEYvdIx
4ajBlTCdquSOxZmga+DP93i8DMSCkgH8UD6YWAlS/JKKcxLJteKKs0EFRY4UTn/2
XKNW1LDIGFHYkyhsmLhpHX3akcOC5RuHzmrD++XH2c/77xPhN4liid+dLER/kiJB
Hh9wWuZoRnaNfVK8sLmt2lnOU/TjvSwARB4yGFDoYcvasWIadKyuI13qbxj3EdhI
QGKz0HycCQMJWtLmgroJAcoQY3Kd4mLUmcK9OZR2cGSHBauCRN6Fq6SBLUSKDOq3
QyP/WCdJhm7Bcs+Qu55sRsBLtx6xfjVWanmVHPB6GIsgTZtTgHn8DnjAWHzHNVO5
6QNbg6+99cY7mrjzhY8WEgfvU+x4FlZwSBdECxo+lwswgP41Ck+kTRdKk6giCSDj
lbek3P+IFHaqJ4TNwukbV+6QRNTz54rM12x8evOAmMWf2/JDR4246izCor2Dsj5U
nBAHN1VD9XndFHgj5vCRR0DaKQr42tRvb7qQWtzwHwMUahGEZYsFl1FuPbgcQqXa
w9rbszXJM/akiJceIFqlcj/x0A4CcRVeYdNy8ib2G1crEdtJ694ej1OEP0cWIN2z
lmXKzqRREgN/Vc8N024J+iA20kqq94/aF8PZzf3n/Y3YreTxfQYjH4Nu82fdXQ7O
e/gWq2DqjPuJgm/KsaRbInJOm1HJV3svJaBYhcajAX+mjOG5cCTtfzX4XDIpN4jR
bDXpynAFYOesXENOX0X/Vkv5XmpOBsBBxWJmKtOu896TdetlEcTTgZPT/XhZpkI/
z4DNTA1xB0czOX1ftm7eQWv9jwtmmZlC3DsnYSRp8CX71BJSZBqCYY+uZKxLBRql
exUn60aECqGEfrAKd0Wd04MgvTnskrF4T3njisUFsMpd9zkYAWJ6+HSFgdcwwsOU
wZ5pJTLKL2ISOhPiY7ETeHHtQnKnSDiAx+peZaTQFhYRgKvCXkyEdQLueRMcu2Y1
Swoug4Y0shmyAxL9weHZN/I8zmZsGw+U1A11muezqQHfjcueLdMG2p7yiMMvOcTp
I0TIX6XDB8wI8wHW9Tnj6ASKRVH5PgPEbVSsQDrIgjDSAGnumO25eSBCR8dGqhEZ
rjtEY3O53A9+VsUGpCtCJfVE8RXvIjUrKERbTnL8a5kOrHVZ0WmHLft5OjNeKPAW
LU7AtocI7xxvG4LKrq7JlQ53jSdKubuL0tpSBaCt4Bm8e5sNFfzhp74JDpEtkwn5
uGD4g6WQKu4RVcrl8TCda4cmaPEMesEDL+iGIPXu974r0dK2P9PjSXeS2BwaqDg5
OpahX2e55rKqjAZmzTLro8oVADQgON0QbLNmvXdq9+Nl4FAR+VT4fct865dwe51C
HWxQzKBWUA3/Us5ZUQSJcgQwETMr35QUBIe6sQPj3lVqphicmCFAaGLJn8r5QBHu
uhCP8ol1QAGnBVGFx67GVyMqx2mHMoqHg/0dFrFxH8kZ3sR28OMOYXMfAJYNdqRG
Gr5EqXGEW1LyFbUb67HyYjhLEc1e/c86086TuY9v+VanMawna8O16T9jqUtrcXu6
uPZGm+tLAs6eZCIemCX3qTqBy+lrdLs9hdGlIfREsFea+6D54Y/qqHNWFz12UzxC
LTPMeJhDCWOTL9wJoE2NMfXLndan9dUQEonL3w2hwie+f/4GBdeh+NInPlfrHrHy
NQ9QjuCd8IpQWSSaL8bbAhWZhecNlSBw31ULKKeRSBWyJy9yKNMHCz9jJYQPbmNx
NmG6xZMFgli4JIZJwyu5F3rq2FpLanNw+ENI69BHq3gmQq+Md9uNiXbS390FufTJ
ARr5yV9+FKUgA0INMzpG3vndg/pT/4Mx/F8UA0TYFnwyPC6WIwQQz9b60anXsdg3
3bAE8u38PFzvSKzp4BWnk/OFlhyGatYm9VIGUqYKPS8OeGh4dGRxkj4J0jP4pobY
CIxTPdCti9qit7kYstNXnQ2j4gfsSDvDwT9BkLZsFi4Ha7CZ9a2Ex6Xxxicb4IW3
YkPx7qAsBqz1l1bkjgXRNgycjA722OXV2705EBpd6tVfQlwLfVV3qQOYsNs7WBdT
wrT069mDPI0fI/M2ZPf0jyrqfq7yEVdl/D9VS5m4tdPdhDcJL3DNIEdX2aNuPGr8
E63LlUy2y30c2AnFVYNGnpgmQFJt9kfPWX6zNVg8qJ4WjM7y88Ckii11ga/WZsZD
ehK/vX0qDqPy++YK4Rt5e6FTfbK8m4I6j8sdTlUrMbqGYTNfTS3Zh+qP7zbM+YN8
Vz/WBaoDd5Php5QkXoQytHkHxKBFYJ4hht1y+nIJ22IK3Voqc0kk/HRybFJnS9QO
MMNNm8zGhNuU5Zj41lTKvBpsRnakUS2Dd6aRJNse4mHo1uvypSqcLfy2EGUAjy3Z
M0EjzRubpHH3pp5Gc+2N0tjlEPnvJsGisg5rtOKlgkiYmc6DDqWxAx9FHbAmtHte
GBEwMzRVffy5sCZMrJzch/uHp39T5RNVDMkmZNoXvKUbLBkbdt+p32SIn257ZJM/
BWaKaMFQtqfg2aZHPB2aEJlhb6DHwuegA/aS2jXOqnS5V1ftNoH3Ax8LTRz6+WZN
flZvCbuv1eUVzD+NnT0VhlwGI4nI/GwpfITBfUQyM8mYwtja7L6z9zJgfmYEhO4E
whgBbQJeEhB/bmTUnTz67cuN4EYMpguvYmvi3bywaZjspL+ANQvFx24y8FQ7sBmO
tcFqjU5CTw7yETgiYphOowhAMNtlFdmcG78Iffljb1yfiC0XpH+cQ8y5VevlpywR
P3QYl7oJmuJZaa8E7BJyEbZ3X87CLUz8npAKqfhKQpeLWF3dw5j4rQqtjl7CtB8h
GWqoHIN6ORWv5p67GwvgRBtQ1IBtab4vzrWeZ9pWbQgLyDbTpuOjXS4sXXReGQMU
fBQJn5W201zbxLTSxBDCaqprteamn36P1pYLDBl++NyZzVPs1xBs1CswooM19mcW
UZAbaqrZN8NH9Zdpgs/GB8sGM5hCTMmKL3pojU6D/OOEbAO2wcinblZaLetsvr0O
Y05Q7ldvhNEoawQJb1FHsXYc/+l33VM24TbIWvD/oOhGgbtnbTzVJ3aOiPoTiKmK
seDTdOsXknz8YsM827OaF9XJK0ycuwN3zCvzU2EYNj+ij96Tc41YaL8rBkLNiKAP
2TXJLpxkyjZQo2F476yibbqGppN+RGcQoqFz19PmJW6Us0yo8Dz0O6LIYPP07aH1
YeNi21ihZkQLX+1n6lTmP9wcKi0gVr4AZUcq2LVY0wZjs1iUM0edfYwFA+y0lsC1
pQh5tkvA6EKqwmJArfxOJld+sUhCBHVSGZs5zTJTU9uYz6i9ryn9S3VIFyD6ecE8
19cSG046YNAAnPYT8IMoCWy+JhGhCK2BJzkrxIBoY5ynapy2FaEuGidk0ez6mAqj
iPeFWlDgivZ6gF+WEt4t3TFR0+Wl064JK6QfNz7yR+T962zS42p1fu+hTBc6su0k
RjfgqcwkEozrK5Qrz6pFJ1AJ2YBs02zyg8M2Oe8pVxMrdd9nA4R5/Nj/SCGcnqMp
tFy+y0nqfwZb+YIcOz0NvmCVGywie+7l2GPcQYeJFh/vYg6CbMia4+YasV/POXp1
ZGlTWH0ggsvQAZb16V78bl2WDkd7EqwEar4PNBSWNfiie8cguj/2dQxN0fr4UlZx
icIlriTgYmCiQmNJ5OqJimHkYD4DkZp/l7n3f6DjBysUR+/gBkED5kg3xVBO9a8D
bXC899ydKkQGrJTVhLJE/EzaBiw/g+bhadd8slBjUbe9qXaAMU2JSOAHZ8WSOkwM
pBJoCSQC+NgPcs8uK/x1rj/uOEO6vCrMSTUqqyAoT6VLvtbT02o4MCijhjLnE4In
GzjclCqe7UKugtaDzK2xn8BoJ7ir46wTrsS1nS49k/mre5g8+PcMZKibzZxp+FqL
2T/Qk3uiJNSefqudHhGMb64DJDTFRmoJu11r9RKsb+lyBih9KoxcwC2tV9JfRcJj
4/H9mdPmaJM+3fveqFyYTk48b+AROaD6slbuu/q/vPgAxUCsRedDzjN3+3vR3+Pu
ujD54hPdP81LUR8phYx19P+eCuqCY92m5m0wVby4jKPk2iZTzuF9Lgz1TXmz2drw
bvBc8jANv5Qv0WGtzvJELcBJCROzjWACRnodJezepwcV/UMnQwLViYm2db8RvKQC
/FxwISj6UuFWUcYQVOax5Fr3FR25W7850XqCuOVGXBSsh59xoH2w9ay80/eXYL/U
bz5PzBO8AQHJbLIaEy62a+pABp5Otv0CzhdXjA0ZnYXGUR7qg3f6wxhOfH3SjmT9
Sc3cPi/MWKYTslRIfqObk/O1RtgDCIKHBFDHA1RPuTKPDNZQmoTdKfFXwV2MdBsL
9eE1jgtmvYVBSLso10Ma/XA4huPxls3b+VMTetWGCy92xemE4e4zxbB7i3fL3pc5
j7uJT2XkKdn/e+AEaOxTpCzOMbchVsAHrO2SJvu3AFoQxSGOIQTRBTgahZ6SYoCW
1OrqSWXsnYP8P0kRe0DXzKv+tmuiL1ibmEaYyAosO5dxMqL3vvEQq+ChZ4ihKy88
o2RKMaCp9AsAtnPtKbdYad+567eFxeqtJyaHGtZMOvzYb9UfdlZ44qp1AEGzCAAb
BmYHQgfLzy9VvluW0naEbiO1wao0X1uMOCeuFp/GWXEOhDeCBPksUZp2m3BjEeE0
/vKjR2GEzWwISun5FcdoZ4QDtgTb6jhOLiuAjXrlseQaywMgMuaAVoQR4Mb/1HPi
oACEidFVyfljbikVGHoARMVvF6HCIr+65uj/WuWuWDl7UuGmUMsYk+zUveZpYQ9X
pOlw7A+9dnp0HYBHiv36/iDmpRNEV6Jfw8d0Hwf/nYwb4AdRDDru8nqTcjOv4HUf
89gC5VDXz8D/ZnzzO217Q3OmvRWhzdsh9Gu9AvhuehHJS8xXerFzx7droTIc97sg
w6duCH30WVKHu0OZ3ZNdtaRP5co7pEh3s+s8SBYAxqiL/uWhttRlE+68r+C/lB3y
18zMSDLDrYu8j3066CuRLuQH9Wgd5Y05rHjkL0uBoQ0sqTVztt9keL59HWUkjJ14
XnBwg0REdSMShY/IcpYVYoBYfLV/GccJyhBF8FsZuu7CkcKutQdk3kCnweDAVMGt
RogRjM4OAjAFgvETYfypyub2qC7l4Yq/BsGoq6FLTGSKhtAjzcC/l7I5pmWXwRjT
fQ+JPHvUroDV3CfFF2R+/z0tN2x7Nyu3aSBoiLzNrn2fnoZ1jfFLnsHEbEjzQji4
xR/khJE1GfH16vhZe4RxNl8E2F+/uj9Gfs1R0d3rENWToUVa4urSA1RHK/YfYlqq
WDpXms2TiBqgcT47Umqxpjz4JEUEB+/K3syUn2vh2zN/3zVVjpUrqtKVq2pRw4Ve
BnjZR+KcROqcc2YxQq0gBtfM09nEyFn2J/jTbSdSoKUXaqRdxih0K9BWqPt35g30
guRO/lKWPvI1zPI9Mj1QPnlXBqE80//aMHejkQ5mNo4udhukvXLI8pC2B/xgE96l
xV1fmjuVwlUxoPMgwiboKoWe8jME5xNaQljk8Bjo7u69ibJNbXLlMzDsl4mFRcWM
FR3QmUrQ5hdH6SD+BN08BJFW7FU1aBenkNIS83WXqypwcaikWXYn0iyJ+FS/VixU
kxHETLTsiWF75G6iMkQdvOPhHx6yOzEbk8RG2CtF7v+sCCmF9Hl06ChvVPRNjPnm
Ykcvr/uVBLgKlN36pDIR1A==
`pragma protect end_protected
