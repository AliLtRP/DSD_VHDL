// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:35:38 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
HUjh3ImSVnug6pBqUvVfw5asFPtaCkkPUjQLo3VXBP9JyTXzr7AHJWKlKik0ALOe
QXcV8b5Ul4q0oVKQp0s+If5KCpNfVvkxhBbBC0j7qaLSAJNwBnfnuh+ErkUB+FuT
E8l8yIuIaBxBFmTaB+A4gP+DrDvyu3+hE2NQ4OpsZnw=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 10944)
XNzbwgk9dCXXEM2NMYp7i1Ax47MkrhqEah1rttAIe+EkBJeBWbMACe7GkYaTxXHK
MzsJYtPzkOPsXRfugFMQ9JWz9keoQ+DOUtUkaG3rfO6Z1mMh36J6QaJ8+5CKqVLn
0ji+fEOY41sSR0BbxNB5ICbabBtkxrtZhHkBx5xKPZA/E0k4s8voQ9aGVw41LKDH
Zd+ahGI1UVNkSHgA8Cn5AaltXELKZl45x5kTsK7nOjiRcdT/dn79XwZv3zQ9e5Zq
ZZRHNLmeQk6NWz6z5aJSkoWfpwiDSHoN+Q/rrAGX5qfKX2KxeeauX+/ZNxwJCOYJ
gsNB+mhBWJwVP/odCCuaA6fwU3i0DVeiGhh5umjc6n7we27tvoscUFcp/vg21y/2
mhKKK6v2V9iWtxzaycVMSmNYyzOp8Ala/cDHJpBp5ZmxDousIXjlou9irjw11ZkM
4oQaRWS6HDcCkCb5o5sos/gsSgIQbs5oE5ZhijA9DRf2XLFFeyYs/icFtl92DtHi
9Li0UyNqh4FxQjtEA4WVoIAg0TyWoCWK2JlpHk9OiscAkpVko4aX+O0cU3f38Aqk
aKsaobbFdWDOMyQHCXGzTkVoh4uB8YRCXXMtcMUVY00jSC7vztzNolD2ZYgkW8vK
LIOU3XvPQ1Al1Q2FXm9Fze/RQcrj70npwzrRYWthH9tTdtaNTaCMlR7AT2ijsC7F
nqjdVR9eDC0oYBlK2KpP8GUvm/FLDSFpS7w2FlsOZo6RU0dmveUyU0vhROI8wTc6
E065ARw230Igt4c0g6wIId0aq/YTx6nTvH/OAbGE38brdEaU0BOUdPzAxqL4pKiJ
azyWK393rY3D0Hpdoyn2ipOIdLT+wLe4NXOoV43dyU6H5vGU0s6cBv6+ONAFFi3V
c1PScxCynIonOu+f8ziq8O51Qbligl6Qwk7APCkL7qEqZmH8TusLdSWw+xHrvKsX
rE1S63dE7vAS/ukd5SfXsM+9j+0Fi3XffjLlmyC55ylXHexlmiFyqHfITP+BHREX
quWMYVcN5hRMil8hO3662gXWR+QRgy8dUwQMD+J/0n1s208U5J3QIKp15GUo0w4W
cbcIuycyReC7fHk94h0KXYMpdqibHP0IzEoyEmy7ZGUWKR93rBXn7HjLMYnRHOrR
8ISE+lR5Jb7MIBWsby6g4OMspb7RzMS0TJ3mniH1fbex+cUhx3fFL04SSZfJO5Xr
/DCw/v8ygWESBWEJS320+5J0dJ0PawzInGBzK9sKMjTNBs6sPCmYUU3Db4dScrSE
VGoyUTAyzkU8n5rznfAaIk558O8PGVQN45FOf+iyFrPm9wFawS6plhgCTeGOHxr1
b+GWrX1awOTsWl4OU7CoTbEscZ8MNUW33fcEQ01jEG6JUUHYfwV6786yBdWYqN9s
pMkXOLHXMJQ9Sd7pXXFbnAFJe2D7D6MZgMh+2k8WIu2QTBtZJQvC/8bAiUm8zsMK
mTaTLK00DHbX09raTbRyrrYSypQiywoI9EjDDDL5t1S2kfwL79McC6UwjiXvJvyg
pzcfkKbMHc/bTvkxTPgZvbbGnFKIYyX7uQyj5etGVAvGpD3b3lMVgFXGVBw1Uh4t
xuFlbMK89zqRrpWjkPa0FCBXvtipcq3Jr7BFA6P7+rKij9eTFxBDOtxsvrPuJXeB
mHMpPAGa3qz8OjnNqHWaV/T50QK/OSVL+tfzFLUav8tpVIVJrMWTvYYLwvul6bDB
aZISUrruTvpdreYieWD6d/viWLDtamO6yF12OviNWImOXxjBfvtcDHWghSDLmDnO
kQM3VSRirRNgQQWikb1ZRAG1STflWDTZ7PbLOLGzzBngnH4RoqkCI8bBAujnH1Rr
WarOEeT43sAhmkrjANIa4y9KXvfEkJd9xGm2SZNrwjKT1VY/rbOeNyGwdRnUJVcn
KI4a2a3JXMPnuS6ECEH4wPgxLt36z7HpiIyByDHUQjB3aaSOXOcOkq4/nD+ucVt2
v037ClKBsCiRnTlBHPA51wYFfMVhcUruYfBkisFQAw2TG7tqpCaif6vYcmmSQT4P
U9VHadWxLax/r45TRX4vkR2e8Hyv+5hm+uoVveuh+KhxzWbxe8letSmIIgNHN7+Y
EbJqYwWFnPzmTQtGGtHZtpdhm+kJcq5+O6tmHajCo/P8RrlKFicrkHfVQtagBFm+
Z7eGBUCfwZ6VhDMAs7BrEflC47S6utC7RO2hDH6o62zxBHTAv0Buxz0AVpHRlLKC
gig3KLL76OKV4cFWViDc4BgC/68+RlfnQayxMBDD7ZAM5YPGUW5Y8CF9q8XdSZuI
G7IjLK+VXrGCIxRxmZcz+qKRUhwpE+SgUzuLsmTNSzAyLAeQ1xE4RsM0MqLI3Nug
+lsZClovs5MKvQP0ykdVCjHcgVmakuFbUPOM/LssHIQEPBUXyy/aW2iORVdBWwNi
mxL9/GGxWPa/E3xQsEYTMGfPAbLFqzeSK+Fl+Thw3vOa5/1My/QcwRw8gQWTvyel
tyltlfQokMH06zchHv/eF6H2Umpwdzd55WR9Io97RkYID9wm0jU/tIAEenDRRr0h
rVu7jACI4NsMtgViOuKIJu1B9UxyGRr4slM50xVsV3d5tQs3l8f9nEP1MorB5VK1
xtVgnAltYS4x6ReKOEsXjQHAt1V1iMJWediVaqDz0CTjv3VFAasr7Y09Lqo4yvDD
f+ozL0V56+WOVa33IaeUx34Mkkdev9ho7Ewwp/X6jiZP6YWdDCpYWlZd5tuT3KZ+
Ws1dhZ5admoArUOrGx3N/JsOHNqUVV+0GRb7+olw6/MFR7jOzlUuEd2Iv7/YJOog
YEFnN2YaQYww/pIJpWhdisO9yrgGORIfyCAOLz7IhBUVPO3O94e0OqQTlz+ewh0p
nWcxI0bBFpFXUCIxUIw/WMBwYFyaqZl2M/svGvuCGX06NMHAvsWEGiSs1rOREK5j
dffz/TfcYzfIFsC49tnQiQHTt6yDSS49it3yUUPRbpl99oSqAnCF9/8QBA8wrAQp
u1/9oEQ3U4LbuIKHXG5m/KyaLBKO8+M8cNs6Idjtwr8T2SwquPvL/LcDGOZnSzVJ
CM3Ve7UDf66uQVgNB3xHaT0RbdydSJLo8g8DKCJYylpZM90J53cBLX/j8NlZgTjv
TM1JPb5psQGwYhW7+0UHQ6XLKKTS0JvEWfMcjhhRdxQhWq9HWLVFHULUjiTfDB6Z
+hvhy18y9sx5kcz9HjRuiXdWwp+2YHdOW282J1ljaJX1r6/HGHnboIpnRUQpv6mm
D86VpsYh9jr466Idae2n01Imv4AL4JDP9gDXzBj2wUlvYG68TubJDSffeMZrXXE+
uA0cQWhqz3u1BnM43ObgYTsoWxsGEez+hpOV2f1/XTx1V0QdWj+uDiyEhuuekHFc
CfdidJLWjpFmD/3VxXGS+eFKAR4eCJP4SQ6QF8bmGA9pegKxZprr03vAy0vKr2Sa
rwIMS/ZbP3/oPeokUgliCpKPYsEwYNauEMP01BcwDBfUmDyumFDr0IjQgj+AUNV1
WpRY3IEmmgS7W0tZWDU5MQo69r/QNxLvX8x6bbFLxb4IalENQsWTIP3r01OO0YGx
Q/76wNzUZB7vJvlM2FEa15A6MzEje/CePD+ISGDsuRgjF1Ktftl7mb2yikJi0jGR
SWy56qnyx1HnxNKYRtEpS2umyawixmANmUXGCD2k340ELAHvFqghjPFCGtj/Lhu7
mTq3MZTEn0kQEP2iHZBgLNgJLbuq0hxw2xfdMtDZ5tKHQnlV/EsWYGPWSZ4zY8bc
VD7YpnlEhoHANbApcSSGxUx4/KKdrthe++kXddLnvb9XlpZyxljQp3jvGeIhoXy8
+RmIUOXJ7INsDvnqvG9D8gsGEKZ9sGBEcZ6iNJO9SrNpOyOplmpaCWTqiXmJMnlY
GUXX/mu9GkJzu+m9KOWnHEkaR1UNcwQRhppEPCgMqF8A01gqon3VgSUvkAturzgn
6qwLqdQb6TdAWSrFhQVG5anKnwTZ7Gbib0RoEUSeelERxfpihqhnaZQ2PgSS4iTg
GEl+oUyEZnGLL4LQOqnT3GFUfaWq+3c/TqUh6FOU9VNFGIOjl63jCScNhS0D1I4j
fMOMZqCvqY+5DA0Nfw89savvEP7yt7SOCWNo2HHGeutpx3MMWvStBCzQaxrrW0xJ
W3dd9QLGSU9SF5EhaU6lpe4pcQrkeAs6DHDTBBxBTPcw0A/6djDnlCejpamYJLHw
s7YJ3Y4URdiurNUsC4PnHW52A3K9Dio+VPFdcmvLYTqMQdklmB38OvwGga3t+3MK
FuC7TaD2Y332NhKD0/tOJqEhNSauo0W4afWY5LtW4pTpx/69Y/J/+bU43zedMWT1
VWPzRDMzmUyJB1JDVjjLq4FbL9wMgDMvDXsZFA6WdOrdPl20DF2yg1tW6k0GLqUW
UWt+CCUJi1EQtp4mFx71HZuokVhzwg6sgWUxRc2Zh2mXMJL047TbwDaOZN5X4jjk
oNzJ9BEv568Q3T5DqMzgbyK/Wg9UqfyTw/PNn4uM1ObrqgykQok9iz37nVB0fGoC
2eSDuvW4Cp1vkdIMBJ9Vjr2NF6cujRxdKjvX7hHwK1W0bqClT/KvEvu45jUKc4OH
uDpd3/l7vekhBPHt85kiFoCE3ydvxvI2kMA+yQJ3e/VuGI8JZ129JJFqOW2p7drx
SK1UiDzWiylY02rRdw2971WCE9tJTA96Ccb6iUn1VMAktKDYOtPMwgqfkSYNz3Pv
95HH4VzZJDZ4HXJRwGyo0rQtp1RMTGXE/pIZOdgV/hdXB+kxr5We2FAjqvAMgPBl
T2HZX9JhiQRDRwSHhogXVcoIyzj/qI4Guimi/Wh9ARS/GhdHlWGofhKP2O6RuE/V
s05NwhHGs+/9LSuQNeCh7Zqi5m6/K11aBfAvrp6gs23ZHmipm0VdU2saxaIePfYi
XUKDtdMwiKxY+ab/+wMvzA4E3k2sZ41EFQFznRarofloDPHM+198oVcwEib0m9D2
mSXj9rjiLeLlOArwf4arUClUgzQCBCdAlKKODorj3JxHVVYMHGYHCbseJj6zM4B5
SUj68/kED7uzKUhOZnkdmt9G1mfqSGfCEN2iVJ+8TjyisHOoYIyGy49r7+F4i8tT
vx75PVsVm11EL8C5vq5bMy96Y7Tg72TmPyKLhCNXxrISwawjn+tZg8FN2Y4oZcP9
oCCroVg8574VTDzpvH2yBMje+2IP9EIttBR72aaVmUi2nFOELICxwxukBuBR58wv
U2CrainIrbrmucJsT8vf5EqcR11oAa7PvMyossugdgdrqVD0G/NXKzKUcCjhR18N
hEoX43mkY2AY2srPPCw7gVS3rPza45wuobKUO2ee+y2W7A4bWlyMObYxbpgow2RM
JKcFDIjebpuySpq57fWQfS6E2EP+8Jp+scCXC8o905qltDuQrnqi34zfwKV29xOF
NK91RZDAZ/gHnyqkFmTjpehntYhfLasf+O+20GLYg9osTJfd8uSlAAcrZQ2Hqm++
nswlR1N4446Vf+zPE4mTb/kKkVmzSQ7K4pw/fe603RaoZEhbv7v4hwNvpPF3lCEs
Rtq9myeo0EWiwOJgDaRkXN2LeetfB90N67nn5pttU0ASuuaTrTNnyTV+jn1iBeX9
9cthlsJ8zxn03Lob1uPX0uVVeYz/SG6XLliMk2IYYk0nBh3BJ/fcIUfs2VWSYxMF
mUUE/TYuo+AFl4F/NvtQv7lfZsNORoV9x5AuY59xUqSkdEg+64IiIZNptFMijqSI
HOQkXZHnZUp7Q+EAwWXCAXD/d956q1TwxuiPMXV5aPJtr9WukPNZ+HkRqTxXOnZT
TGv7lwSt0T389nUKSq+4k5PrhHjWeYSSSxffRV+ZIrZhrN6/rmIp1QsKukIe+tG9
V3b+GEwPORVoNu9Mp2EPraKf58akYEsQLqtnXQ5TvzOsr69NCPiLHO2QnkOnh30c
iMi/A1vEWfT6TbJKtJM4O+PUAqF5C6t+DsMWhv8JEp4jiC/fOHdvPPD5yTAiOonz
WcKZAKqKcb0sJzc0AHhi3LknqZSyU2LVSOnEkVKgsVUaRDbgX9L7htWQWvgU0Nc5
3S9w+7svXCoKfD110g8aF2ONsSN3DUr12r3GlS830orMseFzxci4tfMFKjQpJ84u
GUeB9LJdyXgV1ZUNNLYHmvxKuZj0Dv9Gy33uZ8oYyTILXGTlJBoU73oyNBMA/6lm
oqSuED2aZT7hNxO5vRreLK8cVX3S/Na0y+AD4IVQUYl1J4T+pF3HHaZmL7sCV0c6
pYWsyXdQmHuIhwWQDc7/5GjmVPNlvfTAW1ydzogvEk7hOzMDrTedY9aMeHKsKjmp
Ao3AsoJbDAn/eSamS9Mhu/Ad3prfvonouqucoM1XcVRzH9GJBegD17j7l3ssbej7
R2APLDatcK4UCDOpm42lEwjagwgMTBLBSMXuPOtFLKUGbFkjnzpeoeFcdgPaYwe4
h75toHhcg+SZt/OmfS6ZejPBpd6vjw6NuD9P3QqbxmJABshKyCE3e0tA1TWsd3wj
f1o8jrKF3ZKbjxTrKuH/6GzlU8CsygLq+o+GOb6N7ag4oWCXZhJmlvLGsvErByYU
csa2zbY42a1uOtPjgIMlPGRaKYCDSSN5+yAemKRbiqR8NyflzpXiGIfTnNqhuUzY
5cIZ3FAd+2iO3IyjHeiXMVQ5u7/kpmY88HaPjtAU+iKR9w15CWduvN4JydnJZoy6
SMXlfl6YmnmNx/drHcVUmjPbnQmkWZg8ckJHClrkGhGZTPeGrpQ5ixNcXZi+4nkK
cpyzsKBC1ydfxt+CR7nqD/8GGGP5CMOn+rBkI/dqMGnR2oUqOjTKLl9Zt0cs6ogp
Ufa3WCODg1/lCm/vE0jf2a4nfaJQwwJ0+WMglPN2fWelcqW0NjGfKTY0YG2JsPQa
Va5batxHjsdl45c9fL6WvksuvaQ3NZF3Ll+5MpNOHCcB0bh1RX37Mzz1DgTEHHuH
urlxGuNzRpJH/8wjv3BdpdEZapOXqifhd0I+N+94qukgFaLa2GpgreqtH7XMxdpI
dRocnlQTMlgYqxJ0+Xa1LaAejZt0+6LyudHF1/3pgbn9WxF6yQsC8X2vyW929Jvi
fiS1XcByLidLxppK/Tw/7dgK2cHQ4Wi3wG3QvX1W6+ToWhsGB+X8Aqo9fIzHXv4u
cx488Bs58oM4+yDDt1Qf7QJWWf8c2MtzPncRbZWGwYTPe0Ea9DEONZtm7kxkzy5s
+QVdToWqZW0Ha5m8udWrJfvVF8MxygwS5LELjX7SvlfmuZ0TsKtkvbW9gwaScVi7
Q23QzPTJokDYOxfIr/tG3phCSb/+5EjRThW4IG+eFt1reh2dTZo+p9w5A7gN9L71
XDQ8sjlOacZCvl8UXKRApi6hRl2LVBJ4Ewk4NkrqR4w5908MBMpk0nBcbHBWuZgQ
836AoJsZan32GgPcCTT8Y5FkjnTFS7DdhLtmYuK5pvV/IxLVvH8ZCZTEDrScBohm
pjfVxvfmqFW/br77YGpfL4CfV2IaU0lHqZ2jNm8IeBF7noqEVy4Ay6BPRnghd56U
BzQgapsNbWRVscKM3CBzS9ioyrutwxDWN+ff979fT3CN5BKeAMGGDOlgU1nvyfc7
DvYt0nW30xyMOC7RpFIFFxQOcXbY50SgWEyNmua/jZlE4uEGAZty/JF9DiH3lpMJ
1Po7GU3S6hffEqZeGX6cOhBIDEhTQLLzrq9A5An1TTuq+nRcaMrPiv9NTT31Fsne
X2ZGkwVupPdkmUksGyP39rJe1QgWds5+EyojvuF8QcbXmOMQALgAWYQ34tzQBhKR
aeJ00njHX9GKGQ9AEwxVE2QFJywDjU0Rg5nP+wUSe4Hmt6bhcW7Byj9tTlsiV7rk
luaVymt1ujCX2IrbaSM1IcQVaW8+jTzkBLXlTQzE1iuxYE+xFpOwxG1yYcsJ8eHq
DstNaeIOW2ASaaW7dBN1+Ct+HIhyujV1Is7l0w+6pCbfEI0cf/JgaeXn5fzxG9Lp
Rvb2+p3vuAvVZnyNCfejYyz0K0rvEy8m66PFlCuyVkwbp9QjSGxtyKe5LbUTESZP
l1j/egk1WlkvAg2lbXswpA56NR5wpWm+GrskNf7Z+1/VXugbgmPMjv+0uSeQnSkJ
zcQxalq1LxBxs7oRJHW/YKnD9EY3evRU4W3G50Po9G5OTNdx30fFke47tpbqaJJa
772dIHjKTMW++U2uAqbzYBuikhZkom71tNMdI86NmPgiakk3gu0aTRx4RHbKJVX9
PjHf2UZcfoBkb8Hkr1c2BPf1ZBUPX2JOGd2XAnbjwfluBXhtzDyFetCEo+OVDu/J
pn3i01m2NAqrgDRCBQMD6YPMhmHlWY0b2iPRf7Nw6A4FVF1KU3MV7MXN/OorhUt4
8mK4Ig9xOcgs3AcCiNNNnMdxUG7ZTHjPdQD88O+CS2iBggx61U1QumySdHqq2iY9
FwptLnyPHmD/IMeQ6ommT0jO4H8YJlBx/omQR/ZA4Ci9gTKt5GYO7tz8/m45YYxj
9QyF4j1zPAn9RuR6oowKpfUgAuV2NIpPzM9+Wnkh/KGYztsmUrNFv3RoEssau9HR
5s/1y1+5Y9AQR7prTIois6sFPWr18+lNm1vAZbLkvGEscY9XvuXOV1shCXslJYSh
FHAQsR9+219K37D+TnTyxGqBspZ1ZCDvrVmA5e9ccrh154o8rTBfHvn+WXbrBmRn
82lhnOdTKV8gINUopVQCOu4ufUFM68P4DGvIBCAtzwa5tMIAJF/VvdW5ZoMcijjj
nfh2XXsQWSNGVaYde6aJ5Hs057KlGK45TnxheKpePHHje2b9lwQGb+gkqO7FfU54
d5wMzsBHEs7euNxs91/EY5PZp0JWkkdm3ecIySMNfnnQY0m8BhRnV7zzGKvN8Wfg
e81lvNVt1KKb1WfY2HIVbVzPBiUckpaB+srAl5+wvobWoIbUyn27hGPJMXWgJCVQ
Nr/OJtzv73oxzwtZifuTflBJk8gC+pLjkMVqTcDxc8p4bo83UrAcwb9aaVCl+b7m
E0e4mWRER5XWaIcQxw49B48+daimCcXmHWkT82VzBDfoNxLx9evfCzdKofjRF/pV
7kvK6JqJY1qu57IxdPoE9YeqqXSyLWhVotIZOKgIuR6Isj0xMvmijv7dJyYQjpV3
ItawQWF/0s5MaIdkBJalNV31MufC1kd8H6PtFtZwNCvgRZfRgiwedEc76jUjOY6V
0MMphGBhd1v4VfSqOUnkbFOOJX/D2mVfKbMqngEX2Uag8ORp7eiT7eQxDo6i4gwX
IV9k2V9/G+TQSInm6DXq1PvCnojUNmdXXLsC678Ijf00EW3MxIkkC9KsWEcN7AtH
xkFL0K8owi+vFS+TMnECO/rSG5upvleT03rpG/6ZW+2k4lzMjcpxNUB8XqIZUuvp
drmBPIqO2r3gKM6CYoU8uPbP+6H2i7Ddtfo6UZ4sGn4jcmPdhXHHWBSVo7wDDgbO
IZuOS7+IPrPD6eI4XjQyPrLM7YKnNhlHxmv3lq6HYdyjQ83AaCw9LAqdiXPF+l70
3eCB7d5WWWi6I9iHs3+2ItrKArgfjIH4GqI+OwWH59vDCGizmEjBGSrmPBbQMsrb
CkJqOuF6Of5IKO5fQm5RoC/Ue0ZEyhjXGwB9TbDFFCfexRhXtV5WU4sfVWQksaPa
8HayPbKhYTRqc9SJY7wlyktrA0i9l0B8OIHofEFW/6DOgUnMb/B0FP7RvKYk5MA9
xuvxCjhVqnKIxWrEEpUITGbBuvOqcAuQDNPeZM2ZubfHaQHpDlzHlrxWwLL9i9eE
1NM4gtkuY8ulTqJv1HsLPixgyagCfB3eO5Ku5LZJeKcxYAaPQHXe4Xu/JY/r1Sd4
3IjfYJeOgizy2riov0sS+m3cSjNVg8xuLRnUK0fjqrcQFA3WtWT9ogELiY7pt5No
BMvnzWNTO4vYXnCZDc4QpLnER+KXeAMex/0wWeA0mZX5oNws03yZImmkzXJ0o72D
zwrNmu38GqeTdjQy1FqqdI5wSZTrqleIJekkNJp/vus+q/ljWk5Al7ntELDMwzPb
wmchlNdV0TqBDqiN4h3lIfZn57WjtQjcunRC1yff1DOg97n10Sq8vNhtVclH4ElR
2f5R2Y2zlyhvfVCSBbEHGd/3vv7fTE/7oFfgMflxSmc4g9hZ7WIbGLki02EtjvYo
mLuGc/0pGto3L6uW+6b9q4+hRDHuaiD7BPDHaXlK+QN/BO772fzOyAK6hJRhv20c
0sxIrivFH2TmoNXUua9/mZH9oeU227la3504O30uqWtw5XQ4TB6FK8ErSp9HOwzH
MbCP2cTtIPMd3lYyhp7sQzQCTxVARnlaX76t6DZq0G2LDxJfIaTuS+RLRwnoZn2p
kgXJoROWfzIrsbZFMT3u8BM7P+se6TxLVwKwYZn/L1BwM9UiqgD/rw+VgFzxaQZd
FMucrZ1dYF0MyKmfmXGxibeUNE5PPEy3wrqgNbrw2kkl1cUb7Uo9srHD/CtLTDJ+
ID9bI3OCGGFUK3VumxuAL7JAnpDtmliXFzx/x4NFhiVvGoTckJggqCboAeSEPH9R
gyNh5dKrThnbEy1N6CuJJU+96NL9wlZ14zw/rWO+fidKR4kB6I2XdGgZwAHAcHw6
+MI6idGlZB3BqdUynPyktN3EqK8vD5WFEMubuvgUAjAqaCHjZg4W7deFbS722hqC
VXhz0Vn3hkdXpgrntRQo5Sgefh1k7AP8mv9JceVSRi5xomkHSQ+jhhBaOsaJWmkg
YgKQx5JqrRuJB4FT8dJcIwF/FenwiOCShvjH/Yg4GMEFrcQiB5zMfiBQ0XsJGoWe
nJFMcSQ1aOUBbaoJULi5uv77WhRmHXdk5ZAtoGjYyk2lywYKLqSthsaK6iZv+bXD
lAs9wHK6e0OEqyB2FnJew763d0gFcF1leqJTNV8LnsqMPZSQYtdsktpc3j2hLrkM
5LguU9GqgzwxW9QupEeidpjv3dfRikZDux4anS2bEDpnB3M5rMZTIu4Ow+b9xazs
Rz87Gyc/dr5yw+JA5NhSSqurIUv85KQHdzY2GoCzkHZTNymALEFul+lb5WGc4RWl
KGLmtGyGwIO4HFxtIBRPOXPcD2SVTQ/pdOMVY90F7ag1R28z2Ud99nrN7iW0f2aQ
qm2yeR9gnIVoYvH9oBX7d+2TkTmEOD6yAJfdFRAv36viU8P+ykwMWWeOFfJtWtkS
bSMQ1Lh2YAz2B8ShRwV63KM/+poPpv5OpfCo7Gvb2LRyBasSbj1F9rRH/dXDWS/N
KCvV1lAjqB9bNu+D4xcIszdTMhRJlnwHvYMk7Y/z2QevC8tauzPfJ7aMow8+uZWB
0saapAx0ZzkcGhCyovtevHMd65In04t6WfFYZcJ7N3qC3FC1c+6XlvPTJNPwckh2
T/NVuUxC2QvqiLn9hQHfZ3VBK/2cOVGSDJ4VzItlWtw5CDL3AGUR8bSzBgu3RO3B
lK3WM8fQB/D74kxGVhwLJZz8nLRSe6tIj7L4fn5iMWEdZP3WniW01djvnvD9Gl7u
FkqfpyAUGXMjOU08+0j/tuJCxCaKBnWJSoDygvivLlOUglqnKLaUUzjubVwtaz2f
fNTJ/fw4mtNGVb9vbhtrpQc5d6px6MjxEAtcEXBi/RU5biZqZRqEnBvVIw4jdLVe
y3sbcw+ZKxVSqeepoW7SZExMpK8usup9QFnpcpUvStrcvegLuaBuUMnxz7gEibtu
6P6hwl38lY5hlEN2NrRGgigNLrIEIDCMEftnm0Y9+TY8QqHKt4E4fBlqiPfhQbXF
4BNHrh6s6cqB4FBXD87BLKv784bShDZtlHBRvGYdJq5GkS6aAGVWFRNugwhNehfi
t6Qs69m7GestD+jDVSRL5U9BoQwVWUgmGLCNQ1eATKaUScBYh/L09Nl+OAaem6Ds
tcT0K7d8X8aI0pc/EJK6XlQ/+CuCdQijBayGoIdQVES4YYN3S05fhRPexKJu6gr/
WG+zmOhf5T++3vEvTs6ppJXSiTyKZ61aRPzGnmcWYJTR12DPrk+Y9JBIkq3OlrkX
qwttKerkwiI0rdZ1f4pRguGf5QV6FA9bFemAm6+MLQyOM7CQ+/KNB3eHXxhNUJJ2
e+Yvcdu1iC6dt1WOr0KYoHhO4YgMIHF03V7SY2FfKf6kl85tUFWGzTQVojVry98J
jKbLz2Wbk979yyVFWwLiNPtFOoQ85EO5SxrActYllse80MDqt1ixnDh6UTOIsO47
S4hv038OTdIYRmKUftVmu7T/Jt1iuHPNABVjUVl0Nd9PvFI3+906qcImIahoHWRs
fXnkYAz2SrPnMOjhO7oBZ1J5jLeIFWc/RXDzzZglTDX4GGL4Z2ipTd2cUhgXDhti
qZVyqSjykqELndgJRdg3IpaVDdbDnUEDUy3Qro1m5dmGjrqhMPyHXdoIVESvn8c2
T2piPCPJ4luVY+MfIxPFpzOvYPDZH7U3QJs+VNKmpDnk2KBYehCSPysjzXNHd8nb
2oy69WfHjoCgycpOQBk2AzUTD5H6lQvGReEoCDRtJsEZuRvabk6VHyz1VMFR4l5k
vVaM0GyYf2Hkx5oOFfzui8Tx9T4gkoQrn+yy1NKpPXmw3CyuU1ury4FsH0sQKRGy
y5Nu9hlpOCEMKz/ZoixvgdPSvVHJPmZgvK6wfJcAQ7Zq4oxH2rps+2EgZcZBpbed
Rp2h5J4QcASFxY4Lnb/W6kCYLhEpifNZQ42U5fT228BiczgZ7jKrKp9cpWpYkvvg
zVV1ZIXNAqyW95yiVcvN5MxB+g/yxWnps6J0oCO/94bOUjR45Y7jwtHMsiVAf4ow
PJUICq5HnW2sQDOOV3C2Oc/FPLER1WLwlScf5eOwmW0Q5G2cODycPzm1SmMGqDni
3umdJy8woBMnngW0ZkuHAaUiCsVDL3RnF1XRwLBywZgH0SVMPFNgB62eZ1IN1JNT
HPdxroXl5+wCRBsgm8xLktbGHgrOCGLq5lfyoaORNJk2Tl2AmElD4oKBPrP8OOk4
2IwniQqIv2D67Hy76SO6I6/YbLVxpZu9RCZc4Yp4JNk+GqSKQ+grDx3EUWyqrfJ+
ey6jDpDEV1AKUGaGHCKEA/fKRM4IAcod5MuFHKDo/HTVeVQHuXXo9kJjYVgo+QwS
laQGFQFZsKAPfCdb+BtZM8jXekJMsOSycfZGlN5N0eLXjYVkMv+x3uocHJn9Ysxu
NOseLJD6pw4b4EOKQ8x3HBzCjQPX8mqk5FvnmNblwd3uZsCafuRShmq3BRiXrPse
WcWaViMzkcD1gzqx3TZV8DRVOAg8jMi2Yx2ckylWqmL4pmQ0Btj82ndUH/OfEwHs
hzIIqcGqYMN9c2B4MRZ4KwoTLPS0ANav/oSLJFKKXTULCezZyBSV6WMb5htCT56c
hROo94+tvRE/rWvxJoHr5NDIn3nbc1IWo+PegsBxETdRX4E1nf8MyWDaRNPGaPQ8
Zs3e8e5nQWWGmkVOO5Ejr2t2QCHCgjndwQuOyJfTw5qk/BnbByxpT+biWYHqnnM3
tz12x8NGzz4y/nbJJ8R7s51q4vZwMM2qyaiMJ8rSA6wCAFif0i5ehyjgj4PduhhO
MvtP/S+bbl0ddS0aCBTccrsKzzJ3DBw3g02KepT2EaVIsuwqlXRn8Ag/B+xCaxcQ
hlojhRGt+ATgBnZ1NDIrBAvreosbI1NdALABGEbsCcmCWCLnM3cvSezFlOE0OvSp
qKiHVTRpjprsZwDW60tL6VdzmpinembvsIa0fcrhK/yX2n5ur4pdTYxEmyR/BSBe
iD8ouCpW8Uk8mYMBQGj97rIsr41kbPLoJ6Mkmq1k4JHfAnSV+LRSrmj42yS4jfqd
5K4Y+BoBhpLgB5rg8wkQUkxHKMKQ85PgM1iXsVwEoF2vfFSn1BekDuX0R256sPZD
T96843bYpHAMtyRIxiJ/wXS/IaiFQIzCfZGgOfEtc331lFWnRUlVLzGb0CZCoa5C
0kjGu1n1I0QtTny0jp1YE1kY5Q6ZyRx2uu2QOmdNnLYRJw1OkPU6SGkJ2stZov1Y
KZ1LQuBw5UwotceW3xiu30vSjKa4LEvlyTr9xQtgWtz283Xo75U2p85AC6Qo7/MY
VxCpNgv/FmMuw/zlfIbUnvrhcuucdiKlvs9F/oSa1J7aS56LcHy7ditVvoCofueJ
MisRaOcl8mzEHe1qUswTb4A5JnsVnQkqz5qv0Jkx9lkaPGrtyfe6yL4PuI9dLttW
m6RQ/QTB9SB1NV/R5y6Z1qN+TUkBBhDlJHVqCgKrz9712ks2rK/C4K54/j0FmbjT
0jyKBtzBJxtH7eApdEC4aeY31qhmesu5heI2bz35F2q6kDUU3utcv8660b/rd/M9
f4KiFTdW1CWkdjihO5LWEt13ecF12ZUPbOdslTF8tjz0dAXWqJD9/8tzbSQVQ35E
RI4uu/0QYUiUQvPoww5q2vjr6zAz5MBoH4CcwisDmjkIFBsJZu6caFm8D5tWFxnU
G4yOkesFk/HihmHb85tKTBpWZtE/pXwUaTOpEjjFaMavN4e83WnWvhj6wV4twwsS
eRuT5UAcsRsDheYWRUlIbCb4Y53xl32EWYvctCS1lq+G9wLm5wMZNKVq9lcsVY1l
`pragma protect end_protected
