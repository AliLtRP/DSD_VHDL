// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:29 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
jnGJXfS3TpKas+EwojzqQ3z2ycVHC5t/6qT8Th2AdeFvgu9jnP1IjMvKX2nN4YCM
on/XfxpgF/PAzZTriUdxYUZYRntTsVM6gLinwW7lreP/k6WiSKDy00vuAsazsl6W
jOQf7Ifffi4vCjIyNEyoAzflrBWXKJSfJHNo7qdnQJg=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 18656)
0qJ3yupK47m7Off82h9tPE2GFasdSONNOGSFviWRoiK7JGg2h0cJ+8hmkRR9zU2F
V2N0rhqYxCQ7ABsp1ruh5GQ6kXCAvSHiAmWa28JA9a5Xd1K/mjxecWIINTmRPmNO
8t0UDyrC8VTky4nWAewG70XV6s1y6JOKucU23EabNpjJHZnt4tk+/pQIxBrZYUyz
UeSHjGzqcGL5LEyS8TL1Ew1T464SoT5Trfgpf1wl6WBbZCUXCONsh0x/UofrhcDz
nogB8grmFjHSMdx9AGeRwDFlWVk3TbKPRgUW6nyu5qbCH4aVbwit2daguImij5G6
vjUkD/8eoyhAkxI8JJ/FAAilVYWL4cUnc7Gy+JzCAGBl7QTZcMOgOnAb/n3/7XTd
uWkUlNGd9CvxwAF9h+aLuenfzDLv8B3/dyUKAm9wm2V6xUxB4fifwgBY5MTvNp4D
5OnA3h8RwxEyFFAss9ix+mIbtz++NCgL1uhwhWmLQ7RzaeIkVtiOAU6+e/jToiKj
7kum6yJpYX76dPa8nlF+j0DjVw2bhdrk8tuXhCRBZ4ZkmsHPomgT9IXfJBC/qUCY
zSyFOyF2MBwEQGBNSib2cVs498j5s7fpbU4OpMnIBLsFLZM8/TtTHaV9b9CDC4OG
5omHGNUFgFP/UJ5ZZWHG2HTJasXDtgTp8O1lVdPIB6T71capCIWRecw8FAnqzk60
v77rBR6P9b3hbFTrAvh5jcuuu5Zxnn2wurnOd8xAFK5zIIl6TBJXCn9SgyQbS/ap
ilUNX8hceVnLUiN855V/IkbDZXw8ffeMzV+b6ThhZYmSvsUfi5dSsey2BVhwbbG7
UQQbm1Ja4bUG3MsoKitOvSlHqez/Qg1MGleYlpatI5irbsfcAAwKoRIF+RQOV/97
921yF7pG5QpiXleUemaI/a9Y2SieCxFpQTDGjpMtTAInJPaHPPH339Z778E0XwyC
9eQQe8KWzW/0Fr8+yn96xVSWjiBpBREjw+Fpuk+wA824YTvm5W51kH0kqkxH8X4i
wTFFMdvDnR7vgukb42Af4sICL7F2CYmx78fm2bgxRbvgKoELEhhktaBZGUBgXduv
R0yFBwbBKgJGMDRgM7I+u3qeVdWl7FQoatBl9sAhP+B8DTe/13Q85EwZv7qcb6AL
ouRuX09QpT05IxSQw6wsvzZ8MXTz11Ja+NG4trh42XiLK874ef6F1R8DzvkQ96RM
6P5OBDI7P+UvEua8OtPtJXCmBoU56XdB6rp+k9F1wwg5oFxj2oJz5/CddkMYTbVc
6qewON3cCgSEensKstuOMXJC8g/bijXDEezI3uZ24dzatxb4/MGq2Q89q4xxVkoN
Q3pNYJPbjWu4q4HZbthBH0J5UIerCDd/1ssVV8Ra0BBpAjFSzfv1ytQGK2s1FnkE
MxlHNbKQIt2HwHaUHDPZfYAmp6h/pYXGGuBUD6WLN1iXxCOKxcp67CQtPwWsjW6E
6DE4hNWxCqrM3zKWT+GyEf4BoFDQ6+unwL8/zBlX80DjraVtq+EcVlLsQ711bFFY
4+Gmudsre6shu7kiL+5T08bdFBsQPHbl4pvs5S+w7gSryFRUel1m8muHLtdVW9YW
kmpmJUe2unzE/Wt2b8xqSyXyAwiZw3yiKceVtJ9xpYDFSYtCKUh4l5Q+tCrUQUDi
3BAeh3tBEmOu/5bh4Y92EjQu1Ph8VoHdB1f+pE2T0DsqeQykC4jnSp7p5t/J50pe
utBTJXCv4btVq1WTUGmFdRKqfU8MCmZB0uePuiwO54MekO3PnVssO9tU39a+yO23
Mxmy01FCv+b/xQ7B6Oela6vskLHc6eGmXz+YLun7cvfNM1P/+AeXOK71DQ5d3uVX
qCw/ePNfUqMZsmWLk/MVfIcNZU/OA1FaPkeYjF//8CPrk/zTy+kHU1NYAKeJPENu
bRv/rvW1QtyYHOsurqK7gkawiY7SvzsqXO9j66zrnTccpZYvRwT/6TDqT7XaUFEN
jdpVxQIpCIk5c3xRhf237w9mpb2bZR9v7MZstYBXrkSw1GAQo/WceDJXqUvt46Kn
cV0LVuLIe1mdImJ+yxXIDHYD4L/vbeXru+jm4r2H290tdqeIJZ+6AaHTfFu0MD2e
TIZL6Aadm/kDU6YDMUstX/8hP1LhjxTbOwDKbSYV5G6C9iOaGkAaFJmUtfSD7+iz
EuaDcO30DgIAn/HGiVyDVBz0Yui4A7++Io55tYuNvIqqeRvZM73PNydhrYE3Vp2s
KfG0PJ150w7lmFNFN6A92nwewsuhC6qKmyIGxygzbX3BBgzFhE3+BeFD4kZgOTlD
WP9E3SS8B61fiNRd9WOwfI53LM1pOrcc5u9SekpVSzyfLLZn6MW6uNoA+OfV3gm9
qFhu2oYeVwE3KswO1VL3sVfHttK8v3jtwaoNHs7sKiVa6vRV6FidEhba5nwRLqOz
BzuKjGKzO8p4I+XWeEXonGpkDiM3ffKDcIhZgDbqCn4jjWT+kvhaH+aMqKF1glj2
3YSqIWSbcWCuTWH6ra+WoKwrUKjQOt6gXRLZEg/lp8eFWUzZdPSTpo1O2W6JMwjo
BjyOcoAv19a7LYffsYwS3lbfQSO8wgwr7JWd10wxW7NgKS2XHmAX3FMt3OgdAttM
5T/dFmrlj3zMsad1NmAJrUEYLNmGLbz5dzLg1uXhPl+JOshIwoq+HHSD+WipfNU4
fPJsHvLIEYDIjqyYOzowRL2g+VDoJDWA/KFFXJSvdtjhcVgCV6KsSmulRmqDDu1v
g/SFC8+JaLbRe5dIRXOagT56/kS/e83YfZ35/uovuqQWiZpJYNENWRb2P7jE7Af/
ZEPwpSBLNTLphWkXQ9SgpXH14oV1FoOto2Qyzv4kZ4s8OORYSvU27w5DKksA89n/
+S3dkQX7So67LGitqoOEiIVwj2KU6l8e7ubxfSEIulXReVbc2gtdFRmE83cC7BK9
FnPRdizncYfJIf1jtgjZEgYvgYL9AwBWGLiB/GCsDRey1VIbYY8Fmjp+MT8sWMcc
T/LEK2bGDdgCmUBzlVLoBcJHUE+EZhksZOlsC+/0R61RmFhJRExD9EWMLRqcmWER
kOGGp7sL+yGFuIRJfasSZAy4ntQpdDrEG26w4OEjUpdBTvxlr9T7PkqHIYuNpht+
ZyqqPKn0yEzvqUlTE0l9vp/UkZz3Zs02g3nppXHSY8H7XQ8jzwnGk2juwOt9pa5U
UEFU5gpUdeN3Ng3PDfy+phk+NNUjGOevX6xvSr7TEqnJSfTX/OXwEasaoLXiEvFw
3kuNjV/VZwRFB29DpgCxM3taOvrXSavWOHIUcWyYVUrZBonllo522fl6vdU9XDKa
9bF9ZybUUg3y0zT983rnY4AswX1NbQjoBiNl8r9Njsgb4ZUjGUkwoJCI0/Y3MfOG
bcubo3NVXIr+JYP0loKs2BJDw4epmZsFj96F+WlgcsdFt7Ycyy/QZE9ASNpGNT7o
3aX/vrfL+cNat3tEgK0gFky49/2AAwNcsDjpACAw87274kRxoSH+1T3THNvDRrxY
5v3Q/5+zBFH7ujpHXi+tSQTZQJTin8+nX4x3GDx2WQgcl6UPqzZMnG+Kd8gw1xO0
jk1/OdOUjAwUz03fHrI793DY7yxkrBBp/KUiCZqrEWDRZZCX6KbVQZlGV3j2yMaM
MrTodLqqCd1VqfF9oEmMJK6otKp6n9tGwwf1KqHUG33n0oMUoPMYaWchRHaEvKgX
3+tJDVLYEDi5dQltnJrSxN2Oq/DEQ0TGNLvDgGAGvTHoTBlvfwiDvJJX/aniGKO/
9VEv3dYaF4hu6zb+q91w4lLFTrfXGW8JFKkCYvWf+9fFtRF1D060OLaRG3LoPFJy
SxFSS3Yyg1PUOjQb0cQVdVHyD+bxcAafeuAQ+3LbawGrs1sXcbiekr8+t238o3rm
H9DDwcv1f47CemNlLVAMXX2JOFDfIVgLsGaULEXZEec+t1bXRFpkXs53nbUJ5ruZ
zX71PmXq/1WTia4hpUtTmgGFh1xg7S8hsCaIdYbyU5gDKrkcs70BtOQYTojOgRKn
q0eDogeJhH1t2Pjs2w/nBlP6/aE7dI9OuPhELhPApOaQDqY18UJzKArHB5v85eCl
9v78q4WHAPOYZkU5cy6iDhJzAw+lPl13R3LvqBnttsdB5Tc+pyBf23uU2MOn2PPu
1BdpsXqCpJLChlPECjnqyJYbMjBlNS4pIIjlmMRcmHVaSgNiDFsouWRZLZdK5mOS
1pMR3QQHv4CTNbJ3hypOZn6PnYQ70o+yg+svOy8WRlToBef3rTly5S1Nzln1ITXT
OWJuLFnbksaAEcMgHEb8N6hSCKWCg3NLxNX3Nbr1EXyKk13sB4KazCGO0zeEN1eC
uV50iv6JkoEJpkdvLxjA0VKYQAHNvtZjy1clWpfecZ6Jn/DzQbyMfme81PlTe0pC
SiDKmNrmUlIn0DS8YbFpIVgMt/72UwWvuT9sHgMXxhnexx/jayv+P9ep6uNKv6yw
kx3GL/lST6r+gxb0e/nzR5TGGD2X4gZRx+OBi7co+o5a2XVHurMeKvKc+nYdoPk5
ddhpvI8CrExGK+DwGcaO5znP58dw05g0OMgT4d5AtI+cNIZpNwE7I/7IJPh1V9Fk
+MWZOOucrb4ppqfX1OE6kUQL9Sr3/V2KYDp/yLqqESmNh+gFzue3amArXA2AE6R1
hyaZUfaLLdMOqK0VYOF73HCgYxsNjt4N/NohqzlfxcvAaYBe7Mwj34uK2xaXYOxC
vFh7ss0OZ4FQ2zjznMF7HiPF5jLep4VuMr4Zfdt+8H3iNsDTGf1iRR2V14dEDCxR
zruT8ieWwVyzM6r2/uLcX8hxk1nRB5P8rEz1THN9jnMVNxmVJGEUDzE99fJk/8AT
m4aujCDiJ6vydAfLF9E90djaqzciAFNU6VVQFS6aKJNW+Tdx81g74au/oIxpCH2e
XssDZq0KW0zvVBWeemLNehXALGrZYWzQgLG5eck4/tNMJs2jJe01PKhaKmCqOvBD
1g5LDVNh+HFQzII/HwjsRiMUj6I7j4tfwOGYqchsJHeJBak8V4gFYJfbVOWJflgJ
InXTbdwnYVd1Ry6b5GxSxcuMwmEjNQvcriRAprIjDAffy7UryxFiiQW/UkpKRvUZ
cNNB3Pg6n5lDLYW8sKs3qfMWYkfsQVbT3ZzhJZS1nuS5zSbMmYS2Edur+brGKAc7
+5ZqtLnbx0ON4VXiIG5UBD2GzI7tvMmvxdl+vUbz4+UIO/SmSQJU/riqUNFFR7QZ
fe75O0XH5cbL3oMDg+/TyzfkvFqa6PzUuRZc+GxKnXuq4jB2bNjun5wOBKXoq76H
rMGfBByNH2SKiHX5slU6ltADlKya0whxTmQgUZmdi4LqZNj7SEu4ZEFPPlFtSWOb
8kkLV8Ucy+bGZ1By5MF5cMb9k87yE1UgifErYk9ZxBL8avvpdAonpeML5rV2Fby7
okQZP9YGegxpJTjc1uPhwzeywsmvEXPtnMYLjq2rbHv6kgn2rGXeZDv0/APxYy4m
m9qLXWmmyONx9CVd2CNNaev4vkeCyD2U9hNTYZi3kvLl6ItqGTyeaXa02286FoJQ
/Df/8jH9/cg53nFy228dHME+RTAmjf0Jv1cExX5lnM0dgKbkPm3BJqvXFZ2ATEP5
K56OLFJJRQCohkBhjD+dBRkoPCVIWBHA5zWtwSj5XIlzREkewMkd4h1Qw8RQ1uEb
yb2+nFkcverufrmDPJjWpL+odza9aprob7ijPGWxTof2oOKnnDhWoVWcNpjfAnP9
FB36iSUzeVW8EkJWjPxh8TENFHUK6NHov8eErOmf+TghD8rbUuZFFo+h74KaS8XR
5LimvvxYAMohT5A/qDhPM1+K+0BrLMGk/9O4p3zj+IWPgbCTNu7Gbch2aDEiD9mF
7HQHTyCji+65ObBNOnm2sl+rdaXtfsga3hOrCrw5RfW836cRlEFNqtxOcOc4h37v
zKDkKRDkZQMfWaXyd2f6V9sO12gED8C8GC3EKZbCm6m54zpRGDToiCzov0/GPd6y
Gr2wceXTkcc8RNl3llD7UF15AFgrsCY3IxnZG/4Qd9vyBORqAyvfEwlt+Lj+3qNY
VIHmhRCRlDsGGAEd7V52u6C0z5roohRlGfIfpIG9P7UR08wD6ClObFkrlUTlYX6c
Qrbn32I9FjCzaDgFW1C9N6AGbq4uhM8buYyfo15IuhmCmcMfOnxOzlosjnTlAaRC
RzGJFrZo00/Jo/GhzJRE+dmt7nbaXEWiNRSD+XRtCk3+O6J3QiLXa+iNMHtG5l6Z
yCzV1xXqUHbNHWMT9AaNSZt6BB8l7EazkPURRLXGuiUV1qzLYsYVSPsqOcsF5Pwt
3ydiJsHeyawdhOlLBeFDC5xhQIHfEcPDTid1wnPqwl4KodF4QRvAjo9peX9tT0KP
S9vU6vHLw+y1yZ4A+qqlHOk1f8RqbhfuycxE2J0P2LZ+aNcD7cm1t4jMmHMd0NFK
hYi1qBOs5tCdqypfj3km2s4KYIj5ahq1s0bPXPQzqS+rAoOmbnYpynGW+WVvK5+y
mCZmQqtvl+rvOsrKhZzNd/l67/CY59m95u4Hh+nKDyLX68gUxSGN1DAZrKUvTXf6
ehtQBf1QIHnG7N8NGWzxHD4USx0Yvgbz9MTCIAicP0NNiw5gj12Xzv8qpl6426Kl
vcu23V/qresVd+36fSsE+W16uJ/T6gIBWvTuD0ZY0KSV5gkQm9BSMXkxKDRJxYH2
V9LhSQaCbvxhgTWGac+SjAKFfTdt4TmxohS1RiVDCQoMHZgIpfH6MZuJqluzaPdr
Rg7Kg4bbKAUC259HwRYwyXk/ALdGugp4of1svMy+j5i/qk/L57xH9Ps8mge7p7ZO
bgdQAsCHnehgmZ3ZZxXeei4qLbl4lv6z7V88HaTN7VE0e0dBkG1JGm5rG+zeji6Y
DBZ/uDJLD1rLVz49Ou14+okKJ5eCahiAcYKUwzesahJbfPDss06K6b9tArC//++8
QLHjQRrWM9mZtyS/DgQUinGqtGOMjHs2S53kRbb+zYcejzNM4/F9H/FaD5e2nZNN
XO4GowRYs23cb17fVNYyi0J70cFgIFGpUPdUcJRJRHELZHaRLNh7dAqC1XmmC9Jo
T4kt1/seYbPofY64h7xpHpinErVWBh+2WZ8ITyXD6jfiU3kSgy5wDtNaHvbDJB7s
rivPl5P5Nr7vwYbqPPP66zuUDfGfcIquLQbEyO8/DMYc40/+M9vXWpH3G9FUXDOp
wIRmYSPMR+QVtmd7p2zbio1hkgszicn9U35KEaH36F5EF5LvF7TEkrWVKZ/29rkL
I0UXYfo+41khUZrG1Rqy56xQS28Gbs0/pIvJQNHQ6Fz0PhjHyATFLBJeWFX1tfUx
KI/HshnmXAxko7sYNV6KPXjg34Fae1IUJONJ1XbYTPhvZNva9i+Q4XeL+C2rxRQZ
Ljcv19vPF/8caj/y+GJf24+PTuXrzr1rwk4T/9Y9KUSk3WgoqC6tkymmKez6XhA4
Mi7M3WF+1sbrPeht/OLnwmeIHvGn5/w2dNzGmWyYJkICmxvs8v9ZYRv8dSxpIgpx
5tN2oFezfbrRFA/cPmPY43AK0FD5jHSSCeSiGM2rBjK14AxhlmqPV0LUIpQd096H
hCcx/Sp4OMDwoyXlY3t+PPalpUB3Gq5/A2a7yd4nFRcWlXAKqtT71Gtccl90pZ7k
CTJQk89AIMirQE8qsjiBJyAMX5PeDHlGSEhtXR3W8zknUBQ6sjwy6+nxJyf6oYm7
tuCpkGQvWytljejx54nUaPZokNTr7SFMkO7CwoBHpg5c7t1XdDGkNJM2WIChdYxv
x/c6kQBGd/pAmmETKeO9xIt+XykNO1kOiosw942V+Yq+ctw4APZUvYEhtnp7QMbr
OVtx64JUI0G+ueO+kyU/uOyfRr/0lZwnPPZetuDuAovP5kAKCnc+sm/yCLBLphZ4
UeLuePjg6p/U3lmHz1xdAL1hHHZpISaLoM5lj7oY4TYCtv7RisrG3dXEW91QHdUS
CMqoKB6flfkQtls50j0Bnmp9AzifXvO4iiv8/xJFMqAJBjTWD4Nm3Jzr9w5fWjnG
FI8tZiQjwKSrEMoxN8WjZpSrt3lCeQVDOTBLVwhflA5EdLYInLFgTPGHaNjqTTth
0o3qFBCN4RgJ+eSTGH53qPugJxveSb7FB2ndwQI6GljUuY3mUVL+I206gwv8E1QC
ZNt1nFXAIW9xwmoigHnW/dtAHRj70/G4vkKB4FHPPXCXr1jDqAnl4LHM+Zj0sfFn
bnPwDgJYOoQ6Qz4ALfWJRTExd6gQBcmibDdPS0qIgw74HvNNsVd/Z0JFekZK4THA
p02Jp82cQM4sEj8qQuMDm78BzogKiUQG7aNnav/N7Tccw4YeGD8YeNcblQQlfzBc
glx6M8OKG44XnjnciNwNqUXNKCohM0jfrFuYXKNg+n2w70KpLGl4sZP5qlUWGJQx
2j41kINa8Q+ZDKb4fU4lY4ysBNumiNNbmbWhnKtRhV2vD6iLDrjkMslkvq8ZqOtn
8RNQOhcolNzU99dJs1pgZUN3nq3LlYFbjnk0Dhy2PML/6VXgc7NM1kJl6wzrQaCY
pFPLHsY4gTerFTLHGhh6ZRJsQcZ8h8Giaix9+rP/k59BdhvlV2ItFKTaebcck0gM
yiUajNgcXy0HN9AtkKoPNMvnRfb2RX98VP6/JaVRL+8S/aMq/q/rYkNRm1NFUfq1
9pld0ZiC1Kd4/0ATjmUOBVFr0X+BRdRDCHSlZeBIO/18wUVdwV9krhLfUv1ZWwuO
vwF3iHCAc1f/hXkyLN86Azr448YeJI6NaVUaE4a7NmZ+HOKfE1bQjek6n51ejvlM
VFbSFWiHEZYFSu7Gb+fsX8M9MLBtlmehNinaNRxvti7r7XFHZr2s62c5brt/mBuF
7WSZacaOu3W+3n8KbYR4qAsZsuUzSF6AjfvndsfotwTKO9Z5H9YYe63rtKEJS8Gi
+Ij3gQYYgZdSc9CXpMRIxDUtrLzvG2ZhDozVxnm9JyVjxXsypddtUoBVTiaNpKa2
rV3BTa2U15sF95rXQusqXotHnGuFisYca3iynA+fGhIe9KVTT5B+NwGEqRkB6K+W
ZbNLma/Jfj+vtGg0iyCOHH0BsG5SsWK7Z2tCYn4H+4keO95pXMrTVgnSE8gHU5LS
4UNjxL9sap/7ajE7JMbwtrHXw2oJKaa8i4Wb1WlLe6gK8i57aunGjZDAad8jdI94
A0dndNOcT1qvQ6maiqcHgLQ+A393q7u0eu7+ROXddYA6icTfttdxKU22YOVdLScY
0aqf84YzB2hLsL0bs5vCTkFcBz/unMKMsj1WtLMPEhoCXstFn0nXzVCCt8heCOtL
nX2JzHoHesEvAPJaf5mnDdh+EYADQl6RtO0/hxgeUZUXeH9FSCNqDEysA86V1aG3
GHMOc63Aa9hImLaLcsRRmJls1kCsIkCVA4j4qe6hK0hYRaOhxGyAWGjjy4zDaVqT
2Z1K0bQ/ehlm3+iv+YGZRNBaF56LCV+gH/ogSUVht8mDlOKy/iG9a3ztsRFU9AKf
GVUFD+m4NozfWc13qm4/sW2luOVfrlbj25cRSKSR1wR8m6Tuuq6u0XG03+dGeQf6
1lEjs8lLIQwEvQi4YSgtNAlK1BEIdwjebB0zNsAXhuqHCYucPr7uXyTZGw4X0Wws
m9rd8YUWUpKTLI7BfFJRGE30FzGmL7p1bRl7L+hzdRr2rAgC6Y07/g/sgD7c9nlU
7rkPlgeCV6BZhVFVlIlE0eiP0eQTVNQkqhCr6T6rO2Vx4DsCgdo7hHyJ+GretuUo
PqaFvIYlNIxxKaZ88ioA8bF23E6c1k2z+BuFbo9X9a4CH8h228gZrKiqdgW7//BR
9DGgFJKl7W0CubDyURWly05WjEdVYHWEJtW2CD3muEGzJ3Dzr8m9PbCsb6dDGhSC
UAX9BtD/tpeOIOMYUGIrkUpfhUlgTm0mlyt7RI+Cfd3IwxHIiXW2EtpXjmlnwkVI
+QIIzUvwGwaJkGWVI7c/ac7m1OQPptqog6qID1Tf1zfvKgBUQZWTx02tM6uRjLEK
D+FrT0UnRlCFKW1+M0qKuKDDmL/RRWJNhK2exh/3J1yTV9t2I8dbSljezRGOp5Kt
Qv4EMeIBwqn34ZtkCxcX2Hsu2WIyrGfOlbOW1x2fIVP1XPBJUHwdXDzIe8VaaY1Z
RhRwFNrmZjKvd+ndJywmFD74W54aqhOuigieLKNgbqndHsLpz+Qw8Y811tDavkZ1
kCRQlFDAaBUOnaRa6JzDT9pNDz1pTdcgtx5/jJ24xbzYBXANCNSwCpDck+Gbjrkc
jRme9ycw+CxYasGt/ZZ3i3TbdyEkRmiBGZshR0WFUGLqq34zgGEbW6PBGns2GeWx
QdzRV170GXXA1Pmv1lxeT3A6kLawTpEcRd+GRbvtHQVXcDimidAtriUnBsBy2Zx0
G9qyEbejM4yPLiy+Kvqj0kH0QYyxGc5czBWXzjIREG3CE1CatldNQI9ZEYyDwLo/
BbiUeQQ0DSW0ZEj4fUQycxw0xsgmuDiC1KR4rTUgTsnx8P6cTIu1TJPA4qPqDOP3
wsZQ0cnbu516bH/QyI3fbwWtvEgGX+Dotl2LdIJYvei0qLZJm7P1Aj2ewdtQ1iH7
f2c9zWQPNJePcLxzLlw4ZYgfpy0//Oyag3L6AAH1ZA/wYdX6exoUZqDZYO8dSmLe
bGEol0Kz/ed0dL0XRG3165xRj+VnC5Dzvjhv53C+NvGeG73i1rJbJnujCtso0YoS
LbZQh3R/zL7oEZBzl6fMbg46O5FcDhD9TKMnSbismyv/YbHbU0n0PMKaPgfkyt9/
rh0fTY42AombBfeSdRYSmsqJdosLd/182edV0xsMOb+mECsEfGD62mMDsMRYuC8+
39X/bGUf/g+WBxN2NjA6oCFmZ3Tr05mB9N9l5YxBT6WzFqniIVFgNbgCCX28mjUb
kIaOUsKeAU18MHbgmaFAStDd3sMKZRylGaLILkpECdDpN/HtyNJLSJn7vAEkqrmC
4tgwtVa92D2xtPnv0Falzq8rQD/l1763bgoVC7yb18O2rW6c8PASqu5k66eIHStz
eiXz3RpY96Pg+SmIdiFhqh+bXml/i0Mg2VC6IArfdCF92jHh/idHHTguJX/ey5it
8PI8i+eGokwe+jbGKR6LrVMEaAMbPGaFyot5Ext5TBO7lEQhI/n0SrL2dCFK+0dS
eRwJsKqXTRkhGwc7BQ+dRdPabIMi50DMV870jyLNKHMbg5sDFNlKp1oXGEYJekVS
v5gykZvZmA3vRSHNiqB4X70he2TYV0rJoy84fYahqeGE0YQu7x4GxbCY5bCE+++D
LqHnZlcLLY+3DswFoE/xY+m7qLxZ6U5O69eVi1I/9Cn/u59Hx7eNRqtulj3jDU9G
84Rnh22Hp7UwgxXMHaiMU7cy2N9ViV8x+4rQZr1/J3k0mEXX5Re4iB6yk08t63Mc
H7rPMdLX4Ra8BQRJFc7dF2I5PKRqZ6Uq4Ap4Sw4ltCqpeaEIMOHtDkDWIQq8JdPx
69+jkjG7wxzT5fQfEdkQ5J0d30iAUG3QDwBl4X51cgDDvB/MF7FiOm46IV5LZTSC
koS+bL19zMfp464eEk5M7iFk1fMCShlTQHUrYdOufQqfEnstIPdJT5mtXy0PENeC
m3gpzaPYjc3PzgRA0LeEPoAwwTsTtMOkI+hPlDpeKXVXh2FlhB0hzmefQnpDGjCy
hvMIwjn3l86jc78zj4LIV5RpbYt3pjth9AMswf3j0l+JY41f9cae9w2jZNYegEWq
RHlkeDJi9XLuxJY4I/KH0nWfOm2KSuNxVsMCYmnNLVcEvdX1P0bGrLJEu/Yh3fpM
icvDUErEGNKrqsk5pLr1xcTQ/paxpBhWa16+ufKF60IEA0ZC5snnAd1uECyUeK5R
xxzjyja/of3MCN7muyo/0pthtZFTMibyuZjPdQx+sQFexzBIm8OQhVXd0gFH3wKk
tPIxLMZmdAJYf8K1XaAo2GCvnp38o0PBSSO8UQTwtBYcqXBo+nnlyYkR6nxCtvc4
WmxbPmUB2erm8EjezBWw7cAuKRGeIBeEAguCuzi5xKoSLGniCdRBONhsAZjz9Ntt
Z/N9+BaJTNduYKGtZAowSWasFG0mis1x/OhlZJRMwYnNIqV2QVLTBoZ3SUlpxinq
oBovEdxPGYMVJwaBg+Wxgy1v2mGpiE0fTGH2uf9kOe6Y+L2Y5vmBMNqQX0NGoTvP
v3AU3n/v4nE38wCX02yBU+DJidb8TnljHuJAXsarEQPuFPuhK+JCh+MsIHqoOMhD
N/cJ3RXHFInCkafyoE3dO0kUOz8Lg41CQGVITmzeFkMK4MfBc9F8o1EvCR800yjz
ZmBqsDaaKDIlQfcLBWgDhr+BxqyGW3thL0X0/wCz4pZyW/6X5GHg1ETFkFAaMevI
4b/x6WQ4UaT7PQG/dokekwLEFmlXXQsgolOIEh2qnNfAqJXTLsrQ9yVjhR6gqovD
N7fgGdE3hCkCP0asn1aRCHi67gK1BngvGvQqv667qiyqjZrCbhx83Kt8+xqv2lt+
wD4Sz8x2g8nEaBppcxn9LVgLf2EDFwdVhK6jKOQjgyvKFVkNxVUgtFluMdgZjS3x
6d3fBEgoKxegTjTt1v/rywq5Hry1KNd64fDX4Tdm/wIMMQlKYzMYstHulv7U8M+M
fzhUhZ9fU7Jzh7Pt4DxdKPnEYM3lyubEyqE211DTdJWejGqX3JgjvQZXMppWsbJq
k5rKjoD2KRXlQuIyAOv6MfquVz/Rrwcx96LTXQFenmQLur3zf1yZPa9KtRp5PPp5
2VzLqxosIrh8TqHEfeJwmlZNf8gi4upTadRr+0fEbCrxrFjMjVLrN+fG8iHFofcs
o2V4WqUcHdT4MR/ykJRYbtEsCb8tpFAN9Y5VmluzQA0ArsA+tjhKd3DmNy5UJoFX
lCAZwfRrN6CPh4WxQLcPSQli0jlZXS/Fvq4Fsf/G9/r6RvOpnCI2ZTo9ZfyChwwP
FROJEdmC1UiNQgbFk7TYSSyEcrCel6rafDX5CAIIcViuIHPtpOTSqrOgaQmpLZ7P
ObMxwhTU6YYUX5xgsyQfxRcODTPx/kvhwaxQsewr80dxWbbxnw6OXeClqc8KapSF
eG/TjopwbIWPzjgkZo8dj9nn5JSzaa2Btpl9gd3dkHdBSLIZeFd/86Zsvf/OqxM7
ZRuyuGG7RUZ8+p3qQaKzymzcizKFCsr0R8qUlgcILmhpFZO2mKS6xKXdkDa4gACy
RrG7mDjfz5XaJYWRJam2mwhoWHa2u57g4dkRYy3XU/dkhVz6rKC+nyZvDybcIoFB
M1WpDWepXyy7zfJurPTwiDbzQnjRMsX2ipU62Rqewwi6PjPdz06quZgcp6jzC/Th
UZNUZmIM6FKxSuXxq1UhzwXOTgiIvY8v8vwyQxTgcl9CkStcKXTmJdnJNokjWLVV
IzrczoiMXnZG/byVvZtt0jpqn+2zhAyZYqDdRm9PrG2LLM0X3krDiMjVvZKe5U8c
m2fQGz/dK1+UMsFzYLl994aocFwH7IbGJVsVCGW1xQ70HDLUOfqe/8WTDS6rFDOU
+K1RQpoIkqmKytNCQV5E8b24HJIOepGklznGCqow+UrOEYxY47bKgCspDO+9PK/9
q8YUfDe1HCgq4qITc/xVehhQcZM9E+fkSecUxCMfEyQUhzdwrVey6PpUGz0l1/7J
bSn3zT9Juk4w85IIqkSr1WZ/9h5Wauq6I8HmyRpHVSVvJLYrjLktdPRkbqptYQRi
BnDU2hb4CyvHoenP7BL07vkN3NTdnndAT8uCNQKmAofrBsUytWS8TieoEEgnzO+p
x/lp+cmHLF8vGoNulMnJN09eka//YGUUsxb2dZIfuuyUiv5osNh4sr903GeJHJdm
D+q6F24CRjO/ftytX+UEr9PNUnTdtPzl/vhfe4IxKhdz/pU8/M5zS+q5FyN4Uz8C
jr7vKlPEfYsHz4lQs5hiLN4UJ3dEiNgikBNquwPy0828uVUYoZx9KBBHYI7zSnX1
v+WcftJA0iiV9vT0Knwg0hRMqMhpipWbYiSpfUlcX0Nwn98WSCgApAN5E8zNpUFl
TYVs26WdCvu1oOSJS4fff04kRaysvPaTDDVPrLsRSy+jag4/JoPyqD3eKJBL6CAa
Gi5in8lhEFGjmMh4PLyx8XeSFTCJioB43nJPB/JKLVlbmHpVbkjMClCykSHSqqXY
kmVVdf25xZm5W19gHqB5mm4tL/I/c+j+e6yKYki5FX+R1XT7lmJS8sSaL4Xls+mG
QExoYJ41kGGcetpugjGXRHxSIEqARUKcWcxlIIAF/6ZuDEReDFVRoOTW4hptpRLb
kYnLzx9U/asGoMZtAGKtxaH2tUaorun8kS0BY1PS0dc0X3MCddwAyXpSFzP2qSPM
14K7EkO+87X5qAner3BfM4PYu04MHcDzkvmHYM5oTzZhVydhYT2WU0RXWUI6+29J
hU7UHMIp/SphCagrNtomiQhPUm0MhmXdxj1HTURJP25CEM052iLA00cwJ2k/mKZn
OdMQHV+HYdaxYtIXEjrfy/ZfolLx3j3k98HlioUxPG6NKWCsiMEhbi4Bv9OvlE8d
haXhcqhhRKrO9DANH04U7s4okIX+n1JUedyXDR7GHJqHl9Xiz/iweFdb5GMTM1aj
ML0JHq5ZXgwUXZrEtHEUTrShp4F3fdIwr2Le/WWkm0NKhXtbmWkOtjokaPMvivtq
CH3ynH6zF+0AePV/DLfdIawE+Fg8dTrKatU64UFGSGTtV1Ium49jbpA1GK9jHaTu
KerXUAIvwytfmJUNyJ0v5dQSz6f0P5p5av2sSKvILtM1jOL1C6MXsky25Jk6jmFB
JRBc6tld6aoc9CuyvLvaF7eBkqGmRaXconExdRmB103z7V2FNFrmjyCK1JqLXhzn
DWNVsRfoV/medFPh9nx8cJQ+b5S9D2DxAskHWJrcxdiRw4QYU6Bopy8I2Xy/6fOL
5umbDZzbZC5eP0rWpvVIW86n1u6c5LsnsuOe24cncxNA2Pic/2jlWcBouivPxPkp
jV4q0UqBnbpOyrkUbiuQiJWrxynFYhRC5emnhXewbUcKYbteW0fWo5yPEpxF4i+U
b9qWUtXGV9QWZVpE/dcNSuxyQuESizXns3SJ++nLrlOq/Idq/d/0NiZlyWyhn6zs
xlYiQtrGNYg1S/3jCdJIoAqjeSt+qVQNjLEQmG9c+Li8eFn+ykvS4Gz/Xq/C5n9c
w8B92CzqaukLRl5EfriHAB3l35WL4Z8qeqkwKJ6jaPf4nzGHD2I/QT9tq0xWlFYe
8MTMkDXery8YMbNWUo65M+MhfuFS+9Rjm4f7v3NsRBZhlxwV2HoksKDd1TPF2t1X
UL4M0d40kPZ+rOdg+0RkKWVkuSPdHypjiJ3dpPMU2gBqwC8Jt1ga1cA9X+qVcPMq
nTAHQSNFLaUmLTflv3TxBZ0fkwT1Cxwd3rEMUSiIlbZMuUVvaFNbsUA5kCYkkgqh
XE2uWx53ptAdLvP+zfHV80goGFOQSdlvAbWeXt6Kzh0/a6yCYIBqq3xU4U/pmZAW
EyM2TGBNo2kmXvhay9hTR1J7AhqU/c4lHsgK4yeYgFfoIJXHvwFBEeoVAvH5OWbk
VYLOx3AyvVLW+72RNhYt4F9xJtHuqPOBKbuFUJc246fdJnSVdLLnG3xTb29OAM9N
Sz3+1Twq3v18GqeWlhAgwEmQsbO02o72oddtLcNoawElQwY2OfHlVqdpQdmsDXQ8
lpSeARJQLYKe4DA9PEpSaZXaIbXU5OOZxYwDo+vpJUXy3xYuVtZXDZvBtXc27AAL
BKpGE3Eu3ElW7QqZfYdJkT9Pb6wCXPc/fXMYObxCrOP+mPipbD+o8tDstJBgke7C
ZcJ9IskYKnL//bGqYAzcOqB0TICnCHALHneoxGhQZ1p+FUbga/8P01FEoGUNImhw
1nStEG2GX/VV2LJv4MKmPldi4uLOK285I/U6nWRIj47ZUFhb59DfrSn7EZ7mDf8f
Xyvh7bMRIcyybaalFf8b6+m07ERkD5vkJ8ctx80jKMxpdTLVJQu+tmXCwgjQpH62
vFbn3GZgGMeBeMwNZqrv+RPT6bxioX1Zwa+PXQjEzcHcEHYy7jdgF6iu4CcoymDN
oLmyjgk4QD7VPTFz3/7fP+T357GEenM7FtH87a2o15U784KNVPyl/VUtWo3sxvVX
lco0fSllJKqBB/UwtoddvF9YP9n247TFEs4Ed8UTXY/KYofsCjxcJkrkwqfqHji5
3DR2l3xTfvB6+2eQ52zPYuIn1Rbiq7x3/yuraDG5Cn8MYdxrcGtaWSbEv9PGqicD
SdpvEy0dnGXIagmIspgvJj3albrvaruznNdX8RZpPTDdBYYVLdxz2Oxh8hPgvigg
YR1fNwuwXQTU+/21tO6jfewm28BsdjHFptSnb9ncgG51vKTgD/ZQvN70f0SEk3/s
sMaIG4uvR8SwsE7WKZCIRZkppplEGIEjyyI0Co21ogpf+rDg4frMdx6xtmWB3WEf
soeCpwEBuRTuOKm2HBOz5rkrOnX7y6aXUv/q3n5ng0sRuSKW1pyNqO/ac1vKjseA
SfM7T7JH9WbCBLYgCErx4cKHH3aCnt+emO2RV/dg/KBqYH2ZyWMbqvlkQkwIyimN
C1c5RHCc3uyxaHaB3gKzhFSNPttBcTriClfn77g5TXzY/LQ4W80UlQT3/7lhlfD6
Ql3CUVivgQQp3b5QfZBRjl7/wjHoM1RTf9ULnz5sd+xjIxiZE2ouq5LxyShBIMjL
oJodj+3m1dHiLf0CluM7qOWF8E63BNGAoNS1hW/4nKmKr44RUdIQ7oYmjmWAZl5i
DFMCIw5kroEfrUb74O6S8VFKs8aV7p95PtWWPX/72xFW3Sdfq5susUXJVUROxKqS
xdzH3dvyBsS7UVJalBRAxP66W447mbXsOeM2kpXC+t8PssYCVeTKyHTsskpixEwv
v4ra/VNqtkPIrdzY78cNZPeVf9Yjm1O6p7aIKKhFOfEyveezEuAQ6vTjkd75vOx6
eRMLMzHpdDxkYA6KhYLqHzjQ9q3/nmB8u3fE6YTiMqtbWfVJ6RdZ/xcnmMVEdcGL
7t0ujJ7GBEG0InrNuE75XpJD0u+I3LwyQmXri1Sg8DgRXMmAQcicCOrlOmPDBfyG
NpNIrvHCMrYVCEe7Iv0S0Euq6042joRb3+d8XF566+vJc/AqZ21SViK9WW7TEb9H
RIt7TLRFVH40ApdH29t2UdzVqce4uS9u4LkIanrNxYwzWOr/qOmWO5JR5q82Jj0W
YJFVCNf56VVz293wszvg5vWHBzkUPAhgNmAJc0y5R+R+YrOWTWuPlC/9sdjzp+dK
rYm7o0desGbwpzmE2vla14MfkC0H0R2oUSTPaTBZaMlBdFRNYKhNbFCuTGjg9OtU
JfjCscV/Hq9ClBnGuS+2I9+8kWVBEtk1390rzO1C7oEUtTmLm5LGtRRFUpMUyDdq
kE8qr+ASg67shEJUmWLWq8Zymf36MoUJsNJNRhZAwTi5OhaBOfBgMmwxmuPj7pG5
BZpg6ilZ69HcebqOnGrOGwSHe+pR7UUoB8DffNEzOVcbyBcC/zg5ca4rWOvcYGc7
HDdg6g6sD5lNc+RItsU5lfGZtGDbwYtX+3HHW3GMZa/o79i84m5/BOr0qFDSqDIc
BbxIvkMGEODgEJmd41W3E9rmYOenlkIizb0cfmGR/TbJACLjhKM8FtIkAUI3Dh9+
vtEWjLspIdxWUwrcj5/YJgOW0OMahjaNQ90svGuQo3IVhMVUdnWVqdHHzaNdgsRf
AoBIul2mp//0HeckoyglZSyBP54YtUUjapoxNuYa8W5cEvgoLTNDvv1vAYZ2hYFG
dIV6j3I7dSGop2whVQFbxxsssrgHQbUeacnxNfgQC5bMIlgtSkHag2iDwjdaRIch
LCcj62MRz0ixX2ueIsVAeOodOxByiI0tkKcm24CingaosKSCi+0u8uJoyntLyC7D
4hASbtY4WBj4DGgJ7R/rjcB8QvJqogcLGSehv6fZcrjGLZocJD1rhYFFQtJtrk5u
rFx2etJ5UlCCCPfHt3rAp2TmSt1VjzUXFydHRPCI+GJOCqMc2upuNsKtg9+crwuG
37icWjK28l9pNa2w+VCE3/PvTflLfA7iiCo48tDUCWeo5kbScvTEl0aLkKf0N7lh
ZhLB2HN36/FcxoyxIPxp8q8Hr0rnSfDXVM1jSCh7nu2VYcxVOmpR6eVc8BgEuL3L
OyUK3L9Uz9s4PMIU1UscDKPptqWDzSKTkezcFhVk8LGqtfLvgJ9FMnBXVTXZs3df
Cb6gzVMgzO1GCtLEzXmdGnrf/+kEGWFD26cY3Sl2q7pId5D+y33wJgwSQcNA+x70
sUQqbeBDO71UIUi52pzYBRfTkWSmuObQyqSiIIpmmE78HvUrclESF5hkERGPEWZR
iXr6CZ4bXHg+Y5QdrnO5P2WHEKrXjSVn65DiVy6dFxse0n7mCBU2MjlsdZISUgCZ
u7QSKlJUi+xJE1BXp9+tqEcxJT0g9AjisT8es3hvnod3Fc7Fwz5MCKq21+z6XOlK
xuJMyF1WRWfLIt7OzH8th1Z6/wKPN7NONgKWAUiFuQ3rd4Wydypce76EzNX049FW
/VVUUaCYQaZG5MhrqALPcBy0bzUqNu25WlmUjAScE48tnrAldIpyN4OYFfAoJcQU
hsd9+TSF5cIXD33Ry76rLdcgndFQCb8nOpFmRRFKerJrPL1NWJ4xQQuGgA67kk5h
2JjNFWPHLX1oBTr4GBy6880ngrUckAuukdBN4mru7fyJ9wePGCIsy8k8RC+VaeiJ
etdkdxvdixOv4CIW0yflDozVUI4ndM48vtLc/k6gR8ycgYEQNicOKAiroC6FYO9Y
A0uBXZkmhbI3d6rpji0iJZEJluV/aYm9658lB0qy6OdufRezmi4gVjM7tN3yu5cH
lUr6XNK0GRmgwar6ApxMhDo/2bHnYn5EzPIyus4nlR+RJqaWiIhaa2ANhFtoR50T
jVKdvW09Z1U5xueqfJ6Cq+JXyo7p/hUJEpMZaFS7NCwTcnEkXAfQ676QiMpH3yx4
NWsgnV7eJiU7PlcPw0HkjAg6iqTNcpd9DLzck72e4cTJbB+nCKaRqQS7inaZkf0j
jdD4iNdPYowxeJIB+QBJ1c3KCv90P5wsElDiQmT19BOJlVjNbha5dMs4yKNyGF6+
lUh/rTYPDkt4e/qljkmbi7bvb0Mlu4udKIWlzNGS7mD+8XnR/x2OD2FlnObDj26A
a5/U84iYIdwvGPjTvBvpKMI1I9EAXY7O+9QZ817E2l7BY0XgFBuK/hbe/6elvuj/
vnBIBweJU6+UrFiqGrEF2SDnNNdxPUYkR39AJNSaMZDIUL+Zpw65oD6DWb7iXu/3
zsZgpZi18v9WBuOAhZCmMiex4+ksWibudHfVs3dbXt51XGd3USl2Jnulczc76aPA
xW4pYUFgdxDClYNWjlSwViccJHRt9YGltZSNxFPzkQUKHf+hqna4h6ZX51aBT3a6
i8whLWM4fgq0tPle41rad91R9ECaAxxRepP5JZzGYPwJ/PAbMgYkGgViFDYAsTlZ
1SF0oohSpUS8NCPx3Lt19dELxqDQtyhmZXxIc4gF6N0PwCZF5/je+Y3H5A3D4Z4n
QUbnmR3Pq7/R7Lw6yCMLoGwaMHoQdxKYtSrzQqgll5aVwvfLlRrX+PGQ4GFpyIqi
jQHnTR8ILaH4KKhjupWGjN5v9kiFaZ0UHw3SWC68coSxRjbFOvXKaqYy5oPvXObZ
cbTTjKQi55+ApHBEx3SxQMa0ypqkY9Hrfr/tjJLzINNInBu0T3m8uX2hX5Jt1h91
HqXwt2M+b4UOBzuYSnZ9e9iLqQZPuMXXMiz9AWIbUDWotJILO8/Dilz1/pwKSnmM
vOJp9zn47vVXAnpJ1buTgNBGx2V/apDilQZi8Ui/vq+l/H6XabNi2NEmnTuFQK3C
JVxu0yarYwLPU33SzhcJ5WE1Tjl7CUIV5EOcqJ2elsQY5XNapLWXuis0DCQe+CnH
h/YAgBYNiXo6Bzuovm2H4/a75VICMBBEBDeKrNHU+FgW2DZQMR/kpKqmMta3+3hp
tZBi5pYZ80VpTfpMk4kFYvn/LtOq85eCWoiCLKe58DTP19MuX1hY/0jvUwATbFKn
m9qXfn7tSLWT+tHcJyx3+xqFhISWUDIhrtRKzKYEGLh3ryu0kl53jrG5kCvvzBFr
UZA+KlID6ufA8iDRgD3J2CKwx0QYmSx1UStkt+n4KRBDdppdAxuZI9IKDjclXgaz
fXiMt3abb+Jks8qMXeC5NyC+vo0Vb3z9dY1mJo/XrlITqMf7YpAewHrr0yPaRvog
HkOZ4quRU0cObkNHOxkFArmwqXFqSGLWjajMpVOfXEZmDkdE/sMzs/hOBvEhlXuG
fq5Nsm7BolfclD28Ahfrlz3cKz7AO0MkecQdAdhu3WW2IoqrWF9OcM0SND71xGkB
Lr9LB/1Tqc/NL4SQPNz+/SOTSd1yrHao6H/pksLj0bv/UtkQigdvDe38J521ApYv
iDXs2ynbHGs54FAhszUn4Eiu10WGhK+EVIqHu//41fXsjGqIoF69OLHqKxldLxCC
pUZPo2JIy/Atzp9EGU4fJNRJxOwLFugAL8iF+cnFfc5Hi6vzF6MOkKv9m519V+Gi
fn6PxPChHN4Gd88ZRUEsQ2MYl7VM03hNyaMqpL5CLchS2J5i0Ni4Wbob9jDbUyQh
iq+GYU+GxJtiZJzWHjRiDdsD7sPmP9qdgyX6JXt/42lMwdzsycXa93GiaNQrAShJ
lO4rfwl2RFGfcUEk7AbH0zXVAsT3LXBmJpUogETtj7phaMyS3SwxGSfdqWr/D1d/
2qKkKa8j99GFG0FVvkXmkLdx0aEBBpOe0W3W0G2Zd0qlWATsHFL72v7eiDyAltrM
q5XGEJrcJpxxaCFXVHi+ou0P/LVjsx/yAaLUE+DwBhYUwPGidmfpjoct1Et4873M
hW85VRJQt9jnivepn0AIZvdLjNAbrdihBwpcwXZ8cbVEQMrWfduPdKqYRIKblMyV
n1Ry75NXNWVAv+1pfpE8f+DOouFa1WWPIWRfhnCfzI3QKw6i422lzR1GP3A0ADoH
XiJpLzCVym7AX/avcvzIeq5eON6TrlO4D/6kjo+UlBNoVoiJqY6rq8uQhQ1QTa2E
RlVlPpGSuEK2Pd8OWkFlB4WN5VrcKCbqFUK0S5sofp2qUgDherrzjqx0Qn+I6b8G
/3Lk4X20ESyjTa4ytb5YUIkT2renaVglapXAALmL4I1gDvfK+5OoPPXFZ9sZoc/o
+mi4cRSh6/FOW2zY3xgsBvdiSxRIfqPmZJrq8qnlUIEW96RW5eFKgLmfsKOn6xma
dlWJsUJjhZ5YzViJKo/nTR1yb8nKbkA2sElJYfgQgsUnMpCkiJ3/G8lF/msFwtoM
4ehM43hvf9HLzzLNKZY+S+eZiY8oSQ4+2VRf5lKMjNnU7DH03u7wUWjBBHCcbb5k
2wXoHTfNeCyMQQ/Uld5ABPAoaPzx8w8d862boD7qvmf90jsE0cE7EWDSelwXvDA+
e0YhgxuRjVAUUhXN/riGZvYQTlrj525IxB/xE6h48qatRboaMlmr+b5mD/DuB86T
OtcP7LvH4LSgUUogDAXkCkQzSan37DtFUYTTft8pqTaSiijrLyEATduR6ylyAHPJ
l0143+rfxC1TXcBsgXpu7SMlPMOlCY6y8PkWfu1wZHYB4bK1m2qZRmfGT5eH9HA0
ZTV9EfOaRAImHM8dDOWQSZnUcBmugQjERkMDgofRpEw2/jyoOfCn0dTpvXJ35PUL
9DifYIURmQwMEtMtgxjIDqxgA85Y9Cjor9ZNpOJUg5gVPLsq3TDE5HSURaxFMWPa
IRyvVFjyzqsRnBkKlM/eWq6nuu+/oN3FFCn0Jo9Lt3tFPm+lIHkPedXxJf7FlEUm
Ee9XgWYQixjEPQBmPS7oXn4br4fIzk4I6XuELrAjeMcrEUIGBV07MOK70YHn6GJb
mSDq5vS+o7Ujq7m1asdCHQOBm3XaeCoSzf/0oViFmT8LlvQOcW9SycehJSt6Fonk
UNM0Q0NeKHFSvWd/d+l93i5V6UNz2F2u7zgJ8W1xIxtRlpbP+1wOhSM/3Le+2B3Z
5V9kUzVhDzR5+Zj5B6HEE67HsT/WY2hW5h2LWrXK7QdTJ868XWkD2FoPm4792/7I
AgInOArZ9P9EzH9wakSrB2pcKlmFI2eHH3ItzLFy/i6n1lUYDh/UFMbassYfZuX9
3COoFlHpbUwUpJtMjbOAHet1JwKYKqV1gO7zKQYu4DmEQ/o9TPx2RxOVAwRDEUCg
QwUY0F65A46oLGKZYIuhrbhSOgd0kAmI6bNvkdfpJFdFP+bJrdKtIXk984nMieNv
MTazUADs76DLfbY9KdFsGhB0NTVIGoUn+lmXBZyJQB4T4SU9vS633GIzSWT6FDLQ
CkUhlVIMSX+tzIY4OXLyqChcB5ixeyoA8O8ih40EKhbqOYCJR/Xc7GjBJjqR9jxC
SEqZi0V8ITJ28r4iZqK0UQ6FDv4sDaqWS8xrtBo+WLUHIKZ5b5bCZRdEhtXmqufM
VH+yS+n8on19WafT/pDj90UcuG3s+kyZztCXq3eudGt9t+D4lmre2XHnaHnMxMmw
8Q+eiU46hacbPe3uIYk9w2J/gPYlVB9CR9YNczyDsaP4e93e544BLO9dKJ6bnyVt
FvXV+4AkvC2sFWMvgwmidEhcWYxVkI2A+CimDJotJu5mW9PvQG6Vin0kfUwGZdff
/KZtC+d5ShdfPulfgLtr4fTvxXjntrS7W4dfJwXNdVjX0wdMVzZGnw97y3Pm1DoV
TmGNJAZgVVQQ0Cu/az5zw54j+rnCUAc99Z8N75QrifEzafsRM43jDdRD4oBHJ8CB
WSzo72X5SCf52iZWAHqT3PelmQLdzdbxdSuMo31HtyLQmBFtamF4KS1OYtzKTWue
jWsaKYpk5WQcvrRoKryDvFBF7ImelZpeynXsIn80i8P182scPdeG+b6U9hUwu8qR
FsbW/EJvBO3/S/+Ig6Cnbmj9rDUi+XKk96VSARe6HTFoCTi7kmM3JfRaSoAW9qev
oHxrOwW1TrxFVLfjlfi7ZVkLpA1+2l360m7vPyrRVCLtVhR9hPUMdzJ+Oo783kol
lR3T5PRESQWQII2K1Y3BgtbzoEHwc9yBZ4bGXYfFwHcOyKLWWN44+6+lIIYwn1Lf
QwfFHc98XhEmJpd9yt633/qJPectGFm++hL1QiM+n3GCMLt7VEbkWzMlOwGZIeb3
L8G4MgvpqrscTNXobUvVu9JnkiOZ3NznLdyUQJ+KF9FvApc9DATzwOJw53YtJdQJ
Cf6/8hn9yLh/cHx5/hLRECN/So2dCfBnfs3KujifeQlpdc8VrYLFXdnJaOWkjdz3
nNGrautjeFAkFV4h+qtR6rL+v09yM3J8GhtCw4MqHtTV6rBAH0anEb3R5OSELyd2
lE9bL5XwMm+kGbsmWW8SbLsyCIUraNizVrxO1evnGba/vIq4zW1TUQE6dIdCtb4c
/m2Cpotbd9J61KL7BYZGIfjmvcoVcksDi51v3fEVZy7kE0TaxdHKdbS0tf+ZEX7R
CCFLnxYY60zcHpH0ks9INGb9gjH7vsOj+GYMvjfSSXgkPwcM+IOsZYhOOW5eGLDi
UHjxmfMOIIAgsV7axEVBFk/0QYrPWil5CMmdW/VODaTFGR4aXwpUORgy/CY9CU7G
KemND87Q4JbmjcUYp+BUfzzGmieT0CiN4x6l8OuNijSCgy8ST9JboeVY80Ztznfm
ZD5msp1CRN3SvufEMQ+o1hUyfq6/I6Ft/5T1hH0VsOCd192DCb9ODRa76cb2czM8
fHSryYMYO4gbNCNZwCxsba0Jycn6iZe5qvN0PnPApbpEoCJIBQXLW9XOltXgNMRw
wNvFsFvwyTQp0kc6XUdjZyTixHc2S+2aaIuHz9FXRe3GS3jbmCObiSwtXR0mMzKy
mUHJ+a4CYyhikpEgCpVwd6xOQAtGXt7c4scwMf8QnXg+iuJk7FQ8SJDSoXzybZil
5kAqpIDjdiVTgG4y6e2KBtCDBVzGcuX6baRyIFJzeNiViZtXioXe4YgR6JJP8fnJ
mwJpnAThWZFgtuBQ0zfO1+bYpaYSNdGB3xmMKQGIglgnVJQhLNZD4s4lObAxFT6I
Y7gEVlIer3V88yKvckH1/acDA1DOuHwzWdLkvogZC8WB6fYEKMUg3HOdhfyXJvzz
dPg+XSPuQmfTSHsINnDQ7EKkDbvyjsd8U/NrQn9z/r2vm604Eywm5NYqQBfWe8Iu
ssXHXqjgJ2A7jA6PQz7QCCODfdGJoDh0wEt/vQPVuUkyj83t2D5rnOdp+lJ/Dq3G
aAKjaXRIyYd4ipV2AP3HTnnz0Dk7LkRA+uZm0BPmUQZdO+UL3IzrZe5d2RCnjmKh
XsE+BwboDUddFYBHHV/kSBtXCWD0f2eCiZkFrY1TLd98ZYhxyy3ki9As+1r+WaN2
gALsonI9lDw5HTOoQ+NOavonE4r/oTt1BsRwAjeH9mU4D6ypOeXUuIPuJNlK8fwN
MWvw9iHMoNMWu51buAxKGR0X53uQhUKkf445y9+RtDp7cEWKADW0LxqskbCQsqX+
uRIvUK31fR/5PrtEm5K1CHZqIOEPRAGzMvPoRmWgl6Wg1b3J9zSUeGQjxnWFUhd4
xKCBB2k7visov73gN/BlGitI0MncMXUYhfOnBVK7jDmMYxVOBciRE5+aumw/akhd
NKyDIwT2IBUlUmrjfr9vc53pq4kcNN8TpxJkyRnDpW8LPZjAg+R1GGqgWnHG9bmR
ZAsJ4oqZiExXgfN5s2Oe0Q+/YVeuxr0XRZXyC4inpH0=
`pragma protect end_protected
