// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:35:43 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
DiJAWDN2gpsAe5Oml0oqYRP3BEpiT8CYZb+Qhg6fVfqkHuAma9RpidO1Pn+GOAUC
k8LWvbp4LUX6wJkthXhCjNAQy66haFJR26X94AY6xy8OOh32O4+CI/4LAlbN+WlU
QiugwQa0JH5eQEjbMuOJW+sagHDwt7Y7nWkCucqu2ig=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 6368)
7KhchO9Lczj7GBuGbUHlbIowl3kP4GbgGIuj3gDsOhyXnNg+S9a4BNSCC/YCF2ZJ
14S3FVBZiHSZpLYrFMmd4QQdRhAiUhXbukGpUABB4n1I3mo7omtmxEgaDjTCFUCj
YIayx0P+/kcdiwkJDlvk0dCGmiftDyPHhGEKe0kdgBcje92ranLaCdPSEjGNrTN0
YpB7sOed1MJYrYxyaCgkwQs6kjxnaXU2+ilGIt+dwctoG7TUgn2quoe2QUOwdiFz
+Q+o8PSW+dJAJCjcB559ogk/5Pm4C0oyO009ysqDcIRipZMdM0GuA/s2OnTaUMQx
RWIwcBwHgqcp8EWWcZTu1BTFr0vv0nK7KTodavHtEzMtkMLND7FUET5E1uDoJ05j
HroeZ+conlXsRP0Angr15kjUc1Zo9GbkFa2zhTTtU5Cx8aE5M9FNj0AqncXnBMa7
jqVRPqmP8LYIowBdr8sTpb2Kusa2wwAUnDGzo2y7ixUBWzjdI29K6OMwpvUktU0v
tnLI/t9b2JnxGZnmFRbjw8NMOobUhAOmyOuwvhs/tpN/NoLnGFr3k9gTKbfKBcQu
q5KwLJLynbE56sHUTTC61XAfibo5tYjtDyRe5Q3vJDxycFgQza6X5IEJWDuJnnSg
CBec8oKLUkyUSAwK7+1QR/XHGtz77MKs7liXTZUkJATdBZwtoaXMdtos0Wt9kmXe
GedIGGjnXsHoO6c2k8EOuWW8YjUf+RPaG5BDMgnLTR0o4Khm5qhthxNfd4dy3VdU
qqJbXfR+BMY8aSBrzOmFnoykr4TkbXVY894R2HcBcm8kirAfVfT2Og/MVdKbC2F9
d37cnLxnJBueSW2fEqME9QaBwk+0lkpCycgL2RavAZloE5bTSAeQWXql2Nh1yBnJ
vnwTEHNLVaWzRoc9/Kv7OL1DeamVYULNpDA8WgOeGNChzoOzR4Y0Ph3DWU2ASLja
iatdayqwGBnGSSyMVnb49u1EIqw5UtJzB6IuGUz7GM9iFWZ7NLER4/Ar59JDnSQ4
FKLmJT45hL9Z5FzcV8wRTaIhkmJcF7bcPDAlWznJMC9gD9iZcMMQNuYS1sJHcwjK
1A/RMwsn/RwPshhl87febAw8GZ+2agoT4+PoJh2QLv1Cfr3SVQmIFcmYe+ccFADn
HmGr8og+r49cZ49zGTOpjRjxtK8TllpalndNqBo6SxlyiWMTlMlIpunRymvUcsUT
1l1hm9f2DYHxEFHsED8aedZqpF5FpUbsF6Ru0aJvHNFJsH82Cot20hH/ptORgW9j
C14GLaSJiHAO5ZGU4sY6//0I2XdNgqjctdF1117YxMkIGmgN4lFvp83XRRJJW1O+
BcETL4kqsRcJkUBsTpJTJqm/yWU+8yRrFTi5hTzqnDWrv6cVAaxpGJvsI1swntx3
I8eOBOSVlBdlHUsFEphbyah4CrN7R0HZmK6lbq4mX3xIty3QXaYWYXMGdi8o/ulq
JtPzke6Ubhh55BSVwAehoDeD6B/SqwcZp8CuPmvnWoMSlGfu+oCXUfEOhoRMbzWs
l2/xwjbKMBAOldpm2rhZedfAhL12LSz+nH4AOylltup0Bzf/0mjZdJuVrkAeFKRz
30Go+kX/cYdJe6kvl8TI3CGsLxNeYiSOnYvt8Ga6CNQMxEW6fTddiYqUEvShUO8H
9mu5cB29AxSOh/ZZHSWW7EBIbeWfyChfwC7SKmQq2+CvFtwxCPDDpiKNRAdRBnua
e3kjZrqNnsPAbzPnVEVsF4OYzLPfqKTfALCxliua3svzTS+5m3XZpm91n8/SJphu
BNfMjs5U3hn39U4u7MqPB/4gPS+OOVdOgfaIZScoAVQUY0EmukCV8WvtZHkWKmTF
CmcPuxHyqnhmxsIkWZ9HLuYbZ1ZIWVKUH9bZfAM62UocN0V2RZl+anTijzDN1mSM
pk+ud/O1Qc/NUoW9zguU8HJ9rzSMUKctdA2DrpW0lmF+2vcbK4+GZrzz1Xknv/tz
3dKe92DJ03L22NIToc/Qow7uyBZLBCtMavC0s/PC1SHEgWrB9wOTa9yJj+7HMfGr
WtVX4USWSJkoR3bu9/ClsSV9Zbuldzs9DQCZJzNTuNd0uscVCJVJuixYhOtSbn9i
iwzbcJbvYPLEA2oHElQCqiRFBqc+lbb6hGG+6FkTpoIPCJ9DTK1jOu8qcglfLbKs
T65X7CE7EVWwXG/NUYwvt8ewkae1eTFKTJb2frSClgo8AHaf+6RYc9f99ioW6f1a
tkj9FbXUWJBDVlP7Ib8cU/08TYdTaDFS5sBYd/oLKm6H+5RnPyCngkA/iilhWhsG
EkR49SehcIdiIe0419dZQQ5dvhZynIPEp5ag1zJsXlVnDMzKLxc/kGekHZFjyQas
w7V2a4935WqT7KCejQCPv91adAqzKw5UBvbp52yKSYjG9h+XJ4cNNd+WHXcItvdM
Cv3NK1T9yrUYtHryiuXTrqtLoME/qYE3yYVTpGU0lkIIqjNDg+Ct+tc8WxpeiI/J
JjLGts7jPPvxKiQeD8OYG9yHtd14oB6HwDXdu2gstkCXbnQXS06C7iQ4bc9/P0uC
gNvm2NQz8qECR8T6D6lM2oj8AxLN1rbD3+TCEI9kzlkysKTI15C6R6YQmWJJkza7
yzfZDB66BIAooEYJ6dOEvuKM5PfXEg4PQpC9kzWAO17wWaWj0lVWqAuZnGxmy8z/
6Ro6ubLfknSPyFiCvh7EoSCREbmji/ByBonPJf4HHswK6u28T3cymF3WrqgWN5sl
07ohTB4NaM5LmuT3EM+rsifKYhbUhBOYyDO3xWZtxyu3sKpmaMNhZtpKyjdWmcES
m32gMC/SPbRKiP76prORZ9sPyKzu/i4c4572mMUOqeXClWt9vuE0engurlbCCyPw
Fkn4Q7yvb5LkYVG3R3QKNvTuO8uE775PJq9+5mLjYP/0WBkbML4hXUWugmNbwk44
+RdM2YaOR/i1t7dSlAUXGhfi798vFbBtXatA6fpEa7hotkb9N1wRAgAAP35dkTYz
PtuhsUQQK7heosyb6R3cHnZy++Fds7cg1vP7SSGTjszibesY7LMXc2SWOLIRe0Sz
Hti5ZV9eVQM7AhQn9jBjA3pqXtHMPMOE6E6ulyWlrLtDcCCWrOtNbPTyhzC9TfcI
GlCdrAujwn6JKgdNh2dHrnPOKS8BmnK74r4q4pk/2/EFTSJGqToG2ptduN7Q6o5V
oy4Mqgam86UYJfkDk6LEdzBjvxAFI3Ppget29ukgoHcuY/Ny6s3jKY7uwZfXZ4Fi
1I2FcQOR8OtzB9YQuFvYenss6WW6ecZNZfkbI0WIL+mQc187IculnhNH8myRs54S
4O/LQz6NBkEAKmKb9J1jeWcGPWQrExCenjTiRt8GZiXIODH/nWdABLb5XrlwO83D
O1c52dHTqaqQQsKGaXsl7VQkv0UoLrSqjeN/pIfImu8zgAfvGmspjagN55sOa0AY
dTOeKjpsAmgoQKyBD5gtA8Q3ILdC3FzyEYAB5erLfl7qTZnsKVgP3w/iQ2IOaDHR
pjv2OUQE3UVHJzroW2OUd2ktZqOyf0BgTb+n744n+WnehJZYYsc8+i1BwshFLV6l
eBfeTblsgLWsg5izT3ifOWsu/7mN3qTIrGBM14/TlBh4bEoBcuAGoi09LjLLpbnm
5oh1Urq/bZ12YK7CGIdXheWLudWczwdBRR4MchOn4RTaFPlUFC/jLPQswfxyWLUt
Fmo4YoMZGTUKPKeVE6kH5E4wXDOMgQh9L8Kk17fT9fangLCIP/9p2lnoHwDQSJzl
Nfja4SJ+b8S7+TJVcsTQYSKo7gMOJOzNhY1KEIP+a26Q7scSKqHANxSjuvOqH98z
h80ORC+DuX3pYb6rSbwBKNp8qkHQVs+3Ibe3pFR+L33kPmS0OCCRBId3pfNBP+PY
iKlKGWbJTIi5qnFZtOMbwf/z38sIt6SM7O8fKI6cI0TjFFygIKbf+7DMdAmERe1h
Daepjh1wZ915KmK8u3bQD8smMtTm0rxX6kptZkBBdOS7YFQaLc/FvAoynWW5pi6S
ZsXsina/tRazymwwTHi67Hdb02bhzT2gSGSr4sJwFyMQeqWB9/vIkwmFQqnXJ2Dy
U0+IeQjU23qEb8rF89xipZRQ99oE3PhiDrzBJe48aQzh/UU4KiIJeF4p4s1SU6Bs
IAy3vdnsenOnfPLYMLbiw7LhL8IsWqtwV2zPrfv8gcAWusEpvTODCcDS9Q7yz17r
qUAPnRLh58LNXQZNvWkgizohZP9fjXm7ULJ3vyZy0GP73ZpQ+d59e0kVclGWbLzk
8PF6/M0jlwzImbtEutxunBSFVfPQuSmA2SOSVdGxzDAOVl3sR4e8zg6RDUz7h3ur
tUS0C2y5bem5tqQLMJ74ji6RUxWQLpwod2Brx4NqSu5VU4gEl0TKON8XuBxWiuDC
pkKZGpD6vz6oBIJ/jKM17DVBCmvsN9NmFydBaOlN0DJ+sTyWkzXdv6sTl9WfUqI6
dxnKVO4sX/nX2ejBFeouVijRRbTSS0pKZNm7/hx/LG3jTnefLZHfWMK+gDP9Re79
cELxy0Zra8LCEfja9f0S2DvolIK+2cxQVwlSyfBTwEni84EqejchC8v4VeoE/cMd
duk0WXgoX9mDeVTjCd6wTrEd46ALBT1lmAKuOfD5Jus+7uDDF8U4am+S17x0aJ4l
Zn7/z+DI7IaKo3Mh8SMAepgi+0EWlwlAshqLcmPcRoB2d2Aih95io+wzzgko8ds/
Wc8hAfsVjtXNf6f3pDZ6P46XKc5E10zhf+9njHSyMdu3ldB4b7eYYsYNpzvjkpnw
Honn2I+UkatRlo11ZG3gp8IuTQS6MrWx4g1xo5SY3S2qcycYZHHarNXmSsbGezbg
t7O5F3xnLNMCdbR5U6Q/Nu4sA9TJSpfG56DLVVETFRHgSjGybF+3eRyexXLDa4II
pmGHQItXhXlCM2hPYv9eebCQoRrCWbNYjav0AYOSHqzPRUsLPDU+k6As9nFmO4Ul
nuYE4ldU3sI+9qz/cqv1zByABEkwmxAgDwzHAh2ASwTWSVhWWk4PY41ke9rxSb4K
DcOkC6x48bdZZnVWq7CqSQNGrGKiTBGMdCs0qwLHyJK7oGeqjnYEj8psAZGuqNAz
zouR+w95pZVyMsjg/oEN+4djhAhv4sl6XFPwXTUBnWd4Qrzt/1d0P0pl4EZq37U2
tBP3Aa7wBIyxSpnv+Xb2U3Q8LOkAUKgIfCr/qFCJB3bhVywQlXHHyKWDYShNZuPo
uOkN3xt723a3zSqGLu+mfeLecKmKL3/6lq7jC6aG3rh4aPBKcKxLD5BbJBIWv0EU
JTsHTN2M07he64rUB5N20muI/D8gZkmhd4e03vXcS3FWIU56UdUr7UjMDtNBerM2
51DHugZUSe1YkIJI0QyBie2nEQPQLWWxvNi0yzQN5ud7Jfam1g6GjYqHZ9niaMKG
s5URbpTajBqfkwzTUU0CUei+Q2I5bbOp8JSHmWtO5yG2L/3HnuEuFFFX5YDa/h4q
heJkrj8P+uafdk86Q19KRR5nKV7PB4ZApZ6dTJZHr7vhVuisupcvrfWDOYxWXgwN
a8Eem22D5m3AMATObWjqHu6X55G06SExYyY/HyAolaQpggjysPjJK60ZTB4Sb2Sy
NwL04p1m5pQyc0+V3wtvbRFiy+h6UGW5rIcgYaWR1x35uOsMRUzqCllQE9mrqZXH
khzWLIp5vC6WVZZMyqynkwrxgAfFkAdXv5IF+zE33ZeZUqgoEyJcJhymazZQ9cmu
LdhglpttQec8CMaR2u3z77bhjtu+uu3YtfU7uzwixMveETc9+t6nJnnTrcHjgn5b
qr+1PHExF/DAlXm2KgOfXnG67lgNaQKScwXoFim4cECm6EqNmv+lYuvvArk9pBbU
ZR6Jxk3Ey5204LCzKjmJjFNgKEmKfigzpsmlhbkVMbm1lsQA4ZnVcqGIYMLFxrGP
gbbaGH0veTrf4daH1r3Z+0Qm2gKor6+nEd+DiL7LiMwvOqlm7E4vlO30DjdQ16Hb
M9U+7l9El26+eDHmKTJmHCsDXy5cLb4OejgkW8a5I5eCCb49Iip2BP3YmQdVysva
/NVfT01ig/ZXBI+UjFPtPkgjLrgAIdoP2hDzMnkumODOhvjYLke+91sMGfyyfGSp
T+xTzo3VaxCEryLgdqkJS/x9Bp7tSr+WzwkmsYmiXxJ3zArlT10zD2byz9pnUAyR
OFHckxTRWOnag7CLLNyncgy/Y8BB9VDqA9fi73uXzYy1qK4y79E8aLk5pS82a5/1
kYcg2VCxj0KYE9z5A4q94bITpCkxuEgOpKufYtqb28Z+YMPEzBjsQ74niob8/eFn
gRG5jIHJl1iqZPIdGX5/4jz1t8zvK5xEcjTt36QRHsQLcTw/cShTEpe15IAZwkTA
zgk/EO9vwXuKSJia1ukeNbBSGcvZH6WUoRP7RfGMXhxcncjsLFLCdtojMTk+M7Fc
PH3Ns3ZXHscuN2GWMHvhTF8nM464A+J7+rT8M8Drwb+kbFT6a3ZCgx1Wtug/lvXF
2F8Juqaw7uwjGYdKOTgXedGuI30vDNCBe6hXoCABbS6mdBnk/zpTlSmzHgT95xb2
vW4DR6aN+I+ezCCyI+f09N3bKL6/lnTt95woer7x12MzKLMumB/6/tcB08pXvUoj
D9a380Ay11ypIGFIyG6gGjm75DBmExOorHeWz3B6cPuFA/RrkYhgFZ89tE+3mcl8
0AJ5Sdx6l2eKDLWkJxSCuDNOpDPXG3wadOmY/aAENZOm1q+fw0vbBVRlJ7bc6Alx
VT83iMN7fuVCSMNxSjyuL8o1qUlenPHleNhmanhqHoNjH33o9m0eRtmyGyOesnA0
uXkH4gm1FCc6y4yoTCgOzTwA6t1Ga93gnWIavOIdTFuJP8soMXXmWCum3DlLjyS7
mZGDZjrMddF1jn68BldRqBFTRqSxTvKtQcX+Czu9Bxuov/2RVhOilWe8QtYE6hrA
oDmTPXLxY/Okd/icinsTtFtL/keO8VwEUx4HhCKdQoQ9Czsowsj8zLbzMs4/ZW+x
kNU7/+5rUd7qKKh5e3+x3flYuTS/Be/vCqHElmmncQ0Vl8Z/ezxag0O281PSmblM
AIEiVOR9h2SWuJwL7rIAxeERm63bfFoJayjVmp799wH+SB7vO+DFiiTCpXK2vJ3v
ss0DP/+pH6TmAidXHH9x2HUE21Gf632dqezCHmz6PQKfGnOOH+gaEu5O7mpwK1Q3
KOSyrFGmIOXAN0Ry9bxeBucUwawpQmytsM992+5oi5RXo01QTlr5FB1NNpsb9vGD
PlQQlwDmxEJx/ZvflGztkFz/2N3xZCVWmw/qR+z7VqhBotCB6A1X2uhROTWoC1Ep
iowKOLFDrOFJ0EfAmZZs0WsrWxVDQIhmwu94yKjcUYVAsynrOw9KlJDGBxLCVrhH
Jkq2EtuEeI+yXAasnHKdZCucrXc1djNVDISkoIbDbfSZZtQNP4YjcOKZax+Iyasb
6wK3yDPIfNubP2GQZpajrN/5Lu/3OpApRzzSCniF/O8dxdlkuf/coccTXalR/o/8
sVtN0H8ItAM5IPE1RqgedS9FXG4e6Dsj3V6bH6A/K28vCFc9bW/04fLVmmnjPVn5
392s2tuCnXrfRCgAxIgIaXIZhrMI96g9jcJcjphhj/3GWYT/434VvhxRtD19u4oq
3cQ9Owmrbs/6a7YEtWDELBSh2m30xL5w2fKZTswmz0GmMdPSabwnApM0jkUMb+4L
aKOqcIXq1yThlUG2fFnR1AGMB1cOyIDo6YtqD6KTXoX0A4eiE+XQHBgLV2m3vXcS
G2Nv7YL6QmJYlCExpIp6zshuRK4uHdZxqDmHYQPadYjHyIUtA5xRBNyBescKgtV5
G95mQcTkaHrerVBjl2BNq8X5JhURH0FP3GA1uFni3b2k7pC4LGzBSgyBQ50mNIPf
2gy9e4C++QVVUSIlU9kIcbeaztPUEegKJbhVZ/kYLYtXQme/rQZT05wJKtOKVbFm
yVm5UWlUr3PXqQ92hBoHNTO4d91hj6mT/NQbLQ8rtOpxF9KeOWamfXmEQ9cY7G+3
QqnBNCEWx1goz5iuZWJqilk/RqVAJUr1KLMRFNPjmu7NXCLk7Qf239ke+pVERYf5
BM2eLUQeLOc2Pe4JbEfBSWyjaVVWzkT4fh+eqQ//EFr/6kYsmENV7KXcXVjitybH
8ltUdzKwNH6NObgmTkcBXvRohgizXdn2V8ezvCFPTXmKV/7yyJpWTnhMpRkXP8qM
PUY4I6YIw70WhF7fYKs/hr5WPAlUNPndMsqZ6/WQsLAUdFGZyHudErK1gn/okgJG
LpuWNA32C1Qxb9Wg7MPwtmCl/f1AMDyNJyU+e51MrsBL313W1geDFU5w1oK57G2s
VDyyAbQXpfom97c5tqBWrHEMRrzxfkx1j6gL4gyP/FgGNEf30L4AdKOfjuMBqGvg
RP4grv1WMBmYV3nxzastsc95wK+kBCC+PdurtL6/kPw=
`pragma protect end_protected
