// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
NcndUY70vsK32Xvbz1SF4UTK26EO2tLExVzH4UzAb7D8ZWF+FqX+rFI1TXZRKJtEAQq7qX+yII0B
PKOU/NfDXZIG6/PWgI+oLAoeYBR/WOdgVnudt8b3mR8pZOMvkoyOBmJu9GkZIhr/EMq52RYzSW36
A5Pogi6Iq2t4lHe1ZrpgUjWgcsqSVUo3Njbj9AbZ/mN1XzM7h1SDLOMo1KXuV+rlbQbOqTGI6RKq
Q1qES7uTYGXoa0lZTjvdirqXdUJOaKtwtjxHZKn02yBY0YdYjYo6K2jOJCFGklLyZngEmLNgNgZP
EX+rqA/fVB2289aabL0E4CZBnMy5gF8hvrSLqA==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
fAkPpEkw7LHu7d4niAABMvejxCErVbv21CmY9aVESHEAd4dV5NDiqFCmQUSrStMHyhwNw7bBvCJ9
ArR3g+1ipqLyHt3GA1BxqaKF9ZOxg/qOnXQ1G/ijNLcsv/NRlls/Q0HyqWeMAK7xkkg77y86bEeL
nq42vkwuhFm81wU4FvPCQk1y7fyavkik7QV5a0LsfbG7BpK7ohKLENGsvbM1xdsabIyXdyJAaMdQ
lsYdBsrg/DB7IJipn4vvWtLmA9AhLL2lnvjnITt4jjhdW7ot6n2/y/so49UetWVNkegcuJiYsUs/
6ZMc5CuLw2jsU0Wn91NKm5BlSZrsvAd4jvXsKAGn2PDSQGt6FYm5gCd/Qs8YW+grJ5jSoi9ohg2h
qnc7qQtV0UaJqduUcfxp85f40hRuh3dmEEVNEOZzbfqgjZ+c+oo6BRTOXiYy2MFmMN1Fv3KLeLhZ
dkWSZ8qncR7m8hssXeos0t76nO3frfOA+abchIAgpp0Fcmc+w/hPvviKEh1GzQaUGWpBPyDtdqa+
kkX8xoMEskKnrYuiGcFIVXjjpO9AhH26MxW+jos1+AHEebiAvcmmZdMoMC0tS1cF//tzd8wozamN
peyuFfXFCP4j8I5poxOGv3xh/fpveCNommFkOHTobSwhlxLu2aw034ii0d9+a0kJ7YWrQSmHLJTr
Gv0iEG1NMBzb54lgtvGeCxIqEIK4pAgy5134Ro1WZjn6xIv4BqSLtR0Af2GLl09pw7Q6IA0KY9uN
E0tLmmj1MYPw2mLqezjvMtbgquD7HFy8v9WN76FsymGhjhkNDqmpiMahhuDRX/7Kon+wN21lpkwc
SSVOTCDO3QNecRLF9AkhHd9hypAGssBiD4v1njmZn4H2kz5/mfQt50qUqJTGP0iew95YdjDlqjr0
IMd6FMf9hEKpMHaIuw5o7lvmKEngcLn7fCSfdV73Vg9P5QyX8z1GdTh8eQb72Rn/cO+c9k9hhM1u
gdBBzZdFFOz08f0OwrMzM9Nr8Xb+/xJUi3vvRxzpG413qpeESe8ECNsgbjKXaDOpJ9P1TxoGoK1Z
REcu5KiEG5linOndtiv19Zf8iiGoqA5er8eLVotkMVoF+85RSDYDNX/YurXZQkuHtXxqbmsMQ4G8
/qBs03TYL3gOz9l3N3rpdpGxV/+LREqzHcc/0uiO5xX1qa1DKezMdp2jEZunhLSx81S6Vp+CT/y1
GNao2lnIdJzjWY+U2NXsezTEprZUsXan81JtKgX/tNzLc4w4y4sX+SDdOi7RyQCG5BkmY7iFSh0y
7eKLaUVf1HytFepP5QHUy3LAIYrdcQr3jr5iD4TSjGHY5KW2dng23GPG6DeENDHCUEyaXBUv1qzZ
e5nKkGOpjrx2Rj+Orc8C+cp/xOYzP0MJZArzeAzThJYPjW5s6KLIWMZb/nztJ+XGfWkHLMeMyHy6
t37xxbNIdspT2CtzpzIgRqgMzA5kM21PS2bUY+gmU71np3uRFLejcuVPhGpdp/ZwE88xKpmDGnGN
F+GJf8tBukyLXBfxNMyIqMxfPy8swUcH/Bq5EQIe+1sARW/g9m8nrLbqfANRqceJ9bgnYpu9vqS9
8+hp1aPj/TPVCkryq/C+Oe3TnHxLybelbcPeJJg2VcVOgEZueXYeEUJtYzvs/bJXluSLZ0LONxRm
WsXW0iqZwwXCYcdwwBH9aRTHxDqMScbQy5yjPlypE6HWTjUYSU65P3XPHKknfBA1dM3hyN5vLEvY
so+FR8iFwrTTvMC3iYcLqfY5rmnz/5h/5DvXRZUDyzKugQGQ5/CBKTjDPBgFaaImby7IN/xfSPXi
2fDYFiNAf2nuLx6eJ7JrzAJaL1D0MDdUyHGovdKUMTGh+IIFw4sm/GfiYiPIGOJs8txjbulixvfJ
C+iagiJrHGy9rQNZ5uqt+c7AbVWyF8wUBI40EDVPOCh++iJGrXX7gxaneBMgvcVGMAK8GNty1Ckf
5eQwcGD62IkWvxc4QTOSz8RUoDdiH1QayVC+jRkot1HlNn13zz9kjZ9FKPjPsQu9aEjrxu9Ve/mV
5UoX7E42eLiEFkEADSkKXsp8mhQDpeGwc7dycnIduCDJwAJHfZqf4dWi2UY4B3QwmAzmx/f1DHHH
Z+Jcee0r+3YnezdF6vPi2LD8Ks2ZYJ4j1lIu9tnnFipaOxFlBUgVqzyIToyVzpUZEe/uEZ7VQMUh
ghHMtUfqoz9ooBu3T/h5CD65DC7eHUaaSJNiXKvLeo9moo0KdWTrw3yisQZYKl/Mzj1K51DM9J4I
gQFpnVD27u2qV2OpmXQs9RvUbB8SpoE09XjYFgf11s1cES+GCeaEkrR9yIuir4vDmX3H77s9QhVo
eXYQxliqjg3t4MJBLkk6Zeh06V9mbxUmn7izDwPdt6wXUUWuGTL8dt+mo7dIejrC4oOeNpWwNnKX
8PQrYn6N0GV87vOVGdYtEt3OJKgpaIN+VBXBtrDw8KK8gqPY0j0PbZ5QQ4Q3mdeJin2uRroTIvVX
puy4oFbdSvkyiZwHjF/EAdL4wV4INH+WZXdelOWu9XiBRVoesTa1HEm551F91YSypZg2e9Fm3cTD
xlMJv5TpxCPoXEMEyRxI7ZlUp/od4KghCx42TsS4LVaBV35u+1VcTzP7sUUspLuMZ8kR4a2wJ3VC
PTWf+radLdrI4d+UKXtxI8v65ga0oleGGj2OldFP2PYXa+qubnGiryQEmqzdU+EXYSIelTObSzH4
uYN/HF7R1adO/O7P3U5UfRfrYZ/NTfx+6url4VuYgCrTisPGqvUGUo3FbA06wkiDpMqM9VwtXyAy
oxhk3szi/wNVhW55NA8t2sfKH/DXxmO1drq+sPu1w3Wra/3lRXhffCe/wtdakvyr5651lOVdheT5
Pet5ChZnLll4xUdf+KzBgwL6XqqBSy+1azwgMrpDXJWsN2DqhCXuk/Td/DyO1SIPGZCVjzcSw9mz
hEXzNhb7Wtz/6Rq347sz9kxoMPYFwXYmT7EhSzqwu9KOGgq3OL44lQ7s+VoSQQnhQt4o7gzDwvOT
4XDf4iNsdBRTx7qmREwgJcpYB5PfNMNaGsuvx7WaWcmX4NP4nbj8DZEcVDSoOAfiLHlsS0eBk+RC
28Ql83/GShU9GWVyKOEsISt5hgocsinjaGRBI0je2rXmpGmzw5rqhlcoSVvR2MU5u8+rMiAACjjV
rEyWbxK/d/pZQ6Yuu9XgwRtX4DHApak26WaeQjIdYfD60XnXxVBlYu0SXFHivN6mS+AqzLdLGhFx
f0QOm4HMyvfeibskX1l/2yvfHDo48LbGkYmYb64ai207XUYqgZjb5A1AbqqtmaJyiRKWuZsh7B2P
06IhZs8xZpLvwyazK+ZLztXGfNU62oZJs/DukVz66HTUEDqHWCRWztPsbTQGUm5Lf/1t8kuOV22p
uqDDDfiW+BMkyR2ItKPLUmYHdGxBllgMtbIHhmK81ROvTjcXJnSpFF5mB+60usco3xFZ7DpAmeQF
EMcnLHtdiDdG6nvt9OEGHmhyX9JIttKFkVYBNX9DV0e/nCUgidwcYgRFTEB+F8JArc+igaCAoFGz
30all3ERzNP7ggnJ+PiOlKhv7MQT2Ff0chwmH6+MfpmIYJrjzLOmsk3oUR6cM9JOAfbY2sqfYV/Q
mkXiY9cWSthFTQ/K6yDwMx9DU+sli6ZgU3WyxAvXIMp6JWT2A25k2N4yIs7FY8/Vpt8HxnGyp8mj
FqN2fPJpexRLqs+Qw/gxKXU98/Vohu1JrOzXASK7R975uhyVlpxxnMlVpQjE6Ftm1MEAW9kW/iVD
K8fkqzkK20f9UlNwdsM091ixa+brxJfc1WNSJkR8pd1fCc88qG/hqvT00tWRWshirKFuwofjBoLA
ASRj4hH6HBh/aCmeKGMOhRy7laT48yf9CGz+qnML8n637jSVQj3ehfApJkyXrUQbXBHzTE5wd658
YYl2lMr5GMjp0vHNoi3YxqK2aPbDqL2wXwNkL/8ZLTk6JHEUMaULx7oOYHwDuREtnxhavXbZaUX3
TvcJ80JofX0/4PxdoJm2YTpH2Nie9B1sXRrRaLayQzPgl1KPfVar15ybO0ENZ6sZcXD7Y25TceFD
naRghDb+6jupuvDRBrAvax/prVNG25UBPv/UyMJPf5pe3trtrejlJ/YefgEGHIpC0b9b5+y33TQ4
r+g1hyqGbepJkFXha0pG1Ci9oMIltmijs3FI7UGsIqycCJEiJhVBIvwieSC0zQDr2QNM73AxetW/
IbBQ0v3WttjTfzSpnbdzrP+l/Pj0umqdZxr0pC9XX3giOL5O8r/kPdbplmXyDfol3e5/x26CfENe
FEkyYO68apQ0sQWIRo5lTByIrc87g8vu5eGBIXc5yRaKFAenjjHn38g/KpBpNejp3zIEWkaDT7l0
yfJe7oSk1MnMDbLmv4tRiCAcReqbXhEyXzMSmChVwkeTO/5IlyOyqN0VA9aObZZprMU/9RZOQZwa
gTQAZ4dXe51z0QbuEpfc+8pIUh9mJn7XgYbcqt6RenRohqDhT1/9ErqWgpo/YFWlMxLDfMYE9Kk5
dmLf81BwjBZkYvB7zxLSIpP455L0HGhEGZFFynWg/LJFqgPf/KA6zBUuEpnDu0VECkXDwFbDjvSl
O2Mk6ImXi3WFcIl0TYoLz0ldO2x0Ta7xyjXKrIUoyUHpb1Ek8bSYRFKlxsWesPPkkrzZbdBRYArO
Qi1zfgqHrK4BFIEj0OxzTRKsVFV380reocWGnIfNfR5TrmBI4VTlX+AJxRmVc6s8/W+s4KoG7EyU
PLIiGkO8Zini0MPbhsLX1EIDoHYlDiPuJryisW6trxI0pyaXkb9umwszzKAV06Uv4uirDWJJzlCh
uYmGLgwTIwGXYszICDv3/5GLpLrE8qkGk6Ehc5jzntslXqCPDsuUobD+rW6teAM2z1B146sMka5c
6ODrxXgN3cqD+tXt86GGssVIJZ0A09e8sMfec6Mu1xNdvnHj095Cje9NJOleKxGt2jUr25d/+keZ
8+2xnKiKBIzlUYxYLfi5AqJIbYBNaDqiwcjyahaf8siD4vtlRO51Mm4Fu+tKKc6Tv+j1LtI2vKWE
mSveXUNn7KZ4w5oIylEvLmkQeIv73gS27iGC0ulQv60VynLLshCb14S0yzSTDceFfJrdaiWiBSxV
QADsfd0Z+ktdBhfDnO7TcmHcewzpfkzGqN9auoVS2S6NwAKYKmYUB68lOtUs+qaNAJB7ShTdBUJM
r8n55Z6hUat/21bbdPTb87j8/4JlRc9ymY+KLetj/y6twGl6gh+VZv4GSqOXogQIqV1kvKNq3apU
GH2H7wqDLl/bwwFZDmcmFGHCSo+/fI5Idm9ppwvcH3CqKD7KryQNQIl6Gqc8plc01LYewSXZdPKo
sIN0ILk5oRK1oIlUt+/2VcjrG4rpEGurZLotuMLicRyJr/xZjiyRwJe17DqhNJ4GWAcEu5dfHYp/
5v/PrqavTA/S8naIzAV2KOZTs09AkpS1vtSnDq5I9CM6fcCxsKN4L51oQp1zhmRcd+nu/ed2mtvf
ir8RczNTfAGCJ4KppTquHtdjnZH6dTylQ6ev6KHiEqjBaJuQNzkkbNisLMPxGjxYz7fo3onCX9FX
+salWqRUFh1kRzwy/G3/FQR24X353wZ6qgUwDYHX8V+4tBKz+eUts8YP/4PHz2WTJtm55kfPfh8q
FU/Tt9b4UDd1aepd2Nm8m5qoUMoYeeJT/lhAuLfBrZ8nIMjyX+AH1dJv2m1eXlKAxtglGXCVlOTy
unPHbWTdXbwdYhW1GF6EUmt0vv/owTIAuSfSB0JMSleWoaA4pNbpTARBtF3bJ270hWNwWNEzc7S8
rvWdEDjNTw+0tGoG7nvS+s7dQqGXu2QT6lW044XRoaYr/HKBzNQD6u2nzjfioBgxPeLZNvL8Kmf1
QQ1PVGw5zWlPdl7kGEqhaRvf+sPHa42vP7UAGpsBOiEjwTl0mPQowxFIVictyZTfeqbAaRJVYlHJ
3J2PS1ephY9kuxexJQCNAfF3YGhxvWVQmM/PhVJR0UPcTh2jG5JXb7CM9W0IWTyiHZ5L0HASCHN9
lLZqCPfHtWrdG3bFk1j8Rq2L7F3rLIgTobcXN2pXvqbgd85MAG5KjRzl9GCF93PACgYtLdAounRM
syUYVQq/p2lpjc74tPo/sUEVSTgEXUPjKEqr9DstPbEOFdSmgEylvaEEzx5meOqK9G4tm7vN2n9P
HHIjvRP3qThe2XSkjIdNE+Em5Q16a5erGsnT/ca7u95JlWACUXcyi5Lu6/ynL3Y7nkmkpZ4pW2bi
i17YeooEe5O9l1X/ZVTcSpAGQzXhtNMLOnlsNWVMobr7LwD0j7NVdUwR17e/rQ8JlWMEnOLlgrJy
KJjYIW6fFtPSVdK5BpHAz2daolQsymv+ZCO9GrCkomQeKvF0tR07pb2dUVWUlzF7F6pr6q9/jOQb
gFA+Le5gLvvJPox+sIBLzgi7WISoQ6JCR/jQxOjXdFAn85NsUhTzHAxCXZvsBrzdLABA/kCNr5C+
tl5lOy9KUZt3M+Ch14xFteML6UGFvUHcT1xFJ/gphzYmaeV54jL7OTvHix4XAybVlh2LpIDNQ5mM
gqNY3jYXRvgYC2dHcaJ3hJqruPIw2lKGVrn+zTplgmBUtQAL8G56DmCvwy53EsrQ7FxFjU4fbP7a
u8hlsJH3DdvIysOy0cGDVFnX9sMJBQZ8rcpRDxgRn6ADqXKZyb+DR706AWQt7OmzrD2JloMCGrv2
T9i7G34jQkaIzJSmgt5DMlTIRbZzK+7gsgNYwapWvWklh6G0TWktvkoj0hK3kSUp7b+KZCcNQfb2
SNIRGi1HkXc/iYT0/smYI+ZaVuPtJWNX7veUtIpHRenj4o9KSTL+ZV7d2H9JAE9zKgGS40EhpMST
igDrllxuZZ2/8+GA0ZR/viUT3tEMi7CZh2ay0R5ycAHrEVgkDks1NoqtAnPpT8VGB2pHJUbSM/y0
3Qo3QZyUaDGM7ZH7rNzqJc84tkAutXj2TH1wQIRUvbfzedGHCSzYCJdNOMgn2URqUv/QVGEw8Ku2
0EIEcCkJBXUo7J+WA9zsexxm77aU2TVXU5K5XtFYpXeXTz4QwJkOt2X19MFDGhlZNt6A/RM0ieXS
KIvLGkxuN1v5uMZCBPrlyEE2TS5Ksdk1N5R1KJP0zaBuQj0qzv14qsw+E6lPJYQpe6bojXtc4CS5
GVdRbbrWIxKjHV12HeiIvLGehbCfkQE3vMZ9jWH35V4lmhyzZ5HHbE0DSWdyR48tmmPCdYw14q2z
5Z4P0Bp+kzdtXkBJNbt3SEZ3FktC1agzLs89jigekhjzlsZOSbk//Syki7K4BnWXAaTXBdnbXXzw
yRdca9oy5g806MT0iLk3m5Upa+wr+WKNZwFxbiBfV1pJ1DsaiunDXZT5IF+v7xlNOGeYWqoWxu/i
hofUrJDYLd4CyLQc/DV88VTadMmUuR/dj7Wc/0QoC37fRtDeTtQD4/5O1w/bgthMkyg1dZxiwB2O
TGb0Yoy1YWMpcgdMpzwdgrkr7J29x9W10n1SYXY7XsaoAd96mCD+Ax9TDrbA4FyZSh5L5rPUouST
jEihzvZM9gUxjsoOCF4B34Sdz23DbNfBZzdqRg87MGIaVID6R9jIQoNJbrs8N9NlYrCpZuCJtDrk
Ry2QJg3IaHPEwa7d12oebmztGZKbqmvtYRnWXS3ui6C5wz+cWdwvjmCoLp/UsTZiST9eD2MwV1OV
mW4PY+H5tlUsjHL0dp+bhZl5w4v6MAhf8G5irdj/QRpt3MJzJd+Lg/xv6GTAAne0DN/UlGIr9E3+
UIM0fpGzPhutUH8koKZb8qSSoNVzQvYEt0iRWsIOUieI3z+atx401VOdarjMQwozj9IB2vQmnb+3
5wLHKcxZNMU2WbssfHUvNvuLnPbJLcPk6FqNiW/uCW3FYYDBXm/EfgABg5YrlSdsF+ETtlesWfyG
QaDPDqNGBZSPIR3wO/P8w00ZorfISz7R9/swoqCgQd547RSiBjNy2lJXr3k/1/+pp/qnVISDS+Oi
Mc4oMPaKMcBzk2YN8e47zT+uPxGGctsmhZAoP7Xc9xIraqZcl21CTdt6Mc/lrHr3YhuvC32+AQrJ
eE9VzTGKUD1oooQvZaRVhFGkaNqrepdbwsROBbpb8EXO4vCGZXwoVxG55p5aeY8Wq2PRI5IRiD0J
/LxK9vty4QXUBh0J4XOMNoRFW9/mRdpwhOkt5HQ8MSh7G8309mUhEknnfD3HOLLMz1P9XyyvxXn2
u9Q9u2WMT4gixhaPv6l7iyxifMlmzZ4TrMytXYdEYO3H1UayzfXDoMbgENCt3UjjQE8yQXaMs9Iy
D7HS28slkKaqyXzkXvnci148Bvdz5f88A+n8CedYXYlFGfwPBENs0Vafi1C3704F0Pbyr8xVfeNV
a4t/O+5NdFYJh0ww6x8wfXAXFBW9UZLJfEpf9tjRuo7YN9lIDYmMzDkG7sKGUNmLC38rVKu7oSEV
b3B+2E81rWU98LbFu46QTO0Nyues0DbxR8KQiZYmZS3H8JsBbHEpv/F53AdMYPERnPguMd2kn1ka
ZnmXpauvkYk6JFgVZKBGEhwtGVI6SUnVeNWRxxmQZUyG0ap+WtipsEaI9Q/FNHPmJBQCNygczXQj
oZPAbAT1EbuhVbsYwotK3X96G47NggFaFKStBsWbntkIbpondnw8HdUMW+f9kadDldI2G8Z2xyUb
R9wGzf9NVT+dOQ4tW4tJNseUAl0+eKBgjImbEqE6K2H2kcu/9S5VJ6gcCyxoq594U7revB7QPaZ+
jTOkASyvhNc3sVN1EinClUrU/kFWLHdB8l+Xg+mi00smvYqOMsIK3d+wH+B+jmNUoTBa8iP8Wfjv
9alZCmzn/eelUNBYab+AVRSlsmhudHLWHTseAiF0JwxeHa/unH/AG921fQEWlRMfeYIbpreuiq1o
BO204FIdYTyW9ynRSpxe/B2gqGIKyQ4fiAYhfkUAHdUd7xMT2adANJnDI/eYXdLGoLWkrWd45w6u
GxxYoM2GENtU/4eogEUOEC4o3thIcFEN51kc1ZPe01wI/kFuPanjTZmrboPHYl0RA3BvRaTF7pV/
fhbgLZmBqCJrV9QyueJxJuv6oyuEAa87zaNdRC+k5sSbfejs+gg8c1oFif4SOvXv0XEgwS+RBX79
+BNtZvY+5HcrlGBlJ3JKRil0OgGbwSMxCbd6unVnXiw8hV4UyzodeSgWbVCvhuFoO3hca9BsxG20
GRD/DsTDDDxnDfQ5RoRXQSyBU/8YcilXol8jhAGAlgCUeqXngyDUWcW4F113XhvUtdqtDU9e2aVd
gHsqs+if6PuvZJdTQfyl3c5Q9lNyD++exG0C43M42sVDn7EHZOrMlweMRRqdPFYiOwHMUbibnXGL
Rs6PVTmwDJeC3pOhdH6wKfx2bOQjyr8MzcUV1rvzgMSWKfmhBUguq2lrROgUgI3Q77eXTwztdfaz
05ceqzL1P8GZ7xi7MJYMnuptRFncvsXLCBkJSaAc/Kb5KdNmWrIZ+UyQmoep+XcIepffYebmQd5X
WeNxjZ22vNoDN3KNtPo6s1xibU2/Fpe22SEDhkZQb0MSiwZs8GLMVaHthQoX/MZ31dlIKPS1joa4
tJuBSIrYyJrUY7rAAW/L4O5iiMv3u9wDghEsDxIOsFXOZvHB6sm5ZOgpB9uYzdSFyPOJt/Rx/Wzm
J85sOqpW3mtPBimSD2756p9jO7Ex7OexHPJrQ4Kooe61ulrw6vdkFy1OSrUvH9ykP3zKcBZJ6bel
GseVrZVImdVPsRQe9Ml0VdkhEAp0MM8fJ6zWPJLMNCbdnROUBctm0T8ZEAqaegQT/6v4WPTDwkZm
DWm+j5x3KxhLCsOddPYu4fFlNvMhBZhQkzOxySeXo2NnJpsmW3QHDm5taw7iceTZBXWinOXoFuFS
QAc42Riz8gHVWtgC9aPwU+96XL7QotvdzOuxxYNtuItbedvn2XmXPJNrBXNkuSS4B+/YNu/v9yhP
139N+U1DyTPjym+KDzqnwwQ2QSpMg+/oopcdp2OEbDCU09nq+xCpG3Fkm5TSDdc/xw0xwVfOSYS9
qIyRu/lxsB/tcAtTNm1vxAoSxc7vi0WB9sOfIy4gDTIwIBGX7iQih0cGvPzJWUAE1vZj5KDBkEGN
D7Iho4GdMa+cLabyriokTpvKS7cp5Z+cg2kfBgqwvZtwi22pPtl9aRmi6desOar5i/DiFzozA6hf
Obo2YmT8Z6uJAfah2PFB66FrzSrqQY4hhzppMaiClUzzWB0lnmkU04po7F+6AoABQ4HuxTo4oegG
X1IzR5ce5zSQIrLeXE0ENO8/kJ2dbbB0aOJKmLZeUaEL4ndOt54DGDPS69keoJiVuNO2YOtMS+l5
vSkg61AALyn+fiXXetexm8dTchEi8YbahfsoS4UiaWH5eNd5H+1AZyeYkRItMPyoWk4mEXjqqvyq
utl0ClmQ/DH0sN0KuBumj+hviiJwoz+LXDdKGG2yL/NvPRokLC+4oTPfJiLeXF8v7B47kZAH2dNy
eOpYjvFdZZqurX9C6qu91pvRWfAv8xVHzs90CWQ4bbggjdWow7m+9vu82habyIwjVjk7MroFKrWJ
arDaH9hG7bLgIfZGIapRMWu/A4Lw1Jv+/zVK8qmRKLLa69rjVLL41HZFzZTmPzRju2IyuwVObN7a
XhFiiXwWto4EzYejEniEJe/6/BxKk/VTy19vi3YC0NH8LHK/WKIDbkoaSu9AEEJPt3YbjGUykdS9
v+GZIUlAncrWy6xjtdderPRVZpmEIPWNbECHD0PUy7QgwiuSbNAtkb8R44IcR7wVDDBpXF0XnX2A
9Ci8pYnl80F4LuULQmSv2g8Y3kyDYedhNj46EPw3qFQKdiWh1s2X4WX/0WXPHw/rPseqVUJpp5Qw
E8lVlU3zpaHnt6wxcV0lxH+Ww2gwei0rQqYgUaHO2LbZqAN5KTX4OSSj0B3pImFcHsz1HqT2BQNW
U9GKI+kLsm9MZ04tgUBIabal/w6My21WUWgjogUtOZC4kQNl315V9mEGB4NLsL18hNaiFElR1Bzl
Zq9ltDofpYffx9GyxyVPVEDw/QTs7D6CbujKCrxnbVLXpwto3EhJOwlJzp0qoLdMEhxUzUefP/qT
LPMTH2rv8bCGIqzUa/zcdJnKolhrharZdyEHGwtDVKPvUCEy3CRE64I2OugiLnc7ai1Xja5z7veS
d/PSpPsiUf6llpD/lmMF0K18lldWl9nIByadFHyDOgNRxuFsUqdJjOkbdxEcfaSDq/+BfRZjGhXK
h6AJeGbZIWlXD5Harmkytj5fC5LknYC1Wtbc0XEKEefCFrS5auxyd5tzQu6/+oDAwqRVlY2sP0tP
fef0mn6PqFol/J5T2TT8ar5Ou4RYSn+sHIS7n0fSDmh7Y61O322hMOWNxolGBVl8Cxk9wIH874Mo
HUvRmnDeg/XXG/cQlc/4Q8/IuVjVRki2lb6bwY+RPxEF9IRBMwFs63r1HL8tAlg4kHUKJRf2INAV
qGK7yuXBKe/8APor5T4fabF3LIqybvsANeQB0qSomlNWccubH7Qfr6MyrId0b6FZSFWV/AuG3oWu
fQWaIwPY5kMVfQvFeAgcvcyD1cE4z8JBznD1XWTXlf89FxfTPadtOLtCyt2Sp/F/08AX4qsXYlGW
pAC9nEjZ4UzNEZRHrK66oF4dRXAyWrHmzlL2QYcLuDbbVmwxeml2euwf64C8oRZ9tusZPdthkXN3
v0QGywgeJb2fKvKd/CqsoAf+UFdpgNgUXBROwp27/ZO5Mfn59nhqYOzoH1AuHjwlWoOKMcQGwRJ1
uDVh4cnxJf0A7SIWhSJ27sAdTQtdyaPftDTObnVsuqHwq6mKTx5WObPlDg88FS0+LUj6LoP4ccse
VQL3TgtSDu59bEe40VxNge0pTtvNxr9zM9bIZtJb4QGadRgjJbeOD1F8BGVUTb81BnqKahoCnW/+
hLt1hKmQuEozYJ9ZJ08iyTki+AcxeSZPXDoX1dQySHRzfUoY64XBVoymmVtqpnlXbcCh/WfiOjti
5a8h3xa8IL2nAdTiM134wroTtT9Twuikx7n7OK2ZNK3CxT4ZEOnqttXvA/hJHfJ2kb2rfCakAFTr
dGRdL6sZtvtsZiPfybXbddJVur37135kDhAMlQaPVqmg8K/VReW3G+jbHm9/IML5z1hEfvmhPECF
t3/21wpBHROEHW2tCQ9F9TzXYZCagde9ikaZRT/jsZjNuzwq5Y7nTIbhdXGxYH6S5vt5xvyRmRZk
UNdDLTKuBZdoGde4sfj94m3j/VGxwbS55ToJIDgEjwM3sx7bF3wZeBd7Zyw+FytXMpWfViy8hLz7
LyWxoqnT97eD3hhbMMtrk5HFqPiVWTkCMvcLdqUUKWnjnD0B2EJhXgoc4ue8NcxnKaf/c8wDOJUP
qKZnBccshLX7KKdd5sPvHbFa/NdZHYi2+oTccH1yugrpT7XsljiZQ+wJHLocU9rYZ/r+MO6summy
fAaBtZCriRSk6lHZnUUslGWsGQQGXK5Z2WzRi0vpEuRp3gd3n5q/zNnbQ6px1n3XAkj9cuI/1xUE
6c7u2M/+L0N4yKowUjYBOTYFXLJUfYBo86pw+mNgT14ibtDsAdUVa4cdE/9IcrPuVTsgi6V6Tayt
cnu6RjUWO8mIh3E+A7UBke7CwXWzC8SP28DAjTicWHWE4QjBj86haCdnlUrVfJjwopjZD07WE+O9
mVgEV7oBU8oEJiyDQ3aXlNxVdhdRZwdJKrO2zPCriYQQbuxUFrUHl3brQ4UMHx4ZOyIY2y2M9qK2
xsI2FEKR32K8QlHARrWeEmyrZL/8rSlPeLzJCA+6vBFcZnUQUYE1GRf9z9LVlr1nxOsCK8+iWPrQ
jzHLVjY7+wGS6cdIvxzauxw1CmeqoUc7Mrq1PtbvQbcteWAT/65BfzcSC7V20a8OV3CNP4eRUt9l
YPzcL/EXA0ncAZX3hJier5AkMASCavjzn8tpJRElP+MG58yxC0wJ2O7vTNZz3RiwPGpgLyvjYZ+Q
FVp6MuIOJKbm7Sgd/Beyn+NPUGjUyD8JI7kxg9V+5Ep/H1encggoX+MyeYTJdYRzjQPYHMCauByv
7EV8FlVfXEjH+3/N+JhJDvTma+xRrGFhcrUp9JIEPqRA0pvBoFuCCYV0DLaO2lEgX6mBhd4UKdKZ
5MiGaTJdm3LC2j/LQJmgLGFGyGlgs0VL4pZnVKbTkOyjWdGeCmMtQ3zpH2wjLeXqcx2IsDHXvj8F
sPqyc+F0rcqmxUPbbKecEfGEXgIIDMqoUX2WEp4Igkc7GXhi0jBpuXrVacrU8lVhc6PIhjtLfP1Q
A8kbcNNTwVBgwfOXNy79MYbxiA/aIA6cniDtggAZJ0QEoT/Ly+p4ZnBY77CrVplxcoYrKZ+vQz1/
vqYP6QGGgfx5ex1NoZBf+SrVqdRufplvOi/4VYndXarSw96NPPs7XB4I4ZwJIFw0OHoYC7SYmIBv
iWUUscl1uxvvuE2gab9U30SvAttJLnKgjVwpmDnwtlMW6BpKijRlkfjvfohfO5rxb0LIfKjVVk2K
LnJqj7BIUAdg/kcoesAHK6VG+xjZwmhjLOR3GWdCHKnRpMJ6JrogYAKm18OVonloV8wlHFIEXhB1
CPM58fjnq2wflo0fbd+EiCNiY6LbdI5UXwlzF4RzpAh+DaEQdsLEjegI9eT8GQLwwjdA/9/dhLTJ
0CeEq9iUC2cUO11meqaWgPtkMlsbHnpVENzv3fXso2oStJbrrM6miqwf5zdz1TBqRBsvo2dCR7F5
NdmUbhMNYuq5UTgH2FD2uz3VyldOAzTIYmrW+NzKg2nHcuH8pODC9i00B86XgwIMyo0FBf4S6psQ
ntBk8xlR/4sagALzq9dN73yx4aqgQ7H/z22/MV9rG3x1fkWkdBakG8d3AVCIXcz62GBbdhvfFEbX
umHsa3dsKBy2Zxzi+JUwHf9mnRwISPi81fUcZtpKQlz8zmk4BZeU0gno1IbdYE7OZGPkR2CsXdWB
HJX/lXvx3qei/+gRVWh5WIu90VdW/SLdw/cFouArl99nfEe+XYHaXmmpweL4PSEcHW3eEyq+1oEx
3f7Sj7yAsL4vCEl+edq2+6rocqQAGOdv6WythN1d5jrSF/j35RXKuoYvulBg68pKVaV0kCi7YoAs
Oqr94HsT6G8yVoUptgX+2f5oK7dGyGeXS1BUhFxTlwLHdE43zsCVVH963vm4nKUEzsyvsc6l0hHr
cn1ot6G/LbLNr0HygUEhO7F6RHfEG3PBYvxterrg7SnfJSiHY9oLhqdz28AWj2t2lhRkRIHrUuiR
KLiC6/IshdL9rDurSfWBlStTVsRht4yXZHD8MQlRqA71/kQjMaQo83TLa42hoAPmyJQBA0iUFS+M
PAnlIoG0f64sfYX53Z9cFg+ACFDM+ZV8j37nL8Q7wp2xXDvU5igFXTgH49/rXGjkqptoHVZb5mbj
/ClRbuTHA6OTbnVDIkMepz4VCHwilGMGRJFptuC6XqKR5Y3fJThJMoTbyMf2kxncFSg1LzDTXo3p
PzypzZLm81KHjxTmjukfWfPOb4bJPqAF8/94D+WPNOazJtA3n0432RxKTp4fY+oX6YGH3iKPp7nm
74fVl+M0U7ZaaAMjYVT8ubZbgDe5oZxHayBRWDgMW7G/FDKW/sQRE+Ur2TOV1qzoOTjhTwBMU+FM
myeq3SlavFs40KjOzUMS72dtCnYCBtv251vtkznmx2LZ3RMV/Uu96NM5bot7He5aQFaq9H2cCzFm
7iv35PUYRyNXJ2VRXX8bXVj/1/2ILcTvbNqT9Dn4hxKXJ44JHvZpCZN5cwSgMp2DbCqepIhfko9h
iCTtIYJP1JM7wcckuBB6j+jayMrHHm0lHJFqxJCMtgqbyuv8s+Z0KRBmC71G/bBga3wlFqMkz9EU
i/sz2EWlLPw7E1DsnmLJRiIuds/mXwwzMt+pxxl6hEpNoYl8Uem0bJcSgel9uaXSRfdtsp/gX7Ci
+Nx7gCCxqq0Se71gamDZjjK4STOKiPLrh+lXn/waPkEBXMjMTiDln2pAJk4Cz/IE9TMqz04NhDF7
1vSqdU0JPwzykOoI3hpN4sRx0bHFnkJJL9w9+77FJaKuZkFVd8nuJkxw8+VA4FLkDmzKiPbaDI4G
ImeFMmNPq0xTtIJOrW+jyewE0XfOd+GMmkHRQHiRfhMcsMazgXvyIF8cXoZUjo4IeqD8yzh2qTwL
LOPTMdDMpI6tYeCsEl9gPUIIv9XMp9Kir/om5tZBcsVhQ0FZztlNMvhp4v7Qm9MmPXE/5gFNnkIs
+NyG4jVeNgbqOZQNy6ejUs+1YfaK5uObdt4QS/4nBX9W20bFr7ZDfdzv5R2pY43LmjBm6MgELUle
NM9seMHCFTXtfw4RuZvYhafVY6NNx7cwbcSkvVdJVF3WgD/iZQgujVcurnzEFi0RSbI8lqZP0xj0
xhiGfFHNevyA2pHZl/AQ+3YPBTSBfhIo1jMnMkQAKdcq0YomNnGhtZNjBPWcia8znLosKeatt98C
QsuGA1KSLgf+jXjWKbfBl7Ia0o0KsDF5j4uMnuhk9kNIx6+3d5ianBSmPlyTJjezvlOQPS6V28Mx
cjvM32WzRVNKTYAUrVPi7V/OMfoDHP8/2RVEdtBBjLylvFXsBfWIIflWPSh8nAs6iPqBjaoUXESx
j8nNdpPUx0YigThPlarRZzzisqbdvMJ9cGFrjVzBwD2jCdQmtTFYZDByc/2461roHnWkw2kSjcOs
P5Bb/yhT+5beG7FZiesPeZAaUDZ0j5POH6fUyv+/TaJnjFK93D6O6xU1/aOI16ecZF7vVswgR7Fi
pO+E898+AbOInZGlw++Cr9xixUTd8jURrt7HYaTNpefF3Hq5qYlCTiqpJoJntD4E+80IlOObWcXn
msIs7HcFAEgs/mJK3SMii1Pz2NMhubu8KVOKMf6SMzn9EbAc0XhcL20jaMb0j9Q/mynoNcCkucCg
Q9cOupD7xnfD2efyWrtHsdXw28H2B/bqhhFpGRup0v3QKEUCES3d57IAqZu69Y6KQBxUioyalxgz
6WdQAV7bcmuraF9pZK0xwQQAd9w8xTE1jem1aEUzyYKqeJtB7vFxho6ro17NCkwu4+kTRiT/rKeb
7FWAleOHZaO0QoTM5ptI1dyhmhGiWOiamjqaRXrNNMs6M3Psxa5ul+mf2LQAr2CiCsssrlxT3FHe
YtiRXm5RjuEU3ORQcY5e3LW94YjzdcDHTAg8WDwva2t3RVx73pb4bIyU5W7N0JAtHPD51Q2r+hRe
uqAerLm0sYewilhnc/KxsxBvv62ga3W/kAoPB4waiD/tJvggQ6o2E/qWy5CC92N95w0Y8uNWohhg
IDRlr4GZTJJPfFuiJwMP4C7EhPB+mtO9w5cI3f9XJeBWHGFQF39DDrGDviQRG/UnY/IADfO7gx2C
Ulmp1sc02545cNGMZXqH9FHeq5DuGvxgCx70JiKsUNlN/tpvOSDNXTB1zGfvzujaUiUqBfqph9gV
TORT76/OChFjiBV51O9aIZx3Mv0WDaD/EKrtXtR2vruEsDePmo6GAfDRUCzbMJBz8Vds7FTp6pAX
1r6td7YHP4SBd8E4K3VeO8xe8Ld8fIYBeDoYMTkDGUthlkf0AYVqEVAkq9LJ3f2y8EnEO/4p/Fkj
XwwK2XSRH2Cl6OwoMWDP8qCRhG7FujxXOZjJof5USzER+pTW5DhcBZPE6R5tuFJQIcYMFWWsLjEO
keyRIMRL/SHdCvCC6jQv5nbSe6bycuVWXc3K1dL3+jvzooOflKlDe+uFy1Nad9tByF44/5zgCFyL
0kavYcuzbRTUU/jLSycQsQh8yyjTptfIVsyBjmQFsG1puqXLwUyUfAJEziSfgj84pBukA2UkJabl
KBpFgX/VaVNSbOIbAxOnVhObTOlJ0JnY951ON2jzPdOirC25tNjww/VmuX+h2il1x+h/gGLv4c4q
wY5j5IMlPUX6nsaans1PZU0ABHXQTavCcs12ULmRf7h+D1nXw45C+LwkBqEjYdp/tfzhzPt1dnU9
tK0J38y8DpLVZVrLaJgfiuNeI686rQWZc1kVhgdQNfM9uvvx1WyixvVQB1P1a2IVHp5EvwS468sP
ie6Ym+SVco+xG/Pxckpx0NjtY7Lw/OFQM1mklLxTXtGCb/dBs6ESfBYbA17C5oCn0vgOjyQOV7Jd
4Eyju/xz2axAVOc3evd2WgRivyb+xOWPP4HmYMu+DYpn8W9ghwtQzE7XtjQOWK7yDHhiprta/FQ/
ZEweFlAPUNDzAk5RMwJ/JF7gLak3MeegZ0Zjhx6RpD3OOTGumf3bJWJWzUkogc2mrKgKqMFn5uWj
FNmzEkaqRvRF4km4GDomPv5BqkcVXeKkOhDc9ODHUZq5mWnCIYVIy+rDV16xuTIbBjSTMzeHUwA9
2rIRaE3pTiGjbUvL/9yyuea6ZAXuRwfTqGeJ66eTfXuYu9fDlB9QSP+/ioWqQ4rpfbD6U2yS5ua9
Y/dTA73dRvvotaicNzK7FNx1xIbbOi+8C9b2zpju4gkAZFd1zf/8KF5cF9oyQ787xqv1GgDbjTVf
kNUO2ASnLf0ETlOmJAIcSwoTDsUMq3HPCQqpG2cODVa9aCuIMTXwjNlg5nTW4DpXOvMUbgNnYceK
mfpvfO7+RRchk51Ou9RnrDGZqKnmfb/1xjIYvQjyXpxWzoEyKPJTkDqL21+HgK0NJmOV8MDiVG6I
OmyKq7FbdcZNu3J6VSesINoo1nuKJ3lbZEIC07S/AcTCtQA8yybYhvPCrbfdhWdhiADAvCA5e2Z0
5Q7afXJy/0zi5DJiCXMV8t65yoIQLGDay6k1gomSrUL0a68WTc8fO3YdmhsJ2TEMh9UBs5+qNKF9
4ttKtQH4QS2qgvmPbieRFI2ZUFYsfve9TWf/v7bR9Mqzb+gYF60TXWihl2L0A9rbuyGWN62tAt/6
OI7lJEWaL3Tfn1Bo1+22rpNku4iBhNkUXhEsaCU2ZjX99pW7L/Xthy2XZtWFGzdgKzcC4VQ7mC2G
AwytLh4nCdkm/4jGE/yLeUeAHt2dku7kM7H1vDHzpm2bsxAukrntbS3LF7pTpGD46dm2OSHwVV5v
DP22dwro89/eE9pI1dgt9ntm1UwgstdhgRmrwY1C0LR+vX8ufyHls6yaAVCFcIXlWEBCwhZNDFjF
qujvWAF4XjCYSBenxlH4ZUxT97JtQKMamdfy0sEDfI3c/W70SLb8Rdd3Ec7ymHXgKPDa/0nSkXdt
m197TQOJc4eRea8W48YwZbjJz9p0MgEWHY/ryHMmeQbH8Okju4DMdgpURRQm0RZ6gIFObfdeMQQQ
pNXtrxYBuV6BFQl73hD+ewLoxld33NyrQGTFSr5LTcTBBaZxEjBlJo3eTkex++yE24aBt7FubC+T
etgVr2slcCVXDkYpOqGItOWv+Rp508NauBqbImijGqqA29MiM/Emp/VH6nv9TOGaSyhr8xn5sqp7
9/8zF6vSLCwXX87uROu7O6VBGXjsguLmLckUblFMP8+pdYfPX7LMwCdtrUg1DWPI4Ud9zqJjZ3tw
OrUoZeAhDr8hGOZiwFs9J92wmoYuMhiezHUPKD0nlHE5xvf2RNsJv6uro8o0vmWNudy4FOn/qFyo
Qs2Y2jv0h2YgVhEl+9HOKVDh1jYelvWJzzvLy6O3oiCxfzry2AfFsG6sJUa+Bul9ClKuekNhWx2p
qbiDa7YwrmwkADHBuUiOqWueqh7aLrp39g+0WB3GAtkNxlvWqvcEj+3RYcubAd/PN1E7nTNhJFRi
WmhXeWPoZiOfwucmruDUcJg5iAFTdZT3AQ6/MmegfSp3at/P0UivzvT8BAq4QXK7jPYQwpVC7dXO
1kwhqk8NaLatOhE9X5zhHwxgQMEbcS6CxWPgVxHVJYlJOH8jfj71JQ/SlaGJ2e7kfz9nbpro6EM+
toYM3tWsi5suldWCTc+HgReEg60M83a7qEF/3JDLYCUS/B3wkZRg2TF7kBRY7KCyr3uuX1QBEg82
8RJufsAB3ycaQ50lUwiKPrpd9dqQXmjJOKZ6UyghEpx2t/Vh7+8kYYN9iVirnVdajBs1xo1OffgD
Y1HeQQmUGayWNzDSlKJuKze8yL/imj5xZN3HLtGwhIgpoQRdSAoEr/JA+4m1O4mg+coXeUhUFCOK
ZhIwWLJGZYkVySmcGUVJEDrwFWPRLLt/foJhhDyiNMKIiNfNHorg2Oy/H+g4G46lsGJcPPz/4Bj1
UNUBw97lKJX914igqXN4amf6p2H/bfu3OxN3af32U1mn8pyut/KpGYZzcEVHPxaeW5rwrNBnq+NR
nUwBJBWpgCvb6t583CbcsUVC1/1AKJHx5Q2F4NcAYYQfz9K1/NIKMxzLJgct3gq7oumZorKIlKoj
MKEiUu2B54tTg+x9Ye8RCBF1GAfO41aEvQptf8K/sy//FU5tSmBLbSRfrVjq/zIMiR2bsxBi2BbS
75LOebPV2sw5tX3GSE5T+iaHvgYyflpz+iJsuIoDoFbwdFr/tAgZ9errHchyqU5VYZriRJUB+g49
j0YWgVgewWEin5xmJ+GcjPbq+Xe1LZClgQS49VZuEZUoVGri4g+OsGmNNOl718sUlZ6jRhP0mNYn
680WcbUjz2XOrN5lnNHaUYgL84DdG/W+uycp/GaC5tXKZTGXpKZQfDFgiEU3YMdcwrXDvRpPmMVq
Rrw16FIWk/XU6bKoKFbXfa2QRoN4pwKqY4Dgw5WzbPb8jAUppgfOPXlJbDzvTM8rsg5yfEJQmOpl
YmZgKnBFKtzkIkP9FAM3jpvBwEZdjOcZ4Ut7g4wvOnTkS2IrP2xmpDdvdNpInpBylSwn0sxPs8/t
qTTkWfgBZ6w8YhKrcbe87vcEUbpS2H4xshNBSIR5INlpiIhd6PfETHK/4eCHveQDj5YwRQyuNkg2
ll66XwghiLEDYfUinAX9BYBn9EENnS9ChyPRwmfzNihQ3b3WHJQGTtWzqAyELKKBgLfolZMQRmL3
Q08Uw/1jHfbM1+VXZS3ofDjwFZOxZUzx8sZz0PEi3hZuWeKI1vNsSKEvjbT5BvNlobA8Leps/bTr
m2gxrCutzY4/oYzO8CBv62jC5pxCLSJ6d0x01Q8ynMpuHMzIuCeXmTMiIDyAJLZkxkK/CHh447nZ
e5F3aHldzcUnE1xOkkPEAcQiyQdFGWOqDb2S/el20+Fm8Qu5XD0EBD7y37NwgMQTtYWn1kuvpdWF
C+fLPw1idAc71xIOlN2IHrW3pE8zluEYZrPIbdHtoS8C0HuNRrEZiFxt/jifXzxzWBNgLkHyk3dC
JdHRIAagACPSa4uq56ugUN3eEOpU6Va59xYTkGzcrYPiRYLMiNERpf3pU1OngTBJZIX0CjzYC1Bp
9aoELrjDRdw9lhGMalChXpDawGiSVxjEz7o3/4VHw95E1DhGC5YQRzmPqh2i82g/XooB8d0zNaJ3
2I4D1UAA+lf6s5u64+fjp/zDReykq2V6ortjz1kjHR951pbFnjh8ML6I66SBn4/FlsdtRXwNSE4I
Dtw9E9OpednZIhZoSNGpCRtm/wy6QOwNENtjNKaMD3jMNNUUGraD2ac4DzGe/hpzxdzCT865+ONo
NOOs5DaznvtzVowrAIeYS94UWNJ0r/nvkz4eP0CUH78F8BkAqWoNJP4sZN75VHux4D5UU9jeHa/R
zsMQeYZbZbDtDQxiTHTWwZL5jJXI+dBm+lyu6svjCdFJQVZ0we2KteTGCkR5RUEXRqNcuVhM1PQ7
0jxf0wiuECf2fjVUV43JVoQWlr4uwK7Fz26Xy9//2aTExf0o4rP3+67zqTZASFME9ND4EsoSI1yP
DJ07J1y6evmdunb36tnWKa18nZUISaihzh6w5OWLNmvU3+eD01WSvV7Q9VcyCdbP5HOtUEEciGko
AS5cFRg6BAcfFZAhv2TtO2qVUXulflndeZ3Z5JIanUdoOzYG/TK0tHUNYgSiflR1rjd+xmxBZzEq
CVAjkNWFVvPBd1p+yarITjf0mmqcsc5Mv/v/gr5DkGtMFwpBpH5t/K8vftxwV9IzeDNOEABLEWIZ
oujUHNYmh6w9R4GUeBNDilngAoDL5CzIOClUFpvtjluUdQraabPYzbtu9z92VY6i7nVVavdVK7aC
IFm+3JLeSx18pEM2UMwNtTZMZffAHmaJCYVI954+cyawgLYtFSEmC8KtleSwUgH18axu2lGeX1ek
uTPqK1BkAftZeltbw1xTT37KIXJxVwWfpd7lUv5jW89qVNiMGBEABpHzpgOfyER72ZCYtPNm5oJr
xVt8Qe7B2C2CSW0ECPwT6MBT9LmaIwtsCO5jJ8o6uiMCxc489tcQsTs1Cigtitpw7iVO6n2NYABg
boCv1meVQSTN8ThQz0DvavcKiQzSi7Yhq03hRRZV5fpK4lDNNm51OhQxEmTw36IZC/xVyLGvPbN6
KPOBjAMS+2d2rODev9Uk7tsMycTykqjMSbAWWS0Y18+BmGuX5m0AC8E/84qKcf6THbuO26fqB3Gi
q7pitY7DRBjMNqVRcO4TyqcCaiOclvyi2xN1VNp3Ow0J95ltmAIKkuKkLL2jTk9YZjqF8iW4gTkr
fK1TISOaDP8uJz299USUhvswGYPMpsEYZ3iHkDJW2uy3zRTcyBxtAeTW04u00G39OJ0reoIs6qia
A0rfSsCh6BPPFf6bZ83goqGJvuo+F1GOQWVTF6WadEIEweuHJj+lnjj0F6toP+a1gt3aw2AgUUhc
QuzgGD0kbJIBA58TBPCNiSNy+jPyozqiGfJtiNpywuy0s2zkfIjd1ubW9ND/C1jlW8AgjFga0uOF
AwvcKUV9ZRsuB/4mmX/oM8U81aPd9bhXshghdixX2D7izOOX0L14yWwDKkTdeCToIcNZpNzvKOca
yI2Gzuz5qEocnqvtdgCRI0DxktOlALbXvtU1HRW+OY+nVAdhSO5nhoZPgwt8OkLI1msqJ/DfkmHx
EW3o0wcoShVEjRiGO7ZU6iVkyG2sOAPERHkbg/yIKAxsuqARCLtKF11QbpidDJJyaerglu0bGJ6W
oY8Deb1FMUWEYtzNvE/3sk+Dgnu2vy7o3KBDBYljD1LmVs+AyNywCfumCp4BB/5zpmaEZmX7BnEk
3C60XqCR7/dk2vMau7xLBhlthhH9seLYiNBQXOWiuZNgHLoPB+dkspA8tuujzr9rhBYymL8+EU9U
zLdLpEJ2KPRYmRwb8GhifqEzwnV1mjfaxP4JajFvAiiri9wtL3GVlKUwKRKOv04HtECkVl2Axw7L
WTDXQgxEIwmYP5YtNk6QNir7tmpbggNdjL8nXYTccJrIArXOjjenwC7TnLhdUbzrpwwRRtuerhM3
biiUuZ6WsHrbZQqNlOMMNYYaBj7cJw78TXxFB7QQ7HKQEOqaZPELsUaDHxdOoTv7HkP/3SZLIYP+
td44ECXMguitZZAVj3xknlRzf0bub72VINBMqm0Xkpx9l90P5sZIPIlpREoPrTveqn/fN+QegU20
6a/DgehE9Tnyfwmzh7ZbpEq0ZskOvkKeFopYwyux+Ho9lD2+TZPuxF0D/GUpBR4x9fcokn4Ae/qu
28Tg0iMVyLC1St6YKezxeqYyFRd3qVz8nGCCwBSj+cJMLD8nrOb8xphtRRRlYwUznYw3lzRYONh2
pv03FvvoKcezKxpLVMWow/dTi9n4ah0Nix9eGm1a7VJfbIWoLqe0M9xsqK8qAyh9xIIS8Dy5NB3n
O4N6npp+Z9zZQxS1FyQlJmUv1Wkc+Q5JU/iyTuhw1JRvA11z8Kau5hLs6olKracx+s9iOglaEoM5
PEm56KtGfgQpspNUYQ2jWHdf3tsRrWJVxDubZtudK5rOrCAdJh4USUgzKsjHnnsOsu2r0zxALUAG
h3Beec9jtCoLkNX6y6GRtB5N+Q+kbr83Z1AhCIbmM94hPI9OLfRDbgooKFK+Qe9CiWP/FL3AJqoS
aizmXXaVzKzJhra8zx+ZCuTv2g7h1glFy+0kRuduWzO46tepMlZP137r4cCXp1QV/qADIJgNf9yw
0Ct3hw5D4bIqc1SwF5//WDPf2EnL77+peO4NaltAk6slPs5G6Q3tJ5/HkCtIejF/DJKLI9XiUKP5
tcFpz2qGIl6wKHJ7WhBT3TJzG8WmzGJhSAY7B4md53e6JmDoHeFc5QEtr6j6OZ3qQUrYF8cYYAT/
3Nz/yjjRgzY5Ct+iD/5DSQjlYYdeMLDuqdU0KkGg5q3hhQ4dSwfJAWSxk7CurpLGlA7r6HbEe+8G
g2PW11riEAq9tfjRzn24yKPVDY/IV7kq0MUnxQWOv30E79kQW/cSw053BBKgiBUmD7mhI2qK8FVK
C4Fken4AMmYznLYMvweiA3IYyiNqfSc5qMzi2wV8rm10o1CxIMDtXmiEoMniSf7R3LGDDTmr0/d9
Z0ckU6GAU0cZt5DtZxUNAYF3akeJ2qNhOV9hwdZFv7+HSXnVYaYJ0ElcxQIR/k01E8AtPWGDZtIA
O00H6aF4DvM/67iu8VEg63SkFqgJFYrIbxHv8XTdNHLgJ5FqKsGrufQMjfmpozF/On6+Q5ErCi/g
Yk7o+ZeKPPubAp32au5B6TaK/Kv39TmuePfYyFNty7wVsfDlav/2KPGTitwYUBoecpsWSJX5bjOr
nDINjwBMZfm59+rr35abCg0Gx3nEAictB705ZofhOxyaNGH6k1v1su0gOjEsaNlocPp8mB8wqh3s
t1wyk/7+ne2N/i0TIfJZMWHwDaNro3iBXbS4p+dcLjJHWJuF1P04RBCbniF8GOk1gJmZn+fXh+yj
t9asmmic0Zba+MricqdDLDNHXiT19gz/SGWR5sbUzU/kzq8dY+5LN6cbmCG0J1CjlBbnSWzGtutU
ZQTT8gJJYNJ5yY4Gmcnc89L2ttL6cew6IiemTUHFGO+EnJIDyubjOzfulyWFCU8iYrlBgEke1HSG
MdilH/1zBZWn3YABgl39imM8MXKeB5BEM+IAKjbUOAirFJc3v00Q9FAy0pNn+SUU03sh2iJpbejW
nMrg/SQn5nXFyWN8oZTMigzIwKJ2B0skyixzXn+qwLbuvwMk1VIg61l0u0cIFc0LuMsdVxwdFM1E
lQ2BViHUqe6aV+EI3dFZNyXQCnC22DRyjywu+nm9SGzKvh4ic1RZuMumncKYKTLT8qwbgruCaFUz
qQLBJunO36Zi2G3u3LE7Vk29ote2b+gRLMDWxiOaZUmcio0WWz4xwANiC5kL80iBDfJBDex1/16g
QWJIc5CYVqn2KX+bk+H1GKz7CEacZPu/jbzJCcS0NdUqu6KWbOhpVROFAkrwbSzn8qbJr1YnXHm4
KySGzoiOGVM0pxhE80uCq2j9CK0nzMOXqV8FH9oxeplH5pjXwGB94L5WG6GvNZWLua6lNyDnb76t
0+1vXr5ig7YfFtCGTaXUEDiiCgS5ulJ3tr2wzYmzz6umYKaXwC2xKezjbCyXc1ztC/uSlfuo/jWJ
WGgT9SLeuWT+G2FZhYQ7AkJBktYrCM6zsITFG0kSEY4BKvYE5o4XnhVX9oUwDblXIMUu/5QaSGy7
gPLcYriEnWZH6MQW4YUq1hG9eVUkQs7BSZ8lkM0R2hTFMZorj1dRayDvGRcgB7Qm6W+Tsz7BZ0tU
e3a8ZMaSi4RqovVvd8sQ8DE3dRHvLyVV6K4pLTuu4hH/aJaRsvlPmlqazHlCAO5VZDTc4SxbPkiY
c3YpDnEWt8RCpSMz15waixT7E46e8RauOH4T0Nczsg7pT9goQiftldqi7SqZMUbumbU2J9y18QT/
tzYmWOKLHO9Y725rJu80OTf3tNI1Ic/mHOSo4pMyutvWRu2pn2vsK4FzG+F7dJrQRx0B/VrNC6BJ
xCfpQmsyl4HfAkfClDckNn6o2OYtREeprjZ0G0nmva8xFoirzCK9erFpbkYVFfMK9BBzSuxcYDOw
kT1Tj5dGMal4ejRkQ9KIMfB8WOqrRWv3Bi0IRxEt+UzOkWvTQE/PAiLhvKvz1DBgwMWSs6D3RIS/
jxRfcFw1ZRtKtSQy6kl61XRAcsLocVI7LD3dVTJt7LnEU0z+vDJCEM3lfo39Pg2ZQgUy9btZhT3e
azlVklPWEv16j2aJSTCDzSbypfWQEz8kzWWpwhIBIDvTrdznemw+nsiovJ2AGJjtZ2qu5kkGPV+z
qlvosBgX0v/0Eiqx7c52dXR4Hk0MqrOuwv1AtpKB557fX+H74X7E/81I7WMqbxFJghcMVOzp9BUY
zI2nl+3DxViSHhnjRHkxXxWBc1F6zclENghPMpS3rI9ukhEFzhlymGNiitmPdYWJTFF7ATHlig+z
yXgb65Cw8okyyPvD80Yit366YB6P8Sc+PN1HeYwPe3SsRH/gJNJvwK7TcxIj3rkJ9XjMTdIs0G7J
EHxx5GvGH3n6sdKLa/fAMmv3kUmnhgH2wIL17SVmaz+mWP37wMqAySaXExsX+wM3Qzee6IEUZKXO
AEdx0CjHBnjyylF6Jun3aECZ2JGwFoGObXNGG5lI8OubN56eH0PeIbbyRlF2ofVDn1kWZ/zTGFos
Q2EAc3Vow0N/1shO8D9dhYqXfiFqm1zeGSKNsv3PhPfZrumnHZLwZ/DVShtNc0huRuOFOWMW+zsH
m8Bq/TSg15U0kHCJzfNnmKdL0lqJ8QB4qT8zBztWgYgw4rTUX+jwqxxYj8hQYalPgQ6k/RZlbSe+
C5SHyheM9hEGADsSE0jcv2gETPF53JroMZz9g/DM1uE8vaK0Wi1DFmqfuwLHNQ+7wqDwmquTSr83
SPI7WgkOU3//kyZ0Rbt0dTxH98kcnKaAK/h3bNbldGVpDiOgbVcXTpUJ6h2OFSGy084+Uh/Xz9uu
/j9lRfWEtuRFPq2f8EOr8pmHJMG1oAbh1tNKuJ8C2jlvw7YuJL0CnMWU9qx6LEBf3b4C+r76gyX3
QblJmbfbGwjcjsq9I+jKLudOj4f/hpRXb3KojWfVvMIQkHiazmLoVNTVNuwITYp1Ec3TYnlQ7UYQ
Gm+PH8OUYYN9yR4pbCDOGPA48QqeLj897nSE9r1n+lR81PtDIF1x7SyWPojOqn2Jhm2bDEdBvQUz
NxqRV7xlmyf+679jD/NG19TW8PYOeKGfAvhUYaUAw31/v52y0CIzNsVzO5pJcRoxRgzkcP/F8qFp
w7G3/lTEh2qxBilIhQNpXOQC3u3171pGrRSJJK2oI+qFf/WWtonmi3A7ngTyGdTQMTNaCjkMmQVQ
W/x9dpjNP7e3RGH02deA46xwKVD8e3Xl0Pk2KMpNoB8vNQNoxz/VsNBs6Oo3LgN0WnS9d/kDQUcB
i8gqq1xiEeFQl6HJV4s4Yd9LfKpdaAbU66gpyQolg480LeEwtiPihxLMGm+B91GNeZ+a9I6iOXcS
YSPtdf2hAW7o/jjVLYZzjkTbdUKdrBf6AcjeINer4F7/OXUSL8wjXu3kgxdLKHEPjnx74GueY/xI
oF/OVEcycx3MW1Yh2Gy6IWgDwbTPsfiGUJuoeBMfiBMV0b0cgj/kDuFWvWfRtO1uvQH8cuHOd+Ze
qKr5jnybj1Ls24iTeJPzhUr5vA8hTEvcD3zixWlal43EI2meFo1A8yGyelGX+p1z/kg66uC3Gu6k
tetCvV5VI3PqB00y3t36ZGmlQoE4nGYapgtmZnnvFaLwuFpgKrTYQi/fDIB15Q060O4QtgtFm9Ac
QCo9O5KC6iXgjf1hTHy4u0tuxmzlEXuOQiqPyXm2J64gGfuCZhpK2YzlvLwXMgk2M0rW0jJrKw7U
fZSBeFk2ELbq1hjqoig8oz+WTHHkbVQSXQW+H6MUK5HT1HpxT32bpOwsT+0CR3is9BGMDpcnSfbm
Ho7olkg5x4fx3Th4Z9GhEO2uIBpIiT6rTa/r3Fcq3liqwbxL/+70taF8Jr7HnpPhQ4RzCZ+DDlge
KGWs5MRprhAaIorSidj/PQCYI1voxr++BhzBkH6VvhdKC2KVmJVTtXZ0Hm9yYHUG+0BZYDASt1px
fq0CdnT3o/kDuRZQtRERkMp9W3U2Ly0qmWqsBILUmvyhtc3LlXTjeblCKfPQ5GK+x1dGJ7E61Jpz
UFJ8hdOV3dUwUMnG9n/1Wv4ZsfgCWpCV2GfLMsw03kuvVhzwqGjCautgC8o6vJHm5c3FOWwRcjaS
uXEY37tiKxFTYOBZ5CUWt0L7lDvicitZHkTpz4sNOEieZaOX7EXlKOdlTehWSom6eJOO+fytGid7
wEMct9p6eJaJfDVwyHCAcNUWRh385/68Ks5aViXAoeOfOHbYl+xyn6ozSqUNe13xUqJR2QeqpVDh
P05D8fvgF6kms97HuKjwzjcQ4Z6yekaSY25YKXTZF7vwDVWgbBQW39vy2XAnCYIu5VTXACFtfDWe
LA9Eu2i6iQMBSzG/UvUduXww9reMrY6w/E074vKDSib0r0I6brW05doRX3X0EPk/Q0siBMtQEKOt
NtouTx4UMkvi6ZvrvFNqyZeU405WDHfqM0977gdcJ5P5IHCHGm4=
`pragma protect end_protected
