// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:50 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
VgjM7uE5KKpja909ZqxXKfYROBBwSZ5eZ/CJVQ88pa7ZuKDY7Ydl17b+X1pV/l4+
jGjiD4ftmfG1hwa2F4ZT+lStoG9AkCUub+5cXSzNa00IaYMT3XpVpswDMHNFlL6C
bxXlpcRj3gx0+pHuBViX+DCtd2XJo3Pid7HgTzRiUP4=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 6000)
oJUeyQ0Of8WxBwIGwZR7GOOhauyqIQbi2Ydtiy03iug/5zU2gVyUnCYfcF5AAbLa
TrdzAgUipFY9OedGZk5XWZKQUqYoThH/sVJdhXihFQ1ugNtFlBHhDdbDTD4++pxm
P1uV6rDX2QgwFZw9ntB3x1WZH0/xY9b/jmgCLKVJn9pP3oVq3fgOubAQhSTr349J
mYbA0IqcFxmp2mLSynA4KNfwwaJDtOBKDO3HVZybkiBtZ39yFWikpvRkb5mBZMj5
73lPOyYcWUkSSKY4pojlnSNWvtTpbUI+C2COZ5M3JKKZdwo54bxuaPOm3NZ/4TUg
tseCO22OaRDtXAIjKyWmvl3tRcEHN+oT5MQYrSXSfrh89WPwocfkEW7Q4x05W4vU
TL5ZMiba1CvK/t4L6pe+9A1ig8R8OLjeVIqoJWMl/yAnHl6H50/MsHT7YPsUX8Io
NlTuK03V2SwK5OJll0isOwFJPthHWb6+5s1234NJgQi7SBuYLXUYTf7dBq/+9tmh
2NK7bqekvuqIkTLQrvQMDfSzrG63zVa7VKzR8YyG1Zv5LTKDOBgoXUUqmPgpEW6I
TZTq9WNEPAIG98CmjVYby+Dw2Q5Uoz6adQxTGkf9/cKcycYP40Ry635aJkzVvRug
wCZXe2A1X8MRGS4HDN3V7xnmgIuTs2W3tc15ml1nQsyaIkoIEOs7shS4Hw+hasKC
7wZbDbU3GKcOIqDAk8N6E0gf8bzKo3b1Ourx4n8zNys8fB5CnpajgeB7kQoSub97
YU4Onjfyu3jvVU8j7m9HE2SzCXirSagsrwfZiK8G2+2TIJdexx4ieqi/nFqv1RzE
LDxqJ7U6O4Xl08O5R/q22Y3USsWz39fshwAy5AB7djnl/EMD6kqORljaC4d1b+pR
NaWJXod0SvTqI3HAs9PxVTxcKw3BAmt4do3r+8uYF2PLuokl0IEFq5XYujIlL/4E
45hOfkhotMAVHlfDYnLcoS7p/+g+SA1ihU2+oulrMDqhXM2hBu0juXfbvr7bOzDV
q3JfGtHtkJhXt5R1fyPOBlm2qMWt4ItTahcJn2+d5T4I54yp0Ry1VldvGE1M3V4F
0oHoXS3PT5gE/uX48D6CCIKtFQowJsFp1HR8erYiwDtlZgtoqy5F+ZI7kfhmHBVP
mrQaIERysu+eT4bhc1Lh5PExv+3imFoRvpyeJPGq7xtXAK5REtTr4YkaIbTfbf79
IMW+MOKI1GqmSSd+0bbBha69xHnU/XYfRLLMdXqlmEZ23X0yaDGEfw6gFghwipAy
bvwOd/dTzBLIZXL80rf823D8CsRe/DKbjjeGZXbDvdiOz4g3Ri7B0F/HfilG97HS
vYhDLp9B5g69upo5d/cWjwegpZSdrhgrYjePjO7fluNY9xseH+N1L3d1lmERgQZ+
CS25yXKpxH8tK6ICDIJRNFx4EUBzdK9GaW7IICpyhp0d4fh+x4EE2NT4gyfAX3Et
oXx030nbQvZhxrM4oimp1RXpUZwj5c7qyGrbW6sSC8p8rCu3RzfEmLVZN3f+XL48
56L2Pbc78nYhvWbRBGXHpW7fBroXW5nNh/AjI8TW8TpN8KuYqKn6Cltsi+H+CHwB
0oxxhYBGfJVZhKpLHriJRE4jSy6kKJsrC1me9vmFSmOJG1Rcvk8ncDYrpBuVnxMW
EWlJhqnWRIZdM2o6GF7ChenbXoPqzHM2M+qgjMgPwmT5hDTBkO4SSY4k0cHjOURx
4wgMa38umcPH/zT6klPkZ4lepBsrkj+zb1rLIp/YLauJm/inyB53cvzvZ1MPDVgY
O4j/XlcLox5CLiSzoFMSDtucMZr1FuOoxvtojUmfnEmgXih3ZLGrGE9BeYN4QoRK
96iZOUM+r6C3/bBkLp/5MFa1EHlMbVpTGig00Xn+3TUQ0OLR/606ynbFCdEnmYXy
KOO+a4zRy1S0gKtfHInWAO09MxaZ7mp7T6oj7ADnYcpJNnrrIfV4bRnAzKH8TRn1
NHvVLgQV6NtFIFnI0MDqgO/1ylK052VmOneG9SP2M5rlBgwSUJXIH4mkt/AocXWY
KTp6WyBiLM1IwzgQ/119PuCDSYrAlAXhLJo/le2icVv6AADFZ65UvR3v80htYdIZ
NI3eMj3wxdRTgTzw09xnNKWnZl9+QzwIpWef8yoVlGo8wp7O+frY2n/FAPyVhoCl
z8gi+MwHEEkh34MBOfWidqYbGXfbjvsS/6WLX2Au80TkUnBoFGQyKRvggxE84e2b
isX2PH9pDrfUsOjV4viUGKW8nSEZw7xbqrGjNhvjPx/r+KTjMax52+TRcI4Agq7d
dWrQ+DPTwv3Ah8h496O1TllyUDynzQdMqZHkfL/6V6tpZApz3PkC/1sMWqZaZJAX
nOLJZm/fD6V+C8nknVU/VofkW2KcKQsIjN8FOvCH4NpC4A3iQPpfLED4x4+9hKt2
K+f2Hrhv7FyXlrTOrOcozXqd3zNVdEQ2JhTUuBw/9YinBuM5SlLgbit23mZ1jJXI
eliDGdaKJXkoNw+TW41w9LUZ+HaJ0f+VNvja5ZNRfkmWvJ0W5ShwOBwi8moQj2UW
qvSmp514em8ibWyzLADSYEPtBUOv8pgiPeKMGaaYy2W8cMz5b7iKWxXOL9qln9Xz
zRd3E6MDYTXn+UspnK/IQ7qPYug6wIzS47QG8FLx3z7m2noMBLIJRweQgCcdtkCY
Blna3/356k+H3R3LEiEH4YisdJ2lktyhFAlaecKVCTyCNsso8doB9LjnFNBBvD2A
Jz+2Zh6xh2fwV5K8E3W1SIyBgeCRpwZt04XnaBTAxa7qZJJlunN9qCmR7zFZhN7F
+0iCLkQrvOPxDcc1l6MfRT5D9pDpQRIxtnaGvucuudy/FHzxKQSpju9uPwlWnA9t
F8Gai75KDJvgHmIH84vO3dfYsYWcGH51odEpNDqDgmrcsWw2Fhjja/gft9ieKgrg
AGVQ7htZfpwx7/Na7/fGFn4RTXnbVzfR0xBP23GIN7/2+aKEkm8kYvAteM3CCE2P
2aqJ2v0q8qVWgnoj4MHBJAjftC4wJgVDcOvqdO1fl5ukSP2mJKMgMYYA1b8X9G2l
RHs4phZwjnA/e0WbUR6hjLGOdg9uYftYm3TC2XP4X1HxoH5kQvbppvVJ7WTeYZVm
PFC5E2mQgaZawalQWenV9tSAOtbFSI/ISkb7ZzC+xeLiEDPMflPLn7Rap+KOg1YT
iCexHKu16uEPr55iMbIQTU0iZth+6sOZmpOKPN64Bzhqo77iIrFAabbQCt+QtEku
a/oo4kGkBZKXNGFfLfveyNMIlcvQhVIzOdrHOnV1sZUt3bjylrkUIJrHHnfmC9Eg
73B0FFRmFCYgtnmeN6aAbiePQB+HDn0hUsxA/HGbQeetNZXm04H2dVtXCk14cEXw
+u964OxmE+/QyWKCdyII4ikFR81MICo1IWAq3iOHULTjZHuHsy/sWQ3Z8PxEpAIG
U7NYkxDzDciJNL7ytXdnu8Bfq6lCY4JHMln2rjUtXgjRTU3kyY3HaZiveb5ludls
nVyieElBO9JJSD5wp4A/WWuD+BLzBVjOGGRzXvmQ1FBp5ATIAkAzo1Ov8l+32slu
GpvwKspilsW/sfvR99IhlCPuqJ2oXDotIHs7oYEotBNu75taL9o35CRdigdfXKvQ
7QEgkq8UOP4J6nVo6yYliXZPDZNjhPeJtv88Fll/erdHiR4LrjpYD+kFKS8sdZcR
RVqPrMpBdqsGgvc1K0azaJvALJBT1SMeitYsy//5BL9Hc1VWV2+1fTb11onUmYj4
0QH5Wb61gyptD6P00aghNzC0d1tNVBjw6fbLRQK711+KQgeTZlZAmuU1jDGYyu5a
mrY52mCr1C+d8PN9QQR0VVBvZvEfH6I4xI+kecdHrjzHnWWrpyzxjKjLnuHqK6PR
kA2DJsdrb2+Hg9xnPyDPhtvjBx1wjAmo90myo+GWKpSOjV1BlsMNlg5LkDYYTr2K
+IVlFfyAS8rSRQo2L5VClWDhMFlfd5wzxGxk4s3LZH3ZYkql8nWCGudKOlOeAXLI
Ap7xmFtYeeAHqKuWIJufmTf/bW4V+K3Qi2BjOfKW54I+KD4bkJjA2qQlAZu19NSf
V2QGxi+e/5cEMoOs8Fe71zckw7PRuv7focp8O6woML2VtTOggPg/LdDhdC148o6B
f6eRhX1F3aGE6G+lF9p8UjIsaJrntzLjEYSSSAnOKwqe5ARA47aulG7RfsDZKeo6
cEf/r+o+cvIEEOID6bkimDaze5TiRgThxMdoL8sRtHb4kkgBbMPdTbrUaI7d96xr
V5ekFMQwMk3HDlrdBIAqOXIj46fZxWYilcGir5XdAX22/Ay2V9FGeRcobgKjkiWE
sn/2Zi/igIbvHsIhpg8BZvXXdhlrTw/hGF0w1T01j7VukuRKCOhOBW03FDvqjbtk
uYWXwD2JD8ihUviSMjeCiw/7h5iVxWHYyWqTPgPXg0GqmZ4+1X/Vuxw/viqbaZhg
pp1lytjbOjDy6ZtTFxZGQM8JleMvuXZNsl6lOyfVQBPnVCBF2vE1GV6JqTUZFYW4
CjCJAAtr0q4xOaeAX1RgtjTJTf+UWX9ewyIrbGxXd2OnwnBewIBxB4Ng3Beq7t7e
dCs6rGA5Tl5MCsNTKQWO0T3UTpHEVc1xhcPYK0F6NVsBq55iZLeFRfO5Gjw60EES
G1CfzDy+WUR6RKOjf5BgiNsGqZnVq31SrH49X/b+Jum7DuV5zMq/9CpOJWkmM3W6
oN2gwkGaMSCXT/zVI1aIsUZNmj0lKuwuYuvdq5DGGqFOaUqY+tvtcPHZwgrAguWd
qd1HHKJk/hOcljy99tC1/Qn7zt+nbmhXAKvAIJdDY9usTs6Q8YrQzlq2HgIIPQK8
L+4T4JtGix3famZQod9p7jKoDPbQHOOR7yFKYEZYBANRfZ6O1DCB97le4O/HSPV2
+MCaLtM90L4WVzdtn3Y9heNiWvUmPnixBKskf89nK/wjGXj7Qj6M36zPuBp+e/98
b4pt3CUH4e88UEqY9wY5OnhQhd3MBGe7Y9ikcfJZpoj65k0gGkpS13Fa58jDo2IR
1ZGnuGtlMIaGZOdD9XgIEtV+yD+tT5tnI4wQgkTjgeRCiIuX4gtBtzS86L2+m3He
fD/BaXy2mtFpGO6It2bd+ngZXj82dWdVtHLGDjDsxNHIPo9C5nDTmv7vKIpO+ElQ
w9LJKnGoh0uE+BMAsg1T/wDt6kstm95wQaDbOLnsLlHuT5p2UhtiYmu2FwB6Osll
7b5t7/7XPmj4LKn1LCcmTZrY4aN2r/oPCmMA/AaRaQlxmxtUWiDspI/eRi4ZejcQ
89Xg59EG3fF+yJ/WOSwfIVnW5SOyZorW4I635155P2Z02mzyh39WYU9L54zDsNiz
dEss95xzSib/35RNikVct+BTibFYoaLxbfzWB7c2bqTsP+KRoqq+/luWXb2Ynqo9
nwy9fAxfqvKrcC9/n2/LBjOxZjpbMYQVHucB3o32fSXZ8rz+fS198/RGz5/E03wG
fcZPx8ChPQdbvC06ZkybkG+ANMuxOkD9am2H9zH0tfpltl+uK0fbSuZiicjnXQgp
e69MKUjt8xUv8uO2v80QgkehdLAFkZtspaCkm2xlz2Ct0S3YJdkvu0FciogxAaSw
AoteOycmk0RpIKlcg+lMP23fOH2PIT+8kp270H+dGRxb36VU2reKPdlfOzG5MMOV
9k6zmIrywd6SWW+3w1HtOxUrWtCqDALgMJd5oeV93S8m+UEP/R8ZF9ZKpTsQTcZw
0bvD0Y2HefSt6R1PRc+/P/zNzkYKRlUwsvBqCBGpzmMc0kLnT16X4XGYvKLmu3W+
W7r9NUnjHzgZ7MRnmDf7F2GifElo3huXhdKvwQVMG91sWF2CVqfmcGYu3P9OmJJs
HGZWaYQAL8dPLM2f1M8jMexQa/p1Xu0SbiqHzHhGmkLiIVJHlWCq/ZBOhtt2otWw
gTH+jrLfnsQCYZ0kcU03D8QvwnVq3vIGc4zpGUqCYraWqURx7X5s9MahiPJxgEHk
Zcnu2gXzWGRRikz6jXgvVm5lm0ek7Dof76qI0NBM4wb+C4jRP1vLp8gzr3nvJqQn
+rwJ1wDwgDpxqdBk5fkVYknHR6r/dd3A2ODOZ8uNnCCTa3cwaooQAZ2D5YXWoR3W
JTNCCsLBHbvT5FiScljuyn+dlDLcuQWOkAkkzOSrJAy7fxxFRaZwWQUDBPbDj44v
F6cFkadxrIFdd/1WbLliPLJ4BIbBHdSksbDQLG/CuzpQta4+N/N8FvWfttXtlhOJ
0hjNnUKUMeNbq522+5s/jrEACp9AqWV/MOGO79FbCAdiQ1JJ1qSrxNBTR8W7uun8
viHJ6WMJBrRRcc9Rgqwc49uGAnDdWF9dPO0j3cpERxesTw3vSZnMbU7/kqzb0iYS
mKCKMQ5HyiVkmtgdvcYGQXzEla8nUYn119g5jfm33kKMdjH53zDFb8Ny2j6alE1L
TSGQRyrofONnw2oSZLTGrptqm7+KCqnNV/p5hboOr07JWio6G+Njg7PJS2m6z59o
dK1H7X0fkrpearzFFmooCY3QuF0ttihZnYkOTvxh9BkVbHg3C6D86zeKHHAWC6PT
W6rX1GvA/jBYzBYhfmAhFoSV+Ty9LflcxxUJnbX1KDDlmxBf7FUoaKwTMGstLn9R
/S0KWceEFUovx15ULuGY+2WRV1loHA27edj5do/QaS+gK+yvsKrIKkrxKG8FAiRm
Coe0VCmm96VDLiInzSPWbIDpqbXlxZdtlpa+3YuY58Z5ZPe1CtcAiH+uPOGn0lHO
8EyGjqaCsvyiR/JpjEEcEhO8ogziv8kAOe7iF4WU2S8j1RwNR4PriXfrSWluo1PA
KCp0IB3mXYaR0Kl2aVliNGwLzzwJ9T4RTaDq9bidUIdSN1xsht93sw0fAwcaMR+1
Rqh/2rrMv6INBSg8/OG04+G5hpUX2qLeBBkmozdgqlKp+j4M0Vefpbxj9kvPUCGJ
gvYj3Wgi8F4hrFLhNQe2vWjvm4cJmbjCRfKy2mMAEIfXDBtzzcRK59B0w7z1gr9B
OD7O6bD7hx4dTczgbl+H8cPCTBUaMxkqj+u9i8rcJTRM1lz+nPBXshh9LkO/CSqr
bJhcNXmhtCOpByv69VatuefZf2vKzKCsX2uQindoMDUBFmqUWdsc8yg5X9mQh7ia
eMgNtzxpwWy1upG/4/l7lw7Zpr2tgIcaYEW8g4bVG/MWjcXSMJK7FMTByrIPo5PR
HNVnpTCtydchHqX8mfJ922P2LGyXhDxMsQNHf4VFB0PUatytwjbp3fgFPChNICIQ
D9lTYcmkEVk1Cl2ayujncsrOODiH6irDiItDAgOufQSbMjRayCMruNXGZJXD+roy
Vh2MCu8WT+lWs/QCRQ7Hv9x/49zTdT/CYc8nauh8vQFXpkA9wzGTYEa1It6UHJdM
VxjSG43pVhKxCYcThkFWvF4IRho4y6n1aXCZAim3+sU2NAgOZkB/M/nzEzwee2Ej
IjHwBhLOCGKHWGMY9A9fKk2/MbL4Hlrwar6yFTTdy+uuOYoJRkRwi25MWuYr4XBc
wkq/wrNmGmwVhc24OuLvDb2A+gfZ8qaG458Rk/pIWqwl4lQIvTVK6DkWdhHCj1yw
7y8frGwEmohNf2ie3yIZ0+glWa4o4wiEN18QB4KbJegEanJGfGkvj/qI4dFTe18N
WrjrjNvOVGlq3sgob5dhZxl0+9VqE0jzaTwjZcAnY+kWtFo/qyLxLH110O5gdKzF
HInxvgQyzkHDzcGQK8hDhdkm0BttICKKpw0LkpeQXbVS8BjpQ8MTMUAr7+1ApvVf
R/Aym8nmzzdTNGzqPLtT1F904heRihpEWg22/Q9i2W+7Jo47CO4rMvFFrgYzRFEm
BXfrofR6Wv2Q3p1lEUugBDUHAWdnP2EpArW+wnH2Sefp2JrgQMX4adM6HFDL2H+P
aTD/S2kEPVjOJhI6cKZZv0+XUHYX/IFfnMFHzsKcRb9sS+E5uoGLENCtFJYjlKul
`pragma protect end_protected
