// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:35:41 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
E12zHERlze60ngeTxQDG3fsVdNyUfW6nrlLF9Z+qcQ2fQtqtw1PBeGKsjlJq08wE
LipdlaaK9djPiBioVJ/1KIEh5aPQ6w8oL7vUo7V6MRARoqDz+Y05oJ7eqplEGCLj
LC4FgwbRIDZwpZbhH5d4sOOSMWJa3U8bRObnD/tMb1A=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 7104)
P3Je6NaRCqNId/jmoBl2x3ODuAhmP4XhJ/LHViiERDsBxMb7MbhFWxxI/iiO2FMb
Vqrec8pFIk2rjsLsSsa2HX6sm2kY+g2umNn5ADcAzrkNC4c90eJvQRBv8LQ7N0J3
u0EPRhlSrk3hCM2zGpdTHKgN3cxUMu6jfBxtY5ZpHSSUjs8Gnhn9GED+kwjDbItP
0O9MfFh1YlOMARJSn1sA5AqYdQ6UaHyOULh24XKPvcIaFqgQnduFr0h/sdCnBQn6
bEWbZl3hQmA/2Vj0gOQDuMY6nup6HP2iS5KsvKWe0O86dNufaQqTB2tR9DkhOdgn
bTyxEnw52sK7P0zuSGhmw/hRvSI2YVFbAcJPI6BzVtBcRcXsr8FibV1LLD5054//
oNVSESykovE7N8CBlfz+6RlW4cjACvAqJTQ3HHszPrm+oT9DM9db7nyH/cVMXn+X
pDpCsLHbe8h7arDCwW40fA6YRD91rUO+PPtgAJch7jMF/vQg/wMQph/Q3BvX5kSy
d+nLCtpBN1FTuakyRIBXdhU2O5BaEd3+M6aTUHhNj4InPXEP596yhV1ZUf7F6tQx
auD7bJHmy/NDzQUbukaRYdgF/hza0pDHtMUVluDNQ2AV49Ydu2xxhDrKK1crPFlv
kraiOkyOQ73PeNWXaeXMTv2H5LxpA2xmv4de6X4AnDnYjxW657S3fPxGfQKfmAnn
Npl8zEtK9wjfJCv7H6ARPNJbXygQh0ReOA28wgc5CEOf41dE929PKy/kJZEyoat1
mI3qt+xVH9I2Ui8LrqaWsp18NAs5fI7TOy+cplGp4ayvY2A55gotlqUKlB6ROw6S
sp3skFmD0VNN1DIWAto+Q5t8QNvjwnx5lHUpWgOx5uN5MIgI61Q/HNIdKzcH9eRy
rSUqIWyXL4AcYYL2nhcvCeqhIP6tVKnLAp15vI6xsG0B4o91Uia385Tsywvq5ufa
Y1cVV/GOrbHobJRzKDS3qvf/dijSwG+Jy3nkK3RtY6d10vcEG5H6Uiu8cqHrZlh5
SixlpZdzEOIwTaPAuxnqBGhlJmLKoRQ7hq/oI7H0f3lCxb0+crD/MNTV2E+npZiN
Ngcsr52Lmy5gEpbhqNCv3re/tTpL9g+4OCMqalDgPd3rzl90BJfm50UiYONrPJwI
j4p+iVkLkiObgyP9i0xtnOCKoDmF6fni5u5MbioThPomCXWRJLX3D7xDxkGOB7BU
zih/FO05qG8mKrSZyEviVA1G64rdbdw/hnzyVzBYvBz/6MMVmoQln9ZIUZ2LzAyw
tak2YyjlykUPfYVEjv5JeOlyYDknKbH4sx7V9tKc0xKFLplIQZ4tCN9dtKgitA/x
pCRBGiMD408A7gQC9zYQydCG9CzS7KT67WaSLMWsWt0NK6ukPSJRIvYn1oiv1ck9
gkyElaWX9Lj23G1JfstclYnORWjzpt9QH+pBzJ6sYVXnBgDQy3MtLTcEGXIuKA1u
kz4mePFTgDIQYyViuM/Q0RJjKg/bF6/fIQ1j0emLGrWrFozpVS8LWW0MjO1DI7hc
Gk56lt/cHtyx5rycXtecziTckBa7LbrznNYqo1P0JOgpRT2q4gvWSdN22TQOwZZ+
9ZU/8hhcFehH3UB5+cLlVxKtYIX/FKTQ77PWCLQqiH1arQTQfKWTWNRFwXeaOGvR
u90T53wRkN3e78S+DEzWELFJ72xUK0oxTmOHk3YcfH5N/LVNjqM9eDAGe1wn2K7z
2V0X0PrsueR13cPzCem0Cu/p+fxtIDyD7nsJqbFVgdNdzFZw/sj8gA1AyMRYJzcA
1KmvBX2CNJwNblR10x5AGMW9QDInA3eOxYEe30Sbq984CHhOGpqEN8hLNz6zK1Ni
RAiJnRf29JN41/aONy+ooTEG8VLN4j99hlPJ3H6kn9lA/fYlenhRPBEYHd+KnCDM
9mIIdlYms6Jz+4uripCcIQtMIuj6EXEfnAeOz9E2LlARn9XLCJQoYfQGsJtWBkJk
EHFRksOxPKnkCCF2Cka6VIOY6gVfnCOisvGGgXWviaKN1P/BKCKqoQaycf+GMdJU
Zmko8YZ4ZNlhKIoP6VKuazVHij7yINYaE7D91nCpc4ZWrdD93ThdJ/BYjv64bJI8
lj2GXXTDXK12FwCXVWFvw9Narw3KVVsxNvxe9ZXMjh5z5g5/l8T7kL5xs/u2LTaS
kLe9U7pC4Ljsx3VHaN9swQUPGKyaZz9bIYml2aWbLel9gj2/wOrfqbWfYjjIDPFF
qW7KKxqfjvM4vi5KzOfua1qKEk4hJueOeJdSHT5sCm5zXSBeRQcbuOKpcBcyXUuf
YNUts0DaTQYmuZNREcKDKbCTTuCxJ89HID9RjsBL1oQCJZuS9VKbLT1bGzMVRBNp
ABIIt5qRREymV0nqqDAEEnOlC/IKH2LEUoMgyroBNhHdGKMEf22Q/8lcoTQR8hQH
9n5Uw43r6Bd48ZnaD6nGICHwvuXNQvkQdxR+bvsZN7XXDmaoXrwi9UXq4HnS3WKu
FIR9Pd1Yc3iGiyo8dCcoImQrGrx8TZzFwSiOjhMYQFk3MY3nH6R6V/BrnYZNs0Zu
NCE2htEfRPt4YTrrQT6cn0lauz6I4DEoB50IbLiPdjKci/qCRuQl58D+HD//Wc7+
fVCEnEZ3LhUpoB7GdjHqsmGHM16srPQpUh3DNDWQiqE4YJrced9M/lCeNP14xqb8
lb8m5PRwmwjLKQVasvykpCLLUfAwycjg93R0J9dMSVSh70tJPg+TiPTmVfcuCAXf
5s00zcEVk98IKR4sLjKaWhgGG3jxFSP9xv1a5f5gzpJi7AYUDWFCj0COGRJi9fpg
i6UTbvmZZASX+bjEsyI+C5q+7EMkjpYfBsDgRjrXIJzF5s3ceuBjUo05wlq6ThSO
RJtXiaZZm6MpggCNofP25yqwuEYkplKib4gcWzla4oi/IAWjytao4+heXV5UjOY/
NV7hLWTj60GNDUKG7CPDfZ21tQcT7aytA95ern1mrnxeUTFyjZTpJr/iB4mJPc2C
vqWwgj6HepgmLwN2vsYA6rlfL+nV5F9EbpJZKOqlWrRXLqiPiOi0XOMskBOz4FBe
CwuzpT8h7aL5DPo66bFV1uZhcvWUcYkXn4COUBggtn5YHuow6lN1TtscaFLwvCO9
73dLRG0h5BJL2AE8n25losiOhp0E+EOjI5EQfHnk5VswHk0IECH0c9q/gQDWy1aq
sqeFd9KjWx0KAU43i82OqRFszAF1nTFX4XhM1orw/amca3SK4VCks4Ws34bpHQmm
82SRW3vWDkqUxGqattcDIiBikhRqYun1omW8hUfF7qpZWxSr1FlHqeKDguNFqMyc
XD267G93SOMGxKfN8/cFonRAuEw+8Lzf+GqO2wHzmU1x3zgHDVaZqO1n+/AiYQYX
xlHcOaNMNIJtiGEcPCwL5N/yEHcrQU8VO7MR6o8V+B+Ij6KNRicZ5nD8BimXXw0m
/wyb+vqpwXzKGYC1jPdH5Pq/mlOJYPrenAZaGyAHm/IQIvdSeTQYN+kozlhe7nYK
QPnCLlR8J3l4/wEHXOhTKA7fF7g2W0R37PyHgH3YS2aox/oSGl4J1nyKUXKVfwOd
xQ0QY0e/VPxXo2KCq9lnJDFxoh85Fhq1SN8AWmR0Bjiyv/dGEQd0ZlLn8G27SusZ
4HelWnw5ClLK/2zN8Viz/R/okcuMLA8werKpm/Dw7NeertLaDzjApTSMvKw5So/D
ZlIUCWoBIUoeQbuR+f1WTyhaFnXl+hy8zwGHVTNjYBN60cIshsdQ5NFSbf0b1zCl
OUNZK1K8NXclMIhGMe1nzgy/O5BZ6hEYswPGhL3E7aPgY3A6viFYXU3JcP2LMzXT
4/0JGybEBXrUqyth/RDU/t+4qN3bvNCcCuHeGnLoCvu3dkMsvj7Hhcd3Jqi6cE2I
+5yHBzjcs/S4U1Eo2cEiTiy2SGTCwIBzoAVrttDX8GXmDLCdb1O+k/qdXJwqBjpr
7C7EEbRnXryClwlFKL9G7fK96owwW8ulPA8SsBx5gdy0GaFizTSWNJ99C0NPSodK
OfmPCZEtv9LVb0DwfGT630D/x0Dphe+9A76ZWPmQuM24/4mP8OdpvitcEXSnRzVk
RZE/qylCf/DUnEg71bC4i9CrLqp6IomsPY4HNSQ1i5Teix+oijHU3PC0vPn03HS3
LNtwFGixZ4kNWCFI7OG4t9tyWBikddbqYEJDQBF+uS06fPCgT1x78dGMFPz3kg5X
58UxUbIHLd8GY5kfz6n3DDn+ITdE6kd4+K1mIMWCKYqnggufGpnMury/SVgPsy+G
C7VGmPe4WLuQ5zex9SScQgNNcFRJqtNMoSmB9Os5VAmbRlUEPjdGvvB2Zswmhy8d
uUOpDr0QtrTkF60IiMLtXWlhlSzbrG09M1bfSAWi8G+O8Tc6s8k7hZW2a4dQbTrC
dmBwE1H1C4Murnh2FOjFGMxPEUOUTmCdQnJyBJBS8GoXV3uWHV8z3GbTUysNUbrZ
WiIt0Mda3qLfGYdNf5j9Yz5mrt+PN0k9g0YERLOYPAKvRyXMHPtiK5cjABS0bV9X
QkGviqtCCcNsdibRi5yBaSqd4pIwYKMRlF5BvuL0ILI9tvpgXizqN0r4PbgcaPxL
m2T6ckzJG7fq+qKTXD3vXWDZRp9VVU3A1lLqF7vDz+6colgn1LNOvt+vqVBww3ld
AonSABvgRQ4blM6AKAByhqFfjLEi+YQyf8UneScTajAMUVYeulLnc+vS83ks2bzr
xRfVOINYXtWy26lzAVK2PLUZHpvqS5inu8S6IMwHkZATQK/aqvzn7ovxT/oqfbc7
ixTmn275/5iYP0uVDHvqIQJk30ZWk54My+mkDwwqEzeP5oXelwwKtaJf3NFKoYkN
hwZHHUVIH+wvtw/fzJy6i1NwwaRTgUEfMbAZSUdRU+nYOdGI0uRe6k5Ms25m0NNG
DXWl8d6z0BXoqXIVs69ImXROOvP1Z5XaleuMXBEtTi4hu95/9ilOropK9adI0Wjt
BlrA2iK770zQwSc/n2iX/oUxBBRqIk1cNMZvauU52ObBXuyt9FI6zxUJ0z7uGtEN
THfoJ7CkGeJYwNks+ZFXdYU/yuL177OJ012CagnAvvMtn3PUhcd/lVtH1iy2Nkkk
rWtRxzpTT0+cFU+FsUNIRlU/p5LDIDiBPoFASZ2/ZvXbxyOPhVWm/3EYXvxzkCFV
mNNwtrOYIDWYfwuHpv4XnJOMl0qJt+1jIERy9dThK43ABhxGwOHuaiUInegHaIyW
MbLy0NGpSXOeQ7o62RXcfJNMKf/URR3/5/EfTD+SCmdeGJsoJjQqwXZ2KYDJMx33
jAf6Jsr0BtVyfza10OplswjcG7RPyPgQIL8HKW7XOCRvqXvyKh5mmgD6T4SSrFVV
xYBwAXsgXrZ3DPukJUe7wNkz7Iu7DIdAOAw8aAP9bt2isn4KuhN0avCjx+C5yLuL
HtQBh2UEm65PcVmhrsuAkwSUlFw0YJt9b7aIF81ZwuOmUuYummZqGIB4iHzOiBMg
BDAZefyOqv5Q6JcHxrh4TyWj309//ZaHJEmUkogqi7DwOvMYgv7aqE/QzJtpjaAH
Dn7RAfcNtzrEu9c2h7qBjUHY6fiel1lL+x+pGlVvV5BZZv4FL/A4amWZh43mE2gd
7H17ckKAj6TFIDz6evoNoxf51S4NgxXzfOQ5MBv0miHzViSkBbu+erCiRrYUlTKi
yltIxGSNpESepERvHfYRLqy5VhD89AwYaPHmIBZgZqFkxQ9seYUz6a0CCRIUxw/U
eO0CYVpeSxLUWPQB65EBJ83JVFixvPXWVCB2+SlNIAXLGOplSBxgnCrMC5Glht1s
gxeMejbf1hOzujgly9UeVRJcsdVD+AcwrJj7wLRRwfGMNj9yOldfvaCLSGBYUbF2
m1AXzrb0f/nC8PxwO/O6GqR6T59FjJz0gNVSktif9mQaxGkXT6IO/Tl6VjjujQ6B
5zyAqNggqnSG/IP1cmn124OGT0DTqJWSqjgCtki24QqHf8cEixb3kvfYLOmo+WgH
C/isN2HXhmBFqf0OW/TQZHEYyZ1pWd1BCpGzjkw0qfgNriK9ikV56oHNn6M2F1vM
He40bETvzwhfkVx6AVAh2DsITZ/KwmzumrpsI3Ez25mf7L4Q89KDe6BE8RWynSub
Vtr4gFucTubUFVeaWejaS9jHBisDkJdWwb1/++T0gtbZeVhVT0gon/ixPAHwHplR
vHUO4e0G8zeddHd6axuf6gxCiRIafAGwuEfbSFu549beibT8cmAHM3OTTC5pWmPT
HPFYkgs6pTK5pydqhtNYZ8+XuZoHoH+tBIwBlHY+FipUSNVJ+A4OXAc6iROzqhKy
pzOir/ewJrSrTnxeKRP9mW0z/C0A+8jV2U/p6CuPSBA9GcvevgmFoOBLxRlII4Rs
cpIyJUI/HVaTb8mq1EkSiSiQ/tUAvW89xlJ2+XSjSPqDz8Zqg9ergDUluMcu9oVh
Rad97vsUVfp/6SsN8QZ7M8fMsGuWn7tKA3YEoSg92LAIhsiJmoQWNCAbxc8YBXUc
WQ0erdXeN7YlY+hPUvRAwvMGWBn7tTj84L01brGb8xoctX2mOJI6qwaEwWCpkW6h
bfreggJaCiE7cWMeGiFxLCbM0TsvQa/+C/tZ3hsk9Mz7wcceBoQSG6m5xsg0mj7l
QRYe8HmjELJROego59q155i7RqME/VkIau/apINh4JGSjg8yMaE61oTyXE2emqil
LEKcWk8SisiR6KOdyNx8sfxSP19a35S4ry2PxkDAUUXL9EGgcTEVqYp/tGDNsQ9T
o6/g+RpbOZisdM5q80xFI7OQnElWf+iEzhOMDbwQas/SAX+ZmEIe5YeO/mVSp17A
3npDDFWCAEizypsJ4eHN1OG/61tTUmrYLUWx4qYvGE8GHSFsR+cPLKrS5fOKinw6
FwZ6qJJLYqNWxp03H04MDIfCmoyPHlrCT7dbtFsXhoIkRIpFLRSJFh26OImFX6NE
A+llsRg4INSMo1fzvpwH0ZkPMP3fPLxYN0jHtV9SOkx22Wb/GRLPcCLCaT/q8qgk
mS4bWSCX5HwOPlhLIZ232rmkEjqSBEVhz0C+uKtMiB7CZznRjWkHcrulNffcAHwP
PWmH5YzNLR1YqjYPPuyVZh4K+YiFdz+LF70rDrhtz6X2hwAyXKvE6Ar5Ip0x70Sg
EU2U5nEZA5rv+ZceyiSwOUm/oulOi5LO2IKsNhlsQcTpPbE36IiWCv5F8VNEW8EL
qIRStcSQHZX90fM3bHqDD7xHLRxAdJq6Ca8FgRII/MI3IVVZnxDBZ0RuCtr+shkl
pusKEriAg0BPWAjTNu4HdjugA48jD+TsgZ9LNVlP0kBVdrQbxuI4i7ocCOW7iPl5
vvP90Gmo+QwyOnfXRw+5GO3zhoM7pilmUvJp8KaGSpifthV2Ea1L6abPXaW9aadI
/OXqmdnCMa7kMmO5ECh7y16ojP8AR0mRIxF1MEI+uxQF6oSZ0C1OuaM3sWhRkQ4I
4Tkk1zgp80BlQLM+rLKKJeh78KS2RdVKu+HcLBwDxK4IoX1DYPyfVhAs+6W2L6DD
4cZRzxuwwoMSp+68CGjsn7NLoKJU5PIWnrVeBT8ViMMMBGHL3wnOuwaDF9tkFbBA
+5GOdO5goHSe2zZQIghBX/E+gEh64dzNSluIWjDl93meDtkDH4DPQiF+ZCrW4ygV
U1ONzweqZeXC1yeR7VfDzC0xJY+uGC0RupRHoUkHzfzZJGCyTbLioRa42q6BZc6g
E0Oek259SVAvbVLVwjN5PiNpS/dpqPorAGfQWGZMp1rQXINq6I+b9t1PlshQeltc
1i5fns7RC4ZT1Nl2RiTDcBVn6MaJs2ARSLt6HmmonzDLxcCFesWP7wl7zqWhUA+R
o62HjcrZXcpES7bjmzW0vGKrwzuaNHW3zyc3D2M84oda+suMuO9StTvtPWaG0nCq
YyIoV+U5O+WeJUX6BXoOMCewFZuWB3xJ+60/wTjlj0qKW0dtrNpjq0656bA6rl96
HMC86BonTmBrEivZKSw6XU7bbmbpZ5iJjLFrYt3rI7x6CmQl4+lt+IPqY3lNGDdA
Z/qEte12aph3Rf1P3SaV5TdVuiop4j7aPDIWZ3BMRwnRo2GiCFW2bsPP1cGorXwB
qWQ0d+FgPSab5tt5+3Y9SfIKQmU7ui/FmmI3XwJqZYOxljsrKIv0q/2s3MeMeoNP
fhRJfPkBBckq43jw3SBtQMwLbP5acOWVVolPUfHq/A1yjmFMMXzNsphTRRCqS8b3
B4caaP1qIln9TeML8deu8nIN2OCP6hRpohPsnPzvBksaJuAJeWQY5yvtloXNwSCC
RjxGa6MqrNgfkmP9L/8uNEb83VItPObL10ESpnUhQlBo8aybjWPxUlYN+KoJ9nE5
vVZzWP/IObhmV+7w7oO1j5j2KhJNqmcwI49ZnhWMWoL9aYxVm6RH5xUG6TEG4scz
rLa2c6QR/SixzQz92zBTzX52EmhvuTZzTV4Grh3wELKD/IR5U2H1tI+WOy0S5cIB
+MExxMZNY3p7aJBYcbWxGNl9c5ihnQ6R3d9iQfjR1ZOlKg6IQSqL0u+h28bO296R
L/VN61OwIJxLkeSdYk/gCaE4tWeHFhxq9PezpawfkuioVb1H09pX/0b/oTNvCzr8
F4a0yaamA+sTFhW4qMC33U9tQC2HXjT3L4EZ0UL5vcugmXMulyNA7Fq9ULKB7BQ5
lMf7XpRCfC9pnwQMkBixaHuAHWOqTahT90YC5WUzvbFnsB2cWO6rSkt5/r0cqqs+
F9p94UAUV2bVKdT6jk9YpTpiLZLstWPM/Gt11aJwjbT8zKDEii9zLJ+UXLnxCAUm
3L8E1WPMnE+1rwBBGkrWR8f2PTMn2lyGyENPyFkI9hFdaTRlOtnOSleOMRsq6ZDZ
UxKty5iL5H1YKs/d5b49NaxzqvDqpoomPTx7vPF+ZTrFQuCtqs0TuRmOd8XGP0Sq
kpuAwWakEI4Zu/Q7jVprw5+vmZ1cB2BhDVAYBPCmrifw2yrepqmd0XeQS6FAKCsZ
/FlHB1Mc1gt/4zZaxDYXRi1lx5bJ/yhT/cLx9M+VwFz/bJJ1pAJwcc/qgK/KEusk
2RuB7pUnGDQ2mhJqvDwbtVZjAVSaK+cFOQKOv5ABX7aMUOFlr6kzKx/3FuVmp2kR
v3YJZVD/9iSVJBSziAOPzvRxgaNevrAUrCltD91CAZK0KA/K06QSCGP+T7M4MCxO
IPxUNe6PTJnrs+k6+r57L4o2tH4WOUt54YWNytdj+M6RjINQ2pl4k/KcJ1WBHGTk
7mAVhB8lBHu+Op8ZDuAtra02Ez1+lcQO6+bYDxtq1mzRJR2/0jUFF2nmIYuTe018
rE4m5dC2RdPlvsXmNESpEtSlienZ0gLWAuYRp1E7tTkIhoHt2POJUdmQtBQMWTAN
N05274YApD9Bvy75yyCZhsyBVKv5UVE2S6jJzQa3Ebqz3W2SVm7N5Vhh9rjcRiCe
`pragma protect end_protected
