// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:37:41 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
LsfqAQdjErMQOTwFHrynN6yKc4/OSlcw1oCzPz9qRZOU/1pPdOxzprHGt/kqOF6E
dTy/ShiwbJXFPFphJ+eHMq8OKb1RF+gHkcsWK4zxqr10oE7w/GwsqNCkndrUtYwA
LywTGSSx4w8I8C22xKECGKOUA5R2P4eclyOHcsq0mPo=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 14080)
aMaH077olheJRTqvq0sPHNHNMuAr9uWPFiHD7XgqRY/Zt6keL12sLnAgTg5sdNTl
qVVgEuZYerSsBx6e0IIG3s1XwgZovfORxDzCoLRBVNMSQSMduv1z1KDqSk7+m5B5
I7KVKzPiUw7QLyNUE/0p2v/RP9elS6zgYz0BIGy2xmYehRO7Jd6D7u9zRw4uk+7G
Txy1MGcxLAm6jUBd42mVRgeqwVJK5FhtshxrICnH/e+ZU14OCRQURv77rjjXfdYa
U8zYKjYFrfbhXgTNGk1ew5bZ+GfLnQ2zCZAbLXxL4RAWwx0MFGbO92Dc/h8MkfIA
qt6n/eBeJ1wEqOoYond8aUdLwCy3YaHf/KENiHT6oKcDQxP7bEJ7KPS1VoINK4fq
6LBhR/LAi0TZDgimguX5TpIF14Yj23mbbIu2tTP0o8cm/WMQBoVsTonivzQA0zL4
ZYwVcVnNSe/fkd/NoX5sEllISCIJ8KKmXLQCvwkOTncENmE+jtu2+ZEAD1jbmPPO
VPUXCTK0yyr55phc0mrbvV+6FkAgr8E1CPt4WO3du9BFfYIR0ddaqb/rb/D39qud
D4fnDjl9eL30tpkvLbu77LWqnSaPFmj8VOhgi8Y0TI1janHaXVUErxYid4ysjFNQ
+9GHE8hCXsLQDxeS+AtpLF920SZtfGHwHZl84/HrLX6dBmuNXlnpa7hCn/LPM9BF
ORDV4kvg8efNhJ3563TUhbRXLPI99SijzfVXTvSxkg/Pn7UAQuAafxsID818yA/m
SZcPr510B/sc2BUMMHfsa5DlnzY2Roihe0Z3tEmTkFvThjpI8fzSpZQ9eBAbz/pF
+8MSfuuBS4eERJ/+qN/nmrf9JUDgQ+BNrekcgBB5LsulziurwnyHry7SBXagol6e
x+DURMnczv9HwZAXRzT+FdVKd/VBGJtHFDKBwyw10N4zC7qLqDkzK6FyKnAo5fsk
nL/rS1WSp38aehG93/eUVY4bNYsDGdrX9XThIX4TL86sd1bvNRe6klrNjBMeAwxa
BezZOUqFHvCkXHbd0BZf1kpS4agOU+SqgoRrdNNdgDbLjo+REzGd/ecwCIzG4p1M
G0ITZZoYwVwRoqPqNJ/Y490qDniV2du2VfQyMv27p6bSkGsttL5xBvokV84fjcZY
xwUPhML4kHur0yuHcThXaQ4my3Gp1oxF2E+kQz3DiHAjx0Zta18LUCgD3aw85jd2
JJ6WVbczxa0/kHxSU7cmDbBgDElJVP/qYqp3wcmBK9NusOhyuD4Oyw4XAzGx2kw/
JoC0ITW/ZpUTTy3bVLdj5g9hDgZiVa/LVJETpZBZzXpp7dcpygDfGEAoc/NtVXax
mFN0dMDbjI6LiKCryCUToZKpxE3/oN2eh/m8Bdq3AW+d5dusHkn6q9lEdAjACoxT
Xab3tNSRTsPIiX9bn36kvRP874j+aEJGToLrs+j+5CctsJva5G/BLR6JUrYw4ux+
a9V5Sw6F7ak7wGYJTvvsWUHvBsweDaMCDAxXLXNVWT8WYEPDbc2x/efwAlPU70zZ
g1L4o6kQiOd2jG666B2RCd3XLBeQdVmYwOtr7Dp4mQ023Sby3Te9mXKYEdblqOI/
T+HIUMQkmNzZ4D9P35ZB2Y2DlPvzV27JUaqfQW1Rb5+VfWXtJnzxfCE9335mLHwK
AKn9cwoiv+6jrx71vW+7We3+QJ0UPxFRXsaZs/FRb0ywdOOXmMGsUQVSckGQEy3T
OtrI5ucQ137BpM315oW4ltA35wu1DGsdrG8J7mkUvDa25AIWtIxDJQiJTKlBgxiY
EXVkzC4rJQjVuzSiwDAmVDGoEBqjmFxROBPlyWa6PP0YqlwgxiyYLqZMju+uvQ9Z
YcqGMXjR3Hi7U95I/e6ySTeI7uOeOJ1Mm/+n5l7PInaG/8wwaa177ThLv0x1Gpog
EpJeabnoQ8uqP7T24OqCOfIcS3XiqpnX79XQJ+sXJUWsIMN206qXNgZaRfRuKxw0
d2LXfvWL0LAocncKrdYbgu+mtd+HgjbimXVtAb5krW9gAlCVljN+TL1/Ocqrsnjr
3dHfod4ep7K31On5lpW2XFzf8VElvFHxE/vcF4FhRbwB6AJXtLjHN8O0JDphyufQ
4ggSmPq7cRWVBIYPocGE6M06PMOnbqQTgabMZ8fv53r4/rdFrz+xyjs6Nqbbe+mE
m+a3TzPEzmUnWQeKNLcyi9GBlAQ8mh/f9Idziy8XvIkbM6IvKlGvx5m779xRq7li
2s1BzeVb6rJMpK4pMEBEWsdgu8nmrUflf++eZ5GPZFJRHtos6J56N46kQVOABmyv
2b8qxQGy/6pUZP8Ivgxln11d+8mGRFtVAxHIRIGCDnRvPKIiaDWvG/lCccz0ZpIq
3GYq6ROR0G3+0cRJofS/orDeQWYepWGucYYmsgAVudx0CfRA8TWJzVy1mhBx3EM4
YM/wOjwZwaEjTIUIOpDqB/d7WUkHi4nKPRMn8ON8Z+MKqvIRYTtBi+z2lCSoE0Ji
lm9jZPtwzCMXoJ2k0SG8337/sHfGd5u/56whXTtFDjkKPhZOV4ffLQUFG9gF6heo
4PKD8AWgSrZ3gqYvFQc3po4Y6cKuuqYgqyIawvo4YtO0MzPtIoUiAjr8/jhrG+pl
11fu6Ov20k3JRFEX98raS/ft6a6ayAUL+SxVjXHJHxLW+KfOeMYlj9R30e0dADyh
MxzJ7xc1DF+DPn+MCY1iDrwAdUkB8HPOHWnn+/zW2yme2JjcRws3LpZup8qjqwkg
GGh0oMx5lUx9MTyd4LgOwvY61AvWcVPM+GBt45+mk8Hrzgk+wB9WsOuG1VU3Orzl
5SmkPg3sPQkGwZrllsWbXlqrmu2RsuU6sBNfyZxILRqsanlm5FbISeW86L9tdqGe
WRRlT73ai0cl0H5DcB42ZfIip5zGJ6zwpb4eETDeBDpI5HRzoDGgH7CMTP4kl+5x
dHKBumyLrM9tH22Obmw2Q5LvRXllVjLnnko5XqaZnZ/wpLsK9BsFDbEJZjowL67M
Zp5tZ/au/1+PEALwJBBGcxYshXaT8iGCiaV4U8m6acdMQkH0KsZm14CqnUR+m/tH
f2a5VVDw29p+xBXJisSFE0U58EDRttSryV98sPsLXJfPGkB15Vt7zPDhSHsT/Vmh
k/BtC06pTxT6oyVGVSO7pQETrSdURzlY8OSxoQkxwM7ZUINTGh5sl+A9RBsRCkzI
gD0wBrENCukbD3FAz9+rHq2pXL2NK4pyop6OIGADG7H2jNxD873YM5eulOCB772l
PJnjDa0NHqtYzOe/WA6mQRlpfpz8jP+xdmGM29fLLiqpc+1pXZRY6lUqmJVu7kQP
KDMcd5BIcuUG4VDJgO/t8migil4mEXQCHrBMBk27GUoJkbXuOXj1temFZsvDturK
iCS153EU/vNJ4xwb5RcYb5JhekmVN4yooYVMeeD4Hi6ou9+AN2/1zQIoZaFjy8b5
7xMerA1BgTqKqrp+uVWW/5d4VeR+817vh+0EIQ/5snNXGg8bszPernTd+ReDRkaM
0ZQl5D3aTnb7/nh1r9OLMmTpvZ4/qvJ//MEYs8LWq8/F6KuLIip4MuSRYUVMcL3K
6w5xKzXbUWhDmaDfBESWrVFGyrO3niv7RkMgVbQO+eup8dywk40/ZKGt4NcUWPGY
hCFieTLsZDyOapPrbG5XJFZDPUxTfZfOcWr9yp1mjE0ees/W5/zXkncyvDkqirAG
BL91bTCHUIStAkybaIUOHBq56VgMg9FrhRyxWy2iAPjA54uuIw0QDDHN/K2UQHTL
rLIgJWjV5m94LnnI/iY6APSzNIlCRCbyxUSACFGjUxbWRiiVbeInfJn9Vlg7gGXc
faaXTYuZh7Eg1C8pD56/7WPJzsfX38VYm2Kltjb/eYVEgaJiZLxNhBvkVD5Zhs8l
+HKgrAz2lMRj+1WWz0JA7hFZmo5tHe+4FhIeFXI6fUjMLR3fm6qCeb0go7E9JNZX
DkDy4aAOx7o5lA/5Dlhgjbo4Z8spoV+ni2IejgqZ3esAvFswmFkWEg5YJ9oHPHgH
avBanmIx1GDpURMn5PymIMjiB/txgSN/p/JxLv+2fjNS9DjaFlzKSWGLk9x5HYxV
nrlGBVB8Xs7F+FRfWpaqg/4YYTklwvgXfgSII48wrQXWM2YCQtVj0lHc6RMvDHmQ
tvUUHdS98LlmrD3jbCMfqJvU7/3LFKl6yq5W7he6H6EuGkKOHhVIJVsnR8hDriVb
1sjvGWY13uWnsaEROaP9/fEbmv8AdtvWJFk417RR36AS4ahv94iajgeXXSnFouQO
TmDo8QpB00AVKZ8knS5W2V9H8rz9L+cIV0uKoHkRqhKu6M3iYYsc3P6Q7Aky7aSS
LkgYxcNqDcJKwvxU4cS8212iFI2HsVMkaKVG19ab64hthhAhPOKUPRggOz7ko6gi
1yOY5IxyWH2vxmJZA7NeXaBrCSp7scOzo+qNyFxp3e6lCxLLjcC9K4nGyKx/k8y7
9RGmK4vy3ME+Fg8DEJZWFMk6FUZnVjTitplHXvSRYlq4JANLD8L93RT/jpastMJS
v111JdpUIjtTBTMiAEk1oHRyHgtz7Sc7KEQu6K+tbYRP4BO1espE6yRSsZXX3xFW
fVtuk5COzJ33stCOJQ9uyH6iFXERX9fqtqKoAko1MCZI/Qk/nL4oEdX6CC4EUO+l
aBRI42loLK/mLlLGNLnyC4w0cXGB1pT0XrrVldftLs+WzVaWNvGVIl9f6lYd3PrU
VOt9b+XdR9TUQg639OKwdROuqupvWz0b9G15vwf3eeWNRrVBSKdlcYHdMOM2b2WW
Xv3SZ/x8I3DeFaSJkVZpRchXtXFNcv0MCfALxehV7pRlb3jtGHMWgKTqKljvQuhf
ykPY6iP0ErQSXwdNKPJ6JmSR6MF+7BHwXGnKI3AajXRF4DpSia79qCqxQ9Ta3Jls
552SRV/OcocU4vaXChyB/yWmUv9/EYWiQONdtOPELhS2l32RaBdoz+Ienhee0gII
8/Bbkqym/BFEzzGu+7qCG9OYwGk3DhMgAZ2pv60JY05vJWj3kJ9kb2M4ffC6xGto
WIvdkQa/QXqfaAO+7353LpaLdWZilZj/MTM+/iGq4AS+5CospjsAkwDPiRD+rzYe
IAovf9ZCuOv9nCyegLf7z6+GLkZ6PCMKZJW5suBtrvSkULDLqt/zIvXWA2eFcjm/
N/4YDUVF9Db/rsDzmHGlpF3JaE6+wfGvmIxT+n79r7FecuHC66TUnHzS9V65lP6r
InvF0R8VIhtLSu4yjNY27kEXSpkuKvkFr5K2gIk4vN1lKPaBvimlJDGhA7tLNJS7
PavryRkzEsAkQ7/1KXS/hZlLiTPFP1adZLZmZlzT1ffTuBlGSmDEqOUAzGoEVU8i
ua/eIN8Tf06WI21UC1K1wOMbpsGVAgFjXw5wb4nP6QONwLxRAt4A/On++QBtptc+
88ajXFDemDx1ElSZg2wjB3y/nNiMeh6h7bxN8p94MNP3CoYu0YXoxA15MtaYjCP8
ZbBB58QWQq8ePruiL5L0Z7nqKEJIQScuJs9NdkRU/klJ+O/7waLkrs1gCykDNH3Y
07BP/oJIbfvgxdZXXSvBVH9QHzvEF5OWF6GFUxTLZS2xq3S3sT4cqfWszsPAltDa
V3ORNpRz5AJLput7qdsc1GR2m3eXNIzTApbkFgziMQRGu1xZejQzM1uqPM22e0Kg
dTGP8b1Sv49UHe3IiOZxownmyEfr8WOia9nMNbZoL+gESEWfnJ4YWH21hncPGh/Q
wcZ0RjKTJlmWr6k7eNv6VeY+y03OLUxRb5OsRMSwF2UWmWaaumKEAy6vpVEonRY6
bRxcKpnrBlfF1oKlXPMu3/RS9NpN3LmuJQofYlUYDckQhQiryWC+hvCR+SNUG+jL
vQFAEDeUpWLrMpK3d7nmy6zyJpSb/DIa5ueafJHR3onANChCucmTpV41TA/kPVTV
6Hsf0fiPVdsTZ1RnPHFaT4qF/Y0gCp0QhktickKCr9Nz41fP37ckCWkY+z+GIGvA
l5JuZe0+Ut8yrRtVN3AKvPSlUe1YgPkGi0SsKbTocnoDqoJMxRqcndQI8n7MVaiv
keMrYs6qOE0jluqWp8Qyq+HpchQsIDuDKUYn9oxABYZ2kyIizkGW80Ch+SqVNZwW
KZwlwiTepg0P2kqPqlEnt3QCfW/WmodcvYUg1JtnquKjg78Won6b5ntJC77w4GA0
lnHGUWfm1n1YJKCtrAfzDR8PoclYCYMdbmjZWJdsX9OA9WbbwTxVbbnTb2BozIIK
4PDpZmoeSB8uHRFHAUCVR83dkLDT0tdINoB3JFgU54qXsGoJj9byZaPpfS+2120z
vph9BJek88rxOAGVDqla8v9z1WEH74w1ybhEwdlphUpcLaZL2imFTGmPxA6W5hyQ
nv42OQ3o2ousMlt0YygkRDroYjtEyr+Ag+hSbY5U2z6iwnjZ/nvmKj262k+VQQu9
GqfXBxO5QG3I2xV2XUQAt2WMynS7EJ4jeRYOEPRma9uMvN6GunmNjmNYCeQ7WGoZ
oms74Z67fm6jbp0+6dUo7s/rJu4ksO61wIaOia2a8Vb3dEHCSqqlBlR9EcUCHu9o
dJpC3j02whZAxIWphEkFlzdAht00+UDAmPDTO9PcXdEW+jM5wQ8FJFjN50RoHcN0
jfhx6y53PbOvvVQG4ef9f8HLMtvls/AJPK2hLAMxj88Vf3ouR7jstlK5aGv8eJeA
0aX1zDgv5k7Dd8E2elE1xLl1eyEV6s+HJTEy/ccbfehiv1nBtFpuMusllDKQpI0V
w+7gij/Jid+nx+wfdn4DZ5BZtjGR2oD7bKBjFuvKOo6EPqIaVufVL5MFJJgn3kNa
d1NMBkM3YKc4Eo0ykWUgGfl6MxFWYQKP/TBVkNmqSS8biR+IPxnufbGwxKx3DdbV
JA6OOQmsk+0Qu7sc9u5zBiC7S2gXQSYsDHRN9wtOQHVSjlf61WzP+FK9PkoTW8oh
x+ot4+ZJ8jkd01Eqi93XfqffJaafvFj17GFL1NOZnB/deEcuM7C9wzpOXlr+2Lp2
JBzi5Q/rNVByjXa3CIR2ZS/O6LkA1IuS9j1VfJgx6bhW589uv4kFkGZXMsLgdcVn
mUeSm+3Ido2H/Cuf4t+pYbGAnLE/DXHrLkDXzqVvyS83GMbSs/L1DDZ8NlrGMn4R
w/umyP69XVZDEh6FBC9RiKZ8fpS+u8zrLW/u/P+LpMe7A+qJk5WwK5mHULnqXvbn
u0Z7Cbsg3cp1vEsNB5OWLZsRXSLnHalAeX7SVNVxk2PJbgLunxuNbw5R5UnLdHAL
ZT8auBfyLlUcG17FLGOudHeFLKPMlXaxF2P5Vf/assgC2H0C6f/W1XwYbLE433gW
ZArdLDIHrrEInP87X/gD6D4ObK+8huyOoaI8BENmlDDBFXms5VcUiKbBYtQ7gfGC
EKwWXa3RjIubBsVCriImOQ3dEBtLCy3cTKKxJjOaHIhjLZijQlUTIJQ6dm3nwRg+
rnlG1zgOgnBWbvHQwDDGoInSXEhHj05kPBMliDH4KDhfopxkDO8f727Psia/nDbI
S/LctAB+MaztQ3OXdIlm6El4noCZb4KF1WrQigqd5a8caqgsdLmk8275Ud9C8V88
suqGusGSs0cwI6npfvbe5Jhw06TAgnLEonCcmfVjFz+v8/ZVogdtTfQmB9bnUWiP
t2vCKj/ewZFJ0HRz0iEqbE2+ZfKEaf+yJgHJAsU+ISkt6TMNSvDmGz3UefYLuAO3
PrfuRvWvbTRflFmRQ4iLUzylVs+sD2S6RwgdO/EEaHWC6THBDBXHIl6Do09ha0/U
DdkGhmGvEQPYo1VSKEYutttwrmsJwiuT3iSx6UEdaES2J4Q+uUEfKLs+s53y9eSU
0lbn1ufg+4amRJub5AES+nm2KBS/N9OUchC0qSmMiZftuNaCgqFS3deju66RPXWf
cVKMaxFENzawavxOIMdCHb+MgtZuS2F3tV/zv90tfm8Qw+k4TQzO+GfMqU+GhPhu
07BFlNCLIKhynn6QTgMsnZkavbnVGLrP0KGKbDnc0Xq9VDWXUSgjuj/77L1tuksp
ITQNuXAy2MUookof+vlFwo/3rV1uDAnqOrVpOT1DNyvDWKbQyIfv8Yw42WPYL9Gj
SKOM2DtT9vDOribMQ5/23WPJgb8xlKJDzcmtmhzIn3TLPaNNYnrAsqaUH5DDrD5F
JHORBRrcsFU5AuMY1QVCv3+l+W05n3JhL+WLeO3M42kD5SlkCc7HJ78lv7qO3UG8
12oWWoaubm7knOmeOUhwsFekI3z/iDXghztJRYTOB5KU2Yn4AIIEn0Fp0HSOp5E6
CfGgLjtgw23Ma2EZSZoznfh7yLjARu1yD+1eP6bv9lDko34c04MNr3B8+PJhBox7
DO7AwQ9WU/+ROLFS2eE288YDw2gSdVsOxBOhQp43mrFQDudd5kTTCqicxGIlu9Wk
WGJfELZZW6OENblu4HZq+Cr+G8Az/OPN18j6/OZjn8NirNBJXazTfcrHeQ33rZHf
HVoqdNs4+JAi4iAcrALtYgbo+9vkM0j9nSlsNAR7DYoREYIEdN9O7Vpi8wjMjHbR
ht9bd90swtalOJmpZGjhSioGhqI7r3WecL4EF7K9lmJkMaFPGOAJ382Cp/rG4R+U
LLSZsRnhJ+qRHey2Iq2MJ7+UqQctmNYAcJO9vuhhf0t0dkCKaol5h6KgqVemFWLQ
48GJOWx8QDc9S3t1aGlvFpHJgC+2F+DjHNnCeiFVQqD2Cd0g8sSWyRw9XcLhI2YF
LjpCpw8LGLO4paPzWlhmRq5fWlt/tyihjaTFoUnbtlbCtW/WmrnCqVFYobk+zh3K
22H/CW5cTVwB45ZWSC9LWURD1y3TLApSr8iz2deTPWEdzrQPEvo1k29F2P3YJjBO
YCBnXfqaJgT3uLHT71yATVzpy9XK9R6EmpglmiKKOmEvXZOUBYEi4hIJ/BGD7OQW
tz1KWQ9UZX8NnoolUW52xUPya4MlFJbb4jDHvpz248U1EV7PhrgCn2s47oapVghO
OLD8d+M+ssJ0FSpkjVlcutU5VwLpXMuWSCRSSBCyXEN1sDwq/mERK1GeeTKIxyw+
AyoZKYEZ/41JauUpdm3P1Qe8qyFxMZhQ4Usm+5BAudpnySgHaZJZQ3RMHF2ikPA4
4U6xC+gb2inLp9GPLoxb7qtnfsOm43Iv5MNBvlkZ2kFgZ+q29Mn8g5k7n444Ra0u
/WXRgz4vT0FwS97bneKgW/TH9IPBJLDv9vgw8gLmpM2QUG2T0yXO9OEb6l/DoZ2N
5NA1WgQcqY0JA3e6LrUi43HxypkmStoYg7uZ0B4n8i0mP/1sd1eXD3AGXbruCLSU
f1LaB9Y2BE9vmIdFlJkaw9qwsFGKNRA23CmlRaXuOdThQDrssuEkCSCzsTS9oomk
O39VjSryenNb3GaLx0P2KoFUuMvUpWnYd5HlPtXX/fm9/G7OJV1XNCGjt9A9SjEg
1bl+MAQY0y6XNTGXgKgDeIZmgdsjm3xV6n3cXYEB2rAQuaRRteZmMu8d6sps3H0X
AbyX88Hrvt4iYkMLe2oTSI9K7RwT5uiBZ1dcwNld2BDbrWdBMt3x2tDtnEaL6EiN
/2juNkYbJQZ/6vDZebEkOcc+1BxFDVcobC6uiZait1yZXdmXVNGMpWDuw5NZCqYf
XAwa1SfZ60lDX6RU0QDQ4DnG3C6Y6Q1kCY2YAYa20v5YQzPr0UF0B65tePY0FMh7
WOp/tu8+b11hsFh+8HIUdCdtUP12N+Kh1oNo7fYSchg7CeVU33zOb6up/KIKlvhu
H7G95ySNDoRYBZFAmlApv+L/sfk2rE/O93Xz2qA8avdFccu3NMFviAMB6VdzQnY+
/46f/Nam0BkXqTNMkCvYry81h/24fdwZiZhszWXMGiRzY8FJ63vPFLhWonBNV21I
iSNJR2+c9CyIvliBkaC2rpWVes72Jr8lJwOgYA6H1qabalQ5e9qTLm2VKMphv0lU
q4czvb1NqoYYA/0TLOLlwX50dZe2LFeepa8KdQU1hxJMsLJatprWMP2ZxbsHWbgo
X4yxpgTaNaKUG0XeBfwzrhBT7gKmmlDeKyqQ2xNYSpAdShca6pruWniZWeEbD23H
b0FBHa3h3ZPWBi7fuAv8yuYDEc/wtdDD4PwtWsvxOU50DykVBkf4RHsADomw1x8c
OKRR8XU0zagtHxEpc3fHXffnHFsrl1p3K2wIj7jKr/ID6RLjulqtTKRhKa8ySh0R
rEgF9T7ZPDa+CGO0k4yQQMD7ElsCFu2I86a3ydjcELz4Gs4icQZ+jX275F5w2Lof
vqnO7kaCeqmGT+HzhYbxJsWasOWFG6tqTN+mGhYv9Tr7WPeHFezoMbDC6Na9PM13
fQeOfe+C9ZTlE3SilzuFvYwxWzXoVLkJdWhf7HMupOQ8giVTNGkuYpjrIXAiQhO9
VCU5LiamNnfVrpPHy918NeRFf39ufGsiZbM/TqUbbn5xJ79W66/M1p2zsyXUH5lW
RSSW/o0zMoE1ddMOaRzOrwi77DeT4Ag8Qg/xa8RspGInGW+mDx562zyjPDHa/KkY
EMrrg9OwKAVxNjBfVzw3y0MqVZ/dUA1f8fbKf+jhbcr9H1G6mJKuzFXsX+d4fOyy
ZnX5mTNxV0wOl9/KGqvO4mZ9QlPUAoY8bsDDNUuh88zmPnYL3xSyKijozmEucq1m
HjT/bSEDWLe4p8S8SahoZiskcBBWnHwjm2hezLFNoN/guDR75WkmukalGjL7GTQw
PCPe7jk5vGmfIqmHZs+4fhW411cSbZqHEKLImKmTQxpvNdarXLbFMfeI/y8Tbi9g
4RqVpUgIHDw2OsxtYLth8V7yG3Tu8QaVMHLOZIzmw3yXv+NceMaKM3fnKjn/wdjr
hrpoVmrIBgYph08o4qhiKbVjXy7YvBHuhcL/LGV6AWl7k01O/qLWZcZzFJrkANBS
Ofwp2tWT5qmVWGPYzlRhIKJeQQoLVu/rXD0We0MX7Awk2wyotrOaldIn9Z5m/i38
G9p6GhVKULQBxTE8t3u2098ii4DgItRxdf7GR8UzUw6Nh9rH62t6XFqbG/+4Dbqh
wR4M1JJYQ6iRhOYXG8y3k30LjB3KK1j7Jj/C94fIFbW9IuSLxlXsxh8021+nqNVo
WNoTzDWFCbz3tS6ep4mJMeZF3e3hXUL7FLPgREJhC1J+tc+aZ03tM4l5BpDfZ/SJ
Wajw89KsogNYBQZDNQEhvS+ZxCxta96+tX5b9Kl2AmP4zCR4fzAaJPbd26+aSW6d
HT94s5vUHejCCNtDmCSerThHq53SnB+iExykVkgo1MEGkNsqTzJT4UDtovVDrLv7
Msgfzj7Y7Tcm6MnPUf60hsdDQA6uNk7jy9dSu7foGavH5cD/7/rceHVD95lX5USx
lTAOWPqWwp3TnBK0Nz+zTLYcpl3lUFlNXgsk5EeXfwIXFpPvJJ/h9VFnhbK9VsB/
uWqxhipVh+K4nIZiIts8whFBwVBPphnnIS9FuIKC2ZYVNvzYepr/WGaaGSXrcrFH
5vodmK1D+YfWSO2iTK88e45gmn9eRn28QzBEmSuF3vyGONti2wH5T4hiOYtRrBBl
CCOWmeZtrK25Yg3L/Y1JJeJFEldjQGyYHDCRWSQmZvo5DrZYS0zmRUykT+nHa45f
UctQ4wtbIzvpM7zPpWv22DdeUshhGtHAW8tqbsqqvpmphxAll+e0USEzxHUagRMZ
z/HwGMvW10mj3jle+FAowcVj7nR9MD8qIAc8lZz5jWlJEZ5wAwkJDr9Mz4SYwDcb
A8EcZHScR0irMwPQ5kCJxTPBRyJRbXBgEhnrXZJhk59Y//HxL1e0czE94vlBmTZA
YiaQGPzA0iNwleyYQMuguhTdr+SIhBCyDhIbGei3bZJML6o3TjeSPMXjSjRkpNLK
mgJQ/4hxruGpINZa/4Fu2QouRugP8CnK04HpbSkUHek9kFhxaqFCIyUdlbLUGh0K
oTDLMX0Sx3lDtYbcEFsPxpXyEWgpv2pmcVY75uGy+R/mpyQ9RaJPoR2aR0Z0oXk1
YTVN4dd442WGQXIbQ+tf3S00mC3AMhqpUIx2zbjx6INWEd3AB3Gip2vIyfZ5feL4
1oC06dVD+XcMSr6IlvrKI51TgZFV8KM0JcPTAQDjxj2fNhZKsS1BavKrTO2gzQY5
/xykZLWES2yCEL5H8GneHNS9C02AoJZaBJGtpqiYum1Nlv4eAnDiA/8e2e0R4TM1
Id/uSbfYB7ysCbdOKzYQtZ+46BA5CAgilW7vLTgbjgr0XyplE4lQ4Eig2ERC+d8/
g7mBbBdJV9KBoqQxGFMJua0oe5YUa1qnMyRlgXLQLNGXeprVLzgKJ9z1pvDNUrIZ
mTz49kBH9Wno/sxbUxJg3AxhmWwhUEYmtKgxj2EbLhhy48d2bkVsVSLIh/A/JpzU
KJsF3LwTP+EKQYcoMw/npJT/nBVdpplszehgAntzfC6/vk0eewHhY2OFSj+C1SJA
bYfAEr+apMIkxoyZoef6ygHFJlloqcKBtmWwaW2vEfpwYsC1CApyRy2YPJ1hSKri
PhWVR6Y5/iyLVs+YuZP8vWIrMbc7mAe8+IEmPzmJixwpf7JqUFgvmP3w6QRsD7Wu
gfXDIvjkaspbD+AKxhSjx/iIz3cmDATnCVzfm5mkDmWnDHr8TvxVLFPF6VAdcxDF
2J3hVZHEPeKpVnKhAfccIfdV2D9zaEdwVd++UXuNpbPg/fuvxbEv34j1yeUGq2II
sxuRLuWpZepNhr83K4obKFN+lqUCoWMzqZxtm0UaurMumMAZ6Gr2sC5Wu2fjxZBs
Uy1d7FA3vYh6n9zS2MHUsR0aYN7m9FWoysLXzIXizu5eY9IoFcOw8xj8krwu1mHQ
N21aWrKQtKIB228xpkLOKPTwU99UAPWc+5ULNXVT1JrTqFdEL6WAQNVVwxXXbpnf
sglpK2I5oMV97dlRONLuD9HGV0L4Bx1JrfKV9lATB03vcWZEcMWb/oYtZAzOBf0K
UTn1tCQnNYpcmC1FS5ckWOPXFADeObtKpgtLIDu2f2rBhgrgHV5dY7ZPXfu1RMfH
tPQDqBSuRx3Iz27fpB38a8EA62a/1Ez7DxtWHLqqvZptfjMxJ1MK0UWC196JCoKg
f3XFx/7pFLtZN36D/amcXXreuSxWRVi3WL1zKXzPZ045pX4v2eA8zrJmWjA0WMs9
BaaAbXqGgJ9QmikprX/Q2+Fc8Zye05eVYSoFngeBE0NYmJHeQgOovGjcBJ2zAU4B
Xb7RsNRo8HRQqKLRAv+QCJaVFEYoy0HlLS8O0mux6K+Ovh04zVt5rqCEd2iB7UUa
4VKsOYkeHatMI+fpq/q7yKI+IoP4p7lDPtxol+85oAxZ2oiNaGM3LiMstTRORFLw
0b/rnKEjYy/uFdpIfoGhAt2NqVbeNnzroxyt2zzDO092c/pP3TOdyDbbAxk4//Se
KYGXdpi8eBmB6+n97OXBqK9cs63tAfOSJ7ZrxOJX8cslpGQ6Zpk58R4/fHFH8dFg
uZ0P4CE6tQpPA9c+vkgs8I+8RrhERo/ivuaLwH4gtvTmnh1y6I8WkQFfPWmxNDVL
OzpLo32uCD4DKMZ07UCvXoPgi1sDc4gAitWDBC3YJw9LdYXczfUZS7vr4mzLG2LI
gbIaizshUEIYidCKyY85L7YwiidIthYtG0q+kaRZWKaS5xvQ5+VfWaC3y21T/TZm
X5O4vzOQmVKHEb45tQ1VhYI6dzd+NQeWtKBGJrIfinWkf+DWXGoJFhgyZLAQ7b+b
OyiDgTk+8KvgtzIttAMXrMIAfXAJii3gjg5MsPJjJnw1U/3HLcG79J91hefX106Y
+lFWxu2lstMcD+SoxXpn4TvZLEgdl5CttBo1ZpfPN1meQsKL17lyeG2b6snXVbwV
Gywya1cPKIBDwiY39C+urEIP+Q2EYPBt0sjqrrsIEU4NXZ19RXzLa3DG84HqawvM
YvsPdjDlL7+lOzxBxLxFtB/S/6IP3g5J8/9JfMNp4qUFpwaCwHFccwrGJjAap0Gr
AGPvYNEiDNpfUWpcPuKab38VOh0gXjIAHUjwA65GThj+QU5mZmLCStejP7zgwZQJ
YMuyH/Hq1z7+A9sbzRUyo+ZNP8fU+LE1/+MoSIMJFAGYqULmSC+3UV1HTKXnCgpv
KhOSHmLS9hZ5vV5U43TT7lOWswOvpLO40Z4NhdorKybt6v5wsNpiJ3CCVImqwlDl
FxxiAS4N9omZZOQIE8CBXeci8wkPWa1xoN0l2+7drmSBO50/6PmGGWnd0AP11F4b
olUvOZpHAcjZ1HRug6RvWL30fwTDdWbjJ+CjpKM8fh1cC5JXDUakFKCFlAX3PYo/
Inn575Am00A8PYFovf2OiqsgyitnFlSylP8RQIqisfxkOYWId7RMgXSHibfE5qUP
ynNOPXGWjW8OtEAW8w5LnM1te1+4PsC8eXGo9fuVnfigdLaku6DOm9vHge5HIFNa
cpUzJWNlxfhkwjrRPAMdfNhrGz9kTuHQZLH9N/Lr36nK57wSWTzNhTN03H5OjkmY
6QjlfxT0nxdfeNE8CmIH5kpvThryfXIdYgA8V/03R9GozFBIoNc2mXECMQ4tReNj
eZ+LfA+NrpozRgEIIBgf/A4XOG7+N7vdkkOCbp/VwUshjVCUX2df+AKOAj+o/DUx
fO/Tfz5Ir6CJLLMjcQNDtqM4AKXNF8rVCF56q1fJPJIHzFb84t3ZF+iWbOAcNrHd
POULwVQBZdz7VsGG4guf4tCew/47LdxEYJCfRtPafq1mtC6uZ0LLeTX905infj4B
DmetKl+/6dUxfm86rOIFjb3U6uzaMk06+LmAPM5QDB58J7s+U8QyhOlBI4RbIBsj
F6XQXmiExE8PKyB7/q3ogPQ8l9F2ouwjle8/OC9aL6xvcUxh65lg3OYuew7Gm2B/
f+kxr7J/3AbFF/QBfphuhN89G1z1csv8rigUI5fNaliHlXpoENnktvqTq0SQFzbk
hchoq2+HZEvdnAQY78YiH7tlbkpX4OxS96FP8kIAW1FmA/I2/s+D/yB0olJdcRtD
Jvuuzv//GJ/3JRyCJglBCD9qsC3SY4c5uRWG4ysD9tHZR/rEkiBp3mK+5Yl1eBOO
ovNv6+dRDP1cwvoqA6d+nQ7+88+qa6TbMbdx1XlbGo6Uk+oEvXCE6sutCXdO1VZF
M1ZsXSzap5vDjcWbNSXa81bXGJsOUCzSPMBRLbnkn40w3BSC8WB2j/uLiGY9pEhX
DbhfeA2LxNF+1lq4xexVpQ6ZU9hqpwpVMjUFLskeDuVo+xPny/ld/9GUoYUvYyXu
bRaRI9QlGNBZo6GyfbJD2sGlT5pD/M5ja2ISk8XfK60/BeGcYeFCcdDmC4Cfr/ai
4mLM2NH8fNRFqKin6jEY+mVwMgq651bSUpWi486jSB01fvz553DAHuYtchQaGJ3p
bAqbWoDx/fFwG27PefFdBCXb5NS4CXG5+UVs7vGq/TERhoLAa0etVtcOEpXLqa0q
KSDwNuj0PIUSVsftqOp/CCjNnD71TUFuXcjvZ5Z63UArnfonaQc027aJoRB6uw1o
G1WrrnK4V6GIbjeaYdxHc6Vw2Fsz+zP5fcf9Lvpr+/3ptpaBCQdk/dHHq8hUaLK3
l+IZXNg6GRFhLmSL7oGGorJtugeYk+kTLIIB1Cpv+2RE/sOqftm0aTpB0Kuj2v9Q
RRWiG6ovf/83kchj0SgJKZ1dtm/UL4zbQDNhs37wL2MmP3+uiKq6XG26KAvb4lRp
vwFS9tjQNZqbKOScp7n9ujQhKPXHKR5ohWSQzEp2DYdd0FIB7CZppJtmHMyDml5f
ITVJoC/ASUeA9JXtIfdYDln7jRlDRXvCIu98e/kiyXtQ8JAA/D0KP4UX0r+oQpDY
OhG/bZZRVPg3IgjGAQLC1YbRHKocDY4xfN5KG4tm38PXYUlT5iKoqbgNxkFiko/D
WJfTVgOaXxW72zTUu7WPTiODL4ZnBT811NiSHqOXJp1ARjMqnwh7RVNkk+Gkno09
DQT3+xJ1QBenhTvRrlfy3nYDWPGZo+oAFbceT4RQUrTgxzdsmp+B0fVzMhPea0CL
qMVpxCxF059d2CncmKzaZ7EQo7HJJZ29AvFW9GCxzrTcrcfDxcI/4+wNIbJjFsjf
YRizCrSF9zFFdYq7CLPZMetoCnLNTRbIa/9vU4cgSDrzfxV+0pqSaUjOaah0DVDB
Q41GktPtKxPEL1StqziHGvfnON08NBSNt6yz82TrxNYmnFrC8j6yCTAXdrS1kJzO
sX5bhfKIn0vhPd+VLgURlPRcpCBsSZfw9IepwPE2rX9ptK41ZRFTCdj4sPTwdkVn
zLROYkRHqteEyZgWdWWoxFCG71scnY3Z2COxbapGMZknh125inlLxS3Y6p6EU/xN
9Yd/KFNV4PefsR7bytfTrauZ2LqV5QMh/rXBlAO5W2toccBbtIVXQabA4o5ZqjSm
GEdVSxzboMtxqGpASj+4pX0c1Ev6KFC4W0inboAUZaMkDIcEOpGqXRxU0pTSS7yx
2O11ZoKjxKAAENnf90yfTWRVToqoMXQtikhQBtdxPUWuMRRp1o8tSvj3Ln87/ySo
99WGDTWuEoWXKa1I1Zuv5/nwNhfzFe7DZ/qnLf+R0vmMm6iPrdXUlnHj+W6OLxtt
ATEZpDPOLAfj+AMI8pQpL+dI8PR+4bObc5xS+L6QwnARg+fVhGpM1VIQnXj00btc
e7iuIUne+KQ+dY4jcgCPyBVJSp5hGHdjw0EjtDKleNKDOx0mnCk5Z496sCYE7Tpc
l/laApLUtkFTiXlqnbeFJxgIvmtaTDZdTdFXf1F9KPTdc9fWqjIUclQiNQPw9Mc4
/Kxb+h1UvteSIiJfEr5yKw4HKjn1DFvoG+jhdh5tTQtdplJO7nCluDty+y1lXVSb
5GMYB9dBCnubPIuMJZkYIvkgiXGs1uJ0fG1EPWSo8Lspo474e8mwbQ/DZO32I6YN
vMkxl5WGvWjzUZz+MUnz/M/rYJ9lsWD4SoEMynv4q1IxD4B4MgsfQ3WAzFXEm+8Z
xf6zZx5rPWixm8s4NH78pzafBGWfNHoV0Zk3pjhi6wbLroni2NINUzEcGkVgQOLf
VJe3mKrj/acBIQLlXL6RsS27xtTxo3ZJd12lEDhjWhb1u9BAXUEK81J4ZIc9HM4e
4H+OgNjwFYF3IobgSISjIo75WCnfc+dlu9Jj5woU8IGRX3dKkOt2ALk52kx9uvi/
uQR5DNxFjHqm6qlQJa8MwoGGwf9+iKi1HUK4L5pzxfC0zF1qw+qqWtJ8y4N9aQt1
HOifgF3ISqJfXUmfSfO5tRdO45ldeXhz68/G8I8fcGumfWH60ExJhZPRvfHUZcH0
GaVU4HD/lxSUVDhniatt3SXNxgkPP1vE/61FMqn5kdcjkPFmnxvgFTE+d/plixZC
E9V515CXCsaiZTE+BkthAOQKQEDnTix12DVfXaYpX/q3Clhf4fAXJitJErQyGmHq
0zWbahYDLu2vKebaGivnbsVeaVWmJip1bWff7GYwoChfpUCMEzwJghhkqx6mizFm
tXguz/HHKlbdBFWwioFBlvrlM7LCX2B8Q3GlccuaLwR3A+UKUUbwQcsi69BILLe3
/Z0lXg3OHfrvbA06932F+XKKckyhgC+PuCai+Ke7UWMUtGCyibE0pEiHI/nNbFl/
H75pJ1XqcQRm2/X/o/qiKwCvbKF5k0bxg/z4Krxu6IkNBznQwsypoDre6u0lHAXF
b0no+ZQlFSn2BhV7isJlDDNLn3k+T06nI7dAVurvr6EaU0rJb4rkUlQS0IiRt/rk
VNjxgZjcrdF5p5KV0qN59F4Ns7YmSKtR69YPDAI636W5UsidBU+QrKJsSFo4beS/
4idvhcUxabkRwqc1lo4SDVR8zeH7SZo0E/9DHKXu2OWN+wtWDBxJwSMYOkRuh10d
8jahfCv09BDRWcbUvOWuelM5LuhX00uu3wZZN3b+qAnLgpj8kgMk5GxB3ts2sZEg
KQDctQLmVh+r60i8ioTRuu9/m2vp/potDXwAKijNdpexVqetLjzmhY8OO4HtNrtD
speUmMy9uvGK+CS6lC/CIBtJfBdPHJiqay3rYcR7g86KYNSvOtWs8NvMez/hqH/j
iEPLcRiAejy9BbldJd6QjHInN0BvSx141p6znPdrH84wvFNmRhuYzxk7s+8aha0x
j84rHhV3X8QkGBqwu4zIkc0eX16SFtBT6g+XBfSGaO/Bs2z5iA8shQANi7nuAi4S
ff22GseGaWgaepmcPrpwhokRzUmJwaAhUKs8EmWnsbQmhQHP0J3DxOroVgHMOSwd
kuULW6OhkInVoW9jjUC9vLNTb5pn+a7AfBzMk/DRjwT5DG10Zf0XxjcjhoUuiNrz
b2wY5i80X5vSNgLk+tnyVSJp6qsgn2cg9YFAxO8iOdUzHdvN0Ie+MCFEP1pamQ8b
c00DuYM6WyI9StR/18hKvCELVdnPeR67+grIqDFAofWkuuRGGCS+KvZGP9qSGA0K
YStYLiywn9rzFrYDcM09VgLwFxgsPWLeK2InKCuoWA54aTYDvepKORYXoIRHGwEf
R6X5WhZq5iIXC+Ux0kmcSFRpzxj4QCnWzmPm3c/zz/n4l3ZkbU7jr2vlaC9XvzoP
6OdswSd/Bezkjh8d9NP9whhJSjfyi0eawzJPwx8nZsVly1YM+tJvkGq9n5TCrr+5
NeENDRvC0uSxd7ond3kjAU4Qu1dsMBwdawSPOfdDBKDyIBeaDHt8VGYC2c5unNzF
kCorpyJudxeLLtc8q4BA9Q==
`pragma protect end_protected
