// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
Yth7naeo4tqOBQiq9PO4qjomJKtxPLH/pS34VgyrMbL15F62q5DKBdoGooeJEBM2Q+kteeWT0x4Q
+Hoh3OshxTN3bbvRkQaCfbRzIWJ+qBVMYtKkpysQVyXKCjQ2v4eRrJ1lA5JWHgHFWkz6E+LlzNaK
xh86iCLUEKhTdX6mp8TWCQ226mu0G3pD18apFnxaq74/99rRbd488ZVybclnewROX5vaElh/yWn8
X8/QqGDUTwNt2vW3w1Fqwgwyt6ikDj862TQNXmY9iCxiiH+NGtaDx6vO4LweBXQRx7VD8wilYMEO
mqpah/yZVTlYYFQM6vIUh4BmLSrWJIdeII+wcQ==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
olX5d5DLZoum6rtaDP5D7Y4Jx4YchmWpJqQcug7PMRzqnyi/OTnTV50ck4CfwprIHhesVqNlinxU
MwnRp5ubYSJZ7gnP6ooXQ8CK4tEQ5uFAxm5rLow8zgXITFr90HfPbvFLPARt/vLDaVR6Yb83/t86
FospPzz8VC2EedPWsY4tWvvvI1YbkqiWnKyMaz6SJU5ICBjs00o8NZDHl4sykcL1bqMPargt8RmC
K2F213+DwaezywA+cN9nnsEcdFj3ItJTCrhkMRWSG10lGRLPayogtPcWcGOYLFLlhgLYOpUBmAFK
gnLNleiF5AF0N33zin1kh424jK1yuuKeFESd5HY8jB8A4ThDCWscG5rKO9+6MOlsgad8HNPJ/pTj
KZnNE+2AZKxWyHiCBbeC1ASnNeI99OYW4pxKAkS9YefTVzZbRf2MWa5SFv+VmB3InauG7G8q2RG8
z8Xn1fjF5f1MTYiLyyKQFBO/zK0NtXP1pybNs1HWIpWLP/FXktgo0i+EiAAfudN7JE++IzcaVShg
4MTQPE+kK71mXWer2T/0cQBV3/QSjF00O2wviXaSIBbIgtiXjWOQHAV4C34iSKpN3TPt6Jdcg6ad
xVAMRpblYcH8jtX7HGOYwjnhaYLktdHpQHOXlR3TK/VKebFQ8jQ7taFkx0QjmvkmwoEUqxkHRB41
X3FztjDTcLZ0w6Jr66D4WsepIMwDLm4ariW4dBDWYca7oTBxXy65Ik0C2x4abP7RF3nGlNEl4K18
/PZiiEL9w5BjA/Dw2uTJC5aPVYpIQGOwVK0BpsaLnqN8r5JSsz7wD4Erk7wCFHvM+/7YJfkxsmqV
QKz147lm0TxLbOK4ouQOIJZRf6l2I4oW9EG59Cg3Mg+J2kObIzwQKohVnG0vXoTbijsGzw8pyygv
chqEyD6mSlA6J/jCchakNVw8GmzGRd4HTWz/sluxBHPGdnGGsYiV6Ai0Idbcvqeciq/XFLRYsGt5
U+3NqqSj/c7s/csQ6bd0XF08BQNG+qt/0Pxfmd4xrliCbcbsQ8RLmOTPDCRZ45UIjEWb6wqEysx5
3MULXklOpZLgJ/mqDHwJu/Rh3w7Uh9CEbNOTMm1xa5jAccDeQHdY8EEMy2wxKsjoJcZvjYIdDkiN
VeL4R2wwIyKSSFRWX/1hLOSXmqBBJu/ws3mLABU6I8pXKnMzuRVgIzV0uHsLSPSDXrbM6279MOFR
ZKbCjHDzmCPsemoaM8aaCGCNdB02V/0VQvMVMS8G4XQm2MeiSFylC86GHj07ZDxv/0dgW76J2Ylz
9t1XsAQeYC2A8SoxEMxvMwfelrSY3wtWCs57a4t4EUZq2UkTNu0Pd8Ia1DY+m0w9J3tvILOL/n58
5h/zhuYSjg7KriuLmmmWUIrN9xr52/hWdPN10gJc2raao5UwUiWastx1itNo09wR+mU+YKluzmBp
SLTWN7nXWR5fr3GeT8iAWjwu3eMMWnlraqMwGQese30/BWcxxmHYahz05zsN2eBSbpPjnzKRCCEZ
D/T1PVUDPKiIsrMtIlsZ5IduCZvmVsTTq9XdKRSDNgx8BbYk/t5vvaHuUyMVEz7IZrqDd2b3vSpe
1qJR4CJvcG6BVyOIDdarw18+a0QHpLiE3E7JYnIvUuLF2xlnw6TOcg1jKoFdUf70aBZjWnNVSThA
QP7vtddWvXZb5Z1a4Tlu6Hq7l+UlJKPCcwa7fwqasQrBKMHr59m16Ypz+37khdwnXJGASvvHFIHu
sNGyDiORp8t9ndV7sY1M2QW5JIjl/zFVPKyEK0/XQHns7F/BiC8qitmrEXlNVlTFSTYiDiJNsh8O
VMwt0CMYvc96ILR9L0OZZFgL/HZXYXfsSnMSKFxfMZgWsCBgRBUaxWYo9pIxO5terDOOryXyVF3m
BJcgKRtl+2gCviUpAmMtkqwqM+LOZEaJGGShOsm+syYMCp3LJMSNa7IGqyi7jdl36hLLrQrXkcV9
szg1me5lq1obQkY1vGFRzEGNoWnSIB+99jNuLbrCTWF/lqg1U5wCNoiGVaj4VUDhTwEZxDgRPW5W
R0gTUWM0/DevZ3tDgPjsR+q6DX12p1u+1/tzjuczdaSReyiOh+kincTM1TNCYhmGLoQNPc/svpRb
UzNLfLuXJhpx2YNJD5HonRGzHp/b/41TDu+MMoapF1nkewVH6T+MJ7Qv44U9YwZpfJZPr2b3ZLtw
DSIYXeraHwZGNpvQJBPyAUtL5zo7tHXdn13fP6QH2C5cGbrGbeDPADuQ+gT9/IBEIrbN7TJ5nDfJ
NfPo4odD/HGDpHu/iKTD4gP3/kZuqyFniv4UP5y3PaEDPWGTCCf5YNYY9s6zmuC0WpXo9A4kp1Uq
WzZWCkEVcnSmKtJztz1ra3pliiB74ppKCJ3+ig/qLyeBX4xzio9FQvJpUdmZHSveKGVcuolv6iNg
gC+g2yCMiMR+I89YSS8sxBRNrmBzshfPQdZlLl2ERSCHTbrhVXkHdFvDA2Twg4epz8zKZ9cMRFvh
UaTl7f46TrgfLrWomI7taYruQrU60gpAG2jHPWQ7JekcBNDhpcMaV5qLVz6xcCRG1KWuhgKe+WDW
vkemjdxurCYV7Vt6L+m6l1tBKrV+0DyS9RRjxMlHaDI4r3+EojhQ7hZ4vzdsqWlubiJUEdnJYitC
N5cICMvRDKRaP1uRLxCTZm8h3TyWRiJN/JhCSDl4ch1YoWKg1Qa0qu8uobSjGR9tn9aQyimvHAin
JYD/CdFnZDZYz8cvQMezzKWZLBg6ghbthZgSACt0jvjL37fXflbkrl90tZPcsvql1n9HILZ3zHhi
SAkTwTtTXLUovS+3HfECpV0sXsIjSStPx5xQQme7h2obHIZ6ynegUwYnpsYxt9wNHzZF6pewwfjP
NSO3QP8kq6dlvSVCpENqxVrXfLIXqfv3fMcNTyR4R1Emp7cSSUAip/ypRX7fLU2dJOkq3w9J52MQ
BC1Jq3tYLtqkjyNmpAFuEE1UkiXuRNXyoFTNco2bLUIgBUDw/41IFa6jtTeryXMxNy6vZjjfMl4s
+dbQmy5KIlZ43v5is0dCmQgRazzQxpAlSDavW+ssMsaeSEAS8b7STfIQlLRf9vFieVJmdnC1aOBp
zzHxJP1Pyyo0FhR24ktk5sfQ028p/7J8GtSz9QDXh8CJI0aYm6O88tGlkLxn+A7NgMwfQ5OP26uS
13A7FoWtfc17N+5FFsWI0OrjxhXPpl8Cz/YSA+Yx1rwI1OeVkztEyth4L/hgzWSayxGQ0iWKEl2K
aHbHdI+STvafhk6jb0X5pK36qL9GX5Y8CMVjZAhGoBXVgPpPR6a0FLfuzxzw/rIhykq0usb0G0hc
8avBgQbkXdDiWXSsCefWEmefIu/kdgkQ4HFpKCsNXdLw2O04Si0W5N8TArawNLIhi/ydhZKwf4DL
fkTymYI4VZguN8SD/rm9SQUy0sKMWgaCGKyz9RgC6NYjUHWZhxTKWarfiDi5Ub8gUguTTOLlfHeD
AqVaXsqCrzmTtbsowNBB/Tn/VsXYyfIQnaprmQCqHpctY2Tgp1vfWlpNtXnIDODw/PeiaVfB6zXy
ISHBj6hOmEnj7VmwXNfG2ZWo2QDso2lFqZG4sQHz9omgNpkOzmyvL+NGjb+njnNQf2ji4hrnrTBg
+kH4ERnWfqQEQoEWZdEPKEG+oBrogPiwDmQ+Nt0MhEhVWOojUgCaKgplioBLwyB4K41wD8BV7c5+
JPpNaati9KXPU7lurhOPfLv/IMZT/bED7EsBfGPdPA4tp0gW3IaaDBVk60xyTxFPaSEBUwWpPGna
h2DzG0Dh58bTVUW5WnFVOnVOfWO41PQ1/oig/GuFqck1BYBUOjkuAH9TL0FrCA9AY3x1vCrYe1VN
idVFG1bGaa9rCPURtDw2H07QGyrn/CP73jCBGifZxKBikssIMm6FNgo7HdZBK7K46IHrOzwZalfV
IcipGHXDGp6ft3ms8rgtoOJPRSn7FV3m7n9g9RIm6n5n8cxGancDGL9Fs5GdRrux8YonhRlSlQ/4
TE1JEdpLO4CTbY2ioOmJ6BhqIErakMzcLEDyk7SFiNreBi/nhUsWaCw2qGH3vxbI/FXIKHW3KVIE
4sR5rJfqgyUr2qLCxt7FcrsPlrip3em2Bzh+bQFOJjvHkTSTJYhfQNam0Z4ei8ZrfS/1N4E0kbkq
p1aSsAWLMR0fqi6qUQnC+28c/NL5/5LHiYrdqCnviYMOkHbArYc5bpvWZnniCh85DNfNRsbnIP56
JOTZfLFQTp4spyXzswvibSW/ve28fwF52AwL+xpQpBLszwisR1Izd3x6X2a1vM4RNzUTWVbJ1OYJ
LvXZ2vc5M276ta7wcxj1Sw9w6DSvQXFHrqV98BvMbsdEc6Cv/TrcXtrgrRdKN/NHK+weXkUNFZGO
n1yrAJEMdJBfm/QUrL9Oj34gdVRxtUc0rA48p0ce0MCYq96c2kbN6aibCBuvKqCqA+FYTgtYiwGz
qcJs7tGpjCNgzhmiHrtKHdWZvDHoXqbfytWvXk2oCnhG1KPZoZ0oZbtDHwluUJzYq2R8+ORoE9z+
oCmVT8liSnO6ES/hYbBC3vSJJpepW//Kr7NWKyMghi8UEXhXduVGSBQ1CfBpgckWTCoRnUQ4Zzqm
oh/hVJuCGPN9xtnZiGq2PNpDkOQWSnNT8ghl9NSlCb1N7o2P9JOAUV0qofCvqjawHjLCpyeZxdoA
nzAOzHObxhyz4UvhruYgIK7jOe1YiGVmfkK4DvJpMO0+ZtZMYokW+ejO/ncbzzc+orOhuXTb0PiZ
Et4FCJSvTx95wj/qIW6914fjJXc6BFCb/AWb6WyF+49sW+A0SGfisFLqNfdAh3lmA18Mh8xuzlJQ
qfFhZyZWEXbSN5yE5l3NOmBawCfVXAyCAlxa01VRUiYL365AHPwoNgN75Wwx/IkMX4oHBRBJUL88
CCKTDj1YWGjCB7W5fMudhehh8+QNHMXWBKzA0PV4uOGqneUU0iSp3/K9STgxF4H6yuAwh7JFnBcP
b6uOPweUH9X+nm1Hl0VnOGJpjjZXZg2KYfsxdJMBEoEjOuyKFs6lT5Gq7QliWYp2smgNZXo56ilG
o78UGVgbKTgSAWAbfCsy/QtXxt8i7A2AwGFFKatMNxBeI3LQmcwaku5h2QZRuuTXtjttk4DHjYil
whgZkFgKWeAdBxC5qAWY6yS41Wb5xjcsElBAts6a6FG5wm9yf7LNR+VEQQqYMJ3e4YTa4oWsfjXk
fXI7BlCS3ytf2pB7Bs8YW9xFLqaDsXDx7kOl95LV8IDikGM0gwfEyITV/03WI6hCcttPCRZormu0
1c7W+7m5KfHszlXImIcHLxDW9nEzUlYW2FoSddC/ac5AoWme8g3sNrIkTryqeZamSYOOQnnhR58w
6YzDeDYdvO8Pjg0J/cSQ0A0d7lCYalf8wBhqdW0hbyoIEmDJkcf1pHAlWYwdpz9Zkt15Jf9IKEj1
cO0rmEQnd7Jzsxs6Cb9OxYEx5Y+8bV1mhkaKdo0SeYKy49dHzyaZfbq5mVVe1KSzgW36oupwOmVr
c76v7WXd8bVnW8s1wFvr8dPHDAv5VjUycaahZCXlRW3peT4qH6FHfg30GHBCeDuROMEpHS9lwpXn
n0aFxliiT52A66izvt4nPJHSan0qRgLQhR+0ZEP+F0q+dTJ97nE6tzaK+4bPmdByeik7qKLSVi0F
EOl8qF98ADtIdmnhkXadEAXouvRWDytP5sQ+MaBPAurScoqFeLVMgXXOXAtnqi99Y7Z9w0Ib88Lz
BkVlbwX/GHxnj+Ga6t01jGFjYqjQGYdXWBi3i7UZyEdVDlQ3xpkfamUtd3yf8/y17a+5zxvCtEzd
KEpmrQWvqSSjTQXYeyjDESrNnvHz06t/l8zJQCuwkDHuJKbLau7kRwyNJXaEMDGnP9nR80MBuqYZ
VJgMqVCNWxZnvla1wvU662MsW7XdNvHWsaiBZQWmZqthFABFzXQfSoIhIveW1Sbwi+4OdQLEGZwH
AaQ57AOjRv4Lls/81C28+68QFFcr4ImaTwwdpk8IWJfLoGeBrWtuCVHGU7tPnUA0BsQNjbfe9Tmw
4wy2xeBaVI8ODlqlkCSxEe4SX+LMsoQBPMLsfy6utpYsyk2CG2HZkPUP/SqL3+qf9G92nCwCQOT5
42pWL1mWY6Tkick1sdplxYcdI3z2x+6IL5m1mNpOeYAZbXvjzcpMuQNa3d6FM2aRsS1l3Jg2vAhZ
BrCkX5vMYelxcXi7u8oaPel7JL4yvba2OMk15yJmE1tLopysdRwSY2WlGJXxkL5hkLNj1hw5cDmF
18f5NNQXiHWAybgfK21BLtNTLDngB4PRhhepERa/ku9/04rSelfDXFL4JKB89DRTACu9V787VScQ
qvRYRf9Yqea9vRqaJnpEh8YcqyCfn28WEPA5fKGk8vpyRvJHJw1VMEw8beGjrJi2ZQpu346lEgpu
6Q0kHrz6zH60VM4OkOPMFwD9CMcYUchyD8G2jHeqvHYlN4+oH6OFpQ+DwkoJAtWzNBY5n8FLlWto
NxtRbig8UhbBnpBpRTTlOikGOKMKGojLFSuTaeXuloEFoZBoYRbgvZjGhkWHVlwtkwMjB0f6h1HM
Yp/z/wZdsbph4D18K84CcKI=
`pragma protect end_protected
