// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:35:35 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
V2d/ORguw32SeqFsN+6Y5IBsbmTdW4lrgN4ybYPZTjGRax/CHw2lWG86s2x+Dxk+
K1yOPNAllcAFUjqSXQ7RsM5kFZIV3kDtisMv55dK49QZJQXz8SYBiXT0uGMsfeUa
sMFRm91h81nI15ZdetzHpXweL2nEfs0EkPc7FpN3md4=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 11728)
/vdM2vrQy4WC7XVxGBLlggaGI2YitTsQHDQPCU/r939/CvmaxEz8syw8jzRWSbjj
G/p1kbPnQ2MEddXmMAlwox7F/YdNMOSTtswa44EYoC6u6F45qUUhVcigx7/mRQou
pvwoZ++R1cWBe7xEKsj+YxhgSWb0YwMpQ7G/NkCyQLrdLz1g7vVXurwHr2Kn3Any
DM5rTgYOYLMz0TKiJwDvNMseEWLdiiArSTS+Z1D1WYzBT33EndW9EMDfNaJwh2jz
0LqgT5WWkeqiVUx6GHXTcYsKEFpg0jne2pjaeXK0gPWltdaBu/d3iy8LnN6pVmzS
f7LX+r6/XaY+BwCy1IuvKGVZhlpvi+BLG6d1ygnrLI0/wB2cYprLo3MLp24Sq0Mf
09yUJlc8KGENFuJWQr5EmvzzJurGkQkPXMhqv4a2cyAHnIDvJm8d86cwNdaYoJ/M
nx02KfGvqMBK6kIRUCkPNggwGN+fBb+L6IOfik78290Y8x/tjwuAtyS4WRQmt16r
jRAa1rDOiAzeglqRVisjsy3hArGJRBximwQn0BGVoLxQHPIEJkkD0y7CROtzZtRN
Ry3xUQnXesJwcLOU4rjubg+HWEiNTDrsS1wQRtkOfJPiBJvi612blRQn5XKHIZXe
p99kGxRfLTzkDcrMOdSJcNyohfiVHB1Xf2sb9EFR2ipNtvKpFopPpiOb+rxFKf65
3cYrnXXdLCsUAiMbxgCF7B4rWOUQ4q4DF/Ls5gmlZ67ubp3dUC2eoKPFdYmmqJyg
2ZwKkIWVLC/F97iULMaQKcdfH5ZbTgqK/iqQfZcLASsVJdgukmFmSEFAquhGo8/n
AXjNL2oTRTrZGhTfy3wP/d4pHTVWAFi/Sgw6pVbYJdKnBLExEHGJdAmoe+wjfc9/
E8ykllZ9kDgZlqyNjtGRldqjwV585wMNYQN7orrwyK1eh0xBnge/2myJgLykGeRB
FFWbK3Vm2bUvqqNaQzzLczXtGTbRD8pzlRKXNnAtdat1MZXXrj/rDQr5MHWg1x5t
uCk4qg88GrpLvmveY7ajAjrgv4QLzV9tQVu0QmEcnXaxzIxfNyePE6Nsuo1xiibb
koQMkR15coU9ft7MT6GyWZHxt/LwI/Syi1W5SjMN+zb5CINiK5dT31bVhavkrHGF
EsgJ6J+X2sDKSNvY41MWgYqlhqRXNviJRW5oFEYFKSigOs8pGrAe3WXA9frjNeWw
DrjA38t/x97wPHpzPjTWxfG02Qd+oicPssojmE0T8XPieY+LQuSut4j7wokIzUsO
5sWhPhm6iuEca67AZEHNAcqbc4QFpqXM/SvvaFqKNJtChagRTQ2Ydq2r0bwAUkLZ
7XjMjBRuR2L4mAmpNMj6fvHCHispnk8eQal+JO/hMt5I0CGO61mteJ8Tood/KgFn
DBx9UHM5PIXsg8dzcY/mUpNDvybpl2aSSNVU5Hyg9e+JUigkrfcogWGnVGf+GuSq
9tvLcFozEPseYH1XAseUC6FcF4bmBGIqLmRUMKkGO1g+h3pH9b7p1UCT935nca7U
EX6yEDPnE6xSmsLhfhiWE/p6YzaxEQBAH14U8iSC0Y008NXYE8GfAMzvraiacjoY
e6WA/uc2gTX00ANDXtTUadjC+BJkr3G0fP6hCnajxh3EviADUP7LLgIcfVHDIEDJ
IR/iZ5NH68HTrR6I3rc0mDDwqVKBZSpHvj5lqziWn5oRNuosn4Y0CGGH94Na02W6
435T33S6ph1b7i51rfbAG1oFkjEDq11VJXmnIVo1CP5J4CKhH49hv/I0JvFSs+hK
kQRLnH6FHh3BEe17SfofEJh0B6VyqKQFhSAWWASXOLZrm2b8Pg6LlaGdVaLaLLca
wLW5RvWiN4vzSlkHPbyTAU66lLY3COc7tUlwkV0zm9rJHI3ZumGztAHzHx+k/Ynw
SkaLhSLV0m2s6Q3J77fIr5NuipM6xrpNd1cru+mA9L3O5XLsPPlPO4iW/YF5DaK/
kcEoKRb+UWlUjcVqE6+mi1JaYYZqwzhLCnxIDC/wJzkHV9ijccicbj9AiHvei4+s
MltlMt8CWn8LI5xcKeie2t0o44qtB7pZ8nZRW2GxVRSMXUFD8NSGlmSi4TbsecZH
fj8ckqOKYsHvW4aLFWiJt82GeS7H8ZpEwzA+RX8bVK1h7l/8EOT+rhOdOGHPFdtu
43UuNOrsTGi6aXcL2ukNVPwdbbAd447EfDYCainz97+EwLIoEHqRCqlTFjTWV1Qt
OtfWuvNstmM91BJAEPbhMVHd3O5BJ0ez9mbPlGXA8iLxtcm0TspNZxehSnXXupGs
ZH3JH7J1hE0vmWWua27IITouaM691nxGz7rSteAqxDmnxVRqSWShJONFce5DiX2y
eRJPHUPbGdrUfaWQ7G30kJ+Z8kTiauzGTeXuf5WV0ioBQMJbDtaLiSm6A2J+Wf/7
nTQo/GsIDEfTz28LqACGniKQixUxHwkSA0J8jMz2EdRydO7rRrsRUxVNwmoriMCk
dc3sm1g09C70f+TcfPy7Wj6FPEBRlc+8yS8dAZanFTLu+gK7EBYOivGypMxgKBU1
Enw/oiJbhMDbV7vtMOkfPv8PJPhIaMxRMlgzZEA+/A4dArOyntNl5j8DkN+owX+V
2TbA0dVsnb/9xnJ/GI+tVfTKaOQk9zgdLIAw483BsiE+sALSfxQyLbq3en50Gz0T
H8tR/jUPNrkvF7okc7oJHv9BmfHbE5kOE5GhQW2llR6cELxyqGcuY7f+3Gtl0ic/
MZCNNVL5j5nMnFl5khc3kF08Op4q8hleCwczWMm9lqNBgnLzXBWNSl7vfoNgkDHd
rQ5AOihe9uOTt8h1Zv32LzDQc1C35ToITbHHukjYGdlhCqrY3atYMwHbWPB0BA26
NO1ke8mHuNrROek23awPZ47H4JQXyfxz5XA2chHPzMQHjpvnGAOixWWDsh38l3OE
8QWDbnmEbvGCW5t2anfoSqWHBJc4nKVA9VsuI+ssu/LV/tUPcx3BWWroiaJJajdF
2055c/4kFRhy6DrAzLnePvT1hjHPGg2L1RO3Pb9eXXptLwDcUBhC6EJKz3/0qD2I
M0yneWwvCdnLNJCBUmxYt8sdwvCxYzKBxy6pdCxzhM3W5gYOnaxz9GFtpD42QvSZ
OgLgNrgqULKKIGbX38ovX/4biJexeE87ObSnz9CA/3lDkgih3pbwD4YfYAuONzXS
TvuDyTcCIys//lklJdUkjwx2Ct1D5XzMOxnX8KDa983ADIeIW8umsDUNERsgUssC
TAJS8O9qsfu9AvFDWkSF2PhSRvCM3DQL0XhNG/ixJMLfXuhyvd5LX/7tuuwDYsX3
j0/0eZOVJ7mXrLt6w7CfUqyL9Z8B1EhG2wY3LOfgCoUQNQSOjrhPEc1EXvJbMR06
+nGg4MSCacMSaV9pz4ZfxD9cf2kDQAYDnAgWrS2PlKPXywqKNroKlx5GZT6xEbYk
xn2XAAlqLGulrqrU8EKuAniMDP2D5hBuNZFhEQDCJJtwgU39R7otBsoEmN7YGwTX
JHWJzaW0/nUrt714E3D4xHWyfRgZyCt/xHhU+MYEf/2fHCdihMTmEk6/CJ0Q1gHn
yprSo5dyef4PTKsXYH85Eo5HZrLx0UjugjoYMul0ki1E0ZmAanukyiFz6mtREIMx
hjGbCiCMQc+i6tjIFxww1TsPF8EkHHCge9D1Jbzxnp0GjNijWhkyc9amaF7O7xum
YMyQeo/vvbuMd1KTOCUAoubj2CqipLq2bmFVXn1M94kMPf+9eYtULqWrqrAdHQLm
yuBmSdSUENHR03XPbSEmmIKbQE8/7qlY1hFbwBZSp5S+N8d1V/YnKpcaIKLeFO6J
7MeAzyGpR75jh/2fxHrxsdBxk4IPlYwQkMw3ME2XMT2e6EJUf3JVZ2VHSrwz1nfd
UNg6kyx3qdMYdk/lxxz6UspegiXTO5SmaIkoBlqxijLKrnDCqbIZMhnxmiS2CUwj
dr5W7MqNFyW0IgQgCkVzFf6PMqTNGX36yi395qkwob0gUvxKvKaHUaNNIOAvnm0h
sBtja75Ae/ukAAFuhD9RrdgAUhqhJrMsqt6rP/6WMrus6rUPaJjFhvcpZYYgRXdL
JrJlG4GiScf3uqlY5S7NX0MB++TsEIIRBaefQ0ihLExV2iRIxCEefEgKPQxe5t1+
9U5iKbLfU8WUgcdbxdcAFggFrj17URC4cow6AQTXimzrxmMKxikMkK1E9ZrSwFVm
BwMk6czwd4FeGfMm2/MVbrcvIjsEZ9zdb2THE34RjoRocdTQJdx7AkNYwryc33nr
MeIaG0XxoC0WytWSRZs4+E8dlFuCgAss+O/BYIY5O6zbNOpyqmbXh+yPRfhI/38H
sRe2Te8ah/4KjfwS5Xgrj62ljuhcrNBvdUw7hS2qBL3Eh/W820WmXntFKDdIRqt/
6L3gGR7Yv0Ykfot23shoF1LqmejmAnObfq9zWMbeIgiY2BTOfsNSppL9sL3ipCmp
Ke+I9BPMc7HJRAV81OefQSTJB+dk3FWNPTUiDxmX01ZbiTxAYdiKVHWM8TNapsdw
l20rgIR8doblIgU2ASCmzSvgHX/6YkY/0Bv09nTBubK/N3lbBHglT9TEQd1lxFCa
FRgCjDvGgcwX9HkGZ+8MklwvvNRaqRuKQUy9qQ6QTS6e/332LvApEgpopFzW/RRo
RWQAHWZC6X1VgPZ/Xa2BGwyJDzL9WkRcPEYEPgXQpj3DnIwr7qGCSprTUauuliI0
3CswOXM5eHvAua1EXo5lcz4voUGRW7M6tEemRYkqGG/Sin7Elk7wLR+BIC0lIo0d
gsYDw/KF8RrTjB4Mm6QomFsnqHoHLiyOE7+UAyAUIVnGnWl4wNQgg7gBmCwyu7Hp
gfq90adfuIWsHjXHRQ9m5h3UCznOXa2N2lNSMV9uZGlzPFuITbcfiDPKZawxE6gt
vcTe5/7Og/B9sUMbbog+ZSpI0kdlnm9OQ3ocE99vloAeeSWhecT8GFwA3OUybWRI
sp0LldT2FMcuVi9zqZlS3hSd7sv5ZRK2he/DiSZ4m+nPcv5UkHdCBlTYWgUmn4fg
KPFoYSj2ThzgKa7KDFCo/PWX2rhdVf1K/934Yg+U8nS6HqyYynC6e7s3A/sT5muH
f+cv9Zqy34GHdp9hL2d0qQy25KxhRANWW41nZHrAPJwdtX8Hpv5mmY8ZfrN3DDrR
F3AT2P4a9z1OuM0QviFif9WAiDSR1j/1OVaZ8fYvU1mt1l1aXEHGhfe9Co2SUCxG
Zhw+nyiUpw0U8AJqZYCkck6PlJG/WWG9jLNMpNeV1DJlAesSDJ+M1qzN1RfsJJNZ
vkx9oc+Hk/uetVeBPSj1RpdAlx3jRZxFb4mtt9Bdw3I71RoVd+bTYPAsGVldoL5M
axlo7aisLYyPtQcqmb0GZ2Nj88Ff6PMxzkPGsX3ej5mMisZkIYys0xmi0bwKco54
KkRVNPuPu7MT7TnVSXgQHYtAe8fvdpSq+FHbrn5H7dNp4PCDb+dVP11CTgVRgw0N
GQzrQQio8AmLLt+NOoiBycKsMVaMew8hePXvyelLDd59xSoa58TGPlWZSHJOdAo+
I0qLc3Yb5N7U7c6+epTImsAMWBP3PaOLNQHhLoibbLgmdEYB2pWnKQ69XnsuyHbP
CL/SnWbZqXUJBy/Xh9C0Li6yBTt1CDhPNZrn7uQdlQ+6d9xZPerap/iit0C2NkT/
+PbqpKQiyuRM8UP1YzCxirod/jkfqcOaYuJNmfW1H5r51UO3G5Bn0Kz7EhapXsOb
aJggoHx/lZXvdNTkVUH0YaGpSE8jftIXrLQPngpkhCT+jBTgCuj/AiSHbe2jcTZx
0ZxAqRcpkgrq1I51aG3vpr7vs5xrWCSOQU3rsuLlAyunvXo/VIK0pDjXJ+c1a8m7
szAT6LnyTF+rEd9BfdLmnZhyt3p8t+pHQMUjhCyAZeZzeoyChpW9plkF9Grk0z2I
2h5KobBpoA/Xcr19EjXhZDe1Pz195L74FKwvP0VdrinjmeL+2bQZbS+fg/xZCNGD
ZoV0UqKFS5APjSARzyayMi+SXLhVVk2zl6zykI3yCeljEeiPaRoc3cMyVXk64+Sz
AmK1unOg+ayDKJJt90TIV7xoOgrlIrgNcrLsebQRVr/YQwfXDQjrh9Uzx/1lcJ7H
AvcOL0RXZAUAiLKtQ08+EMtHYkcdFj2RzHEm+3xV7zjgSaknETaHx5lkTDJIlYiS
Gqdo2TVWnnh7xSl7YEYrTOSB0QohV0NteAhWk8xJfipFlIpuWasXEZgg3/oiHUzV
JOlghTwY7q136RpWE6Khy9r3aXZxQC/ZLhBe1er+yewsVrCr9fTfbwRJKf3Aauik
958TTw7i3j6a+Ke50aulPkoaVNSrSPrLyMlDD6TVunrJdnU4wtctWdYG8+sotdgI
hznqWQzFqobiYmru8dU8VriJt0joqvpJ7qBFj5v8CUlziERDW0L/B5jtjZpy9Aph
9e6UlyItlTR+mhtbe59L2NaRTW07auZsqyo6oWqHG6l/ZTl2jmUd0agXO20PjePk
auw8LLP8I6tZXwUxmzYbLQJskk51iHh1Pvsgp34KhJ6qhMx1lpWh0tRooAgaGhzK
NmiSLR1jdB67F7vjDF3iCWwWPTS6l4dvObDjKN7yfT1KPNxkYyUFJQePsmZA6Ury
3MuvI65SvjNfcw1QADthnHMfpXnrpJGh9i0qPJ+iJwJ1I4KG+L5HcFAeoqUfdwO9
nq4D/Zvg8Hd81YX5rQ+0s9o5bK+QtMFGl98vk/H4JqtvOUnATx5jln9JjdxXF41B
OsCv27vMBgquHS9IdymkgOfNE04ACFMmeTskraKkTKSW3DxqvToNmLfBIiXkE7ds
/iBRA09yoC5j/UaSXTh/d4W38A0Xljxr1hWLGpsGt7ENFch4cbzECFkQpDIotoAO
kslMN4caFjKFtfiQCf7aGOHdkK90HHTM/Afix9OqZh/QKyvHyebA3A8F4XjUPD0F
HtSZHtGTyWA5DYkWwtbzJuQBnUc2QuAVF8PD9sqvPvvn7SxOAfZAZzQbjXQxdWL8
tGiyI7srGNMzQ7NbU8zBQNgrsX5Y6tPIb7pFBm5scfnahhrxlPhvuMTuOOxJUKCl
381Nb1WxekQ1lmGGB+BqYn1lnElIG1s01tlQJpjl4PM4u6JgG2UjFSDAL2nu1fQ9
6Xbjs3MEb3BaD38qod87xmBVa7OCY8MtxzszWHd+PZqjGU+9v2BBb959WjiirrzI
tqgtr3GACRQvcb1sq0TMZflzZaFhcvfe+NXp9KnRq8mlq2AbhkKgH9SwG5y1RGAi
5dPtfbLv4Z8e8kcm5bs9+QVzaZmpxP02UnRzGOZKbwiLJJhTPbxpet/6/z/vE5in
mEGY6cG+Yly6Q6kjYpXgjDqOTPsa61wGcyHDFVt/gc7VjxdBVXcBHV+l7iCnBBVn
lazq/XP6T6kK5zSrOLbjwsCjhw8DUNIrxLfN5ucXt6Yecyj32+GPVHtLl3M7Q2mu
/aMkKEPWDMk3NNYpZi/ZXekkp31hMnpmfGsQ6e8sM/W/XFkato9xp1GT4fLJQKok
8Ulb8r7KPOKmLZ/30Vhnj4zwRqE/YAiHVIxR5LJGi0t8hY1O5VRR8h7Nf31OpzvV
MrpG/DIrVRe50bvSljAp4si2ilAABwmCtLuksvrHmoCNhMsTU7JGasAGgY4LEWkn
H94JjqSgQZ2kYbESBMg764ShvlKZxYXV+FBkaH7R5cSN6jy52S+j8mT31HNg9HNF
nCICmryBcv7buneisY6E+Qg58ExhuLb/ea1In1VMX5MZHHm0PjuDYyWdY0fve/YJ
E9JdXp5b+p50XuvqWQ9pxP80N1Rr0QOfygbEjJs8z+W/PHAWybMsvBVSPoHlbKkq
hb0b7EwtnSIgxKHq75YwgJTSLb5dYekb2KDgWWnRGsjZRPUlbgKY3iAPMX82INxX
TjPDp/0/5M3L06JwgN2LBJQJo17Il+weAAcZVg+BH/cqyY/QrRdo3EHcOUPcj8bC
QHsQ+aoSswpT1tyFJ+rTDA3dpGreLspISKtNdsZ+fusktKawyGDCiPETd3XoO++A
VRQ4xI9/oZNNVXOAd38he3+ugvwZ1XYKVWyk23FwDK0iqMnYjzYd4VxGBgCWHwxa
AbomrvJsaPFhdNikjtl1puu+SdFh734PV4aGLIfAHBPHfpZqTkLIlLiFH/frx16K
cS+GxDZ1hLadil1EIYXoTsDoAeCTF7eDHfka1Zkaeo9QuErug0Qj2mh+JgWjYHxU
TcliNN/kK38yf7oVO33HGY3dCwEv3gRFZoV3XLHLiVESTP/3KDD7yB/DWVfGDHLS
jIvTNuvSYRxVicmEV0dVOHVh7FHK8yXUsA8DUCzKaFXtRyQ9A9ua7RdyCrLWXhHs
kpA3M9Dt7i3TdJK6GHfWOE2Dxyerfd3tcmJpxwlZBEsvm+ZFAZDlbBR/HbD4+YUP
QTlDbWqOiMVa5ca1e97a1AlowgQZLM8S8ckmDXwRjt7S89hiAFq1JvID7ub8Fpaf
JJeqKMgKu1yOScYekxhrdn7SGpga4GMX9eOKofCcB9cOCaGXoMFGqMoAhGTw0L8i
bd7U+3Hm7WC29yEuamghUDEBoCXkJj1HyPidgkNxjq5T/IEhH6GNXRwyxIAye8Qg
DF8i1BYulDgrFhQAgznAyz6kEQXcnaJpYUijHi9YSi8kN925H6Oki7QlhcYQWNVd
BMVtN8aqeeiU2jp/nb3svFtsiK3tJiu6p8zBsrL6pOhHrqB2p+7cKMDYNFNPyUdr
oXGNEeI7TKq7ldQ2wh+1GRDQbG2Jda3Dj3TVUc4YaiO72//x2V07skuxXTEIc0PU
Nkn6zi/Cw/3NuAefJ75sZMbLaV0H829vxnq+l8cM5/ey73idhPnrGKXff5gYncxQ
xvA3/UEa5NXSImIn3O8wCqzZKwhxpY436qr5wS/tbYYK9RN5fR9BtwCrfA1eBgZu
s4g8vPX8smcRHuW5HyQzmFvQGh9bSV+6peUOmcPSZCEROVaD57ziMVx+jl/EXGHo
nIZBmOJhV7sHHTRFSt7j+w+fQZnZNG78AWTzwP4e48L0+zq/svgrE3MorbNfMoOg
qHxi9wnocXpdpbW/ZnOjGWUpu6fMT4c7i2ctUui7xfq2adU7bOB8hOvTptz1J1CQ
xqPzlh0qsHtRrsUnvAof+ZgWB19+0k15RwRDWaNr+wwdsxzQ2Wsmgh/ArfdkNX3P
bzr/2BBi0WyyXn7JrmqxUx1eaB/bTcwHYXMzOk7SvPjrGLrN7c9rxLhx1pWV7YF4
OJbqaOX6WlAo4Efz+x1mI6OlF51h3tqpfUZFi5qsG94CF2i6RO9C3KEmmOy7nayH
iL8AOF9nz0VELZgxl270w0W9Tlrty0wr+OtV5ivhCt5JH1EQMNXCMaYQTSYftlN8
3CmgMUcDmlpJGTqtCsjLvU5AsFnF0g9/4zpum2Dp0VW9WXyWYtZfWA5SgkuT0edy
yGVKv4ct1KlgeKaceCseEVuF+7hCw0a14FPc4dAG633mZHvXrOv8zJybGYsdfWq6
i13C8UvROV/qAiC96+V/8rH+bJeAPpzEEs5gS2gn94GqNr1s0JeqcUBFA1Z5Fp3I
vKHu5SbrhBeUx/+SOnLP8U4oFNTpCrruWcBS5j/fFqZhZk2rRZm9r1lmIe/EbkAk
vF9gJud6D7TTLgMeowde+WTe7iyy1fdiwoW/MrgA5mqx5YKwvqeA+QZAkYWRpj3Q
u/hP58A7+RmQJgra9I9wZCx918raPvH8TroX9lwQSytQIvmk236UyDQgAdRCDO05
MyHmIDCuVH0ndx/slbQReYyIDKYMVbtBYcRkeDgIQhjGF3gkdsnrLJAGPHiWNwuo
ez00ptbE7PK9g7w/qg0nuwgsLC2aqihvpB1u8vvAcGnJvFSZk5+dUp0kSR7z8Rb2
pmhGxNbyG3wsfIy/FfCE/C7e5AvoIJppniiJrJ31o/gSb0iI5hZSAIpOHxWo1/HF
noaTJrxlqwL5peKGKuotMxlwkskTNuP2q7VrcmgzKBESp6xEOajZ+gozkTAX09aQ
TlwjYgxTi+WajVKT8NVZtZvjNj58TEghBtQ3Rc3m/OyXxdhvZOhCnsFMOP11TG3t
XMMVPFvoYF+OfxF/WRGWsY6wXAphOqw7+vlfZhOn4RbxESvNJiAivhJa0iuvVVMZ
NqsCt2RReDqA9V1YqSOUQV8L2ESYVgs0ZOUcK57D9HpdQ8l7G9Oa7aLFMDHcHJeB
e/qwnsjiyaQA0YV0+vql7gCo4y2hiKzf8bpoYtqE56tq0TtjTlFcwUv98fkvDOeQ
PdK9jaJzzytR9DxM0BPDXB26fc2iA18Bf7WNw/eOR2iF8z/CCM0Dy3h4UxToBmzR
LuFmGlCqDIa2nXCfwy4IuvzQm34AKRcyjTU5RQtqLLlh6hWYxRnBAZ9b23sdH5VC
IaHK59iYf5NALhZoNYi0pz5HH2ftzte6k3yWCou/sJTgAEVJqyYfXLp9wTVIeTGN
aNbTkVzIZvkeObJD3Cc66KlRnNz1xvbaqeAx6M7XfxeVB0qgtGClf8TDfk4QcX+P
CVBlSuFKLP5oUAA4y+OAS5EVDbWTTvXni5y0LWMnfYliIctwr/5ljGfUWZLQxRAn
Im0ns6FqNhJxAcrG+q0p1GJxzEFJpLxc1KihIoINwXNVXuvfG4hRvZou9AXsTx4z
/pfZroxfa1Wv1wjvLJ60wWez4PfUNu4fcmxhexDkaNRg8srf5AMOW6O6c2cSakq4
mbRBQ2vkTVV/oMYGcPY/6URpeaLz6FWLnOchF2PcHkTby+xjFuHgO+5aVrsa27gn
iSWWGPaAvceSbrtCd+4IQ0ZYYDV+ymRCiabUAGT2rdpFdQdKLwQCPo2d+iE7wZMP
OIfHfTH5mHHuyqMVYdY3ExWy29lTYyIulGViOf8y0/WxIT+5bEOIRa3MoJ6lZ3Ld
lUjJjlJKKxKIn9J5imi6dWQ/pjl0EcjhHiJus4+aOHuCrK5fEr/zu/MRxrThZ8gY
Hm6eSA2vzdKtBuEpupDoqu1pHZFHeU3hQ1VnBFKUnvAxKhNVZrwtpEdh8llW9sOQ
bb7H8VuEsYrsvRsnkX7lSR1t4Tgho3Aw+fl22g5cvnh+MAXGedZ/EDaDAUkDe3jC
BYUd3doitms4vsMmNt2x/U07rPB1xgzme9alDfvfVj0GYVbw5+N9JmuulcbmXNTp
ilnGYicnqhEGZB/rZU2ggrrtlL1C5k+qfIgZiQO8FbmHPbHebz/IaqT//wp9W3rh
DFebUbq9nsCSrgG1HB+/dpf3OGY9ZYpw+gplpz9KfhUmKCEYC/4ApNcfJpKdVzZQ
mgobyETXDRU5XjB3v1O+vRGamNE/OJUBvCc5O9Fyn0jpqavONOdGld3ibpZlG0+/
+k+Ozmxn/aoYR3JlpQaesYX2hMg5qasKKlsDl4ZeBu1/U+1DfNXCcVcpUh9wdP7s
ZQHWhepko6D1p65Etq1jyXna7RF12QNoCMvY6yqRdi/bOYr/JnEFGVAVJmFo3oGx
9AGVj6BW0qRZtmeiYMreTmQhoQARP7/WJffsM/YdACB53lQZeFeHdtEgHSWnRAEU
0nV2VCzFXgc6XZY/BtkaLESy74fWi9KR9BTGK1gVbGtSbAGZPXvxnvwTf0Fo1mS7
Gs5+laCJ3ZAvYFULnpY/DGaZHys9aAuWPgb33/VEmC98Yn8Fb/c6gwEdkK81IKj7
/SRgm1cUidYZ3AczNgyXwHbzVYI90/uVcQuvF4+d8N6z+gfv+1aO94McHPm6XXtT
dCUgIWvJTgMf3i3YvElfB7LK0BU5V2tC+TuYhYcTj6GeIGUtqUbp6Qu4WBGrA4FM
/oesP4gH41wZC2DUCyRQJTA1AyrShUpgFRLPs2kujE4LXUx0V4oQ1sNs1OplLvBn
gZlY6m//6mgDxTiCXixYD3RVmJoYOGHlWuWJhUI+UNIndYz4Ctxf+/8Gu9uWbVBC
aVVB0Dzzvho71Lw9o5+PxHopn0fKKYBAH9gINMEOANGc6JMSIwPK9fpv2Ah4SIoI
2E1be/9oEmLafAdE236FV7XLD0e8v+mHSSKvrXQZFaOns+XbOqEx+9OtD2juCaXK
hd08v3Q45p2s88J1ePrx7And/8bRp91e/yVuYR/4gf83qdFhZX1xiHxrgJPZHAtj
xHDV0yVkeXaiypqOQlZVC9nnpIqNX+AjTVAvVXNGKnnkdBahklf0abX1foGddptB
4qNU5j1j9o03wVPbYAaid4ZjXCZbHb8TDsnMfjo2lGPSSqhHxroi9AFhdorSDhPS
7iYzeIQRZx4LvKc2HnUUYyyfw8JtsN2D02vXRk6pHEwpFCyJt0iQKyn5uaI6U2if
AHJgRRTtoG+/82kk72zu1heXN8Qe/UhEfoWatpJGJ2dqxIr2CsB2bdLpt6fxa0Go
gvVtyDwGY7C583wwNKYB9ItUpVA8yaOSTAlfUR4vuBFWfHINSmiHehbQ/Y7cLFv1
U4DqAUFXRdzuI76QIhjQKE5NNdv9RaasklWRB0XTp1opyFnRp52KBsy15xJk4He/
NU8WnNzSq1IgVCZ/zyk/keTMl22rvU62vrTTA/1VVL0NpucQ66X/sUr/6ZxYbwRt
I8YpNAoS55pOLKtMBuZ9IkRKTA+SRWaYSWz3kcg2W/kWBh9Wl/uruSQo/EBKl/YI
PPCl3lTWiDE0GVhtsNHzssvFLho0jxIRRKfNX6pwmXXz1DX9say5PEsycna+wQ/+
oWNK30gYCLM5EQpWLmvWZdHqVfmNQMOcBiNI7UASPHSvao9SxubTHaMBvFNyYJpB
pCfhN2FecQ/FlPannNdGFKtZ7xwxYV/cuMcflwCpYAMMX/+CDfY4jd1UWh9TgX4x
eXzS061QURi8YoV1J6FPalj8nzE+/zVwT+xh+kmAJI3lqgyz4T8l3uwivNJvEbH3
aITY+V0DfV7ipJf5ohVita2vUXtvAIal68TpmQ0TuLrMiL12BxdKNxfeF2msJj6T
a43ePlfY7YG5B2rsuLy5EMfnWVwXDFek7I9c9b7dRw5WiCohd9S8mH44HPNOEw1c
/TtM+XMEIYiUkxOIGKKcV+IKgWcHnKpmvCu4wIbU9cQh61HcX8K0uNcBztD5S7Zb
Tgor5DkIp3xqtgpYGDRlM1SJ0nO4AYms0YI/rF3D07TBH/kcPBDbkatTgUEUX5lj
js2DzHN6cy4s3v8B+eF6OLWQVMWOADiSraO6Ov5nvhVskPec/f5+o4VQqdkSG3Go
/Z9PL/4ebrtm+C2wgZfc4uE/Pbqf+f2jkaxd7oj+nUptPunDwKdllbNEJKPCEukc
H1aw2Ug1liO7IMsNorF1Zcwtv+/yCAU8doqUtAmpNYHOYhGVmpG56oQATp9tNkRs
CXXJdL8rrOmbbbPUNFCqeAj5HHoNgc4ucY4L7Vq1fQnRVGRz7Y2jH02s4IO9vFuV
yUPROTqBCQZydOKgGy7qXfXbiwn+BVyM6STfGkXBnjbv2Ut864B6vwQrAWVReePr
J4fGHwRbunPVh3z4NZghVOscoZbyEyXAkVLauvYP3EE1CJPVfavrpxu/sJci2ieu
4VE/O3T3D2IOS87sQEg6UewrO6yL/AkwLo073Ke8Op0ldFzql78gmUgcmOfGWJ4q
FX63xX1uu+8GALOy4xwLClMjgw+m18EcSR3R4cqoqzTERCQ+74LNiE198bcTcBO3
luQQrlj1xFyQnXwE2XqW82d0BLU4TvZFe7f9GRTYwU1AN3+/wiY3PgNk7GuJbHVc
8hhWmSsuI4jc4ICQOtgo6Fg98ZzuTC0x7c1nLw9wvd61moA4olZeCHXizagjZqaq
dpizrhhIVpwbnlgs0Fmq3zKrHnh4gGe07Xx57OyvPbLuhhayW/JEOTQxIw56m3qs
zlGI1Jdsi54SQU0ahpYi0CB9JOnEhnXsfmfxrKdcuP0hJI6EffPtU3UKqeIpdign
+kAHB9mCeze9Bp1itjTHyJlf4o8/Q4vvdmsg+ENT5tVAC2j1MLBonO3VScdwzz6B
s9TJWyN248suEnUt1fzUUy0LUFflVUoWzXR2p/gLqzYSaGedc//2Onqvxy+CWZAt
sVzdsysB+NC/eKHshborMsWjhl0HuBTiDM+O4PLgUmmn5EkYd3tMGSxcEstosUkq
T5uNPK4HAqRqbCSLxAsWzRIbt0IjEk7whl8suiClI4uSGMPHv24u0JTVNQcnO3cu
RfGvsJUK+xNH+DUwSma/BoXsj4uEJRl7PlzGFAHN+SaeBgv/T/+fHETDaCG+x1mN
VB8DUlFLZGFYrKmz2YWVIhen9Sjgm8SgACcSW72+ncW317APIaMjMokcEkK4Nraj
l+8ARrQCGLS1v6WQPGkQYcffmadxUhFEOXdQpzNSPONLkgsskQER0pErJfvytPM/
2QV9u8mPVcnfZ0l12nGzY4A3GaHQazjQipvmctikf71iur+lUsiBQKLVPtdoG4hd
9wuiAcLtCF6O0OXFZ53s4dLs0XJ5V/epXdvxGrJTKHk4MnSJUmXuZn4QzoEJMEgh
sGWZFbFY8Ko0uqoB7oJIaAgAhVWmvPYCXIEUjog3i3hk2eQMO+c5JOBhyftS9+6O
jQzNjDl7oII+AmJrQCi5/lYk0ZAzE3IYucojh5Cajr4jB92sNnqCcysZvBN/37xn
Zutf11RpnJirRdmp5xo+6iwpZ6SxxjmISfxst9b5UXSDCHSG3ckMtAQTghnA89Um
YJMrnQoY1XxYOFdUvmw+udwyUGzdWxiF16sJcHjDMLRJN4qzVCSpdCRrclW5WlXt
ary0sMWcSi9ZQfXsQV8g7M+j6wpGLzjYAFS13sTMIcbnttpfMzDbPbsj50Ut7yu6
F6+/1W5i5iFyE8dhEdL+vHWh+0Ke/HICVQHQyGeq2EQEQvym4360+w8+t76kuIo5
cHrY4NjmYsjPiHCByHHMEUj+TJrY0NCRR84EyJ25GK0c0FJVNOJRhb3xvD7uceIi
dMhVCb8rLzNcJoHzhULyZeNz6wcxHkK8/bB+OIsrszHe6XjiwrYewHpHHTsvUKlG
ZR4j6pCxHVYKY2EKO/kl8/K7vVepOu4zB8B6lMyBpbPJQQjoivPq7nTwMNtt7kyi
yaKhdEoIcvZaxDU8pya2rxRSyzp1jgzMvZtZ34Gfi7VbDHxicjeKLwOiBem9d2Z1
nkrO7ptEcrUDpQGMEMzG6Tvfijt90VsVLLh+EvWjxoSY/4KMqhsLFI/k06R3ZBS8
cwKjfWDqYKujj/rivnQ1OxEUQkAbigTTGaynzWjEQQPIvJOjkcpi3Cm1p00lyJUD
D5U2cBNigwc0MKUPejx6UX2cItrnwL56N8UVDPxca19ybsiTKRYDfO1Le7Dup8AV
qWqqB/MTsJPKByyxpLLKAyrXG0XgyC9rF0E6SO/tVZno/gkTzF9s8EG67+ImiXF2
ON8UdF2VWEfTBhcDOGcx4co8zdphncyQp0qCGkOX9HbDpKgEkhdxEQc6nk1A/A4c
6X4ujoTPaAmVWBO+sFovLuUpcvRQ38VHAgA6hYoRlGmoe5G57TVXRQhq31qDyKzZ
88jfyUtWH8Y5VE1JCwcTv0xsY/QrBJoDluC432kXz1XMtccvckjjEQ4pDLTZ0yoe
6lDHCDIVqfsHbEdaNvmKJA==
`pragma protect end_protected
