// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
chMwfU5hKX86AA29KCbzaI3On+vOY/vqZvUx1GGb2E6XfHV+8dPracT1TPQ0UO49EvzScKJ12wEJ
GIWOp6AHa3ssL6JojZlrL2YIvYAxylbarvKTMkC5fdxmaL5Lr4drZ6Uqea6M3DVSDDPnq5FOapLf
9UtH8U6TIzxXf/6iYK2NtJ2P+WbHEDBZNhw8PiJtFeeN4Hh31nCjFuLxybbDTxtynsVewkw9RK0v
Z8XwDC6mG7M6m0jzalNDOr2nMjpBTSBue1jxhm2gmaYieKNFELPVg1wHg61ka6b5yyN/5h4huUwt
Kv9jwA2i45vDZumt8gV+PYJmXKuybiJsQX/aFg==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
sm9wjiqJaNHN3YibPON3f/I9NNbIHgaIUMb3XXmvFxfGRced9mCW8Xk0uSVXol0lmOyzxrxW9256
vPJmg9v8lsPrJEEsENXaymt8aaTD3VoreznSuuqczkRxiIs1hVvwF6zzO307lKTE6WQuLDe0k+rE
KNBedMl3C06qqnSQr54xvezNprZRryTGkA2wF0p4DkjkBwj4DA55GH9M0Ii1wprgKJLSud9h4TDe
3CayqvFUAqLJWKEYht7/yqhCY+99/dFxRC1mwjeqDqyaxYEpvOeEyVK/p0tS1UoDlNZhns8xY/T+
xPFNwfhdjlVxtREi7bExa3q2JNYMC6Djcskc5xYQgipUL9z1j5/Fkz8C/FuTlUKDZO6GD4StyOEF
yxqPOmMYSxWXEuFqPQr7j5cgUQWHCKy8sxUkb8UZ5sz3+yj4vJNrrnO+R/Q0r/km7JZTY9jVXlJd
oqGG5m9w31zG5d7Oj8zXJbkWMuDr4VkIFPZRwCD+qRsy63po0WRv7r4ruXlipoKFIq93ivzleUti
nA9Y6xfAaruSj1SONFstMHKF1G8o7IRTHVe1OR9dAO9VABycLFta/FMCCGzFkRyXzwFzsaXuiyQc
yHUKPaTW/xrqdrvPv24MehkFB5N8dem7KbmAYQOmvtZCJdVnImTfcnnZPu+sO9MViCWRVbG4TgP/
IyD1OHuqwTldr4eE2ExdaG4h0E6l0OSnp6Z8rsaJWLjzf/foQBorqIhfX4ta+wUy1wJ/IKUnDtGR
EYgZlOidrAhvmAal1RWSLpz/RsH+Ulr1oxhePHitdG6go4eIoud7ayjTFOVL9+2sJfndNpFdV/UY
Td11jLNq26nWZonA3m/0jZRJIDqbiTteRaD0DZytsSYtL20NBLzxCQ+xpqJmfp8fSoH/0BwF6irG
DbwQ69SIZTTSJI4oBiqKaR9FXIUuO9nogVSn2zPYaCUmL3BOv2F4rCUcMeoNnfR79c7h02rSUszD
8TdHrfoKi2N7fnMwszlSu1LGaDu50fLITa39CZFGbmEU/bqibiukk/yK0rmOjCbdz/fPPOTr7XLX
eEBNpmismb0uA4WqH7l0O8jhbZRTASjG/2PVCrQlDJgPw2NWUovuiNSUmne+zC6oanmGuBZbW9PM
QfVokXuH/bjwSek4ojyLPp5duDWFa1xGTw+r3xH2EiJtkvOjTZrl/USUAMwVyIHY7vHaB1dvrcEx
I+CzUTg8MBOFkEeTLNcYv2yvdkv+UaPmWzWym8Aj1Sv39JrD7U2CcvB3IXacN2eTSOXDekDmQu3i
NII3Z55u6GLUSvpMXmajco39j0DqDADjpHhd4M+xLXsBXResKIgCp9nO3vWQA7vwxx1fI9mg/bNw
+I8o33yrWgg7OrFD8hoZZJ99dUq0bmAygd1n2yKbQInBNc8Lgvv99xg6bPS42K1veHPDrYqxXQVk
WgeAKJPm0P5Cwo0fwVYVp8xzvlT+z8SkHCQhAJmq/eb8Pdn2KP0Nhy0PSru8xTVW9XugK7FAy4g5
D5qhF+FPzuB/rVbwEaKZO3FSdkjG4BWiLFEcTSxV44gE5NpudA1OfTKZImQQBWUvo/mTpyNEhJg/
epor0bIAnQfhHhVNagLsyReN3FBLBi5qcxdpdAgSecMTlzZjjqjkio9GaiT1KqC/TOJoeiNtnTwJ
0bhn4pOvhnqFiqJVicdIyFu2rc2XvE0cAkrSQYuoODlSsspw+iygT0en9KPPm+Y25bFvUFG9Ka4j
vbeB1rgKj0o38tZxrwZU0tuWI4W4IhuhhNniwPKBM1kJrqVa7uaLCb1FTxvjxlLHrnNpyOXBv2YW
8TvsThyBPwqGYis54hhc1JcTOoUs+5QCubfN+UkmnRn4CxnbmsfswcOtxQ8jpLAXgO/nI5N0iA80
ovrUeMfJbaLve8eRPPcUMY1CRpuGAbhwskNB7AX1LG6eCtdiYmUwtMMXk9hd9a8iLVHry+8v6wgC
sPk9gDZNBz7upa9xSGdFpGZg7rf2uRKMRaQhkx11bAaTIbzgaiuT9iozJAlZG8WoCH1SJbfABQab
5ybshnJ6+adpogGfVmXlLgGx3DwiSfJrrGgVdd0eTZUzw4SAO+9CKPcon76HXf4DVspENshi2jU3
x31bVxTfO2vHUMgqQYffWMKR/guGIVUrmZcxpe5ieqNdgFhn7ts/i18UuDAM7Woy3SHyF1hrpEVm
f1ZRyCHNYPBPv5ZWAtQ2SF8IXTDheMqB6Qec75uQZSe4vO1YGfwqrRdr/Qw5jKSjb9mO+FgO5QRQ
o2ZeGwjxrfZpDi+QxoRVEJ7gq61g8Pk3s+CFO8uUanzxslTSKqu1lnRrZ25x5rQyBDR98H618ODB
6VUbz3YQ71UFkO5k61M9VkgZPvU+ODFnHdruwTC7hQ9uQao4CJX9Q5bXOrchm2P9OI1IRzpHmDRS
CFtgkVbIF9NERKcCzMYvdZvmLoinb68RPsbu6yW6cqU2KtLDqXx14wC7UgyEAa0rfBmQUOUv5mX5
8W5UnVuToWCOglYpixeygn6WgU+lEpkT5QnNKbXuVw5SXWwTIblp1f2k7gbjR2/ORjKlxCjsOXuS
ARwIPFHwB/mLy65HXjIhnXcRDwP0gzBbiZvcJjcZMocE2piRyFKNtqzve+FttWtLP+qINzU0eY/N
vWdVvqnaGA+oMG59v9NHheD3uPO7OHZY0+UR0hVA5/bPIYUf5PYr8+2aCt/qX3ZnJEmnMb54ljfA
3WOHt+OAAtmYEBeNMaHS1ko1msVv5Nh+N4Dt81ysVVfLagX9NiOyoddRUBXgwxmAbTLddgtKi0fL
FhZ6uHXGSl2UuoODECYQV89jWg07G6VC/Wkzfeo7LfaS6YHCXouV2074bkpNCFY0lgq7nChw/1WS
haSsvHyhQahER1zRenQI8MBYpzzLGKk+Nqax7S51RIYg0vpDllJ4RQs5oWccs/sKozfnF5rxBEhA
S2lVt+222twpTa1lZ7HTsR5d+8lnPAtY+fHxu8osJZG2ER0Ia46hCJIOMQsIserRdV4csSOkgztr
U+sPFN9h6MXdkJQtv8cnMTFDPe6qIw5Hr9v0WSaNyGAabhkEKzAAK2NyutCs63aPonEG3INAJo8O
8r+P4axiUDdf1pvDfyZdQlYMd7dBm5ONhsOZbAXgWdFzeVEhjTv2+iuCqiS0G7xo6hYDEq+UxhMI
IIb32mgMIJsf11cRCfKC64lxk3ib366U8p0oS+Pn6JvQF6Z59YvRWkegM/V9fNA0gceH2CoeL/LK
nDbPt81DRLW3x68FgndwmEJPbA7wgYsTyfPLAZs52voD1fda2JtSTGebsAfXup9QD0QFW45/3kj5
wfJGb1ZUzbZXtdrabJNnfNORQ04KAqdUwjpFLazdxjDziLzEoIjUwe6jYSBpHCRTRLNo//GBmdWZ
Tacb27N/AFHQJggbo1PxuW6AJ/Vw9nSy3tLhbbTERMlVoFUqJBfMAl3iu+WMA08CvY8voL1VDGSs
CM/Z7FnJmheAZa5MM7HGOvAaEYLLucCYBbidLGzoKzdVmjTfHwYZ4RWSHbVg+oJ0W7h4Z5s0HEjK
hsmqQ0ChH0QVzQz2tleRLctgHWBR3u2i2OFKjmwNt3m6egKh44vf7scZnO3frD4eGrVHCMLUsPZ7
zHr1LwM4wGnVWGB38K/NHOu60VNCimVByNm7CUZJKL1z7gGWXCrgPbNy5zXfowD8OyfOkKupUBrv
jKvZ+YzCqiWdFMEbSOrRUcx3WDCTgP0CBATGtPTDItohxPIFRfqnDDhsx3mn3WUV+HBqq8+v2UFh
3orKScz1cw1KKkzPyHDWLdkgUOIknwlyJ8R+nOCX3d39kHBE1nn0yuB2RjFVeSfghjE/vGA/Lmr3
RXa20Q4aWLQG8lL8boslnXNZvgeuPkHZxLbmF4Nsm64ftjdICPZzUGkumfFdXcPkHXZJzxsLXPQx
ic2dqprX5+7ahKuNLDOw9VIABcfLF0DRTX3+kPvrXwiKRRKVazPfzw2tlHmneB/wXXSppPdpNWzc
prp3W72IyYIQAfXdWrgAnPHUMRXbjRQ2EZzZG7Ld1/5JUYY6mVnyr08TyYvFQwiH4CUsPwI6AWJ8
nH+If9glsFOCkAxGTxJEqj81/Uo7qoKv4woCGoM5NAJblytauFxJ1IpFz5YrLANldkVrAcaI6oHi
sqWadrMZqGpM7kJgaSUWF7dhuLzRt0lRTL1x8huXNSyGWOubalXctXhUhI9BSpo/egos9SgkUfEp
KsNs6m12FmaGjtAP230OaXtQSQwXbsOnspBOLeM/fKc6e19PcZAlWETDyBqmFdtcrOkVlDTem4h7
qbduO3mTeIcWirXhOjMZXGew8H+xc137jKkqFeqQqyl12RQmr8M5Hq/2LUHC+3D6tpI1ES8bluzp
+npWhI/dmyCmlQ7mlUqsNW/MxlIGVn2Uhc0+iXqOkeb1sef/iYUeLmUp/ITX4PNXz27k3M+JO/9T
CWHvixDX/26dMrWmiyMlB3yroyyee9IrX6KpFsJwx4LT8G7brQ1//PeLteE4i7MqH3gc290Q3Ceq
4r37bNn4KyAAWIXIMUV3l8bFtWp1xQJ8vLe0qxFeoCxQsIeBaz+3rOb+ZL5EQLwPGm9s6J4TnPkL
PZhMJ/GDZVfed1aaXIvt+jLdj+A3AYdjfaEoKqiVHuhrJ26WdyEtU7LnTrMjWu1io7APC9IyX4XU
bA4nHDcEroZg+PWpDXOxPjRLMMF0aSjWc1YEY/nxb84Xi/eZdGQII0EI4YhJRUu8QRBuHwUUpdHD
rwmvkynyuuIN1MdW2+P8hHa7cugUmHWjzIznnFvY6VUlHm56KYtF1ZlkXMKX91Udp6aA+HqEegny
IoWP7CVKJ93QlH0ez/dSL3zMsAmS4ym3bDcaHWSPjf0QEBC39F9qvr8BojQ/Ks4Cq74lpfkBTq07
n7E3RL0vHEBZtCPU/DwjaxH+9/LAhltJ8O3cXA0gJ1LRRPDxiDIUt6h18t+4Yrzgp6FiALly4E3C
t7PUK+NpR2lNfUxynYWD4+2J7ZLZAWtf3jcPYdXED7LZ+J8qGIz6wkKqKV5tAOWSjaizzKw5Zpwm
Pi/VphcaS6nmvEdLI8BdqBM9DMS+olCgukfZ2Z1ErLX9iKq06PXVBh9I1CNQG1I/BqqrzoOKt/OA
0SA+/QOTP56d1kDFJG6v8KeDFpIx4Q1MuOdIeSEiIc94xUmna/gDvQQyfaIkNXONFAVjAwVaIQZh
dGpjvSFsx2A5nLEv3qJ8iYBi6YClTerHj/pOcXLO0ZUq8U8RUDCU5ejWkIN5lmDMuCZncKd8Ll7z
kcjLbyU8XFEjg7e8FXJruHQ9yBxuktbNghwB1tN9e2/FBJe11wsuwofS2egtyBHsOQsJqeqTWCII
tllfpzQopUeilex7swWobk0RIESavEO/IjZ0s89h2q39zaWzPCTm+8gX8qpvhBAba12Tc541tiFd
+sWjL9zU0wmPvRiAYAqzO+iBtf96PjKeVBdM2EAR05OaWGRq2gHflqQccyrpLtl7tNwVsKQo2vD9
w67XftjkwFTyTHmPFBQ362ntYeenfTqoDgMLZUPgrWuJOTSMUPj2V6rOVCJ56orMiCtCCpedd/R/
o9lTGAGR1JhqKjNHMl3nkxNOTxdlgbyFUnL2PUYOQVwkPt6Q/PtNE0+XtpagwVozDYaqIqd8X4De
/7kuslQjS3NBQC+yKA+7DX+7y+hkxL9a56ttsAZ/Qr958BJx1lwb1u3vwvv698bUt/ZptoLyp81z
sg3RxwN6nHzjI6g6H5PmCraqRJexKKCUKFqVog9+jDIVKrRP9v69Uuem3ziPHxrYj8fc8rHXZuIg
ZXafNt85vk/ICgELXKG0oEshreDTo5toTAxWISEkrg2U9PYm/RaqQvV1CI1RLSQDvYka+JO0MZMJ
BD11Y+T4mY8cu/L8ZznYlCyjdHvN4ZvKK0//FTK1pyc7hHXMBVb7UwyAtAmy5DwHgwOr1VP642aG
AsAjeQyW1UGABOTrxRlMU88xfq2VxdEwb3mCx9bfdtZVaUS72ArT5mRgqq2TF8cLj4FFNOgjPHlP
X4JJ0whkgTJoJwHWT79uPMs9kCBEPf2Earp9a7OzF1dmjsbJEYKo78Vq8jBqyirM/Ks30QVSmLSS
rjfQBEYRBIW74sfnqE9sjfX0v85UYMyFWtjSd2F3ZvBvxtzXqiCFEFKmqmf2CpJ0Eq7S2WF1kYGu
vl1bW1p38aJnV5uRr5jDvIgrDFZEZtl1dmx4h/x8pRZefD1AtHmK/rxQoFuExoGZ7aGcIHsjsaeB
CCqIqeMai7uiReBeGeW0P4RXC9OJ5YNt0cK3qfFXkhokFQ0SUldu95LaCVK+8lGkfUON0yEPKL87
y3csIA7DdWN0KvQm7+D6J1dfkzUty8g4z9SCmknNM5DAWAYzrN3Oo5oMjoc0AdMv0uWDV6VT9/o2
YQfFd6zf2hCSypQpwVJWtEyKnNNEb921A8Zo9J6yficW+z1WzL5N/YBQbyi7zf6EU9gbUnCwZ31H
jDFp4mNlhk0Ijy/X3ZKutYHZ0ZAOk1io5+3dPjnIiGScXvh3uXeYp9jjaqfddty4DNEy0/HQz2b2
1KDBg+GUg4q4GMwTzrAGXb9WkjI9J3zFSA9GKCxXlGye2Qw6rGX/diGjQ1ade4+fAVhMusJydDjX
+UjKrd8utwIQ4NyrtdpDXF8/IAsTE4Oh1VvfkqcQdlNQfBaw9P+K+x2Rmgv8EPvNe/AKhOKDVr4y
FZu9P+mwQeFL28ShSLipjISMl2exkQ4AvE7Su2vGMnB/ezPVbeXrriYucvKqlSlAa7057jvwQS1u
wilT9BM1f5GvoW/xmmuknO72JRhNpnTYlSvkQRYsSJ5ALVMXmHmgCHuYT0aByBlFOyb54tQ5QpIc
AoX+QJZ77RMfyGz1nzf6u8nIk4RXhc95f2RQGSwIHe6htZjwh7a/v5SMxaGIO/1LSomx8meIAO79
cDDWRlWgInaQoRAaXV8eOSEahGiJYONV17YFOE65qF19je4NtBqktE/vtd+vkMUDigDIJI9L64lI
vBX8qmfDQcVfnC6JCbxN6aj5p65sBgCQvyHuGLqEuX0onLWYjxUZch+NinxBAhteupdGzhXNJ6q/
cxlEI0krwGm77nP0PSZltV1C09E1Kk9U1oimvhmNjRlLav+GgsjLLSHRhR5ydJxvi+0MPNhcZpta
Z77WcPkjUFTgVg1RN6aFpG3kRs0YTQba1RMr4wDGFDdte1goI78NLDtFAkcMMs5K5vm8uuX61/G0
F4DzflgHvutQ/jh/r2UZpa4HadcXhuWOTbXPjox4rGzTSvq+0n7fDTZqlGtYlJuygzMUSzHKCQ0U
kP1Ovo5+vGybcBhS+jWLL076bcJMVi7NppwAQFakM7MR8Wpw/9YjMtjv1zTYZTsxtNkVf1DItI4r
EduEp9w8EtWB5e28SM66DuRwRD3R0vCzftsDAEJx3e4s+uFnCYxbcUujlnhQNIySzIdJ5DC1vQnM
EnH8Y97L+HUKkXC1QbT12OWQsyJvy8fpiWITPZiAZE4EWSz8InPeBGZkYe4w5PGIsQQj53Iyifww
BBaFV3Hbw19PoTJlXzpsKoGP2HSZuYJoA5mXcAUZJ46dkfinEHGISBGe/hxA+0kMsqYRNdRrTSc9
oKprgNWDJb8+DQo0W+9ExeeMCg+Uc0CfUe0n7yI4+Jr3tMx+ctrBYAP1UJxa/EpsZRawra0R3fgS
BK8+LEMKBRkqWSbDj4ne0SQK/uNO20TFqJmjvQm6ONnkANDx3ktLyJLisea/uOdxnSObQGSqBFk+
wCHcmY8neH+4A0vzmvurBzhEN2W0FZnpCNYockHcz6qFiAu6JJrVlwTYD37GH6+frL8HvpZu73mW
ZGvdb7o1JPyHFWQBuZghJQHbatEXFX+kvmWHax0Gc6DOePqvyRZZcimPza8PWTYIFvwfYMmwGram
6q+kucqf88+l/PBIdRfvmi6YymxCbvFci/LQIQujHu2bpSOQOUGwWFZ16NbUNIyfUh+WWaiF/Lhd
gwnjIht8zu8EqjSlsaz4tEz78Y2sdQvoeNgYfYf75Qx24AJYMxs4YSLFPH/oHEBh6bn7+vNAgr8A
XH439yCEgxbKLQoO5SGpgWXaCDUOivQT6PhFy1seFUEf5rm0f5AhEVTQAeXxyUHc73ToBwCEUB8M
B8ZF6ERfnAI2nZ7HsKdD0S6H9aA22IpGtntOQZxSalYuq0fcHqGV32SadyxHGQb8CsXKJe8i5Quv
9XvTt/CliE7LZ3PSDA7QmN1Yl3qiLAJctrH2fLUMZd41oCYiEkeETOnRdesDo82aMoND+gHRxKDU
16F40bDnGJMKfsrhLrBI9OWISj3UebGyd4myLzIosyamHKP9/88bN9ldtbz3niXUAbM5LxM9ci41
ClZF0uLFbe9Svb9CDDz4drRsCvYhzw4EGBoTSXdXPauyemNOZfjc8p4IL+Q+sbCjjGdxNzYO96Df
0L08k0cyjMi9yKykPEVdH1FxmZH1ZqZ9HkSbT+R0JYXGVku1HPdZkG3PksV0TbD6kB93pqIbllgd
20n5j9kMQRSN8Xx+pVGkh2aana6dc5v46O5AXhQaGUYf+259fgwlwYQSaNzkHE1RxjDdvuhNP8vL
lbBEQlQr7BchLwIYGidJM+qxOx8VQokSMQe+LjhinfiLjnR+xKDZ62hbuKBM9WFnLDtF7CtD6vtX
YnqWkcM54XqOhdNX6p9kUJ8166bmLlx5jzWSvQ4cyH2KuflaYImE+d8f3KzHdgPWn2poPf6KRKgP
34yOhXI9fomhCXQogAwguDR5I7pJ7FVswowoxJRlq6jj3FqBidrMOiqHC4lQe9QLVkG2qa5w0fkE
Kx7rhpv9fUf80EXuEQr/j5B+gcHCkbkIqBpkLmpvTkWlpIuNbIp4FwoLpXklgX7UnfM4a8laKcA2
qFsH7l2kf3/FhYPApwGPgUxvaBhPRfTiPd1/UJ/c2DLjzwhl42ULJ1pht3b8XhTpIMew5F6FoCRB
MaYbk33PRG5dsVPLDbH596RGmNTlM0W4l4SwxgWgpyNasDW4yhE3cjwULy1Nuiyd1r0wmnEayRhM
lmpJ7fhRyUTLpBAztFcs7pNhdsLAcSn2Fq8tTx8AG5vFoqDFqeJ8mdgYL5WoBWNsIv+p5G0U9ibq
2KvvP0KJ/P1iTOJQUlm4i68ylVp3KwT18HyjBPUB5118q8GrxenA7ngT/hpGXxV+DP9fW3BAFC6F
6080+JYHTtM3BEH/aeyRBrO+JBCen3Tmtlh6lzjOaMU7XGfmeUoeZkT8r8z+8JGSQykDfT2hq/I8
t0ZrCs9c/aILv6IX8D/yztAY8MCwTCSMgflVogjWmlB19gJAxD9b+zOvh6It7whJdFhMM0YTm0bl
2s0i4oAeF02x3JLjQ6tL2oZtAUnnrEBtIxYrL//jiql8LDU4rxhc/wkjy3sU9Q1KnA45YRvqRFFu
pphbuKPNiEsDSDLHQ4n8o82OjOnvDXSbdmHg5t0fy01GKky8/CsaVwz+J8JAwVa9Dp4uzi0SKq9f
uNrusG8rz7bU0AnRXGs0bMRbj6LmRnGBcXYsygEppccEqB4yR1Ni3aNv5g8vlNjgBkvuzrztVsYd
kePpg+a4ZlPrAVrCCRHcldUn58xGp9q1D+Uk9zBqqBJFWB6vSKOiXVqB01vR3FzcBbLAnOwJORFD
pN0iNm6jYl9kus5kgeqheFE678u1LAOkEqe7NtFDn/NfkuJ6tcqsi4ZOqJAIsl7OazjMs1Zb67yH
Lw5aPztONyjzkUN2fBYW3wnY+qrnj1vv1ELYNUtq2cKm3Kp6RDe7cnMbBURVU2acr8jTZr8sGNF0
MyM7nIELxO+bjmpjWKGVp+3sqAhj4NC80sPvg14J0djYsRA+8BgUQFSzt/JhdRUMeq8iavV5V9R/
+o5kolgsN+dZprMpzA+9wVcWsl5VBXyYnhx41xRXdPfo2NiowPCqp2NG134jFtCUxC7UNS11zUFW
P8R6f/QG39RvjDdv56aF7x3ZVphBuJo8DeAU7gczkOrABxX2dpgtyx39MWw49Vubv3CQPZNG2tTN
uR7m5i+3C1Y+Ykw9vkyfxsE+X9T/T3W+F0sa2n4TFw/Ev467w843KwyMtB/q86RH2Eabe1VU0IHe
psZfOrlxRALLIjjbkBO1y9OZDfNWgX99ALiq5wAA1BO6IRDu9LVAZWiNONuWKkselUh1kS/elPW6
ieEkqCTuCURk8pcAtvTL9EDOdgL70RVpQTzhc9lHehBRU9IrdsjruXi+KzBVYOmj7KpuEpCe4HQX
cg+UXQMHl3s3Bi5W1sCpQMTSS3YEVR7voejt9KFa88WiZl5nLYJNeLXj5dx4S1vzzv+NToDlLYfu
aL4VoN0VZYrL/NxL7gzrDL6r/aDXACvrJ/WX/4+j64Xy2/1ObQumo8ho8Ya6Br27W2KwnBVweVRK
NYtMXiX+lmUFiBv7CrVy74Wra977Lo+oZcukYi8rbZ4W6nhXPnFR6nMP38A7vQ5WWYN7owN8haTH
YMmv0kAmVLDMiM+EzU1T8PfBPVzK1rMWxU8IMdbEPnmNPwPxWhNwPgk2T5R4jQBWsPvKbdsfdiER
w6KLNcz9uBZ+o/ONTci8rsCXJe1AWkJSl0ZBL0YicR900ai1pELwGrek9TlyUv80QYs2AuFksGPJ
JfR9A3oMkLQpdGnM+jT7cBj+IWmj/voommir/J772cqZ5qoPoILwpE4/2qS304+AA27M3oy3Swne
ep0fvNS9I0CdJIT0jF7fBreMPWtthSxcKp/m7w+3BqhGJ2Fa9s4OkKQYP5/iQRhFbppMUia6+94A
JYU0Oo6nvUE1QdBEcG44azyBvSpqE/06KgqBJ1yEJDhij2aqJBeRO0Kt9+B68YIwhHMsJtCx+HVX
w+SaiOzbqF9v7dPKZGaP4ikgxnORfAG809mNgkR7rsKM6PbBcFN5h/mJH+tEWD0GHXru0anartlx
5NtJEGMwklv5rj2x/peF8laZoLbcXc1oM3xJ2Vv9qcSD5IcenCcNWxxzS9Upg0W+PkxMZktwfzJW
o3uZpUH3Bpemmte2AufUcsR6TLLFEvSyOMoeMxW2FXmNScBltr9rpnsgVsDF0A6BopzbzvepEYo6
WsDpzU1fLwHkqgQ/uLoJ0xgwilAQzGqR3RQYcRq2ongYR0O1kk/JCKX1UQxLNHKk91ASX1iVSH9D
ZA3mzXXr5NrgR/ol0ceHNRUJBSOujbMl8DEFOE/FUaJ8PRFQWr6pFygBgwVllX21+02Ujqm562c5
gxjL2NBUkhoBBYeqUeoBQK7xztZv6nt6en6m1CrfQbrYgpi/YJYQk4CZ6gugvHkvxMgjp2fuwI6Y
NeB2XyX1IcFh1letmBdvlhvcD+gZmQxyAj0hDwsKCYHc/7ZMx1gbEjt2UdniEJqZmxXYmbAh1DN2
Ks7tLxXAKRJjczkOoyTTZO40k7Qp6IVXhOHhtUAMCw3a+bkMjGDzti7JvEBiJG+aSZ/K4rGNp5mu
GWJmHnjfmEKo3PvSCfkfL5BsoHE3AgC3X/x/jFdav2VpolOUJw5CDTijQY0Azshd8NHtcFgVmfPp
LdohMCsCbknqrtkP7zvhTU8LQxxhp1EVrtL27VBySfTSNPnYw/6YBQz1t4v1RLiYFUNudxFWycg+
fOd4wlh+x8bAIZy9buPYSrrlrhE2sLAHqEddACvVmVVnA/XSnbqclbM575Cxd85XzRP/pcofbMB6
Yqg3hSImMqN2bvdNfTqjj/bpPfEfTZUsQWRNm/bHvCXwiIyS5Xq55X/WvI8xA7hZ/nXO6aX1gOzl
op+BvUKWJgd/2rXe1uFXoz9G46rmfYaPyQToi42cGX62sU0kfTwVALfuQ7MX5gzvL23liQH8KUco
r1V9eejwW4hvZJ6tRPcBa6Uhq+hKFxtXu9AOAbJtpGyRXVQwXqOIADjfEUW8dhYy+123ULJ71Cy+
+IRzEH0iDJDlkemdLp7pZKrMaS2i8i8xwrO9WDcdYESgKsB2yln+Sl1YyzyZIX9+279PJg/FRGdD
KNTABXCucWsvn1jvOI/DulEphD63c6CpwULooxZ+AiIyZtOU6ePyd+Y+1TEfQ6ETM6hC1NuJHb9e
77G76Zess6zLuZGin7+qWfOxtd4CZIAXWQuKxOBdAlnBc/pOOoQNnVvBOpAzmHrMJY8NXxenM1ik
sWUctfWzVg1/aFwduJNEp1EXvDH2MR+cYWpt3Us7OLTe9c88gOxgsb3Ip+4MIibK/iB8vajjqe/e
ypS7xScewPNde9j9NtaU79J4DwJzdSTJeqsksUbqHB+AqYHBPT6ugVkG7TNxTx3Vc4icSXRuzde4
xx48dQX5DL8uJhbQPv126RTwjuKgx58iJzg49BhXCBQIWy3az6TfxYjssNbYpSmHDPKH9qajSLMT
vWQo2McRaEQmMZ5RQezY8vfxDEM/ctLHppiyYOgoZsiXBXLivn5nWReTpz8wWT0hcpzztVYRCZlx
qg3tjrCO/XJnX0rd/PAiSQnQWGubg30mKOIfQgQVPEe9BfV3n+RNAI7ihd6y2Nk3Z2fdnFDIaVtV
qrNaZ1R76wWQwm1QaB7Cr9p1q7oIl+T1p9tl68by7n1fAQ6qszo2D4SbQ7vz5xQPxOy5AGVkd1EM
+9PWoehS4c8MaryYPqp+s7H832rttudntLNJOuzfBcsQi8cXIXipJ4eJqSdHPh5xRzPZo9gPe3W4
axGdWgTzj8zN9QYuhjXRypgCYnTrqJyQNV0KT22uoFucKB3mg5UxgZRqp5yjgXcFy7INH3Td5Fdk
tp9cMDKUQVaEYPq5ZnMbbA0atZPyVbH4JEJXEVb46M7ahBZN9dxgx7LIGV1vMWcNPq39qdpwEpkI
o9oS0e3iGsg47HkUFqj/L/eNv1OgXe0vldRg9Ag9sM+nTp6y3C9KbcBXXlG5RVSNRoMyayzPOsXK
rV7ZzBszCzQE58szE0yHN9fpW0euh0wYgDsSkorTz6P6vNvp2kwoeZtXjWlZ8Wv15VTZpm192dGL
Kkpa/MlYsoN9hL2r6MivTlRwAt18iQ8vEP3ZdlM+AvHlf+zICYmuxvg7H/mzNAURsQhKapB/G/a0
pmtX4Xca54hW3fg2aH7ORSyIBut6hjlj6JzELvkVRrwzNbZUF/I8erfFS8Mkkw84Qp490lOrGHHa
dyQWvReFnyx87hAOoOtjbrkO8C8STavg02fGNWR6S3WdWP9sQGNZfjPohyuhJoKV5uKrIFbQG+/6
uHb8+/OiKj4RtQV+nXg+BDF1IBJjvSIq0pV0q2E5IsC3piZmx+SyrDRGrMavQlnimOBunp5zPi6g
80eJAFwfX5HB9LamCcJY2Q7pAqhRHfXqk56fZaQfo6KaeB5uWdQrJvVuTQ3w4HV7vSTmZnBs4ZxA
elb6p8edR7IJAjSdpfqQfekwnhTi5IYrMkWaEFbY8amF4HpKcVzx8TuPgq4h3RT/H8Uv8/KTgeAV
KuhsFSq66vEM+bxGX2L+53KyHiC8qzkmLknic9pholN1ZFgl61xb36xUoNRYFoLdp0kPe9SWv5zC
vGosHJ8ogGTpdufhQNV9pOUwWFUdwq49nlm3gIgDv8ef1W4LLTinJDK7ele81t6MIK7/JmC8gEX+
Jq3FfQyIk/P7uzk96ASn+6NvRAqce5oaE7DsQnghIvOz7wAS8/KhBdy7GT5zAOII6+8mMRKzXRzu
CQ34O4wV2nRS4GTfr+latHdwF/1F2ObbOO5GAkFbY50dbderwyzoXebnNOx6nX3rS0z507NHVwZt
MNnMFiFbzOWqTxSujCGqfSDA8P3Ty+ZdQ/mWGcblAgm1ELTfcMlvSwLRCVD682UdafkKUW4SX2hT
7QhZgfxWcy6NkM7gt+j7csvb1tBEo8/XxAKuIJaWosojIDcNXFCP2s3khNQgTW48tAPwptOcfWUW
YVT55EoTGrreuQ4+wfu7qCdXHllxMZ+P3nLTOm93sPbt0lhTMWR/GkbG0DroZa26rY9xjjSMBX0k
eZUxfZw1iij0fC1zqYn+EigXsVPIoRrtfqDptJgbhpJMeFk9co/xpVXaiBO/URjz2eVlwCqiWIue
OXYNDB0dixzpD9VH58jxJRoWlVXbcExNaZ4ZoZvBLtIAMMxi2T4Gciimxwxs3rxnl1HchI1ye22j
bt9BxO5TCVQ/gmdwkquqHZmKlkD/h7GYTGUHqvncSdz9nKl3nUhjF6uGLYvp+ZYQYGbhC40i5wbZ
42KSYjBlyckccORVCSnI7mwynHCP7ZzaSIQNu5wbKYdnsJWi2dJLpKhmiHhUskRvrY9jnQxipWo6
BS9v0a3ZYyvUbzkr+kE6d+KCNRqfwS4z2oAeNeq7BPoTS3lNyjYrPERrir3kG2eq2DEL/kH2IMQF
X8PQwtUGjw3Ru2Z2ziSnrU9TldigiK9oke1nEK5GDJKv+ptCUQpa0pbmpvKcNWjY2mGZT2VdIRjs
aJLiyRr9W6skT7baps/KtVg4y1B7WrzeGs2/Xf4fSX1HhmzjpVFr8he1afSPvdl2vbZ6MwiTgNls
PMB/u9RHblV8WO+lcVKmM0us8nE7i3wrBXOJxeIFnZcDQ8/8D4ubAetXr9VK+f+T6snP++G784+J
583ShbTv4EnOZe6Y+SZUrubREtwIRexVJqAxIX9J25dRvJoI9YlaLW38dPtSzXIleNcI2bdNHZgT
WHhxBRf5EJD/ejyjmMfTPIyQ63mjU4EcWpUWzB1I0+iR1zAXwSrwlXjFN+q7rSsUJXEkZHQyfRDm
q0/actvYml3Rmws+orkFiytl92eqUvJr/1uM9Tbspr5eYy9Kz1T6JN/VkRdzbk7YODdD5fK4CGE7
feOVqk1CFmS96gRijCSCYU28I5Kjbxrdn8qLi991Z+pVdd8SfiPUwpI4fLK8w6JbgdiaAh72SzEM
5mI1ZNbNqMvGY5nbZwwEoMN8jVZDrYrbb4clhnh7LIBQkkevHhCDgsnBqyGFvlpb8bpxYxaYr3CY
/9jRSeh5nSkIgbu3dZTeeTLI9BujVWGrOYRypQxGaSMBdMkPJ77egXKiQZoTR1rwSxk/eYEkZq7g
lVHpz/DKTV+1lDHza+XK8j3BOxBbK+OcmTV9sjHRIEFcE2bhH3jnbWh2HR7okmzdNV5ZHke0VAe5
6stEk216DtojSv78foP9w7VYnfqyv/9DxkqChBB7dHNHsHzfzoHewLhqxiO7HceMlGnMFjaDcckZ
HylFCJomIS55UklQ+E1zyZdJaAz93jkVmFfQdeRHOpoW5g0EmIu9fODoQ1JYal90Y6lVk4uWMyKz
lpfY8Ll7PbsonvUrfpdUfnZQJqBcRiUZMcsFwI2qUCWC3oYBEjrw7+X6xzPFe6UPx7l1KfzEoKNG
ItrfP6B7NjS03oIKo01wjvNYi/2MrnrPd3wq3pQvDrwiv6esdTQM0f/wdYMa1uGw04D9MDkbzWFG
qQt78CnsrPvjhgMdnWDRHC+oeMJ9U2/i2G97khXwiD/sdZ1PYrN9UZUlg6z6uOreLKf7Sw3+SYn9
9ABZiOD1rW9FpJrkUZPosJGUO1d+pUaM+gHwZJOOwvbO1myBRhIeEp3ObxX42wKUMh3NnIA7WlMO
c0flwIM8Fzr24ew0Hi4dJ55aD+xcjGEGuBvUc818ncCsHnrI3gFy02LbtxDY4zttySyidrH0SGjD
8jI3scuEqkX/HkuORXEUQm8Z6fbcYRypJRT1DgzE65qcD2JPcSTGoGSFZDak45/I9hWEe9q0a7p3
GA3ETw6e5B50yBFrRQJcXEPblZDzXCmlc6JmCunvy2sL96kl3YdO2M7/N+u7qrHAmHNiNFzbk715
GIclWRCxPkPrjbRcnBpEcQhSIl3LHKiP4Kl5zDgezCSeuPD/GVKqvxSwcOEKs3/7AjUYtwGAwJr+
sUMbnd9jr/hxBdx0OgBZ7/I6ihct7nnhVmSa7iTUwIKMNL3aAleec2HJ/Igs9AIIdLXR76y90oC9
qTG/mEsXpp7sajNZKJDnN4OE7tSa+IC9FIa4YAbkksBALnlaUnazzegCYrsQ87NcdjnEl8AjOFye
9/3qxBAjWWWSA3mIPlRUZ3Ychy+nVro7nt9I02BwnRCNHE2G1Snwr9b1FZjnni2vUjwc5xV8bmNu
0JsnJ24lv/H3tzd5hAFSydbYpdC428T6LYRuTMPx24PAN4fPORwPLhKKOkwLL1lM0BEGKlikla9c
4RsZtIvXkPInA1UDYnO31Nr81QLY5al+h7oIMfnC/qRzlGLBhFtDAjg7wXW26ybK+/O5LA5Lj88i
SURZC2zVsOE84qU9f6DiwPhSPBrp4T4XvQRhGiyG0tdsuOnsFqqv820z+TLoKj0hoYUcwyUTGqqf
ZLbgNjV0N6MQGYvJL+GGV8vvvstWyepeQ0b5zPXyw2XTKMW7zylbyiqba8HcNqvFYjVFhFljHCr+
yN+IiHWJ41A61MmsS4oMHq2AIdv6UJ8ycJudB4nmzxLJZSSpaYOnJkgoEhU9aLebWbK7SSa+Cmy3
ghhOzKc30rjPAtIBPl78EPNbsDlTcmGxw2vkpNnxUazyWL8LQya5o8v8B02lDY1yvi9+qhHcbNmw
KyICI+nIgCuEefj69vKmrRBcRb5nDKh2W46LLf/QS8U/B2Pl1CpbyaKKVsFF6X133u3p8Bjv++ir
WkD1vmob74j/scx1KYre9e/sDBSbjxJuAjJuREFUsrsFAimZkw2bV54kMsRxYCq9IzVzPMZ8l8S2
x7CjkfOpX4brQ70Et2WQ9vrAghF1R0059yEURshEt41yV/d2uIkKWi9Xam3Yty7657XiMWHmWy7i
ffwvoFN2GL1z0GhJL8KzDLEeOsZmygN+30F0vklvInJhmcBcdB7m8LyW/KNU5RrBKwEPx9Q8nKmf
zik9OIx+WepNzJl2UMUyZTd6jlkrYwopB0XejgLxdol17pw5gQXKwLIi/0LRJPK9fXlJdNWQ7pC8
0o3+JtYPiDzjWIpMK5c4awLTZiDo7f+g535FTKnQpV0/4t8851pd9/Vf3xINuf8ovSlZoBxPecAA
q7eQVqrg3ioAn847dIPhg9asGgRQsIvHmSZ6ulF6j/ZUBL8bCBm1HOqV4a9xuIQksl2TmgW1jJD0
HWFq0ecMOjoPXp5nVjhLT4EACTYGqsIHf4HVELn/PoXCttpwVyZGm2iLcVr9VkaA1d5ncSMbxcpR
he566Pj/rlsD1Obhcd0MPTCcaguhpiBAwCuRcq+TgxsRVhfWHzA3K96R8xKifswQML53FASCFkeu
hM+IZh0aOXHKRz1iVywF7VeN0kAusC+Ry1j7Wa6E0X0xQnaYjCBCACz7WbMnt98hNU7fYfb3QYWC
lONILuveD+aTwyYihbBhfftTvSUYx5m7Z6XenA6eKB3MORgih+aNq4hKUkL9wOFZ2zhB9MdkY4wN
n8gRukFzVQMo+trP77VHIF2lKHecz+34z3jcJnTduM1WOe2Cv8vZlSRFFU9LPQ2pXWrZs93SRbMq
uqHG5DzbQmowJ5rJtkNdtPsS8CeFsIhbcv0gp95udfkgb414nM7ya/gptnC2E1sdR1vKElMnwNEk
Gt2Z6q4meW3zlQrnW1d5vW4T/1WSbhf0lYfRmml0faiCQBNaxqqbw0EavTe8tX3bCtcVP0ABR7WX
eYhVbmnh430d/PpWVRmw3alUucFtSjgYujrpHukq2SytCLCvweeiYrW8f2vbmMWa8zQsDUZPBmKu
p2hX9sQZc/aCbrZVdYTOI8o5UC1iAr/QXCDwONgqFxktoAiV4kZ1rczncVfLH9vf1usT1Z8Fcmlh
sKKC7BDZMfVkpE2TIDAEG1qewjwkf+ZJpk1pai4YO+5L1ZwDEc6abvK6pqgoHTAsWQknHZ4ymfeE
7F2m8Gnkzf/msJOqdxoGWoKNaDp0ytBIkF0A5jW9AgCn5jqaWPIEmcyaG0vmOuQ9ACVb/D/dWEgP
2EWo8kawg7ValzCF4mAdyHq7gAC3f7ry/OL0nkiAK5RGgx7pIwEBkbU1WQN0bXp8QKEoIstrIBZu
IH0RUo48MbvrPuDLZJKf7z5F6FkDhzbdvD77aiAAZwhtk0INv3Z6Vj38DpzkXZTYXX39I96OTXMc
xc843F/itetdRh8igDyOgYvp6+MzNxvuk1oiZFm85HJ6eT+9JoyvmY3u4JTNAKhNSZ5kD2dol0ya
NMKnVbI/uYz7Iw34ZPt/5n4sj8qD+gyuoMIyfbNpkcQPapOkCHG9BmIG6fPiOltKsdZhYV2rnZBt
Mj2wXSekOCmEn2zS0rt3VyT0QfRL2yj0rH2Jv8qCbehQbbmxadhrA0frE+RpMVlPp2D65wVHJvcJ
3ojfGyeAODqRk9MYE8uLo3gKZKDZC5AgM/c7LI7u1YhWWI2ltYHkhfKEWnEsgPRSJu8ZmIl9kwWx
jqDirGmhjmzT3bZNgDmZqxwkFlVB0PscNpY3ZUwcjk5ZtkJr1QNiztR0dtan+rVwTcQ3ao83hDdl
47i4X+HQml0BlvmHee5BghMVR4tt6v2+Y7jwieUyLjabQjHNmUS/b8sfZIO4XnwEkv7AiPvBrwU3
0nTZ2Sasa93kLbwb2JOqMM82l1L6kvmX5W+3QyxhbTvyBRwtj9aDTjX1q53k/LOe69KaAqQv97JF
A/9qpATzGcqiCI4wFeosyP6C54h5HbbpBaCwebGhyX0z1nSs4n5+QUfOpyTu8KERkniUuP+9g0NL
F1vsdPxB83X+AM25NO6bCILeS+bQqf7SoBY6d8BYQxOW9sJVThmJA83La3IAhHTGsJR+qYrn+7NG
CDeVugMzBPYxQ4YmvHG5DEhb0tajfnnMk0g2UCcvC2W8QtsLdoNYr+JzIWIwqMjAkjIipt8tJ3wG
eYfp5zZ+jqnjpu8sFR83iwoTaXLiPlJEtNH2kYTUUmU2eiyfgjMuN3FihBiNNLc9fhhIzy3ohnqz
OrZPNiX7zkcIaFPW1bogpm4ifc0EFH3HDntOGeoAXLfln/bL1C4Bo59AgALG60K+VhMpNM5Rk3w+
cVmj9E4bhI9Wgi/GyYfmr4VJOJj6nHOVAbl53cp2yO5p9fcCuAMkBoPog0WoZSN1WABFdKVEhAl+
nF2VOMfGqdMWpAFCsU8BB2Rw9xPm1dwPTlORWnf+2ersGZze1+CzUf2tGh3FkpXa6HNMj9KRaPsE
yS935O/ePniAgbC9YXa6wZ5DobaEmNvawdjgKOj4r9a77PzUManQKvZJwHYjN63wXUjCxyQK5+hs
DPCP8bvbu+GsFacnP4B2XFHLUlwrmO3iNhzcM3BWqsIyKk65xDalF3QsFiX41OHA472RjtiMFfeB
2JotQatdFXjTc8rcZ92C1lSVKYwPE3mDRdOuN8z9hbn0bgdwQEKLqgyzgor9SX1Q3+SRPtiA2DZU
If5zlc6tkfF/6gqMtqSmBLDnYaDaDEwimwzMyFK15LnH/XgVHrqOiZmJNI2ggTBVWbAEDmWH95XF
nQzEaIrROmtKe1dXrPpGL0OR1P4bmMOTs22qNKWgo1dEoMa6DhiCjqjR0NCuXiX6WBGaT+V2MKRb
PXvA1Dw3oVx23JyCA4hde1fk7edVDXxh7PyUnfLIfKqcNj7B1LxAu1R301d4QzpVhGLpgtIzPpDP
C7W11QVD7Eap49UGuT3FLElpkKERI+tcVG1S0A5NZezp+UuaTxALJK0Yl/cJoLp/GgEdj7TBioBu
50AmDtQ1lIaq3arxy0tSwB49veJ4q4aSbQQY+t9TMuAHfI+zeXBxUyd/5X4RbRoE44x+wN0vWU1y
WqZlrPV+jzxdM5wjxksRsih6pLxnpQXs1irvB8sAoDxBhayjg0ogonk9UBjku11QT9MoTD6fla5u
7v7K+HovQvU4KtcV9KeYdK51i16ONhNELuFJi7WDms5On4v+zctBpli2Zr4jMhqjUTPXrvislYup
sww1w0fJ3W7lV8mmaX8xxu+5TSL1zxVYsg43jYEvRyIwMi6wHhc7g6fjL48Ndx6wC8omSVEETJdn
G+ckjpNLSVItXqz4t02BfrGxbHNZ0V9YZs6+MVV3oLdUXGt2rAVAjQA3Q9+sBg+uBKooHGzRi2ZE
ZaMy0OjT1YvemTJRENxp8ELKujXaA7fyOmqYexuhEwt3sjoB09wzO/j35Aj0OF55yVC/8+RXqWa5
RI7bJx1yXhuW5VsSLPdSb+IjmmacUQR/jOpFU5M4syyoOAj25x8R7HzKqnEFf1UxABH2IMRforZd
YY432s6GhicTTtkG0FnfeEj9jteZrsVPxMU+x37fJ1qprcVBzFKxGSE+dDuQFHdPG71L2M53HfwN
8IytEErZCGt+eWlITU+40AxWYRV5DB6hbJUi8akvPnc3YMXmAhTpNOQ/eDxGRC1RKD4j0B2n6zBG
n4euUfI4DtaxGqqQ+yK5DZ+cbCWRSsDL5p3xO6cYcoIojUCza4Xvn/ahaFI9B0pY9Y6xgjtdRBGz
y8zwZUP2SN4Cu/3z3wtK97wtfZr0iUZr3lLPKswj8cgBrEAL0JfytQzbxMVkgi5ycDUr9K9mBqo2
MpWaSI4ktTxz862lrLlAZECtkxMM0F4XRPl/0lc1pEfgc2ftOOh1n1T56f65g9FMFd3ywZ+8v9kv
zMZWBejrReJeJ/sBJH0zR2GcmEG/Q7P2ObzFUDXx827SQdnaEThPoIK8drfhvhbfCzBk5Z2q/KpG
VI6mZRMfLkSphcKSUm1HfSOcsTLiMHJoZKH/DOls7gHQ1ZUBh3NUde0GFDAe6CXBq9oC3u/ZOxj2
EVzcHsCUOwt9h9J7sIuerUuR5fP4y099uTJIFz3z7Himb6XbtuuDxx4zerbLGQ15LhvmkI/vjkPY
qmdNmEz3eMEFJZawG8TjLS0Z5rVQLkHyCD+6hsg0kQf02EtkxoT1UjbkXsFYoM45ZYbNBnt0bk0y
ybz4m/x1YPEUkb/mfvtcQlxurXD67+mNjIrIVuSE0gsnWR2maLCTv6SBC+hsRlvO/1bAEXqAipmP
78OPKbhA5UVDzlKD1Z2BxZdSqWg0TB/cCcjgVysv4yH+ozsHsAAcADdah1kbxpzlBLOrpRQ0NPTT
wri73tQ8oW7+oBF6wUQPyTFke7BPAsmM/mLNDq9uK8XVKcK8OPHNohaBb2qTuaQzfxJR0fqiqrdK
Ci7eoxjOSSl2wr6XNrn01ZlAQC/l5xzM0jTS2yW2LXPn5vFId9qgd86OsFKUSvovZ4x0ZbNthVZS
aoefsLSER2gyaUx8aBxPXRRIx3+guiLCvGzXfoUssDt3tRyNzwqN32/a+yQmviO4fWcBUnu0GzRv
9gcaByuuK9qahF7GsMeUqSSH48RorFTkaMd37c31N+8y4k5Uv1cBrkFQ1xKaV8gyDIqsRovJHblk
EnkAJ/4+hnAouJQawRwqjP9jIuIMtZXvnMkdBJ+Zr7pTjbo53PUd64071nOXiXhw1p2P50PtXMXb
nazYfHkFszEJ7o+XtYrpT0jAac1MvKdmapqcRnAYL0+3ImnadZ1iQdVybqTYMXmiYUl7+zcOYScm
+2bV0mm6NZAZxaPmmo5yQiBhNy9OPDHoMwVwBa0rH346mw7FV1CYDqiR5k1ODD8DvNudh/BCLE74
DbclMn7lzlcp4dqPz0BFl/IGtiPNYUCJN9oJZ6jCcVIVI57YvIU+R9VQJTSmGV913YaXlJe/5I+i
+eiFCP2QLi7NT4xUy2fQ0sY/SqtKVTy+1HNjGfNaIFLyJEN1rgJOQ3i+P3dV+qQsSLT+XHxpAh3c
JrdTYkF65oJantEm2fCOe927qCS00hdT+S0wmm6NOT6cBBO1e3+FJ6BHCb2HpLKXUNltb4repAnZ
o8joRXZ3P/BNf/m8rd3Ei04Ndl2v36nnibMT4LnEeOvi5i3RPaaGTkaqaHaZStRvXAiu2xOr41jA
rjgt36Aakj33907LxxNbs2vpaMafIr7GVJJ14A5VVaV/Po2KYKnzeSjvpKas0FGCnuykT10vhw5I
ZJfBgdiP3XIOHYS3NZPUrUK9qhvG0YF8KdyVhNB3j2crOL/k70wXpr2rMtZbaeHAn+htlNlVHL+Z
VuxoykG8PS2Fhzye7Pc3LKL34iQ0+GGYjjBYCfiI1E2tCNovL1uRyOG2YliTZzK42olFJrL4qSBy
h87tIPCKJ9tus6hMpF5VpUhYNoIKWwgvsbycKGpM0Ttw0eqPfd+PoilocNY5SlwBN1fQSQ+zSFCz
Ed4dZe57h2TSQ4zK+DAKP+XL1WfJkAgAYW9ACW5yns+XGy/1nF4jzREPIIXkTZIX6jTA0OOSEwcP
n1ifbH9xaL6FAnn5AGsu1fwhLfPl9wccLpnhKAPjDHe3rNayjq5MUMx8fYnDQe92XV8NetGW/KtE
dp09ld4hcmLASPSgBEfVflJytY4qO3Lba/rDN5O0BWtrmDqD3DYKS7+G2Lnep0ssjW3dJc/ulH7/
tMptnOkK13KroL4LJxhibxA4Eq7JlZIqXr9yuUvWnUuLX51LHSiIYfqIeOusfr2ZJJ80Jlkuh5LH
dIb4JRROgTVBBF5zjZvIPqMnFdSqISO6bD8JY6oBEaKmr+2/1hUnMrXkdcXyVDRDxem2VUfdbBzS
AGAGUIY85zU0v+h50WO38JjQUqfS6R0F8QvAu6BjITutho8Q87DU7EwzurbOa7wjCaPXCYcah2Ja
Cm+wP62c7rjXxVLigbHLOJUvdneRR9L32AYklTGV8MSKmoduT7olgBXc7jV39vrMcNO/gSPG91go
saF6lyC8UcoZcPvgNp/5kLhGwYSs5gx0tN7NKiop5rUhXHyEMUShVdZPy/0bcO3VtBkNPCvjsfa1
acQTSoxpLe4XbPrPvD+VAaT0YrpTabogRNrj2YlyzxijoQ1v5TDcNRpv8Nwk1NdVdGQKOF3mJOUS
+uL+jWWAnoJDUR9e8WvwuqJ66eyrWqjyLunZPa2BBeCam01FM5+7HDVuPHHiWfv9I3HV8QGq1Qfi
4MFrBQO0F7TLkPmRaVYmxyTW5n7M+D7KiVvfDj7YIwuT5JErnlD/yAKELJ62MggskQAoy0qC03E/
v4ewozMhgKVE6wPVgKeCdzD7Txp461Sn3DqxIW9GVBv4zpMybIVsxlgIV8Az2Gf2sKC173tMRJVG
dJBV4nQBjUBOfGPKnXNptGxbpJ79SsjLUM/b7Y3sOmtWVRKOCYBOy19XwWicbREml7ClkkMUPjap
a0xMggLdgSoRSCikLBF4aV6Cb09n1TF4CaKTTNtkrATCB5OHKvzICAZP5odKJKZ63m+6TqGz4wCu
bVT8fRwT6l7c2rfRjDO06SFn5Wy0WvD422HnmNIQ1iOdE6dZc5MfsJApQbKCkUKCv1MIO+8mw95l
JHgB29aiTlFXHppxXOEbnb/zFkf9Dr/QwedkCkutb1XXZFV4KzUi5+ijLuPWl0Y1M9Br6L6sHH6N
SguAm3EczE4N6pJAtUx/2RGvWaoRxhhLto8CCRYurU5V9s6jr4+igDcxpb727p4QuwhZLYkAZcv2
piNhh97ZyrkUa/liutkeU5mRl1WDaB9Y97dazur0UJmQiOkgIqYZ1M63LPROwMHaDgf1uSuJhNVa
eL5SNtDybeJ1RDOUUY3ubTmeS5zjbQPR8tQpKz2G/g20StnZRELdlzRqOiVXmK9V7EpV6oInjWvs
ybNxbA/Ap9PHaMkHbvbgYSwYPRG2R+LbgEI4tOuEeVfOlw9QXE+3DmwwaEOyEUETGMEhRZNItZVD
1sOb9swUpHbGVS3sxVLOUw3bdtdEV74YOFDws8CN/IX7ouezBFg6z5xXtBKW+fJj8s68oxBcmTWI
SbaG/XaXdvjlKCI0UhFh7nan3kWgaEjBNDr7hWPTts9AizBlWm7krtEx1H0Ln5j/x8aeSAgaZPBE
CfQABvwiiXZ5NRdXyzcTvMqEND0OrJ7Ki1eVFWue4p1/relfuvemIyrwR9DFXEN58xlnSmxRmUPa
2NvJGz7b1Z1GZzDsP8GPmWAQtsls+ph5ncw8xylIVvgr/X7nOmTMpFH015aL1ZB9NqFYvYwBVHjq
c4SXf/6eD7vDJnrB1tAkEtPDk5vkMUSPSXEMdsT6Y6voELNvQoyj6bFbcyXRpbhA9AIH/XeWsilE
YbKnz7qg05uf18OANKAsN27FU6t3BvIWgBkvLPiVJ2fo8cgtAS6r6qZCdIr8+5YbWJXbvRSk7PY1
w76balNUZ2VdcdMN/u2Ur06iqRvrzcNpBq692Fau0Zp0U9p/uPEEGEMs3Cad72MTJ1oUsnJDzLCT
yVdy9123P+tI/TeUFO8ixPlGiq5VzZL64lLzURZ03oRVE65oLvg3p2a2giHjLrZbLFoSJ/D+iJDl
lRQlmaetnRQczH6PKuh8hjZYFj0DLZl1aTNFtDfG8SizScHmZniwv/RDO7rz8rTp1RwY4YtyXhdM
dbslzbRC1pMuzT21jzFy3EOnkMuQNZyzv6z/4crfQ3+1bSI3POhh0Wj0FrC24WRRR6D2A+k+6HeO
x+aeZQpqzMEzk4aewAdfjOyHOgqn7UD2VGACOOkJLQFulyzCKI4G4sw98IjU5XhVdE7ttKsEhMHX
FGUY1NhpiMACFD1EZ2bbqtKqQU7IClWUH7aeXx9dAw7E+bq6nbvY1IDi/0DaqbyWTSY4K1TVrr8E
o3YGBxpT6kXUygFaDtyN5XPfeZ60N1lIHj1c8VNKlEKply/QN/DXJLYcKEkbfi3yNaJwx2KdELYc
MYHcsht2BdXPWIB+N2aXOkZkUSA9GCtr9075bpwAli37CoK5fFgJe5LiCFWgHruGV0waCZHx4egi
/vpnEFimECybDwOiKdz/RaZfyhUofXyPTWhL4v8/LtGG/jDDMzjHRAveeSKO43D4GgFsqcSr3HQw
zhmEF9c1nU7Ko8DbLxa4XPfhlZ0vnUlfzyxUMXcnOelVV4f/eNoVTHWBBUumQnOCSim5GKTLwnc3
Y6GJRDxiUSnajKWhq+wJMjE9+fB8lwgvNBRucQ3dDZjl021Yg+w8F8UBAQKBUqacw1Lg3a0WCz4N
XWGV7cxdJ4Hzu/dm/OGmTkbmLHNt23nwusicXXJe0DvOw9cdAPLrPl/k7ou9pYKwSrYRGWrE0feE
nTbkcZdG5rm2FdqqJ1xuOhEuuF+sG1ty8h2Cy4wchqMPCs5b1CyT+V9dkVtcK1/BqPdQr8+u+qZP
/ndSqOnqMQe7wJO1yGecPlRR7HitQKJSFtbbRHIjZha2/z62MLh5ChqyCJBqHKzqtdsbz4C64uWC
lr6d0QKyaU2LWZ++Oov2HvnzqeLqvNfWv3RINXRQIYWE1YnlV9C4+rmQbmJ9APwGCnKZpS9xcoEU
HLHZxbcLhOpLNyiqqWD19otZ88ZWvROCOD3q71Pa2EKph77Rr8+MqdAcBgCRzwZ2owGZx1QUaVqj
DCkPd8iDLPX/Gi3LNf1/MzQkAY/uf60MAaMGBgzlFdPcTVHgT40maCb7m3+nuAlFzE9yFiVfU/JM
j/FAeYZA5W0n83l6wegNNX0aWHUGVhktaV5NhzfEl1cv8coyrUSuVHrPZAZJbtiMLZJ8jlRC2Jco
CxairRKzoYa/Ehm891owJFFL/eFqjLwnF5U4dKr7XGkoF/9dZRtDhyrrB8ySGei0YDNOys6oTBQg
4z63Sf0AH5WfT4sk0L5tPR5zRLf5lOY0MoAa9NSHqYuQJg+xpfKwjt66X4lFOx1rtov7abt0Cakm
nsmeMFiFrUI16rmvjpvmPhSCGBuH7x8lURo4pia+gZgWArrYEV+C8kUN7Y4CiteMx+k4NftPHWY6
oemt9XYjZUDjMqSR+0Qs1sWripv7fzx8/eemzOdC/AY7RNcJqA/xb2//vfWqLZr+buvJ94tlpyWm
Q1JE7pu1/thdRRH+e1t48aX5C3kWZM0lGuuHwRHLSYZHe19LKQ9Nse4bhMzSp+tEf38yOrCDPcN+
sZ9OnCtRFtaJB/sMhxIbMv7W5FIxiROF17fD0eU4SBljMDpXJUfspxxJ1c0uuoGEmntdlr8sG96i
LcGNIEQ0BA/0spgkURjx1NlhM+F54o5/8Y1/qIJV0vC0XMVm/qvOT3EmpOMhUu/QJDtcpUVDDq/Q
vqmqiMnMubvWzi/cOQvN7Thq/QU0B8xJSrqnebPzu5k3r7LktIVder3xE8HBb5OqeLcoGbZmRSS4
8gEwmCdPlG3nrXG61Iay/bgXAnB3QatZdjrhF3bR8yqlpGtlWOhMh+nYIlX6YLDQbidAUuL5FVul
DRoapXGf3aG4pYp6Wbmhl5p26Pd/9mGkBhGAr6oq8VNSrFZSfTgAeAxTQARKlh5nbnoNionTHg0B
DM1ScGfYNJuhjvX/0cObw0aUwMmRhAt/CTrUsOt6X3+hbn3fwlzbjAKeIWN1WsXfqhR84hEboSjd
16PlnD/DxnL8PyFFuSVbrNCWhy4dZccFr1D+cKNEJ5oNXXHZv8eKn1eTIK+OLurmlV8GXsnTmU0r
Oz/R3IpfSvuwAbv/gz0uSu3FIHVqopR0PBoWgKAxiSPtDzAR6mQY3MOkisJN3G4kqHpUT7jWf7Y7
wAd0O3Q9ZAWhQ+C4hMxF3LEN2xTvMwJXzYCFcXohK8T76x+BfNHzBBZPMDiboMHmsLV982qgYCuA
nG8edooySIwk0AF+CZNZQBQZaOtgE/15tdrJFepJpajscvfxsuxrp2FCwsUXbERRWrcLyg9rwZzW
ZPOjZyBg4yapp6ggks3SBF87t/wmYaIV1lN92gMZV09Mh+En7fWSr5jXhtBESuCKv+gx1g0xxexU
lWUDmQtIejzFeqX1LMtiY6N1vTj/KdigYRghtrtnLfnoMGFZGxRX5gvxIPmyCFzrH8wY6yZVoMIu
B/Kxlrvw20zLSZx7UFyN0CnD19yGqf9J+hX+L6LZQs3+7ZZTkND7mHVNsTX0FH+RFYHwAWhcNRaw
LPmQKQzGJzjgyBFkKllqNFaWh1WEldWiojB3rOfgB/e0Ewlej0vgAFTAN1RvjRvXcMYkFWyxkCzm
sE2oE+oHl1LBfx8o4Ka+eoy/74lT+psKeXY7HqCLfTWD16jccyhe2uQ80Wqag/doaXyKEriII/Uw
lrV0rCxic2/Jh4hpVJM0gjayp61MdaiJfZl0jhXK5I8GgR4=
`pragma protect end_protected
