// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:24 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
GX7nFJvkTNDAngeSIBDrgNw1/nZyODR5r4YAzvZPoV5mpOY/LJmflW7Ofag8Cltz
niAN1ibju4wc0dbszxFciPeHqIepi9KVP/9uvlEfaf99qhLjY76XC0hZSnz8heem
17BNilqr//PNVvWbrIomVCUoUYSQuUHyd6FfbmdiWM4=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 16432)
RT69irA4wmfXFDNZBVwEFVzLbQ/uWgH932aIOoTd33nufoblSZf30iMLsAtBTppq
K/ROOMcFCT6VQj4j4i3XSAwZqUL8T2KX3uu973u+2naWM56MtWyBuufEAoL0HRAS
IR84uYy47attL33NIcd/YuHAkgiIB//g2tFbe46+EQ2t7Zhbq9ZQdAbAe7gIJ4U3
UrO9GZOFQuVMCJKN8sr69SDwfjVR7RFvvBqII70M5FO/0hx5B3fANj6Ii5svJxfJ
eupj7SnG5/ptykHBA4ynyeu2iDAin2cBMcKIM8TbteKx8Ej8oJ/CXkKMPQPf1elL
espMsloJAaPWBt43PzgvWSzHQ32xMXlIpG9kKCjrntppdTqTuxORp1zYBRhVhga5
7yEpneU8z5evevNgKDFAxQKXgcY/mkofK+6SMlQLBFjQuwEfvvYXlPU5ag0hB0sj
254rl3R+6LPnFUFEiK27wDUHw/xx0t2J7PqthONO/hZikY5lonvMnCmfbZRE3u5h
DHmeY8JZqCrBRaytxp8n7/2qxhn3eKcQ7iyeDNWk2FOnz0edv1FzHXtkMCAEryZv
SvLQ2X1o82U8daai3V1sLk4250H5SC2QZ5b22oV8q3rOgj1vnkV/BWe5qPHAWjHb
o3qVzM3OXrJuM07dvyc7k/ra1lfV6yivCTXs3xkM26B/fkm+H5vO3YARMIuRzxSq
yRgvFlebBZBYU30VLMNdTrRaEgb/zSV2q67miFQuNWDJJTVMyivNa1NkTnfMMafi
+AtUejfrQG/thze3VMjj3t7kH6waRZ3ESQBmEGX+4/iEI6VGa/pZvdsuI3cc/zhX
+mruaMK0e7AiJKJDZW8wIm2e59ctNeJtj92oQo8EceXNctIYUb6R8KF8QyfdmchI
zBPbVuNCkqX09cJScvYSlqWmcoGILl8plz0t/WZ18n9D8PGmgUwiVNB1cCVAYX3w
uaY0TJ4But+F6H+CcmKUAc2tKc48XhS8YkRdM+a2z/srRo+TwzcaWRHCHMs0ZIwj
iGXEzI2V+5jQUQqE2DtROPOkyy8aEXB7gg/Il2Uvo2+BbcKs7AvtMS8Ocoh2W+Ut
Q7UYufYnIBuXBgara6Hb9fHyMyAgMXG+LG/g0k5++RPPByjlgdM42DNhAfxxzhZL
4753MEqt5Uj31rMOSSM6XC1ESeL1/J+2zcwy5DiZ0tCIa2rD0Zj+5/CE0N2+D4We
nJBTn3+Un9tzl/XB0J66/Z8co/UuPNbJ5CI47pKgJjLDj4Oya5EHeloFd8tA+ixR
qnCDYtXQLG9CBGnofmnF4I3MWBIcY1dJ68EQZAK5KnKv22RrfyjpRhug0plbBAzP
R34OhYE0OcUXumeb/jmPv0pRY1kvgv5C5jZrS6pTKr+QxfQDoYaOEIQTsa+gOySg
BNHO7M4wCO5WxQJnj8Oy7XNlHJhLCsqcYsmIc44f6sxVM3CZpnUVUKm4iATKbpXp
oj6MdGyvd0m2nSHHJCpA9rLlr90cZniBKTAwAyHX+xa8rGgKUORImb+4Az3J5j9C
CujuvOJDU0TqYlE3OrjymQZo0lcu2OqopZW05xNaou1a+Pkvc1ao13nSlauXM961
ZvaTnXA69GMx1d6KyrOrY0BbXwlRDGnRcVXDVsHv0MvKod4/OlhABBhHj21+TbbG
BMjbZgRpweIqvzbxZaykaBxDGiav0sgJXmUJI3hFY9ajhkl77z+T2O/Zb7OZm45h
wK9nJseCfYlgmvaZc6NEGXZ7BRXoXlnS6mqSONmyF7put6QCrOwyhtlmOWEUDjAX
2yLwDr7H/0yFD3egf1tq/KKtn8W9dN16rIct0fbKAmCttOglsI4FRpOIxM9hSm8d
TtLsdS8FPaHZgHIXUH78ugwO44lu7ytm9QfGfpNnvpAgKM8V5vSluri+kGILHk1l
jizq7RDhhIqFZUwpQqN8G1HCvzaG+HV2ZFc/v132tRGutqdRhsIdJrzLrAhIYIoG
YW23U+gEJw00TdQgMn3Yq0LwffW+4hlkndKgsEEVOR1U/AU8fe+AoPEkaiIrStm2
06DraI6jfLIxtAvE9+VTj/4LWVrDk2wSRhf3QcIpGh+rJJRn/53sPxnXqcFG+ijy
bpEIOrjySvR/YQZUoeRlCeDY9EPBE+JjOu6w416+UX9PI4ihWGoyK2ddG/H2l3Lj
KlzgCV8kMquT++w2pTI0pRrztrItVKV7kfpkarsT3k58YmXB4pQ1Y/JlnwLhZNUi
i5BF6bsajjbKUtrf8Icz9L8PsNjpUkx2V/MEt73Sn2JRsgTNKpLIzmfetjx4F8DG
YwhhsITkJTQR2cOVleUoP3JcxS4hhZ4UsUl0kkZiwIjBTUBfc5FuE6Os9TFsf4/t
PNWLFfHTP1iCE1XVM+Pr7URudzbfX2ONJ2Ln9a5dqev9ZRVAiZrU2h3E3Z7U5ixV
66aD/XxRFwfR0E6L2QjvjqKn6FVOCQd9ZZYR9QEjT2FVSewur2JCiXYumvNPkgzZ
p05xJg8EmFhYZlXiflqnW3DtqYuaRZMMpmAPljKMa9o+2/eDjobmavdE7zul0eCp
SUeQrM2RCvR3i/jx9hNusdjQ0p3llaH3S9TdMCjfukyPLU4daYo4Po8SR4dEy1YW
bMker7jnX7lZIwkllcPGH4XoIVIs/+yiIl9XiatUOR0lagHjV2NrtbT9xeRlscJH
LOPUUsx8ib4dFT+2BBG3GGSdEwdAYyjmw4gkUaYXTZ8Z4u2OdcPVF0HkeBUWRUZe
Gto2dAF+5K8E5ZgrrU1vzw7fqyico7MGqF4ZXvdVi9jeWoGcF4b7++i1WgPncVWC
ukAV6EXZdohxV+ToLV1akXdkQmEdEDEUo20WW7hLpbwWaI9Zkmo79JE7Njp786lY
6EaORFrhudrJSSsAaomF5DA8LDTJ77gC6OIkWoNRByVMntAa27jQ7Gi6Zj9rajYF
yOOW0sOZQF9FR3N+KJp0rYbMuLWjQAliZ4E5dCQr18afg7X7dezMY9uc0sNBh9lv
yLfVSzcKbFh/Kc3pJ6T/NMCpPF5BlEa2RQIlbpWRBu1n1ey/DJqK9BHcWF/Lr6q0
QOUYyxt1S5PhZKb1CqxlRFhsgXpaakkW4agXqCWtuNgY+wAyttwQ6VREvSYrGoxy
jHjwcDNzdO5ft2Xve2EU9k6DatiEIxyis24qTjp/7SnGrMF9ljZuLMmF1PIFiKNG
ZJ5hxZBwaOzg7kNQ2yke4KTubaaP3knox2iriUqg8WCGrKhLnfm4LPFoPdufgUhO
5Q1IEREaTSAHJJ21XSiHYLicY7wkwYv77c3GgGEu6aRZKOd2+MJcXMd45N6G+qoo
NcgrR2/IKINnB0yt+LFuc7xXMxIAm99s2/fvMYU3QyOJ3OpmAWAonBeBh1A+G9BX
gaMPZRgpOh5Gt5art4vG8/G2A9xkkbR7gz/BRYo2YmCNpQZ/7SfYw3zHEbs2/1pW
03kDcr0wT550xQWvXNNa+recV6YQ+p8OUQ2CQL7Itg4HCZapYjslzBKGyPfUbNrO
JAGreErvNOhLbi1zWF5ll0me4QY2lBKbwvbbN1Ra/Fo2SeBVwrha4vBAhr5yj01p
xEplJg00jjkb8VmHJb7RcXaiD1TPt39uJGXypEYQpGwoKKdFkGGApxD05IpOXUKe
CB3NDYEsdMtwOCZlJmFMJ1BrZMfyz20ZwLtZ2Ar5PN90L8+TJBDBb1vE2qlWkmo9
4jmdlkgaUsnPMSHIMMF9PWQvf8g7U3y+DKmg06w7vRFbLXMAB1f1PJjgszZatJh0
C+FNLGYZUrxqPpDsuHq+EJD7X44OS+vuvZJclK5LcBmhhgCCD7Rwesfsq0HXq7Sr
HNciJsLX0nqzM9ZiAuirgHQBv6vWR9RLbUqaha3iSLolB3mdll4+K9u8DLwSiXd+
mBE5wOQAxV0sA/iuwtf/uQQVGXsT5AfUaanClsRy1ondqQ+K/D8px5iHscjx24lC
3pqLMPNFWAM+hpdZyHkjRCRpSU7dlU8zwyFIZcOyCPGitRIfzK/5cH1R82YlHB3A
uxZXFgCnvTlQnQ+CmHq1IXUtHZnf6GzHIQwYOnNSpkNOBpLkDTGTSqxl0JUZmo1e
d8OEExp8t/xrAyzUdywqHGAqmggeU0uQp8Gan44BxwQemdFQ9YJ8MH0nX+kFpn+j
5UKmBsHNmzUcbfhHBml1slZQy59Zq3w3urvfIJOJboBST59mceU2t475O3vrp5vb
L3RFqRIS/lYidFnW7I4DSKUdqzkZ4OExzo1JijlZnk21Uhyc1GSX9XIAEHzswUY4
p5a7EgHK8a2b+LZEWhgN8IOEUDX2NaRBTr7NXwIOo7Y91GCz0hqyJEhMHIJ94ofo
ebTTvnMe0f4RknAhS2VHn2lyfFP5nxTE7zPhQRcyZK1YFvEGxfn7KdQ/Pw3hDQIS
H94QoT5noaN4RUaetNCTEGvfxn1OBlTNUfq+8fqZp7QUuLN/uayMxwsLvm7/T8mc
O9cjOei8nysB4sRDVUU5hzMuHEgIkV8vM2nxJW07o7AoWnM0OAOa3h3nhfJ+QPFb
/b/dImZ5eSpxE5HD8nWlUrUcYPHTJplcrNvdo/4FFofbB9td2NXQWHET6XWEcDkd
zNekm78YzooRPqSyz9UB/38uDzPjSDQSOjHNWpYmWGTX180NU66tkGPHXT2MQq/J
nTKEtFDYf8AME/U0fG5+VvO3YPcmfRQHXPS1vYg7uYcHXE/+2PqRPZIkUtSLLpHb
iV3U9N0+C7jslTyUpxhCPjz2BDauZjDZGRFGMatXKjcitNkI2QuNNMd0cnWgPP4/
hrPmcBK/E2j4Xg07sOT07bMlBfqjpQ0wnYbc2CJDV6xTpj+vJeuixgxYPovVwBO1
G/J+JKaUaTck5tjAUAY0E0OvfF0WXty1wFHGBANTHOeaOtcfk7xZxTnRGnllKSSh
5LJnJnOxFidWa8952JjqvZF5V7xyYPATG4wgBV/2KtT3jVbn4kB0gZcEBuqDtEhZ
SLp6r1j78vmPT+xLmk8JyE6LjL2gGnxR8kUNtA1kJOsETnwSC6pCjPyMkOpb13X1
Wc/eZ7Zcg2g71jRoCjtk7EL8OvLspKLojI2hPMyDb3PErEEcCch7lM7RlNO/FiZu
ibfNvuZetKdPQ6U+n5MT3XXckdAN3dXhhBB2kuJD1ymQ5TM+vIwlx5Rrwt2Bm5H0
pDqxNwih4ojlxmWbhBwdpZIFZKdlUzk0qxCbPqcOxHsvGXiyOQDedhZgh+VczN2Y
jRXIz6hyjeTXtIfhuv+SV4GOEkioGIntOGbZqZwUxLGc1zAneQ8VudNIRgQT7+Wd
iQq9cJtpWexje2B0TjtogKDS3Fn+LMolYhJoNRQP0zmj+SuJCtesdwDGI7ZqZEUB
Im8DMskOkD1fzttzdcbh2hhibY49qlgieFVZPt9iiNPheYiEp+GCbQP9MAp8Wbkz
sm0midEjpeVHLcLjI4UtecYbVHFjx0mGwfJjwjIF4O8gnFPKGfVdFv7DB4Ct2A1P
xJw3XEx94k6ejsH+pbKopNRqoPE9tICIVojzFG57nEMhT+3lPtE+VQHbnyYuUu7O
omtFZru2XEWCbZR8AHxfaNV35dLiN+PAJpu2RtzTK3YgGvzM0L6khDGpSTbH0b4S
WIHKumcCTACCXb/nGF51XPnCcmlP5nFQKgMIMcplvO+5a32H7RnAbUXnVQQxLvqo
AKsAljwA6QemTcPzBKY0gtrtYZSbaF7ZQ7kP/bEISVzirft9IHSZtnD/uWXVfEou
L2Jm+OSi/Ln8N1tXSR2reh7Tg5eg745Jt/PeHCukmHXtFq+HdxH/wYinaZOexSPx
w4Ux32wXFfz7ef7T2cmdN70gXhDMdSYs+wYmLliMBai3jkIobfyJwBUEanpRfHyt
CMFJb6CMGnZvVpWqRsIfeoq64cHJZ5es+/5H4a732ntmqTxRa/YObxANgb74Q5Mb
IMCLaLdMdX7HkYRrk/gz107hBdekXmfv8AMUR7spmcH1wg/5QLpOZeCg9HfboihP
6BG5+z7aTI0XVrCCjEBWtISgD+PN2vrNmDxBcZPACl+pbzdaCHfjnASABbn7hp/5
FjlWcr2AlC4yyQ+1ZKgnAy2BrKDEIC02o016VbcevZUE/KY22iC5EfhBrZvLNkFV
KUGvBah8ZeV9V0kulXf8rvUnmeY6oNhUq6Qne15ttbCRkJHY2feJJMpX1JzRkPYz
B+Zg+Gik+pBr67YaxarL2njPI3L4nJR7p/VfHZ5UTikvrplUkVYLBr3RJ0e1JPw4
QyVPH/JDsYPhLVFjBeqyAA7CImDzzyto7/0aExWaPGVNyqkkIZ0wjdqr+sG/L/SJ
DHChTduJLuGazFALUptEZN9JUz6evelNI3FEf978xHMw7Nbu2OW+Cliu9RYWIUTY
l8EVkv7bnLUFaEB2ClsOazfJxksb6D34VFIAhKzJUClvuoUWVX5xUqEqdMsUy7cg
AMaeBwuxqYHaK1AoW14AzQlTJgomn5QaDdR0hZSr5qn0JvpyGSj1xogtpZipKeO6
OgyT8LKXorFrTq5i3/Z6HsaWVlSdmE91WO8v6UzRpnsDUvjjwuT22WqzDkUK6h/o
E1/PEkHJYQBgAS2URzZi6j9l3pjmYRmcOvdiu0E72xlIaKog9bigW0Mv9Ekyobvi
r1+O40WPsNHj7HD31OxFEu92l/xqb9Jd3TbIa4b/BaJit+Brp3W7lFHLghXLLXK8
IOgpJLKbS68eytOmSJHB3oMoov2pXbvlzSbvK3klLqhm00h+6i1eSp0GWgZV/HHe
2qvKNOYtQrdnG6TLmCZ20CopOmgk4b8V3bAX8qHghOxlPOY4xk+PcSlGUusEuzU4
3jisNJ9ttFrkv0OrAnvd6T8qOsKbsxkfbXIzZ2q6pvaqo8roFSe9TKTTu3xFL6dn
Pvlqw0QQt1oP5OBlNZfMOzS4TgQoFjT6e/8GsIT+cMvbLGmRp4AgqWrGOOkIIzjY
ISlg9Yyvk5GtjDq8Aw92SysldENxywOPGs8s6kF0Y3L11IF9LduYQQbpAJUfO3Zo
1urOTKJWmdFZhWQOpUhMwN5jlyHXwOCZfSb/A5hslEi6V4RKN0z0WIFeS7e/L8VY
I/FhkRcq2zXRiOeuYm1X10i1lksdN3SNAmqgGZ85QB3mgD5lzklfeVvaxhNAFCXi
U4KYuPJTdsvG5EJ06wJD+HPNQL/Hl6SIHa6Zn9cyCoFHi/+38d7E//3A8TVmyxN7
yZWeGCN8Ds/+/lypc3gu0BdIkjkUOP92ynFwbLZeHXEKBbHjsZBGGLEAXxeviifw
+j4hfG7dL9QbRhHnSKXifWHMndsjo6OMXpzZKx32vXVvaCesByMxjxT5rZ8+DqIB
QXzSrMoMzj19S3ZmIjdSoLO7qHobatiN5sN9awb9ht7wn/rPS9A93l5hjbJCaicG
msXqw2z2ohJxCWbu4VNN8Ua6hTH/Mqnfy4POeGqwVdYIYGKxh1xur3YHzZapYo9D
PjRW4+e4LilRN7CxGG9Zr8EJCJVAfGWSe9zb67zMihVpS0fjSkm49S134t0ax3nI
7WKaGV94FXBQy8QRdjxBJxFUNyNhyZOUAcXZnCIhY7eH5JWWDhH3yXubkQZIvC01
BeYD5JBRiLIGt/eSoavuUP3JOEfHCjtwEnfLhrcmmXBXloL/zi51fFSthPMiGxwi
Qype2iYrbn7JPdXO3ujPs7Y0rFGX0myXwek+XDwy+GkqqZdOH3hSzGTPRJjnRHBs
kMQ9bF5KGZBxFy/SzpPD46gA+zpx5tNE9SHeKOqkcrHhHphSc9xfrXelFS1Nr7vd
vqYF8Ye/Xe2VX7jAgbCEmcd7XRyPgksjkPXE0Iec23ZbPwH1QqehcE5r44ss1Wlj
1ZqVPZSD8i6cvEfLXLA9rrdIIhCPZ3ZmGIND/GAFjYt+88o6ywhDrsyV2uMJFaOv
Y5W5W72i8KPPd9qcawAvlEnzwVvXCoauYVXy69TcpoONq6a9bMH9Rr9u58ycr8Un
INZHpSvm4HFc03VbVN1/4iJhA+yQ65VgzxSRTTpHM5ZNAu/iwHEJLWWcdOvFLKXr
JrtOFbDzK9BQLzwvwz1xbpSEho3D5gFVS7sTX8qTeNuJSgmtWRC2chgtEvh/db+E
7ZOQiGUlFiJxvrMzuOWxsCTOAWhYlUc1mv1vUu+ENY+HU6cApFVT97OLyjRGwllW
EamuIpnxL8I14ASLkiF03GAoxTSV7FA5vgl7Y8OoO9XGhgWKoyImKbFZ4KJBnr25
bLDIBJ4iJvpouvzMChf3H8XhCgBzNUaLc6Ad88LO2mBeN1pLZDe0x/70WcxQdA07
rIJdVjQGO/rRfG7QsocpFU1ZluLKsZ0vlZq5idOMMsY8zE4Is8sOg8Y1G02k8/BF
IsUh4rtvfH6d+HA3sV6+nMAagYs2rqdZ9GOp80T3f4huKVjAMphgCGZI97wtIBR1
FLqfyc1L1nWzI+cx+8qoTQaS5Bhv84AXTEYBxzpBU+O196mMS8pbRi7YIDyGOpcg
vqEsnsEeoOLVt3r/wq1ke6jsSZxZDnXp6xuV7O1h08cPJDqSSngWz2JYeFWy1ZNk
QaQuMTcK5vHpm5pzgIqpQx45DXcibAANFuuU3Xo8wAZoB2sqgPBLj8TKvNtxQMVX
DJdRlxOuLO9Pds1fNalSbLEho0/s3QWQxrTDEFtZIBZMLK2tzrIbwL6qkNWlx5DN
T1Q75ywjr/bzt1826Ns/vGeQSqKuRD5cgKsbafVIVFoJ7EomE6vS7LO451NDliWY
LpbT+uCSuVa6D8kR3kBXoWt6zAnl7zHaZ0tUw0QT1OqvCi6qQ2d6eQk5wggLP4ld
5Z62jlw1Cg56TCY7NRFsbnpyYWL3JQ56O1CM1cIJ3CpqxfzGSvDETlA45zsVlavM
9vyf+ZnRvd85WdsL4aHv11XfXtonyWoFkZUTkY8j4pH7bRw4FPEYworSFN0Xebgh
Lf/uOUyCkfmDcwkI7zobqWAGJlGuc2gIgmaekuyNIiydWQqPste8j9l7l0+6x9ts
2Q31IreeECSf8k5cBCn30LhfczN/4J+fjr2gmtLQM2snCPz4bF6lmPRSWdeXlNLw
8qQf7ZWScabCoqbY0SUTNlyQBjUCTqYMGF3QFiwwAFyiVNlLwd/99Vh1TLUva0UM
uU0KEHn7Y2MKMApJNmvz+WzFmT+LvRw8Gx2hmgLJGmWeNPkWCSTuECkxBaoiLjVg
txBbSd0K5a31+LmRcsPiqIkCSghMQe+GZ1+F6aMtDTfjotU2XMGsqgFSwKUZ0hh9
AK7qWcin0Ex0iCBjn1ruSmLoa3c5qkEhT0h0A3uetxpEwXh2AAFjSOwulKnQV5YH
3wTxLdwvThaEYL4pXJshlZnrfv4qMKaYeKC5HbFBjjTxCM3IobNkuEKwbubqEPCt
fLMAAp14H7ENv5ObTl6Jp9bLHIbAyI/nMrJd3M3VgUZ4LGzc/l4QkH5lf7Leebht
zyxaZgnlzf2P1tXGV9EOQy2O2Re/0Wi5QORdwDQAtN5tAgIiHT4h1dY/Kexr1sPd
2pUG1GajKnsvlj0GMTDRWglqxICk34zMfwea8Kwdb6mQ74Aw3olCr5AWNYNltOuR
cD/2AIBMOGw6xf2k2KBhpDq7SmMaBbUX6WWqC1FK7oYPoNoQbvFBmdEBPihCuiAu
ozQRVqzE8f46OWavXWn8qAQzupdxo/921KA34dD8z3iwMJ3DDggLz0OxAyo/BsWl
2kvTcWBnZrf+dF0p8zsBZEIUWr5Tpc/fZuIeAQIu+GrOgtqFt1AMV8xutkNzDYEC
QQn4Oo3f81/KsZqbNj8Vam/O0IsELeg+bom7IPd8tN4FWxqavrnVOnB94LCzNeRn
feDcsHjWRETZwF6W9TD+2YMsBqcz7Wb+TaYiigM/DJFTQ6qUESCyjX+0LzxWVVf4
9DHFdTeVTuqHH92DOkR1b1aHVJD9amEcdCM+NijSKLVOa1YyyBpAnPg26U4YVuJw
WFobJOG4XlWWy21JJ/bBdzpxyUPtf1Xz9zowZFi0AH2F1gDYQasBByxFWNB1GhDh
3/7ThqZUuMIbtPkwX0o7rwXOERPhUFTFeLbfhNuCun31fMJvMdOwky+E/x93Q3xu
OvgxsAzY/ORRtGUYJ5HyfMuG0CPEXkeNRc1I3zE+3MPDFDlL6RTQMcAdvaECSSBf
qqHC8MP4mCCXm829y/wwmXuXSWN8bHIsAbn+jN5teR7j33bKHcaqWQ/JCHw0tilD
SDjICIqKJePOgm8/zXR2sssL97KKzYPr5GeaMaefWq4lM1iA0c1WuSIR7MljjxcU
ZqJ1zca2wmsZk5xSKf/CZANnJZKOOSTzRP1TFPhrObzaIReUO+CuUYi62KoL9f9a
h4LQOJKBg0AQv+tAEtfqYhDf77TDeWyJMOe0e3t/4ECmq/Ua5ij/rKET8o3hSFyo
8u9lFCswDTyDSYfj8en0VUf4/yDR8oVSwERhJXQOhOvpZ7bH/L4HPLyDWEgUouSN
ejXpnYVFI1oOsuicja3rRJmS5XWTFTQXl9AV5HGx/B2GWsX+MxGJF6GzsiwbtBTA
UDzvnatUpCSRBGXluF56SLEpfdvTQiUhR3+R2K2wLDoczb7WFpBWArlOK5Eip6sI
qR0O7+eik3+GrK2uaf76L2jwRPVpn3NQ8FThNmtaVaURjzOpRI1fBr0+6BKdxFq6
bCilvDpVtmxh0sWn5ouptnq3V97PIkbt5T3eDsedfHNNDCNXmUAT/nMIbdPvFnzv
Bas5ttpgC8BWNQc2wWCmSht8IXfTR5B5JD2tNt+pJuaUBPGMknICpCq4MlRxIz6r
8wyujVpuYEDwnRD/I6lnkTJVmF46Mjd4JHHdqgJ7Z24qzwJiiWllPnuo6lAIVQiI
Px99n1DXcm1Wa5NN55FEZAwv+KQ1FGAvioamieX6+ZEId8iNFgQhXDINQDQNRJKJ
wXn3L1xXznJAyXp8jZNcwdSjcA20OwGf9PBLo7iTpbfnFRHa7X7lcUHVh/Xau5J6
r8UitCmK0Z3PytYeY9W5GUT2Xs3WahLseuny3ut8F9dkML1iAgoGESyC8NqJOFMA
flIo/DwGabUvFOvydWEZXQr6vC9cOMK6sHX/yuH8qKwBD1zXgyLbXeXySEPV1usW
3CqYI4tp48YLrom8BprPPSTwbe9ARhZvqAMQHWSccRu3/2L4niwZyS2NpE/N4Ag+
uM9IfgQ/GW2hifYSTA2DLF5kKviCyShdBwjJfGnHjjvOPIymzd/Ul50SPR0hFTej
VFmf+GDbUU6slxZ9jyknlYoqaHoapxhJUERfGDTmPjjy3aFSXopQHuFlDF9kMG9e
fZI0MOiZtAYh4w9ibSoBpOQ4GelHQsAny9a06FuG18fn2Th+SC4wqoY0Oup5aGAB
pthcQ2/n+dUdbC+iKN5iam3szSyCi5493dszHpwJDHRe7qWeCC4mNt+VCwi58brB
rckVupRomAxErofFCZ3c5EhEpiIPNS4E+5kgJna4YoscE9jhHKibcCVilTfRRkTX
F4q6q14XBTIpOd++bEKAOqBHujIUmXWhmlxT0U0VnKa/1IY4e/cm7Uu36TYJuuS/
ESh3DaPOFYzSpOMXYs9VufTUEP/LaD2dObltBXOcWsuWX3t/EcU4eS1NBg3bf8c4
V7NCNmnJgeFAGUoIPDcETn0QJ3J3RWPWe0NS6dNk0sM+fbdKkrmXME3eZtzYxqYv
IgtnSTwRhQiaBBC+syXjMGUxnBsRmmCAu+Gjt2E/97O3T3bdnjLgb6YYfZJBjKv5
iU+AK4tOt9B2PDnGyCdoOYQEXfLtDn5Jb95glGSKr18XqF/BDNvzjl7SdNLk1bxL
WpNGF+KrppWFjAfdHosbjJ+AJkYwU5R4WRGWkJKUiOgRkCxT4l7elxNCEyGL7/B6
A2I7pZV0WM3hmgoDBLdl8/7+cydV57MYuTA68muJswtAbzqZgoX9y1aC4uyU2LE3
YS7y5n4Uxy07PIp3IHXcrUCbkruyUyfca4DUGgQlBm/cz8r0MVGP61xEl70elDJl
LJbReF9iUFADJ20pb2/FXqnBx2bMrd4EcvpVtw5A2D7vg7wA6fP2l51S7FCSerCs
z9U35LSCStuTIV5V2mzclQkAmrX44Onusc4Ip5TuYY8RVe3xdN1KRG+3oVg5xR3r
+d9GYZ8hOMXxO8Loc79phg1nS/IDCMuk+xkFYxjuM40ZVJU8BHuubNuq3Qqs+Q+U
VvQqJ2e9YVBnOemU94FMNcygVZUISy7hk/sxHAtaRSUnRGH2GmHLSY6PTXZbO5rO
bLFwWQRXtMlCl2ULMZoJj/7mEl6r4myQNFpMxG1NyjvMq2Zd+ahxGiW13cJj/8Nh
MQ9mrResIUbk6yjqoDtk8hFiiig/JFTXtab0SNIuME5BcwY5j/f4HVEO2RQ8yHXX
bVsqMKp+5wMWXY57IRFoPH8V+zCX8VaZJ7dwBU2ugTE+Q7XP6qt4pa3XnSmRih4d
rOz79fO5ixbbtMz8MMkOEq8FLUHmUVFx1Z+5+mMekKofodoFUo0pmMvt3yPq9H1g
neM26+LoprFip0XYq7g/YabOwoSicZX3g3k4MAYawwUu7u3DboqWYmgrorAhLVs0
J3/FY0wSk2i0QWBcOrcRCmN2Q2ytSJXWQipj8hldDxX6h/M5NWmDvBdRzAg9LYy1
3ww7PmXF+fHimZSBICJ7Pi90BMc1J0gE/ifHl/6HGbqybuvvx04iklCb/PNaZ/o+
57CY1WxrMF/43s8WHDHfZ9iv/5Fuw3dhCBqoVtc9B0LHZLbWFXFu4cn6MJuP5mRc
w4BYSHnz6H/zTjkW5E1AYNByY6DYKCu9+etLMTxpLJbyTspFsjLXWM6XH705QsZW
md7oSjkXavLsTL2x/uB41oYCKhhqjETAZ/ykdI+DlgViv+/OS6221O5YWF+grCNZ
T3l4kr0tKd7ohGPBJGVpT85QK1PszOXIWKqGqZw8OYXTU1ECUbO8UEQEav+BeiHR
n2s2rL5I1DUO0toElvvusew4Wjzp9Z+UntImBsuV+9iyJDSqHLvwQucFoa6hg82w
ZcGiEh6MzOjc54cmi9ZvvbZg/PN6VYbi6ULXJGTA1fDG7WfvJxESFQCXLPeERzUA
nea740L18JzsyqYRXNDGH7MZ06IAlJ2k2NPP/sVy+9m1unaDnyFO59WRT6B6oUUG
CiZyB++U9KMqxL5XL4DrT+EGemUdNungIFrMf2ZztrbuSfWGWiNzEpvtcfy178Kx
tA3H6uO+6vphJoUXxfjD4Qnqn8f9x6I6McUak/FvuRqAU0RLL5k7SQnGMfTf1meh
iJOyRG7s+2n6pRKBWyFtj7qrtoPYAukwMAkrv41cTonr9NV4qM2A7l9qfuI5zAdr
Ul7UN4PrcTLGVkO20DD25GmZk6i5RY43XrENjwyFr4ubadJxz8NY1Rr18DIx05s/
mhXX+DFWTVTKnfEb0i3/gw/Mlt+u85eun5obPx1IbSl6v62l6YpF73f+KreFUwZF
b8knF8wN3DyngZSK2Pk815IriGxoGPXiRZbecvUiy6pKsMH4/58GOhxsd8qOXgA2
NfB+vql3Au3/4zHNOo7mSBX/QuVzpmtzOJKizhJri4OUbZNqH8q2QUgLozrhW0o+
B8CafUqocFxCTZqUfKOn10wGyOR3LEvoTXoIhgIOKDzc8kzJ+ngRdBh//MwPC6ir
JgRp5i+UjamEuIcWdqDbzzbV3cdRMJa2oMtQDW3rD8kA4phA2fA9Q2I/ts61PhNW
2cYjfW1B/HuKI0I0JXJjZIj1hp0Q7IwCI23kmFQPhPG0IUO0gOkQVYIOyNw9iGon
gnJhAsYiuSmaVzUfRwuqFcYuR9zHvTN3rdhoppzjtGeuZ7DrKrBAsyDy62Jk740R
ZsmR6U50zfJwfnwdpcPQEYns72sRIuYmGZd2PUGJKWKgQ9Efo1/NDdghMhXjQGZ7
nFDQTvwIyrEhHa/idSnVSstF/UCv9AFXKURnqO6+8UoyYz+wtGTOsNUX3MQJqJd9
e5JYkjsqOxc+8RkowiSwk7FgrD3WcFO8eXCipvP8OHER4ne0u1VRNEfuNyaflyFj
XRe3zIRJDYlxtJc/MboHGwffFEEYTaYIdIkyH8fksYsYoOOoJ3sVUGXuUMH1Ky4y
nCNMI+rStWZ8cmu/VHwS7uQ/O5/a8U609L7hAZZKDv/4OdUbHVtJpdWTb30qqtjb
rZNY2NJul5h3taO3QcIQNrzfAdptNdVhsnY4wl1XSpmI1gTsqAubhar4LukgQy85
TEDXwy1LhUAZUm4X4E66PnPby2hcwVArYqHgAlr1qUHIcmtq0BND2tLU5SbgrnLT
Q9KCKuUE3TzRKm0WV8t2qezDkdVw4rkCqsmMQ7qb+xYRxSO+CsesyNilJVGwCk0p
AbT9GnD7NUQIOcQFyDQg27/JOlndpJU3GH7VBpNnbkJDvVmmco96WFxVDKfp/95f
+l/x+TosAPCvmtYQWR+RAhB0P/dtplDUgdmPoGBXtSQbqhWgGPBx52XmZfe79jVz
9gs+bg8640sMEE+7ry97tIBrvWamBXhmRjYcdE38/xDiNFR9T8Z5mBRCgwHkCnTk
5qVXlyO+SSOqpy6G3lCJSGXh3kC9BXHzQyovcfaCTmPW+uOB7Nuvz0p6/ayapuib
r+TvZRBGV9pvbFhCSU64s3O3Fb0HFGr0WsI6W/GN/IDjdRyANkeuyvzI97a6vUeh
jyymjCOBBYHocjuKbeYhur3wyNOTMRFULbDEtT6y5ZVyGogeaBkE6ImlGCpfGC3x
Yrbpmgnz7NY7pjF+dKtxz4hIBhxvHiMq8OinW1M7wlmYDV7mu6fZ03Ef7vBEkWkj
3E58kJbo5Q7tjFiLEbT3i9hDniYS8lg1Qv0/7g+/JWC5xZX8OKN3PVrtISfILmZo
v5NA5f+ppnrnQBCgMTFSTDcoFXZ4HaeVSneW0k5KVkMBPFwbZ57lslKkJM8ZgCtA
69r02qDzRbzBQlyL0nDHF+BkrRGUspF1CGe+meyZqXRYgcZSOYVIIZhuW8duoLWI
j3kPnNq+1T7Au6g2NKguYpwBRNsD2g1fNFVVk+7NQzUqPUcklGSC1xr3Wgpov6WZ
M4AJo+wnKPI0jPVUqcZO94iowovZNOjfjpYKgk25bRZFx/PSiVVfUQFuqVxCK14O
Zt58K9mWkv1U+fjCK0R4HBMTXZcifHu4tFL0Zv5Q9VXzUyh7Ru1npaCLcQpF7A3O
aGn/gLWg4n0w0t5HMrCJp7HJxuvpPs4YDWlV0n3qaTPkW7jABfoR4IctCsnq+M5h
MAH450MQldjDT3d/k+ZveOIi07Q4MMVkinQqx39uDFq5MUkExjNKtr9Wj2DH9KuL
NWkMbWPz0KmADnoRevdKe+ZtQl9bBKOkEG9WRu3/G7Dj6TX4cOdrEl+M+TSNzh/4
oQsxw0t1hSod9d9JE+CF096RwmS+zd/UrVNL4U/HPqAURQ9ZD6vXtSbqhzT4CvSG
oCMHNb9lwlbh+JPrmIAnjPmKVLAJW07vpYolmDR4QVzQav52f/YB45HAFbmXv1bQ
Oq9b7dka/HMtmak/kRS027Y2nCaAGf1YOWNfGb92UvdqmUvOk/wWm8i8Kqt+1W4D
VixNSmuxXa45l3hbU+Sii3Vq8vPEKaENQe+L4YWTj2pAln0AUyzrF00wd2NXuztf
a79khOzq+ISjqdAn8y7S5ymBWLgbiCWZQe1cvlUfzuTeZMhfBozKia4ojsk9xAUR
D4Q0ZrFNWWbzzt1y7Y7m+swCX74oqy9rkH4nYc4DMt1OCVaaHlQHp7U/Oy3Q3Y8C
lohiTjfh6NJz0yR9CnW6eoIkrwfSBZplR4zLcR+l/FOQ229M1PrFicC/52zHHP9J
WXotjNucIzHZg40OmMpMHy965+7zglsC2Y9w3AHH2SVbFMUwkstFTi78lFjvn1+3
87AAX/fDbT3j5foB2EZYNL4bvr8fEy/NXCoEAf/+EBjKpkQaZBf4kYJCXcJfns7R
ozadohzqUKIgrH7mbcRR62t1MK8LGldIaugxAmaeZP0T7FGYpFFBADzoYFztCwJa
PQwMCLSQgzFRlSiLeifx3ivmtsINlTsyJEtHsdtw1bZFpqB1LdoRDyIBGVU8tmxs
BO12s7BG2FzBRxUavpu5eDrWPw7NeK2Kg4U2TYg5zZnCv/xVD1GQK5OWvlqs7JvC
jqiFgZGLFiqNaeTmlyDGfdhimeoYeE4aIHRCMVBVfVPNw8obRyK7iloqyzxOF2f8
+pSvZYGbQgC5lKsvzjc5lw6iwUB/ZmUG17nUUl5N1bXDESDwGr0dO4+SqaD7inHy
VFuI7JycpJ+Q0ccisM1c6Uj7/tsj4NTf1znlnbSuxnSwiCWXiAo7sIz6urMKpPSm
LAnryfBzxWsehgkRwMxmsBk5UxL9YFTs1B+EZDUNONYQG044p7ETuHAWfhINFYGr
NGLVhXqqSV5MEL3rSJpM0AT+LXu6L2vrrJWTFKfApnAZKJRmoGwdXIdAbZp7Eap3
x+347RJNWbwje/XotSwvGHE7nXl9yEqCybwpIVkTe4Yx/5LudQHH3u106BHGZaKi
f8Fn9lwmZY/oVuZhQEwYwlGl2eI38HyCOzv1jpK11qEP8sYoVYg/qBOmznn/LxCM
LHK2OFh9nOa09PwGavg84ALMn02et5lTdNWpCJmPae83Y78iZSGhMkStBoF4n0sE
iJ0N56TJ11ojBGCBwt6wLgumm0K0PNHbxU6G+OYtLg4IRG9brvlp4oWmO2WbpZdz
8KNJc6R10vHMkD65B5f+OQLTSKw23pY9UDORdccyLUJAyiG6D1FcW4IGAtKyv6Ab
us9L/nG0Ih9s5JJPDOz0EZSeqmP1d7IdZw2rbOE4ff6Dt7E4Bi6CN4pmWPp7EG25
PcmPslTF/HqaY9/yFhjydXy4VUD5ImNWdDQehedKT+V8q7R0IgZAils2ulTqDW0r
E3+D7gtgJtPEMfUSUc+g9sfEaVoGvn9YgCjFnp6hg258y9Af7EJvDas+NQSuQBlx
tDypwP1IlCGFu2WfG4VN81Jr3a6qbUGP9wNN9vxFOsrTDVEQLusRsc+E6XM+w1In
yZBySMe6L7oTbYSaPpVREHbDC6zYcS+LEnn46G5iGGSXLmOeWf7fJRHaiwHUZfgA
sMvq0cXp/4r+Y/DUsn1XOMtGUUicnemFiBcI1saJI03588VckccHYRpyEd4xhYI+
l4rj07n0sgCvtEmiPbG2HuM3KDSynja1iwzYvKha7DIzaHXl+lOEgjZ8NMC7i1qf
i2kT3Ubuxc9taCwYtG3ZXrPv5Uk/OgcJ8S2gPESLrVm9w+JognlEAP16/nCYhoXR
N8Cm2FreM8gNA6j5NapdAjl1zsn/WbM1mSjPnewYGUsTBYOxW5hCGjFwzkW7RmKE
zmMsmpKHHOzXh3/Eka/LetU05nU89BU25UB2agVnVQdGHOI81VnOCFJ7xZvmN4JF
2NBckrfE+henHsLikGdFKYC5B0eyanjitZ3oqBlQmui6IyfcYvFkTFij98qnnsS1
yNhWi8ZeAyIJ6jbXLb0ulq6GDQIsUHIvU6QnL3cbk6hHBuKnDs5fBr9eFVsi1xKw
dLdz9h31av8ZSESDsn/txV2CKPc8E+dJ82nLZr4lLoVZ8s3OE9UMyMVM//WelJrH
siyGp+x4uOhqXz84p+WMi7jMQAi0JShMQe/5FkT2p0V2ciucRUBufKpj2sj22883
j5g8/XKktQK1Tw+xRpUVVZc3qRu6RuN3E1n/z8JrBwknkfdE6KvbKbsQ3+7L/68p
62yJODala/aeU0hlgTiRZIhRfT2AR+KpFTegNN3hC2bpo91VEtjmJfbtBJRzaX+o
d3XTacw2xGS4GYz1DqW5vwyId+P39xydAyIZGT2IVPNlA7S8pI7e118CqbrW7LGV
jO+9lhwEE/TM6fFnfR7vYNmfHvX1mULMzmJKYjTIFO201hM7ilNqYEfxOFYJk7KT
3vnLdY9bb9RX0hrZC1sJQQVi/eII/R/Dxet8RCuRcubd9Le/sV0OC1r5L472P7zU
pEwA0CAAb5SVq59ZVl/zFJ9ybjDSpxAQuBDkwTmoByGbs4IssIj/GGW5MrBF3S8B
YkSgpsIfD/AXprOKVHri2Q25awATerqehSnDgNDXUs24vTZ3hDSH7NJ4pT2LbhWl
YQTVHSdtxnLaJ8/kipjqnuzmOTz7V/XdOFfCo/ZeNzWauDQ+iX+YTGOF+xTllJYJ
l1i8FqyItORbJLe6CxwHxuHIKDHuji5YKbd7mQMkJrkvjqcqy/Rm21lYsfz0Hhvw
PuRNfMGmTH8Q3mNI7AKC2BJQUz0IBR3LpsrFnwHAAwZ94bbSKYIrc/sWlJMeqiTq
qVsLr3dgJLmZkkaf8i5C0gUBvwWTmZRccagXvdSINNHhWPy+7gefn/s8MBMZ3PFB
BRTqPDVDIi+4w6As0q6M8BrjAtbk/fLUhx4NYme0dGzzAtgDjJ4PF690Xg517q1T
vTm80kjoJVz3zkF6allbjbnCzLf+5xqsoiUYASHyD+a8MG2yPuWYFEwKPUhi6aLT
WmHNXO1wDUGn6wEMITAppAWv0XRTGoxr6NDOBX7TVb6LYU4CRavDNofIbVrecLAE
ppRZYjoCogzCvoGG/wp35IUr4x4DhLqFY2ZG9q3mCGlEZIKs+2PSrn4dhXM4iyvj
csiCXV7N9rDnmOBP6Gp9lN6lW7zclvCaNYIv1CAACw/c0k91+wzRpBzJfoX+xIhI
/LFd6qNZYJc78soo8CtqvzixmWvNBYBF/TW5ZmqamlwRZLZ1V30RAnqoFjKO30JJ
GBIMHZzuzj9oF6smxiidb+m1IigdggnXwrhs93mkYX+owbfDobxksanz8Bx02lY9
MsgARVGKCgLonfUMQrI7uU4xATyzwFsPzvsBTPbk3Hb1mqhpRtRQgribEnr1mhWv
he0jswk5lsWri1fTWr44HnGbNJYtY+6oh5q4J3/DlWvd1UC23H2osn1TELuotWH8
UrN9gHWIVOuaM5s9EJay+lfHOJHOq9TvKS3OUj9SIsOhMLGdGjfNEnzkwUysFMeu
fJ/pWuKTzUwcMfPhBFhOWCt3kAQFQVTUhIyVi4muPjuAaAADgQVxfBXPJLJA4MH+
AVoCGVQZpNUuOs+agn7F2UGGr7voUwRyr3vdcfgKA5mLef95IVJckI9xkPQesQK0
O6+RZaGFAh4AR9yGUUh6L4esnpe+6UPjrtc+kjALzP77qkNDfXz9ua4/xbx1gZMU
lN+VRPLAeTeE6xe0DDgbi/e0TKvJRX+i+Swnat+/iuY+kXxhR5XLV2aKGuS038+2
OM2UQWMwMXVjQPL//BtH4TtHPHGQmeNXSTVE36c3ZJAUubcA2yXk20pzkIlREKqz
5cJ1zmyN343ElXHin/ioQF+WNug6HVNVuHoAfUh7U4f9D1AsLz+V49MCtzcksSnI
WeXpsAYBSov1veh3hv95cboUPVQpLeTGs6neJwS5a7QP8AuibWLywjN27A/c08MO
4DrYmAyvDxLC0npG6F3wRQvItBvGpmxrnUbnz6RDgAy8Nssh+y/5y8QGyJqJBShT
jbrwYCXHC4tMwZF7JuRU0RUifk5h+6DM9o87oCuhPT05uAlVJTx474U9reIP8sxM
wq8/NlV2Q9jb0i1gPeSvJdC0F4SwVi5aoI5hpNg4vTaKjeK5wCjCMC7tQ/SsycRI
KLT6kWsLywL+nlSLGqalqaHfT8TBaLQqIGeOwI3Cu4CYMy/SUynmSBzY2B9z2syd
fwwsD3TQpRWyLl4rlSjl9bUwSUOiaAjpgd4vghfyD9bwnXISt7X18umXysJTUSGS
TquMGd30AD2GuGckr7kJJeUPYdR6izuO8R72qQfyUenGZzecSQKlpBF47tEnzDwo
GNxd1VGteye6J+KKrNzvLmwInHR5WecFAtPwo92zpRVlADw9z+FdPzgVhlU/28Vc
MJi87c/A2PM/J/PEfElhP8fwLcKtRsqcRlM6aDOukJGLjQxs1q1uwYFcSNmNQO73
L3saO0n/4KEQAq/smvsxv33tJkYbsI2Jp3rrtUsv6iXBJflJ/ZVCErUbt7NAvtf0
67+QNWcXwRGTJ7weVRgvT8ygf+UKtLi0LNsb4HlyHvGGYPI7oi23wOB65ULDwXze
EkXsjn4bsNNnCPq4Swpxy2pyemv0pAysTdSpQREAJTUcEvlSOGPrMPE01q0I4Mvs
06kH2Yh3S8GWdAMt8Zuohkt0Rn6+Pvv3xPI/cDEC0k0EVFcEjQbSznrsYedaMYKe
zVYUBMbQu79PtfFx/Zc2Q6pUoIpGx0ZS7c/TxDS3mrM4yarpOT5aHJLN22HBMowx
fIOA91gvEEGnSqyCf23wpXuX0lLrgw08GSlzOC4uxu73KCXcmfrLF9iyGMcPWZ0t
7/8R8sFE+sW6Ff5gJblzi/UxC/jqv1098TEDY89bZXtV84yfspaO0GvZRd2RFXOc
t2zN5fuhNQY7LaNkZTaLhQefcXmDY6es7YUcGOo0HLSi7EIAknmHbzS+FTb1lz/z
MPa55efNavKvk1LTD+bdDsTzVdCpq/nYHA9H8lvr8Nav5zEL0nuylNvi8P38M/WN
4GtnwJw3clwiLK1DfLx0FDFh9VLXD6G6vriyR2ba17dZet05k3iWLe4nrJepT2dJ
lZ5jfPPoBLvU4DNUjHsNm6Io9lop3pEQoyIWBS3/fO9ntyxfcJim2nD1xeMbCRJu
sQiJR4aUdFOdxWqifSIRvjPekkJ6hSu2NRsCX7mSlfTM25+kfH5R3ZKcRl16I9KK
nvSxdSNN9kOKHvIqYSNbcnc6eIB9HkSvRr/8ZU/IJ4wuNbKivDtSnF5k5y+0v7JG
JU7O7kQlUitF3DO9C9fHhzXeVi92GsfBqAccFeCW8Az/3VdVr0Pk75pvSlXLbV7f
UTUUAPbRFfii/RM/IvAZtXHB+YqMAWSB9cmNEu1QoH9CJgc64fnjYbHQMrrTbSNp
XHXJmhDjmooSTOIKblIvu7+XmHGT+gx1Ov9zjS2pKdgFDLf12tBQ58yDzQCkXQiy
XpTl9rVBBZBqz9TMRMAOEAoqmB44jg1TatV24EqGBpHW3SM3DpKrUYi2d1LI90CD
toF4/AbxrYGbrhdVCSSjWsMWNMTXrWhRozo6gDFvfoMGeRbucfhp6vexiSsAOTEd
y/UX1HQInkYJs5786+SPm30kFq9pTczAsDel66ih1ja/C7OiGnRsHnisD9/nBjoE
S525wZ+9VwqIB+jd7P1+Lp1Nnjif2wxAYOqd52+bsZyGVqevXQB9yx13m2r/4QvY
FtCvrhwjxQGdFHySApaHrlFkhfBGBjBQN2NSXIw2mwNjpa2llkLvEVXM+bvdkqsz
GdCDESm9bHKwCe/7POrSu3CqdLRYYEI7Vh2lL5paNPcEeU2skMyjyiwBNSBskvM8
9m7vAkaW3cIhFsOIXHV1LLsNWMXQgTRpLDrNbpALsx1Fgy/lhl8ecA8OiMR2MHzC
ruDbNrTKpDxQahhrhfsbnxzDd1goDHSZcyE6q7lEkCC1n43KW/w6S3TKetUFqjV4
WLFM6ZeXzZ1vMm4AfJC+ZDiEi0c1qPJ8jNJ1jMgaGppvVcxR9MxgiTXZ+xoV1MAf
8sfW/3fTD22mpXGcBrtu49QGkza/A8/6JOTxdl8k7bTVycIaFy5up6uFlNfEeUZl
0BKRJ65EQ3lnU3zKeyX/0WQhA+GxUV9HtmOiDPochMVtachmC/vKgBDX0YIzbOME
eXHSHY8O0jIoUs7rW7C2z+7XbMDEhpKS4e7Wt+kB82j2quMXEC7DB/WXMqnmAM8B
CcRxtOqg6ZAKh+5tClC7I6Njv6wF3l7CQ9S8CtE8BbIAwRZxICWDGdS/+dBujWEL
s01BhpcQP5ynJDxyurnlRg==
`pragma protect end_protected
