// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:35:26 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
lBJRIceim7um7CETr4kHtsD2YnMtefMEhdAVAvFqiNaCnztf0d3GaMwG0OGmD8Q7
bJ714Kv0FyzwD0tvXGL4DHcARerd5+QQOzHv25rO8JJqqvpA/LF/7TSLGhDoIABO
AAPmJQl8jYMiyXrZKntGf7tznaPTuTuALqcTiA19aeA=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 6736)
bIkOrzDqCkJ1d1JuB86oR/kVinB647Wv5hOlSgRDBE1wybdc+9ll5hPg10UpM2z+
8XQtpzkXYkKCrtA/DvM/FINK/omDDcGoGqEiV1gb62lI5++AE60C8A1Vh1RuRKAg
r6x1eu887VjxBha/+GzHBOFmm/GieEamdcUGNmdMCwuiDEJ/cE+oOFq/2FsLTTiN
GaRmV7M2LWbjbMqpe8GDQvQB6PGhljo49MgCmXmEjvBJRBcmdf1RcHYISamUNrbv
tRu6KJfGkp1E2H2SLBGzF+elRSqGoALkO+w3XQia+ySSo8ZFjvDcd6UZI8d5A9Rd
LbQonon0fzQ/eoYld0OAYpUIT/onILPBQAKXZGWFFhp+INUkfVF/Kg1ujHGZJ5hp
YZUhl2N2AO/649zX7y/NPuBtPzITrxkp1dLOrdX1Sx6Apzfg2nINAgCesx8xK7og
AjgHhwr0cdMY6lDsIs+2rYQlH8oB+YtItZoQp567c3IonFL03TeltIy6nn3LWmCI
+xC8JPpPU/ssikaUveFrHDqzqgx8C5N/ZG+FrBum4RrClYNjpX22sGkQlqKSw16k
V7GF7l62oQXOhKnJG6lLOz3NNhnAQnnx1Q6sGZABjqDDYZ4nR3J7V53iKhegXjWp
6dqaxZkPEy4CUqG5gU/CBrs7v/d0A1HhaJrAprXsedNIVklqJMEWwM8+LYyyHGTf
nqIWSV235NUIqWXAiRs5Q7vmEEifg93ktM7tA6n0Z6hiJJTXTwXGjd+nw+mYnc0d
oLfdD3DEg0kIMzRTgkvoCx90K7IHBwZMPSE8BhYSeTYyyWnSu7gve0iK+Ewd5Sni
PbQwK+DN5UXO/YR+g3iBNyKIMICStBIUYnqAIShpmQFBdbo74hs/jFzZvV0O4/hx
98k8MAIG9Rmw2yJCmTSvHQHN4Md+I49OKHIhZFFYva7GHgYvHiVDGnKVyxsoZjoe
X5oS7SdIW3qjJA0De3THb4AUwnUtxu/UKNIdIMkETLwo+rf1jpFWotRV7xRLf6m5
nqCyJ67Id58/QcEhIlEcqhzVMQVZphzwW77VY+uto5565tunICHqzu+wcmfO4rc5
mpAefSaXDzMDf9z2pCF1kFo66f84WG49mepDA8tRppOk0lrg65FN4/gh6CQJC9yw
yzEEZ3ZytOiI7WbE5HDWvgPb02t/y4ymxdFF6nYG9eiopq7AdbQ7CHYsoFZOcCRr
jUVw/83zuBk4Z7zbk7cfFJIIpj7o9o5tyShbF8aI3ToFzdg8npjbItXdVoBjI/jP
9Z+wEWjQ4Lk4zV9CruOymgeWRTQ/dLy9CqCI0k5YieeVNkSDYE6p0TNgRF33FspL
IQzBunjsv36tRr83G0Gq8OE/9C1CJMls9PvkCzkNNypPjdCVLixBpswUmak2HSaO
MXa1EhBHydfOcR1ZDObblvEYuC4KlEVy1K4r0NWZM4Y/l272pVXvzV3GOTYaz9uF
0mTQIzuprX5FYzdNA45VOkPHp8WteosBGnbQl2LY97d2iMrLfsOsIJUSofwexmv3
gzu7YrbSkzWhTGtwcoBSKJDmx9Ql/8Kp2eZxc6CxRy4atSXArvR1OXaxeFsFsyQG
TDreB0HHtEMVszXEzR4G+bE6PxwVi/goCqvWXQ7usX55/CP4ko9VlFuUlacM+SD0
IAZQJnxs+Rxs1yQvfGmUamcwbZPBbJbN+fQHF+qAa4VCuDOOLm9oldrt+rH4EXzE
gbNsXK+vilQbWBslv24bNhbK1+iHF86hriWsABySWQc3rTtCGDT0x1/L9YtrJ4M+
Ps6MnKJqPbIOiVeQY0EulwCEfeNPVqnAYWDxf+80gRmpRTvTUJZ+PlrBvCZ9jJNU
pK6t5A3ub5Kk/puwncf2YSNJ96N8KSPOJRTIa0UlK+bRjt1o6Dmq0W+0nyBG0JIM
ytlAsoSW4vJ9/+cxg2RB/D1ZPPwNpKA4h4NrpDY5fjYWW8nQjNbL6Irlv5rGPos3
TmLfBLvvN6w76nizgj4VSciH3me4cY/ySPxtM7iiuI8RkcSxJVyPEiU/+Qg6JjHR
rl+lwNrZZErcvstxgx8vIf5aryn6/qqj8G7A4/xXpsIwTV8kn+epCLQ6oMckvrJa
jC4h2uLooLmnWOJ8Br/xYubH0lEI9mAYbZMX30/bkaIW2kK5Q4WdhATHevgud4OQ
uA7etT7ZL3z8D5+TAqogmMnVXaQxgfzD07DSU2EuCTCaAoGPgvsCcpLVcrWcZfV/
jNRPswTH5wiVuhifnRi+xap3zvoe38F93JD4NdpKv0yspLeYD8Y9syWx5/oqASWK
QVWBpj9WDhxzBsuyQ6Zb1xDAv+aYdzR3l9ORLFrzl9KsXqJWvC08QhnppN0k7sbL
95nVDOElUQAiF5wmGamKpoxjrepdeMQ5O7sTbwa1OcAiKHoj0Zp7ZctvFR/eCvBA
B9WIuTSBpzEdIWA9PGC75MD1+Es/seL3YTPBU2vdiKbujBDwtDfnXA17km1uspr5
6+S2jfUrWlFxi42Nf0CRKT78CVV0CHyOUS8Y4Z/FtEtgar9SfFhOaCFNTgvb6BmT
vupsuq4fqqhnBjHILXmJJNHt/1HnYVi0ttQDnbJER/FkPMrBcqPqkTTNLuJuN0KJ
cyKZIHOVhMABzk/AnJfd3StEXMq1/v35K/8E9+H+QU2hs0wDZAV2Kz/rbYkj7JSe
vHlveu1rnLzzrdGC7XmT+P1ghAy4hLWCgbOa2tcur2N95QYuz/JVn4Jc+QMtto1u
mT5+uGL5zCuz6ekzm4Om0msbP3yr6CkLhdX7guN062U/5J/ILjLfFA/uYw0NnHNB
XvqFC9NZMoIL9vfamegy4P+augb4kPr1he8TDCcO6brpCnKXqcNKEZ/5hRlIV/fk
49kgmCs7wJIHAF/nzwufz7t+e4yw4EITIaubhAp3kiRD30LBfeHNSuWWBGQn2DxS
yKqELJOti45IH37+9NhqbxbRRAxV34KDN9dOmcdm6psn0DLTh2mKX5g7eRQYYyNT
x8vUlbFG7hpdn2Tjs3zrTYtO8qBKBnAMvQuS/OEnMSfFDEYOQLJYAaysp+NWzC/+
auPNRExDbIFMCNY6mTDspvEtOVfoy5S84TIIE1TucHWaYl14ObyI8MzJXWEsnGY6
8JdocwVUEBljCJAFjobUDWMVny0hYm1Q6xKOBmNXjDiDAS+TbuJv8bbBeORAIDwk
E6Ne2seZJklEuAlkpAAnK8/kVazllVHJE6qWRkWmliTckpPqLFTMdAALMes/O4HB
cfpNjLbuehSmPnjjVlOPUHW+ZL/+OESyWvp8i57wUKIa9bJxAFW9vNu+i6VDYKA4
9hxJkj3ezxKFBCzNW1zmUerCapUkI2+uKyQKdmGemlYPE3E3AmqrBbT/SEPKegO+
sNVEw8Wmgw4FA/W2WxZuIjXqeiYB8UcGHWmYBjKHaa5gwXkpumzdv1dxR5t5YTMp
SFAk6b1vPgop0YQweYOKEudeULeUzF4osrkPafyuPmKnufmjQxUEYGFhvb/benPN
qWc/A4MluhLx5G0vgWAHmqhkHDZrWBtCsOuFMiBoZgL5K0+CBZUNLjCvJ4NodD4u
c37YQEyF3zMbHAiDFet5o1fmiDKD0wmX1B/vqnVLk3RMIH5gLYrbziY3Hz2SLKuR
qs544kjbBit6pb8e+QHyR6AW3tdgE35vW0WjjgBMovVGxVlUv9fcy4bbFB0ez5m/
3pQqWpznptQ9In2gbXydWhcAd0ki2l1BmGoC8KkkSBnheUl8XhTpKViLFGk5Ik3V
umVi9ZNaZ8nNNEivQb79+BcRTeCZCde20UmpPj5NSecOzfnVCmBdftullJev5pQg
/BzO4Vhoo+9fJOcT9U9aBghcHLgABUfxnzNxG5siuQXy4vFlvQ6ypBKYQ3nigaNT
QlbIJQ3dH3WLw7U29oI1yhCsbWjx58BsW/0UIjELz5U3liWcdc4baH6SCxi2Ls8v
ivmQuiEWHDd22WjRuAKYrLe81ZAHDqlHe+1RU51dypV0Tkc6CwN7m52nAmoLspN6
23/MX3TSR5RtI+49gyJBQiQ9C/QfSs6w4sBIhz+XaRmeF3DgolOKG7W16lW/lQ3u
YRIfw4MuX972rz0OEPYrQXGcNAAdXblvtwmhnZmuQkRuaPUrlQTW6usrb6pEZiLy
EWYiewx6aGdmYGFY9x1ASp4geIeq2wiMsFhuLpTvPJQul5yn8MjlVy/DFUwb+Ssw
Y0iLRKQ0BFZx9ynmxbmXJzByjo23AlPeTd5ywJA0BZk/SzjeG6O/PMjS986k69eL
kNPg2aYCIA8fWAhGAp1UsLZ73NhWFvImtsxUBnknBP35ZCn2IaciR3IrfnMkZ5VJ
Sk+XXVWgAH067jvt2MLM3MUodX0TeEFNjh1aZ7pBxRU/rK8OIiyyvMjraIXloEUA
1JYQ4U1RqQvIpdailpZV78WhBddTx+sTrPFpFTTQWrCY0QFx2eIAFYn34UDbYDRZ
/d68RYIJGzZGvTYNHCNJH8sZksF66elhLCAMQEVo/BRDcLavMbq+u3Qwmlgo3r1l
ou51yuyKqDYc6PdYjQ85MZksqpA+tuwqvWQXYKG9EwFWnoSeYNIWOOGcQS9NPe9h
l41DO0QnNUyopv0s9Ydy+dzmh+WyoCdlwBAR+zZgcyxR5qk19mhqtj8Zp1OKp74d
Gkwc42mEorr4R67cq+Pl6tdE0y9PR+fCIw3aR4EhqKphW8p+FB++kUtCs6gakOmI
66dN97gurdRp+BhPsRuzyNZ1VCuU8L029Qo+2mqM8gXloHd8hIvsBtAdh9a2PJGD
2JPuv2O2UlaSsyD2j9Dxq4xVqCkp3I0DpNRo+4qDp1bxlh1GiwNp14sG+0NeWHgj
XbERnxpOxXIR1KQrZSPBHIHeSTp8JScP330WD0p3u5/kFvKHR7aFizuP+nipj6nv
6kTFq0bHqtXQ7U6OLzwWgtVDuuPhUiGvoie03oV2Bdd8zaQh/ku+nFxt8OR5T1om
iCRbI+d4NxeFhFTY2uMFCWpm2HVM8q2SedyTX2qvHSMc/A63JaVLs9bBTsvHhcBk
np9e5m/4eGl0FCUqgyytbv3oO2jXlkoeggoKAmCv4aAaG6cytUD0gCcC5voFHOet
rtKLujbqNvQ0CleYQQkHrtse2VOX1gsrgOgFNv6K8A45N693U+15nx2ZQ4t7LEBq
B0dfdjAHuW4z3nbFnKy8mTsgulpW7jwbylRHtJ1Wf3ZrmG3Xxxb5eeHlN28syBeS
godxtvbI5gh1JEv8Ne9+fKptKnVtGTBYwKxakECK8+2l0DxhkXEh/JGtu4wdxzo5
WaU4t1niR6R8xTSOhiDYt9deacC90Sxz4ngqzdn6oRS0+HqYKftOSSaf/FjffAwN
KlfnabxU3Et3+zLgty4rJDU2ic1nawUe70d14LOTBdFjeMkhTa5sG63IxW+PjkFC
nINkdhBBBjLvpSXj3lDp7qrIJKk8s2UjUKRZ7uKuUyjSSq8bcNjTgEeTf/efESVn
Nd6HdNdFm05ueG6Y9ZTLEpamD5jEv+mNYUjtVNcahlQOuzU5qLjTueA9SmgOahw6
OMO0mQS866yQGhlnmtFXvT0L6XBuHr/0/hugtOEpTiJGBz9ZWm6/pkGNd742+o/H
iqmknObxBCYXNy+dMjaOJcnb8N315gYItNLWPppJVWAm/r7ICM5FcvTDh8XqJu/7
gzH/baIZaOW87/ZpwQkZhyioNSBS1mVZRTOxxS7bv9HksQFr7vhWZSe8EPFAKeqk
gHY9e8mYDxVXk3mD7nHj6Ia4bdgaLE0c1MWXL4kdwT9IaaOyE7beNtu8kURWoJcU
L4xD/zvQCJPADQFlDmMINFDp0CjcDY39ytRF3TU7n3D10jk+UY48qlNnvLB999Bb
hV3+ye2hyBpF9/F5FlAq3CDj704UspRoACG27sik1jd7KB2OA3n30DwhrWTdWdSp
Iq2gKHCNYPWB7FevCos0sEibpRa65SxlKm6mBiTzgE5oAH3PjPF4EEy5TchfDDdF
Ek8Gqn0ZAVTMSxUHyBPw7jyFFFBYs3mcKSjwPwg4YV435e0TN0HQeeBDiU/DUlEz
q/lfXEuAOCj32deqLGRnAtPOs2RThBuq12WeneNUzwxFeqIaaDGX3GdfciEFzkHx
DIjfrlVqJLW+UZn/SgpcJBYTy8Hey/VP7mgFNo8ZLFoe9wXkVZ4s9FE4Rhkq/Hj4
Bp6wBrA6umuwyojxGgeSXEfWnYRJ45R3HBGiOKQoZv8kCx8wCrfIbI7PIa25YMP6
KjHOpQHX3JMt04W55smN9nlP1va8Iwcx1MzUprlwzbU7vxekqtmQjzt27w5tfZGQ
lTjlMG+QezqUmYHRmY/sECbHp6hDmxIOB3WUi0qdScFTgzmMFGQP0KW4mwlm/2BC
/QHevklNl30UjE4VAM5nuf4JMa2Hib2Yq0rzVdxXgusqU/uXijw9VcGwiSa+7i72
TBZN0Dmp5LCN7kgTt8djiJZ0gjCvgDxs4Zq5VoJC8RCFbqkt6xkcrQ1LmyQXykDl
jY5RWMEdN1j9/h98GBGyvOS3rPn+/knuFjMhTfcgicnlbi1pEf4nTf9zpjQROo2t
a75jynwheZuV/6mPXNtMBIp7ZDrF3pX43D3Uzn5eY2nH3ox/7FOIShHmL6r63kIW
0XzmEMJxMlHyhm3H1P5irgW05ROFyLva35KknKZVWUFAte4dgtcrsNgWpKXa2J60
0I9lgqEblLIHjILY8aji8PvwrZYJ6k8QJL8xQISDnXjKkd3vDFPL9WWMhIoQyoL+
bI37hrf8gNY30z7eWzI/1uHAmTYMPoSy4xnkvAQ7BqHAgaeoz5BRAde3SKS3qTyB
UqHrcpx08XcG4OBxwX1CBLMkB8EtIGQ7mti6QH7y0aTJxrJ9JnZSunDLzMoArRAF
t2x5YKixN5A8AOO6QJrQT3G1QULXf5jORGmvIog30coPDe/RtKTy0gFPADCiG+rD
rbKAWBvGtd/Z//shWb6XTqAFOKFEtJ/W52PmJxHtXthHe917qt4xZfKwIKgF4KTK
WJSUnfTmj1YM/HNiAxZyIPh3pG0iUK3hm7LEwkFnvtMEZ11QkLu/jpwCYT/jeNCK
T0NtH/6wg1V1MKpxdplj0NyuOAgKu9360vGcQfDHFr9M8QUqFilr+LsurFDxRVt0
gbuPmwM7ecBVR4Nugw2NsLRwtIt5FlNFwVoCMcxS7y+TWw4MYLAHM3IO8+qqoDci
BwhPNan/8s/bx8fUzKqktyR8oBJnGZVcyNTYQZ5NF/uMg8h0E/e3yKFUs0RHJaOg
JepusQjZ15ezjNBUyOpVxtlF9yInqC1xAytNSsf99twOBHHkSXRqWQ4+/iixN1qN
O74BVVIkIoxpV6vbBFjdFnpI/OwpTVtnT5ptqG68ljIuWJ7EZCjpk64/Gamv0tda
k7/Y4sEHm+LADiCRWvBUkT+e/9wI8YsYCiZBE3gqSulhveSkJ8NZMNlMsgqqaIVq
6aP1mad3kKyRMPrBEwOOMSqBUMzLSbpYCTrJ2/VSkAY8px9Fn3PAE9YGeGVJ4SiT
ESRz2zNESi+RQB4TLap+2izltVtjAVV04tDMGkwqydDQjszurS0K0Y15ftBmttth
IEk+NdjuihEyc8arQHLIVRTHonBZ4p3lIuoXqAT3OvOMv87wMxF1PVSmwbIjRpyi
X6NsJR64FxQFXmUx5pItQpSXPYRz4u+0QhmK4bEDLrFneGbxJXdHj6eLWQIFuabG
PKOivFv/lhgBICz5R0X91uvKjOewT7s9QUSW1MIpvbmRSXTZD81GveF3r6prcOup
g5UbLQN/f1BH7uE8CnDevzlv8wziJUg1WoCcVRVmOT7PPlhqpBZPoSsP+SuOmrEI
CLhuNqWuIGbtD9fUrb8/wQD8FduADwtCa45n2EGaioxqtiEJNEmoKwyOaX9AYuYt
7zUKCgxbyZUH+jB+yxVUjTTyktbW/CpjQ6mYP4U8ZkZtvmOUF//Tra4qEoauQ+iV
5SDyweqnMSuli2Bix879YinNdk8isa2MmlreZ5eBhKCN5oD92VlClE+MEReLhQlI
BYbZ8URQmMT1DEy1qUnsuPujArlDL7CyW/GaKqY8wuNZBRtcdcko1TYAoFHC/Va9
UdLWbnNJ2VOvzu59GbkiUesAOcDzx3m2QJLc3mmtJOIJ+Ek7sKaJxDN5NAhJMEeG
eP+17AIRKsGLQSxFhAendbfQWbDwmUmYfC7jNAC3bzVV+h9UT4s2RCFNdSTD2aVs
WiYTKhfKF0KflTdtRNhyaVFb/LB0S0XsbUZsOfU2gQDMT6Lvl9HIpN5IwCnJbWUs
00z/o7QVZDaUpkggN3fxT3D+QF7me12KFHUY4Id7MllP405gSgxYqqn3F+RF4f0e
IAGtBAp89g/eYJNppeusn7R2Fh5EnZuxC0R0pUFL9seQ2mbPtzOi3k1zcFtHyDDk
SWPZAqm42FzBL71jZ5msh3FJmbBgILXBBGsoPu1HSQz/yuj3/8EYicwwTn/F4TKK
sJRpadl2moEDoqKBw41tK5SXK7A1Cj/9Exiq58Yg35Vbibmwo31sQ6pp2qn4/r4L
1st8WUAceOWbnQDPTvvC6XgH8wstEH1Rga0ws1QnfsNY+9k/ACfIqRANsXN3FsPR
wxFSbSXFQNPi6fJQvCd/9oyHFwBxnaoaJ6I5YR/Nh85FCv22JHX7m78qGqCvoqBX
8nr74MF7CmxnI0Cgww7S+EfHye0wTjYa+McqDMs7HfJglxMy7C4CdOPL+l6iv/PW
GTyurrDtMtLo25ZgGOX8ybfb08MVYOXPnbwnpHPxUg9FCKs+aQWm7/dmJn30qpdE
gY1HU2UsklGIYJkmw+J2OoXFSF+K/kCwHndm8cRD+YMqME0o5GxQhfqjVLSQAGlO
Gil8PKvoaGTnmqWHoUaMLyfVDbn+z2WRzahZWKZu8huWQQFLa/E5kS3zu/FGe9gl
TH7jYwWRobZzJmPhpNSKdw==
`pragma protect end_protected
