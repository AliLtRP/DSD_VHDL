// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:56 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
A3dLTVbB7nG8EsSJD5OQMXf5N5kQ0sTmuuAAGqolIT3A5k/JZAc7lLxNcoFQmbaN
ohgEASpWkB+SYJXpBH+qYbYSprXXgMWAq68Tdt1czc9A+ohQHHACTK06pEbbWw5i
bRf118YAlzs+U3ib7XJdJ91PblShQfmNAqvwMu5PlVk=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 12912)
MEBQxS7WcoGlVIMchZ0PBNiwYmYjxHqOP0NTu1m103udzu/tSJWsBAnVRm3yaFJa
WChIqxByj+79fnXKapz9E1vm/25maWxeGGney8CstdoQduToy+95ge1NY6/UTSGu
3+NTLL3u1uqxDFoMPwr8VWSSCNQJWfnyNiHMZ0aPesuur465y4AfQHWVSocqVYw2
+ttNlAeZQ33LJiBjqdH01lcYIKtB5wSerg6k5hQ6HihT3j3LYSOHAxiVTpQ/ee6V
6ZCsy9slvnudnhRh1RERNFpX/HKGVmlAL9Oc2lX3auHH5z2UQItVqTeSnlP/AJlS
ukYXYZ6Dkw608MfmPVCZBdTDIE0sV92rDYCS/Xf/QDx3MbYT4vkJ35J17Db6xoTS
0X0TRSktGcv+uz7j+aIFyuh/4FVGMSFxjm5E1mWKwGr6mvZ/X8h+9ySH9mPyDYhK
rpIKD7QP6TFWy/JDsCRnYRVLGTNuEFfPulN8BfW5yA/yjzznrLvMdtyaFFPZZqy9
r2zwhkeYkoFRfkIicJMUYitNGA+FD/v6BY3qfXYQcaMmacsqrchFDj1ORmOrEsEl
gLqXGU0yJ8nM/IfqJurdyUC4q01H9uNebipXhzNJf5FesjJpBVdJEDYPnAojCEMX
skjRqlX7sreLQ7gTW3pxuzT79vZEu6QHde98L5gZFGUeu6Ptb7q8PYpby+iCAxvb
ly+/TyCu1t1n/VfVO88NOzysblM4dm8VhuR713ebOKmLCwBG33AfpNVklbFfDmB/
akAfmTbwwa660m81OpB4dmUdo2lnQPj//A2SW8Yml0jlS0g7cVgxHUXHNjICM0Of
sAqjgjjy4sjQJ7/WTf23C/1n9oMyeLcUQP3vYlgUO46+c1BtlpnKW0vabi2r5ip8
pM0WSMWt9lscesMxDObEUQQqWi8pRLC8WRHmOZI2F+MUGjVARMweGqKNsOzdzrwW
611b4Zyq4bAV9duXNe9qgZDPuizWzXQ679+9xFyToAigZHtFqW8UqhFoqWQ4kSQs
wDzE/RNBZyqfQpqRq05nP2Paesiz/VOYFih7IWId9YiS2gGkzA1taUB1huNTp6pY
XY0hKmvor/A1QbW38aJZDSkkdAMXCtLc2mOYcH055UomQBKDPpZmUWgaWv8l0jLa
OeVcJQVp0rHsPsd/fR3Mf1E2pcoZFDdS86LmNh04NVfQum6J9Zz81znQETH6zIP6
eWR9D20CqJm22Voa3cmMPEvZXSYv1x/vXHqaRyrV3taf+Y+rAXVUVA0pqgvUkuK/
Mc0QgvAPihADKa6pqda99wWghnbghFJn+ynserVVOHBMYuVRGD9rm5F3kksQL5HC
oZmx9hp5uwlKTopcygxjqdDEV/HgLtNeogbpfEQu2n5cPU6QSQZPM9lJC6pp/PNI
/oPLkO1oJoOpW2IkvTChOxxvC+AeIDKiB1jivZzulWZf2HuBz8PHmAdkdaPhKdRV
RiD1D67QNwruWKNjudLZoJR80oMTAKqOxCvk2rp3Xa6/uo5Vr7yxjqki5XSkelW3
LZxnT2RfKwGzJJ7c+FhMPI0Axl42QBwcXRunlMI9sRsMP6xkMR920PtFYw1SWesM
QVy64uUNikfDmB2DAOMthYuM6UGhY+S47hniO20h21xCqpk5BcuQW1G6ZFQ/3v9V
0TAMYnSjqJQz4go4okfBDGYD5VY4J/v7Xp++wMvmtVxlZ/IFlIsmm/35JxBbtHOG
83MbLKvokkWF0Jph03vTNCV6TVMJ34iqPySxGlDHsvGvtrxqY1TcNj/mtwNEopmb
auGQeF9mVQUzZv8TZa8TcHsPX248VaQA8mcw5Qu1lQMfXQk7YTbRjECt1Su/xyVr
FMD3/Z/a/8Ml4AdrZUg1H1A1KtFQVmCpl8ncoNVgtn6eyvPToOGJ6Qg5Gd9E8xld
BRe0n4j42ZAE4GVmG/ymrUoRgcNWMi/OdoTanbWYi3OklFMlcQaytg2Av4GC18a4
OUVxfhj0h9wgq6/ifolmHNAuarNg8Elz1Lo5JvKTNNYK2Z9A7yqTY6Re4sANFZrK
fyw4klzie6/oVS9zNdXvZ8r4Fxy63X/Bi7xG67//W73YbP6OyNhyVz6Ti976Nuq4
a86/dUfVx+0KdTnuOhPwCTifmp9cp/2603U9zKUns4GIt8cHgr1C20qloIdyg+D+
V6jOZhudlEvrIwHjqKB6Ef/tXgFcS9u6u5P6cEF/sFjuHVTOPRVGfiFVEi9q5ata
7QqL63n4a5Dl91VFmfSRR9cHjqGrrnalaUaCBCDT85IZepdMN14bCO5/fIlhfAsu
F3WN9Kx328jCiklLLjUoeRVsQgBsj5OkD5IUbp61roI0RbnZwaNUjvWf5dnjAoCk
yrOKn44208E8szHtpPDIiSA3T1gleOJfLNwtHoUlA1dRyiGrZps3PTHswnx8z0Eh
7yU1M6fgMimJ8nYFtj7zHbvVgrTmARt15M/mJZYtFxXszi9rYxatEbFEWw4SGKTN
3aPTop2xdL2IIP1wY75U1tKnWJreTM7ceGt1kSMQx2nyTbwn9/YI2I9KcNX9FVZq
abk/IEhMgIX5bZihhGkBl2lYkzYQ3bfgdj42HP3/SY61g5fIOjOjBEf1at5VF19X
KUMmReR8bf+gzT5VLoe0OY+RnEkbMovKgQhjsXV8RrAHeHkFacII2kVuCWkWndUM
muNwoEV3Y06QMqNbqgu6wqvzw+cLRqrVANhocyVOLr6Z35136uNxrp36ezv8N+NR
6fyP4knF3UvAAgB0j3DF+zKmHBG279LMCdU0RkQY8UpZGtnWVi3IaSo37QFRZ1sV
q+f2Px/9Tl4zfa1jmlbafuDOXNBTEIk5SOuY4EXsXLapxQpeVq60LgcyEXQFR9vr
ka0qs3H+t29Tkt5LcO0cwAl5sdMeBCWG2629mIOX5xy31l78InAI1v8lrdNVFMfu
dgKuvhbKht9AHru5m5Ps5MmxYDNnLqdWfSdKz1ImfSSMuniHNba+mX1WXJJMKzOO
dEE7WHOV72/wAWY63j0eq88dcxF1JHWX/prdbwCdzJY4v7QZIQCvCKgkd8S8yxI5
N5ZS+AsnvQgpJuFU3JlDHhYAat1zbV5YRtFUX5av8UHB4yswq8UG1Nki+ljee3m8
0YCNJ+Q9K6pf38MZ0bozR7i4H92KB3GzDW7XsmYQQV6N6hHd3BhHgaaQvkwcNjYz
fIf79J8PekiN4jSWa4yz01BPVBmRE+rICK4fVxfWiI9pCeXHgQ1pumG8RZDzMzK7
I8yLdk8/4mEILD/62nr1VGdDhdWWt0YpL2TyikSpuBKF1ua6Aa0dnX5zne1Hk32F
UZ5fzLquxG9RDOhe/d8qQIL69xlhzANg2LGtyjLp8VHcEKaRpJGN9ovSxlHGg2iL
TS5wqebBjQnvMEWw6BSaVi26dt7ektdU0SsyNEBRvxt6ciUxav61rQznJLNrSteW
pRfj5yisAjy8KDlJ/yV+jIeB2SMK6gddH693kbz8jqWwZ10eLq5rUObyxzvqHAXP
+vNwyXEnyQ3WmWLSec/m42TzIW+WTBCdd/sJSFZ4+l4H0hVNZoqGir3PsCcDQQ0h
sTWnBXZV/Vj9FBm8nPyrD5jh5tfM1WRtYZwyBIdTtcYiQ8cnlr4MZASXdpJ6G2wi
EPKwyPNJ76GyfaFxw1QYohBkI5TcYuRQGJW40cWPWCcmlKBxaP1ssaTykaf5Kqmw
xuyogOA2SzVAw5b45LLLBux4y4cIIegkhe7hEeK6U6xBr2hN6p0lICcGe1y5lzyP
cLcfxeaNJ8VmeLDqK4go4B1ViG6klGAZ1N1lLY+lN21GnR6jLPnhEThi1x8vN8Jt
nRJWt8xgAkMf85SlWtS4vIqS7aTwTrBbpdBVPqMij/ysaEurnOJ7zdTIVV9OjFff
9gkkaY9BqaiSPfgVsHZm3fLlsUkMTC5zREsqX0/DKgxH4tkAJBTumuzIxqRPAQJt
bQItXBwVyOew4L498rBaT1VVyN2nJQwO/iKG4JdEHs3maALJwlRNPQf6mpcNMY09
j+AvoX9C28ah/7xtl2Dc6J/a6czT7/QK5qvU1tIqcW4Mf7Ug4dGuJ5Pc+Wbc7RF1
H776uyUCj5HFExisc3inKihSBqPU6q23RmGgMPDz9ZF0BNElQNsUy6loJTVn/Rd0
kybYnZm1DddC++T5ksEBT1AcAiUxTDvyJmqn7zgTtFkJLjrm3Z2cjVA+gNzdAwNa
sYvWXSRry5RIuM2VvSig6db6MR07/xl9AqqLXF+UhabW9VHrF2oRLfAa8tleaS7t
wDOT3p3z3HY6AHeE/YcLe1UNTFekhbBA8gLdyHEqaweTham8e3xn1Jo8NFsIrZcW
gYCNmmv5CcGRcva52dtPHUdWaOrb146uRyPFT736cK4Nq921Z727GGPFKn9a2fPd
e2M2fA10/0HcnzCOGzyZ9wXhxhm6hE3KAtBhEN3eTQ8rkbc8gcX/STfl0LPtDzbK
bqlpuZ2YJ7Cv2o2SORckxIdL2b4garfBMRn9EYAPRWMyi+8b/1VI6nWoy23ZcVpK
TEL8RsTV2s0zBUNRgVmvasYQnYQZaH3WLtyg4Q85MvyXtaOF3rWO0sKn5zdJQi61
Q8lxD7aP1/wGQ7d0bQZUXVxolslchk7dNxz5nrt+tL5Y07Zk0otVnoU3PyeLtlDc
I4w5vzdhTKgtpEkS8mD6ZKeysKrrrjhKaLc8+N2W3n5B4Ega1nurpjSedZRwOaM1
XFktI3x0F4ws3Xbv4BkzFp0fJJByLS8nv9UnDIh2BnJDiuJUjZJxwsTNC17hhtGr
D9pX+6QUW7BduyY5bxIWPHbtqIBm2rHS/TlTtgmgcJzYaY68Hm7hTn9BnuJs0+j3
Ul331p77o3/QTTHTmS0pxPDOeAImqiUz3HO5HpnZJmNwLQXvp2t2zpiPtPQGtCgH
yBmhLFMg5eTfzHIqWbOZNgj1TYlq7+IjsR8lhINlhpMNOJVHNV7S6xtECBHStO0+
9giIwuHKw8IR9XvV6g9yfc7/rqSaNDfHlmHDNdDWezNqy3VXmqxYxtLNIPq8JhH0
yQ2C+rLjBIJpKQ3FDQRXtgfp3883nUBbV5FF4SIpEVQD4uxhr7x6bG7Y4z1Lnuk5
ff+dINgk55ZD0cUjjJMHntKsuCdaUgzDlGwd71FYimsboFcqhq7jJKfw5hds8QSD
w2a4ovcZHxrBwLROpeul8+IPFRXB7rSYuM7YYYydo4FCT4lFrEXZbMN6SNfCXSZX
VuwTJ42iSXh/8wV8TnULw8D0Fn44PX6mOae/S97IhKSjKB4bZ40+BkOVYHIR+BH+
Yf3Tu/+l/54tG27g9stuPrAECNLy+WNUB51RcmKPUq/Z9tInHEA9mHsia/MB3M4r
ZBO9p/Bk69UZM9GpPxgmG40aJxkfCBLf91nQYfWtFIgrWvwllMPGOiSq/X8jJRrB
dHZDb/1JTnTuxcqky9aGJXcrvv9iTEl2PVMgeII3CPnffHckrSpBFksw/VABivOE
T6PnVMDHHXznb/ufk/cXmNh6oS+guyO1HWFyX3xqhwPsymlEdcU9x56FKE5bH4X+
bG5PDG03SiNKEGkxRUaIM+Dn7dYMJ1Y6NjIlSjLyh9pi/MWJThX3b14PWSPTfpr2
wGuXj3tia1bYLeHcZtDmUPSsmcYbCXSSXIi/W98Ms38ke1a3iLN4YfS5u9K9Z4aP
VDgjVk1pY+//BLlhhMqRklVGiBrKggiCfXMmJmmF2f/aFDywELBM5n91j6/BLkyO
WmCXfOu4MgjiQKVe5yHvUBwKD5n0m5AmimomCM36SUd+o3w2hR7WbahDBizGwy/I
B5kyWFO7VhC8rARA0goJoY8MrxNwOfISZsd9SOlJFc9bIYCWyzdNJjxJ27hLvpa7
X7PsnS2n83ANXGhWdo/XwZPK1C5Lc7ansluZkUNY8E3enUoqsbfMHuZpCDYCYTqY
2z7duTmkdrGC9PUAsVAJ+tQ+INfQJCY4KjuYxQYhV2m2Y53f6tGU+fkKA1ISMF91
q3lejaEdsQA6XyNHFcdiSKBLp8i5+OV/O0j1hS3jVe/Y8F/rq3JMKmcXsxFN/mW6
dXLXuZJbDXPRUC0jzx5V2pYHjS9PpvTYpXdGVULIVKV51R7ckAU8gS7IfqTmXWfV
CjQYvdq7LuOgZkKdSmMWPH306nIX9o2MTN+F76hG7iL/PZ9Ne9vYsNvgz67tab30
Hvx2WCy4vPk1AaxR3EBsAtAQgLcga8maXK0XaORCcLDl22uCaDE0rLy1FYoDSlra
qEwICPkeEaQbNFx9MKfWHZxs/Tj4gMhk5NvrKK3bNN1eppkcMFNRR3o/bo4gmLYP
g33iCvQXDNUbqOI6L06S49DyCi3D5Zw3gMD3R6AfP93NFDvkG/6Y9bdlCKOQiJ9e
Z/S8VkgkYPkKAYSZjx1KH1L/0+acgAof15YDPtqITOkJo/4zVB3KIEe47WKxG17q
iwOk9UnbNRAkZ3wopHbB6y317g9y/ugQKFgl3eADhz639WZq8/Ix2KRs/RVpBKUw
aSXn2IF49bccxNPH6wyw9i0x+e7cJO951pF9MTo6Ltc7wL6gYIK6ZS2L3ylnpUWh
Ff55z7zqjSRJabmk+ciPuWqG88CPzVhJmYYIjsoQ1anABHkUQvX64ZVUYlLmIC6F
eUHvInduWD0pGLaEwApKOtE+yajkXx49avqacYNHv92O4SUqJ34YIJ7wkGuIXhHG
WIHLbX+4ZnfngLxq5GLODgwe87ygetq0MaXY1bq6wWJKjuY5ZbrpvpCo3jSYJfFr
VRBsV+xuGjAPMIGWJ8lp+SmCIl8/MzKD4C7I6WrQktFzIwFCrgUEoIfSPe1MxgGC
gKdfXAbMFNfLOq72OGGxTVFutAyvdn4FedsaQ6bt3W8uTL6HO53bBNqkblTfVvfV
0D9P9VUe9BxkkAtjn6DBSDwPqWFZ9FnhNZRWzNieZvzGNi/E/+XxP9kfAb9wra0Q
j7XIzRt0pEThughQeDsFw4uA3Dk6a6TwSNlDzIZIplFA3AhwZ9ZTwX71Q9yHL1wO
VpsbRRYYbtwqed7XnT13TmKC/cnwm29x+gerUyUdoSepE5vLKCqCxHmUaAboHxIT
PmQd3D5bcXRheiZKc1Rno3fYsBLjYkFVGFxXZc4G2POvMToLBrCe9NP6OzJc8Tyf
PILcoV/Y63yvmF+LuMY8La5CVtQI5CuFB8EFm6SGa+af8FDY84Cyu7rfAyaOfOtK
6cK/O4igUSdznNH8ClR83LuwxSo0fpUjCoxhyCMIhomrRceMDsq9t3i6hHlRM6go
lEVhWzAbdAqfpvDTaX/l1cSsLHEfqRgxxSoLI69EBjTfQBGOQkuDTK9J1UyIev5P
iszgoRzYbixfDMWXt44y5aXLGezCUjARasszOdV5fX8PuriJdu6/xpnlB2hi0B5Q
JPcrYckeIClS8IdzvNNgDepzzGQ91HOijayRSjk+u17i2jQAIW1sMej09RbhhDWN
4r0keiCrmnQjgXD1j+cW8DVygMH/RSABJm9Ffg+9ld24G1UuonOzLLDqx8sCmymN
8k8DOJ80MEcE+U1L5JBbq9MzPikx/8Rg5tvahl/NLM7R6thZK3aYf1MqvleEUqtg
mXC6f1rwTuoORmuBpYfHitdlsRPFy51UTCMtOryX0agfi8WgxVFqMkPpswCqmNoX
897aC0sNKo2rwZBzGSgaLMFohvyXtOhsqvTKytHunhPTh/GCZKqJuhQQtaryDb/y
LABAzUEoHAVDklPOh0r7PJivmQIjzXl9MPgam924sjD2tLseqU2h/RMK16Op/ENb
ZHXHoBYvvSZnYicBtT0YbzW84pl9Otn4xLKVFKhdeGbVE/86lsKOhmqPIX2A8Lre
WimP1uI/lvNPuFmWkuBQcOIzzutQvbnkv977yY2nRayl7w5lqJ+cmsHCykfPH46C
09SsUj0FB2CEEI4cW0EArijq2HGvafuQiYubViYfAyqmaGP/LdM110hOAOBWEeI7
LLCR7T5fDpv5LPat2MbFlSNsA6ymlZOE1G2fiarHwuy+uPNz3i/ion+06qjB72m8
aDPi21tHuYgJSAjPa2P3hb9sMaB3FP0SkT1rcP2HuIgD0KHpxorfe5522w3edoIZ
obexd8QlwhCpNJazcSmvYzImmLwct5y/6h4bEdrLtwm6iY69NJiHmctBaNu0yRAc
e/GgmNVzYyVPNCGEN4EjXoKw1qy4UBqVVg2CEao2FwlqvfgdX4pgms4+XpJEze9w
P38osQ7FYBDvB9Jx55G4J3N0tBxVk7f3xnoRiDMIlamw7aKD1TFhbGR1ge2qr9V6
QixK1bijT4dNGa7FgXU5/9PLgl/0s4Z9zwC2wfLvtwFXblQ9CetiWa1rq7M1MhnQ
fr56DW+9FA9PJr7WUxYrsTN8Rz00cx5QZNQHocT3oXkjjgsQOPDm2LEdA9VcIniL
YvqhBU6z1X2YObxem0Hn6nM2k3TVZefdppBaFPxs3AZWGPFYJxkUi7fZInn0lP8k
8zfIhW0p6++H/hiJTplrbDTgRMOdNuEteJxSJVa0DzMgY8OZLlneQucxe/RWD+Yr
UG1K770bYWqstCG/LxaPm+W9TKfHTT1siQJUXgNuw8yr/cr/3UkG9bufPqDlPp9p
wfR3MIXGw/4iiKVDW7YNoSnUVXuUrPbvq3srqtoxBDp/Qfqi+6tHsVZY1l6mI95N
C7OZ7cl7zg+4jpJ8C/nb4ni3GJEK9dOh98NB5tzdj+CS1pnBLQH0SSU7DzR3WVbj
70lVcPNwuyqDz+o8BFhvBn8wIoW7Ve0RkkUdEvULIofrfuh4PC1c+WpTUnaNtZYS
P8slT2cRHxNB4Oa5CpQYHF+6zoeL6IwSgZ1TIyxWTnh5Wj1qpquCQoWL6GtcoCVc
Q+0sqcJHjMm5Eh8R6+9Rzml5Sq1kzj2Tq9f6YcVFOByx04jhyFuaUno5s+QrHocU
9vvSWvXAwOu5T4bGxNzXQMlxDIOSSX8qhRuSzGTn+eOAteOFSlyGMX10RZ5QIS6f
EHF2ICh74iTLpsWBiP0ZmzKLtQT2Pes0nrV8rIW7GmoVN/3I0R6KUqNcDN3HrU+R
QkNwHOFKhvFp1FIHtn0iq+rwEi4M6G0EEIbS02xce6puIyjPMFZxedDOCYmwN5C8
L6hNZl4zlZpnGaPwYJDss8p8PLDfyIPhnz+++CO3O2SSEjdcuJctgcMpKdPMvbX1
Tl4f9Hy8hWY6A9fcI7in/KVlvUYHeXf+nGj3CqtSTEKWlybKHUM4xHTby3E0CYMF
EDEsyWaKcombNp7uf09TGudUXS/n+BO16rgzE0UIt4mb/D+4+fQM+RgsikV3xiUX
hwCStW6toPJb1m6tG/6bZl0vvGBAY3GdsBDDDgr5TyXHqmEilqT10sQAkVNI4U1w
9w21o8TXTCGp4/SmvPZ9kpAyRRV83Lu/m5kUnhK8aJx7C8nFwWAoiSbLpuL5L58l
TB0XTohF6NMuXF8asNOFHYOW1nXTSXy3TgGbNiUPwg8VS8pLQYnQhgo4yeaaFol/
c4W+4HsEwMwyDBBLXTUb+tlSirHHipvbAUx7DUDbQY3rhSHVUYr6dWzPQFhnkWm2
P4BheRexJ4X7HDZbCNONCxs/z5qh2x0hef0h+0YtzrmVEoDfPoDMfF4+bfURWIlU
Asey0KcmKWfX8fOpHGPrx94P6l8m+uLFfakb1T741iE2WpyNYNtYk0iAHd2ATSb/
nIAX03Lx09+7qyypiL/dOQ0hr+ngWUaRj7UQ+FppYLVgMSvfUe7QpAJEhxLHRVda
DiPxdM2xI9mldMzy6b3YZqa5BCy6F6qLk4dD9obq3L6Htsx5tWeSfVQENcxe1gxr
Foz92bAhKzZeWUhWAXmBCciEfG2oO2504MYUJIIWMB1kEbTvhCBMshUWI9Bk1jv7
hZsTc63PCYawxwR6mZYQI2RvNDsxF1y22EbWydQXcvp/DuutegnDdpmh8f1rX6Ry
KKcnWgFKXKoriqwHLS5zhWwgmTdNcg3hWBkj1INF4q1076mVyk1qIFII5VXyokZE
BW3qjq64Jh+DMvpKRuJO7oHOS39nu8c11KPL4wqx9qnvfHZTiVRtEa5v1ja/rs4/
vOULRKXLcnCUMYtE5kid21e9DeidGjws5s2bPWPVKBJ8DKObBmCalUuuAT+xRY8f
3MBYB8+anY2A4JOCym888IRYaV/PlpDGYXIyyDa5xv4wt7mY55Il0G3OYO65y32f
6kD7uZc8Q3up/bOf4qkWvIhAbDmJUoVmyXxh4lPuqef782R+gXULthi06yddoYTo
moMtiVOjE+IU2MThnEFo0pOrrlRoDm941WJJ+rt1l+tEhvAKH9kF4jSEFKeCAsGj
KUhzDYQzybgQVZAEPqAZJV5j6p9c6ACwRLzbMqOSXDWfvtKA/OzNL833Di2xe4Fl
5JmeDCsdwD47qkdnrzD0dstUWNeRhNLmozvXsaQBqztjb76WuF4KgwMsbGBhvWuw
TDQwd86dgpBHnrKWodqhIOGhl8t6FuWiM9YLgkM/8UXD3zByL2vHAoh5wbgzZJfZ
TgBFre5cT80Ue/vKxK+Gmc0OlBygrIFjRTRIqQLlusqIzjP6bPOfCK/iUp7fGQzU
fXgKWrHUNy/RA7jGiVMZwse2vlQZC+SX6l6NvdYvK0PSOwcRj76bQr7OUuHVTrh/
ChlEYjyimcY7s3OLDEfHRd0hB/JsMbZBbXPZ2jbO/0ua0lN8Pjmf/qxLE73oRkLN
lNjDCUZGvWEdqp9g5M+ZEmrAcxFqPbB3zDswVJd9XcnkYqNyHyT8iKTh19dy2T0Q
z/zJlFu2mB2p/P421jmvt03hPJ9zAT28m96W1SjDE6dMhW1bsKxQCnBs1QfmJP1l
de0HV2bqBslzOS9yJr8fPmnwMfewGf8ODWNzKhXlsOBJpR5G0QoOhyOMVehM9NEu
hYrvAOiqRQ9a6Frx/wqGhzrRXTZokzxDWKlUhIbXyop0RkxQcjvLrKvqV2sN+3NG
VLnEK4iFNYEH/mGjPbfRq0NQilPtBa4tW1gHP++w1OAwWnklrrqLgOlksaKhmox1
810iJ5f7pI+aWOHYouelaEIze+Apd9qUjUhTK3N6dXRzVFwCUXJgk2jpmlaXwkit
5nmXgaO48UhrqxdX73pprMXv9X/iF2rIMacchCAHxlTNFuVHkkuGnEbMFCvbXgkJ
qrpYNsCYIOGKwsjorZDspVUjX3LEuiaqMGjih0EOyes6hvfSq7/y6JzCHdzDzW8Y
LV22TsayVlSgrH9r1soahdRJLCKXeUnr21mf4FgIN1SVJXfi2F9hBxmvnqgHVpaG
KpthBFKtbFzYy09PW1IAI9Xebputc5Ah7t2LyVGns46dYsA7tHelzcVjZHMYCB/G
j/Eynp0zAiCtXsladrKmkmK9a4pUY6a8pbc8U3j1O2KtcqpC8LvnL24nMSj9zJVP
wNucVjXfVJ2iN8kY9KEHrlhJMspzxjoupNEp+DGah30N7SwGh6tYLpHF/9Ekg961
6a88HeBlDz10T/7NhHD1koSoNB0gK7Ie1Ux+MvbQG1JZRcWJEQQ0SJZW47flhvZM
3YacsfYdihuo9YQwcy+8bVNcx2r+T+6aX9AZQ3+gkd1XDpL+q8eoqYD/e6ICVuUB
86e+8KrBNfIOQBqZns8XpmJfSZ4bfTAo1ymX4bYvF4FHsgBRVWphtZg/Jo0EJRSI
X2ARNV4d+7G1vCZ6/vLIMerGF/4BMDrCFp1yhVvxh3VajDfUZ20xpTGCJQTQCnL5
W9Mtvl9LLQGWqE4Dy490a5b95DqxfRJguRsACeWgYddtrQSktn6SCa88SZMlYXx5
thvUXp2MIn3Tf0C6X1OnX0FT1UxZSSexfrYaTNH6lpJRd/DJAnf6NeM33bGKVLnI
mywb0+/mduybEDLoIiZQZlY9gLDBLdPc3XzMyjKKw8647I2YI2TqrIiO2BJtPp86
6nJNLKu177cZ7q9RltmisZU35llixzMlcYKQnl7k6ygzY75OFv3nSvtCPhnp5BK4
GQiAtCLqdj/iv/PwlooCK1nIELnmB1t4vfoNoaIxIB7isM7kcQbRhP7m0SmemoqH
F9tdbClT6OriqEUcjZWsO4zf8mU/aRqNiTmLJZ1vvtBicLhDyOjXWWt0hr4I9Fsi
DnCkhbq+4VVXuX8YI2c7qYGtB3GVNPWa0zBnylthumYBeewGz0BxgLVcvIH2Pt69
Rs7ZChEKJDoAz8xaq6fsbAi5SQqP6rZf0o9A/LTBMQ79fqtDjKeT+L3WirmtrZqB
piRDUn4iAlCIG1grcCc0WcH5HQIP5trvrPsfbEi5UTgwNbhklgLt8BKRv3snxoNn
Ws0b6szKGMd05CuayO8kkJqL6bx67W3nLTiTbPOLb+DGJ2V6cuJ16Fd55sD2Fiw+
ZjE3sBm0RS99j5gvcP7Xwb37W/UmtSLlq1sJxZ3tqEQX0A2uFW3ArKdAQpvg66tt
sFu++P+Basgow0fjAvVPNOdUgsxdqqmTxb/fgrbA3V+dinscDh31R0xlepDrGkvp
65PXKi7xCsHxfOaxeAxdWIJwz7UGB1yhnrKCgsJ2eAf89fqpYYBSzNCIZXhIa5UB
l386jMPX8+Ph5hF4VJzkPJSB3kDJWlQSluZfqDJpaI4hS490qqPlD34Viw30vwsT
KSRHt/uCoUqjbcLLvL1F66/3UsonxCKYH8kcb0kx8y8SwVx8Abt6PpMS80+7nKjR
uxzEP2aNlAdwrVYuE5I4rcy0qgrN5LYl2WTqxJW/SgyuA8e0x192LYeq9sX7EMHV
ufkXwe+jHu/9bfb99t9cWmB8pwIMp9kEcISTJwIgpDi+oxtZIO0XiM/ghAiLFaOY
OFOILL0AvJ2z8vO3xYXiqmKZs9uavfW0FTJnwv5Bj/cOt9a+SV/flc+371N8MKal
9za4KjGg1JWbfpvVbKEoVYvkYYsfWbLgHF6SUl4EmYzqd1t6eiSz9LfctN5fLQcn
945HnJr0IRSYwTBLHgEQ6F49X50pUN5WvnYkd82Idus5co6O6oL90WTox7fAQcVI
OWjeVUb1Zt57i0x/e8QK/p/lG504sQmo2N2IFDoV8iJALgF9WfCdDJHxAhI+T95b
eWiMLKrPfrapdtr4HNZ1ChRqYBpAfdePBG4MlsFCW2qIgZtm9mOtlRmDYf/LcTqo
btTen1GuVP8oSayg7RzeMGPuozziinDu2A+2zk21ADEcJxzHOAdnwSAot4pwjh9e
2T96y9BFvhXbmXQVjA01D/eDAo7oKDPg+nqIONH/i77flmuiFrbrwZ2ua64AlLAU
D6RubAlZ90MLgrtSvyB7IybhTZxHESX0S0G13QTNlxNDQYWM6mMnq4JOCeNN0Kxl
faZ80kVPpjuaZlQod9ULV1rUxbKwDs7bZWnkgofAv94hxudSFJARN9T95oxrPgvd
GuF5SfnAgvTzrBJmacquuRwF5/g+Smp4H7AnQx891nNJfEUVEIy+9QTnqyq0jbVM
aOBk033ZNrmcFwDcyMbojWTFDYZADqpm/2WpIAmFwK/w+V9M5zXuGMcvq1CFo27d
xQT6FkH+q1UHKwiwM/rMWadAsDBo8Mm1BeMwwxpV6NLDVQ2vYlcrRvstXjV0Ln+R
6WMi+dhDvJH2wzylpgXxmqhGW8WKXQM8sOq5VJslKpmzD+9IxwQ4WYgnrKHjS+jh
T6s/U2BmKxsKEOJ9pg/95YrE+fPNQGmZq7pJ10VzPstVwXUGWG/bFD3+ceas+Yh8
vBaZ/Hd+WAwORglVbMOJApf4zZPwIu7bocpfPFfykxDS0KpjX0VMcKULJNenEGcq
CssvUwFRkPE+ZWc4M6mVZ6FYULqDt1WPRypczbjav/J1y+2i/Is0woWeCnsFW71I
W4ZPv6mQtqbc0n/WQCr67Xj+NGXOXATXQyPVaxWuJ5eO6P2nZFyLRZZbJGocKjYZ
sYn1jef89goix4wjp/5MmD7m2PqzX8a14D16hSt/yePjAnvR3bC22key+ZdrDECO
1rc/iJaXHYjJSQ6G0BDQ7jbbKZrmVsu5pXB4H61aNMG0s3uK/BfsWFPLx0HH4xY9
bGVbn1gVpl4pIdtW/A5z0rgt5SDnXyb45leLBWsH6MxjlyV4wOA/Az8jrcUJqK2g
pLP1nmTLwxLxqhG0+ULLk8Ps/kPXtaYWhDO8Hw7qJ2PO/mtPeFoDPtaeQK2XMkr+
0TTwMzvTgcxrNanAxsBF/oedpsSt6vQ0v7kNrX6l4ht/7lbnnlYBhpuIB51384GX
xS1D7J3VxpB3wfJ7wC0L/AsKHMJjG2QOyPIXVqu6nTEOSpWVfD7s2/CYJb0I/czd
EEHOoa/mMfGpSShuN8wFrfEuX7CJWxUMlVshdEUJ1TVR0azaflOTEL8W68kbIjpO
FSs25Gos+bkwHBJqOGscCHty9Pb+dLT7+QKnrGmzIrAF8Z6Ntk6xugmTw8rWcvPe
KCrxlDBg0o0/+WentgDAOa/N8pPrVKNQx2DQ6YJBXzULDtgBPTlNz29xeybAR/0B
qn2rzmqMCa5OHn+U9Mk9P1YCaHtfWuxSmSPMH1z4dVBE3fkvbxRiEp0HS/DAoLxJ
BETGU/rfdVPSvSAuJ/ZXAD8+PkDCaoMS0MF3qw6d/t3xvfm7beTgR+3BwAbZ86pQ
I+4SpoaTT2tdwvsdVb6IiosTPV5eCKU5qa7Fa6nN2Y16IuQF3YvpVm1m9A1pobqk
2tYN5ugYO/rmwFHXZV3V4Gn4Fp8pPZpa8VPY/p+Tp0mkJAkD04d6pPKIcsOWCDUl
GmYpE7ExsHFnqrxzBpw7/c5Z4Ktoj5L/s8wLi22D4SodbMpOqLSv7Lg90x2Ga7yj
Mn+EOejfVewOugb56XJj/cz4GZzJ0PVlkLOA1XIWl7b0jIwuuc5otH/FXqg3/6+8
/JTglz607l5KJAZFm0ANvhzRkiPjlW2kMvTreRgLSz7SNOlHa/xWRRYBzweDHhK0
kdN0LniSrAkD39KeoB3bE7792gQJ1yOr1tMj7JyyUbMo2nLTln28X7LK6OWr9zH2
f0x9pzNgnxCBAG2qxba9B6T92hTQ5jNhm9/r9R5Cqm0a81Atksy6wVnlsNk06LAY
Sw9lLaa0IMKxzcFaxonQfCWz5ibCxj8CiuS5jidaJPsa554+itrsB/w5l4fOR+Kv
vcMbkjrSuVZxs4Ey61DW16TLzoGPEgOfrgU/nwzB0gtf8GqCDBrCN5uOUYkS8KnZ
5Nb6DBilTc5VIuraPZ1qCeknTVXuoVtGSRJHnKeE6nL8B9pB74XsqiXA2jeLmJv/
w/UiVSXoJPknR3hC4dzUEAinYNeuD6DD60DlOR45C0bDyY8Su8QWh2QfwSE9Q94H
W4XzI+8igeVmkBy1+L9j/c5uGVeoLHP3YeG06oqfMAuWmoCWK36446BacRk0hc44
hPesPa0upsn6eNyw+BqlYIAIZUpbT7GFFON6n3qcXR82IsPm9bAY9U01uPGStop4
I062GRZXqWKYGQ6YOzGJ4BIXcXGuCApbHWzJ//IauT67UKVQewLVmKPstXgPTEm0
5OBjiAlDJBx6VlPjlZpQGhv8nY+WBaJ2idhCMa4O/4aGFGIBwzHo4jjtR4jkFIM/
tAAKS58dcZzFX2ZFxsUonV6IsMR14gT62/LmrneTc1aqXv66YJ6dB8xaiD8JrLyY
sTdKaBhOyiaAQKzKLK3NLOJiSPUq1jYmxnAs5gwiI7alOK9RrRVCuitXpUH/35Vb
VsDuflMZkPZuHXkrXAua5cCwm26zBWpOFT0TPiYYVVbU/5JImLY6YYPPI8QEzcJC
rv+j1X/wAXRFi2Gu/tbIlzFQHTZeznEXAyPWcYwPcqjXy0yhy2TSlyG/+w0vzWEu
4+I7y6YyXr7bYmnp4JSvTwn3Oq7E9VXSsBfkiRFwFQZP5ksRLzhjvGWWwEMZwAqz
ABMZm3rwJbCQ3M8KBZ7MjjfVMiOss8ZdH0CEtqRMJUJZIYRo6NUmERnc2YLb1u/k
GsdWOWiSECBTLYCYkMwDk7un9m+g07P7kCzRkiPn1Gb77x7EReyUfmYjhNjy9zMH
zW43AwfFXNFeLh4zoO7AUEo3QoBUsv4rZ1BvYtz1Vzj3+wgXoi7iwwanWtYuAo0P
W2X1zDBg5QZDJgL95ksILRVkKcYBzEs8pu4EUictaBEXh098GJyLr9WkfA9cT2F5
dpCcKay4Fiqdc/R8oB+rKDFVYYeK6qeUhZ+rkNyGkpxZ2zLHU1mSRs6pCKhIIArm
13wXkm0Pr3DNNMfTWKLRFmfcMalF5g0mJlGKWPTk64fhHeUes+gdaxwcaVcH0CTi
Abm9gNeKndc4PwPZzKlvMEN7y4Z+qZ8OTzrBhZ1TfURtZpUL45stsg1mS9Ok0mHQ
HZWkVXVBjTAAts+uWUlX+LWknXb1/RmTGGtL7k2c+KyMg7hn1e0CmZBTedWgDf77
5T5bH8WlcIqKFrZYH5xBTmQ0V7FQYdd1xB77sSIs9KwFFnYEhKMlu0+uUkihdDuc
4bLSyrVmPYDH6fq2iDm6ai53yuP6MhfpTDvxYM6rUtXO/Zy0vwHc+moIOYYkCiy+
qjt4bmPHKRkXK0fdGBJU7vsOURMpj3XEHLFnM7YA47SfL0mIIThjjIEYhn+qEO70
wvTjD9zwdWRfZ21FNsujWR+HHw50xqqk3w7SmqdJS/l0Xf3P3eJWf8eIDItxknKa
nBoGEr9fLkA4Dcvl+XdjMZVkVcviNmuVt9WnlJbtJ3dxTf5Uv+wgvsLhe/TBLXJE
cSRJvoq1s3tINdYYHw9lmmi0ZaQy6wqCSOlnhh3aV2YW+zLdOZC1qcFmy5Pr+qCx
QfdAcQwxRPfZwxshbz2B0iEZtWQFovmhYIqRF+0xqubhQyrqiHAGUxo4/vlyL1IH
CAcX4jSbv8K8qqRgPxoAcaEm1EPBDaxJWH3Jo61TuDs20JjiZa+pHuPcBgFPZhvi
ez25j1b+a9ZK1nzxDigaj8GqgtdY9ZMsrj54so2tYLMeYkF6VpI1Tma8iK5i65bl
kobNcZs2vbnQ7jOiwJd43isb/cz4XENtNn9nVt1ZFU5LdwdVHBNLJR8vPGGUxx4Z
4CCWv/LWNC1IWYxNGGXpdXbxNcNrk/5AP8H5GsqMRDvPDIgtY19u1wxb4Pf0CneX
byOBQmqHD+A891hyugiIr2qGRyCzmH97wE5Us4x2DRtuqFOfaWBqrr7RiF8yj0+e
`pragma protect end_protected
