// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:42 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
tw8FG+WG/UCoFvrX0Grk/FKTC4KYpNqQffu0/9u9/PqnSmW0U2siad9v1WmDCiYI
66WagSlKOdootfaKzU7ifxW/CZ8xpcLXA/cwTONExsxN2zHje58KbQIT53LZUcb5
K0aqTV6xcut0ec9XYAhztliDFbuZicOpQHJUtLC1kL4=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5312)
nG5D/Rq9+aDvhJPloZfrVIbo+TezM/LL5Wc40OH7enMBKQR7E2FBxHmk1B50JnMa
hs77NKI8+SCLpQmWN24lPI5QbXLZcjxReGlzQJjT8Oy3xVxJcaBo1TY8+zgxg+zu
PfPfmQ4mdvwR5poeDlHJOayj1O8NvGYuJhJl8EZ5zlNRh7sDTcwK17om4Zdc0pBE
BHIFJhnZn8wo5BMKKX0IWfa7ETcLGEHSOEXNyT1G9l0wpIRkmFmYfFeiGjfT5m2u
QpqrA6J/CzwX190IsKeqA/pUmWesxWbHi70mtv6wnB9vbhBY+LFMYLROLrXD3Ks0
rAiHEUgF9yAKcBI55sST77O4zObenjiaCmPU81JUJ6HRlyhYadRH59H/P0LMPHAc
pRhHx/mtn9rDzxnc948gj3OuRmoU4+mhc55pqf88zrhqUwjZh+92BNyUy6w1fA2E
hCr7CISsX5QKr2NgKF7cTw7GTZktitzuSFrKf2Q+Pq2Lml7j0pPcsxeBhrsi+a02
jo35NBtd/NiVB1oxdnDigjaqFeyzoxwOxn7iODHf2IqBNlATc6XJJVZ0nlLbbV9C
/JTojNxCnUnE3IeBkdBNxwBUqErLSv9W1QS6O2jH6IaIaIHqOmgobDgqtT+O5mTN
f8XUFedCxz8SgUGO2wYgeleuFhTaOIZjQKeqJLIOMmm1uvLSQrMp9cUfHfqfE1F+
f2hhCsaoYmbXea8D3JCdQV227bblwRfAsjBVyVwgQOIVSwxR7LL5V7XLzPE24Zgw
UoKS9FD+3gQl9MozyNqI5RnjP2JBGGWDuRyyyIQB5udZ+ONjVfq8eHbOiUhNEyHS
IYpax2OevMMTXYH6CxkkVirTg6qDQNwesUHVpBZTkG5YcK2fvptMDaXxXorp/Bqj
I0OwfqD9JWYArpdT2Vc2FU80v1ushO/EoSAzrcClZ09JdWuUUVhY6W9iNTMo9VRO
3z/FtKynt1nTOlmAxDCpmlPOQYbmiWxupJsCMke9r0c71PaBKryw31m3cmG8RZO1
+juJcw7O+Dz7dcCgfoa7ZURwpTJd/nn1kyr2QxACsRgki9PVrOmYlAagvA49u8d2
ErO9+kJ9ObZc0OEeN6YYfKp5ngXYWWl9xuBivUMkppuDi7Q/p8vkPhzN8FbO/8TW
rE0qRX6eS9E2K8786i41TDpCdOx2W+tDqGBcHtDWxRH8RFLgFEZTbSnwlLErO8K9
Pu/Q+IG65Yw8JIcG6Ueq51GJnhyw9adCrBuEHXnZQGOLDDGhNPGwTxChjDsglCBL
xUKd2fKestDIxzlAncuRgQxft1+a2P3vsLDkY9C6DRUpMEAgMpleKxhfa3AFCkvJ
dSl+LO/uhA0Sk+tfhc9i2729EJ3hm2FPUThgBHbS439JpV6fr8iCb3VHN7u4R+F+
hzJcc6WVNZfHuDlZR8GHb6GbN+LFWk5ceSZtN2JkG3XoWUrVTkBzCESohftNR8+e
q3MCzP/qJOzWtHLC1JS8poYRBXu7cVzZrhEO4cWRYhUeHmYFL2rE3ou2TISn5DlG
nxmk0Rv2qHq5rzXUuHv6HbhrQM4FsXWnixLOGdbB3eMD5Ev51mjVhez2PID45lx1
U2MNTZfLFkSsyyaIAoZWYlvGjmeS3tn00vOicu+u76RZjdQwry+76FzsqwsqeKUT
WxW5VdBBssCjK3YDUexY9IvyegqUItbLGYWefMBq9SmTXXfLG1zsTpCTi5QmdsiC
MskRCrxNoQG+5nzRlV2i5PL6Fc/SxJIN9vxriiMBcN4lzIwbhuoBxPyoegZ8f4b+
Pg+zw5rW2zNh4yG0458IG9zuCK3K24tRDNa7uVpFwGaLhaxmolEzyXGsNYqt7FmL
z3sHja12GI6/K1Z6U4FWO9ZqDHrydNLCpgYZnm0pEH8QF17Cv8VBkyOnqDLR5F11
qJwl10UeVMwR9aKPtZGkcL4BgycquS93R3tper0pvtgt8QTBXTzezQoCYzUsfHfj
g//4UkTcPxdZsW1VI+JGXcGhrXtI6ql9WSZ1rAHOyP1LkIArPWgluZoHLE4Ke7N9
1msYFKj4ftGfKJ2D9RmFGsSisD2iYknx83rKS3nMU/xcoypH0yHbMi1lGCB4gALR
aTkNlVQ86Me1hh6UtDvZtdqOHt3pt2WYtUMSKVKKyGHUizRfKoyBkA0Rtop+vXZ0
EJpd7nCOHmRKdgUQxEtaBtf6e1j9aLSdHggeYahyY4jvxvGK4LKo9joky9/7kxz2
Ea+9thYYfRbscIZEGT9iOgovD9Jz4i0MXE4dTr0ma+edNjU/MSe4FS/P5qkXSVcW
1dafcrEhieFYYlobINfG49pL8oRPRBSGn23AW8mvOejlKNBU6S2/yXYVmRy7p3HT
oJBRqaw2NjAbSEYrTDL7DoQshBQnACQVRbEgTYJIcgCo7h0vvqMhc1gToZ5AginE
TFByF3bfqJxANQFYP9kQxQxe3am/4jSNeCxRYeJzOaeM+X32ByqAhWXx6WVIOwUY
ZcIb3ki6Zut1Zz50HOr+9yTSkpGfIICizmWPDDSj9+vFg9ygrA5jCG3kL5257W1k
LuXpzyMQT2xGgaSRPcrmLIrcYTwHAQtNmjytiAS8/oxJCTyFrmtgHU0baf2wWTFu
9MihIYU2OuGJ1rr47e0jc+MkurjzKkSizwZ/j6lQvP8vZOTTN8LDkns9VDUOt5zw
Q0Lto6+QMlStOrTVTkqohNc3LHt7c4c1bcnVH3Ygo8BQTNj/y4IvA48HzhhZgT7o
5GqTsSW6HIZ/d9C+5Yks1vUfN2doxjwGc0RftzqQQwNoNVwrgh5mQXV6Rp7F5e2g
4vAZCvvwTKffmFM1rYmiI7W9DuafoZpib+7r0tJH9lMUM82EDyJ17mZasygAulf3
EC7xQsIGwQJaUuzRgrtKazYp1oan/aVaruZLXZhZQw5z+cWkdsU6h2H8vpizYZX7
i9G5oX+wJOv5EnS9Lozn7lzgCQ6DbbpbPW6l8C8DpainARlaJ8W+/1tqkjvIILm9
U6PSh1emHprg+RegAqt+CVWS7RueLNfx6VTKNCyunrJG43VNLsJk0sceXL7XBvhh
GDG56LL1F2nJIftkvY6DDJ5lZoisdAFfrVeyLu9JnzBEFqGhNb++cyYCTYAiIcIw
+bqbpZTfcKGKhnNOHQf07xW0nRlS0xPzmX5ekUJXzMNBuehB9zZgqlOZlNQLM8dg
bihdjO8aiwmAxGzQ52OeoUz4FedCbKHWeFWb2P85pHjpykSwogNSqsYKLuiuXep/
BA7IbAekEgHbULJQCnYiqxfOKOr/Te987m9WAA4apSdmiIs3zHUyriOaXiUTLgHq
Opps7TKeRXWZ/R/1NRSsnbPRl6hsVEJAAvUEBUL8Q0b4saXQj8ZNnhHzzBquL0QM
R+aEGd9gefaI0spz71AbweVzUjjSLah6wZW7pCHF6W/Rt/p7fA2EPuSVuocbCIHL
SAoiuS84rI12QnligexZQcyThx7NU97LBDBKY/Exj5DPgnq87qItM1lmXeW4bqb9
dye+nmYnYl4JdIDxB4+jdRwxG0qzanW9BYFHGC6tr/3r8I7MMLBUAvAUJ15rhLWn
fh7CPS84iPV2dWGfJzwdpmEtjybStvQYzpoOwcS1+sTr+EQc2EB3vnGfj3qJMFAy
07VSae30gs79LLighCeOk28t64Fn8AAoEbd4N3FLoWCz//mKfWaIbaPIoV97aKjt
1+yr05GGpHP+lpCnO6DBndcgRWMXVn6ez4+2HTBh+TXEeCa4J4sv96c+HoPZdqud
Jplx0BEq3vRSLAfzIedR31vcr+YAFeDBv09m9B8EwxBPYRQfajQlukvQu2N3K7xm
iEMxp8URzn0wqOfUmpk+/j20r/DAvjMY/Y6ODk9hUqeb3/yFAc0jNday0n8xL/TN
WnfCdrSklR0+8spp50Xi9RYpoZeFBoFT2zpxaU2y7hybtHzbVytve4Y4CmZ6Kr8V
y8SSyhVpU+ckfbeahU0l1pM2krJUo4G3IjH2UEbmjxkJ1tIYPLlcqlJSUEbFeqIX
GtQYD8aaaq+Bwd7wsFW8BaJ6jeLf3kSznpXmpKTefpN5MqgFQgaT5hMVR1oKEzbd
8VLIYR682EgZm4Sqpl9Wj3weZ7gDYG/fO2FNn0njMIeYcKUKUWx0gPY7+0KlDazf
QWYAN/B2LE7QpeFjGKO5fh7WOdlvc1xLpfi2nIhw42eixziXrdMvs1BZiNTd12hr
U7lg76owzfkS/da2QNur8+yD6zYozeEs7QLzzr1gNnZZftaUkKeTFIYk3K698rB1
vIDm6PLLM4bNXojFC1RDrdJbSagzvtpy0/7RQ1kXmpn0z6Wr6Bg/WobnnmtaO9qE
A1tPSQ+N1Dsn/INSZSzqU5ffkftRVJLaN/Klj7+TL+PyEOl/L1ri+ITsA/88Yp6l
wNJ/qZVemlZr90TBsCww/cwBCpfGahn3FRSw6mq5q5GL31YeZl1EVxjSLOMknPp0
DChkvXQ6NqoyFiKJhNhfgkMBdouPkfI1lRpEFYqrHEWt896tIDnt2xw8v4L4nQkG
0LqbTWUX/gMUvaEXGK2tkDhPqAh1xnI3rCNWipELPjBpXQP2i9Mvtq95jfXvUdXY
vsJtBWpOrCd1ZSuEndq7UKtYEtmOfJIHHx51LUzHOUjRCsVFjyUuMRriSTtN7qR6
eELIy72007dZwLg2ZKOElhsM3BX0kvcDF822xthnW3ysTz/juYunuo7e0Dd2disA
sdjeXlmxRF1A00wT9N9F8AgsHIkxEbbsy9IxxIVhDBwS4MEg/CBSrb65Bk9+TfR9
WmnsnrpCZLzGJRpYPdBqY15+O7ar0yaEgQ/1461/PJuHM3ybqFpN6oXjBRwtK2zq
vlkGzcSt6cjX3g6zc6mfF1inEmZ2V2tzLOfIXpQ9G52L0vaNMqKRSGhMaL0A7gRV
itjd+GVy/ynZ7k/ClPJu4Ljycoflua/qyIXwqKpm16TXAjwG5m7xIMOBYx2eBIvM
aFPyHty20pDNg+iotZTw0+/wbibaN+lsQXKC2Dou51Nk0/Hd+LeD4jgZiz4Ai6yg
PzobzJg4RDYdjADaj0JoJUJynME45ftY6Zk/EOflxRCJN13axIIP4kcfShU+YxDs
w5BJhaO80fDnsEYIpnKSsfYxQp2YLUI2e2cG3LqeV8hZprfnlAWeQB33vhj/U4dk
+gcwKGwd12MxprO6tbif8pWHYonj7h0+KP/6HdG0MjrLxvm/bXZn6NpQSLD1ATi/
3FDDY/FValqVR3OU9gCeWRyBDHbgL3f69j18ngqJVvDqt2rkUJ3F9SPXMv0IL7He
DpoG0+Ww1ww9c3s2vC4hYy3V1YLqgKzwMhu8BztLdgbPxKIBRJESV0MaeJWA23mO
MPnhg3y/SZ84Bus+mqkaWm9PhFxMhEMezK+wdUzXavXNX0k5d/lOj3ypNI/wxsD5
+oTGhG12HR5Zznjm2S+GA+BUH0CpVlddSlwfm0UlWXjTG9f7YB4YHY4PMweShkFa
Z9uo9XEUqofiEANdOou00WIw+LbZ08tPv4DBL56Ln2tYrZjkWnCPPoE9/hVwxdM1
9dq3lwzdhtFkawX/bLjYnaF5Oyt1DRjsTG4WAUFDJopoaW8c102O/i2dQ4sYvjwo
+ShuDYSg6RKJF6/cHZ9Rtm9RKNJ7aswBIOqGEgFMgZ8yB+n4PZx+iB+Hjzcv0r7T
7Tgx2RNFnwiPw+o24Ks84VUMD/dA7BhHC3ntZbgKEswW6riR1S5bAJzjoo+V7X63
qtE5jDVQEVurMkoXdRzJv65HzYQZwbYBhZKqq7W/54RYMzK4H0vSiy0zsJw6ame+
ZTp2tOJ6om3iAtryy5/pLOVcYUfAxMMN0VGHIn6QlQy/3R09DBF6BxJEK1YjUXOy
kTPHji1vybjOao9WUd05SdTwlp84/6NdeCq6wQKyHf9Dn1nk4my4QH9G6RpryQDh
FMqHKazOVJoe8z0lsN8RYuxMH+O8ADZgQwsxH8yzY7WYoKny8P0+/tOXMsh0rdQd
iZ9E6Q9ER0dUgFrrzDU8uN8M1wCjIjGXTCexMZbm6Sc8gLAiSsrqRug9L1zul0zl
ZJIsIFKMEdvUKTXpRDsA7EktQDOCznDHrkfBu2NkYHnA5ikBVGZvYu7wGPHQ0swG
n9EnEo08HXPCRO25nwrfMVI+acAzlj9o6C999dX8KfBNyCU0iYY7PVyPakhAiGD4
FdovMF2msDb3p6fFCCpCPNJuz3Bp8B96ican5OD3nNWBSV+DHo+B89b+1V9Y5x9Q
I59WqxUy+5nV+fIXM0c5CSZ3A0BKWvNHURzcfyqA4bk9dX2ksU8nVKkmCQUoBhAV
lhfxvhBNIo8ionOGd3iQPWJjtw5D7kcvKUqtA3J7FI2IBbpwk9wJDCEiZ6Im3Jva
SvwF52+Ro8aIDm2+hhRgoXzmn72E3QVPAHjwIi14wfVxVDJDymAxAPbkjQ/3zi2s
S3VjzWm9pjE64E/ap8ymlWb2ClUCd9go5R82TMB8RUC4bj2wzTLfsejP/z+/UOxE
6KzLpGegzZxogndNz4nX5e9uaYk97684GF27wnjqwp2gkQAYXiRZkb6WDXLFYSiO
DzzEZuJ6VCM2ivRhPB+xfyvMmUTDzSD1ZnTIemJKnXCdRCVmm3VA/NGrCm4pTv1C
wDmldp9Sm1ZLuhd7jDVjuZMxTgkK6o9RmxEg5KfWPAmzlYbO8tmKGw3iaczcdY+P
fHNcrdKdIUXlW4OM4z1SpmxHOfD0jcnc7Nfv0aoocb+G5KpySK51v14gFd4yuRB8
kL3pe3/y0BRbSYofhOHkZrV0AwR8Mfn9/LXGmM6JWlpDkMwDuagmKgJ1dLxdoBN2
EGk+Q2izuDBoPe85F1rfU5tcVnNPtQWdJ5H8OclEyXVFsEd4us0jTP7QxbV5U3+c
vrkRm6ZtmwMQzGmSJPoKqiQx5sDBhMnIBXxzlmaWH0JrbKW5+wAC3xjDX5EJ/K5i
WtdTGg5F1IuwKEDdyHSjWyX0hD2LQhb3zU+kOK0c4NiXpdFKKDM3TsY3QBf/PsZN
ugbuGgz8oLiVtPAUIO5x9RSlPjuE7+IE+jJ/3nN66+k=
`pragma protect end_protected
