// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:39:20 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
lefNl8Vutu8hbMoxb4OAMkLI9Pmw5WD4uBM6gE23JWGaUsufQEdW6ADPJGMHj98g
92dLe6DPZzEynAa0SlAFQtPazGZmSwGZbzoqhQvvrdeTVTzUi7i6jH9kA8UYB36I
r5YLq2GLGEpxG3JFeTvJJB6vFP+ZT1A1N2IBCKtKQ5E=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 3424)
SNkP7/Kh3N2kmq5WAyyIT4ONzVcLKQwYQ/DpEJ+nR60K9r+K+CbXIkfYi811DWTW
AxhWNxQuXlwbtNhkQ9W2Zsw7fmoYQQbacB5K/488QOlbBRXnmlEZ4ros5H9JjXkC
7k2GzGiEByJswLXdOvorujEU+oe8sk81V0uMEDEy46JUzt5Ldpt3tNp+kpOfkYD8
Hvk2R8sRnlEkNTYdzPqbXuHD/SBHwF6ewkaVmdsTNE4e+uYoCLA1x1TnlhRJbUTb
oTjia+LbO9LXHz2Lo3iUPHOjVZsVqL1INSjm2a7Rop1WjM34Zayc8t7spohL4cwX
qn+4f9SqiVaAXjaf7PWkO4+ogQSYDnpbYl+IvpS6FFD8UuObVFf9yBNBAf7eXEnx
YeCTXSGZahZwRp3JunLOjHk2IbR361dN60EdQBGvEkdZ1pVUFPRjp+Q7aRo5OGMW
NVjWIrpgI0W+FNp9aWPTngaJGLNquvsEgfNKYOM2mQBBk66uLfrg7PDcXEWk70w5
In2y2dV9nWBQdwy7YTBmSXEQJxtNyUDjvpFdu1XeW2up9Fxu1lqqnA9iDXkbm2av
hPxDW474cqVrjRq0P1R8F8uYpmoKhhMoIU4OurUiKlbvkDRYHnncmruZ+KgU09Ui
EL2QNvDm3kUvpgzucgJkIHkXpXwonWt8KfWkhvtPMsSlgdpYsfy/i5WSof0Wyxdr
5KygRGkJtUeguJQQVfhGiJyNc2VRwkJGLEL6PrKzH6ChPXi9Z4uctH+DsnV3YHfQ
iJa78TPDvc7lvHoNpnJ/F/3O081ig7+aEbCZfhtjAEnXXmz30uaUtKcZFVK4Mqqz
fLvL3YN8F5aXsMpNwsJSPcPwv5x29n2jfn+Pp4cIqqX463reeKf7wXMTozllzTzw
Sr4TJV/dLUhAE9GsEQt58Lf0Tvs8D6NhkLgfKUEHc2EudZE3W6O69h2vth7lg1oG
xCxanDfdyXJpqU0bw/n/ZYjQXYKRUtH8t3wrS+Ypl+7AixxMnzsVque40cXWj4DZ
E3wTgGP+udEx2ucpzQghakxtMZZZwMZaNhXkosCX90qq6TrILRHwGJsRcAu6P7Fg
FHPrUNtZFoil4AKQRWkg6hBpN5o5+w/lcSRnw0/BpB1ch9UBNNwnFDb7TvBf1lVt
I2mztRPqV8V9uwjuBqKkwq60hcBB2RHAan9htUhBbxjgDCKSxpVrpMwtyovHM8Gu
IOK8zWBno0KCxpqnKWNQFf/6yREpeCnlTGd0r0tVz1TnQLTj4NNYI5zB/EhXKcyr
h7qnD6yJllQp1CjAxvzw/1F2vUFbUCFYPnSMvJaD4x2LPn3/A2jGgPlXP0hDiLog
Nt1E6AEf5HmQFjEIUf8nRZLn10WX2eqLFms7fe7QQcr/K5+xV3gYI4TBbKhLtGAt
zK/ElWr64Qj1lubicRMiKuhCFcXM62Z5S5ATOsn2rIGW9kaMXEMkf1bdZ3lepHjH
bWkQYTyWCJBh63/ymm29wJQ+IhBjTDyvJjWf7KdbHKSkJ690nPoHkxMt+gIVy5FF
WZPsRiUEKRXn8i0GoGhLSD73NY3L+iTGBpdSx5Ifw5yOkDQ6mMDCFj0eNqhFX02O
C6Hz1jaG2+rg8kXuQ4K7dbr68K4HSk296PPSBSPW45cSfVItDjLxh5N3wQ9lUfmk
yT02VHq6m6X6ARMHb+fZUq9DTkxhjmgq4txxFkQNSgtYrBov2TSZwPQNAsTZImIw
r90wcUDOmkrqEK/u2EoakIZp7Iw0KnblHRuwqtSBMf4iTq9eB/oa0v9VREDYInuL
w5d+eGjpeDcqzea3ZkFU4OH8+9vWKvCfA0S7xUxhWTCwMvMCSrWiC6Ut6TuTsw8U
cNiCAPlHecwWWTrY2EkpNJ+wvyozcLIJshkQXCtSEeP71H+E3GiXhnUbtRzAuUUo
+jpnInJP895F3FgQlM17JO68Lf1jaoaHwrzHOEv4YPe+KwQY8RN6vpKWPfAfJhe1
qHiLPK6RiUSBn19dUdU9RJLqahQRI2zEZKBlJQ+7L0ROntFVnrgI8ZoQww7bBoDc
a0lmAaXmcyD8Z25k4RU1LFK6lkbbERuDPorGvOBYvb13MK2L5yyS4oq4/Lxn1XcQ
Ko8yx7QLcnb5/mZ+7YD6KcbEZyJ2W/1jI8Xgf1qWGg2D2P/2/xK7/UgkoU4i5nGH
lJ/0u+25dFvbwJbpfuiqpPFz7iwLUP1DlBmElew6ZsrlI8MfG5M+0TRqr7MrRSUr
C4VJS/snBWv1tTcqt1Q1cgpXWiScn2v7FbvuAZoE3zbdkSKxUoulV0pFPf0312uj
pRbL9ZB9fLfLWnpdqPJn3u7LW27nN8uXqPUPmHV6bBJjo46azHsRbXcd/enqe2a6
WgjojXUPqRKaR3MnPHxc5nnYFAESls+O89so8LdzbUDZAFNSZdIIIXBZnf9ScTtd
FGQ4msuyo9tAxdajd1CbDyu9UF4DghGPhzYGKaGj8t28nwFAdcPS2sV/TrYxUnNV
JHvOHaSrA1LSIQt372nF/tXbhtIDEL+JaNW9ZT06tRSN13OGrCRZznzOCJpy3mdf
SXRfvhWzK4xD/xn3fDQwn7+nLmcmFWlnyAXivH6Xm4iLLLXpC6KGWy32XcUDM73c
umbDqb4oHlOFB8bxzmQV5ilcBZZsxnfR6J85nv4rHq5VyzsZBVBCFLo7qk8esF/0
BymM16p9GgIR2sEAB1pzG6QdFbk4IUKf9R1zjfbQobBKUJYqo8bADEdPVXgUGZ56
NLlaLzjG1fFWKjNGKRTJhWcT+v6Uf4yJPPbSoPIQb8yrIa82c9inBnDmNB5JNO/U
cfP21F9SLbJSOefgxl7JuHlidEcWuPQGLrybEnWtinerBRZnBZddUJj7tKk2WX0q
a8UkDlNYvAbonpBgsXzFec6LKeWphV+1GX+8ox3U0CKY9zASD61oPCzQmZPOzjS3
P4gg9sL0Rgg6qBQ75YNe0eeSzvJjHSxUgD/7ad4HMv+9vDl3TXdkWFh1P98fFhrz
C8gIpEy+WIJZGLQLTK6u431FB2zAwxkmAdqB4A/a5vSHUQ4/V4bwqIYYNLFPjMed
+v9M3W1tFcxeGmLPkCS+LWgnSAFbQTclQg7VF41dCVHAiiVbU2oSEA3HtuiBFHmo
46gVL9zxTDiQ3ehEjXCe/r4HT2jDo3lOna+vPIYaTlqIhIPgpslrDvcEdrzAwZxR
wKfOP9m4Tx4j2+0d6FbwIKKma6iWy+YXsqFK7yGKu5ETmRu4hjlsFAfGGHiFPoxU
c9JZEABsZEeQ3rL8InfL1CXu0iQaa5KHuOAc7Kwn22szxYn5N/3QIHNE14SG8kPO
eMvFnzDJMwheGIFsTc7mqPCRgFU7TgpTXaZeIlyWEaIBdDJnvAr4ndzhxGOHe9EY
6Q4VQBR/GZbSyQHVATYz3dqzlaIuJgiVZgeKmLfnLiGXRqTikRGSdBd4pIuupqfn
rEfwp1oisPry9SEqTDq3oAKNgHJb5YMkFWcaL+odnplhpeWJwimDDnOYC2uWknOC
jIRTWQOLXL/ZhgoVIhjxog5QD0tn0l3jfgkAYie1LmYMu8Y59cVAYW9JdC2qdctu
J/x9Ulxw92Oq1pLdp9N+o6+8RNQ/uvjLTGWS8+WziSXNLeZ+Dc4ffSY+LSX+cgPV
g6/5jv/dIZVt0z//YzyOoC/d+HKBF2rHf2hRkW22WgakhFJvt5My3yV5WQ5QTgne
7wJmlLE2Kos/0hHsv4FukQ3uGj6Ioz9Ki1thq495OnwMYkY86FphAMmNsZsyQOaN
upstCH4dm27egpmzEavWrDnlNkkbzP7LyoqBcc4mRNlBi5xTqssl4Oawf9wDEsWf
8KcoastQEvZUl5pgHAoelm9OogllWLkf5TyX4tVdmjtEEjUbIS8k1jNwrlaiCvcm
P4VWRHNUNVFBRgRw2Gwh1LMUt2xzCGOFRnqrqcV5IiTxz+qhP/PsqyWDBY+dtKvv
e12zFHrPVnGmvEVXLxwgz0KCfyUZyTcKqX4BpATwUA67pXWr8IlWobxj9ybSlxdj
A5h3O+73Mv1Mc48zZwMcV1acsGy/bvU/fD8GPiGStDFxMNMPQF13TVxBRK2gU8m9
LXbgX86nmuXWJV+m6AoWL9bo2uJfHj8dhklFr3u5YVTNZ37TzveMFMEJdnKKySL0
wDjKmlOKlSUQesKgqz+e47nBhdalo+qrCbjgdO8+KYyEejJXfJAfW6F1nXSXmVwv
Jla/j62NqI6o/fuOacUGEqSM1faUeDTIPKEeZ9k70cNkPTk/5MQXrIfxRyIrexAu
F5DtTsMxwHhdZlFJ3gGoCv4VTQsTuTZNpNSE5YGk4l23ShxKevqOLG6D/Q0H4Q7n
bjNIc0iilX5LrlqXkZZdO1nhfcP1meM9Dx2VnZAfsku3JXkd9umJbbHUWYV4eiyL
kpKgjlHKQecHKDd3Xa6m3AsThR99BwuLVHQVKxdkVzmvSxj3pUyCcS7TI3mPDorI
yTHJpqVZPfN9IpVID2+UFFptK4ub3O1M401Igd/v5FiKh4wVa31gF8ahCljk/iWP
ViH2Qk9p9doooOMF+ugJQA==
`pragma protect end_protected
