// (C) 2001-2013 Altera Corporation. All rights reserved.
// Your use of Altera Corporation's design tools, logic functions and other 
// software and tools, and its AMPP partner logic functions, and any output 
// files any of the foregoing (including device programming or simulation 
// files), and any associated documentation or information are expressly subject 
// to the terms and conditions of the Altera Program License Subscription 
// Agreement, Altera MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your use is for the 
// sole purpose of programming logic devices manufactured by Altera and sold by 
// Altera or its authorized distributors.  Please refer to the applicable 
// agreement for further details.


// megafunction wizard: %Custom PHY v12.1%
// GENERATION: XML
// oneg.v

// Generated using ACDS version 12.1 50 at 2012.04.24.14:58:51

`timescale 1 ps / 1 ps
module oneg (
		input  wire         phy_mgmt_clk,         //       phy_mgmt_clk.clk
		input  wire         phy_mgmt_clk_reset,   // phy_mgmt_clk_reset.reset
		input  wire [8:0]   phy_mgmt_address,     //           phy_mgmt.address
		input  wire         phy_mgmt_read,        //                   .read
		output wire [31:0]  phy_mgmt_readdata,    //                   .readdata
		output wire         phy_mgmt_waitrequest, //                   .waitrequest
		input  wire         phy_mgmt_write,       //                   .write
		input  wire [31:0]  phy_mgmt_writedata,   //                   .writedata
		input  wire [1:0]   pll_ref_clk,          //        pll_ref_clk.clk
		output wire [0:0]   tx_serial_data,       //     tx_serial_data.export
		input  wire [0:0]   tx_forceelecidle,     //   tx_forceelecidle.export
		output wire [1:0]   pll_locked,           //         pll_locked.export
		input  wire [0:0]   rx_serial_data,       //     rx_serial_data.export
		output wire [0:0]   rx_runningdisp,       //     rx_runningdisp.export
		output wire [0:0]   rx_disperr,           //         rx_disperr.export
		output wire [0:0]   rx_errdetect,         //       rx_errdetect.export
		output wire [0:0]   rx_is_lockedtoref,    //  rx_is_lockedtoref.export
		output wire [0:0]   rx_is_lockedtodata,   // rx_is_lockedtodata.export
		output wire [0:0]   rx_signaldetect,      //    rx_signaldetect.export
		output wire [0:0]   rx_patterndetect,     //   rx_patterndetect.export
		output wire [0:0]   rx_syncstatus,        //      rx_syncstatus.export
		input  wire [0:0]   tx_coreclkin,         //       tx_coreclkin.export
		input  wire [0:0]   rx_coreclkin,         //       rx_coreclkin.export
		output wire [0:0]   rx_recovered_clk,     //   rx_recovered_clk.export
		output wire [0:0]   tx_clkout,            //          tx_clkout.export
		output wire [0:0]   rx_clkout,            //          rx_clkout.export
		input  wire [7:0]   tx_parallel_data,     //   tx_parallel_data.export
		input  wire [0:0]   tx_datak,             //           tx_datak.export
		output wire [7:0]   rx_parallel_data,     //   rx_parallel_data.export
		output wire [0:0]   rx_datak,             //           rx_datak.export
		input  wire [1:0]   pll_powerdown,        //      pll_powerdown.export
		input  wire [0:0]   tx_digitalreset,      //    tx_digitalreset.export
		input  wire [0:0]   tx_analogreset,       //     tx_analogreset.export
		output wire [0:0]   tx_cal_busy,          //        tx_cal_busy.export
		input  wire [0:0]   rx_digitalreset,      //    rx_digitalreset.export
		input  wire [0:0]   rx_analogreset,       //     rx_analogreset.export
		output wire [0:0]   rx_cal_busy,          //        rx_cal_busy.export
		output wire [137:0] reconfig_from_xcvr,   // reconfig_from_xcvr.reconfig_from_xcvr
		input  wire [209:0] reconfig_to_xcvr      //   reconfig_to_xcvr.reconfig_to_xcvr
	);

	altera_xcvr_custom #(
		.device_family                         ("Stratix V"),
		.protocol_hint                         ("gige"),
		.operation_mode                        ("Duplex"),
		.lanes                                 (1),
		.bonded_group_size                     (1),
		.bonded_mode                           ("xN"),
		.pma_bonding_mode                      ("x1"),
		.pcs_pma_width                         (10),
		.ser_base_factor                       (8),
		.ser_words                             (1),
		.data_rate                             ("1250 Mbps"),
		.base_data_rate                        ("1250 Mbps,1000 Mbps"),
		.tx_bitslip_enable                     ("false"),
		.rx_use_coreclk                        ("true"),
		.tx_use_coreclk                        ("true"),
		.use_8b10b                             ("true"),
		.use_8b10b_manual_control              ("false"),
		.word_aligner_mode                     ("sync_state_machine"),
		.word_aligner_state_machine_datacnt    (1),
		.word_aligner_state_machine_errcnt     (1),
		.word_aligner_state_machine_patterncnt (10),
		.word_aligner_pattern_length           (10),
		.word_align_pattern                    ("0110111100"),
		.run_length_violation_checking         (40),
		.use_rate_match_fifo                   (0),
		.rate_match_pattern1                   ("11010000111010000011"),
		.rate_match_pattern2                   ("00101111000101111100"),
		.byte_order_mode                       ("none"),
		.byte_order_pattern                    ("111111011"),
		.byte_order_pad_pattern                ("000000000"),
		.coreclk_0ppm_enable                   ("false"),
		.pll_refclk_cnt                        (2),
		.pll_refclk_freq                       ("125.0 MHz,125.0 MHz"),
		.pll_refclk_select                     ("0,1"),
		.cdr_refclk_select                     (0),
		.plls                                  (2),
		.pll_type                              ("CMU,CMU"),
		.pll_select                            (0),
		.pll_reconfig                          (0),
		.gxb_analog_power                      ("AUTO"),
		.pll_lock_speed                        ("AUTO"),
		.tx_analog_power                       ("AUTO"),
		.tx_slew_rate                          ("OFF"),
		.tx_termination                        ("OCT_100_OHMS"),
		.tx_use_external_termination           ("false"),
		.tx_preemp_pretap                      (0),
		.tx_preemp_pretap_inv                  ("false"),
		.tx_preemp_tap_1                       (0),
		.tx_preemp_tap_2                       (0),
		.tx_preemp_tap_2_inv                   ("false"),
		.tx_vod_selection                      (2),
		.tx_common_mode                        ("0.65V"),
		.rx_pll_lock_speed                     ("AUTO"),
		.rx_common_mode                        ("0.82V"),
		.rx_termination                        ("OCT_100_OHMS"),
		.rx_use_external_termination           ("false"),
		.rx_eq_dc_gain                         (1),
		.rx_eq_ctrl                            (16),
		.mgmt_clk_in_mhz                       (250),
		.embedded_reset                        (0),
		.channel_interface                     (0)
	) oneg_inst (
		.phy_mgmt_clk                (phy_mgmt_clk),         //       phy_mgmt_clk.clk
		.phy_mgmt_clk_reset          (phy_mgmt_clk_reset),   // phy_mgmt_clk_reset.reset
		.phy_mgmt_address            (phy_mgmt_address),     //           phy_mgmt.address
		.phy_mgmt_read               (phy_mgmt_read),        //                   .read
		.phy_mgmt_readdata           (phy_mgmt_readdata),    //                   .readdata
		.phy_mgmt_waitrequest        (phy_mgmt_waitrequest), //                   .waitrequest
		.phy_mgmt_write              (phy_mgmt_write),       //                   .write
		.phy_mgmt_writedata          (phy_mgmt_writedata),   //                   .writedata
		.pll_ref_clk                 (pll_ref_clk),          //        pll_ref_clk.clk
		.tx_serial_data              (tx_serial_data),       //     tx_serial_data.export
		.tx_forceelecidle            (tx_forceelecidle),     //   tx_forceelecidle.export
		.pll_locked                  (pll_locked),           //         pll_locked.export
		.rx_serial_data              (rx_serial_data),       //     rx_serial_data.export
		.rx_runningdisp              (rx_runningdisp),       //     rx_runningdisp.export
		.rx_disperr                  (rx_disperr),           //         rx_disperr.export
		.rx_errdetect                (rx_errdetect),         //       rx_errdetect.export
		.rx_is_lockedtoref           (rx_is_lockedtoref),    //  rx_is_lockedtoref.export
		.rx_is_lockedtodata          (rx_is_lockedtodata),   // rx_is_lockedtodata.export
		.rx_signaldetect             (rx_signaldetect),      //    rx_signaldetect.export
		.rx_patterndetect            (rx_patterndetect),     //   rx_patterndetect.export
		.rx_syncstatus               (rx_syncstatus),        //      rx_syncstatus.export
		.tx_coreclkin                (tx_coreclkin),         //       tx_coreclkin.export
		.rx_coreclkin                (rx_coreclkin),         //       rx_coreclkin.export
		.rx_recovered_clk            (rx_recovered_clk),     //   rx_recovered_clk.export
		.tx_clkout                   (tx_clkout),            //          tx_clkout.export
		.rx_clkout                   (rx_clkout),            //          rx_clkout.export
		.tx_parallel_data            (tx_parallel_data),     //   tx_parallel_data.export
		.tx_datak                    (tx_datak),             //           tx_datak.export
		.rx_parallel_data            (rx_parallel_data),     //   rx_parallel_data.export
		.rx_datak                    (rx_datak),             //           rx_datak.export
		.pll_powerdown               (pll_powerdown),        //      pll_powerdown.export
		.tx_digitalreset             (tx_digitalreset),      //    tx_digitalreset.export
		.tx_analogreset              (tx_analogreset),       //     tx_analogreset.export
		.tx_cal_busy                 (tx_cal_busy),          //        tx_cal_busy.export
		.rx_digitalreset             (rx_digitalreset),      //    rx_digitalreset.export
		.rx_analogreset              (rx_analogreset),       //     rx_analogreset.export
		.rx_cal_busy                 (rx_cal_busy),          //        rx_cal_busy.export
		.reconfig_from_xcvr          (reconfig_from_xcvr),   // reconfig_from_xcvr.reconfig_from_xcvr
		.reconfig_to_xcvr            (reconfig_to_xcvr),     //   reconfig_to_xcvr.reconfig_to_xcvr
		.tx_ready                    (),                     //        (terminated)
		.rx_ready                    (),                     //        (terminated)
		.tx_bitslipboundaryselect    (5'b00000),             //        (terminated)
		.rx_enabyteord               (1'b0),                 //        (terminated)
		.rx_bitslip                  (1'b0),                 //        (terminated)
		.rx_rmfifodatainserted       (),                     //        (terminated)
		.rx_rmfifodatadeleted        (),                     //        (terminated)
		.rx_rlv                      (),                     //        (terminated)
		.rx_byteordflag              (),                     //        (terminated)
		.rx_bitslipboundaryselectout (),                     //        (terminated)
		.tx_dispval                  (1'b0),                 //        (terminated)
		.tx_forcedisp                (1'b0)                  //        (terminated)
	);

endmodule
// Retrieval info: <?xml version="1.0"?>
//<!--
//	Generated by Altera MegaWizard Launcher Utility version 1.0
//	************************************************************
//	THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
//	************************************************************
//	Copyright (C) 1991-2012 Altera Corporation
//	Any megafunction design, and related net list (encrypted or decrypted),
//	support information, device programming or simulation file, and any other
//	associated documentation or information provided by Altera or a partner
//	under Altera's Megafunction Partnership Program may be used only to
//	program PLD devices (but not masked PLD devices) from Altera.  Any other
//	use of such megafunction design, net list, support information, device
//	programming or simulation file, or any other related documentation or
//	information is prohibited for any other purpose, including, but not
//	limited to modification, reverse engineering, de-compiling, or use with
//	any other silicon devices, unless such use is explicitly licensed under
//	a separate agreement with Altera or a megafunction partner.  Title to
//	the intellectual property, including patents, copyrights, trademarks,
//	trade secrets, or maskworks, embodied in any such megafunction design,
//	net list, support information, device programming or simulation file, or
//	any other related documentation or information provided by Altera or a
//	megafunction partner, remains with Altera, the megafunction partner, or
//	their respective licensors.  No other licenses, including any licenses
//	needed under any third party's intellectual property, are provided herein.
//-->
// Retrieval info: <instance entity-name="altera_xcvr_custom_phy" version="12.1" >
// Retrieval info: 	<generic name="device_family" value="Stratix V" />
// Retrieval info: 	<generic name="gui_parameter_rules" value="GIGE" />
// Retrieval info: 	<generic name="operation_mode" value="Duplex" />
// Retrieval info: 	<generic name="lanes" value="1" />
// Retrieval info: 	<generic name="gui_bonding_enable" value="false" />
// Retrieval info: 	<generic name="gui_bonded_mode" value="xN" />
// Retrieval info: 	<generic name="gui_pma_bonding_mode" value="x1" />
// Retrieval info: 	<generic name="gui_deser_factor" value="8" />
// Retrieval info: 	<generic name="gui_pcs_pma_width" value="PARAM_DEFAULT" />
// Retrieval info: 	<generic name="gui_pll_type" value="CMU" />
// Retrieval info: 	<generic name="data_rate" value="1250 Mbps" />
// Retrieval info: 	<generic name="gui_base_data_rate" value="1250 Mbps" />
// Retrieval info: 	<generic name="gui_pll_refclk_freq" value="125.0 MHz" />
// Retrieval info: 	<generic name="gui_tx_bitslip_enable" value="false" />
// Retrieval info: 	<generic name="gui_rx_use_coreclk" value="true" />
// Retrieval info: 	<generic name="gui_tx_use_coreclk" value="true" />
// Retrieval info: 	<generic name="gui_rx_use_recovered_clk" value="true" />
// Retrieval info: 	<generic name="gui_use_status" value="true" />
// Retrieval info: 	<generic name="gui_use_8b10b" value="true" />
// Retrieval info: 	<generic name="gui_use_8b10b_manual_control" value="false" />
// Retrieval info: 	<generic name="gui_use_8b10b_status" value="true" />
// Retrieval info: 	<generic name="word_aligner_mode" value="sync_state_machine" />
// Retrieval info: 	<generic name="word_aligner_state_machine_datacnt" value="1" />
// Retrieval info: 	<generic name="word_aligner_state_machine_errcnt" value="1" />
// Retrieval info: 	<generic name="word_aligner_state_machine_patterncnt" value="10" />
// Retrieval info: 	<generic name="gui_use_wa_status" value="true" />
// Retrieval info: 	<generic name="word_aligner_pattern_length" value="10" />
// Retrieval info: 	<generic name="word_align_pattern" value="0110111100" />
// Retrieval info: 	<generic name="gui_enable_run_length" value="false" />
// Retrieval info: 	<generic name="run_length_violation_checking" value="40" />
// Retrieval info: 	<generic name="use_rate_match_fifo" value="0" />
// Retrieval info: 	<generic name="rate_match_pattern1" value="11010000111010000011" />
// Retrieval info: 	<generic name="rate_match_pattern2" value="00101111000101111100" />
// Retrieval info: 	<generic name="gui_use_rmfifo_status" value="false" />
// Retrieval info: 	<generic name="gui_use_byte_order_block" value="false" />
// Retrieval info: 	<generic name="gui_byte_order_pld_ctrl_enable" value="false" />
// Retrieval info: 	<generic name="byte_order_pattern" value="111111011" />
// Retrieval info: 	<generic name="byte_order_pad_pattern" value="000000000" />
// Retrieval info: 	<generic name="use_double_data_mode" value="DEPRECATED" />
// Retrieval info: 	<generic name="coreclk_0ppm_enable" value="false" />
// Retrieval info: 	<generic name="gxb_analog_power" value="AUTO" />
// Retrieval info: 	<generic name="pll_lock_speed" value="AUTO" />
// Retrieval info: 	<generic name="tx_analog_power" value="AUTO" />
// Retrieval info: 	<generic name="tx_slew_rate" value="OFF" />
// Retrieval info: 	<generic name="tx_termination" value="OCT_100_OHMS" />
// Retrieval info: 	<generic name="tx_use_external_termination" value="false" />
// Retrieval info: 	<generic name="tx_preemp_pretap" value="0" />
// Retrieval info: 	<generic name="gui_tx_preemp_pretap_inv" value="false" />
// Retrieval info: 	<generic name="tx_preemp_tap_1" value="0" />
// Retrieval info: 	<generic name="tx_preemp_tap_2" value="0" />
// Retrieval info: 	<generic name="gui_tx_preemp_tap_2_inv" value="false" />
// Retrieval info: 	<generic name="tx_vod_selection" value="2" />
// Retrieval info: 	<generic name="tx_common_mode" value="0.65V" />
// Retrieval info: 	<generic name="rx_pll_lock_speed" value="AUTO" />
// Retrieval info: 	<generic name="rx_common_mode" value="0.82V" />
// Retrieval info: 	<generic name="rx_termination" value="OCT_100_OHMS" />
// Retrieval info: 	<generic name="rx_use_external_termination" value="false" />
// Retrieval info: 	<generic name="rx_eq_dc_gain" value="1" />
// Retrieval info: 	<generic name="rx_eq_ctrl" value="16" />
// Retrieval info: 	<generic name="gui_pll_reconfig_enable_pll_reconfig" value="false" />
// Retrieval info: 	<generic name="gui_pll_reconfig_pll_count" value="2" />
// Retrieval info: 	<generic name="gui_pll_reconfig_refclk_count" value="2" />
// Retrieval info: 	<generic name="gui_pll_reconfig_main_pll_index" value="0" />
// Retrieval info: 	<generic name="gui_pll_reconfig_cdr_pll_refclk_sel" value="0" />
// Retrieval info: 	<generic name="gui_pll_reconfig_pll0_pll_type" value="CMU" />
// Retrieval info: 	<generic name="gui_pll_reconfig_pll0_data_rate" value="0 Mbps" />
// Retrieval info: 	<generic name="gui_pll_reconfig_pll0_refclk_freq" value="0 MHz" />
// Retrieval info: 	<generic name="gui_pll_reconfig_pll0_refclk_sel" value="0" />
// Retrieval info: 	<generic name="gui_pll_reconfig_pll1_pll_type" value="CMU" />
// Retrieval info: 	<generic name="gui_pll_reconfig_pll1_data_rate" value="1000 Mbps" />
// Retrieval info: 	<generic name="gui_pll_reconfig_pll1_refclk_freq" value="125.0 MHz" />
// Retrieval info: 	<generic name="gui_pll_reconfig_pll1_refclk_sel" value="1" />
// Retrieval info: 	<generic name="gui_pll_reconfig_pll2_pll_type" value="CMU" />
// Retrieval info: 	<generic name="gui_pll_reconfig_pll2_data_rate" value="0 Mbps" />
// Retrieval info: 	<generic name="gui_pll_reconfig_pll2_refclk_freq" value="0 MHz" />
// Retrieval info: 	<generic name="gui_pll_reconfig_pll2_refclk_sel" value="0" />
// Retrieval info: 	<generic name="gui_pll_reconfig_pll3_pll_type" value="CMU" />
// Retrieval info: 	<generic name="gui_pll_reconfig_pll3_data_rate" value="0 Mbps" />
// Retrieval info: 	<generic name="gui_pll_reconfig_pll3_refclk_freq" value="0 MHz" />
// Retrieval info: 	<generic name="gui_pll_reconfig_pll3_refclk_sel" value="0" />
// Retrieval info: 	<generic name="gui_mgmt_clk_in_hz" value="250000000" />
// Retrieval info: 	<generic name="gui_split_interfaces" value="0" />
// Retrieval info: 	<generic name="gui_embedded_reset" value="0" />
// Retrieval info: 	<generic name="channel_interface" value="0" />
// Retrieval info: 	<generic name="AUTO_PHY_MGMT_CLK_CLOCK_RATE" value="-1" />
// Retrieval info: 	<generic name="AUTO_PLL_REF_CLK_CLOCK_RATE" value="-1" />
// Retrieval info: </instance>
// IPFS_FILES : oneg.vo
// RELATED_FILES: oneg.v, altera_xcvr_functions.sv, altera_xcvr_custom.sv, sv_xcvr_custom_nr.sv, sv_xcvr_custom_native.sv, alt_xcvr_resync.sv, alt_xcvr_csr_common_h.sv, alt_xcvr_csr_common.sv, alt_xcvr_csr_pcs8g_h.sv, alt_xcvr_csr_pcs8g.sv, alt_xcvr_csr_selector.sv, alt_xcvr_mgmt2dec.sv, altera_wait_generate.v, sv_pcs.sv, sv_pcs_ch.sv, sv_pma.sv, sv_reconfig_bundle_to_xcvr.sv, sv_reconfig_bundle_to_ip.sv, sv_reconfig_bundle_merger.sv, sv_rx_pma.sv, sv_tx_pma.sv, sv_tx_pma_ch.sv, sv_xcvr_h.sv, sv_xcvr_avmm_csr.sv, sv_xcvr_avmm_dcd.sv, sv_xcvr_avmm.sv, sv_xcvr_data_adapter.sv, sv_xcvr_native.sv, sv_xcvr_plls.sv, stratixv_hssi_10g_rx_pcs_rbc.sv, stratixv_hssi_10g_tx_pcs_rbc.sv, stratixv_hssi_8g_rx_pcs_rbc.sv, stratixv_hssi_8g_tx_pcs_rbc.sv, stratixv_hssi_8g_pcs_aggregate_rbc.sv, stratixv_hssi_common_pcs_pma_interface_rbc.sv, stratixv_hssi_common_pld_pcs_interface_rbc.sv, stratixv_hssi_pipe_gen1_2_rbc.sv, stratixv_hssi_pipe_gen3_rbc.sv, stratixv_hssi_rx_pcs_pma_interface_rbc.sv, stratixv_hssi_rx_pld_pcs_interface_rbc.sv, stratixv_hssi_tx_pcs_pma_interface_rbc.sv, stratixv_hssi_tx_pld_pcs_interface_rbc.sv, altera_xcvr_reset_control.sv, alt_xcvr_reset_counter.sv, alt_xcvr_arbiter.sv, alt_xcvr_m2s.sv
