// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:28 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
p4UGa7ECECzE3zDgKSqLOsM+mnu2oEmgG2EZwY5bKSyPieDEP0z725tkrtOeiV4a
OeqineN1L2kg2Lrq6BqwiYZWtAxGlEbcOGvESuvXMGNXzGxtnpAojvij/jBpbF4t
hqJXEMyeaLJ+o8zsWsikYapuWJY0wpmnAyJ9iURito4=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5680)
IvLvhpJjfR0HqwqDsxNQGawGBtLdSqEV1EerHgZHR7CX/TzSi8MQpMvavlj7Vpr+
FcuZXA0tqwz9BZj3DTd+U1GapJ/7uArvl1NIlsZh5souMZWMD4KI4S0FQVcfzTIG
3YX+sFS3D2rAo9dZdgNxzzYxugoT8lGFuLPfpGkSi5kdtbVQOL9tMr9f/LiNL7zn
ApS/T+/sSLQpQrq/3PZpMWKBb8d/ogUOF8bcHR0uWuJmwi/GKuAfoyzTqVUjdX77
dmZu2Wej7phjy8MkaHzKeD+jcl3O9llSjaVhnrotyccsP/Qro9sePTUXclqY4Sw4
horyBamsaqm57v2sXLWtiSc8H064YeAitZ2h/f0VhakMyQcsKexN/dIQhNEnJK6K
Aym61vlqY9rQzH7X8GLeErBOozl0CZl+tTB56FniXpwOPMJihEPjB05uNwk1M1la
YmdG3HptudA6EO4q6ZlqB/mlN/QSCs5m3PK19NW0YrNsDpQO+xRg+DgaYMKKFQGl
c1eAEKx0fD9LRVEdeDAMdOKTIYAbeGcZz37XQchLuKB7se2Rp5hsM3AYXp4Gi2Fm
2JSdgOHna1PSpNCO9NnuNba4LA6hWMf2RkanC5AWd0dyMByWDWPfyhFc3lrzMLu2
xbAgh2OSXNQiK7mPVPPW5f+jGM1utU08cwNdAmXNp1oXA3PcaBpH+e4e/j0BWL4g
gZxrsdNpxP66MCpS+RNEPzPJvles+WE/0vq6DBNEKF6YtWCxcYsG+qCJgD61oSnR
2j9bZYSm1azcZB92tbnVaf2rllxkx1i91HU1OP5jUOdajwIQTNyzrA8ybONr+Y91
zOQfx3lmVcx5KQkIuugvy0MzqGIWE4TqiZzv7/v3mIL1XHtPvlINdEuVgWjrK9+r
j3zjTdFvK+LItj97QmBrDL5tbrCM88c5Od+vSTzLi6guEaL31feeE98JwhumyK5s
wist3e7NNKLGZ7WPVZc8PZS0wT/jiRuYNfAOQjP8vlJMbPVnmPp70+j9blnrl/D6
SsdGe3qegP1Us08ouXXhoNWlJcz83Ru6/gPg6SfIiT1TqQPYwK6ZfUujZfGOCOiI
lq9ruqh6mr8a/WLAJTKHCP6wH4oADQrHNUnsWoRJbyDE9HXq+28l6AviAzYopUIW
66TsR0X/KFlk9FwN3gtdreMc6Da2+J+SyoBTz2bQDVOpSKgUk4+IqgH2gI9lc7/0
ETXAhz1l3W5XtqeQknz/VfspDpBGJbjKMjQR4EwxyK4LcocYtacJAZwufMzDXcjl
6qLtSaKiwQTuT64AYVWxZaujOOrjVGa8Fsijco6qF3fqDU7vpt+A76mS5NWama6i
TANAUNM+C5Lng3HDkHudFZi+ScNe9tM6zEUafAvHrmd8EXP1SZgGQzaMT2eVGV1X
ihp4kt8upbLFrD+346UO0S2Yl4mDelIHUWgAgPE1HTnI/oMlmWnyLtrAWnB9xqZc
cMQkEIEOPneibGRDcwFRgDV1R/XorwtglJhAsJZlJzNuFCHncB//iO1y0RyVgX2O
LeuqI4jAjg7mJZnoOniEjEKPuNaLf5r/99Zuk6Eo6u6ttitWeKr8ZwVNU5XGGAwx
LnJkNbVYtCqqM/2wYO5M6tJgrxy1ZTdVeOuZ38j43FJDWC0q1F+BUwOuoLrMQz6s
pEBJeYqV4x+/Spfbs688LrVOF7j5LD6+dPBF31KZaZcRbI69dhb7AbYgwjhON8ne
MipN6udUSFJszHiLtBMN8nReVrf0YBhzF6UOOwWkP8w00aT0jJi6LNrRGXHXD8Eg
ZDfLWVVaoc6ALcySoFRenB1LDXY1f5F9BJXsobCBi5JV1rAvnxzU6bR/T2R7xkzv
464mkrLEhjHN2CxvniVaep7keHuPGk7I01ih2dwBAJ1HA+t8JSjDn+8kGVlBHfkq
uEcbUNRIL3QnYFb1YX/dEqRnkbKiAz+pzSozy+kokAiVCirMoFXy9e4nCu6qgbfk
nZmQiFZDSryYceaLgqYZYk5MdJ9VAPm7qtcnw+Z0arOXk/3YD7zdjhQ8kTeT5wHa
PsLN/bXdqSVAT5GtoVbReA5tvR24sd2MGHu2441wK6g3zVtykEU+FB3P1Ep7RLoq
pguf6jDh8nFDDFwn5GALEuCPHmdFJQJZ8hcciw9GgqT/OLTT4rZqUMD7lbNZyyTa
1sI4rBVWK8ogsHcCpIBIWwzjbrv2i9cAvCcKK7mqs102gC4gqCsBGK1e3LT9KJd2
0oQvdoGgpB1QgoPxe8KB/p0+n8UNDL0cKzGGmKSSWZpSZxYPtJeqkKxeThLzrLGd
PoHWImYMjLJB5JxINfJdwnOhgRhcRDQxweJ5PK/lraEZojqaY0fdfNIf60r6GmBN
Fzo6H6cKe5Kw22t8Lc6EVl0prGkatCZNGhMOWee/bBIubApjJBF/evJgC6oExNg4
Pvy6BUmeWgIlloPv4jYTd1g9ZCcmzZld8IX0zWpP71zTBp/xVPPxRMjfUCZTPlZh
ScUYHm+62p8gfDasjXEwNjtoMe28ty4TFryirBuQ+zZWjOd6M0kqMS02qgxP9QeL
RdPbmXUoG0YafMVS5qKfJiRzmMlRlx7xmL+P/8IA/rKvZYTEyMwS6ClsX7ZF4KF6
ErNi0BnMrVeAUD5zmiHCRekjRIOVcEcUz2CYYHyj429Se5rsWv6mKZQj6Gs9scTu
eKft6a0FBg5/oTgk78z0QRU0zVd/Uhw8mIyMDR6FhYFD1EDJNUBe1hvLJ47KjvmY
WLjNGU+J6J367Z/Wt7X9oGP5pBNAUuwROhuGUNbqPUHJ3ohfOI0wE33RaOfhxCBa
YGO0uco8sIppEHDes8jBlOO4h2k1KZh+JxfcEsYUf7TvOpay06s5S+tXnNa6YvgM
Yp/rDzub0lmphkphrESISExrkUhV7UCJ27x2+reUP8DD7FC1Q8jqmU0pD5Oa68tJ
4tnsnsY6eyD9BzrCMjuN1hBFWHDn8SHgxPndyx6bFfHW0yciWIQz3e7d8wHULEwj
+6Jw6/8891AHi+lsAw+ilbOVCtEb2MUwRtfDNUnU/NKFAu0ACjB5TM2Xkb+b2ZuR
TLwmZEAUG4hfJLcQeWKb1lHP7CFOvEZ9gziPll4PxaEnonRZ3fNmHNBEDw/RXCqx
43qznJjskytYCmcDgP0w42I7BfQqqDILgMkq1FgjRC5R22eFuNEssHR1aNeim+MD
PXHV4xEit++uGU6jfPw9Nn6JLY85Qip+ZsjYzFvEXELe/Uo4fbNJiTSqSqVy4FDM
buKcD2TD3grMXrYfrW4qA9h01gr06wP2TD5enXDWdxi3DaCWj8QAKDR5XouT3dsc
u/7i401x6sKDtMwDBi/ihp7cO1QLkELu5HUTfNtxRb45GLMYYCRaPZMegQgmxFme
kYh3P2HmO4soIrIoU9dTX4wsRmncwvK9O28h8avysi6BpvXkDf9YTZm6E0IpANFp
VcMjKKiohx8i+NJ5EeXE6K+KBH8kvXKioALE8ZiyYjiXPqSJhWeORHjqFPJgs1N7
Bu1uulhbuQas5dizJgMIQD9bgRq9d2K1u2sgIsGjP+oXEppmiooFxl4fMb4fiALJ
ef4jjSskclh4o8qITkMGeo8p6kMQ/D88OfsCOZo4OwifazigA/iznEoQtA6phlUg
Zpyk+bQCeYaD08PsxKMUZBxQT8/WwmjGOols9vAUS9+tRA/SS/Opc6cApBvU0zOb
7rrQ4oPeWR0RbM7L4dsiXPD6uCsld5v5fD7AMwWVyceGbvFC/h1kSvmLQQlL0RCo
ZnPpbYM17ZFx9vHOtD9X2ncnxx2wGvwpWZ9i9G6pT3Brlu1NvVjBOKNFHD/c6w1W
cjhKs5AlYzCjjrZDRt8dAUxDMv2wjJGD62fMIG0l82Wx3418za21th4KEF/KSeSB
2vlPw3mVFxU25ykh7gwDS0XTBUEQhx0+MBPngHilG5Z6VvtmUKeDhqyFuQkiZ/XI
g+wCr5NZgDkflwVeqqKhJg89HN9DraeezbYqMahI9yw6K9LTHDXb+yGM9KqGmULY
Jt/C/Oe80uJCl2EyMz1alGcZZJgp1XDmB2EQF6KLs7m9uStww7fw41zRWjmqcROi
Mr2ucl0vv59DuCKQPhUWCPAlpQdDqbMxwdCnCGrIBN5IMuu7w4XbcnRjsfLHEVQ3
PrcvPgrwtybTpknuMJPlkYHlVQ3WWFjkuDgy84T9e02CKYwQy5TctXvlPfLBFDEt
LAMTa3s6znykkIgTMeKtwu2rLG26x1LVHRJ2nhKzvcH9uY9RlvQtRXR980SRfUFP
XPAy/nB8XTD1J+NYsE7g852dX+8CoLqFwQ7DYEM5LbIo5q28wwn7akX45xyWj11E
BDtgVJVw7+zec6BECvLugY0fsEsDCIWnzzE/Ul6EoeEtHmy1/k1vHYdc7eRikoCS
PkShtintmSe2eFm5upJL/0b7KTBt5yi8fotVsna1cuqrP9CqmgK7JbRqjFRYc287
O9PzGlDBrIz9HJuv0rs08AHijyB3Iq1taPONP/FLS6oDlfbu20HPCoA/1+To2aby
lggqZ06h3o88ZsOycjtHvc5jvP09SSBz0xrXiqgcS8w68+3uvHKm04/db+vhnQEN
KtvXH1+VX365HeQ5whfudcTtS8VTaGJjmr8ki4O6n7arYW0f2FaPYSZLfzK+n2ny
njwt6TZ1m0z4bpel//z5mnAYwfvt4zDjzoETZrG5kJ8SbKCern8Bxu0cZzA+stjW
KlRm9lIAX5j2lIlYjVEY6NI7LWZEefZMpKRixCQCG9rJH1XGYpCkJBYT/lWyYKlP
O/+9kZtx4jeS1r/LTg581bqwxc45jmYwr4dVzYKNXanOEey416/6lxvzoJyDnfHi
N97381PsXcnYM6NhkbX9LvH7bGK/qDQHSnk8S6kyNNl3gyVPQAJjO/2oDtSn11BM
26nr8+dSEiHiEKMbfpFhntlFsiO08+ChqQJx+jCOaJv7nyvujzYIQ55i5U2IU8LI
ystG7kQlg8Rwd308ongRAro024n3V5MHh6aAqvGdKcDvNjNZv0/iMaqJ51zuV2VM
7UkqVa89Y/GeJdnw4/dM350J7Ba7Y7GvEckq9BJaslUH6JiMPRWcQFw2lmG03NwZ
KmMmv3Tg5kBK6HkMsQf4ZmLpimI1qzsUzWnqbDslK+ta0N6Z89ZNqEKgLOZ/hNRI
PgkqFOkuH98Fn+loxrIXvdyn/qCftew5FR0aeKYTVMprHwPjmYcfdWvQxxKia8Vv
EZiyUanqVamSrz7x/sXTGjNkmNGr696LDzF2Ob8lsPopK7xTY3KAAvhRgheWA5oe
CTjjocj58T+bgjJqfunrOj2C5RL7Qv5ghvaGsb7WyXhfap2weRjzMqmXUURd4Z67
uzaKXrCyYlYq0CLbkcNjAuLYMk74pgXV35UHLch7hefiRBpaL2WLFNgUVWVxwhc7
Y1l7M4IXwrSXLF1vEALXkxm2FE6Dbc3UFGv66rUY1IMW+BBL14sj1Lt6tN9BC50D
wSARFaYUk993lGqH9n2JhaDtbjTtNVfGWIsoAriAgdyVg2eJShdRFepaVEl9C6h0
fVRpND6inG+l7dKtzSOQkLygQYqlh+VtbUMc+uymGF6qbsokVsaX0sH+HGmzEJ7L
09dVaQ+gxueKou9I0oVWWN4UwN937WwH63eiD30cOXaWmQrpdImaE3kqZMSb+IZ7
f1kxh+ATglLaFIhEX22lb0EU3D9Q9kyHlOVGN2uPQJrC+m3PNrAkDlmLMmNFuZo8
aUJxpvAR6n/ru8hwX4ziE2Gf0dY8iZyCXy4Gljs5zJAJSwQ06nX8RXMhVpW9KrMM
YirhwvLG7u9L8g3C2rEy+WAmw047Ib6c+hJs8ikKHteh1fsITrznGUxoWPpNKIuo
zNhT9D47QB0xNslgZ4R7ZtgMk9/h/BKaT8+xdaIYxJJIQrXJ3oZS/JjNxgsGbOto
TB05Uv1G99G9UztcweoFPi/wQZ5PX40PRxHhPsUqyqQB9iQ4zx3vxhyIc0WzPGy/
/Kx7d0VrDlF+4vBvFGgXe19tWozr7SSUoteGZ0qzzD9g62lNhaTkE6k1lmZ429Ji
M0+vgmIUxlMs7qjR6W/nxb5cU2asOPN4XgWlG/9Xx/JbZNdpyIrRj5wtxijDNuG9
6wpJ59qCTPdvPov1Cyiyj2/BjFyIhhzQAXDJXVU+8liae4GJwNRt5zXmCHLX4ErA
Dfvn35ZoMcosAj/Pr0m2RzfUCG7c5YgBsasVwYgsAk8+YC8VpF6ZCmDrzuIkj1Ps
KOY1JPqPd0oCIzIcAhNXcNkpnh+T3pZFHi/Xguhtc9lsOGxeYx55UVLkSl1kbuA3
n5AsgG/l23d0H+rHwVw5FEVwV4NtPeXkWY1ursh5HzUKdJ73KtNnzeEOkp5Rt1dd
YyLhtFwydnqDYtvcxoaJ6IpfZ32dVqF8O8AUa55gJITxS6sxI3Sfr+TEtRduli6p
NIGzQH/4cPZAkZSfAdgzlhpEY1d54x4oB9aye/eug+jcUvIRZsi9KXcw7EVNRdNN
Vm3yLOECwX8yfQGRi+Rt/rCVc3sCP3jjcRtGDxKIosb05Y9N79dbnQy0zlWe7cX9
VOKaPsvxMe/yAeuA1t9fqKZeOaOdFTzxzdezjamAjuWWXDA6GprYRv8TF5NUayxD
z5lQ4A49crlH1LtWX9j9P0Olmdxfvv+iXUK5HlYW5DOTVpOs9mKFYz4QuB9ZE7pS
cDHfgWev/mN89Pr5SiwXvXu2vg8tOSNxVvjddtl5UbdM7gg5kGPujGSp4rdnQ5hR
dM7ByeNdfZQSyaDuFQpFKnN5ZdgSYOHlkfYENo3Xy2nfWYajr9ekzBMeSnxMqXC+
oaeQQI5drUKDj3BtjEkEsdl+Z1y360bugQ8zn8u0Fg/SM3DsvdaOeRQkbowMzIeQ
t7mc4zzOy+D43yN8JFK5mrC1AyAJVwTSQ9zz+t9ksYezMTDqVVzHdGPUbZdAZJIx
ZpWQsVbsY/imeIg5ICu8arhNdpoQ8OuL7GIVEdzMzZococXZ8UYvaG9TzxybQXS4
Cf3cf1lGiHpORKUcVkOMsFGU/mxsv/sEZJuQ5Z76nA4ynRdlkJJlPjdOgwxnF+HC
drqvtugFYozcoTnnfP70vRbYKpeEmuFJ4HP3hGGJW3LwtHSdL7V28r625CHEjJan
19lvyj+fva2xirV5r23fQ0cJ4Etjqxaq3MJoTtwc/nt8ObXJ7ecdXxP9hFAA0frd
Tc72V9h6VaKgZio6GvMESv54/Hl7ykKxKBDoh8/dsmQvWr1Trq1DhnBg6gXIAY/X
tlsZCbplTRbp3x4wmdlvYMhyB1tGOluSvDh42QSNJT6sT6Af1L6vgSCagHULLw9D
p+RL0+LNwaInDOc6cSQrRV8eGZ2uofln51RuqKWgEBhR+qDpSFR8DYxfNPfaDVMS
Zg/xofa8RDgQmZcAFjRZDbCFhMJEl5yc0nz9wWipjssaP/EJVqADC9q/u6NMtBmJ
+Fy9rlGyE7zlUxZzMVHy14SdnNbo5ji2eNah0PwKcu86OlT7ih+KkPnzZsE1ft52
lL28R2hXoFY2I5xwYIpwfw==
`pragma protect end_protected
