// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
oBD+PCQJJ9F0Dvs3smwvqYmoJ/nLDOGRuLrKR6k16DtKHii93PPORlZi8LVUaDYx+vLLyav7RpQp
b4r7QV2URTGbGb2IBtBDscQUCzxq3ES0+znwrvqD1wl0pOfNq7b6ph6kUOMiiF8yggj+p16yWr6Q
aZXA3oPYDLh8MIIhehyr+AViJQvM2RiLijukrlE+I9i7yatoq7fumT+N603aA4T7xqzv71mrzsfj
/SNFjcy0nH9JB98DonBN8pb9MjGDOuEU5SrmgBCBe/ADkweW+7IGdJwq+sU0/CAp0jhmH6R90O6F
JPENMcPG9cshLINFjnRZGiydT/exLQ276FwQnw==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
u6MQxOXknHLtBcn9cy+XHFVQDFyBp+6sxt3kpdKGNbrmb1hlK8ilhKkXyqnkangA7w0ZQ4SgssM3
PUSYbR3yApLYIHItiHQeFaxfM2tBK+bUFCxbBCa28c0cfqyfCsybvSo9XNtjFlMlH35wKrrnESIE
bM9AXmbENCROPb/zihuU6gxYKQGdMgQ0OH3jerVH/0OAXK6tsFckw0Iqqj1bumBxWs0X2ZUgDNXP
XB6+GZT+WseFqE7VACLmWvucMRb4zti32BBpH1PXzsRhhO9jXJJva454Eh+hwqJLbOv0Hj3dau/M
D9ePqCAovciJ8KitI17zoDreOqJqgsODbyE+nYu7aUxMr9TYRR7A38cVqFSVcAe26RwlpthYTtix
lsISOEh2rAwGoJKNPZt88mKyUTCg9nSy4q8ivlL8L5ue2QAqSvjD7pzlx3u9E0WFhgisRz7ESUAv
9u7R4Hkh61eJ+d7AKA66hH4BSW3jAl2RSq10+AUVjAosMjHfNhsTesBSoFF4U52ZdCRJkx5EaKL6
6uSTFy5kTq3OfzYOw0jHDFE44gL1948mR3zCydJqTfGNFQjQ1MLEEr0A+Cd92BmBfterCZ7xmfnM
c1uwqrMdZ75ybJ9PbC+QjKmc0Xbu64dJm4TCeTqbl6L4aIDI3i0Q5eo6IdmCAJy4YRwzqnC9RrlZ
hhhFOmZt1Lw+Z/fgjkpD8iyeD1YsF3E5xmWa/BRdHUDfRGEAfHsA658hzdWY/Q03pmB/7Ns6/L+f
Qe+4g6rv7vh/RUSb7vXVAeQTvIbTOBaZ77fK+TpP6kop/5XyegnnsRRy+BmU9LCe8JsRleOHBGps
thQNmt8xPRLbjq2c3aKCblEhgPSV2qhR5f59l1snNjcRxuz5ECQPrqB9drKkiyaC3QRE/zLYF2Ni
UG/OBQbkobtgi4HC7uBvZfalBEPHWZedqS8BNwhcRxT0GwcYzIeu7tl0bWjIy+TqzRwYEvgRi37m
qcX0lYARW/WLWHRGm2xZ+yJB2qDcnf2tvwyqjg1sOvGO+x+jP50EX1L6G4ieGxhIbICxKvhjsn+H
1r0bNSt6EZ4O1Q2XzCGZrXf1kgKAyu00FevUQOaeKeyVicmP7QM72wrjshz6oAbQHPg1K5Jl/iBX
kopIJ4uPwgNaN+gYguFlxaDKUyK+9pSgQgGLtLOAoi+CGSFWB+6JxSEdD7UDmgNivdcPCwypRLiL
hd2kYeHBAUXb/ZqfA4OKBscJnTM4synwcQ/ySRyiDXfPLKKDGr8JSDn1fYK2SGAWU1OxbbNLDKL2
2pDYEox8VRdiIQkpb5/vJhfglxUtmcrpulGOjXdICscPcEigi2p2/8ePWuGl9pqEsrkrwvXl3Dp1
oUDI4qyRX5FEtXMg2CL/qDeLXbcK/+OsqgrHT+LNkn7X0rUoZWtpT7vsSpX+8JTAmZXf+Casc0ZQ
eeHmyIRKVKL3KtJIwYCG6oHSjWvk7QoeZY8wirZwlH6nUvVlhYlLj4AYhx/Sa2/ctFjli0acEi/e
uS+4pSedeqE1qbV8l3kobnILMI9V34j0Fy/h8wew55pzZTxaOY+21Y6c74Clrj89PYXJwDg8NmFb
8d8VLUfYTS+I3sJYpW1IYIJIeurgk+XM0TOI7ydjp6FirTRZ4BPV/tyRlQ8lmhiVqlvPtRphRfs5
Yodwl5e2D6IBQzGu17V7Vps1VVuRE81KjWRZJDM7gmHuXx6u+J0YilvcirrgcWO3DxpvH5Y5eLsz
Ml4OMLzZQXrHmNo1LRQm+5qTjKN6W6Qq3NS+OS1B2qAmNDEojgBfX/PvuNvmXVx8TQ2zjpphoGG/
Ik/+7mPKyIP6UAJTeEr3lbYoNWvLw0mrlt0HmzSEIAsdavR9Mz1QZ29ZDK9KIFqpQeJw4d7PNRRK
pacmk1In6vEwDg6QAjUhlR10kcAkHJcMtia9xk0l9+T2jV5N5g85OoHZPGOI36/+x4bY+rAoCIuP
w1SHJcG4EFgTf/mhim8Uu84vyTTEy7mInZdns9fDJGGmx61RjSebmyON5p8RTn7E9jOh7tEVDPrC
ohlbhiJEutkuwh3F2b3NHJNFrsoEB+KLCDx8X6vwL+6zFlUWKu6Fldm2YlprpZbjFzmd7aWlTtH+
SLk8kmDXvq8j4b6z1JE+oVUY+uJa1FZyrywQ/d97WhED/G0AK486y+0YGsPhri6aYctNZzCD4NuU
gqeAbaQBbtfWzIdFP9Z+ncbNbfSTzQyw5WbBY9WDTvIAWe+2ptWQFGv9GiaCTjChCDCaCJekomoo
RqlRJpZZZtfA47vDXIiYrq7CFINasYRCbTCTa9gALunWjJeUfe4rPwncae9cgpMhADunjT6v/jUF
0xVGyX7t9g92609uT9lnbvhktgP9VCQ/zDF6K7DRyQogMeE8m2mHjZSpnIsesWXLo2UDNo5S2jB8
qokbb4jx0qA5+8ncHIhK5vidy6SyDFwjWhnAZvuil1DZkKUwxj9iX/ZfVdvFYLdT8sLX/0FtOvbN
VeZeCospCOrMzaHuGnvcD25HtlqNmVZ9MQU2p3O5YRb9TK6og28q+/p133Z6dNiur2RxicF7MFXm
1t35JWk5g9toOtEdSvzrWc1t52GcXoYRZCtfr6b3yC6W5CN3TmSQ5Z8B0cNx6xznadwW8i2PEPuO
Tbt72ffUhSjYcCuZGHZzqFC0e1KSGTPcaLitN2vmdZEfZVyE4Z9fruA/DPVXG7uM58O/ai01BLzG
Fr45wwUws/WbOunXyrOcnrJegtL6eU65KKTjPFXKPSobkQM1NUHtAH84ByUhg4VqzDNtxIrAfbEQ
jGLrGc0ugQ3U4QyDjswOjHYIEgvP5NC7xCaEd4rvg9dOwV+vJg+sgsgL2dKpR76sXjHZEmTKG+NZ
+1VQcig19CgS9V31NUrTS/Dbm/kxC0dzlORK/b3QFNcZi9bVhboSTkxNM43eTo9yJK3A81Y+FKDd
z8MBTzKbFHBwveum+Kl8vx1doKJrk2hJd2UN8svno5mE/Gx+C2OwMJ9KII4KmeQ49cFWsmf1Abvv
nGip8Lb10FD/amg1BoVhuIhTua7m3vLbL1eYpAfxUJj3izfjayzZkYrf30YGIvsf9DHscoVsg4yz
LgZPIb7Gy/1+0hPAOCOw8FVqr+MNSh26yOUQF7DXYtrm8bwv7sIZxuJTa/nD6ST/l22hMVT9Q/Qm
FZtb0zrNBM7WjoyXNL7wRK8UnEjwCVqDu/wQdvGKsodTtyUOBJUSA0EViYtjMpeP884sPz/U4pk+
+iGavCaHUWCtneuOCaxz27PeB3W0UYFZs+b/Al/Mly7fItlkMYWKd6kQl7TO4FC5T/b0Evce3R9t
ay7m2fHDwpWhLZJ5+T3ICqafJjrqQIfHxUC+/6xwRdhtogQdTwULknrPbso7J/70N8o2R42Xp0VE
ixiZV3t3nAp9Mlp0u5u5SAr/DlZ+rhL/FB9D+a/UQHJ07ZgA5JwVT0u/LMJft6Ju/8wrLi8EbYP7
Y83P4yGeVl+vzEiHE9niMV4zaSDMJay4TUWZXYmGY+Zb/s89z6j559/wsSSFiN8Xy6NoQ5eq62/4
t30bopAsFWM8mUWp/8ZKz89h3NMWckEehRUqVBKICODHram3/FomF1BIuMtdJBWU2Ocf1LaSBsBj
8WmNcrmLwbjip+uLAxEWcOZYENDRZpyZnJfySN7Ss8QOmIQdFepk+liE01YTPBWD6noGp7mCptLU
+4VZX0qTtgnVw1AI5gJLi3K05B/UskRzcyePWTVZCu0XjcKItB//MT+/7os6AmOcQRrfRm5sz9Au
GTLPO/cjYr9G2BCwXD6+eP09n8NdG5I2kGiyikGSXzQFo2X5A92ghyXlwUjoqPzHuPmfygvqxMsx
T5qfBzyDKQ2UEedYCTabAK0xhX/FDrcdZo5y6LVZ9TNY4tNqGpjMJxiJakvLwPcUzoNSdTTCjNFD
NOk+Hf6LF1UDj19YIcLcvYEl/wv7Wm0WlmcFNBbGTlkoe5ey3xpw6h/FJ6M/++eGRpNdCjuU3Kqh
h/3uxaLVKf9OaQW/KWZxyoM1u+yoifoQLGAkYyV5HvpuPAEdhNSWD3HDmREc5+n5hteYP5BL8lMs
RlUTzRgeivY+AYHlpl2pnZp8r0webLKKa9BNhFDxwg1Zou7TY+7WjAsEw2w33CBToub6s6zG6CDu
0hPt2FDAys0U8jtQe7j+8WH/mTrkh6JYm5wq994IEEIlzIEO8JdZG/uUQe9qDJpDHPdncTEeT2zr
JHkn0ioxO1aV8fs4Kzti0gqQU2LMuZYAALbw/OOswVmmNenFMZLu/UvXoJN52D/JVWen8GrGE6EX
f17kaR2DLQIwc0x3WtKxPcYW9Q4cQE3n6ys0GgMhoMknc0fBJQBtWpGv2FtYiqmfifeJ/vKUY3Ur
/PpTfW+DonUskVQaCnzvf45ZcjiLnHRBCLZeCO7/nzBWsDtrtkMCCy50KQFCHKAbIBs3f+S2DuzY
4Kav8t8M8dtYfLX9CRHRouzWgxh0pHvp9+EE/Pxx3WGOUp1UCNfJ0iOthbOICA6i1A9RrX6IKdvS
aGtefHzf1m75lbY97K9338JfoFc0X3PbpJMM3tlNkNbvDT01VDJWfdy85RJ8zR5+IEpooj42ll4b
1KQO+xrKIxRs3i7JejRMlfPPAC4urXi3794MaRP/uJpx+L2MztluKx8dvCnCzU3qESKhSH8Ptz+F
RhIGNbyyKFO36KfRTMVzuJ3UtmDO1hTyPo/sBOiSzIodg/js1sYY2/MSzFHQNb7Y90371nVZLRY1
6aBy7xbgVWEA34+b8avYwK+D3+dYfbgIxVITw3TW6wukHAXcR5KWEwkvFPlseufTnqW3vjU6HnjA
LHerzdLydeRyIpTnD+T5XXtgy8alqOkq/Idihp5WU5WiFDcZcZFzTqn+tmd38mdr3AvXyqih7LKq
PEfN1/fnMuR8ijrmXlD+N5Y8Xt/pYsCc5XqNB6VHzg6P+mEaybrbK+xiHgm7EiIcTF0+1gFcWt5+
2cU4zG2CzI57aEJfbZCmxC+fVCJy2pu4d04YlUp0iGjXUJKBVZtEkvH04242t8W4VI/QYoMCMTHn
Vr8q+BNT8lXgr4BSJn7umBtmEczxb0aM2G6F767GnAQKDN4f5d91Jdr+Z0VXddjCN0tZJ9GXB1uh
W48oXKuUGhK0VQ87LVil/vhUF6HZvdyNyi/ewi8dT/tbScFX8njTTGOr9QL1a7D5Oep88QtUGI1q
Jgb3PnABzW26ogtV7qEf0+Qk8fkBx8vjPMhtBipyuUvxhPpFDUFOn8wUcQrC+52ix71ItT5Dr7xX
s9TphVR02x3ZRGkhXxKxRhUEjmHzAX1X1PKCZwz61mImggW2/i1FosqIgHEj/djNIUgDczXTuvm2
SkMH+lrKZrEXFt+1Oqci2/zO+B1sOyCJcydYo+JwyRTiw65E0en+UCOL5Q8yPs+BDnfHFRhmCzFZ
+SGdQXSx72x8bHptJa4fQkJybmrInkPP+jiek5iNM6U2+q+cedPSEoC0kuUIbtbxwN+XSS/cq11Y
OWonumzP6mrR4aJBsT430/ABpQ/d45ieUaW3HVP5YChczcMOn87WqvYzKaC3cRsZk3ZAK75cs4SF
gZL+4kYGIq3UP0SacICG74IPNqx4Jsuu6RGbstEWkcAI9YMRrayUcG6y73Bh/+4AJfCPRMP6QtI8
AN79sWxwTGUR5A5YKInoj0BMdfmyXG5QykdI6sVA1NHU0ospVmKzJxseiT32f3njZ/gmosL7fIbH
e0mydyL/WYGJiGqzq8hXFgubqzUx7d02FJrWk0X7m9NMlY8Q47abK7GVdjKW+AkAy4Z8D0zjOBKm
xGHrMDCP8yXfCBo7VBBQCa+1hhl7qC+hE6sqC5Hd/4zXRKqreN6xUccJVLPlifX8cl6QZWWO4rm/
URSDFE7Yv5Nw34po5KcQclzG4HepSTo4Qhap1DUNr2jtDzb71Xi4CJHUp9T0FrSB2gLWe0alxxuh
JVbXK78yyDfQkClTpPKfBliKeG6tfXXV4ElmglFusS+tR1vkLvvWYceAwN7dWojV91lRTK8FgVle
pCfGvBoBdkwnmW4l59/46/cNwh3PFXF/EHZb348t/xBPrk/QTZGEOZ7IVmFPM2Xh4LOLG1TX/gDt
nlp2alXL5b45tMnqP2EesDnV8QxBRyc+z/jIsaQbXZeu/Zq+oegmJtSPIIJw9Lxb1b1yf+BAaaU2
f2wzGDahuuBKSB+PCTOjs+vYFv4FTeWl0Jiq44EuKSK3VOKeSPnlzc5se93Y6COLWam99wMZvkns
RqBdGjnJj8Cb9Kn0i7o1JxHAtUxJd6w99FxEfpZSfxjqOJiIYGRhnMACrzZhJt8sXE/2qnYL98Dy
m/wDJ2qSaUjsCHsoX6paVhJdcRx/f13rPmqTf7IxALF/YjRXR+4LpIatpGo8xAVRybKpA3dxys+W
EbQ8lDLuUHEHMAeUQcuyJ0vTVIUQbqN91oqo90dlG4WQJDN14we3JrbHqMJ0cmg6sitQavowWTgn
xhcPka1RZrzDH8TdnfqVGRXxu5j5zKmBGwuA62ls5DwTLyRVZlSCysZOurpMMyWaXqBgRQnSNFKH
UYtTQ+bQvBWPnCn/kO1+KVdZ/6r7fKcIfVz7LjCCWQbXCfkq6654Itl0vYtEj9cy0K7bjKNhbVwf
yFRWuD7397dxvjXvFIt8ujYbXnzmevnKtXkalYRoF0WcvBhMwCy2gBRNC6pFZCCvCh1tXa9+jVEA
P3u/jkWZhgge/QJQE0nUFGSXeO+FVwoHSGhWnKZdGVH8R2+HZZ+Th+t/h+8EPzKjepXn9nCUqxH4
rAT8bvvTZ/gIQIa0rnCi1yfuj8Z/pLP52EWRij45ARJiaTUB4Awfi0Ep7Wn8y8ZPawyxM8feXNJ/
0UllWwo5AC/togrSNN/Rbx2isUE4tFcVseSfi26WktLNU6p5+LjDS9v6LRJpiJtMs4iM9jMvy7kO
HP5CUsOXBI0uuPZ9M5+CnvPUIWFJQHCMV2gu09urQV51BBPbTJ+eGNdMCD+rC8Vp0wrd+wOKZByd
dO+vPB+A4WhgkbKBQqUOL+AH02ucZ9GfhurDtKuBWfgqtlm+tr8IuyNCl4iRMzgYyzz1OGSPPQvd
i+ErOBDaFQmud7hkMhO7MeGc0DfbBarVmzTGQ6H81R5wjhye3VbjpbA+PN1TqSYNnWYks34ejCtb
jbrgo1zO/vha3EKaWhN3pgoVsp5JbcFraqiiCIkHn8m+AU/sssEhzR9VyPvi//6ME6Ij4oC6892R
EGHtMQjHwVictyOK4FYiz0r3vXC8mUmM0q0Wr65Pb8S4mTVClzo8uu0XHK18FB1v97g6sApxDXXJ
S9OROzyphVSwDo+HL5X0fWwrax43api5UuPsq7+I1Np9eaAB8U4zBNl0ztLQ3KgceuKyNaf3G9De
JFkEHnIiw3ijpg7rqhtItzAtCo0UKyfKu3r/x9VZQ88Nl5qkjEkhUVf5tJ2708Y5r/FjAtFuvZSq
EdttqImRXajdihaKN1U2Ach23/7AlGeEWQxx3FJT47FJIncPfH1lyQ89xMI6uVS8UGXD4wCBwE4i
BbX4VBw/vnQZjFwGfOrUuwweJdjrHi5AETHVgBbmuqfGrQQozhGLoVD23/MgzfpbeKgcGL9caPL1
gMzBh2krx+fuFcwqnIkn9/sOgIsPPDXWZkjhdF0OQVrRQMKMLILI76+uE9f38nRnErsChvmhK6Vy
GzOwuW/pZpt2G0zBIhmyT7vwzSXhGBPmxK9+/KxwmyvEZaJaun9UV0I4+Em94Uh5GnPDZ6yOFE6j
u3tzAQdhe3hShqoX33YRU2Zw91O2XHDYQT0J8IhqmMmgFtPDQjGwIP8rMIvn4U8TzcFCxOekVpAD
Jff/HRfv/B8GYploWzDaIATKievtw+9nX+DQnrO3bjx/34KHEjgBHQpkT07mPQvN4DCwg+95xFfs
3MUBVODIFHmtAlp7GTjMt9g3R1i/BHqLYpfAdPtpt13cFcg5ge0Oge9Z8kAqKEFru5Dhi0FcMhuW
teZpVaQAeuXIvvtMXYcdqsm8XUj8m4h6hSv84RN4VbekMwNhLoQ3UgVJTdyY4/SQ6BM4yQFSLYMJ
2oXTgjrs2HeqmcL7skE2Ulp7adFIp5ml0cFqjY4ITll7WvnP4da14TgtmsFGMfAaR68QKrMdaREN
ulT7ze+gNpfZxUYpxtxJDB1u7M4xJ15brsKH7h5Wxn09TPmAdXRbjbCXlfr8+tlOwl5Ayoxw0bVk
aHpoICVSXNNPWskKtMYrTcLmaGW7ECTu5wemjtvzLDa9R1+uLy2TVeTYcxchMwB3nCJfM4SVI6NP
n1c2il3rmIlU3B02AaxvjI/8YXpRWI15RCQwySPmHv85e8/2Ss0ke/rA9FB+qo6eU5XNPRdATeYH
9l0iFaK6DbFJe1WIXkR8ETJdtWT7Q7kyinYLdlSJPhQZ0pzIrQWhCZ6rU3p543oW3cpkwpgyWcZi
M2cE8e47AErl89h2J2oT1P2fvGwJ5KlKtf+2jmrIh4kULQjbLEgVs9t/hbtUmBxBioqEVdW99qP5
7O3hnD8ABHlE89Nf7e7OcATrWLBlI28yByb0EpmKvy2joX0Aqi+hk32s1ngpmeiR3lYQBxIW9a8X
3MWbv/43Sw0W6lXDWnJetiUJUnZK3nYsCl3vyYFDazE2ner4vBKz2Z9ylhej7+Ry04shfdwH/mmY
5lo2vv+TKOYhUiioRXAbypGi+Yacj9MBlJJmQUUk0AGFRBtSPhKczpVMJQfLRGR9G+IhZ+GIlR6W
DpaJuFPbFxX3tLCO8xsX0Og4WRsNJSTw0zGsjeNrG8Hwvrm/yuFAvyh9PJ2rQ2PkZsC0DTn03pKf
//1nicClZKyur/fzTT0A2XxtFCgF7hIt+e3fpzeoick+2F3iQyD1jifbz1T5ys5fSi+Khi0T0j5g
imMYWmWWDqBvG2JsB1HHQz62EkuaOyLZXo9emPf0JOU6pVO3QzQeKIkgOUMG+5VegW78ZDxkfOyb
iMpjocMXi3hOVnEoEtMdtftOzHEsHYCNTi2vqUFAABSRK+Kc2VdQs8fl27PtkdgzGE27CHx9N1N+
eLb4w9xWYugoSPfuSf456tJGNXHN2ajdun9f1keeLFYI6IqZATsq8133VNtMzDLXuqUwavJBFbd1
A2G3OfTnXfnS0eDVgtr2i0jNAPLzKBmCkd/OUuo44dm/To0XJEoqnRhglzVBIjI+G5V4OclGpYYi
pFBgBHU6XZBjeTedlA7ecR6lkPdSZsbdywjiPdK98HyD1DGFV6l3x4+rvf61SBF9lZa6iEhtulpe
Zf4mDN7m1vC9LQAR4SxPQ1fQV5ifsDWYGboBbWivn2Qn5t6Dbrj/6jdy5afrs90lvJf0VBHj2/GK
l/qqLOrm+Pkl7vJ4+OpsmTgOBjdbJeaazk1raj5+JnDCsHF1D1XldjEK7tY1uOYG48e26OKn4YZR
qIy06yTfhA1U7B8FAUfUhPzNjpEhnOm1flZguuIDNPGTwVOHIzcjJ6hejawMz58UQNAXhMdRVG8N
FJ4bRvYsUJMajqkrGnvKAmRyFhrDX8/vsM4Is7znpBwUOpaTjs796jyBfHKaN86C3RRXPgiQuuW6
kAk8LLWOvCzB255LCdcmFpojCsOQZdHrBrHdTzEjo1tF5sJLsQr03mB7ysn3Re/RVlaktz8y0Ifn
A77CyZrWS9ubMNka5JnzaDmo5KtoiYdShSNvnw804keVKVixAJV72Ig2GgKOFJdmCkii1YqFFUSo
FUFnMO+FAIA9AMtsA5GGs1EujIhkhIKXGduSI/L2fanGhjXWkq3yAY7+a2JWdBV0Rl1YbsgMX3BF
CSAr89o7b0QBSI6jGS3mROTNMRFxIcCtKlqQ+DuTynflO1D9BTzT5ZRXCZHSApUWVzsd/YVZ2kbI
y8LlSPB7LnF5l5rdAKD+3dOWhQNWfr7gZq3nhGA2t/TWF59qId1Ppo4OxvnYlXRmpIJDMcvWaqh9
tXr2Z3nPZ0/ImoW2CtpCfutH6IWRdP1Tnn2NVnMUHJr/46cTWHWpwPrAef0nVWyHPAX2GfPsuPI5
4FbIgP4xv//1xAVexPPrwI16iaK9Okz3bb9BteR8duu5VfAT54fW8rD4S+SKkkM+390b8qrrOLvb
qBAC9PKfnjxay84ier3vwZDZZqKoW4TOrJgOzMRV+WvqvuFNiZ7fT16fFjQ/LKaUCLcmhzxP222U
yZaP1YoRgjBweO1wsVPEk9CbLQ+wS+dqve+8iwOOVYxnYRnIMR87L9HodatqkDG2CBKr0LSz360L
dmeoHZ5Pn3hia5cdn7RlAjKf/IxZyNiV9XtXGvxaFuqwQ0cFml9csetO+qDEUSdTqGWxNfXLbcaQ
riDXQQdpRc/9kAbjCJZFx2xounTMH2p9N2Xx32A5SZ39QFHwy7wgsYZTei3hSgl5DB5NIRNcVcQh
O14vqxkBa/MgzEEDe2XK/lh78gNvhbtk+SHcnJKXSFWqgnjWGYIY4QOUA5aaFFRwoSNfiDq7xDF4
qB6HwB2w0lPCHsEkIKz81MG2A0/LA+CtzW5xdDbv5qKYKTC4pB24x46pqpHH+NBu5mVUyGu5G/Fh
3UMXBTUs+cmQ3+85cXZWeyagT4pawY9GExkeKPrzY5bEB3lTmumSsA4ggzECpkW2bmew1lNGe7Td
nm7EzOgFNsI6q+ApfKY3nx75Tc4l6nBB0f0d+j02v2ycqaKrFh4NPfHFP4rtm1yl6Si0I34wbnyO
scMNU1kQhepIlCCfO58y7bPofYf03UqAdtnLHmonA+DJQwkoGLgInSdip88tcPniaHuV2eFuPauX
lCj+muPdH+M3zaq2qL/7FThEb+B4rTg6/XK3+i9yIdO9ZPuooCgzk9dEQc9dExenePpvUBZ2NUqV
u5vYu3tpLrLZ7CDPFGo9fgwADB9KHLT2CjrudgPhnQPy2C8bcNVB7pa81L7h4xsti0BK4nKlBnCd
e7zywklLAZ+wReWd7ozzFY6hug9wIkfXtV63w6TNJ6wHtTzSE34wa24fyIBTXbfYsHtIRA7smqyO
f4VkwtfhuRbuxTIsjYgqsJ+7wr81eCLFNfm2lbaTUVEA/YxS0SYwq5DJGnj+jkfUYLp5iR+IUynd
NcVhTiY92YR31K0QhLt9GLLBdANwoS1lMjWfTvGE9MnugXVRnQgovrqewzLFM5vWfnco3+3DwMgg
4NZJ0mcnfZGqSWpqboo4xlR3Sdl8VwbmP+J4oCojLOtheSN/noIZCu5SdZ79GRdjKz7OxnZxvWAI
In7tgNXzxyCymGx8S28MV33tQ95DvsJlm1FpxT88W3hQ61JzC218T8PCkZc7CgBivg92YhIRm/je
JzHKIyZV7K84XsXx3MQxvI/L6VOnJrqABAGtzr3h++CqJSZbRa9iaXcn7b+rf7AYCrQM6pYSJTi0
/4nX/6C3Br8cLxV5YRlaMHZ9n8W+VowvE5x9OWoC89OSRe05I6T1+Ek1FaF/GPi7OH+mS2lj7n0B
qZieXDwxRvHNSzGp3BXX6wttRuBYjT9Q/59JofAJTpC/2nVW/ZMbOPErX5NwuFLFiRg3cDH2wWAU
+jimwNt0IVouZ7kTLibgLJe+k863j87iRQ/XFDl33aXGY83ZbYMHCb+MHDy5l9mVrtRwRXNb5vU9
nwKvh4xxQlanmam6+ngjpV6UwoZ5tAItINV6Tz73Z2u9bOC4IXGsfSCp+iy1yh6qKP0lmq7R6Pqj
CS/++ASvN89g/xJEuwQcgBfjq6ZDwEMGQijh+DRcGugXZB4LBhu51YmgCWeDSKM83O0cS9O3sQZR
rX4C1xBn+n4PSYWkQQLDWu0u2hxyFA077JZPV5IbQ3qX4qwnRFidm0rVQskEgaeTH+8qOZb7FOcn
B8N/lDYGzg3exNgHWMndQCGXULMvS3j/DxEZUVR3OqA7DnMnGFTEa+56kbx92Suokvxg73f97IPc
e/pQVMo3JfTJg0lt+rvYBo4GzkWg3GwwFL78dKDmlDzMdkrLfHOwrCecCcz14jWiBv2O0EunKEXc
GyGUGJlJ+Hg8PbCWmbkgvDbyrgYdmkMlNSIt2d7K2pTvNf2V7enj9A0gv9H1hRZbrD0UAUVvY7gG
3p1aVMwQAQuhdyOgxdOhrD9A3UWoJQpv1YjcCEYtO/k7JhqwEvjuNdrAZpoj9ZsctQjT+KD+2Ocd
0Div7TrmIdCljOv+bKSO0ujIjqheEuU9TT04xRW/KXmMN3PRfGpHPlfPfT4E3ey26ZQOCIrMXkTN
tEDqV5ujXgSxeAFKfvY2ALdbYFG0sST6F/KGYfqYombu0bSBncAEHOMus1lJyucC08PPwtY9A5Ex
TuKh6HZ0QUm9KqEZPnBUP0AxlDgV3uA0nRjkVYK/SGG04saDQXn4WS980pfXl1STLKiU4f+iPfGY
7BjMWuF+e5O20y+OVxghte8Arfvft0uW69gd2LB75SCaMCj/AIZMgtK3gPA1MxxdciIFf4MYJDL+
QTCixkQhPgSOTsbWb0sM/CaHWf2o6QWsvkbQa7KPHdwdZE8Q8jtDkQvDbCHNsjJ3BDbdGeWJHWE0
761QTMkJ+FxQ/U1A/wcFcgRVIwE9ELvV8Kiq+OVwn5t9eXAM+umP6cvAlV7CZSIvXOZ85wc28ReS
qq277wMS/J0xPNgYXrxOUaTqNKYnSUZEUDXwPepdGxCrxe8Rw7h573xK2knFRnwkyva52BBZA+Yu
/aIGR7axUyqrOoZHMUsDcjwECeSD+5UL
`pragma protect end_protected
