// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:26 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
iYCZ9hfB/CJWzQ9BNOhI5SrcdJBem97GfT36ootqLe7gKLppsjIrs8HewqPPRxHU
zAGf2hf33sdOhvodTTE9bgtXJOU4ZH+FzeiGocHxfSooyNa0Wh6n0ABU0tF6Jjiu
J2+eG3rJ01SiYq9+iopu755HTZNAdMQlIqaQ7GNq1Bw=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 9744)
znQwVsUyx57gzyJ/5wl3TyYXG3UUy6UhS7GhWks9KOvWOabrjy4NRyERCIOKRMd/
LI9xFDMCGCDa8kbwjGFfMlfo0DM6HnsK6ZW+bQYvGd2aDXm+Z4fmNJ1Xh6ZirLaA
+E9Y8myLCzSTwtPDvgB0AmDamF3H7wa7QODbtRY0v50yVjkAHuNoE37HPojek5Y7
KYUeFiDWJR6CXwqnzMmQF75+j3bF9Lp/H/HiKfU/oxttu/Gnoj+9iyXTfnM7qssK
vz2TkS07FVwzWmAII12IfaiaB07/NSaRV7F6iF7oKQ6Uz5If3/ueO0/O3NxbAvVa
7N+ZY7d//XDt81LnrnP/R5Dd6zcPPGJVH03obVaNc4o+u+uSMvDi80ZzR0lT0+nU
E7wrYHBQixRRBbroaR/o0A9ztmHZqW2NkPnVRGQ6zTSxKoT197ZrmkFs2gRycdDM
NW8r0qpMNnOQibbujid39t18PUX2NHiLnMsndpKYbrS1FpZ2E9+pw2EWjKUUgICa
93RrMlDvd/S25LUdbPdqIhzog1ALXXxj0bPZCQCMNzeoDincelSNalwNXR4OymZc
0ynAsJrur5uZZlpWESJsq2YXOEycSkaEpJTE9f+16RbrafCg3IweTspwx6Al7tSk
70rjXVmUJhyzKp9/v2ldyVVV5C1qaQ/lKYuoy9dY7ZMDd+T2jpglPufLni1AkT11
qxLzfYPqXON3VLenfvZ47I6oQ36tMCj3j2bvQ3TkaT5KmnQkMdBPWPxp2L3aigJ0
dIgfr6otZjhL0iYeIvx5EZdWSFvHcUsJ+wIdz3XJ6ROMFYDm9SwJOCUinZw7cyMi
iJIUj3p1JDWGJDnZdBImVgjngGX7HoqS6M26kP8i4uYGFzi4L/f4aILhEh/BSDy2
WhvKHjEoHK7R3wLPNBTOBEilvi1RhzAW9jPNhfk4Y7YadeHey5uSUnG2D3Skr35y
q7P0axmQ45zIfBf0uiZFYjRboLB1cQFOuCTiVxxaa7PIjTRgUVWP/6LkbSILBO1L
W3GLRD/ENHFSW+EEfSpiSOPCyQLs9HOkS3kTUdGgUiqcQxeYWohyqti7XaeYgTWs
GV+/kmsmWp04PLFM8dL4HP+3Y6F+vkcUrYaMNBM+DW3k7bbFh/64/xUMALhgWrTV
gkE/6yLS+FsgvrSOUJ4FiLRFZ8ENIdMmqZCCryCtyPsGFlshmZ8YwCIVEVZclRpU
jCLbahyDYDa4DJZkrSrKLEzDokKPnB2IV43tGV1c5mvN2Wt7WRM0LQlY5q8aV3M7
1cti1hvONKoMUX67x6se6sxtJoas0Ec770UmiijZ5FyWtsx7tFfZ7eJYYQmrkphd
4VjnKwAO3wxeX/6yb5I5qD3WXgCO/1e48pGXaSdVokVOercsS6YINwNvO/AeqlpK
d0PNPDaGjIFjOD7+H5mmkQIvKcWTz8K6roU64XImkNr65HpgbRppb0PVVE2WKXUb
H9WhAWCsgXcBlRyInkg3qcl+75pAlYl4eVlgg47LbPDIOrxqc3dTGGzq9oWaPVrM
hJ9E80YQaEM/ecAdJEcyd+xstpjPM1MxEOgGYl8SEMINjzABxSJJzor5SjB2QwcF
J7jioJaFQWHo+ZQ1+INz5YFKPL5nsZ1H11iXbZPCJpVmsJRjEOTEy3H5/n8bM/9c
jPFRMDFJRWZwb/WDshfjoLtV4DxMWMp8/zBdAZhXX530zmsO/bpXijAwKqrWUHGw
fco46RN9v+R+YE39DItpuqUkJ5qjeQI13inpDyXGTwQoOi+FXxBDqqWyuAeAiORG
/b81Gj6ArPNZP7zhDvzFk4tx7tUg3tSi1+IN5+vQhyqH3RrwoDHxxT4FPYowX0uJ
GJR84gfTEEhFePVFLNDN8G0HTGE+ND/SjAKXSUgAgRxhJXhJw48muvrwKEC60set
4VfCJLMqSo/0MAKwxlrpAZOmq79MzoL8aaz2U2nkg+cBE778eHjjP1ogPA12Wm04
EUsySJwWhxtI5OXstGPDyajzmJTCOjEehkZqZSM4WD5HG69nPqXxm8IUDoXrtM19
/yoQmf9vnnQXvy8x/L6MZl9FQrLJd5bvlunEbJKcIvKGabcMEQBaZsuyGXR7/T0x
DrW8QE9zf+/Wb98BKIzhoi57vQqHaezxjkKz6XV/ZDzFcty2jT3cYgvvWlPV1bSn
4yxJdSzhh2l3sK4N9SjIq0HAsKl3lLU410C06o3Sb144N1irteC1XPpEkUirrpcE
IK5FgVlJsn5f0Bixp9cdPAJoRCpIVswE+zM0u9MRHJVGqW/tO0UsxNkJ5C8bfmf3
w4fFMmmBjyRyyZl+aVETEgS4jVdiMTxkHZSNSvNvhC5rISiUizqxEK3pxYPQGHg6
g4ErKumtbcwuHjVhnDc2XRzRH/Z1deADwtjBDbg7lrgZ5+aALujBMT0BrWCobjPK
xb3+qUPyNAM3W0T0Ln66BsnvlSLUWIsfBGohRFnUIfExe5ti+KbNgDoi7YkJ97td
qvuN90JqeWpoQlO/Yn8XjeIAPRbtPFAdNg9DwXG4o3emFcV10fhEzYrop2K3oFWL
3vrPnrV9DW75Vy3r1yrS01LepMtUMOcBwpyFXYl66MFRPLVPbHQdLv1UfLTUAFSd
XdU0toBMIARaHQEKxNQlKGS4BmyFNoyNAr4BgkWv0YTB0bt4hnPPwWRu23oGqaCg
NQMgbaBWxCreXlJhqlPdO/d8Yk55lR/1yJZUoF+HyLuG0zwohmbgeOkLq9Kuyxow
3lQyYdvdB8UMhVNAdrbYNN73aO0R/zggld3yOBTq35yspOMphWWpJztQ5dWNCoC+
UnuMCmKFQjJtZQ03qZtuqoe/YvtSWeHt85ZAIduaC0i8eIhyagRW9Ro541IqYlk9
zJDIvkkM68GVNVWw5iRGueQcYiCp8Wk0C8c4hWiwxmko4oTVV4UHNtBGejEyR6xS
dhIvAjf33JsNT3gOx0BvuwFoiHwT3zIJRSj5vs+omZGRIWjoK8rmp3ww/7bTVd/o
kCsK9t9JHJGQICd5mwcZi3gi2aiWQchBFjy+1n4TH9Iz4VLm/mHRtUu5385Y7r6a
wmw5CC54lIMxkRJ/Xgl1WEaFudiHPB+lnSaU/AFGN8j6y6jNBlVV44/8DOx9kSk+
mNFQjKVEE133lBuZc4sTcFkwprg9v8YGuqEWq9Lc0yfAlGKlesmf6zz4ytvOQD6y
jPWAfRs7h7l26lt5ewVNJiJ/Q61JLCCnL3gbEXdrR2yZuKmelT1DPK6pSL/Gg0Ab
pqAHAyStPAAbz73zjoxwfEU6KUJ8br/4F4HJydb4DxgNgqawJg8bvEznhU3XFJmn
FiiEn3NHBpbpJGrQE05XPnv3QJpmpCjzKi1tKxV6eZVzwtqQ3GPue/w0uQBOvBZH
HPPJpmAyhb9lzdIgtgUnusmsznaywKsZyaPmaJ/h5qVbbkfWaUGk5lwamVPBjGNR
6LxVv53Uu7JB8tuKx3nXZQ2er6cAPGVGB9YQXt6pWsZ1DUWKBrpYejEjuoTl2yMH
bBlp3OhJ/Rx+HECzuDszyyCEteQT1qODNyu0KxLbS9JiCPl5NO5qEzrdoNCEcnuv
kN49E14O/qpFnEDRzrVvxABeODohXMWAFb3BgYOuq/XZvacCFiayHfUEMls2HBE5
rJAU1L7n/n8yR5Cg7T2zalhL78sQTSNDKn1p0bqQWAGhwbjrztTrGfKbAf05K0Ag
yG9OeTFS/ciGy+VXKxDdoII8tc2ARO1TKJCxaYeKPNp8iYAXlS0T/tx2+BGiLIZ/
FXRWqXZCyfy4ztdsaBgxDnZf9lIVub4C5vBFgQSeArZgOVi0qD5yheHOrFRONR2n
8mNmIjBiVkbID3LDKKLZkrJT7+nwPjo9s7HpydvyBdjfG2VFLtAoqVg6jG2IxJtK
j0BNr5evdcfEkL+KNtUzPWfiIkA70L5vSgApaClLKyC0KWuSA1wsF3GL/yOUXD4O
BEtzwmXDEjPSwfjnDn/rg4pM4GUlqB7F5aKFqwLPIOSppnEj8oZEUYvvWwWa3gEU
sbQIxdIAi0/TqRjdfS65aKQ9WKKLx/x9ul752Urvnpx8S+rtWCGgkL5pu5LPzp+T
4znnFp7n1RpKznrEyQfQ+4y6wmkfSyhJeqTvjsoygLxYtLcLYre4JW0J2P92Myy3
I0rkOlfo4umoh8FR6isbX/2IFYm+m9cHX2Jax6BIwnHgBOICsq7RDBIl8/WFnNrp
r6QezVOthz+Nvl9Taran1NLo8lYH1Je9LQZncvNGhA+wl0RhTW+I1I+wWjnVDtqo
rceEBCSzUw2IQ2StJfk/qMAeyrn8o9LEotkeOTpDesYtEiGv1iGT51UbmVt/4V0a
1FA4NsmVQplIXIQzv9dp53P54RIe1ke842VEIvUmc+upvGwZupAC1feuUGEBYZdX
AwYXk5DcrUNpO69PUYn7WZ9kuNys5/eUWh/yVUVFAyn2eCdKcOFS4CFzPAYewe3y
f5qUdZMS58N6abswsOneFawAT0VvIy3DG1OPpDMWM/DoYQwqkGKUmDwdNMJmNIGV
EQkBtCTs9qDkH62zTpAafW1t/eHaynBK4PkGXbiia0Mw5J9pRbTeaF3SfrDwQ0C7
UnNvtyABttLZJgQ0q2a3regjyaRIBuvEkaKCXcKAoUGmkaVZ3gQ6qqXugiTbrcpY
Z8SlgLNg/L4ZC0QHM9tUKuxPs5yDMQkzeAfR9+CT65tX9Tl9/EwfQkxnPQn7nrof
X9upXuFZj38NfEev3srXMXrobCpmrq/U5KRL+95/2kUAKehbIaZOfq83vuW3qVtZ
4fKL34kswd/HfxiqF5Xuc9AirX0Ag/KzhELJBqA+Ff26nyYp0yIOIm4dG7xp2WHS
qt03LfkjpBZq4hNIse4sLO4HnAzLOJUiIWPhRQYnPqt3o1py1uedM6TRW/2WrVtO
c70NgWBVMqL6Jslw4/+LC0hBkaTbjvw+jsYlCXx+LGZTP0yjohIUQP7ZVU3F1ouk
opLEjxSJ6qtmVHPtvDcEo0MjbsROTtAonmP0UzofzZ0S1n7QJ8d6+tXqt66+slJq
azRKBPnuDnDb57Yh4PcRds59vgDA8Sv0bpJlcqBnShb6RS1iuvCkFvxAX1cxo/0c
IWPSHQ1C7KatXCHwNO2S8l5l3C7kHvJocxRB7QKmQeeh3Ck3ZkK1vqqpOMRuaLwV
1A7OipvsuXa9XXpCYY7UsehvIZlQnPqFZ2OQNSaDZRgD883Qm6341DwG9Irc/C6f
JBULhWH1sFbDhrhWOLdUBBg1yvB1PE0FO3F4qZZhv/t9BF2nhlP3lleSg/9hJ33z
Fju3IyTIeWWf7Uo7gH+DKXhkLz0egO+5IRRRM3rYr8WwjdV9qumGXM4w4MzabTgl
G/lTwRDSssgDWwO833BqlSCE3kSc2au53eXoSD9LFrC8Wj1GGRxC9YpoNMDBtniA
RuGZOrHGl+LSzvVAdpE9Gl+fSRTOX7r9YFMMrVsNXT+1lz/XcmtjTbvy4/q5Y6ZI
neYG1lAUbftAzGeBJ20EAN6EjZkOP/y8ZHMWqXe0B4TiF4j6oDP97dOKFzM83Jfv
FWz94wDKyrhy5ykzENovUFsGVRQvvnmZ/D17jrs/S16P4FmhSalQ2VUMagFOrkLX
Kf+zS6PHRiP7x5YqdLIapiVXlMK9RTORSUDRnQk/tFKdpUn32RGnaJPhqTkAhgct
58323FxlboDWNbRZHykCibtqXq7bPa4b2Bbfo+m0CWGqX1rdlTCtgwVmzVKnNtan
p0g1cTTeED30XIvelK1fSbiWGMzOEqWhfRti1EW++ZYGnM59uYDubrFOV+WtChES
dJgb2OWjGQhpsu5P82BxyEV+LCF3v8uKTNkd7dR2Y/EPAz+FtbwyhFs5f5O2VGmX
tRDj7ROgXwUgmLs1RhgPbept1SoCRcjGxm192iOqqF5AuwSvwGrdvc3QuKUCVfHG
4SipvcBAmca9ybfGdHqg2PtcB35rY7a9nIu6XMMLlU6me3zkgmDDqGFWLjpSgpoJ
Dxu+ztwKt0Es43UTkdqX2+2g8pQoeu19S+AW9h1jYX8/LTVQxIkwB1d3qWOBzbFL
CAwdcHOvNYYyoD5M4ite/o7XPhpasqQ/sgosxaLuH2NkYXyTnnTlTap/ISs1bRYu
oIs7ZATBpyjPJMt3jnVgBUKhq0LpN4hqgJ/nrhhiBHMjYvMP4Gp+BQcvoCOaZLIr
j3lP38E1V2RrXNbnHkBZvxL8PpaRZjvB40bLTDcxZCBVj/ATaljapHq0SzO+PLCG
zUBlh8w/hbOXWduxuHLy7dsGpoxR/zUXk9F0UphLwb7iiphXFH54494qPS/DeQKR
D+NkWOaL4xMgMaLBcz0dwScJbuP65W5KgTQkRWrHf7823RrwaNiw4fwZfd0j0fM0
19CAjY+MkbOikin9S25WYkBzf0ozr+OvKj5WLBQxhZI0ddi0ugN6RTgssCGtuznM
jhN1mveezHB3senRQAGRgTfh7J4atmbp+U/VekxNTJoMbfT/kD+ATB8NlaC8goaO
Bds2LSjLP4ENR58a/KjuNefYRl9wPMdWXGUfk+QHy9pJGZhNIlMuDEY5AXdZaIsh
BCt13K74mTCa2qV9I8dHrt2NmKobagnaIdj3uqfHN4cEANpPOShjHp2tb+QLdEkZ
kgzouqT8fes34hcIoIaTqOS+7z5MXQ2qXCI1KAPgAMDm+CgfZb/7jCkE4CqvnEQA
RzsdBIOZsplStTKZnV/k/Zz4U4d/kNuypTNX3c45Ez23FkjTJ2QnHAyYiqp+eGfi
jLPqt6G0bnllrzCAPUpp0pOrytVpbVq6mi0sStUYr8YnrgOV9GkEQHNBPRPwuJfh
MoUpeaUohSmst/tg6QSBZYzYEcaOgxF17iorh6i8Z5gzPUGV7tL/8QTNcqa/Ue+Y
2qn+gRIcdJYoqOR3E0qLJntxctjYCew9rJRgOFJNe8xxNSmUJHabAhg2V97n7BGv
8nn3thxzZNNtATQiAOcrk5zU/Ek2iQPMuiB794MOoYDbw6QNuXjUJ+5toWS5oNR5
2VKILMEtmBXyeJ6PCoeF9QlV14rXGKpeR5jiXIhMD+c5CMQyZdod4YEUMLTZ8ZHB
fDubclMML3jhFe5I/rIMv4iGC0KXAdxu5hM9FycyqOJ5CsQfxqNRTDt8DDXTRTEN
vjDOHFnG+afC6s88YGpsIrsaFvzY8YL7qI/C3YTb2wGCRV5IYzOPob9JbcHtCulk
3JrO3qaJKNCoBhM+IF77Eb8pItjJu/Qo4WkzsmirynEllAAiTs4INvB5MQTYJ4w/
2bNxAAIGyPwcj2RhY/RTPRwhVtH72zxYDez/iQuv4lTfM8r9CWm34ZHX3aU9zOWy
4OXls/d+EbdNotQioadxdFpbpzE8FpBepo9J50rEsvnvmzgxHVukzBPD4zpLwPY4
eHHBWIoGg21aeTKthgdNMjgbC84ZwqGWYwTuk6Andt2IuzxRAc2k0NrMG99y+mcl
Sljaa4pT+yqq6rTKKv8warDGMpqJ+TLW8/aqQko8UxdE8TC7gMV+gUfPM+f/ET7T
ok4qKo/ZZfVAkqsHqKrENDHsaiMrc/VGs6hy2gDB1uX4mtiso1+mYrAtIXWc/Fva
48Y8QwzhLKmSfXC5JJxHhw6Ce+QqGHPvFMBqclhZcNTHZZyfq3IDo6LdAmoBGAmg
lU+aYTTh/rw3DY1gZa3oovmB8eyBv4SRlfP8yfpAjjm6T9rP0gDRL0pHr6ApPfeI
r38wysTmmADMjQE8IPwUS/NkEEHgKAZghxlNKGlW30H2t420t/mye5paM9gejyuV
SaimiOTGxAQS7kpCPiqdSpIUz5m2MSYlE6MH2bqa47/f2w8/tgfQk6Sy2gQbEq7+
Jm1TIERso5kL8GDzhjG/CMMoxmTWQO8f5broxy98Nm6mAapv5hFnRPBfuUoCiMDY
Zq2ewUTaRAAZUiTdGdjrpRfK0U17C8kxcG7y/eK4efNdc0IE4rzzmNCK6gXGtJyT
XiH/qe5tfXt77J/1tXduIsnjHlsUzUo/AL3JYhyQvqyaW1/9nKH4jKVMZWjaiTIj
wfN2zQC+T5pZuBW0s3eOE2I+5ZGE+di3TKTwzme8M7vyQ5TvXCeBbGCAhCECOOLk
D/dZUKx0LCvi3t3rb5LXzDmRcgRWfdxdcKzy/06JGAr5JXqn15YOyUGN7vlBODN8
q0EaErsXkdz+yKNqMlQ0Bd7E31i29aYOLX3fyoDn8sUDQ8OquO5fBaFSLgbFPOp3
CeMTS7jHagP/6nVmnxvZHa0fR2MUtCN0zoBZbexJHsDCgLUWM1l+80dCsDF5sFxF
0Db8gtKPuoHgdZ7Udw9Z+zd5wNNa9j0LeeXebVdKZbJtlVVn5yJV1tSzdIn8dSJk
cFj9RxSgTpbb4cwgwR4HFquILcXemspjdoACyuEfxRNQPuF+fyMjLdoAOWX8E4eD
zhC/yaO876pVttHJqnmQQ/IB+Eb+a5uU6yvbGZGPaj3TKlCV10zsXQ/gd8A9QBfI
ZQjFkngTUFQoC7QhnnIItcLU92z4QtxV5rGt8s0DYBT84bKtCZiUUSsHPp4cqkU3
sKz+X616RA2VtvnHY+A1d/bZRWsTZ5QxCbJVyQKi2du7cK94bjR4jW2Mj4IAPpk7
eOvabR4V07Pb6Gt6CCgEr93EIuO4A2wt5UpPp2ZDH9mpF5Q0eYL45Gx+AOXl6IlF
ZnLqOyY4TDNEZiFpl2YXX+eveLfHQR4rxCS1V9+AJbI+ijAeGdFp0KdSaFS/F3HK
Q5muL3M3CueDXYoDqqV8h9jcrI6VIaRHcyVx6p9ipG2HZ24wYZUipLmH0zfwPrke
i7UueDMRc751d4ZTzAUrQoT+zommLytsA30HTQuOI+b+wNhE5Hu+2UNP/M0Hqh1D
tFZzEntKLM2QKUKGKBnSk2WGvc1mJDWslng7g4fjPojHzPprtPd9WtPpLNS4ihuu
BrSB3jR4jiB0LcDmKMkz6S7snDfNhGbu1vK5dIaijtDe1C1iLJPELisP2gbwO6vb
UsuK0vqjafJes2lP9ske5eHwOZHhtzA6XQhux/+QuFqwlq2f/ca42Qht/1zptrzV
Bs5WdHgIdCl06LB0LUISJ61Xr961OSVF0NufUwyaKdOZWOgfRmh5yy/tQP2WTLRR
HsZLTNnTvUcMvwSWb6xUhdZUqcXH4Ull13g2oisgCfetH8g7AwK/mDX8njPmY/cZ
5toRB+HIh5M6ZXg3pTtk4j2d9zA6NZwAmhohyIK8UXReyps4XiUmLkrxpZsBa1Kf
TYPpqeXzq3896jMqxiY+LBA/2gqRvNBe7BRdQJ98Gy8utDaPPLpXtEYWfQhmDBFe
fNCPbDI5eZ7Grl/PED8Bo824jX10i8ZKRjX4NsLxAMQpLoUSJyCTUf4yEM35awnI
QZr3JxMpgpe3xkamtTklfMm5sPRe7sliOyNyWYzRQ7zbsc0pqlmDpBKIGDyjjPx4
Gqc+q1JLwrtMCLeq1OPLrtXA7PQM8p07SwEN8LITXvQP19zmWNASCvyo1KJiO1em
9+jpsXL7R2LK2OWEImy/fDVBZ9oitxqx+APU13IwHLCbtjWffMs3z79vrQkVz4vG
LcFGo5IfWZxyMSVIOiUdTnOlcENqYOzzPeIZiNyP3azHR4QmSxABJirPbjST0wPz
Uu4rW0SpmzTzUAWW6+leuTjtx9ZXu5jV5jxu5TX6nHzBpnuorKqgmriSLklEWGMu
3krB238O0KLOE6TOPQhvUJs/tH9mHnIpfFPcZf7qm7a/eMcdjRM9+B0EqyjWxvI+
vV1yqlG86x/1pEXPYurRokDGErx+jXuoA5LAHlb2zrW3e6+ajVbBW4Y9Ns1vRrca
nWr6jS8RTB+2qjBLn5eK5aTF/nu2K5/bhDNeu1SEzgshfeCtzhS0570DjYsMgPwl
WBUjYek9g699VpwBIzyweFZ1IQBBYW7f2uia8gY9+WQMP+mdtYNo3JhEBWesXug5
drpVMGQeFFmHLmMa0A5W+2yBEfiiI1HUNZME4IakaldNQ+LY/lEndwm+r+Ysk5Jm
UQs9wDtvkux+DYZCLsefffTXR+bGkrSHatWJzeulxLdl2RVDoxEg/GXuK25MqrQP
DzMwY6mOkJsk32bpTBFMKgKDudZia3fIzxqAfv8dJGbrV+pc3eK55KOBRxpAsnkh
K71C/u3l2EFm8gbLCxkgAWdqR4TZLFF8iIMb/pgXazvdYMjSLQ9sE2pSXLX7XRiw
FZF2zyY5v9S+jY0zjLZnJ1Y4wV1fmqHQsOP45GfXarq5yxloilWl0zULl8R9g1bp
/+NjiM/xQUdISwHBGVNXBMDaGVT8dS/tNFlZx9IfqDTHqYetQ0Bot4HKyYR0E3nr
XgiE9kLBqqVBHeu49y2t7H9VTMR38vN33/BNMM3A/KF/pLL9VHm5EB7ptUo44bkj
bQz3AamfbUqTH2lM+WrDQh0St6lQrBQaHW0VMhdl/64MrL1fo19UcpFECpwFK2X+
kGsBaQN7Jgprm2VyFtA26Q8qmuhx+cEMcBrBjVt5BtoDO6xcGgn+LhVFlxyzSmHr
aUHO7zqoX8aNIJLNew4WSI5lXHxgRYMshR+ZUX9TLehhJP7z+rZJll7W+VbRtm+x
tfIX9osLlmtstcd2eNTdp2LojJnx2kHHC3bx7sburRegRgmpuCf1l9B0XbNXWtmf
XALyyrfsv3Yfm3QzNpJgtkZHbQMelayoQm/0DnAWFl+KWSXDQAA6jgRR5Tt5XKjB
RRZAvAkZ9xhHEnTgMgqhh+xa8OEAn/7VyfPEG/XjUjxWti49Liz6dfvRS48hpbZz
AP8C112MKqUAo4ERTud82fk1tWrLePx4nyoPT068SRj3yVkeYRykhw363065yk5B
msyGjcshqXOP8+jTpwRdjM3J6DEZ//KpYXFHRgrc/XSZLpjFEfqKcnaR4ufbc/qu
wgUHVx3n2E0bXg2x/JVZ+iLBCbdG9UZO9mdTT7J7ruFBsZpFU9hHQVCGcADitzau
BdcBs4Ho3NUasyIuZs2t1L5DUpDOpHO/KNVk6q8jpVYVLkkn+W5792i6O8bcmqzw
CQmK3h9uhKLN2412az0YekPqls0xHpqVF/pKTXh8ep2cWdnVq06X8E0IUFsSUEz6
uukJUE7ofC81uIDlVLmyRYxSZGu0JlD3biVq0qQevxSYHQJ4uc6Y+s7SmjLOOd9/
8bIGUopdiXmxeRr8CwZKIIji0eGoEzQ7jyaNN4hDR6GS6p5dEx9Q2DejdT7sxL6H
+DVoIqkgyhP8LVOtZ8r3vl/2DX0KDd3/K16BAEKaoanOJpZTl2p94BbztsTAfA1R
Ug2II4v4lvGprh9Ql0893+To0SgwNSev2V1dfrjQbDRJyDiLK6kxuHCSgfSswsF8
TJNbpMzriQ04EnGSkUJOW5+DKZf9vUdMSjN9CNiSdx+DmaDkGcuKNLkkFqHnqI67
nIDSwSI0btf6m3M766EMyAt3wZ02CzAcqDtBvncwK5QBD6nKkA1h/U5QKJv2Uild
yODwiO7sSb9FKd89rC2Q+jttfrg4CtSyXJv5fGF1KRkI4opamTSK0gA6N5pXW4/x
x2Qhh+PWFcfuTBdACvZdQ5iUHYzUCXDLBvkAshmyTJ/7pHeHK3in9TRc/ch2U329
XPkWwun1ndqsc08BbDZOFLnRSYzhLHn2OdBV0EvFCjVp2BlQ03CGLunSI6e84oV5
/vpxkTdrieLfpKaa0wvxiy6SAUw1JSvA/HbLjRYAbvfCK7LaDLfT33iss1AN+kTZ
dVDepdupZ0VbY6dS9TkTMwfbqS7bQPOtt1ViTKCU1lRoGz/YuaPNyknGpI9ZVxRp
sah9xYXsCn2xpym/GSx2CvSWzXWzf9q19HkOmCB5OqW1ETVitIJOBuNDN7Bmgub2
wiV3V5eLFge9+7lOOcPeL7H4nt9J9gKXpRbuzi5oxJEvk/jhv1JimFE9TslbDuKH
Ja7WVhB/SR7lCaupSo4YbkFd8RSQp1rHaGca1uDss9163Pjzb/tthYVXxA4K0B2V
4jXMo32j/9ycOpTl6+UoXYGQTjI5L0cGPCXEE30NkK1h/oU4Gvo6GWxyutbuoT8g
eidqwC9PYuuNorK26CmHqvJu1DpMHMAKJzRpTvPvUJj22PkxA91vKWI6QOuh/Ey9
iBzPBwwoTYBrwGrbyHRmoclOTAVE0yh0bukBtm8TACWRAnAb+21/GOs3Oysik9pU
1f45OkPsbOZZ2Knw5IzfqDX5PWmxZpYVnpCeNE/TMCX5BmMXOpUBW9qpyWis+GMT
sdzdlEyua6af8uwNkyLauaHJ42wGk1GwXg8BiUg7xDSSE7Um2ZmaSaD7Pfy0/2HO
8DkVo4RZ7ZrPemwKPlQyU6IEwWvuxVGzEHkPRJQcXa+yatyibcJ9S94fzgRPKbyG
lKGxM46rhkevuxk7cXYBkrXc0nPOj8dghkCUnsOdtXjQqf4Tot8kUzwKGuShvC5F
syHsrO+C8v5aCS01PH5LATRmuvvGsX0PZuqYsU93Nt5AqXYdhSufVNW3POhrVs5X
7pCzpBdcO5dFUnjlzjWXSSXxMRiqy7RHE/Q2HQrOtJ2fUIoOqG2Q+ZndEG+//IE9
3pcpfiq+Pt2MiZiIjgWjE2r+1LznbfPd7a1zpBPdoXk3EnGrAZ0w9qKYG8iDhfkw
UqKQJ0WAmcMH2NFZW18lixcx5c7kCDKG/5onye0jl9mnWGOQ5hjYbf3HDEOp2Kkz
LdY7e78XHpLqW9rK2I1XyBv1pomUlmbvysb6FW7kerRJKlHNR9NxcC7sMpNgVCZ6
/k6OuYBmuuzdLzZtsU65bFvMA1ldYGoNUTkHVcoEedEECiTvbDJBq6TXbYV8dqsv
YIacFfJTHwWjizmV2f4P4ivFBsnqtRnyNFYrIOftY679e/Pjrk9kdVP4xeLRG8S3
5kzPiy8FhGd/H61b6GKa07XwGhImM5cXtFXMMDmzR8EUoZqfaS/Xoe6XNojSE/q8
`pragma protect end_protected
