// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:33:01 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
lrUip94j7UTDDPGEPA5gmBEAN/99z39SeJMlhzbDzuz4xrZHxcxLR8hq/j3VyLku
GZ4oKBodrPvohZImre4RQYJXlaNU1P9N+I8E0UoGpDiMw4q+AjV7w1y5OWGZFmTY
BfPVAFLWD/b0A0ySQhyWfs809uA7ILJIzKBuAe2bFdI=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 17472)
ZtLVhJR0U2Ilou6eea4xTLrsP0rVeclcwlMAWbmVM9xKhJEFD1tMz5+E2dJThVQT
OrlBRR1izXMkiMnpZPr5dSUbaO3JCfxSMBOmdqsuD0Z8s63llpAb5F0vB+1D/ZsD
Qv5qigBsrzNnxVJ/9QGHlGk8N5GF7DTBWsBe0zW0cgfIteKeYwX9kMW2AnRxs6ry
flEqxwetV09Jz6GV869rhTHED4PpbExr/gcbHd4zvs/OIV/AOTWugkQ3Q4bRTSGy
4Y3A3AUiSXUINNmAoW5uTYKWcLHb3/Ce4ZuaLqh7nfyo5gK5sP+d1uO1fCsINgLg
H9FVhk/46EPu0ATZKTlsyNW9oZAUBRhTAv+apHDsR1bdmNl48DUqjUJYNV9PeqdY
F8PF3Pb0sjqDbX3j6yK+Vs2MNoPT5Bbiu5EIzqKqEcmDoMQPaPI9X96TN4Fx+tY9
LCwXju7bmV9+UDr9GbE9rR0C4HJVNEJv7DtGNvAcYefyLx0ElxrzmsqMFKw+TsOr
Qfkx1ELK3E6duakiE/lPXBOMOMIaj9QyegcFptnX1X7yaN8SXHsByEeazw8d5P0E
Vr2pfUMeIBebXC5TvgQNCmY0FmrbYLueW7MPF8DJABpOoxYeppjkGoujYx1u8Zo+
jeqK+w4K/StuQssdO2iXGvzivJZd5fduSRZvmOKAJiZiziEiZ/2ybppdC7XPQWEa
NKNqDXuKRJ2uIYLPB9LE4Qi0iea3X3xBIWsmJt729xad51aMGz1chno8xSh/adG6
qtqMYHB39FlJShwaPRwHbRyNvqJKk4ZQUsnQ0VU9UFsbTKHg22LvPPUJjxIIbUq3
PWLYetZq889KGXgPc2U9skmkogEqvEXph1QFXomshK6GdKJEE84uVez6I89sptgl
HWyl6B2qpcHEtVUeFvKC5brhPobQg0exTvF12NdCRcF1XtdutFT50f6wbj80JN8h
m5V0urubSmDlZsasYZVzcCQmgE9bL/iqhU8rUAIK5OOmd59IT0Oe01h6DK+EhNUe
6vfD/9bnKMdwxj6jnrb/0CgtSldFu3gM1vrggCJsZxKFpBqe92Up2PNDyp7bvtG0
oqKx4CpHYMOvlfCQJ4zDItaeTpnX/jRyg0xQExInP/fppj/rxmzt11+8zC+PqCAH
jYRH+K9cOFSuoGLIkUM5aDHP1EyW8LLhBHItQ680hPmzL7zGiA7Bx19rOeu7ScwI
yxyQLbWMxoPjaEgRXkY4/6DZWf3rDvGYwbIrDKibSD1lgiUTjFF3UPbJ0VPKaSta
E0hynlRyhw3KDiLN0CeWHCNuCyULLDw7c9qVqM2s4GThFHJD+joQuBMwaEip0CDB
qXQE1GFFhzat2sHfo6cUHV9rHC+NH+2y8jbtowg703M/9CYXMfZZN4TDu/jRzaM1
61ylXf8rvyMZDqKziFoFBcrgO1LcLs1E7tGznY/CdsRBtHKxJyGHFAy5m/ZcW1vH
cbkXCgNDJgytEVcyah/Wc8kAFV2FhqMGAP7WiQcozGgeSFMA9v5ogK7L732vxn3G
nXam5jxOGAZYO1K9IhlgEo4c0yJAzTPWPsfg8Ynyok6SZXN/rvWJ4v2TNNtKnnc/
8ft9jlhQZfs0IuM2m99BW8J2fhGioyiJZ3FFjHX2M8ECkPzCrtBrDW/sBZfMsKAH
GPyY+UmNBIADmfOEj+Xmdog4GLleSu5/TQBNmOzcn1lagLmGmWu+VjHwkyggGwgt
Sv5oBkc4rk19h2KwodGDJmo39Mf3obcvQAH5s7KC7YlBn7k0YocDAf3KBSe6QSXZ
tpW+UHNAb6FtEm9rfAFvZ+Z7V8i1nQNLB8nCWrt0w0OlEOY26DGqtm3Mf0/lT5mK
HvgoHMY+OPwFwVX4WUMCeD8BmZPbLqZV2B3dmtwhWRvjTC6kERIPQenf6cSzyYBb
o22B9UZn98JYqCkzXYHUKjoo96mS6bdHku9WlvUsZEBp8UkkkOGx/q64DmjTyTXS
EPgymw1V5MyuAtVOV3GrhOamOlyieANd6bXVAFVpbnCMxq80NPcmzeT0kGQk0Sfm
E3cLh2Gz967AuhrAvBezpREoAwaSFlEA2IAVauo1jYT6Rht7EZ//PFPj+kof/kfZ
giVfK6bHZS6pbYDOMIxeHMIrp40Bsfhq/c3jC7wQEkL3ffpEiTKgVnvGb5UqAvQF
kEYtDIuOdHD7CaxkYBnnLlXG45t0LUOed+CI+W0EM86LnqL5hX8sA7f7LUIY2t0D
TYfHg1jrLqxW0zwYLZhUv0VXBKsXIwwGy3kRP860qle6pywNG2vBfvzmz3Q+Z7Hv
tFbCIHjh98dIvCyMQfeXLKLBMFopZmmHr1I/9LJs8m1uVk+OpfTsk64nMfM8feID
ItBpIAnYl3Z7vvlR+xOXHuNY24pj6YARdQHXlwgxEucm8YwsmyCmcsjN0rDgBWgz
NGaCStEYbZ1gpfj0BCBV0pCufrIhWUxcBSWZKvkY8pk+R2Du5UCF7pKVq0S3TvY/
LqtPf3aCe2zZOxJApT2rFe9k07haDbiHix7YNdXU2onyraFDxr4olqAZuzFiKHJw
heoaNT989m+OErTvz7j1b/fRo7ExYzMav/mPKdoQmYzer8O4XmtUXCLjocGX9Idb
qCsLKrkvUOi5RE0f/mralbndfo5t6qTU690xtNeZR5hp5hS1nG/J039rVTVdJPQV
RMFIIxAkJOXC2BwbLnTU9J9Kd84zerWxHH7jpG9m+V9hXjeuMKi/dWsOmQJBO+sN
2Pi1vPHgvqYCVSpAb9MYOnTH9WgCExzsRhUh6reiKSuxnC1YCC1ZPUalCZqibLA0
LHrKa1JuYZLF3eY69/WRngB8M+7RG1H2Dl/UMwFAf+0PEcwUq7z+EsoDHP7i7yN/
WPlqydwjzcQ1c89ygWdSJnLk3S1hAc0CAXmeGPvt97glqKb5XgxPTsBLwMB2Ud4A
ONyhaGGSAAtpervZyiBQ3Ex50BtnS3TgQUEYdqBEgsFaPCdjlYyu6poaAP9b4Zby
vwXHj38Q/93/wO48IFEF/r5wV7QQiQhXC/POsvLDuHAubiec5AYHFyMh2z4SF/DJ
lpHO+oeJ4ErPuli5L2p6ySR+q0gCEQMGNb6Rip7P3dL+oMpjEUcNRAwCP88rGKG9
muIeS1FK7/CBqAubABMBZTF4ogNGA2uDykQrdohLLB/rTh7zgab5GDZHrLxG5md9
YKcyeO6kdkAr1MYHTA7aS+wBA5erngMxK6Fv9p2ZcyX/IY2hpirFLj12Qx3hSEmH
ZTzwqvJKMQL95k796WIe1h6mT94uhbBq5pMBab3zivonJx7QqlwBBVGHsKUrV+lj
4Pk9GnkjHsip8OrK29Z5YdSuVKXB6jxknORH86VIEEl+vqaaZpXKp/al2V4hePLm
3hNaaMpExpK51AYGufiTqKKFJjhmgHwddYhscLWMU8O0iJnE1qGsC3nVpK3Zw1eU
BWDsaFZvTNXqwbhcGhSx5TJ2XWYdiMUVQvBB2xliefpUIf8NN9FQpc7+VtMUx8vI
ByeS0kdkTACz/A3Gd9/em2Vh7+BqfGn0H9jdB5A9SYpN2YRf0b2/MfqcI+nwG8Ii
FgKDvnBMF3Q9ledUmLtU5PyCgfI6o4dNIb3nzGUnVWwG2yz/zIWAI/6EzIB8fBq0
YrRENDvo1MZYODmj2AguI5X6YTXE/gXcLrNgeLXGw8BwSVGN1t6Xl7lHKxb1dfRV
FLfmrZiUHvECXN554OB6Vt7r+iS60K6WWC1JmPupZdFjMiGawa5WhwrWCJw7eOGy
d4+qqcdN9oi0Oysaj/IjPgIdSDphBRxzpj/6DVkeTRKhkF1vuATj5L96JmpRJNz5
Q28iNdJzndvQzVKQkYU/NianBMTPG/kzhhd1GziJfTGjvLf9Qv9afKIYkYtYNGO9
K61kIH4WxyeBR8RUhsEBwTA/uMi52fTqB+x5zirteoQw0Hq/spyqrGLWYJ9YWb0f
1XEcwwlDjxvEuxzc+LUX4+qEchETYm47J3ReiY3b1xRrEJO/og8V5R7nELgriDJs
YnKCvAPXw8fYrHFdLnrSbaSrJry0A+2pE5rp7lVqTczsdJcB/55ct/p3OyvFLw2i
DFpIH6gQ3AaoTs41RDx9D20qSdWWk9ujcC2y5hd8gzu7VIK71ejDMmJ7IGly1o7W
CvLqF7u1cy57414tnxdt/FQ8NWThV7OhSGbnxx/veZtmwj1W2GQdLzkh9U6ZGlyS
cDnwvQs3sKxhdSCsCywxELddM5rm6P7gvO4/UuxyhB76mHTPuBYa3wjKV6GdxyqA
tvqVmagHs/cefwuhLG6CQkIkSdnXbE6iT0tBRXGdR8YIpfD99+VV5qTrKfkTFWWT
udyT0t3jB4j+9bwrZyHFNC/shgbx9k5y8sJaZqGJYErhfjXK90J0gRiEgEDdR1iE
UqzDLRCvkDY3SmFpaycRcnGT/K/OfTkSMaKgwHLG4KbZPrgYjHAYNeIWynboKP4q
27s2NNAVli8Y1SQ1hKE/CHKJAQcX6sc4qgH1JPsg0q3Tu/QlW/sKKl/8b0FCRlMF
w4nvXszKu4TV9Z14VcAgO5/3YEKcvDhhAWJ+kh6KLwq/ct8mkhDAM0MENMGLKDx6
03o027o1Rw1yOv3LCFs1LSkuWKS49WrpwaZIag/gB71G+HNgzV/kkeWkKSPBYeJA
ERq/5TKUk7XIAIsZoP3TqiMMwMPDVtYE1+ePXGRHayWluzRLg1WKPGaJCCE2nmF1
KnW7XwS+W5B1ji2gfRa3BGekXcz/RT7p7Dk9ps3SZ5Bpj2X4116Bz4ZN1R1B6bh4
qvfxaGxgOTBGNYgyPFm/UfZ2j9iGBl8yGBeKcpIItCbwUk/LvFIadNxlckxYasTc
Uja4nYrnac58CvnzNn5v9g7ZoJ9ugYfzsaxylJSs0ZU7G5g+zrNoaJ7kT8GihevJ
vqfFTexoAdOyS8QEaosw4ayR0tLQkhbYBgvUkQyMxogICsRvayIzQVcEqGxA12ln
LOSr4P3+FFs/LXgrJAYsAQIa1mOW4PLDTT8AO9/B57GyaLDqznTdwpLdLbjOlnEm
c9+wDkd0DOz8qZ9f6nU4Vba8RmE+SYg/Ov78/8sF5urfwrfe0z3K6stGmYXLPMF2
klz64EcLJ356ryi00+PguJvtQzStaw6vZOgYgFkiOS38DVQs4wzFFQo/vWNnjBj0
Up2VXORIGZPun5HudazRpFhPNrPIZY/z5HVDZPxKWliHZax7WZrIx7U5gtDmhh3h
IzTzF1bitgQpw47k8fMyLYjsbGVxhRowFZfDYg7bgNvegTHkve64fJlIYV1rkqHM
WqhU8Oh7VjrAPz0MPgBE1FKrqGbv732pKu8AJClnC+UXbl3xsyWaPWc7HttWqezo
MdmqEb+r6Icmi4v5LLmbzYWS44TMBe+81ndsMHD+C4sHoTMxHmALyE8T7FQ7VwV+
lPzPqPyWP7MGKcItupqGMMfUoxz9ncssuy3cru3SMiJSAkCkMtX8h5jtQsyNLsSS
psYYcmxQKdzsQkMptbd3oV0By3n7DtZcoiNg+lv3oU68gjNV38mibqT5tfaCEyH/
Yi3IKYGr60eAhT9Bz2lavO3Y0K8UZ99jB6ota4l9jVH1tfwKCV7k6yxs5ea/IKQT
R66dsZ4eL8s9dCYtXgMd1WGoNSI0M9Sr2WKS2I/spKaehQPhdqi9DvY/yHzV5Sk9
EfD7kPGK0x4rkpIxvhw6zzRHbBGzpmwtuN/YkNO9rwukzPzr0Vn/Z8v+6duHBV+y
Zqs7er7Vtcz44lsYtUEhI2I7UHE5r7hxWENO83khpeo28q7+c8GeTcCvSkJTW/64
uDBuoEBoP5eSmWCqEXmw+0OeymwmgQCtXqkGO3IC5I2eSgnuiIoV46xY87YbaQYx
yv9rafABNSLMik1dYHGN2EQp5dgtOdada8TTMMKrRoIrmg59seyYHDvDqmZkM5x5
UwuIY1WwXaaGoeCp8NckBBbHUjwp8WI2X/7D98JJsQcai2d3GeMpUZqyVztKyP8Z
/OoZYv//onypxkx2REaIYDC0M1viQ1MVA5w61Oh+tu3LRU90fSpeCfVzoJJ0MVWe
cg0Jvc3F6TCPlHOKzDBcXLVhart9lGD68aCEqyJfzMhL0R0ZuPNC1mr+J0iAsb+/
CPTFZslKlmWzkBggyHHt/U6AQt/9Jpcb8w6hZ+cBdbrgnzMtkLwcx5z6uN0SZe9J
tdtyi91T80394uSisCYi5aiu1tcZi69lX72DTT+9tDQBa9ZA400aFAbkrFV9wQAv
eHBIQ2zcYSv3773eJKXQjVPoxOA/N5fY+soclc9gi6FlVUDG21ReUXIVR6IKFFlu
W6JgwLzkDPIzC1Qk4jHEehko2EW553+wW/c+OhGJby42omJLf+lRSd7KTbMteiwE
/QC8yD76iO1cddAUMvk2vtZkvO5f0JST5jkKTGB61DIqoSrTnbCBChQ0cD/BfP7y
6Z6/2+Hr4lH1NTABPiA46vToMFDdhsQ5DhymYDIMT0Skh/grkEW1pk9JWy8eq7hg
bdZR3PYVkdR1coK/Z1sgBxv2/eflgRHGX9524/Tn3/OlmNosgC4XpHmrEt+QuT+Z
Yt1pItmCEvRrdjo8mcufQ3RxEnhif9Cyd9VAGi6qCpIxwvXoP2GdiLttwSaPgEIt
F1fCKvJz1btREg6ptkrIDNzZpTpL/FC7efiFonsIp/aSvRSR7VIWzxvH+4kx6VpY
ZK8bHIoarFuw1M/wb72zn4MvibUBKhOG0Ym9ryCYOGR/FMZh9JaRYtqxGAJkU5K7
QGNhYF8svvNmTugZAREsWQaEdfonX+BOXg5m2+SRfjuUOCe40zzXT4FGl4s9RB32
lSnBLcAsYo8ZN2j1FIUiKBUUIank5W2t0sMZujfmNCR3J4rb7WOmbrTU91wOZ6qi
7AFMH06XZLtapRK9qhfA6gM4XTB6Pk/pB0ndAp49m1ZWp4PMZOVJyNUu3mhCrXUV
kMpqokC6MWunQ+K+CJaU0nGo1ztdP53u6DXc9Vn8lN5RO3RTran/LTroaCcoUIVO
dskdqw+G/mlYtiIkr+X/PsbR3975Cvp31x2Sh37iFfoKj08FfVvvE+4PZAmOFikH
Ea5x46lnkSK2Aknn5/RCZxjuxz9SQohSBShElDYaeiilAUaLqIndZRizynbUpCP7
8YNDP8RVF2gPwBwiZg2AQ5X8Rlap61NICXaFXLUVSdrC0bzlXzyNp/whYrEVHgA/
qA7KPOw0Phk3rcM7bpjklamPjvFGSjJ0C4MFrAf+iQY0Q1kVuM24TYW1cty2vFS9
ira5AcD/D73QBoaWQ6zcmooNg4RzazQZzLGiGTnRdgGW7cbpQWZzRn2HqT22fZ4A
4tk7f7Znx7emmWeHYKFTWv+WQm254sbErICZeI039hNLlbHrm181nayU0NOLxP+u
VnSWEmysaEdIURw/KuZImUlQpgZKojJXEfGI+pLB6tCX2ooO0nItIBJRKRuf1isR
M930vIYMRxv8AHGiMJ0xtpV/LlH9L36VZ+FvLCp69rGdYJxV0sEYJicAoLOJsOQ5
4av0cT/kKrN5H/QTAn3J98U7CCGafoG3aqszunzmXKxPxuz5fmXDTqquN0X3aFSz
4Gtqwqk6yR+pRJtz8WHY5+9Ss/SlawXFlobNItJHnSWvKdlpdv9f/Ihx8rfO5n80
vfR/J8UI6Rxx/5bhwA+zyYXc6RTKyxoXCioM4vEn5q+3FP5Qj/RPdiY2O43inVaf
W10kB2Ab/0A9lHJPHHTmzJys6qavBO+xMF313plAK/VAmaAL2p0BRzKs0ABnbq+Q
fGtaZfNvqFUw+HtVwzmRXTf1p6WGzuh6/ObOtllLQPBFVrZH0Cpbcn6Jm8xyjw7T
6WmeUuc2X6grB3bp7ieEFLKE3qwv9kgCHym6xUBCZJIZhX7dZLXBgKEkNu05NtGu
n+DgBljQNBO6zlWZb442eJ4ALpUz7ybSB8oBKzY2RJmm6m0DWJf9p4mEVIviH3vx
rbiBcOwdGRoBnsTFO96IH5FCVc+xonpCvpvdTAgbNBjTy56xpiypDGTodoxK/WHZ
jFATL6SYPce9/xR3SoSFBzt92w43+bypR9yFI+X5gbLhoh20T2i7afE6kfI4r+8o
GN10ReYY5345KQsKZE106VzljI13LA7qA/uVuLZ2IZAqMp906/xStd7zhacGJQK7
yUA+jI4wflyqTG/l7G6rBEBPOQO7oNkp1duVKwdvuA6ESHs5UAe/6jXlgTHRh3dK
1vUDTkhSMJWXreczzmk02au4DRVKWm8DTtTiEbA78gdS/7S5oKGSU0KNELyU9KVx
zUoMeiu1RJsanxpQMwihYtgREziFOcBZzBTAcquhMMr+GVQRIeeNnEaBcagm0Ho4
Wo2iBMlsxKiXtgy3m/Yk9yQNghwPEgFSIvkcppQepQhJo6NYXFaUqLWVVPHBF+xM
gXCoeLMDhUMiBwMxOtT39k/yINWX4Orx2LsP5Yq7HqDk65TKqsmlbOzBCnDFOuVg
vnQLPr0P1kl5EYLAZdCTIMAbaXdDKxAwHcZpSdECb3Mof2wy/1qCYYPKNIS1QnfZ
gnP/+aMoEI5MTVbTkse0P3WHg7VdBz8T7CrQVvpDBkwDYA0KDFn+XpbNGr4jFiO6
NDU+KSLUKYa5Z9gBWITYm2ccSoJlIQ0HDvPxZWcrUOYjuYWRHAKJhqGj/RbVJS3p
teFxtwI2khsGh2W2Qzhtbc1+GYip4DCPp0SxHZXpZpz542RCjsK1Q393AtpnopXH
yVf2iIKTLcPUxfzQhuGrKcZP+uXEv+wXbO7ZUSWFMhsqx9b/VGeQvA8ouWTNqwC+
4zGrPtlK6F1NIFTCR3wIH9gL9p0GxoqXcQ3Av07gPacYOp9AVMUJ/55sTSDd91k1
sR6mYRQ8FgIuSezoLujgec/CGnI4h3zDxykG59r32/FIy1BOD4e3KPPBANmgkynl
7StbIuJUjDW+Z5ic2rOUYA1Nwg1E/3In9UEaG2QYrCWjfezzdfoM/ETF9lnp3nIb
j+w4slWXyf0TzvlODX6G/zp0cASMkFyozhGH9yLlVZFjZMJYvAnLz9WgV7XM+48a
MjGi7OEwpYCBVSXneTmMP2BFBHYS/hIywofJzgGWl00rbq7xAcC+8r385WwILZij
Jo9H9/h6BgM7q8uoSt1Cyzl0phxZdoOOiMZ/J5ib4XIFMuhteEJ9BBt63sG645A7
PNVp5kTp9QWSRA9QOwQgrNSznK1HcexMbKf4UeZGsJ5wN6Mq4mQodY71UN5McrrV
MtS8RDm+l04wvGYy81RDcM0NYiRZhFBsXvfsKafw/bDFdgaSA+/RmBMdgK9wZkXg
BBGbWNX6D1VwYPiA4NnU4YL/G1+7jJCnbcJ3PQ0Ws9sWy1eZjjB7nm42sEzuoAmL
HIzWttXqimxsAQZjRD+/QOvHaNePxLis1LvezaydclEBz+qPF5Zpn+zBXrCwnEOe
kvkIFrnNiPT07xaTavAZ9AvBjlxCK5AZTO/vSDAkLLo1Y6UhZ0FkXiQyXYMLa80X
uvqe9seYMrYiyUZ1uTZJQZr2iSEljLWsRRrk7pmonYukP0dkNczc4HL0iEhpmhJq
i5OQRKF345/RrQtMzSvFFh7eiOdbXkFZa2a5cfw1sXgIXHm2L7aIbUc+PMRVnoCT
124UfBIGHQ5B+K+M96b/QbhBcxs5X5tHOPzFbdw/NVGrjWrgD9Sskr3Qop90LQ/6
SgmiYGSHr02IqjwgZkAOKOfxYiMDunYEx3YMQQupYl6bLNJwbyTIAkKspVbEqxIn
CSFYvF6MOduW4s4vnFY6SHvgkRs8De2nkY7hTbfPBk8Dgi5ZDvwmxzNqObTWals6
Y9MaF5vZZt+qXUC/2QIOuUNDQMt3oANpUDcKR76pKBnJHtB0ZvmEcg8wd+75FmDv
6vJIIdn/VBhBtV41HSxSdiy/hQADR2hD35hJS4x9/WDFSgF+afCQWCNiEYLpWhak
XxxIkvFWS8IPXs0XUOUZX+g54ySK8xkaTM7cHzPXuPbKY3gFEHAjdkAU/VF7K5KV
DVMsd+6Hd0GMswFEAiUzVUNqS8kqKVuADGRa69q5qEqEuz4yoH03RnG6TZD5PaD+
8KiTDOKOckyFAm1c8Aw0lpJo//MDVXSOgRwecgCJ02wEvhrDBox/ldZ8cj2nHqwJ
kyVLy6MPWEaJ3AYLn38dvXtsiEYrIe1r2mpAarRZLjGCW/pEGB3unMVSz/DwowIU
BFhKxP9YEiGhnRaaC4PnWX0yA9KNXQkYn6GIwY0uqsseWo54Jhqziabe0ALSrCZl
fQqjwqbHz9kqbJG7ONujFzjETW0Q77apxQpx/OSHJgNaByRR2sP+7C0vsHGA72V6
ZG6R3gj+7gipMLC9Tw4Bl3+Hqhmre71MXUFiMKdT2evsW9HpAZWLOnsNuYU89wdV
HhtXrBgSQ0T5PuWZo0dF0IcHRN9eb4zQId5TtS+XvuLWZZygbr0GIH6bDWpngQ5E
QlevhFzmBYcyCwUQ4/7VoGMU7Tlv0GwqvIRvkDhU8t1iDa75CpfU/1cIT/s5jbRL
8nFViQJjGPwcWLKgQ/34na10HVXkHn/5qzky1J5AKlm2YI9PpaXAMxrcQr9si7hb
JX52PmOsXX1T4ct3aMDZx4rY8DRIYt82wjsA5hUtVsrQHzveT9rwTe9IfzAzhg2w
qfs8SmpDKZs9zpYrfPN9fjZ8l5go/ZBtM5n9nM8O2z9LaBRckMKcImliLmZxBbLH
c7IB/j+5jLdtKzoY6kJS/dd6RaOo6hIE8KyuWLCsijB9ESrNygjlRiHv5lgnh+N3
q4QugfacQipFO+oX8vOA8SivWaKnV8jzcMwaDWBT2AGLdPNE4T7xr4QmRe/W2o2J
yIVnwhQCZlEB8b+gFw5chemG+hlf3k65vvWIZVcW6flmcV6CKXeTxmPdGkNVj/8u
G7OsH9tPqACm64u6Zzq+utbR7sYEbmJZXR6kHX1OC0bwzkaNxrywF2VmZWmMqdM/
Lquu+aQGqMDOSJspvoe5VujOfUDlQFojOkNivdbWbHeMVuyAgl+SFbEe3VA10ptw
CENxESTMN+4N5NnBviAdyKHcFwf1WIPTR6TLFZwqPsyNdc7gyFYOF2uCXsjxphm8
q3e3ILZDCYxEFLgJy14aUWUf1iR9kstlYsiX2R/dVYrMxbAcByMHfY7xkO2RJsVy
Xiu6fqOpqc4obvL8nXB4/YeAyvdhkiDBPniWFZHXwkDilOEhtKAM7NqSEo4/vp5c
YRyjoujOuPYoUet9ER69UvaKJMIwJoAO6TMS3viks3OtDtntZvsRyJe3unCMWiBs
UdVM3dxQdQk4a8EqpJlrbZvRsXyWBo9UH8I+Rmx7nANK9tT7iAek3qVQHm2nF346
m+A8XTzcJZIrhgvrwGBeoW/4q3JKDr50hEMG/MOkeopEp3mAsBvDGC+WZCp9uzDZ
xX5HTEHF/GAeELzsWSzIwrn5YIKLqVmK3K0AOjgilVJyUeKCOCoq0eJqQkcROxim
SKWKb5wouHuidVXguvFScHiICisu10+AmXnbPG4MfWKwc76nuH6CZg/amoyJ6/Kb
oD7fTsEdXdDt3zj5aVoJipiqqz+5gg/6Ley1of77EKl+cVrmTLmZUHG5OIBxRUnO
NGllJtFRxGgRA+kqN7m8TcH9uYH5cT8VSr/aFX11ojC+flSeaVkBSoUrmZKsby7n
e1PwpCKBf6+jCpPsaq9BtVBNVq2/SPp+g6QfT7kSwjabcAtZhIYdnDhBa0KOJFkn
SD0TxhKFkYJ2bJl/CgvSxOFfB66vvuOzPgcP+eqNrd0664zRVLLY6L0RDMND7aUn
Pgi6U2Bnjx6ezyvZ9sDRG0oqH5mSb+q0Kefv2iKZolM4mu7dY+QORTihzfWHPrw0
cx4V5sHhejfJdbvwGAfYgAsPMeJedbtlCpJHN+b2o/VJ5z7kLVra9R54e52O29PR
sOj4PIWxHMH0TYo5my8xWyZLoEvh39f7jUc8YaqpVAi0TQOS4sP0t5e3c4zHJrZc
fo0vuTLUpeye5TPhFEimGtvnwZq7MEvJk0OlHPy4EfgiqiKtQbXcdnrmraRGm/E+
qK4VbUzAA35+WfHxGu18ECJlQKE753cl5h2U+lHhkacPjL/Don9w+g5lm9kvG87B
XYiCvBN0gUcQN0v1kDqheCLL7D29MPjp3Ybrt7lgoEzIbK5MXuOz0lypvEB4TCnS
ItWluLiGXwpgXTDdAvitkkmlg1dkhHrQWxjNVrywFDqifdBj70XjAxmLyS5gDMmK
MGL7gn3zvMewCEgDYmpWnVp797AzIMbHAS9TyzP4UjKWI9LCA+EMrGoSkJ+uLxTT
Cy8DfHZZ3RJzB7S/98RPJVuPCCKcpJBNrqE1XQf3B2EvEO3JH1w0LbFiV6Vka2pT
4C6RfE1TuUWC0y/LOr5LTbj6mvnV0JtxIYW5RCgyCH60V2OMFhZqsfWnZqbDlCmv
A4WiwgRngVmWrvPt2/ePIn1pwsbxw5OIV/YnsjZkSG0sXsfdJ+bHdMpcMJ4NtO8i
1w2YhB8ZoupJBfJ30jkWyCyDdg7B/xhyYVZiVsBN1bt/m0/Be5furknudgwRFaAX
0EmfH3S5WOLIUNDsZJ7Smo8or+hazox7tKL17kgTAhyP/p+IoW1nXfXcpWbeOE+m
GBICcwn7qYM0Im4tl/y73lYF8oxcBiIXVqRMrp4o/C2RgOba7QiOPgoGMGPGtPOs
B9Hcc/3XaSZjb96uKxy/Wvxf+4A4lUMWGQyq9O66smtNk89zLGjArNcVwyyFSuS8
QrtEbdpPM5IWBXwm26sBbHgi0VeI0aNS9pZPkHE9tKeVKzIeEKghdRduiShA4Rxn
I/qdPHlkaQfI3d6OLBgeOAl90CUbOM0+qH7zsQdlTNOHqKQ6Xu8mSayDM+dWYY7i
jNHVlS05F2cRoDX1M0qT0nApnvtnnPDz6U/widXlyVxjtk19sGkUzxBM8ys1mEkz
kDygvHJMPaS8GZuUsr7WJ+UoegyseLI0HITz47UcVRKooCQTI5EaWRfurTvkKhr2
l9VzWRS7fpYpCyHFJaDUlgBclzOR2y452oqccavzY3elMXmAVLaAcLOe4PdM2ao/
vc95iIkORwxUtSYU7pEIQp81ANZ9MsViQQfr3Dhgys1cYJjTgW0GJSHpsJSkx/3u
2zilrlCQumYu3hmT7S62VNkEVXmLbDaKDM/WVqhwwPaeCbvAIM8JMcc74gyG0eTD
vT1cq2Hs3aOka/CgGt8MeSgJo58B52vre87MBsQiqnh72SknmzBxnb92Pr82/nve
3Dl2EKv3uUXZpeKokeR2eT79wFufi7BWUeBi57GzJxK7trC9YSdxUmTkt1B9h4S3
vs5tbqf6Ra+T0nYgqOZe8Xv3Z8ubT+OfNqxxy9HmQajy+102PubfoOjofblpKn5W
VFkpxq6t+0RIpveppgUd9qSLuxC0xlWv1l7zVye4/Lf0+IkkOEIJdGlY/Vg67oJ7
O4syCKSy0mGgojEZJFQW/gnLbXBLiI9OihFCFD34JaPjx9XLySid7KywNUUK65jl
QG+9gLX0Jwqwef3g76YrRM8C4lTEuB2eN8ZqOhivDmUChtnoyWxiv8c9RJWFR1Nj
uLzf1QUcW+R5KrC8PnF7excOr4DKTSs1IfR+XiBwFZ5I/RwoeifpWQsf+FHLXR2a
8o6rdqmfRYaLZxX24tNniZxcs4AV9z+b4m2xjqKfGhxWcu9AEbvQ1/FD3te+wTC5
rqr87teAcvCaoeAe7l+uafMqPIbXlUspfNkAjCGj9ilgPsQv6uy+iRFHHWE3wZWG
F6lXw8VJjGScA6+NAtlwwW2FSIxau9NgmShRf9pKZN32cWyo9VTu7I99uMvpfbe5
4tJo3F8eWZywhkUSlAHgK8JH8X4Bd5wE9b16+8nqBT06ittqQHa1+SZfBYqPBpZ5
Uy8C5Y19Zt7+vdSKkqlwh0aX7Z3ppRajtnWX8pNX5LpZdWVGDx9mNm2b/tC1cvPT
wnuVR+K09K3vJLcBFG9nBBGEWCxPWHsEILY35NkfPz/nqn57korAjXar5KwfJ5C4
1Irv/fKlDVoOB4xYJeERApBxZnzlqHO3o7UXUvRAbgnTtssU7BsYTP52fh8DJFi3
EbqXahEhRfgHY3KTlNlKPd8majb4zEqxaOw7P9t/97i2wWYwBSbg9Y0HNAfqsjAv
Mma2LywjqbMRzNBtU0GeMkFlv7fg94pKbSIL1jrYjP6yzQR88tiSN0U3SpysvHVt
tEiNIvGt9M0tLog6OqlEAJBCFTHjxli5WsHsehqkqwkPfu/p+v+beP26URe+67u7
JmS1YqjyNLRK4VpLRtAKXiv6Wd0ZPTq7CHUBQyB+ENTCzKLIFfMZRZ/K2gQkyrSH
tYzahlZFwrRt96UtEyHTNAVoT5wAWe6HLQ3jvBLIkpjEgc2Cwj9WI2S5422IrI5E
oX78tMezdEzUFv85Bhe2K1sLUzC2B+IKkzc7CBW+mLUeLPXSkPF0R7WeLLDGsF/v
j8DFUQ4hmvWcYXcS3qXrvCHRA16m6hHQl6OO+iSeXHxsHBwMKyIq/xzlQtGuFsxl
Hvvi6efGsnpWcaX8X6NCyziG3NLfxYm/7BxCa5uh2K6c1fbNUhUUO6R2gTm5OF1m
khJ6YHNNpnU2Xx3KPWzRyWflLK4bDRFBgWCNrQadF2lLDA7nUehuHVNbdJFAQYqO
UPVznFQoPUsSYo5bsGghlQpuZz3cNeUFrXHlL2luL95Hph7V85XAe01aS7UfiYTR
NlsmCfk5pmqUoU4Q14Mfa0ad3gJ0nqkfrF18HMJi0bqR3/iTmhl3uASiz9QHvL53
J+T1ok2AbKGBoGw8I1/Y6sEAAKoqxVosx7a/LyZrb6frEAYjHuXFWh9tf3kKeYnJ
D7IQrPpjUQyUIyaTFdf4mdxP4GLLM/f7YLn2geZEPJboQBu4IuC3QocNOaoc+YHo
8GlJPP6tHJsX9YKS6DYSrL9XMyTps9onw8nnLl8vHEHT3KSb2tuHMi6GKNLO72XR
Ms4u8K0PBDCtphqUE+gvCMiDw+EUFy25/dPZJnRLx1BfMjYZ4Q69nfaecpIP/GUd
FIuEf9MePqt9MaBkMTgy8qEvLxk/n+mph+LqwL6hO6U2VK5rqMTfp/1zCiSvFWru
1rHzlEpGd0kACxc0pm7lr5PhBPyzIKD8CyFag/zks8nXTSo2d+HITG5yHltreki1
qR6BqmX5n2sWVX5gzvBUJa3Fwyt+R2SUQ0TcdaataIm4BbbuCQKmU77BMN1tqcoE
4sS8ZJVIDUsJUIc91ESqz5QkowtV1XNquMdXQ0ht/HgUojkAg1rGHpAil37QWaeH
prCoxcYZdjFUm+NGZX7guJiPcaT8SHO9cCHVJaD49KhvjN5Usig3HqYvN5befCMg
NVa1ifFvevy1A4yZNaRXJhSn2/wz13fTmj2FsyluqgeET+f+ip792V7ocP+aY9Cw
SRTHpZ2ESFtcyRRpM2vuVVsHwvRHeVAmo/rUryQzu82EzZynUsH8yCizYjA2zyb6
i1lz+IhQgxT6LxCTJHKOKjQ4gAoi4eC2K3wMmLpIIloegQW5nsgXo8XPjy32W3l9
KV46+F+t8kQqPl7hx6IGO/la4AbSQNcKvXp/lOo6Yps0ebbgkGiSWZzlwzg9GBSq
Zsd8whhMIruapcqkbIz1PvI+1Nw5FyXuRM3vEAbcoEI8twDqbZEssecjBGL1Pzht
hl3Z3kwf431UyS6B+HJEX+m/LZAzIwMisgwpq3TzGfKLqWf5bTRqW4Pi+qu8/mYp
2dXjygYcPKPmHPr6vsUYQIKiCA1noI2MLzVYKEwAn/z9xvs14oAwXYVjv/zuJ2oG
sJOWy5agdo4CS/96yIw5p97VpNeKCyzxZLt33K4WeCUeTiPYQvIqok1uztLpEQnF
5uAdLfFY9ckdBFxMDHmK0JEwQrkAkc+4NA9oKoraD/UseGrrxZEtc1Ayt1/iqiRj
8dS5/xIT+JjBMYi+nzNsS08XSnvrHmpFfpD2yxGHO2UWS5z3afH8Mi0Jgl8MTP57
PPGKAChqcfm55nKEEey8m5984Qv9UJA8YrSI8PG/CURvjcpcD6ghnSjjfUD9WXyn
pUjqTQtvS+O8Dx+/qD3cRQ3/hDI32RPIm3c5p8Rf5EcEgWvfLIyZ06teHbq3TB9V
ViUPOdolZ/3B/KdhClOLId9r2AkeCNiDsHiV1H0jNQXXr1J2ptmNhRrdOp+eQZAC
XhCHpnfdFJOTTCeKHEK3BDHxFI3BcdaDsVHXllmtic0VUi9RqxxGuG82FUl/9HUg
ux8RqvGcXk0NWdksMtg3N9NW1q8EiY/sExAV9SeDwlH/aOcJ8rQJ1WqeWetuGCCh
6ZgiEm673KmdqWQrDL1/UYTP4P2nE2ECP/heZGSQEznh2f1q/9srMxefjul9TlYF
VyWBSnj8XZvGEaAmw4DXIQ8ypIvBgqygYTX5mpuo9NEkQiXZuV9N2/eRcI5X8vVY
BCSBXq736vzBDztD3zXVX7lBctiL3+bJ4RpZR0i2L2cKtCrVTUENZmuTvWhmPhTL
pcJ1fcv2YncXdvAE8qpI/s652Wg93SxFkyZ71AaqwaxyDp4SPpxkC85fw9el0nXm
HI6Ij4IWC1wbOa5OkifewU1zPIwlhuDzXhVBdU3NKUD2f9itUPRIjnqljpdk5oWF
UvbZQZoCZkQIvsubryrepE88OcIfxxwoLC+IITq4RuNiQjvOoJEa4IVBdsWvxCEx
4nV9rtnhZ7rg1xFYWuhZr3IKBLZQChS5ccY6hRYX58VhgAv9CI7PHcHiphMniY3D
i57rsyY9Y/zYrZgJxKhvAqoSfDkYiKKmpOn4+NhWnmEWFZ+D199UCHSCJApFNNK5
eTWtPNukTCTAiqwG5GufNlnk0xzsmgkc+UoAgDvJK/a5VinGf2Q77c4J3lXjt0fb
RTP1/SSNh2R49zcrjiU+He0DVUyaq+6WutGkUJuGTOIox7xo7uJHChSFMNa1tdap
1Ar8cCBKEsZn3/ChSFNQW5H+FJmQSdt5b8JZPEOYsY9FQwNAaVmf0Cys+UmS1I1D
2x7g0kaPoDRh0pf9uuh4H15Z8GRvRMGHfzFxUbsQo2Mu1Y2TdQCyWR9GZ9T5uUub
+bTe1sCMtvrseXYr6nuYLyDa9MixHQvNOvLa6CKEP8ybtwjLJIJjCJfD2lvHMWlg
Mg24xOC6E3kfAnOY7IBV1xG8lrcqYOmYPJPfvKHe2fSu+WwdrM08SSOuUsI+x5Mc
ht6TQnJiTNrK0mXeWD5H44fKQSqnrxZdXC65CGkO4w372pmiSGLdhXJCdzZxPkKp
l83X0kb+yUehsMfbVPo0vVQGBX/7xpVbCsPC3P9XHOip0NCPGfiz2oh3j7fPHjAx
+ZjvUBIvU7LlIUgH3BJN1Rl7XZV/JoC/6r9Tr7brYa7GV4h/T9Cj6o2umRImFqWz
grh2ZjrTH53RmGKCTqHc+N61s3fiqKWbf0kwXgbt5HSnDKb6+nP2ZZ2xmPWxopIq
eW2rPtxSrnVM89xwPeN0K1mM+CFHvEHscbL1H+uITNP2+MsBnUWuyZ8vQ1e30m0D
F8vjtsAIUnG/sf7FzLy4dflGGIqkCFJ8H2XxQrtllBwe/NEFwf9XW10mBjTJ2tfZ
DTeBBafj/lCfmPBzmgalE8oqAGPt6BkcB/0BVgc+6jg+4LhBPbDwVxoI3xpp8U/W
+Hh9y8J4T15+9yNYdKBcL3T+LOvvfgp0Bq1Mof7DnAMVikhkaY0GSDcEfHZ2X7k9
eWcoWsPFtY7RFBgHkWoy1AbyXVpgavbhLgwgNMmOQW+fP5Xh4RoQattDLGRmtU9r
0x1IgkkUdfdcf0Wf76ikZYb+qAfMj1Pt2kPKNVhXyekEdWFjH+esVUiWY/BcGD3/
DurBo50YKHW23jyMLR1z+x5daFKQYe71Ub1LaCokynZBs8aZ80vhTILlQzqlPmWb
vGTMxAVdINILowNaeXefL/XGdvI/tY6BY5Opp/YbsRFBVliG3y+PzzUUpCteZ8Z8
mM3VjMcCuOAL6PexwBRddXTtaZMd5mCMBKkF33pcpElBuuc+CuUGWGxEPqk3wd4M
B6+Gn5WSZRdqNHF6HhMVwTG7apNyUr36rs+MkPZr3ve6KJXfMr9BAyiHR0Jh8UWk
OxpObTPlBO24uo17ust0++A1EQUQeznlF8KNfzEeBQQ/ZSQYTCLf6Hs4uvnibAVD
AY2YYo08bK6Go5iqvgcZUNZ0gRyG3OvsKBWolsxMsPtXAKOAdMWHW9jR9MkIftDY
73Yb50e/30TToT+SWMGvHwQwjZ4vhVJY0X8MSJM80spm0J3qnxpuAjFlohJbRrCB
bfF9ZeWVSCt3d0dprlspDBMDuqIEXcOuqIbxEjoB3tLqNGDjVG67KgOjT+eRc/hQ
t69v75F5bzbK1qeXnq5a4P3Ye1sYZFDkZ2q8eB5tMnyY8azFDg9IHsfIQabRXZrc
yRFH6foUEbhV15FDNea4J9XKbP5o5LyFEhnDa8vsr/YumWfmQe2u1yQpXc8AjFpt
Kd9+iEiqVw6IkMNdPLTMno3OQWGS7a3TzEtkBQFKOZi/ybWKg73onA9CMEEb+LTE
K/JRvHP5VdsE38+WucisJwDQ5TwTbSlgAZAY20zjHNRD1U3uZVOvq881DJxxgxay
f7qYmJA+1Yn8f1SYPvptL7TncFKysQvfE78EOKcuZS5V9bAOi22MsGfMCegWu72H
ReNXB08DPIvRYFwH4dMSuGU9EtMkIO3QRczQZEQvEJ6GAjb+PcW2T0BHwExkBdvt
8dvluJ89fektY7p44flqJ35nZpPHfcObW5XanBiGivw25vnYxe/wfxZZT5CSma2c
lSJ1v4Xcnc1LI1X5OuT/XWsdeQXzuPU3do1DRHdKHxAsbaenL4ZI4K33VGTvWd8x
wZmyxp46GY+zyIY+QTsJ5YUvDgbFXEmLXBA84URWx9pEPXgEOCGbosbJ2OBZAKj/
XEdDINAc7zo55AZn3qu/DrCfiDFLXqU1FaDYn7uU9qK1Nkii9SdIdS2lVTIVdqe3
OrZy+3EhK7R7UQwYg6VuvFKKkOFpMvbrxwpdZE+qD+0O6NEtEKvy9PUvX+rnyPco
9SQ5ognvHJy37nE2oloXVDj5llFwkW/mxA+xDSAjKdjWZM1eAibucEPEhsSPSFk4
jMDWyMZpQm6wh2dhuk9ApqTI5LN2+J97rg+Gyk7d77kzLY8mT73Wa7H3qr23moMp
9UQqUnkHZkW+Fj+sw1bW8e3p5XiRlBXITq992glk2TRzhGlnYj8v50av6qd9uGZ6
bLj1mjO0JbKD04EQndz5dnRCg/Top1JgTqvduNK7C6uy5VOhljpu2iQvFE4TIJwx
Neg6m160zu+1kFR37CiCU0u5oCI7ZECbPAlmGKOzxgn2Zc6L/PqQK+HRYW/P3HEt
beI3UzV+IkON9v9QJhS9tVCs01NuBfDI9QoaPr2JIOb03DBuWDXZs64L6xgdnhyO
5IEhReBAHlDvPi9diyVbMQObeMwj7YImdvuz+zT9Cj22etDo7gzjwvGcolerly5j
SVyPzCWZbm79PuoQfEAijrFXdy9uy8O7Zd1pq0xjyV7jYvcGjejQPMAj7ZJ9hM7Y
VE6EQtdgTiKgB1bnKRNwvX+/Euk02tez8YuvJzzcabX0/lWPa+ny42mn75/VGCxl
0tYfNEDAE80vWf8Cduc76aLmKZGhc9rUFyjkt9EFkp3AabqoTZfMZKhpOMZQhdgw
/ptwQhvtHahNiqyAszXj5tgKzTao9AJUJIxhpW4Z8HtTG2Ws3zlpn7A0NDTamfui
cBdaUZBBU+31AmpFT2dBlVT/CU37CfaXv4CR1JQlt8lKqnZOTzf1vTrQxFfVEBsY
1Z7gs/MBEI8tvQ9rU+el1tztdWQMNt6hP1gVDJu172lQq+g0S4GQ5VYfwV7kZP8d
lA2bzP8SazdY3U5yL10dr6kLUgH+O7P8ITRaKEzSjODesVka5r88GGU0wlRwGvsq
iO1oWqAGCFzvvpYzG6TXT3LM6XmbPdu8pj8U0zZLCJa8H/M/uXWr/UZAI8GXI4nA
x83igZavqHGN2tembBd98tEfmSKY4BY8zDtVCcf32hWphoq9vXjs0i/5LF4C/j2E
KemIW0Z7KeziJGqKWgHKLTnhFBc5kFgOpcWL5SAY2ylWkWO7Au/wsJjPukk2+Kcq
ZK3ezIHDO/PNBJfQgskUxRtGx+VWcYAkeVOafqXmSOkRqmltNHO0EUPA642ccmyP
nqjLYfNKoQJ9X0eTMgIpV06WlXdBdHe5V8gNTynPpfJCd9mwtt6PSu7BGwOArY+H
0uxn4xzZkq1plJnn1EuhRSzqQpwQBDl4KQVlcBdA0i+K83MHyKVXIYmKdhM0tiiP
gUxxRZ2+JshxDPgOy3J4prCx8G3vqqfzBXbR9buGsV87e6yB57ZhoVkV5OZw4KdX
6WeqgRDu59B2LlhoJvuA7DOfQAYemWUh6tBdXCSYXMh2spc4+30IbcVGmOizLTi0
PPZu1YCB7syEWHWQLbmlwGOnhebEx2FSGB4ikRHdPP8T7IJTbz9cf3x53XM9SLoi
GAmvrPWfar8CjsKzl84IF9Oibwu0kEjD3qDOev1yJ834UQItEzUcQeMh8c6C+pD5
vvtNoCxThlseNNa9VZo8S3HErFxGxn+ySG7b87rqzF1eoXHvyJPUps8kvVEJlICF
B42FGZgtdMSTGlDn9Xcmj7UtBBxdZ2c6xRt+g6ANQew0YQRfPVlI4g8yjvlL4xqB
t9RpW5JQUu4/3lhFTXwYiYNs3MRQD53rN/8zfuEmBGGR/ylA70upfEjLMdE9fQ0l
9dP0nxB21kiia3XCqdWyvF93lCWz8N0XSUAtdr2+k4V8WmexrmG+35XHjDJqbqlb
s/JrnH6sFB/yiSqQ0fZMokm1qRP2w2iThsAvRUj8TR/2k1+sMRhpVfhGDxy0rCri
euELjXXtGIjg/THoib0Yb3c5ZALsUVh0orQ0HphSplrLyCzA6MmuTdIPBHfkptrr
p3jdA/B6giQK+SWL434+4EaeuDr0t4Ia1y9OVd/Gt27DurijT3gnTbN4+j/RVath
htOoOUlROxxf5k0bBaA0AkvTc3eKJvoKSmR1iNhesAjRWaGlWmL/t7iimt7LmPgm
bvcsjWNg8E0KY+kxBYsp6cp1ndaNthbmYyzDuVNIKKE1qKZ5I1QIR9MQv7iVNLez
8cdLeS1YVp0Xi+B4tp8jY2PR5VRSPHDkc5/AtuwmtN0ETjr7HhvCJDL1nJaq7wzA
jvw2WjC9RK1aMX63OP9i8kqUR6B7rYA8icDe3S43veOHfO+YYKc+dMtp4lxBoJ3N
dZ1BXL7pEqbYWKlhpJhH8PaRFFKg0i54UEa6NVQLyKtFNE/HNMcBtxFw8tUaLaCp
tIE/WJTRcjCFAYUqjkPAsjd8sqCZwejB3JJ3+iM/6xiwvuF5GoFHIxY+QzEqXjIx
BltUX27EpddbL6bknbI0HsDvEo/TAdnNCkAk5NV8pzGZQApHc2wz6WZbCaWKC6Kf
b0FIaCNbjH7hHYsK6Z9Ewe0IT/3pNsJvPfVlic8zm92Q7m5MEe23fKHFyBYaHjYi
miauH4f8IP/m/BEjlUgxNeYE42uk4N5Nssi/9fEuY7PAygJNB2umJu5TCmSwmMkp
3EYse2EDhT5RKnKHGxEGHwckwZvkifA/voTb/d0i9UwSPWXDplsNzJgiBoANQpXU
V8BqXDM31M4Cw16xEqIricS+Ofd1VsEyl6rIod6asOoYlRPREk7tl98oDjAyNOs5
mow0akOmg/q/nUYRCcW+rahcv6p6yxzMHpRgvfws07WlTowmup876bI6e6d0Ph7k
cHplrazopBxKslTWjbHraA2cYq7iq9EfKW0u78w5ERXZEPZ96bbvYb97jwxUvw86
NZow3AW8gXJzO8KWxKnENMLmGlw+yhSgzja7wGd8XO7XcSTFLV+4e7cDtc2baaf+
4CwZBBX0PFW64Te12E9BelyCketloK0olbGKtAxCS7GIBQhQnNYpgic+kynI1dgI
RTCjhMk4EjpblbwdvmdvCL2z+JZx1ALy49omX12jaZ0uTJtPgKh6RZ52WyiTOmYr
VfK6e8ZgQtjV5xvwYiOzAWwRtzuVg9ak4Cj2pMOLevTblaziEg0+Ufwdwr24Sb8J
yacOA2FCNZoZBST25ev5GGGWILYRjCvW+9frsaY/tAJhWHNnoOsk/nYlJAZV1LHp
kj91znIS0X7u4LjH/OYwL7UWrjreF9steCDDLXY6VZ+qT+Bu3jbzyZxfGGH4oaUY
wghEkF4WSQoHmKE6CyVmByFfqRfpbLGCVEQypIk3ucyOGu2VxLRDsyjiwJ3hAuXT
oRmRTAuJYjTj+BP+B8EX4q608VC5EjGvrvglj4UT0Z2Q5UMj+pZnI/B29OAcOB1D
Twca3535HNom4m+pn1yaw7CwCXMJILzKbjRGoJ1vrxgq1U0fa0ANMQ6o/iG3yE8e
gV1c4fN1Z4Vtx7qhtKMrHKCy9LYS+cJsTHGJ2FvhYb7CUFFhxL20xovwCqDq4yZN
z8WtUmNAs8vix+wzzbCHvrzhU2m2pBZ4vxiHYT4nAwuS/FQtoAOKT3JIuRLXfbRb
aSbmQoBOFsRlldh7/fd8no2bxV7TFsqlTDDyM8Azbn37LYZ6yXqCItYRIb+VGCep
LUenXy6YYemSuvjFMkQOm4RPoHqhhrkKwJibJ5CX8W3fIQAaFXh1mEwYYBZAxH8F
S4vwXL8hKlwHxyKIF1ltcYRZ26opMJxFZG0EgOniOFINgJSLqRvexTbuyjTuAfMc
4uwlRikDUrNEmfBcj9jTnmRvR3wuW5OiFjE382NraI0Rhi+HXuBRdzKDeFM3d3gu
3FVyFfUmYAIqadYFWZ892bJ9W1Hvw1jt8uxMNqilt5FeM5hBO8V98jPrff1v2TyC
nZvjizW0oAd3HZAOqxHbCz174IZ1+S1gnGHRgSAMenGJ3NOwzN1C5LkGeWFbR56T
Zd40FnHfnUAXIfJGxaogaJmNvvHvfcNvbpEXJrQihC/3oE0/VR+9uSoFJECe6fQl
SqZlV0ZxUGNYIQ05RZsgyGrBa3NDpC+HXfQgO2Wyts3t6EN3MyFOgkcKfU+DdK4L
VpM3uAhd1QPrBVnH36i5trNnbUekClPVg7rq2eMg5xWDICvv5+eyBryCJoem9Wxk
X7weQY103Wy/4LiivzjDMr4IXHLrxfPHJeo74eIJDdPSu9hbWn3vmsTGaChJjoMn
`pragma protect end_protected
