// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:35:36 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
kcnY3r0MlEJ0VgQO0QsfLZ6rAjjyZ5mdNbH2wUb0dEHfCLKubV7WhQKShgX+KOTv
BeZGBRWcRRVHtv5E8TtKofvKL0znqQdHB7pRWIQTxABhTP2E+FWglqR2ukfeMbkO
49ebqhFSxulFeszXsV1eUIxim0ZU6yQQCmltq66U2ew=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 7376)
uQHcUD8mUqZktUh8803uXh2HN9bvLa8K0GfgANBPggi2gbL1DYBOeiRpg5MV0ulK
P75ESFhE0bnO02Fgt8CSTbpKbw+kTVvQghC9BEZQllEhSb+w8/GvtDvCsjcyqfSl
XXqNwZE4cYQFGMdpOnEltCQmuikzUrc8qjhR5hgydCnLj7CuiSO7IIUIxLr/wdSh
W/INs1ZLAZuKbM1aCMkiJGpC0FoZmhA03QQlmLtBaLN0n3XZKNdPAYJxfHyE0qgB
q8H0oh64aVE0A8zWE/BpVSE6LkWLKtUG6pHTIoZ7J1thR7KnHg5QY/mbUh9CEXNS
Ct9r2VidHF2OZTqnAdXJexCfz3D23PsXYHf1gXcuKT5w715fYeyIDSRsdIbH3H0c
eQtreLG+H3xbVfU3lQ9UCYRCsnFzMeeDohJNW+LNPxSwgnyL9rD0p44x3TJi4231
+sg4/10cLD25VAW7wmV1NAMPZDkzLkDCIEr/CHg7AVY7Oei1UuM1czh23CAB0sfP
r79wdGQBraWDC5UJDqYzC0RYq6xr99wOlqvc/RcHwVPaiy5dU5OL9v2CBPCjROKP
Ji1EH9WwVjBYasPTNHO1gE9lZbqmpBMasUXUAFIIeyG9BWvfbBEe0p+VjREGBbSr
6gWOJARPUHzN6qqmcgeGtFqqra31N9KwxK82tFTAOSWcfQpUEejF52XToOjEWPkZ
budRp/MpmwjrWguaW43fuI4lyJNjrJIvIW2F2OdvdJvFHeETahxZOncVsNkKSgMO
MEC4kqjVxhpAddGNJFKBFFDdOEnHfF37joEvH9+1zVL+ljYUj2BbHzEB3kDZlwCN
JPJEwON4opftfRUpkoEcNMXeF9s35fEsgiyPBYjEJuTCyaVIR7hXvLut4dGNWjqx
5dOWDfRkRygByEkNV/CMUBo189b8yrVIivZ2bY+08icmgyoKNYr7FwWzE/cIGRPu
t5UeqJoeCcsSas2xwOg/i1dXHLr1oRYA8VFSsmm4YEz+5nmjhBHmqHWi2TXrEcBg
lSevnTNSo4QlfmlJFdxUVq3DvxJMOqiXsIprK0QsydMto0FZA+AHflVuxR2JrULV
x5nY7D/al3PCHgTx13jo0x7QmreXZYVVr7gLSV48USXWlUNIwywCmzkssjzo1yrU
0S4TaaiXnWaPCn7KXIRWBg2WV+Aeh+9EcEi0C88QjO5jl5md6dTHc9T7M2VjMPbv
HK+TQI3iHhDX+hmGUcsUI85E/sTtA7M082rBZxMknvPsbe1/jRLLkVnjoRjB3kCi
5YJkMZ6jeU9NC4rdumiCRgg1ajCupiKLB6GC+QdZ8STg9m8YyfNplL1zvHpp47MC
66c5ATQdLr0ryq5OFwDakpxA5JHhDi5UddQpX8cFT7WfWeCv0MGupLlT7IRuCk6X
gLHAqOYWu/9G3NATUm8fGnoEwT8MubvD+NlaV3n3IStxfNfkd9QJJc3/P4QEP8EB
avpJ7LqZ1umaLCA2y5puGCMX+CmykujPpBneMuMgxyLB8UYxA5NlzClQzcEGjMA9
6xFodzAWjue0vXroRqDupfMQjZElbp3JeioY0Uncwt8UXS9HVMkMh5ZM8WJrN932
AQhAt/5aaPnRMv4p6WsPDnPHWORn5fQriPAefCay4ChCF3BCEiPCrheh1opW8yYj
jlvMlHh9l4MYAFT0n9et3Zkn9FlFZVFPXJvvUvKZZ8iogbaX6oDBoE8AvUQ2ci65
ZfWaKcyvHkTvoNWhC+NhQBcrkLyTGmWxJx5acE9vDPNvXaF5frB+yzqBZYsj/IC2
tk6B8omNQQSTcyLdYnyTAn7KolSxgq7bui0LKzNkUi0epXy3d3a0wvXpxOzDs1Q3
bCgAf+nuz1GVa5jgMNeQ7bRht2OKW11BQZ8CGTWm46zjnIisZHAUnQJkUfzYcBtB
Kbk/dmMEIWkZYa1A+2Th0OxN8eKqOZzpj406B5RLPnW0fAsa693CMd6WVSI2cLoj
+EGqfx74Y0mXvfnoKF8RnKIFaKqX/XNGwv2r/0IbLpoGqqX/OkfJOj2F6NxyuMfb
7vxgDDpotN3oE4plxIVzrnEsfOibyjdHHJ/IKx2bzbs8z6Q+Ilcs68MNcV5w7SZq
L1yX4NxWNJqRoHOS+JW+QfpCoNhhX71LXiTX/nYfeyssWB8L81h52A7/3mXOY/+u
35aE9PhrFs+SCLztqlre0Xn16ukJVXt1LOfenZeGgtGx7kMwFDT91H2Ah1dlC9UU
jjAUaYVmZnnKMteMdtZ/sRa213uhiiApwB/bYaXXD8KIV51xjbjdMwQjGDofnhcZ
CAAU42UpW3tcjn23bsUXdjaL1clCjeIcgAzQsrIJI25XLRp0d4vtTQ05Wu725mBv
qPgvVOvQMdY8MmfATCxx5VXh1eHDgRFTXEKZ7FS3LZczViA2m5bg14vHx7AEbehf
TvSukSz3aVmF4Y83PQsrLMviWFdEQkg+r06dG2woE0kehdLuoVBZBrO0U1EUFcIh
7U9V0u7fu3d4fTssiWE9kqLWs2Du1I053WfvB3TE0a3cWWvrjBuvyW6dOaH2jDMg
pd6GzrSxLd0XorL8THNcUOpqNZl6qZ5g0azGdLBwPR9jUwCjdjjH7+B/UZZLQTd+
tbBJaCDhMOs7bOf3VUKON17wfmFKdnubbUdAcCoviaJaisrtHpwMrA1QWnHhHZAn
wrC7mMSa/Lt+mLYkDYuywv+9yTUNfrRGnp0y4yqqSKEnXS61DP7LLVStejuP21VF
zg93g6P7YrQLScuf39eZNzhZ/2QwveI75YcT41bfKRmoGR41mrPwdi3pJPnswUoc
XCiqawU6+yePgewFdjRgxH3NLqjhf9u8ut7tm7wHSLabXpNaZRULBdanZRyPJCqv
zWl9EoJJEWtZikqBTWKSYjovSkVkmHPnkS4dHaLrDSE8u9Lmlt6fy0GLxJkUl5jc
DWdzkgMBcMP10mGJeuojiytkSHhV4HgoyK/D9SuabuWSnYztxBiR8KHqglPE58Ep
zZpn51eEEXF9bZ+njXse9wxL+Cy9o8j+rpBiMM8sTrO0Umz71SxvOxRYThooeNaE
ExCam26R4KQoDWtjPbwn/p9nMmFVfyeZ34iFKFyfl3tNjWrBCFl7POAdspHog4dQ
xFSarQcGKswPqF9QbEyqft5gRyXEMQ6EfBlxam7JJI8yAXLvM/SVrsUwyc8gqjDv
Csb+AsEhI7U5WH+ic1KoTWVr45sMDdvn0ORqPIzJ9yO5c2UODRJutN+9oWv+Nawu
WXqgauqHS5FiW+feRCn8CzxiRExwxwrl+aLRoiRDpUL/al7HXH1wRstd+Qf7jt3E
X9wCwOijyCingz7N20FYLAuk9BlXEzDFh/5k/519YB+OqMlAjBTZacVzH1sBO1t4
++rWMpcd0t40X/mGdaismYeYbyNXsnEeDRx0K77+fcidoCr9ErZLDJEEl7ZlI2nz
+rQLNFazUfnhFRjgIOMXUcBOTQim7LYSpd988RG8cS3SNYavxyKw5suTdH2GR0Zq
WQqsPClsX/nNDzTRqbEM+V6lKTRNZQlRKVNnSpkWQ62MGOg/7YhHFOEXyZJ6UJ5T
PTFCkmJwFlEk3jbUCwE42HTNEF4wSZHfSmVKBJRgSPqYU52PIwSLfzGoCUFHcLzQ
w7uNSEcOsSup4+7PgRFrswdTcpOum+pahio16avjh1UKeS76d3/r79ODzV17tgEG
MFR3FCEY2IyvObBA4U2UWKZbjFEVctbvK2bUuoWoFps8vHvp00EXl5h4YHvF6HaC
oNE9qC2kyD0VYHScDD8iB2ITiCvsJ+51Pm8/9LRMfrnLQ2lgzwFQI91PFa+O1weT
ledGsG+GX9sY8Gm6iR/0bfKvpImj3RfhSh7Hw1Efw9nnsh8qqrNQa73flkKBCYpo
//tAQIFlHDRo1gSmRaD0QqYJAbmjG5XuEyrLX/EfaOgJe6+XFtNrl44kxsqavhLf
eFseK2NdEphmR1gDW+wIE2tneuYB/PtgZ5IgxBhUOHL4CTXPoDaLcZyDocYlMzbt
NDuFhTmIiPFBQttEhj29cqcooG7kVkLGh0x5WOaZrk97SL1AJKgUL0aXAlGQ/jvp
SQ3YbQrcxnr6szfL2p8m102gGpwOYLRKQyP5U4I+z7mJduS7lcTM78l9JiwdCCJv
L1POskWTBp1OYneTJ/Srzl4WMMUquTuaMDYCKjujpe4EGy++dt3JFrm52NSxP+yH
DFJT93gM9BgAI9UaVnCrX/dSmF+AYjLrsXwQktE4Y2fT0+wPRZxwGjyaGwB/459c
pBzgrDwgsUhRmqX4HM42dXo8Bs3o4SrsGJt3ABwN9i7EStaB/bvjwXTwXintPHAQ
3B0rKotbvJH3lnTGxdXMhTOm32wAwqq0/XitUS1JtyFA4k4acwKOvy4PyMUs3xbk
Z5RG9JrU0tgKZGxgj7oSEK/bfwa01E3nqVtt+VkCYCPAwvfnGEdv9Zz0oc1m16zf
1yma3hf2vNaNNWhw/1aN8tZK+WjsS7PR+djkIMlsSj5jsdV/dMTnuxV85P79QHP3
/DxBNbybUQuTd1lHVIDDVupxRbEYZtoXdYVQz4y6nZuztkX/bU3pOFejhXu0RRFP
3a5K+bhnNNY1JDCMINXMWdmmO6z4CHCXTh8NsomUc51QSBPkqXOHIMngDZA9UBSI
H3hY/bmZIjux6DxdjwQtzQpEKWqWzFoeLotShpEnVKGFVl/IYDvRMlHSWyDztX0O
bXHFjTZMy0xwGqvdP5+VxhoWJBD7QiRVLSTjayAMUp5GVqJPjtUXK/0gbO45sYx1
CmrkUQJfD4yH9fwd1vSxhiDle70Jg3EdBO380+Jl+arJnmx8Yjsl2AnuskdYFOat
be9GTKfvQ1Dn5V5LZ+km/vIRPiNFiucuLSeiFT1fY6VOkpPfea/Ujkac6V5YuZLz
5n7andMXqKtwFgTHpgRgha/OQ0IzmVAlvIWfZ07WkWbavcjfK07YyBTFTXgjduxu
gfU0julk/6DMPDxHScg3GBJcqkm3s6i/ts5OR8bGAOmTusJ0/5ANfTO91zjnvRsx
3NzBeyKkKQZouwI1rD6gHzgFr8ASk9CGOyZofUlp22e2TRXPClFnjSBobz4Q+CLC
gls20kbnrbAjUUHtGfcqgBpKynPOF3Itg86UbCL9TMAUHVYdPMNBeIAZtoTA+Y0d
aIRBcaJrR96XQGi/hcTAr2pBzaF8GOP2QM7z4eMYkAFksKlyvFFWpU2h+iLE68Rc
3VhdlwW0DV/V5/eR2cjX/0w8UpOqYAN/cCPUg9eODtS4cvB0Pgd9ta+szi0Vwsz1
YfwLpiWGWK2HAUZUkmozD9fJfodRSbzBaqIvHxoNaGU5foSOwyTGJtrSmmdoT5MP
N46qC7+SgP8wOA4lwTTd9SNLta4Tt8cffDgFc+Pdq5NAsjs08QG5wbbBcyY4lsDh
M5+r0/bDJvc/amP/+7tVfN89Z3KNuKIrs7i4KkLmzMHKVQX+zIPDsHpF8ZMmJeu3
rt3GcGREVhG+u96Pu9ZT7SOG1lBYS1LWo236YvdyFYE8hsLZvPZsNmNU4xkQTJLB
HCjgRbV7rxYx/mwfXVIqeijmYXBcn74bu10LneOcGIGXCUTv7cbCAQz6ljK9PhU0
DxFGQdnR7C18PWD683v2/P8g4zRN4VA8FhVXyqoMDrbb0swuzUmGT3Djm/lGtGKh
2ZglI/uZKy3GEy7HSWu6FNKEOU7+an7bWdUWcRnJNiQ+RiHfLJEXI2yqBjEWR8TN
5hb11yvp9DPw/+KQwZ8JBBr1gYadcn+mJ++/MW/7XFzbW9Vtl2LyMJVIeQDSIJT3
+aDQNtus/H/ixE7aQwvheWG+afX/o0/Y18JocvrDt5nfcN6DdZwJERMPW1bUo7cE
aSw+Pw4UmoR2wliG3rI7itBi+I8FjgEjusxOlexc4Fz4QlDCYx0Q1CQ7+oxQ5LoS
VOZ2qO1va8uHwr//ZEVnt3fjNrlWeU+cMulfOMMcYGq38gpk7WMbRiUqNdO5CubG
l/XD8aAq1BrDtPCa1YyI+CFEJ+eG6k4yIYVn7jRmDH1B5dyaTEj422BcOPk7hDfn
HbwIW95Ow5EnLSDx8L0YuO5aVvZBKVpQlWLOsMOEufDyWdB3o2A+MrkYychT38yZ
FYl9VZWlNXXH/8LE9iBONlySf5YCpO8xoOJKzFEShKq1TD3cY//qywgJU1ff12z9
elSjBzk1OYsWB+5MYOlZaXEgeo6Sinnm/X+VNV9Q/iTiqxsKR2USeD//U2wIO/Bj
n4sCQe6nwR+GQ+NSRcdaiotB4hKm4C8NRbuKpluIkmeyD6lb0xYrC6BxvlZiY8kU
BC8QKUlvplPMb5gwk/lNA5O6Ay6gD7Gef3jNYc1DGo4TBorEDOIRvDKauDMTPcoO
Hzs7oPA5EdjuvlopyCUDJjAd21fH/KjYf2Os8GvhutkOIKPHBQlSnfNHGt4B6l7I
ffgZw63Ul0L8ErGudWDR8hkwSoHNuW7dezfzHDiVm1rJUkYJgkPfazZdTeT23uGt
p2aq3++LOwJioEWXcGLMpiSDh/StQqxC+2IeNeNzX3NJUngdVUWd9CCAXiM8Tsyt
+85M1Tf++mb7RrnqIbfaLl0D8OEyYU8uCjmm3As+OfsOErrBr1lFzMizDNw/UknV
um44PgqrwWr9Dpx+W/+zLnqHGGau/3sQ4SW6Mg4bGXvjx1TkD8e6qrfcy0iDQkGn
LwFo8AcOpJnrsPTAZ/c0UGa7tYHwZ4SLfsyMjBXVBAzWR2m7uoqMn3NLAjbQ8+99
TqNW6sEwc5ZpDWQ1hQfNwt58dpGsPhGkVatlMIPj0/Doj0344+XxrtSTe7Q4gq+l
ypO9mlfbH6mtbR3qvBt0fKNQeQSJs7cHIKZdi2SY/n2umikWgjoUYCH0I46G5Yii
UxsWRL0OLZpePbw+ZF4yF3brjmgrU76tsSsj+eQnel+btoSB6brEM/cfrZ5F19uK
VZMzVFcqkzwSMmt+nNV6IUm4TwQTVxMSCCxS9owI5CsyHs/1qpRTtoq/8xt1dQGS
SE5uqlHoETD8+UAPb2/tpXfiNAxYNSoHglYvhV0Xd86zaplTvBsQCiRyG8K5hNpa
HAhxruq2yErWIZSE+2nOtMuLkrBsD+nd1eBZuqtlADo/gSgGhVUfwga7/r6/8LFN
n1mqfgT1ULa74Pqkkf1ppAHq6FzwkGuwH1UmNDmi4xMCcSdAzD6zXs1N8ALAwAxX
eyb2ze6Uu6CIeRVuOSFvOQiVEgFTWqAffvFrW1QggDJu0jOJ0okxDwY8BtLEmqEU
0Er9IXIZdQyxvQ5NA41wySi7dD/YGaBoiSbFYoV8Z+YZV6bmx4wj8lylrSqJFob3
GZ96a15s0OKz7vuFcKGTyhiYIuYAU8HK/DJuNInU3xehM8yGMq/8o2jOf1SsIr7V
YLpeIllrp65lOAeazHqzocLtEB0Omc+MI+2vrmUcdh9IRlzmdhP9q0GHtjq9vU3N
OjtpRPSURJ8vUdhUEkLEy8xGkGje7XVEFvyVKA/WCo53PzJaHJlldJh2nNTnwVUK
mYnKVFsEYLVxLdqvAEuYMdf7t71ImOrXm4U7jut8ZSIaPBtt+oW8k+VV9w8dIiH1
qZOaMNMiB+TWSlzX/3BP/T89CRacZAaIeQmIcDuOZKRUUdDB0+vh4/kofgDlauiy
HCSFatbl+PKbKkR58lqHMER6BfjDov42hPYPyk9NKp9MgDSlJ/weyacH01DvnY5E
5vXWic2sKNitFMA0/KaltZX5xRr1dqHw1bpMKLl41/xE+OxXutZEisr5kJ4+PesW
pYQfrUvmeairimIP0BQjeV/um7RR9wX8qnLvZ7HAXtSWnEghriJo1/2+eKj8aHxK
KR1dCM626aJmyLYmDmAyYJS7U07eRI7Z+x5nvDK6FKYZwOWLCG69igAnXyT/x9CL
EyZ9JaEvYgIEeS3EVhZyXTO5se7g/ryBPJlx5M3ocBR0vKzFct3nmrTtB2bS0wsF
goBqTkZa3DMsoc4JJLRSdNf2IK0uULD2Pd1CilL25nKhxtBULnQ/z80s+AjIlumz
h4kDvO0FUD50eeloFEfWokhrLnkRgnNTbFs5wNtSAdjtduPO6zlpnqCvk8PpG4Yw
5vq5zrZ5FxdEOTSakHlIHLJhfLuri+7gRp8BG8ZNnWg0/ANQliuBO8NfR5LOoKbC
djhGX8dfKqylMYs6QNcGH+CL8+wVQQZucKBI8KSIRhiOP3o75MlEOB5zUJTIF8kO
2rs0FHWT7uInBYIxQSYlFpA65WISfuZVb6epkkcifzZrcB/ZZa9E9oUFNk0Gi+36
1OE0us6bHLq/xTDTf0LPHmQviKzVJFlF3rzMBB/TQs2uP0LPOWJANDuX1aYVUvfA
7us/u+fiZWgEWCRbBlwVt7Qk49vXn7LUjI0QTZUmErVKxFMCWAoXyzYVuZ8XmuC3
fklBwGMPok0i1tW3MtFjCq6Vr1u8D39osQYkQGza1J5zfIiD/HezbmDAcuJF/3wb
iqaUyayzftvNUPGVkS3rgCCA1tOZ9c4jbjGjJIyQUFovqGyrqww0ozX0maMIRQA4
o/0k8BMBEHOQn7NSxtF08eTVZOBGeqV9B8am8iZ3EltWyNBh910WkTM/l+YLR5Xm
jS3pQljggSekYKhBwOQFrwkcrH6m5JI20UAJKvf7I+Sq+BnrJXs9XUVF/7jGk+Lc
jJH6F/DbTSLEfBbheU05/9Hho6SeEy9vkk/vj0bOEVcxrbChETxlw3Y7tPTCDRf9
PUXFQQZZSSuz0JXjcWCcdoYnH6qMzj1BfiFSvzzZBDsu91FUpsgGJmwW4gwln9hM
aupKVEK4+lnm7E+ui9LYO6s30o4XthPUtNjxIahC+SM11yHs7/94hGVk2ZbSAnto
XDspBwI6jicfqnUrrd5mRatsgxyhCDAubZH+ovu6Ut923bXrD7vNZIEpwA093I+8
fJiVTReIbp45a+TQSyzePetVOXpnSeDbLcc3DbyFng5187jR641uWlwId10JNQLP
TaEELEBSLBI+71kYfzXA9ssfKH3hhz/R0P7gjnFhRm4WEFAy4Bw87NCZIHxuZvHy
WvKTq3wON/O2xPZEUrAqstxOJ1CVuLLo/8GcfrEErsnC0MPOxh6gTamaIphv279L
Z1CZcHQOX0kluVBfeHEAv8l057A5wgKJkYrKU6JQyZUx7dFGSwBFiCqVNJ+s08I2
WD5SUq1NKz6cCxtvRYnYOYene8VndteRlJtj07gZAw3GxUAYZeK+z9sMWUykTbRe
FT1gaNVSx6bLPJ4utS7N1d/VfjD+H7Ss/sUN3+HdEWDsZVp9YWXTtij/7B/XXKDw
FtzgxfJO6g1Ez8ZcgPgXszEEIJSNLHJluEGiglagmFSPnIh4n48gAOil0fbkgcLj
TowFwnitfKfVNbBuM6tr5lBgoC7bRR1VKQZf7yJyr1zxzmL7GPh8yLqga1qafvEa
0qe1M1Y9MGuS89N+Teyz5+H+P4oqaUqrbUNY3sHHvs8/WgAF1R5XsjipOnRXilRz
Z7mUDPhY5qQkx7Qz+DJ/sFmjjNlY8edfgaOiJQwUcb9+bxi7cZLjNHt6KbC2VP9h
wy8CrlrWG6ydEgbAN+OYjx73tu5sbUAXIUOUsXU5Mmx40Qb+0hdNzGJq480Agzk/
v1/Hu72G7rlk3kR+nVZ/HWSNqr8/I62aGQoQrgbzW9SWBF6pNrAkmt5DW8Uunfdp
v3C6z8yfC6lzv/RpTt6j0fTMkcyXYWMXn4Y0ZR/8juAcrFjFla4iM4tQG6TfoMHh
9FiGkzE4DYBTVqaYeT/HFEqqKN9Yz5cut+d9BJ+88a8=
`pragma protect end_protected
