// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
OCAZpiSkCffP3tIw8f4hkhu7lLBoUYW3+TYBWSh5hYjxj1DeHl8sVbtYuvOD7mxjbvtznHPcsCLQ
g2UfMT5sM7JLaSuVqHVTOjLv4rUp1YJeMdkMe1GuL7SO/Uisgav4pwlFiRmLTChLX15/HYFPs+4V
q2hjRjjSiRk93LNYkEd/T96i110eDr49uihIUJhnXLxfgvtr+p3FcPM80HSWxfrhrCNUi+W0cjFa
lwVdw9+Roy/5LhXxPPD1dLbdsp5C8AXxN5zyYLTcMtYiWPosjXjgn06NrrVx/tqxDOknj5azcsao
pP6o7B2w5/CRs8ztPN43jFbLrTA/ThM3dJhzHw==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
MAhJiotWwvlPVegRGPlYNdGyPN1x98MeuhOyP3jbCqC1OMt1EWOrW9vh6aTHCSuvv+fRBlQ8eDbF
NIPAPei1Ln4XBHRFB7MZyDZnHO+ecXbUVabRdawAX+yKwzSfKZ4pinBz9mz6+Ml6h7kiC53twtcJ
uuPtKx6mBeuUYnR9QV5tg1+g2urQPKTuZRVCWbvBhgP8Hzxq621drVxIkD2X8vpvKm+sfWV++dfr
EcFfi2toivNTupWxuer48K8w6BZTJEuvH5QDph0m057RBpoXFtJ3RZkcL7UeqyDQXSANuepy0wgg
e88J6VPwH3GGp2pKC7XGKitXLZts+xs612ukNG2hZlFT0pUHuI4nZMDMJ7/VLy9jm4poFtOvBOQQ
csiiVVy3FydGg30BWx1Vj5/X9OlsM913CC2c0P3pXOV1HlxkF9v0RkmgL86H66kBKkpFEg67dUfQ
6zrElKg7tR/iC3Ke6My0tep8bhepSvKDhK7nxM26WSzhHFMn1rR1xIu/ecA6jHJaEj4jsktaVX7U
NK2zJlOaNQP1Dv9ADSTKFuiVJ9oVb73i8RJ682Po62f47xxoOCDR932bFxvYc8MgDzFcPfmDp/Kq
Lk5pa96DsGlKw/9VTMaSYX2HVhu8hR49YMDQERYhtewuFOBIFhG3x90wVn+CidRGFkPBcAdmNq7w
5wisTCTXVWkYDNbB40i1B46OKPxoLjMvuM/D77HB4yRIArqe/cy50/wroXMm4+uTSWNCZru/xzpi
qxiEP35Krs8uDjF6gWNgyJ1MKNnkeuMpenatBOdK/cpWxbyNqI09dpzo+IW1HBmTKMAqFyNNrwDb
+xx/uONlFxLGQV+Yf24Cg1NAHBFrD0K1zxdq86sDRoEROIsKJZ51UZT/vtcC+bkv96pHJIUNr5Q8
klHSv5HfC6F6tZIfinfDNSFa0dYJEFbjPTruyKih3IDG+yCK/TLXMIL6FQzp6bEGcl3/3+Ip0Ui7
8RVisEvm0mVsc2Qd+aFAdCJqYFaXwjHauGwMyk0Brw4gIqG4TYUQCLTAYf/ztOaHYBTtUbK1IOFL
KgCclivb6DOWsvYs4qtPB6CZfeRIU9ndUepluEByxRPVPKKdAZiJg4D8zYJfiINbrIvi8td0UMM7
p8ru1C2jLtRzFFiaRVMy+HqyME4DVM1P3wPSNMdJFU1PvDMo6BowC/LM1LT+JOBJpLuGM22Q1YED
wviGtw34/0lis79NTlDydc3TNDb9uH/0xVk+e9ZP4jbBCPztUv23W6ry/k5DtDEGX6yJTbJZZlOm
hsRizxrUtrWm4w1dwOGHDR0e4FqwqIo1MJpRlOKbXSoZzXr2G0LRjOGf+VjJC445VxLipcoyW016
bWrbiWFR0JnSWGgJYGOoWnCTXKJB53GlV4f4DbpQsYxr1CFu7H27W4j0zkeJcy5kFFrK+GrpNxz1
CQPz7ltvGsuUAqTYBGLLzkVmK546mc7yRIPQ323PCDIpvuqEeSp1AycAui+qG9jjMGO/Qs+hpH7c
PIRsg66p6USGOj7909RbSbgVbheg4uqmtPPxnkQ29iHOv/97Vxj29NYj72XuI04tA4acq3/KTybI
XOAl3VtGtfSz1hfTVBy0y8CoJGR91HtW/NNnA8j7E8sPUmwfBO3PcIgf7oonYoYLrePQzhzkpG94
FIVgIeObrZ/KvfJ30EYYmuXVPIGt7f9K62GCfidghC8u52w9Au0XXjREEupLZQoZUPGDx4OakhrC
YfYQs+ACffBZaRVo+BNI/jA4aGraheP0v61aHowBZM+fEm5UX3zi30I9V+OR7PurjSkXPtksyaRK
/d3iTczUga6rLCrrxi7+i95eR6ZQFpF7tpw8vCfv/omsIQh39gUVQEAdRE6Sn9UB/cDovSmZ621q
G/6onUc8MLIokIGwiFcHtdRgCc1SBSNxiXcAImuVfcLmFU8VWUrLOuxmFW1abPI0SzXisVC7pCPx
g3wgTtS8rxNRzB0zVrbA+qmLBt+lCigmC9t8CXcOmXSKSkXH8MZOWlEZnZVtRxwCQ6a34svFaX10
Fpa0YpiGxMFLad5W+FD/XPMWZ3aAD8lRRjaNnhJl0ogwDAwPvd+jpTo+6+xrWGwWToXJVe/o4PR7
VBQjh1rfeClwj5Usvbj/vrxeWDOml7c3tMG5FbZEQ7cdBmheIg+cbi5/UF2MsJKvaY5hON5W0r5z
KFChBEk3t9uxyaLwjoXtA9Uu72knqqhXQU/W8GlQoG8p/Yyeya0+Bxw+rcxjyZNbjZbY+1sHRVWC
TdZbRrIlSG4rR+3xNh/pYnxdmFbfbkO+9lI4YFuQFvwsnKiqmRGzD1MR7uFjcpyQ3W/9CVL/pwkl
uiy7rr1DgCdxUmaW/1OsSZmypHruevQ+AEOeeoDI1DaJNdmbUFNsaBycXeKrOzaH9Qn69XXlFHTG
mea8e4/x9gLgyqsoxTlsxMOAhOd5SWR0Ga5YRrfX7VBaVj1ojJAhyfMrZWBql5A+/mTnykimZUcD
I58brKbiWmNyBX7PE+pmyeF+RMnBdRnCYXqfq8LRDipSv9IyL0uRI6TK2+30DlvJkYLen742Szi1
P6AEra0BOcJAx0D5EC9CilEfcWhZi9EMo+weOAt6IJtwRjf16pRRsiwrlpVVJEEy5Y38IkUwQ3/2
LgzDrBLWP/uY2ikaf0qCplwNqZ0YV2XRZ6hwRxviPqMSQ/xByQKssa5V6wQO5lZ0GmKkqBVRi88t
60NPzQfGvjGxnoyxN7KJi2O3quFi2lI9LiwGUrtEpaOs+vEKLH1nT7jzHgC8A6SUufEInYJ+4Aux
rdFmbYmvsvWEXgEd+jeuw3olUZ0AruFZhpXmBYcj0NpvlhYaecRySPSWujCmivwmR9W8bsFLG0Ic
KLKhpkxNhU6uchcrZzF876aOX+Bp4e3An3uTvRqUz/22h3LI30EXs2LyW9L6R0I+xrYzsaAZ6Ji0
rLfdWcbaJarULUDEC1x/sLYIdq4ZLUKfnsZYT5AuDi+y0LcQXpcBzHh47kgzNPwBEi18vba/19qa
G6I4Lx7DmunVqLWyTpCOnvHgslMtv3EWJbiyLjdomrVQzdWAU/Bty5l90eTiuIRsnK+gB9kuuCfh
ytb3AKYPloehdnpytTkXhS1g1bFAbQZ4qY34NgJcvBimtFq1WLsQXe9LftIHLuZKgqzRCV8LVyrL
YM1UeR43CqTAFYePlC+mAF+FGXekKYOdjyJzusxK6XVFLNjizNsihkuwsdwknpZBMhoQ6AqfDNL3
PeRgyaUG+vrwWfMtfRToFcJOWo8C5Ee0nQM0WztDYbmh5KfKCv/BY/4oVOn8YAX5vFdtT2z+rIBC
5igEBV+4bo4Sw44ThaIu2DwDkMFBMOc4T993wAKf+OIgFCitDVGUwVskwJxFLyWWjS0ZmQb/EgUV
u24/j/8d+0t73ZvDmu2irF0aPRF59VzbqBFk6w3CZ0nJM8Y1NRmPXSupnyB4Rf8SDx2aqmrUoECu
jSFA7Jx5xgUW6Z5ht9fjILkEEf5FgSpHc2tNK7COJCFrVqXMpoJ3jVfoshn1kalWo04h7SgZCQI5
WExow9iy6vKvjMUGuYy3b3XmS4RXtYrvQgSz4NYYSZ6HESJbKC/AmDIfIpjTPeRBKDlM7KBUhXFw
2qCWOwoAe+wdLJGb7mpnz433AtO1wcvmCFuRP2gHBJZsVi9UORDuLd50yydeMDa6DdRaMh4L4FBE
gVdhiJZ1HMg09jDCM/V3uQoZMHMwPUAkVqHz3eR3efXjKT8ivgXZZZAi1cAPKysdsTbLQRmGwXIn
o0TzdBx6GLXwk4h/HgmFkGwayZ6UpHGAomVZrhJb3hWLOHZcHBpU0+Nd11JVm3WxzL4uYwXKoo/e
zdD6ziOGeB9okcZWjPrHX30mZNmmQvC08u5HNVI+KhHcwYzIjpF0obyI9cgLnlLuFME2pSU5vF1Z
OcMNDoQ5ZxXRulSJQSjCU3teCrdmXqxbgwPNXaNp+NdmaNUQ6GDTPCqHjdvFDeejKMKWf8nxHVU3
y1HIppArSuW20OaZgWinYJAUfoybiLTZ0TT12Aa4ZoxdqCqkW3XPI9XutvjVWRUbzod5ZGVuIg/g
my5M4fMXS3nVqb4+K8vWovIDZIv9ZSeizwBlZkj9UZuV5Eg/yE1btFQZZ+satKtxPRXgtb40IgmZ
3QnHp5M75hOj//oYnDbgdtu4tky3SfikAavbCaUCvr9x02kSOE5x3iYy+t+w0/ae8+mUuEN0ml8v
Nd0zn5E4fDXlnfpfzfNz4OFX0WIYE1NQ6GAAv53/VosMP1d5zpn7/wrChEEbwoUrEwSwAuWnx8PS
uYh64zmkshhFeBOORXdcLX62CcRvrYJLC3xB1waEw4Oy6859eFHb+uENnTMEp8sWXfXf89hYHlEL
gnK415+YuW/xWgJYnSakjxR3fwQC1peimffR8sxS+oRHjFy5RyY+3RtaoTTqXr+RnNaIyuu32f0+
MFYJOoREbpOCaoreGFI41Be+Kqx5N7oz0nRv8PfRS+lag1qmhLA4hFGgzA9c+FlqRkE/1SEvDL/d
mI1sF+CB2+dRmqCshwlS8GFLgV4FvF3oZSbxRVn9T8hCKYVdp8zHBDZq1cqVpPCijh9yfZum8cDY
yo3ztxTyhBwImDlneCKjhNTMQBtEbwuJvKmVcNVRhwSBOOkAoiGNXiJcbMLpxYLvhU0jAVx2GRzW
9cm6y9LEczkFPgySgE6RcNaq6PXwkfhoEACGys8x9RHN3sf6oST+CqKzsF5hwHf+6phiFP/Uh6K2
IQDyG5tIXZ9bm0AncRyJ+AdfkYhrOaX6D+B6kQi8dhCN5lNNnlX4Tys/IPxzE9alocxKmVPMS5WZ
JsHNUqnEMxEPg4SlB/E8wjI9AN9YfNv/rYYq5aj5boMHSXNgU46X/b1ESE85crHHeLQERgzsqkrv
6DE32OeNsGkDMUSri2GMrLIgGwFF6un0its8iymVLhag+cb2BZaeCLQxHtNAHqiq171R0nvvYgFB
3On8PaT/bph33g2cSwbZMpHidgrFxgkAK7+hF/j6d5IqP6VrqlFD0FPbVYSb8vTTyLutUQjuMixp
xrhykNCJwqWxIpA22Wlt++MuyWIIPrfIWRQf1rZmp/lWg+xM+yI4LdgiD+S8ykhWODYuOYZAxWiL
6sQsj6+3Ao3pMhh5It6DRk9CADMU99EeiOdCYUIOkXmKt1F+mY8148SUH+1vnEitrA+uJyAIa0hV
jkJSrZ+u/k1xl14+LYLhm5QW4QbBtFSb2MQqQ12cJ2SRx7kYwCLChhU2x1tQkzjT0IBhj/UXRyoK
Y/1zMR0KG36hxo9Q6Q736jJAY+g3Yf1vPPhVylO6s3GaJIiX4oSfsILgxopOxzEOCghTxrEFnEyK
LYH3VS78d5EHuoHjJqMsHLTrPNkJm2smfXfxYYBSd/IKFLKiNhThxDpuMh8CvuymosZ9/8bdLW5u
iDvnvYi7Mndf0rMVSzrwc8AVOKmwa/YOzSaOgg7D93cQhL7C1L+jmscvE3+fVvRfmUKIwM5eyBuf
3rFV5T5UuLWDYuwHYpqdMer7+fxxscB1EWnTB3QxmXoOGy1jQqJFx8Op0H87T8WWxF7vXvTyWgAX
HCRppc5M2qCo3axl41B9Lwl2AlyPQDW7BJFeBY4kJQAuM4TUiUN08c9lYTKbH09sFTsoJ76W86du
Rk7ZvFBeVJSUB1yRbSWJvmOH89FQQFdB/7erbTG6diTpPvXnWMyRmyy11p5pz0U8uHqDz4x8a23v
6ee8C5YSAZtqyRMud0fWjXJ0AaDBkrn8J3o+yt/3QJbrYcI/qYWkRjo+ni2WsU3gh3JELWLif8P/
ALXoZSl7n/4IU8uWe9Y6iDaOCzawV3p7LtpNHEveM+gcNvXoHOHTWa+VkZVjjWDBifp/5pLVhEa6
L26V4XcwWMAGElu4x31X+1RdITquxhzQ6gVPkJsPBRVt5y6Qt7ei04+9BRKBbcSCd7uAev3ZJtPY
Kpuk/OUiOB6Zdd5kOiVWxHM9ugfprSZBRA/+ofaCKi2YeI4ltF4EpjruxOTjjViDJEreVIoY+/Do
9ImS60ouMLDATCMP/txTPNshwqdFpdWNKN3FRM+gw9qihl3NeAJAZnykHQ3ce6BK2nXV0gyvZnt6
u3gOnsFlQdJ4/Dpf25FK0tP3YRYvEFjZ0RXNFG9YsvIJ/eiuB1dFBnxafSqMewjlPDr+QE2xywWg
Dsvd6/TVX+0hLi2HMYJnmvQg+cRRH43cZcBkKObCvaq8p8nRiK+XIlpjdzeeSJntQJW07Is4cMeW
5jPLr4tFnpeG91t8TP1Ws8zlKOPzKYdJ8sePnFZ1e2n/V9z7kooHpwrEpHM7FRLiLzmUw1cfcYqA
+w2SDASFpg4EqtXwuR1IRWvbtUcpmKSj+jrpHeMKlMPFtZBAWCMbT4dAn8a0uaS22JnBfEvKDSDG
GeGXJ6UHfavtPrQKUa15SO5y+GmqQFgP4Nf7qz2ULfqlpNi8jKFhsp4cKcby4s0cIp54oGjR1IJ2
7LSaou5txywhvxJ4OSHPDCiquGRTft/njZQh1j7apIbhao2u6CtbQ9QA3zfpooCIOPAMKkBQM8VE
tUJ1OROhKR40cJ0tzBA/ceMZX/XTPYvqs7WcVLwDlTenHMquB13bMKX0Oii3kkKpbLcIOn1Pd+6v
lKoaTR+0m+4YpKhxI9FFJ9wGkeTG8PV7oEftr8K+GYvzXSOUpWCH1/9FBLBX0Kd7IFpKtbY+O4Hn
EQPg+luSG2aNIdiblMW46+mojExJXt/P2eBTAoNgochNJT/AABB2L0KMRCzicCfcJ7lrjw53it94
XAlQXb2S8JmiJ+E4ej+vYiXBtzgJhTAAcZcs9K47zR5Cqt5L5lJT/4gtuoD39EVikh/6YQJkJyd3
yfPFLdsGz8XjPuKSy2a+Nvz5igTEHHwJ1RkYvz5qVB+/EkUSSTvnq0AGrboV2eXZKB/lzLjuumkt
affRTWNc/D1MLIQNRctOdf5TJmt2dnKGIFXEInMeTGoE3ISsRdub4m66GOIRTOpbdzims4C5AaP6
Hr30QdjMPmHzSO9ocSiAuBkdrCfCNvc50ENbcSggM8PoBeHdO/r6J3YzimNP7K2NvXl3yadSg2Wn
OAdx3mngyGvE0BfHyh7AIi3BXCJBbE5TDMimoTT6D9iATb5f8DRFoZt0Xnh8PFOa0/Odvs+h6oex
GNJNGv9n7+459/C5HlChdV7rHiiDBsTzLKBfkgOgIpcV8vLPirQH+rFKL2eoFar1xVKZSR1ulFhq
WNHnCVa6k5U6aaw7JQCTkCv2XnSB6x7iWzflAUnWzKzRVvIxU+bXoXksxkcIq7ws8XWkA3d8gDWF
fOQf2Fg3qmTeShm0ZM3K4JGPsHvhY+/hxGoc3CW46rPlxprZcT5RTlKGtLa/JHg5qsbgJ6zS+aOq
opFwIlMfzI+MeC6i2aGL7In6QOyHfANNxfc6Ic5texp9iySf8sCdlfIEOnN9Jyrn/bWUNHf3ghO6
671rE7ZkSq8PiB/XM1qMaC0U5Vglk0Q2ppK7bozOuRoEEFKTLGjoPTEP1VvXeI1sP6MrlaLM6zZi
LUU/yFNgUx6XWp5q9xd8hfLGLNqWzuw/B3fOyJDsx4TWzbpflxNtNNaFpvd4daap4SFEE7i8Q/sK
kAof5dNiA2LRaSLK1lj17A7avFdWueQb8JR9bcKCzs8ME+adnX5UNChlAYoZU+RhjJhMyKIhcdLR
13sU7ozZULsijgGoQca/6ekA5ukqEUAN81QqXNSn+hpe6Cna8Zavp3Oht1n7Jzcoi/YlM203cFvT
woCMw+2yjznncOi3Mgfbvwql4/5FpWD1wGrBvIfk/z6cqzwAifHyx8mFQLmU+dB1kw5+dprm4lF9
xtgNQd0Qyt6mALvuANRk6UsTHdnYP71o36hPtXlH5iEa4AiU8KUp+Wcbh24sJ0z/PRZcSpG0FYMs
KRaPxxv+j3NOLQdbEZpB3dGniS5wQqekECUF1srXfwToLKWnmpA/XbRvqpNDQ/zHCv/vd+HQPgqT
XaEtN0ogL4Wff+OckxSnmuRSwhC/Cnm0n4g8iokCczuj8R0r+toRbipepJDr9HM3BJh1UIFMaX0J
gwY9Uet9yR3REFy6hWXcpfkOQ2p8tF5+enxmQ5P6GfoiXdT2Vj266Aabpb6sSV/HM4Qs05P0CU+p
lZaq7LU6ApRCnbwaqmkmO8AVcTOAZdtEpzC76dMq59qNKDMdCNURCOjPCqDBJjeZBguFOlndWgLw
DjYHyl+Q+Hn5JyIMsLcq33qYkG5PvGsdDHN8NZCSg+jtKGrcczDCMu/NjzBq2cviLt82To/WrI7u
H1hSc5O57CsMF3NndDiR/7LjInDV9Rm1DfWmogJEcmuDnp2Z3eQ+ivCOfmhhuZ5rPL6x1XJV5R7Y
n2m2DBZQA6rEO4VKebhBB5Qiyo3z+JLivam2hMKbF17g46mdVs1bT9e3wd0NIqwmK5+KfyqBSDyu
euFmstEoDe+Y43j6ObsDlMmg5hLOG1Hg6RH4S2WvYKjtBqubfKXYrWJGiynxsVymE2nlvyIFr/TW
pi1FaYz/xtgJ8BRZJj+NepwFG09k343GREENyCe5Y8W12KcA2HPnO/pIW70wULEnvXjsZuoZJXTO
csYGiVo9fYQBJAT2AeJK4ax/MfDUodIXrAIUj2DNh+Bv8OzwNoXzegbUht/3Qm/MdRXNzkwhSfZZ
WjhpTdtXZXYCqD2N4Y3jB1oWUN2f7ljgWFCS/0sW2GKNwNlKsCutdLbSS6NlHOBAIj0atqdSeNXK
AXNpawJTAkLl5xXmdm7JFa7MqTTBXp2m/z+9H3b7DKNUdCmKUMIKdvqS8AnevFWJN4GNKeKjhjc5
ZXAFzRwNV/rReQ4+9FF2cbofCQ6YmS80HaXfmre+H78Own7Ypaz4fXYCWlhBA/RVzB5EeYT1jXbw
5iyG4EyBILRLr8C9iayb4a9jjgBCxHTqndmvfO4iAIuR/eASP/IxxTU+YDibxgO7GJYb+oReK3e7
Rlf3Q81lQYb9u2zo2zZ+wqh2yx74OyOOcZXU4yE1OXsH+L27Vg39R2VWc0Q2kfYggVe4+UrqyEAq
f7LQtMjfWAvG7Q/+cROrKhIAPQ/NJ8ToE0l3Aoeb04yzzDKGsjL1Zj83zkkAxn/Zd6cIb1fWnc4e
ZO8UsmblLxDKreRGZ2AjZpVNSa1EUDDvi8ADvM8KoU24WxtyqPdyPX0srCPfCNVNoBtRCd8b5WT/
fMxolHdmZRe+LmeGTgQu2op6VuecXHvIdN2+UIm2qcKOZojNY8r8KCkqA6XRbQzQwH/Ff4ebdIQh
RX+ABsks312T/3i+6bvpJQlfT2MSc6ed+joxoBb0BbQcgeAdBi5kht4KlFkjoOWnsir2OJTU0DA4
Y7qHj8s3ZHzRfIVBl/4BWxogK2Ad0kMpVqtuuwzxF7qwZmOhIw8qOP9brM6jfiXuGN8yQLVK/e4q
x9cJNOzHu0coZnYAFS3PNqa3C0wjSSSkKrM/Xe0jy09ZvT4TAaJirAV4eNdlNPKy9sLwQQ6Fgdms
kK6aMAjCCFRaf545duSybble6HDi6cmEbiGCTT0AthnQkXiEqWcNddVC37EBM+JFYTi0eZy5PYuQ
WbU9bep+KDoUDFlh5Ubkqvb0p5rimxulInIr8V5BwwsT4YGzqyy4Fsgxe+qlhptVmSXk57MSPCC5
/6TBTX0M0O7SqsxgnHMTckjtmktzoQClOu80C9T0tT+OvqCY2GBixgeUKVKfs11qxXeAQ9eKATqu
xQZh1Z3OjldzF3pqq4kF2nRFvl3Xh5bXpnuV2nBqf6/6SAW+pmMeXihB3RSnCdD6Hmjwoht4jnyr
cWm0Xh6Ygb7RBEZ1bWNHCNneGZxrGWxmvGI+b88tQkkwJiGmRbhjbhwK/l/4FFRpzbmz1v5vNGXw
ggRTYGd9SqTxhIL0ly1XdpVKfrAOUZrv1exasuffz0Htsj3Gi4rrzCAeHs10dJw0PLNpOcae+Myf
2sZ5p0dotEfQZfLWgliGfl5HWxtq5EHCoETe2IFSZh85Ih2I6VxZ6AjtZ/Ild4WGlk5JCL42aqEj
aZqY05NAQe2JGh1jzOJyQ6wkIMyhBKVkHOokhqvA9NPPzXVYkw1gZnIkPuZWZc7mIrV7PrzomF3H
EwUx9RVQWh3hCJmA0moAUI8J4xitzK6JVHo/JhO9oInXF9YYvJKSRDJaPv0/k0qVe7fwCCF6pZtP
BwFYS9DxyPG3Gkj3nm4LreOilc39kKL79XgjrACGu3NUXelel8L1c4wVhKGURmDZs90FwRfnc9SC
QiMkupqNq5YxXYaTG5s7BIsW32mWYE7WjjnP/RMKw/L/cbx0eOHI8PFtyd0p0bu5t/eVdgNpec3w
Grxyiond/Uf0+06BIjfHuL02UPzv6gFEpnPEq2io+UOV6lpTaGxBP6l68zfvxPL0qJh4sC9HFP3Y
iW9IY0qChP0FDCmm7Xjmd6CaJeSp3UiMSisxKznI6Y5dFEACjPYnoho/fXNW9t5U0TdbdLhf7wqD
LSX9cwBWMGcVRhEMRnDSsW+O3xP8ZNZ8eoVF5z394zu86+iZNT7rzoIj2jzlFBvJ6y1ZhJyYrlpA
x6AnqLixuRvOEuZkdG7cTDbt4JmUwNku8/AxbKI0SyBYQbMmpxtUFh0Qq8nVZunSiADo6j0s8Bow
zJ2PDWTWMYTfT2bpF+yuNtX4DStDVHuJNAjNOqgmiQl3Q0EkhwVa+RttqzTmh+a1+r3JBGzGWkMF
W9el45Ls6Gs/eyDb05fKr71C2UVOk3GIqH6WddAj4uYu284442Z/LvrUNUevrsr3ozDeswBMEUVW
yWnrcnaLMkZGiij87+GPc4ZANGzhv9nsHwEtzpjxV5lORt2NBQADdi//VwNQw9LbBbC8s49LWZKA
kpbmVV40wPnSzq1gyfLbuNl044oWuibkaNHBDeaGiVp2kZkLcH6ywJNP2xhU0CwR0B37n0c9S90W
4REE4ac1sbmT8IRNnj4AfibBUeyvw9ggwtae95oTqzmX3oY8ompqCPCf0EU/7gF72kyf9heyjOgY
v8+OphlyEX3QApkzDheunYLpLZwa0kG3lWcJYoVm2L8WzwAkt++xWagsZPUW/CaLI1swDwNK3xFD
0r7mZQws+6bg61PEUT5XCb3BUrdDpkNbmxP5kpz4axdloP0SLGEfLDSDK+4YwfMB9+gy1E26NUOm
3rW4eLIO/1Yha/1WUJmA/C8A1WP3E1sSNSzc1urBLooPrMTUmjZeciAj56U6HqvyBIEB12hdgR4z
w4zwZ+2O46wu4Kby9N2s/Bm1EfXgkMPNo+Yw0XrQVt7UyZzYYm/TrmP8DZbaYu4w79aQpeR4vzDe
UiGOqeHDkqdyEtigDJ3spy6dFvZL9sRC2NbdIBl+dsO2FjOfBPNjHHglN8Ak/BEaTzpH4rF5nbVp
8am0C+McNLLculoH91oUZi4VrTvmT30OP/QzpG3EWVGfOZtzMBPq7gOXNGqYGvfMGKGd2JroIBWy
cvacPJU4BjJG2eeXh1PWSK2fXuUKRUQB0Q6CQcOzyZGx17B60pk9ckDz/6QB9eH2FupTsJkmzxGU
2LyPmkOdrSZcq3Teq0bF6uZX0seGomLJXSAMkFGgt63OYggd4P3Zf0Whg961H/gR3dmnSEoAzpyz
qjQYV4OQhuIII2Rp5XUvo08WpeGqynr5JUWNaov7TZEcH/sSuwpswvsG6bWXaBE8eQ5S/7AEq5qE
lM+dX88c1BSukFugg6epTl15Wx5e9eGP1uC3HgbxukLj2t1czv3MjPIorYFTThH4t56X2hTzGDVs
JCWr9EI6iQZ+/vRMIjyoPQlX+2rHdUF3rg0W9/Wl5W+qpCFv8YKqBkRVdJd+BwqUMeuE7/wmTvGh
x/mWI8Qc+6n9FKzZ3HCoWjmY0pL/B+S5voABaTiZ9rWAivhb/QrjGBaJ6hcNmgLULp585ts8cpM4
7FAWvxTj9g6ZAGxk7xUVkQgPCfR2cvT1ivjBSjsK3L2hAYAHNh0dHbOhIG6dGm5wUS8db4vYyVLC
nJceueLXC9P3KGPt+3jFrqUYsJQGle6uGXcN9TpLRYYNWwhCAer02+9vo57FwTzTPF8uc0pDj/WE
Gnx9YtAivk26SzU+qtt4fbKCoTlBT17IBEeIouTrgnCQn/7an5R+hq/vRXEXPj1TasWk8kDRa6Bv
HuaBCszxVRPP8aooZsb4XI+JQ6dMwPmYdtRJzWrxTiccYrxXSY1Puz+V7Xcgvi47ZNMJkWlexXLI
mCMWOAEXqN72AVaiAo1BYe2lhU6s3v+QmEy6FB3tk2A34MBLyMuisiB11Ofph4ORaFLDOjVamjqm
tAGvg4t2XmCMqjdw1zkCzdp1FznWuc+/vMuJZQgSqQ6KZixszBKha1YrFSycLTO8oJ2KwsjcTw1W
WBj00DR+jyukRFCb/+/Sa2gRKjvKoG2KXXLSQUuT4uJzz1VyJDOmNj4X23xIdOqtHAbcT3GZg54e
zItKM7UTXfR0LniVc5z7eW5JatOidn9QnP98MMcj3J/Y4fB3CvTsBYJMjj2rmK20TC5mJHWndj1P
jEVM/oMx6T9LdI2oW5oYq3kwQDS/ehmZgs7mHC0LnQqp86edvBarsCQlhNO19CKEgHKEUJPzxO2n
Oitze3cJJOEx6LYHuzFwS6a2fZMsw5nf/qzixrYExFTAn09MewMISyWrwB+0mjZsCmbyuQfsg5Po
DGrNlnZ6wOlyIF2nuD4YQkNGUHD0y74yi2VsKMGizFFSS4Of2onHoda4Mmy5ofDFL66t61zZhdD2
8NSWp+5pMPObdElVh1T0dJWMlZG04muFfPDOo2V63xsowlMbC1mk41d3FAF8Nm80klBRrCzk8vac
1F+kFBlIa3Dxodq1rt47f6i4xR+QqTV1qCpxiTJ4h42Mbty7UhdRW0yYNSzVYQdI+0KWMAvIZ8SZ
hrk3DlV37os2nNJx5i70Salo7RUAk4IwWQuLl3Zkt1CuNfuonx3i9mydkxjvERBA0xggLYCdLp1t
8dOb3vvR1c5AaXjT0zB1T1ZjXlms9obd9s/UB4qTjBst8tdP7O1Kq7MZWXAL6PzlSXx6Suq9ihsk
22W8J6dJTum12+Qb2M4509VpurTfacL2OpLCxbU18T1rTia/gwHJjw7Krzjm3lDPBYCjtSEwWctY
bRPkxJol4oFQDqIXOHNoP0oDrZVyJoDISIdufemBepSoP06BjgQAkiYJWZqUwDysII0rzLMD3Eyz
o7tSZyBv68aCu7WuRli6blCLLbKCdVCtXnne78LOeGzDS0rGc+M0lO9OR3slFfB4kljZleL/D19u
Fhxv8ld/TM1fXM58OgTJ3bm3yFPzUVatCDpXxcicj08maT0YBjWYaJKPRxS45Vc6AWAh62ZI91wz
8OW1PbRLsQ8G3FNPAKFdQPV/JTNYwVKLoBqFxL2479AVs6qOl83ADdWk9RvnQFxyvC/FJLRn72ce
AXWkec0JW8Bbx7k3fR3+4A+lvjKHpNh34i/1bZLxLSXez8rkm9tizseZk8HLcTg80BZWPHw4gjrC
UTn6zGO3oVvAk18bBqLq4OIcmNsa2FqTlZ89+uMZ5B9JuD1HCDIMrVGELoFizqb5oELMhFeNpkuP
dF0wkdjNTdkMzqYvgzI7zWfZFx7wr7AV/K5bTBImDi0DDPwEmU6eLOqmj5vWRmhZFQDrZ1JPl+P1
0s1eW7Yx2XdnCVvSqbjSrElBa56EhGUY4scirGR6cYNrMgRyIu+3ATN0Iy/SzNCPRfsycW9z5qoy
sNEcvWp6vkdK5nOaNTne3YfxHAxpwwQF2pHiHe52ii49WaJ3r57c+Z77iUl4x6qtOJg2ntuo/aqh
jF0xxrM8GwmiU6QU8zfW7znmtXmcK+0tVBEqa+i6iBRc+ixWvUujJmfnJT3bOs9h4otOnHL4/bFl
GavD9YkP2foDT49yNy+JuHez+rNkW+DIAqxwb2eHQK95nQD5NfDx28bgx+z8cLh78js0+s32SbpP
2B7+dDZI+9RaADPqvb/CbTmWK7OAyrlIchxgO1pQZ8GfcjXipSRFSn4XJypvoZtTDiTPwM+QjegY
QkkZhFqzOuglIjv59RYhMsj0v7a92YIrnfrlhhIC0MIjpohjUT8UqgxglwqwXMF2+1/6e0Aasjg5
sdRb9h7nmv+gQUA8OWVBNB4fmxOrQ4mveLdMSsi/IYTYnL+a0QOE6y1GE5osv7tG9647VAYTVWA6
74ihCIrD4tNGTKwtitQKGuVaSzVkEp9R/9jjPy6s0ylhIFOd1d5CgeGLLL1Pg2GR2N0RZNkGhO+z
4zbEAFVUvkRq4GlOMNZ58zjtk+IZn0i4COC8K3nwynN5V/GowPJQsaRR5NPUPR+jT9xaRhBUQ7en
97wZl3+U2cyO4LV4v7wc6jmTF3AhkJHaWvO315WtD5NhlgVzFLDA87UFcVBHJEQdvSqD7FJkbI4l
+Fu1vYpV4U258/BuguDLYFzGlrK2avfSkqi2wJ94mDx8sV1q1ye8fvLgKwSxFmrLh6aT3P+7L46+
a6KMrWlVtuQqM+ba1MUJSMi0UdIlJ9pB1sqy84nnYyfR/aIx2jqJDWSxIP4YBS8lkWQ7oZEok0Pb
UJPZmj9cZqpTC7HEey/mpxUvnz3y3gl71ruocgL+VjHOffl1bp7y585xbFKM5Yk/H79p22aaZmm1
Lu7VdamyQUhcbwC21sqV5v7YirYUr5n637mFgBQc1d6dAqrqdpTwqkQMXMXBwYMGyrIiRYZoj8oQ
XO6/+VpxRVuJPwbmUKfFAOTsSWGtgCcORM5AwfUQN5oRz/2u6EBVvTDLVPqbinN538OLwigDa507
LFrlqAv5jUg0lRHd2Eh7PBVuEprHwoJznAT9LS6+Z1ZnKm8EBkOlnHUI5oli1xb4YEguQnfsimyu
jz96VPVUyIglJMqa8bmCaRcrjhq6lVs7lvXKygatwrw1fGvW3Z4TKhX+N+CEn/EotRGGWHJQ2tMM
cQO6ALvAUAWN5a756gIVXf9VTO94uU4ZrWBUb48c9pC1DAYid33AdM/4GXHVhCvFmHSDegeXKDLj
6JHgsmThTgIGuESEHv1r5XaPSUvcFVLrYX82JblRg1+MFGiDD+kh2789vgVg9mIIjHAlFCcQreIq
VbjhyA2zT5SrDfoQ5SvkYqTqgc1I+uI18pRr1nzuHudlAmZqb7fV1AaoR1srRNkYJKnkTrB9efa0
qi/7Ti4vsaX7Wj6um8+KZJskM/VLXHLRof6/FEyTXa6S/AMGk+IwvAVyFSqiTaD2QXeGhKhqu4GY
iXDnfZPP79m/z0BfpsFtPt3E8Moju1lpc3CPVRjDxoILhTxsvrHkZajRAydqvULRCPGPLL/kczym
+seazoJCYs+kWf6OrfI3zJ8nOpXFcaYJj5Ytl6A6Sy/R6etWkiaF048COO4RavTtmlQ3atgzBMWj
nDqvHwCizmbI+zfLG1nnVa24rCBr1tnQYdmDx0JryuEOvSPYOkDshN/osEh6B1hvuGKTZeMAcmro
S3/uODLGS50VRtPqefwKpF6RklWR/5XO+mzrksSXD1Gi66oiTR3al9B/f1DAIZfVy76s9BZEgoSk
2fAA3pzFU3C57svLF31rd/HOnvUsYa1TffoURwAtKOLCnQ7HOs8/LiST2LahPCohOfF1PAU2pM1E
ZsIzfWTjia9S4OipR+TxYsko2zV+L4w9/OTCapYanDgQM0JIcpupChh3+S9k+Csob4lFG4a7tGpJ
whGN6N1TdyzQ3g0/YMRO5QDYkcvShvbAyLGABRtv/HOzbdxC1wme1mp6UMofrMeQirV5Lt4So0Oe
GcJixQFmU/k3Fl3QNxlHeQt+zIkju96NdOUgDf+MX/61wMrX7nszXeiA7Yz6fesuNyhqWwfUxRbL
btIMAsSW39oGw9jpYSJUH3EN3q3RxgWRdgGBw+iN/NtkHKW4nEnHTf1MVWKMDYvep83682StVrsC
RPWt2HAUIFAI0Q5fky5K/1tmdXSxvG4zX6RIVoejYblYib1jWMYMvnz2pPKt9hFK9YMsW8c6KxN0
OeDHTOZbqoHpOkKpT3GMwy2HZ0JWSmWanjO5eFEfSZk22XmwURXHngUgrx8kDsbMIx2CCOAArpCk
h1AJqlZ2tBdWxYy+LMWp5VT0CaNj/hhWl8RRqCa4RyeBIzbzxkuDefdKlZm0XiPCOSfldRqiKkS3
YUV/3+29czTTd4VphdZ5qHdSvQpB3IQj2ok86PlpwkUFvT1GeZA4tuV1U0yiYeIwa2jcuWjGnvm+
jLxEs4WbvXtC4VposBQmpuknZH6tuNg+cUW1JVRnWCldSrv2zBpZpcYVt1B3yuvsxGzo45Q5Pgop
xrfFKNPJSWyxYBN1KqosgloKKIitat8E0jwv1dkpPGpihKhgvkkZg/os+9+S8PMdOTwGDT9A2zuC
dwuBhXKbpibdOJmy9ATf4HhGGoSv6/0TKQMgxVtXzkYtK/2aNklX/AzV8nXrTjCU9A5tNZ8YkBwI
QBvm8RejyS13zXnf6M71xUQ926Ey0TzczQX2i/zzl4/qfKh4MTRXA68FhljnvN+bnKWVtPrLfshb
S5LMAxAi2Rbtpe503NxUJUrzQDF1jS5E1KMMxcTXvdTgC5s8hTxx2kLJ3XEjk+AysUJQIWGXWTo6
UGoZcqpLzTPpAsP5kft/BzOmO8m/yWqwavF4Gf8W5Ss+tmg0LvCdK8/YflFFLXFKj9p0yESNyZRb
NqAWoiRDNMmJTxuIyTb0yLFclnx/w/yXFzKJiky/njD40Bx463YoJZ5d/U9g04MbERm0EqFGSwYX
mNBxeTrqaqZIJSR5vFhArn/Ygt+yuiFmMBLbDIPPk+EUEEBmag1hK/Pnb5rCoQgUbIbwRbt8Dsja
WY/UXBK1TJqoWer+vqkqnRNUU4RXJVNZfslN8hCfHkd2NOpN6Iw3/UnpAQqQBBcypzn4UHLxU/t1
A+xhDcVcAi5RzpSE4ZlUaLkevMmOusbDqkRPKKqN3oWFrFnxO+xy2126jBJt1Es9tq3/as0ZrA3G
lBzoYsCVVI0b1AdAvrM3xQEo7vcDOZsZzTcOpyKDUi9e+1RPjLovpJo1YY66ihGqf7mrHT5tJnhf
JzWS404cSNq/7ja0aJHljrN244ZfsUQrsN8QfRxnYHXtc6PtYPnBCph32WiSQxo+/uOFsdqNQaK8
wQElBMz9ya/V5XTlU3lAb0d9l0Cno4lxwIXaqDVQWUa7Y5Urcd4ATnvigTEY4cp2jiZlWQag06uA
FfV/6wmDH93aqp+cTcYY51mzIHtB4dPHsXYtKG3wlbs6aiPtU5pUEwJL5c7sOw7DJEjjaEeftzbd
fFTTAmAxNWPYZoBsm1UhCs9Jxt9DtELDBPkjsoGzHRuRQEflqGWLlxECptOX7/ZGYcZu+2J9LC5j
wZJ6MsbFzNr/KDHrHabApz3meo/ejzTc5FY1Z4dDR88LMqz+agLwra7s4PBfGx3f1bMdkMt6Jagy
A09IKmRlZ/FakLGOIFU+sbWxg7VwJZM/L68ibqKw5MmjbrIW7uAyWO/8lv8/px4uromwcWz4XeIn
2KP1VjuT4HJa4idtEeS8lBm6zxwahidptBfOWr0uMbxQkkJ7CB5rqeluunh0tFoOWFiDT+Gy0qNh
TYRKjwxW5G1AaVV+Z6zSc5/xqCupRJ7q1U8cGD9IB+lfpfqxFjO/VgdYR9Z4b6wJKwYbpMI9SOFo
NqsaOys/j8a7mi13BZ0bMCYJBwsZUt6wRcI5B/LkKAudRWUtYkGIseRZ7YWNF/JvjCwVNMXEBi6z
aV/BOC/ZIzCIR366SobRxtIYGyHWvx1vCj1FjCkxzxZgoR40Bn5tCuxaEr2q1jiKbvyn4DlrI82M
p+K8d3K5BUt9MnATwuj9BQ97EM20pJhP4YsP829ISmYSTnMp8k6llSq2WIH7wpJdk/MxmXea1RC5
5ny7AU9dw0pJS7lr5ewRjpcvXZ2qmhzjwBUNKgRYKP5U0I/FqsG8vA23StZbFIHl7zKE8oanbdh0
fKoXO/yydQMfSyul0bzUDf2vrC3JQPO31WR80p8/DoRs3C413wBglhb9wptp/FClmceSXMgFmzx8
vb2S0SKpQTZXkbHh1tU2mZGqij+UOadlwM/0Dov6Ou30AIycc4EDHN8gVRVG7Z2I6gVgDKRbVrzA
dKXX04cJzzzb0gy6IPzfIQYORMAkq6Y5kGFLGfeWnmUTCYAqgRCh3NGnPCOwxSUIh0JD/4d5aTUM
niBC4fZjbNI+ciTpsha3FaUkD1JyMKk9KceCRWYwJz/PR3HdUTafUD9r18o6Yjnn9qnV6b9hZFaK
Pc014Hbn3DvX7BuFSiL8ObwM1mhicTb0YgT0Z88smyd3RSRF7mY3lt6XifjH7RrKfilwnf0mQmfQ
NovZ67lRk4YhFu7pZ4zPr6Uk0OmylC3zI9ar0I2k5IMMk/UP6wFhAfUgc09oedlrmUm+xdnvk8bY
fS5ACk55fcoWrNlgjHdtUpGuNwPC+EQ2n8GT3bCiIGqsAUvjv7HM6TrYHDnt2RfvL0my28BLJDXB
y4qXsKZnxrYLS9GBjw2/6IdoBdBoNUweFr8sHQGH/7/1WFcVTYKSMvO5yL5553HmpvM/fzhwvLu3
ocfIc4yZD6Zw9gxh8Pvqjuyqua1o9G1OqePR9XN/a37g8z5gZKOy15uh9hUL9b3ujGsn9uw0gC1u
DprDYTDrpJu6tqnfNC7gCWenxwgpiAksHdozxb1UnRop+fEZz4RxZiX6GXWRxv4I3oK7n1gTmFLt
LZ4YSKPPMiJwXGaNw6lt8Jns3VVeTmueRFZQwwIFfXHcmMVIv/8m8Zwj7GpRtdQYGAGrMMeseXej
rWTwLRVxTMLAp4e0cOt5flOzM7lkPjlMOCkiZi9HjLSuF6AeUVMKe6y4vsMM5tJ86opYKNjTsZQW
xDyJ62KGZ6QofHqGrlF2eKV1osEADI4WVBwQjRKdn8VgJ1brQOxcAt2G+WG2bqaZbmFzFZ6hMZaO
tfaxtoZ4d9UiWkigXOHGAUTmg9kIy3dRza9kQEHn7hBeOal43RL+BBRANukKBT9G9xlbTZp5Gn/d
rmqOhNFZIUfwxW7PAAHS5UGvshQosi4wQVHpeumbFiiw4/jL5jL5YiiLYmB9uxxTWmLTRkDVrJAP
yJr6HRr67UJEXQIz/g5/wZwbBHbSqbstp+mScHjod3rBZGApX6nQ+qFMYa9M3juR+RqcAjPLz9u2
qeE1zefsUSHlZYclqD0jmTzcgyfzijTSPNZ7jvknjWQRynnJLzTSlYK+A/JNxtO9wbeu7WWYWCzp
o4aUS8LvdcgWNYFSrjrPUgz9sO3FHJ2CRUohkH/O2vNdYxYvz517O1Gc+mIhcuQvZY6gUZERri0I
2KMkvuGnB9DwlUByyzqnDMCLBe6fFc7VG1jnncupGxIqncX8io2qJY+qrzB6sSkYkWqQjw7NpPjo
dqkDdpqltI+PnrysaLIM4QdnnwzArU8u7AXHYH68ldNCbE9DLNuI1jKOgloqQ5gpi/ZWxH9iE20E
N+VaIH0JElc0K6H7T+loliJrrxlaxXy5upLTqrRskGI7sez8rSda9ZAXqcdJhdQ0G+LIMgoGlB7F
efs4QN05M9mR32SKZUukhDJiFBfF0StKKi43lgYqxQRqkdVz2XukJzkN99iLTZe8/bdPz7JIJkre
M1W8oLhh+p5wNYxZjT22IDGHbvmQgZnqFo5YbvXttMf2UR3Gbt0srKnSdhcyqm16sveh/1cVh7fo
xt9LIXnyPlHzSXWli3b6pkgQET4PFHsdy3vvn2He2s9ilAWoBcSxRohvHNSc0Qe5d2muU/XapvxU
XcQpAe6OQUyb+lN/WecHdSjQgI5UQxKVNFjXvlD6khMdgUKcpjtWZpfFeKUT0UfT5E+y6qPSv/mw
gz8zn4bcoZ0TUiZZDbo4Sd9tibkNkbLpAWv1ca6RYKVHePHa9TyCMK6rLuhl5ALHbdqXEC1HrnOP
CiaWmN6Jtce317wYkFyViO7qghPGtujbaWDcUCs0+cn4l8VZas5LE4v+UX8QBpT29HYOr8ab9aKL
HvBOQ3WmamkKLH7Gj+NGpVWXqJxjvTXxK2pmcIaLGgurVeJs/7VQ4+S9RYEOYQVTCdFusuh6xgn/
p2VR6PSuI+7ixMdQ17+nDwUOadQAMAG6mxq5SXQNGSE30dVRgJzLMVmlIH79atzaMruS+UFgme+S
IHU2C7cHoFhNavN8VkkHVVTwbGSor+W3e7S/EWJyOskQwUrOLCXfrA9bbUZktykbFWZeMg622v+i
IPtlMvREPE5Zmy1JbfGvr//2cdGSRiOzh/w7jFs+mXo3uV17Gk/jiOYAmx+/1VcYr2SIEbbcxASV
otkNPpb0X198T7pgTYgrQO5ZVOGGTyipC8Ip1OB6DZ5Y1yTAbaaHXrotV9FjrUMEQTLe2tUPjeg0
tS4xTUPCOVHlW+BDZcN5I8hjWH1C2yUaCvj/aVhIK5s8k4DUth/v/JVKkvPQPWgzmM8lNeScWwMs
XUg1ZpYriTFm6e2yTiyXHbO+Rh1z0nMkDS7/0v1XFUZY2HRoqqRKI09VfUEXoPxRZPd3kcYEYgx0
7pi2YCNmuEX3wvBsRhfn3qcksYnwRUt6DlOzR+oCD/34W/fDzO1aPC5DdoEwm6i/xnWnaeHsP3L3
G0h+OF+0kFW8XZqyXHJrUzdPNXqb0yxoia4B82NHUh7LaGcqvxTesz70qjOcw50b8Fyvc+bfs82d
pH5qVnQcwt/UFqAqf6Y6s+LZu66x9pkCX82tMIYevkDHGEFQtxSnZ0QrJNlCogwNldmx3VUERyDs
kXisxbO/E8r4pWX+E8kvAhjodXxlJb8JFIJlwpmEjAttQw+VmPMXywSPApwNmOtralL5Ryp6SXsQ
nfJxUU52URrqt9tcFh8xvZ2hXcqc8zMExAOUEUG1uEepcmuFsRRx07b3Gcex8kh6qwzeEv7Oi/rv
JVV4NAFxichXqrsVHAATumRKLEhgKqypgSW9UxHUTEa6eYWdNAsJFrZZklFHYt/rndmTwbQQB/Lq
FxVhOElWU3Oh3qEOo+ZXRbPKa2BIsVcVOq3amzK7LPgV1ex7evkOdDFwWz7j5/0AXPnygKbMDwGE
pzbsjt49Z5OX+iZDOldidSeFHkAi6yFAHIwGJmiYNRfPr63yCXzBImJM6mWOPtKdrxNtI0QhtIRZ
TeBuKdmZC91BTlUppSgVaSr5CR/Hmm+iifuPMyZmDsVg1HG+J0/p06SWMpxBd03t/yvNfdUnf8KW
TUgaiMv/7MW8PQpG/GJ0mbLjoIrGdYbLiCG542FryB5tn1FY1gWp9ajkBj5CGho4ueZ8tA6pNRmv
Uo2z9wNF7gEViQ3DxOmj7QhXMHvU4ZoHTa0SUndNKTogBnHX0cPthuXtBiqrkm5/jbRFjZ9NnOwy
rKxUD2Ph7THhEs6iY6iDMq/EQNLjDqdR2se3f2pqab3cIoQbRpBYrl/0xskCQZJh4TZqhQi94zIQ
ysIwCpquhnfdeepZzKxvhFevLI3WRXTQIgZqxmSZVsRITyj3nYID0Npc3HhwAN2GZl7jYHp9mUap
RmYiXROJyE+RWs4W9EegRyFDUs68GEYBSZxmeiUFW3Z5eLAraYGekThIiEfm0tLn1CYVQq00vrIz
7CuShN4txIQ2Z7z7FbgtY/UM7UIOSZs0chpS2D/l7zSISEvKMY9UcDsHEioySZoIwe8KfYToDADT
Wem5WuXi4Ls6jsnYquCyCJveBPXLRjJ7UO4s8TD4112VylF+tYcH6RWuxN6gfJUT3JTcSfSqepU/
kau1rK09w/vK93OQ6u57mFvKTp7xOrTogW6VH9/TGZKeLDd3GfuYG96Kkw6oTFdkYLSwrbjVYeuR
zK8bAoyt6XsPruVMCOWyWXxkY8DkyB7bKqovADL4QZXLg3Yo3A6sWxbpKlMHMQAi84uOfnsRPS11
ECgLsz0RZBVw+bJ2Ct+RtyYQA+G34S7yjGHAt7XMDwehTW00xDOUvxLXUe0A7sTW1l2hZvGC1gLW
kmIwXU3vWT9ytoqggXLSMppzXWjNcFXFgQkisbOUgEj1jIN9W0AjWp0npQQMKYzgtrlZt0Y4BJu2
NJj18Wb6Jha2MHtlMeS+OyHLYns9Kq2ZzU+45TJ8XKMazgIbAKOr4R8gwV1P3lnl+yvdEn6SjHgC
SQawZoUwEdFXgfiV13u4Qj0e3GjOHCZSrTcCvHHvFcZHhUXEEVC9ZPU66kjXyNc+qGCTy0o+LG9O
XEnjLqNGuFygdhAiCeu5S9m8FrLlJrVbZdqeOu3OHLQIN+mdbwp9+XlTmK66Y6CKdB7ZMWztW4sl
NvM8cnfiCGLS/3Dlenxp96GxqIeSye4UypvuubNx02ADhTxyUgOWncD1u3k+jM19pdUKqKMog3FH
vN3SOQA+kzfaKWbVueAAuJi3G6edwIdX52x7vTQN4umwpLu1XyPN58ISPk5kjKf6wLlEMrJnO3MY
mqs8WyArmhAt1H/T79wCMel2jl7ulkrBjyMOwrDbaBZNsfDDe2wNaVJtH6M6QP/QBeBEXlAJmsoX
7y3PrwfV/v7VRRgQEB/9sQSOxTeKfQZZheJXzJiHjaA/u7IfuSMvjg/LA1nY2kLse9eJyjbMMRh6
C8glF+ajOgdvsTzpwvEPjUBuLFgfHDKfr7fdAqWob4BQ95RKi64AXfhvVKlBHEkz5JMuscX6FPGE
vCdKxuRK+5dG2rGW9uhrlDjlcscdP+oh7r4bxp32v5AQ2jkfTYYxfGBrgvbUFwvYf46H+Gbf6Q0G
tQNfjmXpAGCQ0XxvCr9ySHs2Zhtz5fiYR+NuO798D2GfasqDBA0l/2JbvY/taL2irM/kdGEpDf5E
WaIl0ba/iewfWi80LbbvRDhjxe0wAccoHssHJ86MUts3aeF7OFy0vhWP72RGik7hrZRMtKrDjjzf
wTbVp2oVJvPrZhunzc/gsH01WXcaZxHiZTReEqWy6z8sCUSHAo3UTemsYvz90KfNtcAwbpY/w+B4
3+FI8Jg7OruuWwmtcdFTQalNqpD6+tHlgrDCKHa8TnHoqVQ1pmcJ79MNBMYlCSG14MEqQzK4p8qz
Du9apK5g3sPOAUFec6I4qoZ+Pg8W1se5KTnKWT1vawwvLMpxmMwLwQJjO6J8qlxSCsS6qfJpjUCz
lczFieJDTQGQ7QcyJSiY+D2OBuq0FOZh7NLfzTCHGwyYDeNFFE8/KdRxLvo65RPfO9chIho/4SSN
I37RIipts89G25meNO22+wiLW2e58mLqoTNcF3Kx8MkhMZGyYXJszAnbsUex8jQkn/oGs2OugmiV
pZXvI7TG2nLQJD57YYftxsjVaKW2Q5VMRSTxehbpofFkU1xLB/d7Ewk+Iums14j+VG1Go9WBHBGm
HXSpKMz/F1lPc/6MJVQRMlkdEuR7SKb7hq4J+hJdCYpJVSh2lJ2gRvmYzPpIJ7e4gXdrm9GyQQgw
vK9U/vqu79E+vjDM5YPyA+SIvki0cWyUVrH4fEehpum+dEFZ27cZ4pkm1eyteRbxOTIvUEtlcd+x
BzrVTN7iYbgSPc+FKTWSR8OC54/W4RmPT1vAJosj5mLQ5jLxMKuIa1xQV9CVOZ+u0Fyq9c0CDJes
dLhiRvOnrzY5jpZunV07l5NDtPcc3mpOffOa7lQZcm95uujWuriJBrfDi5rt0ZZWWhIZnsQuG9yh
rAudXtRDH/9HVvRzykYAwAOiszbdhJvYontI9QW+9R1WoL1UA4jluScrTESLngZSMpfir+OKGoA8
4+kWjcC1ijw7fnvpQmpAy5GXsoSzv5lZ3YhL33rTYPQXZjfCbW2dMb03VaqslfXc8OHF3n9EQpZC
RvITOc+v4mBKPJbzkp7kFYXxWvFe6KeJWc1WMPdVb6nbiWEap7c8f+h/kaMTl6MmdEv3C3l5nQq1
z2Vi9hQos6TSXo1Qt4QxhCBX9lX1TOVuLiCUhnlaxYjtiH5ghwi1gl5qm+Ltl+Uj/3Ql4hLCBNzF
VOkxTrN3g+JUDAauXFY09e2V5OZotR0gJjf8BQQrpao8KdeND6Teoeyhf+1AjoVViMhcejo6OwdI
wcoOjIVYLbqeIdF8gjp0UQ3/UlZfZYI68PjKOPu2tPfkmacUENolE2KRXExXlFZG/+AdRPZOFmxj
nPDhdDff5gjNQDbo3KOxeK3fvt+g47yvDyIuKalUsE+pZBotkfmBRn5MVEZrNUeVMQsKY1BgZiyz
QiTx+mGqFA/T4a9P9Nukf6PPrdsorVImlB6BCtaKOmkfgDIxAN9oSDrSDhmEDUHXoiz6SUZ/sUCU
jn27pJZdhzJtGS0mcQxYS70PyJwyL1xgXDZR/1tNvLNnnNmUYI4znoBcLzZ0PP7kmEqcfV8K6Qug
m4/IT9L1gHrLYd8olhIsvThYCQYdSDbRfc5tZvQl8jDc/B/7/C4EiUeb+z7/+hLZhK/SkOPhY/g8
V1Rz2hZhjCRQGPL8x3EQk1mCC4fZPidJgEEgwEs9QYX2e3J7NUnbo55p48fQ9m1ugQd76/Ih/Oe0
7mAr0PpDzgH5bnvVr+8yaTS2TRnCji/14bNdCWv+TOV63DXubUokhVfegMoaEJF5KyOkAdOo3meS
TMwSxWREucERmXpE6qYCcc5mYA+Fvw/JegEzUwz7oSFg+DW9NOYCJY+iZ3Xsnt3P5N44W42ZOKZN
r5F4moNO8RxR/ZDBkeArDYBCygiudYeTYQv2+WlMbt5HeGoJhG8Mxn7Nh3udEBALFVmX8KfO9HG+
Ap5LPuaZYUZsvqA/w7cBDjTHZvDJNbsjuGotwc/sGxem9eOY0j/8mEALSCYkuxkFxcT1millMfIu
gNp6c3pYATgN/Ok54tbzkayoOUJFrfOV97nvulfqQtLunjolI59TnBjk88DljyX7fVw+sXRBw7Kd
D48FV7CsR6vROPJgws9LE4tgw0agg6Bbp7nHvzBceG6zsnetxbnM9wpfWVfzDZ6Noh4d+AcBpsKL
+m86sT1RIuFZqVygRaerKcemoXrHYPwfKgkXs5mAJx2+vXAtgaGacyJgoaEYudshI5qo1hQ2i4Sk
NYpn8o4wi1wN/GYOfD1EpaAjjwFpiQcP1J8RMVD+u8x/JC0GiQ+ooJcl+fYUdl+zp8UZwygdrrhr
RA1ii1uVaOAlvPDx6Dcwi8O4Zg/psodjOoPwz4shVXJgs/4EhwySqQDknR43La7LNhEYEu/v1dJO
+oSiH/76S6vJifG3iX/BHj6Nu5Jz0syH65XSTPCzReTiv6ko1yqonC3gmNGs8t4QDSC+EI5kb6KT
gZ8SVsNajytHeL9dpo0ek2lMyJ75xOuni8qH+FdbrO1WQ4N9S0hayugslV+ihoZHic9Angv8CqR8
Jbu54d8Zm2xvTUlgvL/yOLf/dhj/8+zFcepm0b+snKU82vuDi7F1YvRAmbe0bqyNXI9821ZvrPa5
mjWzL5v+tUTljkg1Q4aJ8Qvh1CvCRhN1SzXgf/OW+v0s4NfZYlcLRpFJU9z0UTX8NZY5kNQATt1j
UdEJgcKZMkJsVVWQmC8rh+2tCGPCTPDCw+S+7gShac+VFEvTFn7whnPIv7e0qAC93ARQn7iQ3xz7
TZKCWRgYWyrZZCkb2b2NKGQZjtAASfxJoA7LZvyvFNhgH9I/GBbMYKP4xRbB7qD5vFJxl3Jl1qtN
eltuBhbyhKvzZHbFpD7VKr3yygV6U3pZmup4L2nAfDsLQLv61mveZapEVzh7yS8e5ss2XFF5hQgn
qWNpNBRMK+YENLm1R61WZbJScxHe5xFcbiU2Ruyb8nGlLaFAfIa72Ft5iWjX65oesYjHtrcBqWc3
Uu8EgaA2vrBX4OwQOKKD15Bz4RFLRB5A8craToRKW/aCMsfkOuAh6c0URKrPSPn1WdearfRIzsLY
87Pn5vVIuIuBQ767hftH1G3tTILgUOWru0UIduCXZa3dI4YnMrhg+D6dZULE4LD3ESy0zA6eVVWw
0B9/ZRFOHjKxfGDZIK9YonOZBtynuXLx320miVc03MnPnvfhiHKeUsF4SY6U4jRG+Mzz5zR7jmbd
GpdQ0zMbCMUimXs/xa93miYAjlNij0dmfv1PmKfQivBMHZw0VoaJzLYSTDug1WhHIYjUMRtpFSNU
DbAECJnKccnHVhuuwDU3vNk6CA9SkKlrUKhqpb0XTUlKv5ztZnEhENvw3sHEroFjKDlr59664CLY
bTrcYu1M1BZjHjhFCMqJVdyfdFHlJqBFJvdedufppyT4K5G1sqZgHk0ikps0yzUeR6yTaY4KnWZF
XxRoixWCHAyZB0AsDMWAlRGaT7Ek22/sjosyb7kX3se5QtXlBT6FyMZinku9aks8881a19HWDFlD
VGLP7YQoKI3y50Eho51W1ucW5d7DuO6erMWG72CFMIC2MmRyZ203MOzdqTezcwhTUsR3Y1vSKI5y
vB22O/2VJQwe2gXCGBe9tGQ0vcb5wT5mvC/Yit1b/Qgxk2bxG9uoMVK/17TvpZdkzGYf79DH80fA
v7VlFoiwB2w+dNXeadtVh73214kEbvoLgL5RMi1cd9Vie5YArtmwhQ8HofQnoI+L1aDqv45x0lUr
+LHHJn9TUOSaOWNaSxX18eSQ/foZb9KZrfcGcLEDPUZ93G1kFiytTOiFW2d/7PRoDgYbVOXQog5k
okR+JgUrRMEPZsuUmjX2CiO9SDsUKt6xCdkAciyR6A/5ShHivrlegFeP4RGHNv+o5nUYWJ3gtw1T
qa9fqCk00APAcRDmPY17F6UwhoxlbydJ9AOL3I7cfGx+mR6G7c0nuwMBO8OZnDeE7vIAfzAgXe7R
7tNX+CvJ+MRD7tGdixW65/y9dv7ZrJoyI9ZyeVaVM1nJ1VvGUUrEDWSqWhRMwxVyNzWXD9srVgSz
cTkFLuxNqzhe4r9Puig39oybN5/ncwyAB5qMNNK+RsAf/zhOfwd+HNYnkE8j5TaWtd/CFkz8ZG8G
TOrEFy1a9ndnBYDbOp9nGcaSkz/AQef6BORoYKHb8o0ZqlK9JwN3ACtAUCSlNpG7VgeyQQU2EsxR
X+UPLvKBntyCGiHr9ziJkmjLotbuQxDV4lA5mz6fhef8FRBxtgaGnRIKzPzR9Ph7Hf7GgepWdddf
ybOlcpZzUSXEJ908DSxyPTExj6+6nO3wR7f+IeqQ+5+BVCFLP0k2K3ZDAfwKiE7o4lo5qr2ZYEVy
nKeG40xDQzcBEhxLJGl/94J0Lo4AOI2bBEZDSIo3bc2kD55atD0dGcPcAfDdXp+4OjWzfP7is6l9
kVCxheqs/lfYUZwn0zwciUK1PiJyVyuE1BRCkuM234vgIEPncJU4K1Ha8d7AsBcM+79+z8LViqQm
2Uf+DZbwiERCmQW75oZ0CJGsKpwJKibQEzsPmhFyFgWsQArugmxEfcBjjzxQhVg/YVcQfkVP6zV1
XM4uIsyAiVYz75siQPDB19jZk/jC9vlDvpF+OpAvmmvipwzhvQHaNzkmIutnozT944ez/XTJ9k4o
rBj6BtWSq1eI4H9vXMdqmtqLeVPR2a55B58ctELB6kPqZX2PVbjab+fMj/oaDGCOVI5XytWcWZ3j
dskEkuGty5+r2w0ODH6lnbclueB0utrVn4ocf+G1HietSKZcpDn1MCkOVhestC8kTtZwyw0lOpT9
KdPqTiu73Ir2c4iHppAfiWIaflm+LzBlUjE8BM7lIl1l49O/kPaeBPGgf83kSoEZB8qjEPwNQ+R8
Wl4ZXMHqXDMVa7gzM9VWdzpQVYz7Le8sutphJcIwdmc0/SC6L+UQFZBWHUGS7OlqtByPnQQUD0jb
S9k1RJ67noXgY9cGXf6NEY374eFGtM5DX08PSslCnZ90w+q3CSZNFcfJ9CEwNuovvOWJ5rCzWXQM
0xXN/mwNaEXNa8rY74v1NR6gaP027WFjRg6t3JdYRhpJ7S4BTQkCcEGzuvYOUyQ6fl36VOP64tsf
LKfsH5wiks2v2DgjMuM5SrtWtqSkzSi1K4YTmtKy3im7U/7z3UgRaeuwHzWOldKNkVvVDyPKNeyw
dy7w0majC5ofcAuCth7K6Dd33jRGZRBqQ2CC0N0TUp69U2GCfPMGTswBzd+Y6qCgL/yiAeqsoZGZ
xRsaTJlf2D6hfTMUT3b4JRQhtZExGZkDCHSGudsrezif7amHrHo0ALSPAMC+PshKMJd0RJKy8yPt
LQznKUc56qJ674b6LCD6M+TKRHb98jC3t0yMyziuvqeGYIAzjSilvDtyHd7IRCfkVQaBVBoR6Lnn
1HAPWV3nhS9CTAT+Zx6fhGXffbA24r1vMnf3cyDVHn7vfSfmfVfVB9ZhlyFmbuZShtEXEoOKYysp
2PYQ4ICiYOZukWjoY2YpI8bYAdZ1B0JFjrBOzsb4RGwBfY/tuX5LGzulOTiguee9WYzkG7q8XIr5
aNKzg97HEPilKFoQ87d0bhP1WLwiaYZVEG5gLSs88swyh//cjIwqtyX4A+rIdiIG5K8wbAKc6x/m
6mqdV+F9LkhzSxUKPp/LHPPdVulFCn97H7BKS8ehuiKn7r+YzApBuODVqch6vVM+prwl1tK0HF77
pL51Wbl7EhtNCF8i2bxQuFJfVe/JrrCE0ryKEK90Nf8YMh91+wcTcE87aTwCRBKL0MP8Vb4WVMwr
6aUIcdv9woATrwHeD+UTZphFg/Td8xwscTVnjlYIjsGKyfAolhG2FHlB4jAYyypV1fFRcvUCtBit
XnpvYuHUCWEjG4X9pqjma3dkLjIr2B7lN4jIyW1LqMuemFyr3+qdFD4EuuRH0x9ys0DUXusC6fTg
JKGfEYWGFLq8Qg6JyoZmcFxHlkMqf+2v7uc/lVl8phYcGfMt7rj1gixWruGPAcD7XVOEAKrx2Hrg
2P7KssbzqbOBHq1Z6S7c3m+5XFlMKxM38PIlZ5CcpEgA9MKoI7NuJH6BhSIJmMa1/pgQwOMtpHpu
RHEmFjmal45aZbIRwizqIHeK0DYblR3nL+PHWkcENHKPVCqGzU4lFiANUGFhWuVbkj2kLF4QU8aq
CdORrP63SN502gzcfm4InZrfxZ4n3kRBpdZhqUGSCe6WypZ0q7JuMDobDSSf6gVDck7o7bzriMEz
+ujCgq7fcY1qw0zwpbRGeagV549rkYPocuMjyeT68zeK3FMD/Rpe57sbHoKrTG8OfPv5Y7YPm0Pg
a5wERj4hpJ8sdd7KUFMWpC05gC8qxW3VmuJHKkFw9B1X6nYCSL2E/eQ9W89S5DjrIKy4aRmrh9PA
ukX4NUpd5Rj3ToZNOocPZ7H0AJwIP7n4V82ujxDyhtyBWqdSuCMu3ae/qU82AKeIvlwf8S7dVG+5
GH6pkxmzj/VPbwCwBKdl6uQqrxKxywFCc32BzQgrWCRazN+1j8pOJEwtutiybg/UNUmVzs5KTu8v
11zcmY95GSzFb/TsxjQnPy9AXTUXHa2DEdi7ulAC3qm6LYqp7gfwl0jwrsJD7Nc2tOXswMJHR8ie
f3wd2nGGd38m9f/KX/gklG5wX052Fh//C+7CLMTggFm6XUn2E8M2/GoHCru4A6L4y5u2U22aYxJ7
o4/InDnKEytSjPCfp0t3u5qmWgbSqyVxgDhbmza6X5sUdVFtK2lwpwvlvaWdBuWiFVQFYjXn87u5
/AMR0zDRvsbBDopggDsOBZcZbVLL8atP6ghL/lWEVqmfF+u69z9pjKQ3hs7K9cwx97d8OSEHiX/K
0KGS8hlC8p3dy5IRrP6qQiwb4Uj5LIA2KH5tU3Zypr0UFwEwc3fbSnsIrQV/6VuemjpuEGEYRZrC
jTKgdPsOx9GP32YYi0WTmDwnFhn5gHXnuJorESJzUJZQ3Q8w0Suz0vMtyLZIO3rY3Jj7YJa1Imj9
Sm4Y2lWVhobrAzHyE3kQixTjNhbdrCW/J2pAo/vHWLJGRPw6OS+Wqi7xzPVp9qYEZQM3Q7mbwRUt
JEa9TObMGmMhVhj2AVEN2s91DracfXW7nIlvJ0p48FlMmoGZnsDiXpfLyKDf3S0aTfP44YtpKBKO
dCLfrnLmjh+bX2TGdcTedEd3OkvdoNUmgp0/pL5gJtOjCs5JB6jvnot0csN8RkpEnZqrY/dcrfnc
xzM7f5SIfJFTlBj3js8yNoIqvNZPEI51caS8cBnFG77VYCWCDaijaeiVm7qVBE9CL979hGvrG1kZ
SwrBJiDasdvzEX7nyL2ZXXGYQCyvC2sxmZmQxNdA7Y/h6VU0XvvWYOzS8VIum+1Qm72220U9uxLe
x72SzymsRg85oqMXwB+riDUYHBk1vYPGCshEtGUPkqFHwr1nYAg9LCRlNIzLxXhlR74iBt3Kdvly
9TAomDBJdsY2ea2RgGLEOg3lMwROeQZnPVKjZ1uAkzHhFCOWjW+UC2RULYC6voTxdh9kXAzF5mNP
qK76QelofCn00QOIkRbmW3RMjj0R+GiV9HU9gnQ4RKVydmkT8cL7TTwmXrQ8b8eFvnEt175LVzVL
c8OUibBiHxmniUpmq24+d8Bs1TtfdTeJ3oiEik0efYNSDhR1diNbPSJo31BY/lVr21Vm79FcDyW2
whp99tsqMm/QlvJsmgF3UNsBR8SXBL7RY6pDglAWHEo5yIgITkoZl0Gzh/XMMUBGOxzny9VJ1btV
bpxDv/Np8YVeZg1XwLmd9iUdwZ/O7hVykZDYxj8DSz8JuGi/Pie1hDT7ONJIzg23Aw7LuAC2Mdjy
zCf4wmS99PlJv/zm5Rye/iZixh0SlaEutgNjIfjBvUmKgLUtb29DG0zdJcpVx/gNWOeXMuGGHWTV
GA4Bm84GnC1QS0MGWA3uBAmqQgPs5tSH283epkY4g+JJkrxERnnpkhMZBid5WE3NGS6koIB+aZy9
PmrL00V42Ov3ZDYvM1Q4moyAwlGicprBOmQMQ2mUnc1a7+bO7JRRMSbEGF483wbGLdm8UeRNZYri
8XQ2ZI8sBnPh0tVPZVKincULTJIHP2JyBslNs6mj3RbdBlvrhCaiz+WuLo9QNGjyKQilO6yYn9xf
abJNcuCISD+NboKDCzP4qj8MFb6QVrM4lgdYOILuisGJnHm7TR//IzdVSb+8KsASreBBJh0exO/n
hdIUQtT/TZIhXOKbMeqHs9McK3UpNqppVaPHN/4vgOtNfcy5ED4iQk0UaxbZYXwAritOmTYKt61G
TPgkjzlQqeFO61tLQsqg4LiXQdeIb9E/Ed9MQmtkFOdsHzwFxjXV2LXQmdr8cn6+Q45IEyh3rTmG
OXKiqJvxXwGWnwvusmL0TLLS5JUWQY6Pz5BUKRyYvB6khQCkQb0ji2+DAZ88NDgfZqFqMH2X2D7U
qwSK5PT8YyT/OX6WQCzsztmaFAE4ngvacuur1JqbSu+iQ8QZY7bx2FOTiDsaU9Fv3eZoMRdZ25PE
6QhziuypvK1xkkPppPmFVmHsnMnWbSUss0ENZ1OqQiJT3e4BbEv5s8gBk3+sKi682gxcnMgWYjdW
x4gVd3PmS5nvuzwtKGB5aVMrDYkTs0/REqHCU3YUTCqv8WVNW6dzatuErYtHoFUHLf+8rPDlWVvM
e+vSN9+aNgIGvCCMTwYLe+ciGAOe0Vzuuqe308oAGDXpuJnESKs1mfArPAD2hFSHLO00a+OSpd+/
tVSjfPGmh7X3mf8rhA3bbo1YlBu60P+BCsmb8fMlgI+7euEGWhUGJ3jJq8HPplxMrIdXTttbaMNw
2qPbiIoGGo3QtBbk48hewcSny+iisU/jH8LnwT2upzRVzAcCwvBnF3DX0W4L1ESYFQxZSMZEspF/
veO3fb0fu9b3D0SZ2cRnTLoNY5z6D89kOqkK41QAJENX5JrlbNFTgSTdnQ/jyxsfJmEVmuETwExW
ZUUs/bwhRsVuyZosAA4LpkeSUNmo1I/IW4iWLcdyp5aEIwZ5y42QrX7i1y+BTiIR/lTzUm1G6fPi
YNLcrGfK+HAR4uql4xSDmuU5C1EdPptTIglRNHMPriCuucx7Sr0ykSfdtUMUmG0+Baz5u34codJp
sdVeU2xdOLT8GKMDPUERv7ELVXnbxbBp4hYLFB/ideTNO4CszQJzZjm+lrxZJRXjRBygrBhN2SWp
nt3QMeXGsueQojz290RI2jN0NOBB7c6QLhieXtiQSOX5wxmRjPYGZMIFRJf7Q/wR3WvI+YKpD3bk
Iy3m8F0nWCnGwEbnxUmBD7hESNmwl9nUlJLqjqp+5HUIDYTmD63517QqZ4mOO/bWCjOl9pD+5IXe
b1HZjZglDjPTo7geLBy9GbCLI4oEfQIoIFsvsidBNDV13iG4QojXiPzFEr2qKQvH9yvLYODwTylD
gTQHQD9/rBUFXtsz6/Uq40cpcQ2EnhukkuwsZCm/mg1zYJns7ClxJ1IwNGdXPZlxdbFZzyN2ui5D
srboJ38jE7iqaJ8OVqSWVXoOVvR3uLW5Vxzj2Y27XFEKz76D0ZphG+KsASK8DeWsSXpfyvjOVI5V
vcE951RKDAaQ9CiTc+3Q96ZAu8K882POOJusWvhLBJNFJEhUmMX9vs4sltDWzLNONzmxd9tVwG5d
3S5RfL40iM9ztyoqq8QNmQsVM3rhsGIYWYLDp2WFj0+kJ1GkuNTD4v2to6fqQGUsu7s+oELuBJbB
7+0M43OhGaVIwRhW408gw7QS7r/77CwVnRbOAPCh28PngmIk+Lbq5ZyLpXz8gGyV8DyVgcXsHm5L
nc1uIlnTrF0nJG4kcuqM3MbyF1GXv9/vdzKnJF+Przo7Bhvivz6ee/1XltPoCOBRRT3KGYNwvqgV
SaityaK4+lr5scoVIRKX0KK/GVtIKnF9oYwVNPNME88tQFTCa4jKGVZjUp5pCE5/Ml1kRBivkgdH
HwSaSkXq5jkMYiBUImBwlsAmYwQh3ZP3tg5UVrcT46lZXuhX4oLM7SOg1a4y18M0Gx1j2an8H4Nl
LQuPTjeRMhhyLaVXRFUux+ZicsFUC4TikWU5urv85nLt7qDovFul9Clu4WMDn3mOWg7+z51yyu2+
yNJcP7vvTRyrbncPjfGQD9iS4lNR+hmIYby1DesIXToEH0EqXjsXMbZMWlWWarlEbaVh3D+m48m6
r0VJ2SeWryW5QLGSMcFUrtEmV9BndvMlZbdKBNqbFI6Ael2AZQWGgpnpTBh7g3spymSeF3qpsuKw
UcoNGKGU4npZvNTkPfwD8UMbaN3GUpBmiV3Hgn3upmNRHlLrDG3IebggJx/jTZRQ9I8oBoCMjkRX
xEVB7EPj0ztwV3wiuUbEC23pOaqwGyqe4Ixs6od5GtjajleEk3OVpGoJ0Y0gqO6PMhn0Jetxx110
JVEuYNgGq18lekTiDl6lMmJGTbRZHRlzTa7T2voURQhbBSkrJtxjdpFvwnwG1TzFphdSrRkftr4j
IoRNpnTjd7HDzFTUfBbqv38cwwd03D5L2vvS5mmegOniiFqoNB9A5kTBRZy+zM6gKZsuDYC/dZJR
a0OtahUmaMCEsR8b+9qeElxeq8V9wV6hsZ0TyjtmrGRXloLzOxAxBBASTLjmVNK0CyGe1udSREHe
vkPyBu2KOKJ8miE94hPTc0vfQ53zmyqNeEi1O0rmahlE1uCEUpYVW4Pam3z4xQmw//EGQknEj2TE
O2I6JyFcHsM2W2W5/PAzw9xkDhSzYXuZkdXByppQqMieNY7RaG9vzttsV2uc9c3pevl/AAW+TxbB
A4E6Z8nnbf9aAcUcPu49df88SaYj/+lmeHFtBT/uk3TRp4zfUpKKbTYPEuvYfLiboe54g92yYVNw
C+nwRmMBH3ehYiPzC4GJil4wLighAbyU7MRqMzZ98Hj/3T5sEXWORxxIFxWEZBPyg2hDxBf017Ov
PrsLDN4TnXXtOfW8HBhjXdNBED5aX562eRwTyOWpPJZpSsW+wwCgx6T3vYVU2Ri6r2DEvMFXqZuW
nwqgD3/0xABRmeh5RPbUOeg6QEmBMDpRGksdNERqj95ljJnvKhWKEJJRfftMYDTB0IalBmFUc+9c
4/2ru5rxk72eax9SN5XecVCDNxgifD82bgb7/oGf2NnKKmfVv2ndLSRSsMn/QjpRdbg+QnsvLEW7
2mngBKHFZbdHLWHm6Ytw3mEhLtzszfJ+VZlxYKDfjfuGLxU+ps4bcNcQt1ywcHKFq83BwlAmHDtE
hECGOF0c7lPhaq265gd61s4g/HnvOIv3kRaXWrO2f6zywLBxfDNdJiqIMOn5TRsDNVpqgoqKW9BU
rfedfaZStugPehodXsTWtNKpxOcHVyWFCUqEbiqfd84Vbk4RAuc7ZZinie2nAvxXmZQ97BTi/EqZ
YEFqtbUId+83aidJDD/NhJNgzsVvlQ4ieS2AzHzwWmMlAqDZxRi+MsnWg+ujp2ZG8x81ewlmwjjs
H0kaLpx7KZtXkPEO6bEdK6KuPJ1mTpAfqz9tO3mHOw+wtjPAxYuXPVp2ecZxNRh79iTNHZba33Rt
BrUdJRlSjrLUv2HvITl7rj6Vs6imcWNYd7g4GJuyZGXFMADlvDSHl1MA+VwZmbO9E+x4vs91ozLW
3EYgOCXDy9Gt6BPF6NSpWEsUjjAjCRl41r76AWkVKtg6ZnaHpHunjFErnhnB3pETFsQzO1kvQOf6
MH4H9sDCdtchHeW9bKUi2QB2lhSLdIn9/T2PxfTvJYQXUx7BerkHly0Ee/21J9isAh8K2i/ujI5D
dI0IwpOiAJ27KMXp2D3xC7mGsnsNjA4Mk8/8FtWI1bFLJuFM8RX5+Vy82CWs9k43UhedKbW3FSQB
5C5/NXbDGITJF0P6ztIypQr2p1AzJFThAfWJtkuu3h+3EAtYn2lNhgUw72miLjwKkGhj7xJ4nkH2
b5JnrNFO06bhoyKDxIjscaLFrxiGBkqRInRTh9DjHImjIFbc5gCw5KcR4c168DzjwUKnynKG1+q7
Ig2Rv+616J+Z8Do3D1CIrfQq/C/LJIf1zQ/pLD1a3SDeSHwG0yYANtOlcGkcSSdmnVu0brHAsNdJ
1xjSRBe0OY5v/+IJS3nKR3E+KVHLXI13U+3XkZxznIoVD8qGAgHjRKrAMdYLzlc7F4wG4zGb6T3n
2O1g8cNJ0iyj5Q4QmeLjsCntItsDc+GpU0QrL+XOUy4kPDYT5qkAwk0uZSKm1nQfFCtJgVm22vEF
QTd+M4qDpVYxnKpXZey5i204cPoM6VyE/BsD31oP8lyhskbFVugUr61cl7eoehU/zrNA8dcbC2Oq
kEyBKVkV9S6O70hOi34sQo537+A1Z1FKtMfxU2b5yd5P6ZHd2JaOkYgih7ecM5zepNbmkmeB/BsE
kSiROoRUepV8e4l8GCHymi7kHEjz+nkKQ8sEJVwhFh2ruuPA7O/vqvdPxt2FmfAtCrLB+akQ1ioj
A3ISCqGEG8LCRePD83hM2UjoR5zf/A+rsg6ktKTvmZNWSmPyGOXsUz7sz9NZhctp59Jl0/D0TGO9
tDJ+g+puOkq9d4ZR872WeH4efP96bR+6s9l6Oq24LmdYT+ggAIfOn2OBtnT413831wQmiF/rKGU8
NW6McvxMpIFhXQwzw//XRKq+iCkrPT2pCKPWUeEVQOoj52wSzicNVuy2AiRu710ttk0ahjaDShRZ
095bhPjBklKRjUAL3veLB9prLFr6OxW0o2Whh59YGeXkTrXuUNHe+ImK7lG6/GdDrHLmjhgEmk9D
gkZ79dCzAoc+98D2XF9SSd7BbOJ1AHVW+qbS3Kr32JIXubrYijCt6QddDEloys8jF27bUP4GenMZ
S5ZHl9CzeGqp46ZCIH3z3z3QEUK3Th7AQBCiB8Qy26xHITYMB4pSYRrWriVTgFm5uX05VqRvjFUR
AXSmdkoa+VshO/Q2Y4bghGKt9uC4Rh6DTGZprMkOObdP9dACr/94s7pTnu9/gryR6eq0Te/El9y3
wzQDrmEynNpEFS67ruA8uyOqslulOT8IlaF4M03H0bPAXpeSMkrE3auOBdgmP5MfiwvLp7Aef6d6
0Mvw89RWU/QTqUuewQ/uCzCaaHG6/B/ZbK0AC/Q3icWiEaj5iRVo2pDZHDQx8gEdVyxkOqlm3tBj
H5k3HW6lH9zYgv2RjrpuxV56TcJ6bIweEDUvrimrlvpI0JdDsWCnxQYd0WR58JkTJZvmWs7CvRop
FeC/m+HuxgfoIpOQL9GasYidsndujOD0EuZ/CNdWvigLGsbF0mFskZsJjjLwFSgx7VuH9cCQOCEf
+zVNpwcIERmVnPUiiEGWCqNHTNua6dZf1Ygpk/DAFf/spmkXDHsVToYb94bX3pU+UWKWP+GfvFXz
yd0CoyJwb5M8KhCcjJAQj0m3v14W+Gg4BoJJyubRD2rFdtoBVX6pWgXnExLXN6XQvN+0LPeUfzPy
7/7Ib7npi0AuJaGS0h5R5uMScM0cP7cWZimP1MiDrWsJJ8l/qpma2sjPWCUMHXiM516+MGhAyYet
TBSx8IiLof2qgxGGSR73GPMrp3Gsp/mFMI8EpEZpYvXeCFlszJjUXFl8qD2I+bctCltPBCHWD5yC
PSlyKu+u6euW4Q4tNQMwMDerGN+/AMhNNnSc4LS2ULcNSg5GEmUxtVjR6Zg31RjBznmdgq30pkQo
PjzRspfiqY8+H42N3MywU7oI2hfADRjrIxsKjBcXMLpKXzCNftXA1gmNxBg436GcYrsxx2+zPA6L
8vsDatlBHrOQbcWq/9PVD8eaiO7F7J/rqVcmV0Nl6N6wE+l1n6H1BEZ/C4TKR6ArK18P/UBYwBBr
ZbhY4+1s0OjoPPjbAesPi3BIUuz4fgmlztaQeoOxIVZlvaeeWc6X1kjxuEVNkhA4lqBtdCJldFS9
36o1ot1iJIHRZrqHEpL6KktHsLys5jaUdwCL8db3s+bb4HF9MwYkjUEWsWOoH+6YYHmXQTLGukO1
2nuadqoQFdJwX4W6EZE01p6ko0Chab5Ml7mJTWh9sm0iELUB08n7+NBuwebmM1b669NTObbQF3fx
6KFJ/i52ZB5cG2ikkVqx98sgCa4DnS/T9v/RZH6gR8iQfeMwGA/FFwe855568MeywQ==
`pragma protect end_protected
