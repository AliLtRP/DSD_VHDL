// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:31:58 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
gSvrJAzY3m7FVx2HWhrojP/WdNqrOqHfwsD7KOhPATaNCdji9r7xPDQ9UHLvr1jl
YNiGrSsmZbA8MqILgwmlHF98bjmq626NrEowJDXSiW88MgZfmfpzURicxCQWFH16
6WZ60VKlqLAhtg79e0sET6r4WECnTDfi8ZGELdKOcz0=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 6000)
YTtZ5IcxsEm349vPsAgy+U5MjYWyZ27a3IIv3ntc5oygsmgDyvysQNdHlFlU4SMh
w8u/go2bL3QCmcSH8QByCLrPbXquA/StXTMdcYMD1a+z6Uoz3VhvzdfrkLV5Z9jW
oNY9FroynvXbC0HVmnM3o/ySBBqt/qDh4Wgz5zqVh3tw/els3KILPSI1gDwelN2H
TrhVeydg3Z/zG52vqnR7hi6HfZwCSF3lHRpgzFJasOZxhz+3gObtrE941QyIx2v4
e3Aol+K5dZZgOlC5UzrSRbWP26PjSNC52Rz5g2Us48Ayv/7pwzOPxv1H9HsDz7w7
4UktmWudnutCID/Umj9bReICrNk6QC3h3Bkmq4qmfulVDeJGXoYOrGtgktT/ih8n
dmh+j0MVNiHHlSQvjSVKAUhvI+jGWfE+OC1tg9vOoYJxgEXMkQ2PuH7U/NY7c+Y9
/aJ/wkqN4Gwg/wkNcI3Kc0YFoxuZDZMDsndTEE+kC2cdcBkoHVB2OMNfEv9ki5mX
7Yj5WHU9ranv/VIFJGg9vW81Fc44Dc7DJh2mp7z4qU/JhHXpPYUlCl7p6z0M8hiI
8hlzYQT/R/xqSnf8EMyrNCTQT7KjX4Sz4MafeZvQBQbBYCHtjnt4K+HzPSD2Olg8
WmELchzqy9v0sFOPtMDSa0ecT+y3dp8jDVjVduNTpcdeUpkNNTB+ECCGIiKOUGhp
nFV90wYfUH5V5gRMuKh+4+ANsAC1tm2JcH1gExPFlbh4+cuUn0P3kATIbT5XvPST
N8Fb4EtG5BXea1I5pXfc2sImjknLJrZzK8hpp4hA6OUuG36ii94pDxlOJOpbHx+x
MHfaP/W3I7jM7x6d750J2YMET/N+0xPc3JSXhEe0HMCqboSKJ9i4gRtnWrpiFQJK
VkhJ5EDRjspiOo7CkDeA074jKID1LfbcHW6DS18hHmch9pz+aJ8EwL9Rjph21C1N
FRi738ofjcHF0dPMQZr8a9cQ36WSte6xwl5Ed+sBEPRWb0v0RyekAzefmovrfv1X
eD37gpnlTJZA5WC8//0LSAzN0PzZ5YRI/6BfM2HmtI2mgt6RO9uAvc1W68JWxMb2
GuUUGlbSkjsNYBQJfEXTW5PvnCUiWJxsnfsRzsK0jJ66KGt/KpicoFeuiEdI5F1f
9//c70nEYjZQufNnhkE7Q8D7dk7JkIAoY8Earsfp2YK8SBSyd0TcoY73D8DF1NcI
9GuIf5kk/CTasU3AN83roaiU5zZ4O3ANLMWqaM0s2eH99NG8bJpM4IpaCSDSq7nE
pO92f4oMf5tkFzMe352PYv/1fWhQgZboh+MwKaXHxWWqqBaQwDzGk0Z8hj/UXFeC
VGwpsqYj2zftYMsdg20TiqES076coJJd+zRsBU2/qekgMQ0pPf6B4CLNlhQBbiby
8nSPEAHolHWKD4YNLbNupKQ56z4ZTMUbSTDm7btufThHB5v0LeacUVNNY3Ay2FpA
vuNDKGjtkJdM9Yw6FMfmwlRd+QGXHueLNhn4AnmpyX0S05ml2O3OlNHeyMXToF60
c1ApP9ij5BUhnOxizG6Bgyb1mIqWe2qy4R14wmh6FwFnBJHNdDLU8k9gfSA5fI8I
/5y0cdmzxi1xidhrgOZG6Ojn9/XP/atEUTG9b9EyJ3T1FrFrCPq0GgOdiGm0tcXc
MF+CjEP/7B7MtNKadeZZ4R3FwNrbAFV/kNssLmqqLp42XfFS7OrTd8U477Cq/ZLW
2hVUtSnvVUkltrBVzEwYO/XBrYH116p4bN+jJDi4EZEYrdFtdtddndpLEsyJOKMZ
YdU1qWLvSU7KSoRVNsNIKppekdq4xNqsQkZIRvbLdPBOWRU1FyTQMAqYtnRrJm8W
aqB7UtbkPDz/TZNrk4wbH8FVN2Ncbm6ej7cEBwK5rXCh0fuvs41oKuOA1/Zb21IH
LAtrhhSPEFedJ4TYU5xh2/57U6c5cSfKpdaIyb7eI5jeWr17V2xs7khuik/9y4aM
ZZC+0ALRJQLFEkSczngBuzMz1tK4ImJCvXccecQE9A3Ao2K0Ll7fCRLM5eszAAkL
OPHpof0MG7W9j78HJZNMJNd3l29hMyTeQIhVgMRWkQVmLghrH6RiUMqhnyTRcr8n
SEyqhAB0QX821QtGr5+UGA00Qq90a+kU/EFA/LRoMQB+yewJEes4bkW8KfCxTDsx
/oy4KazVFX67QDUQWo7lnzBk42J2YXLX25SFyWHIqpFpaIdxexwJvYKzTiEsaL65
7JvvXKH9YR26y/w07RHk7UJIdfBqoBv7jXq+YL8pImulD76mmQgI/EkxCVuJlG2L
o6Db/TF9yFRlQkabIGRd0e0M/FZq+1MkowfAz5h43q7h060c9K+x8t/gcCUHD0fj
qWivgkbK8RAt/uOkrOEEv2YdNNU4MoRvk6cCp2o8VOklaKNp+v14AenvJbdE71sr
bNF3EfqtefdQ4D4g+RbOgZ2TFSRgmyFrkaYPXAghGPibB+Wicp9w2DoNC2GFW0r+
m14ZZ56651eMnglsNG0lhzSzPEGPG9vmZDSzLrMReP2LKEZZ+rhRHEOwc5PeBbKg
2DjTyy/ZtRXfrai3Bbulz++Hk6TsilrCaSOow/0or/vcgBxAMIxUXh65bTY9pT9k
RdxEw7cmVMwf1xojPhIf+dbahBmKqRzOMUNXSswxKPHkxGDSMaP4OK1KGm+yKQPG
L+iRrKfGls0ijef2xZE9IflasXB3p0E+vYH0h0xeojRRK1WCEvBCflx0GQvaKpql
tbu5/ghDxupKw1CBClqWuMWW2FbdheJC2rxr6Dnesv8Nr+8ZuxGD4JzmlSQsZr8Y
EK3ZFcVnXO0PCTgntrJcL689/75gsxPWozNfU52S1r5iDn8KmT0J3M1Jkh4i4/n6
CvWkGbMPhy8KiTl+3CQho3IMoPU9W1sp61RdpnoIHNrSfVpp0fVuJ6GHu3u2WUdH
nnr4haz5fbRE7uMpfnsF3JDcNEtwk8Uvt59WnHnd1JYQZtnNLFCKjsxxbO0JPjeK
xaSnfyRTZ5zeq8a2InAPpxXDLVPvxLUTSQAgmpv5XabTnLSkkyzxhlfl6a0KrTyO
obKN7jC4KSkwA4hha93F5RUWpt1FXk3eKtaFDwZakVVX6I3T9Aneghv1NScVySFa
jrc4UXeRbW3hWRNi0kfzCqX+EgvWV4JZk/QSE8z0YFwl94jC7+lw0Sra2yi2ARv7
XXgGYYUjfScEjluh+uY519BNwL9eoWBRKniPqjnEaH8vlO/D+xrJlSu9IQ0wAX99
xhqyxA+KO26qlFhvPumk/r2yUAnRLhtvUxduQCCDJZCFmZCaruR6Jll/F/zfk3b8
2NBPrP21mxU3SuW+6k34vn5pL++IJtn0PCHBC1zOwNhLAiJW4w7T9SS2E9D6ZSeb
goQpyKMvfQyUirI6yOZ2AfYmP+WMV3WbfqEeoNxRwFXUIp7VWWBBy0diElZarxrh
8ABRm23R325pFY//KXo4Tckje40W5B9nASUfoNm0IIqQk0/u94NfzZYgvPpKJ7Zm
6S/BdfMpRwNsTA+mLCqZyUW7SWePXEsTCVizrCpBXHHMKKH5sQjjnZYOc4bsdmCh
3euea4hw580FKr+x9hWOWC12vo0DC6b1bXsuTX/uVBDUIUcSwFoHn2K9m6fuT57e
QNqK5VwiBmVsLez+Q+Vg06NY0zO40e+uXxlLkBjEeYdDWM910IpnWvHNETfOd9Ae
L4smODhBfxf9opJ4MxXYjD3QPG+sZOFnceXHrBqR5+5fNjxKNybEATyymlzDcWOW
PwZIGcGq8vNX3/PE7nPI7ZbpNNYE3Sl1tS5yvtkE5PPihWhYKnViMQkjJLW32HfV
ZFx8YVJ8kRtUkFzf/KDGghy/aXHobW5djNKhRvKKvgitLYM7ZlPIr7BZojeL5fDi
NOeaPt1iowwJwN8HVd1YLoOyBKCDGbkUtXXRgC1EgFJvQLOVIFIsCejPmEOEkIto
xR3qB0E93CA2Jx65nwdcZX5ocHXCCTjULxcjbgxOqBNGybLRHwEQaZH02czFT6rU
hhF8WAae0xQ9t7D++H8S8Tk4NAh5v763+YVZkckEU/1uHW8otFWyXO7906Fq6liC
eZoOsr0H86krg2HdAeJE/EYdZP7vwyVgnBEhgYkxoT+lSYyQ5qzfo2TUgogOas0y
ShF0PtJg+Jqb8ZWh1pq6QUH1GrPd+ZdgAWsC5Hxm8t2GjxDoHi/5Q7/4yz+EYt5A
nw0HPN8eGLV5+UF3k9z2udQH7pMao9Wpio6FMS0GzGn8nWlGEAblsY9ErOKAfaTI
w1zyhQ+rCK6B78H3j9l/TVJDNlQVt+zFUyZZB5Tn4AH8LFbtr7rhaeNCCz3b6nF8
SPExS6JFW7bNwH9/nbUDtHU0vsOSsOvBNmRq3biimqn9kS24LLOC/Mqa41+kbJ86
AhNpN6dL1y1wlRF/4sR0P+CCC/AgWaSK63+W0p+V11ZOqtlM0cvahIIXp8fRZZw3
2VSZXlJoyRVqgpd5OJuw2dVuzXsh7+N+W+fqQFOlixdfXvzEWiPT33TmNla8i8Sr
LiW5dOqqjUyEY0ZWqp6EezQYn6uUcX3Pt0BGO8iCG7M7JKA3lx5qRloXmtf1C/I8
7iu46K9A9eVEMwwYJwM4xec0nGCWJ++QEbyhg599WDa8/u7AhlLcXmn70CrKkP/z
dO5xy1pSdZZXE9IqLdTIMyKeUCIKIt+8VbWudZWpOWesGm58yCGhJ6K0pBTaIgny
za/uQ7pWrE5UELVsxKXdt/BgkfnZVrZTvfGOFhO03B0Jp0I3fDjm7f9e4NvSEVGF
JBlKxIrksR1ctW2B4Rq1GgwvQq90QrlMS3wU2LE4TroaNdMr412OCxL2AMArgDJ6
7NuUgaPgCku667H47JrkpQDyknFugQBTh6EunMuSOdUsP8gYo8Q/nHYibg7+SGrS
OoLEDQ+I0xWtM5qxZKzVqLAnBFEW8xq6XCJu5pzZ/peH8M/o+V2T8WH2zG2pTh2/
ZGAw9/Ctig4nc9ruYCYbkiuCDwnVFK5OO87njWlNyX1xLJD+p310RYvEOwMQBtM8
KZPJWbo1LYwyTh72U9hRkYCj1HSjFPxoqVpWPiX7D8Z92PGvil37RMI+c4UFfra+
QEYl9tah38FKkYcPzmxlq5cMXd1V4mGfaBX3EEYWf/JJgU2lhzOQx/qvLoqlwydd
VTjVBDAFvJoXWPVHzHFK6PSwt3S/OnVBGW+kldME5EgUwqqaA54u/VuOgkP4ECsu
FD9yFymdp9+knq0kDxbKDrbNQJnw7YTBEeKbmNIi483BQpaHK8S94AvwnGF7hQIn
gdrrizUOrFK45xPnYG+wQysGTbfDcRdkdFKh2eQVr2/FDtbPsxf7a0Xxjp0g26Tn
lY+zwaA88cbsGt2tbYzQqZakgv5lIe0loJOV3q6uUQhf1Aj2G2TQzqU75uvTgx6d
lSoVmx44tIH5sZ9+HNsj4ahQdshArYvxUhvJy6aDCTQXsQova/SjtiQ6GUiSy0uk
HO3+n7AsQhqI79U53dMvJup/qyPKRyAO3PNf/TUxhw/n8u1kiiPuHcNQhyJegxru
thl24FiVgGMfZ5PQ4ia51wvmmxijl0cge3vdwPSdzl+h4rqqMZVf8yI48444CKKR
KyIuRqRseXP9lLccC7An0mKjdO5DDRpbFHIjdg9AZgxpRGW7PRsXPV+30iVP0PK+
JYPWrb/3qZHerfbMaCUlDu2e3+FjkGjkSq82z7ocupkk/XkJZS2faSVajS/0GJPn
JSOWqi1mzg3qTOKSCu+qXiAFQ0eXhbIFs5zql6JHUHMabxgEDEi2K4NSqQKmzfuQ
cyF1Tm6c4NYr/ldtrInUcTeBhO5Gwf5lPdza2wpKik14vGp0bzN3H42IbSU/Z9lP
U7SjwE8sb4QsU6aqCyZ9Aao4stefbl3HaiVrTpkDLcu9qzfSTJEQpPMowp9KthAk
ux/5CGpP/WrtrX08OHATIgkU+nW9JTq34Cp5hWepjXRy52nD99SD0MNTMzItiSVT
C0zmABnvXsK2rViZIo3KiNe6EgRpAAFKfq/HQtHECtT2jpWIglj8cGqJNJ7R84Ln
kp5H65gvHxSvGawPVFxQaDItFRbxq2FzAZYocGrFlqs8pY0DVChkzsY8edVDHNxu
8vlJPgwCxG3+H4vAfN+wDIh4qfJ0pT3jBvNVA1iZ81LsfUQtrDoElvOzOWGJZ5Ta
/nO2MIKOoOZLpSWaBDNfnMMW0rzB6eCIxgT86EJtPNKIKbrU9iYKW4ZWU4B1wHft
9rJNrQ6WWG1FzDXtuoBySq37Q9YaeYuN/cz+9mZDM/2EDEc5O3ileez9GJOeZnge
MgtZwhKmKsq/+PPLHsQkjscfcRPst+5NKTszVTbqHmj80dp8aCRUdYoDHqbLIaPM
ZSiLHLm3Ixk9FmdYbCWGYvIXMtTmm4wJOJ2Jsb7eL21B2IfOcHSVOKEecajUl9ds
S0qAz791lTIUJD0YxAalCoFziDC/v5Yx5wyjeAaL7f/Eon4IU1zoLwv6HMzB8EEq
kcNtaAumr1bKiBy88TZWpuh351ssV1U/kF/Z6014DhwXUWViPKKPPqviiXqB7zq6
b0BWeDnrlr8o8KaU5DZK7Q9Dw/6BErgAcehBVhrTYHdr/3QGnX07vCo856/72yEB
p01HlmnZVcqcBF6I6Xa7oXmzGPo2A7gOalAWQ5fx+qer7H8dFyQjvACclldppwbu
4YrYUBIY3UgIhl9uiH809EfIWtiTyjI+lF+HnXMOcbpsuhlN/RJndMkA7jqp4njh
4CFRqVP0PPm4DjmgmdKwqkD0QvCXlmwBYjtDH+xks19q8kEOtbTP6U8Rgs6OXo5Y
W0+XrJue7wuJjPWUjbRMvgc3UpYsjOSELV4YLLVFAHlbsopnMVpR0dWuubxWB1Gz
mJpT5ARuHAdSw1njQ+65yxWn0WdpvVzCTtonsANhR8vYI9l9Q+/bdOwnv+ubquWu
fbkdtEXnQljPIM99aF7Tq1D3bCX4W6aeMPYbjuy++Xs8fFYsJeq+xAI+AmzlcOX9
DgcYNrWpSrn/d18JsUO96jvv7C3Z+xhCmsR48CslSOZd2SxqTIXv+9Q5iIBFVjQu
r8J2XHijzgYj4kLCjYuXZ7PfvKYzoqor0iRPprJVBoA8xYTFNICyZCSVtcb9vKqf
x7UnjMOge6IFitcN2xK2RlZHTYQYsi2HqBug9CMId++rK0csk4qk6OIWCTE28eoF
Aiadg4Cr/Usal1+9c+TwQXsUfYnwaAyBl6FLrr9D3m1ULx2accH8QOQrrtN4/wOH
zmWUAUubhqsCGO5k3wvnLd33IWZih+zmQJlUbfJ2yM+K7Us51AB/6HGYbCNA0bGI
c70PydMlXDba/VlvpYxiLKoT12bGgSuJs+S391CB5GCFScK+TBf17CaZI7B0HoSQ
fJqdWTQb5g5w71P0hMIx77ilaEQsVwZJVfgSS1yt7LHAOph5Ugot9vyjWB3qaUdu
CtUYcrE+kRPXnaz62zp8h2SMV0JPsXKFOYq7cI3Cjv1FECsrebXN+VuYN8RblV0Y
xjzU00RLU8SYfHyWgZaiZgXce7GbR0n5MtSM+2KhTkgBVBKd3CH8PtEEBMyKcIze
vpA/XzJu1DXswGnc+46EXiGo46frtUvIK7sIspSk2jbJZyiPrIq+xHN2KnPzMp01
0k0+35GgYiq/i3qdM+Si0jZLr7I19BTqigrqSrsXuzxEDDL4qhNOvMMhE8GRY44V
/nPg6eslbuHZWSf6xCaPNObsCM95a57BU7jEuM0UmNtsB2Mq9jwF4xV71xcPn0ME
aD+XDbKyGYYzpdL4Nv26tMcB+QDkSNinkqyOJ0tYzsaJ+r8/l8GQiCn83vmN9NwE
8jhWdc+1WEUVxho5DVE8peonEityZSYppkuPI2oDCo5O5xgKgFCzyQ9Uz4W760lV
k0Ir4/KvqT5kVxW7XiGclBDNLUCOyadtLWrirhzauwYWj7nYhkmpzRaWiX50/p3s
`pragma protect end_protected
