// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:35:48 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
fFTD51pCXPyApt6Ouu9oYHxC+OwGeeDLDgdzqlCBM2jCScOcTSH4CylS54xIxk1p
PU4xzHrBi8Ah+qAjBtthcm84huNhwkGhbuPPiCSTfXockprCefpqUTNKO1Ha5j+G
+N8rtuw/LTlvsDsKc2blWIrCwSu46O6uzjVt6jW2XY0=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 3136)
Ao2BLd6SPmOXRpzO+I6CSMjPEqB4ulCXDmBbq/H6IrrrHqZ9egIBmLIvxSUIUKkG
Qet4/3nUog65qCxZIt9GO7buDIfdSVSgBKFopa945DKtuVhIjg3uSQjwVMidaSMN
/b2FRvjMF72MD1ppOX1JAxRJrIvHYd4F/iCrU07M2aLmD5rzQCVqpptBmlohaEA1
RTIRkN1u/PwBibYrL4KJgHfQuOWGX+ERkafLBBDoQjA1Y0MIo42mcXQPpKf+oFrx
xA4odVkM2FmwQ5ssfvF9QsrzGZL4WJTQpqSsJlMOfztSZutW46gqANEqzYjtjmXo
LfaKJOyEcmtVwglcolHebuepSogrEVFSa63WLLUtzJURDYMttlfOPj45u3AkH7uy
tQ0New5cdHba3KSWYthQCARShfPRoQPcRkpKYlAQcJpDnGVrLqI3PYe8fBXsXwBN
PE0kXXl6WnUCss4SxaQuBUw5RdJRHOc0y0e5FkcHSxn76wfwXSAeTY2BQBXkTbz+
jVnKs0bnkE+RzNuaS0niL95kFQmrGmCVLLwHGqZWF9vZ/mporhpLq0kA+c2uETlA
2M7d7TRVhnVr/pOpBK4MjEZyuKVozbDjeFmSl1AyALeiE/onKxfZaLPxdeDP6trY
m16FPW/ajuzxgGL3STvdicZ1rmOflvjJjSS8qNU7VKKzQBXyeM3qeo80d4nQEG3s
NjGD5rVszcl4Ee3zuTYi21aIM9qW4FEMpB/bu1TvtIK1xH9dFLiRG4A6CSsB4LMa
X7+yBVA6tFUVYG8LT4YQZQfkNoBj3WklGE/1w06BEx9dDfuMr4kfV7EeN4dC1jLK
JyxZhh0I0DN8gzgWvN9KoWzygp9TBeuBzjUOVbEW57sZ8zuGpzKahdS68t4Nzf2X
ArzL4COXu9aMK8bc1PgYMfjddvZTJ+tH6AO0QJCNgPZxE4/4pfuXDvUvnMadxQh4
I1LXl0kPX+7YqxUjSeR5DRBuDL0ipqj/Pk32ifuZqa5kit2BM6oA8/WHcCA3wmE8
naTQZ3OQr4jVOdYnj1CnlCWBlDxRV8AVA6jaJhGhEGz3eIhPsBjYyJ13iVHEiFUA
zsAuIGJ6pZP3yCwlLdGrMdWAbudvo88udoKWUonf+blolVzwtjWkcSG/4E5hss11
NhZJEJ3uejtc6a1qzuCwITupvGFbE/HT5XvgGKo/o1KAuSJnRZaUdgoUiV/sC/6E
o1MI++eiacNmDhpz7g3xxXgomHnzW4fXCJ7+jp2Q9j2BJ0fULZp1dguB5KmO4zFL
8JOJPVz3pnpYDZaFaAas7rpaPrXkJjiAXXRh1nkcFCQpXD4KvhWwB0TGuihJkQwd
tAX8sHD+AOLy4QU5w3ckjrXdHDrGciF0n5FAnLwl77XmgZwkFLmTuxgTvoBH1CPz
d/wOQ7vFsAOBzMYIP9IVjrjX5ViPloY9E/1N6RjdLqODP+552ts0WkjLFnUdr3YF
OLh6kz7Np5EdZuKg8fVp6VLmz33LD9oHF9s8jvKmDmsTbCutp8DixDdgANbb8crW
Q+kXRRO/KvkzuAg2Ec1mBpYxFsvnDPTkCQ1/pgxNbfp+T94ilK3ktUrG8N+34SU7
5rr4/eOOTN8ie3w38nvXKpy/GYbfUOvCz6rScgq+0ojW6XudeiTdbiofMiIFAVgF
3fFofNN+a0lcTlV8ZeBl1yVQ3mZrwp8sdiiqauKp+S/kgzlzBoWqS7MhoeWqkQ+G
hN+rnLlXEKV0lojVSZdVqKtlLzqtzKx6YSNKrHdCBdoQz5reSqbh0YS7NQxkeCcg
/ZCmzVyJ1eRKfimOC7r8aT5rkFxbmv9rg1HqZ6BJUNwVGeJk8Xnk0nbQzy7SfsK6
3jP8LmKhRpWgD7/bdE+Ajmsmpea2E5hv07SUdQLYWAhqk9izRxTQwceL5s3lzMR6
Tya7xS+UOaTVUKgZZf7QIbYrJ4/EecDa9MePvKXVTVRtb/2lHCvG8CnkA5GAOse5
KTvXuLbFqlH7vX/FxyTUTfAO2Ii3aMUu5eJ67Raenoq9Jsyfa3hIvLgydPZz1jI0
FzJeKLZenIfMa85tV58feBRb6OXzKq01woykTXsz2jrOblIacpkAiLgha3dkuAe8
mkZe/pHJZVkJFVZlLJLCie4nAKj9ymBdYQzXzgJhTzi8yXL7psgHv414EljTLcRc
p0ixSXk5YNy4vHkGrineP0PYhT742vkyUNjywPZhRgDUR4nnTrpGFiUA0g5Hr2UT
9bs6dgKzpgcQFEUm6UJOTf6TRRnOwNjjGujKUGDdF4aJeLFGqsUo/ihAs23UeMB2
kSXACv/C23JBxdQaR8LNiLfghV++KYNW1Nn0uxyXubPxaO5mX6uvUOBcZZGEzhnC
k5XIZTVkub60NGe40A1pCCMP9QqG4cDpsiEErK2YXWW7vsyxr7R79N0wY7nbXzmV
sGGms4pXaCPSLWyJlLtGIVQVyTik0OVJGIZHAKsi+/3FaQnPICh03CP92auGZsXo
vIkcwkB9JPN31LeId0e0sQE9/4PnvedEkFkP++d4jSedQTr3wpzwYhA/h660FJcu
ikPBiPC3K6UuED9T8t0nkrOJ5gPUYwfdJa2OYpDhXLZWhJsLBO/GiBDFYtMUCh0T
54Tgy6stPJ/xZ4QsaHvU4xic5rLwpkz/wk0rRQ3PUudc0NR2G9xm4TdNwfckoKQS
LXhBpzJiCGiL34LGCTrv0i6w2Cjbzw94AeOgU9Jtl5EfW8NoFqpb2c1SwRXwh1N2
qvqHFBCvQ6Fru/5m02SFvUS+ZOo+3Oxq9rFzsV/d12PcAyYBb25DYhCcyioy8JMO
TsybLzZ+oZIjBpGmE/asyOVOJfRO+uHaWOSPrYfFjBINaNs5ohMaeaM6pp9envLX
2VVb34QDBmlwHlfFM8NTG43jtAiD61oDN2h2OVH2OUnZPQ6hKu5Ne1qdHXaXTT/Q
9uWYEo+3LM/nZspnYxXWtpTnW+icpSNdDp5S+rcsgO4M3hFfpckcrMSiqm+fPzij
v3/P8sc5ZI4o6XAormOxQyUKoJ+le9vk2IPADZbpBP4pbNRbH2oze8uUmfNNJQ1w
/TLlW9R9S7fhkwgS1vbnEJ9fo3J3VZWQyT7lJoTM/golcW9ij0NLOfQi+UlHka0A
KA8fJ4F83OlLkXmQTIw6/iUVp7nWFa9umJgj41Fu206NdXgJoJeCOhGiEDFzLZNV
XaO5LqgZbrnGQMLUADLjCOK3OjABgn/45EIypXnIAhu9XupUIsMGH0fJMd/vj00+
ceppx2/aeDVzae56Ut73zCJsgaw42vhRN57GLIINrrJRjPm3mo4JF9jEDWulQuUd
4nAfQOMddjINH/4QO4gcLA2YYBzMpiEG3FLwCGYScf++jdid9rG0hwc9GhNJuy8t
Ror0QfqGsyjh5C40YkH/atZJka1fJuaLLScqphw1clT4LZKhuHNf1aHhk9KCCqe/
uoF2AWgBuJRXyYfw5YIOXOrYzwahMCb4NNFBE4C0XK5HGA/fAldFHwKN1MV9VyWP
49h+nOmxRq/fOo5Te3QkDQNGO5q4BqcsLcY6CXlVQ/ip3XoKGtPKlBcQ55w6yMkj
G4SpiKtOruhnfLzupk4SEarT3Z5aIqWBGqtDpkGZfvZBeA6zC9aie2FfzM1PMGwU
CDxcl2QzKjEA0HczezSnnhyDcRBEX2ZkX3lUSZMkg89iOtC5RWo0hrqOFTjylwE7
xyGWRPsZsNVZr3v4kyAZeB1zmvo38YMN2X/wabg9jwFjqKK78S5BIxrqFPPe/Jen
j3lMemnEBEvhnB5ZaiQcGSkOnouJBoV04QxbJGwsyKrWksHKvj0v6lSO3rGxb90Q
kmNjPAPzu/+sP7aVw5wS62/K/MlfA1nVDHxTPpbiyJYBG90WmqUhsf36j5uRRlP1
3nVn32YAr7boH5p9dTFGc0svsbYSntYTurJSrqEpxJWJLNgEv8oIPX44oUexXVm4
sw2BIgk/Z0P5moVuxK7G4rK57hq78gsqeAp7kkyQ7jD5whM401FbIp0JMTiSEIAf
RPtzmD+GRnJh7mdUz9zhVjaStQmZGEy3VsPa3S4Jp6trU4YFER1pRtS1KXy3ul7W
hXlL0GWoVZBhIXXuYUWzn+UfaQEOo0HQMKY74NgcJ/D0ta6yl3FvUvgaK4xMPQnA
st5RCFGjnu7QRiF0fp/N9A==
`pragma protect end_protected
