// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:31:48 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
HBd5wesxrexPWBwjYERL+L0m6vkJ4gLQ+yKO+P8X/0jwurgqSlbet/p/Of03/rJA
qOxyP2p7g9zVkmdnHovDy4LQrjP2a/h1QChTadpOGud+WSVBzxL7fWvptl3TpSLb
vZIfhBNUQzITUr8+NfNeqrxE7fmwSqnbaMnc5FfaMZk=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 41440)
HHEd06X/jkeYykCBYgW3SgIF4Lkk9Y0KF4QCgffeFU1QG+dE0uOIFn7okKQsFlOS
SnBtnqWNtVsURz2079luCWpZ3RVOgPghjWLHVFaO7p8CleZUM7ZwW2Jcn6wDUsgZ
RNb6k1krUouFTWTNmtaT9hKm0vIG8AKRqFhPb2/uAzV3eR9ly11DKaNMFyv7nfk9
GZjU2Y/XXbpl0jYnb4pOVFBGvv5XxmSkW1M/owxOni3T3bps9q7axqiOo9aNwu1X
bEJb7fM6y18z10+tCLNScmWN1+mIT/S7eBDA04gNgLih/crVxMzZbM1NGR/oIJMP
Ncsf9NwArQzShVhEZR7dGg0yY3fMPhci6A6HgwPvPdtCs6giNdf5Wdvw4i7ZHHKQ
BSRLmqd5x4tj97J1QRQqJA6PUFwlnrra4pBCFrzWHy034pZRXTABRRjQsQL7DcoY
PuLSXvN1RBdaa/1DGc8fxpmY+czyCHb3trxlIS2FGVbZJfpljbFXaijtLF49/s33
iOuLJJQfUsLsoHJF42Cean9m1lMovhxDvfFFlLOBEjU6rq6XsOVNzpEVXSziQtr/
m8csqOS6LZYWdR8QINIoRyGeNBBqo8c1bsTkLhoR4RI6wMzZIkAVcN1saJxaHhJm
7Wlep+xAd4ZYgvff/oALPwtloSLeB11SQP2gOlSzVIBcsRmkjzNgSpDOQyAaevu6
n3XVaevbimtH8wuRgMye5H1mefDDVOeJwPInuFVydGEKnYWwA117c5hrZU10r/Sa
NyCu//HnfSWYLSYBxlnQIukT3P3edLOYLDYts+xBMJt4Y8/9W0WMD2p/FA1JQJAs
1fsZOvV96zXnndVN+NlSeA7LUsBACJSgSrk1LfgQkpSs0VulkBXfkQ2Fa6Y3sr7Y
eBNCPYRv1KlUIIcezI+C4t6wrar7dF7WHQLtDM5PwWZvQDvTV2Cxd4RL93wdfXpz
Oh42B0v79wAyURY83iQLdxbgpk6T663k4OerQKk6gDefLOWiCNNCjHMjMeJJiCjD
miUpgDuRM2x9NlV2BNtRAkVHCInapXCR8DKtBt1GcvNgKdgjaQxZWwzNfa1f6Afp
YMJzelA3gjq+989efwUtMVnVcX1qBhXpjlPL+5nE2yo432ymf8MpYQUsxoC8oCe+
9oepUUKOdrwX9T/WQoHIVlGbrYvCyMBtjPczYV/CcVoSKQYLjUS3k7kDIXxmTXUr
MRhzUtc3OM2fzlMShuJfVIOT/ESmfXv2XGfWIlImlDd7Bf14IFc8nb1d831/v9q7
LYN6vnfaB6PW9M2K60GLZ+Oq6Qq3Nke239oN2t+b9VeqSzU/LIZKMuB8vMWVQW4H
ygPnGIwYulDbwRVkIL1BPQBPFJ/vweCj9RQHCuokWNJ3H0ymHWiY6icSLyJ9UpXG
X0yU9ZWSWYLDeNuTnqzL6fUD4/Wfk7IwZmrUl5/kReLZN0PdSqwGHRSa/pPMBz4z
RkmkrWOQWJBi3+S+xir9UdyQvPDNmKWpsAIJp7PrtUcWQ+SXE9K0e/EdB86u3SES
KphirEtDJsVm8yWi8ytJjaG2XaEPRerPOFxn0YP3k1G00/NAAyuwiHt2VC3jLxMA
Fpm89rihLhiWJBa3fkdYqGiLXl//h3AgrPbo1EXnnQCHGgCk7RkhTSBO052aReT7
QnwKLPq5cnzfHgFflHMLAERVUMLJik3RsnRVL/wRi/0Rb1a2FQJoBtTwceRmhozV
f8zDR061xFEQ/A2EQFq21L4TL51D9m4SAfGoG6qbBvkZ6sWeec1Yr1qV81Wx4Ciu
vWoAsCVOP4mHaMJNFyeNG8UJsEI8hLpOYfL5IndCivpFkmGKQiV3atZk7jAk3E/p
mf9M3Yr/qDD2bUXaGs3tjot5DKLDK0BFxsOoIyeLALfK96G7UXtISwhXMWYxr/FZ
PkKA7kLpBu7OZIg/Uosbrt85Q4ylonv8X0gKq1vFxaabVZg1eVNwOLwk+XcdZeKB
Wp/bRIOTJ4BpCMSLhpljjoUIjKZQGhtBjFAohAPnctDzSleq2vxro46x9nnfJL1Y
Vb2bGcS1N092qUUGcWZSFBS2Dm0DFNFY7r52LHPpl4lXxVzpBsR8Iti2ZgueVCaB
yr8UgO1dsfSDjs3W0ll94kzawB6hzqiQ+SUBHNPcAEnQSw0PkdqKUvI04bkRA+Lf
Fq2QhI4hErdCZYDnKQ4jgYzIJ5WT71o1CGmxwHnUaxw3QA8EQH9CeYMNxKy+oo4R
y8KA/4yCiZC0Hb6Qft9YZ3Kt6DADVnmwEeSj+49QHMv5Yi03hbY/vxKxuxyRfFd1
y4eiHwno3DKiU3esZuM508KoCn0wpZVpDnnNsdtIXW2fPiAjxYTnqGZHeKmH2psT
YxOz0bCrLk0c54gYp9PLn3KzEuRruKalNJEDtw/poi40HkrnbOEhjWxI1yLS/7MJ
sA4H6IlcDHU6haJ5jgdCB1OwiBDOdFf8lfeShE2QClgDRdKxRGLvpDLVNC2ZkfYs
Q49NUPyaDqp3KQensRW9DvpxZJSAvJJSQYLOL1qNx8cmm0TD7ND1PAv/mPo1yWhV
+Yu+PgcrVrVFH3DjXlfRe//qLcKU0eofvYh+2EjyPKxaJMq8W45rwwcsx2hOV3qF
iPwjlMe56aQm8+HquBeYj4SZUguNeyF6PbzTPP46V1XpwkogRPM93qGrQX0iCadr
paYIM7axtvZspSLF1K9Fki6P5Ucjbv0Rdi3DjgWaVUtC14ABDEeDaOCJOsAwFn0Q
ZuIwWQJjnFd8f/CQTKoOHDbkbSB+cI38CT95YbrezowDTXCstN2YBGZMqKH2K6ct
LldQW1aRPA7z32RHAqVg7tMyUh1RGJCvp9e9XjoDladbWbLcbv9btRoHPlINzS22
YdPjcbrkurHYNZc8tTNizA5BTRscWzOlBdBbTb8SQAIuQyUxwtgdVhEb6Ir0q4Bw
NzYIEw4Od63GifD7/5swklp1vbYql5XOIOSbVYbyyStNXV5jNk050wQvaqJ8+6go
YiW1jcBQDVaCoPsMFgkUytUFjDAREboWFYZBhhT8n8CB7HpWDd1BtxjBE6qVP99k
t/ju7v6lzIUvIS8DsDk9rGKh/+2EbZBlB1Ij4emEA/bgdM70IxhpemVhQ33p6raV
xxN2PVw6rCzxhM66T7uduTtf/2yFOxjZnNS9iEEoi9Jja1kfEQxYA26moOGpXZ3+
uG5aL/TIFrqgyulMdJkJ2UtJ57AjNPe9U5ev2LFZpaHm5zjwDwt6WzBpBzoF0sET
2xlGwKvUYDHCYZjZP9T04lo3ZLiVCVIx+5wpXGeSFZwBMxWo/hzwO0ZKUopcB0t1
T6R/fHBdROcxEGByiU3+DavGlRGVI+ESBuJFgdamAze0c1OTE5DO8lUkZWksFib4
iIruPGpMNrexRNcmlClj85VcU+PSUlOZJc79QGSmlOIdEBmG+w/qd2SFVlv27hXo
UD3RYlRXJxzV24GP8Xknv66N5DdUeYmt/713uAvvPLCWk/i4LwNMM1693+BmB5nx
EWwTbqg+Zq8Uk5kwiUqfymM6VTXB9Q5wS4gvczkRwIv8ex1rPoQQ5cyPZHM6lRDi
KodASaeGxEFr3cY5R6ayWcQoMr85LFUOWd144uQR8zd2LPc0l3F0CDLF0YNrNTyt
vGb1Oj08YdhKdqAQkzBuDr15uDSH3ig9d7YPOrRrSvwfT30zPGy6HfPnYUz1sVnI
Hk3Vr0XqNItQDuL6GpIyzFnK/EnWTm5fV3CsRwfJcDFueMECzuFCoj37R/wIlj+m
TDfjKfx3qd30Yi+kZiaiBzXWTJbDrnrO8oEgvyZvE2MuVc2zI+aU6iIiP2X6wi6s
geFBSyrezibWfKqbORok497x9am4OBknsSSjFC2VJb5stACykv9ANH4ybzmZKgJP
ufOCGBXl16kWTBA9wxbMH6+rpadsyxVI/g/E0A1EMY9h9ABlqJo/0fopZjGKdJ03
lrXs3eGRnhY2ZU8dx4tJj/3WVIy5aVIRKQ6GS8NaOSQDnphCliQLPZsNFF10YsNp
zJSab6xG7dqrlB175L/klg4jBvYQ8KHShp03dkMipw1RC2y9qdHFjHEeSqAKCsVP
llthhmPeJbvIiWiv8rSScsMef9TK0cmXtbi/G+vQ8YKOyoXCehrJxaLrzRMXOphu
o4nbaq0FhtxIrkMl+KPCga8xFaqvGO90Bmi2hDI9wDvfZZ5hrQeaRdOts5QY0uir
QO/uooaD3rHpUjyLrc3e43UObEzjzYGYuw9JIN8EdrbMn9yBkWeDdOLY+EyAv1yA
A8P9vGn5bsIPZAEoaJgx57nYThtui810hLB/u3GmyRnbnyRhbMJ3PAEFiE011ViA
KElB2AT1W6JPc3CF4fWZsxcM4LFwDUt/aTd1SXsOudhCrI7XptgViXSzm569LBoB
ET4fhfTCrKol0tsTGqjz1XitO5NBPcqCjxCt3Q2egnHQv6Tlnl1iwEz6hDs3L3Ux
CIopBl6wWOM3b1hAbHFGLV2KiiHaRoDFY27vElL5N/JJ+svUxp0jOeWqodT2XCXS
sdswFaBeq4/ynsUpAF0KEHoTkyuHGmC0IIzTxzTZkXcxmDfKuLjTmkjULLcCIWLY
olyOZEz7mJUAGicGh3UZvwEy9uIsK3GmuEcHOwiPHfmfahRExZWNxMGMXWe43MD7
z54IY949s9EbV+qnQSoQXxqHq/8Uvy9u/FsXBZQKpuC5x6H8JJPeRGoNnbs71SX8
lxqeYJ7LFdR3ym4gbllNf7ru3/4gm4831jbYoqbUFJUOB1XC87+RTXmCUqfPJ3n9
3GoYekjrLcium/UYNicz+29KDNYKW/hQux6KjrVk+WRllMY6cyWSH1SSpDepto60
NoEJS1YwkQ+Puk0eUklCe0EAFjVhqp/ZLuVymfp1yO9wZ/cUOt/frnR01SYCrMWh
p1+tE3qxxbNomjFf/t0+GR7oIil26A3e8DIhdw7ceTCOLUxcT1bz1Dy46SEFs/oj
8mySpDqUaikrEf0LC4phctxEN6NaincysaZ2zvEK9Nc1AvH3v/gAj/E7P+/8nzGm
9zptW87NqtoALsXI9kGenZdlz1oI1LudNnGrqo+njqvGRh5hKlmAepr4ZOOZ3OqL
nihl0c4B8jVxiUO3cvyM5NXsQ9ZHCLdvVBpxPovgZj0e8G6VCaFVrUSS7ymlY4q5
L/PvJRHQdfekdSl8yLXgjvt20jkmlo3RTlKdxaRHWlcM4OaTjCSZq18e0OzmzneH
6Y3klB5AF/2Ido185UyvdRY5lMsuuOzQuR7Zg32XG3bzf94Wumo43fZGDSMmAjvA
qUgPrmal60AxeNQX5L1ibvLolS6xSlpwk/5ahrpqzI0Sy+LqQqQnT4yeQIEjwmYg
agdEUP9m0nMNE5kirKlmXlzisU8jOURKV9SFGnvdkrPiv/XjbHqk2pyn1zpGFMAi
g7JyRON3LxMYe8L7X6xAt2uqqKps/Z4Cz/awfyPybzx7lJOG9vJPdDUXGvfM5MLN
4ohoTpjhwhz8JtufHqXCvW077AIDNPeaS+FAHThVBCOcyE3TTqQ1nuRuwxwLdFaO
WnytybCq1sa+Ws9kPBNd53AAH9xu4mJaTmyV50AWAalr0SOmHyvdphg3wmtptPdq
WNaKVZUUs62APGvAkw37yQ2GxFdMC0HM2b4M6yx5rS3p2WvV0uHQKrLHyxCObfpD
zOlfyXsOW9MgiR8vlCDfqsZMltF2nxLbQthj4XLFLSk4+jd948n7I6elk6gmrTa7
y6o/eXAo6reeW1ae6//9sEe7FoXTI6+AauVyLh3JhR1KCr9iSzaG6z5sZgHjrXOv
QmAPYbQS5E9qcnfZb87emCrR2IdU0GQtfqS2oeKt7NVBicJVf5RCkn8BW8tc4zUu
9dR3DJXouPENcjpzuxwqgb6O1GjNugPlgaNS76DmvF/l+jBhQcE+5lVHSmJ2oKIY
DScJkdGxyXegWTtWfXfUbOq+N3axGqhef3U22yXRrHv78Z9lDQd8tOGeZWCHE4P9
nSevsoaHYLIoeDkDWS8Mf1Eg9glEgUuAANwV2VIMglN7ph8fTGPNilERgz7cttMH
E2LpDVV00teosU/xpRBl6pdnccObw/CQnxJt7VukpVVD5O5vsYOzjBtY6oD7za9a
o5uJ0Sl0ydIBefN45yaAyTx4OHzCKdYk63dyZ7UYtYT71/xC9A65jLJqnABUjEVP
Q9WRt/xBZxYqZipFzWY/H9nuD+E528obGLJr+oHqrG6MvOQNxh8HFH/bipMiEpTI
LWE2DkieUtYJPwOGmYTnejBZi6yHywEFmbCNjp3zLCwyJICVGBA8PByCaZi6i6OU
ZACRhrk2ACK2m905cQaCraLmPFPYAY21JPCv+9oB9InsN0/3vP40o8rm3xRusFJR
/ebHrEj5gqtFvI+JOmVwKMzxyMS0Qt5m+wdhHH9dLPrZ9qamWrO7482xjAXsssKb
EyblMk/X6ZdOZEYfkDo5EkPNxWSu7H94YgP+tajmyWM9pPBUEB9670QejwinzMR4
z4XqT2IuBhcClmziow8xzOIlRlmPcwc61eSB92Rm3NSh2NrdccpkVputqyY8YsUM
hCsUSKT+spREhr+FUJ5oh/sCF4aqAuVF9XFdmmxoRuYa7PkbvifnA/zNpIcsqUjV
0bixsNhBAU7lCYDjKTeB380ASSOJoRgIJoVrQQFdX4L/sLSVz/1g5IlVzmjIgJVS
b2gAVIWJklOKZ7neqwlvpUj3ltB8CwgzsOHoA5JIng+Ggmvb9SexIDkhA7f2YjtD
ow2cSHUBZOdu49nBJJABjjBBK655Nzoth3c3w8Qka+YgxUy9w8snHzLVSxK4ZgYb
/kps5V9fH6oKgkf6vn8OZmU7o4cIOr/DB2nA4O0bZ6elxt0KiFZKMjVduSbBjTmY
X8eBu3Ox40dgLbY7W/ttdNfgSK0hitbM69uyMLndtTBB/uuCTZobQ4/oIpa1H2ow
vK2vMzHAmgTrP6I7eoMpP24vdIy+gUsL2fOnocvz2RbwwjBzCWEvkkvwvDloeHLq
t1Rg6CbWsdvW0kd0X5Z1HY0x8L+Z84t43dZedapbipVUwwuwrsocDHwf1BHSa2B4
qIuEhRbx9hQYd/g5c5Z/8WpYk+/GnXeBLkGq9A1vJK5+Gt9HeeD/4bVCwUXQ6fhK
b+WDygiSW/z36FJneLp7T5g626hbcvQsUGnVxd8ZafggdxwL7htt7qUxzd0F5A8J
BwI5pibkncp9mk42KzmiZiiCKdnNN65jgJOGK+UVbjAMrC03D1ryuv3sXYN36E0U
9JwwlxINvGCEsDleajE3j7RFJw1aDRJxTPiildxCdwKh8V2EnxNqtzYHPgDvndyc
J2kJzjYqlKGWKiOQu3rw5QruyaM0sA2BdfI73Y5viKLHBI12ezGC/Qj65oirz8zx
jQU6ZSuaaHKpSggqS4KdLUy7/aaGZboUZPAeuOPsoQbpu6CFeEWZCLGHdSCF2rdx
WvdAAgm+YGPDwOBT2B7QvZiYTzCbIrwlZfMEX4cpLpvfQxLjPwLknc37MPTTgJAy
u89+ACau7w0zfiSRzBw4h9xEBUwX0T3SuIQBZFfGOASu7t/tc8AvI+O56reZWkIO
qHRCz7EsFnyexCFza4VNd03zLi8J56wPGgf8+7i/5njbppSBCqxgKhHOuJcg9zaN
mUYmFd5T/Tu4lnk2jSM9WMCM7sOKwFD78XSDwz+jJS9H7fucknPQ67y6miRAVZ+J
dVEqfUxNqF089CA56G3vfCKU59ZhqUdZhm7xMECS1B+yS2RXBhc7j5/VcSF94nND
VsQMbMd5id9xVmeKFwCZ4Y3geu92AtZ/r40AuvGMQPXYb2hQhaukIq+8oCNwHlEd
LUF51oQnzkeG8WSNhOeDprldAZm2zkDjz2wzaiW+iq7mnepG2D5B2YwjNnmYkeIo
PilgnpUwwCYJHUsTfo4MEmiE0UtmyqCh6MjWKdwQdI3yWmjMcOnmS387/UAiJAAm
SD81YgzMItei1iwDaWcqZ5H3A1cvcCD47BKccvGC1HILGUiRqKUmOpnAT+frGCXt
QA/HOdQTwgYAmD0CUCKfSboyFlGT+KY5BPA14ZIez0j1GURxoLk3/LpnP4qq8EcT
1dxM6nfixtB8raB+YGTpdWFEYW+NawZrm5iBclzMjhXIjRAi7fYXbgt2ZiYw0l24
MdzZAz/bOU4HHJLz/dcU4JEYZjsBIPBjbXe36/qi2pW3KoI1q9edQLAQrgRv/L5h
Rq2DPeNAqoYmVPTJ8pplxrSeuPHy/GiRVUhI0GV8xeEFUmxQHWz3FVFh2QFdDaOL
EhYlJkc4MkkLFjHsaCRbULjckW2TvxqJNEBWktonX0CzmSERyWg+AuVj85vlvVep
iYFdsNAy+6nbncUD6nPEH3FnNtZCNyfyl8pmiZYihR4jmMrWEmeAkR/uqBbPncIQ
HjkOWJ6yKm8ls3TYWjoegvbu4mC6jSEvjNaRPJ/dkZyI9cvw9QlAe6dK2EXAONJf
l7uMXhMTR9JY3PRqc3UK9K8902cmVpCIoYeDyntsGD8kH6NdTyahgipCQufftFfs
PR43LpNZWrNTVpOFOudgTOcgP3hKo0dJgAyoNl+O1kMSswGfvISQols5vNUBgp9S
Zo7hiZCOMauqeG8IeBvmG4cQBAkfgf+HaHGeHvbIl71hfQKvLpNlGu37PiD5w+1h
2e+cobpH7//dT4TPxzwgdPVgR51uvGcvA5RP8HNOk7dxPsmKAoPBYvXdMKTXeHzL
oYFfarUaCd8v6Y97lAF6nSQ4VTeVAp99WL5w7QenFpK7ywEkG1M0TA8+kFF5RPwj
L35L0aCFfboYJE+2eJEssPDy4adfzKP4ZzjpfPbSeYAaJ9hhoFZFvmc9RwyLWIdv
373TsNPtTZCq6WoIw7XKgooR8/sTwrnc8rojj/MdAD/Idt70+h2pIqM005lb7lO2
15lejs2K8lK5iUfl/H5OZhua6CwLLm1U1EtjMLq1QpIfiUCYeIWI5gur0zZRYpak
oCeRIo01xov1EFoVl3OqxZpZ3IWhiW3UNY2MycqpopQQduQHnXLXpREw2WrMJR3f
wpzvzgaqVyyWC4o6jqbEhvUIpWAb6BBaTfEXrPuet94yLcyGKWwavvnLIUzPvv9A
17oOYjM2K6Xcq/UHAluBruk0lJclu5vWWit21oEVxLs+f3d8tqkOFtrFPHT0dYlc
x2IXP7+udaw1c/joGcuSVP4XPImdgEJKtsNiKvWYfjBimt8bYiqFr/EgR3G82Hf7
o2JRTtzelJw47UAz4iOI35Ck7HLksKyItiF5t4xamOQBi9Jth7aA9t77yzC92x2k
gE/wCGIL8xsRwHMC6a4tO9A8X09y1iP+73ONQlSQ9lhd+ng3ctSZM3H1MwQJhZkv
h3zHw6NUPoQLChDGEqkz8DK9lD1RDzKB3xDKIBYxqaHUyYe9v8wsXzoc2tEfgHzP
11ASAGPfF2n/7AbbZvE/yodMd5j9C9L8v3DRgEtgpUeZu9W4PY5Fa0pDPDdTMVrN
U2p5pA8q17RccppArdsCCyO9zeSeQmXhG9MdUCpbfwhn6HAzEZB6AkA/o9GBnaun
nOEjzMEu4Zal+Up2vV4D4j7dZtAvMor+HHP9/TllZ1ULvxrAB0HTf1/hYAIayUV7
REjI5rSP45DBdEWQEOrj5c5zIdysJLueqhAaG1D6M/GL/3oIQf30qmD0b71MQ70e
GOtPm5GXfaQkHVv8wjNDYptdAKIIVRcOAJqrseSrgj4gkVS4WIm2GCb9UQb4m6P4
+U2EpOftB0IjiG07Bs4W8tDWKEEYaB3pabOBVD3egD+EFAtOGFTfu7E+l0cEHI+y
M8NbnbvHSdErjVw/yZeYZeKH2mIo/Ph1OUuVzyzq54NDTfgR8YMh/4adpN1s3aZN
Dexo8BekdstLx84SMcgMlLmBrHwZU1qcUND3eo3ouRyRM7ST44plNbB6mS6hKVFZ
ay/xUOHA6COENEqK8IpJRjZLru4HGcA9b1OUMBQkainoSEIKFNgjKo4pFOHoRN3n
RDipfGwapJUORko8TVIz3iCviOAIPadz3MgyeK9GKCNP+rIMo8ArmdhflmbxSyuo
8AH834r3Q4mELg2ZBGeJeRfVInB3HQIy9M9sStZ+vdiWTDa5CR/EeiIj7+AgG6n3
HRn0J0XkigAIw8wU+hCmYV/R7BG9DxEey8Xpn6PlBsk6urxe/2GKdgTLJJ8NQJ+t
Um4M/mwKaWgki2z1NdIUYqEC7bYQqf9RH3gZlge6RZhPjkdNbX7oppk5I37GAil0
E+sW6vMYXV/fJ/gtsQ3k6ZtK2QnFPI8YendBXjrClDv0mc0IO+pO+SjdoBc9Ucwk
n8GFtowMk4ABopPJ3iQog9Rzq1KzyhGYSvV/uX9oClT7yyUTdhaVhscJHPMdI4JQ
bj001Xu63DGzhIU+g7dawPfE8ifiaAG0tnbS4X1ihTHALtbYguy52v6yh410flUA
psfHdrY+ZQOYpPVEdjEkUYqbxycJFp8fdBXV6o9nl2qRuup/roZax9pugFfoiSwh
I5pw1oeC+k9Ol+LmZhuOWDPe3hWvOh2TrdB7JWSaLmKoP75B0sQS6JAG3s8WnvOC
qjsxteq+LOhq+tH/HNvki5Ufce/qhS1qhbYmx3wIqST13kLhH0Jz835/NKp8xWar
dHIhU/xDwOGHR7qRArqmxSZHz3jSM9dulrNrk3EgV70PqEdNsTA2pkLkmD6imyRt
LkRcMssDofe/EOYg3q+FBh4rzw0abibxpanGEv62+yb67ZL4zZ+6cdjaKuIvnbuA
uSioIJwDI7Qr96Pslu4RFzs1ix2Kka6mZ1l4g/GgmB+ypc6Yd45mwcNvaSc3zRDl
RFQqbfjF2FCOL2t6QDuxbrK4hc/nJ0ROwRrrQ6PHaedkvoOHdwF+1OzPIR8lPAic
BSRzifvcOlAHWJ9R80F/grHcysiV2wefQgmWn83Jy/MJ/SPANJD3lZgz92KcZD/d
wMTckWuw54v0k5CGm5fXgicsTXvIoweOobVcsfou8pX7wz//ioGqAZ/mUH7peB0E
ARcpyGZ3vJ3VqEnnFS9ykq/r0apJDgpPq9xMYF1QkuI44be6Edgs1dFI9iniiGNk
eRFFQYIbrs9a42bu3P4qpAzHw83ZBsIAvqJm/eus/VFkJcSxMbeNDMGaEMxzSDLY
809gZNUf9n1TTBQ8GJ1Go7j69r1f8ZRsA/dz69M6TU54m5G0Ts8iR3nodHGtukfO
N9gSUmUF1YT69wHnkVRbsRTMOQIeZkuXGIveFkcb/ALig+jQ8Bb6K+i2IXtk4mw7
kNpkrqBWKp0z8SdcCAKdsowv0hCuNchg1R9UB/ynOpffIT4+8RJCApwzbB2Eqhdl
zpg8IrY2H098S9Y4+mQAXpya2n54iQwWMW5PN5SoZxbfJf2i0tZuA70YDUE46Up1
nnF8z4H7whFYieqZAbhy8IfQUaCJG7v32jis9D84aqJqTaNc3FRWiOinf5AUGbuU
rGQlzYlNO4sXEZ8DiRp/ZM9wEyJe/a89iOXU8/mJyvkFRbVxlQ1Enj1cyaaZ1e+I
0YuYX/vPzhZ/owK7aiVxWBKFkGrVWcf1ZdHJxnKS/c9f5TMXZdOOYS9y0UH3Qmf5
YXxeDu+XI4x4Fp0HfbPkZvBe+xICp7n4fb+ZVM3vykyoO1Xqqpew7L22oWLiZ8m3
9Prm/MXcp7v3Z62oRo5Z8bkzPvCKAEkxIzD1piXnzoq2AaIXlJp4De+p0c62zg83
VD6y6BJV3tvNIC4Y7cJdbsS8sGtoOG1SS4aDL8XW8ee91NH1MukNAn7q2CR6jJ6Z
SQmTQRmZcGpdOe4D6CFuCi59NP1ZIwGY90UN6pZ9Q7BIqnG3qDky+Ye+HaESfSo0
JnYUIkYXOWuEw9JKbpDgQpH7otT5aQ3VdiwS+soYEiLl9N9+TBmF2P0V47CKL57P
DgOtAMc9Je8jdHu5fP4nE5gZRVS4RLb8LMixZ5hNoNhv3VjMuW2ipSz2Qyj6P7Gg
UXvRrfh32vM1gJDTMSgCEksNGqHjc5puOHDQkLSYVEf0rqBzjno7Gmxm/8p8HUx0
mShnJmJL3tlri+dhmEd14ObhTYcn5u+zVVRCCvYzuoKfYN43SCGE+N6p9U7zZ6t3
9aeo+PY0mu8JzYxLkWMRlfS4z1gRPu5IdjLSLNw/zcOSaF42SABpk7WnkPgBNhNI
SHgZ1FgpSd9CjdH3aSyUeFcsr/WfeVQojTjNrfNdRJRggtcUQIfOUqHtnWfkC+67
Vlf0LH83EbuakO0BLJJmyt6yDD1HdPeYY77fWW8Mo2JQJyoCV3zwWLizf5N/7xUN
/uRGETyesc0NaVH7n5tiKl6lCfIW91vMURCS5jJWUNLGGWauBp2BC4RI7LjqpSJJ
Y64fA8ANCJyT4e2bR4FAx5vLa0P/jTKmzwByeqmXEdWY8RmThCD0XKtUaQNxw39B
6lK3+Op4J3XnNnu3ZZ1pq4HZbxFuiMb4S1/kLowexVnYwEffB0xPJcNYlgvWq45m
1ZguPm5lhk7CZkWmMMD1YxUEClW5xqij+0SVrAeaeUXcDlq/1+DLbdHg5nc3dYZJ
9e1d1J8QDBZRS9HLF8bY6alskup6QiwnZ2EG6DDF+wlt6ql5gvt/SRjhhVpZFfxO
DXlhR+nUSau5Df4f+aZHobAFu02TlcBLqAhnistJb0C5TYgaltK1Kt5M56x8JdW4
ECCJRfRHSXfOLZ+qP1ElU4DYSiMdCYtwBkL5vXOEOoBVtkRU1yOxk42XcqMNEopd
0Ctof4xb9KSYEGWnn3u+/w2dzI6nFIXYYtKKzgH5qdP7Z55pSlseyCNyTrO8FHuo
wUgL1VdpaJ+P/hmd91W/9GnfAo4YWYL7unxgihBPErc7fLes+A0fpB7txd+Gd/ev
KFYRpC2L/gJF1XR1DoN4SncB6pC2fHydaDQGkGGmBHy4kjPVYYuDRruBkgU5jRFs
55p9LhOmtWfXXr0r1eCShretM61xCFek3zrLv+b1FZtlN3/zt13KKxeSUoVyKTlK
z3Y8f+EWksQ3+eQWUpdt70BY2sYqVvNDnBDUfsfxZnbGbRQf+xqkeG6ROV2SE7Yd
t4Vyaer2gR2u69aImn6Qt3AbxZSdJS2fCbmQAaBGo7yzTbOZ9EGTBh7mPD3YIlNA
5zw5JdX+buSC8jNc1APL1Yj67XA0SqU04kuxJIkL45Te2IpLee6LPwYZQUXhen+K
/f0dND3oOY4DvqrrEPQTP8hvn+3Rs2x+aq7SfAnunCR0usNU86EihGERfhqVRFm7
LuhHDtjNrtjVosbWk3CeNLSyuK7kneuNMSkQdgkHUKZhNn7USmzGG5f9tk+3a1kD
DbJAYehzN72ewk30Zg+kWg7hk4M0ttmk1fW6kZw0bSx8RquIaC2EOZsF8K+lCf4B
7EIg7IPA2a2zk/sHEcL/fGe8fa4DBC2KGFkhITlt4+HZhbiSS+svNoID3kegYAd1
w0E4zcyPETU+wCj30M4vkPfa9TZgg1dblPBxV5+XmVdrENnAAWrWKbmGdQKpSVWT
fY9mEES0YaUCM4kk6asVAYv1dro9KkAtY+AlbQFymQrSKNsoXh+PYJ2i13khc1kG
glrh/25w7308oqomcSO/2nDC8qM/JHYMhfya+ynypR+oW3QnWAbkO3N7bh9nm3li
0EyF9w1oVp4eZvHM26xA9M6FaC+CGylfyVstWA90aKDf9Ff47teG03vLrj59JA5E
fn7KWJtbVVknAojuCSsuUU8UYVQfqVkFdcO9U/YDbC56KSv/3Amm5UyzWpgfGpVX
V1jUa12u/vb+jyESsua8gCnY+MEitFRdP7cGYjq8xdmR2XNDxxVsWu9e395FcKj/
3O4MfdQndqZ8BguwhjnlJNHwd40o7VhGyq6YCFxzV4Xkw75T1R+MpA0by8floVqH
USo95NUNE3Y+X/LP8+bKaEAf87xIJsqnEbdYfWMlYpmaBcZlmzpMzPkDHj2CxqAz
/NnjVFXy809keAjdFUKc2YWUk9Ffb0va8N/VIxv+0Ci4lPnEgejG6w/P0MyyVN8N
BfLPI47MIot6zS+/q4xYcbFfEFqEu5mkzoH8rXmHorU8h7I+T/hCNiQPBtlIdHWQ
iHsTD/yh2N56pCXa+P2oU7+tfhtVyDYlEy1EW2aUyFUj5bA3LThABDVn/9fDNf/Q
RdGhZBZ0YxAChi23AJvlarU9oQn1Pttce6ojCObErQkFlixJ57KFy3VUEYbKj73t
tKfIQ9nrb4/q4lplPe2Px9OH6hnYKwQ5ltgYNKRZ0/UAOL/7lICUG/U5oaRrcduF
BfKaJn8JBdTktZCqu8Mqy5oUdC8qmTRkuBnJJFK48JVK6IXfdpOFU/F7ApSx58Qy
RyUN8WXpEvdwsThBaD5t/UpZk3TH4rsaBxAypvm4PJGGQWl1NuC0NPOWuapY+vc1
CNGNtqoJqxvJAx30204wtNYhBPhhMN+hZeXT2ivGHFYTkoOSqJqeQW1Dx4CJzHtR
Xr+YdQt9EjSwFTwwEitmxUrePXUd99RNmbTKu7s+Ezkm/I4Giy+MPR0XZVjUTxRF
pg9zMx37Eein216hS3xLR44ZlIySaPeQMhr2u7HTLUpQS4ycbhaylvXJDlqEQSYq
f7l7IaIHfu4hQ9JY+XA2jJjNtenlTlIODZoW5bkWun2k+ckSG+qOZf9U1xVuBrmr
vHYRumgIG9oOOZV719eeh9ue8Ew66rr9/RNud4Sn9Hwkbgmprhw5pZlWzFl09vgZ
JAh62RpxwcE3+Ul1WHDRqh4UBSGPfRFSMi5KIOZYJCtuXDSsoVeiQqi2TXSJc5Fz
cIXRLNrWPZs5SB9Kpm6qnR3zcg5BajJh42GA4vOZneNdP2+W6lS70dJAfLFSa/9/
X2U6POU03OENB1FdJcdxmUYPEzkC0pcETtvhsHTNmQEOCDgO2GTtGsn3zVi8KsWw
pBu0N63UQILCfIhhZxO79YxLfUynMuRM2SwowSq5Zm7giCWgjImLeL82ok3tI5at
bvj5pCRdRVLr0p17g8ISnjq8BfS9Jl3Icc4JB22N5NkUDjWiLLFQuyvZ1hdSpF+Z
FmukfxgrFWUna600JR12sOH6C3iXOYAyr0IDX0WpUfLQY6BuSQ7hABYCDr4X/F5X
OOWKBQMiX3LO861VnofHgcwrXntSbGovsNjW4/0J1X/ppFFMaiXxmiy+7jmrEQNs
CaPOllMwL1B06L44czyAdA+c0x+ayeJ0qxWvrCtSSnEC9W/oeiLO29ezoa9um9nf
Z2G7t4YwZeeOYjb+PTLTqCOlQJv0aDHNvEXBaBONkFW8mgD4MDWG4x86gkYvIJcr
HfJvrXRnzUys0nsIzdK50zAKrE+iYCwY+1s/O07dW2dvqFyqJR3V2Og8HkGarT3v
ISgZl++JM3DqjvMqcTLjNGr0Dz8jpbn/7i6KaV2Yd4idUvNVMqt272IVGpkF6UtG
YeMaWWWBJKAHV8zqf4nxvpwg1NQPyw1b4Zmo2cBjZ5e9/HWqBPdxPS5mBJ0ht7kg
bpLxwn+bj08bR5P6enSW7h/PKvqhdGbKCxphsAYcGokVuwz1ZwMcGMA1caaI1fcR
1qlWMG7zFNetqbIoZxL+L7lOMN0nisLVIRILfuIMmdzYxq9bpFqkkBpdLupHIyVC
vLUoATNxLsXc4MTGHZqdmv3RNUQb37M/8uLpjdSbon0aA/o5Hjz0IKTcJJe2Ym7o
OB83+k5wi09bgFp4+33W7JbHGIu8kdu/EQSZqrgkeIv+phrLXwbfMiiHGMkLcMSx
it0U6r10mymWLSdHTgXQjFaMd4UmV8W/IFX4POBypjUlvlsR9WkTYSAMkgFRgcJO
KSsngMbqywmVUpNQBmJQKa8wvqEXa/iFn9H1lJfYTr8bqz3EwMHzqH+9/jwsjWtm
WEuHv0x5O2R4Y/+DUSl/Wnoe/ipGm2iop0AdcK+j3jgTPx1cQrqc4KrOBNcPXryn
C/ucVQVDV82joE0XohetDACdehj29E717l4xUeBwf4dkBvbmXzfz/Rve0ezthP5i
FfdzQ+6SR5IQZ6iKX+7OPe0o03mwlmw2H6GpVCluEfa/kNC622t1Tsiq4Iilo1SI
pewzVLZxmQFq1qxwXxwn6JKKA2xiqQU75zmSXFp07XXVBpRD7/+r33xg0MNY+tkg
HkfPe9sYFaan/MdxSe5pDTL3e+MhKNB7xOv/h/rPeQrzrJOi5/a5mwB9Lr0WZSiP
SemfFf0XvvBaE9kSDV0qRt9FuTLvcAC6juc9N19DLhAlLyZU1ua/r1H4reo0Nmh/
bdse8Zfev3mV9zDkceJqbKVuEa/Xz89EqT6Qx+HGy0mhpqyMZtuSTWXXFP2uvpcd
4S1l9rCa0bePoqTO4ltZPsEEnBF4HWKdm+URHksvqA5YcOTr/GukQTaoXRMopg5U
XqzihSKVGsVi0ZYi0ZOt9twEjxB2LW2IUVg7ddnttM2u5d8oBmTitpJolrfoj9hm
ut9pXpYfqZ5CJs0XvoBOQxCQze6NWWxUi1XSykwVF5qMwyvhalJqBite756vDwVV
1EXPl3kFKUwamAjBiDpsI0Nzk7eMXsV+QkPwafoq5AzULX5Khi+FFgEJDydg49w2
zJtMKQC5LPs4JYkEBowNfixy419ZPIr2WmE2+kgR3usadVjM2TWlkvXn7O+DHa5q
kJHVN/fd6ONEl+ZYPc1ET5xflPx0L/IalkQuD0P84GBwoyVEnkzXOvJ9RU/ypGja
Od/851Edfs5XBllpU/6MXtaSKxH/SW3v5J7YG4jRmK+8ZFSD8sN+zp5DhM716pRz
63p/KgNe/Kjpkhek+7i1jhCG+i/LC7fiFd1rYp47z3hebcy5JxiORGAOw3068q53
nWUj9g7qNEI8vqWK3X2K+OjFO1VuXnORLgqxLaxykBbX6AyIbP2ZHOnSvGAQl4Bz
pWzsAejycoFquzgWL/h1l4O/DpzEDA/91qU4gaRMmu9a9naax9VSjY/8KKszhdcB
ntzWStNhU7KKgqHfRDXALq7TRjANOMG0cDe2G/OS+exWtsMr0HJ0VsgJTv1YI9eE
fL+OGX4GORtFdRqN4kAcQIokHPYwZArojqcMne6eWvkEIqf+03yQZCoSrJOLavaI
q+L5gi31BXOfe74EpOG2jcECXdUdBDD1ekeGuO8GW4lmaxBpUdWTKsaL6n+7DZGm
cgWARMq24XkVbNnyzHOjFVH7HCTBXYhMafTDqSSpqPSMZjAE6e2Z4tGG7Cc70QPY
3Meqi9bP52lODO0z6eXARsfqm+6jGd3uzJm7gKFLzlDGgJlooqaIoJgOfMqAICc3
V5Fr9BYoS8WCxqjeGwFaQj52+SGBJS2i+ZBUeQMGOhsLzAGdb+L6JI0jupjXcqIp
z2iUNcJ/3Bg4FxeGJJmxBb0y7ewzuWzlZ1DPfPv2fkPMvp0Go9KqUzbK513FMJYU
Fq6eb8UlkGVdbcpKCvEx/hF3S1kOKMvHRjt73oUPzFiQLEqzQszepWxXmyrYZk1R
AL0negiILJOvlUzeUsvRdfSXzn1zcnPZ2cGa0iGsEfFD2pYvm7HyoNpNWXQVdAbp
ybi3xoFDe9Zox7EKM3sgp8WOomKNvRArLhGcCJ9WfUyxqJXKWDC9a1YSFoddHsI4
1m9ylaW1D72OGRuZtKADj5N4laUNYYiz0K8hRjfy55WlSRPoG/q5OYYTXq3XOW2n
7RHgue1xHUx/Qxd2HjWPbMJI0IWnRGl29GuHCfyrmyPxq5Xz2Jhi9d1QKVf/DI7X
2kc3xhALWkYIzMJt3S7Iur1LCr9zLCrNQZwc+2llC4TRp2vJMij3a+Iw+6IuPNr8
eToPLiesWF4gyZMAEhfox/y6y6r9X0fd4RxqqLZbDSWZOzW+knsKZymsBECf6a7Y
4PBxTTqkMlW+Y7ur9aRodE9aTbkVTHDC60FVnZZTwj4+Ye4uQ32ah0kyaZnoG5qw
zmjJ41ePLMd0teRJmWgLDlBUTRTey+na+UaE8sxmw2KA5a189NcUnExzVom77Ug8
PJxrFQar/rpydfAnIBrqWLh7/9GmKv8eUMi7f6lIdnu496iWm7bnkaSYwdC/XB7w
YaQa5zr/63nlcdAIRB0RKhSgyAP3M79lxqUrRctWoNYkqRvHfdRBzECnatjCj9VE
eys7pH8IkOSwwDrscDfc8DDtojIQVusj8gGEiqpFqw94bcSXRLVVK718XI7Gl+gs
o2eU1Mv3pkp8DWDo7jDGipAnnWHpkiGTPfvVH0NMAaJeGAI//w6Ig66CgduZACto
NVPdcsWD3BfrkoxT8lr7bBWv/ELwf+G3jsrTO6D6KICIO/m+eqEClQIqQ45T3Ulb
Zokbl0XnfafZVVMaMPPZMwBlRUvU7Jjhdq/dnfFFXKXdz5DQd1HtNKMcKlDpg3eM
F++2T7sT0IjsggHHF+JM42kwlxUENRdhI0SJkqe1bdrukB+mFE9ffMLy618dE608
Ig3i+unTp5wn1e0RSqmL7TojD168E9lWHKCOau2p6yhKS4AWMj1+QQEVLpJ9RJAu
nBubaZ8XW5URgPSXnXthY4+9I13UCLy8wJydbif2boKsJ8Z2YbYW8x8dSdhOR8F4
PFT3vAq9Ie68ShWvXBVqUTXDE0/hdAYkubkDQ1Rc/zAlZhu4NUz+IVzw8QvOEWQ/
tg7Q7cSI4NWGGmA1O6BG6yQLzcRIPvCKs5Q4oXvZfr/oJzUcNO+YEqj7XIy7WvlQ
Urj6X16jLWvRCWmxYRzjuSf8QYW23zefJqs7Cmt7sJzTh9Tkfu+Fer7td2hVSlJy
2xnwJTi+ju82SVmIevQMtYI0eKYTKqBZt+BfrDNcuKdjOh3VKEvLEd732aHXjpSk
VD2Q8t8iMn99BJMUW39BMN2QjUJb4GT55qaouTlkpcfNxyVmyDDEFfGiwJFYpdYC
nUewUK4TxPRbI6mjBbVAveXXBMW6PQfXtHcOv28HDs7sWp9YVfTTmdZUO6JG0QkH
S9j5+dWjmSqrhSNzeMl17iDPGKMTL8DXbyKx4SygCYXazJANAmAgwc+3AImfalmw
wvES49pgqeuF3RxPf/OBKrzK0KGzITXp6u56j/YL7+Vcqiy11sBjzEkQmAHSGdqZ
fwPfNpEvuEUMxakxtUjjDKKeaDoukd/ZqyC6rcFEX5LVSMR+nTNln6Fqm/b4HlRO
k/xnPF5o6SWisoo4L+ggpj+fTRbNiM0vIsFEFGsy0Bfd0lgEXoxJ8uoJ5L5lMeXb
zZodR/yOGgdTzintXb+tsPblpEg1BksHx5LNXZMhHFfMBlmfPRIJtjNUYtrn6Mqx
KBp2iOD+uCFD2O9Wo19OQk1aXG8KBcTNWKYyGpxyDxZkfEVfEIZs5TMb6kDhh4Go
0zBbX+dPbEUh4G9SrbFHf+lFMWUA5AFhwddv972NyuKrB8jNrVOgddpl2HczggDb
nUlOeSoqmFIsmzz95C9F3huAVAH4ABEU93K1bwMaq70JnzMSiTfw1GaYlQFMT0wh
N4zTjVEQZ9S22TMmf8Ca5upWbzvWVF92RMrPHrFEW7UORUUynMTjt9uqa77oP+6q
RDGfZS+1i3o8uLdYayviaOnyksjRwzCMq1bFM3lS0tkUn0EkaerIv07sc8sLuP0v
8IEoPVrzkKSKr0cACV0XZR6aVwYZNCiWuHB+dfYDdskABQyOpt46J5qmAFWtXVNR
6WbjrjnIkqQXm01l5eOUUwKTMsbIIL6KWAy+xpujj5EwbUieNR83H6MjdQhP30zP
5GdbXHMW6AUpo+alkMVnw15zSP+SiuuxpkccV7BxWs9PteOg9dyQHEvyDOflWf0E
wmyb0a2mt3ILrfqb7u3L27QyzDpxORRjzCNEVKGipweYaskjUQS40UZ96OHIlgxJ
cQrgVV1uLrbLmYTuMek6FD+VL2nzHemTzVG9hV5NK6Ej7gUPnDgwjGriq7ftFKEU
NEyD20xzAcbZ9GyImYDhggGVJCz/tKxfvfwMrXJdLkNnrn2OiPa2l1oIKuU0QJPe
wa6TAIYxQrjiogvAOyM89Wbih1oKZMxyHQOQrWuEEc3K6tRfutBv6231vuS3GEs7
NSQvuf8h2QxpSDsT/KH2knTRcTTrkxzciTeG4tTqJs2wBZVXSo2Qe8eZR0DxjJ5k
3WJzNERmaP4OqhESelYSQXKZoa6wh96ZjzqUwaYxu6/xx4TevUUUNCzb/HTJ7zMI
rWXsLczza7Af7XOB9+HJWUEPmGOklqYthDCkPqDt+MYZyvqliXK6tl35CAvPD/jE
JDJXZ4A32HqLH2RF0JUaaYqX+kSlLrn7oHMsczILCp1j2wUdVuKuD7hnDrzjU8Lj
3c8s7k0Axt0AQuasu9KbtgBJMShXRqUeVQeE0tzC0UQcKNWrEt9h8XzP+nNOxm6Z
t0+cJAe7LKN8u/EvjEz/+1piGW1/379B6tWCJpxDFHEYjl8a+e+vH/+kq+cKUPsi
7sJMgyhMgBCA8UY2Al6RWMf5pWwk2+NG9ycV38uwkMSUVUBq8Wzo66/FhXjLGVMB
Y1ZT96joeT8Kk2SibRxpPlq9tiO/cszshT1JWJPvXspXFFmdx9D4dd0yDeBZd5Yx
kytJNfXXcVjuisnFbXuKu+fcqKy9HfKOAOiLEaKoRNq8T5RW7W4l0fs4lxBhWiGL
fD7jWvHDtTjYp5Gmi7nMgNhtEc09CmBW6ZJrRMpGlHIr+sHzqoR7Bl+1q9ilW5Ay
mDy/qclWIZqBx39orh7Nb3sTdXjaqaorknM0YBB8oTdAToDnYjEtFTW7mP2atVV0
16kk9lfPIsgA3CQJhxFLnuDF7UaOSkYiTDsbqmG4GespFF6CYRFqjcf5r7U6+G8M
xasxDN6t1C7vznklY+SOeeJRV6F1xvYO4gTBct6x5o2eDKzUf3xomH6sGPpYqCt2
OfrOFZjt1zMdq05HERdUKbVY2Ovmq+WNAooCvY6jD9u2b1R2K3gNMFiil8nKIXbc
YrW581NknlyX7hAXt7Cisu7ZTKgGARJoVAWdYVSxoCAjObR01gEfMc/G0Rf78lYI
KN9RbRhpBoL6U97bzVZiy7t0+85I4Owl25UtTuxarZQ+rUBFRgobo8LWc4f+e83S
YBJrioNgopl46Mcpixby6682loN/Lf1OH2280Ao5NM/dhMpXHvAka2l1f1tnPcok
1qxW6ji0Rpy34691Wudg6uxkRrSasQwa+qjADJ0fBKP4zXUF1pKppf9D13WTObiR
Sp02iVW28YvrSkzSASQd3K5edjba92BWVDEdqUBw9qQNDFMliqvYY7WOQfjRGfwi
VKQX7rDVoThXmHl3MqT6Qq8h05GrSSNXtwrPtumnHsCgqDleTTIwa9ZonlJ2HxfJ
gF54HkJ3/C65JFC65A5JZqbwZz/5YT1+IGdwOOYt8xMO1ltyCPDLt834NXrLdI3d
UVoXwW65lBxREp/JQFkfIcZQUErfS0qn9bS9t8Gx+QcuSM/fyC6d4ZSlsRpjwsAY
jL1tFjsyC3eWwIMkFtHlG9AYu5/8VNC3g46a1CvkKPvGo9GbSelwQFhzynoUzLPJ
Sbtf5afVDGvnW1n2HcxryfiFN12UgYAb4zGdmZ4hLRJ9ZD3ztu4o/oevBSkbeaUP
wb2RToY8Fn5wOHUEqY/ZXVLIFcvu+m1ZN+CXED+c1wvQTQGL9cN0ZK5odUpA5g0a
w8DSFOJH411qa3RYzeDEc3ZIppc3aKHizzI+ifYhAoUi9fgaDy6mYS8OtMh6qKUJ
KNzl/KvGqNKoV1TyFLRe7/rfrzJ0OY0jcztzB3keVZvClTpwXHQ2xknXTJxx/bwK
w3vhCg/79MtHy5o03cO3MqeZoDmfG4qRZ8fgYlkNks8mBuA6V9p1GSB6B8EUf4PD
/Vzi6sWfbuZYPCQDuMihJE8QMxiKzOevmWUQ88MxPDXR3DprmqP3LOZEEsz59hTo
q8T2qsRk7vKpUaqKgysjLtCwpLIRxFP9/DpRVp+qkwagB0a5lS91Vyy4K9nyaqTU
rCtguevopfICUq9LYeiscW2uAu9d3XpXRRIj4wLmoexwYLD8XvseTwirro9jER4P
mV3D6c6N/qESbJr6RdGeibxlR+0gDOJV/UP8/vAosg0IImNQ+qDZNBvwkBeZaOyj
AZaGYl+uF+KfhzVcw7zFFzg66JxjIEP2/EnIji7zQnc8GACEgvUhHHZCcGHht2Jr
/cPNZCa+HWp9CSktENR5JkbF/tOw4ufEL1kwb29hIH05bgM4TEbOlnY/nzEM+Mxv
N93pojGhTmqHO/iYj08FtTMg2Cg+FR166fPiMrv1E9n7eMev7vhmBaRs8ynfSiPq
yrZTHevoetGNoGK/Of7p+rMdiRlr1k/lOwkGMUxPADr6McZRUIU7VS6SUauGmoJe
VoqFVb6Lzxpxz7OSDMnZjXozOm0NEak0UuBt14EJdodlDQSMUo9PYg/OQtsfp/Dz
W22oFvCGFo4g2s0GAa5yAml8qXspiIu4+7XpBswD7SpTVQ5Y94x5FRIndYpctAjQ
J93V0GaJbrqGVz2ISTFofec+HTbWFZk8bpvgfH6ZobmAcTQ2xrvf65lQC7kkY0Ky
/7lRYuNpT4IULQUYL47qSsNSjW8bT6WuTZvmZKHWk0hCqmXijNDy3slQXgNXrVjj
d6dT2lnMw7dZahxDoo7IMH8mjAb4u3QxfLcxyHO97+3sPbvgdH97VjnMWmjUAsDD
Hyba6ljJykDLN/lutvenQWl9QuEe4FzylrQKtk776XRbK2fZYGj5Ae1jBnAeI0an
rDzMp2D4aqcaX1VpQbnUv19NXWkEXfEZnblazTKz3gW1So7jNFGy6jXCzqfmskJU
0ZpZdRj7Ys9PnCbq11CYEC1Es5BVIG12W6sLNJ7kWP5bMqGKOm10PZCYslHW8t8/
Eg/BvtzIo0NL7muvjgSM5IEbh1DvnyKwWrKK0pSRu78hpbkOmskW9MP2phydqLLy
RyDIlvTVtkdrmI94J8GPcL7DK1riK+PXRBchbNyBEbNUgqkzkQXsKthEJsfFsKaY
w0XcPtZ3sqeoaI/PgFmSWZBfNOyFPdaV5BxK4H3mwqA7GRRuAgGFW7sPjIxTm+mo
fQ1yftAgnchUaDAKiVW9sR+2p0EczqWMvzWdHq+G3wvbEkZF+XcoJEWwA6a1SHJP
L44kKDSEQH6JbpvpC6IX8L5tRb3T5XeAmgfnJrUw6ZLM+hX7Ch7A1CL4OiDV3lvW
wWx9I750CLNB6iyfAhCpdTzDdwmcqnqn05SeTpCSHuTEHl603+F9C+lDitF7rsWZ
8USfhmeCXhDjOd26Ni4GYdC0SWmKngSK6f+W6yoJVzv8oh9LZ9hXD1yBgQA6UX5W
RL6OLJXS8St03sm68JkwUi5gmdGSli3MFMx0ymlPtKrjJAxR7F9wXczdLHhNCBTB
Iulp1YMLh5Xbx27xX/ZHnHJAzaFulRQb0hdNhp+eqas4GCm2JZstWQx7mYmExP7D
xg4+73b8mG6FobrOZquFyVmyI65aJXTWnIv0Mzs5l1tzV5VCEvMth4DQbN1siq2M
vtecgGj+xQ17IQffqliZIOuZZw1VzeSart5AHhZ2FVJ/eQujkrsN//gzK/mSdAHn
//fn0k/TKtNkclWwgTaEJApuIlNxcNmjxzh/qDj8Ye0TqlFV4ucU7pmwqaLaRhfc
3Sin3729DxKk+NjtPLMwBJ9ra9vh/BMo/3A02y5t1tIFD+13mpP0GM4DVEgVmnlW
1lYkq+d6RiRBl+1KYqmrtWlGuZgxEQylZ1nijn5EBSJWnXiT4cK06IU9Z/ZrmUaJ
EeSvouQetlUGIi8RpZZdG4I9/Ja/SDqXemdp64UunORLG2eBr658FOnzkaOsXMc5
S+o5uzrxaWxWl1lCNuRwCAnaAJyXo7a1PWtTPi6tH+hPy8QveHChX/HMiPK89obd
kwo0MoA/OIHe0d4NyYB9WkKQpjfWYpxcAiJq6Tv7LRBLSoirPcXdhRP0jzTwgLKG
lOJqFgBbH66gZVRd8hGW1pBBUAXoBFxSR6aJytjqoGxRhD5B7X0IlUHPZ/hf92qU
NdjpOGcm+tzNmdSelXtVTHpyVpyhVVpkl1EoINnSzaW7f6VYWUkgchM8gjf/ZnZb
6C0p6xNtlmT4cvALujlA4j65qWmxF+dDE5+pED3xfi6PggEZpWfjIwKq2eRZrlnu
GE+ySlt1symgzJxkae8ZFt0WUEk3lORvf7N4UgIeVCSnEm4EzKj17truUa97Dii4
r2kRF2e9zc7RY6td1S0A3pBzNPxF3IdBtkNbNTQGXLezXT63AhgSF4+/F9te328i
v7b1XMclmsl+/uzMzsJyaUOm5Y204Voh7NLqwdfl2fmf1B2SeU9ql9IISnli4+Ku
fnUgpdzfn5lWo5qha+mOvEkUED7eTnkvBsBy50qwF5CHBUU8G27pvK/1VUg1bxC1
ohi0gREWyKalm5O4gF162oMHKb/Zye98fOsps9per438WNysHx/q8heQlsfkKNFR
crBFN+pImLCD/AureIgOMyUCEO4/HJP5o8vmHbCdrynctUJlU4aSZiSwkhZ4X24n
nZSPJDft15AlNFr6kSRRwdSIEyz9d1HxOwQtW85i4oU/7FvbIO2Eb6uQXPn8DxIE
Q+LBv9N2BAAiP35HabA22RigbMOuHsxDYHvXtK940jk5GELvajNI1gvX89mJSwmF
r9xNaGmcBw3FHv0aMiLQHGHEqSLvBjKOsHKNoca0rXAp9lJzT0nudOXTwCKTFVqu
Www3IYFNJCRQ1Fa5brBMgoSyJF5ilWsCXQOUCJ4JUW4hSmhxYCWsQHOKGsOaZ4dR
SwBIGgiIextkGzr6vCBEvkkjS+rqQtgywELvYkWkYCEkc9AI6bLkPqtC657E0AhV
KQuwmrkevTPRkoMRh73ZDSn/aU8GEHBPZ7BGaElHKqMm+ZdTE/Cq4DZ+UF/HoItz
J2FpYpTeJABw1WoYnFU52mPM2ObRHe46RHaQe/dpBUeaX9+fwcds+Q6KYRy6qNAY
f15vLdJTNo2ULiVgm5JiZzanIn2GCvtgqhFvDTrO17xBB9848YGKsXbsc/9tejdq
LTgwXWOtM4sVYPwVSrWrNIAj/UAtlxmXA9KE4wfVs0YDxyYn68DKuiDZbi2XryIz
kSbS4rI1ZKUtz0bnrVhzdJ2GDtHGLjPQkg5P54EDUelvAgh/ihl42zpLGMx1NzVX
ZGEaOSFCoDNBMErrLoi5mJzPndhLcrZ5qDP/2hAsMFBkgu+lJvv2DmyQ7b7fQ+1+
wOpk30CHlhxCdgUPudWKwHi1lGMpEWJAoN3jVam+O4N1OuqL1NAaYw8EkQvaxvwR
QKIlwWAR5mB7lomUWRAWUO8xtCGLNzNWWORpPD2wzSVSzUixrGy7S8m0TIyuMZxi
3poBTmux/mRzI7h+te/cGpzKerc2rfdTH36gAkyEMw4UWyzFwNs3aLEbmOeAn+rI
3LV4NtfuWFvnzaYWGTaJOzrcksDgBe6gveIXAyFPcJgW7wEhLcuwF+uXB7GBcG2I
rXvWV03d1rzddF5ftQLplDNZNFxoPJ6AK9pGz+aakBOlUF7WyXrwHF9rNrye22b9
uCHomA1Fh6Ct4FlnccCa7IkshoS5BcTq3dBtSu0gqyOZmEUIiW8GECniay9W/BsO
1dG0bq6qIfx9Q0dcQ+VEJzAguu4BRx5etpPC41C5ER0+X84RXa+aUzQBG3TpCsMp
kIOhKe904TOk+IbwrIRwfnzFJIEGdWuCnf2PZQzpODofk/8pMxzjM1Ivd93VKjEY
UAwsyKcVIrxOIoodzazY2QKv1JDwkqFPOPgRKKP3Kk61RJ4QKUJRSzORmpcbXsFk
GwrFuYtNlWQgOeretlO8kBUoZqDPEzXGtnoJwGFoVd0rQEA+Th+xbD459JcKWjhF
drfw44RedD3xeVxBDk9FwyzxCIPBlcahDP4oOb94/BNRDwyE/Lga+5wzwfxZYA0u
fQookZRoTesz5w5akqiqVWiLAQTaCd3yeUpaLmxT5AKO/+kxcwPqivHxtppHGfJA
J66gSdrACOa83x3yW2ctUq1T1Rw3+auxCQwgUdxM2Eva7kbFSj88Yfp0TuXNCTR2
KNTewkWVLYaJsFpVwUGNsQMiVlnXyJbyGsuU67UNOcZAo6ZAh7x7ULpa6sibXQja
XddxtIY+yRvFjz3gCtCheJ6HLblUSq/7ELOVoiKh3ATfUAJjo2Gjsv6VoRne3mY9
02ZcSJBYV+K1gvQP7j1WrTyvf1muGFBfCaAICFLJFXxtJHwe0gChYgw7P1PYG6M9
qb0g7iLleGRewU1SzJ167PVXNTajYylUz5UEvR6LAQvhm7xO8uPztEYdR8AUk190
PJqPSP5KdzLrP6Nr3jDhvIcTAMoF3R8a2oSxqdLxP0LIGNrl9z7trTYkr3Y0BECC
2/E4nw7EklUIm4H94C6Zhmw9DUUeQ9fPV4brSsGdMDLkNMsZcsWY7mx2B+4rGfIT
TrycsKx00T9mmfu6licGeE7SO/4cwrSfX3mXg68dx8yxigfVt3CDOC8JyKcy5sTD
fOd2JS+k5/3xFf41hLgLehCC1A/eIeJDdw1P0vvQXHUVC+KVuRxFTaMNQHMsuo2Q
yJomXHpW+Wjz5DFdFeJQkkMWS9Otgkyl7PA4YhJI8VdCZ+QjcDF4gIbeGUkd23V8
Jp/xWzi+LbEH14atrDNInCy4MN7gpqBnLC5X/ayRnhTkzfPwco+MPKIimocHSCEk
XkEEUFVpWf5wHt96PgdSfpIr0yBVaU8pLS4AWWwdSKP8XM3APdSRHqO8nv1+CgAC
FxTCmBV/RXxWLn7VjXqQ6roFTOQVqAg+lAHZ/s0PFuQpOMuNfi8FuNy/PR4iPSAG
vtrYQ1FewG1AOYqtTwOS1s/lPviESpt0hydzINPcaB3rS14JHFVwrGGslWrinsP2
JI6jKCK/vCarICvW7vt8tlcNcUsOiGW0X8V9SqCcv+5QTjI32gABV9gw1pXXexrt
p9OnpdNiB3W7j1gaOlVWjUCq2vNJX8kb84NLL0N99S6604ncHeo1SOp4xBcGklGy
DrCwk+XZ2NSByDc4bIbdgKkhHfnt4biwmV6vFIylrwSBaZzm83BFCJGHBDtQCSZZ
xSvQezbyrlcmvFlTX1qM8NjtArCl1hj8Colf6SPKf6SAvLTnaVNJQajlQyQ2PGkU
o3+Vd+710Jfu51xz3XvXMKPsJJd2Fc64J1rZybxNkxTebTaRMqxud4Clax7HvH58
mq870lUxJCYLvoOgtzFXN3n0P14MOy0bCHr2DZr/xsmXQFCkZ2J7TttQlbOnvKeU
9WhmvoXrd+VnzGBQW+ssPGxHS3TJfhNJjy5Hb4HhpgQ/tH/rf0hPcgbcHYU5tWhU
C7ulciSjZV42uRhShboXLqZapwtew+LzUZYM//Qd820A66TlPw8J7gG3bBV/OOdI
+YMpUcQ+O4lgr4MX09scJC10Oig+9hjxza9yqXX0YMsVfy9fp45zOxl4AKYLzg+7
6xR5CiVUSa4JyMtF2K1FxqgYn7TPaSZJJf2dOaP8tI9OG+TsVLHkLgXu+lrzvUWd
S6End51Alqh1qPX4i64xrfRaZ9sBIZBpPem/oU3i9IFJRLmhVv+o45kxH/7FI8ET
YYZ3ngjZcWt7pXgvlBvvmVchA1G4D6LPtx/A8I5fkLZX/rqaZGCeFNmyabTKa9hx
mFUjKZvnWqCvF5uVSw2BavHcw3ZbVZbv8C/XI42aV17ZUiqd6COMrT7oz86Z8+l6
Rp7ZqCmHDUHO6R31u97DMsK7DfA75X7W5Rojqfuuzct5/IhN/N7pbDW9lCeS4fQF
MrfZBbtZMSiiyjPXEQmG7w1Pc7xUkiAr5YVUhTG1ELOmkyYqwEPrtxv9A21Rx4w2
/qQfq9ULIfBcvHvX2J+lAKm0r4q2g3DqYsH4AnzXVx1X2deg/IQ4GDFD/xS3WJxO
sm4TCac3sJNki4aPtq6ipeiDtPUgSlTR2G+iXg9esEvyrJrmT9RUUiz3Z8FUknJj
xJQ3Ka6OIrstA+LSlr5PA69qOWa/DXKIC6O4fkVs6ds8FD0CV7tBJaQm3zJXLLyD
bRQ5sty9tdBguShJMJWYSVFekkvtFQtz7uQT/kiR+kyVXo+ZEPw9WmOafEJbgDxV
SzP/kTyYH9e3dvT0bq8gYrP+zdkO1yLRbx/M6xujU0Ta5KnyEZXhOfLI969fuov1
FxEnln7CRA3Ya28Nw9N944Z2vEDLYgZMbB6tZzEtCj5QohpruHOZC1hwMxnaGDWd
1sN0PO4Jkl8R7pcBJRNAFwfB8Y6+98gj1oIKfNn++AawuucQVRbS1y1hXnA0blER
27qqQicYXqvUO43pg7UxY7pHvqQ7O+10iMs9dPKVVuJdlUTrFAXMuEUM6fhqdUVg
g5vX8xdFMtdmub9fr1NLjvlAapcxalQ+k/za+yHEfKIdRdPS8U2FNZo5hotngdpU
v5GBrrsoA+V2Tromc1itFKI1TNrCNvV2HAQ1NfiZcYv6rSUD0sU3nd0KvB9fBz9I
t1mkmLKDQ9o+IbVQMabcdtR8SIOnw4wLPY/DbWPZkBQRsaaUVmSiQ13Zp0wn5hEv
mhkPiLYvON3XWZjGgKZxYic7S0D41zjjCNer8dx6sSbZFiHrvhfXsJAWLWbUVrmZ
x3FHSR9EjHrPtk1DrLLbZONtzBRzOu0KlC0Jw0PhUYqwondEHEQuqlITUx5NJ3LR
+WxcSyfHqUo3+th9lrF9Iekz7DSFWkC3c6hD28RvWK6q0KJHEk/Tw2hNK9dp8FrB
U3YRudso1vOSZvqxJDlQRW+DK88RjlTL6mluzbioNNbuWE3p+0OeeFdk0cNAkvwy
Q7yXsJkw3fOhMUP3FGXD3Erv8U3ldxrgUXfjeZj7K4QLAgW2HQxU6oXOsZyueX59
wZFY4HuNzH7ZqKEFJ/02R+SPPvTjnm/Z5JV9R7H0oAw5yYpyxVC9ssNHy8nh3sxF
kYWfzeUm6OLzoSUifPCHB9ZPh8tkJaTtVxvM+Gc/taiX+FskhEta1G6dWhQYyO88
qcWo6aE09d//8jTRD873htaeKhHiijz/l7WcVklcQsxbjeHG4G/lS4dt/36AYZcF
Z30ewiZqTG/Gl8KQkHr+nPnrfib8VOK9IT9EEItaMLb/6sQYin8WkYJAKW2axdAm
Gh/OFyUaP6AMHXrh/DR4Hsom/IRWeck0Ou6aneOI3ZjVsmXV39s/LbqRcPXp8lth
tXy3+7Ts6Il2Z3ws0Iy3tAzZHfWUYEXUUq/Sit5p2B+cJK3QAmIcm/ja+agJkUdN
uvKMT8c4/etbk2GKMERCcIVoehZz1/UGEJgmiPlt+vw8I39Kf3p7C9dsFcOP0D6m
inriUglrdrC+yJebndG4MkTr7KZeVCLIUACwmtX2y61ZLHhLj0QPkjDajNhbaGEH
UE1Jne06m/e050YFQ9trp6XOMTylZ3RjEuwclCbSZbXeSQfcj4SJy305xjVGs4aj
F6Ng/9QODXFz12g44lPHvi5jFn2im2KAhmEf9KfmEzNpnYwivphqv78bp1CaZ8u0
4CHtBLhGnf6mRlkEklVylmmGYIQxlgc99fKvBGCTPVNtXwdDOMAqFLCOOJ5gSClx
h7tgvw8baqhBsE2agMK6HdKB/5XS/CD4UzfvkxTh0ohKHLcymr8SKZ+rqJ4TvLnB
sqviYd9SmgVD/t6/q/GuRo8B84MX8UlYA2PdmcnMS0XeC8oupLhSnoaoicq7CtVQ
iISgVMQ9ppsL/ILEatiSHOK5daVokdyDE5J7m2LkJILWm0RGCvcv+Tt+WV/DRMO4
d2wj6NgsJWq4jjL9o+JeQJpfo6ESr0sYzMjLE1Jl6CO6Q4tn1eUMZKD0pYdVRQS3
M5ScIRHkLTrsTP7ku4r48P/Dgg0Gbk+CD4puDkE3myL2feF422qC8s9PzPlJ2lWs
4nKGMNPnGJzzIFxV5ruVAzdxTUpUqQNNdJUZ4aBvHR3sRFKYE7l+OcKJIkX3dzH4
cUwBvL+oumj+N/LsbHJc8gHnL+ZI2tdaMcPSKdRA0UEsUYqkKq2qbjB++RdKedWE
IBLYtwNWm7C55IH+mRPdkGaZmcuo9mprElAO4NYMQf4AaC8LFj1ofYK9wKSlUwiC
D4AINxs2getwBO3mAdUFIjsbsajYaQ2QQEdiNkealCqCfemSrwVZZwynLRxb9z1O
RUz7l2+LKita68J1IvXRsGbP17JOf+ZqLzx0YNnmhI/tUYRpvXHXJZHoQXBGLELz
XWsidlrS9n7uWVTKio2FSKDt6IGnip0tY5hH7MIcfPqgza+loZjLMoZ3vYTYassH
3erGIJ0OZukqbQtOz3sOCSQyGI5nGxZegjQ93tov4XiRjxe2qwQERiNdJ8rqjn+r
axuD8KZGYysZxHRw+RMURC5stl3YBVqWni5uYQ+s9CPPMrRGhr0vWFjqPb/8wr99
9PYxqmaE2z+5VEiUCZt4hU3peiu7wRfEaX5j1WLo/zQ6QvlecQuUA3rKPntxKEU5
MZOv9ByAWkQ/Nw9PKd+nC9cbj8zaaZhxLavhVG3p4THVUDgkF/WotbhNwOxh8rEY
MrsIrB2lkarS35FzxXeEKiGwnXoQU+aS3QhOxVS/bp2qzjdOungi0C4uomeM4fQ2
2Dnv78NjTUwbZPHXxHXhc0kPDKmEBICDsGKBexGYVra9P4KZWjY/KlQaAzTMw9MR
Ls5U85v9wYqbZJ2SZb/4GPC+CrQePdLqRAbM44xuv/O+Tox6Uu0ZEM1c/Jke+GvL
hD9Noh9dieCmEtKdIiLPS25C4ssXD4jZrsndCX1aRZPUVFk+DD3sYVpiH+3yVkQ2
BTvBgEY3cGflf5s7jG+5aOGXoElCVmEAlSLSM5E2b8wSchrLlK+yDp7eAk/ITHua
fBNZmOWYgf2yIHVVgKIaL5HKu1V87RIzUQ7b8XSOfQeEwuMN58hNNqUzJiv3DJVR
8SgjO3StzQXqaGiBUGgdHmFe/c8U4zOMW6ZkvuGjKuf1cD/2uWei/YrHCoAjwfA0
T+v8h9//bqOqUVNSa+bUBH7vDf+B+q1+HK90uiG918eR7ICY8JyzDoGJZLUpifEC
VDs2cPq9fJXTE2EKPz3NbHE44uXkxpYzGXTi3YEdYsMnM7VQpg7eqI5flxfmlj44
vQg/D0e3XFgjodK3OM/CHaaSWpwcO495J9EXf1iQ6Z5QM83ogz6cpwIi4nkEZ+Xw
i8CwoRM8NEd3aWAAsimTf9aoPQzovO8SMGyIcECFeCykE/pqH8hDSc+d4DnubAAg
zucxEFpP4NxmGoSpqlxBhXfGprTeMNUZFxMzJa1h+IJ8/iNuWrT062ZngYXs3dy0
DfcJNvHWO3mFTsRRY6XGsl4osFGD6gLZQbDOeflN/cc1aZ3unPqB4cXnYwefljyj
MlaKr6+wKSwLXp5m7Po06vdti1cafRRtJ/1b/IEwVuH9+8LijfNli6ciZVKJIU/u
IKTc1R5aH96wIwX9iOT28hntUJCddYiqRYZ1R8hZMM9Hd22n4WuHeMjA83ilj9Az
GASt8yVPIzXuGapEAiTYxvYUCFuapz6uB9kkiQbRj8+KixprrVO7FF00SBsMMYU+
qWaxe/y5cq/EvPLuqlnRgtABz+NnJqs9MIK6Iz+qBHiPKg2a16IQyjfMC9PVOm8J
DQ17VAIVeP/n+w5Aojam0vDvr8l8xZWWtg1hh1XPXd2chIAxI72H0fs2PSesToHb
sNgLJw3xwY2pdgH6WzjM6bMCH+RXB2YnwjZsSF8fs4an8MUbJOeVt47udDcRAiUa
MTp4nHF9GEI9ETRiLo4w7ApNyECSkipP0naAWaWlQUDCnIgAqoZfKMXTlRUWdgbp
J3jBgRHK0xfQlnvFf4cRMi0IPG42jcXTvQiJsFpc0/VudWQtGeTCWPIPHZRHlhcG
lRT05dN0EvsrRmhDslQWI09c9LbtYmxLnKsGLfQDtfx6sMSXAxMFD8mAbQKPVDRc
2uCwsUEyecccyuvbGoTPTAQf0wEAAqlIXn0yLuoD+YUI0HoFPNSa6NiaToFbCnE1
glM+yT0bcA5FIepcUMAaQY9Qxcmyj2tN7cYtq+apK/Tlt81/fhF6RwSSjgYzvFgF
mwDTKKcYE6mIsbJX4vffF0j9KoGbW4D2YbPT8v5fN5L7Y5xTEhyTfOpnklbOjqFc
tBzhFaGXlh6M23X71S5DzbF33ppaMrDi9MAKIJ9rlmVH399FTBNwpio+Hr4a94Pl
YDvZ2KE0b9/iptosmEiRrrRiFCWY5q/9PBb9n6bit0FiRzyrX7cNMlvA+OyUVMYB
sIgaEgGYYXpeOJzsNdD4ZfrducJjPrmjArx99WoNW1U8QGQZC1TJDEQa6ypxsRzM
DSD9M7RkvAYkcedIFgVe86IB3uMuMlCazPYOBVDO1FLFG+YRG0spcXKfwFvx66xQ
YVbANUOJWbso+IhSRdVWI32Pdh3vcnnzFHs4tAvf3AuEPXWoZQxVZ0FQHq3iB70e
69Yndr0YX+q5g71f6FkSgJ1vGZfFsq5Z/Kp8eUGpsQ9UGUe0+xOcXfMOH5c/NI9L
aqXVxopAVxd/6fzcGCZhPz0HwBRM4/F7WC1Xn9W+Ufh5+nE1Gz2+evkQL1ZKLmU2
hHsPUUaNtyPCf/b7Ce9GV/FIo3tBfnjr/DovexBnhUJXVgo9TPuPJM9OPZ7fukzr
2kv+xOFSuAoIKq7Mk7jQRe9iRR9yuxhz+U5hk5Gras1xJKyZefVSPhjrH4R0hQuv
JM46MdJ0YiThr7eim/N9hnQuSkCq3Uj66dMHtqFy/ejBt6MlFLW1EIQMOrNg/QFw
h2XWI8gpvePkIWYUw1vDmo0MEPO6sE+Qvd8h/J8SOVilGRCDNIMwQINaRLfrp79i
nu84WSjL0TGS3HwVudoy7mzoBk2yNj+tU11BzGFkrHCZ9G5xUeZPyMH9AQUz0Y3Y
sn6jEISfINMo3Gecw3iXr/8SyxcN7Y7cNZxpZr7/+XsLqankUa6tQN824fG4BRTr
LyDyEBPJXgppHJ7VL30Z3953jxjNWO4vsUknH44Si+VVY8grAhtAZdcKAsmAjYL5
dqiIuX1l6/tJc3zk60LI0KQLJUh/RrnkoNQx1wAl8Yr3qQca/DlotgyAaefvDYh+
FU+oRgEr3IgV67fZdFgs3U7iKxqb5QeBKdTswufUDZJFyD4uG1viM/LWsABI1g44
Kgb0tGVrxhnLC5fdF8cvJfgQ7hUezg7RpJ/bnrjD9NA3hSt7UovtrP97sRjUeU3U
88iLuzLkmtJ21tJBqbxvcFS360k6miPKUE0s3vV0iP1m9zPVS2aRL8CaYz4WI2a9
m5Zl++NxN8Q7AC0klXO1Tv86dfZXOUKefFQg/wDzNnsAexHH1GPEePgvE2y2uJRU
6i9Zlqdab6gDEnwM8wkKL2K2C6F0S2MHPYhfRZD+3pux+j1aQP6N9+k4zZlNdnqF
SSvrOxNQwt0taETPVb6OF3PEhBxzIqOopyyn5iE95YfZ9pQ0N1CtsWI5I6tm+JOU
OlSfbVHuCqsX9XR1wGHuuXAEDFJhSQ8leBljHzWc3CWi/XwqZ87dhmj6oib4qa6p
fDWRY1aYF4BOETymHpPS2A+CWD789EcUVZkJ1wmHyMtsju9Gt8O1WiOWfIPb2XH5
wVUJAw+j9A9rECK4Zv8+PuDfJwVx9eoxbrRMPpE4ozN8SpJSLFvT3Eah3IQ8MyBw
PHIZc29awV0wYVGWQsAgG/WIPLfKux/OYu0nzHs54AwHaE5p4fGN33/JjF1ogKXv
2GNtpTSwTvGCKPwhmDl/2q8SmrC0nC4vPCyy3y/YCyfY1AFXjcNi/gZRLFSro0yw
uTiLfMvApF3xxq/3n5a01ImRCkHFR131NpAWmtn4FKoV6Y2frhMeUe9fWIYsESq9
x7ELBixKMHsdZ/yry/KjJa69jiKuL4EqyAkgIkfU4w1JMfxEwXqia5id27h1jCGw
3+lQuAN5VjBUU9w0Y9ITxfMvMpDhEo1x8enwiCxtJWcgoiHinUomilN2yD3JnzgW
SWjJCx5Opplis81f2z/vwEO5x3vrn+5dwgpWImJXs9xfpT9xMKHa1nP6PbVnXuta
XqhO3ftD2Od3sPHrd85IbGoKLOMBt1TJ5RZQDA80qiDEtK/2EyBS+KM114zx9xkE
ndlJrMg2Gorni/RDRE/k617H14KjFq7em22Nt3B3UETrwZCJDBjGuW7tMsergy72
58IHzA2csj+nV8OSjOIRGVPZMe8ZrxTYRrL7/ehdM7HLHt6+koqc6Axr1G/Kyyb+
vEE7Co4Dzx17jOF7kPknfrBYdsNP35O54waIZt2hczdMxpSmETV9tIyukJdmmiLC
6Rye6/nvKFtE3CgikZgNJT3tZ13Ndx2lQdQr6eFA0p+QZd5PEwXlBXgtZ107bA39
uqGv/jAffx0F5bryaSvPJG/2WFVwPU+LbSoPZUPNFYDfcxlQn73/TVeVlml+K1ed
dLxo84gMK97i9kSlLxbqR0xHSKhCBXJJWVwRJOzuWTTo0o7+4gNWeIJ6YnJx/GAT
R+paDCNdfIR1LZf6eIwZcyijpUHXDM5T5np6McYmDD8w4lRjbA+KQ5WEWHK3M8QU
7qwvTGkOo62NV/ZXSzXXvpv0GMePUwoKtVGHjQH9LwR8vvgQZrc3EkivVDVa1/PA
XYCidmjOwHyq0uXz3NxusQXOQefVRg+L0ZGHYO4/39Tv38oeCGX8yEEKdZfGT6uQ
qAaxj7R720CkROzUuccwZd/1JWTtCGvz4O3P3wgnmCZSSMWnhLixeqMGjRF9n6TY
A5NI67xGSPmJN7R4PtG3ItV8ZDAwtFKc24sLvGJ4XdXRW/Ni7DAWjh4zf4f+gWIe
4jyn6I7prkW/WcGJx0JHSbbRLkh8CQJYeKuUzhwaWd4CfxZsqXbLgVhSjr5oe+cW
obzf9jplm4YRAI+91h6epE7G0DQZ7T+96zw8Q4uTn9VAQ28zk59XV6aoLBY5n4QX
DRnwTzibC9wsubMomwGYdsJuknzR3PgRH9q4o3tQ+4tTrjrBLgie8qy8bwixDpx8
Ka4C1N9dENdrFsOqLkutTznCB3DEeIk4PZrvL6iBevVILualyVNaGa85ZCllRIvI
woIl5W69sHHR1EIkGcI3VSiPyrXHk9Xcex/LC6HOcqhfpCXQNurcSgmp4OEHch84
jpljXapzwi9O2aEEcOXjeo6hgXva1Ie9vDBIqt7DpXMPrg8uE0tLSMyEbkzEt+/C
lROhhtFvc+UdjAbLRVukpKSmEooTswx1uO/C5WMaNzhvjXxQkkbcmW68eVUHWo29
S5rvCJNr+iSJjesxr46L3JKjJdlj/B/Y8TZzG0kH6VIvtXHKv9+/aIsWE3g9SsOf
9CuP3oUkXZIn5yPNPl1zSJAJsvTDchSE2Mueqjb0iwsem7SiGl6OikxfPaUTNvWd
Fy4MmeVFxXbS6dLiBe/r2ON/JKhkqZockFXTnS4b/r1swyLXCw3ighbUGU9iH/yI
/jxyOuxKiaCyvLrCpzt+D1ogxN1oL6Vx6s95yrSt2I/CpRw75XPLXHBepwakh0PB
laTqDVVHEDvejOJ43ZHf6m4mri3do5qsX2SId28709EsIFGswPC4owTOlqF8TiB3
FGAS7KbyMQR9NqG+/0qo39T7gy/YSXYolvvS7BjIho2uzh1wUnVknjeWiQa7XEF0
67tB4QPV9ry6VBerNuMZzXDXfLxr6TrByJSEv5rp/uO2NzbFqGbhmguBfyqYNH7U
eQtE4lca4qxJmBVRxTGKfK5mVZ4s9ZHHZJX3aTsHOw2165EDOXW+qidsDtp5kFgv
cjhEZjQ8fi1LtCQ06Z5w/RQcujwvHdzlRpyVtmx71XFOfpKBKny8T/17VYlRvycQ
z1kqzNUFDAxdqrnzXbqyPBM+vN1gruj2unGi6q9mXzk/qt/53oSBEf0wwTdsAjI4
DQio0ULz2ahKBd2vZGevN60RtnC4ipIQTAX9gT71TMbuL/H5frmAY12jtvI1mmPd
wxTGQATRo6ArzGuiLZ2pC7FrhPdJ9x/PBN/YI5J9COEE9M7XTg+NDACzljdVK+mO
nkAzVceAIMZcQ6qqLomspcH/3UpTlg6babgfw8ipV/R0Ag7dp+cqkJP+jKCNrBY3
2Cen6un01oVnKmyUSvDtdIVRsQ4WQvK5xm3epNEDkWaWr97lCJW1VkPiEpM4DlMz
3fv6asIY+0bt8ltqpXonUJOhJ23+QKsD5T304nbSKM4lCAXaAogL7EQL08M0UV8u
cWzJWfFoSKDKcOaA+18I0jubPPZyfXgzLQLs8T7jiAitkgZt+ro90OJ85G+9Tyti
iGA2fhIBou4l3mLlcogrStR7SmQe7PXNfgzbxGwA1/WBq7FQL8J7lJ0xuFDP1ZhZ
qkskFgN31k9QitThWRVsaNDvLiHugr3bpm5Es58AQZawomI0Dww8A8tbSCYb7LLZ
9lG8tRs6doetDpskaOplgXtQdQp1f40jlXjycCNqlQkNIBUnIgDUrm6IuVXJR1+7
RN1NC6+dX4RwFzjg2qzD/zk3WDJ38ywqTnjzSBLZb4ZaVeZ6aAm0V+OAgH8M7uWw
lGpoVDVGlG8Di0EkWTL7c48PQiLxrrIr3gmPvhYbocV6RhqEILInWdDsxkl9J8oW
DVE2LUkHmVqZMOUUqPOMhcbdXiE+1kRDfD3hv5OG5WFP1rQHKIz1ZM0ybA5UdzVl
JVcn04Xd5aX+wW6NsDFeI0SZw+V7Dd9zhrPNGvbP7H+cTqVAUZMrSkz1eGT9dIru
Et/0QdqhdpTBkHdiEw/N2jw7embpjpp1URwOXsLj54DDp7o9qFOx79nUCHNdrYbW
1adUGOOeKeWlxEqPWmODCofqq32wYALnJe0QeC749LClI3WXGUrledekMRNKS8XX
tQsNk5FFp8Em+mI13sTAik4kdvOSnaVt7I2HWMNT1k4PNPWnD61sUWCdlHgjMS5e
ysX5xbpSwd8jbE1dZszkfGV/b00HRYoBgVXE52yrIUUv9jDVpbbOttfUK2r9AzIg
hXDv4B8/A89Cyaqd7lbvvfwAkvnQMw0akrSLp2wGs6IMvcIW+ME34aV1kTukdoD9
FAcXRiFJp4EhttXq6qfC4QiVxhr0MX2GS3A5OBGFnoj7FydVgH3aR3hTvQrljQiZ
ygyYWE3nJx7PpdnkzvT3ijvWfLkbhdSh2YekVSB9dmjBQrbJsr0K+knQa1I6NCof
WYA2ReiNVekEj4QpbG2GU2rGAr2uwriF6rlWZ2UH7DStvVRfvbZBJCY5BXg70cFU
kcR672LVpzkDfsI6JUnWjaI/VARGOHEAFIfJh69CBHN9XfkzkSJVT4i9AjWqR3YS
8tG6gLjhNq/i3GpAqZufSVGOudSEmfeY/raba5KFTQ7LaglDaMaJ0zZgYM8Vr5hU
qa8eapw0B3xf+PVV3KZIQ5o0l0C4yEv5cFQB1t4MuhHSJ78yXhxC6MY6iOWIh35P
fNpgFv5q1z50dInnfJZczslPROvBLafwCzvB2z5pK5s/hn9kslNAlrk8lU2Nn0f6
TkqH0kIDxq53NKVHXQrRkcDKEBA+/vMuZeKH35s0cjN+CF1JpelzISQ0s/doId4m
NKtlIs+TnFOErTjd2u62lOPe1fpLmMyyyKqCuuj3rOhvHokAwb1+I6Z8O/7+ZEUr
HA2LfcKvdOxPHQ4okyAgnKLsuKrFLy2k6zg6VSKW1ehfUJK99WvRPc+JVTYLxfGj
Xlnz3Ey8TJ+kLOadrtbBdNXXwB7DiYl6wF2OusH6cnRuNNgSE3L+LOVDA7+1bCxT
AEBMJmWonU0rpEI6DqeMqd+9tEnAcSP7+GJo7VWBJgpZo9W8usGoA1zWfeQ3pVdn
/tF7dfLEGXqywuSh1oloaWX6S2KRiwxrtXegmbKW8DAJyyMrn9GSHIxehbUnCJZD
aRpRqp2cuHSO8ZMXWUtUSQB9X1AcGksRj7OfPXZoXVVi8Eyk7ZVfzNOxlEMyrIlO
Z6Nj9GeCH3Nn4VEWQZIG5nI2bXa2KJAk26tJ7fZ0S/ROaIuMLecwnM/MlRHY7yit
GPbLWQzpedgZEjXEGs1/RhVKZzalbbj3LEpmHTcAmb0FHnyxcWu7k479cQAumWsB
nB/9CkHiANPZ8I8R8OSJe0XkgwIi+DRa6MXnPo1+gZ83pwfpoPhXi7KCf8k9PkVE
sJ0F3HtpFOtsn5ZiEnJSNuhaETgdohLYigp8s7RrnrnX/ohQzWlZt01nsVS+Dj9l
EFV45L5UVHTHW1mjd1Oxd5ARlexZkMBpiwrQTxb3nJxz5KlFYd39at6L1cUcOvuY
VXJW7+vQfT+X8z2EH/6XJkn662ILJGdHNoB3aaXbeI+N1tHUCAL8Px8ExSfEEIuC
yW7KRo9zqS/4agHT2I+uVLnndXSTCAYMAGM2Zk9P6iDNaPx5LYaRvu6NrHoY/9k4
vKGdql7jG4AOyJk5RLS2GYgttHHY1deH84T3EOcAPMASf9eM+27j+ZKE9lSsp4ZW
Yh5rjshGlNsoaZco2IU+hpS8DfBigisW/m8VK3rOF9SthZBFSK/L7x/99jUbkaao
dexqFe3YPqwEqIILxasgzu3IGDUUBs91pVHCAqBHNqgNXObRYv0PTgJSvxo+abO8
en9B7hC5LYgS+THdYxkW8jsxIiZtNrxn8HqbU0sLXYT6WSNduM69Zl7AwF/QXmCH
MhtFIqnljxKquwz2fgaY5BAfEv0X/IVj6m6vF9ZQFDgsc6V92GoOoRpyo10KeY6t
dxTlSdNmy6FQiWigjkg2Tw6+0MmhtCw+K9mZ9y0W48Kc26f6Mr0o2vRF/FWy1np2
0wNFI98cDbvYtGbHiCgIOCAUskWeteB5znVuXhj5XEroAyjSHWF1vRZPNjePn4KM
quDgtNSxX8jseFFamtY8sysD0I42kowrS12H9STSbNUKAnY5iU5QsYxFByYtktmu
0xGLrEG39phZ/xrMTAHj4028IwAJc398imMofogcpYDi1KO6ird5lTqcydsHCZh8
dey9icFir8UAnqHbyP7y3YMWz53LTOVokGS3BeL44f6F0K/k2RZNXPIlQsZ3/Hpl
leeUyQLaz3U3nD6P3Azc5INHO6pQC4OotuH57M52l7ESLZs2QS+3mjzD8pEvftXG
tTBkF9MVNxx376/zSSrU22sox3OlPpbhanYjNv5G5cz65EP/nksktQOX7dCh+/oj
uu9O8+ch4n0JMuorFSXmmDtUTN6pMIDjTHyyIvJhQHxoQWD5J9061wQzSl2+OTw9
XBcpIeK42WGVcFD9RcfqSgK1dIabIM9LB6WPFTeeq/pgNLplyQwp6m4VpVKeDKav
RqKZIFMYfMIlm1W602Dfx414KxXX51RruwCHExGh9vv+TQud9lqCD8kIkrU2jQ9f
cBnE8sw/z2sncKqBlFq4aziK7/IHDPbncobhGRI4bkUAjx5S60vsyz/pWvEpaj1i
h+wnHhLm3yoElB4dokH0X+aVt7qh5zX1ITITEQJR6k0K9U6IMM+zU4Dab0Uc9e5P
f8d5uJ6h7aRh8os9MWuK4kfPxugc61mpcc7tbtI/rK+o1NH1Dw91pP0rxpV8LWX5
TDlXlzZK2DGuHv687jNxH20XCQefhItOOv1Iu/urwOegyztPznt2jkevZYEDRlE3
zlmTGEfx1YsPAV2+zvo01KO4bfky4+4CgV6ai3wA1GWFbeRXAH9gxJK1m811g4kj
PoYB1RkMN3pouv7wF7H0GCOrb7V6UbjJPSmqAewrHIF/e4MknHBKxffC+T7dEgRI
qU6FXnL3OLXl9dfipZNTk94scdaLczUehSmHACZyuK68tBzdAi6GhngtxH4WpWkN
7NVFcHv/g3UAzEYN43OhoIEaQQXHJlIW4itJAsl1B/6HQMhkScjwUCqB+th7Jgye
DyiOICdQodh+F7OavHZOivQfTLW5Fv9Bu+NqT/n9HtBBMnkecpjs9xp4kl4oOL/Z
Lct4HsOinVePQbZPeLtEpzu2OVBAvKy5TvS/qcUoYMRpfqf5SGFc/Kdu5+pTwYmL
7kgvCz1KFgsW2WHPa0jqRY2g5LE8Q6e2w0aqUOerlA3k5Dk/15XewwKD2BKd24Wz
uAO+cDI2rzP05Ztr0Xi+cQJONhuU/LMyvn8J9wuLdNb6yJa/h15T3xShg2L6KVUD
jqPUj8ihSIuU/NJr5L1GMFM6VFka5XttA07dNPJJYeIdE+AoVeRChzlGrKric/FE
RxVuJSN4CEPo9Av6S0IV/EHEAIRRxJeNUCQxvfBqZ6GPz2QS9KmUeW1ZB5z/N/8v
G8jc8ZPRlC0k0rjg9b6Tfi4OuYEzDn1dR1PdraAN11hUj648vB2i4P6c93T9niJZ
JWQEZzTeZ/n/AYKnfAbFSEherBc+bCFlk3006Pm/Ml8iM7xgHBf0odR0IaofQYE2
3B9qsx52gLl8NQKpZ6Qt0JI13OpEYxHXw1OnAjxxCCmzsBrC5tnPgFi/kOTIH6m7
DF+hZhElHTba/xOJ15xsOPzfyRTGXurCryfNejCj9sdHqT0+VRdFLSRFHgsH5U9U
a/rs8cFiYePRq2G6aTfCkuaEQCCc5BOaeCH12NryAtmm/h2a0kt3qKNct2hRev1a
FYmJqy6bp7kCSlOC8Voe8xRef74nGXzlQH9GCI8XuqFQupJO3DJ8kG2e9PWmRuzf
NrcDElmD5UvsR2iLXb6C0rgEmUVsMHO5VzpXQo0Q9pjmUwvq/NcAsJ3gu/hAwHbv
Z+ZXThCcMHDcpdWF2X1gOFe+iiJrJmchuiDNH5KoC+c48tfvRUAIvuPoySFQtAGd
H2GN4u4vxUgNrFlFA+BO6HUTmClFwlDHPXPed2z92YDyDMtbvsqPnmpA9a0WeYWC
WlOrH6qFaQhnqyUK+xkJM0kUM+0QUg94LSUltiqpzWRn/X8AqcpzXNE230rLwfQi
ywQjcMvOoAYX5usQGWhW2rf2qJGMn6sDI43S/FVbzRS1zuQIFOmF1q3/KQy9owoO
o47K0vKMi2Vmrq54YWn4A0vJeLHNt9Ei/LnDEiVG6CWPbUI7uOvDkw/fIjnieS9i
S8EIF/gc8uoFQORuPy3QH1TBIbVxCZXniRe/QAVq0whIx/Qyu/8JafvyGwSSrzE+
tpiCqZXayKrUdw/ll2wMbHsiHYx1QvI5NSqAbltXm1NdGjLls/W9dWPDGfcFIGw7
hYCwqOCGdAiF4sCyzetpRD2mkDnudmGhUm9EmDqZu5ceSHXzYxQ/zKmxhu0PLheC
P/tEIcPTopk8UsbW56zrtTdpOOEzAzr+nS/Q6eUjP9NpAriMsEfPtODa5ryG82bm
p/b2ct8SmW0IhfvauYLtBFm+uZ6uvPLbByzgiyuqmzuJgd8DzkMMqF+OwYGhZcKE
D6RrlmAOrhUeYjJpdcKDg8lyuDlQEdHPcUUjiVrYQovyVB1CajHMxIjqHrcYYR1W
v9OZiZIIHMWbiIiJm0Jx1K2ICU4ezZvnPxCc8TnC/ZnDBUF7ZXc1zc0//OaiC8Ft
sGs5HEMrM8a5gd55IvXdve526g+FlgZgT+3QL45tQO97SuzP0NU1uuXMt2WRGshc
EPr3wPtg2tK3/WOv05kN3vb4UrX7JXDts+qu7ZtsYz6LsivhhDCVikEfvdSq26iJ
zb7GXW+eUItDDNuh2552dRpgtcWfW2WPsRlVznBvB923gLCWWgYvIszDBPXfhxLW
BZGaYZ4GaizvhhmYrwzMAWYEl3SXxWWfeHW4hWmwAX0gfVptI1j2NpPcS60hwqF9
4PyWJiSU8Ky4A1Rv9Txg2Duq5z6R6j2Mw6Xbxt78qm1L3UjBH6nwW5qMiGTFjPFJ
HvIufCxDRdl+nPVytXFaxMzhhipR3RylQwwCnRuXLHw7DLoe+2yk6SJxLsxcBvnc
obk7gI5NVnDy4MwpR+jh4+QGIIltACFFNUrk5cLz2HXNx5D1viz/BPhzKwc84ts6
Yf0Kz/QzdQFVJnEFmQP1hf0YbCJuu0roMUX5Q45F+amEvmopgUtTnw2gpRiUKXyh
vumyE19Nk8WrIBUQfqMaGzYowSjkOY7mvD5vPn9mlQdoIRGgttQNyJcxXb1tFi+m
U89sZr34kHcBQ1i5d6ErqrqyhepiWI/FTOMaPYUhwTDuwAbS5CfOsotP2sRqBINg
Oudfz842dOfdQNrc3zRSHrbq3WS1LnQW2Xr1RpxXDpHZds/Jf0Nck6gwCwgq83yo
KL423vZ4cDDfA9NOS9sv/a9pl2Q9M2HASbLZpRrMYJ99bx61mZQfLfyyjJFp9ymI
ouAOrywzv19nrbT+GV65iNvEWSI3JAzXnQELtlxT+/9bJQfhf+uwetXNdh65Uv6z
bSElNTDFOpZUPu/nujRleJEmGXosMJl2o2yZr7IxzOV5YLAMXleKUkPOohaiCFfe
XetMl4ZQD9YdCdTu1h0eobUuLRCMKSeU5vHAui4EV5KJQeUOSqG+9HPPGASSArom
+ezuc3S63kdg8D9CaYKrYVi5+Dn57SzynD+cEHI2BzU6j6+8aWBIgol65b0fX11u
Dj49z7sE0qwfIynCP71B6cx3cKBjYiCeDVExPYuGZpT8ZDFFaydYXB82oFXXyWYk
P2Ag7U4JRDWC4/8pABZgtnRyIO7oEqEEEr3Cabt8idLnusro15Ge1IZnyRIo5Edq
y3ggOECVqkuMmlgmyF/WqKWT46Hj0HFqdA9+ODh8gP4V1PVwneADYGVZd+Kx0AWA
rz2siOy2bhplveKx1+maZvRvFLVumHjdc7KnG2t85VwtDZHt5utWHY4czgVEmx8d
y0hVN+PsBEagV7NAYNFPfdKbViGoBStjKOEK0nF6mMyZ5QAOg6UEBWhCEX7C0ZKg
xX2Ko/1v8ZZug5xCpRFhtCR+ZCamh7gZ0z55jDxJes5221qN43sVMfHeR5hiS9+6
LbafEtJeQiaumoWb/txhpbWjwfxZe409WZY6HLSr1aWCgtex3X0FWisMNxKbQdgd
0KdZo+DrRx8GpPqkOgKYlzPNMYjxmpbPEITe8i/T5HQ3ghdVnuCB3RFiRE6Zkw1a
BixN3t77gcjl9NARsJs1tlQ50FoB0InwfNVN3q++vuEI/tL5Kg6xuZbn2S51Bt8/
2qW22FSOJzPCdXRhoruBDAiwp8GMmfGWVTrGsLfZsmJ6wiAHRM5fM6BSpF4rnge4
Rq5JnZEPtEufOJ3t/k4rAom8HSkCYdcaL7rhA0aYUjrVcZz2UNmrcRwk3zsMK+J1
YB4VWoqReQyp8tMCk4jqSasnTP2aOPpJm/Bdbv0W82eyj3JUSenKFv+Mhw2hYx6U
Ql6W9aEwEE+BWDAUv3atbafwbKE1PlejHpzVPUAROU9H06Kopv+Y/lBrEcLGtj8W
pKZxLCTK8VN5MuDYEKL2NT15d/TKfRlaB6ktFTsRyGBBCY9CuY+hrukvVT7PZ3pd
StTLWUqt3++y4KqK5g4No/ccqZlqmbe7W0TgyzyGm88/4aw/nbH736E33p6zXGhQ
/E+G7ql25huNEWwmKNyAZGBa9gCX8XqrNNg6xlbV5MJ6ILks5iFUn3GLn8CdG64J
utOzEHKGJEpOeHBVLO2S+MACluq/oRCo+k5Rs0eh7WWJP8B+sLtL7Ck4vyB7FloN
kBqgOhU/cOvXXFr23uoyw5LO2A2e3rD4ZW1R6/8mEwvlLeZyj5LsBnUb77SdjlB3
HppT56wWyG2IGQaurfobK6xyNftj9Sbl0SQQi10jeTk33ItEaKjsfxklTQ7HPZc1
dpjr9nY3SfbpHG5DDHciwOBTGr999ev+dFYG0f4vHEVy+8zkw3R/GFSikqhZAoRm
m0ao4qV4kXnRCXumKOnWAqk1ZnzzQTD/XHsHTOJh6KqixhZV5JlxbwhEl5XfNV2A
P8b9ZPcByu0TpNJn8OpXVfdLAPlw8ab9KLfdwf8FfQYRoJ3v8UtFDoc8Se5ZQsl3
dMl/3IBCVUV38qMCTSBzFNM9n8wXj8RP96oObNa/v3xctt6gJplN6bT9rUgaGmrE
tLB27ogX8wi75aJlxc5vWjxLu/N1CaOB+XtX+w7pKMkiUpv9MvnhKp4B1kkEomCn
W93Td9qjJT/4IImZaNMG/jQugYgZ3NRJ6PiTwZ8SoERzFo8XCrb0GxlIAivXcciu
Wv9dLmCYo2YN0qzkMF0yJ0GUcw+V9NCiIgwxHJ8XzCMfWEH3cqI9Ri6SdmvXtoAu
m9jbQNhuFK6LDVRkSJEVImGOcDhIuNzp+3oVale1aCPLzsfSrzTEbBGGmBApMmuh
yckTVMLZhmfu7hS+2TuoUCM/1TMXvx+2PVJJ9huN0wKFkhns1uuPhOUPlLL3JXlo
srJS3HqfdrhbdY8lDP3HJQdxVzzdCaH0iSl1Pt7Qp1KTlWajo17213SHQtBdSqPG
jTT03mwjph/9VoX5q2hD5rQw2hMOdP4h14AMXTZdgxdiEXVG9XLMbdOQO4HdqGhO
FzLvw/+ps25PWC5gDkwVlDUw4PkabbejL45GdAWDEhH4VEqtHu9z3V9RGnuRSuSY
KOoQTA8gSJu/RegXAwPmHri1cYtVG1rulNRC4nwi00QNLHaXevmm9vCjpCQOszn/
uApQURRIVF8n42GuEmppP6fPawBeCU2WCdLchp+INJiaom1N336s0MtL9Y/lO8T/
hNiuG1D/aMHScW5YGcyKHu/XdSCHKfsLOf/10+iiNTnRqlZQHW8m0fTwivZqUeDa
b6rOO6wvzHEPHpP9XBqafHvnmcDcnFJmlNufxB6lRlNJc0xG/JiARiO1IfzMIsXM
qj03E+aKrClms7RLPwDOnqZhbClgWRow1So9ykIZdYMtfRQKWD7DNxr+ehFhT0jl
COUxlnUOCZJa+2xlVr7aYexjkZMTbQJxesldqC9jGONBJ4OxMmCU66sITTEsewEl
AA6sxsWYMczAt2jXYQa+L6vaenR1eXXPWa7q4Olr9KmDHYTGuh0GpnYn03/DWFUQ
Iw0ekf+v3FUpknPExOAMg7/Hu7TiX517GyHhaDFGEDsawcDoGsi6fzuqiHdtEJMn
9McQ7JqaqDlTFg65HjEkq8lwFwcTC5nZmDQ1oQV03b1J2lyrPEXHIdqGpKOjhVUD
VnE6dw3+JAmPf8T96/w4BHgSLMqsEYRUY5G+OFr1M0IwWjB6tp/gSswd0d6/danS
oNXSKI001HssjzS0Gx30j9DepNPfvY4hW1oYMR0pRo9iVZ/Iw4IEOBzvAtaZxeVn
041M0ggr8Q9oTW+jhFe6fGeox6EkIapMJHfDG4/Dcb2GjSx0fEedF4NdITZk2RPv
cDF5FA61XmvopQZTILjU6qWzrKGpNJkDygdArfe94hRopVCyKjdtXffbZUUxb8re
np5UrFiCh8F1MTp4KaVHkGHJLzDFNuRv/TDL72Yi8eMhWplg/cM972tHvW+O/T8U
T5HZexO3mOyT4y34vpu7lvVYHaFC12A5gfiKJhuuADloMVsl1Pr2ZYuYfEh2gVDv
cU5e+vnYu2KSTIMJO4rtbLG5yvRHJbNqHTo8jkuhMyomIoNTjgGs+3IZ/dGkxsNR
v9NZ26o2lpItndIbPoAPEd9nJ/nw2F1t45/F6yEAySfgTjuG7P/iLJ7ndMIHb55S
aXqAjn6PvOYEKWb26iCs8V2ItCO7LBII5OQfFt0kzoKZ6oFGi7VtULCapb+YYKaD
vkSFKDAD+QeJem0fzUKEbKunXDNURE+QzjGCuMY4iTK1rPrlffDeB0ko5WL4fxiS
bCOdeYEO0GEa4TGfftqNDRZlHhNM7QoyY1oXK3cnZMQKoE7sXKf2rdv82DT96CYZ
i80ZPI/NtKXekImwNOU3PvlMVx52Eo8V8kq0aMbRIrnAlv6RQSbqE+Gv0hfE/eKJ
xIVIagaSPo1NlHgsQDUJ+ILTzmp4ClrvsjDl8xYqlF3sSVB6jYLhrb8FRrN/Onp3
rCXPy0oUY/jl3Q0gH/0DWw5c8RN4eCoLJvy34ZFnPIbljLT6OHvpJYMTbROGVue7
e6AwzK6MdxP+uqsMQ7+UM6f4MGg0dfNQyJgJlzICM5fiON2CEmZN2Rukv/qAccNU
a33JuBf0xE8EPXJbb73LTGfjmqHWR5fE29Z0Y5AuA0cYGogSigy+kwzCI1eeUPFn
ndggNOrILFtFM0FLy4afMyhZ9Xaaemkd8v3zW+ODM8xSJrrhM1xsRaGx99zaRhq5
JkuMG7/ekl879NBcF3ssgtIqA52KNo1fDTBBrVqKWqx/V2BbZZxXtS27njxfgwzF
GIzmoTCFggAxBrX5jPkqDX6xhhmKia5HA0WUK/O/l4UgUb8fp02j4dIDh2tEL+xe
b9o418eZtRpavDTBnqkX1KwfhZmy0ADxzviYI/P0sXgAlVD+fuIKIMHALliH2BFL
CRlqKgs78XCJpqAN5l1AUFik5/IpL/NBfLy662f9JEwMcmFnDCWr8R0RKPH/Jmiu
IWTIyjr844XdlVyZcDLhqHkePST54i1g0ej/Hc5tzu4IbKLgdZ69yYz1zX0znJD8
0pyxfIKmZuxON2YkamIJLRa9gXJ1p1Uu0jFcDScyl2yGsIjepyEblJL5OvQhVbHp
f6kHfqwmzStKoMzRuQOr3/xO37FLXhha+9QosR9UoFmCsonjB3fQIXyQosr2MFMm
LI5ytLPWr7A8JqfxP9yRRz1XrVTRnovBG5kT5TmnLUMvrBVNojO1i+HD89ymyv9J
plBoCEjl0NgHtQa+9j0k2FUSTC0NEDBe3w226zXDwAMRZNyjGVngn9WoXJaZtUK9
9cMt3MK0AccMKm9daQ9B4xBm1adW0prh/Aj5wUzaGFmiJQZKQ5Jwuq6Ts5oniUd/
B83y+xzBAm63j9SfJlydvCBXF0PvQ015/GNA8zY3ZMOOLyIWXvgyhlLvrn6i/3oM
m1q5wk739uRapjAdweB5TMI13rZX5FXy32Mzhl+7RIc8kMqMP3MjgpLhVMU2zAqK
AiDzlkC0V370dEEcxKJjBYe8m9BhC8EJ9XhHLxHvXpjQ08KtN2jtk+r91jffkPAw
GbVyTozpNkG8EShExU7OnH4xB0ukFTwYq+mV009dQFvIjifUVbUy1QO08YGca8N8
Sl6+c7DSpenINCA2P6x4vMkrtPqxEIxKXnQCVM9Dmn2bCWkQtd+OlX0kgDqRMmRV
FHsupP0DsDezGQU/Y8ejVP02s/y7Ws4AMmGzE06yHUP84OCfLsBWg4jS5IJO/Xu1
AYgydJmFS7KPSQCaDSXdOPs0g3WOdfmUQ+w/Rw776+o3pYP4EVHYgRiJPCpLE50Z
jw7DvP0YksIny6Au5dNN0k82OnY20OhIRuCX10D27J2JfCBeMp4J+5+YuYO/lFpH
Nff6ybXzwvF9O/kyoVUpp1wIHxR2lmx7athutlhP1EGzqS8MiQEwJDMehb0H4xVj
b51DoSEI6Mw0UwcBz3PNQvlj1AL+1t70Ujow1tbZ4wgg0aciIs9Gb10ZbXDN0mUH
IGZ8La+3pt2tSEpjivAkJdxZt/AfAtinwQwH7fjj7tYphn5kgPzBU0+s4eYYKSyM
Lz2xmt9NHRqF2VZU3Qis7J8uOfTS69VIG/ZZwywGqf9w8/mj164y3AREMQLc0JBd
7ArPZMGoQpKVUDoQ8ZOvZDkNEOztkzBFjW7s9qAfyx+/32jnPtmk4JZz1+kaRTfi
HGKsz3CnYvUyLLTyRkx0PZRkpViWBndCXuJqalw7q+BatU8r7N0scQ76jBbcCYpM
tAPzW3nkHXepbty7yZGnPHDc8KmDxOooaZqqE5ll/PDx+oovt6FuA11HY3gJZIb4
9DnIVqDO3dlASHy/SNuTWKOlv4obOY6NsFQ9hHvs4crUUmkmnolQ18Q7ovK3Mi8S
1Gdld73Mhn/VdeQ9B9QS0lI2zJM5mBYbJLsPdTS0YIlJvMmZARHYyseTiKxzjwqi
NDAOSfQd/ejM44d/cOLBBozRsNdN8aRD232acUSeTO/QTdUxcWVjDzDmeXO8QkBz
aSHreHLv2dzPDeV83dwMTB5Kwr8GfFZYZnzWI5xnvy31hnlA3jf57VVOEB1dRLAl
3WsTqKdqNEvpDVwxKHFoiGYM/bNWxcIFzEvEOSsERmjXdr3qJ6caewW1crhnZ6U7
B/cwnMaqgaevhpZr35R3bg54OUuirpedcf6smsFlmlo27/BlysHhIzXFVqgAX4BO
7SICNihHviQEuMbZa+1BCO2G4GZ09+PFKKuip8BZPV3hBPL7fmUxnkmEXg2um/fA
pLmdM0TgeRihcNSgh4UiP4/5WTJIJi2xipw7w52yNuh+TWALhCC3zA1ClV4tmkkR
/y/HzjbmWNRbVFYcC8h3UEWVIloSuOru/hKIJexj0xcGDmtMMGKwLbzqxJq70M56
x39mJaZFuwtyDdFHTjutcXFDVyHGnKaNB8d9Y80NZVnG3X5PVC2m/ZTSV6LrUBls
xdo90Qe5OI2fe1ieHpx25v0Zmlil4rsxF1vU7rxOitp7k83TlAYdRcq2+Ytpp+n9
rmM6iU9ANH+Dfqhh4jCTPyEYn2cD0Rb70JWmmroDnuXJYmNIZ4c5NYOaORE3B8AW
7ar9hjsonMXyDXVLj4GqC2xwm4LtCcQScNo1O0ewe/5R6dclKcUBPcUlrYUZdfnb
WYznRSlLgrK5cRxcSxKO/N0sYP9W8aKre8ZPc10uO5czAxF2I2+K6FgNe6728e7e
WTVsHxxhmBjmBVCvcgoHBG1SjCfbXYEDD+vnZIvd2U+iiiiS76dAy/YOCvTuutaB
FzFBw02AYct55EL3G1asQ8bBxo5SjjuZAaav+qa7fzv6IUdNrwB0rFekT/Ky8JFy
6ucEqNFF5Os0htpg6WMc1bgNfpkijovhlCnIrJAgumbCMg8lVb0HbqBWaM6o7nWL
7gr259eQvaRaBaHUB79lXtZ4RxUSGzBatQinU47P2lWFkEoWw0wARayGkTXya+Bt
gaeBw1d3L7pCydwQjTmPuZ8GhiRZ0+UGLNzz4ZOxpOhYZkqZOeba0f39IvgJP4eY
EG9mhIjw9UdtTpkdNr5zURHscoSppvfQsTN4jaeAYk468xeW2XdWL3ZQXMxhRpCR
3ahZc8MXjheE0KJm3ptWP/NS+3cikV8AhEjLMjrJ+IsTBS1AeTZMheH99FSeYPBV
OIphNtHPTrjvqOTr6b3g7HVk95SBieTPbWxKSoSE2ynUFvkLZJmWnfkGzkzL/MR5
H0oQVh31l6TdZFKYDRjyqK1ohO1+PxO/CPCgTcy52HXUi5ZUUSEgVlSHfG0QMNFx
tY8DI0stBVuGzX+aH1z2RPGvFm4BITk1nsE0eqAhwJJ7teYecrg7HC26FHRHxcZu
poZivkqIajEhiMp4ScJrt+1LJf3kL0QCXYuMcuQVlAUxKHSNjZuI9SxKUV4g5N/O
0cHinjLTgHwbXa6ZfG/nJeQGJpcW73RSKELiYFSEWSmO80GJSvUX1A2ogxZHqfIu
+BX5TLd6cuOEyCwX01ex1I//KV/1rhTLP/u+IIkIO4UHsyMfoXs+HBhSe+Ji200q
h9eg13rp6KdQs5Fkr7dX0Za5ukJaUu+oSUZWcOW72HQtJCdnHjozHqA1gs4KEWlq
WVjWTcbOTmuXoGPs2nCjVbVd0VwvaGgwsu9DasgfIrKJLShAqdZGj3iWYdT84V+T
GMrTxhxqR8gFoJSxZyYr2i0TpVMG8cL3kAJKYawiipWGxwJbNT7tkANIsPD/uYVD
KTyOS2vq9fT2gNvMjQIClhkH26bbxMOxIGgWLtlZRblWRt3p/S1O1mpnBuS2dhCo
aDWg2TBRJWJm+umDrfMNPbnTHT1Syaoezwg+OcQoMMedEc/hYsYw/IQY3Qp7C9gK
QDMYF4dASDKOirAFGprRyhi7Gj0GHLcIJncaPbsPmdfvCsneVvu2ARmOTmoKeHCU
HIoFPJsq1kS9RPHXPz8Lj8dG525swf2zAHy/jC1j+W9fxd/ugTo9nEmroXw+7fUg
reqOTt+C07MbbRfSptkEoLvCrNXyu3HuQGhvDoIqNEjKhlqYk+CG24MLgbL23ZDf
SPEz3VwoY3BvVxAAmF1e3VjhRGg9tSCTSb8fyz6mgPPx/gYYMwh8J6e5HPT9eIut
B5Vm1JKpMCeWg7JyVhMlqIlLDsf7EqTWyaEEG2rN8kuGhKATE7YGcL6LeqOVXmX6
5QnL+0j1T6A66Eu3RE0GCj7+nJimq18ZoaUO4SJ5lX77WAXdpHrF9yqEDupiKNeH
j5Fq+xxZXSDISOgZsyBzKFnQ8S42xEeGUpS81+gE4enGByWOq9rbfsQUMHalZcUH
Vb5UkloUi4JuVeJUbhCRyzaSKrJ6FYSV4yvn5vF0c/UAmiF7XsobHd8NOksdb06o
4fdb1KzBxIHXz6i85rgZQqINnloyP4fqdKXiaROWZ6wJw6Q90PROmfQqlYNWvC4Q
KMb2MDIKZBJ2ToSS/j6qI9Ga9F+1iDCi0dI51u0jFAcg3sXqwILcbPfLJHn6+7cR
2lZlwK7aF5IRxhDULBO06syWaJcqx4qVZSwbRVXbUCyUANqfpTJJ3cEsKG/lheRk
ydGstaZEGPxkTuEWiH57q7W3JFEWs8z8iAKRzkVYLtqUErsK2u3i2PVooabnakTR
Pe+IaGKLzCCwVdJU7D7EowtJZG+NnDI6u37Yr3Fwlw6RVfKsUTR08EkKMBZtpWXQ
jAYxmIFxu6mtcUcmp65wg9ShUCyT8FDIDc+CetVI8I4B/yHH5yo8LX01b2gKFOo4
YdDUkvfI/PgQCtVFLsUZ/8eFdV+IpCYtyuPr30dgdee5vTMfWKs0DG4FmOYgCf7k
x+8qakvPBJPURXNEVH9dfrKrLAjTRT2lWEmkzQP8smNJAfVF3hnNxy/nTrN/1Eh9
DnnbtLtGXRBI9vOyrb8621pu+bnsQQH3uQhhuk+sxY3lRodauTUoZwqTUXYhxpz8
nmMw0j8fxDxOpq85/MWOJ5ND0cMH0Xvp9Jn6sixVx92slE9uYj8r36uPMp/7NFZ+
zNe8x6jTWJx1Z4ogrj6GM7GxCwuY/Gr2w77P6A7UGg9Jfyuacls1r3inPRCv7IAc
czudK2XUaqZKIHB1nGJE7pjTeRpnOw36yN8us4S2acO8Nva5gEPMQmluX9fBHvH2
1l7vipiBdmfEvDgN6zIf2po27ipYbH+6JYCpxD9DGWjzhcNIyqWAxfqLOCiFuHGp
DHqy/+2LwO+63m9FyEeAFeArXP2FE2nIaN5cZDvBIArBtAgWeIawdgLbdbkvHlwz
sQbTkmG9e7hob7kHH/6nAU9tR/r7ZPcGBjKAzCC0kSKWIiR8PRbBCw3YB+htbcZc
p6pg+WfWt6igR6SsVJehYB7Xc1OOAW9PxC06heslsENAdxh/ojHz1pqMcb+3Wojd
aOR7xAc2eL1oaLyTrqLHEwYvdIR3PvNuIGwDA3eey79/8qnNJP17+gRoFgA2MKfj
yXOSgzI7HTww+ddwgcZOjiuR5hSf1dZ1ubwHcip1xnh4Cb2y1sXGQIQk4v/RgAqE
7TT/lbMfpupg2BPFPFl13sxXXnV7l7hgMnJmYguPnTpsEFC7d+s9rsWlplBJ0W9R
MXSseZY40TfLWC/HraNE2t4AjlVk59ZybwAaXIc1RPD5Z3r895qM7npYL8fNJ//e
571TnPwdLnTDw4TlrPpOUrB00/lCOESegtefKzzPlc6BBMidJmSb2DaR3SOHX/sA
HQC5MslNP6p3jl6ZL0DGTAMNX6dsH3u6v00OVSVR2R598LAV+c73xEIHzJxjLsvk
Vtfw2rEN4jHSztw/wIPKkVakLABQ4bFRXnnNWR4gACUAvPwvHY24+sQsa0RptTok
dbArgK2jIw6HTLzDm//f/LhG2nj6/10zjWEknmLjwnNyTJ3NOotcVh77C2qkJagS
No6T4pgexroN+snXhDsCTpIbJCRlBaLkjEiBHHu2gMLXWYlwWRW/QlW+6bWS4s7y
aZ6O5JKDIwUzb2EfxjDHhI6jD9KoNdfYhDdh+8NES5gOjBHb05K/2fMqPqdW1lt1
wPvqj4JCp70EXe2Yk2pioI0L2qr0/A/oiq/g68xaToYBCPytIhL7hXNs9wKmy/8f
XU5YrOyoU/kJNMqNpVyy5XYkZ8/2CJeIHN7SZIbSRkeXxEK+5ZazXYwxukos7W/q
x5pFQUoBrpG225G86NnHd8gzXEXeTtIcrmPwfkSrM92uf+QKaDtyeHXQBEuS1Sfb
jB0WPvAwkFp9zBZMo4kMeRKaZHt5g9U2B7XC/2RdZDWP/KSsHLOqonIYag0kNU3r
fTq2SyqFETdcsfnjnTJ1JQ25z/Q766ZN/EWqBXCy5vgDrvs665/HP08oPn0Ut2G4
H6JCyVU5c0+jcbCUfQGa7yk4twy99lYjbcc3AmrgtmNhztH4H+XMCR3N0zPMPKrW
Ex2/129M3KCFYVczrD3yoBCmU1LPypIKHXcNs5TO401k39RJ7/T1WynW6TICzsOn
x0On8T+th72de+MxMJbdiUlSYMxJ7SA8qksPeNkoeKz02UEEdcjPecbp0ci5Gc8M
HN84gLmpAY7XSUDiW2C7BgxHs0ujpnSiEo+/Or3siUw7BOVV21VargTA3ecNBx4v
RPpOTDrXo3bD2VSPpHYvNgXKRqeNyyxFsuaUHj9A9tdgrjKcqs7t6Pps0hiLpKYH
RphHLaX65Vofit7h+o64Q1BZcFQTz8ZJyTvt918/uy2cVaQx6CJr62KjfgJYRsaz
OFySLgFD6Qj4tJ/FOgEP5YiiaP1rsalxk0N8StvGRD51qsz6ykLUbahCEElvsjXC
4NJJciJINuy6Xv/wg2VSOCruha0au/XNowuEz5GndwsZvmmZ8EOHcjmRI0HuBbuf
4SYlFFXTG2pngNbKtUAYg5wrwrvJcFTn7ZN/e+mdJ1tSZtsvhCeuF1cp0hACdU+2
lQuxipoTAhf5mVuM0qtqGUPNzanNBbF1Y5RaSuYrKVdpGy3ZKTodCqH9OMpL0LM2
UskndowUJ+z1R1jyyPZgZThirIO0pmfOTZQ1eecULLW2HQGCeQbnqp5RCuE6RQjG
i6re+vchHU0GR3N6yb9o+i7eevsRQIBRKU8Znpk3s/HIVsmMY6Gf7pLGMEPiHPIq
Cszbh9TyuH2nlbVe9WCKs1sIRyPtYhi2iOmoUwG4jaoCaWl5gR3RDQXIlNYrzoAl
/dLvxFoCibt7A53RcFM2vr3ie20XANc92sDxG8lc9EYGd03jFJ2/spzwTg1TGUsL
9CL/v+IiNhaxQRiDxxGwwRbRVrPtFLPjlAckxFK1F3rEN8GtmZTZTo7xmHdVSKjt
5LfhHofVatFrp+WgQavjmr382dVq1bgSHLX4vgDoT61KjiqW70EuSfYhoyA/rJYA
Tt511uw0d/9AKEUK8ckGpjUO9kH48skVkiyweO8t3eVIbUZYtNbVcR04uSCzzyTV
NHROMDT0ZZcieXhuW3KpQhs/R4woSJA2RBbiBDGkF5wL57jXsEtvkk4eL1bkAw9m
cYqQyFafnUxEyG49rw/TKrx9gAMNoOwkDSWEWAB8PI1eJFGhADCuGnFWhNioHYZT
cCef8VWi+NcNkBoXAP4mN16FutWQQiE9bGEXi6q8+GFY/GcO3j2rAHcjGW/Cd4iL
VKxPyRHifuAE63A0k4BH1KgzRl4iYs0IcVbvG++4hICecYpzG5eKPsPsisuX55qA
Dqo1AANTFUHpXIJKME/k3y62jn3jHGbAZf68Iy7Bef6LYRdFX4JFg1ZrUuW7I0Xm
gd/e+QxaSnZx5VozNe/8d+2NJB3OyrLeHaofkY21+XgWl4DhHuCr8he0JZ6n61Gn
UziryIvzIzMwTYIG6A1i7JjYF9/04dNU1jXR9iwX+TuNmz0DLke4kE0YxYwFt2eY
gvOe5sT69g25+fm1VYe35HZHY96dqZ+hi9cNB4ixY6RuzY7Or2+tr1CMeqgv5R15
GAct9bGKMc/6j741FEKTe7zbdBPZ5q3KpJr2afUbKcvAEw9MGN6zCYHtY9pIng/N
NqC3sPZPxtpS9Bgpyw55qYvx2J67SLHxKjB9KeqRXrxZeIHYiN91qiUlh/oiFDO0
MKn0nQ+vA+u1PaldGGf8yOolAbdsFdE8dl7unrFOoO+GKSfpfBsHMwEWOMlw2X3i
SY6BNuPt9vqBSliP06UaZnRylcmEn5XjboyobQ45YvRDVJ10neZS3NpbETN8asi+
yLpXLFzUu05OiB6HjilanzE5NUlhGDi16kN9Pk1z0OIMFZVzg4CvI/BWEIKkf7oT
/2IRm61E8KuS/uYuMYP4+8lpjOPywGJ4Ee0R8uihUbSmsxm8E7XhcWW0D1sJKeei
k/5lIS+IqK1pERh9kcdaVeiSvsBYYfxzfKVShBQLZOkAgwfAXtDfmWCpbBsByQe2
c0oNoIfq7QvV2SI7/ai/n46zvpjCdgcH1Jyy73C9h4JX3WJOvmo68hgv320bC0el
/W5qv2cG2EgHtSIcjre4GNkMqNKPD78O3V56VYWY9jQ9pRd6y4Pl2DdAJJIIdVDN
2iF2zEaYSmxGJZAMXA5TebKefY+884WasHTzaCgt9QIxDvQVBwAeZwved1qnpZOf
HZHVFDmhmLMYMBvNeJsaf4GBggeKvZDH870lcI+7eL3s+NTda6mny0YUQGkU6aw9
No0A0lmQ2ki4TuxAYUCJE6Vaf3EQN3+Pg62w7KX32wxk9aNAguayN78/eWpJ369w
JHxIPu1iCYPMLBTZa7Yppg4p6pke8sABg5ZNcSzH6IlTZ/qy1v+NIYSsw9x+coEc
o3lzBn4IdDUarYbjEHdz33638w1z0OEpNt5osXypLJ0y0fS6TNtudQozsdyd45eq
kHKbA1XnFSkr84JijzANdGD5m2AYpAKX61AG+2fVwCzxsVRhK7k1hT/blcoMmcYi
k802zeT4wSjJ58IbRgrc9Adq/IOIoEcHynQnzzhJbWgvbXJrkM8vMiqUlzVpuyZi
bvR1d4svt+HCIeNqD9p6ucHdTCK3p7bFJQ6NjREuXewwc5CaYX1lmTRKz7aWxdRz
81hWMEt0CnEb2Gbd7+UuK8ULxTuqtj5NvpxHhbFVJzTbhG1LYyyIvDcTiA9boHWG
UkHLg9lw+mTuy67PzUdqqFkbD4Y5Qry9kAlcFy7w5tuoZuGHeBY/BGuwEFhLDAHK
SRmskbjeAJ3IhWl8czPUp9+yNMk6v+pLttfnMNB1bU6s7oDO3IAd2GV3QC/h0BGZ
w2XsbOyYPTi44vo1uaSjfg==
`pragma protect end_protected
