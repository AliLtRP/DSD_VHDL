// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:23 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
ObAnz8tJvNv0mmKXmsJBKSBQn6H80dGAJEDSi2+hoURAmHjasVdiRhv1sRYY2T5+
MbJp7vIMhB1DDAPPCALoe3L19ycPKELeRn/tIg5VahH6s4IGLQIhu8l/497jSkLP
OLbP6eBBS7ChA//+boPClYwuKjirgkIsFK99Nx3HXBM=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 30368)
v/rl4ZRNuwbmigsJlwOXPmU9CVObsJU4PPGClQIJSOWHTuxHjYQd7AhekcECH5Ea
TsaU6BRkRS0G7GvHMgT84/Op9oDSvlaFnL4+xLW/5LWVV5fhTSjfDaDhXSo/2ZNR
vlhq5gw9wkevJDllweBdJVsEIhtAnOeGlAi/ktNtbf5L7b1arzT8oh/76qT0/ajv
++MkRl2dLuzE/hcwBfN1KloPMsatuIdOO+rwcvPcPtzhspHKupifNSYxaFaxrfri
p3p0cWxskWQSFvUxgwZkFLoYdfZXGA9+zgjJbJ7lU1y/FhkpuiGCZiLJWbdBcWfq
+fxll1QasKAiNYreNYtY8pqH1BYkILFYlS4P2ilVjqyywlHLL6SaFAReywTX39D2
3JO2jkes1q5e8BYpTBpGv5h8AFZLiqDOnzT0fcaRao7m8mo99roTrhC3NlzZlU3r
NO/ag6uuR6VsyAR4jBeuF2EKSF+PlFAGJ7GRXHYH7tf0qYE7msqRCoG/hY3eIyUY
fUJDFXS8QDeb+GRHfwREfB9upG05vWM9i0HhGRqGOcO0IzK0o5R3q0wAFVpR/gpf
jc0/OLle7uIZH9h9s1bIxgBp80QISP78Tfoe2BIbjFT5A8IIlAXoGK0Xo90Y6yES
4z0PxP0QfLx/uQpLa5jvOdJyVuiqgp76OH2z+p4mI8pHHnjlNrTWljpF6KbC5s9/
Mt26Ct4Jp6GS0bw2ja8kuvI+fzSy+BRY+5QIZFVqkVJ8cRFcYrDWyLQwmnkO0Q1d
E0osmj8vPWi7r6osaBbkxEWCJb3SIhy6iqpyJkNxUNvDF0eCd3BdGBsmY46u0Eep
AOEq7l1LD7of+DlbUpu6A7Rho5haYH9QjXl+H6bICUyXL0ftIFoHdsZsja71YSNQ
RbL8ns9rt+yXUjwj1k9JuIUY/cbjTslJ9e3WMgNTJPJJsR2Q/N986/X8+WnvmtkV
evK3Mqldfj1c0m2HQeDyDYF1Lvvay/z6wD40ZPh6vkKmUA3t+WutqeDyvW/9+kIX
OaC5q2eFzbryEY85Bu2VzH1KluAkwQyjw2uj8LKkWM8My/GkhR0Xv/FINuYh0WSZ
kjwplaOzsL84fTgxNFYOZlMMsrCDpHXJrf0cbyGs3NdS31A/ZiVwYRCX6ZOE8Tqd
A7B5R9RO5sY4o1rV5Bz7FrBJAtlNYS9BXunyMBSXAunUR+ryiEcjPYFjNnp2uF+w
u9aYVUBY9gbQTbjx9QEVCYOW6tCtZEqtLrsI+1MbYCdKhJS0pBFrYjl3rw9Wz+Kp
3MYjmYLAFfmVaP+/O42IEjEH3SZk2mJelZLx8ldz43sIOsFJG0W1o33qb368oliq
Rd62GKdEu+wn2VXIFCAJNCj9zX/oQudT1tMk+fABbtL4zQpUtWbePDDYwCm7vwNJ
zadozRDg7I45Nd0VEqNtJmZQaJTXIAL6ZRJYSfcwNc4OwNPqIcCV4u+Oe4Ysyksx
kbYVvZJ6uuzu3Af7RqOQUR22bsQghb6bYrCRaiStwynm49VFq1MaWZkWmxdWSiqd
3M4IHVLGN5Ml4M91z3XTTSTjW2RR1QvXwVG+zH5cOeIkdgRi98okRXBL/yYOnidQ
beA/tlAutasNarkolRTVQZTlyx5D6SNTinw88644Nzip+ixXa85VVgCJkXBjpS3j
XAknfwfxogxt9Md/uo77E5MMzWyxl7QnOruI7u8IJZ1oaVGZrMNqqtQZ+Cq+TX3k
8JquEcppfGq05U08Tb6IndYRk4L0b8Xhd2HEfb6CPCfzbtu3pfjxW+CvANR/692T
zizLbiF2EFbdT5NQ/YrNWEOQATuOnkR3D70y8zTyaO5ScDi9Hk7SJXNZDClSz9Zj
hgDLAfw4XuFjMxVB3CCa8IYjg8WiawiTAkzXYPYnVRaUpZoC9AnOXQ2tYtJMH4DE
r3rfnz9RKKDGIW63iUwR1bBkQsIZFxkYFgVa2SxPIs3kKxbOgzBpsUEwzNnr38X9
sMz/UVd3zDkKxkxYLJXN0esbsCNW9rJYYKk1iD8jRfDtpnvCP2hY9iGbmp1Dj+H1
BiwG6yl8i+G2S9xIFY/KN0AO8IAD7f7pqJZuOYW5ipDGSfR3lawVa3wloSSlofNc
RcpTGpkm+4xQBw46euJI64qCkAzLUNOt+jkb/BUy7aA5EkK+N1qjZw04SfRwsPAT
pVpRy6gJCDsgurOrxkF/qDXN6/xkhVoldq3C0OVLrRbgLimcro35aL9Jvp8ByFyA
f41+t4ozuvcXybpKnva0aY/h2y1gG9ZGRsK0yqsshXLPeNyFEJWO/7SGqwvRZUtI
kcxaOKLnw6xnlGXWhPaUdfMNB8D0lTyaPwFwjwbydDWnZIkOJ1vTvX8v5tkeiCi0
0M/WfB3YM0pUZbYoMxdlbw4Q3gIiMojTuUOSxd4QlwVaBmiz+1B7o5/LMKW3lglK
WytB4+xB3nxGvYkUTRIlRfy7MsGP08UKGrB9s3vDHGPxEAi3Rjsa4Y9nv1ugxk0p
mc1AgLyWEHw5FjQg4rER3bjCS+JarRHKgxYMFfsDbLZXthEXgZzX9gWJ1jnVBL7X
1R5jV3nhS4+/NmKjXl4FUhwS3UOFgsQ2pG/ieKeaVstJ5CZM3Vap4qjV5XBPHuzX
671Y/1l4qpJSAL9+E/NgmPSvb8wbkXOc6UCtxqqKyRVzmMiuwPfbq5nZRbT5IrV8
RebEqVmx7ZnVC2rU2IEukJi+827XYAkgBHIHHAmM2sXcWAblIp9ivH4FVj3g2HpC
TcIZfee7jXFxOARsS1L9FIO7Sxt9cf2U3VkNeGV/MQzl1t+/CDwTFZ7DJK1NR7vV
qRxE+BAWRjB+EOKSP41nQczHhoIX35InKyXA1mWpA6XIYpcgO+MZUET9lVNSxTqW
0gSmQ2vUAhatinB9Vwhv+Xwv+Rg7SZmG2cCS+7Gind7bXxOsH4H4KHRWUfnoc4F9
tyovicdOxGmNZQaI4ax7c1LABqA7pxPs2ZaDvnaC1Kkb7UkHzOlkhvVih3vr6wYO
EqqBpOIPU1ATHzuy03OQbYW+vobrJi51udUcH6r8xMXzySjPakab1lZiAwY6Pq5j
AazRsMdLl2INzQuS4EePYBEUM6UtPL2kakL8mMbQCYaDj1uuGgAFNWjsF5LRGYs1
jV3vvEVWm5NbkiAEyUQXKvbPB3hzJwL9ZxInguAJL443Hl6hH34dI4BEQfPORv7Q
p3SeE3JuD4n9rRXpWwZzFcTIq6NK0a7wxtLM/in2vQpkDCM6JHRvfZtKFPIwuTNj
XXDWLlmrD+iHaJpLHbayV5ODFbW1KObphkyRiZ72WMIfv78CRfgBmITJmqCPb6Rg
+yzChdJgiy5SUl8/choeYqts2zwBtD4DXFCd/SqQgcTJ5+SIlG2Okuwdei2SPfzO
cI+oq4xptXTVhy5eyapITf8MJHH6DkiX8YtK8rnPce24I/7xHN8nbRytCtZ1T9wl
gH6nU1/IgXKUBKDSKPKuOsQcnpb/J/sl8lYVf3STpIaY8PC+h420WGdJhoz99Xyf
ilSLl2fiCbYodqCmlr+FaWmZc6cSypebqRJ+iN7nbjSd+BqcB+7XVY5WTvYAO7kr
1JJ0TvetIbjMTnjxvHzmGMjqcMShBAyW63+hy4VjYB9eAZAVjSGVhy2uDpGfMmaY
/CQr9gvnP21KqzQ4pYAZ6LQ3a4wdZUKGAbwEos7nh5ZWz0o7lb2L19Q1Q8BdCZ8W
P2NkIEOk6nf1TDBHdNqhcVqB4GX+X4Xl63BWXxCcy3ZtJSO9RJBd71OLNMQVMBRt
pvz/cl+jyWf/X2g87a/BHJAQNlOw7k4+r4jCqh7oWv/ZFpLsgmbVUt6SQ6J1fizt
bhwG0P6yeG/oKfwSL2aBZEsfqFRp6tVNOvVVZop82j05AJUV1RqSGUmeJIwBl00M
RcJUW+Rh2P6xMljkmxShZz4eQFRGf3WTvpw9m/TYNl8ZauE6ZVB/B9FVohXY5Hps
QLyuCFcUBtfs5YDWFrccZa2uN+Gf7y03ryPjyZrMMk1g53iQ+NDdB/USdvwMgwFY
DgiOsbFFxmQuaUPQfE5anI5Fv7h7eIqai9lQFgSgB0CKY5YOZmOK/tVs6JXojoIH
u24NLhGP1pM4vrkCQqg230eLv9cshx/7sMor5xh+n+1LHVeyzr4xRfA5gvfPIwnb
rYSZW/kwU79rXWqExUNKfeNOoCQVkuy9J6lUepMXtH57SIjT6T/4KseF17jxp1li
ln/WT9xIXT6danWaROyvpzNO3IXHjDUOWAGyX4IlUq1S1MRf//Z3xfmhYVw7vn/H
GNTSHXBNBDAEjwQJEIaBqU20r2nOzcz/8LLIhVi/ALM9vxSIWZnoFkCGHv8MSHgl
CeDIPVpdKPjovEjhkfVmnyV5zzy9s+3tPcEWqOMfgxtPmFmXzn3MWexTYVU5XeKl
t0z7jyVv7J+fIGszB/aBgFpkFMLArvIkSf1G9vf/p+72e8TmywffCnOWiZbAZ8Ci
YK0kdgcSNmmZpzr/zovOkNZ+4N7DML7xKLbVmPuJuOe/rYAhYJ7Jx1ljfFPushyx
emOTEIpi78MiYQxImKJ2n4Ux9uoflduhsnMeirvPIW3HLyDeYqPSeLzcNFKCy/Tb
Lm7rWRjuAATXYhAsM8YPOMICQmavJ5tP/ywCR9fyfrdT1MfwBccA43nnX3dbtK4J
15JePtBLVSzFJPjA0Jmmlq7vzYqJM6wOKFDdCRzw9DlSKTqLl76fdLg2cBJxAtAA
fauHqOuj9rVwDcyzyg0iUiXsiVxz6yOLigBPSY7EmHNOl20RU6FLgh4HxDA1g0s1
MixStMqpjYKjvzqxZdkH0vJlCGWPO/93jGTVwxnZyqwZTmBHOsTSU2zqXjr+g2ip
3jV4j85XsqidUFZ42OBXmOVeNJG8umBmcbu8WnuDKHPGLZ7dZoIT3cvg2qIGSDw8
rodRU4ekYRtA/mDmiZkIGtfm0W/quLmg3x+N7HzBv/f8ta0aiURnyuTWTeGFJo6s
2rpDY8MjIeUzMEYCqQB00hVMk8ibmTEu8Nn1stSgO/w8gQT9OWbKwxGxSOZYEjng
rHNTQmzeTiPOGJOIsPc9dPgmoRg/ze1aJk0uPClAcq+CfYdVebnK1gpgozg26n9C
Jgcwd2qxpKoZQJpQoOdufV66fHo1WiKKrugWVmcbVYjYV51rBhVm8O2v1yl6v5ll
qDbyXHUt3sx+zk5ReqAfQlBWI0SMFNedNRbJKK/AK9Y64Wimi5ebC0IlQwigzs/c
6IRsdNL6Uih9+mFQhMYw6B9luqQWhmYFHtOqSxa6YH0c4bnTxA70lxcI660sIgz0
7y8LwrZfEFyLYoi6AYihlm2gMk5R+YW8g2Cvy+iqdZqfNlGaAifBWTm++w5DbLk+
612cW9pa0C0OnZHjoEgWWwuHaj6TkHoV/iorIwLpLIFMCWg3f3XYnUgt0GnkjKtF
wmCLU/px6dx1mXA3J+fUPNUMpxBw2E8ZjAs+laJVgw/sxOMdzRDNfEb+hzxayvqL
LwtOSkUyQsCRohP96XsQ4ivtyiSL1CMdtlKAizy4nNbijxbw6oHK30OCfzWNZH8D
SfHkSUwNYNfiOpkfRbL/dPalO6iA7L2d3L4HlcyynYbJO0DnTQyILaTzUKfE466i
nRU/T296Kgw41W2sjw/ez3jXyWy5nVuvKoTouu8IMackiTOf2SFslZmN7lkwcpq9
xY2QcdrY4xJAItr+ktaOE/asTLS1TT43r6jwRb/af7zhs5MXwBqdjogH+zZAqsGD
6bJyMFNZCys2JMhm7YqsCByMLOkfBS7bFn8chhA2RFT9QeZPJFXqKnvaw0I8y1ac
lBu5+/KuO8U4KkIPlrdDPw6lB8O3zTAhY3b5xOgrQgz31tBypciBBtu3RJcWfpgS
+V+/dZIP9eV+BefEzri8qpmG6O/F7YfDpmQ/kKsy2tMuaL0/m8+/O3v9V6D2EpeD
bErgEdw6px+8qJCbu/i1nIBvgp3wMERmd47Kg5KJtoknybdMO8f1VD4cuTTYyjfu
yEhuev0C0g6+Llk2Gf8psPo7SYE7nZZLr7L1pXMLPnwAgINLdYoaMJCM2O5Zq252
agjOdsfXzhwauI09fDlh4BgdSyGVHT7yGLu9HnNoCg9yK6PwOVU+NO/mFwbwBpok
VGYYWZ/Io3Rir8favIErG8LVO9KiOUQFX1VuOSvqJU4Ks0ysynclpeeS9r5hn9t6
Lt1d/rYmC8s7Pzz0R/lQxQtxbOJvwcAvYBm4Kku5Iuarb0lITnMKnXOhDu/Mk9+h
ozSP/ApH5YC9zLz4Kjd4OBqvMcZxtsqFrL66afcl35Ut9tcEXmO+JSACSKerB6l4
/yuFIOhRpWTvh0jXC5iZBrR7RiLmlUvzZQvkirlnvEknkzYLyrxd88wTCxNIgVBL
MkIA+vqDWgVhdKp4J6h88AGOGlJJ/ZklQs9NlHossEd9/+i9ve4Euw8LCE0vw6gQ
9gHWLuZrIBHEdMI2cuenc0O+NUt9+0E71t77IVfJzSP+JvYbUrQaUUHPb6yCC+7A
+1kF/PCj+O4Mmj9FTTyoDilddfwFHRFDfa1lndbWxUhQeCDA0V3dHWLiP5LPLE8A
RAhMFOa8OLQ8L4Tr1PbUP03GvrvU5gVwdjS1M/Od6AZ1lW9m+mUPAmWTwsSMJvyw
68mEfhHmepQKqnnfz0Zu7AesekO+tZPze9+SHmeglxIzt/9zjBH0j541EjEnQFka
XTaMUsyvmkdQBEClhqi95ouvkCUKAh5GHy9A5jqJ4VCxVOkHeXvs71JwYa43IpMt
SeZ/Tl06ugSnS5A6MBSq5XeiJwn1xqpdqkmX2d2gvawWzuRXM2/FK1yL7N/nQsX7
+FKj/h6S5A5FVgpb6RCSaaVLUhtrvjC4DaU7cA+VrWXbUQo8sPPVweXoqMRyF2AP
bKiU5dSJj0iAZ0MuBCqnYV9EiAfHg2wzLOy0GMh4cwicyuudbaCRZdrpTtCS3r5u
0KQui6yOICr2bkJNHdMV0i7IOKDEgie6E991cILR3w8klonN0k5PHcImn1ZqO9oe
onRnW3DSZgmtwIIKaoB3zV7LUYhlpy+EfEreVE4gxr42sPLePjD2tmFfWtszjc5g
PKYn2Xou/h/sF4e7IAuMhVf4shS9Z+BNsWSlIwPeZtWhjnMw8oG+PYmhFBr6m12R
Tn8ebR16OK29mxVqgR0mmrAgskSifoWtyMkR3L3Op8Tc8sfLNRyQide/LUlA1ltQ
yio8miUMqZUkOKIFWQ3BV0GaMAvm3l2u7akFPhhE6zv2ne8udsJFZRpLUI+XhVjX
qAAY5miLBnm1gmWDo7XMkoLPHiChXencLDlo8Wbqpv/PeZgbQoxzOsXI6MQq+wi9
yP39YIpGBu2qHWj6+SaTDApcQiiXwDVcxkVvncFjm4YiTLbda1btrLhNTBfgRy3Z
lfB93wurBDIMjJNnkeUPYNGhscXLNGbNMvyOy86BnIZ4fCUVdUDL3MmDBwQLGSZJ
if3yLYUgZ5eaAkZezagaS2vohwiczgYB6eSmoAOzIq2dH39tfdMZ+Jx5E3T71RK3
BVBxAawb+fLXXyK9lGPk2OA53wEaVIrxR83Tr10ri/SHEBMlVYpvqsA28MS8XJLE
iO74PRiiULA0W1Nzr+fa7IfwinwEbPJhuXexSz94bd/58gMo3XU3P/4GXGkzZZ+e
T2ojwnrt6cFbbZQweRAdy5c5bOjD4VRDrrXdPaMYm3PLy5WSMwMe90BrF49u08Ue
o8h2SgOyHsUQhjh4YA0PNG767JC4jGtMnYfCZEHz4NSutX/kRA45en0quBWpO7/c
l2JC1oB1fgaC3v+AkFBzKArQp9QsBfVzTjR5nqjF3mjdWHp1vc6qPjFXGrVGI0Ro
xrt0I9AJ3aplqY2H4Rq6BAqn5dr7s9dHIi69KDd+RI7lYvPzizwSVO4FG0Tch4af
gbTJGdtWcwb048rjvHvuw5+kLk/RIYY5bszvOA7PLBkEkwcpgRDb77JSaydEWXYV
bnA2oQhVOKxZYV0kQaaBDNi36x8cOU1cJWHuEYaMun8CRt6dC6IlTbz0toa/uOrh
FL6Mhsw6/45acoOEGAuKnDE1ZoS/yS3MqfEzsBvGxccXS15Sh/PSewQ5utOLgSqA
qz5HW3ezKrFjPoBV8nhAK4hkatVicT/eSInmZhaJ7g6ldHIkePV8P9SzBjIA9/X0
0/TYRpFtpu70dNccS61lqiQv3tNy7sowtQ75dZsoo4WZ2/cKpwgRg4eZVbIdtzvx
YyN02xnQqeGOyGsCsyuB7cnSzzUdol+skkRkqKs0yNS8j+8r7FcyQYZL85/8gu77
OfmouKP5TgMSH2u67cZL93Q8Y9aW6caDPsKlDsqX3dzxeE5lwkJ699T23abb60FU
ObRG0pzB1ZViV6cRafLE1Ixis1Yx2YV1mx988qd+Q4fHc1xzBt4u42mfUBrU8itF
f0NjOmHgn9OqgRPRoKSPORus0tJahFyFh1SET4EeQqHcm9zmPNiYJ98QZSw3LNs/
QfDortiXXaHuoBKI/zGEHI0RyjmYjT8GSHK09ZcV199AKoywm8/QPN/2QvX0xdbp
YJ6u6cC8TNCwPq+p/GvV5B1FTwOOgGrHw6tJu/4DYkocqRofI5YzcUXkF3YWS3jo
DRJFH7w1W3K+KKVchNjiWZoja7snCa7EkRwebCn355thSk4TyrQGGKicWi0ppXMz
zqIbTLwB3Zslj6SsBpeN1cAg7dtZhPWePMgZ+KMaYSYEmHqEUoFZD1sMm529tTEm
idKU1BAT+6Fy4rRfqSApZTzMAB3KC7eMGjndIaOTfR6Wb+9tEq6z9Ulqmu4m3fwD
4pv01bM7Z6OFEHZZgg29FlQuZmNuQMgJCto268OOYSal09aHiEFTX0o9DwKd9Q98
G9F7ypOJaU2nEbqriCIFP/yB/j1JDolms2zgTMDovR/QQiW5zIL103GykAfoqjZM
QRDZvYAbe7OwOTIqJuoy0DHuQfX5XbL38clpnY9N97wNVWyTmZ1EQ1vzQj+9284u
RVCnjKAnc9U+BvlHSPivcKEKUn6qSOKd5Gn9OT0RNyXMeYzD3MEKcBia66UmGIYG
ZcNcJrt5UgEnNt3laROOeYhjy2R3xS+AT43K15qc8t+fpVhqvIF20FDnUOGT/R6b
P7nkI1VSOLbAgXgNy4jloyQnOX2y8Fd1ksx4aXRxEqQlQLkWEd9VL7jKpdkh+ysf
ZnsxmVMYUSoZ8m7o2KCbqlIvgsgkA+rYITeullzp6doD/GFOTjXelZGePk4OA62B
gdDTooxFOd7BWMTFxutPFDYjcmrA07KxRqG3HnGXgh0toMfVmBCzrk67bpqkNiCm
Oeqi0nvwpY6pnyM3IFGyFlstRGLGu6LOiVbBjjFfchMew1TCiZkf46nlW6eQrMOM
At+aR+xAs5mH5TWm3uzqgcNSzoOB3iQ3TjKC0QNZLr5to3+aeUzgTUiNTrrD3ZW9
clF4r2J3Ct1ndyyICST2WBn+S3TTf7FNxfSGBq96Q92XTkij4jp9kAhb9NyaJP8K
5NZLkrw5a47AQkXNHxbG9Dojh4c3UN1ga/mFttcBscfIVkFpUwexB/W8CP3NcB16
drNi9rms8T2p3hh89rYMgOiKY2CfwYl8lthVMlIHRoommlkCLKUKHM4J3Gshve9u
ytPaADQS1/Wo6NDomLrj+Kjgtikr2LU+zDmr2Y+k1ufb/3Mi66XTL6are4T0M1VQ
4glfkx+tUU85yEUiACx84KnyOTlPXL/dK/twkMITwMGw+gbbb20Av9vLR3iMPex5
u2q/gK1y4vtSxycM/SV/sZMaE/pGpXRTqhesz75swI3BeoM1/v+hGvda5hKqWq1m
OleS/lt8A4m39ThSmVniCsGJ9bu+cUVsQoZqyvEWIiiIeXI/1jfaedhAwel8KDKc
0VAeuEipNxXzxkrQ0fu4dViKyITa9+of45g5mcDnXPMv1IjvU0abX9f42g2wzfhE
EEMVSm2oWxqEuzradKGyi8+AnkWvjTs+ASaPxpHZo9SxKhJ+XpCT2++jJmppmhsj
dAgG+JUpQTOu0ZyCCgt2bXNzxSVsfPI3aYF2Mi3oMc0YsOpvMIJk1DrcFnvyth8f
a0yPEri/K+FWFGFdokE9fO/LnJ/JypC906AjZYiaXZ84YNNbDe4eKzsS4kY82cOr
VqbHxLxXguPMU6CirGlieAW+pLsN35+oqPywM2yUdl6HWJ5vIwtBCGOEbF1NP7Yu
fchZmuPhzp9pvJ6p2YEUpS+h6uJh8g/kEv9mun+yJ0sTpPEm2HSJZfrfSqNqj+BB
pKqnXZMfq97opY0wJgOnbz6Zdhx40l7xC0VVoCNLM/dCnyXIVRql29eR6l2ngEeV
VIxmKp7H4AR7qKzKRhWEqutxK2LvQlVBrzUBuigV84AHzY00VPxVrt39AetZWY9u
bSWl1uywdenpnQX3eIszb3aeqzwDCH1jVY9moSzgidXy27jU27jqkz/gxLwV42e0
IvIRTa2yRUr6bcFaIttbYznrD28fT9VShbgasUm9BGmOTV0zh5XKSmfW9SJHzwk7
Sg3ZNQW4bdM1JOeInk/Kiq5BWEvBHH5KMd/24o25Y1RSJV4Ep216qDZkBsIRvCHj
ryYqLdR34TQnuR6Khjq9gvx4qJs3SCpqQcVKmwbK2WnTDEAS3qkCcqUFvVz+I9Ot
17Th4zuD1h64Jge7HEtfHaIbTmJFDlNW6ZxPB1BLU5goxgsMJ2/NVj5L4kxQmz6V
xrsGcec0pD2ASmVSPPLTEHvmstMGIKR4KX08k/oSSfMvs/kW7HCnRN7SlBcBciNw
qm3JT1FGpsomG06UxH8Ewn4lPfCzumROfcmXnv8C9c2iXBh1JIuy7+pEHZEQKLbC
A8pVyCUzgAaaaW8gRBCwfdWz91Gd3M93/LqVHfp5bN5X2waWHe8vdjiwAhB1A4GY
RM7oDcaSLlOujLcUJzfUh/Zu3XTKJhs+CSPubdWiM4MyZo16mZ2yj+tVxv9PVa2C
xoutYByeDzNBwwhOxgsafkyEhWrtk4cTIU7/A62qcpioevZ6lc1uqgPz596LlEJb
UPvbB5XqhSDgiTG9H9FGTVw1CeGmbeWHYaFzcolJmh8rp5XqIycHKQy8dwjCKRBz
vZJPlovP2Xxlzy7HZ/qwF9Pl666g9qBADQCaMVzXZQmLye353ak+00iHOgAv5pV1
kfndaa9m82JpdBjSe6jbXfn0sJMy4Mtsag0e+0SOopiiswRLg6xDlg+IMKFs1BmK
lvyGMWLiw0LHto1b3cbm9OPzjwEm7ueoPxz6G5jFkxSCxoDFaBr7vqz6MJ7nnA4K
Q941qwhNbtrD4KCJtJa1xOR95iQEoqMGiQh+KNAYwFJokGmpJn8GJ02tnEHuy2GR
NBGv+XixVJxB666meFVhy9AWMLkWQTJy3HQM8tkMm2vgnNN4BMH9oF/MovB5S/nL
u/KSHMZK4S2D4dH81UP6a0gUyizAJYTMk4W5O7aR8e4oV+PfOOjXJ8SqetMAmM7m
Np2ayoIKzEq2titIBMqnEZL2F7z5MudBF2biPedrA8TVkYNr8y1f5b39vrlCGFIb
cRDdogBDeC2F4vUZG3rKcrxiyR3yyVi7J7whnBjCAtQ6E44uxEK6XF08GBF2IWOX
18bwzDyNIntlMgUtwM8SCZr38TbUPqp3GrJYiCm1gw5bxD0xhe0jnm4BINDnCIBt
uiNtye6/MWlWhsJLfCMpAxAce1qSIrd+D5uK6pamxA+uowl7TpPv5/v2uQcg3o5G
eUn3jaZqI0TkvP9HAyFKEl/9pXDsBsdpClqr/mzoXjYEYHxxRkLsjkZGqKGAF6/P
mGF3oYwnNnmdbO3P5HPhaKCr0pGOfPhEZ2j/YEIR6MEBQuxaGyRCDeeVWIvtSsoN
XI0OlU9Y/X2NBLxjelo8H/BFDU8i/iukh0gHYQMyfUD2x5qLANMJvHWf4uWpOo9S
cNyZOpxgjiq0eLnHuD4EtnMANKzqMun+Lge9fIRgKhZOXqFLo5mAp83G8a2QQtpK
5SraCkl55za63N0xRhs9hWSo/VZeNpaFdba7R5HP6bngN9+DXOTWDMt3uanAdN2D
L1OQEnwUXO1BCp5iu0X/nmXV6Ab3C+SGz6fa796pcigL5Sn/otr0liWOuNZjkCLa
++SNwdkE3tLjHiRRqQG68ojrqm+LkKswZgpACqZ39gllIpl5AJR851ZYPW4SiEoZ
rp7oMS74sMhaxJwlv/B7lzEbxYixKXwwBBPMBXIoVp2S6S9S430S78xG2Uvt31og
EWsGD1HVYpccsDexrVL1TshTKve+h90Mk9AMf+a6FjIsRs+LI2t8Hdb05EkHr8qJ
gLXNBX8TxgfJyLZ0vmPcZtvypCaLLuVGjTn3mPzShwfH8m/Zf9F2h+WPcQnGCerx
A+l7d/R6pI418uHXl3Sga9I9lzGRnHsyjFrLAwcLR67zcZAw6jfpI+Kekt1Td1Zl
xhxdK8RA3LvKekZNOoLqZaCVNdUBemV6hsmO8LwitzAj7ZoK1/Cneo+fY83ghDpl
J3lGuzGpRgRjTBePj86dUwaxnGxs5yF+y09z0ygwEcJf09YXjjD6NwVHsONf0ohU
NhICTyvupxImV8ZDZYBMmPuR8OKGsuXs7IPUjyMJ4J4AU/QvSOj5Erv037j63Sc4
+69F3G9rrV8xg8VU472y8kfOAbqtqCHrsiMAdSfEmFXfpvjz2GH6DIjcDHEvq+DW
nn1fStxbgT0KpW5UxiLtE2GiPhbAaap6T2Wob+cuOnMCc85PYgMZTqj0iEOnSlIb
CX8ISVGzneEaaZiNWfBfNMIK6bBZFTy4383IJsRyxCSDNtfkpjhAqn929vG2gi7T
NYqCLVWxKSJP5qwT2wlUkDooOKOQC2QfFIwJB1s/W4fh99IBNalb9KrZHZTXZJ5P
151ooAJZkA0yQcqwjdMh1aODdWICWjb7jOhgChbflEThQ7LwwjSQd69yqpeZDH79
Fm9o4Nq9uU5R5zUhGbxyD4SwmdDsQJWhTcrkj90DUgxRQgycPemqSRm8GjM/p+ns
bX+podeBLHMpugdUyU1HwECXIoXm2LKoYb9unxY8XVwTylhy6rF1KlX0aY8ndvRl
MKwlPoU8jm3ECmF0htazaB1tj3Cd0+jHkEV5+xwk4JEjnnOD/v5y4la4X4oS+3U9
cCQuOIWGNtDnoEUA7OXFoEXpSo8iiaDgJM2gt5MAnBJaqt53yajb/jkISglXSCNi
nFOn8dq2smKvf9nYugMqulJNQyYcg4BdQN+xiILnYZuyQ/Nq0UTM+r0ehOJpAQEQ
Db1J64se8RAvGF3Q6TXJsMj7X8u7bDw54G7zHTPuMBs9VCph+31gGVLv6phzEj/N
FsBFZIoNw2uBrc/K8msfIvWZn13gqTDCuzmvFt1uU/IhmYWtdFqgHNcPuXTKzAkM
qogsxGrEsN0wWjpKyimuc5UpiU80xTti0QJKBCEQa39oBFiaS4vmy6S/BPP1hbH3
y4yKVfwesEobhJKD8JetD0ZiByEoCxr0M3NhOV2vt3lsCgvOcaL8IGoWgYOUWFKj
zlXMlipAQ8MH9AMvto0mhOSIt1DysrgpoBZsdUhmCm1S3BhQo8pQ8amLsHAOBXRP
Q1F8fjgncHEfe2BR6YGbjAywePakD7Et47s7+S0gcRfS3Q7Xyx+pLUhIz8CORKKp
y1PtzaQZU5kYeq5YG2KwE5XruVybF+GtDudYY4lmbYg0IcJe04+bjZ73Cilsofo3
j7QpC5FGfryeOkbU1di2y+DkClZ7Xgpx79kx6wvB8cj+D9AMnJnZeeZwPzrRfOLE
7m1OsmYyAH5YFRqy2qe3wTFrQgkC80MN5GiJDDWDKmcuYs9xDzt9avr3qn2f/65G
kQw5lU6xN1aW6WcvUXR/fgwlcAqkLNwPMVYDSklnSJgtARty2ZTsIuKwcA3IvzrS
7q0dCPIXAFQ9IbySz6ctb3u7yn6fJ1l4Ay0CGLqcMbnzMBZLtOauPtc76f0UeqW+
YcwoTnhIuhri0thafUf4W4HB0N02gdDrPjXHckrCYn3e5X3clP62zkU1eTjOnfxW
gQXtLttzwyB2VeJtdkVTKDMmk2WkNFbQzmFtkL8w1tfFsywK1EiKyIjzeTuWr4TK
v4/RM71y6Yna8j1CW2Xf+XMjbTMSZ6xWdXq/YpRFQ3yCUS3ODgCbPo5lAqq9AcDX
qx3wYkH4xH0AAAasB3SQGP4jYkax7LtLPSdvtKXb94adPn1EPR9nP8/rL8jVcXts
kYRQ8gAKUv9wuJY36socjbwU0EnQDmv5pA77cUmqjIqqFdersu5zVse/ocArBlPc
ggE4UAtLDEp8dBxYecy5zg9YgU13Dx/nS5l3Fbj9V+Ul7VoEzkIJs3b0YQyMbFxI
FsFeWrtvxkbAq6ACt4p9/gkMP2ZDTwcjxj/qLXGadunBU48S3wgqCpN4WfPQZ5mE
ueACcP/WFC1wzqEQdRYXEIBQXkbidSPD30FT5EG5cEkJRZCzaaysCg2xyRvQiF56
MTgLWM8T4NQvWElrz+8E1+PX7/zRyFaQjiCCEF9Lc23qVFY+5TrUGEE0EPZEDXcT
IwBHKrB9pDz/KOhJQZLo/g4P/WmkQ3sSt89Fq1cIQxNONgi3adivp9ASntjHaQK6
i9sYY6QQPEQhKnADgVuTKgwxrtzcg265GeXvgB8oShH/IzDmywxEeoFOy0rreiy/
ltovZovfY7bLko86eIvp28jN9EkfYKnIeC0VOZJJFZtK6+PM6h4eEJcjWLHqnifI
okGCteLjLgFLpPD+vhu5BE2VjIGIh624+TlVfMqqfJnuzU1VgP5sUemEcxdy+6LN
fFvzXLD6mhXSebeBnX/o2lR4zsnZwUT15t7W4S+0VVVhBheeEYW0X4vsml5jhd9/
3a0SEJ/bsIcMWLGWDTwqaPAZi5kUX0t8W8ax2u+FHagFOoERY5vl1Rb2wLSvEsgs
lJGrHpUH53ZVRpKJl3hyvnttNHiyrh6dnmx+gpDjOypm7WlTjUtLUBpdInhxJ9Th
y7rQ/dcmmyLFAeXM6jx2ItuX25qkUHzVVSg3h8318MOf4WtKOL/uwDcF+dePAeai
ewO4qfC/yFjZJAFdxwdIzlXL/EJ+1odz58GwgMY/uUX6SerB4FO3D/4M9pxYnexv
vIQvrb4ff/EXp4bz/63YRGqfal8VshbHrxUCd/Fk6FZDrKJhL06w555Yas094d3r
o4mIKX63pIWVt+8gBbaYW/V47kRYmwT7yVYeQOx8Q7dRrxFhM264320HoXfnI4If
2ysR+17UC7B2kquDlAcIcYh1VToPvUKw1vAvlb8hYdG78JyuqtjVoavb3W6Z5j+I
iXHFWEOXHPga5hXd/ahtwC9Mnx5TsiIwWHgk6EsBiLafnfmzG3hGp7hmv/e52EUW
E1wK2Cx3oRV6tTZCBZJk/gu9N4D8uKS5XbUdGZJ+Ms7T2xNN/s1Q7ZWgu2qO6aF5
KMsFiKwJvuIX/EIFgyp1DOfjYWSjZhmsCuhyRi8/0l6NoYxFeWZYaYuUcGLd1j58
7VTQJkzSyEajy5GYFiZ0VxxyhV9vyAKi3/VZLpVmVxYAp2zdP+TJLyyc8E3/dCRE
fE7AyeNPMFl/gkRWWfXODinohZQVr2hjNIGtsl9PI+mCoZymu5mTOTFBxCXKY6qm
69pLKOYxdsP+C1NE7fW4ZrUTYK4ieavg+ghm9UzSRt39OXMD8h05hz98DFnSy5MC
zNwcYFiWADqTILEwEp+Ki4bwnrM/tZjhYqzn4IIjLBbzAupCM68RBDcp63dQEKY3
dDsFY9KdksPuH+areTugN8rcPYuQbvNUX5JdZ9RF9Tkqed3gyLW0FsEaXAtVF+EE
EBRmFzvBogxMI5Q3h2/iWZ3MX4SEHb2KXqp4hNVWFL1TYXZ6VrNODFlPA/Jy3kf/
xn0yYz9tG7CCmRjanvSI/uMI23XGo4QIGl7g1f+pRUQK7pBuIdSN0IXbzyqkgdWs
Qo9XLzUYSQlO1IqG3P0/IxL0p3mhaf2nTJTvsCKLi090MQ+uDmu04g00HaVWRsGL
/cPBziZ6/6t8zmnBErX8pVP8CIeJo33GMD9mRAkKOIcVwLX81VXQ7ZyiKYWl6FPd
amekKbMAGAprM1zlfDdFBtf025n/j+mtRzA2EzuX2oRaKzteD1riBTbLD/i68aex
zySnhUPiXSKVt+bQ/6pqLKuFqG6UIgvRlY1CcVfrACKzx9fL1Ep+a1iYq44Y0UPg
B8EyGHHF5mrpz2TZXxwUWZeOohAwTBgKe+Qv/IK6Jn6OBwCnp0YRml5V9Ls92Zj+
6sGAKBYnGe9Wu9u+YnCXnYXm/sH5Bh5dJsDi0ScW9ZEFAzz4GPQ+g7sMaS+FnQjp
9rBtRkNHj3MXhDvSl5WYYDI1IT6T/jS/9m5ZKjsUGxWt/mGghNZAd6d3XCIMVTxt
uCcPn2mQ/bnYqm4QGn2ba860gh78PYzAHdQZCMmVyYbi5Bs5GaYpRvkKJZ1x5oDj
iJE6AyEIC6YJnL7v+w9MTL7Eo3EHE2eAq+YBCyctxYDIm8WcSkV0mYzyvT0yM/5r
2YWfg+T05UyEzv6KaHRZFkt0QM4zvGGPzb3GkO/KyRSjqs3tDi5CEliU8Csokn++
YTcPEp3sznlexL+czFleNSOFHncETpHhHbo5IQgKryPYfcerh9ECQPm+PFm91WEl
K0VUut8lDRYhG2/IdEyrfAeF8fqX+hR4JfQcTjY4YXmsMi/tXGtiNT19m5HewEyt
HrllRXpLdSyvu30AgTfluzOtRflkzLamaEGm2NUkmg1kgVfQ/Hah4pkx37wT+kEo
wu6TfeClTisKZy60QqcR15M1iokZCEfe1btlX9ZJdfAkZTPRsDmia2LEbt+kSjlk
9F4Ka1J4oYchJdAHYh9lG6W3stKtI39NX4FE6LkYcAGfB3PVhcLhOav2Dweg6Mqw
nEUCtT5yByU07UoDTnBNeKV8L2uVA0srQOn1L/77KLRvB4Y5GDd5HEi7rD6B9yDA
Pn3ZzeKp4/YTTPTyBL7qLsAq4NG7CwDOwmyfiJ5Y04c6U1h8XzFtchqZveXh5oCS
6OLXcyi/exbQyZzk5AezmMuwcjqDZxUDZ0Cf94X0rfOVYg3kq4v1WwlgVqbAATZ2
8JqnNovozN13vLp56uBrhsK2oO2H+E7D8SnAoIS6er4pKrAqih65ob8PLY++0rrw
COoQs0f70Sw9na+S/JEqKOXbE1NUPT06rSe/OVS46ZDbFP1gRCndakDcpVtla0Jx
GiKf+3+bLEDU/bYZd34n+Q3YWbzTs1vmvCDZ90cnnGNA6RI5roUN3dUs4e9Pu3PD
1I5y0aWVlDcSTNYB5ryfiGiyUng3eo5hfygoONw43B4gJmYYTkjGXKI2GuuUyIco
KHJPEMa65St5ySvrPI+2s86eSukTHwG/LrbRm21vKtdcsGOPDKu54TrUl7HEBtZX
p/34JlNw5jy9HCYMLsngv6dZMcxQ+NHovzVn2Q4B2UIbCErRdSlMIwI3nqYIXRQS
QX02tD0H48qBG59s4eDepyKTX/F8THPnQBTewm0zoDCXMRyT5oenPO2h/gkCnpCq
rwIp2VvyaRX9gu+3lmsHElHMfis/qRRGdVqv5Du1Gt1zfBUYFd6ACGt9Jki8WlPt
mzCaDr7CXDuv9d4Qe9dBbrc1Ws+54qZVDUzNWeFDHtwVJYLk2TZqFE2hQPozhzpi
jLKqUAoWy9gxf2CEib2HcUUV/vPoIkUK0121ZodMjr17xsAapVmSi0mVP75ya7VD
eZA89V20gfZANLlgmOTreVPsgy/TP1XKMD/gDSIopjzDs2xroLEa4V9PXwgeXDgc
xX/4fqCN309fErWN1w0Au5AcGLwoOEb35AMqXbpfCRi4nbPoPuGAT6OKdnN2/+65
O/Vkb+5Y3q9Tx+jBBt9fwOcz8JE6nyGoZOxn6CnKt1J6HO1B9GLSiya0uTKms6NL
Pst2DZWq9et5sz+9yYrKPZ/ecmF0RIYI+slTlR+aiMC+44/vTTnDzZbex1RfRY/S
RXvT9rvdvgpDbzVNhDu+IGaURlwP6+MEc4CSXhgix370HXnnOSo8vTps6tyYVlJl
a2TbqwPAGrbf4eXDvqGYJuLIqTwPnkSB7xzMEXhTBs/ix3mZW0M+Zf/wLSUgcePe
b6712jtRY3iGXmfik0V43ziDhvv/Bs9xlZJIe+dROZi3Ud3ENbuGHC/1Pkep0Y74
ud5lal7SCvmZ/XGkfYjs7g3iqooqLHQCFTXX+o1Lm20VpFZdCJRx8/zyycF3w6fV
vPwixfBcP35vysRbSlJEhWsw/Li1hf9mp/WRy12HeVhIQTceEMdSJaYWnnO8aiGb
Fq5ttSgailsi2eoQVthXoYbXCf3YE55AlEx/CZD0eOCOE0VNxKhCHp6tOZlOJpdv
n3oy1QXV8bDacDnMN/mTkE9Zsfas/mdKmlo4SjG93UdKusZ1xlVk2NsBYo22EoxM
A+cEY3MMSIekuckZi9bneUOUea9UtasG91RCy4tzodExkInuAkAnLL3NuDlLr1uq
XhFVBEWNFyMPrBsJXMzEkDcaXBk5LaXx4SZYqEW4eR1O0Jqx3kFMhgPiqQYAd3+Q
3aZLF3vGK+XFeeMwqJsY213j/0NuY0bymKlF3nqLbtLJ9iCFCHGCyrVNs82q73q+
Ts4Ko4/p7QZ6N9l6jq4J3b/IPcdz13IBDJNBnfS61Dqi2VnDTSzzTgAXBbnBm2W9
cO/LZ9dMPkbH9g2ua0kmHqv/AYjsDNMs65gDdaDe7KPSagQVpsDtCmcz4TnWGwbv
RPsaSa1zlKF9t94gry8nBA0zUGh5/5uDP0YvKPs+ObZFghBRvHZfBMRFEl4Zdn1F
a8TwO+D9XemfJE/NZo+nMkCpqgHo5LugdjOccTJQ13II3IMhVIuYe4857hQAtPSZ
VB8jSmIbBZzBiYSmOqEfGJ4HgETZwDbPk/CyLf+C/Y1pSKGYpF+HGrxXhqYAOoOy
o7P2i8gK7rQPKoDKYPcm8gcDq6WaKBkqeVRJ6x0/DVzYQEDH4o8SNfzo6Ko+bqiv
2oK8e/7ANwxoOzjrwIfgsjtvQ2VjymhmgSJHLoXH7n9g3nvjKCWEZcQORNMs0B7v
/7Zg3/XMIKY0Ec045C6WrYxw6LzlJ+/LCZUIcteKQv0O6H0929kTd/NElPjdQBrG
IdVjjUEemOaSs9ViX2LdISavWk+Yjv61S8+aKSMhjj1C00gmBjJF+54v1hK57yyF
IXmDYlEjKqc1JaajcU11eaz74bXgWUyj9TiNvxnHJm8uSv3i2exqP++pmZ52gAcU
g4DYWG5KW/3E3N0Q9Z11+94xZ4ZssKnyE3bNlkk5G/MTCXdlbvUQE9IxQS9EKXrj
F+F0Ch6ZMI9ugd0fGR8KzJFuzrGhydFYWasiTjwjrM/ZwvnEnbrqe+FJiTNHVPZr
qRGRApVZSKRFJXjcLaKCH8hQ6SNJjX0dyRV6EESMfO2bWUjPsoXFq2c0tgF9YQOD
muUrvbvDRoHgTSa72zAdJ12fqco6hvFArK5h6D1TE7ctcyklKUYRj3h/Hi7YDe/C
ARMamK9O9zAdhCTT+Nwt1lKYwHK7iF9Q2flxPSlQuZeL7qYNzjPdM6xj7KhT/rOW
Z4GD8J7LDKRp7s2leIMCLurOFzfF3rnQLKg47fHKoCzNgrYNGJS1De5ZLK0hOVGl
n3gSovf6D6DyipEdinDUlZ+ZuRTNZEl4/yrnQlfk7dxswdvjEp+ZMpof5xODfB8N
nwNqkry0srS8dzsOflRc5MTn6zilwUGJ/JeZmQP9DWEhXpSyo6TPo+yiuI1k/Llx
VSYzsnIjr34sggDbizOc2umbyD+UlNMQ8E4WhEvTis3ZSQUuTN/uxCALDVT9AYDQ
+PmwmJbt694d4+S0uNqoh+JXrOlWOwzooTcHUelK9o3hhpeIV+9v+8mgbpMw/SrE
p0aSoCjl7FOy5k7bY4KVq0tkSAR8zi+PZopHausV5oooRMerFviOzJBbv7XORHSB
MS4MgWut1tUAQ1qv4EfgaqtaYOL/m0TaPPeLkrMRpxJZCz78quercgqT+X0Spxek
7ohtc6HCHCc1pfSJnq0FQnVEcKFNLUh/leHijZYwQ1XbWVhDXzmYyYrxs3jMMUKh
sArpFZgCmJQqJsUc/VUXZWbjk2KTyYDrwLlUsrMQj5WMq9TiQ+G7sNOy3Zaeg++f
EmxCuHf/8H2l/Lrlc+R1XuJKeLr2kAvRSccrqPs7H9vWpGOYLTe1RBSaMBTb2GE5
mng5ZuAOAMDBmvbSUFWcs9Gqg+VUMRU/vAaMciPg13wWjJGJUP0Qskl+F04gDYSn
unofQu8y+z6dgRkfuNluhFtGofHXo4eapz2GwpbEy8RETZOdkwwfIL822YFQSnXY
07MtG0LHry1vgXbUYbVYa8GVO8pd8AGt77wFM/YlMT0P4UrGcdJT2bTCUhRgtk+n
4UecPS2QzHhuDjYa6uP1BJO0FSmirVxQ9H4qRv5KIDr9+7gKO1WLgKaQnnD3U62V
3GQi8N+d2RYY05PsggfINKEQjrF1u08UuaM3DA0ZdD6ZL84U0eHRwWeJWoy4x2NS
B9/PJBcKCcU7bJYwgj+JyGcedMDszsvRoLEpWc0to+c0B52gE9F8eE+kShYsJGsO
gCrxhuEWkG9DqdoVd/cjxFnSE/meCxonJw9CfjeEA/PtwzinMFFpo+dFASrZmJSR
SE35zu7rC8qna42wpnnZKbMlkBZBE9AXxojEHGw8nv70OExA7ka/zIYh9/r5OvaF
cC3dCkgq42CZoD+0s/DTJNmU0wWHhUTXYLDPUo/qfo1KrPMs1VrcHz3XyUHP5B2p
sMSL2DhbiNkkdD+93i54tcHBC/8b9Im4825f9iacwS8qAvgo2QGtRBBoK8tt8sfB
AEwiRd7KzmtUWWwebUAcIbEFR1MMpEU5goSCpHn5juHeL5Fs43FQ4BIyZhFTxezp
EfUCJMzuJX2aFBG91QTtQVwvIEBB/0vKwcT5nsGWBpjeZBkJLA7VY0No/cUpsmY6
i0TqoKur+9BIJBL88Rc+dwINgRCH99QO7sN22by90L8x99smE/af1EaaHZk8K+Px
hBmhlykylnUIhxpFxTZPYbkXX2R7z9b2eIXqOpt3KxV2EJdSar874ZGZbAUeBRQ1
GEsP0BX5efuapDeCHZuRUpeX0ngkJ5U+OMSwUqlkau08FB5Y6wIVV8C7UoE/ropN
IPaeVkTOgz6PJ8f1X4uwLO2CmvOP2vOtT1iu5z9KSCc7VDOch5I+LGyDeHUMhrfo
3XBxvVW5XQFDV6ewDClV2PABIE4pWNFyLyeW/02vZuxhgmVDkym80LfrUvemtBtS
+UVwOQBMshoJO+kbZ8nY59LkZA85+EXBSlZQCt0w8Ns4dO+NTPR9nHA/UTlgRdsg
XGVmAAmgW9u60jFL1YrAauh81xjr2QwkDoqQt+Hi9jIZQBZ96twQZ2bRhKqkGKKK
xdZCuCegPJzE5coP8FxQUSAYwprBgKJKbZY003ZnDlSQFicaHbMGM5kGzKEr2vrU
UIM8whVmYpVyfXl6Wut7R3I870EPQ+YHrPFR/SyFDBfgQPGonZnKSVZXvHjy39h+
6J59Og+4M/b2cazVMZ00wYqsebRvLbjt6oJ2XBa8YIYx1YxztR56zTrQkNEc8ZIi
BFet+Qh0V1rBOufZbRRh7NMWyiMzmmFCPZjivfTMkhL928xPHERrgA3uYmG8iD32
IkUPFJHADKJQGWoqdppV1V3uoFllUa6RrooqqH0xhzxfRuFg2KVBB/C1vD9tfryJ
roNUpvGRten1Q7k1+E2qT6hNUBdstBVSwZXJZV2AAZUapAEFOevDonj6gCrT3xxG
60r1q8EvvLlVslPgseBqE9b7pf8cQZjQotXyTdHd3MpgSuafF2Uc9pCom7KDykOq
YgsgWF8eqROKnxiklxRU3XSlziOdwEmed9xLjPIfL60b8Pcv+Ke6FBLseR1BQJMM
1O/ah9198bExM72eafGUNkI+DOTlzt7WUR73KrbuwHFQbjX2VT8aWuvTwpyQQBc8
99o8zU4ISXCZVShfkPXCRsR8aiyGHLe2thUXspTmiZnkEkgTgUHwQ3YSBneZPnGW
x2wtbKB2XGd5OFaM3JzMNByVvCB+BNtjvL8C85HRMAPaGoZV7jHK6++DZV/ZwnJo
D5Nvp268I+xAY+4KJbWToLe27AywR+nZghto0Vp3fXjE6kP1p8UrNAdZaWm4lsLY
EA3YTpiUzWAvJlf/JgWTk/Lsdwhg6SzVhUbQ4+IvrnlL6OLIlVN38a+XM972/gmJ
Bls54mijyp/Gw1OFFUdiIPaMT7K8EsYaAn5XSAbWXeJ7CurHUoHRIa9Ew3mSJPuW
k1dTK9y+gP/iCafY55Xi1OJ0/cbmygTp0iNxAoKhdchMsWSLK1QeSMyrqb+XLrJT
6UR2zPBybfOx5rjxYwDA5WO5srC6uTcbMBODbM9ghwwQFSK6AxC47XhTcBlbKVdl
5VAMwEF0DLlAlUByItam/CZ0oX+urxAYbXRUkKonNZKatMySDAkZixoul7PA9tJW
14ShdYd+K20fGECf0niHEC+kdudr2js7rAMo+hs7hqFd2KsX5l7VwJnYJFPMsJ2b
JNY5J9goN/8u6yACA2GYz3tE866SijWmh5FKDw6aJpZAn2PuyUZ3taLBjy6efdlq
3BmIhCZtQlUGLkyb8AotaphgfzCjdh/8Sv7bmcwqZM7rH46Ahk+bvRuFHA1SeJ6V
qhBWWRYFNMFE3bCj8RICo+RCoy+TJBqZUJDDu+ZJc15ycizqXRzqiK3y8vae6y2A
3ZQV68gxso0ZUDnwQk7GJWQzMh5CfLO70aj4pytK9WTzM9OYzjwosHZwJlPF48TF
yGFY96bzcir+9/9aLMBaehVTD6BU1RMp+3l9JN8SYksBTvywNrEPkPeVeBsIPNUN
WWsWY4/PmbSlEkBY73VyGZ5gwJcjxPBwqpOPgRSFHYDrRCuP2XN65pS8gmDbmuNR
J64KcTeFNz0dSryB3+XLEAyKh56PrELaWxcmONSHVkcJIAV1RxdHvtXtKQ3o/GyF
HEc6TijOSl3gmyuITr8DNeHq3y73tBtZXsnnHJmQdhJfjqh3TLx7wIwvhdP4w7Tt
7MFCmvXLk+lzmUqScQ5JB0a+bRd47DQmq0uvq5a0a9JJNLKsoljD3ZvxYQpIQeMG
/OCQ7DCZoOGw4IsLv5FW2bxDlk+Qcm1MFopi9+4lyCx05WdvaUDau3hJdvJJQ4cs
4K3HxvryKoFhWmr3yEGhglI/w3taBfp5KbKQzx/zcktFlx903aCS1Gl5xyDtGqaS
54qn+gwGlX4QQudXOKrGEVDHvajB7c9VOnNhXhCbb5rSb3NaK6eObFX8LLRvj2cR
TeoI4ysxYOrzd2aRo/n85VL+5b9ciovoiS1KlFqqigBS6iDWavBT6odSvf1hw0x4
pz2ejtC4/4A3rlTPWJsRh88wiZKTOsjIaVDmjqp/nOBx7/ppfX8uMCAC/NTvSxNl
ba1oUVH9/C9YdEwwFILoKhgn3f4mQzvTqPH/dHPkLi19ZKS254EN+pSoOX48YxGF
rHfKkD0E5ihzX9BVRLj+wmRxlhWr88uvGBzf96PPsakkwqIDXiGb4YiQziyBlmSq
B95hjPlzHNhD4yx5/DfC5AhF1uuabPmLFYxVrkwLDUYxAfP5TA4Ws2RPfLcLSd5N
ZT8oOvB8RSdh8CdG7no79fDHvY9iCL6pQSkFP8rtx18gt7F/X2rUN7VFHcEExFq1
DEIRsadgo9maSc+SOtAG6Bp7RZmCxsKbxDrg1b6X2O1jo4fWV7ltXQp23XDQa+kn
tqut2cfBBFMQnH92hnxsbS9jfRYtJZ0W3yifm1k4nJME6hVt81Mfm/yiVNs67hvU
XdmoyKkpXvWZEwC1mlX3c/h/z+BXka7OXbIhOXUPOA2Fe7+WF8eYURYm75Z1rDPd
NV6ybQnUU1UllBTXTyMrn4v4eGS48jT7q7PuuPRodVzWoNvwSbE+N3EKtdEnDg2x
yVm3b5U8P5neTw5b2HcsgP4Tn/3yQnOlAhgfHkcNPa2g/d98ZRiTE3lTGZPK5wTy
/1ek4x9r1gGSiIN9CwIJXsV/MCAqnhW1dYQ494aUrhPTyNsm0oXlyvCbKNHBkzhH
CBMFW9mtIA4Lvo7n5E2I1WfXTJ8Kiq79HVb/juFvvW2FTiiMCFwrGRfLTtmZOne9
HG+nuxO5JbbNTt8okiOE+HZsI3y/6KCuERte656ir776rJjvfZuPSHXdqeHZSGP4
jUi1yE+DFsH68kHNpnveLJUbGXcG6lSFeuLq4mb/soqXVXMkCpYorFZXmHxCSWDi
0i2kEooK94QJ6VN8f+YAfL1m62cmhR95Yu/2m5YHexJWQI19TT3KLZPcdiagGMgS
auePi9Ai/rhzt1eGRF7JazFLv/xcWXc8vUD9zFtpoEVOSWkJ/fbuV0iOfIQZzZap
INK6P8TVj3MXdvU5mlp4mpJ2ZHynRPj/39kmYduPOdu3elVge1qQ1VK4mKaRmXMo
ym9KQ3aH92Vj7k55B/CLTHR1kka/N8An+3ka+o3Pv9jrHPsmdumWMKwULXIW25pz
EXtZfGOadkyWip4TkNGVy2akZFjdxTXxrQTLK78imUl3MUbMZB+h2VKZPaSsO+de
iSaEzpXhIxvUiPwFdvajpKBb5++z5AymeqKVJDwCSwf8qZ2HOwo6MTUVLEON3Hdw
0lVtnQp7xUyJ+5BivqKGPgRBCOqts++2c+ubc4Ki6SAPo+wyYG7teHNMitiSROFB
icTxjec+Key/gEY+12y71cNTy7KD9sAsetOm6H9MN5RPEmhom2R8cuWyzagfMQcv
+jqiDvyvxilfXbPeBNphjbOGrjNx2IZ+s1AZ3IADsc+b/0epLbELbNfbXAICJzrV
aIfFT4nJlTHpCL8BkBxSD2q5i6PDj95+Hgr/M8r//r6IBoBikEztZbd1bbkGecrS
Xr32zDHSEcooCBPXej5mjH2Q/qVp/T7/w24l3Tnm0gTXC052+2cpw3RwPrGZ+jWc
GHsrd7QUM7hYLVujUHYtoHhpLr51W0UN9urhsqw+dd1paQ1yMjDwcjN96rR3A9Tb
u2GZLY9H7ALqH85ppUqvHdAVFNQKEHNVD/qs8e6Hos3WAspZUNRqhiM2PmILILUZ
hXNOVHPPFNElcazHEldk92lxSDGiW59+gZMzrkwMiTMTDqiILhr7NFsS2XzdJ1MV
DzBPcEyt3evZwgd8sBJ3t44nXF+qIxIi6iPOKhugikDBolDOTxmwYRXou7M007cD
qDQ6Lt470bAfO624idBsbr3jyPGbQOFDNoBvIYD//SP3LKsRTGEdk9JQl44l4woS
1eMGrsrTt6MFjVIpeYVrN8zVfVy1xy30Fy+L+n/PWOLsoq2plwg9ZuWxTBsTTcoa
Gp9XC6ILiiCoIR/hdRuOikfqmwnIsqhp0p/f2oyhL+0WHuKTnpsN/nTDwUCImaAi
Xz0RgZKodHkV3PdjWkKHj7w0DtntxnarA5HDva0HFj4e4CEOrIZ/jL3FVx8ELiuO
/y17CNopaukCVQve+aKgiLWOa5v8o5/9SCoDm77Fu4/i69PLClgy2c0rI4socFzS
mjGcT35epagOvqx/7Pkfc394M5/yLhKFyntvgq2T9+nEXN5C0dE/K2yDv/rSt5bM
NsVYzqVvxwaazjf2WYQmrEzH11DlTN0WOh6iimjaAYoVT/YTzQxompq71UpfUftA
OfDJI8fkY4QVXw4yVQx6w0iyemIZ7b8V2Bdne9PX8bKqjkxjfezVrfCAdd5Buj1D
mXZT70FeuflIbjPElrrRHKgEYr+D/rKmdfeX3uG8Q3nfUYP4jj82p+0htfslN41y
RdIgR1ftu02asaJ2W8guRJweH99l0zH7CN8T4PHSSsC1HnkLk2x2HjSxG23OWGJ9
QguoRKwe671NGb9D1VWalfGsFVtqSeCAfaBYFj8DwsaCX+Ev0KLQogYw3YDv29Ii
p2Ltnangmyh/V3K4AfUE3wDF8BYPMKqgrD+D/xdBP8Dsx4b6HxjPcWqXaRgdg5u1
vtG0V/t6WxnvY8MtKV5mZ2pK3jrI9EAHBi3DVX1jhOREp/WywHNyGwcXCuO7YD+J
iPqpfXnCr2huYVGnKp6Qdc11B0PG/6g93hGZJsEs6eT5RMiiGKg97ItVpT2e5A/y
G/ThcKI2/nijWIdxma/cXZBeV7w9cm+jDtlahYqpoz6155rs3jRA5ns6q8ehW8Rc
U1oaSp0TR0Z/ZRpbxeOh2BeGvyT0hFzMNZr1Hg4uUxmMBjwY9ZeYOYZvwpyf1kpm
cEiS7ximqPqNO56c/7/cWr716GZnZrJ1odgK5W5vAU1IlmtnM/3d9E8p5fXjsdX7
ONyXl4HI392FjhOISCD135ArKRoPIMzqp25uFTjdLcU39FT9mM+U19XJQDHU0vBe
6G9E789nGwcAOJf6XK1cZHgA9tfEiZ43Hkfy9XWGfyZD2Tqi3bPRU8K1Z/aRxsVU
ywHBrwMSsBDH+2h6zAubTCvYmsG7VsEB0fiwvijDi4Leu8Q88c7bNngFAQIOe+Rh
UZ2I+Igy6jHDCJzvEsdxhn3G7QqVjt87HNA4SyIbtT2hGutLTk+Hw7akQdM8ahiH
do52ibrZGkJl2vsyM8lBZyHqEw8UV4r8WD9egCpqltvx7boDJIZyYU+6r3ewnjh5
e51cBgHQkdwxYuZ+sYEW/EuP0g6hECY3Uock2ypUeJ2dic32r8TfFwkthLWBxtlh
P7rfrwpFC/1BA36xtnohowkNIksI8ejty7Le044R5l9Li/i2tG04noc6e13w4Bio
sstx49oI9CHTfc64f2/yvVpkVJ1cQzSAH9F6SYc75CNzn/TkYfRpHNm1dtHFgmqn
zGliAhC1QgbGRJLgYdfb9/iiT+xUBB+UwQuKVbd38B1OF3zTX1oZgi56VN+CHFmR
66ila4q9hRzeqBskxz32HWezPknIzQYFw7JlsamC3UGix68TnnoCp4iG1i171IVJ
51lXzZuNyV4P+VyHjId5lyf/boHsKKg1FIJjuB45sYAsgiCcL5oMRoyFmyOkxd0f
Clb1q4hG5EbyLupfbH6Y/tcSZQ0tdIeMLW27tYQNRzqsv/jRnI0rFGS2pKFBYLdV
kKBbIx/ysd8bzZhPFPBdZvV2pwsNsWYyRxnA42YRb93DgPAaTmi2SqHtqgRUdThS
SrUfJ2BK+O86qx8uKbuxMvKQz5Knmmd9D5uZmASkGdl4ohdui5pknQ37QC30yAP5
mrNyLMpPtWEIyoJRCDBbHXldnW+5tkCOX1jSLXGX1SEpwN86LYDFVCVkmoqjO/Wl
NcrKsv9myZaznB9Qu3At9n8MpAotYmfWbf0CuGbgQ3KuXXrjjKDESydPFgZEJiaT
xe6MACPfc8iV11k7NQa9jA5Ibqr3fw5AIT+H7IPPFFQ7y2i2yenINj1Qid3QOj7V
IsxYgGTiAs/Pv/5aYx40Q+YDFgjA5EDG7RkE4Ko56hcXPqXjKaQkqOK8mkfpRchQ
+Wtdyoj952vevP4XZ7jL06xOLswHpOtg9xAFQN9f+bdb1/i3VL7mgO1c2uapcZ1a
9DUin3bFRDWRkLxaKB2xfdpahuZFEicTNVy1RTYbH+yKuB+LYk67b4DxNKONYHKb
qDIYbg6Fx3PLby/fX0S4ZfRmnVzSTCYcvgtPaSlJHp3p/ZMyqqLg+kEgYAVN8zBP
GJkLlYK3fq72Dm//z6w8D+aK3pEu2eePYvM0zehc1fq47KZ+sNdRSucryppAhJsf
h4njJQje1QMxvbuz/tCMK9t6s3njC41IpfJsMh5oEsiLwhfd1RJzZrJs90LarlZ9
qsU1YQ+EKbpF1jAqN7bFWphXnUF4riSfz+WLl8PvwNRbTGWP2sVbm0WfJDdGFxLz
VFca9znjEhUMJujW0VnUWJmwKRTStdvS4m5ep4iv9kPuns5eJvpKrNJ//H+RqngV
ZVY77cWD1IGdCBOhI8hjes6s+lR02ZnF8BItZwTL4kUtQPB4a84YxYktfcY9InFo
x3+ACjMJDTZAgFF2mq8y170xNBgXk/Kn5mm+cBWw4QtO16Fe8gLo2Jmd+mFErqaF
pMRlT583R12ZBsPlgLrzW2UsFCRLFGj+TQwQmDNw5CmQcNkYO2AZ6jfHjHb+PwnI
uyZgYQY0FPZ08aAY830SRonNFOt7T9zjSZO0wi/9YZX9Epj2QwXbUxupVu3/MMqK
b6AGbtbCCXBlL3je+rgqK/Bg31vfK6yLFWC8HaQoVapIXY+1AKtSmODF3hVpUrsw
jt9Blfj28suOUWjhfj33ZQ/Wm9AlgoClX6kSSGI0U7JaRpYVB5Yn9n2dhrnQLKnI
6XxTnbD7lNpUxsxC6MUR+nIaaKSrxsUYfCFmF8IoXAN4CH4wR7e6yM+Vrxr+pE13
28BmAKkEetEYSWfWG98IwZefTd3KZ5sg8sVyFrMiMdgnO6sMaxa799DJxfAyOde4
ZDiaIfbLDRXL+bRx4/KwcQSgWvMH/iQQ4Ty5GVkafxoF1aHVQBQNsrZN8C9TcL6i
g93K0Od9HioQarcfrBmMUA1cP/d1YzWIuAVp2oyiFQnFCpEp2n7cRqR8KP8vZbnW
OLONXtVSl97GmQwDji0toQHqgEoxtahk7HXBybmW5BzSEK8IaV7JXxX+mKVEAwGj
d14o+ZubA64LpdHWNbpg/Rj4nhZQey1L+WzzkPtTjwmnmrUYi/YUXx2AQ/+26BZ+
MAQ4acelZ/iKKgMcdXWIrB45qpXVu5o6+J6PQZYztVoZMfSRmqDVzLWe54R9Upia
rwbfanvfinYNxuLswqjZyc/BeMLOlAVS/P8H36jGJMGlVbvAfGCOhHe8b5ltKU08
b9V0CULrDMDsQdSBExD95/eyG+ufLTngOsm1pZnBAuaTbqwK0GnShW+xXQ4zL2FM
vKb7TdHX3tg+2hW+rUqSvgiKlayzvFRJ47wln2ZaVvhRqHlHQoni6jptbSWDl9WR
xN26fk0kK/vji4/a3dqivumRl0es9uvA0FTAjMOvgJnu0llMARysNuzvoyZYZGJ5
j+GoP7eLcRzzQN3y31QaHROA2m1lfjsKB9cLrmPrrvL6jFwBSOgTDN/G8I01KNAc
8PoNUNXkA+UT0fm0UvyDnfQCqvOT81BjUqxj7NpWDtx9UAdT0osK1yj3KdrA+Rld
7/vk495IQqav7IceEu/CjHq+XzfcsKHHiEkFpXunyh6xBjSmPIMIB5nm/2T2NpHI
jtsc7NsXRADL5+JP21TH7lXbUITjiKPaxnPRYChWJVXZP+dma35UqH95v5ZZpfmd
8nEY0I61rZpCc6Y1D/JSuBwy/L74N48b7aOLM4DYIW/Ry+Nhphl8T69g+V00qws4
1/zluMMuXhjHzukX1bXDha5cyied+tZx+jbXvcM37jO2bXMV9Mnf5cHTwis1ArA7
hyoA4AgTNs4vs++Nl++f37SK0w9Ce2sltKAwiXSujHHvEqewcR+h9CcF5zgioQDV
Zcw6VGRcxczGTMzhyKDWrSLsk5JMOoF+UwqXpmXciOn+PnO+Osy95zlZVU6g2mb9
YQqFmAX6lguV5LYgg6tHxBuuzfUEAVyicKDbX4nfKQcm2/F487Rs5MzHVSJOAQFb
2NDKd9BFeBoh+WUNvLgXJxgHpEspBvoI0S+TYhGHQAs+RJeY0Z3yQF6LOFSCA97Z
0xwlq2HmxKORmTchEfVs2gFsS/ryBe9At1ggHBojDpcaj+P1IlWNSQcG6QTc1duy
sFPD83o25TUf9O8ioklxr1ZBG0TVb5DyZfmJyhfnb2dsD8osbe428ykKR79t+46U
6E/qWdcPwmC7cHZ4SgOmCxk9u7kb0JrV/Wl2QB7E2aHCv/INyV0niVWZKKwvBvkz
E5BsCrORAq8co+esKPzc6f2QmaNUsVuCKEehX7hIBLpj8G2QdZP7HVi9azQJ4BiG
U74d/gtU8g7XQrSC5Bn4uP6yp/w2LoTjz6wSjMiMGw6qhXhoYa4c7P0qHnM7Jmfj
RL+JR9zan+t93gCTdiP1NnStPAZgDAeIV3eFgKjiznLS+JcQ/ATtsnBMRVtV4GHU
sgLNsvwqRUT6NSfWxhi3dxckbE5vF2E0W8bVMvW+rKLGvqSID2sFx2qZxdwAgKz2
KGEr+cRbno8kIHecSFEVPbfKzu8tPJn+ojD8EoKh2OLY9TvGNg/TQDtkodXe+xwg
HTeMS64KG7pMeSR6UAm7x/kQQHIN9s21q1k+vFFDyHG7Meyo0gUZ5FVwoOykpK80
jmKrAn4zI5Z9T6btFO+srLKz0SomCjcDlBZMQA8Fvq+dXxCaESh69JoEnBx3Pwju
z8zQzR/Icqp+DspU6JQTOSqVyau8Kqa/eqSF/4XxSf+At027Ow6MIiSA7//bDrHd
g9HrZMqF3W/xvh+hVLSwX724Z9F94S4wZneeY9KUySUGVnybPufovqZTRSge7gJI
oFOH9mejUTNSnY8NURcMpnvRw3kXwTcGSj6Qy8Utkv0h7lTA514RdFB5h8jCY6qT
NO3h4KrHAMKxJwwLO12kHV17s0O18x4Mdy8gn6lfl1pzVhZt2aapuUjqDK35ty1Q
3gWj/Qp1mfzX5vk6ULMLOmBXDXo8K+FE5fgicf4roHSaamf9dwI3653rdWJgoLJT
opDXYAg7BUiIvNAa0qDdgirEvyzh0i4hIvzgVFnQS+8WFJOiR5hnSebOa9K3xx42
9OCb3eJp8kwXPKST5XGQTSc9qthvmKWnCQQKvoeNtqUaYqJVRkY4Rn5aI0AR6h8H
nN9WP/Gd3gCyO2cKiUL1BPZ1Ez6IkJv923p/7OEw+b9ZKKeL33lBxBR58q8UpDnh
JkmzIeQBqlDxuwT90peL0h4ti7MsV2hoOHzX2k65fazF2480JxTtGbMxRIf7bMTK
d1OwXRFDMGRsDIO1v7Ouy1K1q6IlTBZC4sXPhgjGvEILLVRPuTbz6lnIv8v8x/DO
657AMy78arTC3fJ8YWi+kwzgi03rwzSCPCdSPQuZvLGg4+tHHiBaKsggHdA9K5V5
IgFr7rqJyxCfRKo9MMrh8kjUXIMWZreoQLLRWeiDFwzkSCCETqF2YJNEU9KLJ9HA
gye0QrodMJ4Jp7F2BQK/9IMCS6jToT0OExrkdYy+2d8RfUzZFiM95Al1cpJJVVBA
nMqBU6Q3FMLM1VCVqMZZTtwerzw2qD70MS1f8rfFY4ewCSf1NfZBtY8I+B5Dsd8j
IyPK/LhiyZByLsgrrLT04CLJI/PaUzErOZBMOFXSELlVVtIFuhY38l9wl9cqIFsI
qAsSyvkywgZPvkz/PDVcH3opzntlp+x9sXryXNhrNt0jn/zca7uVTd5BCy2/WvVQ
jfclbqbLdXQBw7b3D0DyGtgnK2Lq8ouvIjLnPMHoWOtcDn9hCn4+cNcxmwM/W0i0
4uJ9PMa/mZCfCbYMJS/n/JE1VL+Xxlr8bmFq1xwpPBw0QE9PtBdat3LbLLPW0iYe
oUn0c9bbptB7yA0SR8Es98lDtGI8Fo4UwONy092dBj2v0tAiIliY/za+NH9Vw197
IOK/3zK+3O6aXQkjmjrRIQldXcIz/8dn6zaoN0rfOCOpOYcuWg9TAeub9n9mj+VD
eR0ovzoz4rFShX4x0WGeRy27thbjZF1a0bA2F6SgJAuZk3teFWPwjy5/DIgZB3pB
jWXgSXGETYst/h4b8pqdYbKnLG2r0nWOK5zGpTUanZbXVHtbQhrs9Ppy56GRCZhG
MBwHrmWZyzSTSgt2Y/Ner8ogveWpACWFXk/d2EFd2z4wtt85I194IaE73vwN4NEI
crm/r8i9DEW254vXvD9K1NvOfo6/FK67zfKn+qjEv2KZzv2sdsO/F25qRCpWFR1Z
gA8u0uxHpeFSkApIzYrRbAIAYTkxYJXqC8W+8VvKAKPr60WXmV1/UZb8AtiYNHHC
8iJ2mn6GtMf5XFlDejEXejj9j1+5E/n4lD5dVWJ4Sjb3kpUlhXy/PasaajXTagwv
bOx6gRP+/ZQMEXuJlLo0EoXrGTLQHUlBAM6mPCdMbuXsp+T7X/kMQR+u1jlkfxdx
avnPxNaFelLkQm26e/aXfQKWq9onGpy7DqaL+dNsPLcz99MfXY5/+mPs7Ih2hyAy
oUl2XdopmldMmErqxO/h3tNVts01ZwRFxYTDpvIuR+vvyNFXRj13fSV6FSulIeyN
IqV5XPhwCuCWbm76G5uQOM5uv60cTLdII7BY+QG2comEMzWT4cDHlqPDwd/moFeP
iMiqBf/Jl0dDrf9A+v3wDKLePNZbbAXhQ48/Y3lydtYF0k9eZOyr0OrUZKrtj12i
uW1RarKCAfH5lizttbS1gHBtQm6aKI6Mhd6jM+MvbtvtMWpfVi3n0Oz2TOn49C2r
4s7ZT0atKJtcon2pehi6dh4tNzqZTP3qblrSSdjWd+sN3HP6+tdTWoUyCGJTfX9X
mlIgW2ofyMbyZHwihYtqNTatvD6DMz8tGqaLqir/S/IsxHkKO+zfbVKEzk45lLYJ
AL/xUgenk4H0yQZbMYnco8aRgc7f8fSWzYPK2zOTz6Sq2fxOdCbIQzzq8ZtR5Upm
10CiWSK8JoDBvHVpY0lLPCRskDZxQL7Iniq6fLgqxO2r7kOW0/34mmTuxFOGNqbY
a3mbk5Rw5soLtH+uYMLDNaYSXJ+fGMBI2S5N5nSr4tka3M3VoLH3ug9RmyiQPYL2
Z37sTMjsM+kL42suRkEmw58qA1gFD6vXgzWdaeNeZiu0/ySdi2h9+he/kB1Di1zO
ZOuuUeZOubJwB+iCmJOOChzoe5WQICPOtaoQkbzXRhootmgKh6LrdolW6tSCPpWl
oweRq4qdHo+9zina2D2QeJhh2Sg32CcBaaTfUF/U/RKpZmdde+xKSc5vQhF1RUY9
9c2ezkN5HYS6Bq5fPLMtKuRR1wwauMblG2Xjl/f1LBNDHrRT4iSh9j+tYYtkFXwS
+6j+D4IC45AcJZh7gjN7t8Bu7CuPJsrMeoUckKPIMTQUpGOyO/oDexorFCuf8qhU
W5Dtm+IDvFbO3mxa0kczmsPU4Qch7gPorjoqKP5mMmBQ0gxtgr45fneHL5a1060/
wCdKXJDYf8rUQTGdDfpIcDbDwURywIm1fpkpuKZ1XCKu+UPmrrFRg2ZAKIBSVnvA
QpIksfS8XRXLgsdxGPziqKvCO5gUyRZehnZ1Uosl8PwsFTZyxdaYUX62n0h4XBjN
qwpffZu4fuCJeig6ubP52GKjg/NkdpRqv3zbNK7Lhqu4Yks4j2yq66YlOJGRMO0j
oCUT4BWB35qqS0pEXuZdda5ZvIRKn7kcXCyDFOCW2KjeEFRJ/TU7mZwUifnuuNTQ
IbjjNCHcEPkxfwaKHlsI0xXLq9ncwtU7Uw2BsjJZpt2GmKpWtUcbVGTPYvk3eqV7
0aVcUkSUgZHxxcWgqVuTZlZDT9erZgjU5DwyxFK9ujLbTcDFUb0899rcT5LN3Xvq
gRUmxBIqfb/WTa7JKKxkadKxEaR2lgj6oCMRkWFROgFP4WGBsQMverCWGH4EbSPr
F/D/Ms/8U+GMYwAx3XZ48GifB59z9xeSyU+nVfxmpc8BxenzRm7xnfeX+qmAZDbT
INo0ImFdakb9BYTq1OHK5JqSD9Ls36eFcLzuytMNEWOrT8GAx4c5Aa46+CoQ5Bsj
d/i21CjJPYCpH+RqxaXHH8nGqxfiN6Q8Y//5DMXh8PUV1m4uBoi2mQh1vrQM6InI
MFNilAdN0zs4nAYIJKjx16cH+k4Eft1Jcqztv9IPCwX6Vfnumy9lutDeL8PYJUg8
30w+3GfSiOBwDWYECN5xJptUiLUzGA/Xtnd3OuOYJ7sgjaQcTPuyIvO4YRDuocYs
A9+naB5QXToyM1zwgInTAsoAoLp52Dcrhut9cOQPMTeMVlJe9qBokRnjKzYaRqJ2
0QzNVEOunltvycOYrS0SNsKl73blLdGj2lZMWXb70xM2dAJfgpHaoE3JgWvoiGZr
tQ92jjeJGPnIkQJdymMEcH4DogyORNo9Z4qr84BDdN19IRjuWjQ2lqNuyOpixscr
yQCHqaYi8F7/hURxKd+zoGMTBSVbRLR+kUaqaxMEmLvbdG4q972ZSvxG5G7Y2+ot
JqdvimVb6Sqog//nKB2L+Qfo9u72vwsT9PldmekrD6vLR9rfrgCpwmmMX8vqpdm/
Oih+ifr6/K0VmpGXwDJF3Pn5i9/um7ITGxDnsFaI3TiPhM5BHRHnzrqlQ2KvBmxW
+O2l9tvN6tOqJscUdM2Td4hi2c8UXvA7Xj3JpKTA0MQs+WEGfdpojvYNIh0zqNjX
MAeLemzB9rA0oh+5GtJm3e+O+WIe3mqfTu2m+8MzmVLt5SUv5HA3RLUY70dsepIW
3KFgYz+5wN/P8Kd8aVzkXHLTSa1cD40ykaJ6DRnfSo0qFLj1C0Ay2qmHlIX0qBi4
wXVyQeBNDLS61qAG7kk4w4IsraP9+jE8LZ2PjmkhriupYoPj2a0EKpCVqE820PgI
SfJm9yU9wrXmGP08lXB2mEGDyZ+TdSQo3lkID8I8Z3ZraxAZrSyjzTXt6gXIXpJ/
iDhNm8pIdKh22v9Mj1B+FdNxCYkexhN+irypn+3+ptunUIrTpIW6KyLoIH+NNeI/
7eHnepyY7dA4fJjRrfkJdJ/50T4vnp8fvytPaerPK6fpoDO970YRlptXl3/ZUMUc
O35cnstSjuV+c22cHdEWiT86f874SKgGzNkgFt7jU7lWSEUBNmtqwwqxvJDPzfyk
71QHiuNPjumQGYclFGwYyWgsmSYgrgbeiU3usIo9yxs1gnL9AVKt7Aovv40to0SG
yI0rler3UcRy24ht218vvJn77j+Ei/uqpjAGTFHS+uUZRoLP/c4Mzq8i3UBofCrC
pnWh/JaUOjMkC5e4dmH90aINx+pkOKSEfm6QeD+4LfNxBoYxCpA46DNMWTf4tmUu
AEu82LyXvZA1RA6Kx97Fx/Hk1B+YHSm9EtqfpY73rk459XVxaVIaTIKjzZlmMcn/
8IlxP9npN5BalKjoSLT2X4xawvzjEnXqgbiSuR+zkXXP/fqnr1hzGqlKMCj95d0x
deHWn/9pOJ2Ym5/M8AtoksKxG2MyojaXPcKMLJW+urXnwkn516HdaupB+gyIfQXx
vvh5Z3rU+9Sb6K9ryM0KBYO8ZGAU0GjP+QOdT7gXW0DoJwSgoCQzaxLp0PLe4Qp/
SDimVyflHpNEGE2IHGxJTwRlu+zsvXDglyJ4mD9l9acfL8kzWeJtPeK5XDHTH85h
qTWHKfQv8hWd+YX0WIa7sb91D0p2CnzfExcxmWdDCP4ToSA2n7wwV6p4GyLYmxiM
lyEZqWxWcSpME33g9RU4IshD2/ouHXaUxK8Kz6L9dm3FOyX8769G/f20MCfm/cQj
datZ8KVQeQrR09Oje1AKJiamx9LVzE8OnBnb9XZSRZCQQvD2+kI9z9/zTqvIT6L3
rLUz4a7K079tw3U7gPFGXhMjraLgFH64ZF9E7+uivFTHcRQPxzOV30kxvj+O43xZ
8UTCIsHk7g1c/Yo1OSh3iNCOVBR1tmPWOVYjkoiR5xKqe9q9eyAq72hzvNW5t5oq
rnaomW9cxD0IjJldSpm44SuKlPa/EL28wUK0IwwwXGMU5htQQjafA2JpdHUFAOyu
lA1mune2hpAZOm7iuBfGmUc5KFoYUJoaECbBN+8SPO3PRKjpZQMR/pMfn2IKSLQN
vLwtAvvKlPTBk22ODaY0HysvxPc5+e5eHp3qywjzBz2Y1UYx28IX/XYyksN5ELMO
plDwAXhFREtbrNrd6KB4PrhjWoqLaNiY9QbMEVuCXhR8mnpBj2obBoMUdHGwhcSO
4/xe/5lAmvSPrVCxeFvLA1ro+QWS0b+UZPWHW3CJfK34SFdifMV35Izc/kfQ4Idv
MubATkVLB7tRUwDtDEeOMmfJVcyUX8wPQkTmSfGsFENLTP6ktNrlaZDeXV5QEUjP
51YmHdkvdeFyDZoICLobfRsGV2NzEKFvheTGoozrYgKTer7YbGyXkV/g6hZ0pmC8
GX/efr/OmaXOyvNmV27889Y3MxwopoBlWUVlXw+yFWMrd7y3bFIeIwVn1A+4K0KW
BlGYvoH0eQl8R1WRhEPeqD/yZbtYFwm3Zfl40cf1ZkWyxk/XOwd7oFPueVplyu9a
+8kaObdZzPVRdhag0rMprih2END3cWXpCbnkVNSTs65TFNT7IpM82NAiyIlpi3hx
QdoGY/bQVS9GNeHavEBM94fDVxa2MsaVwj0geFKoy1ko27IGVYctxgcBzM1xf44Y
QTn+fEAqCgh0SLgi/fS0UiVavrebn7xwvMfZIt85NV7CU2rKlUWC2tQH3J2+A81k
EJM25uJx6Ts7UdCxduwrOmUr+F554cO4PjYWHO/hceVgPW+ksxdvo3yCA2uyVqoA
5f6QZKJu4QUlUpeNaIzbKqyZIpOB3iU5WymEZ66zJhlIy1sYJx2nPoE66ll/XcGz
fKOLOP7A/+4xik0HXlJIH6eujYCjfcYex1hNQhhX2SnS2/QjNiTq50CsHDrIpaaV
lXwRiqPvXy3Ha9aqSPN66jHyrveRqls2O+G4Cef7Ymidzt+I6wQL0tLP9XCeMo7i
0f5OTMkLNIF9LKX371TTDL+qqGYQdABPaUoZB8hlMveaHY716I7DHTCy61+6gIMA
EAd6skcg/9iPz9p6pY9LDhgrtwlWaJKIR/nqr9htMpn8Xo90tNsml/E9df73VPPR
oPfdcby1wIAMwqIApMxpIk9nPJx9Nq94Bsm/Lv06M/EXfft74IIQCvduIxUO9dh8
S4d1mzj9t06AAsc1OUPv+ExPrCS8eGCgRzOCDZS8vYoFH4F+0hlS04FZwBbvdT+y
TwdfpaGINewYDFVyTXJEkgjEJJ1nYbtyAf2qELSeAd0OmiGMRVyPjuDkmqHfkDKy
EbR9LaebHNdxqlWcOXDLYK1hKSV9JY8o3ru3SfF1BZNaBafVghjmtLO98GUywvag
OCy6KJVZUnJU4LyU0Lk1PphaIlgGdlNLG+VuJIWtwjrbWKmEfJB+jA8Hfk+GXWNP
OEDbEr6UK/yj2HTqBTPNjPKOfuOILGxNGviDOG8cWvWheMBfqk3S0X1RGR6m8Bv2
4+9BPheDAuUDeZtsHch7qB5JpH8JDd2fEE1rfjHgXHjWc4cxUsuaZV64N2+3s0Hz
rpDK/yiAtFL76YqR3HLLa9KBApDO699UkzE+uOb8VzKxvRW5R5A8Hccwbq2aGixl
dLrgmYatc983yaBE6yEa/UvBgHHchznEwzraNWYW55xlI8H1U9OUhuIW+BYNifn1
4mnxy6WB3jrFNmNLuhEThO9CoAQomJuf3x8x5Mx4o13mnF+Jq4uQuIdbOzCwfHjz
Sv2hGNOrDqqFfXRioPJSYtIferFo/dmxyt/A6bjqk+VUlpB028X3y6Y8RrVYF+R7
TCqVJwPaea0vGgBGkr765lTHRRGFhGmz8cw3h61LXDO9G2kcjQxxJnHWJTxiZYow
W2h1D6Bum5g6Wd7qnlK8VlokPT2CJiPwgsv0+3BI7Nzc+p7zZF2tIzpcdLQIRx18
+6/tWjrxPiVYW8jlz5lrnLRUWXKbQptBIzhNOOFRChKKAcpNnLIgaeRaOb6lywhH
uBno88SEAYkhHDAjuStPS8ir19nhhXD7n3PrAhsmzbaNwEFWBNPvrMMOD3jXzYd2
zi8y2gPeBwiWrs8s5O6yBu3iCPlP5qYWAgDj8yyX1RvKl+rC9T/VhRVbd16HAklL
LbLBMPSw53FfK0omOxvRGriWK+5qfnonaI67bhS9FnDbP5PMZkYn5uAnc9giebDZ
om9o/C8G8tLZZpRS4n/BtZ/NcQAa5VmJKrZrRLDAxxQwofcqVSo3OYVduhdA4H7s
UuOVcRA29HTanEx9QjjUTdRSMfcYA5hjOLGTgcmjp7ETTEysYcQDhNP/qn3d6FSH
dKG8sDDmpgleGBIb050fNVLstWXL6ZHVoPLeDeBjrzTNENMqmKBkkDYIxCxuUGvM
1vwd7SDfLd3kebVGu2WCCZF24Cy3TShHpp87gD3ceCBm8La7IaxERC2Nwr4VUrac
ECbXjYKyQbuMsaptFgh3BzICEMD0I3hAU3rt3PRWZsVgOPHJvh6jiL6ujKyPfZwr
2iZtiZvt0KiS0lBs4MtLZ6ru+sO8TIrrrmS779bZZIz5f0MS2fzBfz7aKUJ4CIDR
viD/KaAWxo0aopHgYDHI/aULEBdZCY7sWpdoS9MVAgJhN1EvbemfV5lPL97I1SLz
JImNZ/26VSm07rJOS4UHB5X4imgMcs0uApzSiSw+LLghSewb+DDWLXBUraDjHNyN
sMGkq/nXV/ybNJGuRALhXOYfpNgPpIltbXFfbG/XgTJxRrI19/1y6GQ2LesaNLmT
V9B6/k2u271ZPEe4o1eAPlqoyIP8gcIvOWawlDxi2rodyvX4aPQNOvjY8gvaL6xv
l85s5P6CtJ5FyVSwCbdBUCsiKLulLwvhElVE7c9laxUTBnqNzkab1qCmuH9Rrq5x
agCxwNnGC3ADjfz3KX4AL7RGOY4aTlpJ7ykKnugHgmosLgnlbhmJIeSUNDID4H3D
q/kbHyzFm4ZrDtYa4di9aKKHPO4jPADz7JiA8DVxNm5nRg6yOMIT5R2GvF8Z+dqp
/ot6mT++gLLwkKgghXSpPo9wH/dKp3eMOEx3sb5Danl9Hca239pjO/Esd4RnsKPv
2BvD0sfItZfsBStZT+ktKlz3uT/cvfRblb0PQWt4Px8AOtviHTNQFRXY9Jb7uoDK
weLD+c4gRX0lTkcwzk3GaDf2wr72T61os68sZhXnsKrQ9YrXBgBOdY0T7GMn4PUE
Y05fkQ1/Akc/zeEfe00ForIxiRevtfGS0atzVs1qZWvnbaAp1ypXQWaseav8XBiv
0cPI20jTVufK3rnILLTG4vlgpRHhNZd1WyO8E0OdnttstluLwdl9j7A/gh6ZFBgx
I4YzEvROLe4NuVsaV8exhls2WhGPgru8+kRR3putLAJ8CPlUp6Oun9pBgnmDP59y
PG/gqQYctDwaf1FSe7ZQU54+wk0h4GiCQIy7xKpuESraStq3a5It6pFEZBK6JBSl
DB6bYjmbyJwX2RWZ+glNUnT0/HBvVfpfwdBq7VL40G8UHhcMwtjpwUqobCSv0BPf
Rwfc6/oM+oVyth9euGA/ifFQ9WfY4UQmSnIfKHi3o5UIjUW5NKegGO4TdnW84Wl6
vyPk1Nxr+zTlQ5MOEY5+DmPs30fQkGQ7hqY2scTEY+cRNlZl6D6WtV8rWS1vVjE1
FNMrd5HwPMc1P7sY1g2leg6V5fTLoclfXpCE79g9VgDwvKXh0m8DiYGYh/mGZytz
0pLKetSzfjIwV+lq7TsNe2KcIuCOfbNFP0mMPGj0bmmLsJs4Q7bhn5pW2Cf1KREA
vcausNZO2Yp9h2VrQhT/VeYJNK+3IYQH8NTJRRywHh8iN8T7er19waL3RH8VSg9X
Z3MDBlInFJ+16jX3hf/zOKupo7/PLyfoT3LQV6ppi9Vt5LB8oHfLizTC8nWSEOyV
1N93yRV+Jz8SkV7d391y/VBtLz6D0VFSCdR/dst8EFeITSSD1pMhstLvG5KS/Vc2
tfxcUgbIFRfYjQh0e1NunvPRd5FhRkn94Dehx13gMO084o3ioNlUNpPah8gSN6Jk
qyxWSZqsJWlr+UbuP521rB3L1yqqlSyTy9chV2kSHcbuY1LR7lK1rS0CWjrgsQyM
mt70LU3EHtvxHTyz+36VUvCEGo9n8W0214qZrAdAxZDfbCeGxER3kmkImsjT0rFj
rYtt/WI8NVdlWs2inNriZAUBQ0dCYuLFdp9ysf67lhABaezc8A0CtT9svdcEuSfN
Jr3r91ZVCBiHkG0Rr8e5kGX3OJRs4UbR1r2Abydxrhocn3R081QcJ6lF/pkAKEcO
VL6ulhC/xYJu+1yPPeCo7B6e0U2XTmnyLcRf8+CZAkh0bfi2IITYpjl2j0IEF0H/
R2tT6VnfiushqnzcS4BHtTaz8Cz/CwO86DtBAa+ffCgQQLzAA4Ox/WWVaao36efL
ZoxMxz/wVGsswII/Wqfjf22Xp7g7BLHipRTWBItrxjGIPFdJx0wVP3LAnIe2JOCd
roQ2Kntzm3cp7EzQlUpeeYzr9Pfm2t/Od5OGAgJWH9TZ5nKfkhj9Xo3/JiJ5scYa
BDvdaPR7H3IfyFPECflKDRkUEMfSVDdCl0V9smNN4366HvaRdRHRmV4Lzo41W9iD
ZfEg4NLLSZAJxBfhlsjviSTRdiZGX7jgP+Bt8TKCsDN9jHgVpEk5iMMZxvAVsqF9
fqFWEPuZHj3/NRSJCQfqy4RVctupeSfevJY2ChV0z/a2mdfX5Ze33SVLtnNUEI0u
DBRg8uewoi+R1c4AJQFB7XEF/gIZF03e31BnqklggE8=
`pragma protect end_protected
