// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:41 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Wcu0+Zv3As3uxcrYT7Q6UcWOgLU9wdEE5eYDG49r8BY7BUSDAOHRLScwho586+Ud
Wby/V3eOjTrRuZ+aHmO2M7zS+aAMGaBTA6xu51Gvh8wrDAeGqVwN5fuNXwQRYzeB
xVxK8m7OaUBblie2bl0pQ1QZNVdnMo1p0Sbtey91Bxk=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 15744)
l0O055Tg2jy4vT871K6MEzfDQA2Jggy0Ewq6al7GHbHmg9FASNuddk69xcTDhVFS
q2D95POFIAaV7CcWqDmKx9Je5m6uqDzm4Y9ZEvLe18F3IKSGNqZxxSNHOJCk1UYJ
GT5vc07UOjY4ZJef7rNGwxmk5LPjZA9QFLPgK3fgXxvJ/lpzCDrNGNQbTwcE4Jr/
mdnSOIVUg+PickiWSnnFLqwkh4ZdomDkmqeLYLvmGEG7T7wKk80EQIP5XJxxLLeg
tj3EL0NbXzZ6SN8d3/Go4PJ4e2fB/thCPKApjj1UXtHWrToADUY2wR3g5spMZVy8
gL/UNiepN8PyjTrLY20eMmv2NA3vVLOpayElNgfhimLAxorzqOCxuEbqN1QREvsx
CHw5/Y+peu/jBg3Mf9arUayMKoDJ1YO/LcmUBD+sKhcAxoSIcXh47ZpTXTi4OwaC
G7kRRyoxDQ6wUSg6E/X0qWcBV8ZgiGchn0c7oGr7RFnyF9gtIiPsKyjIBKv3ipmA
8Z/HgyOJiUJOlxRyal6yl+13psu3lFk6dl5AwG0P6UGkYwVKuUtCJfVW6J4eWeVN
c5BARfLu8bqIIStOY1oW1Bdm/OUyZ8KBmC1BGRFLHf4dMfi4qOht/sE9ge7e4S8c
kUnWrTKMJ/596QCQjR76GvfWG80+Ph2Q5Jti+8AsmQmPUprRNPHmMlozUpmk/Iko
1/enKW5tGTeI9dyvxrkBO9HydCvMQHhDb96fNvXmgJRvNrosHZiWmZCVWfjiTSvc
YOA0LhlRfo9tUxhR6DDUS8/r+PYl+oH3jbK37bYUGEdzugSJShJHAXYSb2B5VoIV
oV97NSJ0JjhjQf4qI6ZjR3YeIwazbAD1a4zaloOmAOiyMqoFJJ1xh3xqWT/643XC
jf/NaUsb2KwXwm3by9ZRr7Ow5OfPov4w8ct7yRCfwOM/riJ44X0z//IGWOjGUrEE
qf6PMi1OsRv0sRxFNPG5IQ4VZW5tihxxUYpdkRp4fKDBhKrRn4f+ho6gdG6Y4v4J
8G8KcqVXKOyyV5ZBYMgQ2ehVYdoShP9i3bRj/Kex6hVshpv8kYJ7NN+FZ2KibfCb
xGuDxVv6p/eLJKF6NftV0vW27AR1LQPMKzGNTwrUwttKT36/Tyna+S7fU9G/mKNo
P1j5kn31K3YUFG0Oscp9RSVRPuApGX30KGgcuDk3qX5vIgZZ8urM6Ltnpys1zdKS
f3SFX+FoIv6yARqNd1LkUDSZuNsddy76BEA+eSr+/7M07yXbysr7ZVLr9Dnd/aEY
fh6RvIdN57ePpRwxnUaauJjbiQd7fXfgJal3c9hF8okgmq1feUvFXG2zlagcpcoW
FZehnCVusD8jdjZC0HygBUB09hP4SH8jVpxccc1cxjGm4WoBLc+cVZdEYCSv9B5X
y2D+k5Qtw+rF1e12aSxGXCgrBJvIyqCCacbSCzV10aXUYdDw7qm5UK3TKm1Qdo2h
Sw1LWjeWlUIN6/5y6XU7ya3k2RpUQSU/mEg3qDeyNbpw56ymIGaE1jUf5hWZaUrr
NLrqYYKTqJfivsIAETJ0hkbOaHnFq2Xc5x7t1vp0XQT1DGQMfTvgtRJyV+I3lkxg
1UJbOy4YLunTDz6+zlKedgpOCYGWtSTIy4sZdQTwbnHKE+RWDQU5L2EFtO/ZCvbj
J7YRUo6UV9UgXH3WEnq8g0k3PwKD1gTY4mhT4EA2+KgFPSKRScV13AKe0WiboPeP
NIwoABKenw2sj2tCTytBooe6JXiPRP2GTJtpSR6J1klg9PGgsYPxRrHIPIcsSL82
tUsd7Q5PIIWhF3HShdE8DaaJg12R8mlTThVWnNNrebjKh043py167bT9zkaU7ANy
lLM/fkEvHIQLUF3O/4B5pQSKCI6t8PpC3iBGtihpcYoe1CJ235tGRcfnXYswuBkR
5z+42pLjSVvO02BsU0Ljq0higsHZsXnSLHXHyMCm4WZXf4xCLADWKLGjaaWLdcXi
u0D3Sj+gs+jS7CuA1kd0f7VGrpE1qCOOK+NIlBlG77CmcrIQ6S0k9dCpbT23HyTq
xF/QdA85V6jkmh4QYCUovdcJC7tPVdZ6WmDBuOErpTu2+xarFU2DC7jHO5ZrQwVM
H1gDZH64rMu13cK7mgQNLPxNsU1xdjdf0/soM7tj6xwJ7Dm4I6hvIqnG89rTVCO9
/o7rkUa9GY6u3Pyp99tOgltGfrBHRbE1mgnn44ZIpOB95+Upu4pC2MMuxZpok/sq
LYtDG4vmHjh9M6QlPsj4yALzdT0YVUNhP4jfup6S/4VlEZWHS/eIEGzsjHZM5Q7K
QxQ9vUFoQU+NEEUmF3tRaQiOErB4pZSsqbHEBnpf5p98yVbSJNLb1tQkcM7wuzo+
srzQb81C9eBVxk/p7pL8FNI5JNquY46cL3fL4TnWQZEDuPen9fZPZmuzbKnPJhlW
W8+Z9SAQwYmuEmz+G25KC008p12AjsCMpmXA9eNhUeSePkE6CcnDlCmj6cT/rBBa
ItJFEggXhq810BvfFFIpieS2N9yBMXEk+8AyB0QxBT12SOwN8Ov597fxwXhWqKkL
WGOCjf7gkAEz+UeNyCDYmaM4HYPLuQTmL+Nb+xU6qa33epUXW3brq7EbTOf0vfiB
bwm4gVfWrFuldOeeQQqf9xj7gvzL93WpTR9XradsbNlMOCnp5zgTMEfCf6vaIat1
EY0RyPqJOls3FP9V71R/n5UKKcKS/0G8OklBjMtr5lAXxyFlqHbvEWZplHMEx/vR
Ax0+kM2LlXF9bxTwW4T6k0aymhXS/p9w/oL5RXB6yxbCHevyiGEZQn5CU9kdRfm4
DNVeqStKssmJYNRMz9rtER8hkfYdGX6ipuSjAjisC3/6oqwwCjP+LFxdKYqgt5KG
F6xBtsr27CQPli8v8Vo1V5Pyq9EItCXlir7kEgausqv2nl6S6IfZa+1lT+dfGPH3
aV0yv17wLMQhGjR+N0y9nW/EXX/hEm4UJhnJBmxgbByb4g60Viv4Zjn0hhmDqxBw
ndvQ6/DwWkMAd6/qlBTaTw1E8UGaKvb0zcNDh6oEZe1NtZGSUiu9cad0PfuO7HBX
w1zt4cmRC3vdB/DJ/d05mfbLf763uKy4sYYUaKJ1P54+p/DxdGZ8lhrAEf+77YAP
4YZ6sGFqqfgMxNUcT6TJtiSjW2q+7npR4qe//HU3eXLLrOBLs236pQ7DnacyJFxr
7RswCpxoUqkURbvCx9FNTQp21eyLKnYWXdip+4FDITmrwf8Fd2A9ZvslISd7ksAf
MpsuRr+hKolxWRbiiThcRU06WUebaNOtRnDz7qXf6jjvDGE+fVLBjrxbCVB7veJp
NBWa3CDNF3iQqSOxsiib481MO8tUr1ByyoDcNB17mH/a6Zq4lkWYskZ9ffNS3Uuo
QhifH99o8U6X3hJdokvKfFyJ3XtoXe0wqun3Z/H9WpnCBU5XRgdDKLynx3G60ZDz
47Jfxu2Uht4SewsKdG6in/pWcQZslpMFF4OpYf3mov47mCDltQVugITfOlC4qcGp
4thXWceE9RFn16Vy5xM/z2YIhpSLSP4pO0+AcDg1QytkKMCCJVL7zKEYZucUQuEh
hoEjJldTGQaX4GERjhIxr7XGnVvGO9wEj0+sYN+SfjW2ad4pj8YVaKcicl3ZSn1F
HGil7fMTfJuBCHWVhjQGL8rGqfNuF7nykkJqvEeB8jnvRvh37X3Qs9Dxab7HO3Jt
BsWzEi0LdvB2COC7OFVlzMXMvV+r+AJNtKFj2vtq9BXVIF6kbQfJNMxSmOS+NzcQ
Bk3V0Va6WqEv0LSBt7hiFW1O2napcQCxHZxFTsSLrB6vHKq3lsfaPF3OmOEtmhLb
z5rtRTHPapwgnBqK1itoHHJhpHUie3aLU2cZrwaUIDTqEUGUiUkBrby/RLKGv79w
VCFSN6P4StLQ8hJVdtdfXpcvgFZoPLC0aWfFBl7Cer+BoBeYeZtGlI0rfcaf3ZxV
cyqM34NJo9cAfGZuS+b4D8ppIl6IKqBnj7Z1VG6mA2J6qD9aqa9J0ft9ZQgZl0ES
T5YrMy633d5bEV5GzaAjIaLXvStsO8+7mYDgkJ7sFIatseEBWTdytRksNs+6ir4h
cLSE7hUikadmWFcAh/ZpMx4n16wSUmTIAYGYF5q1YLRADDyCCiQ+o4WpRV9dgBgG
PNddGmt+tHQjW1PZT9l8+HPQV6qiFlWx1mComJt1BmEpM3EBFMudLqqd+8EbFVMQ
dvvOu0Tv7D93dQHiwv+5NG1ejmuLJJrMG5lBu7873TO1Fqx8G6Gf1i3GCFi1/Pnv
Ackpo5IOZxt1GPF8Gp39bcO1USlwTyEsHSOUOXAmKHgaoTguapS+yGSfW6EnW/Bv
2TnNX8pQjUsYqyfbcZDjYvyhtFvI+KfayMUSlhNfqiKHT+IaYPieuhiLTsxaYAJB
QFujOTF5Fp1mcvrq3Z4iT4qelxCUXfxvpt3JK1jnB8LBKiG1K3GQ0EM8GmaSyH7n
YSrRBe4QOtsZMcYtpHizV6dTTdrzXYumWClnwLmlfze7q0AWzflqg1qY4LsIQ8wK
gyZunxiiWthN1Tyr0RmOOpeBmXZ6d8wayJWDvknyky03Cvmkwk74yA3KnCb22/9h
eXUc6yEXloL7pfZena2loiQdLiDA/mKbeLZQ3AF2up49IlD4HBHYd94VnQ9vLXII
3MtrbImyhXzcCIcP+aTx3EWFUuHQRg5VWdhjpLUYVCTg6hLoHOJ0ti/xxwj3BudZ
kXiu53bfsD6+tFQA4jdyT+ncrGdNH/Q4QirDb6vUITzA5T286W+xT0axVdi0Qg0z
V/ZCP8J/XT5di7D6yB0a6+zvhr5jA/r/gajVeTddZKRGc7TSaYuDxgsR9DNGVkuX
3rzMMF9whUWn2TnX7TPOT4mhRHlBTmtsp/Ub1GY9AKMl+GfSXycIX2NhZ41Q+ZcA
QDJLUnkdiut+dGsqbMnSabOYcpZLONJlCdFEzmJetKTUrKH7Y22lDgUvcB7G63U9
To+XNcsF/TGdBsNUD7RNnJQYp+vQyCMxFf4r6tUwajiu35d+t5Kckg0HukE2kn7Q
EqEg8NQTa49WCDfeQnUW1/g+7TCBtGTA9cuYizULcT2CNBoMTJTXxxtJhG/1jauD
8AIMfhP/de+DkmLSj/eEhEokgfOUCliWz4Ur2oP9EJwYZuIZKD/2SMpRqgTrcf2J
1PFHRMhyvYl8ba7BCwNmcIjrsl7J6L6pIAReTWpSbScKgOwzRdTTHCg0Bv1dewAE
5HxJ3Pqe5HDH0bolLDZ33+ySW8RET7ekspdfCL0UiSNF6yv+VDaJqKhoFAHqnKoH
KO5yqdDeqyANCaJxKdeUAHvP85qz8nsRSrFfUyrCJFsu8J5PI98hW+EM12eXEtcA
s0+tr73QFjuT5QOkza9eAwUIMdFEv+XdlC8kvLAaqU41dKAW7/aUJ81ls16Klng4
vJZCLgeLicY7Tp/9ciCIsmNI6JOL+/sKrXW7MiGkQnGYpap2ShEADCLRNRtNZWA5
/N91OZeLOLiEwX2NJwFw5hHKf0mTDb6IvdWOp4IG8JBllEVWjQGqZPuyj9kOy4WB
YrGQlT1dIJ6CsulJ01tpHmSublNJ6hISej4cqmarJF5Tjci3Ult1ciGOtJ0Y9LuW
dbGTR1Gd9VnKIZFdUw4BKUjX1AZgyHo/XRAQObm4xeqjnRsm5wP/K42H0hkNN4VN
W+wEYenCEb4+7X7MpYHSVZA7bO3/RpxjPBeKDRB4fzKxjrotTKCw3IOkVp74iKxi
nng+vHovyaRPyvais3rHy/GLPeIPTqotXCxe23ryVY1p8gAp9LMW1qjB5vBqdPf+
bEbV37dV+kPQM2cRjy9YCza/0rUBhq39AqWs+dM6b1vDiRuthK0/Qt3EIHAPAPjz
Ugf+zEWAHjTfAESMl99Y4EiTkyBNb6sXmHQxGtFySxWGur8Y2xEuRH0+rqXDQJlf
m6MhsHnGYvR/RjBmcyVTCgKOxiAKECzOPZBOD9EvTAxSy8hzZoTsVfqyxgaU10NN
JYSFX5/dvvtm2H1CAXYxYCQWXJhQvsIz+CZegd7YeR4AkQt+2PvSwG502rh/Rwp7
TOKQE8jFEzb2oLxc62eR2PkAj+TPXeK8/w1s+zuk+kItDZvIfmBhj2WeEACixd+u
ohzVfzXOQMrDUkklOEEp5zCmsVDCoDW0q6JiunbaMmJtlXjDdk+1HAcDj92OfcW+
D5TXihLxFvlDHwEtLiKN8yKBVJCj0CksCczkS3H1Qyx+pQ8ab5izjKCAM+Eoz+74
eftQkJdlw2b40ocTs4QwoWkVeNJHAWOIR9dGUxLCfjH57B4b6j08CtsK0mJM4rfU
V2XA1ePV9JLt3MsT7wEpsxLQPt1TV8V4BvFp2xDtapN1y05mz+hVERp6j6EYWSX/
cIhziD2sigWXmAgcZOx2kAqchG1zUSSP+9Du4T47z+tcvzqAE08DkjfTEqt7+CjT
yN193e5S2ZQrIjyNlCctmZT6uIkPsDERUcQqfluo4nEC/zfD95Y6ExgUfAuUrwRD
NsGWbC57qQR/LchZNvf1bKMOjCYtw4NwuhLRBrV9+4VJRUmKcQtkaqZh0Mn/rhj/
Zor2Hhrdb7V9N4p7JByLsd3FsXg+vo9i3OmBi10HLN0Rj9e2tqWnfQFTUhkbJJpc
BXme4qV3E5KERyFWaXDG5oC/pN0GeqJLsEtMrURprLWs4JafICr73cWE35dm3XUg
5wRLmbrK1iA/ccuU/wI+3fRyM48WM7FWwuYHWdOOguwr99ult+/ZB9XlSDdi64hw
gjK6BPdeabHC4E4V8yP6gZB8Sge0qr755RGoYOC5fMGgUYTYSHlWwAcS8UTi1Lx8
JmUVqZw69FEERJ+1pkhDpOjxw11RbzvRJrl2dvKXfEvSFCxnddEKzZuOtdgVvqMr
bPuXjqDW/7QKgHyO1u98HWJ02Cw/LKsczgdLOO1thB4vpx0WmA0eZVcznVMjaWYF
da7944UTkszCqjZ1Tt2r9hfatU7ltxgN4u4PgUtNJcBvC2T4tS+9ti17i4OaotTP
PKrz48ET2/ltnATukptJDJ7H1NK2vyhiBe4DbIRDZluDeyacsEmHA84gFRQaMng6
sZAzwFVLybeRJP2D2cT7GNc38DYZVIgu1rxbV6GYXFli+Sb8nwbDEJ6tz3A2vKSC
aX9cEzzhEcsZSogsOJhIhe3tDpd2Qq7m6fDCpz74FCi+tPQYUxCh+5lLJG+IVgQw
Wrai0DUPyzF/ZuALRRuFE1n9AD0Q2IfTwa/E+ak2521TUmSR17TtLHcfBx/fHS6D
W4KNz0T+uYDaa/lJUcqIauTiDDYnd26SyAzIG1Enh6wJOrMVB4qqsaLBTZ9K4mr7
F5Viu4XJ1c3DzPPWAT8QC+8BgV1foUxf1+x9KptMdLGGl91WGKfsMMn9LP8KHFW+
3TXYf8Pntlob29tZ0sJKWJBpNdWrzv3ILeiH4TJvql7tIJCH32MSeNUbV1DGdIgy
Im8Rfv5ObRUGq9A/7iwSw6T51hSDA77i4a9grWCudXU6vH9xvDc95qe8u7RLKYXC
1f0z1KJN2k+NelXW/j8R2ezbM3hezSbab4GKlfQ4cUDFhTLZAoKy88dLxhwBoLFa
u1TGSoQxf4cztNX2MHL3B7GYl6luurb/23587Ehtlw+nYi2u6PBXegs8PVGjhbwB
KzbPDIhBVTUzcHg5B4AKKYVK6cZtW/KEGwD4ZEZmxMszoDEQg2X6BoBLIsTn644y
GRlAu9fTbDJov6GM7r7DL0JRwonCHCk1h67v7Na7TSRFTNltmNH1yvIRkprOoWZH
daDyYt/qr3MjNuZuYi/JifdrJn+kNe5UxRfIfZ3S+k7tJDfQHFZihYGGd2eI8yPV
RaCgmeI3pBaWVcA0FS1vE1UEJtlFuAAAqzfTvP4Zq+u2w67uWxqy6+PFQojUUcHh
nuMcp3ppajyJYRBGGJkFTXmaZS+vU9BbkTbQizv++iamT/x5/aoPgXL9g9jhXdcg
oo3bCKzaHul7olgE13pz81BBJzAWjgQCBjaQ6g0PQcmgStuoOHdjw7ENdKK33R56
ks0QftGq83NEWmFV+bXb4/fidCF5b4e473brSC0ZgdB9W2xo5DYehBLjg5vpqpLi
qoeEVOq8Yw+2APdygACgxKMNTcAyHvL3iYhpy93EvoSlLRMSwSY0b1Bu3xkbcuqj
rg9EJ/HR+om9KTmJQGrpRdmBhTOnul17hpAjq2lTzk5fuGvUFJBCejqEr4Wg/7nn
kNXSoAdbSS8VZwZ+OOtt5UK5ervG6ArqrFJ+MlBzOS9X/8XiEKJDRqU+wcO4qsdr
Ec1OvZZC6EbSCAav5ozo23QSBvKxFiVH/Jlu7lOw+5R7D3isxGjhQ9nvTi6eYpLI
8ryNhr6uoqPm/IOM3VZDjiGdcVt5Yx8F60nf5TzMSLrTWIFAtblkAQl/QDCuh8rr
n0lAkgO/c9VAek+MSSwY1FVdJOHA7W/DrgQyiMD0d+D4exvMmWu+QdK5u7WQXcv+
F3w7Yul39WUWnWmjiTBiDZj7EeTryIz/8ryCjEZ4fSQlbUOjJWhJy6GDKoZbDGkq
IgtgkFlPi6hh5tykDiZXBORPLfd6kuxzpCD1VRUksca4OLryZTVv8VTVR4bfTssC
REW45uHGClD9scWTJ7pPschnCYZsza6h6FFJBhZQ9LpHOY40rUoUOc5QxiZMcoxU
0cN8kBH+zZa4bhf7wauFrl5ylyhfulbTcGs8xzMqAQvwr7WdlsREbqnXLfSUj4M2
z/c4uRDdrYQESFxfx3qjfrJx0jqOC2ZqmR0tPrQlMdSpfRyzy4Zb0bYgYUD6N2ji
ATAAbfXFG+rE5Lq1JbOQ7DHwk6yebO7CUS3jKLfBApcarcGS0nfWfGJub/waQT6A
NGIYERLpI0ams/FNMNU/Lq2Og3PP4hEo7I1mLspx2aNnC+OD/f3ezqWBghI4kLYu
LvHKJi1MvE61PnLrI6VxrgXGUF4KUfCmDMoVUI/TH+/7tRnayAoCvBeE76ExBl5Y
b9uUC3ZReRUIUWyB8Z8JH0MzC1T+z5Djew/p1pIObDNQwrZRSvLriImNqDanhvUr
VXVI9yj2Z7LL7/gXJA+nGdtNYkpbJQzXCuZN2AmISOx++03PKI/7vY8mHoSnexF9
ZHf8ZQMCc49/ryVkr+bXa0BtNVZDq4GIzdHXawMUxq8M4ha/01H/vqtqxg0x4+sJ
SkRc7cShAq4EIndPg9vcKRh8DwDtF9RmSQTozJSWauq51bA0xeBsoDdW4iftqSN6
pEenTJEH3c492GSjuPI0QP6i6OKHMBuHjZaQ4/ghGdB7swfyKiHKLvfzWJuPkitg
haYHMGhLWrfb1iitpOzfgzogxxIDNHVKWt9HR12Z0hIZceEE0d5pKXSgv9z5WYYI
wM6Gh/1xOWKqtGcBWPhBHp37mkmVm0xfL731dYDJ/op08fNkTCHwMj4vEa9iuMuI
r0cz2DbIQuUT0Zt+04PVf/0n832To+MWjDir1PGcC70Hse4U7n9AQIn0rQ0DTyzz
GePmDyN7W3+zhHl5BD6c89zHqKplPFzJhPeaKQy28XUoXEWG5WDLGUtH84M3dn+7
K19A7aJDDnWL1jPYCb5kyhgeEZAtSH684RzmmLp9UGpIqg6c5GZonCT7AKd1JP5Y
BHpeXSpWqgIec5X78v0xs4NyN/4QKg+rE9SFxdKCST5ShcHcrfOZU2s9OG1Mahc2
PpAEgErs0DklSl0/o2puGpnttHzDDEAbOKDbiQrq1lJhLxLNmGwT3A8wuWqZ8vzw
em2pB6ZfxmiaQ/oY/HBk3bDLPJpSn7Il0LjcsjB7h06qrRu5C3xW0CZXGXFbJRKZ
l5jRuzW4VbyhbZiGmqeREwknsY6Z5iT6kka4q5ZvE2VSaZoZ/PaFYlfkZK5Mhvpd
GiY4H1W548mPsroZA0/aqVw8kOF9Xu06k1mP35Ct14aaIKZGEe0SCET6Mpz7liKp
QAD9l1FSvWqETrbln+PflEdfGMANVi+N78zGC3kj0QQnC5gHzKJqvaE7ZSqcS8ks
lmRnlBOx0fESxdfgfhDkXhqL/d12jsusQIS/PmTiLMIc5XKXIUPQsC9azrI16+T8
OKv3JHevDHxGU5oAWWoW+r3sipI+uDZ7FjKIgUsMLkTvBns9pDYagQyuVt4DFAGg
fXed8odUUfzE59emoslCFhGWSULuo67xq1132STmAycugpO5vkVTB9Fk9buOIqk5
old4z6XbQ5nT/0D2WSZKhztDVh5tjhECSybWq6LzmycDvep2ds1u6IqmkN8v6lq1
RXLA0XATaL2i9qOw3CFd/SsHw33qAHaf6iffOgUIgN4+LCNYoZI88Kdi+Oy0aNT5
F3oDTxMfoPy/foFh9s8+vVk62IwUV/JwZdFYGyYWROyV4N64WU1Yzdj/3EfzQHd3
v9bNhHX9bjCLKPpb0bIeVokL9IGkdBUgfaka0ylhKcgzdxHlBFLL7+hUsPQz26cx
asfQDLd1g1DC2nnuVOS+TMqFojitFNPxZ/HnP7PBRtTYuCLwNMockt5f2rdoqaoB
q0IJrFDxW91sk9iCZz4luIAya0H/kPEdNDiLQEjA+9q6nptKeU1MZevde9kYGNaE
x43J9xWqJ5Eblg4tu6O2UHQrirbj2OdBB+X+5sDMunCXnx9S0Uz9TedHk9+/v/Q7
mJjFPwqr7Q403U3b8dqBeXBKaZ/bhk9HgcvaGC2yZln4jWwGp4zKruanSWUOXiY9
VY0+uZ6jFfoeIOc/sO4TBrTOgjykFMv6GlTWjaY0ETlYtEP6G4eBRbi0G6k63C8V
KNy3/57okkXKbNBD2GkDd8xrcYUpAqW/p6QnGXKJOO+yZY0he9hdwN5FacNghGPt
vz9S4m5j+fOetM0ZsjDb+THcDpgyY73MR5dW1Dc8Kos9nlkPivwMtiktHgW9hyg7
VhGV/lmLf/tVm64efin5cws4RWW2xxyQi0gUSirKMxy0rEGO8aM+Sp0Q0qQ5pwJ8
t0lbaUGReKbzhf4/WNleImJ6DWASXYOwkbh2EtdTMuX557IrfYbgEfvo3FbG0y0l
lexgL+skvEi2SrprRbT1rrP/MzrQ4ZlrULS9lFIYDc0sRTwiaZ/cKiytT0YEn7nS
ftNHwAV1a9FJ2a+nOuyVNEaYf8ijhOal1AEFjXaX4haqpptjvFWab0zrLpagUW2x
9+TNxdMboksUbkNTe1UgGomizGbGdKT9PVV4CFWAraGyKuxr4MtgbuEDFKYdIEXW
+Hh5xIyFNR05+XRTf0Tp9443dfCJ7+oz2fk5MnaaDw+HReq5c+P+/yi2UVUzC7mV
lQo0mQzipEF+aTQFUQDZNwsw7di3hpdH4rBr0fknxfBmFS/hYilcTgX7jCV7DRsY
+YVFS5JAXaRzBdviqyZQvFOHfwTz46dB8vQMZxhfbHjXrv2w7mfUYkFIlmhLCTZn
WQ8SoFlAdgIsCnTwS9NvC034jXPJP+URwJ/hVH/JJjFv/fK7pIsXg+yxgk9m7979
0kDQqo5bXhsP1xKs9Sxc0YfYqxXBMsR0EuBnrtNlkrImM57DXV9vgp8e7L4ZIl8L
drgaQ8CRgCHuY2by7JhFI32ZNxNygDEwnv03IMqd+GW53jpzqSRWmSFp0mOsAu69
vaaeOQcJN7VdN+InmVdJn8iUZjnzrdRGaA66SO+eDz6zOTfxClNxNLcKhwP6XJvx
aglQWv36RXUHEAxb+w4jf7372g+mZBMNR39dOwDSDp/0nEwsvMPmLEca6N7NQdvB
HVbaACDzp+OZPl9MA9UEHixnp0+3Jb2Sk/S+dkC1KO+XVF9SORh8SKuwmNDZz4b1
LzIk/ubssz86K4zSWrdK7s3CQmp4NyCuzC1rHhx+tEY7pLrSbYApo7SYcxjufthF
Xrlf8lyenmy7HUt2MXSzDGrAKdXVVm4BNitGGXM+MUi7dXWxBhAuV5fc9rVa+zHL
FMvZE45pwAG6gK84fXiLh9fEV+f0c3MSzIVSxlaBp7xIwp63oSaOL2LmhINn9ESA
Y+HMdP6ROpF2IRhqrZL46uoa4xcu9ONc5mUSiUwEPwktPPpQMfruFPOoL5bBhC8q
lZAmolG8eEJLAvzbe+e6u8/Qwy4AxMpdTiGdxEa4egr8oQAm5rSLrKvhY/xS4oDb
rJLiBNoBYil4r5I34kUYdU+D/6Yv915N1BCVSmubjM+4dBtBE/czBQYSx8DNHgUT
4HiuYHC5w3yViAIUiNQpKew322HlOm7Y2J6MnpPkx3Dg4at8aOLvCf6D2QhanyRz
Mq4BEOJ7fLjyOT5OlUw7TJUMpi3vIdLdx+MaAuul4vECIQlh7t8CgOFwNoDP3Efx
lkvnvilxXZZlkbnec7Z2lnLUBvkM1kGdiFSWWrfvOnW9m6HzWRNg9W/MqzZK7Xsi
EzOTU9vzShVuPvQaYkMeAgsx25OzFAKWeuzgCoRc8QYLiEpf+lIWdIbqidU4NsOM
cFDZ8Xg5o4SgJprNru1/rKfdNypg2/+Hdwgs1sjhl9Qeo+r8HoiPxfULZ4nTu9uX
FHTn5QbaD/n8UZzrJRgkvwILDO2+5OHtMkIQHeXMAvSLXM5EMWVxrIzOtw4qptpe
A4yXq0BMMvjaF4I4pc6LKDh0dDYzwEAu7WVE2v9Janpy+mzSNzicD+Onlb5l0CXC
3RclpzIkFy0yCfJP0E+UySa6cMoWfC5swLavgH54JroYryPnmqGFtimkr52V/PzW
iP9Mhhl/F8ID8CVyRgYGTVNl1C+0v4SSmRkiUmdhvAIxoxfk+LqlvVzaZTUKiUJr
gSuww6lN3FABxsWzBYKP5vadAfT3j08zIiktzrXSXOdZNHnEJ+ssU4ruiVPTOZUu
y2Lm8jTA9tdh8Yh5KgE0TzlVEX/0o3JNo5Y+DXM36Fbn50A/diSUT5S3IipnGg2l
ASGlSKZxYdgHY1vQFbW0fn+lp6tU4mB8UkTraAC+2/3sPsoYuzLfVXed5k0qvQI3
sraqB7STHyzWN9tXQqkT3qx+KwM/Edj6imlYH+kFkxcXXXTGa/nlSG8SJUPbEJ5G
4XKstdPDZgXkQAQBagXv7/AP9oSxDilmDl8BDPsyet5MUKxV27rCDbEcjXvUpXxt
QW2KNKdVs2ccdA59Ddxk2Rkat+zNKflzqRxTDi6Lt+pLHOOBzzAoZ3eBfMP5Unk4
ufhqQayyNHaRAjV+3KgyhDG82+EDo7ctx6gTkCiw/vVnw7bfrTQN+YtQWRI454s3
dYJ81NYxihQ5ozyd3lMxQRhATR9BDLh2K9B9hgyNRZz6Ia62T/iqibOFM811ARpK
CD0V892K/emjAVuTQluu1OboluqLHiHz0XFMpAIIhTZPgdeoZHvpUmefinYBeslg
aVJzn0VD4Hbg1gYl31x2St+x42BczQeMmCq8rfMX9/NdGVQ7bAXBXY1DvsoBYJWW
XXYmbtYOtKL6WptMqx3obJBPRFB/wot8nR0T9TvNzK9NXrkmGpPljhx5YhmMp13a
QETEC9mILFtYn7gvAfZQPxW+dTR6bC/iYjUOG4TBt4TPmeYj2Rh83BWlEScqseoT
XKtzPRCstJVWJjL58mpq6JUTB2/a5mpzD6G2yzZj9rEGGZ5/s5ZIC6InMVenV34A
H7C4f/OTtdLQwcIZx0GWcJXSaAzrYDP+w+SUCx5yUJ6yzSuaV8hhHxe3goC6E5zD
vL1HVrqcBelhbQizIQAtiUgv9vcfGgTXW0OhaFTzrjUAkalYXz3GdEu/wXHp/Hz7
UjeNRXZ+69Dtu0F+Lw0gyWckeX1vQIYY/sc/i/eOas46+XigI56OUbtvuewHk1g1
Ca99fZGIT1oafEQwVmpWMFipt0ndS8tzjo5MBrqoxr4R6bwR2Ajs5V34tZE7HJ1P
BJaR7HS4wlF7bI3zticOYeGUQYWB/czCMyYQXYzTP0LqmkZnOp36Zf/g8Vgg8jYG
4/mTfNhU29AZqbroauH6VW7yKDx1sW09jQ6OJzGWN8ciu1lrrh7SQ/ETh/BVdCWW
aQZ+VCesOrr7MBEnAG5tfglppgSwxnESzSU+E1VN7fNIEoC0deqvKDT2FNUzbXmC
7nn7IkQEpT2X9V5RqiMqPb9Bt/hPDmcvSG8DKFPbNYLNgNYdhKskV9/wat3PvONE
K0E6tpKoJcz/Zdv5d9R/FxGrKAi2ffP/+lZfxSOTt8dKGZQPxpq+3si2pwz+ZjYd
b/LpNQ0/zF43u2eOQQRkLxxsaKo23wnwpfrfinQsG92rzWmuJAkazohVV970ibMI
bXrnFHnnLKaepQ6V0NA9A6eTXfWukyAmgf3fGDjLm0W5XvE4rx8rlsGLq6uS8+ZP
Q2g95uA9VdJXUcj3E/mM7FgQ7jMW94+X3S8g0xCJKAlEWK+BWunVcz3nuOZ19dkp
hCs/G2uRxe0INQSjxY2G/q+RUUHTdc6cQHWgELsasv4M5C9nWm+6tYkaY2zLW4R7
jLRB/0c+eOtgwHOAJ9LWYz418PVW9YmOv2cT/6utLsxALtoEpKET00oEnub65Gq1
pPODPTsZ45yEYkaohA6N4PzWDS5wpZnESsiIWUU1CVBGuht44UX1pcuvVdtP6zhI
z35Zlh+vWn3zSn+hTrWWrgHHfDTOHBihB8MHxpSLJMezhNyL+pIC2qI1h4+Qyc85
jL4oNbGEHXouIF9nHRA5oevlfQIggz57v64RbtivUCwAfxZHku4ED+dvbFMWeizP
6pSQVqUUkZYJDxgitgobKn8uQfQporrfzasoOh4J8udOAnQR74BiMXYA0dwkH3uj
8TxbSS1l1i91HMkB2qJ0JhsVUzF/IfTXVoOySrFtU5quu6J70H1rS0aNDKXGqiV5
MlJgpbk5MBUuX6bsOD/49nKazSMlS5LSCmyzpOkuDRt7wNmb3vw+HDOFeQrANlpU
Y8BfyiZPolWIkvatGL1c6WQeSp4MmRi3Mp7d3XfGNeHejhvbGOxdTJP6338A9FEM
jO1eDljwDF9/WsfJZdAjWJNAplE6giQ3FyTY8deC/hSM7GIShQM5VgxUrvTsufLw
dPrEoh//YVq61eaJen78v/7eAuAzl9/uzTAvRRuQSLa1tCdm3ozPUqbU9VNb4dDY
BJODQaNvUSFj2mkuyRTqF3y7PdAi6Hf7SPHgDylCgcoAd4miIZ3O/PJ9Vtbw5jJJ
i1LCO6NgBZdwqcO1ewoxBfEKD4J5I7dITud9K5q3ZAYifu4/g8gJFbG8Wjm/QI3o
jdH2EL9o6/4NhH7ku4Qq5WrpGmLIVbyYgi/gzEt+EP6Cx1g0TEegJi7SaF3EFVMy
Xu34P1mpONKGaj56NEJ264djSQ07g7eASctVGEoFwmix6cVntnr9NivX/0xFKjTA
IPoPSfVc4T/SiBRrM0yBFIwM9cYiJxQjvR24V5/0FUne8+o9dJ0517P4UXI2BfYR
ZB9lMwDD27c/V6QVPjkjqZMQAOoEqwBcXrAs4zF0HGsdw6VsBPIWRgeeHoxV09vy
F7X7CSeIlDOwFHiwNLhHRoyhz/7G2dxnysi387H0op2Ajg1hWc+a2ZNFplyjKyA7
GxwK1ZVV5X74rTxxh3hT/FWBH/wIwBFwv6hSag5oDhqFEaP06+C/JBUd5XvuFYX7
bcsUEx6+MVc9l8TOJULXEANwQfogdWjQG4w3bGgqJ+ggJMsrUFmmMOsiMTvUeedo
8omD2k8okAgdSlB5YjTWQR5UiSaSZpokC/JbWfQibtvOqJUngrA1l8/V3cwShuf5
1SwH/X2Jf7fQ3Lk6PoUAFXH0cAB7JOML27h/BUfsOkbv7UV14SuHqSHn/sfwBSRx
ERQHUNQqQltdU59x3n8PJORyb9u5UI4aFcwj5avpM0cx1z/5rKzSidl8G9PWSr6o
cURVUGxbqd6llGtZCKGt8nDYxrqbMkfjLBm7Xk3ozNsr2K9AZzDPgCi8ATgx+7OA
lT//2bfpJgwYwxaZxSIfzdunafPLxWps4nITtGxuvSnj5V09Nv2+5iMDdgHrFya1
fdETViTEUX1jhucK+kQoLGpPu2PZubSeIFr0cL3MhiMufntxvRJOdse23t1mmfLh
9me8vHQultf/W3Wko+YIW23LuqCJcJJGtQQ0jPPW0kO52SeP6YfmbGqzuG/oczGS
1lFuTdK5wEYOU8gmkp/C5CBetx1UXUclWqLsa5xV/Jtf+2eTVe9NIV5dgen27tas
WTdpJzD/1FkPw4ShpYGwzwcF5D9YICRUkCSIZI2jXEou75SaCaUU2m9ya068zjSy
RqhWrJ+9Ik2g4uEN2TcmNNG4czSY0NK4e030YN09BPRigT6AaL9KuSjTY8rnR4wm
G5HP2HbLm2NjtwSt9fTX/BEJvSQH3MDyNSX88fRLXhvwqUktZe4vIOVKyFBF6JiE
KIpOes5mLfbcZxacOUgJPIctxrtyWQyUYzPgME5Vk2G0wHwhdErTfsqMH3hxvEt7
zYr6kJTcX7MMVfH/hHZBxaME9L2WKkOaDvVl01h+3kPhkLUZmmKbrs45YpM2dGro
8ar5fKusNeHi22qK2d2E+hfp2+DYR0CoFV3FMQCXxkWU4hv/M0+/9cx2ta6+Bpx7
eZg+Q3HVk30vXGDXTtUhnHSTb6q6eYfI1lVYz/YFiPSiBIJhMCrZ5lz0XEvEtktq
yRxhfeYnhUNb67LzDIrvsqYq1conPcOnHS2ffydx5W1jkYihmUZlklOxNDT/TbwM
m76HAhHv4WT4obIYMQKFeVO7iiP1RrJh6wSoWcL/pgCDUJwUbpx5adgwwMAtOd/H
BRyGV/Eql2/nOOWpPjFtUwH4MhBOCMUXueIp3WrGuvC4nKQMo+94TLpNini49+vn
ClzL7seovzdPVfhPw3WaIDIGc+7XA4NiFEERFMmW9QZhydva1mK/bfJOYnUFVsLU
Ss6GcT6COQ/Z7h6gIgopj10wIrBapW8+4FCCK2pcU1D85y8LxWzRRv7gxw65g/F1
+Sr7TfFETI6MQFRIdo1ohkRHIFNDjJWF2G5pkOc36B1pZbyvnqw5QgJYNqDu8ZQl
TQrA4Kw6jKYlKRbCxbtI+NfXANIZgQwCET1FPntUhi2SiYHfhncN2ltpcXJA6z/+
zizzR6hhqr7HFi0PhF7ICc/DoP3JxZRKSWoe9IIR6zaG9vbRo1gmsEVjSs+ZDxyk
disYaBbiNROgpTtv9L8hE0QrpXeKKXku+cZqo08TnTDh/DzOqvf4ycH6FI6jB6Rc
2stXlgHLxwHnSGhg/HW7G/pHnSP5Z5A4tdxhM/asCsjziDhdjunOS5PLEMmjITYK
9Ji28qvC5u3CZmxcG4Mm7A5a/WabR5G+6hBvTTkkDgOf+IjzAIB2371RTORkryY4
W2cXX9hKBPmgn5FW4L6qOT1YDmN5tgHdmKroPUwYm27B1pA9aUyPBkvqrMYpIz2D
loOtN2A/BqtacI8UcxQyZ+ZBLw7+XsD5voFEZsRcAlXfjt8pHKz+I5D1fCOlq7UR
FYGjyzgfCoMo1mpLFjkB7dWz7Y05LiRnr8+OE7B29dgP3MpSTPc8UH7EqrV79ati
DVLAciJ6bP9woEJB+psMQ1vV1ghoPRFzpZe/Jlr5yfOq/ZgPuVY0rYEyhsLEXrNr
7aME5wQgn8VVb/XPRaGtOggxACtQcFDcRrGqdUplD1xUa46cdtg03F+emPhx0yBs
5mdVtznk2zlRT/8U6NdgUwt/fzIqqmOluttsoJREAo4PMtW3nU5u+Ql/XT6RdFt+
XMFmbOSfaw9zHtStYHAXxmPSE0EWCfCoAlmIjJaAQPZJP8bkEpfTH/VsystAA6T7
L0saH+f/bOBTJyivt1XjR1PixmE+aSWT28Lr4hJcUnXdirt7m/Rh1jxR4NN+9wln
OR9ZPy9Pat6Y4P4Whm7w83cGDsS9al8SqYWH6a5bsq9QQsmSSKh7M4tEANLazHgY
RsoW73alh3amkYtkyt4aA4qSnqyp41XzCgClRjYUeBB410kHkOpPYijhUCPY572G
8VzFftha0m8C/VbxR5p5TIPUW44B5z0IpJ+pOzi3MlcypIrWmJYl232VaNuR2zkh
PmH91Ij2XHcUJU3WMWTKL3JifeQW450DkdbQFHTUa0wxAth565ANey3Z0zWSfdZa
dPMumOPFVToY8i+ZJq05Ft0SQU+952BBVyxI4xKjlMIxjqCT48veax5x1Ih5nLPo
qlGJ9R4CgZpltpuv0L7w4CTwJYKPmFHRW6zRAMAJm4jwgKyf6cpVAoXKFXLWGfBu
0Lx/W0aozPH3dwU1XUEV0sz66+Op3crY4H7QT+X4zZ0y4fWEccFeSkahL3xi+NMJ
8ye1PLFYT97Pya3LHvF1bNzBooMPoBGTDcrC7TN8pGdrkJyAb/EN0fWrrlDODdl3
ZIjNmoqgXxqUmYyUgIUDDPtEL0dDSGUd4DwbMs2GKjpn0iG3JH2pIbEgg10nTwbO
x5T7X3zJIzRvtigBbwUACcUcGbox0Kt+0weVgB1d1kJa9jQFu9ZxjWY1SFJGEMQI
mJmDV5P34PwMaPZ/+8JIHjgzH87OTZkm8FJHjeAWnMbrGk8eMblUtYTutKlmQRwX
tsMl2xyq24bSETsqUcFVB8rGHJcNnwe2TVAy30dAFrIzfKh+rvrI2OdJShT32PmK
H1q44LWsXhmEFeQvH8rKFhRU3AteKq1sw74mvZB6orL9HlgHZR5DFy+X+XuemAuF
EKnaeKLzRVgWmQ48hU9mcw5kBAmExQJdd+ralxPUDgG/06mpvEVA4E612Mgz2Sq9
pQdGnaZlvIJ2rSKPyByobCtVKEcw547AeXiN+xfuACJM7w70g8B4wjt9eSgNgQLl
dmbWltwPg5xM1k5VismCOh1RjdX+36YaMDzcMUGyD+7eGkUxrevrlBk7llPTmObo
FXyZCI5Ct307xJW5APqsaFf7wb8PimOw+3S6HdU9FiArNwsHeu1r8lX6bBoU3OlD
3Y3UtdPMpEV2SiiM1I7L3C6mJPPKg9Gk9l4f1PCQJnReTxykMTXfDJK+GSxYn+Sy
5j5nUYBIqYxV+egtiimJ74/0GH2BAjbyEwLctojiSvZf39jBykgEpY12OljyxL1Q
wd3vEr5nMsPIlzqm2HW3GnAtDYGKW3dhT0QujSQvUXHDqAhsjUa4WwqicNswRi1Y
KztusCpuuNo5CNehsMKMPEvd4JwXLirc4wBJGxZgzVfYvnT/gAggvGfKGfe1/ORl
54eoRaU5yLQ2ZcdIT3PxAwTmYIIYXKOMo5pLQKN0WYDGMG/f1sVSbF/vOLA3ymwW
apC2H8z0L+RW6VzoGsPhCPe5VM8xjkGYH2emO/nxfCWLrySyME4aPDR2JRK0sgBL
22F7JBOMlymJDjHoN4UKZ4wQufzOfx7OVUT0I80C6BIUxemaPGGx1cUZ1ro+8jU9
EpRs231lv+vl2bJ4Yl/iePauex2m13dSWW4q8P/B8rO5tqqJr5xYEKLq/uKBLaj6
eAu+1r9NH+yTgY7YL7swFYVTyz6sg6qXlw7/AardYxl4LzfbkK7d9VPxghzvlOdo
qkwbAhuiVtU/Bnl/t0oMb3D6uq3cVQ2w8kqVtWQY0SB+yzSBFjo2uWRIz919woQp
+AZ92zY1qcoW0+8xz5ZwssLfqF+AOcFJXFutV3n1HvC2K3YC6D8/j7Apc1tZhAT2
WffxBWO2bcwjnUSP+MiZXuBdDOhhjR8FIxKEf+F89uGeXGmfKNcugdyjQYooMK2a
RTWBUdkAm+nw8P2AaphHOeNj8unOozuMLw+5/aTblGdAYbESuK2j1v/fE23AT1Op
OGGU/4uGfw2IiDWoIU2VI8BgdlgIyoxbHJKdWTPTGjNAcniL8ZX1wVnLNzTJwuSA
s7Aq6iudrS6QVQxOW3oc5LFDWc+KLJ28ycNJN20cu5sVS7OpoKs56evoQKgx9Vxz
QbUcS2drQtEx7YHk0fzbAHXtY4kpnt4BSKdhC3NKYR8TnTWJgdxsS/zez0IMp4fN
18lBGlpF+H3Oic1kH4Xv0doU8N2/wIh2h85SrmZff/Vx91slq048rqRjuVekcKI6
xpnPSvvVmyyOAF5hxuVSoaSDLpv8pHHdIY2V52EPrzJvhWuFY++jn+IipDqsFdut
zmqcekL60aU1s0kgctoF5GQafjx9MHhj3SE2WQdiA3S3yrBoYEHXRNCUnQ1aS0Ip
2+CNFWa/vEWqORvdPUzushFx8fj7m7d742yz5JQVaxulQxCN1gMSCKTlkC1Vh8GE
38rJIcNr1hgLQfSRij/QOXIpBhLZ8xDRL4nyogtHFdBDykrAXfcPciRTnQEr0qdV
tTqeSTjBjP1Rf7jJO1nrZZFUrOp4Z3wGPTOqEchYqRl/KK4TitbQrbjk1H0pU+XW
QaWU2mKhDwI2lyXkuCHzgSJXmfnNE2mQtdovrczvQIFlEVpOYyDD4Si2vTtHkPoB
VaIm/Nh7Q7uT1l5C/AtC8AHwc0b4DCJ1kfH8q1/NKHP5o1GV+0ApwGdyLDg3zMpc
AWj+uW23VQ2/+lzrwM1ZCbrOoOIjYVZTzxVeEejSLdFLauqGVIuJzRClERd7RFRX
hDy4LvtvBKeSmnoicQo0xY4/Ww8ojiMnQw6jP9HZmOYE3kaWlcPREr2IHIor+bv9
VQDl4mH/E4X38qz7s2mZzn59yeZUcOMVCvfzKSo7uj2nYjOvizFICPA4Qye9QrhM
lrMoUJ+ROqPLcz+Q16DcIn9Og5tJjkDSHyARWzvUBsPddMVctMQHsmjokEGwFi7A
LZFwwM3/YMeuqG5h8i35RJ9QC9r93IcgmWlSyHF6WmnHRJJT2KQvfELgV740xRx8
hWr3fdYmX1eY9MyksfhaeRHlHrhXElDuwz/iP2WLRMqi8vI9FPo7KsJLVuVYTN08
3gKPKZWgTJZVuZ6Xucy5uAG4ZgFyH3WU+vhPOiuIUd7Aj6Mm9id50+AO+ZGWLFAH
ZY/0p7340N2ZVBt6laQNYgqGSpuXSY1bCvmHG+7H64K/g8HHU6R9Muo9sHbUhodH
`pragma protect end_protected
