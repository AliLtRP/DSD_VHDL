// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:38:23 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
mhJdKxoTEPvfW0Vt5HxqAiPvMe5NSaI7rVRWzIfFNNeRrdw5Z7Q2Aym0QS9mCafn
T8NL4rQBsr3LO1fNJUW+HXynPOflT3aCUTMuhII4xJrQbGz/Ni0HyyhteuOZqm5X
6n0u2S0oswh1QteZDEs6LJvhOTcQjxUP64MEb5AYYZU=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 7648)
P6gRug5WWW6glKOr7IKlIpsmsZUIRAb7psr9yciuyuH1SovaD5+yYtnuDj8ujot6
CY/fHpkjNIS5megCmXOTicgezK4QsFLUy7qXvRsYMoMWh3F04r0KaX4E9NlnHdLh
CqOm5BfgGWUqf7r3/xjcvePhAkgkyMnZzBB/lvqu/i6HLXKUo68I4faPXmuEX9Jl
uoHTQdt+SgeFxQCj20jUnAvaSXWcxQgB74FhaU3NEENJ4wvGRedUjSfbn5lMPgMX
6+PF+wUfln4RDtEG0YI0LCRZrDT3dzf4U4FjmrxQ8udIq5hWt9iGz40Fn+NMp359
7q2g8Hz6Q/SG9uVuKluBITb5bTpZmhZttLX1B3/bV16P7WYgcjaEdGtkHWPZ40QR
D0vafhXtll74ypGSsx96JDS3u/NmXTf60/mwmdIpvmn7cNwQ5xFE7UROgXKGMVDv
d62NAKgVyJZysO6+swc0iR9uxTjmqXrBiYElHymaLlTM0i7MJo7ghirzk4/BEJIx
8BOz6dsfDhgTCy7LmeF9C4/8hhcx0w5vb8v7YRJZABPT/JfiUmHrZcb29zG1N9DC
Yvoj3gaBEHeV1Xku+Wv1tGC5FVbvTYm3/pWfBPxNRR/7IWz22jw2mckTdQqI2vn9
H7MNqPkpmOiEqh1lKJk30bx5Iqe0yYIIZIBNvoCSSJeHxPWVDHgDm4bprJ/7xLPT
zrCsI0GNZuqZNUac9viieJy14syYKlLahsDxJriNX0pa01pimJw5uFruPYO2iVmw
/HwO82DZLqUYyT6nrzPbeRtsv1Adbx45K7NRNzfbwWQdCS0Mxpnv3keaOQ05lkWh
sSpclSgznabQNXOh4lNa0+R+WZZvh5HqlD9pmt/qtJm9VESVDeYTb4gRaWjFpLvn
gzw+hVAq5ZrptFwwQo3Nea3I+zQEJSEioYUziuq1cRkIC5NuvI3KfV4krUb6GeeX
W3f03yYHPM3D8Yu5OiyaCrItt+/NN9nNZNW054Jy2ZByrFrIBTPsdy96j23d1Oyq
/4h/LETBggbyWT/+Wb8JKoDRlIV8As63TnyCE2ZlVM0OnzTOjnb1ePINCdzjS+ek
SRZY0LoyaD7ULenH1RyIESxZ2h2KZdMdkSFJ8iKus6J11sBVh12NRYSguDSMWl5d
rjTbvJ6JHmqIkvqrIRyIXCUrii3SEc4Eg9mMp4SvjKGMfqSnz7vJSEZ/tCMoTUVF
3gibYM/ARsQq6jrwIynrwOdcnmbCCmfOn4sLGMH9qbhnfsKybyqmuhy6cqxdQJlI
3/7x/QD9+oa0LST7vbJ3TsacEnelFhVZRzGyrsapeEXBetKiMWcGZYFpXrXv0S3O
m8Kwu9BeMhfQ/7izUVN+K2fvLePdur3DaKWZ4F4toTUSSQaZ2QpDY8mgHamFI5sB
QWQTSZFWl0o4pBiw93LMzWMJRPIAQQZbq+/kFX9St5ORIhHxvgi7ei+9YNm+Q2QR
I0NSrObiuJq6STMcKZsqqyNRZpA6yy35iQ9bFpRTIMIyCgDUKugZ3qlGQUTPj8e+
zcpQEPkj07FJU+QFjiadJn+IY/wY05Zgp83CdRWmdjSriuLm+rcJ5vs6F6poe9XU
XqjvTlNFwLy/Zve64umRA1p+Nh9ur9Y68/GNEvj4Na9lvG0vixJTrguUcHlmJ+3G
lXD1vZkN6kPazA6PrDoYhFnUqeTTdvSWNd3Pod0UbKs9fKXwo1kRxML/va8ii+XJ
Wnu/sEGBkGLSVzgKSVEON95Cf4YnROcLzoXm42Df8KmH+fKX5KKwnp9K8J0r/jPZ
28fBr+3QQSjR16NeYtTwajFN91AroiPIc4Lrx/fIqkVnMx150XhbpzmGrlRtqRx2
m2ekoUULXOZzrIXEI0YSkQb0gNHSKliwq2SJ5O1gHmWW/v1riMU+4HmV7KL5Z5yV
JR3yRcju5NZevrOOQRfDp5W+RtdFVluQkl59PN4yxZK5Fq/nX6sXBq7WPGjLXYDo
TOQWFESQwzAz2ziH/FA+Y3Lem3YcDf/J+CLb8nNBrS53sTRRk29y/K7YzE8gKL2Q
vfuP+zokr85AfFLY13B+5rCDNYq5JxIeDPJIIERZUjdxmYUNF1DbLdtvACaw/KEC
H4nkBy08ylRBfYEi1smzYf37l8YkpcFXLovJeF9T3CoopByIkIxeEYGz6efyrS+q
/J638GjYhyV4dxv8wP4DO8waT4bUVKqdGnNc5IQB3JnRU/Nl2faUmo4DuHn88BaF
bunhhcMr88cpbYqW1zbNPenVyvQQucJpbyTOmrD9XJNGdUPXoBd4T13McwyRkPnt
ZL87rjHKHBNOjOdxv6WteMYQlkkGArJxW3nJhLth6Mfrbfm2EYsDWekP5xoFHaEa
WMYrQHG1tcJP/j/EZEzGbVEOqMmY4WbwaNDyCY6ntLIM/IUp3THhtwFAD6waYjJJ
LgrHRQ3iKrxwawj4s/hhmIwGXo7+THmOXb4yRYTgkg0fgI4WDUzlhieVfptTGpz7
sPyvb5JIs+MtboF0C9zsM1GEdMvqwEGezUXf4riWfivtao392gLJD3297NzBANA7
+OJaH9VYBE4Oe59svV49b1W4g70Zc/QrnEZ15dy14h/Ia6t7A++3FrRDxs7nFy/3
nV95oTEKpXAbAWIX1C3JXIlnA1S2OvFdUwxEi+atN8v4qh8+KUHOfw9zEXY90eig
gJlfDQeOnqOCXkvtkhRgqVRoyKzWhqeAWg/Cb3ISScQwmfpiqLUMkqZbQD3/g+mJ
bwYumICG87kmGn1prv5r8tP1YQEkLxBIID6wIwRaoNk/kwFpdcWz5mF7/4gbcm1K
gpYGrxj0ufYZ5dgR5m34XJzxKVkLaPS2frnj0Xxk3o6LUYi/bLiTVFGmVcUz4Cgs
DeM4Q4EkGkRI7iJo42S2ps28e72sKJQhtZTZg6VgTFlAJ2OqaLRb3oX1cOY/TOsm
tbIsStTFEcb7FcL62VeZyZxdWZVYXqWy4gR8PuHppymqt5Ov7X+auMqLwbT+0F0i
ikC+qSOLN3hmbpsuQXhVn3a566n1cWrkwtmm+J3l5lUK1v4YGH2xnjg0TXlppU0h
/MKg7jlgEqA8yfgf/NqeYV5qUDIirK4CFKILXP6eT4e83aTqK4sxvb0QFk59Xs9I
Twb5w4IJTezKNFPmARs5761A4ib+ktSniOeaC7HPhUlAGABMJIAPrNeUc/L4qm88
kSEqMU2zS6c9/TuakgSRJIaJ74d3iTxa0yfIKThfg+ORtCA/SclxlBn8yc5oGXGt
05/I0J5hrzg6i08WZ4NlQip+mghnktq841Tt1nqoT0OoTYpLK3wA9tCbyyvAWt4q
SgHxyefNa0b55gNq2OrHP7A8L+dx8GFfYpmQlkzYdA/Q5IQAPuK5l0UQMGgPwX0S
86VeUZJhtTvXKafgj+C/YwiYazfWmd9jk3i+4wfLtpFUu+Kwv77HUOM59n4w/xd2
or2mO2GH+NjD/kupmlqQXWq/HXZSmqQpwrmQG8fwMW9ZIF531pzK6L1OPcv0DaQr
QW+Umqz6LNJi/5+HGelJ+dNkEwYj/u0lAUPOihpBXgsWO6Nu7nyegiQYNVcTD74j
h7lCM1AwBi1S4kvu4N6d86YIfT946trIhTRBS6tGYJwVpNl2dXFjgiSklQ+K6DQu
0OFgE0ubgQp3bwrPbjM3OuK98gpmfapi/fG7ruD7+i5TkA/3fwt6l8CwosR/of6R
wHcMp431RXAKT3T5cPdRCstSNJ8tzL6v/1DXkM8ifi7dyt4QrDDUY7KKYXhbcvb4
sizZnOQ1r2IzV63L8gAjwbWWJvwfYn1h0ucYVdDbMqWszQTLVX0HaQERe1leoroQ
hr9NZwlZ8cYCiA/eQEXoWuyGB9EhIIvOQg+/F49HiuHI+3dcJmilQ+dVAatfAOqc
/DM2oSHal+WIrucHqVITO2AMi2DLvLIiMDPa6L1xUVqVVDnt3UTdWyWHLA8X7I79
plF7V1gv9hoosBfDdAEThZdvn7qtFNbFDEdYh6wN806VI5xhjg2vQoSWmpaRaWA6
8XGHUKdZx/rynfKwxqLxXiFPucWgLetEAagrGXZu6WlkChtQBcq+bm+YE+m6bscn
N6URi7qA3KK6JiayB4HFTFn4VVOaU6dfOGuUDmFXaEhvy0BBuDfXERVQdrZyhVTg
FwrpYcaz7ldc88ncs15vhKtzPrmdOSg7TqOF+9FQ5IpZsTnw2Y6XjgYMeEGdLWJi
FT3ypeHq97Ni3m2lZ0dWPXiaT2RP2Fl768rSKoPx6gRfwfeOcwiYU5vLWdyJCffC
1kiQ2zdg5dwmhBwOSwFzihW7wEXugHWqepjm/G5CokszXnbJqZBKrAAhUREZzWWV
/zfzjn6zTx1IFayHXf8nan58w5LowiGd0AXMsPZFEh/jg7Dl+2nPD1FzvZ3Ne3B/
3gPOKE4dLeY7njQNgJ1MREzV/ZTvgqE/1v1OmzN5s2DRpq9EYHT0S0qlswko80In
f5muC97XQsLErFLQfXYgx3P85Ma/Yp8a7CclaEoa/FC70wVYXJJ6lvZKeMIMGGm5
VWrW9Qr8uLrsQKg0pGVCJUbmLnXnR4Lph6RBpncxhG4KQu5VBdCMMdE9KurWplXC
v6Wc+jKeseWZh5ddQcdgIVtin4wBIYinrergAJuU8sDSoQKQwHD/O3kulHzsjNCw
GaaKnDwAWB2tadpE7fMk8WvZ9lpOdJvgILARbBpAcFLcS512WS291pjcLaGb19r0
CmlYNqh5C4KaLRPONMVrjJWrBRaBO67po3WpRd784ejSnz/ewxXPkuOGHzOhUnkq
0h69oRa3mWZqW62JILDHjAkL7bjI8uRHSzHDcaYSjFqpHmCXO2uqRqEf+09FLFUY
uH1QedqE7+MCsLh8VdRsVK0+eSm0a+H496CgPRylMRCCX16Mo6994MlWaRAi8U+K
C6zeQEvA52tO6cN4QfJZbHjL5DcZMOiIocp0UjzdkzGESsASseBqoqGDTzwb7O6s
xj+NqC/vc/Sjf/wk0npjyY9O7FWXOvKGBwWXS0Bh7JywBUG5Q3wB+RgYN6QKpFVF
Yf8V/bE6CANiv6c61ZsES8k8eltx+u5jzlRV7HdAw8SbDsJi8N21NlWH1Tn/LlcB
1/eg4+xIBzo4sXlpLcnx9UN7XABWE8zub3hD0+JT36eTOAcJI/cvgrYl3HCp50ha
DKYLe/j2UOFNROJ5oIEFoEKj270sOQai5KkdmMgrXT7piBM9Dh623+6d1z+Mwyyu
ov01yVfzW71Mmo00LSgAGjhq86eNpqGtGFasZm898cx7gAUM5OsGxb5dfxf5Eio1
tcUVs09GG6Zl1CciTL5e/G3bZeenInTySrtLRw0KGjxLtrPxDpOFyusTG+IPm/1k
9n04kLnlx0itrvAseF95KsYHyGOPh78z6M9J6fKLA7vG4DFV5z7fSXijKDTeorzo
Ujcc2xVXaBcHcrSOWLD0tRfe4Qa/Qoqv3AG2ZzDt+378CxB56fAOep7/gvlLJ9jY
LmeJjTnOFFpWWjmW7UeGq8Gp3OJi36PyH0uRffS073JPYYMOfc3RZ3GdSqxagYed
gOBrnuyFL9NsL7BLZVtbZopfgYyKUJD2LMi3hxe5rjGdLPYiLLBNEFttti0nvQAK
uVR9KZ8NhC+FxIXCf3SjrCymycwaXoIBCSXFfQ4LoGQpxkLs5eZGQCXC0a06p+kQ
mtJsPB4E/eXXXJQeilOjeEIJuzX45eho3xthR2ChsFzeWh94EvMnr96jNvALQbgg
mDQkCWxhLT+te5hbxQkkAF2D7+9MGp9Td9JAXKGqcRnigXTa0jukOvFgF3HjIVnH
pQxO4Qs5CQYsN+VW16oZcy20kxID7N11eHtqgQP1/MMzOS0JolYNSbJ/vJq30rP9
HZyJFTPV64ehOPg29Ny5B5BG3fnbM7wnJHwPz/XJetXVY4AF9YLsK67vYA/NQHmG
6Kk3v/yRvYJkm8njy6bK1vtI7LhLnVkq/wnpyGQS/koQhGIWWZ5l3PthZ6PkAE9w
ojMkXDRU89qt0TscFfmL4po4ksZiTbfqP3Z062TGzOjBrP5PZkx1f/h7ttcJTfjk
cRGXvyB1gsl+tFbIKK3Cf4RMMNQz0etgtvebzd0cJodyYUtfseqxb1gqa4t+H/tZ
651QUZtlDR5ohzJouGP8gkEwtEtm4a+PXj758Y5B+FQzz0vPGj2ksLDcVWsV+qY5
wOYkcykXUDOsN2h1nQma0TOI4xun/WrwSr/BK3c62D37FoNPlC//Zg6U3gDyL3Xj
dsKduQsL9qpcBwDGcEBQ1EqZycqkBoktLTPt/2M8DkMtQxOjEryCCy32UOP8ijWG
fKQxxrMvrWj9VDoDIj1D5Jmg298uxGcqHYl7/iY7w+qspOVCrK4jfUPo+wOh9Yk0
0wt5FttzWAYuGqJppJhJXpprs/LKVqKt+0mQ6aksJDffUInGf0Fdyi/AluR4M/ET
jh1oHrxrSnk5jxtgFhzbJR2Jhmb3TZ08wqlXqzjMU31sjcoFcowtKy0ZHh0hUkKb
6b7xkBJJtxMDDb99jk4tOCw8Lm8JOMaCh5zLcMxuKoecFyfdU9L248WH08/9f+Nz
qKFYH9bRmTV0hU09fbf1Ai0f99ZEpEe2Ez0LH5ayKEhvG9HT065nH2/a44c4/2CR
PYdijUWHuwnAiRBtRXSjS00RTQKQhiDACRhzuoY0X8OPIvvzQFP+Rm2iFMpm55rm
4Yct34UiMU50po7KKdux4IRd2frhNnye2twEid1Qo3iQg3yGSHdeg9Jff0+1L2TM
ZcUaKTQe/n7NHdO3VQuM0vg/BzzqMyY7VlqpU7rL6H2dTQC2dBFD4q8cCJqu5EnN
Y+An7iSWIiONik8xYfp7Wn6saRFYP7lBCiO2IV86zOPB9rIljPCcO2mwL56BwWDo
1oUYILEbDWdEk6HCxbg86qDNNKs14raNXH7wHnRjlAT8kTtyy8vV7FlUrCwlS61e
GAxVt4XLDwcWTl6dXlPmeUM4mVZwicKUG3+IGFpxwGDtzNWHdHSGLdMsaiPwjdCp
xBE7/JaehBR6wQmFxlpZzhs4dScS5FEMis1QpR6nymEbWdcQseV5nLujFY15sfxZ
hNRlc/GmHR+QhSfpcppo9GXpbOOhFMcEryrVVN4OHmNkz5O9i+3mrAKCJsb0l4Ti
HYtHAG1hHYjxuRCUpGu9/eQrjN6CymPlLd+UmLcd1elT9bSU/1wjrIw0yGJPwEt1
DAswqEbTP+0r5v0sTu/klzX8qun/EpoCmaFH7TsuhC56qIKUTPaxB10dEt+Z9GCo
IvXpdttzrf3srSd+QlyyeMG5Jd0q8iMxf+wgjOx8QpQFWn88SYOAGXV0Qvxnagvv
9MIcPh8QhrI7kYV1MK/pG2AH8E8b9xa4GAV8loGAN+hJRfm/XQLuZHa7kxvIA/1L
wiy6kP3t+2K7C7KXM9olXKfg6SZzwdWr/FMjFcEDXPuPDOZ38w+p33JsVwZkwdc2
U0jsiqUyEk/ZSTd6kn4puS2U2KP24WJi6urVHoNTJLyaZgjhpMraVOy8AHz3AXNY
qQ1dN4+ZFtSlbEHKZVhSvJIF9N+MuqP3NV2PfQX7vanBLiMh4/UY/NOJFEZN/rrs
HDFX1Q4U4ZV88jZ4uJG8OtyINQP9+DLqQjPzw2I60vfhtKnoSbMspiUE5AJ/BG7R
Pw4bHiOB7RNmD8A5dsMofhjiJXhux/1dXS7mtydCAWeTXSjQKgjJ9p5ewDsD5Kxm
99K8+yq03WkLbpqZPnJJc9fp81xgCpuNuTIoBXVMgDPQRJIakyTG85eD+T+JbO0t
jvWubLw2aSMtT1NB/gZJy379wOU4+iWp5RSPy+M9RpEuB10kZ15IRwIrZzbw161w
Dtd85MOIFJ/uuwugc09Ay3b+YRO3Fx1t54/XgVOnck1+HceKv0jJHHypQTzR/mIx
2Q/sPS8h7zXuktCh17Gn1XzRdM4tWVBYy7kgr/DNIQ0DxAP/rLvjgUXtKqeSbcf9
ulJk8TojSotzCMui8Y5AaL6fQh9ZlVDUJpRvgv6z35dktHeUcTNGYMgtdw6XOJjH
ZA41H85ECMZ4+qEQlo80EYRhmQhDosnZExa5B+Asr/2LF9YJWlRCgIYKH2Q+AusN
XIIhLP30d6srE9uc8DQiOuX41jJFLOsuXdz15wtMSLYnjD4hOLajy7ugUssgBtcA
ErfdNUF47vN10AKRuDSYONJXSHmSkj6m1Modryg7eBHW2WoY4N2b5CNzWzRvQYFA
b9d+jgAJAKZWyNpmA5SErCsbuQ+jFZCp5kVjRvYJS0BopCM13SxU8kD190pEO7F6
rSiYLpGVr8p43I4DV+VQrpLuzo9q+bU7cSbOD96GrfGi4rEA6ezlHT5JaXqHPT2N
1efV1GUl5dPQfoKrsGRxGiajzOFGV7uaXVjS8x0edctlgax0LnSwraX4UNs3LYw9
wDncFLm0OinNRtGI0lxtKCa6KO/75tAvCCVbyVJDZnyoWk1KiuMbxy9GK6gYsJ7q
0ZK3CI5ATSMI95DwyA7uelps4kLnziTi0p4dSrdyk8UMrvp3GDA/KhMDLovjX86p
PrQbKFfGiXTYo9WiJeizIPtmfiRvMK9GBrsHrd2YFbSW50hHXqfTJLapWUh0Z4Hl
JwJwMWCAYfcabz9ZaiOokPoJCqHqheGGMI0pdAZHWiKRyVeD+mVHtxwNasN4XuCw
dAnA0wr2aWydZZDzV2qcQ85w7HBdo/Lk5kSw6V1QJl1Fia+iz8eh8prPeJlSfvo3
5dSDsabWOcBwsfKK0xdJzyI7c7hVyqbzhEQGruEfFwtt8R0Ret4wNkmWvgoElyl/
E0R9Po52meroNewkWlPMArGr3T7BmIbkBeh2yiMWClEJ8MKLZr/rQ08FiBNl+R4Z
0nfR9jy0A0VHE4CANveDyuMY0MHGj5vSpv6BdvBFgvYafQE/0oLFVZnbfBvL1qYP
YqSNTeKYHZECGSpISSJOmPaS2A/MNKMt9QR0juJ4OelUMcqzL+Eypf8HxWeCBjgD
9b9JfsJsgbBbclho7/7qOpZyG+Jf06o2PT8J1Ng9tdJhRCLSOGq6fUA9to8tBrve
O4ZBk6jHzStgbOiekH023IIdLdbiioIMnlXz498rw33/AqAQ3HKyFb+nl+fZCqaS
dVFEUdMQCWOatgFLQcvPD4RWnVMzA4wz+tNx89/90m0zecwkxkEpWYnGqcsP8qH2
XpM48p0513q0Ap0gpGJEPbdZ9T1l2tnbgb9a5ws6hzusnE+N+90immZk8CZZ61Qc
QbvAI/rGZvfj/DZtIYNsTlRgjsyyw6HqRvz4L9C7OhlqKyBYpKlAWgkBu24/FyNH
zjd+09EISkbp+SkfYbuTobrH4/qfln9uNyZyJ1c35XSvni0B753lexqsm0xjzGCq
Yp48OqXXMHTAW2kaMCoE86/SIvSqyjwlP4onUdbN+hMpeB+LHq6mc5mrTtGcnmUH
C9rPlzlpJLZqopbt29M8CYkd9kYkHoNyZmwxoEdWiQd9zrbAhpAnJbNtJPnDVFr+
oIV22Qor64fODFzRlvM4rkC1QxpvdDQjzTyNaSL+AuLTOMW/SyYUZgdXAdhY064C
gCAbc2nNIem+MiEjjHcZC/BOkFV23RzGRmd4G2Obr3g7by+OimyImMqlXgVgU0hA
qKLBDeTi8fbXYpclTxPtTfMXMYlZpeoHg3suLtYkXzbZ3nm/hzGm+muC2upWWUEh
j9YojVqK6KfqRP1GK4XY5hT5twJHfkVun90IuCHlljcX3tPaHhCtxct1U3GSq3Py
AD8qO+nN0dUyNDVjK2JFn5VBiH3sYQBqc5FXlv83dxWEGJ/S9TEK79flUj+y4dXt
O+3wlu1JyFOesC84ogtqHXDnypKKGExAgCHFwM9weAWMHmyAKbfG2R3HiSIMCf5R
1TeMO4pnCvOURkMI3p3pWoIlvN9RbTtUSNM1ik9zmJMLRop5BqCBY+dF8fo30uWj
ySPI2KyO56JWA+12D96B0ZPevB4aFLUas5c6WKzfDXtffaTlRBfbwCybfi4k49sM
Y5x2Pl/CzJLyes+zUyYo+B/2jK36S3v5reBwGrUi44DUFlnVlULTl42DlTR8l01D
0c39LLM4V6I/9p9NQn/QQn/+Sofkl0kVrHAmpxOjdNRxTWw46EKQt76eQWPl52EY
WP2Y/UVsP6zR99pcrKyuVA==
`pragma protect end_protected
