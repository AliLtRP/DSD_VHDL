// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:39 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
flI4Trl2UJ50mQcWIxQx60gwhgtLRIg0B7POc5xAsJe0+MKHzrYP8zgqbPJiELse
3d9eoV7964rHdGEaba/rXQ2hDLC2uBjDXoS7CpivdRWyVpI5jDeUO0niJ4UTn4IZ
Es6qZCK+oFEpGTMprGL/CWsPh5APfzqBUoemH2Gphmo=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 6336)
Rk4J1rmiTISE2U47fDYR16giZt246Yw3wSeeiRa5T5kxUmwL1wqJkYtupZnC8mZM
xrdHrYn6sb606ZvxNnofItW5520NSF8qF9psixnQQ5a4spJMHlIqf0mm+iYX7wNy
Fiz84RP0wWkJ9cwyb2TTmq2rYvJu44S7Lq3WoUZJ0UA0qAkDR2JWm188E3h2S6pD
23lmpZpnV92R0RNZzRlynKIFIXHY+ykvGcs1hAHQqKVtpNBWM5sPwVuImsGbD0hV
/m0QkHz+jINDGfgW8aIFpPkuJ2GEnKYDI2OC+bKdj+0fn0qaZSMDgbdI1YYwM6q1
o9omHHoHWOoIUXjjD2QDquw9FfuUR0NCcMPZ4OTZ9I/WgSblCs2KKeuq7hdNmyjS
/Z28OOL/D0nyRQ5Okbg7SEfusmPT+z7HqhPNu4RrRyIhQpXCcD4eJE40ABZdV65Y
b8zupqhYI+zS1SiueyBm69kTRJmg5I2NoLkoBEmDPbTs0xB2BoiebBODXYx77U/C
BlARSYKz+E2hoWp5sWldkmU5Yo9BmW/XoIli9UosMUqordGKbXMP4CiSAAbgGywD
eoYyssO4PXQt7yMXY7L2PMMQ8uw+uSkMr/WdLfWSv3qt8lLRDlrv29tIdqV5I7MV
Kp2KrVC6m81tHoRjluaRLMIOV9vbouXxATnHi8mNUKilBfkhQoJ1gBR3ZJoUfseC
S0ACU9JaG//Y7QBqc0WuHBZ9kVn8vxccu9gtZaYyfzVYW4HRIRdSov08al7BfKNx
5bS9P+4z9zpGXxdWLm/de16o3IEbS6f04pDIgjJcNgBTcG9nOa3PKKh8iVGZf2cs
Gv/JbCUAJDUpOUurhwricuQFXLF6LXL7Xy6jX/qScSgGSjDObe70qTyYbTxMV3M8
lWD2b4WleuNDSUI+hFOjpd/bXYo8JQF84ikoCMjrUcQ8kQ3AygkW/IV3Xpai6/xA
xlYXU58OTa2UrjFM3i4Gq3Nn/W9jTWdlZhwjy8NUFTv8H3DnaNvilP0sX59k0Rw4
D5DJSpq3XM35UOlAej5cXmZRvHiTa/pi8+YojZ3KkNreCguvu5ZjAbufp2mZucUt
Xcm42sRENkcWvOfWhtnR9Sot2WPHV5hrxEoxiDxKIESPDaVF04hRZk34QqdRkn1Z
vl6AM21AH3YPXCbemqbDHDsRKLygpHLXpmFREgEE8Bp7oYNuXZq2M80HPUFpq8P1
PjQMc4CNlp3pJQE8hjWeT6UvlGpCpZDPZGSRzl0b4SO6j50fK6Hl6a2AeeiiES/t
pRS87qhXRlX2mkTHCE4UBR6zCDuZ1nkrediJVGBb3sydZs4IhvYXoY6NY7fLsmWm
yn/GpAWM7fWZjah3/YRG78jZu57YhKcM9oRBKIc/zQuBQ2TxQFdipNlT+wEwrMg2
8B454z4Ch0exUVm/H3Fzb4HhZyrDp+3uSPLn8z4rfliznwN4F4smmEuJ73v3XXfY
jrCQFchY9YDFQuoclBD+OFAeSZ0olRgT6weHoJWjnsCki0wdoQZpHbS2LlJPWnd3
g62WEsH5e4vewm+RelCtXwPnuUOe1SpbY3BLN52lpt9HcVn6ZtLW9WuDrxo8rtp7
yNHMU8ljMymIJZjXVlMVgY0yZU+PHMRKc/BgnnJixUeq4DsJ/wiBObQ+FVm3B7bO
jmwxhyl6fRu5zxF3u0wOP2x5tGNEItJZR0xwZGdWX9xIuVoroSY2bgEXdGVPbSY5
VV9+xRqx43Crv2F2JtYPabZblEGy6180gLgmEMJ0AEEof2je5YGAuT+w+MVxClgF
TeEw13yDooqLvxJl1O85mSHQqUpT2xt4u/QrEcC6OgvwEmj9V2kaYcXEXaXuz1pu
NPqKVOeOZdvKupPnRDwEp7jrYL+vC8IWzhwvjUTNwf5ZEVYQRRCOKjbcZwgE+mSs
OUkMDvud0kAl9iOv7yH2MSX+D52YJg9tyBFT/niizrlzhOJ0oMPLbs2LklOsZFrI
XCdG8Hp6R1AX7JfuUtWImXhbip0Bp6SVWerJxumyvUjCUpZsvzKQeXchmG+XXZah
Q9V1BFid6DOmMRwzUrY7Jyu2h23Tuej5srid51O/Sd9OF8fY7K8omSwA6XbbCq5M
9ks4AMLO9up49HjMUUDAuPKjWxE2kP5WumOaZQpB4SYAsM8qzcT2k7YmagEg2CQB
hfVq4fi1QGKdMy+zPCZQbHRSHSWk+2rpkrXRzD3pcuKd4Wtfa7rDt9sBuDdE7/bP
lxjG+VgocZYnGUAgKfpbRrjjdE49sXciK7E7w4HGfJCe79b/YF4dKG4EhFJXVW8y
0GP1rjT8upWijWqPEGvVim1v5jJXR2GLs+zq45baMiK6MecYpx2vlvZMSug622s1
VExDpHam8YH9+IUATUO74lPAmss33ggfd8/3uMIXTp4ociU8ZiyZvtwQyuzoJTlv
S4IJm8fu1bm3QefuReIXVRBGESgu1eHqxap+PaNm2tg/03pqhlOGY1phFUp7+xI2
2JHHZfwWwiZf1ruKNDB27JUN38D17KQhrXwvORXc7zWZ0I34+bDHwNTIqACk6mKX
aA1M4urTZdmhoeVnsQMqd5rHTFfFjpanCrsoLFfQ5Ma9QSrNF4jbCfYphQZSfCCQ
jkcL4DiCGp5X1dZZkhWBi0m8At3pS7OVd2Z6DYkXbjn9OaB0a+gyxFpNQUjSE+2N
V/ZxmYJPA+2oDE5x4vVob01pE23PGV2rLfVFfdglHSxAYf8ozyiG+LuWO+VgPAqE
YJnmJQ4HnHIhzyIzRS1eOalk7ZAf0jVwMf+Vd/PW7Sq+IzdwWjmdVeCXgRHHElql
weIF4MeMzGZBQS7z3H5zT9dFViUhz/Xx49MxsjCPAoTsm6QkY1wKrP6Tm/jMTz/t
gEvqYF34KGaeKuHIac7wNWPrUpW2+9WjRENcPWtDXSfDezRQwRUgJVXqqkURpMd9
cXfA1TZCQl0815V5vu9oOXAazNpnjtrtmwU4pY3tVv53fsx6FuvQvnH26DhNxRf2
Zl4FeqpcPdEix6RO0E72gnPZDc89S2gG5Fih+g1hT8nxrqlPUuSiMXj6V3Qi53vE
QSzAnGuSX8CtC/io21jHH0O0jiuVByZQ47JuG48Zn3iaVTsUVfNSYnF1ronJV5AV
tAebI8qn+o8WPUYWyREqii6c0KKTDvgIl30ZwHkKN5imy3EdKVKiA1NtjOz8N/6L
lhR2zM30jhAw38ZZOuYCOZ+mXUoEuMbPXlHkrceExOw8ipdc2eGWUmeveIAwH87y
CkgBVuj4F0gIzt0f4A/8U1Qjfi9GjQOZiUrdeSd8tuQaFyEp+9vPBFXfmKkqZYQl
1XJ+5jIOvoniGcLGbDtZItQUiKYe9HO4kWURfhhlk1rOQu6DJoDJ/IsJ/msX5h5/
HIa7BYOr3d+//cpeyHV7L5tHyjMWamxmzXj9Is2Ba/HJ6gxoD0b2rIIElFChhU8S
xJRejP8+y8UPVDjvREgWnxb/nLPa84ht2yFhYSFzu6WHOm6+WYKHrx66+36LjOgO
+6ytSBpjEfrEv/movR6yU6x6TYZq07KQbM7v0/hzkcz6i579tnlrRmlzEPvZ+Y/s
Ku8liuxvlBrM9dcM3xxpaHjbn90RNeHHH2xJDvHtprEL9DFIxSoPXoGfM2oHgtC4
//E70PhSZBlwjY8yqddVa8JwB+F6Uy8K0R73R0B9QDInsFk4Dk+6r+J58EMXHnv/
0FJJQPzWGNaGzM8kt8ci8uAv0vt2CK218Qd9gkcCgzUIkbHDLxW1jm7vvyec8mkx
DMYn4HDg3xuUrgrk69z4KKYVZMjVTczYpXvVT8NXWCn42Wrgt88kEho+wQVySbCR
EbgoxROl9D8K9XJUZELPcTI9WqflURpNIHnzYHHTLGqaVxYZZxnGkcoF4IRZ9wqi
+/IRkTvAltk/NTPyjYbkKuxo8krqU3nJaOh7h4pJ83jXMBq8vdfPt6JFkCIrwYV+
KKZu7Pf01rnzmtPrX4Rvri5mPwE83Kk/UmUgWhXbvOCEncdRqrckG3/cW6Y6hNER
DyNwzVeWqZ0sof+Cr2RWfSIALgkjjukRqnAPRsSZRvYrO4wRCDXv7X6rbnyS6uBI
Ymf09PlDvt6Y+4xNuGo/4N7Ktim9X1nIsOFQPmTTWQjBLWnSRax+AF7pxAJhkT4u
o6gfLSBghvEol/HIAgINfZnyx5FwUhzLPW+zGYwW2L/IOOu8KClVnnvMzTS4v6s0
1/MZZMLBE5NZfB17IlMxiFncvu7lEWtvqC/4Y+CRuwI9akdYF2PZPyTyXmOD1oj1
KwnU/U7TQ/7Y9IMyQblP/0V8aD9RGLS8z81AgIfJoCF15g3mD67zeki8gMWqd6Ft
l0cSj69PBH36lku53lMCi6QSGVLKDPnUAxJZqpTbJQfPuW2RQoI9ki8MH2Po35R3
8FsZUS3A3dflXqYJn818D9ovC8FoqR1dgLg5XGF6r08GJKLw2pyg/sVRM/oDeQTA
S6Yo30XjOYAxoGE8BNn0ikwprXvfIBHu6jSHzhV0DI4ZOr+Tx7875rCqZrHhPohi
If8rCTtbNPMG/68ej2kCz2+GA0EfVXd4LWyFX8+3ua05F4MW1CkzCriGnG6A3MH1
T5IHSHyUOeuWC/YWIyoUhrJVqJC/N91al0yT3Gt0JOB8zzNFxFDJf5/It/GuVzgx
F0vXoxkx37TPOGTMqlKcBW2Fo2dZZHJIipp2U/rq4AYZ1GvABZrkRDmJdYL5geKM
nNf0aIQO7SYz9wmFxHEmyAs17seYkYeK/HC+5DTeLdzUv78nZNn3UTLCroM1Gxb+
JLFcC0aeA8yLCC5IUfkaNt1shaY/+gjCoXOeJ5aZM4imd6LjBUlSMnLpoISWT0MP
oeW8hAPnTJQKUdHuwLx6A67KEx9jR56I2bgl8IaBdOsKFjbDXZwes99slQSP7VWq
9ENBJF34rNuvnr/5hyUkgQJVdBT9Vv8gGd2vg5389oc81dF4Yww4aF25Z+m2xD8l
vI96FXDuZwqs/CkzRmmqQavhZWI5OwbAPUoyD5MERGOUsjbr066+efEZ/j64A14Y
Kq9gOy5xxnjyb0zTb1LVlUWRCRYJGqxLRaKsPnQagtOtVfQSWjGLjp2cuaWvCrOz
EEbtF8aYb6LcMTrf0Xog3ZfvfHurLhu13qd5BePRHlz3gASLNMj8I0K5yWj4DAIA
5zqEGDGNIZfqzwW0r3h90U2yUdO6FhB5pRlRcLeFmZxj57gdx6TopA4WPj7dTOsC
Xd2VAhKvB1YX0nMIL3N4+3Ox42zEzPurDWSQG2ofgvxiTmYIQ3v6PQoZrbZgNRrG
Ad9m64r595bDbI4VfGfcSN+KciQMdPrxEBAK4U86mo6731FH5eC5a809zr4UBTAC
WQEJ9jc5xL7tmdqC87FeEMLHUvx0m4xtC1qJX6r9FOB/eK75OtgDxnV8zo3IXyqS
bihTqV28qj36BoDuP0rKxUOqki4d26fRr0wpFzVSExAQKdHRBYFkmse7Wwq6i41N
1fdmg2vexxG87loAZpqgJS/jBbJtslpLnRhuwe6wnK340bQ1hRGTCHWi2wc3ejbQ
OQdEhj9QtDTYreXqIPY/oBKN3G597Ut5V7M5ltxs8iWUhFcyj6IkHdBM2KjvNtqc
fEZ82GTZ13TT2B4N5S/lrBUgOe6HP52jRLdvEEZZFsPCLorwpgi+j4AHVKiKjTHu
uAAGd2KvWaLEMod15UOBd3qP/GpSn5S/viiUmcdNGtcN6Z/7/1bScPrTrlXa7HGH
davEz3ihd1pFAYjkAkcJ9U1rc9PruBjjvlopHKX4Bq/vWZ6XO0EE3ESagaaU9MYw
HcQzi4gEtTWncQJLiiQAnS8ZJ1Cm10vaCrQi1Qo9nVvrt7iWHv7LvDDyEgrZ47DN
cQgoqmce/ui/Dvv08mcrM1TvfzIzIgiS39wBLgnPB1vrrc+shlTkKf5dfyg8UZJq
Oz3ivgxPklB7vOjUEOg6KSyXw1FwmjSWaIxGHr8U8qjrp2vu7occK2P0QgUbKJ5f
65qvWTpDs6d6PE7Znj54Mn9OMSgydCzZtLtRuaxnniqLBz89JnfRwAqWJwBRSThJ
dL5NRC+BHPlN/uN6IMwkzyBvbTI45xITpSh4Z3V0kwRC3x3fj8fgIJNmKsqXpylt
rwDGA6fQwQarRTrkj3rt7ODCk9bppl9+8yubHwH0EnjeUS1mXVuLZ1vB8s6P6+ix
9Oo/PmSuLiuVEpmn4XFB10/vIsKL4TPlbVx8me3VlbxTcjaQjdm6Wx5esGHLV/8U
FAZx0GBWWBWdRG9D73Cc1md/ZoAmpTr11+45ppsCkbukSfSnstZUMLaOccnXITEB
5lDf5LEoTzv20JzWKE7/X1+r9hZpIzgLClu6AvkFvDniQRV4qttcaOn3v2uMUX+z
JAB/PgGVD61P3V3DMlLTrSw6LzKkjGB4n9gGKUAnr74pix3tazn2Fxw82IWWmBsh
Gc1+lMg1gK2Ld1Ddyd6d5w55KViF5hNsHatGpbYYZEXbd/vV1pZlwnnmlu12VoZ2
PyIx0hbyuW+19W3amiCMQGA/GwMTkt3Tntvk0Y/GMRz5yHPod/ys9zAV7cH2XW8A
gMQBAGL6uA3bN8teDbbURTIT5zZebJ6S8TSu/gTV8pziHD2R6DDxCcVczAoeVn4o
1hIg0KRNosjRG9ajdYnoIdKzcO64LccDNeHAowHqT4AMTLN/YRa2kinyQ5OncIWh
2vppIu8XAaEPZq3pJviUrgDQDFSee0JvzPVj5erjpWNsnM/hQA10XNcENvYVavKf
PzYbE538hf8IVNZ3iFwm4ECLyU/beSdJ20flQOyZxSO6B1/605zZjMLWH2o8HR0W
jhgrIivjTSlOPtuMHxbIZJK+zV1RF+mDeAOF+TrcHBt6KcvUH6OF2z/1HXF1VUE/
otF8Py99YFrGEvFo0cotyCgYdkSLI/DgPEIfE6mwlAucgyFPcRs7Yreq1Hgq9PFx
cMyk7YvU6Y5oDoCqQnnPaVCZODPc7fxS7GzEDCeKNbhl828aAsLu+zBbEQHMbmU0
ohGzlIPgVoHxPXx1GF1WEI0VGgXE/x9R7h4vqrSqhpTs44YycBSKe0ld3bDPltfH
fTOX4r9VMqnD6d4H2gvlI5e3/qpUYkGEakisuVbs91HfdEozxGZwGBCyR0GKOtK3
FeqYAinivNksXhOcl+MfBvSxYx8O4p1tMnghqJCfL1yLMtG1ljq4EUEgR4ssJl2s
GCXwZ6PenxQbsZkvYbqPAKn6oxY4OcUd+h/UliJ2vI6Qc9irnREV5T/j/BNfkAwi
RlhprAPKbrs9Y8Egnvb7WjAac/uGagTqzD5nfaLpVebSowiEjZmNxCV8oTdsf8Y8
gFRcZ3ZyVXmAC8MyB7vk/71B/LlWW/QimoIFh6nMlcxGLXG62KXccayaUSjTEOZW
laExbYgC1tvxRqmD1TtsMIXb1kRWJofaZOedQpBD0OH7vs+lWpWcPK7l387/tXd7
xOYAqydYcIo8BiZGy3Abp6D726xyQ+xMBjxeqDWJ+etwguymsHOsTcYTaMcv4DsP
wivX5G3qGnI8Vabqj4qU4oiwDZg7EK7YQA+DUTlJ1A/PQQgU6INDKSmD1/G2UrUo
fklHXyc64sAbUJ+J6vL42nHI8maltsnkPI3k4kKAkKMZXEErYuUXL8dQphqtiFK+
HBGh/1ZChr+EyIbun7TLRxeY4V+Djamy5QyvjGmGKxLDs2scK4+NIt8yjkNARJjF
wYmHVszkOUghRIxFUMwKARxM6Qu3gaOcsGcr0RJDXEa29mgnTKzVdI8rrbaGqfxq
F+NL2SYdCCQn0GwB3yvHGGXVaHwaXHh9FkEEedyMcNV77ePMT4+ema5M4DAzh/Bj
h09Jm/ziDO5V3RUnYpuAnbZUjo4hLVXlhglrBJBNa0avGjbW+dfzYwMbrUlJ/1nu
nQfjOjncVwsBBrCkW93sRPSzgB7VyqaVdGTUe1jpgo1vLzkkjJKYHqElx6mrfv3l
JJ8faN4rqC2mSQgb5zSeLbWetK+blL9WxO9p82dLBXXqD2fp8wQK9cMxfid4Hze5
ctyRDf5lZYztkpaka2J3Z/nhMOdNOaU5QnOJVJUdzd0jq8wOfck9rPBqTm1wcf/w
LUwDMooskKYbsoazaJnJNaCTY7sf6GE9PmihUUUgVRbEdjxLn5PyO2Vb4S1X6HLs
q3u95Qjp9cA6xKWH3o6jtNGCpBxnLJnJV/QQaHNChRGG5v+tradjJRG76cvbfJEX
CuXl4Z3vFbFibDgpNvKBOwirrxGWR2CXGr53v0UqUQM9/5M/a+nStcJ3h213s4K/
QodzpHk0yChjIIP4QWNd3dIHCz012ADOv5s1wOA4h0KcoQAchA7QTA61NysJBVc/
9+Ph+0dmPF3Z9huhvz/58aBGhTEGIQOtFsEpJ6mTupgABjcku/cTP12fKPLdIq6/
`pragma protect end_protected
