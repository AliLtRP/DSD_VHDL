// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:44 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Kve7Lt9ft8aBK/dDcHiRhxl9Jkbr//Wq4VFDqGnS3lreg58Of64CauYQst+O8BZu
sLlnn7PrvqEO+ww2tiuKRiF8CCnQHFlcWjqrSyTL1WHNP/8UvJlJdhADV4NkOzkK
neeUCh6Ljd+r3zNYUiY4asFUA8LREiQpn5r3lmSsBjw=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 9056)
nJb8T3cDnKcIaQ5lJGkAHXMFF9l8DGyl+4Jb8SGZKZOIah4CNFvjMaTELO+NhXcf
FHCDBfXPbOWCGQLYeIFWytPZE3Lr60QOUPOgccou68cqNKFlUipjnb6KDEqizHS+
Ooi6SqaUOIIAIZcOMyl475q2tUTzz8VFXB549QfGkMmx6+SQIu+lLDr+RmAPHsDO
VRW2M2q2Dr2Ib2pwRJdYEs8aeaA27oQkzFMqd0kFXpm7NukvIwAdlFShNdtf1/cv
6jrOIAle6ZyP895+eoWNG73yNrQ1I2NcfgP8ppI8fkrZeh4rATOIYjdn/JhangVh
L3ECj0BPhQGhp1Btv0iVugG8RKGvVflSrvxk1kWvTQA/cj6m+sl0mLopoSs7KTLD
p1il2eBf4jtr3YUKCH4iTHQGO9YtYYpCXyXtSBsAM5CL2xS0qOW4Av3H884PZ8mJ
fZMuvilrYQYu4j6upXeYJz7XhprhwH5peHTtlFknjRquCFqQvRzH4/7hL5WdAj/b
mwDuZpmp/y6IKyq674/Jrmtz8VQA5igEr7Fwfe+b2XUWtioQ7+l0Foh6NWLGDGpv
OIj4WwbqBufLHZP0psSvt3hb46OjUBsxQors9vblXeQu70NV8pD4EDpix3tTZE67
McvQVi1MxWnr6iPjscv1Q9aA5wT36rrYfjyUmOtCop8ZCV3VYvoNJm9OPEHH0QVS
sBY31r6/rNBCTFXM1LdnXtS4N44spU32hnLBIdEzgqSOw5I6oH6iFpcaP9T7Q1ld
+YOwZUWaUpwDfygkzpLNshJyMEvz5AXRrLjGEqZE+gnks63Uym2lTEDmBR3J2NER
XXJ5jg2cSSKWFbqUcELU9UvD55iTe9Np7qbhOixIdk1zy8DMsZGV2se4us4ymNkU
cpkWmigVCUZ2hWLQI7lzfCQUwGHoPNoUyvc6YtPlzPtFQnV9a2JzNPfd2EujtSrC
ByhoSoDQqfWaveXGlqNchSi9zQ5OeHHEnDO+oFx9c6/0QsN6oUJnsL6m/5Ivb1W5
QxaXNMH0VAJpRC+oaXJ1qDzZ6FNhzf76+oqbN687immQgFp+cZqiBJIb6HZcMG+N
CvehfcdEwbQb4o4i3KMJHSnc3psOs0zUPpKnJWbL3plA/vAyljEhhsze+1hNSaBb
Zt6YCTPXgE541YfQushVImF/BcHRE1Hq8zSeSGWk/2S9sxeghj5vGDp2THOXdC5L
/LVdwPqF3Dv8rEsma4S0kfawB4Q++3y/PCltEQjmULpMSMigtKkkIBZKTN2uUSwW
fxP+LfCADfYqMaJ6BVW7dHqNk4F9JR6EyxN8wpCUq0svmSlSzjVsODaLBRLL7H5z
nTdD/iL/oVAsYIzWarat9wzuk3hNw0xGRTW4ZP1A5VT3I9lSgA4AvG+0J/14VZ58
IiaS6VGup0ayK820BOzBg9NsllsBKYRGAt2ry+uyuPUq4glgPX80OlIYwOrhIIJU
GaO9LBJJs+vVcP/DSdvvTlOv/yxYR0ra0aVyz5+zb6gEWb7eP8crJrn/dPqlu3vZ
5jSi4KqbTMTym5b9SAnW6x0sVfsidbEHNqb1l2gPPxZwhRbOtjqrxqXATzPh4o9A
+WeUxGm1JPAeDgyVOy3Cj0r+rLESH4zgyBEThrIgwM5xILLuiiubK4PKpa4BUkTT
zShLhSXdZak1KwWBbpTRb1+yuhIpsXZZFcfT+auRFMrTZ7L9E01PXsvUg2G9mRjz
LDZOAVl3m2FprmPEw85pjvEki96PcQ7yM8k84Rc6VtXq1y4WzLdWZSRw3cVEO087
aiOufSI4/XcI+551Fzm/93y8T1EaLkzRcRp+h9rtJtmHNk2mZO/DMHeAPhP2EK8b
bWQ+mCIUurHvgqC3/olfJd8OHOsx/yyB+XrsOpL99AFNMc/FteVcDb8J47rnjRt0
Abnt4C/WWin9+5dxwlnkkj9y80rxzBpFnwukkyohFL/a7z6ZnAhvPM9dn6s9sC8v
+7rzjFRovl7OHSTjzAdd9sEGR+WTlog5UV7qB5nuazc9Y9hhW4d2uwN30B8nZ2oH
JVqnMENUG70wwsn/h0mqqE6Ic5BnZV6bdaJFP4GtA2Y2CT3l8McdZsEkhCp+6OEP
BgkTYE2krdZ0GV4Gn04A4/9dErQLfQbrPht0KCRxfUVsAhH13IOLRLNiDJLLIy3a
ZRpv6WSo3hpv+CWHkd+c0aQgRng6MINQA0TcmGHMnnVuobAfzqpTAIr+RYVueeGP
NfmlCM+hgg7Dx5gGEW/9TsJxj6tJBQQ1YOOwoEYR3WHXM2QNm32iN0u2DFtUzmXA
W1rFqhq8y0w0iqGdRIZT44wf8uWW8BUa0GmIzs4c2h+0Ad2Q6E3I9w845a5vMM7g
1JQg1Nk6WkfeGUkh5pMRqNQO7riZN9pgJ633Za/7PDeO/onnVpVwRndmxVUqxITd
VX+mvQZHTehtTJKxo1hLvYBNN0xuqpmw68OHExipteuuq/5P/s6M1V/MzTzx8JtN
w7QbkgSoV4cBd0XezHTM3wDkdDHwIXTNvSTVxz5xHmXcgLq+yN5ZWunn0rts3HXI
oMDRXTCqDwpIeDHgKOSWP1GRxAYinpU+JmKBt3A7C4cedymwfLCWYPxNbDnE4yTq
Sn+zpl/IVJItbSjIX9Dp8mfORkt3bpLpNVf4BaS1zDmf1Oes5RzTUY/VrX9GrwOV
+/AW/YYi4M4pILZ1hdjiTn3dhZezBBitch7PEAnGLucBtlVyMQUFWY3mSqnpZs20
X0f6j5fEu4i+YjRtafKpoLCbQQKy44EvurNtsXJ7FtcbhCV4H2LHmDR7+1IM9N4Y
/46cq567CUWmGYjc3QCK2EYgnyIbcI0re/iPo/aBKoxsUh3jqhb4TJ0swsatTIp1
wuEpQQHNLjo1hjOlTd6rDnXLp3QzvmqfKmQWb8VWG3oZDQF+sZJL4FSGQkDW1vLo
lR9d2EMpMJuSUpCryruKxCZX4o7sAhqzxtA5IyVd19KajYdqMUfIuyF+YZMHWMUi
dZvWsLdd58QyTHoreUI7T7S7q4oUMfshGUDoAubyThIAJOsxfPyrVxp96r91QdjJ
XbbVSC4/c2y+t3TPIRUnKqBdPyVRCnuqnfO0Uh10ombnBna8CkzsIAX0gjkrkCTG
q2ZecMTPAszz+LOLSCTj/h7ZQMOuu9RYpgWoMIghNxaRszmlCK/y5gv70ZvNdRvr
YWB7IDRWWg41bXOow0vq+yWmmltLSvX2IE2pgW7jcBlR9LGCnTp73VLGAb0qGRvJ
tTquAbOm384td6IEQqlUBvDUK0m9EPBDGKJKd6NQ+M3Tpn4Y/zab9pqRrhja8dOF
rBYVwgrANTj+5/ARV9QrGirJjXV85lcUlL0Xd7tfSoThHHRsvIDkahncgVD2Zaou
i0wT6RpwFvb4D5hOLsKw8xDbWLCHDKapbJ5G24avko7tW84rWG6qkbUAf0XJ5Yav
Kl3hLpE9GRvJjupoPNojR08TfgAbWHi2xGF3vfx6XrbBxlysfsRAMn5lIKgtGcYn
VTpmSsZk166cvQBhqE+bqQOYJixoabYUMr86NSH6ma3DDgindbPjrzYKQ98+cWiY
tFSkfSJx1F6EUtxZiS7vv7xRyF0NgZnUkM/Y7xAXFcMUYNQMgjukCEotA2dcwcKI
rCNY1LhKcZNAyrXLk9Oi8c0z7hdDO9qemf+UwteVHpJxNiP18EJoj1Y+5dLItiIy
LvEGU8lnH4E3QEa3ZeP7HT84Y97n/BgIpI6gTOJagBYUStoN55NoALozQt6cWnHg
aZePjT3ZPNjO04PYSYnDmCbXdO7Fx3S8CjuMoUKygObvb49ZtGIvXvhu0d6x9J+w
Pr0PUXRmCU5gBq8wA9NqyfRLqHfON69JmXo8ZfkZyz4Mt4NBukS7xaQ7ugOiJgus
U8r8RH2Gs0kESAqsCdviKAFLBY/VExGIwRoBkDLmcp4bJMQCnDq3DT0cUsUS9ZpZ
68+c2yC2IWZ9mTwG8Vxmhz7ySTV1ZhNFHwXZzG/SHOLvDAozv24Y5xbPZQU2MxD0
xEOIDWWJ3NpbY5d/dQS1i0ZjG1fav/IAbSg1lPWuKDVdvdE+ZVy7uBXtgMNbKdf+
BVCbYmrTo8W7AuL70zhZFVhjISVFBPdO8jGJ086C87em0B42brZ0ykRacWiq6XFO
qsFp3lxXpvJxqxibeFe+z6jEI2BqQcyACEpgQDSKou63gODoPwFGb/JNfuZ2X3ZV
uE4Cje4Vz8Ub/b3s10u6pn5VBu4asa7E/ukMSgtQUiL57nspxGzI0UjO6t4Jqfr+
G4jgCfgmo65O9Xpq9mnLHS1ssDkqILQX+3Zz+4DrAbkctrOOoLR5IH30y/dDjgaw
HjaL1S26qxQyMnNoYuZMOERzi981u0fD8JpdYWVLMrgj/rjH5pw2Z6Aozk73mUU9
qdPwmzr0KFSX9ZQ3KMz+DbcsOxa8akRrmJsRF5xzXk6e5KM7cDVeMq9Dz7fGBDmD
CxPqRTup7lfTrE9SU3qRD3qP8PNKmUpW85Vuig/e5wY2Fq3KMIRDCQr1lbIhEP9t
fo/qF6wWH5i0kWM5jdtpaTaL3JEFFDEs7qUKlm56wZZ0rv+ENj4q+YmAdjWxvXxe
PuN5DqW4xgmNpEv/i/cWZ01L9eWrzYZ+v3i/sahuIAaTpzGApdZTKdq4JEA5K7kY
ZTlagCIMuV4vDzrwCbpuhlL/1kr3glfCskKGTIYXpXwIT6jVhcN7ZPqqdlT9g6d8
raiw9KAkYGVLW94xrMquSLCdmNN5pbKcW8e5+USePnc968a00yIyen0ONf7MN/Cx
8/sh1AKdQqgNV23794zqY4BuBMo8u9/JD6FxLPVxW7ZYUiNDv2D93U2+ySye4D02
5pTf7IgX526ymOch6P4QNdV2Wwrf9cqYnDaVqMa9V9UUXBxg3AUDkNilwAaWBhWa
EzXs6dRnwt7dap/uQKXa81q8aTyRm5a7LF1+gbMNy3IzaewbWwHuv107D9ckVTRf
O/ImssfBlI1WpsFE+X+wXPZQWRjmpIfDYy/n9GlCQna3z5sNmAvK7c9E9jOXIEyy
IvgkN2fBybNzcnQ0eVzSFYnxoiaDp8on5dAjF7t37sv+QJOBPrRpaJMimY9CNmeI
t47cHfk5KDgJlYKySW26PMAsUlE7BExkfoPr3B0XO1QDQfzJmXkCaOIpS+yKp1Oe
JT0GTO8OlOHRG8zO/d4krh9/hc3j5WKXH5tlcp7xT1lIl2XCdp0VyM9xyGUFiI6N
8hPAwMw6kREQ7zijteAk+6E4NrT4gjBR+RN9lf8UoODIqzRxDOfrphxnGcjcN60q
yKFyEu1tAlDOdCRkCJq09C/JyJiIMuDoGPQI92W0yOLvibHWkdI76AT6wMHoYG7Q
AMl0Tpg8bk0O9tcgRaT4iFnUVRi1G5asm2ueDVhOjynUBRdSlnAOuckRHG6ymjxK
hxaJbpesGzFgYA8dMmrSw3ZJn1ncOZpZ+pKD/bddTfh3XySDAQtEPwg5Y6hWkUdU
etbGHDw2qT/ZajXm/owdCSGN/s+AKTR93XUGVH8uY/OqzzcFO66c9PwGlTrVXP+j
7q1CnZQL2bsKcSw0rg3M+opgaldzmY0NX5RfHNBOZsgpS4icsqjcm7ks/mqg8g1l
xaDBBqvYaKl1KwT/wTlSgZYCOQxttRjYHUiV1gvDbvfSE1y/11lxdG38Z1Hlmw9V
wpDi67ke8fHEyABNpnUE2ipCpTH/J5UvQ6Goeh2/n0n5iwtJDf2LcmkyYkSPMzBK
VSQjaDEEK7lWJgUVbYfuDW9LMDOqS/b5KxtlAXFXc9bsS5aAAf3W8axzx6+2QA/Q
yMyHA8PlUkcRikh4EUjqHQ8pyXCK2lgvEBeWgfu8IKaRnueKan1XD3M8iP31HEdo
szwM+0lG+rPeJPVBsJSAvtCMlcnpLRlS4e1eajztHQKdl132nx8+We4qaoSLCsry
SwhWpfCmfGyhbyhOZWh95PMnRk49En4kXa6UEcM+2+axrtN/XwV4Ejaj8P+i580Q
QulKcox7b1ChatyqSyomIJ8dlNkVP44eRKKFKjEgtVUaTO1xXyDNULax0DoitotH
G2HxCwlLtzJ32c73z8I48VXeVunFRWGA05f1bO2SyONTy9o1A4T2YAYL6JyIkvfA
VX4KqoZd4451PDJ7DUIbutb2CPOAgSSiuoszhhXeocw7Vn71JZEzmFKvpJNgl+dM
pCfVOzPswotlI+5HFPebR+xCiIa/F/Zyi75k+1J3usyn+hluwPOGxM+mj8OA/P/j
89/Q9NTI1whi4HjCGlQUPv3k9wioVHQ36fgCg3G2ELUFtRrLheyjPKXI4ycN2/7m
WZRjVv/GvuGZrjjxzNTjtU1/XdeFUnGzOPg2rvbbZFlWugkKs6W5k2enHRQ5J84d
p59WjePLWWjTXseAOpeEwe4xyXjRRzivd0bqAAYPwPdUO5Soi+6Gjm1rLDJ6AMoi
lcotXgcUJgLKRkDG3lKx7EXEkRLaGi6dDhCgrg85Xrf6G5CefG0SDI9F5c8qFLLn
q0NRpFAlZg358s17tzmFbbwBKk18OanMKEyMSbyWmdW96DHfBBeHiNDy7QVIPOkP
9UlFURJipsQetPGIpDRPiyiTpDwR6DyCxdzDyncm52QiiUhtNAwmlfiT1a8Xfe22
ray29xzyov6cxQNW4VhiHCmXpfEeSju8ttnxCW/iZiL5Q9bgTF/9MMgxKEQDPTqR
f/zPsWlhm364epW3nlUjk3DOOJSx3yFHyytR7KaoQ6OF5NIs5GN8Q6j/Xh+Lq3IH
2/1Pf93qQKLQWRdVSkdi/g8Mow1dznTdg9gM/XtjZx2Qt8B7UabH3ww5Q4BNZ90c
6092PNiORQB5aZ10Z8/YkO2ANPPYCPpXfw5fywMSSJSKc6oU4ZfqHVG3/DKLpOsi
RxT0m5j61iFunkrflaBwBE/jvNN780O6RCdt+/Kkesz2pmrSX9XgjNsN2B2NMxBt
SXHGj0Td0gv22POJ6vmMhVFZbaNdNrs+zVKH9rnSH5STFRKKGg1XH5qy14H/ZkPQ
GFsiL6bVUlPELVTPssI7K7ha0cI5n7rmoUkfg+QBJejSPVq03FleU7xeTPir0x14
b3/Cd/pggyArxfkqsZHnLIuXjTe1ztjnYAjHYBbliMjtqh+Uf33rNFy5JR6+hJps
29kq2mfVZv+wZqstjUOFdL2j6/OI4H1cJG7jbjC2EYa66v0DLI8T4XQseHh/R4aG
Gsj58ZhxXfoiqIT/nUYF8z+GT4a6zbL9P7eZTNJMiAWC63KoM/4xLy2CgIBDuijw
Dm3n7JfyeiOFUepEZk7kYBwrNQNNWsDhcOLA8it+Tiqtl6IMI3xv1/a5fRMWo7Fz
QYH9z9uVXz3Wzw3RFhyTFLOLDdQO98A0W9SEu2OMwQUP0BvWolFK3WwVpemGdvQG
g2iSdIkqVF2KIkElF6T5/L6j1y/a/0T0OzEn93RLS0rocGPMUoq8TceJMd2NgkLt
rjhBRGwY9GJe+6R7lDH+gVqJvUzKgrOKJIc/6Gluqznc5rByAOEts9kUdPc0lZtH
XlKkyRJQ+h8NSQ0BjTONxMHICIlBM1OFT6jQ5m7jkziDiENkrFcGBhE4bOe7PSBy
2Eflkjw/lkm79fuPFkGujX/5QMj2tflhL4JY2suKuA4AZ/kX4NhITyh5uYTU66Gm
lK0TqVz0q0Wst/+xavjeNpFc1eXaD0MC0r+Ip2AKjzfc849BJKzKj3EE1ObdMw6g
TxJ0HfEDBu7rlW2Tlpif3+J2Y5JgJPVR71GteaMhqP2eSe9bwKIof5wA7LZv1q1L
+m308UaIP12LyPGnSh3Vx2pzVavCmcKdxk0iihCjEVOzm1z29v+seqsFAhhTT3ZE
Rc3eDgv6N7ePn/WUCjj0cF7+QEfQHu3SGAI3ueBWqdmwinshlB371dM/zSTNQja3
Obqm0yjoJ8uM34wnCavwgcxIDd+Zi6HgRlclHLxQoQVzdidlbtS1ElLwf8/Rgw1v
XOg0YYvJliwl+m11uBq33dy57v/E9KBrpjjaOhq+b/bU0Qmzg24tZK3t2hj/9C7i
LXbHAXFhLOODMrs1zIKJN15HmMgzLM/2WhzA0uvG7KikVHUYUwli0xG1BNpR6EzT
GODLVV/6O2/maTBi4OTNcPjK6cGuhJiiasPjL5ndWje1tE4gdvnUUT2OzTQfzwEu
amj3ToQ17ExiIhj1Ys9bA64DFtUR2C+RjtgE2jV/uZSXKPg1Ahr09FBIdezB8zpi
NIxQUK4rnjTJuaeWknxOpxQHDC0XqWp4siPpnMLGJ0PK/gtV96ul1Sl47J7Je0DM
wBuidycdNZP8BHJeMx0NIldRZroiqh8psn9PSYRlig5IF9ZIbhwRuZS8BRyjj8J0
Tu5A9NSVVN51kfhJZyQMOelUvgdUFAVKiFVte+asG27mHcK3+LB9yoKfXEqdwMTl
qYIWrQB38LtOBAx6Z0upqI8xgHuWpW20iS3GYEC/yCPYuB+XcziJzipHVf1cQ1J2
Y1LoxtJ0bb/Y6BIv5f3S+1Xcv580yIJeBNdZwA+aIRr7rF+nmObqekvTiYqkkZv1
gUnOGAbD27qSbIvN/1C8mlrAlAi59dF++kpCZAapQDxwo8o43qk7Z/GzRn6OwFTM
pslDFY5lbU5r+lReRbHtW/Fc/Nvms+inQV7zVP1pGqpt5pLo3tYTA7yV1KY6/X7B
oZiFJMCo/JmBm98N2d45k/zoTCkyVWucOCO5PSp0KG9gs6MQVBE7prZI6sXfPiYf
74aoC06l5xDk/UrKM6czDaTvaaC8P5d0Itv0AOTo5yXmGLoDFZfbeBayxGiZlkMe
n3bU9bgErn0xGG07KWm8JKTQIahhOx9jojoUrDzVWe7FU/xTbg3rzTXnr42MbWws
NdComTLdM25CrcmuUIIXptwYcPtzFaSEBgjkt3hdKET9aUbSaA9GTWbVhJfkMgLK
CfwmnIXOknfF78lpHYRrPBF1ZqvurKxxVZK+q/nXcSswFf+i4J+/jyhz6daXwfGE
N/YRBiim1vO21ZnIKC3CzTLs8hdhXAGxkqDv1XxQl1keoIcohWmRu/r50WluGioW
zorlgsaAziYfKjREIofUgSorlnIlr+P7RpYVrQZXMpztUv2CCD71yZRQ9ZWCW+nm
EZ8l4bZqIhxmzKhVv/B+haFwRpCSCwXyd6eyDOFHkoCFuW9UIBN/PnajrPHxLGeX
aaut/+PvpUQ7AiRSMs2p7p7YTuo1fT+h73u9AQg1M0NpBCA5viXRE6xKNwUBMIwE
DwCEDys5XHYxaBE0rZTqFMcH3clVDJpdYcDgY4bOQ0IozPeEhRcbs9NRWhIyL+xF
qgjLIePapsuRIW38BjDq56pKpYlDwjnwTcwSEzs7yKCq6HqJXG5nAhAtPOumTz0a
2MJS7btwK6yH7Dlyg3Lu2cXKn6aXo2a2cDJOw1sG6Pv1Am1jxm9jyTpuD9lUG7oY
ijpJZz1CZguW965V20U+pgF3p0Ty/GJbcHLdxPRc47Wh82asdNvRpmW8pj2rXasT
pezmgJ0I2BerhPloWrdFLnP2vpx7bj1zhTVBoyYrCfIK1qErJSjgcIpdjH3XkmGW
DcnOyeIBsZ/IldVLvBDAj1xnvPbHWDoGN4Dw9HuMVzMac5dVb3HsK1fZOhzSbcRW
H0ensjvO+v4p+5kDgZx0Auu9fDYIbXuOiEmZ+wJmK4AKFU1Ib+Gk4/iQTedrIVAi
HNkzj2J0izE31n4qaqmMyn434JfLCVh3uOPB7VaCr1z6utraSsIMLpdWa+IkOjOu
gwEKOWrAytDDG1hlk74jYYzK6Gq+hnatUZ8MCFeattFvZRD4mFVebHqbjID6mzdL
tOtW8pr8Uy5rADk3dwgkcMr2drBzWsFFYN1OdpEa5PoQZe4IEKUKbhj1E1YK/TXY
lh13VGt4aPD2vSd7IuO80BdjsxMzpuuZSgZdWH7MAg+Utob6yXNHyG6Pl6WnLqWC
6bdRuKTOgPiDxy97+5jaXG6t28kUqRgip4pQG1k9FtY3aOwHiyqTxjfFYv1jabJB
ZGpYkLpCsr6kr7HuG910MpRHJLDDyRYjxYeFlmU1NQJfhyfUphgPtD+8woeT5+j+
vB451vN089M9J5OOIXuuUWEwJcxP/VnTjA3Owlvazu2sUq6nL5bsa4egpSLGqzn1
HJxy96ulLuBrqaHAmjYM6RohTI0XoVv7PU7k3P9hDxH74s4mOkdUlrM4XO6IQYHe
fg2QMs5X3ZQTuyCEstJogK3bu7ibF1VOf4eGC4VzR9h0YxXKh95QrbcoTCyUyFGz
+5N+tfq/FvPxFAZRnXxYOvPb3HaQtdJS1AiIrbuIDsWInAtRmIbXCvVpbCSOZ+ru
iuzNReniSJnFUC7aem31T2+rcw0ylCKr1eKU/RAhg1CHB4lA3xKLXxZM2w44dvfS
hKJsN70p1Hm4QSF9oF/ue7jLAh5JRA3YersAy8HEAPn5Ozf3T+GULC15ezFz28WN
0vDKX8975vBqcbS6uQZBic+H7cSgJ7qJsn9Sm2rHRGnODH1WlWobVZcpdVu6mJZF
RnGoGqvDB8N4lj743oZQyP8L2s5AQhPoJooRbg9nRLuSf2hJj7AWjGARltUTpQM7
aLkW8DwR1iem4BQHWYsWQf6ma5qeoy97aheZLdrT0/tjOmzS/vT3ng9MbnZ3ykhF
ld7tqZxTErtiUQkdbjXtEmYuE6zS8EzFNfK5PX33OqTfcwdCNJsP9I0RNtgWtJgZ
UGQR31EQjM0aLGTro7h+MVd8/PAdRmuy+WBwiL00duMR1nGpC2BhoYwb0wBVV644
qXhyQfaNPdmiGd9DMh/yaKSgFegI/GmnSLU9hgDLnub+Wg2Lx0UwAHwaQITQQeES
P2154uP8QKkaaqBLwXkEbKT3glGYYhs55kWJn+uWdZ4FkVsjSOqDcDFk0EPWyWWv
/AG3koyLeIBHOd1QyOuzABN663GvCKIayX2GeaKNz1T76Vb2ww854ll2TA0k82gx
YnSMcYA2+/i8TPBJFyh+9ZZaB4ihhioLNK3GyieaAhOSOYlFNYTnGjUNya0uSmn9
9bIvWE9hoiP4RrR/9rQeGTjm4QpPQyRCdxlFKABtuHIDNgy9jPNOzmuhqynYrXlj
Ktpgg/nUj01aYRHjThH/sORzAnALc3i9VPW1PKek7e9T3bd4MDeZxz6Rc4Vd9C0A
S4PTzMZSaKv/hGneV0n2ACnu03kI1jtZPPsdYZZsZeOsbl/QiEqHeqPn81xMeZE7
u79CklRHE7ZLDahaxm/Yhx1yuRFp1fMY+L1gKH56ymuOSUVO+tdTEKw1vcJe+Tc3
UEDUHaSJ3xi46uHMbZALO6oVUFqZErhY7R/Gf40YjiOg/RPsPLh9eFyvvPlbR34Q
HNfjv1z3sCPC0fS5zFXjuo1ivKK8+HMc9dkblkjVqBmgmI4Zb5HqxAgBvFyZwjqf
hLXs4x3nCricj0SkS48cUP0xPOb+iHEEvXGOQqc/wVaaxPTIFxGAc5hEkN2tOTGZ
lEN6MxXCiMp7SKUnE0o9VFBYB3c6fRvEFFGwvSpISjnvOW19/ZnK6TRBRDwwJJkO
fSq1JL997gbf07dtepiXknmxAUjuRDcd94x0MvMBTXe0gCipE5UJcfjHAKme5gCa
OYttD/QD11ZwcN2MCXVR4L+07lRiLdwbpJE8m7RK5BbecvfaiZBisnQvR5cYWndr
FmZBjJx754Wj9q0HU/smZt4lZjTeZ21Zp/oRxGRhQOYtV+ACmczQCWcXFt/Z4bza
l+McqATdh29Hwq6i5SJYp01yASb46UPH6DkXi99csvf/qqY4k2d4ZdZWwxlEDIh3
Ed50ve0yKl5/626QRQ+muas5Sp7i/8S9IO38YR5cq1/gwRNiYxczhWQDgybcow0Y
siHvpsJwPzKN7WTlEmdF5TSLpnSb+xF6ih3AWm5CF8z7Cz4zIa0yxPEgjSPMJpIv
A5ydvsHWL8DVXSwm9JxEOp1JT7C0q2thgScyUyVHmZqkTDFkSCaz4+q4rF/ibML7
sgTPaDwi/uFvm9BLLr7jTce0xVKpXnAlxbt6F+U/nt0=
`pragma protect end_protected
