// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
s695BwWBLTGttXy+DYSKOh7OdQ2FnSCEVtE+nK0WM6nGiyjf0/3EQWSso4/sjUwMAGmPuvs19iRE
8Wgvr7y8FsYhNDonjAYisW+ljpaN4cyJlOmyTMKNhxGaj1EZV6zZ47tFLMhllCdBRc5m+gxJ3W28
GQq+U43JdQStiD3qAeYvYoFFZhgMYrk7H+iHX3qJ7ej49hysd+r1EV84G66TVUjSX2NRWqWRaq3E
uwLcBDJDeyoJJnvzXwDxZXYxGlGfb9Fnd8w3M3NIef212eB49Cdv9qDlWqc1INWpn+H9BmcfeJtb
uf0s0eMWZOH7pWr2tLCltCzbggcEUXchbQjVyg==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
EAeJiFVgT5MWVpHdjfdbF+sB9ipMSsPZwS8OOzZl42rqHO3cKvzoRnJgYi1iD/nma3mwDjUr0mpP
vNetLb9eMgRc0L/KWHgPTPYQikearzomkUgaZV7zBM7zCDLjqFJa2Q6kbIyLIXaxrTEyn7Z+1UUY
8jIMSoDQ73SjoYLVfzl+Zn5YXh8gLFgtxK093U1mczC16M4eaURfntNrilx+EI0Ou8sloRlpt8PR
yVXHYTpQU07CURys59JJQaZTZddBqeKrfssXBJTmmKXwth9cy4eZDnAjH3oAjgDJMt9hNW7Qp1xp
51m5JtjWObLcpJSl3k2U9R3hxwydfYiIoJOq29/SU0K2Twnfk8sGJ5IR8a8SRm/rKHZr6St8fTRw
ABLzag5+4NPJTYODTYfj25cEymyjYmUAsffTCmNyCOxOs3DRBvdxleYEsWgTgkB57l034pE22R2Z
pp/BNx6i46mwbqQHoL1vH4K6+pnHkYHmjTgKvtapD8P1f4XxdaY9xraGPvwezSfpfgeyV3xmlWqe
y7b+bYZWhkarJJhq4HcajSeTehu0sEtTEOdfkm6cuUtYxAFZFgbboE0IIDyOfsjzFIWLzItqDp2Q
0RLrBF3RvksRTC2WRYm044tagpWtHKRaxcNQ51Rq3+ZIxmezYOURdOvm1qZ2o2XXnAPcEyqcmgl6
UY8l3RVQbYFM0tAhk0QitfvM5feHsXiU23NQJBuf1Yk5PvXgxDji5Kf9pi6mae2PLLeEdYi48dow
Jo33q907KXUzaAIZkykoLl+7Jk5d0VBTsoDwJXJLN6M6kvq87T26jzdLi3HkXSXEF11l6cGYMlKB
yAmHm4bEIUmp6VSLWjpgxbQpscRLaQR4+opkFuBvC5e8DHANpByR50YzjzkiuIdgbr+luhvd+LkL
s4MhH6MBioEmdyf5TP9hXQIoGNsj9u+4ZKlMLr1cWuhx446V86SxUyIZI7UdDWr4gY3ILUdjyyyd
Um3fCJiaMLX70AXYZ5vjF05uYqI6FDPE8u7WpyF9NZ5KLFU6dKzO4RX6XVYjsAW7qEzebEWJeKmF
nSU0RCUER3ZxwjpAzDiDFMTbQMW2zyAAnvBYeS6b2c8BIz75AZbec7WApiiONLcTjAWnzUOxKMi7
bwCLB8mHVHRfauF0t/UpEyXireB0nWoN+OlSOsQj5NMbBJfJxt8FKkYjHDWGxlmPu8TYpk08fyiw
/EhGPArjp+mBTGhtgOogzE/z/cMv2k/+oxcX6I955vpa43n2JqZ8hNIFSrfprS3TRFbRVycMYQ4O
prhct/1CJnC3nJ23TS9zfn5GWmqDR1XeVXu/S01+oo2rD5QELo0UbvKd9RF6/nHB8Xp4WtVHwyJB
XlLHE0u+KABk4m9xvpnIJwNqMj5mjT/fWfx75Q2vNzxGDTMefRTwS91C/Cbin4uemFPeq8Tkg3W0
T2HiNpLDBjIjOKClLIvcET3zIN+jD5B+VU/04zxjnOWjo1UHsHl/WfEkijFlkR7sU1B5FxpnVVO0
iV/0gwqeRGMBIvWss26NfSdCsoOmaWojnptW8ARlJQlly0/aM9eWFYY7PwjrS9W0VH81vHu5ChKo
q70WB6UMlNwEXxCaD+nueLLCFg950mv0jDQXuA8upvcYN+dQTKQi2U1UTv3Q2Quvtd3j9QIyCKD2
74yTBeMnIFhpEe1pRAWKO5jm8+vwnRi3ZyyAeqv0LqI7z3Xm1cAee9r7T2LfFUAcWF13vvWaG/hv
lfdSUVy4efpeiF/OWMJUfp/DTsjan6ne2QQH3EixE8ZAo1k9H/s5RUUVsaLZmDxzr78zJacu6GYx
IUAnfQX9yCgI8HUQOTpoB5qozkv338P5nNVIchJ6l8luCl1nOKr9IVJYh13KyM76KL18NSNaCtj+
nrFHETbsEYoqDbwCe8m9KH+PpqqMRyhJXte4+lIdaceBt6lFVBhavrge26SfMreAP5WtQAU8LRwD
qIttukImama4W3FKk8eUc+k+f9OzcD1a4idhegB2YVTftdMIzZjCffJyzkRZEbfb2k0/rZGzIrRg
YRhiT0XyNcYEiZ+NRP28Kz3dlTqU/5eAqnVrsjSXU2UR/LjlghLYItKo5Vr7athl0eFHiEafyka/
FRY+kY4zDPjyHVAaG9zBRYDmXUAEMhrwprEcbWEmE7HtRnGudg4oPk0QVbzipKnZaHSVe3sYUYo3
OY/ylkLMBOU3phWp38NCjM7zM1rXuWIJZCfjHTlBLxw59BOM5OYLg65oeNVKwcNGw2cl1DxR2Mad
doOff3u13FO3pAX+/QHp2dGytWgiA97C1LtrS46/OgkevO+a/PM5PgCS0tb+k+u2ZD8J8ACmOGcV
geTcqTIqcoqfajmA4IllaQ75GvH/EkK/MQQmzxAJxwycGPASfFCUSEOsxXzk5b5l9lgobOK8xzY4
F0NoR/IBJ9fx80Iyx4P2xMlIT/IcUtrM+e/9k3v2hwkOMVsqD2lszhoKPzLkMQ1BPzAGqDL/oaS3
pWl87WaTMAf0PPkAfzZaycmLcuRSXx4w2Gp9+PS3Za5au6oIk3FhW63tjP6g7nZBKOispa5BAqIn
tukrANt7iFvyLzN8rCBh0D+J13Xt61bcl6GMcawzCzeDspsFmbPJ9z0pUqpjhj801fRdmDrBEwcj
i/lAVVRv58dOKRwJBDwg3F05FRkxDP9yhuNIcA/xxZ0nn91zcpuWNi28CP0+qccOOYIalhITdGN/
c5qfvzvyZPnUz12ZZcti1euFXxUnX/FrhENAt1Wf57/xL7EOTJI0ICaoKcjh8y0AJlBwtRe4Hh26
wps1hCC/HiAkfAukPg3+uQydY0hoqaPIn1gvsa3pkOGe7gFnFhAyWWCzxI/nkOgLLeC5DiCQxDNA
GnGtFG+zouqAjQNL1B37QzsRWJtg9YjIN7JIQ28oVMi99guuQqw6htU9P+h4z/r5h4rEUTtiwYnr
grNT+nGNUOF4kDgs7HujTDFhyE2kNSERgWA4B4BrjhCFebs1cxwL2vOP7r5MvcDiA296BPtwvyoh
emgcx9BTzLiF62xjeAtFmmQSnivPCaq1CgxLZRUSZHpFWiYj/vg73NMyA4n2tv/9kwtsO/oYSaus
GLpCMG29E+0Wpkb3qDiP/OZF1M06cInq3mK7C/P88fS/LQ3Uxp7XfKDxO9dGtzi53O9gJoZaPiek
GvFPnOsxj0IS0PzB0f4saqZz56sx0C+RXvFs4IoRWo4bPoJ0K5HHUw3ddVGw7yJ7s9n5c5yVF4y0
nEIJJjto9nxC05iDdKmdqnJn4Yhq2Y9ITAI2s0WCSYK+Ail3g1Jh/byQyOpc0I/Sfq5ngWBgvrEg
1yJRERCDJiwrTa4WkJ6sZ1Of1blJjanzc4+4m6q93CBNIre018a72hfuU78eWLKhXLsKrfqaUP3P
LmMuhnbzFx1y8x8unK30dR8U1ANiOjaIZ6lLZSguGESjAVCQ6GFNQZvCepLxwx3uuDzlirOj2I/W
j60nIMRZ4WfFOZTQfzoA8ULYAdhIwxZjCAIUKPtTpkCdJftrL8UhbDKyi3V7RMcJNb6+BapVdqeN
cIvUZcZc3wS2XddKQFK4ktEeSxYVCBTRPCnK9MyU+QyZf4noiYGPDt7Emn5z+iIarRB7H8r4yUTB
EOrPs9GbZA3VysPECHW+HUYTMhfkNZ00wtBWKynaiow0l8wv6eLJjrUhtWYgHWa7wmvM68Xv1MNN
BHLU+kOw4jsYwDBJUhs8RRqrHRWr9Vl1S4sQBOcN8zof5FBBYN9G7YT+tEmzKiPb4SpP09HfJNTi
EXQUnaEDMULo2M/hynbGeuEJLyittM2AYoQ5LSzhiMSo3Y8hLXHYsQaX4g+givhDhOwYGsBTMuTv
WDZhRzlwIXDuZk4O7s7wHnHtGjZYgEfVSqC/LLFUJmmby3JIciZd0koM+G4LiIx+02dAqjJnTGIn
Uo2bpb7QXV/0OrlWx368/iyHJmPw6wBjVdCUd7POIy97unYQIwKgsPpRQBjQjBk4D06bqtt9FaqP
MjTpLnetiyswe5W6Xdl0aePvwxGSweBZ61G/bxrRWjy5REcxi8Ayh5lsijxryP5hZaiGVtA173qu
nxQ/hn6pGS+k4BRfjVfgRkhZTqFZ29toxUFWt3lJBvLHWJa1RpKOFF+PZwys9w0jEGP0La1AXdH7
WDhNDYUcg1YQXJE6JovINWRgAGTZlGqLpl7OIGvyD3VnGjOOrDdDJPGXf1toTqxz2LsxfikKX/sv
01EpuFYIfAaQyZRb2jWsgKVLdMNH//5eRzhw3YJx7SMWKkiq1A2sulE5T6fsokiQPtRbwX7Od6AY
wVZA3V0PorcZw6L9yULRarcpBGWOW2MaPixMpTDMrsSyUpCT4hhl0lQkkZLHxh2unDuNGu+2e/F4
PjgYFDjhdjok5Ncq4BtheKfodrNEOAIcsaodpxccEegqbYZVVhEnXMy5v6V6qt3EW44ULnf1d1Av
rKmPhxCqyebQ3zObZQrpr6gbzk7b/DGoDx/PRWQiuuq8wxRkDT7oT5ulvoDeh7vRsC17VLrrdGAD
sdRUekyZjC0HF415AHAWRoCjLzs+FhU0G7JcOUOjE+mE9bmjeNHpHn2bJFk/peO4RejC5FFRzq5P
YLjRAGm4+CZS1p5mF6a+fsLEc+0IbhBK3ReMFdEIKNDVdxxLQ0e7lpfLB1P7loXjlSC3wQi48/5p
9utnrOlX+UWZI/Zr+X+2Mg78C/yRFRmqvSEyT/EYREA0/8c5rmz44/l0hGUWgiBMK56+5QbqoMW4
Yjt1aVu4CkBs+CUzweyPw1QvF2IQhSoO7SYTYq3mcdyWj07x8rDcqDRpOFBvSWVJnkH9bWnNaPWT
T9SE1SQcQZQlXd2TRlyDXYUrFy3CPvB5Jltz9YL5kW05p9X8SSYFE8aEnpp7esGvbXCQgv38o9G3
usbebP9R4DzNJbCzTaQdTgv5vwYzveytba+byt0ewvc+ynvd+sP94FF18j5hm9q5hfoAcbmUGTCs
BtXfr/ZZDu1mD72F5+BnE/dqNB0mBgJN5i/LahNdYxQCr5FGtiBbBwjoXy8EC1Ji2dobVEAOHHmg
vVr8JnlQNUMnNI0K06olhspqNCUO31bvNYr3GmDqc5gisX+DB7taGonFX8I9InmkwC7GIZOCiP+w
C6ACZ2YcaKT7gVKBGCAS5B9zcbuYpaQXyitv2QOe8HKDxXw5fnd/i5Ob0ZHXGT/VchHsZrGHTjbd
yMCPDGbucd1RDvq5G19lazfxkITLF27b+UQ+63heRHyY3TDn43jDwYspSTswS8OCCis/8O6t9jJ/
2P3bEGJRVBUGmgqHImMNph8epSS/W04yI/X8ZkquuRIAELt7kLC8/dniGTIDSHB2ES7Gf5zjSyqv
jr+GF5rJfXB13FRlseYs+54p4m6GOyBN8rRx3LChizRa4rNESCQsQcBmZLGVv/hloiw/RkFF88xj
tmEOd70AJdxB7htlRJzEW0Ewp5pOn7tLOQbjcCWRvOv941+xHl+v4C/stzMeJEe8tRyUJi9Vjiij
38rEGgvsJFH5xpxmuc7+eiBsGERA0C2S3a/wnR5DMMAKCzuwtUFfHGaUb6nhxwunaSvvF0lCH61Y
/HU9JH7JSLyTvyhSE2KNEufELR/CS67CSmtBIQyHAmIOvaJicRGg26yOQVMZPr8m/iszNWd6FMjN
VTYi79AM24XBqU/QCbCVWDBu0jZrCacvkaRMCgoEZJ7DEPnrB1i9u1ifrQxvhu2rZ5wCvqc+iCg2
VPGG9odKQ+CMREz2kKVMckHYRWehZ4wWSLvrN0Yg4LCASWK2mpu10/sNh2o7aeq+tGDtW8c3NMrj
xauu+LsC/uT/wFK5cjMhHHV2dciu4m8MxG+eZj8CwTzCerhM6U5rY7fmKAGklojQW225ddXeFDP+
KZwubFIXtrWDmHae4fmH2SHU7LmzvE+bBsdxvrWONVmCyWspnbX0ez680U2X0o6IMf3Dz6FuYLaO
UcRwgNgv56su6+x1bboYm8kxXFUYSMHololxHb6ORmnszTPKQ6sKvIy6TqkVs9Yd5yAYBMIaLgho
gqC6QE0pZG2lqEsxiDfGdd/xexEFIpcpC/aRbDkpTsrHOKadcGE1LS+JppbdEVHzOaRivkrvJa09
xZN4nzeHdYlcX3IvevEi7KsHt8qVHlS50UFxCvfc9yAJqm5yj6LM9sTm6M7a59ORjkWFJLJG2aQ0
gzzgh5rpYtlluVBD9p/rtRMaOrcsSPxsWrMlVOJABAqZW9lGShR7AtQNkra+hmwf7wKuNpa0YUXr
2Y5h2136G5Gc5DyNdMXsu6VkLQHdy9A/pHnze72J3A12NZ4S+ZNAwWRPEUvbXmlNrKaM9o/VuZu3
oTbBUe4zGF7EJfEeHp8jlQNSS9be3D+aaBqEdJXH+wRzx8V/knJM5PLMkzjYOLrDIDTz2N3MzhfY
SAAXHC7xF4xk7NmBNHdi9trPHNuoTGz2hq0Psgp5LHE2HwVgpquOenQNYg5pTm2Y4u07KsOubIlp
cBknPzEoZQSy3Q5/Y7COgxHAn+V9MIaXxfdFysB1H2pF4fGQRP8Aads6be4QkEyudpiXeqMxk6t0
Ag==
`pragma protect end_protected
