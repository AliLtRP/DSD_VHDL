// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:34:00 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
ogL7P/NeDfl2qmApzYtoEPgY8+xuqi1Oz8w+Yjhedta5q45U9k8v+T0ENlGifwEn
jYtKWRcdNXQsCv8VnvETqEPW1t9ED5HqZY1KPceSWti/hCIxDt139epLAwdJ2HP+
S9zyY7VafGGiD303NAN9yVn/Mr36IpTrKfMcORaIQN8=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 27536)
zb8RHk1BlO9BSGj42zQpkKQWeTyXaXvqvCNa69O8UFzdI3rk7eJrOiEicjVJ1c8i
tEKXIjEdNXg6bGUXkx0IUrhXI/SMNlNiW6EY/qyr6VSxlHq4RrNTorBZWMgaxTqk
Dc8Zj0oD9gVz7G1OaAmsKvy2n3zadI3+u3HyQflx2SYdW8kwoB0poMK89x5rw3N7
oI0RtrcnUwG7Yj9rxzWmA5WWjD9EqZU3kUhLCVgvM9XgJ1e4osTP25u+dMLiKUAN
9kaH2gBT3TpcA/U2LhNvFFIdrHt3AYGs/MhXDmDn5ICfVq1OmHd0PcoKY2zR1U11
5I10YuHhEgxKHMoJrZ3pk1Svx64atvoNxFgDtNukRhjOosOTtkUdU7URHzLBbQ5m
RhBaMPX+cNhvk2q24g0jbT5DqCbwWn+dGKTgCwHTr3UuzBAjh4UtC0vWUNjWJAqT
x0fRO/79OCUPrIhIvZZTYuD2U95VfD0EyCagD44LCpK7kxedUMSbbN5mcnfIh6Cn
Z3sNRP+Z4qG6LxsNkK+Lxrxxk41ykQVcFCbZXSPypR3RdGU7XzFgkuFAkrMNii0a
elVjVheiGDxA249zzjUgunJaZuYuUzxAXCu0rsmfurNOiCg2MFK7e1TSZh5h86Cc
ngGHxVED2rcENNfNNPge7vMxzi9hORNMfRCkm0dUUawCqeJ9eQqhx/MDtYqjIvoy
pGTWiTYGJW5bpDSS+JuP2NvpFyz2Btq3aQ71zkDcIVEh+lyIf+hkv+DeD0OTq0hq
9vLQ7P+gezDeDZs2O3e/NvH4RzXj79f1U9Dd4fivl0gRCx2Xc1yHWhb+vfHNfJOu
Dc3WqvimHGI/OQg/1U/1jk94Cmq5XIyE6/cvt5tdBBIEBNRUZJRN+sW4SXji2R6j
HI4sTqoKE4qpD9uoPmBPqEAU6zrCXEZI474DFgWxo+fRDRW9HLL2/9mDHUuSq/vC
dGToWwVbX94hhIiAu6bkJopajXexA3nauzxA8mhpwhJbCESlXq3sPyUG9390CPFp
5sfd7PMRh27Pbrhj9aM22EWs3DMnmMadVtJXMLmzigQ1Pno+cb87Dp8/AgBr/+Vc
2m595J/R0Hj7KF0HlROTIlgPQBpulnlafJrctWSxW07IxxbS/F+J+s+Unq1ZhY7S
YIXnknm5haK9GvDnMXzUlzRpgsu/GR93OBuToxC+BMfmD86XwaYDE89SqprhtYuW
ns2YzfhAugee4pI5TxcliiN4l01LWbCqVVVDkF7tysvlQoXyCwW1SDuYxkrJgW4X
VfN6b0nsauL642c1/voHBQ/U3S8qOS2piqLjqOhIraN4meO0itFevTcoK91QDVib
5coBhmEbaVlldFTSjJKcgkFGXSBdwaM/2qFLr3RB73uLxypgJQbp56K68ZGNMUKk
lVl7jNsppV8GCjYUlivBNJGt4kXcVW9/nv2ZTRijce/UrWhK1kf+AyqaJjObZ+rS
hA5Q/GS7maGpAuUCbABwMxetpxlDzfiLqDjajYvv5kHFOOfybvfjgpAzo9SDKr2s
yUfFyU/Py6oNLOQerx0gjDKrmO35IpKKhmmh4VpSUp86pvxFAyIKuGUkrxiTEmv8
ud3O3poFuIUAYt1BC9PoaphIU5geEDWi2gTCHfhrEHZ/OOtoysOoDbYYOMBiQAEv
2/J6qGAK4No45dnxwDDDMUmVjNMzXulX5E6jwcytJLObOxOAj5pHtyese6+o2uSD
WgEhmdL2UhGD8o4lCBl49nMX36CsvpfB/0dMFu1MGUDd0Dr5dsfje5GOzsXkoxWx
0enH4rOkV36QP9Amj0EkKKMigc0rH/mLSshQL5B33DglS2RQ3+Z/JTh3VsZYMUTQ
2lEpqlJKWdwzIrFhxdPplTcQZk2W3JcdyNhUSJBKopRIfC9LJ1/rlQudECWjgptZ
euaQRyHXYWvNygmjmsEcgWgxNPja+bqZCksyvEi5+k8nZjJ7hRltcfEqCy1e2t9v
hEu/5lMtbqajvpSEafgaEfH9DKnnVhIbn+fciGl5wQOUsnksDpvNV+hwISK40wFw
RhTWGmzsF0GpP5Xb0KDiDwrHC28pahoMci2AWaKYLLF53uiZRTDQAtlklr6GUP/P
RE1HFx0oPmEAYRJZswnUCu1MH2zy/DrR3eoEAk4e3P0bjLa6406eJE3xFKyi8zMA
Y+q/OwZiJTxW1m/TXsK8gYFLly8RwuuDrjvMH5krv7YaTpwwTiZXLXUyoQdZiPrp
T9J1/zqPFqSrbU/AneWdg5AjI6aFF74vrkqDrtHpj8Q5cyX5aQvnkq66ERQzCv9E
2XDpgQeDNKdwnbdp3XGHaubDPcP6o1iMZbGSfl+oqWRnZA6LsGyIKwxmJcsoJrCh
ORRr8K4GT+eUSDv48s7yjwGZuxmabhYTRF/EpefWLzm+0J2LV8xRfdlEBCmGfmEX
QxYkzACXSHyg7rBIuVXZ44BZ0D5zUCGvl8dyCigawPP3jlnMyl7icHtIE24kIMSX
EJ6Kr2CmpkFhN7dGvlI6qxE1wqA0yMw1HRHmhZvEUp1KBIfTYdVj82WqZQec1YsL
+6bSQdlrtmNUtlWtt+ba7cfjmStvlQtseOehhQpDj2TkUQlQWFlV1bCf3aFsLjsg
EaQpoSb1ER7b2uwn9VdJJv+6tGCqSC/kW/yV7K+7JihC+TO1zbwigvVX8bftDMcP
9LsNIQRvkbNK1KtsIJ1QcPi8/jKD0lNIWBglI0NNTwGXqbhmNdxFSUTSaOSlNFec
KTcsWj+53vjjJgWmjVdc6jHeRl+v9qLcvWw4E4ZPBVoKTchl0Bnte8JrsOzpr6A0
PD29MMEtaT32qhnlX0mp3uLSsCmKJMLGBftyZh1mDLQR99z6fzLxf+rJH3n3GAcm
qaeDWt57Jj+9ezcoASH3Sj/X+FxL2AnqZTXUNGykLGodJOz+6ltEazy8n5yLqFYj
NUvNn6nTPFGf/IVvLKPXA2HEvIaXBXYoE+iHH+hKNlq5G+r+G+NQ1vKg7EXL+Cpk
6SHWWmf8rjhqEgCJi6v1xpY4FwY8HPkDGqpom2pM7JmCIMS+o67tclkkBZGBAdlU
0OYyfImnok4cED3IVDulTaE/b9fZA1UabUSXZv/pVHEy3pWHl3gZv4sbJ+fIEvIT
cb3/ccjYJQdsflbHn39/Enra/658MW6SITlg9LH3KJc7WXLhgJsjvsohC3rA04TV
kvQWPj4OCIrkDGSTDdZiS9iqQusflYgbIxRtbUi3r9S1MkpZxH2zRIEtq0V0/0CN
Ibp694QGIWnTZinCOPUTGFi9PjIHmZ743yawEiY++dZAqkDmWX2goBRglPRwadIg
5RGnyOATcKTUVVvYswWd4fbUvBUpKeITeRMfzj0RtQDiZXq2VQp+P+6up6wNZEAG
rnaCT0Zwmu1qOBSCnLgbOMKZxje+IF7DP1+m4qXHNX/WpbFEvkEDGXJiXCqHqRvx
T6MROlBUT5oXkFZmg57Ym6wjNrO59tkLdK46xEwcfz4GvYCcHjSApNsWwwSHoV/r
ceMBWsCdDuoI8jIaiKBZy99TIQnFOn/Bg48wi8ktybZe4E+NRFcIcbKDE50Ga4J7
UsqkwFjd3q9ZrmioFWCs64g+W0x/OUaocKWNeJzNfaenGrCxcgqSfg1qtBi7iLcj
8boilXsXjzBGcrUKZdYkXg801d+468eDUnCz7qQ3JTdQ3+E7eKKmBuAhaLfvtM8t
yQA7slHSCmTSkg+9WlT8+dtlEbiP04aH2iWuXRdpL6jt6jkE+cH2Q6d+TQ+WqNbi
Cu8CPX6fd2/9EA9tHl2vN0Fr4v44+d1I3D5W+5cApjIke62XHIFjwZ9/EqKM8UyE
n6dlmaKFJK10niant76N8wx549XsbxYI0iF7WtzbBinS2NQwLmoOU/KAjL4IShy5
3fXsm54d1Wo0e8N+Eyu5bkhlCK2NuUOxBM1Mqz4PsdwhLtRQGAcsvnIaGg5TpSzl
Ugb/glWZqJEZukRt3//vWX9LV6XCREmV9VoI7S4fyZ67UoJP18tDKxjNlISRsyY0
ftCkN0XsJ7wfuFuZTDDQMNJccF0ur/GMZJgmgB3o0WSz/Jd6Idak5enuvJ4EC8Ct
17ZgvocWRK86bM98BemBrWOM4Ax49ZkmTEsi6VLg0Li/jQNVGnmiqg7frgTetm5a
LeJWgPcQBLBIG/9bB29KhHQzAwEsVgt3Kk+G+CA2TiQkbWcFWpikpyflm2O+XoTI
tfFz5Pwb882pCaIiJTv3HETrA/zUkvS0aY0sSvcK6vVSfTUpEmWjf4ocCUJsbl4S
S5OjMmzVyqiFJE1q9oCF+NRDV3vdoDkyaLYP8EBtBBVCESoo3BR4MryZPsUF2Vcr
y0rrHYn5BBWutrsKDYowoUfgzWfQBv03n8+nvBZ0p+CL5V6RacsJLB7uBSaFy+Y2
qdHzU+1BlF2S3q6DULLMt0Rs8nO7WGDv6xprJDgu6boDBfO+0AY/HdxGx9Oef6Wy
tBCN0NmySZe/h0wKpz2Gr44FQpPmW4wnnb9jYBFVh8B/gC0Uou0+m1l2ttzEUYjD
a9kLNcg9Lfntxk47PymrU2Gl1aI7pV1tX5yfMVgFjLQ/4mpxDvSAGHM4rFlnkQdF
8iIeN3QshWavzwDx+ycNP9jCKeKjAdadPkKWTI3v5lmWkaQ/YVOtpQqOYKKP0jDT
vdg0365bbTRTMYuJ5iDyF+PSZKqBOI9yiQo/RwA43Z1nRHEPnjqVgZ+jtgDvHq+0
KRK1YLZvnyUDxobV6RHBe8jPXtPm3a15qB6qvpkLttk1kH5oJrx5loujR3R+dlyv
I7GnIM2mksh8wCQqrfDW8Cgd2ojP4C4oal7aIRwV6ejYKG6fAwn2SursJszNMyVY
c7hOa/myFJsvCtuBN8onJ4SoWFS9GSaHXM+vwaX9Mxr4lVdMjh7shvNRw7xmQALD
HpWBWyMil1LNj2t2iP2urZCYva5RtA55vzSgBTqd1aBdlwapPEKhg2JuLm7txbVD
4kCi4wHI6yweFMbY9mk6BunWGnkmuqqceC9/i20257AFQhEfpNhh0SctKawZFrKk
dCoOWuveyPGNKsfXNiKprFsFNOOqkujmzP2KVvZpTTUa9LygCKeKSR6Bw1N/6aXW
BpvenEFb0gyn55tMqhY+BXlp9y5IcXotE4p9r2JqQ0ySMCI6hNyWk8MQBM6gwMfg
nAIJQQmMVhNsSTvE5JMb6EdmdfXfV7RxyOhpq7TrJXvPfWOR4Yc9urkWOaJn8Vlg
YHA8PK5xUV1KYSdsC34Rnmhv4odsPcMStxVikrSywHnyf+PczpGi97lgmDvBk8YM
JXT7fz7tAgTeshIQxeFBDQhBOnd9UNO9ImoYNbXAEjPW8CUI8u3POqRVAAMffqSt
/YkkGy3Sg2HgzGoEx/tEVw6Uctsx9hqxYoDXeZ+KiiZK0+giagk2fvs7CDtv6eIN
deJmEFmwiOfX1dD5wUrL41JZ6aV4wo17vXF3rtr5F6+LrXBdbRW1fuJDnxgSPFoC
DgrkdN/3jcIQExM5C9Xmst0pp38j3Xe1FjAPS84uO1y6H2eMMcAAoRxKq3vp4OQ3
FSGU33mA6tyBIC6OhpntYSylo8EsVCYtsVwBqP8j2VlkJkc0bS3WGb9QaWx/Cmw9
Y5fgIaTs2+u7T5+GqFo+bk80tnWSd66yd2n9+EchpMp5VBsMNoIqOZZTmnXx/WLT
+siPh9L2bhbw+XS68XMz1zWWzTu/9WPITQhxeaaD2dWIahHsp+sIUdqSewT+zwdC
ZXe5lhPIcX5Z78+5t15h4bjVIkgNB/gPqNGkx2UAPRd0H8acgDjQn+WdK24mQ0eN
0jaMHhfvw4JITrIjr1aDxYvkPt7Uo16IBGSzpKh2nR9X5mVJeFMDDXhq4PeAkwrv
w/even1YTAq7UvB1QI2WwDDtvnGy/Gg0VY5mCA12rzVBEnh3QhvDG9EJk945/qpb
tjTQD4ocdpxTlzyk+jXIZVq058Jgfb7cSbAN+kFfSVUbyBIcvALjMqOOfdEr/0gE
z93y24tCqpLf8MW173G7+ESxMipodQjPHE7/gL/RBra2EiUq94b3pm1jFTlJ90KK
7Xb7QqiVcsf9Drg3BReMWgF8t7Cg2TQzrjo8Fpt1ObJG7oJrBA13CzIdO0av9kZf
1Fl8/lPTF9m2oIi2zhIQF0QVlvfxxOCp1m46FYivgfMB0g9dSwmyrblVpL8uZCiN
Qb8WlPqo+GstZ5mp9cOS/wpMrn8bAmCm9jSwrgs7yQhzkMQ0nCzu14vumK0eAJIF
+YftPVntI+V5VAYD+ssIeuB/Qpsr9BTWwRQauZfOyRpWu77EXRNjqjLydYhy0SKG
bp0qLUCaqlP/U9wOXhxkb86G6vjiRy4bOZntMR1DDenc82L1SoF3u1p32AHvjhx1
W29R0pIzCRUFJp5JVl2f1og2hYD8GB8XLqbeOojl1qEG+qSTKyzwrp/sLSu1WsGn
waYITNlisZQQWh/Rz97rGTstNQ7VXQpAzaH5YIM/Xw9yNbeisyKygFuydXQhF44w
tEYlhZnqmTs55+jlqK05rUzQgV3B07xgk/RoR+giqnuoDI09hHRHMfC1NIEP2R8E
it4UxaqDltDOZCMafeHHIAAwYJnwpAW+/uFaAKmrUpPRRhsm7Kw+2guEAb/BSwL5
MVb3kuuIrjXqRd/FgXishNqPjR7gIecU/FujD3TJRZNBQ0oavfrZJbyY1VVmYUR3
AdV2ZuM+SFVyQHVNi5sWlQlSpdMaqWsJJaYuUjNoGw6a54aLu2TJGDuj63Z0/aei
tIIR9TgynQnt9geMcFkS1XwVgQxDpi/XH2ueVan4N2jZlcLcWGThvVPo1Lt/yt9O
IHJ0DzteQiudY4NVjNK3MhkDEmlBHKwNk3loFjn58I/YW2iIc7kh65SbFSTz2W0q
JVoNHOZXTSjQ+8waEctmGBgAa8CPc0sH8sy7NQOWkR8Y3cd3Ela78ueTS8qA4Ncl
lfV5jKNHdUYl2EG4O0jdDG3m2cL4SszqbuR3srpRGHKRWORsWUrm9O1S5vCa0/Gb
0TenSwe5ILDt/6kNvAaRQZgudd1QAVCWTkP81iTulu85g8EuEizixlTe4DOh9Gjl
I35pDlnRln6qPIr3heVtSU5KBjvU1Ia81GFisSk7uKB9qACdwUr7gaanhqALD2Jz
kABIdTWz55ZX7husmjwYZgNjaDeIoQxjP3yt6p+QcMFHv0+tYUD/AtnjwNjrONO2
Y5w3eTv44RBFCEnEyzyZK7nD55NtRfiSxJR6m7j/y5lVw+7C8EKyMXDm+IkYAd/c
ZuoTFdbC/liJxYkSPnnlEecAYId18ywfpAXE6xKAmXr2Q2aSJR0F6mIwkf0udm+t
NIdyCc3aBD9vrABXrYZ67ksoG3aQuzOhcLntxCMSyfFxB1AwwqGBixoaCPUcsxrI
Nob5wqRphFukpV8jYr2ugli5fJLE4KN1n1we3p8eLlXJVdDapXoioYp95aVYrEUR
pUxSgGFRk1t8o+zR4LW/ViVKfZVOiAXSK3L7BBk/hNC2LxbDVXgDpDBZlGJQah1F
IEcW1RuxusMZgh62xAP7Re/DWIzDUiNCdH4WhArVQIoU72OGpwZv2x+iTECCHOf4
NPkhgroaeGtmSdx+EkiMYTBppzWQU5hhG17nzepGESL4+ClQWMPg6SP05j1tlN/v
McyhJU3hjSHNonUcwu99HmEhJvZW9v7m6K8fuug3ki9+wnY31WzgYlDlC8GztZaf
MknruTo0rafeUYppBglPgUPnwV22l3Z9ly0VpBh83rP65NqJuGl3+smdERRnpwXT
x3eIqWYvX8I+OaF79TX9iZ3vXZevczjkTiI2B1SnYn1PUM6L+xbPEAysePV2Iqj+
+T4tnOUcpeDrwO5dK4sY5XPWs3OsNKLcYSO9yY3LHePkOHKauKBkD1cvcZNqXmyJ
3aB1psSIOL72NophDPk/lLhQehQ1RZ1l5Mk1Cc7uiJ6ffc0tCBKUZuLGBnBtKdfe
JwSeYTt58+KG+SH0+YXZtDdcxFRkx+5IhjsIXulkmjvn1M0OQv3+kt26cv3q5Ck3
uUjdOHN50nNNxt18Wr7mb6qGD6AL6LKDfrt6uSj6K07GPw8Iiz5Fpou9Dc2LrzTk
GbadPbfG0TLOb41F9Zi/BsAirzfITTlDItCU4pbsC6NnfS5ZMoVoHrwMgFdfXgTK
q289f7K+h08Hv/sLn1Pbi539JLg4RNLwzfN/lHgD0n75uhz0hq08YlahEr+B4Q9U
5Nt085ynFKVyUJxjHnvrHEBWer2nLpNGIKcIWhGHpa+9XLcQYsMgzYnIaFyUWqzm
dBmWHRI4n37lXQL1gwgHBOz98iuD2xR0IAnP3iNkrqhI986oBILKBlat7ZUbujjd
CB0HUqMWCnvgy6kIlSedIubGvBtIVTJLPKLC/pJaXIDq0nL41qWcHbIft7LTmoyh
2ov2ZG+FgIiMJURil9ytU/Usd8s2MaFe2pvAEyoVPg6l0Z9qIn8maAZ8fKS6flLz
LuuTcM37jOX979X/EXGFP3CKYt+GZnujGVIQkiEzjozcjr+9Y2xToCSrVFgZWQht
6KTzj2ivJFaoDdwNZMKic/2/gItiU3QbemNVfchMaoTuM6q4464pWVpu7WfX/CFs
Q+vVdO5l3trHnZdB7cEVuEeyRZrFK7CLH3hR6s2U8z85S3+aEt9gUDsUAEo5TQ2h
ceEPk6CtTMfpbduE46Oras0YKl4RJFNeLfv9K44JAQNgyXravekz71mQDmLcHFGq
cn+VFs//685nwAwjLkV9iB005PUkPiYuapP75u2gYwmhop6nE9Bu/yOwsEA5hByx
NGqXZM6TYAU3v2yUCBEct78/uojJyxm+obVzxE45RqqoJLI+fhkM2gDsBJDd0JIa
7w1SRVEgVVGdgFLy5CDIrPaEkoYq9vQRKB8WHZuDKFke+QUhzheP9dozfbmjAh+t
aHzDPxaVemlPREst0EPVRQhcJOLZQ2C1a8HEIZ5yS4mLD1RoHFU2EcaoghBP8/Fv
p1n00XPiYsgIzl3niJCZSy/KP3HkILHTqK1rJgJevzJ4dAIF/TJiEkKHpf+NwSFn
4EZ1PkEIa1NWM85UH9aqndDVM1Wb0q8lp1yLfQl7ZiDkSRABbZaX4qdUFRaPHmRL
QuGtFlj8AvxFb7RDLE1M5IrykZY1c1eoUQMbtFVg51YUVlb4c50EnmLeCJ5zBEhq
qatcraxzFrJV3NsmkKN3XDfA50gcwQO6EprAdo4pQCt6nD5jKpipS192ZsR+8Qe5
GMJv49sNJnr/K41+3GEhqRoh6GHbXAX6cWBsDDVpgZntTFgwrECvWOSrfrVFYk8l
SJdqFVJTQN3Ltj6HNxCwI06ZCs6nAFRJsKgkm1vbj0Ypna+YX7F7lYllxwrrtz4f
3KQjRKOU5YSo+YM18JlAlUx7SvrVtldLUne/jXfE67Xmb13yG0C7oGVifdIe9oNH
aD4yLLRzSUQ2eXEgXDn/DQURDm4nKM4f3tafAOkLeHMvQ49sBZpRQh47vE2kiPc+
wnHwbhnhcHjsdscrJdr602uAMvPSITvxPMeMhUzv/om+clC2iqiuzzKy+nOe28Gw
E+CmOjGcWfkGruHm3yK3LOMpULF3euS90vK1fqebADDrd+HfHFlFRIhYHN7NCxPR
8vjH3hR3stULgiGKs3YDD4g5sdlFgDG6NPQHDeIrwb1duPlbCOuGjn4WFQcuSWS4
tCveI9rpywqSiDv6Zp2X+ja+gXqAtXLP6kcm5R1hKYeWzBL+qSPQhvEBEy2cIltZ
f6ySdI2kgzTJlYVYIYZrilIqTQVHF6Lbj2xaIDz1hI9+TwIwxZkxRdM1XL9gA4z+
JbRa9lreTDaHciB578+RG0/Lcq6FxAzsto2c4SBiU0V+YSVjor7LgiCzI2uu0F/w
T05wmEpsurBRMklUfStEA5sajykLQLJTyFL1EI2LhM3lnla/+mUK8SYzJ+Izqums
D+9RI6wRFf0GDHsIi/mykWSaymsCEyvwleeShNndi0yaQGHxA1wLXxipjWI3kJaK
+aBkfx6yS3+yPX/jPnwFeXzwxoaSv3RLiJVXzKYvi2VL3s3D70swn6Fli4HVXSrl
exO/0AZ33rqTKLQMG9S7/S6M1rwTgxioxUfg2MbMQEqlobslKSVkuKTD62+IO+KU
Pg8SRlwzEMKuGp976o2iqzpxtzXU+kxO3KDphrtA6C7kMcW1V1zMUtpmhQItDTvN
+p70p/d4rkoL5O1bcamPcCG3xeoByEnG5H3ELQcWh2H1feUro2bpu06s+GEjHpZm
YEihm/nCU7j42s9oXFiRnRY2dRZGJMKAeAp9FKOQGAOkd7AdTHDeTWUld9CDAxQx
AIQcM2S7PKmTkWUID9Kfpls954Jo+xZDsrB+yVNZbtxYAGRGGQKeJY5hgjrgIpps
AsSI+nNqcpzn5pwh6XK58QxjIxNMWr4bc/FKFUBOYzxbbLSCaIjMf+zBzUkJqQpJ
ILNZl6XX0Vh/XgdTXnoskuE77tcubJKy8rzacluehjyMms4S6Lk2h+oVO3zI/kN3
SBIsla1ptzPm8ZblZ+7Qd59JkoUHF5LmoM2NbsJ85negowV7fMHfyn74DgzpX0vX
Gv3VS3UfWsUWe5JQdCyePFG8zSaJuWcLcEOeyBxWhtfa9xw8wHxsOxu2VF8G2/3Q
iV2LOPb+kQzgpv9DqdwORyQGTGZHEnC537j9pV6J+XL3VzKC3fNux09LIsqBnkPf
GoXpjNnUshYbnS+unhUBEK3dFN8WBwjFQlpPbItdtOAxhfYaeu7BPYWTVnT0yg6Y
e4rqX41aSaHZ5NdFRs6nE0MXFslwgq9YND/doPPUlHA9saeAvAX50JkA3bSCfyt5
WA/FxIbrPIS+S5NpwsgyGqva/h7tRVF9CwXSZg+1vlwAG6cK1BbvCXFZRpOp5JBW
XWW87o4bIrjwrHYtGcC3ZfiimXXC3bVJcnmDZLZt4X0rwICjuw0sGVDGfU/KuM5J
9mSBS1wjDjwNwFm/hUWTDAwFAI4ewCmvnXkrhsXs13pRMzmPP5Grq54XT6AYfEmE
5RNuQJgVtQtcYM2RvfnyicdpRTRc2ka30SLUtXKWolOvf8SCTN2mu5lMzBTPz4HZ
ztMtoaFG4tsStb2HMzHeuJHBhKgsB8gTKI/qHWtoFz1D6P9CtemfEHlDP4JSaGjo
Pz9RRkUTlj5nxeu65vMoKvD4Din/us3tqdT9xOu5ki/HiTMx7ZkZ3Qnz3FOnTYh4
YzbgieSi7aEL/Z22xGsAmMi9qO3RsCLjV6UR+T0MwjctwcH7NoWxG+WEIGsOi0Tw
dlhqg0ozpTmzNtDgJVJRa5Z3wjt2v3/9RsbpV1bK52gCtykLLuHeReXLUetDfHtI
HQT6diFrZyw6d7L1gdKCi5pITqOQEm9pYr5ZVmC9QeHTgq19Tu8Js82xKVzJ6nqX
lx7H6YMBzlZ4OUTsMXSoORO185s0sYdsMcm4SMnDGXW9kIll3GwVQ258bMWaZIDq
D8Q8pOUSPRkWfSuO6zN6efvIRJGQkc+IZsg9xuKyorWPLXmGPEigCBPedta55xmu
uOR8QNJORseh+42awqu+G1F9hy8kALKtYF9weNfA/8dT+E19k1fZtzAO+wDKIIvY
d2S8BE3Yxfnotm7OwoAyGiSQt/p4I8KFGWIU2MuVpm3z5k570y3fbX4HhR1r/uV8
RK3zVUF/ZKuKYXed/E4wrVFod4mj+R5yhqlq6wzqZ0Y8/luC3RDM7EHyKX2P93EM
OeHP/xazdHn2IjBvR7ipU/PsztAj5RsZsUMrxYH7xJuhObxhBg7EpFKVFf0ZBslq
7aScM9KNnmT6BS7nl8IOckXM8vh1CTGXO3tW1pztQF8PFtrz7u9ze/wyo5Oo4zYx
GJPeb/swpJAGYeO7HEGqaHmO2/CNh8PCQxiKsbLUMYbBmZUtR/0tBG2tKMxFZe2K
0illiqpoZxu4CoG83dh3EOoEzma5GeIlPXLBf2gwQc39Q/pvRQo1dsfkhRvLGVgf
8ftOCa3l9SJ4sFGRxTAinH+dTV2eql1XSZbc+a61J8uhHF2rshS0IaVuFuQScOEC
UTwNIYsbn01bOGiA+29XUUnEY9fnzcKBwRlx9xTrUr54T35NdBdZLQvXZYdkD5y5
LuTfuD5fPJ2MoYZIC0q9wmx9Yd0uMG2c5UuNTPNrYEivAkx8fY9JvrBKHqDbVRWm
RDueg5Vqt0Naeh/L7YmLOo7l+9nVIGrGy9zZiu9/RRF+lnRMsZ9MP/2I8/V1nM7v
9vPS7g/FZoJ/dn5yHirx5/z9k57xcfVW03Ds1iajMInbs7Cq4HWzMn8hrFCwjfFm
nO7U6b91dxiTbgxP3ryVuNBxsagX99HG40eZRvpqSlns9yn0GyiqkcGcS5lqc1IK
blndArvySbjXjakZvGxUYxBMBwRyDM2gKADM7BA143VOdfkeT7ip2d5oq/GSjQSn
QddF5HRi1Zkhw+nj1YlIoxG//eTUWeMLHUaU0yYUG1Fns/aXWZygCvJ6rOK0zD+2
ZmAsD/gUQ2iyujV4IFtCfq8bWp6pGWSBkRafluoAKiawOxm41v1csvxj0QqZxMB1
PQJ7K6XOhPPTzGUjJxEKbIOMoN56OLR/CBfWxidK7e1ZkMFSGydGG672uD46C1Sh
545yhFRa1feCZkuNRHaBOfk7TexNRk1WCe4wOpVhY66xlEUrCufFn17j3Rw2AjmS
6hhn1W9cU5wSR1+1uRBnlfPTJvJpj8UQufzbWUlxvkBTBCVx4usRd5s6gOOz+8wT
1Yqd84M2GAh3NuHfJ084N2syQoJww5n0O4p6L9caNGGepYSXf35KQA1GmJ0lhP5B
Othmc3pHj/yOnDgLX6fF3XXBzJFyJZew0ANNj6ZlMLfQTn/xFHzdYREiD3p5G8ho
/Sg3B2dQKiWwvjkFHZvQp092itdm4O/tvPBPkGXAszatSpR850wiAYlsiqTBLmgi
lAeJ6m7RH4V2cLi6+tHxh2pgk9Aolv/fzAOabEpleDKbGJwFsbsgEP5pgPIvLfRM
OpbxhbKBiPxGWd5mpMf+4VXiNoS09ihWc5ZTbDT/FFaDX3hehQeGJYDS6Or3CDf/
UCiih9RfiXo+xebJaiSTB2UojrWY/UVByrTEntvuptXGXGAab7/Qulu62bS0iTtd
EUkq6p0xNKgwaZNLFK2CH8SastBblpXN49zqef4ZCRdA8/XYiVMOuLhMvXTaXVB7
pYHCpqFXlk0ovEZRHkSrrzSlBeWoNAOJci3ZksjOldC8jRV2ce31Vbn4LZHea1kQ
l96gqvFsCabRrYZGDlYTI+AOZC7smuSHbl9aamcp6N2XPDvFfeT5xz0ErxOnoWP3
anCNk7oB707IZ1+idfDteBovFcQzSl4NC6kCnsXwkGlcM1wZ7uPX8oV7mo43UrJQ
hYCW5WDWeGciNoeiKE3m8iZdwefZ5nuxDeiFuycLrrZzZlJIlfUQT0wkRN0z5lWR
Uu5KJtypP87E+YA06xuTtCKiR3QQgNmpfUP4vA3dX3YPq9qHLwzqYPQwcbjfILsj
pj7T/BKF0KzN0ixcMMz/q27BK6fNG038GnLzX1CNbLoYNUPmCQCASq6Llxpl7sFO
CSOG/CpFPy1CSKbl/koDqziL/Qao0DrSBbhv9YcgP8EW0frzRjMQGa+PxAn1cjbr
mKKmWe8cKQ/1hRecjD7aMCxqXGQFjLnOxvXPCD6eieYRPQy0K4jg7K6Cv69/dWSs
qHExiMZGC85/7PkAaIy2/IkgpU5ZPAqX2icQjGI8Xngf37T25PhQWbF9ztas1cv/
rgSGFd8uWKfS3DUBIoXhO9VdZxHELHJ5oiWFtt20oFSgEGDMUdaX0OkDwfDMG+xp
oCr81S4da1EUo6peRDVoiwXDUOm8cc5BHpLNK71Qoi/ucZMpGvOO46DSJ0ZG9P5k
4nk59hEwDRyLHDv3qnnjCcwA7Oxg4lin7ztSSOlj6lGE18Vw77DV6RR8c01VyFw3
HHzapSFc3TX5j2xJ1pOLuZ7rJ78FRoKa/BAHvuwr2JnX/5H/GMA+CyIFDstTrhZE
6VkGE/pVO406lpYCK3+E5KWnytE938HkyuXpQ8bb8g5d1rpXW14upMkyGykce1z+
vmsSk6/qJ48nYpBnoFkoUiaM3u0E5xyy6G5TqKV292moo/Mdl2q0Aw8bCLS6duMr
9Ye8hb8sULVlVVXMoUtFdAk0itGmQx1ohz1LwQ7QuFInh9dedPTOvNtpD/4GJPKn
Wbk1FzJ11mmLWlXYAQVBhW6OEBJIjtipw5j5aSo0JHzsJlAUGnGC636fzweHBObk
zLCIe8Ym05vvu+yFq1awuOGau65hRa3pMYbqyBwAtTlKO4we83q38MArqMj+TJP/
dpQjfL4YRTGlodmNcVySByBj4PIHbibFrM9N5xd7rGMi/DcjzyuJ8SylUXxfA7kw
cyo1v11J/i3hCOpPSxab2OKH6KfL9VqVxhv9ihDhXV/GyKNWkk8qofz6yP97ChSr
Ok9Z8qRY24rW0Patw0kzvquyTOmdFwAqnuhq/To/uj1DV0GdAnl/uBvYE+YqtiwC
Lfo1U3XscJmQ0V1VlkbKSNTfV/s3JQ/xT6zOyAg3PC0uNOI1hWt5SLANr2sYp+6Y
YNpmjqss5Z8ae/G1UFg+fLoRB0egS10YJBw0PhYGWUiRzlTIhpVgf+X9e+2nNN3+
b0j5V2r5sid3KOmehJJTf3umtLOxLTdhMyZhI0cQU7P9cAhxwc4VqTyZx3X5lXOD
fFXyGGniZWcSNRqtbmjzxCKG3EBjTjdnZM6Bt5I5r72rRbAAyBh8ppl5eNfD1BXt
6EdB8FSQZpDVTr68MBrTaIIITed4m1fRtNk8IrUj5YFp5tTAePoiEnnFALiYEn9x
eawOm6Ug7gH5vVIYjOYWrJ/4InzE5VJ333CnNQ3/vMm6zNMF04c67HcBj49MNLyb
PmOk7V0lisLptilAUYBn4thWnirN+HqSz+u9YQ4YLDIDycHQ3MBj3q61LTBgk/xv
s/0d/PSgjEelHB+F2WfxuPGS6IU2vNs8LjvJFdZgLuR2v1MFUFKckcB1Z7CwRahL
ObmztLamg4Mu/Ub0y/qhd7PMzgwH5BDBADlLdmuERzzLyC1U538MCxH042OpoHN2
VvTKjCXPAt8eB1Zo3WY+1Wjngpk/hh7xrJ4+z6ioqHK7xVJU0Nq5Nqe3x67+AzxE
WC6qfRx8tc621cGNL+0W/5/5GUhdQzBPGDWxaRL5eghzR4N07xOlKalRZ4W8ToMj
uJPs25i9+zmgW129TtyHczr9GE2GiILJdG+6KJ5eRiEg7BozBAYipHhDHOfQ9rPH
UMNGxNJIGt5i7T+q9sB5M5E/leEdFZZDR7omjzckXvt+N7GVKbYP5wEr3ROkAI1w
uAM4s2qUXr7yaMpcF18KzAdCps+6BBOfArTKPM4/89sOESPfJNT1o1kme1RKrBOX
47UCZqG9YwV6AGc/PkFrw+GpDQTf1bkABdZbttA1ud2BfzXl/tigldgjsukHu6mq
sHx2cxwwGV4qtDIKw1gUx0Mkd+2ZYyP2oE7G6zUdEA7x1js/JCO4+N014wHRbn5X
gpi032mE5cIFEkcuEFmrs3GSIA6S97C+Yu26m1yBZl3eRnBEPwfWED5/cRQThTON
BW/cNADn9HNFk1ysJr1KB41cVooYlDzKglJqg5iTKh9SM+J9RwoHQPWnGwFE2877
CO2Jq9as4CuuADcDwNzvLDINIudqbVi5fGdJp1nVAg7dzt9Wprz1VOpGNQx5fE+6
F0eXxva5TTdddo2T3OPreN6vTlltzs8FfTlbJYdKldbIojYXxNGrBbp9GjMZ+6AT
x6qbKQre+p2mARqPp1UBNityEESiTsV+AJPJB8lVfJSzeuLBMAkt7RR2dmzOkHI4
L0T5ji+qOh1FEG7ZFxgY1JFk8HihFvmgSfrd+UNDeIKZTvMewahu0oPGnLTjLC4G
/UVpyqB6OsdrkTizzymVATARAx+f3CUROk+mj+9bFYCZLWZIp2DzhI7bX0V5vMz7
P1R8c+nOFPGZRPkE4R1whrx6ILD1JB2n3/a5SAfKDIdtFOB8Vd0ASCe9aEZ3lVLA
ese4ZTiTA0KmTSbBjxlw8GRRwHhcO9+pMRaK/jpNmg1N/+bDTiiQOgWvz5AyhVG0
tt3ActbeKp6GK6x8L8vKvkmVOhz1uFezlzb8tAU5+Hn5yuslwEzjMkiq/1FsKWUy
d4BxfouRuPJD728zyaKqXTOsDEgRuqVAyfoSHb3tB8u+oSUawYsV1oCMLAW62VcU
D6SG6Q8uPN1WemdARG27rrot1GEQTaiA57knwiQZZayrtuyJeFk5C/fxXT+5kfOY
WM7KGa7XI0fTj4Xsj6vkB6NsfbZ21tuQI3VlrEMXfgjG7ohLJ93GFJo+mXJ8ACCJ
L8Uh9KhewGSZEjEkTG7XxzPPeKSWg9zxLmDi6q0HfGJMf8htHz9MrgUL9ot+newX
jhGcbXtNJYpTftFH7KAKt6wqpPXYw/HBTS9kyQvrawpbNUgo7lj5YjTNwNZPpRLU
F0o4h570isgKBgC70nqXLG0kale7MkJ6To7mIWCpCPtddmSadyOJPCRJU97lpOnz
MM1yEbbKjXNOuuAO/JKJwVQd80Ypla9aKslNFmNRJSFhQpRlLkh2NQxgD2L5AG4C
NvFCshrMhPTMu8sAMEsmWyj+GryfJ0wxHVuskBQImo/OWTHFrHt42dWCeZi9JT/a
v4ghISzgoDafQgjLPd8ItGFj+F9JhJlA4vdaxYPAjcfuoQrK93dR9ua8/mIV6+2f
FOmWlNV9TGa13LrTxu3/zGs9AJGpQXcjVgddQ82fFs6xR8zEXhIK8yNuyzKeUGhf
2GuHS8YSAUBSfV8uhHq016nXBUOfIs+y49tyahL/P7Xs8Y8UhXVezWC2yl0OgvDG
0vOvo1iapiMOIPr4ZKbcLAn+Wov6o7uqYI8sp0CdWz34xzAp2WDvSYuZAvnhfCxG
P68wBm3gFFNb5u5iYyhq8GbxPzwqRLQf0o+umXVN15Up9OydkpLiv5hC48RVSmGX
vRxh7K9C68qpavNQ6bp80U/dJ+pukEfcwR53xNuAELDsDoqZ4AhXGCmferzUDOjf
GJeKkgJdHA9k5r9+Ir5Om2Kn26cj20lgUfxPqXUls4RdsUF79YXCdUpSkzXiW6eX
inCtNtk8+9kRw8w2aEG/2fhX4ELLAHNtNrSk4h0AAH1bIjJ4Ko03T87SaI2mgSOE
EDkeHdHbCeJ+6KcRah6aPIoI6emHTQZ3+kvTVJBxMtF0asKXHtoXzgsA0yZTxxUq
AHt4btR14WHM3nQxzlZjsFsVOA+3x0EXrxqoH38zLXbcNHIyzXCTtNPqM4MdAdQv
oN8vncX4z8Lv4jSJIU/5YckqcR7lYdA0Je6AvTk/Xu4pAUuop3Pyj7c9mmysVxbt
qSqgzrWyGECQ/zqjvgaW7XfdxIFzb+r07kxxyURQvUWBT/bTjh3Le7hr83RxPLQ7
cZ6ps8yVTJXpIlcon0BV79KovAEh4+HryztOPPuol/zNkcu/54SQhWqP6YH+Pvhd
Nj68xTVqzEvdlaQ4V7TzsB9TUB9dzGvjflIAu3p4qoXOKxGFTE/4tiJSLk3j3/23
tEJ/GPJpa7h79Q+va2WqCvQx8FR5q04ikkAyBS6b+poIgh7yrOAGRnRIyrZW3zrO
bwsISYHJMQCMkq+B0GS/WUqKy6pxwX+pDp6xe0049Pb0zP9J1+fVZfSOOoP/9nHw
UHVNYdtKwTNhu3SsPgt1mANN5uyWyrbTBs6PpPS4a1g2uJLOydXfMh0iSFHTbT2i
WnI+olybB5GpFPwQ9L/cu2gc1QQhfa1Ofd4XnfOEFc13w2cva7giaoDdbbNm5Ivi
LVmVL14H/aPgCnE7vgW6cOclfl589GuH0h9FP1bV2wyw5OCIhF6vLcz1Sb/67HGo
UscH25SPH+xDaMAMgBCCMGYww/5SCmSdwZpXlo29HyoNRtzapHTz1snTGEak8c+a
GOgnpb02KVmieHVowCqETgGqJZY3MLqaC3evnQ5H6mRaIbyxdvg3+7FIRA8a7VjS
udQy3WDI5fykw+xnicm3ptNff0ZVFGTxqccA+QlDqZpzos1DZiResCykmxR10KvK
+3mRtfsdqQj2eAINUP5fwqIvm9SWZArK+6tp4D+Z/WeLaEc76gFxl76p8XOYWidl
nN+ZVg9o+vTVNnnrlO11Wc0YYPAEHldk4JBjBXlj7eAVlc29hQ0VXYD/esrrHQhJ
ROwm9xKSgXswHK4PQb3zazqeMUsqZWbwxpgYSO+mwV3g3wL3o5tAiJthzcPV30Io
xaD7Z7SpF+OGoPPinjt3UKrhV4CmGC8SAToOZ/iW21I+CsMjOk4Cvg71pFINi7+u
fIzwIACPtKshEgPSkb0lu86eudVVs64Gpa50nf1Olb5Fjsy/djj8kE5ENDKEMJLQ
nAQ/gWgqxi+EqVip7TylyfEzgKcTLsdCO/LqWsjRS2670lloetJ2FDiFdp+gy/Cx
7lbixSK+NXQqmd/JrKHVfdVXrPbFxW3rsFFsvH62SjhRfyJ0CWAUDOXPLe634ol+
PAKw7PD3rQCpvkSR9DpGnTAezmYX1DOdFBDexJt6tcB156O96l10v7mLim9/Q7eM
4YwXT907WxWkENZlBNFW6zDRm2MRMErHGz0fHL7I5SpFoJiWgiwaOrTQw8dEZbdB
FiX6HmH77JHfcp5tfC7C/JUAeK53eD/ioxNQJtNHDvA7Hxu8pXlfgV7IcWKGaPZF
uMFQHz/7ZX/y8YQYLihp3HDgLayGo1C4ymUASJPPYTxAdxMQ5LaliVFH74zNRjHl
ITpnM/LrhY6stAgUHP4pvji5m9v/GEi3brKsJNLuvJ875CGnuFnJ2oKjqKCwHp+8
BGNGyCw2Wz4+9lBucIgYPMwTEuGy0O6ok6LGU36MVYgc69IjvFumBvMov/zifwBM
Vy9clIlk9PpvGalTFQPCz4GkzClsGsJMv8n7QifAiQMVhU+3dW9enveBr3bCVB7A
Rh8Ue6zipHNgNrjON3sgLdMivVD2j8OG2g6SuJxOM+7nYPkgHR8VR2ExdhS70E6f
xuIrFeJkRYNz9gMRy3UNu9ki+3xs10Rad4jOy+PC5SnqfAHRY0Jw/PKulujEWXbz
CDNFdhvHl7y+AsY5smmge22MlZQ/gcwd4b4zZuu0eOLLic8TtBozgP6CfEs213H5
CSoHcftZYEAhKo7F778gT8po264EEMjzroOaEPcriQWwYaOs++s+U0z29Bme/8DL
bQpQdYLSceeaqguyQB7xSUAsAM2zGK7aZkAQRrruDU90v2SnZWtmjHu/DXLltRK0
y0/8MSL4XFWVb3TmYSU+mueKDcln0eQLH5BG2RcVmipFb/LB2iJfS/ptn+8G97K5
KBODFaBh3yyKm3h4yEeULnWBchjJeFaPsqS5Gh2QXXE+TGuh5B7cazclzpYjkvB/
MuPpEVJE+61LM1A5cxeHTYxMdQBeWdBsI3CPlFcAmMXnTiJtktm1R2R/S5gbH/8J
1Mhc3zU0J6X8MgMOhy0sUOO7D3EOZNlOBdPe3N0V5FrokV5eJSD8S/xFR3DNq5JB
W2zz2aidwypy0DJV8FbgrXgrzG24zwFe6qaqhs14CBU26X7dQMcZHyPd+rEDZDuE
9nTRjTWNml6EixQH78818h+TBHWIcMgpnu3N9OHiXEY/2FWt84Q+l2Y0qg3UIQqY
dGiUc46GC6IdqaKXhPfr/KiLyIFR/++/TCjA0hgjimuGkkAFyTvO7uN4dXpNC4mR
H/t7062FBi0MiLtXOhNEUDdSOuVZx43Vvme2u+6kCiA3v2Vp3ihtscBzihH6uMbh
ziKFuCVbRRSJKYrdvV6dBrOyCVkCIwXeU/F4aQwxodi5iznBZ33Tf61+DWoXX23g
n0ZjMw+0UPDzehwpj0IjBM3ArYIfeH9ZwhrqvvmAP2g+8/k3zas4ND/8cFfOnRD7
g3sabBMZR6xAWlf8olyt5Wn+RWr4uNXo+BROo1+Skn1iaxQJLZbMEWQUXknqvFDz
pEHDW4QwlUM2r/sj3ynXbM6fk1pBau3kkLv5zIewV/w4n5ddsXYIZnR+V+bZCPWH
OLSk8iYtaJew29LEmOVTnyDw/p0fq22GDTP90V4HweQwJ230ncXkiK7XufHwrcTn
yGCr/J2YzqPGH6uTYIDpfXAM+QkxXFrfhjSjiRZF6mp0bLBmPr9owBuGxHH7gWQo
0JWYkXSVJsJMnEAgUjSUNRyVvjNvWtZnhcadfv4W8SKhyhTBV2zshGMB5ze6OcfW
NfGxFTYqU4eBiCCWybhZGlL4YvL6y0mmRmzVKUS60JCS72T9aa0HDqykdjfkfiFu
7RMbCBuqQuuFM7VbFZS13S3lgBG/UNeXC6LkJam7Nsk4bTSuO6pxyEahs+ruQR1D
/EHU0OkpNaSdnJ8rtKpVHLwgNt0xu4acb1K8mkTXELSwT2ofk3qLshuCqLVJ9lYF
ACnbRuxvLrC5hXrlRzn0/crTgfjRi0tXrOYxbrpgm4EJhspDkCmTGCkOUAIzHpKS
ZniGnqv0m1UJdX6gGHiz7/unTjbc2Dmfadc02u5pMUaMUKswD3ReFhgTuBRZBZjD
GKsD08RZ2/fpctjw9h5xAw3klE+F13w7JMaDZPPsMvZUECdhp0LFoJCDqtp30MVf
GA62VUhdK4GLs+59UrDju7aujeri/2ThnNmE6ao9YcN6S1EZBoPs8E0Vn8QE0Ebz
wSsQHqFcriiAkRDR4f89NfxK2e3fGt3s92xPR8L1M2xt5dFJ/fZV6by0k6ouYT4R
bl2bFzfZu65xpXJn8+riNyMYm6kRlaVXWfvGxhnENFK03v82ig5cCDdr/Fv/RWAo
PN5tnFJxC6R32+mmE583UFVDER8tbBWqJcq46FMmf/+dCJEWbM+laYw6+ZEkmY86
+D7Q63MzxQHdUDymypUx3ehPN1LLgEc/dTrYfv4geP9Lp1tX/wM74DT9Vmx3BGBp
LrKRfuIy6sLxZUSagBwH9z3IFrqzwGdB+Z7qA7AV5YREF/HBZ2QseG0+ZjC+JGiM
qAWZ2s77sz0maodPPtLpb43PrktA4etYC/3OkN9DWriqLSp3YEmZEUPPBnmBCKLh
LdEXk0t+MxgoTeIlRDd/tZUa4Mpp8Imt3RxtmgBtuZLQqJNSXYADXn91vBVzA4WR
fWCUZYEtm+omq+qKZDV5UowtrUbxJ0x3F94RJqC20RllbJM14j2xPBe0aSZpOef9
i837M7q+IjngG9WV7ra+lR10Af2I7FN79xA//AI6YSIXlkbgFpPjGnxzRxelK0LS
tR65qd4c5PRtqpMdUs5XPwLDqsfa2z+k5JYbvF1/CGWYtDyv67E85+jlA/wOBHHQ
9Q38lcGUMf5CVsGO07m9xdqbzTW+5+Pfef1KvHuit32CPAj3nx0geDZ8nEclrT+Z
o4lH5TNGPt7VwXWpqlfKFIm+8Q4jKkDcnCt+Xjgf0RzHdLeol2WLKLccv9jHt7ko
kXwM80+7BTwVOQQPsRl+imsrFHkLL8QgOG/x99bxyMOp/PAGxLDBgVsgih+hKMzW
kGhDaRclgrOUT+zvZoQBEz+4HwGlw81xuEpVAfJgXkyk+/JrTDxnJDauK/I0mB+P
sOM6HKHd50WGogsC3DrP18qQNW/UeojnCBZHlbyeXQFG/eY8BhCmxKohmaO4TA9W
j+k6Gzny/QI7uZIl20fnTzLHmeXHsMqo4lgb/nuLfWUtWMjYHFuupD3mvwKs+GFV
StvpEHOSKSSjoHG/5iETXOQzC8PtDBcZMdTPt71KEBGl6dc4Ggy1+DwYg/It35p4
KDMTBdZAfKTeR4V30b9dxa5Il4M4VVcSH07ipzGGmpz4LC2o9agAdUtAA+ECFJxV
ckeNsUCYHwpzawe6R4fqKDTJcdm+69f4d2KOiiTH5XrWTYVpochTd6AJqIFBRO3o
XQkeXp+oDii1Ns1GCxSRwZG808Qa721R71GMvVgbPypazqFfqfIyoC8gWJ2JIysy
tPsMR/Cct3eg4CErovOKDVXOPmPLE8/YZkPMY8Yk7gqR1vkrp59hulGYXqcL0Q3f
PLv6OCSR1Gnb4kRT+4sRPpd6U009sW5t40UwHEHRX3igi6WEckew6O5FuxDUnCFW
B/8a/5hM8hDduwVjoE4D9Bcg/AisPUNKx3XAOKhsvvXOLOd6dB770VcB0A0CJR+p
Ad6eG9Oq34Z5RNULDKRo2N4o9ZwRBGT/R1C2TQ4tcAJc38jpA044k/aX/jPFN7FS
PPV39Ddz4djKfhiCPcfw1f6xiSBqL4VOXrPzTMkYeYDxxLydWa+MdgKL/fCSPqL2
XRv05qWswy1wTVQ5xr/qf2uTvYO9YvcukjabHiG3Jo3kuXD1vzqLZhiiDupPKAhX
RHjDhF2QcJIW/911Nbh6DSx9Fy7KCaTAzM/ky9qufOBrlElcAHsIMLdSOMKl6SIk
EE7EPBbkIQWqhUSm5q591v+nLHmt5QUszRrblEmaxA5nfpCKCJludCsq/ozk4s6J
XNi3myD9RtAXt3zxgJwZagb8xpPcG3yMHwaUtC9wSkCdW4TOlDpkmnxtzU873H6W
OXjmZKgPFN7yQIFodsdhUL7oDt4+BBU8M/4puj3FWeF4Pocsxj8G68C3FBoYH0zc
YR2PVJAchWYAy9QX0Q+Pc2nqx1H9rTWexthCX/eb6kuyhs+qR9shsNny82jPEAr8
0nGOqYRN2q5Ey3wU/SIdQvkftj2F1Ouj5GJEsj0kAd0qDhratlHoeFevKCTmbdwL
9Cu1+/mUvmhhg0mPmIJ6wjTHvmk/lLwO343nA3HMx4VBKXECysvTjqcFGyJkS1UW
BZpRtLpgsivdZzfOK7nueS0mqrW9B89zvyBgmleuO+ULeCAIxbzvJ0Sba1KS7Tt0
MyqCmzYSz4Ap8IiJQGnoYIJfxeI/317d+ReZEgQFNO0vhPjT55bLdIaff7wmBxUf
CYu2BcqRJlHZFLNvhwoOdXqpINTphP27l24SKacY8bmAtxvjAbEXeX3keKbiR0sq
VSpqH4koDNGRbT0W+vmuvvgPDRtSAhKFeLt08h/ysB/nO/l/tCvkAfI8FVef/USo
lOIT6pUz28AWOMVg0v9f/aUAS2ZNufmnc3mrFOE1A9vcgeqa0OuSa5csJjEipooF
FG88JdL45QawVinMWSA/TcERSGW7ECRWp1pCoYZwyulH+nhrN6mmuBkGJ1d6hrOb
NMp3pJBEEdpK9KfAfSXbo0Sn4QyREsfdkFKwkcks4wTByw+18r0c/Aim98BwU6DD
pbhVY7ZvvAa9bp4DvjjYcDwBVhRjHAuoq9ubAi/0VM8xw5ZTnx9RXi5vr3AS2yxd
fH6Lo+lQiPfn1L/huromrsNiQ4PWiNF+zzbGjLsvG3ttFo9yLwLwQG34Id39vUGQ
le/un21iL0znC3T2vif6ev9KRZG/83YgP84lKE9QYDAQxQXtAF4qIFOuDck77tov
SwQW+3N+IglOnuGoQy3y5A/j/FrxWRC2zjhnNwBHRcVhzRyNPJ6QNSjV5etMO8nd
CayK+8229mY5rRLFu5vdPusCxRfZnYnWSMVu9S6BenbGvrg9OFGcMCbmubS0Le/M
PJ8rhNw1KNJxMQGMAG/TKD9eynhkn8iWUQ/I7AtZXnMIOivNQOx0bGoDL0lqVEcw
nZustb2pUFZv9Wfi03Njo+cDuxVPWwtYOJDXWYKd/nEmnKUUXXzj6BM3HVdG2Lhp
KFUUrst6r0UkRKKoZX5/TbFuQ8ZgD2Hi+oJOVHSDW1+vX/mWAUbwXbIl2ry13G0R
JBYworl6C4ChzK+GedACCiqUTyvG/Jn3wXOJ/xl8EOAT2AjhRzLS8bG8OSiQU+9Q
CQexIx0WL7C3moLa9aguhawNm9A5IN0RTtea+1Ur/MEOYnu3R0mw6nbNuaGL+bYV
Olw8/qzGseq/qevsaaHfZZNvxC2ysKEFjk+FSdnNv6sUyFWNYnT+aWeiLHn9IJ8r
2yYxFY5H2YiocqdMLIDY/n4wams6eeHnaxCfu++NSDFrerHBDh5IvzWH1MkYlzfT
vrIMzI05MjiNOwRD3JSsqTcWg6hBVUt18SQZaEspycx8vh076c0FctMvtdQQ96P2
+Bl2wQ9EMigSzocmot1snLDRPf0alUulASVEmiR7EIsxWky6rLYHLI0Jox8nubvj
czbXVZBvTQ0NOeyGgsha6XZVjfQO9QRqNfA2+1Ov3AQ7Yi/zp9kX1/7vtfVva5ST
Hooono8KpNP9/6h/6OmbfVmWuv4osFLniFHwNNeYcsyZwFB87IYZJ9mhbV9jxaX6
Uj0lSV8Vr58YwOt/PthS+8lM99NeQmGQAPt0YBGVlVfIHM1iXgqEFj+t2fvBk2SA
Ijf2QwbWQpI7s+cTzPWsZ0xdyg5oJZI5S8LBmCQQ9QqnIsSXMiHtwdDo5jG4zWsw
4WMdzf4NZ+qf185rNA7nK2q8Dr3ThMWZSeApeRsObf98f9obODmt6jlBqqm+t10u
74iQdZ1KpaLrE1HVSqkUhEdc32LXI1Ao3bLeKVPIYpOyh8SSKlpVnwOAIy0O9k3g
4rNWCXQr20Cbml7l8Ab+7Gv2liB+rx1/a1RD2OFOaRYuoWDXtOcMELM6ORuAG4m/
+arU59zUlJyuuLoE0hr7y4b6q4afShGt+f6q5sFt6r2wyRntmM8DjruMfn5j4qBB
048hcw/XSBUaWer4ELQuWj68EUbWKnWgBrVM9nH0qCtpkXrMnDABPX3KizRZnSWV
BoDTjRA6jLHnW1BdpalwtqWMwdDyZu1D1WMjpw4H3xsBQrJjaFm3vH3feOubOy+a
+umfuNBiLDt+g/MscIxEgcZEWUYWU8pDShsQuj+U6Jk6iL6sIQchAp3cXCRmhOFb
wnqHHQLrGgBzJHeD/f6IT9HHrOdBFT63urgpj2DUP8LdkcdMkdH7JYa0TtT46wZD
8m3C/8QKAmP2ilLyHaUUOhyhTb79UKPz5w1damZHp+P+/Pjg5UBoQRYjt1c1hQNt
++bBjeCjYij80mIWmIwOpjroVj5DJS0yT2GCtjY5cm8bF5ngEngfNAFaQtMa3Ezv
dz+ng9GgxmrElSUl5BJOVzv80qEAlyAar88uk7+OA+x9gFSjT/Cg3Q/OSNvSv6ms
FNH9AD/BhdyarRx1rQyk/FpfvsH+zYLyOTBAVEj02xU2Uga40zWOoGfnmkj7d7ze
n0XdLD1FRNvli/zufLPSkESl2mNWrDoDDXL0lkYiKSUxQ37+KVKnkrfbvh6FGqTr
EMQGzQtGvhG89FyRIOgkXihFQNLU7BWAzoSPuAnEAI409dJ2k5uj9jakdyn58Qwt
DmwY7RWspXLutMCEnrg1vZt/hD5YSIZZLebnOfL0M/PXnArnDIe4DVfYmO1o3xAk
X8fD+JTQLFv5E+3BJCO3hYfeKnrYuQCifJHaUp86liQO9jKThecd4fEiKTECL2OQ
YIfqvy6rovJZ3HyPN2K7r88bJzeOB7MdQRKuLtfcQSUG7xeBVPyWiVfxirC9rDq/
uj0c+KGrY8ecFqCyLynWyatCronyldj9OTGyEBcoLU52tBKuatmmOfRFlg5ERgaB
H9r4PZNlSMar/6BzRtjE9jH8ExNw7OjxBxAQRnCThqNBb/Ze6O+AiyPU9bY4bHND
2vXMTPRXqKfcqYY3sFfkq1IkoFXkTtgYlRsurIuW3RZKFyM4MPhqbQKsKa1apiEq
fORuPloZvyw/A8TJMfDmo/n3hdvDGYipAvU7z7tup7Ka1U+/kRSxvV1t8Ssp/8WU
vV+lE2doZNEb1Ii3IvH9N33JPFGTwd7zpbDV1l3jqH3eRPwNeDoCeUNCJLisZl5M
njyY4MbfI47GZn9FcVUmUjBiKwmvbf+s5JG01WQ8k8j744m1bMYXNyQWBTeZT59W
N63U1F2Z4KHBKYo6t3tKsKK+g+LgSydfCARSQoL89PlkOooig6L3pRe169QBSjGF
qEYCcPs/KiqWKlAchJAfoYl8mSkZp/HYVMwHCPsVCtiLngYFz1jhrBTRbyUu5weC
pSPHnaDyXcNFlF4+HFvocebLUZ//EmXbT347HAA7DuxWkx6ix5+SZoIiOiKqZqui
uzwVWokeHIVfqZ5rcUq5gpuxb5nTatUfo5o1b4n1wyLcl+LvmWQax1dpE8VwpX2/
IdN4c1cop9CAPEFiHvX6zylcaTOsesZWvMlR3lPsjMZeUpFXizUwW0c2lUqBs+nf
mOHSVAacSS8RHNO7s0vfUtSSA5dZEcvUFlSnH4eFqFnOOVCEGSUoWzWptZLH2/Bk
WvVPCAHG9zpza0JBYeKDoxY7OwX7YIdM6PN4VuzWMgsBzybaIkWUOSQ+tjgv761C
q326+gAPkK9GqQWK1XKOKAewkC/aqpe2jeewlWFFBvi6ElQd0DKKzdmm97gfxJoB
rXyzwnoruXtwHJr+yMWo2aXBLmWDcupsvgBQOBaWzt0jcQT2CzkXMZ1CbRMhmh2f
VTYsl5YMcyMUFX8zT2wDzckhOkA8OZgRFRE/DP1B0VULzx87eISzifA0pp5OJXps
UrEPd/2jaVdS3OxNebaJjVmZDUdBrQy2Pwh5MxjWKKgvP3VhvivMoMvXbXYt3RIB
2bpMD+4CUvUKN8IRRIPpgYQ3S5NgOH6py/3Jvn67pIFCyC28CY8rSRUmVVwcUOUd
Pr6+7D/AiYIPs4VHBd78yuI3tPB1AdQY6mt/d6YWkuAyIgwWUboERS51dQVqdXWu
Ijg0DPL/Xz0A8p4lbmzlDYQSnwNIn/RUfE7nIBr3LKCPksGP0l1YUty3Mz8gFh5e
4sU15BwbuJAvhWjnzW/7he87RDDJwREHTUgJJFW72fThPU9Bdb+aPk8y0OBkSp0b
4g/ouanawMsSvmfR6EQ3DEqPrDgjtKHzF7EejwqIo3Q+xsmyBLWGL0Oimhl6wci6
ebq855cK2Ov79XZTPSPWcTtqZi1WqwQZVGmLo9gGuWt7AsygQqzXEr12514zm8e+
zj/4cqFJGW5BEvGoX15Rm+kWNhuJa3OjkNzqIt9CZhOI3IfHOEw5OgAE5jX9vPoP
5ZBE3Tzhq887hfC9p5poXaCSnb00KFuMScGGjsTeV2AIfQkotnOx4pTiQa3Sm2d9
b1HAFmnsrieCBkS0Mt/rIOy0zTl3oo2VFhwJseG3Q+XLu3Pa65Gt8NopmwXwuQll
2dTGFvSLv5ufXGAzbRoNH8eBaShl6gFqxrtaO64fykkc5mtJNRSplaYlYpLAV0uG
jUSkvU0XXvtUkk+OHI06oAEfQHqh8dQr+m0liXC0k35BqhQFOuYhFZ1zppvZPv+9
wUgQBhhml9XTdwqH3UrLkbOKHO7f1DUPK2lr/mdMTZoWyC/2i2rDGx+Pq85cTqzO
CqSK4ZWEWgSLpeFWA/BPP8/SvnZsqpTcSHnbIsaurSkbyFuyBH/86dPxicvVllm5
O2APxPNmFPJpzpKrXk7kzkgHchFyK4aRhjKuTQmRFz9HALqTT0s342bUUP25zUGH
H5GeiswVuY577gNgt894flf++DJfZ2K/mvZ647vlWQoyEjhO8NhA4HucdRg+gdAr
cw1wijhUy4aXQLSuqhTTK8J6Nlht/yajovfdfz5Ib+MC/oADJJQvbWa/toY1WZwx
MPCllQ2iREB62LYHwWfppQuWabOz3Bd8zBAuv5I2dgV5s1UCjA1fQTE+1k1ssTrv
qsWLuK+gKAgShbbQtIOvx3t+jWhQz45ux0cpSnXOR6wwoS7a+uuNICZRUykP9mZ5
od3PMVt9TEOl6Ey7p+OGAYYSm7XOKweuPSSFmJw63mQMU1oCvTuSmJVQyxHXb4bR
r2f9XYQq32q23jMPGoOawHHuM6pKFRtmPpvsTMaqFTWbHHxXyOiAVJz3VY7W3Z8Q
QVOZQrYz1g3gI0NG2YyJihk1DeIVf6qWsImb8bMR29C4YpFUtqlrrt0mej3jHoOo
bWtymHWYbr3iAkwG1KZJlUEJplvkv3Pin4LByNc67cE5Hkitd8VfuxjwZz4Uq31+
oXKXUchViJXQAoymZFNdoGxuXo76RsMMhQew/JyvadiG/Gldfl7rWnCuodG8Rabi
FkxlIJiPKSK/R9DwEFhTddjSsDNLfanlTWJ7Th5uRk7uDrHeAhf+pqJMnQ1QQD+Y
94qVxw8gapbT4wfQfaS6mZWncXuqJ94ba/1iK+WzoPq+bxgpiCUHjPrnGPbnnRHB
OAD0qke0mmEeYtmEOr7x681O/GwR1VMRal8pmersr3lJZa1epBLxp09RuZbTWlTD
d/ywatpe0hIrwG6yRXnBprQ1jHPngIEC7czpqHMZhW/uO1aBKxB2wT2qwtZkzUT8
W8GqGbytVsyRGiYddE2PrXg5XBtNBiXDqvw67QLG8LHwwKY/NRnHhJIcsWkVrp2f
D4dXgrhYzTchiVt5bT/8fnigjnGx8Fql/Jkr/b+uM1rHY3lCyJvt/mE/P4Eabh7Y
CALA4XXLKeykz8grjpV4iEu9pBsmPVMNbd+iFrLrTQuWUM/1XKNAMswGQtPgCw77
oDtHquEwmOOPdIiD0cZM0nuDIRQJrpjL/d/qkIX/9+P0QGPyPeqKcjVB3ZR/6DlG
JAeP2xJItGUXNOuzWpTBX0BU9Mb57LqFKRyQf9JRKEggYzfV2VCLE+99N3chZ84U
dSCIh0nBjSCKvbvmdVTVSTpEfBJCR0X+TISWkSnUkmsLRd8AM5gPOkI3/BAPpn3Z
kAEXm9611KmlOVsgevUSyQP+jmmNS5wg97koqWa8cOkuRhztOnx8IgwLPWNC+I+z
WvmeQ91GN3Zl9n1qHWz9HDzCvo8/8UTZTVAZUK6zJRnuaok2g7Pow6EMcC6fv/QD
3MLVSIJoOvNf2hrwG6YsuiKPna3G4tiIgiC5YTnj52zvwtwOzkgXBHIwUoWd8e7C
j7RtZHomAoxmlFReoscq0U2hOR84wIFtbI+a+vnBGXUJL3EeN0HsIErBgJ21bexe
6b3gfPfikJS8+2eKgp1nG7btBpy4WkJ2/mI6qTN03O9aI1+l8DayrhMPtEbisClm
44IiA/FkAkwE7sI7vvSudR5Qi56N4iE4pMtUVwK6JhRSImVsFZXU2BSKLcavF6VK
zO/gPP0CqLj0Ht/QkcRObm9V1gtYd+4WCBT985NuX9iFhXCDE9AnLDTF9nBXwxYX
FxePeOIFpsNGeZ53neNYC/z9eYqgIUecJMAVTBuI2R9UA/SmQZqzXW9930Mt2xNG
4P+a3TzrvPAOE/w1eK6wOqQdWUkHIUez+jmKrYuupVSP8hq/+8U9Stq56qUKUT7r
lc2cR2RRLJhmMhYDYYK8ZbHDxlUAIBoIQxqpVrz1f7sIJxEaAgWu/iSXsR8qDrJc
xsK4m7KMpG30bqXoWigiCmBnkIpAKkW5SKDyWrG370jKSwKsChlIM/jpq2tN4UtX
gX7R2NgO2grd+dFSTlwmPm0bBqzcKjNBU2WdGqi+OVZdSyDWcOS6yk3KQIN9WMld
GrTKzSbiFbmNtjHIgC4xoVVJUm6cd1onKyuStByC4ZlYG6bA2x1VBKtbPct2nPUL
xpKXQgtuVYV27Q+ui7C9AuvLUaKPw3Yv178oZbwPUKJPnNhQvaKUMNI+NUlfOId5
tpZ1o7mxXIs4QYqqhs7hjbz7NXNM5LKJgpEKLjLAgVeQZ6M/U+0whaUAd3Iixi78
f4FPVCsRNzbnT476A0Ov8rJxNJtuSjZaSRiDaNwGPnzW4h0O3iAZKIOX42wsvdDo
rB3YFUpgnzrGyMrf0Qqde4q8bWa9Gh4HEv1J3gEdOJUn8Wu0FuZafcQl57m53lnT
ukmxNRa27LP8gTM3WG6E2EtmQO4Yk9op91Jchgs6ndGJtx/3c40cgxNjf2AS5Yr6
XzNXDbhzGizuEOKwOExhsZS2s/GO5UG4jwJR4ud9wYOVQhLJ4P27ifPFXlDogVka
MS6H6GvC1uyaXE1JqcOsEhqvJXwlSVhzxz/8uP4WNlj6X2zifEeA+WdbXFZJhFYd
NxMwe3z6nvo4mNx8e0EGXQ1TBiH0yIO1FIgLeCajagqGkdkgh7+GEiDBFnHjrhUt
iw35GC3kjyI+AS3ozE3wG1O53lNIhmKLsr8OsKmy0L21BLX3KzXytdKcHf3PkU1N
3nBRk9eR91O0uYU1fPjiIPXllBBlttcZsrkp6mhkjjIVTswvK/UkLoT/YM/ue1RL
FWaceqCCaEAvkgdLsAPJtuK8Nf5W4aQIULrY5ZCbXGNAj9GB4mySLkMdrCKTtZ+7
PW45iWH8mUQdCTzPEZmQq1a1dn1DwWu1B1YLrRObrdN/L+1LBmTOKwB/pTOHC7Ip
Mwnspm24y7xTY4D9MOIQZQN0gLztZLFZpn4J83oONnhhs5LgZhVlCyzbDLzjNh2t
z4O4wrPpRl8XR29Oa21p5ukKy2c+JGXnROcSnBL3E0WSMn33s4Qo4obr+sqP9T1a
tkT+rrIJnEYqmJ2EFX4oswRSc0f+05a+PXqzQioR+CPTuJ5AdDEmJbhVq0QAr+wJ
QC8sLYJZUD394hWAhWNmjjSEPbaeitAtuQcmcg6vz3n05pcXr5NVT2PlaI7NczQs
jQMNdfVTncpOdcYfUvdOiZ4WjtqK5my++2LXcH4nu5NCp1ajWIlHNNaNtALXBWN1
f9NmRO7YQ1aYyRwmt6c+xTXN0VYhkn9C/lbyze4QeBkgQ9RQqQVCSZUgUFXXN00q
Uj0iMGB40WxGQp7zmg3n0yp16hszVcuvMTFcDPBvnJ3Q5mICy3SVXFoA8OT2GBMD
4LxdrpSYVhzqiC0NS8e4g5nXXfzylMNafTnI7HwemhYKCPK3HH9fdYg66/CfLf5d
6EjqtEAnxfQJ2BzUSYbl9l4sau8bu2qnHvpPP61cS5VoW3497rQLTHQWGu0zg1bF
zjIZTGFhkTjkaJonvWwPD0WOMaRJHg750aB4N459SY7XMF486AsxzBYdFnCaaprV
KB7fC2sHXZGqz5l9srUedKkOvye3VoQvmM1N5qOiw1Lk+gjYeLEOG7zdXMMe3e41
+miaKNHQOf7A8yy/fE/tg8spMjkL63uxveLISkYAqkVOdn/Q1TwxnGLhuVEA0/6U
3TkiDLrAdOTZAq7YP5unZh0Biz2axjRDQj5+OMKR9FkGAB89HHoH+h673+y6+pc0
bP+7EQv/4NBhP5GQKhAIx9OQ+iwXRwLO4QR9+1H7qI+bl9Z9jZo2pmqy5HsaxLk1
1OjUgQRR2x3Def9aGOgIq43+XDKQY9+VqjeQOkw9Mc0FCFOh6IfnFFBKnJawZKgs
3nYoUA0tWoi1esvdXu70E+mAdeSHgWpRd5XSD7AcDdAkxYN1Od7Seeab5p9Wvq22
j+vxNzMjdxEP17tFpPZe1PNwErYdy8LF3akiVu8WiIDHSgbXK+aUQk6CCByV36gY
IMeOI22fY3g27ee4TB3tXyqzxwFeK5qj9y0zZmFHlkkqIN4xEDWdWjtYKII8gSr6
IPxljFk6gHf4vVVGeKD+aU7VV3oB5DPiiFH8ypYECqM7S+pseFhnSd+jA1fH+KaM
P7ACx/DGpz1fMyw4foL3nkMJECR5l+wbMgMJx3569w6rsanBAezGozb5WjUjcJGj
MhAqNFSPmlPsz0V6Hp+3w06npaPtDMkhH/iGA6jLe/Yexg3WcKcb0MSWSDA4DXro
NkSu4rMfB8ut3MbSz3g1lGFRmnCDliU65xKNAOVUOlwFx2+dRntNMDPCmCa7Dtq6
1cbbEeau5BGjzGP5uBK76CUMCsA7e02y+sTEku2eMP6xyPM5NLYgo22RjDUrbELB
hYJ00mnX4deHF2165xHjG5Lz2vouWI11ynsty+LQlsXL5Ih+jWrnuklHDItVD81H
bO4pe3b5QPR0Iyq0of0r3idFqhQPOm5JcmDFrF8vtMVjyXu41XgEFXYnJmWA35Z0
SW9O8L5ZY2n70DX0/mmEAvXx5djJkTwrAPfB0WzS0V7qgQVifGilba1hvEzqR/xn
tj/jpFvnVbXjr2XvTQPMGK4GfqOnSjciO+lcM6OSRPOy4K39UiH+4+tcDvvsoHX1
83PHxE3YxRr3RZZi1SnfKP09T5FCrkbVxCqAPiIke7y4XgwueADQwK6TzsHBrlCI
BkxREvzRr/1Y5hFViqnZUzCW9A2GAyjssreUSROVYPbgeR4dvowhoyssyLqjuLoV
1/MTAO3NW0MFOio/x8TS04F85tBTudid3JpZ3HvCJCZCZCiJctPHeGndOpNgSsAJ
TFB2veFCCwKPHbL9G/Ex2ZePkJ7gSz3dvFrsbQnPGCKZvGbyi4euO8HTI4/nhgup
q2HmxVhYzPwKpYiBSEVB7Zr+wOnR/aeGCTLBM4wyJt8bbrWBlDm9tXLCVqTqC9Ll
NN5SpD7sTCh9Zt91xyRrGRbW/liKVEn3jrZd8VWbbCICyEoIvNXBw01jPOgEJ+6d
LlSixHCigKg8+k1civUIgPQmJP4T6T5Qy3oumACbLpdJXGjvD7oHi4xpI3xNkSGF
6UbeAgUpUlRaGDd4jG73/kWGSD7mthIeK0+FKLnPT283iP40+SszFtCtZNcv+2bv
+xyazxFE+o3AYJJp6gbQsyPTA6E4C7rGyDe8RiG4ozLNWy/3WpuAoXSJFBBuo+If
EZT0BRxmqM/9XGqWtB6Bt7vG4kpxd3hRAqJqcJWb3F3bLpD+5W+zzLDBDPTh01rI
nPOt6X8qZuyKWb4fqBaFPALQ+YN6ODAQu6l1EVFY1NoPoiGJ7xcDaKWc9lRTO0PS
5XtrRQdGU5y3vGOsZL7xvJA/Fc0PNr/VblkkZspsZsKMe6ziTuZdMhPg/Qmwl7by
hW31iIEE/zVcdJcoamuVT0Vc973onZu25b/e4avvdqvcOBnfNpG0IC3UZsC0xHcD
kxtlN1NB+XqHQmEmsHJD7MRITF7UG254ogm9r8xd4sn+Jvzg+2WKlLYEd9gO7y4k
HjtgWT8wMDuhyIBV6VE+d1MaS6xxBTqpb98D5XfnoxvqOY1Hr8/XdlaiE7U+rdmy
J90Nv0FtLgvZfxQEIeWASkpJnbxsorHaZRLC30ZtFWX+P9qyViCQSuBm96/rNTDD
1Pxc0IIdv6WAgBvBRi5b6K4d0Am0ep6JSLSlpaqnmSmXRFUBmTinAH0sCTYN31m5
pUXJBKI0tMBVIjq1kYyarhgHGdRcGK7YQyIOX6dQL3LTkW4Ia6M4C4cG30VuUJxJ
u2115QTF47B9DA5yOQRWu0tdQ57N3ZJE1thr/0My4zNG+PSD6VTTNusn9hpDsmTX
xvjqiVbGy9Y471KJWBiTd/48Rp908wU7wKWBN1R8Z80J8zWWDJmyDspyYHL7ne2s
VB7oRbwkHx01dqSPCUqowqUZ5z+1qW9BpAuHR1uzKFYAqjP0ErLg8bb+hiuCivsa
rL3fVrbaovrC5moYfSJdrC66MDACgooGzRa4nCz7JQ2eJVhPbiL25BQpC7heHAo4
cJCJ2eOY+si8OuoRFh1R32BovbqiRc6vcydJZtdAL2rMiECYiOQCNmbun/fuMZqM
ee/eLdydFnNtk7g6sbCwiUBGQ7rg9Oe/DgU6NYC8zaHfk355I8B384fgpdPyVuC3
5RBDoEbyGI8fp3HkfY2kAGPXODlE2XlRFpcRK2U6aPVWKYZW6UeYBE0SmWQQCzhC
Z5nijtL/1oW4tVBMDY6szijW9+sqX0k1FvxIJIDJ4DajdaJ+XMxyKc6Ll6iVslCq
g0xGYSi4B8cwcZWZ/iF7ucgoUkXrar1eFVi/evs/OJe+j8natAK8VGmzHDu4xLhh
g+DidOFL8XcogkBL61yghWzYNAfJlIHulBFnEG+WvpiQxrfOyH8awMGNjJic9YG0
v+x7fIJR2VIH5t7AI4+I0N2KVqWWq5Be075dgx28nHkalSYvMElkU4ayTtgFmdWS
PqnYDwmsg/mYFyMpgZydUUT0AFYJFqn4FUq6qYcwt9eSHCZh4S+ulGXGdj/lO9Ti
4Ja3sIxFDJQjgLUW6hkAVbYR0HlE0DYVpFz0wFIJ5vE7b/KrQxo2aUyNqGmHyMGb
5BoDlFTnwGJHya7s+jIBa0ZV5GYizbtQ1BhkDfpm5N1wC93BKhB01DgvDsgAViy+
l4GFMARVV/H9m+HHfya20ubtUBEH7cx59l6ryxOafNYq9p+eQkPj657ESdXZ++U3
DHftUBmd9h02hKk0S5B041ciRMkg6r+3I+EAzwzFbhAirpI1YXqehSw7LFz6GfcP
E/XYbIpJt94Z/M53HMNaGxqhhA9pjfvTRrLilxgHrL8Rwh9aMLojKNqGKyeYGlYB
4pSQseG/5xhy4ELD1CiyUhk9Rhc4y9Os4JnJRT8oRy3eaaMd1fE7KTVKm03k/xwS
yR19aXiBd3UUvPgi4ndtYj+Ls8uzkJ4jS55eeJmw+9vfXqap0wjgZ2pWQa3OMNUK
kup3vNfUvo9ZYuA7reiGC1DIbL5s0hm2y+qqg7clh2NzlVBPC0Ppa7XASh80RgUQ
yG/oUu2fP6LGgFreUcjGZiFGytxKgTbxpSqhsS5aHJyXg2Zqr34qKtBf4jgVNcHd
febG1kpuNHKSecURpd/J73LHrSwqnFQkq5xIfTdRUuHidmkZiPh3Xc1XD6pIWvq7
wPfY0AH3IBZ429GpZ2zYZbBOqVx3kH+RaxRjklB9daztPyP+e2f4FTPgWq9pNjdD
MwbqbgVgzMQ3QHp8rRti+f/XHmfLHkH1tIvaj+GeOymWYKLB+R62Fqd9FNLN/SBn
LTFoNDGI5oWenjPCmW/5GfmgOg0PF24iVX3s6lew6rQHNh4JE8JGTL2gpbaaY4+1
7T++Jr2eM3FmtV8CYlNPLeqWhxopWgWReJ4rCerGZh4yPF+RLo5tjiMO9SebH4bv
IB7d4gSKDPPu+aUzPZwUl5ENVilC8LganOwS/vVu42GzZpSU5etx9h7nQh9GJTl6
Qb6EFvuYtyt8INGmh8+/YoiTHsIJHFWsPGefMF7Q/0nckvWH2scIu54U4O8p9dGg
xOzNNm81+pDlNGwacTU/VDkbpJvhtZ5BhpaKJoumQY+LOhIRpewDenXTAWn/Zft/
NqvWjfch3y4h6qge+BiduBj6LHVzrah5f/IFk4qt1JsgPKpl0kKsiR/AxSOcjg4l
TId8QszeiwOipCfSOi5faoDuAnhpfSmbmeBoH9ri5EwhgvXIW9gWanW3QDkhF7mH
8IeAC8ZHRusSsmyg8gQDFdfhgtiVyVQuPwdyTh2Dvub7FOGW3QLmhkxZiwC097H7
zgTwdgKVAXW1+kDInisiXp+8E5+BYuo1t7MHj5TNIN0uvNmgatl5y4w+R4w8wMA6
bmukCszUSm6Z8QeUOp5W4kqrXc6iXNcliiqycpi2p1/oMGSeVB0dILSfJSxTbhj+
cIxigsMCplS6B9Yp0zXhAtd+gAad9+ysE0s55lpQ14UvUDdoGJ/E0RxgmED434Fq
KL6/ULJ89YXQ9mye5BA++mIoaVEPiz9nfFCNy/bSLCnQavHGS0fiNHrob3Fs6oJn
q+9/lrULPuvSkCjQ19NIOJmI/NVIlB5mePoEHY+Kt5Sq0KpKs+OWHUKx+9sTBJZS
fHnhcOXJ4KeH7EdBJrePK+YxVM6xX2pzPS/dv4h4ZzpARSm74iq2au+qYYePsP73
o2KKikdM5/Ajtti3Kma/7+z48T5kDqT2ZogAbxDnF1e4glq26ziY84PPdxM4Xt1l
ia3NZO/1tNLCUdeMJWwEI8vzNMmQLIFhz4Hj2F+Db+24uN2ARlDSP3ztobTR/PRg
mf1g/CFtnU6aj1oT3qwcQE2P8Y174RKA0urbKpQfW9AQDIAPN/pGTg7wzw3Xv/D/
CGiHD5+/L0Q9W38MYsVHF/FHBHmjWDYugvrPlVrK+BHqdG1+aF7tFrsEYKiYdUWq
2baHk1Ten5vLglfksL813rrJdf3ej7wt/yNAsylSQRPBScrhya/TvfupLpjjO8Eg
6HPwrIa4uHH0s+xNrgFqfHPD/QOzaL7zpME4zEzyGaJTsmeaOxUusTibXA6umNr5
A5kWznOzqUYNNx57Zv+XBFnF7En/1YN+4u+czwNfSUFUHTZDsq6XKBfaeRMzS4vk
ToTzG0dfRl1eze76Bgn+6/af6/f81UNaYsryzPrbQhef0i0w9PP3rqI1RRXrNj33
EgPnCzU9uVC8nisqGbsgm7irI02+79REguUM3Ive4P+4fP/axPLcRqbNYgtG4KBn
cJkpp+j1Nj03ultsvBY97mQXfukb+iyjubHJuknOyN4grH/682vOPV+FvPPizWqv
21DwVt9S0jyyOo4XNFT1ES7qZwIaGH7xzjYSyLyNH9lN/CMEArOhedwk2kF4FiYT
F72QLn7wn29U8+Zn2tXoeZ+zrEmMw86ACD20q9jrXzZutgKWKHTTxJv4gCNHXee9
a0w5gLFIOTNbw8zQdY/YdKbRMDBJ87TQfScMbXcXffHI9wmda+om5UlHhfdse9eP
12cdajqu68ePnUEpuobpjjyhGOrhLtlzmyhzKAOHr9aInNvH0IWjfNyf13KhivHf
MxkjVzJNGC7iVd7/1haspWpJAuD374bsIhunkV+yopExNbIGjNYHFdO18WrmBA53
Yozro7k5lbkL1R88JVAEknFqhUZwnWMCVN+JV/DfQNI=
`pragma protect end_protected
