// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:39:05 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
lBEKl8d6gnOVz+6CBrhkoo1+vr9jS9txh1Romiviyueh4M51vt3NWNCukZoqSOJa
Af4yAJQK8u/iVEUwihdSUxz5++Rfn0Vwo4DNZDH4I1dlHwAAupeeEHGWUfpZsJCC
CS/aAiKhWOLTOkM2LZkU3/EJKfRJJFNKuGVxrtxBJJE=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 24640)
QiIz0L5xWuCJMArsSLLR1k2yaZ70rHoSNaLtt7+drrrKlhJxW3aqRJYoIv7ODXZR
YHrHn7Dr/cvzjl3ntwtxN0sctzOMBvgJRfNfhBLt9G3KGj94jVqdIQhrMOYK3inc
boB6zXTxRnRbHlT48NDx7kGeu5vkGeRVo0W/1SKy2HSpvPOzm1+QW6Jtuyh19viY
ZinCfL85wL0bHQGFCLdjLiXT+zhOPN8+6ybIa51c4m1d98Z6qta531JblSLTlWxH
+o63+GUUQJGBZ3GhYbOQHaYZRg9jrzC2oIQ8I2TyT8BGmuXgDDtbfAjW5aO2utQa
2YwtM4l0wSiRV1YPmj8GqeoKBNTrWtvLW8lI8AhnBwpSNfa+BrNFIFSw1oNlftkO
hBhjyHIlwIKlFRwRplfMi407EPvtlJwn+2+s/M9QVbnF4ygccom2dAJwLEzefKTK
UoWBLm8j28wDKwrhYZYIgE39jsAMfeJaOT15B6jCuNBsPOiUJc7wQ31Dy96dWC1N
imb2cMUCxj0isgl2cjOdrPEtigpnEEQJWUC7TKT/I6lqw8jyIa4Or9PMmY7voRVK
EkZQ2r70mmZ/BY2G+NnU8XHgI4R2wlHqpiAKVd2UnrBTfir52jARwWme02gB0ocZ
grCv4h4IOW6IPDBw0vuNk5b/ordyyq2Aurcn2QGZkfoohB1Olp5Qr5bayhImuIsC
McMb/eoh+vmeVK55XHKfnVkvQJJsX7/L1u7mqOJN7N+63JT9z6rYFpj4XisYczXi
Jk8AhV2zVHltZasKW9T+gPiaNfYuzVQXo+xnwPZDMsk0Fh45RAwJFrR9TdTvZ13C
PASmNxQth6ms/gc9ssiUQro67ZdXeruknwjSDi0UBCrJUBq3aUNq9PllFnMH8/WH
yiukM8JBfulya16cJkPZSk+D2ZKFaqKQwWA8wEfdYWGkAi5x417YpdeeWX74wFj4
M4xDmqZLevAmawjknhojePjNSy1SkAne4L41VXTqPruSsi5Ywfj6OHUgnJYJ74jN
wrrrpqA0lEBFAO64bxRIxQkwtmDDNc7BGGTE7tMpDhUuzFXnwTAdHJyErFjHDxkH
vgtTQ/b86CYcHCzUchaJ4ymWj9FJ/9b6/5igo03Zi7Jo7guf6yb5+haseucv9Z+J
PIIBD7gOPZM1GHqzUp8ltnZNccOpbwNoyTl1QX3DgKs8bwqevOP343odBE77qhwD
+xCBDxgilNAHFUiCNBU6G1n/I6YkUhGeB3jvpNA4RzNsVdHJbI0XpBVfvqBDxZSh
CjPIghrnLwdz5asmJpTUzQL8cMGXkvEnsICRzcjzlOPft2qrX7kLdGcsysRRCVCu
XWFHcmDQRdrGZXqVTsSDM/t0BBgwMe2C+GdkPVSMdfJFy+84l+MaRia0StrOJQp4
87jPsX7Hd3k0ji2NHLEbvzXLIByZWeFqkFXE1lrYoKVuShDUM+O1pMgnW7QURgB8
IHig44qt/j8Qv/FRUjnbBXnaVNK/n77jJTgahrlA1IDPNNdI5olX+J/9IL+udZcZ
OxESxJGLSZa2Ds/p0wa2ooog/CKaxYZFMdKBrkAW+P5tsnYRde0ePUCnOeVe2Tep
J0Fb8ItJ/hCRC3KVcM5V7qA3ereDA+Vsj/OJ0Ou9v2kUy1zn2fDSr5RqoCSsoPK5
r0OLikTOA6G0NeI006G2L19Ysabq2pou8VZziOoXu8hX0VkMNGAJ2aa9Kl2qWJm7
djgJmYKoPDMGvaQDiqpb4KRTc2WWF+rCTdEpmkNtAzxw2rlCsLO8rvKssPVSKwNC
al3y9ymR3in5eWRzfkV4U0T2GWIU7MxFz0/EUurfKj0N92cpumqmuJvI27Duh+o/
RBJCNFBED/FXzGS0zgA31aStEpDaB1riVpg2RlRGg84hqdtwL9gT4X2vfdgk211b
St5SdoDcGqLJe3tNxRsXjMNHSmUmrOIUguxBOJ0BXyZXZIRJHGZcS1NxWGdo2PP1
wXkPqDoCfRlf40P4avTamELp3XoCg/l8VVXRvw+/p3GaiXNXoJK4Yd9qDHp7Ccy9
6E6WZTqCeBesrEzxzIaOahGJnTUmRUfyQL6nwd8SPgggZncE5OKsnJR/bFa8fcgK
sJIV3H0T7QKH5nbk9jDVTPuL8LhcKinFhCDSTzZGYg7G+0G9QCoDvY4AolGc2tt1
S8nhlFiGrfgKhFf1UPBD2jlIuvlI5jnEgd9MMXEb3waGyX23Z3+km+gfFM1Mm1AY
HnjwwYRlShHfn0zy6HDdh/JE/kO3LqUwKySWJaFqkW6HiYgqhkbAvHwH1D3Gl83u
kHjYKlb9ep2tJ+fe34ps93qAFy34RkNjVTKJ9nwaAvLFzH2ZLqeI/6mJtKcOergZ
AMSPKiFusosi6EMCiEEJW2dwbLM+VQ3R+AESIiLQm7VB1qUNNq44xijvP4Qln6z5
vTO10Wv8+FsNrRlcim9D9A+s7hTCr+kSjyftByf6P7J76NYNQdYDLW158UsTM7NR
jd7L90Hd31kfrTTVZQ2bkXhAnv6QcdZckzIFSWj49yWXnGoXNG/HMLHouGGGRajB
HqjdORi2bjX9IrPCdthk84jBh2482h/qdr0gFz2Iyl/crcydKgViUCs1U9bOkTks
CI9bfmsDnux4eCdj1JTsMVdmJO73YKVW2GHl4LdLSawbeVRjhXDUJAFg8XsBRfn/
dp+3JHznoJwWDDxvPn2II3+vLvnSE06pkFTUOsZTRl86hf0PBm9t1YHDOlXXR2Qn
5PrmAKZzu5W7kKVw8riozxUvINoKFY0h2t91GVB7iSpJGVnQgrlgvF4uylD7piYG
7M+6Ekr4Gmyr5ZgihyjqvvAdzEKeaPDe5Zbg8y4ye6m6FRQplMwFrQxiAFjNqfcg
4BdDjv1DMD/ZNfEue3OpkzY5jaLwGK3dj9pI+orpwKkEr4x2GRax4Y7m+j3J7M/r
1GlcMYiq+UT0I4sJLgs6E7/m3YrvHEenfuwyIOLo6kfs5Mf3FhW7DriReB14ofco
yvuysKezjS7xCqLyar4FdNfYjLA2pFcClO9HIZ2fmeEb62AgDy2tzFBygGDpjRjs
gfjR07ds5hMHtBPgYju5sTBxbAtNAfkcL3IcnFKbx6xRt9Y5e/vUb6SBUq1nVSYW
zGFzQPXLuJxzTwSBgsDebH0NF6FZY2CU/k7aFuft1rxBqTfeoTHZFmd0323oLNm7
dU2j5q9puU1JS8MMJ0dtnsgWvtxwcvWIUatJtwu7meTv/MEPvE4Xc/T8C+4O2Gao
CAPwVcUKa7SL649ydDpgLLtD3H1Y1draPuwk11F8vBCZWN9PeZD7xYt96waHZs/U
ePt+EwqXMKziiq/cHHPdjy2f/iwaa6Rocl5esaQR+G8PYMfLplKl/FpRubad2fTd
7lLAr51bfcs/rlfFmD8iCqKnV/EOGgjM/3Q8Cpp/uWUD0+7EG7cCgxldrbKN2/Hr
2HNbznpy/f/9vSDgQZ2pI9tWelleuB3pqq+I5oWrv7CAtl4q/Pc+G8bswesqL1Gr
RR1kMUrNeb2CciZmDUCyhkEKnHIktjOS1NQZgQlM7jiaEc6ZSobfmlSroiWqIgRN
MwLCu3AigAgD7NAim7QAw1lnAVV1D7IWsZasVhzl9YfPTJJIT/6NvsHfLcMADgKP
nRkFVSKNhbJrVnGH+obLMgNSV1SZv32A4IGUKjGJHLMyHEPlY3BjYAh0YoVBgcDG
c6o/7aWPZ0lya+2qimg3Q58Bj1wtK2PiT1dIuDnwHZZpEqaE2tYsR0TCi6kc9X9x
ZvnduROGEQcGkZo4Zzl4zmNwPojzNVlhHcOXgqPEAkQdQ+FvNcrdNXY6gudInWA4
9dzh/fi0dYrPUIciXBz+qWY72INK4jRNLs8iw3P5x3Ft7nUkkcn1lGtydYuiEtvD
aj5F3GF3CA+Zxoblp+LS5OYuHgKZHgXa+vCupAHkNUsrcjVpbVU8zRRxZYcdLSPs
N16LgsPk0CVHthgAgQhd4sCymSkz/9I/Iz5uIV39BwTHSooHQ9n+oJlkjAXIKteW
/JaMyBQaZyhK4eVHuD7BM68E/NuapFLZka5cSqN2tFf5SWr7cOIk2DJjBfeD1+QZ
9+6aA+rKBIdm/r06+gx3hV0iMhamVirToVj+IN6Q628f71F5Vf3z0InbGnQkCzP7
SXaJ0G6pOx90I9MHfgKsoLDalzUzwG6QG1NUhSLD11tR0Q/LETdvg5mPvNCKQMtu
tqmfXl6ojIyi/dedegrQewYDEh3SZNJq5WhJQ3vafF+AakNcIXfGe1gr1HPX7zZE
I1OKIrB6WbDiSR9IRMccgdW3yqpzcpbu/qnP07DxU9oHMZ7k3KRt8x1wryOx4mvE
aJzLI4WRPi+EBbwUr3HXuL5lJW4hKXR61kgV2APf7qjNtf71OAVQCdYlSSb0LC/+
OzOWIE4BzM9P1osDdRS/9xPTpcbpXYCa46MRD0WyLivc3gmRwsuH4ZKuwgELzSQO
gUSq8P7uO1zs7k0ov9AgjwgMza26UkBHkZK/GXI3RqaIvM9Z4iQhcjP+W9kCYHp/
RfM8OUz7F/KOpqK63q8pKcLF2jI72ZXg+gg9dQTNsbDJaXrcd5l2DPUlC9O7o7NN
PGZ3nEsvVPvyfNnNFmQlMJy0fengm5ivOJ0HoIrI571Lmsyht/63wAajl4jL31JU
heH9qF2W9Su0cGalurmjgvi1RkMwUg8yrlAW1P7N5X6WlO0l9wqzEkvTQMoj+9jZ
kzTtMpH0aHcvMGNjJ5Lxm17o8mo/HZ2LBUYHHGNCfbPGDT+9LgBhv62jSheAhk1U
fgeEG9AKEod1WCzjTorlDtpfYjoXvmXWuMyJGbmM7Uyha3PlF1pbuKUxcxiQOl8n
fE0qhJzGhAchUOHvi2ffVW5K/DqBHTvBCfDz2I7kFwzklvzFF2fZ4AAGCIZ7lfk8
0Ga8/4DAkNvzI8VXR8wTIlEd5e5y/UWPuBCbbGpi2eMZ7I3ut0yng37ODFANrLSp
5+qzUTUfGeIGMjz4CuU1HdiR9w+4g70P/w5U3ctpHNPe0/uXT05ypa8+NTphroTV
Amrst2IJfb+nAtxZqr1QZjYK+v3+hCDL3gduYxp8gG1rGlHdbxdwUruu0kAfoVyx
VAUAzemuDTvf77YtoKC4Kbz34NXomAh1xbjmVVyi/xpoEMnZHi39j2U01mZb0/2U
bP2AM49XWZM/7xwZVTlLY8ri7td9nv4Rzl93ghXIIJ9WxZohHTx7zDQ3aB4NcL87
TDW8EHYuDTJNLZxsC4kHSwmWWz857CfzFMXB7XEXH83pPLd7O4Y7uXsIE4jLRODZ
fgsJpFYYGgpK9xnH9C+F5Q6n9eFNwFx4vB0ws1N/m41Nl1yi+FRhabZrzBXYdCRb
PgcFIHZRVSS/Nw530D2wWCzY4jH1st1qCAuOuGybci0sMCKypnahYQJLp/KpI8Hk
cUXqnssTkdsCDyh/dNlJRc9Mp84X5EY9B+aAtBBKCDk+t3A3cA5/P08WJtgogzxA
ZuGHwUWZ1bHz/5Rr0yagYM5lOcpY/fNEv8392IKqLgwwB+baLTN0IydILIG5jUIh
Xk99R9ixeemE0kUungGzzcmnGHdXQZFkntDhz1YF7I4Ay/MrQpVAyBMjQlfoBDNk
TrLHzZv68yHT4ZazS1vwDWGx0eeV+Js3IdOniIW/NrlU/M3gg6cdlXpF6+i12A1A
g2jEdeZ12tZmO6GzCoOPkBB3AfoaaNsv5BVeB997ekK3j7csmr4WeNlGnPxFF7TG
Yp9XoMcv1NPEqggq/Vsw1UKv6vIRdCV+0+ejtX3H7f/7P90Cy0/VWvcBZQeZ9qin
nVu2IFQ6f1ITy4NECI0sqvN5jqlRGJxs2qM6PFFAYZVh9ITZ2kLfhHjIX9zA2YsL
vV3NhiwNvTg8DPFohdQrBxJAvQan86ouJkY42d6ceWYftVwToKxkkK3zMeAl7sHt
tdRJtS5+TwofXKPth48kho2i1QvuTI4U44Rs14QMr6yKDD+JQjb9WesxcXLNUaAT
cd7IoYtR1uJh5PAPL6qkew+mGuGispCcYB0qv+h3Wuyw0murWYGi5OZKkzPwKM3P
z9ebz2FrS18QVMlrbq92+sNpnT88r01HkAfWkQUf+c333vd5adcMFA3ID8Grmf1H
GB6mY3K2AcTyqmq554e9aI+YhfOwfYHeFawdyADsKNgZndY+7fMJjpXL2BdHRitc
UX0/Ei9Gq4ZtH5vRrdYZUIyHwS8JuolwyWnhi69AvvnjS4Gtef8Set8/reafG39O
tGdP0MO2BAQTonF1MWw3Pz9iKenngsG/cMrk9D0GEnC1Qf7wsoi9ru9ZqkUzDZDb
n+jEN06dDRgUmUz07R3dviIVJYlEspTVae10eRo8JG+facYYCnQ/HC8e97hnlz8T
RRmUelooHm3yI6a/rWDrZ1oHQEb/fj9jRnj8TD9d12h2FXM88b/JZDWjmQ9oxuAw
sspjMnSsS4qNcHmN3eAkO2BOMeuEOgvSq9oRgCBwUSWoC2WwRI8p321OCvaaCxQP
ZfgLoW8ham78nOhlGGlUKqHIcjS2o7kHsnLqb4fIBDCpT9x2ReyE+WHPxaIBWc5E
Gn/Iymd0rbthsRkmw7Bkw8OZLYzNCvcnKcNNwtJr41Ux4DxfRFCXk+x2H+Vw2dof
ywwLpB2mAlgajKX5vaDBMO11O9O/EUO97pu02T44a2dQIfjxiFkxsca1kIa7KKGB
HiMdPDDlbGcgzCf6pIxwNin0B62NLIUcJtdDl6V1oUpCrESmk3ww23u1jrMraxmb
zvqkJimXqIBmhJpchxva72dFkzDjMilOLzLuuXNOnzqm+YfEsWzDk7LBK47dHLou
JiPyRNMmNkNbW0/QPh1HZr3YN1GABpZyEBHdeKWoJDpelZ7cRNHMC5XDly8Vjj2D
v2D3OQ34q7TRrWmweVktmhtqmrlX+RYWdRIeYsEYybb0IgDPu6bGxvTXuoWp7UiB
hhPdPh24vWzv6NmlmmBlBD6z0x75ePx+w0nB9IzHLhXDkQ27Nw4OtdUlgde02Xkf
TpvLjn1KOMoYOI4XS2Bxuweagn2Eu/iRK4CIrFOl7QHdb/tkfWCZ0K0z/GyhOWTT
UcodH+gkwy4mK/0uwiXFbOFfaWzCRmNht393EEeFo9ZR8NyxfkiFcZER71k80CB4
5Ou8cWYmb8738FrmvARxJ/bvciiFTz1fQIHMkM5YisBEKT7OIInCnXTP2uzrUQMm
KG4tmaAWEQS+CUClSBt6UH0C68Ueu3bpxDLZzDdhsftEWZ8QhhA/OkhM5XH1a2al
g6eSngM3qiZ0hP6CCSIb0kMECbevLFH/GQLRV6pwYpqZlKzQjRVQMhzLU55rrnFw
ucoLh9sbBbn8iExr5czUnMYy4pFC6IKMvHxBoSEe2IaTI7U/B4zV1LpaIH4NgIzi
vdsTv5JB4oECudqhEkn8cHPwL6kuJA/qE82LSAS5LbS38ToEsPj70nhmXu4XYxeb
ZbT1d4Ustz1u7/58gZK/tPVGu8ZeJSZmIoeUMrizPMLN/43UG6JZYyM09oSWHsQ0
dSwG3Kzu1bF6blvctXiOHH79HK362WHepLhn4hEnFmkEG+ZrNclTAEdgoatfxM4S
raJLwkF8fWq9AV2N+UOvKA3qB6Z2IiimIun3rI0JrKLqzz4Y1MTVa+9NztycuLog
B8iLKzA64f+hWykXkhhD17PdhdbHhuudTCqSd2I/zewgUZHkLXY9TLADyeiPEdIa
ucGrQKq+WP+RqkdN2ynnR/LrCoxB+CKQvZfMjZBzI60YAQF5JCbZwrr68VZj+/V4
S0Fv2i2yB4elBgZue97xa/OUu7l59SEbbbk5a73sYwgVcmxwVkhIvMZVq+Y6SKb2
se+++/Vp8hBwp7dFa6gVdUf7/M5fvetVIwutk6yIU+h8PloR2sDyF3EIpIpAMnOg
8Vl5EbL4m4TDsEdoFaZ+PTdQ++eQ6E2oEOyNJal1NCoZPCRkNDJ6CJvEoExEG1XF
5NE5RwTQ4qcOYKijKXjtcof+RHc6t6jRyo2jeGvMs4FJcaQcjaCm3vkwz1O8J5Cq
5os3ivefd2SUsU0LTl7lHKIXkMWnRDy++Gqo2GqQorKQRX5p5MsToTM+98RjwTrB
uufDCxA9o0sqppRx3ieirX6Sh1zUnnfHJNWNgR8gr7pp4aF5BEzatTGuxeqX33Db
zjKeKWiKb2Pw1WnKe2G9t/XOPr1IsWcvolZjdX4T/ZA6jfmY+t7QYj5Srp+Q2IeS
GTLlGfY2U+iedObOAKDXYL8gVpjVXeLw5WIJ2J58ftzsTCPUdYnVlvINYwYQVJ/N
t5h5pXdZtqv9onMfvgrwu9zC4YNLg2gTTATGJUG/2Va3RqiyaRrqvn10Nrwq8pi/
Oi67VzpnZ47o9JIhgqBhs/STLOhTWe9PbFinAjDWX9nABOVqGJMxNirZdcB6OPkX
5CDlKz4O+byesvoXw0MlUSVkwD37X+Ada2UE8kmJertetgPO0wQz7uY3BuI+rbdX
Irdlog5pIiy0EekGJfDPN/F1Lay8KbuEhI4CXu74mr7NPFhIaVEK0CIpiiFYkUmS
euuOLzXJWo2jrG7eksXSVQohPma1k86N3kT2LMe5wOuhNBHNm2ZE8wrU3CZAI5Er
0n2svLTUt5ovI0P40WpgvVehaccdsk9zq3NrkydG5q+i+5xk5jVrgVa9OdRKEtSe
RYE2bCiJGuGzVIdnhw9/yHaqdNPnPgq8UP2EA+/Oe2vNaMNnVuu80ShJkPSyq3ln
w+hXIK6vidkaQ0PAPKIAOnTrfTCoph2L/qB3L6bjTuswXe5D6f7o/5uF15MHbSjH
grlCx3N2SVZjfBHTDljP3xXxnSpqOWQ4O+AI45UESn4/Jh3hM4gq3DXRawMEXLTn
uv85caHxhTgOIvQWovsTwMSBZFG98BSDUPTqp3okPDUQT8YbRkZey/cLvDSt5xef
1eAdQmItZkddY2eMW03ri1IVGW1r4/AzBWTNqzE7zgPFaNG+VFW5tr2V++ySY1YA
2Sul51iJ6Eb0Q5EgaJIFCZfIpvtakkVVcc616QlBCOoUO4jWH7QLDISrjOLN2jXf
iJfS3xT9AQM64/QMoCqeS9UpeoMQ0/bWZ0HhahOLgqqHRDKwE85zvulF/hxvF9wO
xh3Xhcv+rErixfW/ZpAJI7cQJi+VxjO0m/lf4IqolNTyn/BIbQYnejrbYjSyiHTZ
jlRLjTJW00vgNnCbMScLk9SB2qduoCx9kwI2r7T2iQsoXg7z4Os4jMI+3q8fTBi1
lxU3bFOwJeYgdb8iCw01aDMJF+65hh9q0gS7PHOXxQOHg5tKXpnhXlmgSW8xTsHo
K/k1s9p+aROqH7AyqEMUXQw5Go4QXLVQuJ/OjPRS/KB6uOXy2PVu+lzwa296gJTf
4eXkTyRA38kKs+E8/xQSDSZ/EJOWDD48PBbomRGifvx1AsJHh/abWWVs2SSyvCK2
nZus6NDTAEnZQTqvOA9L8uqHkLS5Ewj3yu1gcTsD4Al+dfDKZVBGLgvqJXZB+bZr
+meiW8AP4Pkr6f3Hhili0ofdum8RWn5/R6AQXNezpxS0WARtxNX/jOUuJUCttrAA
dCa0he0htXqL4tGEdnoMlyYC6xFqhLvw3WVQjQDyF9gjTLB/pMmmJTDUBKJN5hDr
LOVI3UOWdl9wfcQT6VepY1iFFh0+hyu49CqRf4NPz3/M8iaaNyKDAiBPpZ2hoGRm
cebOZcCjD3DV3ErAX95Z+MLa9wqgE/FTDJEgk7SLqZ3kdQGsRdE4UQWqNBDHIgNW
crGIIIuvcPIauJqp5a36zDBTPAS9emNfDNwVjTU+qzC+rEH+FwPW/KMgl/cJYiwp
Xw061HxHs7/QeLW6ntU/c0KLYKimCsiTIUIk0vMoH9LkpBzCsIk9Td+lNfpBcpl9
888bEcVA7sg3qma8vRWt8nUKVWhVOmnvZbTAPd0Nu82nvC9CDv5s7+Y9M5CPg1h/
2DDd9+6dwNaWSNrTYh8doq86Kz/X2NE/aFXFs8lHXFFGnhny09AAVunU4p2NB0zQ
69n6b+OuyUWfQUh+PO6FhRd5ouXJbXsnjnju7PmbRTcaGWTjx8m47lpwd+vZ5w/V
ttykym7VVavLDq1Lh5L495ZcBGLbosVe4Mh8mEnoXHQp5lUcRarfxTSwcHKUdTga
0weQPvaLx/vE0lOaDowWPLyXDWO4eMO+2Cfdi7q+SK6ZgTBheK/6lFHX0wAozkjK
MECqGAOMFmgAyeAQjWEs4Epc6w93b6OtgXFF/p5Lc5QDSi3rvvyNs9MaIZZB68zr
MF5qSvnJMSrMv2nd+03rU8BGvnAliUA/zs5KWD1DhQh4KDWygWGdjDMO9GmQBBYB
D3+pj3u95L9yoVOW6ZSfGMpNO99Pc7SfAr29q/vtg2QKb1yPTnuZU/fjpmLiacys
vlYXBlI7EqvZnvw1ZrUq9sSmtjh1vNc9tk/x+2LTGAjjI2lcGOdTlzgskSXEjdt3
GBphRv9ZI0ijYkb+h6qMezmfE6UUs2QZOC5zGwPJhi2Ds0KMvOMrixyCr6YOBAKJ
iubyov13uBPB5VA7iC6dDbJWQpD0u1blOqmwCxtAJo3biYmYKQPFV+qLvyiTAwCp
iDgdsSU7xsVjVatd95zJtWS3sOW62HshIAn9f2v53TUfPiY1nDwbClHEVti5gFXN
DNQ1heqUsTK+OcC6u2ZqkI80BMCVZtL9vKFrPAiozSAsuy0jUR3PbhEzJq0NSed+
BIPsPUKuCJvuE2Vb8t9XFEYe5pCwAjeH9+FFjGcFpxQE0swvuspmZPbiKJWAADFg
FQbPc7qANmCuaQU+DMFRC/AHidDGpAiEZ8u0ktYPThALiRIM1GLN7WgiE06gIHmF
1e+U9pwJ4BlnZ3OCbzBqb6PDqcHjnIttpwN9tZ7iaOaR4biMZNToY+Yxg66F5k46
XLRUkhixpbiWHYLuCPjkNBzr3L0uA/ciEck1cx4x4orLNujRhUw8NMoveC/EKfIJ
XyJMuyD3yw5W5k62i7fToLwQObDWgoEQg0HUVew8T9mnTpOIBd8pCd0x9T2RAf9P
8sN/nQJgE+aiDS45/CoAchdXSUfI8AVbQuHvBb8oUyIe8T1s5zq5D05Q4c0pA7NB
3i3yBRWMvilhc/JLo9i30nEHeAf38HaOaYkusKKuuNYC2rxi1cvySXhyId+LcjvR
Mf+o7Bubw1j3g8jiOuDUXFcTv4V3uQM3hWX+v1UICc7lljaQ1OZCifSlh/OqoPkL
ZVOruFwFWb9o1Rpf9vi74Y6blYY0bakmKoQ70Pgo9NCefUgIHE+muicfFjwZGhtj
RLFhUstsUNKWIsuwkWTuNZMejR+BOdhkiCV5MfUB5NzTzHhzRUSV1nD+qY77pxL9
ToAjFHD2tZl+ZDVEizcziu/nNbXnCLCYPf5/LdXm7p7ve2HcNEVR6ioutcNUGYxf
j5bFsH4BaL+7aMJ0D88+WnCtoOl/Uz2/D/CthvewbqWcjMisAhwwqpy9tcMOxWLE
VHWa6bbBJxSsyTEaRZxBuBosWY3usFqHmVriB8lgj6qx/H1qg06TKCt0vKPe1S48
qCjOeJX9zRPN8jLYplAYwLiIEbbdFqxg5CEjYqbjcg8GXQ2cmqnUlCny/OY83G/5
yIAWEDW7OCqGQ4mTNfbgSJeeTEQ1hugtcKkGM+hvbmwOfCV1gU8Ig7s21FXLrFGE
UF+VlflpQ22GWSwzN+Oq5uj/sp+SY/QrlcHL2Xw4F7mHRfQMWSlO52l9P+nzaJ/R
X4TZV3TYmpDHnFAdDyZYefppSD+0dAe1tpzpeTjIeqWwC1z0pGLNL+6/bVkO2UCL
zX/NJ2+2qEZn6xo83kkg5BNaRRm9Lv7H0u1n4s656hSHOABgDRFx49v/tnBwCQr2
DoPpPbBQYTYm4WuqUBtEOvSEQz1tX3awnV20uLiPER70/rOqR/2kAX72VLTtLtgs
xNhN60o+07hG/KViU93KhMnB22XG/u5JuMhHrYUFBKZJ6qdpr9CBFuNOtJrIONkv
k66bprLMC51mZ0B6bEbbQXJI9SvQHPYNIU044t+HMY2Q+7h1xWgq8RacOaUQVonq
TrBr5/KQ17cB8CKFhjb+4qt7MJWI2QJ6SEPteKdARyS5Djx4o8DA6j5PwCKSds/x
M22XVAvhX5axRKvC/ayO7pK4sW5B7Kh98gXv0tPXVScw4gYFeyzH7h+iaZ67Z/yp
UPkWJ/3ADKln59J8T4j2C6tWivcAte/PaXQ8kCjc+LgsIfrCABtIdu6w0Z7PcH6E
ev3JVaq7Clc1zccpaXWgmkkQbdheTk7baGh8f8C4/aJmA5Ff9AGThacAtBEM4Vey
+Dl8dsKvLhQga/BQyKDasm1Zjo5YSz4YOciEFBv58ybrkCIVLbZTLocKFzF/tJAB
kY3RU5j7/XCngtEF6dp9byYNfQBT85bUm8qPUx4Urlbhn7xX6/OZEImXE0M2gqpa
1b5lJkJA4grC5pqOsbiMhlYwrEJrvMrw4LMa2wYlx4a4DZqSczdkOjZPis0245rE
hQyGI5EGQiIE+FhpP4xxnnMZ/VN8QCf7D15C5z+hcVAV6HIn+XBs/n13hWgCKTT8
kn1x+ALi0uLI6agpUFq7zXLCRq5jABjSA3v0uPOspd7MYi+ZUw1KlGc6PSusNtSh
5p20iSdARr7dsUGk9x69edBGxAkvqJ6++oUEqJbqtH8uxokreMHfB4NfHNST1bRo
KRa2pSXfPH6lO8gF4uhowvd+gY3Zl7ATb3Jxth7Yi6V7k/v0oWbV9+MYTCAsN0YZ
W/AU/nkTxmNRxmlGEEbJAHFzPCKyKJ+KPfNB4dq7+F0iTsaWuF4OyCgr9l4cpI9j
wdrR7oRVsySvjCFFVImCSNSd+XS4fe55l6LUFu4Nd53muZoeVFYpYq2izvf2WMqu
bzSM1+xCgDQQTetM3XajxUzOryu/HCWar13VDIW9YVy6SeOF/q8ZGiChu3WFgBzl
esoPr2+dPh8iGYH+9zDN9KJ7vViM2gSwiQ+TPoTrHamcts9904VocreiVhzZ/3B/
93WQkMJwiFgvhGeqczu2hrbex23mEWLkahBas0sGy/KpP67nAUD8OUKGwfVn3MUG
moNjHz7KecXH0RKHIHTOFD+J+9I+nb7xh5PBO9o9baCAMir+SYpS6KW1743v/GIc
dTXqD4iTuFywdRbrJKgJkDlPBJiOhgOum5LCGF3qaGswYAmt+I0TS2fG3HFU87tJ
BnMW0VkRzQvxx/nAVaAsMKzI7DsKvCuMq3SU/r37ExAvGiUOi3wD2snN5oFQp5De
3J4q/L6OgT9J/Q1TBUjfw5N34A2fZrek+PjMA5d5KPNXEYCD4tUnzDxat25cI3zK
6fK6qlDx0luX3yYS3KckbUid5MsGakaN/Si1wrtWNxPsC5FtuC6gtVrQoSrZcvYr
uuVAGryQ9EMyt0NDo5uRYNIm3Dx2eTX2PdP0wm872VdCMZWWkrbV3+OhH/ZkP3cA
2PKUHqW/jpaMn7zKGeyRXn8hG1FWmS35/V2g04xaj/poZCo+DYEnH4P6ERmhvLMC
sx2GygLWG8gy+wmWKD9WkFkczOnQ227OinP4yOrQ/osSVzgn36+XgcK49fIRnfOV
8FcBapJWmzEwh7Af1yQmw3HyVuZerwOWr4GEsBbIZP51dDn2hNAQkKxWVqqEx53x
VBj26s9xXuyA/kWMQG1LhmVthPoFqL1nlfzDx/hfeSNl/SuVZdRPDpXphORRLUjx
0nFIiNe6wj9+5/YGJ4J69ycqp0yXf+Y9FRsrVZA5pIR+UCoj6ttRUrzmtfWHIZxe
nyHlGFzsU+lwD9Dh04sjlhAAFDHhBJ6vR2JHtfPyVw2qgogk/tjZpQHLp2ydIkXU
7WWdEFvZtqMpCRxKDWvfU/CYdCucWCsbmuLddgg34wOo8c8a0bVVh6z1n5QsIC+L
3Ix95YKTWcbYO2BUvrFF5DoRs/f0RFSC/acBO1HwIiv3H1aiL6a1y7VE2ADVPtJB
mvc67aoEryA+XPWGR7dx+xvxUmSvSn77RM1b236W91DeQMLyGY7JvpBo/SV2ehln
z3Lcq1UE2fHE09R4hJfRxQIP9t97FO2lZru7RP8YyhYIAdrm7nD4nhLNNPiqnf6m
UtITNYfj4da2jBn6s0KZXlQSOGTbkp3x2lrkW50JiB7huDZn+RgAswGxhXL7n82d
8fSkOnNu6Pb2qE6jEImsTu1OV9sYRZuODh1VW1bexouejXcrD1sbwNyMpqV14uaw
U9dI7VTqLLryMtQaD7U2qNA10nk0qRN5P2C3ZxGmsRWE0ERjt6b32MaGYncF8H2m
hIldktj4lu9SWbIFYWFn2+o6ssY7Ic7DAIiPWddEqtj8n/1Bx3k6AIMpnMbdV85Z
1rkdzXxV2HDzz3YVC4aoAJZXoEVBV/3qnizKNTaBns8ERVKI5iSdHgAQq9N7i5m4
wT5iisW1wmZbrzTssfaWEqVqISJpt16iiKGTgt2SmNL7HWHAoWQPloDb6zFKhUB4
2OxC0JNnbADp28GCnn4jLHu0pNhslZvUySk2EQ6DjeqXT8FgmPe/gB6Q/bfsHovY
LryJnXIHd6Y74u7ZUvkf0KVINo8j+McKA18PLHcSMeoz5JtV3scAghXJ1CMTylZa
QC3eu4Kk2bYbOjJAk5jU7FNYucIH37WbFevZe0EMnC9mICfSSeAUm8ALV+BfLWcL
WuKGjKsy9SNT7Y86pC+G2kB+e7JTF7/sbSmue0fXqoKtDV2leF8BaJ1WdIIKtzMK
f3Y+WI9FF8aCX09blO95MV+qvWV4+aS7qqjA+NnI+f0IxsXl5k5AofsqcC1nEsDt
Bm9igPYTHp5siq5TGvlxwPZGd+aMXFjnjgqj9XrS9pUTA1HCmjG3NN/nvARffByA
eRmspSBYyXG1P+9UdMEUe2sPl74AZobKXV2Xgt06dJrXdzekypsgRUBL4lXiuSQB
g4B0lj5Tqj/SKzyPzkOfKBeEgoVD0od2xdTEpyiEBdb3k0I+TE7baGnHSVfmcMdP
/Ej5/u6c0X+vjNQaWJyO5d2TpAPXUukflMw65F9zt9TbMJR6TlxNhnSwOhJo/lJc
vl+SEKD1c6/6EiUeGP8cCKmqcJSlIOZOP23OrWDxf/a+0mG8cBJeO/AFedJxyNGW
XP4DJXotqjEa2rzo1LFETpcdtpS62c5QpQ8Z5/dd3HICbdS8nJtpQW/qNESHE2kr
ZBOsmZbkZPguSKfyLB4+A1/LLy5Stor+BU5Xxvd1+bWpffiTlSUGEhMIHGF2fWS/
TZ4ncZ70jm1v41AkANJHoU44V1J+yiYV8ATfbk+TNzticOewciawX1ZaMhQc+ILN
awtklbuMq2viNV1Hq+Zvq2enyDVzsSIvqgQNB3uH8FBj3tUEje6TIAfAQuoHa0jX
W8xCSgzurtzBx+txQ8lc2QUIJtfmmJ0gKEzq2aks7d+W+Ni2rKUL40S8uOZOm7xv
5n5bJqaQLBK5iE3ooyTOB3l8ib+aM9kk2jZzcbhy4qgHgRm/NUykQXkVEECP7u8u
yQDxZ7TSng0qDjcK072LSj4/AOF9XQuLZAGz+z523IVu5PRt7xPORrxQPG6YBArs
F3fdGR2tN29XqC4nNSi0xg8vOsTrbpZXARQKMni0ycs7V+VSThiYjboLvI0FBXBx
hTQ29t6gB9rxJ+FDhG30Rz9ahmYIYRExRj7PC0V3XXeiIdTOccvtq1SsEwP18slx
39v0m81memOh4Qd6ovFE4JMXJ6C5Ut/mznPKJvgK0osia1WNb7bf7UfNyjUT1jgj
KVdtmWcIBaYivG0l5cUIRZC2mAjT61jGZakCpPeiiGJNGM8kym1I9jPmKOHIx/yI
jomr8xoSc5+1Ow/HuDUnMF3PYYI0KWiPLcVc+U70bkxETYmDA6kPXbblrh0IqWty
TG8dIBV4X8PLdwKnGM24pqg1cbD5rcNBhG+/KqeaxnAUZdh3S1zGo0S62IBujgTu
Ry36rUXmbLJGpb2HUQXtdETTrQvKGla2G21ZihNKHikt6DnqUKUMsT4cFVApWz4o
1Ik2QTrhSUQhF5VMj1lNM8Ewwa5BYu81DnRA6gRKdkWk0+EiNNE8em4hdwxVLbJK
4Qtgwv4vV5HBE4Z6h9V2RdbrqB9aADk804jScSe9R60dbuzi5I7IK0bOk63fVp7l
xkSk4lDjyYfGQD8+ZWmzbi5o8lurYP+NIpbCLinFlzR0vT4GPyhKg3m6ESJz0dqm
+JoNsUF3+2LMSZf0g84bfRnTwvg/PDd9PjJiA16otcKd4LFmr4eUiU9HogAVDjj3
E8hbGONB5xXpuMbusQwhIoke3Qb65pT3tnURobBCIdkgeZ8O4ifinM/7MTJjIQP7
e/sdIkMfbofEV8Tx+f6yq95JKyikjBP6dNHInlOS0llIF+r0WVGfLJQX3yN495sQ
QuJSl7VNUvr7gHc/O/O6cfkf/vkbVA9iPQBL9BL+Ifvglc0rzEPjySw1xLbxn7Kr
nyG12wuau2zsauiQ0sn+Q3Qqid3Xj3F3HBPwKaHXLK6wnfBfTooIDzqLyZBn0JHZ
XPR1CDTG7NUeLSSV+rv6xoXrCSYHxggISu0ECAr3RqJq1utZIEZLJ5yz/IFxEUmQ
dyiDonzuFEshUxkrRIylUPJAStpbTWVLN2qeWcmKP0fAcfQjA5w/ksR6pfdFgF6t
xZh0huZZXt3upwV/jWCtCcLotfONEOnZVn7cFKsgUamWiXq5k5irXcDQbjTYvb1r
u20EkYgKVtssffnYYmTJYt3zaFedDrYBG7HxXw88ihU6hYTtRDe0jGouqhwF4nB4
z00cr8IOw3kCU0lpdznfChxTz+tWuzkUmC+jgTIvmDsQfGdUf0YY37czksHqjJW3
HL3eB9BKYfGQxfZcfZmQo8n8dbapGd9kQ6r/2pYjFBG8NZem74Kl8IclNjxrt/1s
xwU98ln9PdU4OYjhsoeWVoO7Nj4XoZgaDarVs3/Ic9Uh7ow24x1pSkBJ3Onu0cyO
sPkF+ffTLPI0jCuU6k6i8qHY9likDLi3wdqCd5+2u4m6fC0radkhymhy+ar0mYyr
k9Or761/kUoX9ZIB1GjZ6Scf35RYsJVeyFPi9tcaZ8hmQ8rjLh2MPoifRSVuAMBE
QRe9WlWJi6rfb5nkHQSZjzDCCO5Dv5ZPBA1nUdYk51tZk/+cDGXAox6Vt2KRTdh2
UUd9RSbHq+v9z9qqbNpDWqHML3MhUVQuGsqXpbLMEfRJDQbiLnST+1ESG81+vLQH
P6soOGwi7F6gBwDD8IPBxTKlPjAb3r3Gte1rKTyTi91X8n4Ajbp7dcx+FPftuX5Z
tR6o9QxJyIPBJ/4rklCEAmYAQt4tPciODD+HD+zivHA/fAPJeGNg11Ih0amqZ5xM
90I16Nh/rXNBWU210J5XE3ZxLpNpwVhWprRdBosth5G81AJx5hY8LIUZLjmXndnQ
RzqRP4L9sMWVzuYQIA4kZM0MGgMDG6e1xS78ucfcdqm/UVIA07zox5a2A9X7w/wN
2OO4H23RRSQPGYPVA40y7NPkj3u4rwY8k+3bsq6uSm5SQ0qom5qmTCsf7ErNN4kv
PqU9goC3eID5IpNGMfsaC7xGHUiXMhEP23vCFpUSHJfPMwMHNzWLFCZgm8QotyQ0
s868Z0QUW3cgCbTJqHlw0ACSvj8I6Mj6js/z+FD6PD60yxZ3vZ8SN9hjDc7XFzLZ
Wv0/aO8LYxITfn1iNk/vpu67ajk+mVtTbLViwqSIjVPYYmHnhWYgLHD9a4ymr/u0
szndyN798pQx9lz5XfPSrtrrj/FhW1D47j65AB0RHsQgbAMqEkM0FTg+8xeEwrs/
ygGo8uG8PKsKtDn6/yLEX60O3BjjvSWVex7OktU8g6Y5B/LJZn4GE22WX6x1HR6f
NXWO4/vItJcOfkTB/rNsPC5wzuZ1nUTN6R8vTbCFzeGl0oSPWxYQ6uyuulFnTqzd
V09+q1wkogzdJSnsGeWjvWpvxx+egvp2I8kkq+51dHlXOXxW3Gzg85PJsQJuRqrI
WatAreEeGmhJ+8kwER4k/8Viu3WxQeZl0K3X/KlPjaEqNsgIOzXvBLt/sw6fGzgX
46m4GzZGLTHRBFLg8OM+/ZTob9bHkIKLT4up/J2tyoe1csXtso5Piy8y2tGKnF2l
+FQclsi4sk6OK8lYre09M3ekHtCwTnGiHeYBomWwZsYeQCs+PSZqxTm0UYxTfk2E
CSW+jb7RPXLz2cb6MAvaagvGxCkeZlkgrMG5/r+YdUrsVTP8uNZgn4NqU4/FCo/d
zfh8Z/68xjI0gkCF1x5nU+TN2Azj7bzTMDT5h3dGV3kwcG7NlZ00i5MWytDeHOxQ
CTIEQKAkg4/Ijgm9LUB/5sZHHodZZen94sThvYxuan5PrRYECFZxUCUROrDuHrjU
7+IigsucFCdBr85fzG2oaubM4fdmY02oix+orz0j0DgSkHzN0nLaN7gjuEpqIhMa
K21SZN66RD+Kc7vlNue1UrR89jPTDI6hrLgtsudG2LQNcPDGpT/Vas/zheqM52oP
/3Hxzu0WYWjORcOLUs+Qa0MTNldYcdvlCKJkc1OJKe3O/JBgLipwgPP89R2v5SW8
7pwZzUI4jGId/mOAsfKSMEQDtwJsCIsraiT+ogA2WL8Sx9Gi3pnn1bKWvWd2A+nX
IcVEiSrRLC/lAnjCEp5ufMpCUoRTfcr3TdDIuCpAbQ+lpXSg39orTUGtQE4dkPqS
7HByX10Dkmp/WiusDm/NDSYFrwI9zxAjfN7zs3/7sh+HJFxTun2VNcEnf8VL0LeG
GohUPcJhrTdz20N6Q8uCrAps6NTpQqycjeUIUcJH401nFkndNnyQ8hWYM8sS7IFM
cG6fd+zCefeeiGg3k0EKa4k6Q/Ei90yttv0eiTNHLOwiolV4ljxgBW7W1gmsyBDD
LtJ3Cfj0E0WoccmaKxueVQEQqPvDmuNalqTgR1h6qPag0hSDn3tCEakk3csPB/L2
OmNtIl4YCiiFbkPWziC0Ab3jzncx5m1RVjmoFgVV6SL7t7FThlfJRFDEP5GA4s/6
x7+Y4yRhh1CE6/RaXEhVsmFBrG4kFQQVLptliPDXKGW9vTcasbsFk7hCfxXAHWVN
VRArdfyXyFQQFnnbZzEJpPxY8g3+Tpb+RhqeSi/3nRSrsGYVelRk2dc/nNbVrm9X
pm41N4Nsu+cexeDXT3DUmo2GdbAkyafICaJgh2bc9quhV30cm307oMh75XrfR+aU
mYFDKG/jTs9E9MTXJzEDdAkj7Hcvxidm/dmxENE04IfTAK2x6CVKAlSQEmYDN7xs
NtQbI9SpQTpaQ6NDvISsfuEh14rlAozRluyx6GrsO4RpvlscmxRX3p3hXLZ3hykz
8yHivzsYt8onLjkTOr3Nd18mvRwURM4CoS4kXn+0ESIUcR+HFGWzCorxnUugIzYa
bouUv35GyvhYDgZoy7pPAXc4MpxNP2cawY18y3GQ5Ue+hQqlxOglp79w6c8cf+Np
0etRqYPe3faUlqlxCGk7JcQ3uJY6Jw+JQAmkzOkTJ7uiAOuOg4tvJwDtbe+ZXBX3
jjG2tl3yUKQ0yXw33J3C3WX1ZZ4YiKHCIjEPSwuHTYmqTulsVoqOk3uhXy/bz3ct
RyUsmszdFpMIvQVvz6DiGltJtxm1DtbNC7gWPjGVxQpHsq0GLo5TgVGjJuxi44sL
RfweSyRGb/N3I/iXZ4gpWBbd51Rv7C3efAV0d36aQRpnSiJWxNAl1/0eFwdlfoUd
4+ary1uuO2HdHGBNqjHDmsJJVY1vfR0UtrVDB//kJ70rIQM1p0xSZVnmLN8wC0aC
isQ1M9YH02vvVmuQrMwSyqTopH9B8IjXbKKcwduFEEwDj2veMZbzpGEGCv11+4jq
aIS5YQZc8GbDotHzA3IJtZ0fkv7116EN/nWjCsJXPdDQ4tCLThAfKYflIPa75DpE
cyqNmpajNVb6O+QezZsiStrgQm15yCfLrK8b7921lcN+TbYVSYZOAC4258nJaJxw
rMAjE4u0z4+Xylj3VuPT3bqp8mXWfyR1O9Q6daeVdefBlcC6sBqoevn4RHft1c1F
JPQEgvIgNWuq7J1BxKuj/t3X0ISSkOQfYGWKCYarXhg+9au+ubGbi50HAsr/pnbF
NhgQf14STF3Fj1CAupXaVsyiwPfKGk5LFkVx6Hbht7f3hJDj4EgO1bbqgCcCBPFs
qghVt+G5+8T/Al2CLVGtJlJ5KEh59NA1phDCzb8och7K/0MMfsb0rOz/MErf7xeA
T7/u9ze9SadKNRYwibr2KKBUp+L/pyLiI4x1W3O5kTkQd0LOV3qPge5ujHl6WoCv
8BIKF52yiyB3uUwcnP9MKjHbbdFy2OK/pS0QrBiTJX8DqJJBqTHR3ojnEUL4ARO3
X2IYsE0wZxWaszZhtcsIvkv9bCmgcgYu8fodCkqcxlhCjN4dppkKVy0YOrg0qtHM
4HE9ORyTtzFNf6cCz5jvdeEabTel6KbPlBQkPhAR9lo3CX+ge9aEneY0gQ0u81Qz
+lMLE6MtX8v0U7Hv51wINCzIuiU8YEd+HSb69GZKioI8zxgsnK1u74sEOodU5zAs
4DiRi+jDhH8gpYCGYuRt/kGl9/hXF/fDP4pHqj3kI9ig//HdLQpogRwzjBiBP4lT
4cVoBlzbd1hB6Jv1jx1AzkjUw5bgZ/EHALe92+kv8/fmXybA+rUETo26mme8zFG7
mh8pESMSG79fkKR4jQ1a9JxSGoQI9FssPFiNhWiYieXak/vZl0ooKyofZVDaTN9H
9qRUKB+BZSAPSzi2e3VGWo/uPwXJ892aHWGmmlli8lYjpLvXTaO1RpUnxa2EFwG0
97Roy4Yu9G+2+MVvUII2V3KvfKKGx8z/cmhcLB3UdhLSjnTujILatdajf9gmG3qO
gx0fjScG06Oit64S8GEV8f5Et1es24dZXunuO5NF/5rtEhuAD0ow6OxVmbh8mNHu
wn1SQOIRyG0I9lwOiSJDAmpIxPHJ/61se/8NuIl7UyVs6G1w/MIKKfzmKnSzwiIX
wIX96DQGa4JYNe/mKwSAKcSHLjcfdYSlqOkWa+9gJT5XfPmg0npDWpWNgRXFGO3H
hj3LSCGiiv17m+rOrAsIJfKNsGguGCS0V7ypID1claoBJGUdGnfskxu2ocokFNAt
xcVu6Gy2uq3FQyeMYNvpzfMOrct6NsNrwFgsAn14QSnewYLhVTuXJeOXtSqpBhKT
ilq4iZpr3co2VldHMfQTSf/4YzYWYujCxh2rbOsPmb2Zhr7K/DpMjhvGOv8PwIV8
1Cn4dhN7eGCV3tDcvZPdxgxyU6ByaTYuZvXxmwtDuOXvHYKxPwz6TqMoMduWtvC2
3gXV9pnpd7j6DFYsnFLQ1cqnWfgfQKiwevKC918sBH+onVlMxGAujV/ngK6J4fOF
ioG8/U4NS5ijrqsxCXwZuE6UrzodgDcUx51ukyzeqDTcsg7+ONPlW1kHHzzw9/+M
iju9HXnt0TOP7kX6jTSTmpfTxPj6Qqk/HJ4r5IcRIbrv59VWFxwKHatKv5EsZvmP
bgkh6atq2eQvBOG6QAjvfD+ydeTbeb9LLgYAQpjy59IiMLEoXwvKkCyCvuqn9mpd
IoU8n/MlgV5F9XdJ0YzWG4M5HtOwpxnrMCs30VkGBzF9G+W6rDPMEw/FGywaLDha
u9MweIAkHKYyN1DQYnrO/3DB0ZpEEuSTLASAI70/fh7MaVI2rxXTqyw/GHX9RCuo
4Z6SC4vTjqr1Qrlx/sq1BqlO6xV2TZQVj18jcSQAM5mvCcRxQe9i27dr20TVwEJM
lMNpEjCHVPpNPLifn7+2oF3x23kcna2jcd/b3HcCpjs4Us+K2ooC8KUQHCPm8gLK
Rki6u/7gjbrdLiJtyxb97CBQkPWymxp0Buey1dtQefIbpdt2fbMW3UGoXX0VAH62
fANuWF/qAjPBA0mifAu/8LZj0ujKFObG7aBXvupzf+CAMbfrAH1UXKXAiHsZHfiS
7teosftMWuAQxczYL8Qur1Ymld45MCRXOZda2AFU69yawRKuYw6SOyM/epfQwdH6
n3VOsqTIl9vS2rKgYeQIxbso6vnfUYxjD5ovkLsxsf0JgVJ3sniD9j4MiyWTS4tt
EOpeH7XP2aAgwm6HvSw/Y50M4B7SZofHlRWHxDBm6r5ZVwqB4UHI2vzvEe0+AI4+
WPtbkrwnoAzO8jo3EgxqqgUyEK/sMHK+w3SSs9bflqo137MYKpLbkZ2eGITroco1
ruedeamiaKD5oKdLQx5sparc1SmhTTtuUL6MH0CAh6KvrqaKJkBEQluRbj7WD+Lh
TmregPYRniFJZHNy/wUQAClbd6/GhXgYNGH3ALJEaw9Ip0xMNibg1kmN6xm0XEu0
+g5n5k1D8PJuctwblvBTEtDcKRjy3K38beiAxuTDf4gr9N3i3eAG2/jamoyd8rCA
166tm1qRpmgm6D20i2oapL4eYLsYGn0XM+V759f4+te5w4AZmS7ylCb4YcziN/Hq
VMgNvNsAc8JBCKxJdGpP9NUBWb+CR21VX5pyAG8IoQqChiOLwr1/gr4i1z2qH10h
7nBLsQkKB4c76T3oZnKSOwsJNEpv/rhxAUSBbuKgEiVKHNVpxngJbTgwucs4r1ml
zXtsqBQkxyitVKe/eOdG6SK27SF5wbVT2ORxIqPnKDgjynDqXXioX5RQaCnev4vK
EDrfloswmCtpHZWJTriXcV89vr25VmqtFy7CcTssKt0Se1LwMpZHySQhiYmRZjiQ
EQMojCwsD2nDUqiRN0GWvy96t7U/OMQBJUdoc7DbM4NSvlUSxgjLKs/B08iE/U7N
vm6o3qhi8FKO1SG3lNqms9Wc2KrfvVZ8R51WO5BOiUx3UKRd3DYTiycRCSAmuPBy
d0J4UaRtYk6c8cb7PhjRNtaLlhcLP6T7M6k1VbkfFDU6ZoEcsd5wWVB0f4G4g1f+
iEddUUq902+Nu3oJh/1dzXrFT8iWFaxrTgJV4YrTuGZR1kFZgFKLN6W9P2+DpPz/
3fqEEglF0neOp2HttTyT5TGHU2yRvNBrEZ158eOGqrnOvywJ6fHeUsiZVa0tuyJn
q/DwuIbUjcS4FZqNoZyISp+rJ8iiMiokEjLzP/W2ywkPLboCzEw3/DnWjWEZrLJx
dOpNdr22SNxWmyoiVSFs3qUd/+YCEU5xi3XF56T7K3M1a1mNXGUzcgJqcnb3EewF
jlztfh+8R7ghrRzBZ5kcOtiXYRbGuN6/ni/aZOy3iTmMAHDGwKTXWZUQlpBL+L7O
W3PXM+DoVqVY6bHnhy+6nHtm1a2t0IUHbD7//7kZmsazRzjteaQpCCucLW0ekpaC
gdWQKt8uGwDfEiSD2EL9YrHg9PUlkiN139Io+1XzhGyjpfEGZDHTqsh/6fxt0vMw
a13bufpl16mZ7oUZ15/CwqpoxhwpQKeHYOoV/nOpVJVgIu/T+7Edy2RqnaM8a46S
oRXqP03CkI2Ag16ouPmfSyGvm+j5dQCnGdb0Xtq5sIImpINTI686NDvnS0c9y7/M
fwr3Q09GWFzQz6OoWI9SSFDP4RoTRV3/LLJpGCaunxboVbInlTIdOCIgmSmk9SLr
hqYKvaAvxjO+Tr3SqxGU6iEHag5NfzYyNhB4aiBudHtW/kyhxXwMm7WYKF7QH/zr
UXmYGwQyqavDCJRSlMxjmmqI/f4rtq2LfPfCwodPtpzuJjyo854cTtRifIZEqf1N
A4SbxjccwxKrN0UvpHl3YDziLZclWkSjr9WEXFqvgKTR9MD0IOGAFG7U4KYS4yZq
PPcgBd47cMTRYVjqovondxj5TQds0EG+w2EXOdMZLnQgK84Do3uWL4uO9as4RNK3
d00Bbi2reiYHNRniuH2ByKJ6KjlqeHcZ1Y0rnt9Em9t//1OQDjeykedlzMRWhJjR
WUHVggxH7wc1NZD1E7554Aqe181nj/HuaorkqHcXIZ+JmKwixqrssa8MlS++Uh/H
c1F8xsruBJOGZX8G1xXX9+0OCnknxIirSZfHkRyMP2hkJvh8d2n22X0RzuDnUQbk
TKRny8zxO7Jxq9W9L6RmdIUwnrxzlsGVaElS3b0EBNsOHxoEoDbxwxi0WhA8xhxE
FG83m62lMcWcUODabyPq3swIqvpsnr8MMul1tij+yPg1uJp3sD0y4DYDwfe8s26x
bSrQsHF6OWzooyW2O/0Y5ysgft8UYPHNsRKPHw/w7AwAH6+B3sDMsNOZjVYy5xoO
Zhfp6Zy8T9/wjal9w5mrBKNzjbM2WCHfWr23Y62EucF1NzlTP/DyQJ8ww8VZ+Ygu
S0x081anZm9q4w8sivtUuqpmr/z/NVZzkM8ann7EQjhY2oymAWV2eQDWLyAhc1us
wysyScTOGchQX0WEBKBDGXyGn7zYpr9Eogupi6KUTEiC3LJEhp/nXGVq0QOyCKb6
H+kBvb+vsITUwhYk4VRbOwCjDbhaCKe8lK3P+gpelWQRrR0tLogfaOI4/OI16Vu8
R5GJWU/AXoyGj+ah2i08vD2zjKdntG0CCMPmrY3eAtXZ68crR0CNhEZ89pe3Mo/U
dl51bM0xKkDHugpr8BFQFuqpXYRGzU9MnAtmZKG2Ts3sEEHF1/ZP4qc+5p49S2vp
NKZdLuh7pKOF/z59KW5BGwNSjoozKKIF6MIUtH0DyeE4mWrQPkXdS0nX7QqEt9pu
aAMVr6icujAg0Dic5y5kPg6kRN6x73YYXA86AFFY9+WlyvwOR6IiEb6r1mneh9Z0
JD0jKjcDwEP+EQ/oIj3K7agPir+hssBfVa2gA53cq3BBf/Rl7g3pdDyY1YotfW7o
vdmFo4bg3IS79sv1rQUUsYr7PNbCvgA8jDLVvf3o9RgfSBRtSBkHCIVca1WGsvC4
Rw0J+eL97YfOqCzFdTcK1DZnri5CiVAaDHi07PoUVSc/M4oTwAutPbY0vs4vNmnn
rlHrerFm/ukoqVx7544rnE27MDgmmmGaG+EnEPDtUkLM7GZ/9381vYksK+DoTc1x
vi+FAbsrmkEp1ssfSVu1Y1J2ThCNK73HLLVpRUcQhuLVkhaGBJTh3DF3WX8mk7pf
ZTp0ECO6P/oP/f5K/wea+MQIfRgTlAGcvFy0QJuYRAUidFIyAJvQYsXu2Loq9zNh
f5LZvcrgzmaeYDcrMiXhqaBoKE007mXF96S2TikNanunWtnlmd/+jikwarL0n2o0
L46jDp3JO/L6DRHWdAdzoNvtN5YfcvRv3uKTEqdayIyghXYs0uX4/1sR3JaHlFf9
O0EY3yHr9qCopoH8uKCBs0wMY3D1V2n0QKxrjZ9bvT7JzehvtDPDpBMhhc3VbLmo
agANRFi3pe3fsqEu/FNl06EIpvKnLqRjjsU/5rF+8xHLcxD1R+CPNxW1f41sqjnR
qDnoP1TOhdq6CboPeFiVphsuqyfCHQ8LpBpxhymexoq4STqZvex2rT51WoivZxaM
Oarax2bIRTL/8F4pDR0adZgYLJjb4+IC2KFKRQUGr37MLNasCgZrkwdaruIy4O8Y
xT9mEFRy53treEmNr/qlNXaB4e7Iwhd1R/v7I+9I5VRo0vl4zZi56O0Yzi+B6zLQ
w2c1ukCwiHa/E7wtxV0+PITlRLx/HmEDDH3e9WRuHIAF+5smlYjKAqwSfaIzi9w8
1n5hwK+ooXkSjiVS7NzAXRZIM6f00jwR2ZN8p00RTsR3v/NZHewyjfjhzgqpo8Ec
Pit4o/72XWd10e/5vnMTr5OwWar1mGHke5vbthKX6lIFZUJjI9Qhb+CZhfTfhn3f
TAc9qDHlykn/IKdAEm/PHAt5QP5kzu9GyP1N2lcfcJ/u5uRGS6FyuR/StoCFI/FR
4CD0wgzdWAc5Sn3GQLAKMWyETCfxNs1C7Ho5VKSjekGK6zQvDgK9dLEhMtYb1jMP
EbHMRdbvfwpAdcKrsRuQRYxdp1qEL34UFKUzp/rc7TJEfvqePd6IFKEihcTVhZSg
zm/EeHsNgnK5miZ8pIODAOMbQSuNs/rxbLp8ZoeLpAHaUPktdUttIF5Gtx8AtjtJ
s5Ajw+foT5ruEfDe4u0orVWzaf4xBvofPLmN8yQsxDgavbXz0yi43tnCZo+KNMKm
otSqftSDD/uAhcxllN2y+tKxWVHOe0PvuMKTsAtLJnAcyXu7ucEDoq0H4Bu8r1vX
VMI/fCA/E8ms+VGAsH4wg/GxgAMNhTm24LtKrKjWVurQ1x6qFY6NBpVVtq3XAZx9
bKEdwdizNQfXv72VsROALwrf8WRMmVGAHcNBtB3egPuOU5brkQYdDAmBFiotdVkj
KgAbjCC8Hz+3/Vl8RSIERz/zten5pH3Z2AHstjBiI1rPm0yB8VnRQ6zNqrOVS5Ly
HmO+QjGHBxHARHrlTQd6dJtBrIKJJP7ekjlLuyOiHuhm1l5qqo2zMi/qnJfKGIbN
/wBVHYBQjSlCxvi48HmOb2nbMNV7f/8W14jPszJhqXuw2bAZD2f2aXLKR1RcMlkm
9lU92BV8b5tbhZLQZeVNC55PRSfmctt/s6pd+/3sN+2bujxjK9O0NbOKC/AGozMI
iYoLj58EpgBb1lAyVznU+YO/sbGAinYtlpXv87PbWREYA0x4flDhMw4u7BQGDIxu
sXmFuQqtudAAmcfFn3glUwnQKQnXjiajPErmPESV2TEbtD/dwZEh42wgWNfIvpK6
c9+7Nhnbp49LlvP4ka+SAeRJqTuzm79TzSpi5QS0QjEcNrdGZEckx0JUR+15jSFL
EflqnnWX6Qrtz1h6cR4YLdUa50V17xPKmKpbhF2d5NY8eD/K4zo0ek+VY0Dr1MUG
p3i8MhOT9ygdBlWrpS4h6g0YS7Y2rhnuGc01m9eC8XR+We8Gdy6DtEMiktNhskZ9
2nEMcFZEhVecQsMnK8Zyh+D6Md8GtyeVHFN0ZvcsQKzELVm4/nfWYDsLerIpSE2k
K/3eb/Uf2/JdeF2wF07ElubgEExV+8En9gSzw1aBRuPNM818wKnUkotHcDe3snwT
Bt61C5QF7Ve4IXIIYapQVqDDk/Mw+ViCeyAshrAbWvcUFa+1/ZsWKEVgsVYfLuPe
1W8PrsLTEYdcKjAWi0AGBKu7l2oVpoZQGt+9+XsJuoccHo+hh2OpXrM59GQ4iVjM
cP0wDkJ83yhzIg8hkQc8VYrnOx5LPnGSOyW0tLyceXcmpNIf1EnvAwipY5I0Edtx
lwxEEF+PQ3RID93kwe+tH2Qi418kKJjrECBFi7wLTsgtW+RC635WeDBIUpcCik8A
7uziMsowwpC7k+4/twq1SxP+nUR19Hymf2wfqP6YdAS14s0yH68/EuhkVLQMWM0z
qei/AF85RjZgCpnPKWUpIPDTSL1OBuWt6p305v9Sco/PfaYbwx3RcsNvb+mR1tIR
8hnRhpkBse8IfqHF6fzPvMJIoq+PfhP49I7fZ074W8QJHPJIJP39VvL9LWvKNoN9
7FOvyYKpMp1+AXPK+BPmSJIqdle82aSp6EB9MF3CgUxsGIuY4VsTrdEQiNaZ1lO5
Jg1EoHbcZgrqmDyizjysnYwDGKjR9iI56/OEtt+3R2mCOc5bi45L0/ObReyVmB4C
R3DgrhZfCpu0lzkk7Uu3n7OLM1Z/ArOYt3BXjR582YiP/tTi/Blba8Ak1npfHvb4
TJPlp3ItdK0SSzf+Rcn81PYSk+MLn6k2NHhnVZoVMukzRORQJf/Q3Epw5swLfoZR
5TtISLX8nqs9UeaCMADvxN7xCg3ihrAKMzPTjae4WdwD+qBUXL1iaxIEBx3/vKy5
8gY58uGYlsZdxletTLP9D12BkEEVbThVA93zf0dlsKWNpdnJa+9uJ4HvTVQtFlQ0
NEmOF6K6ZVSTW4qWfcFkOn2fY9vY/tZgdNedbYdaxK+rLG9ZaxDU6eAlSF5rrjoe
TEwevPV+cC8vSXth6CDUObCxAgHDYTaEzQmslyGv4eUF+eNU5IikxtZKQPxFDlRz
WfNFHxTt7jzujuMOugD5GE8uQei4X54dEwFQpG3mFXjxk2TO82WzGmBoW3Wgt9Ly
Bl22xd+UcL0s/mFN35G4gDd98KJgJrXL6MvkIXD6c39evLa/S2cQhC+6rlT7pqWA
Lj6PelvoFkip/4Hw61TQCrJ+49lfWHwpT0VQbajHz7vGYJZNqWw+jo4JxCgg6v6o
zekWyvRcwD9ctzFV2HNqMGrJSwdfB3uYgjaOt9XTgX883AvY+1O70dJ++JoQHyND
b2fLk8pkfB3CfN80okkYMQSiEnWPXQ6QmmqbKCtgKd2Kh4Py2t5xWd5ZiZqTOQq4
xsHr80XwR2rOXLlbWX6PzkpS/N2HugX67SaOqRRNfSeqtjIzSIhas1Ut0euexCq2
DrXCzIhpVCzDEES0txQ3KOFLO60eOEAe/QhsoOxUS6rQl51Mqrzfh2mOidKK1xnE
wEG7CjqZtVukUPuj65yJQyIZm7GvtGrI2QH0AyoIRbxl6y5sgKKuN02VQM4lEZKN
ucA6QqoKwmRfdQewK1GBZWiEo8vJhNvefPc86gOzwb3M1Qe3qdYSD2XDSfoIVmtT
pmBRnYeteO5MvfOoAA2uCXrYraLJVUkqW2QZKx3WY4gsqwNoCkF2Hxyko87kiETx
p1EsBvjBPfLRjqpAj+dUcS9Py0zdCn7plNK6QBXdHN5e9CJu8eU4JXgGqqcvP882
55wcXCVHdw8ub6mXYhy+8ub9Tsyu5B0cita+J6p+Byre4KVb5pozOZ+j+81tpbb+
9XyffyNGPoTrsuJavjOHFpxyw9ja4Zprp+eDIrjRy2Z6MgCs/78OeeY7Py+qIsI/
MaOWPQN/6BzjDmqgv5TYoZ864HInKNqPR0y0xPnSx/826u3YrZSQ/p3EnJTHcYyw
rPhLFfA+Bo/ZIJ0ab3VN5IRihRpt9O4H7WtO4dUrz5G0A/FQhIyzSIyqW1Sib/0S
KMlPtacVBmnKqiL4MK5RZ0MbDKVG/vWetApVVYSxmeLMSLaSJmnvir1O5qi9Kv5i
ZG74W/rTT3GyUz8BneAXTGwQUN7IvNtkBofkyJGFmLop62TlJnEEJo3Qeczwuws5
fhoGz6pg+8am9/88OxqtG1vCAvAb3uROs8CZiIA0hy5e0XBWQhxQKGMORhfueynU
7JI6JjZfQSMxfagcAr/bp5lYda8jEVDs0ZM3Fyb8iE3C+PqP2WWfasdf7H29rdrs
qCuBU/VqAzfJ3ENL9E/YjvrBlohYH8yCWcCYr7KD7aXjIQ0c5g2ZltpTuJNkUMN7
fLzfReMPcsBd4Hot2mnVL2THb+lOEtbAi14DnqfWJwFfAOIZekY0uDkkabM6Lpn0
0ZTMjZMBUcP5ve4tBIznPIJUGeqGX3Wde1ejF41TU76G2hAZlzyzUHKFpALwnDql
JeIOsAaasHodQOflwmTjyoXeVa6/N1Bv0BeSehD/O2/Cz5eWaT00/G9FaS5jP+1I
61ig+MKTCcF5blMoB0HwHs+rmqPW58eBlfT+q49PFOtwfhL8P1LJzd7q+u3UD9wF
FkTnCRNzSNfbRWn5lejSqMM+0wnO0ZjgWnl2pQFJnj5AwU72XqLXsuC2963WtLL1
Q09NTYdKJp6A7OR5lv+Ng/yn4Fu0jHLdKGldP2IPOS4PUynwQqGHg1cQNX2npYZr
5jVU4t1l8LasEHV5OguF2823aoj2UdP/pYGbdcf3vn9P7fLNfoADCbN8AsTbmVGj
+933J659aX755Qrf/4WwP2IhnT/Tuzpg/KCfzfjkSxUBPMZsRBwPFbIPixQbKgXR
Ewqv5yMP77xVkl0eOSogHkdE1HXOS7XO92JqH6DNdEwaf0+w9YSwXYhC43ekFM3k
VXdY3HbedQtlpTmTx6VlVFmBYVkO+tXmRseZoJ5+I5JMZAxsetNAD0xvSkjK8Liy
pBwkdImlOlpu06e4rsX8hVd9L+8D7DcMm7gzUNijCsAitUPSuHTqsbe//c0tCgia
CsWdV9O+jmUAIkejJzijrpNHj7Efbagu+8vHDE46Su8AFijhqu3uqIQfvauWlO+e
w7R6FICddclQcwXDeVCYoIlZkLJAdh8Lg+CeTCYWmTWJH/DqrXZKpB2LfFjWGEIk
Fzw6G7FiF4DQ6hSvUQpVx9INDRjQNzmC29gtGE37u3kQgU0whYa+qSx1hN/qotZG
4BrLaaTZzV2AzZGLCJmsRE22fgxbirV57a2E+yfdlPPkYSZF44ryPMNtn5IteXn3
e76QO1tGdQdSAsrOjPj66Fa+cNS2RQljYpu5peFZVvMfArexTU/OSPPOMRaR0hH5
8WRXirK85GH3BPTdkAzOh2VvVdvB2E83ANEnaGxWIhGW1+XaTIjhyLsUETUt71Ty
1MAC65HPrc4IQTXkiZ9PT4t7ZTxAUVVS4bUE7oISVwivrSbNfHeza5rBmKzgAnk8
lBvrEr+k6MXLrz+4quo+cnYO/b6DCPWYQIqkdYl5VGM+TQ10oa2MFSSlNt9eFW82
48TWQSlq1GC4y463XYVNQSeqnD7nbJgc6AE0ts8HOmXhwgORao7V6m7H68BDr2Y4
GGnc28Ochvx7rHU7sYetI4njyZg4025yY8JufDOWeXDY67l144q9qiOEhLytDg7n
rM3pTdUos+C+uo5WL4sTm0q7WwYgme57QnFM3oNQVpcW1KbTwWtpQk0hobfvtuxK
y4GfUidqWLnuiGJf9URu6umTZDw0StBy8P8P6o5ey6gNLjDKqCpmQVvntmFA5ToO
aRi1uNboXVrzzDYJdzmRM71B8fZAz6P89ffBUqThUTuLXJisyboIbJiJBSuwcAq7
IiwlmiCYhP+4TiIE3fjwlKVubhVoVOgbATA1iEx+hTULvGL8vQhtS8yM7OprNktV
a2vYhpdoPI1Uu9ikathFfxV1bWmmWHrQAPb20zJmxREvEICbeagfY/18Kk/bVFY8
FFuXnlrhiugHtZfGxdzdCy68/2rZ+Q5OB1Ne7SOtEXQitlZ/7axFpW+C1ArsLzQ3
XCCkfD5z0ijLGE742XadmmoTL99z2j3KTqzwhrjAVNLo3+ZHOOwoL5+4WiSDSCPY
h4oAox0Nmi7CTWd4f6UBqzocFn9ILpsSVwz6ADoBx7+KusWQPV7cC3Gu8PHYof+T
oxXl+qx/xPH0ilXHUA3KFW3qlre5/ivioP/X4qH+/b1uFRto1LJdpNgjbeI9wVxg
UT2vxYQfRLC9O/UvuReJEN0KBeywDhqdN+MNLQnBO/EfhUBQatyRq0QbKwcGgqga
2xFtPVYOi5jZK2YOSu4qR6AzyTByt+YHfPmyxnGmuDxqw3r0qwD4SWmWqtXKsS8M
EF1L5Rkr9wTrT6tcwy4CPGdlE/u9Ta3OunzZUVmIlasZxwrepLsLxz1SdHQ2x4MW
n4ufc6lmqcjAI89m5tl1YoeRX3yT/ph4/59WcDXljKF3H3OnqCRZofF3OaBE1c0n
NAjDXKNObaNYvwc8B5eP7fggSY/F/mOPsSwSfckZSFPrAV6tn7BZ+VlkbCLP6iJr
iaQ+pNIc8xLLY6j/IO1rPiV+YGyGAJ1Lmp3Ko8efnYQvtpddsmE37JK7QoOMzKAH
wL/3ZCTSGEyoZlORSHUoKjQh0NhXdPEK6NK8H1K9dWGclV5UZMobZ6bIdTXdh44k
M+89SS0uwPkF32cQAkW8fa1qMQZSbtAUISO2tUgTLuzS11WJfl+KESzF/toXWdCo
+45VdeBHri5Eb+ToAVrjNA/O+ChRliGlIuWsfSggRHHJRkHyVZe4c+wWFwlatmWV
MjoS4d6DpRv825TxTvsaen/PfQIparfem4iKKWBMnkkF81BrakM6IPehphGzS9lI
PJPa0Bg5puw5p9Gb3OVrjFQNJoFfySbekzIZ9EuoOpTjn673UCLZDJLUbmMd2Px6
W0t0u9adGhRCiA4am0i5iML60lfmf3CDRHymPZ5UP7BgLQfj/ZjNHJR/csytFC8W
a9FAv7vy0EBHzC3h+Nz0Hiz4TsFm1YFCFulpRP00VlbX/X2q14MVoH/upP2ME2js
XDebi0RTdR4jqBQwH+5GLsc7dp/N/VA1ywSsCeSwSTwh6QkJ5G1+G6CNSMdDbVKZ
7NAfiKoY7hdwzRfgJ3Po3TQbUCsZgPQ2QLZry6M5sq6ZmDzmdoxhbPhbHZ5Lg3Tu
o+fjC0lETb3iF8tKLZx3rj1lgba91paKryX18L0LMb0DRfXUErLhvjHkTEfZSadQ
2Kg6xXg27XnhLYR0QMhLfhhsJyqEWA1q5zxlc1gK0SCJe/uUwKSZe207ZtroUxC8
eoVrSyZxHsRtlnHU4HYPCncgMCVMG1KfXLcEUIEoHp3I4cLqvKRihEPVGYLV47qq
U/sqlLSomwsMw4/b77xNFqM9vjFneQO54HluvKNkrjE27gm5ZmGSrCw+RfC6hfR1
P5gQjIXQNs3rr12Ioqw0pyLR1LN1NFAuJKIsTqKSjac5FpvgOdYMT1AB+uzvTo5P
d6O/b5PxxjSxnsDOST2dIXi8NDeYe95w7NFAXlPBPCYrEA388U2Bhy06hdN5ws4J
Tdz++FOEAX/s1e5V44/2r75Phlj5WLURBxvMy1rQsRCoZbfiUHSlZRKc/7uVDRM4
Cl7tgSphCreemyS1lCOWgb5BaqHappNy2X1l+32wYstqu59bkGO7qHZer0o9wZuI
PAK8fQPovmflvfkXq1qeG3STw81fZvxOHbNar3V5FFjKlgvSq9l/P/iuQj4X/uaK
3T+oOcYkwZ5ZfVOb+vc967gBVM+xMuqYcJWV+Hn/THQZaJ+NnjwRKM56krDTgb1o
e+lJh8gTlBQLDNwrKDAwD84MdeKOP3Ngnr5NJvyVECimrnCuHiQBj6WtLSZYC3EY
mRh0iSYqcfT/r42Cew+sgw==
`pragma protect end_protected
