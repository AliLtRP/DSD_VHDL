// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
l7VeNcXtPhIfYVDUZo3Vo13wv/2NB5Kp5aFU4DEGul0x4Wgy1VnEtO86SVzvOJKzEGePjGrIiCee
WIGDUz5Zt7DrMUHYBZVJp0eWpLyZwX5ftnvBfFDbzEnnlrx3cLqilGQ88mZr93LYtx+CJGvDrz6A
7lxCtfWvFRyZLTZC03k2AXav9ueE5wgTDmaLg4rZaJecGb5D6j/9AsocPbvAsSS3gXKYrGmHp4hg
JWiB5+7PU2oEdfP2znLSe8C4AyVhhKROJPNdY6jEcc5c++fwO12F4Fbq3tSxg7tV0j75VQGBKw+A
cr+AkX5LstWzybvaRCx2a8AzjYQmOEQIdGsoog==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
+aHr6beOcQpQVtPW2Sg6rk0zghmMWZYd4k0LuAUE1bjKMm998TU/JbtAkUGDpszjx4gwuDsYDOF+
SbyL37xIHXRi1h9YwWZEUTfnOttVje+7DPlLQ/czSaB+OVo/zMZHMTXBGRFvd95AWEqns9c+g2uC
beryX4Rx/gPjChD7Z7BAXWH+3t4oNSAmv+DaCeA9BUOAT3K8VLMoMwrK5hbDIbhCXm2tDrxsxaPk
ODqd9kHyciwVe0UHLL/dqi+tomgLEEUxUCEMvmgRJlt8rZqkVAFF00Opp9lF4K1lNEyOfhCvgfdv
7IeIkCYIkxH6a1jPWaGghUkmfsq7xZXf10SYR5OfP5I+tWlNzPAK6H/dJUiYwUFjRfuWDX2vD1fJ
n5n5KK9sjWnfLQwk/Yb4DDRAPu5dWu3SmBn2MLG6iqDMiaDS2eN1zlLkoI8QsaS1HzF76LuY9jy6
wefkf8djwMmXBPGEArFCPMctyUP5eNEX/feUknREU4OX79GW8d519riJrr/7cmH5I22ZQ1lFZBLh
DVxooiYy66qub0UJ8Ms93MrOBiNXIfnogv7HR4AqJWcO4bqnSvng8K6GYjW9Oo/N0PenOM5IxHBH
PjBMXDPjMShiIU+iLPRej2B8KuyQYaAtlcCzxU/+RBtOKf4Ae909besdW6nf5863yYCMI5SP8aPG
ZGAC1HQYEhejEFf/hb82ddZ0YcNsYIwXsEwCbHdkHV5DYvONgUPzrwq9Pknsn8jTaKDMOhz6dZ0O
D+2mtMBt78WlgkXn6emkAlQRJKjiYaZApX7IdSathLY772Q3ojcB6N1QTzIgum+Av+SSNIDsH8eK
b+TqAyo1cs2YW5ZokqaUjLvFRHttaVYg0VV0kF6E92seFDQifuuGjWJy/mWWPhUflkolF52Iix/N
hQrJA0O4rAMHf62VO98YwyRHYxuyFavp5kAHTLMjm8JG0fJaYEDHaZS3afPEag411KJ7aqRvtIeD
Z/NOULkDJ+MQrQLl0iw5xMdvJYzuNHGf7vbqbH/+Un9VC5AfkbJibdYzNR1Zty5F+N6MmJWlKoI5
KSK80t0isIv4WT/2Co55hUVuRuTGYguY8X07qvXGYvCc0YY+t9GFFrpS6qFe7U0KsmkMl+Ucj7ot
s8isDI5YrOx5zlB2JA0fJLX3gdUqgaLzBHEyoXNBsvdCH5cxxL9oDmV28VLw1K5TgYD8cl10r8aQ
oEjEGx9YybNXVuYnhGGyWEKrron2bhREZw9q6dA/TgfAuThN+rxPlYDR4I4cigVeP8BMuTrfFah2
HBwYb0ayvfY0w7UVT4HGQ9t0sEM/e0tQ+G1jFvcBBcYtiKMj3QKowkEcqpOlHpQNkcOQR2hM9MLG
79BU1qJniuQl/B0Y34t7l4c/sgyusvt/VKPyChHbFJe+KLjmhoYysYTwbWX26eKDXIdvUoOIZ0jB
Sbt1LwJkLvmV3f++MQyxWhMzOdqx53EG2/UPKRC3cfX0QcErcp2/ztkWyADfuZMKwzXCKadpwRTy
LwrpkCoex85avMyD9bw8v33x1+257MxTsQkpo2WANuGIPonIRBIbDCHlr8EAxCX25y4JcKT6spO8
iAv38jfTsAHnl0OIFyfZs9Z+UFDVBM8nLjD6zQmvxDR7FWGohY4bJiDYQoYyssZ4HNMzsqOXf8BP
z6pcfUBQ20ceWr0lalYZtX7gHc5zNhzH5/Rr4nxt7mDsGhQ93siMILqPD1xUfwHk9GjoEuW1mL8Z
/0ygJQHsB63/PYfwYrZCyoYeXOWriZPalafS+SgMvdtbA18VonUy/svT6l5TwBh4K2n8SEHxc6yZ
yFBhv4nIUUy/AbaZJMPsNdnJam3Ui04tabxOxxVrwIHKifyxCdAiSOhWPUNdDFEMGKAI8l0NC3lK
Jozmy901uohWhWzjAM6nA1h5+UF93yuiEYYXQfbManoTJWTmrA/UM69ZBV5idD8K96hEZ2YPuEX5
xKK7jYUbaCPQk1+Ck3nQTCycEWbH/SmS8nzcNQfHAtXJ+LLBTOSOmBBXZznDp/CJ1f3XTMXQvLTf
s3iakCHY9aogppwtQxcEkBuFH2LFVAncOhZK691MSFsTA9snQ+SuQbNf/ANNyXObk7tM0+EgQmVq
Fb54QuFe5wO1yAyrqZBO8Indj5IUPuXWWWvltTToP2uVwABnUW08FL6cc8Sc2W8AUCEpx/MEbwrj
4qp6VSI//qMUL7JRlC1fKB5P08iCV95zDRHyDD1ari6B+IF8KGe7c4JyjAjigMR2WItxyvxCerRl
h3DTGJgBHC57F71M/J4pQSkhjoySbHbOQcM2dVUiMNKBjh6X7Irr/HhdFIsFkCnxkgIxHC26UvTv
tuSYXPfjhKkNNJFfPD03FGrIYtUD7uZUEfDVsGkwp0hsjbiD/ApNbYmVj3lR1wAq9qatMyUkf5iU
ERd8IFXwmKdSHtuQjcCUVEu/xJnJZnP3Tzujej+By3bnDcN+8xaOTGMgFs2dHor8GEnlxtXrKGm3
LDko7qe5QvTR2ZlHRs0rNft89q8RZl9UALA0Jpy3r8X76fK/Qh2C2otRvbNZbxdklcsiusN+bLcm
XYw6GKKe9lhym3kVyv+hmSBRqLK2/8IgvtbVKji1ZRwY/6qTZsi29TqhrfXuyrIQPyPtZnv4WoYM
3kwHTU3++FkvBujPZsZdGQRwdOnBs5AJrNMBVVSXKK+42mLo5KByHn8Wmdluy7IB6AafegmuodEb
uTmn9kc/F2mB0fDKkkWE2ouTozAFmXA0obY6Kcp4UWHsk5bqETsmXX0ugzCrDrkFqLScMzuCyo+4
Id6nAp49XK7cjwQkt3gNyIteGfKkFrqJb80+J8IHNoZEI4Cj2dSSNUQ+l6vxd8fCP/6uikFPpiy+
LFyXNCf4cucZyH72s0qheDXJrqNU/eukdTa3ni6ahtZSnJT1k5wI1UIfM1Q1P5Deod1nGoBdlUAN
G0YgJbBKnnTfFTdGih30k06fkCnEMZ7EQDKHkoKq1doDtWyeAe6mFiWjujaTBCD5+yG0ZZWVabjJ
/SRX7hzsUPG9jfDp7rWA0QQDWEKy/fRK8K0bZjJ7wPs2kIE6GRUBN+Trqr0IbWL9f2gmEMtZAsbg
saYBuh5UqFDX56tC9wu4f+2p2cjHlnnrIMQtNrpWsVMhtuwINVkfJa/mGBQRVfN7Hfw/WepJyaI7
5rRftfUa1OqFq2+BPoMwUr+WTuqDn2bQ2Iti4X/lYUv3+sEQptbZ9ruuf8Dg94Yb8ZtaEoiheqTr
KBr5OV33+Z5O9y7q8B0FsQBfImd3Zp/itq7+YairPk3e+6WkyhVC3YoY0YHwOZtH8H1Dqo2Si8j3
nvj0BvR17jO1nNWRKZDmUv1fqDN1Fy3cJOuQSVWC6xBmWHXoBdXmjzEh3lEI9A0BW0nAKAnlKsE+
sQBVGGlShvNLWM3QnfJNJJK5raZAg5n3ywpAC6hWjsOmOLLgxvSwUTYomZ0VuQ3Cp7r+3NlG0VoK
Ar+VUbg3ZT3hG5X2FXuk1fEsrH2PCagYTNjKev+n8xB8AHhULKsXB2Zz+hpgjW3VQNx3sDJHST4a
CKEZoeaiikqQ/O3gF3CY+W1Cc+t/MqRqXau5WG9fxWuTbAPiM3LbQX5nl07s2ohKWkG+Ng7ZcWqq
+CPIAsHN/RiBCACeHQp/lKVyggDQH+yyqLSMNeSlPtDMSMqAl4hOMGUvy3RLYhrzPuMICUqIbnl1
5nA3w3fUUDILKMN9Y+gQoc0LMA+izM5hCb6fiYu3WG026YWJvC9NZVQGogey+ajC8lRaKw4ijSKD
8kvFyOeqAbMWHCYgtN5B0mvipgH7BpD+JrPL6C/ivTq50gZ2X/NAEJgEbdxFmTuPvH/iucJ2MiUl
yJ45tOpcfP7oGsMoxaET74jdDGeLcIMIBTjKhlq/LS7qxM6PGQC18BKtu2dT55NV0miC34E27MZ8
gizpWWIjnrfsgY1wHQxm9oQ9h3+ZYiWZJRaiW8E6vaa03t9Yn+O93bsauvWUzuzqr03A+2IqdRXR
i3BP+0H4tlGQpXzC0K11gqRFSMnNnw5Q57ytrSyM7Dmf/X5FWF1p6JLi8wPG10wFqNDWnQPVdP4N
fAUCY76KQyhnhYNJ7MH7rbPHha3Kdn3hdBr99I1fOEisF25ytB6Chk7mnJ7o+yKVNNGM7tHQJYIl
7oN0VI/RG0dPktNGXo2MwNo3iHcdHFyKxiPZYU+FwHnSCa5huohgxM1VfVng2K9Vl8qC6hAAw4+I
Xig4F4AmUcaFuWpWSkmXbIGAWGd2rDGBezqCYY6/OOKlGSxvwXOb2TJxwKWX598XwKFM+T4hoc5e
51wXv9m01ikAUUW7gYF1oFEsSTBekmNdXuBJSXVIEcosbJf9LldJnq9bmWc47u2Vnln486wN57Yw
SzOb3XldnLYkcEQblkQHR/vMcmeXx5IWD58ptavHeDb3iODr67KpZqIGA82rh+QSGTa287vx+QR4
4IMTJvbZn+bO5p9R1PE3eXKsWcgXAdNf4S6NF2KBLBLulwobvvAzaWLpVyt/CBUNxGLOs/IdQsB4
J9Alj16Ua6neA85pimW/uhvXja3FbIEm9wls4M6/lCki5H5CCuOkrezrpzirxv125eCG06XBpVfO
lzqE8xBWxabOSqs942nUUX8NJ2NNqWfw7PAOtdfwZEGyaFr2KnG9hhibEBu/4s3Y/jH/UnW6ya1A
17Vm8w1xzkNQOv+kykvUWKTn9+W/jmOVoXy/TTyEygve7U1O3/HTM5LjFZqtjYj33PpPXBt5d+Mc
7dIwBbLGpvboHr85Dwp9hDJpGF9RTAhTz2a59FA41VVZ2msVOR7vSGUMicn18vTpG0qzOKQ0dbtC
oz0MC22DirQKF40EnE0COQqywtCuLiypAY0vHQsSdCTmWknTCSY6QD/KwbeQagdyK68Q4P6JOMWA
YIKQWNvub24w1BJOt/84QuzZQ96ZRfAvpeugbywsjoBlhxd4mGoRetM1sOv2j31XwW5hdjwholCR
OBhage3rBOls1OvkMZn3D5gEAy5MZJ4zsCdCy4gOEE9snXMuvusWcTEoe3hatSXnvmzoF1OgZi6Z
cSGV+vNPDw/89rMgNW2JRoiF5nlD1jeQA9AxMw198WdChS8ctK86FGbPgT8CEVa/6cibEIjy7N3k
EH7Lhn6+l78ubQMkwDScIz55ANY0UhJc5y8ku1NsJkTgQ687JtkV3qSJKU0l2yUZYPNUxXXanQky
RZ4VbL2fqz+J0zrrgRMLR+oUDqXEtalVz1uzxZ8F4Vvz206WfNhCFyalEdgkHp0sJQkKm8EXGynT
mCpCvcaIstzg76m12d0Sg6F8eXBLAmhesY6qhi7W5CbHmoYQGItBwY6ITBI8uGTaU7wihoktmTf3
pwJDxXnSRRtj0GwhfkNa8MUXadQCyVq98w9bkJzwjvWGxKNwmpzVfxgthiqgujTDIiuX1Qzlp4qZ
uuziybLydHMWkyctP42n0L3O8DuE82HSqzCRbkqzzJeo5oAgwydVxLdb30o0npRXJWS3zMe8cjKL
tEtXbkm8+qD6EwpA/DGtPPwqzxwefq3y/xps82lZR3NHcCnjMNR5eOBZSNdBWEPedk3fXS+EZC5Y
0am5lf1hgzpfzr6xO4Zk031GfwLtZjx9py633w6avk7oOTi+S4RmIDq6tu0adXCTePi87aGR+xxX
+h/vec55e5o8jEdVwTdoicYm5wUnMldH4u9P/k/+dcR4XchMjwYdXtFJ8/2vvw8aLUf1PHi4y54l
0dr3WGcvCrd+XGzQmQy02p9IXWqb+OolFKt1E63S5tcEwBRrksPLW8umi8xRd5R8Z2Uq44idhrWu
vY/lk5N1c3kPrYDdFJraU+Mong8CrMNzzIONpcaLk91kvt0cPFsgynqFP102WNVixawX7i5lHnv3
ykcetkEJKwBYlLUC5oPJhuOocYUX9byBICdD/xrVsrmUuFSSxNpXTcTiBOs+cPZpwKqkPaEifxxu
6eaeBQduS3M17XYMKjLvPibY1BI3dyZlCpRdNmMMan+E6+CyWJ/M/+SoQhJwGYsz0ocVCN/z3YBR
zxvcXTObmxuA61rs3qUfFAvOBVkm7iMl2X9M70rLBh+L6iO6SrBy6hXQXKtDjMQwYVQL1uBvhn5X
4lkQmB1ekUTROJD6BL0RcxxXZHeYhOiGC6dVnlH09sGMOR7HWi4VpOTIjjgGhWRfWgFqJyfdtGqN
qx/hWpMjGygPUzM/3JmDF8eDoyRMyN7oxBsaVNjJC1sy0RDdgJ/xDiIMOLgs/9SwRJpjQXqmy+ot
Pme6vXTID/Jshb2zUoJcGOXMyMFaSWdcPXQSGtkTQa/JWxm2NlW2wJCFNtJJ+Jf5xY3IpA9m7P2r
YjyU+NokLVUmrHr9UJoc8eWTt+IwyU3s+wlbaSVCt3lCQtAVp/3bAYhF5AwgP87AKVu8z617vY7S
TFGcO+pCpmsavd6/gofDVR4TGZAL/zkd/Ffjt/Dc8+gq9EGNxeoD+f1u1Q5jIVhZUK8quRm4Hl9m
Bh+vs9LmPPA82LNg02oy4AijzYepgZTyAxJAbF0f2WagWaAFenYV+bZBSHh9dbV9aOeQ7JtMtvJC
9B3EHZVOyTb7Hbf39k0KAq8dT9Bm/YtTZhvq0d+DJF40U1HDJ2MV2LEKFdv8YIchxImG0tXhtaWZ
PWDtkrv/9tKINmYJ5lbiNG7hCAKmPsgkW/hTPzNKsHn0YNtMm751+JFK6AzI20ZO8Hh2wxl8a5FW
tVMS/KKjduurZFen3vlz6ta3K2WP0LBIymKQfgeqglc0FQvv32svdYBjHoMppS+lBBtXd65x6RzE
UcOr6/Atrwn5NrfcBDgnkkfKFFDSuSoyIV7XUwMhGqI3CpgBT/UdIl2eusbAe9dWKLztIEVLTP0U
rh4gkgiJTJg1yd68ejieRvR6HlFOvvPPfniUyHZoiwg+abF0h4dIVcYIutwj5W+zgCtze/KXZNh/
MHrvP4WRhXuUJ/W/cmn8b4XuZxIX2vQXua8Kf8V9Au0U6DadcMYGf+CU+c4hKtpp0W+NhR99SEK4
a57dgpvbNf7nnOPHvowX3s5bZ216bECV7fDDQ92Sdkemp/2EZBAh78OCkQ2ap8va2uG4MAdUiw/P
WgtSlVuQik4NjFQLvzLBGhNdy2Ntk4Ahug9BNhAkZCMpD+TBONAfl0aTVHr0BQiutIgI1VHRl9Ih
6nVUcuVAkqQQJmy0EPGHJ+uN9jyD9D9sp3RUFo56aqb9tTPa6JQWZpfcpwdXT9yNOovjrZUoDh4+
/pDtHg8L0NetNydRU4NgztJ1yihPX/peYKdguAlmuGhuhuU+9KpshxGwTZQCC8wBNLrinnYaHnSb
Ru6/TQoxy+OxGLSxQOBEewmcb915ki6/1Z/66QQQjwFQb6zMgh9FPd00jEIfHZnkBz2GYjLjexaO
QRiIJD5GrHrkxnEfGNCh2uG83u8LFb69ZDGfaS4kNZlX0refTXEe+AnliYGGa7feFKg8Vh3hgJiR
aDFvs2VEz3/s0WAxSCtHbAP64/c7GIm9gzN58btFZXerF9f8Zvenw62y26mbur/E9rbLHz7QtgQt
M8F++c6rg+d21CfWptnxPV3CvgL2NWXV5STF4EFZKkZ7eTjlfeWD1GEfl9uFLMPB6jTdPM99zeld
V3tyKLpwfw5h+1EDhW3+CygG/kqEPrZrquMLqGDnKTp9nZkjyVYB6RI6Bzw4J5Phm+bbKlXJBs6x
xXJyvtCVb8/nLQdKRgRfwUO8FnixtZ+eC/ZiBCqZpFukDms87guD5Z7OtnMntdaU5L0k71aHPORd
eheV7QZiHC6/a5LIgAPZAvWbQTvRzyMXHJtvQuU3t7XjUGmMDBjvxt1p8EFMI6omUxzxplXIqTOU
FJJt3qzCC8CzuXGf2IVB6GtBBvQrWVvBfOAh0hB53Uydx8YqgjkqIHHsGABk0g9BDaZpagfgdHUb
7H8ai8NY/lPJnKLdKUkZz40G+vl1i5J/3oLaesvXiEwnZLPzEzkJP52e9ig5gL/L2m8nFfJNHt0y
TpaLjpaij3ts/AY8YG88Vy/xenNxBcogcBvTNuzMSMSEEc5iXkq6acyikdOtrYk2nAeVLgLsb4IJ
W/7g+dNauwrgCYKKJey77/bAPQ56keIlemSyeJKvaaTO77lbdxTwEwmYno7jfzLjgEUg8z2gtzL5
lJmYpEKbgzMl0WpyAepX2wn/+dovbYUuFn+vk9EMTf4ZVYMqJgxeumU1nC7MxqgOkn2L5GN2/MB/
+sJF6ntVpjhSBIw6qpxqWbxaCeXrAIJfZC26Q25icTlYktFbGXMtuvgIywULkhhE5F1wunMUUGXl
inow8NIbdPKRdN/XBIqYZkSddcE0eKIztaQASpks+Wv1s+Cq38uiwqntN6tm+SrffhEK3vy7e124
ZFH42s4ZBuwpPjNuFyaenyROHePXABPQUyJgRLKwUAZiVvpwe1Bn30STeVcz1CZG1CD8lQOIjyFD
cLKfKB1p4EO9MP1kWUXEByBoA40g3RA7QmIUsjEtGnV7Nx5YnfINf1fGWKr5oBFKLAY+KT9QPKp/
i5lrTOtUzYapxcGsxF9gxxPchZQcd3lrlkOO8ZOoWJ2Zzzk9Y77phiIYHFLquqXBajwxDKZ+Dmih
mBhGVYB3UnWE5bIxsHu7YtEVvoLRFt5lPo65CToTiLQnuHdgJ3Mwh8/PMfy/ioqX2c+EhRMlJoD+
+YfwYu2pQBzVscwkhF8nUC1+nmqQpriOgFPBv1p+m5UJb36iMA1FWrsVCbGVGtZGon6TDWbvprGy
in+9R4TMI1RodvLngB80p7pzUDp6DTWlgts3PVFBqAxmWh1NhBxFGNjjRpBNluQE2GU5tp3zIw7z
mXi57CDVHMRDNDjS6DC9kG1ehuc9dPIDwKn6jf4190i9OsTdDud7thv+eNviMWbYm7mKDi9LSqwt
eSTMyZL0oveSJfRCAM9y+CuOvVVPK5hchEC0SVN6IkmkNqVwIBUm74pxmjbnBfLU1OxurNUu8BQZ
WM3HZbWhTN2BnFKJpJgHitHov+fEvt7tIrHeMdbYQ6RBimfzfuLcvCcECLYj2ejVIpjkMJ3gbSNo
bEJxXW683KkvA53T3MKTCqfvpdvHvW6CQRrqapkpN71ZurwmfmOTKNx/j/LvuNDLxalIFfhLWJOO
8bF5O8WWh9TIbhpn5N8TmyAPLObQxIgFpDhwoyZDwntpeno+GJVrZwbmdxCw+oqEbnwlcfZDzn1N
tlKdOsLwU+rFi2ihcA1UVMxgle0zI5sp8krrp8FXsv7RYfjiWDg5hrbs9i05PuBdB7OShvdy3D5h
wDufi5WGoWn3jVpALgEVrguAH0oBQ7wrRb3lj3iA0Uw0+3iSzkQqvpHGQI/2br+YrChYmf1SQcQb
O4IZ8vyN31BbBFj313v/TAKEge/SZmWvrPWIs/cTj5zRB148IrAfaiOKaEmDLXcoPlH32mQym2/B
gbhswNFJdNLqBrRxLXTvQ1ntu0z2OQ5FmjuLL9CvruFSM4h0pYtcZdwp/Otip4VNuwMZiAM8MpGp
BgZ7bOMy3GqTzxbiF77xLQxSsXt8Z+uwOr/4hND5NamBY1FfAHaCaNfDrQO9L2WgIWmu6IY79Xzd
H8Jr5+rKRrog+mT1D9H39/5hZ+z9UaE9TSJwDD7zctKAE+FdSz28NYXne9p1tgcSokeuyMVJpD0p
cgqR45Wyx4LxH6kIg45wc2Z9qSBlGEu3W+chpQDOaJHEb8ozcNvT1BG6rRAccIBdEmG27Q9ulO2y
3twp//87ty+bZXdddhssAjGnOUISLXCHAV0trzyml9cRJ5vfdjASTxa/g76TXULrNwKMBbFPB922
NVVdhWMORa8Y6u6nN7UCwoUpDKDLl173s1XKFCL8LMKmpN7ay7Kan6dLIOXo+xHVWP+dfdroa8CU
RMwESQJcb9IvHxXm/NcTIJg0d4icatVYEXs+v7DX3W4BcBEysQSW3YxYubB8RFNAsdwWT7cWIaWS
xcdAYjf6EKQOARGwmAL2QjE1PQI4VuiVzPKjTPEExcd/fg8ygW2FJWCqhGWCbkWBEJjiSI7F+GEH
EYxLtsGcA8L46TdbWsIrz13JbWiQoDYCmt3QUhRuip9Q9a9z97dikKTFmgYoECzUVZp+B253eey8
RlrqAlfA3pS+91TBxDN4ac2uH9SYkaOqVVaaZSfNAMr488OpAkg3PZavN1knl6HH7B3+aee55KCu
p3bxgFdoWpiqDRHVKJ0ngYfYqXq53/Cg1YOoKGL+iVNKyCaEkBH/otQIPC4PFvgDORXzUKvTPF/C
5eY4e5iOEZeX0G+UKI64VI4gkAu+DRqvI2KcPbR9s2s6Iumg8sDrBgfF3/O0R9fEVnoEtq9JnOQd
gfbVSBSHpXok98eFh44lq5AN07m7StVYoigiPM6Ze4h6uF+Bl2LNLf8pUl8+qE6KRGUEThAJb2fe
uYTUB0QNHRSD7yh8VihHbmBhQAkjn4hNAP8ThpBHIncrkQCNuPBE4BmnrmtD7QKZlo1Vtn/QgPSr
w2unpD9FeoBDXjAwQI5t9V6AfkqSo96+JlB7i0+LsinqlRFaKx0rNrH8gyVP3+pXFbN0zLMxGeQj
zmnegY4sz8ZyFaA/GrQQP8iNlMypiPiRCF6bSgw+RStqgWpfyA/9KuHxGuzvwcmnAd7klATVb8n5
zv5uYq7DHlbceHZkZhZUQbGOKfGbYPZLZAdmdUlSCyc36AGBwnLWMSqIuQG7tmYuTfn9UvjSnpIb
E2BBXDTmhH5H6vDR64ULxvy4CMKAxjf3183z5TYy5Eoq1+0YhFwTTVd2w44J98LPZ7wx3Yvx3NFl
puVxXZ8IWEgmoTOvYFrd0R2equzZZyB6a1pyvJ3xmskur18U8cxOZA5csGqjT6I+9g3aPyIGdgmH
p5+dkRnGUG3+vbgYjNuyb9AOSurBB+gZLkenDkfZAi7/5iNgndhXRpM7N4PC0cxakLuJobGYLpKf
JV+effsXcPRQ4mC50Cfzcm2NegO0gXmhrIIZH1c/JUAGjGf2QOby9dcUenBsM1oGOU8AMGnZgop1
AALKGZJ2nGqHXMtcDU6Dz4s7upPrkdKZrlNoL8fTkAXLjhWfHcekKS8sI8DlC/cxQzSJgyM+VYkv
NHLsuWh2PavgpWGOQSpJv0qfuB3IPlQSSe83RSu1E+TnVVtcnHWOR5Jlu+wReb+YSvSeMimpM+sI
lT95244Xlron9hC3li0vrhP+nnE8i8JCMHWRQXx9tObx1et/c7d1vSdDpB9FJjvrDK5V/d1kpH3h
S1BKyCVEXlfH4BZXVQm8r8leM7G372QxWHX8L4Te1Y4bRyTEEvXosHpLRT6HY6U7YA+7tjaWMzIl
PSO4fCZ5Le4zxYNIVS1B150EWEjECqykLRXUWb2g+dmCOBJFH0vWuTVb/Ktvr8+EXzuFAzpowO8K
XkNrEXKwbYdazhxADJbfm0YALiVocrHFvTAehXKl2lYXfOIZihwBTasfMJ0djXhwWYazuY6ffb+O
8ZVZVYyVbtLXifIFnGJlfBc5eQ+Kmr0DTIyQ4teHJ0iJcBFgp2xBvIw4V2WFtcbWALfP1rm75XcF
VIvyeYgBU3gWUnBQLQeP4G5k/rjfsGhk8T3pAz6dhtGX9queU9EreUL/uLnNXjIL1QMyin+9ULYb
pSl7j9eNBWEZJcXVg4Q5L8mf4UK/Qb+6omxB8Msan7b1KnFeRjeDKPhGvsoQgkS6Zx41PohLlTwk
asaNtzK/QyRPBW4JbWsJjV3Gzrg1IGcUvySW8wGDi6ftnXQ3AJC5rE3X0VJg1ZAEjyUJIqfK7e1H
iCl5j31gt9j5KKgU9awcH814pZGpp+j/oEJR01r6lhlvJTKuN4D0THD/hoRwLYYMkcD5JP3AsPUi
i0xJRxkDqfNkZzZwjTnTer6w2OrriFJE0FqoMHyRMpltc9Y06Ctar4ayzlbQIrg7YpdGYBqvp3zJ
MyBTpz2xBspuRztajjJmwzarL8rC4XtdaKBM0x2SuMhHekVxCPyWF42WNNB2tQBLIu2FNWHodUrz
V44j2A0jNC0g13ILdseYvTSXsUZuiaN/Ydoet7t5N47Eq/HUaPl1CZq+ACZhRXXM6Y/t5u2KwePQ
BNOyeADmqs3Wig9CvZgHjLD5qb3OgXTmp+1L4zkYlACPc6HjC093lJWOl1w0sjnx0sDMtYqPDM9M
EgOoMskHTNorg/gtUcPkr5talZLlwYrMBp7DAuRjOj8oOjOCW28vi+2lCHk4wE9LzeHAI9xOQHSM
jR+lblzvd6hmK1tQcQubi/M7FymEVm5/Gnod9QKCynOXsMHylpgVUDgPEYhOYuoLhxLu6BWOTYZy
bwfW+vhSuYdQlx2TkI3QQWJrWLq2kO/ucL+ayjpgZVj5rIvg6NgXYX9bzKlbC5deEI4Dnks83w1T
YZkyuPXgbF8TlCPWIPJU7mm7bO0mdraNvC/VRd2cZKoT+eePtGbAX6S+41EGNj4wWxrfxF4sEiMu
rmTVB5CWUgv1XDEI75q9j4LdLhq7FSVphEuoyWIn5uOcCexSNm7GckE3hLcd7EMlzlCS
`pragma protect end_protected
