// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:35:30 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
G7ozUr7uGrWStfwnm1x5+6X1AmdHB5XZn0TfZBqo05cXKP5AJvxUlg65bmC4pp6y
aWOSvxPt5dZqER+19wJswTR0mCvi4aSZ+cCjUuwu3UKbYdrxEEhBPaOc3rUInrn6
crYV7HRBUuHCySIOH57rE7WCtJOoyHZayGZLO0lCrFU=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 4816)
V0zwPnOGrLWAWO4nzzOTTxs1q8KhPU6ju02jxEqXUE6zaj3YkKP/6kY4H1VHKt0E
VzxPApcddKBs32BbJWJCsTHTpRhwEkeDTH81sk1nARXDehcoypQeXEmAL9oiWnWA
Ua7Nwfccm8J0qhPdRN1OZNDVMkKo79msEYaOBoPzW1fPg1zKHCa6AGhxtJsQ8lvF
TlhUWxA8ed6zybD/4Ch8CMwLWzXyUw5/jTaa8l8dChTVFJoljDm4NUdkMdE1JnyY
CUxThmVR7X2Cxa4J4aivyZcU5GMA4AU1VTTPYQIIzdu1Q4NBpkQPffEpIdYlAU37
0AgUCvnmpQMrBedBsag+InVngIQ7WPyNymuuao91i8RHjOARtTu8lxuWvTnw1bz8
fhpcDyBaUoY1TfzhYGdoNzxjxtHxDS6PEJzMWfXM/rPYjmoIUROVsL6vTXTNvBKX
2Md9WKy61jkVjXnseLfC+h4icb+1RJayvTA1ZBKjfZuZoJ5SwUP+TQ04Xe3vOKQo
nBKzHgWT9CWoS29ZO4nHig0i+IK7MRHkAzBMPhxs0R57js6ztLMZAXgHTNZcWeUQ
DmHIbNbWI0xPjhwxojkwvLH2amWy8xGGu7KqvYoqoy0TDkVSIk59uZygPcIWlGIH
HYUPKburaQpPK0x0Fb9mo1RKcpNn29v23cX7R3PtdJ/toJ9Uw7AWX851Z4eYE+nd
/V0Yq7JzTtlhxw8uFT+A5mbRGU52BsC0XV1rKZzHsfd1Y61PAvRSCpBoBAE/ESfc
UwVlqftbL9Pfk+iSeBgPHJ/AO5chdgeCfQ5CxhGb2lzaTxZuTB2lTvfKHRMBUoEf
vi7Yb22rQMSSFWSli7v7bfO5TlI1hG57JahaD/BUbCjt24at2kmIQyW/pqlvDAaS
Sd23+CcAxPnEoscH6IRNb2fiJUoklIPFdn0ELtDGvOqksUGjozyUV2NJGAKv+Vug
yr0lG5ypRxUil44bFwITk58XsqMKrP9Nbsp2/JBCj6Sz/vT1ROhqYsJ+bcU+dPxP
9XOa1f41qZYBxUAgk2erFIu6BZR/IHyVFLkJhqgg5stB6DqdtOzoAuXFIVjUBRLb
eBhEWnmWjh+MVje2IWtjK7z23LNttF5Q3cH0eTyuSBIw2S9UX68H5fnLTNoLFzae
9LOaly/vGg9ZXUpMp0DX/gX/b4slrZA3jnv/uc00YyHNE09YEC5wbzCa4eW70zg5
BDgKGJ24af4XUzbJtslP9PzTYaBJHyN4p1YA4HPmmc/vIrnnPQkwaMV2VFxYWe9J
GLb/rmzfEWXBijm+o3cAF6DVA+N8tEpMlAR+oIApoGmza4wW11wNVqLgnDcYZ2Y8
zhKUqMvNAm/lekXOrfvebwoNHX/jbLaEZquNHyuqdhconW84NxkgApg307dgOb25
+qbscW4rYMZnudxJO9mXqFAI6IEc6eq+uwBlewtybnZ01d5Y0cQB5jUHlbFEkVKH
0/gTKEuy6LyRE13QEEBpCQ0xoIN+1r6xlZTzsQXm8UpdmkKiFLdSATPQRc222NI8
vjSwPKBk/zMWMEt+TZ0p04cdZLBeWjyzxZY07PytKGKqFizT9nECVDIhmT5fpP3S
Sxpjsk/9Hj3m9FOojaLS/CxuhMrN9quloZouP8S1RhJ6TZziu2WNGFZPZLgDc9xB
GSTuGr8M3v0BMNKNdOz9ZX+7+t9C2WdaPQ2p9UcFnP+UeCUlKy2rAm+p8uAIP5Qw
y1QY8L0qSl4e8vjiEwd2eQKVxTeW2gXZIKuC01oClj7N8EK6dAbEuJgR9vYKV5sA
rfqs1UpxstLtze/8t+8RH/nid4dBZ1Z3oKposJASGMXH+sPUuzy8zUID368mflig
67FiSx2DlS9qJdH8HSuT3ceNQ60CMDbe5dJCkZFtZUz8Lqnhr4BexgcDNMowzr1x
dJKiYW6/vr7W8Iz8GlUkKQiB/1RkHFwSyZAKz2c85O+UMzYf45iLyO7LoeCL11yq
fl0VAgJQawbpd0m/U9i8lGh8t2IV+W1TEUyoCQy9+nChLx8JmWtpRO2sgLIlLUqF
oXQsHoVJ1Ey2YSL2QkCPMLScjvQFfgvedMSCH3icaLCz4qAP4is78c+YQep/9Evh
bOd56SHly2PBL0rOKMmZoFjsTu0TyGWbA/kKHjK8Pf1+Cn7qjl7q0Y3gVzuXyGA5
xhXAYZ485btD31UJd2nutkS1bCqjQtmqG823hyW3qjTSlT/E0gfRncXEX0XjIucw
Jed2phVNBxTPHrpusEksKU7CUBx3WGpHa/d/vhkQjDdV64zvDUHl+kaUaeWj8YQo
BiQyAuXaHNq2l87EuSROFnzzR6yaAuuJA7KrYGTp/Q+6X03ekdjuhv8jmp58Lt2l
I6GKU9l7OLXfz8qn7t73Hl3/eXxf4Q0N9P7hmN9XsBMPHOUvhbL6FqpaOf94BKIJ
SASmg9VXaDYEs70a0sHh1xtiznEhw3Ko6EXO6npO8XREmcrzEcX4yNkrbxX14pGU
P1KUJDZOHBzP6d05J0fSn9jTmd7azY1cvdVDXQFnenka9v9W9xNSCp/sejLpafIn
61FO9THLHCE3TulbZuiIp0o6EBj2pEXYp8Pb2l4FWZIhXgEgzHcL8zCCTZEy9iOb
Fo0tHk+U6kHVka+AMzu6IiPfkgyCv34h0BPvDV2btTKQMTxDw7RsytSVK87mCM+e
MEuXB+CTGQQlCkFYeMa27dYO5ahNGyhVfpU7jKYn0XoWIECqj3Jh+4BZ0gNfhePx
ZTFGH7HgNBfu6lGE3M4W1Cd2pEF5PkDdlBZv3UrpGDPz1i6YPGY0DqHkG7niroat
qjPlAgnbmz2x0swpH9xCsFvZBBNIGC5/42NolFdBWCMjiC2ZPTDeL9h44nkomjpG
SBIngvQL8k7rWK6cFxsLymhmhxqcQtwKWfT7NWsfycFOAEsGhwpZlZDqLyuTFToL
TeYLQJPUOilSrCCBu1zf3m603QvIDegEAw0Og8ZTpx82U4Y/uNxhBJ2C5wv0gjbs
Z0bLs+paCzNqMipjHyeugSf61/+qpV1SoJpGwqHPw+mbdq20oLqcH1WZo63x+VdW
cLe1onOx+NozW0ODOzDaljBRcwm7xsXNnxPhpfu7RVB5jODZDjn2DGGie59OVpIf
rMfqZkaJlj0rPyFGF+b4NznggfZVHLkqZKgDOLrltgL9fy4W09t3Rnnf3DqCRIFx
x+Q9KxBKsili0NOlL0sJInBoGuzNtZ3xtZLMppwBwWZO4i6M/8Xa+aGDXYjxeXkC
0qUWLiwb9WSiCckOoawXwwoBU5OAD4VlGOU/nS+DGQ3GDwKZT9vR4Fxy2FhS5U4o
zI8DSCbTbRgPCJw2fTfDNoaXgBfJehx4RDmHexOdrptQcIWPhmpXy6QG+1mwtNln
fnRilul+QjrNHIOTzG3guKgXQunhn03J/zdOxJ1Fe6I/X1CjvIerk+QUr5Nb09lI
2vtM/xL5ZxuTjTQ9k2cBAnTY7y9DGs+zT9sfqnxEZ26O8hsomqpxBDnf0vDuYv7u
bNq1XlO8A0mUt7WFNnC3jXXMw3rvctni7TjqeqxVt20Qtgjmp8zl5HMK/aT9AlN+
Md15JKSWPR/g1rxqYXuQs7N75+6bjU/BS1Wh40+kGL89/Y8APAyZlv0UzbnALAf/
bM6snWuKHNYk37BC3dqBu04M2SVjOdxW8fme+vZKkjvWIJQSPrY4KRiL20OrUmIz
wIwpM9CfBLoqxoacLuYrnmjoNlYxGoXw3lNEJ6tXWv7N3MFBix8AffAS81yXbPsA
aon6pchraMLlpYBIxjK6bfi87zSIGBTFEP67bDqoP7x6wQfL3L5onps9O7X5QiGv
hWxpz/fCqKICIatq+vAdE7kdnsVhc4LqBvchEorc1Xqiy6UYN9dJ115cggsLFklo
kt+bdSXJJNnWMXgC95Z9yt5lDXoOayTpLh56QH3S4MCpfkgUDTqG44KNvkxoLTln
ozLZo0LOpVpbfUjhvp1eCNUNYP+u0Aj+K3YO3uTCcWiZRSrSE/VFRZlSQXrykeGt
7A8BlqR0NN+0s4mhJaimxsr4Yh57hx+xTk450adhAAC+7+d1SHnruYS30TmKytyv
ZTlIviGiPeR2eSpaXzKFMPVRyJaSvO1ZFEHaGog9/5kDYvh+Fnmu8Wq5HMi2+pdd
F5RZEQTNIlO2HewBVmBhAcjE/vE7ijE0twPwbYH9HIAg/rq2ZKWtMh6Fd7yFz2hj
sRog2pckHTomXQjcLzAu2xC3RoKL5CZlSpGFLN9swPC54P0atAhMP0bT75ymMQw+
wCD5UTXBdt4/bcUMJRX2sSryo8UEDwySzkbaOD6LWSwLVNNqrq9jH5yfvTA/UE/2
qeO+c1ZzZS1oEheb68gauv+MAX6eNoN+1r5FGEh96DBJbiX7Z5ElAElcWics4zoz
6Or4ENlJfRu4bSv3tSdJbnSgfUPfP1dmF6Ft0ff37ibx6OGvl8gCXSmFXTJkXf/B
Xp3pKwJQA/RyyBG4f97GY68vDgEi179bKf2bV4xWS7v/q88VAgLnVZmrF4iMJo0m
mcDG5DDG4cDaANgtcDDxrjqVIT7oCusFQ7eEFTPf6NgA39iP68moF+8e6J8r6M0E
BQwGQrrQrUD5NfpP5WnYwfeFCWqy1/xkCgR4l6EsMyrHSnIR7jD8iX4GKn6QTIbc
0UZWCDxs6X7zOvHE6SvVnRCBjDgNV5hKU+U11MicZpmKU9d1PuucCxPyMCCxRFtu
E4zlW/LujkF5YPVsOtuqo9C6b9xvZs95qx43zuXifRJGkjjnKQNPfwhX2Wil2Z0Q
NvS3WDiPnRX+TmR/lJUm1GRlXSy1bRp+oe3mr/SGlCght6NtUFLD/pXhYv6xnpL7
6HlNQF0WV3GxngcrteuYwMplp59R/SLI/TLxlOMsbTXZvqg2GgaKCzCcLu7qhpr6
inePn3fhBcL445wbzai06WhA/pkrf0EMuDAaL0nzsITDCx817ewSYyYtdpOIQMRK
MiR74mL58TkYyRWxZjrnl3WL7QYogsHO+VQ7u3MLexqPeJZEnd1bVb+wQj11FXN0
kYm/3AcDmc9/MJ707jDVnR9TGtp0E+Q2Tl2SojTBofLw+WSoXKZRGoQytLOt5wXM
IdEw7uarcDowF8rXNHguUNVA92Tji+8ruRRDbr2Onm030o1YjBUjKZmGLQKOM5FS
TpJneonkPZ7ccj+ZWSPQRslhO7MDQkGgJwlCmjuUoT33xDCQebg4o3724Ey0ntL4
fCr25samwh90j4fZN2KeDYwGj3oeiB+7JJesMpyR3FxaaYY6eXGpl9kcq7ppp4Nn
kIQdv5gTfjuWEhiCp3FLzxDf0iu1XMhhYLqQCHd78NPwcRbpr6rXE1HjjqRbGSVU
Jcz8C8/PlulYDHHCBEDwX0saghNviFjl9X3JZiQGsi+u/3qxpNVmLcTY4Sii1hhr
oZ9wJL3+eWXtdrIYocu7Yu2WC077mEf4udvvL4o3UYI1w8yB0yNheqW2wp4Ieu8c
aakoyYCF3OigugStpy7ZQq+kTvmIUWclZ9NAMPfbLO4dTQrtEgp//QgIcIoar783
ZOSRncxLmOf7qBl6NVLIRU6NhtgAm/bfYbcJNdIKXTK+IZr3s20ht2nyQ+tQqCI+
8ldXeMwoTo4U6BrYkMoZkxhxdZungQtigioZoKnuiMEyMYcWaMNMLn7odOge/3Bz
dyXNBm0ukHuABCavUtChOxIGWb3Yd1qPJ4cO4M/hSLSlNxX4zAKhxjMYfiV3e91D
ibmg/4lYpH7aKSMet0EwosLbzHcWHMwIcMi6pBXsmZ4kXUf3yZXYMZpjHSBam+Ik
2H8gOVo/My8uWfY7ALxZs0tLG6yV4Sl5h8vcHyyY1B2AXNi6txjDKaMBNUoLHnSx
GU7AoJaBWGrEReoMqg37fg64FXL1FzVXt7+sc6zGJ4zEnqCydGT87Kj5AVV56T5O
x/0u7KQQGMW0d2aZrfq9st2JHOgjUB8+eoPzVubhOzph+eYpijit75wbZofgCx5f
M+GhqSXPInsvAvZgxtWAD3WxEXdYiHrMwncmgTWp38G0UKw7tdwvZY1ocuYGt2ll
+lABv89abw2CeuJz17Nk2gCQkZY8/dTld58TQXCTk0hIhfiEMuuE1CT90PWuooXY
DQ5I5E7mPZrIBWiMUX/wfIu96p3wY5ArR374Hy1rZhiJgkZhIAUi2BCgmHSJmJM/
HUw/l5OvtFHgt9qhgqrw08LPCY6udbTy4M8GGawvrjh1zuTD7y3zS0t1ZJOF4Bfm
Y5wUpjuoB5a+P6YmObifGrKAXF3d13v6svQcOLDuGq56A4ClpOfaxDxh48A9jPbx
IfZcs88WTjIi6zA7XafrCw/p6vQVBTYVY6JaA9gsQy24Qi6cqTdfx/j/nxLG7xES
wyOG6drk4it0e8Vvg4Dxrw==
`pragma protect end_protected
