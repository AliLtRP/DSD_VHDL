// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:35:41 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
AAXMUAO0fvNt2bc/di8o+LukSQYcoHiOUwjOUQU/kLfx9awYL6SDJocCC+N124XY
+l/jvCvHqfRRcXhe+1e0BdZTyvV6GlmrqbwG0jL3xgDCUSgo+P1/q49XMcqyLkxX
5CwlGa9X3yMB6Rd+t9q5dhxrjyEZw7kmulA37VJ2Ezs=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 7728)
Dge+WdEtTTEMwmuuy7hjMkdwxKqDXRlsNs5a0M6rc4IRDwnT9qaqlpTVVXSfUwat
O6LQkiyXczhbf09QlDp+5ilHbQMDBXVIXoCGfGuL7KruMgjxc2QJqYPWktohZESF
JychBWh/nOsm4hdZn/YJWIuZj2h+pyoK0UL/r0pK3fbSvHeeRtT2cTPHjAGsQcwi
jq+fMARj1JtnXgz1oOkuuvNg+3FA2oB1Inxwgt3JV0KAK8Tu/JGqGKl3M44BYZPW
g3LqJH4irP1rMo6SrlwxqNHzKBrZ0dguTU5z+jFxEvPiq0PNjwxPcGtF01cqrStw
wZazYQlfHUClvF9tPJ8SNe0c7HXjdPTlxX3JViNpftor6Abelyt+/JIcpWtmP+AD
szjl2M8c8j9HNSBHOQ+9UvGiDm2iy38FC8rxoEHrCXm/MSS2S4Ykdt09EDaHF1Lb
pMEGmM0tdS/bMm4RH3G7ycxRWVYoiTNCkRd7BRsfi3HlUxIJSYEOp8gttTB+lqr1
TuxFGykR+UBc+oks/jIRU623TrRbSAsiLs72SIW6AiAG/WpPX5hKP2Quj6KGKjEy
wPBz4/FpGAZydyZr8g1wuusIwiXLB0xqyc9+bje4nHcYOdIpiMrtIZ/YzF+mPYAG
ve7pd72DG2J7u3mVsuAfNLQBjBEQUKQ0BzhZmwwjOA2jgpBD2V3bVmItzWmV65ql
HoDOoQh8+NQlMDgVxpruJXrO4VG5xARrvB67wL5gfhfqTntrpvZZEBo4meJO4g9X
zmHifLMv98U30QoG/tEg7jSGPCXwWZlDTkonMll3dApcEaO5BwzTgnAcB24fuI1n
1nQklNNfa3emwvScHur5rmELHbxxOcLJ72jJxop4tIQ4/UndEcRZhniBvRzVO7NR
qGAnmrb1tPNaE4FOix9mpvecNaCeLQFyfKY2QfQLXD07eefLwZ+z8ZO371EhncNQ
ZRQFVQaWERK/PwuTGtFstHNvM27zLaUAEHIfiCFnaGGAQ67dAzW6zP71gAZy9L1N
KeiCEPbcD6g2mf+2GmD/ttwuwkzzleYfF9kuG5kV46zDfQXLRdcVqxtw+hUmVoef
lP9U3cpGcbgEhlyXwNTvtIoaD6yOSE9hvBnD4yAw1yyzKK1Iec3/LEQAdRN/qvA6
4d9K7ycrBLm0sPROPSUelDMExIldLQ03aCcKfEFww9EPfGSTjB+LvsE1FRjI0oua
mZ0mMqDRP8tX88SKp5zoRAvV2IB1boN38rkD35nXi7qT37DzbNK/mQJ7YQWo1IDl
VM9V5dUGeLXuaVz5pT8lIoQK52yEGVmsA7G2qlAB/OVXsPaz2gAGx17DjWc4Ltds
qlICnltuDymNUDD7twXMeyTj8Ei5swlSiMRBY/LrZMkZ85kPhFGfn8Rfd5XAcakS
9J4mYesUUGkvllfDDw3GoFTYHS7Fg28ZcWWYP3+oPzswQQvljEDS2wwVmzTjJjU2
x0Ich89jKHKAnRCsJgMWz+CqWQL/sy7o7AQWTkGKblhPPfufi8z0YNXNMMkoulaq
PU6hNG3ruPD2Y6+4HYYhP2GWVtfP3NE+elNY4qp4V1YtLcuVKT5Ju2qAVX8Wlcnq
z0/y9pl4UEPZn+4W4u8L2zC35KKFOyDBv7nstW9IBXnbCpQt4idHLfe3R4g203Ho
Z0bQOYuaBiuqBO5CwRCM8fITCzX6vLDBAw885VbFQ1gXwuyItiNsbTYdx13T72U1
BwL0jFaRCQOLtQpx/qJYYLNL2PuDkCECBPKgDtxcnDorp+DwoC9Ydx2vX8AsXWsd
xytMXooyYd2yQXtWmRjigr/tvucRC+xQimB00J9QVixE0MBkVZjsbQYluJ3vl2xg
C9FQGygz1v+87GMcrZW+dKHKBzYLVF2vcdEsFDreHFBJAXX4+mQDmoyIA5VKX9jj
SaEsRP3A3YGZ49ZJuep+6rwikxSOwOoHoj4FiLvDDPoEb86GOSnUxYH69BhaoRkj
PzBAhL6NSqwheCbL5ZHJvhmkD4K3oCXgoROTC+wukRb/FHLDoiBV3CUfC4uvHst4
No27YoZmw7VijAz8lHfM5R70rxbtIkJR+OcjC8OyDVOTZe8J8hJD/p0TjtjAB8Lq
li/x/Tl1ce7G2egbp2r5K9jmiRX/6hFe4kYT77ITs+t5KEuCHsvPc0HP7H6kQLMP
QLQk1IJ4XNIeWN27ZD0bmILxgPVDc1NxZnOhRfDXHd0Mt0sFlMEzyd6UcxvbX0fS
qC7u+osFMf8MGKbNUpqiomDdXU8jjh6aOFRZJfRPh5fqISr/Mm5sqlHy4zYVTKNz
dLTR7OgfwO9aLFXvECitXgyO6sY6+3loJiSblemrXPCYTIk+pzwSmeqOgpkzwJrt
7g+4lrXG+Tq8ybOllHKkOYpF7DB0hoMgAu2IWFa/LASomqXvzKiHyrggxC7HQyTU
EABuE4N3TOMUpOo435HPSV1n1ZkYO8vK3VLAxsgPbjqGOBiasFXP2fZLvnJXcI/l
qswdtmdAauKTiFsLfK2C1uOi1mubSi5WZKTufD1R92q7sl0PajPCyzVvuTZHo+Xt
VQ81UIiT8JxmSGpOrb0U4Kf9bIp6i37o7IipBLyN5DR5dM6u4FsqDunup1kV/l+7
whRDdiypvhaJCcwaZB3qf1SfE4KShxYxQxM9MAxc9CYj0vd2a8W3L1ebYXxwqtx4
V/G2LfvraoL/WWXf7pdPvDWaLRz0H6OEy+xjRZhspTIautt8xoAgpSJQ3zIpIhjq
LGVLEE+nGjFyD1o/6edpMC+pdBVXlJGz5HIzOwl1tskzRK+2MQB3LAkpexTgT+8m
gEy8rTxVYgUb1lyY1gkOlC1Uy/JdvFevUJkxxwopK5N98CBfZc6pu7wBltot8d18
+wvV6y2zPYt7F2JEEETqftDzEMz2o3qA4U0osBOw4+jfUIxKNv0oNfikvBET4cxf
6cn11yPrP4a9NoOs3ARsRp/Ml4OfPgxnu+nuzfTkSyHfRj89yimUMomK1ILSTh4w
XAr4CqnZ7jsFWHczowcZCT2n5mIGj1B6ICj6Ip5a/wWypSgI/ErSbgeTcvsuG9VP
LqDyDjpZQgPKzSRdlLUJnIODHpxpIr7LvBiarrVJ3ladQ1F3gc/pdl23VBMdXtp5
556TXX0MquxnHOztZV+V/0s9J/JjL2oqbZialhcJDHmUGf2B5XUZ7yWFZwIn2Mb9
2nl/A4o/el3X1mP62/YehuJlwFRg6thoq/L0pEJoRvtzXbSii7/FyXTgE0SoY1bg
5hGOeRrfNHr32pBdCSA5Dqie7mmHZSh8iaCdGVIBu8Fo3FyXlJdQ840VRF83Focy
9eF96MlptMPnt/RseCGX8wSJk2pEOUSW6NQZyGwOX7yiHJrYh7Qo79qUBhl19bfy
F36LrZKwPJW11XYfvT5gJJ3tv91WUtHrCZ4e4Q8zh63brF1xAJ1yYYRF+r4K64+I
vnLN9kYoxWQmrVGOFD7Qz1WK4uE2g90ZbKl3825+fGyDPnsLrYVIr5M/TZoBgfMu
4SfbqaSNXtjl4PP0KHmxBmAe3pUHn5B795GmacbLPrQ2W+Jg3HekZ/LqVy+5vJNm
hwpZnYfSIB2c+ogojmKuK5tlS3Y6uqj2OAyCkFExB64V6qheE65pQsP5ZwkTuj8d
dbqH5/lM2155Ar6sPEYm1tBkke0CBcbMz/tcrv+7WETV1bFzBc4ktot13uEOUQdG
N/DcJCC6dNiWnx9vA91zzp0sMZix80ZtQvH+l21cAeB8fWqGBryhHL2GHxgn1+cX
2g1DSxIVX4BmKOMLPceNBORFBrtgg4GGDG60LOYFUxWNbEMHjaAe1h82rhTqEQZR
sQ6juZP1rjLhMx6du59XJ1FtUPoanx+JELSaRGAsfKtSmmdBhf9vuaJ1bwv/HHSp
jx2OEhhD86f7j3y1lV+7wEVtnUWOib+b1rt7OisBkDXRjCdRtHFfz2KUI4dZ0iP9
kxWib+tdxsK1SEMXZWIgdF4X1pkhVl3j/2VDjA/4C/X/kzVMMIt7yVlV1oDUlOxB
0kGLNNJWvrEqtRnTd+6JLNCv/oXcrObaGXoeaydVDEzuKmHJCgVXrdfrUQyxcd2R
R1WLzvUEXLbIfploFpmMxyhSJW1qeZXkt0/Jq3gBLX6zjpIXYnrvZsOcYvG3OsVn
QLa8C26YzgktiyBj4wRhnzqJPDyCNBxqBFDWiV+ZE19Q1rRHfS8R1Cz3rnrMD9ep
vt0jAN56ezJMe0jXdWIHavH3xuC30T1YcF1qdcyNwqEBsloFewkUJDA7z1bg4vS3
ZJUEtL9OkIwDFaFWqoFqHU2Wwb99obmNQdfO/gx2EB5TlgOtzgD8v4kCUmRd4O7U
Uf4Fwob1yk1SCs8XAHMTIRJq/3eL+6OFXGF8zhTpp77iXbsE/CMRXRUKc1fT4i9s
+mk7QqWNEfg2etA8OKBazb/PifFdoI8mTY9Xjj48Cb/85X7dVaDmY/vnrRUjA6lc
0FXayXX8Nltr1LZqowgEsm9rBFUreydkwVoZYJ1qvokPyY6dts4oTeqkm/mZvdY5
/W4Ygm95yWhkPdgaP0pzYWe1v0DknQd/6AriPqvB6bxZMD3j26MBXcb2DC6fxhrI
mA5/C51dqklQmmkws1LudqRHQneaCfTMf8vBOxhDgEgBg8JHG2WaJl6LsU0Eb5Um
sKITiF85k3rDxyVKXn93xlW+rL2TfTXr3Xme27vek7E8C8NC/uOeEY5fXw57DCqC
Tdi2iP3R9/j9siDQ0351kf7DuNWfVV2UQ/UtTMQxYzgP8ig0PXxWeMCm9DTNYdEG
3KK/K7KkSq8LAqx6titwkGGU70ejhF0uzCLuvTYWNJIZtJ+HMqhdFDS7v4ADt6YS
lbN7WB2linJspDwz9eh4fhXd59bntgTQWLiSf4kGN33SrjNPmfw6j2G3vq2u24bx
EE4+N3CwFYK9fAgS84IFaIOSnO1/i5Z0ZjgEPes921pWyCqhbHV4MGN9Fy1XfWM2
PSRMrmkVcQOXWQOXNADjW+NCK8ByD6h1cZDFsEeqwZGBD9a6xVzfBAp5PriMcO8d
PhjCNVNsNPlO7D643bStUru0WK1oeIw9p8liSt8DbG/cksZWlUMMSKA79M8wM1Nd
rE5BC8ZeFb5aeh1g6ECRQU/UNjCE+HKwtupZ7M8T+76psCrZ3CbvHS0DG8c2QqTt
ACLQaeTKpY6ZtREyKWB4K2OGaqSAbt0AiikEdDNZrw9ncbvsnIDfifvqlKh/qmDT
UqRPKlvrOAx5R8uOPFXaIW3c5ZhK7HbXQ2wVO2gIWJc4R/3RZSQ8SgeFRDofVbu1
gyhBjEYL2YgtOWGDULf6cPvNKs75gAjmuRecA4lz5umJ1gqpsLi46pQ/hplVDJOn
quf5df5wS7EG7VaJTt4GOtZLuRCzv55DLR2egy2VPLIlSg0V82lmox7M2pWwnoKd
0+vNN7k8xobaoSMQhyNBu9+Gc316mlBQXwrLwpVXQKRUh6SWrDTo3JcJm8zY1Atm
vHDDOYxnz23bXgUA0Dl+7QCMLEM6Xc1l4p+M028c745w94h8xAbuqZYUGQpwSq4c
z4ESnBtyBR4nMTYnPGYp6MyAOW1hwQGYBGF1Wkf85ZYj8N9Q1jTQyZmQB0Gw5cXi
2qs2WtB0nKPO1DNs9+Tw11DtNlKEaXbysCoH+gMnvjiiCVzI/hc8j1okAhWHP3mP
kyv7SEomNczARSDJTqNDsuJCYj2/t7u4QlV0s6/u9YqY4Iz5A1xbHHxWv4X2fi1T
or+vjuU/LkxgPXxu7rJ+dHRV+d6dm5svfy47GBLDhXZ6QBGVLIvXsN2/0AbE/Vl6
YfzVEN4KPCGTAR32KiX2wo3caxzm6/pWccqwA5+UTBbPN+t+yHy12db+nOMcOurm
XpVvvgFH9NQBURYWmJrec3+E1fCFeP+3lsQnjS/6SqGdVBRFW5G53DSFG/TYRlbq
gWHsXSMCD50Ub4HClS2qTYXcRe9mRgmH5o6/fqKZN7fGRaQgCicTXX0aXgotLUWc
3iZVJw6lYhg5gl/IFXIsRfC70Jj0Dyh0dFUBAzQMR3Rs0ZNnc+Z/hk9TECcCCSJO
M832FADVEZBVKwHd/WYiWfdOv2wvMdZnwcjp7SHE9gUzj7l09xqh9aFDaEUI7eVi
p5RaX2wmkuuHZ9a6UJPp8HD1SgzQ4Iu90raExrlMu3LuzdI1ZVCRKL4++HkoqDrL
+vawaVob9pV+D+K0IQYFMahBxiPulmO5Vzfp35oNW6QtX5NAWCh8uquf/RvX1YWb
rIAKPuHfomiCDb6Z+Ca9O6/Nie7WqcbKImK5ti0l3GI9uiavIh4lRfAbjZ7RtOPy
+IOsBsitYMjzuOy9xb17+r1ZIIFrtl2sEAPwNGTfKAwQC/CmA9RaCRFAMnIUJFo8
uVrRwi95nWMMsW4pdj0byzNyS3G2oNJWvdGZJn7Br6QFYCdicponfwb4qhcSLGTd
8lYNaUjqO05RVi+SLhFR3jnOUykiIE6Ahtx3Ifq6AgOGgl3epYvq3EctJK69DDYE
G7i7FXzQ3AG4fd947vNw9A00bKFPvQTsXXo4z/GigVg2EWgRvI+QCdCk3IvjmK+Z
pFJveRSxjTa2rVFa4qFQf1mIbEfm78AGD20R0aPFM4fCUz5mXYQ38GJ9W9OPUzuM
kQQYuS1rcOOhzc9m0PhaZJA/g9dTYAE99Bs55SfKHjaiaVmD3hr3+yXyLVlJIdNr
1TR3UZ8DYV2V6o4NTUuVwvZsXphUG6WXd3oQu9HyOdtVL5gI9y6vspz9/1gCoCFL
C1uvWg6VerSa7qxBqIDa4CuKoI6HCgh8Z3+MgX2Nu3u8HdRhzs9J5Y12yLGXpSaM
3ilgxYzQYzQxqZZfxhQ0X/UgZEZOwEwNyjdnvgzUKg3jjlyo3TGD4eGeAjxmloiw
APZ5+ZPTxe2tn+ne0wBdq4V8A13Pk7hTrosRm69x3NWZtg1rxBKWetfkgrfzyvEJ
RTyC5OWh+yQWJPFw8TmWfYJ9xiQLXt9AvU8ALne6jjI1FgGj/DIqgUkzFfAPVSUP
OM57yAR75oqNipVsyaaN5pLpuuuU57sbe7VTqAkFNep7lwynF/bNoE/uUbkXxUDT
cm6BvB3ddMAdHBt//2v08+f632vSXvytNvjk8vAuSwEUiQTgebbuBU0eg/iOJKW4
EHTiw7DVokzd6+/uIXmCZOib/KBUkkS/B+kkY0jadG/apenH7VqrJ+4qF43d78ZS
DPsogZcVqIc/MU9DIrp55F7JWDr0F0xcWz7K1pL2/PD2q0joQVqLzM56a38tj1cZ
I2XH8y6ARgYvrvolylXDizG20cu/vLTLAkj4vdcGUL+XldRIiXf7wkqc5pWYyEiD
ibaXzDoykvHNx2XdVaCTnrCTyNhJMEhhZDVCvajKKcmeSyQsMiZRoanuTGmvbV9I
EcP1wX8NUwfw2GeEH6qSlWU8ZuR/EpXihiK+4TRj9WrwZA1u5QVbEoOd1JmV6RJ0
wL0f21jvIj95GNLzYOOnahAvILjkv3jWC1LFRncadrX8IyZAfMv1N08HOPI45z95
Swl1J5neGdZ4+E7MvO+7KVE7ook4S/pKyWAVKK22wCGcpDk877wpgbnrZKqT44hJ
D6z5Ceca55Xa8OawFf/6rzxoryhqu2W1jUBHnUORxG2Edk8NYFdK6uaKH30HYP32
eZHzPoMKG+n+gy3Mw+BDf/t+Lp8YQtFIoR5sJs2jIgMsWcGUl9FR6TVsQa/WW7I7
nSbT+lj0IDNTD/PJn2MMeLVRh8EwuaDy/QUWsy64KxgA7rdc1jrHF37DjVUHb0A/
4wP/ROD8CbeMbuBBbFZBXJOCvi4GsASlnMldXLmLe0rUMC0a+Q0gLTVga34tUy8D
2//cTqm3j3MKtxsitRfUFkfLgvcCrI8Vz+fditlvF58c5R94twX2VjPXOGZgoPQm
PZqBYYLQdQk62UBdYRuShYzxmi1qXiLblLSeaG72F8MZAEcP47IWn0yjC8NjMb8E
Ba68kWE5ETsL2QahlJS63RDCVexeJkqPfgSLJAP1Q/FjvIUG+dxxJAZbRVG4d4Re
6d1DMC3VsvB4dfDOdFs1GlhtnCgT2wtOjB6rBe54IBgV9iVc35JbvaeW/c+62vlq
WM/7oo07JxCL6qyLF8tuyyVwtfAADTJgM/KcAhuBiMMoqQkbNvKwPKxWUvf0X70v
w8X8NyuBH1ZcmyrlcJgRgB4XoUOK+sIf5tQOzmb8p05tYlvMiv2nhW8bREhsw5Rx
5pOQBinIRmAVAdOCBUhlZS6GubZrjh8dRDW82MCfPmA6U7s3cWs/IW+bLGqQ8EFU
AoDCyQtvNpAXWOpjdu3oUjpsfmr7S4RnA645tMvjCBKalcKVaozGkeoibXrXFgZ8
DBZ5OxtrYk3Y2r4KcB3pQzAa/DxtGNQbQlcolNt45WMDKdr2IgpBa9GDu6qHRvTS
3B6IBLapZGXt+YJxy5AIUN8LcLAwXqWCQxC/gzUXjJfc1QtB3tyYEdTVyiX5h+t/
a7fV/hKbt1S/V9ilP3aO0jrE8bJ/459B+eQDAI/jjCuCrKtNfXgDdOkPRz9pteyG
cy1t9KR8vQ2CS8f7t5emB84SUAnkDWvh58mXo+tKjP3h/ZuUnqy3fgjX+Nbnv/AE
lKwUhosGLHhtL2Xhl8c+cczIxlfydD5Qj05w6OAsthFnHRD3MnbStrt9PVC83hzn
guKPPRlpCmZi3lhrpICZ4EcX5mLmKFvjDnoqlx3FsjpJU1OufCifqNtiyCjtdZHv
G5EgU5nIevc3T/zuhyES9r8biYST8QB1IcQloH4jdW3gWJmEiB6R0VMGFXmYRCTA
gBI8lzs7fr9i5dbNk3aa6tCtptLnoXFYzYRVnoYA8vwe2YtkfKpWek9Q0Z9ejGS5
v5BnfpXIaZPkBWuijPu/TNinPqCsCgtdJGVuKXzBfjEAPx/dYDJ12AA79/qcB7BA
UvX6c19djLzYgcF8Zn7Ks7ss/yaRHW2x9ODoCw2HGLkjPEH4t8wpU4vLtZ+AiwcB
1W1fDAjRIKwxSZ9/wqE2x2egYgWc6Ig0kJ07sUJAApgnZjGaR4MKUkedWmXo+l1i
mDEPbehz06afnegi1SA8OhVyts4N4hGCeSq2Iy7SCop3nuDNjqixIzZKrHeKX6Zc
yTK1ztYRHnAmWMpOa+LMICExfoyoLp6IuULRYjt1h35elxTQdWcLiV39ScvzU8LX
1ygShzQhJNo2ZL690YdjAQU2xxF69/AEx4zG7n+9ukDmk/8iUO2UJAhZvsPgGTDZ
z6o9l6wIlbR621quIoqcnwv99izapKdF9svKtz4rzU6RPy6S4f6RnL6qGU7QY/aI
TLZRhM4lsTawYn7W2iwLWxQRcuNs8WtlPs+F7sx8d0FmlZCeI/qFxIplXGRPoWr6
Q9V1e1fFC5PIOMV0DphJCl/3b058t8zD0oAxpSU2SZbFAUfLfZ9GrpF26hDTjpCG
mtpGtMjBlBhqw9cEnQiyQ1jbVyKepkhoXLBYxok1C8iefSlTZwhg3zJ7CpxdRGXd
u0/m/kLwJZ2yRZHmqIIe2Tm7vWO5lxYMyvJGcYuvcLL5vVAGL+h/J+W/IpBUYD4U
az/hcjfoeJscxvUjv6JYhtoZGrLMvhZeWOO2qPFFRt8o+4x2PIriODN3Fasaq1AK
6MJyDV4kpf+tAUvdU5i01Rw/raR5cu1Se7wRqF4BiBb8681rTC6QSmyiooR2Alc8
7nDBOPepmU0cQzpd+VXjnSXhR8UZ92MqjG2vpMfRnJpNAh0p9KGA/A4RXn7sM02V
fSK1Qea8+IPu7yQGTVYO3P03QkhCIzFoxpI2nXeHhIwI6xmoCRcjzoGC5vTO+C8A
DXt6KpEoJuIt83WDIEd6SL+nq6JJv3qBqQSOzMFOra++B5X2VLgAkdhMi7ZgmkJG
yLX86plUd27JTTeYoEO+biXd1uIhi0oR5/PmvARZQjq+XNwI3wXw3w/HPSXysCZB
PnrZQ3kSh5L05mO5DBDOCK+faToRNFaqdBXPQWHMIeg3Ej1p3wqxWYsn7VMsD/Mz
WSU/lDmSrmGO91jJNCPru9pTicJTOHQT/2oHmQ6gyEeFzv7KZyM0WCKcH8Tq+hMl
SRCi8Ww8dbDY6xi6Reyb6en58qacTIMZ3BWqIjhVa0R3NOYrS9ohbQf03oKVRxwh
SECs+BP3Bp2E74yne00sqOEX4bvfGddKXRQPXp6W7YyydcmyvTs9XKZf5Q4IRSdS
qchzcgDcT6qUMxp1dFYaHMgOVicgYl5dmJ//bMlb6NkhDKEdTaMSoTLCxJQYulyZ
`pragma protect end_protected
