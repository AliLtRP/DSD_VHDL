// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:33:33 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
tA+LQQIP00Oznwda4q+T5QQIxb8FTudHrHvjhnXYZUUaZPA0HbbkpjpcFvOCiEbR
BFsvSeyePmyTgu6j6kQU7MkPY6cR+WaZCax1Eg3wnYKDWSL/j3ILmvPEiFaGa2YS
HVYGQBi3psxoheMq+ybGxfluvXwFrEqTu9UScNKxCbM=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 29344)
tL8Ph+J9EbijGLVjnvSTRXR9zfyI/dQ1VW6woEQhFDSz0CYdBbfwLPDpemfpNvAK
FELxq7VxwUAZMnqvlptBMZ7LYAsMwWoV8Uu4TCgupVzmo7xTNlSOhd/V3eSq6ylr
gkUV1IODO3AH35+0Wgh2UdOdmYwj2msoaFBS/FgtiOGgnKMvpiVSO22fQ/sipiCU
XN0wfnsVExy4gnhy7jwrILlQf8IfTpQOmnuXEWiuofZ8G1tUksQ/u+oWu8MiieOL
9dIH7ooaPZqk3nW6YlDY3vBFU4K9CYyfDMfwq26uDVgpCbUBEGGDx6VEvMnnMZNA
Ht7K4hr2uwwnC2pEHJn4k4f+APu0h3Lu+dqo0EelHv1lgZqFzXzWCau9Ml4orQV7
u7/0tOd1GZ1le+1KBEV7fN6noRom+7Ylb6iBgEqEz2mzWiQmPqn7M3Ily/vnSrJY
uNcFfhiAC/qAppl8eZ6Y8bMpVOftjRzU0aRBEty0sLfuZ9pBebSEQENY0893BU8l
VAwC5OWIwRQOKDbLwbExqzoxeY1b+5Ub7nvFWrYSyHnEEVwOgikBlzdT8ruhno8r
bAWv7S/TL1W7lHY9bU8Cpw79qwcuNDVie7I7UMc8IKCJjeRuRWq23zSyYWU8ow28
tC4BVY+tjtTa1HGfQW0c9yIwqZgNShQFLZdBbKlUSVH19QuPdlagnPEthpNurvCH
A/S6pg+2RLKkW6dPCasIlRrltJHyy0rmnf5kHujFf9s/vchtjLYVENtZwVoSwc5L
mADG/L4we4V9iQ422Ra4+xTRZePWE1gH0N+crEUGaTmoP8DXk7pNib7sFYKqgBTp
49lRPOJUiBfiwGG6tqYoIPe2HWwaB8cbuBJ+Q6ryzAJlFlc14xk53Y3JuiEa5zrc
NK9QjFf7jWEIzvi3csAfWkvJTZNvnjbPnpi/eUaazCvVApHSmXVUcTb4GPeRJGgQ
9MrJ0u7QCSctNAjz38a8tEEK0CAdTEo5eGZ094mvMBiX0ylRzK+zzrDqDj/arLQT
SvBOQH9QKt0S9xO2+DlofPhsAAYxjkM2KrkpmSgFo4BJMIlQk6sZct3ZmeNOQnCD
shIiINE74FwxGnkWiHl0Fv1v+8rlwXamo4db9LG3hrqG6pH8wg2mWeZKBMxm7peR
ZOSLSR4zbx+/v/UQkSuAwiCTte/UZz1vppC2Z/qQrz5Qp9orRKqKbtuaMGK2gl0E
sQDinwTzW0L4fyfAWeHbmVciTovNq+ALMd9/j3dZNn3fIQfAw3vteSkcNtEiJGfu
62lzZOLFG+MaVlmnBMZ0xOfkFifLDRztL4ibpDOy61GzfTZEDmwvkYbuyk5u4YSt
dnzozjv7SDpWSPNt9InzaDIeqTRm20Z+lUgxmffT45NahLI/KSp4vDbCCUrdv543
1nK7fI6zYAxP8h3H2jDkHsEkEMXbgSRZXG+qm7sja8wmp8bvTsEQUx1e9yQuAAz+
peaTp6RnISJuFgIQDja5HiPnaVI5yFnzYm7M5oW5pOFBZ3wJ94suRB2BCw3oIt6F
n1OS4QhWCQN3cYI7EzWmKGZZ/zKA1ohIk4EROEAK8I16zWfxCCMG3NUUi22QB75Z
+YVumI8xbaG5oAG+VEYNifysqwbyCGPgGOpIFUIngve2oYDq79AzQKperiVXUlvp
E9nmRtJtek07MDBbXZOSdDNOGPe/izJdwpyCz/s/6lAlhIcJC97OuO1p5HA7skR4
1rXH4REbyVImBIjTP4e8Mk3ujKmaLHppw7PiPzQCHlkFj/BLiaTQkxDa/p/4XDgJ
P9LxNnsBYqaoqB7HgfooPr0D9iGutFfB4CtBms2Qz6QNonWmjejPDUH0BEocAdHQ
F2uN3eW0qURO58ytP2b8gQVXOGnQw9ZM2+giF3LtyLx3p2YHgsTcDlkB4HhX6YNf
rIZYiVucxtLlXDTtMd/qidopvdNyM3uMPJmDjuPQIj2XwBBAkcw4VGgMtZDjJp0g
MjXPqik2ImseWqmNlZks2o4Qvk5SMhj54bGA0B3U4KHuc+nGytVDLfnLXQzkEONk
gUTLDp8bqVMIG7k1INUvLifBBN+pONrePwONFscKR+MxMBgXzn42yX7LT8G9Uzz0
9KH4TpRUfuaKVVBMaEmb+kv/jEfTQXo3EHth1QCMr33WqtDOuniMU2/oB8bkGHsT
R5ZYBTZENCPLh4W+eGyYUlkM4sET3GSqCG9Q6goSSlvLAsuD5InxRaJ2MqtFN+cx
TQoYx0S28mYMtQYdRsLlnQfOv93pFsT+BAqBPv/IHK9K09IIogDuGUNKim5KJMxG
l7IF35LlCcFV97n4ARHtnQWLtmfVtQAbnSQEbTkxhSH2XAnt7kfSgGwpBpouffHk
J0TwpeXS5Y6325vEKNHyfSIKhg/PbZg8+cKY8XfdDj6ohNCMko5jj8oJrzh/V2fn
mODkAeq4keGDHuDqF1j0wfr+/kOOu3mn0BBXarJsmIiWizLuxYP/qRiZdAFCbqP7
AD+u3Xd2/Wpn1d4lhbJwmd8gmd1XbPiEC/pG9AS3/a9xnMl8a92zTDv9qSjGIIaQ
cOh5d5MJ7xIY1bNLBJqWZ3t4MnIPf7k9uvtNJd3pQzBVsJPT3KPIZ7pEIS0vq2Cy
ZXvjtSsHg4ArmN8qhHoozgXplQ2UqnR55VGiMvs9wU/EH9i6BT15je6/yFBsldiI
bcF7dADGb+B5XBS17riWnGZuFDq5fK/f/jw4lP1Q1MDZLSDz5uFTkZB1uvqVAXu/
TvNyb9PTzUUthoBpV/Sb2OdHhpHN+gZnuSOCXvc/lICxUS8/lACOGVPMeq0tO5Ih
3N2V5sxe+6jJAAd+8IQcAKrL8/hvtA39iqD4c3/PTJLEfyLX8A/f8oYu9MXemEnx
VDTh8xiOpxqJCJhlure7Hd3GNeUW/7+cWiV+KIo4rQ6zDh+zeLn1inrdpmlOUprK
gJ+c3gBsST+VIKdnoPi7caRFjEZl2TWnXBI/RLviT+sw6cKcVQZaOzRCAzJShb7K
dGN7DEN8epD/EstUMGnZrOH7AFzjbERTW17LHFMTAACn9fnEQBIno/zKJ3kss3Kv
/YEwJkOPkUaojqM9qrSFh3R+5bgYw/feJPB34XhihmafYRHX0psOPbVi+ZM+ktp1
UMX6IyCmvOtErXho89tudNrePZxjiYp2/JGkPgG29quEEf8eTFwboU6INp7u8Oqd
ccHCjDlX+GP0ZqRSYwchWFM+YgD0S/zy7E+cEeFpNPWwvoRmJOy8Jxi7z1+rCvs9
g/ygI/E3angTbZvCd0HmqZFwr9iRhB3uFhwNf7ansSj/Q0ffMSzrWJP+8ydzhgas
H08pwvxKICMxm9nbVCIOaqBCxbG5NdeLZ/8Dg/3szTiwY5MVgtM1/fv51+P+kRn/
IAzbkl2gjoAKDRQP3wjiIIzcxN1+7Spd7bStY8Bq5RCT7nL12x4ROZ/ekrwsKiLd
+Wn1AxrPpSWtIeRflxsbSdMLfPuTsHXcDsJTpzPX35EiZBdayiBeHoeXdJ3EFWUx
7IqEBWY7ArzNfS7uMgzQjsR3WPT7BMPa4WIy4Qte5Wgmaj5Q0iDLiu5Luq0X0l5G
r/9N7e79qLvrvowRewOUGZRLJoErpwVd8Tc4VwnCdSMnVfc4gfMVA8FdI5WexCeu
8IC59IBF7byGhZ6e7ei0mNFmzqNxSYA3c/OPk/QTj+YzcalTE83u6OL6vqhcmm/1
yFoNKoE05L1+JOYgVsLi68tnXuPBslGJwjui1WyuFEqfKUEHb50lXQboD0vB6mka
wH5erT8qWGsGCn99jYxcUtzEjM47LoRnhQWLl4/kDSw3gFBJVEn9oCZzE7TQXjMW
b1T2KSimXXpX3Miu0Ys8ARWER/Z4QLDKqT8dOTD5Af82RBJfe5Ey8/ccq0dH0Wku
R48Hfq4HWePb53wODSkKNqq79mQoa7HDHfjmfw08YCBr0JmacihURp1ijUpExJ7k
Bp1NzA1ISU/rg/sXoddnsSSutoQKP6PQ9RPeMimmz/5Amj9tbVebcdJMqZDOb3QU
sHxUdzxwFWga0vYGSt4UI9GKh9Jfc4ger29DgodleV9p/J7wcodSgRlU2ySLplxo
BBfAuOxSYfRWEPU90lAQu5pjm8SKttP4ZRWXVNta8J6VqkN8ua7DmqZlvqi0Vu//
DtSA9GQUiqC9017v9kOPkI6lC+XV6LWlMruRBovF8k1OQuhRrI3qbpbdZ0KYyBiL
uihAoZ6LhBqTryzsQ6+7ubIa521bRa0fXijRaHQEbebJO7h65mV34t29/KmTjl1h
F+mEtz/4qkkQyW8RqFxcsbH8/cChjCBLKCCvEZZMsRQ73vEFYlcdgHxqxo9YIQuX
ol4yqOkkBjd9qqi5ubUSoWXkM0VaFPPoWm4fB+K8V7F8I94tc84cZ9AQvCTfuqeX
tu7yu7T/DNaCGmF8BkjpXQtp5Ymd2+/Sj8DhWcnKntb/BZlNplNxDw1hDUKk2gyn
8GG0Tm2meOR+138UsXyatPBfdFyVEQXCddcKaQhvio3t3spS18awKN8aSLPNKoOZ
I08oUKfrT16ztRV5lPblkWQYBeyZOZhj3oaAkNLOc+5VW3cR+rzD34dAvF88vuYr
SsndD7rZ8HQrlTAntzrRBWuMSUwAFyA3ts96HWiivAW13G7pM0bck2y89hHAbU0c
0EE9vkbbakdFyx6QYCG/77RyAQXdAkbytIfoG/4bTzPMFabvQ75ZyyHIY4c3Nut4
de4gPwdHz0kwdlDjc8ipniM/q9uUE87yNfZBSDpMABcVC3Akk9CamyDF/rTWiBoS
DhQDjADBfM9E51Uwo9Fy/HujGoz3scQSw4bIgPHjxyMJgQE6KbLRO02UZoVUkDiJ
oMN4Y8kWS1W3IqZ++w21qDGyELKYGkj1AUtTMNMHbusLYBoYWBg7dqiMW5dLdDGS
XPYZu6RJ1D/zv7mpP0Fdl5yBcwv3nhoQO14ZIWqzpjiBOYIxxL8vugH49JmjF5dA
V7G1lnKsazlEZUMMKkp84UPC/GIq7M6QhG568SQnG32PfBHCXO0GtVZ7+IUcnP7x
En9UG4AqT6JO46FijlEIS8liH+cMW5rCYhOPoiXb0tzcBRDfcZo1otvkjp3xR8sE
ocoYtD4Xs5Wt2HKS89tEQLlrv+gdLZoEUiE5/ioVCp4FoxrxpwN0TFGa6GMfmCug
05vWHRBQHN0QsL7MqhjP+GrqswxJRJpyvMJXJDPTb0JXXjpyRTiblOuSCRGPnbVD
IMzDLvgEtBi/vMdxaCMhihVhbXrFUrlH7gZKt2rXcya0an6N352ZR6ix2vhcrxbq
NQ2fSsAN9il0vEhYj8Nm9uvgkLyH7h0DFZdTvklwm2yr7AKNBuLjtOaEKHq5mbEW
76etnbsY1dVxse4wuFrQuqZveJTnTaR/EfVlevW0nC+q9x5SFWnE3yeBNbr4H1Xg
rzh51jjf1MbGko7BivB/4HRUFyoL8ZG2W+gCjvXvWHn8FLnMu/fuH4HNIjtAzotf
xxCfbo4XS1jv2pOwzUhlVsWrRn2wMabltMGqoToqFe4xfw/mdccBGOFrVcsE0n5h
yMXg0TUJDvodYoLEMQWWW+7PeifNGwEN69E3Z/LR0+tviv+zkBu+conWN6gZn76Q
dRKkOTdKZFQJsl80IBllN98RCtPPwTQI7p+nrqLaOyFoy1eQlxhlt/5xBsVQL0/C
IPEqSrUjU2mO3OgcFu5Hm870/clH0MgQZ9zIS+2fuxvwNQbb9WsrOK0LGv1va3kv
Uk61B18G0PECsJ0kKUZYqtIfac29hmKGFbp423Lc/NxIKbaANwm39ULAirl5QJ3C
AK/Dasyyf/Ydi5DGLjbNIL52rICoJuRuoHJGCK5TXN8oDuZQuXeYnxMvIU7eylEo
708mZ0XQrEtTRd2NFcwrac5FgUAjJicm/CNacLdAoqkowndZ6Rl/YL2UvfUnmF2H
lPzIOV2TJlPhdrODHkNvt5JGiw2HQaCZ9JxbFZrsLFf3M8YjoJDc3JoEFzK3wHsf
L2sEecTqpUfgzeNujXHXL0mQBEZ3i0ryWieb7cCpZkV+sMHm+N8RVwF9l/5d4WB4
Jd1/QisclVTINKezJ4dwyZQLul4Ow82+EYiT0JZKtHIwdFYV0mR6mr8619v19+an
4urIVnNC9SjIgTzI34TVy9M506Rhy8z22puFCzDUOXHw6Iu4YQhbqKPDlyf9SYTX
sO+F8ztuVm7DYNeiM0DZEzgNnu66kGqp5mcS0PY80+OeyeW572dOZ2drSp13i/1n
BItJ6KCBtSMqCF5ON8AiqOMp9rv0wJddmwncdHmCMjT03ExtYY0KoG9MA42IMvH7
iA4Neb0aZ65ZaperH//98AHiC/TVcOC8ZDDwLACD6gEvB4lV0DMi1Tk9qzT5QMVb
jdbyv013OiVfXl6tQsCz+r9nhqH99TeaRa8gVcn6EPoKZdmShL8iJ/j5VbYHGnnk
JYW0Cp4n5jSW205hMqCpFckanUZfXZpAuAiPm8crWGfZYzXwxPxBBWMkyDgbyzsu
plpY5UCWLNiqVLRFnR6WSP7x5/6akJJ/KelOlIt1lJHj+VxzGeA86Fn+7QLe1e6P
NiJvhqJSMS0MjWnSNemXCLgbawfx0pewxcQcjjX0WG8EAB1rKsBar1Yl0rkDqN71
1Jx+8oNtJVgv1LbEwdSHLEq/1Mi3JQsrzzMw9qTELw0AwPAz4yK09sybVigeBNfW
H3XqbamLEJtFoxTPPqIYLe4LzBOA205qReNOaaa6uZFJXsDEbc/hqfj/dKvLGdrb
VkZ3mLnb4cn/lEkjlV44cBYpoLk7dZ/DzWfMi7fyCq4ISDW+vBbUZrYFoau/wcKZ
i3Wvrh0wOTFz6OOk+ZcIivImqU1sd8aGBhs0xY0VTb3uPgJY3tMGOnYBdJ3QgN/h
LU84QfSYZ/5ZI3AvEs404B6a2RZOTJ7T1YL7HGBmN8TcriOfHMm0Z0iIZKQfY6Sp
qTS0LUfiWffihSUHZmXCBC8KMCn+znrQFP7wyuxvom/3Cc6sQ2ZpPHJjuPMFrJiF
wnP8LNzMFvnoTAS74mIiYI5ZOggB61bUzBqdjKOep3TB6AyINQMsH2Udywgbrz1B
fxpWm7tXAk27I55aR8d2K2ft1ACt3mF8wuA+A3PGps8Ci7Llp53qzxFpouHj+lqG
FOv/tSYs4NII9UkqQooCTzxXMGtOLvC4CrqLmxhDqU3U8f2i4mMqS1rR36tS/UH8
//syg1h/4fIJOoOkmCJZRRQBnHTVv5JhA5Z6tUPGHCmLY3d9eMGyQiYpZX5gxNRx
r4lF13+cRurty/jKtgrSyzBManmfpRm66ksmPHbaydIyNBOqCEUFiw+6f9UZLKkM
IG0NESl0/9iKWFAeBdEWKYSz2CV9YjEUV1WxD1wRAEKqmTVXsuemPEDPsxmzbdSO
K1NRUct4XPTGCgyI76vzq2zV2IaOpFhuPyWw27MbW/unvQ5bhmgYU1q07PUL0c38
vPUdSS94nPqUahf5DaKPVuSc5N5F9e4sxyoOB1AYjelO2yJYyWlRZFvEMcEj8wYP
KpmtvR2/e8eNx9W6DDDjrTRJMPaWnkaK2v6ZkNosjSSzlMdEgfJ6wccmLR97NsOf
9/4XhqRTrA9TB3ydNZhIF2VEoSweOKc3Wg6c1Td2k4y2av4vD/WLA0y4QLwQq8W6
76Dz65Six+Vah8iDvWtZYgom1DTfYy0p6ZjFEiZEjbS95gyQl8bTAc+Ijwc19KhY
kQUk2YMXUXt/100ow/t/EaQyt6jyNgxkd8IWumkAG4XHoPytGXpRidHkvTFdyW+T
pVe5XMzkyUmURQ/ZB9lHw6gHaBMssy6huNmv4dPzGTrK3F4D1PCmt3oIMnLn6ojR
fjEtBD/W00vulFutWNZza1TY1jPZWioySQKb4w4GzK5Z3vFM9bUhyGInaPm02T0Z
2mzgE39IPAKQNl/RxgDml6fIirwTm2ilBRzjG+cxiklKFuHwr/6fSPHr4o28YrWq
CIyq6Rm4EqD6ibHxbYSV8cbw6cQyEw1mjj+9h0YkuXQlc1QQy7apDJb/JEAOfE2k
xfeHPiMVgLuptb7uJWas6u0dfyEPCrPo9H/QhHkkPQS/hOQznZ1dsb251a30AhHR
NzTQdO6h2bO0SKAUjmnl93enbTHkpB4YlTs3+H7rA7F6GAs74SOjpumWTEBXA/45
CzVCqbM70khPEdXQxKVfbMu0QrHxhYVz/fjLDvDbbw9Otvzbiezo2MB91i6bJySG
+uu835H7T1Z30nN52sXvQJK129pWx8/Q7MCeV64Y7EmcV4MhFkXovgm0JII/J0J3
QMrvqyjXUYibGuCATnmCLxDwhZhnO6zqmw4qXS8HkEnyQc+vttR5GZG2txdzjQo2
CPzWGpG/Zd0iudtBuKKa1y7ihyRZH72Q5bZoW6iEgjwtiyNKe9H0JfRtxtXNocLY
TTkBrJweOPuMhQ8cfFn3jiGw9pVQTcBfiWDTvaZIcSdZtlSXLgCeDJNYM2fc3GtM
1piTWgQjtS6o/cVCuJu9JB+3tR3Q6br9YMgzNePMN2n78MsB+bUcpDQF9aISpauv
AZiGIgakDKPidnmV8lwncHq8g4b+A+QljsvZmjomgJ7K0UX4hkS2gxIshuOpZbAE
2nw6wBQrfPBsZTL3AblJhKMGdslACjn9St3jtRys4YTmpiH0mTaVpsvJ817dHt56
lrDfZBBHoqMLw0/OXamxz+8oSqjoecsun+u376vuvpDzHCp8nkN4y+akWChqUslt
iwLINFEYq6zK9rVsRLWjibaXaspGu7VY+nS7aUcLuHHw8kGW7PxPEtEo4JLQVM4L
C/ZxSNWT/hC10LMgbXOVLxHcplKt5EDUOfcf+wsw5I/4AEEB6eVb0RiaqQAK7kXp
nwLPWUkJYDYVB/D6H24/t9tcVCyf6BdLiC6RhHsZllIa5OhO4Mv//1ZgmbjzeRnJ
8CwiIbkHVLdnkNnRZKCDned736O97d+8ibAWK7Rty/SvVOqVVnkIud85WQAUT0Pn
muhbTj160ch01hPv4d8AxhGPMY1URrtk7EdfynOErQgosDTHyRJ4fUpSdfmrCufx
ABVf01GbJMAuu9R9wF0LjCRaQJsiq0kHJHt8QZ4S5yzC7fCFwIQliWdhnZ0NuVPM
lSQdBx8U7ezEFwoMIAtw75Hfa4241zrvoB5kolo0jsU8mPAzvnhjjsxVlKcE7ghC
umIqLUA50k3EAyveCRM36yoc0JmIC9A/EW23+KyZwlt+p3wVpCsaN4PZykHHF3OD
3oLkpwZiDIrzMglvNDdQEzILREZckagLUYiNJdC6M6Ol9XYvA5yvQJEq+6Ss/FUZ
os0j2XW0/y5AtsUCmSCCCwVpSL85oQ7E4PfdK0IWbzjwz7lsNOA7bx6WO/d+G41W
K2MMAybD0mCtYDXLaDdUGdEn4c+sDRRQxlkwsqsnIpexjaJeU2wbbDaDjqvW6+Hl
DP8pOfPm8x2bw0Aqfo6b75CFc1D2TnovQwyj+pUsZNs1JsXpDApPZklJUwRMXZIn
3+EA+INT1ZR8rRBvrdeYqDSezsLqcT6dVGEP+3uwjZmclq4L4QUNNP4GNp6XruLU
TUqdwgXRm05LVkmhnvMpKUjjE2lmd0ZAnmT14b+1k11txUyauJOxQ/UHdkuS6OcX
LT8PvPmKvRvJVKzsvMFQkagD84e3uFappSnhu/BLPivsz0rro7+tkICXvCt+VgAV
aSwk2Yw/sceQVkFOThoWNTaxWVM23ynfgzbGBKzPDLjAUVdDDZKQhIRiOSmSzSjy
yQHjhvpjvnY4aEXJvfLPS0WggVclzCPZAlUyOPifvYIEjdJGx/el6puj3MdmCXm4
P1B4oC5b7q4vgnLZZRfW31T584p2hxbVbX77pORPw2ZPhje3cuZgEf++RX6veFgR
wNKPFOt7BTJKgsiBTMujMxl2nbRctBYrgeGWWtx5dkBRPFPEtbMzsQcxxoa74ASR
AQIe0cyt/2ACYTY8TVDGh/BvPXYPLo95ZWx8x8M3UfrgPE/Ozu3li3UqX8vlZMdf
fecM88Vr6WKXhu5hffa5gwrzYl92c2eP3lwxfSOdm7ZIBlygTcVNOXOoFpfU+ufQ
qyr4btqKvoODfhZ1rm0i5FGTJnxhmodtIdi595Z5TFVskwE5eTj+3q/h0QIAisSH
TATbBKsJjYrCrvCOeohAIE5yZS0qvUH8K2tpbcKXtRUP6uK3pC+Y5QWKo288hlom
jQiLZ8wfSghNW8ET4M7kox6GrQDaOloZOCj0gItf9voBjhyu0D7/+tuRGy8wFlb4
8xksFYc7wlZ4RnMgtJWJXFskHZ21LJcHy2RrLTWlbfZ8RN7xAO4q/7Iyjmoj03Uz
gTHc5Xa8FlmzXrSIMepZRtab9Qxfil6a876m+yzv0ONQVk2d78nsVufRxGIzPWbN
XLB7BnjE6OdvLv6NcTXFcLShMze3fQj49PgwmOyrR3lg/AC+8OdnD9SynEejRmGx
gZt5q7eKVIvim0PB2mJkknMIKxMe8p6/i4LQk7OSsgduOxUNIs5LpWhSsV47xzvx
Ru0l31Ch38TU2UaJ2CKRi8pyExT6aeEsfEWcwG+vY4eEDaPMlnhUIICuHgIDllQG
9lUuks4fqhijiyCdBvUwZnVNOh2G0bVcGe+K0L2Z4KZXuFZcnI16rKMIDZY+r7Tv
rTLMww1dv0u39HXndbhbBOVqJe/D9QXmtp23jNGVZxSmLwBs6X1NgK+Iwi2Kqcvd
8EeCnSs4Apv/N9/EKpNh5Q/TEy/ClVakBATa7bhSsjpQku9hBhSv+oEKZI64rgoJ
yyiPjmVmBK8SLcnmc2J+WrPHS7Kd6AjOeueAIbeS2XhBn2s6522DUb9ub9rZO65K
Gftsnth0RU7ZCAMtpOUC1gtUKhNh4lGeZx3UFtp47T2iwOywOXJRhIA7kMo9xQ9C
tfON3/JoAoFaEfQNCYS57oSdz9hEflogKQgIkCKx/K0+pYS8JV8eEm+8uw/Ci96w
ljELlvAkOFHldiRAG53qEu+r774DlSxGOKJo/lD03N1WPl+cW8NF+scQyGadJFSf
TQp8IwWhAOqIAkgE4XK+k+A09KwN6QV4GKFLL30kZwgBS1Nx2ERrgWukwY01DhOP
RH3lLC5kdxbtdchLl5aM32B/gVA65oj4JQ+sf7GLIXpkNsf9xJfGx1aJ9z0Ji1mj
Fju9mgLurrdHQrFhDKHXISpwS9/W/4oloBbQUtK/H7ZW1Bj8+FQIdw6p559+s2OW
Bq6YJUdTE4iJikEAGU/lpoQisci3CqEwbAWE84wYuAdV7hbGQ1VPZKRRj8k5N8tI
mnDnYCEJ3KAQ5eQYzJ4XijodU0oq5W16ndT6s6r5WJwI40X4W5q6YncmHVAuuGSi
rKAwJQuWjmdctLtLoRiFihsColNU8X6MFZzj57tJEhmb9pZ2Wk85z23hTSH25BZl
vJTOlYkv0SkT66rUoW+KtkLQLERpE1jepbfxMUgbn75m/XKTAvrZ/cRirGrTRNlN
KIYG1BH/xTKum5A52ErxSOBnzk5pxkaldKTqWaF/NcRlUz8oJM9p/Eff5gi6KnSU
+q1kh29CULXf/hGhbqt5Wxj9nQog1htdiStgys3GkBiYT3hFlge6fljvaiMZdHwv
HVtVpYq+fj/JBs2rJDMnl3C2MC3qqKGObyOtE37y2HxAmE+p4htTE+F63d8a//OD
S8ZWcyyJgHwWJLF0FTkJegiP1xVRvxMFbjEOkOjqBN9fR24z6h/r3npFRIEb6w3x
2Bi2qSyWD66IZcS6qQ2rPJwxLs+hcpBu9rv3Sc7jJL/wjqAO6czxpHWAN9N/RYoT
UaYen1RGMDrwj0jErjaej2nsLzXUWIL+KfQffoYzaAPQRKfifeHCtFQAW4VS7J8F
nZkLiGR+nwZ5wut3+vu2iru3+Bw2O/+3+VijXgND7MJjIDkDZ+B9j16gcMpmoPZS
CqmKfiIFHjVhqQoY8UmUR5ZmTL9GjsObwnWGfImre5KpDU92QYY57pjJMCpIV5Gx
R/5xZEThlFaFwtZEJDsQiLJXVbjGGj3J0GXpsaK/UWT8q5getyOJJxUtQypfFZQg
YCs4CLF6W0PSKpejIyw9/vN2WmXI4lSnt4nd68nA4XY7FjqXMC/kZZa9yn/OUfFR
wKcoyWrCzaLsVWEc0invwE8gQd6osv8W/vQ+HnRSN12sCa5dyUAgCtd14bAGaxns
/aZ4MEAhIMD7863Pu+32DTgo4Y4kNLBwliY0imBMmtZE9JhrUbecav25Rxg+x9QO
hFmUlyv4kFr1JZAGkuMg1dPzsc8hLfhRvBjnQR5liuWH6Gx10FQklhQpIJW//yoW
tAA8U2EmRHtTylLA/5SmEvvnxoyHUZxoDtPU8porubfDhta6E8L3NVw5vWCW7JyD
tWLg2uKfmJGwVCmgKDjKqsReb1KkJbpKdNbKGGYqHvhwSCiaY1dob8lKAYulBeho
aU5CW8CTacteFPcSfq3zl6qUDvLMHJIHIqO38ePnN4fbDgh5K9tgnC/kxkEiApN1
8p1wwI17nz1hkZJpx+Q7rRLEhqTuXruPqYLZd3D8DBl7+vcGloGib58g6ySNI26j
v4VUWolb/IZut4NCZb/V729MZvdF91jb2WRooMLFuGWkiYW0wTtHYVoYgzbPA7rB
C61Fr8AtWakIm5j8jm7WQ5uQtCiyYj+8VyFOGQotUNDYG3fnwgD1FnC1MkHKjVMK
WtPKphD9UDshz1fDzbWlzLtiC9aFGWT19KE28cQ5Te2pfQ7cDCqssYNrZJnlumph
wcMJYH4VACOh6yVhpHqBCSY1ZTQ+X7BX7QszsJn5ND5/fsNxOewi5U25HuFCtvhY
yBwc43/3a2R3jB8ldBInpPgeaVvqj33xPIkCt9EC8LShVTVS9OieiQ9S/2WZGtJq
qc9ll7zrSE8IcfB/qH5w+D1oqqE9yIserXQaTDQ9qnxQ7rPVQDUQ5+pTEygNiJuu
6Aelv0EVd3bxzknVw2wzgiE1pWie1ZK06fZFExQ86Ia5dJp/NpNONBWUUXqAc38F
lDv2K+P52+P8t0tpL/0Dd0+epuUEZD45hujXuSKZnYmZV+q2eM/M97qU2hDxj8oM
hwUA0qmCneRLjkStGIpPX9w2C4IptJG4bl5XamIxK5JfKx4zfHM7LZqq/4QU5jL1
geIXLvvTDjCN3vIf7Zoc+uQ0f3V66wmVgr25IwMX4Sj5UlBRR6o1ML2VmpvvFHIW
AOn638kDf3xw1S66FZUCsObRO8EwdPUpwAWKZTFSs+mdsOXGBWqGM3V+nbwOBRyh
E3hmvpUqCnbYl9WYc3F/nr8zm2lSXGyXWRPa6o4SO2TB4ds0vZFZLdW+j43DvDjZ
SCWEk0SM28URfhG0sldFvGhGcVXkIXs7iXPpEeeEXAqLbJ7/ChQs4lKVXDcU5QeO
Eq3MMsWvDmtQV7uLfZZiUr//SLKOzM9st4/GrUThhqO3E8LkErTcG4rmHD44avve
nJOXJI0833cyXIM3BhOagPW/hzn0X+v+rKYTQQrj9+hMcSxFdEHtDsXyRk3iygEi
+Qz22RTMYeGNcSho8oVCzt/gdXO4GIeV+e2FwRScZ/kBBUsfXRDtRHRjuNv4hQhJ
mm6QnAtR9uk6FaoydIWJjQr7RGCe1tIFHNPcw85qaa4njLOGEIGhizu4Pg5K+PIW
55B8Sycy1tx2EdbGDcsbMfEFNOdBLaWlpyW0kh/8ioqFbnpenHSi7UErbrLqkRv4
ccFBf/BZVAFtjDP+SAfc5REDBaKZ124H+NzFUbMK/6UZC3Hf1fkPGR7AWsTxqlf3
e9gGqeiMeC48glKAE6GW5wuwFxJXlowmbVbA70u1Fq1q4XcNeeuuhubH/aJK0uRi
60/DBcsraXAA/ZVRpAq6ZEBouZ0B3Dnhm5xU9bmi6rrDNeCJBvqqHyGqVWiUIqMJ
lLw593bn51pGgAgLVpybHCttoCodBqnbeWkTs2xHlLBD+5Au1M0KwGm3wO+IHj6k
TltYeD6l5WwgwTVIZ/hN26huo6FAnhKEMlS8kJGTyqoT7blhoc3eFQi+swOCgdzj
SyYDiBZxnPqDeEMiEC3nAXTT7N6AqKsTt9+4qKkaVtIoHcMrzK5ZhqWnrFJCz8f5
0P4669B5VI25jTCK8Y3KzuC+GJWTzoOeu51DY93chGXcelHXMr0rJxX9/uwHII5c
HInFJjgMUFHrwrfjTBYClWQMSflDxuv2gEDFDA9o6sFovCPLM2sZW4WUC9pa1ijI
jIVuWEjXh7WchFTnSehRRrWJdyzCGp61Wt1/rfwg9VnevNZCEVZ58sLGeb9IW6rT
McUFPSiZboZrSedfAOY0c00wXNZG4CeeFeSuyEnt8tw1/4lqT2HvWcDE17oFQ47W
yeHnxNm/vmOBSFQZYgBme/4uo591QDb6hsLRCBTW6n7Apn1YitZOBfycYRViBMds
dgR8p7yJNuZTXBSXO6v/F/d8/nVcMWLyMciBbvJwvTRVi/+OwB8Rt/J3bNEhAH34
qjdXB63w6545FNZYAUtEvLZbLgAeIMwL1a4ECJ54AKBdRBiCYkilzBt2EYEkGgGG
cEyBMrltJhFIjanNXKXZOVUXRpdfH4FBe+OzuIoYUywbjxZ3n97nIR1aYwrOcgkD
efdEHikx9HHtXBWGrOP0RrjbQDGgkC10/FyAnR6Ifzbmg6RUj4arjDZDlqgBKBEf
s0ZxxJq0vxu1SVtzVWFlLN+POPT90LGAOtBZdBApDoyd2HX/7QITJBal6ksLw0MI
hXpwrSqXBrRtCAD8KiQ2kgi7X+JY4n4gw9768BI5/eO1rSATvawZ+/f3t3xj9yu6
p8oRS2vbCQcGzGNKDKeQOn662RhgWHMv2WdB8/GFF+6tjeD5hMLAuhzUNdrfqjbO
ykp3JSrdvwhf9HGtwo39vMxG3y4afZn69oFpjOoT+sbx4mfB6SqTsWc//mguySWk
PbKUlCBC3O0jzO4//qjjegA2ll17eyDUelTfAm/CBO4r2m3w3jKVL820riSrIM4n
jLypkoxaNtVxz9C83RTB7yyFpG9Cm4LrplDo0QfsgBSEwLHUKTFZxeyZT7EW/PSr
3zJ8WiJEkFq/skCgDEPQcOKjiJTPM/zz8UwnNbh0Xm1McblILdDfsU0xRVm5R3vV
AdsIDJbryUfpS1HhYtq0Bn5s2ViDhe7bo/8rwWIGbek9r5LxRPDLuVT88pB0aOfW
N3gAw5l1MDf+Wda7FSXLtdzlRNTWSzMfMQtnRfMWHC7IxAWijrEU/k1DgBBE2G2E
n7G2pYjalEXjR/6bVBaGlCPRcy4uBOHlIuGdXz5jK/zs11VaRcKfpGNLoOJMXT5v
zzzOD272gsJWpdv027dDp/J9AFceFbOlU76J0UuBWMrPTUph1osUZkgCHibZ2JgU
3s2ziA5aluojL4cIRncSf4iVzDfpwngbV+vsKqjl1C9EKSQcIgicy8TYdUYvx+al
FI2yiEsqR7ieSqlCVYGzSJRyQxR86DXqQveJ/SNvHVgsCNZPR6/yuzpM6FyFdedL
dCwiamI5S5+T8+zuG6kd5JYMAnlx1OIiG7HkXkhbJ329DLtRvZSuXGQvZ6CaLtJY
7BsmrAq9uNeRR+VUsm0xGcws4iLyC+Yb52lWXAd8gEHw625st67pRBNEwt572lXp
02gmjjUHsaea1BmsS8aHMjpSM/gLJwvwPFFt9fGUGwB7jj/7UnST2i5BRoSTG3zd
3CBVeM1DIpmo/OmU1FljuuidavNBSmZ9rkeOj62jJqYrItRYXM6jcYdztw3u6f5m
PMsGI8CWUjxDCLHbxP/xsAxHv16L9M/fTVKbdqnG6G5lkMnk41ApnupaD4hAQc+N
qImdDXBt6+OshHQZ+3HUVYLy68O6r3Px9QWPbS5+XpbOSuwD8RDLgOaQ9gs25LFM
cerz64uRSLBEiSoL0tkbAU5mgHHLHy/W8xcaEMgONTLrfsXZ6mkhs+zuCZoU55Fx
T9xH05IFVlRvFxCbpOu0ExGZGIzyMazZbTIj7cQ+ysRU2tEr1THu+nRHhunh201y
H4P5nRiKUfpUzc9vmhufohLk8VPaXjZiiZd+O1JH3zr3dAANE7AXhxjHzktEN9NK
UpR+tCWOXZMMz50sqPDPSvw+fqVnWegZVpXu0WG6DeGgWSuVJ3RHRmPYN7nt6Rr3
K9BmtEytG75VAmmgqsDKrgaUDfs8iEJ3ZfiQi+d8B0lGo1vur2+/I6U6uYtlR9xw
hjriXtDBBaDnaWiNzIG6P58lHftzETi9R3FN1VDicoaD+fBa73cL9/tzohlUMLf8
A7FBboYLoII7FldMsBQAjLN+ptpRryvIRq9/TXk8b302RBKI/Daf5sPHsLpiHKeC
YuY2gAE9xVnLjMFvWYwb+LuM4jgEwi1OJnez/CdiSgOIkgOSNiq6uOzK7yk/ill6
dvhM97/PcT0Nf0aSxtBEZMpYo49LcQ5tg6vpzZOkvxMxSPTJnYRxnbox3BqjLZLX
fCjXT7ewnpkcjnhA8ZHY4qAUw5YUlknfH9RCJEU+MylFs4IUgOuBVERS9MHV+fjg
FjML4RKnrbAfVgCFQFoLKkVvtKg/C9YUanTi98e1GGYsMTaquHO/JPct8Ot/+x0I
rfjnUFhp46QS3Nx7mAA3ISsFC6K2tnDqV6lhFe2J506X13fq/xG3wYvxjcc5v1zD
KGXpWQggSIAJIauGfqqbbRz4uGgGNUNHEsntYXlgZZWTl6jsxQq6pKJ8Q7/jSgXC
mGWGMZRwuDa/4EMIBgyp3SDP1/emlFtiUswPlH6PANhgsgSFQ9UTdHQMcQI+5jp8
V6K3W8ngLdqMeXfnkneqgUlSOJyAkcHL8LKpbLI2XspWCsTn4z6vqwCyfOa/VXFM
T4gsmEdRmob6JIWJ/NEar026V/7oQQV4sVrCVz+zk1KhnDtrOSQGsmgK1OMKMBtN
DWdfYeu+d2zP6g6SpGkHknX4i0H3D+89STF4/SEV5BukmrBqgDusB6FbGvDh9L1F
U7PjKNd5atZZQ8uB6mTB0BFhn2xlYJaIoks9rw6whkDYPnAKDQyKG8dG6amZ0sW0
oN9g1DsMC/OyEbk+gTiRicehNMOCYRXOFNWkZi9OMF2KvxRml5kk/vM+xuyAjfRf
iXM85eW07lljLmwJ9HkYAvoZzTcUR9k+mA8NjHeIGCCCCJetzRdGwXIZPlWKB4L6
gueElMelLb8LarISZMqgjsY35nDCtcRlhqYyHxXgXHte/yAjd047bKWVTz7WnY9t
HQ0AOsFcywD2QYSsopKJMo8CrBB0ZBhVzQzJMpR104KXKh0f9vuPHLgsCmp35Hz2
NhfmmHZJfKx2D3/e6bcXB5hWydmI/nU2RWsHqI6JYN77HONBS3GF7TVHEbKytb+x
wVLVO+wpxTU/Wbwzw/ie6mOdDRe2VZl51IZ82Hx7d3eXF5M/qxoUPyLD3PA8kOOX
+swcnzmdLvjqcSRVLOQco2PDzDJbV05spd+tAoQmV0QpQGfrse00sFWq6AFnNxqO
lKOc5mEuDpXBL3ji/eE1vFAfnE9off1kbOsfSD9khPqm70oBpLWzVBc8lHtBvKcy
pP5as4o5ZF9j4RPXjwvJNnGtF5zk5K6iNeVNCRclB8X3qP/h8d17zEHlw7oNyyYQ
p1RU5ROYCY0b2ImbDnOHO+d+WzIL9pSQ4YuSzJWg8vPokjAdzKG77KCXeOpRMXO3
TM2X1bz7g5hJXa3/4jATV4LhtrPl14TMN7xbiJWqGRbw3O+KNEmpWEIVP+7yhpKF
u70ilwIm1yNY9L380CxjMLGQmzPzJv2Zxyd40US5vUUBTyQ29AOjdtsEutTmywhv
qWIOrhLBRDd2sbVXDTrkNY/gJf0Ng+oyc8dsOhtS5ILpMfxcSRPDSSzM/8/aJTUF
o+bsz6YY0KOcsuqn5qwiSCe3ICSD2+IjXKauL49om1lQerNXa3N7FBX+WxpxXXfY
lhI5YhrduhWUQPwsrTNoyS+QxSK7EPP7ZL6HwHKc5nGyqbC+M3AmYM1Oa8vhGNPd
dpEJlUTZb9Wf4vMGVe3wq+auX6jnUVBLIdlcOh60AyWaFyh/mmDx0y8sX8InaAK1
mPvMvJUZB/eARI32l1En2Jvs9XxV4xXqFo8tZ3gQoKJ/m8aqT3A0aurl/qY5skN1
hjisoFEWMW6hNNnyvgwLhaQcoNrekXb0SyFGq3i6EpiVYvSBkcVDYuuh4eGh5PL0
K9o6T1gfC7rWrm183AOuOXjxFA3rssWUUojb1rU9bznSP3u5zM19TlGUr2wJ3Qhx
Qze/v1HledYVSSd37mgMR1dBQhu6szirQ2Opv4jEWgXhsBGlvGouAOX9vwHN2INb
teaMWVIvJZ4wvbt5eFmGZN5ZQHuQbc4ysBMl6+V0sHbECoZ0c+iXVMRqXNSe/qbU
GFWAuZQyfR01g69kef87q0BGrVVJZUsOpvck9V6SKLyZPbdbi4/Ly4on6iUICrn4
YHFSRvTG8sTYF7pfVA7XcZnIM79zQp3MHsRkKgdzYOlVskgjZEcCu0U4MMOfKsG/
fWxQOQXAow7NIdVFPfG9FF3s8miCX0BkcvZTXNGcasFPpyEdzhJNlo70h8lJvU3t
/UHnSmjqaOyhlxfEAZmhWrqj8zHMiqGFwKybwbo3t7CyKu8aa+r95SA6CzegAErt
V8GppnhkfyLaVM2JNKObrGbTuxYxPFYPmuIfuQoO3ERiO7YmCw5CpJWZh29kriGf
YBi4iE16Rj1DT+a8Tji4FIAeOjaDDFqzXvNFLzC1ZUxsHeHgM1B/fXkhuhjtN9ap
/VnLy2F5oWku2HWgJfwdDtW6Z17a63j/SFwGFyQz0pVanugLHw5XTMY12lOOvLuh
GXIlHhh9CVcdruMerYfq4FsxrS67ajLUuU2lTRohfjSJo0vO5tGJQ30TlWY8d1Qd
7xADSD/0goR3xn072un9waCGvxaSkL8b66PwadaJxwyRI00XIMiQ/6disFhzQGHp
/dp6fEFW/JIwKIsvZOxKXuIu17r20QxC3FXZt5pCkynU9QWWOzb5sunIPkWSW2Ui
5hh1InZ/g8CAqFuh0FtsrJblaecHqwLx8ivoSUkSru4R1IoCdbkPZOK/LR1ZQrTi
zvP3e3jWi73eB/azSQLevwY3w5LIKt8MPzoFmh1Eyz4gt8zuwlGHrW+q95HCQ9mr
SWoC0Wiouq65IpM1polHEitoZOdv0F1DO7WG4fg6SaV5gIe2Ska9EPgIYQTXOdEc
Df7EGdkezOsxLK6EBcXiW0Z7yN+rcL/IKvg3LkVoSlLDsADkQuQAtx5F7ZEwK984
xwUoS2GryfaRiKKtkxEBQLHHsGZbkqNiurtKagPPPUn7MW0of1DuZsUCWfDytfLZ
wqD1ip3ruQua20jPD2s6SGXohNN5sXZcxk6jSQ2S8N4b7VoBd5cAN71nohaWwIBQ
dg18su5/2DmDK5mTgzqa6EPcwJrTzVql8UhUX/M6MTJBuU5WkN+cZXa32HoX4HRn
p2ozDmLPiqftTW2cDhjW3eFdEf/M45Q68YfpZmtAZjowZHE/t/V5vn1V6xXS85lj
iN7tWwqbZltOZWSPgpg+7Tf8yAblU0py9q9u6MzJIhUy1HF3nprJHxEmh4+RQIoY
JJn2Ogkp+SeysR7fgs2kOwSmuMr2rc4F8IsOxFtO1HSyS77GFaAeGtl+JfbtfF2L
YME1J3zzU0mIp7R6Heo73SHL3dhZg+bwg9q+7HhGoQT4Rx4+Sjfv0PTD1Qri1W66
5hZFvZlbF5x6zQUAfAZ4lBvM3lGRYI42fUYbfjWOxqHfBZy2mJz5CKE38yKVL19k
QrNQaNEIyJVMCTW/8Zaw6QF1nQ0dMiLnlPPWXONs/EHhjBePmmMsuXZg4OVD/y1F
WrnsAUpfJK6NGOtuK3kfDLgHuVauPgsYaGtNWdEh0deyV7W8l2cbqwbWEeNcD1/M
oWcgT99UZZzWUI3EEkEjsgRxy2w2Ng26WAYNZZCn0Z0V8kIdsSjyIe86VOj0A3a9
3weKrOSOltHsfza6fyYpyN/Hw+VItka0o8aVkK03AOdqSHtYgz4TgigQHEmf8WPW
CePULcfM3KFycA/6QerfRtWt8OMnt9xYjlbftf0bBl/BwvWf8W7AtT/QrRTe4EO5
dtAaroHuSOoPhqJSae9W8/2e5/r7O8bdY8cwzo+bMWgWU/lXDvdD9xATZ4fN79+3
yVogkfZH7axnFoncrUjIvseRQ81FRrExHJ7QannmqiFMX1xpnCnDmZw13nKZ6yTY
L/DCfW6weJChrzyMBthSxlAJscf8Pe+WSMQICc4TOzzXnf9ffXoT4H7ntHHAUpcV
QQwVW723e80Wui0MFjxzLiqDGFRG85Kj07Nj3rrAZBc8ibIO5eBlpdFTPrJuUp7D
CUp9Gd1kCV8smR/jqb5Vse35h/8Xa5pmolD7WvXawHBlJRCtFncOzC47RSix6TPc
KatHtEHFVOGoeTVJEf59DSdvQ1STqC5eSYZL/8uPpCTZx5VWBauc3efqbPnYfxla
b3EY3xZhCxPjftd7nFnNQNIDG2e2mntHcPU+bcBKYneJlkTrXBkMyKG8xLfq8HqO
/93GY7zGL+7n6HMicu9NLH4s/LAJMC5QD1u/Zi2nlVD2BfWqjdb7ZZw112oxdVgO
WXQ08BThZq+0fCSn06hzKEvqmXqHgc2mfRm4WHSR6gapRmUrKov41E6uTqU9LpF3
yr0lL8wQ3/nG73Q2h4VH6Acuv00kSx6KRNpsv77wEuLoQJooFEWHpAwVtOk3XxkS
gxlrgArNVj+se2qoh3kAJSIvY3oFKZDpAcTGAXJ/BZat5H3ME3p4PjY00EvfFP/X
RVquvxw+lqpfE50VcRBgDVSGAZY2rB1P6yzBJ2xESfNPIOqtW4IgZqblJ4+M8CMh
zStUXJgfhEKzkFHfcXDR3ns1PxlAmmuqHK/nh7FNjx9gx2TEIlowSUD+d4ifbdU+
VpVJ43p3o51Vn07nOjA7V7ODEtUwgUPyb/BZjgR6svaiOi3qrr2kwPFjv/lyrYAD
+vx4VorMAIlJlrAv5OC3jvymBDdWQw1W5ohMePZBiti1NLiy8Y5bfjWWQbijWMwB
ObzPKOESW/ctiPzIezjjaV4bZbELJufBPy6/bgZ11LACWoTvtq0QuibTpzMIlev8
gDAQJVkm8AJjREhTE0u7TRbPYwRaUdwbK1UBo3kvloJBOArLdBm2O8pcfmmhuNmK
zAP71dlxdLVQijhVhOTKHC34gx/K/SzY84/ICqkVSNvAPbhZAaS77iUrO2VlDyZ1
8Nd1HAU+abP82QpPhmC9EnxeYlcclmozh3x4D2Fiw4Qa9wBlXajV5XY8mEzVnDZf
UZczW0aPormt9oQjsidH06cxzxJm7uxvEeLQsmw99PlMCPUPZrX7i+ZTHQKLjcoL
0K5CyNRQqxXkX7Bhq6EBNgO74wuzZ5FkudFy9DIjMpfUDMqX49vIUK9xlu2zZWXo
yoKusY7LRIXfcjoSTUz4qftA1eSGQhgugljbHTox8Eimo+ELCsuxtEGlHs/QV6dR
dSkHgxed8RovpyoJWGFIEPzHrMm537TKFVgAiz5kREHkG/mYo1pINQTx60Ous3s0
81FKLDStzB8j5oVlvhiKa0QcF7FTxbT5QA28mNxHRTVKMg/kuBNhcW/yPUsIVVFD
Z9X/tCEH95Towldp1b2EoW4GgWbCQMw2dZaQautUHFkAKQxIwwoVzPNAfeZDecoL
udNvV4BHB1IhpY7toVGDZKE9FQ1KrvP9Y+4SzrHw98Wo0pKUmkR8ZL7VuUMV7J8B
P3O+dZChsKZtYiyQFp8LWo0FxU1gOzRB6kTocZU0De25VkatllmXjB2qLatUUkmt
jCU+LdERV/LwVVn4JUTSNMn/ia7dPRHOjkRr9yNxTQQN7btU6d5adtWXYKw45jp9
7pVrkkiHY6w/wNvbTrQffX93lzDCDmrYKpS7BR5ZUyx2LS7+Uy9HeDPZz8962UL5
1dheG5O5N1DtApUqMxBh86w0YPAR6+4JoK6wlFTzHwbjy07/rsR1Ib1BIKUc0KQx
7EPma3s0O1ctUe3kYx4+wAMZ/Pnf8QgdT6yWxKf94Ncu7FNijXtQEnkSBLE32NvE
uQCKN8+0vGqjIZNnOp9qsVMFWn/2i9vtsB9TkwwhNhobiYiM83q+rtDUipTIPpnh
ol0mhadXRQzSSOVC+rhREWY9nNTuxrLVqI1hnCZdwFLfPGGqm7JjdfzypOfXy7Zk
c7+ldqJrJbtq/yqw0Rjt1xw+9oMIXGiIJYoA3tLtUynk33qmJ1aMsLSfDZWbIHYR
q7h949JxCFDHfyaOYMWnOro/cK5regdgSl6Xfq7ClVEtnrVyeR1sVq0Kt5Pw7jQ7
JYdx0bjiahQ1g1BrmGxWGwL8W5qSqjeEsbekeDGz50MjLIoKdsM+WUo8x/3xT9Tu
M262ofH8ae34iFH4688XTqiX2hQP6PzEoEwaZjooCHkFrF35YjvKcAY3BLk1tgUl
Uf2j1p+TYUN9nhX1uaY6bjMVvtXohQQAZTIz29DPCPPD3ijDq0ENWU1QS1Wj86G9
dym8FLl6FUpTqVmNvJPS0a4YTb8njNAzYl/LaELK3/1W5r/ZR/qu7uplQSlLsJsY
0LyiJwigIQSjZEoNu9+eGffOxH3imAysT4Vpq+7ssyj7Gm32PwjHW2osNA0LCfEW
intBUy8PwJixCEy624OJCvWU5CCxlY0Y97peMiMjhc/0KEMjLkL3/mLiZirtKDwS
RkmY8J1wLIOoglP6PGq4+iV8SraeKafPNhrn/5FPn5ehMOsrU+RJSSPN0HzofK3v
l8iXr+hms4sW2miUAdxirrIfSZyNmYSsBNfsD40clwpXEIW4O3kSM9UA5n8wRwSX
XluIGsZEkiZ4MS62zNEyRpWIEv1a1yrcz42fvNlJ9nXp9Y36krhYTshCHybtet+c
amMJlxTeVJqU1blB/M5Jiog61a9fiKKZXdBveqOVeEU+mVK+GtBcTpTiOHucXP2z
sQ0VX0hllzS+H9W33otFkTzedaoBMosIhTNt/IkCjcJZR20n/Npv0imbPeLkeQpf
HGrGjuBKukFM3PkmwwsElXWTRolpjyUkZQFcT4RNITe9CC2Tlvin6V63YYUBZDkl
lYrThlDQLHMF3gqY1CRZO+HWiQpXRs12hBNfUsBTr/WeK+OYFEnEdm4IsLVMA8ft
pL0/39C7RCKwhjkECqNPxcG6b9eJl6BDysC4kF9BDMuRIvlV7O7UaCn6Xhc16apL
bjlcT1AwbKZI550PqQ8uwJAT2/r3mhHn4901V7R+G15nOcf1OrpXhbGnkLgI2swY
UpIRfzIPx20Bgjv7SLoua5WNJXIKJv/mlMEtf9B0jFwSTR4Ea0TjazXTeCwEQ8K1
FzbUJlsUn1aGYOrzmUyzyIcx1vcourSNYZqfYNz0F1qATbO0f+6CPHAlV7BNik/J
gl4gB1wps1xIfXbvlsuxgOPvjVsQClS/icl550TOI7wowwEFPlf6b3cXjGBcIfSL
qnFTMuAn6jek2aiAwAxIAFEEbRTMVwXYY/OH1LSz/MRvCiBxd3dQlGKF0V5oGtSY
hYnJm68tWVKhZ8CGMuKIVAsyAR32/dCQ8mvS2VB/OzdeZeZJkYZWF4JHSfr+WyZJ
3X2t0n4qENP8Wnnjk2KI5dd/xXTbf0/jmvGqDQ3lXfJsKvH0IRmHjRGHY9T/2K+m
/MXLM+72zxgYh7YmGzNmdbujVPiT31XBRcCZl04uEZDVQnjz6nlmeKIfrcSNSpFF
3QaKir+puWr7rEapLUPThJYxwx86IOd/Z1Lw9DmSIJ+qZ5gh4Gqv1ryVEmTjzXRT
4EYzyMp4+IeKQRjkuQpzVsm8/KLcqPzs052clNxiuZ/mXLWEIT5oeqanH5oUKWgg
z+84Wyl7bQRnt68NJzv10Y2cmEhtGNOuq854BvLYHHZOHhd34SF9Iw3YNHTijdfj
TxoQbul5S/9YkLw0QdCoNC/61j8fLmdCrPDW7ydUt+VY+BCa86DXTKdqh1BxXxwc
9aUwB71VVIrIN/nN82csETyVysORQ6cd7yR0Rv23G4dI9RbjBRLLH1xBQNIy2U5v
H51Op2lrdGQTIBNjupbwxaa9UMn5AYgfi0qcBfLZvclSDKrCBzA2iX/k5RH7Y0uT
uHZqqfTnBFLnX902uFZdW/cRoTlmg7oRirxhtLk+QJiqCBILIgKQ2vnCVyO6AH7v
2RTovQ3IOfWxP0p2mN3k3aa++K4jxip278DNRzkWa9y2YF8DLI2wCmpxJIaXT9X+
a1p2cuiS64b9vIcpqCEnSi/5+GL+rHxiwY3LGXKGC7pqWBI0JGBs4WsK/hLkJPwf
+7ar/pt6Nmwmrq/Ajl+Fs5WtSo3qQn4/PUGNa6MVWZfS1lsLOhWyvLX/xIDAFPYW
Ig/2OfUsS+UrtnxOo/IcJ3KuHmZKQdcphQU5c84YOVfyoLgvOLrgh/YOKA0qPEM4
1dMgQ9VY3olK+0VmbwctT5iABekggl6SUWGEqE8nrVzDXLH7nHO62y0hzISi7Hkq
NN1wNTwDyFa3MT+Cj0s7YNKnfBuzlN4Ox9TjEaLPmua41//Ck7YakdeineDaaa2E
y84JdYuAf/ZuAY3nl9vkYoTHDbTGSoFBEVU+Ig4kRH3xVHszo4xtlOahpRtLbx39
dc7QG3STRrbuL0HnFgJw3gEDt1Op9oE7YRXdE6AdxzAvqpYQHp05PxSphYr0aDAK
nYLSVM+jo9SwydwQr4AfsKCIG0eafZohrAuz8eHZoh8B7fPYg+O4at2JAf7T8fe2
M/JhTilKFRaTA/JMEV/f6hn6VrOsfnsPpIgWH+vwUm1QaCVaCQywHlilX53klHA4
9c2rcuhAZBdNKjvRy5POlEY5EcAqIlLE00k/1s5qJ41iSwxntx6ZOz+lctkBvhR7
dA/12hbE7qKEHcu8TyOzDXpPwzwfTbvQXjSPQdwICaYnazQDPUERSm4xhxMTay5J
QjtholmkhIfWbn2MZgqCISUbFZoouv63VxDn7AsYJ8xzP18x/rOuY4X8xgBLlUWJ
XErGOoocFXbbYA8niW1AcNmrxJr9zMkJZAPiK1BxJFivrqsZ8V+Sp2oLlkBuxJ7I
ijZ5a171lgb/AXhE/A50Ltwf5BoqNj4d3KKZomjSAkjqnLxGg1QgMRvNAZqQncRD
ZMprq0gZczxxi/P5nZ0NvFBhMOQ3IkCeY9HZsf7X+/IbBkMoc/TkdKZJbdCuA1UJ
1pHqiJcGtj+OwnMjoB87wr7VHitghYM1AnYkG+uGIIk1pH6mPBo5+5MNmPMu7hMN
DFp8oeNf2h2Ao34ugVkCeuZBIf6XAZxQLBm2g6gNTCZdKKR5JIk5XHczLN7LzwHo
4gEnAtBbv4eqP8SlwVfbR0nZU1LlfUyZKrRiJGfe4e7C0loKvBJMKFo5PCqE/X/q
h4RVBWzfLNdWRXi1MIptCbbw5AYKw6e/8BI4XH5ZcYN2prjqDYLEUyZHY89L4D0l
ddFjvEzns1JcD6sEQGFiTRjLhhXsYlRsrvhkHesSFmsKT90cFpCslGjlQ1ELjLzW
tPybKbMNhG4RUTFntoXaJf0j94+xHfzrt4VaBBPGqVIyc2byzhrajchBECtaXvk8
02FaHpCbTrcKlt9N9F933GH92Vhd5OGmM4EqlNlGCLpQuKtHFKn6FkXiBcKo8+fg
dUI3r9VWN6/9gTpqy/Mkhn01xI7w8btQsqdL66ShK3tH9BvuyKKGTKGgQelB2mJe
wX4kq5kcHV9qImGVboKQvHxKYMrmilBhIRhoHvtWIg7DFMCvrMJl2f3PBo+1tehc
+1EAjZodQG9oCt1Qya2KfBu9TGYjC0XdSv8Hy2Jp3Cgzr2IVLACEY26x1VfrM5oo
OAwH1BRMcfoxIZ+Sm0uaZFM8xqz+nNdgr8OLpPbhSx5YIHXIGgf1yit9ZEpDoVBr
zmM6i+QpdlcZ2Me8AY7FJyEtQXV8L39HNk9W6TVJ4fc8V+EhpgXZPzbD6OxHWpR8
A15FHwMpxNpibtMquydCguL1R1JtoVNuRhuYwFAiG6XnAcLt1moeiYWiKuN80h72
Dh19cd5ztPpX6lA9mflsqCAUHnqp+CQMwSLVWxQAQA/hKwy2fxor3/pIYOBVQoKn
ovN8GkS4OkLf05aG6BN/NV5BS/u8eFKBE4znph00pgHdytZKw6xPebuK/c8YjAm+
vpmgDXQDHyjTclqEsDmAqBWdi6jT5zBJ0tj7lS+K+Nrgm8ES9l8AkR+N88FysRJP
0s6Mk23Mzw2yqNA/eKEEt7cOgticZnnBGl35noJvtJ2EudZKXSb5VWuW8pVEzpUL
JFKNYAf8y+rGECKJbd4mFSI0v6R8o46+luD5RB2CaLgKnTnrf4J5w4BRX0OOG7Lo
yJqBXkZs/j3vNK/27kJ+tuFy6FEUa/e59cMP9lsKO9IigyaEpMt9fLATSKyqFgUP
3XPA0I1Yvq3eORCzVmobV+QsJYYQFbsWrEbKfsFvZmeTm+9X4BXFRaRwlKuJYCfP
j8zqm7K74jVycYjExMoNEDwSCNsv2UG6FFEqPtNWZa8YuK4F8Ben0SgnUoeC8yH8
nSIhRHB1SeEDeYllUE2Fd7Yi27CX3ReHl+smtdRKyHLHam6YWGSTMQkaaD2LKgJX
5xQwinXU3bAz77gCzkez4MPyw9l6uJHbu5a5M1Uj7XRE6tN6sLAOCD7073EMD6CS
DqIOhVkSidazfkOE4j5t5ZMmISLSpPYOlHmczh0BS6Aim37QinMZ1aO0hBI+a75k
rSLSIoGRIKJrM7R7LhvW2htMXzJ44VWIHV/p6WrhQPMVhFiyRGdiY+8hZ7nm93gd
w72cGFA54Bl8B7BBHjvSoMSCqhVCt5kP/zuMGYmsOM8AqymByUcl6a9Ac2TBfA10
fPa3AB7CZlyN/ufr/NfM8G7ru+ll+Yxiurt4PlO5hb0ykR/JHKcvLRAedtzb57lV
NEiDK8+9x/bwvkHEEeSIaUMmnoRnN91vT9fLqk0QsKsd1AvF9EnPfTJt1rRP3r8P
WEv57vYD4cP/jHruLtJ5aRNzqNYQ1R2jhPfT8QlqVZqKcGBP6t3RckS2CRx8AdI8
zGYMIPpJnxzaG2AQyCxBI+aVkvjbF2A1LIvVpdlxOdsayG1/+lUCjoIB2DGmXMmB
N6XBxaZlutMyVaz8+P5ntccFLkJlcDpKppFyHenD/Sn+I8GLCi4Z81WI7h7vzEJP
QVGCSztDlVLzYRkLJTSdpkGMyRYaY7WdzVdpak/0XvZ4WgkNXMGrrODDN9hPe7Kn
cB0bWvrAOZcHPUQt0U3lQNjUghhyM1+Bj/hfFQCb8W/tGK0HLc6aVwptZFgIT0Zd
9rGRwpLcXaNxiceuqEW4rpwEh+NGqTjjfqNksxCpIO+GYMxNF4+HDLnpE4+NjDT7
+C6KAWuWPliREXGSckGVq7jAjIGnKqXMH8TDYt/wkk59TQ7OAEk38ccg8pL6dv3G
ZjzqYhfTFB/zRMq8GTJC7NjzeqhEMTQtu+SZWaiKQJfdvTbbRpD1luBxMKo1VCbY
OesYUfS9gKDtlQgTdto1ZHvgs+fnSVU963laa1MUXltmUYR6Vjyt+nKVudHztr0U
v3l/z+Z2NJEer2YLV2JdPWlh7OQFNydcffWZv8LlbEJ04BBx91LAyhw+0QiS/50P
gwGZ6JJEPBKCamNK9lEG3TJobBTEzLi3xEsnCIHEAickJs9V7QaqtqEWsnxr5ocn
NqvNWeCfKjGEXumth/kt+Sl4rXeysJtgcsW1469U9XNT/c6kc0ZpUqxOVficjFm7
7Zl7xE0zH8KUQEFGHTJmy2ReXB+J+zuzzegAujJCPnndUqtrvM8q63KYoad5SmFM
yrZ6h+q0j0cfxQhlFU6q1A3XRsdAVtyVa5TqZNDDb51GpAHttyVL/eW/HYD1lOB4
SBNe17Qx1/TZvnaSOO8S1qbVrlWJyEzGHwD41hTZh+vQwfILCIwuuhQ7+QkHSN5B
ucakvFo9NA3SvqExTJjG+UDIZVdxC4MoUnEhUbJqdrmQKa5nERnRoCo6lP6rXnOa
H29PKooWe8hngcur8+Em1iEJutnXTDin6ZT6uP1uKlT4T6Oa+AS5r38NRW4CH4LM
sWnRpW3lkYPy7J9U4YCfDv5eRT06ixQlkPTq1yEos4v8iRq3vh0N417+qbdmtCOP
Wmb/MybsEMHg5onpuO5Ji8WdECxExW7ZwpuP/55N5h/+1R+W4DoqW7eBZWY1DfjD
VbF1zHNhaRQ5y4XdhBdv8e+Au6i0VCkbyLZQ2SsxWVRpWMA1VqsN5HHza43sbV9g
JRuo5oDcE+xqTYCA6DBmowu2GkS3pjfJLZRGjgaN2qM/NMUMfcSLMelL6e8t0NAW
zcXOrhb1ajlc5Stntjjg02oFUVjytZ4CpTsec4ymd0hvj5Cxn2D6lqcFNyMHLWyL
uFAYLxdo/Y/dHJn5OrkrtwDYWTTYMEak1Dw1sEQbGy8VPKEhXVHEK4AHGOGZDwlF
7m+YGQFC8HS52CkQEuzV3JtRFt6SasGmHuRqJ0D40tjVi5alIsBphHi8b/etoUW6
mT3hwvbEqbIxtZgTvluLIcpOgAEUq7tsD4lPqcMdNNwpFYcxtqqZ6HbUhfRg1qNC
r4ijkG4u/N0YRCMNirUs2/N2gT3x+VvL2wzvWj5NZDVX+lauKnz1pTo0wStQMs9f
AVWostBUYz8fxS45ZXbRTazxsPMK3Wrs/bD2yw2f2Wqc2y9mYIKTQLLzts4rBy1L
uGaqMdSW6PEyfob5qpax7UyakH8rDwzBOJDwvXWQAtIHnX/sGCgNRHQT/gsbV80V
WktNxCMb/Rbb2Ds40qIDtGNF+/4OQV0KsD56STvH5+4wrO8UZ1KPQ/ka5jAr8Ahl
T2D5kiw84brDkc+SH89G0JMBL0StNM1fWJyku8nlpF/zJ++pv+QYzdjBNVamVDmD
KlnzEaMkXfMxeg2OV2tREHgCKe28roEgnwQyxgWXMb+pJGnxjmtz8qsPz3U/DtQx
XpOMxoAvEm6qLqSdDuj0OmBR7Em3ppJZmqLeA7XZo6GqToDoxlKIZ2On5Z69RffM
fHsjOP+SPQDVeOsujBOl4a6YNONAYh0akREwfYX9vpQl+L/MEV4DhReQIe1f17uk
4UnJ9XejulmBWtK2KtrcbLcvLLYvhpMuaw0z4cN02p6Elw2wBdWIPG5BsV61oC7s
dt3nkNbpUEz4D/5JdaK4z8ue+CnhmrczghT/61OMXuBVIFPIPWNbDCuqKFR20Sz/
6Cq2hP5G75G2kTdLEulJRxNjbg7rWCLjFhYllxxEPJqqKzeM00Eowtk4dTs+ypTT
2qc+4MzdV9JREs/iyM6DlhehYErHFEY8VgT+JTUhAyLDtqPNsVozuXn1Q0lySA0l
VjkwP6grKKz8CTDQiWLuxaiwLYcjEy9JnYJoy8TO6lfeXDzIyUideSaWPwuR/IAR
LRgfD+zeCUHuutaXYppZjQxUOX0Jl897EArGl6DB6ebs5Gs7JUKeGO5WcyX5dyUw
bnRmekqJLCQtFYPoPDpMEEXE9oEf0N9DvJTLkVDRGhT0llL2uSJ9j8JvX2nsT1AS
hZREl3rkG6Hg2GPDoSK5sljYJ5+PJ9U3g+DbcUfxT5nrcntIjj+sU9t1VBMIugQW
LKp1KYRgWzUKcLO1ip+V1ByFXMM0mUxcmpj3n9cM76DfJvuBRWKdtebayMPj3/tb
RRmn4zZJqAePnUHahvu1JNAsDrpnAlMs7xDRo5NY+q3grT8QEU3X3QcjJIA9SV8g
BYQbOXBN01UhKkUP9nh1yfwGob2QxgTuIk5rkF2mkmn4j8yBfDEntD72eoHhjD2B
yEyK849BKH0kIkLB0xm0aAB+Sw8Hj7y1pM3j99coDNmP0FSpkWcaAG75ZgDMPVyZ
B8+gNwIPGgUntcq4KrrS+C0QiTr94QGifSGXSHdhsd7gcGwEWe5lYxNMixGoI/2H
RNjGj8zLuk3alkGic+lfqYfhYxd1w/yID4NnryfZE7xAB8ObugyWke45yuOB2+2h
sOXXCeeDY0gW2njqGZaYtVfk+UgnoSXn+0TSjpzA4RB1vYF+hedSPBBL9qA/6QJB
lAM/PqSlkBz0gGwli3BL0rNAASEfpbSAWOu2SuZLfwTkCSByNfAsBAsuajMP8gRG
+fqQke7nqKRFZzKf9y1V9fD7cqODLeH4y1ui8abdOKpHQpU+2gfWb7G/oXxz/4Ni
USLIv7a5RWZVFa7hmPle4Z1/DqJcsmd5mQ/X9hCoM9TwBDAaBp8wNexpHwQWwVgj
IojHDsYN661jUTvRww40sAr2QIkJoRZsey91ZPCY8Nf8R3ElqybTGzT9dDcRZxWw
PBWGK2n93+5cF3aTuIHo0+pyNx6MUY8B7GzS2HS4hg3laI4I9ZHi2vRVC53V6FnV
qB3lAOfcJHv0HRU5nHcSVZ7mQ4qvR2cLbRf6lirvweNvwyvVgXZ+a5YqeQVZGlrL
tJ2i29NIBvCJM43BNcDS2gtepUzAV/PkgoBuPYSLrBKVQKR8EqGWRAx2hvaPv1pG
MIu1KiaPKcVXhiwfsMP05o2MWmLR69AJ5QASvAeHv3M6CNqZ8OBqQQv25oWh00mK
2nU51FV4FIlzn0G1AP3k5NJuRPmwxQLpatocUqSQVnMnxjAvWs/2KCfkOkfeWEif
MLnPO0W11dKsMatIThmCDmhbpkge5SDpI9JlQIRH96kQhGUnr9L2leggj24BdA2r
+ygFpggBGgvDnRmNS09EeGtCKDNuqQRUEb8eKRA6l7O2es/ueHJmG08c8dOSb6n1
w2IU7INLW9DFOcV2wt56Dztuegh5DkuOyQYh1xDPlLRlaOWQPebsoZomCIjKoccy
/MPRnO5NyFcIgM6jCjjFcoTKYZZltjQII26Vo7swjzxv/vmegxcfMeW9ZXezw5c9
jOVaAsRw1UoMzXzTL913dtSTkgB3BBfT7pmLbDxh7/IFAmR1dD82W3Yl/Bufg1Oy
WI9di4WWoJ9K9mWAq25VuuzDR9MXpHNvjDAvlQTOR4uqkDSsXv+bGWP0wRYQVDQH
cjwhdW6h4KBBfzeK2AsrvD8DtVH3e8GvMP8jQNfN5qnt709E90no/OyLm5yC+W0E
BXJWPb/l3Xid2CxYwHC9x5QyEgDEDaQRwC15cfkdPaC+O/uzOveh/iPaXfaedv9u
VyLwoRMHMxt+ilWtmZIZFMmP7RJURpWjnoVJywOnT4FLLUyT1Y3Cwq/hCV+lgF1z
aqi2jxP1YNfIaN2RfTGY9u2JYIgznB+VM2eo09Hf9lMsvRnlkVPH4G9hKIt3DQlT
KNHZKExjkhanqu7Mgs9wU5KeEzrBqAhFtrWc64c4kJV44Cr6dSTqrWVSO9ORK0+U
fFJTHckKMu8TKdEOEW/GTsqO5YhWwFMXcmas5mf+4i+C8DOHcNnDMBCzKalhAnR/
2M9LCohic1QxROy2f9oOkJmk/ZjxHl7Aqjm6eP5wskcPB61IGu5WLhQX9MC75UYh
wXNQhYcbJMrvJVsqIola5iWfmNBF4YQu9OkDDuYCbARW0aeppDQP1JaOndtony5I
87obSMOk5WmSrxFqLlPiCR2Vs128UrHLqrnZ06g1yyAozQyNkjU8shveMZb1fXtf
xEfNwpPiW8qMpa1ZS6dM0jiCt0wuPRrUE7NgEuSIWaIYcVpaOlWcnEpKtj2twr3E
SFz+Lhz3HVyboz/ldBByrSjB0R6dhx4UlDcjMQUv9FVUxjbzZzHS89a3EUphSfs3
dbDC8u6pA02DRux9MW1Tn/n1B/3rEda7noouudQtDK4QeU+UzoZpotUDPI5Wl+T2
YCPdAjctEcct4HcKk1e7G/M8/e9CTRh9MrsW8RMKgM9nZll9juvSy7m7Spty8CgL
GvG4r6xwShN/uKDEwsI117sL6GEWNuA7YJJhYrnPqaEZukCJAjYN5mdIjQJfLxIJ
aE2u5UpBZdevO7J//IBVNqVphrHHUvdwPwTRwRIVYYPQqia8as74pRbOYjmwR/Ic
X7FSKIXON/q7wsvNhev6E+k4Qtrx54KYrqXAFtqWLOScRMwFqdl/CZi420cOBqwX
22lMcRLheXW1TtNWRG4yr1keGVW9DKWeOWFGH1ii5h2jEr9EHs/M3gpwNWWEOWp8
6WaV2zzOcrTQk4liR4PONO7qckGe7ZxwGXJhsgEUXDDTy2+YQE2MivVnrwykUFBC
TJlwZ/cTy+WSBGApObNWt88MEtP9JfVb1fipeXss+H8wOeuwD+9UeWD46WiYtIV2
9Q+OIYG1oXBaf5vn6xYDclbpZHAIIs8eXnelkoSq1uEOI1CAuW4KqBVD5TxOMVqy
H+oyRJCGL1zKCmrIKwzptcRwmJh6xU0MFNt72g3n9Oj/QMpZ4s5dEEirJWtr02mk
vVWqMEBs/ZLfQtvaa+0P8YJiRVh6PJ3whg4akp6A2A9jNb8vVccdiy+unAsl1EIZ
KYQHuFxhgBFBZ0/Y3/3Ti5fpXalNRB0O8iX6h+vuYt9MKjtVrYTVQvyhjJ2PWKUF
qrkQ4llDH60jZeDfZwendSNsQTi6lywuf4pliFKnPxrDSM3pFkFqdaJSI/TweGLM
WYpMY3iJesjBbwNn+zLvPqkldnr5hUTK9scsjhqmJTRWQmQmqG1AE1qbMpa2f7Gv
vJylg7SzA1KY5S6LP0ge/mOGpxGIvyfSrJ+ynnRTHKLXS+sTFJRb7rBn0qulnnak
H7o5+OR15g6kn6RNxgdEFeqYPNSk4XNqDjS/DmeQuuSE/D2VRjo5SYpmHe43Jqpm
QgglgCnSReqSAWR0WLgxTTxiAuQ2GfvKoYOGLRq4lUK7nbcIn5bu05HRp3obPNHc
Y5xzCXFB4/L3A4X3vPxD/mIWeuIy83RONr5jgJMxpdteUVTqITIwmEiRlQzrWusn
2xaFlsM/B+KF/aUlqdcAcO6Z7qt97v2/CiAGhK9U8Ye9p34/tsAlo5glr5yBbn4f
r+1THMsbn1ELSYXRBHvaDNUlCmHnUEF7TQa+RNwDXXYo+6Hu7jX5K0/TYVO0OV5a
1sJyz8RYgR5vOUC+IJ8Y/CMlH1hn62rilYJUyFrLUUFP6f2nS7qku0Rph8fu6+uF
PgLB8a4ezgUSvyC2AYbTfOmhZfB93PcLdTGu/ZtdlgdKZ48WGMD6XKLJIxN+sTFt
v4V0/IMqciP6HIrSCrYhESlLOn/eKqtAQI0qHOS98vcBD0C5ggzOxW94Kfu4WQXx
wrIwPd+9OLDVYFwVTiGbXVNMWTA8LUAJIman0B2eXM9Vpn6uEs9LtO7F7Eoh6ky3
IAZgz5VCnQIEG0y5NPFnhleqyGNmJtMoMNbtuyA9uIwVmjzuXy5fOfkrTglMnWjt
Z87FUSjY+iizAmhkFBhqDNc3mqxiIP94gfI/iAs+9/vGYi6gYiWlJ13Fj1xKJol8
hAUy/UoSrlhqhtRGXw1hgpbvIZyzygf0/MNzr0ZoRJPk9+O7goR6RAwv5ymrTYpV
OG1Rl2pk+rWmkP0Uy7EzdtJ4W/v689zoLeX256sjfqx489zVLB+h60z+nJjrKBEb
wMNHmt7qtAxxO5KPKBIdHIKjMwqMNH0Z+RP0JLZB/6FtLNMENFt3Vl7phctv4DOB
Wiy+zxm0zucPUW/bfllVWQuvd7G9K3AuU5ywCNKfHfhQubVMa85cSXz8XAdvwazT
swoZ7XOKl+yHLfaGQpTQokXKdHUV5dARfi1zyLW6XYmla8PFMMrBKx70TJzIfmf/
FjNkiHdCuXFv+G4pQMGsJbrNTqVUCpbnj0XRdFa6KtXB8N33kEgYHwxJqFrAF0Wn
OQ8wUWciUmsQJqa45eGMHy3UMSYapFBrJWx0E/1vUd7usUNBkmjjPYdt/U0L3tdG
jU8q3HOkE10F8orc5NL9SdcpGevWcOII22NgRCOIgWd8BoPidAQYTPB5Zj8w7qsk
lPo211R0SifV4xw3XscG/GRoKtUR9H7Bzg92LoFHKfP08gD+SHewGrNiFTFwxOZP
FoLU31SdpXNEL9XmhjXgRUXFxK8YoN52MvGd9As/zkzQZ7yJSKdnx4j9TFn28V5M
UHihC23DPOCBLfT0YEB1YdzlDyCTmhdyXhDx5V/N3VOsE6Ir4HAX8gTlDsrVM3sW
MbpHkQ5m6mAs7oHk9lVt/P1MgXe9ho9g7P4qKzaRx+CEJFdDuotedzkUEsb1KAOn
ZhojBBQqCrmh/yXXMPE2pYH4/zrTINPAkL+/jts21xiBVHhkQLy0vyKXilvqwjaV
CnacbJvSS3fotkDmAkX6TQbTocU2FMRTXOhpiLdkPElKMibQn0u6ypqHzU2KzrQd
F3C3Tn1/oJJCKi15SSXez23/hNIpTXVYS4o2RNo9WpHunC8YUWyR9R9s5uYTV+wQ
sk+6kEbV9pSAe7UujeAtZH8GJinWN0ZfFi5MOGbtG3ATdfq0vX8r7p1xzEqsu+jt
AoGC2Lnk+xikMjOj091zMx0Mn3ohsVTBJEZTQu/ooKoctI7GJME/ocOoiL5VQZ/Z
sI4O6NxfM/xlZagHJUYYmKKwCrtZDvqwrvG9EDoYPybIgin9q3VP77wB6WzMFtO0
juYE//IQU+1mgSlR7uCvVFbHTAINm77M6AmdNHKzHGzIpe1OGLJ59u10uZBBgEJB
fzeevNaK8ffQtC8OWatRGHLokLryrjSmzMOU26sD1fJDobV68Dk0nTILbSsl7aXa
mdnF/cw7vaNNivbcOdOR47PFBggtnznCDCed0d1kV9AWHHCS1pxsaOY1dFRgM0GA
KXYxfgejKwHXziIuz3rlMw3523hvy4phmIpyya5laBCjZCTgw7KCLfM/T1WUvlpd
cWxojcwO9JsiVIy4S9Hi9JCCwk7bxGQcSX/eQMLOaA9fC6KiE14FeVRLkoioWJ50
K6JsruvXH3sYzUkxLHdbgzWCNvS9SK/wulrkeso2OkQn2tUeJoFEsdQa8czInTXf
GcmqLOREwViiH23bwZ3XdwRRFw6t8/1T1Aernw6T1ncdpN9SCM0FhgYTQRGc/NgI
rhq/HY4pNLJ9V1kaMfeGzYEllnBOZgsq9gRNtWKfYJHubYXlbmW2v7ammK3XtfDy
EDDJcL2Dq0MgIATYA0xz1RVJu85c/x0X+tvALomq1o6pvLopUM549NlILnwp7qrZ
R+XX5tgR8QkbThEnq7D8cQYfqpTllw0Ok12Wdf7HvUoQtcrJmzkHuwsYBMizZ0h9
7ZR7JQ9p/2Re4uy7NyO0PaEsR0L2yDb5ZCUF1t8YBZMFt/fIXITUc+wx/CoTPAxv
94SU5TlXtcDncSZBSQAPdvyflDQ2jgNiOX82m3HjG6ucPF6lenRJVbkjV3SS6y78
X/AE2YEoK279zt2ZKqpFSHw1LUJuVehrv/On+qGHCBJGxNCb+o1m6SqsIkerorJs
3T9vwxr2itgNOO9oACqz9+Z96fMcxgqYyzCiRle12Bab/mb1Y6095kl2+Bbx4kjD
sEg6R7uVn0X6CaS/gjeot+PJGOeeFA7BeFBCCrZK4ASg2cCwmnS7gtvOai9xeIvG
PAnNhjTorPhyj0kMPc3eLhXmBW0irHoWPLavwPZYQvGbSwnjJSHBoDP99qMnna0q
3eDKn2se8f1JhOdiDSW8jTgOaIy9MErM5fCX6ahchi8Rp4nKKTbUNQ+oAtmjp4BH
okVkd1vaC0bOC8L0a46XfaOHhHd/o/26W3SdFdq3EDH3j09m8u1CEzG3BSNS+nfh
1V5hkHjqsBTNDpNB0QPAPMMRtsl+7af8Rj7aW8l53K3vO5d50qJsn2hy/MY8egOb
+fW7bRIn+nMOEKSh7iIvS1PI7zpm7zj7o+LDscJ4YitEmvA6N1ixBsNrzlfRFBRQ
AIjm8TsjkdIRWQ9/I/TB2bLMKFtFfaqXB5utc4o1n27J4sUgHGxtoMt601jJP8Ob
qXO8OhOEhAdhD4HzOhcxJJe1n4r90TutO7I/kHogu2ihpyXPWNXj4629vhR7+g0Z
LdRQnStaHLhL1m34EmRitesF+28P5WiNWivHcGMirSJy2+o1ygBNisO5DBOX/xgo
d2nCzOBT/chIXXs030gcAg3NRJPnHrE13IHumET6T4IiakPYWwg4bHUJEweSBZ7I
Jn9IMgInMeltGha8HZWDNGMdtUt6BUU22joYmDbqmDAM1jMxNShidlMEXXymNGlU
UYOZSZPIEEUWQqpaOHXsxkIJkOiYBeyw7W52uiAhlzgvstGG46UuAllG7nI84dOs
pneXGV7XKO8qXpEg2uecezltEwJ1N/u74x6KikBee+0oJzVbOoyQ1pVYfN/pdvkq
wAQpw1X6R7bcfkf6VjbXI6TkK5BOzRdbr8fdRWJoYPAeKZaEJbswhvO0AbH8Z2m5
c+gaB7GGtVCP+23zO6b3zS7qhOnfsYWAlsbQ7CrkFmqm9s5i9yzvfuSIzCw5EWXj
JWpGn6FNPG+Uh3Co5yeHjiUPOptBn1btNwTONI4yfdzpzv81PmwVR5W+yCQ+SFnG
IniStDktgaZT4BVb9rcQDnR7dVR6CHLtsB/c5ZcAfFMQ5RjbawF/EauNqSf3ZZWq
g5yn5cRhBkzE0LuJiPkYPeZDBM4YoQTqnwzECZqjmIUAFU48d9/LVejnngMY8cnS
jnETt4nrUiATo+wnhPJZBXR2q/NyMTgna7xQUIUZG+Kr+YxLW4A9uzRkQmGmD8YW
pUyvfKLpxLg452PmPyhN7zCB5IXIDrWXT2orEhl6JKSVMD2Hbm62OaIk0ZZSdLCf
t/msY9eSG76cpX6qV+BdtF1XVF/MYTtUaqhRt4wd02JNZeRjMdVT2JyEF8bI5un0
T7g7M2PsLbY8eKUbQJHoN8fkOxLvyQ/gFLWPW4pJa164em6WczKVaBIcUSVtscQ9
t9bE/VOOcre0gKT2G5Z0UWn/GA6pjn9HMLLq3zGop2K7IaU2D5DDK6/tajbtQne0
pccPWWN2EIAiYc1jr8iXcUzZ/QcBIGOTqBWIDEBpFxRIzD2+hrP2xrD9GNkz7pWj
0Iig9Z9jsWV3+gWhBNjYBFAoHPScEaR3oyOnvZuIXWjcCqFooMZkJQc/7f11OnU0
BFF0pTCYBOzqc7ZIKZtWWjmQ6iABdtir8jVQio1W7HzKoOxKRilbrQeKUbfSt4X9
nTeec4Wa5QzkvfyR7IbapbOPhFHmHVCZSr3ErS0Qmg4i3sxaEwYv6mMKDGqw2JOl
0sd1IeJJaKFc4V3sEeRA23yX0FFAU/sMbNY9mNFoOpXq2/YoShKd1hryCIn+/2By
NojBK15//0mpj66GMTXy/lu/wXljCXv7lDFBKVnnzT3PB+D61yqZqzJP6BxLCIs6
hWA3TfDSjW7+uFCV+l//GekdlYcdKSPrcvDSNBqjFLBaX2FBkptr9GdZXyjBYQhL
c7EvLB7IwBlJDEg8Ihcvu1SSNQUJV3i/xo6vuKF/OQlzGlIWeOCG0VdnYQE03BB7
BjzuXyo8uchnbvqhltgP7LSYGg9Ux3YgriIqYZCUUWsPtlZveT8x2kCuV8sJkGOs
8HKbynBFuWw7EdomC45QguRiKlwvFUg4dOxJ4/P3exPYmkC0lrFUWgcCG7DCGhmn
bLenx8x5LbtPQFWnQop91+Zv7pZeRUPQxETCR4A0AMoatroN0SMujV2ZCe9cz++4
0JSXYOszS920r1dq5s5g3SNwrlGsaS0cRqHgQ12k8n8vT4JFYj1nNT4WAIXKjEt5
9cS+V/H61vzsUSm+Qyv1gPE1EERwQ4k0LuBj6oui/Jj3AHmBc9OAn4AztHOb2uq0
wjrtISUKAqq6oQVhaTbE+VtyDr30AVp31Mx/a3W1ykhPFZUeKWr4PuhcKTVysiDC
aNwBuY9iebChbDtPkE3DqG+pxsEZbhsulf3a8k+EWVxq7M9mSgyQ0hrSU0cQotvm
napN9PiV6Z94hg1UJa7B/Y8X0uv5zy2B0UwZwBEnqeXgeP++Lu23/WdYvFjuBaij
o+OgwYBO7z7ElpjmJMsU5lS/oeqzwOY6MO/b/qIZfl7rH2y/kxubehbfd1lIVcFb
V/jgTBT+a/GkRRmAQuSknOzsSQjd8O0T6vNEJ+4R57lnTgyO8sssxmLhibE+em6c
INqoBz9dn4H3NhXTwA2xcQWhE5nVMr38bGhayvA1oPCj54cwNqCY7DK36t/or5k0
VvPd5Ok0uSSCdEMmCxJK5C0lC/8yBTLIvUhpwihMMpBCS4moTF36U0uLWzvyGJ5y
GiW7KYrL5t9tIj+rfaelVycInDZz5Bn5hb6Sj9gsZfSRMPdWj20y6Y4ULwe+y2p+
WG0DYZdQ4Z/nKEeJJL0q+xO9EAccn023jVt4ONmYQPrR98rNl/pfCuVdNbemgUiZ
fnLatFE2OM9CaPXWSNonyuHjU0vAuBm2Fu1jUCXdTQCiIkWR3SBPwmiw0rvvnnQR
fL4zvGIsAUShdlJDeS63ADouAI6cWV9uGtRIWlFQ+3TF9gkp1PT6+f+7wAztpJuh
b06giF1FSdHoz8QvjMh/i0rHqYbO1drvjNkj7uK6DLutTVoiYbtyp8ZxLNM/Gnbj
/GKBczZ+DMOqsP6/wCcjljPcCvh8PK+lQa9/0lXsPRa8+W+Fi8d+joSxF6+JV3my
LxHttYSFyQzVZp66Z01dYfAZ2d74m2KhGFcgr0hexQ0grkFm5GRVncYIf4M/PZxV
9rgIpGmU1+B6hq+tvUT14u8e5Qrtcu3pd+yA+ClgVzoBv39ddiAJzXcDmdNDDAgq
2M3D7uSMJaObm9/LQgoHPo5i2FEGzs4sCGIubZFAQ6d5aQJNVFbAbcFrUnuuZba4
+WCSR61sWd/zfdtENtN2gWP3rQ1kHCi6UdQk3nGA7T5Vg3OgSyXjCQY4cUr1M2u/
EtlP89J+zhzMgXZtXak+eac1JFNSVl4V2fN0+h9RQLIsRIjxX3tdV3fyg5VTVygg
KsfFtNfBHbZ05a27saS2Jjju8dTv3A6o/jG7DGF0aO185IzDWqoYtt6E9gvs6E9u
Dv48vYO6bOJJ0+y1GOyNW78lWAlk1j/zZDNHwNt46k7SyFQmnzKr0H4j5FR/dTqa
yEtRaJatwsEzrg30ekO+Ug==
`pragma protect end_protected
