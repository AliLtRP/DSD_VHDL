// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:38 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
KvVDe5tDupFBb8HzGRMZJkl3Zd378w6D6aDyUAHRRVgp2mFGvX9C6NKs15OcbR0z
YDaymoLkszoP98JOPdD9Plw26gvtphAS9VnqfmCW8nfh1Lr9Vrs/7TkFHiTX69R+
F6CZ3b+ij9KJ0iEciSZT1snmS9AmlM5bw1cQg+1JO0g=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 3520)
NQSHIDQbFsJ8akkrJIRMxwmsNTQoJvB6id3irrXNALARgnnSKrFLUQigeVn9bEhY
Wii9ZLlW6609icM1u/91UsCiPxFN8pBIQhqIXkISapvkt1H+w0KprAjgMXcRMZuL
6haKs5e+1nIvSJcVSR6n8z+SD/td0vY2aCZxvk45VOuRHuwOICOpUnVTTAsXX17Q
K6TajstL6scCYPoCz3Dg/OnUgenWYrsYus7m3ZO3FzyS+dygM3iyK5Um/Amr3vFe
HAAJncU2WCDZI6ulihf/h/WZ3DqTL/gl+PT6jqxGg23lgRTch8we9zhrdhko+Nz+
NQSrB1szrwWMu3Ya8QuwYB0bNkDkK5of6CMl3t7BWweBDia76/hmwCy+BCYRHRwL
NbctKauhzTMuWA9RhjXbpNioLdZe5q6CmifwPif7jr0RjcsFpvZzrx5kxo0FXL8j
A01l6chHdCN76Zj+DhlIXZf3243T/QXyHpBvZ2QIDMO751p+dCg1scoqpYDvSZZR
9uZ18qQYaWGsJMguwslYZJgml+ieN6mq6bBhXKO9gvVrbvPqG0I41moTanK/RS6v
MWclEpMKcly4Rwjqr5Z4k3Ln3Q+1jA/uq28O271OxVEN3MTQ9MQIwhYDOdQAU5NG
0jjbTv1WVVfZaCiWunxO1A2Kb9IaJnU94H9Sz9IKE7k6eN9oek+b1Omk4HDxcd5n
8Nnlo/qKA5O9TumLVGJRm3SGIjHDxQdFj0k8CfTrk62zcsFQVyd4LAOr+VV14+6l
RPo3gV/UFWEeoWb1XMK7zHtqHVZsie9R/udOzS95cJ1fY65sVKUQZQbgkdBidETn
vfTzWqG2h7lRYio5ERBZsiYygWu8wa0NAFjvVZQvjAs+TcuExpl+DaCNvVLftf4c
Rg3RCoqpjrI0HhLUXeZpVTyd2uoq4QNFuRGbgP4LSbM8j65T96DeE2wGbvFpXBZ1
UliIOaKMIZN3uLu0oibPYFqQn7XkXnJasZwxg7YJ96iWNZy8Z/1vLzDNYEORGjXR
gMNAl59X7vI65lnRK3iUKi1ok4rxLARyZcv2WaDB6CX2Mnx7I7mD7CjZ6xjV+eTB
7wj4RjF0PD12J+pnWRZVsTaftM5UIV51gf1C+8a0zML3pdQ4RN/MIFG6k653o0dp
HRnM4aqJiGQdXl3eGP6FeUYL1W3stP8+XdYJPbU7HDM4j7jZ8tfBRkOdA4oRJ7hZ
OgydQfpY8PaFI5mFhgwrzsRIjOrtJdI8OeH2+XrBlgqbvSv4/kzpGjYHtU5BZ9Lu
sWgeVGUn6kRySdeDrG0VAUhzd8c+OroKXspn5GZKGzo7q1YyNuASHOuoColPiJfm
8iWC0un7bryi7HRL2jNEBeh2Cq//ikKZayTQiwGzJdcvDUnyRkyzy1b9fK6j5RyZ
bGmvnvY55zz9d4Ifp7KMT7KwYtoPzmrNX7opIxsgBZb/O7coUCaWApbgZTgxMbcd
nMXlsJXATZa4PuffwmqncaIaYmyX3OqAeJM1TzFanEXivQ+C6F+wVBW9hSRb7nNK
AxOjMND90q6Ewy68xoUlwfkcYe3V3qb8E1iPtr58XD66C+K1ACWZLPXPUqOEUvp3
0lgf70nWIFhTz5xlciZeXjpyEqWaigvHurMvq6BtnTRB6czOlLpKZZD5nAifMc85
E8Npggjg7laGEgxmbuVNVfm6UkXyvQq0WoJX8yNh2y8faryw/kBlujP1mpVlzxyG
tjRDj8TIxOcclFbPR5tS1kmTeCTh/5WMv+OMRIPAfBOyMdxOwQeOxd/hM2bhSap8
l5gx+eutJuUMzCzsPmDqF0WXEGY90n+2JlST1/pIrmRuLXNtRrjwrlDMpF4QaMAn
aVOrYTN19T3+eJNoIJrkmPvXF1ggbBOhfwUn6eff1keJ4UXnqg0Jp2LkHPK+PrN9
656tJP6fkB3nVGW/rYo7mp/t43NW6lZJLGYDjSeZyFDVm3wU5IUem1Ph2rwZlZ+C
Htb2Pe32v4Ty7W1vazIlTN82muqR1/jKMNZCAUaMQiUWj5Soa3R0ruARHVrnMq4t
3nFMQQLo5N52n773t4237BmD6D+PVUlq4rDShvo5ETEr0iykL7wvaLPBMSUDBOLL
YlpNUSKziaK2QoQZrD9AatrVwG2P5sjpLjxPeMBZlh5RsLyu9ydwkYTAihlOf1KT
iJHP8axMR18Tr6GX+oIhOATXV66zxu+vAJarcMdc259+uBeVuhM+sUInJp5hMMDr
hZ0zmJ8VjkoykjXPI3bI16SLzJyZYyLeO6tdAdJqiBjtqVzDvskB1v+xvhdEIpI7
MfHlWSrBwyAktNW/6StWgdA9PeAzSVktGgISUrvNV/XAbSNK7tvdah93SFXuvIsj
HYi4xgc6NzskxaOvn2EwGxiaeIF+L63suuEdE0UgS/vDYI5iBesmjNQM60rCtA+e
Pq1rQGr2fhpQ1QCv/u3VDwV8Tjxlk8lBSL656qPvviFPIrdPWiF3lLLubhvsD+bh
ErWKNavBSEaYXAKuPsdqMGMaIROd7GaJNuhn63b5KxyIgk5l76lFjK4KAw797Uvo
vOsBlykwXt7vouhDZssiHBEcU9wd8TSdEBtMCuR2sJDNXuBM90Osq43jgiGmkPeS
C5LtM6c1xjirlmOUqYDSQsEQ5w1ZjUnYxPRCEm1Z3JeZL/LitFYUXnha/Kd/+nOA
/gSfYRcTfN9KPEaJzBpk15bjhel3HuFY0ze86ficULnJAhGr7qSBel3qbcWLSjOI
nL3aiOPKFOVgLul40KLUCpQMDS6rPGtZxNAeGMbluIptLqUv7U+hAq3G+TnFc5lH
87BnoaKXGKdVwiYwZAXJG/GqvpAb+29CIZqxN4XGXpUzCTTZFYeSEsxgTU4tFIQt
myCpGDhlBDWEaSN7uHvW9dYmA2ZL90EbcWJucdRpZ8D3onoy2wFaPNqTshx2p70F
WRoh33yk1HOtzWem5NmZnAGxoOZCOAR2aHeEN4JJKkK7qT269cDm2tIqdKaBQwFm
pP3EDVEUTBbRX3wxKjkBdIje2v85GRZPizMkaiOlFiehN1WpraUU3+y4b5g19VH5
yXZN2DNAptgrgGu3UyHqmCXXcwxRUwnhbTEy5tmAKbhx0ucFsZGoBBJFHgidOLcH
t7uQpQR1hz3s5e7UNWqEP6vooVMPiL+3EMYUVt/k6Mkd6VzScqQyafmfIaAXyAHg
lPnBFmq0kxvwo2HVQmhTKpIs/TLClfkG+n4LZI5d/o1vkXLMqF+T8z2uQh2OccVm
X5LS0AWZhfFZxPDRrzPVPKaRBS7h0e0BV/+OBw3OmtXnWO+hFfYU2Oc6ygYUPBc0
a3I0xKy36xXVAqoOx1UubA8RpB4ReUA1XnRBAGGA4a8b17hKeefkVwRvHbExMRGy
9tHJDRSMcRXxq2zDuMiwCfoRI7JFm4h6YJV3Mi5eGMIT0kc7JYHiVAzcq203yiGW
Rlfk+Y4lZz/CqFLLC+Mfa1DPKojj8t7gNPvTC0DSe7KTotY4SAZIP5XzNe5311mi
50BMpqFWFN09fYA2H2OOmNEtWfmzEBXxcvlA6ka0Ea5xnv4zBM1TackoVwSjejmD
dmgd7GzZnmt22Ii64js/tn8gBjYEbhP+UuRY2qADxQmKWE8nSBd3i/B34dqT0Rhb
Ig32Yfj9lV3FcH3XZpBPglyU9/5Az8hL+Jgq8G2vPpKWsfO8isaN+ixrrN10syIl
DVP279Z3i2nnpkqO2gf8+LKerTmdakKpklBDDzyrc35yzO0FnFJSyuxx/PRu3/xJ
l0sCl1Xb0XLJylMmKt7WY0JYrLv80M/XVOHdvmlIYSxayTFqDoCFXM7rWVUvMPXn
vzw3TT20UOeCIYX4KhZyjAEuDx5aIDlwm3f/I6Aech3A/7vHXo6iqdzulMV6oj1Q
a4DKUHVbGwixFzjtx4hRgQ0WTNnW2n2DYOchi/WFYZo1JL9VkyTxfm3pcFkcjn64
isfi2C+DPrK0DmPCeIjP+wF9NyGvpW07MT5SahHFYFw1jBjcaPzrO4GdhIaBmLs8
qYALwaIm+C5m1yQN8az+sPkYWFm5ZLdgzP10fn23gUpgrrplB/lt5iDNVIGMhqlh
tE1iD8YdXZuXr89nW8uHLSePvrBRwPNAhnfWw0z6O9rcggV05cLy2BzW/dxkd//v
YKj8gsmi6MNiACA/urz+cc9EWhriUP9cSsEXYrXuNlGyN6Dr0kTUHCrgGz2JdbgA
HDDVol+nWITy9JmNez2CadNyrk3jmOadxt1esTA/4JKvYPUpSYHUX0N5LPTt2+By
Fjao2yVclX5RvYePz32KHa16peNMLrJjxMW0aHU870uzKV4m6Ek5fbCqzCDQv1GO
60xDrTYBf4yZGvP5Km00yqaIHQugzvBIL6bYgObllfh0Or0kbBXPtFnCP6AZa4uW
wcSrM7JRMrT79jddr21cQ0u+RkuRO8QUnS/0HrmudK51W9r5/EjtmNaRqGEGmH6/
G4DpERJMUdUL6o/Om5r7u4OxlfNeWO5W5xF6uNgWiW865DOWTwiW8+BuE8TFDbFI
ebKwkvhHzEOYLJTM7YXXpjegc2lOzvNebbSo336lRy/QiDaNsu/UXk+EQYH/WHJG
SvlocjZcbb7kRuLrAPD6MlOWqA8PywYV8jC8OXTev2hdj48YlTeghWjm4LBQkpxR
Cv8lc6E60WyAV0lN2hDHGQ==
`pragma protect end_protected
