// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:49 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
teVAgFRjTaAAsc7KDd1LBBhy+xsJBD0TKQfguAX0kLS89XTvWDm2Fz1CcCgFucFv
I9aEhVGVmd9+skG4WTvnAbtSs/5QhoKWcY53voHtbgZ12qP0bhqapLB2tTmbsrLC
HNeuvONQlydIbhTZbY0Xo9Rp/oW8Ug843a8Lb9f7HYA=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 29040)
28Sc7PW+ol0J93vwDJ9tfUOVjUmFi01q3wRFUnY+0wLYXA1ccSJf95rmwlwogiF4
gSnxBM7d7/gFw+CX9YVPLu0YQYbJ8ZODQgeIhudRalMNkWyFkDsFsOHceJFMIQSa
XMk4WBlLWZu5c3zvFRb3fysDyxJ36Sh8Bk8htkftwpOfMwaWDDwYafgSPjd02hnM
31uNlszITD14LalcBrsKc2v7NEsdq2mEKzMc08aAOLs2HhrOkKoyl5OZhV/1ldki
c9XaY1Dlr+6Ay5KGDKSlHBsDXf790r/3HJTxsmDG9ug9inwp5oc8U4R3VgQI4dd5
v5Lsxx542iCjc9yF4tNwoI5k6HooZ7hvqf7pTXeMiqww2HJspva2iClwgJe614AQ
VXRlvv4tGkDCRtYgLcCNXYc6WUH8K5U5zDkWWtLTxSkofKukYu8z8FMg3P5+2+ux
HTkrLI1Sgms53PEcvcymHlmfWn8uWXC8wg3qE0fBrGs/+uNAHIb7LAswVrLltGKY
djuOwl5fxoQo7MSHBMp4ancASdIHxMzuGWwfQHzlIO4R1YmQjNpY7BvFz79TEPjJ
UR3GziV0r8yEabcpMTVz9bPhHiMhPmlgcWWJJXaoljHt8/cM3vaSpDOATBt20MDU
pGWEKV1f7PJiUtFWcq7qj9ZpTbF4SUNwI9X1xcwE2TLbtBpeSkDjfj39eGwQNldv
01weKlj7X9G0KYqVmOrl1AJxAC5rXsds4Z4+b9trP/22BvmG8+XDg3wneXT7oGlI
gSHzltZ7hnNmU10mby64YvWaq7X0kz7rpLV/TlJp4Ub6Bi7AM9i9x6Bav4MN99Aa
yXpidvkzXTiZPfcjqNSqH8oVKcCXRbzM7oyrGesmtcMR7fll3g4WqB7L4G3Pxp/d
SjvTtJsXjcp+OfM0if/1bVhy/YA4fmLRlXh2mGiRe6ZhBxGNvf2/YBJdwrhpcWRT
Pp736G2owDY8pFLs1xfo4rEqSGbrdNU7GRKe9dcmjuMB24gtp93+/NaY501qqFu+
XDLwQmrtfMed+vYn0RZO6ArhBK2gYjxXkBv16IY38S2jsVJCpsMAXDKjTLhdTWVk
pQHRmCJNNm9eP0eEcxUlUrXhyS6SOBm88mmxLNciqSGJzO9lmcSS4PtpyxNacvEG
nRIZ3Uz7jyP3ku/5nwF/lJJzWaDTB+YQfSPEn8L5ZgQALXz26/aSTSb/16mt/TR+
o641UhqSV6/tX7vbhLBNRwFPttq0vpi2sCwzGUct9LunOHTiuD3ufA/xWjcm4zbs
ABGKsrKYvHrV7TXVPl8zzf4oubt3WZb3OaOXIdRFV9HK9/jF/HcUrrDqO7hMwlt6
sy5PaZbUa5B/D2fEVxdD95xME+h4NwIOoe/dKVoBKhyqrm0MhIldukIk+T2rYmnz
yaQ1Ddgz/9XDduHx9wkGfhBf0i0JcdHWpm63EmwHEmPhbTuaHKQy0mdd8KN3PkbA
uuVuLwyRDYiHpXvTDkVY2g8H4eu4nvMwA0WGQOyBtA99d9KckYTy6ENPve+2KTeX
2xV99AU2nbjrggOB4T5rybit3wJg6A0T4gG7lXEdxSs5h3jFOiolYBpDxvaxZfnG
3cjlRQRTk26Ib33N/fxtpz4AGZ1WuFQx4+/ZTmpxAM3UUa4ACvn0HMLH4sJUdpes
YroNdGUqslkfV2ARNx6KX1vrbKG3gsuad9SO+GollkusqCPsaaBe6flN9NXRKkTG
pQHwI2yAH/my8Vx5id6DfPW8PyYSLRruK7weVmxlbDSPi+tEl6wVtCYtjjv76DzF
WSYhZSHAe3hiOcNfmVTmoAHtrpTbgwAfOE5OzvG7ZE7chYKNKyim36F3o798fnP4
4LcXyhx1Pl+n79my0P7d6NM/g/Z/odDyoqgxw3M9i5yt61lyctaACyVAduf+qbPP
+WrWhtuz82gDDJ4yb4x3MV7xvMSfSa/JjZEvCfkrBpno42N2P2L7zr+bsXIPfUnT
OG/byfzMkTgK4im6ucS9E2xGTNShsBST0LpXz4Lue9IksqhLtGpGdw4TQeiB8oWj
aV7hzMRXxIoT4VVukVQa4E4b68wj4aUP0KRrKTlebO5COvs//KewhknoXzjdIrB8
S0rCPO/aGABGDWvDEy4Vn0oNwbxp+9S2tRSFPGzaKvi74hAHha/cqrOpu3Lw7Yz0
PhjSKa/9c3Y1RfFbG9OjzNmRPIZxSYOEv2lWWWPdAMc+3icOGj0rThTn0/IVnRiD
lXabsZeuriA97bMP6y6ijq9xuyLYx30tXnRGpnsbzNQo0/lPpb+MXdKk11JIaN1s
ZZ4GjK0e8dfZDm6eHik8z3EfuZ60o679XZWGVGpX6dnwrH23G+ZOrol07DCy2VV3
EkUjRf6+5aaHobMmwJvK8O0/aLugCN9XvrR2tfgW7/GzCDpaDHTV6mtCSkW6GcFm
fWCaQz59fLYV1q1A43b3lJp4Ds69EtcDFvqU8UWE5dAq2FcFrCnY+kFrwz+Awylh
K6qWM+iZ9dnJKV8ig6sMzM10N435dl8pcQ4A6S16K8lRzjxwjgJohXSd7T+Zmnxj
2l6TeuSid4Lpdrq3hvMgdqqmQ00I2XwAggrGrVAHJu1mRpYM8PsArDrMOl5FfWBy
fOz24p3GUGdKvs7G5SSQVecSA/RREbGOGJMTrfBvP85I8cJBo63Twi2x3VZdVuzl
KsvQ2nf8JTgqAr4MSolJ1NQCrdenE7SNxxZo0lFmz/PSF83DVap1HTMEbxrf2pIN
Ym374iCjlttAFzcrCE7CHxtkaeta+g1FiVrUsQilI4qu0CwBiZK357L5GiC1n1sl
z5Z50DN1Y7UG/sOzUNDxMk7wLiqmZdrF/tepAtghXgE0t1eGszeVO8KuV/4W15CY
tPJLkExTFVK5m3l9WGcBmebkPVeNg5l8DlbvFuVI2bhcJHCDiowWt2L3eHY5ij2o
GEKw6KPS0wUKZI7U3YfVF7eZLGLIs/ynoidHYwhnp3p7+HJgBE0TAC2MnWmtmJOv
8ERTE8WkYZzpQmX32plzlLWS4UnVGk4075rqy2unJYiBNnXk9H37W8zDz7PCtKRM
EjRccJ/kOfAgdNxKMJXbQnimV4jKKqr+4fEAS8ufVtK7WluYhdn6ymDVvQuUDoEN
BGD4EUKShHrEdDRXwGxd8Vprtk4eqSf62M/vayNwma9eFNm15CXX8j5OX77efNS6
DUVl1916LT7jes8XZUuGS7lS4/lC+3pSSm9V94ouWZN/AWuMuVlZpmnjqGM1t0sG
VOOLwFnSNVypzKiWBZ58hxyv/vCNSNWlhnJ2hZcLFRrdvj5EGGvUxbVDcXV6L5KG
cuKt+hoP48Nz3WvW1YqJS6IgB4TnYyw4t69+OdtOwLWzL9Z+URj23e8JMTuEI9N0
8Nf+6J/GJZUCXqsGGdD+CWZ1iOx8WBtX+ttmO6klUa4tzYOnStTtBB2ZssvYlkMk
OBTroSrJeKqEm4K9o0irJyvK2DAVUtquZlq8TcyD+A5kymet1cERpIn+QTuvu8nK
GLsK25kcL7Z6W0ordDJyxXF7y7OqQHnJzoK9xeW4WS6eiuhXugrblThDd2fbkScT
OwOY27b9ICYy89ks6Dc9MkhRzePppWKl2uRRLKGBy+ctK7rkldO8LSsyEn2YzSeA
g9fxfG+AWW6O5VP1Bq6lPg1o9GYDTAZzdYvnVNvFwcV+RHnCM80fb6FCNGGPGhh+
rQ3YyDx/ij8OD/sKc8vU5w4rmI6iqgD4z4OEe4kMY141duslQLMoF0fpYfpAlzho
NYtn8C6ATVB2z/diAqCLPP20+RUaW0sDQpGVZCPKpNaI1ZZwpUV0Ao/RcEZn1Jny
WNuBvM8s/zdEd39O9tlOymn5yFq6t5a/8KMzmMemipjPzjywFkMy5mSz4D2/wAmd
DkPh1wXgJVFDeQRwt/QRGXADknGA7lQYqx0bmrww9i5S4NYAs0FmqK//Jiqc3RjH
o04i5Ry7zDd+2RPhiUuLQPT+rh0/EMmlN8bGWuN8OuQL+hc5GtCqFW7c6vq17DTR
5zyttW/9F/hTF4YD4pAgotGtrLnoNbnE8w21JYkiv4F+Feu+aJ9l/Ebu2StpNi2Q
yJEEY3DHrW2yoX+lbe0xkVi5P7XuRg0+TpIeW/9VdcxmVYWLmaU924GNVqpji1gg
Fv4MkWwKuV87GsBZhJqC0H6i7NrV6kDvY3GEgK2vyIKyo5tN/lz70BWdY4uiQXOK
VCOdFZ00+RTasH2l//BUEYDEqH3KCC14YoQAzFs78Z83Z0h+hC/QwIxdunTv0Wpo
kUGtZ/TOEs6hL9DwAHM7K8PuAgBO6KEmKvrHXse+V3ACK1xos3e4FuffwjUhbDnH
fyIiRZdrqdKCZ8SX9IsO8IYx8zlgIQ2BuCULigCJQFHaXLhHlnd/JbdX9mPxcuvM
oVTAhRRKZJaVfY/DQs55Gis8NjuiBqrvtJTUGo9S5BQf9U3nDH0ppS7k+8ZDt6yx
+fYljc+k6Zk045GUSzGSBEyBz2ccnCcpvtPVOmSX/IzkUjRle+/zwrUhUrsthh+/
FNmtqBK5vwvrkStW8osn006XkwJVW6KM3+Mn4YY8URgviZxHsUo15nCTTQiIhVkv
1yjp7akqM6AweQHv3gW4Rm6DH8BUFCc6eA6eBe/i8qkp3JC8bTwecj4rymCM6gnY
pp8+SueMuHQeFiO3qGOe+QKb8b4uOBAggopC1FqcXOULFbR4O559YW5J28hV1gWT
yGuC5D29CRZsEVNxBGS8Dhqfpr4smeHNevDxxalzcV5YHg5tqjbWRA7RWHhUHyTe
KSiv/58jBFrEMM5kNHVBVixlkk7F6+iEhfRVRGg8LG7hWS0cQ/bvTRem+D5bhAYu
r+3JKyTA/9FAaR3YRGIJ7EcnhD9ofPYrBHvuRk9Qt1h98JOLxw772X4sC6fpcVOo
cl3qgm5tC+uJuUpCz+KrP90ZTaiiKSD4onPbuVEMJ1dUGZvK5x0VhFegEdd8ZblP
OLXa5QTw4VZ6HijoVmufCcrZ0vKpINn2bZxaMk5/YtokD3z6XLtHDLE9LjSYjPkP
eydGeWnba+W29j/y326BQBeO25Lc03XBKWwBngJ52KCqp4v6aMpHCInte+2usk4D
VpAC4Inea0MGfe4dbDMbpCBXDvAqm7M6ojJyN2r+4NjGVfbXWGgvARzJWOhpCx14
wy0Lx4NTVjQrC7IR6LjuOGjPSlcSQrIh0M+vld9/Db3lkqXAFuJfKPogYMpZRPom
ucmermf8NTXtkPRAMK2Hjrc9hEHZpgJChVTg7tEjXUKusfBCW+3qHzQ+ICYPkK7m
zO0pWUeQq3YCkE9Ju+tQa9HGKLXbLCtxV/vngQp4nWutQSoPM7/Hxu+4T5KbvxC7
KHZ5alQIv5FnjX0DLpT0zUjFn117A5CJUOY3mF6yz4zEyOyzDJgNhMap7tyOnSoY
QI9hGuorInWdFJyBB7k5nDN50AWgRL2UyNak1XaMHBjwI1iGUqgOR8t18LhH74IH
w0GjIx+TrnWeOSB30HOgTkdQoMuXSfKi9N+YlOUjTJWVkjqjNsWV4enWAwc4/1oQ
p5c3wq1soE5MOVrY8xGaYLGTv27ZqKCWxnOxtsu/CJNqa73K5VbxHehJOJrKPMr3
yP6ixYCDXPp7d9NjrQwef7Q0bx1KSUdtj/ZNwNDjbhRN/SlYDy5VhJPj8iIGVFF1
DjIWPRBEiaksl/tuukh08ZtRP0I9W5saOWZxOpkk2TqxMRQhuNPT5EvCIPeeRsLt
mLyOdKOoweK1cTxmeH/K8DrKskJvN8cT1NsOYtQh54jjHk+WewYcHR9LcNqvHYFW
PyucfVaY2BJ+ziavNt/zkrCvn0dBSZbq88BLkhr582vu7230juALOqBiNWd2tubM
Y0J24hQzRLzP6++tjJ3OhybHp7qpdScZCBB843UTY7283Z0PgveRgOFj9RTCk6Wp
lu5CeCFkTQhdOM2UZlDQ6xpvqtRyA7iQAnQpN1+Z+vt2f5EMDIYLotcxbQzOzize
WqWLx4YkGn4DITvgXX1+mAsBZvmgDrBDbzk3I0zJSPHnt40JVvYaXAfUXhXBLinv
mgQJC5r+Lr050Z6nTA4Tt3cnV7ht3tiBePK2pPInHAV5Q9gH/dZTIHoSoZoI8ta9
UaNj2flAqL8kFhyf7iTptCOsxmtmMVXTnLgK4Ddx9VZJ6tgw+FlPCFfnHuJX2OK9
qW595nDfVKHBfVrBzn51VNn86nkfn7B+PpTppVHFcniABD7LyTQqJMbsjHIdl9ta
42bGZ3sj0WYvlt7ZXlPOF9b5IZKlkh2q4OI3vpykOgN6+nSUWIcnpO5ULXl/LLk8
GlDGiZV+16+U2kdYWgKT1Ezj8epoAKvhQnsBY87JDH8Mk7BEjVNwYoVHX/DehrGf
1OFaZrUo+6Ue6hlrt301eaezgNj2U9qjXiSUdTr0qnn7rRNtxruE7Y6Uk7J2wWxc
i9rqr8yaqEg+fzBZGV31GNqHPTG0OZON9ATw3m3mQh4ucvKEsqNB6zLLBrxnc0Xy
Q9QDzVesNFG7Dd4VHZ5SBAd7CFIFUf8QgbAX8g7rgNHp/a9W3J5t6o6clavxM2r+
XPGnVWsDmjbNtu70z6jaE1xoAcdZValPPBT7rcAoFfAlJKQI9pySjTXhDtuV42Yn
WV+IUrfEBxekWlwLOiFtpwJ242RA8ckTj/sK1nPIx4zBvWhkFbuzd8l3rs5rbD1i
feD3Z/whwYgwx3rvTAg6Kg02EFMxa4FFARnZrLNLrvT97pLI8sUwx+3vi16rYT8Y
Aj02RXO57D5qvJdmBW+dv6KY+BnnGURFvWeF4WYj5XDSMgIrBxYEjgOIgGZ7BFeJ
AdO2/iZYceiVcpN0pRRTzMqe4874gMqXvTjpqbsXLBLnxe/noPpAQX7iw3iqJCIK
OA7Vu8ItfO7JKU2TPmD/zbCGEZjA3/rkNRjxNcKtUoC66e5diSAyQg1RPncWabjZ
TsKAK0XZWDktqIMdNlWa5ZhJ+CsjSw9w4/pLLtfyYKOYQWl0+97/+KUyRhWjrgQl
tzXGBwAy3r/TbDtw/LjEpk3DO3uCj4jDSWOP8VetEccTJBs8dnWm+L6bSh0p5GnM
sMs5i4vVHJjW4VvPFKvjDPPaG4RTJc5i0yrjNtwwITc0lm+r9IHyIhnoXiRu/2bY
WVyn6x5uZFLynllX45kiP/gp4NjJy5I3aV5owdWbOeaIiN0rgik+p6CkuRTLUpfo
i6AgUQPPI3OHX5gjkHbpZw7tQavyKKPdATmJvi/V9ay99oYJBrUyZ3pI125rOekA
6ltmHMi7bWzlFt3oLvnfGDdqmlUZFolgtm0/J8qs3vAYKhWLigXBHz0yw0jE7xHR
zqweSFSRiSChGfhpyI0k/hiRtoMWHMR36sRC0UlVcRUAhMvpEGZ/l3Hu8zApl0td
LztqY/r3mr1zE7Kg5ERx4I7TK7JGJK+EA6tCd9NXp/xJtpV9EHxISlajRSkX3GcT
DwB0oSOTBAUVs74ZL3tngGYbaqadUAf73m2POjduAMfjjqs+xn+2F1kj+sIP2Y8Q
UHu1DeR6spiQ0iGTbNDyF9knelWZi+RMhz8byuc75OwBDk+W5YPbfv1rnoBbafpB
tNi/XNlg301luJC/Cw/kzPZePY68GetXPRN2W83Hdn181j+ciavun9YtgQhf4LIR
PfvRe2cMqBOaXPvyCaxG4s7KC/uly/vr37FBF8qsr+wGQHXxOWWZd5bZKWR131tc
ddTVrgeOGRHsceLkRlRC0OeJKg5TdI2OJ2IhUBl3K32h//4e+6EoxafZP+fyWKis
7kW/jMOMo7mfEcLuAf44jj+sV63jRxf9Hjm1jXNlm2lfkThVPFjcmVvKnQlxBv4E
HFZf7OqGt812yg30ZaSgBf7Awj7n4/dk9MWXL6ILePxRqxhxHR6ial2fVQy/N3fh
hQSnt9vBfGTDVOf6OaoyCfGbE4ndVBqkqU7SbUfzSz36/CcM+zz/I5miw1+UMA9w
UqDdlBGBebu/nSie8PTrDi26lMTtx44vYPn35BLlqNF3LRPrzuO1ud2U3bR9pg20
KEFaq5cyvVmFIlxNNhE6uXr8IPvcfaJaFqVQaktzQSc1sFtvRNY0VbgE9jd8dRcw
jP+p9mDy13gm9M7Hl8Qd8+05GCAMySe5zyo2mKehEN+vee9kjhLgiHT10GaXebUb
rqhIZ9Yi9QvF+PS4wFdcV3MTTtWQGvCSL5IpSHEPDiqY4YGT3kdGusF2wreoPkbd
I0HkqdYj2R4sKuV2bNvhUEl1sPYZO5s/7B4uc8haJZtCrDv8d0p37XXzFMcXjwTc
8obARbEBVReIMmWoooKsTT8tT/71SZhjU21/cMhasvtXzL6Jl75nYdclVho2P3Y1
KYytPBqRGBMHxQuptHMjGAqZjaCONTPrAvDEytLINJwY55Wfr5zCEsdoSsWs6438
HNrHveez+Hv4SvyALdUtetDOZsaxLVJIDw2vLSncJxAfOu6cQ1Ja1SXm+p+wlyb7
mdlzKQaUgOgK8gn++MO2F7hDRvqvkG0fs6lELapg8lqhQKy6fR7hgEczrvA1WNv1
/Egtdq7z89eUCBWhM6mgHF9iT7ZpvU56d7Z3hLfAebj2DxRLatym9hQg+lfsEw+g
h0V7QslxfPaPdspUkmJ9Z1I5huJZNOzlZhuKxx4rt3EYvdxbfl5sUk6q5xaP9JBQ
+fjzjMaIJe2A0rDq9+znP2urCrcgyoiIK+sWnGuYDX6FeTJkO4fJQrtT9wL2UHYG
omtSy3Q6Cnxw84aGSrUdjH2l4IhiTiAIDmVl71pSNV9EJueZaB7uv1gylXQy+3GJ
eGj3xjVnYQ14Knq6/tN8yfl4uxJ3qc8dRsNnZxZ18wLopSmMpKwV8s3CukHBPSz0
HtoggTN1paTz2ARgnMwuyIdZ7Bug8VMH2ZbhZEutt9WdA2ln3C9k7DnhO/M8zJMa
9yoJqJUb59XMnK4zErT7ipNI5qzsTMx1eSkJJXA31/EPIQsgz1QS3E+5eHlpUdBP
bK+fhUhRBi53iVLJ2to9p9SInzXKuVQw7f6w8FLZnfiZvMLhczFzllDw1GxZvW3J
mLxrf6JH9s0xEh/5aRgsHeZ3Qjx4zN9Z5zby/623SD03oH1t4UHlnfdrtCghKsrZ
Fij7X+qEd379MnrVlwySgwxo/ZfSfxXviqYn5EgQw3mQ1qufgq7Br/wVbbtz4gkf
qnQChgJMb6aoXU9qGdLFeIL/Qzgvdy+ccf1yBWjFKtjQjyiKeMmSOf1fPV0J2zzT
W/Cyb6PNuiv2DO+R+44UREUsJbQwGHDA45alD0+BkP/V51MjI2TfzQM8zoEKWUZJ
CdHP+hwS6LW9kvdfSXbKxd22JqQ1uviPEojxEuoCeAzrCylEW+qca8Pyn9GduDQi
VUd8J153s9ewGy3ocu14zACBW2rDA2HhbvCZOoaZubatkhSzyG3//VnKZodOZ1o3
tQeAnYpKA051CDHjJ+xpCx3Nw5r1hXmYTUKkCFt3fHtHlLI7qkkxjIdbXBaRFgK1
FpXJEzVUOkBwHu3SiVV2R2GazrYTZgsp0u55FjpoNkOVN/+itvCUyl77YaBLa0vJ
OLvuAsvNbqyHCxpL4zzzq5zXf1e+jkUNZ0ECim9y2IGT+/V/8tY1PIQHeghekpQA
hJ1ZTDayKQsxTUUHd1nFvxHeQTKL64w77qb/YLwDDa90R9HpHVQklMGlrZ+erV9Y
6qUcHvV1DTw5q0MR7+h9guU0lQqNAn6vX2AhhMpsK0gaMhyyjyNb+3dyK4bx/k94
tHzmROivkdI7ps+NXi/0QRBVYsJJQ1uPh7evDuP5Uy38clrG9bIrmDkj2wlgB3sO
3QtGzjnGC+DOLJQfHusvr7DEUNTmZlo0giK1UrShokCeC2juPTyQdq7DSc0N55AH
N9tjXJqyt7R8BACCst/M5lYxTuOQRzKe8cLXKa3jXw111Pfc7k5r4LxPV/JRxjhv
oWcJwvSXMtIUB6JilOrUw3T9XUfLZl13JuRouw5z52oeIpqkiuA5KqbPXWSTaUfq
UjmR85OtjHSumUL+tw01qaTo1uxUpLt9BYlH/o4A+fdztYNAQS4RcwCeqH/VEdIk
Lw+BbNp32Pqxmek+1JXQC3kdPJmx2ZH/hM+AyxSrQxYUoNPYD94JVTsVsTU03mkE
3+avsZc7L5jXqY7mSYd4Eg4G56c7ISiFlwbInuA9qzdhH+9/fnBd6L/f7vESNv69
TXIqvYpftorf2WWAmfmKc63psr5yzfqahdPmB8UVNc/O4uVFtxjizDAROmWKJXR9
CV/Is9mfarevlml3S6OtI6Q5Aj0zGztM/eSnrkqTxMbDw72MCROPy/4h9ixY/E4c
4V0RDhPBFrSA7r0j6YvrKEn7Xsub/1p28u/490SH0H81OohBCPlMneub95Z9RBkz
3EeHdd0gjBAclj3NC4zJQ/tBd1gTzz/MENl3VugdJAvMVLZymqrcu3u3wZG1oZq6
k4R66EMuq9GsIEcFWBMR9RJMpkiIb60b8W8nHYtGo1hbp/4oXzM7eQDootsy7jT/
RncnuOefMu5+j09by6xsI6uNp1gvoAczH4u03lBJJNwRYJt3zt36xOeIMKfN15Ix
sjyY5VRGLdzxeNRv5FzjQZb0DjhljX6v4W8OrX8uvfgf+corWKzSuRrqXoLl/+iB
rQhitGbIACKiYrqfvovvLUefBQ4+JsnWqY0VAW4pwdfzuBKSK2npLCJEBCHAm0d9
w/erWZqutZOZHfkdeE4pWxG7sPta8N6WMPYSQvcT1vtgsNuobo9xufhNJxgG1yPB
5SOH/wvjKG/LUH+C+oPIGc8T1lQCqslQ6ASEzZUpcty7AUNSz8X/3wuyWu4itcY/
G4/yKLwEttyphqjMPdWUaJU37S6CQ/OaCZGR2H5ks+qaEe66fC+8AfAomuYb+lMm
Rz/NIPc365ZT7S3mDPwYiwizArEchE6b2QamiHvxRK3TGIKIPZsSzCYWTXiKTJwM
XIhrR64yFMz71f0tDXuEb0U9E1v3fN8RrnaCDuP8JtM9YdS+dY+yiQN96QP7ozYC
AkZIJChpyBZU+NEjBGpty4ciPXGq4V013T6olzqIqnr7429CyAJxazklEBaVb6TB
nwqKs8g+TaWFc4o313fQ0RAAYKb9YzZVqn6eFR7gKBMiq9jJSETuFP+RDzUD3rli
GUbTocg4tlOY13gRvWlOUBtGqRnq+qR/cb+RZITjU2GIWiTX25NDHM20jI7euYIW
hDCu4Pis1vC5uo9/8hNyDfiJRj5QClAnNpk/KkZSOryxSkojL6MLw4QwmPnTzcIl
XLFgpGOBqWzyATOikjCBSZuGYb3rw4uVdvqXsDK1UBmM5VgZIoE28lT8MjPgbry2
3hAtxbX2guf4hP7AnQALKKYhthIHLMVxDfCW5/hFh0VQaKIVjQjTnD03F+nL4nc+
sWwM2Rm0cFeoUJy1xpgVff/CUApJndDqrDtKgONQijctJQxVgwTf6h3ZI5NCdpXu
4zfWRENfoBTTsO+DlWVJSRet/gHsZ6JeUPaJqVs5UuPoandXwNn9dSzOr3uGLo0j
WdXXhWiGab7Wf//fZ/E/ccFg11yjNMbgbHCgN7hoRU5h8RIziQrnO5gUQuPP8b8V
KKgEo2xnDQcNjyurDjWAvQxt6DcoxmNkCDOUoVahoYGLUCQk4WyK+DerPrcagdYc
fPZXZJ2XTmB8O3UCAWjv1AJFSS9xtBa4uWs9Tx1pRvHk2vT2pRG85HYPL+uSQ7GI
+XwKHFqtg9jgCmJgQTkwJD9FZlOSAoPy5DnyEMIGlhw0oNRV4/DK8WAv/wvNhLpp
dSB9SJJpCxegSTRKOAdu4hwZHz9bi3Oje2qGSS49HVklctc73JF9oG6QgcSFr7Qy
NMie8kssuwLO2ZF1zPNpsRIbFtxJu6I7WdPprPNS0PdR7nWpFZT80niFTLSx1WeB
W00sERLpIjB2PapBv0Edgo8gn5i59kjdyhTxsdufIDv0hK+/xs1mxH077HW+nTdb
wyuVrWo4gLMX2Ds0QuUjr0v6eXH1z1r8tTS6a1t+AoDdufhFzIlSkJYQbIec5YPp
IQPSdlphIhiOBm9lpyd6IwoL3TOWoeyHnQfS6VQD1sswcREPtZMlcJkUEitm8Ahh
tEL6D6ng7rq8HVgnTjGTKJR1a1k5wkNEAhZnGq77bdEvKEzYBTfm5atOhMYTf5rJ
/ENyQoM89BPxUW72raGGrE8skjPf1HY5SBaWEXPRwEustUmco7J0WSMbHQd8kj19
UKcdnByqy2HfuEhvMEqJO9+wH8Csu2V8/rJTkd0kCIzecbNp1poTSlh9fvdXlNCX
7AXp8deNTaCbSXeYQuATICy9QdNhrq1HTxD8a0MzIJzzfKomlsApMZI9Eio67ocr
2Vrrj6zIWInwpfLimJ30mvijeLh2xL2+hk9I72bnJ3h31+9jpOE1j4ejIFbjrR9Q
ueIBGKHA/TG6qbQoCgLgr6k+FqoaLLwoAlAFaJ3czcMSMZNY8i4qA1vFcW5/h0j6
WEtKG8l9TG03GhZ8x+b2HPrvJm3BCnXudGPccyUKseKIpeUICh97rFFeQOGDqpr0
nS8Jemyj2+RKFp1WQvFZXBNg38uM5kbmOF+8E06GtWicZGU7MgBv0P+W+Libbeo1
tcsXQWY/mbsUu9lzfr9WovQNjDlIW31FvU+mBgJMYD/eAp1c7dl1dXRFaRxO3NVL
q+3G3Rhwa4hM/ZL6kpr+Ch3fnfUE0JhQF5InOuFGidKKoKPSp5KEXWBCaOxyLU/B
jJNjGk6a0jPCocrKpeBU2m4T3dhHyPk2nOmm9qULxyBUBd1NJ/Wzhrlk9cr7n4ib
wtFdPxi/PADDqtl6kQCht/MKa95YrO3sreg3qLZn4fMp8vSLO2Cd0wwe/DeO5PV3
rPqB8anDiJ7BSKGhPLhoyCxjjNhHMPbDyKqIwehoUT6jnQxKXqJZsCofqKoJOPk0
Q6Fz2wP221J050us1uRLALitavjTmpe1bY5h8SFz2sDl70MHKDzBvsfYsXIssQwl
MNI/2IR6ZrozOjB1gVUy+ehl4g2ihkD0Y4maiFfnR3gAACBq2FViuLD0j1WykrUg
ECVtXhGk9/84Zg3bnHtvJ2e45sBsgQM/bzHz+j+2iXPDbPCOb6Eh8oaLF/v+VYyK
XkPW/wywxK02dKyxOQWjTec4Z0/OrdkObp7r6tDotHT8+0kG9nFQ9PswyoHUvPmQ
KQqsZFpuo2akh349k0mCSKYDN/qOr5tVKdVd+X/AkaNt405sQSsR1Ew1DfJGhntO
41CWmniOL4XpvGzMQ7kwM+j8DMKp0Net5vdFfLn6lG4HfDRgC4tsEdforuILyQpQ
EIiCYlqLhT4aQpceumTcmviMnazaqxGTTThOwgZcn05ExZgV8Fw9SopSwsmJOere
wz0lyLfhRhGuO6cEPbqcYia2EmlitUts5Uzasob6Vae1XFgCy9GnaVDFY/blEgmf
p54snOqKQRAuPR/XYRJYGEfu/TKTLVcNVYqxu9c38Ey1bXUapljrjT01KTtBDqZe
MXDSxPk7EKvEXSPtiINKOaIMeWQGH5uH2WGzOCNeqDeA7jsytx/6TyxyjsAcYotE
cd9813pe+okcCvVTd6MutfWkPIySu2F+W9jCNoUiESnQCrd+YH+lUiaJY8rhU6vz
L79D6/OkMk6lv5Qy4xi2stJDtAdEN4HqOkYBEFPxYuGXsurrr7zHsF8bOniHXK6q
2x8ECmZYY8w+8qhVCIx7noNZzf90MJ7FOuyCZRFyaLBbVtU7s48ROUy9xABYoP2D
RyR+QQxX6bPgvBwUEwpgqGSDiebzE6xA0x3HTsn/9XnBs+fyq7fEbwR6+DzMcoPA
DXxHMubcVi0YRU06KbyxzQcZJGSZxQrk6f9PFsAUwcTODNKMoXCzk1CC+cVDpyK5
sE5qthLUXzF/N1CtVA+DP83Lp++nz479WFOcxN7O4+wQfUD6ytvqku8qPT5FH9GY
TSFomoa+SVZcYusZAuuBIn3XTg5hZERswY4pZZ720N9MEfSaex+vVvhCX73vwl8k
nEkwayqPgqqrOpSgek4sHKMe/wwREPEUW0cdi6P4jaixFaeMuUJqB1QZ8lPtZSFN
Gt/3Inrh+FgGpeN/W/bibcC4cyA1JmCGjWU/o6fAuLQMwfWpUFWS241IB5/2KXV7
LtdTQDFzHV/I6JkoVuAkqATTnR71rNJXxFOSnIiy3o2XECguFRsyrzfjxR6vzZ+A
MtfOD0sKGhO6A+md22cLrJcX5TuztZlxYl46LHW4DhBjyaSGdfVhczavYHojnYIN
xPubRKPnywBZujTb10oh73p37hNEHR0DUTMQGSJr/ejrAtRT8rFSVdB0xo5u/yVW
DpRX43Z1nTpWPsdSpVon1pJbdYH6d80zKSTWWOoveYUCYGRKWVTgamSo81+2WvIi
6Zpf0O7vL7YAGl91xeJfF1TcksTlWsdFLCScVdTKAqnle+saX6bI/dElnP+mEkfN
qmpeZU1IN5QVVQ+yoHp3eEeXPY4/yL14mQUiNPlJsejDECoDiqhuKrw8hXdcGoE4
Y4Y3ZEuiuVNp0F3wvh9XC9TUC4a8w/6FYWkzD/k+k/kUEDo+RQ+8tGsp2a7MbWjq
BqJaARjvfj2kg+A4ypfVPE+DMkGc14qqlRRJ+myaUgHhdj38E5bHP2juxpaNXGnu
Qojm6tPu0EsjH5RDz3c9Nrdp+fxJe2NHjM0k1x63cefcJ+M/hLr8gPXGJdvWGJmj
la86EeiJGmhz4Ivq6ZJOjB6LXoQ8b7gzI9wxfgmkR8MjAwo+DfP9UUJPanR3YjHZ
On57XLiJnAvzxCp9AbczkuwxBSUvH2q3pylrNmgnx0BSoR9RiWVLB0iH9f3b3l6I
UXqbeCz02vSRZsPU4VzCjuRMEPYYoZyC7msFajEK1fUH8QAD2SxDXXlkDIEfq3y5
T/ob7FoJNpHmBh4P2VH+g6YHzlnWp7c8qhwyhJX0RyNTw17ELdFjunrsh/tmkf+J
I3wmUxwEvLhHRGBgw1KonoNFOSBP/inoFFJYAh0uzgl5qtNL8CBGlkGFLSxwLS4/
i0LgxVGOZKPFuZPvPq4evKlH2bwl6WpshtCeps2HRueMUzJGIgV7mHEIQYstiRux
QdWjeGRpppReCnm3BWmSYhfCa4thxTLpv7ro7RJZuxy3IAz7vDl5oQDkKpf9fgKQ
Rm0OqfMbX40+JgJmnkY10750TwskVi1tXGP+7VUhQGyBTGIYbujfbZ5+zlnpuzPw
IWrYKsztP31pW9ExhaPvUj9F1A36UWCa3gLHOl2kfZncNJgQ8VbHZOHSMkdKh6k+
1aF3e0X66118gOJdkpVXbx37hLn0+zewNi2LSDmmI+xcvOWMMhJSAIVCFdRudXNq
mpUxTuSUgs5s+9lwQl2ohZyTLUkmDlLM9q5TPnUgAVKT1n+KjNTc0ETqQOxGsBUy
ql4WYjXgBr39EZ5+ZDwayjEHIV8SH3OsDXCdNf4T3GfDEtS0rGi6Ytg5V3rJLfgz
jlG/ukw/marciUIzNvjtKJS3oHuO0g8Ld9L1DaNBA3NrXTrPM68SzSXmHxb04XuR
uFxjcYFR7y2DHS0m+b8BvvcqnoG5BDvJn39KLz50iNzhmuM0VxNLLUmwtEq4MZDr
vJ85V2bOUbbfZp9OWg+HAP8qTzhgajPqwYPnUmKQT77BvfEwdoSraDHzwonZC8VG
B9DKkazRrzjxM3bYvde+IfPuI6b+967WLPmGd9JxBnh+sdRiDiDbh4tTtsuuUf4K
Ju+7ynu3Jq9R3c+6WBXl/DP6vAfC+U/rJrnfDUcSLsSS4apip2dbWCu+MmkBs+qG
0hSEq1GIaOokCrXyIoXdlV+7aq9x4OtrrM2zN0l5R3jUusxsMBeGFYm0dSLF+dfJ
1jn1B9ANvJwAwyHa0pDsPbPU0KcW9PfPtticqlyei5TN/lZRPtcdJZ1SgwDu4X1z
Hqm3isN6qM9JKGVxfQEUitvUfyO/Ht3SlqHvVN6QrGAg5uYjbo0pkijZFOH2zl0s
m1PohZImEPsoJ5n4+GXwlKlj35xJheujqbrK1YIqhoxm+SQNd/vSIrmeY1C6apJI
uthA7JlAfmMcGB530XwFKoVopNCQU9WtWhEbPQ54khurcE/oUAMUD/DOC1X+Dn9U
eU90/YNBeoJuoUf2CKQ8lBaz6i09VG2Pjj+2Z3BF7qiawxXELXoW12oLCAGg700O
7HzcYyqr1wJYqNRaeuGFYQ5bZnIS+cybys/Y9IuCMleqPNoSwyZfEYuZ/QPZl/MY
LmcZSLLh4kax0W65CX1T6J/1e2ELtdRmN/4GKOnzlhc7EZPU3oadJJmbi7zU0nP8
kQ3oaLzaw5vePgn+/bOJToj4hrH56micgzxnHYq+4Yyd3xqxn6KHk9ivBP9DGCGN
LWQuKf//gOlseOq78O2ojWspzUWFK6Vjuvs2q2ZR3YXrW//0OAp3+It/lxpoSwLd
2GKj6l4dG+RFfgHYPCDmS3E33KztHlQ7fjbgwBPR44EQjT7xEFH9YUkR9W480WgL
rFnzx8Nzy7fogEAQN++WhsLh62/vGshr8dqrMCo1IwidMVhZaHnyVtjDO3N1fpJQ
Y0aiLUZwrsQ379W6ZpRq5ZuIe0OEniflnIumO8B9mKlFRQ7Umx38xn7DdJqPD3Jc
1jeQ283rvdGtZiJOrTL8yocG19TCNYl9AO7nkmOQ8Nsi+mq5n+8Iom+7vhjOx5Lk
qFx4tsEDDxV6Y0tXKYcUmON2H84X7/lIq0QyCPawGzyXLhS+fv1kaLrShZCItbzu
97UW06SL18pqzHEIPsJJyiK02xi4auxtrW4RHY7auoM673apEyAoC++P9OOziYvl
BBFHiexbcCIYgXTz6Ce6G7+a1pPXmTaReGCi8enC1F9GgnvDtLHAAhEuY4YqwzdI
e3AlBVsR//ms/Q9+JGMxmF4wOXbtTrEvcgk17DuxbHfL98jrykBdSpxp8gcjQTam
Xmxr6nMey4IoZUFedfdh6cRUwtBmqzUn4OC5YhA3H3U475Hn84iePbKrMDz+6oAx
uLPzVO5a4qcbZToQE2f06M/28fmaTwS49UUubvB2Ru3m58Fu9motVDk/nulr0dm3
aA3it2P/HLW6MOcmYMG6HkviY2KY0DONoBl7UsEVG4Efvtx3xFeQ5UZaH7UgHbka
GIrohMHVvS3RrRjuE0LV6xoGi9L9hO6/9X28lxolKiVSLLGyc9irUZmzE1awFIHW
zGyd4gsxO6GYc+Uq85tNI5Kmw8o/7Amhynwk/Z+yA62tZbIDYWC4tnag2nolnvtS
+pHMvQ+sAEiHgLO0KwHWCTM9/9nMdVxj1QipWrGNeg4vq12xV/bwguB84r3kgcmK
5ThKcE9NlBAgclovODWJ2+Ibs8Rj+tvD6edC9sOHReOGyL+JqIVKB5KPfcvYBFQQ
lCHuOOBVF9OoIt1Bv4SYw9cj+Boepo3H6313LK4Qd/C0eQ5uXnQMSrC7Vm8fnb3j
+GurPhvwOkW90f+cRz4R5lOFkoCJui92XAqSLtIhZKLD3vmTP/QoS0ZMxncPOrfU
VaI+gMDUdweqFKO6a0zenJiaGikyC2pTFRjKLEsmluV1OqYKthErgTu+Uo+IKoKj
Q92zc5XhZUev6h82hF3Wgp871dzjQ3P/dveAyKFDzlCUj/inyiNGiWKLZtgT/r4b
hIJFhBxlJ8yDv7Wlsh9oHPk7wwXtxZoO0NpO5+93gt/tD+xzYs40QTHbdNTnBgGI
qdCutZZhDbu8vh9413rRTIs7mEjo0TfJn2yioLpLmtYT7zY+9LFQRpu+O882cJj7
rC6IIdWMLc4NTXHB3cPCZ9Q/qSIC2sq0zUgqnw6fhqGvAA4VCb/LgowvsU8+sPMW
2rkVEmBE0xlRvAsaO3iq5mc2UxK93t6/d6gKW4uUaH41ciY5EBa7KndmNpKmOhx/
riiF5UvfZlywIMnnUw5eKWRJU1eKJBm/WlDa7NkTSRKIaiT7vUJ3LqcNKnM9+JJU
KBe0oBISB33jqFvb0/dNtRvQKpEA+joXIprUp4Rbub4MH+9TeuqvRMxoeafkJbQl
FmQQtvOBZEkxcHy0FjGNINyrvaMvhQbVT+HtBbNke3K9nUoVbBOx2Mxpkg68j8Xl
in0CdE9I+dQKbCZqLsaMPAJ3WrK9TrzmOuFH4RlBvNlQfEa7EGFVWE9xhJeRuWi3
YJtHIxj3X03MV6czQEHMfN0M8sxo9GvsqxeFe5BkPgrX2zjgcZwISALkWjpunuVE
dgzcsKOIKnaVUPCXeOftTcJ0NV1unOTFCslvd34fHw68BFhAXllrfTeyAaEI87NF
dEt70Leedk6y71fVb84QpDwBXEPKqwfNAjaX/Be14U5XRo2MDZzk+Nvb1ikI4O0O
uGILE4Icy3/YYQxBsal0Ee5gUOCLnTMSe/UPEIDEl0qEXSqHZNbDPkFZ3oC1Ec/3
uCprPOF4zHQTpX6Zgn/zZDQ2tnUsf+FuBfBU/PZRv+LEV4QPsBH1V48WMQVF5DZp
aRGkDRUY2pT52mFZ0MAaQn27fYDSU6XS/1WlkK2KOqX3wcjAd8f/HvWf/3UhxslS
A1fzQRDZSFXCRN4I0cC4tpfKCDLY6j5DgGnvQcuewvayh7qmm/Ds+5MU6L6FGL+w
oR47fYw8mtaNphU3Www+oIh9GuEiJZBR7n0VJRXnD0eMXVbhCETtj1od93s0YluP
8YWpEDOLsjVEuGqZPINaQy443SDtcVJYaK5I3ufY3t7pgSVsn8TGBxd6B5Rg2Hvt
SgF8yosngdyBlBYY9bIuSpuEvzuwTGM4Jy7uwgV4k+iCwPSvsYvXhBWIX2+d2Dzq
p2jNwEas8EEOhsehFpWNFbiT+7w3irDVl7LxAmxHR93DH9SU7LGye6Ru7aZeEMtq
kBs1b70gx4fwPZHJxAdqA8PcV5wAAf85VyHk7A3UIXrAreK57nmeyVfg4tie25il
nPgjAhjvvr0pKHGFYddKoZuBq9ziGjWIs7dY+FcNpIwsVeIevHhgnmuInwJLBXD7
K86F7xR/ct7jfzgjElTHP4cgKSDtTSzAMVWj9JrG3g551wdmmNuPTIehcHBAU/Qr
llYzlj0iXx0zMDtAAeK8C2GdPN5Osq1dEMLS0uK72JN+OUirchDrJ41HXxRRfXcx
KIonr0LHLI/l41aClaDwW4AcCBvTr2ajgOtJOf750k36ndO8xJPHrE3wz/rdOFWa
S+BVO1cIOzu5rr4pecLhCrXbHQf5/c0kTDPikIn7RHJa9qz+Iei0jfGdNxLUyYjr
xwy8ZfAhgck4Ta0G8c0qIocPKrLVNZXV8tHoCYd9zPYLv//1XUiJiM6dcFVrKola
wQjfoPtIP8XWQBtZE2M6s60+ztF2gFxWh2rcpJvMOp2nKx3smI18XNrwS5gF0W6t
CWN9OdzBWENFjVrsfGreUjdSrOBkjHbYrHfa2dqdp030vNsYu02J2uK37+oybViK
B7VCcSTdS2PQKVQ+m2WYchRZRw5XyfHboi23zdcW19hr2/I9vb26NE9xPtTStAG+
HCcHgipwZleJAIlGt4F4vVbCjb1WCfMQB8zpqzQPJ1VUtC0aoQAdDmXz8tirQp2d
gKZfiFu2cvd5vZJi23EPPsA7A7b+AdjWeoHcGXFzLEVTxotgkB3sqbbWhTbYiA9I
bvmJorFRJLkpjs11itHPnpAF5nVHQcK8CivP3lWq9RxgnnArJA+520CcpGgUn4nU
HKsOCc/rtw+sivYwNU5tgOFeXr/i6aSkzH35afKC+XhoG/YGAJw8BUdXFflaalJ2
QOfsMc2bF/FdTL3GiGAh5zqNu//j+B96szBbg8t+tAgyKM47IFYX2fL6yiFBve2M
83hDaCtyaNuWmHr/GutQo5iAwKUzprbwFYDfEa8cOIJ3rLoNgElWBQM0InFH0+Bd
qIsEL5/AwPSF2v15Kg9HlcjtOXXZwFZ/IzP5qux+zZOg1NnrxnBDvjmVoHm8efrW
eyMdQcmvG8DUrUfw1WqmhejDQ8M1J2r6IL23ypz42OETOFlU0oTvvg8E+E2vBXoN
5C4PD0OI9S7T6SRZIL6y7y98C44O1VZdcwaNAChjRYE70nTuH3mNokYOBYnTInb6
xaWX5sdYumlXOsssoPLJpv4YuNqtIPhH3wtDTKepm3qlB2oWzMv1fG5/WUkbQqkv
pP6JeVWQ2Cl448vbg3a/jSN4DRrF9+VjbLYl9eWaeJQEK70OVI32tvQRvqJOuDjG
7r5EhlS6o+C5WOtBh8pHRSnryzPvTIW2IFszCDl3AQNe2puwMPvk2wmpJYTo0G6s
xNrlDTY286CvS+yWQFMHVaiYMO8Vdbo7UnPjJHlFiFGm4PzAv58IZG8YN+iO1Y1y
weRUieqchreKVDdY5RV2vAQpdoygjrIDXmeabBF8cxJwL17ZyUivETt4DTfbcu7/
jMOztBbfAwCBUeFJVwPxZaEIeo/yu09roqRMX+5vw+PmoU0/D8O2VkP0Xtxmfqom
i0AfMilPu+sRrYJnXm0XPKF9g0wgisnFddMI/vc5fLH2WM0STtq7JCaQSFKGt+gz
wIIhbl24zcQR0u6s98hwVK+eyD2oag3xvdfgURTtC5Z6xGl/nRs00+KIUQZT/aoX
s4qSwY+Ibh70DKXxGA5zV7lY0gIApCO8ej24b8RmlfjcxKbohU+0IC91460Zc2Gx
NfXSBXXcSH5Liw+zLaDM8wccBsUf9bPYEB1/oTmZo/k6zBhqrYKib2L99pCLZYmb
W7s2zRBjsk0NeL397NKJPHcpcXrOPOR9DnQYfIwuJAEudoUZqkuODhz298GS11Vw
7DM5q/vskHIbeWz8L1oUe1OJiOJkiwqS83PfjHkVT4o1CgtDLOuQMlpxoVMuuUlG
R7Cp2jli+XuJMN19her+6DkVz972mLd6oKFBVg2kIs6udbjixOivtiWRcK//pI6k
S9PDhBr1M88GD4M+9wDr6J8bIYYTUdEQEPTkELI84RLGY1/ljm1Ch5y8J6r+IorB
Q1+8iILmjX5e+ZVMKyY6YLVM91HL9/xJ+/Foa/St9kcL9JPJkE6c03L9AegZ5amI
28mvLIdVqdL9Lae9D7SjdcJJztCTOYmjYnT6dpF+tw+1zwte4peNh+ALYGDyxnmO
48i8eAmprp2BKm5GW7IFgPZSJVui4QmEqx2UkPdu/rPdcMJ48IlnqGgR8M1f6un2
7HqbF3cOJOiVyA28U1gwSwbantu5J0TNcTTneqxsxjBdKqkQBDDfJ2OGVMgHltHR
P5JMBov/t15eIJjtP5Vvq6jVqiWEiMs1RMIsJ7df4Qd1DrWLVAOB44x7vv33cuPY
wjLfjjDwYjl/EAPKQ8irtuc1xRNCt4p7+0TCBNdZOB+cWs3hJgu1ChetKD4bBt35
f0sZriZ957whk4SSZmIXnjpXTdQMf8vadljIhF5K3kPh2TC4ttNJjYm3DHqSHvMA
Ah9I6eifKzmr0K45GdioQtCLyFd8FcOi4D3h3/p/KGFQkiHJcsz7gw0Px4uHHiDM
ssAreT9dxPGYc41IqqnvlpRONlHcgr/zmKfzUQWzX+RteDJBCY3IhXZtPIZDWXGd
CK67zG5u2nHpOMu0WkhVnZ9YcKoIQzpS9dQurfwN8PXh3j8ClbMhfctqL6shxLSc
PvUMk4quqcNrWWII3ETwGfODWqI49ehvuyAwAMSCKbOT/Xzcl+ssBu1rq1/Qd2HR
/vs9h/6GaWSTh+KlHePihAzVziq+IhWXILnmMsUVbkNKOG+JhtUW34RCEPlQHloZ
K0LR3tmKLNDDedf82sEz3+/FZE1QYZ+CAqfSJQ5+9O4bZMwB/OJsO3ou5tbc2p8T
qEyGjjUm29WJpr/cgsMF3kl6z/gDVABPMTLKfC11aiEdp1UGmB0BJ1ZZIqtNS1we
xNhsicLn4Hjvud9P5boM2vbIsE5qbftJwQ/SYKf1Eph+XEu2UIir3v7QwLhvSFzc
rlvENbmRtYlmNsTg8W8oNPmLZxwqoThYMHjdDroqk3nZ3ov+8oW3mxyympo9E00N
U09MG029LTTpjL6lkZRRgiClCoCgXMlS/OaATYt6n2rRImmCUBzl0mPqsj1jkqyH
XU9l8v9+m/EkHlu6hxgZ9zhZieqnt+tsbjXQH/kOS1tYORizriNBiP/Dq7hn+vrT
9/jFCyeLk/TAnZiJLqM6fDqqFTx0E7I8M3dQvDv5UnDnohBnVj33KCTOJrEgzGu8
CzNF3vupOYAGw5xiOKVEuO04pwICkCh8JQ82CjyVOwYRY48Me9QDItGo02dgBYtd
LZVOZFQgU94KuSFHeMINZe3zw3dKmsPUQarM72ehATLvhK9aAx6ueKxroLddaXu9
FJ52oak3clmSm7BO0j9R9MBcOHWGpez2khM50MUpyJbccMQW2jeyqZpDAyclgUhX
9/1SnX3cgsCOIYm4Y+DplQ6Dk8oaAlDXrcsip4AZ1z/B1VZ8Jpw3ZaDb4pLhA/V2
nDBxj6GAm/ObDVw0qCbStu0vxQprcWinoX8jlyxEaDDq9EgInQcVBhHUWvrph+Rw
T34rG95SyK+XI11pzrWuxTXPploRiDqCoAgDO9sihLQdcGW8d+FRUAQnapOXl+4i
RsdXBLNpz/yhqAdOO8AWPH1ML27NKFsWsMcc55Iqxbr2gSFIgMZ6ijeCOkSdLIKs
3hKVAsLm3twn9CsQTaRrQBN4P9fwCsUa7mfqoWrezUXm3quajy9ktXeGLQquKU30
B6QountCAQOZq+VsE46kXxXmSjBtm61317GxIazuxO6U7SgFM9x1Z/sH6oKusG+w
Ns77yIFUY14NwHwOcfCQXJF2K6kmTUJDsLZoYYi1hJbbaL4z4h/naMT4dCqntCS8
DYGFp+NoN5CG/ed4Q+T/nUKYMVN7wQZ8yDugYP+1Yn3gTdX/9F7XsDpTqWWsXZIk
y9o8nuRO6Nt73AEOZWF00ZaPs5KJIyFBah4tqvhr1hYNbh3kTr0rLBXkWdARevkY
Sq9y9LjnB3xd2T5uk24P+qwBimaUBUlSrx4IwhNCshbGOgvhIvFu3ty5VwbN44ve
D7YMEkvDLBmDgrrpEXnMsDDyOi6wmkUTQ58iCLr5P1eo43SBAx/JVoSuF367kyjo
Y0YKzG+js5T4sbSQjolhjs1uFchVBw/6LmNa0XCYaY+wCOP0/0MFD/cG+7oTB3rc
8vevK5RCzAkrwS9ZgQj6ZiVLxpWDhrArVEYjMe07ttvHOvFUsrhwbJaf/Jf1p9T0
2h0ul3yAER98dpweW2Z2I9Oi1cQBuSjV7ZfoiDfT05QzIr9QuWU7uxX/8qXfJrbN
vvEsm2nU0foHB/WNMR+Ke1PpwUqZvKXkMnDyF7eAiZ7Taao7D9WrK8JefZu61ZgQ
iv7VsVMShD8kRHlq5ekjjh2w56NsgCyzwfcSO9YXkWJpjsAhZ3WoQ88ViXinNfAD
P5zLqOmcEezvk0D2HM84OZTlLP0+fWFVx8HYnSjrrw78+EuYqDTkuEB6SvfpWlhY
Hst1p+/O1hCg+WPE6TDUSpzpJHVXt3WOk5V0rSI1z8SyAxijLqGusVCEDxq9/phz
EgPcxJLZh/FLK+yKlnX7dKdlIMu0NbyfsY79ynWzgje0PUB74iaXCofAB3yMll6n
Fv6v13LM9SLfSr8+qPX+i5Q/GL2i/6y7iUZ3ooGwxRBdSd4rok0Kfn7ZpcBJ+caI
Ux1SpEr/PkvxLNYo9uE3FWjOyhE3XuyeT+UO4/DvCwmzhYY+hy+BEi8UfYpAhgDJ
4xsPyim/OCRFU/C4nr+HvXOEqIB+bjQjfqyx6m1AbBRc28qg1E/L26vGtKawGbOU
p53zT7KL11iR09mNtIa/7TFR4heXQZpkBDeXLLCwD1Z8wkyetyhdYbw5W4pJpYLF
mD4/5mkuUq5EqRzsmWvp+9O5Zv06g9KdeSE830sCwLCDT54ZrEsEqSAi4Xu7UgU5
vpyWIZb1NciXiTiqGmlArARdgKhHymb9Z/Vz0rVJvBX0PV4c+VLrOSuNq+Om+fJk
rOhE1kDdMk+BjDOT+Ei9WNw2wV6t/1D12xkgEbO76u70oQPW8Nl6W1P3upjwbxL0
qTtAL95Mv1rfPXjFV0g731jvOrKG9hAi1GG4jQyZJ9W9d3tKV3CSzGkw45tyWhmK
HbXUBf+Mh83kbzqi12HCKxOKB88ZDMNg9j8efylOLLLqbet0kl/XlTP6/G+2IEco
9wSNlwn0+a1hqUszccJqrZqmx2OT/fqhL2zdQdCFngKxEcQ9zN7EdwLl4Ig9FLV5
lTv2/oVT+5evZwvKeAfxUUcOHfAd0vQavH6pn1WnkrXAHhtxUpqwzE67DVBSaxiw
Z+6YOLexkiFTM13IIk4k52NlGCFpYHqnCsDssF5QU+Tdgp/Zj75IrhxLXvaTO6D4
seFLXAiqq3QbyjPCRpqEZQxLTik+75IYrm2xOgZFhnFuLu87wI6zmTjcveRroIV1
f059fN+V4O/Svt8C/t6wH13t3qckk69QBd/Uq7IVCSKbY2dFZ9wCVihb/mspbWKg
pDCkWZbVA4qEqfrOQdKKggokChRa4Q1ZIoX/abjhrIOs3SHiuTAG3uEODmu9J4HG
JKeKBJaGRZQAV3uRWW94gAt0p0NN+13P6r6Sjv3y5KojVrUYMRmBbysO32YQ0wPq
P5CLYIZJEC55gm10/SfkuTBUAndQG+vvfqaekVptvx9eaTCClJm8eXs8xRUXuWvM
Ulx7kAus14z/am6dFyDcKiZDljIbut8BTEHZFz5QkO1MhXVz6SGxOJB+Ou5fHR1f
k0lk9L3zEV3Tvc/uAcGnnPTyK4JQqmVW47KsMt50xFD/V/dnqqD4gU0xNxUzQgw4
hYHSeFlOECqCGITS0vAlt7xEOiaVQwnhPiv10IYrO92E2syFQSWNDAGkmO31yvef
lmDa/XUa3wpuHbeTupojaEfDInEUudyYWcMxHAb/LCoxqgfMUapG71qcjFNyjHOt
B4eG9iyYt3lnADRC3w/0GtwBVE5ifonzlyFhIvnUmYF8IOn+RqB0I7ekholRIZr7
kh+faF0vlzXEuinulwKqp8Hs+0Psj89xh3bmg1nLb/uLEAzydWxMuw+1kVeReEgU
8Lapfq5ugzBoVHeomRmCuabG4wFR3QHwuXFm6fubeXRQNqCW1iVKcX4wb6S7LyJk
vOny0+C2xqZUfxxZUxVusBovKWSoGqHedh7hNsMqLJRuNa+ab9OaMix65+V1ijU7
6AvzisyeS4jg7S/vvt8bkIME4kGV528OuoKQvM+D1FGL0hznzs5cwhfyD28QSmqQ
RGdF4y/Sa89Xr+Not6nMrBV4nf4t7nNtuneSc9tSvtHVvZrEzILSy1AD1b+N/1IY
AleFwr1wTYNRRJyoOyL+QnxsJsEwQBHegUV35URzNq4jAQDeYCn32817MyV7gRoF
ejg783Z5uwAx01ZM5jVxwDogSZgAu2XyKgC+Lyv4NIU+6Bq9qpZAz60hLbY9ODIE
8BVzKu8yEta5klhfT8w2v98EjlfVBn108Uzvv3+vnxywOczFvY7mqMnssvqZjMqe
ABgLrsdTQMtpnqusPlursIv00fkfspFftBTIDyDuOJ72zRTQIF1h/EX44/cUjTBo
8I8k2Gy869FAYbZ3+ijJLsF4rIyc667cXP4CNeC99Tx1UxyGxEbdiA5m+bqnwkHI
LhoRNVqiN0SG5PnCopynvR65j700ySMSyuPsPWViRA0XBoM+RnXV2tBRsrUClRyA
LMlHYYovDgrpwR+To25YGt5ZNRUzu3qzJspAt0rKShdZfeZM2x4xqIxq1aVUB9MK
ysCfWQO/BqjdSZeDKVn5GG8tC3MspdDqNUhbMNT54AWLXyNgnVEWOxTpuMXuHJbr
CKq8m1FQsKUTCjahjYsdKPQQXn3Rsg5Y1XUIsM33ep19XIw9VpyZlrohdfM9kaAG
+tgTDzOJ2geAo7O9b9VLcrSOwmpZledODBn9U4zJ5e3YQv0Sv+v0S7x7Lgf3ynRm
fJtwZgDsleYDCfGxox2f9/8URRiCBIW1UI8IHM+FgZffVjlq1a2CE70hxiUKfHvd
MgJkzMrhaBtcJjBwyUTJgNjGdTGsgP/wPCTD3XG4Gu+Y7VIzhe12JTHofRryewZL
LTJ6BYE6rjTOxiewtDd9NtGUNZ4kqL4xxlHDToh+P7LoaxMSJ9dNhgducP9a69MM
UZsO7vz+MpPcATclJNQy/xQWCS9u7lMgaqcT9F7/JjQPD8Kq8HL0iB3caQqVnYwH
lJBLHMX6Jiqs5d9AoFDvdwDB0PpeDDDk+R55P6FqtMgsH134Z7+wfCdN8jSSp+YQ
7gvdggFqLjZ1BVN9tiVsRmtodVf0dB8uRhTcu3VOFnGA72KhrB7g4HcHUge1ly75
wKqc66QuxdlKVXyIm3OQvaskr414XfwSlKJ2fOBksPAAJ3KcNr7WCqBEyPkoE94P
ZQiRAGzzmSrmiOrb3GmlXJANNXBVi/ZUMtBMroHhj41zOU2UUam4JpLhoKRcUt4y
IHIewQof23LNnsRruJefTmsh2xZIlUHySJKkyz70iNM/QZfyzn7EyfVYWUDUNK6I
B38hvylZvsbro7o987WnBiMDGx3CT5yGBPi+jQyb88HYHbGRVqzE3f1dvTH2HQO3
O1ctJRYc0F/XlLdcsGmttXEB5/p3WBBK7pT5ZzcjNwO7so86OaOsy6ABK1QgZHti
Tfst/wQeoqP7SdF6UX0ar9zjJU46ltSQ7B3+RzFO79STlulOiqT3CMT2RpFX5ZiB
MhqXGpZcBM7Uzed5XRGK+ln9Is7MTB5I2RG/CgwczUpip79SsxFo7Au2i3H33Kxk
y2myZNSVadDTzwLJizyMxk3SU4uTa+UUg9yCJo6/x750iBu/3oeiWwJwzNTRG234
xul3KR17pYIO9btCSxEL89QQ1Bpoqlqo36nAzjiXVGlQjAv8q3ayImmkmrJffx/B
VyL8if2ROcPtke5OuDykPfOErXADVLRPj+vIGjOuAoAW+qXhh0arT5gGSxsT/2DW
Ixq5JKnaGh0ovd1QdmdOyE0W4XPDwqOnSclLm6ACIvu2jbQJkmzLdLcUKEzlqgRJ
O2l0/6lds8O1biNOKwKNaeu6WzRmW0USQ7uQh4IeW1ndwCpP6Nm1vEYEn9F+gU3e
gA1CyifVxkimKk5Cl7UcDMNP4wle60i88n3FyIaSf3tMHAo2erZs73YlKFeCRjxg
4x6tcbUIMvjmaHTu/1YuWq57m1ODiZrUP5iecG2Qn0gLff491jPCsEcfAGi3Ty0e
O0qi1Wd2O588B3jjN+Rz6f0YjnduyadxaEuqyPVpidULQT7GWy1TkKlpBDhvWwmj
OvQy7AgpB3Qq6s/Yga0iXUohIiHPE6svjc5vCoH1ICmj6y9pjjoDQR/n8lE+GsKe
0YJ5YGwjtDhX6NJ1HkzjtD3KWJi2WZldP/RnS9S4tDwpoJS/qpDT3CjZL808OVV+
6j8KkDkx1C12ZFF+SZgTRWhd8x2ORtFiIb0ngfn2RFLOxFI7FRjPLmTReWoSsUIW
SUbn+rHxwqM+CeDK9OTmYh4MGFcT9Pkwlh+ThqLjDot5pIWz/uJEANftOPyFkuBM
bdF/FFyxSTUgKQ1Qx52jbtrJUi5j+sQ4n1oXEMTKJrjhmHt9cu0cT1x/FquJ11dS
3QhgcRS9UdUS0cnCu+q4+3vM0RCKMZoHHbrDOxBntdELg+mnLKkBtTAKOJUgHMp8
SiOKHydSDUkYZBBj+Len39ZBHBYWasonnm/UgPJBHdyPEECLNEz71NCh4T9NT3lx
NM9ib9mi/yHzSyoOkvh5hcgPU7W68Dqizb9/uC3il+Eh9XpiJSAsKNPnzHa67csY
/rTFUOXJcl8PQgf32yWJgZFb0IK3Qchc8yFOeAl8fn71jYOZmQf/oXy9Jj/cuQ2v
GJDkjokZTXTYgM/x+jxp+oGoQxlWn4FlK/PesVXDKHlv/BxcgeJU4noKcwU6BBee
EefYfZ2JT+m2d3FgMCIFkOkL6AL5xdQFiQPgv8/gVlbWGM3rSjj04QFlbqCEUlXb
J5x0xCAg3XlOKBw3n7xiqg53AR9ZeuL1lONAVmYDh/KJusXKdsC8REey95o2emWm
moPscxXUeQOwlmoeFyOdhb9/RKiesbT3aw2S2pC2wdRbvOBmnFj8zbg6nSejdI+B
QUTX0l40aaQLa5n6F8az9CvQsQkENCXD8zJz5uIEuKZF/rCqP9G3HBW3isQWe2sS
luDbsCRcz+PPdDI6HXzurksT60U4DVO00d+w+teU4dOzo9gSAsSh27blcAsSKfdQ
n8nZ1pQIcrG1tX4qQlG0ieI6edXAAltcL+28nMRsOUAmw6vz7xmAfjT0/LwqRTkn
FkHf6Xb6+XcgRf4ouHGL8TwA1ZZInSwjRQcNtRvPLHSJQfbqvcKtVqK2MaP+I4ef
eS3E0Ujs/Sp941aSWx2BglM4cxGQp8/Y2cGD3QvvGexlgdL7pVJaURpz2yXa2PdS
rd/5w0ST5VFYL6hrd1GpWpJ3YrtOLiCwCfhmVWW4G60MFuNgjQbBoKaOvZ4/rgPL
02iHwIgJqHc3idfBOs6wQJ1LzcKu48fhX6XhDtpmbWNYX+n71/1ovI4w0rCAc0Pr
8PzkRKxsCO8jHqBqrfrj2DAm5jjrnpCu4ki1rL/D+O1t4FRQdM+UAfn0g2Wx743O
oKELX7CLeie9VKfvNIh/teia0d91M4DqTH4BMfscVyOrDlBNn8BmG8crDMWg3VYK
Bwg0ycsFzLoauZN//AuWpQSCkN5FNB2RnXQdrEgNRJQDd5Npmp+dkXUyhSVQ97Zr
goprm1Bjc9kzgljnXOMhqtDrJVoPRYfoOB7gB+MyRt+JN6J0ynfiB1S8dnJ238S8
x9vFOhHfnTN8/rvoTZQFcB7IL+Smh1Rt24GWUYJCcAsa5byh6glTThHYDruZT0Am
vG5a21IJhZPi8aqm+ID6Tp4F8g64f3nOBY2jz/lUsmtwkmSCnyOBTU6IOfODVO4I
2nkWtrvUDcynpGpHmVncPMQfLu6dI8diFulEAImUbOShFtNeBuuLeEBiWAMX08R/
i40szHFJ/KQFDzgJkjL554Ys4jtcQJR4m96Jsjy/CxlcQln2ycM6kFB+ticWuaOh
vlgsHxK5Jm+LU5RkFF4Gd4xkgdtZM0VoK94x8ok+Ooh0OvFZ9eLlUD8pSit3VYa/
mv1XDlWuztCknA380w4Vmu17rwaT6z+kYB0fhm4nqivRgAl58lKsd8CtgU19HQrx
ijbbXLYBCkfg5nlu/L2yuXWb5Qj9cqvwo83vdol01qwz13EdJ9clUYH4napfJaVm
8+lyFD2tvF+Az0zDa5e0pG8hc0x6nqlmwaf5VFuRrWqXXyaO0akFWtoxUouzo0au
jT+IzCDnonZK4uNu8e1DI9mg9uYOz/GT9g+Wfky2cgVJdaWnVOm/W7ZFAW84ekND
a7DIqg6kjjeBRb0jJF8XJhcQJLmXoGCutGThjg0uVF+Xq7GyWw9lpFqrGK7y9fcb
5MgvXYwt3875UAlpjWRgCW2DC5douo8HYimb7IysW/tGJ0jLCmWzv3mN7Fd3KiKL
8rqFB/g75JH736nt2edGVgc+ZibsvUdmOTNOZFeqoEaycc25PcEYOC1ynBPUuQSt
Wc0JId5hS06DgxVpVeNuJ4q/FOe5NZ2Pik/0U8GP5iyIwYI4cAAsXffp8dV06t5v
/M+Iy8i6AeaiTlH2HE7ksASntje4XbFznt450jBK8av1z3NKJM4A2XkEdaKUYJoZ
3UDl30yRvj+Q+Bjww71VBhY11rEf/l35mGyuVpCFBzvSU/gLUk2Z4FQcpGwEbOyb
xkBazwqYGdCJK3e2UTl773jm300x9i2UhKQf5UAlofQq7kGno1n5QiO/ScUPnLea
BaZAXoFEopfzr2lszN3L81J0owBpMPpr8dRrIngTOr0d+itCAh4dboSq7ux9TXOX
3+JlaMQzDKtXM9UG138ED9q/shS3zQjv6kvLw/kpTUyfMXrhbWA2RR1w+TSV/Inq
KAqbvyhtqZWPYZfb1qw2vkDo8lP5WUU1DZFLEs29VTdX5UEqlCcrzLx8eNCLVn2z
7B7R8lq2sgpK4XTgOSF4JLUP2g1/cVsogwO7v5alPMeOcf2hg8jKe/k/UAoI3LN9
LqVlJcMY654BrmyncQu8u8+RINeT1iO06Rxx176pXEhcINYZZJ+4fpa659XQosw3
4/uORq1nTlvw5ScjQLKIIIyL9pMuFlEGFzNCtTRJX2K+Xhf6Yzj9J04uxpCWJFkm
HoAkjy16hR7POhv+UI+8delv6sBca+MAp4M9TQS2zGhKosa32JVonbLv8gSMv8Ev
bRdac7FO5Vz4MRbr5hVx9E9gjmZLk/+GZl9c4ZlgOGvt96s0kMvm86Cn8LeHz6QG
vyLB3YWqKnfdyj2g6F11IMDvgrXjpcsn1sVHSdf7YMZW+AJJgdDobB2d357SY9x7
iU73E1T9eGEf0AcYV0WMZCrIm8VFU2eMeXWunyld3a5B9auyROehxkOkjGDL74/S
mNgRU/8Gagme3Bgn13Mq6XBVwUCH1TsjWiZIzouFGG3HYrT98bSnbx/UXaBiQgHC
x6P0EgFtB0DWNinNFUkdLrraB/fi3oW2uMhjBIY6K7oB3k4fToLS/HYsfUqDZNIa
LjsbykKqQe4AZDXy+bwrHIdSKiCwQ6Rt4r/wMoOtEVBnKByDKI+1Ay0ooD5KhtUu
oV2vAhHJOIEboRvYThlFlHVOfsK1qZ5PcQ7+VH6K3F4CGGuCUe0IpCSYgs51WzIa
b/WFIoySLZ0a/zZQ2CfFiEKtsn83+kLuqjFWaUasGz0b+KRa5BnAavScyxXrq68L
qDl+KnfBG4ZunOrsUISCV1T/otk7x2NF1WkwqxYhFft0v47PWdPf8GgHGxkwwIYD
6IlT3Fmp71VgTJ3pRNoihmbK1kbD8ETzNA2c88Vmac9P3LGrkR9Kd9fvSRA46poy
Dd8YNHMrMyqNoESVSUrD918udJIYC3nHXP/l+BZY9PesxCmEMcDD37XEHYCc2rmd
ZVu0czAkqiXokULmr1Km0kxuxvW00jglALI5fjxBJPJfzS5J1bkh3vKZtlBcf6aU
8qJMTEsENb66vwkIDKCRW4O0AxEYgobK9TnMpZxMHVVHxG7Vc0A+37Cd0SQw1VV7
y2i+rFuuE3QPIaVRUW4O78oqZk+O1Ohwv2QSUl+7pIibldzzsim1y5QsRBA5u5Gn
nqwr8hCBclD86+LDQIMY4JiEDX9QBulPlpwqLZhWBjVuZ+ki/fNVvvSxF77AoVIA
rPUb5GoPWPw7a6JcTASS9zyk0+tAH0U2vSiIMkfa5koI9OImhSLzGxx4sh36fv0K
OdO3yqBTikUQO+QmqkM6ihvYlw+GsEJUHzy0B8HVPPuM3XOM33P4HCi68XshrnG3
soDCfDXyKxYZeNxvCaKwKgCHUFNm/zO9U2WLNQA1WcEoStj9fL6t43su2SNHVyRQ
TOO2Yxb7AzqZRMdCjl+QW0opKwhAuCvC8l7H1bPvyQUOJF18EZ39/XX5OM51d0KE
ysW3gv4dlth2NG5DKwJMd1Lni3393UK4BltwLCnNHCRs5+K+ePwaZ1VvzKFhnRC1
pQTdvqHJxPdWFwq2rbM5aMO47RXpZPe1Gy+Hv8q6oYJCPdcZbuKdRxie1iscQ3ik
EJmiZRoT7PleRvRSPQYIBkcpOF0xgLkmpDmWta8yiIKwPWMm5lEIAcsfkwJ4kUfW
oP5WosL2Idl8tVpxohiQ/5ugfkrXVGvKQrEs4obSY/Zsh/jqt2q7+C/xGc4rCIxC
6PIhgRkE47hw404+4dTr8QMulZUqa2x5Nfdq/J1KspAaUYJeKlK0w7JeX1sL2wof
mSSeU3m3v5MR4lPZtkg0gWIQIlTXxQ7dkNSwfcHfSRYjdk6Il/iRT5f17G6zfN7Z
WX1HutS4ivycfGiPVhg9AE+oB9kS9A/Emuzv2FsbcrAzoHaQrC+n2qch9Yi+f5jq
d4sxY7fSDFJrC68SNJ7q0QzmHMkYJpH30E7HnNna7WoNbHKTXfUt/cRIyY7kuMKq
aAL7GSutxDfO0/Sz2LB/1wJcDXVvHKSeY33iINL91AvhyNt2u9L7liuYQJ6Dr9u5
HAu3Pqt6cOUBqQcdLyP71UsAD3e7JCsKX16uKKdrjnklU/LPyuSliUQ/3vEnYxws
47H0ZuwdbOfoL37WzSu5y0loMW9xU+Wr7FDom7TR8+utdg2fVmV4y/Tzx5fT7JoB
iqBLpxgogQdvMhDMc8z7LV5mqQxDYM4XqSjir2jeoarBPMxvZmXco5QFW3l4LDKw
4Nj8HoTre//3tHOg2orqtVFSjIBNZ8hdx3aStHzeNN/inNCbUwnynu3d/HSNRChN
wlDY60lF9tFkMeYS2KN9NIuctWPZMTiHfpzjyUVVtUrrgEnoQlFxVEUmVF5jE4lv
QI6Tfmemlow9AoNhcu+HsoX5scP6E96hLAXqBk5uKJkY8qKbRkak9/XVRBVcCUC7
d7Psb7IkBq7f1f3jUxIJUpJKJm5W+nao8Creec7lI6r6HK/uv7ITFPaLqP/jCGsv
ZZeRNi8cun9ccexyASi5Wg4MEpI8aY5mst+bXxI8Ww/HEF8eTw3T/NQpHtoTQYy2
5bmXD9qmSjO00PKkDmmJSSXh0vvHQSHcEppmSfz9VS/k7vNU9lEqdOgkRDk+FT64
hkDl9M6kGkyGmMHDMZ46TpMdZwZX+mNgG+cY89WJWqW79DeqvFmh0DxLCvCunZaY
pzJJv3on/ryciFa4NCjl/tq4+WbNC9ai4QBQWEHIhb4Zp+EE3HPLSfZATWEihN6r
f7Smy6Jniq6MspAeHWg+b4QaDwP1Nq+nxgVNcnLtd+8W5mgrVjd/PWfmx4OZmeeo
UQtZAPcRywjcQLTHQm77DSBMkRbQ9gifOAhEhwJist1QN8X2/KtnWGCNva8kQFT+
gEYJfCv+HRUifwfCk0HLgwlR47cbJ4b3ST2G6MHPLMhrztNf8FbUMAoLoPCGqENA
Q52gi/iOCu5alE/t9CWGSmEHlr3V/N/Pdribn4e1eZ5aUWpKdbMhVerdUAqIS9U2
Q66M9u6dI0sQtMgkJjhrWYVjseGzhz/Of2JS68Bf1astUn7E6gdjYNN63M4RTiuV
kIgbrUc+R0Z1TbYX+zVQIuqVLwv7tOKDfZFaCm3MlsT5hZH0k8nVi9Qk9wwJqI4x
OBYWiG5vhd02iv7L17do9zE5xiudmm3AZlECAqxTol9HntCYTihSVHBzQKIqwJyu
PMzdTcznavo1LfmtuUN8ioAOp4UoGcZUa2xxuaCZqOrXnWofPbt7tu3NNk7UWA6h
noGMXfXlRdRZgPoDnI97nUHcaerFw/olSMZ3hCfwWHVDA5rD0Io7Nann1LKgJpCc
kNf3yhpLYNpzAYvJ9YrnqOISAcVTivA8kcdhJhS9sm/YWqJonq6n/1ilpgKLYv0e
rF36aNKLSmhsWPtigTicN4gXBgEVY4tkzKiTXCyIbubHHNCr1pjEiKbcbChH70Mg
J+1WL9TKZXmvmwXvgR2Epzn8Jx+rRwu/tQy2w/xwzxqbTlGOuRTbwc1+Pi41je0m
vlR2V8OuJUEX9NL8yAk6PIY9Dk4dTiO+x2R2i/Cz0vBKG0/7PiC8VhhMvdP5jZZg
jCLYxaGZrBHUSZhucjdLK3rP7/LHur7jtG9m/a10OUpiCCTqqMX54gNDn2ECqI00
S7YxY/8RIwpHrDdfnqPOmK3VCAi/qPrJc8TbXSLBgXo5LT4SvYa2DNXQdXvMQNZh
kB90MAaEiXd0lEnUVh4sX1184igSMYvV/npC+QJN2fna4XUViAyO7xzB0r8zCZZI
9WE/Rh5nHWdQkePJA6SWfxVfQAx/FNHNrtqGWluQ8TJ8u0hMwqOG5uzxDFf02Q3X
krkNjnC++4WVNf+eapEBeuAWzxJ1we1Pnu5hbVpQoC2CmHW+tdH8yMQMYLA/RY+O
goRoCjJDlTdZb0zcUeLiIjr4RCWwg0iP12xhkX2Rg8XXete/ckqY9dcs6CRQrymZ
GtqQkVO0qKCXJDDRKcehybhYmU5bYKb4Ev4hnSmLD83umlPryWxWllvFKl9HSMSF
X6coTWG0K0PqVNJdAVCnSGTdRDN6oX+oA/PHXiTAW3dJmTSckZuE/oenjWqJ38Nt
mwiyjDRPoylG/0rbM3jFfAgEcG6ldLdc+g0AvZpUryO+JvyLcCJA3Ea6D4w678hz
BtOqEjNpl/goADP1Enw1P1K0WbV8zuJavB0Zf6NDofy6cQCPZyq8hJ2u2ZZUJ7wP
B7mWrlRIGaIgkRl52FeMulvXP9F2MP9f7vK5aq5ByjipOUc2ms5WhQ0abG1Xe+py
bm9Z1tId42MDY4hVo3S3hyGvLzqkGU/7KfTB8ekRkX5RlHTM5OgecK5ZF7qGgFHe
AuM3vD2j8Hjoj3k4kWhvCg8+8sdLriWRmvk8yNg2kyfmEOsYuPVUXqUqeoUGm5TF
EQKhIL9zhh/AnIn6d6q8o6p/AKaY5AYHSEDwdSKLYTakKCVBTmsVWmN/ei26n7Bc
slCYEA+nqQltMW6O1NajW5EVfXGrmd0cCaKNEkcdx63qi4c38vyIAiq/NTszu38C
cb1QVwTjA4YlTuf9jRr9NLE1c2sLsYDXsqcLBTDek0vIkTkBFkbwKRyojGOgq4Bb
DMfUv33TAZpYYrXl3alDW4ui0hHr166B7tjEYiLTHxQFi3Yzai8FmGdx8Xdh9BaU
brAlkoZO/RYny/VAKWVPAxAJCTW15ca80ko7OKBUkNkKeYhLurdoA15uMWqrnBM8
KS9mvvQF1d3p4OGxqweiMQmTlYMsqQiunG/Nb1vWnR7LgiRnK7RmGNo8c7efNIC9
eQbhXoXX8gaVFeECwU2PmkATslGHEwuu2epkMt/RdFOtnNZWYpAjY7X/Cevqqwyi
17mQ3iB3CAL7EheSMKsmsKRmLaeEE9O6CI3ymfxWhcYgMBysasF9an7M9Xnm8nTl
x4wGNtxBW8Pyg8VdF9BQoDo1c5ns4Mc2Y08/6Cz4qEuUjgy/JUHmkDk2pTnTMmfA
tSy7VsWEDGk2GIkgK/MNvdL184Y+SRwgUWCUcMJMrOfulfsaIU1TLDqoJbieWSWB
1CtGyhtbOHCHTfYC1Ek+WgPrrF7S6CU9HuYVYW20yF5/EsL7kC6vv6XXnJ9YGYcC
LKhSQWhF0PVnGYUvKhG9mwD35jZ+OGpQzvnU1SaELkOa8X8r1GaljFyR8yjmlMrK
/BkbqLqgX8M0Ys+mJXW7SzDDTYyYgx9gp1PuMfsVoPZsrqXAUzpex7VUMTRyDmse
Bh3wzhrdV42RZ3KSzHUEZKLr0sKjX4sTqtm5o+WQ+E0CLxLBVDF8zVGKNjybmjMN
E477Jv+8KPuNQ9UE4WPkylHlFW+ntaXMCRh/2Vm161hrPkwSWKMSHwkmnrecscEc
OIcpjQf+ieBBWTc9dsm52sP3ygwXtWFudVZGpMYccWj9Xv7oAJ8XP4ALoQ03sqLy
ZrWslIDgIl9b1BnZbKXjYoCNHrtirH+HkSgmVhsY1U7HbrP7Pv3JnnVjIkNpUdf0
EaL9A8vrD2yIoVGmUQJab4IU4DUjMaFaEUBkmGmAfpMfvHacigU61Waj0qUhovC1
xdxbgrFX6UJl+rNreptEvdIfC+zNaYMi5vxaFSoMPWJoHEYed8jbKA3SBZeEmdPG
To7DXBgX/DHbJXYNjU3b8wze1CGoWBJ10f8RAeGRYPVUGV8f/7Z1lckrVWs/ignF
sSEmrGq4EN3iTEs2Aiv3fiSpcRBb9mGPDOc+ld+1AyNhT+kTc3gmDAtlbmp8sgaP
NAit4rrLhgiSgEJdYMILU7nYw1ljnEFIRiWMvdHifbZwmiQIi3u+RTLDcbtes4Pt
9PQIyhm7q8xGaa9uHqEcadUYhvDG5Y3AXK1O+Tbmcdx+RaTI8/uipzpmAFG6JYDc
U+xTKRc1KmxJg5b8OmJHNR7hHVdKwOfetp/T8h7fCwPvyGGTKYLYBQWKyDagi0q0
/v6o1lk7/7jp8695ugdiI7f+foqD6lCnNwov5Hzi3rptzeRQuGjgAs8miFafc74Q
QwPxhrG3IwGe8W4+7Hc0ziHP903Zrf/BTuiiEgMwPzTc3qVnYNZmcuTYyVtRzyGf
Yn4+UkT7SaNZkT+p5CeGrFLFHyIwVKnepWgNmpHPt/LhALYBcg0xXu0NR8jvWu1f
W5EnVO4zmpiQk7vLUI1ks4EqaB3O2VfdF/m55DYzU/qfVJbslhQ4AVBZ2xc2gLb2
K7vVEqUTXfuWChTHCB04vQDhM4dNxhYvxo7FLAYH5at5miCnlrQz2yQgOFdAOGdk
VN3ugDqz72x7lNwoz2M/5wTarHP7vlx8bC3e+E0kywdnYUfS5vyHAyq8yMAOtPzH
XjaHWB4CHA1dwaqXBHuZoN/Xtu/oHujaoDmsgSr4x4q96lAscKdLfkKBTUaEQBAb
YcO0dcUaeWPAw/EMrXHwF58XkNS185CTQ5pmrAqLGh8UcfcDXjkFsqxVJuor4CG+
xaPOehhHJLdsm743ACkADdO2q5NwTX0McMCdlZ+azLDzeYnm+L58EwI3A1NBIo4k
3ZVTNfp/1omUExjgiO7KrmOcjlA42kJr1D2/S6pPubFHyS2yzBaW0xq0qpUEzMJ/
ftOVC85vHoiY/kKpVC1UQDix8DeDjSdz+iB7vtPjzdLpxt8REMVWi9+qGG/0hJID
aAFobv2h85LNjpxuL7AFFowmwr9fFKqePnf+Yh8IPPsl1cX28nvkec+1bQnmGpw9
Vw/SehD7AYW3U4R6kcfb1LLSfLRHj4nnH/LSiYdi3E10Fv7Ara+HpnSAHdnQ2rAc
uv4Sa//JSZP6gaOgEX1S1PahWOD1972ckHQiTI/mb+yWyAbkwaq35LKKLywgzIAT
qqcWvqcV4wYZG93F+81MEkSQk1KSjv4u46nv814/hN7VGUH1f6Dmy3+EV2hHhd00
rNnZKADTlplrYWUW4nkD5ya9eI+19a5MOgzdBbMFQi2lHl/r+fi1x3Jls5milbpy
uz91jlIl3u0ypGAUsn5B0Ux9Un5Abe1ulnM3xJK0foVQdmtmbQzDl/+DQ8qhkZwq
OTdYhO1qq6uTMl992jVb1bpmARsfPS99+elr8yuqSU1xwn/jToruzdovkKbpUBRw
WJCZQ88qfQW6RNWRPbw1nFunXdH+Y2esPjIKHMhRpOAcf5dG1kX+AgGXY+1WzVzM
HoaC6GYaYe76clbzTfcKJ3uKJkDlZ+NDdRWH7K3Qy4QRwH+jVLZJhiIaYdbp8xkR
3NHwCgd+0lQd5iZz+CiSYH+mhJHwQphM9mo8AO2L3pQcZtzYKL7vD2o7gbk3CbRY
un0PhXLR6Jiz2YgHBqHusl2ZtJETvYdnwe87BT+SeE9vhEWkO4n7zG8S8DCQFDaO
DsBVFMYafi4/R+pCpb6A4a37JIUnd2YT/3mbFlfSgtJM50FcfMM3QVF8uU9/14aG
8RlEyM2gE5RyGZ0Cbod79426oRkyOIxGEblGoaShb2PpcXNNeEgX/fXZzGYLpAAL
V7lES/Swb1oBZgSDUUf/lYB23ha3uG8XCWBq2q1SLn+LLTnDSFcq3fVWq/rtKET9
gZyPprdU60XEmwG6VZInJFMrWozqbp9n0k5keMdRfW9naIdM/62z1FU4dL2al6+h
+WP4Lcp7iZ9dS3ISJDNLRyOxVxmew/Xa2vSI3zAbW83dO5z1mkXvwrntCahV4eyK
4xFeUB4mf/MLG1CCAKfrDSimFRcWeADsU12ky2mF2Kke/cAOJyuvXS7V351bUq01
sXxh3xXZ9NudvttEj+Bc23LMCbIBXc0dqBlFRkSSsA3lUjIzDZ2yUIoa87DthtN2
xON9nfAGspO5BVcxQnA2p+LloN3UUd961sg/HiS4PYuCKRQGULHZWp/TJbF8Ssh9
CIuKdky+ay1GooXr36DH3sQyC25N801VtPRRWB1G4qR7f05Gd/VBsMwHUQSzjzbn
F1guLEWllVWOYWv71dHf8QQltosi3WzI2KFkOWPVlaatvasl1xmx4ELBhwffBbs6
TrxfStg6jD6+GZtr+jQ0JzWKkLi6eOa74/wF68a7UYnjX3+TEmPjnh7dRSkQLiQH
ZroU/waRdZ5ycDDsGbC+c0y0eESi03k7cmTJX+gIPHoL3X3Hr1ErfSNERcoUHrq8
yp235LHqHGdp504HvMhWVcws/i8+Oxhk/N+IVJlc0fMMmmuunvHjGZWhCtRvJyBK
Pot/tkuXqDowdgSVp9FiXj8Lrb5Q77Fvozeh6t9j5YVm7wU6XCGrxdZY5xitaNFU
9oOqrg4rFNwiRYCPqgpNI4820tNxlK3JjOJYVzNUL7+GLRtXoAIec0xijsJalcd4
hF6eSvMG9bz6UKCnFx+3TQ0qhslYL6rTJQ8Ho7NDTS+Idaua9nthE2nWejHf+RkA
SUyg5g1YCJEyO1Rj3PUqfmRt78SROEOnU3N9ZDhN+8J3pQA2JUpKUTnwZ8hmHMuc
xoR2DIlCPDspZTct1TI1ab3Kjz/YHxdn/ZXs8fNe/3O34ZMrsS4tGJelLbeGBF1t
kiuiU5sHge580Tst5bLGSLN9NH/08kuNQHaqKrrAcE2XrJOuVGzJBRgC/8XpjVv0
`pragma protect end_protected
