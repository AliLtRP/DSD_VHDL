// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:24 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
VGpcBW7kpjFqGLIGVjCgfYFrxozRFbE0JffpXCbukMUu8nA4QeL+zrpCMRp4qOFD
w+WyNQn0iJJZm8F47npA5H03b99CvSVZGndawHOiP9mJZbowzbdVyLZUrfePC2dG
nFPTAzkGZGA/1wmiC+INxHtQ3Jz+joqpaViEoH5/Brg=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 29152)
NqWBnR4DmInARXZ7QMplzErqcZoV7fskXiyvapYKrRDh6ElCORTCDQc6d+OozVxx
66qjB9FPpyOz9X0IvIXOM262H8KzsrsOp2CCUOlPsPMhBnPRqNzHw+qgXFoOnIIc
oLry7Nkoh3qnO6qVWN1hqgnzHc1Iq1sNpmZWpVyhHMsB7aRhlf8eQ1bQOBc/0iaj
TgqiGjHs+JW7rPzVmOPz97D1Uc3z6cQ7+G1HlZQlPU9v3N8VDKrWqIszShDb9Cu1
gwiVIB1ZECXbKdiiUO4skM+ZPWYp9lBvHsObmnc/hkZ4wBqrQrOft4/fUoHbzUdi
PQHzqJGcSoVxe0wQ7m8oMdGZcpQ1nzdj4FS426wHsqEVFoQS7MXYDdjRdJK8AEkY
csUyRqtbyNtUa00PCjKczvyzHfHhNWXkFBRjVZNkzD2Lnc3pRHhH2xvSncUrHTCF
f/GgRc4ZYEP30NXxhqvSpvtrBKR7MpF/euT8cu1cgHYGtOErV8MKGCe63eGwAnrY
QD3busNrrdxLGfIra4HUCccUF3UH7+8UbpO5mptRL86pxuJUZbBRUOp/Qhcy+IOb
tzcjLQWYbHPrBjXF46s4VOKV880RuapElVLR6jITzHLdArKBfK8mQKuLOxjNelp4
seMazJWV8xjlUplFNuEnGmg99pW9pTL7y9i/+ibRjCkjRcJY+q6yImq1QWUmOdbA
khJtKz+g+J21yPRXWnRo2mlA4j6rWrf0wyDFCtVrwTnOEwL8wQEGl0pbh3F1Py34
SWuxFkVjNNp5Ox8DjBlKmlt678W7eFZxyp4RIk3EnQJanr226Wcl+VafPxJ23jlx
vpUZnaYQvORItkhSSscKFB1+mwlrXtUhuN3QOF3UZLqFkPOl4noKjLsRAvuNwNaU
CDwZJq1WgOTJB7pEVpmBGZ+12guCpEg8mkpBRG7kbYK0dKV7EqN48elQfwYS9X6Z
fLm0KgUzzXVLOgRfbBVpGOeNGsp3IqUanIsvK4ySt9CK0XsXwEelQNzKJ3Sonf0S
mWcS86wABMh7EgpU7koIXmAGK+MUI4eJjT654CuveYX0ShpKAn9uB1314YAju+SR
ec+LiseVpI5OppGq8bED1MfkG4e2Hu8DNV6dtEsv1fXV/6rD1AWjHMHuBJAHHSZs
urUaBWMNlOHqULyfJn+iVauZ+mSuYkROqGkSdhKf9BgnzQIhlKoyhx1/ILF/OhFD
/BVbfMQiE+43PfiZOba6X4yYyb+Y4Gaxl6l8UDPZp25zYuZ3vup2+9KYmiE6oBW/
23cABzxNXPTLoqW/QZ1AEmBb1DCNzofXPpbeppgR3RwyD2iUg/y6vR9hvkf8Abib
Bkv0in19nORFJkEHQT0zYZL28RlgEp8plKMAajSx3EyHaGf1BMsp6Au0ROy9bxKt
dih4ydG9YCSmAIwoaMucjOQsDSna1z1/QmrITZeBmUJtT24C6ciKR8ScCo/P9eB/
ucofzyEde03/VWwHKJeAVL3ewiGyRqDnbj5A9dw8Yr0YEAUGu8djrjLTgAOayUt3
GDmWPG5mPP650FjnImPcDQ4YmEphhyV/S/SXqrupF3s9BCq0AJ9gtgC5dEe2GVVU
aKooq+W6HEvJI/pnAg6JmYn4fSxgl9EJZBmlBTaSF4smWgtZgtOnn452k1cELnwO
jKjpESrh2EJNAhm+gfsAOkLtqv641N26WGKB8fRAOZWCjMP8xFxzAxGuNJRzYSfz
RbwCHjEcukv/uHGYfFU9gEGXGqWfT2S4aA/UJh9JGt62+XbSuH8hRc7GhdUQcCc8
Cl4XaRhgpRjjJrP/XfOdQxV10U34D8WIXv3hVJugwUFPauBBxn68Y+/Z4x1jtzA4
a9MUQgWhS1+4DkOQrdujK3MqtAqmK26SaLEK2MLcc6kpPvsg4GhZixnOW9sDESXq
VHzG33P57OGhX1pxKlahG3nU4namXa634fs1kbUnxm+vZ4JSkNKRA8mPVzdiWwR/
bVoDVXO1+0nxe6Lw/XZIq6ToRprsMtlnyrdSouGbnH7FsI0dwE5p7Rtpci50fLDc
OPM42hrhPFVuslIVkd3XPaCkvK/v4RxFNzVV4nhz6D0Lib4uN3qmQgIG/2neL4rn
+cEyW5i6Pn3yF8UVZf21TD4dbp3xes7riwj8i1Oyh6QkMW9U0YDkbmDog6g8GvLw
XEsoYMlMJTcV20e3pR5Pyj2+crAwxdPWUeFG4yKAPMmo4pW2Xib3uXqxGDR2L+gQ
ua/Ox9Bj7FgJ3iMrbG+AHaAbliYLUCbzcfl7FZfH4Mi1I2cCL8hWGZ8apJbafznW
6LzKWhT2tx5OtysOrSSeRyR0k6a+gFOy2Uxw1pGFMRCFIyJFPYXhshpC1Nqf+DNR
7LysbliyVDR/WPD/P4DO6TLYpouSuQiGpotmn2A0js9nU9UiW1TZ6kWm9v6K31pI
r/A3y1VpbWBU5DjQfdPR82STHNaHv287gkysIB4m2nrrQZZrz0k/Sj36wbTpfg+q
oOSA5b8ypR8/JfZNv+pBkOTRL4f3v0dsh0LtIaT3p6hj7exZafG2o2DOHYDR47yU
0XFxRrUMfIl01WuQTKt4fKSXeBvr9g2Qm73niiMluSb+iQR3ux63S9vkJHbB9hOf
C0PjfR7xvcTrS7Wxr8G+9m2Vv1tG+73ECFDiIhBxlNN6jpkLqsyCZKIVkdOVv+EJ
+GPJO8jRHHxT0gAhFE9/2DU/9XebG6bsY/QfFeVqSibnt9+EhMM+DWa74o+NJiEZ
xmLIXi1o9xN73KQ3xney5/7tNfYHVCBQ/KcuevmRT7aMm2L22QXUiAr2L94/M8pN
sYSbIoMcg9fksHrW0Hy1j9XpYLUUAjPc6Nt80mZcFxH23gFAEpwJIFyGS2T+VlMC
1SpayuLaHXr3VvYuNRD9v+4QXUYe3xpa/CKeNroYd6GVxnyCNc6BQ3uNoD0LMIsH
dQbfrsf/GTA0ULfK8e8M6A6pRpN0ceGMsL9NYi/DHrmcHw1NaHoyjj8yMI8bq1fN
zwrVbBZ/2spaJN9pRL3za9ySbzrvp+PYIOawX2Asb3cyiHmaWeotY0SH8YgUJAW4
Cs7xIyQomsi8YhvVZx8nTDrkodd9dpyVwU+nBXxf8S9RsP79+0XAiwpBuln9mNIS
BXkgbSf+1pB2OHWOJ3vc716z1VkLp/IgjqzM+0ZeADb+bR2z9c2kdswKn4yPlhdg
YKyLn5ijQ/WuBMCkim2LYULOXxbK0u6gerBv8tfsxU0SmD86p5kwUY1LgUvl2ufL
jjWMWM9HOymeErupgwh8d7qBdbduGlRDT4AgsMOz46EUOKgnNGJN3EmU9WwsHEyD
yJKtJJ3axnXqcQUONfleVqqbjgP6vrRHQD1RtKJ2O8h59TmHv93z60RefBjX1kRi
dg8BU7OvgjmpFxwd7x5QcWnNNcXfU6ucP7HBnla09pHrurcQ7iFgxy/VUh7iniAz
zr5iqQX7yJ8ltDtusK6TZZClCaEUpx4EjU15MW8ZSQXHjWtiEvBXEN8I2hOl++PL
zNi9DqV3obsiKFQYDragbDVy1PQmyEHepR10TCoSfeKvQnXuSt/tEEnJ2D9oLR3z
LcV43HVLRzjY5svmniGQ4Oo5lH2R/VCMdLLm5Mr2FWpw1+NO8cg+fdoHnOj+QcgB
hmWBeJhDG+Ptu/axx62HfSaX87bBQb9zHMKQEDLf3EUzwbelBSdsPLUHoKbfJb9E
bdFu5URMF08JTi0g4ex1NMm94I+/o59XCMl5F7WozmSMym/RCHrhuXeNaz2yUdGv
ZAobzFihZN6uHPL1v+pgnfdIAtyZSC3Y96n+u9dpFW0dfWkLAKfC7qQDnt7pvY0r
j0Nzm4c5lcQXbhUS/H05OQCIfYlX5Ai0dLkGrUMgTW8n2HBuXtW6PF7Z0kywj+HW
qDB3PwXIiAOPOaXV9bA+2t9PsQIr9DWA1ZN5aiW+ONaNwI4ZANUSw5qDPaaTGZOU
q+vQJuyAklvUIIg5QCOPJmcvuJbp/5za4QCCL07fq5LlPxpGitQMSuv2V+ZyFHj8
TCqjYLPz66GHL6QgMz7m5zQEbL0EbaiSt0b8DO0ZbgEilcHoG2jPJYaIJyWiCjBR
5nymtIi/SCvlWlY8mi7WY7FHadvIq5+TF6Z9cWsPcyeLjrcANEXy3OIiTEJk5TdG
H9m2Ox8CKEQ38wDn+J5/Ktlt0btXZRy1IR06nqtEd3OH+YNhUs3a5wFHUGAW1H/P
nnurjKhXbLHRsSEMiAB5ZVP3Ag8i60eXsa0bkPfHIGpywJajyV1IzyaqdwNVfp+a
b4KkFJ+WDAlgcbTSrq3RoXocybw4i6AxMvXj2C/U9UUFnZ2V6dfyQ+ZP4JwnDw1x
PfZE9ayRrwT8V2BHqJPl5n6krbRB7TnIPzwmBagD4IwjLBusY+9V33SwOx8Gd3xW
YGKMtfF67TVWDtn3CClTm7wx2NFPAp6rsSkw+V+U5dym4AWsJbBoGlT++KPMByXf
kFpKgRGu+9AOaUL9EdXGT20tRfUy1FGQAU6R7O2JdZ1xf9h8WB0XSB9zUqrQs0FI
Fwz++99Tpptq4cw+hOwzli0ZzU/us6g3hBbH23NOASa6jJNCq1gVJwIzhNKLNgtz
sq5/9ojKLkg/3jDbQXnPGuvZmlZfcFV0Gh1b3r4HrzutCBVU4rzNPWqJ+ZEfD2OE
oCfrxtsOCScbvNlBDmtZ/alecTRzynx/z5aV9lzsNCOV0H6Dj6Uy43bBgr2BVoD/
5LajB6443wFh7bnIVQHdtC0zU5/xhBLBeovc7JRngAoGNjbQo6nTYyb4mPKgpnOB
AM0AeH8mLzHQkW4FHG1st+Ahel1MT14Nc4KSuuyeybRkWSLQAv5RvTUDIrgE6BDa
bVB7QcCMwT17DgS/gk/KSFPOYh5K11JOgVH55EQEryxAKq/WuS6wsohSyIee68CB
CoAea1fb+M72UfuO+SP2RmtkMg3st6U12BARJZwApSwW5l8m1Iy1vtWHuZeiPf9c
1ExI0IRNs50nB7sXacRXd1ME1J82f7jWQ879TLIdMPozNOC4eLOPkFtbWg6MO+Fk
pDJTrE5j3qi9muxK2PDNPjy0PtkpOvMjzAzwQedI9y/ZzZ7fqXLR4pF7p9bwLmT/
2PlZg68hhB1dQcNCpSBDZQRq1k4P0CI6ovQ7wjiAgkmcxB5A+38bOAceuKP2FeKY
pdXTvv4nxOWgurgK58rpZiTsXwlbvSf7LXUU3BjnL92OUZmXVdPzROtLyitUOQaz
WTrbeA4gkHgJypdYy+Zo9vadaFE2Tvpk+kRociNryc6aauZIQes2rFALjQpL2z2Q
N4v43H4P0J9mQHmeDpuLcOAzXuga34qagxGJyA3ACSY2l8k5JpEUvIf4mlU4JY0F
zBWYm9cwBXD6SI3LE2AasUN+lC2p1/d1NakcQekLKD2KfrRSp2vb7esCZuOJ2/l1
z9YP81twDhYP0J9Klikyl2H0KSThjAnVixRMejUfdS52RLW0uW4mtPmivWmk4RUa
jBl9EDQci+jF2op5zEOetOY2nBrzZXCmIWFECSAZbC1XmnnJKRPc5AOQ0USBkUDW
vW9tFJhjE+eKtKZF468TSsxgTMXFRW7YZoMY8HKPsYDQJJKr3Hl743bGhGWqy6gs
Sds4qjgCuLM472dCIlxbdL59c7avUVZjRxv6hhyb9+WMLzgQk1zyuUiXdFvOCtYF
KePeGZnPpvMz9LMYnmZqJdvBmZkeB89ALHtq5Z5S8ayZw4nluSyfjy7FErg9mmKy
NPAHMO4w+ZB9vjAnGuvkNKwhLpfRn0zfdox+cH7dirdNiArIxz6aceLBNPYj7um1
HvKOJulT1YX8tMy4AaYLtBj6sfBT/pK0IY7BUzQtykJElmm1RVeOgl8+Wotnnmse
1tAg9cHE/bsoDdRoM4PQ20d8t1VU5p7waqUoXyEtm5o03rUOtOq/IWHD5GOTmHrN
r3VJFz6m52M2JJ0S+HN3RiznTQnBEguSvuv6UKkpYmyF4QOqTnga23RiKYaIe9I3
Ys3pJefsNOzHhMrR5LP/ntz0E+mYEAVhzZB4HELDPqw1U9WgCEYHj9iNcl6tydjW
YvqWjJke1Y/03+HUn8KGA2SYYaLS2J5z4qJ9r6yp6n4n/PWa0rdleVGNfz7C9aEw
mBDI48EA0Lc8Y7XHlD1wJza785ZwBDOTpU9+bnUyWWI8NvmYwh8dESp7jSYxiYH5
1q+Ckc8V6lqLiZOMHvgdRfiQaRXq2TC7zC6+JKKfLWpH5ToCARDIrst2VE1g65GI
peOLs98oS1TB85BRfuml2qoP+6lM12/wvXQoz3gAnjGycqTRsEbAxFbi1MEJfnV9
7/6F0e88qqJYptZPxG2XRCroXai39XyqEgYVBcxAY5GlFnYc0g7phXUXL9+cau9i
JOErY442O6Ft/WlzeLMTNNBgCz5u3uDoxmzsSXBsmUf6xZgBHvEn6w22nI0hCf90
GYqSmQXUS5G6egOFfKCB3VkVcz5N0SL3jcF6d8VzWAJttPR6dseFt4jNkV0uU2xN
nWjxTWPWm3kpYuMvBfAKH4D9KDInfjoR7uPf98ev2dXtQmGfokjKXEZSwDrMqfp4
jGwdVn02x42uySJGDlIhexyjWr/lKJ2X5VmvD/vx6BWhItMR9TME8zd8FIBrgkqa
nhagZZH0BKHDucLCh1hvLemhq30SHa5GUQjQreIBk75++qOWkWVDWefdsoQWlsgu
omMbRgd4AN0uAhi/SSov/XrFtVM51z8gb1QLHT3paO6yRacYLD5WTUp6VvYy2Wt0
IjCVMBVpH6wVqF6MaSSC7hVwD5ZGME7T5/G9w8sQnSTs/Hz94gdIpW9hMdhe9BfF
z2gbUPUyF/5M3h6ZaeZKOAZ+CIN70pGafbNRA/tohC4qZ/qdoo3q412kbZAKziy3
eSEMPdAlx0goVErWcv6OBIb5NJgGwr7KYBvNtbG5Q2nTNdHotlSdI79a4avCCZ6x
pQxS7aDrh7WEfuFnNw5U6CH1Gp6cBy4m8zyjIwuWJhrZzIGMGwhKYzbvmBqZ8rXh
A8niEzBmSocIqViydHAfQ+spUtLlJ5hf86Y6RE7dN4p73u8jSWcpUMVLC39unhpS
spMALcpDj79z3APE2GqBDQUnc5v2bkCSe6ylXlXmZ1Ps2KoTG7JrTthVUldyJ+Wc
FYywPBH4QWQwQLAEaDa0zFGg3XmCNXlFO9RO00LIIWgBemOmXSKYEtRiBfdPBE/Z
hcronXr6vGeJ724GwdWTeY+S1TifZhTM4btBpXiMzdkL0kO71h1lcCa+j9vxswMj
SbqfFlV9+c7qsNps3iK19pmZp6qfnFhYqe1qQKcA/rml2rVeAgeGTbxtxsAMMywO
j2K9zz7g9bWshwvzca7Y31/+kes4QY4GFkyZfvKOH7RvVxHvV4BYByJ364wemw6q
p4PMqxUkMufuGFDQAgvx4Z5q7Chnq1Dj1T8wjh/uLH83plPIPSicgSFQlyEbDPVb
kwTZigA6S05v+SgYvXvr3F5IMKYRrJfwcpJcXIGsVfpAqPjTptQsMEDRA6i8VAPu
PFrRKZPkwe0LB1n2+4rgn7MCONikzd4B0u4yj6ypAC1JEpsna65VrxBTgLHsX0P5
BQ2Llwb2NJ+prBCG1AByAPXg/Xu3dcPpswbGl3xddbTeId2vy4N3O0nyVn0EPHWa
+1pkjD8TECE0dcW0cyG42FMxH5X9BCb4bFRecmjOr9nAOKLp3Hl7nOCuPxTGGRMA
5H15hzsvovrqXAV7RTfKoAvvTFNvz23v/mWzf3dIQxQZcpt0EWG3VF5054Mb19Ne
9cEWvjwJv0/EDZIsyoFtRC6OnvrRx/k45znNKdS4YaR6BzzdqunK8yK+8zMB5INB
D/LoOOq9pApZL+4g7IqHJ5JhSIk1cNzhbva/yu7BeULf0ZhPfwXsaZZjhUpLZySV
DPMAHRAVW/bcZkaixGPi3poD41kEanNR1nK1Ou/OlK49uZAb/S0BfTPFNL77k9Rb
JpbL7RVd9joEnLqzwzzSEUGmgKMYl7ssb9vnMPUju4/2EdH2nX/oxvT1xpfBaO6X
US9bGHkO3VFu9XEBacTvJF63oWGqkBk9sPrRyaZSYPeQrNu3acdw6JStHNz+cpWR
CX1TqpAnF809KlXGuMaA1qtsp/pdKULimENC3GihHjQc/IEVzx56qljdZ9pUtYJ5
zm77mK8YTLl26c6ANjvPqzSy1Vb6v720RnlQom5t/fw3cpKNO5mdTudnH1wadSsy
/vLJRdVt9k8Hx6h/iRk9EvJ4fg+KpfkqDOjkFycoCT23XP38BHlFu44kqErwSuVu
px83eoW65QCXeAlqMnbKCXQi7NZbme6bcHFBWoui6mnCMnBepDaUDXy0akbsKyyb
PXidxpcieea81GMZCVW0VIQBzh89v55emoKopQ48+zqblGl/nr5l9hX0rjLw6raU
DEkYU0R/Qp0qmxoRUbihlFkA8vMQOy9rUJ/L+N/DGVVbAuWRW9wQfw+SDnsPIqfx
D4M0S3429WEdH5AVPoCb1Ltu/1S2fTsPRYv7RTXy8xBglOt+gpqRkZIc2KPP1BQF
aggQV45WDRXIq9Wh9tHW2Px1lrN8zNKhZ7twzhWEvrQ1xAyBd5HNfBRFpm27yvfw
1X6DoIa/UN16/PKD1S3V4hOIgMbpIZdkp9L7MdQOKVyOv8ED/+IU5NZY3K/hf/4P
XMDkGPBU+2eG0cvSziP7fihekaMT0+DEYrWprDO8xkrSlrY9ll6u8v3Ic7RxzlEg
Y4DCSJn8FSHlCjlsYMCc0narLPDtmEWX5CqLJle/p75nxLZP6OhU7MT4yurkjR9I
Ntm6d0iQIj3OCpK0UTQ0sEc+3jyY94y6H6g9EhkLNuPpESqK0RdOafaK0zesyNHb
ANyxC89DGHl0bfc/gqasFXYMrsYEFrr2uitO/BIYDiWKx3LFyqSj9cXzbX8WfLUx
L/uONY4nDxWRmRRhGrvfUlodr24AT2UC90hPdwLHo/PUVcsXt6k4ZUwJw19Z6Lze
Ohjv2JQvWexJizkX6wmiH1BDOqbTgCqjtPM4ooWXbpE62mjGm58iU81IVF5UpSwN
SHs0+IInh5+tLc4wGuzHGBWpf/z+g7zR9loZC6D7RQnqiWzM0zxYwkZ+F/GKsVEe
NyeW/zpQ47tNtsaXSTiWoBP301eDENskKauINfYtmRRQs+6aouw0u0ovb39pvAnu
1RhWYNIjHZmTxKqKGzfncyMi4oe4p/zJrKhar9fphBpRNIYylN4WaZlDZsGFcSir
MeyAiECrOYJ52BDHw5aTHwSQx0D6VaNLOvHGAvaL08qkgBxH9pC4HL1ncM0F5ulb
A2WsZS1zCzb0NxngQiEr0mO+bB2bNFQs1hVMc3d7CyXIZeHgVI1l2tsalfhNQ9rw
wj526DBvVdJQG8bdlHRR0RkZsLXxq+cbioyZ1LkDNs5IbrWpMWxL7hhSYnGrJPDz
vAy1L5O4679fuMrfHfd+rldXFihrRjZno2uPXmNzO+wPbwXTJK3ZWfgpBAb1kDfM
8JhTj0cnLzPJ6YvYora99MCL4qf1X+WMci2LEuZ94xHsXJ9KjTcunCQP9UI0Wz1x
SPE/q5CZ47Dvw2rQ5UQS1W/eYuaNs3SbbT49m7zIReURgehYsJPOsGcpXtjZMPzy
8mrGe4Ss9zM670rS1KTrv9VfLYcBUfXl/HH9hs2DIdPzRKzbwT9cDo2tHfrGoyXX
XiEK0vX/2I3b+tZv52hfT4M3yjTSGgs79WbqzupiNYK7aVpj73jN3hxbFhOJNG/m
lqCAyt5cfA+CAlwgq0DcOXc7Gzh/2dgSTkDW3ZE9K9Xt4+hChfu/KY1PVnwCqtaW
9cQPG/vBEb9DA5OgsA9MiiRaHST+DT8wfwv9OnUck1jrNypYsYanBN3Vk5Q+k1bX
I5HPtsikqfEsmwjzMKbjNbQPubUVonKo4Gxk1V02N9eKdBzAQ9ML1JI7gPVZqVQt
/Mfk89lxtzHKKv2ad/ZB3V+NgjtuBSP3T/uAQPrrt0/xDeXx07kBe6khSaZcrwfb
If3vECHHGGeoQI5AhvbKk6JHoLpjxC4Gp5gSdncQ/mgha4iatHzc1GbfODD2YOKJ
Z2bthuhZ2IUk0590XzZfSCouQt00xXi2dO+Cd7mppxbOw7tlgI0KggnkJxUBR6UQ
YTM+OF12JaM7yZa2S/GEHnGw+f4//8IdW/km6U9Wq2wqWskodbKUHgwuL3+jRdrO
VY/Z6AbqZU7IZlsQAvCWvqrlWWiMBDRcwwaqyuTxzKJwPvMnaX6UDTSAaNN9RgXx
ono2OXCfksXUOjWDmbSuXwra0SwKcCgQHpGNB8uy9Ks/tc+i1Y5cpGOwDRqWdPDw
VwkZKIVja4ieL3Q+yN3/pbz2ITGts01XP2SJR6SjlT9Z9qnqS2eMuYsdPelhMjTp
P27e/P/QbwiAjKwFEqyQeuCqSG8y6+6zKFEq9LzlVhn5yZRc9bQVRevBRz/FdeJn
bjN99C7OWrywwPmSKGv0gfMb/u9VZeo/9ijeaU3570IAkfBVo5wJCJv9XoDDSDJe
B1j9qAT79G5Du6xE6ypoDCiT2Vmkn1CI+iNioN02upgCHXqIzWQufJaig8K4hzQB
rNV1k0K8QlAM5Kq3QuVQRMNlit5pKOr3qrcKBNIHVmo96h3D/HhiOWtpQ9NeHHmb
uZby0Uveojd5J3nwEy9ElA4eMvlX8DeAPJM+2CL1oAsxxStucHsCzK1pQfqfyy64
HEbkHK68UNbKpkuIEeaYIlepqNNgyOwVlYp5htYzQbFrfI6tIFhIOpP1Nt1kd4vJ
qJ2E8/jeSWqHNNsjXE/aoHlOrTKGs/zK6/Lv9DB+mpUbGNcxmQFGEyAQuOiFOy1L
bzvAnfgtCOTq198j631rrMbH4kncRP4+V9BDZE7ijAcLqgpsajaNUM+vmXA4xW3r
n6UqSERDIeFG2GA43wbKNWkb4BmVJjDDBtom88To48xQ46OZ8XP0gdUAfX+LIPiu
eurq2S5g0RD89HiRLiVhl/hwRyavR8+DENBvHpxrR7yYmuankEGLSPf3cDyYhj8Y
oldDQ720w0pVD34K/lZEZQwDrHXl/LpUEPU8zrmcYU8aoWtQBU7BiyaCt7rjRUyT
BrFVKcbiZquJSttS3cB0YUJRfG4ysqfiJYlcKEEPDhcNB5/EZOFYusnimpll39hY
FNeW+iGvKQeK45+Zu0Lb8cCAcPRPKVUsEPY3l+wXGjwMaVe3/Ic7UF/rWzpKgQWU
uKocvbowPpjaBuXXUgNeI9EEoabM4JWUnWlwjMS34oH74ddc6l7kyHKUzkFQvBnZ
sg2VYqSYELzEo8qto4Q+29lEAl6T87l/25goMc1uYrDOEhDR9f1t3XOHztVx3R3d
7yqYS0WEhvFPoO5xTPrvJYdwKEA/KS1JwjTjAXsrxn3rVLOleIST2ECbLAg/x7tF
/b+h8TkmhiCZhDbOc2i0CPyG3kj+zjzNRX5nC3MNHEGDZ3wEjyEQgkwUd0dKnq/7
FMk/HY1xSMOKIb2+IImtRvQwwBi39Uuv269HVn9mCm2SVVESZccOHRO8bRlHC4vS
14FPUF8/7wjw33cgN91Hgv6EI3GJjNc7drD681YCGeeEqpWZCPEp0axcZRGWw48V
uWXgpE4T39m8dWHadIEOOuBu9zKyrqwJYqwPv3zTf8Zq0Jf9MhqOd07tfnsAONpS
d+Fp3PMUSLsw4DX4vfRWbLu9QRhbu86fU2+IdybMeBniJ+OxI6gyoZjS8b57fzi1
6UG+lSLVs/jhuJsyGiS5aseDD+pzRXZ8KR5xmBdVgNlBo64gzvYLfJb9Hoa1ZuV3
bzgmeNjvbpSOjFdSvtpI/ZrJi5nk22nW5zogJ8OGLtE8h1gMaHj8Zypx52TeXPgr
ZywW2GPRhIWUze4KotUPixAyAM/cLNF4QiCdssbvFDRMCYjqIQJAGyW2nAuyk9Zl
9v9gaAh1zc6ccMNnDamYXIC1OroWcA4m9aDyKFEDx9o6GKDO+2hk65pnw2owZlfF
PFz0Bcxo+0aiQh16/ZuQR47EHC+r5F6RZQqKYiROCvDa0Hn6SjDJ700jC/UbO4cV
pjYqo30c+PyPV2jX/OEYRXOf3W/lP6/tPBNqe3ZkyvphGtjg3I8IA6j0r5QZLSsw
qpq+qSIhehYOtXIXq0lA4uC8PoIrsMnvgfaVOrJ4CHnP6C49Cl98/C8DIiqJK0IC
pk5XxPE2klJUzPwxWkDCkvDXn3+dk3XeJBhkMQX8sU1HQIt4gQoh29t9HayFfp4Q
EGN1wvPwvvBLKU6IWaJhsdR5oMZ57f9Llf2zBzt8NyiNDNrVRswSfD+VFdnDL8pU
uIFPinBv+1ENb4H0BfYce5zDhYvy0oCD3LOseo095dc7OddNTd6YiTn4+/MQGISe
pC8A/3lrlEA530bLTgwl2z7QaddC/+mxf8QQ8+9OHLKmqlNpLyf2Qfo/yHH4Z0mA
RkVVCunqkdq8e8+XkPnRlm3ngumnmHhjWwU801/Fyf9ntaZf39XaRD7GvXu8iksw
2a/1jgTKP5zhrHa4F4kWBPewVufjUWgnLSoTR388y0cM20iLvDV5V2sOS2WEDPLI
dD3m1RDiXRRwpb0jdGIRQPtgPXfy5tbTvJkJo0QXNTBYYu/YlHo8oVdZKrgqwGRL
vSczDmEkJiN/EisRQGh0er+FO9PFwVhI7rdduiUrIzFJOYUqrknAG1Sn0t5+N9hf
QRwxBqPQQjaYY9oKXarddHIhduTvApvjST1q1ukbLKaXCnpAnRUzejMl6gpKSKlZ
GF8Q6XyY3EtWT8DCjpZ8trxK20QQepVwsjJHEmypyguLZrRvoASqhVQzFQM4LDGK
MS15HnUiDpZGAkqe2ZDOM8z1rlEYuDusonGdn5XLCfdWZ93j5qRJZ29n/yfC++2x
cm1nuh/B8DXJ5TKUi7lIOGXwHHmu/4Y8ehIfffc46zvQgURkV5onEW4bKFeaB2zK
GrDWv7nLkqwelWvcYlsqPcdbMuUgNCEQueecWyj3aUfaXumjBY2osse/483xIv2j
Fk4DmQ//Y2wKeShtQT5HxyazraUVjo/iGVIMZimSJuhq21wljIB4Vg84iQjbfNcU
T78IYcNfTi3ex20xs2htDZ1Mi1jNx7qRbNYmgSiyTytbRBSiMrMvHlkxeYMyqL+u
OUy/2+fecjHtjNkOi2mlb0A2M3GDCmjxT0rF0+K4tJE9tJKU91tayXb64piCAITW
lRuEz6HMzzGPcG3Xh9lIw97OM9VgBuB9pPXDaQoraO75wZrJwrBcIQ/gGwnvFFdx
STqOTBaj2Qui0FmLQFhi3NWi7FTYfTYF6gCzlRm+bX2Ygnq6rpub6EsTt7NwOyW3
nCahC2XPC/e0wR79TrQ5OAkLDizEtI6Po8lvYdsMLK7m4+o60ufmm7UKj31Byac2
mY7SlHttk6jpMtc0N8k6kCfswQ61eiZqHUhue0WftIPouRZfQdYMo/ERW202fTmk
4Gzmg6qcqZfFqjpFur9yTV6tMiyJMsWMKY4qgDGJPT7/Q6Ct5IppZIe17Lip+mpr
3p7rL8EdbCxzZsL+nLfvZboDS4cIqpozyT3Q1PzvF8E6IO7XaizkueuNuiG1OyBM
sVEt3Z+xC7BCLjfVqY9d6f67IJSkzDweS7cMEQVSJpi3KGyVFWGgtLjjng64nx1r
IdGWuwTkDnwXavhRQZtG7EnKoXE3FspyJzjUzvEZfHeDkjNZNux5eAPa9Qt0AcoH
Up67PyKUu6kDRfIp+6+DOUXybqbxKBaLcavN+Cb9HjlJjiyzNpRYN/G3DZ62+Hd6
Q0J5hLQdpAF1A449O7nZo5GtkpFqWnLe2vU/fyUz3WA91kSuGlcA+6WZjmKhhQrl
1npZ3zSvW9eJj734fYPoeCfqGgZRIpfWAsxbTnjseqIjIgFH7uAAZwvI8elpTdtC
tRX0czvSMIc9UBbhHF+OZTQZ99C16uP2z7vFGQNCIhMyWq4nePY+y5EEChZAJTlO
t4ycda23+NbBcgpFXOe+NeK2WGomQJfyWHVEVRrIDyo9ofWR7isGdiW/13MLDK0+
eUba0ed65nEg2SzKz8WggDjwmraRj1oai6DK57sLDp+aP7a6lP0RGwn4enqZPC0e
lS+mCnu1KnyK6090ON8+xkH48M8xPCFv+dvY7QC8KTbNyHqabEzl/Sivc/EyV+Im
giLcH0iYj6hgDV9eygt36JPvxh0uMP8/4t+Y7HG2gsua7mIl4a8FXMejhr3QW0lC
4VixreekANwDkmCZyqRHiGdFWLqO3gSK1BF7q3mCIrnlExgjvbklOMUT7yfz3wef
x1ubVPtMAAT4Z/js2tMNetbWhD/yRUUHXo+xLdMugIEXt4rq92cc+gUmNw8AwZ7e
/2O0axXKwgX3dYjR/f9lOXw7bVbeZ1I1e5+LQNtOgN7cmTx7H8/24Y7CT/71lzi+
au4uzci90e9Eg1nhDXZInM+MChbYHm0RqosSjBV/i+JB/kxuD6x5llCiZAYxTaGt
6c7AMWg0miqvkCHf/B+hy5e23m/hfuL7aGLOqqMtofFPL3FbmytbCVfnzAGHg5yu
r1UP0MKppvd1nxov5nbUXFVdwLWbrO8tlK1qJlwhRjpBrcy6fF7MTnXM7EM50Iau
JyfH7lPOJZ7eqAPVidRd/Ruy0hx4+jQEIwasP57yJ2PSFhllI4ddP82LVEsSBk9Z
UaDMytzEF+7WMcX1C47N2TQ/R9Q1gYiWdnkGZQproeolfh2TjXPmXD/PJRkPpPRr
RlvjAhHr5G/j3+vJmMeMsjlYlGWsMOFWPGArychYKtzkE43LfsKYZrwP9nKckjtC
tcayEoYX3wuHqh3wBSWVxWeFyI3r+KBlVL/cSi5yURLHeV3o8kLt46hFV4gA5kYq
dmpXxJjo11gekSKmCOHJGEhNc3mPhkCfLUYSaYCs/FsFZzQBd1WFS6Iiiaf6CdCN
W7YGTjxY8c+664OD5cumGEGEhI4jsLfWwiCGeBcN9sDK2rE6rnyp5X+/pbI0lqiO
qhwr2+bjm1464qWEDm/6Gxjy2gsG6SsTa1wrs+rUtz5ap6kCBVMHmM/3xZIh+GHJ
wgIRs4VzetUZftnR3itL0kr5kCl8UvVAu2igJkiZdgvanbw2seLjhq+uR0EZpb30
Ol884jJOmx3IT2jOGH2sozUAgil8XZoU/XSEHW7unYDSJ9y9KYnBX5chAnegiZ7k
bQ+BHNJcoGTOW2BzWaMcZnq5Th9bpBzeo1gz6ULf3uXUpRBgC0KZOsPGctNbrHX8
HPxsiw0AKahTp2LuyvXf7nmmuS4VH8q7kzszLt2IQimD7jZJqOrbq0N7+4d2+mVo
+zNPi6at9l1LXBt1zADhX1KfqrOCZm6oNjes1l+CDog5TuUTmYg/JkA+CfD/U7oP
xzlZOWoJXtfOF7jePTbWMNQCx3A8LQRSlPkk6I8Z/4tQB3B/wPGtcnnNJFygU8XU
5jScqAtc0t+1JqjJx13mKWYgkmqRNCK0B9mFGQJs8AJHhBdPkimZAi89JuZ293Fq
H34sKn/ACN2HOtQs2gT3IrrZGqlzr+sN35BZnBG746wOZ5/6BHfbEBkLLmZakMzq
BKCDUOA/vxk6Ubd7Nam7OwdFg58HDNLS2wLHzEtZbR5iBn35kLjRLgf73IZbcOZd
4wVqJz3AvuKkP8V0qljcySKl/k2T7c+ZzyAsJs3XZ2J2Wk16OL7SfXcdH75qI+c1
509mxy/JFunGrNm4IHmqA7oviyN245i8w2i9XUXkjwprKPa7tH3eETNlJyWxFG6y
gItetDuc7GZ6MMLyZvQlFMjgYeAs+Z0+aVGzMEFWC5sOhn4H4d42X91eXcag59kT
bV+CCE/gEY9q+ueY2linI8CnrZXwPYc8FqRM5rZGlm3lrrlNOct/BXJ/F+S0svuS
/dcbLD/ivbCGjJJ1ZPYPK5NN1xk+G5TLz2UonfCtiEtpNGW/Y6UER5eUqsJEZHhj
Fugcc3B3zxoyErUkLG2LZCzk9dYul3ATsPsQar2BjWJtB3yV4pBb6mx5+YbBVCdf
QdYspXvuvB+t8Y41iZa7riZz/5sqdOH0h9jE9yQPPbd7rM/IF+Wb2SSwm8ucmOG4
74lyrnbBvt4U82JvxLtOG6RGkUG8haVrKN09Wuudxarpm4tEGu4OzsQdcb+8OKvJ
6D+jIiUc5pO0IQut6ZLTY/fw7WIgYDkEB4uvKB2SVlOpyO7dnpsecBR29WyJ/BxR
D9458//E8BGHj6cQ2bqMmBRCO1dxNjWq6LKl57LEXELW4dVU+JgPCGMidE26L7hS
8pMSPpJY8Z328/GiNdKjkNTGRZYYd4ZHJ2c5lTgMWX7QuYBP/1gnwNfViBCk7inU
sprS/oNSe9OVG4A+6wHhJ2c/coW+ZZE2PnE/w3s7iEwWdU+NqZ54M4gq/PkSGRlb
XY+08PoWn1aVTetXkM5UrQzVmpkXQ+pTilaq3IjvRfGtEJK49ZW7ye098MH1nE48
GQRof+XrGFeqsv0RDrP//xEN6wy0DhF4MfoSYtCtdyk59iJ4rR2YKxINdhtX75IU
yRNImqSZNCKk96LLhzl8xKsGnhCajzbaREZjmFGQKCmwvlpZS/4xi/XPQNbB0/bS
HdEOOemO4BocM9nFAcTXhY6Yk+b+dxT5HM658K6d6IsAGjbViyw+bpBsDc+J4b+w
K9m9bsyzWvJb84NUlhY/LHyfPVjydLVQIwxbmwiljRiUxdhFUaGihrnjeqUx8/ZB
x3r4x0nY8b3WKoDzimyJDcfKEPDJ7saN2BjZcnA/L9XmI2vk2OHQOpAu7HwyY1Fz
1ztsP/7zhexTKoy1tOxKIOA3ENEdAr6rPy7Pktm4cIal+eqksmTsUOjMWLVaUm6C
liC4Fd7y8J5fd/mH42X6lXFA5JqjY4mxn+a/RLDhn7DvqObq1nQih3BMfiruaO6u
3VVlmCWic+ugHuLYmSM1l0/wfPKwNiIEKnrnAgl+7IgM7eSbqFm66f/tyfYg+CoF
tf6dEyBj1TnAEevMqYIqtVmoFp0HDPYBiRnU45DAEu3O5vGHF7rLtz+vL609KIXc
+tUw95Im5q0kmX5rXBrbnAasaOdbwZ4jNKt5fxDACAczac8fddX5y/xhWUusk6jK
bTm/8J5nMNb8xpYy39ZBKiZq+SXhc6AFBo0wL4fmhpGBa60FX7UkYPYWg+OG37ah
jQg5nyzfquEqL1i5TilcKJ7W3fgGydFpSGfwEZVOJZKbdcC7YEnLlSnC71JD7Avw
STCJ73R1EFmz2Pl716ivDt/OikQQDQouIDZ2nDil1gU0MigSkwsan6YuE7sP0kCv
NCdQIg/TdQv53hDn6VJmfsRFVT+5QqSwy3KSplcurr1BWCAT7NBm6J/NOI4+OUw/
98oVd7fuSC9rDVxDgCkXuQ8jPSOnC5gJT45ncadK8lk3CHLwfyviLYOZjcRA+689
4Bg3Z3nCambkw+65SW6ZXXzq6z735caGnYczPvFgDWV2QCpXwKNijtkuJfjjejCK
OzeGJVEQuufrVXCa6YVat0ohuKN9MoDGEGX6TNyK+zyNP6HvvHpw+19jsZ6KnKFH
h82StQvv+2JWAAtTxg6AFZYv7uYjExEeRlXxaV7xAlGqIUgEq6+3enOn7vZyH22t
KD6w9+XGEGRW9aHkWxvgegXZHa+gcqJQ8vFhj/p7gFLdW+F3JlXYl3RvYEjvIbW7
T4QTrH1HN74TGf4IM2q2RFZ0y+vP9WQ8eiZg1QZw2hlMB0b8s+F1/83a7P11U83j
dJglmPBITpD5tVrvFaVC69p7qksngBCj+KVIeixv4waM9/hPaugD30t0whu7iqFz
9gg6x8oYHPm8H85leZVt41KrelolqYtcdtSxaLvSXAkDH30JbBowZ2kM+bnWxhAW
nMzUuPCi6k0XkyXJjY6kwzFgvzA4t8YcbTsmkQp5AGUM7waMnYqYxRVJgUhuvbHR
yQ8OathyJR+hJH3XOlXI4x6DwFrqF1JeGPyd2CdlKyJR2nN4yAE1Xr81Nlb2xDGR
/vGPtLcL3uBWQml7tHAvdV/FPyu1GpKEObjrPrfxRPUSfVsDC7WjR/18mq9eP6I1
OONxVjm/26Dn7O14SfduWtNDUrx0eeRiQXxjWjfL8vdPuf1aNzv8yVJ1rUTo+yJL
PvAJ++BKqPAsrG2+eNLvpvCpIUnNqn9enhQL3noMwYD27n1b7zHFObdko/mxSki1
nFg9Ut3QB5AdOWpozcDkEqYcv4SXEBnGa4xBdyvRWPKZqZur8kLu6VUpOXIXY9jb
6t2IsmND94LqbOnd1VZ6WS+Z77mCVzxnzyDkbah2j0AMm1EbpdC9H6C4slb9jrq2
n/Wza40Kqf4Rw8zkKYcew2Hck8azFpuHh56FerpNypVgU3VGtmY0OpY6GxL8imJ1
tXDjpzMP9iYu48uENVTn3LiKvEsbAtuvG+4h1ftaeXOo3jL4KrvIQg28De5NXwgV
++h2E3YU9j3FJosBXW9Zy/11RVD7RAtjR4rqaKXOyWMdoRgourQvNmMt+iDtSvWA
YrdbPBDRFXUVheaYilH0cOWLbgxqIhEu+tO+b4kWXNvc6JxdV4C9knfyj10XSCjo
sHqHkDutnkhV1oMgGmtL8Sg/S00llnphZx4yBhrj6cmyHRbq7hOjo3NRHMuepCVR
bi7dAIQDT4RloIWxpfs+jVZNKCW0f7lR5j0FPMSttkAfmYeSJslg5hkzsBLXafF/
woRDDwm/u8tBQ+01WXJLJ1nmTHHhIwCepFri7IjRn2+nsoRzHGL6KyGidUGdolSY
TpioQo41LXR8aLQCM9UQunkzl0Yf4t+fjSjhuzZvFcuteRDT7/10H5h+eF4hyxWL
JtmvsRYgp9kUtqyN55PM5TCVLrKZlUn9FKWpnxZnROnudGfb6nZpgUmMdgeklWCQ
mK1SaK1Kh6LwBnm7v/V+kQGJbvfFQ3W8AoR17JeKXwmdGJWINJEVHZpWk6vPWGqL
g2QaVul5a8T6Yzl6+VfctJjYh/3Iw4oESrKC8T91oGE0OuLzMplb5RbBUmPCyfyg
udYo+E+DVN3lzlSPPvK+GNtpIVY9dZHPk7pXYrfUBDkWxS3+O+FKC/SaP3yDKAm8
4hbaWkVlqxsCDzSj6oUO3/lFEaMhOak7qx34cw0c04D5qGn3/ijZe0eoFnTeQpdK
eVPuKV0OQ/vQ0uAtcbEEoQpKfGBAxiobrFNlApjmWLQ+LwoDf2flF5F/Tejne3NW
9v1ljhl5L4HW04KK0P/GYIwr2tDXlrr+z6+kddvB8vWWyLzDVC4SNqkTsU2uio2K
T13JIIJM3jSW25U5XjnZhTQ8LQLahdSWHZYrbKqH/QDSbPekdMmwzhLzUEDkbEQR
/F3Y7bomYPSPSqZGj2xs5OheFpWcyALDB8h0vBsiCJKl7shr7BT/p07W8zWwLAXZ
hKqBzN6A429EA7oSXB23+elDNDokDfYZ9sXSCquRKhvGUgL6lizMDIt+waTBoxBx
uJdYOsMwW7QCebojQxTo6hwCXiFY1Va5r43pJs0ZRUkBgldOW+GD3nMM8sNrNLIB
uJqQGkxpe/rOlzeOlNBo52KlUqjXZr7or8wfw3NeJxLhqCVDBqWRRfcZ4Y2C1EHZ
ft4RXkBnqU1gIS+nHqHqqKyJi0nB56hZC4sK89ChkD4FaqWn+N0a9v8FK2Z58Wdg
sAoQr7TQZG21s+Q0qz/Z/vYrc0zNhi+WW5x630N+/yfWQJ2Ov1xBDtd0ZieEvnv1
Lg2IVyom47QF5Z7TYCtkggdOJ21GZyWRmkFAfScI/+EJFq8O9dB0a3T/tMslgJV+
iNr9v0bFE2K31HXE0T5ihpCsHv13ZRn5uBLV9oKScAmCKjQyiWPa6g2FI0yCHMLJ
Yrx4X+LUNylRtn4EaaE+H7CjYvkRO678KIso65Jsx1OTGVA2TNwCI7dmMGhT1M/I
SB8eWs5A4vsO5dVa2KJ+BvRPwrI/OFNRJEDWqt2m3egrpLtBZkjd3nRxIXljYGW4
nasKfcBOYO6zaWJ5Cv5n/d5GNU2G16Z4TGbYB7r10pGWFqjYFr+aw/gaYZJi5zqy
Sxd+FncDi3HxPxRpqxWf6+UU7a9t9XCfHK1JDfysBqEAgSb5Qian27r+I0i2i10g
BgNuZMA3Sw30wpj8dTekZJLa1gCj+wfLpFfLujP2zkCGMtGa5vAijOLaKxozEnFS
fQ3CUfq9Tf3Zr3ANoGmwq8VxSlS5z+b/UwC8ZP2JSBTuzWV6ZUBoisp+d1912wGb
5kZkN+YYKI+NGhYXIs1I/rNoRyc0MZyaWuq8spE/czHY/RRBrZDVwx9kYI6Y2clq
FGtFXR7KyUqtt+/NKlZZENnYVJPGRso7uQZCKtLuquGB8RcRu9pzssl0Ugi8YIHH
MOjJtvlDi8UthsvP8KIswD2kboXt9l6vfG+RvNMqgY7xa4RLQOmvNsBhjVnmM81Z
1r/B9Fvcz1DqwMJjIBvOvR3sqx6+e/u+MW3PYai6NtisAioYOXYIQHCruvrWRoZM
NWRkWRykrWhmOTW4r5mvEsxuee92L2QwFtK2IE5gN9xzXr6I8U2K92QGgJZBCjbP
qEbOrvB+Y3Qw41/ntFd7nbYrUZSsAJ+CQRdJHrR/OlKpwn8iQmEIRL9XrgNR9X9H
hoEzycVqpiDVgBecC1/ui2TFE4V/Bt6WKaybViW70RAkVt/NPMG1wcCYLF7HlvUv
0082ft1/i/cDTEx2ilT2wFFrTUVoN8zQl6ujVVaMebJFjQddioZ/X223dhLztbkE
WD38WEhZUFRl8JIt0UXe73xKOWeml9asSaRu9uLQ6YWO8rInqLPTV9RkOPzZ2Dpk
iEB/rdr3o0brdSWLMiCn8mi2nd0yNzLlqjf3iYAADrnyXwGvBm+fPA1g53TVd6jw
L72TFb6CYmSJBRCFfCT11tV/RtZ5pUPRByM4tI6GfkxJ+yv3w5dWvCupB/N3QNdT
fZJx4TeGyz75Vkxf6hw9Pi9WI1+IaB8yJnUlHuZMC92oGEULvKK0ze41tLkt2ZRj
58IGGuXW/kfSvClN0mEuOrcxPaYTuatzITE5QkUJ/LHLgcW66sacNtJyAQFcCzG2
p1hOkbnB9wlPuvrFb37BH7BX+D9/DxBnIBAb8wrNn4pMHWgc1pnERtZKq0THMdGZ
t0ZXMGdg4qPTUCJbsRiITpimxdFUyB9XmJiX/yeeC+/jorwqOx+r6Fb+EmLtAzH/
/IEleye//lYDyD0YPdI1O4iKjBW+z/VPNSUoGvKHqIKmwT9omTQGlL1I2Ktg7b+K
mi/xX2zrXvVE+eU4g6ZIJff9pfbyFpeibXI9eGgYQYNVuzO9EWP4Vb4UKA/7eUb1
An/cbAru//xbR9HOpW/FyQtMLaLz5ad+D9W2s41kANpPLvyomo5G8WDKoNIhdmek
xSLwJuhtxY4GCVDFjalMgOldic7t0OB747GdM6Tj4to88Ee1qt4C1o9MDNYkV5E+
m0xyaize0O1hbGdAE8Bbuwc5Xwp5TNsgKYSERdjYxMTsJlB4ih4z2YKVHtLuxEvu
eoGMI4pRK1BDAh0VQ3BQp48uUuhvtuNXs3J6i2W3L3+gN51+YtvA+mWn2qBLv2UC
yZqRYtngeqLWDcov6L0G7oSd8P5f5LoKGIQL+6LNpfW2FI8K0iUMtQYp5Cv+JF35
29hHRdSrtrRaypawBEJiAZDNbZ6edRNsaqla8YwQeLSxJh5Td9qxX9ezn/l7hAzo
aeCZFB15Lstrq7lEQU3e7YfKNptVvmJ318sqHTbHMs4GxiwsKR4AOl/T2mFNsK7Y
mmsU+hFGyCnt7nKRh0/om2FIPTsjWd3qHiVfbJsTUAwGkdNxsDkAdKUa/3chAFLR
H/owHZu0drTUT2//AB3us21HKm+0zv52cRgoLl+exv2GsF4RITTSnWn4QWBzSiIR
wxUACfVd7vZsk7RhlmnUU3Q4JYL/T2WEKN0ERRPym3IxX0OOzddCYGgvvyN6M3ud
RbmBaXBKcvlSI+TkaAsgynm3BPDD+qj5JPr4P0ECJzzFmr53IrvkUEKq7s8Uvj2d
WzaQ1QzRnS+/xgFdC9wX0OqdoMXtqxSu1yj0acyiXeiiYl0nJosWZCMFNB66aA9c
+EteY25QzU2A6WMw3WhE/qGRRm10Lg0HxiHdjYN8h8MSsEmESJAFyOGZNnjjGRrh
x1guHtS0G2rkAWBvwzGCxg4lMLzllV6S7a5YfIvKN8STHh1oJKJK2kwljcFOuugR
hXIRvt5OWMN1NYpSnrXL5srl1il7dxO+zKd01uLcGoRjodXTFlLbm8EsmQSGClGQ
JdjvVadcXB9Gc2rsedAKkbm3+25YGoVBVz+hQjklsOoj5IRKCvtxKvNTQxzfP3vI
IVbOcvdZssIXe7m5+QurLovKDRxC5By8N0oIuhjG6m1g2dQt7ukmDM2S78sCFt/P
H6pzHgoMkgo/2eWHzvnf718XsDX4GJ8E2FUdEIJaTweDjscD5h5HQk6pmbuVm+WG
deqfGQSl2dbwKLUSlpl8Dfo5E90fJm6K4SARKhGWKmawo7Rdkm8neR09MtJbi1uE
bEab0yAiQGG29509UeXYv3FH25LkJvuje6VarIg/1/UaeANGc1SlNbZuaRggJnaM
VpFmBcnpRX91YPSCGcbJTN7IZxj76kt22axzoQYKe2nUeZkBdmM9l/lCZ0j9F1gf
CXtaFmF4Xi+8pdCHMkltOlReaLy9p2KV/E9zXAVRLXwvpwn/hQnOQrIsCmGoZCXj
yu4rdjqNWTckWw9OmufHCNZDZH3Zw0w0NsNgHKtj3Qi7z7bVeeKc6dvjmO6hIeSo
nWl5T6wUwYzJOnK4pQuwVcr5wtn7b73GD2yvZi259+zOG3oijuEFVVKGoTwPxMSp
aqbc8EGrbnIGi7AtTIvhHCcqZY6KVRacGhWq10PTBuU5KETLhFcjnSTUi99oXHwy
xfWJVNz5+mWsNoV24dJ0q255l5f8e+MhcNYSx4/k7AzE9fmJdS08XxJIPKxxJSZs
cAI/RU3MGIjoz1Mgrl58HV+GZHsvM2pUch5DUIVw1Ez/7E4tWJketisSYMm11zLJ
7Xb/48evg2y1efWg9MZ0RxWjFJJ303WUUu8JDP4c3/S8egomQNFnRQylxI6L4pX3
c2+6UoYyP7L6y/nPwZbTHyDPplzuPRYeU5EafKk+TR4HrU+tNLP4Fh3ce9Dq4eDx
3r61VUuZHQ8pQ/fyHoszruok3y8xy8XBxqJNTvfrmBGI4zFrwbAFmqFBzL6acxmz
1JOdx8dRFdhZpReq0148ipsn7sNURT6CEckIzWNOTSK1litcfUPjbU3jzd6N5NP4
umLJLeuP2Z5AiK5/r7IB+yflNPGlsLPCwqBMNGSo7B3ctdLqX+tDt8HjLLX558Gg
Et9wQ5xfM0kkQqclCHke03zvIJxn59e9V60yKRitxCxP7LMFGM7KVKiADD52ioX1
FwHYzYem4WqhHuEnTvkpHu8u8HkN1MbqovMiDFcTv5qdbAo0vq3KDlzKL06FeJxv
rLoFwmYCeIY63+G9EltW9cvLegS5UzkpyGr/Z11/eKrfsNyLm/oXFdZa2/qw3lBG
MbVhmmxW5tuXgrKoBPOPQ2PtxGGtDCpD7yJy+TNfTRkJSjjU2w2Uljpb10xGQVEl
O88e8Zz3OmX1qkM5qTsA/c0DBK9VVo3Tzt/vkIgCaTP8jp0NTgSCpbpO4uCfU4lx
CBU8b9ZkZQlhkAH9D14UQ/qt0CEqJAZ86hjvqO1wWfOhQgRrfyPK6jp3I7tPMgHq
mj+Rav6QEUpyWTNHBwt5jPfiH43Q90SdE0+F/LUfqwUy2zYLQ23+/PFIEIdOyz8N
dh/EHZpMnUBPBTs4NzIe4otx7aYFgaAQHj41beZd+TvI1oHXnJ8WU4hK8iSJJftZ
y4oxZA0OxS+TXmC2HeWIRDhlWcwBcL+4S3Jp+1GFcprZ/ew2nLxnXV4KRxzrkHRi
JsiEr/wO5jb6K4R5WTVeR7elBlUPG0CQk0GKjDNzGCC7fldkrHVANb+aLDKTV6yb
k0NSjx982FvfYufCb6uq2U9AAyYlwd93fsoF9bNGDjBdaE0FEl8mJsILS7YFcQ7Q
Ki5jOb/p7HwvG0jE/I8EHam86fDwNwklcPfmVdGZIsh9DqOzqbNqqQJZspvZ+LiE
ZCNr3xmYBuGtymuG1b2b9trDQibzkpbPEekybcN34shQB5228d4hjGhhkSL6b9R6
lpdnNr5wy7YqB6hK4Kzf4ensfgaaaDUw5BcNT8SdVOIzWWYtSDgGXd4o8EE6pzWG
Cueau6lna10Z1kB5wg5Yo5Ha7juxmQbqdqKXh1kiH9pvclRp8gfP7C7tARA/Clkx
YY1hTNfOex4Q/MaGaRLBr/TkZE/hsTL6isPY0XO0v8BqngBHrxikuAY1YOAU7lMd
TGMa7DEq8uCx1mQm4ncL7LC8nvbB02ZQRvgXX2+cb6rsolh4pSMYmCG/57V+2cye
B5mAuRgaZpVAScN4T36GpRhIsFMh1/Jc+6TN9Ewe//mZerUZ+lCeCJrLp4kHRA5y
/nwXD+1rm7yiN9eNOXgk2mi3mpCK9Ou/Vayz5OC68c+TaUmtqIxjVl6S4OQFyC91
/ATNhff3ot7D3FeKGJBJ2EXPMSiBdZGdsSe9xDs1z5B9h1MkeDWElwxW1+hBsHhk
adci9vA71kurA3I+Sq2qNnWgLsXmgvqAEz5XvinmHRwdxJD2uN7RLvOTTeffzcI0
9XtcHsbPFiq2Q/u5BLZ6LqIN9TVRUtHnTH3H+vXdIvyJSJbqt1hwOZzwRPTIDkQZ
V8igZx278EmOs2DpayrFnN9mpKsASnSi/y5aq5BFZoaF0porFJDosytIqmhzDhRF
njFrkWyUw3tkYpmBMKqZCYbVfnpfrrb0D39EM5LiCr1BQylRH77g2+ue5c6wu+J4
3Lm6Thy9M1uba8/OC0nKy36Nd1CHmRTUYLbMfQgH5+mGjxH7fPVdxZvo2OuGwOom
v80bpLTVhde+xtSCfAumcpxfysoSkeoJE/YPXUtq5THjWZR57336MddjaNwBHBqD
paUml3spalHZ2JhOviCXDt1bRFADjPiPeDRbMtQ3WBYa9FZ4fyFNEnUeJlPWKLv8
5BS5bBiPKNYpd4UOeESndeLd6lai5nU6Nikx2KunA0u8/2V4nbykYPbA6B1zEE95
/m33uMWT5k5rOHUHtX0yBfInz8hWMQhEtMGe9+tka9ijlNkHXSgnCzVEw4H6AzMy
IR5Z1rXo/p5DUCuq/30Kyscgpuk1vkQOp/XqJXS7cAppXMiT0FaPL4iDeM9iNBxd
JNZzMg+YioHE9Gf8xAlV/L2+emUiInJR8Ayf4uOOn+EVOagvm3ZmC3ZiU4CSkshz
V9pOwZ5WYaUrcMzK3Zetcjq8koHKyzB6T/xPOBTuOCQr45hTd8cyqbf9ZlTWCJOx
jvgWRp5BLlRBkSh/bngiQ+p5MXnlr7/yR2vcBWE9mvvVjwLKkdmI5o7b1pXAlh5H
Em+nnSKx8XUTPYN13aPagvLWZQ5s/ytcr/OnlL1dOtN6UuiWVagPAgCOqZ+sePYY
TaZa0jnQVcSFWeFA+Hy6WUtztJT7t7gYM8lY3IUg9UnVRRO2KEZXr1uNut9uRlXr
Al5IWKz4sCWkmc8DrB0fiQfKZBd7ffNBjhmEGjka3A7tW2k23ZAQ5C1qJXgCNIRC
vOcN0OZ4yEzIEX+TzRqADJLwambWQlTM80PPhOz/Wz2cIIf+M7SoYGTY6tFX5SiR
EgLbZYrHwkZ4F7jaysZAwlvXFqzAAt2EUptIU6bHd0itJ0fj0zl9Ifn5a1LivJPc
29JuDr5/11AgM04C9EqeuWvVWrX3n63SSOIYI3rARek3eQOvcUPBrcs6cwnAWKwM
+5nUFzt6jIQwILIvpy/CPXDLjISNGAb+koQHl2gLU5VWaww5ErbwgjKFfVd10Ppn
ka4L+eL4lLXdZfMoBv7UdxoFAxNdNMvx0ccNfiYS/0Fsgr4jLUDzXyaxlKRw4Vpx
6FtorJ+DnbAoom77cHtwvIs9zPe5TkB1FXd0wrz3fIkf2ALluqMzM/n8amPds+Vx
tzsJTCeNUsAIkfHoJD9HlphvIwSyYhlkH6WeFiUHXbF2LpMBQBsksCrmSVWM7yYx
Pe/xgyIED905s8sTSLF91IiAh0WS88sBwXvG4aFfFGfVNMVQprV2VcrLraty96M4
L6E2jL6bsdHegKUc9QHhvLweooxJ5ZHNf9hQyCoNMHWBQj41d+Yi2/wF7hdaH3cD
6HBovuP7PcYWjAAm9IZME5ypzcpuA1GxSx9r09R9X0yo8+9EnWx3uMlrugnjMCDV
YG35qMzGMUyADjwbYsACnqESjGHY5gorGvwhIIWzwQsTWVW2eW+v9q4CJOnwV6Uv
zvVY6gM+K/Q07Fsz4BKTaqOcOI/XXDcSXJoEHeysDCW7KNQnYxCj3jyN/uaRBecI
ePsj6WbvGg0Y0N5SU0AX/CF7YEvSSz1lcYe3fZfaELe/OHSFaPlFtvWXqerux9fy
2HEoXVYG3aZc82EBIEddsx/ny+mQS4NXyg1melYNruC01MnkoHJvCfoFxAF2HERy
Q6ju8Z8uYkvgkegH2d1qymulAReeRZv7IcHodUMhtml4Vv4D+XKver6P2Co2LD6j
Eu3I+We0xI7ONpyTiYLJhjQndvQ+prW/tfeg/CWkXCpFXsyWHZTjrYvfJ4QcnCur
WA59CWrxVkijIsS23CaISXogAYHI8SyOlZE37dRaVwjGBBAZfgtv/gXgEoMQLbkZ
nm785uZL0Hl5siJcWg1RavGHMEB2h/OsU2ad1UWrIrl0znSww0iINJwXG4kOeFXG
DOfZru90CmjEpok1N1+V+zRmtfkFhyOsP/lfNnHZcjkfGY1vX+wfe4JaS71Q2ON6
fXUiq3Y18jsAtRzyYaxzjM/AtzwcjvJINnz3qsP/QFJSQuq6kyImT4gwz5MgpskN
OtuHCaGJdPidVUG+ayGQJQWIVfiKB6uP0Tyud2SWyMmz2iOkUXlZa/GoMVflV1uQ
S44DKIMFmSztEjAz0BK3GzOl1Xx5voRX0/7aYGKKYDHqju5xQmxCNGodmSOGEav7
6IhLsgPRNbDoMWgVJ5ZQVqVKuWBRecTPbP3Vr0NFDaIvfDQGWvaatIxGOFojRNhd
FJZxsh4WXKAT3gmQb29b6YK7n1ZwZc7pP4eE+4cvBioVjbRuGHfOt6LaO33O8h0e
Iucu5/jpSiZdR9WBGnrV+O+R2tdT3JpIhWMwjg5a2HImA9KMTJuUx4y/QByLOYH+
17OWG5bIUbc7cDO/PVwvBf+H5TIqAU9GzQ1dH69MgjU63zYCD0Tfe6knJv+ywGI+
joqDa0LRBPVTuSxPpl7uPNZqt6yQ4DVndXuUASzXC/qV9gquy2i2SjCA52OOO+U/
ajYLUSqFgSQeaNaqfyUoZOVFI23g5OrNfm+898/UYMhyY1iJ2YyRgp4fbvv1KhgG
bukr5hNbonHkNNcksULuKQcKwMZhXyRkU4SdIGkuGsA+JwjdPBtKB8blYcKdtfgn
zLcIvNxwcFF12jWEWb34epkVvEUljqsFEJsUIc5TjkfVyten3SOch0f82tirObEi
OEC1/u+mv1BTD7gfdyBZN0lrPGQ9GbOPsT2JjTtUBeamTmR+5Iow3RruBMDe55OI
oSGvYaNoIdLnfZXd+TDHS8Xc/TpTgb7631whWw2V9sMVebekKEAuF4JHOHz2UBOR
y3ITgH9piOqhDk3SzAoidR7YbgdBEnxOjEFg1X7mQgUjADJNC558iQChqPe5cho1
4JAV5SlKY/M5NSvfZfWilxGYAWyF8Q3/u51TVZ9bscSSSEU4ZJWnPGqBkehVYHIG
Pa0nKf4hSAHBNwBP4NDi97QkRebgYtFVBuUgiQ17n29WHnwSbXz6TsvlNpccAVal
N9pekDu37anwWqPXDoNkOIzZHFPvtS3Y2nlosTstRaEpyqgy9qFE+Zret1KA0Dju
E/nkVqH62x6KwJnds4bQ0cz0qwEhP9vjW98DXvimWky88puMBx8+7Qr6yYwYLqdc
VESkRgF0mh+Mn6LdoNhZh8IEirodR24L3atP3HKANN0wDi4wXpwcAJA0V4c8Boyk
v4Qwye4GSbxV3SeEP3cOYrgnoW8VkiSOgMWkrMvCD9DzpuLOgQ7bu2W1zgekPRSj
flDQHg5ATTbPOsjifGnsUIzUnl0bmXB2m9N/WgBaRpoeL0rQw+u5G9Z8CGdeWx9u
DaqeUmSmcGW3dL+tqgKEkzPooGPPJhGqAv7izWLQskBAUcB8rkIPYTPPWLQK4RKr
Bw9s0xla8AwuG7LnZ4lVl3DNlzsbC04pj0fNGbysqQRoL4Xnr/1rKKgL0/j4Q16N
5jiarrgoecFn4iE52srSFNgPuzWC5nYSkJbj49415J54tbCXFPCXLDNS6fnGlWjQ
sezRnjhLC+TmQsE++kDGIwce/O7UVJ5pmLdfsDxGn7jNjg9kxguSuXMB6WdVA6Gh
/QnlcJ/c/0iktZQQhxynL68ir4h9HzDBmXV3X0ijmcocsgsoYsHxkWwiSZA0+3Mk
nOQ8kAG6BjxdhJPll/q3j1LVZTqfO9foi5vBozRRRVUeggWZhJbCXbRNApu3/Op2
aczx2NnfE671kfoB97fK/UNT93Ul94CTgC70aOyVMVjMZfRgDxYOYkvxbb+lSrM2
wGyPiunGhpDSQZwlFfFT7814WRY/+1KPvDg9C/0tggp79Ok8Cfp1EtGpOmn3J/nl
uHTT+9POKOkR5qcGP3pQmO47RcUSD6NFPhOmDj3O8gmubnDtUG21GcsaHqcJwSFY
DU1/0gVWt+XKXc84WDXb7cv1AzHWqsuD8m8gWot0gDZ0USfb1zNqDCczSf4mAJ+5
/sNRhevXseZ2w5i7Rpt0KyU5yeKSdSniF5/In0a/VxQ3ieRNzs25LQXKlL0xthyJ
GTk5zc0rxa3P7gC99RZsCdmhhcto0dKvRVu82UmAAMSEg2POKm5dgjU0oh2Yhsje
GEwylUuchdUkUcaePxupLi7fv4j6iMsWf81k6tphE6xUZDogXic4ms5yy4uGBh70
wRgZhSZ2l4YpW9Bc0fO/Tri+oi+bF2JL1JMDJRVDujFcm0DYs1j5jN9DdlZ5px22
hNjPrYzt8DHLxbqNMYr2SswrqIBo/sDFfCbLKwMFg5hqLf0FtL2He7iFOYujtJhR
FzegI+cQi9xMRifNNJZg1TSy3QYmDwwv7i8HkXNAu3EdviAumC5zvrPQr0k0lRAv
Enk1hifC2eCVZ7IyZ+vEydujiyOcZfg9mDfqvsnKrJMio9yCiJY3f99+rSXfFTXi
JnF6sb3idG19Ax6bwlY7mlEvrMClKE6gozOZvTPPmgsYRPrA6NFl5opoD5BZlsct
H5ubEcmPsdJ9Qd/reXiN/k7wpuPGaTDZS3biS1+zhyB2RRZzlCU3Y/tZ//k16piB
knx+ZZ7TyRpajsIuDml8DCY/HqA9zyJ/PyYoyS5fcRafLuBslMpeor7tQmeBk1n1
2479zAXjqOeHddD4D8ADtz7BTn54hIDdgpujxnE7rKCHaQ0k6ezikZ/CsOabGUCO
RUnYU5FKmqCC9+u3a0VruepoWpMp2qH1XmvkZDLrEjnasWNrik02rKIiTO6YnCmu
q6u8Yazso8gm3RO5AP23cdAF1kMu0K+So3JIpBzixdjFZuTtrOFQeLFntbyiTtsL
0q1DZeObesulhFYiVfzhfL8ZvFlU30ZSUZDXIJXrBiyRtZoqffetKrfIvDfeWmeo
0d9cM+k4dC7Ei59zoFDCcmwIe0XqIkpkxV48ceAXUrnqxiS5loRoVNnYRAwNYxvU
F9XcYzv9ckf0kk7nXp30AmfvN/ETm3DsZjROOoWA4bm+XDRMiAACXIcduRp+xQ4j
Gci4K88eiDAPr9VtxX7Kmgoc7zIi1JLlZXOAzm0gXT+Iibi+cSt4ibshujbRGK3q
RqGZVc29gTgT2l0i1cskR8cVWE9xQNbCFO4ByE9Sb/OQ8Q8xxs3BhPFqZnMa6jZZ
QidrcsnK8a8Tb/vQe8oG6HxqTANcZgz0N1TJUyKan4OyolkTscG8RJcEJ1EA+IA9
pWM4OBY/uGxzYDYrEqaKdUpl980q9/mIoXXCigr7TwBovZHjJrgCY4xFUOng7h6g
nTYFZJOhVpW75uNZRbacJO1s1z93LtmYjB+h2pLJxvzQQfeJu43PvJcUNkXwQ/ul
gOLTrIPWKafav5xmF8OfSaRB6aNfTpJM4W3X1Q2NgwpwnZH0D3tUcWiiHf26OiBR
TXL7/PtV5BTykZJA/V8rjES4wY9V6101t7Jf16tnZallzVuZtQFtqWkn2pBu9NxZ
ETEBdW0B9IhAAB2EJfvk90XxPOT/Vu5r+jukQu0X7jySoEJaD3w38TRq+W8QnW1r
tXi6MNhdrf2q0jkG2eIbPYmoYhtIED4DVlQYybNStOVq+Jmk7s/QqtObe8r4iaza
r6m+ILbqj0dYGqEhQhuq5HC9u5WRwdpn/sEoExPEFgAxAlKzTqvZsu+kLMrsZO08
uQmdZ6I+Q11UbVegm5HaRR29ZsVwHfpPKHZLyTufTYcZM8o67KcPeyGjWN84kuLu
fFUMFkj3cKu7CoINlotKz/2NF3eGdKdaHFgmNcHM3w8AseDsE63W4QXMzT6SPVLo
8YlLpEnDqLN70NsXsX3Gr1YZwCgKY9YUeE2fHK3sS3oms2+BhPUSoidqc5vS2vwQ
wj08XtCy8KngrgWl+EUzr27fCHGXDxvWkwYH9b450UgSDxgycH0FQFyKTf9YJJrt
vn9yakaCGM8Rnj9xSytlpkECRi81nG4lA/xseCo8HtjHG9E9opPSjyrGlTgSiQt3
GmNTiw88kEXc11CIEpgVS0YaUeu9b1tfBhBZeNBGGhqOZCh2arpbdiKH5Hf8zyqd
0PJBpb3DLquj6PBcbJYa6wv+1nScfAOlv7SjzByKKxZeS6XfkN2sQcwXcnbqsOwk
5abpWdmdQrldvMeggL1J1AqE/y0MZ3OR79yne9d19v82sULEqKXiABwKnuq6qAb/
dENasfiJt3orHYLr+xA7qudF9MgXoNh0TKK4W816Vhe0YJy9+X+ZNSqXtxnwHlv3
cRlgQEk4p6dpwjyUfENt1XzMzJjKZCr7Nh7d+AJyYf6bhHEQRI4GTxCpgaQnEstO
kUS/4z1+o2qV9e6eWicWw7IOsGp+KA5EnNty6Pzu6conkNTsJXMoDsfQrf45Qx3o
NZl81pzMoTMwSwajXmE0qOoVRUMl3r/6GBLErZM6KI6NXcANet9wvdKg1p4nLMRq
meh4ovoioJ+f4asUA9tu5D/YurVF5JL/5mOkgn74NaQzHMcT7fxp7U8u//KL6lgC
Is5Md43nDIed3oWVP3/l6Rg35jCynUo9UlamSzuQLjP5MAYHQlqVlYrVh8UTou85
M0JsdC9xU3gN4ya++uc8tESIS+4jm7LnD1RJN8kzjExVI6Dj7Y7kwFPtYzXZtgCf
AMxZE8SBsChYOXwxif2vXS3pYQtk4CERSTtZLbUKIP2LY69vEUJzDrcDRCNOXY+x
6sNxXIfdaRawrGqGExSTwPYAFIs2V4aQd3t3Sjo72uOz9XuP72I/FbNF41IlvUdS
EuEcoMZWT3CRuwYeHECPVENsgeo8rYRhwk+4ZuEr/Ez6txcaeWiCiJGdMFQVboZK
oUuDq16D2ZfvisDZPaV0rJEzWmSoiY2Lw7QmBugT9rLdStFlVB+2Vl+7gFsvZwj7
3oV3dtQPZl5quJXJwhZ0YaY/pyeJCSCYC624tnpou7N0An61SUzlKk4/NZd8VXN+
f0FYi6KUxu9FznqPNcmiq0UqQqy900RNDuFr7RgUwwunBdX3NWjxnSCPgUByhGEx
qilXx7oP1dwgskxHT91owSHltAEG+RoP52nH/LeFAueK+H+CFAubaeWuK3sRpDv6
pwEHmZ1fRpDMOCS+qm4EGTXs2w/pSU3DnNwj9mhGKE/hpzspqeu5i4meUTsIpAwl
k41mojoZtqQE/aLkPA9oyX34KuNuRGaNy+5K7E55cIr706+g+kCFEgUA+ynGIOb5
w9kdGxVeVnIPxef2OfuJmyB4HqjgVGiaIssQPuKuO7UjPi7QDCSfYDpbD6bfM8i5
zSMaPWS5Az2jaKdAsqbmIcLDa92hVWWrPNs5Mzn60oTdazIstfvwCtKuFGdYYXRH
am7/zb8uDGSFRllGJU7SAozjQvkMzqyUfsxr+A/TuGEJQZVQWkW05RxG+Y8ruFKg
Zf68Iuxl0HSRM9jWn17FdSZxSBPvQSW/XZ4m1DmjERr2QbgC9YnPaUf2+QbB7soe
TyBGtLIGQlloU+dYtvqXiSLPMGW/AE0L+vP8TK3Ytq5zHL7HQNHxcGNHKOm7HYcY
XJsdtZbYu/JiQabKWgFtk3jkeJOUGSZ2pMcLjZtOuW3QF7KqzM/2gLj8m9ORAjto
MT9VTKTkIpbMzOHmsr2BVCV70JK5et0+pizo/rSl40vavYYlX+A5klSOz3H+WVKn
t5hsM6ZeEZGci+VZrAvscBexr4hb67ZRqhgVDqpOyxozOUd8QpE7LiiYqZGVSgWm
OxOfdvQMhYs82iSNUeqoIM4pYy7KkWK/vkLoW24gwDwf4GF2UpCZV+zdspaMY4nr
UF/SuAAh8PXKhZn9ezLYl2JkEGETVCo9JjffOEmdWrhczkon+UVVhlq1OeEfsoQ0
qRr/KXyaZDIqvML8vR6mFfyAvIr/V+iXQJCg17829gmgyIAoh2jh5BDV6TN/fgml
PAulFV+vbGt3uqUm7WWr4uAyQGq74MFrff4iV/XafCQSCPbi9+9q4jrqbnpjmNub
sE9xXA/QUSIYJAWIpOLHzry45CcdK8xGuQRdEEhbDkhuH2d0Yb6g59iyOabddBK+
dXF3QRKiiK26Miwm1fRedINs+fRnOhtYZWm4TOqAdBoeiK1P1V9ponIhXrcMpvkP
Qo8uzJfFFDNBwZx4N+XX8YBD+SVR0xN3Owrvd6ujbRB7sE3l5MofT2uEl05iF1JI
FpuqttAoQPbsgsJNOEUgvb2qKs1mrYQACdQ1O70a6P9tsMR2JcvUlKNaDD1A1Ynf
X/z5hsvGxCd4tob8wIPrMEKzpyiI98ox5gXyUD1+XWxbNqh4PpTXTrh+CLLQmxo9
GVUydoLGRzvzk4EBpnGn5AxivXa38Oggf2JgXg6vKRC+lQClQiuDkhfxno8OQHbO
HwdS/dyhZJALl4WgWaZKr3ej98EKr1z7X2ESzuw9s6S1hEDJGzlEQIhUNFADdbRs
6SH2p9lqjC57QcTAEwMuH2ev1lXMcS9a9feXmLqxgKTFHkzliHqtYxhyCPDlubO2
dUc5vyz4ET6fiZuDaCuwynlr88eBehUmWYmyzqV+B3qFKIvgV6wvdV9EWVQvzWwJ
daL8aR9vQiK8SbxhOo1mMR92nvpd0xkQAQMrMdppTVLi1N3WlgOtliPwHFv3tU87
ZLhHaWREezHj0IHDkDUJNmY4tKDkgc8emYIZq2d7vsYpgyhJbbsF/OVOdva29eie
ZclBFG3UsQxNtK9TOfuAbHrPodJc2kglZZzRsa57Wp92FmEKCi6YMvZ7NOVFRYFt
lOC4f3mhyefUyEuPr/DKq5i5JsBTzngn94b7Uo8Nudd3GK6mB1ZEn5STl3kJClRa
c9Y1V3YB/yVVRJFBrJpq7JFLtMDk1FebMK7KU8fTZGeU/dIWvvSzdunSTttY5bOW
O9jfwZ5XWPuDgHeFvSu/9vjrlA9Mv8C7CNf/GUXGg+rAdSfE3umFL4868WzMXeyP
soG++nxZngD1fgYTAh2CageSPV9NQsh1pAyNax+wZuFce3yDU6rVRNR2E/zoSFhd
Z7RmXIz7WzpfrI8TaaQ7uBdRpL09U1CAsSTCcBetWZIpUAzZdSCxQN6xFbJIWGF8
anfYapvIgied0+R0+zx1asiBOswMjThIzuBAYmnY/IhF3pyjyXz8OgQ6+2oJb1+R
BXZRgWMm/02ctpytjf2qN3BpJHxVJIkcjv5FAnkw5KiBmSvHNgTaai2mCR98aNyv
FXyedMiQf+hDsYqZLYerT4yu+NyA1SR5OpYwK24ybGZo5s6r1Ua4kEGcKmMJPN5u
92Jr+ZqLhXNTN13/ptSDCl6lHvrMPfi4qQNR0oez/RtCm55ukLGRZ3j3fvuiTWzb
tHn7qzmYVU2rTH4vGqeqn8OScB6WxDWm7TQOf1+jlzRW6X5RuWjNcUrSa4WoxdBK
I8E7VLAScN/ZvZMaTcWpFo/K4pspa2nNobzRbHWVO2igyDAI87V2VIwaXf9vZW2R
I2y13L6qu+0XerR+kZxqXwn6e5AK0r8WiuMZiXFwGpDrKYnJcOZyGwVtXVHRWbDr
yNpHBQi16lxrp1Ih4PvRPZJZJ3xlch/GHL5gv38cEsf1NimqjBkR6EqXfi4NhQOf
ZwvwpYIjmyOSHQi558lN54UiXJm0TXJEV5gGbXDafgYCcz3Wq7QxcUvX//X/5ftk
+1e4G4IIar17Ir9xdMAu7zRjBWeP/DiNfj2DlrnV/E117TwWR6hnXbvqwfHLQmv3
XBm9s7vmnKwm0D5BijAqzu0jRu6swmA1OTlBm1QKNa2KjHeH3joERhdNRCK83G9r
xybwcPtm4SBTQo6bnPqqgoicPWV8Gc3rsVf5CfNj99Dpfgi2YiJjmpL+vYDxnimm
cm9thdLq4DeLlMhmlNy7Nn9KnXyUVuCRMPeg0bCI5vkuriy7cLBpgg1Y2VBA/MYx
TA7iPNJAp0Fi7ZaFd4NpHM8i7MOo2lwv4Vval41n5zLlKUDJW+SJr+C/sXwX/R+D
8Q2jpdbo2JE40fca2J4DDJSkO+dX+IZDepeFR96BhNxHnY8JCnH+gF/YTuHPuS8l
CfoXUlZLooUZueTGuuf74EsGTdkfROA40hVmpNd0OsUc7OSe82C3dcoYNv8oYrTF
n/BJ/1bfRSDTo9oed3CfGUXHsTctt+AwWq63uojRAt3MARUrBi5ebD9TXzKp5iNQ
6OlXEtURsIOJdtKkaRttHJWRfhzGZbLuQSYOygjmPC4X926Hwx0Dca3v5BttrEiO
WmbRVh1ETMlyEmemmsV5vz9TDCTRTW6NFSqU93ITq/ZSHNduq+zvjAMebT/Bak8u
IDfW0B6IfVFgqhMjEdK+tr7v7sjqRQ0LjWpwylPqNq+sS6/03kFKE3Aesl0vHF7R
yVM5UmEJ+AqRZkETMyrD1byQqbMD1SjcdLdPSxIcU7CqY6Fz//dwHg8kaR7ZB8eO
LlV5S+JOxuSxxUDOy92P7uZ6VtRk7iQBqPEocXW38YeiyPwNIgyUYPiJWrvPY/vP
quu/W49RBkACDdT3S0co5cWBPMBHySf+4vD3xjerjGq7rFzqRsIdpTiSvpG5mp43
Ju8XVzi37LC+XPeID7UNFOZnZEJWNdr2ZCGzehx6EVchzKDPwEWPV5Euai7jOGhD
h2U2TfLrwaD0/qS/kz5m8pu1SO9HOIJ0QAfpHmqsxFpsDbRTOzLscfKzJaJfEDOb
3nWA7vcdHZKDlNmYXlW1u1/uk6L0k5/rdUlHAEIGro9hyEpElQVTzKccxvyVZSm7
4Eu1vOPqAv2y3XpJN2OZhQQ2/qGRyXRxOka2B5RMKg/PK6GOWykXVRPqh4rowkwp
+sez3+HLATaOctLCJjmrOJTKWC0lIw1a9TvpY3WJAgizIXdFX2HTZ1J40p9NPdtk
fjnkbcvJm/6WMqXTP8CCcnAe7NZBtv3ePQnDCze2Gj8sQ3lOgOmRYF/XBQHQy420
QK0QA5/t0F4h1L44RCG92MtrfWcOBuhEcTtYG+wUw7J5v3TlAPxYeHFySkxIzDNk
5u2TrzLM3sQ4o5ZhZAoP51nH9zkSJ7iBgLbxT+VN8Skmr8SN0803yzVsEAfXyDHH
qzDTsgsNkTj5rAPVJTH58yQQAKX3dmnQzhjg9ESa89is9Rb2UAvPDu7grnM+f/Ir
5LjFpUR8KratTZcaRV6A40gDFVi25qNSS9WJJdp3Ybj0orgKOYoFKD3AmSdP4ae0
KpJ2LuEsFdnLzKEX9I7oTGxl/gadBdZ8OOhyQPiw1vZFeR9+i+ngdyG+l0nEC8QK
Z3nUjhTwWlpNKhjtAonSjT6AsV6Iq0Rx3dicb+hR8YLzyB0aub+6qgujlukNQEN2
v81ds8ehF0JfmF+NTrQ0q8M01OSH/rORP2r7Q1tjwqZDORmf+yKP0nNKCEJsbGh1
BVyDlH0CNFOXA2t+/xxq87C+Jss7N0bghm3a+7zRacxIRRQctG9yuj+gL3XUbmxv
TyPWioj8kNiip3e4IQW3V+mqjC0Krj1CLLRUBqkrDZ8joeXcFed8GFbVVmREbpcU
y+RXYuxR+ZzOIeMUX+cwpMkpbH7csTfzuwvqi41bODVbqOZJ4fDuptaJ+n95RRXz
2cn/cRU7UTehEe2kgupGKrWXJMAKVuGk7a25F3UMuNopPUphAEmDpR9okXGSDmgL
jn/Yptbm/XLR2/aQus2Pt9Jp7PIB+ZZ74OuYBse+fLjlTd2I1hv2m+XlR/Emv5aA
XizVjRWQuRC/d6dimG41GFi1CLgpLzKBwUqbbjKuJkX90IQrJ5LiqGgiEFDvNFTy
SDYrUVER18SBkfkP6qw8l6jHBrMYP+JZq+Abfvb7OpvDMwqGEC4dHyAu+TfqYTeY
TSWfTqlCllU7kLbH0EGEUPc9O8vSxz4WkG5fKX1xpxbjFJVzhS/cRhxxy36UI4id
XRIro3+Kq7JnurtJs3+WRsVJSVj2s5BRRp2ijGn1WDxveimWuKdpxfkko5HkO3GU
UQkV/7b+VT3dVR+SdT54baah0TKiux9Dz2/iI1/cI8PfTtwnWH4xJC0SAQorSPuZ
psjPw8HJ7IlhBsyfktbGB7T6q5VDZ4I0w1fP2YFqERQlXuDu2uZOtCtHmumhQRaj
PTzWARLnx38+6NX2QQ3tBD9vKNWqycySLQtlNkDa4qTx5MvhZEYLfpqHvzVPGQME
+S4WppNwVj7Fl1hHwKsKI/j/xkU2SNDiJokCDshVQtEz/sU5iN0xYDziTzKbG0Ei
F6cmKYMfMBk50KR8jhOMc8Wg1Lu+BX5AvaAWMdK6ouT1z709RxdqzSb8HKhqO7bX
W3nnVMhVXyRfjEchnJTagoPqy16s8/FKRAtpAGb+xGnAoQywqwRied2wm/XZScFy
k+Y+CXBWfZk6hJgJCIl5Pd0H8gRvZWeCY2lC4YVAI3s2XYratgL6Tmvf9KbrjKyo
2OU6ybMp+VfWvGeSnArj90+uEnitih7FKSr8tUudoq+PwbPBeHgF4DUD5oeCBLjR
yV35LlWrB93p4YbPnmzO0eixUukX3Z1tVtL6NkhyUqdQjyvvgBGs3R3IdVV9ThUR
OQK7HI1YtiGzSzQPsmkEgxwn1lBMnUA9XxGiR7YQ6y8GgI/v5+lIRTLAAYe8bGvB
LDBCzXe2Vm0uI7P8EGqL24XYcX8coVmmulbaLKOEKb44dpD9OXIQxPO7YcVU3uUc
7FFIwwnNdkNUcYDnhHfBJPUTVjhyoEUEUZeglGr+YWXhMmco1wEWdwWe1aWlPuQl
0JcgJ5zNtJR4ANaBI6bF3CrcYkA+sFoU3zsXJ0hvutFEc65uCXPzbyzm+qzg/35e
wvxlevPh1L27tODCxrKd4496DmpJTb4Bmfev3YlP8UkN6hCC+26xESys1UMWzeZU
JJlX8AYjXEWVMAOrBWYmThza3Rlgv8WadHLsjlzD0wInb+1Z+/enVIEFbIUbps2O
EPfUdPnhbL0Wqyyd71VloWhJwrhVaYRwENVIBu2kXv6veTgZu0gZa5aHllKs8rM4
wbi9KHOlyaro3fJSG7s+gYDV9oR6Cpaq1Y33lGvD1xELcs36GEmcEsWq0+54YUr4
Kvkw3fQjulu2Vi3DtSlFda2jm0Ehnu+nB3F/sjiNVSsiIKXGvpXG+5niKoPVwWls
4hnnelxgtWWZ80IKud1j33y76Q/Vk/8CWXeKJizQya632UBeE2m8PSyAezQyXtx0
hO+IJJ7bLKJCUROIUCh+v9omIvKpSqSHVnDZpP8LITu6ectWGbgdIbNHy3wFHjRp
CVVN7dwdBXysDsqFm3cFZyQGxWyc7IALNcEsBV7nacfsivQzV18SB2YefrB0krb3
KNmmKdiaiM3nem3bssHFPWaLi4EhtHmKlQ2W4QW/rNffXtNVXOOveQGJdxYdIuMI
znCHbu3/mq5Ls/5xbUJ1GBWGhMOeP8fetaQyC5WRTkE8M/kR574l6ntqMV/5JoWf
DihgWa7apfl1NgAGRwskH5FwElvp1B32ukAZEUDh54eGKUj/6Yxs2w+cuobdQ+TO
/YSP1+TzpE2iwg76F4Ys5i8K9G3/l5aMfgGHmr/n/QhkRc7ZU9LC2bH81BpDJiAY
UQhzWfuNLWCR0Pck0+krk5l6PEfi2WX/4O2PE874dIBCzeBROVceRhzqktbxOQNq
LQl18QAQmL2c62+0Hpb6b3WQzxA+TX5taQtztS0vFd5aLq48SkYV/mTd9XvFMlyU
vzEqJIC6c0/w7BaTmyGoC83JjCqdbnScncti+fjeEfJ22wHWqlSyyr0cShy35Nnb
pO3C1lsOH/fzRmapOB9NZsrcU99AJGqNl+/dy2j3nR4Snfc2M3gNYkQujTKK+pWH
DjIqGOkzd9BwR9roF+sxXoC1V5bJCx1OCpv8iSe6f5znzNdhVmrlSZ/g7REji9aF
JgSUmzmayUOLr6qK2L3mb2zoCcXfPPtRb5N+FbcNvzK0NgMfOSk3oz1+SQOUrgtY
tgFiLF/ExkyuW8+HrllH/Q==
`pragma protect end_protected
