// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:35:40 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
mb6Hl0MB9/8xDIWZBXZC6I+jogzhwzpE5dFatFc+4SmLDfEIfTWjhg5hxFeZSCEk
kJ5ARmTYxgLZWiaN4gN9hvmSL4wBgAu3u5L7EoyV3iMHqGWIitwHnwiZYEIW+NsK
12KT4dW72K8RgF3YCBgcey9NCyWidFG2JLd1m2MSLZY=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 4816)
cL03W2ONUVrdUSy7FqTLpHmT2CtYvI7AN0HknSSS7pVIoN2CuuZ2Dz48QTwtOhFH
Tn73m4G1c/2rf7FcbC2Mh9FeYfxRYmLtf0+CNXlUndnEyWcKq8p5HUJ2eyTgU3x4
XBhcK3/AELajLtxcnw0MzC/OG5Pn7cEjb46NQWLUX4PzQ1Ot1+m123xiRuVzPLh+
YFlAT7gqEj3yMu4DZ8q9CHn4dE7pH0/lQRjppA6lji0bWEFsnQ4XItD1tsb7+nb1
6NRlZn2vqKvJ/PKtMrIe7BHPXgTBrM/0KWEv7tVkRMbzJ63M6QF4QbxnaG2gPBF4
YVCMUXBGH/uW3HoFEoDYMcvKkR5g0obuq7EluoX3ccdoWym9tAP69Vy88g/SK+/u
I9O1hTEAvi/uGEqiLRMVIdcGI+GDM2XkH8Yd22yOpvSFvewhGq326yUAhAzW0CVS
61IqOHgrMS8uIlRJe360KnKRjmA5cOFBe0hYqoIFo9FrnmD8bJOyIhDTaG4Hk+x9
hfWw5xjDwrWthfN7weRmDkcvhVZ7puQwzJlSV+owutZ0Rfj1fGG6b2efO1aSPP0L
UZH+lMcjLPUxKLhDZZHoiNkfbw5C+ORfZLAQVqBbnYL/wD/J6kJARcq14/iHc9qW
k6RcdkiLY01Pg6h2JmVouvY1IVl3uxMTz8mYJFWc/tFOjFMORi6a1LNONP/59t0x
Y2z+2iv2Pp2i2JIfg7vcxBGR639IP1poriZzDz/tRj7fRycc9ZEDa78O6y+h4FEr
Jy1QcM+jPcgQyPaGoUrXykW28Y9ooBPDM9oGOAcQAVwKE+c/2B1m5HdCKNAPl+wh
+hF1xErfVu8Y/bk8zb4Y1sAuAWWEhLPP87zuOZUugU9nh2eFcdAlW6yZ75Z+iQ2e
9I0cChSu8R/qm2PEvD09NxXqHEhC28kd71kvrBg4uumCV9g2PRflR+T5rIpEZxzn
K3S3GUz4LR0I72TF3zahrA+6WI6orYEV1vWcLNXEG1SfMG2/k4AdjKKkn1j3rlPq
eR7tb0DPMahsKO3CUoEgZwPiX8y7kWUhfiumcj0qxHcWPRn94NhcqTVPgr3sjrcK
At4YWJZ68CjtjtFXjpsf2W0iDo0sbwQLjGiV6zrK0uKdm4nMnlikiGc2B7jzvMTv
zJznYKUtEFzsHkvec5krBrCg99+d18ZIZyC7kl7at5C7TkfO0Vk9c6zJjzubFo3R
AsqBArD9DNGUSFbz5DMVxEHNkCsXwtVXiKcGHooM53GgjiYohiwSHw5q+zTrb0j6
q1fkFur5UCwYXg2LaljXT3ss9cPPr3juv2TOgEm8uaXUX0NihOwYDvwYBGabaByQ
DUMZ0fRbUCBNKyrsMCcbK8wxVpi+eT9eqHdLVNz99MDcLPMshwIwsYlr+2g/FpIm
BY+poKXUpdSGcIzzJ4kZ/xX+OD4rm1UBTWNM+t1j4u9UZxQAaHSw9HWe5SGUzMAG
YqmWnfZEQNRhKkkmcR2crmnh37nwjVnOp/5uQRtLKEJxcxN+ak8uwk+mDIEuiu53
I26LMUNN4K5FkSm4yCMxtcl+SU9tWgYv45neCQ9eEj41On50y9aytSe5/OPsfp9T
nxqOmKC2m0J1uPgSvbt3Faq1MW6kIMzXxcsvYj8uV8b1sfmJG43WIqfDSZnv56tH
P5vTrWvmvXr3Y+1obL4+sL1r/Xt1VxuJhjciTLGQIHPdic0oRxCIhw+xbsVeCxNs
vkqKCHHNev4LRsMz9E971w5LnyclWF9r5JAlMocA4VkosuUkRzv/AA//cuYnfrr/
Oizwyb0WphNPrVKNzSy/K2jWonNyWx41xyWQbDVjW4+I+yls8VsnPuA4huQSLPcw
3YDgDpWz2n7LtqBSue7gfVwsyFi8oKhv/FDni/QGEHCcM2RmlUCePz/7tWn2FT9R
msvugSqdn/1iFiIC+vhwUs1b2eNUUhtbNKd7DtGhaYuqRvYuWmchWJoUUkFnoD0y
yS39HcstbJLeCj3y6/lSyOns8QVfC7gzK7lRkZU9Lttz/fgDtXEOfINyg/A/BngE
gFBKxTBN5bcEqB6AjvGOczjEiAyQ3Sz+KCY38Bn31NRJQq1TVu2IjLk6pUnwdRAM
Rl4cE6vV/g7LnL9WALvnUjSWIk9/wh5vPISczkwRQJb1qXewji4fxIvUyiWI5ebb
MSCHQ/u4ELyAT8ZbNrb1H2+PPTrmL7LCKx2zCfefxkW8+kB8bhlAjGi0gewnhat8
/Q0tNoCxD6jNvbTTJs6fA3yR3wyRV+TzXgbJdwehDvJG3J4N3rOZR98iJFPxi72I
ba+ZTCt5B1Zh4KQywKXwE5FPI+k15qv3mlIgWUfVIP+xV7ThOVkVuAT8pRBJZua3
CrGF7pBtLLoXuI+Jb2o1rSf5KoBkLJV5pK/nE0Q0alOdkTmIkJgKYi0UzZnV77tI
0MfgMpfciZw592QaddIPc7tLbSJKor8pzYO0gsdKWKoW2b3ObK8t0VJw3rPMm8G7
UKVWrD/tgzrwGUHMe4LYY9pWIFY5OSM3oDb8spX3ZmGPB/sfshR4R8DfuUeoA34B
XM9E582tCyeGGOxqnLW4kQ3VVQwXoaFzqndjvI8T+ltILknOCANYvfXLG5NvsgHs
zbw9oHz7/038CZiiScpm7z63RUbxGNfMtd2ShDCMxJS8bjS+re2B6RWjnkcgwcr9
YIMvAEKfyp3Y2lwheWTSs7fv80YQvGc6KC6WZPf5pF7RGmk1HANdbUh6hHHNN10K
wfB0djiQW/LOa60NJfTpiFe074PuwxdjWzQxc4jM1Y45nfuYq6KGUkkXGk2Np5Xr
ZrUlOtEHsEVxCWX+7Jd3jilmVBFonJVzStUkatxUidXn1TGBRV5YaOiXxr+eHKfG
anXR5j+UtxHwo+rEf/8iJgw/DiYX9uxfsbi8TQxCrwBddGUvDEaaOKp0Y8kGp9Dx
fz5f6OCYE9BNhgcnTOCsCfr/hKqnDgVqsA9GG8HeOVchE+X7Jtfmw9OJCGhLGyH8
/gDK0F6cibwEm32cJKKbocRrDW8RiVFFhaPU19TRj1VRkK6UpJ2eKLA9mBH3NNPT
a7/+1T0lnTT6STyl7L/Jb2YWs564E/UkfO0SYRRXbVcjDcWm64BXr+PbkmJfhqGJ
a8yh/4KcbSniWYFY+UPBz2V4xo7jtOyM3w6G/xqmmrpLfwWgki00yHmeY6/jBcUj
ToKxI+YeqjcBuiw39m/yA/I2jjW+V33r5xCXO9H0DXBMn/xi6RACS+iVJWIN5rxq
Z4jtQ/T7t1Tzbb0ISUgv2j2rZSZXvIZNRToB9Ym5qFCYYLnbmG/+yhLIOaoBLUpV
vDJv2bmMUpvbfQ5hPocEH3qDiQvb8+uviOJ6Op22gFc2ctyMpfO0JrXLEY7osMoJ
a+OSU6FpqZgFvxc/D+VjCe/wvpBi0UiJgyPkpYbzQANnDDlW/KhL8uuj7qBuTCEE
eK2b8YnFxzjyPctCqQ0xiSv2D6mZLZQYwtzyJ05qEDiJJsgmPuGebP/pnf1TgYCG
ny0Yputt23doz1ogXux+TDuIcPme70dNE188wWCF248vhkdgO0f3tGen9a5lqlv+
I/jZM8mwvpnmbWGCyF/q93OF0vCrG7Wu6uRR/ZkgwqsP+vDrtNJAhlKdB7D0J6yd
wACTERgW7hkLqafBtnKnDWhYUQiwZTXcc35OFtmO4C0wPtcPeK40k/NdCroaM5CS
uIceIj2RTrhWEzdk3YocdGnaisZTWputGCqmOmPg+zqCd5GdT3cfyKB6/A+74TuI
67anhSA03K2xjniNyjGQU8I0SAX9/rufC3+N8xgAAQa63LSxHswX05tyvmHOGWLG
1f8UBGwoBZul+3vOYIwgv3BdXp0Xmd+g1N4GL95XqT97g0km/Yi1F77C5+LeElF2
HvW+Q/MCXjB46POg+9Ddnu3xUkSt8EQcWKxlV8xJBROtC2bomD1HrPMAV4XglGBb
EDSqCJcCNXvmdQUZABLsSZVjXhIecg5sm2NF0n58oLnTQV4Y6BMmatdKw/qvBHc3
za+4ogBWkW3RmqpQl/07vp03QATd5FnQ+7Fdu5PsK0xubDI4TT1cfZxyHfPj4SLP
MSrOxvWkQe2LrZt2kJ47i1l0MzBvwRZLY1YQNd4b1Cb80vUNdfdmkZltW3nKR+Js
OHVLTuVRYztTsVezDU5bRL+sx4y3xE1AGm3mISY8dBf5m5oGZfub5sstHBJjK7+S
01d7FoVqLtTMSLLR4VVH0AJXDNKEnRHYzImBP6L6BgSXFfBpFO61qCYulxcBV4a3
cJOA58qSzTuJ3PgNeqIjeF5Rsv/NRfJOaD4TSQf+jC7rx9GZ9oJ3xDetwg+mtc71
+dMV6zKFVZypfoPJFDRH/zHI0+PnwMZ5yGJpr7jqVGQns6vlnSA4Gnqkx+Ddg6U4
hi8nBb+PELQjBzM62Mk10wJXlLuP8NRgMbXacuHYXh7QGgDsMX7BAbGTruC5x7Z2
97mxtc7Os3jzcZNlRz2/sQMVYVrQrw1wagp1oISsZYbeKUT8fV95MmcNlPgvsF+u
WUGudWgzeYQq/MSRLvsL2sAa2ls7h5lgOJNLsAjNGMVApzPri1fPRrvSucQr9BYk
jMhf6Hx2Grb9LOUCZwo/XoXy4DD95lxmkyxZA+MI3NfF/DtA67516sNaAZCFJm1j
KyU3a07oMLiVj5z3DBMbIFCP5Y9w/frJ7uyQKmf0EVYLMvvXQXqe+HjbKHIZ5h34
8//0S6RyMv0J5hgRW151r4S5gbHpkr5sKdY4sjwo90TmIcQ//RAFOhNPIgwLQpLm
6w/u/YhT80WsMxOWCc8FDR7AJN+Z2Cd+2qEbuRSzaW5GOsyj/7/Y6P8o8qi/F1vu
iRYifLMCsg6ACpJj4zWwFbzOYODmjTh1ML2DxMARR+s1gTpss8myyaBzZc8LePEw
buERUaTMJY4WLrCAI6P1EV/cOx89YrKMk6lLlNk+xQcGpVienbXYzhXnLOYFn9GI
jpJoNFF0jBs49Jf9XBr5Zhg7SzARx8B1x8s/bEKrHrC+a/VqEZt5RAKc8YiGQIn+
IrGgJYXd1zI+u8+ACkph4TGmENOOXDJNsHTs3Mtoly4XaJE7JtCJq45Sl51JBWxm
lHCtFKvj14V+INjdyL18A3YOt+DOkJcY7ViNFC2LILFCpWzNlfuv/MAgrdb89SFK
38exzoCtuYwhswkMtX8KkjhMD2gBMLPCThSHKGOfq8A8dkUo4PQFELGRkbcQyw+g
uENIxa0U2qaes692bLX7dfpYZJKmPimfsBNQpGf+kX8wpX68wQUAMY+qXHPQeUzZ
iNQE7BVycDFGwZ6MtOGtPYR64mEr0Hmv29o4hM9zPTT+BgU5CYZ6bCDXWWy1kxkp
Ih0kICSO9vOXRS7H9uV5OZo0JtkEWvH7gQWbvHy9X1pb/oHNrGXfKjAAE5AP+S2j
TljTmUSPSC8eJQX4LJ2qfEv9a9jxnwXIT1KgTtdoYs3OuZOng5zpH4Fb6WjH8Jyg
px0f+Qken6VoEHzvk9+z0tGtQZS9mBHWrizeR13bh0xF52MO/JTVMKDr3A84USSz
oRHToxVFhkDsuMPcwHzGfzLVKYS/Qw0baBzmn5/ji3Vnx8/9PglJAb/S4ecgmbgf
4gVxk96QN8hminYka72ZTpi6goF6dlT4qTGJvqqqX9fCijr15fUs8V0CYMt/fNzp
O/jaFsTgLP+J8rPvtsSwBTvhZJawLrq6i3zeW6Zl/BrfUsW9jDeO+1jugXCX4zx+
aoj7apUDFxoGjBBq3vZkwNZpZm0YIg9bESWGlZUpMBXTPI2V8p5bl/zc2fDFjU4x
b+kerOG73w737ZBH5QO/DlTzS+MKsCgbDIdzsYrAV7GDxov0VH2emEvvtGmEUOxF
LpCYQXJ8QaNfhmY9gYpm3NPautbtgpnaHLD56AcxfT9yEwDC+W8SIgyK6HVPi+Bg
45/7ceG/D/XajgKXjEICaTec5iJv3XlG/tcc5PcdAIWADUGgsxUtlZTza28mWoVF
VLG5Mp68e8N3QWhKPe1Ohig2jPDC8DlEmT2EftL/65v+tggD0oQeykYVonae121l
VFFHtS3GxMQbTUGVFLUl7aMybGOY0Ds7xK1zaLkUYanI7WoSMZnW6DxRtTE0wGcn
UG/dtMezd2WVc5krfITpJbNktsA3hNwdvW4S/rFiZp8q8fVaLNwGYGkWU8H16qMi
jdwtyvuvcKmHFJLU7edxvhN3H7XW1UBppze3AuQ512Ax9hsPVpDA5BgrFyXyTXmE
0qijqsytGJvVx7k0ThWunbwpx1/RZ6od9znGsaIUiLa6N1KDyjoWrcPrXY0r0ovx
F09r93dS1I0k3sLdRCOpWuTlSP88WNxBsCEzDVtnLqjY0xf/6WGQ56suVVnRBiZf
u428NZSG5tkH6LVNTLM+xw==
`pragma protect end_protected
