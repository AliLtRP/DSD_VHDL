// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:49 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
hIG2Ssw7JYADS5kc26WdHpeZLWiFxDULH4fGdbdAFImbTfMNWRzATTelPZsf4Pj1
i66HVNBSY++scVjNxcrar+C4NiuPEeD5ET69/txxp/hkkHq4SAG2mZB/haBPRpEW
WHtUnCAI1CVb8kCC2//oGAQ/IKdZLKrw40IXkRloP7A=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 42576)
bzfN1vUzdXMXZK5Fx3Vy5TvfW0ksPEmJ/ikZMH/xxPk3ZkWdL7dKeJQ/N93Gljgi
HcrQZJsxNFX67G9tMIAOFsjUeWis4qeJLpb2EgO5fH9jezivS9BqH7UFeI9wXjzh
UIYS54tyIgnzV1w7Dv6XLIopg8kbSh18leIdQeYe+A3VQJDRrseSl0gM5pujqdNr
6qHQcslY14Ftr08k0kbKX7AETkyGMiBqjlQtP+YSU4TLqr4xtUjqoKyJLvm4cYcx
MselxrdknUlhZQrR4Lf9mwmKCPiEJ5b8iGUHV/QPNZfPWAvRAXwIcD1kqcwx+QJ5
2trCx01FWOQE2tzmAFnPU8BMyrKwGtfArl70erG/OYAf09PYGV5YWQjMo/Jhi6dG
pua3OssYBfexzabShcIznebZZQ5rPjCxbpRTLLtqhDM6BHk+ERmvmtl2PGxyvXcm
mlmQMBmVFDBoMszO2f7AOfnG3y9We5vwkUTG4R5xEKJzxsmDrmZXQWNprjHL6u/D
rVvw95+yUe1hii3jZOuxiPhjJrVGW5U9BAMvY4oBC92oTP+zA1LALpTefsjFbk4E
8YHtMGqAR8omTS7wg6PklyzXhLEkLfrx2OLUhxde733leVzlV4AMSBkVo22mP3js
ysNfqB5iMdPNla7dqgS34MtwrVRlWzagJ02mxKiEJhY+sIs0nlkLVopZIFGS5tAU
lSZY5ZFUB+EoeKEqQR1IbIStkxlLlpJE+XNwtf8vGCn0kXkIOO2vE8GHq8rUDsOH
PKY8JBqtX8+U6pIP0G14R49Ur0i/66uBXwlDSkD3QUVuQ+Vr/YCYEpZy6Hdz0dSe
1IfGwpfRsIFpbG/Qq9qN67krl1cj6dcTMKZYfl2jz3gwlFjsqi6qqeHHf6LnQgfh
c0lqOSSX1Zr3SWTJMO5yOwICeG9d8+LK2hLznKjRFtpggEUYuU8SBlxMhzGgZiKA
MyRKJt3S07TKS4mf0IXwzVUooqUfnPIgUSb53SlWNgiRiwK2sU7swr4oFku6ULLR
/JoeQLLh75xthUG73A45bCJ2R761/2v3iAjKbrb29tuM+WZWL03V1tmI/srbIs/P
+6hIK7Kn41ulg5etuo8xusDeL4QPpUYb8YoxZhnWnSoGhoF8Q80xGkgbp6kSTF3J
+QRN3t2bf08OYqqhpTs76m5pXHovY8/lXiFVHanH/49VnvKAYLS8/xv9XFqiwP2+
bwh+j1ccZYtLWnhTYxsDIG7AXz0HMEmD300/QTa8RetqOrdvEt0M61575bE7XzMt
WKLgjwaTATdMGK1+LA0k8VwQy8gh5EcVQXxMP4Di39LxS/pOny23FIaIvIoRYUs3
Ekedy0z3vLEoBoiwAl4JyValQssZdZYWZQHqNGh9KAUwZy9b5zTQR2sJ6mQ20SY5
V263NrwJactQuGtd9IwICDqOUSqGqtYyggKMvDYmj3VH/J03+LnwUzgDFVI9tVEq
tXUvlapcY4+5wb6325SZqXuTe53kGXhITsryOzBukL9m+LFjHg9oATKLYfIKbMMu
2JS19SSytyvHn2NeWd2jCuxMdSHALd2lkS5Rzn+abn4Fz0KR4PAK89WERa5D/uv4
kia5Qt6JhtjXGLY2S3JVNqs3mzLCGGiqwsnM5LezBGmQaoL1f71hBTwUXxhBnJFS
7J9zkxomPYqf/0JQUvuYy5gWwmRHu0/2qHpqguhd49YWVxvZAgeLS7P52OrWO0ih
/1TsGerSktAXqSkgzqGOv8Da4Vrbgn5Lr1aSYSwVq62hNfUExVeMR8R6p3IRQa7D
vxp0QWzo+muV7u6Nh1inZqK4lnk/zcfXEx+DmdzBQgiX5yivk7JgRSfbo0h3mxQ9
sT3w8rS2yPTcN1eYrNv/OeRUlPLVqJwN/tjQ7jYx2ADkhJk1huk2apE323fMGlY8
UzJzkHHjeFj1TRrSLGvt1dj8DtkNd+7Jz4RDguJCOMM1pUqp3O3y6mDRk8YIifBY
1/5W3/H4NgMMGewvMrx7qcTLClWiBfMpsxMYkW9flS5CTh1zNzKXo99ES6VDVd6x
ptyGt+Revle7QEgOANSsui58aaLy1zd6JYD47CxvUvH0qY6L3r2PDXu+MySlHwiD
Ujucnca5JsxjlQTy+C/uoEHEtEzc9Ee1t8iWktBUd5Mp2Nb7jyaSG/a9f/onzEjL
k1U8np1jkfCKUVw1kcPMsAtGWZ/9SQz/BQhwSCXFfYDah/yhanMVncVZpOLvO2HH
/coTJ+GSY9xIKgeA2/Xjwt0w7DsEdqT4THZn3yMlAwXATnZnYDQkz/enSivQCQjc
fSU18GgdKtaB4/9haTYlyHEGR/36heTXD5/XG9EZdIQchLx3EFLbOmLqOyNNZlSp
YR3TVz1P3rZDw8vfKhP5g3PlQVaGbnppcZqMD1SSdl2zX0bdW6OVJA+UHz0zfHUb
OMQKJNxs6Fmx4ZkoRZdkCV3lNmhtgcUZF2I3YCz037f6tIdF4AVorQLMnuL9hEAY
rVHnjCsyFYlvu+lm4yynZBq/6Zkddj4yFTQwPlfSRXBV9mefDpMesddMewdVuU7R
Fxb4sl5kYv4/f6YXw3zI1tgCKBeDyQfW+rbQS7QUAU6JWLEKzaTg+l/Gv3Eqaals
8fdVrwcEliEPfvKFOfkpHIJd/mqOESSsBbsJx+H9HCW6kxYXKhG0QWp0cnOjzrgm
xK1XtibwPDpavSPDf1uo/bfEWX0HX8DAlP1TBfjji+deUFr/tnXieDuepkDk3w18
M3rgaD5qAZdPlW6jqpudR60xd3br2MulrQ2lglx+VfQzWSEHCuBdHtBrwudiibRf
51bNQBYodVNLbqJU+6rdphBlygVqBOECpzG7ZjliYOwuB7SKIrlcg2xewdqmgmUd
9VWYDMtfNhcoheakGy9AWdT5m81EqAsAtlR7fEuBcmkv+EFyEHdF1SplzjNRDY+r
sFUtsJJJFn3BzHF93U2iXDrkPEnlPkKqPKykpf6ZMl61a2LJEu4s6CtB9Qq6TLHG
47LZAv1IT4jOCcnydTHienpZH1mGYZost17hXTEwqSRkAydrfB0yvgzueqH16ZW/
+t3lKCf9NMGyWrrbTWueMYgf/yPSIOHmY+9CDMww0FaIqYxt8zuRxwMwrBanmj1b
XkOJlWRA6mYdKYSZgPPvRege9WWR/LTC2FkUrOHiS0J0+u/jK0a4Mz/Gp2Y6k+sW
5M+gBT8064CcnqNbcpKnfx6x3RA/NtdzwUFs/+DnARt9VRs9GeCYja95Qdobkxp1
Ut0YV46Z+0qqG5YTn4lHpQME4RFDufHw38jkNxarM3GycFuOVbn/Ul/FLF2IovQq
Xj0VcMA5Ah8EyDiproZzNqoi4KxnwVtwykygMd3n5vxqtby2j4fUlctkGaWIwDdI
UbNI3gW18O2dtP+xZqPn5IU4IOhlIy8a9+aiCreV6i+fJxnfoOHLiq/HD4XH42y6
e3FwjwfWwXv8apSCCcric2To/6WCW3Vl9h4A+hGXYocZNm/gJDUNv2AftJe/h1A7
xIRuHs9MrpOnJOgbIdMymbKio62UzHsT/VLvj3/env5k2OAazf1L2eHs1+9nt5R/
FduVKC4L8MPb4qmatJz4pv5FlCOYEtqEr9Yt+Leq3qIJJeN3paG7wBGdMZj0CfLr
Ca1knirvkiEfHgEwtLlo4Urg0WQsKKumAuBcojVIwCiOsMYKg17INJYUbI3bDHgQ
903yfrZy8AOB28XzuxwU9SUcdkPWmEmZ1q9Zf0zewSoyvdBI2XLLyGMti1g5sp6c
AMwY7lQnP6/VeJOnN7qKpZ0BgGVqt2ESVulzotyO8rs5sAH38NHoM9xu5KqqE2Ki
8mLvHF3tW3nGX7j27YdVG7hks0bmzRrFhK+BCiBFJ9MEW9dNK0QMC31cQ2TD/DjD
UUVVB1fpTuvB1OYC6oVww8v3n8lTVTqU/un1LDVwfPOdjrYIx7VOIE/Qo/3MI6lI
yPEuBpvTRsioR6GW0LPO1c7lRD/LTwadCvhRAjw81/SZPiFl4Kje0R4gX+zN0ZBc
/3diSJSOuZ4ZoqMhd0zceLSgdgahUP8HgwM04C4V3rNAk/7aoqBaJaDxhHjKku/Z
pib6NowxpB8TaEtm59MczxxicWQA3KfpNCQE6fDhjV0/SJ8e9Ven9ojg6hpLXBtp
IHWpj0sDbbRpYS6WfV8C6QmkRU1aMm6Zt0cAbeN0aLGcU6XZEXzi1PfmkVxZLAjB
8tqR33vxtNEsmURxqaSoWfLMZGr1DlZCHoSlgYpaJKdpyFdh9MrGIXM9siwS636S
4RDaftbpcxBkqco+Wu+ICxk1Bx17HJvpWM5Ka43dXVFxJFQgBYiZpC/75o7Kr96U
2/PgTqpWCSdysv6FltbYj6ryy6hcslAoCe4ltADYkO8g0dHUqA/geeNibG+gJhnV
j+8AXVvBeQz7B0lT14Ih/JEre5/RINzc7AD5SBMRxVGbq3hRAa6e/q2iWnw4uj26
ySLlLEtHsYL8DIxGi8zwNAGpVkYQhF8i2q0Z9gOdoSPgymTg1djr1kNsosEsFGwG
MXQwhXpw+s7+fqQLanv2XbRhCmRjKNKibd06Jjfn17ORPAUv4Dc39bZfgOOXSGcF
yjnCkFnlVi7OUIfRhIu60i9g5ZjO2KSpCjCmkCkQZdWST3yw1VbbG4qiwsoRy61r
pgfi2jC4KKBRHWCOSsTi3oKqDZ5QgHBD8CIgqoDje9EGLibYdEjZeCo+Cbu2YqZK
DoOqOxActlPsk25h/gIHX33pJQ9Els7j6XBOC2BLN5PHyDlXO+kUKMPrPRIz5J28
Gf337bMYFV4H3elSE4mCTadkQwE+MSHEEBphKebZraWkEMyCIPl61Bk6Q4/Nm14s
ZfyDXl3foQcDMxZNOMEdOtVcsJ3Iim81G1lNTAX70olF9TaafHTnTU9EnoCM5LmL
9Y61D4gn+8RB82OchTqYKgrRDkXTeBn+etv+bvC3+E/zurFLdWO/682hEEqTtxWs
ZPbBGGKlb4YnqQ7lICqqBhviKfNRxVX6Eq8YmBWtTUjOXFjCEbkfIFshfNDo4Lo5
aVzSJ6tQ0fmTPMGWOlIO7VqaThNjP6c0w7OqfUSu95McXWMQftopA45dA0aLGcJx
3+jUiJnxXTatPvuJo4ERjddJYzXYqeLTT3Wl0L8tuA3aCzEof6JWlUUHCH8Kmobr
rh9zzdMPJDgkAWXCOnmrPvfoFDUifQNDVsPs8GSelEF48XEyk4G/UWJVMrfqQaHC
yMQ4HIkcDR9TAe/Ic1md+iHi4SPLcQJTvP1WdGAAZQ2STZo2PKV74T2TsiM9HpAv
XLAAHXPah5l84KRx76sVWzoRlxfvJgRpM4GthlT4d5zawNe0uZG8qyp/T7mVtJyx
UnLalpjhQ7WOEuGsbh+0kZXUtm45kRjX0JYeTa2Geu+IMFzuw5ljbTy3Ux6SLWPm
BuUIDha9gMH6UYVbhzZkX1vLtIoaL8qA81lbzQmi0HDFcs9ncQ4uHS7zv8zMl5E7
GInxg346n0MuqfofE/N5qA9yZJlgtx8KBaOJrwyt2cQ5jZoMnOTdL1CfhDI15B9e
i4YsNs38bK5Exm0vkQneD/by3KI7oWI0jHEfcTgSExHMu5/C0eQuzfiEbgQsIp06
+4MR19hvMeaedM8ZgY15EwemE24Yhw2gPIsGsM4x31aKNdCzh0CfuJi/M6KUCWJH
ncD7xh+Du/sqGDoCkl+7Vy4Ay/b72TxXCrCGon6G7V0qRXk0eIwIVIGH75J4Iwl/
shwiG2GK4eb9uxTeoAuZRK90JgkOrMRqGCH9ZPwSyS0G8NEjv1zC9vNxLTLY7yIa
omXN6H91k1okAkqFE+BQlwlAXfN61TyCzchl0WGQwYhFywjY9QCYBwdTxUOaZOmM
kChAMaVjxuQ4rnaeFbkfEyV0N8PCgVV3EeiA3jETcARlfRtGcIk7X0gRwQSD7+cM
7c+//Cy/0thbY5D21LFNG3TeXSWy/heoG7j3fMp/7SLWnPNMzjaOBLOJEN29fpqv
JFKfPuz0yeq0IB8Y6MpjxjTl0y0bPPzcfl7fE8nFq9AFt09yr0bx+RpsAicp2EqZ
Nr8VhzxZz3x+ZdsSJcGaJWfWYyIPn0iulDTNoUaCJjR4KSJ58pHltLS86+jcgxQ2
HBHiZYB9gSzZJ72/JeY3QgFwyYwzSlAvHgIaeLixKqhYkoePh9JvUNtJu2/r97/F
50HHfNKKe62im5NS65b/YOlY8gE+yZrq3QgPFe693ZnyOsLBgJfSpTRv13GNtjgk
u+BVUGaGUOGA+ZOgXnGbZkyEAPH821TNBNDLk8j5BiY+HZKKZ28xYuctXTeGWwhA
q3kut6612uXt+5EdTelOs+1G1vpWTxuJyBg6RjEtrQcBq7a5wDEwdZrYs6grXAaR
UGV9XD2d4+vHUVNsPkaBDg8lRbUoon9gcVFBWelLj9Yegkge7Ohc5xS8kBhyR0El
XhJCnDR6zF1C1MTgTelVihoKVc5d7vJOjzoUD+zP4UWMkbPQcBjsp2Mc5RySL6qU
S8gyZe7hYKWZfmpCq7Oca/BDhhkUmfIVoBOlm5K3IMmwuG36eXYfguOWqsKN/HXA
6/RTh1ycb4VvMTA4qpV+fin8WuZs+lFKKwCWMWj+NsD787jNrnxOkIJLKwMbXAWG
Mk8Mh83Klge60xDwybMRuGrvDyvMVIF2u8+TmGrASH5Aq/9an1W9mf/cSQUOWJHf
vqdyoOEfKGxF6J8xIleGDonxjgNv2zc2ZfViUPRrpGp1J0+RNeUA2jak4MtwGJn6
rgn9IHlO20lmmXXLf3558836EHLvQ50tdRNLEmR5Mn6P9hecsTO3nAX0J5UZ1Tv4
G5yKP1XyDEUlRRqE7Q13cRPoal+0qjAlF+jE+frAzYdxFh1gyQx5BGoCn2WTWOdR
xJIWNow2zGSC2v9ZstofwzJAaXcrYZUkxzFWag4yYsxvzTLa7VpK1pCKVt7jzwJW
jIXFocPIgPO6Hk+dhjSGMSNw3gycx/JNuJeteNllr2qnirBKHYdCyJPNs/mgABjN
8DQngArggfCWEICjiVTYCnuuoxKlY6bnCcvCxQ+WuR82vbsOBNNb/nf8p75Pphpr
NCIR3b6ULzn/y1Bb153OXCI+VivtZnzAUbBPhsagHYbejrjvdytdE650uOr42i8j
O6Kajd51Swv6DKd+nda98a+WHZkmLY1Ahq4X+Nt77IkFrGMEM8l+S4MRtt3OvO3Z
ko/Xcgdwm2sNvV0zPcbICYrLd0fg65oEBmcoaIa2wk2Dg8MdJ3JNdJdyyQJDO5S+
o8vojE1Y50cUeDCbvvuQv0PKRyDImMTcDaixKFZ3o1pgxe3uzwustOfgukJ5Cgdu
CvhayWEaW4WwrjTU6nBL32KSpnp+H78YlgfX1z9TWc44UZbtSYNyRnoNoxzgg7Uw
D0gqfvJTWKbpCVWkv8XlERa4D2clWxsk7/kysEQZE6bFn2Bdg2zg8x5MHsHE/GOQ
BiOXrCyCn5zDiTvra8+hOA98S0OMlKq8HxhRHc5lYMirTbaiqiVmKDwzSMidtH50
tklW5NDTOWj8o3fxc46nRk4SuSO+4bC3u4ab75bFT01VYpmjx2pYE+l1iIh9gDQN
wZxCNtQ0LQXesOH40GeGu+NF9uidrWD/CUjwyOQbwGW98RO98SDYeWyMR/GGxIIs
7PlAjyf/grz+WP61k7f+JM/JCLDfIGANjNi32FGSbUKXYTF0GiRt6S9dF8mq1LbL
uq91eaQ3MFV5eG1MCTCWg33l77TsWz/8kB9i1f2D6zdQEDE377Zw94aGw/rC01em
r2Jp76MFVh3fO7widS1XNno8pnv7Qt6q3c8RS1vdDEjzBieTAvI4T6AUc7LpZyhz
T9yBhEiUK+LcU0DOOe/QW3kj53eihv6ylD4NqzcmIMhJtWF/JP2nhB5a5dQ8VjeT
UQMp+SY8Qk8MOVhuZPaxinqrwcayEQ7kaScCy8DXXHP6BMA1P3tdE4F2oYmh02yJ
XggVeMtbbMMEnDa0DvlGMtACN00WhBIXeeXkV8gVBtfpABrohVbe/ecjcg8JptMq
EtpHV3OYM/XiGw8lAjjjgBVqiZFRvLVOV2p70PqQwiPLcMy8cwja3kE3f+RcDZbJ
zFQRcgdf02L74H4keapZOT6FlViCmiCLEutZXMQkZpI6ZJa3qXm4husWKUe3XsdZ
AlfHmHG2TghU6Mp1j/qy59E48CwL2vOC7wVj913ajkyXNCoxhcFEvov8tyt2rvvi
syHTVK6rpUjpoOSuokKCte2nkEOTEG32kKdvlea+5JRQZzelS7n1jYcA2pa3Yix8
RviF4FYkFCiHwq8EKWCCnCOZrp/CCteSPZz99YF3taYVwkfn0ZxcLtuladoSCtVE
EFvrpw+yETd7Lzz5+ba+o796AQrbs01ywFkc+ddqH0gn1LRUy/4O4uGHcIbejQ34
J5XUlceFbq/uMadX+u+5nJ+DtVXR7Cb3YoHwGrL8l5g2mQNhGfcPRB1k9H2NiKA7
03sKjWulv95XVQJYebmWCxGlQLuQdwZNKJo8a8HYt5Qv76NtWddrcoUQfEfXX/nK
DXaLw96npUSxmDhz+/uwjoHn99HMtH/wOz61OnDV9JFLZTKCSbIOz46qsCrPUZD+
02PRRkQSljUoGyvEQ2r6NBSApD5coYRxa+e+2tztQVY2pd+oqnMJs5oGn6Ebt5Om
p1eCv4rdfcCYyE+G0fSyhr9pqli5sqdckXqWK10+tVNcaAvRTxnF4h/vvmktLUW/
ynco2BU84UJIHzgfPYPf2KbABZqGo9CZGuFDIP7nPUuSxM2PuvQ7HhJyGu5szuFl
SVbVFQmsiTIMTV+2DTH50Q2BAQp8qullL/DxbfrDlp1rvKqoq/ckMtaiLpPoiuaS
VbQWbpFwn5VOjy3jIkurvnSSW/kLuTsH+kB1xDnmaCxp1Dso4qpLXCYRuzxVHsG3
AgT5L1AUtKzL3+98jaAojnGKKFb2Tl0JR07AzYp2QkZAVc/Rv5asLGY6nn8G64v4
VdyPg4stoFWt7uZFLh34bUDXObPGaPbrKzob7AecO+SXP1aex4/KYXiiDtqCpdnd
Q9KIrp+kdPPvgELH3rDjbSKp5N5z/2GCG6sO9wzE3PEHk5X8ljvCiXpcDr7hKZzE
ZOXyhAY2+xpwRvDsZsKhIrXs5yKrjQv5KDSj1Nw3emvkv1P9YQaBuvuPnW7zCn6U
ILVUt4c6hJuA1j6smBukd17oPZh+A7LAbRFQDIm5v0YrMw8fr1bs/uqDTdTbinq9
TEfnGdmtPF74fK/GMWDlqqm6KwoPeK+y74ZYVcaxT+NhSg/451tWR5xrRDgURg8d
XnwiJtHOhN6gQuKj5hoTFZVQn8meNks8Yt0A+AT3cl+cz7ilpGbcr5YVN/JonyLW
upBh6HeESUh2ENUoSgLTXsdPCqovVKo864u4JQcSsNIFJ19nyvGm2YgZnxl09hnM
YHkHj1OUli1cll7HqX1QC+GeqTD2w5MwSb+qzT8OAktbCaD1AauT8tR+zN4UtCrZ
s8GLN0OFccEn6+dOZUkz5V1NgsSAOGRvsg7tAy4JV969sjNYr/WwaNxSAY5ShClc
eAVrpq15zydosszR5k7dkflbqbAXmvLY9SEQUF4IaHP39cRgkwms+2x8mnK8mXQG
mkCugxanUtWFQs7+uCGsQax3gaF3tre3OqRxFXNy6aG3VkbLZMeYpe+N+Wstm3+f
xyBqDrN7c3W4Gu4meYkWummps/fQL4nbkoLES1v1s4aSsU134g/kebs0ZIViv14n
AarSde6BsFGmrqMSTxEZyL22KoesFJkKB0/bbZ3fQoePFb8Lu8r6/0ms0eBEat+7
nxNo+dbePCCyw4Ojn7sgcfmLEr8AFYK98EYenJ0u/XZcgPCYWTe+atrOqduJmOq7
loBNyTQ0a/fslhqNIR7bgwbvIqsfvfNqkxixB3MRR/mD8vTFOpWNrJRw9RNn//la
PhuOJpuXvITfEd/B09If37QqNbrabjZTpRN4T4L+4yEE2Jo9lttX3digqmr/r4f2
/5KpvfkQLNPrTEjfht5vOmAcEpkzFZwFuC/aK7LQExUL4KPLwqvhdCcABeBCWApY
9QokpBTupEzjsdLfR1UBgfaFY6KzrnmBPweI92HhteGyqR7An5WIANXA5uzQV+B/
fuxcRGM/SuzQYKn7ozAVsnqhCxzz95CgfSimDzsUxGBfSwqmahE8Z4VlHQBaGbfQ
7vfVmcAsc1BOlcsnbyv46aYS2vJWC8JBBcs8P8Cf4qXTAVvVJTIyIiyB1lv5e+M0
YbgthF2IBLMQdgkkf4+saBMxOfv5ftaJXeWB4QrCqeTRtgCjvWOcyOHLMkUYZR/7
JVpH5GAwwqA5ZxN4gwb2c2ScxJeEB8JOC52/KiXRk5o+/p8y4zOL1PybWy8DPQdU
o45ok1AyQTozRu1SgdVqU+ZGoZBZa4fFzykejr6hrm5iA9L4Q3dLOBfxKgMqYF8c
mHJ7Ka7dzdbIH130H/oS1aZU1nZSaX8cT5ih5lVOtTBld4nd3uwg64bGpUg4QRWH
HOMtEqJ65gIviPtLfNng7bd2WiUR1/NhPiJDAg5WYd5Cjlpcsf2By1B9cPgEOMC/
0GyJ65y5ZXzUQQPe4UXKB5/27HCO+J8qsFhgsGFDtZTaqkSasgNdGZWrTBhIvZnD
RyymJpCh8Tc9q+1nv7yDPGNig2a14UuZzxawqn7apXcNTS4fFTAjvj+ITBtTMk0L
H7dkS16vQToyg9/MhRrorIIanqp178CmtmPegkuPnR4grGrSKfDnnXFloCWFXlIC
1e2t6M7wlTS46YcgO296XNgbpYJpASZONXbmy7gLsajfqBLCblBlp7RZaY2n39WE
ePik7X2c17I3q3nMRxCWHLPk85rthde0Lo9KBmrtFARKv/Tu3k8qmD0/lDfufuHN
QI7hds8E5VwzHS1Y6v/mWkyRlQ4JEt2W790Y41l3Ys8FSITzv6TCNCHgWqNM1+IV
ebk+DQ4CwsqwFroeLGTb53LWE1phrgbhlMeqezcPWNKnEO3Uwfw/Dzv6mTo5oZmt
zjzYkLyjXAPzJJyvqVPYPOdFL2XwuLJHr8CqcSIAX53xgTpBhGFZo7u2suMghuMi
YIFQka8W6jxEz3jlD513DdzGELpGqXbcq6ia/xvjH+TTzyEHyp6xg3nojcKD8uI0
9TbNZFmrgfG7Hq4yVrxcsRkQj6f16fg31GDmYoXXWvefogAQd9sK70vQcNL9GK0R
V+BghFjnyxQc7Ml4mgXrEEtRD5UAVuy8RGSXTBIuWw2SzXPS2OQPpmUnZ38T7kki
/Ps6WWvZXwFnDV4vZMldY/H1eZ3kwOnPHYMtVV29AAHMjn3U+W3TOEZoLaDyrzUU
FDm5p+6omWQSRKiKDo3Kol85QpSDmqHig9yQYAmpGiT5TP1arrUFsZnQEDW29G9L
peCEEB815eYUhFdP4FXCAPxHQ3dPkdGP9b4ZZ3+N2bdatWJ4+gKX3y5ahtgJ0pmN
66WAGFQ46pLHodl+V+EssNRiR9zEaml2dRJucaGkv4gaezxyNOwbZ9utNpfpfAw0
fNL/UWsaHZlud6oOzV+BDIi5OWKrr8/9tuw4ynVYJBE58yWpHE770M6eizGe5vOI
BuyQW84e9sD2zWQMcKZHmTJUaAA/ElVGcTNa3Q4zmbptCQbsNNGXiK5U3fe5Ocod
mxmszjj/lb4tRfcnL0B484wGbSHainDd2wV3OoUottsNwh0WqUoUWC/T+lQJISqJ
olKVqYt1aZSqYowmIq4VfV3ymlC0Z6WpxlNkEgtn1LiNy3AKPTCj/Ha1AepxQGfG
5bzUGzRbrkgW+6PdUyy3kBelBxYGt+LBMiWK8J8V46kDnNzqi+z8K44DvPN7Wi5f
SqsjG37vnsX1ryqJLjfD7EmaiUpHy7+UCSAiMQsBNfiR/GQvZTpQUVe18/2fdx11
07OLuNTapTG8t9Xo3Lw6sFxQKMzMPyEHDRjwYNLLB09DM0r3njbBW29fNv5fkHDV
GLSQ4XSIcodBDf7YFljlNIChjiPqcOppSk/K6oLAeUgv0TrJQ6t4fY9YYQk7bH91
CvzKWw5dTP43H92fi/XMA4jwDtbVYuvBbgkm5nfxyawPLRVqQzJ313f26GwRguVK
VDlvP3PX/1GKB2bSjbBn9aAKP6p6YMasUohQ/HgaDaSo8eaG14dL3Lr9HVFR/SCJ
LKIeKiZ5s4A6u9F3EBLuL3LGYwFnqKs8ZkCrWCmX5lyv25EEvFPhnlz0fzJfwydB
NzcHsRpS21v57unLOzrlq8EmH0HCNoJ+s3A8/rjIkM++xtq4iKnquHR3QWE/PVhV
yW5UmKv7VAfYRrPrUardDVt/elrpsXiXGAPvLIcgFVb9vsWaA9Qxh0hU19ZtDr/5
/oriazlQJnAhbwan5xdhSCu6gfJZx1gTVJ5z1I0JBUEjbkOrPTaLnsnvQH1N6npR
laM2094977KUv2qgMxs1h4cgSul2aFF+PqTkRc6TGXA4kVgYiLFeJr6/XX1QidCF
l3M+CeWfAINWh6bBEOgy1n/UR1pbyU7Fij0k4pGbQsL2I31YoFjAl0RW1nA7VL2U
v7QIB92fGfkz5g52PvtMkjmIDGeizPyNBt2V0Y3q5CKAQs0Eg8WVLsOt42BnmDpu
NdKoMkbSJXrP/IjNBDbpSUDCONWfghAsVp/2CO1aqdVZlP2VtasnUV5sfT4JgX/3
PjhWR6ySy4oOjYoysp2tnbV6Qv2Sqj/LfUay99phFoGd4XkotoLyiTWgQ3W8Qt18
yvmVnRc/Xm8gXm65CMRCOW0+fE9gO/Exn//Te0ZjeWwh2hokfx2bVmW5WSm5OzUQ
zfDXP+ko51d5FpgC0xNV/wmpDoz/31q7ciBDYRuT8MkFURisRQsSZFJbnPTd3KVf
ymxGjW2/GcWvug2Gfr31garbjB6YsSO4s+uuKsA9U24oCZBvd1kvbggJetkbK1Mm
1FoydYqRROfnk/G7I1nS9M6E7ShqLXB2s0iGW6Xl8CKgBDPsPIYz027OMNTtovL0
jCqzbAqTvzXAAMAV16a7C0skj+UOLu9ZdV8X5/1hvSlIV73lJsMA73n5/ZGHq8vV
7e8JVTOUeSvKAKUq4UAU8BTLaE8uvJ0wLJJKuTvQyIEn/NXgUWt8OmFPAEzfah3N
mm/DVKVDPjvDlB/nbxfZh3sxnGbFKLxTH/bGcO++671MHxFolZjtXi7B+QGgQSAr
neVkY81IxGpCZW8nbW0pFcaDBWvxJTxH0YbHcYwCeF4lP9BlzkcYyx82zFf7aYOJ
Fz9gHakpTuDEmsJkcIRwUwLwJGhaDPujsIwzb4dl79rXKp57mRdHgDokKaoG4q1z
ikOlphx4rZ0eHhGZODr6AYNNMn8wOOkBenKU+1t901A53s9BVJWhb2u9ux03WgRQ
+TN5iPKcP4Or+RyX0PYjQkFNfdHJJ4wqqUAP4JgDdGpRT2V3Mbx/H9/tuP2N+NhW
Gk4YaM7IVPoHYza2agCEBmyjAQOoTV8kuOJU4NZFmld6bTslX5l1MzIu2nFWlWUI
u/Yc5rauGzmOMaiGWCKlheZNb+9sTU6z8ZHCWKzsXD5nxkz2PeqFMzdMIG+Lmzwg
0kzVFwGJF2bh6mhwtvIF5XYV5URQ7UB3o5YTFTviVJmcRioJVqLRf8Qh1iunNNiy
3IW2JJrNF2HrBiwkHE1LWQl/KSJao92w4RHxi47vyy2vKKG0wiigzdXtypXmfXaq
2Xg0+U4XVO3sTJI6r53rW5gh63mJlEO1nVVhnwB7f4cDcgrO5LDzatH2e+WJRH4B
/eB564TJWQGVNTw14SPn9SQSAJoUrDEFjo7P+9027RGF0AiHVGwpHLA3qpctLkBy
XdntXPEUucmWrMgxKzMw4Kyk+MetWJRv1tLKH99cbfr6HPLuoTv9EHf0Weo1N7I0
diNGYTWbUIF6C/OIDDX9LsXf+EQZeZvrUkU5Dh9LPJUEdXP7PaVP6tYM0TYV1rUf
Zid8ZDXXL9V4sRgk8g3Azlr0tavMFropHdk8ciC2bgQbDe3OzRnKWeqRQiweOtY7
1v9nxf7XHCj6C304tYHqfslW7lH+6XlxUQM50xwUdZuiy/3IZz8LEMkwqTb4SbTL
c8HQK7S4WmRA8cjD5kQr+HjlQCHVFGaPFVnqHsxJeow65I843lHE9K/nnHVvcxxH
l3AtQNwsIH201Qwz7wyLgeH3mUHxtqeYW+CYqTQXLVDAcVpw28yjnvYbFwQTTd6T
CbCIYGU69XjvDkjhoaCwUOaPoKwDtwXXGtk1SgwhgaVP6mxVZKcw+puNRJ1B9nrs
aGMDnPBTXHZr8HlEuxQAbYcjE3yLuhQhpFWN+49pYacBXnGEd2onkahw6gUJdYDx
+3617YA3+dG1bqX+DtjInD+q+5Ge4Z6vrOM1Xye2INo9bv8x1It0x4ZUA1lXRg9m
uaklIrGBPLxWDwsFqysYjSBc/B1Kgkd3Y8vgvpL8EKRSE2m5W3pTLt0revmKuSqu
ihhm4NgNrDHzpAih648YpxyrEXSkIQmM5G6Wwo2fM/hqCdRu/p5e9/dbwRhSmHau
MJr5G/oyBjO7vXflcy2uCizcKd6ZBllLl0IchKIQcmt3bY0YB2yuHi5sxSyUTUaQ
8VEwXp2zeXp/naeQMMZqEod7cpYk7V9mXuY9+CEs1oZfp/0bR5pBBtL0fpgUWlgA
oV/mjnrrVAsjVRr8yb9g5gtChxG5fJNKyVnqWUn5Uy6+sRHHFTtrYykCmNiVAqoK
T9PhHn+LsyMLPyYt+9Z4QDHI56/wSMfNTnqSCDxJdAz0VAQl3j980NTC3NhxWq38
AUY9lv4kW+kwurNyCMhUypAoFkSy4qnXMnQrR3c4GZYfgVOGbFATc9idvIGkUlgr
GMli1kPHwmRwyzmxkllYPe8p7LNkTmE8kboB/vFX2Q5pjMhtX0NRL6R70vsBKBXb
SJMyADTkDUVZ7Wfvc+cyl4FhpDo+z9cLqS4Gs9Y8OQaNWND9p7KklAQowyjEAtnT
af1TA0pTnzNbjQ7FiGymLVCbwq+crRJai6XFzc5dMoGW+h+B86+s038l8sLzqSvR
hSD7JscO4PfVAZwme4IglFBx+oudG7AzV0H9auEZG+9l15WDwgJuuVBIGQ8nyJvx
QSFoaFewGzEiaMd6EGGfM3G0maIXM1eOxmMpaQr1Wt2yWpc+Lgnrv+jwRC10Ma3m
W1IDgJfNRgGIr72hI4IP+9UmOs0JHcyI4hEJwzTSk+9kv2GVfsDQIi3N8SzoGBJq
Atmn4TaC88Iwa6c136x4P9oxuQposd3cR5S8gGYjIdThudL8JiTLxvA6rPLFnffu
kyp/7cidgp7ADkN6h6LT4o0VTL7rugD6k7s/CEsljxDVpCqYgwD6er7J2DQt2/TD
GWjDsmVMcWPqTmXQlgoGuSY51khov1vBzHY6jx/JWG2y8f0rPUXZlx0lwp+ZYKsB
xkPMlnQjS0fwygWL4U4FG4KpALC3h5EsKpegWHIc1mGWMctR3MtqM87lw93xQay4
NRvYmLPkEtgU0HnjAT6In2P6qBLLLo8/yKb4bBc8QMD9KTr33bBFsbx/jk/vLUFx
/2bjbwXLlS8/17b2fk24wIWk18dRqMwqQCt62MrCqsnol6WvHuI4ZAmmwGyGTKth
AMmkyui7fPViS1/NRgGzvimcs/V0ufzN8Me5R20zr4z7n9VOj/D1kAokCabgUF6o
a9tSVZeBx+ZwNzs1Ec0GOajHCXapqT9Yct0Am1RB60SkRAtUMHPpj/yjKp3VLf2a
Ra6eheFDt2Qk2iTYk4bnaGht0THeQxuKkS3oyUdmWrlNaAMDc+K7+zpnhCnAnnHe
lm8oOwQUOAN2OXqNf/sfxWKGzt88OYkfQHFFMnXkrfpPwJPtRh9G8mm52f+qyuIS
vAEzn+Iqn/Z3rsJUq8JqFJSMYLYpZbh/YL/uFGY0XyNBhDnmFLxiX4F0+VwF8DAC
uNO3oAdT5hl/Du8c7Yaiv7Vb9XFG2K5lPvn/rVO7KFHLRt+R9kX4jYaYX+ryMj0R
COFFbqXxsaLCPuLzIhY4vRnlQoND3PKKJxrJPnzkwR1QuNNeKhq5nzinZmzVgBB3
/7Z9vbdBuzIP23pCSiris5DOj8p2USjNGQJYkaBUuBaj8yHVcrfh9Vwd2unwiThd
VmCtudIr3snYx78smTdmf0h/2yRbpOQ/jzGMVHfc2o+EUAAgb+zfG9umRh/xkwHQ
vOgwnD+7Tds4NEI/ZXc0qGmY3jhJ1VVqGOgAdrUZRZFmdgbEj8o0SFZxXK1YNjAx
AsNgaYAN3h/pEhnAzuhPwnHe6l7+e/Tt4M36elHvjEVnVqzxTX52amamWSSPPz+B
WTQKVqyGTMbHQKClRdMRPoTIQoS/9sjbLbIspQpvQ4AQVZOT6IQKfDwRkPVGgQnB
0DhFg54od5RItBc2X3ECN7ONiAZxn3xAh0VkzMqmehVgRGn/emvGTduxxkW/YAqn
E/x8hi0WrR8hQ1xKWSVQGcZWVB3lB0MrCkRKOfP1dnNcUdKisbrgdisOeCaXESip
KRUueyKph127nJ9V18k6N9i+OQbrUug2eJvUDYD/iwHUL+Ad+wv/wl7nqncL9EOm
W8+UxvmM9+y3PhqU+B0iqkL3d+G9zBH7tymQQ0KB4Hus6jW0B4ymVOV26k4UcCsv
fmvUMdaozwcigRtq5A47HzggfiG4EQRNAJirWSp6vldfe9LAmVpkDIcBLODpN9fM
YgkHNBNCMWy+Xe5cpX/ro/s2JgqXthh1rW4ZHMxT9nJvyoMkDAi/F/o1pnSg6TOz
yQqGvphhKvKD6PFWm3pUOEvr9vNffvoSSkSJHt4jmsf6gDqIMSuaxqTAeGYmRUWH
mZitgeyBp9w4OmYq36tiUjBsMY8JGGBBp0ftB5EEQIMi57A2EKc9ZM984Cv7Bo50
x19cgoeb+UM5A6eJI+P6NBFdnvVcRm4p/N1BdtbLtRePZZ4XqdXuJKFYbICcojyd
Ydq2PSEy8VthLbu/zga9rLypHoL6kMMvA9KSZKBPqFXh906MI4kzajNRcAWOy2M0
uQyk0QqGbR4uVtXSCq1fM2lJsbx5W6yxm74taEZbhsyHTpEhNhc2uhZ7/77Xi3wi
FFK7OZYRcz5eKOcNoFUCnKoD40sqKro6aBLvtWFIUxc3fzPUVVu0NlKNie+El15H
SkQD45aY9S3aMB7pI1NuMEerssJVd/x7WKX36XKSis1QR6dwS/o4HM90blovAxsu
3WIPCNP6TfQdJSTOkarg4plvPLalleAneqmotSXGeW4HRwwgajkmL+uR9rMHLXm4
njZZYLfildoHe8m3mmvH1PPTB9YUTNfMVjGCDvfOib9HWTClghBw7anQQv91iM6R
rVYoZ74pdrzLOIOBgjomLQY6PCm5lrWAHhi2HWoCK8w2c0tq/WypZnc8ZpCD5BdB
TBiO29uYROpDmvCNY3/CfgfOtHubbQnfWSa5Gv0nP2RIDBGqKwpAWPPr5sX4oODa
be0S2xz9TFWt/G0q6XPpF1ysYKHdR1WQf0lMxhutIRWLS1ltd+7UHUpo2tMxPD8B
e6OFyMadMSXCvOW6UZ3Vvc0O8O/+qCxfOr1l1jqpMVQlmj2THzsBrMb6IKEhQRVp
5nS1LjmywZ1ba7t9Qku/glOtR0FYUnZWfjKA9J6uWUUBPuqhG/CxpJMvqmlgUEBT
tWj7z004FxUw9G/TjU4wMMpR5nLthFnzJQ8dM7zXeHSI+AbsubAnSF7gOij3/ygj
JXMhbPwCHwBVhNLjKch8dxdI9cs5FJy3YdJEoB9JLJY97oOBRqz9eZJAp+zB02Xd
nqBExFrZ6pDo6HlPTeiqsbok8bcuynRsIJjAom6zodoq66R5VG1HaJUJ/JCKX958
yEYZE4c7OZ72q9Gnw6dXoocigIzfbOxrHnJf9+zJ7QQceDt6sjiF+/5OC2BH6Y+J
JYY8S7yVVwGCB9RMw5ABwizbOA831XN7NHT3brKGkmJj4zDf2XcTGgwhcVDSZvJL
7kRPYMO75U/fKc+k+2CvkQb2V9lDQEK8WvFB6Zx2lLoWLf1Mfts8Qd+KiAQeLbFi
uHEscm11+rNQuwnZKO7AYohseKBwMlQocKhLDLq3H9SEXFYr4QcEhvaLH2f8kDU6
2Cwlh1NUyIExV3qEOL0YkHGhPa+qrlGCsRuRObMLVHE0Z0YapV9FX0fWuDms+nlN
tLTTvFykxtK+WH7MGRCgwBrX9AS5lpBQDX2/2p83QMAiLMV4AfopS1a3fnvBrGcE
O797Um8A2mi+s088lIW5E/+h0RC9p8NuM7OiGAcbeil2qm0TOM5xYMH3ePViYgbt
oLOhVRtd7lZzDxaTeRQGemKLxhdKOjfq1zfx9y1s2YkarQoBS1mLTFCAAgtvJw0N
Suj8vd1wotdNQ63Lo8ilAc48s0JZUDUw+/TBMAuc+L8DwxlMJw4UQMdkyPDqZhlV
ap8BkY9VLdU7Uj2D5QrVLP7UwsA8ma9yU8/C4Y1fki5GI9mEI5knfnVSYEzN1twM
0LWyxDLgQgpA5YOn5RLjhggU+WevS0D0aPn484B43pootCaGurarJY9TqeUx/1EJ
op9lsd2HGEtPpFk0zseELK+rRFtL7lrReAR4jBosvp9mjrtTLdONE5ox2tSPj1t8
xeFA7tnyypaEs5qlZghcHC3qz1xdHnbjpR4JDKE2F6y9rDv6KfC2YVuZpj3yveEr
fgsqPlmf7Sxh2U0lvydGTRV/gDjDyU2VzssYlOxdC9W6xdHOD/OwkXPytLP08GiI
j2yOKa0thV1A/Z5DJweMFpoEddtE1noQsw+9R3io9hI2E5VXULCYwpe01ZFvqy8C
WOsyfIugLIhUVnifgzhtkTklF6NNOEZpdEyROWdSmjzJ3ByREdIz1+Hc0pgVf+S3
qilUeMn8vlSxgczPnZ4VwlMCKbrw8X0fZXNruJ1/CKDcsos4JKz6qwpNJrRrat84
kSWQyVJteBdhm96/XNgK966/epBwDEowGgHHhXA9RiFyYtdPDr88vvPzPKnv/MED
/AiNSlmlWBdUe8GiPMnhJouITAGvRR0reuA2sG/r9h2ef01s2A3pDazdhb39f6WI
AOl443nP9fj0S0D0sK+udOVXciVW4fz89FrTGGQrzl7D0Xx6XgMS2f+Hg1+zZeRJ
Jd7Il63C1Hb4hb3tdyadC5UvZniGbjC1XSER4ygNghtZ9ny891F96kGMNoYcBS6S
ASanVRjL7HYVvsr18q+o8VwyHOIFKyUQsZIlIPZAI43NgdhEGojgQeiYoByHDWww
9dhLjOtH3HeRPF/Ll4Aibd583twwnq1M8sXZMigRFcI1JOGW57YpOyHai40s8UeQ
F3X3PdzHt1MHcG5CsuByM/ga4sGlvhBa3oaWEdW4mcD8JNGtIPW65y2KHh5dS6ZL
DVdqeVSmCDNKx7d1mooVTKtoJS9nFiI4N+OprrokZnp/MBLzm4lzsWLaBqJcEDzK
c0Q10wL001+CrHnx2L6yJCj4Z8caHAy+noMUgkTg3ES6uuQKTLoHOEP7LeXGYBKv
Fpzvf0jE/HUWYJ/9T+R7Y7ar4JMgYgFwnIMoB6bYsLHYrd6QLzGHFQ9oYAlnC+ZS
KppZ/wiZTcvXiFIk0aUe+ZXGUEL1lY3+P3+AC/QRxxP7KEm2VmkFKeqmzMgo6K92
Gotcvrzyt6At/97CsU/Yh4oLo9wKQuMrsRgpd6v5Fc9TzwRGdFedUhBZK6pl5XjO
Go7zUreROkAjjy/85YVaoRqpsNVCwgTcbgaJEOkP5p52ZPbkBoQmNtHKoAsvSaHA
g/gyHapPYFPcsnCRlx/ONr9iHxbhtcwRPAMa9fWJ4l16BQNviqcSbgQBoRThFg5U
uA4S7jlRdHi+NOIitR41yuKgdsER7xxhxODcoMCG5VzoEMmmVvCIHwTrBpxS4z2/
bpat/0p6NifTlPzc2IB6yzsRFYc1uchNlaXapNyjXk5Y2Xh5IseAUMhY7VuMxzdM
QElbsthWP1dwaqgxaLp6rldQDUZlXLeKP5tkngKBdUOanzzdFQN6gmTwGihVL8XA
C3HJz9suzUZjJim/DDb54mZJO7oLUwyze79MOdIc0MDURJfQJLm2A+FMTk0OxxQo
jHWhbNLSmOgGrHAkRAONQqlpxIZIUYq1YpipyDkGhvcvuzc7OVElSPuUVIh6SUrJ
SEz8a9ASPWuZvFtkjGXoRzY7/Z3xuhVoDK93v1djKIlOXM2GQ4S2i7rz6Sf0u1XO
WHGsJVaLompcGjq6KYDBjgFeYmqv2cckSojbWiazRj/vJeN3CmXa18LdFKjv0pNY
oSANdtS+5NVgtXma3NwbgZqMGl9bTRG4ZjxGiOI2Ny2bSrhilyqzwpdp2OOe003j
X3zCzWIO/nE5PhweMI1MnIB1UTQt7GfQkOG07BKop8YkyIMHF7vLZ/kcjEpOjLYS
jKTX0FzdTFyOm88Sdfnn7+bKYXaae9melbzdyYvZTMA+saTpTmpSemh90Qt2OSUc
zsWRQhsQA6bI9BKxgBBKS6CsFg2Tf7RgtE/3f1Hw0/YX6BjLhP7A1dXh9i+juGeh
C06FPTxp1sE+EgRMuRzeJ03lhhJPH51qgP05zN1qJbTOa0mhGQw6Fj42EKLUJOFM
JTn+NSkSzmMlqFKbayB4j6xmVX3kyCvnmKKLK7hazGWUjrhwLquaMRwvTbfOTsvi
sOfbK1e5SceVn1FbJGLEzg2ilBpYWiHZ3b+M0PEn25yS601ACw/Rzd9IN+EwiWP7
hEAlzAsQPm1Yu6rfrEwl6YmXhdQAWqZTDEt5H1dU6PNOt7x8Zbd+5CNIlg/BXEcb
ggwCdi+e8Q3z/IGqAglt4djq8AlgxahBgzNhJOlFj4EbP+WjdggxiNqnyIJlsjgj
fYAgzAL5BiL2RHUMuvjCB6beA1hVvC0QdZgc12ffqAeVJLPjAxdMHwPgW0nKGPf6
MYwGagjR8T7/EG4c+jDmn8cV3t0wtp+PgnKTBlHiwvq7VybjNzLYqRNawvPBh32S
sT9KZFD+5L6phkwgvGTwjgC7kpHsZyhLzVZ0MeLOkbVRiqa3hfROZOcdk2HMM6nF
J9Dvg/nlgrheYV6bJzeUEjAl1FvHpuDXDDB9a1+DdOB88tmVIiU8twwQ4y3NJZer
aIHhcB7mffwYNuzo14xZLamXPGADfnWpYUDyt7bOwSRbmUNV9e+jfuKPrrFcijo2
G/7yUSGdDByNEmKdCnugabm+Vg9LsF/jVEkHawCt5W3OJPJdVzdJ9PUPpn+EXVwt
P4NeoZeEwPhOh6cS8MuMdrCK+eT08AOZFN8yM73nOg6phK9vpq3yCjNgsOebbcn1
Rr/1kMvoCuaHQT1mymjGvyOO8SVWqDXydgRme+t0PaOoufLQT31EWoMlI9bazLsH
dihd0IHgTYJ65ZL5J6C96SXU5oh4+Bm6S7AfCg5i/K6mfIlrX/kAXIbA467hCsqC
Zef8KbBpJQ71UEW5kdu5C1OMod5QHSDp2Avw7H7Jvmv1zyV0CUNvNVQhKp1OHhbF
sA9UVLiEfvGSP0NRPxXmutd4Rph0zDEAtxzHIzy41c58jG8KHjkJp+cVExYzy8q8
BqkdC7CNF4/QMGfIXzx1B0FSDweQlAAN+T3YZY1BVd7+pR7rZJIt4tjRlMZwbuTl
JiBpoagdwdk84KmT7nKqWHZEQjfqmjboc8UAOf8xAgLH/yLNd7ZJ8TWRWh9qntqR
xb2JwfvSikwloKOPGWRpGA3k9wyY118dlNjII4g5KbI9YQINHHS/AmDcYMk2y64A
FzLr0qlgRhbVrkbj8SdXog/IcurcgbI9u0XcyiPLreJ5gvkqbUgbU56we8pZ0uWx
c/Mh6QzWmuiAtYkl6Z+Gm21nyHPo6Rp4W98PfiPK5c8G86BJvdROUMn51X0+gcQ6
CpFuhi3RmR76iJpCHbwJJu3ONBc3lXawW6qFC5174WhdnEPvyZc1P8TtPrL2QNko
ai7yWNf7O+SIPiJUHVx4UT1P2cs8EoXMwh4gfCu6IPosaGVwiturcITSiJSkkCl4
2TBoOWTEqe6Nt3A5SGHMXJ1k4VU5Ic0wEwQWh+8qpeTfPVlRCG7KU7Dr5wWCBFVM
sTpQhNTZNCehN+oDOnl14bnc6nYRqA88pk7tU8nePJBdZN6S9IEgBwiPM8Qqz7OO
wvv5dpTHIU6EAf1ZDj4DfNLfgGceFOCwOKGtTjYn4tPbirAljAuwYxRfaV/WdL6E
Fv80owzmi6qZ97x31N0iL0hqwDoS/ZGSsD6v8VRQJw3bzhSpHKue7JlHdZY4wWfF
Lo5KFktWGbB5I7g/HKTJ3NlX2kjZBYIISVTDfaYHpayxbafT6gPMdiAXbCc7Izml
NiipCb58gqFqj2CHpQL7wY3w+rVm3sfXMDWEXuqNoqiLULqongDD4OUfD+szuXPM
LPGxqFbgyY0ci/LbLxXTYM+6xrlaTnVMhbxue2+tfvSC/9epgYJy2evX0wPNMCD1
pAWE03rsdDt58yCGCUwLdveoJgSwQ2QTBGyfEfM+dbowU8us2dtZ4SgnxqUuL3Oj
OndnUClq6JmSEXZJoAEy6cCfSZR4DhbRUH6q90hfuxQcQtl4BOfmFnl7QA83g8t2
jWhUV2JA0cTfSce6m13Xsm4OVMBbTnmUgE+fA60HAdfihwH6jmB6EYCalkz5XONL
H3OUH3uUgcPMWC229AojWm8TXVYPR/ByJqUTSMq9cvyBht2Jd/JopNJqhIV3NQ/R
Xg2OhTyHLO9HxqAewYz4rb9hG8eeaNEvhnXb3XMUY59XmMrHXJjDWwkur33g98Sp
72SSeZGFI0aPM1g7AiEDoeUwIen2H5EByCd6mSULXETWAZAuRmnJJG7G9Mye2r52
0e9qNC0yv7KAFiyk6CLbIFQw5MW8LGlsQSmfSDOFWm3qOAJQvrCEY1WgXof3x4A3
D2vhEQTTRuPG2ieLT/rm7Eu6Jk8GcpPWZU0SFd9kHzT1xm21PxvtgbsUIfrNQIOa
57u45Ij/4AHEDo7G1KP0nFLnm1vVAvrUfN5IMUp9BHEziLWYzfpLY/ah3UXaXaai
zNV4JQv0z8Kh+bblpUNrAf+KWjGi8gk8aAM9MKHXzaSFMPHkpFkzyoce0lEBoDxI
RecfW7uxZoTsY7fNXZ/XMoD3wVhMqIC49Lh1jfF4tPzykWsnY7+RdqTTzSC7OMGA
8K9OECjOrIoDlCR3kFegNvz+zh9x9vzSs2+RSa49Sly89qNzL5z1dm0b/iljzJXb
TelWeTtycaSigKjs0hoPKGCQ6JaFv4KfhmLqNaOz8YjBJJNh9YwLBH3TrcQsXUM9
sRXQLELjHibs2+2KLDU6CHZLdE4nswGPt11rvpdz5kpZiQlhvdnYBQlIhXflPXmF
b3iOW2u31oNbzBL8GdTxCc2s5ilHiVjSnQaJiJoWA1C7t7CNTYgbrfLbAVmq2OdO
Udot6ZGocgIcNIhJ16Hvakz4wNOSn9zHJLqL2zUS36AMikgeDQXpbp0IRTPRpji7
Fp+a1ticpF34W972o8IxiXMWyKYMIjC/oA3qTtfPZbhCOwsx3AqYE5/kTmjTGJmM
5/Qy1tv5WUTBJrdtzMCbAL24R5sWev1kyz3zSIzBCsUJ+rS2wKrCfI6ACoB/aDTg
YrsdEd6/kLHo5rMnUn4EMmCXe/hqMwTDvaOwOtuTnUQ+kxK5wNJMfgPd4aivUdEf
JrozynyrhHOashFbv4cbkbotiVPN5koV4kNdzzjgOIjl2iY5OmWHsJiEcFq3l7/6
T6aZ+tzF4SrdgiFFTRy/3P1EBdsRbFPysiLgThAGuWHbJ1/fC/J82loJ77jJyvMQ
vvQAPrEnYJM3bwxPDv45fif5Ado7wofx3oIIkvDZjzaU5zLu9t6C4Snn5xVSe1n3
g1aebumzdtur0BLg03YkhKUC6VnfRGCkHbshkcF2JTrH1B/znioneI99S4YUp6ux
ASuPoqav8oWkboNtYsK66vDSpFUsqhgMUL9/xCMwiIPLKBpSO7Z/Oubh8HECDYMx
nIl0aAki9f3jZENydpVv/inuT8rcneMjEmkgkMtM2m7kxzqt2bXBlBhyluTB6Ax7
yd9Lh9e8rczl3w2kAm9fjN0I7FnqAQP20LhSxQzDeSTptCuacoGuzAxd4jKlYawF
cTliaYwLuwvvkDZMo/zUw+PZxNt9QT6qNKNNWu3l/fOQNmMgzCq5eRNAHRZIs4UU
f4oDQwRPoeMQENECSnXGwfq/ovQDN7CxMR2AARP82HkpclBcawmGkNtUzyPQvb6q
43vaASWqe/W/bGAwA5bmUsx7jNx7IwOzXR7L7a1OG/Z7g0f/D0JdpAD7WznamePJ
w9ZiowlXZaYGiyif3Gg8mwCxeAQhPmXkmH9rtM8E6PH17iemspA21EDOp5cKuDgJ
fv54Mtii/il/uU9S4KUZ5Oe4cKTzNk5TVce13TGwDlOQdtUNfrns0297EUGlhnN8
PM5qsf4M3pnCdXv6b3UHLA0nmCCdK46ofLGrrEkbBk6gVeRVeRvv4xESoofeM/Qn
jDmWmsJWqEjPSLlxOIfeF+7PK6cHYLjpu1kH3C5NzazY4aOfVnBKUZpStljU/9aR
6AalXnUtf59BF/BLUWnrIBmbqOkp6JRC76f/OJVWtpNht8sfldOjjY6VNbeLBSer
7RKmjFwjGhFo8zo3a9xzH8fdpmDb1GM7eh2GcFZJwENMmZGyvwrf20r5ddBhDiWa
ZUiHkgf1u0zDOauSf3mYYA5TJWnw9YlXbNxsfx+sHIxLq7vu1SafCdLvQfm68eDj
z2Kf47W1aqumAGS6Dh8h73O6KDkjh7aER9/Lt2QkpgxvKNuNg2ar9oI2VaG9O6nY
gkyyDrKHf5Tb7i6g1C/W3AjseuxqzxAfk+bysS9Az2RH1AODhlSez7k/JYHoUC5j
fo87C6aN+QXjGJS+vnkeV+3wQbU40huwkc0M/GsK86YeL3I0Llr60+Dau7BLp8yX
2L3O9mUGDo3t0tHbT77MuU1g+a+Xke7u4MltIhu5wsS1dmzc1dA6c3KeEWcrb3I6
UJ5curFrZuE/Ekf7mE+hut1VK7qNwMmyN4OsLk6fOyPcKSYFvvUjeZepfL7p0/Ee
YxK6OjWMHkHAuLLHPX0LC7v646BY0B+J8Le3uPPmb+iR9xhN/wazzWosIPbpToPL
7Xk8mawaLmBJlGzv0BgWpLHDIYFpMdK4ZCocpCk3ZPJ0VN0iS6L0fu/ASW7jhwAN
MOR0ozAjqf3no+iXUaCDmHUUasRLXD8e6EjmY3DXxeunMEkk+Bt6WIB+rwUeJgmj
yT1ejV6RG9Apdzlmq6wnexU4dwXVHqvLZ1m+SZl+XqjZEJ4F4w+ZYLQWuaG18oUZ
Mj/8R3BmMMWpMeu718f9oProTDJjTPCtQ/Z0f4GGtN1dbQLxN9uOoOjyoPgcKF/F
E2P+qNCshQEIbSrRZj1g/TL8M+5/8vVPfJZw0+i4z66JaSSHz5JhdPH4a1Mf0Heg
5xo5fGJ0gUKsgdeP1lS2Gya9X08uZAPKCL0wxOM4Pp8F9qFla+EpTRFKZmzUII0C
xSD1uiDdO6znYOVr1wtaRWfLjZLhcez5N2cfcLpfKnjM/AA0GBnJgY31ku5mSouc
DFn5WVwb9nSY6jJmEb+B69jfQPuzXlRL964iiG17KXIEGfpRuh7kqqiaFwM6n08g
iLWbREMgZNM8oDQZydDnSJiT+2KBX3LjLamD4UQMb9ileueh66chuCK5m2KlFWEU
XNyPRpRf6Qv65K1LbgYwTZD49PA5hSGf7hbeO4QVuXec7wtDL2jWdE/e4ydKw3dF
ZqGpLOQbuJAcSDBJtwTrowHsF5CgSOQhfyMjAletru0rjIsGF6IxdRLJIsvyufdP
AtpGuzDdEUGeEnLg6pHAghvwSbHnT5Rw0GlSpBfWEXyyJX/aBwnqMrY1HWzZF3lY
rEBddvFxOndLRdxDTYJvpRwo+RO/SLtUPgokKAqTruul1mspsqbfOUd/kdV/pDby
YTCCL3cFZGa7lNm4Oe7HOtFPTy1AED4+cqxmWB47UmQ6/U4LJoVlx6J8OPidsJKG
N11SDb0JTX6sKHcgq7vjGDMCzUaUy1ksJKtMhOmsBO+puqKkHRDe3Bx3UljRDurv
HRE6GTv/5pCDvcYK218lh3RmgIz6cZMhej/0U/vnL6QmiZGhP6LPNVyAwkRv7Mq3
Drx0XBj+t/9yBvraf98pFcThxz6j7DgqbrCnNnIjSU/Rn/5z/nuFxKET2DkWYWDy
jZd2nJZkncemhYxVg1uosOSdeD95vs8ouvuwZo1uP/DhwV047lPpWG1N6OYA7lq8
lQ8EcG1S0Up1uzMNh6BJvHtZyMfqFfUS+/y4C7wSJ34eitCIY6/BWJuc7sy6+HT0
bRQoegNocXRUEEM7jqM+rXq9xUCJTn1CP8esUEJF7lQenxg77QJDIH1S5DG6Bpfo
tSVUfeNKwKWIk384XqtwjGsATpUXkXidhZ5tbwPzDci48L0cceTCf7KJ2V/x6bjt
YZvALGStQOkc7YvNqSH4dtvTk1d9pxzvgZb6Ce0CFOrdd6FIrbmN+BAJNNt3o25j
K4xqhapYPP4RegzOk7X+JC1oPdvneXqJi7UC9s6ijwbB2rai8bRoOCljIZdkDpRk
OKMlzmMKehj03xJ0DTZ3AmxywkYQuNnapbNqIKVBECBvbhFI3reHOFq0GpPdO+WK
kYUoeWGpRszJtlI/nzn39TnX9AyJE2ncvCniuPgO84BhtzhWiY/PX7WpgAjNsrLg
NujbdFEAzE9TvfJ40zqa6+uA5FUxHCY2X/DSvXdtYdQS+KTWLKu6EX0FQD6xG1PU
2Ajb4oRB2JYQcEo4Tqm68fTitipDMgXqAWGtNTUsaydAetgZ9LunWniM14mHQckA
MhHY1fOptEAjqpGrWrUHBUWAe14chCvftLhuq3QsZtH3Ad27M9S+/3g+j4imtg/p
pVI8lpPKGraiO25DGYYmTfslgxTnguEL2mYoFGh22DuufQyi/yzpLes7PDDSB09+
+T8Wwgec9ubCL5Pmw/+lXjoGp/nqH1+5vhVunw0MQM12xpMxljfTxQnT2k2wTpJL
h9bBrF4qpdvTdQpu/DdfLGC1QHPQ6F/ftZgOdrZcobnwxy/Np23r955S7pafNJV8
ptZbuaxDxqi3rDlx7JHuwQgx5ARP9dYCIptK8SIS6e+yNAQjXoKXDDN/vhhp8w8H
NDcbrcH9uphITJdqDIlxR2Box/YnhZIFNptLTfgx3pcV5zj4/Qscp2iDWRWew0Bu
ZzsHo4gRwGTqW8SBaojwRZ3IqbsNIL9pZbAsbhZfVtPH5k4t3Ro3elJHFPM8JhxK
hdR8kgSX1lMoSbNGtpBntYVHL/vDVO5aeaOiN0YTN1l+vZXZGEWAJX/k3KkhemUp
MLeplzj+NA+b4ptXmPbhim2+BLGHIcGDZQANJnxL2meeReoUSRXUi+Qa2wG7l3/F
Na90RenpsaiDoA0MVJuQtScC4N44X0V2eUb4ldzGkvI0WgVL3ETHW4PKHDRIdWWi
+9gIdzy/emPtxjTNsnqQphIY1vk/VQup41BHOTuTBMBSD1fi8f46YS5mTMcTk5vp
GkLw03S8BA+dVB1KfbdX415pOKSYJEOcOSy4yL+SpbJmmEVhlZsmaaBybvJ2ioO2
TQYkJmb4KKvgngpged401zY/hcyatMXJHlZPERvlTnj/DZURaRmXuFe28utnspwO
yAcF0YkFpMNhphbCHaWi7gpEuywVRCigYe+4q2D4QhL6qWrcaa1XiOJ7duq0bBp7
gGBvgYOAfeQR3q6+tqUB+wKhqDKiMoL6Tve7QY0EGvdhrb9b/oro6+ALPnvLIejy
rJMfF1oH8tLSV26oM34BEi8nfe6NivwSQVeIIOeWpoA6PQqrrvYat47PGpXGOlo3
LFnDzVucNGMBtcAlJ4limZBWXbKMfSiyWsEKXk50c8TQXoJHcK4YFGX2MbI632Sl
m6zMYFPOte4/2yRGuHzSaiPzrvaZqQgfueXxySs16X90SfbMwqmJLaSklIjrtF+o
0BfhdKBbqpWHPAzDuxmXbejFuZG2Sfp5MyiXgL+VJAQ45VtVmgyjhj561qxAhsNZ
TF08EasazLFcyfyLZ9dAVwpPNnPJcM/zyKlidgrIh6YwZuWS5OSfL3BSuaOtRB6B
mvUuSIU6n7+OuG3AWb3EG+fdWMVhKmE6FvgYbqEGEIX2C2CAwDAG4zMeuIy13v0N
Rmdz/ryvOHGNbmWpEonpTj/Hi9MhuRzQRIDvDTvtcFGpZco00xM0K2uGZmWdQr+Y
oaOlZxUsDv2yXyiZewpx0lvSSEy8An8Mp6ZeAr6B2SeTj03/GCdb5zLZYWviDDZ6
hMO4C4P6R8HHCWIrSv6ScH9qGwlSLUSPdB43aSPnkbU669ZeSvQdNBdd2VRiMnjG
ptNO2hlAVTBaZMBmk06QS5qDNXOORqzoCzIvBDVvcb5cgqtNsDyrqhT2I1KE88Dk
olZmpNJV/Xp5Qu2vQMZVTOAZp7Cgrq98DWFGVsd7HEaUn9WmU7p02LfuNQmBWNia
A7lHR5vj3Zs4Wdk7fvz2ayNzmlLsaVktPvjgtibZlD7VkxBRhMJ+RCDC1XfceGQZ
BBw9Zx6YX4SugKH0J/h+s972TsvTzyasomI+tQB0WBm652Nl//fcRplXnLi//Lir
xSc/flFzNKnBHIBhP5vAORDUUNEHt5waFrsCMlFSQeOIIw5QdcmP7aw844ZP79Me
C983tEWatutnxS38z5tdaUmWVMXykmoNeF7fL7OtD1sg8RAN0fp9CeGas7DVReA2
nzsucvYPWsoduIFbonMKpf9QDmjQLRqAUXQz2lxMLHB4WVtDbjSgzfRbdTvRe4bJ
4G2DT72Ks+gojqfAGO/HXIQdLiNeOiq02N99ewEDQDORKn9K17tlndnvVkWrUuvD
1rM98xCI6NLKrnuSSn/wVg18wfAFzIthU/DMEUPcU16E8WNDr7CMdVl5/VjWuG0i
0IPi+SntQEZ/MOVsY3CyMCwYrcefefHfdrjKfByx0wlcZGtdhi0Wj7iSoGRLLMaf
rY6bp3IQL+FNO98e9rCgvJj14AqwXuH9l5TjagvaD6lxM5RZh2f2CnbR+amNPtil
iNmpu/JI9Ycjhz3CnGkZV7CqTdqOiOUQbCDjX3nZX33JAZlrMmJIkjDMgYWQA+4z
DeoOYms3qmDqNv+Bjd/de/bTBUAsxEJMyoj6LB9ynCQsuFoy5MStSB7eZSjbajsz
TS0UPt9VvOjnSA2Q9RTgv99VBV1wRnAl9HD413B306blLkWDbqELBGJJ7tfQXpW+
Yr84Q58PlCRxiwFInP5C1bUrRi8t9v2iwwuyzZqIH6atOjE7kUdcEi8LYitt3n+H
cQh3gGFe5CMTi8zh1n91qNmqxG6YE0t7scyaNrPJ0sKQpV56NqQR4eyDdcwsTjEs
ygftH9ZpByMtdgfqnqgY/O99HQl4egjMhMxeenbYunY4e3uOeFays92r7Y6n/i4l
zEYCk2od8YYLV3DgdRa6/WN6+IebyjpkbqUakbjEzPpnBYJmvE8LnfT6Q3vOEevQ
G5v7KeBFTLvuCTZYviSrmJBvq8EGM5ARuWBzjiK1kvdZBENoSKYPoYEG6bNUWNMz
g2NXkK55C8/ob5TjV3yrU5iuve954A/C0IEYHr2cvpiqMepA83zcVN2ya58PMKcM
sAKYZ5Z5iPcPAgUQV3SBwPYDGCyoO4ok8l/bmi8Rk9jjL0vnu/DrN+nHGSx3JJVm
7n3vNvUyqddGTyzdvnS1VZB1Mz+haq5G/x5bAofhMndG2LYgrquVJ8xWvyfkXWT8
XDrCr1R54oPTN0jlX+IhlWUjjHHXpuG/F7Ev+ZvY8rgBdenz/A8NB7juG0XwN/aa
a4wXPjd9OAeuUWpXNEWvSDr5aUAIB7EXlT13oPngD3s0LR/+D8yYanfku6rbcsgN
y3nTw83Q1l5UfBd5lIr0cHdHFys02UxCw1wYRW7Dd1ce5fAZGmSHEEWfZ0orGTOz
f0+lMLXP91/ZUnMaAWlJRkX0LE0F9ODdLAwKPxeoaVP3x3hVUv5R4IFCOFoqxrIn
Of6uwZf9nrF+E7vVx72n64kqKgj5J6xOSKj9RwcG8BqriGnaeFNNGpGfGm72WwyZ
0wAOCmSumFPLRxL0u0dUQbvBhZOTrwm7y7HUtily0Xeog+5E9Qs2kaw2j7ZaaTRq
h8rRSFeXtkFDJPBGqmclNCpIfPvwnoN948xMTTuhk6/t9K3xtpgLY4KeEZ5Hp/5H
xhbvHSJ6+2PoUtr5rpPEbinbbLGUS0GyrNuVKLQcujDubmdkN/t6G3W+MPGttzTU
wllWLWPEjrDXYxDX4tYxAGmC8DE5W3qSuBcQQ74wNaFMXsEWbDBXc5Pu7IGO+odh
fmUqOmOxuNkZRImQqP/7Pi2DBn+qMNTZoBKBuDmEVb0biCqmQubaS0Z6Utl3B0MG
Ya2koh4YmIrzoz8Nqr+apzHubFtMxX2CGtZdaOG4gMtUVrgfhYRjhsFC4L114Pu0
gKrpDuiYL5FqcSYccMOxU77JZrqTeZRCMkTCRhu94KmBiHqs4u1qCJDS/1hhOmrv
oQNHq/Nmc22Bpp6C09C688ikKtcpTeZKuLrqRUwWzDYP2/r0LAaCHIbpHD/T+KRU
B+EUxXZ7KIgf9u05hiDSbJErL2hr/oSBQMS1Dy979EZ3a3Ht4p0SRpxkgv+LHHW0
7VSgwlqxFyR79+tDgnSn5BPU58WcTJcbjr6LNrf+FKKL4McSZ060DDJqg7vrli7o
QrH1fLMv3k+L5S66zDj0Hon65GHS2EX++m4AFMKoF8Y+KPbteGZ5w6Mna8eafwAn
yGVCcDFoy+dR2c3VJNjdk7BdrEybtu910S4XHdJsK1ZwHT7p1vcwG9cqi5CpPfGS
5Id5rzfB/ttpK6qt85AouD/ltdeswKxyp8HeV8D1ac4NHvF8yZ6I4ZW8Nb3NFzqT
UmVibfn+eJgnXM9wPFwEUeybjA46IFKKcIHZek2wgNrrQiwcdPzu8ET16MTva2w6
XuLL5+roCJ5QIG9+43xP4/gnA6vv7tsNpBGuSr12eJsPACxZANQu90X2Ay1Bh6hC
20ncPjcQs3KH9aQp14CDKMORzgbrlaeDi3LX4qvwHw4xaGiAcB4BhaHqht4Hfg10
ISFelVbkAIxScMtnJy1VgQ1ismFuHaaiy8zGunkLL9G8OY16w+ZspmtVMrndVK4X
5kkYQZ/Q5xSveuLx9iSaOkwNUH0ovAByrJ7AQOMvwGypjauQVWKdayFYelZl14uI
Pd+uu2hofPB9/VPXfV6+JlYRPEPhOhjyAvlO2znduitvyIwiKaL3V05dAS4dL4xo
pcN+r1AwIE51u2mUjaDPGozdlyf6SsOsbLsGWs/2WLqKaK/LYNHnrySxdvAelW5j
60p3OWYYgFpuVHIBdvhhHpf0HZ1cHzKsx47Poh0OpoQAxEp7ek2LBa//Kzqsr6bW
UANDlh0q3lLo8IuM419KAGsm6MOhARru8b2+c3pICINWowZZ/hJ+VFKoAjwXNY/f
SHhVvakVWeE942mb8JTwDslHaZMOcGCF8wCFT2JJok3FMxN51qHUFVBA8Jkwivf8
LhkmgrZTh2epeToUEc056EfyuS7fxYdbTZv20GiaL2F6zdqvWQVzZUMrlXcJKZQs
ABDgdRASDfqlsdREBVqWHK8+YBBG2lqRO628x6eabTlrlSioVBrPqN77VlaKqFcc
iYvUlOpl8E6EjjqvurChL5qyxAQy7T0A6na1R2/+loumqv+Ngq4zeHKjP9WRoWtS
4156ajL5CsuuGvDxXJ0DgjfAxWORuubxz7Z5vpVuW0lJW8RTvHNOnqF8JChBxuju
aODBSzuiD4e1/hXdjZorcwi1wKphhezc1aNNXF5g6lsmkWrDF37SjaYeZ66exLht
0VLUBrMpBLFrxwwSRlO37jyaXiwnefL+g9Y5Hh+2fjdcAO60+Q7sfBFD2XcVcaSU
X8NHuEBElMCMFy/Mt9HWf24dS2dmCMMgrYOiT7s0C9G7VX69dAcY98FPDoGab9Xu
WX/HbNMzgidkWhQBDiVVSuzfVdT1ZZvLw1QdOxNf/oYpSX3p67q9iq7YCSyjtBHf
rnlBdqQvyPto2iBOqo7AA6wES5dYr/pLMKUnBL84Qjfu+23hPhRiVsCCDvohvG85
ZuA7WeaMlWiBFHM2dqAUVdRUQOqqOTr4NkN7q9L79Plk/mwInLH+E7qu8EBLG8ar
pxowQT/MF1vLiHR187lNjJimr6d9tjhITdxP6ILhbL779xRyuiNZvC+IkiVxVmdv
4N7tjK4HFBHGnlVcLfNwspfywPP3G1mVqH39j93fLr2JJHWYRojmmTijb33Am+Hd
X5C7S3cwCkwKJ0T994Nmn2h5XEu9uIEtT+Kd28kuYl6EDesCbGOQknim6Kl57tFK
XwOLenSoRnjerswbHN3086R7INGpfuwzTcoFVjW5gezvSQTTzB6s+W6q9oxJCOrI
MxbYajNk/vcqdA1NC5UjZTbgLOPqpqNOpeRHXrbTFIQn3YpTxoi35oS1SnuAw0K7
A0zkc7Uw2UD7HDg2dek/eMP+sXrXr7Cu0Z48uN3z/M8FDbqS5P1xfXhfqkyeDlbk
N3ygKwly0fg+GZcxWX24Qxe1C9p02CovOQLQhkIzFIHwtUW9MQHZTBX5m6l1OzGd
wXb0A2DZeDek6YZkXN6BJObA2FzxdesTBFbY34Wy6PVZNt0cU+oVQhA0iYCGoFI5
VzSHjsM7+kL80FN2B9LesL1wHkIpsdqHITFEFYl7iGh9TkdpyXO0CLQaFg1VKOSZ
FAvF7DUgAP09bPaOI+2L/C3vGu0Vombslz90rq5h7ZVWR9/bix7as1JhvdZDbZb7
HFc3IlqPud7DB+sk6UyIDBvyZLvUQYI/CaGUP5FZwJp6SQkNsrB+9Pq59pTD/3hF
rTH0JHeZ4L8t4SENXTzK8ntygkHrJSKA97D73O76WOa97Pl/AXVLBGx9DBEwLXId
7dxIlyUwBY38Oezbiy3iv3IgJQiHOhGtXpB/J3GHXiZs7zTtjVu7b54k1hTC1+t7
mlssmiTY7igqoWhoKSTKOvktyyjFRRMKsmXnYcn6eBgmnjiYXw6HVgS/0Wxy7wFA
ZRyB2zkNi22+q369iX7uOA9BjWtiOgJvrbIE4Vh5PSiRzcVPA1JASpbv6qfdCCKq
9ZYZo2J0w2dzAfO8ahkB1hdTlURp6bcLZq4YQVLyR2TEbU/lfKTNQI3PB6L4gXVp
K/SmDKqngJ42nX7Qed8aiOgnjRXiw2kwl+haQCkpvn/JFJNpggitQL6ZogBD52bf
tbeLCsUvGMmixnDt+JmM4diEqdb1Vcvf1BaDDDw9jdNwv/US/2ZOA2Scag4JAmzr
zfefvgVM8XCQxBE0fGGKy0Y0LEZ0DbWuXBBwKmlbv79HI5nBaKG33QSrpRoMdRL7
84Xe08R+OswWMH2h5z1B35dDuD+J5HmKckYoYMZ26ivC6Mk3ZwP5+ZygvmNgoSL9
PFiWewUl76QG9tVrKaxXSyRSouDJEBKT9nieykuzEoa+FXpmbkO1CtQP9YIRGOnM
3JKUeaOkE3Gm2Vvlb+ErM+oi2oClX29TNg9s/tjd1ggIcozfwUFvyPWwvf90vZrV
VP5LvPIInog7rG4OUWChJN1HyWcOXfPW/AHNR+IMUYOaxgnL2dD9w7Wqxj2gUEvJ
vjo9eBOgHdUqdl9r6EQBpsNWMkQcQKQPxY/HNGIetvJKFEugkTD3gr+8RunUofv9
6PZfiJcD1Ehr0+SCoQ3DCvJ3SaEx6qqUY5guaJY2QbNlwFsimC+prahTKj7rChTr
SLaCsy1AVq6OLfkwIezfl94/hcGRqNyXP22dOmw30uKkw4mscZUyIEztI+VRLMUU
VSqKzKvf6CzWcCbBNAXzT8n4AxxiyKMAU8rI7Vp86NQsTPAL94P8AcPbCV70ZnbC
RC0F8/UzJZsHysjDRMa+nBlSepaVuxW0jxuXuVbED3f92lYgBCT4/q152HS09udR
3E3zWZy8+FfpKl7h/iZbft7T+tjfUkI+IZG/eNCUJ1slkZHj1HerkCJer2d6rp3Q
KzIWclf/DEojZrMdt3d6J5arQ8JK904/AHiv1J38S3wCh1utnC0vF5rV2KK/G9ma
6LbNhkKmSsuv+1pOn0HBqe+ZZmo6Z2B5w/VLlPd387/QE0TwEojCvbUbQo6anWcb
SN4eJqC25dqP/k9ca/MWo41txfEoQv4F8v/ZuxzNgKP8MBMKuccEMusLVucu9D3e
XO3ISdTNa3kmaIRnf8YyAe8MTRLheAwWdtNE6thSw3ztjJEgAzkshlf7yudW5La+
fzgdGmSGm+A+4sjCRqvZlY1/8zqFjyVEbUX/R+2gNnQGyZm2EkdVZI6LFB0IXmLR
/jsh8HxcvCI9eRv8pBxiI4TZ9NiTHgYPYUyukMG8OF/u7Qy3bRD4SLvlrTUHmAfI
0dW2Q0Qc5Lu9YfAHwBHRiJRvcGL0x7ZAPk33nNhDLQAtCazvEyT4G7wXT84IXt4T
XvDkJf8B5c6okBclTtgBLqP10r35UWIXiHXZ5j9gZM+cghr845p6FlpyLJ/MWsh/
54sD5QXI2X+ZdHTrGGo3tHLuWyuieT6DjudeRH8sUCimxz0RC+aioJOr8LavDawB
G13bf3RjFK+zm/uKCNzBg1jbVw/lypozpLER4e6GgGc332GE1eGQUWjgs1u1x3Ms
3rpHONKqHwH7UkTJoHMmcbr0X7/kClS/r/9+yIS+oZfg7t0qQDiY8NogujjJOBIz
IeZ8gULnEK3JN567F87Z87Fnsvn1TVsGQ12hFC7dZ9cyoUlk2ZRLvtJEE/BM4L7g
/iAXzqJki/grMsaypXPpP5NbI/oLySQUtsyKpHeLCTxPnC4UcIRfsXs8K1DEUBS7
dJ9VzogPz9Q2CxHqYMs9de1wbFDY+zyLYSJGPL1/Hpb1o34zZliPTI5H/Biq688I
wiXdzBZVuCOAAmkL1awmDxlGlM6uy5r0yEgeE4U570OXqDHqXHC5/ZCrsfFDOS91
SbyyjuQMKTXBIBLowDFXWg35eNIZLNn4oF5WcOYudIpcEwzwSAjhArlFNCTmWFYC
iDuB1mOu81IMehXkWTSO39ObmraQUynpCL4YymUI5xSJsg1WxXp+dl3vLfSgU8JJ
hQcX7qLEDjTCZRw7d1ROSfkAOF/kXBt8BWCGFX/XuS7DmPnqq6aSd6wAO7JxgcdQ
rrNnerXxne8TS11Cl/mCwEqqRyeCeYvc6+02ZZhHI5tQ8LUWRUOHks2/Qfn2qIth
YV2TBenCfB2f/zE5Z5Ah8crhInj8X/yxEViTOtt+mTgYN07Du4YarsFUXUZ8Qq2S
yiyYFdZ3fwA+8CqZ66U0DBQTvPoghlQG1Yktv82kglz6CUu85BFiHcIM151b1qn5
62q1gug+qUczUZfDQv1wddKmcZ3ecfoArf2QUDoEiSuNoMk7uRMX/5GA6Awg4RBu
EHL39L1TZmdEb/3CGaeWN0bpFl64Q8KHwu9veVcEUWIPgcCfwhPGxa9ZKKkX7de0
TyQqp8oKGm9RuxmeaYk5adxxTU9lX9KDEAw0aqVNNtzU2f18cbrNagJovb2UDzQy
VONGKlloRWxqEg3iyK0DE7OrReKPNMz4hVMKgOMM1d4Krf3aydbKbuPPzmHt4p1+
cc+bSmdUb4y539jV1o9HE+kA6IV1XtxUJiT9pjMQ5dGh8Usjr0Hz/CC1+iMLIgQa
1METa5233wem881w2JiIlKA5Bf8CQKmeTAZG2B5/6dNlfg0eESw9YI0J1Uavt7Rs
Wmv3Hq1LnaqjzK1gTPLy/pSwHsAl3pJ5Ip2aK4F1n574VdyiNY9W2tdcLqpq3Hd+
aeugKxkLLBDa67tgdsp7jEEHyNWqMgYaSu9fdYUqj6aZ5xVoDkB7zeLcvC1Y6Fsw
o3CsJVFS4XvU6kRiGk/o3pSPLgIcbIeMsIqZ5aDVAJj55zB35PD02N0P9Y5QsWEk
kUw6qUrnwBGLTozJwPUsiGim4ppKd4NJ/95b/dM2yseS49iDWQJV99dd8vRflnb6
k8QmcW/cL9cukerrfxpW44I6Hd5E37NbvbZlse1E2tELvEoc88jZOptT5LT01JiO
bbxzxjtGAV69YPicBQtX1/42LIkWDOI5qVc8CxCRn2iSYPWQX+BmahS3g7Kjxqxk
uv/6zmnyZuqugPYJGjUTCVAnTa05+Bxnvwq3cO7ZqOjNAQl/jPzLwnx7TPvf6BNM
8bezjB7zz1WSuTJp7/YOqEl7hB8BqyguXlfVspJSMOuOy9oxiVVXPIIK4+kg+gGy
VTXcYT/OsvGhK58rQND8ISi05Lq74qw73ODeUzZkimfoNev+thyHKJC2+EAQIrXt
dD18LA8FRSvJnC3L8hKFHRd/XYbfyADCVRdLameZ4g3vR6fvujlRuuiOl3BH6HYI
pFalv7U9FcHYBDWcIAwzhIhDhxhOct7WnNEeL1bY66nB9HZ469wLE4Isc1/iy1+q
+bQNstGc1+A+OPURunqC18lhxU7Ydhw252m1kz55/88bO1/SjeuZBQAA8qrZhbB4
PxaWfGv9+YjfvzwYoVJmUhqhApCgG8+a50fxABUqwKRXoihH0GFYuNz+tw948EtK
vgSZyMxnsKUbR6NF9nYzlUHcB43f0XihTzzY+9mTE88Agf/d72T5EFIcUmt4iYyP
79eoPQXV4Zc88aFdMqO3St6qN1E7MTUZ5I/C5i6SEys9FkS9UTyQDvhwLbBLJFGz
ipOblDAD5pP04wdUgRXWo329H9Vfcc+e4szw6K4WT6A3h/BCqX2KRI7HqYq5SuhF
zX2LGW2XjPHBrFNkiS6nE20qo6yZxUy83syWZZqc128+Xpjljlzw0jgWfiOlgSLM
G4Slfcbgv+hixBGlVAED1HFgDNyYWh9wyHbduP2I9MJR8ETYTyFOP5iRQKhAaAlk
zq3xuy1qCpKQ2GiFobRMeGTu3vSGSZd1NVQOiPFEQpZm0XDoeB0UkulrVTUtLI+K
gfxxMBZSsv4oukQ8Cn4cugLHNyYxapuxUPwfc8ur3Mvu54a2XsqsfHkAYmVW3Asb
4x3P9xMbc49RLqldBokfvIoxihhaVwbdHUEzJHikmy71rRHcE6JeQ9hn0WScau2T
lz00Q/HSR5Y3DLW+ZiLvI4UTsumwHrY/9gRuqEJialt89JYKnKEyLeS6XRS8MuWp
K5mxA4AJxqwwNOoEqqTYlZdhjLJYbK0I+mroSF+3265htq8f6dE1HLXj7I/aBj6I
LB5E56zUA/KnYXrEk3oUwYUe3LEYacGD+WJFWVEWCxyemNWj3/SlJqn8I1kEkuRR
Sp1h4ImY64srut7rPxLu2faiI7QEmws40pb8rCDS3Npc9UMEyHnMoy4a21vjdeJj
/Um2b5YVp0hVjwbbOZmQW34gsQxXvG/BFK3awujsFNVqVINkGsLZMlRPtR/RvhCm
iVgW7I6BFZ64NhADVCQ7BkGm17x8GlWtQrEYaXNvQcPBMkB8J/7eh3TxquiXLCXY
WalpxYZwVCpxEssTs4Eoryu0E9wOcAFNtD2GyzMacknjaAYS/YZunCB0S8k8TlU1
oTv3NifJ9Atu8lsaF5FSQ0ANbkcvWJJ/8NtpWcHJWoY7OAPyYajdbtzwMtHbC/ye
OJCs5uCGzdIEyOUUV5b30O6w6Jy/6Wa+/1e0MyiOHCmlYEhfh42NC+u22lWjtS4V
WC5AmMGhmTvyujeE0ESrizE9GXMsxnsWFp0VHoabQkIG8YNu76TXsiPgeZcvdp9C
lUEHAKUnUvr5KTHs18gEMm7ZGylMSewGBLioBNv93cRRCUK7k3VlE++6+kSS50u5
8BU4tJvEnm5eNLh72YnTE+1e0Q/k1OkqusWPgheOwldmY3DY+OVSMmdN5TlhXFIL
tJGRWL+ZmMi/5NnrZLZLrF8XRK8ArfIVIdu7EfDdIN1ufxEf8wJbhqbe2lqmUthR
7SBA3IuCxamwK8W93fCsQF5/+2PG1gAZOhAXkq0SZv/4KcDaRajsaxEpGr+hDzIB
VPcu4dah4bvT+Xb+TWztqXnayHAG7P1271VeCbHiqRWHde3pM5UIq/dHFb8Ys5dx
n8SXy7UoQQlE72fUHFQFn/8JN+oH8SXbKvmfZchNU7UCsM3EFGr6BMqQyLsdbi1f
YAOt+TT2g0fYW/JPAhSxmdcMHEuxjADMM+N1WNXJGOcVZhG2rwf8fwecnIHelBgc
B1khAj8Ft0yKILhc8SwAxBzTd6NUlJcRexB6nmeJC/DmueYnErQCXdn76N6QHNZX
AgJBYKJEqCid06sYb5iYiEkF9IfpVwQR8jPvDMjy++t67NxPjO5pwi6ND0reVLQ4
/hYz/qJeYrozgKaA5O8bR6DSPrSdz8ks6mqsrhpJmImuksQG3yORsY+Q1nkbU104
cWW6wMEVRxmfXyycTo3qJLa2VEBWP1hKFOSOfImMtu/gqqB1VqJJUSZK1n/csUWJ
r8dPepxIL8iG5/UWDtvJNhyuq+Jm6gBjRiJM4OJTMTnYDCsGo8z/qJQwfais8tx9
jAjUFxg9ZjO/Q6V15KhtHK89CDhvILsomT1CpOH/bvT1GHp2Y/8cvWE9jbUS8Fd8
x407S9tqE7zZZ9EesDMFcSNtbPw3oZajOMj6FvSmdecBI/bP2tfg5um0XObBDy0C
RvkFT7msgWHvtytDqaEU2bLwrWMLHnFlsZv5tW5bjouxsh91Oxo1yVJsrs8/HOWC
4lGkxr/fHD4NvftsgtN6i92xrfbDliA5+0rn8QD35mI+SM/0Z3GtA3s9s1sFMsgc
a8P5KSrvU2g1h7/LtFoFCIzETLrpF+otvXbfoAqIWq+0UsXMyGRv21mL71NyOtRm
utY83GhY1rzTKrzbYseDbLH9u76ouYJvD9bFXzOXOgSbbZW1LUbLVRDjD94e6fgm
Ai/Q/AlWo+YzbJQjVjW7TdAszIxWF8vhTAVLpGjaDxP3cWpmOMER6k/Mhsw/vVfy
2IiY3KKXGmB5rnwbsFOIB2/1GhAa8Lhqg/KUVOBCQsGh4M5Vi4fFwO9T25j4vaei
1RnzhPU6z8GqLigls4ifEsuZdwgLYIrmw/lq+wZ/tPG1tcwzfE64mg+BuRX+myB8
+iB474y7BJ23s0eI73PJTACfQlNCug9qc3Wr9iMEH0ECoi0oaNICnWtGp3jh0JTG
3soCQnTNu9/vVUA1AvXtwr4OI15a1gjX+/VopOl3ul7Nqm5wwo8QrQ4FLbPnF+a0
o0uYpNryt92D4dJ5dqh6asyP0TfGXaStbBjD91j41aBu8XIzdSd1+vEDaUCaE42n
T869j/41VgXtFxz45782OGlfgzA81GDbT8d9/dzvA+EKnvoaMkGu+j9MXtGDtoWr
Kw5Sz52Nj5gsrTfRkXeZuiKvbqN/5F8ToWTOTWRw3JBXmkuvt1HQ4cvGGUNcZenZ
sc4BYvaRrNv9bH2XY6IpYqKE62DxduUukaZkD0qDR9DlxPjlTQlxHLtAYs4Tyop5
1rCeCIN5r4u1z8eTyQtnmKYcldoBflCued+shnemLxjY0bNhLgBSFAIGVz+I2woh
SNvWcdZG233A4lw2Q8IPtBtrSb2yoVJmx0FawHVaCPET3GrexJAjLy2uVusQ+pvF
izb2sGBz5QHQzDLSJy2/lscJIKcw6ayYSZmwAE3DrI7adW/f6okeDVxRCSXjTnaF
gtyFLFAganJwX266p5j8n9Ea9Kn8ZqOVNSZ21GXqyue3Uvi9eF999jXow+6n4UTq
mOm+eo1KaQKOMKdQTtiIuOVZHajPSYo7NMDK2T2hlYJ/2TzyfQl+He4lUimjS6SP
oz6M3NJlQ+TZnctIWDwlrvq6eUoN9m2bueRd4ytL3hZO3L0Pien/nk4IGDZmk6QX
Qwbnvp2CMfzzVbPPya4n+s0cvqGQ8LuRYdtoXt5Rqqi9S5LZdbA/G8vtdxfHq67Y
6wlGGcyWvmdCFLOihd3cyhono0+dcOOenss23BZmWDiJ9aO4cOVovla7lmqA9xhH
REfK90LpVEYYlFFB2Ou5mxVDjImxqicCkpiAOCC2RNlJQ7MM/jM8ZXMYdPjD0w/a
Ieo85OT+VR0ug03uifrJa6mMRSUqmDTdMrA07bkkn24HgBBa7/UPyRM6QTHqTngW
X/buFdWobECd00sOBnte+k82KCCtrcAbjZnTft31JI+LrW+cj7cXGtJAbFNcGL79
r6Fngo6YPQm1FyH8V7zPmnvujPf7/7UJyP4AnZBf7qN7/Mj0An1c9lUxgxo/WkNd
4S7MnYzX/jvCP8+huDOcV5Rb2S+qwnEG160gxulQwYOn8NdRxOAUnq8Z5Sxcs6os
W7ULbxO44D5JdxCCUzWhFoq0w8P2N7Sq8Jyr8Skopymhi418eXEZ7Z1pJmY1r1tv
Kxky8r2OhC5Yf564jgiy24IzPCDacWueqZlK5RDgosP/Xj5qh9Mil2DXKbKsSqhJ
zSesWGn1/VtxTuROTf5jhxbceAib4YYMgdHfbhdvOhRiL/h1FQMOar1kaaTZoQhP
0vRs+QQ1/WWoGW75Z7Vwc2A04N0K/0hhiEV7J3ffNoX0CAbqLz6SgSYF3feZ1LtK
CCtrWpKQfCNEf/Ex3Ovmax7qp7cXYkPme2ixOLBkKh5e8+1TE/AqqhMB5NlMnCuz
5zu3Ql1JwEjNFqSWtSqJ7bWvg81KK4At0faQZh/7DxI0PjRulLfS5knVNTC9GgrT
W6UdbGf1ANKrnFGRPgDraW8vymUbFAYZsSPSD16xXEjhKvNeglICxaSp0836eYnZ
/JVD14Dok7Tltng16hh4ts7wZ3PSqUneMUEJ64zI4IxZ4fTFwMJ+mGCQfpwO1V1T
2Th3SSXitNaFy4nRmjpgdJiKeZvnptcB/S0gNFmhlqEoCc2bnbs2UJIQ3LMdORW6
Au47mrOjcUVlr0M2k3/c4qaycW1JjS2uuhyTSyPGs9KMNno5Y/VkLohGMjBWquvp
g6gpNaHtdWIUYe3WzhWqvxERyqIwBM0/A2D7RlpM92fd4Z4fgHWyE+4HT0H8pC4y
93MN/JY+iZpg3D/5pq4NebWqF/DNF6JI3eMOrU5qeTn9dkzLk7PGWIf+TiXn47u8
XUZHEwlkSkQ3hx80+icXx6EWEA+AziMzt5lzzUk/aoDzQ1wtoaa1J23A2Ztgr6Qg
xPhBGKXRBFKl0LmP3XFHE4EhzQ/3CYjk49J9AXJjqEEBCXDUhwuJ6rqD33m2tuZ0
h6izpjrkLugzVDyqDDOwpDPEXT+b1CkAdEFReVkB7SPz8GAolPFPOdWYg76rk8Yz
EdlGQBDMNPr3wIigaOxdGTY2XUQO1TrFIaZ3z07YoZhriay2kCTTEsxVf1lwJdtk
1wn0eNO7i8aawUtR1Cse3zpZg+ITzoumfDToyGiDnKf0RPS6Sq59hrWl4WEMtB6g
OQkenINMQNZNaj84uEVfnNCqGuK8+2ih1jz0U2soWjaxSEGSq4TM/x7OFZpVD4iF
bhYm5BinoFojLe2bzBa3Soi8rKfhlDDIQUkwRLwP7w7uKxRLjf649URs0a0CEBVd
gya39C9A8AnfqwdagFbPHX+gsaxtk+qi3OMPvCbvsID5Su6ujus6m6nZmD1BQ+OB
NSrSyfNz5bjapwMaJgW1m4vAaeUuZJZWJaclNajphpHD88HjM4eGg9S1gKr50ZOu
SOHNDQxL8ZV/R5VhrHrofsmu9T0owCKA298bUy2SFbuM+CqWV6AgislG6+d7OIYw
KdyeBUHEdKtptcubmiKkYI0hU4CEeYi52FtCcXMuCt2Jl1w0dWf0fy/TvPCfDvVZ
D4w9n7vDahSghVE+b55V5w2pq/9L8ZFi7uB73E08hzgeTlkNaQeaKKj7+Z/nXXPU
7cHUoT7FkXBru9CCYsoli0eD88Bs6K4usBoUhDSj2viapSMLlS9T1CxHfyMcj0Dn
i0ty5R8YxT1bMwms20TiJIpqECKmHsbi8NfIO+sfVXO9f6UK7lKYRzC6TXCCaiXq
AZCEmDoEXCByoahmFvB7r4DjeJNV9BY08tXWJokHb9j2LtW9iYugbWPoyoPpTjaV
boXBXCB9reXtstALi4hb2ZRZH5HvHb/zEarX6+ylgf5IVCvcBBc4hIZKq/zwAIoh
ejqbEFBnoQVaS16WPvaE2umDNO0JGj+gDAqS8giYkOP4+8Q85iNv1U7E9hCc/egG
i+hoaxkScKP6xbnsBVCB6pLjYvawZbZVXMID8U06vR+J1XzGfGAOnqWy8A9r+bs+
CmlBlsvCWI1R16Idio19Ur67DN/DwjrjakQstn5gEWnf7OQr82tBQO/AJd+R9LPQ
nHbjxBruqTwq47zvbW1oOSKCa2nWJ8rsIaO26iLvcnZ8OjePcmV3Q3YArvD6NXXh
9gyQvqnFip4ExkAv6H3br93Dxb/TE8nSlwWogyxRE9mWm9ZJqcxU8PFTm24zyOiL
Yj6+SLIXr6Hmxp0t72ngAZD4JKqxrOm+IcUtyML8OLMfoqdMadDp7MoAQQlzv7Yl
d3maok3wxb4b6L6kz1Vk+mch02bsSXc9e2gtjBPjNp/VrSE95sZnmbcoGdR5RfLj
oTVEmXuOUU0bTMTOnWxOMQDe0nhD0ws9nb9FNlYtN6pGoo342F0kKkRIK4vT+ksP
iFEcEEJvn468AU6jLssbMRnF4bxj2x2ysn6aVcYy/LeeN7atazH090Hm6qb0DkKg
jxFohaI9MvX5dPzMyYlmsjaWiqVbSui8/QTj5bUvCkpZmvkhWjUxdd9NHnAlpapt
cOJz4eLMd99g+IrjDKPrGV+JYE8coRloCmjjPnwDSGUWbjxdk1RWoRSB+RTeY67Z
HNiHTChP7ECSftilRtlEPF0SHW1YnlB+3tzHDxBZkP0HXERRwMP0up1cxzGW7V7K
g3s/EH6reX7SCWV1QmHgse1D6o+ziMNxgr7Ont4eVx0oDxDHnG2UuCnJ92x/Elpm
giwp5cLDwZVcBqAqYGXOYitdiF9D8m7Ma8OqIAOqJfBPdwX+xv4stZxUx3ZcjVds
BzW5MEUwRHa+2HTqmNjN1OCpbWWX73u5YesGR9EEqRbsrxj3Z2gWepkwRGG+Xwft
cpkU50Ci9odlHNynGxApYYhkLpk41cOTdLPXJGFTh0z+24hH2qC95HLIhANvuOxz
qbEEVzECQ1M3Q4UfRqyai2w2zpTNILQYMNeZMtc/Ms1s6Ut6fDgkuVHvD/T2Yq5a
sQbD+4SCgDtrBNYbZOBRRqWxO+Hwc1ISY+YVS7LddPDZgCzVbGFwaALUJ2tUZH8U
FAyR8XqvH/g85bQ2DL3FyYFbxY4aZ5OkUV3mR7z0RbHGVloRt1RTGQgKTTRT8cGu
FShVBtr6x7mfTOD2TnlY0HXEvpWflmIkVBxduTLzJw8XYI0+d/M51bcMY8XiTQ85
LTS8a2TdS+3TxfQSG+uT0eXczlTitKJsxq33YR7c5r2tN0TCk8VGQbeBfxdyDncJ
+Jq9qGa0/4jmQCXdIj6DE8UNvpxFX16Br028uzMzXYaxsoBwlYWm1NNsr3BYgAlz
CO3DIM9KmCoAcKwKkX1/geaW5H4tXO4yTfFgB4NiLuGjpPZJtlfmSC/i0WZwZRqx
AJ9r6NcspQWiWE/vVF4Lui7zOJRKPKDGCZ9QVMQAtYJsx52xhU/lwUD8dr/jddif
REhhr9EWPqPH48rLpaULqLt3H7rVRHk3Bob6tZXxoAn18Fo1y+2+Ug/N/+klZDZ1
rsBu2BiiLrck+mYALMCMrI1+HC0LWykzmLPFHG+P4ka/0qNCavDejAZy+Jpe2JbR
74UKoMZpevi4k19t/9/WAgw/tNXsK1lTJ/+BnTFnLMOLAxubgtHSkehi0VTGJBMR
6GPL0MS16EyZc5MBy8hON4Q+YhPcdRJxmcO0j/e2pqw9TVW7JiDE+Den59LIzlfn
XG5z3dYzKbsHgS3DXQ4Q12mU4wrsQdgjMmfWFlUefTBvT4krCXAqqyPKVOAP7qeU
MFGkExfRg+jxGa+OLiDZ+6ar1dfoCBFguGRWts99uBPh6seLdIeTz26fiuQtkWTy
tbK9jdQfMoXbU8DO3dOx3l3SkRCyHkKh25/5d3fk0teaY/7jit3pWWvx2lUKxswE
cWWyJPhVnBwYWTsggUv9aBboB0nw70PMB5gHQLuLHYjjYfbbP2fK68FOKvurP2nV
h3zODN/tym8fCsxdpc4fGwNfs7OQUfP7YKrpgnxgKQxegzDV1ci9E/tRB1Kiy4LU
jxZskqeH8C3Z2c/be0UJU1Mz6MaIvjmQLk4tKoSqrSUQHiNPkdJYfgwCPHmTQ/E7
FKzdviDWi3WLq/voER20lnkH1douWLEN6vDiiz0GuiyTNr2hG0AsOxv/0B9q8//i
j+JWQ6AfMvtWxhu6IcNbd9nmR1ExrFHBBfKXCrP5RgDu8+PkSjuadcOq7x5x+wsi
s0Ur0YVgbvaVs34lyr/LIkuzFUfIgZf9jwNoTwjp6x6OXfMuziACNxz1Z3Qo5xOi
LGvz4w7Zuu/XynB0BVnH0cDj5Yggf0Q26tHjwEjPnBnVIIEWgy99czLShLeTWrFZ
Jirqjnv1WbQLd17VsdWTw7uCB6pS90sEyCjIj7bsJvWGYM3ac47o40LmXQ6RZHhm
2eyzYkMt3xzR+bdMR18oO8NvpWlMWxovqz3L8UmacNTy86B4SGHr9DU0IcT1qI9k
7nCW3OoHT0oJ9iAwI6/yWJFzfEdAlm6FYGVdpA8qNZAz5EdgujqaAZ0dPlxD8OHt
jNZF2sqdrkvPZ3hdToSpy7XGlnHnAXbMHdNNOpXjuBue362fKdY24BZmWlHR3eSx
2WLldl23PM/kw+GBNO1lYhq6lCZTCaS/nQoBBDEQ/GMFJsKhf8pJZtHuhAHKvzSL
zcVuCovCEP1RqKl6Q712Vmga9HpsHF7hjFrI+JC0JC2vYQvom2p4rn0O7RoNqaPR
Hrd4wu3R50G3bo8mhY0O5Wbv8IzPWgM2Qpy2/+JK53alRdt4EsxAGYmpz/yD3vYH
bwENELTXor/4qwFlHspICF+RAHYP6pgKjbJNNYcZWJRnUddl5A9oU6yilQnzAa4P
tcRuJquT484GjEc2wkoc22/sRfMNl4PIdOQp0jLmZUpP8Ueg8y/KjytOi0veI48C
F7t4NFbsxH9+WUbDapIoyeBOGvGzpnlpFIdbR+fUaDO+NAwRcVNuQ/ZwsHtBSRu7
SHUyrH/cqoBqTCWLN0MXbt7d6zisWPZnbABlxQ/+FIbhVXObjeyyvzl1bX29WGto
hFLeLVUff+xqZW+d2xZUVvKGIiiC3kNzcHVe3DP6j+rpTWqXMgxXku3KSOHYgD3+
CIdnIXWLlkbrfu9CppA9m8KJ9nBRG1p3y4k0ajc8KtK/WXlRk8/JgfZ8i+vjMxqb
gG3jfO3b9IMVZutQE+LzXXevI/AO/G3xRMbkMt+PWjvIpRC1X+njagzfqUce7+J2
RHTsEGugBnPFEbOepZPzheDp8BcELVg7AP4QC1D6EjD84P/wTfuvdNe7X9l0G1zb
2iXPWs0w7vuWBZCNSRkSAxw3BR0zHoLjjehdsEaN8h5JNT1H3L4TvmFF6/Urq12P
n2bH5qUppdJWs9lv7jx5MWrENoRwk0LGub6n68crcQKeJxTRMLzz/ZI7uFoXKuqa
vH4ylo8o57uKS4Mc5sSKMJlm6mMa+UKEYmWtUkYoeZjYd+DtnARNDIW+8D9HTg3J
+5PtgIQRkMBE76eXv9tGqt7wBRTLhXpSsrB3pbxGTNibBF241LVgCs+zxZ4gYSv4
5xIshPEYqyoPEN1x8yIthuhH6KBPoNGjK5ah84zlUDr+77deHOqpoCMs9obCkISA
FIX/lcU88Pp2a7qUWzd5Kv+/5gv9YFgGTA9qX9a21xmSydUyCdKfxvkoJxUA83sr
FxWc5gHh4mXgzSQ8NpTR+ez7yQrZsDEdPmsga+od5Q/cPTr6By/kX78BiG6en4Ek
2EQaAohDLFR9Cbr8ICAQ3znn6n43IzXZQbRN978+ByuqFL5DyfJ6NSRbwi35nXOr
jrFeMm5juTFY5X280F0AgHLv6ZJY1Sl/oOX/IeTYz58rh3VdtcU96nXto0d+JcvV
3UjD/b9+nSpoU+sh9bCjORnxM5qLJGvtMDmTFR4u9ke11O+/+DvslWN3wGdPZhgd
SdK0SKlc4G4C7qN5EHX6UHaq0aaHETQFDITSATT0Tcpi3qNGgHf2LpJC/i+bmbpn
LUbdcHHUlDTbmc6dPlqIbJRTeVKTb4qyP1XqF+xx8K9NE8zfKVJDPIkHk8s58YAW
La75a6s9xUKjeamGsLCxuc5wAsfB0npP754EKLIdjMcC+fPA1z+EfglWaz7hJ0H7
uuuhWwEK9qSZGFJRc7k4ui9HJRL8HMMSj1m2GcmPYpG9uIxVkyxKYogowEV8TKyi
d+vEelT1DWwH4azWuxJtxOJSOud5D3m8JvTFUR6XjbLz0TFKrBIfmB8h9QDgkuTG
IEN9acNU0f7IRq5fmFbRJZ1uyoNAkNaqD0GuovfHdpfkvbaJWEJ15w+9Y3EfNB5u
i7v5LVxzD/O7Ln/pYdMET0ya+7iJ9HBuk7iMPzTr6WXxbNIUasp0kN5nQwfL/9oV
8xQ/dnxibIWV3UvJmsBcapYn967YWzJF9hU/1eDO8wmiozjBTz1i0itLw/v7vOev
/M9fVGY+6S2LgePVVYLZV5NgxG/Ri4eiD4PIAcpZQPFbYaA5972yokvFmeuO4C/B
RqU380sYCTr04eLOBrQq7vh99d7RL3gIY/FyL+Ub5CwzV3r9bWlhb0mgNXbkJCH/
yVGRFWF+9lBmtxzo2eWCc02cCFtopYki47A1kUfPS9zvszZz2i4EKwb0fWbN99ho
+kwSTckhgYh5cQSGEnU7wJNYflcF8uA+BjWhiHShsLz+1WYb9eynaU8EYeL92dMN
ngrOh2n1U8ZxRKnXykLDub3Pzs5bWRLsi7lqFaxBzO4o8JQW/HKF8sJ0v8qpdjYg
IQ+KUvn2phNsX1WUzxrFaRPLcQ1OfLQzGbLjIekuPcslYkB+A+L3ZVIw8VoEz3K2
wOUK2BhhZaq8OCDIF029GoqY1mud5SVbFwUjMK3xFs/HNaRWyPApgqzV5MBEBiSv
JXgkZ1+QBfkRIf4ngfkocfNRqeh1lXRSH72J1QtLc7bP9S3vCeJLizge6gu5FJgC
nOAiMQG1N+alWjNlKue4e6nxy7JHcBbfR9hz+BY+C1/jUgAUFLWnKuzPY5P3ffLe
uvGgz7UtLrXeJcW/tI2+epzyIhEIAYyTOAlwS0WxOVHcMsah2YN9tjnDspmE1tlS
BTlAZiUhCaXYLWpihVree/NPTuGS2/owrEX9toO+q764Z/BD2TC8mkqv23Zx91Za
p5kbX89iDAfNhZrcbrbFxAQf3cz9R0AByEfEWzq6ItZmkALOmwpriX320q1aDdue
yah342YANuyj2haQK7zlFklxnJV5oeR0wrWzEvHct9RjAAK1jGBU4WMh0sKfLQS2
8eQ4i/koPreUJ4syZGhuNjN2tAsFGL/2EtWnj/K9MrzZ81GKmrfPsAjhYtl+tYEu
x+jVFM6b2PQSBsLfJcj7/rRAGl1e3G7yYflARR2+wqnvtc6ipJ7ZHfOzOYfXQVZU
E8REQHZt1OH6LXeoqkgSeej/e/fx1GcROK6xXa3WhyMxH0QbX1UzAGIFflCngYnl
3H1urSeYuQMaFz0D4RV3a5QeTHYY3Neav3aq69WX9A2iw2Zu/5Elvca/XuxfBDNg
2+Q+dk1vs2qR1/AmBXuXvAPyyUalTpySmngGruG4r50aL/ZpJQ6nou9k33pv+6Wr
TZ+fDEwp/tOFG/FwzVSq6hJ3yUarBfsTsEGS1QxrsytnAQmwpmgLOBikci8kD6JQ
CG2C+w4WEQaqMMK5lfGAWEu0vW8oq7Nvi6+qgvQZ8seLXVwUWsAWDIGqKEurpdvJ
U0eCqVi6FmHuE95plH/hsGUig9WEt76Hv81KLXNgLxWWyiUmrSANavlPTkoAJIay
CneUC8aPc4+E5iJGecJiv945z1Jy/FKidbQBBjWwHAgtMo9GmLBJBGE4UngPL6sz
v5dhY5Rf/7+jq7H6UQBScjFyYGpzwfLRyuirPGnID3ybULFIzagXRUgeD3OwjxGt
XAZDf9cYzlvaVmc9e3YcLHP9KDQviD9AUquc27H/7yDe4hntw+/l6kIu+k43E25k
w7K293xadbPeslib/KpUjCTPpxyRYivBvpPsieUdtVJm/QvcYa52AJspTGLTSsPi
7ekHiOL9OTA4pWY1ga2eokQFd558yHP6XBOj5jP9nSajf3VKLuWqhXMik6KKmOes
Cv8VtoeFQa/6f/fzMzQHT0o4SuwEG94ZUb64cas8/N1ayWrai+FsNRTNL/0ph+dm
qhsYJTUkTm+dC0HljbTLxhGKKswCRjY4f2LLiAT5qQKctibdgK0tnywfCsuTn0Gc
iMmMbEb5+13iADV7HABsGYFnn1iJ7QPPxDeyh61ZANWoraxm2EscTWfPRt3wDyaA
RVcJgNXkjRVdt6+FrescXjIaJAjek7qPGIvwNfhg31LRrE81Ezx/BH6PquPBCwLV
wP+TePm2cAjYSzA5eSGWq8UIrNChIng4OSRWAeubs4UeAImS2U1qytKG/5lU4MhE
zh3FmBnB01E12FY/C1K67BwM3vY0eKFnXVyyxi4lpDjYU8OXTnmJ0+t0a8kF/EzU
K6XDScUi6kc6SRQecdj71V95rvb0IEgDHZpquUns8m0XFdA+b58N09wmKO/bLnbT
vE4AYvJ8mCZUxhdoBpMW+7ezgpkYGaQWa1d8uyubjwlYlQxQ10dbLA3QYf2oHWzb
XmAWgcdHX0eM/Bb4ewypscugVGxD3wsXBgS5d+wTrwD+zXGb0Xz5++BPyAZhJ/ew
Lb2R4LkLVkZZAKNsKbq2jZPY2P0D2X8AueDvNTHHoFPRu2rhRkNPcc0qbZ3h3VJx
snecDC3DKepMzZeMo7ox4gJsGHwotdC3wJ2XyhbhTsej6kDW8UlZe82EYQBByGSu
riCiZNhr6WMhOqkaZu0KL23tmOKakZPQlMrwgR853LuQG7ZYAP5BybXAiPHFbzsS
5qW6maSsJ7GAVYr/JOAyC1Dat/p6lE83glHkOr9H55nMtk+J3ZYjRf1lKUXGVxsP
2KzdSj9EZV8VuYq13g8p56QlzQe2WYkZNqFnnNa006anYJDPVFXb70I3RsU7foxH
co7hjD86y/DjfaLrLvpQP6SD7lv9eqkMQ7w70pdsgO5dFQP1CXj9+xDNFJfvD0FX
FVFEgXhWXTFwQCLqvc/1cFbu9JyvGBhhSPK4wOcE4SdEeTLzGo6E2hCiMMKFWaCQ
dtMtHFH53Y7YtfRbk6aIbFlNviaZmn824AWMq/GL1ZKrFZ7jejg5nsJGFvpVI0YZ
L5CSPKvfgqGQojac82rtXpNinQg8EldzVjnQZVJHxh7RLy1pzGgfREdlgflBWCda
cVfx0aVOhOlPyGdIxQUo8cqyIQAKbwrNkRMrZwOWRyWCcrdnOwNAV0Lh2awD5Ikl
PXIgU0VOQXXkFKfDo0xOR7qMDooKK7Z2cUMppc7oip5Ji32c1X8l4yUw+njtrOF4
OOYn0iGJxffJBkxU23ce5fJFCkCgPc1nOIxFKzVgo9PedYmXnGX5mHp4/vMDvS7a
bh4A9f7oneu8pCmg97tDusXbYgq/QxiI8jiibYK7ZazYKb44/DaAA7hCueInsfcV
SJZvo3C8aRI02R6eFWDV0K68kDMtDiCoccx042kObglqk0RKmFFpzrqIBLsS75x9
KCKRLC7390Ot/HewXiycIOr0lD0KhyW4ezc8N3U3O+n8TuObqNx8joJ4MVICYy5I
LvGL7Curv5C51sNEo20sb4uida4Mn/uYFtSlR8pYL+FYURrL344way81cMoru6Ps
Ox1+q14/uMo3Dib2H3EzFwTaSJO1kHdVOkuSHsFwFThBQoTM3HzHxadNLMiJ/r/Q
70xgqwP8EWXzzhe1hQ41CQxdnfLyLXiLceIfh9pr2kMuX623TJHWXTXyfBy67fZ8
OYrNAmdw3trRnF6jYE7z+ZUN8fbNi1//FKjBxIf8ww+RmPqRrl7JSm52Um65R/pp
QmQw8CSiNlTy6ZWq2qiDtMT+J19JO4CP2/yhBEpHMKia8u+bnQ9cwU84FMGQQmRm
Jj3c7lNK53YR79g2goHFA1f6EpPFoAXL5EFIOHmnKq9Sy1hANiO+PYlLVdDHjvwx
e5z4zMPDj0GfuJFiiw5+Z7GoKlPt9GpE5L+61i34xkexMDyhHJJ5RRUknYkDUXHN
mTC9IQanGRL7nmvkGjV5sHVNujrKhzerEHiEuTlFnZZwnInVFmWjGFRp2WTRqje9
0eI8iX8CA/C1cUoQ1ykLP4oolgKytjOnv9inxNkTn0NzoPyMe4zDybvZHplf8KhC
nP+75qF2WeUBXEbYmB9bg4pu+GnQ262A6Sxc2xmj5VTPLsKHNZ30BgzqI4M4WKdk
janLhf/9RJvVT6XnOwCHHLqn8qkzx1jfUKbnEOoWWw3jtS0t3OvZyablBz8mS+PW
z0PC3OysciXKk0z7Urj1K+V0IH8PlenMZ0i7jbEQLAoXyenUNAgUuKN3F/ur5CvT
5Xg56lruPW4T3J//yHY9v9p6IBMx7XJP7zRHlXfe3wbKHDT90hF8VUUH11wGIXbe
TVNJNH/WqO/p8PY3QRZnTMbS1tnqPu8vepI0UWA1PRwZdBQhpnXddorzGtAhDVTv
EGSSyulB3Y0dnp/Spllt8PjA3sJJREsVW+d4YGoB9ijaeI2cvOtZrqESDXBZJr+0
ROixHUDc0d4oUz8YCpHLoV5FwyazXSUN/Mec32Yq8ZnU7qiad4THimihaGALj7aW
4+SKvsUskreqpsnlZTJY0knJAWN+BuhTmuBjZNpgYQhOdv9qWkB4RO60iU57zdwH
We3/I7CnH9n77Ox9DPC0ZgPzpEDWgsDtTRjFBEzopBsqoAQNuXQ8vQVvWJMahIvB
WHWraiB4vYl8/BAQOYWTxX/EJv0S9ijzRYrVouEzIN/bj7aruI21YvTcqksYLVIV
PWpI7QHwL+1MdYu+nF3TYCnwGu0ItshMXkGUK+Vs5z7zjB5Hz6fzTHeGmcnMSF+l
esKV6OhW8VfkcMCpvqPCVSMFsr5/2u3i9pqdAONbgekLdqFgcQC3lVc7v1+t0x1a
LXmhqLlPOgPjTPYtCqYfbNZNmaGowmJZXqe4Ajp5cNHp6JbgKZAVEF6VAoYA9x5M
2ei1TEXdsLmPBgtzgMAKkiCAxQhcD9AYXHIjxOBjdr4KLQC5w3qOp4k8/02pzE6P
jMeXaQl46jOo5r9FjP7f6pc3elU53z9lHmfgzDQx67erncrHkLVX0V0XGgj9K1wD
LskSpHLQ1xcEoG+3EUTRT9oHkjr5bnv70KOxVMv1db+JAqAa20Yu55vX51Dq39uM
RUqKgtFhhoWXfYBKnZY/VYf1gER7nhIaE6j2KmZV+IV1fok8e5wN7TNb0rDxoNIo
GpeNOx2lHWCRG8jSBnrY+mRLG3qxD1q+XKlpqsQUIVZLwKYvD1ABFx8K8Ygaev0G
bFooU+MystOCom/1pfXuiCON7ZJfiGwxDjQ7oecJOWtGph7gshdk72k3TWQMtxxA
KTs6vt9JJfap5mFppMFOhL/hPj5GQ34T3Y5gUrWNeWQpZruRHH1r1rQ1bZQSD9k/
UBeL4pR7QRAs7tzm3KYfuL0mBeO5yl2265vMpDiu/AjG+RI4M4hj9BYBeIwD6iMH
2m69K6+ZynQgImb99zoxkBweMUcV+NlQq9gjmbAojudfd+xxrZ0S7NMgWBFoX4l5
OXGKfXJwJMxpSwtMAs63kup3mKgDLAv4iavq/2jXF7mhBvtgtZCYWdunQLq6skVG
ZkR1ih897qBll4E2ynhaQ8WiYH8SHcksJSOFHmXMlZaM7G0ApTej5NbnL/vs6fvk
8ItjcJ6VLZ7aD0w8VzYj1hc59860qfVg2GCDlZ0/yfYJULwIojKpcJr7YyLIqUHn
DLGgYW16gAcHPNzyMhebGJRXqumq2JfzJt7x7QPzS9hF6pyTpmS3OvIb34j555Jn
llf6CpQk9BRVexxqcx1X14PbyuKdOJDOZQzmp2yAXSDjiXmL3jwaYbLX2qjZJqZ3
BNGM92fGCYiCAq8xckmSHWf6pBjpBeARuhYmQWSOglqb95dbbBVmVxwW9L70ZbgH
wx/S23dRR726kPSkbaeLDfqbatCXSi1q1thmkpCPzczyoJQ0JrOH/BGLdAJosKlp
HfY4wtz1Clv1yBVxW1PkW4/Ms7EXQU6ozWatQzfikkm0/78ktiIt+6Y2Y93pxwDw
BY4bF0lVnFJ8c7EdShRl+b4QWovirkZouOcAVTxe5OeuUD+FIDwdfekBd2MgAUtI
pFtVZdKLyK6XwCYKVaic2yZfXuhn+qRF4FacB3prCX9989MAsmEiQuTbB/2lrojr
ScpzIt/DVCEIxuuveTr5o8WL2cGvnXcjQI2QA/JjaZoZ3S94gbPWKZ/DpXhfrJ26
iTfT7Gn4NS3ZRBNl4P+iEZmcOf3aK0eLRoVdHkpkDUaTBkdP69hTbGNOpakSYieY
ThN/PnrCIhsJp9zbEry+DZo+cFwONhJPmfFX7CPXkDncfo5tJIt1BNYvu3V5fkxl
H6T7xYwX1WgilP3+qI0n0v4lZKn6S/ZoD5CPa2Bno2aq7W4bvHR/TXwyKc0Uexhi
zdvm9K5JJQp825OtWPmaguvFBnILj9CsG6P2W+1tQRWWAAD4p2GqCjPBf8Ob7nHv
QvqJ5WeHcdCls2QZGSz/EgcaUC/avjUyeHgFXaSN7GO6+skatdACZlKwUFXB878g
Dy5n41oMI4SBGHrOtnBFJaaANh45ACqSyCpe5fvQtMIW24XvwaxU0OxJDRnqZQS1
aHCSaQBJbM/AI74QpE/tcoi4YZ2KJ3MtvvJ5VgE5CDdbB9kwOkJtKEE5IAdB3icE
tEIxA1hDqkdYbnu1VUzO6TsTboE5vCEeVy+llGqrOe6MWAGkR8fnuNOwfEC7GVMA
6Si+cdP+FU3nehVgJwiC4awH+T3Hy3ecUUA/XFkXF5pE1oEh400r0MWGcFdy2vs5
bbtakh6xE2lWBJcN6NoC7gj/xfJpcHOrCSK/0jheJVJwTCBqgEmtrur2qjaOA21M
0PJjvOX2WzWlJE4iMGJkA/IgNly4jnO/xfFoMyqETfB0BvQbTESvaZ32F6qhN8OA
gF8aE0i3ln0507iO37E8Ks+D/xe/RINPefdPxRhafbk1+Yus7+aQ//kD0SsvRAou
qxq4c6IHk97v+LwfcNN6pOd2SSvjjoamf+ieIy2qtCy2CNMgJb5izX67IWSDm/VF
AkyC2Xx2b2YMUH/fAruBACtFZhqJdu96JcDatx2AG3P95G4xrJk2tzSAnrl+Y94t
5JrMOfn7JNZsa4lgAoX+X/ocRqXrsu4L3dgWPEq1TMWdVLOg0C+gET9dFBsnj1Rj
OUboPHHCwThZRLD2kWXW3jvVDlJ/9a7VC0MeSLScp4ZQ17/Mm5fVKd7TUyziCnOF
l5SDpNxVXX+SRGHtLNGREkwDBm5vqAxNIFt7EdTE+OHDwmGlXA4Yns/sixoiAgc8
vIo8ZtQKGsjf2RojJ0xUab+oxqw09jMFprEdFBr5BflLS3sIhtdAkcuXjDNtFm9A
t9OGdUuDy/FAntKKW5Zyz0XaF/xwE3X/F/huNvc541EIgq3c9i3JODJcLYF5VNXw
Vj1994eg5NdXd0mCNH7pUIySkMq+DHtmCedUSWCshLw0auO2qkI6XAqDnn/5nq23
BxfelIPBuCaEI/mJsZddgE48G9/MU+5plLiUasLnbDJ3SIFoyz929DXQYg3Kz11v
zfm7u61/uG2E5frE+eGUjNI7T6e2Lex4tLjPUmqwk+y7ARwJueSM2Vj5g9akeD6S
EkiuWzy+rIc0C+bzxyXus9suFnio9p3rxrQPZGFJyxvQw7rwegTK9IbF0jmrEhod
ryssMyNKrgZdmilvZVsBQyzEyHavA3hp36Bpy9PrhYJbbQm7ejboNAC6g//yaLRn
aGCPRC39jiAZ5lbrJeaOYdoMjgvIJQ32BRNFjrwAiUpxWq4Sork4zrqfsg2BoL9T
3GnPXkGyAh8JE7b+FL66iqDr+HHEsPGM731SqxusJBqV8aE7B4S4e7B1R8yIlqGT
ah+zRjbiZivwAG6eaJhMzdK3QXMu7gJXLzk9gBIr2QNZqg8BeaxybUWjPeEgk3gO
m2VxkpIdetsiuWhTklE36qxNj2OxkCOoAb3Co9kUwbpvnTk0XNDpD2sSd/vXp+8s
CKkkaprLvXV2y4MPdqRuFjHnQ+kdhvU8kKsDs48zL2VpIKaU7XSG1diVEqzSTfq8
G4eAVxXitFApeyxdDdjazK7vIN63BnPntw5afQ5Hm2BUC/qQ1P+5fklTJej4j8AR
UmBd487JlPme3sYsj1rEPc2kHp66pNgfL8CZvRlq1D5DWRKvQarhOtJw06wwvCYC
F2GH1M6+1rIhsv07SeswcXpOaQPJHSloYBwQPE2ooAzyIYSkwelCPqU8wrKMkbS6
2ZS4OBmGV272RetEjFnUhprPiHXFqB6flDvm0nWwcO4vJU0lFYGktOk1WJboHj9L
5/ZXEWJXfrESFgqjOHeKWmAxBiDXbAXaKYVEVoXKTuSLcBpAtj8uKQbcPgWE6TGm
mGLbH6eURXzUdHvhwFWn4U/s+HuLtbhVcRuh7MFH0Y3GEJQcxA4UjocMGKr/Xpj2
o8u+nj//q8sNr7W9Nx5qE57M/qWuV6QhzdMP2C8xsGqs4wmAlgjNd6RThB9tLbuK
O0OqXJNTYeN3vDbWNe+PGdreMKGZDzRwj2A1C3Qt+V/zVuKob6sPOPcfHHs6s8c5
INu6GDnnXew0NFy7Wit5wMIet+nZFr6EO+/MvzhahMeRqypW6W6P8zJU2EE160kd
DMyjRn4X8NOLd5FC0cYljQseGmoWsI7f69RLvQN3Qc8jiocnd8Ai/J9XZQwdTi/a
QvtilB0UaFDmELNrN4qEMZ5SYM4GFRMYcOgLmlzAZNK95RCi5r/VNdY9r2c7k9aA
OGUYI9BKdGxfvznliZ+5LkkvTZEXF94J6FKiKgdk13q5/HelzYom3EvED89Gt23W
JAgqzqZFSMBXBYS7I47grWHgobmB0aWl0WzvQ7NTXZRV6GOxaZFO/KRNijtZh1kU
ePvALYZL4OHErTp6YHw7TQGvKukGJ4aOxP0QRcEP21C5OMefTbUTupv+2VbO/phe
Hkd5eo1KQVtV8OzUmYGP4TbdpprRFs2T7XSR4kFgVIQjdOYqrO6P0eISkWxTYJxI
gnCCzuSw1z+Jv0flvACEQd/bXJ2LFkrXNb07AsZmQGwcIkC8zBllgdXR0nvf5+yn
U9P91DNzq1D6wmZOP5WHkUntfTZkeSJ6ljAw+F/2tHsA5q7tq1a/S0ClBR+q8P3L
pA8S8Pa/yRBb2bP0f+3W5hVJUnAi89W08rPjIdcyeBRUkigX0cusSeIp+T8HkuML
36o4kogMVqrByDOR2S2Y2t2UG2mDNERNMu/QrOy1awznTi+blgv9TkaglHIIbFvf
iyD8/VEMDm0CsFuK/RYSANW87ohHcU97RGcxd55y7uqJTK6xTCssJ68Nf7dxwhNa
3OtHbO2rIko848CtO71HwP+jIDK5WdBtlBPpF51pPl/LjWLiM6rfOucANcns7YkF
EbxMrr+Rx8HOKpUIJ5NMkeRumyGixA8+PITUvnf+aVuFZfw4YL9o0/mw0BbjZTWF
J3HJ0tnpYkNKF6hYNauzpEfLuvS3qIuD/er7V/Zm4XN8mUG5mUjKWEwatYrjBuml
YKGbA9Aek9EfAcRkGNKnkJEEJMFP5mW+zmfErddQysGn3kg0cWEn+66+lSnhA1UX
NdTlL6eEA/iWZI4x/Bn3yWdj4xymQyRVQQW675vix8Qcfk9J8DtCkPJ2V5TLMTpS
GTDk3rkYfXeiMmQMmpCe26ZYZUHeQO5JzBSkMxQ9xzTdZocilVXhVcdkB7jiv+WJ
KaVgYRXsZOWUikMJKhqS741+FOz2ZFGdKpAnblncDTpMtX6LTgsnS8xnwcvVhT/C
klTU9J2tr3JaUIRi1o1vQNY5jh4rXdReLhNtDYV8gdonM/EoUS4fG8gu1kGrTwyh
ce7v+fX8JsnSyx1GIePcQ5uQJpAXZNrHKmHlPZWeHfr0DI6RAPAyLEHKHDsPPdGX
GLF6NTCA5bNKxZTESNOtq+pywBvIdHmc8HXaZNV7PNBw8qk+sX58zV+unuO6SPmg
n8e9vo0nIwgHmhrng9Nq/FWaTPEadQFoLaO5s9uecB1lRstA1RuSEu2UlvN7Hl64
33xruywjqoi8XOU24m1+8f7nwgl1kejtKD4E1/jyFhiVWRPSHjapBHY6tG8125BS
MIEOei+QGgcNiSh67vCLNssFF8ePN1NzD/cTbRPW2Zefl4CajSsvtwSCF/sJqJBe
QhgW8vtjwPS+oM3NWMaCv77PUSD++V/PuBrZPHaLYp9zMCSj+t+GSI6pPJbIBXYH
u/TltywB+Z/oS89oTY6hGwiAMhaCNXUaKdboUEmJ9cXGw1OWcLbfeaSplIYngaOw
`pragma protect end_protected
