// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:39:14 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
acksTX4uRLctdL7LHqiF6YXvwnP+PyRFPhJjdhrv59qCfOctNwF7eNrQiniPTBFj
d0FWBcbaAqYzHJ5V/ID+Ss7Sp3TqMlyVbvRYYpJX8SPwv+eYZliGI3QRaqK16GA0
hkcFglcFifl7UCgBWIx+mSG/yAS0CbV/gwwmtLZPCrI=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 41344)
GhQMcneD4TclTlOoRxpheNm5qB+W84p4UaY6WSckGIEe4IbzGORV1GYcARSk0uC9
xOOIu/kCEmZ1/xMuv0/nnolayLjcZr/ldeBt2FBuMrCtrWKi6y3ISvQjlHMAVF+p
S0M3Y/KtJbmF7on6M+3AvQ1RvrlKcHUm0ibSVowjRjTq4yV4WkYQjoq2FYjG3KRo
5mwYp/VeB5dsRC13r86SeCfYDCaJKlwvfKXvhc+D4bhg/vvV3wsbRPSvP/3zsDFY
yI+imgZRfSpi0YXSLn6vl3DuKsCqHMaCmU4gHjdQQzdnoTDwFk1afVGeF5aKCJMb
Bqg9Drt2d0h2wLyvXthrJETMJzfGYmBFg5IJC4W1k+ztyxbGKTLXMf9p+iTJDTDa
YQvt2eU2nujTAWS3d0xFzoXs3T2uvDb5p9ZCxodZ5/vHS0fidJucXbbT2fI1XbhR
+eanfVEMfI19l4qZ562QBTaoNAfOifh72pvmENwvYh8uIExFTzIXJ8jOySJenC2U
75bvRyONiZSAEJHwPZCwfqC47S18F7hWGzYaxFzg1fBD8tFmhoHfGay04UT+NM3O
IWbiGn4lUKRt1V/VMq2pEr4FvzK/sqMAusU75tt/dXbea4eJ7aTxx2aCQyM26YDy
z10cEFvNWQJum4yw+t0n4oWLh6kdG3EONO9JNylJre7JUE8vrlc6JE4cX6JtkfNr
tmztwtQrBsprn6NcdiZKd8CFhJ3K44G51nnxCbWzHV7E9Dn3Rl3FtNCB255wNQZy
iXquWC8QGjv8RRU3IhJxVLIVEzAZyNFhl/FmAfIKwp4fzolxjhgGGQgnfQ4tOqmi
8LlQhRDEs6ofC/ncZZUdifMggmi7FZhqf5AILX8zEodJfvopY9QcCIVbs/xpw8Ly
PF+X4KwaW4TKvLGcTuNeJrpCT15ISAHOZq5Gi/fEAYyTyxWFWi6fznV4sXlLBmWL
g/c78/Qc2bkzvgsRC2a7XfSqRmZfhVgjyJZhuOzEV75vIop/iFcZInJl9QGIHh3K
kdWf2gFOVsB6OTEXxAKZV5f6xH6zLU7t4WNWDkvDMIKBrOhBAo4EV2W8SB8bQ1D1
OAfJdd/WF2QHaejlmIi6ph13ClIjmPja2/+lXKBO8Bf69EcbgVt+jI8+HspKY9cz
rpsp3qljpH0NKTpi6eD3Kcr6k8TXSgOASrgWm0+05EwI1r4GOeEUmRjixsdbfC5J
aYNv3o7yzDI8XVV8k2Q++aLthPXLlQAPVxdr5PhUMOchjvBvAjnDxZ+JW5vu4f69
ETjoI0rVxF7NwZHkVsDxp7COraUMRw9qQEDm/fjmWsBmV18hyVEKGCYOA5P9x63t
reFpjN1yJS2PG6p/bBzLk/4xpjLFhxcFI58RLVLaT4TuLaBldPlS5yDk4tUxaWFA
8wCGMY22M/7JcwXfbgB6IYJN7q12mnWxivIyDhUooxgibfv7vQ+ujgZ4SbiYP2Ic
58DCYI9H6JPkkzfLuqoyXVEDCGA1sUcq5zQcyE/SmXakcsq1Jaww33WxrKVamQhB
KL9JGr1CMz7l9U9eF3HFCKAuESwORbDQjxkB3cg+tUEaEXxSgSVC7sM3/TtMw5bH
ybQVGBasGLeA3htuBJWDU2cXi92q4TbZevSJ320WxRbLLIxX8905olx5CHRldZBM
l1IYAowJZwDEDm2ogT7Ch2s0cOhlwOOzXuOiLImgrdNtEWz2uHL8WN7SKuf3eJtC
cg2XEDLfsFQVz+Nb8+tBCF9/wATvzE7mYyLCN5q9HSXomesEtfcvqOZwGhUCbbaI
xhgFM1m8AgxC/CZuIwFZQnsMmZz1jhYbexv0EKanPJCTycbCTf5XpeFdleOFr/yJ
bYdkDkXZ+0d1r6bWPPdAXDqMecb6TKWL4SpY4+JM4mU91VqLMambnzfeLIIK1O3w
2yOFhcNFFueRkgdmAmsacGkeXQVLfVYeK7TpFZSj3v4MajKsFq4wtQNHWMJdvH6L
jXhXA4qGYia94ifQ6MaNmPdEOiG1pztA75+r+QgBUbdyOVNIQIWHS76Kb/uB0GsK
Z0P4GMK+63JYmmm4e2YP1wl1OgvnnkwfhqjFKh3nzR287IlNPxJ5k7ioHcTnO5fu
0++mfrMXA4cUbbknA39Kj1mRhLtJGfWVygeUbGxBL3oFvMehOFD2dt9gBAOC5L4h
9JH4mFtpQ2ucNmjZ29WOqC1OJlbpTtbPkwvhdnoue9woO4UmTnycR7qX23Oqd5/U
bM10vPHAzzxhf978EQQY9TyyJdrW3oa9QB6jauhemRUi5qgP9jlJ07GcvTw7HhiV
jtf9keh5FTVS0qU2UAU5daj0JhWVeDAk+TqaXYqlbG3+U3LO9Sf54R4kdkIh2OCq
4iDIyIWHiuAw00QSmdeSWx9lqebmmHiLEj4/gCAOKUzx0oL6BqmON5rbcMPYjBTp
cFYtI41fBx2CgrrY+h7vOU/GsIKX/XJKEZCRlfFO9zxq3rJf5RZMmQRocfdR1Yv0
7TOHLTFBxCTXTo8jujnZbS22UJpu+bPcTugh8lbVziIlo/CTL1q7o468juzT7zQ2
1pTq88VT8tpebsPk0GBOv4ybaAkmeoWY6OatMbTJoIY3ZB/UZwFAS4xjTf/GuEhu
V5oIQ4HPasCEUftuhGRbwFpO3tAicna3ov2ncexQT3XgaYvuxuvT8iUPPSjL5Ulq
D34vCESmMF2YnVcrvzHuWHndrv8rhRGLhOEAKZk7JEmr9AxP5mNv+txYAVVkvDZw
gfJy1U9ylysDVqo6p72XaPAwEaDGJf7SD+9FvGXzGTXatmp4ZKvvD7m0huHbAs3w
c18VsmhE9qVviwEgim1bBN+QbPJuwoSyT7Sfb33iRUKi25pYdGG+6N5pfkAhCKJF
iX+8oaIC3mDH2nh3wjD5s29PBFt2Y4I7eC/k04kxiEol3MVC1icXB92cah/B6fLz
TCSlSF24xx5FB6RPQn7eibCZQZVyjog/4fSpHZZVkowAzPib8AkP+0ES48jI8qN8
6/jzHYcabDDKUArUYc7VTq8hklk5xu0OLP8wc4vM2GksIcRynmJJ4PNpGWG9MP+N
semDsUxJwq77fksOnP8D0ru7QkGx5xzuTYCVJ0gIee/4a1c9Pc41vpgAK/c0vAq2
c9DSolGHl/fEp/GF70gRncp5LXyVWWg3751seQt0iq0WCZHpeuJbSdJg6LCBQYZk
oHbmdn2IaBXvR4VXupTneMV5jkYosN/IqHkW98syFcpo+mtAOj8T09b6/AtmhblZ
fvq4qLwYZE0mztBFbRZtxfzPTC2nBGDsRkAWpsCpzTacuxTx/WIlZ9k2GribY+kb
TzVRGM+vt2lH89EFW2wYok0PiOKYzfz/jQeOm/dqzZV5+xyRcl6WiUQsKRLDm/lh
1I8fdhraQYBAQZBRcwafYykpLPC24ruEUkeRfPE6D+MUN5+NWbZKZeOUEn66EpF6
DVluT6n+yL3AMuNbs2y4ejtSzooSQ/SCJaEYo3nNU50qU+kxyZ5TFV/J0ncTJu0E
EaEOZsidQgPAK1ORBuQ+BfE/mgIpNW/zJuWnQH78kJkl0kogSym92XsvtcwTXxYd
n2UNk90ZNWWoWe7bSHO8w3h5648uYR01LotqXSHsUvD53KQJ0oBV453tKd33E7Ci
bc18HrK5BNYkV01V4MTWcqvupVQ2oMessX+C5jI9DtTq9Mhr4RmD7V0/rMmJRqkK
+QKPMAgPDnLJvRaHcU11/f9DJHYPzCg7gD4LDvd4f+MyJwFWAdP8ZV5IzMlP06Qj
hcrC8Iny/57PM0I+ImUpyB9FpiIDY1YvLG9o/HX1G/bJzhiOB3DqDp6QGC3SQ6D1
Y8+GCQiHfDCEU2hQiL87e4DKXT1RPeWXkT2rekjN9+xU9In5gjJprG4fXqufHxiH
5kiLbDX2ZEVxRmoKWEXi+QbGgBwZFBBhim55Enny4iLQQ+nvDN+4LiEpq6449SNd
pDqd6mk+HSF8KpGj7lzQod7l61g4c6CPmOiWmwdbXCKkR/BIwFWUGzcgqfDpzcLS
rrfy9rA1eAyP1HCsy1RM+gBKHly2yRgB/JKxXZYxOrQnK8ZfJ8nocpBZCjQyFZTS
WbSeDMF4NUNUnPWUv+c9+kBX3amXqqPL0wskNXTDL7C2lRDQ0aNHvwH0nC1K4Zx3
7my2zFEHrCTbX5UwIvsg8mXkRdnM/Ro4aIRbECE6YLzqMkDfqR6ouhgB1oJ6SP2O
90iA4kVN9noRAGBT2Xe+MO93m1Aj42Q+35PpmPBzOoKdNsco/xq2/7WfNnDh+/hE
TBwMN6WKptk3SMXrO3g0bHTBJrzrveBBG9kBzpbn9+7WVWbG4irV+HqPmxZEa/m6
z61bje2Ht0qQs79VRInprhfufNvyPcEJF2v1IsbF+01DtVYmcFTmIsJAiH3K0xHR
R7GsQQykwHeEuSf9Up2oYZHEzdisGCkwNuo5scWe3kpcnwVfqpgDH2eWMjRBBFXU
EiJ+/aGcS/QmBWIY8CBgkCUKR8jbeMn6SLI3MpA4CkFt2FhzIznBQAYWqTacwyY0
XDxh2PLUFmGevB5pQE90lsD0Ty49T2YxY+3kbiYBXL0ik1/xRMX2LcDqS9T24Mi7
x1To5s0Yd9oI6PlYNYktfS+d+jB2q/I9WZE6LklQ+Meu6z6/AhO3p3LjuF6kxXfI
zWkHQvLL1Z6rDSdx8llFBkwcToZXdXxyzLjKxXpZ+16FJ+BiZHCBBpJ8h0qCzPZd
tse50/wphp1oL3H+yd1kgsQ8cE+DYE3VN7XJ6A/WjC2nI0ojLc/ByqzMtIo4a1QZ
tqbETua/4GPadh4YxtGq2KLe363u7QBwNAiJkHJ1PcW3oHaHbaG+OVrnp8cdU3S+
P52tXcS15q9CTuDt6GKqfvgvQLvvvNcrecjHfVclcOun5+AaYMlBQtbVZXPjsfjC
BuxjwGc53gLwHzqd7QZDg8iKOQfzBkNnemt27xvEWcTxmfUAocfZOT0c5yRT+sWD
zRil3bZONMn4gU4NCdwoT0BrCZTnJIPRg5hHOke0Wzo1Cbg+d9TEe5aDSoAIRjwu
3nwOtNNVmGp7zytxTp5lp5lDYNfn8WTa5Yd5p8OJztPLk+vLjR34Y/mDi4eZ4hh0
mo07f1ErzepXklSG81Rl6y3TbHm2UdjEjV9ZaKSylJIMVI6TwTFuA1wCRUslRjCU
4IDvPmmfDE1PphICIFCm95AerqplFWlqncGVqi5UWunvIyYjtlh3qgeIs/pk4wKa
illXMWyqANgZrE7DV6nN7CypJnOSEXr3GYJZ3ncAlqnA7tPoO1Py4GIr/yn403s4
jrTAUDX5KGDU5T+M7Yx02AEkBexHxH+g3SnpUY2G+IS/pao1Pqf6vk6bnQADMtrt
QJjRTEdz6kNCpcg57HP3wI4QKRpibwgUtlrH2yLMQKrstRcBGjYp2qn4M2GC0epq
ettFtIUN+ZnHkpzyI75PMe4W/OY2CY6yHOlnTS+tesKjkdPgG/4eEesVxHeUQFQx
rkWZVqekkrcxcLzeeJaK+s+Z9nOMHRcNUC4rdv5lL0RKIooKsqceW+xfd20ngSr3
22cAGHRVrmn8qj0hoWwDTiPmKcMpGo0IzTQshEd4Qkj9XWju2iCCQtgryU1p2i2b
jPcjyMtb2hFF54Z2udhH423tRfOPtpD4PKmhaUAyIu4JMO7UmSbDpGed5A65zAPf
6h/hRJ/ONfJES+EjaS6MJ9Q3i7Ar2KrTfVQxgHIqx4pt9QS7DHoLXq06IWokA+3E
BEged3PlCmFMulqJFSvpenY2klJg7QxGrGzRZRZmgylNqaVQomMaM/DNrWxP3LnV
k9VXEg/HyJPqAzwDPR83h1dxaFAWaEhxWb3Lnd2mrs7aouG5d/CTOfabI1eUv/Df
HyonJzMN7Kjq3f2tMfMawEgE4iFbDSSqgjU2u280tk087CtsPFfoV4p4nzh1H3Nj
HWITBByfElYSjfMQyU1d6v67aLAJmiSIZqcQBIE5Tf04oeH2M374ql4Xrk6sHPE7
KWL3SnRN4RXta/KyTFIK2PuKD+X+I7o42+W3bMV1IatkY2k3LsrLl0CyUvcZ0mAv
CKDwyIM+ts52kc2x7AzlUrD7xMJrrVNmX0mI6Z/lNiuGiOlRjwMuCQUgA+VQteez
CFwzu5O4T3UakYMYVRZOHXFpfgdDzyb182WB2ssGfKO9fN2JbtQaL50cnL/NV4JX
qLrlJhJ6f5/ocRK6QPZgqgMlmODkKDwlocKb5xRqsiY1P/vXFpgsH/cIp6s4Bah1
VWR03RQTal5edP4NeMFhplcfyDdQucKjf9gpZ7EOhHkpIYFF+PZJDpDkzPAOmoLa
TTQpPish+KwFwkZRFBs/B/W1McZs3iOql46bewdA3OZl4Osxvf0ehUQn9ed1gGb8
jd67eJ8FzAwiM8CTduDDT15WsPkE5kp+CKTOEtXHTYArsTdA9+YecdGEkd9Sq2lt
7m9lGtzd7DMtPvbZPfKXcVOriK56gJCHPS3JDW0N/03r2Owm5wLI7kpbMmxkYkmR
s2znqZmvhkz5NaL/6+sDwOjFxn2sXmprVsRU7rgvdhJBZxFGrjitr52tFuF5rr/f
tZX0SRodXzuunx4LuY1x9hNE0C1I47Sg+j3HcRulo89dRDPdCqwva87TUG/Uej+e
dRXOAlqrTcjsbFj71zWy8fSTzz01Ic8pazHo2V+8fsACNO/M48hAtLcZx3FmFBv3
8jz3LM/KG4gBV0XMlgzzEJWxt0a8v40tL4qWXFeLs8P245rwf6n4z/2hXDefOaYc
WjPTr0SURatDYf5n2jTwqZG4hfHOfXbRCwOOF59c6gQTk9yocHvN+GHW4DgiNmHI
HmQHrGfo6wNUqKSPQ7/lhwzsZJYmrnGS5TxU2m69fqqc0Y0IPtxU7UrReylq0SY/
r11XGMc8U+CAN8dPenxZXF63UlumWavF9tArkLeKSesvS1Cqkk301Gz17Y4+4vhZ
LdiF6cNBV2gy6fOa6IRHLi22nbRyduIjqD5fj2drJVV2G4xeTSVuRfAu6SbtyBZV
yxwk5pjYQ1hF+8WJPMdepNWP0qWa/yqKhKfLn6bRS4z4+3O5pT0jox2C+nppMZjo
+JSXxZDrqffmpfTDN+iP/mGmxzEOX2HeUE4/iR+XVt73cyWjn8Ef7TiQX6rsO51N
dpJNdues1t0pzlT7q/iVfjtsCJwKLwI9CtcJXbLqGGzU7AkL5ju0PkHtH/TrDWgG
v8tZSPyWQhrXfvgZpuV2qH7Er5sqfwjZflFZhhD+FCCBBYoqwKcId1uZk3cLD1lw
+tIblCdeWN0Rilmou7Xi7NtWXkYB90Ftlx/aWh4NpreCo0nEEnaCC3MUdp5NQf2B
pD4JEGGglU+RnLXI2XNHUtSvlrJvED3k3pEZs4Go1GN7u2PsYhs9VWrZqKRHAFd9
YR1G/knHSaflOcYJ1maDPoAon9GTDv9vzk3SwNeUTSKRstnMbFKq8wdAbCedSrb6
Tcz2doxxZpNWFk5JkHK2qB7wOMsFgsFuR7CtYFB9aShHNtrcyNLsj6RfXV+u/X5E
iw0a5a2JQyu9Pi/pOFb3uI7IcE0UjC68iPdQE6+YBHTdqFLHd81qS2lOaSYvBHbF
eQLn4Z4kwHdskifqA/Rxsh6Fan7Fzn+8h3LBR35gxCMlH0m/XnqNJP2V+hQZMp7k
1uRteHixk06nVwV3Y/8WZuahSvj8QZValTb1hP7CqfpFhNpMl7trxG6PSti9cdY7
KBC3yTMVMpUSheUipChPYFgPw0C+t0KfLGDkv0uMSbDkkw4NZSSJD74jsUY1khb4
v6Gqot2RCaP8fZSfip2KBBjtyA7CRbsc8JejYwh3c9qdOCWmg6RmvoekIX0SUcoE
q7lY1wOQWPb6WVa2FpScOUvbX7/n80vASyYO2doe2AmXwcHks4skZcQF5NMAiFSv
99htRgm9ZNYEx26M58oyXXe1j5l7cFa/dmC5GcoqR4x/BdgDq4gWKHaBGujZIKNp
hSBJml5kusKyz+yLLbQo7O6DrV+UwQelp35EP98d7xx4T1FxdOqc6xsooW6isCWJ
pXA87aa42mnRNAuCKCm96eDtLNyCMBhQi+EJ7RXakDAsBvpqi1wRGxD6DOkdkNyI
uSV7+jOrojc/6c9n+NRxu9nhchx0F8i8YsdqF7uANke3CgFN34euTCh/H5fASwxF
uCTnMF63wyaRNKwItFIviwIs9JBCxCEy45XpGsjeGNlyuRRSt3Ngbu/tSUAYasmQ
Z0kazqSf0b3/7kcMBO4A3vC9ckbx1+3pdVGRtISY7Js7LH1jlMIuh/oCKF67dmRS
DDE8oAoAKhYIj61SIEsXJp69ypUG1/WNlax6OfipZZ4u3PDLWFV1e6jxAJrsOVbX
xF4veEllISiFffnMATLxZ9cn7BC/mja1Mg0sMMfyzJxBXOyUhALw9kARpGeHngZl
Etq/ILuAQWNQnn+La3xPvYe7cJc3oJnQGN0iS8TTH3vKM6H6cGrVjkXBypasDto5
5JjPt/UqgCHgIiJYX4Oi+ZtNvVaoPJNAF52Na9aJsdsgx9Ok7eQDPtCuJj3xR7y6
10O8xOurNr0ho14S3N83caotkE2IMnrJ7DlHmq9PTppc6OcntFIx1x69psJfEUnO
zIarIWCaPyoHafSKX/RNu44tSt19N1AnQx+5moYXxC5i3yofXN/oum0rSB1qo8Wq
NPB8utHqermfhPiNhFCtefhO7OIApO5Wn7hBvepWdHP39RXVJoQrikad32EjvO+o
DnqdFv2nV+gJyFRNRmrvVgaH5+FMVVJZukQ/g/CgafTcPb3pegvA58N/dgJM8Jf1
j1I4Flif8CcvhnDqylvGuJ5qInAkANZyTd/1f2dBiwXixxaB6rO+LzMwEspoNupP
jq//4uvDVu9hei1HFoqioO3aeKwFyivlwAk4RnsqG5GMHrV7Cge4cRsgNguhbc+f
JewiOxEhM4sFEFDDtQpahoKJoVR/t26a8+V6ClrcbsFMSqd4o1tLtbywoPhnRtoe
qdPtoF+ilqHj5AglIPBMH4hF/2iq4RCOTn1RKDHeKkxWBCOhd36CtysFtCTBr1gr
hCg9B6Gb3QoT2YHqjqumdGCnjTD2W2j1QUVT6aNxP2BKe9Rb4C68kz/TeaHkFDpR
F4plBf7ihWp/++y+xJXlD+1kTHc9zguVsJr92ra4Jfxk3ZfPaejdXxCokB6OGINe
D+4ralM5ZI7NGTF6BM0hC613bfzyNZbdNvDPgR/vW8Tb/5Yb/0vQYQMPTmCwhABl
hu1zsYwyTU4MVBaYQJxlylrWb436IVJDt7B9dfHgpHc10nupyt7FlDJ3VRaZbQsO
5t8D+hXK11gDMZ3/y+OJzt3Oi/seTAAh845fnGlgkYKk2y+ZuXaOV6KJYeHxAm6r
2hafH3o/CrwFmt/suSCaYT+jy4bP7rwaEL9C0FdabxRo0xkdlaRWyUQiy9Z9tWJw
0vRsUZ7smpgKeJ9eI1qoFheYrmG2pziu4ih/spZdcCRnD5IJDxM2d7yHX3hp++eM
TZicMCot5i0QgttdHWEkoaQobOuUt8zlDhXAtzMpvbkI090+13ENVUHTsnSJV3Yu
1MjA4PeaRBOC990udF6WZC+lWnejk6pxQkF86bbxDU44fp69QsooU2cRcShYRW9r
CKWJ3xXKxqk0xJ4EwmZYJsWM7Y9n8JmBYO5MuKkTbV1mXi7kboV7/SkC0pXJyhEG
zfpImKVX6wB/v9fAVaWLktNFFavO3nBEUP3IVj5tMEOtfpw6uOUE6WPqfINX0QO8
rJYW6KWfAy5E2wWzskVlBIWAVyMTGb4l81/hQVXc1NUE7FA3/fA2r3VuAmCQQBKr
RRAHeArLtHtULw6BMAQam5rPI6Jybd3koWiL+XG4I/zVdRFKP4wu+aGr/mEvAkLT
QNsc5o3dnLxvXrb3cjdLV/hNU0nvNjWwND/qKB3dC7roxAHxBm/bbdCseM2MzQH0
8mfHrWffFUymyVQLmz67vWWfmFpw6+5cVg3k4yJ9AQWlUOL8HAnyZEnRMhHpKa/N
Ei05AsxORbcxNFxNIDwYnNuGzxfqsJJwkbEH0U+iCbZycG3SKhwVoZxuMZ7O7GVA
sy+CjsmywlYF8snWrPZeNhblnmi6FvqVrtmdPzy9XeGVcoxWsoytKU6G7nJ35nOr
y0StJGheEvS+53ndWJscij2FlqTTK3gnpV/lzTd9w/7v/80vt84bFhvuknC8sp5K
PZO9WLFR5OR5g4888NPNiJR0cXMkuWb5vWtMXttHx/dfiIZ4bdUPLzYBjOFQgY9Y
3cI822OnQIN9x+CGx5xSvvfIJVU0qi0XjcgvMRoHdNSy2w9O0lmj6r22g9xJnX4Y
KrDC/kRouJ48upI45wUrfpxIdJEIuddIwdgdw3Df4oIPkfb8dZDtbpSrQz6VpByH
cCDc+kOCmD5eA9X4WW2D0veRuuaBPkhOC0V9J99nnaiuZtYORpqX5xJX/jTjWoah
VHX4yfYee3dRdaOLZJMiakEfao3K1AJSFOwQl4Wl/GCWD55tsBbdtxvGnsySAYiO
0TIyc2l0GERRO5q923RgHkJRGmgOhMuKICw7sTqYYpaI/QZ7pagm7MxL3kTSIOZr
sFCNDszA590j3GSJR/eFXFrrohsMN+4Fq1R7MRWDDPO85vqSAuh4tzfTw8dkE3pI
D5bMbFVt+UdWcSlRjTfWV1LU/DNHrvfiq3ay8ZKcAWHv0xPHuOCbceaqXZMleO+D
ykmk6AaTdrsbN43uGLyaUtkXQl8sCOb3e/m7bBmhxUMEVmioRv0EnfROxdrs0gAE
qRFp0NI50Aez1UABMMYB9aRSuOfmzTZxD4n0aCmJ0aLTdD7GZhuCoj2pX6sLMMPj
Axtb4U2lqxaUPnsW/vPQ8aaM4guCYz2QrH9+peYSnA0EiE2PazbfJhGXQ28yPknJ
ylhFFDVq+9D3eYmRaxsCGkLLf/7li8QsOeCoFut2SCI+JALpwKVOvQ8xqRed31Jo
//tcywfjP+TO77bw9TDGR1/0NWuzvDZFd9NVGkmdZIsWBrwYix1UDl7GBEZvIrLy
OBcOG/XoJ9Az0KqvtFmSrvuSCdoDNTKWoyKC+FG9tEMmqboHMJS2XrOMOThYZPHm
iyJIM4K9hUGt4F1p+2E3I/UxVWgY8tr3NVF4ox78Ygwohu6sagUSeifenk/m+0L7
tWYZEw9WX9+/1+8UXBZcMR8ATHRQu6EUuPt2U977NPkC1uQxitLv59/DomaZ6wuo
yvbKyurC3wDEFcmBmt4SrUPu4WBWAyQhlX/3pshEJQ8ESCkxYa92Nkr1h0euM6wj
gHTE2beR7L7BMG4yIxk+lihjThIxOt7VVIlVWU6WtfnqpCrDh+5c3KWDE6z7BQZh
GnUHiVbGxygblU17fiMDLDGwrmC/JvjRJRprGrWA9YgfVUpPnsXeg4+afSP/2lMR
FtUZPMMmfsdgeJIfJ0nRIPJ8KBHOZwdVsMDkklWnx0CqA8Sd8DoBLUVgV8bX3BOV
hB6gTubrV8TpJ1t0SUaj1sGx9ngeG+NzTzLVlPh9dW9b01XeE+QQfn69s2fLE0b4
11XE9pezJrGWpQn5p6A/FwL4dKfVB0cY01rTKvCGwwTNVgKFpngueq1+IQMXdyTc
4BPFFFwgtIDbuW5GOZ0y2J5/BCvVB80j/AmTjdCD7I9GW6u/pGMNfow84h7bSDxO
GHwWnZF66hIZlmwIlmnxwkcRZAbL2rBL2jCBJB9itgC2oyDDuR6unthdLS8QzVP4
Ge9Ox9Wefkil67hi0PiKkvtoym+uwF1CUAH+9WOl3FpYzSFIlwFXKtWXEPQJvOsL
NSugpcSnCbcfpj6Fcpq1X5yLJXNEFq7u45GkTJpbBt5vsYBit5FKzWpZZ72U8wBJ
Is4G2W9EDqiZnZQbPUee3glYBJws9/Wmp9cQ22OYys7vnOqtxQKOlnW2IFgG7raS
NacvdyS4Xw6NIok+fRLMUz3dzjZPPV1nmydJ+IT1zZqnaH/IktbQ96tViNXBreI5
2+sjnEK7g1xDBFkkGBCGqnk1UhngO2qa0E8hjus7BOubZDXZs0OH2BNF6kHGQHCe
ihvIn7iEQLaRmbVk0PaDyHaUZP/O/1I2WwUXp7WHUMlMhtOVcO5N2FlS84fxu/9x
ZiLURhTUgCFTllpuNH334+kpHXjFMQZUWMgfVDta+slBOdn8wgUQtzGjmwtpiR4K
6wwJ3VMcd+f2lHOiHhlSIppjnob6Yn8DWg6X9A6kyLGCItv9JPJDKydVg401Kcw/
T5W4eKccuOcD4Q+O4E0zo7qOQAHpBmyGpvrQ1tld4pxWMzEavvdmtNMTw7S5YP54
KWsWKKYXD6RtQl/T166Ls0ZiqjAn3bklrGrXhjWxYyNAWJJ3dcdwfmh8VdZzPFTK
asaJqzoNuwfe3hA2UzkQhAP0ZijNBPBvtOlKF7XYOzZTz/ERyChhfi8tn2b3gfzV
okspPBdJgcg8lIZ3uUsnmAWwAJSqeEqaHZSnAUaYZiL96OV/Lsjg1F1eVDhahRax
RF+zv4Pfvx0TngIINM9zB5aQIDnoyCyPjRpm1Rk6LQHkh3FlAzvW0QuK+xQ+JPEV
SQNGAUgRcUqz4f+rkOnZe9ymvXSf+xOsTnLVNJ3Xb6TcZXy8Wr9wGwDgx5fcS+Uz
FCVkHJbBteOfkIOR64KP7tw1pRnWHq9L3Tq34CsD4gUoqMN16cl1zpAm4W7VMRAU
dkblcEuwJ7uVjsp7uBqjFsiIhv4mbJrtnbZjKoh+VQuqdL6PjrndW6zpoIewIhrT
sf/wYEfzar1T8vUtdSfjGahsWPSXuNWKhslwPU8iwlisY2e50d8ScdxPDLRUhhUP
/08TeuuhF3wru3z5hO0Zyaj6fzYioMHh1yCp3z3i1x5HpGKxlw1rKwBfRWUPy+HD
WrwTGdJsRoCk2aPdAzN1YKz8K4VieoZKoLvcb8Nrvzs1+qHCNzc2OU5OdrRf+d8/
o9IzQdFfERLgg9wcpB1nXSPN0h2YORBUtdea6MwEN1u79nu3Pz4VpqpF6oLFiQbc
7MfB1wtQ8HHmoi9LRWl07AXOgr3wNqGohS+eHgklRGYFrRvuYdhSgkj6TOV3Uap/
XfewoNfDB+8hMEDZdMil+rH71NDwVbshErFyYh3dirBpc3SsMoiYsIj35wxHQsLU
/uhcoQ8sh4zpt8cOBcT7DB5yPbUQEwQhSSDAJrz7d5qBpDaCgPBtPluje5oSjqTa
FrRSCjikvEmoenXGpczT8t5lJPa/q6FUZoTchfUmrgzqC4/Ks8M7PF/9fNk7WZ89
ILoPv/GMENVZl9fB0Ziocgrme02t/RoyyjJPvYGn0Q7m6sq6tcX76N0NEYc0qxKw
u3Op7Lq+BmOMKdu2MaWUL9WePAWtc65aNbabdjLjySPdqchWjix+SsFZmJXcgMDv
lEcXbLWwYWnvbfLV1+QhvFmpvQtrgujRULJJR0nJi4a5RH8l6egtcgjHqAw6n9Dv
ecELOSbtpsrwWp6y086Z2mUFW/RFBLh7UUpoTFUZ1Fuu93X13AGLdNOsboKFZPdo
GuDdUvPDr2YLODPYqOZz9lF5ryXqVOmNW7SUVYsDEMKMQ/9bQqJ47p579pyraxNz
uClvBdVDN4aGkcvIg0yDILhFwxZFB88Sx6qC9wYXqL5YQ9bslKnJcJEctjYBpiCx
c2Zmf1tZn6hPkIz9mvi3LFXyPOyW3A1moqMdR+4JxIgIyTA+LLysZHjbt8YoXKKI
y6PGrru2KtF9V//pJHcruwEEpr1+37wzp5a27WP9FSM4Vgt8izZQkunOGtGPUFyG
cq4lGlCWkyMgqRAGYjbjbfIX528nsdIlEPe/uX7XTrak2bDCr/JUnoGaT6qBAhKC
k+y82OFX1YUId+y9KbsfGmjjWNo9VJvclkZhbEZn4yP2juAbsUZtO4qOttFjawr4
Cte2XqX8LcEq7OHtBZslaAW2M1nbEN758gO0/GU+947m+TPM7QIM+UKZkxIIvl2n
qg0JiPnXyiGRLqY/SvvZlheH8l9VWQ7FQozzaBaXlV6QQf2bdi6CHYYRZTHhuCIB
1MebKIv3/4reaBouHjWWy828cJMXDDCOBgCnoaeI5z1/jDAyfhCH8ouximGbpWLz
DYbxlmWVVS7Wow+AbuMZbPihGMorRLUqOORK3w58go0tA0/iMsNdm/YyqDGdZnyq
FBLbFtB2VCrnX7iep7HE5YDXt1BXt21f8WJ3CMrJdxW3eCqtBoZQ+Ex+Hq6GABHY
4s3HFHoNr4gNN/ZPRwBjtfRWE7J+NhUNIShH2vhL7doJBxL7YBlkNYd1uT1E1xbE
s+1fwUK18qobs8x4oh9srfOKfAuZ0UxXyKlwg99tlKqLd3+EfeVB4cv60G/275q6
ei0gPKEPuUPOtW/IRgPvYtPizzcI+neKTaz+Uehlzb/FLSA7AzFqPzS5XUweWWT+
wMWqnVsnPOz0hd16R7XYfcMxgiwuOp6010pbJOJyM6Tmkp0p4zXuG+A1/zGkqTGo
uvJcEEdzGe8NgndwT+IqU2qN6k+gOb/iu5wxcFyWGsSSosKpGpD6BVCSkZPtcta1
oY4X65QayMZcRmfdYI2p7w0yQLqtAx6CSS6GmRaSDGZXTpqnCFo8PQjEZdqa3Y7b
tUgZ0wMH1yxAq2meYx+lAS+5cYqPgW74bb7+N8Kt0Q9yop5cuZvXLehp5b3QPAtT
WEfIdCjYY4AJAyqO7Zw2dY+4FhQ8l2+Itoy0SW1cEXz0MsV/GKLkXLkctYSNaa0W
C6P1G5XVjckTEu+U/rYtxaE7ooM2UhnO99TzX2OdT2v7+kkHg5/pWytZUAYX5soO
w8is5lyzV0Oct9YzOyDaTA1O6Jm6wSurHHUcXm14PScEg4uUMkPviprVSpmyxA4c
u5FV2dgc2SCvxYcsJK3GhQkDRLfPOZxf049LAIrv7gbCutfimkuonyxImq2ZLx2v
hWMh6/6mCy8pQdxs3JfxxSoGaWL3W/v5MMznbjCQTj4KlfO8SIL26SviMRp45Gat
X5OOF6Zs3kgbbBNnthBb0hnc1O/lgaaRxLOQcGeSE8eBBki+lAhGoxQiPj+r3OpF
imDW8Rk8cJHcbvdr0PciqxpBmWqqupwns1+fuOE9dBNmEtUt57+4aSZ7v1YuIesK
CM5bY4DUvAOv3h2+ypp+zqhwYqZmYQAFMWVVht7xU0LcxdCJz1Mf0p6Ltca/LqZ4
1AR0vsWLP5uRpJqQrgOv3RqU9QJv67/x0GkrAXyshfrpe8AL5FgVrA6NoqRTenVH
b98L2gNhFF1zRi19Ag+a8SiqFvpQBCJdE8XitMvyFUFz6g61I5TDyZpidIuDhX5t
7S8zGYEEV4130MzdpK7TRvrOkyRBUeWfMwd6XF4O2u/8N4LS664pKInQPo6ZhVqg
nELQyBCOvzqkcFLmlhuz8/3kdxxbBjiPW1mF6EXekQgMiu9nlJ1LW0We6nQ3jzlj
/5t5kbgmI0+l+OYPnn2UCvsEhhBGEyc80J+JD8Ic8iNbyvBYz/VEwkCnbYL9CRGP
0TIE2CTLkf5uD3w4AO3C2IDk+FyN21yGJ7ekD62Z0RjD8sEaaMckcaFgtpOznzMT
gQ9X8dkNPDw1NNLAslpKmBBzNeGrGq75uikDoFPoLH3dASoSjlAJ2eF0h16bgCZV
Uyrem/mndlUPh2t8RlS5adMMvwr5Hax1ni9ZzPSBVh9oADUyLEo26LK8UpmLh68x
V6WS+i1mnefZymVibOzjEy8x6sDWq79Q9yaIP03rETDWRPwS6tfffxfD1dMNKFtv
xkjmrEmj7iF89Qm7VzffYVOuuQb4EGDFGtWYMjKRcKrIkSy+cLcu0pz/NB/3HFV8
zEjWJvCuMLBzUi/EGJXYPGJk78rCNhBewD69sMFbREYzQUTUf7wAADhdPPfSF46B
N3tEynXpSz7CW5yWObMkC6YXTAj8v5wrxU96O2imVaJm49gHWQkhKLXO/mJHEWIk
4m7CvP9ouPMMMu9G1ZNG6kEw7pkLC7505zjRTYw3YDIeAf3RgIOFpON9134iY6rc
I8hluKmKrKKtSZsZtcMc9jxPEgvX+hGXCiRez9jQLiWFanYJO4nqXPiSufCBEEo0
lGx2UfPEeVxNIrK4sU7gPlACuD2ZafxtlkLSlm5J0D7UwNO7TUo0OoTBNx6TEsqX
Ps4ZGiP6332iUyyx9J+S449sk9OiAb4pdR6EPT1cbzOz9pS5pIfhIGQ+DOQbmR2p
vMfJ9ry003JT9Iighzl9O2DSsbF8TjhfimhPh1aDYZJ9LV4Obp5qrsUKRFJYrDYG
BnHl6AQe8AU79zHF0fpQkvsWgeeSYcj2OVUUOpR0npFZr/9vZ+F5jnMJyeUPYuk3
CL0aiBBH2b+lmJmj26yic43AI63hn3G4Tom7qT+C5/O8Q+AxW96kjVx2x8XGB0Jp
kvinFNS7l6BxwdS4Oxh+oe55Nn0SZBD4lxAfJI2EYn1CZFeXYQqTPTQWZLxLSNn3
1mi6F5R1nqNceqGnYvJDWkBMumTVtxkT0xhG6hErlbr5NINkdgJlw5P85TXElXvz
Ud/3j+W+PnuHPnW48dcsg8LcY2FLu044RFvl1N7Eb692boJg+sH4ImT0pjjbVSaA
a9eJx1jHTvKvfJWZ/AqBJ0nHwPFfOahnXK+EEreXTnSsZxVhhmco1dMizRhQ8xGE
uhtt83ZnuSS8q2HGYuX+XJVqSy2KgXVXrjhQrL7u/uWIdJfE0BRhz8ZapyVUKkEy
+QETKUMTeF4oOwoDM6l/hJdoha7cYtxLAdGcHOUoeOzj+oZ13MH62X2oVrqmvbOs
todgfwX/phqhlbq8MPZmwtK612pZFEVlf5BaJhYLP6XAmmNwkmWlSjJeMhYeN7zG
PnVbU0WsyGqiRXerQVDsHek2c24ZRXVURCyX27CN6EWEAJHeiN3XemzvSVGsKAU4
2F69A0MY4h+ep4gRIB0b2/LJ+drGgnHgQ9WevZNM3eBCmTWvLG1+4Wof8YjXqfmt
rgPx30IbIHhlCe7FTY4V9DCY2kRDD+6NihHgvlhZP3I6u6uzLMcFKEeVlUONhptN
niqwstfbm05Bp08xSp8UE+95lorLXwqcbgmz5OH+PaV89CcJa+SvJlhqbgWFjcSq
sOFpz+s/AqHbMwy4wq26+vCNLFkCgr06BgmG7Q0ZNYLKCKZNjZz0eryaK/Kl1fA4
fM9HuIwv1yk/Rsvqy3Z+YPfPR18w/ieJ4eKJ1bnjGwRdggyQmrudsC30Gf3ucEPu
vPiddnEQUIodk4+XGBglMoxEoBsuniSM6BqVnlvcw/+ZGUbuZKM7l+EdMcTGzivE
y1VFmIF/w7x5W94RjXhtRqMpkQKDA/tCoK4r4LXkb7S3rU2jwF3GEPBRjyhEL3MS
NTpAus+f4XXnZhNjeUwEC4fS1YplJelzyxMSilXy6gHwWR4URUU7icVJiULt+ayo
iTHu6yJmor99P9wKHLJimHm6rltLJC8ZinTRwnjNu7j7lqbRxhhhOP1auYH9nIKQ
xXkN5WoKa4WdoD35mie63IDNTuS1IIAoRfaqvMbWxocnedZ672kbZuOMFHTkkRyZ
l6F1OhRTE/jSGyBE35zGBz2i2RA3dlASKxL1wqyagbq7FETmHijCJT1GkEnCczMX
uxAv05HpflP5LlhnWgtUP+vmYFw4/xvaDsnDRpv3wN1ythXgzNSILmfZOnvnpi+4
DBOV5wO8ibUNUFWaaKMnok24NjwW4jUGhY1sDLJr9V3lqrQrP1Kuyd+rYtvwV7h8
IrqvMBNzmsQ0ZGGN9/QA8L59K1qK4DSV922vpepcmV19rJ+sMIVeycilKqbZwuY8
X0yLNeOYf7hZn5JF0sqDpZR5DXApLx0iYiG4Y4tTbCDe2wTKn9FasYSHWGzBQceJ
JxQ2AofEyQQS5FiuNgXZ2eULZ37W2/R1G4WqxLSydLfRxb+55R38buWQA3MeIZMG
HjJblFoJ+Lwfmx7Ce+pzLz5y/ii/t+RSchtUHHh4S+2XZAGQH1HUSzgXKGDH1X3+
50WDUjEIQqB+Kk+iT72krJv5HPr8fBK063+/gWBElZDQyP58Ty+XEpmemqVfhNnC
Y9k4qg0xGl4rUTvmRwKsjPrFslZdYi69HgqbWlhSwUC9vKkND5u6ykz6TNyJV4JR
W25/9eOH/wucjlwJpqijNQhB6gUxhBlUZaGd7vJLUrbeUF0Wf/3jIlCbKZeEhDd1
CIsjTKW63Ye0qWEUssbJSmhLy/vGuMjtbF93pgQKdN3vLn8JZ2eoeG7CtEapopo0
yY5/ZXlcnypzGSUQDTTVOyDyhq/DzJ/w+gd/4w0kB5JK4MqMquvJBwDIMH0A6Fwk
b3S4/kVqEyPFdjwKZKCn4cSKZelRb8ttY0Jz9eTh1eQoZlZvniAwp1SgRdjUBmK5
Ik/CoLTPrCZeXuvmYpFEglJ2qmZogyeF3CUObufR9tuMC/ZLUxQG9ezk/dQlaiT3
L/7YkImceL4XzDg5v8WCvt3tXuHL/tWtLRTbAz3guH29NA3eELiBo/svbu+lLzGL
xAe/4/FWfM7T6bSGpvKqiyZk5etcgJBMHfYSejEbECrVxqk3bG5Q0jI5/+ORr2o0
rjoZrc3lPGu5+1IOEowUFOZKwIANZTEA07GYAMEbESB/TczBdPy8fg1mtpy+n/8r
49zrnrE5mL24llLiyB/ZuZkoz2yLY66APHZVAPw68KlS/dOMqKDydwXwedWNmwjs
3wHgeQCPhzkSpVyHwcNwFazr0S5JY8isBnOBCLBCYyZbQZ8mZRh22I5zzx0p68Gr
+Znx0Li05ce8PFyWowl+slgFyc4Xv4JMpi9Decy2IDP6VhuhZVZ53sLwwJiNgCwY
AwnNmdbXt8f8VLPSZJlEQv+sRgC2379jLuYiZu+6kP3rrZelzlec9IxT96vAlRr1
WW3hJHbDRalo/CBIWZm79C/c3KgKKzvsfmXtm/PhcRmlzFydo8qH/8uHTP96eofc
qfhVZbuHjNGHu3zkh05J23INkZkJZWEBTHPSaFV9C8CCF7/ba5oMm/cvf6DcGriv
X5MWwqaeumWvRjDvFkjQP2qK0MuM0H/OK8JdCciCWzR1LnH4wAJZyc/M/4EodKUI
9lbNBzZUf8dfuyfsfSVd/l6m8oEaSsxZ3R5uLmJom6O3ebx2IzQPn4GLP1Y2oqcL
xGUSCgpPI4zXR+zWmYBGmucw4TysrPrVhXOe2WafqROQJHRXed5M+/geOphFTqxz
p3UrnwxqLNO8H2BHvZPzoqiDQF6hlbrSQT035xifxT3gFkVG8yekcvRqfG1/yBF6
c2dBMTTdC5fxDc198DVIFGYvaViMr7jDlh8mz3zQQ66L8G9CZusjXCZ+xdVjC/eJ
uP1mnN63GXti1VIggFAKlTt7drFjuNRIjgovvdayGpu1GHRfcv25ZKAyffss+BZJ
zcSNxlGFbdmm3mzVaE0o72fmRqbSHwHsFcMK62eEQ4syIF3PNyptIkweTnrloaUv
6xpIUbDcIY4EESMCJc/3/6FaluBouf76fncKHFgwIb5xFOS7wHmj9GD63KXBX561
YaPJYtX6ve0EarAXDgYMTAe6L0Ykt9MYGK3UJ/gbFGJaI70E3Pi7B3sBwWqYSe8j
Yk4zdScluJGdjvUNOJ/6FYnMBbBvLnm9obako1XKA7/8JEXhdPe2ndCYjCxnuuXY
no4TtoyE78TdP46gef5RYVfgn8o+hOA8Pu0HpDaZLp6XWtMcvF5ZQJGsFuKOiVeu
2m12IAhca9qpguOjqA/UvUU9GMJj77m1X3BcSsGYGGTV9zlQfeF5kHGVjRx0XYKt
ysViAuzYRdGaw9i4rmDH2u/8rzOPn/WDr3R5+973Q3SoApQBLbkZ2MxTUhT//32d
hdUCGKngsmQ9yK6YpoJP8MGHYcFDe2E1kL1suoe9gxxYiqClnJiOyQ3ciHrANTVJ
lstFd65VaSFGp0ilzyZRg4dnmDpdrlAJy87ky28HF1CHjhbIPkvYIOOmCkrUe6IB
O/ML9YZxmxlwo0K7x9bY2dFjTV2ryDVG0p9qRZrmFPyxyLZ9uLE45dO6SQ4CQJ8y
GEq0uu/PdTEK5sApHD4AJk98OZl5gHenlR5vi1yLtnvc38SMOPIWSdJZgQNDF8Ty
6VgV0i8kfjsHy0uwp5P4jJArHrGx97GFAK1DpLzXZX69ZaGkMdwDnfF1XUU3E7RS
nSvhsuGzW2nyyOwGhhphNBd4nbSMcXd/mc5qPAzrv2/jUQcPKnatTUoEwDcUkJpo
06mC3zBcgnjsHffkUrGOBK49QA8u7Gmv/98JrB1MwBD6V4L89VdQsbPnyo4xSdMh
QJzaRWm3RgMT/S7Imtq6xt/0+QKSx3FoIrt1MuPX21V1VzuM4Z8nnXZeyklembpc
zigIk14mI3LziJxtxOYUKtYgYB5iI8iw+mx7DobmGrF2Lw3gFR7RxBmdxS4vrWZQ
HgTCQo46CDIyzV4HCk5HeU/es9IDr67FZMCfTdmJ2i7rWY7Vrk+lH9sLAYF2KOcO
n/30r+yDJR0F0VAOBB/43KeiaEKYbXR7vwY84gDOJglMOB+h8ahXMzND8qDsVtoB
zlX97x121fwnc1Ad/xhi66iv3U5uIhZCm5mEf/w8k9GArnxH9UnWVYtsVaiClph5
0Rev3hnFLOdvRxJxflKNJ4gYgoqN1LmkaenQkJOE1++9RW2+WwRu0rtIvPGsdM+I
tjm4nDpRH3/cBEfBgGEIhV2E/NQzWg+tqjdlv5fdj61Snojsz761xlKOlu1F4u7a
nut4RV5EKBf3A5ocERngjYXCH+ovqyycBFG6x3MXVhY8iX8NDwMeXRxvF5Nw0eyf
On9B6VgVeCtloIsgJ1DXGYH+gmP7sdbA43ajCNfp1htyIAbH5h/CQ0ql0fjFwl7E
Hm9oPAQA/rc/OcyhqvV+0GmrbNYKHKia9WFc/RHViF4iUwHLTaLfprSgZM8FNpMJ
hWhgNz91o4YL6awh4M3773Mca22rUAJagZz1WtjMkXnY4H/0bDuZfQm7gDuMCqwc
kBYOhZV2l05Oo3jbYjmcCiJGO2MTWqosCJ7nZuA4IT1x9swW82CQIAHFymG+dyJ5
bORAsVmLROXyUHcpb7rbnv4fxZuEFGNz08iKnfAKjL8t40md4f5EmA5TOHibPKUs
BAYbDTc+m1ukI6gB77gGCycaYI2NrtUIurFUNQdDLwCngY8xHu9KkAlnfQb1VWZ5
6bC7jZxwkTNKVZ4qrfHxJ9pIsNCvAdEnW8QnokEAoARzApQv6reQE3p5XYQiIc65
CnQWgWIDuRXyJVR54m9kPJlXh7689YtloRJvvSo8ryTYT8Y8YnOnyYwIskXdP7sB
Bj5Daie/6a5I2ozPHUXGnugxelaag9vHyg1hcrZ5juJLT4XOfMG4wmHbEfNH6lgA
fkCGDyAGc6Mp4rRafTu43oj1uuw9D27hn2hEHoKKYyJzeKprU2oqIL6TBWkcz7Zl
tO65myl62DRnez+e5Sf/ALGn2nPriSZiYAyRqA08veRM55SN8G2/Rwg9YHW5P4AQ
Rm52kbzXcEmt2XuCBIkkzK7hHZI0yn7GzW6VNQNxOLHH9+z3m7lGhb3RjuMSgJ8u
/2/PDRQXoFLRjXYOGFS4lXa8fmpoiLXa3cit2s6NSyfHvfIYHMDH2GKZDeUBMEnC
9zzH27reBG9JdXq2qfL5Td/6bhMvVAf5xpg464xfL/LYvJreBCu5R9xNqftcx7lq
CUjlXArAfHSKc7GlI5o4FhXCpuEnQsSPtu78dy6HfZsVgO2POodxKMdP8oiZyuEd
kXmemc9/rk2dbSbON3uD9QyQxOkLZr4hmLxdeZ3BPYpzQP3U4w5bgkGPj6ztVn42
dkM45rukVlrQpN9AqHb0OJDqyxgUizqmt6ivO3qKe1fUMMMsw0EexqFPRWLJuvs2
6NywuJjqWwtVX+Szfx+53yjLPPSaMExRg3xeWGvdNahKNj57F95BxL8v84Io0r1D
Brk6efACuNdDFCVZl9Fb7AYe9EvE/B0dPnWvFLmRMpY8r/Yxx0p08b2DhcrqGDoc
u/+OZQb4hiHrpm3TlsYrABOUHlCtCWfX805ai/Bv1/9B7cFZbdN0k5QzVYPBF5Yv
laXFhYV0p/fOMAMvICBLG1n++dvnHJWj6FmwzM3s5cDaivqO+g5VScZWm4LxF5vw
eQI40zDTSmKLOsIJhmhAPF7W7cp5ZWHTfOXLoriyJmzAITilof2Dpp2upv6CjlCg
lRjdWHjmJsa7HOPwVvU7ZPtSSC0NSod3ZNUTm8H6PdbgVGgXFEMLbBz8qRSo7Dzy
L/tPU4B20Xgmt8+e6pBX6+gaJmtyYIUq2KqsOIBOYrI8DchrRHhYRVEOJGb9qyJA
2OVKpW3iG/mPtyZ64dSXpya1ZttWTfihKc5IAtCE5+Blu+xqEeWNai5zFQDch93p
wpPrtdmKeuapQ3Rf5aSNRzGTFKu3c4wiUQzz/q2KLA3WDDNQiqVLgMEhIPuN2d5K
GUU/WKSGyoL3VQE/onULANG9sG/KKr2/ORaqogfG4a+ME8NtaXsuXjTodsmT8udL
iKkYdnCzS9yn/fNJ+RVBpVKL2J+OiyZQwuRSmeFLa82uz2eO1OUSCvAb72my2TUn
GFrF2CWEnZPtuM/E1wUZA89O4MTk7DM+CFc2VFBFFHyaP4OUUiwEtdl8X4EN25va
HFU8yppgeRFthfMFqoxZ4KL2CHdarZlWVQ+FYV+QE2lCtm9ney+NQBKgL0UPvbs5
VtFtle5tA4ni75egiAu20/0387jRwtC0wuo6C5RymhXcTRqu8Yq+ml1aYL7sOtnf
6FrHAHGRtBmvzu89xXu4jARilEFPQW8Pu4oWbnM8C+CSwTb7HPxY7oc23kLrV75+
+hyuQ7w5sSobFSm1q4RCetNV8It/LMTECa3IieztTXnc7wgZKTNjMK1RCCnEiagG
76YLjafY3ejh4eX4Jw0zwQjjEP6PAxYRJbQx7V0kF4cWLrOnlFeTUski7qbIupyg
NJniv6l78mylVwQiJR53HzVAZmoQWYzzxLrABP2i+TNAVnRp4HGAqzsyEjeIvctf
v38xTuFCFLa3NETZ0eSw3bTApuUm6Pv7OmeuK6997dvVDACr0UtSRO7HfHzbxhfZ
Q7OodSiWRUjQy1qSW9GPzXcAUWjK1wyP+mem+dtVXmvVbT8+HTVmMgBgFQhjYicx
uiRtZIq8w/ZKQfDGTb4v58nBf/YgzDK1VRGJGnlBoYOZKjlyFxmjLsme7IyuUJg3
cMYMg+SHCnzWuZkOq25PWP5m4dybaxVyZWIXzOX5+QDEUGbIxW6G0NQHjBVIwDcT
4Ts+etvL1Q+xoME/ISwTzdW5GyWhcxwlMIHfcDYpF8qrrXnrDFpy1tnZPafEVR0h
SQWL24UU8y1NmAB9XPuo5oGOdbChRzFCKEa5DsFiChVDuo2KpVN5XyPkWqvFWwvj
PURK6tBWJy7WMBG7qOkqHdfU8Y+IOBLPsTpi3PHq5UppghichiSFx0UHJbmQHhqr
OjiZswjkzztn7noFwdVILLnZ+RtWy45eE38/VYRHXDPFrDT/JGvjA0cpRhrpeiVu
s3Fx5APmFwu56eJs7v3zsLlJlkezQyDg76VrlQMVUGcc2kCPtLwAVKPRpdAIuFfn
I997cHY98iqIrs8IkGZIzxJDilVLS2YQka6icKA1YHTy2B/Rjhi6/sxpntLxQ3m5
+xPbavOLUL0tpuRiC449bSvWkI3CFx7sjNTCciCR3lA8xH3P1oVCH8WMJ3YCx4pt
aPu4o7VflXP83py1uoqPzs4FGgdGaOwhsg0dbeMQeqoWc33eHgzD7OpRENZYxPPb
AgFNFt7uSEtVwUWMaXIVq7D9ufH8fDZYcKA9kj6G3a9od7PvsknAcfESo/ej7vWH
a26wjk+iKpg47x1Gbr5F7Q4er3K/2cpLa3IE47BgCaBQNc9FMBple/OBRuTcADWl
klqWMIrFFmLWZG/dpzYuyRViuOWIPvr3Q3xdhKBkm42+1Gnc/G07daOYCajR4wUa
sSwGLDhhsofWxijh6O7rTL/npveW/XO9PABQ5Pc5MVpZuIWNwN1pXq1nPKScPjqc
SGZJz4BfN8JDjEhZV0gLw3B11/AmuwE9ZP4NsdvIStIMbEy8CQXX6lGoWoHalVoa
/E4gRLj+jH24g/8qjj3hSBEMPRkjbjhIjX53a+ehc5A9KuGqvEzcH+19JsBLE+EH
GqWSJB8M1RXDi0gezwzXj7rD7DhJKWUJ3nx4SYh8lJ8TXtQzPV8vlW9q/Y1j+mCv
l+2QDc1+z2X7sTlhGxbiK66GWt8Hum5wHgN9BuoiBtqbwTmSsT5I6YAULGhpY2Xu
Lgh89WBsuqsm0ZzVTefa0pvID1psD9sE7agx6hP6nxo2pAeAdmvTP+udHnXpdDfT
ViX75OU50wvYE2jqi3ORBSZuemVctaui48Ibo82eH2pDJxSbmw3cHYuEk0Dpa8VO
tdRAUVRQ/iZ+QILvaJkdrMlIHIStDYCzfQC1G8jZzGSbBQQzn7hcknM7WOddhHqU
m5LZamX9RHWCT1++Ej6WMgteXiJMa12/kv11ZxvSD57608gqKlGAyI5meLMAA33P
W7d8VBJYRMeHiro+AcwSZVJboFOv2XA0cCvbJtVg43bWs1Doc2J32Pjf84620TQX
hp0z3MNOGZEFh6XGEVqBZ9Jt/5vWyNt+DpUBc7bnLadoiN9OT/WoR1k5VAT7nUu9
pXnQSmHAsmr+c0vKZIkiDCWvN2NzhCunqZ0nWfRY7OTlPvaUD5XhpieN0SWmzLWs
hZ7Nu3X1aH3jM3/XmvYMMancr/m8ZGdTw7m0Y+4lKxYeLPIirTcKSvvo0oQ6nFnf
7jXtq2i0I9YE8GsqXJLqq8WP05Rm57k5syDFRWNGSF3XaEHxHFT2JFtrInu7c1Jx
TYSiEAyfnnjNxw3loKUmMismZZ/pHZx3JnitqAbu5po7GlSqsNko5Z33mskQ2IBp
5Z7025bkyiL/oL9Sj9pVg4tRaFvNOP0rdU83xgnA6qZJQLOmW2qlTACP6WlQ7DMZ
MRVrbsODVmbKJtKiNGxb+Bv9U7JM5xCRZH0nSL9LbtF6jcl0TxH3tDHungxkC6tR
fRwadjGzCI9Y3HzGHwnB0DHSZg57EZQMCVMwAMiHmG4snKzMp/Wx/y8YcuAtDC7P
HKOW4B6Ubb9+v0LYX8eTQkV6dJN7Dm6zQ+4ME/osPI0wLLOr2N3I4cTNyfBwePeM
7iSpkC9vu2cN4BOpRLmjNK5DqPml7l4heu8mtHkEkAPfl1ncxZ11lfg5nJSLa51T
UjWnvg32yo8Is2hmkrNnJnVPTw26U3WnpjrXArwVwiaXJsWFsVvLnE/Ig3o/8vUq
F7DaBCheHIfGrFum9BlWeW92UNbheWzDdHUGlcXvZkM598vxuQTB54Vg9JDim8pY
fUR+nef8Xn3Ry6hspjq3Z1RYJHNzS/N6uNlAlB46b4Os3sCy/sTDfdZlddlc4VLm
DtsH1qcu1+syuFtznjDnK1puEg/u1xM0HmCO3Ns2w5yQqy0gXDUvNI7xooWGk1lE
U3sK7EHnpzVqjkC3W8m4OtfwdDJz7q2B0oiuIpCH1JnatYJa6/yC5Ewndn3I3FKP
FzXfednFA0BUdopDalbNWbtoWUpSphiyVKEdQKmVgcAmUoVlu0qWPAa3lWDhbebB
aTui+eLeS0Xs+BrwLGI7/W93Jr05ouiU/RWdU4GazJx8aKssgvz285DKnSgqtmo8
MCo0WfXGNUl7WnMFG/SKBuS4GqlLnOo9do8OLbBTs+CmLIl4Rv2abiCGNfAHoxXZ
J1tN/S81nGi4RIzXXSxzIrL7uXctwTvF+tMF4oQr/tGhY6pgwOP0I/rlgK10KmjD
wt4LvVnLq08cbxGVk8qQW7SZIE+l/tSilK3SP1SR02ceUNSZkjRDL1YjEkRDe3pr
C5P3lIyoouKHuT09cdoWzdfxjeZjNC1z1bwwNtAAFsOcxoWVNC65mpI9aJm/Cxgp
9+rzkftmDZGrmfsFXTEWcJCbSEg6W7uWG/R9WV+0/BLh5oagpTCQ3HR7RiUSG75P
kydddfalUrwrf+N8m6KuHkqhFjlmB0J+6pBTBZw7Vhmv4wST4t1rxCfihZMMLimU
crjc7lf9EEtIrFGj04+d9eQRcI6TVOyKXrykhzz5U8NBTtBtqOhXEd6jLq8aOQVr
CVTM7YSbs/DKO9M/JuNdgv2IRryOFW+enKj21fy2HJxKM0qkbWTGVzOye993IpYC
7MbvB9X7YVPKw3PphxfSio4LtQgAFw4gpu4+hYgUYFw5D6yslQYqHsZ7Y3q12JCL
iA2IcfBMyTnJD6W+bjGvvjJioDt3jdbsHe/83TBZAxOKY90wu16AXYl/ftgvMXtU
nOLeNIL2KIRj6+ZfBmOlTgXWvyC41Wq4O4GQ5Tf5MgnYnja/9rKQ2XHiY2a9tuiW
DbjXXF0U/Wv/4FdCRuG9QYdKuiF4K5bxjiYScVm787pqGAttTtw5QtM2iOLkmvsr
XbeVxbOQT0q3dm3SeKbTXxA0MbfiRkRMrpx2vJInc3mIeieM2kUznsLzrfVzxuJL
X0acCKOWU9ov2xK9NE28mVR62KcrWzkjbasQ5jROIlGZ4DIEnTLumxs72hUGsm1r
uyeUKEZ5WzFOkypUOsuJpGVNezqsjbPu0enDfzd5A/xkrinmZwBtpFw21JbyWOu+
pdCXFHJw64lfST6XCPvg+MJxnGHqQshTXEasqejB3pG29O1d9L2Sernl+X2ZFKLg
6Qvi+8LdsJxOMmcToXAOo7wH602mQJBDk0zVtPaaly5u6ErJg7FumMGr+Rud/fw4
flBL1Ru3wF/NFjGi/UjDAC1kz4VjrKrOI2BqtkFOHTXgoTXzSpezJDs/6gwpXLRr
55agD6hyhTjVI97GnYXSHjCgTB+fBfI5GD2N04kw0ea5XbEs4kimACyB5rw4Cgpa
+BSsOno3ufpqK5pETJrRiUf43z1kxJ54JAcS/n47bQuFOfetvjN6gH2uwnpn9RLd
pknRW1tIGzm0/XVuvOPtxKNLXO+QJ76z6O6FVDRd6AWpsRGUQuUPXnWtnNwc95cY
sgNypvYMOnYcqzJ07t5t3caxY/sBgwEJeTSASfdMfLZUIPK4Rl7qGAakQMYu2sMZ
nKg2aocVnXdlbpLTYZMPgvqiswqwmXPt60hEPMaOTHGiECLR8WW3ouYE/vD22h91
4s8kS1VG/CsA1aLu2h0FYRMnEcxy2FfrRum5sQFFLHVCIFhGaKW8s6gBG/lsjBjg
nNVewV20T3DeRz/LofRzoZmW5ZggH2GgkQH3ua2A40PvMxZ20Nuu0NjLyb3DiV61
bZPwL4aVQoMqLeDm6ZDGFRzSVkSQWOHKqv+zRDmrvQRiCq3vFmMGvXIkeEuehsy6
hLQBmfLzTRZVJvAUiJcJY7V9CTQsXplsETwzzb0ZhMH5WAJfQJ8zDvJC16JpJgUV
9Y3THqeBpjyhPBrVlQkojCF9BAsxICRqucJVLWTihkZlNkWKpPMrNEyba9VZCfTj
2kRvkY1IZSKBltu0W02bsO8+7lTErAMRlOWLJkLalQp1EpHNQPIBlauHZeyvr0cU
xHcBbxdQIZ9dgmh35Bw+WdMXgArwP+iJBhSKo1f+NnZAWUMhPs9ujM7jpJ0lZ0zy
zUPI5Ur51GfemxQBRRG0sIrTrXkO8C1dlaYiNg7AvE3lQXOzzK1r6w2lpa/7RZ90
AFhJr9kzY0yypu9DbXdALK3aBsjiCTW45KBFDzQrlfB2WXO5pSYhH597DOjNmd0J
o475vgcP5mNFgskRcDXO5fOKBWxBxWAcGlFQ5YU4B9XxX+T0eEMYhYoXqk0Xz54M
O5B7BSa3dNx1Rp3I3vk2HhuHW8s3k8k5zosjT6OnLy7P5Aw7vDP+VYrPhYWZSCWS
lr5nnmFQHyQkk9ASN1cZecsfKPl/1Emp9utDPhd/ZtlpN+rUElYHnnCw21zCEiX8
CySlq34tNxLLaCRF46aUDuhxHzk1AWjmi1wNuqojhsSpksBIN8k1OGkY6XJhcPi4
w6YG2vleiCwf+TlTh4xRJIb88r/3m7Vj2ahf5IDQbyzXThZXs7tBlnRUZ2jUKVVm
zqPkZ4fTKUPVNP/IRigGfp1lAUc7T4xZ04jiBypccF356i+daLJqbNyRwFJywpAI
tVG0K1AZa5qimGVxs71IgXrN6aM4HRY3g0cLZgKAvmwkOb9MwwLBGdF+Wt9f7/R6
t5xXkSlMe0OiosJHsAJTN1nAZ1Zof42v+EJzR5VBO0ohLFRdnSrX7jySgSvPBaeD
nS8K+BNe4Jev5oRf0fnxFQSiYG8LV4NL5qu0mODVsrNjJP7wtb2xV283F0r4M/lF
pVIbRtPZUBFrf3ifckNCkozpj2Fo7Sdud13EyIIE9WA9+KsrP5Vhmqfthn8yrSQk
V5v3VJ6YChANi2VA7GLSacNEX7QrhL+0pDNUIDg1+AgSpvDKlrqLJMxH0ufxv2RP
MQtEs27C6L46C6HirGZzT0r6oLM+KQ7KwX7kC8YAmMWo/CQcC6eJdp00ycvrhZVE
tffdpLuEvkl+qynHBHQpohDvnWlredecf1BfaDFONZkKuRif7Hd3lcURibnY7Mto
Nb4BUaYA/oGZeXUjXXTwpzFsHT6cm7DYnoR/xfPX6OIc9YZ75MRbpvMpyG1CIb9m
4+BAw5qpFgN3MrWerza5ggNCKvrdM+RVhH5vXEIGJ3OMATURShx7yR/klcM/0v50
CjBkp5Hf83rDVECaFNu8/mPByx8mEyxfs336RPGPLvei0ewWQOABQ8gO9u9w17Sz
VBpiBtLOGgAJ5J0YvmDXyD0ce9hqCZ+KK8SdraBKye+RCh3WPrMhL1gQl44jlYB4
SWv3FKyqiVFO5EDokc5bc+QykIYmvI3h13+084dc8cICsfrxCc9ppaVbYJ7zU5w/
mteXSf5SrPlppYyKqIf2KuuPpq6zkBs05RU0qeL5qUhCXBYnTXZHxgH9Q/1JRnqU
axUxzrQvBRMlkuM+B7I1nw/XzUL/oICx+QQUmUtxWE6cx7t9IPrqmM+tCMAaosB7
3Ro2p/xz2Uolm+rUSz9xaxClF5rf7LS3doa14ClfcdFccdjkuxaPF4gyoCMRPBio
lO2xZkHR9NmNmEcJnHXIYw+SUiYM1bQP4fWleZ5apeqoLiZ5KXxkBSYL38vQok84
PyuIY7jaKpoNDhljLdpenwmjGvWaPa0v8OFE40G6JYHsToGtigQx8jRSGD3WApca
rXC+ODaMrl13Av68EBRJ8lLvwP5hgnkV8J10tHtzS3t5YMEAHnyUc/gqxLSjDBrR
0abNTbda7RQvSAsb/3KTVHvzwjQ7e3v2loAafNuo6XZ5Ot8YRigf+r7ih/3WcQ0v
LlQROojLjDeBaIefFKpnsuJkTijqO+rpoYFjK0GvN2Nnv0PuEtuhty4w8gHg8UFw
1kLtxuHgUZTZ3Kbql1rlizCI9s5q4s73t7rQe3J25QnXN+NB1/nx4scppnuy55nM
QHZuxlWg/dO4RctfP3Xmm8Vy7mng8n0KuZALQCWCac8RoyAUEHk9/OmLEtLrkSn3
krF2LFMBT5N6TZcuDGKysrVHa8xy3fDA+nAaPu+wBTbyOlsB7GPQVHRzbE+5q1KD
KaXELB7W3mWop8teCjzqyvP+M8RyJUa5HQrVZw1sn4f+Q0jd3/hFJcMhVemQgF6v
esa7hvoEMpOsXBcMvB8N8YaVGsqfH8kjYJte7m8EvVWdFfR5m+BhBwOsN7KshtK+
SoDeWVkLugBzb+Md966HdmQzug8wCgKwuTtFWoj8mQ9T8D0j5kUdmeaxBeNgugAw
O575K6QhtGV5/iwK5JtRb3v2KBpvtZ4KqfcVglnZuJGz65jpZxR77R0EPG8AZqhb
+5VLIL5F0otmXKju5n0d2wlihx+Nx5uGw15bob24BrtDFIFBkEdCdNuCMzoUH9Ry
C/svUr0V6MjI5ZujkasrinsUpVuVGVx+CpmLoMfcxbJKl3Fmxw2Me40QynJ9YOvT
y8KDAH/trMUJSzZJeD/QrRZv+pUFZtZ5yRMN24U4hqzybEXD5zuM5jYQa8CdeyDW
2HowEwjiClX4aVcBqVnAch9eFh4eqoEZ0z+uPFFsmyXjyw5/JfkyltsvEGCh32Qx
gy+2FkRPDwcFQjdb49KSHrPJjbJQYq9OlZ7G4HlCq/D/NAZyEczx5QwM+b+wDfPe
Wunpprk+EAQYEvu34jgpbmZgGCj2VUAEeCn/zmpPwNuCHnBI6nLxbHCLwpgqsHB2
rXtakOmM5l/bOLb4gPRe3SKIO8OJM5dx7s5CBA6ovONiLOPuMYR9S17xumg8ZOh4
OYKPOwNGyPgRRoFFfriqSXTRQlzC1tdvnzQPqfyFFtDNr4x6zsIQrxg7GhEGH+lE
1/ntPwkv6AXUopR+7L/WmJn717Dw68/GRM26ZniSDFaCE2b96cptHN+fyl1YwdPk
Ci5MqFwiteetbQ+5cyXQsSLz4ID1gbpX8FV64fV0W4olQdUHoja0bbJSN/3eznJh
Y2tbfYiFOoR70+h8+nAwjVRjCkErct9igszdSuYvqzcC6Ko9Uzr/ayo4w6ywtzVT
pZG5H2jaQswHZdiNW13kcd5qA0GqnalB7zyBiEjYAqATWMZYkmRB6DZe1unqbG/V
SpCvDRWE3uKV0qvJY1QaLBxMtpZHVTR9JIfZ9D+OhLQyIhGdcUmWEaybrgIk150R
OXV04y55Ty8CHSe9bjvX7ymv24ZF0chQs9e20f/HmBIm/4vCaxjdHgYA5l+Zj4i1
5dLYzBYNuj7tZos2hPJTxYRYlmzpB+1dsAsMhxfx4ona6b4J5LPlspbgIsMQ2niB
FVaEwgHWCb605xPCck5T1/ak+ekgG+PfFGaQXdQu1vac396OeV1hRI3uo2XifAqE
65K00VP5Bv6a/uGJAUFRNu1JIcziYilc7LPQCB5XUTs40+O/Si4jJiPua0yoTUEM
eAZWO18k9qFkFDrhZn+hX4fiyEMs6LEDLd4L046Y9fmyJNopeuvcJ20qyWcCnFx3
Ni9CFvIh/ka5y6jFVyZVvK/p+G1hP432UqSWn4myUPIBVQwXlJmOzHQTD0dySf7C
mLt81PcuFJdj76LSHBuHwrc5fb37qnd1sIVTdIB0rKGoB35+M5yHD/DocJcpKPZ4
dUIm+il7aMUfnf2OUWqoGpCAQ2xXyXK+JT2GbDsvarOVw7zM0wcqgXRICXFb0iBD
23zyj6M/dFD/weTmQBg/fa2PcqIlH2SQF0mbx3YJSVIoQS30LW+qB9cMGl74J3KL
JhS1ycPthRQ5Y7sQz1SM5WMNRp2fjHyed2wqGcoxzXWEDhh40nBls6Nw5EqbEp/3
ewpFO1pS7l1T56Kcg3mPxz+T/uFXDI31xKgF81yyNQAJyKfi7ctPADJuF1AiFUwt
Q/7FHfDFyNSBD8+97uXwAwIoL8+T27uabwnpa52AcETtWzRTajotTnW4GSYMulmM
rp3JZkruPSw/JD8XtkJ2msbz74s69+I3iZ+T1slFAXwlMCQmG3X0ITuHpWBkBe27
t1TJTFd+kMpIJgf70fp37Qw21mTrCpW0pdnm2oDrk+r5qI7BTcVrhVbhsSg/aMuI
3bBvhm7hAM1KUhb5xGaWuD+4qyy7I7wi4lMqDqsmWgyGg8AxHrfNxt1Ly73cyW3Y
Y7EwQWh8lHyHPkoVfIJ20a7xf6nEZUjXbNpqgXYuofhDaCigebtM6QngUQgrEcGs
Sfj1SMCmE4u9TTSLR65Do+NLy7usZif+lLswNKYgP69V84sJVXEPOtXNkjrpivS4
ZZ2FY24n1hgcxl9YngxRQM39MieCpNL6IrYy0PL0qJVde3MEeGG4bVwk4yzN9gOl
Ir95+lp9wFGeWEZ3deszRivR0NjZ4q0sVZEoHcxbk3IyRbGxVZJcc7s/o8WisQOR
fSgiNwp24m4gnax367vdDEHyJl6Tpr0Xyglt4iaR6fGDsgGCl0zjOLTA7ucxb1Px
aiKVpU4gg+lWy6Sm11CZp0vDYJQdg6Uu3W+isvKCJMg5nLAHJbnOgJ2z13D4hbKi
sf8S8cpn8GGoOWpkwiCiGLNRkKs2Uv08D7a+CYQLmeSNLgFhoyKF8fDuwM6UETbD
5NINT5O+nV0IU2E2ClPqs/XULREn70dhyVj4JuI03/hzZ29BH8KjZo1qquePvnJr
ce9c7a2I2G5SLQAK8aS0WexfD+6Y4mhg8rH0zBnzEx56D764X8IORHFOBGSKDOcI
yt8JytMI2Jto/DJiJkh9k1cgSX9qehAOt2HH5AWEFbaE1Pc639nIPJhytABUYEp/
ijLvuOgvXWQOuvKAGiU90hJvZ7M5iuDZA+1Xyz3XxoeplFOEfaNmhOTh+u4I5TRC
wyeZDdNLac9990Q8qKdwt9yWW9xPPIwUy7bFdTpvmgEhfVdF6vo2K5iCptRf4KR6
VzWjPUHJtw7xxy6cYk/atGO77jI2RCkwQE4GAunO4BbiYXvjQS68z+irYhYLjcnp
McAyA8/yOJ9gEiaHASIHGI1MFBj2P3McIeO6KRGQVkEe8y0wqziAvqu5bxpiIVOg
xYPQ/M9ehrOXqC3BrmTdXUYD6O5MleUB5nGsWpyWOUjLZZTepTzwgSwxxzQpAxJC
PZgGAXGwC8Db6kpb4+KM6DWB9SMn4CKgaQXhKyPPtbnfi9geD06dI0bTDwTtYhBW
lQABSh6qal6hItNvQQmpNONbNWUOjrS82zqjTGX7dsNn0Mm7HZj/3rJ56MjcmYlI
IdEKMVNcIquybhGk6bMbGBRYeYFN6m1N0idCxTNE0HM7MQ3OYeG8EJrrdy01iP/F
abtorAMmnMaM33l9/gN9Fr3VYxTW0eZ+Jo9gzmTT4SxRYE38eLoDNgae/yfEUUcH
lSFiPbrMmna89USOhhW31lGuJx6ZP/gYCW00o9Q8uwY9/KSgk/z3qqku4IzDA5VK
kmb+piEsoe81QApw5sE/elOaB0Fu5Bh9xhWekYki9tMyGoZzqz97MQsstrxYyXJB
Mi1chBEA/LOgsi4z772PD/LGxzNuOoTclulhMVKZcQEWZQI41mJtJ21ClMu9S/wW
yfV5a1zj/xNmPC1Ax2GNe2cwyUGHUPgUSOW7XDHiliR7MBewrFMXQlysZNL+asUC
xCVt1wxhkni7GcWhEcmaiY44QmKYpqD4IJoyCaT473HM0l4yjrCqDJPGUj0lonXF
pSkSxgta1ml7ZeM/TsPhUW3/R5Zq3jhkTwYMVsSTiSdwRJslIfe2ygVVfaNVW30E
3VqfpApdcoFonzKaoTe+9XdotxUR3nPIOUE9g0QorG5NKXJX4oePrAZ2fDGlTKh5
4+Fan33mXfF7QVodSMIc++VTD01wMSLgUgXELboPqDiKi/NHN1MZ0LsNLzxdaIV2
3euQUL0u1n+AaDlWD9bZgGlvmQTl3dNYqt8fa0QNwwM2giUieOVU90v0vRXwmXtf
l6Fbe69kOYZIyAY1EAxEBdvHdEjtpw1SYbHmNsof0XwwngR7UHNSZjJtuOPGyZco
vwYfFGXWq1CBE9V3KujqS8/dX+EzWiPw99XwlmXVwOVrfIWbHUPZF6Jg5mzSyndT
OcJl+blDOzCcqv0UbbYUKxWYAQDu41vCCvOlXrZi4A+TORe/fox4WktfHB6zyG/E
7nWXYvM1OTidpUJeYV1NH6qzduMOCsO7dHm9cENcQQY+tTofonu5mpy9V2gNtU5s
mU4fulp5dSKFxtxfJi6e/j8oM3oHr+9eFjtAJwUu4peGgDPfJSxu7KkZf+PDAimP
pjpWdPq7gtONn6rElVU73ezTNlRWruXW7h5gKUy6MK3azokNOUG4MgNJIC6JYKGv
dF86XF9P1zuKDVB9h6CqWPzGtMLxQ1xOenUH3O4/QIvJBAsWM2kVEWcZfUCIopDb
/rsY5zfqcy7Xq9iXCQquG2Vo1JHGylK7Gc/ocSBiPEhZ1YRC46xpm80OVPilhd39
Egiu9fu+8sOeHNOPeqDPAkfuKjXMmJf/k2/V+61E9FJCIjOkKNSqW0aAesnHtGeZ
cO/PwL1sayswximwz5hhIS5T7GnJfz5UpNIz8vpTWWROU/lV7XthhkN9yPw5ufeI
sccXw19CU+DL0qpXRDBaxKvLTUr/nQaQb8oTemsemda6udtB9uxD5MIxiEZRm4V6
hK4D9Y/xGU0xBpPwQSSooX/RfRwcHJgquu3lSBvjgt4lKKI18dVoR1IadLfBLVpB
+TdvhfGkQvv72m4Rjjo1uFyF17O2mSwasft0LQtHEFMp6EoWfsoy8RWBuxJqTXW+
DgchXbKKi8Uu6g06kFs6jcQnK2rLbNreMtrrR+9yzrL1C5skXuncR32vrkFchx8e
fd3tmsdjEqsio0BO0PrnSXOfzJ9D/k6wYAKaeYZ8P5mCO4uS3DPScspvTYjXHVs0
DNUOxABcFiuSlrzFF4c/qXxPDlNBiNIrukRnKXSvWAB3f3aWkH+ON2PFGQLitVhX
7VdT6emIWSpNQ0+sMEafXoeKBKUBciHNcfZfw3LZY+oTq3Wl52s1MO/xC2EpGfhr
Rfwls77a8mlviGMiOJwPL9bW69vZ588XHAT31Dv75otiGGR2BVa6Z6Puk5fl7j7s
wZCAgdxbqwenamQPccZ4WFA0RFvZBfqRMuze3/LkcV0rvcF/rmBwAqKc6nlRT0u5
MvdWpYU5toNDvXVHby7VnfXpYOQnIR6GQfLQ5GuzMM/P+YrjF40OHRyeh8nkQOqj
yV2NEaMXBYh5O/YdXI06goGWaD6vzdWi/qwRBCCBwUP5Kmdrd52NgTfe/oIadw/r
kvHhT/rv1BPsqX/gcsU3aomS3vQdkmCabYv1ZsGXj0KxPmireN5e7g6icx93Oiku
OeYcf52x4a3iV6APR2ZRqf3l6H7CPJMK7R5rqOBn1frJZUZoyNNzh/UNCvS2mz26
Ub72qHr8bSOTa+4V9lHFWPWtBeOgBTcRjVLLDVVSEkPwOTRMe2YhsO4jHWYCgZ9v
sajXk+agZcWiClgH7X6rq4eGCwivVTSlGEpq8l4Wfd2PU2IjRO9iwHG515frbhjr
nrMYnyv4qNgYRGQcWYXlH8UtbNxoKdsmjPab+yc9hnleXz28fozpzDPPycpo6McJ
ogaiTaeGEM5+0e1ze55/3vAGjZXVwRYjfg8l3sPiIqYq0zJK2r59+BYy7HqiyXQs
Gd9uy+haOj1v5+NN2sdifwbgLnJD/lWfxniF0rdNvWGwXKy0SniF8ELi8oapUjON
Jz2gGINZLhhv7Evcdc+xoLYdKxTGybMrwMhe0+hZrgTO3rIbKKo6dK0CJfJwF6LM
I5/iDbU9LPOpsiLnv31GaiN63Xro9S9gUwC0x1yImrQydCKaeW3vo5W+rKMYtXdT
ufFc/OBeJfcbEhOKyEpqGH0vq0Ge73BdoIKIRFxz/wmvbvsg2jOptdTAlM8J/qT6
qJD3lUWoqkwBGmqziEaiuUeGSEP0x1wac9IbHGqxx+j0u18jANRHyhTn82xiXx+B
A0OKhLQdC+ExirqZ0HsQG7PjkYwSE8KgDFJYBmEuL/VGJ6eInWZ07oazbPvLGPPi
BQRMhQCkCAPlkY6zrcIjnoZt5+Za5yzVi52Dj+IJGw1ZhpZxmcDeXmUmgAqKuAxG
XsrPSQTviBklAfmoqZnx65W01UZ7ylhZMNz+vIyOIaDrekyaRPbU2nzzxyeyagZu
hjT0Eg32WqEjhxgiocsgdGlDujT5hwDSBbVXuvuNnLje0udCBiHoSU9k3jCxD8F+
pIqE3T4HnuUVXxTMwoICwdZh+TJMERGxBVgLDL0PtFbMBhd2HkND/YRgPqNO/dCY
C2Dsn0fKku8y6gUkbWLk2vvmqvf7TVJTNDXKkSRqbyQu5CoTa0iigX+TRe3i24z+
BqdUAQxe5hVRyGbo/sJ8YpM5Wt+jVNjl1F1+4uIjMozPdajolDNcupv4FzV13CfU
5vffBuZnVSRxW0g1UCvrxzgVgM6vefjfUYcmfOcSGP5WSIvmWUmMdz0i+VL3Linc
kBlTEFLRKNHURMZE2/IDx9LzHuR6phrfrI0EkjeVhA4EcI8AARQ0CYFcg9EUSN/V
3Kmb8CrxyW6sZRkxzkgPbebg/ZLTZCEUzoPDM4WmP39DPQpR85E43JCpHeIU2eGL
aeDyvsKUZoMs+N0NyrSYGmJLD7bJl7GvJRk+Rr+LVGK3cidRwb08ifisDtrlj6ax
u8N57X6DWxn+/ox2nLfDFaCiOh+bWM9nHGFXKmHdRgRdJSCIWvYE8KRiGBEmpNP9
SQad+sOoeZxte2TyqpOOjQDnqG+kAQZ7ntVeTIbyxgmEQdKiCwOXHxU55ZDHDi4K
n1q1+CmrUuI76FgqR8y8Nz2gy5K5yJjC9zwg+5FzvIwuVvCgOSF/UAygXwQMFP15
sLnGFudHOAT0N2LR7j5K0OnN7pjNwLIWxdyyIZnmWMcJ5/b4TtuJq8h/revf2V7g
5w2qog8AiBO9aEZ3OFcUKf7V6QqbTsAj4AlVHQcA+jI+yzwwK8sSxjpD2AMKyb5q
IhPze4Q6RJMTnV3AeSTNGHoNEl9VFH7FDSHNwz/FwK5DHA+WdJTm1Xhko3GsgR0G
M1nGNTFcUkOfEmz8/IQAx2AqnYON3Jvy5RUYxiTIx8R5URbS9lrZzEqi5q6hvbnF
ime4TCIxb5HdaZ3lUn4LMri+foPumL6T1UsKu4tE61Oxeo0JExywHn4qhlxkSS0a
lkH9f6a6CDAk49YKTgkMbaoXagMBc2dtWK3Xt00/lrZJ4u5A4JXAXdPyupsleA6r
WbSJ6Lw35DXD4BFtyvSFb4BO89I5GD/QWsgVga8XSqwvnYyjMom/bx4sQvWXaBGe
/tkK+Q9/vUw5Knr1zUIFNJgerqqCOMxkJ47qiaFOw5yNwN6iMM4nIi462CCcVvl/
Y2YFLMEhIxYQhJeYhaJ9bvJPpQUkh+Mzu1Qq1GcNWr/UdchX6KXs5WHZTfuciLfP
74nkfTflr7pWJqTBLdwku7pKWCx8Nlpp2DVjxyQE3IO8ZxtvuFmrJ9BhnUbdRlNz
biorv8S7KyGXHKUxAlm+FIfV1OH3zFjdY4aURVQVWxGbRf2r7QmotvUJ1doT5ILb
Min11kaONUnEKcI5IejfQjLNKYRSY7lhVEozkB95+jCODkzTukXdlRtqyw6/xqAD
V28Gfwo99OyeX+tWbYkv9waqaKdWnx9uDEYj+Ul4CVZ25w92SXcKEiGuJmSW0nqU
eIKmWA58zNUs1F1UQFHW3ulTPp+jcWg5jTzydqM5GN8CERqM7zNGagaoihQJxhA0
0U9F+w/rqFYzACqXP/ToOhbiF8XzNQYGBYj/iWMR8GAPqvjUqJD1GYjus3jKwnqT
qQPnElhOYy8vVBL0RqoarLNOHFXuzWfd/NRI2NKjEjEG97hc5wp4JB9jlhSZ4qn5
Mqh+1e+0Ma9bKLkAYv9kUkLLDyXIlE2uc1iqZ1DOeveM+cy7p2/1UuLuzeZ63khd
6lhrbhTuaJfOvuDuYxF6Mq6j1IoEkyCqkbf6Jx0r6JslT05RcTTV19aCttbxXFWf
NV29sf4xiQgPb+wcLiQvExNhEDVhVRU0iSJEzAFA3urNUNMNteU0cs13njt2O1ZR
VwalMIeXQxJNAH7GDexHCS7hJg/FEMP/lwL0NR49SiCcXrGBBIITADzgIYWdQhVz
ZPT+jeZ3qxr0+JQccunPWunn+svnP4pDpWQOqAQVPmEfpexCJccIrbhAbsgXEPFY
ExwpAsXeMF3HexUbkGqDNKTuq8PjeBUQI3dyM7b39FqnjlR86YU76+p8YrorTsvW
j0CNl7s4uC3O/oAPmtYQDke48hZQDyw/jeKRYKHVJGXklzIuN9g0csxmEeRIhcNv
SI0wE6gapZfU0ehtw85A2l4ytCzcdi912OMSx56WUnqVTPle80V4I/gr6lRNrl56
tHCofCeKOn7UtsuTEvTNb0LfwptY2ZkX0W/4c6v9I+tBR9hMV8Kj8SglVmG6Lmjj
tP+AIhputdH1GpngjvUcS9RPllrNGRKCXXZidFGJ0y6gdHH54OxB7PwtfBm+3zfL
j1/rhC0U16iAJiADQOqoxWxQ8naVXfsh5eX8zBlZxvDiz/Nipux50wzA0rB4hMa/
7/Lsn5RsWBs8iRHxzk27VT2M/UjnufitccG9FANcANUqSz8gPgBnb96VgUUYOnr7
bgeYwbKXLJohr0fdN+cgpLcZySzHKFO5bxr4J9eTlmWpfC4cd/EwWCaTQkt7RTyB
3Q3Fbveqd54/77bczwbE09eTIOkp0/FHTXlKPNVarIuIWo6euf8BW+adQ9y+QevV
FEWVBSWSxP+7CRuJTKzLgpwUURWU6ZkwApE9i8tsPB9zUQBEothMhuAGA1Hv44I/
dTbQOwsbKqMaCLh+6lllqGKhbqPFfjysv50bq8k10iaV9Z92xeMzDN26DLsis5BY
jb06occ3m26St9zH6/XQQd/aLpZAO6/xi5ddbwnkzpKVJknJM/Q7mwJa1fgoKYyW
kcX6zu+Y6cmF5ldQw5SA1mRY5t+VgpU65dm4/62ECEXoRjq7dOYPt+YtlVg8gk8v
BzOkXxLjF6pSf8A8Yta5Wg0wsaNixIfp4I74+xSDkAcez3Jya1QrTlXlMRXnEKvK
VGLGWLJcWyWV6vP4OR4bl5kc5C6DiRwEVOtJU4Q+kvnpLTeczBbM7AS2RaKhlCFo
IhREvJaibbRLw9giwJ3tNb51yJRjAAPf2Tyl45O3D2NVK5H0mycqofSudhMQXM1+
RUBm/t1ZNltmpaqp5wraIpmHlJfwrkjMXGqfOz6okZjY1RgT8pk8FcmNQ2RTH/bq
nruVSc/jJ9CK7eGqB8qM70hzT1joM2GYKaFgW4x+dfGdTh/7+ZYhFFaUUCEFNzgw
oFNeOeDVzlyHAh+/kFP19rlhVwBv9CcXLOwQPpuypPXly6Vz/wQ1blvoZQ/fZh2m
33GJn3UGY443NGydSidrzKU8mgQF7HdthlCFn35nu7b8r0rJ+Ns2hNkoc6nIf2y2
s9xrPRWSS+naqXjWsa9NdlKwTMn25WB/1gWGmjDbvjjo6sMsJTzajsnSoHN3tK2t
d++eqloSQ88hNEu5hHNFmdppgLdNogsNaZasDdh1HijfM/xtXHw2CO3WSF28ui+y
3loxqv1V1eYeYstXj4aPb1ryTlGGBPrFKKRK1mnEnwuvfQD2a4AISFXR7fae3mxg
0fnvkvVFgh2StV8mbK3IxMXCCM4HllKfayR0q52T5iuV7Ki54B4v6xg4EBm30wWM
GborcVLStqrcGEaZtToB2vwqjhJB/b4xg9RjMYoBUFy30dr7RrxQWasCF7qBDvpn
w13ZVlUcVvE1H/57/hLh0SCRLtX/UmIEBs8EJ5EmsHKaSdJBuI0NWNQ4+n5CqDXL
aUk6dEQwgyW9Df//GIngAwXSjF5PZKTuJzriqS/jyzyi9d4dzaUE41dxdGHpQBUX
8zEyXyM+duDoBr3SuxeNFlxP3Jn5j3cp03QD9o+i6d+eINPmRUxIVKy7A7QA0w8K
cTFvfoDA0hdN807QxDZjn5B9SGLaztB9gsvPyElscZMGUb/9Z2asr2EHKRUb3wd4
o+k/7IpPJnzErQGoYy28aYOr5czb62VyMw90VXHqVuK+9ZZ5ErV+dqOb1QMlNn2h
bpLZyVX02X8kCAfGOt5vGD46b5XSCYxK+NvhuUnPttbU+TQFNmSB0Z82ywE2PIpi
ijLlCB4kw37/ciJ7KjtyE1LFIwHw52EEmGEtk7sQw0HyEVXgwE1/VJYI5oJMDh2N
1dLnZu7y6lRVgQyKMIkTPPCDS6t6lnbHmhphO0tu0NTX0zF5mGBGAh9e+aNgpiu6
oi+c0Czm09O8/eygB1z1HiOrEcJgg1pAiS3qHXIHRsNcIs+y8V76i8GRj40h9dAX
mRht1uenb4w17SinKY6vh5HGLp8Rs8D9YS7jvwFM4lNk3w3rNelITXwsbK/a5MHJ
KgbvRlhTkkdHDtZhYlWqlZMDOnCW6y5udBwzsMOeKDGQxvZTzmFcZ7ytB0YcXKQv
5gnmOM4nHjkCakQ5trIZ5vhcgJqz7oktHvzvJeCUaBNI1n+VPBUCqeyd7Al6BbWS
TyDtL+d2I1H1jAiLiVY1svp80E76HQ/+cl/DMjkGUk+TKNAqmebhYecC5GfJzgi9
Y3khl9TCxtXrpdy5G7fVSljaFPW/SIcdGgjweCwAqPROr7e2fBc01hrnu+CRspJs
e/+AtgIFJgf0zdlNPNOYeiq/3nFrjnPzn2SMcovN952Xk3S/bCiT1KTWnW0u8x6M
LgFZ+nsj1qeJn+nc0jBYOeuPxkDCtnWROM9I0nLUFDgckRJsaMYpDo7N48Stg0qA
xdmINqEWju5fuVPNbRUXNhOy3C2VMnyYO0pujv5L7Ib4s5EBoFveR+rTlA44J6po
S8aYJHP0UGHwEYq4cbsecqOvth1Byx7zmsDWyoZI0hC5HxRjURGY22vcDYsUc5iV
JscJpWWSicq2OwQhXKL95RJa3wTbKovFd8bLidpcnSYxUgbh7WctMBephNBmO6+M
39wSULRAEAy1+Mg1uv/IW7BLEiUqglqd8pwBIxYGNeaOKmwu9+Ipjq9rq4kbzj32
DzLyB1/rW1S2OAQaRi0ZNh0Tvnv23l0px/fxE1YmA+mH0NOxxPfWk3IH2wzRIQJn
pm0qP8no2aJXn2YhvR151PavKAdXT87VsbTUCmQ56PSpttde+SY7f98ALeY3XSqZ
5H7jgjcurknf4vBG3zwZ2LgZ0GhlLgrh0GRAcyQYObsDQzIB6N/7J22Op96zLvyO
Bppx+o1TljhNEehmEC5ah5lg4zMCMzpzX8vAClY/qsMh6XZ0L/MHlXD91NTjaONj
NeWZpTIhYDHS3js/2Y7XX+sHHz8dJXK2oyh5C8GkoMUyROrmcNoAMk/gvr07zzJd
GsYAlg7WD4nG3Eqc1vwN5hIuIJx4wTL18+CYGQ5RndVKyw3gCrL16Z6znRjUSU29
u9fxsLUVXjB2ahvmg3K5pvFTudx82ZOkBPkA7I/Jv0NZk+hQ1g2d7dyAI0zbiV/F
rJYD8zZC/n0nHg0AThTr6Bf9ASPKNVy5tyArklQYUa/6ge0/EMiX70w5XTY8aetK
mm5k41++rChjik9nxq0SzGhgXgUKRFzxvxhF5brQFRVCuheSPF+63AXwRcJoVY4w
LyoXiFB8aFgBOOI3I0xgIeCu0Z24co5/IDFfoitEi1mcPmoIxGmkLhHpiVGKT2j+
i08kkjD8ipmljKpw33W4s61hstWmjdbFCWXXrXtRFD9NPxK8/lt/IyhabfnOtq8G
XFjoNhzcnm6I4Mr/Jqt6bpREP+7ZSC6/pf1Vcp+2Vq+t5sZeTT8gCdIv9I/bX2gQ
J55BwVqe87QsRLfqCtJ1tg4LsrkxSKsIFxqaWCYKDJ4XNNt9PL6lEB8qOmlNbWYY
PXj4tMQzwZegAp/cOmopxkSZHpy3aUs9YceQzDyWsglzcLFWo6bzrxsgL4sbKz6P
H+u5GHa4PeHaRo7RYGDA3YYg2fxDEKAWAyMe1HvTefh36FJ0tvEiqpvBsGgg+wrp
JLDrS4U53zBB0p6soaFIS1hNVk7nndGne8uUqYjrTD427F1XIgJNrUdc/sqUmrIh
cwlR3R0Gs3Mr1b3Tw8ftJfuJAbAbcMmWZJHMT/VxNSugfwKy4zuZBgHEPbXRmMVI
BIk2UhqFerSuTBRHk1uqAIFuai/CEPVhSRtXgyWXFK1d00Nbc2aVC0FQO2T3y2/F
VQOgsQro9pdgt9AgoKiXIwP9soIJJ8p7LvDaCEJ4ttTREH3h5cbC5oacVqdrf1cw
17VAHBG1GfHy/68eRTFi/AERFluLU6KZvYvBd2WeZlWgVXijR97EXrwJX6fb55Tq
8G9vASJ7+iFh0ZLxrNkj8plzLe5n8x4bGcMRgFk/k2piHVklWf+uFK6nEnOfnMR9
c3ot3ASQRESJ0h7VgOl+bNyw71hKXHbhaT9X/rkp0mB+OlowUhfHGNtj8YhsnnQN
vRSqpxX/XZCmRxUZ19tQw+5tPjhULIxqBBMnxqRQt2YdAJLcMXLZGkzv1PkLYPn9
xaja7yqcdE1a7v8M2ADn81fbK0GOJ5tJM3pt9cu0n/7IvYbfFDbnsSdJ7vDHSj5N
9iFIW9XdM+dxWwA7t5Fhjv8Rg+Jx8Ho+KiDUmnK1l+eiOQLE9/fbvq8F9YPSUi5L
cMeWvkEPoL14Bs2JbXOU+RJr6JkqGxhx5GApnOGxpvs9ozeI70DvFUUNG9oK5C8S
JJTZM6sz9RxMyvdNQPMPDwumUbIfSwop9UPWeE2PoLogFgbP6EXjOiuOQhHRUUxV
5uVG4IDPfPDyYidaUjH3qjc+KEo0yDoZOZ3gK2nfIHIY6RFSeeOrMIa8+OGfW70i
K/EyyIXp+0QyH8Gg4mrz33auCxdj6mNXRl9pXSsnfKO+75GDb6p+DQ9iU528JPJi
6UNxRZ8znnXN2W6tDETWoOScgKoLsQVMtMhCTcbfk3JfTcz0PoDUoDBr3MXfYa76
xiUtKQj3gYW/08YVnNxVf907E/1TBMe9ftlt7G3g31NR1oCPwgS0WJMxFDImuzHg
KUZcXutanJ5ESQLikOWeJd+SATdAIOpj8KeY77bK5WnbkwJSl0SXFpBOx7jfU2Gt
Nf19ROHuzPYsrBpuoL66FRyZAd33tum+2/XXKrTmUmm9rxqZBiqaLiNS267nPFXC
qAr5im1VKeErON4N/zlvT2tub+7Vw8ROJNdt/i/nPPohPBId/I7X8U23voDeQ9Xo
W81zJzjDGLGVXuVybljr5Y/Pq6B8vN8HlKW6PCfQ+lV/8SKwn8eFLe75W8grBlzG
rmCL0PjaLTeid3ssTyG0tZVID2GK0keYRonGD8Teo078mSjmtQLueLmn1tpHo844
3JDWFAxS/y4cYN8Za0p1iRxTXB70g5ytlgnCsZ8PCuhhq86dOp+MCdpegMMEt9ZR
saXpJK6r8CvZUFbWWuvhXJp+EcnN4gIDAUWKRxBdxcc1/wYWBtekRMhQS7btwg6r
JJUL3QfU4BC5DnYQrkfO/ZKg3i6TZSc8HlivR0CoWZUwMERHCJhfu5DT1UZ4rxcW
RIfWQYT4VWzRfSoJin42+q7BiS2xK5SxYxsVh7FBxBwS7VKeK03ZIxAObKBXebDU
c+a3wkBwh0cypfG9TKXAIoVMIhw/Pc9olrNwkJyFx68y24wMLY8mcvyFwovRdK0u
seYK5HUF4BRvO0bKT5QYZ01qCZoSfR0U7yBFkQ11O2f3fi9/NQjiEBwqpVavm8H1
uaVrMVXpE2ubH6tYa9w1Hn3UqrSJsN1Ze81LTH5slCHq58tXozRToF9WP+nG7lEp
kk0tzq41oHjvYZ1E40Lwo3WlzFJhEJrxtaK8WfgXl32K5emz27dWs3BSEdJ0w71X
kJYKd1p2mM7dLnqPlqrZmeLzGSGw281sq42L8By5pfRdsNRK7kkyw7gOR+6kqHfo
//DBlpdnDEgP+FpTegAD09maXPKqYm46gFLHQa7MhmXWv446ZeNCSS8/GB/AbA1y
Q3QepvkVy2/bjqT69SZrkXrYudVScJv0FAkHS+VODFBopHcHsUnguGkm8IKmOqzC
m4T4Dfmi9OsairZwMEhJsXFO50ZNTWd4t9xtanJtIe1loKjaAIGJAlSOLgBpLgvU
O1FTrd+NhbPf8OI+3pdA+RfT0t9o6qy9WGIfEnB6B1NM9Jg/N9df2FdBqFuhq8Wr
HxB3A9//MnlsYrcVN1oaC13VofS5Xs1hBkXFMJVnCMGKhdyAOKZrjAZko2bz3UqT
v59sfVcD4P0aFUxY++AbeNkQr6aoR2Ht0rFTtPdgPi6PVvRSeF2QMP9cbTwS2f7b
smXCuC/ACg2v2S+ksAPGUQ3GNm+yl/1/WDxUO9MqH4GlzCnmKEFg250V5drqxK1F
70nFShI7z/da7xxeAavr72CVut4qFfuHReqMQaaX5L3uS+f/unkAFv8oNU4nGjbD
CImKO1DlKuIi6iwZy/XnB308NcgiTXhs8ZDkPNXHfRoh5MpQUKQqE7vIAhH3DXEG
fBB60Wu9ahlUHleB7HHPOc4GmVy/60n7WuvymvLe1J9soGp2Vi+yXoYAEoGcNeXu
WFmFs4vDjoLCKCrpcpUj88QEA/z+/dynIH7eMfbLmigQmFdS9T4hrdPWm0VMu8zP
7ojvoKYlqpKT6ncTAbf74AfOHJCZp8i1eRGwjgLkjDZQKFvHT/DPaq2dvE+MxBQ+
nFwAmZ0H6oryVOGwKkXYCY+HfzaByYL4qYcPfwc91vrRwgUHYLciDgsZdUKsJaD/
Wic1yRt1/mizFhqmatnaEsvxgelDfGRjYo91BG1vwVEgOEMc2goY6NI7pdeX8AqA
5hcECJOpJ1hFqLkyhPosyB6a9Ona5csNyZdjw7CTzl9g3rwJZ59wHLfT9aIKzaZf
zrZWIqWAQ6zCeUyf3blECtJLbAkw56iF0v7tnQzD/CDFyLEPekdBqyqXgnQ99jhy
K+uwlNwmOVte06KhWZyUtO10RJiPXclpokXTaVvayz1ujhj1QNJnIJEBbQ4NrnrG
+PJnlpATktwr8rbn+2FQUo1P4Gg2Whi2knRhvTqJUBuXgtrpqx79wPHgwY55hBrq
KJtik6U2kKzVNxjhVRVfTjcLjZCH+1FPW0SqqG3xLXn2+p+lKTKW7tC4lOoWXvcr
BcUDX+GRSYwbkwqWsVuva9exQu//8RjYW8ykXGL+a6tlEfU0c0oal4n4NcTIryJ0
lcGWCHV4QXxE7eo955JO3e3+evElg6GEebUVqBiuv1xcGmmOwc2AWpyShFd4zMAQ
5bMNtArchvxs4s54YfvKqriTfZGG0gfO42I//8FY/zKS9/A5bXk+u36ewP1ZfklR
xU4ayyGrO2/8l71WsoeTJg1158mWyiMl9SdN1wngg6NrZzRQMZyvWgjEvkYGcwm8
d6/IdHPz6SYlaM3gFMrE2JdJMIFEb/K5zC78FLwcNNAvC5+LTTVpuwdRiwG0widD
MESE3G3kWBmV5xxZkhMvDbzWlFiuPn0UjIJX16FEKeyochD5c5QyHudpvfjvDqRe
KQzfRoXRcN1Yfdz9XqgtU5tby20n6efXM0f7HXSuFOUr8rjmeZYRkEWZvpu55YcM
ZXZ284JDARP5qTyiT6VuUIvSwX8gvYt/uqmrlFIFgHQnnvj5qQ1GqkYvNmU6vgGR
uhXQhcjzGK566HLCG7aB4s55y3Z/gsh+yjgklbLeXdhr2sg/c6/6z+kPFwQExfNL
mUtx2pvZTtvbEjFsD+zjMJyaZUVsTZGC8RDa4ntIC+5bf1KN7nHDSk0ZfZ5+i6Ev
8Fca0zEF37p6mydTPYQoBLKLid5AqOoeM9fZD5SuzUFLu7eM2llHGK8VT1Z0HuiR
0+rHVF3FjyFyj8/Hc7GEB7NBnuwcJ0tuiT49vIuUQPFG9jQc3F5CHPArijPuWcln
a0BV6UdN/VuymnUloRPhjv1VxxQTfPTXxPmIJ8mKaj5VCuqok9o1HzpE7BTlF1Sw
7IAwFbBEiEA13dK6//OAyjYN/7iNoBIfdPA+bgf6LdqcIDoAPp2r9AzC1eLE+GPe
edj9J5Ewgu0iXqngpz3YZsrihL8fTcpL+qZvMmKXBYyfe2JHBdUQmqR9jngC0caa
wNviOYWlUD+dDZoMv+Ief/oQ9zcU98wFad0qNbEeWvyiJiOodIi4o624yCKxqVed
iT+d6NbWV6oSbXOlKQn32devjDObMgXyw+u+J+PSMTdYPdY4kEeqwtBVqI+A4WAm
o0dXZY5fk4na/xnM4xbaWUos7L8ewMdAMGJTEVzTe3zP6hQfMRl95As5Y3enmvRC
zM9pPzfD0r3US/XoAIQbLFVh8GZ1Rg83KhR6XCV9oFI5M2GqcDpLcY7V8WuJiBPZ
/WPMRWatYiBKn5Wy+R/QxkTjLLikpz9skWm3TKQ8xiyuaYuSFaCQlEhb2z97CkER
GTfthYaCkIm+7nfGCJUNQFsIEuuZ75DsqU8YRQFb9Hq1GCJdsjAwyxYnDwjeFvia
xcD0L8Xmb4LRXRp/6H84daHGPjRNXTY7TUwNNcwx1BHYbG35DNAjYyDFBrzxeNiO
hGhmdadecsxywEygtPzm/wdqriveC2xdjfMMQBCUexubsE1DfBb43MNB028dx4e2
ZJrM+Wh99MPuNQ+puyq0sbta668pGXNoRZb4Sn1sev6g9vZqnuecOJPNnnC8SQsB
H7a83NKosLM3w7GiU7hGsWGUYVXeLpu0HHIMcaREpVYOytFquQtfLNjKTWc5G3un
eEdDFbEl+2VUlNuY3/s2W9+XKwawHTgYdofwPt9xd2Y/VePjwW5Eq4gTU0vA8oSs
AR9ke0MNe/HXF53UgaUK/Fg7m4v4bsQlYIU37rwrg6rG5N5pzn8vhWRkcxrIb4ac
gjCn8jFaVX13UTHKhysFnr4yBrFm7pd++X8cR+nWRRdMT6eRcl9/J6tAZn6NAoxQ
DRdCh8JeYp4XLqhP0LhXvb2ixkyihavSWTZm51blyjOfgmp01P+cljSe4fCq6lHa
LFyb9EkIeI+T+xWtYyWUlO5tNrauEVNGQZvOoCet8f3KWbMt1agg27fXwa/YRJj6
lKPC2dHkozygbSpmsxmq1z7Zw+v0bdeue4oW3U5Ac0GmvN/4cUEL4jeB66MXE5gv
+J0AwCICDIPsFQ1AmPPqIeGd0EKIg7mv2JaJx4G7a7YilzSCIITzVWOWiAqFqevQ
04a2f9ShEL+pEmgatZMJCOFmuxxhUN+nXsFW1kqa+Gyloq+LAsdrrRJhTPgyxkv/
o+/yVVw/FipQp4F7ayGHnfrFfm+FbzPR9XwMCcZCHGYSi8+c5RRYroe7Bo+UTeEq
NpR108qlQO9RI7rm8S+Fn859JGyg0b9nzi4eIeOoUZOGrxTyLmGGnpVfNDDKeyro
lzGbM3rTz6/lEmJTMXKISdAMMh2/yeB4Yvppl3tKiTUgZ94OJR0SNXZhjNTa7POo
fjtn3NoZ+xlpmXTHvMnWftUeUQ6tVnVIQIuWlOcGBlq0w0Y1x8nlK/e8FHS3fUdD
jCvseCjy5NPQrHKRhKtQR3W791zd+hkK4OogTTzdkaF41TSY5X7CSqFWjXeoUIgl
R8X3boR9ymGNF6+X/cJ5Zb5gShUCGmLZ89KeQAAKQxTVskJDkWsDM2UlIuM4YHgY
O1NHd38e0SUHWklS3cu+VpQy/s2fDY7phpuNIwzxTi7xBCBhySfhDgopfcgmzZjT
Ai1nfwKloy4phbKbt/CHly9Kd3/DUanoRczAf2CT+3ovK8H3AQkpbzqCoauGLtan
Rj8ZFgAGpakhNp+gGTXJ1vGZcv1QH/Y5OvOwA8QsNKOjOavggkcM6fOXPbq0f540
l+zf7C2IQxbZlnajMMCyLV7xOyQY556nbaIaO+KtYeS9qyEINtCgO09CqXrRyo/m
qnStPDtNPj96C7QCJXpjT9JpuCb3gRxSCqlf5C24jJPhr++W27IB7t0xmwulN/Bn
6cG0b0bwb9GGUEFzrit6Haz67eB8cabHHrMeAUIKxi4voyV4ZbPj7r74FmiKzCIE
YQatPFA6Tfc04XAaPePd+OvgEPfksqBgVWaV2xMxmbGxXqdX/T2/nIquUvodJyFw
nOiQ25/TJxY/UadNCN79V2URgRjo8fcsqEXNfOOAj/7Rex8JHdSlh99zU42Rk3w2
0WINFopWd+pQ1YUWfQ+Snujl9qLz8B14xOtTKBMitR6+6uL7FXcKnw00r1tGxYRz
svcFGtWxrmPWllb2TE+hWtUAb5yuaUgq9KXJ6Rbsox6Ki7jwr7FwuKq2Cnl33Eg+
Z7gq9vTCl+RXx2V4dtpGdnadgSxOCb8a8OU2FuBCID02bJbBfHw7o2noYHKwc5RG
AwKVr+cfAoCWq38inM8T1f74tZvLOMjkJSY/jKe2QGDouqcFUkMyqDVBxb7wdfmj
pxBJI/SkEO3adn1Bb6N2t15kj0M+mDUGFXhT9ltg6OduVwj78U0b3WQsazvFTM1f
untoXNnSinDk19S3EKjrd3RDH1dowIn8SX3ij+32qnuKx4cgXtQHK3fUvM3Tgwxg
g07HQnNIhd+z4/gQ1jPcXfsplI/Ll8AGhlGMbJDCZIWRNSZDvbq4pGrpiuF8b6KB
Ki1qyIhpWNnqYqpPXesfyejDwW0FpABCVpdg2D6rBujXxcKZWPbFZpxtahwZRgPP
t5nmjpv16gZqyDot6hiuHd0yggVrEbwhqxiCAVmBuiNGBp73RUGPUbY0CXESP38r
RFk29NbI4vUYuuPn3QVkAun1Li/dAR7xQZnLpl0xHqt+7zGqEkSVDB0WCX372Lmc
tgXCHw6YfKJfrbY1ODzpBpV2eRUS+UvmbfgzUchSDdbaDcfz2MsCsCpi0LZRYf0g
QXCW+E8M6lk3O759sHc8mlNZ2WMnyH+a373zfN078aIeZIbfC3eAA5pEMs+DwYhr
aP5ScbWkHQHQlwrgFjWYbstySvCiu7q6Y3B54PQGdbGXlMUsEqMMQFttPLuJSAlE
ry4tT+nY3ygws860b6whWGPLRDUyjrgCh+7S24fUYW8Bv6dqQY7rOepkjOZBbI3g
8jTeIq3vCSo4d1rjOgbwplUmFNzihhCGYYodOK8cpX+n+S8miwJZ1fGcQtQYpoP7
oTglrQSZywaKHFNGThf3INMSGjLgjiADRjdFSqp1GyUn72mSRleUrZHSezJ4ivWQ
UuDY0Pbq07bWO0DAgvdPZ00ZJ9ZokuqDgCeftWBXBsLXXxWVkL1MIPywBy4A7pYY
8Un8++e1vqOToNBdJUwULIk/MEzsjK5l3mPgPh8us065C5WpJJAmgPIjjineP2vr
9sVEynZGXTCTRwdnprANOO5GI/J4AAs/NDvFLlyeIiPz+EPGnZYgUnBo9/NEJuoq
kxVb1KHoUCFFdJikZd/NeziMORHbp8UsDaHLz+v/U4nh3HOygkmMB3wFa43T4e1H
y14hldBf/M4UcpYcm6kM/KALCdlBOU/BHVQkgpAgJr2pCbvdSaorCiji8u4qAT/z
fPYHOd7xTsxU+9GmWdJgIQSNsmq8FfmAvK0C84DuTjDJEFlPj3+BxSXk+DsHZOO7
7l6cr3O+VInHtXyBwxY10a6RHBm8mG80toD2a+7MDVninEriIzvLFF2WDs7pJriD
IoWventT2F0MfYbwpZ73397XWa5tfR8fDXW0V1JCIGo5H2ylhprHb6nDDMu34Nn1
F2L4PSnEEdFXEXu9xsskmPi89AlBbibh/hlJjmTfYJ3HMf1QxJ4u1EClr03nGs4g
vV/nCepxvNgayTGAKlKTEPZeFV1WM1bCetsDsSjHL83djq+OmZGlndZHINVgo9Ew
H8iM+Q9fJD8Ca5ERt6pxBGfKRW+epMlik+anRFqYm5n1X4LERnz7auH4kDowjdx1
Sr+CrPPp+Um3AiPSl8Bvcp7HW7EKA3mTxm81B8hyEHXbAKAYltGWMrEH0rhI+dXE
SY/llIegOqpZuJl0QfkWnau8ETIhC6e5x8fnyCBsrLVpMVonFL4I0tpokZKCGtr0
izr6vt0aR8MTpomK5QqY2dbryrIavMWq86IclM4IKQCCrbn+gEqGGk7vMzXopepz
5I3YBADptvTeclgIZ2JIJZ3FEi2eYxEuxa/oGyBouYlAy9XW8633UI++NGTwpkwN
E6qZzP86iLLmhKdiNg7z5dKOVjG/JQLDpG1lHoBD1nkX0WinRpOiqt24WCnEEZXF
E3oDeqL98uq1cwmsTomp4YNny1x5DO91OKA2NQLNwAXaac4jcrOXveIVvG/Zsmx/
4a/nRwrPNGnsToSO/GZ8pqljRwr1pio7EoaaUpCbb1odlyJBbQ3JNOFQNFifMlqY
noziBdxrgyE3UKW/SdyhJbRE63U3pt7dwX2cUJ2zXZm9DheC3QY1hP9NZAHlYa0j
Y6uhKsHwVCUVjhEKYj17xjgfkSeTHRHiMrLWLcOXHvFq0ZQZsOFSYc9FmMtZ5rkf
43C3H9DM8pk5eaAVSmCtC/nM0amqhLFTvnVlA2siKSQE5001WP9V9s8+ZT1wSqxg
2DQzbg6nkc/jJ5QZBs+YTHrxX8vJKC/7UUWMd59zXwI2TSUSEohunsFYv4KUF0D4
JxCPypU9xk6wXp9bE+WpyZ11eSYCxzZAWp7DvbDre17m41q6KxTx8qB2w1ohW4Fh
TJiQ/8sIm+sJtijSQv99Su+JFFNEMCYhIbm4MZcpZ+Gtxea4+H0jA9xumfQTNXKN
Qpr0kxgjXpystryVe28OCvBX3+beeHtQv1R7PfdclOborbo/Ol0Waa31E2V5V2eQ
Hcvxddi6swKdgWFumnBtcIxe6g/68FwCPJAkkrPB3qVsY2xg3C2qKRtW+m2Z+p3a
A4M6DS1QN5VepWoh6b2kdsev2slFY+uX5LHgCZ4ZzXkHYhH6obNK1/8oQYzxl6xN
InQbwf//kwcJC3VpRAc7huBTz/3f3iY7XK74xIMfFPBTyOzTYDp5KkxHJ0axvnwC
p8CAEjcHq2/C37EY17oaSpsz1Bb40HHnXRXUwddXp7ZEWJljVQov8vGtA/F2sHWq
ak80U0I/CZaZFzgNhKvucsx0whhouC7wRq/IsCw0aVf4wB+SkDeLa7R6E8DyB+4Q
sZAnAr0tUrPG3wZicujA3qL2+3DbeGUt/0EgVySo9tNx8z8L2sRr4yPmwl+fuFBm
MH3QJqW7JH//Bn+SK9ZRTfMNg9lJfNPMOo8ughXg3n746xQS5OqQvl9xK/sqcAJm
P9hbMp1q/OEyuwuMg3hVmMGkc5ixc/hX02uTEpn6mfc18nvc17lu6OJ38IIkTjxw
56Dbngr864KZoXBNEEBkCrdrqdel8K4cOoVeuLpcIJooOU2SV5hCIii9wwGQGRYP
nWSTiZastBAgo04TLYQUN8mX7eYuIctV25SRFXUqE+cQVcItNLyzZTiJM1tovux+
Fx7I5r9NvUmv+2lsappdxwSLjJ4m0xsSjYd/mOFA/AhhdNyg4vhksYQV46hKVn0D
QKvLv6B+JpqEdkKM5c1jipfVR1wQO185e3R6HehzX0hIJ8GbHa2zdE3oKCpQC8BN
p+e1ZvF4CWd8eJDtf2TTUC8vf+S4QQW49CaDSSzWoNbP7jVe0N3vSAHl/QpBiM+G
/JOsgB1Obm3VxIRb0xfV9FTqsJTF1Hz75KVXfQx+YcmI57jJv27j2JUBMgJ3AxVQ
/mb51Yhb2F66rmvZLfcClVMGWLGgtiHPQNHJtiuQAaMaOxWLU5L7nQROsJZE7CBl
7yUL0N5vrjK6fwARwDnjw+kbIxvh6hlMYqX7yydJB+Wd+e3TbCSzMPuQ7ighkXfM
vjkOyIpgmbxb/2pWKPguEV7zwz2rPmzQMPqhb25cJOSGNBDrw+JKBZUsXy5cuzns
0aBMR4bNS4bgvSEKvwjKidfmROzBTETZEA+QOUd+bKsSMT2m2ay7hYN+GTvgaHNV
a1srE4RAYHjm7q+EA1nVZ3nkP1X1ec5g8g75+bmoBFiAITrdeMIP9IGRj2Azhdpj
yfVhqZydRtdp2Hjjea0CQq45wED0/FLmGxylgSbKqXNNsqqTA+3BFElWAk+R+rGL
IOnXB6cCXGBLagGR3rBOYmTIK8fit6bWA5Afi+EZHWgA/VTFO8tmE+Df+gucZIPu
CuYgvlMpfmXz39WNitzmAzBtW659qVMocREKo/J2K+n/Tx6TCatHYgrmBVrrJGc7
C4PygUBoCB5pd+GcGoTAjeOqnKzPAjBR+9yBIa2pNn694QZgP0IUpZaTlJIwwsHK
udQljZvsolmbEZj/lOy2wPtgb5W2kd5JgARchcYBUvH/g+cR+sSobS8S1hyZivba
8Qf5Q0FXj1/oM0tjV4B4A3vmmKVO4VSU/jaiciIXF4o+3Fp1aZ8aHGrwm69roOld
LOSCekoVeo43V65eNqH5PGrr7yyC92Y2xoiDpcvQc5vXLSD/riBa3L86JX7hXSwu
tMPWUCVUBU5YSf8eEvBSifkRUMRU9ViZh2xfM+YnHfjD1PfjF2GKX5rXx5NYdXoF
lZVRxGwokQiSXozcD8uYz+TkvGFYP3QZja9AIqJZ02djb/7gVGd1Xd2o0mMcDQQy
yyh0qAQmmi99SbzGXltiNi/zOSGHVdZsbw5WmkZ4mAie9fX669AReRJs/d2TVJxE
oHcm0b2QLR9u42cZ/RXGHpIUMJJLAuCMRLv7qsxL3YRNAcsWeChFqz+Zu87tboSv
iFjUXeUciHmO+d5vFzFxp2OckWFrFE697K1zhiPE01ljb4HSfLUElrwSlZynQhH5
30xgCuchw5/vFydiPiJjE38znlnQCp5grzRsFXP5RTpLFQVY1FO8BJsnT/eBRjNT
GETVO6XC3wDDigv5NT9adz44bciuCbOqVSNg+WhEERQhQmpx7rh2wXICrBqM/WUd
WvYfHLXlOre0lzJEWoolqhSOCBTgsqEkUqQ6oinGx42kAfE/hKO5/jCljjpMk2CY
FrkkqoT6pge0YD6B0eP+ceNkBbai+3V40b43zhMREX8KeWeewOui0kSgVjMJA0vE
4RKJacoAheYEBp/7fFo7ul+j2ANArLvxjLel1abI+6k70I2sH7XHDpGc+9iIG0iU
AnSzF5hnuKidwI/Nx+5IIeUNKUthVSJP6F3cLo1HZH+OK+x64eqB84GwWTv0aa7c
aXP8tCLMFehVImfwvPffXyZfqgZTOLD4D8UCGyB0W1YY/7ITvVV/2q3oj/P76jws
Gaqp29AEaoW/iaq8lbxYrJ1PMYYuBTDTHdV/T4oYq+UJPCJqc3U3pNU8yDgq23FC
poSkkfAkJQJPAjXO7fCNXbKMTKd0vz/rXcGyZryejr8JllphczjBm+9mwOU54EDz
5G4Pt7rftdnq76uE1fwnfvqY55f1O6dSLpOnGWUE9o/mtyv6KLjH9H7wBrZR5pbs
O02a7ewRlYlYjjuVeRmlBTmmid+UqlsSM8P7Dogkgtgynz0RmTeWFW/xZ86dzyjQ
QSHNpazTELCHiK7m+sYUgf0IRXpT+45f31aqNA2bt4ic2EcAcobZHrUDXMRARIks
Ffm9onV8NDEjlMvGmMOWIuInwJjSY5eR9t7IMtn/eXus1gtcSwZ0TndwI4aoeOEy
lJbzGAT/0bbSSuqw0EkOnECOP1nPoW2K/bk8lfV6GjSakcDlOoOtwfg+EehBtnWo
4Uf+dNL3h3bZCPFdU+PIf4goyT5zhmvVyCg3A6FvmiZd+MKO8wBiVvlICbp136QI
OHRX41/N4R4pivOkBoQ5ep/+ydYNwT02PXhLaclw4edTVUOLTqcnuAeTYiKCNQn1
hs1Df4fr3vDO/vfmUOiocZAG/ssJEp568i9GlDb0MheZg1ty1UFaUHX2754766F2
UTEpHiQGZYtavycKubK5yepBHvYo7b4tkwDqzxxX2+zJBe/IsDeq4WluqyMJjVD5
axoF3wiv2cT5yY6VfogrSIcmFnPeX/8cFtZ5fFmb7Ig4WDiT2AOGFXjaWt8x1y+W
Go+/QinW7HoKbIWSoV/nWF/vWFckXcUkABvNiAmbo78sWKfnriG3q9ETS51xrNdJ
MmMbRy88MFmsPaF+Wx74g+yLg2QA6Z1UQYy+4donQdVcn35ULrxWl0rgRHGcplCc
GNyAZs1crDhdLzWMae6upS4Wex15doiJIOLlssWk1pRjNPwQDLN6w3+k1RRqdznQ
YiHQxjOEfS/bEmcL/10tq4K4Z60oemAuYcBSUNS7sduNnmOnrPHMcCwtaik6mk4d
VPH6E1ePuaTDZC7FDyfyHlDw4y5vVEquYXeMCVP1VqnYsr8U6HXnHBFJAVNbOAkB
eUTjvn3Z3Wo6DZRfCJXgQjJGLTN0rwQ7F+9/tf9yjReZ6KVkxhLodN5+YGATNY61
MnNBIwTeDu6Pr5tM/AuhDJ7ul3cMtpS9gKQszM5zW7PGGKmUWynegPNLPVcI3wmP
jndHO3seHHZNAY7P0i10ycZJXqCzed9da2+bYOmk8MOzLPCL2TARWXdx7spGfcgZ
KHOJyPjeGQrOLbkcRyvremrhlt9sbFht/hmdb3tVhMlGclulEM+WoTEir1KxThhP
2n3p1SvZSTSzplTpJaOGu7drYJuGJvP595y7OOkzSsDOKy6wEcvgqOtT2XLMSZCg
zvz8vcFulvopzosAd5FktSZUir0s1H9Yi8218aJQfeO2Jp1HI/6EoGugIMz0VNNu
zksS9Ren6J7O2b8YIS53DRjpaw3HqqXgXapqmv35vfcNkuMFxWwKeiJszAi7R9Nd
tcxeW7o1cQRVGaE7d6dFJLvXdszqJpBPrzszv0DleuxPCi/O3S7JST5FwCx6Ttqg
DFJYItKafabSNH3/ylFxpskI2TLxMO0cVKs7G2aFi0mdnaLzYTcWJco+hTiZlmpf
1qw4CWJ7wGrhHu1Saju5I1dubTjWfICFewirHNI+EbzKZxEh2LvSCY0swJmAZ6Mx
lQ8F3HAbViNW3b1b2KbFId8v3oOug4fk08c8XHKPK3ofwpR/Wg7hNzly3gA0xj+e
De88f3nNgiy06LSWtZ+V7H6ggUXDmKkW81imIw1NKmNGKhgRnT1cDLgkkSXkzmVS
FDCNcebPkRI85l9PX6ELOuZv0FwjQg1mdOdMKkbzRbv0GyNSw2L1iU3SCbew5E1G
ndm1BNevHgLrBfyYOVs5RAhDNd1DtLYJqRkZUC8WrjwymO+d0MHFg/SqelnOOkwK
GZlqgxYD9BgXxTr4u+Pot7QwkHw+pIk5kpS2WVr4nwmMKDtqvXZb7HK6VMUY3PyO
8xugyhuw60YZsszdOPoSQUYXvkKUIkjJYzsf2pjuLWJdi0xHEx81oSHyZJaC2hnV
XP7uqDdxYUvleFDg2I3F8vYTLVsAz/CyVNHL1mS1qBSRYEKwqnrtv5hm0Ts/abgV
yRLBV0YV44SqeD2v7kBHYjneUkvADUByhXDdek4POrD5w47G2pXSLR+R5VMsoF3L
EU3XqweLzVIzidd3yql2Hg==
`pragma protect end_protected
