// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:34 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
H/2zQnpwYcU/dVLJXu3fIc3YjmFL7c0WSguyU3rlC9hyBR2EnJh36mDoOe0zHQVH
P2N1csYAMXsiwS+SzACNAKNBs0GJd9mGCsNuDw8Czagvak89UGNAxUyzLsa3JaPr
jL/5BQ30jKx26BcGKvSU4wuyx6PxjMzKY+DIq4HvTsc=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 8224)
8dGmf35Uq95wCiZz3FX9pmKTBwPjEnbruCT4le5dZLvpzemxblpwSMOcGm7XPefK
1TXogqVFmxEg30H6mYVkN/ppcbibf/vKNSOFlFYpDSPm4N/X9YbVnWRoJep8vE+C
ltVzpyRR8pak9Tqa/wJ/aZe6pgXlWKtBU5slWxSvPtMLlZl8wrSmZIxRPEd7QAqr
Ihcxnv+MZwwVer6ftNzqnOCpCOKqkXSr+h3+adULVxZAoA4vWv1sUUxsuKvXuGyQ
v7QPORni9xWgRJLs9BLZFdllCA8a0zdAEU68vQZPfB3XHtC/sdEXbAS8RoIKJQJw
8P5Ps4Q9MLjZBmxS7MX3KdnJsrYzu2kjQRnbogAbFBy8Oz++fp3f1awQpyvUj3Wi
x+JVXwlB3YyFT+juqK2M6gHLxbb2O+Qtalt4yjSWzJdiN/usSmE+G/7sr4QK5ozm
rKyTOiOPy/mSNaEgnAyDfcs1khIpRrsMyfY7A1VX4VlFMV8Q3+/Ebg4ZL8Uwup1Q
NoP46U4v3pcXNKVAvPlIqQUWA1MrQQzzQ5wwxVZN8XmNqpCvfyLCF584agREMcO+
gxy8ynH7WtLD6W46p2v58W3l5aV7WJFVzE7DZjWLsmT/D9jyUZ7kT/EjXs7zViWi
jG8+aDIy3gVgWUs6sbG9kopYUijwRSY5kYdgPVrao+XN7uVN85Gg3QGIKo31quB/
dQvSaJeKKZGsx7hf5KO1wffz+hqOOPYnPjJUuKWxX8F1egCSXqQQjt0kINM4c47Z
Mw0wHfBt+oqQuJDhoyBZZFipIW9YEA7JZ8U8rAYZwPFg4kFI+MXmsS1wFwiRt4JK
tX6PoPKmF+RSRfMC15M6ZjYxJcHsPCGQEbU+pw4Mgstk01BAAufCktQcTVFrGqP1
EUZhrW5sPObP3sXGdl/Zu82EMgYd02prL5Svif4FxtJ+/wqwVEt8c6OKc/rHxpUJ
G+u88kjVgGIAl6T4jgiETex/0PhjqRFkDF+j7jDPvSznRJ+Z2j8b/Tll+CDrSN2x
VDvE09jLALThvNwKoTCHq0hJCr9exddO04yPAfbLvsIroSPitKFOXOPnwoIsCnRU
99BmWtXL/VMPXjKUWZHX/mZZIbT/7ZizYrZ02tGAsODFUkoG+0MH6SRdhtkXuW65
ZkVmw4CsmI6kHL9v8abNPlc2UyMQ+QoiPaYdh55JmrCaFjDUm8y2mLnnc4iHJGv7
S0HKTUyJnoG+jHNjS+UsmpucqV1QcvYT0ywhM8O9C10X2POTdrxvYHPxPIb4da3C
fHfEnfpJ0AxZIdRaThnMGYBkbmGYrzi9fJaJEchmcY2zQp8BH8ArMspU8CB+lfY7
iU4W7rq0gyR+YFUV1QlY2UH8MZ7/3DdrE/nxP4POK8sno15KYfuPdbvL9xUzzgxM
U1eJtgvCsJn+Il6gWyExefk+XvW9n37eO7Jw6jSTbfsZ/G0OvmmTywYxbLUANhdx
CZnTotNAE5OXC8keo7b/mL2YSjg5Y+9AvtRy3gcL0w/PwXvlu6ntOu3XynfbrbcE
JnlZeoG+8fqXFP8fSutcUxFDteH+QQvcRiEPu3xSvyHr9jZ1E2kJWo941UjXBcIH
XkZ21uy5lDkAwwswLK9GA2ExmPbv7Uc5WRHQcNrgjVMfv9T1/VYKAhwheeHIcx/z
ma3mk69LA+qzB6FqwVTEryRUUcvu1wRWXXkDOzhEadYAS4Ov0fdZvlT2kRPvq46P
a6+40qcDRA0FvAzFw6PgFUzSgYe52M3w/zphyqqM8FcMbwwT1bt+FTV3uf4EIFho
l+3FdH0Z3akiEOE9M1a+ep4Sf7RslBC5drVIQSjVTadmlu5zhu2ZjLMkDHgCar2v
wFA+ikzn6wsHh7ubfXY59ccVbb1NUlwaP89KTwbZyqW+19rKguCsoESKTsenlEZp
UUU8Ds7AigMySyWXPd3eAf2HGh7uLGzxEScO2J6WAQgbkrV7MBMi7UOqpLiOLfwn
9uTSfodBcbpyC6U476qSQjXWKKxOqGLuLHbUUtucsq3ZJ3SaF/J310scA6KBqNdW
h915ccUqGuiPOAV4LQ/0SlK2usyO0Tr9jxFUAaMqMPJQZCHVevlarh/TwgtoJ/3E
Z+gUzRX0uNpAv1Hlzui572mQ6Xe+LahG6Idg2EXAvIst3VxuaH8vIWZUMOZfJ7FI
Lzzkd6x2jvDc9fXwcXl9y7BSa6R6uhfFBAgav+XvhpLXOA7VSdyXZv7mKKQB6XRa
lUYkhp44owsWs3D/ft9ETawcLg02L8OMa936V/zq5BrFJ+y221VfrO5GDyhXvNX0
obT6gVjYeK5r/9RqdhvfmjNbCamqNA4Xd4QeKnHGongc1g1ey3oVV75ohu/JOAOB
a4pidPE/jbj3b8Ik685yajmIfB/EFVrl/XBqT4OlAZCAOO2/p7JSHnUi3y4IoLhG
0U1BqH2+nypUTyx1yhQSDsGfj1XQJV4B5vluDOWXV3upX840ItwI6wR2w46Vt5yc
DZRgpErmazoi7nySfMLUpsIpMZwvrwcbnsWeDjDPZviGHdBK/AS9pXEhKrOi6kVM
D1tZCrg98IkchKWWTG2aUzrw4X47L9PizKD2IyAIvb7/f2SsCSu58MuN2E19vIbq
H3uUzclhjfo0eJ1be46TOfCiPtvHxd8mLZbmolGbLgwMtLfN+ur+T0+2+GvwK3a8
PQocOG8GnsYJT6J9tXhcz19fUSIAdFwBg1AqMWNIyu2+NJqRXmUwwkl1DZ3q9kqz
0Y8syp+L12INd82WOyU7dpxffbXd1CFN0Zo73d2u2HjDcPPGJcOUXv5FU90+08iN
PKGqVRqxuvzIBM+hjp5UajotdtN0nsGuud89DXONTdaihwz1aujtE8HgdAonLNEB
ROC6L4jJSLbaKedO1oMIV9DXXtWdKZ8Abc+ALEsJUM+m8Emb5rGtCPXzo72pxAXP
PBuf8ZKmtAs1xLtpxHHm/TK9OewR95daZZPcrhj6GgGBTGtUQU6rn9R+MrltqoIx
KMn5Bpl0E4Gh7vtt2Ge9Nv+T5oCnaJgNtwpQv5GxVvB8vkdMXcPsmMfQBjO8ZDC0
KZF48J+Qr94d2FAzCpLNoi54kWULYCCDJpHif0VAUGFwqL45oHEVw63DRau5YL+0
m2ccR1mIxN5fydCXSDyXECCA1fOEcfaUrxjYuYWTjB9V3VDaivpZEIrqQHbRHxZK
IIc2NLnoOr3Y9BowrCMsUl7DI9i9h4ltnul9fWzJTX/pSOiWklP+LkQUVsoPr+Z/
RBWEmS2DFHvZLywUHGA3rGiNbn+rjVKXio1krgkVkakkhZNrX1MMJuayfF8wBmEi
aUlT+dmDJE6azL8Wvg7keRFR9cEuQ/BkLWVvxoBlPQSfgY19D1nxDgS+Ei5EXyHc
9/NVASgYB+Tr6cx+3vG24GyOm4b4+ILXjXiKiNBSzUfFVxnv7QGAseWRXjjeY3pV
gD7tVy7ORusXA5moRUali/qirYZ9h5msnThPZsHQFzqfLpSKQSzxW6KvqKRqV3Ep
06LdFy5eFwuJBAOo+9nV7jufiZcjAMA8iR/3pAzUDe8IPObQE+wWqm+FEmiRiWCs
NnvRRTVcnATlfwMB/pKcUfCyCN90uhZFI8eWipLGUp6y/DdmN2WL8Zz8IaLyS381
n25gFwbR1WPfVAripbFIsxlc8aXqaqi02fKxgAvuLSlr6Xc+GpmXXUS15obgHHdW
B2Cfell2q8gPM1/3yKmBxaZ8zVVXYaQd//S39q9CXgU3ibAdLMjsZITBYuTVsYvE
q38FLhv/dB0iPBhSNAMvLrdbGKAmwFEONKiWED+fuf7gOsmTvVPA2Td6M0ngrTZ7
tdnYKlQyhZZ+SVw3kXOZj3Ctk1hXJbpI4IlnzKFVQGrNhBuz7PHgN78aQoWyiU58
oVxrrbkRN3bXaBtCreSN8DRNKBAYIQcwF6ynErTnrJdZpc2Zvd98RWoJBeZNvfec
B5OWWv1irDafN6g5En7WfIeFc7O+j42MtFmvPC5E3y73nwYyeGDjF5fw9BbpFQft
Sw/HwUvgRiXY09duzncVoWDzJujdbDQfcptlzgGjmTvLWNebslZ1IL8POeO6Ztb+
tLNeHkD5taUpcYnQOMWLYa75qYQHUdYSliFkHFZDRamtXFtp8/dnpiJ/RKZlLIJ+
V5jnXvrJddX3210lXpb+wcYhG0maYtH9PQAOnb3GDh4zOqYAo7DxEmTD6SZtDm6C
eRrBZHI6p93OOIiY/WWxWYtq3sq+xCz9iokpttMMW4qTg72doCRWmaplqsza1i7N
GAh4pwcC3fkc8uKnu0l3lOlxn1rdnmd/6BaWOvB5NRhfP+1iUkIREMduq4o/Sx8J
TWGU0vyTtczYHAnhGRQKq3Bof66S+FSLdUdnw/G034KxAtLWN+f8g4JWd+AL7Q+j
pD2XHqy5j9mWeMjXDoWHbI49JX8E88Y5chtq9682CAKXAJ/SK3BEQvXNT4NZcg1m
FzUZ+X7zj8wh8AxG6seAZHzT0cCiWpBrkCzUb2QD7R5SZgPOP7rhS5M1OmDkQgie
3rVQz3IHR9cPxErwUhv9q6ddazPo2E/V6JR9cVVKrvDr62lT1M7hA5iU7jpJGfwA
4qC46ZlJ7tNoupwstEY/YuQEd3PZuF9IZLRU6aDCGeImsr0LrKDZuRuVWO5K9anv
IU9cuvWLQtmC8bGBqHbE7mM1MFouK5UNqUHTqKCT/IGnTm7NQc3yBsQBTbUCrGgz
JsmdCBXPhaPG8+yUsydB3/JM4x87cn1+FMOwHOVzC46TocV+Kzbqu06mjmVoHLhs
nj5h99psJ0IThvje1PLpYxzp/U6rI5rv8qTsl1hkeiBkVl27FRrLuT1o/Ky0C2Ky
w3nnxbKPKPJeWY05VhJAD+tOo8gO6qxpm5Q6kuSqlbnyujN1qPPn4dBcFBNidoCr
Thr39KEWRRlaGUjJoPoPVCg/uOAlFWJrH+jKVaY2QbyUlsXWH8RqgKgyxREVzPi/
jk1GxX7+DoAl4A3m72c2+KUhK0ZTg36cpBbGp1Oi7HoN0msl4MGwhIW0txpJzyUT
WFWaHaBqV+mhsq5iz9ViEdG1QdpQNbbTQnSz/K/kuQlNiOgM21T1/O26Kd9wp9AC
4MeqGnRKQH7igZS9l5ZSo3fFa5s0UQgUjKr2jZRx7qmCPWzlSPfjB25DiCEy09sN
Z/m1U+om969lxB7/N3W8F7vg0AF8B5sqxCsFifWCwnEsSkjO/dMcJ0OWtVPxrjQ3
LVejhP3d1deYdLhzynvbcLhupQlAlrrKezsxb3A/yM/epU8ILTmW5IRVh7ELA1MP
+dlIsLD5dfxhCc6yGNdhqfOzeZWy9cRpkOMinnUbzrkbePEWRO2ZIzXD4gCqsrEV
6pKc5R8BbRLlQcx+HbwyGnjr07wxbxopKfOZPswTX3xV98/d1ArpbU2lPQOn8EyR
IV0HvhEbOW6IvAkcx1iW4gUXdDfZ5iwjVCGN8f0ASALbY45ba0Ti+cP9Vydligaw
hDu9Caq2dPC7yZjtUjSsupeTthpnZRSqc4eG6AWUtVmfSQqIP8nNEg4ZPYqeSU66
+f1+Lu8KfvV3L0t+OLTXgShdBPQwDTnYF0bVD3SKJoLpd8/O9zk1qujqBgjgxj0Y
ZLeMVyKJP9VILUINW+I9tTs/aindGfhzOY1wYtoZJTNTEmmQiypZi3DtismfSgqL
eJBcx5yxMzqhfVlwGbc5SHV4PIY9ml1B1+5bLLgVIzlsRG8FYa9OI52a1Qxm11sT
ICGdM1t2Z3qbIe+FOVp1rxqPKmYQgdemp1USUyu7uSlwmM9w6P4A2mxWCbf9a2TX
uglBieoTZhxtk2WcqflcgZUg3ef0NCxBntY+fHWWziuIRCeoHY1VdUELKSxaQDJF
t4y5tqlcaI+BN9ICx1edwns4w/4qqjDSWNxR423DCJgbJ6kSY5Zk5tv20n6kOnrZ
jZdeJ+lRJNwZ1ngegXIemutEHlh/iIBGtrOvrWv98/kB8WSXutvxLHWZt1LlHYdZ
NVJgpz8Isqk6kAYdQMqrmHYcUyrzHMpyUE2+vgMyVZ8rPHhDYNwjGLjEpvQasExa
RoF0sWjrBjPzvIJlveFulBP+ZFUSNqh9n6lXGqqyGHfVvfuLgsOI38DtH1JUM60X
0bWm5zkKYJxXb3PxPekFnHI75/XWiIdZblT0S+BGUf/JdXjENCs/2N9cPV0BWKPy
ZeeXiHvcVIICjEkrn2j9Ckhx9gdFlJSLBIvVbC//71w449Qk/ZSOKz+KF08/GBmX
x402Al8vKWfREFurPwbNluagusFL9YgK658oM/dF61WEw6ewfkH9NQVm6E+j6kka
qqDg/lgH7Fmgk7/hOEG2gxCsitKV8IwxijThS+Jiikio8PaYEZEdYbmZ4e7XdIWl
aXLulAbkCe9zdF4gWvQr03u/VaHwW/T6i/+TZ4DKY46uRX2vrpKXj9FTzQgo6syy
YjdY6A2NzjDM5XnUXRFofgic8CdzlszCVt6qJDQRKWl7WknsJLE9VDNn8eEIlEuS
/Iaa8OwYXL4d2j+VkGv/XxShE3XEkj2G3x6ksgDiyIo5SixvamreL3L+DnbDYzoF
5oP4VuoqhsVZftWiByQSrIx9D3tkccxgH3d7h/HwlmmIhqTsn9UzZJ4wRzW5Cu2g
ZB8dio+H54ZgeEMWkGFJMN9CboMfteiyqRoDJ9yuqu3Uq3EykEOAOFdOoTGIebP3
n9RCFShjFKQQINPjtjh5zNkGpasnRYo2EIA1khO8pL8D80pooXvucRL66X60CVsS
Hq4hRuoKVqQ1cx4ZdNfzxVSMOXH/Pat4tL+WJ3SGi8+AWNt/8mBpXFX7QB/cBBrh
CvPhQ/sTHNDp4JDdqarLDcvkwo88EOg9hFJyWSTVsOsgD7iobayAOAFz/v/jFMz6
s82RP8b2dnCzumkGLNB6jXt9pF6YSusKYtuTzhJ/V2XaAREh+M5jqk4kFQECFWiq
6UDy7C8ZlnSB42ZrJSJGYlmEfhgRbdthTa9RCvfiDyGej8oDeXrDNHwpEU8AmAen
e2ZW+AA8BvPzijXQCOja9wyfgWI7hvGHJOY5DHEtfzUQRdYSrZtx+ZadI4rAYr7y
HhzBOaaokBgewCX1rZTtyRI6RSvx2Vx0StwgmQCQhGdvQhDh2S55bJU9uETRbXzr
xKmjsds8octTfKgxOBXJTvu149AmaY1hRjE15TIeLFFAep9BRacjS+yGYg8wYkLe
6K/MJ2tU+hnkDdQZrljEklv6fWcXJdwkkmIY4Zl587nPiwsNtEJWRnwVsPm2FT1P
2o73ScpQ02kyZR8bD8GP9r+CCJYujzPhy1jNWVxVr3SUge8drDS/m4EoOKGxkBq6
VmT8ySOna3+k2GGCBtzie3n88abQJbtR5lkoaZi5Eut9S4EiQtQHK0P8GFYgvz2y
28WnnSBNypgLf4IxGHpc3SjgnOhEdHm99ywKOJPYm01ew1x53RwK1I9t2tNFPFcl
XdV7R7N0u8qw/6PHTjR9BJJ7BrjL/UPdx7EINRDKSB9zLnI3qq8FWhXTUE/uZdoq
klEziGuo7jrrU+J5uPgjGkegqdhqskLHfuOxcWyjxTgt0LxaCu0tIDAk/JWZk2MN
X6FAYAhDPMF6ebBlGLj4LPkQu8Gc1CIiAW4AgW0IreMGGO08vx16aAfHhCgYj8Kl
1xwshj+pUoCjMwQVDs92qsYtw/7UnKR+uRtZazPppTLuhsK3PBwbcgYc1+rQ+CIM
7H8muQb6KHg7kUIFrabRz6tnxxpQs1tDQoVD5wkzLkYsVtkbsZCE384nb+vu9X3t
JYXrauJe6gMvfgEDRUfnbzLktK+N4/sCycv22fc0fppEE6KcnIInKDcsGGVOe396
7WZDjeEPPzyj0dXFX1O9IA1yySeHaIkiZJyPwApxPRmZUbcnJWAqS5+BQbvRYcEK
zgMyJbFU42ONPev3rDlEJJ09usl8o6nVpewbisYFWGEr8HdmpuqJUQoWxLTvqrsz
1a7uNffsZxiRVx21lE8nZMI8cqRjVIYLD6ySOvIfIRn0sJGJbL4g36/CBsP3eedn
d0I2BSHsWn6lIcAyFFhpdR6ygjvmEQa1PHt7NcPuiHnNzFWIJEE+IuV7R+AOIhE3
pmzE9oaesx3Gw1uooJUrqdlXPIxMXzCmo0z1fJPTaDN6Sp0A1QajrZeGO8p/2uB7
eXGeMhnBINqpOSAP3W1KFHlmgF2LiquDpLMF60PNplwvE+r4aOlgsNGSLrQlPooY
zA0E8M8AXpVgh0DeEeKN7uDODjOXRGY/xRJKp9fgf/3QuWXtuqdh3EG3nS9Kafbk
Zx/AJu487umtiX6d4r2ekjwpx66YcbR7pelpacPaCQ7ColYJwkyyVm/Igp5ydtun
j3utEuOiDqcIS8BHTM9dRam04zpoF0vuosduU3hMEyDGoXSkYcYf6XB8PGwv8t7Z
abFR4QONEnbXI79qYXETBTmjcpqz2l1Debu24iwJ9mLG2eWOkVwd4QrsHIcq0/rt
cB1qGHXb2ImvBS1zLDVTrZrASMnLrDIiteqXuRXex7ZeRtLQqJv9U2CixJ8d/708
yXZIgFKwYkSWNrtgjSYXuGw0atVm9euG9pFzsC2/Y29tbJuDVt+cOgytXnFCfwQg
/yfzssF3xH+D3Oz3TsSKNZMNCk0c/cXj5V+icoDIsko9ELI0wcAGb04uBbKbw/ct
6P/NK9hIJ3XXNcVn2FHP6kzcqlBCxD70rfzE9ngLSQH4jUfNdUFUsP+vrfCRz1Xq
9kTUVg3Skc1DrWIQgOpLV0As5QSn0e6LpnrUrnbhGK3BG5kJpdA0UUsy8XB8Zokq
n6e8Oa0M0p2aeCKwqu/xq7Rc/enEExSe6LX0Tcc5SjNw7G631wzwFin3ciBmOfTh
3AblsJhWPBfixsal6PmW20ZxR/YErqF4XAuAQKeKyL8lTeyljHdxOlPtbm0xj6bT
s/I3S24iiLsQQ/Hm6erX37OeRcKLOW6b9VR6N96o/Zd5nXSUByt19FytPJU/3cF3
waZ8PbYDnhrvX27Lxck7ZdL+LFQH/j+jmV0cBYrzJWvbzOp59kYKs86LVx28hpWD
tmB7HxDkOM4XSAL53G8DdcHD9wPpgXdJX2USsfHa4XBYQDs9M5qjaT0WpQ162Hpd
gkesF9Lbz5JX0smPINqtz2sVRwqns4qzopy01yg4123M+CmckTShMqtUmlXQzaBj
skmzCx/bLeKBK/wTfdNBxk95HuEz2zWpyXcyfKDH6LCimDfftImIVjQhJ6IDO9yv
dpdaiuYV+SzDVpAfmQyVZ+3/xFQ4/gh67vFiOsQMVTY2nOzX+0CuSwbkI4dJu7v/
ArI1YD6Z0ir7H5SyGbOinwqYm2RVHRaGTmLjse0TD1rtDI4RyQRA4mTaqlSsPbWa
2RY04DHNlkfYU+Y1CNDIlZxMPjiQ9ug1dmnn67/7psSpq9NSm18G+M9WavXj5Yv8
hW2s/W7zF/SGOWJBcIE5F822ElG+q15freDj80uAFZS6Z43pdbWrmZ11rIKWt8c4
MREvc+/5Fn90lExmeluAOn4rfoFxTO3Fv/yOqHwaOyqhzTNkXe+d6ST5uU9EoTP8
hmcCkc0dWskASZe5Y/HjaIj7J63kZ/+c0NuvOroB8ATVbr+J2BRh6fCnrF/bG5eC
NR0DMqbJ/wk41TJPwTK8ZfK+OAfgejX0yHSSOdLPjJAN8wLegOzKACPVPYmLE2vd
/dv+mh88++tEQKkU0zscpPEsRLgLXA0eA4PKQwEuLNidvxkAz+3IMm2vNpW3GDN3
/np8Vi7yAPXNE3LDqxj9wxUThqo4Qghvd9uehnBkkHFdto6U9Rp50Pls3a/TtO44
Deg8j9ZLz834I+qlX15S91I2PBkL1CxWJRpRpiH1azFR4TGyzVwhMw8s6Vh9tlIv
KG4OasYDpT1M/qidHlKU73a9kxoOJvjSQ+nIwN4NIyKQAIja1E3xT6ig9pn8Pk1P
LdkFKEStt7Sbg7OYOvnZyE2QdX0OtgUNeTq8P1cKXs6B7vhvvA0yqsabYEHQlmy0
XI2nh6nqOFPVGoth6sRgcLlKblNj071gIpIB9XdPJ3L+WgVYznOxqKnkBBnownm2
WJqdLcK1FKz/6vahror/FiS1WR9lV2OWQgGXkKgm668Ky0jJMg8pNuUYMhpC+Czq
BbTuVG/vAev+CrB0NthjvJzACapxoPzmHiyXoAgWKWtBPmmCAriCh654UZ0wlawP
F/PFQBmgcVX3maADPM6DX3ixRTEySjEJaO2TgJHhf8XQ0vhJz6uMoKCekoPZUrJu
Osqi5SDCJAWk11cjNprW9re1S7OjNStoHC6ljdBaVJUSEkzmyd8wGO5rl976FzvG
Y7ZeBKHmXAVrs0l2m1x9cAngLFI4NAnTFpOBXh3mLFywOv2GvJu+ev0P3EnnZzPK
v8aSqhl46Bw+07Hw6/84ecvO3Kb1BrF88pSprmU4AYh5hjDfuuZWXdVX7jQF/UZT
DMhGYS4U8xobUPfCHPp5M7ZHK2Oc3MonK1FTWrygKNh50teqUpMcpbH3zUG1h8jz
c2d3n60SMLOQQLV146vLiW86OyVB9XUdmBQdXz0BblxSuJ/hKWZqhZ3kWAEyxEvy
MPtfOW/6CkVHFVu16qXj20/6amNZm2TbfK+etoEgnuaM8mAm7H3ZjMWgHd+JmRQ+
LW/jvwgOvwHGN3ryk4o3auhxEgySNR5LEv0WrFOY1o1w/SsDpp5acARqfqsFWSF3
CQXDphVlZFDs9ENJK77HM/RGXcDIiP4qUkn8dIlDCwy1a3jaGlS9eMPfSt4bgoEF
L2ZUu+YErvk7ow4iNA6e0C5LvEF9b3RF4VATLuFN0mfDZQQaNZGQuMG3WfrFGdHn
jshDqr1T8oCiBpXBg9847dCAxhNSsJAL+ROArVnUJ6Ubr+OOtSzczbqINcRdWHVx
9V9vLQ3BSWymUdh8WY2zJw==
`pragma protect end_protected
