// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:39:04 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
IVaklsiUDMQVcL5ey8T5Ph8ELcAwivsuw5k2sA8sw4sStcu7Bsri56OLBJ2NacB7
i0hMuWm+aYtA8kDhUVDEMRgIHmFdNzt5QdAv4L+9H3klKq6sXri6BiF44XbiqBO7
nYFc6L7Rc05QRWwTcn1MGUQpNXc9yOOHpY+7yVdRpCc=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 17488)
FHg+scb4XRo0ZIW4L+STumM1cZpqzhjUQGn68ZwHfEXhgmEtuq7B4pKnBtZJk0Xd
eg0ZLlVcNidzs139Mpriyqb11KoVLZqi9K3XmUSgaMI/hMHfnVKLymbirKzRNR5V
dGfeh2Pmln+IPhUZZMuJCy6sETFXUDl41shOciKufOJFJvaxnLIruD5kBOSjCFT9
uIonqPVo/1H3SZ/OVI/0r3aNxN8ryfjZa7GIpyTQwUPaM0GHVAc6B9bG6fCarzfg
eWYmPGJXSRvEcSj11/Pt/TOXQx775AEsrNhwwJ5TbV9NqQunzh8XjVyekuh3M2p0
w72n3t1w+0M7lVUI2kQFpyEy68j6Q5W9cznqAlx51MAdNnvmmNzQW8jNt29Ra45V
JBLSsqFexk/CdwIPIO8nC00rN34UZu7o8yXdSLh5S7f2x0JaNu0zFII2RzlqZt0I
bLuXNfTqsfjxxgMQVGQbIMGtu7KpYhjeqjel0MdS85dI3XaNwu9bdUdp73lEy9Og
9spv47rih3OjOG4/932+zZztP4Apo22jtspflOOR5lJQuoNyhdjE9X1z+399Ya76
U6ixBYRagxRasTXbGi51o/uNxWwqxGLIMBr9e5fnVvN42g0/pKBLO4QZtDuI947E
griUAwOi95IZc6Wh4RVjmMQy7A7aNUFar+7Uy5q7AQJtW9GP+GqZZ+jl4boRvD3Y
khgNzicuK079CNaoS/GtZsPzK6hoiRf/XTbJJM3Uw6yCdKBvTDjWeYz99Xk1S3q/
rWZg5MEGww79FdPW34hNwFgqybQjO/XqDakRqff3fD6t1QusTrsksfekXBI3z3gk
U1YtroeozXLs0bpygGNBhihThyPZsII0+QsUC6tg01UVmx8cqEsypewXIXlI8xiY
CG9jjk70SlXJzi5+9dzHfDIvNAdAZHFI3OoRQQzhgDUqsBROXufBw6MT5x1Z1U0K
/mY1nHEGrkWEzxcj2KLSEuYmQ8kCsWGPT4irXYfs2InZdS6EDaVsGwSakIF95yur
qQPqjY50UX7FMjcNfUxt127xXmahUQJ6PAenksQHLRuV+Fd8hgyavTbZWkWp4aAr
4MQ2mElzVP0z+fL0fyNvMOsbhkYB5gb8CPem1NvsPj0S+sKOPvRxDbRd9Fq+ruuJ
kQOvOVP4uoII0XzkDBoofKuh4SlyCmI4a/DLQ/9EGUYV+hJXXxZPopwn0Btkktkr
Gpod6M/6NLM5AmYRelg4hAkpMwISw42LlazHvHPC72coIo7eWEa+8RALU+IS/z3Q
yWXOd5p027JIz5yrJbKA3yBY6Iltsbbr4Zy91NJi4a2i+6wWr0D+FF/3ZYT+zMHF
aY+gF75JePSxtrLDecEcTllaH4tCZJtJIyv5jtZ3ZdbScZgnn5hnkItMA8knptaz
4+q7u/7DxgEys4u8heJ7nLPDC8QeDmC6PnR51EpR8HhIOJ6+auls7zmflpgcogYR
mMD9Da2G9jq/qJeX4mL7ff99CvPlGXDab0hTLKQrnXQlkMflhuyNVWfMJbY6STyF
RozcUgg3KJvppCJpy2a8EkuV/HPnQ19Dt0oJrV+UtgIjy4bVausQ5Ctdf+I7jGD6
9Tc4SZ4vz4s3NXhcEAasVNOBTMYd3lot7wGqFO1lvJbSeyAzdCxwoRDoMamFtxcM
6HIO6P4zJrPt/XX0EHGUTQWkuu/tMVq+f2+m1e0dCU0NLme4zgmTn5OnrTaohE9m
oN6F1wHlPp2O4Y8WmUxfxYX4GSZL5IAXODFn2mQ+HwFU0EjXDnVxlhl63kcCF3hl
UPshtUmIFS5Tpdmz44cC/WBHnwG644G9SYB1KzZfkh11pnqThW1Vrb1XgKBlTs7x
vmDO1/W4wPx9GiRjI0hIt7rZNSuWUNfNsgJOZLK2nKlxP16LK6860EWzduN3z4+X
65JBu1W/q+R9LMB+wikZsMro69lPWmtCQOynzqUBMhf/iXMz0J1BZAw0TikPkzQn
QObGIBNoASrChNt4+UyKgyc/06sNKDh3AEUI95f9sK9BXC5mwpwRy+qduoo8VC4Y
Z5Pk/UM/QrGVRHfONKFriyIbdjVADIhhW1gZZ8OU+Y5GiiIKUFKytHSp/kUL7SKq
7YhW3mdwgN7qgTBU58Pm9gsg22s0XeK1tA9xuE7rqdmghrEzF1cEFCrZyud7RQSu
2MmeP5T6uwF3EK/vMy+cIcLL2TuZUUJoElVYsNvf/DQEPh7CbKBautHHQB4jAnvi
so7yud52sTrA6JmI8LfzOQJE2pt2GIgGry48oT/X7x9/IetjmogbWkzYAafvWBXn
Dzwbfndtvilde3HR77u0REfAp5AnBGC/BhmLeSIMffcaJ5B6pcKdKdecoldnpxQw
J9fsPZ/h8PewGsj13htsm3dNiVEB58lR0vGPIBXNl5b3NrdZmaeXW2lShJtO0uJA
yC0tR5Lv2WubzVYFcfwy1G5Em5gqbFhh1o9RaAb1XJWmEWV8H7bINbaDkpWas2ZI
5AkESnftHD5k05he+3OJ3HkdOv2yrwmCm+7IVjc8tNf5/Qkxdew5nEYQxPQ1LWn2
DPjUBD6IbOvCDGMe/OKxo8S+kIhb9OOxYXHVkMVsICI+vwXbv4M1K6nwWWTfrVs2
1OaLM3MPatBBgjZNmYVu/S5tce1W5c9LbDxkP4z46ojbbSKipKS2yr2wCF7dkcO7
9r+DZIc5pnEXzHm3j6jfMX0KmxShhW66PZOmRtlswKIMg7YqJb+pYJ9caXGMpApK
ej/HDoT2aF8YMXqq2nr9rSJdNEZckGeBmlRrksEYiw1EFObjVrLudw4Si/WKNuSd
BbKO92h9KYJU3S8JyqfJSwO2jmAaHeVI55QabDAVzwliou+y8+1XZ+E5bBv90qxJ
EgJHPREk43PYPxz6Z9shirULPHe4XMdcJ94vNgZlb5jcRGiWFP2m0YJOQSHDfpOw
qwV6ZW6LlpOQ/WEMMCOAMxmxgwkHw4RiMl5Ich1QXCmTG4LsDD+tXfoeDb53Q11C
VgyYw12AS6k/Y3IKICBcbNon4EHA7DeaBThaoImuk5Ox3Jc54Wbjbw+fuU0xumsn
aA22jBgzev+LFdtokK/t3Q3oCt5QhZ3aL4ru3RorqPfYDShyEdm250rgT1HqbiBH
tjagv6tzMWpin0JOBRL+usa+uml/lRke6iL/+0Ct18K1XwL9FYc381D4WopjADYw
pZBV8hzgqbVOCPhlTTTBsVS/p0Qc3j7qK7RwQRcpLlF8Y6+2pcExu0r9ZhGttn0r
dHrSC3jxo7IoqW1TFjzfF/kBSmAqZ+CUTdJUqLtD9u7nVoIeneBQoNV7Ujo/8IYy
ZrRBYVudwFXVZYepbq0skG2V32TZ44TyT7qpe9xn3ENabWOTmjDuK9cXbTAyCjZP
JUkjZkxa3XtM/NPzYaz5ZuIfHDzrWXabLDeIyZLIn9F7DxSeQYYwla3iJcL5nKj/
V4CaTFIbp8JRUe5ts737BDiElFSF+dUVJkA3BBsrWEMDS1Rc3wVy2uUAezKNhWjp
DRvfg602rUChNAwWXtaAkwrJTRX4YN+FVBx+GbnNSLlPeAAl5xAodcKMYkOhrslH
L8uUlKPU0P25RnUT7GX+WH0Q13pRT5e4TvWy5OFRTJXEHgxotZcV7WdV95iuOcOO
fkLvnso2alFwg0hhonGlzU1i01Wyr5aJHqOIxSHwv/RkEXdkPdCQ3yjEZ+VTMM87
4T9vWhgHaB623n1Ts5rWsq3RcjGPzRp5bXXRrxZsj6MOU5/+aYxEuW/qKiBwts2e
xzp2jHySulagJP51Gd0Kc0plt9Z31kF5CsDSLI4kh+vTfxhjdDgD/o4tU/Fcyohj
s3dUaeVZHB80bCQMg2DV1C/VriLTHrWmi9We4YSZ1+HgwtpU+Z325OGJSsls+NAa
V7qaXQTSNGLYX58R/uwPtAFyROJlpWCMdYEZ87l/RkZ7bxuvec6WI6bi/+paQ2Es
EXdSutQZF9Juh7K8qzaDu3Dz7qPldPcUbES4o/7R/5MutF7q0zdJUa90gVbkfLit
w57HFDTnSM6AOQ28mSi0RoEFMwKCpLsItkx/mIKi/LBh2qvgU1uF8bqUVMVBaD24
xXt2/BjoqAdAEzze3UYVRjRK1o3zkA+X0ycx3JN3R9TsfzbvXrDVCCctQgcNEHuE
BVzjtyZVLaAwOW5mJcTO/1OjTvOv3ex8zOrXe9I7svKnbzUqy5SlA5XwNRKO01Fs
clVvB3qTJxdyAatawvp4YylW7S7Kgxg48PGIpz9j6yrO4MSkSZZUln9GuS6bJ+nB
RWZvwHkahWHsOT7FRIh3//kv1gXxBEvT1T+P0jL7LyyZq9fGTT1ggkvaK6NPKlrF
seJcO2WB8bMEPkKxd/U0sAtuMYmDvVJoijgGiDXWbp4eqBBDuCKvrWb+VGRiIwQg
6UYLDdj6HWT2i545/2Wi/rmDroGPNRT+5xC882IaD4u9IJOre/uGbXHCQWzpvihy
SwGLOS4kgysfCC3Il1eW8blwF4CY99KETljgn3UGOvqOqIS7vYpg0YfgX5EWmrfM
T8TOdGuVPJQPzAUp2DGhy19DIkHoJ31VSNUQA8bRUfh90AEyylQZJa+CoFyy5oFy
GmUbMGrZR9Q3KMma6LLNdO1PsUJhdhcSK0LrmWykYfWot/RS8yxksCe/wvFdnN73
n8uaOJ/DRxLr6Ii0Uei1N8HTkzid0/XdrRvVcGZfv42AYDo82TxyIiUvM/nBs3IJ
aM6d0x/M85A3/XwIALZb3U5Aw2YfVefZ88zXdDau/v5TH48PiipRzGNuubIMbRC1
/4FiYXySdvHudiV1oCeUleHlXaa4t1RiTk9ValY11kKHogJdSBk2CFevcRruuj71
phEWU3e8G7PMlIuVqkSvsrMl8fcXtS6bDzJgMIVh66zB/8xuoj2yAto8RsURORJX
4DTfkd2pfRxlGmhd9G7IAsGslHMsvkk4/Zh0hDHSdWjWYcDoc5YhY6dR3UrHa/+M
2SwhETZGsJYf/MdnY1e+jvP15ylAVbhOVm4btINMypEuhKyN3DKrbi/PP2D6WiGd
b++aS5lmxPqNXlGi0tFO07JxZC1dQjpOtya51PDNqyAbRLYU3lbfhvJkkDOMqKkU
mh3n3CA4fXOqZgLHqA9lmJw7EfLqIWzXCeICZ+68NUVodDdhpCbTDKxVnYjmoZlb
FDVZOrZ+JHjRM2fW1RWNKKmmQhp2IJy6hArUxlNc4E4zX9rtLsFO8V2jLP8DfMUa
LbAt3cjLxQjfkCUGEyi688N8MId4abDyvFYJcb1c07FbU8IQupCSe/AIX0vUWnH9
Nk9KL0G0lFycDpKPFLbqsGLuLrYHiB+mpXzMhkE4z4m3mUK3kQc2qnUwq9Ga+iCP
qIW/g7Awfbunu+u5JrqCB/feKXzO9kpnlpeDNk0+UtabKO0uvdTVKaYTKQqTG5S9
aC5UWjjHmw9nyCAEXJc9DRUSpB/+F/i7+4kxQ7zm2/lFspWhg0x2ydgm5uOUT8V4
Qy0YUvzDlYzI6Hst2gr2SEFYOO1SHJ61s0u0GQF+PoXQ7Lh8CxDnE/cggkPvecm+
KS+DeOyh9P59xn/sBq9hYpSpDVny71CkaokmI+tO+bl5XyFQzVXJl7vodj5cOikU
w48A8l0GpKjo+3aAHOxTyCkdcvQVCJXlQ5ZNIfpE6Nb8rr+Ut21wvVQeVP6qhFsd
K3wLFx/Hj2I/ITOTkcVV/EFYt8EIt2KTitQBn/RrNh/tepTkVx1yGQZLOmgbw8vb
jH+sBIU/BlWiOKnUAjuDrw/IZ9Til2qeICITsnqh+1yA4sbgVpHahlIcp4HefFdW
1G2eQ4hOy6utmWz7tXRfh9GWxZOJqKvpGebErhwCL3B1akk5rv6Fsgi4y8qtNIAF
76Y6zOue9LeuaP2Z1R2TextJvD38tn2/ClHaV54fIYR54h/Jbx0VbKK7teiHp3Dl
QLspYGatY7EjUygF6xJT1LIsYA6r+e+SOy66KS9VsJ4Eeq1O3kcWOmdHy46aeKuj
f4ssWEk7GaRjTv1GC3JSxJzS1fesYU+9fj2x2T9JrlFNPBZaCfWHdqh8hKAGK52e
iGO9oJ/URexaJ5b95+skV+piaBNv1cdxslhzWn/z/HBr434dw7owfbqszhzVl+qR
KkKF+iKF6dMN8iCFrxGOjp/9bP7AMVCsYh2mD89P4aJy93k1qYTlT+8ysNczqsWe
3rO5eWoz2b3MWDgg668Tm0h8oSQ5W79N9gnLDijLEFDinazhWGs45Pfyb+pISUHT
jcoJAitYZ0BIWaWevljV2HyFm7CIIFAlz3NNiMtl/+v2YCm2HVdoXufzVBcgg35K
GlXTkK4Tvoe7UWkRc6X0FoLwdH77R0jyAVqcUZ5M554olNv6+O0Zkofj//F3kIB/
tL4EVZ71Zk5dt1vuha0iUp2NyN7PHCEKHG4Bt3iiHOBHKgLcw5uv8otvmpzDiCKr
6Xc2EwvaVT4+16wBUfUOprYVNXKQN4DeOe6H/1cvhYvZ6BBjyLtuB535Vz2FhazT
9plUsfxgOY5H6Sw0/IXNdvudfMWAwOS2QRM5gBDCLlFvP3oTRH+Dn1qjU7kcQV+3
TuUsjaCB3t2uvBgHxWQCDev05OaFcAhZ811UuecScPiKFRtakdqDWhjColMA8/fA
qDvRZnlO/d4Dxm+jZpVIdhxNsAUaDVahFibYHFP2aYxKXu3Ybo3y8f++RvO2I+zy
ONTDNqr87l7u/mG37klbDkto+RE6gQgQlwDqraFe0nWrW3Fv9tvzE5XMAVbnSkN9
YiwO13ERo+gdnZMdrlo+wcep+fLwEOt8hlhHZaZn3CnJIdH3SPv/en4Vw9Fvu1L4
NKP547I8qbs4tRc4Mtgpb0DSggUSn3TtZq/18RVEhfgMau6yU58JxTz1v9HhfbDr
5ykaIlIx6I2qMLmhB9Z4hMDLOxXwngbtp8SuKi3BYBxCQzznTwvvFEcGthc+hb4x
4/XikyEQ0du6pdeO9mVV7FbCPOr+8nhAE1d80tyUACVTsd8PJIDy7anZD6Q4zJ9I
7j60QVeu8YoIRILra+tCOMtGx1KID4JWegCs0xreohHiWzBlIiWYXdUv7qKDaQY6
LNah7dz8A7f32XkhyCsR9h29Oc7GYfu2SEuz3fMJdLXs1TjJqRcgS0/a86jRQCIw
mZIT3dErQx5mbbhClZjy21D5fnGIsTkFkJRFiBowRO42YwAnpDOzXAvo1+3Ra4BD
EuaN93U2EbMhSRKTNjYfB+Ao0Or7RxT6os+E6nx6nDLFeCIaNMY18WZe9uj81JJW
1hi5D7rKNSishQAFnvrLx2dBJjIPd0bZfVRCWVwA9Wp+9btIA61OZjiIYIUqnXf5
VlfDOfFwGtyvjpNgdbvQgVWJhL3Mu1uU1MEgMSYFFQRvt+akZToztCyempbIvMt7
U6nVYpB3nE+dlEXQPwNT2Z6EfHurwb7PrMcZ6YsHutca8L+P36UKtvgnKjgAyR+G
aikYk6A2MHQ11JMqonZN7QV58Z8PNCdBt+9MyXgV4uWfyzqSkjrSY83wsUGSuNoz
7HQxGxj6JE9sCRr4TcrpHMahz9XEts9DHMtXdu+ayaayaXIqFRt05jVw6k00eVXg
40X8NbdU13UY0ldiUf6hTdZWYMcvz9BIEFps3EzkOw+nIjfiIYgWKOpedTaodJLO
Vv/2HZZYzRiY+HX3em2iiz9sUtZsL2q7NUS5+hTO6Mk51a46eQQvHtphGes78sJa
hFsszkIJORejqvLADy6DOV+gyLPyu6iOfxD83LGbFUy9qPXkjkxPpNCx4UgzuMbj
quChTxLkLx93/2FSgdH5G3xZdXmsREcVZu0wssXyxhMMX3tohqehOfQ/OkMIXFLt
jp4bHbgf81bQwdIEjsyP9GdETDdf6flHIBtQgGGPDYpV0eEu+koYRt1/5nZGixJc
csbU8wtIcOSGh1dKaX9ZFQSUbgwmNh55OGiWI/fNxolrMMtCnlmbgGIc51cgBXQ2
WTf/w5hGLk5g3vlcuMsIHKf8YNki1+PHGJQ0Py5Rb04mDLWvxfC2iiYbxHERFs/4
u+n78ygCbaZ5XlqH/R1eutxbHYZoPa75FsHio/BUU5Bvym6lIPkHBCzCxiyTvgTW
zF5G7jZv40bs+p90Q8vfXlfr2QIVBSPYd6nK8BoKeGDScTJtZzTt63Bk0E+V0IeW
XPTT4uLQXoLUi8tXLe8OVGkMsNncl5aJtkdCttU1Oh6viG20qP2trXzV1NrdiLuu
h9vybbxar3aV7DOvEuBmyJa3mozzAS0o7I+EuM8wpb94l1iOs0bq8zLz0o00M+x1
Yyv2TC0/vW1S2Z6OPFNwtUbqPV+osGGdtvkUvtGPL+nw6VCnmjr7OF5Dc2GRbVZk
cvBADQcsRUDFjyCNDB/sKkriF5kA02zQNl1oCkwQKMgsi1FAKDrEZSeA45Y1rZVI
gpdY+faC8mh/e3QgmtIJMRNC+qbxAnLLZ344wjLp8r6MwhE46P5c3Cu/oIUaCpPE
CEXRj3R99isATht7DHHsfLrAzs7qQjY+KfH/y2Yap3cOLC1ITmhgcMnwsxnm+V4A
SGu9qVtv/WkSa2X7Wgqcw262acP9g2C6RXjcRl4BS02kafBmcGx39ZR+et45yl4+
8kJZcZzOw8RijQdGoFN6NPKnDhqkXO3fVGetLPby3BGfrXdwgnjkeQFCwmg9Xm2O
Y1omJCTLsT/X6pQNj4pfgcGi3HJiwsfK+t/EYrYPSF0GfP7PVKx7OIyjI3xoyBf5
yqi0FEqeMQJBxaV8KcRvtWUjS3rlkf/xoK1yF52wZnKzhk8ab9kdPUNnsuy2oTs1
P7HJ7XJ+G0aIAYt+G7Y3KhtxoeMSMm8xGawvx0UWeDg0iEvf/w8iolAJGZwM8Ymo
P+YDKf/akQ4HMGM+XdjW1zBp0k5AToPkaCjcpklPA/iNl80A1aO0CGjkVQoAhXx8
VqSAqAGTMWSpejdxNwjWjMunOMNuz8zTQTVKvHsXKBIMGGk7Zuo+/xL1NZAcY52x
W5jepHtVl5OHLq77o+bsFE6saQ8xaIgpO+I5yl9/A5CZWHcmZMian8U3VdafQfRE
x+TGn52l+OTgLrfGDAv9Kpy+0IIHqup82xSx4exMPQGHuFV30aF226nGtiv+g0Pd
jiafiuME1OYhR+OQ07Z2W6JZyh5Ya6PEBdwSSHLKqY5sr3Mqa+I3iY2KD+8Gt0XO
SdZqMtXOTIJPlCuCA/AIq2UpMyBnYdQ5K98kvb9CQk7uVIfPY2ixmQ/MRoKiy2Va
dLSSHMVN9eMjsagsl6PiynF7841Hd4dwtxi/Dwc9C823uQz2nEOp06/Eu5IGQPqZ
xo8nKa5N8DU9vz9V0e6BBCkzoWpM37th5BmmVPQwtxQzbD+YG3UPagV3jVGrT3Fz
9+snlTDUnDhfdpdminGroQ2/UjJOyLcIyCrf9K2u3elYzNiXXaS7qU38gZKSfz4M
oaMApudcfqV4XOlDWFTEk+NKmUHq5dpazB147LZoBUNF8MA0KWMTRCsqsolVOJGG
k+aqUff7wywXzrmRtSu30Mwm66rtNJSC4D7OJi3qwoSB8dKny0uO5/swcm6mG74A
6ctIgpWYowU4fCvRr332YOueaqPlgQs+yBG4e6ico7+ibQopWW9XvtLCTJCMdClW
JKJAvG50rsSXTNKLotboiaoSSKIpHApMmED55YZ0HO1+QEgBHPtA+ZgeddEUs4ZD
AmJsZn09nqoCHBLRvDecW543UI4jM/TmBfN15Gb/NQHoaY3oJPKg31f5sLsd/py0
TDxhxy1zTU7QEeS6TGuVwEzGTpUWZsvf0zcQf/IxLHmoNbLMISBw5+qrtmrKkCY3
ZoL7GHSEI7e5Zc/COu86+P15UpoSf/t9uv4bfH13VDqGcucoqelVZwfwavRmpnNo
VgIRulPqegk0g91RVMduFBfLDjxjcb2Ve7knQ+mtDiMjWdgn9Q3dPHtT1z2XtESm
P4/rRZhsOhM1hOlP/sMVvST4pA4Hc2zF1lL/D2LWDpqeZZlyq8oP1bQQSN4eu/8f
LEtgUTg9B8Ljokw5su6kEKd9VPt6zsV0ki7xUUMN8CEhgzx4PA8U666+NRmMlh39
UKjO0fuIwpVOoAL/pQ8G5aAyfiDZM4KmIFUIvOwQUAEy53DZN1BGlE9atFCJbLZd
v3iZ2+wAwqnemVbm7GPC3++gSfrzu0+z0tI4EFm3+yVO4Xgf55+kjol4v0sXtoig
GBebXpkD+bj0Dirg0eWE7tOi86yolSv7rJ3IPkDztNtHEdvhRKwCwHiOSC9jFk/O
3L7LSp7hhhpzgkmRv4Rq/9PzwhRU5K63ZDMCbvbFUQieiHt0v4xRgZyDGwUYP1IP
DxTcifMdQZkbSTuwHOCSbltfOhKIb4utUzGw5kIBi0l+kHR/RhRD+Q0keLbdpEvk
NlqUXgSYEd0Jt5x/OzIENknZefwjwYR16qzGRFGYMG+u/hnjxFQIVKZKarkCylmq
B/6M+779X1fn3aEPcxheDnGHz0IYK0UDx65P/UjBeZC6afkz9oXRC53mSZZL4+K4
krJ+f5ZgMNMFKDAMDqY3xWG2nPmlHv4D13DE+Lnjy3or+GgQ3gg2r2wb5JFLLc26
ujkMhbM7h3HWptv8hG5WnVl7w9IQ/rPUZ16ePvK9eysnwp0lUKTJdb31YZ+ccGX6
4l2/sGz4TaOvy+eMmH+aFvGtLxxowCgyuSfEO+E9Bmq4iNZXc2jWtxzQ1qK5E+q3
YQxM9Ve0b3krr0XJ4zJn4NedL1TZVC05GVukjzn1z++CluFb3lUx2GS77Q84d2dI
WpBQptnbW9yNuflQzvdift+FN/ZMOkZrV9cRG5zlQ/bV32buwrU2j3pm2jkSU3V3
L8N3mV5YbKZMa63NaGF0wNgMrbqyHNhu8YVVbv5dkzRimQsdGJB84T52cHGl94mo
VX3yo4KGSyeDKq8P4Tuku9oNQ0FADtFPPQqES9pZaH8gIJZu9OjbVXZUKgcVL4T4
0tF8rQ6R8z/uNo/49ANgrn9sLe7KSAEex2Ok6xCl7cmM6seNIRXHa6QwFnllJQrC
Gz1oJuSykgrP9mBcuzye7Xr57e9SF9BE4vIUERIyF/eO6+ENb+J6tjJtbjjWL2Xa
Oayf7nsnHW/GWqgrP2HI1QYpy8IvgyFxIm8XBxgl4iVylH7RKLFsXnfQqrCUifg/
odHQsyqVVo4EFu/AeFRXYqoD83SNtnP3Jn9OBNyMObGCHomK/FgWEAPeA31QwfXG
PPCaQb0EjPqIRFMqwuTGi70w2FtiI7wiFMt+a6pUW7o1C5tah+jLWK414bmJbyJi
O57I0UusD/bXAmEtrrM8JL30ZkoS+PVIv7HbJSVLdjyjf4afM6la9S81lA1zUuDN
HGkIKQx8qqv3X+59JDeFmeWk8NUrAyYLPOopFbHez6rJYAUegtlt5lQKijCz17gz
8cs2g3B7BMX6qAe3xyVcnG8gUH0gFcoPi/K+wNnTomdmWsXscI1cqWXDYWe52tWa
eUzQGbtvwnFvuuEJ2QfcwJ2jNGaCh+IFOofvYeR6YzZXVY/7Z10CkcBTTE8MpLsf
M0hBw9coVfFnlLMvj6To+9egLssSruHHNsBPHmE1e5qv8Y4ydDqM+smgemebBl3v
3RUocigTenwk/+ysEiEWCmzUM8xS9OrnFPXU28jb9YTx4SXtie7I38VV6K+D5tHR
vqI7I7ELdGEmDfUNg87gJQ2EKIlVBvyeEIm5yqhwflxILV6puHIrRhEltrp10c3s
O0OHZ7VZcWzEHqeI489bZrJHDjW+ksmftG9x81jUVYtMpBMqLR+UyKnJPPzl1Y5F
HtjjjmDHSHIT/m5n1WBL9Ov14Xe/dghMujrL0C/tHjIps7i6ABuRfQxERQYk/voF
ii5vMSH1X2T/ha780805wtKav26qQLLeRgFPPITa+11chUWJRiiVXmgqHZksthlm
ld+5esjeh7PGrSko4o5P+I2E12HltzJIcw710LL76e4G/cSNtN4ShtSTyfVOgAc/
juUsra0DtkJdloQTH3kFxEUlSeblXcS9cFyIIqp02TdqUeigknIM1y6HSh4WP3kL
50HlZfdY56e25QnGEgaIL5mOtVKNrbOw20l+13VFnpAwBlZFsRQW6GC7gz5RlGKq
HMXGNPvH7NPpv1ZjENDKZyTAvL/r+h/iolEOxgh1NeAYKoVzJLbo1HF/K3AGQLMo
/MWlE+CBwkNup9RrmgF3idTYNSl37BbR8/Yz3CbHRhT90zvAuYCUlmyBPak5q5xa
OOAzgJub87GZy3dgjx9WaEwDjL6fczi8EelZD7AOiUN8oRpvrqcpIHelPstgi1vi
YefbtnD/x5yfBIMdYXCKZu5FDCujIr9QhLa0FfC8aFCViqG8aOO8z772AdnHPP3h
ZVRHr3ty59vvQszqWeEpLRrobk0XeGpQAseZ/cshdgN76Gf1Gf8NMTh4zdQpbSNW
JuGihERoCKjqTbydiHaiSgtsbS3Z3raYEP++ORfG5ZWz2xdPdfX7ebYObTF3+QKF
3Z+yWqActY/4tUkV/i4N8Lp13v7HaJC35ntD6/lmcjxMZfGTaH2DT5aWRYCIEvOF
cIFfnrzeyGvGHFe1RNqhLkUeDVAS6PpNVsuDwi5W6v+2kkyOsslqJeBiMfMWj20z
HBaHzpfI/R657b9RR215mcllNwV33oTGNDroV9EhrSC6WefBbiOIOBBqVE+MBXFY
Dnf/YZ+A9S9FJ0fdMCh2WkrTb9Ykr4Ps5MNbx08/VWrZhg+5OnWrybcxeOgvRLqE
5Veibc0CRJio353Y9s9bx6WO3QmgGklkDM++1RRx4qUMoQUKISzfgzSevuruhU81
AOntP38zHbAku8421l/PqaHtWFE9yZUDrCa2sRHXEBSVLKdtT5aJYExVAofBnR4c
6Uj+Kr6OZhWuiyrupYnqK5L5hH9Qnr1K9lNp2e1PEqkH/jV1FI2B3q+opl/uR3Gv
25OsIbfDZHFi5Ay1/wz998A5HuKcSWl7FRqnX2BaoHhdOwkm5pLygjhAeUuzGlWV
cmx40SoPy4yQ5nkj7qwNbmvX8aKi9sq7Fy91qAZRmOxgPEbzE30zL8plY5iQ7kf+
NaUZcnMAHIwSnIQMYqE9xUGPRuBk1pGqpSvXAKMS+VHV9K629ILMbUm4ML/pS23J
Rj4qtWCQ9p0CpFeuLeKFle6rzWXimRCciqOJwHkxbyo5IklDgWRT9kVpIAPTkbmB
AtU92BT/cBC3fl4tGmKPmx58hElKbIKbd3w6xdLfD5x63eE+F+jHHeBuq4xkmVNt
THEeCw0CdfwJQ3fmm4rVX0jeqoBtK4N+P2asMVrAJ97a0NDxghzeCYi39n/APT4m
ju9NoYphb3w6HlapSTDWjdiCcoFAYEAsVDaHo4nynz4MJIjc4pj6y5j+fjtX5a02
SunpKetr1RFcO6VvikYm5fnMh8guijQ/1gojB7XNP2eFCZ613Rl8n3fNHECTOJvu
FxUtK/H2bbeFocTgxMMY9Q3jhscvPss64pWTzOuSePi3EXjqEi4u0UggD2SjK1dX
zzWM3BexLu9fLNLsG/uEYExmineUVdAvacrTEaIe1LCdMMqQ3cXxD9tvd+FG1wPX
2UdKWsrw2ChpMqZL2Gb9nHgWwfXf0LyFtm/Wn0V/FBKU5X4ZJv+vWr5iV9/32FEt
nY/oEk/uuHdzW/xF9HBuHtDEg9X4F03vtXv6i0klc3iKLf1pGtaWr0rbW627eOTF
HSy3TjHFAKed7nVaVRG8FXVekrjTGRcEwzMTVYYZ12Q7fnShe2aUNTV5f0dK2dbn
4KM6OUnWPk2pHDv2m/B1Dy1VwxuTAuB9LxiVlt6wmiZHxqOvwUMj/te5syWxW71A
9GTEW899ME0VxY1TF5n1H75qdYBmG7CSBLGZ0GoaVYUtelETXZYkVJpzMV2Xn36o
bKw+0g8QP+uywKhLqCwIvs63G35sIV4Fdn4vBPkm3rUgd/0ES65bNs9ltRndCZbP
/upJqp8gTboymDHYsmBURUWtclY/aGzBrRltMDSksH/Vv6v4cT3JIeuTzZRAGwx7
jTKg162PLtUhxWs1c235Ja/SYSaBA1BsDfRgWslo7zstwR7s3ZwcSUh6HAKjEHT5
A4JC/7Kv41jrbtQ/SsD79dIIRTNbLCHCrUwtEAQv5/6I4kGUvsrNwQRx59blGHjr
J0WYvaEdGtOo5cVN+MAyzO6Mw4MgVaGRqVk64l/g5PzPGsJAun7UfQiWu9frSWbv
eFjNfpDsIXSUG4UHcN2JSvvyD04qRLAf3yQo76i25ntcosefDAso9cGPUgw90lJ7
MVPEwMijPV2Us/a/0FBHuanGDc1tjouiAvvE5aHTk6hViozhdeZ0SLRIKdLeN53E
6THTL9XgYvr/jxmN2T7mkamaJij3TRu6T608uUH8YAl4ejFdnYZLAxVbAB8GXWMe
RfMq8pjgQ/wX0fgwRhwcBNXD2mxO5PbgeYRVhhLO8yF3fTjx+lLaerQBA/IwMTJy
LpG2GWGJ7qWoOx+7LL31B7KpOdpyquoH+wFIvSixN5HE5KNUZgnxm47MSXpwVT2O
R9YzbgJ7+qU+lhUN6LkkeDGdpNCXos9lUXA6ixFnKcx13mkcm2/IZIsSWAfR9Uxh
u/WoKv8mNI1sl736ZcFlYgXkOPV7Oadyr/Bi37kg0v1INklRV2TWvc8YAveUgLiK
Bicte5uoe1dO+YUZXViyHvyyIGdMhG/CKMn0wLLa2XG7ETl83BTuno6RSmwZqu+b
1T6oXTSzUgCQQi01+Uoa0P2MUU40Zu6+IV9mgsRrMh87C4Bs6VG+ZN1g+xUh03N5
XiFArC0L/es3GL3wyf4GEfruEbCpgUcsjMADOeZsdNRvQFDZ8jwyYbh/ixYvh1sM
MsR/EdX468iY9pI8Iy0d1fnZZ4jJRucQubISTTJoi+OltKoy0Scd5bhGDOCRO1T/
YnT8Wv4lEIQRep2+jEf0p92n1kkluAUrrycyeb7Kd+X65GwYtqX5b2lnrsPYKF46
QFq4SSxaCh78IXGWECTKQqKw+sFvPL1fxev0kdNFhYn3be5Mx2Yq8Hv/8WYDRJPF
kasXMXygIlMKWeZIrRTobVlQZlZsrxzf495HUQrvv5/0tVnAdnoxPsEX3Cmu7F4V
2bI8vwRXBP13t0nNB+QPBc68llrS2MBw8+0cvCHCxbN1c0ocQ/1hiC2n1KfCgITU
XBWY9MODBo1TUyiW43KRFegJSdDLtpIqwT5PvGRy81LSUvikdm+DZrkfmeUiT5gj
WWS8NSPGrmv3DcgBaR4shXu/ytYHPxJLRX2Bad2yEh6UkM3VvUQt26gVTagQMkJq
kAks6QfVnjokTj9cDfI/m6UAlkM82NvMtBbyXU7hlfLZ8h07m8gxP4X7CyhB36Xg
NDijD1wtTemj75AtjaISXCBkoFljlN/W4SCev7CzRx2WmBojQqjZELLz2xvKimNY
3vb+Au7ghjEURcwl8OKPedO//HJbLZ12o2NNWEmUE1UFcOO8bChxOqRC4LNxVIQW
YY3vZXMsLywIsS02m3s++/HeUOxH46/XKVIItCFM7SptuuxNiAqyJ8ZJivCtpg4C
gjGFTH1eyviVqqTcb0hG/qTUcS+VlHk9qmU910VhQo1+rlsMIwlNFd9xhjdqRxBY
O5sIW/1jdnIWiJrk8MCWBfj101eTw5vUk5cFLACaa1BF2bO+NPVS4x+HeCTUttcW
s8jUwa0dyAvFWIz1ZmgeXWowCdukrT3ZO/FkYYq9bIwD325lxX/1AGh3TYXECaPN
nP9D7womJglG4881JmJx+cKhVq2votlL3Q5objZ1rsyW8pQ0NcjH8c46m3xMmqA1
DeYX3587wmKstL5bP/jPEwrMrF+ofOxankjnaplzJiRERHHdQ4vyB6zSGsIsj9BW
lGWJNNjDJ0bW8zozozTKscMEBkgVZKha97QXHAg/LXWNK0/nLHhgdXdwEpBoXI31
42P9YQ+Mp/vTJyDnM87sx0se6cSak16oBp/WuUY2MeGjrzBcKXdYXkoK6qgTJnPu
kw/R/X5eDFf1tbE0FaAlYkVEF3hVH0CXW1qvdxmNvMT00qOfsQutS4sG0HdJcojq
G3yFPMuPuL6rcWVld97gFSGehyPiJelxerUSbO7V2Y7DEV1JjPJFFjO9IvXUpias
NaMPECp9ms8NsV3HR6AVZY+SS/TtkTvuFqmPRqq/hhJm1Jl5JZGG4v6FqVve8Lll
2aiPUsoLj8PJU83F+37Zjuw7MFUyD6/fTgSo3mRAc9hTZU4lUIr8l1bnHJkL7lIF
5Bf16oviGM34Qd8GVuiOfvRNdjDWjwDE/65uGktWRXI+3bsybNo7+9a6PxuMEo9t
d798gn1vWG8nw8J3t+ajJ3ohfjL7yQQzTjdsht5tzwyZVlklkAY3MUTiX9WPEECV
LHveC/C1Cxj2TCd83LGuJqvZtNHbYMQwgv+xQyn/oIeo+nHhAhmnsQ0d+C7DrNyP
sqVTnC9MWhPTg0en0M1gq3h+QAaivcaArB4toAcBG4LPmrZWOzum7Blx4SjyL6/M
xfbZCYCkLrhdzs7BY0ZT2iw/7ELZDwHRQlgL5bkDeQ0IAOtYbwL9rUTQDikQW9FK
4Ro8f3R6bYg9nAnfKnoUdb9RWg8vxvdieEqJIqOXEXKEaESjNPZ3jFYFfTrEC0SX
NUwIqP0n6f1mTL8MkP7Bno/IUo3j/uYjP/RwdqAGP8kFcb206rRoyx2znC0EUOEt
NhUgxwRt2fyXDbZE6IXdnRxr7UabUBU1VGTL2s7r2TeMy2BaNC2ekdvWHE7b7Pvl
AM0xWnVYsFJ94dMZmGbayssW8dYL0E6SBPhLgmTh4ix5y3LDDiJmBHwUvkkvRTU8
tyfdmX1Fb0PuxJ2vnpeun0NJiLmAJYfO09hD4gJwYVZdZKAIA6g+T+8d4l1H7RqH
fskeuFUNK6djFJNYJP7OQfCxhPUNg4JTS+vg/YXARPsjoVayw/SjfnSMVjRQ9MqT
+n3IcUyRnyX23uA3gieeDg6Ar0F17Kp4sUBJIcNYSlX/d8Yr0DbLn2BplF9pKAPi
Q8OFD/M476FnR52pYMom+CipTy2KAxrSHuAwGW0l23QYK4Zrde5qkZ3scbjGebZj
sJIMPlo0AZPYc3RLpfX/xb0DLniIeTg9KKGIAxg1Sbl5k2ba/vliNgXjYZtDRYMw
2N3UElC5VfxmBX4m5vY04kP7Jsh85Ycojor0JsU+pJBldPC4PpC+mw0J+n7wwYAi
sfGlaaTgDdfD/u2WdRo8RLmPQF6TRq/1fOUrTanzM7fE/1NGaCYKGveClN+vVjHZ
9Xhg7rG0Jdukij/y2iauvwffdBXcdbyKTrWHcyTQq+WzDgXgA6S4hsdH+dfF2Mr9
LdZXBf73KJPwBnC4/SdKl3SAlqE2B0iCdSlbicRKBqJkicyucHOUleriZv7FzGf7
lZUw5Q0NLphg5AJ2Y6XWCpEPeZ8h3nW9U70VG2fnPS+0xZGnBvsy8HY2yPHkYAe5
Wsti+jN6kL/ZdaNNPyYyVKn/EY/Ssx8JcJDb0FOm9Ikb9Ek6+wHwvpVGNhiNGfPa
tj59KdMJVUjhAdpHFvg7WI96KE1yG/azolmQzOmHiw1W2954r/LWDD6dqugSvZC1
8lsFX1rwGX2g/Y+AfRsai0sKwMrxWbIH8aRSrINyB+C9a3TWVyMW/BStJcEGUFS3
ynslg3FrwlEnrHLq+fA0HPp9m/+uQoRKfruMT0cq+9KmcK39mMH+aRJFZeK7kcaQ
MNe6+IT+s5jqdkaWKI4ekFfXecqpcWlyEm4XQxqH2IirC8TGGw5p6VXS4E4kfeGy
aUGk1mgQ1/hpIgBh2f1ZDQQbXwnqSYwXFLVmlbIGW+Fou2HuRZa/SVuscc5vs9B5
LNSqAb8lcnTux3WdA09+xIVy8OkTW95eftdaVg5R/RmXzG0UpB2TlnE+5laYwj2x
kDgrv5rLlBmwGP3dOVoPJ/UGnANA0k+4VMY6V0QZjb6DlW1FQGXElWQbWjofoDTO
GKZIMWg8E1AOjb7tn/vNLbeZM202rhXxaSR28sUXHua1pddH9UdfPt2RXIIeajN1
pooCaNHtEHGBBArwDkzXhwSJr+jui6hTvXPYozcijuaTDE9N1sy8MmJTe3MDlBup
7T7JzZOM/mOAS8Z1x/g0LYLpIdmnpmbKRxE7u+JQvvGB8KetR+GkNLkMR4gQzuq5
dzsG7lnrfsAZT95idlynUL8PH5TrPpKlNWuHTfljEzM7FwZKGIWeRcfuQSUvuqRU
sFLqLQBnDGVAsvcnuRPjqAv3K5afEMKLRqF/mbYYHK3/r+01E8H3hUEwH4/k0+wc
hirrTTlQJVjoWKXJ4Wb6hswECubwuNMm+pVFkjAZSbFH1p95MvyXaOrrKCJ6f0nx
u3fQEWOsjv6Iusqw22d61/jY9ArR+BO/fiGdzp4oUTZGPL+v8wZ7nIYZuLCbp0nl
RGzuzFDOaK9LWznBfp/PM70nFAWfroYfn/iklhMxuCipOxUWXqjSjLYUxttazKFr
5HvhDGQ9I/yHYh264kGTjrvBBbgaRgKcCtezaDLgu7PnExCGKiZM6PtMAZusQghQ
JUEzQwehCP2TbzZLmlmHBe237VjvMMGOhsa+ax4+GVgYAgyAmjbrAizpKXj3QbS0
JWnDm6HLaJYgCXE+D4q5TrltxbKZV/q0S9cQB0ZW1Qq18tds8OViXKlGMd6HhgIt
X3MmrktkqFTtDykUrlgxCt68GdQAh0DTDDoKHMSTr6bZG+o3CanCI2KdmkcIvzWG
gIUZouJy8RYC1k3SJyHycMn0EzbPCfr27noiyriuJOF/Oq1uLiM3vMXf+SfTp4gS
nPbDFKciSNaVxRR09/lU5o0O82ZZHInHTY4bRoEpmtLQ2a04qCFgwADKsl/CKp+V
ripKkHg7dxXxPgnDKM+kn+DNTqc2gh2ofS4yrp67ZnrFqy9vf+gFEaqnYU0zw/fw
se7STK7HekE4+fjiydqg1UZ9w2Q33Z6jGpYyBa0kEdivJ8MQlqHyl+X9yiM4z/l6
HfGIAQIRQTbGIvVPexzw28Pp9ekmaQ5loZu1rZ5TaxeqUFD6sVpaiTbwHYbPIWpA
MBeOre+8RRRNAIXFbpNM8XMVSZEY09/k2KBTIE0BYwC1N2ciGQMe6UkEQrLpbX+e
a/O5KYPz4eK6S7C5joUGsN/F+5wTd7pZ0a/C7G88K72An4NI5vv06QdzAG5Px0O4
UMi5rGHx6JxU9JiU3ENhmDAUkp8gLLhk92owMZRKqN2mjATyYHu+iTurUg2A3vRw
owWzzLPb/GfQjWhTH7mjRNw3ymjPrt7vJP3TlEeLrsO2NdV8+zveNWeyAbqb1RYQ
sL/FDxSL4cO2OrzYftZig5a7fE2iRT/f1eVdNPQI7fcJ8LIl9fvGrDgUfyh5cDOl
aD/tSg83ZR4gAXH9tWrzF28TDSXt3TiAcTRL8r4g3SpYs12fmwz+b7088hS+FJ0o
irzCrSF9iCJlcL+tbQf2pvVoAGpjK3x01/O/YU5AG0XFk+VNMc3wG6+lZ8jcijvI
kLtZ9rck6qyRvE3H/LmXvTb+M0ao1dY86jidxnQ/RfouZd1THS+gEEevCukKTaRY
lleAeW9VMqVIQLOdC+AH4oIEGO+xGccY80h9jSzVsyzCD/XgYwCq7FIR9trx0fK+
Zvwh/K/kQ5nU/tfWIuTs1K5LPgbAFMEb/URPjoHjtVGMHmUWYvmElp+9AO3t0x6K
qbwfF8QiIm6efLu2pFsLrOs0or86qqgdIUKsRereBMi6EW4MHTqL5aARjSOVJCM7
kzYmDKChvR8jMZu+GeclSVsASR3NbiOwaJHnxhfdm9dvGs0gvWEnc9/A4kbpgfTU
9V/mlJV/s3AkMUQKeKfyNgxVE5o5O2P7B/cgU48GOIpoIYJYh6zWl0sPQGdRUfv0
Vr16xNG1rL46MuxFvj4ZYXnGfhKMLSLTcWIjrJRbAGDM7W/AXd9nbfe3OgG/tHP/
PY5tXq9E9m37FPq+MKbfO3TYp31ah+tYIiLT4EHevGxNsO7LmVjWb2lwuW3bvbPU
/SjqryZl+9BV1cbdDMPiySdQAO42WynZ2KO45sJ9FMtaBgHnvFK/DZzUQFd3/1IR
WuNCotTvowU2lvHTjHk2xq6sFcr32M16NUS/Inp/3MssI0O83mu9EQRBWuoTkg+z
SUisCdoEhCd8awrVFWJmpuG7ZmlGXq96GTXa0rULFuw/V2Ly60/bmpPaTqendxxW
6D1+3E84hDrDHoxfMmIPXo92d68WVcDSXp58qe1RP9FL+G9TohyLvYkvMz1gwnWZ
6x94AbqAyG83k3445D17ZlHmcRtEEHo2zzbn4e/PfAsHgIoYi4lNGP/OUNfPe+EV
45ud1zfIUAxLpbAtcuCVGreksfHLheg7x/FP/CQnGT32spGlilREGbKzHyEJ+DMW
eRSwoY891dEMCp9qHCZApYVilzY4X/lki21gomh5RzGkfHYbyiGkJgquMKY/dw+A
YQs+GSjrE6hkpnp4DU0yGjvkWmW/zDrwo6qtoUkq2KDm5I3sxcmZCMNZFpNsX8zm
1mIrXLQveCajYWi4CroMIaxjxWehuHhrGI9Phdrf/l/Rc/JoFQyrfZ++GR9nufq4
629xE2z38CbS8i/ANlr43n7aeHp4SJHWzqujgfU+RxNdcgfQJVtHZT7nawVHm/7H
buI+ajiE8l8bhTdl31qNTI4zcYE9D4wS1kK23kl0yY5+LSIkLs4Mu5T0BX4IK1pv
tQrqO0PbVckIjgJQdR9l67jikWEv5SszPS/hgWpySZGryTt2BI8AX24Vixg2jhlE
8bVt1mNAQps4cpuyJqC/yb5pxJSLh4QDQJttxiEkaqFi4Q952UD1zTNun6SmlIic
EL1buMNyVZKhpX1MBlqTX5djyvZ84e3OylK1FknTPrLZD8M8ybDEunRKFduud7up
j1vLC9hpYzxBc+XR26JDmIMlh/azjL7/5HaSDppmRMLBfiiHCXWFEGj5fEF/UqJH
TDhXJlFTpECPapOooUKS/9GMAw7M6cahrBxB188CEYwL3wk8JCHPECivWjjgutWv
WdigNmWq5hdeWuTYSGRLy3IfmjLAz+m7TrmF7LOatBit6h3BXcSbFcN0SJxy8Q9o
qK4bkLNxjipCINLQATPbJgcFgZoBWNambEg/50hjq/zWi3ygGdUp0GKXRP3pyjuk
JWJ0yKSMLvtIAA3BnJ3U+6OtoqSjCTi5oTX6340jkUGNL+JZFZuebBdg3gTxK9L0
9qfLLbZ3XMOqVx9pW6VDC1bjGY0MfOHPTemSXROasAIQ/P8IwNqTZcAGLqTH+pSh
ZpTCGLM5x2xYBOyqzCEEibRpj8P4hV9Z6voql2ryt8JqjcO4uxnNm90xGeUbI6Ja
DQ44YLEk3RkLkJGCURQe66wosGrNNMkfgJyqPv6fDAJxDS/i2C54u9lXAesTGnVW
BlTXolN+XRKeQgtCHKtu8Ugu2khnqfdKc2R3ZXuuxPk54ZOJPohiH6JAhDt9IuE2
NTB3dH6mIDiGmTQsL6ePc2dUEfpZIppAJYZNwd4++D2wCXIpuSHaNYoXeghmAMvE
L/OZMmSwdZYzsXh+lwE3Qn3glyJ6a+2XdnfYN59sszAjV106/iYhEJho1AvszmS+
F1ZFWUFOOnLuh70vURH0fYe5GPeLJvz0Glv8fdBh5iuhi8ELSMtphR4yoRwUactI
BUHQaOvHoX9QTPw/ITpMDwY2yU1ucIA/rbtP/lz6UvXQ+6pzJQH0r/VIDIh8dJYh
t5PbFcdv4pCVHj+bw/VVjy8Lxtd6Ii+MVxakBnSkGV/KI746I4ABKOhelGw97fTZ
VjAqbOCRg0M4p2Jcw8jjWFra3d1lVX3h++VuKHwVyngdKg9QkGsu4YcZAOO6Gq57
xA+O8EyHGPc/5Fu2kZG3lYPHe08sb4wKJe3TOOmI0WMucRNES0fzSXwLmUDoFr7J
Xu3LBgsU4QtxgpBE2hN0HguQS9qR0ZoJf6/PzfFx7BxIeydvR7rdtSPYAmx1/jtr
O8qUkcVgK8bJ/2M3qmyf7Vp8LkhIqYKzlNW5tPieKYAqRLco3ORu4Ar431A3I3l1
N2FlJLJup95GuVdAvgk+E5FpRECdozhbJYQWH+NsL3v6A9BtMzMgB6BcdPoj0g45
S7ebjPbE4Tao1H+KInLZ3Va57mdZksACVL+ZYABI5WJnAiVhH/Ha3lNyT+6XIRJV
QVlHA569Q0kEjiV3ZdCm6Dwmrm2GLwT/xjUz9z8rmc04B7D3TQkzuNIVB8ldQsua
TzGfrVy5bZRyQBMz2CJCirxWGBPDHkc0MhBK23KoseZw3YbNCYD3yd8KXf5sGFSi
QbLmrFJ43JtWGmQ9yddZwhhe9oyGaqWoNG8l8DfWlO4TQBFORxWNd14fEF6H00VP
7UasrzZm1HAILsh/U300ZKjizkeeSWpdQK+bHrDotrKtf6doykk8X74tX7ywoYPq
Wc49AWXdE6ImWvzG+1LXQG+KE9ISZXVzReMNdJYYexXoD/v30x/P8wWk9sAHo1kP
+nNStOhLcGXGb0KEfLmUeQcYSDKqxe/t5cP0u2t5+dEvliEidqyVlq7yPExmgYvf
WLuLHjnYi1N3m7KxRAjgBinUpxCJgrKLAcLMIK/b4q5hkros/wepUmt9dzPMAlcD
ucZFyn8Ngwk9GGsln8w+3VkIOceRrQ5G5Kj4IzFeUUTz1gX+b8saMqFRGIPvqr/H
3UsP4SLFpYY26K4FPV+73XpXq/qjeYrTTqgEW5ZD9j31DtJiALQ4FjDmalaC8ixD
rM/KO1NBYc2bHZBi+LQOGqmRqU1Mro0Fn5QmENxd88dXxl+kvrNu0MJHiMIciq1w
KL6TLpLQkjBsa9Gb1GiXpJGm1S3gS8H5CHtz22PkhaCzDXviGl+0tRYZtpGXm0Dq
8ZHoxa1zYDeO4bY5xn9PoHbMgCGrdllspPtz62RwLcD5cxqPkMxsKT4e4bhO4rUl
GZkW1Lj8+bJhscFR+F1L2yCGbVwxRfHBLg2wLKzs+hPxtmMH220m2dR/lv102D9c
lvGEhQ7TBllRIfN/4s6/jqY+ki52AzYR8tk7NaUFyU7TsVfbsweu8futngAOGMlS
7apaGtjkmPxXyIiJZ7RzL01HoFbmnQRYLdD6BWmxDqEBaFR9MvxCMx/H3PRP2Z6A
QU+YT5QYQNXmCdTLjKy3pTxGCmSguWeSYxxZkrUrtPcGh2YuSpY6JAbmQELqbfi4
Te2bpNS47UGb0u2JlOJuyA==
`pragma protect end_protected
