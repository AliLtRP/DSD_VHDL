// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:35:51 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Wq/8818/6MN6iEdUdkkMP7I4ge+ejVdFLdnTMrGUB0TuKYezNEOHIP4MzwvR4clx
rV2opS951dTCMS/80xIxYGzWrbLLD+e5/JFOIN9lUAqU6ClPWkPAUoMNP4v5dbpn
hBnuXao5Fbgj8m3YLwGpKnXy1bREHvReQDAlADBzrJ0=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 3920)
iM1Dwd1vuyjpqS5ZHd8nNqMWNE6VKtjckcQQmXEEFBeXCJlC0HZSTfeKCoVqN28e
IW5mfoZHFmZkKnBiIsycwmQrqTQP3I6NaWB3xZSvP7717D4swoWLYKvKXRnUCK7K
YGzg1RV9o90h6iD1n4P7jQ9znsm7RHQzXCzfz+z+k6R3kPUMzDaLPWzJFItH5KlL
YQTHVIecJor3+LOKfbz2TTpmXbDolBhXkNYmgdcUPs3E0A/cRLT862nkhSDnYIIy
O8YyCyS7jGACDLA/cVUTuKPjvCPzkMLGRyR0cMqo4B2ybTmEb7Gm6gtaO+ATltn1
He0KxHKva+EkjMlY+7pJKIU6jYRZYkSQyOBzzNKQzIAv6Tdc03EELIdatM9CSJUw
HqRlgvrvhW+Py7B6PAw3ITA9V5Bkgh1UQgq05FdapOFAxgntZKz2fWaHZi70f4TN
e/62f+cccOoohpMEt8VVeA1nvINexzQGn+xH28nG9ETOr3QUl4veVgSsoJMpTxe+
smZdk0J90if/Ibfa3WJsj9DwkBjf+6AF745Yyd+V2SV8IMjUEjUvRRZBu9RUdznI
fPwZ3Kc5Q6Yova8epWQ+tFegYxnHFR6vB/E6sTg2DYRQT+fA7PyZ7nHdA3W00ZA0
8juQ64ssiIDpjoPTafoHQXtYL67JGTtCCcfOPHu+vR0dUCH9Ie37rVLPU4aYBoLf
EWbIPRnvcXd0bAOduUc1AMtbk9n3mHmMFL1yps13X2r6SpF1gAieL2SoWgeTeLw/
2l0bk7ifZMOxtWIcfQpapeVkMYXu+GBC68Bw/YKdODdrqt3RMnQZ1vy4i+xqS6dt
x6Xp649/uxSiqF4RLZTqKCNS9Jjr0KXHKFXqlUAcR36DQxG3jLGHNBDLtwzEBY40
mKBfgaPZbSJbAQ5N2LnguD6aYTpHUsUViYhgfk9bKNoA6p6YyJSW0QGLXRKi/zeW
QWRK/IT6PB4ZcGPn9xtGaD8OviTnkf+Wt08ZIPBrXCSvkKn6x2LAyGQu8pelW6Ue
m5ABjdb3R/dHVG+WY62sPQF3LF/c56ndccO/lYtFs7nMYchDel0aW9uhx2ljDNfV
CjkEXG4LZSivJVJq/uV4G+7WuGFzJAU/dyenGvCvF9FH7Mudo9mBjiInUz064Ci8
7SoBdZCrBgZeDha0j3xkFB5yal6mdI615c2xxgDoGZ4qDDhrEOl/gUfBiAPkQZ4F
PY3+/jEhZoLGkCBPb8N0FxxVV3gAuZ75wGNc0kXDE2TEIb4yrahG8oLCOZKnQR7D
j9VwIPTkCqOjgY7ZqlUTR513a84K6ACbY5AglgGAV5bfqw7hnbYjhIkc9E6LYIQG
oIMRpl8tufOlkaeFMW8j1fia94nvD63bKv02FaY1IvR+QBTjNl+H2Zgr1pOljctX
/ij9/86nNWGzHqmSoVsCmgMUIAGqP6BaIva2o9pp5BqEesDWTs6gldO65CbmdX5q
dHhSj3E5PNxm9F/LGzBYcY6esLHsnEn3Zzw5S3WnBU71j7/AUMi5UepISnJ57R1j
lmQbNFKIxWuhn0BKMlyufpQVlC9g4eAKZ22U3Wq4QkzRL6BPXYHA/fkOWUUOrmqU
RY+lbs0bTt5uU29YGLOH8smrvYXt/APF+JcHgzMGx+vahpjhUB7iCeR4f8Jq7Nyv
6vcwN2v+o7M7s9l1nWD/I39AF1aNYeXyqCWH4l2KAWUhcvbboVpSOHnKZHzmfFdb
XQt6bbdmgWQ/93iDaHVgC4f/fmq8t2zIXnRgvnhdDXBTpxg5v+zQVhovHqTnuDFS
rOGg0wOtAXn3/+AT/hLFv5aLVtRFB4t73sEJyGe0DFRWuqWwQ7yRLTftN4jodhSo
LuoD6WGdihYw+C0J+SOK5L2FVhnH5cJzYTBBko9Tf7Gy3hfMwT3wEWhbxhtQrf1x
AUaHBrMG7t0fdl7KD6kKyGAnyA699kQpJb2zmrDR1jESuZLj6xWHNGS+kHlGAID3
Rsy2bgoKybH67Hn5KuI3TSG54hndfWpf11zQ4hZXXnJcz9QdCm9qCELxXRUn6dGr
dMYDO/FoXUrAMKBwG0wlTM8iLegr2JxwouOBYZ2euAmgO0CPCtOMAfZ5xsmX5J9Y
YCb0VtZZVESjQ7qrBS9qASpu+ucVcTF5D8u38KUumjEfVjDy4KWi9R4GndCYEXUt
0zYsQkrk3e+VQ2CCGBnTQHpcBbh/6rBQPtf53WUP+3+n0gQWdUYsU17kOPhwwVMJ
UpCgvZwBwOCPeeFGTC/qW0SmEvBZfxQe5PGIsgTqf0fJ8huFkb6wvNsuOzuspMT2
dIXbvoJgkecWVT9QDOWyLjvTfRKqmw9KkdYULrw5WJkxMCdQvNBHGIFQG5w2Q+xg
UhZ1n1mtawOENOiftIOYfR/elCx5PSt90UvsfotssudgbeDk3ew+93BUdn3I3Qgb
2wDoK3UF1PZ0KAP2i1dHNdEjfDkDxegIuIIyzHu4Yn45oeZOS8gUttqakZmeOi+K
/etf1tbK5dfrZljeO2dzH/hJlBBl838ahxx7ppfjJ69K2++b2sd8pl+lv9tsHWK1
ArwwK/cWthLUO6efBt/3nhGqVcM1pg00QI2zvTQmJirR6NFOos51ZCmKWH1ZAeP/
k6LKcsImCl2KgxK/hTdIq849Da8bcSiLKrNVg2afdJ5nainosFKTre44xKiaczN1
7TUcDH227miRjYSoaNxyNnDmEgK5i/5aW5rmW1TuB0di2w6CubzoMjQlHWTpmyRe
rQ5NWfZ6rrbVRcGHPaPZvdoQfjPiX3rqDTZLCnDzlNoNctqW7PJz3dLp/d6odx6m
L1sJRaGKmWSYDk4ukZDtmCofxAbHT1BfSeerw2AexWSpmKS3yvV6P3TfJZ/LwTek
41DF2m35kwa83Po3poEklW+qPrX5o5ZLMggOkN31Ra+jN8CDN882284OgoF/K2jL
BeYvq3+u9rnB3u0KwyVcIHyljTUnusaGeFWTNunnwBLMpu+yJwtjH09NvHo8SqSh
RvD7Hyuz6wbVA9aEZVJNQY56ySHRS4ABh/OxqXVmbSU6Lc0oZbTrpBQA/oSjl7PT
y4QdJM1bP0OYmgeAFEF8L+zZSHII/OSwluL17R+hVk51MVb1I/6g2TxGyvGz44MN
JOq3p1AUc8ZJfDhcRPCZZJ/1WUxvstKQWQkyljxa93OOoIiP0URAi/YnIYiCnK6+
+/GngJMJ3zuyvYa/HjcXkwYVQHggypu7aWQdFFiK9uRvGE0YE1Gx7IMwY1w+83kp
tGtv/Z3g684L3V6FJD9pUpSO36ujeAJ6Dnvyf45oZMW7N1F/3rlUOjYrQ55R++55
5Fj6zufolcPGxhc/bxzuBhLlNF3GXIVIdKSyg2xW+NxvQIAeN+t4cBzW2k5iKM5z
5qCpFyBlxlkhx1+OtdOzyAOFnhWHQ8KzEzOAXsTjPVCrMF8dGWqhUQI94wS8zeDF
NxvmYuCPQYeinVb702So9J/RNNIzbGWLBX1eqSoBzNwuL3A8ZAYH9t0kN7bGTOPC
vkk/mjp9oS+7YjkIoj/qncXQLFeYihflBIHexdEh4OzwDavqZa0HgZxeb3eJttoP
XIc69zMYK9NCJuaU90dhxDb/LtxzRS6VLhFpnG/E1fBDZUz5/KuocEMH+4le1e1h
DeFrESIXEfpGeZyanR/pmkyHAzRxjmmYdaMoz/llWN+lVifkiEliEZ4lNhf7x4AJ
ltC27+fDDDo43xCNBR4ujWHaAIiSep5vXd6zSWEUyBL3+E7TvKJM0FOMNsW+0/DI
1uAtToYr9e/l4cGKzbaE1UiIOekUCncVIFQYsuXR45H9etLYcKjQdmba8xAfxWZ/
UzxmRzlr/wfBuG+ZTHK8mqtPV+L0IybQ5vkgYPlR2M3845SZhm0l1+0mmAf5R2/D
D8lQoo/ps657WhXo8PTp6TbihvQhmyf7M5Az/18IXbggK46WScAOR7czGx7n14gt
jeb95ZVvFArlgjUDLRx5PhVdmjaNX0bhCmNBxhjGdggY47X68TlUBC9Yb3QpvI8i
XzPFmRJmBHyKfDKq0XfT/2/KzReQbjBFI6jHO463rfSH/Ks3J3n61EbnR9yY5+MH
DvOyKgBi4U+EBUTRLtodqDv+ZINcm8I8oUkMUaKa3TnaXDCslHM+hiz4vayxFHIt
8+Xb+306OhMn0UFiM1jwfRzWwCGB27TvcKyZ4bWv6y0UJ6GnYQA5ToK6m0eNGI7J
FqEFBs0qnoyHxJ/D/AdhRjF6idt+moG9HvlAzSlh6X6HjrimtnpJrqoSOMWEH6Wp
DK9cRQ9nH8W7Vv+57OSwnUBIJjikvnKCbImbQUE9z8TMpZg2uATozdh/u3FQVdIj
fHVWgyZSAJD+eIKr6Q8NJwpiP+OsGNmvY5g/s0X8/h7GHWcNPfthfhZoEDn8zmtc
3SgNx3HOH/4wFEJAPJ9hwOJ6XBxNHiZ0pwlpWYaLR68a278BHRIRQMWWWHcfn2FM
Pc84T6fn6EhINuAESaw+/fPpcHZzoV0YvG36rfHio/zuWf4qpvuMhYpQqgflDQ1s
dfth3fjGvX4qzzBQTT2MuulEIQWE7HtJZ0sFmi0+3F2yjNL4z/uPgwIvJevIiVuy
XwI7BdzUyItx/GhuxW7MQOHnah9AUrLPZfDh3pnYtpLKS1QV0yQjgIGP9fmD9ScY
jz32vXuT47ukMaoKUiYrM57PTfUM5Gg7gC+vxdU0DgyzrlutQhrBeo2X55EIZV7K
H5VtOeFhhbxQD2h/9zU773Djx8C3QV16i+V1qKjvduhTVUymUqpjXYJnlfmLQrUo
Pr2k/9Z9GzQbTDIVi0CxkvNVJIEM1UpFv5lKG21u2S3pO7/WBDtXP4bjaLgns9/l
B0xEb+rvf1z1DESHmBIl+1W4YEy2T33/GFHTBfiUPsLH5WkPNRN8RYFQ93y73CfI
j7XAvvSR/pZVvlK5oetsD6Wb1gHXCw3gv9v9Su9B1pBeFySE7f3IqtSYHVfiEwJV
d8zLvZhaUL2AE3tLrmnCok8UYQ2meZ/V/JlFrsJPDUcy6LAPLqQxL/StMWQRAQMJ
H2N1nZkst8yDE9cQehZy1fusvxK6gP8CSDXY+uTS9CvH7JfN+VAyrXYuQeedxoyz
4QhqWRdjOkfrKOTJqwRoY1hJrKyVNxpzTf2KQv2mSPwQ4q8+0INKSbLjQkPvKhQE
sxE5k8zqa1RnuczRCTJaDdYKm/jI9FNnRDtIGpaHFiA=
`pragma protect end_protected
