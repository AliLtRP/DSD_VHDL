// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:46 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
WghHpF4av/2JqSRtuiryz0/pZSlOzzbBX9wzXrMSn4E6N26TGRp997/TayJrHiVK
rjaRMVZTDqvTr2U/gF3ZXn4CYI3rQ+VKgr4nqd+i7QgctsOkCmQyg/blsqER9/xR
T8svjual6UmMFVmXyko7r2VMrBxD8Pwlt5OMk8fNbCk=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 47680)
AaN0TKQR0q9AiYcGqEtzITy4x3Z9w4hy9PpBlWNYPFXeEDqY/VJnJEAZp6E7d9n2
a7ZjEFAMenY5e+85KaSKSW9yi45nNI3PaGphK9RKd4GYOk4vHgjYgReRxGlF7tTd
UdXUU7zfJXKOOsrBWmT11lGqsne0nrj7aNo8lgOvi8xLh3bSE1lg91OSTBLUXlqQ
/Tk25k19hP8YJrFWwUawohvAOTDIPHVDexYJp2CXSPTKjGbouq1flo/RhL4q8DHA
707aRuhUXHXZSSKCYLcbHl5CvLuet0ZM/gr7S/DmGzNPo0Nr8dW8xLzpaX5McQj7
x4DNGxd9Tgr2bJPcU2C7jZaQa6bNcxGy37hexeZyslgGLFGuOQ9qsX8HbzmH+sb/
YJdrEyRc8jz9rEl6Fe0YmGUZRkymhaR/w97OVYjPnuKh7nFLYPr/JODNHfp0o25S
/ChGc/Hx3m7mczth0GmHRy1Z3MUguD8nfL8YgyFREXt8lwrADFlSakaMmCdI3ePK
3AjcFMvXwHv4zGAOvYoqlqzs/zzBbjdBZ3O9DMGkVvCU7F36miQc2MGHU8d82zUg
Rg/BKaQVcRE+3tVF2d4JZcN/RG15hzz/HTFgHpjgzq6A7Gla5L5cGwsvKkJbCh6H
LCUOw7++3RavTukg3VKHI3xO2zuZzrcrg8hVEIvWD8mN6ktVZL0WixzxZrdkBIX9
FiuUmanyJ7wNYqe8Fm2xlB1T74rwN4XIdrb878MjJo6lH9XZrTbohv4QpyemZvGR
AqpUnnu9oqDIeqoVisHjR3fKyWHeYeqWXKo2rnlByWHEtjA+IHTS6fvCfpFmI//f
vreCGS4BuhEaqXml7WOBdIof1evCk8xIU0Cxget4ozR9vgqOtZ2eftpZR7tXCWL7
HCpmFi5EFvjphq/jleodqKWlKUIJGQUhlBtQRY3wXxRR1/0De1K2FdDteDI67BQt
vJ+xEDygYf3RTd7/ZCEkrGF8MmRqlQh/v8u7p/Aypcb7HUIPuUosaV/ApbW9XD+m
1EQhEjPVW24Ql6yFI4B1FJb16xGpuO0jc797GDaOU/W2MCrN7QQdAL++DdUJjIOB
3hlWyWZnBheOzsdiakfep2KCG92Jlqg7wWGDwDh2RIGpt+G8wIOx3ym0Eljvk1H/
NAliLkGg/rRpJbB/dihncRi6oIPbEj7eifKw1tsoo53vPwgc6lzEoRJOGzezOS2p
3D/M6oCTIXViKEWhUA6smcNmmoGwCXV6fJEPzY4RQx6QmAb9Ozus4DPfkHKZKnkl
D+i193y1GcTdMbAOB3omX7YYx9u571QRHa4qJVQZOvzbhM1lqBDado/+zQ2tTvRV
Sx8cLVmXCLyv21sWAUI93MI3yTN62R6py/Plb6jN9uIT6PuIfjKNSjFpTtvpSlaB
81q8z3GxaPWLzxYOhXF2mfTVTwgfCMM4WY73846wzJbgEEBAC+mRouMRfmi82Yef
52XV+fRtB6vpxzFQkX+ORU2jdhhdCPCjSybdho6HFqGvJwzWZZSeBoCc0pfaPg5l
CBKFwI35QIz0kz9iuLLnnfFpPKP+EaRNKjay2yd6nWFyp3LxfDIn+Cn7fgj/zt1X
3/73Je6OzukEhmKpPw1+rKAKspGMd4/+5A0YSDQB2UxEaYJEdea9tq+g1LwfLsHR
01CUzk6KElEUKhr+xwnLGGH4wxu2tmKp0Bx9pqIu1WYN8Bd63qB6garP8Mi8Eyjg
c2x1NxWyRAsbV9JgZqNF8RBylrzbnP5o/ev3HzxRMGzB+z5xAkvWaek/8hsakNCo
zytOHaSNB4015E1qDNdErtCcHEKdC7ODuAgAz4Ht/hI4Ds1Hw63Tcs+0BT83/fSF
ujdgOQbC6oqIiQYddBiXb4xIot373bWzaV7dgUpHEx/BpZ1n8U7V4nmuZ0haJTMC
n5qwgT4SvwJl/8BMqyX2fDLw0j4duYyCVkw8EEMvK4AR7wmwPvNnqqTMDDcd455f
O62w/A1HeAkKXY2iSfCkPseLGz6zLuCkqpgANq2e9j0u4luerZQIw9nnQbpPgAZu
o3TgEU+cmPLnbFjGr22DLzXDt1ccMyNhyiKae/1kHFfzhVixfLi6ErBVLYt2+vU8
UdgT3CzgF54ak4CnFEFS6tZAWdTjc9oPu+rTBZsX8rBj3SLqhNxdt32WDQMqcey7
AisZYPHFPyxCoAVlgK3AQ6AhJ58XLRWbuaiMSU8VmM2p8kq9sL9F/OH3xqJVjb/G
t7OLkZ8VOuf89zz8KTLzxj8dVGg3zpw/RrH80n2JntRxqDVZq2ZnuH+7ct83klT3
+WMWB5LzMWlCQ9qmAXN8ks0m6KK379Ci+ZvqI5zap2aL50qDqzcjcCG+NjlwNnv1
a2hUYO/bk2nBte79w6CZqKtG75aOk26QLqAqwi6qmaQL6Om+UvK6dDS028ev1n9b
ruJrnLPRrAMdYxedy8B0ugLGRmNeXqVd0ckxNAORVBfqj+o2S20Im/i9UULgnnWM
NEyMI1RXyuYdfX0/nEaD6vlZP5FxPMEnauFL8UsV4aJTb72PcgTunUXz4iYSLBsv
oLrEd4CAgXlBTgoURBnnWD0G4b0dqnCpGKef+NZC+Px/oeEQjuT/Klo3BEx4AH1E
f6FPPyDVi86sbtQAaAtRTRZm1MVLgUz4hwseLoOt5BfUGfERcZEMmaKkoPkkdJsG
a+BQRhfAy+0azTWX0jf4vw/Htp1FyJsphwuo3aEG/86NqvzlLClWzKka9bsyni81
NTZy0I3E6JWt9AM+QEGSc5RuIke0Xk4aKEexDaGcny6nIsqJ8VvnwTE69SGMBcK3
iKLtaLcW29YKB7tWL5TGCYatZX94hH+cKwtPcdp/zm7s1ZIfsoXonWRGpIMfkQBs
KNpBwpeAMM39UFsdz94p093ifqrVu5TkI7gNB6ozJvl+j4e5VsDtwrnpchcWrcZa
in8AlyZYN5UiuwwFMPvJyQk+GtSDK9CBmdjoDU8RTNlyICr+CVQ1kC9yWHsJQhW+
YA+KxbEdO2qJ9dbQIoc3o73ix5Sffa6lxuNWAgBVQ8UNsd21CDLz1uemecmeyeiH
e/x/kp/mjSCwE0QnLsqDB2Q6/1OAuw8RcJpLs/U6/hsYGdlfkaJvmn69/0UqONDf
1ZDNVn+vDenFw+9Mlb9UZhDkpG3DaIHIjUIPzi1fWx7RQd61DHxmKyb1ULQ6mksv
krIRW10kR03ww+771MLX8IAVddrk1vkZpKIaVcARVa7sZsbKHw31kB7zoPFas/cN
vQSeDwS6kzeAAyrQ+6AftKzha6uHUQG9foPw0+nrA68p1CUxw/BEeLYBOQrYeL8Z
3ra8Uhts16yPQt4hQeVvZuA7R2f5dmx/H6ZuzHCo7yQkVG6OkOf/19pCiHMD4njr
s1TRgK71X5Pn+8uzc42cueka5nkifKaL0qLSrsOM11SQS3esS1GVzWntfu2+A21j
xsjbgDM3j18GQ3kULI/x02fuWr5hv88Ncx9+EYXCTo+7PS4gZlvSkW4KEGf8oUJP
qQraoCvStjsWBvlF0/60cFBYfRS3etL20XD4OK6VluvQ780Q9muz7POnuxUg/g/f
I+fxJpy+XEeGnCp6wqyjRqTwsP9Bl9VuUNIU5nw//+gaWnUQW1pRgwhvwZQqSSPh
/kD4AMc96c+aC8lAZeJ/9EhA2u641AOScugwpOTkPbcD6r9zjdORCug9BunTdpn+
KvB0wfoRYGGUIVvIuO3lQ/6VnqcbdyqOSiPx4uyhf/mJZwN+KfTfrEiifMshTPP9
kfTc3CVAAYQrdF8R/tgROhoSvIyHG+pC26ylpFt+sfLvxsTOyt3Q+/HCjrUKDRHx
QbYfxZWNU/MonRvW4z0R7RU8zksyQRYPc+LbRuUvx8LB2MNhZPTuITApCncXoBT9
zZzPltugNoOEI2GBunXby/aVt7WZ+WzBQ7EGpjne6LpbvZNNnHsdUw5MKr1Vuah4
ajr+v3fp8dnNTU7VSnAWSIuCBHIP+HaDSkN+t+ZHwNlmFf/V3WoZGTAWvLd8qOe4
fBYyeBvxdGxGbxaI3gPLgN5oG831Zccj5JzZ2mCSov+1U2QvB7XmUi2or1KwhBxL
4RbjWaHJ6TaOpfMZSoofe+Bk+JQuWuY6c0M5ly1YyckySd8k2agcebnszRJtaVCu
pLdMm+apw7CUsNE8zH1Lc7ytHniRjIU2RywjOAV7KZ0GpNUgEoj95t9F1sIyNx4x
0JZ/xoYUx8tsTojH6ZVVm606dCqiSyBTrDVMU+znRdxmNgw8LQ/jknfUziP5w5ls
hXWGvkw4q09DlNK3wL6MW07wqjDf7KTzWyllWTUlObqpV7Nmy/4VTF1JkQR9/Zmb
EFc4NcKHsgLVCfXhzk/6Au3x02Zw0xRobVITzkvTwpQtG1BNzS53zorluz6gA1qR
bjSZicdc8ugTQN0d0KMyJCLpFCzmDYiMxuM/Z/zw9A7uqx2hPIHNqq9D8zsByXtd
hpw0ZTp0TXLRd0Rvh+kT4rJ2p8gcBuxzYFDeK44pUxKEjoN5k42+2rS56uKCsoYL
Wb6FtizaEhYcKxRt0tPUA113iO7FPxfqPlE+QrDuMXGnRlqXptUMhMJQnmGaRyIo
g+lkP7b5+xUVnjJhYK1+tHWF3dCc+54emlwsDjYMjsDK4XM7C2F1N5z4nQ0yTTC5
/Kw70p5ZnlEuXtJ5dZSQpXnDilwMRhOaDazikYDX3VM7bTuKv0z1qT1adpg+FY7/
5xS66PyaKEzaNyTNwraXoG4Co44MHdsK+aNoXAVY/xKRHmctb8caB0IN8xI0xHlY
1iISod/XsCnrP6QWdxJWeYdvvegdlIRFS0Kx20iroPkCY+D6qBobqPUMhimuhsr7
YiuufQ2mL9wVg6BXQBkvKr17N1qR9nacSB2Nl81ZN8BxoVjcrYRSDDEPxeDjUumi
qI5KiQdPEugEUver0ZbIaiVokhH63N+3ARTaAEuVFf9jcuLo7zupZOPe+KJRTtqe
fVzkti8b2k2KMwuSHcz9CbBzuZa81VSusWV7AdbLd3mx/hVXY9qgwdFbtSbj1Tbn
4ywPMu/Qm5SgxA67+Y9v6aDDxwmOneElxqD63MtjR7bdoLo6g81Dn6ri+9Sy3Eo9
7STFxoRHhu+7e1yGfx306B8IGzW4L0dD0XYslFo6ys1IVWw/Q/BBZsXjCGavj2z4
/9ot1XIT3XqXASookIUOhswJn2X7Rve1Zh+igZeqUx1mMk+93/QFfKbsjRWrO0RR
kwGofxhf7ok5TU8NOtLV6w9U/QMk53kolmZh/y37ECVBMbg9j546pRZ9eK/Iv+YF
qGva33Vxc/SiS6JhUBof/gmd3aZBPjfLnRP6Gn+clplGffsDEBEE31q3vJfzkLkU
SgdY64W7cX06+a0vTyPtnZ4KaETJwOVRBv+1+OWSOkiV6y2IRGwzzewD7x3eGPHs
jGPgAf9byHzdUElvpvZl2nuZwVa16nEYXFadhzd7O44k86+hFokVvRs4ajOIFHHA
KkK+XfJZNmCTkESMBrLontWZ+1ny9Rpt5e6380jeRafQ5ugve6jOo+GtBSlZiG6s
9yAGsEReGqnnizHKLOFemrAeVJ9H8iXDsamIa2O2P/tR0S6LMXrq9qpUI5rjSuAS
oBsghQhRK9wFR+x/hXb7tbj86VJjfoZUExgrehnS49HIxz9ovXefHBBMJtgE1H9Q
kXa4lPcmjz4g5t7ctM26kpHf/dA0EuLVwk2VegCBzf1gYvUuWRjXgTrtIFmPLZWT
TNduttluiXdl3GDZJVDh3KBTYrcgWIerT1QoxvOU+dSpV3Lng+LekQeLMKINhGdi
cN2kSKxgUysfcySRoi/FU9qehQAPkjLaRF/HxvmuwVToVTJDkRqOYl2SoLT0tuW1
XI75WpI+dyNfBcCKsw5ObUmv39RDOewLzsll0QKx/hnOBKq4cst+q9FDaNoXKQvj
QX89rlYkuB2m38qlHnwjzd4c1lzTO5vEjOLXBqSRuVW21C0PLRa6WM79ivnGVrtF
JzoUQVG0xRZ8koyHaInopZmBNJc6haxroF5TxMchiHmmQWAZT2gf7l8d2idtGsp3
/fuvGqbqYh/U6+O0hAoCuNsmuhjIKKo1XBxE+2oFc/N84NIy1jGHCizO/jEIplVP
LXLyMTKD0S/5HIUt8wnx3GxpV7GIp0MfoIRsE9UOi3sYZ6OdCsQI5O+9QGr7xoXq
h505lVqNeWwhI76ukBKaCarerYiBMdcW6iJUl6yIIFCJS+3s+r5hjooDlUd217D1
CMjWrOa1w8krv2SYqk2mpCsNVt6ABXw5xi9f+9zBAXsKwl+R7K/EBaTgBaV4Zy69
wFjD2gBHXge3k6h7CjQr+efF9j8O7uaUcAZGtduBBru1myM+6rbsxBzS7ypobhnS
AsIosiaEd6tTVH8rxwZa/2cZbvgc2wgZ8j/lQ/CKRAk9BTV1tvSHlVYGvntcs4kW
yHW8RkoUdNc4dRRIrie3oymvR1QEp/WfmT6d6gklA4sJwnnOWno1Z39V03kCw84A
Pc75WMSA7EK2dd5WxGldoQNEQu90xJDEPE1ppZdYIM9I3VzNwbx1qu52iPBpJ6CS
3Xa2D0gwBrq792Xwcg1vegZyAHCDGRJfDXnw7XnflIE/TcTZhfjtVfLlgJSMwUyO
XdQQgCP/+1oWRV3O7bQwJ0IggPqDijFol7RNeUhCfXZ2g3uEjlrM8MteWYrGeTff
BYXwmHpWm5wqYDf8acdscFKqn9ssaF1lKS4lrejT3dKssvrXcGNzjvvKSyElJbVw
sbqmOL34SRKp7YfwG1jwSQyeI2fVZ3BBI6za3bzMVfo4tinELJWGWxnCCBjQRxZv
A+590f0a3gTXioMtphk8hEj8+q1UEbfejyddEXJrlIzfuAnxC6P3U3dzMwOrZ7mN
yn4hdQe/00+uPRutvt6UrNNUJpo7eWv5EygPbVpPA3hcEyO8aV4dybOCVIrZJKsb
TRv7QjZYuWhgezW78yiroWInvLYCeZVPyEaHLzSTHz7n1dWBR0SmVnsqnIMFktBr
XIXkeww/1jSRIdFphpA4HQOv21ycC5DQJ/0f+LuKbTp6tR8oA6JNisVrk+zgB+sb
QauWL9nHJCS84/AhQd+X/C1kyfKHYejcr/4zNjTwC3yC2cRjYmAOB2ad9bVoeEUP
I30onm9c5P19x8p3jhXqtH4VNO4Zyoz/R0WrpQPIeW8/Uj+EOsUIXOpI3KUkWgrZ
rIF4JssDTgx93kRKdee7JbysPP8kyaCk7E/0VPOy5jfAJSc5+AunBfSd8FKbJ5la
c7N8TXg+xAmD+Lf/h9sgn9IB8/Wgqagr9XLJbO49twGJI8uHYlVz/lf+3ZNgiIB9
MOyp+2LqiQtkm/1a7OVtvI66gwmyM5SOnO8+mj9LLt090y4zHFhwT/KGfHN8E7cY
afT3+K1opuvJhkKZmH9l0IfDvZZtfaiOjZ90jUfSOqjHbcF4jdJVMM507x9DkjYx
Ge5LI+HdnELBHEpwvqp4/JHjF+rOvf1XSvz179jc6f1jMux/u0zN3k/2HPN4yaRQ
x4N9S83V715QEEzH938htGFdUBas5FVWIOX4NavDVota9Ji9FIrga1gp8pXT78wM
D1WTZY1bfRAiCDfftvCnEq/ns6DLbR6Jo1TLfRtWQ8gcHNmjw1Ec1dELHfDV32xx
cFe/fGLFiTQFpWAAna4HaCUoz7B+EcjfTokeEAaqGNz2thGw/RWeV6ytfCi8ZsNV
1xxJmaCZe+/DmYBsZOO0xTBwBu+/kQ7ZslbKOzAsWCnbk36FDq1dKsYKlNo5Tyt9
Mk949o3yv0Svk42eP3VX3FCJ+tq0l0dUVCxTd99I6ufaO3zWFyk+hdkXmr+DKzys
RPK2lAIs1AYQBUAWzIMeXs7PuyX3kXNak0ZBh7ztErXl2xeVi98Sq/1zC+GtL4YO
t9srOQo3JPb8dVAOpuWmR5TaWhNL7lqgPodCZ1wByn3kaG17yRnBS7X9idEvIiVT
FSA4bGsULKBVkRcZ5Q3DMXKQH3UaL3U+vCyNYccrn30Ce/AimfBGHX0AUutJkm3D
SQzr+huNlCVQby4Xn5ir17AcKB2nCdTM5elUnfR3dGskT63FWmvAvzyB2vyIwYWP
taUln8Jslp9O1VIiZRpD8T/3KzhUQEVvZ64F25//RKqTV4UL4PCj848TdqYUpk/B
B3MjJ4sL6I5KeMQDILaQpZ3u9scwAnGSR+8xkkuMgpC6iaM9qBrCh5obFDBCxdMj
NkqiV4oYXVIiC7kPFgjJy2hOfXGyNCeHNYqlZkWIil5cB5C+iPejUalCHoLZEMDC
XhkVqp3MADknqcFZO165twxRvPjiqGPLoSxz0WlzoIKKXK4sBl+vd1inR2lteSWA
HhDdsyDrUPqtVoidfTR+zAB+MzhAPY8QXGDPxOaFP6AFiDBrv+j2WPeLvcQbDSBi
6PFeXETQHZ8U7D5UkdJhMrGEJ//iiKlL/QBNMNwKmS+5cyHh+rX1hQWG11lRTOKY
0Ys0WdtGwfmiPxO2eeQud0rK73Ee0vRsk7ysw1MimRvP8cOqHtJGzTxvnjcVVDtN
OtRft7CJzpWOvaXdbNjJOE7VTXYtGMUjFlXULJRHktBDQfzBT5R3/RTOz5pLOWH4
32Bswr6rVGGtOr0b/yJLju/NxRmvt22ymiLwl8xBIb6EPHMMHQ7TR9ZuGH1IhWDa
+bb23lioUIRe6gh8O0HmsYUylvHaOZJ9kZuoA9VtaL1LhG0uiDhazrgqftS+6j1p
Hda0Mi8lqDHmnVs0eOHZT1nMr7gRNMXqwUCfmGbGJ6sNH9jqxSqFUxRjlyvT2DbC
lf4cOZB134lZfFivIxz1K21agZj9iyDjPyb+PQhrKE8/Y+RClL1G2aPcI80KCPlB
1olg1VbiLvaq2KN5O0CyY4j3EkOVts0+BDdypyDOfd23jYHDn/Oh8AcGQAr3sEJP
+QJ/INxLBp1qX4sU5l+MBxEdVorwWauR/nu1XlOo+QARrz+T0ECht51AueQjIKaC
4v1xkbfG+vWOqVD0pgOUE9/smvb5OPYKsWnQZrHl2AURn5XHOlSOxDRZOy2fF54j
HdScctBd8rDQd/oNqnjDFw9ZT1P42N0aAE4iK82oSMxZ3qcmK03ZbWDblOE5TNm7
A1OeZb3lnqez0W6shHkR0sm0w9JkHrll66wTqvgOJuHIqP6ES78dsUfzKlkx92JH
gLGxgavoBugZfbi+XN9PX+rEpax6iQJKo4BZGNgwS2ms9MeDjHMCjLeI/vXV42sf
jkPNE6I/RczNQkgdgYvt1u9xz4hE4rdX4Dd4gcwxehukihjX5kPeIrcg+sO9UaAr
z/abt2Chcfy9PeYJ2gbsADh4atAZGiJ/o85Uy747vEhAkfPV+LyTTQI95BlFGj6N
6J1uLCmy7lge6X+iMErpWBDJDDWcx8Gxb21WmQZvsHI1ypbt/ygtvWpPtHSWD6U0
0XruZeOFG9wMCCn8oFCqVS/jnGfKe741BAR9MAXVP2kaOJ+FKeI9ro5kJVGF6ihV
4FBjFbXGybEld0HgD1HA25QC0CsEPm6jZm3wCRuBAD9BckJoCaIQyqtL2vLpqFAg
7QjLhYyUmGAFFHK9oXt+sAaQ5PdCre7k5T1pken45ceLu7nD1Ux1RAa7ErkTqanB
25SPDpK613INQ8gmFeZEhJ4mfXQSY76LywbvKcuH3tERtckIwIUG8R3ns4ShfG02
cJvyGQnNpOuniBoiz3mJOKF4WV4ctplZq5yqLYo4y+3K27R8jUdDTQ1Fc39sR0CP
HLzbdaq18+9GnQ+HC7ndSSgCoi/GHFSonmjFaGZR7jRw0BNbfbp/QKIMK94GXd7G
MzFrhGkTKkmXo080RCU8bKgRc2CLTv5R6cyqqYe9AwK3YN3GViSZZPdvphoPcyE5
hil/R0yTmINFvEJll4VcJ2JBD5vGuQd93BhZ82Qye6WevP8IbfDHxYw+FslQCVNc
iyX7m5zRdgjEJCneNaHFMo3UDAlocS7R2xZMOwez04W44tmLtf1yQl+9Yc/PO1dh
EAJk3t9ONbXgcGBgE5D7f1/l28OH8TMO4LgnrYXMLzUIX5gCiBd6AgQzyTPGt7XT
vNyFrVYaGKA+Ua/HBRXZUi+2PQ3yiZd1ristOKioRIuvPIOKhXsXf1zRIBMbwcit
3h/Kyf47P9AB1kUBbzs1eUkbd6bS0ZgM80er54WBPEYLPEv34eSJ4Efy+z5aLlx+
W63uxG5XOqqRIpYFZxtS9hZcIztLiPrvuz9BQPIuwka5iTxt78DZ43uhPFgca+3o
5yc19tB8IAJwdwDo1xuRZda0PaI6d1Wlddo2Dqv/Y4fhVdSTUji6z0yL7Sm30aZa
SDgRvL7+Nf+5VN3yTBOG62ubgr7ReP7Rs7PBOaIz7ab0vByxv6qMuZPkBJgRL+Z7
kXWugGJmZV2P23B0jKFoC86tHxfbfhhpYpYPKyQp7rc4N0m+oohB2Aunh65lN5oG
AWExHeW7G454KfBm/eecnFaRxtkaWQcTluPVaFovj3op+LyN6TD0E9XL8H5WPqth
DWvhXwy/+6i47HkqwruhjmIc7N/OMyZ7EM2wIcPk+qniXnSAxYpBMkyant8EveW/
/Mz+MnuR4xZSOWvuglCNH03nhrjXVLMeQ2byCw9KVzJr1zejnUIrUXAzLs/aWi7f
yVIOuGEohK1khCZhuHFOR6kb3VVGoIXTC9mtzMyrKYGe5s2Pdf4Y2H0DMeKbvX9o
ZxDrLrlsn9Hrp/UAKJw9nFgE9BV5pCUBggwfkXxyF5CIZS4RsyUohAXCFPJyniGi
qasTKfqwzJK5qWXcvXAtQUGSt6okd65pT+Jf5HakSlwH1rGYZyJ25b9NfdV6Fq1y
t/cVzU4TLUsEAn4BJ6lics0TKO2dEH6sqizFFkWrsUd/DC5ewq0Xg9gsUJ4nS+He
9tDP0ZnyiaghUOm0s7ClL0wKb75NPVDLWzRwUaZgWBVVNAZNUlP1QABpKfAPP5Bz
ZxBWzQkYz8/kRfni7zTd1lt8/rc5QP7Zka+nq55RGJc1XXopKCMT8NBkdjRJd5pE
Q3q478l8lkwvq4EO93052Cb//MmvM94K+K6YD3R3txdWUb7nL96LMJsDmSFNI5NI
R3SF8QvSOAUqwFzeC/A0of1DiEYLceKfQdJ0zJj2VJdu+93afqUt1hAwy0jXn2ML
3k8HVL4sFvWhXb+ZaoTergG1O4mvnvQ7e9iM8TkH4+5wXaXOBYa8oTxDlcuw2bsI
1VjaRIZg3IJukOR8pxIPUCCiBYcGbbchSvUBVCyYEVYzMEKndCX2mnA2ND79prLw
TVAfkVoUjyVOjc5tABuVcSoUsOes7sIW10X6DApd5eIrnez0eekuVgxdFemPSma+
HvqeLCERZmkE+nrDtPayeirYRQmjwglvnmBhk1/Q9prVk3K50+RJ/ATstc3OPVqy
tlgVZsxXDNNSNwqoOvyq/fGgJoKrCvTEBodIJJwX/5MyQL8iPUGuDiDxQ8USIAxj
PojlXG8o9IiUyCRbkMZ64P18qmxCu7pGWs1Q8HbvSHtvgBx2RfdRUHyTzuZPd1ge
8EZ7YlTO0cYCG8/Kig8j6N9up8/PrQNUl77vgl5sZ9h6+r1z9Hssixvh9lolPZ38
ev+d2d+5DEbenS9nAi+1jaOTJbY/RWenz6IhaUjeKyWixfNNwOEsyAsR5wwO49uA
kJarAdqXHM6ScbgqDb7dD1mdJE76wiuOsdIqNKXoVlBC6bbjpKubDb6u3+8ldYhn
IyXj/fjod2tqJzaFbe9IF5LxZL6tkHPBwC2m4fdgUHuvhqSQc2+oL7OP48QZLbTY
vx4sVCAAfTHE6wO41MljvnZqiU9R8GmaaokVYU15gA+AyrtdX7Z+JmkpSZ/FIR5y
lFWgm2aSkgdIU0mSYCiTKLBARefET369bEz5ca0hGmwBaMhttgL/35TPCnq1Aucn
8vFBY4m555Gw73VhN6igGz0Q5kIJ2HGE4UGLvMxCUudymYZm5PB7XoZQOlQmjHk/
ShyOskv6ddM6rm8rYLnKMwXZlBH7TzvXkirPXgD+w7+vEIl8hphPqNTRxmBRlEjo
SpsDiK4T9L+ZBizC7IprS+AUUX8OVRPV5+KMx1iQ2XAyG/HlJSXN56BsVQXsK+jL
pVNZnWhLFIfHbUeMJSR1HDz3VDetRL3pyR70exgHVE3DepeGrc+szvSJNgRJa6OH
Kq/mXkg1xFN/aZdwW68MTzGYlutDS3/eXWPE8depypXqAYrr+zqEHTiuMPBmj7Rm
dj0RILwBciuoTYN4gafG2tJ9l+8PaEH2dJtPFLvo5z3OY9JUM8AYbtxO9ZBd+6F6
FIG7GORXEcXWqiFqsTDE6rs7oJ5VnZnKwkXr8bv9Vdjj9iHKv2iNRf0fvX1uznWF
o6Py/tcow832MK4X9Iyj+i50WiWYWbN5ausICJXiyRa+shAgGtk8khY9H5KCDYu2
bXZNx9MqB/9levB9mdr1IDR5j6KAHzniXQSJ1lsMuW6UHHrpZTrjapNoIo+fY+XS
GjiIdPDhBoDI4hTIcvQOUFjEiXfXkRHr3X85FkBopsBT3EekfSzwIg59E2sXH/ZH
AVc1Oo2uoqUuS2MG9pZzzcSOnLtPUVzGQQfJSEIaDoLef+ZrbS0/Fupg3Ipbmt+x
vg3mU27Jg7cbwCFsCkP9SmyZ5S3POP2Lwp7rw9WQeI7r/jo3sOFCvuprNn43Z85z
OAjjy8riXoTQubE3O7p3HrSFhrdzvHKpssaa6gXQnZVpxh3Ak7pxb5CzHYNuB6gm
RCnZfDexL9p70GWEI3eK0xenR0tMbeFstoBSIUSS12p+fANgcBrVyKzbJ9UxmmIk
3d9Pkcz7V2LbET6RzhlZ77/+1GSP/eKFgMyk7z5x6JYwEHAvmhx9elMI8z7JIAIT
mhWNYupLqzLj0/Jhtsmlj3anwHQf3OVMGyhkwg7B4qLdROUoST3ZW6Ru/wpKkUwv
0jih6L9AMSk/G4OCllrz8BkGhuxq21WzyzAPREQ/3aH64/tW5R/FOJhxQzH7h551
tcrhiyTekBdcb9lOCytOd8kJHyGasjtIXDbQRAuSfr2yCcEhY2i6X1VyNV42FRcP
sgHCdNZxuDTMZH46Y39NFKx1psQ02hO7gG6+n3+3dOxZnCQqwFRzDJX5+i83Fef3
gsMhYDLjKyIJkCmtmnex5crcvHOx/Lwf9oqkPR1YHv+v8tIvN6cF4ojPAlogMXVl
p9d8/UP2bt7axYwEqtvkp+syY1Ef28vfUyJjK33tGvbwPlHA/kqXic2eNIj4KhnN
aEIxFgql4dchGGFnRRxx26w/OWl/UhaqN/Ab0qBGmgBL+7ajEjDe+5TuXGWtAbhO
6Gh3HY0WduBjpQWDhoaIYJEXH/mtmV2fYFhure8ES/xu84EymP00Gb3fw8rc8t/i
2LGr10Kiq/aQB59xydP0DRwxD8c6/buAOA4YlfOogJEt+KpsKjzyhynx9tlJVAzt
nEkPtzqkSLt9NNb2NrFlLl962ghBv94kbSMsbJXRhhhIgwA+XgFkyGZLZXx1J9B0
o7lfrj2gVh3pLeCqmvdw164TJ/3HgTwC2P8wE/ov2DlgiJIEMocdIX8OBczaFS03
4MOQYISKyr5fWAfkqoTbQmd2A6umrQNIFIJYW4GjcYgPuEXXpebZjJZ+7dUWW+Lt
RhCvVBQL8oX9VPGVSk+wsEMbqfRJg8Fdzf+KthBvu1HrmTnAnxedkQVMQqBR82Pn
JqcdC8D/HmOaDHLHnCfgtng1UcExLIXtluC0w5TTl9/frwvJwDcOcQaRsjFUmq3c
j2nYqJp1tI9gTSBzV0u36/IfCuJIIi6hbSrZVXykkeyAh5Lwq1GO8ClDqRaiONLZ
TVo1doo1R/uEREmt4DoKKvIsEzi513TOUhrozILyi5CF33pqFR4j896pldwiW8N0
KERD5tzcPPqyvYSCiii+XLVyLXHGnqsFEBGJAJRc9VphbldC8BrhCX8cvRcDfS6r
8hKiAwq1RXwXj8nhZcOi1wBRTVm/MccLwolX6ZiYds85+RUB1n64RNu9/7Kwsos8
34Tz05TE/av7r3UFU6pHo9jGm1vth64WYTZX76ArOWPI1xBMBJk1xg8JUdIgEDOw
Mzcbwi1pM+VrJEh1aC2QFXmNbP5QnPlJbGrmULVq2Udy5xo/NI+vxttkkKRSSMkm
HRPj9CeWU+PNPOj9Flj8vwzYzFoR+wGtlQEB3PEb+wamTi7gJEWVekk8iZjUJ7r5
7PpwSDa8gQz6/QcyFBU+ALozRQ0TFhzMtrPS42eCsEo37CCOlL7rykgbknaI09pd
IZZBdGZiju1wGBn5a6j6qAWu57qSlU5w0Qkli7kYR477Ea42LIQOUkc80MEqmmaH
lLQXnQ7E2gRqM1TpSV2pHviYvSA0gt3FiEmH411HtJfxw2hT+mjNkJNIB0RkOf6O
w4TeWzAbe0u7ta41wNakkR6fzHfIZv1uSViehOzHKCESqDP1ot01R6eoONiKn5zm
p2cdXbfIiSd0AiB7n0laqU08xwO4SDrznUhaOeKy3puz4TqNfOhETWxKeJ2Xr3ZM
7uU4d6y03Kd1I+tCtRa4GoEnTKb3VYFJXs1g373QmQv+Xf5Ls49+gFpDKUHKHIWb
+lIKzyWLVM0IQXqBVGT52VX5yBZ59RoWSaBeyt2uyGu6hrc24isrut2F+kK2Xoii
WIMrp/2p1hoLuSJn/uJ8YyIhsJ+G4Z16xtGcJ6BxWDocHov3qE5n8sVzWD23QUbV
YAKrkFUvBToisw4ZgILPXHM6ZnsAOntABnpHKYuLzws/ErfJKww4lmsqZxAnOfWQ
UcNygLgeVdW8tJB41gzHagFhuVGH0eGQex/k+60604mveVGIlfJyH2nSMssotcYZ
S+apFduBhmAgYk8VyawNByMcfJyPP9Q6qnDDyJ7+flJ6wt8sQXPE9Ht7EoUdSsNC
i7snC3J6hT5JDwYbRI5zkEFsS7TkBX7U+JpWhCLRpc6yZ8dVu4ZCb4fs+Ec06VWA
MhAuHdNRVLy1gWUdbkdBceTImvkFvpEARCAkYUT6dSrqxyyhwMcmac7KhFDTSyIA
xLRttvNUB9BmHVAHlzpxpfE2C2Cnr6ZAkYlBda/gSuMgdBPxr9v+LzsxpyHwJCjk
zOk1uQQKwlBKvpp81nSFr6X7MPq1ifvAMut3imz4YhsyIenR/iMSb68Ro/HnyIBa
1UoIEoCJLKPJIep8Dkra97ZuCHXtHHtd3qvN79dS7Q6oAh1Bjv/KJopeLfTkvNya
XYsteibtzZdPsm+c7HkFO9ViFaIAt2jTVp37L9W/9rYbTIGA9FmB18E5k2KSUfQZ
e9aXs1+5e0/UGUsRWk1hKHceMxm8ohChj25A2luRn+Vyk8J5h4LnZd9AfvlYfnJD
aWjeRNOAsiTPUN0TLyBtDM0S3C1S692Px0WGXB2uwFvYRlhcwIQEG5eG4irz/a3Z
KN3Ql82A/WSttvLEDvDvEDltthYTDr3VEFR3IVqzoJ562VVGKm8B58ATkWcPgeP9
Zs7P+1IY+YX24Hjq4eMVYviO9qWvQzo29Izm/ewuOzTqRQjnYgZ7BZhXowrJrfKC
l20Vfbc0aIWe+OeykBPhTlhiUpvkkVPNCP6zLZtUTJK+KwiaiDa4ApjPk3pEcR64
/YzWZNMR/p/SQ443pTsZPEFb9VDbUd4jvZGy56U84YZ/Igm08KCElHQ6o+B1pElu
UOLmewdT/1lzKfmPTPsGYKvk0z6LAQZJ8+TbFCGrZwe3AG5QhRLwEhw3zoe3GG5g
hF4ME5NOXKy7v51zSjYs8u2uA3elzwGhr2MnoXQaigMOkk1DJRHCvx4S2O+S7/3Q
awhbT+pi7LtRmbfiA9YrtaXSTOj4ISoSmARJd8z8Dd72XKIhbFjHyuIM0H8p2kuc
TpK6yZ3Rlx7rJ0y98RaDY863ICB9z/WoylMX28wybN8XwZ9/f2UlzuQqSNwN9v3o
TrlBqnaEekS29jrPbqY0Qi+2oDmYd+bwOzBsPHbo6FMzDQCrFxbVvRZ8sDtrNUNn
eD40ASNxdqhuc5+c6oX7Y+GrSyf8DqaJ93hVWyxZAgd7jambuVD7dUq6wluVfcfw
CnirkinDPKuZ1UbeVcs/JptN41RpsajkXfZXlh3/2NumoMl7Z7jkeVZzFS+lCCA2
pGnEngOaEICJ8+dvDVX9YiRxZQQP2yaiKqVmKSnXWqOPvdXR4hWAfhm8ScZ6AyVP
Zq9o1Fnfk6Yk19M+ONDaXf65Fa4gY5LQPlGc9gwv5WOjoZllP2FmZGJK81wm3FhL
MWzb+CCSTDKg87MoL55D+E0xgRq6CdFSjLfQxn4my/Wm8ecmjOeEs1lehfZXvsej
27uOrbqJc0W+/opIrfQoaRqtTmB0QMs3tYVZrWaa7uiynx67c4UPckYm0xdjzLjo
UPTYFlnGJXZfnP+4Ro1HDiXvp7eiZysT9fQRLiIDmiUEJ2K3zpDa3jiM80j0PA5M
qNqO2RFYndZezuUC5gJCP9IgtXoa4GtVB7MlhjNYD+lo+Q7W02b/GKOdfuuFk04T
hEXp1WXnyThywk1PQ2dr1mBVusNzaiPD9kUS53QNjoBHu55/Gqslc/SNA8ChXr54
iX3HCYePpt/tvDd5FZMmIqG4lzJN6z27yqLzoc/lzEclx3uG+QfF3HzKSU7N8p8x
vU/hMJpPdH/xfMK3ZsJm+15A+qb0AA71XbsTBTBJdgdbCzI8E8J9sB3OGLULReKD
9u/cepF/2i6vsBVuq9rTA09/j9FNHO4zIgeJIK1KDxNYNDqKJF4uI6f6ImPwqiu9
LITcB7xjXwVKYvd2N2vrR7MJS1hqMth98B87f6PFc5ZavIAMtM04NshgerSkeAn2
FTGeVPWooycoXeVYfq4clbUh1ifN/WGDEPSdRFAr80CTPYbQxYV/NyE3pbEBTXN4
qnGPx+q8xwOPEwOWO6cXqhc9/Q9VENn/J20Gz+JySxKtzHomk3QYk44epeCfUy6p
WP5EC4k1bQA6qrOWRUS/xJuyv+wpb5GYXZrdI8X/3H9K2RzONrC3Wlay63phowG7
xCe9bXK7ltmUG4YfCTqEBjZ8rNk2Nda34yuI49XELuVYIPMtqAfk7huMUPn45cA8
Oijx0j35V2tAj5EleAheaQkIiSjz8W576AhQBIraARirl+oUV4Q6oGQP+XIoKDrN
QeHthkR5LC/Nyws/ewt5Zg2kZ3zqysXCsrzPRt3Uvt+MpwQqL/ivcuTWKIerb/rV
DdBUh1DURdNh/7uVxYNR0qbF5d/yBg8liWL8wGWCB91w0DIvonGe2yt5s1zAtFe4
qGSPJiiYH5tv7Mt8LxCojIpjoYgT75LKWuelIfyXnh1ngeMcL86hSEInOaSuGI9q
PC9dchqB9Z3BmEjQyVlQLVInCDiD4EEePI9BWNbpe/jTkZIa6LVxf2CzhNLn23l7
STmuVuVN0ncs8NiLm6WnqDQRXCwlDqDZLO538uibMBZ3I+ma4gIto5Xi8FuqX9zt
pECXHGFVxq06OUhs2Aoj6iqGI5IRyhCSj2o0fT6YNv0OF0qWQkRH2ok4fibb8sHD
5zFwgUQ/hbyttIB3/vFpYDUkFaZoKWVtjBgnLsEXcHuQ14nfwZlQrJEqNvmBg4My
ZjMb+dSUaYRxLhoxcfVFq9JzXv1/KqL9d6DKwKK3uSuaQQYsasKha67/Ounu6nEj
XBc7VcImM2xQRGfDCdBGC6ZmouQwP+qRzsQULF+0Osg3Z/PigtY4yzgE+Dzt+sVo
5mg2Iv3FDAT+i78cjJQ6atI1dU1UatNJZQ7YBdsV82vqA2hK4eH/uGV6VQeGBnti
GbGZqfmmU9Scaeu+O65O0M0xlAY3HgqbrcQDAlYpCxjByKpF8yWoDbChUpPPuub6
clFWk1k5Zx/Rqzqp4A/JlqOjIaacQWUXQkhamhIvzZDxwPn1rVs7Cypcmel4XUJm
u3OZLQ2vZrLPHxu/+lLav8fibtaQeuGI04WK/+JXb3Csq5R5SXJL9bKjxSSklUcZ
hNimJAhdrH8eZHIuWBpWVl2TSYhCHcivXe+Yy/G/EsXikKsRK3EgTWxUdRAqOshG
psmBRvmRsEKg9DQ9+c/FaxTpah47MrxR5Dmg0ysBSH+9D5uZoUvGvuSxmm2AaPVE
SCwS8jpmiu/MhUMEpEOe0PQKkw1NdEWM0Dc1d29GZ3y15eVeXyNgATbCa91Y3DWB
FZ95ALU32lAWLa3yow1gDEWMKtcDkdA7gK5VdiLx06A+rYFL96kxQWiOM9plnUgI
YvH9ibpzFcjxex26QMfCNyocobcAgP4OJR/mE700olxlpL9qgeylNDyVQye1fSu+
N1x8EgZAa5CfNYg7zyx/54Kp6M+mPglBqn7JOnhQwLzMm/cMJZTnarlCDMfBdZ8J
vDXasJTCqd04KlO8qC+bjokY391QL1X8A6bu6Jzqo9zkutmWzCYkQSuhSyL7s7Gu
3XUPNaKAO7NYS+T3YfHr++kvYFuN3fID+eqKCWSbosgW04/UU2W3m43u4nndumtd
9mvXMsC9RIhKHdh+sPlbt6BoqtII49u5XFXm0jXrD7J98ub+KepC2981ATTmXejm
DHJhNEeccSyVjx9mC+LdzOYe7m+h1fUjaXM5I/FSNLtClFUjVLNTImv8+PfQNfNr
DwZ9eiFeb1i9Xl2wFzLaC0054CUrjrJ9CVGLX8Hx7YjPEbWZ+Gk27RBCvkn+kK7Y
SGhu5FfyhRP6EeJFOJkg0MjvAsx4VgCoXkqJc8kuebBDtb7gkpJpZbD5jsZLbR6z
MWW5XE7WCcrAxfzNTt6XqXbw1ZJpMDywyFWyvPLYHhTA7CD0LD/IC/pNcbKU2ey4
YxhlcFr8KtCozg9VcTJRchY4dBQ2zR8mpJign3zSH1jqneGjpX5sFgCH/YcU3gPv
FtwlQs7lGdgSwNMsau89BN/YKMy5UvaP36MW1LsBkezOKKFGw7KGQ3vsSb3r0A94
3AKpeE5ZE8gkAnsCcdfpLuOdZFmlzpVh1BnBIHfOFK3tJQj6vbnCbXX9V34sKgp0
obrCFeI6zV6hqa2fWqSnP7uy94ewMGVXa+E0NGmTRWOq2ODt1CGNwUg9+HOJ2/1C
l+E2dKiT4mK/Yp6LSyIUqmwLlbGaKxDZ5fwx9ih3BrGML+2D0MljI8n7WOqfuYAZ
odAPA9GhIU4b1JXtxSHMxq2elZrlRiQLStwUa/LV1GMNhBqcDMPj35CkFmh4mjro
kJj5QMAzf0KjZMUh5vPdm0Wag3apntoM/pLFujxT5fuZV+bNMciU9WAyg3R5pQuc
SeXMoNpQ9FEtdYy2PwODqgmuVjuhDzbHyaefTAG2ma2lTq1nfMc/MIbSOxk7mSiT
KqMrSQ2MWP0muHOVSxriurudHqlpCzbdjlUGItGHLA1tOv/dMnwqRWcJ5QO/dvf0
PeGSsQmdIEU9lFdyqEgZrTUfwcp5pFA0MsAOnThuj4LKjdezt7Vp3ofL8tS3ppMA
79AkS9Nfv8q7S1ABfuCIgopy1635/uhJQSzg0KCqSnFJt/wzWMd7S0OFtQMdgFFe
5ELp51bulRqf6nD5+nvgN5I/NHoYhfrNRNdiL+g8aBC5W5fF4Qy6y6yxTe7e9y9Z
g7DsncQ9olX/91lHgHvWo7Doiy6QfnV4kKMrNH4MadEk8HIoONrnqvKHeQ1GYYiP
49YgPXTC4C2yHwTNMNc0F/nkYSVx+dJU7KE/avMzaZ5Jpll9+/xtKDs8S+8/hq19
jmPJy3k+VbePLtO84sP0xxVnbE2cjOiI2b9x902XcTlxL5iJ09dYcXIUxDtPCbOM
epiFkB1cWE1AaN8A+qWhKaOq+9EvqJWrxVdInRBZhMeVpThZg5s8M4fbSO/+dR7C
FwCfUxtaBJcQZYH4OV1SHV34/Cwkv2EbAGYrCqhdHqVN95WcTw9BrDu9cwp4xA+w
BJPF4nUztggiWAYTVBStjm9REOysc9788ZEExkXLsmSdWcTB7a1xvl6yVBVlXaf/
a+6HFeYdAv4vhUZHAB4zOK/ss4BWjAFIw/AVEp+cpawuhcz0vUzzZ5X6B1+nl1vh
wUJKKCUOf2UVQ1oDMB1oBcZRhMt7aX78qzFtnqlaJ22tT/nqIsqgTVkcjaOb0XWK
qJFpMtjFLTIBXN4MnGimgmHU3MIS5ftpbjoDejpl+1VmrczUlebdRRSXaPKt+8pJ
M1pKeEltafhV1yTT+zaFr9gxdr5b6zNrx7RVLbilnFr/lBTP8c7muOjvgnTE0HPg
5lhECyNP8qzlEgFDOUTbKUmPsocUTKAOadpBAe0M7A2DaijpXYTDVFBMAOe5lk2e
Te24HLqX8UIS733xogR2ToYsprJrJE9bOdNO9smd4094FbRWbssEO/abnJy20KkB
9PiYzYAyvQ6vyc2fw59X4rEb9Ra3prZv62Di9MxyqLOb+vJiVm4eCw622sbyI4OO
8BnHWY393mRffWyZuUyR2oWWPo5aXNvT728986/nJNRg7FuO3zS74GkYuYNUqfIG
6+Erlz8ZyjLwif2Vy4MVBon4WPq/7QWxkvT8L2s/e8V6L/IeDVJx6ojcNgRyzyab
Fi0AEuRu4DN2NCkwRfWOqoLCJzotxT8N4DLiROL48NNYuU1q2jq8RPNp/bbcQlpz
sU6D5LeFzr81QTcGuo/XaqVZl/q4qOTTf9DKncZQD3QIk9qkk07/9ynCbC7AuroK
s8oVyGDHvklWcUGHXQU+PXGycLOjxxfc1Wj2YFbB2ACQyZPBepg6P1tZilX7rrrR
UO4n7eCvZELuZnaoSMXLGD62ELGar/3koJViLjQFugDRkzd8ELnpyCtHq9LA44VK
EtKpteZfE68D5gqkraxv1K80B0QLZKhU22VOyLJg0155/61aPs2QKF1DXWVPuVLO
n2Q1d60CXNFybb1qeI5W6nvY3BWlbIGC0SP1P/aUaLz/jkl/EGrxIdFyhU/6WtCH
1x31mJcqSitJoQlPbsxa8JngpjjYcoij7RBJP8TBFkSwOrhZpccsp28sVe8ZFFFh
TGZ/LPiO0s71ss+h3RKmQ+R0XfhkKyukeNcoAn9rqFjXYjJYpqarcShL05b4d6wZ
hRMZhHji1TSgpDISDjpaDNfnNsZxZPa7AwVQlZcjA9rl2MKP14oplPzTglKzbR+5
0Dr6j4ghJ7scbZLVT6jy7Nb7ibkMDtQ0cj5tB9To6X4QZFd06ijxf3fqLPFIzhfs
ObeXNASw8IWylPu9iLqB05QDXawT73DI7BYTxM2xapanDAd42r1dydXdOsz9aB+w
S4Ut6T3XnHgqkWv/QTnzpc9rJAmvC+ZUWXaO7IFo9vNJHobGjJtx43uyB5SgJdih
EkGtCf4CYgtsMMT+fkTGECeBMzDZ6TPmYVyHCvzMIqf1+5LcNRA8MnKJTnsyJX6b
xqGmX4ZOiItHNB54Lo5giaCD11/6YMO8Xk63a/0j74rlC66GnnkJZzcsB7IBiePk
rIyrUgHJnVHfk0ZhRP8VT6YUAWn1+99JLathicZldqbx4e4sq4EPOObhrs7ALUjQ
q/KOegPKDFVQ9RR+jrorGBsxJfDGBYxgydd+k2NC3fYpDwuxGGbLgo1KQEZER7d0
Q35yM5mQDh/DzX4mkvHGVUen9Dr1xfgGDYIbWC10i/nfLPAnABqyfGjnmdyBYhBS
8O+t4nFbC5fowpHMsQosJFh8zRbxoUxDAv1ZMsaqBEJrdOpCs5u9HPiGmXjnslnB
b/L20IQ5yOyG67Jdj6Kgn8p9APL14CpxB0vfpJ0ZkTsqkYM33f8wjDsV9Leyf9N6
45DOq/buojqhn/zAEOn1qE8l8gJrxT2c/AXSimarpOFSvfwPFNixWRa+sHR2Kd+S
8yjlbyONKrYeK9ieDj9KLWPxMl+/w3ZA+U8tdHoRH58qHXc9/8fis2t0A9JVUZzm
gyw2SVL7OCImtTSvqIUq/kgNFAhz8UEROn5Y7rCKq+p6hIDp6PakrdVol/mB9oRQ
aFwVynjYk0Pklq7ZMc+riRLKD4wTP557EHihJA/QtdPPmnf8l+a7ZRH09Eailv9k
7R10w16RLPXl48X4uNRmVCFal9dRLgsCFPH76JB58kSMBVHe1n5qaVXtv97dlKuQ
4xdaFnWnhmb5z+lrEBXl+7ZEhkhnS9LuXzVs4jW3RSVHs1Onpmw/926dr8HeIRGm
24y6WlVjvlhTPD2pC4FT++As23mNNxBv6qRJP98dRDCYKp+MKVfGLocrtW2uUWVC
wzCIQy4tDZA7CpxqTWXqRN0KUlA6pLTqAxgRdKwantq+xErpEiDwTIYBUzsHSSCo
BKh05F9kZ/Or8r8UV5ZHcggVHTMiGMTafB8fAyX87B31vhmYSewdzhNf+Ck2XmDC
jgSORoJSsO7q63hiWah/EHhn1iwJSG/vJK8XtOjWDjJJh5pNqXhFSE/G5n/yJMct
v3z5zN4DmKajbD3hP9Knu+CIjWnmyhOo6EXAhijghbWXBTWlTUzMmskSA/ZctkRW
eyKENhyN+MbBTfJ15CUTSk43GYoLnHOexivGXd9rCQR9p7FZvNU6RyBVDDJCvOAw
yJrtZsguBiw7J2rrkwWZfxgOsaQMvtYNN8eF+IZT2VSCj36lLc4q7yY1xrNW5OCe
U6quk5LT8mCApisBGz9vY2SbS7QVkFXdVjVmWXJqXZSwBLSRthFqhbnaIK5p+mjF
rT5jvzzqVrGGKHW0YVRvy7UGklx1T7Em9ZpMHfIIA1q9CznKpYwTeGU/cJ5Mp0lS
RB+MWyi1LM8JoUK/Fh3KzIpZ9hfv8gfiOwgM8/6JZRPLZGoyteNXgt5uLozl18WJ
VNO0cVME/y4asMxxs6LVB6lLor3Ee1BMLwUPPKTB/tgvjUI1jMj6oIzQdKIf7lqI
1J6UU3gMfFpFn07Gd9AVby82BySRz+F7KgBVeXWPHsbNdU/1QoXKhi0e/tMKzvwt
Zsrc38uNOAePMBpMmc5d3y3hGaRVHLvcTHj7DZP9/mX3yLBA2MGluFgYSsJZlHNT
Lkcy8wTUKB/kt207E8zczbMiEPZXIblsVvCm3mhHdyphWwWU6dBoMOjD1ECU77UH
7ez0KcaHZkk4gZF55jAHUDn8Ykjl9mlQTiL814+wUhF9/pOXGXyLedQtIHLIGbFu
/nt6x4XJPm7pyIl5LxFWw60QrNaS+286YRw7fxpQU+NWPnIrL4/GIkeAeOblFs6Z
aEFb4gfw19zCTgRVnQH/7S0nSWtkZdOZBNJ+brJZKVSMdDVfNo62qbEkWpPJ391k
gnQUifp6NGgtdrpeyMZYngBlNqV05ef09CVS/AqrqhWrnFalNtkg04FNmPbKNAIC
NE8Uf9Od2wa2rwnc3HqXXVF1c1J2ntsuLvbBzFE3F+c1rOacMuqbLtRXah9sepoN
UyLH7A7ZZq+m5B59rmVGNfK3uoEA96byfAUBWudY+75b+nSoTpa8oEUCpRPNKVYa
s5IbB+pNvMxuuAJZ6LxcOoHmJc1Egr0WftIoFnvhKEg5OnIOyFj1cDPkJCPfabVb
o3UXfPeGlWO8EWRPHLhPLFmt3XuKjoNW4d36HSaSnVEGS5Mex2V1IqWGrmQ//l2j
voarLQlrdQ39p2Him9qISd4iIvT00F81FxfQC5z7OwGTjVq9+tI+RknGYgSL1rI1
0xKXgdBNWn+EalvwXf2iHUBvdfsnWWoAzZIiTJoXdJEOvKPUqAibfLupxmRoS2/7
jTSEdMfuzSrxOXtX766bAkIfZ7ypVSxzRN1Ij1APe3FbfAwcZVWUPJfsPLwjebBM
pcykE1vraEBQQjnqMCFT0SsjhdX3eZZgkDNdzaOas/41pftxW0ZIIVXB3LDOcYjj
5kn+wiBGugCn3o4q9XkOoSEbB/PG+VmgeLi/tPK/akYx2L1Rp7YphXyfZDDspS0k
ZglWsZCOSFnrr+06QW64KXLwg5GLzXjR1uvA42UMEu/k96H/o/BJUKCfD5JgrM36
siUh6F+m3tRnAiP07l2XgMskh26h2B0JuBtOIhkjTqLMXOANI6PsWd1ZghycwEp/
BZAJoHL08p0Wrzv7ol18q/sMHHpP4T60yGXRPPkDQ8d+LKZ7EP6LQPjTZ4fpxlXu
Ew6by3TfVDlEAQcu3ti9EscZzGIIQNe7T990CRicEF1OqxM2pKi4G8FSm+LyI4MJ
QqckDi8YZdmqdHhLBcfu7W9gBb9EpL7kIGzoOmygOb9L1rpfkh4RU4LkAM+Y2oPP
SJQdj0i4rKX6HNMUyNxGj7viiSHDY2w5FpxgkpzNhsJEENkq63/Sfvd2VTI1kw3t
U4//0VZZtTCdjzUJXElTYe2qIzYU556wMw9+wNRtNPRKSqgDBnoS8z33M+Xqo+Z6
BovCXOv9W3ArNFu4hIqR5fYJdPUXejL1mOy9uPt7jJrr8K4cF8TmqSmo4Abpm3XD
jDmvRIOrKW1I5uzXCAAn+i2wlLzfTn/0x4J+GAKY3e4YzJ2YLm/8NCXRNo6Eu3SF
09GVhTbQ9AQL9uvBulUhVEPzrzCa7qbyYKGbIWkZFxAyERex3muqQIkMh7BAzjgX
Pv8NUyIwtg7dvA4GwLFWFU55ueHpZf5FYpR+7TJ7wh1/qILi72ohWNS/p4eV1ZI/
RKRnOc0zxhfJmi+5XGjDMFE8uG2hdx43kr+3jOw5lAmTU3SF8I5zEOb2UN7Qt0+G
M8hgH/bPcQLw75LWBQLcH7uO/T9fo3VtO34GyYHRZ5JYqZOo/X3jIdCuOmc8roVl
tX7VfSv0en9IZQGw2CjpmxQDuu/Ht3uZ0GvbaUfBr9nYg9h+hfIYdVD4xOIdBKWG
HmkF9xbnhYj3EC5T64ha3+oHBm8EULZSG7OkE1qPrOcoc6XqvVBrkRv2mD7riSka
5a8Y72r8761AHNEAYLx6tOx88GWd/W/AEMzdQP7/wYPYnNwdBFOx2X0FbI0pl6Sh
NerVTaZlJl1GortSKUJRRe3ApREqk+H0rt9UtjsGaYwBsW0mb1W5skVjMUTJYik+
KQtrOhah90NQmCVefl4Dwnpd4oDDNHuNJLH6HTylw0ChdpoluEmMwh9Uv8I70Mk0
QeT8k6lPOmEVS9pzTOo2DPzEvq5FtBxnKzW4EDV7EZh7fONaPtRQ50KSqZMhVy8r
oizKKYVYcGb1Y46Clyq62WPUaxEva2JMq7RPRx81rUy90KSEUD5iBHb20UPF+B85
fy3lTMszMejiyORz1rRlu/dovkNKcI1C3q3vDlIGhi9IQ+8RUYYd/mVLiIrmQRfy
akZWuG96nXv/xScUzKn/jEpB6ytuSAMeV1V7TwNBRKQoRUd9J0mwNiACfi3UHbyS
U4L5feB4gMtr/ZQ5/GOZzhZljHOIgHrU75gfg5uD2vHi+90/54LJ6lv39I7h1jxn
U/xyaIeGmUInq1ItrZsH4mVdxAYCMaNyP5TRJkO8Fy6C5jOUQpuY1+fz85ANnuuq
Q7+h6yjEZeEaZhEMWrm26/IqyQtd54taRy9fTnWVhSA5ga9KyYGErVSqmTnLpk+X
pCU7E5uSGwVQIRRd9Uudbvha+ODJ9V/XH/ivxEEf8j6AEbkPDy0j5P7UcYio48lK
qs/k3p8rjFyVD498ofWCpkJkmu61ECyJOIfiETaLIHb7izGf0FwoHqb2by6WPFhc
80B9MAObww/geZvAhrOlUlx5wtEl8LiFDHkIABdvqFsA/KoFUXrMJZ2qJbEsiG0P
oiYiDI+oFM3doaQamGbSBI7dsQs3bc7R0gha09uPRRwz40SlzM3jIvrXNrak+wzu
qJ+QYXT0yELrIThxHAHNjBEKMmUeBDTg2LgfbDxQWo/LWvUNtgRdZkC8mI9mJf+d
UzXPOAtzAGUN7iq/9GnYi9hd2vD01TKJbzmxfD+3shTkVPPAmhisC4FxgNkkbJJ7
qzDvPPuhUlpScvTXDu3TDIxnZsfNicuTHDHHCZzlEyPqQrRQtKXNNfIsaG2Des0z
eh70RGSlo/yzgPl8dw6oajgA4aqA2N86Risk71mjXiiUlFBbNzWM3dmNQo09r4zy
1fUk9v9HteOe86kKcvysD/Pfy4pvktl0VAUKBy0w2/nRN5n3QgEgdpK5KDEJiNNd
1XbjSdRsg9CMyqTHMmiWXSK4GyVevAd87HEbZPFUzNNJbEZ11Aspmqrx6qAoLDP+
oWU53kNiZKbmUN74lOVBWk53srcwglpHF5b7Q+NYOBP6jGitf1FbN1I1j0HdrSRc
xQOHUx9epGY0nVV0AsABuZOpwwiPyWwv95T+JHtuWSKLMzm7RJWXr5ZkvkrVytws
pIsjX34CqrRrkg/aR/G7HEQEZ5MBxrXDQlczW0i7NDlyWP9l5xiO87rHSS+M5TJ2
v7k5gPPB0rLD0zrlepQcL6FF4yMvUTovkc41E05UgYHqjfU3Vd1JnK8kYVJ/CUKc
OPTEeaJeBGbPLnWdxps2BZXUs2U3KkWWZ4bVHJMeF5uts2rX8KBZT9oCQPdm8AXj
J3ErgVIucudH/pJ+TDV7GQP9jWJjLRoe34Lr0ELtixMNl7PTLsuQK/R342j1QzCW
MZPjYNtutFLcuDEsnCJGEqFAGW6BtyWPG17x+tWoxUPcz5S5z1XwZyD0u9W4YVyl
xI49DJ6oBqWPiJ2/IcRT1U+hqRLrg0/iOeJn6OV7pSj3o6s/lPDiE9IbMmkDx/2G
mSqwVIaMNtpfhKjGSKUETzeLOkV3f54Hm/bTZHKLeiHOuDXoMpXAYzkaDE2WcWbL
yLK4Pp6NOLSJgdrBtvwDl0ZdFZiPf++InLNI9CBRa3LDw0KB02+beDsLzOlwJ7GC
JygnINWw/UJqfnwXvX6sdGfVoPcM0JN3lmTJ5s3n0pOFYRE2GXrptm/8X1t4byft
vPHYE+R5e+ExiN4ZHdlwoWpkFpXcS9K82ClZjz9peIPLtPTzf3OceqUn5hCMyTFZ
sn2kY2O8TO/tkQQy7aEvR8lnLS20qkhC4GdV/D0lBHePFADgioNos7TSs4XoNblp
I2HjSZ0SIYK1YWMZvnAeO50NQlrzP+DCeR+L2oEiumEwcUrVevvjsHtiSYZONq98
FQOVwDYtU1aJIT7GugHxUCmQOG2ewowB1taqPLVOZ+E0WWdLKNBbb5NJfS2OdBwp
AxGLje4tZEudui8Mg5QWAhWqqP9/bF5bv0fiOLg4buMisSXnBmxx57s7BvGnt0C9
mUP3I6jDZCvpuydY4k0Q3Po88/KIFvbEVKQE8XLcsUX9L7OOO4eSGf0MZexl2k4Y
lAjreeF1w/crqCyTJKVVu9yG0+JcPM5k6R9KiViYZ6C28D3Wk0GAIFCMzBnzjTFa
aPz/OteFdj5JdohXXqt0ULDIYPni8VUDDhCc/w0G5lpnx3gG1s1JX3/12+bq/hQU
wdJiwDAWrHJbTNP28J9UJIjt0s3ttCWZ9R1tpkuLbAwM4K+UYYzl32pXnnezUXvt
tvDNLdYixwcdTy7RUj5Wz4BHtqlN18/5GHyasNzhVJVRhbWFe4Ri1TY5uHNS7C3i
jlYe9QA48BZQdzWeh44Ok+0/TAYU48pEV/oyJG2QOAcUr+VZeC9/wPF5DFxuWMhM
UcyBa6Zno7Kec2VyZvFeeDLkh59CnAnZ6FptSU2dYcQBHweEmcznyK+ASoXbYd9Z
fp2wCqSiNBR2M1AVwCn55wWpRYYCIzVZpxzREi6ti/jM1+2aq6LVhroq89JOq62W
PpkuIV6fdpCdYuJvH3vZDjBH+vqBgQF1ZwM13GoaPFo5UzSmlCIlh3Kzg7b5e71e
5aDrBKpMg1SP4I+gvwqYUGJ083BBLa5s1j6Ip7Y4QahOBKzmOam9ZG9yIVCKbEmZ
RJqYJLIkbn/J8Bxg4Nu2Ir0l6Q2IGk+hip9if1ZpcairEs6tz1gCib2M0SbethG0
z6uGD0T/d+hzQaypVnkntS4u9xzSZBRy9AtZl+ZNDITM5xVFa1ZjU+I2E71vVFW1
6rssoSJMmHsxCrqHKLLZ4gh1m2P80kN2iszywhMWm9n1N1zk31m0aY2yyfmeG3h8
wwVdG1h4Da4kxTWtzZm/M4pzE1nPqaB5TFsaHNw59WsVgw2vl6ITEaH7Z8jqT5xI
BDzeZ5tFKZZN1SRTTOsks42NtZUMrB52JODkFxsTFoxxwvLxDlW6ST2AmsjGvQa8
Jjo/QgWb8zrPflfoaoqtqHbr2GVI70WJ3b1VGmFP3wPbdGQTOVqe2N4ELbXE4igM
nmKLm1Qj6GqxgRANrG4SAvuhK40vJ7jfbHl2Njy6v3c3vDQE61knAILOAhevAr1q
kcLV3veCO5cRzQYYw0rdiPL3BfKJCnnL8HPOtIrlUwNkmXJC/c51QQC3SzWc4MIg
Eq2mjGN0nWYierz6vr3OH0zBZMViUoyq6BIygPQINbBkAbeja5yzh9X3Jm30LYFy
mvYLTWVe2ShpK+zgl9eRbCfejyRu8PLezU5x61Fuxr2d786u0kOlGkyn5K5UexGn
MuFMSn/7Sjr2sm2pCnsYReYtJ3dRIwGGh7b4nnWfzGRX8Lht4wpbA9kWhIdXN5My
4wJGU4GedpSVbmXyEDUKZj0UYMo6ZuMXGdxxHXo7dSlNNc1SfaiYyMfRgclXVV5B
7qD8DRPlKHM5TDFXeq0CUN7id1M6/R5YMoj9CmsnCAP84rkF/XQZXcnsGyQJTVXU
g7e5jnyIUDfMQyr4cMmHZd4MUs79XEbMY5YRL5hx5R4OBbrToIXCjB7ezfEq014A
NZ/V6CP/lMb+8X/AFFziJf3JClGMC8X2QknY0/4rhbPjykLUaippIm5wWvKMVf/0
iIHLrE+bcDeaZw7SL3SJ1490AnfF7qWRNM6r2c5ZP7posh1h0LPnka2MEnf933ou
c9qJIfmwGOrperQSpqi+t+a8p2e07W6mAKl1bwKvlUxakfwXSzE8TfvaQXQYubvI
9QwTQKD863BbFW2z2rmDQN9Vdz4PCTXBoqQ2Ws3VfgibzjpPcJ7mG3aGQ0YuoNyD
m3IcRSLw82q3wPxx+5lCpDSZ4kA1kzVXiakf0EfsaKwlOUUXI/VS/RnFQ3C8TJax
7nX/2EKhgpbEO0FNqCTQC0JM9DKs7Td3fOYHMBnGDRPiiMUkrwkSoiwRyMUswQru
b0824sKlGWYTytVXJxVy6mXw4mrb/EGnOnyjHN4aGTjj82JtHxyjYuta+/puM8A7
AvTpCaosN0P8XpKMW0tITr9XC5LrhnQ2G/ci/j3DFhGnZeY5IullLCq1lH+n3cnh
JyIR7AGt36ncbqx8PhNgmFOTmDMnRy1Sp6riO/kmFqrxK6JOSGZWtst/d+r79+Mx
j67BjksI2jc48KX8l3ymEGl+1SYgoKiFol/sbbA4RjnHE3EYvuyKMvDop7Wh554U
JI6C1QIgmrP5PAYFwIwTn3DY11bdWuwzA+BPJ8qD0rAjJHCSM6qKgQG6AXEVTqqa
iwumfl55O0WwjfIwmt2uw90A+f7BhfBUyM0lN3/B2t/rQKV5Xg1N19WjkMNtu1JA
rlKWutJZ3j2drl6lB8GPKfm0u4RQ//7nspTZXPdTJRDjD0wwNrxk0x2Ur950XXor
4eKzxtUo24XJae0/gKVClLjoGTN4mXq8zL6Te9Rsmy0GuC5Ve4KrHsSZEb6EyMxg
ps/cSGuxLHTJuCkgj/fSXOzjweuo/gvI10lICymB6RsdbujoXw2VgafVHdTZwnCC
auaS44jZF5ZnlpVmWK6gP51txtk+YyuSedd1/NJ+uuRZl2w6HWjW48XU5WmLSU4w
pU2ByjaFkpjVVYtZoI41tvu1j4BZNaK4NLSFrWxcb/5XRQgIHVGkF2YvDhCfQLaP
JyC+f7cPB9r6rfBpg3ZW5qTMF8PfLiJDfoBmNXgoahljd1nGMkGCZlzNrG42IaZa
baEMTQ+s35rdsQa6oriUKjx2KsFnKwMdKOk01+Ed2NFLDHdrxbrSuvYnRyQ4mP74
nYz5LrucyhMS8qOvGPwGnmEXY1oOE4mhHPysh77HjT3VKk9qHQCzoV5ZWHZtCWdx
mbiX0/Kc71DvYAkennpY+7Xto/9q+Y9KFtMozCdj3nDllJ+fzi/VLMsd2uwmlaEC
sDZFaRV8aWqiJIFYbvlZ/7xtW0QZzdEhgrM0fBiesbFqeTo+aBJJCHvWcwAUzA23
gqn3AyHY/p0Z33rAfTqLUCq9qrM5YADc0/kYJJipQqvrFxvjgbRkVyTydnIwmOdx
eQYp1SxYY3Iftg1lYu572zRvZutPxtNzDnIFdAxkCPNHFSSCusmFe6jssNslYzUX
tbWkXE+M4CYoAAkLNFpMXFrbThNDYFQcx2/LX1HrYwlLST1gUqKEmE3Hsen7IhGf
yZLyzWv9gE6AaSVW7fpNvfo+BWTWXT7xuPiDmyUXGI+aKhJGR3s1/WLfh1VvtBIf
oSeoRHq3XgVqfwn68tMAbK1UC5fs4PgTGpI9DegNOINRbXHhlpa/Z6z6V2g76iVG
Cvk5Pk5Wcq8SMJ6ZYgNqWVzZRZ9kI4GaCY2e8Le519tcBVp5soSzK0Vp82OzjlXR
mE+3nIdmy304DsVyS2wsO2LdAh55cOemcsuGjKvbUXNE/PkY1aHyLzRC0HfN0eOa
FOtuG/cqr9l5m8Wsiogm9BBCdS06lQ4cml4dzCp421bB/S6etdWUkVgoek4xISiS
gc6Mjd82l8cRuA8R+/lgwk0KN/6riQDqooJ3UEnOeXrDbfNrdqVNF7CkOtpMWUxs
B7AbYA/9BRfjhetZaIBUTDX/0YFuSE7BDhRC/urWBL4qNLp7ba191nZB4TuqU88w
d/jFtg/1iLXCvKAoyOjvdHy3nfEfDaYVxjPommOTxVTVpMlp8FwT2U5PTfhatw5Z
ejjPcpBWq5eq4Y60xwfqGnI8WpnbL8tuLMW3Auw/lrw5CrckQiC4doDfAjuy3+Vw
sToF8kNOoG+vQnWsJIhzl3MhLVTTMXX3IIc/Xw5COqJXtDB0yf71LNlSD9JC5xYS
aSm/Qk48kVfg2Ix/+Jx3ig+8wLaA+uEPbXmaspwvgajoRIVWnk2hkVGtMA5TGwsf
d+FgpL7xV7L+kYX/Ok1UqR0EyquKbb4aejdzdid7JyQXhINonHIDoqoUcXarg+gA
kqkNBnRDe94AbZ89FFMsicYjaE07pJXJ/gJmGI2SWZo7aZTnBGaWKuqccFIWdpr/
7JRpWf74NshLv50QUW98RyGCXID3v92BPOQXFfgGy4H8vOTCHiJSkiuQTodwbKdw
+3mkxXc3C0H/+L6g0Q9MtyS4q781IjxXXy+UarzBwrrsemD88I94Pdf1pdufCyJA
Ld3u4srnguYFrdBjnZEIQY7Tv0eYZ3W2NA8OJyvLQKXTouLBp2guYarkCEZttgeg
0MXBAxt8iaBartfrqlC9rkOimp8f760Gun9m2gGgp6MUFo9WJ+jePX/KrRAMToNY
pCHvaDAkupDjVbGCd0dFb22S2iT6IMNBLQvI57jAVBOx11giv461GKWh7TGU9Qug
l38l/enQGfd+KG3ZYD8NKO7G+uxhdWotvRjuBMoMxgByh9/o5ynN9gG+htP1YB2N
uB70o4dZzYzmqsS8LC5UqMsU8Bg799Q1wJ8VeKO2+dzTvK/vA050CVWBt7AS6MVf
0QDuEJbrZOPTLkSquFYBzRbh+rq6/SoLxiITUy8XGKjS/qySybf04xiFVApOv8Jr
MVZbatzuCn2QlXm7pwIdBDzsaJmMa3hXIXaRzw47F68j3CxcZEqpM+yWDLEa9nyG
vgNdIs9O4M24PbFLJ7S/DKGky875leP3Fvd9wb+HZbczyhMh3yRyIiRFfG8XLiWQ
6RYo8jJECgEnPyVKaqr38FDfcqOFaujpXtb8vCLelDxHAZel+9BrrWv3hQvzVbRc
U/1XUyTxE+2/wwtik7v3Ba3h44HAgShXXXaDXFY5qfpGYMmnaVUCv7+ifEpDCe5M
+FQXnE5k0v5CQIQCtn0eL4S0RsYaorwqymMssabJ/Spt1LvRJ2q42fiZUWRtUs0U
rgEBtlFKqU2XYjZdHPz1ge493vrbUOWJW/jOfhF6ov6QeASA5Mw83mbKLOr2Ifcc
Pn0oHGFZtA6uAOXPJXG+HVg6r0HCKo/cQel5E7g5/hMuploTh+NDZT2d35kaL5j6
Vea1EdqC9jvALIa07F7KUAHXWvpPLyepkaI5NF6jGPnGai4WzCOWi7P+au6KoJ3/
wfRdaIGCc4kkXkgHSQWmqV1R2cIlJkuJgoaGiHRsYWYIRlaGrDMaCnm51eM4ChMs
4IwOAR9ottRfRZxPywCyNdQTrrLhfI1IiQUzF88u/oyIxKnQmHgzJpZdmRNacUL+
Svq+3U9BMzDsBmC+8r7bqeuOJsDJcXyBAumxTCVqZd7wDPb8m8trwAR5FFOvkmk7
rKMKgAFeQ4Oq26ow4DUwWSiQsSMo01gsw8up2p6okH+J4O0Z4+Zzsd8DCU6rHexm
KnpAJabdwWbnPQqwuTgVI3a0IF38qzqpWF57Yx5SuOxBRoNbq4hx7bRtmgfSGVgc
wy01vFcRpu9UkgnRT+jrogZDL9c2JZAs3z5O0Cv1n6nWL/YzBHsqQF84JDUT2pYi
zpt8Wt78toKO7o7Y+FeOFYLrjZqy/HJrKQAZnaMIUbv/Ppc2m6GZW0Dz2r867l7J
od482WJKDARoD5+bvbmFbOGxro+JP8dVuKQmr5MbS/MKkdJVFTn+ILCS1VZPT9Z3
kV/iiwUe/VQhDfMPM8A3MHFp0vpNv2bfjIu7HU+YImn7821RYpLUwLd7+IMFktex
RBBKy+/D8r+nXTiEmBQ4mv3U1QXIF/z/d3+b7bvqURw9ipcdIx8gxWAWY91MyvJx
iiR5PKcGAOrE53HNRN8Kn+RVDiFIDb1vE8ia6vQZGAeaCX2JWcHcD9M7UwFi+JMA
QCTOKGHsiXa1S/hRPX8VRxoHF8RZbeSYg7LC+Ynl5A8EuIY8wLOps5N4dh1TcZwT
0JJOo/Q1DrtPd08CfhFLf1t5cj7fOxvNMf+7I0uI2PKsF8zBmsBaMH03HZpmtj+D
p2Xt7HO5Vib9uqTLYic8RFyWHNt1OvN6ZgXSf+5guGKle0ZLQq0aP/gXhPT1qyHY
4UEtasa2qm8B2jSXkNoKfv7/VV5Zt6LEWtD0xIOFpo7CRE1dTwm8GBo5OkKw2SOl
EpAeoY560icC2xLhpE6QDrkjMJygQcW+1CXUQJe7P8ZnGh43eKBQOEbeWRGnS1aC
6c0e36Qi1a/1Emm3NM0kBZPHL3xViy3GcE2luCLcKNOtd3+Qw3OQ8fEOUZ1bTVZx
1dTShDDuxxhu+9UztTW9s9CN9OTWjmoqFaHVqexBsBwugpnEFFoIArZWSFjtl7sv
QKPXhQdL19aIfUg7SMPfeB6f/8qCbG40isjiGsczaEFD7c4OlXWwbEGpK2tD1ph6
aMtYWFezP9bTHU3vrYue3wZVeHEc22+zjf5ymajdDYruGRtffCrUrWRrr7/Hiygp
52sY2hAn9D/G9ntan+5MkLDQGnVcDSZ954B2zz+BhPtqFSq372IHGjFd/oSvonxj
O9TS8dNqQSuAgW5+JqufN6rpGVE/Zz/dl3rznkZbI0slTPkqcvguP3W4K+XTtPGf
HK3tCPXk4HhrdZQVHdmqA6dWGjHGQESYjFjL68ITwkfDZ2LrJxc90pUxIoQt9lv9
fLWqeG+duLWgoO1jFlol5FmssgvIQM8MeE7g4EmslTYopvjWc/ylpkBPOXPInvIS
wVjiVItStMBvF/SRczuHZztCJrIXEDozbe+uOpjGrfcGXcG/sbNd1Eork1TdqZqy
iDuGQTYEde4BpfDPVAwqQEJ/tC0C40KQLnFdQhW3eYi97QOUf/q7qfLT9bBTMwVe
crROIlPHS1XLnqz8HoeL+uYjL1nzscrI3I4GAl8XHLW+BzxfPJ5QUNW1jrPWnXN2
0paF8ya6fxy5IjjWPGRc+Vu0XyPffIpShEmtJIbBcMxU+4w27Wxxu54fTDbogyn8
nYGCizzWav9juUO++DSmjKX/ZxathEviGcfXEpNnzzKxyPwwUqUHW7fGMufXsjBI
E9tgyopgJi4mTBMxfEHJ/qTItWtoJLjHUKd+jvgIeSvDfX1cN+e4d4zT3IFd3qlC
hDegiOv/YMLl52lirTQb4Vw3yj/frHupoqQTozN6P/cm/5/NRkbaCIitVge721U6
7xJbXyM+i6gPm8Yp5sVON6BHIPNmQThz5vB/cBOL+dSOF+pHDAU+pUrMYNQ6faCz
jfzHzugUlOK/8L+fA/c9XUZdMcJP6bCgCrN9y+UqL5EYVV88xmxS4d4aX94F1Xmn
ZP5+Bn9NUAnJoZbKoMQFD97jRKAT8EwK3l2KcpifijecUbxKRS9haoFmUzJQ5FuU
L3BJ3WACB4GM34DQN3l9c++5rE1tweQKsB0ECL+YaZ5DS7JTcGFMvHVK2+kG2N0N
PbrcboC1+lhidZy/Nmvs9PmOwHKJKp1nNQ+dyHV93XwZ02sD5/aVoZ45OF8mxmlo
nBu7g/97tCi1eHQq19wi2qN+2tMhJ8gKFTSXXD/qrj6hwRSTLYJmdpQGiJs+RQyf
l0j1Tm+tBvJ7PYQj54UB3EqGIwueUa1HOl26Po8N9pL2qmZtfRMMLfHrT087Od7g
BL8DqTe3Mq1kAdvaDydGLjTBjiy9AIqUBvarjLrf4H32c/Ox+pe8NUQoCM9Y/4gL
g7JZapBdPjFAsM+mWTB7nfZompus4NZKQSwnNU/mTxXsbPG7/K8Z/Z62fimyhHYh
tqoglYkoeTDQs428WwbRz1ox0h/MVZYMhuf3oACvLioJFom8+m7GRko6wGDU/Oue
RGma+phN4+Q5xFaaAt/X6DN1SwMJr2JOKiUILHRM+dRsUZ2S2Pmfrm3XpQ81bG3a
lMX6jMRUhJhOW2S46LZmN40p3PPY5vmzX1PnD2/Iy3jTBcdDw6WxAYMQiesVJ6mx
2MoXe5dWqhmWH+0FtgfUuu0gTmCSiS/z6dOoD0fvFK+Q0NNvt/pYRmSUEJrDFEfe
WdTEcBXPKpJ6Edy2RZe4e0zREX8JFBAdMsz0aaR2Z4/LHbWUzarireqIh5FPvRUL
qCaUU1i3WuUR9zzea8xX+6XbEHwtLU6fvvd5F0jte2OMzUX7OutvPi0X1bFHXo+e
Jk+Qru80mm+M+HVfHselQPaY+q0fTUNjM12+JFhO1JG8psegIFKWtpv6AjhqZ2tF
wjUQT8Cb4ZFc6VfSkQiVEB1jyWMSoS5l2cYKcSl6c5YRBFM+AeaTuLUsUYUuy3s5
psQTyQXdnbwblCwZhh05QZyP+MQ3oQCy8JdvKD3S38npnusUwuHjm3pmsZQ5wSob
Tf8Zt25P5geDSn6GjBMx8CPC9lyD3s4Mu4wJszY2WjdzsAk+hQN3gQt+ld2GJPNq
VAl1i6Rnavw6qLy4Aney2d5xHvYV0Sae4KWm1ap3GQa1WVknHdSk3aF5++z2bWOn
l8l6EU7rVZ5OVjeXT1DdhAUQRCn9sACSCP+mFIcNkZRXzXxdVUlp0y5QsB+xI/uY
VpQ1YeEZWth0qSS5LmZwx6/loclMQituFm3gcsKhBfPcM5fEkKxjquhMH8KQODUM
W7uAEy7eJGT25DnlWp+V6pr53Hr1v3hUXCW935GzCnf33M9xGWUqfTFnzTKjXVUi
i/3VE6XC2b0ycSKPEbNawqTiWr25uHF0C6eCmI12tn3xaZze6yUncujypkelaiO1
N9mnerGV0mfF7AT30x9K+SoPyrlAPCY1DBbz/5zjvBTBFfBPjdyZSRNwbUORC67S
3QEeygn+TTksNhNSWYbvUrOmmj9lsVQGUK/wmYrmhU0QoSWgQBqO+artpjtUwkaj
td2bOclRBzmKnMDRVg2VNYe6N8Fvs2S3Am6oh37USjBtlyba5LoRSeB0EtKYjS8K
iNloNicsT7JzwBhR9A+MWwJxT6im/Dx2B07uGUTzibkXQcHfbCNvF0Dw+Jd3sJiS
fR19gIzyK9m62CHofa94cK+zwSdPNTbkb4HFJWMwsryHitSpJfLE73VyfZ05EO0g
T1au5X2LS2l/9F7r3c/UWwsEikcpVPAg/WOKlQIj2UXLW9sDlA6BKtFS3TJtggc/
cm3Q7JApkNbx1FpR9K3ykanr2nSFPrX/gEEd7KaM/vMJo5GRYPKFAagg/7VjJF2d
e52X7EYwff1vPqBZRvYbQn9DqEn3kYxIask422dBZochcL/lKwCfCZdOIQx3d774
s4ZEeLyY8iHItCtY/053AgUfJMFArjAEpwbqBARQwdTuHB2XH5J4sUl+pKL4wOkx
DnMFJoqhtH/A7fzXG4hV/vSMtHWmATre+wT+8nLy62XoNtrl5ES27gsCcC/o1beO
3HqD+wsgecwE971JX1fDgH2h/JayOc/7F/c8Rytr4hBMygMGzYipeKlr46aLOvf/
NsxLXn4KmdWE/Y65qBKrPeORGyx/FTSqt/zRxL38PkRJZFDX2RqYza/dNQOSz+C4
U62NQ+XoZbeIBvcN6Deivn80NCajrE3aKx5Va/ieSRjUjnNzksJK0hxOBQY1pSKF
/tUpmCXDcqpxcXS+I5ZQvztxJiFMzfoZ53kNuCg0B81A9l4iah4lWboF8W1kjz0U
I8K2OY/642gmNTd2pCeYo18HpgJu6pQyPiT0HW+aWTuQ79Wg+7UIa3kGZQbxXb72
iG0vSQlDkFcJknBTGmqc/FrsvH5UkaxZKjUePVXMo4NEjbv/le17nzq8w6myFmUF
cNRaKVHGNlIkOiMYBu/tVMIvAwpMHeCi6WYNI6ehHbjv6n4DDPKrjh5M9saYFLsy
e47pCLa0iUq0CETAFxwwPbzND0BCD+k0kgaj6nowww7qKDG8Yg5ynhhOotV/QiZ7
5DnpJMGCKWuKG1mNWn3phUg6enjuB0Mkk9ZzULHLp+KW3f7pTuPd/fnZDnzooajy
wTKR2PVw1eKFUTN8Ftzcper5W0cQtvrv5eY+CtuaSSzVviMLQRzH/hnU//dbfA1S
/O9+LNQnFqcpcsNeVrilu2yAn/JnLi9nHKxtrXcq6wIv3Dh/LglQV5YoYXB+U/lc
nq38rFSAYvDbIdrzcghIBWdBGKxo/CKDvtViSP/I9L5PMHaogil0TKAaRuGcNcES
Ypd5jGtz2174fu/2FICL6q9/d+g9SD+v4IXqmLUblJMlaKADa+7QlBjeDXrFtNbX
9mnCpavV0EBQ10KR3cYcdNUd3vVirHulG6DQMEY4w4LvmLLDHBIFoQOyb86Idozr
9l/K94WILAnNqWbs4RN4R6xGwZO1Y27WUFnsaV7SvnXtYcirBmIAjv1Ejr3XGCYw
oGiE9T70nc+L+yDtYQqqo6M9TPQIYFmpgy3gXDPQAZc+YcAXA7cB8PzizERZp5Fq
D4vPl0Z307pVFtDiclARD1k6ZFr5z8SjVtlwkZMbYwAJfd3IV69g3LMq9R7Oh7gi
hHAcCCFwo3zS7TVJqqxqjUUvu3i2o5Tt7iFquZfKDD7D3isyOkjADIJNYWyqa9SA
Mm+6Bdhj6oeqTO3O2k3irgFA1nV9GMAJOaaSIBwyr8rAEEyCSQnu6cmvaI584/Cs
TDgGBYjsID9QwVJzOF3oXpoE7RvvkmvnO2JfbH+6/CyLzxNy8SiC4IlwQaouvKvk
boJS5ur4Vhxj+T17g3UDQ/VHZsoRywXBRZ3gCC/H7uJKJx8F4unulgN8b/yIeJZm
b1snRDKbTNl8kbXD1ZKB9/m14SG8Rd3CEs14n57T8j1gKrPl7JaUOCSJbC3eSJGJ
OgbrnRcfoXe663Y05lIhNmsEtdjviGWvHVYiSimIs2Ifq8OYLzbU0BU2nJSGD48U
TbWNA/Dbde854XUvzF0StPfLtZ1NrA6xST05M2I+dWDZ/pNRWX3M4pu2atQiJLka
U2jUR5b6sXVwB89bHRyUDwigE13Mcs7atok0a5oQsAgL/ftXvy57xxP0DbSxKf81
a5LC6YALFK47Luggcx/SLDRCD2UMjH8T6YKx6/XBG5YCPv99hM6+nXTm4fSR5D4N
yhQI4k5Np6iUn7yhUa2xSmKW80EuwuZrJAYIaBuwrOKHM2I6A9sGwxU/f2Zbm2Dr
WadjjkopmhyL4Jj4ysZ+SMkJInLI9/Kf9RfZFyf/6kFukLo8s7rKNXW/JwHclddA
Bf+N1z8HTXSKkOACeO8qooWG5bsxhSGp5L06fXQAwJmebL+UxRarBP0UhU90iKs+
jDdvuZfIzQo3HgDsFPvT48fv8eR1DtftqE9hFGVjDkIgEhB2MAOG8+bDPyzibL73
orjF3Hxkzz1viIc4mMKY0rh4EKEPRQmwu428Qoul/s9Tdsat9yjCEy6gohgHcdbf
wpkioFMdMwNADlwd8Q8c4Ebf78MKkgwDgaN/DkCiyRevreJlMQKWs5BaGaKwHVSL
5fREYJfR4nDubV8bct2BgOvAwY9V+BESRPkj+aTbZ4hpAlGzGUc7tSnbw48gUQSs
8MlixLeTqZIgfrs2Vmz0NDCBea3aFjWj7YnxkEyDsGeTTotwyj06A+tIeuuZ40CG
ga0MaGXc3B2BuY9Iez3RxSeoGHQvpXeVEYRwapiV1N/xr9nNuMxmgim6tk3pbjvH
G76r0bkC06+Bqn3a7K+TGTE622m7Yy/QIkO4+1gI9/oNx1ISkpMFwSOsZ1Q9T2ah
c8XXyGp6UZv6MkN9M13Gzhg2Q12R82iyBWmVp38l5//Y4+z7lMcn/oNPe+K1sWYX
i4dBsp7BdtZGpGt5DOfW+vLNlA3q18z/CfD06JLGhAYshk/mp+knhzmUFEmm2rx+
roh4FUjKdPdycqrY7No6Ll2mKe76n4fZ5j1hKIM/cnV3zTag+nhAeOqKJ/TSc4YF
U87keHeRT0BHE65mMr0t1KIJa0iVg2fuXwZT9HuVrnISCUDFzga8P8mTRe4wFnGI
yyWMf+TaXkZp/2LlnDoCGHYh2cBJoXQ/UMO527iyQu/8LbkTQbJLBExBu7kLZd1t
QMrFp7cKE/a7DkRELvVSnzLJE0jZm82hjBqukbE2W0PhvdUQbOcgaVjdF8cC+xZp
9+PWH01TY3Sn2bEOqsUyaCm9ClxSe+cE+Jx6qj4Pv7+OMNyUUlSJVx86nQ02HoGr
8KItT5FNaHTxFsNlA36fcguw9xXW64ze0RrKHJlVZ9SlO9w0u2G+Hb6EYlxJKh7F
Dki8AUc3nINXJR3yexr5HwoFzdvku8SQ3iVTNRubayhZ9iAlnXwWJyPjXnertYLS
OUh++KO7BComxBB0trmS49GwH9XZli6W1QKLeSqLSDRcB//UwMJP46ZWOQXsYmUS
5HOdlqno2mTCAC8FOMwok30uDpBHgMRmerlvTy6iNY2cLjXG7npItZ4nudvkYVw8
oYfHAHQbO+eV+UhBHh5bvkPu3WlaVEu3riHDe64gyN7FHt/UEkcGRKYe7jbBejlf
MDUItRXrAXrsrM87KuxwKArmg0oL0vpc4dQjhTY0Ay+Avg68j5ga0ujPId5yEc2Z
aqa2jHskYNBkAYlip8ZSNBOOTWa45Rktf2MLZD+LAJT02okge6l0LAtZ1ct5Tsk9
+odA1ML1/1svVGlju44wslF6inhJvydFAFnVg4sDdnzo8FQdvaCGNAMpA2PJ2R/x
ROs3DQmBl9JBdYlQi7bkIDZTiGvxv+LHLJNFShnF27UNqVIoUXNzvBDbt0PfmBqi
Ui09lc6UmCu7ijM90fRQw1Dfco20GTz2M8urfhffS/u/A6vFZFMec5X3M6upN6NQ
faI6XthRNO8HOtXMGMhqKQN/0Y4umqerQMkdiH5CqYA/fVoc36cvzLDq3YnZ9qca
mAjw4wRAZVZpwibL3B2LTIsUnPzyLoHSfygPKjGpYA/pinG9Q+RgVJbHS3qaRSnk
GnxeKTJOeFDDoA80cbyKQZcDNRO+5BdFByR41JDpKLjqu5RmnbRN2OwIh5LC9+7+
/kyFwME5UVyWYlW8FYC4tlksz4qNcjquCx+8LqjUjoWTGML2IdKLNrkH2ofM0azV
uBeMs9ZpJ6w+iJ/x8ADQ2Tm1zutyk1EIXgoA8EQ5UssawpKplPKRaaKNm1OdhRPQ
TO3Liiw26c5/ADXAU1jUux703YXEi6qcHsAMyEb8FELg1eQnQOIJCc46itCBca0/
wCETJOc4gJvuVql5N+ONmCaEXWb4Oi7yBy/6CxIP/Q9dGptdKMJ/q6iS+TQfOxCC
LGvlHqtfElS6ErT3bG6N8zrqBIMWwMloDkztvw+NnXE4iqJihpSoTOPiaKuwy6qN
oCTetn1RGp1y+aACWTV+DP6QZIoDc+KX3r67/x3ud98vF58LYZ5+K5vnJnj1/FWP
WFZsnOHQM5OBbE/4egfvG1v5QriZLTpmXjTUvoDSpg8s+0gad2mwh7crc0cS2eQs
Get29A2/tsL98ID8oZ5qT95WAdTXg+7s3SBd5ykPyoxTEWLOHUG5LtVyupl/6JrC
0TQIpMQjNXiGYdc3evT4QM/IFZ7YDuK9YldnLqCU8fFAYXuorT38Ucb5oGJ0XpL3
OvwnDCnHmHxIdL/bMuQGb9W4m7FV8ED93Yf4I3x4d1WDynfo4/gBZCR6yXUMzWbe
l9akVA3vOYJ/rdDiViYue3po8z/RYz/LI9uoO8EA/7TxutVZU+/oRP43mxur5Eku
+Sa+lDJD8wOPigUPD9C4Vt9+ae0PXolbsiAyv8EJPlY+d8hevwkqhBuvV9vwZhE1
vaV5szFJIxRIl1KacY6qh8hvxV+/NOauZBPP5SrDUw+uGpyu/vkL64cxCDrvo7Pw
Q7sf5/BghooEjwYYGLOcJJIvVSWN97SCkZFkcknqSdEAfAGHFfQehC2iODuIkhjy
BHcdB+VVdSCE7baDbj0xjcdPF3MKPcA7EgepqKzsZbhtdW9Xm6AdCPRQgD9lVgnU
M8oW3BFYUngkgFoxYNPdWF/ry1e5/FUhe1xmscdtaihp178Sm9dCeFjHGUD6JjdM
iQ0c9HFZDO5vH7P3Q8I9RGebvEW8QzZh42Ze7QSq3PTiZAzpeW3Orn/vqUJxRyaL
W+AlHBdpUUdTYsyPiaITDubIztVuOb2jTEApN5TCuvJ/3VfWNp1gD85THeUdhsdP
jsaMuE4VLnTdm6ZnptlXpdVZWvQn67mTh2rTSmGLV/4tnPPDU4j8m9W20J6tvRQ6
218eIYU1aJDyRgdwX9Xo5MUG0IovikwDQ+4fKDIxFaoDZxPR8BCD9jxPSHwl+vkb
nLXzH+aWDW/ZPKKD00S4xIzWMqhlW4FU+Rvvgo4F0Jjx6YIjK2UTsS4AaTIWRr0+
JXj3CsdacQwCEZeCVMBH5yrC8lr7nr892dUb1b6LMpFkf3M7/UjjxP4eYf12ssOc
PYmUcEZVyWTHRFXmF3C4Mv6L0Y1e+BxtuR2U5gVRwDAbjRUxmYBqam+rF3YaQP0+
SoF6VJU7gEbvE/6SkQS1NffW47t8iOQYoYAUTMIfBJBgmZHX2QeAFs0GHyFKL/0G
F2coLTpqI00jWKfmFevlLKTqjaGCeweXDmkAk77o+h6tJRTKp0s18pDhPHkbySQy
PqYAwpGJnPG/53kUk8GLJkLwhgD9F1sEspk61zwAvt94kbnYc0k06nB6VATgdb/h
bJz2U6TCRwDUU1X9sNKyDHNwmlrHRtcVBjH4iTHzXKWH2SmsMRQ5a2N7s6C9Udhs
IrMMdk9YyGBH4pfE/1ETlj3+wx8CtCVQYk6Ob7YawfIuuoMx+zglIyGvSU3vFG89
rWbBTh5Yr93V/gY3QY4ifvWDFPiTFHC5Rcf7p9ps3dBEo5u+wlBO83szdjg80GPs
XaXQGcNfor4+PHi7K6Ny71pvWXkrfRK/v/SmiEHZgXm4v5Tys9ueoNvRLsBi9lh7
R0VBOz7lE7dh/Oa5vgCvjBbdICrP2fOjHzBYzmRNTRd1nZFas1NCN2x5fy5FXB6i
bOpvP9GU7MrRrRLdawCraB9sRgHEG9NWM4OgoojZU3L7Qd+jH+Fn9voTH95UbWHl
h+pWDTEgEK+qaDQXPL9uBZAKDGTuufQOlt673NISg3bFMWU9Dq5HHwGt8EYFHgzl
3vZf0ztyG5WBgrcW0kA8ZaU5z4JlYBQCEQe8GWI21xttxdcCANm7lSkXvzXxb1AJ
iG+yTdnxRN7nG63CUZPf2xlyzD35RM1z3PSjQzzmNUKv6nSdhctx+UK9Rr9HfSp2
qhlgpLqU5XmpvVFKLPlAI/sFzdvCaKN9SnfRvx1tTWqGDt0TpL835yZHGSWwjx/f
Ab2OLo3iaOM/XWch4YtYBuTtdYWNOWuWYf4m320Qqgn6vmBmfY2I+vFPPGgCaJ8j
xYL5tkIsu0xjN2Uf6Ej2ZrBytSNNxTHn6J2WOgQvVHrvimD6SsK0vHU/3yQ9H92A
S8zf9ujxyTlIT0Jf7RihlYSKkHn6x3zDSII5XLAVC7KPg9eYmewHeYUJjfi/uhhU
r/MSn0obFQ5FDjelQVBloduAfrIQVi3Joa/JQMAiiUFqxfZKpC5j/VQTVzyoKcPB
TjQIZfIJwGRTcbM5WFnsNcAphKPAzX+Pqn85rizdwWlcswzBngF8m7BSO7Qldhd+
lnGOgPH52A9yw1fleLguO36Gw6jIhks4EDki1g3CkD0DDEGt1Y7KayKa0IAgxFIR
p4npA0VskQhkrPfgxM8ykwkLoG3URgAdDaJYEBeWhnzm3ZBO1/aE3wfkIspLSnTc
EMUtkuQcFjCTqiVr5MeHEZ8X/wKe2dkrFNxY+QeKTLG70266SVuNE9f1JglhvWI1
DHTjkrpJaeAyGPSqGuGxIMxH+Uez56PckNQ7htNHm51ab2yrIabeV1WKdUleLl4C
tNWs68GLswwnG0onDTrjpg0UpD4BB9DkxX023qSp+LBJRbIPFzmeXej/VJEG/vbv
bw0O+sG1sXgkroO0sV3CVMP+Pub/7cQVKvQifsF7RxzxlqKxVr445cdfnOhLro4w
P+2tB9jWuTi5h9ntztzZ6NOWn3fft+JK1FjZmZTCWOhRc5Zm2BtAWr/fLcAXDS1e
g8ljOyzeYEpwp/8lIZ4j8eA0XWNX12Dng82axJeX2NWrrwGxrZa3Ybcqxxu8tLCq
5ZlyBHx2QDyfpMDfHnNk+cRsmIx7xsfvi5LJUJEvmmVev9IhY5yIjvyhNVB0FDul
YRxgzX1tqqn2IomxyJKgyAprUw9flAMBESAWqen4drilfLKNm3zfOk3A8v8WhKu6
PdTCSYhsecCsPdxEci/ieBjcWN/+lwdEMe09v1IGkZI94nzlByOmvtXM4bkHS38m
csoM7HpuHebmhYdn9WbptRajO+iO9wLCy6YH0Tnqxdgdqw/YdKLgXkPdPkbbXQdw
E6BVTLDVTlXfF26tZWpdN3jVdal2uqvA9Yb6OO26xGejO4VBNetjEbUera3cugNM
DHm6/lH56cFxM7UNHmxsNjYx47dxw+5AE9yoGHjaCuiu2xjsK0fyRKj8W7ZAlrFz
dhw9yewno8wmusAbANcVZNfv1loiCn89MN9sBEaSW93STg62so8xkUfghr4NAoFj
4dgnlks7wcD+lncBcm9yCrunDW1QcN7hU+wBCTm7jGDNIfoHluorjPBeQYooit3V
L9B7KsqigA67kpK670l9xS5+F7kiX66bPfl6cFs1D4Jpc8Bv95NkRW0wXaXZRGE/
H9z+0vpN7rzB0cEXBf65aoThrZQMsLingUUuovsG6UBvQjlyE213Q7S+q1hIBtX6
ykHVCtLp1qRm31voWB2XXI+8FKCHH1XbHFsXsTPGpxM2qG3iMSyULVCHkCJ7X979
yZ+30XKo2iE4+nZ2Uo7qtzwnDDpTF4eu/yymsht5AoOhB90AYDUucy57dXydlySJ
XpC2gatibF1Y5Fq60FUARNW2RjHEV82ClaOlN6kX3mcnjDf5tAixgj8yArWvH5m1
hshYIpvYvuna8WkZPV1Oyh+PBzTOYIs/YWdgGiOYGVZwuyLyD1mUC+SNt3wJ//4N
2bbgEVYrMGws7Uzueh+dWACuq8dfTA1q/9+YEnrhL1fgA1dYZLjiIEva/9/sLKjX
7yhsLNF7BtuOzCrg0C5URMymnNnnvRPqPN1jLh5jqLNt7T3b7TPJy/bXPgtwcrDP
mOX18MbQlNNdurvTSzMaQPq+Ceeur3sykvcsSFMNl/tvYrJfHO1ayf20szBpASQs
XjWOCG7I3DTkhqOk9RTeJMe7Fuq5S4d0iIxsz1wUGeHsSjihfG68JkYj2aNDAClw
3xRxLWR4tdWCgo3FZ8jl9v/tSAEIhRZXuYKnZfzIfyvmNR2I803MGiB2VU2hgBIp
+5Uj/nJaqH/3UZL+DcT/cmR5Oex64VxKx1bnFfwfs4HRMnoejlEsTe7Frec7A0zW
HwCGnQNolqPUOPI7LPNzWVUaAM60WOTmRXtNGEcqxIa8zi1X8Z41+DVBizuJ6vMv
jXn049fQssbEIlKh7uwMI1ZIDw0cv5WRif9pNgsWkab8AOn7kIBJyjxnC6CjTnc+
VuFEFEV1sQIEBdm6rGFP7hoHPT1616ccAyqQWTRR8kxQjkc2wzsJPkX7CRyqgbs5
BpqAmKDktci2Vh3Imhh0u69ZpbYj/hK/sUS7s77tMXZYWK1vwePcMtfZCgb4M839
SeS/pMCzhOnMLIHflvV4Ty+2WVlQVmtgMPzyv+W0gRwznX6WucaSsA3fxUNHkD2O
hxUZJ+GPmPTf1s34USGdrtw7msgQ6rjlZa9yk54FJHn8LXngNxSFAq0NuGVBP6Wc
u6C2L/VGaHecyF66jvlMOQdGBOZoyP9WmNNQWGBpnSl8tm7K7OI88NqLYVEUNqEK
M/IsdGKtyxKuAV2QsBzkni1/0380T5CiQKLBQMA4P+zdsg1A2zT1Ve4gxnJEzTtV
QEA/RnwSnGnGTfJxVQ33jrCyVvYwXdwx71Ut2Xj74iSILqRPgRL0CbtURQMEjLXT
U495Vtskgq5/NjkqIKtiLxVW+BdloXhwrp50lw8v0Rxmw94HjYcCePRcngXZNEhY
nU8soUAU1pI5Al2uFmlhB4/m/RljNfq9YdOtgQvceChEq2o15GrTpKtsWXgCTsgF
kigPJX/hgI4NjpXxbJpaKsp8meolRBHYI5m0bgjFC56FD66et+717NW4Aj3PFlW7
s875RlXgNCVG8HpTPxtEbiPy0/lIz3zYsuNkDFZZbL+LFN63z9hLkhzm9H8Wkywd
YKMLGIKgPwXCyLRTY0Hf+ENXBPhWo68hkZ2nj3ddGYvUzydv/nAK3LOn2Zf5RQKw
d6Xy0TJasEeE7CCaH6AYQpptxxFQyQ/yb1H7XoSUlAkH46Jk4bA9qkiYhuNUokaV
6Fnq73bJFkETsflAEUIlkHmLAw/DQptwo8am3SxMRJgr/68IhaJVn1X+CsYRCgpy
msZDrffhSjHxSuY9DS6CUxn455pWZHThWZKJv/9eBVqUy0/OF9/NRfBek8Sxo1Wc
WBJ9+y5F+rwJTNv2pR3SD6cHO4oe+MpN7eJ7GXD6RBfigTRaguF9m4DTnqa2bhEA
C2W3YEDsA2WGdNe8z/z++EAsGZ00+3vhrM1XHZ50SOxguPQMAJsBBJl4VVfrEKc2
/1ksq7PFBQYJTU3lExP1aTUF7ev64iqUKavtxgnmCV6eGXGfJ1Zcc8TCrQyMfsIO
TaykDWWAxknYZu+2hnWRA//C+CXe8rm1H3OokrsSFHhdoUAxCNjiYv+JIMyO7jge
hDOaWt/e3nRidzOf8PhzgQfalkKeESY+bbHldWSHbxneCnD/IQLq25Xqidu9rvRW
uSsNNGmzj/2fznMvyiLUn2nKJNMkVjSCp7kTEROLLEQvM0qfHE8q0Aaedajisbqp
rAdVQnAijfXJ329jiPS8N3YkAvlB2PP3SWlNs1i6LV7GxddiYh/tGgvXG72X4bW9
67mm9WrdgjSZk9UFoWjJf0rdDyS/o/X4bZt/Bz70HJp3SHIhvKe+wR+mJns43afX
RSxnWLI7C7M6xPBZmlfqjID35XCIsjryyVa7T7Qh9G7agYuHOEiCcuPzmS679WG0
8iBFjuScMWI0y/FeutjDdcg6VoMQrD+vzlRBRgBjlhQdvY4JZNYdXN8rFSyIYCkH
jFZzLtih3IqDj2IFpbWqDysBhevWScCwAEwRmkopw1b9ZoHniSYRLCmBctqSoMm9
fZFLUq+9pCRum5EEMTB+KC5mSUzyo0eeaGUkZ+XetKinA5zvVrF7ExgYpdsBHVeC
s5b9srHG7Z6AQgXJGPj6scuKT+u3tMz41QgjIiks3pDeLypi7qQ/MH3Ilgg33+rp
AQOYi7CPs/NNmf04APc9Olybhk+JZMyNy7R4eULYIJjSyBjdamLlrc0q/jCYiLCT
SmyWkjqXjFwuNpX1lr823+m82mF+qMH9bVG/Voe038/nAJxsyMN95u1H++pBbwMm
h3nzgI3WB6aqTJbg86hR0mzZ16gm2YUBMeezRJcIJsnzgDQMWNkRZpdYrT43AlIP
oIRL8tvsJKhCpR6eha5s+2x1GLugE3cigt1s9jBssTx5RXuQqFiW9i0G6pcWRfMO
USYwgU5SIGnZG61D4yYqI3f3esbfY3W7QnA52xF07HQnx0zaPlBO7Rp1edXgPxkF
rDEFzS8nVOgbDFL4Vug2MxIWwXZIwGXkoF9OCgM52BJ6oU63y0R2Gbtrd6/bVdzK
EptPfphuPEJRCeMNTubBheVRKqbxwx7hCo1CvjwI3bLrCXhjUDokbSs97FyO9pwP
4FMD4SRBFbLW0dYV8q+/5jXZhEMW7Xn1E20N4S4y//ZyG7YMPXZOT2IxZeMXapfC
AHOiPw+uAt8BTTiCZuOLsIplAcukWTMIxqJ1DDuc7x9Ri4/vMGaQkY2rHxeRWVhs
DXfIml6q43+ytInfLbkGt+zMD6qx/6rlnpErfbCB6C3Dm35OgkCSfSd3VSmBzbrL
EzL/1+eQrwaQmiiy8HK4H2ie2XQrrIvPaaI4f0ZcNT5hl5fswwlIgHVxnfXO6vt8
2CWmSsqjamyiy8MxPG4Vpl4GXOsVE9ON3Ty2BQXYb0LQGNYfazyRReACxYMnZfLQ
ZJOi1ODLRtJD1XJsF340XpyYMaevANnFQV3B5xdVSKTdMl5BVvySfClHVtzwWMW0
ICy33Djeya8tV069hmT7Ydf8z4IFkRREn1E7vn3LQ1E2Ix0x7M1mjYngsiZDSW+1
P0rbgdgwzVCdev1tJyvqRx67mNMK3PZnTK5yHHRHIxF0KBlH4tYuCOlpOWIe4hQn
7arByARgZ/JvMTA+/DP/ArA3Jnf8SjFYFYXhzyC6E1LE6HSFjmGq/Lvjme75IKpu
qbq5UNikRlsXQ0gNXZ1r6bcIb6rxDbJio25MQ6aC5wpLHzk+gfzvoSz9L6o/kti6
6p4Ki2sre/hlQHDvxLIBzXyFilRKhuCGqlhwMfdr1iY0H+tZi2miv3MDvUNlhdDQ
9RfxoeN5UN/HwHR+C/fQjVv/wQk6w1+LGheJKLi6i8OKdzHr6LJzQXdIpb+mZl+M
PRvBU9Odv8maM+uvVh2qKu1r+ltPx93DVZ97FxDcLwv6VQxlS6MwLDX8l8v2RZZM
tDPWZaPcrsfVF2jRPe13Q6TNMoYsJyQ40doU/SKlyqY2RbJhfnKCEoffgxadm0zm
UOBLKpNTLU+mmjiIu8JxFhwFhxAINqqpEHeabeEX7k0qS3FJtNktItM7su+Vg0Gh
Ldkc6ehYT7Y4xOmBezYSOfvF12G6LnL70XjU6XEfq3gdq69AKBISC8WaaPNBdC0Y
8Akqn1ZOqvM0xnmHtYakq3/knj7T3GfzVUs01nobvCIoJi8WmiLBobioqpFjjDYJ
csiUC65lzRs7r6iQHGvShfcWewvlibhWV0WdseWdG3gEJFeWoG0g9uAmHM2XZXnq
azLIRi4JmNUeHrfi2/CjA+UiUCeauoh1znp62iXdXCfvdF9kNQgUKg3krsK3e8+1
khUhZdsqwXajdC6m9tFpN8EgIjGxZE6dAO1kdWnfmtpDT2WGQJoMOFe3shEQ2YnY
/1HSAPBVJOS8UmwZUNjhSM/MtxduhHmD0CHvmSySU6cdmsSvrezQYuZ/yUwQjiUO
mmOYDPX5VM/JgXrPvkrnIwGZf9MgpZNYgDwOOz2C3eWbd064pwikkMJGJHjbfJuf
h6Y+9hzEeSAutClM1YBHzReukGaYkgp/v/KGvUJV200xptWYyIJ7L+t1E90dYn5n
TpaPuJzWBK7NvuuQP6nHAu87eulnsFvbEpzVkDXN8LReSopz/GHvQZ6Aaqq7Jdy2
8Px9ZSYcwDfANvLCBmIofdaqLV6IbbL7u0srgHL+pKaGej7+4oWiApTSz1mCLfFw
qUAbJUeZSW7y/vI02dmQ1GVf5+UlATO6cA7cQBujpaP6Ado9wH4ApfIvSEkjqXoa
rcFIa3jbe+oHInTvV1VmAl0FGK+zhE9HQ1klR79fQcyeqj++crjjUx44IgVBhPbD
IvaAu6v24eVr56eUGyrh9GtRkVpPcAht7XVWQWgEXPu9rUV+WIcCadSqxlVMgW7t
kUSf5F5kwZltfhj43VuPJ9S42Sz17MQXLj1kILIbg6YuQiyF4TrROAnYZbmK2M5Q
ZWcM1dogr4CFEOxOIXYG1kR5hW4b/4UzXK/oR4da+sGGRB43XFPysRkRkitqFbwM
IRamyYfXGChl321snSGSKc0cy5+OnRIz10UqLquu86wRtqSZ5TIiGXRMkjtZjr9x
KnQilM1eoK8YRpbcZ3RdKcklXC30JolhxZFGfv8wR2i9p9f1g1IPVtNgFh23rcee
oDPhLiQjc9G+nTSd7JVgIXBdQA5rmeItY2zzjQd6Aj81Lk179zY8lXzOd7yFNhnQ
cAKnPeX8RQ/VWkIgccA/TO0NFj4vuiQbVL72I6U8RgZi2YbdG06ACOjwRA8KLyyC
Ynot3KeIokHjgrlXOo1sNG4UhzcNI74p+bac1Ke7BO3qNJ2xPJHSKyXSRcIgjdjI
Sr2ak4oAOjLjs/VXXYpc/YpJgZl6JTJi6qsaU2Wn8u2Ot2haBc/pV9SxAk7/2Fvp
+R3L3EuOxqIz7t1oC2HpeWJwnYrh2GmfZ48JgBJ78ERYXiUPrKxx+uLEdNJ0huqQ
vvpKKk++yknLQRZZdUP8dybquFrACvqeRe7JQo4C+Jzla+M90V1PA8Eb8HgwO1oQ
D+DE35CN2zeY4//CKcmlyTP5CR1sRuZPli5FAV40ANT74q0erFDYA5QlY4NpBkUY
lAgSb9Y2ONu1N0U6vnQlIE9vooXo34khcXn8EeKlReSAHD1KZn63kApXGJpsPzra
TIbfeRPKRcPRUfpq35w8UdoafKpnWs+6mEfxzmHcGb5rEUBFLPy4Nyt7ELMJogr3
XZoHsZR3hFDbQs/GsO7Qo5XKBzCjrgnFwsuHBH9IdhMRPa/txWgB8xnVYPRuc274
196gXgeVuSNurXV16zOmRMvq+ipAl2yLVOMP+jqTGfycnZ0y687U80z0PB1i+tLe
ZG9CQuYTe3xpFe8Dh96nxcY7wqZz1Pwhcu4MHTkEpaR5tJmAc9TnOZPPQgGZ4O0X
z6uKTQOzJ13VFMVJDIOuCYEcLZeXyVMuNUbZ6qC61Sr1RGLohgSdHzdUlrCXGZ+A
Vuh18Hu/wLe0RwzEeO5x4pGOg/6rY3AxDjsqxjz1op745IVW7iiobBQUiErhtWCN
3YWgOzevkPCTqjHGs/+80QHMSQBcsBH5iM0paMLJFdbEk/GJ8ccgaqNMOAYRN3E3
yagJjqpxgD368CmzPUxdfu2IksvZeJWBBL7S2Keh2TGgxWblTqB9DrxgG+AHezFG
t08jsbTsKQ/UIYjTJgj1izWtlKCr0s7QtQ1cBUFLPQyl8dQvsnuCadEPrFwq85bX
6Q7MdUP6DC2wFqPPdrkED0IzGWLigGnXB4e8eHMUI4sjiRf2vxJieRFakdWyIceQ
8KB3SbQwGFp1SOltP0BFtXWf52n+87GRtuwQEPv+It6/7qvKI5kwQ/r0NKgLutVt
trm+zmQ3VbGWzeLTqqVmwhS7bNivXG4UwMxHtmliEf2ylVTzyogAX3axZvRAUw5U
WYFENVG601r479gVvPk4UIzrZLN3TxIzhCd3pW9bG/MZ3+iLBuj3Ew3Jh3SQX18h
bzhQoLdxIqgCVY1Uz/creR9gJ8eLEWqNo6GiWSb0+BLMy8w4q4si4N9bBBlRo8o9
BsP5ZIEIGkzolZzl18BIo0uJYszv+yodMALO3bnlncxtagLID2jvrmGiKcdAOkE0
qO7g8Q46qzZjmJaSWuPhIFdvQiPUQqAiWsLm1FmmhAyYdMBZ3F2ZOqPdZs4E+w60
8+HM19+0GD3O9e/TYX4V+nXwLtWQ9k2DwFq4D6JOFm1wMFUus+pOd1CZUu8bNEqv
boIFCiOSiB4ZDHkNDJdRoHzECe5jLzL4ba3BN3Jwtsb120HbbvUhiNKyI6gpn/Eo
+lIaOgJkvKQDWNBEhMMzojK0WUufVVzOP4yY23RB9Egw/o4uKxvTUYHKpMWBS1V0
3h70lPxbvUnrFdGmfTEHShPlJi+ajcPRDiwdaqf72shOzPLzxkQNCybGVz01LmEr
5ojfLsNCsAMSVW4ATb0lp/d3b9uoJ97gabl6g+Lk5UDFJ2cXcrK2mqRUOwgdduQD
AlfRwdRYabo4ocqABqyWfmdFWXyhyK/BaCZZbj3R2t4J7bQdRyvtxSlKZxLgs2o8
XLQvdB0H7NsjNsIct3+npJ+nKQObTjyyS9QPztEppp5sxTKpspnUt5ESigEQuyCp
Sb84RCwL648DgTlbMnq0aMTDW3LO+D8OwL9JJlkTwvs1zAzaTp9yvKC/xzvILGaC
VoK8e7boR8bDC8NaxWx3NZeimGHJPy0CaAcDJ5D8uKfECZs9L+g8nfYfEMRgY9r3
rLOya6GDPev5tJzaMbkyH6jRmZkyIjhHWU/ZfK6QT0/9KJADm2NP069lBhe+he35
UPY6mAUMwmZmUdHqGcHycvqLkHYxTjKwoW5Yr25z/twAMahNRUu/+LfrFtJBzEF/
VZPs+5PDYnMrHrzrH+IOh0SxoG9KbbIVIX+H6CHsekg/d+duBqz6NpzrxTdG7/sd
l3XKlD2ZHIppvoVMQRHFJzyE/3cIl98fmNhewxLuRLS+olTQQinq0XNBrGEeesZi
XYkRSIdmF4QeOFfimP34b3DcNL1xicODRSwlQxrKgT29QZKMDwvxLFXzC6I3/Bv3
IdZcqAxJQBTprZ4uHkHKsK9Edh2JRpdQbX4Xj+Jnh73U2mabzWPuKaMSlBT25KxT
IFW6MJmL4OG25JxQ6snsfDpwIGPrQ/TeJASJFGmvOwz4LP0XKkG/NkTYepYXcWSS
1L1miWfL/TUgqDT2knZDH/SRkxY/DBjNvPBhyKL0A43IvIKPwVmLiGKDjn+UWPMW
w2Lv/fm18s4SfsmKefSD8jxDq8rHJGmpMHa2TEGqmAm1kXmoNMsxX3WYqGHphzCH
GGztleIv9jQSqz8UnOzj0mtNqmhGpsfAGWT8aJNEBo7fd0fBYo2QJlZTbR5G5Zlu
3d8eCSrPWZJq/gIg+Lu56R4JA3k9Ny/BL6ImAIHEYRNEioZOY2ZlpnyxtQA/WSZn
iPrHulPELPPx83f09w1yDaJLWd/qlSQaKVD4kh7Ojoo1gzeSsbKLJeUl7AUpRHbf
c5Te5YCR7YrqZV18NnuTqzfxQqJZKw3zo3WSSHfnpiYRoMNjTK1hjo3DFiTFJAre
J2d7cIBa+7bWUW+b4O1VfOUVCBw195H6Dd89ZI/kUVtKQeTqhO2rVaeQCTeHiN92
z4IXbbbho+o3I2DNwup6fzdgMiEyRJyIQHF9crg1UmkRWRtfnCuxgvrCKJ9cAMw2
ybO/Fy1EsMosziO1yJMpfXNxsRbx0BYQEH2UeOF5zF5Fu3kJaSRZ/+bbV7Nf3Wd2
qjORE5u1odER15Sa/HnHEGyBTumA6c9t3nVwdxyfaRcz3CELH+NbpisSnE++xP0M
FjES5sDR6O4TxzohBrcggvvAFZG/QWP/Tgz5xczvR1XJR3rWBuZiR7pdgFxrQ2Od
ux8c2tIr2qvGMYlHUBp7hJP2dbkkhiBCv0rdIVC54eBW7dprcBdNyTnr4dYspdck
ADrrptjahK2S2m/ShQOg+B4iBoAvsbOG+0myy7p+ZY+QXrxgQS6EMGGwCogRywFt
um23jg/sjTsFN94PYUooHG/bReSxvyBAkMxA17HwqK36YoKHXU4yLVoyc4OLsTFs
hkQ1zfC+FyAV7H6NYah1goi++aS1g783iP+AjYN99/v6kChZgrTXiEzyzd1pjujx
MQ8ULYveCTxiJfuDErpM2m1xcpZmLF7sM+pJwyzrKOWUcnGoyfhm/Ei8pXCqHaMn
/UrDg/l/GXTG5KGYhsChKuK8/NNFS8evbcuQMORZ8Eoua/1LCgiOvl9uOew+0IKw
SDJN8ceqkt2fjaTeGR2jpCmXAqsTzIsUOWP625ptdIh0C44YK6y6ZXaZvoyNbwwo
+SJ2LBR7aOdKsLc7QVNnodyiFTewJCanhBsa5FsiX4ONo9rHBrBS06dfGeZKSHA8
u5RUCu4XfzKq1Jgk1hAMHPlSpmi2W0M/8g9nqF6xfCpQGqulrXBvlpEhQXhoPGpR
SRT+6fvoc1si9nUyY/Fjh5j4AUxHQLA1/11yG5QuFWMOpl8zqXyz2qZn7oWpo7iq
IY2DSBTq4fOVcLKSUv3HqBbqq8BVIAgW6LsP8L69qv5Qo7Eo7bjvQY9ntS1E8gx8
vJ2SNomkMMV5p4gKBIeo86RMbpIHKHVKSpGTKU2DhPZM+6kA6z58F5PobpVdOqhM
LJEZPByY9UQ7CUV9Ex/zBTqi6x6FATYKEypX4kOaH/ri9eM6U9i9igOC8qqKr2Pp
IrQMzHZkysRf4kJI7rkzGVnTni1T2cHOrBiex8Hju6dlJEHJkpOrdDjaZspEQaSm
H4aowmaJ7kQRHM06IrXv62fICUzOePHghR1a6aSlbYWbMf1x+bt09Zc8WI2oMOKU
zIDYf/2jWTkQJWLTRnXPDq8zdwYmgiHbBCnFyoxZC8ONQToaxIM7NBgCCeKHxjdZ
onjdMZ6ZUAUHAg2yyNy2rnfFqsCU1vmmnj5DSvH5I7pBt5VJQ6ec+b5n44hxpnNU
aZ992GdwIQ0f9eRht/mtgYrvb/OB4K7up1sYtub6UeMKvVtsctwgQ0o7o7O1zTO6
ImqUjVAeZqRb76wKoH02aeiTYWJ9M/5klVv5Ku2VFnQj1F1yYcz6ct+3Z4hyCPKX
akBzHWWMmpPaMxnA2KSnKvRxrpnI2nMHGoJyvphcMhaN9iMsN8vIHxFKZeEboOUE
GuXkTPUyVnRRLYZqRlH4nEN00tB8cnGyYRhNG811EH3GZzcFVYU2KlBmKS+Gj8N3
Y0WjhKiaVUnEWUiCunHNfMofMaWj8/enupKnOAR3vryyEsjM1vloS3vrTYNM740t
VZjZfkNT4sUOeSzVZAhbLMrPkVQF5pD2W/9kPlTw23zi68Z8GzCYiO9j5WPsQGXM
FT6bQ0BJ9/nblIbjSsjoko7QOS8hMI35PUnSupGhio9pu8mYqx0sRQ1TiX+Nulh/
E9u42FEX68XqwrV2/msZUEPoq5DyPGo3HoxMHog+PwRAhucmXu2e9v5TQHyfaF1r
/oRRU/ZGhWiTdGOt0aeWvJLjOjeoCO/faFGeDai9VJWnZuZMdwTXvuZiJ0f3DTsH
bV0qoGK2QbP7GwUguiTs292NwPXAi9ZI2kdR5wbo6agfJJXvXBliPsbs46lAVAeR
uYTi7yv9ZMZVNGy28QT3c9RF1v62KXXZgZkFgIcpekRV3mGwyEXYMK0mqEiYvVJ+
+bIahN8QOl3BNAOahIVO3Bt/bxA1JDs0usScGF98Sx6vMOWoT1UAE5S6d19J9hBO
9ICbNplJrtxLx4HeezATIJnN/stlMEy/uLjHcFrNAoSqpYlg+TYqV1yDwal5nlg5
ru8Ihv/XQk/Ve1UCvIPqGwdz0HkJqoXTixuLOxVfKvZRIXxkcUqd13fFcrmd34tr
Yd8oGX46YVk9pkr3vLxdRQ0DVNAKnlNyqnHBaKeTMPTQjofoMVy+65tssz4VeQqp
Nc0hqAoHirUF6O4kM55dfXPjaimPe3YAeD0CBok4wv2F6j5S1GjkKqE3oq3T3PV7
+CSV1HxlCJJi5YtkeitgV+Jr57UXUqxAQmbcUG0if5Edd7eVW6GWMpCrERiCw8Yc
BBZ2I13YjS/VLpCuQQ+/cuDNUAsZYibo/1zRiFDxAQ+B8en2rbWzTGvSC5CV8bX4
XhU36Pv5O8WAht8vopcOVEgYOn8UhqgbVekyT6cKV8n7Ly1B08GeDVON9GNIEWnN
PmlZfAAB9GSP64wasDaBraq0L6ItFqM8uoi6QU1oI/paaY5UgKhvcUL7IAsaaaf1
u+xRCj+GqY3kH2giAE74lRl4VfJ/Uaj7cTSXytkgVzo8sm43+rcA3DAWEQMOKitI
tgS434yKGeZ/5uEzATjjB+sn90TTqTG7Nx1umY4LyzVLDVVI34l+GyBcZS/jhefa
ju+hxVeVu97M5TDWzCcPCvkVatYpxxmYSKP3QYkg0TMBziUpZGty831GeJTA5XTa
oHdg0q6/aQsAv8JvSrQ5l6366gf87bfRobaTRpEITR6+8ieWzI3/FhQ0hbE36pmh
LitVZPFk22v0JFvPfIpSi8Cdxq5wUOoVbZeSEhFGeX30gEiRNTbaU+84NdYQltV6
QhDcG5eaFA3Z8HT1MikLEBLAtIe4EICryOUctxeEtmuilF9OEOazNa2lrOXteTFJ
DjHcRTVPj5HtDndA/vQorLu2zAE+5xcbA4xoP9eOYM5QODYhLqKc8rcHhW0FYbWV
0nPXOaHEUqVPBjS9M4cEmOdEy5g7fygnohSUf85kjVtipCR+cJBBmae5fFFOB7Uu
SsKZ4lhI7MUQC4V2OuhaQ5ydpyRmaEhhaE0iocTWQv2LYweS3Sw84EW9bGwAVrJ1
DGGA6bhvfYCosJDVeLt/f6Ift5Y1QNo/WDyI9skQXctox9p0HBDyFBvcMB/k5ojR
29HapJt2FuBjpy3/3s7+VwIJY5uE6v3LC6VMXsTpKqn4WCTvNwfaDcdT1POiyFgT
PeFzTf0px9suU7HRRHH/Yl6ZjeA4xyrKDKJ4TS7vot6+Zk6NInRzjWDy2+vC+OfS
hfF2u1Ak3u13BBwgSzsVKAclP1c/dYKH7nVJQbstyl2Tf/E1HMOuHv9sEvMtfjb3
2vAJpaCB4o8v0QsOFnzT0g/pfMDetEMve7oSZvIPcuDpB9TErzSx0hqmLv9Sz3qM
wVj0oQlxH0oLc6OreflZAoJHPdLDlb+Py+dungpcxeE72SsOC4e5aaK0eszGZxpE
9zbPxKBAOA4Kn5t7ZF4s6LyPeJQAkawrDkqRdFEXEDLPyqicX9gjLyj7ctsYUsAy
KhkMnZDhMugBCV9JFYBTtVwxPid3tZjaaeRmg+cz5XnGruc1KFLeMKeBHWzQi+RK
g4LxFwp6AFcPQVooEAZrdiJ7cpspGXx3sZ5E+FrDk1KKuezKKkJ7Z7PMspt9/Qwy
hPZ+jdj8zwgIn8MK3LnVNzgGrYilLSNBWw6l1YHm3nlvlagYQRgILe73/sM7UCD7
T8GP+38Y6I3Rd+CrmGb+iHqB9w95SC3eTNoOd0g496/xG0WGeeqgBhhZEI/uFCOu
iedKwpP9H1U4L/LvA3fA0OcokAgQpv4vjmIHVYgLwoO5gaD9R2FjFQHqzyzm12pN
ZPyxaffB3+BO7p3s8Mg5FI9+X09l5QSIJ8UAnFWdzrNTATVYTbo3VR9FIiskuskj
6cLxdzCcPYAakNC/KUtjf/+9Iq1I9AFx100V9emqw0B93lDdL6vDUMi6ShwN3AYn
N87jt2uE0NVhi8WDgIcRmH2Zai0Iww+xc0EYEVXEdOj9GU65mt7xVRWtaOaelYbW
+KqMJ2r7TXk7sE4zToTDR4xYi5vRKwp39wbXu/GI+zYXcKSxm5sMC6EZ8v87LELX
2lATtbxodT4tGj58OYV5tHLFLNeSTggDy6/MrwxwV56AE86JU2vq+xgr0OokGNa9
ryfa1+zHzCXvI5XmEzMt2SV2VSklYpkG4W8Db98Sn6f8e6FXB67QUsZl6Rhu65Xz
DrxqHiv82B6R4+w+Hy/r0lkAiKCOLi+DO/yHoWwORqylmMemuU8tcH968NIxwMrI
WKV9KiWhC9i01JJG2gp8EtEXNMDG5cr4tf0817kQsM+3tn3HLxLrMr3uL7iJ6szt
DQCeC8qD5fGmtl6irHMF81MVYJALvUVryh/DkdoSQVCg2vVpri52vmx3cywpORSX
0TUz10iiZhBUHI78BnWcYFktTSMsuOqAN+va8yaCrJWZW+0LlNXttbBh9Bd9OJlo
zw4cF4BpM5iu92qhOeGwG5o8W77pe6m4eK2Utv7aPuLGB3JGuzUyu+/bF1tXkCMt
YYevUvIw29ETtCEIsaVWX7M2aWLrinHpt4nKcgAqzt1qkYkfUHxjaL3JAix3oWb2
bfdIgA8WiGBKNIyRnErhmcEApWzPsi751IKMS9QBCNE+pmD9igJ6xPbTOTi6joDJ
yzd3Z1rJs+QXImvRvVMksYwsHgdWJ3V6VmSmKJeXayx6/dYX36yKj4OdXTruBt9I
KMt3wiofc8zYWkIRJx/zItVf1AYaf7kPkPeXbRkv25OcH1s7dr2KgkENGAlG6Fvu
R2N4Gegm6C4zIrZjSG27X0gOi/ZJwDdIFhLjNo9B11wxfsMQYl67aLF01/uO8Luy
EUyYIu+s0WXZzaswtyE/sBtM6ya6Q8eyOfoOPpeDFQYJPPhP7D6N4MySwHF3L0Os
YmsTEnpJgRQT+wLQAku9veIE/rfjfWYpliQF27dcTtInWwe7NIj9E5kcEnp00kE0
d12ZHSluHwNXnX0cOSHgdTJWJoK69s14CVoQRs983SwhzrLzzAeOEYd1aWjdufQ5
BrnJRKdtHfN1RbtKv3mJJjNkWCEKvGvdi96o7l4e+lq48PBHkOkqPiiXNUE5pZ0g
T2KPIlpeWDZdJet/kVJ6RCIQlQLZehaice4mOh8Vs0XmYqzr5/KpZm4W56RO682o
x/jMsps5mqS4Olqtxo9F/9JHuzmUlGkcD+cqjfABSLq5YXE5aj91wJi82SOpbJow
Ml+I7FnRFaB1WgVlCIq5YpLgLwvbTM9kZHgwtFTeBEDA5RFrlV6qxfUeaHXtDkGv
jBSGCNF3b8mwneRouQi0xxxXj98ShVuGAw3j+ghOFQ10CBaPmwwRevr9sHsUt5PG
avaSfFDMxKqisiQTWbx6r+pULxic/RH+AZoC3Lk9g+2M9BNzGEukfINL7pYJkpsR
lP2NUn4vr4pnXChOO1AR13TCJeqVZ1dG710nbGz8j2+4rO0PMXpp3kkH+BXnXccC
allmnVRuw0UERjzpUFXMwov2YXgnDjRzVHwXU/n7d17HgcfjxO5Qr75c0lhi001k
S4gPni32e8r7SyXnM4u3E214uD0LDXHrlAsiW6dQifwPr90jx+P9cw1CymwUMdVM
NSPCKDyWkJQDzWjR0OzNanBB8VGWjYRT+XH0knx0eisCWknlUUxXfNYi1OvSvVuc
VhuekmtrOVFcVRM+EKgDFwYRXdnoOU5huQD75nifp2WkWhzFp4RqfxFzP8vdEipb
YWChO3HvHQuKeutM84/omOamC2VVaVqUFlU63tC0JT9qoMYh8Qm4j6csjZ/ACugo
g0JQ3uq61ULXv7RxBnzuzqFRKBnl1JndfK1ieCtwmjOdeqx44CaTWmlHueew42wm
/UewZEcjjIuY1JJhqFlwoHHB4nYdLj5Mj8OtobSlBQgX8m1OKVoKkUiw83L0EjNo
F++T6jD7uTua5MO8maSXW/OJYVedVCd5NkZS9aOHPYw++MrkafYkELXm1sVhG2ue
RBwcWvq6qd0jeVGqM9untcoxvL12Hh0siapGXYhXhx7g1mJqIDo8ASJSBT9qLR9W
s+/e8pAQgYEW217aYyIBgKGdnVJ8z7EovjJAfrcUViJFAQ0Ymu30outNpu3BVryZ
ROlAUdssSB/2JLuiyXCoQvV0MVa8FYxotI8KXJ5EUK8lli3MBDCx7Ws+C8II4Y6u
vam62DQUlvWzoXDW94fX0d+O4s0p0fWnCvPYG5zD82hsiaEID/mn4zeliCXC+4vS
7DyfLYvexAN0rVID19cuKPXwPwWunAHd7J+DIX5Pn7JWi+/uvVsWzg3otWz6AYQq
AyV58SB6RNve4X1zdOdxTELh0oynmsKn5bR2vuj1jXxgSvwROM1rnlbLTTf2FRTH
HZdvQOodNAxOuhBX/m8tWmTAgfXcBDc+LGa/KOe5Atyu/vY1MvYnfClSDQhIUTj2
fsQ8KFWXU8TjM9R2+JIGv0BXl9nVT0+D0GyES3b7AfyNC60JtCGOOl4V/Bxhth3k
S7DLdPm80s2UZSl7bIfA+wQq8oX7tKEGcAc/wFq+zhVJeyGEREXSN8O/mFSXOABw
+TZqttgWDh10ul/N3PNa/ory6VUEhBjIY3RY9Zee13HZ7tVRh8Iv1MTXT+5ODR3u
BHHCPl1mViQEEbdaw7SmWnI3ciliRbVIHrPvhtZWwEo4BOeHYAnYYFsndPRtRiBW
64j/RJ5laNbAwma3WqzW6aQ+ZWwwHPWL0kViU/Bo106BB0reWJae5au+/EgEYRJQ
wOathBS+J0LqqL71XxeDXnjVEM9htfizhBXrAjnb/lEkHpErOvrL/7SseH7mplm2
pkqdNtHudpbCGZp54I83x07a/Kf/zZhdg7BfG2KVvHZu6m8JV0AQMOXcGqwf0kDe
qkYi7NNMGiNtuHZHEKkVF9oDocviL5IyVAtuHjUM9z6teA7fT6q3Z42nwuN/CSCE
lsVF6PVzQWLTrVGOGnimlUkZo0se4uhjXCNlOERlWKJl/dGyDw+em3D2XGjMd1SZ
k/io6MSXbdBAaiLQdpfJHOW5+NIk6WaTrl0k4eXsiDuYjv3aVm7w6PpmosyKwdph
1/9wS8k1d+1IxY2G41NQCSY8WOtiHfksexN0x7EC3IWfMpBdctx04nWntuNHImg5
EQqIEykKnoLeKQ/RhDc2IM08xWP5Dmvhr/ly2te7t1r7VQ6xOSvnvUo9uEJtl+B/
5UC5HOyTW34P3JHOvuHIUeaQcYB5RGtW+wySZ60kYjOSURnB0L5LKLnaQhOt1Jx+
taf6Miz2YF9USL2/oZmrAAed6LB7XI4T5KJYOluMiv7q8ch6HBhJXZEfhz5R0O6s
fClT7PtbZsu1ncjvrUaQlEyBm9Udxr1ahbE3CJNgqZtpfiTKJljV02Xbmx5055v3
CyaVeRyL7VOUDvffbqF+v0XIeQT0H4mtqEUVk2nzUcJSXR0G4sQ7kO5XKQZNqPNS
ceCMVe89AocUSw5d6OFfjFDenw5MxSAgCK4SlAjHkczxPFMYoYDajucHmB6TYr2C
QaqeKsHkDyv57CfwKDgCKNFICDNRzT1sBQl/ttRb8zbg0IF3X5cuu5WldwOgmdAQ
OkhSonulf/VKWzRfLxDAjt+Fv5vGZDpDpfcPmcBa+wQ+QvqvnPh2coCEvhLUHIkT
Vur4/8UD2oCHPH9VQU8P6zLwmWY5F6PtAoAwSrz2V7PFvrCTI+LozHmK6UERdjbt
nIyHI8YFsT4n5zHC3xHj0LvF7fE8szvNfbrx6B6E4I86iwYQKaatNr0+iOVb0MQH
5Fef4ow+/80XmCZl4t6v+5FgVUdzFafFqa9KGrstlj9xYlSUOfkzIU63LeH5FHue
qMmAKsklOirolBF3kd9dW91sTeGySwsYO5iapeiH4UpL5MTA3EvFMAIlj+C7FpdG
Rn+Rrff8pb98mMzqBJIsEAXwxekgoiK0LJ4xGSSW7F4paZiv8YqT4z89EchcsK77
aUYTUIfYYjnd080dpEPU9et8OdTJ6K5ia7nVbcQp4beY0/SqAIQpZgqvIRBlk/Gp
PHNzUo64mFkJC8s8xjkyT63/E+GUT2F7sWtYIXl56tNWmKdzX1mkN47FLPvVCiOs
2SkHEGphKfDAbzSrIe13GS1klRcEuepHC66CHbXSJ+pwWuUYmkDlMTypQ/NqCgyG
2q/hI3XAalILiAwnG0lLXnIinLN3o8z395KBAYy3/OqMYCE9BAssTBT94EDJaVq2
hxEaWPluL+TY2e+H5zBahMnJKuJqoPQ24smKlSFgkRtKoqhmkvOtO1qxQ44mgpfX
/4lBTMSpQZSOOwQZGUsrRLJx7xH/nrVUV+8ohFUW5WHIfAmxsolZCvj8lHbHAta8
dDBkhPukRJYLZ9hc/1XV3CJ+Yz4YpWk9KvXwbLkzELez4pGZ4dI4KO8RkqCVcFRn
Efn72gTO4qHPZrNRBdeG7E/EYEj/iz5B1Qxp4l8dR5XjWJhHz9+b0niUhne45ERE
LHzUmWvu0xntPVosZe14m55ilc8KMdSC1rXtgc5M9JautN9IO5W9p1cxwxovR/aZ
TM5Aofejn4BpLfYOOXzOpowhEJ9zQmp94lErHMxZzbgqGpKiI6lfi1A41ob5G3Cm
fW4NXZOoNuBmS8yvQsNRwABm/YMT9v/NxmcKvYfZT3iZ0gdZ/jeqCQlQHlvuRKpY
6eDFTM2UCJOyaJkh52T0DSAU84aUtUxGXPHOHvbnKlMkeZkhEEOkAUrJhl2VCUnt
LOTzfIOYRHLEZ18BWMc2h+6aynqoqplwqdG7QCBGZnQjHl38UPGztmxbtsZMcUAM
MfLGXsvysyJG9kuFBtkr4LpdocZhu+SGf8xe9yjKzKUj/RBOGOIPSCNvuFFw7IoI
B2xW/Jfy9bBnrYXygBsfpF5J4/rYiirz4RNI3ln6NE0R3TTfVnuN23DEW2RlD42K
BankiPDMaUwibMIVKcRQtgeN7ARx/09guwaU/4KRLCf4bF90JSwX7NOqeMDy3xDP
jIUP1qHpIjHyM+ipsIHRBeapITfmXdo47gJHZaX4fnN8nlpl2ckA5sni4sbv+IeF
mDs26ytlEbDo5EyDGL3lqSeG5vlE5QhwD+tCY6pUMfuP7iL4MZ0rS5f5GRQVfoPv
nR7UmUvvfamRIWzphXk098AmKn5TZS4oN1Tr23L7nj1kGc3TQyT7VKZ2IuLSOBSt
wKJATBAQEJb+/NtuiEjNDYqr8xuxJf2HiMM4z6XyXyPv2n708Rwvvi5aqh3xc8Vq
zgMM9ghggHOrhSDYtmhxqKiysQKd3yaPdlJmWGPDQh/RV3SHqQLuv05WO3qSxXSG
9q5UEx2eVvT7VGT/T82H8kufet6GrAttMr2W5PjuSbRVTtw7DJObByBabE3dGgS/
kx5wJ2mjI+/CHZ1Fkcir0aMN8Wxf8xR3vwOmvP8zzb13gV5w5zY2Jsv0dkNg0Dg0
Zpz0P4UUYxPY4dkwofKYigc3CqjimBTgxuOpvGDyevZnhiCTxeqWaJtIOHm+6qw0
Ug/pydK3fgstD58hUIEeKuLuRd6Xleugbmc88Wfh5y9SG8ruVLEqGsm9Tv443ALy
jav+vt85Gjq2bh+z4r8fEBggO+1FYdOJ7OVL6H2APDhpYvL4k9BMeZqyoTmFQNq+
p1pb3dtO6tOlIEoPHQ4mzfDbuc3TFuX9qiIcdgp2zWa2CvArcKzVuc3OKICtvw/7
XVB5CduOeLfrG0b9I5+V0C19XJ6an3TZTm1WWAxw2/WCsNGffxe/fZ6E1JVt4PsE
02y+SZhobLjzonqRyCvRVcGsCb9j+N4faVq9vRs4X/bKvZG3g3GjwO4csK4iOaRF
nsakUmgqYvZN1u0vUq2a8MUwzTH4TBuuJJiDuIHPs8osgCUH+A8RzqhYX+PmEVOr
cF6vvMeINVArB5ZXBOPWSp2tD3PhrDqWfQulNPMu3zGV/jJ4OuVOeraIOSFqwdpE
D6gIm35/d6ZaMaoXwrtIYL9IMTHfuLbhuCU+sDs3iqPHoywE9Vfya3FpwbFPWrFy
yNUV4bDByrZH2vfHvKqJ2cwT+ftObdLCPHntzNSN4nUWrxVM8yXEFz7ICQn4sTRl
9CVbQO3wcDoT+/08D6lzLCT9XXSynbqG4SMluWU0mYYaffdv6leCJHy2GoCVZLIQ
NKNPdoOz7LlqhgZf8tde2DlqMGpfiU/5pijkD3wS//Scg7sPE0i6XSHRnamvnRlH
yOySVJlY6DhZych72Z14P64kixzV+keLHZvvqlL20Npmgdsh2/h9iwmseG7vFmMF
HQsjM+nYKP2oI3aVbVvEKKqpWe3HyeGmaYanzibQZoAxrL5Ti9IcymwWU5uFWMU0
SdHFs0cBtsg4zkluAzRJpm/g1rAICSjTb9usvrkLP4NWpqKn/5PAZerWBm1C5ImD
YUgNaVU7ozQnqh+Qw3diOp4FMdMBvRPWpH3nzjb9V50iTTvXmPTVuKjLPRi1ql11
P92Of3K4P7vX3QEOKbj3hgtLJOAVyM6C49JmtkTMbSM6SYA66Hs1HzfCQWDNU2Gh
8yP/a91hn8Guu1ieSvAtGLWDoXhcZ3uL1VnhBuhi+Ra9EZtwRywAG1JV0hY/35Gx
MrmuawCydA5DlkysXZyCP7mI+3vfQ3FOsfw1H6llrdKMyiKlE7o6fl4XydQCRRJZ
QoFd0YgNtEJA1RObodoFLuoVk92rMpFDbyuk6DipZMrzjopeL9z1ATkXD1NAe8wv
wBxAs+RCGJtIxmwheQp/mdURaekdhJDTDZ/6+z13EFnpJxNT6S8HEdT3PCbm8Qkh
7i8AfrcxaitrEsZ0f9lh1ZneLLNbbYW38BDW6FVu4xlj7i9GdpHqqoaeER66rp/M
Tocjk1bQ3/tBql/Ry9WYgThrlzUWUHnkTxp8IgMrcvtmdGIteJ6lpW0GyLKHRXbl
/PtocTb4YU5+DkadC0XWHM4HskgIhTG4Ku0GcMd5uP7zusuQkKs35qmnOykSPEwK
SVTM0cQfR7ctzHBqHMCyhe7b3Aa7ihWbv/5Xx2I4HuEGSJd8erGO1u9wpdKaLOQT
6wo5s3M2KllGIPIc39qDXW+EDTwSrTT+5HrhhV/zeTlGq8VVsG5gmw5912d+Do5/
ImcxiTpGDEPTd2eOmvdiQRI69/d7b0lW7k92YdJ5Ps4rg1dLYkMHbbI2T4yy5I2I
Y7ZLIleT7Y2DG+m/dQ83SBe9VEHHo/jVH1SGZJqAFyYWg19+me6Ih14V+Woi3TzM
C/7mXzoCfundtbwsMjksU3G/zunIouxdwqaCosrfCyP3cWUCZGDWMfkeRlwDeI5R
nbNINHF9170HKq2m+Xs0yGQ1ihI3diKrIZCw08F89FYEO2pxAz6feAV4CQAQ/Ks5
tD49VubOtTszfPXygGjBJGVV+j7kDGhDvKgOu7L2Gn4By/EuLF1m615G0Q6Rv70P
i0wbItDQHq677eTog1QYsV5LQGqS8cjdaSLLC2iSzyEPIW2hjb2DxcT00Ho4k4hv
WQLHsXf/gt1st6Gd/BG2lGEYDfHd8F8n/LLL7JTZw5p+ewMDPydqj9PlhVNo2+SN
kkdYVC12DR0t7GpkC2Qu4rgZRA+qrBBoMXbb3cCP78hfoeV8CGeZYLmzFow3oLZx
rsheV/6y/FVQFXEJNGrTZg==
`pragma protect end_protected
