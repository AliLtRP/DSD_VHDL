// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:39:04 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
FRsSKMPw7v61iOSqhjtGKVMFUPkZBvbvquiqU1m857g834EQjx0LteR+6lNfAv0J
tsgRA6CXOO+Lq5h3Ukhdl1VgjXy9FK7JPEe60U/SKT1vW8os64Hnxk8d5gJlDKCS
uaHLeCjgSoznVP9OFOPpB0o6N04cpClcIjJoMcURtgA=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 38432)
90v7WNfjuwuqo8Qg7xJdQD4ZOXVofv/F58YFO3EOlZwfmHlAhD/coGbJRGg4OHkW
OBulI0IqWvTjdmcebRG+QoH49ZW84yC+ZNHaJi6whA+Foac/L4Si00mbhrV1/Im7
BzPZWmeCHDlx2CowGPy5Y2wVm3z6vLUmycM1Bin268sAf5XQOWxlbRhVZyx6wo13
1q5DDQcqVhiP1bnbNcDcaK2PTW72fpIJzzKvHq6ucJJUdOy/E8Mf6AxizFAc8Wsl
8qVhcWLEnWKaiJ/Oc+rMcHsKYeqGRoxZN7foLEJvbW8Gv+P2nbK1zG7AfFKHSUjK
pBG/Dw29ZDllH+6Xl+DCmY8TuMHLYqRF15eXFp67h5Wiie2bZ5/oouj/4g9h/yfT
09IruF/taRCToHKXRn/g/2iTrQfXp6wB4wLK+8c4W/5ml0rFlKYJC7q0eyiAjEIQ
fCCts2wDVZhVC+Q+uvqlY8q7rVB8w3bSByhWc02XRHVihjMVB7ZZTVxC0uEO2C2p
4yfSJc0I+R2BKSWzaA1O/lZjcmH43zW4j4ThkkDJw5IoC3g2xgZFqWghB2lEdEed
yNZ60Ybbbba1ge7poywDKKDFJHyLGL7rI2J6Nx4ly4xYKdleL8BV0f8EsPXEUSPb
kBKYKA1nbMKaspeu+WtqsBSIP9Qmx3TCtVlQKrLwH1uE2pORAdqkYJcR47lWnJDV
C44Hx9b0cbyaZA9FmTrv8aZM7sRkXt7lzypOcr1QArYzkujK0fJAYPX2r0HoduIu
rvbyWU2xSsU1mqdk2Hyige/mjapd+wGK2vKDEVaWqXfn50WyYlPTceXOPojoquky
ZoYRXo/8RkSLQV/bBR9TKw5H6La5WU7lexTvWQTp82i200Paa3vd06NTU0vrX6cq
p18IjzvBJrAtOaI0NkBw3RjYd9yK284habwPa2pXXWp2othgBJUUYRbLA7CWEiL0
pgvDMT0yeoqkzxDSPFyu8LbthoOe5yY2u2ZB11FbzFO4QpOiNoEJcXKyY/vIkL1u
SDeZDq0cHIJxnWXtjcl4R4JBgkouJZZmV8bc+nH67RD5e0klVi/ohXEBgtIIjpsm
DTGsMRL431+RwAAc3oX2XvfKh6KY+NzMUK/VM2JrVH0ZN7aX5uPasoxBFGQondOq
BLWqjQQTeV7HPvjPh6AgJiQl/MS5+Wz22LnvvRLz35Vtt1922OZebFFZWU5CMs26
dbVeCBPZvDt5QQnAJJx07NfbcPLdcgFMG6pWMyQMi726ziaxukI/TEPdcORDhAI/
ToOi5mY2VGnNjRHPozuyz/wt+QrXmhrrt53if1x2UbidPugpSoR1DFRzUvZoGrM2
hViLF9bOcN5pek5y9Q4OddrlMU+A3xrNnaJh8iq5pjtu8Mj6YftM82wfU04dY1M6
tlL46hv4ebJSBrXfCEZuwOgACv1s9Rv+y9IATtRiHFTeFS7ibLzkYJg7pkDFU4f1
jvynoGEiKf0FufhjwMMgXYjuCH+lvgJsmu1Symi5gKLGZCbJedS/aOCMb9Wnl7Ar
pLzpf8Xy9WgGxzAqlt/EElYwD8o5c6aNr68UCTXx0e+JafYjWgoMlY1e1hZCq78X
M4rp8Jxtial+vC3kycHr37JEBUvbdVJaoGYFmXhF9YQD85F2rjh7+3S83rpwPNvM
+NmbIv1iWOK2ud7ZO0eXPXmd9NBHkxHAhcq9QZ6PYTzWHqqNO1b9SdsjOhuEl15p
LdaBNjaqfryfMliC5mdFG+DR6NkB8Dzb40A08yU5gw/S7QhrrMCFEzYrrXeCfF2m
COXl6mbr9LW2bKt2sqV1f4pLYvNz/eSRweq56sKLnvbCAZUmO8sPKAx5dnuO40z1
YQ9DFmSmbovT1hsVK79AVw8Jz4hKm4msH9xXMuS62E45gLRruoXmbCgiyC3j4ilz
UEIYff5DAFp8r3n1MWO/BKbZEuxpouUPh92FsUxVCVwXL7nJwGr0Qz4LxpNgyaWP
/qxUo/l/Vv419W9iInH7DIyvSEdTEz0S6Nam73lA2W8fBKA5kHNFK2zqdVUcZSeo
0EIJHRo9auh6FedZ+F1eqsH+Nr3hMePH4cO5oSDIEx48nQ4c9logZdrvD/y5YTwS
i22Eeli8Wc0Kyn4JUADs4LzQfmM+imQYbK61sxHz7lRhzh/lASRW/fQWgX1fTpwz
n8sXkSy3XKgobveMJKpgjO7JMVi9YJZfxNlIRIcb3n/Dj9LSlRUi8HRfx9fY0lK8
Bh7vdD9Z3ncwu+2q1Gb79vT3cTN4qYJU8Wuezktoav68GUqDJXaDOaxPWfcdw5vX
6XiwpL7wBurddNxellwEWU3aQO9agepn53VWOqTQc2bMyWBk3uBD3sdmvNGPkJOG
QXSrNR1FZRTo8Y/8qkSKsecHWAEffJ9xaBRQAsZHzDyQMfE2vtef5A1bfB6rHs7f
2cU5XesKka55IGnXGGjNqPA6ZNz051X2edmqhXfizFN+O/v5YIB7cJMpypsAP0F0
4qyZMSlI2yzJXQmDsaTNSFhFpb6i/I9M40Gdmy74dlroCzwAoIm2l7JkfYPsbVuu
4TdniWy+ipB5KR1ymP1r/Yr3vdGvImFAy+UwtIP0u1DCIScs3YnPEyYnQQDEKFbD
xKrmaR4TQuc+iHsjQCVowuEirjDLQVs1Ig2TucNlVzWo+ei/Qxm3qBrqBE097G85
QfimpQMBdPAuoBM4wUbsq6DtOo3WBrqps+MnBzDH1yEMfCBOR2NvQr/5NSTmclfe
482nTYtHaEKDsqAJJYFUpaBPyEb1bgIbCd8pGIBnEeXQ7Y4s+dJiGTE+jjg1ZXz0
chH2+aN1O09upkAChMe/PiQgXd8BMhNtCQFaUlmp4SfhrDewt0QKddGHMo8UZL2y
vNyvYx5SSLrFCGVfS0aHoqiFVShayWA+Ej91v0cQJ3LohZhWx5ES+gpWnUxYSKUb
kqyPkufDSXtimz40IOC37V5i2eSuIfKwukEvOzLczpEPFpEpvjlMiUzSo1cyuPIN
egWYsmOOSPu1H/+5N+HXFfnUoAEV7Bd6L2UtjIIW6sWUBmFJaRc4Yl/4kZDrVEin
PDvAL4WExmxSXemUKpw9NfDOa6fumzwGxDS4LVfIMRZbzSa/T6A3bKWNdvVut2C3
q67B+G/bTBqR5LKWp1Hq6Kwd6jsErspjhjrQCEJnLFeyJzacdGD9iT2lrTOdBA5i
DRMpBam8jYyA0ycTzHVwx7IWDO8G3uiN7eu++TW0+BUqUWf9XzITXHF1jFUEhJqM
UH1SgBjQmLMlMVzR3CrHFcMl0g0D6bRaYKRvsVf5VevqflAfSf/MGudhPBS7vQhi
ijq9rtFAsgjKCa0TRABa6B/oEbkMeUxblTW4hFM/ZatgZ26jdyu74/qXl0fk+7Xn
D0RqQc7cvDEYeoCKwFixBgI1x/DTCX295s59X24r6WmALldXdtdXsiaaYiASxUkv
49c1AZ/8oAW6RtagyaGX/Ik73Gyil6Rb00yswAm3aZTAuYbGsegpNzzq1adhci3S
1tZEww3QyySaGFiRY+Y1St/iJomEm2RTKjHejzBnlgL+uUmiT1bTSEPcF9g32qLD
CBQA4FJJtkhbVQZNeT4lM1U01wyfoP/HWdZxChUKT0q6ZXgs43rNF6RljMIQLxD4
IhDJ470oAotK1KOxSgeMof4m8wpVwuN6Bbf9+Krj+PqYf8lvv3dmZPZIqEvR11eT
vlwScVlJ1b0vQAx4aqQL7sFN/xRQyzjrDDUBi7jd79rmmk7/Pfr3Bz1F93L8BysG
27bdxuCvbhOXsbyylYLwI/BwbwTEv3zZwOED02pKSHEgj7ya2wGDKEDe8jBe5ypY
xJLH4Y19QceyA614logWyySxlkBHPRnCna3HgG+rPXpTMg36WsttmlnHf9QPvI26
L/MqJAQtOYR8Bja6nh9ZZBHSZPGKYZGi1bUiZcQCzVkDK62rc4RUrSirweKmfoOB
TbBYbdWEB3unTRxnLXdwZdlQSkNfcu1Ikh4caj0MWivbNxequVeynjjhkyUm6axz
4FTzYPOKRAohVG8KWURDdpTc3C4vf6TUxicNvYylZVdA81Kf5ZnlS8EON6kte64/
jD9NO/nMck9Qy9myp4nvOS/Oj6kgGkMWspM2yGfuA6Ubmvm07WMy3RkIzLnH1n1f
Scgf6lwz/f+SGEdVllFCRJJ1k//xVcTsjeyV9ve8glkooigsZxSRwOpBwpAdIyhS
hLGaMruIACvDjanWPvrJP5MHsu7x1IAfkoSWY7MAo1FSwd1YrV9HGFbmfIwHWUUX
y/UkUomZhkaAojqCecOYuSaUG7D0UzOrW9goFCAizN7UJcBepGtl/cwCG3amglYG
fqV4Jn7JpfW5ODh+mRQ7pghVlmlcabu95I8tWPgGX6UqhXKDp0whhGQkYQLVWctL
eFUI+ZOta17k/HAWzhyK2rHz6sMSzC9RfvhlOYQI6jxibzg9M2ViIaQ9STda0ooG
/Ds1iC/FX9T/1hIVzKliHhFoDonOvB4Sd8ad+39QugGVg1u0M3tjv6ZLDhOdHBaM
qCwKV9ekvtWLZzJz2VK64cN9us83upIry9t2JMaf678QJ+ea1FHumPqtzVJvtsNk
QSYVdm9PwbSMCuru4jH9uSBCMgeoIgO7fZZMyOBckVHHK2EY40ynYlKgofsWEA9k
Q2gmulWbiojg6UC2CSTJRQVACUumCuUSPUtHngYk8M694L9KWLuKev1+SLCbpnn/
mUD5c89e/pUreIkOT1u1IouiYsSPQClcXH7fCnYkEQGHv4iRVs7ZrP5pltkY3e3s
DEhkQA2/2vrmTOTenQ1lOMouySa0RaKf0Y6glXmaXZ+k0ZhyrXVmfsNHg1XPYw74
nhcigLFbbHq4beIAF9K0VLmJ7mO6rnsZO6SgnijQh+4shqH1lyMGnbdY2t5+tJFy
TA1BFEcchd757tcQNPP2ZQE1efiv8WOtSTIXvkvFCPmDP90UIV2d+aggZUJJADAV
Ggd+RWIZAI7ibvT+wxzaJxaO1weKYS9WIiWvIDe8akfacC1GshMFKQr7Ybq2pX8r
a7lzDbdGUqBbumHejYuCAEX2u4t7DO56cNMM0NKpAxmbAqH72RXHMIjPfTF2Yz1f
TRZhRx6gsttuSXGx9N/HrvKCRhsTQP9bHCUcERf5nt0aUZx0WOnhtNEs+wvA58hh
K9ovGAWBzBnX/ApKH9aTCGpB69k2xY+7/lncHRS7L2mXJB61QyqvstjcEkye5yBz
XvAo7OGLLbVdp1ybRstJ5w2xH5CM/xm7k2VGS0E4MWgcuQO18gYntYTRW7pfNvg9
a9sq48NfDgeNQWT9cV0wmtbVORRg8W2WqiTbztAzbq/NcefZyKZBuE/z4tvv88MB
Pgikk2xEgTH+ANIza/Sb5pH9iOOGrnggOxY3+5Gqv2oopaJAZWUxn5TvJSbXxmX5
ic8hqUM8biAx6VWUrEEsHMPmKa4azPo+ePEd2ob4FN0C0X0AiZ+2m3Nf+bL5Ws9I
6A3lDYO3Y8swpWrT21S4X6ZJ5EtMtH2E8zwGwZHmT424ZmXB0vNn/aylTYIZKcLk
gvOg9Xv2nj7IODMNkRn8cDDWcCmG7qOYu4a38+NHjGXN2zffIo6uDhK8OwhP5H9u
vKycaWn1vWjWA9+W5tKhKXtAd8EjoLakzaHHLFyJaARBpOfyb53Osl7hk+KX0xko
3m/ZdQ/HUisW/GoFPYBmEGEGYpst1UVzO4oIMHmi4HBiN41DJ4gkLRPQ1+5dQiQU
ASZ7vHe0+GAIKR/jK5cmn+XROOmBVHi31rPctDYtTYuGEa6pMsTNJs+tVQ/C+Sje
XOyhRIKqnFBJH4QUWwrLLR3FOJ4/sOIKzh425h1Waes2iUvffo42Jq6YI4KNH37o
IYS7KCGMl5zCr++faZalHXMy3RmC1i6GB/dQbjQUB+AfGRX4PbJF++3E90G9dRrn
WnGNfGhNdvBmtS2YExEGlbYuY4KZ8MRWkCmkbDHGEyb7Nf2WYZWMBw4bMlK4kgfl
RkG9gpX71UD2S9bgCPjWLVE5CrC5MJnQLOKdhVlgQiemRcAwHf2sXa3r0tJRfXQN
28Rzpp7AiUt6JPcrJs2LCbFnpOMXttDaPyNGeMobbfV3nqfge2Oy+ElrOqkyV1Ja
3avtiZ6+bveg8Wj3Z6TojihdicbHyG9Vd5tDjZAlPtoUf7p89RcpS9grFw/9EWcU
CaNG5aRkqS8ByxEfyPdLWHJSaxVI/WvNutt5ymPUyKoOdVB+wgr24YlfwTqYg7XU
kbxTs/VsyOzIYYNP7fJ5SmpSOfq3ANeIE/hkn44xcQkOQfzXMiIHwS/LJ1ZREpHY
rn+V9HZjAu80jsMED28xbcmsp4cwv2tf7weQOtGodmrd1FsOgkU6294OD8FxABdW
TnGNc/oPH1e0DR2Ea9+010P8H+WjYmcqy/ny/Bqyw+UOAsuLttQU9cJ87y44a3JI
OjqYZZLRKY6ijZaCGGLsA86iOAvgbRLcbuuyZ2E3BAKNwwMN9xBHexZEDZdW7348
NY65dMPKf/RFWaWjHZXlkQT06wW8/lwXBJXewEQ+h4PLttrPoa6v6Gm/kHH7hK8d
azfB2BzAamA7WpJrUCTkTZw/BgIPTJg7yiNwfwKo8kHktuO7SLFWwDFEQWoxT9sn
KTEH1UwweC24rPbQheS4r4BYtHJ7Dz6b1PgguKo/lGMteK5SQUNq/yntzhWqmeru
znpV+UteCHu09sxZMeISf7bgvusdTIlMTdKf2Yqw/e+R5P6K+BKLYfrHgH/tovcr
ng2U5wI8PhGf0AKqeYp2ZKOFEpQRc+bUxb++uPtNOX8BvTqLyq54zdFLrUTII2rg
qYgOjBZeFy9KyPJs8BpZrI6fLxLyZNlsVtxMhZ2NfsjMMrZer6IzsxkIt1/aPvZT
8gZZWQFHXbAhFDVnU9SUJU4GXeR8FYFDG4MHGUZg+oEfjHArmUn92NCWHOCyEii6
aBSqDjmTpji7tnqzlVVb1kqQvSbI0PJ+Rw7yTpY2nUy1gupRsiyLzcNox8JrMrT3
j3dI9HZ0Iwii4Z96W5b4ShRPDloGb9juYOygKp2/uJzu00J9oXARy6tiNQOcExDi
htk5IOu7skSZqfVYT4o5gHdD2xmY4UEPa8kdU2AgQ6h6b2qbe6RXcnrVJ5HcP2w1
Iy1A8jQxtpFUDGDQ2z2ES1TPfDUndZ2ccEOo1MKrqLn2050k+M3hhBg+8BVvFBIE
gii471gjUdevhyVSmADpbCptubU7P9M+TkLtzEXl8knwYWrhjgMcu0Xawu1O2I6c
v/LG+M0qrZ3T/N/xU3oQEUWa8/FrDaG8ZN9sMmZM+T5xCHmysWczgReR4cdlJETw
L30wnTt4HXnClz26H9WZuZnHF7cDHGkrfwrpe9KOcMh4Du9vNaYAxhbEEN8hPk9o
uZx7YGKkC5zWbnYqd3D9Kl+jnfj2B2N64AkM4PR8YfRitYg5ZaAWCfonMHMqBFQH
ovNUcmjyohfLkWOwquShU+yGr/dPWa9Oibl5rp5cnMQOYqdUFTTkYOQqJp3GiNnX
8v4ntEhXvk7m3pS0BSCF4V555UFSuEDXI9cfsR9Q4xrJe/p8e9VUb93djSAdq0Zq
7cSoSez9iWpCLj4i7YQPETU5vO7WVSYmv/l4W4Rc8+f/yHkRLbe5brBgYiqZ/j7e
tiYJnyeKIXNBQddtVRiDcdObgXIAlzYSWRYRrJCJK+3LNDmwMendYqxcUf7zIgBO
J6wHBi7J9tD16UTw1/nnSNkL7SQNzJugTj9thXWh4wyJ7Uewlz3yCq5z8L0emTwb
er1NJ5YFOeL5LXb+Vhi7q//ISLimC4cO16dOzz2JNeVY3EHCqXWMZ8h3nf+R6byb
G+a3Fzq+aA5qJ6lVlQNVQy30aBGqo3/4aVVKPGABP4mCmzqi4+8jjx+22aZ6DBnB
d+Mnzk8oN2K2/QWLAmkqhbKn/1xKVfJUy1SwsksqTcBGwoFKjx8jnhMubIEzmIO8
N0wSZQYWqSWs4o+zh+2cAdvju9Fm0ViI2YkM4CYJ7XJyyEM+hZrhiIHAfd/8M/Mj
dLaRNeO4KD3M1FGa54DwNHb/fwCbgEuJZcUnpUVXjOtT50CsdnAEaTZ1InGw+YpO
NdS7HSEueE1vLmaXidegjXAFdeD3fV6PriNM13vDCAHaeYtaFYsdAu+3nsKH91u3
4urA2pTvVXydEnLtJlLXBWFOPWPL3+vm5oh9vSTzccgHjHIXE703oTn9eOHe48ld
1H3b9UeFWz1/mcpX2ryHYxFvcFNlZW4bpgMY2g4PGK0xi2GfJ0lc2lJDDhbBtGmf
3h+QpumUXAxm6VE1FXcp15ZMdNJDuqgGWdXT/gqxxDPwfphcPslims6uHgPlzyQn
slcwkHUWyFSupke4goiRhSzSpXHDjAy0Z3t5jhoL5J96dFg6KkB67n68xfS4P4cY
Vxg98BuqIBq6wuF6I7n4P6ORu8/cA5vTq4LKk3ljxuQN78FCOhZsJf2pD+VoeG0a
Lax3tia/cVBEQR+hIX3D6bZjTw9HCjvoUXc0JNHQv1JnW5KgYpr5iDEVuLNggLsi
bZdrK5TzLO+0XtcKmPfFeNd/MpWC5Lrs4ivsytpAsC4AcdC7QX9B6z+zylKVQOFm
0lICq6feUCxm3Suz79+CYiXqllZcmo55ugj6N9KT9JYQDkjWYf+oc6ysJTfDwHeC
qMLEY5veLX8z7SnpZgxwvqqBat2pHjhqxWsJgvxR9r9RSNSr4z/Nzt3B8EMDeCft
TQjvG/B9QQoD33dRzBiYTrElxIXpWt5awVC54e41nCN+mCmFkdkvyHYSIF4h6WQy
QveRkDhBlH+Cv/H1y0VLu/nAL7mlInfsEUZpIBJZBjKYf7PTr/WohjF8NzAeASco
JnDJZ3czo87SoW5rLYRw0dmBqS7df/N6l2qKgBdn9d99xmc638xPELiLhNdYIzW+
5V8RGovzz2QY5Ov85Q0p5ZOzFyR0LlLRhLshksk08VxrDNc1IwXLfDRJJ/CA3y1M
HvT5d++lr8jgwgnyBKGgd3TU9VPp4JWC9HvZqh9/xvp2uJGd8PEir/By/Ta1W9LD
1ck0S4OPw6/IZyA3kV3QySZ0vAohS9xeew1nnEajn77XiuHzBy1Ln9Rwq7JCRC4B
nWfaz8zUHcTXnusPG/fCTXpTW+pE70xHw9ctUS9G/aghP1E5250JwVYRknWmi6R5
cVrfuFBkQaDdfxnYwvktwDvZzqEQtOwdGdmy37cJVp94WNOxqI7gh/OgrEeECnki
hDeoaIadGMmdkQIrIdaURqqqe16htdTfHTFkAODSpSDafJ4wwODb4fLJ9Uu+kG7R
J/2nMbJwGbMqN0DE8GHo1hC93UsT1flXlDBjl49+ebE8LjVymVZ2EbVQoCphlkRL
yupV0Y/laG0RhfXMIkEzj/yPzqFdAP38eo9ImEQ9YGSl+B8LNcp8nFomBdjxmlaI
FNKDbznEqfekRoGmcXVaFo+jVSFHZEN7fdT4F5dtY1E6XPlgtLUg1+amG5OdrXhh
7EYgLxMSfb/s6B/67pUZVPQBkojhdPI0qt9rByNnGewR4kHh4f33/mcoE9yrGG6k
IYQht1R3jqZe9K6JvpOTlecw+L0IuCuiJd8xWoEVHBvdkHDGECj5cnE7EL7j7dB7
tGvUZITB6kUukHo6dHQikHM3vWq5Kfq9vvNqet6rNWebU8OLfM7okInNJYsdcs+R
RcdcHRoXRwpcsCPfoNCVlmrUgXlhD6W4v9sYnpNz7YJv0kkUIBhquwpIPgDrRINJ
kwNejJP4/eHsrYVhYLzlC4lsgA/NxHI2184pJ6FkdPQxCAeYnc+VDKcMEIicjP2F
CsRYYgvlTRSAk1ht/eak0r575yV3vblFHIZ9KEtiOUFQMaNxtxv2/OuUX6VLcZMD
a5WCEDkdM+fvIenx1EyrO52Gf4+X5wQq6mS7gEc38Fdfaz7ODsR7Fk2mdahMNWCD
JG0lv1nw/Hv0pOiabL6N4Bvpk6/E/hZyG50R83TwKbXHNde6DDWpQe5mrhClzt5E
/1ddqc5+tlTxcAvbSHjAmWCPsxkxgCbr5sp6S6tr7nvlR7zRoJnolHFlhvdBpYbd
XeScsL+JZs4wcPA5Nogi+JScdggtHBTke1f3m2zp4EcX36/jTKYEDCmGpT0I5hwU
exgC2k/qLstNXwKzWozwuUQfxadMQQ8fT4/ZbTNHcJFlkbTBHKb+WEJztsDSIBzo
C5WLqbeJoL2pvKLxP48HK+ePyhcH3qLPNc6LEyfzhN0oNEzF2d22fEPcQY8tzsMn
A1nEKdgSLnqwPjunP4eGyLXLOeWkm9R03GeX3GwjvlPJXkXr9bMlGJos3p9xkcgK
eiEHzcCJS38tF+7KjYh0NBBEKJpoOhAWBtWYGbtmsoxTKohQ1UrsafmtGmmPgF8p
7JzL5CP/9wtvZBi77tNVmW3JziQbQn+x8zX1HBxFI84Nd9boyXLKGA3HMgDVdMzs
dKfP/cMNOKnwIr5yOUCDXu08VDU8s+zhUoBGcsZriOB7+V7ncEoE0kNOYJuMnkN4
Fe5DZ/qi8JBKtlaF+T4ifomHgbsAnAzu1KPToCg4x31r5UcURPdnm2oj3A72xbit
5nDQBEoWfAmytUoMChJYMuuv1G8i1Dm0L8zK4NXWiJj4CTTImM44cE/+fjLASWfI
c1dbGBas1PIcRqSVFlNvjkWgiuZCSbAOAUMudjWcogonHDDiRZ67KCgquCZUNfP9
ML39kA5xdoyQPs57hDb4JviuHP7QTJyyWuESJeSiVee6huWK6z8wTzdPITPiRlFC
wil4mfiKja5zlwm+DMly71bLdxDpt4CW4+y4Kt+/LdAJvxLLW36yLY95TnLnyDTv
q22t8gGrdFErh213gTmpdrUbHR2tKmRdkKg2cHkmPLVVcoAZMCBTatjtUp7Pa1xx
sbUw41o8LpGFGpT/9MJfBKGUu3er4jSxlp06XyNoICwIAa8ZDusBynRxL90c4CwY
7Tb4I4vxHbAWSiOSKdUPazjJwEej2gpWl2A+esbPFHCq6dNhRdcsRX5fmd9O6Ra3
yNIZzYc8Nf6O3doZ4QlK9GzcTGWiRrM8Moe8z6q+/lGseqaugInbYy/ltregMaQp
U3WZvxZ6wgii8HzPFs3p/7uaQRTRU4a1VhK/qCcpd0q2ri5oy6U+uX4d0e3SfqUn
c8+F18/o3PUg3YpVnYeLQNu6RjftYLGPpl3z/Y3LKtRg2a/5pmXjZwL1kodeYt5G
97uJRnfVN7AkkssDKIIsnVotAc1SJtvQ8DZlsiiNJvqiv45s73IKbIcrUzhuzCu6
sVM6MqiG60mBLLOTIkmAw399MQXJncdpaBAaQmU9aamn9Y4G4s2KV/iOrctk9FKg
z9o88Hntcchz0qJUP0PKgUixbfxqZBm6w/jW7Fq7rPEy3R7/vN9l9DI5aHETrb3N
VwSI7SBYMrfTOsefSAkH8S35hSoD31YZMgbjuSQj+PnYttHov+d3rtZjPcZ53LAh
cRjZ38tVoviclikc/LP/efUSdIJYjZX5RZmoqAZ3nv0bWUzjC4hnC4KBHyYiLZnl
gjTXDL+Z826WgkGbjkJ6InYmhsncMWX0JesY50nuB3I6v2HKOwZGMkkLQYoyAhFL
gjFKYqNVqYdKuluF9keYJHdj4MjhTrFrookoZInG1G6wKl8KmWEEIO/887QPdDFS
R9ZI7bXUpXVIacvRK4ofM2BUz+IVpdfE58jFYfYOVfAAW5GLi/BKAGh1lp1CadRU
/42Jt5922Vba0ajVbRyTFIluyQAvl9j0xjV6G0ZGmveP1Py4/I3eCF44prUjVejM
doMyi7aEQn5c0BxTcrBp4MVtA87qVVBsCB1RL8LL6gN8t4yAdefSxOQs4NqE01ek
Yp5JOkXHMzqC3k0oZV+g0nVwEBTejXZQefSk9um1O0+rDFit5SixWVq1CjAtOEML
LQbTRtOdJu+wQ09tRAuAzWm5zjNU8CAz4hbnXrZCFB1SV6WcU9JoRN85nBfhtoao
S+HMimAdncn1l8KC8C7VgEdR0IPzE4DJN6Wqe1uGu/x3CZFtJ4zIbQvOjepgqhDX
4NUHFv2N0c/+08stmxiUe6HGa32XBBBWuNnRK+ZNeRzgkZEgK9e5NfFAirhsvf8W
gOOU37Nyq0WsH6rjParWdR/DC6lxpMR9DClq+LW9pA6sz7eeWnXXr2yzvcxS6CHK
7S42f0QNOv0188s52nhSgCyOAX5gWNBQUphQqQ8XIbjblXOBJTN/0grMBvbAiK4t
csEj0T0cakXtgvtYpKR9HSksKprS1U+xC9pUlRbv2lpSzdwfh+JyQ2BD6/EXXnrZ
pC948rXIZYDDt9uSsUL0SI/6D94nWGOsljJrvNnJhMBJZZEpcF+kMH2NZW3tjBwY
x1sn7G85j2QcyJZ8yrFt6yvafVugYRImnWardCn3rvpd1jge9Z+iDx5kgL9PK0OQ
8suanrZQsja8Uq2zGDXGsq6NW8Efn0+wNkxwWO/er+ex4GrR0FMi9RH+Ceg5CN0D
KAGQvL3QysIPDqt3LRx7xa9Lvu93+7T+ZqbhQUNOF67mNPD0NYBWvkvDBJOKUPwF
UTsaN9I8HT47Cz7KUAvXPpzkIPFdwuvH4taMl6wMfIDCY762/UMrENKiKP1J3ZqI
1JYh052CY3tuC5oLVY2HcIZG/8dJROBI2lZZio+6Eq8BrB/kDKvCheVZ3lTG3LfZ
EI7fgqjBlhXUdIFGqxWGeXaPtvLK0a2I3P+ISeUVemdHCyTxOXOviIWX/aMh+Tv7
XPMvYT3dTlMs4UrMlBTdE5njdoSXwNRNfvuPmNvl0PPZy2Jwe7yYbfgK6OXLTzih
54ZCT5Cq3cSSjz2o9MyVtvm0g7HFJ3jIj+heY6rOb2+jLhf51Anu+lLKeZ/peOU4
iOb5etzwZSAf9xAEORI7qr9CD+/97BRMurT1g2BIOTWIJkUflTkP5I3UZ1AjaYeu
gZ8AGiorXecQQFrRN8Jw36pYRDSBOrzOyNsUhV99/PM8pRWdArH70/9LOuyiNx5j
ATkXPhkD78/MZE2XFYuPY1G93bzDrMU4XW1wTSIOEVRfrGxYq3d32zFkaBLtPaaM
fU4/TP2RtgcU1qa1e2YrN5J8cHNIfLIlgQ1GpgPhw9lefjVsRnHgFL4bx0YyNq6l
6rnmmjwFoL/Ah5gUDfh67ZV4DrwowA4pbv5rX5WibJca71thBCzt2qxuo+U8MJh6
cajJL+x5RqhzhTYRR3H7SBFaQzgGi8qzko9Kk+2qToCxYtkKuvsgfARslyLax07j
7z5UVFqnuakmO0IRGpNeA0bzIeLAnp4o9Z9sJLwMo0lfb9Okvd6UQgIz7kFC3DsL
9kyGW7G0ymfU06dfIAR+9e0GPv7LbtTP6ZsXbDg0F+WnYLqTyqp/RtkYOsGwOv0z
FAXicckq9aOo/Ax/f41uquOucGlOHNcd/cgE//29q1Uy+HK9WO40ae0UsYdgz5no
HEJAFCzrgIWjQnme17DGp/OmSfuALGMeIS29ehr/vht6RJBDIKbdpL3ixVWXWO2h
rIAwi4MUzHHgAutVuKeXg+W+Fcxo4yXlNbejJ6GcERhQmSV+4MDkKtuQEiHYlfSR
m2hsKLOV4MjCeKuV40dqeKZIjkMJGRRpOSVrg/OG4eAoAsyNzC0BTmh0AODBbihh
QHoM3elmWRWwneDLlBJUPrxppa9oW5xXdpm/5uhQ3slukgTO9jIwSY5DxzTJZ1K2
sddtPtRdDWg9Bb0TqTJkcoSzhBS1qlACoVSzbykHzcmhWI68VOJrdUIV8OzuEBpP
EpWMBV/tBgUFiZnhjpJ9hAvTq+E1EQxrw8kM01IOr+SSNTGUBQsK1KmGt1u/h6f7
7+au9F0/mYMLoPinImaVdknPWcasSQi+iW9K5ew98oY98AEnV/tLFQxJKjePWtzH
Z4VZEUdcS947s9SD7U5pyVbomAufNWdEKqVm//xM5qaa7+6rtESaBrRruo57Tsg1
lgdW4L251EkK4cqG6V4KOq9MzHUnpRYF/41e8r3s8Ecakz7O66QEnlWLk8UwRA6V
IgV236xJV+OyA1HzrWx8IDGoUQzZHAqJ97t+7XGgBrvvKCjCUhJMW3JIuSshFSld
CJULGT0jVbEmQK8oVOo49tm1bzDoQ2xP7qV09iZObiX+3doKY+3YhynsEXoQEyqp
EkT62wfOcMPYmvxXGdxDPbYZgIFTp+O88t2RypSxUM2nIEw0qFmj0UN8tkzpReH9
RxqC4bS4dUApcnasb9q3/P0bS/Enr6I/sMwZ5Xej9TWxb/kcGTj8W3lGaP0xXPBP
R2WUaSTBKCvz2buCQvLhuSjZ3mUzaepKeb5N+12Yx6LmmCzFrh8XaXHrkcfnUKRn
+bT9mXuHlDZh5bilW4dWzsD2TPLS01e4wjJ6BfUq8xigHQX/QBw3ZSg/nXytE5D2
7bJ/mBOeOSrzjRxc8BxkFggK4txjlbI6QNGQH+SSCWMLUo9iKAKEJLmfuFD3T9wK
B4rpiNun56kQY3AI5PKVQ+Y+lIdnA+poPsieSAd3UJZOdUL8LpTFRu8teWQG5T2B
Zf9etkLl7tdcR2JD3lWCt6W9jU4JKvezztjkEQpZTDaFNqp9k9mYnxukgCi/dv34
I35W1TFScExH5EiYKPX3GFFaq2DUKSHXwQp5hewrG17umHQP7RezvJByAuYBW8pJ
wgqXpEQ0YzYlrRXGJIDJeybwZNF8RjQVQcAusTeigikVFd6iLYLBh9b0vdIu5ppL
+kP/Dn4fTMj29EAJYVg50FNeeaMJ1goeKwbencLKdXxfR1XHoVVMXF/rsY5+LeK8
Ae5WZnRCIXGPpTdRk1Y20Pm0CTKkUcDrqMnRnBPICluE390RrOD3AitFmkn97fB4
6WaG5iJ8OMy932Eanjn27YJb9G1DjUqGX5Cs6rdq36WLhmADx5uNqQJUuIAWx6Gv
QSmIJhU6ZeO42ip+ZQFhuzcJqT6aoybR/7dlxE3DCk2eFdw8IWwtHh5pgmtRFZ6d
UbmETPcSNrXEaS/q5ej1E35upGDPkAtJxjUY+YF0bduAt9P0Cxxz1Ze0915eRa5e
yAcg3l9G3ps/7lMly4KUFs1QIlY5JVGLNw24rO+EivUCGmGGsc3yKuhWawEiHWrd
iYwj1ap7JppMm8ziVZnlyb90UF+cRmwUvRu5aexhHOPAHKHBQfwv1/sHNzI1XU02
r88n2fOh6L/C4XIDi123cPA31BEKFoHdn8SFASWr5MZz2dOe/16WYjF5BqM8JsrI
REoUd/CsjCuxSMaJMY6irVzolfC+S2LenTPE1NvT9IPxKqltO1iKqHUgvd7K0qGW
D91FelYU1CBxJU3uX14Po/uI1d1iuZUSZoAFhk1wGIdTrUi9ICfw2gUVwvzz+EOn
jL5N513rO1nLOIEZU9ThSjwFTpuAgwTuY+PvnRK6NAndgzXzze7+fEE1NWNY9lVL
Wi6/pdIiZDJl7zZUvSmOj2oPN9NfMvPv5J/64rkum7SK7EWLbf9M46yDsYTAJkgX
e2dN8NpUwaLKuTULvMEmXJviYDfXfC9e/TslxnUKIB9KCsVMk6Md4+358BIsBjSR
hR7ECO+PbXn208R75pJKnXWhFlnZ9AAQuWKjQ/j6u2dhbXFrKx4INaWEszYWaHOp
K9lJj6Uqu1PIfwr56K/klw0PZ/WjfhjcdE4/ZNY/un1P0wqGwwa1gyZumvMeNAkK
vPaG2bdcDOELrju7gWAihNP1SgSrDHGKJk1ZGqzB/AeW5c589abJifw9fY1THVXp
KJCwJTRktOkRoWEkRntKaUo96Qo8O+dHSPmi4S1hYYJCWAUvbIFVkbl+5gy04eNd
nitq2RzDqxoeY3ktJMpbdgZhwY2MyY7z/bPul6gx8xArLJ3syVp0fpIEFRgmtpV/
Swqe4Plr8aIew4UF3EeebiKCFALigjajKUPPsW9nVaypM4Q7JrDgm7DYsldPb3Li
ZT87wPUqSwVCz5xRbe3AKe6ORnkk2sacFZfRNojhoFJJnuT301ObMzz2N4EQn2VS
1sMi/UYPD5DJqT3EEIRcHJKJpaqjL1Q26n3ZAbIBftT1or+xsEIbK1P2cUZ8I7GG
PkarzyvU5kz35vRdbDPWgKWvmNxl8HG32XTkIVwM5MzRAF0hlgb3PhvY8axwAgtp
TIGS4iDOea3BXRcBTvGR/w9m5dGKQ9jvP9N/ae7Of401SphwhIgv+qbvNgz52WPU
ZeaPIEDEyWz+3jIKXbCSszido+e4rvqlwTeCvX1JiBIZQt0L4Rpfhe+z/ItdlLOv
eSdsiQoV+O4YdaTourLQxpLaPm73PpivoaxU9Ci+SuTYYEEN3bbDJBxxJQw0oPHJ
vzrRi8d1B2ri0t7bxdZnjwFYWM2LV1tdQ5oLIP12GK/fQEDAVhjgQJ+dX7r6RT0g
IhtgD8hqndixwLcaq9oLjwbN1Tm+goVHjOF7oGs8r4k1VMYuaPzWoASm336tgcG/
OCVlUPa4M1e3afTm4QjXDCqBg0NFunhNkYXglw12fHl2zkhGuXkiq23vfu6Ei6aI
6PTuomEz2WxfphWAyQvviogDvlo7Fy14oIFjENPKMYypxqxPt+wpuIL3luuXfEag
QWwBhh2yNO5/uhpzCSsYetq8kuS0LC2egQITRYuSlljK2SWXcKyqG72TVke5MXHO
aUbumn7gKmDE3tWASmYm33sjxmTEQEx9Gp8gpaOV3bozYaBoPllI3+kTyv8jnvzr
25SqHhz8Vpr8dbx/SBRpVkIO0FOYVmW6Ctepmna/3s7HM7zRQXtXxUDKHlahDIbB
WsspgdMnirrq6vPvw9CUf2/8rpnL0lLg1xuy8bw+7dLwM2Sj31SMEJ+p/YXG1auG
gm7QiouOaA9Ycjh/HBOlPv1gKTMCjvAzIhOEHGiVBfVcl3CAWQWLqFsaICSXahW6
r/QkUTy3ERKYE+dfexUsI46PWV0P7EurT0hucTzYnZDkpTO5q4kliNOAYGTJdq+d
eWtJJymdKie3s8LzGKSqbN/sy6GpQHVDHmZf0UaGN7btgHaBYd2D2bl3aRl0vvT3
Dbw9955VX6gvfaSRnAnmN0bnzaRhMDEUzR8gTQXJ4xMybL9UZeaXuGHXdd+Kua0u
nkmaQi+sCfY0B5quvt2lkqEHMW4JyH6f28VHv3d57SMoeIXADHnw1jTj1T2efn4S
PGH/igNHvwGdGE/pXVf8mDoJDLzg9mmMWeuQ7G10nd27uWX2+RUjum6tGqwXvJWF
2bnqNi8M8LIPKe6eaLQU51OjPM0daer4Cs/i7Ys9y0fEnNEthVbFipXWV10ikBMg
lYjV2DOO+GaxTmIWVxppLBWasXPMeW8PNdWCK20Pid28jP9jtBqGs9fZ2LVqCuzs
96YXWCTyNyDpAFqoi4PYnjxG9HfG+VkJp+MHpZs1njFCQmE+Tlwig0FUNSvkDQrP
+rjsfYxDBo5+FlQWBgQAO/axJ7sZoqW5OJgth8a4oKVUanhqWqzvFV76clrCbpFl
/6V+2FrZQH/C6Suu0oi5z+9ohxXmb7Gj+eZa+9E8YL8b7dpxiF5apVc50F3ZFchz
7+DxrcUVmXZ0HRJ3Ulj/uCoOzJWjQ+9+ORYDnly4OSHnbLVHlUb25EG6Grna/mcA
LZROfYl9EBJOims2YwWJegMYgjDzjk/y2B2GzKmg51tgzEkImc4ugKsDAob3P/kn
meFvMxYDnbsxg9uiYRdzwcxU/NJlvI7yAiYIG592gueF0QGtZ6EV71Rtd4RJwufH
oh+jMhM/EMgg8Qa1ZO3rYaJe619498yWUHQdkg0YxHVrqJeWeLBIsQWYmeyM2yCJ
/gR3iIup6ZEQfLVe0p6YCo+IztN07fHE7fdct+3UtM2CTzbc2CRMXZ6iZoFEWToM
L+2sqySJ2mDlDsDghzkacjhHq6BwutF1QbgxQqYqqBptPc7SWytiOo2NFVAmMbbD
nUFzcPPrb0GqT9B9wvGF69fUl4iXW9RE9yOwphWbCBN9AVXwBV4Y+ys2hgwBkue3
En3/hs6EmFA8hd820UnpeAETZ2Aa3LKCFg9kJEmQvG4ogWaffebSK+E6dubtuzo7
B1rOBi1Txt5rxjt5uWhge+pr0SuTbu+KwovTeIqIE4I0epz2B3incFRiAQaIDQL+
UX0IIIsbULLnmrvNKFCaeJ+s1Y+FvrpDn7s7WHCAXQAeMe7Uidrru2R274dNlnIG
biRP+7tUfmQDuWlFr9FZDx7X03rc5azLVkOfQDIjGk8QK5b6wXANOYACFX6R8mgu
MKsQOPFffMizCHJGEum/Tix8KSlh3HXQ8gIDdmphMhpUBI2jkD6hBu02zjnQSb7L
nheauU1+XxNykKxtEy5qSNm3j/KLCKXVn3mvgEVRHxubvAWIkvJG4vx1osqBzkZI
SHmmFv7KXWP8owS/j5pbeaBlaQI/oyyK/WhURaLWCbr+11kYmrX79G4wQJ8x0hJd
WeCNxI785XS8PBt3/bRhxbYR/Vd9HUIC7IaLS0bkaKzJ72aren2h7J15ZME9icnf
b1KUu6zN8Sn5D67mvjJP7dDjDmcgeXrKPL4T/ZOUADwyQOVK2o5uiwT30Oy6hRtO
EdUiVHVDDdWmryfbWhYWSaM75udEXU5huTNnMCnpYENiHsTUcB7u/jz1FIa5remc
8BSQsf0hUyhz0Za1rxMV0DyeQ2RSzJMZ197dHh56VEY3tVHOxY9RzHyQaZoEkGrC
IKsXMc1+ieLCRvfCrOZK2Xceo0wnV+OIs+mRW7NiqzwIXVtxqDM506kMfh0hu9rn
bSHUT2d3Snbx9InN3D5X/q7wNjVqJkYmmYja+4CvULblsTt3DDkX/hrSUPCCgEsS
USZ9e24g6JM8WDl/iJNCzpzJACtF7fBxi2r3ICY9v9mwTfElEkbxS45iRQivEjNI
KvLFeUjY/DNQeYaTdZh+sUSomlPAqmGKDBX2Lw0noOvqEney/Xj+bN6ZI3vtYK61
3nXZJhadwtEZHwL9vKyNi9uhRElXFF5++CBhKZjvtP70zpylWau1RODtE1SizMMB
RL1YexefNffrmhvBNwvX9odLW+rXailTZGVQcaqQpfUz+Pr9UxbMY3JnFQBpPwii
I9rNFzowXoiBqUan/BRfQ5lRXEeQLSjMjgwTjiIx1eLFvbpn4fGAx31qcwUuHpBW
ScNpatTlYYiacFHrRYCyMU+oTyxOZ1ihTeI5FtHguvB049I2cCKlvUXE9k/Gyotb
/WeC4GNmbF8ZmkY7AJspSTNJs8DLC66ybyozmxU0jQyNfkC3bVgZ7Owl64BCOFYX
5jwfuEUjoje3XNrA8Pu3y+eFT0fxhhgbtjjSLLwml/+jgcHeisLrBQ/N6S6n0ilU
g7zGITn2TjH5OT5062DPPa/+U+Qm6TvbsE0kLy5A/sw6awguVAnRQSh8ZMrxGvUl
yXDUZKotpqwyZAwbOv5igqybNQy78C6uIfyRC7Qkbn1dTFtb0xMAiiJEmyujBwFo
Aus0m2ndLoGGf+7YmmEd6dbompxxkiXvffWzNsbSAjZJ7XMOKMKIIq3AS3YAt3AR
8UF7FyixuUdanFf2leO9mstHLBh6aM+xrNBa1UpW2F8RFYiBDaju1LsOJt1HB2Ku
uUvh4oDw5L++EhMfJiLTds5chP44YO2EoHfvhw3JGHcNjApSAcRCOSW0cxAWpr3p
9Sl3+TSYEtMYSduXLOKhDBc35NW3WaH6oezjDXHs0C2iemxCX7vCqU1YTI5qTe71
A88ZmDIoqYL+n12a8BGVk+VwV9VzlE7vKA/g0NsYD2IJU70GdWjpbkYF3xcVZjnM
LywOjqX4sc+mVCqaGamm+NwA06D5dc2js1SwOlZbtd00uGCV8DpyeVr90Ku+mPgC
260wJclStmyvLAeL4/o7fSGiQyDHMzAOSLG3FRuVx/RFHqiOTLOPPbCbHhoQnrlf
2L5/3ZvJuNyxxI64mJKCP7Fwm4/XHhzOvIP/kVLIXCFuwi0gRKkN3iSeKnWr36wI
8HUES+RuhcWf01HSZBqPTv+975Fc+L5TJ7zC1WaZ4VZx+8Hh0NONVfkQ8E9ZpXhj
d3m+kx1TsJAzTHDaE64BndFe/TTymHkjvUQRgB26ULyqe+uznm0/jkV1eIVlVIBX
Z54yl8yF9fQZkPlf42HFULwINnl3LaIa/z3BUPiCkHn/psMCLJDdQLK9BlhUlRdk
hFMjgZTRY9lKjIRHUARG4/LPi+GCN4AOk2lK4Q/6nlYHFlRxukn3wlBLjnf+Khou
lGIiHlHKfOY4iEAT5HUQ9JeruXOzBKFtjIxgozGrLN5CMUFRww2E/FzLBa4Ezcd0
B0v33LNXC9InzTqsKplqzYfYj2vvvjIfXjphSY4cZQps+W40MdLJx8bLLoLAUP7p
tw7kPSzrZrqzPCY1fUGBsyrY3OFl+tXg3BOccUSmzYz85VkK8vx50F0YRgPSFWw4
tr1YzOC81DVCpirNPNQ78mAPYVnqeN9F2RJ16aXiu/w17A/xu6Iv2oaZAvCLg9DK
gcheTfB3OtRV19FKr6VCGnIWzWWeL5WQk2e6UpPx9tJkdpVEYjLhsSb1ZySzCEZe
Z99oOTcLI6YCVlK3p05AfrtKhEoGLLaRYA0spVn4thno0YcpY19z7YYoxs7CLsGd
yIEp2kyAY53cEs/+arFdEF1/E9n07/mV0MfdkgdQLkuJJ4pEXKWnrDZHVtvNJzXf
fphpC1QRsga7igubNG3OrZmA9fENBBWQek+zUbvt0u+sYeTEPfMcO5hO193lH5cj
uMRdoO/IZYMmh22FQtRnOGm4mAuO32Ao0uEBFIijVKokTdvZ8CETnRQlPkki3Sbe
vVSF+AaJ+Z31T6Z1VWFlYczptwrr8ftzTiXHqdUmEo8QDWtPnshbyX1IGz8UeQn5
GMqH2VYQ24+Frh+QvPxNgvoHQAnzehIm2tAGPkECdA/XJ1uxgIzlogWCh66X1tPs
9tb9rYL1XbdpTXTpA+QvdbyZBHtY0W+bNipBMjUooZ2vPBu8+eMsj8fO5zxVyZY3
Gv11PusiaWkbo5+IuVZjZF5UOtr1wGlP9hrz5Esx5drEYOCUleCZ7OPQlOW+5+GR
FIULmXWX9FjEU0fb3rgZcGWc9j5wfuoQYwRSKKUz2TjRWhJUawBLM5xoZIg3mzPG
+Dgj8yYZhNccrr+VpXUpjUBqxOW6GPeRrRgU4Z5QcxOAU9fPGzwNkYLBNu1KNBOI
p3PtZKNUzG+dylT95weRZq/TLC82da+nuorSInK1zy0TNrXLb1kfe/NJE4cQ6Bff
+7pVYPJckpVlq5+xgUEE+nC0cXrm2uuo9wC6+6R45SzK9wkBHYGJ+yHe5196Ck1H
LO3Mwb3BtFQeCXimOupjks0ye6PMsOMD4bsAkzgylB/YMfs8ElzmfHkJVaAotNvb
L3R0SDeq2+XUJU/pFF9u0XGwtMGriMmrqUBO+q6AS1Tmk8wphNx7uKPv6HrkAMEV
ieJ7aD1360Y2OshY/gqRj8qMR0JnWtycH/qKcoMa5uiCv/sGvPwY/GOwjVtD3kyD
eZMJrhMSgAQMOhaFuUsj3DlA8jmPRTqKaB27cRaGiQanw7JgLaMXUi2AEacrWXz2
6l9oHLhfLxzro4Q6DuIC9sSSVvJI/j3Kicl1odDkGo3pu8/xOjIpCG3DhgKIf1pR
JokBT9eu3y79hzjhv8nTjlbmBJ12KHEQRfJC27VS3ID9nbSjMeSeTFKCl6E594Jl
QzAdqRiFChsX5ILefs++OzhqLrb0V86aBP2K9HvLEMLsHeGYZsDHJXFlje1IpJD5
CJJlNf6t3VZqhDEmZvuJD+1wrCv8Xbn/pLLbA404gB/3weNaC1Kwcw7uGkbLJxOg
Y0FhxyOU1SEcCILImKCynzfeYfEhwtVoMjSDHwJWleeXZa5QG5pCISUIhgYIK/+w
EKzmdGp+l9arq7qmGXV0aTngQCnJOj4RUmxi7Mxv0dh5T3W2epzLpzpBq6C5f4F1
ImjOQPUQ67KBqn9D5huiJzImU9OyaS0S54KzRh7NCHcla6oaZiMH4qr2en8sEXNW
beIig1xWv971TB7imiVcbECHhCgXrHBb1LqRHLe5zuIsFFhOhWd29j7Iqiov+EA3
+sTErMMapEmesPmRr7sj+qWNbL5MtPPkxQW73n0W0KXfjFDCnp6lh9PoA/lXSRgu
D1vUfCqW/M4vE6TTQbwBNzFayEdEcGejPagJnG3qoJfcbGfsTxST7YZZTfSESjA0
GSBtqlY9nG4FblJAH0AdcRlPiUJ81wT4f0RIpQqwNuxAjTnEc7HzkzwtHYoVpZH8
RHTB4TErQ8L4p6BeusUK2tfs1RoLbKwhf2lvVeue82U7SXVhouVlK+jAlG60Yf9x
eZavyM4B1jtU9LgbwEfyrtb/VWOOzmqeo6hA5RfZWLCMOpCjfYgbrLRN9RWB52uA
H5GqeSOFVtvFIZ2sBFqkj1tCH7kcFtQ80cyfSq4i186OzftxBWvwlMQn9+b0gi9G
a0dGj49RrRlT9SM8SWZj6Sl8/WDn7KzmevkwMjFlbDlKq4e7v2Atvf6YvRT8Xya1
8dGqDrkllpf87A/5Yw5dKngbq3qUp3nnq07xTqCSi2LWgmyYdIuRB160AT5giWnY
iy79RYyv3gNvCzKkMK578Y581XzWwZzdN0LOHYN2GynEcuLQ5uJNM5cTdvsNZ0Df
bTkc3LcjaD/O9BL9Q+RIuUBFrKk6E4wIfwccrsoKRlD6a/mZn65HyQtt0XTKh28U
U4xnqVBMDMZnjhrXrouEPboQa146/9EFYRfnX0QyhA1y7KOCEVNoajb/LEQ2ZuD2
LB8yzO7mLkj9kRLxDuodf5KOMpEj88L8j0Bf4+oZIqeDj1GkC18pd4mgKUTGNEzy
qMt4sKG/NikyDccBVSOGveNxEq+tED4EaC3QnZtlDqOoru7pMCwq6QwDI3+odAIA
oKnErQIUT7EAy6TdXoQSBEviVFzCVREgYr122Sg+/a8oqqA4NzQTD4bdTxKLnMSa
tS+1r/UVt0n+1aANLTCnucIPcXErd5WzerYdhMYpheFRoSuERKalaytKPPzdFzir
kiGvjFh9TctFp7o6lFWE/cKkrXn+jdCR9em/PIBMELVC9+rQ52Z3dOPn9b/JDxwl
RDb/+z0NGAnNgfkm65697SwFXp6XvhZw7ciP7oxFdOQH2emDPEmoM2sZOWyYyKdR
D9drixPHlGCqvrPDd46mNtAlnBgGdZqzO1Bg7y6Y35EsBtR7owOHcTyjvpV424/0
7REjkSS8l66uYqIYTij31AxRSRurdPOVrOvcir8qtgNFLHJFbOR4yRkp/GWanpWY
E0KCYzAeyU2jE4NEX/ud9O/DVuKGkR5lcpxB25XcXVq3M2X0FmEhGOZCKM7gTjgH
jkbnaiCiURv+VklEtDjheXWgAtI/NQgKRPI/a5884+LrmqEQ9HuIGkMBP07YmJkd
XHUJUFP1K3SBL5VTnqJaqkpq2NmEW1FGWqmFyB543H4ktxbmwI34j9Eo5avSewA7
AUHuM6QHObt4Lzp5l7WYKitcefLBE5+5myxHRRtsPy+jSQioh/jQxgEceBdIwjyx
XZVVCIssvjtPXparqyYkuCN87siIeoMg7KN/vAe1ABqpxpAuou4JO/JXw+UsInfY
r418VM7EdntlM0Ejma7vSusz9lfNt+Hk33zDlLVuOAta+0wiO1B99nQVk1GXT9o8
74zQzuljyV3a5rqZBEvWJr4NVBwkRxV0kv3+uVo5J17c4AKJjXBc9U3WtxqafISV
qPwlmcX3dI8r2sziiVdufohpc8wHNBbfNxR0aUCbD4SsK3kAlgwQsT28kmX/hFBB
V5a9g/YwsH2yobjEnh1d1y03DRUk/9S5xaIFX5N59LXyT6Rpq9lvikf/gPRN3aR+
8ZjHbWViZtxhYQxeBNP7fenKiG/i6+0DJEv7O85+EfvzJ0tQloAekXKZttdxi/sB
9SMPm7nlvH60FUNymMJi+OBtOELnSB4Hn+UrlZp7ZCoiLBoPk4FBoKl9XycAPcli
236q0DIgwPpeNKALLqFzfzMMlVfBju0DwOcFFA6rIdqt11uLxVG6Hgf5Mz4jRhb7
JL0jqdLqn0//qC9oRvSOIsFPu8hdUuhGSAkKE20IAsMHo/alUZsU9nYw6eiNTSQX
Sa7ioyXGkNtnjvLF58HF523XzhT3DHWZaevX0V1KAJHMHMhQvI9OAKN5eIdM7xO1
BSC7X1H5apjuEE4+FoeLGTmFK8S17pOjbBUpBH1FDyfoISgoRFYNN/GvIvENmVrb
0R4xKDSp3B4IPLLE8svXVfaRGIGzOXfFM1QV0XlHwcoLaQbNua+IJs7SXTrlp6Wl
Pn7GLJ2ar/JX3K3joX4w7EhFtd8fohSEsA0WroT1ouT0JK3ZhL/wOdr2VzO1bGB+
VTC4aeqXpqtUHxU1WFqwOnYF9iUqqz+nDBTDO/oXctgk/lpP3k/vo9LfLN2++aJ1
1CRZdchUqAkvqzegqwv+7PRKj2O/FTrnOn2e01HYIdqhiyUD+hzgi7vL5F+Fu0LW
NmgmjitF8U4WXjNUG+u/hHUukEugSwBprkoIEw5VtcwOTPC2AjNvTurXxYbiAsv1
yxS1RvkFGuPy+UtzSi9Tht9ZMY0b1kGRuonU+xcv0Yh16laFGqp2YS58mKsNsUC6
fzS+edUM89rF60Q+96I015oX5x55QqUilISt0UDHPeu7qbCRt8K6eV+13hr+0s4x
/VTXbeD8FUAQjENWABCwNwYMgss5/rvZ+IdBFFi8QcP5/y3flfe5KEGO2OvhtzIT
M/Hr20J/wQcMbQSePmKgIXo9SYW6MulmZp6IQnJzBNmgMjmNpwfPB34sQcmuO3gI
VPQYif4ICM9TqwLncex7oXV08y2eYXBIXp/TEl16DphChdjk4L3oBuvFVyPw8nqr
OwNLwqQkfwvsARcuegOEFejZeZpbzSavQdIFb4kHghZdZUOjBRiNZWXcU9Zxk0oB
rTp9mgejeg8CzCQgCdGPieF/eSuQt3078mhYZLSqZudP6MUn3zTfWiQDAILJl1f6
ELI/IhaqtX4f8RmS0tvKyuDUv8Te07ykWiOtevuTK8regW2RR/Ab0c59cECijI0V
gcVw+5UScz1Xa4ZSuJwm7JokzgfxWEKlajbp0TieLxoMXII87lnDjlHlxKjWZzlL
eOS2EQo5l5tGg3PBqMoMGMvLIaHWsO+aGh6WazlD9p8AkkLz3BC1Mv25hUKRJ5xt
9NH+IyQJFMyfShkhV49AIdfXax7ii4OvaJkBmm1OaT1W9ZhFReXnGPFq5VLOP/qr
ACdsrgkCi03oD4zovP+n5Tw0L35AscyTaCoVMHt7zptjo/37vsYzE1ykoSeB0RU9
Q90n6jDj/QGPSz1yxUHqOQvK1XakoPkeyx5kglV/MDZT0BPhpkHnGl7TW+pHlfko
qVca14VRzoZDQphm85mjc1rZp0zaoklkh16JOgvF8BUYiwO01R9K2zYMEGWNKaTq
l+gCrKBolsDUxZFUVIbQUOBtkNMVjq37g+XVGKNC5mQtoqZY4C73I6MgkmBrqjZO
GXbGhic5HPrnP3QBFNAuTgA4/dGiwghABHWZs5bcUn+ZK+XDXVv5ekg8qAEH/rqS
kHswJDFbzhSfe997BJ4PXFLK+lT8NljU0ApYybzbhopdQbW+xMXfea6kxvmK5kRk
f3WiKEnxE9qMMkbK0SFSJ5LBxttMt4tysMCXRB682+H6XJLQGLd/X4ql4dxWU4S+
YMhGTrJZwf9TAMXkvC2iS8CnUaYWDMAEf+H1qLUPzVNXgO0aBqkGzuPd8on0WHwY
Y/hP1FH8knQPw14QDzpCsxcVaKcSAmeSK6F6P7FW1BUcR1xgzO/6knaKOcT4IKFW
IWWRTfADafHWLsCbkPwRtyGaxkPCyAfBg1kO02Z91Cw6XNxHgdAVWG1HstKMiX2E
nEuZMl/3U/eEYxG72g/Q0fa19zyzPXk06JzwK2XJhezF0Lh6AQBZQdEaf6quLXQi
LTQ5F+hGX6MIDO++YAKB59d9KiKH9ifp1wrDtae6WXywETY+Rd99Ar55+xZuCYKH
0ORxeI3uAz+0LpJz/LKCdob21G0mCXnwylPXu4aXjg4c+OgL0t8tp2dXb8LRIvx8
TnT8e9Mu6FIUGJQi+8wAg9OHwHulExUfumwqVaRh2IHivkyJIaG74xUyceJ5v7wu
oNKRV6GRXXfxWtnQPAUxK1C6Gf8tf00mxidUVPTbXS9KP8cyW8AAc9pgxzjv7kV+
QtkvfN3seopK8s6DdiMoteUTS62IBACMChLP4s0nbbaFC8tgtx4RPytKRHmEdyE9
j0qMKXphJloXZcDFI5t2Oi+q9gQv1krxvzp2HyfXXETK5XL+mMnWQGnjdvSLa40P
0wE4q48itEe6ekpXzmQaVK4efsGIOI4H2VPN6MV2F0APmN+psO+abCaC92LoiBQj
9kNAPAvlOBsFGEYrYHRZeGG89Og7XFbcUjfbRrXw2quuRgSyCMeKf9MbTbNhZaKW
5fW3f/Al8GulVjJ3Nj2wirMlkh5JZAof2X4PA0sMFgDNciCcb8Acx8pB3HaIoXZ3
og07ctd/8XN9tGhse7HN9QcCnh5GkMzx/N3Xjg9xvUU0hUhCC7mfsZcsGK2BJzwa
m0H/uZlWihQOBrmQP07WXVRnqa/TRVK53ASdDc1UNMebutsSoc8QzaJoCfpgSYdx
X7xiAQhC462HC7DRwUlFoW4lMiKbzwvcPG6IahoOu7dO67lb4tsGO36F8PKT3kbd
qB4ml5RXNaF15hc1RSQgpNWBttwgqRwRkr4bAmpU6qPyog6qYUd9aHBy++45H6YI
GPRuNiymGrGLo4y9z6YiL3fomH6vMMFZ5WC2WulJy6EgIKymFv8q7LpWOsxmEYX6
5+oPxDI6S1V+1wo3CYWFydQW6OKzK47802zFop+WDh3LrL8E3IyYFamCqZajpOor
dVOmrndemBzgkLBegT2FyogxPdOzjwwjzSHQBzNkIa/zLNuChTnDlIAnGuImbeS3
amFQsk/eHysdnRHrfVngsSelJd0ysEbC5ihPNrehWGFFItNsGj1EmxSljeQH9tjG
Lq9LwyPv0TCBAgDBsDZ6321gtiXg/UNmzU1vrU9tSPKbXjOkIQZLbrG7IflxfTGK
UkWwQ4osUKixF+4rziCwjEIHCjW3gHTIWeYfCrI1atG8dTOcvNpaSaHkJmGrYJap
iVrgggwe+7SBYZU3pGvM9gH9CYD5moPx1BPdpfwv855fafaP0/c6MNs2qf0IvKdA
Rp0dbzMOYQPXH4OvCZzfYbFJJXi0aNNgKxXwq+ndJr+0Pc5RbjCz8tsgKMo4GLzu
zIAZMs6BjMarrnxBaLdslaj2jTMnj+Fpq/lH7LLbUgh5kfxhbQ1Czh5pvfzSbsRU
YJK4lKAEz6pNPs5f5oiMIMyd8VCp+M0jEDGNZnviZMeOVaq4dCu9sFuOOJbklE1W
Sd1ohZ0U0SoK1p4KlIqm6TQFxdFsUlkdP9jEpYcWp6fki0zx0u9rab/ygPis6cys
KbtxEcC1MiH8NRmwoootwRxKLUZ/RyPJPnLC1h47MyHedfRUwx8Jujd3oCIkA0FR
GvDJJjXi48t12jmxYkYUc/MVIQ4jy+uNYt+X6lfvvt3HL/GGzTXlujnu7Naufu5Y
6Hul9Q4Ngd2mpbgGKVgbgiPIPdrd5DjzmmEaDnBYlHPJyhTqm46XkSzuJAwHQkjj
xx8O6nwKJQlZmMo7D5nubrmAMtMX544altsMvtk1QjP5UXIHDz/gbBD87r1+3EpF
VCkxcvpLbCn7eZg5yvv+Ik70PQiVTLsCoCrF836Lzj3DESu2IitPW8K840T1PKqa
LmkA5vJ1V6EIrnzxDyVjyYsozBDs+VlkIOwHhp4uVXDNYHBY6OK0YDK1+0iCq0WQ
WxXv86SSR+OG+X2hgS5VB12Uzx89xI7En9HUpwbpzKN2CwSchh5maTfxed/pGFiA
ROSMFFShg8vIECNXTi5JQ5lcHPvqH/kgNLmK90lKeevfFkRjNJnDdymvcmQ2Js0L
epN2yyKOo875N4KTinJgbriNCeMwyKaDG6LoT0Pa45et/Ra0M3HazO5Wqz+SDMux
nzhWMrW8SRfdrvWX23ZNQMYaA7prRwG2cxwcY/zYSRI7wQ8Y09m/hjgNVhE/KM9Z
+fHwU308Va1qbOh99ryBnqZ+/kIu8FiNDd4x8dDBa+W+Uv579XK1DW7oZzucLYWB
v6vWMrL4uu1CbgCu/x1viUYwvcfhnLlKbvnOwebJcNRZK6LEIbdq5Gi2QNdIV7oz
IB71wICA2dK45ZppT/68oqzAjzyiIQjAS3tqiGvlFcGpMgzcknOWV94KwO65J09I
F1PlvYcFtBmYfjgM6aajCnqxZbGoMFuXLB915wLbC7ywKf4PXzt+km61M2ZD0veO
r/ezA0mJX6TG2Zqnjr2zZdNFfE5J2pHp/dHvhRgVaW7jDhFp5i3gUX2UpLIInB6w
DQaVHeRwbuU5fnp83HINyN2Vx2h7zcUh/DRjsyoCcMLxxcb7jF3yn5mv5BIxAVpu
Kf5daW9MVZKDJ/qHQvneWNyP8EfjYgOakzxpY0p09vWQCCV7SkKwxAqmOhKTXPXY
65vYRF4s0awabNaXToNEiYWwtsMcws7rw+Z55d3mqKqXIuuzTFA7MMPh0GOBPuJW
haiQ0gY7yfyH8Jswoc4znZwoVax+ol5T5xaH56qrnCx+KsfP01/C18N5xoOQkqVp
TNO5NLXezbWuQh3ojvbrvMsm4jpfTBAfMVO6s62T2IgFa5TjEuJncmw5zJ9FdLC0
6v5PZ0TTKi1HDVtcOikSsHtsUR3fFFNa3wY4xK36ZdanpfQAFC1gK/o9/xbJqHfS
b4Kzq751AxuPJkhhupgBXShE0RkRgUC8eZgsJQfYhEuO6kie5lFzVT4fa/RG+o5A
42m3UmHrLwjx/ItX+WD4EpN5yQpF2bd0/1sejS4nkI6BmCv5PB+MsmrbKScFnFN3
m6oytYk79rpYs8CDy/9qHAeMbItHRxOGV1HnI9ZxsZS0IfV//fAU+i2eCza4SL6N
D3Hloxnd9cZReMHMBGNYHDP4hdAx4MNtXC3ar0saMpol9c7Q6RIxcz/FmJ0kxR5L
QTQOStG4Y7no/99OuVCwtbFdkoEYxt44IvNJoz1jxZGnTgaSAXWB2piTfAwazAqv
dss19oNww6fP5XKhW68YYXz9y0Fgf2SXrQvY0iSoM2bew3zCc8kGLate/c53J949
1dBIGlYlqkndrY79r/vv6ybck3HtgLnVboGBMJ096GA6BqFz3LKRmASEQdP3tAbx
6gVN4az0kSUueP7EBI9fPrDPp00Nbm1LBTzn4bq71+uw6ON9mHadp0Xp6VdKMawh
qMGv6T5ERzRqm93EXkmGTVe6ar1/wlprjOpP0snSmrvDNCo7a2hyDCQmMPqUjjml
7Tx29EZBRThjrpktKpICVyANB+/M13kqPj9nwW5eEH4WlJ8ClFgWAMv1DJuP0zSm
TtQ2EBY2A9mMmV3wv5Yuq2vrZvHrxg7UDLdVVuoJfK8sE6NvbXqxf/LXjqs89Chb
XTsWJNMsq/usnYkd08/WqYk+xayRJhgE5OYt9DhlsxGvq6GzTJq5IUn4Lz1VCZQ2
eqshf4JZrREIdaylBM0/11nzsJojpmngvtv6mxm2CQO+DMRdQD4WKOggN0fffA81
K1bpGAJ7k+qQD6+x23UZ1Mzr7Us8h8nZpTXvt7oQuo5ycA7/3hOfKoxhqta4k864
cHyrqmYpnGHW3v9xeJ9N15uS7sPK4JYNk229FJXqEdFdhzOmYJ9jKSM/Ey5tONt2
l45/s9XK9crlq/GlilTqf3RUtEW5/QNa4paOtMZp5gCFqE/skTobaKUdHrylHeWk
MQc8tXuSQcxSVpCMw6TSNnyfSduoA8VK1zr33tWHWqcUe9U6jDmA2DsqDX03lcHH
hTwg4ZmTOiHEKfy5Hpr1Jq64ThCR9IJVbD8/PuuVBO5R2+NmGVR35gj55/G5IRCq
rTxT3+Po+lcyEk5IL25xsAA+TmBtAKYLukurhTz0cSMeM5L3by99/RU5ChEKYmAq
2dshCME01vp6vc1oCYSe38ecv+3y1DJ+O68iUkPZkiSNdHkKnsZFgJ6KSBTC+OCB
GDFCMM/FbPgoTagxH8kUu/IwAnRcpfygjDRxlumReVGrijlEFKqutIuL3yNyASGs
Wyo2oPgH+5jiZw2kV6L8dwsPz2mp4vxU5tAAJjM8TF6Bp90TS4mIvDLnKBnHT5ys
CKSfXduk8CPYV2MCWjVT+xOAQ895231qkwfAmpdDQONZAGeY1vXnytEz4OwN3mxh
yU86xRMzfDaFGithDebbdWSVkaqxxee+nVQrQpbMXUqE1LxerB8juHFpJn2CJe6G
bpni35wRkeGzecV0eP3c7jzB92no6+9yDEZjin6aDsKu3FEpYhkVBOEgamSb1V5i
vs8LyFcz3ZUWJbtIN0q4fk1GNysR7C3opZzitgw2kLBPtL57eMtaTzQadkCHN0C0
LEvof54qCzBFvOinVHQ8bZ67JKaUZAGDh3E//gLrMlI3jZeZSelgzBmTr8TIKC82
B9oglkUVHqXdwGsu2g5zTSkeuMDlUJGUfDRSimXwsj+nzlYTkv8UJt69xRJO68vc
J2HbPoz4GXXsFvzhMTH6CAwyVv4cFu+K/vtOLz80T6UFpco5QDdK9x/VAgP8mOnT
eU1qnsDX/75yP1cV+ZrKC1i5LuiPTPCqFyWbmAJ2fI4XlK0tzEL6kw4qs5DLaf1n
e1LeF6s4TD2Q/ksICqfzZzSlA0sMjDN0ux2MhqtbgvQh+MW12hapgv5VgEX6ZiSH
0Tt3g7ZsxfleZQzzdheb6wE0SQTWqPyyDbK8pELAwuPkrsFibpNYDLbTvyDEGjgL
drJo2o/Cd2bvIpwimGLPHEPuqHXcdy6jG5hITOUqR9wcTOdk10sGGObPbX95t67j
kBQUVA+lEzn/c26M0eRNl+zTVlfw+mJsI+I6BEH0iK3PLsfePAdcH4NzVQLiq61C
CE8K5ygKpYjfLD3lvbSemMqLxDcevyXZRxDsU4qwsdgfUw33MIGJp6Qk2EF6lfQ/
rXorJiHAp977BRxdzxqDKFzuWoSXHLwncFBQUbPzevaatfk6vPZpWk+X7HAvAzWO
jSb2lxhUUQyyqYdgad/3MFmWoCUfTWzSWoi3fFmbSIi8+WyQPNpyzeWozkJPq0Nk
I1IpMPfDH+E5AcOoxmxp5sWJvAjFJJeXq1io6tPdmU/xbxxYXeQDFyBILaMRz9D4
Dhx+ppfA9oqsNy1B7iSVotB85NN23Ey72aZdeo51wgxiXi+HSkmDn1lz0KkMD0SZ
3sb8HH2PQpgP/Ew05WPKrJVMNwcSQuNvNzn/iKfu58aE5QH2/eQowPJYVulZ7jCN
UVv41AmUH9yTPV9IXvPg3AJ+OFReX4sdXgqLCMZsRRm8tGX5NwmFhgLKDlgjJOpa
+tUP6XVctIeLzhtaul1RxlDpEmYTQee//F11fYVRSkkl9TtcBzDZ4/2aGU/GeD8n
ti6yXEzL0E/WLHQOA6j0Yhlvsc59i6zEUak0cCV3q7R7ZLp8CSi0eo6eFEF1Zp2S
jIgPh8CxtVnlPhkaSPA+gcjMyTpJuZK4l96P0IMohAcubTj8xJGSHo7YuVuqWA/8
q3Y7RNzVEIXqr54OzyqzYCkGAYx2619uAUkd2rK5fUB/XzJNTqzibzspAgNv0t/D
kfJfZfWrbNgIm5vip0t2zeM+6VDUhfCbQL/33V2lh5S1zfdaxXr2p/YhItMj8Z2r
ZzeT32Y3voNtoiK0nFAKA6MJ2s6xjz0aamlgtDPCRNoAM4orDtqZDBdXMeM6V1OT
pSy1zqBfB6jaq9taCB3P+mQXl3Bu4tgVVwYScte+SpVC9dZ2pWPfwhsXJkG+fGoq
fWql/D8TxQ1c2KsAmNxD/ZOCV2xJAVuIhtYcHZ9vwqjao3VDCKmiIYSN2eU3QKB+
ID/qt/Ivjz/Pb5BP9OGCKVocrFH+5cpZOfqj9RzxI/N/lQbEOECnj43g+zFLUcA7
RvAxkVSH/VlysMtpeAWFSimlVq5ZG9xgWRJSWuic2aAQ+yULrSvo/iqnC5+dsV3R
bJTMJvgzN1LZ/14+hXGjCpgjaSlIyKsSvlWeykY+HPevP9XUxldC6vF9VirBK5Vr
rxCoRGbplwFebFOBPmjEND9Pv+8Vbm6omyp6SAv5EFaaztnZjqyIZj8QUIiHbPzM
hzB7nRKXKnO39vhMK+wI+x+9VVZ8GJ9098k7HbUGZYLfoiV7Bo5MO0xsUZjs2JRQ
OgpnBiyjBvhXrWNuk8+52eoeODciOpGCuX6OB5v+BtiuqAW85l+/sqCNOHDyZYap
w0peAjG9xe2NQJS0uygnK3O1wW1UQSUOKsAluX5pJ3fUTBxET0OdTxnAJxFG/wJA
7eO+1dfx4H8bqkp+Lgj9ppynjM8wr8oI389rjq2TZwK8Vc4wKxlBiIasfSqdmLug
mcLfyz3n4CaY2NTbfP5q62REmTSN3K5e7OAjFv9659TdGjWPAIJnEafSzPDjAOdI
BJUOvNTQIY3w2bittSqPS5KcPjlI8Vc9lyNfJoqLV/CVvegPyteukobRTTnn43g3
1PdbYfouPRrGSZnUdF0vgsS4zIknzWCDpdatEPkyIZtuXTirdrRLpCfpsAfuSW5e
9b3+KTsn97fjeynkDt4rObc32P7nAjZipDVcmoCHklHgMnnAfsP+/K9+FCtXzZBN
e7AcHnbylDPs3jUTU/dpb6VLJRxCoLnT83fZCulLcM/LbwG7RpzwTiWX915lLZuq
BByCrR7YVpIzKVCsdRi8RLYYMP4SENo9buADfal/ZGwwpikb4LWkz+6b8wjpBlJC
sNWOyRo6vYjQ2pUbRSxDO//7hsKpCO29p2k5nUanh1/gaiOI/iCSqitqsy9Kov8c
o1EbuD3clgj1o7wIeZv/GqyE/IcU4lV9jbbO8aYlRIhHvoBKBzsFpU0DnAAG+J8B
WTwbkq7zDb0IiPg9b2YIoqmOedSVSMu9iwXwQJWl/AKcfbp8/WvSMigcgfxTgkSd
bjXn7SiSDW/2JPU5FMc+bcCFSmV73yGFO7qEo4aM3ErW8O0HxDrCvhs5BxomUVYo
hYofeOJECCPNBSIwZOT0OArjl3Nb52VFpA/xYcH2vezH/ndGvYyax8h0FkalaHso
wCW8kq+UzFhLvgdHb0qFUM3rmthEVoq4QAs9GzysNPmChQs3GbpgWAadLmykO214
vVgUwdFyYgO/iMq/dUwTcxxQrIKNln9mCg04+16+pdEmHBY+FgsNM3lvM4KPXHLt
/OkHcW+3Fv12lWRXC2eRAnYAAPJCY4Ktkg7fzVniH+JEDTN7OhUo7CdH/xJ+PuQR
ibrwrBnxi2GcTVQa8bzHLb/bkw48SFQ+JfKUdp6tculwphEsY3ZU5q9qrwn16u7I
Sa4gFzh5cmBrsT845/VNni4YUJ1fOJMf4G2/q5Kev3zYk6ORRz00hAZQosw34bxQ
4VNef3c0IrclxsV+Q6+LwiljH61/6qiqaN4R0ka6eamwTF1a3Zc8aYn9XeICfEHS
l6FjGsHqdhYwoZDeC+L/Guma/7oYo/6rUO1QHDHlZq4fkjKOarK+wluIuNaB3A3w
Lh5HtO5QpyopDwJYUoYgdKo865ADtBpoAONFkX2/pIsaxghwrvRKLbD3hEK3baHa
x1OKdAY/733fKEIno51OrUh/xHx7r+xhbZXxwDvUrtxAc9osNm8T7ZjKyEJafbh1
KR0p63V1BfcZwZlSakek5PFxOdgrIRV3zRByWqqKZjewL2IT1k1M/sksKgwCdYIn
ASKzFg/ttOzA/BZHHgiX2HncGYK/oj27/SYyd9suMj+6VPz/+HkJNRyfPkJZZ8wK
a/qEKC9mYt8WAFU9vOhZuxuhRouMulMpQxNQcv2e/3Igoi+Pyg99YCWVd4PKzd7G
eZ1Y2ldls4+xSRh7WuJ8PRdecD9Ww8ju5Xef0MuYw4HIQ1Vg3PVT0Xb2ceQXmpQW
deuNp8O5QrQ8N8AFmoF6ISyWwiSoQRRqoy5rp4Nx/K4Va92vwgY0vM9oV0enl8W0
WuyMDHH8lQpD5U97p7DRNCEKTjgPYGiaCV1n/1hRmY1EKjI6vpohXA+S1DrJYsIx
omt9Ld5WLdsVrGg2DtflW4hFNvsdZvs6WpbS6NBkXxOciycZD1QUL9IvbnkI+siy
KtjNWwNibtnFvFEezz61tY2Dyhwtbe8VlYRM0Thx4m7bBiONXOQYXwBoqEHYAL4l
cSwqBqpC3RFS14X6v8QRRXQZ7Sd16AltRJghUv/geXiH+VQswMQVQ2MgYFdyYQ7U
PrDCf0to0eWwI4AOduuSJdxOGeFddNePOFV9z7Wf6LQ9dy+iQAc9ME6kzazcc6Rm
Txl6CpF4AgZPOPIGzOUDWVmCQ2AozOK6EsYmKEVEjdI8dKUIDIBllBiDs9qPAzM0
EqRnDtuZ94XbSnNaRUUlw+eG5/A5CPQq+yy9VbVQo58Yeu7McNPWrVRKndr0q2YW
c9Ehe0J4c79x7eDv2coebbT//Z84FuwAjb28cSP2XpEwDjwpW6Dc7Dw/tIaqrf8U
2zzTWvWI3BDFBycRoYuxaLE6pR6rpimcxxqHSsae6DY17mvo8bimT1+6i0Lp+Xq9
GnAPWeTy+5tEkZGo8Qsy2MQAcDmr2uZze/n9K9XmCnsh8SJqWwtdbH+kNOtqlj4A
aBHx+H4JckT92nsXqu1OhcoMRnA9aK4Ro8GPMFip/FpljIiWnT/PSwHGhh/4LrDl
2e4pd8Wi5N64YdmX4ROU68HiBVPyYwnFYOurLtCGNVfJJwri/vaICE79eYGtY8F0
rOG372PtcwAsAi4bu5a6BzuWdUxV10FjguiT+yBdRvqYKrdocVt3jRWhSF8iR92S
soWNUXH+KKcKufBsbq5HIaT9NUDSw1JhWnYc0k9ZkgI+NbmkWjF12+WM+Dsoaf1D
OFbuuub+Czzcq980EBeaVDa0QkfT3jJVaINJbOGZWpVJEl8jjorNvInQvM6JuE55
jzH2yS7C74P1WqaCohNTDn5uJkyI4j4/vktYK+EIWT6/vPUYLF0NyxL1jVvZw7A4
krF+uKwfcOg3Guqx0phn9+Qcm1C/2Q+eivmwgQG7v6bACLfwq6ox1kURNH+BCOjW
OSophRH2gbC0w+J2W63iehvqBqRL3eWNQ+l289H85eiF2Z+2WfDT8pHTIOOCjyrB
XQnbQoDB8rsQ0qbB2/WZzBNVf8DdqD0ANj4u3tr/Flt5vMaAtfRFdXYyHQUnurZp
kUqX4WELXOl2RoQfjYsjA0cBaL2j4//+jV0NPK9q/ad29EKXCsURWH5FM5gejGfm
+KNofIR8tW5gdhpSnMF5QBpcDHeBRu9Xak0/8apdUCOkP6QODUVKbTipX/pfLgI9
1yjHuFv5uhyRy6zZhRPp+vST1rgDxnj6fRejiABLXpnwADPn3QDXOYaoPTN24jpp
uEnqlmZWpyNF2JJfKv1X122zJd75m9znt77ZMkW0NVx+D6hk6sup/k211p+pk2D0
+TyFmRNBcS8H1syqnKJIdSQs7EpBmfee74VNvozRZRKFyw/Z5llHb4XDnSTCKj8g
0RnYlDnLHhvKxFVE10P90imDUsS1Op+YFM8nxNslpo/PJ9D5JNqNJY9XUpkdOK8y
Grwh+NAG0ZLXHtprnoRGSGc/Zeqzrke9hfj92zu4YVZRv/UPssm9xFUU7e8e7C50
DPbIFtjTrHHR7kBgs1/5iLG76IxxqoNrkVN0ASfKlqrz/Ayy97QfWA0ux0JQDfdA
FTVRiUudOuLBChqwKQR1KoPA8ZpmiD2u9pJHieO+9WQUcOSClz4MgD+KTYzEcjUX
Ha10Jsk4kVg4rp7tWb3nkB4OjCfDJ2FsGtVWjlbYPRY6+EDPZW25kCPSM50OcmbH
3FLhStjdf6pLUQ6n/TThfM2obC8xL/QWJKE+HjvghCWxi2WE5rTuI7DVbsSPWUcC
wq6j2BPTWcI/lyjN9RakHdnnVDyUc5IVpF1aSJbkh9bxEjVGmTVk33zpKIQmcdDK
0kEZJu9SA1QvyfPLZ6SYd8OUOk2zjyiBkF4abaqjiQnUrOxfmhXjW3Gak+MkYjYu
0st+ZhhpuXR2h6Lv24yPguoHz5nXxlCGrSrQppCi+6vuho4KruloooLNQcDpiGqw
KK6t8ZBw6WG0cbWI7gJFWHsImP/BzMCbiOtFkanz71XJ8ymfp6d7y/nfZglVxMRf
vuQMohisoKqOI8SnVXkMEHpZdbCC6uZEz73h4TIcyEzz8Rq+0RumZMqOKCrEzxuI
ne8vpDXAflJBmu+6eQCiZh405UYSt0KOSAF41tVM+mJjyVe77YeofR/ra3OQ51Jk
9RGeSRAeqfWHfgmqkG/3ZkHjiv68O0Toj/2zCNbD435O1hGBJzADqrS0HHFXPpbj
fc0+gCkB3hxMqzvghh7ldBXH5pgVRKlBBhP7ETN/HRiG2hyrpaZ/cMtHxOkB2i+U
U/RieDy0KX8uoemyKbigeUa/CJoCahfp7KIQ2sdjIztz5FoEH2zyzF9FdwQ2+hNb
lWFBiZozEi2rELHKNQdf1WKSpS8HzwusPOH5OG8a/Bf/PLr7dhmflzNaAS+FdEat
5RvvtrUEqT2CHpShzkfkY+c2bYniakWUPBNQzLWrO7VGOYPC5qBly5LXb1Gei9Sy
r/Hg73J6kJ0weNBZJ/FsrQpkpOHnPFZrxivZWfUc6uw6YBmFkzzQzDnJgA9HdBOD
Z6OzYApOKxfZffLHOHjSjHyXE00Q8IYs9AlCuRA5dq1ahwbhVUhx/Xn4I24lDQrD
x6w2HjtVAVSYkofm8jQ2Bcmvf846gWb6Tb5+M/XsEnT0VtMsCDHtvFEisjmhVlnF
7k+PqmQZmX57Q09kauUmZp9boFm7gzow/wEkNPohWwF5v7FtBVGeOK+vdgXVUNe5
+CpTnROb8/LAnQUMbjnUhhTyq2t/RgvQSDXu15Cmp/jnrqozU73vLM5AnwDkXMxf
bt7/q6zZ4jbbntSdREWE+Ln8ncRGo2ZoQ6h4Db/pcZe7WmrsIonb39AumZg4ti12
g/4FsM1WBcS0Ttz3qJwcQM68lsZ/QizTv79q/f+YOHdFHMtpBnPKgDyiu+dJLuoy
VpTQq7RNShwF6vaxhmGSDMO7Mp+NtbYI883Ow/s02U37SZSVT0t0OkWBDYaxprsi
0wlEBcUzQ8dHtwYJp/RrDHPGAOLYmXrkTsE0aSLtqLWpY99Feq8xsmWpwnQ+C2Lg
61cNyhdnwWkRoFirldMYJahGrFOk8fXg32M1EamEOzHwsbLIFgwcSsc5oceCCPRD
42mB5eWALE2QUsXegv3CVy4TR4XKtom4KSkP7JjlasA4bnVmOZ63/QVjLtMP/hf0
hrZ9+I+VMte5Z8eAVhb+HPmSgDJsOMQI8tvCWdSa22ru3XFMuUoMagRl4qAgMlKP
Y9POI14lAIUJeauOyrY6f+YYhxlVMprlBI2QhdeBUcqD+M8BJAXnucXxpgdJqif+
2WusitfQHjkwWzHZuVtaYhJWLYt8/XH3r9dchE91P1yqinN1pXRBVHv8ondUIgzY
5qnK8+ux9Fl/3o4xxO941Evh6hkcSWzEQxm1qEUl+3dcczX6kaxe7mFDwlMs0mOR
k/6qkM7drAVdA+vp0dIu9FALLKVUCUUm4mG4eZacJAsoo80J6dP3RsfT45MMoSjV
5j6rlREhQew5p0EZ9T/kfl4lqSb2cWq8kUlfc5MMCPmxccOgBGkhDQMrzf2B9mUE
/GFLScx6CecyxAdRSefoEdXzCRM/BCmvJKWVGmC/XYtI/i+hUzuyteBwWTncIJOS
zuPN5qHN2jNANMHhMp6fcFaAaDX4botUyaIafL8DCj+f9vrdrLgV9yNwo+Gp0ND0
cNlSpOkJDxqDo/V5f8RSyCkJABhhegDh1i8nOCbtGkdN5bwgYg0C6vYiIFE4o3UB
Xdz/2zYckFo03oLRUTsQ3jpiyrmIJw8c6VyBC6i0BxkHtO9ydjAT/vRqnFuRV+hL
3YzSYXLOk0wdTvk60rBdE1goo7091zCFSAerAq4ZLZHAX3acPD1x4z2j509b+Y2g
4agiXq/Ln06bN31BsuT/JP83YL7UyoLyDuOvv0NjWidYqvjndgFQBslEIQhFTbI4
H9Y2gl2q6eoQhy8QQsBxe3+diNNHHM5HeZ6EPjqjadhAFwnTpGKT+pZmwopQSu9D
jOt+fuqVMipejJT1lFLKM5o4MFneU5SINiYWFrjo3UQ77oGPEgYjoy48XbVuX0vE
V//Ev7Lr3kyX2RbysnRq1WUdqu3TywlVlndBlP50PzK/CeR/kAj7jxMu6N6VbDff
dABZOHy9qi6Squ0tR7FNfXfIoLvHricJFZV77sesMrokuiMufUW0hCzR1ksncivv
RlT53wBNfF6WVb0Kc/Ab+rg4TU1JYO5V80QdgRcKAhUHTIxkta5jOCvo+z0s/0cJ
7MG3FzqtKW2Whm39dWYbm7Nwvz9hkIhf/HvNvdIhSrn6+BcFGlHBZfJmLT5XzL9f
rO3cNzsahyu37I/9jlEBNV+xL9yzmtR68WNIuyssFUaHDz7NjtGDxgLZ7LhYS8HQ
9Lmd1/I66mnhTMXo+5k0UHrvG80N6ZCeaXjhCRzsLyLu2SbGV66EoEh8RtzCYZCc
ybdno6yDlccLBLGPT51lGcnju+vGrU/pSWBp2MaeZ9VLVweKX+XiWfpfgljO8ztC
oxz81RuocIsxb1QQsrkD2I8WfpaNj+RZs55PbQ+rZqE86lWooC9hVeqfex8ISJqX
gxHjmS/vHi0n83uK8nmwd0czfu0bhXLhly6Kc1itSOBE1757dSNmotsEqqPBMPBH
iiIN/80W4DisKeSDd1T9Mf4HqjXvfMTkylutJ01zXpJgc8nwKjDPSylGG0aadhOx
1nXxIAv5pJ3m7bZbQDajQPLmAWtsnKHzFqC8PybflHYGaS8qaMKAoJ7OA4RIcagH
OSUvHzi+GQnJcwMf1jD6wBeseCHHbwvNZoIja/j3VzaiqYKHsNlVCGSChF3sz1Mz
9Va/IpSj8ac5LztHkbK4YtJ160buhouVdad0jKzCTl9zW9o6w/Ss/u3WoCtpFcTb
ieenaZt11dE2klzAT74gXaOpCEFLj429sR8C2ElX6/JgRRPd+mSjDi3daKmHfLHT
iQ0SAIrnA15rFyElnABLxCksmg5/cNJSAluBaODm7ikvrC8tgrDdgyYw9vtjicsA
dytovWH36aWpYLhFQaahXiE6mKTtWVei/xXBItWWKhfMa0KWaBFzl8qDq3m+qElv
8yYp/bVBei7a6tUDwq5W9UcA4BkGyTvhKvVIE5h5YeIEMQUOQVi8PAqCC8IOcQ8M
k5BhCgA7siJ5cPdkQoKAlPGXZ4hdpUk/y+Wo6N6jlF4uWKjP41CQi5ILFh8c2/VT
5T7fAhoE6kRRZKAAWDgdq4OE1MW6bwTJkrX2RW4ejPkTBRdPvGsD46EBEphUDPgD
J6yK6Ohlgv0KwIrjYWtmnPbu4nCKJf6gv7cJJ3VTDr1SA7M56hkZcBtdR3VCDMPw
ke85SWso4myjHnWqEzrMujxSFMtp+mZmMUl1fTx03fhi232ak0OBfKxcVTRPnXf+
U0xZsLvBES3/Or4AieBeZGcmRKN1VWFM+uxBBAssciWEM1byb6YN4+gobkjjn2e1
IZa0RGuk8loxLJ033WnUcUElKPfxgSNpeZq+dsHT9PJPgzmUxwvVuoaEnuOZJqHO
s35MCIGwTkzOobIQfPlxfCfe1B0ntB6b0IsVhHRGaeJGERwWJBsmkYDUlGbIERmA
s1K5tKrAnYWl4D5X2dyJ5EqK5CNAFbJoTqHdj31TQEHK3DGLo5iFCKt6JDwqiYD4
kql755Ldf2SL9fjY2Mmn5B7hggpIbg0QWW75BRDFNNMgRNpLMJxralTax80i5uYB
NN4FE8TvuaWLdyt3+sAuiKWe+OHsERW+OPjgMh49JpKEZM4ZFHaFDjqX9/Hd2GSi
aRpEzHwo6PLxH/HcxMxbKWV8JnmDiHc3N1YQB1AZs72x0xxVmduPJz1sHLgYwADA
wVtc2CEVYQ/ElNFmblSQerEKFiurNRb+uKtVodFEsChQ26icfe92XJmjAx2kyAUx
VK3nSLm3CLbitMTcyPeexBowrBXxjRVsQFs0I+tLYdF/mitmiSSbFbuTlMQ764eD
xyxH4RRiN2nSckD3aVQMszvtYB+hX2mnVysXsyF+tfslnXF0xVbNHQ812o3/nVar
FPSFwuVWNe8XBsVsr12mPjmJFvZGD0jE49/NLWxtNwzBy/zSTkv5LX+aR3hM4RI5
fY0Wt/K7r8FaiCkxknbpi5VI0Gsv1btNrX5VLxNcZbW3jDSoCiCdpl3Xr11c/OZh
Gw3kKOX34FxbjNFJVHWutXFR/IUSXN/tMaV3kni02rlXLdxx8NZxcb9zqQ9mXhf8
PKYpMgAo/9o0O+u20naanrsbucy7Li7Px3pnZYM9YaRmE8dojG1S0z6uz6etmdlX
iOMhtzfANEnQasUD51Ru3OhQMeTMZxtJTu3iKfeDx2J1YkeHmpfbuc+PnJZRQO4m
3zrbsjlImQoN3HoKO6a9PosccD/vjNfQ5pGAK3Nu9bkOpJgkVkb0/FaTE3HPtXHd
OuDXM3jfOLpVkDZW0ShCjtpPOYWQOYX2EuCSCV5kgkdPlwrfEw8Yo9zoJDIWXZN6
t6xfNKt91f1V+oMdXmlGdh5MxdjimYuMlEGT40tLjrmS8RYhpSB/Mh0t71462avN
n1hmMY76h5EL1y7K4gQwYg/3mzfxyVlt52iq/qKBKGwgsylKwJUtZGkyV4nHaL6Y
Hkk5j+hE3v8v0Pqtv9m5yjmhXVauz0bm9xUD6J2QM9eQwzTb98Mzal1CT+Kuuis9
+C3JyBwG1Slu4bzvGIPXsWit5HGjH17I93lsn4oSLy+nSjZE/891RwZWLYmtmeo8
NWWKEwoVdAxyIaLIAMM/p1+boIBYsjA77p0VqkSgxA5hxbxr9ApwN6MKUAIJovJr
czUeEfaZuZ+OV4r4Z8MLKcIPzxM8zdIaKx591EiBP5vt9NeBmTA84RR/m9DDznr2
+hc29W2Gy4cVPUvQlQlYS8dQdw0FEWPecOmy2YDKCcAPh49JCKPa9yPiklEwZtU0
4+wxOGi9xfy0g2w6CMMC2WfwNfC7ItPugDLgLLjo4ljR52H/fOB3mTIKOLRmEJgs
SoQ7Oo9SrVkoXepSSxF9LIi8D7aHxtK1NBVh0euNMKFhZY0M3ve1TOkiFNM3gTNS
sXUcC5U265oxwHHtwhIeaGS8c7hl/Khb1f6v2TvJusFU5OBspAMLdOp0NqDZb+uq
YAxa97Qt7CZgG7/TS84sncAzpqVQW7qPUfgn4EF8kVoXqNOvEuwv2mu7cF7UexZK
3Ik8MPQHs646TOZ5aGkUDb3TnPtEGjvpwMdgUfi7GMT3in20Y1PsLiydMwtcBhLs
CGmTYEVTK8P17QRdlNEpFtQI3K3TWxvBUYvv5kUcawPsLnQri1skl0g4tklG5zmc
SZLBtEfEqgyJ9lVrwuJK92v+PvOZIPMvlmbG+QjwaynsQy2yRvqT56dABcSDbR5D
5v4VMCDXjfW2RIzt58l1jM1aO0X+wbSsyzfJBr6t57Wl5StDbxJh6B6fpKK0sx6e
/79ts9ZpTB/0tARNEow1RKW3ubcWqvtfeGA8WSqXH3EACi9+4fJKmJ4WvCCZnw3e
rQ2KJlkbmSuehwGChrRfFTegT+VXCV8JzXl1n0BMd38Sa7FRmRMKq1f+FcQ0UGRd
xxU5QSvoiNjFU0L89SIxKYjRFUtj3/tscJ/bON8gBQ3gl5UMubrbLNBfC7QcT3BG
aV14ro7Jrv7b7bVQYY7QiWOneaHUi2zAgJ1HKgAY0aQ6W6XpfxgqFnpSmorIqRya
IZ51vgQfzBgHzFDoR18w3DdJTT+YDu+g4wWKoVTp+IknryHGenlbkrpR6hpzYwEJ
snLmLEK5T5s9/hk1J1N6n+i1DUAm1o4rto0wG8GBFvRyhOme10M29Fts1FoXJ2AW
VmwQbJAycvjg6Pk+i5Dr6A+VuIw8dtMDzidgr8D6jAWa9CMgrGm+ZO7T9gOtUZGN
d9lBaJTReNZe23fQWlgrrc+XDMZi+xNoDw54yUn0xWKGgpsuqPZXbCBhCR66umaX
YCl3K+vc4EDF2F2vQKTbekCxqP2lTsoP8iQnzMNlDIZRNzx8NBbM5kz0grrRmD9y
zuOVilGNjLnnaA2i77tnqI/pfnyJQr5zW2RIYT8N3vQlnOZ7MlTJ/KoSq+/DKAui
BdjlQWGwsjrTcivxQQR3SvASuj1Jv73SYAaAITuXFd5DLT2HRT7jG2Y4SPgiausS
lsT2XVRGxm3ej2EfrCHJkH3SVVej0TgbxgAVyq0dSWnhn70DovwrtunyDbGq1CaN
T8pRHJvBbE5y8IXfUd33doFf1tR0sM1BUGLqQNdJu7txqsEw1uGmkhg4zQjupsjM
FPl6xBlRCx5TVeO9gAkyZ8NTMF83oL8RGN2+6v/gW7dd8rQKFptQ7kjfstoBtcUw
INHsov/WW4jn9pIevqZ2CNxgQzJUzAdSrAjKSVcBQ0N1HXKGic4V2Lwo+MS80kBN
Znlp3ZEf3DbaGT6MJwYQjKmca8ovffWDWhxTNQIMu39rqSiezjZdkMYCkcn+Nw/V
10YCbvuFtlH0jn6+U1Wy8WdqXy1XpE4g/CDlPRDbLm0OcERsoU7bmXHOe5rWLffQ
+j7q2sYZexJnlLP2jn32zYW5IiODSyfdZDcWeRNA2vSSoY2r2gKpFEZQz6rAz2VW
/ni1nOA98yebw7AmAkTGoq9PH8CHmrCPPxkq++W07CcZxi88OP4IoClm8wm5oASI
XWa7F7AIsvYw+F1DoDTs1z6IxnohbmkoeV2bH9LLy2LwiCBO0h+HeYveUMSDUPcn
Up/mbLprjB4oL4q+irAV1lvSyXWCkzy2PkIipjJK3IIJDZEXOM624yylKejrCVFU
tX+SWc+13hYFMIzKBhe9rgcKZu2m5WqCOySpahaacO42QGmsiv13wN4ydLS32XmV
YV7iY6cBNaYHsIwbHO9zbOIYiNg4HGFJuDwqoNm477FY+ZlrfRC1VoK+dpfzsNOe
ZSVQG+i8FZ7KV1pO3zoVqyjP4f6Nk+X+swtqmwkvhjQycTP7YpWQX2z2RSSKpz/i
iK4vuNxejPD3qH7FyA+jfoo5angliwWQK/p2e3kVX3GlhvepJQuJTCFnuJ4J9E36
DeGQjmrwJnKbLyXhb7VRmHCwc6sHAxk6Y7Zif5igwWRlShTi3RiveNNraWiaKPsK
F4YRchI+o3jJIME6ftbK5MN45T6kWjMX/PIIStwaoo+Oyzo7jx9GJlD4ud85/Qf0
1BhM0XgxZ7i+ABTvaE2FrVAohwOUFYddJqZE/NBuvdLO9a0mC9mmhOhiCXZo9Sag
74UriZUn3nmWTY5AAQDZ22UF1UdPwJ8khFnEhSmso/50DAPPgVRvNtquphmFY+lh
Dv0fxJMmlCPXpTeOvsxOBx/1KEbvfpHSJWGdBHA6d1i/igocu7AIRd+GFGHogmCy
zTQNd5pQaZj+ZGN3+3+DwOHRxmo1LaHR2uWyOa+FmZiZOuApaAWrCPSGheEOzXgA
ZbDD8sCR6rxHLZlqNaDlXPs4HYm3e5qmrkB6ggua+v1WoH8fvgJ0TVn5673krwyy
BCpNPeH9Hqszt+x0FL43Id/MtlMNyyHAIsmDhcHaPSO/xJWM/I+9ezICNmbcmf9z
VgTcAmFC1oXSKtZJ72URbpI+7cHH8ZbaRPpfOxgjk7TOlu88dQe46vgfmo80GNE8
PQuakXFlOFPoUqgM2tdd0RFaO8oYLwQppUubqqyZAuNh+oix7iUSJuytowunRsS+
07d+Yr/sG74Wp4/kq60pbnyWCfpzPkUqLhBAYXZFekc/N9tUuTdeeHZ0sMAVTToM
F2t441h6ShkgIb2158gvGKmjvnWb3S/bvTotgiIePy4HYN+dk51WgWEbnEg0+cpQ
sR+CRjPhId9qvs3UDadnKCTDXBgjF0dPUnnUG5ZzO0/yGyEf/j/M7p6d0iUryJsG
RTxw1txRrXFCeJ3kGx5eRkVuoPzYpl6Qutj2Z3pXxxplgWPnMjkoCXfyEAQU54Ro
De6S8Rv8yBfAYkNHaCJip0b8hWGj8iNcpl7AjYyYVJQK0uZLwRA+VqqEeXj5kI02
IO+TDzFCKueFJ1k+FXuER+m03rV5T4kN+BcxCzA5YCSjLMcLAaAcp9J+QYPm4ArM
OOz4Wbau1H4/fQKSRVjH068+dqPh1bC70tFk1qXhS78ppIUZP9yrsQxsxwiHGcYE
3eZcy506MwH1Onlt8aESj2K0QcPbg36OK2tiKsjP7HfiCopjdDV4K7o5hhkeCesi
jlSh+LaPTl20F4QkQnTbnZAr2Z4mQIe1CeAxHTuX1MJh9z2UQYsXq9sA3INoOpyj
mK7W2c9Y+h3HOvkziqQVflgMg2akd+rElBE/Kfs8D4x6w3laClOf0COEOAwWh7pz
NBK/ge0UeVYP6EU8o+cPRjmGFmRtkHDbkSRYU5UAgjwEk1IoLcpYLfpWjz1VuV38
UTfp+8tJGcxOLF+EaH8ZgMrGW/Ifl/iUEH7s0w4rNMqgWprh3ilcPdmaiG2nVLRH
/6Dh9AFkC5/V3m0i/JYIvvhXksd9T+tGYuXfOH048DvImiyu3ciXKqjSH1qf3Yti
hGkOVt1oerCgKCTj2jxKL0rXr5mgDW0OhdUuhRQI0L5iKJd68o04b9DQ5fvwwNvM
B+4NhO1b7TKp7Z7JHLDkZwiOV03AYYL7v4x/BsNR6cqHxDdlJ7EhP3m2uBGczYkW
hsRCxbeh09UPTXSRHBqin35PFy2AiXnRKh8jskjy2fUU+eg+BgI6EijbvmFl1ddq
DsLLNbJeRD/NfHmpSn7JiyfaQVQ2UafWOJGpsnDhlF1gI1s7lzZ7pniT+Ys7AQCL
8Irj7L2pdGONMew2i26dDUIIBE+lN3bISpwUgDzabtfVn/Y2sdEmK4vrizwPk6Ax
YgWVdZBNBWBTgQ3mYBT+cACRSDn/e3M2gREQmHbf+vO+3Yve4N1f6L1UhJOO+wSn
hxfEh4vvJlmPzOzFOSs0RX/sOX5wEag4+0IxaT52A8Un5MN0RBlgoN9wsPK/DpfQ
+rRfy9LDfcZHTkIJEb7fq9nl6f21jEK5AMdAmVlUffnWRlKoesDDRqLnaY0r38va
t7HCQLTC5eHsP7j3u0A4/8sIcLQwurBXjgE/vUFOYqWCT2U7KGNRgviVoncGZpQg
plGAtDNlw9MZFPUm1nEoyg7jyKQCCOXyMQS3D93cIWjQSwZZemsgJe5sosyagFzZ
ZbOlMjb/GqpWMWRxq7KrkoiKQhT+63WZ1LBHeOB7OxnnrXfu0k+Fup0RYjoqNp11
OtswRXdwkfPrE2QnuUuMUtf03bnKPYl0Lb/x73SkW4e67tViHNClt1ZgOfc+UG5P
uX7qEJ27ExGSxN72BghNxa3TOx3Uo+mRIgKEuJCvM+zhA2t91Q/SeKpiCgLGl8xO
pa8NDVZAASUNfI9G0D9nTLCG5UwrTZLhFioIdwMmTLsiKLLQwcph8easmZTuamiS
mD1dbSnAJu63hLzs+gpah+ajVKS0rGWA98tMo1zXCzmewiM89mXdXPTb9oTRetvO
A40whavREkHXPC3sdbWZo2ccrD8zA07n7NGN6yQ9SO/tP1WgoVCV7KDkHckL8SeX
A9jQW9ZcCX5jarXRcOJco4CqyrTtH8vziwU8SyWPX8XjKargYGm/jVo6+sfAK69O
D/SQy6YGPyoEj8ItaT6AOjSosgnh3dD0sfmD5yzAOmU0tIHSWpqylC9cYNpqUHCm
6L3Yd+AUuGRrI/XWoIIKYUyexUORDaOdOLsPvOfvZ2vmhn/gA2sszhS9IVuxWRH6
Rf+4tsRh0YlHB+CvXcLT1CBhJe7uNZB5D0dRo7JN+XlMta0Gz+L22a19B+dhYSc4
cZn1yoa4fTFeBykca9fXqHwONXKk9YGtHdI0mrKDIgCUWEhsYtfw7FZObWA38Dsv
XZQv8WKsTzrdnAC/Zo00Ca6s+apHUQ2pZRLKkqZBqbfo34WBXrAJo81SOvZclqLe
t+/H5mIG5512LwiPvyq/jNdsThcdplgAP0cMebUyBoI1Yilf5K7JBgcpaK4v0coG
OPX5m+QUfehtjCM+Ty4uwvFwgMVDxwVqfao6HU7pX5IdOUqpOUX4/PgFtuKogurj
xxVBW5wmqDK1EHVZzResozHt6Cbz1dhltlbD0wzCNFbQ8SDAP4nNM0n9k2X9+25W
LIKvhmwvh4TRX+rrrLhCnNtCocPIwCT6mGCwwH1epRQXHzZZpv3zhS8Mq0aLPETZ
g3yuph3AlkpupOQPlfqWavnX7tw4ulJJnZiv1QY0gQaBCbV3nWp2NlhpklEWPYKw
38qM5Y+bTjP5Eg4DymmDkxj1vFBKCGcNgEgUVHs4VxRtbTO1OfD+TA51s1kwQXV4
kPNDjiLakfaJsHXTZNl7Nrz+9y8oLYdG3vv614bVoxgA7uDo6xMdkwg61iy9bOTb
QLrc58u2QmSiKmssz6SfYhZ2V83zM4qoFF3XPg31hq39egXwcrV4nefW5M0rroXs
Uxyh1NU096CPrYHyV3jAax/ifcyK4/DgLjuf9iLOy+RwOdtXHLMf/ZtTL/qyI8ve
L2R+winzUQPSrPHiu5Seig9TB5cKYAGoixdFE9E3jcanky495NUTs0ctQtKnCKhb
jaBJ97x/MRC34woWj3gWO8Q7tc3baqUE8DnobsMji19P0JcR1pFRKk15H5I2pe+J
F5Uau9ODTQXVHKcJImXceByQeV04qrmrJDavU9SBrk4YYNtTAdvRIT2PPF95P2mV
pNu1pivASZF3KiZpMDlkWfDR/bZlsivRc1PBvB5rTlXR1UqcC74kR0PINzmN9B0c
8afH3W3n5ANo0o4B3OwyuMGapg9Rk9Ve1Y940cg8FHawEDXXKZPvdHPX2MhtMJg8
lc6mJBHv575pNH99TRe4Ko+8wYw4Q2RcpRKanBHK4Qoz7XY6ydwy8DFP/ZLQXz1E
qkvprcLxtJNXQ4QtjRVHPwakILCY2vMcOM9th+VQtgSmDOD6l51k9c/Op0TqKuP4
pxnlRuwSm71VlmNHLSjelmbhfT8i8NiyQHLpCgF46d5510T2dVaK8BcBg4ym/M89
0/UfNrjCJDZd0mhxnEkMQHKe2hG0QYesKACpnQ+7wRpGQqrJUv227U7k/dqPfnYu
mvBuJlE78GOHfpXEpp7wiLQX5F9l/OtBEjzSnPxOKNg62rnQ0Y7pnL6G6dCctyGS
e7z4t61BkkJlLtE4fsWRiuvoWCpv7fEQHkHfb2dRkvgsAUk3VteCDA+l5cgv7Z5V
48IWrew9lxtTP5Kz6aTwBeZymWrOr1ZFln6L0Y7yRsxnnMWLLGYmIUdHo8HweV7O
VwA1azYBiDiMcG25kL5JYHgSjDvwkxGBtHDPSj+tL+s267PKuCQEYxz5bKswxcy7
uVV4T5P4d1VRAiAz+QyKqSzTvHjl4RoSZXaQidCe0k58EfdMj+mjnEt9vazYK4c1
2xqhcLTjaw16R+b8rIZ8QosEcRSDfIcsW9ITtqwb/jp7p1n7YEe2jdRneluMAc2G
E2K+Eb/he1tRcQpZVqpxCEl+UDAMVimzoszZ3oHPr70l9Qn4DHWg0Q0mNBsiTmmb
crx9frQmr01A3urJE9sGAjxsaf3pBwRHprR3h/oeFIrhZXIruFWEtWLoA34jDStB
+XiNjs1cR5ieWlYB0n1m03QnVwaOIkiP50WmSnI/1fSihDovwY6nAMrstOZGcs58
GWk5Q9Ri4mtkltpzfF+XGaoA1IQjLW6BOVgFPyz9xrHX23ZR5Cy3UgyRUbH20ze5
9j+KuWBLSNHmwO792fuVK6+vynqcSwrIdS6mKJRK80nPn8QdTcdc8E/Oa2RuCs7v
21M0UhCY+65UqqB8Vt4aB4r5jBfWLOoW+CujB2wiSLDsvEIgBfvE/a8O28eoKlRb
uCx8LNP6+0d5lBW/3urDCOJ2JdSwegX+30iN7xNeSIO48gSsJEfvXWriJvhqi5VY
HwZ/KGXTq9pq2hvbx/pC5Bd7RQhHj2346eTHXknVbGUwycDrMVm8vOJ8EopN5YJD
r+W3O/yeldCEUrOS76Lanux0azhLGg325z7k777tjC8iy2i77IkZAY4SnbImPw4O
Z5S8jx2aNLKBh+uEqM+IEXG9+zpW7gqAEm8xoiOo6k+0lj56qdneBhBzN2NT7hXu
hcXXbyYV6apqF2FD4BogED9cBvny2GO1IXZ1FGRBxzdcGdKITzzXbsnrlblw5qHS
bAsmZXbOMK/eYs8D9OP5Q4x9r9F2+ucy6U/xvDJoY4lX7Q7vj/0CD7wwAb+v8N1m
YuYG3vXbjTryU7d8619Yz/f68RcfqSURflPqOcZ4NMr+H3Kt3fN567xtNqTjMu1w
JXO6wNeT0s8wbhgpVFjlqntHECCfGGAnCZrP81TZ0i5SM/Zjltc1aRzXdTz316nf
IqoPSEeLlTfBUSUERwvqy9X+6ehcDMyqG3LS7Mn1E4tbWquRX3Q6iNacRzfJRxyx
tivWaXJ95pew0OHDLb66vQeyiWJ2tFJt3xB37GfoTvzxmgAOll7RPnqs/3/snLa2
rBWOv10hR0ZR6WKV5hxRwn1VE1NC+/0lVMNWuw+A74fpA8hSFuyv4N5SWhiKgbG6
2ohyWY1ozqC2aKInvReAK1FQwtAFraPS1zjBjivZdWIYfuZlpxKIh40JyrjZdKy6
X9NvmM7rXFf6XuFU7vKYIEbcGmmapwOtiLZVPT5z+zI7ToPUBEQN4gqzaag/cLGr
T1erD/QmozVn3ngihEGVsfHBb97S1eQFNuxK+cbwlV+2BxWYDkgFRvLScJptISuP
NgvlTSZJ+MExUq2zLCZDYDjarCJvNYKSJFhq1EO0GcoJvG/WsgyGM7pZCn4t8/Am
OpTKxMGX/TVTfKlGum8K9941W6vPmQj1PZ+GsuFaYtdqQp1V7pPdJKV5KteJo0/k
pcbwHUzaj/05UFHELc+0+NfNgboknOf4zsav/l4mRmuPUse0kN2Nf9xkEiC6IAr0
VTSJlmnYX099DThh5kxwuFjGyvuz8RlQw4/3/XUc1MKFC0eU/oSwbKrazxw/wUuJ
eShFc8bd3cLsLdlCaBc9Omq2sec6yAX8UNIUTKPrjUDwdHJbP1Zot8nlI3IVQaiu
t+//TFHwoYWM0tdRbZXMp+AVxJNKVnc1j7YXLwYkAqPjnD9jMkiYucsEsBuJHCPr
sA88q1uzCeHD841MBS0E3kf1hpGG7A1rz4FSG2xEOnBT/snHMzrp6uOfpodxwUWx
k6t605pUYV35Rdme/veIDkakN5WgX3ov/7dPcVbyiDoCM4TFh/JH5UMBikn3PL50
lmcJlWBPsGNqsaohw5W/3SsCeksCAgICVOZGSIDrMHC1rV+TkDv+bORNcUx/NPgN
SNLr8UFtkfLreYltG5kAu5U1K3S4mGs8+sVYBZcmckoofuwrvGX7ehfT0+fCrNdM
+SseM3teC2In8SErLEl/Rusvg9mzP02QmAkHZKyJShRdbIshgZWuENUNKJgtnnxg
ouDaFklKETYombCD6eVQJ4lgEiPLExCaG5UEg+na/+lAqa62/i6qzJB2VAoNlD4O
8D637NnaHV8vSB8VQoxUcgq2aaW5+0BNM73dd8Y74rzOGn73jOJ9F3Re4xmqRo97
GIPuidb41ZVxNLaGVeQF7tmlT1qr6Md4FiWwX8Q7Rl6UAHCk5r9cFmKb24Dwn8Ii
BJf4E5NqOXP9//qtMRCDTVg8N/jAXiMB2rn9D4edu2Kf3bPTrZRPQ1PfwyqKvdDh
PCwl7VDs/Wp0rcvR1kb14XDSyBw5h299iB/Si7c9GeWMShms04ymtIQa5a1Hbs9x
kBgVQ2VysiGRue5kOQEZOMSG+1SthqQU5GrDSEOfYiXB5SuVjnlbLRiGF58IwTbs
4vkeaGWaLR0Xx7cILYMpZ1pFF4TwlwUFvHeDyAxyL5dyIU927NQjA1wINeKuIzJB
4HQPRUqqV01ZK1PrcrsAgf+T1QGuX2t2xPoZhn+8Y5/I0uTSg3FHAfW9GjwtiNxW
ZFSyLRIQQt/rI6RREnupcK4T5IStfR0SsD6A6pJ3F1mY2vauGGvOVa1EvQgrAYuo
0fWIK5zvhJD5Jsnpi6j89JS0TvHmNHBQGkkhijilAQu5A4xx/7ELhEvVkopK4GL1
HJCFGfkvZTgt6G73wl9ICXyyfJE3oYIKZjv/cvz7VQdkabA3/Nv1Hl1PCuF442Ak
r/JSur1h+LarVeQ0O/i9FTfoHc+6B98/hN9pbFxRg2ud7QPdyHmsTjBv/kPm3Kd5
vhLVggL3ouA3phwfM46iuwjOGFFiYEYcOoUT6sUfFkPQm0E7zukFiISH/2591Kmc
N2mlFIOwTBGA54g5V4GXm6p2wN0WFPyMRXFwEdBZZ2aoNmP2Py30ON7rwollLjEZ
mKGt8rMU6MDE61MvJ3d5rtnEeXSfx3Qr3Fom/jEVZdW+m51uyLskl/1ZwcWNuIkC
dvHWpKbFfdyQeP0wj/TQVraooLSTTwwHpBkybgZO6poPVqE/Cno8OGhtJe5tbPIj
l8KNk85rab8W07vZrP0IkPAUuspy1OfaHlJH7kLuREw6ybwBENuITLy75I7FgAdv
G4vVyg9F3PqbA60P386AnitukL7FGUh6wduLV0nIG7N0FU2Y67mkAzrOL8z0mP1I
SV/nOCQmzOF4vb6omHoF4cmdtQboLkBmwZhF3AzQzpoSg0ne5Kv+LRUaINU000Vw
u8eB0no/Zu2JN0huXSTnGnP3K0oc+Cii/6VYTNxnkEvLtLkl9f4nHL1RGH/YVuRE
IwPZmcDFDQN8D1Z52XbbP9TfE1lMYLOnjcuJD6rJauwhDGy4TBLRDOHMeYjFvu06
wOXyVriNDjvuR6iBluTt4MYM3SRMGfxaJ2DyEamrDwONIojPzHKQcJf/g0nWgNiq
B3iOt5k4q2fqzwWroNTZoeVFC5Zxnn7KwaINfG1bgnw=
`pragma protect end_protected
