// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:56 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
KdXXFK1OdhWsvi2D8kbfVCkHb5p7Rt1MCi38ciGjRs32V3/HxLaQLOkJLA4j9VFN
Hbeyhb4++74mGfVkugZOXP0qqNDVoTzT0wYI+XxTO9GX0ZIaZzfRwrFT4hJmNVjM
Zs/8Q1TBy7g9GA5zkthZDRC2ApLSMpNeVebgXg90Als=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5200)
fLnca8OO2qELYFiZxjHI8dsNtSF8wxNknamh+4ybGs8S3f6JYEgecYHgRVOyVoZn
+AMX32o4fso0EPPAuMe3kaMRfdBfSoruu8n0HuXnyrMVqbFGSdhqrjNBwQBakmvd
DFzP4SsWCo5fclmXNNhvvWL632CMrOL2RU8z6LpwrWxmq2x+BF9oK7t8fkTnXdnC
vZRDhhbNFEnHoyCifHwqL0UOE2tGbRz9YREJLzcpKJbsfzqCDLoE/qLhku/AWE7Y
mlzE41filuUFsq299Ct4NI5cFa6CZwgL+v2yFHkncn2NEH26XkIVQCe7SgFaw8hK
NsUCSbm8K8DakrwuNW2Zb7WdtPB18uhLDboAdF03YUomJ2tUaYcW0Q614vEqrE6t
aE7ByFtEQwcvscvqfAKums/emTo1EM0qTvMLWajR+SGMxVsyyHZckKTP2+uybrUw
oY5IUjiAyWJYd6yQgYsy4O/R0gDz1UJaYxdm/yo7BI+6f2a+nCLA2VElLWVYyCEl
ub8i1ItsqLAGNfqZx2aBLW1hjt2Xi68ea2HcsQqUusUu1mavhg28cccmiITn+DHv
r1SNDQEOGsTa4cjvUkpozvVTkqKKQ25kGAYWbXDRf1MqufnxRPFPzgB0VIJB9sGI
ECNfd69DluL1612AClKvYSjZ10g/elzl4+iOjyuf+x0CSdf/uZH72HeWr2hSUTct
P9SBzi25OeWjWoZYYKTUr8wq/VksF2YFE1MTfqY0J+cP7mLdbIXXSDpM+0g9Vf1Y
rwfSlP5AU+3FsTfZyV+fmXvRU8FTJOL+IIdJwguuNio6vOV/zknGThQeLhBpEQ/g
PqITFkKLFqrSxQUlgiePI5AUYT0KPPPpcXvDr272VqUyJPAfmSB6n2NYYpb6WHyT
CETsYsbAiVCl4vrFZSEIAg3cGO/fNgOaKUtLlbxUuWmJlY4AwruQy/sYbZ6PlEMt
u1QG/5RqVXPv25t+0M+fy2z3GNSgloc5rQ4JMDiQz33a2v4PwQa8YEyFSNI1RmKK
1Afmn1j645WubGihYt9DnZdhP5EIk7aOyT/ZxGSINHEbSRQxXDxGvwey7/lLdyYP
QVfAQv7KKFrZ58ay9gBuwc8BxI4d03TJvncFTYSoceOj660iOw/u/ugi4+eFJliP
/NI1eOdIOx8i+MbBcbcHWESZyTue3aVXaKwEQzkGQoE5u+hVgih9moGyZIQZbx+O
PeGW0mJ4ZVdOvH7HNHVR6RfWxvVKYDC43651glEd2t/4HtpC1gHOXD6Yo2iCyO4D
BlP+RDt4ultKvqRviz6qE4IX12EzsdOUU1Zu2B8Cx1QHkoqTDuUZ3yyq8ulFuS8b
TP0F9YpIsvJ47LbYplZ3MbJvXFt9R4ZwO6afR84M/lrNV6Spw7kXfhTLMRya4R4u
yNVc1NidjzYJeP4+Kt/yo5Y7txMCxXi7pLdNAYczlYBmygCNYq20XdHwaQQMa+Eu
ew1Ogx6Zyz4Pb/MMowaoa1e/Cl0FaL9SJV+3frclLr/wIAs3/KdX5fD1JVvQmbpa
W0BmkHCfiaqUsOeS31AoANdIfpNwOe/jEgOAYxM3tJU/Zed6T6JRIjx9OYzbzQjO
C4632h4JUpUlprhsqTwwRcl76XeN98OjtXRIa5vLCkEtH+8BlLG52ApJSMjhYZbU
aGdzb/ysQgCyEJSaiSl/qSdXuyxP3xL2wszXkv5wAo/Mbz2L6RaSuLJ0/JDeIvYN
zwzdvE62RBy//UkFcRAUM0vfc/5siLUTRRFltCLCaqhuRcbn3i22MJtJT37YG6k4
peP+DiUWCOPPpsAXEr9xPh9EfwoM+IVbOzradGMLlIV6FWBakJ7YEo5ZFP5CXE6i
Q7afp1k98JWcMN3QZfTvm2xnBr/mNldcepEPg8r7y4Au9SqBd9Eg+DcqbUn+Frn+
CStJvo15pYZrSxSEiidAAiJ0jXTHrTJdeKJLOEMzFU2lvyVV8pwuBJdF/EwYmxIv
d5EWazveLzBqCi3paaEyIngkQLYjbQhQeqeVzmaobYHazYXHhRSuh+tr3l59Ke7H
B9xxFJUQ0e1m6lxzNp7ciqebeRRXSE4aE1uQZgdmYJa/YUY6DWy3gCYC9IarMZGu
GH/X2fIiTSrow5ws3YJnkhK6+GWFoEoBhkDVg4t1G7w+HcK3nb4yTSSrkU/3WyIW
HkaQhYDvlXv5IO/g+zHu6O4AFKMyE7IQzq5V/AkBinIvsg5rIQ56YfvJJh/qEjOm
5KH11XcSset5TlC+7JZiIcArTykpcTAfD5UkpmoKtWw2SFZcKEB53l4dcxv8uqDy
tgQjDhskWH/j2pelPb5UUFWy7stYqsWR7ZcD2AbLvBT8ydRrts3h2bKNZ2SI79KN
iTPRBfr/Je2iBnQ8Cey7rMzXdtORg9/1187NYSgeaazs6oY0U/y2AVkooQmJ0zfz
FNX5rElV4uexoV7pyFtjiBPpIPT3hM4bsmKCY2SMX+faD//Wov1l/iNfbotP76D5
yQCcmOGCi9T2vdvmn4bPtt12/gRapn1nE3qVbkzotC1KGNzc+G5PmChTxQYKdUL2
8xnWwV/np0Ryyw2m8Ci5d8copOcauvJTpdzMaPDbg0+kVlHaG2Ee0TjOCG6yIDu2
cZJn1rAgW6icYjNq7CgpiO/e4E6lnnK1BLy1P/6H8yp3mYPLIeOoRpebHEnn23yz
eeH/zxmlsB+jltLGWB8QFM4ftjYSx6bv+9QTpwGgLYDVTL25PVAs51zvcAcBBjCu
OGH5Pex0Lx6Gl2CLsuWx+reB2v0Lz8P9Lf1ntXyw+p9yUwVdoNkXB30yX2nluYA3
IXlvci5EvVqfFTZEqAZqY7VtjuMAATz+uETIVtFNJzm1yx3kmaANFH3UEKO4RQ9s
m1Y3ZBDzloOhIEDhdiBF70AUJu5J8nOXvQKj1Qi4sldKP9wWRaGw4CCFN5dYslvj
o1mNENGxedL8TqgU6WFh3rYOL9SuYQ1XD7i6s93WgFUlsVM/pI7HbgyVJJScxfeC
Uq8T+A8g1G2oOaLBl+u/+YLzGLIkWbY5/ZG/SfdGyJYLx2ItRLdzRYqKCLuRFsB0
/cMvCeoICBTJbkx6BDIlc5AOjUPYk70QP3lPt6lXb5F1Vim3PQj7cS3sXoOc3Zrb
PJ2Y/BUHkbZxsORxwV7XIsA5DqnWcWyTApXCP70cUol1zLhRU7X0uLhk2cXgihoa
ITvBSls75AuBwNNU0+HV3oBI+cWU9Tn9uejqt3pXBACHWMm24BIGMOPmu9KG9pSw
tQGZwF2LpFFLSkmql6pj85zcHSbsjrQOdOgrUe9X/yr53uc4GNrk3wc5BbhLtWps
QeAHpiXEfmGdpNbiVwAXhDAKJF/OV471dAvnY599/OXIowxSf4zLYaNDXnxj3RlD
8uNSXZtkih2PPRkKkq1vjX9eThA+TwjP3LNFilufw7tXrABFjafZYUOkx4EVP6R5
a8Nwa9OiUFIwylq244G92a3Y08C1dFXOmKQhJOD/2a6wAuddPlHrIrJ+lPM32lJd
MjAMfFGf4R68L1Sv2JxyUwUenPYcKum59RH1Z/f8ub7j1Nh1KIycDcDuYSkfY+e0
gKAZcxplXbjrYRkwZUhXGesll7YTFbEyselqOKYyIISj0wXXbRaPZaZW8pzCxcBf
0WJzPFd69USaqNBrzKb3mGmYlJbiZfju7T8Bcsr7D6A9kxoNVP88WZ03Z55csPtb
FZVicMze06N5d4r/D1yiR1iTTJAOC0dyJMdqHxEh6mQs8gjJP/Z+1/gv4/8UoxYr
vb0DCHKU9M9EThLzVPOaFFD13UqjKn2UVcT95Y6BtwwnC3b0wEMQx6UwXWaJa3G6
LEoCclxf0qo1pNufwdmpRH3rdhKzxOSzhMmE6hG8WMpC+GtY9GpnwB4VKEMgaRog
/WBcwYlPKDWaVVgGk0HyVKZxivq5TaCbW0aTmVJUhJqAUGX0H09KgkH5ba8YYd6R
HU9+Nx/Vc8t0cVOev2kd0LuFlhMRysAZyvL9E39cAOlhY8Sfs2XTioBzGQFrAPik
J9UxSmCpMhNkVn3YValAaI5vojSd8/s5wLXdw4zN0PCjjarb6xW40xBuS7pgU31o
N5mUOyHWyovg7ol1lQtgh79I6QJ2doWw2n0uUVZ83bjXuQM7Uul6pHglQKKNgbXE
kkuE8oqAAM4PYYn54+csjBemq5P2fcWkKgOF/O20pkfxVIZW+ng6H/FVtFbk91A/
UKi4+vpvR2+yWMtmB3gbP9xGV982umqB2wzw8Z3oXScJNMfADLn78cfPnmYrUPwJ
BEZtZNDVUJshTUztGb/1VUJf5VK/brJ6n3gJ13y1fDj9kZwcmwKP8XYusJ88UQNH
vW8A24FZZnncQfgz0w9Is15dgDGr8hLlIQFiNGxiaVZwBRkkGY53a0I4WdD4uNU3
qWhUe5bMtQUmIkI5Cwhdw5EwIgpA3gRun6Yl0QD8v8OF/jR68aincK4JoaYmqmH1
VSGmBx9nMm9CXZm1mWiB718ZO9zQ0PD9uVTIBXuaKMXJPse4bITKsMDglet4YGcF
ZrBfldHXu6rxitRsoFvqgLc6/Nvlgqh+YVdaP5PffHb6jsdC2g6o39zbB3pfJxxR
7hjELiPV9sio8LoUcOAOrQAUlAzTcJdKXATXd5gzlLrp3VU2i7hdVmw0hp0zPt34
/e9d3AHWBXAQIf31wkHTYXTZ1eHMCqq7+ecWcnctp0R0K/sWxt4coQPSYMmGZF7U
edYaFi2Kw7GAOYlconIK0ZHHevGCL0ALMzSdIyQfJb6t6jzNgn9MPFMVu3/L0Xq0
vHHhZHApVYI0XwhsmFozIOf9NAbmN9nPexOjdXx2nuPaYVTVY42UZsc13aEYMqNd
wmwRtsZ6IR9PQPcO7+6duuzVlqLKfR2c9h3W3fk1xYEjkqVsCkdoxVoHhiY8od8c
kFymw3zJ8XX/Zw+vzYQPA78WUlB30+st32m0sgXQ+TU4Ce/If7Vx0vlAKSGgoXlj
RTYaXIYEFc6JARXNlB1hYFDdNF/F8LOeALeTGsOpJdLG0WHJgRR63mDUIQpUBHmu
m83ATjxmaffuW1V1Uhtn5btmg++Gxabt/oyS63ZquqSDzjkpkkV3I7/pvzBQNSMD
XTRLHGwKzfEbDNlKVY2/QJK+67/3yAjHljjv7zkyOuiJLUOhL5TXl4V5towr/9+n
sczvdT8snH0dF46dCzCg6xx3G8AcaN956F6mX9zX7KvQA5rZCukGdlhFbcQEkMoR
k8pyAREVY3gnIbC9dXCWmnKFECnvTmAfkYSOZYB5TjaduzxZotlEYRBaAlmuNZDy
QkR1bbH4wmDjTuT1BWKl02BPlm3IOCqD2qtLL+PHoi8mIilDZ3B51/KYxTsDjY7f
SFUWJA7XiJnjfYriZyAuxQgsS6e+inkVv7UUi3sQAW1cel+o8KZwR/vmBLyru9pC
bojoY92drsjKMxui57QoXJwAaKsnhSg1EBN+RiGJlrMofXlmGqBl4NuuwJ2WIByE
7ceDz4wcEoMRO7aiuW/i7jpCYhrtbsVvN11jwoXVJiyrEkr4UabSNoe9fmQMyDgx
B/uQyN6Eict9azpeVjIcpBLuws5UdR94mBGcEVgtdJWXcH5Vd40HoFmEDS4L7+bJ
s/lwn9VrEAqDROX77gfPOnCrNknOnMmD9cUE/Jyb9RRCfIPM5loeIHk68Pu18fsm
tWXw1kc3Y/imQa6uUrXZL+8YYqq0vh9E+GvY0FONE+q7wA0wG2h+VBQnXeXy/qa3
WJjlpVyNabf5sRljMIMLeYve2XpzU6A+G5tEEqm9naXgu1QjVwXNzOKyriC1RHz0
ZS2kL7AKwk/VUBDggIhI45rNJ1u1xanOg6Wefht8XQK+KfPmFSMDL2CQxw2APCr9
Mw6AA1a0pZYgf+OlHq2vszm1v1Q557qxWfpLwJAdAVvJc63vflhI5yaIq+lInq2m
VdFuz1j574Lq/2wVOd5a0K7FDscbOLUD0i8gt/k3pRnLSC5Eq8Lxj6JxzJ5YOvKn
pcCUiWwtFNWtpJ2XCy6dWfcLz//c5fsRZI8ZkdwRqG2xv+w1FqUWqNtRgl+gMKWT
ALTspzEI0ASmSTJj9LXY0eok5UyJbfoUfp+w42qVSCJrqSQXJssugNCBAu6xFrrW
zrPNQq/75MwaLSVmOms/3eaQ3Y4dUjbbzv22cSFkoJdIiK444w7I/Clzel4r0C4h
734g9vKxv3q1iX1TrdgEavEITh6AXWgtmNiMKYU6hA5kAm8U7Cwr/JhN18BlG+6s
fhMIRMqrrXq8TC3fzTR7dSMcjDluouGgleglo1CPcB9Y5Age11Rc9MSEqtKDOkkh
eHQRyZsz/PQMx7iPuyI1SKn36pNzmoP2C7VTpyrZTxfi36SmdFK85WoetLZPs+OW
228rYDkkRFy7tz6gpmhqniWE/bBLDps/NBQldw5Ka5TGYbPwGKZsTjbz+0ydHYum
0y4ggyQtrripUZXzUf5uAJ7Nr4hKJguYfoNumCY5rYZd6dEL1WNiHUgFpSx6GIMM
dVL/XS/FmmSSB3JA6TBCQLjJPTc3+voSHjeXopvH4C+La/ii5bvUT6W7sQHcKFww
1bdE2arIWSnloXYqvUWqsl/LpfE8SpuT1/Qnu91OMemZxAnYTcH8/swMznEoOeJz
YrYblenj5zOTYq1T9u0RGlhY8MMzTqEfrbozKOCdXAV2/CPy71S+zdAE6aUvsLCw
HC+JAw+rBbdlN1xDmBMlKSTGng892N8/VeAQDlzY3bdDSfipN+WveX7Oi1BJoquB
S4kbtm7hjhYhmpftKJTO1qcQMjRLH67UHbr7m5c7OKiXpjjfTI+hb+UbG8uY6hTk
/s/mGnJK08zbo4BuY/33N/lfPuXJa8NwdaHHjBBAZdgOn2lFHd0TaCIuonMcZshf
QfDusKxYpquMLHWWY8n6ZA==
`pragma protect end_protected
