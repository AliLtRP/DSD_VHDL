// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:26 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
k5XOiBcGgOhTJeYnURLosmMpI5yXaJDFIsAbjg4V0luD5lyvndgn9q3aEUnrthx2
ZcpyUH7kFF/i6s5fctDsrB/uO2x4/8dJ8wrl3YhCfGIDOFC8Ixsm3m1qtHUW6I5H
LBpIP4QVfu5QrttJgabF1JwpmBaVPMGNihxwwZvCbrw=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 9824)
PE48H0RvdpV+emxcxGqsiKLo3ZvJv7DkdoIGTX1nJUTWqadNDDjqWeUjd9Ro4L12
qLChA039UZEYAydLBJ34Bk2dSdNJzUkqWBFeIsY9Pv3h7LWEpWI0NkRq4DZo57oP
oljgKEDJJusibOIivjhlp3pG9kSWT7huHZcM1sUEwOmkA9UoLUDjkU7FTuCIg0W3
kNBMccKYK2bg5M4Ly+FkrVqZQbZCxKy+UhUwQGixjr0PsFDdDuiF6Le8Wg1XJK6q
tL+guzBFGdriypCPE7VJUbcnpqWS/zsvPfU600/sPKfHDtEmHubSd37gr8i2dLda
zLuEdKk8b7LrMnzZxuVRKiHdsatCbMJNmDWjE/WX4NqzqVy0JNn0Nj7WPhW4fb3v
Tr+iO+27r9SLJenbTxUp2Hh9mia5H9c8R9xfpE1hsT+QG0z1Wuvz41UCd39GrQmw
p0iTVshGaUNqhEm8j5KPsBImfe9xzgVfDAzw3yG2dmXZweZNLAWySGiKgEcEORKi
7xyJqi9nr/9wnhkA6PVihuCMzI+LL0+Hh3jtbI2BJIi6Nrd4e4qWs+IYGQlCskoQ
TXIdlWzrBkEb8e7bLTeY7UFSQkrDqfqpT8G1Y5HvCUZGRw41yd3lr+uRmFM83gb8
6Hmjtyo+NC7FbXEaD/BWm1cy6m2CFRodUFK58jovxo57TmgTXjS3YWMj4oc9WCJA
yCeYi3/aCb/CXa07iN3k/k5I32Y0M5rOT0CVCjOnv6Q8mCi85FvmSj5HTPe2phYJ
nJeUNXU0duHMVVSx2xY8TUn1rWIyHBP6K+pG2gi1+lAKlZxIXYkrmN9mneseOlv+
HLCfGmoOCtIFdjg9d54cX87ZPON0ZT5FPofM3bnjPyr7KkyccjSi45IgpqBUY97F
qZqAk5EFupXUa9aodHPkgoDYzLkONQwpitz8DvzQyO23gPiZG20gR1IKV5qXhGaa
MrDBTW735SCpttgFMh/h6Zg54wasrwqy02nLBeE/pxl0FqFC6+uFkdGAvvEpYD4l
Y5wFdYYskcjrcK9AF/tSkxpWNbpsa+v9z04vXimVKtSiSjxVe/POzBPRpCYZc0Yw
BXv7YTxRUlvfPzNzt9w+Y+hIvm9/x390RzwKM8a/f9dRPWWAre1cjasHmFTMSNU7
qCZ3LGyuMgGwyoB4cEEhiJdWNxi+wF6Qgkq/0bh/n2a44ayPS7KWx7tWDO3WVsD2
RuXi04GwiplVLiGafREBdj+xrWwWFf6hrA0W+jmZnh8ZbluEt1wyztxGb6SOfmJe
4Hi/L4avhDOvvDgOJrW6hGYoBYhW+NLPZiI3O1v/VuN045BRaUIsSiaRpqHSBXI8
VuTjopABYSFaPFEsg5w1ntL00cZE3S3D6g6EHhqhaydIc5ZiP4wyPmcL8AV0mBRa
bvFNN7S/QFXBI8/WH5T3c29PHF51MhlEHpB28wgT1WTOfgM1rcvNe5L+CB4gM4fY
mNCuNM7fZbBs2lVdTEa3njD9+H4tJFNa+scSpAQaPOEkOia2ndEZQfrg7qAfGmkM
WhyQcq0wnCqBeLwd4p6dQgFlDJhwLACiafuaFfcVwX+MGNRYaMBa8+cKrHCwry1N
aa9H1o9cqgVvwwDvHnO/ZTrodBTrJybiHYEMQQcimg7dnbhorZPUacU70k8WAQ8T
0ctMMb/pFtOd/iSVIXiZJlb56UcoAmJ5tgqc/Mn74oyedQKuY7roeEEK4/EuN9FP
sq4tgMIfUTIIx4oA1z9P51eSMO/0z8ZF3HWwH/P6pGpJT9wzNLES4nodpJdHjMWs
BGtW8PXvAJcl8C7OfUdaxOA/sbJVXhvSspC2ScM0a1e9dXfi4HLTuTFy47jmkGU7
0snSDTvbtSj2kYLNwiWDrfHcmgwW2AHauJ31zTtXypu5K5l+HAtGhErZvbB+UM+Z
ZLBIetX9gRJlek6w56FaKgXH731I5GH38Ey5S8PFNxZIW7UoT+K34UPyd/OQWO0m
Dfuh7q6LFGvQnEdguDw/gYiNmfyeNnGxhtVnVNKLCa/dMclT7jDtUJqBfQbkukLu
B/R+kAVcy03SWkaRGqcdMs5Sr2GnJRq8oS5o7xBg6Q16mkqBzZAO0WySMUOF7GnQ
so2Cu1+Dx5kql2WBS/cFtw29V64BclrDh68RjgBa7otw2sygxRD6/KGAMzRpe+7M
HxQ70E+EHp/8rs2+xszZDPFGyOJTR12J+iMkSswxiuTVFk40FUbaGYy95WSY8bNe
k7+iN8rcRsm+M1uOHKr07obAFddsV+Mkm7fS4cWnMcx7xsNd/XkYXGx5CXt5ytuG
kk/ZmBTcZDLsZHHohD/sY1T4HBh0ixPwDE+h2Kerr3ZAGZFQVkKnuYg7neZP+uqM
6v9MQDYthp2EaMvWn5d2ikNlhJ+K8rW74xMJv5nlMeElggWXiNPkwGpYlj5s9Zi8
0iRPZBYm40mlBip2uZA4G3cVhdeDauu4NtnxrX7nTfkkLi7bhfn3h+2SsXVOqgJE
pqTU1QScYcqIH7uQ5arO9Gj0h30FlAzgzygjLQHzddtLtN63KxTxs3U2eR4vb+FX
0TggHRkGwqoCMnb+olIejo4V4tGHtLUzWFkZcOsEEK1278zheW1nZQdpNbap/G2D
t33fQae5NhcUfJKPZbWC6SlDlXphIxw4Jk7VzjbSjyHxP5/9ide4t7QzTUaBnul/
avSIItwZ29tuxmgqfVJxrx6WUP603wuYCs2NarTe1Y/ppLh/rRmQq7OhHASZRwtg
Ne4FKQqp1MsXEAAGGpgShocNVN0/+7X7TnH/Y4AD8V1TmUFKIOa3Pk4kHrnQwzXG
+gSeR66Jy99XqlLKyOjIDjUBOSwbafscAVPCxUy9r07n8echc9oZA0Go/ScqOb/O
voN0ZGxo3qzpNV5eAHsk//DHkVC3aGkOPHxvyhp9pdPGg0Trr43Ld7LtRZ/4LTCl
rg31ZXwhOT+pC8142hn8akXID1HOm3gV+GrYY9/KWIF9GtO8biC9YpQ4YfdwBQY/
XbfCkbEYgi7xvdiIwPR2kkUR+aziBEgXx6MzPUr1jysOwKhGqCm8n7nsEHmyKKAf
ZHc0m+KHAdDxq8pweTp/up4Y2PWLvFkyql50r0qOL3F6xlebYZOk3eFf+ezPG9PN
ZI2m6+lfuZwJ9HsrOZrKDIisAFH/RTNDlQI4kfqHAONFw3IHz9Ufcl8WPJKwBQta
ZBt2yXXZikO5Fawl1PN5e9TclM2UFSqr97V1JraCLOvKLrCI5J/K7Zli6/wKwMIa
A7UczT6/5O0kJosd5pQZhoE/SLuR5RBv8oDy6efhB5iTgjeo6qFN+enK8Rrq54RF
Sjkl4g47UycX4lkYECeOkhvaDE5VAeR+SIJKHGGt5t3M7ZQb5kYNd00TVX4txcgK
rPJfyRN4223p/RRwTPuOXKKUVms+7+SzFJL+DrgsDUod9492PSNKqr6BW9DiZXIH
zKKX7OE+qDRgijZTjJw2gMO/0rHVEEIz+/4SrNu6yFCH/hpzy9IrrHo8cFwaZ/xN
XOd3kGKZc0Trq6QeDTpH6pQT5UGBvDSlksTGllfOd+5mBAUoWnGIkETQRYcqM8Re
NzZlrsHk3FhWMkDTc0w6HykRf5lm5+kedpUrs9TCXxEoXshEoynQo6XlGriUsVyZ
NLZciDK7/S3FD1Bs0zo6kEZoJQyLPh/jMXWzCr3SQO19fW63UnOZ7G2AFyhWh7RB
DbPgkmulYLAVBEFAWc7hKqGz79a/KSHt5DSs9bteq3XF9JO/kTkE3bqjEKr0xymN
9WNV4wq7s27q7jpCynzpwIJ2pjhjZqTmE4fW1NEznEE6nBKp2rkqESNhiLAar2Rw
o2lb2SHQuucV9ElFj+yzsO5nDeQCgir1DUkpYI2SFOOA1mSImFPZ+QkgU1QoWJ/e
8DQamrgPXH6Tw46ADGN86paef/6ttG7DfRZdr7RnggbuY9tN8W6BZjkOHA+Js2jd
6fh6uROWT5dgp/c6zsYc8MqufKsC6VRNU1iGJ9dDg1M7Sng5smu++zPWGocWqdji
s1W2lZrcVWJr7ggqDR3i9U5ZuA4CmIiX/9O1H1flJH9uqwVhVLzBiK9zEEdEjC5S
wldxeXA3yyYt2GCOt9SPSy4PSObA3JAqm1Jsz3+flug675ajjhe4q6AK6NLfORdb
Oj5cJ8xuPawKVT4askcKcizq/i16bHmgUdnmH8EXKo9oqtL25ZP7Falgo10RQWCN
kk66qJPLxuPmLPj1NvhuAkVJ/Z5rC8Iq3Ezp53FRICJk/KQQ6IyXriX/OlRnkj5b
hBxFRqPcXFor/9kNovUMOllJFNJDzeSybL0LDq2wt4FhyMhewPl4TabAl0aLhV9E
2QRUrWN2GyLUlxwW0Ripree637KvILog0xsnQaHASmAmEs7nKKqzQoQ/DOcI1sga
1UEmegpDlbmR7WlqXyWsQNmq3OgSsawnSsSRNGEMl0N3YacMRZnn0AlNg9DKry5B
Boci10jPMN0JEd6qOy6FKYRK2uQ09fy+/zmTneGhHpmkOvzXZ5hq9417SFrtY9l1
fvbXGraniqyocGIR7w5F3T8PSm8JKjZQ4LX+cchUEnP7FMpkL4pNj9PfJBAuefhO
TCK5vMJRZ5XXpbIhM3mrQHptGh1n01+eRb0HYKHv09oCOafIRgBFKRtniIbLKRqg
MCRfWZA39vWzI0CRuDl8HOCcdp/rRGOQLTF+WYMJ4AcDRxWAr5bposDY/lL0/Aqj
MIiGkSvx3au8XU43Gm3eyEzIAvRvqyaNP+tAUcNXoLrgDqo4XyfXLLqb5AAtcIc2
QJRmfoTUu7q/j+ZXNkjZ0HZ7Cv0Z6oLwUc5cTxq/z7j/W7fFFJ+9TeaZWvCRHyJr
orXvezJ9ZO+0nq0fyl4y/IKG4IrH6p8YYxw3rH7GSq8jWXAm+EWpdTUm7fqYJrgl
CQivIr6PsFVrs/Ee8XmZNgl4mBn7pfF1B9xggi7r10AmUkV/VGuAOu8UX5lFR82S
sRKx/8EdRASXILhH6bbIeGXh9IsdTl3LPTuRujhPxy4cfIAs1EBpByDIGqeJoeAI
gpD0fqI8w8V4PK/OzcQKkgVU0fIzWu8X8x2hOlM3+tkSvpO2jCBA+0cgDTuu/H21
zo6uRM1a5laItClRfXssF10cxLwzkHZtWTVTvEZ3bynpOPK1J0+qfAb7tdYwv7I/
L6X8h0gCyPtwLx0oWXjW/40CNQLXJSvkJWJm8Onb7VNvbxtOJ3Bo2dkCVeBHvFMG
WF0SNnn3htskIawk00OPjPIFVXMBAX4j1oqQTjFlwRmuo6pj5vGphmjnCHbPwkBD
pkIocN2QCCoaLXWqm+mgjvS/W0ffDfpnjmpEnQuBVfCNQ3o7sTQehFW2/+Ph6McB
o0B9nQYDR2gHcpWy0l3eqk4sW8opp3KojhZTGc1ZHqEl5n+RWiaUZ/sga0SlHJSw
T4my2TznqwIw1p0aOOhvSUVy3Ra0+PLanOluCRWp5wEJOkYQUISzAix4PLUuOimF
hnrI7AyVrueF4RB1GiXoDSEoVYs8U2V4Xm9jK6ZKeHEyNQC98bScQzxhkwO/Hs3V
2YOWUgozSjz+5JzNWxFoP5V3S+ROBpCY+RW102nyJFMvLwYPlxh/TypplstSetCf
XX2c7rVxCmyi3w8mlqAhjX5FCB0u0atY/X1N5t4jzLVE7f4z3PcVi8r6TDny8+JC
mZah6yN56PMhIGhtyH0HkXFCLEzsc+wAf62UomN6ROQCnVnCUIR085oniqH4Xzvg
yOzlKig4EpV2eQN1XSNX1/45y69QYWnfZfNMEgtwqDd0oT4NQegCMm1gqZoCjk24
c6JMETX13cmKik4AwiOv7tKBLh/KGbPlu7bKtLXFEyLacEwohYDZy/JahgOwrgLY
vmwN+6NtDJVkJIal4+CJvZwrSGGkNqHfaraWWxck4PhzHmwZmIKm5HqKkP+X8ByN
JaokfYhTqImg08ZZClDZuAkfa78sbGi2svgvpeKQc/P3djvi02oUVpM0qI3WITKA
MfJYfz6oKifLTH1FiT26R4CVz8H7CYYxiD75Vr+i0KAu90OCmQyms3Ey4gySuR2v
G1wHJCWtkD+UisjnVjYaeuCZH7e6hYyMsLl7rz0Lyt7ASARWqxvDlRmYUY01KRhF
lfUi2GcBU48oGyfvRvh7Ev5VA8TB13QBbXBklKuQ2W1PMMSlFwei55JNPG6qjR2t
H8fpW5Kj35qRGusbKzmPzE2HfAT3hpoteD0OXVGgRPxklRI7rmoyUtmUh9t39dm+
WV9zTHAlG9Q5L9Yu6bG03CWKiPUDpIu81wAF4va/Kgwt/HyacKEumPhghjHNa/GD
kt5rXSs302TGQ53hdKCqxAaRsyJ09IvFM+xIDk3ndI0wtanI5+rk3mR8Ui9KyacF
4ISwSbOEN7swWC/21vF9jzGHo6269Pi5ooHZDjDUl7QCkAskFZs5riUWmI6cb205
eAywhjSIy1rHFtvzw3Ojp/2MYb2vLOf1lpnybkI1ZgvpzOyGSUiVKlHNM3yLtk7v
QNmhCPHBFG8LrDvfNgacy9tAxt63Uer3ryAmyRXW0CY3FNbEUMIF7iHtUW3lzwFD
EVDPlLP7nLO7gW7QdT0jsLHVj7D+n65ezfjDTVX4SBn6CRczJZrZSUuuLnCXX4Qq
TNuvLN9D5S0bN0ilviPbQQNcLF+//fqKD1I6VuhE/y6Hf+3IQSMcnrxERWDk3DsG
QJ55CDZepuCcAJcuWM2f2FUi+FpG+YzGo8RYj490BC+ulckfbDDaF8imM/0sCsfr
1TkihAxYbS1vMNqz3cGyaNjH224gGvg+/GhZPm9ISY0/U1KC91UgeVZFSbEldGXR
sE2ONQ8DHaIshM6IDhIOvuiyXjEgj/7mpDLobnnUAfbjK0gg7X+BLfHUWYuF3f2R
E7c27rN0k4c2kXi6U+f3VqjjC8Uvsz8hYtICpeXLTETg+2w6m8DfamGNm/JBbmev
avAF7G7fsPvPaZjkcUvJAEaL8941c1kHDMTQjAWUXQjq6NiCrupDe9Uaxpxm3guw
Ri5gGuA59nznHw1p3Gee2tR6nMAV3UFGc6/lcXhUuBssMsREyCuPJQ+mvST+qFdF
IbAgXRbwRKQqEXTmYCcRPqLrJyToAzTUIs0+YbIN9BpS9MaBBnvdurPHj0YXguuN
QSqFkdK2aWBg2cg6hT8EkeN30YwjR/lWuOcawjKBuslQtWci/n0frGD5GY4tEZQK
wIYLPyMqpkytnIBi4bj+ZwFCxdxWLrNGinNrZM8aLVog8Ao+OYyt+83UHd61ILr6
7KXFA1lXJa8MbZVoaDJqRr5Pni1HRRg0TXjzgVB5gQuOHTK9+kAMKSsgtB8oRRlb
MWXauZqCHMzyLAX1Jv1hCYU2lJXnhv4TwseVVw/JO7DPzfPT8ESajyq+8hzP1lB/
F/zvlIEtbGCgU5vLJHClE7zeSJOnUakZN1Hw6/Rb+284PuDZUsW2l4KZIgtu0ZlF
BKLbelLqPawfkKIQUhixMAEQ8toy9eN5SR7UnnuYcT5U9qA4HejmxApcgo3hsnqz
rAGlpUOb1IKCyEyeHP/O+1mIgbTUXbSWkkbAEfn1Rtvs3dJnzDW89ORJd2zIfWuK
jm2YHim12KfC1Imn3HOfwZUwS8o1zSOYwEyNSz98KFZu6hQadls7aOzXm5bKX+8a
IWv4kjEAzBVr38wpB9GZQ2qDtw8I1gUpe2G4V6zMoqV0RKZATWXWMY7PX96AHMS+
1hGVQvUDBuTFG7Y9xplJP6/eCZrbXFw+4J9GmzCLIwIloIvwAEEbqPg7Rwgq/M+l
9zgg8RLbnDBAg7qgjxkNamuyYBGm/vYQ74pVSAB3kYRf2DJFEsD3aRYpP/NxvR3p
6IxtmLFi3UF1/IBFCorW7SGY8zqJg+SSPHdxITmmPmHqT08Cko2evZEASSmcO+7e
360y2kA1j6L07fnDgRxRu+6OGBzUyy0lcB5w+WQeaGhlVRQQbbllwZDxUOHCI/lG
mdjCVJZ6O/Ylu5Ox30UzzWZuwcewBF6acLSmh1kwY0Ij8vxyd6jha30kn7eihtc/
4fktrMgap91Ra0gR3pCc/dyko92vkILrOOK34UZg8OJCfiwKxi3jbqH0sr1bfIaI
tnYGqswVLBU0tKKvRfVp7iM4ai5PULMZDphSMsufavlc4FlFYkKA0wAHVfW8fceB
yPvFHAcpyhKWqJv63g1iBFAMogiFYQ+wpf1qZPS5svdkk5K+vgA4C4vH1u1wveKw
5TsBjJblnavqVeCTTBDLmekQ2Gqa9LuLE0YNbcyEVZTgKZ/CCH8PPhITi29gUOt0
SE3XTrR3OnqpfBhvY1CtVbR1bMFarz43ixhNqQuYEZ1xDqLc9NOLnGSXWhUEBQ0B
EGPOpj5UrMEo/g+4TQXHmKx3vXZhFV66Sqn9YPOpYYS5KhLiyofVkDIDtOCG3rLP
1b4N/MLZXEj0B6EJ7geCnK7WWRJCad39oEZL0juoALXJtndBeS/QVzpVe1dQhKVi
ymlyrIQEB3nsKb0oSwPoynkD4GWNblIkPo2j+7bMlcpBTFv4fLNhYD6kPAVnUqYX
qNieoNUzm2E/cQnxDzd3yDIcWrAdJXzaufWMFa/ypgVCvoKiJ0fkl72y4wFshKrd
F/QNyIYf1S0Y6YAUDC+BivNhCacSoQD3m6zhf+/1e8/Nt7s3RbSaPpFfUOl06XpT
oYSxYk232OWjTqrl1HmFWxwv6dmZ5ur7nBqGKb0FJCOVApEJkMIVQXharaJZE3b+
M8ZWNP1l4GAx2AbAcWqxEnsDiIZiWEOae58PUzo9crkpyp7dfDp9l1GgY6Ak1Z2q
BeE7LqyD1+Rj/HoLdmHTR/JtTAMy9VitG/Gq4bj8MMGDJ7c3oe4ygv8QTE6vRLz4
EHbhCcCjC2ZLat8AArzws/16vByZgjRO0YREh4IhkQ+hOiugClmTw47xiVbcIgxd
AMdGeBRWDylP5Lw4RRZMGOlT9P2X6P3/6ACFr/Inv4V46z2oy3Xn00QIib5vEysL
n70Tw2xeiwVm1TEeRmPlK+KgfCPAddTWK8bI2lQPmDOwuTq2cv6NM6z7uWPHtUUJ
7NdgyLxoumQeVT9y3Ngp6nfMps0sJOadgVc/iGrbwmiCbW+y9f5y7auxlU/kpvy6
XfuH4R0Wj+OMKOAH0hXWgucXYz7kE0pGsOHjKmReG0+sG46dmaz+IASkFZYjNe8N
mZcJ6j/0D6xUAnps/w8+MMURI+mleCeP6nrvc0SLb7d5dD84+mvGkrHKIBRwHS+1
57TrikYvQOBQExK37H7tooZxnZoe/Ik3/8OTrCZhoWYz6IimUPhi/hk5lW2aACGg
TQNdmAEIqvMFMBRPcPJGjwIh3zmN/GdhVMJgMUZgG42MITIOD9Mg3Y6cibxHTTUH
9Z3cpv3YTe4zpXMA3GyqrAufRHsqRb1abI/hyd3IBSnufuUGhKvqGhSqIescLHmY
rfK8aqGS6vU+MjPZ1reqXsi8v+Hu/YHA0++3vVsFsGlTNmMNtTywSIuNeuhBYqgD
5RkrVNQPJszpzp+ytkzJJUd9UjpDblhODymrOmeRbv0Zl3fRDJTR43LnVL11pwEv
hIrbpyLwPUcuwAZuE8rMe7Mnabra2FR4u9ktQdBe1DjBpBeemGcXt+o8Lede9O4y
SyHX2RV5tZavGpRRkQVmfotbwiP3J9i58c7myuFRz8T2bNs1EMKzxPmqdg8DRzmg
12Yd6rzE8eqnjXpp35ccLSSCpp9g5Zt7hewD7Wxr65WJ+ODO67CDyrSp3BwCtFLz
ExnthpcvacYPUBYx8h2SH1PdENsonLIH7B4Z9v2wOMBgdtGWbu7h2nRos2ljgQNj
FaJM4/uAszKZn8OkG1qOOSPjAfqj/ICALyf+1iUCbwyqaAnn7Ykg4sqhEhMJntpp
fUWYYWs4uirbJlEFUhoGky0wCoW3hoWA+BrSbkC1SeNJCOmP/O51OmV/YC/aQwSp
fiHhpveDg+fbEGF0H52M7GJhg7Vo0fgDnqzvnS+GOYCoEASoX+ZUOE+5ifroWAYY
wOktVBCcBZ+Ulz7hYxzyMJEvf0Vo3859+du10JXNQ8LJFFXYfZCMAa5FAr8xb6jT
DHK7IBCVxHmAmSYVZYe5qTDRYeP65rE20cGMbHItKBFGrVOQHqC4jmLgRANMxH7D
ZIDmVYeVWULMNxR8+YDV3XxnKjWtCf5UN61EMFYWasAhIJeDAUGSsfuSLdpXbwLt
DvG7JPn3iI7g64ZAO0Q9sTnBDBz+qnI74Fd3tTw9C3z1PVNxJnWOL6rjME/n2SDu
qmXHq3N1qKLDRzAhxCi4HmTHsJgMY/vSQEXJGzFOFrVtXgxVM3Ae24avtvz//mse
6hRsf2f6v9mcBQFVKu5BDIDByKjzBIOSM6aKF868DmYbagMkWjs1JU16yvaEgoga
Sa83d+X9kJOj67goXmP7eC90cXFdFfiIqb6GrlzqpacfP89xRqHTev2gCQrKmn2T
MrT07hUbTjUDmyewOoUGG6rv7Fu3cTdHZjtlcGef2qt4rBJpFze9AY8w4IMpEE8J
6wxHrQWJhq3cTJVYIT6LnCVVLsi5ovx1EYr+GGhs6bAN2SMkp6N8Cz32QBcOGeEw
p+dtRnHwWB5unY/iZrSqCeBt454LlNfolUlZPh/HlbpLhKRXIzE7asQ+dm3QCTwO
sUDWEOlGPr1ReSxhDzSUm110da7YM6XYf7jRxFEmwdgs5TZoHJj12LzKHf+mcCZK
gteFnm+bjlyYYnHkg5TUXiUn6Pzx/BmThWxaFoYqwa33Afz+FtU47XQAfIeSAZAF
FDWSYGQAPaXvC4yxNU6hIf9qNcjOluZzWfCCRqRBYDqQ2vZQKyxOOVz6yDoTumWb
KVU6RVCSdHtpaktzist5ZHG3fGvDcIz8pCmLlY6oKO3RvjXBSZAFO08cmnEo3f2W
dbUAEXQB+sekuzOf7XHf0RTLQlJmnIUqbcADRnwswof+F/BM+d+ktpYt0GaXHU3s
dNDd+3cQUX3wcFBqJzTUlSx4t4tqB5J6makXv5LKAuVOor5fHxwGe13A6IXyqsLr
OAm9vfYZCiob20gUn9Hs3uKNsMvu0sySQ5ek155KGOIsQaiFWQ1RbPU0Y8P5R1WN
W13E3miiocbXWj0nZCFimm25oxGyqNkhIZF3HX3iun+tcQE7B9lhGLkg04sdEm5M
6hFLuQcOleHtlyXGwNBQRthiLaK8u/myP39lteOcI/FpdU97xY8i5H8v5p/zWI5B
aWpSGsHpWig6mE5gMKMMOdCS0EaFJBJXff9fWBDw1Owj+wRwaDErxM6wBWN963Hw
UJATMw/I7k9VDr/qKEwkmTFxCBFllK3YZbXx8JeDBHcLa4mZmER4vl5MqzzBRtsX
LhYZf9ugq4NyewlW7cEOyUsFBVyjqt0CmJOcrELyJ9FqPNlY2i5ZQ77AhNGoLNfg
RI2qdS0t5ZdM4MyD13LMNNWosBeaFInZvtQzl4E25lwBEGdEkJ1avxuiuYbuXirN
n9aiWd9PAixbUKuPQY2P3IfMFxyzYcCdhkQXIUa5qTvTd4Iprq+opgxDX0Yuraa5
cFEokpcXRi6+IMZD1Qvxf8qETOOn0dHy9+eDDyd9Y3rqK/quQQxV8OYnmCC2Voyw
yR4L31P5noR7WNP8Uj2n0nbNIaGLI9VhG0H/VraI54+V1Y117z60AEy/bl/noKoa
plDMCqW35VgKmH2fpos3IQc+/B1qJ3BK8c6sm/ooWMnYhgIkB4kT5SgpkgdcttdF
GyCvjcIzABdCk20q65ruOG1p/L5CNQI/oufr/KYREd7lZtjcsdIkOnV046QoLjtN
7AGMJ9jctHulyeg1E8fm7WBic7rE0tYI70a+VlQx4xUwS4ta7GdpCp1i+aM8nju1
+VanJFrlgX3oBLCXZ26pyzIcXNGXyx78dUOf9ZS/rw6xd0B7bckY/RX5+ucCalX/
2zIycKos/A2QFX0bi7EGMhgeV8K0RPVBLomGPAZ7YQcI8peMOqXw1pcMnlsYHT6V
psWu6/U/zou8Xt+Hf4NYElKtrN3cuOvVU3/o+fXHB+w/k0g7EA2GZyUX7ZVB8zWB
NZi5uLqWj84zpb8A4/jAE9ku5FbuhISkw5mM3lgcBNx6LRnyM3jSyRMU1sLLTRy9
YrlyDQvKF/HE0EhkIbSlL0OwbjVJDVvZEGIMJ205D4OUIS9sb3KowB/+o1s7Yhu6
PuykyHgHDzEqpdGf7YtxNk5KsLzifLWfhgAI71yMQ9cuL1DQNLkWtvO8wFVLQmz/
S9GilB84czxOa+U87EPlkfOv/acFYqXNMJsgJtp1idozWjxZbpTihwbAvysRvUkX
U9jgomyXRf1sFkchZPuUzWb8dY9/kNuw3utjrnI5GeoTTWe7L696Lok0vJIWYqjh
a8qLYpsbqXRoYt1ppY1ciWTMJGnDFKsI4Rv8Af4jjwLzzxNKTACYrB+5DbVfxUR+
hj1YYSsTcTS7pHcQ36YCJeoHuJSBtGEtOL7gU+u+Ys0UBwlXd/QxE7NX/+zUOPuD
xvSIkMHmfNMCS6G8ASAFn3mpy+vyiSrd/V3bG5X/eNaaJvn/8M2zIiohamuChl/1
7tDTy4wdRIiYh+meYGipqPD/cBc5u6CdGPJtT3/+SE6VNm7iWjybskZAkXzb24Lp
wHoA0A08YN66RTzoFoxu+zIWV4mZEIveCefTx+3hIbo65YHGhDOw35tUg0s6InYs
vVqRNPBOx3s/pkoxBK3j9AjwymZ5tycyCtO1kTTZmCTBUssAQuMgm5F5jtwDoB0/
es9ShklSojSM1dtW170uk8koc4rEoI/sJi3Ypkj+JdqfHwWIpYfpERWFodFI8BzU
wKs/8TItzgRurfK0HwwUldUYKdotY8depIT2wAdbAqezEMS0yXbjJ6acozk5YRc+
jSCUMcF2lQ1aVCvQaRMS5TA4DQHNO7wdT1VSRlCOqlK+hRnPRQ5BsT51nakf4X7C
fP2UbsjjBmPmJGjyTsHC3kxfW0/8W/jXMZUC2XTkpXZkVQb2jxIorTReMD0d5d5k
C5SD5VQOOI+r9D3L30eXBSltjh2CjhnYWSiYHUlg/5g=
`pragma protect end_protected
