// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:35:27 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
rgNrangxMh8ggdevlpyNNYL+qNOFGNy++ts7HkpbwMeDvx42ZLBsBZ4HyWh64nxs
anEzxp/xGGB/E5HFbRmOdgi/vKXbRRJ4rSTc3tQ1Fym8T9xPq0JWkdxozlCQZ7g2
SmEHvU+Ah0uOS1CsKMMCBxpGW5C5qJoBReUC5rt9fDU=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 20240)
bkXRjGi5qLgJIkg+dgfG0m26AHf6357YOBWVZPwc0OIks2Mw27OdHKSt/7O13VXh
07zgkWGKdxTGYeKc2N6ACTddh6OnKerQruszHGu9xzzSqYh0vKwmql3rZMmVdRd8
2tKPF7ccw0Jf33O+4PLDn1VDS3CQqbvsjSPV5ysSrj6EvnQBQCkz1K2LH+dikw2S
pBXgKmO/3TlRMGFltZAEMsiLfAxQkIp+8yZcMe44ExdYrBhAwrJh4BOXlwBnOIMS
lGFRQ0Gthqq7RIBfhD+/iSq4V79eQG4LoTKK3sMslkgy4UgU54vzt7XkO8SRUywy
/QCxFq37X4h+uVinYU6n6dpJUhqKtPB6EMmRZf7HRZqqQTouoUR8CZaRWSZdkkmr
3SOKF0Uv8YBKmvhDmefVmDHjFeWAp864d/mUW0vL9om5RAZNmRu2kNYcQ9a5LntZ
E6ciHzc35Dw6LY6Y28mWsTKooAwdubIfRUw+20BFR+ylODtNACkzTB+BhUUjJCeW
rWdbGefp9PxSBdIpSRr2j6RXM9yLQbtuWaVFs60tuC4VB2/D44uGuJPtGBsST9Dx
fbv+x/Xp5NosD4UF+PxdgtAF+lbQ2I+8/kT4QbTjsF2Ir2eyhizC+whP5yRx0P+u
kBIuUDB+EUH2rIhPSUZlg0cXiehcWnY9nC7F3S4uYSfC1ULmlSWgi4OZbnAmQ34P
EnIMpa/MJI/xbI/DXvvu+OyOHiIuW/kN8M8oaOeSgACxe8XZXcuf3jyl4sTzmL/1
3B/Hl6t2ZySlMyt4KAh4cpf+sEhr/icsfVELfMnkkWxQ8j5mTmxTmoOBmfFL+sHZ
wYw5jAgOlyACZjOIj5D5LHG+eGF9NB7AbXLv+tjOAsizGwqxy/l6WqLPUSVaQuc5
xQQvVr52jvVdt+Tjez8SP5P+OZ6UkwLP8s1KTTTU/pr5f80vutmgwKh+9JGQRs5D
YjgEeoAO4yDoUBxwjCJpPUQ33bChbu7ekscnX9pIwQalg9U4J8/SEj4xeChz5B/S
JHbUWtHNQu6kKgj0ntIVdrur+l5eTzs6qrUMwErREVZJUIN45KAh0RxoTBJL/mnR
BXmpRSo7o/+0r1KpyRbGh4Ui+iYcPmFwTgxnuVdeDBHgwWQhfJ/wRrri8cxbnOvt
X3p6vjsS2+txNfDDR3BBowD6KFicc84FTL9tUQSEsXsPfz2DIpkZ4KByEC+zsIcx
/V6bQFjLHWzYU/fkjB4yJnyxGuEaUNL3y4mRMOOf7/qlymqfFqxvlBvViKe6zZEB
iHzEWXravq1WbHCpNhYnwdTyumA04Pm99hsuMPkeyqsgtjS0iWNCPu0cnjT868l4
aJuSlW6a0m3n2aUfJwmFUvM/5OGUv2N0LsH+PESZOL0LAQREyTzVHOaISFlJuTUX
GqjeiVnYgZsoXcm0q4nFbCR8EUfBfZosR3Pw7693mRs8gixyST2qtIppLtdlvWbT
/QE7IaIGvhlD0bK2rU0tEAXYMfvRfEsfVQQXa1DSMb4HKuN0gj1FIP9PvhoTxVdd
EYaUWy/Ocl7GdQ4eyRLJpMh9zUbi3SGxgcUa2TfVzQ3kL2G+rwudCQckjFZzr4+5
SBWsNCHDXL4i9ee6LFQPguN1bbHlNLrtqRKiyyYUZUSD7lDjduv/Kl3Tk0t96ItY
zVMfMHXsF2NbIxvKxz+aGRCYRBYTQqI4kYGMf61y6vLsph7QioMbOXaYHvuYNHJ9
AWTOO0TIlAfnTiqGp0HWrE4yF6mN2yDAI7XnJ1qZZu3YHFUkzttoEQat/A8dpRq7
h2DiPWSlvIPxMAX+oJrmhGqSoiaFcxLZtWWw+m5D4vMrde0EzXnxEraCW2Hl3SOh
9OV8ipsKrlvbNzD4L5nG8CQJ/NKz6nxOx+94AM8vg2tosVk9G0X10AH6019zCCDb
89IaEXa788HO9021/9PKU8P93ljaoWn7lqMRDDXjcFfe57k6v3fDPVZkWNnJ1R5w
SzBw5NvGwwq8goUXY7C3msKsbAzftXYIvXKuYsdVzKA17uu9euMUix+Kg3S+5WKo
NEr0RHHZePdQ1VDj59a2w5P1CcHRUdUGPRyPdA4hmyHk7Ed4pLoyVVxQCyhhWK90
2ojBxhifzuThqtYpRwuxmBepaGtg0swnHU2OTJO7fjgoZgBAv0lulYOqUSHXP0YZ
937s+ewxTAfIOKWpY6imlKwuZEWVhDfcdsdCdospw4lKJ7kB/tVrDW+yvKUIDBli
pn8G6JglWule6VUz0swPpVcvUr9qXRlTChROrWUOAMBtiioj+euqIWz/K44G3fr8
ip70h8E+DlZlPgK+4m3uAWr3mMlMcGwkNDzYD+mgjEaL4gi+jlKxza3xLJURiHwp
/RCPHJi+Vo+PKqSaqxoNMnWhHTh6RvoZk++Xnl2j55Jj/ocyy4GE2LoB5rCq456l
vDxmjpEcJuPQ1wPqmAWutGN9dEAzcjH9e7xwGWrRaZ8xUXsKFxxZZWk6cq/6P/vB
YIbH/cAG19JVDh5brWG8CJSuqMU+x/Uc+RruE+00qYL3Wuoa+MREJf6h1EjClq4d
doKA8UMJOWhY6iBVUyE+JS1G/hVZ798+wr/hkzFfPILv6B2cfKzuyS/I5hDEqMrE
86+qzJXs/pVisl/7P28PcgToeW9UBwS9SZhZKwGhVHkMI+6Mkc3K6Q2DKQwwjDfP
IzOId5fb3mVWzlMJ8sO1bgwi7LTgZpuS1LzwaJOytXFNZ6AVoZE25ukLwqehq+3r
E9UjX3thr73u54qTWovdwkdVJth5yx91uepYyPPRhg5ZxvtersP7t5t5f298FOSR
7eUe9/NctwjDDFvS89O2b4rv8jVC6aigyZx0aAe2zvk3hZvIK3VSRHDza067vY+5
XuFZRkEbsGTDpKkdMv4ZISyUPmtDZYlwAxadcSAlbMcgST7xWe7whIkKPi8aZ1Cw
9ta2ABvBJ9Hrv0gs2QjmhaiHrxpHAuvSIRTNcyJ5AXvmrwrOeDWVUbNYX2CYTQmu
hUxMIHxlmo7aKinu/Y/2rmy74XaSs2RNCLqdvdxv6MH5QQIXs6okaiWw9KjcPaTo
kHMzdeH71nMIazRg4nqNZbC3xwtXpJtk58ztKMfWerN9xy76FKcK0ied33S5LyRk
bGXBDH7GxDW1jcqF4ZkfK0uE20sL0VfuzQ8Ju6xiAbgyOZkaxglx2+DK3UM5eRE6
4q5NJMGiMBU6OBcAqueh2J2KeQk5c/wLGlVIhzACOPhp71QlMOwmkZBH7UnOymSu
lxfNakH84XdEuB73Mbun1uM/MlpnXWaf+gycReCgZs98wc6auSq3bMoL6XaYhXMw
B9N+YgVirszK2yBzTqqRe+cdR/tWkE2uA44ztq5gMUJT2w3nf/ssHaTSVQrtpgdD
azJJQJrxOkuUxhAqyJTPgtfGVCFctzsq7mn0zz/VBTldoVaM1h7bUoLeIEwl08wN
RWMbu45xF6PGzxFpQ+O3qVQeul5ajfaKvGGkThr0DaD+oKQqfHWcEr8n3gXovbPb
6hmjMdTWUs01p1GlOc1j2NFeI8zWwby+Fk6hqElRnsiKsgQsgySTzA31YOlNdQzL
2yi+f5K7zluO0CitGCdO47LNZYjHmNE6fj//jZr0iy4rvhDWdiu33PaQE2s3vsc6
yNr5G3OZwgIw5qHFJJGYJK/5ymJ4JjOFxM04mgw978dDtBJbU+kZgDmRww+94Cr2
t/RuTx+7tiPRxGFDxyp3ew3sn+aomJTJTVM/vDf/xM9LVZdxQlbbo9ngNun7p5kd
6zYgjtLvUQY4FP3DiB8XuXpF58b/4NGNE3VKCpNpuMXhZYtEdD6pFI+OMGzkCtN7
m5XJ4tkIg277RHBN9F4HNGb0wm9xfSzAXSpDDdSdH3kLYI6vDygDgWvDMM9/DySL
AumFCtOhGDt6nidMT+Iuus9wYUCiXiE1jal+h2AQVoZRehICQd41EYB9ofbCQUbJ
j8WDVOu41AEgbZIt0X2GGFrkZPqRgNO+b/cSIg+YFFItqKIyXx1FzpZoUSfQtwf4
ikO/gZz04ce/NdBS5xVYw07vOyODcOc/APs5HEv/vcAuCFSQfWCv5/CkoBZKOWuQ
YFTQXGAcYnkxwaATL4VDZ+yUdYof4wU0CurZ5+UB5d6R0tSVPLoYyCvCyfT/LRFU
5DWtRTrGuGbSL0dwMzjMijdmHhqdWzjT5TxXBKNCPbzfDz8rojXHx/QHm+Fzo9Fl
XzWNUZ9wwsG60By0XNG8OOnvSYNNbViP72ByHMyuGEf8237oiBAslbYk6IMvjTJ3
8IYLmuqdJAbKx9YgslvY9Lyc6CUa3pBFTTzYOiHt2QxI1b5kaGqtXWIFPTkn+FBs
5ODO0N6gFsYH4YiY+NK/gFSmRQ+9xOLA5QHzRotU5hoZSx7LbHCUfdWprzsoJgsb
5IZXFAvMa58UcoRE31dQMUes1pMwS9TCiOhnto1ZFvior9+05/MhdJGXYlQJa9f9
7l8EehayZMzft6p4peYrGFWRrI4NTYbWl/dEH/ddbitL5E84UvjRJq1e/Bm++ZRQ
IJdV10Tjw/AFDEcfobGF8Rr9PMrCPtBLKhpGl3vsAbyV3/h4/E39a/cOoepdMqJt
mAQ4tUEUTrNJlSweRYh+77Ki69KUtlx+HxWU5dN8D6ePWRmo1qWn8K8phgQTFDA9
7du4QutAz+iXNV9SCtTTBDloEMI7yoYg3own3odDtam/GIG6kscqR8FjKXY0oGrr
zu0NyU5hNoLvczUA1T/TRzHy+Pq8AyJuWg5z+GbKx1kYIf/nwsZOYKJb7aFfnlke
x0ESocc+wZdPZyS+5DWaxNq5ahakeeg/3/gBY1MQS/PFmrZTBmoVpjLoiMd6OmCa
Dzre00lEGzpD0SzZVQobu/ycvXqn3BX3fdQHof4gnrmHjhpCyA8QJH1uVrImMB+u
trHbF3VxoY8FOBWusg6n7Ss3AN/UuLKzVJS2jI7F/5adJWoXPys7yU7o5tlYPafP
OJUxdbKM9UmYVoSV+Gec8WS55VaE3LX6MCLrf5cww29wvXwp0ofWCvS+rHyUsXsI
yldvK3rdnwWcuvABuxbh4mxSpgepwuFjrJ+tGCEUTbMEWT0aZ42LtLYa2PjUkdFF
tyec2HKYLLk+l3a7LnmjvubQaAO7tMHiUM7RCtNfMFMTm4SrLgLpIbWvd1IFkEqR
U0Dz96Q80L5ZhJogvrwBMWhmxTnmaPExxBRivrhFjTHleID0MtJVFScpyAMKBG9l
VRqi/D7F6hVEitv0a8TKtHeJEDTp8iX2NkaTyVPCoMwOMHQi+P9maNVeFLkEK8Ju
RvRJrZC3ZH1QpouIWqzNaVPxS91ohs0lebZXHoveHbomXKGumNR6KANE/DPe0xHg
FzTaxN2yISrA90h4uTWLCKgUud1Ah9KERl9kL4rkMUiQbiyHgWAkY783bnziP+tM
OVVqMhKNvbf8v+xYRBqAS7fNx2FWwt16KuTuC10M9VBwlL+bVdEug9Q8cbbp+NyY
mKpmq2TKKj5kG7PXA38UbyVJz9MSTYmTq3l9CYcBwWsMiqYln02UPYEtI+Mll9hY
ABob8lAf84xm6qq1HOKzuRN7/+J5Z1g9VGVV9W2buiNKgYNzTqxB7rA5wX2QNMtf
Jqcj7/8oQvP9u5A8ThEBrIyg3ma57XtYSLvwYFPlYmq6zAgSKJh5LYqZP+SMVxoF
rfFLpRibDg//q4J//5oR3P7Qw98hGVN8ogoeclwB6nybIfpsFTPz5FpcgacZzKpH
7nB7j6dgCXv+RCVkT6kqrFVDbnkmp00x6JIOyKsGFkT2wvXTMOhW4Ah83Lz0Qxqi
ja3W/jvICZc5g1gLSaNoxlLauf6XWf7NWnXL3mVv7oI6khBl/MVINcZkLUzVQhXY
WNn99dYwcozO9/e4pg4++THHIZOOaqN5jEF4lQO+4RdsPIW6bcT6ZcA7uLNwqdN0
8XB8Kp1lTSoT/Ky/CqFExiwtSdu/aJ4WmEahuxAIL5FfP7H2sHmUWf4xNyUXsstn
F9L0NN6iwI1o5O0m3kqMbmajrMSOQ/3Tb2I6Tir/ny1W/Mr1yLScGmva0UXrWXtP
Q293bwKly9qd6O39N0hypnr96x47PFTlr+ILcurExMNPgW5mzjt+o2q6VxB/Vh7W
7nHEt1QEIW10buSvkvah55qOusvIU6LtSszBA4YEfr1XzasxCmUTK44S/2umQDxW
P69lnflI/mrcv9RUQXUfr2nmOj8U+7zfxq8pQGws6nFRHKSHbqpVBfzApQpUaJEE
qW+/lYxcYmoaPu92DnOzPj8Sh6uljpM3oJqx6CNNW8LcIqcqtajyJUjVmYip3/Ob
CN5jClS6/odY4Ni9PmxHpY+sNipFzvMEs1RFb1sAMxuXPx/eM3adgNA+AAuQYD6+
/YUMFyLSEWC1h0lHTXP/qxhE1P/8+IY2g29vU9WdiwBEFEDCjcIx21rRXIFDog7S
tuSHOlmlZVg/AqdLL0QDOlGiZ8SIR+b4KBmaco5+vpO4g34wXSvM/TENZsqBF/Ww
6dSRsCRjou/NdjEt9nU/alB8vOXS5FAN9RYhk08jV9pef/kBQzsFAUWonhkmZw67
tPf4N+ZRybDabt7LfUpLigPT/yckELQsP/lcD4DiuRXgu6gNl6D4/VttovRTaxsx
1LKCJVFCaJdGMI6h6fShgMH6U2qXIK/nkCZEqOISoJaEidx19Ti5z74IoWNi0Nkc
tgdXY2LsDRZHlimchIAZjiWQ+UHQuaG3jBhReZHpQPMVIePpdoQmBGXwNk4suGud
NrcVCEJF0hvr6A63uzXybvqvOTFseP0d46d8MaZ3L+Rjgw+qE/h639FqXU2V27oD
Z2DF5Ib429QSKj8npGSJyz1lSVHp5b9W9jz/LBLLgn0sO/oJsK9PJ9c2rxH+xcKW
JN8fV3KeeVmnOYAlmt71UkeFkt5TMr1xWJOcXHko9DSHMZap3ARuBcnjQJB3h0p7
s3ov1hXP3BLmMJ9NbuBOganDpPpqSpC4USf6U5vIFjbsiEPbo+mb5CMSp7Bln18N
vc2i3v3aySnndeqqQA3PKuiTERVt0EWCUzORwT/OiulDBg5qvje99/rMygZBNY/a
uga4WPHX0v0esPDR/DovayMLZbM4VXNewNtoc0LtAxRWgk7xOCvqy4UW0G7YF5pf
JxRbxQcxvZ+g6kuBpkjJh4I3vAlCDKKCbnpKZGSJgKdLOx4Lro0wWGyW9EQGkp+W
LEUDnAhrKjhL1DVyLQ2MhHL2amfJTGGCTZYJ+bo1ynkTDrcVIA9deoD2ifYtoFmg
o8YC8CwcqoZTZXO2nKN3H8C/XRzmEt5L5eItbg8AMDTZbeQvyZjs1g2wLiFZOZir
wk7mp8YedB644drOmpL8eJ7OqgbzV3R+GQ8/KdOnHlizl43xmhQTNlvf3EHlYkGH
h/p/h/7tvUEzNJpLcMEX2JB4KDRk21NCCBEMGzUvq6DELccf4gkc9RhyPH6SOoyp
1iXnC9cbg9CH5lVEe77oGOYIHNLKaKSuNrahyIUct7vZmB591Ag7TKL7bXH+m7dw
/1rO0PY2rOvJ+hgvWvsNQ80lNCVfDGCmYemWV+e8+0NjbJmHG8NoEZy+2MwPNjfS
PckmJzwXvzY+fzUvKtyuc0A1Mi0nT1F1smYS6SA2OIWAaXozwRGvOBIgIf9O303e
HUYflZjMsZICUBi2G464IA1yNFUHvzB7ODTicFJxWRNL3ddWFL+v718upCCMe+Bm
Ak3GkX3iKuY+0ywDkoQ5R5kLX8iSTx3FCNAvLBtVcp2qTv8fH16uT2tN6ZQJCgc3
VbA0x7/axuCS5PFyAh7ImYx3ZD2SGRM/WGMrG2l2VNH/DzjF2LchT12A5KewPGfu
Ir+Kh5vjdqfSbr5XjKp3Rw2fFxG9fNF/rNc6LTH6xeoDuf9MoWv21W2AMRZ7sMSz
YIZNsLtxFxQPxgir69zGcFSqQ579V4EeCAjiP2kEV5LGl8voue5wY82ltMDpmlqB
9ixzmkizYgtOdriNK2O7UqW+lAY6nykpnkD3U+vCVaRWqD5f0a4gluiXr8FPWvg3
EGTg610kZyvQwdJnv8FBBahmct1Gm7Qyfa+ikqI3ev28Af/VjRvoKB+gkUA/dRW4
9BJqxfWvhFVHomDIleNuEG8cKUrFKSn/bGmAt5ymLK+60WO8+iCZSHmmWN/L+xWR
W6cxfQfdS6Z3C2n+Z9hb70EtjH+mjNkw6ugU4esxA+aFPlAYBG0v+fYHEaay1Ugp
69ORQMGwERzYRAFaG8PMr8jfw3ssMzmQziUCqzHEdG8nnDJXeTTd9OO3959EVeso
TZ5rUEGtNTP5dQuQ3cPyQSUihDChsvT4M1fk4bOnSEeNCbz2g34rDEgOwoRyQLRk
zSD5s+LINewMo4WSEsYVAaepC0HOW5r5lvBCIdHV+Ga+MiMMHOyCMqmb8ioBQpkn
e5SHIqBUUPnVLYHbSwWF4GF4WwRQlVyEHvgzISsr/jErBhkW9ErtFJT5CCnQTSGM
q39Ft+WNeGQwbusyQwOzhi0UFd9N/8crKrpPfe26AbrB58wwCVztvfqftBRHOeoP
XpZmVVgW40GEtwHX2Xf6dIgu/PnTzQX+s3XSGlDnSOKNeDfCiPszDEhSoRSTY77C
i0UGUqVru4M37Si2rDFUBS0wBjuoHXBzNct0Yda30AdWk1D3+9kfWaQLot9Hdzcr
uajvtCgGmbZ3H0LxHDhYCYRSnGCNVYQVLZu3MpHe13o5zkCwjHuRk6ClhQA/TnX9
Wspm0EuOoV2G/ssZs3nTeZisR4r51TVByIDK2IWwclIZYyuNEon6mBPQnvQ2bQaY
Y5SqtmorVcNsrV++GJIrL77n5U0rH/lDg/BVSFx7xAOHAhsNkQhowbMbk02Os1ZU
+n+H0cf3m9INYrXidIySZsICYREWBylFYY/U+DBlyLWq5ngW3PC6SLSwgdreNjWB
t+jzAj8EsbkdGoL+OtGJ5kr+AxuSFVLtRsuqUWj5vv9u8c+z0EVUPp0FYvCUm9jr
JoATdAaXbCeAKFCh31SLIJ0Fr5pypUrmLAx7fDWFoE4urns5UHNxlcVG3Yb8UECG
BLwKN/JOK51K4N8Jzthnx4SsKmhHcRch/z5c7S+VTtj9UnRwxifbLrU5f9Pe0L0W
6NJB4nQozJKAuaoBGaO4QXTZubr3SHxYpRjBYCLtxLvHECXuhOv6SVUgzbRdjtPi
bS35b6X/y+T7Rszyptb1jokcEYhV0z+QankloBEXX3AGU3QnbH1D8ENnc3uLwv4V
DjBqOy1VSyY0c/d4unwrkQTjRkPZNVO4ffKjruL94q4ensC5ve22vKNR0q11kkDR
wblgPNYXt7B/grasZt8w4YFCrN+XCN37P8pF0AElt1M0ysTH3/OarY+zRNhlNlDE
u7M+Z1tAdqvetUea3aZp5v5EcJWXEN4EJF7g83NHHiV42QWeVXxAw2071XlsUPLo
PJ+Q8yuyOLNAAsY1v+n2IWsEXkXI8tI06KJhzBkfZwDbXm3TfDJj7L80Opv9XP2k
WmyJ7C2TTcQGI9HL3juLssiNicZihBPHFJZ2RtK36nvyQuX3ZuWVAZ2nkvuItfo5
bco2IdaYe1aPQq5Wq37vU9GiZAGsLE5i2OW/S2nYEmIo9eGl9wNCg8iXuEMMSSGt
yn5ev5Z6RRZNGP3npnbgQsZDbxWOfV16jTlMmWcibafHqgn7QGHp2rwdi7hxRgRH
kPye8/8wprE1cLgj/NZtGggi8hBQRCSL1kM6MngdBO0EN0v6xkg4zVFAPMw623tL
9qd3Sc9Zz6CPbGTqzvlxpLQFoN/gTrw3njg/9AR8dO2ju3OlxVLWe/NH+KQ9YAsT
/sVho+gNElfud/hmY6ukVzcX/LAmHBujcV6t1fc5lwhAfrHDngRXHwhTzXPA+8ta
qZMWOHXU65xLNLIswAYUUKnROsJBf7wamwDhsmvn2Ag2t7BFp/NvcZdxkXt6avJD
s6gBZ5mjyE+whet/pTRRfxsmsXZf2yqSHhS/3NO8rgqdc29Yer5adpfEvlF/i/72
vmlxNleXLzeMZ9fdSCessK93xn2/jr1ChshPTYEWB1d1zE4LSc/qTsaHO6g7TPY+
CIqMtD9Eo54uC5YHzsz0aT/nFPpFtY/d02yYipcW4X9LlXOtQ7ANB9MfZN2Cg+I4
73BaIVxAXdYTQ7+jm9eyCyYEYlrmBSDaaUHQRShGWdwbKNc3Ia1aq+ro46Npl0Vi
tcKzy7TqNKTKBsiSA6m8P6QiWxsw9eGqjKa/7NuF/GC5OF63i6lQ/ME1YHmzFoU9
WHvUt24f/41MKy5AQ6aD7xF69v9gTQmzNQDr7nEhmoKuhkMLRxIuV30GerWWBpAQ
2yAyKuMjkYCJuho1oauT+UPNmiMROs0APyrL6rqQCWF6FYQ99KCn9zU2ATsysUKX
vQLiE1C3HUFJgSWJJCBNL+OUr2JrseF/XwCDr4ajZp98I021iJcBtduPrCcprUSj
7pm0T0YdKtTRPppPrvJOzjtgcQ1tG1vYdWWdWMuhDwEhhm9+X0N4juMrKgGob7qr
h69RQvMcAV8355jQzlPXNELUcYDR2C6BfqC+B6+7Fot8W7yzhh0Egr2GcRQAXRAq
dkBl87EneeckX2PdfGXyVCxhe1ODUH+zRqfzVvdMJ+vZUGjZZ9t9RJADIzjaYqVL
GhvUW5LPtmJ3Vc5v8i+/x77yd/nxCRs0Uf8Et5CTLsbrvvCFLEpSporFoqa/F0/6
d8yMjEyngIZ2sOB2UGbh4pJOvSCOAQ9ZixOaeMoCsam4jM5iokHLaVp4Z4R1itpi
ASmzlIUXYYjtHilDMlKDvmKIVuhVDWEV6IJZU6uWK8RklNfEFtVgtZdPvpbjAoLN
ofL6qCaGsfRIFOMPcwp4ke93kFiOUIKf5PgVAtvS8emme/787b9zaytrM/Mg3bGn
tz4y35SaSrChAFQN8+JDBTOfgAz1DQ7h14RjruTiLfgS2IcvrKt6D90uEszJ+ZnU
6XqPhjtoDXSzQSLVxoAqH5IRTfTmPK31VnOK4bYWfSbTgGd00AUCuB2bxY21ogKM
EoKDbdTELanfCAueKNSZ/M+mKgF2huspSSzk7I8C3dr7tPwoDWmESNSSV0r/JjAw
ZLPVeCNHkLSw8UZc9pfiZ8LwthZ1RuqxjSd91itFEiajF1/jDxpE/uACTPv9vCow
zjZOCeXGugvqJt34clnRkwILvLIgMBPGv/LI9ivIQetvRPkc+4UKdbPWghevgMLu
Yvpgh8lwlNfnlFTdymr+rVHd1NEIPXj6zUXOZVxj3aAXeyUzocQilaWZ1dgzlJXj
U5KuSOTA8VH1ioeaVHnP90N7nOoI2Uh/HokBds1Yean531zLFMMKlfKNQ12Ez4s2
IuTLlDU6lZM7YWDXjdQohww/E2JAc734rBtNOBuLyhlltCi1FS42uVhTIkUkTnYK
L7dOHxUaFJDbPKZSwgMEPM5CIGdKN8UPMd1e1Wr5YJccppbailvLZW/YZsvE4imv
oL0A9xDK6/nnVQScmArHekUqR+VxprjCPaJlitQMJMCU402Hxw3KLDHr0MRo7ciM
VE7JW2MkEswotVB/fjPCoe9qUZ6bJyomRYhHt+EDT+mC3Bq18+3xm9dyysSF2zsh
+TjxeVv3zJI3AKNMyHhiulY/GB47FMFkToyxJEHu5r3D25k7LpduFMyzigY1wEsd
atMqcxmMaw2LT42jMvhyWgBw2Uq6rukiMTE1B4SKZ37YhZPNuYMIERSsHwPvIY43
Fznu30N17OGazfj3/NV5n3LZ4MtYwbmZWkFexOo2/iRRqPses8qx0P8IimBjgsq6
goI1C6v/x+gJYnJF+PfG7k94LX2/zs/xDjSkQMFGUvOU4cNTfvtpo3NibxudZGrM
+LA6OD9FRYklgVjbT42R2/LYuE0zG/10n3DvThUpBF78i5Jul0SSx6hUkU7+UTyj
ADY0UL9t+gWoXlSwo0C/QUemy40Y5bfIfB1jcsKBsIv9U51GqVwcnhBS2b/4orXC
mkF0XpgvXfB7yWLc7fWbLPN/f9KkKKQpfajABR0aeOGNYql4Br2buZm2b+FY1zZA
w3dc11wcOm1DFMUpNQyBDDXz29DqljkZCeIWZVB5b12N90ObD6BuK6ST1QdTLesD
OBDXnLYzvDtqI4R2Ta6A3ddDhSzed+99CI3gxHdY0+oZ2wKFNZnzS8djVNmn9j/i
myoGWul7iiw69JtnBvXXjMkqELh4xZjUZA1bvlhNyhaVmqgTEcjd1+oiCFe02bUO
xlu163HHHUU0dchIRWthN5tNDeEahtGFv8xKgTl8pcJZ2/z5dMk5gMD4LCrMJDF4
MhOaCTf8d9ZGvXHAepT/RKnTOMXu1cCdnJoWQ0qtQihft6swh1DyPqd8A/RusuIl
N9JyeuPCeIvHCb/pY/it5hGJyldYkKxZ/75b0eXD1cWEJ16gJRdpRngagyHymTAJ
+s2lgmRi9IY6N+XpnWnprAEak0KtRONJJryKBt4ui3JXyhcxcRZICtjVC2v4k8uU
i7N2AyaMMCafh0ZZYOawMMUqijVl1KOxcnYtKMZVN/ILuNm/gbMEiFNTwW1iMuWX
8H0PvGEAPrMmhns1nvnlktAMD0pkEocGEohgqo0MVolzuml3ZSh2T81XPTPVFPp6
HwJwv5G1W6B8DsDmlXKLMfmYELRzzjN0DlCqlUCTzpQXyOs+cSXzldWKnQIKQnMj
gg9mq44WjknKKZCK5kiKF5l0BF0l2Ab0ksk7cmKtyBMwlGdaHUoREFShNFWfgaao
MkvtvhZiYW9Pgqa2WcLuWTRif0vCgE0dp8fygztQCRZpDjgHGYpGTWEJZK6xdLdr
KxK44xmnk3btG/N7fZsYQaMvRwwOEvrCf7N5u527hJOCmrVuGq0ReQ847r+kP9vU
aP4nOjJSgGJLjRlYIIjHYihtQUlmhODBazDCwXJE+p4dvxELyP1/adM1zH9Ujb5E
prac5pjm4Ri7QI0s6pQH/NiM+9EYOVCxAASXXP7e8AaA5DBjov+04jLFz7M8PvMB
fBHCrdPrFZUVYEcNyyDmBbPMCzTM92eMGQ5AZRxRT+10wjK+low0VFWFhKRk4H8F
mpyQqGVmlQuyH1gOmV5hIYkaKS88HdcjvzW0Jh6xCJFLlxJPKygl3nymZ+CJOadl
Z9i+6eTDnPnjUHhrS/qxWQR6tGp3iaD4/nYVNJLSqOoVUT6kssYOem+ABHuszpPf
HYhXQKcCrPkhGR8Y09tqCsLALtMVBGcI4lGgRGzpeupxEJC+aCkwSxmZwwUC6u6D
FMe7Iu/x+5UuXoRM+DYad79RyXMygf997MuKUTsxXZFvHd9n7yw47B44GGqftV9t
XZYtQu5VIRkx+gMWoUJVlDZEKXdRK5Gs2PcO9KFdbtiwJyOrcVXOd9VHIRo63Yuw
XrYWcaowlPh+ylLwL7c6zUyJ/vytnpa4CT1GIqHypO4a2vUs248DAsjhFsyu6Djo
ctMb2TeXitZH8mgvEwjxTQr9T4BGrAZIij6ZWnTcgwZl4TZ0Ni+prqmRjCvgWxm2
s5P/QgvF0uyju28Q3PkkFoMfPhffht7rs3l9LSjXKrJCwxlmoSvCASGm0fnpoK/R
jh4oUuHXGyLFh3USo2DlidnG9Pg+ccmyugvIlnt+EHSaUBN7Sz9xWwOc+fBy09GK
cMeTr8hRuTPSxwhHWztxmhVcgUDOhK6vKIRsboN3WrO4tWieeqbx1zKdxa/RRZVm
e+at97KC5jo+oWYP1HL/VjlPn2K9Ra3RKKo+0yODqJGbdH7hwO5BceWsf6fTObhc
v09FPePW3REdco40DdJ1DnFnGaYpAwd9Ibbf5ZQHShqW5V80ULVhzFs1wk+6/FAA
Ueb0T6kJVaV2IdAEjhWj+rFcICF31jlS04i3rKF/TNe8RZr0zQ1v8AHzXDyUiWV0
s9Hhfpm5fjWXr+ZrWSWvIVn9UhLYlzCp/vIdUXIjMQvRzrT8VykqYF3DLMSvGIra
fxyYW92d102TtX9JXpQpjz9MTxAjJUIy+31YgsQ7ZLjWU0yYd2KDgzMdC2hpyt3x
/MRM8FjJebW5GLLKNHxLph65rim9Q1Bm5lOMILPdR5TUfNWo+GPDrwG+jaJdcD6V
Ql3ugArsfNdNo1jELRYL4VVLq+ZuFj5KV8vcvVoYh0TixWFexFCvyJYKV49bRgFa
TikoslYQkpWp71MAjClfYkS1USW3Ayn0R1++Xx0A3irQIBcmVeSwdey4S7aqLuiA
BfuRXPkFZZdeuIw/Eg6SC4fCIP2JaP+pR1IneN3wCh0h1Xznh/2EnH95CWTIWUz0
tx11+1hQipSxHFAEZmbkTg1sHeRw2djx6tznJUJmNJ0469epuk4dGQOCHVJ+FsdG
70W5Pwf82rD0Kib26weClsZfEYsG4htJ8NGIRJFKBy5wQyEZ3PzugEYYQNJaeCDr
M6x2XSVJTTq7NNkFwIexpzFckmW9vkRhmgDNHrRxwTvYLYuEUecD0lnt8a1ItNua
d+rL71ozsVDySXwX3F1PX6lBtbbndpP9F11RUYmCsRuptkLwidsBgEwDg9S7kcZs
e5s5uSB2zOZse7DLIZnjJhZwLmuP3xUxsQgyOuEIb+nTumk5DrF6+BA6Ln2YlDIj
+wTWl3F40ByRLuXcDqHym5Ihhh9DLZM0Rf8bxDHcAkfJWOzyoYgWGD3TECJxxtrx
l1IF5Tal8lQWzoWHbyIJAvkHrWA3KZ0IXZGJH6SH/Szjcw5OA1v3ZmrG1CylUplm
dlwjhFcmTKMBP2keIuRIB5Yz+oLAoRrQNcOMn9yoW8176xHqwGjv8h/DdyQfG6dz
WCz6VgwGFg/QTyMLDVN6ajb8FuoTtKT0KWm9IrDp/1IwoxFZFByz2FJozSLVGsy0
dC/BPRDcC/2m06ZQpH37AU/+/7QuACCx6z9Qe+nS9AA0Y90bsSPpQ/IXIdG1LZap
I0gpBqKRBUROg5zKrXPtfdLhRgigDuB7MZ7FxdY2kJWP/Ed+2iU4qXS6J/phSssz
2TP99iXk5WPtswkUlA+7Nsl24CrNJQgwDBPLbWAbUG4azDQso7ccEgPJjby3M3Kp
f7PZ0+GmVMjV0gQNo9ecJXdpo40C3jbvIK/njAdraagwhNVPAhSx0fN9OxiTT4u7
LKHKw4qOnTDJkWM8HsCgfjJU0Bp48v9ugl0dAm7XSG9Hhnq7JWIVzdqmzWHh9JAP
/N/ujSnDKEqqppUBhGUH6OYC+rt5k2x7XZUzW4uazPVCHMH0q3fWm8iN8X02Tkfp
+hUGoeT96/+BCdx1AtFyDEyDiuFGU2aSxk4NPs+4lspwNFCue4i9pyJKztn1HVG1
BomfhHyiNKwlutRU1nf4nZqhETKehwTIZ+RyCUo4mCjpYxoz6mYvJJg/utNPOqxH
y3g2f79sxMMPtBIodmyMM7zn4++QurJC7+GYovsO8ugaTTqbp67uqoi2/9QdBqWe
/4eC0L583xqYO9pMInviQaAVMxG1QA9s8s7ybuAwgoy+9kiGtJGOClYwBwfQgywO
hOEhUvKLqDhVFHFRvgg1Eu3hILkYLxHrEADcIB3pfhEZ/NttTYxgYOPoAqBrPjn7
STle4NFi1sNRleqw5IEuT8d5QTvJeA0Ocf3TxDGOol75dB+ODa0MRm7IIblZeoNa
DFzhXqe2fqSTS7Vf0nNJGXzO0jJjjrobphfVhv2wVov6fqNBYuBFxq96Mam6IXsv
Gr2r/RyQGqVy7ZmhEyvwwR3LH8BReAkbT438KauAM4bUSf5l2JxyZpyruyALIPyM
T1uODsOV6LDVhqxxX9XqZp46KEusTR9VvDCCrdjl0/qtGZtvZSrfttQUbSPLxAQe
LWQ0Gg2TDXwMu5tcKoEwbTKtTEhlI0y0u9FDwfscrDaERrDaOubKfWuHpAFG3fQ3
vFINtcCvQKLNM4XmL/OjV8y6astocFTAWx75Ez7h+rwxfaNoxFu7WAUjkmXhLIHy
WhbUim8tcR7iCGzU/oCDqXfNDqIgB0/RlHI4dhgWge0RmhqaEshcCd3fB8WXx9pL
AxCvLAUk0U8BhEMZLZ65L3QMLa+y9k8nhkfO5BLiGjCGTPg+tWgy2fVZuTMQzm59
lYWf9sTKHiyFmRebOqQa5P9m99ek5eY/r1EIkPJ5BIsKvHTec+mxCVA8dLUPvJlK
oGfwCNoPDZcSrAdohCnhzY5RFJGfW73meE256UxiTXOOTiIsb4relM1Jyuz/GdQJ
NU4Feh/peIsWWxraAkfdCdhUK9dEQDsN92IqMf0XTpa47iZntShuxCiFr53fqn4M
zEomhpPbUfOgNVApGc7zk8GNWAwn5D1YMiPL50xmK6N8+j7fahE51bur37+OoXlf
Tpggx2O39nJl1hOUufaXw1MnWhEO7ISVp+SPMTs0DhJrNiZWtVRB8IJcnWzHH7CR
9uZ0SK6QP9rW7uZjd+alltX/E0snUgbu9dJWWr/4nqw4bocs4nvlHShFT23w7d2P
t7O6+qOSRfqdlZ0XSR91ABPvjEfEaLMOn/GLfCfkgOosCliVCyAfFixTaDGwdqge
9Z0QgBYSCDcMEGKZYXN1hye3yRW5wIu1Imhlj/sH7+1pCDWoTztB9pXe2D1BRtsy
9h4ObP2CWf484tGO9WxweTZaAWITmYr1iD62hpcklFMsgIliLGvh+5K/j5Gkn3z0
xgx7NdGVugZLi3ukKWbBOcVhDUgZq6H2/T0+IlFZU1uEEM3NcgVcz6KJV+8rY7vt
SGd8DxknOyvo6i82RDsGJln8dSx3lpUnbbP2kgUsTr160TzVSig7Rz6bUl2EVcUM
ZEnsx/0hzFu1aS1QSgttQImhJecBWTSGBQRs7l2pdCAVGhkxy8OCVgunKnJ5JCDA
rVWZS/zQYJeAyJhEKzkUulZH/kYFLEo74Du5PrPlObalcmarbkJpnCx6FhsodsaO
4IQWIxlk/k02kv4xmLD2E3VGvUo25R1hZM4HNZclu3o7QMEZN+TGUHswjd/c6tf3
rI9vUYxcYkYrhX9PAMJg4ceHoWP0gLltffnf6BX5BBs+Gx1t2JCcaupPDlPHTTLd
hNugVZ1OZ1wc+iTCg1M2qhxg03b3p3KpacfqVLG6W5j/dIHgFmtqaUOkHFUL5VxH
1nqoalANtqiMKGy6Vwv4mmBTUdsDcaNDJ5zjwOb4V/x0Db3IA4uX63aZyyacp1SJ
LeF/hQBWSIU7vbctZjGzlJe6oSORbVHqD9SKgdjBEMputK8Od4PHb3FkyIsGa4+j
xM3f8oO78lw316TRC/d8WELQK4izDgfUMUMnRkjPVmcVeFfYKv4nR3jzTXY2SJ0h
837W5p3+KVU86K3nWbrnZnJPz5teSV0Z6JF7nAFSaekSfbAJBX+uLBBmNxNfCRNf
+vJ+Vbg2iTsbBsK1pTQ00LMpNYU9GC1ivZF2AcM9rAzNOl1DIK3U4CjHZFMfxzi1
IO+o/ShOe7y2vT0CXmfPECwWYT2cUB6g0/uhLwMNe5YJLmWVGiw+sVIQNYGgK0lE
sLcRaymuAsSrgMU4JbHyrDQPHYw3re0WC+fg6psHKEFY50/Y765rxqwrBN9bZslP
0m34Wx7hufW3fXLkIcukZSlQAEyjUHcQvs43wF7GCJGAgnAnVApFlZX9QXScvIMN
cX+CWRGGe+tIAmEuV9cCtmGUCgnDLXWXX4owDJt3OUXPJkavacXl7ZqpqNU/six8
+irg0Z+Vxc4SbGYyM3xi6Zrs+ZtP34ECD7WdppZk0mWdwyYyJISchHlwfEFilzQ7
f5eUAyFJtlb2zBLOjxDY2HJ6aWWvHjCdyuZ5qoZb38JtrlG44N1QwEQgvb1zGbOT
3qjAIA7b0o9+/xwLPPN07Tj4HQVjmO5MJwcR99Wm2Q/bkw57mc8xy8Yppp0FLW9a
iEK0GcC68OvHzsk8SZVGlL92ElSzKrM0d0vVucsK34ijGYKmc5POsUCH+agdUhpk
kqmLr1tWOrtr9U9LUjMwbET0/cziG81o+6MSeHXK8yY8TZF71WvVTEI6X1Wb9A6h
CGuIDmkL5RZYH4x8lfPQu+1lWGqowPzTEUVIhuY7GCVow19aVYZCxL0ZAgKWLppj
EPvPv8+6yrcZVxIr9YUlWx8K202uAY4F5qUgAE3Sx2DaokgjuZLPthg3XIjOQYUJ
Yr4DCypgmy8QBMq7HkUsccjBcuIRThJloB6DKCqJ2cR2dL5SoeC+wd14V+SXHGA3
ZQw+BTn/LcQq8F5ceHclyfDrL+lXeTKN3GhjvFS0/Ed1ltop/IpvcrwnQ90519WF
BNUS/oOUsnRXWlth3wJABFIIZXBU1FMajx0kyswzj3e7yvvVfOwNHW6bKSVyy1D6
7V8MWdawL0uN6oX+oNl3aKotAJC9YZma9uyAA/UNLIcsC20uoS/B1Y1r+TzjGxcn
VribHI/h9+Jd7oPZhGQJA8EjzwogR5GtkZW1SEB/NBB4pKUJA04jymoKtVOay7Mf
LkRm8praRUaS4RXOn8pXrC0pB6XRgkUQOmC/kbOa+v8wGGhhJAFjsW0li/7sjTo/
sAXSWWpgGOSdRjvq4xaC+S44zNHRElGbzf2r8flx696ZAitWIQOSDgIC4nWswgj8
onvbM51FjMjBN8hyhGW7jQvFPkXsRx4zXMbQ3mOxiXriqIFSk+fkK3KbuRkgs8lq
RF/tzbUUZkTuXU4pjrigNq/cG5jILTZ+N3kAUG576Br9X4zwsXrYEqt6YgWbKrUE
UP+XP/XVETs3CjDf0OQ3wdDpyZIKOZNtJyYnepSZNJmXHnjcL4vv9TDRSDLFtq5p
jzF0EXehCmSQInDe6649rPx1yUDw5ZNHJr1HGDjGjPrlzE7bML8Pl46ZZV/nLNZt
n+gtP54Yu+a2WaENBD7YOhPVUJY/dpln8G/oahGVSZIy+DjJtJliLJDpwokyyhbI
CKUOSqIG3e8kZVjOzBNJX9/9y5vvFoGCGbmiz45q9+ZtqfXeMCaylrq2Whfh6ItG
GseqlcU88uXJvOBn3Utgzc/c0HfcfqEECJmeIPjoErgKwks4aiuQufLXiZ5YZPBC
MXApwOs7StQbjVBG85TQQKSbofvLUga5fl7G2DaTrKfW7ncWRY/iIjkZIH14yxRq
4BXtPVUD+MY7LFp8CtrDJyo0G/lPsGUEdWV1uvrHnRG09quvEvfdU3ZXX11GdABW
QJPfDssbOq1Ti5NSV3ba+lQ4KclFowV/fNeYkkyxMnu4cYkyfpAQRedA/p5r6/e7
G6fISR328bzCK4fki+WY01jCUufbMam4CEaMpJwX/TMsAqQoGxCyy0FqStYPncLb
dkRtumkNpcGzBBizYlnu9+qQSB2kAw/Uj2sIiMaQ8IxwNB/le+gxUByod9OnkWo7
UZYnfyHKPTQMgHWYlfuTvOi5LHPZCgUomwGOtbcRXV2mzDWp+x958r3U5lbkcM35
1A6MXnBtAJPMtRgLElrNDqKlsJ/iILfhzG1qLaYwhz+sBLryg6FwxSBKxeVQswXo
qaWYebd1mgs3Cw6+I6lPxJnTjt6J7hxfdf/JG1GPbmLCvZkfg7St+bZ2GepR4eJ7
uAqwbmWssMOcYrfjc6zVtsD0Ym2/1X9YbdFjKOuPxZyLUn4HpCc0qgJ/SJhkhB8T
Xjf33QB+ajF9hCry/tKaZvCsQxYDeLW9uDKZ8e/iMnxhTt400I/3X7zhgZvKJ/iG
oik7f1tq6IjnxbN+fex/HD9YM0hcksc+CM3opM16Axw/uPUoAsGlWkAn3jRiO/kd
SseNhfcV7Wkb0/2TYkWYBq9WuijdTTZzkyAjt26SYDOWSSUycwVEqufdl5STXtZJ
0uHKAb5henwpnP8AdREemtbUYrNAXQpu4e+TQbfVbuNj6GqKkd03PT0ADwQycT7m
nbFpntOBn5WW9e4jO8xLcQgnfMjROAmoVV01bbi88O0cnLuPYriG1A2mD4hGawms
oGsgbrLviMEotyOkF1KtTBd4lFELPxsqclMjCaoH7Vr99PVGbqKae1wXNePfMVwQ
p4V9+EQzO8R0nrrDUtqflOYSuqtTc5L4lonOrbxk9qqZo88SP47RW1oaXbzpkr7+
0lKf7kqaCi6gHO9T8q1TBH4PSZeJu5gTTaUSOGDBSYtE7Oa78lQ35jiei+3OV5Oo
BuyKNnHKcm2vUlJrq5iI4REZKLQTMuFh/eRi/ybHuZR5qft1u5LJFDYDownk3XoF
ZHRVbCHbDUnGi/4eFF/TrtzB/eA6UqPnnuTlur9pRB+tiXqwcFz7RV224a/SadoE
kDYDs05OezLBWWXC+fgjG4RHTQkfVtzwpJbioDNsZNRseig8aj1JQOmssuzq9wDr
cZ8dfNpnN/z5gv/BLq8xyx78127627Z+9kZOj6h/i2tV8OlIb3j36miW+tUWeNjZ
09ygiXcnELptWNrBhFQu2o0JN5OA0Cz/6cHty0ph22k2MUTK6O8YqJeGqEa6IkdV
/J7MI9QX2DbjGUvGIwexDJKhBjRrlKmLcMEmREqRX+0uTyx8DEwwdb7o3xwL1w/8
WDGQ1YErIzzUAAWvjvYhUEf9V5DqJM0QqWpe51uk787SHHAgSIlxWn4XMbfxpC61
swYIbelvaE0noTyUyVsql/h/6n+dJgBE9kOR44tWjy+HsXLhn3/pBCFuoVUKFJ5k
hZCP7gzsIXv6e8USaOcGwGTFFFv0Ba3TnJj8M4aGutdKNKyZHdKEWkwKNcJxrveN
MQzz1VTi1FkCa7PfVbGgbXS/gvQvtuD3Py2gp29icKjiSbBiewcUqhiLccauuY+6
WM0gnVwWsvgLFuMjG2WYrfg5mZqE11imNPDbGKJZOrEtcQb/h/mxe4VHrCZ2Eq4x
/1qrIQho9u0g3VIHpuVZNuZ6AYNgT0Lr9bpveMGSA+tzdXx9WuGcsvs/beqc1eGY
amuM+48tKVPv0Z/9fu6dUOikqrSL6u6d4eKm1zdhbAcUbvDzIEVMWLj1xSlIZbZ3
/8kOgb1AW9kzPR3IfSUTCrlx6yQlAYYadJx2ccWuN7XUrTBkc/R0oN7hjjbrQQu6
ln582Aip6MJyZ/mrqxwuih3RamMANlYdwbH9peZ7/gPPOdxPtwwPKxIMgtX3N+hT
lBHfJmgV5NvroIGMiTzjeF2KaW+1pOe0TdJ2uYAPDN4asAiRWs650NzdOB/a/0md
PhCuF7GeIV5VhBYvRmOvIwzE7cx9XNOFeQi49g3aeF5fwZmVb3Bp9PE5iKaQ9u7q
dhJwlCNt24I4vJyIqgmtig0DDSb95w9TNJucCdH5bh+XRC3Utl5byJa8SitpwAUR
ur8ub+K2LZvvC08FyInDCoaU6fyMaNPQnWgsp0OQEZcOnmglEykRiYvV35c8vocv
3BVKJewGcaUAUDXls4aruTilJ38hQbw7nlfrJAv6g+zH7/ZbqHBeiApULzKreJTL
jm5naeLXyECC8IdpQQuf4whif1mbbyVePzMzblgsNrZpvaFbAodb7EtW1pjphEVu
hpEmqqj6B6BUbas6+GW1oRoS97Qk1y4gnLrwoxBgTzf7rlQ2Q65Zk8oqQ1IxjsLs
AyXhyw8yex9pwLEARy1HYkZfjbibS5QKYWYgQlbQ15WpezHURwNXySBIrhCeOtp3
6LGk7vkUmtR9rbn9NlDg8AuPR5Ph1fa7+6UKeeej3vlnMxG5EKRvYSWIyMbVdGzm
FLWqxYpapdhcxLyg4PxmSRBTBcslY/kUUPfA182i+V1DQm3k4YbZ160ymZTfW6tt
hUzYFiX75tZj0ANZizTq/LEox5CViJgmxEj9fzrLb3sSSTVOsKxjJbQYhqPpjX8j
/sCdfB3K7h3mFKVwcZyoRwAcnGa9u7gczqFKWWvZpH6MD83W8gF08cPUlC9jlIyQ
xo+H5gQGFHkIrt0+dX+OVKtRdgJBqmBFPnlxzUpLLMpHGQbFnIOtYjblutEIQuTQ
igCkh8JZUJl0YZfgjOYi5YhZD+YkxuEhmTKbVnmn3bxG6112ihsxz36G9L4iWzR7
3zo6xFSXu64RE91NZIgASnx5J+aItVxgPFiv/C1JzzowNf3+Qolc6v5KxlC6h7ZN
mTkUbM2ahwm5AyyC6uhOzNTGhTuONV22ZOkTPRTvzfiCWqaQlgXyUlv5JGkWdTuP
CrpmUH+S3+nLOyn2bi2PR0XgKJc7HutuSYwXl4+3V+c4/qyyk45AfGSOzyHU9t0c
tmaL9iFTZtBLc55tCV/+kSNxLxszYA64dyfEy6YP+hCupRB5yjXMUU+fRCanJzV4
OJ1+32bWWyQsjZ6pAkUTyxbr9u3Ww94zCgYSkC3HJ6IuRIJjHMzBVjW3ijgbo6XD
B5j6BA7WOpQ2HH6FV56zzNzzNDNDzGN6A3+fzVjn5R2Vzqml165WPuw7nbEyWSSl
pd09xJ9Pl3qBfJzuiaUSPKzHDYfP9rCFAsb7qaMLf7m4yLKXsKJoyU3iINxAhbIk
wPiOWwSDMWfZabpftBRb8FL6wGJRuwAH2gJ8CWLWYNloOV52WwkasNPzBC5OuS2t
/TcUw+8vHss2+Kue7ua8JGYg705+qgCtb0WNeHpIbLdBKDWnlmMoIVztrvwUEjKR
WwJ9t0jyFrWJAQUkK3UewpFppBTk7cxPZT71zZWvm3Cc8vckPvgM5C30LYvFbfn3
i17lkvyOMiVhRKPjRGEiHpVgyszfjzry1Wc99yXZW9HxAvR7hrDpbuglQ4ya2tE5
qw+cdiruoMK+l1QDOaXhu5TMnel/0DqHDWoNvdK4/2cMyRhJxV77qxCZa9Jd82DY
Rn0wjWwznOpTjUD5yA37jTNVhmIV3HNN7houJEZ7iZaQdlqIwQOV5hJg/LLYP/NK
ggOqlEIlLyXtk4G4VJabB6Rtr9+e0e39QSaC/oBlhMUoQRlYalJu8rT2Qb6DcGsJ
PeO6SyO3Dyn34dDCngwcW8mCSDcbwQH9HK651TKK6sOFjnE9McrcZ2qhDKPAClci
MJQGw4tvtFb3JlFNcpTAa6wzQ43VApxQBqvNs7VaypY2TZ6kmO3csj2EJ8JSzG/5
FMzjsktcPXQSX2Wf3WiCRW6mP+LkLC3Za62E9sXRpRX5asENh1H6KACwp6la2Odp
VD42N2FqOk4DPscEOsOXuJAewmTEErPF3DO+HxhklwpMwVnxtCFsKpzoD9CXlz3H
7GVzZNp7eF0ui/RYIL5qgflhvImbwtvH9aNpJq4NlAd2TAXFkUK8v98r1UKoKadf
fDZd80OTk456lOukcXn9n7hj4mqhCHqFyOO4Ixo4xgrf/MYm3Zu+IDyYSPaLgThd
ivDJ25QsYlSPZoBEp7NjN5t2q2vPgzD/trDTBxKrMlcX9p8etfvg9Z9FD0i4U1az
Wnv7BwjqydlPx/xrohm9LAdAUoXUooJZq9CtkuqFVg2n32xEbrW1rwxWxzRyPL5P
Eqau29jnVD+3Fc52E88GigVlHzTRs9wh1BzA89A2hrz2OnYjkTbjY3nfknn8PO7I
ka67WyoWL7JJ5az5t1/ICIW/z6TQzkRRkT4PPrM6dSn5Tr4Nc4GOQdtmd8VGAIYR
h4rQmlNcUALgkUYhOWvlLbDva0QTCrdPIwXwzHcoBk8KnMvL188+P6eejd7Gm1Jq
B0AAQp5FU3CRxsi6kBIjpdBPB6WnhP0t+mcU2H5muKjl/COja48NXxziTY3VR6C4
TiGF6skIXFbelgq1ou9GCIeHezzcCPAmmhZuEeH1qVmU3p2JAhjcb05vcl3KX43H
VSrkd/eCVgH150OMpUofvbhiVZxj0KGUnr15QM0CgqgFkWue7UU1How6C9ITusPU
Zo5xcewxz8uZjYkTbg8TOV9VdLPJ90g4YJOo68pY9iEfvag8a3quKVmlsqWdSomG
JE/bpFZMCC4v2khjUg/A6CrXUdooKyDVXMVXN94X+DU/hz385ODLuxt5qVDhwVfh
n88Phf/unXpHt+BSWLvPctoUbh8qV+fQ611uioL/jIzleQUKhH0uFm5A3QDEzwOv
TnVejls6nZ5LKsxmVCT4N7OdFkqaJeWCONapoPdQluP4lVfaGde8kp+g+VZeTgBb
QCI8N3vKalA3s3lpVcNdB8zgWhGtXWt0qEIut80YUWPv/IbseDdv20F9e35/5h8o
CaAo78EwGPYwdl0Y+4jHq3YPwyDeobdr/HwhuXp/WK0Sr65FLqtzkB8XnqwCn86E
nee+s3dzbWabuR2psJhgxzhkGqTJIaOm524lTESOxLPssvgGnECVpyhJ3DaiVEro
wOkOpMSkw44pbTBE7OgHUpP9qjMDYpy4ygts2ekDmGjJPTP5C+T9ZGOzQvaMzwle
jpDI6ajo0f6K0Gv2Zphp8NyiD8m6gsatbHXw+gBaCgY9VoLdCq+wqCR8GJzjPzKr
pRXBihBbx21pRt/e4b8Y5qDjQ9a0uKNNoYRIxtmvxxBr/Ju1A5CNZfJrZOF7mZUk
fF16wmqn8qD5BJa2xi0mOs1O83bErnEP8qS2CvA6qjmQml1nvoXEaA0quy+/ANwf
bmL+JplWRkkM31e3xqAEV+T8fqt67qlGs7E1+CePXQUpbycdFUSdvQ9F+zzQ5icD
7M35pNHPOdAbloPkAeTUE7z7zr5lbJ/xmtKr+Ev4Tglz19VAVW9JbQqZdS5eA5UT
SohZhGPJTv2k+qlGRO7aezfw3jIRA9tHtkklrZXGJK1LXsQXzOlhvCnhfumf6NNx
4T2nTqp6zStKxZAuGNgRSh8EG41AigHSNLcHeMwBpRLhjYRzk4C22exvwuofpetB
Tn6xOAzE4DghAUPfdRAyIXnt6rw4IIRhfaakgW3mgEfAE5e6tuAWgAv86anejIBw
CZs4BTmRE1OMFTq6GCAhFKVV6E/iw3OS1x/PhDl57pSnglIlCF3LesLFlFcr8NsG
28jmK4AmUhWOdItkq+K4UtNEVL2u69RTK0PpqV80q4sBDBUmfOKqmk4auPDKBjBg
OjHS016/D9wzB1B5XuTqwzJydIpivvI5QOhE4ADNe6VMxg6Kilt+RI8g099GlRGV
2rw/wip2lNqFU46V8oul90fBt9ky+NwP/iqj5j6+MJ5D8yr4NcNI3I0ErmMjuFho
B3VnaSjFMxutw73XsgH5zFHoTwTX9c34NuDezX3izvaI6BGMFMk9BROzmHROturH
DHM3f/0j4OJ0JCfX5RaOC8dKptj2J0E8LYtFmb4g/1k+2amNcdGgPyoNdo0fnQln
g8xydZhbilzow5SBOOlzyAmA+7qkqWrMA7mSLOqzPT2dATtvHgd+JACionyqQdl/
QdS9bU+srYrfS8bULTcyzNJdGW8c7Y70ACrUTUkFjFuCJ9j7x0L/zzwVGNiGKuSd
2rwvvdiHdqvGPJLrWq5TByGaYdn/5TeIMXsJ0M2OsAQ/pTZrm+fo+FAtlLjq0AgR
iAySo8xtJrCAdh1fHEX0zzd9t4qPzYpcLlYh5+JgK06elJRBIayZjADMW9XuefaX
FZE05DytbKYMr3Ln2XyItJbb2KiInVd6r2XIyTKTvAqvIJDU3q/9mS7byBLtKVxv
cK8in1AgFn7yt8b/Nfr5p+4ItCKtOk3EzRaUky1ElkQfjZKoN+fI9PJ+5mEiyaZ7
dJOJtNKl9j5oR+3P+vMBD3ZN9+wqISBy38wc+GDza+iM0zlVn2PppkWO2KXT+as9
bNWShAVMJbUxefgicn/3DnRcLTuC4fVsE7KCElXftXnvQx4xDBawKsJULM1Pu+3M
ksgoioOuV74J6N2Ge5n5Fa6fOijt5rJjXxOQcv4d55DG08rmd7ytEgMhnFIgGxBF
fN/9TzvADfY1vm8aVhgPJ9j9ikouhJsYB7+Tzdu9Pei/DY5BqbjVnd4iDNM5aWX8
YCZGYc/nwns4jN1ynrAgfSO7xT7uKMQN/TNVSDtraeYapNR0Mo+pD0nKjKTXsm7k
6CyI4p6EL6m9Vz0IUCScivvTH/fzJ5kNGYy/b7f/HXLOP6MroEWXdbZr3PmvWdhY
CMyh5qbeZSpRXVzw4vNH1mfkUzdXRZjaYReZUMqUQOMfrSu7bCnl6fG1fzP20d+3
kAj6Yv9jg7OgeV1UMbj670R2cad6yLBZQRo8h2FRNDz6fIaqyGBBRZovQrEhkCwL
sFd4E8X5A6fVV6NoTmEizvUqUTkF9qm2Jylo0peGiGLeXuDTGF1S3qGPMZBmRwCy
MjZ7lyE8+RdSE5X4OI3NZS+Hc71ZaEwce5QXkzZ7w9IqttZrUAv3eIATlcJNzAhV
+PNsz+j6+XVFDq+hJ4HCQm+M9Y2d44kbvixCW3aDClWt6VNg2//P96CSTrPnya7V
cxWsNhMHlLtDqflr81MdZk072vXDgvUR4Sz4JmJtPCmQ57onke/pWp6OeBNNZVuy
wpGnoD0pkmRZYpnNmLB2LFukSllWpH188MRr1Xka5K6/rrST/AGjTl2VMe8xsBOw
kR/41bjyQ2+zX1TpF9qfLXYGPgohluh3m2+2QW/jfNWy7P+Lsv8Oy/VMD/4NMhDu
lLFvo+HiN7BqEpV5k4aJ/RXNL1WuNHsJT6aTD9C9v6C71SRbsv25vjB5UDD7O1QS
eGaha0U4oS0je4pIQY1d2ftfsviyapqTtlyRCZ9OBa/YbAKmpQL86B9CodDdrcKj
U7XEo5sq0i07wUlmE0Y/JkcR04rR+Vbcw5Fdcg14PIZ0uDeAYPR7sfBa6+npcC6J
bReSHppgkUS883RDhlKtjx0NKY9vtCsBIZYQhjnyZ3pR4JiT0oBjnVY/O7mwXvG7
sqiD/F4sc78QHHzQETXxk9Rsj61S4CGFIBd2VLCimeb5ZiCU56n9SeGCv9gSQpCO
2Bd5f6QQsIST+nKaiR32m9LP1GksWbZNVBrJMti6aplP5p1ass61xmxZpvqZpBJD
f8kgMffY3ioYXwsGZAhgArsb9gQWMr2RCegM6KcTc4wdqx37YmNiqs+O6LYgWBJm
l5+sA6kT0ieEwlePz4JLvdpwOOWGaj7tolu+qUeM8YM=
`pragma protect end_protected
