// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
plMWg5+p+vs5U78iVzGJG7X59S2RqvgEdL/sGqc/E3hMbBqWkzGnrjKscYCtXgqH3+abcsjmy67W
D0JGTPJ9d5S1kAK4CmqQf+vXWbd0n+kki31NRi6KC/2G2yDy7mXHCl8z1HDe1Cq+Fo5rgNstVAy6
ffS+vF/zPxH8Ykyc+kZCeVVlYth5suxjpdmYjwzajyxbISfHFJJrkzANSfI3Skef9ClerW9/KdDJ
rSg5gmtZly0RUfqw0uRNMgqZADC8nUgQnefsYdkfCCb0xyJnmu7n/tLrSVoQAIqRtxH6QFsXzBGi
RZZO6wR25i+NT01Vpk1w48NpYewiWHuBnT53pg==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
ZtRZAbQK08WQnVWuPev9DraovnljXDfsP6WqDF2bCOisdxxLLR/yJcFSRX/RmI5vKHpkNhmXdo8v
O75WeRbTwU3f+Tlb9LPAYOnpTFqlq8r1H/IMkLzKvRR2gw0QkjDZjUEfIPs+ngNgZHt2lwjy8i4d
k7EDPNgvgfDeAAEE0FnAwLLfGgSTehSTYg5vfKNnEtyMWEdaFVgKbxofGObXzIsSENlvQ+1gyaav
sQzCMrJkHUV9Q8/dTpBxJqR5Kgo0iyx7TXN7Azbae8+1rnKkPNHbKTzg652YPZrJs1/OIMn7mVTx
lJ6xHwIfDvjFb43PdaAZ9iM/cTxy2n6K95Lf2VKfg8vY+PpA+vd3+k5vNonQj2JhSvKvrGBp0kI+
wvGKDqGQPDGM92KmQQYVpAVcIpw/tPw8wx8KMuln9/IHfLnxblwTW9qfHQAZverlbyDc8O/48W69
fSXBAgnZrbdM3VftbCIA+n5aWTWocH36a7XGTp6nrclsf0UvkL9M9eSHZn6X6vFz+2UtKbN/trmw
azCFXrBEsEeup6mE4LegC8IhDXXaB02TDsSqqy3uqtuCNR/QiOVh+gCsU5xwrUHyPsWK3AiOtSSP
RdVTwqPd9xy1Zy7Vr+3gMNglIP4g3GO4iJ6xOn7oYcNk+ToKm6JUbYOpy2zdmhWk6s7j306duHt5
21DwhVxTg65Hs+FC2ON3of0SxmOPHlUElh6vw2PJzHMq8SpdBZisJUx3DOV4FagX2CohRIGq7M4z
ugOl+GTOIvvv4SQSNft58x1Nn68UWX/Tf2AOVslqE3Y0/mqU2FuS/Yj1O0FqWdztuQCXNACrY1Bm
ff7q+F5FzVdD6t49xAVVlJAAKx+Ig13MZiHP5RJdbq3eDrb6HvpX5XEDF7a3QVXBMdU4dJDN28Yd
v1ZcaRzlLCR5OnGxkEx4xC539nvMM3/zbRrcoR/ajYoCRj3OG0zjvBnHs3CkN5hpCm3CblwimM6t
dAgsxSSrgGAYch2ZlGQwwFEeWaZz5WTCUbDLNHsiYJSJP49lnDUK9TPQFy2lQz6LlJFUEv6Oo8Gl
D/oJIYSBk9CeibWqt9vFKnagbbiJYfsVK5Udc1KeGE+vq6IVLupVf4LfsEgEJ7jQz2LE5xBx4GDK
RJ6sUaDPUteFpYEHF76rW1PhHx6/8DcEOke6/6W6BY4ef9oEkAgxkI8rCIlcNZn6K+2lgL0T8uxU
L/Yt7HV2HdJTm0tV+YxO2kvyfEI1/PF/dYCzYaDrt2Vr5cXlcrPHcoQjEudgVapNn7WZ6v+6iO19
N/fgaQXMKu4gGUXCM7m+KEEo9aX5Invb+bRknBhpf5UCH7O7naf6Q409GRrOjMK5RQVGwatcax1M
c4zS7b6z48SI7TdK75xn//AQPkiaW2xZfKFCuBOBOgZdDlPiCH0fxjDf7Oym2oDWJqEws4Xf6MtH
+b4nt9vCOMElg3TfqC3jYsmmBioiB5U651AcIlAGg3N9gaF6MdBcAEfF0d5cH7tI1nyz+UMH9XzA
IPaDG0d23HC5XbLKjl7hR1dtb+TaWOy9RoILqwzpLIcW4QqZmzzmuQ4DHhGWkQvJx8Jgh8sqn37/
0u5Q9JZO3mNBJYAt8AyyAljYMlLvgRtnOR9sMolmTf/Zy6FGfk8xGN3RxgFHQQ6nZsER2JbHHxlX
uQHHyGbAUvePQE9Me4Qo40CYL2AdTDPh7KwPAllYoBi5ya5a8Ug8jgoyJ6SzK8GXwSWmLZJzqroD
Tqnfpv3ZUIhl1sVPQSgn4eIf7rkpfqnB0VwJzAlSmAjOUVYbnME/WKqGCWjIaKMemDC3mQ8o72ds
QsLHAW+Accay1dtV+RRjcQ7v4UAsG/nlG1wd2f3mkyWIWqatMgq14m2m3foRn9d7q57K/d+HHa0j
yaACX4Kpil48BST213+5Cj5ymFjwoNmGQCmzh3zmyPZj0Gd9OcBqlYApJtmUFx/1Ic/uIrn4ripu
7EsC3GlrIaH3l0yPT+T5lyUaCqE6jQR0z5LlK/hBsUKEKD1vSDl/sr5VFDaHHyp019yDHWlUzUwE
CBrkmcjHxG/8eBSShfqaDbN6U35/AUnbiPelClFG2wU/afZPLsU0A27nblUVtVNZjcNgiR83d4iy
kIIQ7tenv/KJK0hYlXWV03y1JHSAuneFnLXrl8ecD3FiepWxpyzu+4zc1rRVBleRTJXMufgODmkv
tuahOmqf+3PFO2Z4SWCFKXpxzd+gf0HfNVLIfC6Fd3nZsjW5o9IQS8YEYEVbH4GqJ/kmslCHE9RA
H9jiBs0931OKHa0SbkVlFk7IhLfIvATOgRSEQAVXFe3e0jZ1UtjrKUN2qG18nTflsfJFiOguSjsw
7Ym2MNTWRot1JW3bGKXzRj0Wdr/XUbIpydVUs3OZODUhBYWp6x4btkLQbfbxBWTXcouW2dX/Jpgh
kOJXWtG7dNVnAIP0shH64ReeVfhAkDe90ROD479JQMpszx90aJvbq26PU+RMCYV1uxlKmoUwBzI5
DXN0pbFs2HMzIvAtdKWR06iHEoq6MQTVBQSkDmjzA3A3nK/eZoG7CpG4lnrbW8146YW62AOlrRIi
SNaSH14aIfpczhw+NiXyt63pjiJiop5/3W8GsVCNT9XdbsNA3JWyMZV6dZXljTUCzqh+snS8B33u
8N1mrb0DFbA/tSmGiTBGyw2NjpHFpFZiHBWH+mb4uSWmaaUYkun7/NkjZXvtHf4Ov9NcEFJ6xv4s
HpLM1JzZoQgSSPOxZbrZlJRJn26wdf+AeRkBRq7gbBjawhHVIZK3XokFgUBd3gHrgMg3BE9B/ERw
PWtABHtoTxp5A9Ahz0UyqDJgUH5QYbKyYY3M0S25MB1sidjEiewgS6CoAzLvutKvWaRjieKukbTy
hVGtMU44pJnZMWQABPWe2amrO5/Ib0gKxyLVLK5l5Ln4Ck82Jt3lAw943U1/d8vUq+1B74G+IE9h
MWyQ6xbb3syOyMo+1c1Kl55VUP750CemGwuPGw9RkyKX/Ic7PeNzeInkOFOkdphxK6mSHVN1OCay
vmbAoA7TolI7qK83I0QfbdgjOJ+ApZfHD9Skgud9HALmaAUPFE3i1V38HBC+4h9tASnCO36PZzdu
yB9b8h3oiG7hMMS21ON9XnRr/tGGwqYTkngVdJqB30Jl0hJuHzcV4CbRyQW1auLAIm8l8+rvaGkc
x2ziZecGZovE0wCJl7WQIF1kJZF5UibrGau2xmOsL7L0JbGdSEQq3hH9x2Zb+rHqpItsatD2YaUn
lhy/JO5iCRRGgidittlvJM0/3Mt18Ds9NWPg0zDH8p6TcLJZAwUYdqOY5GFH0o5LwaRMAoycdq+o
FU0ll6BQV7tZmw3HCpjflQ8wuM7AOgyIFMovwkCWqz2SxFfyqfDwazipSzO4QvEnRkfkg1XNd3Fy
FAUThY1MKNfq+XILD0IOjVMY6l7xdXS1d8YygpP9pO7pnk0US/IHFCCMGB7BuCxlIASRVsnWBtzE
F2PhPFog1fKSxM0XwUINXzvrJ7VoFJ87rc1C8hq+wkZaZgzqN6NAl3mh2WR0FiOahkPzwHO1c23t
IH4zlnpU1xzHH1O+bVERzcimwiki4nfs6ydw1NBw9Bw4MKuCUHDtt/cotRdFbTcZz1zk/iqRVzBW
fLubSWmpX7EcBAnoI51i29jRN220o4NYYyMffp/UhDW9Nv4rD2GQmecCBirJinEB8q3uKUCLvJPV
OYQClYw2rawJlu+jkMCEcASXN4L1uoi60+zvQDSvDw6Znu1jYjpkSp6er1CsC1FoqI2TgRXQgHqz
TjvqpSboby4Z8uMj7MkTh8Sm2gqvZHxf6P+8HPlxzR0nm26BYHovOWlqjgICgrb0m+1JQ0+tc+8o
tGfjrmC03dKyUzSYZbBn1TciQI3miw7UrgjYWzEDz5wANcfrdYQinJhBZwouxl+XGW3F1+sJqTeE
1FIeb5tFBpAsWQCl0GI8dEypa7Xe9EzMbSNiqAsaYe2KP6oATZRemyCB6qY2eHKR3i+TXhCHrGsg
tuJkgxuSzBiobwwUF2FkuUuNqcdx6Q5oYeCUGk0wDGMAjNCLf7R3PAcCiGoq6UDE8J87iJE+8ND1
iyuD3u0OlsWDhOVaUV0VUAbfTFGDFEAqRB9F32CDf/ti00+3cw3dVjLQ+JoXG4WlU2O3tmXpZ8jn
qVQM3jAijPgekurpVyRWvCR8zDl31q1H6/kcyZPYQ+pLu4CFCgMHmfkz9qpXurgdBSVzHeJunIYJ
Icix77e7F/ztJSlpUKJZU+xqtyMV3JiUK5QPhJdc33SVWQW/zx291zuglPPQ5qSHIP7lAqyeo09S
WaK+7Tl5Q8mhu9QXCwddF001XFCZ0TAuex8N3NKvw+PBBGlb26ZqK2ye0C5TKJsUQeb2o6sKESCl
u7093bbwdSBReRv6pO1158noKOGImf3npCVOoTbjD98XDYbgkiCy8q0zxBmM2pFkOY5wWra4Z77C
1bwCbKKYuTt2UZl1yRpWGeLe0yY7W5EA+HPVdFejRBaRWnumxuveJtwLp5WURmTh0UULlPuVwErO
61X3/amCRzoJ57AhsvlgKy0IRWDl4nnWHLcGLAFQw61YaGJQau3fZlfqB2IXgPbCgMLbAYqWExTo
36HvHY13pkb4Xiea3vAkYI6a+uyJHHci8LwLovDF3QNSMFfkZbevBi7PP3hMeoLBZo37IFEE/pgy
Ek5TUL4a8ImJV4zyPy3RAHUT4vDzuNZ2TFHJiQ9rlmQrgKO2N+FG7q1xKDsNKyFSAZ87/U4aNdAZ
MJTX9HjUljwK6GIo14VWRB+amgEsepfpvJXW71kOEjIOANvX0VQjD/dKAt1BN5gpttylQrijnGoA
V8HsW6MiAKolPXnwtv56XEV31TxXpZ8Bp+7uQThFms7aeT1kwOJVji2VBfyZIsxPVaTDzeyx0Srd
XQLYosT/nlA+6r7r+c/qRFwqXE00nf/lDSDavrT9hTEBAKINDO3J2AFzzt2qjIWROVlMXuw+JpGw
Qfg2Y6Xm4d1D1AxVL+WM8gzCIMRONNvYMu4TppHD5Tz6XeQDi5v8TN7mmJylM0IKhHxhaWJ1kRCg
THf5X/s5LARrxUJ8KUR5oCkaAwG19A+KAF2curDvJ6Rd51Kv3gcTSTnwytuoZdectq1X1unzHVuk
+EJmam6bv1Yzy/M7nMMzAH14PrOefQRYAiM1TFvbONP1Bn4ag02+HO8vYS8QstD2498eJseSpuSR
klZ9jhWc+CsugLrdEh0f5it+G+eVgUZ6Elm/JvYkja9iQo6SjxjGAqxWXnEdangMOmSYlzvgnK8u
Ulii1GkwttRF9djWM1QQlqyTJgE754AttQY8oRU5usQJ2mRLyhCviDS7LXGC2IBNdAU3v36TFNZD
npkgI70hQYKo1rACNcsqqMptFUFu8Tvfq4/yLHj0yGAxgbHpVDL+2RyLWYlh1TpG0CGmGo3aB4zK
A1laonQkeJRKVAkmzbYL+6PxAUKb2FH3UPTW4ZyMVTO8qY03KNbxgVV6P0tnThAshQTepNEXsYcU
zFm8rt7LvFygjRfVoYs/m7N+B3oCFJbkjKCu/nHwHT45IX/E9uYFPWHqu85Q3N/NSqzk0LTHGpSC
/RdDNZEknShVNt4Ouv/bY9UHwWj4AIkv/JPk6qTpkLvehkc47EulrYA2qlH6OXCXRnX6RouV16I/
0cOtz3Rk82I2FIZTtOagQ4sgb5npqkPF1C1Xbrn9lFkbmJyqQj1TqnXs0ElL62hqsmqmeROV5owK
WBOkLwxKBVdyb/eEi1yDyHdsNMzCeRtFby1GG/VoV832d704KnhKaLzK0eeT/ztbkLIcJVZwqrFy
9mSLQjYDwG+M5q3EYF4qe/6DjfDGtiP/2Jx8//yWKMqA2WKsx8jeF2C/xPRNp3op7pOrzQqxhFhb
VG3qIpoFZi5fdYam4cjE3DvkvN7ANw2Tcqyx5URvRb162FmguoBzqIDiSrX7jYvx53ygbyvbJ7ol
qVz3GFudDmhxIr3JaLgPRlcbs+0S+l2f1qUFHpNBQQ9IPcTwaapV4UsvMguVRHRTNCcvBLPJ2jw/
yNR/Sf8ilOUcxyty+JR1EKdyypumcbOrqFceEkMIx9n6ilUrtKrr5l5rEFN797yEGHN3Oljt4/qR
8+yFBPsm6oQ5uaaDgAC22orFYOxIqINjwfZy+dqzKsfj711yJBsYSybKjldZjZ7XeYW3zd/tRmqk
9A8kv1swVsTdmGCepjfNuuAqLIYERvzHiMeMi1HPUrf86wREroYrFzmQHhonrNYKe9G3wogUWzsk
omJyms5ujhYI0tdrPSZvktRJQOvywqW8OimUe5Y7S6Jv50v9tKbHJql1ePyYx27BKu8TRv0ZJtzP
NaazP0nC4C3l0MzdBCg77Vdc5f3tMO2VPmomA+I8N9PQzK0fRe4NFg41toxdHTSJNVc3Wgd/QEgw
CU/zvs1L2V8JLxoJag2DKYFP6aKAhlbW1UORdsVTXcqm/yi47Nr1YBlgSYbvEZ/mlochD85iv/YN
2NiAFZ+qy0L48hWktwGFzTwPc8StsoSPVwXPihUj8a/7yaheDCcj2uw5Tdf1cTRWknNLQInLwmts
tkOSnMdk4sc4YNGXCypDTY+XKU/P1w1B/13fqik2m+LKP/Rij3lLOlomEA+BJK2mXpwimrRypfOt
Hm6aD/gEV3+IDdX9OZQPbJ9giEbANYTmOUjfw+c//2xjsqGVdcCGfYZw2eEXjmOEfbaiW7aAXJuJ
HYHCw1rHSBeli1UYbtJ4u0hestMlj55yDkP+apPsYq8ZD3dgnrckQbWowlVzUS9Y7RdOMFYP/Jsk
GBnfvIzUJHSuFSdU52VzDhXxxA1C6F7qKKnRn5AnfZjw7Rr7h+TCjP3ZNsxkmXNe2SHYlw9UQCns
asSwXF3oN9l5+MG5oicreHURr5SH1cwXEEC+sac8UQEYC6OQ66M2SLNtGP+JCWKWqeVAiVCVMciW
j19CLkIYB04wdaaFzsjYFttq4qitcc30iDjjpGQwMKgOpeK3EkXgdIJ+OinYzUoBW3P/Cdatw+0L
R+4al6CDelrmk/w4rVyZe18BqC85Z+zhb942GN8JU+e2rnL2WNNrYaFFzLVcpmQjNK1Ynnto/mTm
c/4YZbJpGw5plJiQtkyus4qlaATqK3M58/DfvgX+3fsQJ1HEacHzQVXfCbsb4mmzbnuudWk1gehF
ebPQB+/MYsfqJztpmSCA7/vXgkOLq00FbhXDw1kUnAo2DfKXHGAciYBP2xriXyVZWTc+m9tLrXUI
+Agezj61EE7KDk5AkhQ45ExExv262kuKuDAp4aU3prqa9kpDd2EJf6saFBhcz1UqnRytdcg6mTVU
IkK54qQhS6SVuPbwX1WPM076Zjd2zXJhzycZK63T8HO4ZwQRLqyUQK7taPFlwr5gaUqzOalpmvkN
mNTgcOSgzqPcr45zdKFTfQw5wZgLre7QJPyp6X638Ii9SDruHHnnLGebj4AdpIwdQnCGVc2P6d/e
pNDawSypwHVbs+UsTk1C3zPrrX2XRBHR5A3kyjgq4Xx98+dv+TgBiGOmb8ZDzvul6CoqLaSlcJtR
P022lfugEu4ehTBPoDK3cZcnjjdVMgt7BD9heQ0oiIOA7/zHdzQIdpsxX4yrvZwTjS4NTv5SH8Tl
1+7t/IXIggJ+yJGoGN8eG3GaHI1mFWGBvxn+BXCiHN7pssSvSB65q/o9VhEFESH/eJF9QnUwOPLJ
NERsBnfv8/SqFjkpfiNwbs3eXWmSSmTLPU6QQtWyV5ROMNAbxvJmVUx7fDe1S3N6Y131bxo633aa
+Leu9eitP1TMGDqo5WQnddHwEHtLtXHiR9nKoewHo9qcjJw/tMLSpKFNvEzI8NO5OM4Vj8ylNJxh
9+Wx7WpiLPD2EG1wXOaFp///jO0JsSBCxbkMdftem491XkyslgFi1Y5BZYQ+wR8+w3a4QQk0sV05
Yofy0uTRWJjUkdvTJ+X6urmn73ZoMVmfsnS6HVmUefGe+RjUI8BgX5AwfswQ+1uJ09T5zEKvYwWR
JX2Hh1sCkLTMATt38Ri1yahhZap+FV0Fn9sxT4Fwf3/4vY9I62N1ztOQxtl2xRybkY3t/ltgpgfw
C+bVZ8l0g4P+TY4IDBhrpLnUEvLGC2A9TNgtgOoaLvVqn3oeFDvCzQfAXhJihgb2x9IUr1OP24UC
g7f3SHZr/fKoyMJQU3iZ9k+8PpqVCrfjPBLtqyUs6AnFGwofjOqJhGsXapQadYJGgwBHN2p7lIKZ
+h+qfOooLEabEM37Cp3aH04LllLVFe+sFkzq0T4Pn0OfRyyIcOKYQnXCc/lDI3Q7eTGZJAnYU/T6
/ckKN7JwtF7C400PJpLne5ll5gd+nRMo7pkHptnj9NDRdFsFIUNj2F9L5KdtcYo0Rkf2TFx5xyJG
N/wMdTwsRUKRtu38F8c9pWQZycg9BW0k65ldy7LefVFv09swDEnOor1m/08RxIaFA/JpaYL/K6uB
exs3dv2tRT8DO8vE3d4z3Ax68geZqwilTbNtMnTC/i87SmEASOGZ2QGP2snT6FtyYEEwRmC8NtiG
OwBj+s1BmtRhj8CHReDHynEvEqN8HWxBp3LjOFHkFTTAq45ltUyn9T7fAcdpNwQyiCwGvbT0KVOI
qnzuTMJeki3GU18PvkwWkfUGXXE3GcrFCbZnctZOdVhA/d1TBnbVPnmayKZ5ivmQ0JvO6M0MGXuN
5EWT+M3KD4GC7BV51N8DMxa5Dti7VP32ddF6gMfPZDqNV1wOcCe8BIhDKEPHyQ+NtoYT5Q9XhfvE
UmA62tR56rShFQS6Sf+dD9TX0JFocxSDTpOT5DU3FmMb/Kgib5HcFmYgEEr95XR2dBYJ6+XFY+OF
KwGW9ma4IXY5cBv3ywpWANMWYR3doSeJ+U6bN5b1rdXmCQ6xqnTRgwfwh20Ibx5SmFaM1pNFQl6O
6TFtq4dI3HODkhsxP3jtRvXK28941NT11lXo6eU4kLZPzowyk0xkU+S47tcjndi6bz6k+Y3xdPCY
s3zaYrQZmJzk/mF1ogL+Ato20bTwlRV6i4MVyW2X4qkuG9mZdUA2hf1HItp8E6BKTWHvpIxgpCcK
+OLAnGhdIILnCxy5Ma1RE/lOxr5zfvLy7ChZAdY1mDvojDuRThvhJcH+Ldgdt3QvvJJdaAeoMrEx
Yd68Uh1Bq9ISlHU/Pl/Sgnn4EsI/qAJi2pW1cAN6qqHSfXCtxoyVAqw1twFplJkYqoJK8zUgIrr3
pe4UZqCRlp11MZvTtz1Q+k1QGlRF8Kk8m3tvo0e10uxGU2XpM8dsQICRHZ5qM+8tOsJbvc+sw9VO
NOYqEB5tFKyFalEkv0K7Lv0rh/N2q92xHeQHGcqU4F1bEB8tSqd4JP1rG40LjdnAnhhIblSGlsXJ
GpAlX5vKoXzpNF+d9818VgUKx79Y3WgpByrDzFlZ9ykNBr9rfeKxPpmqFOKfORAc0e/b3YEDX1Ld
+0PyY3tvLF9YpFswk0xQzX11eTqdv8aGN/ao+YgEYxiPhbtUic9oNN7fl0lAAL9LCwzaLI15OQvR
Szmxi1gGUPoy5cr3cYoT3yj5FK7tIw7+PQed67wwIQUlH+bZnemhtVtg4HN4HvoCuKtc4P6+hbPC
N7W7Ix3pYTqxCuMvvBeR1Tbx/874MPfxvZSNja+dIDc0rgjo9XSIn9WbiUpqsGvsMSALRUOEfMlH
s0rfzqMbzpEZRMxUURV2NiqDO6voElX/WvBRRlny3VEY7yAF76ps8lYLsXuESn680+Z26skRGCCi
vGxzW4dXIAQTfNFBmuTav1BSrOd11gzJNbFNhkro93slkRec+5YdGJT7QzAAwHaToN8VCw0PLkK1
JlmsvM7w3Pizt1bbJ9KUprAtWMSHXXR0qJgqb02ZalU+Hy3KUXFwPj8yes6DhQjYUMml3Ffa+PZi
EDyOpMMfVmZeGI49tkqbB0arhTifcAUELPt4IP/pTuJjw1vDumTuRmreLC3ETVXAPY5ExfafBOxl
3bGQXiWHEoQ4ZVTM8azNNCKcx4Idkwr4z3qhz2l0yAqWvGgUleAbgFTKJT68ek5wTmWd3zZjikus
K7mPA+mcfuWei262vIzyxfNjRsKYjMTw6Gi9NG5veXMj7upwoRAUTglwEz6/QZ1hovy85OxTRU2B
gkkCI65BQPl/u6inLRpeVgo9ctzkdTnhDuU=
`pragma protect end_protected
