// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:46 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
jvkl0fkkNbNPKTpAJ9WvbK2dDcoudQ0PI1LX/4n3I6QiahlijFaGEa6k4kMgHmjL
KqbtmwGpl5qQzbA9hdShh24QksyWyrEDtyrCphX+HlXbKgb7Ie6ot+7aurmBY6ms
YH6RQ9CoOR+LLk2Tg1hByFnVfmIY58laLOQS/glGhns=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 50720)
tToRXrFkOFpf5n04HuWOaSoLZ/1IwShDbOOKF8aHWb/3n2SNqMGvzZ7D2VRJXcxq
xbDQphKCr0vcUWvE4FU1c9EACMflpDiylundR/GOvjyTlknR8WWh7xdaWPLM2CrF
/QmOR7c/k3wi6WGKwsRqfgaR+oBNPxRyagBgMTec28IyMZWKoz9rDZ025cDJKgWK
srB2ZDDUzVhwziTN4GYhANXVGyk2WpRFKaGKrYZntN6/c3ZPE+bmxZoSTazsVnl4
MaUubLXCXRe/y8xnMZB59GfE1eQJOLhYkBsqkookfYSP8H95bJScI+vzVWMzfIJu
JQDX6SCu3bVysJcHpptcn86yyOChK5E9sIIlh31/gKzjNpNzMPP6jYc1JPsi5Nz7
qs6swFdA1UmiVLLLbkul02e6FUh2LugI6iiNPyXk4z5E6JN7e71J5X4OqyIRzJT+
xR/1lUFmzb47H77u5cQLqhNdCcZVMRv3SVXESDkv23WZsYnAduHIiUaJkR/T46yM
OLAjV5hOCmnvBAC1Whje0lq31LMIHsqYz9beNEQQ1w8FvaoFBWwek+ujv0C8crMy
fbu/1SunOqLdyN9Ksx6d/cDXlCbrmhia7L6sujcpzCxHlMieZpPCei8jZYwXQmFC
+UTOP+gXor/8dpm5+njZQt/gRC7PhHc1iDImJ+HN2uWoHVkoyC4NKuYCNWZ7bHLi
WLbRKG/lffBFgVX7XdRT1BnuZt8v5SqfNlsmNRK++LuaO1/Pg/dDbcyip3dY5lI1
0jJpchLAeyr3yXcv1uUc2WJ6wBu2H7VM5voYLzrHdYsriKYFgD0jnFNX1kddPY2y
BrlL9JmZdsxxFNTBspmQEWaVl7Agxeocep9KGCscEwgqOZsCK73auEk3pqTcb/8a
47DDPZ6LTswLHwqwIY0FvSCQUwVk9SvVSTdYARQubNcxKd5jMEmzJBTBMULqmgQu
U+BYpCIGaCm71JSjTDzf8P00cGRJFfIDkuiKPPxEOhgIVQFaGZdfsEnbFAamNe/T
FRu8aTa0iQzgAZVr9kEjjqQp9LyKG5nl884X/lB2xcn+osaTHUyeQocXZj9OdimN
setfpgEX/qpApIVUzIuyfG5acJVX5dAh007jw9wCbwG8JmCp7f5JTIo2lc9m8SBH
oMRfd5NKDXa4A3lp0D6Wh90DnY20I89I+UccCy5SWSFlttTT6a2EGTod9APnbjRW
j2npW2ydvccMAFgHC1HS6rfsp7IIyXbtzsir5JfF8L7jRovuzO2jm3zSDquwrTtx
EV70Z5x5xCcrhpzMwmOez4r9IwgiH4Ry645roomcnA17pdAgwIZLcNG4YJHOQu9e
f5QH4EVTt+fojbul8aBHIxcYMDc6QiatmkT6155rf5i2kj8UDyVY40mucErfaOqG
HxoLfcJ0cT2RUceNNskI4674cSXvjCCSpBYwa7cKXEiRLeBvk8tSIuO7k5oxf8P4
l6KFLTGfuFvvpDtFcjpt+bWkbZG9yJ4BWh8/GQKK30Lr3GHcP3WK1BBD2lc+yL81
kpyI3lp8UsRTMbjkb4PhYyd4xmZ8TIJGMOmIiWFPP0acbWXVYzAIkFBuHT9VN7Js
rnGovF4UBvNy2QQpLtHYlRmufHn9y9fqfsiG4lr5Y5C/VmR9n4jvX8QGzku1B3UD
LHjOCWxUB+mifbumP+F+wLXqAlCI2aRHu6I6A2/sjejMenxBF0qzMDHtaotK8Hi3
Eijy0yg59NJVXA4/ohNVABL0ifMizaF6HXADmqwv5wvFtynte1dNol/f8EFp1APz
qHSrJFNWiPDfaTrmBfKYzeACgoXF75/KvJOnr2kjBkfy1WPBDwo34XrtO6iNNQLK
cHwVPYjOCoq7j8qOMKhitxGX2PzvzcsukLDMMnHMiwVkRaGke546R9y1IuI6cFjX
9FuXCjIisCoFyunviaqtfh+l1ebpAEneR8uKhuD0KTktJ+Q0y5f3iIeyrbDfkJsa
q7mtm3emkQPk2swSfrK3ZgFdSt/dMV+jUXQ7yaWGdzKkCocdyFmnvS2ZMFZVvcLc
tYdUYSBpUsZI1FI3ZoFH1dDW2FSE/GnNVg9aVAA17QWw+ZwFlAsRQF4LVqqvIRai
UzWa7ce6F07bypqap+xAM178M5C6I3O6X8lpDxcwyf3fYu27VQyNdSAGo31DfJ2H
LuV48NSX0neyYRghZyRsddYds5ORxWVP2XL+ZfwJ3n0Vdm18iPEs7XZWswNtuue9
PYiRwtdknxykFuELkntFzqt/76/bsnOO+uhgTqIruibUwz6pV8lnvBb9PpGk0MEo
6AdRunatnIQHF3Nt3d5rqNoYLrjl2l35KziG+INhc5XUAU5N7eAy4nOtaOkLj2CW
e1FLpapmSS/lhjWqN0DBRwvy1zQR1hZeNEe3eov6KLPI/pAnTytAU0t7EWlilDpK
ZAfVJLrrAanO2BTXotfOa1uUUmHFAKt/BFbYBnhU6HtJYC3mV86dxEqxcv6Y4rRL
H77wQzQgT58QySFnvJC1nJc8wcA87dGYtOuWl6EdbcGPPdoZ9uft2XJgtkAV/BPU
dB4D8MkWMB558DuRZd9b8tBp2kovpbgrsW3UWgAJ5no8bkp0yitgWbXnsIBkSS0q
n3EaikzPoXL99DA7uErpXKDM05j+GpQwjpdYs7Lq+IvPvhT74ZSeqq8fpZTWmF1y
svxDhq+iKEyIsxyXDWQn3JC8qBNbikLoY3z/YguPITANA4MN91NEV5ucqD1vTC/6
s2NX4fFqhwdZUjxk1s2/c5ybYn4HLyH/bwICaZrkeWJIQdmGAHvYCW/Fx+PSH82L
/uKEDvicDVJiVXiJFeV6eb2LHazkvLVk19ItWNe+t4qaZQHwgHq7TR2RCo28FPwl
Oax91aQ9PQP9cydFl4BpEYZA41nPxM8f8XFQnokxCDMsFQPN+bXotXI+q9T9uoDh
xU+Gw/sN+DVGhWPK4IXRsBOeY4QrdEB8eKFpW6YkgV8w+U2+h7igGxilseFziak8
poD5D5Bjgg2kOQ26xca2glzqIqBvabLroMhDo6gbDGz1kQ4qwBngKPb1jJMoD2E2
xDP9WZF2FTwXwbXlxDv/41XAdJuc2XS/WV1FpAYWazkGfKheBLPX8/Px7OxukYCB
za5ep2zoVE9i4MCX4z2YI5BmVUgmNeAg86Iwvcpuy18qC539Q7Ez7A5vBPGACkLA
CiHb8VZln/AIAUxXV2o9AvIzUjyOhZCX2VwVNmscpzhZ1xemCzJKj57aeQaJDZ+m
5cX1MGsm5/NmFEsKy6hwulNarDZfaItWO3XJW1GnK+TRC8wmoO2jqfPgSdQ3/hrf
xIezaubyk7WMWxaN3T47I5zs+GRmnNqhY9lvP78o5JdYoSQiCsk1GviG/lKiANgM
CcPbRLT+izstN9xxsIjip2F24Zvdkj+TI0VTaxMG7ExVNoyEYOmoOg/1QvecNnSJ
Kg10Lt62o52TgJOHc8+vUqQAdyoZ2Tz4/P0GJsDzq+Oe/YqYZJMv6bzi2inXuqU8
aUFkykaI/adFDVNXP3FKtFWpmR2+zx3GStnqeTJGYw56ey+tHy2FkPU9D5f2tWHA
D1UKiSpFwKA7OLQrQ8wGPxbi1FErzWHnjZtAtj3EcFm6D0rxo3OSa/OUroIWEV5a
8dYBxDVdspdgllvN+FfP5pAHIXOXgPL2B9F6m5AocoIN0v8+9GQ3hwsvmUZ+cPvf
aUbfvk38nmDVB3wptY7jLDKLn5BoPAk495rihWH1SNuV8bKeLVMi391v6FVtp4bf
0Zdh98zlmBcqXElwC+6nc7ndi6ATtw0PbSbsWxM7Be+5jcQXwK5h+x+zozK9+83y
WZaQlL/pbB2ChRZPZDOW7yjJr2G1K4Hj9KMPP6BLVyysmOaT1SekglTTN4e1Zdq2
eOdUg2Cb85NTmn+McitJGqH7OIj6hVXWTNF8TuX7ZeET3S8NmA30tQQ1xoHq8wob
DYsRlRVunBqljlBInbgfXIa6qSX0pK94MJscf6oANDcU2yVHYvuagyY7l0I0CEB4
Vw9PuKVO0kYcY7kpESYEvScQRMF42Uj/inRDy/KDffV9u5EdbIV8vE7d+DAD3Kv9
7hkebvj5QAkJtIuV37hoY82xo+j9JP695o8Z/PlcGj+2vHxVnq1Ad3JGFQxNE1Hx
7QbjnDhKJQEp+2U1v5yEu6t4OWLHVekdhdVEFKz7e3uL8Spay4PBTaPSy1CorGU/
R9C75EKn/fegGGshX6LOapRYZ/WOqJFj1RWRgxCCN2+qXIZTi3k/UHHWVmfvbd1W
qwp3nrEGmSebxyupnvVlnenGinIHElgxCm06IZDDpBiajp0eelhThOMeWIXY5oXv
N87GTG+5/qcr7aEnYfB0J/qp4/wvtvW1+fdmziXdQeWiyzmPs/fEoYdTUX4h5125
2TPajZ7F9+D3Q7IlSh+X350ypBEXyGAFdSNXBYbnjnnK+LtOblbJEq/re7rEfIK5
Rkdd+K/aGmI5v7FsvJcOi5PvdYa8mGOmj8HzS5Qvefe1wsVUnyrgVmbCmffu0FN5
Uyc620vNrM9rV+/vIgnkzHjArYO6s1XgzoyGQNiZCzou9iMZdTIXSdoBAb9iiN8n
Kzts+hUH0XdSpwg/RbsBTSmxxbFMVfwYGuzYxhy5rrrgb3s1MOZMGjSWBRwCctLw
jCdJGhxjaltXMD8MI2OH5s2X3wjORVj+0OR7cU15MOZ01xvJcjXWllD9YEi9L3L6
AWLjNsqKmymmexRIeb/ZQDwLk5D6cnleZfxT2bXW7JkAm2Kb037zTpt3Yikxo07n
xQeelcnQsdj6Bhwvjkh2VTm6i5MNJbqWUYr77MyLE4CPiyntDeE0knE7nhEkrpMU
VCU46dtEuT1F00FZloqWs65eJ5JpzekcAtxPAkJoO4FODufKVcBetO4d8YOjOUBd
nsC5BIro2AWC37RNpDhHg/k9IGr4gqvsbhSDOcwghKyWFaHwCYgLlzB+skXPh1hE
Cxf80npYiB5GL7mI/YMlW58HlzbSkKI3YkAFvTNyL4nTNHevPE4rGneeDQ1JOroL
g2ReBAIa/+t7k4h5i4PLt5I+8BwL6gJNCOtyB3S9DmDNtm62XLe82mXaVlNQLofK
CxfQqsVioJ9V7k0RoweqCyCMvt0gYqB4fg6BZEOwEX/NlhbVth55qU7OwyJljvNI
6sCmaACrW/O0lu+ySdcfFMS292GEkdH5fMBBn4VvF9VlPSYfa35OYr9wsp27OrSd
TFWrinYE42je4aD23tJSVErThzuJzsM51Z22Dm74MSG/240duPZ69qVjpKXdUPyK
cDCBRa5KJxhvFWo+hzrMMb0Uqw7T5Sz+OstGFUUK4q8iFuW88AF/v8wnvOMRbRvZ
OmdQHw0RRs/LtundUJ5MLm3zldJ5NX9iQ0XLePFIzaFqsilJ00i/QRXcJEsiD9Ze
Cv5Gwye/ChXsv49CEBMNsGO6ItQ3nnmHhy51uUVjqoyLZ8CH9yABnjMIfmbwFaLM
376W67O2wUHrOPd9ml8tYODA9gy/DhZDcAMVqE8HxTKeVJnZAxOyZ75weLEJfRnS
eloXKLRZnOZZ7G38X5OKqpRH7D8AfRRdy5aLOWTq6+R2kdetpZR045ywxi+Q6EGm
zC+yzvyewpWFXTSTkNnmz9UuzjLuwUbekhNv147jbKKeZ5T5nQ8xzbk0PMgLavFQ
xt6k4XE77nl35SHVDzu/5QLl3swBKhbztFUZ+wB1zFLkQPGx+MQFX4syThBksO04
xmb02a4RFftBlzJ/ZrvLiqK2VRRNebUFql1/uUY4oMbYjJSdYkbHLdOpWdiCAqYi
q7aqnRWD0dAfrJ7HYhk7HjEcQK8qKn5WnCuitr1o1BUcfVfR5g5C7Pbn3Ha5iU41
DWd2CoHJN/lYKntf1Gug03R5fEBeIMj2QeX9itthW3S+JBYP7wocqKgGlXiIHiG+
ff/tyrsCS5BnYuHdgpDpYyj0KmEc1O8J9GW9QWioQYJ+aVwCEJkFmxjpEdrKcvrh
L9tNfHLY87xY5vN7Q/v3OqSXYcewbaF/SKn3oNAvreDAx9nOG5dMo4BHlC0kNSFl
u0UpaNDw53hSNqthWv1vKuQaHk10a5vGt0NHqZHhFZ/xffAzGIBTIvM/DBfWPdRc
NAdYaYdVSb6ElAM0P21Ll2p8OIop0q12mjknMvbrg2qyNTBMG8gpe+4yqEVwOCNz
dFyJ52jK7o/LrGg1K7mry6UD90g/2mxE4VvLtofneHfKBpFnJOS5l5GcrnNs8Ki4
a2wo2UT4OdjYFZS9iJnWa4kpSEMfHEqJHUJJerNo+qmgf0aCyYkuXv5dEsi+ltXC
vhkVji6dW01mskb+sHhPx40G4it2J7zaqaOfmHLw9oP65NuEPXZIU2jT7atHWPAI
SY0+h5WvG2qClXv1JrDw4o47F45G7NqPCOlSLH6p1Sfx9y1LegmvExWWR6kbyBUg
H8OCbk1K3bYKQ8d1ZisbYPHkzJl1RDNpn+B9ZBc+QDTHEgwznWbBUg542NI/YByA
/Tj/qABxNjV+eazNKx8xt8bkk3FSDrP0DwX3+/QUlyRn/xbhXrp/WJbW9Kvy6FJw
ofis+EnShUBIcFoL8b4ksKqoE8zE10zZ1uT+uEe6tlpd2coMTR9woO889+ri3nug
5Fiw9T6zeLa2YrtOxaZHuafIedMzjNWpOBPSwk0WTThNyVVpgnldXS5KnMJy5jh/
VgKPFaMLBLDg4tv2/2ESPYT5aRVZBZAj0o0V1YM85VkLd5D+UcgstWw86SngrebK
w+L/c5KsVfKhq/2ODnPdOvxLrU8kF4w1sg0K/dfZ9/ZAzs0mRCq5LC+XUmu5RaMy
LozJqLFBZoRtaRulUXqW6zfpm67CkPr8j9OqP3ZKy/GTOzO284C7NobvEK3V1QWO
P3ji1c8zID6HwyG/zVW9bE3XeJ7fvDb/YKycffqdp9RGyTEFfzMotTx1oAlSydrc
M/zXt7Agvy+T5kLQvkDKxJga5/rTaq26uI9zDwVcVK8ZSj60EftoEszeeU67/Yk2
wAnZCsBhwlU7p2h5t4vPRiZHtdwiPw80a63+qffmH9odlCgJ3ypC16+TFHinYr/Q
MJ22IGggJrnz2FvbBp7LHj0xBlEAp5jdpxDbUu/5ZupRKdzAPrn+F1edTnFKklTl
diRZqH7bk3I9xs+KMfS3V2YolYhGrr4dKGXJRhewWhRnnZ6L2bfDDKW1cwuy6vxE
NPfTgsP7uzJTiDLAEGbmc/GEE+HJEeUtba04PbQhSAndAqjbbax8w4dwIQ3O/tXD
Cz0SiH5hcuxUS73I2tk3buLhQpiy+dH3n3DAH2Wj9yZPQ9BgbDOXjVxH+lkd5/gz
PH62U+/qLnTyyFz+D/18rvSB+0fEv6qZB9pjaTnC/B6IFdh4bCDOc4/UfVxV2OiJ
NIGP5Z69QT9vAoJrtaCszoScjXzxrFi4b6Cy0P4Tn9jWlfSo1MkiQmXi20fXv2zb
m/v9VRAeoQLcnVc1lrT0zoX55jj789mzfO/iyyZVuCkahq2P4eO8IXoIY79J/5Zz
zWEW4O9ZFuPd6TjxTzzWFvXBX/dwot1pLnsr24o4AZcMifJMKOQ8Lb3h0h56UgxI
t+DzAo2PEQ3C2vUME9HrYXOAx41fcZ5NUYWS/G0pKVWDScOZUzgx5TdXzdDthPz9
mFtmSuKgSA8j33EaivZrmusm5dkIjLVxYCl9n7ooRRswS7Pnk+59H6oD+30u63rI
5w6QG193aEoT3uivoZpSW8429SYo4hKBifjD86Otaf/HYeNPQvMo6GE6Ef1w44UM
wkVXi0s6/+GrvOC7Xpu+YzJUO2kC0BUdAG/I0Fmv9AgPnCYThZplUmNU6LMtZuAU
BYGcBA3z+5Nyp7gWaeFiHhptt/mEL3P/A4h99FXXchIpX92j1LCAaxXm91U5P1lP
RD9+dO9l/xr6bCzChV1NN+mHwAPIaVhdCfRh0cAWhwlmcqq6TLWjPgnkldw6CQBa
KpKEZE/QVcNzLU5w32z5OiqCgGVGKu/T2eU8AwIPU8tm5vyG6ar6kKdWPGyPsDsE
m/PcJQh28r5GY3b7g9vexaxvDncRkoBd29RsNTMmotDUMuqMZLQEkI3RsT2nLz/d
oO5sWKe+S6V2RZl0nWnvIztw55V6G8ZIHbw/RMsx0rbuRCLYhNJN08uV+U//8QqA
NL0fb4xQ2ErmDiV6dSnFbtdZYJdu2hzM5pzZzduDSqrjNZxK5ZDJV9vzXMuFS8EP
D26rOpC5S3VvWMpm+rBfho37aIPmGx8I/1EAWGRqKyB+OO50IfK58Hudd5t7S5l2
/qKHpc4BUAej1trGCGaPc+QbFFokiTK51h6zR8688o9vlzekQScy9BSwU0gc06Jq
bN13wV0KSKL2SlcvG9gYfHBbyQCHuhWeRcEcA58/C+O+ZPvQH38Ckjo61ANxQMl1
VSio2Z9zrCeME9Kdy0GKZrGMyIEtMXK7qXf70/79hcbtL4dxk1sGlNb+S5kB3Qh9
UTxTZ1OhqCDp55t9XyXh0u6zSQmjKeuTwCvUkANGQj8voKKt1v9mUxUp6l5XmVmg
0cs5HmhFRb4NomAccVwNClEcX/SJNlUY3YW5hM4oBoubu9rLsK5VknlWIrsFdIFY
FxzY77GgkZEmrYKIwtb6EeZD9auScuViVcW5GaBSX/fepuSxnxdo6nkkfuscS5rI
VopLW8E9qKsjiCftSMAxbV0pA0aXlPVNdNdVHbBDrEVyt5arBsuN78lSuDgShfH6
rTA+vqW342zyl9N/vtrnjyMlTiJFXljO9joeoj/mI4X08WGPTsJhGkbQH0Qkaxlg
A8TZViQX3UZZcw68jfyFCxpH2UgeLdQiOtHLxhXPIZTP5B4uuSI+1OGwpcMfkUfi
101iMDWXQMS8PNElcwv/fJ5wieVbnfFW2irTN9hnyGEoQTaJ0olqXrujY3eVwZnd
zz6glpB8O1hV5p/azfI5KvQg6s0/q72WH4FXjGPu65ayUH2l/pY+8dMRtZdEaBGa
XVTD0JJYk5OpIt/wcch9l2aMN3D9fQZNAimyClvDwEhK2rjBwsITPms0q8lGc4qH
hU5jH+teLbiU5YdrM5jP4Qfd3wJA8n6esOd2jofkh6xyYMbSHyqTYreJOxqnBAIH
TO0qF0coJlwOwFcL55twpQsgIcgfJ0bs2Btfb/jM8iCfPsayR6B/5nduQ+sw2x6n
Anfm+3jnjRTevLC9iJFQoh82eBr4RFQxkEMn+/LCdx41LivnJ0UFotH/UD0DR3Yh
WI+bJcZowoR4jYKSBp7CGSB8kWyE9eNmbpio9w299dMlyQs3l5yiNu0R6HkKsjkK
53QzrQ+2fvhA2be1Rpu2PPqAtKbyZKKBSkoVcfa927BLjPWtG5hT7AZhseSWG4Go
026JnuOv3oEKSQJSgZc/4DScBuX+j5HVITWV8rVkJAq52DPdfi1/hIyHLV+B4VOC
fV89gX8a0kYEZpr2KdxW5GKEFS+Fju7h+FtbojB8ivX77rRCGEYu5r1oY7vSWB2c
nToXyW0rgHMNLyDU+ZdNNTgS0TGuDz8ja4YrKyRjwdZ1W3Bk4cTusFSYR4+KliFX
VINkP0ZoXmvh9rcPVHryt/mVm+9vvn9AfS8Kn6Vfb1uw3wLRLCZkKzqeGDxd/jvn
r4D97BsCRoKiV3rmOLv5p3iSn7kHu3HuWEXObCrvPmW95spiHKqI/J43fcxRGZhl
vUXG6/Gs2XycRvG/jZfWiv+FkwFqn/bRL/BjwK87nH7sRd4pUUC0TvGV/BeCxiUb
YIiqeGVilxkutwt8GupqIYldCPyWZOe2OXETbqm0iG3OAfq+j8MD/x/Nkya8Jt2i
xbfNCF0CG964W3l/yM5zL/4KJPSzZOI09Qi0yFyUnSOKQMh8R5x7l4jk2tkW71xL
dCMwPgu5IHZKJWSvsXaA4L4EwxH0Ubv2kdA0Iuc/lulBuf9Hfr0hQp2OIxvw2rqm
SGPwcJJr+GR76OfXhtgJHTKMYhZ3FRdccHWeTVzPZyGmd6m+K2xTe8oYO/m+tYyQ
2CvZfwC80Nwyh0mo+oWYITQ93sfb+soxYbenXzHQfymRRlzPlo+x45fD0i4Ey33f
9KwwMXibuIS50dgx0/5bxbP3X9tZXpVRFt5ED+QdAi4mAA4AJtoMG8sXWoAAt6mS
tVDaXuNRBPrSvh3vQC9mOvRT111Qh3gJsLNxgv5u2kHEue6Tagp9j4MqD6aRcgQQ
q3g/tpVmyzcrBdkbwXSiCvFJ7YJVpk/g4aIFsBRHAh31A/hVfR39X4hmWD3Ipb76
6vQzbqjxkjjd18Rr8xUlqON0dGM6B5b0X6MNwZ7QiR1tayiZGV6WzxYQjJhFLizR
bbv+tS3hktXhtrcUogsj2FWGZbSLO2CH7vhRG1hVFu9q94CSbJBfja+ofrFJA8ra
dLhlFNnc8OeMjPWnG+/Oro/386SXHdsiLGUNMbWf6uSSn+aL3iDEszfZOp9TLgEi
hllVoLCrQ5rh/HQDmTOaA+1gWCXHQXylAfSpaDx6KoNkI1n3X4hOBuTx/+jPztVZ
Qa8darAJu5+o22Bpibpu5i3Xk4SLKcbJzVtulmPzeWJ+lB+7Y51t7QbLS1DrWMYc
pAaOkc+sej7e9Jk3acnbWlX5hP5sphbOAiZYNz7ETmltZL0pT+z72xtS1YQdMcTm
OXJ97EX/+PNQ11iNFrX80iLCj0JPLG6mUuQQcOWM62IYovUfYXVarYQGj+9wS+/v
1eK6xeG4RQA8evkXyo0eLh5C6vDKCgGFGbmIpGclvG73RafMOiqBvppoAsFh1Nnl
uop9nBBEqSP6I3RWwbFOYHmKEWPhGEzlsMsPDXjDnMQ7CXEEy8oBEAm7nOy75rgN
dFSsgVvsrzp+wmIuByUjscBKYUVd+BIC8gVp31i9qDfHDcpk9eG7MuyUXQ78Jby/
vljenD1T+BeK0NKagVYb9uFbaDRLB0H4QRl5oDwYph7iLjm+Xcd30w2vf2Hd+tCt
zC7WZmux2uLyKRL0FoAeU8EWR3CiFap+YnB1UsrkVh5no9wfbYy98A+euFEOi7yp
TY7D0+C4ORd4KHEacmRsSId8HphGyEG20xyiM5Ycn0ZTmKEC1xakK9IMu7wsyxSl
HPGx2gqZGDGcdWnAbv0JUvlwviL3P+jnvu6HVR18PJYO9Kssgp5yYSFY8eVfh/e6
RC/DNXt9el8ZHtWgoVWMCb5fayu9vA1I3BannKcR1BlniNhmLoaLEJs8CyP7hFEe
s71fHUrMDWIAJrHUv5FihfAmVZUUzxElOzPjfzssOpa+ew9j4B0NEWNqi/2hxGX2
zsnfUNnsxPUyACyQ5XIESz+RSUfV+eISUJ74qgSZT3YqV5Bb1JjRXEUmvEEmsS08
d660BuDpc74U+Ngl8JRXi1V6ayyidKWno8cUim7eD944hyNjPe5wwnb2GUgncYVQ
SaHVxXMM6WkNsVbxV954xlWnDyGayUpQbJ3JpB+6N8ZNWFFXsne05M5YlBnXCmG/
s+5aRH7GF4A48nJXHlklCHrFC0m4yCv/rP5WO/TlBkQdEO++VEFcMFJZQvSCVG/F
3MR+zNRB/2tDPhvV8U8X2hV6Pv42jRPgVmaPSVEAn04FdrGB+6OlIhApFEA5X2hO
kX95Fp6BM/iwOpj0kOWx4ynLlekDD3OnpNqR+1qaQ84xHx2U8C8vXSNYYqy/kcWp
4UGk164s8oDKShkTV/bL1z9E94/ICustU5rCvcYNY1yKkUabRW6doReZiH2yjDD+
8aBiH/fIx5GwsHegDP9qH/pAk7siQQgDWXbWCvTqe755phtaS1htsxDv6GwKkRys
GVq6EZyEoryM4EFij2Fqelb+MLulGP5pcvz7USVLe5Eg79ApdTmXaWZzAI+5Tgp4
tTkiQjGN0PQ/N2KeMbz6BC/ep1UImT/FrBagJj6aHCT8xcRLj/e82JzEMz1fbZS/
rSsX+LpzCCL/1a7MlBbPh0ynvErxyKSQLBY1ahiaNKy2Bk9+ZoVKuzVJEMMO/rlx
s2DGjWkJEh00wUni/rSKvW+KVGNFZz5B+xVIiOUptks113gm5f5Q8PPR4crDE1Ru
IkvvIhjS0XYqr/2KKOekMnADufkzMkXmcZ9iXM7kAazuiJC3bJiu5PjLEXoCbYQK
s+woxYWSZdll6H+R/RNzEHiH9IQcx6u7oxI8L91ZLm7nPq5H+Vf1hkZ+PZMWTXOj
xyBGOgYZLQGYK2FA/i4jPfrOtouuzeYOxcZAU+Fi2ViX3wpdD/lQ3+bIflZ4nU9P
OewcfBxz1gtRW7UHvwS0sFQ/3Y2T3Ah1Hqk4lv+b+eezJW2/SOAun9yieAG622nm
7TubtWVn54EOi0LI0kVHYk+9tdnOZeZNdvdKHir9WtjuJI4+jgLrH42/Cvcdvc3o
x1OrOWn9i1IjouOGb33s9m3p8ARp+GIIWQ43AG55qldvyJf7SP+4cVm6V+wh8C50
vBKgX+592qwlenySxSFO8rIBWkBjwkEBVPNKtJ3UC8jAjugvGO47I9p1HegBcDZX
tA3raviqINL3TNrTtM85oez46VfDAW0BNaQkapoQKFfHlCS4QjUqfAJp6SgB9juB
cZWXXQMN+IEZftKQcj+ovL6P3N4T8q0XwBJvhyRU48Qr2jhDRVJ1v6qP6m7AjLr4
0b5bvld5QVdeGh4Wlhg74vABj0g/rAMpxu1Ngu3IorDB9SHQwtv0TGmty31uuoSi
zBYhbAnDz+7VkGRI6BbSepUt7NEpy56k+bXyU/BEcJajdRNshmtzsPKfvYUpbUwD
BH0tcIH5wM2kyvSMcpDEsQiZk/tqJe8Mj24K+xnNnbwJddanlwVfnaTjA237YRND
CRlbGnh0eJpsDTOUoFCck8YyE8UI5IVHLL3SheItH0PqEvswQjxBoNo909Tzw8ne
/v2fgHlrxcm4CD1sDHgRQjsqKoPgQ0C7IsA60ekKvEvuyzuxwBy+AA4/vem3bSST
ZYoKXKaxu9fKFgpsln31m9JNTkCAynTIidsmZ02S1krCA0l+VjH9ErqDifO+0MJ3
QEwEwaVrJhyd5ccNWETSvjQpaRtn7f6FRtEIoiBQD1LQ12CYztTZBc0jOPK1t7FC
tSdmIDywgzg0euF3X8RJOYpcMQzx6AO75sCZFj3JW2ncX8bcicAYGouDoQ7762ds
X+R2ePe+GU65W1UbHqB3QF6/dz+OuFLHAeceQjALBYvpCflgEUVmeEm4TDr5N1hm
YLarwS1nztwQf5mvrC7MjL9jjxSfRuAOg4VsBDLG6jEV4yMBHWH7nh2ppl5JnOnK
gn6t+y3Tk6WVKu4t+MXfXk0QXpdQ/6423QjD08ylv/21ydsI4HvQrAYkHAaWpr4o
NGeuss/aCfa68a0xJjWZSiAhE/uiFep13nONR4bTeKNjf0Zru9GmKJC4F3j5hz+V
Bn3uxdfgl5pc9Spz+SiXJYb4zLnL5tWpS3NkAZh8vqgoE1U+S4QUqjz9ATUs9RFY
KjlrXylDOdEI5jaTIJIge8ps0jRgPsKFDBN3unLSQyDbW/h/uPS0iOepPY/3EEmx
y5hmQWY4JUyg6DBjOJaZuoAVZA5NSHVUt1gX+FWrfu9drutM4hy0o/FpbENO6mAE
7IZyEYikhx36UabWOvM4Hw12u+gBv4EKpTveDNLBjQizQyOSpQ9X8p2cLb+6gL5B
8K7pjldFIdYjc+/W8i48eXK+zr3ZPGINGR4ZINl1EWYkYUYIFbbLthZw5eY/uAKq
1B531xBrLSmyUIk8x6gqi7Z4W4jXY21HR3XX81D35n0zlWRurt9foTCdP0Qmw4xm
wfSiKVSU5q90GaMbtOd9dbK8hKlmkM6KKQoUdDU0hmIfaaN5RqyFOosKeCTbo25A
B0IdgkQ760fUp/jmYJ0mp8rsoJf/bCkgdYvzyCV+0PZu70YVdbhvdkd3Wulnp0Dv
klq61GdN18uFoOCwzO2uofx9md/zWucw4RlK4N6zmgtl4BoWnHruSaBP13ZmcXBB
7K18q/hzsCMc8eFn2mim4bggnsfW0VVcDi8KzPe6Ew0jP9hmZpjG4OAlkk9//VqM
Sb22LMaq/WSTNICFB7l8Xkh0x9x9q7/mdzWxFhgB4pa+TP8Jw5mImwsC8q6TodO2
mjmwUMlbrhbY+OWO3HOxFPjQubCe85fZUfHLktQW2jYJo1/Wwrwi+IIHuRHE4Ss3
5uEIJ61bwnExX6yjSoX/7y0yXrJmCoDXtJ4/McLJtO3+iHoYLy0thSv9+w01b0qC
4Xkj0mbRBO/TOneiZ7TbgFzpQmybv/bMH66dapeUHbpWl8VLHqI/C/MvEweMQdG3
bnMISxXj1F/0ZxWZJMNxEKpGdbnrCAiln9ffG+Cqp9nJLpiaySqqpgKhFohs6ns0
M7OB/Tzb0wIeS7ZwGrmx3ND3L5o/d3eGSHQtfViECS8WYyElRHFxfvaRQmjlF5d3
O8ppcIEstzYx1lPcIwWQBZy3d1Ga8XMsxY+rYL5W6TOWq1DhleCwOMV1HXDw0oJt
ZN1o1V9ka7CISkOtfED2jsmSKgq/fL02zqU4mWZA6E4RIOZ1K6mkVBaiy9pBy3pw
gb/4/jFqwJYPfvwV/b6b8SPguF49/NdQk+TnQwIdvjDJlW8sYjbeeACaMA7VGIOv
3+d7hoKsw3pqUkIzMz5g0QPOXv4w6yp90phjvOYq85RdADxUtCLxJ2GynMxljQw1
vsZ1iTjuojV857yzNM+XFM3Q7xLDds2/oCgyN1eN7OvWuFf9nKkXNkhcf5D1f2Ve
qHO+OcVhLRKHjJALbiWYhAwOjybkYyWRp9yuWe5FKleUZAXJ64vPAKAq8r8Pa8Xo
YS6Gm+nNj7lwbimPX1fjPDzvLO+Gy2F0Gxjf/D79srQv4ZxBB6tivy0bHdDuQ0s1
pfq4ovUy503oHrLdG9+y6VJclWtQ3UTVkiIyaWMW65jMNx0QaN/RT2NDEwar+/75
RSXlcp7DJMbFtMzpnYFKvKqdpoHDzP1iRXkUHzoZKDY9hPwB1VhN12W56FVLcJT6
4j4nH52jfc5kA6ANOb0JvnSKp/mQYEW2KovS3X0H/dC+6MLOsw980MuoMzFc9Wi0
BQKJPOcLjrziwJPlDH6GYO23Uj/LdRGZk06MnWjqyaSaG72GTLSflz+qKJChC8ZJ
84MJT8zzBvENO33mrq+S8OP0Qu4dGp4w56lhf+c4WY+Y+EJPAFSNOLLjdhxzKDZz
r9RcVCstkESjxxgsRO+xacBZ0RwP6w1BqmjJX8CDON5SO/H47wUSMxLI+TuzDBef
OOQzGjYrqDafmQ85dhDOBjY4yYee4H6V+WYIKCS/H9dnjPBr5C8svGKCc6oNtAUy
0hdaIYItG3ruevfu8kjUB5mySF7nxyLnrHoVobebhMVXe5aOoZSfWKPb628/q8mI
fXDU2w3wgcCOhC8Ndwd3fsONV0wAG7lxUhs8KBV3lVXrmgGnT3T10FPZb/0Fq88f
FJDfJBXYPhr8uEjQFG+DFwf7M0EdpC02aQaNJQW5soKJfMRBAZZ6S9yw3AoD4WfD
XrX2LJ60zPDAcHGFR0oJ9T/WzjY39NiG13UUhT1dtvW030dQjtBGrB3vFVNC7k4B
bATpxYLddODbKJx2mcuqGr3GTgRKMK04Od0MRPUfgc7R1IIOs1wwkVyOYoEr0/Mx
m4u3evKMzxP4uHOnAzgfPDC+NUueSFcCI/rusnE+uyYs7la4s8nypHq+EMFWIope
vgPcx0pCidxeRnwZFAnqCzA/TA2Kr7HU5WLsYXAaiNF7U3i2eSgdDPoGUFGEVggu
NGyuA6LKoBfB/ZJ78MaWOkHb86/d8gmYNWvLMEE2zhoniTmyZ0/DiCddXyZI4fDo
qioIOD7XQ5ldOXCQyegUQzrrvNw4zkhiigrff10eK/5d/LPvsdIT680C+sCbrjy8
qU7uws5mLSj0sQ6g7uMvwD3G7VuUaSdSFblzC+UXyyXPX0J0yosBg6dctJaHpOpc
7Lvtv3JCjA4iwh0XODspUnIzgVZ8CvIyb7avXCKLe/sDJzrM7N87TvUSL2oHOioF
zAO7+fVvPX8v07Y5dd77FY2P4fsiFOJpz84SsCIMZCVy6HEGG8t+3vECSHWUUiMd
82J6iLYdUAJuohwu38Pn0zSpcK/Mar72jR0MagdURZbjKDjEoz2l+CZjn/31gub7
k4n/kFE34ElJ4TYCsPUM42kuw3OMT/AdEEkbtVvH2CYEAdUHxq/G+yrdBEuGO4sK
B4zgh6eyE5MW0QMZYaXyQ0N5XXyg5UdnLFEZHFgq71cQw3ePpb1ncMf6hf3S+LXd
X2H0lN5IsrlPkcsoheM3zfDYrwr3XxWTpWCihgU7IGDVek+6yvFV4QZ6lNGW9UAd
UFTnkwwF0HcdwAWEr98ihgh6JOg2tVFi4NnSkosnf4+y5cRGUqI9PDJiIh2W/RW+
9ILuWfE8slmE4Ivik5zgj4T6fmmq4llxaJFV+M+OXj8qLG3s6zYjUU8EZqiGASmk
lD3Gzj9RA9dn0gmxrX4R9SnQt/VyoMsM9qCQR7TW8n79/P98roIM1wA+P4R4yjZS
Xj8q0XBSiGxQ82/t+CWyZAfYn27yFRC8QGi8CQlWbQtzWbgPdWBu4xmR8UcHSjsE
lDmHnjLkIIru75E5YTf0yTytggcPXSAPThnEWDV1zofDn/HHqnq6SzkSxWMre6fT
YnsusnhQLv2tTHP0+hYoresOhMD4tCepy9amR0pHZkFsdVNJgpLvt2ItTu/kvJPM
i1lnl/DqzcZg3bvAWRESePszytFSBQDlu3FoD8upuX1w4hboAJv944fD7dOaRxnW
ynMe88wi40Y58Zs30x7axtHxkc+ROYc7s1QIbNc8KdW2K4OZWNKpjPDXnSm3JLvf
LaPxv4ffwYLdXBLvMsEgkkEtestNDJX+XtFDtDLPuJpM5fxhxHxCE0hzgf/aMRVI
uKj4f95VRDNiDTd9mPbqQuYx5fFW9IDdLp337FFSQgKD9Jl/lzz6L4XWsNIlH4ef
mYFZm+WiINFqhsO+saioVNrXFyyu6JpzLZ2krnUAXUMEPyZoTS979Ge91jJes+Em
7lNCEdGFCJ6ZO/Fy57ql5GCuhHGweArQ8qJzQMmT7GQrw1+iuTHYH+D1ppq+w7zY
3m+ZKSeUk4tVdClY/+sDMpx4bVrou5gS5Bcm6dJ4shdmx6IPA6yGaiXs87BYn25/
AETS5VByAchB5zSeMcNi7L2Uvj+ql/UOPwqkzeNlyBvRmco4VT2MVNA7Sz3Wd5FW
LwhQJsc8Zc6FCpQwOjUI7kb/E1RNxZ1tfDOIFES46/Mg78qtshYg8TPi4VoS+gI9
dLsAYjwjW6XQZkgAmAu54pSYZ0J/LRF4Hi7xRShRm29/x4myn/xhHoe/Ap1tx138
esEZcmv3vpPkHJ8h3kmhi5Q1xoEIigA82Yv57SaFoPu8ewnLx/NtuOImvTDYO2l5
/I4Qh2zUdHERyTX0zCViy/9fLDYZniy4FiYYDdpTuFMTDksMC4mVakcucAX6Fy7w
6DJRtP8ga2vHc8ky8rCHp9iAHTv8wTC10ih08/MSfI5W5eBlqV3cKIunydjeoKTA
Z6+10730rIIH6G0NhnTXNQGM5Rb23U1K+cMI4M0DaM4/wVEzohn8uuhjPSS0/0r1
XGVoUQLot7PT79ji0UK2hV+WG0r/u2015/LPmr2XIuQ94zMGUenKt+wzx6UIYf+k
M8cMAa1RMWrR/NJ4IlnaQAxZQjI5kkOSWSgFuJOfkVTKJnuYL5OIXU9B5ZQHvzxg
JouqfsWKABKvnKPbXNPqBoxPB5lHNFo9NX8xLfy9M4KVLJ0TApyIor0MqW1tz0jB
k5B4EZoQRnWx4bFg5759c9r5Uf4pbDj3o/7sjTP2aIBG0KnfSZ4jmtNnSJC8cJOR
D8ES1ckCpsFUAeTTE21DX1bUmIa/3dT7TUHxTd4S8zwW48EN3xHYzkvwj9Dr90xL
BgWYF0J+WQWKdu5rQYScal+2AySoE1q4yUPu7sRSr/8vCFDmYnIWa27DyAvDrf5T
SbbIo3J8kCmwlhWi0IvrKvkH9VRk3vLtBaFUgtX+uRE6BsZTF2vamIFLylPnT07I
RHNAfl9HZyl/SMS0UPStgaeEg1b1qG8vptFaJmzPpIxRWmoF7U1K8HJIl0WZKBS0
VFEccXarLBvcO9Vm4wctbn2UeI4GryKNZRLdGvmNe+PfxTmurNCEDG043HyNA8IE
c0WYb2FjOP72tkCyUF0UjwYY11WI/MRQUQvi7qriefBTMuInYLpvzpAbju5SHFHm
ZodWVOrWkKlfFUmP3S6PFKAksrfGcbs8SfqcWu7fAXgN9V6O9Us8TE15XAWRddrd
hlp0ey8BmbeUEyvHHb2LfQS7MG0pi26yQelQtNzZXwMXnCl642lMV0vOJ1qjNIXL
l6LPEaAXjcblxyU+AtST+kTGxdFVL7j24vfi1jOLEjpmE1MPLFWTJXkH14Kbo0J9
35xU/EQzWjDeonuk+MvMlSyaGZR9G2TGF9ZR39nVdIAD/cOMRjzZW/qZNmrzcEG+
ZehAsYrStRhUlMOlWLZWNsjM/iMv/TeD43kQzU8y/WOnzOx85KKH49LIGTNF52+q
rHo9RlrjxCGIQUOh1ieHwDR2+8A8CtZ0WYaiu0Kl4hPEctM/x0K0E/fZdVo9aRPC
jedEFYOnO54hp+UWfKhnpc32j4hbziRHQzhzoiY3uvAWRLKgpSHlef0L+OrzNwWd
ogG70NvXJq+taeQ6pbG9katY68gU9oAnaBcPZgT8r1g/GZjwEUQitVXL6OAAzKoj
9NZhMtbY5dbCd3kHU8/Wrw3fpzt20/AZe4XzkepVS5LzxNOZdA0B7FBs1vstExjk
89y9MGN/8OJSOTgTK8NdDMGWFHXWsmTPrEoAo3WXvAnv+L6QTdmtTA2z1Ujrd9pX
sry+m3X2EyVDHHWIpYZh79mY3G82IzQnRmUSHMuYxS+j0bumeYNlbn27fvuWCII3
DSq67+zAbmb7+Q3yMoLnhnf4+ptGYzW6fs+v2LSYVQKIYP8n8z6zRkKrqJYivEmb
6REAz0MGRHiGDsTzz64GOtt4ZSjHirw6cbPqpOu4s1F54nt7cgOCPK/mfZERf6yb
ZEIojTqVqCTIFckBSbEhueW4YKAFMO7QctrRH6HzSZvPRIkZrThMLmMAkZleWU1b
n/PNOB6pdtEvP0E6x50CdhkwDeIivoSn9O55kFAZAlzOTDFVPQE9RsO8JpfJ0yZm
AsT5kMYVBo3yknRObfRsf2shGpjkCSuNDnV+2w2hkpM20gu13nGIfewptmkaO4AU
IaO1knidMmHhl5zi7365N6PH5+53/62ilA/FexF5DxNRQ1uhq1K+V2kv1AS5u/iL
JTOmwP9hZcsbR05kO/4QrjlVPr3O7lMT3Dj0pMJ3yDHg5l+AcSiPx16qrOOswZgc
hkc9Z6YnFei207tSIG3DLtB0pwVjcXlUO9snAOvEel6WF9foURmoOF7rjQ6d5Gcf
3NYH2fwIPzPHSbxEmc7hz97EMmfGfWRiCUpgiZKJEYCb0H4kdmf+UlQmAxikQPQH
nzlBp8Fj9RNUbxJAIxRZorHR2TmlZjgMlHedShvhCpnxzOpgcxy6YVymYQ+lNSYf
9h5TDVXSj8F5rlcT8N8TcXfrAJJEThfSfnL6eDdptlvnXQbNnPzPOCMabUgwLDFJ
kKjTFSFCCYJRezBAQ6RXOIgPUbuNmZ17EKY6zjEfxI4M5zy9HAN+tx72xVS+HosC
VCV2GtV6lN6wynpuOS/cIr42zBQDwlQdfovrZgF/xt7ry0GqHrzaHJ0vyPGuwIT3
d2LF7Mjdcu77S4gS3NacbCCGfG/I7s8b4JGwBAvG+zl5WqKCIHoYNAejFFRyMCHW
AT24f0iCrC3fWauxjBJYkzL1eRbPXG9E4yVsDDT8J6Mz5GQu3hZLUEpvseBYQiLm
xbT/wLD47DScUXCy90uCPLXyqYM3SIuskToy40SAgYoDvR4x5JlGBLSFMf8Xtila
daHhnTU3c8NhHtVTolWyFQdx4XXSWcfpxW+42EJLFgL9xdf3X8w8ui2h/R1qBt61
iuvIVf+0TXc4Wm9F94xEah7Foi47Ual8Yo4qu9d9HJHYb2VEWZgrokSyXDBzDioM
1vaMXCkYJcZBNbPcl+lFYAhLkSxXPw7LUo21wQalx1Vh2ZovdfkVeE5xj6TS0q8B
46/XeGrBdr3XA5HrVYaxnIHAvlXx4rXxSZvhvcXJfFJdXsQ1UsnVYJlwPW4VzPH3
5wZg5666JCCD+HVRr8L0FU5E0G4Z9DrMVxDDiXSMLra55iHJitlBlZUUboL1yKcB
tJB9oMFJ2Zi7P2xyMRPIi7nCAtwiFz0njOyggK/tA2r3A7mYh8pPaAAMHAkU3EIa
ynZ8vmsJWQ+7PXxh97i6LYGq2tebgj7N9NpzPojzjW+mdKjcCHYtrBZvL1CnNotL
oitPR32nsdrKphUZ+TKjv85zZBxg1Ui1aHVezqJW+1GBH8uvP5pFAim0CcRfaGVU
DfnjxIQd8PPShqEWJoE7Sps/+m9p4wr2xiyzl7AG1MLQUV/n70wnIlHwMpG3IOOh
h475ZALgZCcG45W4QMwqVKzLLwJcw+brjG0hEoiXxauiQZLOlYBIfHM2RbaDbomE
0VdwTCmRJwaiF1p8A8+YN0ReHeR6LL8jEI14MynEH/AasEvPdk9Ooi028kYTrVrw
qG4LWzq9d0hUWKOComsdGTpnHT6T/KqAeKNpsxL/lLsFpnptAMlWqsoAOC5IGn4h
xI0N3bXCiflj3Uh+v589Tp3EdSC2/UoKun1LTIigWh77d3hGEIPNPGjYLGegOpOy
YYOxnE9z2R4Q8kAvNmoR3fY/3sa4TeVd/jViVECTClqnwny7tqJi4ozDF2ZzEAU7
Vfb1FcfuLBtdRV8S5ajKlC6fYsyE3XHmODlI2g15Zvz/Ei6j6dddzaMKOtlcTPLF
n/7UcAemRa0W/rEKOKCKcV1fxpvLCGVUIiDb5sJqxJoqUKOGu5dEO97lYnpG4uCq
zrp9+ehGsXp55LcNKOiNe6/ZwaVEuYvdEcLjp7tKETUcCGt+uOMIJCfBpn1wdTqf
NL20lA/iOFUo7gwnX6NeKcwnpeJ+en+ek33QWdaS+2AJstM6HPxIlqnoC2xwW6yg
OlW9ZtixmLfaM/xRzivVYWpAuNSxpVfFfaOriaWl1wqcjT7ysZdsqxpeDVbJKGum
/mjJ2R7tIH1Ypa/xgkBBzH/mjcnqLsZjOdCgiIFp5DYLAbnH10bHPtUeuWozz2ZT
JAz82sIyWOl60rThQjsNZXSp/B0gbvHHK+LDLkHtllCYMgyv2dmrIRnwxTf6AD4M
I8HFM4rDUTuUgPH9A9IW9xkqhsPwxSqzfnRrNGO0XmP/VnVhnk5W9/z80J01ChNh
Cah8WG4Luewc2gabdFaLc3ll96Ny1bwbiP6+SkftwUfqucsR9fnWRm26vCmrnhS2
ltTm/Dz5HM6KUui68kgThmNTW+/id86Lu0nuuuv/NlhfjXmeFAEYh8DxNXhMUfMq
0BuyO9BeiUwpEQcmUE+Tb0v0hKJY+PF1eOVBM39Po0sr0ovxq1Yw1UeRc2KMki77
R2Vdu9P1n4/eyLo6NoC6QJteeozTwzrPAcXqymhGmlwHOTlpy0awUAAHXsCGB6X6
FJr+2sJNDl5NjX2ZbWtWWIvDHJDRAfHVBJNtAcYwCMtB0p/0c89pnM5hmRyoIkz8
g1OeeB49T24ErIoaMl9BdREZxSpEdRqidqWKdEsaSuAxdB3lx6q7YPwqrHP+78Xu
bS/HvWiQT1pub4H3+EG1NQqucBOgF90JM+V6ZeAqzD6SCGCZo2ryVsm4CN1RFiyq
I+VKotsAZBhMcONHYmIJyP1K07bxCtWox1Md5arIa9DsBo0/Uoce7TTNJL1YsgF6
68pTpGvfPEqws4TSY/TDQFAxjGM8w9YHrsG1/YIcsx5XfZAFhxrGhutLZL6gWpx9
2GnsKKad/z2K6JtBdVzmD5fcQ2papoyrxBoyRqhvyGqbWBWvtl2aq6MNqST3mpis
Gg8sfG7uObdgKkSrvkqlxBIgYDMWQA6199BXTnVyERJFwXPOzlLgDy2K8ee56TTm
DBP5053Yr1FsN726xrLXv0s/qtnQurVS3uhrQ5MjP787yuZVCYe4VNOKcDqxZk98
OJJRdAHLLHFd2Hzu4dxrSt0J6Fe+2CduGXNeRsGooX51Hl3VhvszBwsuzPhs8UfA
5rzJ/hCNnQh0MNwbe3uguYEs+0OjW4mNdZ1DIE9x691pOdFnQw9yah9rXhrVIYgs
p/c5NDmbzpFE9giOn+izAGxa70gdL1HuXDRrEyDmMwsvxkHUK7N1lU3RujsOtQzJ
xIQar1L2ju0eNI+mp/th45WSLFWUEb+DHL/kOglnAlU1m8TahXTWBewfxjL6q97d
5gxRha7YPEccJqPmXKgohPlIeWiWrRFzLNLGiA+vgtU6ih+NLsVYswarQfWcJk6B
L/06HzOtR13/nH9YJxNK4P7ycTw3yObzW+kyBtPewlei2uPIiBRpoAYji8iZHsy4
2Vgke8HE9SpWWDdmWVdwiSEFaOEHzeXz1WukHrA6NRzksNUxBMxnYBIOxXi9ZzLy
pazKYkes5fIYYY4C6bpgHDVlTD2ZxcTN0wZ5Y/4H5Z8mIrirjyJhtsKhgKaOoLQX
50+bgx/7Df9NGS2NfMgDpsC8q+2IX4oxusUkU4Ip4rCvxFdnYtc7QQ1SrDKXJBXL
b68R4x75XmAruPfxdoUlUdXwVf3DPVN1wksZ/CW/BPKWEDLnst907QdYOftdV3T2
gSBL/i/xS4MyHk27HAmPqPugLy9+Rfu74zkhSsUUXxsPrIfZ5L5I6jttiCHDz3el
CUDG4JsHLxPEr1/0NrbtM87+Npc3j8ODsNd5Js3AFfM8rinuxY6PExmx363wGjk7
FWxl7tph0H0/ukBcy05TzFjCvOaNu0wP/uxEhcRfu5FkmjF/v4KY90U8yR/Ky7Cw
5PYU1YUkYa3HInIwg5S79empy4tYwYxVTlDJgu8OAutv76/9KxNDgcW3iayvms9s
k76kaxgx6WGg8VIDvFcU68hz7cyTXxpoCGHy/gYXj9vhmQZatqFsvRpc24TZ36OS
Gu6QQ/i04ERhoEjTcHr51ZslRE5a3KV1AvVMfwI9rr62gRAxF6v/lkEj1dX4ZaTS
cVWbE+2BNju7Nj3LDAZD6UcuZMrmSNupzrTdbjfd67U5Wv8lRaYXR3KDJr9SQw1d
Nt9xtckv6BPqnlYhVdIDAXCHUSaVpjJqZ4m37rvaZSC+nRYQZt3oRWamDPOxA9uL
e+Wg2zlRg5AATNn70c6w14pzOmPStV5yK9TBOUXYrChP7Ftfid5SjUBHq0ZThThR
d91a2Nd9Ks8qnlCmwbsBbg8g7a3uzu17j419JhJHB7+ij4MyqmuILMMAtrwLm6f2
DxxGRUQoFOi0N3lHfliG5s3jIlvsJ07IRyRxIXylGPhAJ2ig/5DxRMfLorTOwWYM
X4Blf6pOuLoi0mlQTljUoLdQ49fOPE8/ZRc+cvYx7+r+CIEC2MpavOct0ksboLGL
gy6n7h/Lg3LHl+wQ4PjVAHfEHcYtQ2jnv5I/3V3/z7bZvFM7PlWP6b+v/NfPYoAW
Sbb9TeMYcccXYeWNP89V1MNsFB2yOUQyixvcJG83C1uiul9vHMOcRYYUgnXZ3ull
DGr08z4wSMFC+DEA4zzBo83Fp9ZLZJCefgvvZHzfTce0fjjoDi//ufTq8EO4PeJQ
WS76PmULZfn3zYX7lyQzGW/AtOyE818nVr5YV+CLidmzOicSR4EG+H4QtjJgsbm0
tdYpf09yeFskSb1WcjjzNhw6wGR/WuUtx+T3WTF7MPfrdNaWaRk9wYSmgy7DwBmr
Q96Zw626LBmKe9MCLqXDYen9NNu1GdTu/xep80PrAchCBO3GsT66SmgEwzwV+2Ij
weZJC4ZsT9hqot6PHuPqcv6tEh94r8xwCEHoPNFwQ0xSNHstSNlx2SnOq9EUCGex
Jg5Xtracqaenf7ihUMBxeE531IPZ1IxaY+Jq+IhhS6IR/D8itWeg5wUonmFPF0bH
LuTnxTRAR+hRCNWG4r5TEEc0BeB0y/RICO7/yjoywHiLuHuXbecyqSeO0e9N4KbY
uRwgl7S3KBL25YyNCbDlag3Xn0kz3AIXkoFl91VMMotXLojNmvC3ZmENZ1cNGpAG
XJl1Mr/QzHufAxAV+NatHpo7S4Z/XEGQ9Casl+ArHKp3r2kU8tK52xOpOheZt8s0
5/VKtANGDdh6m3OaJrK0Y38+LRD3Lv7qelHhgxm7pW7m7O4UtQzoX/cQavEgGjYg
cTO/G9gU0okwiO10UrN+p0R12/Bbt8Cj50/mHi6WSXkNBvHIHCzhgEhDZh8DpmGO
rN1ctSbZlGhnCalQ3gdFL80kjYmixGFn1M6vIVonp4c5MYXHfYcPVL6ZpxooD6s5
MqEJYbNqJ3w/TaUPBUaGiZiLzyMfGc6r3hzvgUb9UJuSEw/q4NIGLJfBQHK9FuLC
T5KWF6TaZZ0qcWlcKDIEEmJuJ9r2Zc0M9xuhmek4BLrUb60uo86G5ym1H0Qywo34
UthL5aY75iNtmF//gNCTdwzbWpDaw0kU3LTip3D66yIMfrhdAqut0jb/8txYixrj
F/c5Ij2o3OrHPfX4v7SBNeIp+fT0IRacBTvg657KA3N1WLECc34JC0OVtFejY+SS
U5oxeucTKSO78aRvxgy/U0bJQvPJlmdZlkJgiQbPHj7XhsAWpwcTPe7vEd79uu+R
UGvnr8zPtHgC9QlkoAjwCGIAt+4+2twWKn3NcKGGFbyXojEUegwJ3QL24/7/S54Q
fjdDzE3rfaxJNypZ+JMS7pHwrnwHzZ8HIGG0m5H6vXdjZrIGnqF475cjnqgrN/Mu
06Emi+PBiF0f9xGgLDp8BC2wEjiBhckqb9pxPIQnR+2NgM7YeyXt3omZ8QuonXsY
Geo4ArNSVuYm0PP5xouHMqdDPKE7stywlKnA9QXiiYQos5qPMwkLR0b5y1SgVjf5
S8i6f5F2rAbOS7wJiVEE+3DwpZ60wor84+w7hwIzU6nq0nSTWuLtShUq903Iq540
IfcQc7u6NirMRiXV8HCJK6Py2cEp7HOU11o6jBZTgwyjmEggtMaRGy6E23y1mKkc
q8gNoeOZ8zAH6WtijRTSucZqMXpjnjgHE692xv2jvgUL+m0k9BSPnn0cDz+8YXLk
NXnBdKi9AFrDamB4ckWxEdbvZpk9qqfMsWelJQCugF3fNmByO26OP2sQUp7jUtvK
Sez2Or6HCs49kR96KNLmI9LTXukPluv5ogkdKAlfLwjHguBgQjGusF2WKTdiBzSq
fe7x2hxo8E/MWedrXOQBlm7PiC09mt5rw+1dV/hv11peoXOE996GozfvwUd5Rbkr
Krbzdn466jCvwDHzQtiYhICiwsAsB5HzMcFK51MAhFhcuw/vGWkjjuL/1nd8u0O2
XuJ9k8cJQmrNwd6V+NWCeoalz7BVr6NZhzPIVlk0Y9+cuECSBzUbOOXD11eNCM9s
xtoMSgyBkIYvLs5GI+E08u/sEOA+Fh+wvs4aomx3xIvFJubeKg6DElWHZDCWIfE6
PX5beALbtHiJjze8W2B2gBz3UbwAzBCGjTn9wKMi02SXzJy+Auw1zLFmcG7ptWJ6
e2dxBcTfybyOBmVQ5UfN47kCgaoYoE50Zs/JK8v8EneCrS+j+n1qxQ2VKf7+vb2y
N2JWdeTG7f+HWwfO1sr1CXz9QtwaRMnOuO2aBit6Ai/Gohn9XwxbWO7I/gfbHS/7
RFbrY3RGiabH/1L/sxOiNQhC+kyVEzqavbkCgEAWltrp1dCeSYC/Q6ldq+od8iqU
MakxqOuqroZ4rGSgqpaZym5suGpJyd1+7H+MkSS0QR+1FYhfo7+SwFCyXYkTCNmM
HRqbSCKB0nBgeXnC9YFuT04xq7//+s4QVnbA86IaCbfIfLlX3Qgm6lquTZeidA6r
x56yMFVOOcvxDAIu6+jM3OHly4ffLRlGVaWht0LFA3PBDa6S8cNgUL3DsOMqVAsJ
6Yxx2vZaBRwyOXgvgShSqtU1Sj5q0MQO+TADnPr7ICQUWAW9GB2TsdajCBq+Ok2n
EvpDM8daW7T+76+NLD3namWfa9GhoViSUzxsDSORL2+V2BfA0/Eoi6vZJqipSn8P
QVu5X8mxQU1bVCakjIG4xkQsKFg8l16RolEQ5PgkXMPsEcimbo7XytfyBGnuQouQ
cXgU3g1NzVQULQKg7zYEd3T5aEeKyFd4f/gOQ8j2heGCvTWd4URfvB9rkfVbWUxA
52u5Q+Qj7oiCQiWf9cHOZvLdsyO9dnGsRcWTT43Q/sQDzRtorQdyIpitKvUKUupv
jZfRd5caiD0cofk+b9lZQzKuvz4fh7z2T40ptaswYtgcK52LbHnxvH19add73td8
4zKMy7pTESh44Ycy3UCSALhEzL8uhPoji0EToO67O014y4yQVr5s4Ij5dEnORMhA
ec7riWJuVyGyEWbx7NALbZSu+EppIZ3IUmccwHZRVLTyHuio29TEiC4szhdBpmZo
uPyjZKqS7CKUDB/PZ/jtCXT3MkOrWy2b9b5Re3ld8KXrZzqClmzuuamEaySn4MNW
WJMA0HiZe7y4hwcX6FopDqYI2goshdmIm7hnJdfVoJK2GEyv+pBYY03bQLoMJpus
3YvIqN52pErGdqUsYuucNO0O0jQFJqelhmXCg/+kD3q+7/mEqDNABXAdXSOdDDmj
Mc9+I70d7/SKMODrdlKX4xYWw2zFKMfqw7yf1kg9YJuon6bIGVjGi8jbEbqKW5yX
qoUwbR/MdyHSknxA8sYgSR2zl3MRhmr/1QJB3h8zcTI2HIS8l3rAP3z9hhjl4A+o
VDFxzPWv/tJKyJWmuoaNGHhIswuQJAnQ5Ev0AQwHEB/aIKYo/qYjYutLTL4lR5xr
aC8QWx6mHHO0aTJn3/8BL/g5XrUqLTlC7OlfNWEin6Sfsi9dQXkjTRi7n9KWBgo3
qxleejqokZnZgfESjxrLmwtSs9VhoCKOfpRmkZzdE0T2LZOB62t91HnelLOqsXZm
OxTHRSrl6WlB5jV/wGRNj//9UCn5heQMYgQGLut6njRbUR7aPM0U4tdzEFkd8hfu
ks4FrPoG6i/nEhQHfo5mwgZvN7qBGBCCPi81DwpN8oF9oos3yvcMt9EaFMMoTdQk
caXeLg2UcY6Q4kvHnW3CCOdBFRC9nK4lgppPlBGFhXYJufj4fMT5OlzZm2MKK6BQ
8h2pCzkceEE0PGVmOyYNWzQc/T6j800k5XBMUtBg4L9xjSZTDOQbPcZRibnbuhhs
zUVhWhh7QwCbAGgfwucRrb9S8V1Bo47Sm8BR9tznlWIJMDXVBX6GYGPccOsFlGND
GeOwMVWV4F1Ay4gRWlAv+5SrulF4WASNgk048TRxn3JmQILNQ8P9+jDBm/IphIfS
jU5W8TYVDV5WZVoQsWrkgqcygwEAeDWu73CPFkNVch3sRioFavKcITeJg0NJ+ncV
cyQ4tHqUdTjm+69CSgj4Bp/ohw1StIphmVAsnQ4eqQ/exPDo2be38y9Ln2Hpf8s7
9ncj8KXFP7xMoWzNL16zRNpr70Lqxs4VCWbk1hO9JABZesz2+NPzklNmQHixEY9B
lfo49EDMKIY3jh0dweM9v94gPOxXetbekSpDrj2AiZ+TKcxMTwqz9tUpmCulyA4k
efIrB7tVoucRoPbhTNQyJEVXoDWgph65SwYIiHyL2NJx0wIHG8/w9111Gv7zKZtV
OmrMivZ4I0kwxSBtYALAl16pKg8rVpNP1bTqrfEC5sBLMn66PmFh08UXZIcF3SOT
ov0nXG2yuht22Df2y48cYfx4++H9K6I4XHcdcc3TBIgRL/0cHTwMwPaIj+e1yoOR
9L7srzcjJQaHHhQwBowyfa8dZ+9cBZbev1Jebm/GgvePQADr3e1zr1JYUjwyY8zG
FXptSW4j2/+3gWB2PuofOI4+XYkFFrrU54EsTsjfR3pz5vKNUOql7Q67tEJMU0J6
s/dHwqxkAnXEtL67WkjUPGlMuTNOiqIiEQ75Erg55MjFQtwuIKK82WE61cuFHMPV
tbptXDuCuHulGJGLtpTuM10m1TteSOVgAe/QUCRWrQDnHKtp1UFm4TpMA2bct67G
jLQ5JXkzD7lHbLAZNDfXQ29eB9N0+dRjDTyARldJYiP4zo89yhkprzxgxPQErrq9
s2n5WjoJ7tJN1aGPdlHJwVLIHsLoW+Fa0Tzl+KrIh2NvfbV0+IqQsX34kYs7FWYt
1jolQPGKCNrX/jADnqedXIO40s8NhsvgnVgMOPKr9mdGPeF6sBa+XDZgpwUJJ3J9
1ysiwYCc6f+WN5PB+9RY6KFHJJeiUcWJwqGXnTsChMeLN+EdEKI0bhQVuxTj8uXI
AZNddRSQL26VmzQWPxRIKgnn6c2H/+hQ3KxO+Of/q/TpSY/7JImVv2CmC6ptsGuS
2D/8XuLs5M+k6C+TjRLVrVvqhwaSyrY1QVETx9UMml7y/gHmmMgDN2crpVjTwHeS
W9p4cXkcY+K7Di4BMVVId5d5kAMzCgQpjr4fWSsKbkPHb6uC1Wq0XL8nt9oLoHTq
AVICRZWX7m+TLSl267QCmEVNiEJbztmS70PPFp465AKa5licsxxlFhBFC1UCUOmy
XFAKgVhT7MDlzoi5XRUV+pEX+mF90Ea8YHqbzHIkIrNsiG0SxWPmWg+j7NrZOT7+
RURmqXma6opVt+IeW8YwFk1jdAscct+yaz5IEdc0sBHlYf0wb61tmOrl2XiTBgaV
+YqtJulHmmCkN5qshWLEwBTvMwHZPeAIr11Fbq3AjerXZox6ZSCHL8ZEM+lR81n3
we5BbrOmpBQ8ZcWe8NjQCkeU6x3OoHVUL6hZEfvWj/AqbOxuHmNqHB3aXyUyIlYm
uOETvdGy5sV+Lrs9Kzv2G6hDlctoe9gUJ+3mrk1vk/diOlHCEZRPGKx4XGz10KSM
FDL+IFa7HBnyPT4p1a9wfbuSynBsMSgQ5HZvmOFRlLyabuAxMPlW2ndaUKH6Vs9b
9rT2cDg6srMOqx2BeRFAN7QzDk23OvpS80ZmZ6yJJmVuFlfvgr46/53fRfVnj4gz
jUD5GijIC+h+UWbojWC/LOXjApDC/bv2GTk5Izu5Q6FE0M7/UXHIO1hY6qC//r7i
W+Jy4ed5rgp3cdjsGthhO9uHv2QQxmKmJkepRyJ7aPt7f7sJOSJ/ZX9dNUbd4OgD
FxmV+xuB+6XVoMXA8uBXfx7BOj1Q1J94zmSPj98di2WJ06khBXVKDxssFCZeHswg
2Orn8JWN+J+dg0sbS3uXRcnPHq6dwS6NaMf/3pWiUazQt5W7mQVr5x8+257eZHKO
6BGN2nO6+jUTr8anQVtMK1+F7b71H53Jrvh3JNhHR8pRuSX59rk9EK9ifv8/je4r
Tv8fEKYSkNaU6IqvuAwegTKq7jgfxfzUbAvB2THcU8Gb3UVTZ8Qk/EwNVi4IYnky
/HZ8qJBZfaNMVkGB4NN9lc0FHejgAkXXl/9pU2AhKp/DP/GzH7SIxkjLEp0ho/Ew
Imn9t1ya6idpShG2eaaD9sfBna0F82q++aO3DFRohzkAZn48v0P2QDPZOAZgdbjl
AXbsN0PEI54XokVgBG2x0F3NC8ixWUXjRmke9G/YFnrp7BHCp8wQWc6NNFMUwPE+
Iwv+8d29WUEaow0i3TZCW2p3nl02mBNVFgzZHqRqGW+qzAwJuChdERhrRqj2sCOm
2QCiLdBOXBbSNaACq21ybGeDbnw5wo/KeRmCTJLk11NgJbGUWD6/E+7PriH3CBAL
fFnumMrOJLOh2coousoqI5s1TebufrnZgejByOldl1WdBfD85om3AUB2ChYk8fFv
C4S/qDlSE6S5cXk57Aoutg6/LLt6H8iYTtWSeboipBzjFXbojBsi0N0KbxULHesv
RdKQjvpylGGHGDGm7Og1JAvAKM9l9vIdNAy2jIpsXIxhd/Le5aXi+5tMauLEIpvp
l3CP5Ibx4Wp4pfwuXyg+SooBR9WEg38ICFCh/r4CSdpQHpgvGsL7UvWu56UygJoK
gUwUvwltgNP9aIMyCiXpaHsnE5CVMLbv7h68/u+z/J/8AANdPON+EiGSxBPYqR8s
z2AHwf633eNd+ybAyMPaUUX0skFOf1P/WAbBtIPLvzIS/FxvIxurgJpthgStuG+h
4pAjRQ8/d2Dlf9EcsdwL+2i7MfXEVUOIS5Jv7B0K7vlpr+FNw71JTBjAjEInmQ4r
/qe4D/YoHcg8L81Kork59q844TnjqrFJUwZvoEIZFosTWhBnywV2aAKlv0JeJViw
KLLS1vD1PesgIioZ6FHqAF+mtAlCbnQdHTncIxe4i7bW+oBZmuPHqV4hVlELLLbv
TJdk7bUPADgraK9oHExQ+a9GbU4Dp3plt8q4vE9pO4RIfj/BvYYYqqeMv5OmrF5l
AoRt8eUnCTWATBjw36icrbs+krZTFWgMnogQgHQufU4XJhn+cqwEq/rGWhZek1hJ
tbBo9/EADyjQEi/xYt+oV8P8lQTk/vb6Zdng91O78YKv73Ooewt+/zn/qc6eLeNv
uYZRff2lStIaLvRzzQeN64sSFhWKMzLCj15jePGPMy+MRCmqH5e9BI2DPvuGbl43
+2K+PUTYfEIvZ6FE+NpPBYwQjQasO4vaMxLliZ10QLpQxt8U47aPaQwBRoUNFbOo
OGh7dpzMkRAQ2kpYAk9b/aNe0tI7P9deZ06/DGhfQQZSiJR1DchaOP5GnZ/7O4oB
6aH+zgoQVkN+2mYpfn1pIvCznbUOw2ssK4Yi3Q7N778l6HagekT0NvTbo1jrKw61
oMnQLRt3SXli92U/g6giawikLHGEOz0QpRpO3YkZhSffOuGzUYWA7ZfKu+9WJsHl
B0sRrADDdwGa1MYC5ayksUVCaWfBJRYCodn62OjvDqKXL4LPrm2g52wrk+i2juRV
yTxwrNbuji6TmBNo/xGddiRH8LULAXdtwS1kv3vB3K2aChywotQC+mpUIRCy23ux
LIaMAWD0nBoTY1OAizodpzfGnu8yMWnZDWVs7Mx0IS+3w8HgUHETCVUgEBvKDzbw
VSLIBo4Rlsf0czJCZmdTRuComvwUK1Ou1+m00jmgzQ+aDYGABLlWt4eH2Ejt7Jeu
4rRKvYFPk2WMv8fbJrNovUBzalEnSRUui4yNJiOBjFvTPThQ5lyXWHvx33lawsGL
B5wpAThPIZy9gLhPsaPElj0eBlKqGpJpG7LKJqamicE/BWFtnlZBs4hZd4TeKCTx
GS9oBJKkUVneuITOenlhvSRdGGDgVybG/0A+knSl66K8XaejfzLeaomgxWpF4DZw
rN1wLc/KhPoas/jEKfTzETO6Jfb2U5WjocHh21k2NeNB9pPV/+r8Qe+/GVSlVyVO
vd0G2/ieg10sf4AmRm7huJCiOsIHMtlFmY4pgNS/WRnvMJpi5SPRbx8ujWLxfaO8
D+K+bqjvf57VRvQPx3NOlkyccOvmL4Xu+D3mgX1AxUHSbJbN5NbSTrrcVa+KfPre
87RKDLDUrpDOSAC2zo1F0Oq0PCpzEYw1RO2u5FAnpo2aOQ6jq9ZeHNa0raXRzAL8
XoyeNJwGH5df9qRndkj9eg5S4oyA/NWlk30jKMjigYcjIZdcguwTgqL2/6E5gYm5
diNdvUw1zg/WT3S6JgI10CJ5XBdEe+tbJu9HVQlBB9OHTxR0mOZr1IBFPdBvp7sD
zJnjPikktCS5MBziUXCxtV7Ts7AoJmfslSs//Hjf+o2uIGYU0OuRi8PCVIdlOd6O
nE7qQebbgbYN/hLJGvUno/mU/yz9FNtOUUwMS9V/sK/FuGXu6zN7RTve2HXQnsAa
R00VTAV7Vz3ed/+XLniCj00FbzBAq2pFeFgpefNWDGAoI82eM8nP7FLd4IPvQA/e
AE4ZigyHTmNiPgd1IKxJqZ6K8A/0XWIley1IfPLc+dO3cqNENRuRCslvT1zsR9d9
8x/1xWN4b/CgkwOVYWn6nhfXx50HABanH7s4j225Zs+x5YduLOSlg0pp1nlta0UV
bzrYgajZra+QMZ6HHrW8b5t4MY5U6/a1+36Wr2SBLxHXmXFjJx/JF92bHLG3eXU/
qTXghY95283c94vr3/e0kwVifHJed3Yb6sQtbb9vs+QtVv7tcNH2KmJtAg/lmyhP
duqEoCXuDfg3igFFoDSsKdbz9c31kJ/7kaF2bJUK4kf4/9TJtTNJGy5KeVy4A1ve
1mWntL2BIjtbIw0xyyqjCV9QnEh2395+lXa5hZ6A1hC29MlEZtweP/wcqRhCP+Xd
9g2qptoiAi1yBvu2I/fzLwTwHMEJy+QEBfLyaxikCW59DpZw8xzDXhK9ojTPmtYY
/GmCEXjsdhzAvkReMfBzPMn3mFMHkI7LLOchdDiqGQ1Xk8WqxNfkJPGsTqbgneQk
Ai4BmLiS6jSM5Wv/BUDbTUJuQ/ujF8V1aJnQypmiW9cwNBbjkTY3xtuQTNnjqJWb
Mkk5LpBqmNCadyXPDCh5FeoqAsUbrvmso8ltjkeW1PqX1Ad0FpaHQLdyThGO/961
FU7IrrF24YGgNPtUh+yLGxfuTMd8NvQ+ceqHeX4nlKSaHSyBdRImYBglp/WjBu4L
Ty2JJ6EQURooWTthpScIAdQ8TE6fZbMFrMOrT7gLQpoAaOMcbFBQiT3eP2Ilrf9X
5/f0B2jRfybdyt4pCoYNcEDcsLd1re7nUBjtzAzjd9x3/9Mi0UIYV4nJZSCtt9aM
FCdsXLMJQVrujC77W9wvrsECki1q+h3iKQkITggWQjxI0hM8j8tmlMu6BNF/4Io/
duubyW4StXYnAAn5eBpqEjyqfTCPmrjidlLuEp3vQkrVrVJBklTY1iFTmO8hY6Dj
q+65HZJA702RhuaiN3JAqspzS5QQi77GBFbqc/ZImxk3YC3WR/xAOOUFsmkNlIiA
5jxGyZDBjg6ySm3JMS+u0gbUg8jZA4wviqFMCKXDoj12TEpJoHZNpAfpWBfvW7qK
aSZem/HSIYANJ/heuIHsw7g/Qf0F2gdkfzmV1EGw1eLLI5hxxAFTsZWyKi2VPjzS
cCNkZQkEg1XMYMAfSRpdIIwCvveT4Q+2PdGilKUN5q47dMPISxNnpg2rvjrfFMcA
KvbbwPl/JFFIqwq8Bc+kXDiOAw+6JFsTbHesQbUWHvxXOMPwSHaYHGglDlTfjQOY
XQuQsrxaiVK8Uaft+SFbhR23C7DQ+b3EW60YSKXnCz+AZRr0ClzOElp2c7qWg0q5
Iol6HG14zpjcpj8OAbLL8vPvRTwEyFEZ7Qz0fHAdAFXjredHyWxwPsSYFMuTbdqB
u9hiojhDbMR9xb+NrR297cWFPuo69fXe0oIl5En9wXlgFp/3LN/rlBOYj1X1qRUu
rBlgh+UzW+fZfg8Co1Oczs2UW8bYBqZCyjr7wzyIp0ihDKI4ltEsllBrhrpsGbXy
CuZ43VrLW93/7BuD7I+8anbgD7EnQ8MfvKALEmyUL6q4SBotErE7sZYhdUo0bpoK
VXA4YOnhkPqKU4T++XMpwDDwkfxCPNSe2vw2rB/xJn15UvbtMRgHBzxue0GfzcG1
cvjPdJ51F2KwkS53di2uIMJBq/gmWyH1S4ZNOJGSkas5ZSAcTI5pEbM62yah29Sk
zGP/smXsxEb7WRxXEn520lm1lake5pE+GqGDpq5Ju31A0TPBvDrI47FDFBGHYGGi
2gtGjda3ORjzopPPlG72qF3MGG+jrEAR6wQWaKcPLYg4Xn/OghO2EI5pSUmgkKVh
eNj+pfMSYA3tc8HbwMR4syt5YHZU3OCV+K1JTWq0+kxZmr9aJGz0bLaOcwiSmqWH
CaN3uMsxZUvEiUaWTlFgWnku/yAQZlYdoSBO6PHG/usbRcR9TxbHB327EzfYO/sZ
tKmDWmWZYpQVZhHzQJkT+3CX662zJGOXa8VMFpGjMUeBEwRaw0OtFfhp5uQlL0hr
WF0huXpUThHXASDz0qi4vjVu6Wf8+VKC8n09pwHpgR9s8ts9cMbf2IkayLZ0TfWz
ruiykVP5ktPW95Irt1NmwirSgtCHIENZIDZbKu9ZYgq4gYpG0hM2JzhqfayNIXgb
sIKRTcj9UBWhidozkDlIRcBy4JkiUhB96wTaA4wmOZL+pJeJtzpGLpcB5ckVoeDw
XG5zAurxN4mYsEm2maTWbD/rNULuPHlc0kZGRNMuyyTGwCEakAwxVDbp5GivuyBF
qGpTFlzg/zMf7nPZEnv7DrO6AF27GgIwLXqJ/KrFfhJLzvHuAmgJrnfUfTtr+CXw
0dyDq5BWjvgfh0uvHBiNkuiLSfVqC/sgVAIlTULMMZq2vydFFsoVRWp0HChGSn/l
GrtO1cLk1SuaJRQ9JS9OxX1gf02VNaYwNbUBWMe9PbgS21lNP6EdhV8Jenp4SaOl
q6HryqhPOgJV8iyVRQm9sbP1zUlypjn5NlECQQPYZSNf2kJmCWvy9e6ksnfX8Nm5
fDkFmy4zOv2FQ0uDnGaAws/tnxkw44uf1Rr/oewW24vDcbkaUISyifVQ6x++OCr1
g77cIKKG3a+QjWl+JQDXiLBX9zucuIsDfAj13aCCBOm8EKF4OHo3fV30hU1V3seL
ViZl3k35MaiMJP8Ijj72XAW0HhxparQHEVyfWaJ+8AIFwznwN6TFZKjaTStOC9fZ
j9vocTydcAcLLa1KomArJjAbtIz0APLWSZpuR8oKp3uZ7d+mGHnQeTjL1u61MKUu
MpGyOpg+vofiPtZoEmcC4Y5Oal2M51EAoNUadQk+QCInk7P8yo0nYSXjr6ahz8K2
bufBO3CAUgKPRCoaRnmRItm5eDgcMdrE46q+2f8X3r3gA2vDLqvu+u/HodNjFDgL
a2cAK4uGyer2GBhvk7e28qQtKAOQOfCzDnbXr//X+My9Pzn6/fACPgKBPIbkZ99d
bQt7w5X/bWgvpCwjjZdxXoasXpzMK7WayiKwxQcLbjQRVSpU5CUsj0w1X7BJVsCK
TagvbwIVBghv4dJgQ8JV67BkMIoLDbTfkfuKoY5NbceqzcWfz7sMS+AVWbvKFJUu
8agclMigb1fZoEClOeFS9F5zfz60TCCSrnQGzAENxAvm5/k5i0X2jkQhtQFKZ2N+
RB3to6Jvege7qriyaYOG4aqDPJIetOFWIkcwKR4+tKAbGYZUaG6/VKBWIygMzJ98
0BBfklBxP92Y4pz2jJ4Y0tL1CIuafOfuKM1fXhHioIT1Wj7poid2W7FGs+jme/dx
VJ8s6jW4csmkRll1+xQhot29JRPNGY0wztHxfdfpvK4s3tcs99f08Jm/RA8FxD49
CL2ZoAJekuGpZrfc9aMCcM6+bFhXJ/lDYuqYp+XmkTa36sbOier483Uj/5ySYA9d
mx273THlOYzME1TLy1S1nGGGzmj2f4oXSifqs1ZKg8p3bHOcTx/HWHpismD9f/Ms
tUppzFB8XgcpoFhnEoMXmaPOQ0XsMO6bM0Xvr/nljZVdP+IMCQDmhXky/DZgVf14
DYu0zjrO1XofMkcLDUgGeZDeB3WyyOEmHKxziKwO8giWleg288sHF1VamuuP6bkI
7WzaBUlJeoUPgvSalFD/omxWhzqJMuxfYKPs+oFtCAJS7g3G86+8hEzi0e9E8Lh9
zk7dy1lN81iG709DUc4fs2DAzHrFnfFtz9QOcmlLv0NmpGKEWIt9crdDM7N4MInI
PttolDYLlrKk+nlfVZQSvwyQ4KZvUtpZ8wGt7r0/4dMlOg151z6sMDCU53x9l0Ny
Nt3Zf0iJ6Wo0zhyCOoE2n5Vjxf839G1Xq9xq9GZpIaGTyVJJTmoKFSMElCRjlbX1
M1yPu3vL/3ER8HzniOY5gtD253rOMr1MHsuRuOVpOlgAr3G1gG+2sybjG2/OblS2
MccUI+lop18d1tN1PYUqwoYqmmuC0Js6f52yPdsFoditNH+abJ/eSWT0A1h5HpeO
zGP9Vn5S3IsCj74OJerD0qLXnFkKG2ugrQWMBGkm2NdgbKpRlOWm/AZpeiY5qnyB
2jyqcWg4QL4J+QQtbHP2PR6M0WKRKlKPzlrwoO6TrkeruzRI5dTdMJ2JH29f2ClO
OKkaRtF+liDRWhwrSDUpHFZZ5xgELpCzcFRFdCd5YhzJzm8bMaUaVgleZrxjkqIr
eZDIhurlg/XVqpLJHLvYPme+/th+ya88V7gvV4+wqnaXkZJRC2tvlXpbSf+G92Xo
JBjXjXi5/CLogwy5iGCWVMMPz2I44l2eFWE5f44TZua7Smj3A7leUh0/y8ypH84l
cid/5VwJED4QdrxKIikHfo9o0NePXNmaoo4VsPi42ZAN4S4M9l7oow/JS7Rc1NM9
iE0/XMTfjyu4KwsS/OZ3His5aEfSQucruJ7vEpjaM78KbYDyffc4bkKKxHq/fanD
xVzY/HGqxJ4PYH3ak6j1nQlQz9omMX+EIr8o2bpo5LoHOM4W1gw6q+yNTUlIT5KD
jImhPN6wIAwRNyzZg4Ml1p1C/rl5qoef6e3YSofG8fS5eNtGigKu96H6i1Pe/o8Y
IFNyewLcchKr9FBjFIgmjZgxeZiv6hLPAKJDS3t8s+U2dPytDTOd5SNKchM824zY
e3tf0YNJNfF7CsTvmddJ4KGdCmSkvCFoHZ47/HTCW2V6g+OTgMVgXsDYxz6Gnne2
0oHxQf7A5g2o0TgP0Hq1kRBjU+dHBDqQ5+j37LXCb/Cm9dmUadAgwJqCACtQ1+4o
qL4Z1WSq1L+K6ftAu7p38DP1kIK9RSJjIrnrPuFNw6CD8t6uuX4TIKObvZ+Hlv17
dD7Z2i67JmJiF+/tK3tD7mqPRXAaYHbBsBCP/SZj02lFZeMae5Otk5v02A4v+LXs
t9vcDbRCWLs4hGkfHPFf6du0BUitd7SLY7yT0xsX9Uje68YHPGwPZodfA/QeJtn5
OoffldeIKA1JVxo0VIZ1s70OUZ97eWsvutGQteHTzfL517RzQOOKhKLXzVc50jqs
BQtScx7n//BGqbEwM0L7/GD57KY2FjWlEA4Zjdwy0SUulTyBlBZcyGVuNMBHqKas
S5ysV6sBtIdzgj3uBaq15nW+ny/mVSlwVRzfbzCcOCJS5u23qE83p+c6MfzogWNu
0KYVwLhn7cy40KW/VJZthLDNk0KvkSr/iEF2ILNlNStpufwdYFsKjn7ttCFAzU5a
XQBr5+IAPJJTFj01cKhwU2DVwy86torOAGXMkfZ6QrvOVIROLKLhLP0tUFQmCVut
9L0PiUX4Lf9Qxu60H3ix69fBdX+hcjYXCzZkyF7f68eU03J2ud1Bus57VKQiBJoO
bIHF790RlC5ABtxedqZ+tmOfVlXJlDnAG2covo2YE9XsKfDJaYDfmmgN+uO8nZsj
tMVRNYGThCzc9RZqvmaFjE5JQC6L2Fh33mlzHNPQuRQb53iTQbuBtCmkbWTCvDMs
t7ilH1ucFChexTc4tU7LvTJ9XxbuKtZmPACDkAO+k7LMBXNaxmm/9Pu380vclDSn
y4Wc2g/VIjMs7qY8f98YmzDMJ7MdrJFsRDuPjHj1csW0C5W2hwcFZggRi1N2ZytX
Ilhr91UAv4rgWn7Ddh9jc81I2kh3UcMsCfpBfOKnnJ8YupBz3Vw9c4aeyORRn/0M
QkpiMn+apAtLVdmOdPH/4yOxoPkcxpnFIVhlAngD2Kp+3sMxTJoZMDcNAdD/CwdO
X7UJIkRks6/qBfT3T+7HqCWJBg73Ak9B+B3Hn6aLcYJJNTYpeIULXXEhITUrOYPD
Qr9Fzqj+97c6ZGlxhvXLHHdiXVwOb0677x+kLCY3+d8QgfDFL89kbOoW6hceVTc1
mY5VWVRdMbM5u0KgimKlKonZe6moURcmE3RbvJzDRv0mJnwDtCyNxAdXQBb5Lgmi
WUJmcv2YS5gfOzup0Z3yuUXjFIjDDo1RoO10HMbVmnCswTsjhg+mHOTtr4oxmg5Q
Wxu7QJFxsQnvyIX5tN3y+yazypjjcs1kGGa4FT9Y4YoFxSPS1GC/SUZMfXANVJit
zFy0aKNcJILAEK9RHjuLcXESePEi4PvP9DU44LQWEY5vS7Vqn+zT9PACS1Qcqi/n
YGsPjLx8eLC2nbDEQZ2zXfsI5nap2Y0n2JrFpNm3Zhnn28kQkb8/nUltXzZ8ixko
gutW7omiRHrF+Q/ZHkRby/5ZF19t/jCdgBQkboc5fJBtCYc/+uTD70IWAUT6HKFo
guwVyMfmzxbS8nepFS7oOaGPw3WGa7S8Mm/iunEWC26S7t6iwAD1p9w/CpNaUJEJ
2ycgyU6QQ1tVOu1tQCLJYyH7oe2n+meVi5xixmxzV1E1aFUIqMnA7KdGbqX4rg7t
oHsM/wwWGp1NTu9LIa7oOltbOO1QbEUoffNVLykEe521oFjzPQbHJ/6QwBhgwhBu
Cr5CR5nm2e9zj70PcXHPd5vvzEl63ZsSvvUfoieCDYYPqUIdvxRYaeBL7CKIphqV
KABdtPVg/YuOKYCBzf2JuMu+oHIxA0ecfxREpZ+E73UR33ls2OuTOTBnHxDcpkU9
ISMzw1WY94wQYo3d4miqvmI3dqYZirQ2Abb5YUfgqyUQMEz3LKxBdiobji7oMjSr
TrjOHnCFLWruNSlhqOdZMn8165z4En/D59HIpIP1lGXT0xKM0QVwOyAHWF8Kds8C
rmupvQfHTdRcTTZiLWO4kyctfsOlxqcelifY5+LvuApof4p0W6PMUOpyg2f3fmNN
Oe0yFYiGxGhyezWdMrC9OjT8i5SKi+p0K/40wYQo2WbJTCXkMaVOXX4xSxjhFlom
Pp42E4Ve0ZJbEiWmQ0ey65ryFFOwMchixaQfqm4qAEOmKykG29F7Xa9aA3WQn6D5
Uwhxuq4cYH10S5Ewx0YDMtUTU8s1VyuNJc4bS11K9TWyowmJ3+Sa57YMyYzqNkIc
Z9LE3dbkq53nfy5SXp+wSphlFg0XPRdQ9i+GZX62Z/RDm3TsL5n2iL86+pGGnW/F
XYLUCQVpT0jJxj38v1c53ZQTh6kdvz2gOfEqg4z1EzI7JZ5PxQXYRT6YsbgY9n+r
rDDP2kQT7X4uCahP1zQC7zE15nR1/ComNw2Y4ZwP2TPzEecy4J5ZznWbwPFYLAQs
ajEYsQaZtR5bdbHRXGDTyeplt47wbenrk4wF+pppghmNLEC9cXlrv85nv9IBgXnF
k1A5brrqOskgK0DrqNBplDMz/4o9IbUeInofQnsUjsG+worn7fOSo+xmeRwadW2x
kkM9wY17wpYSNUGfPYLBPGyb3sPvSvDmkQNhd7R9KXKdCDOa+t7wD77GfkjIDx6+
s4Y/dquGU8lwm1Ofu2UpO8rkOIe/kzrYHi5Oc+x6UtkuN+UEbkqa/KtfW6P086Ej
yVwe7q48a4krHWqaRPg0VEbcwSVG66ez5TqIK0ehYxABS4Dma9FOSRhjCEzq5tme
avYGbXkhxw1nKkzYJkS7ccW4q6sayytcVjiF4KmuqtLaCPrBwTfKMorTTmXKxjFa
8fGCfEjZqXNcYH5PiP1mSdGdamjeT7H5i1C2/ERRxnEsKLqenuXNkn0ktzwpPZKz
y2UCevj8wAYb3mkd4inejr8tbSeTIs9xBk+MuJ1Gg2gjofHWgI8nQlM1XvaCiApS
UzqXETrZTAXjbpmcc9uIF4SHNbhqq4Cs+80axTlNOZZYSEpVGgC/Qr2sGB4QtPaz
81FX47IryHfBz7qTbfRQVlaW7d+n13ps/jcWrmTwwCZkIDhsUzHd5PpNpNu92w6g
yFiyxO30HGuH/UyCvUcnnk1jsKJCb/BVeVmJiDyqtZ3KQEx70RIEJXrh8IjW4qgq
HKgfbkjSsbs4OzAGpLKF3eeHjApVs40XL3haaMBFpMQIFmBexv1QWA74cYv73q+a
mb7dokaqT2ZMx1DVXsNEQ93kSoQ5J2c6Gz7nWwWZuWm6YjyUkmmRJGwU+H6mKX8A
1xkJtybNgba5/NU/ycwx4wS58FRCZg0vhnoPu3t2onuSCeniL8/qecqqWVpUKBtf
fZZTN6m+yIYuMTDriG8uSX3FUAWy8QRYlaCwTiBWn6BaCPy8VPSnAoBjfRePw9II
igDOnO0KttMnSHRoSCnZEfc8WxK3x+Bw8vcbRRfWK9YLri5rbG//xOrBZDT3gw8V
QRhr/GhuDBbZg5bkmtX1JWlE/978JoamjsDhl7tH4k+ihJagrHHeEnXfDR1gbxAI
EwugRiiGPEIbOJDt2/LB4VLjYancUwa2CtUdN4gvtQ9WDsBlHOb3fKoOQTlN9lp/
E9xxw89c3LA06wMyARSHPiBj6ciAMVKsqC9z5mI7QbLRd+of2JRy3uAIZSNNslnd
gGUXCIRTnVtybzL7GTXbd2beGEqRaEuLTC1CDdSzEFFCiVxwtxPF35GEvHNGYGkC
PE7vEr1JldSuSm+odd8GIBVTyJ9HYu6pLTEb9JouMStyvneYbDQocz284WiG8ugk
Dyqqgyn+4zYGPZh0EQITfwtiSglZ/c1gf8UhZBsAu71FK+iKL2A9g1Vv0ruwsHNs
ZI5D5V4OBY4HPSPkIQt0xRUeu7Z4JkXYDsMlXWAknG7rDJ7muPqTV4JfaB2QDzv6
KUm3F+7dviLwYpnly86sFBujjU72LQIMwxuT67yDZ8rSCMvWdN7ljEPgGlh9KOts
MNJgatDxp3Ubz/k0TVniYjoIHBgO3jkMOPkndyxJ77O4E753va3hgNzn7/70eM60
6h0C3k1LywaXo+BR15SUzpms1TgaetNuRClpHAN0JNy8pocTbk5fjLI0wyv6F5K/
ZlKUlzcAlvXbw6WkUp3jr1XS9krirXVSRq4J8yp8QG0i9wf0SBCZ2YROVnewdU30
0kR+Fn6gLde5a9weKeIaNOSmNFPzQXZHAY0i8TFA1miIlvmUpKQ3aK1lVroiYCka
JJRdjDlivZ7mC2ulo1HZ7ZJYg7nfpae43UX9RDLEklIuBa+QxRwSOu+DGlU/qIp3
ei+5F3XDU7H2Q19OXfcUaH+PgivXmDzEiH8URQ2b56nN3v2soTYzZWGSSUzPH3fj
fZJAaSnyjnZzoCqPwheALgLnhFqntIPqkV/iqaFpiLtx7EYnA55ObjhJ4S92EQf1
UzIc2ELgqpRSA1poc2fqJgXhc3YTne1JPtmT994Lt7s4oqJkbsqCVVOlkja6xYWw
R4Mq2RrONYuqat779mbsu1B7RQz8fLx+OpOlIklbDltYiNNbQetWKHyEOes9MXbY
QOuJjgcLANXlXiKtFRzsi8lOUFGfXZJ4qJ6EjG7aAslv1pBPQSzDOXtMOB1lVjIZ
Q0YpMvPAVBIH+zfdL6E4NrehD0gKt2b/HrocRajDy+sW1ZEhQqJSiMeq+Fai717h
k/v949M+lKgxtg12lGG8uzbYNTfpBK+fbLXW6lLbWx9VV926oio5jlqzIdHxBcmw
iwYY0dGLJEPednUU7lU8qYL3F6Gr2k8rYVG/DzN/My7zClMRNcDZDU2+X5SesBsz
M3jNRih28db3PhS3i8+f7xtcTSvTt36MjCAk309snty0/nXWPju/aFsCjNOULOnw
zEiIPPh51y/2wVFzZiFHHHGvP+KRy2SLFtR3acGxmFNmRdwZo1XA/16vv0C7DwWB
Qn3oih5PQlWIkwaO90as0CI8NlnX5h0iS5YrJm+O4bfir0BCUJjEgvkZMFng2k4X
Efo6DtnoH9Xahg9VrEy0qVpEyvjNmCjA+nBsVUEx6Y5+zzVxXzDQqhC31J0KcdeJ
7U13R6hVXdEHdS3XvSPoOfBf0RxjG5PD1+3L25lgJKDxYJr9jro5wMNq3toVhP6c
1hwxEJ8MHK3yD0/7LEjsz7RRRCRu5dEZbXQLTWG0ZStiKzMPRm2NYISG9zIGS3L6
xAwoEInmESDchxsDTXKpfWiqgKFlyhBxCxTFyUj7z7uHzjcLprCU42VTNkq4ufZB
dOxwq9M6OiCrKxu1zyCXOI7cbZa2ceV5XPcyvzpXjxppkn2/dhfqMX8lEr39INER
O1OxrL0ooA/4Bx0FhMo85ugcxhowrKbUw173gBDf/e8/cvYWBlnZLOHm9uXI41Sp
zoXpkoyJARmVwvp3uVrM9kmdsI02/M95CQsyp4Bv38pX9PtNwzjmf6XMS5Grgrch
iAw3/xMC2jZcoFjqNQ5AQDN8WbJDQ2XDqc4DaqbLztvcMdQjNjP5HUjHLRaulCml
neRRFVGCllCIxM6auPxJjSGPFSTRwUWMwM8BXSOovq6hYGJjIItTX2X0+hWgSpUn
XhAmKuwzl8EaBVLexll3mxfTAl3HG1zuaQGwl0z8OO1Rm1yvXm4yLlytYChhUUK9
CSgX4Ntvv/jJJ7VcU4OMQVpa8MLW0/eOT7BFguNOfJptImCURg622ZEecA+8+DUm
Vgz7CtZI+t7wW7JtLnRs0jHqy00qFHg4MoowTeb7BElAqk+eDAYDIiS64DPfRe8M
db3DgLE+kb15VVYz2Z66nX9lKTd8bR3nxsv8GFjRdPOCyheU2APXEAmntefcs5mj
iJxtfWd4rRDL5zWsHXcAPnMUSKeREjerpQCW9+5AAweAOzQCOIJuNu6Hbw+hTBtP
XPwTb9ZzHyHOFdajFn9ZN9nPbbKnChceuryK01O+Om4AyhpNlNjf9jNjqgkOd3GX
53wnfNAotOA9m40fJxbw2jt9XKv4g+TaS3D5QKlk0cfVCXhWEMcjh60931ZDKGF+
eQAWLGXmgvXTygC8+XNzP9iNSZjd08QsrQ56RjQhQTnKsd4IUzcfXMVqsWkdpGTh
5OcZa186j5zR5ljFM8I3FXZC6Gn39E0Oq/iCqoWGhi5GPrUQcVOUJkZRX0nVVtut
AJVoeI2dKU5p6AFJaZZ/3I/yLSf8DO4Nu4AsST4Ve8x3YsNqNYNafJVT6VRH/ijw
KLpKivlwHGLPHN7VUgvwf/+3gSc/al9bAal+Bc5HKvt0jpGXy5+9DUj7U8Zol5F3
pHiezrtNBb11ZZktomKZC8CBSP75MmGzDVQLkonpQ7/6PdEMS6RgNaM7E0zVWDEh
qWK/QVtbshKkvpIctPsPU4Ijc+tWyHTxcWFPcOCGaEeOXUOCJBwAQudlIkth+rCD
4H2Oi9DMn85lYwrSc01obbZVmWtFbi9DI7SC4d272JgdP4FmXRCIWEPbjj5klaLN
0NpmD7uhZwRB0G6IYAWJZ8wgPKU1SgtGGEbgqEKrP8BSDszgYIZRCOtzxOkwOsSZ
vTXY3eCgCTVfhO/VR/Glac36spl5oy+lrKzDL3poIzph9VsOdrgHPoRWzdD0u/Uv
cZYW6xoSq91y9LNqPq+812dub2xl9UkUrj/CztOHcNmOxfTc/5hNSS0uktGbkQIz
CcZqhvZMdA3tRA1wNFzZP5M58ganI7I9f1NbqnPUjX2n7rgkAZdCYbZS1AXEfMYi
jlS4QRCrW4lsczMKnJ1XDTD2hZQuEFVbB7R4gUg03EKrEO3/AVJNujmLIqM7/kXz
z1vRRZBFMkE/4HTQiR0gHrfuCz+hwaDTUjuBFmUY74viQhvdSxewUdzXXdJYnRrN
fdNS2avTqFVCDAY57UyArrJdRCFfQAlsj2MjcYKG7CIqEEEqtiGa46U0XRQLsn+T
ib7Gg3RzSmaKndKFa7ykK6LfA2g4p/ByYMZf1r66RRnaja7gjBQ5+8mcBTztnNUV
gs64z4BhUC2nQFE17jh97n+ftzjCfoSJyG28hmeZZQgzSA3lrK/s2jWjnIRAmsp5
u+Jb5XSdIyuZ8mrQrXsgP+lTN3uD3gSjf9DX+ZYTuLu/U/dtQeA+7vEHPnOmp9jK
QL7Qt9pamPOGflxEa4rfPMs+F/0vh88QMvMcAG/8XcXLSUG+fSoOgClS5WBHwbdA
fZoUdlsEsk26FyxwKOVS/0uzxwFW/AkXPubSozjLP9jwum4BuRogFL7x4p/HQwkz
S8DlZ/0i2kvjGhNDvZNP/X310arMBl1lVIMKEe6My3Gq2G8/92xuMr9UJJ2uUE1u
91UDRApoVk69dpqEzz9St45Xx4F3BSUPCwdz5/eOVFU7RAk3ZsoMzLX0hQIRUS/I
2hT04o/ftztXQTuKPZ2YtQ+Ez51fYIj2p808QQwM5ls4lsaMNSGFCIDAPVXehLFL
AsZDEc9jtQ2rrVttxYNP8sb5tS6yU+TTY+o4uhWpKCCoGL/5zgZAjudCO0JtQDpu
/X3CPRcDUzRyO0qg3McY+bwCA3bgnyi/Bn0gyqcN0co0WCI0NW6ENeFPRJD3bwto
DAtLbvKVaVWN0RZVPvWJMLU4xKauPIWEnjSvnJYioBSkvm2EQS3ZwuqZVAVVbiax
FWlOFfqKsdhC1AyoR0wduSG/XuDm1IcXclA288l4OtrSDs6+oW1/E/yQGJuv1W7X
1SCvsT5go6uZlUPfvzW7Ijl/s/1gGQWpP8YE74+XENUDb7cRuXzqDsWB3ZCPT5Wv
sj0be11kVOL0bWPc4ftXVTu5Wwiz3KYVWdatM79o8nmQIqlL8WqdhRtfW104B1br
ZUpZp5NNeXtCFpJDHVsNF7opzKfMxs+F+KevpT0qp/YpGAsJ7SVeveQGYD2ugWWe
uEB6c6j5Wzo2H+lZ83mkoGHWmeEIsa0qSkkMRRiO+C6t6HJaxpaZw/S8mhUtSbzp
BqaWFk4rrYVTIYgQgkX4hMyRhY+v5wGW+jcqABI5woDLLPeD0Oc3qmI02NFCVf2f
7eiTQqNHzJz9fnr2CN+JmW5sYtsQOh7lL8uSXzL0glEWKeBu3ZeRYeer0usheDdL
y/hjvVvs6lSffdDzZrNmZECtp2PCyTgk6ewclqZgc8/U1zGxAU3LftTjt6wvdDYz
sm1jpx8OrP+nK0O9z8KZ5T1FNfm8UvSZqTmkubZbf/OTyO07H+EGtDjuKqbGkERq
DfGGH2C4qwVsX9hWWfL+iVCiHJxaKDtmnpgX0TtPy6at0/XW1RE52Bez1YKZaNLa
tjYS1JF7rtshRrS/+LkZJnLZJbwH9ygVSl9/txzlRluiuu4z7ptqu7QF7DmmW5xZ
e70Cl3MBCD35pf/PU0rqLTcqwFVd2TAsKlWXe+VKDiRbs229Bym4kHRL9Zii6SmN
VS/mzuItD01rVKM6eSrEYym6J44WXAbTLnjVXsMuTOAG0ouuZ7er2sHahdi8zw5Q
NhAJy+TjRFkMCI0s+AMYovfeDLJlhtsSMA+c/AcZsP+ivz1UOTuMk86ceeGuXhNQ
2ERxyPJaeN5WPPgurKvKD+rtJqQltEULCqO3HSm+wxabYYKCk9K+4qtLrLz2X5Ru
6IR3C6rbcuNjVxffp7lDi4dqOWZ4+C/pD5Q/CUkN+N2R/lErOcWvsKF6pHBp+M/T
uOorwT2EUU2DpZQVeKIUV+HUmGDdJEgRk/BfzmY1hdxLaQEVFQKqgrRzeVfgDaSt
U6jK8S3OpbBYMYHWLACqTJGfQHQuG+WTBThsRF02Gu+XjFHyHTmz4W9RQ8r6cuqi
Y3TtVgwwxyzLV7toppLFCaAm9E9ZJHXX9YFQvE6fQEbXaFYdiR9aLd4Cbe6nHkkt
+d8bxqU6SYUd1aOCTo7pzRfhvENnheAHcYQlXdR19azn/i+zq6QnW8mVcEYBOkTF
6LgWMUHrnrmcHqriNJrn5lHETbS4OJfixqguOZHI++9iK3lkohUunKRAr7hPY0du
tGHVFJy3YH7x2Y/mwLlVjYJdwtkVyRrfkiGlNtchBKzc7xqcjRLX0lPzyP5ce0NB
6+JaLyCPdSDBDoIRQya7SV3DjZB4C4Pz5VfUUsnyER9ySrxODBsWIjlvwQZa08Zg
GpXy+ETvBDn5xlb1Oulijado/arDOohfZy1EzqrdGPJ6EUa9ZdLclSIF7GTX7TuC
lWfvldSpHTfHpIJcj/4aMOysbC1GpVE14Ic2AKbLPfLv5T81og1NPpHzX26ro3Zq
KoEc6TmilK3fr6Gi+ZICTJsVD2I27hEHTO8mQVXJp0y1X0zD5Eq0Hjcy0qORQLo8
mUxkyCTSWDo4QBeje88mcV+yjVT4awoHZA/iLhwAAe8PdaIpZ8fZYLV3akdMAzMi
wmHTbxTaEKpQdxBV96E7ni3aIb8q42fuzjDIpURyCIVBteMN51LE5QfCaiBRl8Hb
KBRHhi7iswLpDf5KcodbkSQT7zCE5VUesly8n++RO9rWFmi48XfE0WJ1m+MdesnO
TGlstbWC8/je6yKwke5qin6bJxRIlexrOTP+xKElRXSPQ3RtbE77M6mkKorQCizi
rewKAPB66Ike5Iw6snYewiMzeG1n58zcnFGBK1BcAV1jBVbzzvyAfYblCzLRTrcY
IJm8FjpjfcUbe7CKVwop+mzrv8CTatEmBhtYDhp2uxuEsHJAEwqErJu1XxAxDS5p
PxApdjpkUHCh5nTl0w5jSYNW1Iu525DwYzy0NjXbSSPWzD42UCU7hP3yJvzYoIFJ
l4jT6WmBWgAmpc9vLVsnoyNOSkdZKUcgxaUpNXk8W7Rbj+gIArThSMxyEyoRyoqJ
4IRQv7ZT7yYIeznuhVfqrdK+R6ldhcXx5u4dt71FuPOLvY05e0O0aWxOcqIIpyHy
OLuwUEUNyA2TpsgcYmgbch3/fNwTaYkdEasvQHZyzxFRp3ouz0dxQFDT0wkPHKZj
0fCdnjtZuQSwNr8SXe0X1PY8Rkg/9zAbG2/63ngraFBxnC2eog1FrqxW/Qs/+xik
1xs/lBunNH5LTzOxQny9hkuKy6232kEa4HlgufGyD8GV/JjLB4E1wqocJOxhdxrl
4AFZpgyYgu9kfyj79rHgMwOuuQkfWoTQ4aHJwFXLNLwG5q2oKdVuslmhYYkNez3L
35kJYSYWUcE0kIeD8Xge1ILsX1g778jWoRo7SrK/2LtMpjHwx+jM2X+Q6lZdwKwj
woalReFwewF3FYN6OCWRYUttDaAl7q0+84PYbWQCvVqqb8ty5B0LN8lIZJKyYt7+
p8cV5P5pLx7TlI58CAJgvDXRdGgiguqB/t2DMHDuS5VWef0aTvsL/ACTtZdZkpEm
qZaIxpg61lpJ8HWloyVtr0rKwNGCtrirI795SQADwf9+pQJZFxwM6976rc6FIu52
wy6vusiC7Cs+raSjccDv78WNxZDQNmQwo51ysiE/qyaeRSwXskXxmpOxJs7Z/Xe3
Uiuyq6L8wIdZFrpezbsjkQNLKPqHuKuQwfgfqN02+CxtCCKW7Wx/9ITsSmb35Pp3
cScrw5z7i7590Z2gFnIU2zkuTtQt7nCCwqQXxI5T2nM8HCXNXDO3mrmzG+HPwHjO
boWBh5PxazlETxMld8qkXVEvEYziTs+9a+yIEdklDZoSJKv+0bE4gwDnKYiGdSWn
4uy0HTD6hQcb2G76HTj3IAAr1LbbigSL8PQa2tMi+uKPG+PCqCObqvIVDGyURRRz
8vN9dbFSpa1haS11nbZ4w1GnBmiyS5uEY2Y/4VIj3ct78jWIlcCMszWz7w2+uIDG
6U/SD+kpZIOrvezheRozU5ZEZM59Rj1xhE2DYxPr45CcFx24qdCyXX34lXP5MSHg
BxTVSfLIzlv9MWlpFT67Vg8ZQ9coLEs1g+neTwAF2pGtmGe3xbpZpdiEXA55I21K
ZwRUf/6Tza7aub5aclCbaKTyhyuXO3oZSWi5aob2pEKFu5hSZpolL4Xm+LDlaVCB
/j6EeOkPrwxfPv4ahuxr9yU9Y7OHv3WFaxEY6xQculsmmmiBbyOYLW69rWsDSqPb
WCbsVhLHxD31wrSvf+kNeYicXIbYwMXluQfae9kJun/MPbRVcnHqFmOWhT6oU7Jo
9mVm5T+pdDbYOixrzoifVjVDzGtcntP7NeaeHm4fB09Z7Agg4UeudqiNAB+3H/Ai
S3HDF0mzi0HDHBE6v/dC+CdfwiUl2PTF2rWc185t+q2kre3lzjl4mff5dXbsWsDL
utuTIlNEDwGHNC6ZqoT9yNqu0+rpF3Riv/hdZEbu6BZ/LHWAlCYQT/6lvnItGtoo
yx+qxJytsYKWaAXM1Rf5F20Ocv/K8kNUkQUZGHKT2gtrblS8gaafJStRc++DDVD3
3o2DYzFVIc7RvqTxCUf7vly8qlcOpJjXUzIorU8ebsnQe2nlP+OOVCJ++GnASwhp
mwrHiSeWdsHwyonhVozzae5qPOWX0VipbVuMHHhEbkayVNHCISp/vAKk+ynZL3UZ
kNJ/xLKj5owx9LdmTITQlKDP99LcmoYk4hswP2SBQCxrqPLfl7fowixeUUQz2aQB
ekqxFfwtxwO6zVp0omZJsJWdqEDPQdffqmnWZ6Ld1MtEIGAKyjAxqn9ZSh1+jCuH
fynKjYChETvzTeu4jrUmvChp+/KhlO6rD218Gv6k/Z+3yh8575jztBvb7LyGmqrz
wZ08+d2KHysTCbimik01tlieyg5Yn95iH91HrJMELXigy/cWbSok2Wb3MoJ7Uwv4
rJY3og89s8rsL0wRwY7HQRlkmIUrXXG+2mDv7a3ZpdYxZBkrYH+pAgWnUcDhtfnz
RRIL5P1wvXDyB3/5HfErFzJjGwga0ruAOU3KSjcmniMv61RT/5LAEZGMSKXMMYFV
AElHp6lIGpFnYYiARsnCISc5cxJZyesrwsC0NS9sPdE1N2soTXDqqH69eA+ek/Rk
UlUCH/rbGZWwh66KCWLV0B8+ZY80waxyuXw3I6LH0id9sBxdHf/D13dToTEPHa62
SmkBN11gYKidblWzHjZrxUp/VsZJah85Ph6RNW+gI9aXHLo2pN6y0hG4la60J5Zm
fro/hfjKJvl/nnevJIns2/RwXkW0Mu6H9/3f0c//oL8uzf0+QHI96VG2JMW/KXhi
Nt5pI0v90m3Pn7oZbfb3fOZ5AahxILAms5fwuSv/9KUSodh3UzBitZOfKhaUjMV3
MGfyIMPq03p92lEbLAgc8nawHFR2b7S7AjtjxCjOpPoC77CBLDSxzp8RWbPeAP53
n+eF0lhLVpWxlPPln9CNhFmmlBrpcOR614GFoYVeGyUgA7eVX/634JXeTDldhg7L
A0xdfovti5gFIqw7JEIepQ2Lr0wncO3IWcJmy5fnf7lSXzFYqVtIWz2zbhpdDrCt
xruOx/z/7f3YOxJ1EXl8T1YHoSTBAUNi7571UledWcWBu6JHD3BCUMA+A+Y2yFCB
vusDX5cgPFfue/JMTS3QKVBljyyK1yYbrGwEWMTC3EgdMxOJMBjhySiWY4GNLFOy
T4C2itDYY24gmDAwHMmWMuOmHBltsID1/OfSssioP3LuU2Zzq1rek2c2Lt1CLwXb
MVtP/rgjKED3/6hPe8z0DD3ss3uyYP3Rc70N9jqA9hdRGSEeoRRZAlL9owgrQhxR
JvAd69jpOCKLV9CUNssyHievHQcNG7HBX3brtGDCzDdce+DBTM+EHJiUlcGsBlzx
cGcbyTwJtLC6xEyItOJf82DXJBFD+wEZC4imgtqaZOCv98jTfPJS91stBTEs9mPN
pkJ298+GN8QsB+t7LwjE6YXaiP9ndY3DJmSD38toPxsDGxx1nq4pb9x4zJgnKVz8
c/OwBn8AHDA2aPU8AF1rj/PDWa4Z5gtWBdbyUgaTr+HHv65FzCJzD8eJWv4XuJo6
rSiXlE3POOp3EhgQa6/rCPduuNYCcw5vt16bK8J58QPCHjjf79N5gxkoZQZ87ezh
wexjCt3f2bZq9nWkIyWVV2nAIpOS88rT/Q/fZrmFSs+0U6tc6UW4cN2CLxj8eerZ
837XOf9mUS/0C6Ob+JWNg22AqYKdkJ9W+pLVBYGjgRmQ3eiARpniYmDuGM/vQN4m
DU3qi67XzgHIlr/XDO/GpHPkFPVmiKzWIU7EjbhsvZlQaxyVgefhffsQ+oKZaWbT
rsEBp+X6DO2wIlARKZrDnYicyI2YkclP9Y3jpI7YwCemTgoYEnMRFYhpvZP/xUHd
ILNm0Uh2pdzgV5oN1keDMOBzBeQIXgXvu1rXjUC9E4kdmb1+FQosJUW3mPbi9ZrF
jvkq8RTGd+QPDzH5nCAAhGgqO4E9l+SSeaTRkWFRaVq/9mkUMTCEcZIiTRvvJXgJ
0d0IOOARM78bjIiK+cTBbIAQIzCyevGlU2IIwyz8xRIVrDR7XmHVIx1dZRseZKFe
j4PdUi4KHMvPDf+hhCTnT58X04LR6zoqfTYkBycPOQvLL4+gUUEWRyTW07uCDm+f
HWvhq8ynFpWEiw6t73LCGMee4JAWtKu5DelodAVc2AjcwLA3XA4F3WfPFaUOc2os
iWGme6qb79lI8xn/Xg9VrVB9qeUw8YndxjblDHyL3rZIxPeFscKtmRwFstGfGCQG
efMT3zOeefon/KRqSCI2As4Tvv02AK30ArJ0KI9CMlrKTUw0pFH3k3MtHehEu7VF
zfL3TduXr1p6Z9tzpP9qaoYnymNKfhKjXBy88vH7R1+jbwlUtE5OJOF73Rt+pkbU
oA7Ze2MbsNY4y77MQWOjJXRW4GK58UoeO06JDkJAP2sVBbSVFSEWnxCLH7NBtfRG
vygAYa5Ozy6Ojh4MVo9lZ7ajEjD2Imwv4Wq231e0q0B/c4pbuQhsiAkHYSvIQuAf
dTqFVhHn25dcwKriJuzwn7gxXCDxHj1iQv9CZT8RY7XpWPcmSaicJu73JWt9aPI2
JoBQ8UO793mKbIxTfRqGk9/J3cvWcv3elHONnWuvHHW589nNY41BdVis8TuFX2vX
WONfLvkaqfJIhD+0rKtTJPrAw/2iIf8Bl6Z/NcgitCBKBHmcq/uaICNpDRbPCE0u
cfy3DvqUf/b1AvTISs1kbFyJZql0+63xvqscdILAia6twwMFDKzgFMhjZZEmJfZv
hXKd6Mw8ctcEIbaEQVMfXo9AjG5MPtKDx3xOmu1BjdVMyb1KxNI47JgjPcIfm46f
E53M4so2mSgkFVc/h7i76rj3KVP3P5tZ/95oQS5CBDwzp4yg3Wrgizpzgm9I1LYD
H/ojtAP1x9y27xD/IqpJ8LYJZyf8voxz1QBGoIehkh91S56hN0/oLCgH1VBH6RSm
U0f5QaU2d0PHFcdO7N+I4NmfAS/D3eGdAiLvxoNqzUn+LTKrt02iU+hDNy+an8kc
E+OWFT/D4T3fwc7Qc68FQ6dKnSdeL3GnYedt7Z8opusylmtIb3puCWYSsze1u5qP
BiZ6cofc0GaRgCrXplq+aG2Y5g+ot/S2JkOZVpK7yQfMzHZKBswVe6JsOvvMu0/w
Rgu+DKLH4aKkBc8TUs9hv+j8mNgshMhkrLRnrqK8n/hh33R5A8v7N/dFLZirOUlg
sYnI34GhEnfhXoR4mcnkhAsQxusNj1DxFAZziHG2sYWKlzPSatV937Sgvl/dAumX
WO2yPSPAFYNWOp6BYcmzNcoI4qkJSFK68CvVyyEcDBhUqjY9fC6lpZrAG/yMDSGq
zXQ4Eh+45KvWI8sfm1n+gF3I5j8tRAAsrhKTUuBCI5u1gQTVEksa8PHLLZPlo8E9
qC/rYMxO3Op7cKiJy6hJRJl01BPyNjHDevsq83QTCk804MHHbFMDwmkwSw6gdFFD
KaS/g7+4y5mMPJIfENN0qM5okSJxzSYe6qhmQgm3ZgK5fVyszdk7UfjpyJ0Ls5IC
ybFcHj46GNpPIvQbdjkJFNJrugk65OpLx16S+v/FdosVqofJeJov9pmi9GK8MfX+
TJH/LQALUZS//Lqy/2TKelpV1izyeHAuDZFq6U1IdKB5e2G4nT/k0+wVKHDY3fSR
Z2qlR/DhW2zTXidMF2GjfNHogyNGtpRZTIkJEw8nvs1uI9i6DTg4qMZ6+XwvihBj
7m6b+3KBreAsYTcZnO6Xgj5k1Kzczo/bvzC64/T7z+9yUks/37Ra3gK1qTY3k5hc
po0uv2wVcieS8bAdJ84od1fSS/+ry8Yl1GuZLtVCItqcnc5MtymAqv7FlbGOFt92
90GFvdafaqsyZ/VeNTnATRO3DusD9CdnACLcNBy5m6SvrJqqewRw4FzfwYd60p/M
K/GnTsTIDsEftIUKNVFceMUADHHoP3YFmMGUYrXfX3XSFRZpzvScA8B193xo9h8D
wcMQrQmj7FyCSuupX4sYIHuAsUXA9PKmh689dnQ+fYO6587tnVQPztLwFVPjw4J9
FtrwhRDsYrbXHXKeTw6iJFCEOicfQWGK9Ao6yyivFecJXFQgvzw0va5OS2Go1TC9
ZHl3CxTXSqVjuTejjwGQxoc643yPcP8ffCgQVC36OXvZyjFPMRVV+m43cq9xTkls
ommqD0GgBmutUJUQmijCp7wsIPxJ41u9vW+4ZNUyOySsA7ae1fasCe4pnJz9/Ygg
t3qAsLcSJ9tvCNUM1CN5xVhjmucMe7YIFYb6TQY+2/H9/8lrqRUAqM2wjJV4GTmQ
hLGTNYchNAvbxSDRlLfD2mpfG4M4wknMqdJbVeVAU8grPtyL7Lrnyqd9oIB4gNAS
HBrdHIBmUXWkRlLvUJ/VK7F4CZ0fUnvKddhC9VavRFgUVZJEjZyqyPEA43CT3ADV
LhlcQNwKo2HSW8leYmiwkPa0DFraAA5Kh+5OzuC3bVXgD6jk6we5aOntYX5kYLiu
5n59h7hTMI65+LQfLnGR76jqUvpbwoSpaZs6eL/A/XuuLBTDRxJY9LVi3Iu+HgSq
z7NZzNk8Rk6tKRfhl/HJn9BVfU+c2nxfbRUrtXbSteo8JUCk8TgkyhBYMYbwYuxj
i5mKf+mCGi6lYrDVknNR9fFveOd+zEi8B9ipT+OOn5X1dsaOPNvLknqn2Q2aZQ2D
NdzrwctP6pYgjugoqwdCua3rYXl6IHoDluLrjGPFJXuECw5cs2C5aGb2PxfubluS
3ahrg5uy9la4LdLYDOhmMMNQarv3z0K97I6Ll3iHnim7lEGjyq+CzsQoHlQXoXDa
uL4cimsawHv0b7Ab5B8WCCssI4fXV+bRbQmojH2oyJVdHSw6qvBjCbfRrqKXkipG
5OZ6j2hvdX8SChIc3ufs5o91D6tdAIebfrqrJNS0Rmrtteet5kFKjEUFSZVvK4BZ
zf7zbG7Ano6upCJmMhOEd+3chmr+zUBg08v4fW+buxGV6RK2KqRC1WakzAZaJZUv
BLzBsX1HjZWBUSLEZ6kCTTgjuGONip/iKfBt1nvcc1O4DTmvcXhlfCaQ4OFzQX4C
qSmBwYqJnrxHNJ6XwfeBH2aus3wYZp+N/gsbu7JR8s27IEYrc7VINgJGRtyNqHvb
M9SvSUN6310KlMu3BnxPKSx0HAdMgNqRFoqT+R/iClcAxAJdKSBEgYW/1GKMCdUD
D2he7j7aZHFw70d55V0GReL6fDqBSNDH4sK8AVynvBNqBNupNZrcLR2G9Rlf3ulv
MsDz+eibFkdqkmwEzYkDkutTGCF8ECitdYRMA3HTOgA0R8+Vp/X9OXyHR1bJ+N+Y
1/KUgaQiPeN2KFaWNvJ9Fw9lfRd5bQWkrWL1SAY9fzOIAYwyl5oCqjQIGxegBOwH
UG4o+5B4/VkbWJVkU3lH0uEnOCVbcVEYc9dmC9FOxnvaZI98EB4htK1U/4ioPSxV
GLw3FcwKLZQar0hRRMpJej15Jtc911OOeoJsgHWO3x9ohP7hRql7VOai9GpV0C2h
vE0e+AliKRtk/yfM3YSdS4aN5MviBeAbK3fFlLR3hMZsHr7f76KYVZfwJY1Ov2ng
60QS3974HsBnpljrsPr7cfcSkmzArIe32hCGTMz/hQ4AUvlD8tI3cqvfwuK8sMAQ
745ypvUV0tEKL8ThTOz2w6KlRFohU2sInW2NNo2c4smKL4Bw7PQrT7Dgm1UZ8C04
wiqN37m5XTHM8+8BOlrrtijggK/n0n1+GvMeYBmZTpEXAaRcVhahqWcvIxifLZXm
mFpV/PQP4bNM6qw1rsGDmOkHS3hV635hvyOL9CjzxhbHZigFCIJnCcl3ona6DPUR
PxUKy8xj/m3St8XRdXuIlnTAQ1LTU3eULAuU35kIvVqaXkFz9d1UemZwYynt83d5
JMGEGm9qLAS1E3k6q3+DwvX8v8yUAr/46tSy+Kn9JxM5V6+S0Tj8uNoVKB3/GDNv
AK4yi0fa6kBVXuqysLpUeXiIgKNG+7X2K13L7/fLqdW4R1nvQKBp1mS9LalCQtn9
G8+Il2oWy3oJWJclvYhVtH7sm0O40R4XUPDdWCXrsmmXf3SK+pF7XJeI2Ge5D7je
lSJBxAdJTebZ6GvvICNAxiQG4fDw873OUnT8cOeDAl/syGboJ9Z3+srXGdAiqCO5
egGKhOHpq7M2fUwL2Th+ZR+yAcU+zTAfxcTFXuMfv/BAN2nnfiInC9f4pTZCXvyZ
8A0tEpjX937c05MTcQZQ/fY8ryVSpZqXenvRfRQpFAD29cdVXyfOCQVhq3ytwtds
EoDdupAfCRD6IACgIYJsw6W+z6Di2+qTsbGCxwEzqQeC2zVjuZhRmnt2REbh5OTy
zU7iobl3sHpb3IesErwcchjJ5xoxWmy0WtN79mguzxp1Izsv57U8gWY4bkGQO6Iq
pBvxilTBs+E6FIyIl9kwzvb9HAG+xnZrq+hAGznBt1iv3vwur2PIMH2ew1z/rLbl
7kQ86FK7BmJP1lomvkAS2vQ7s4ltkmeboSI03GrhtEE3Ss/kBR5e5LMoQ9unnBGN
U7GJWDbdNxZoN9qMmJT56bzo/f5VoGRn5rsG8GWwXAbHZwqoLasadvq6+y3pbJJZ
Fm2v2xXIa/lZyE+M14f8GalPTMDZ4O51X4YpougmhsurS0BPk9qYBbSAlaCxu3lo
69RutSTAMmBlEgVS/rEq38ctLS5rsORbUxvb6S+gW0XUPRp1I8yy8KHTZshm0/0Z
3Ac3AUor4envq6WDvkRKIfXoBB/1LnR9BmgpsEBMihtWpzuwDH6IIdRo5XJWo++Q
igHFFKQ2AFU8r7pBXJLJF+PLwaLKDdXB4P/dCgURHHHS9wJTz20RlcQ+TVwER698
T2VUyXzYmTz5nPc+UlZHtH1kl8Jo80TXWGBTR9e7kNNAA+g2ZDp4u55RBVhl5g25
79yaCnfYc1TihtokUGsHzFP2fNPPJCrvpwBQ31HnZwPqGrRR6l+fjkQe+WzMWu+1
x8maJy7EIumFU6fjVH0WSTyT0dgJYaWFsfZfhuq1J205/sGTJrTCM64shpa9Dj9m
+5M6M26pUJj1679zCWGvgu5ZZv6LiCYmPFZoldQQmZ/o7zeiDVROKEWlxDJyAhsF
c2qwu2Xt8phCQPotEQp2KUWc+A664NzIMEuYB/W/vA8F4y3o2+A/1SXt01FHZA9i
6G8BJZCp04BG1VZW2kofOEXmWItj8hQa8U1jUodhA0n3KnqCjC0QowKWiHZj0d7/
KgFFFVNmhZqRftDCmDsRzQZOTdFHmFeevqV9Yt2wGH29SGV/CJZuxENJQXpdNFc3
xgyNUSdXEiuKOCYSDcpv6UfScxmZRNxgJdqs8DwMeoEb5oDkGcfh65qlCjpY23lp
sYygKFem/dfSueowDlhV4ItAct1obOQzcgjjrXPIhOj4PMn46aiC06wXCTzgF3vr
ZbIRxkagoaaSPiAgeJWNkysB2CI/pDjA13Or2XSCASrdT2f1fXoBpOJpI2F/wTpI
CEd8iNY3yJsbe0TSSYO3Dtd6fPcK3jmv4AA5rkGQewdgP9kLQlqlDaLco5S4LmdP
aWn/4t8crRERKHP9lKPmloHrNqwbcwH5JPart0G/h30sR+dKZU1iGJAOtya2CAtJ
s9uAYzJiw2Ex53NszbI4PXCnd7LrzZCY4z79Ahhf4pLSR/TQzP0wc8iR8wSHJYlO
yu20d1Ttz23+Gjdils8hGwHKYdY0hLIz9g5l6gm42NVNlomcVw6r7WRf+eaPHW4F
xPLNYcI+KZkXH40Feq8a19nsbdEU/lWoC1X5FXE3t1uMQHjE1SifrBr53G6Ej2k5
4YR1NjWpG26Q/bivmKUjOtLjj/e2QFJaigqge9x6Sy8WrhMflMD8uImBdZ0YTXtC
R2GNaY8DbxYb78X5HNLGG5xbaDrA3wqBT+ZyzhKVf+FkYg0Jvz6bojdFF8mWtEDQ
6ubOvlM8eWFnNOuNPdeUQWsz5+j9zml27hH/l04wBGBonoHil/1QslgbNm98GDVw
AWYr7BQLzuuGwPWcJ0qUrMQv22UM9hmx200Qbi1xyZEnie5ka5kvV2WDM1v9i694
Uu5kN4+aJCjemdMgutUn7nIq5+3E8neEoEE7Q61jhUgB6Dyx4wDSLM0F2BXw1pPJ
ep1aiHLSm1QA7PyRGqJaYsH7K2kkY9zPkxqJ6wax03yxewict9LBuINUvIx9tFYS
CSVvYMPCg8tNl2oYqrBsk5G4rv+AHP/FAwOJeuqw8Hg9kVR/seOB+6mf7itSlS8j
qzibFQkjXZg3g0Jh7LTMe4Bpyg4ULcIjoaGvtfi7oOhdhvcqLayEUCoJ1gpt7KxZ
lbYBLj8RJseGWKLpReOCM5MojZ7jbJ+FhKtL7K8Ze1Zc1Xw/03vmRRFRO3tK2+Xa
Q1FOdQqLVBpz3EdVAfh9fgV+U/DVDyb5ezqse5THtdvXXQHgIU54j1AwNfhWxTO0
CQg0p8tECeqesQZv6w3nbJM42SlceDNrVAS2ihs72kqbxdzQzyZ+txFDdkeP7ebK
8iPzCP2GGNzaxsqUH16tSGKugoiY42HqQT9x5hGxmzPI0wIB4Zb1L6pKsoMvk1Z1
JUIdGm4yEZ/r3DqjwKiWRc+fNhCqzzy6wz4dEEH6vd7bYMHRWFlCXG31l7zvmO4u
uamxR0wrdZdScMoWt1yUXF2YuWFejb+AeEAERAEugFcAYEsiuUwObCue1N2CgBIx
Ok7hc5jDUQyBMC0CCbsTGmI/sNs7V0pcAiDXcrKR7Wgm3pHIhDK34OF+WsgRSibq
PINEmf0uZDORiBvkyGfhyLkIMmZPwJkRWK4kIb2PPOWorxhjCDvN3a4Yo8SHTRKL
pbGLdYfNSC/GuRYMamvk98p75bABY+RBIjOjqYLLpYqug4aqcPfSr+Wyp9ayNnmP
9zdChqfMqJDLYGu9Zuh3Q8qIEyQJNmaOo3zTSoDNJS85UFrjFIYt+35QS5no/bLe
07W92n+OwUGTF1UDgWhcWiaLJSFcQuAwE8bDya1p7Up9Ng8IwFOWz9zajOYWBxYh
Zoz8JJb+RyIYULe85Y5ihA2WHtaAgqEHO7ROT4c02Ls+QMV6ID/6ApQrHYR7G7jR
WsHQP/72ot1sgEW+iVbYe+4LuN8Kj+sVzfkcICgywnwdKBPzG3es9q9aoCgKPydF
JR3MqOWt4UgTFNGTEZXQ0owXoupLCTcpkuPwbYtvk0LxctIQuBMJqMZM+wgWOts2
jHM/CQQHyo+UbygDxP9PLp+Xj9yCKEnUC4v6AK7ium4cZkvG2NWuELeHxamlI7JG
kQg6CmBN8kd0CSDokyQpK5A1mhruWKERvLtWXoTsqyZORFmoCSmGSsG1hdz445Hs
u4TXPhe/+DXwq2vJJ7Gf4wq5Kw4SKdbjuy97wv8DmbxaqNK3SDngfxuAGnpgHoVg
quErQjV3dnFvnyr+znbwUCKyIdVdUbMsi8rBVBMndGpnE74UL/iO8a2rvwc3Q8cD
bKTKnGAmRNM0YidHxd/Z7HgjQdkA/HvCykt+kDmmk6FZwTQB+qAHqXY2503h3Ub/
xwk3uIbW31qvdMLmuePRecSTMc6YRL1YZLdYVWm4k8ALjJuHIfscp87zjZTjgW/r
NqQeJIHF+4u1SwZQEVKAZ5WCLl4sS8HdY8YNm//UkERzsSYIyFT+o61GHmElZugO
XYnUwPWPT8mPPxaiElW8NTjJcDgG9Qv5DrJutM1k72esrog4k1NliKqJ9yPkaC+B
EAjgZPiXkKVU6GE9xElEqB0jq2cvgB7K3oDGtOWn+qC+8hNb0BpdUyURN2O67I0X
3cRoY+56wtGunOVQ4DpTpSAUMl0hZcSyKhJkMa0ncW83fycS0soLtQnzQCGyKUmW
rn/vVg/O7p0mzSxl0Dbx8W98LbWo8FS0UvLlmehRm9hFwTdAcSb0DtEmJbZ1CO2z
pKF3hP8q7OEcq6f6r28+lOptb970/uG3o+tI0KJTagrXDzuHymIqACtSXTtUqjXe
qatmMkyrYQimxG1q6SWWWh5CF9gwFOK7TUF9X19baiDlLJrpYSrU0erO2Ac9o7df
6F8SIVeR/ghC6ab152OeCAp/SQKvMz03s++//s3Nwy7S4s5WScyZdho8XolPep9O
YB7gpFnpw2tzUb5p2Heg81w/JR2jz+d0j7rCryktpUN2KKKYaaYzB073a2XHh4vf
kEOrzHW8+mYajhipaBAH7FxABJjaUnGEZvIc3LS6yc00qXDK0YrniSneRCOuQkvy
gDedYDrrscsYZD9e3DvnSbYlX8aEwx2V7SR50Zhi+JhaNz9Asj9Sq8oiWWvjUpEO
RzAcRZoibxuR+s8wbCwU0tKomRVFYTuQ/X9TOlIjtow+SSb+n6gPsQ1TnIGgtnGO
grec8oEFJbz2krnPCLe3BvwYgE4J9MD05pn/tlXSauBY1OVhWApcJzVoz6QEUM+8
ZnsYSEnPhhfDwwC0KP56dssDvICSQ1Cbt0DRd1oLGbzzKqGqACE0Eg3F+mtp9/h3
1U1lB4A0E1pGjIJYrjaGIL/f8Sbi3tF3fKiRfPh7+Pnhu7NnHGvbuO3poJvvHhhV
DNyAbhY05PUpaecrBXOfCwYBnlEhrpVOEhRfsc/8sEeUtdIEBonTmQCL6zj5wQEW
hcJZxvCgHnlbq0rxG+/B4g81QL73XoIf+BQDoMKOQWyxlJCw6O3fpNID2T2cWLcn
CjDf6oxwe+7b2gJHn6+ClUXfaFlMvfy2PosEE0zr8MasoshTbPHtF9I18WqxqF5M
fs1YD0LODInZTQehMhg2EqbQxhmJFWq+p1HT+1IinxDywcODj34K7ZBY5O1EJIVe
+FAAuPWI3VTJcDV8gDgqy4NLWYK928mcoLZpaEfeRYhaS5eBOxDkss1KqYF9ZXo+
7DYbuPP5d0ejau0bmR3+b/E/m7kUZma6YH/+niSegF9xTr7ZeYqyCF8XHJ7+2+Xv
d3jYrdFS9UbgzII4y/Z7CnUfJlTJJXyn1/N2i5tGauSsDT0BsQGGD0sXVzEy2Vf/
tBPMYFMaNJttvqX/PimK8GtkXQ+MNOtA9jCYuEiAuiu4dR01b2OCPCyWRNVuTu9l
i3DmjmnWRgej5HHgxAV776exEFMtg5DkfR/U9l7W3iLYI0nJ21EU8+C4hADu+A7d
dbZIa77qoktKgw3h/wQhhxXaWmPt/gGw3y7xrDSJmCpqByYXbmnwdvvpN01fawAK
DaJUEKFaR6hcd0VQ9/XGl02MNeYH2aKl1jQ6leI/QwmIjbqdfY3bcdZXyV4DAqFe
8qJ0xX5FEP7fI1m00HeklGfM1r5IeCtmzdyvtGE2HfqvR1s30+z1c6K+V8veuEon
6Yxu+AwsB9Sc+OuVZ4kWqLoB5+XRjTHpjnSoLMKImBY+KDdaqcRWdmO7f1IEGaFp
c1oRvrsiQ6YfslBQRI3+nO6693uAvxCN2igurB9K+0fOMIJ9hCdBiQ+875+2QhWY
dCPl0sMfpEBNRbtq8B1Dg8TnUvjgIr82dfnGYfYT/axmPUOZ+oN5j2P/BQHPzxaE
5OHp7U/bovk9j3MD0u6diki8DGv0reBAk9fhhQ9cJ18tLME0hkPCKKOapCyNKiHL
aiZzmR+IWg9VoJfPpUuUL2X0hcHfbjPSECqDM1H1ImMPLVqkbwyVPr931VCCWja9
5CLvMFQWtyBtY1l5mV2pggNdgIaX6zXbhsmKGGxI0S45Y/c78gythiv7BkHdUKQA
Hjdpq37Yh7+/MTnQquodZIO4U8KCX8+QzsUr7JQ8jYOPa1D5+8V+x3A8hB/3xNeb
liDAXMoGWDYk1r00y1KhuQdwfOfTft57/YtYlualF6cH0omZ7ydB3yJBH8j3uIOZ
OWxTPuVdRSmpuDH1vmXZ2cNx+B2AjOkbornv6t+vFq64MhwQHixq9KKnu3QbcQCq
avS60iO3NtbTkgfM6CiMKcwKA7dyUZcBWg90gj9eJcfsZ7z83O5WD/nqpdk/kcJr
wv6sQyIrqwLjy/QtdjQhwQPFAlKKrqKml7FA8kPSoM5wTUaDKYzePeMGNNsqG6ID
9SKTAN2OPncd+ZvfxnivBjsNIXd/3Z7Zcgm9hljs0tiPC1kf0bsUJ2BPW1h8QmgH
Se7uTX0aLtUWne7M9B1fbNX+KdBzd4HU53fOVSu3G3o3llg12hBOz5SOktsWoXe2
WvmB9VZfTIDpzYWC36TonJ9mcaIK32HcewOxfNkMMB/SezkQHztwn3pQKLJDwk5B
hXO5vz6wvhFX+wmugfVSwkHly+HF8il3EhTsdC/SPJRn9iuvDHhwDrsa8vcAHdnD
k6heGc5vTIgiAFpVfPQirLfkYnTdbkW6WScDxCsGQ8M1wHa30hNJtqxCeTSEhj6W
9hF5UQgLfZevXgHhF83OqmZS1FNwUkr/CVCfnyd0tyf3o8t/m6eV2RcgYL7z6va1
ze0MkKNzIrhdsRm/Tsg3ATmbUk7W9U22zcRXwtefK6GYZ4BPGE2BHIB8N/3VwQ4c
4OUy8GRZIeJZ5ZSbPNd0anmAqW6lSD1rQwi1VcTuNNGEud0xCsiBHxl+33vOe/uw
SoCr3ogbMM0ZZb3EPeI5/u23yxiY/NSQ0Jg+YRzE8CfmQDBBGzWNcoj795WdQpB/
JpTIyKDtqtvdUgZZcapzRlfCzIOby6a2eUK+zHBtI+sX5QwaKKNENL+tzgNXwmAS
r4t/4K+DvEvbYVAHVEojXqD5k60Zh5LUkeRkt79LxMgcv0o7Cao5sRFfmagNtMG7
h0yAxZ35+grsDJkkpFOq9A2oUO63Ra4wntSLW10CQTFSyGUB9PM0msMDd6w6MIoa
xCEMBAQ6JFH2q6tsjQ90u76tOCITlzw7wz9YHeY0cE4uZgetpqnc3zodF41nPpxu
/JvkVTtzcN2FQmaNvHNqlQoybxKtj8S2dpu4A3ut9LsNZ2PstWr+VOtumB5+NBlr
bSWFfBueCGE6L5iUdwoZXW37XJipSovrBYBRft4EMJ+CAIufdbrfXbpmV0qc0VWs
emX65Tt3jEcfGhtqCpVy2PcZZsVmPx7iGxPlCkGFhvy+kSSyNdrsc7dpYAXJT+Iq
aTbxyKyeB4L9GSwFQRmV94Dz/5xVIrctFq/5PSVSsR+wVtUxTk2vXjlpvNoie53Z
tftBF1+WXrt/GbgQ/AhMOsEaepFsadZr7FBEytP/Pkl/LJ2DqBheOeEF6/03b/WH
LTV+9BNUQyuJQI36IVpDXQoPqfBJCcNEDAhUwRjdNmDnuqM3xXYyxP/U6KNY2aiF
I+WmhGi1KNjM/wp3uScMZbcIoDaumJT+uVRPNfwlCHvXdm9dTk7nV7RqVFHeknwK
bNR4EhLq5mxqaRha1SvPdQaR+zKVVPO5H48/d9BT0HFTIakSQt8sx42+WTsLJjHR
K4EpLouKK6PPHxGVf3eI2SATMHah0bn5L4dIiErhGufiHHEoFR2vj4gw9c6ZiV6n
5gexbnLS2AGbDVIcuPK1if3q4wUbPBKK/DHpiwTv6881My1kLPCkpv+gE+tkM6TH
bkukvefaXHwrwwnkdHO3orQgmGytNQLlawSJpgzfMRyO2ivRTHRMYI+26+kXrgMk
yOEnF3WjHNaia5heURDo8kj4DY5u3dKUQDeIPWwoz3+IaIMh/7kiJT6BfiykOGWO
sYJe8pCnWbR6F7VgxHg/5sg4uEaoG96YoCqbWOctcjnS1bpVBJEA2xksWQK5mgir
VELrQ5N2jLageBVhwQa5hYCWnpdhlxwtLsukiP5e/THPbKBhiEVl0PINp/hNmq8i
2rekhFmyG5DlljlxJgBR14OVNxzO/2eXtwqlT+E+qn1Cdja66ZbBDExV5N1AP95B
DvAROF5Dkc7aZ45anA93I78NytADohzQ28Dc5v5aXsx0CtFXqovMxuQNjhI0cbMe
tfTE89rhIJ/Pzem0nz2AJMRMCFhc+VfMnLgStLIp6OEGssRvFpaZuSIYAiM7+uT+
7gwfWO8tB2wKKPA/9tqQjCrVjz0HJCAY+b6wam7d5iJ8/yj/xKAJxcKJ7U4mNePK
SNY9e5EA7gOMBuqmMBUQyqukgZ35dlORoZ4NKjW0FkgCSag5bYkJvbDG/mJeZ6kz
z//zUwkwm1E4Gs4wiUBrnDmpSXI4g7hEB02JkP9HsDANKEf2ThYTzKggp5IaP1mg
NX2+4RW6sxjwnTfs6L0IZdPniFJrt+UsPHNXKj9u93RuUXskjJch57BaIfmMTfc2
y9+TjJ5sIacf426nS6hCIX8fr+xcXAThXHcJQxOQ0JJ/5ywZDZiasQM7YjktxbVx
1euC6lyoWQtEfzUuL+vZ+gpPz8Wogmz+ceIkfd+yPTLE3qi9sVo34GxFopb9Frhy
c5xKkWc++RgZOtJdVDGo5hv117l7QrN/pzxh0QP3uFmQCsc1ftHQEcaw2VO9Bo8q
tqsNsmKSl7Wraxr16Mk4gi4WpFGGVMRMTHpLoR4RoOefadtbGCnErAy0XQE+n5X/
nqTtAklYhC9xgf7uPs9ftWJvoYd+TGfDasFJQfyifVLt7EphjnSy5WvQ0tT0RxRF
0B/y+nLxWkeikMAmfQVfe6aHWFOocVAg0NIQHSFcqzC+Ok5DVUVntKN7QZG8oXda
PHCKud+xu45wf8GBhphvexNjy9H/8/vHOM/KcwtdrOIv4QnFsHDvZDV3t2KkiWWh
MZPcHSh5Grrwn+TMg5euXMpKmtcd6kYxzRHsr9AdzrsMAUmqjjCDpg92RLLMGIRk
htoRHKmZhIZBT0828dXLfXN1JTb4FSJB4mBaoEHzLfnQlM1WSoklX4B1/Nedcjji
zmeDAkRNpnL9CeCZFOuGTTIT1aA2ju6ukwOby6jBYqha5nMu6iZ/Afgdy9XiPFhL
CH7cSH2VQWQMRpUZslEsNORyUUbKbtNMcQL0bj8qvDfxLadEUXw+5IA3+IsdxIK0
jOlBFDTRGlstNNdXvGjPcoIBM7N1464a9HbgXgLoC8hUokCONYtjolHUcdwdZ0fZ
sRjDG/2Oex3LCtgRgyKweT5SkdNUWIW5nh2mGO4K0fa9/fKy3bqbJ7bK6FCnBWUV
q7hBKWz4Lje0w35l9gCl+21Pe9uetzmsgxVzFHdKQMmZAbPDyXNqVlzQuH7YnDMd
uMDIRXWiuWcmBOj2eeXzvq7CWm0uPzjXjlYNGGoIMcTL0BeIkrHDbo4TCSMymXN+
HToXAIMwlPFCgsQXju7h2kiWO8jERAjclfO2UazllGLs73EyTv7jxNCF3CyfYh2B
auyM9xBKHkHEloolZ2sRal7XLuKsG/dRHlYIDhv763/MI6bqFF5M5gf0YFfPXIT7
yW69yft4Do32DlmaldadvFKkWKai4k43ZvouScXrF5vP4VWeuUDdNFAqhFvXi0Wz
PycOVkjZIIj/nOeVCaIngsg56GO0YRAqq2Ol4wcxrhbzxMSrn8EUVkG6NrEtrl1s
DDicKRBsRsLeie7K3ItTA4zdIGDJaEDIrd/TMM6IkHBsC+XjFRBIg/+t9DMEKMXP
UaB8uKB668R23Q7L/eNrmwzESQTlsrBXqOw4UD9ELsvKrFSo7Q+BiH9XcKuPB/0p
rCs8jfpiTiKf5PItL/bfhlOBVjkSfQwfPlQcZN5DOzRIhO9CBa08qpaHZFt7W5sg
J15goIkQsFXpBxP58/LpwRtPfY/TxjPDpHxqagxmNS2JnfXinAle5ChQFPzIQuqG
p8+nIzQTeglwA1ZCavxgqRQ4k3rgN2K4dywmDK2GEw+F4s1rhphjnb0GM7vrUMCx
seI7BjOKW5MeS2Cbrr8DEmqk1zNk87dPvR1ZRzvtLrzPAHimdPwmQ5ddoDFQtNOr
ZkCywXSeYh9oFzDJaGz/YwAfWFnqzZ1z06Ldrqj0XMAoorZl++68pLOkkUS4NIpu
wbhjHnXGLWurfCwJ/gvBlqF0+IjRsY692Bp3gvftD55XAkKodp6pLVNw/wD5sdpJ
7CA5D6gMYVpy2Ow1dJgohY3Bm6J5mtNb6deMh9ego59ki+cZw2WfR4iJLPezCHyh
7Lv1hPjHZunrGwKHLG/Ak3bKHb2WU8BwKmBqzqe9n2lOr4gC6Mzc736Vkf10hZqh
jNNourhV/Ng9AgVgICHuUKYWwqE0TU0ECSi9gZdjX4aPa19MahZF4WxjSJDEB+IU
QLMXgyueBRBIcAn8qaQhUkpYoq9ECfHyMhAWqTzvAQjp8OpCc0CBMqISzFoWDRdq
pCyd0kvSZMWv7JbuSPmjOI4MBNJ9UT2Hq+QceumzxBoxrBFySuEdwFplzkWOQTn4
QkEbTiD2lD3sBBEcvykD4NGA/5V7qj+zsvfTok2GwMNONbjI9Jq92vmFN/UrJ8cs
FRbFiPzXUuVTshxovfUrMQFZf6xtNZK2Kv7MLE/WrGmIH9ueH6eT4XSPTTpAXix1
hr6Ag/5cZTPkbktI0HUe2G0nM2AJeNHX/LDGC/noikbxUz7smEvcfKVmiiVmFlsR
F8EzAnRTBe38XHbBbqmWFK3ECydTTntWyZR6ZrwUteFkL+QmUvze5UGkD+XanK6v
TRbIBH25885eZBRSN45uVv3n4aRgoqp9jROEsmGHxUjx59tm9NInXdMP9WtHYqP0
RIaS3J6gy/yJ6rwTg+vNrwyLD/yKBPbohu6pBdvQWX+e3GDO8hnnIjT+6d26wRuh
ts/OioJX/0eqiaKXGYx6tTS7HTDGBT5FYB72UUerg18RcUz1TIWTnP0yOpQNeEXr
Vgner0hwHnMfQGbNQ5pX6H25gbHCT4+21SQyOWRLzlTozMcnVAG5ZhjfDNkSPdyE
9rdvd2OVTUpUyaI8A5Kxo5FU4uo0PYhj6iyZw3CQujEXc9qzFvd4jvVl0tQHZ3BS
7dv+qFyS1VAbcwIjGttcx/5YJb6yUDJLxB60AMoe7gSxGKzh22Oa81Qh1EuqZgSP
oTrtPBLxnEdB7FBo2tVfHe+g0f0v79UJVT9uRGpK2Xnb+VhUS1PovEUq+dlbUsxy
bGlV4kXpSQJ/YrymDK7mEnEiKBF1yWlm9nf+9dScvmnR5bN4ikfOOHo/R2Ws2mNp
FOC8JDNSreiFZ4GsdTTfwb87SCr1L4u+6SXLG2WtDV0K9MZiI7DIj7xTS//ZyrBd
pQ7mW9xRyVfJ5xzyVtQyKfTjthqvwrvowpcQdmrBcj+TmwnNI4iWieb/pP+iXoqB
vnXEnpgsIlwBkfN0dQSEgApG0wFJrOLoLAQiBPIGHY7hJDBJ1/RGEtngGeDvH7jO
C0IPsfx09TTSVPAj3NrzEaOmCKDaw+Bnpwq1M8dwJFOqhJhuDOiUZch+wl4SlFMR
uTu2lh3tFhtGc7GDxs8IjLxeHs1UjeRPiRQ3VdYfZnqqBF7nGoNRj6o8R1vckKKW
VlwhsHn7H4A/4OHi2Wne4ZTHrQ74aT/sxdk9NWGJNb+U7Kr9ytA5R3etvf4jwuvs
OxRYd+YWysIcPCNpvtVzeaI8MHHMF92o0k26DapF9tHdTa+D6+cwmbQ4Sh9dk1AW
9UWOqp9hdTadKKpO+Khp6yTM+w1UUeVuwpX+tjqw966ge1Yg8hbStfoMPyIVeXFm
aZh7Wz+Rs9xqq4wfqTCDRQXujL+nlSf6dbcegJ1o1AN0mKa9JTUmI4Xe2dsooFh8
SGTjQdtBIpS2swmyFp4J2wQ13/fN29qCPPR+Np8Gq9slkoFnayFgO33aWaU0Z3TX
MM1XK4v5H/DMIyOgrvZxAh/DVsJsBMwJhUf5r93qXUEV68sUvzEmNdnA2+JhmXFq
stR9VX3XSfXnt5fKfeYCbGNrTLkj5leXRP8FNW8z7M+8Is84bU8GV/XDrBe6uGfF
0fqgJI4H8iW2nIlEDlifOWW9sM4hZBkjGL61Uxk6bRPk6Tf6Uul3rSjpGR11M9G3
gtvI/fpLCeALB7y0FtVXXF7E5KRZDW381+lKGQanCkMDHkmQ7s8zzZR2jhOhYSAQ
o5ibIaXB41nBBGUeH5XVziOWXD1T1e2k5MVYMmbAmINMqrLYrrz06Lan2wlo85Kg
aBq58fWDptsCHArJPrvMvR6r4ekOMkrAe7M2Mds5t9L51++ulRJ3zAV0AWAARVSR
nH95xF69k5/s0hrA+rW1ETkKABTmHMdXVh7H3qvBYVu22JNMdcmdxuF7gBEucq0O
mfGg/vSjr4cAFeqw8x8a6jzF81TgXM6o7UmSFgzivIUGH0vB/0Rf57ngDAbGO249
SWSYjB9pk+qkKGtTvepzLgvdlN7POhYj/K5wi6ZwkG+68zt25CBze/g8Nw7Q9bcP
jFxTm8xHf8PKDKLyVL3x+ajIgmZPEgd0/SxsVyXwErF2QMy9lH+MuG3e4d6Zj/tS
HV4R2mN/jWJCROzyl7s/X3x9qeDkSXztBFgwMnJyTX77fxbju8QMl/mafv+hABSI
AFvBhVRXL8dMK8wZ3R8FU4u59mdkg0HFc2MgeWm5mbFuDLsmv9vm8zyfzGwCmDyr
J9K3V/uH8U0RdpnowIP9VUkYpYDgkFqBBrxoICUiNIjzPRBZ4flm6xowufycEtiK
pc/2W7HpsWTxqPQfJKmaaw/2fUKtU/OUgaRV4t4M2Siyiw12Ys5KE6/JEAQkLM1V
5KMfkUdl/3RrxCTBI4AovSkS/g9r0aJxppNCnXepM4ZF66jKWFC4pDgIf0UNzot+
sz73nqHD3geHlHa5WZeM/skJqmUt0r02zLM2v2P7Lar7kalV8WsbloVukub4fKXo
lqe5OqwOXl2YPyt7dHNLX//aOgh6lEEqk0t862bkHnPlUZCnnVmsxz5u1pUdRSib
E7+cckzyBlJLkqf3NB4Z6ziRUADFEnHpVUzlsxpW+zYoN6hx2xRd5HrVJHzLc/jF
peW/s8Q16nIIB5OmQM5kl+ILTjc+Td0iRoZe9++VPWIPcqwYuo+9LLIv+xAH/AC+
InknmCjl712+Ok9O1uBCXo9Py6s9PJpFnii/HACqg43xiSVb2WUXEf+orUFYipKU
zj2JCyuY7h20KQ/K1zMqGg+YXQYBXgvJDXk4LkEWuQIOJtSV1WWkIoP38jUZHTNj
Q2stUpdC2lDUb9DAdSv7oQnLkJ8rb6wfPHUwjtRmpbWLhhTtPzf1la4w8/kn5cGW
MZW/MYh0haOY9x8WuvVd1wjjA/v4zqOOc6UNp1t5OkqtWlRMG5sT3H9lewQxRUzZ
vwudvuZAEj8puYLSed5ifsmar+FtSTm6OC9IZnjDe/bbPlSkCmgjck4PSQFx91LY
vRPbijBS0g08v8KXTWVtRkkvclXnd53Hz/abV6EZeTXz0IYdLEBOPbC1Qzd6RFFo
pqCBYzjYoKCo2LOogdzOnLeHx96QHaZ/Gtv1TFOvh7N/AU3EMubos4rmxYkE6L8V
zPwMP+jDriUfS1surIkP0u7JFTgysEtlDH6/P6DeXudqGk7vjmeZTeHUIMmbG4Tk
oaXUGVDuGpncEIAMeaR3TcaKMsKGfs/YsdO0KGFSTEfe+rK+1lDkCilr6uqeTUPN
RvAzS+7dgKSk33AsZEw0FTv+SK93CpakC+Y0TlpqFCByzG+Bw3pdBN4d2jkYEDxx
6BsuijneIUeD5I8FdRbYS/uye+O2Svw5i2g3b2JZY+c=
`pragma protect end_protected
