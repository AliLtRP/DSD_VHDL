// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:35:23 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Nu/KQw6YvvkSUQpj3KX2rxyAUJQb4uKyVivk+WV3z5g/nl1lO3HQZnzcEy8ju4Rt
/gZuUZHFtX59vttY3EP3lZoaNRbNvXfuUl5Wss7sU5KLQ9mrS72Aweke42zTyKBk
+CF86To4W77SvPATrXjz9IBXaM8lU/1ZWhqDdwKp17o=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 8544)
pT3QFwyy8v9YOyc3hnkDLaGG+p8/J9ep4+MTyDwDHycL7Kazi+NGvGA6uJ3hYeEV
+NtMIMb88C3OOkef1dd6YtOhaLpzmwLZ7S2Lsi6B7MG5V0Rrw+NXn2CuD2X89vJQ
Srjnnvfm4D4XxN6hwb6dHD5cyMwzgiXvJjYnVvkqXjCtgOnaMQVl8PiktYvNUh4D
Y4Kj2a4jhGGPtCXGB5vOumajhqd6Dg0lj7qfPfY/Ne8TLX/fr6nWTEnOytZzs1Bl
XDzW2pJ8dCfeczJPR6vw9lnqYMBQM7I3WstXSTBIerXJlILmz2sQ4aYM2u2/Zjcl
qz8txMRMW2Z1m9PzenP6NKoZyd2ZuoG/y9MhM42znHE3aZbmr/y0FwV7hgcZxT1F
eWV/xXk8Yx2C/N2sooRDQniSQDivKVTdOpqs6SEX6Hkj/DwW3ela6kmc1uEDqW1P
pYhedBbd3tT1LEwV7pZ3vhAkXC5bdaKM7WmTH8aMPdsXoWtEQZ49R2tlGF3JyI7w
hdJ+ionEvjYAc2S7sKn6OOdRwyMEhDW3fqtemNL2VSaDAo8FCMg9Gike+7fihAFv
ujKLpQpscVf78DslqDkO27X1cvkTuP1Y0NxTOXkzjWXjnaAfYilt0/CypSUgiUQo
aRAE72HNR/9b9zqcDlbHwr/S5xZSos4JBUMbeZEP5XQh5OXaVLcrYSSld4L8jwk0
Mmc5EnL2AUb3qHO7R/Lt6Apz7hnOpKKXJlKsUy3ZZrcfg8rl0WMoPgPcewdaBd7O
RYd4YWxY/3FzqQJGP/rC4NJa+xblpBe93N1rw6K7+Q5QxPbMugsKVtl0h+lCiIug
lPc+gvzCuyTVo0+c7mckpgdn5vCnZ1R+uIHWyBymfEN34l3gOwGXmWyXtsynCdal
QFX8b/l4N1STQ2fHLCgyJ5cEnXwTDwrx/SCFdJqw7MBB5z+q/bRHtZ0r8ituJ+8H
E/3Vjb09jUOU3qhhsx7G43Jx/LRQjHgCdKZPCweXXhvAYCulUOwJpxJ24Rm1SQE7
RFcGoQc+iqCLJK79R8lDdts0FqQosZqpU/xovNVUDeWWBX9Cg4lOh11o4liUJYaw
EAO+gNfuzRSlz7ljlPKK12LgdS4jA1teqp6IWxwS9xcZNhN4If8C/0vQEFz4wJrK
51ZeLglYhNpk3qZeKAtzBmZqE1aQlWbER0iDYES6Z41llBksx7C9YyvCliqloGph
qk01T/ZnmN8hnGmE8YMWL9OkJcSLEqCgwXEy/adC+uJUe3zscye/TAZY7sSfZqzw
Od7p9S/a6FtK4fW5U1Q/8fWWmYEesxeY6JHcYSkenVqeVqUNd4vtk5kQZW2Y3BlE
73LrKD3aDP5uxowvRdRuUyV4wm8jOIJjAOh4khNMhM5MLxvWg9j3XybreKfJB20C
xh4ydjzwG38zxiNQwD/UMgBROs0lBY4xC4xsz2ourMrHigQNqlZ83ti+alIU1BaQ
c6RyxC9DwFpMS2zmqtpNsqzSqxIU9Ixm26HPPCforQhmDfyNqqDtpNdwWHLEtNAl
2NgVWam7PsSK+1r4PpCWip+AI0wJCtRzLiQZ3fwCdaL52qDQMb1gIJ6ltnZkjkaQ
4UTD2+298LcONR8ZwbJc3OE7pO8w5QmUR7q6vD0fVI1uidn9xOxoNjPnfNlKtEd/
i3wpdZHgTQAMMsbf6mCN/zDJFR0rR24QO3lLyPw//qMPOT4ZMz3jH2hK+f1U6e3O
yDktHfiLfh7PQeNgjxvx2LLL2wkKqR9v2/vo2tBdSkNkJtb7suOhT5yVGd3rHlGD
LHuKC4tnmLR+Klw6iICtI6VhCWXzLh7UKHjVSZbvRAMCA7D38uNP38NaNz3GCCIw
RHaNt3F1cVCzwHrvtkndA+8DHV5WlRe1kE1h6kgUTjAUsmKiPXtK+t/hSjeW2lvJ
3lGGSC/Oqnvj+HCG0YH+jSrJNMLytUbNjBB3hTsDXFwIGKLpdON8tZ6u3DPzhFhl
+PgrXmWkgRkO3h0kfHbHGTcym+qDVp+NeVCmuPwOiGi9oMhVge6eysiQ3Ayvgbkk
6ZvuDv2SGw2GdNPSrzSbtazrSl+IbRrLab5S3qQm18GII7Gbc5TVcXuFO5BSp48R
TPx0r1apngZ3gl1OquPHXvYWeiuSU/b8WuqfQxVwZ0MxL4Zi+vpeQH+5S5LyiNGu
g2tgcc4ZBDx2W8aJOJ7FLpvEiw0zozkrZH1lJrznjvrJeMIzJdy8QMTwSTRVpJhE
KoB+gkFPoznZY7sT6xhybRDa1ZjI7R+Ql6dpdetYS6yjq0212ZTIPP7FThlyar7M
bkjsUeW/04pUQ71hqONhuILYHRR9awbVb5wAH7QecXX5q0TDM+TN2NMbFHvLvP7R
evCUw9JFQkemrqzdKyP5PAUhgBEtgueqf03kRH3elcXE0rTPdeljln7M4zyWIjFo
njKb0MfWPcwujFPgTYBdk7EoJtf7YWbfBNtmauGptX2v2eB3oHKIrpiEyHMN4xHK
lThZE9d/c1k893mh4noDjNYljLtGMJTNHeO8Ag0xbVhKsdH9ZGJGs9K9lEXTFnWw
p6ojJhKUO7JsyPrJH659m0cqMTlx9WGrTNtPaDvkRc6/uLnEJqAZDstr7iuLktqP
8shwxuhf05zYT14WuGUgBk2F7gMwoBKcprPQ2C0dQzfhoUQ/660Ke8q8qHGGqQaY
kFswKbCb9uEArSiAtrGriue5AgEYX+Xeg6+nMLEc067osR7XgRsCyhgJQss18g4B
i2E8OPH0ngn/GdpGRk3WhRQPWlBYgzQl21VBbDqzESiyXuXSmd0vt7JWJ0hsnDw4
Sqw1oUUTbFJEcGfD0tV5pyg8RFB05HxPhnFH/PnrzhsVfF1ksUjCp0gv4/+2UBR1
D+s0RX7fJuf06V1Ae6AMmQrxrg99yRez/J4sV+IGD/PJFGwbEPRaxTildcERFzgw
IVY30ER9vniSb8JhVWbio2yeWq4TYQLiyFmSORJWuC4iK3yLyJnD2w2Ao9ktEsTb
SiG4XqoUgie+0iz5zvxFmuTEZLg9pPcVha0LS2wyyNzHWW7zs9/BiZJ6dqrGjbbb
jI8/XhryrdR5I0YXJyBT8UC/S/K6gqlr7dTvcBbHxM5Q62Dq+sIwZPOS0mWe+CZM
GzILamkd2uMSdmoMRgGeFoh/V408mtbMpy4PHVT7EOhcU4I/NiXUhMSYCCdHhlSI
cbvl6k0GxqCuSX8Gq8Y658aVpKbKlQ/6ujbh1q5qcLgO7dfwcgRSp/LZwslQztU3
Inju9tq00HBjAdL0P2jSlbejoFf/GCcsHhaMP3t0IiWJagTG2EGBvpo44XA/I0Eo
hVUYV7F95SpyWNNls64uSn22Vb7QE/oejvafZRaVeMe61Pz0PtUx/GprfFt2un0r
k2pUJv6mJ5L3Gl6wLoAFdIR9Ge5DzIoAfXTUbe3txfJyILggpos5FocieYxEtrV8
X6N1XEjhxRnL1sj7s4icO1BfSsT0Hj/25u5X1EQwrm5gwac/UNkvCLvgPQJd8xH5
xIXS2liVhmFlRhO5BGY5czyjoX9GwAjNohr0ItvlYBaI16MBFpWReee/PS1VzSBO
UpmZxW8OVBOAIDLeyheE8cw5x6zuQQIRHGWv6PN5NOpzCawrE8IjsVEY1KMo4sia
oKwBVZGR7dd07RgB1Fq/zi7pyss1Fka8V16xXCRCJVTpkNn8cWEpMkMybpkCD9YU
fiwbeRkP4tLZtW0FlAuC8xFHFG4eIhuuiMZlk0mt/G2WSAnSQU/MIL7iPKflXOy3
YWTDSQ1ng4SGkp5AvwvG+P4PeFy1JHdhNTXkVIp5T/C5qsURPOiafENBITTJsgfH
jVyB1G/d3ivSXkIHtspBZUgiwrgQMFy8ISFEdOQURuttYUCTzhg6H/WogbUPkKWr
jXx8AwdKZDTG1tyg4r6nhc3GwgiinifG0bLAXrx24kPR5bLSRL9YD8Jq/B2LPKtA
WvtM0oiv0QyplvvMvKW6YKlkOpzVNJJII/djsjUg80JCusm3QJbXRPgrfIK/mbLo
+U5jCPbAN+Em6B7j73hT8l6QICp1rN3IBjB7P1DCkbD5uqugz9ijXDkltguaKOFB
8t5bEo6KjXkHZTP1wJHBYonG0mJB5Edazy+JdflxS1pCPym7EMCwvuCPBB37wtPk
+f0vMRlx43bvaTglIOBmC0EC+anIFxPU8VN2E03pdlQcnNCDGJk5TZ7bPMBQbk/K
HuIte3d46XnI6lvIdp7o9/OwO0qS1eWMYnkg9o5vY6rmFqOWp2XNgS0R63VB6XrJ
Hu7VpFU9e//8WxGKpI7vmJ2A4HrbmRL1P8yjn2ynKqfCPI+tv73i2UZVxbKSp6wt
/XQWyTYAmqOhhWJN7ZpvSpS7nkrjPnplaK1/q/kQ5dUFgsXHbifb7MnwVkGYB244
scmhRmhZQSgitxz8rxLKyHbt6F7TKA0R8+Q48p2vV3IGcpsTTP7KeSlAjPMWxASZ
TYCDbE0DgmrNEc/Teevfjix24cMGRvWf124wGzpW3s7fJ/70isCra5/kv9TiZFNy
vAHjZuhmgCdyTVyKHeGX3Tdq+BGt6uLbGf4v49pZS6gP5VLe5eCQGwLMeg3jDYj0
N3f4VzvwvRVOWiwDworMZzjSlE0dUYEMu0jaAinEWQwVtHwXxQ2GeJiq1shgkVRh
rsJ5jGA30EBGHs7izL0mI3SVhJh3/Lz9WcGJD0y+ySkeSJ1KP8UCn7Zhtqv4FSjj
xdNEmFYgpk/Ndo2FfdxFnGT8+qpLejgfC2FnC80OOp98b7RAwuIZLzzQBA/tKh7L
5ZPVdpxlo4K0jXiTj9ksuVfRWchksbW75NNkCBBaXxDLtJS7pnyffgRdoeSMcDDn
r+m/2EsGIxzXvt96j4C3dHSKK8Kgdm5yzInt60ijnZUZgwnDsbkqC4s7g8eKYkmG
7QK4K6aXbDxd0qIrFwrJABQwn6LlWFOewbc7AMuM5s64/U0siAeypHJIILfMJa9G
0oNUMAfiCfnT5gJxpJLAOO16HF2Z6pxUTQsloGgj7jFkx4H2evAe7flKEIvrL3LW
9gs5fUQkv7ymQfDSgSmiFiU6c5wCAfNtqhTZMsUa932HM1kPctWkToQ8CtEUOaxS
ke5tvnqBvRM6pK8VLkaZuO+lRX7n3PRHOuHGTYgrGIirIUu9potxLUsooVU7kKGA
Q1EWMnuAAOjmqeHpaz/clWDtLMubznuo1Vkgv+nxwleCeEJViZxMYa588ZMf8sjf
zlrtKSMeG2lO1OHfTEzZcZzSkGs4HWwu7pDRrC/3BT3z8fjutCQPvfI1VQ+uc8CO
hk4hmVlRqFvfJSWLRX0DMqHK6hx5bqX35svfgXQukiF21XyzKluLp5c1z+y/6djN
6d/9UosHhz3SKH4BQiEOlnojFQSBlyGC5PDd/KhdalhbDWzGFvBM98iue+94vhv2
sZFhdTwIrWDE58dMx3kLTTbLrGc+3tEy9HPADzq35EyxZACt04YuKdBbAJ3OfSq7
OpzRR5EKMOWY7+myIB18LlVkhIqmX4R+CncYXCDo6eJIpu5RvlJzXt5zdMSFZT3I
yZ0K5miaT8M9fs7QjooiFNaNbswvozxwPnwPB4VuqQYfx4ZWfP26n6XEGt1eLJ7y
Zr7hUSFkb3+WDZSlQb/du1BNO990fEhb7pKRKHgypaAqF6guOxVjOBjh+nZjoNo3
OS8HgRhWSKoNq+UWZSIoC3UYW006Uxie4UDM7aLwxexlvoNXHPunHfOn1SYfTqYm
qtqq7kFI5mN1cMpXmrJfYNvN347Q1QcC1IcopOQXxJHLZHaQVE/EEp+erc5KOuin
kgDyxgxbKlENxV/DvXjWM+Vyad5h7Q8Lj8nNfQCSxIGyKOosSFUcLCVUO8LKw5hY
xNlmQDB5tNwJdJ4onDGTKyEuVRp9yvgCUoVEWUcaCJ5QdyknLMvVC5NhpuXoVAXX
NKkFJm71ygCgTBsLSOS6MF5u8cCxOk7S1+Uiymlses/voLygvFPuN9NHr8Hp9aQ1
Yvt9hI+17tlkXic7Yq4cP9lgnRyxys9ICmd7sxDEqt5uxdxLCqhqPJJZ1gUSwWqb
dkqvvdcev5Va67qRvpVkuOYgNiPfsqONANQA6GVqmlaCQEdpJ2WbakBGazpe7ICD
Ifbp8kjWCG1k3olQQvl52Y/YvMAOr+Rszve26s944kxCVtaIK4U7iOgTDtMF95Oa
loTVhvsoUi198h6+l2HYRX490/vnvxqgtSmiaHouL5cUAjl60IwRbslxCVNxBQVi
CFoC/DvMSbWTG04Y4gzN2Y52wiOHxLupRxiaZFh//1zXDCs9I2OafgZsUZgToBFw
gjifMLJe8Kt07Vty2Jcq+dYlRmpI335EzXJK6U4tm0JgOF+AsuiXigGfXkeJFFns
ANPvpRSvKkpupHSyT5jdMZ3J1FTC1StGmfIhmEMYR9xU7kiGC1D8XlnYTUoqIWuZ
eMsKjHt/+6MwYUUn959BgP2ricMZAmmbDxbposMzH6G5bwUtDQyflk8f/nVD5LRU
UYrCShNQ/a75NRR6konOWk4VJMbZj9Y8/o+Z7HHsPTiWRFdmAF1GKL8SRX2QCDg9
by8Sgj3ywE3rZJBNAVe3pnWfbK7AfBBMVdwKcz/g6GnexVzOQqwN4lU9vgWnqccR
I4Al1hg/mvAkP4rcnAcrAyeJTTILCNbc54pOcUQoiRnUNwd5oKiJtnGVfokeWMIF
MnJMEgkORlF6aD9hy29XQ/rKAYQiH9ABfzRxZmFt3Cb1t4FDXTWovhO3IdOFo93a
Fc1vrZkcEtlWRI3P1HlsT3C3kPUOwlJyZfJXi3iPKXTRF+COeaWLOyKQJUH1SNBk
UCB9CtGy0XloBl3WRcjFw/SB47Up34zipwqHR4jH/Ar/8YBolPyqajaNehNExJqD
DvQIRtJv1TS/IPc+MXZgft3MP4d6cCI0zTaKS091H6U9PGLx/x1dCytlYQN+Kp/N
XUZe3xpRMKLRPrPPSzCF8kHt+vIWHN9GvAhLRMsOagYwx2Ci2JInJJFVjgKj034J
OEEHrL3SkP8hCBjMfg/ZVq8pfaebQqb+dNcJxZJRAwghlrZ79TiQFK1ujBd+oufn
7Bnl70cC/MuPB/+fHD9k06231Up9K2qzI8/YiNwDRHKdklNVBv1qpsxgboeQaBSe
REIbTZt1LBCjM2UzXGa1IMirbVoC7WqDsgyoABNW5Rwv9Ba7oAkZNKmtWHKW0T56
wa852cQCFPb9G0GfOjhBRHO36gm1g/2PVs+9EHSo7ewud6tr8cMNoZqzgElRg+6G
d26Uw2CjhK9jllQUAGB31RkN7rJgt6BH61UCshmqdvuDA2BIyXYbcUcVAz2xS85g
9tpG12YxXqYMfXYy2fH1cy1f4M+5JQNaI8TBHs8z5AmiNwA18JSExfpHRVckaPMu
Ab3UXoHcCQbTn5pzzWIYa986Vmxth7fXihG7bQLnaDh8U9RYjXKM2jG1f9MPzefl
coveazw0BSvHxhH5hJnyv5ORtKPRpMx4lVI9qgt+YJh/HFnGG0Lnugzb5cb2pqpz
4uHeNPNgq6BOsPPzAaZBpq4szFfcvntqBkFeunfx+t0eY3iAr46OaMeX7OtLQR0e
LsRFO1w//yYrX8z08IFOi/V709QgOawr2MxoB7D6o6OgMYxiwjUMC+PzlxXbZoPl
xY7AIySbOhOHZhg3e57qs9JZHHkrg50oklhbVLWpN3IL+mykxlXYAEU6OV2xoLeN
2tiSBOPOA3YCAdoOa7LwpxfmptznAZDIQPEsUk0v3yfadQMZbMfHaRMS/DSLZv1a
oLVkStEMuylmXoXBtRx7A4tCQ/Ns7okYnyJdYE7Z/7jSnNF3c2T/DeJiV5oV++sG
+Dak+e2K0+9aZ4iaeCuWRZb+WHncjnDlDSG+DWo96kpAQ9La4y1yOVuPSO91tEoR
8ReZvx21xLVQE5nyqmhyzqWJoYXVuvWmfYKy3JclOU50SlhAYy2Jy67GHRN5XPRv
TpThplYDwlaWsX9xWzck0qKb2AYETBkmlI2ncMD4hoiz8BtuiiDtY7GKuxTqiedh
dVHOVJrvg4kTPW8hD4jBSr0Pr3X1PA7hi64Z76tSne+v80o4NCPwm15cBVWktfR0
25TQQMU2Q6bn/LNG3jTRND2AVOhFA52LxoGdJ9Eg3RzxIXwcq6sJfbNkYCZGNY6D
+Rvsx03TUEXl+ne+wN+o++qduXxR8KZvah+D4f35izkcAEaB3mxmTMPxXvZQqPb9
a5Xkc30aAnTEFerZ84wYZg7QsKw33EhLJs0mwyWBohgHE9KLVDf5KkNq8MvirA2H
/1zaJ4FE/kl9idqf4AR/ZghxfEGpw45LHRZ0w9fJxRKdWMwpxLiZ3+HGVxZnqFSh
iD3K7/PLUPdmFnC8/+B5qyj+pHaoDLmLhgEFvxFptt1cmMapiQV7/VlRP/O9wwV8
mAHYu/EpCKeAxckZ0rzBimMnkt+Kn25NRSNdjPsKvpbYYlX9uQPNg7pjY39yo7JL
2fk+0zv3R0jE5kQVDvFkWqTLcO6rh8RiKLs98S8cTncvede/gHFIt/BhEQ4PtuAm
eQcvg/o1YeUVHgEEoY3ezw63w8hgD3uPUOpvd0mWVPkZI2lw8LXs3N6n8k/WHIaa
tGo2d4V5hP1YKrwSgj07kxEbBSs0Vi+06Yl+ct1KU6ncTm8UKjot91oYjOvl6LTi
r4y3NhZEL3XflkO+MEDl1JUrFSTJ8xRfhxQ591EVVnbAprh4fcMBQCCpaxznKd30
cky25VW39j4aN3VGR86J92Ku4Uj3Cx0TH+vd9GwCaBztN5buQ0IjNeFNMKumdwdq
wvNfEcUFkDBwqR6Yn7buKAu3VvidH9aLcTSI+7IXMshehiwxFPgTD9bkSgDDzsDE
DGYGj3aWoL7scbNf1mAE6PHjcNy8PgLLkN4bIOgE9QUYI68PBtpFmGdKBKBD/2oB
qnyegxmB9YZ8+DjQu0CxWQjJV+vyl+FpPSXvTP/t7p7cEdfst6Jy6a/DylpQ+8Mk
X3Wj7gHmdFG9i4WgZN2GW+F8l5d8ViP7x3uGK+dLgfaOpQu2zSqj7ydeso7figYj
XJsErxoypZi/B+8IlPySHtxnDGnJLNfnb/lFgm6HhZ6jEarlbMeaBLaBcHKaapmp
6H1zWpSs0N8Y99UXb2Kp9bxIGE8o9j97SgJBRmMXICW2PfpPLrTR+qA70Z7QWpp6
0216H1zx7FLh/19teOA8f3sexEZYkkCnIZeQWwrrOp8NQNygs/OVbsyjexY3iMHh
dBOu8LWXwFXGlerXLcym4aeQg31KE1PmG5042Rd77BFtMkyMJnsymUsiCEWSTKpp
NzfOgtEAvI5BZSYfVdBGrTt/fIvNf8TmSMbZkVEnTrSFzJIYfFji3XPM1+hSrtai
QYqi5faMbNtIsb0mz4R0j6xrLhqxReVZnJUhQ2Rf2Nt94juxSkwrZlwy1qO02OcL
LKzx8+7LHyrJtIU+3H9DsIgG/tVF5oKYEiwcXxjyQhGl7AjWvEEIkOydSEwyY+vk
Rv3A6AGyI03jGbbdMVJcMrtDkuvFXvIWVmfij+IdQJ7AH7rnwKU8yO40ZaaJcrCj
9uO0eTxhLTl1qXkwqlJiVp/4JaG6iXwr2JKIafoVH34aSTmh5LWDcIV5HwFZWjnx
+5jH12nxVnud/K/xJlw+wx0AIhtQEvZhXQx+3BdDOC8SUpRWTS+0vPaZ+2QPTzdy
neZY8puKfz57YKH+6yElMfLWd+OBICgN89ROuU8NMVUI2WrG/XVYJ5zNcsjQeEXr
co0XVyDwafXs8Th3j2HjrVO6WQ/a4rjorNKSILEP03yPiH1xC0jT6oTcTPjwhTG+
gZmOjCM3uariOik07xn6qPgSGhkWaCssPnGtUr3yL1Sde3nlgSjUOCQsPMDz4lu2
wW/vhcYs63vxfHrCG7EWjB7v9Xf5pFGt2v1jRPsxPHwOpSysMWQ50x/MGxMdiz2o
o95duuKVTje+SsfVje63kcezhzW/21CoKySikXGjyHHhrPk5NLWDJOA/yqC2rMHR
M+cP/da4lCSvnNlkxMN2YGl3aOJ8FgTPj1lnyO1OhDmAuq7OfsTYVxzPr+PAklA1
UvWt0DeBS/2N5h49y0LBTHzY0yDzm/wRuTkjeeYcqW+0tYK0ZJ2K6a3If3pyWCue
ptNvvzmMIuhFyjZuV/gXt2yKvlqHF8Q1+s2COvurB+9LkUe42DTKmWzCXAF6Z5vP
Pub62DKLW9dORtLK98sl/0M9EmVWqjfg5eBr1cVt1sBprcDfmNLOhNc8rhQhiqv3
F2h/9MS4Ui1jTk5RW83ttwWWX1canWtlaeaB6QC4pBcgGAjwi0IjzfLrWTnok+fm
5irjQaQtvi/2Be4m2ediLRZj6kCZaENNS2GOb37jNgoDoS7R02hjseNSr+UCiPgL
DUFkGdX6Ux9jR24kGra2KI9xzvsz0t3yDN089BQ65B4ra2txWI6XFERXn8+rUgqo
nxzIai/3vdKS44XgytgbIFjO+sKDn0daxjNIMZGtXzv19gilNkqb3gksIlDZlxU+
GEQ+luuCbzYA7Kkrtw9zbYQbf/idD1cQhAQ9v5iB2uND6LNIrjbsO4uDlFAiGZIQ
oEEJgOBOvm1UWPYg6UP3DYT9YuQ24SmFKqyIU5UuQE165hmaiN7R/JsMyl1tS52f
rvp7+LOuQJrsmIi40YoKGgevH2nU3NzQ1zk3vvY2YiQx/I3Do8CJ+UIxcYNwD97g
8aV6G8klpyye7cK3jkoSQYzDd8yOkxZDLFoD9N6ZVKSegGWahWBd16LdLjRtm2+a
W0A2BEPyx+OuqF50cdmp78xE9F4pULk/Ydj8NNmsdk7pw0z89dDInP6SLhyqzsDL
OlwaK1euxWoUD/NJI4rl76nUuHT7GIv9sjDNSnJCeiQEnxinqlyTTJ3W5yoS/7oQ
eF5IvRNblPgod3vIAe5KvaZZEpQ39EdgTDqaCGFipYaaBRsPvIomsEBa5CroH9Ji
Z3ers4Go/uiwPPzsF3qneBE+Fv7cAe6qNSahvlJ5usKmYHAgte6HtRpnIu5cLIgb
alUDif3zZ63XibHN8RIGmrfjHqnwlgo7J3tFOi9KJcrfpeimjHs0z9W0KUoJ+GdQ
YRlfwuYTYzwmlDL7VCElJnU+ssU8Xw8umj9OX9A9A7bgIctK/KjGHXV4UbRF39lZ
OmDoT5s7gj8oZcGVg3KUprEVDfPT6BUxIkBSO4lagTcKqbWWpXha1fuZepOz1yp4
I+RUizxr8cx3PW9BvCptZdA4pz+hXvcUcj35Yx6y86tSvfl1EVXurmBWEHWof8wx
qBXd9ZgBqmWKFkDcHchqJ+DziZynTw7/D3nBStleg0dHPfqeYLDUncqzCJ2mnxBx
`pragma protect end_protected
