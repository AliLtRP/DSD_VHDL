// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:20 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
NSketRC3+gSG3ooQlFR6vgjFSmO/ZOLd84wHb/3P2KeOhjNbIab87ya84rwPm0xN
7V80nDHd1oiiSfU9h1PPsSepGR3tyHqnbttN2fL7YKsBxfqAPIramI3AxMLvTmLz
OUiOU5O0WjmPZbd6UiWYZFsel+pmTzyW2S1Yvl3I7oA=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 112368)
HhVFkn0KpyuaiXYtVnmrJ6/Zg/569IlF91i0Wtr0p7KJ9GUjryrnmO2lKdDVfzR6
JKKtaVOh1cwcL7g/xQXY1IvZpG06d4X9sqpMdqBh4bfIXoo0ku13BXKXmXjmqaSa
pQLp3cPFUF7LBsHL2kOLWHjRL0IWfm77Q+t5CqUN4XZyFtaGlR6UD8d/DOCJtzw7
n+CC2KZJluV1uhGOQRYB9ozZ/WPwS3krQPJijxY04I/EoqwkWu9Zlzol3JlHSIYw
QuIg4gbtvp0yi386OqqOuu4S21BfP7/5NKNw0Qf2nDMlRkk0RZatOG2/rMt2IfHn
p+V39QR6ebncf95s81YDmaQr1nuLW0/I/o9dDpdgsumrx2ysFpWacNO17bMGcJAv
LrimEJ163tXVgnZQVQ9mOmHT/Sm20TLQSof26efJDKoq10/DS2rTMb6QpDPBmf3I
P7r0tKmuEGrq/JJ4MuueSlF3EAc3PanER+LIRcCZVRJwiwwPNBRDTeEVxOP+5j6o
HgMeqHNR0FGYbUyJYZI5K1SuAm2D8EwlntkFH6Im/YeVF35XYrVAGmhbixZ5kzvp
jUGcr24z6stB0Bs+NGopSbac1Ks4iLZn0uAiQ5PoTkc+7jDtJBAzIJD8ha6srllH
h5N00vtx0rKvDAmr7XE0zh583/o2iz9OhJc2EqrZSR/wrkFY1wgotOowpvO/IFUQ
5k+h4tLftm4NoChRU/7glBENTIEsybRFHGqOP8+5NYrxqfQrLhtKrAMwLc5Dneyy
+f4sZGv/vTmdJvJRxt/3J3/A01/2fYA3J7WNTq/HgYoqTgNKugusJuvJBIa+wWkM
6FCVNGf7yI2pUiiYECeElhZ9TWJNiiuRIMGBuz9FY7bf03q7h7Y2AHHrTqR9KmTp
1/NAWcF9P0mNqMGK6HjSVNpNvw2Nep565J8gQmE335WT/021CEf7jIVo+001U1az
5l81HL30OKgSVHDi43O8ltY67lcdvkzZfmxnmaLjfizVK+03uiC1DoT+kwy1/LQ1
7oxq9K64EIeSdnuEVyuPE2yJXyzy/HnmrTfVn34G97YuGqaFD/PJ1PAu6XZB7GNq
DRbyHmvF5kETLqrzRouY9FBjw5tL0BusZ2m+cRxYEReue+pixkkgIDQ6xYFJ5lca
uO+G/XiGiIoJ0pMqPFuIF5ExbSrkNMqhZh/57n9oROEF4KP0YgEiwEwu3nAaqQfE
nQOltT9oh6kYhqyajAVnclyhLZwFm/71JSDV3b5+E3qvCO6ddwHB9aRZ45GdLMIk
crgl2CHUCb2+78m6R3nZ2oHLJoX1Hpw7O8HDWtJzuuebP6za0zTw1Nu3rZuLj98Z
yohaBEWFN/0xJFHqEpzk3mB1MdLPtQS0lhd5DVzaiweljSiP9F11M9BmHb3eaK/c
nJSOkmRMOra7M8lGz4BtMl+JVwSh7+6En6MQxSfvo7nOTalDBdvcVv0nMg2o0MPk
VvzYRJQL1kaKPlCLU2NLDT9YsOPd3bTKR9Y18Y/GJCpftn3NycJWIyBRI3nfzKrV
WqvSYjr9oJhhqyR4Oe3nRUCSXLvSmhodp3sieqNVwuoxjcw3II09eGWu2J7k1ZP6
UaJdbtKpIQJUdfvrjjVFjjcGnl0IP0/HpjDChUE7RmOz89Lbcn4Dml4ONE+CgXFe
J4c+/VmfxJONsAjsdvVk+ayvRKlrGTFHGq5404u3t9ABLdBfYCJk5MOiYtOPjXBx
yt2Zm5w6XvbN6nh/3cJOASYMW4h09RpY4AnAZPQ3zeZICSapYrjR3jmmx9+10rES
hs727Mrd4fZDc2GANXJik0vltsddFnnzG16oiQu7RThQuARqzs4VUlikP8OFlFEJ
XEDx4a4xyblnwuesMnWf4PtLHr1NLs2ohvmT7rPo+g1S+Bb7Jw3muD/DsVIbol3P
Cn38YjfyrVXreju6HvUzK2RCtcOYOfXyITho1Sc8GpE8Rfzq+yY+bVhnjEZo4AzA
LS/YLCQyqLYte+lkXrq/j6r9oKcRRWf29A04N2M8jP2biQ+uZmsf2w4pRtzD96Kk
PUHiocl4GtjEa/Q0Cx5AFMtThrWVV+PBB7WT262uT1/2Bz4SOR96ICBhToaZKbHJ
VhY3EYElJoh8LIzgbnvYoh8Bw4RdIo2JtupIZm+qAm/cZjp5Cc9yEkEXeeJHJ1a4
XwgRrLl3tTz9J1wRLD9dwoFqsodAyVFRdEtvL9mqzgRxsvsdJciKbxXR68G0PNGZ
Ku1+1bIErULMtY0bYGYKBo24mYAg8U83MAi+WHa2p5Ky0gOCfBXHM/bvb/5MTvSo
TzOxi5bMuA3TXZ/lK6Xgfle0ZEj8lkbwFsDcReGqEpg1z8d9i4vVCgJrQMxQga1K
UYkR5EsOrFFTqxmQIDPi+pj+fwvbpZLTcxd7diX4QZyItDoFc8ItWERKpAiMqDFp
Y34SFqnbFdkneLPBfxsgnhSMS+hWQ1hAaDCv3iTc37uxwnkD5rQiw62jLt+K6y7I
wBlVK+3WWGkwzzLkzIqJBJah+T+qwdp88hOwu5rt73opmgyg3UIjV5exoPVmNgJf
xzZQT5f24sIc95jW8PXGkPSAPJO+hUM254QsFAH0hGrCY4b9SKdE/QhkZ/0FmuLy
ewZYwXhCQ6z/aAEvb/9rO3lzuN+xuG7ghWqNchH7jaah09sabEPL2256gjmMQQvM
z5T6KxuijGhmTOs1LWvzGvYPElK9tIcMuYQbisng4/rE5eywHEavT5W6H4BBleRE
01h8uWsyPwLSfhQaOkax5W4TvmAMdpFZ22hBIuwSyfzd03RjAdpHB49gmzMCz06r
JV2Rzo+LCHpjVLjJ4Ay/A4j4M0vSxBxwhgkmLb9Lja3bKzM3mBPDfIFRhy9qvzCH
sNcK84Go4hwl9Mt1Q67B3Y7KK/sz8eH710GKI7/8+5+WUpueCe8wpWv4o8BVXc9f
L5VvJ1nSsqxc8vSlnLoReUzLM06etF+95Xe/7YKJfJ23q3+WjW509A0vz3njhdU+
D9e6xUiXx2cDIir0/lpxMroRGSdHYVuU3YgoiDLVLM3RPwhI/mfE/7gBSGZ7hd1S
r+yj5yDo0Ba3DzUtgoc5ROVtQEJm1Rg2NvytH1+jcSmPCv/DbZsNrFy5yuu2B962
fohu3sAuNEEGM6tjIX9brmGzFBz67Bga9w3BFTyvh7zR6sFsotAlXm+bfqqr8r+r
Pn9NgSrhNqOyzr4GqrLe4RsBJ/RrpFhmZlcMMgizTmEd2MFIrIwmBQ+2MnxT0ZWu
DFovmKZMfF9+RTMJWu2TvotzOyVUUnI3TlF9qCZClUB4qM1CYDKGbD4Wl/OyJaVa
6m2ho5f4JAgiLEYXXt+H8D0XwROY/6h6wfnNruvccXCjDMzw5LAKpyFwHK/j420s
TH3c+cPVY/MScAXDmZds7wPZduOjXOqSWvH9+CYua+7iCRbzysYLEVoD6jpqgDhu
XApXkFcSbhtwlxZKqavSWMi64QmTR46MiPNuhIhaeEyr1A9MM5M6rgdH6xqiOtmc
pEhZyrwbtoOIuXLC/C+5ItqDoVPuTFu8iVaBFusEdUIPHn56QHhVXhxtySx2Y8yg
U607hUhQauEcTNa9cuIwiL09VjXhvRKmczMo0zaIzgpWW0QhICXg6zAM2lXGpl08
DjQ9JqEJ0V5bbwmzYUkWJyHYBHKIPgOexHZRheE0P+uxyRD0yGbQCVwacraXDWvV
h6shYXux2U/2RZZd4siaX6rRo/b33n8i5fT7NMv7ZFWfGVIkan8qbaPCq496czCD
zJRFxhk+dFpyddWWvYrV1A060r7lbZaz+FSrK08hKGblDvKhH/bvxY+iWLKmc/YF
91/Ev6rUjlVxNXrWWHO8iURB8AMjzEaTyRctKk46nrovYBr5XdUxO8bm5aP10t2r
g4+8wuSBVLIoAGZR1XHfHUxQObNgs6lEj4DtvHFOcl7CT9dEwwH1/epP94CKoRlW
1mMPcmekCiBPRua/FzAvNXQQAbig0BSnaL8w5EUG/o/JwHdU9DJIqTvwaamtTluo
/Wdxvc5e13LEk9fl98NB89xvbxkNWdlYN/t68yeJjuPS4tG60JSG14mVU+tPVepZ
QERgFKmIST+BW+h7EUc72OhPC33sd5s/t0ZUp+Vdp+7j7g7LLOG6nFCMSwtT90HC
wS3j0CYl0zHobFZy/mqivySkW5Zo0Y6oJewiwVOseN46GbKdvyO21jRwog9ZPev8
bk+1lhzF82H6rA85xs7gW7ByFNgFHtvIma8gprg781ebevQ3dO9354el2+D2ynhG
Bn0iDF9qOBkUeeSzW0gVKmutBBFw/zh15xZ7FckmZwOb0yQDJb+u/L9PwO9JvDGA
p4XySymHq2Ej9J2sUJbXeSj/HcEY4dMKyw29hbAnxdFFTl6urizOIzP6SU0Qxsll
zyXTfRukxQuia7w1wXT6GN2bmN6VZbZkgMmlE7pqyf4ILa+i/JoiTxLwo75U0lkx
jOkpkeK/ibt0bJ4fLM/hNtM+5Gnw/yca+KmF+rbpJPKC5SuXOQZQPrsa+5bbnmvx
Zv0cJ6lZzOLCUfV9SvwV4gLSLqPc4P2xf78/agle9YY/EyHk9Csm4okACsxf73Ph
7Z7klnAbV6+JDtI/WQBvdi9hGCt68RSD82cQPUej/Ask0FR1pvV9lQPDOIQSPHnC
YxBJ1lTwRP08D4yekLvSqK4YcLsx9yM4Kj97bOCI0dzTN0Jom9jB/w3a7vHkdSzM
lBEzWIFpjtnIsPM3TNOFBsZbTnjYLkzBmvj6ZnW2eyhDBnd7Q3VliHu6KrzXvD5B
QbW27cI2qe2Hlk/ROzVb0GJ4O+5DqfySfdz0iRU7LUWsc+UgwYGc+GMXayLChjJ1
YFxA3oT5UPA9jqf/5GBbHgpk8ch2JRFLu3380O38IVYjQvA1ewmfmPz9Lh4iDliq
gniCD+U+AZ04cki3QO9c29IfLBGk1ZFTK+QOnEoc6yAAymAJlyc6sNa/XBbcI8R8
SQnNPh5qzpZ6nBlPDoB5iQ/lHNp/+QJRuZrUOWKLQdUAWkmpypRNEy0A+s/OHN5E
BUIM7hbl1655gtdVZozzxAuXn1G37w6TFa7TimbwO3ho5QwSbsBUGjLoEk1cPYP6
3oTWBvOnBM8D03Ow6cJJkfkZvlDphUFnK0q5CKNZoFUxsG+DkmXUZRKjwq6PCgZb
yBKhPJ8r+5MSYG/8CbqXe0RFMoKZxEre8FpTf6c/9bE+O7P/sWK44sMcg+hba53u
09YvkaHSLqmlRzzTczc5KEVbY3snr8M83ZHvIQ8f72uRXbKHi+qZM2BKYQsV/2Af
Xvq4C+h3vp9EvPLJAps4CxegwTy92HBPeQUusfDVe88ipjngk7YwUUepwjFrfN7q
aS9l95VwQluMqKHWi/elJ/vqYJL8wPD2Ll0RIcPlOwvTZdn52LxH9EgqtkH8ChEL
HGUjFk1d0sJA+pg5v9rLPJh8obrSlwGLObVD0NzGnD1BTGrtIoGhysVlfKF9nukV
2RnW8O1DoCWocixIixUiCMdkAL0NtBhYkmb8hpQDhVY9yb/R0DiXNISsLo5UqdMc
yG2R9DrChfbLlKAHaikabve21da4lrGqvRkpAfkgeUI8rUpi1xIYM3wPsBOCfwdf
otaDf80pe5D3VvzJ31sN6QqozOtUFCmbvP5TMu8ywTTbue5InYsXWJft0FI4tscM
FR5e+kvCpunZZ5GSkbgpvqxj6xr1gHWT1vLb0hSSqEMFS84/FeD1H8/WohGVnCha
RAqH+CbUHxWJu8lf/CJmCJyzcJE43MQTAblR0T1YbgH+3Si4Jb+ut5eTaxSjFijV
JD8iBbIwJjTHERrpxDDcyKNpHBepnzZiRu72rzHnfKUuFFAY3LCc2rwgUV/B9Ix6
7+PFQEbex1rv7CS2BWE0uDePNSx/inynctJc/oC7oj3A3+ve1tCKYNA/oe8ohKD4
kPqDZEmRB/EPHgG1W9JSfXoMuFWjOCvLNPIv/Ww5U59qw2xuTVWJrjlWljFRirP/
DEcS4V4YYKiDZjCAfJEQkqSJl77Lupm3RcaAd7WHd39cyQU5cl01yRXtZAngBiFr
l46XL6Y0lRwCEXVYY+2LU/D/OqyBl8KnAfYsvEjGcxbAN11fDTOKIoc2QFO8R2WL
d2tW+8rpEe41hnayTtl3BR+KpZnnFJCgEPF3tGoj5XmjOSExIpwuNjyjxYb+Ldd9
6jthoSFL8C6zu5m2J4ugrAYOtlhB3E+FDEWuWnnoA2VOFVGTigga8Kc5q5wdjeZD
LlpyBL3c+F2JCSebp2jEVWbolUqLK20kP/oNKGNrzWQ3bhinDQx7lJ98ChLY2g3f
PCwRT/g4ixWYlXqzseJWHZVqZpFEDGSzWNpAaTkm4eIXiN4XCend7R8foOiGkMWC
oNbPYzq2AZDlpu47SNuhbqwB2O4UVciOAmJnXTi1cErkl1YOZCAG/X2VYY3uW/tG
ojChZPlF76GSGwGXofIJ+eBg6d29jSTvhiXrOOz+X97VxARUsvOe0N+V6YsrZ0PJ
S9GDd5yaAD+doF/s7ZCuJ9L2BjLMNkPewrrRS+B70kVI0jjjbLiKOnyoeRnE+TES
Sm2jp5cXv8Y/f9g3IprCHwar8BP+gbuBnRrCnXpyCRFT8Lu+GWnr2AfuvqeCY6uY
kX5RmegUvbs4Gpl4bfR50wYSqkECh3FyubmhN0uZ5NGNQ1w7gOOLLoZjgQlI+h45
T0jeNYSWh7M9RQL3mRfbDmpYq/g2XzYDiPq3zDd612aX+xTu6u8Rq4HQ6k8tmNwi
jPwnpPfi7m+EVDVzI8uqRXNFpz2vgqVkmaIdhJj86ZQrKggCMKgaaemATy1U6XWf
omOzxENnpMLIxMlVYFK/LlNfkv57DlAS7E8aXkx4NERzI66TEYKN+q7QJAfzrc7H
OvFHIkdgfMbTd3FoVA5pDr96T67Iih4+nttHoIAybRv2aAtEvpf/+xBHf2Dez7R+
B+DILYRYggZmaqocYekZ+2gup1+s3gvKAicoSOEyBYolk0YvpilY+CHSTrN+PN4b
KRLQF+UOkkH+naHMYrY9H+3/fIbB2GWgTZSai192WHf7E9TLk11pc4p4K4u85YHR
8s4qZgVy1EbDFseWKrPV+GKJYYbedXnjqKvXKYZgtYHrzJL5N8HbU0euVTP1OZ6Q
Z3zMCcIR/noynnqM/JylKOfo2lxJlEnlgxQ2RT6WJmd1mNujN38eFvbS3FWYG/P1
Beq7nBM0ZoLlRGqmHcYPFGuwUKG4uc+PqcfQBKntufaJqQt3zCTbRkZfwKeoMXMJ
epNt+pAuK0qqq3tFlWrbgFUXwO6VorCu/mJ/FaEuMW2ZiJAfX19CcovZkFBtx3ZZ
baXaeOx994eLjGNO36vlioSkbZO86s3s4ge5OgOthKAcmOFpSCvPc0gXxbPc2lss
f9q+mf4RvHBKb/9/vhhFGjT8KcC/qFBjFV3V6g3DelFk+c9UA13U6o4bV5NrQ8kG
7tjcywn231xXM3Ixtxf8Sgoh1dXQUn0r2x+HBHPwqj3MNQ3kcdA0utCSzuginaKA
O4k8VsEYttPFgdRta/W4+yTKYub1Aj2dq1LK9EZNAIvmv17+oMe2d57xTI6L2ixg
BxCrXhRm3l1k1RzjgKupgk1ldogdNwZfUMPoYGWdgeClkG7lUjxJoEDViV8c7Uga
RCBgMCD/d2K/wozCEtIhTm/M5c2hwTDUxjTNUDEvvUQUfkyc6yhXRwOa3+p79s1G
rqBiZ7D00KJ4blg6mbLhw44VLhuqS3zIQ8h0lLPkKvkdrBI+ZzU6iZLCINbEugle
QYU3rze03lS40Oyo01M+x3GJN6bZW/jamNqoyB1fKYw+2Nvnps/lwxims1LQyNAK
adTyKSHKt4H+RlXkx+KK9V7C4g5zP0jwISfdJNc4HtYToEW1JAWPv2Uo4QGSZzW6
0dEnWAxFP6s+EOyTjpYB4iVXalzswNDujY3MoW2XD6HLsuvLQrE+Lbcc/loRhk6E
sQEtbR9EIkWm7L9hVAdBI+h+Z14s2SBmvhkktkaiEnC1KDckvrvqW+0vJPm+Bxr+
zhgsVtPkm5RQe6jzPNU7/Dfpn34cPeUIz15Wxg//CvT1SLuXbut0aTf4KFjYBcLh
tkNd/aBM8iqcByK/J66ENIA5W+3FyWFkG9jbk6F8F3OAxaADVHp6M4jGL+O19vk8
fLALwnHdescpsUFQfnAjxTr6J1R6z+ygjh+x+OHjAcbuO9GLVo1UZemDqnz1UCoE
NOCijFk9eKY2zNtOc6I9Zn1l5tZPa3ee2lmNpzDivHRkJsg/IlrfsOpYCMwLo19o
TWMUifbl9DggcBOLKZc9iSXUhhso8fFJD8nu9X+CdlsKMkY+0IGgc3Drtj8wjPq1
6t4XIbkJD43cpvX2HpiE2xKYVOq/7iLGRdAmU1n1EoiIoY1J7zBNUlL5PoyDQu8W
s0z7Qou+kajrReiYzWmjg4XuXzvfyJ4IaJWV1KwUnEgkKZjqS2JfMO8lsYKFXgvd
HMxfyQyZPl2goLOWo79sqr+draMkAEL+Jz//kUc23fIHj1tkJvtfsYbeMLobOscX
0plTnmh17SogO35eSsmJCJ6iz3yheBdvkjBiycSi6sNVRQ7w1uGi72JbbbqlpU1W
/fPF6AqH4L09bFk7UkwwtCKn3Mv3JImzX1APpljCc0agvFBpxq9b4IwUPEJ3siaa
KAdSIJbvINo0DbVQqeToSZbqVhQv6ypPmZ2rkMPm7IyJSf3/GFIK8oHHZ7odkbom
h2/u0Db59H/Jm8E8RbQPLnTZ/mkUJV30VYlPw7kcrW9BWoJJOeDWU2ObNTYl2aK8
540ZxZ+LR13ILZV3bNoSAixpSXkdoieyOMMR1jYPT+IIQTDcQxhLLdzg5Daa2M1N
zCH7i9DwCIE0cXC7CaKaR3c4hBB+IXBwopIExIW65mkdaruDUSS622NophCMzFCG
E9gcAfq7xdACnyZuemfl9XKb4OpZqUZreO8jjfJtRmrsBj6+ceeku0oDiJogXFlb
MOL3gR0TzTrZGv/9kORPsAp6qt+tRgW2mSXJR7rhAyjXhsF/2ipvgSbnaWLLpSxg
AZzfGfnkWMBRnPzb5U4yxKDHz8G0hE67CRWuWMKpYJHcGFFGUdVZF40U1ryK2E2D
hCYWVnE7NGyC8KME0Q/NfdokeMGFfoQiEXmFyi5KPcTcvaO5XgmXe1cjIj67lNyw
Ckh5iVgrXdPsbuHJwBYA7oCXGcBSNpuNlg8tGpwhZMqZu5ZvQVIvvKGRZvYWbQ2g
csUPpJyjdsw4S9bnBbWDLNhvL9/cWRQqvPmJnnVqE+fBK3j7wxAdLDnc9z9lzskU
EQUpsIippAgzuCX017MEcbNtLBjHBo5EJABulJJ8y7cEUvlJQKahGs90SAoxExdS
TgNMQELTXRzwkLkVQScIVPsQ2H2eUVzQviQNCdL6bJegP+9Ad0UHvV0WOVwfJnDH
byujV6EYA9i/VHwuXPO4XJdsbrg0rsl1fWWGWcAoB7f+/a3TBbHp92YhTmXuXF7L
20UoGwo8VB/n0FH4DeCKoZ+fDT6mYFef2risREAnMyFrcibEYFegKIp8jCF600tH
np7hltqa+e+apyYEg8gFtWz+T5pIWNI/UeD+dM/dfxsIRLJePqplrxO0EUIb8mdw
V0M96gULH7d7HAm2hyi2EHeOldwq7E3lfNhifwaHUtwVab3TGz1zmoVZzupnCl1F
vWZOwqz8ab4WZolO51ADEkDblaYekx2TBZjFC91Kc+9N1XlsZ3nP8SNnik8Kh296
+WbC70Jc93X6f1ENTOWeSOIdYfuH7gNTNlwgc5gidpJGKiFIQPVAm75sHUgCr8iD
HrADhKc1nXYaPe8DK3TQAmI8XeAfJkQ6axvEDRtWdQunjmTYDv1TltZdCWZOW34G
cRBfZEoFaXaBNxptflLkM3ogWA+gkUveE7nJ5PLWJfzmeci3wUgfS5zg6SzgrW4k
gMFYcRYcfRK1aGvCS7SfZ6pG6qrVT0DEp8LwWb1JVxRry63FYUibigKQC96lreIs
NgXeWaqQhmDg2K8czB7+JHxgXvRqqZeriKKmKJwPGFwOCvAmgHH/1lrF87f1qgFa
RJv4EPh2DMn3K73YQLzzjB3GcH0AKGkmrom2pRyr+8od1L509eNXommJZYfo2WQq
mn+6qSmKpGHRPg6Tc4JZQ0Qt5my6aIPgG9CdEZOAwrIjcX2iFelbs5crNhSZ8zMe
2TQnri+CRxR3s8pqlRGvci1x5tRKPZiWU39mT+CdkEEaHKq4/g4SAzWjVZJgiZ45
r4rhVToWrEqTA4ettMuCTA4WXblbfp3+bUaQuMLlV4OSKy0h5UwbYgfomGzQrMIn
Iej/Tq0N+OR0DcsuGGrEo41wyAgpsYCt9LbVxHyTyHqAcDD14itEdLDtj/CktmfN
RQ5Uj9whja5OWPTufhn5oIa/Ni9oYIysn70DD90o/dWM2/REPX/jB+mQmgBfitS9
enjuwrucOUujGT6uS3MsF8fGGAuXcDk2fcALogyPlLJK4UazUho77z8ImiZWwQNi
gMzp5zr7VLfF69G1a15BG/5/DtvzjK/bgZN8oHOR063CO+G3W/fQ/j7gL496Dpn4
VydOeGtOsNpM3cl2EeMjFirDfO5sjY/yI45E6+NjPU/Qf1dFFo5UJoUiEAgAWfTh
Yhq3nZpm/1CzE8wCut44u/dgXYyG+PryOeoLNTPSo5sYBe3aV2UPMOXuBZ0vT0yq
SfvkeW3zc6EYRe0OXmtH7NrC/7RrCQhoWQFp1i6otmrCjfsciwBJbDbjnw8lOz4U
7eTVYsv9ldtTVFJd0sNhlO66SMhJn1mNv786vuuSk0iVcvcRs15NCNN5O72moUNI
oNuPWiYuXeHyI7gmOTmJ7njB3ZzPVGOuHNXwaF8e38D1Txbho3A5oyJGXrDot4Yj
iadZqssI/o+0Lv7bJaaHsC6ejQ6hJRshEfeNH6rAf59RLK+2yXW0C3KgeuL4R2Xh
C5l8k3N/7zc/T4EETE+1IjW7afA/7gjAes9sCwUfSYe20/QzP5+8O5pvBlZgGlzr
d2/hw+2lo2i64Nx4hYoypOHKunyfAC5+g6jQn3ePqRF2czWaCZX3aCBUjMv8oMVb
nTv3AVUtcqycdanp34bvPWqjTk9ZzSCN0ybis59bFPXv7p9U4vC/DWEesoGAps2+
4QTmn0gsiAi0NgycI3TKpGKyDTYbrJb+M4Jn8IvUSS2GlCuPU/V9Hi3k9asMgxcv
Wxq6fGuNxIyBpNZEfnHdM+1c2lK/uqyI+N2dKrFB/4y+Pk/aPxZvV43Sm0x/Dj6U
o0ekzYKS7O0RQlqG65sWUNnjNtQ3jyBfQQ1kbq3U2OXqcrWzvYw1Y7SFv9La3ypD
jIn0A9JQE52hUxwWxSXiHSoGRutb41fF/zguVSGWZsxDjRObt/PUFEGd9Fek/Ypk
vA4zfT2aoMz6t0rLLfhHj49IXjwZZkkKShesBIFYsaoVUzBHcUE/eqrv1ha3SYGz
cxMdCklAJJAXMhimEEQdj4oJF34tqtODRCcxB7Wp+Nn/nOpa1RhKLXBzET+dpJyn
YpljhUdqZBrf4qE9Pd8oCJKiuGltK3j18KvdNF0GSjneY4Yv2NIZe+wVTLVpBTU7
g0oBIFzxA3EPxRP69jd38adGSuiFv1u6P26txNCdufqj29/lNgd1ahJWExXM94yy
4PPJPdBCn0ZQNxZyccgdMKOFX9edaK4rPcGkR34GkAqyoETf4WcExn8uXt4H+dhk
1dITf5dkuFAeYIc70ISuKBH/zb5HEaPWZZHyS+wHbuiLkcMDSERlXJdXLDoCfsfc
kSntpBAkRgPYt102WMlvgI3bm1YCjfbSRfwsUiXOKFGJw0/M0ENir//lHCRv6F3g
eZq9CtvZ7igvVz1yY5toqmtdlpkXMhcP9nY7xRx01kDomgItYADPC5EuUhPe9fvj
mZPzxxiioKGTkniBRdvBRf0NAtzSe3KC4IUvcFEC5W+Pncq/U1iChAZXEJVllH4/
JhEMI4D1d+rsglmfRZl5w5782iFB15Y6pogDUUYdlXK70Bt+b09vfxJH23+b09zp
sTU6Ltww1xGim3vhIYz7s9hI99qTmOvv3yBgVPO8ACR3t1P3A/bDXQC6klUV0KjN
07zct9gs5x9e5JqxC+H7keSeNCx12i5es5PQh2G/Zn4UOxspR27hQ+xGdPLbkhM+
cG4TE0NXRMPgBcRX/6X8o+0cEXGgRKgM6+CF7qehHLJLF/YgYl8PhrEYYUR94aQ3
8DrF4VEbN04k7XxMpsD4GSTuG14sVJkDviQcTKqlwc76Lgh31sVLJS9rhxlzVriN
LxnzfKSehrHv3vODj/mAxyuO+4JzJYrBZ58Jp8GUjypJ/XPVYbsAIcMQIPtEJZ+0
cj95hhTF7hmyv4qdVOn1NqZvc3Wx8dTsa3kBtvpRHeZ7PytwmIEM00jfbBXlezLk
kBpXqZ7retlw9NRy5y0nzlAAAos/5G4g8zesTpH0JK258UVOa8mkUgT//GKgbsbR
T5ta6jgBxDbggYHfFQ8oZEFZMaIbOcZcFBcHDXb3ainRN/MDJDKg1wgTsprhkkv3
UAH7otVmam0uwatSpf93Sxbhp4V7GH0q5F2Yn7Uwvt6XS2gMLvskpxUbEIl64muE
/Au0S8TIizKAEFImuN8RdT/Wb9fZjHYIKzdx/uWo5sXfj4qwQe/uvEDl8zFRC6/4
pFb5LZCPPzCFSIGUoLjZEn7hEidVXkm7orKzdbvKZu8hDNbz4uyZLpQHSMxPirhW
hCE2PGHyids9XBAfP85aD5F1niuHVvqqs36EOF8Mpt3LzbAVvG7jRigxv051/aVq
paxllmm/k+zcRwoLiFMkNE7yt/2BQw1Zq0BBUnSrXnWPq6EGP0PXVQWzrxs/4ewP
fPoXVbl7MOMvgeMGeRV8ORaKWPXmBIYMYIHlwNNNlrDXB8oZ3iDC46PxwiorIYtO
th7MJbzTyw/leWMaUO1O4cax5Xtzy6VqJeyKNQxb5RJAd67Lwp8US8tUWqAsnXcC
1c6NYbDN/Oo0o1IV2w8z+bb05TmPFC5b2/rvJNYm11R/1+39MP/qlc5tahzVXMTk
Q7Mmhjx0K98uxF0+De3zy2H/GCqbdwAPgNssT6SqwoUUpYUSKrsD3oSQp5cnaK4x
ZU1kHP+WI529irsjoTaYfcqyfut1Wm6KVaKBtZ2eeZgXGiUaIjCL+Ahtb2XLjvLX
EZFBD4TsH+Zk/mmu9A3VlmzUxxOX0Mjr0lHUxZgk0S9w5qTZ/fzlgjyrlA60Btp8
e15xS/JIGCTt2WGS2YgQfn53qZbygylxvT0MDCWg3EYH0FJUUIUBygz+dGx9qtDV
N2fWw9Snrwd7PjjPND7gJmHZ3fD37K3lECHR3NJlSHtdTCk2tIK4lFtpDuvvorOr
aoxWI3ch63PkMR4cxNkdnw80dXHBFpBH9lGqhIV1eDzeYr06gSBqdpcLzzX4MNvy
qajzngMrBFTsDzQUo3aTWeAS1/q86RXtt1uM5hr9ONizfljuqpvskuAVR41OGXgb
Io9Myz7M/ttxBi+AFnaORNPRTwWI0apY57LXWx6mg33/lrxAt8dnXZ5XtetxgkjU
tnQo/dG5lQToYWvJEz29nQpQurrUGwbwozVvalHYJHkmyPKanMi6fpB30RexQHM7
aiMEWa9iUNbKoewFZT0IujPCEDjKfwfAYGa+XXLxXBr9/YNQ0RqyrH4nBFZjjl1Q
jW00xJsh60YDlN2AtVu0izjngR4wdCjuYkgMJkK7Izk3mS+volouBrOJXO6DilrP
38x9VKTxNtZiywi9oqj/Lw6UyihiaqTwKYMfG7T8pEvwuOWz+amHDJpEBtaS407u
VglBz73zNid3iRtNRlo8lwrUzLLOBlf2pxl4xof/Gto+SzpRcXZVwDbZTVc7sRJX
4IkByMOFBY1KQ10SiIA5owp+UW8eermadBEI3+s+inbG4iGtBAd58xFwl6dERftm
ieZmVTK13sThS93z2kqCvMQkN6HMqZ3jVluiobloOjGa11Z+whSnY00WuRwCEl0Q
G1If1Jrhp0zGrzkBef0xsShOpMlBZ0Qisp8ert8QdgmYid1tYFuC636T/0i/kI6s
EX13BsUKS2TDh8SEjOwH6EtbzJN0nf9YIsNqVQJApAAUIMhOz13oZ/ua0UNBF4eF
rx1JQpmYb+VMC6wirUKoQosEWJn+nOYBmYDDHQFQLUlXL98jU6/TEyxqlOeEQeN4
5LeR4IrvdS/VNeZ+3P8eNxy6zp0B4VFdRa+Oyyk+YKsm5euibJlFXLRtzP2min22
vCU297SZ5mDq10oSoHbyboqv3PfZuH5tpljlSXfVqP9TTHowWrBf3z1OTc7GpqQP
cIZhnxFwaF5yz1nbxHhNrL+YVPr1rs8fuac8gp8EejnfCYqsGpC6REjLNE5cs3Ju
vVWwTJAt9buVDimDsHLXJqnH/JRZmF5YZY3HMmezVO0w2+N/HbB98N/dZbt9OsM9
lTLkYh3ObGUOrZCac26rE9r7Doofw7rC8hCQl3hx2Sr2Awoi1auTZcjpTaWpHgtf
7xs235Bz2uygxH4tENHlZv1tSxfJIxzqvepl//8rYgkGEmaP3ti8W8e5SODkdQvd
6TXvAfxiYetr5tV4K8h2hN/jPOiJyYZtR/lSO+3VszamYJwjhnjzhihb4WUGtynS
CxTeWxi6R3irNdOcgKAj9sfGT3kYHLJE2JvLT+L3KylRrNxK6YsQQytYISxq5QJ5
+7dppf73VDn7uXKWKFheLkBAmmHftKpTYR4iqHA3PKIGOj3zmR+Mko/p//YHFqnb
a6k5Te6hdjYIcrVBBYLX1dudZoGd15qnFpgG60LELrXKhw7SXrjr/Cop2vZFB+KB
RkHFW51YhRjFQf7WfPFz7U81UC6V2zE8rYz6Cc4gKkGzGRwwkqdVb6A26UGpxHKs
HUirFpIHfB9PJ8ne6nEu3q9AkdG1cSU4d5cXD09Bc0Ws6iNC7UdoZcobtbia9eWd
osDwAMANiaQDhWE3l0BAM1xMM3BWcwSf15u8rzziR7KuRmxtubhVVrCiisQuoPaq
2Pjkkkt0YE5FVIataSjbhbZoVbB4HzYgHjLJ7gEsxnOvTshyDIkK/Kz2xrRqe2xP
bS6cM+UuuJUmK+a/IAAqM5lNxIMXrLVVfkBb+KeWKFzpCn3MiKDB5kKFp6QAobtO
kPaDn9+FqhiJGfgmjJ9zqkDNAkiSR9F/Ib4o2/jgL/WawtJabQ/NfShc06DbzPX+
HKfQmcLUZLREWk6K3h9rnLJGDyQBkl4SvKd+d2CQcbyUDOT5XEduNzu6S2fKwXwG
d9Ef6uVdccasOj5pVS5UoeA3sHCc27yS3upe4lTKlxWKRDh43QVbMOx7G78QP/+a
2nkxejKG6Hbw5Lh70Be9m6KtpHUtjVKfLikTxFIDxRHa8EBkW+Gf/jCcVV+wiYBQ
BVy9EueUqzr5+faShI616xk9ztvBmq9IW9Yx0nLPF1TJjoNA/v0vVMoDU43TqyWp
z8oqDq4sBK+7YMW1uFGWWvG3f4kEHzMmyoxOrgnWSa7scN0XIh1wA9vG9zBBzCjs
6eaYiM4zUi7U5pMzxM3YVK9k1c1m4VPADE/GTb51gk+ywHciXw1Yq4thLLE4qWFO
knT0W6kWXijFe0SQr4D1qyWJsyi0WKmXn2bkRvBM+r3bowdqLJcpBhxna8z0qrbM
GBXVrEkDWS5JCJtUrjJsGBX13xZC0c3Ntu/gqJDUogBhAEvCH/isjrB4pNiM8E/G
M2YRj6XSDU9ItpBueW1L9BF5mFBuYjHCmPcDuB3Q3lp4GiWpbtzL0h9RCa89d5OS
RKMQllnXcUCbmB2ib8Shf7aamG+QQm/pCJ1Ei2koVUHdlJEjbBC/NeRktzgoJS/g
Nh4YS/z4GX23Btr6oXQLpz/eA9ekHG98DaCO23tWkAzujfN47JrcDeouZqxp8R5S
k7K1AX89uDfovozAjLAfA/Y2/N+y7X4OcsH8+vtYxmnEy50jZmwnEQJzVCndEtKu
PzOjuTDYjzbFfgzWErCz37JnqxucwyM49/+dKV5WwMQ3n6V3sn+2T55z6OT4Hh85
EJ02AIHc7Wi0Whx2ArrHWrKik0bkNviAUXDjkT6OIpaVM+mGBhwp7dmL20BqB7vH
1TzxxUCV/Wpy+V2agBKzIusi7kbji15t/6ms2iAhHLD7IVjh3zqfgtCK21HsyTVp
s3UFAmyIO6YnH4EvfkrmsWdw5R86e0wsdn546SARtpvhsIaLPvack0lMMQCtmrk+
LRM1PvPGhEeDNFPgj0JWnQQ+ORvk1lvyKDDclu9Ys8gLabdeld9hd/fj21zon/QN
iUwTHj2EenXOkFNW9exsxgwd3buq3UFF9rC8y33V1/uYiNunl/OKHpLBOqs3/I9m
d42Mtj5yizES0lwiqYcBGbVilYtGWo+OH/MiKJ+hj1SxlPaHtxd5h8TvgNdsl2pF
D/ldDkxF/jgON95wzlAHx45QIvkVLFBaFdNrQ4o07hZwP8Hq60nZCa3EnF9/Mvii
A8/NWwSgw8UItj5H38Be8oFM9oDMGivcHpN4NQUlxJ/u7HVvG8kf1U+5Y+MLhByx
4Hgxd4XNKmMtWXLuu5C9/m8w+oY1GLbrPf93BXCvcC2wT/aUk3cINGofGRzhCUpc
YzvTLhgR8nDfsUUopmgjEjMqA5Qag4/ulqjruEl4GMQq58eqiKFLtMDSMUWg3Gj3
ay0x2OEMz8LNDM/Y0xsjVI1wm/9bngEKCh6ucRjFoJoK/wDDjEiWvWwVFtXCLgJP
eFow8p7vxZY62MGwXRbpESzAoEo68MRwceUYSwvny53/HHzNv/DacvkqoH72Ugze
YG994asMXN7TL+qlSpdykJ8SK3q1sR6rxXTMTYJoG1el0tf6wlr5909qlVwtdxQ4
K73qAuntGq5ZSAg7Jt/fQnyC30nI1VVIX2kqgMHyo5Umr2qEeriDd/1fVQ5eXD7J
MCxUSjFJeyPDUud4llwVlmg/9eqgm8BD7GfW1hhP0irWJCM/MUkTLX32Vrhxy278
MTLqJ5oR94pH1DnMy9PZgo2ldLAkifcF4VsOLaypoQpIcgkDvVRj5TONjCL+tezO
TGG/UXFsboAxuJxBRPCdB5URHcJoXsNSLOx0VmXJLJmOA0C1kcHeX//hkGDcwtwJ
d9BVbGdomos6Z1t5o3gsp54S7yqqDcZHZetDpjlyyxgSJHz6IyVJD3MLaSciA0er
9nDs8WlxG/ICNcJQ1iSum28xRgifNKfitdimfvDcd7ThPBohQqIMV9izwF0Hmay4
2vK/GzYOe0U7FsAsjTwKr68kPSTG6cpeIbaEp04sVzrXRbI0SWf6gvT1Qc4CZ+gn
3or3veVplWD0ZP/0zlhvM5Y8f+J2sLvF/0zUzNZPAOUdGZHGrJypNwHxD0cPmSl7
6uiT9+NNMxBoiamtJk064SePjqPL3GfMiyY6DVTNyi1zxpu+Gt+LWX3h1OKUZmMk
Bex0Mrr9BEJONe1tUUEkYedIsHAYaY38/SsPXugPVrephzOk6mFnBnXcdtJLUdNT
zodTciqT3QZMBAQT2dsBXAeAeBFTs8u1ooDIghYTlZtDy0MiZ15wVcN9oI0TyODa
E7HTCaN5yJMcDeYCNdkFoTIEB1KaF4Y8THUmfprPKg+du0989GXViQny9z6hqKuG
3qo/GQ9VVHYNrRUrh3CDg55+PiXhVQXAJkSXOIQ1799ZZr4ieTcC24vtZ5KnAlIw
Pwbe7Qg8i6P+A8R2jrAnTJotVd0aCz09TtV7/JAxW0eC0y4PxIqyZziWaLb46d4+
IhUeIU26qG9Cq0VJvhh22eooaTLoYLAPKrqpR4bxyQYqc6g65ytP/USDWhIRKdYR
IwoxkTQKonNh3U/ESu1hV/ounaUUgynO5ZnfIqa1fQAIaaI+V1A2W0Y3P71kqCU3
F4nwKAImIZWbWL+gCibeYsXtIySLYoV1Z5ldvUUWE012Y92KFBmKFdpq433cEnin
NYV1qTQXQtc2noAD9D+rqLPlNcJcsA3VhTTdxwOubxNe96mX4SomvVqaIwfQJLSM
WM0kV0I6/ZjiqLaONQC0vEkB5jVArFZu9Zefs7PPOIdQ0GD0EpSYKnUYMq5RlsNK
VG5RUr9OximU8miP5iAXbTsPTOA7g1soQ2iIMaNCCKA+FJBOmw3jp4bJ4gOlUuLo
dOJoaeH9kmjU3tbMK/hKnAQMr59MuFiOUSckeoHYqs85vJcGbUO1stMb/UItKeBe
Gtu0FDfgq5SQ7biQcEYE6TWwWzX8ZBB+BbtWomzzCAV6cd1ye59v1S2zcU/+gpso
ZylXbBeT/FqQfJkAPsYdfkG/bQhWV8LbziHOO899aoHBlUwVvVMIHJewLfkAm9so
/54wX7J3zk324rFz0ggVbxqkNr/BnFwJ5xaNmabGJnfuJraY9gGzWWIaddKmmev9
k/ER7QW1JTvRqt9IDvW86sWxSbYwCaGEFKKNFhqJ/QqYftpn8BBqQb43g7OZ294s
iMbmngd9bmPeeRH+LvCSqOuvHzNE75sTfV9FCYRHmCAkfShhuEuQDidUQiQpiQPv
zWKxRzTR/HpAlasyr9gaYyVaawxNa4Bqe8G6gdOVCUmfSe1x6p9tvDh+9nlz+cYp
qFUJCdobPdj2KE9mPhjqV29oNC+lwY6dqfFDN4dxIXkdkUJG2pkWcrli1arKwcVT
JqUj6Ehe5KyLdZrUSMUJuIzCb/pnIeKLXu5t5A57E3HBXCj+zAxpBKhd0iP29gLW
WlrqvhmouQ4ZwcgS3mb0nau5/i+6t3IJle0rQWsy0oVSpLbe3Cnorn8R05/qOpww
gax+jteNh+Wly4zMOmwbo5gKamOoklAh5FiDMF4FzEG+np7iTAmnOYWHWxv72dR+
EO/qkceHFoZS+alxhUhXAyAyKl1jADRnb5xjSn6j3U0UNH1PpcmrOGDupqxvcvvs
3P2p/3unhKAfSp8FsOcVG9nxjizwzFChLwvH2vjCzFoQ2c4wrkZWwdItkgWrM9Ft
A5JmmTKcrlBtDSqxzCLDKvoazZMVoyg8JvHssZ7iOi/xN82jclSVFWCJmox7amQb
t9/dekyl85gKRTbPmsNgPW00YiX36pDgqZ8h8uhinEB5qAS5PMUHfZKvlZROG6WY
WaZU+1QsTO08hGxOzgf/HaXzbfnukOjXN8qNHTUia/0Ui0jmMK5gyLf+O2/Ur93O
xDsQJz3n9+ikfWzek8ezw3pZJ3dZ15Jgd2RE162UeX3QeE7dygdc+jNtKW9FQMnM
Q8h9PNBrzKLOHfrcENjIbU+eM1m78ELtDivaz980Q7DaYFhT13/57ah4sCOda/Oz
yV5VxZcd2sCdfYnBlsi6HroB1XQenUI0Btt1DNO8knynCxB5YiMnY5pTGpE8CRvi
uh0wkxhvZ87g+Fj4BamFAkM3wCSnEk0COK3Rzicn8RNmCFYaWHO2KvpQLq71Bxk1
Uw4Aus8SpS14ly9cLvdjbDQYN1Z4dNYjBpbjXxQwu44I1YO6BKkuIGoGaHlRwENy
q9Bw5gzsUz+SxPI0ds6Mk+ncr4QJJNNrlPqT1XLpWMo9dhTewv+SVh+0Nul/L3Dh
stHY3TXA/JT+PYcScWN2ipyfQNaAcqDl9GZZoRq/qCFFb+clUoG10rdr8niNIu+m
WzagWNHAQSK4NwAAG7vmEtkux6p8vF4Ziksdf8yxS2lL7ZZ36Z46ujXo2bMKm0Lb
lC4hMzgehtjh1jo10t8qSQWxdIUiImWnuYm6iaBwgTM+bftvNRy/Xzr5aqzbNtYZ
6hQsKzHejHvnVN2j4FrVu64NRksTmcpcoWPqaL7gZ6A/nD7VlEyMPHrcD/eRj5Z4
0VPqka73BUdat/pMPJG9MukGqBCgR07DKH8lHe1Lh26vuJQ1JozAkHse4MpDZdqR
+bVIsLrKWELEQt3OA/2gPyPLXCCE75f/6I8CgmKaAahJxV9SuUnr5JpPAdMzrvX6
CH4nr95VLsLTjswft6rK3LCOw+fHfo/Pf3Yqpbr8mKdGdgIaZrVu4NTRtVnTpD+l
CZJW25lhZntkBD6mZF/2DV1VbHOpzovMpjiYDviKXLsvJr6DMUhoL4fK12RgveqY
5rULntEGxj7byengwICyhHCWs2dp19XT9gTlt8jyrkxX24c1yElAfQ0RUKN5dNjg
a3QwSdopBsXDZ7c8giceFqz7fWcwe4Tv/ceb6/y0Wz9IFwKRuh3Jl/W8lYhGFmBO
0ktl+qBf/4q4NoI/Ctjla4v8kxyiePwdle4mjUkckIBAU2XBgWHB1CY/RsGIuCBJ
s9QE46YXz1r+PE/yuiryYa8Alt/h8N4IGwQZHt03BEu3vSWBMvLJEkBJ633mS8p8
8OsEJOsjmaSSqGZ3WaR11JSF8LFZGxQTo/KhXVQYtHT51KGAdh9L7vyTyc+xRLLg
80y5Ky9ImylRq267lXU0VHjqH2mg5biNyQmtIxcoqLYqmhUGzJPfE+GdiMdw41kA
LmMXYKKMhArU0/0A1budPlVTy6d+KmITcvzgxqpdAEBxttSgRxTQTlsBBOun2CM7
QSC6eEV1WySd2sdpNdHL4DaBnYxhqZe3aDpQ27en3sMDG9pqZD8cV2BGlR5ZnADM
ABN6QuFdLfBYxN7585Sw+miSHmd1KdFVymKul2voK9NI7qntHaRMFqWOmnHy4DuS
rkG63IPuLgaCk7lAx2U8nNX6rIQOdkZI9bz6iLs4kvMKN3xOL35fCl1tBhPSOJbE
yunbMP/UoM83xMbt2LrCm9eq7q9hXOMhaU09MtvYTU0t1OhgaF81iVy3NI69K3/Q
4xmXN7cDxvyYImy9sMHboQYnlJqjPJTfoyOergVlI/Ots1wiRl8sGwCuhGET+rjM
/2rghyTLE3E6LOo5nMWuYQ2v692uwcNysACMofkq3Wbs+1V3Bd9HGlN7XjKUv4kV
wVYEvjePibaCAiOIE94ShVm6wHBHVCmbElYT4mc0vjU3Xd5jTu98hi3PQT7HjJ/p
1dp+4zoF/rGozRw5tGWqpJjQiNRMAVb1PI4wz6ExjTgJl+4wqxLgl3cxU2drcahB
iw13y6tTaUpsdeC8BrT+cqSAfCpAgOnNJa/IEH8eKq9v3+OwKGxeEAREGLMrB/Ac
6qm5QhuNOdzmiVoTdbz07/WCAMI0AZ0XCn0X7/xbneEsmrEe+RwbJs8cLS3tMpPC
6ygfxL3g+spAR859WYlgRqrMRFhezB0IkXrg3Rul4PHWB+9ypAbg5y4wFoMF70Mw
h9aFHnLOir8NTL9zJ7jhYyzGwixfm8adDTvJpdDKMOq2vMqzlnO6tlmiotgVdhIq
zlihtZ87GrKT0x95y4oQW4TDmimuYXZT6XxaQrPf/jqWjdzjA8YENqER3cl0vgGK
nUJmWsr5U4HJZg8scxDk8y9X8nhDrhnupA2vAVjK656bn9m6Fq45BUj8bzlUvIUg
qctq4OnrQSAhfUwY2xpSs/I7N8/BrLkcdj3u5EhX8moXJrYEiMk1JpZnz6ZtBRKm
OOVDrMTeO013vRZ2lsVBGLOTOYQxa2bi592eZf2cOe/rhumBwbTucIvBhYH+f2wz
RG3XIjgj+6oZL0XF2/3lV/dQJDHYM6ywLwXmjXwLwusfL2bh9ZcUe4K1iFD/TDnf
vtt+TMJa/eZrm1+qKAqotNW+x44XW7AUxJ2T4fGZVvg5x5h7jV/vwqcIHhuO9rvv
9+ZKNSnkvxoU21F1HtzEvQ1PAZvu/XRp6z0dNfL7Y0ckFt1Ti6WRTAIVb33tImnI
l6ljvcnpdHtjGxjGJuHqQ1Y32UcIMoELd+bGMsa6VZcNW2+a9hWHG8KWfQklW9Ut
9+cbJ2pO1v5g05tOsob4JYQft3DvoTkXf1GWpP2x25uBYJ1mDSBsASRYZPAIILDz
/KGMEEnoAO/wTrmqPlxejbhhuLoDNnKdv9JL28z9LTa87Wwd12l0yE3KZCfoH1mA
EqVweAa8JzxJR2KYQDWpycsDc1p7i4EDlnWr6aBKN3KNfUfSfT+eU9r070FFP3gI
oH0Tt+8hUa4pcbXZo1iJ2B86gx0PZJnXJLnQLWpdBn5QFKeePPS1EUJDaOQ9DPOF
J8bdojv7rtoOSQhYnWNPB6dWXa85fP3QYjmALtk5wQudMc1EVKu+jIqNHjnl3uez
5tzbev4QOZ90rTyNcakMN8a4o/ptBLbfwamAkOLQl1XBp8N0ww1hEEGPscOQts8/
ZabXo+yuqZGAixkySwb5idOaPG2O0KdG+17PkyA3ero5c2O4CAbu76RsXvaFlZCE
cPd8c3neo0LFybXy3EU3SefhueMi8+Su9XICHIsMHjcTvOHy3tDVn7UOCULDpbWr
QZ3oD/jDS1xmcK2be8bpASVPWXpMJHqmcu120UfI/5c6pyKrlfZ8mewWE5Oc1MGj
qaC6zO3OouXqq2M5I2hxm7KNmkvnclKE4Shi2dTqICvM3xX223YQbBBqGzLqW5CZ
KgYx4u6EIxECAVHMfFme8koT3LWtstZFndd38tkgPJ1nVt9Su0hnbn2HuLlq0Hlr
6DRifZAs6E8bEc9GzIu4MLGez8AoIeQBFEjd8sIddGkrcL+1MZmleQqsZxBgDbzp
oQLvPaDpbklhdN+kQkm1ZDT8vF93H5LC38jFFcUtHO/hb/t8nD3wkzAnbkegFP5u
5FRf+t5ih0aQyDEpDh108G07X3P+Y6kRrUGYrv+nyBGbIJf07WeJauwXfhAEpkZa
YAdsEUcypYBjdzC34uwFRltSUatG6cW/qciH7UTePK6IVuymgEmIWT7Co+y825kr
AO1Bx4CF/88p8r+g0qT+OZRruBdsaRG7F/ZgAkw3o0N1nzkZIT7tfMN12FoI5saQ
z62aM9lmFmOHXJxoXrgvb+O9vzm0Zn+iVajfj3RMU5Vi5Fb7brSan+LgfKkQoHzN
qcjVbN3csAbHa2iMVGfX98FPbmTiMZJGK52v9FZ4rJ2NJ71VheBL7bIjcdXXZbR9
C70KtoLsHG1WZDcNwFLhI4d9pQ14iWhbOzRuvR4X2zQp08C4dmPaLM4sq4jZK06b
RpqWK3d67RO1aq1WLGue/qAEe0HkFOHX19XuIymlFtTVHMzDiDRLwTWjpz0tafUv
Jht8C1PG4BjMuJt7L/Wd/r61C12vzkk8IdKspzMafiuv2Xm6vdS3SJcSQ/F4HMJU
KoLNSSc8skQ3NUCO6KzRinEnv6IdzNlNumBCi65aPc/jqj8L6eYDZ3EFUiIqZunR
o1fJ486xoiQCB9ChubFOK+A/xybqpQc2KdRk09WSTTNrQWAziS6mDhGGdbpKYJj4
kjXUvpRLGfFo1ih7b6JVwxhHhXg3SLrJF1eurQ+I+R/lQ6W/e45GI4I2+aILjm5X
sgCAXGPvDQguZB1jqeMe1qn0z4tYmFrXngD3Hl3obc/LX8Rby9Jce/B2mDfp6XyL
7QJPRkYJL1OsW6H3lkSCWZX8oVypmPRbMEfobeiV9kRWEnd3Xw7gWXTVGpCQZ8Yz
D29d2SoT54a5O8A38Z9HwLuvEymoeyB7GOrwUtL0pwQkXXLZpVt/j2bqg6LPuZuY
4/Kprfu19T3N3IqB/dirh/k3+N11RJkdkC816C1dQ9/Dmc54IGfA0ZKbkxDBogUc
NiSoxysTcwYkVrxXWpcvE0NdhifjG9Q+6I60xnUtAD4kYG0QOoudARvcNkOXzgCD
myIwH56R7bcUWVaMYjljCUA0R2KVora0IsrJg77fou7zv8Y2ZlKKx0qI5/cCs0i7
5E/bSI7AsfDq6ZcUDGKmno1DxN2Z5u128iiTNXAmpyn7tk/OeGBAyx1ljzB0QO77
lPW5Mt31PJcJD3djOjN4xSEY9Q6GDD9htf5C91GrBo4Y1XjHuTXSxpSfYjGmfXrm
47aWUMHZUttSGcnADMIjM7ZmA6TLHdppagE0TUWhL+0Wqw8/pl7baTq4HV1xKhfh
lNcQH2eBZcfqz9F5vihuAtfTpLfen7r7GhzXvcddmFkZgjcK7qCBegF2N5tG71EU
/RnpJFyg9Fmuntk/WZ8K/pUQLnPvURjjotsuTz3tMkcVkdRI0Nl0W84FcTtfpwiZ
9Lv1r7/Jcl0+9ZL3B4d900dtpAY5/pH0Z65XTVQLmaoexQGI5fmWA8JMehmKfU9M
HCMclDtDMIDrXAgmslVxOD2ydMDCcf3xcr7gXDqM96qpuGxIuV99kt5PKRk71X0L
cgPcGoM8n4hoMGENbDXCkaG8E/dE6Kkj4dDr8v+T1ejm2NZB4gUDovTIqX9xPBOV
7MQii0hFNizTj8raccKlVa9M7IWHDHQX8uSnGAQoB2MHkJDJMzeVSMWogKwtLo6Y
B7jvQzsXY26NJUQa0EVZMzchPP2fIBXjbKPOy98H75P/B7bj+t5F48mFJZcdxF7h
3ln6bKZpZS4g7kNLX5GbSRq9x+dkpZakay+BnDvY3MWk2JFdX1bhjxM5RoW9aLDW
Cb4l2YbPxPyNdorpInDDC80lARelHG0Db6DAyiWY3UbgHXHUdi0SqmZ41VyKlJ6l
E6eR93lCGFiyTvn8F/Li2T3mRj/gWw7mqeDLncH2ay1ofLX24zx48Lk8A0aHGVjk
99o9DIUjfWUIoV7H7o7Q0sTpSCxH4iOjjq5fNYI8rzvvCu+a5dbDG0aFYhEgn6eE
oPPzd1f8/FiL4MIdncOO2nc9R2PpUBC24aWRPOWY1BHNM9wu/0orbam3+jQ7QkHy
Yz1jzVgqgFo3NmfuKhKFS0c2PvR1eVJkvqIltB+dDuAVleWysJ6hKjuQRwT+mhK5
TeHVmhwcEDVSdG4XRH/1yFFb4KAyQcqMk3sHHYO1mWMPL5/HBjnOtfJIYt74F9Jc
iyt3IMh1RtaG1ZXhr3YKZok/0XgJJVRZ9bBEsAdY92/1/bqFFc6oQ2rkKIm08cMw
zJZwK5qHcQe7kOC70CBkF6pA3iAHBZX2cGVbe+BhNzA9/MsHiwyZ6MXlICo+p+2k
TtHE5mZhHEcX3TTlDzw5+RUGZ5w9m7kHPS/wpG93uz6+OcsdWAVwAjC/bO++TFpu
sGeyS0DYkyInRgUNdc6U1LL/IYAoUXyaxJiPIsNMPf+4mIawftqjfG7hFykv1mIi
DwFXHB/Iy/QZoHJ7hx30TQyoZ/n7zzGGET7IRsqY2UxnGsixN/0PmNCvpIFhF7TI
ErRxuQXduO6rmHtoUHnBfU81aXc/Y0Gzyh2DqM2uhSTeODb1aav6/xtAAUPdBsCy
tzemnXs6vw5zmBF7dE5Rvhxad5LPPnVJlwP01KhDcwP1TLBvLs13G09DaRrALFUn
RdhtbjlTU/NRrCQHelHh+WNe6Gc4H9Z0WaQ4Yjnka2JN+Rmq1xi7OAfeyPhUIsti
WBWFvTZeW+xRG+QRwl6KBK9qRcmorN0Qr1MQv0rzJeEQyIEWOcyA3Tm9dK3kE67w
bT0jFcO5hnp4AqHL7wAGQEay0OdycRG75ZmFOs+XrXAx/i4fC2OMg27FMK4lUczV
67g/aJutoJcRdGrWxqncxawEBqDlM7zZsIx7N83tT5rl+uKYGVvKlb9bKioHv4CS
Iv0JnYdTKnRCmDVVkJwNecPNT+VN4Q8NqunDaW3y4WOp+H4qqiZ2qS50Mf85dbww
jUkeuIBuDlgYUqmR4DhUARtzrCdnh0gR3klG69igyRRF+yRJP3dt5JxETamepbgg
EBOPZiEbg0ridixtwwQxOW12A1rCqEF8kIjuljWexGbSqIBJZ+9Tk53jM1ke9cAp
lret/0A4QC74Y711YDjQZZTIDZV6gnXQhlrqHlso1KBlyOmXdTqlZJsJIFWPtcQ8
mbc13GfFrVgxDYxxyHrQLqbxeeeFDb7J3t+0bS1L9Md5jIxOpBCAACoiFnuBhoAw
SxHFQ+E3Fi62B1Fzv5MGCRvjJ3q35Aw75Y7C0+xgeo0/hT6OsSwFGjNMgUTu0+C9
UZYN/HV/IP26hxj2WbOfgjtb7B4ux9UibuiraV7z+0IR5+Qhu03rfbet18qQLdgo
ramTyyrt4ALXsGPo1lAVx50guMgpwEBMGxcrJiJRfkz+vSFTEj+O+1c+5vszgxqy
3gzy7kOfu/M8Ra70kTWXFekniSeUs4iwUX0wgAGh/N2P6BQSQR+sVWoE2nbb/IGF
0r8TkLzQwCyM8sq/weuMC7MsSo8r7DCqs8X3kFuM2U4mWjaVV1bVwRSFAZc3lWHk
GDs4Hd6kYs5VRX8GwT9XJF7LmD4jczccus0c72QNYib7Qyn67PUJ/KnTMXd3XkCX
iDBxuvqNBKX2xM2d/lfjhO4PZIdWHgnbU6gcnGi0hcXvtWXXA9EQsSo/YIxc3QE3
vEpUQzCpCfLQr45T271gj0G7Y44o/DFetOMTQN2kgSDN6mJxdQUhkEh9EH8YfRg2
JWTXCB9AgbXDJRgtCyA/IaHiGypFlCo71hRpJSA/JCYLf7ppOlo/BxnrvxX9nAzF
OkbUVDoHQ96ifvdH/wDtvghzbXpNRlHXJaVKNsFFw4rt4q6y1qz6hMKD+ty13BZP
s6jmD+FYb0wEhqobii/4CDf5UxKQcaExyZ4UIlV1r2OKCrG7kIMkPw3f0ZtxDbyy
pKgkwiv7PvtjPIXXgy1WZNRJr+BrSql9WFg/wj5X/8zscBmeAMaa1FGMq51MKQyu
uhUy54AsaOFCrhm5L29EJpixmaZLWtkkTPaPY7lYy4iiLgv1n7qupRl3pGPv/D1Z
jRrRXk7Axlqhixd3zzcinkKn/khNpmSZBcK/A9O3RPSRRkFSa4D4cRgfrMRmAtvz
QK1OXOFgnkfiDYn75d9DqN35Yvg4yCEfPYfsA9O6NvBJpQKBCHwx9JX2qI9bcW+j
hg0pd9vDDAbqlMkRdoJ6y16ZLHVm/BGoTijyccPpqKn1sZsyzeUTc1+KjYsoIMmH
CtRfNmC85SmdgoBtgUHJS3j8o3AY3EdKK8NbghxzuSFt0r5N74uZw39vjWcQB7Uq
ddQD6ZCAh+sTnzfsOxxndOYCxiElHgw1uKY60WRYk3Xjc0LYXE+SjfrAr/LXVnJO
WBSj//kQR3ivmekm50esauj5vVMTDAnC53mCGGQhbFrm6L8Q/R5hNgWEu8Z7BrWy
vBRrIRYdjGhX/Sol2WNoD9cDDRByso5GA+KIciiHnXM8163GbcVgSO2f9AHyAVJE
+mQvZetdMFQ+lcUocXKXIdW18gzKk3NvXojwiZk6xdRZw9K8TGn4mxp/7Min47Am
dqwqt2PHNEvrMZaEDLZw2pbHzVC63Antot/fnW6337SKZmD+ezmRpKJHUUDOjR56
60u7JvJINDUEvkOAwu/etVPHydfekhXMlOq8ddTksD5yB08yqUxZkrSM/nn1zv/F
eBXD8iHKrBbynV7x72UiDDoS6aJo4NjcILcuf9XZX+egITlX3WiFccv0NwPdoFB5
sRPNL+Lk/X2HGMSw+EFwiTNb0n7hZkP7pYldgLD6b8j1IceigGfHeakQ1lKSnnHm
s+YXyH0sKKWTpETzzjxtLaxamLow6P543Clph6ICg/f4IFxPcueeO8Vuk8KOKRNi
FTzDYZ5D2KPzkjWAKXH6jkUZoFKDyTs2pdH+lHXVQErJgjBle6rJKBtRQ8E0lsFl
a/Fv6NGlqbh3U2TopRery0GmmAgh113FSayciJQf7H3IoFn2XCCRqd0cJwh3gsla
pmqF7bBuf/GaQ/v+l6rek5TQHvDJV3dr+HDcO3+zrF5sSLKn19mKRsfFj1/ZUvCY
mdE27srYOdkvUT86d6NzGw1gYOQDlXJaxeZCcDFFRQmlGWliTRk7OJ6IIEs3EqIz
qZUBZT3IPiGfa0AkiPr+TGarqiNoMzfx6+Lsup+LV09phRyHyTsyWuWQtbjTJuo8
IWcQefvY/wkGRe7ren6rNZ6cve08F4WKMlq35cd4wgj0A6OCKvFuXe/a5JDw2YnA
htbDova7c7vLi/YkFvIQDGYq0+Mj7g9M4eC0ZNUmgl8voacWZ41I31N7DEE0C0k0
rVPDbDNesIJZJu3RjjCJvUiQ+QMrHS/dJ9bejA+TnkFmYvlvG9qhkJ9J6uiBWiNa
FIijiQdagWt9y01HxG/GF+j4dAm3kI8Idp1lpYVNpALvM/N5QEW2UMTB1rbKW2Eg
q2/779GHG2SBHd5VRRo2y19/NQnRJbqtgtbgGqc3Mcbazj5LsnQb0ZzfKTa/x7TA
GmK7vJS655XwiD/IAatfIs/WzFk2k2XIvegarKpleNJ2vMMF8tJS04gpSv7CUJg8
HG4o8R/l0xqmBHhvP11YLsgORkzY5I45F/7r3KcjNLOBG+cIfmDUHt3Z0KG6lQ+b
++3RhtKTKlz1K7UNZnjwha6lmhmJJd+HEp4KuiQrBBK9xwTWf+7dewwP4l4nYNf6
aWkAZWspskybMMqzPEtZL2pK+OPxIzfGOroAOtMO2XB4keFY9PpSeMstGRxXbG3o
SoTUfTtL4JEODHUm7Ka1ex82uKcD1wKFP9pS0OmErZlAgN8TXCASCQaEwHRH1IUB
NhxECWEkNEQAD/HX4LKhqaZVlPXK11PlUxom8H75xPD9KhSIFBO02m5GCRi9iKWZ
9Lqq50B2SIbX3wF1rYTC+4P2snQ7HR6Mpo/B3JxA9ngxi7rBWAPX1bHrPaXBsTln
zUtfouvgyUpiJxHak/AWu+F0aG6FbZQuI21iKZkaetZDrGAgdT3kvT7K34MzjOxU
A+jsKgVjrxc8nA9nY+nBehd1d7RjnjhIbmVR77ZVA47jJc5C+QVG1pu531o0sdLv
b40WR308rFkXynF11NuBTqFS88cUmgWt7JMYZIq1QeHph3/WaHIoE1ZrKQXglTJi
WPG6tZauqq1RQp/SvtHCoeKFibZO/07MYXpWAYOgKigHv1vPFWaqy4zYLa6zyCu4
gr0ngV4oV+WIT1jTNZNjXOSiCsjvkMBeRWkDOttTTrNxOZmjmk5Rf/BIyLIVNq4U
GN8YaEdz8uQtoaaQKK+CQQyjleYZ6DrE7/wJQX3AMJ2Lia6O+clwhiIWj78eIzOH
I8CiPnoFZbfKrsFslePl2gIUrpa+Orr/H248xv3ztcX4CFO4kyQ+xXeHvnFDWIgp
rovBSWzQt2wEnfNZe1u7J/mB9r9I15ZVI2uJ021JRSKK29nBBCnKHyJqsLIF/0YI
cYTVzBSxwVlkpgVutWJWyEkkhSIiJqf0ZRAMnOyW5duYOuhw7NLkTnKgiSLfjDmJ
g9OfxetvjlQS9wDA392xWOFOOn0rUETQ1+8A47uUPeCYPzpJYim4BDR09cYIN6Me
X7c/NlkR1arwyQnDpVfUNsuSYNeyDf5f3mcX0O060Bz3SQB0hxfFegkvJ//FuhSK
iUq1R3j2oj2mw6Wb29yRjDuHLoke9cKHbXF2LPfsYine1PVBNsQ+E59n+LaZk/PL
quRDs/df/eO+3dvEjLekcTB+UJdlIgwb47r1B6cbfC24Z86GbqsySwtwomu4pCvP
9Cjf978fJwSZrLZnXZt8au2LcMV+O14jSz/zQiFEPWwRt/GYdEXlvMMjDuQXNSsN
0mqiPs6Q9r1v4hTkpZZLM0oDO0pRCbIvzA9wEjgiEeKCsIHeL+V5lFJxMdpqHd52
lXto/1XuzEfJTm9KBwhaom/yswdhBA3znvakC4JR6HjSwpnaqoK2wdcoEwUPaxf3
qjxZUODcJWUe8rLtnTZgBkVApmHb8YUVxatTvDygKPThflA9KpABEaZm6DSkbpUa
Bw50hoQJYT3gfXqCQIio5sr7SpUcqk1jiISLdSLUjxlXOKCIMvWhxgSbHO/jc/y7
BBHSLdDByU4gxC1JqpJI/Hifp56AWQCfKogkcQJ7YR6/tTl6TJz+pMFSWW0iBH0F
X1gY6JetoLVSwr1g21j3D4rJHUWVbF6ofX8p4zEfKpW28p4eE+a/ZLIhtKyGe1pq
PLO1/zsxvcJQKssSH+eWTd/S211bu8x9xpAjx+/uQtM74oSwpPxS8VR01hKE20Cz
pYAJ3MlktfGP8B7NFJCpiXpPxN5HMZbJAbmolGSdQt/8xWA01ykf+49job7ifviG
gEDW+GHEb2CQ22PGzsmvgEYnbWpEnPAW3ocw/nKJ3dK1BtwFv0TaYvj2JQsOzjkr
JfDyoRqvSOtXbspgpeJOP8F1pgqfZQhTiDaDl7wm5OYENhC6Xul30poPPankdYau
LU0ICw9abi9vBPhjs08bzgL7+X+g8/nGQ+WXiD7vrfsh9AJKRcmQTUNUsFqWfMp7
NIyy2FZf4wBgVzNUO3DQkBE+znDanXapHM5zvTKNVLZmytNbAmeUCadu1wLRKFdU
qBnsY8N+OboiIiXuCSE7D8VHatPOIKQvVptlWFBCaEdU45BUUCK66FQA/QlUVgow
2xJVKedmB9vSttK03nkN30Fw5QLe/xNGTg60+cnaXxXNEzjFoU/HBPhFi/RgaAix
P62mOCdm9sih+W/FFuqmYWWb3sA+ZnqeOvkd5nrj3KbqibGIHRct5Z2Vg2PTblSi
YySHw4McHPCsgnNTSUmZz8u90M/4ECsmAGWr5BgDoquS3nK2ErvSdxc8LpA5WW4p
W6WereyQp/yHdYrLqjuH0REce+7DlD48DpxqpfOKEGwK8DAlFuYXfFy/PKOCsRGt
CcNZ6ZgQd4UDRhvroxWV82xp7vMCFfWnWbd3JhlrbPBhlrOD0pJ3cvabuUxkEKOc
yBJ51XnGRqr0l9ykJbmXGfybnzsi8JtGCfo+BBVYYMtlkQUSG75FH5erKDtTwwgs
qgB7Mde3U+9E9KF/unRLzEuQr6rPQvQhB2UWUZKD+7QWjeL5jLIT6U2MpjmsrYL4
PflAvsLed1/cogGj57/4sUMauUhkVKMQfNW5KZReKf9BxUVIHiy5LX7d620EcjRw
GzrtBYugtibRi2WEmaFZBiuLG0ZeDw/cECajDaOSYWywARZM3NgP5Nyc9/hyjAT6
I4r3wH/QAJGc8MJovRGYRtmn/BWiSckYICoC4IT6v9BdKb0CZ9ucCSR96fiGpCQ/
6jHKHLyJPVs2yfjMm4wdS8qJTAdj4Gddg907JmExi8xmtqiJ0M9HVrX3u3Z7kdwC
uCKSbDDbDq3zlPLyCArWp2ZqbPjmNis41ttVADPe9zH6mWyuxja1IHoxGKUn0bNd
8KWETIIm0BcDAAHel9IXRq5TZgAE8ahF+e2PLEwdYsazc4s+gnxhXqbZ52yrdoaO
hNk2uKoUIPIpcaylvngmPGTUf7tgAHf5eL2VUVJ3HAj7Iw99FjH9Dtw1n04E5+0F
/O+ZR+Z2EVr8x0iQrPYmP9xfHXc94QadSMa/vj/hbDjXVrvQDWGNIVs5LhcWJNH/
E1nhi5ZVFxD89lh40atypLT+DKbn+Ns1CvHKIEl3pOBN16gl0C79WLakTf3PvpKe
3CnRCXyQ/0vFZp5TnANr82OsiNVLgnJYpspKx7m+29rsrG/mIAlyQsSgAZo9H6Mo
k+kCpyabPkxKXpyFHbXRpg3iDgczfPkRKo0gl7YU/QERmKk57DHEqeg2mTrdDioY
56Kn4ArosUnSCAzJy+tVR8eLX+sPYKiHk5tbTfC+uMb8Uv1jIb+2tNpG9SMmvrGw
rhi8H1L4CbDwqm8/pOSBXmoApbg0ie4CxuecAajNMg5ILL2PAQVClPAHJl8wJPbj
Y08Mdh2pJ6Y0yDXReHuhzQKaMdguE9KxF0iDe/1qKX0j04MFaFWSovD4bgxL2Wri
DOzt84sMgx8QrF+HPsm7jb03qllgLHX5pJdJr3Sdfn7llDoGCS+18owJH0xqyC72
Rz4Xo3g1Zrv9PkG2p1fh9z0I5kQWqF0K+srQGQaObfJZ1P+bZvhChh2NOTU9hm0E
asNgLREZF1fSilQdPZzP0uz4NOXyos/ng6YPH3A23ykv2miLQLRLvhakZm+Nvmz6
hHSiJrAOET4HXzaz50NrzoWfGVajpi4K3mPaBvcBdR5QWGQJNsKtMgdalDJLBY4z
/EMk2ouqwUhwJwfbXT3gKYeMHSHrXQnGnxPJVkRN1kofgR9WCsgoJ6v2BbZqFukb
YSausMbl/+nmiGwLd1It5Z5mrWzIs02cKtVITopclTAmRdAXaPvAcS7WS1SCOyuU
V0oCJNQYzhKxhJL59pUE6eaja3OvfQFdCJ4OjWIzrw8TdKSw1UTndfZTTrC3pjSW
xiY/LUKRWFEp14k9YW1ZwwCzB+be7jn8TV4pB0c9nj4MHzjVUNV0/ojOsQa+vK9m
0X+dBkAkixhTsNH45BOp4Dfwz2/BNQRQ8T8AnWEQ64m3qRwogrbnhrCb7LHNLpW/
gi+KgKMltDDeMBnJXuxxaPYesY8anOWAnnyiog1QJOqkxDutsR57DVtpZYro2NSO
tx4gkSKv3Cjwuc1rSpJJlut3wOVAMsc0AO/DUkYT72Z8SOgC+KnvyB9bWSTYTQYW
WX74lYpXGD8XbsFxnUMZGniJjMM+8SgbYo83gLv4IMGXI2d8i6UlgXyjesiT80LT
d7qzQQVXIxgjvM4r7hcllMRowYknQopRtElHus2D0n9Re2iDeZeu9i1AFXiGIOWy
oyRfoJO0Ez+byAzGoyeeL5ii1zDUY713xjC1mqcT8zX+mFGMiiOFWjiBdmeKs8PU
8eF8N8j6KW0elKys46P2Pyk93krLw01oSQyNHSZaUxaIjB+abtZ7EzA4Pt5WPvXY
ymeU/hTiXB4MWuDgfKMeCXCrQo1OzsBv535s1Tf/4lbFSG0jmQFWfY3cOyXliLq4
AOI0mYGBCKLcp95LVcQSJdGgKXegC5HBbMjWClTUQK9cpSTYDTFW9/xf8xLo1ugj
Jb4yZC6v8EM7+rGzFf1WRrn6FNuU7Sjte29cYhUrJZSKYtvK+Zw1rI5KjbXpjBm8
yats9QXmaYvI7mC4ikrH61Q//l62I30nxR4WBVSs5ofBhDlpTQNsxyxMc5srvffw
QQ+FgegsZV2hWGEXSAFklajPZzWvMqD+kLBLb4hH1nfU0N+L85AzX3z1E5YC9XiB
amtg3w6mh01TbOkkrL9OzgqnKnCLl4ulNc3tpzNt7JTm+t7/9xmf04+5bhiasVQV
M4YOTUvOI2NkH2VfIR7XM2vL+D+wr2GRqfH7l0sbznf72pBTG98MOMH1QJY93WQT
2K0RrQKu9ihfDR7moXvwuMdlUaEqbxIg2538J6D3HGIONsu4DUPF8uYCdjb5hgha
pS6P4A0EmUL087GIlusFNn01agGrjy5tPjH9vn3fshzvzjOXOE+KT1iUd1XKwMAn
Vf/JxY8/xA4453sHtdyroAi1loy+0L8f7cswWXcVxdIeJ+mdDFORcuzzeOOlsMva
u/8vlJ7Q6TAvy9Qrm+9h4pT2irrtTvhNXRQbiWDSs2h2iLCGW8PtKeXulU7OGZ2C
zWMql6PeZTn5mjo3qCrevDo0qY+xvQft+S/soPUHbUVcg2d2PpDSwzoWpfHLNlBT
vIJ7lPsHLdRK4p92O1OuUIk0ckC2S1PEHNDd7jk8mS0ymNbg7FSC+0YOvtUbz1U5
WCiRyOheQVPTP+R+qnxKlx8EIZ/8wlruybAY2JzEb9rzJ6Ibb+QGrWE0ElGU3UVp
5GUC2aZavLI8wkKF6+GMNpfLyCfTSvzUin7CfokY3Dwp5lPPW4h5ZU6IRQXxEeQX
RrkWMjM6REZ+pq+md9zWfnFx5pjt4E46D3NE3X5hQeQd+BxkjeK9iWl5lGPqSLWl
NaPIn5oLO7w0iETXwgnPxZJf06VoPIWTrcXph0Z0NcvIOYY7+ZqfgiaXIayIdEXu
DnfCyzvHWMC0ACxt1TzCHjwMiIsaVJOKBWSq2vpvO7y2iTFZfdM4ZoF9+XXQJv7z
lgZg+QmX+xrL42N5aRqCNO5N/9mhW5P3jzsssjUDMnUP09CcfOsMBAevWLDLhuaM
vj34n2fRC2fElj8X7yqWZXe0i3j4XM0fplB4bn78pNtWtprDNUuoa7+P/Zu9ltYK
jwCOwwTfqmJfeIjuEN1thQCbgmsOhhMnh4wZAPU1AsS4oSNr1MQRPazjElRBs5Ha
O7js8mm64fMThqJYniofHIWJAzZRE1lUSF6lfRaRc3PpHyTJrFW0mFKiPq6m/av+
80LjbWGB7OlJxrVZRDcm/dD2i+IxurcUOH79y4KFsG0Qih7QO0hLh5/f4rbXYaAd
isSremQkoxF6GwMOWlmK9F0Pw0J6QlW6K5opQaz1pwltrunYVKOSB15SoOilRRN4
wyU+t5Hk8gbS51emz3UEohrfMvxwEsvLrCYYEAtGqAdVMFVng41tZHrxFqj+HlDm
urBrQK19wNC880IABAHhgZsf4bRquqo/YK43i82p9LHv8u9bjBdl4aeKTlU0ifN/
uXhiOLjrlWwLCj/ZlPIfwTVTbgRGCDGWAZh7TPN83sv3fZTV667ELQBo7ngs1D4l
omle56H1kAx2ib6OFZoRx8ww5hyX5E8Ok/zAJksi59UZwZGGUMK3D0PtcwOTthCs
5NxtsJbIK5qmA52WUnPoMIs6LNYt21ctiOQDBbcJmnS+8ZjnO3oBU+ICAAVg/B5r
vUyr7DxPosWL6NUNXsEQLgSo+Rw493zHsrK+hSxeIbwpaC20t7N23C3WrroYTmRM
IBdhzDr5RhorqVht//mtl5N+9y8Kje/lqpZWmzvOIfmhCLfihPy4cFQLKp+1KgwT
NpHDD2Ulxn1M9Aa4pjVaxgtsle2a0R/0I3Td/HlFlxM+/sPwzhQ2yGy4fW3tdn45
gn/KndH2r8t20w/zApBMLgwZnB/3y3FFFBA4MtYhGQ1BFZt9Vn0/OHI4sT9uPexc
H2qH02I96JK5b0L2zugtGX6Dlzq/DgmnC/+LiIaI9JIOBqMWcofkt5dCYGqdtCw6
jZqtRrDBtOSlO6DrN/DJrLKVHN6oOzdf7dRv4e/9R8SGf/Oa51vmRRfmZPzGazfG
TLQIUHKnbWOaNN+7gfhN19HgXJ4zrBm5K9H9pMOiSCf3ijkRXa+cHYL/QAPhmizO
X4HJrN3xEc/fCv+OLKgNcumE7V6Eu6Bw0wEEBAMjJ7Dk5vy3JeSouZKN4f/3XXmj
JnOeRprAM/Nfyo9A4A83RwzinhWFouKc89et3VokWyAClF9xrPiBV0OzHRiKxQH0
y1W8J95z1r13rXCOucKitDn1l7huN7FJXVx1b+cxzkEBzWgh/jIjfI7tl7EAt0SU
s0SlmJM1/nnAjwnO278GmdLtxo6NhrmGPowULpK10Vq6y2Doic+WXk3yDD0APJZr
AIRHHhqhinjtrUXBg69WLANWM92VdiVjZC1seowCAgaP36u6XDGPlKGGzQwWyOrd
E2BKCbJiY2jBKJf+uZIUVdqrtamAH6UWl6FWmWSBfyAiplq4Lxju5EUiR5JemGt3
ty0MUr/PaRMv+ZjCQZZO0h42GOZf/MkY65MGsfoOXIf4m4LoltUYwm8I1Ov61uLf
QrAdaZMyvipsf8N8erzlHWyNzPRggDkFzjMFJVwky2dbLnAyME1Zfq/UIAogpRdW
iv+ByH6+KbAzkqwA5OWqxt4wDsQgqw5BnSAkb3kqrWVqfJuHk3VkWZAEALVL4ooq
JqZmDSfkaWIVDjIystX7NAjBrgXFh0RSvHQxWdrHHqdSo06pcHHBjnqQM+ICGYW4
baAuj/P4M0ovFL75MJhmF8rI30KNXE7vlsRvf6qhT+s8vSTeyRSKvYSFYSoT9H2c
/rqBKLw602mY7jyNZNGB8PYd0lYkBCOAtZJI2M/EqJm3OwopO5RGrpbaFtxQvA8O
OIcU5Q/puG/fQmka4EwlztjuVZQIV++Vf3Xf1mM+KUk8XSaVYlGtZc+xVf122/y/
aQJEDFERWbw+FjNRgcN6pPl6NCejltggLLHoXZmJldPOh2P9fnXGOonEfN2TjeyQ
Jul+ziQZZvgCUhfinjCo86ShRCPVeQSfQ068kSyZ8ZIZlo1+tqvPLrB18vqN57Yq
fNxA+mBWXkzjzzLeg8FmdQ+HZv2xIyAaOn0+jlNxGYSyhVtNe6lCwTcS/HZPgokW
R8bSH3vfr+SlP7cMjY+sgr0d3fiYiZMJFlxWRl5NOfQquaEXO87pOB2F9IEpC2tB
TbfuY/lQQw22DMOUgoreveNBcLRfz1tAWoguczTA1bwYShNV1akKQQhJg84rxZZ7
DTfqfJ1HRinKDBCAdE5JFLdae4DZM63c6m2eJ+bDfW0AgPAe4gA1kEZQpRpLzaBf
DaKZtxoem4K6GtSM0oCwaskFbe6QfX7AeUd8Cl0LdtRbgGgbce9Rw/Gx4B3xF0AE
+oiFLq4v+JYEN6aLaMFvFtmcnf2y70bJnCpfmGC7FVOlG3kmGgGDxF21zXd+SHGv
2Zf5jJ41dpxHGtpuydVvTLmkTOCsCqIIIDqJ5iN07p0pj9xIxxrkqqQs7T0So4/R
cQQZLvQfspmvPk9Z9zLGi0lNK4q4eACJ+ut4Q7ESvfwrlfoZo5V5YczlbLVoRGBJ
PWDFXdJ3ZoZOlxy/sJWPDBMBXrQcEGBvuF9EFhOwYxSscMbCwcQGQ2Kw1O1OCdIL
rnMlOBSBEiffoRC7jIvL3i9LZfe6GYlk4PosfiIjnt3sKat2egbV3k32DDkSKvq3
WeOXxYrN1dtk090qwEI2HEsWcyMfh6T61C3OTeASwnwsaYbFOAdkZkjHe7S6KYYo
Ra7dEVzF+qmSNEu5zUz/mH//YlChl4A4WTkpacmIvfFvMF855PEQKFvuEtGUr+Fa
6wavZVtDhv3Kva0il792sZj77HO1uH5VnG1I3w8BACeJJweeg02sdb0uP4JF7fQV
p/o1h6I0UauNS1I/4avQYSihy1yqMkspiU/ltj2A3005Iwkw5vApkRAhwuPmn5yp
6TSpsZ0X4VztUOcT22TGDkncdfNpRG7gmwlsxFR/5KTZAlN7rDga/sHoGtUcCsUh
UvH/Cc7ZrgrEfC9eQhq8g+P5YeOJvPEV1XuSfJm8wntcrIsOFdy21b8tssGhL7T3
OaZ3GAF2dUuan8PgWs+6y38Ld02xMNMpL6SJkK6OrMh11fqrcVNAkZbg9GvdrdwU
7AuV+o+C/kYdm4hKtWYsieoJQQiy9NiQ182cZ+U14+EPC8eZuRwpzeczdk2lGN+M
KZfvzECO6JsitLMRNoD2CX/w2MiDg2kce7jD5+cbSvVCkwLI4kbrbqoRE0kcxHVF
RmnlfaUsJXA1J/PzgV7tzsAdDOIeQH5wpl+NaLIpg8Rsq3rTzdymOhbypb9DU3kW
3mgdxggZ67sDIe+Cg26LhZvcj4Gm/6DaZQaEzopDCQVsSclZX3foNU67vduyDowC
azT3i/vF1H+Z/XnRB6BvHJrUH3iIX12G4ipkQE4QrYgZPm4wZiCSWerxoA78DRE9
cqOm+HsMZdatk4Gl1TVrYJKW2GBSbiPUQlu2wa4sONY4CcA92bbLUQPWOvl24sYR
OTblfelYAIizOCih7FnFonztf/UgItvg2G2dJynU+xLQSWkR2zGTiYy6PYp71ct3
TaZXHkh5Cj2+YTHgkibrbTMOjuNw7yucJ4srquFgzqu2ASfOQ0v+MddRkttpJWWn
aW9F1x5W5EkWqiw8G3aXjIx85+fOim1nUHEw4oRDGra1LSnBiooy4Yxc+2t8A9FI
4/bFln7cNHI/dExzkAoPZb5NJkuiQ62wUIVupugbT7ZsCZg1BeH4H24SUs1d0PmJ
SsOx6MOhYlYw1naczIWUuOWaGd7vFLcmanLF/2v4TE8NAxkr6ZeltDezZC+mtc3S
is/FPKF4jhxw42kA1glDVIszfz+1gyrETJaKvamsVRefMPAC+/SbpveWAf8J0Se+
YhOnnWeXlbG8ic7Asta1UfHrPbwJwRpJYFHQ/n9WezFScl2eeBGN1mjzswoKIv9+
Nn17rJ8mZZC1ItERHgdHD9bfYGJRrc+z7ZNIw7A2RfVUNZ8sL+dJ6J3gb7O7Wu3a
JP/DdbB3xTWIvZf3XAwc0FdmMpmp+DbdV4Aw4GIAoFhiaCmKYAlJ2zCo7sZZ2MmI
2aSB9jjL2KAbZF1zw1inh1/bAYCyGjeiX9rZXmCT8M1EnEm+dgahxPdNqZEfWBcq
WxF5OfQOg9xdBi10T8lIMgRAWzbaaST/7naErPFukNolm8mkOaLpuzsLN5FbdLp3
df1q1VxGt/xZ08L2RksdJhVs0kMa5nE/zpyajB3Tn1WNESBTkEnXRo2D8yNBVtjx
U+1h/p8w//X9g5zsiG3ROH4n6pVosvWrnQcafnqzaxEpSbuD3ueY2ifi3aYK1vzN
TFrfEHUAP0sZVwfuIiv1G5Ab3P6Ij8vHuUyYVrZ44XKfpRXpUpRsplSHj6riHZc6
2/JGWL+aBV+ewgWqrHHS6zx2paPb2Sq/ULcU4v+NgXLpcL4V9+Agq/myUzy7cv+P
8FMD60XgEQ9XZuCAXfZaah9MNVP15icGAzwjhnLA7/nBO+JsamOyvuz7s1bVoX9W
pPOm5hRwzhwky8mrJ5NQi9hWjer+Cllcxrk7gAfZ9AVlP9DLV1yxG/fsLgvlkkLV
ykxxBlWeJRvH1loPcWT9HNbSeKXdWE9f4UAc5jwUzfGiljseZKNElRwaQOVxWcOE
02WUlPu/PL/5trVHxCT7MMaNtHEMahGO8AOxlROte61envTJsZIhB58Pd5JqxcMn
2bzF5Jbs8SiIOZ4B58gNDu+NSItZ07l6740vGp+we1Jf9Z+NGvRP5aEqZxgE61Y/
1X5lBpiPKnt/P4+1fqpwARPmM0YZu5fL0Ez9yiSDoHcb+KSnDPDNCkVz6JYlqvFT
n3Hcwkqc42jb0D1kha7D8Sjd+20CFjaDALI4p8I3KhfkIoV5csL9piuZ1WwsvKq2
jJfHgzRSLE0aiyuC9zjDm8zbW7nJX28XAfjcjodEmMJqMeOLMwg5m57r6kYU/zcc
/C9C2ivYb0zv2aksvfYRK4wu95oJcnzl5+z2G/tjiCxteykbn7WQDph7jOD6nMCK
tcFrIBWPzYWc/xYOY8FPadIVHLTrv2InB+pSXsnBbibs1xPigO/N6kQ0UZg8Da/w
iBP55sp8a7pVoMo/omNqjZBEyeqICD0v/qe8dlIi27Tn7ZYRthOub6F6n1rk7e4w
9k2WAMa7CtWtaSxo679HAbrs40qWQjVvr36H4HgJx897TcahxQzp5/55KuSTbdtx
8LPqa5t2vB6LDMx1XZqm9UoLaOTppaV9TAs0YZarhh6qJGuLjJL2aoqFxpmoOkdA
DfscbnCj/WmmwV9BRuU5zGww2hWxJPqzvusS6RDeXfTozN2PDZsUFN28HEgt0zu4
mVHDzhglahVf7PyXTxveziivUUqvtq/09zj77vq5+s53yKLRMfIXbEuYcFGwRbay
bdksljdzGrm3EIEGrYQcxPV4Zx4WXDw5DQtptoH7eVg2FPkBJR2CQA4t0ywgvAsY
FjiC8IJRcEe8pOgwtBgVUIXccCpLyGktnMus1Jz4h5chk2/64sw2GBIOYQZH2DPe
yltQ1iCfsBfxypZdmckEevUUiBWQkKa+dm/ShhKM99rhUvZ2s4/2B8A1bgAktHwl
DtG2cH8TGIR5MQa9rSiqjPgts3Cek6GiGdF16uODzZHMnhWkVMLBqFEZS02i3XGP
yXNBeyRWnk4RSQasIu4chIjLADxhVTQIU1BWy6HDNT9Li1cT1RqqUbE0vqublO0E
vG0qZz2mqMqJHnGx0YwLVikvB6+05+BgAlIYVrRFxnfaUtq3NAsGlPBen0W13UXN
rgEMkYfAuSB2BLu2dfMPbQlV0qT7Ziq2iaGTL6aVJ55J61POBI9qIppJKqAoL/7W
TtgOTa1YoidyG7+ggi5lavlF8ZfNQPbUOzTqJ3sad9aFv2+KajROW5ZyKwDB0rjz
+jPhkCjJdQuzVooX6N0Kgz+zY8QriXbi0huAtJhzAP9Ykl4N3rSlM9iWZB4f/dwJ
jF5RXcKd+RDMLXCPg08En/eJvdkfl4E+vUrYU+ONdGNP5cy/PqOD7LjEhQWxIFup
tUEBWwt3FtD1hnddC/aoIHdrs6NPA8cmspHyP9QDfl3HYNHD2CAKIPXXOs+9FIze
Z5QOxbHzL5gGsbrOD+W5m4OH/XS6k5ofu6p3FgsMk5OwrblgpabKfae8zPmSlBvu
jXSrMRpO8sa2htR2d/z4fJA19ngb24D+BXGITvqOewyxTEoA6YwBK/41LvAtvusR
xCh64z39mbyvKWgqM8hGwMH+SZhZAJdmx+skI47UR6ZEk1AZErn5AYUgB/3Hojqc
xAwae23iJwONRAuEExzLrRIhyRKvTfISpcPsP0lu83r+at+cqOM6ZhWwzHRhrxFe
ONM1Gg7I1akpSDZEjn8evUtCTDqCnMYy98tsO2AHdRn4pjjp0O6TS49iGP6JoP/J
+rzMvh87CmJJkIbpUmN8fKKlPYS1g1iqaeZObTmROsV9V+x+CmpZETtgavgr0t2m
1QbGOZQ/o6PO3Dr6tngogo7cP44+kw97RbfXRBevdmNHevovuEk5rWBuDiGsrvxp
Jvuam5mcgP+C/oVosYbYyiJc/+k7Ce/t7pKKVjdWtMR6Z/ego02dtxmIkkcUuxs4
qoZxQOCpnm74WbAB9ONTqW74nw/u3MyqqiXRM99Zpokg//LYA89wgQHSoI+EDnln
QAlshmU/drP82axjQ57c7+VA3fhsIdMaNnrec3GMeUnH3cdk2Xvzqc8FmAxFZ3fQ
2WLOvN41/X4lIcaL92XdPsuT+e4TTljtoUl8zHHuhnmSvLxopIEWMPerrLgVM8HI
IUgeVQjrmXyTY8Uc8+kYC169AyXXa9dFdaRY0aBKGJ7E6oAUKzz+JbN9Nn4QDJgK
3xFi+2d94IwaGJjOMAwl8H+DQgopMxEf2C0jlH08/CuDry3XcjQepSY3i4al9NfB
vFSPRdQ1cPPvKrkyy3JhZeOvppYJCyik3VdOjCNwJBJtvJBrABZzw2o4zp5eYbmj
xXU3T0WjYMXS5TXSKvxzmbTkeLPLzfkfQqdAz8YV5nJ7Qtp10SssRnjV4Wm8xed2
Mn8vPAQQcpvX0Pllhew2ky7xJmvTM1Uah63Tu2a5/g6PkQBnsQ14RtcIM4MfYkyT
9pcG0fPQGv2slZoA1pwhmv2qoO4iW2d5BRJnJArComThhozcO8+CQXhM6w23KkCV
ADvF9YamPYwQu49UegyCAU4scsw+a9gbVzrKeGnJVaZo6Ww/qUQJhI62ClzUkbDp
G2XWyWiZrzKMVlhhO1zPihXKzi81wLoM0FR+l2hvqYMA+hHXcGHXM3KUcLrdrv4l
YerLvM9zssH4abi1mLTy4+gde+ExaRvmUMnM561ZRdETrBqKf4LyVRRR3CO3AoMG
1Bzt1sXJTariFL+4nhrt+Lxe3a5a943YjcBLHAdzo5FAhfQg5kx0slC9qDJhJml9
CE4m4VlcxpitsqckAtZ0XBjcInaqUk2T0RH+pPtPsT8VUmFJ6LZiTQD/ZBWbN+vt
b0nH1bdd3JBMnOuKcocVsvstwKKApQ/ZB2g+ZdCDk81zulAnQ/MWtYTKZJOYDRuB
5Im1PW9YKPyGHC0msV5DpUJvAS6onyJ5IhJV5peDUYFbAdtTSVj7JofmrRMLjYcQ
QB5gOktNOe3gTIyL1vKqDQXs2ovxeUDGhSU+B7pehownwdmtRWPjTay39cew1Q/2
yw6/5qUoRJHOjsNmOOh9uxxhUrKSRuLPyW1YPzgB2scM3xK2C7CRDPiNjwqS2OsA
kf3LTjciI4F5FBMDYnH9EQOJ28qLZJ0godPrebv7WYkZVXQjNOUflMyaIChFMNx9
hSxpjZ0JS8JVPslke9uLIoj/qHGSAP45tT5OBsVakcElvyoG9u+dXdssBE4YWJ54
r1ZnGQETBr5ZNp2CGl3oHapZ71GiLXnLVE5zarkRAXba5+xNCCPgHSB+Bk0lZAIt
DujSekR0ds66c4+2ihKo19L4FVvtPtZqerwFCqndEVKoqorLvWmaHg+/X0plSi5R
rD7wJz92yUqLywk4XChRQqoLqwo0XbCsoDIyDVH6dmjcrckQDanUEOTipVbUVV4c
xoPbvI6Bn+eAJz7veOokR+uR4GZ8cYRA2xhSYTkCrVIX8yKH7JMWAS6jCFKQtWAy
PKm9LhYA6EOAe7Q4jNzz06kUhPo6mrZE3b9OnCeWUVvTZFdaI7hdMFkWpEEfutlW
JXg88tatw/uhV0qRSNQMkwKqfn+xSP8sHFLc1bCwzeyzg34PQewALTi9jpPcBgTg
9qAxrWeT44hlPGwPtBn8cvMxwHJLgIK0n44sgAtYKb0sMX5ZxBu3pcsB7YaFquG5
5DiXqezPs5Pllz4mA7ju4fZgKzwAuOIgHg9qi9I2uUfRhNcmfSpbkv8CDLFe8YzT
SHDnNRrnz7X5QlsrVPlmOHaNG4juXahTY41Yb3nl8qxH/bIRpnNYzsp+Mwwh2Boa
gYy/2ocxivZDqUhV8i11V8JxKZZNGrZj8KgJEYsSV2csQxLE+psa/bSTabPWzB67
Ov/DQLRpEAqePK+ZNXkTddvZQXzXe1uc69bWA+IUyT8H/pRg0PjVYtl02LGp+qOz
fPXGHJO/Mvn3tj7AJ0ANP13c7AlstyFWMTLmMaJkW7JUelHIRw6BSYNSUS5TZqg2
HMQQaGrl0OenJPOyt7BG+8RyagTMJa7W4bIAlUNNAoK2aTHtMJmc3H+NlFb31D/j
j3e/Mu0R8epBNR+agbHd4do20eTPUptiJ3l9fxagyNcbUyNTleaiaa9+qkfr4HlP
Cx7rvYe1CFz1jF/+A46m/p1IHJuTDb/HJzEQlvzNVfKOlpMQAWy69HscofGpKfXP
sLHJMbUIVZPeKiIxa6geslsA7XadRlgo20JF9J3t+oFEvYLZe3/WCZbCtC5osTpz
Zp2Cn80VFf9ya7b54ol1hpSIQNEBXMSknuflphL41b+yTx9HARytw5iq8e1fL8GO
RJxKx2T6B1o5qnpAbyB3Ow7txoFe5IYySHlNeINGhfnXR+emOyIDDr2mFB5D/Nh2
FXhKPDw6oOisrzO+MiJsiY3vXP4LReiPORCFeYVDkf6ZIgOr4yA5X7jUso9XEh0L
VC33rLca4CASIaUY3d2mipAjvq1jAGhayIuWnD6w8SFlwGsQagWJckAdl4maF0gb
bqTLeJFdKngM6OZlyKqRaH2UsgjbtXZb+8wrNqV3pGJlJSIVd0pYGfgxdpM9i+gT
dL+cLC38qwp+lRz2LTtyQoyl9z4COzWiC++9N+6LjWP9AJdCmGL906ola5gLfTjj
juXXGolQVQ3uP1nIE9nFTHw2uskbcJYgOf+Y2xsVvVJHSnMCwonhZhc2dODB8UZY
O0twQgKL6T/dF5RiE9nXrp4+dvkUeMSaWdq+x9xtXWwy+7PaQp9VPwBYv4oCBDlw
gj1FIG/qn84tMZ26LuMCHQhCMpMZE6Rv3RUlTvmYqFz4JVKwmjEH2OPfQle8yMTN
KV4H07m2ktoiK0195NH/7r4uMIMEM9aJWHJoPx0m4myw6IpXnWEGzyM5hqN/cjED
e2DHVIHYHCJmTYPfa6y8RCvLbBukonXQXl86CLvoZDLk1nLTg2qKqRjE5u83N6Ta
UYUJTFlsd7xitxgbjxyhB7mZAuWPB1ISdz4ngA85s1LqehrW1LmzYud984K6sLMg
5v1kTeGP6megNL7umANRxh3VmCpZNUOx9XwlzzhXRrglzRFlyppLxDp5y6+jGHrV
J0NAGsZtNQIqFtJy1BPl9/WvAIUPCIY78pDVjH0V9RM6Mp4RFj4O+8mjupAQ0skK
zzWVr9DgggngxEmyr1ehyjZo+kqaEznTj9I7Ku4CJ/V2l2QN37XtLiuVVqj0Uc1N
hpTHxZ6a1DbLb3zX9HGN64GOcQZD06QmFOit/ySbAAvugDKvQwN5HPbcpZ/fQPgM
r9Jh3TpEv3SUPhc/Sa0q80dya7iltX3tTl9HIEGne4Xr2Oy//JDgy3927RsovBD1
GpS9EP7gR/Ij84+DH0lL/VdcEISXYk78+Vs3FTHZD9SjhEmlT0ihG8393/STSoXb
yoL8fKr+3XFh9AIkGIsB/wD5QLHpQdFB2FCBx/DiAU2CDVq1snvrOnwZE8m7C51Q
hOxXdpzq2AgTLEV9mSAgqAsfjQVYgcuiYQIPQ06zPt5dfaeR/Wgh8JH0dacit3V8
m6FSGXUXySYlF8wdvWvIWuqpQ96kEM3BCyLoathAQfXnBFrWplS2CJ3ddplngrv+
2Qgbdb/oM83VEHx6uZCWh/6ZsRnZ+YjSirAivbSu8bJrfsZRfDWo3jzaXtKNMQ3T
qXtyolG0HtLPgrq5zEb4nQSt0B5eRc10ro3mpaueP3ibbTFY5llINptLbMQL/LuG
vAM6w53Ljb/KYzDg9CnUeJ/S5/VN3ZSq9+WQy2lNREB6xajaHyuVJ5M8RZqxstkf
+KjJBoMMiVBcZ8ZUZvth6deIZzrgmYhoJAuho/H+GTyvid/GG6Lmg2Z+FySA40vi
tUL4JsYCDiEvKNrJHuYTo5ZZH3fLEj5rlkqgfHmEF4aUq/y5MVu6YLzNvpxB2zDe
5BCoCJnMP3+n0sDjuhYHgfvYE5aa7tT+rpsCOmm+VLFlbPnQcWqt4ewmJP2rreKf
vM81GxCpgNJ4oWrRj2SMRaHJilATtMsT0RjhBpADCv12VY5wBefJUgj7AboMgfYE
x89Of5OSVVGG/i0UTfe7Dtrr2OECaNKpTW1OagbF/YcF8DvBb5wk0AOXxkMTrV0R
jfhdyHKDNxAPB5ITkue+AoKjYRskb8xHMLAenYXzp40fFOhTvbCilm5v1PHepP37
mFAcZbE1AfvGoCc+YwvRiurMtTDxUXARKiHKc/WABQMc7+xFgC6FNRNzO89DDlYm
bqxZ6R4tlAf9jTyT7PYUu/4yJ8m/bBWLVUJfuSucGIL7wfnen9yxPgBnCYb51egQ
htIG3ubmgbFbosH9GradEJu4fFo1Wpw/N4ASB3yB8gkBCNo+goRF+mAvWMuj5fkt
tvs0LUs2miTjkFhJJZskZpwb++rL2icYVgH+MkGkRQXZ2TFTXjYiFQl5AqOlwV4W
WK8/jutW2iu219NgIk19InZzrEgsupS5ceNwxhXedsSXj+KZC1482H7WZEoklVPJ
FIBKt5ihUUu714wiT6j0tDXwsfOIPcUdWrwkEI29l/iP8AVlHBYUIF4oW+6FK7AW
152XobhRs1AlazQwWwvfsGyYB2syd+VmDbtCn/DfmWMGX9fTlmcdglX90qCrzWOp
MW0kTGCZszJmGP9xXX9iQcp+31C7wz5NuVeU+FP/IF6MnpkXS2V7G7aN2PgzTwVJ
iEyG1PEkLAJ5u9EaBneGZzTqWKJwiNMAgP7bWD0hGTx5067uhxnxX2Yp2EdLRkTr
8cEGx13uBM7o4wQUepjrEN9mu6AAtG08/17jHcCaxZ9QnzuTQfw13EWcRSF+s3X1
py7ivWOTSmN2UMZkyl1IMO+iNeW5724N/smqEm0ZC+4lcbh6v5saOGyYnfdj1I6L
DVqZLYlDoHNDt9FI09eAdL9CatUtLG04BfcpwnwhuPcAqbSLEvg4Lhg30DX8HvUR
MfW0GraTIc/sp40YTRAv04pmhTDhISwVBee71sz1YZQpnOTTy1eCmyTUnKB8ngdi
QTSjmMMoAf/vgwqqoXA0a3/6d8Oq6Nl68edmgdhc3a7eP89M256Yf5aXELHVu3Mb
8TkvySJSHaV1U1XAZnFLhA5drOrwxxUkE42MAx0E2PZ0A5P7q2mHTYZFMwXYMBJ+
LtKZUN34FY5GjLLxStZomGIqQ3jldOS5BtL9BL1uvIipe4SW9TLvXFhsFPVJU0qn
2ek2gS4yG9TX3QLDcye9QPTc0Nb5JGXMUctPaDCHnYtAXjK9FKSSYF+eL4SHcL2F
jYIBST7gd7Zjp8rp7s3c9gIb9ciaPgidLjxmfaqsOJvoZUSf+EUvgExJC5k7De3f
44GckM9PVuO4wHovbMWoN0E4tS8gAgJDTA0HRSsnILIp6i81U3q7+/fSsP2U/CL/
/b1w92UK6OPOH+LpdmQhUH6LDat7MtLLaZ9pWNBHf0XXYxwpHvLr7PwllyxIH8OF
ww3wXoPaLzNbVBnCaCeF7XKQUxg5986BYp2cjDeC8mXZ0AtsCAZl+A+PQhEM35P5
93nEMT9OIZop4OGV4iZRFH1FxlZ/I/bwphRrPQiVmoG5lIkxElf3EVAjS2JwmnBr
56wvhsCgZhrbZAG7QJPNB6Yuqi+oXpVwFwykEywks6UCXSmII6AmKHUcp0ujcP2m
bEdGxfVyhL1JW6y0/h4i1GNaKwNZ94l968pJSH7jn9FRYPAnPnLjj/OAhu+TzIaT
HsCygwjIXymVQylNsS93FemXzgAxqBLdUsLqglNcbDF05NyHndFFmy5skLhLwlcl
GtzzIM6pnkLY5wmP6Zskal3aReTtVELsrwoK760RPuQLBLVNc8NhndRIt/N5JOk7
sJsulLNx1KHbBz5YMj+2kJPYo0IM4xvIsKaC5jJoUskgCZhK5fCeRwkwXtwyZB8U
1qAgt0jGC6OrfgAGgiJh2cLIs0Z1yUqnGXDR8cNNJ18UX6wraqofBM4hGvU0vUXg
TljMfwywUAW4btk68yoxS8BPfe0VxdRxKYgVzHZnxlac0xBDWul/B6dF9sQcgN+z
b5FPkNeuzw3xh1LXxuQgkU3QTHHfK4NnqQkKE+DPP/ApLDmVuqkRHNJSSsTbywMt
z2p09g5/FhrP+HepcqNUU98e9UkHJI6d25uBmr5YaYWcFxTiAJh9XPPunLGGx9vW
b1iE8IrVvUJXyruHpwWP0roLRdxe8LFOVTOEaUdz/LpPMcorHv7Y66nF0m/vdHQs
7bOQ8LeqLhNz156ORG76EpYpx8MF7aih5W4+yicSwsIFvc5blmlKaZ+bClnzPube
n3aJYzM4XAdhh5TlJT7Q38/tWVpkVS8NzoogTJKd0/7gEPAm+Gyea/Bo1y4mQ610
/74DJp/goe4nDoTs0tMi87S9ykjWlYNd9aLrqps0bsxJGljWmXQ6iSnOuOyeCyM3
0hsQPOb2IDIQ8K31E2D9uw+XSSKwXcmFzdN+UsVzDsDJYDmfU9a61NUqlelvcXZQ
QadAuSSkNJyPe3vD/r10RQ3OOqP0kvkhOnQjQvF0ucZqGqqdES70g+uSuytFSCQ/
fyz8J+OlvN3718yvq1sl+6T9usu0Z5fMHBf2j5whTB0m50Jdzrnc4Qtyxgiq/uNt
i3uAhfod+Wcw8nW3jp4Seo4i1zm0jnC02hME24oTABo60HHjrHWQzNNDvmenzRsw
PBhAMYF8AoFytcDmiXia5Xa/f72bw54Ni73sIQ69gkdZJag9TEQgN0AOTxZiMnbe
sGu7EfgkQQGsbGTAVfDK6vFuFAH1gHIXh15u0wAxsIQJK6EVZtGrNk52BHjC/wps
4T00Q3cVs2aIoeuOM9XeFbNkSIWbgUCkdoDijwFdyqEnRWmYt32iLfwEmsxcdKgW
KaQf0HQzVJ6EQSfWGdY7c4BO0dE7Dp7/oKdzN/QTd0iO4KmwHEJglYv2CZjdXB2B
hSYAx//Hv8zj9O1oq59l4P3g0CCgg9cpcPjvysZJpa4a60r2N+D95gNGMFgFxNtQ
hLQv+SkuJJJCqZGgNUiT+gENNvXNjqYGWg+s3FUFJ6drrETywCsbHciaQY1Vl5V/
VS5E5omoqOfe3AiHV7GliWJRDnC7QhCpRs6MPJdKasLLLaU+1CKAwiEx4KWmG2fJ
fihLu3leR6dfpREB5tTV2xdnowC55TDh/ImrUlgb4Yi5dkXESkA+KncOvbrKXZSh
s1WmHSxGaV4EVT4/VBoilI64GWWEa5pOAr7yr9zkZIb+d6PZaTwulBsL82dt8W4k
rHHjixfnNolwkBipiGQraVig8VaLkRdbvjx4+Ydqf3kjDP9HOY006zhF6cZyIvpI
tRs1p125552z2a578w6JJnXAjVuIMJqkLyKl5iS8oOYy+7OMO8c93BPggaSWSJnN
ybsySWn+IwtVfHvm/KPgCpeNdOLIrFNpVXFfTGzTky4iD12t7eCVsuFPhVsDUd1A
+GkR69r42i6B2GLJT2uaYTn6qdjV9Y1sRsBlXN4vq1RDidb+0O7gmsetqF7Yk30h
DBENbqpJkKNBDdvV1UkM9HnFF99k/yFIkiKi9spQLCm1MngAhHbjq+l4WcavXF2q
RlE2unagQw4T+bMRAENsNUl0NVu7siZN1NfwB7l92Vb7bxK69d/FbSihjymyGRwI
d3kzIQ6Ocr8ORDUbPqNTC1Sw9uHi4CzpNpTPmaUFrcZX5DCcV9wKwDjvw7inPmdi
okJkVlUK2rDKtDdQEDjF0FBYgwUUpc6u+dyaPDQKlZvediXLXIDxMIwDHO9xvwXE
kPtQgTsBO2CYlR5C3HySsH9/eug8M4onmELuRYi5uXsPbUuI4BQrR284aAW6+DHD
YPIssELh61rJhvVPHNksgCo6WAhKksjAcXTYceqjivWeqw9kKaunbSdSfo2Jn3dG
f27V6YbrmO/j1Q4iOCrvFeVEmRNPvospnVgFuBkOHEhDeuVB8KlwV+nPKbUMWstd
6+73YsRJw9niiUmibc3iir/h90zMyNjNHnHxPg42YBihefUbjNzTcEBeEadGSneJ
dvhhILPprEAu12SZ9OoKzbiyNwnltkeIP4eZNq/sMieRzYqkDDEVHau19rAu0Xth
cpJkeyvA2Q/E+3Wb/hQ7+08L9cxbHVZLzgrAlpbLlk0bb7wujvVZ70n1ai3f60V4
p3WfHcZiVO6IhtfsLbZuGFsohIH20YzBmv4qlIcStu39urGNXOwyO6Rbq26NprYN
jNeiWkKp4v6jWV+LM0oOEX9Lrr88nOBR6ZEl2wHgt665VgXqIEtFAE6JZRzpPuJM
bw+e0CnBAWzU/NXnvBtUUNsdD764pfP8gPPHdMXSZhj/y2hWxYrkmFqrk2TX/bYz
FhfsyY3IJeaJZfnFfhUWhLzbIgVjgGB/txjs3Uc/HI4N6m9875Q84gvk0g9ervzC
CzgdXAa4XABTTR7e0NOsfIw8BbUIIdWE57Pne26JPWxU01mE35E7C+xHVCyMFHFn
Tk0ra9sGHm5+VNmF0FG7q8WCQaR5eRnnxrFPth5c7D/jPU65xxWsZ2PSriWb2+zg
Y+i9ZepjxHdMVncTs0SrBciS/qOWAHFtkKtb19N4e2lKMWkMqWyp5RkwIAg7bL02
tWbNx7c2Zb5fKqHhhDS7rcw3GIxB0Y4TEYl1P5S2JQij8/zpHR82zZGXxaz6yMjm
LEl3tUXFa3dOwvdDfCuW7D3Yu+ejMMZyTw783oj+jlLsrraRvD+t7Yi9NI00rDZP
7krZjab7DV6nazcTPhyMkjzaJv/KknYDBl+HFJniTkjrJvC9RgxDznPCjVB8c7T3
zG5Yny9W4MQY72xwjYqSw8hMVpSX0rbU/y6DjdYsi/drjlXLfyPvgpMx6FkzcJC9
QaIdJgFoUkrjZLj+QG4+GU8gXvHxRREUv99Ji+Q/rpn6lnQMHv/t93DmZ9CnwEXV
Qja5MHrQn88udhTr4UXFhplntVdqLwacoP/LvKLqEtzQZEvOftjvPHKFick3e+2g
jzA+1Z4dEuWHWRTTzf0TanwDOMSBvbvd1Qm3wj9ss9+GxLntYRlVjLHVgRW8xsnD
/AXFvKsX3wGSAyb8ug5DbHNqsh0BRtW3WMWFdijQdtc/n61EZnpwJMsHSKhueYCZ
VWtmArMsWPvqM7wzOoE/natBKG/RuVT85ykdyiOlP0t/pNFmugz8dInqGkNLTg40
39LvCwTQatZAsU5tIxvoYh0sqjbuvLF1gopuHQlS4lN+ACLsS12FE3Ox3mRQN1L8
ImR+OO00e2E939lPXw7tkIlzHYAD8yiqtJtQuBgISRBkt8r1HdPG+hSWME8QtmaR
aPWHU4vwi9xCQph6/BYwkLxVBKd2h8bQfMMHwt/08U5j/YHvEKZf9o01wu18uMp9
/KBXa2aM5mCxo8n8Dk8XZUZYqbtwKH0b/bP7ESyBR7ZC+a53FZQfOVjsaVvdTKYY
65dL16I1CThI/oQaX3okf/VwyZzS32TmAF53R6hDeSmUvj0OSjNhVXsUldUlGahH
WdtLG9bWpEVK8ALSwJfxj1ZeD1p3rnuDPKQt2Na85kOyZ9BCBgDFG3fDmgMRPxsQ
47EMoJBtVVjRJZjhV1TuK1ncfBXdwFM6JOOavLqRFjz0Yci9x9mtpM16Dg/xQ6SN
WM6SGZXvbP6fL8i7aLs0VZgA/BUMwWhMGSfSqVvRakIKFPnMsR/XfmjGHMV5oPTj
5uW8qTinxzJ7tiurzVV0BJgNz4uB+YqMN4rAHHx+/fpYTdWgqR5ZfKWy+riSlaE6
7yIFtSCTlujhyDe05XUAn+egVn0A6Vs9+QyT0rXdx+0lHnVjTLqRfEGVh6GNQMK9
mZs/9A6mEfSoQk0dA2CqWHVVdXcaIq1dyG/yjfqlJu9hpe25H0m7VetPzv21XLTu
itzI9xhej/eKg4P99TuUUO4ltmQa53+sgNE26oGbaxN9dshpOY19OasGVOPH3bHV
WNqTXQhv9JJKnmMsKcJ1BLcTUSl9do+wbMQRa1AWK4QhnHCI2HAHvxTZMICw2DVI
n0pralZP/uTBwby8/gpEJTCEYF+JDPRaAXKodEuduC3AGxlltvtqH+5T4k91n3de
yGnHFR40MFnUXaCuwqMUK0pOpdsmSdt/x5vOEkdAZCfZE+xLhFSiItGMkmm1LGV5
/YP66wdnlBrE0o9sg7SsmeXdSuwcFeI6V4eaEZgmbbCAlWGs6nDnCBu2KXtJlg75
wUZ9dSnUl9A1aQuepcsp96c+/N6V8vt5oRiQmpw3tI0KYyRnKmYQKgBgT+kYeOmf
lXnEewm5pkO+GTCLtJ0EYS6XCCNSTR3UcpPvwvtcSsJvgDr704WwIgstP631ErR0
eldzw23eXnMZ5i7ej46O3Fy2RF1ab2B4Ljfn7jRbJJ+XZSrrj6N4tIX+sd1mo5aG
lItqvGb+8V2CFrCin6YK64fdxjIh6FWnalh0R3dkgPxWUgM1fPjin5pUDiUOjhVN
0aAUdZbRshK+4CvnHJ3Cl7oFheCFo88vpUiATptln6gi2poOn9lTem0x18/4JhjW
TOLYtr6aM+3Bp00oeLZ/AK3Wp3Bfv98r9SbUcwnui2GmwnXE+JAWR4f9vJLV1jdG
Bgwr3cD8zO8imNR7eBtttzv7zxqRpcaMfB9fm2iAf/4lC5Tl59RKyzCT5+c4Ilrh
FNPhVx5JB7yvqWitYJDAbBwH3DqTZMXxNfl+VGUAZH/3nysKsNbvUNKANjvCL+7i
5XBmZFXk/t8R+VvDZ2fAZpxqxUpRbcoQBxRD6qndKmzBVAn/Juz13mpLDZxbDpcK
2XRV1GEqK5UmnhD0d9PW/RA1mJIE+lIZ68CkSKxhiXr22+6l88vo5nKDKXnRUFN5
1enmcpBTZRYjB2nWOj22MebTi3VWAQXL35KW3YqWAwoomQqsB9I/r8vdQMkccNT7
nAoaToHZHJqPzQXCWvsMoHHPnZ6Ss0xz8CCXSyIxUJSPxABiKhq3JAgro3ofS1d8
sdqqTxQV9H2mal74RnO/94oNd+DHfhVkKRJvSq6+MxixhVVRHhUBKCdhGnV0IzXy
dCaFDFfQiQyq1Y4qUEEnJYhV+/TqkYka8MoGLcLpaW5fT3R2q67PzzEP4vz8icST
QEQW7b91ketUrFt+T3xF902n2piOAYfpCrMahqzhRjzxZgX3kE6cpeqJ6MWu74wY
qd3pAHmjlwMiY2QNu969wkSQSpfJZ6TZ/yVpAPPdq6ljcBWRaDC7gg+Lev4YIYmY
LEu+NfCBayDmqPVbt88+RamEPKky2AgecFRyS9r9NKZux9EZw+ar+yXUnvIkYWoL
fIbMn/mLcoVObAEfmDS/ZvL+1GO0126x1HzVs5rSPgr4cKmOsHT05bcNh6xXPNMh
1nvs95SM7+0QcL4h/aXR7DOOJSGY4QlRpOGu9w7jKQuEJUVzsmY4XvDyfH/U+hrl
HVrC137sMANW8DDljUxqSFPnMUv9VYkC/2uaC+kDZI/6PCldx4aIAwrcYnyvOXY+
pW2py5EL8mF2R/Hg0O9bmXge/c9Uawok774e6bBqIE1mgjV/0DBZYCIK6VSSe2Ij
qdFabeXz9DkpPzl2S0FxLp4Vd0WVy3EzHGDpYqIeQ5MNS7aCdBmcpAUKrnTzSVby
7epByqW+sgyj7uq95KcJq71Nd0JPwiDhayhZ23r77mDy+9oSrei6t6/99VbH03Wc
w76Cej6jJkZvMA6lobgIRwycc1oVibh43tNZTaZlfO4AGWzeG0bsfvCGJYorzccZ
QsMkaQy1y2uuQNCBNBZ6NOzE34aQL2hlJaI950D7URt+7vC/rBSknrLZf88d4hyo
vnSQmb1cQpCJMxlytyqUDCNuBn5R7LsxZiPcqAeQIBHvzPcMqKREzZRB3zK3Gcfl
m0ANo7wUWrVKxtLoEc2pyU66TU+r7lp3QR4f1Aidvi/gwb33yiMigbuq35ZZi6bQ
WHIYtHUz6tC2paJr5Nvi8b/6owN4iuUzXQfJIsQtyIMuKbt5pK3FNXC9f980DYqT
vlVChDM1L7uFXGBhCJYEiB4s7/rLR4eAT8raNTAaCq293+Y7AzPxpPAIOsqd79MY
k4dSWidRXPF9h5AQnVnAshb6ykX/ujUsB/Md5072PEPRI1RKusd/tde+NGjs+1qe
KvxLPLjW1d7Wqe5lJFS0vmWVFD2rpnxu2ik1YBR7tpS4IwgZYzqCNvofaWGDjxSC
nxg/qsvs3zeqdE2Wcr4umQJ5KZSjQTiOGCZzvDgjgKh3gkGbC2D8PURRWCqY+wyL
8YH7g6CYwKAiMbLBmcG9PhjOYn4LAlm+FPAhJrFwIFpdJF4bz7ngdVcvJWkUHlmM
pG9aHY3Ytdg8O2DQvhw2JRyoCOQESzCGxPNlVISIpuqf4EloA0N7H3QkBgkdizG9
4BEZKh0oE9QrHUPVm0O16rChIJFNqJkvJlsx+BDWZRGsvgqIZXpW6HlQ4xhWEgNs
0WLZWYUNoqucwjVmSBuWxvycFr3HfAzB35l1qzi9KRRJx2G7MHECNT0PyirKkHAf
h0lsssAFhyqttpTrrjCS01o7ZDNB/IAl+vNdTX+f7DqOllzsI1b537roLmsiwEEa
XjKEchQTZ3YKG/S0RjaymGelJr6E8bQ0Vz4a+gPMsR1KfOJ/114QJ4GH5GklIDUk
juEyUpG0LJ+428SzjMf3JRFSZyYacL08mt8HnLxYm4+/bVJArLwQW3yebLo/jlVO
Ud6UvPY45PUIsM943o0MGZf2H2dyRgc+8GbSv/dm8Ro0g9/ELmOdKHk8vQHec6UW
X1QtNehS8vtuuiAEZv+Cnj/E2mAbaHsNNHa0gBV+/9fwX1un+GSxfIczrVpf8Xv/
lXbp+MNLt9hoDFjmvKHWTFT+vCemkHB5ZXDRfXAJdAaNg/4un1r8NVm6bCSPvkXa
bLIXRVihmowc9SVJDJA3jP9bs+5HqD1zPbwXa9WksM72uH3QTkP8nHDxZPeKWlD3
AV1vuyiNtTGaOuDoGpyntzRmq/BdZUZ43ra1QJHD2FQLVPpJ7aS7tjRLfa6C63HE
4O6MkLONFl7LOWMNWVXURXxBf4rWEyaTWh0atFyJVtzaYDII3BmHoRk1inj/A5rY
jt9dcybX66jhGTHndsz0xjWf6TpDPxnQtFIcWqaIxpvkM5BRSfITJEYw9XD9MONg
9n/CkC9C2NUg3qM/dEMIv6GDuVqQVzNbpBhJG034DdqdjTYbCzlLlZM3QOERLwKB
AvG47qMxfbJcQ9k1L8Bhnz/oIYU1rakM7Qva8XDNnmLO+rgg0+1Oek+DLxouPaMq
uLfpxXN4SQ3DViwDvusvp7/PaH47d5nzVFleKnIHBiTne5f55HNmSuIuy+Jvtrfv
rPOB+mtm2DwMzRFteY0zutsz6nl4jWdGrErLeiOhbsZ1Z4G6yHHSmBXVeLzIystn
tZpVNZict3uDtkWQUYBN6XsvLMg4Ik9fQAyfn5l6YC09n59IaegiZnnzBJJaOD/7
6z0vQkLnhpqK73BK0NnNpNCNJjmlYlHqcibgNcE5dIufCxk5TqO5CeTToRJnJR9/
q/2d3EcQ0MlU234qEMtiNzydjjuooeiq4hZT9C0vImFC5mcIA/TZ2+r8X7WySxga
BMewZcYREdoaJe1alV+Kd0uYmHQqa9IuybP8FWXhfBQgUw/hPf5G589hr3jMzkqP
GPM7zYuZvKk67N7vHcvb0INYox+nNhpFnMYGvvXlZydAEf7Jk+NW0L96VZTC4Tcj
+BcV5d6msJPjwWXN/Qs0/+qI33fDWyM7kQ52jW/GmnkJLnG74XzmkQwGDPCYTNTY
yZWrEt0LCSS/2GeX/W1dxhS6efndrnZwO67FATA47gXaJpuyLIVJi5U1+hNUdb0F
3PEzzeR8Jp+f4zmShTrX3HixtdaWKyB7CtzNjuX7LkRH1hdqPrCQwLOl1msL4Mqd
ULXAiEmj86LCHXKXmTkHcyOP9cFDpzbq0Vg9PpsFiGFSqwkeyxHhHhrY4vH8fUym
QDAkyHiS2UQofaOgUkN0+qpi3ewjvSkuGe/9OWIA5VfFD+cj55WYUw/VVY6Ea7Ro
84dLlaeHh+mnNBs2IWACXO4HmClBiWz2UmR6/afSuJwWqz1D01H5mWgwCGDl8mex
vG7JpuuRgGoymSaZxUvfuW2XpCDIacqfDgh6SFXgrca5/dhPTZADAoGaykLDqPzD
tCTA/rgFn1D4sFVpdogC/zzoN+01yUJyz4lvwC2oWWHnLSIu4MI567Ev+33QNtez
rXiMxC9y9a/4VMMF6Unu7LkdjjUGWg0TzjUpgB1MnddtTAFBt4e6Cn+0vqLOF7z9
gF4ajkac3+V2JEMCirjstK8UkDBBzNYizlnmm/eJAZp9susIb8drEDxakE/QYMxV
OYcqiKUa+M6DSBtzWcsPQNwiroHmrtH6V8wa+29nFz8RLNxopWyZWEg1b/gMXBVV
0vyGTfc+BYcvOnoX6DnDypDcNkbkiphqRKFqD+jXaGu0OBHezmTzyc4v7VQQ+XE5
+mbrrO3ed0Y14xVFbnyD+3f3ap8mD1xRRtsMRFRGfNGdxB15rW4OqypniQFhEjeB
mFV4kODE/77qY7XyiDbHp9pp8lZb/I4iwQ8cynLBNmImxVc0zE+kVPy9mFUUHkOr
TAL9wq0up3FhoBOwS+9UsvmJlWr8PwzH08Fsnel77hv0p4zia/XkDZAnN0aivzuB
PxRFoq9auDoc1a8kQ0GjFTopZBzyi6tFTlxJ92lRumIQykZTUh6D8csMnAtlJllG
PlqrVQXlGt3JGHW0IUmD2Yt/lr1voIRJtPgIjEHWOgxlgznJH8daHmCQIzco/wQD
HGXh/iQbAaK3OQ9R9e1woj4o97wz40zc7TWnb78O/wOODMBOOWLQ3O4Iul/XU+kH
fOMwhx2X/uGlg5NHxA+9a0+Ie/zOCJgXskczwesJ9dhmpLDroOpZIYF/m4T2X85D
Jkc+9QAX/ugW9N++aRCi4/vw+taOOmT2riGyBlWvkNQvpEOT5U3NSCIl3XPW0okY
trNw3cZZbgB/L96FjTCvTH1wCzo7MqcADet1METU0hkAyyaj64RoXV3LQS0CNUiW
zu+okoFQbg+r9msm2MrgTO0qvgzLqOOt32clf8u9Bec+W6Z9JMmyRpFTYjjfDebP
hLcvssYRVGOqXCm/ORj5s3LAt0HQjVREmBq7Ic+JSbNrSlf+VvqM1450yGxVTndW
9Gp7rVLX/39LmHcD6AVdKS+BdqKeDl22oaM5NBSORfmxsFSqByLHay7k25cN/EU7
3cLHTUSu2YnljwFd5wik7rroMcJcBULjWYIUMC+bz4jjZqV6FyHpopBZVuCvNaaq
qndPm+t/jnm+9atX+T++JzpFJPuyM4twne4B5bC/WtSa+ZzsRK1PrdKsZbIbIzLd
iArR6ukboxH56MjDabZhk0TK4WjnpAbAFWnpWVVXEbjdXwhFVSrcg55oDMrcwaQo
z31/Ue7cppRX2IPh/02vWVvu1qB52RW9z9GADqlnLP/fINRY0U0pnaK4pt+rEuoz
aoMN/iYhLj4W3S7+YnH0opzEsOmbnxu1H/LT0xcoiL7iF0mN2S8OYAd4AASPx+xu
HA4HzAx0hPorP+FuzGbJnvNs9EAwMDGSmdOneRT90SwUPf1si+EhsrU2MKf669b5
jCsMfRpqcAi9qpkFBbT5DpZO+YKLic/jKBIYsqrX1asttrQruF/uXjHFXm1rgpbl
qDrC1f9qa2H28q3revMhD4pPo9AW3ZoYv9XPlwnZK4gDA6aEOBbZ3KIC77p+kYkh
dqAA1vYWpnPfycJYZKH+RQYOaOEF3haZPoXRCeLR4quDxmaKuSpUIvqLvkhIrO3X
df3jgJ47WP3/hwv0hN/g5OXUXCn/pHK/N5FOxxUPhrfyd7f7CeDTr7/AyxwIE0cK
sMb9OHCo23+HVzLgokUM0c4ktWyaFuTLbIXTRfwes4+ofdiTawwIPGb0r+nHsih9
6xnolFg1pBubykj5CEQIuRcBZpsKPd57+TRu97fF5tOxqBNj87aeEY67lIQK5BJS
QDYhDJAPSB0Cflo111K+FlKA2ctuy/i+eGC4luLtnT3Zjmyd+GX9OZhB9eiNVilA
KtyN+ikTLsUf/RqaWhMX5SRF5CNEAhsijtJE8rQFjU0EszNaIBoVy/bShF97LrIZ
kAsUZvhs3VwWCuTEAA49ae+0Xq8l3dMBKd+1m/O9mgprusaa2YScVQh8AVXsObOZ
qzbKN2IEeM+5eJmmpWxQ0nMQW/NPhmet7CxlW8mBuFZYlNqqi0HhVYqWYsh8cUKb
QjtyeW/cZBNmMtS0OBSRf++X1+8A55zr9IiGLiWdYpUDFYXekmIAlcVXbuaLFQ2v
Za9QdpVYUVo5BdyIPmmtBf9/uKjYQYdf087AtiktxrARLzqMLt0MA155oYJV0iNw
fdgdDqIL4cxcfeGdblzxiFGv8rXsFRi59q8NOU3n257JyCfJeKWQ+6z5xpVv38LL
oHdngWqL5y9jrhMVj9j/qqBuWnRs2fZCheZMYwfLJre+tV01qtyeHnkVMEvmYe6o
pmZyE18u+pYYfqxn50UF5XdS1Fb7SYxqe+EDUZwTV2v9W4u34EHmQNorgk+jycIr
2F6I/DbVclVCk3Xj1jtxMKjiXOmXs3pPR0iQHjW6OwOR6ZH11rp3fU9Yb4SUF9pL
YPMFLxyGqDV2Ahg06lO+GwyErlLHdiDzz2FiiB1YYcOiyWJdrsCmk+8odi7oQ3fY
ZTOn1knsB58TddrU3IepAv17/Hsykg5u/mTCSxo49I9RLBHqycYX82IITc/SyZMR
9Mui+FcIuwv68hgOCOKEsLzVemf8gSCnnPXPr9rNNB8arbsDYYr8AwHv7r75RViU
gy3xB4bC8V8qhFlMRKoA4PHHlybmPIAk3GDX4/Nqb5nlWIaRSk7I5nbJfTBJatlo
u2VXG1iPF5hvZIS70ZL7af10UEd4oSzYkZBZ2R8lZgeArt57Uhz3tmxSdXzi0oh1
50Z2j7Rs3BKrMUx+7mvnjOzNp1ueh41k1ayvJgWo/yNULeeHHaHNuUl7SW4J1i0M
5kY9V5izVpaq6NiruKYcV8bsfHkuKxhHeJpupBoGqE2dIm813r7nhBYYX28X/xcB
xfBW80UGw1sjN3yjUOt+tnfwRWynOvShkkg2zievrWUMbIhIaKP0nrWJnRItk2UH
MIdKtTHGlPp01Gv9T2ifhbybFQWkxBjiNMJWj2+ANSg6woUui4QHpG59RuIc9uTx
tyyYzNEe3B6VvMpYkZyrzLvZLa7iZ7zBogKTz5ty6smAaQ7Iij/dHhuwcBA09GIr
BkwDeF/y8j1yjxLDQy47VtSoPkm8UqWbpSe1SlkkQQaEErHDloHTyTStQCrUovh7
T/dU3pi+oi6swZJDiHyAQ0tPXg+d55Peh/lLHrLeRIvY/uE9VEyXzgqxxmphNhRb
ucB7/7HTDLP/KrFY2Am4uUXwhxrHf/dfuhZ30oqnvHKH09TyNUBdvLaD9J044A8m
VcYsQdmwRdOoL1s0EaRIlJPejiNg+mO1NYUms/HspXZ5AnRVjkan7BfFT2bn8KvT
6QD8dRPkaGX/GSUbCLlH/+OMGS0ggLmXpnSdiIBCt/rSDvSsHgfKpLUoJKui8DHe
T1EeEvKYwuvtHTvzwNEfU9XeGqWL03XbdtrOO7AN/9e1A7VKI1ikTK+OANJhfx3e
alXEs+oyLbtxME2RnFCVfqjWgapkHu9HYXgzbOR2abC07K7nmh2SwiNe8rrYeayf
ve+VEULbeBnEaPlxmKCsu+alVC8GcmsH5r/T5Ljf/dMmyTKnIYmRHLVecRYi/w+e
DduHJACrrQ264HjuKGUqwxbBvZK6pgOp2fEdeWnRM7sm8w+gDnYUFJckjNRh1j6x
qUyys7j9/cbm2N02ooh5zGtprPUm6j08wInpibwiWX4parqWmT3r/roNr9ojctzH
RGFc7QJWpkYAunCofIO2+ptJr+ZdgSzCRoLPuG4kt7XyBQ0jRaVe9D/jd1sLFA6A
GtfF822WeWcBGVtMhUqlPmT6NzqNuTtxUB8eBjDNziWcS2ds27awRTaOi/p5+/6X
CH+JYC6Z6H7fKg/fAN1+haQrpiNPeTxowQJOHLMBYrfSooQj9p/3BXIrBzBO9Vqr
LbVYCPKXYdtUYBGHIAQjFHGLWoL+5jKLuRQMqSj9PTIQZeua5WKyN+i9Fr3OG2Vw
qX6/3sx84Uss4/ciGW2QXips4X5CjReqvgc8GX+Spvh8rgULQZJaiGHQzjbJ7Msz
TW6MqhB/yHTfcRI0hpR1w06Ih1eQamLNE7hW8MYgq/hEbSl/W8i7jz9WtOg+smLv
Zba2YDUMPmv77WXv1+Sn9hqdbU6sRE5SKE5C+OYuf012tWBuB5O5dD+N36KWfBYm
htWgFjfK1uQwKPTCwtxiZz52S09PDuAt47g1Z/RWRW3y2a2W02HLdEyPplE4vFDX
8LEjRV/h2AGwBc4/C6gL8X6wPyqhjZEkmLU2F9uj8TDe3LZc5f2jqMkoDhjUdIOZ
Vz1AyyBTrnLD6cknrwMilWEMUMYmkd651KFJ8Bz5jcgl2Qq//l3/G9Aba4fIN1IB
2Hm22rjX+Y60d5SeBh2BGF+InbIMeUxrdxRQmH08hP5dF0UiQzcP14JoTWUYePSR
Uzx9naIssM2V6k34i692WXGBGEXrhnRrSXwb12FlV/9rjCdklWJ2T8RHJYL2uHaW
GqxVvVY/Bw8B8FMCcYMZ636ySjAFJ2tMgConttNmRiSsQG35Tb+3sMcbY0n/sxi2
I9LPBoreAW8oJ7Aqv9tHvu5Jyunt/i2FAXsnyQ9vRTi6N+Wh5KR4gEX2/Hl3WDR1
gGi5kr5980Rnzg9zQ13dQwT5rmy5nh3kZ3sf8N8zC41uhm/4sI1FbhsfZgPSvbVR
oRUlHBP2Xx9v01fADJGhQpe3w+d6vhIVbNKzr+pw22ys3Kqsyq2IJgm+a7l3xzZP
uqjInbkGq9qanp19f8dN5zfeanU84iqQ8CDuwe6sWL3w6Ou7GCtUb5n8sBQ9Qzfr
D6pLG88NNemCo4paBj7OSPuaEbACF3RrXSzyDtf6aXAF2HOAYzXmd+SOZp+KOgDS
kIAvSXv3HJMeZQ2JOyDP7TtCMXksF0NPpdcNkXbnMJd0elAVrLnG+ygeVxQmqAOr
1OkTG19KmmWwPiK25OCJOk8r6Em+vFFu7MmSs8orF6wnGEBd6cBEXphfLoUXqNB7
/RHvKUNDulszQY8Vuv1sQCEow8seDtiOy5RDTuL+vLEKnCkReZwf3jdNWAywvyy8
RnakYAbNcio18T2R5fskxrlaNRC3sm4XA4dUoR/TJ2tWJwJ1fgHLUdEtUvVrX3Oy
Qlyl3TFve2t58ZPUnQ+qaxHOfKt7RR4YLo5PIFenxMAtB1rCe66+exluf0hc8Ii+
XTuDBTUkFVW4N3iPF/QUccYmHLLopSMnjVCL9PdkT6nLB94BtHXgiP425zP2muB2
rYe+w4J3+dCQpt2VFzOHLVfdEgndMj7WA6nCVPEkaIawEF3k75ZaGdQivOyM0gj6
CGUpQ4vibPt3kTa8Mfb/XAGVRmG6VySEkRyJTU07+6YkdVMTdr/8F48jRFasuYYj
alJxXL3MuPU6XXLh0TZtycwQD1OLmJxPQaEmdaxl4AudULCNjyh80fod8m1r5OQK
n6NG2ADjaKRtPvNNQyfAxSS7pyfphGFZqIZdPzo+vA17vIffiKo/tORRog8ff/3S
4yqDc/hunfIb7N1Cb4s0g4jjAHlmHxdiODdsJZ2HBVAH4r/g9BZAsDgGBvDJpmjg
abA4QQgd7IdJmeaysN8e/bRL3W3wbg324ITMCTQ5FPWJhjgYFmuGDT+gSXXvyvnC
CAEqaRMVWsfzubQ93R/udxb3Myo5QhAKzQI2iYfzy5lSMqkOAiW9w4TuR6vSqGrC
Es2/v93yGZ2sh5aJEQOzilLjp0cH0j1hI9WaMgQyL9G86whE+qaiqWN1+DOwtQ7g
j7GE827kK820xwLBGXg2QrZwlwXRQjltN+62CNlW/n96gG4EaUBVromWkBPmt23a
unu16k/hxM3C0SOi6OBobYpWktLBZppALmONW4GfgHRQZnCkNebQDizK5Wr0beyT
FFCEuiPir4yAyLg1dAGrGHMkZaie3ne2YqDlkIKXDwEKVgzjwr+0oreSDxF2Zo6C
GTTc+N0U4lR9YND7uQ9G7WjvPJ9fRsL7dp4E7l/reaAkvrbyX3t36FSoycDxPMXX
/EGNGyIIgFeqxSLeBQW8rP/lykDnOdXe084G2KpM7hc333r+uX/omnXADBDnKmLK
GPqwNMNlv87fM5ZNmJo0epcDlRTaQPQdCrfuJZgajhRwEYjpAVqcR8z3opG+Yuej
oiVp2eV1zUNOtyYYaB4wcKtcenvSPGSRqShi/KCxH9EDvPtoL7BRLJUIKJGpFWvT
KOZkAqoAKvy4JlrtAEMgoiAUm0n7pD9qKfg1WhwlRq+eI4gyCT6Rbnda8Z9z5rbZ
sR67dlXotjgveANLROc7VzAqMapSaPxRCWBfq/SuyG+sIOSt9iRjBQtS+v4Fr7Qu
YFMgi13sP7j+Bz2FXH867Tbnfv2S/D0tz8W1tnqd/NCotIzlwYQKm8pRJI+Jk/Hp
WtuISNt2kCUxA6wGeDcyVGG1JCPQB4dvBy3fuA/K+eK6N50WX8EA+RdXELBhedYk
buDEmCdnjM9aW/1JDrx3DKhgLuzQjopMkcfPgMIJJ02pPESbcbZ726jCI77lJ0Ni
F7GdWV9/RT1ATZ5PTs7VJJZ7cnANN/tS0Bfb6cAXMLss2oTFrEAcuwZnT5YJOAjp
dVPVvpUdkXJgOQOq4EPSOZs8V9AT1s1cOiL4E7zegDQgE+R6FbZnjEGuz+fsVYmp
gBQvDtmIngJQo3hOWPiGMrNDLin5/5cP6EBjbY1Z8ugU4b/7MlrR2RmspKIgwhqc
qAjTXch2eqOSrF2Zj1SV5zlDR4FaDZpwjJt4JXoLfGJRjgLSpXDdYveSW5/QWIzc
XGxd+f5tJKxI0usCuOpa24DobNyKvqo392XkhimTkwwiS1f68dDo144lDmhM3s6Y
zvLNp9kt8iYS/MBln2HIQq6MIgcTNPszqgIsPpcZEB9mJ8rDRwzZ1dRXcnBrcV+n
hlfGS+7LOrkzvqQr9c5p1rYhOwpoHnA4/8nZEj9KqKGpunDrtcMsvdfQcue5As0G
aimSkE4y0CVGBruqi/OMzuIFDAxj8QQ7fBUm03keschXTvctsf8DismHV7+XBo/r
5XR4Finp6VZ9sMNdVkraN5IQt3o18K9pJY9dvmnBmQTCow8U9S+UVPDsDzrAxf68
lisGWtBb+W6HFMG4UjDY9Mhfop7YfDXeApeEoEP9oyP525OTNb0sDLnBIAsq8i5q
22a8JHxDhaCBX+CzSlXsCcJU53XO/2MqUimQ2UBuvNouR1yRFFh2cpLvFgRhRuyo
tWMEvcvxZIQU/4CdG3UacyCYwJjRJylgxRKLwUPXnqbr0Hz0HUZDQwarjo4CyXer
o1YEKAOCMLkK9PSgmkICiGGiL+e4OaDrfJG439yIfLb2s8JOg63Z3GrRWn1GAGJN
wJ/GSYkAh95DurtmumbJIvEJsZfRXwLZmirpA60KM7jf8fWig/ap8tTRNLSO7ntc
CuhHAIDSvEmVDyNOtfjjuGQ174hlvMTeZ8AgPsBxVdorScExZfPW1tPgEVTvbmTm
dojlfXLa4GElKDMo9MpS5S6R+pfSaImVPSVDmWduB5c22lrHCdhxegQLvmMauf8h
SD7G0roJtdNphVc5/NHf70NAgSRollDRgIgtIIhPGsvoD4BR2yBevCUimHYfvArL
se5NtZEGQtTDPTOagiNElFI5HIz3Xk275l5EAswuUTD9GgAF50+Th4NhUEWR8M5t
Z0pxf4FN/xKfUFNw007tB6dfQhGpooneFfwPgs9SLd+7CJdiShj7Q74lhXRTDz3b
DBDOnr3VPUfdeiA02U1doyKhdFy6R4vwzXuxLDF+ek49/pn8++PPqnAeOWrmkBRR
B9HcqB+nPDVyZN9xzsS/B/V1lYTGqvZ5O9yjnMAm/X5Ncuo7kx2eJJgTuYKNMx3L
KCqOUTh0Bs/aW2KIO4y8oG+EqDY+2y3jieXUoB3ajvVoIKwHM2WIB/EqVag9gxx7
iUhfvRGllUTyxo9y6BVlYu7oJFT89q1SVOdyKiyCdusjk96G+ByckY6BsCQEQ/qh
lEb9vVCp/OgXABuKcMY6G3fd4+iTa6mZaDrTWK3bPocOn3yTHuYY0W2Lv5sixtVQ
e1NQsWQcdMuL5RCDcQXvvzqvu9wzW6/JX2ocm2jj532/2tUYDQo6abAWQ7Wo9SLc
0O8dh6ZPk98TKcvwdxGogyanoLklfSEaKV8VGbgGBotgXUAgM0a8FOLgbZHdto8r
AbsVSKcVwdkLpRehTGVHntJ64eQjb3Ke6f/44Rfvy8VWm8YLVB1JEl7dzxUD9FUB
hvw98mEXu0QHxUoyHZlh728xvnni9Ugz7Zf6tcdJh6W5QODEaAoaX3LfuFlCTiVM
2cjdcaAO9n45jg/0agPUdO4FyNAvc2fYxnYRuc18xqlgPyx7PHvfZNKdve5DqZWB
ABoV8+zeEVt7B4f2AqZ5cPH9xIfKruOH1nxQnJ3ZCtCLiFNI5p+aLYj9aRwZZZQ8
fohF6rm5nqidUYBJ7lj0EFyvbB69AGRAZUX+69PPpZEzOQRMBgkp9Fc3gdueD0cv
AKz1E+txf/2IEyw2HXRPsrG2NhbELrygIWg32GTiPgb7Ug+wt+lLCZbk5Rgw3jLX
AvV29aCgdIKJ4RKmWsv/LgfesgQPe2HITadPaNa6LKjut4BFetxP44xxm0++t1d4
Xx8ojkW3PZu5NnekJAM6FDkNks0v0Ppen3o687eEcG6Sqe2ViNJDp3Cedx2aPt+l
Gj+cjlFX5b+Qj8aK8iP8exmhfHwyuZ94JBpxrzboNgvMO+UhkpxYrrYNNllFr3Kb
TweL+nxxyRY1fkB8RQibRibfqBsFhfx4rSyqg2m2XpqJBgrMfOJ/90ZDdZfcbgVw
L33QJzOlL+Y+ZJV4yfEI1U7jMvJ/Osr3TGyqWGqFkrqajlvFhIc07HnzkAUD63PI
2yw0U/hOcsYaG2liK7KqSxFcyBF684K0OkoUNRjD1XBLKius1OfC5iwarggH8YhJ
7rUfadianqkvbS/6ObNjDNg4e07TZs3Os9NOO+vCxM/89h18RBrYJ+9babHaZ6lp
GWdS74JgLjEEyfznITsg72rztA72+PBZH/v6UBSprINiINpzkigSi+ONsNywcYdC
hWrF/XUrVTwrPdEd6oCKgjE1rE8uRDT4nYe+vSEznAJvBDHtYyUo264xishDHxGq
tKiEsjSrOW5N3ewVD/piSO9EoY2rnvC4hzf2saE/vlFa1NVMF07zYv6McgnHWL8O
Uy2b9w+7GDwzgYhycqvQyNa1N35M+e1SsiWQ02WOkA3diqa0CgMpUoNEkumZJjd0
Ahz+vKhpdrwE4qZqerMs+LxRB8HDl6EReE3etpsAY5gIgJVNXS5BwMKO6WrTuEOq
A4CeROg2oe02AUOdlCqBXrBqImgjk/4Z0/zxt9WgzPPvFpsilkCN4W7jCY7fHQJU
vUZWcw7nSQu0TmvR3LSaK+1jliBJn73WCZsnUQYk0Ua2ysTgImGzJcilpTOBCAyV
6ncUcbyxUlPffEJiTYW0ep7EF1CeoS6591D4n0WETbVbcDtnrUAuzGypAVnMxZnz
PkyVJIDRwRVzIhvKiPSSxKloSA5lNzyE7HXN4/3lYrAP6w8TvYdXQ2WWcgydC6R7
ErCGcQlSovvot0p3JrgfxC8V2LJYrvr/8GnXJwayKWMdo+QxgCKXBv77lqwv2GeG
XGAZc93KKf/0BEB/jYxA/HCgN26IhI18LdawuiBAio44Sk610bTI+0Etzck8MKhP
ZLAAIEaF87KOF91bzxck7KkoXQCfmEqsmdD+4YjsFKlXQtsecjqzzDjwQ1jZ8lPh
7rcxGXsSkZimdmzH5HhomoYj10pSMuB0K0l5IVcy57xV9CITO+65O1OWNKiqxQtX
EfCyHJn8JETDAVTrBndrK85Hkme8EVgUTpcelSh2DrIdXZZukzUIabUvM2KfvQcR
tbggWRtMNvx07yP3RKzw8WwCBGECdJWoNblHEQ3AMzdAyq5RLj3M2ysACSTg6+Ti
lNbXXWkw3yleOcuVQ/3Yp7nyHPkiBij/Te/7hMTnQsfuyYIHieqJbQl8nlbGCGhV
+ijQCWPqvBOIN0ONuxsfnLXLEbJsueG9L3zTjYt5j1JbfLimJiIENlDyub2no+hK
lCvoqN8NaPmVINg942aFKJQ1eAY5Z+QzG78Gcqots9jq7s5FrI7875Xyqc8bVWsI
ck+GVG5aqpClTzXIK1mMtzPsB5VZghGaHNz3zaOpZynccPt4pursYaScC8xDDcy8
S30q/o2rRwaN3LtkcNDTITuNRK5YsA5QhQ/aqxSviFsHBl9JZ2iXt1fadqIlrNf2
M5ZLl614utXBXKxqV/CcYbk3K0NIB7+o00O/dgDjKgp5B3AdybjokUgKqau9ONMP
2iBOhEKsiTD7EiRgXaWQgnZG2fmBLiYAbe16r2Cu4qg2RoRocuD+PF+ctMd1LTl/
0bw5TX+kMlYtvQ9MZDMgqZQdUJ7mdQuXvdro1c4BWoR9MsvgR/9HVXuWVwFoLm1i
P5wbAFsjSa/mpqBokuSlvylppGTIzm3oB5aqhq99FFRiYG8Bq3Xq9Dt3kGpxRXcQ
h99dQQ+AELOcTrZcfvfQgplvnW+cC5bN1oWO2VFVYRChogMB6FJqv+wAHQ+dn96r
x6OT1ULufmLaSf1xBe9Qb/7/EMBZLxaxgYJzY3nml+q7NZQgef/a7xJpDJIvumSR
LqmijPH8rEVupI/BJWg2g5+ail5m9VfZKHjbgJ4Ie9J22k6U6QA9NgZOKdLeQVEt
IQw90lfxHCekAQOdQBIjMWUrklNMVsoCRd6NEaLN2QQ/30s18tXtsjSiYUJneBm7
n4zNgNlJRQDnlsLOgR71pnRBWn/+Gnc2GYzQ9HEQOkhr+nsdedTTEsQGiIp9uqg2
wBDI1IWlBJWQWwiU8e5UMkMyoIhLSfJaFsJUTEObqL7dUUoCzxNGQKKRrLVO4qO5
9SlmKd0W6+0vkWQghJTz2x0DcTzYHQ3DPgpcTY/4qfYOd+J3B60EQwhbMVb3VPiO
uCHZqin506KpGs06h/SBjufQNTWxvTAl5w6kCMYpbyVCXZ2BJYAOoy6Dqg2+KSq3
owpsXCwJ7g8IANdyap+e3MbfTHDthyrvI5IKbPibXw6wFlG5UD5Z4/Y3zQAHzbiu
j+aQzcVlDADQ4BQCu27yxqPFm6Ec8JXF4eSz+l6pBd8KxPUhsF2S6eLdqrs+SrWB
WHo+YmGbOAkaUuitdlfnLzqZgldtCOpfbOIe+wWiaHb0Vnyz6DsJcBT8m6/nbRa7
jYVvL52Z45y4BezbDVzxWt6RnB9k2wnrj4uMmO0euqNnFKUkZBIT6OsXSSVNfbWA
gH14NeU+v88dBOamD35wmof8yoeoIezqBbOjuauFsPyEazB4ocrbrsQxP0fRe9/b
GPEFotRvev2r5BNbZVSu4spmW3q3mUiljBeG+joA8AWLZF0//1tbUg+yXZT2UKNp
bq3j/CQvFx7kbUzr1p9iuSTtp7P/G3WIJIbD+F/BS9ddru0vnxcSzc29ss2Qsxis
5Qu5bABRzIy2q9GLS4xp4zNOi6+eGXpuqyH/mRuH13Y24vzkrcb72YL82izSyG8V
Nj2lzvzOTlT2VxS6YOkgOfyrnJJ2IRo6+mUyjHrxovgjEbqSRrk4aCj22FaD1b9W
5U3EZRSZsf5y82r4nSc3TkxzbtXmHKjeRTVfwgX3mlWS1diMQUkpeG4iglKszIaA
6CgBZM4pC3yQLC6wicAsSWs0J7RsXH+rjIu3UhPbLvL8ucXCwOBYUIQV5c8rDvc8
4bjIyea1J4Q+LSQj+jJ5BDMM3M4y+bG5O0EOBzCbzKu5vpRJEpyxWeV5OMPiDqL6
1K59PAOnf3z3oAugL6Sb00lO5RlHp9OO09rySME7jDr2zTGRAJ54V4qTwcf5hNHy
ewdCkiqQXUqWWlL22DHtsVMRS07czCHIZhoW8wRcAYwMqrmpRWeFvdWgkmJiDRdf
BN62ei6UFLsZvk70XK3YlbAkklKkz7VPil/kVRNTKTZTLGGFeCKs2v2O/cCeEMgo
OC59qxBid77BT3/HBJa3xRbo6M/X73T/5Pa1eWvRToulvdeKUdAGpuWliWUdVXyA
UnMxmkBMPIrKb9xh0bc7V6mEhinw/LSuVVQsvsEpkjf6D4URaIWdRUcuN4yA2LEX
c4xoUmrAKgnkb1uptD13V4JIag4XbtwGPV/GnMJdxEudS5IivdDMw1f6uhgrdvSH
wAl0MHcfzMOuRg2WIYTN6GUrvbax5RjdV3OQYu4IgLcutpecNHxY5xJP0nqVEl7i
uXWyv/KnqAZkUdnXPzuINoFIGZrZlMj4Fo2zWimtLYU5rAY+IbRuqycDtQ+qdiBW
OuJCvIy4c4FsSRc5OZbQ6V5ZP/e9gLiX7Qp0d10pz/vUIXIaj+hYNVQAzrvPp0dN
dyTZMlRS2l0H1xDLpB9/hNOMz8q2kcXI9eG7fvxV1o6vRIqJLpEaJancqrRIKjT9
c/5eNdgD2kMvTUG3ZGeio0zhJ4dG7brSQC8ldzjJNapjUODW9UNJ/yGgwubj3gNB
AkXuGTawACeS7SkrldMpzXrlWIHVu6A27kpPQLalyZK9h76E3/67EzbShfTP/Cti
QH4m8FcnULs+JPULET0Y/x2LV/7EoNTTO4E2lK3yr8vLFel7oY2EI+D1d93i9JmS
kACgQmdz6P1aRQmz9gOauefyBcF2MNNEc+e8WqT+fIlVXzPESZ2duR5NFJoHmHJT
vdZkpLrxb/xitHo2mHc+ZWZogg4HYukXYAgtNxlaEJbRsmcaEcZhuNM7rvqu2YMx
ELl7CoK9pjyfWCLOM+pxhNH8wWsF3VXUcSQiWlQkRP+4t9aGNitST/iHExnBEuWU
Dc/+NGTnn65BQw+3NLj3Ia7WZv/jqXFliOvaQFsUCi/q0HA+YbyhWHUeUYxnmv30
5/QX2i4FxKNnQpjX25yWrGJPkhChPEZy1ueu8WC0c645tKuiq3SON0JdqIWIMvRR
31A5gsrwHx9y+3XwXf3mvDdhuF9k7t3NT/aMGvcfL0RH84vMlOR6qsdESiU/mCbk
dXxRIwOdYngWDImydfsR0HhsSYI7PpwAZJEOPt1h6OIe9DAMGYJATONnOwkCPAYa
iUysQpKL/E/G20xhiWlQv0uxtIBuTNsinjgR6ZkjBI7ovoGOINe0BirHQRPn2zpY
gb/rTa+MgWrautdTg5gXBstXCRMPjtvy20p8p/WIQFXmOXurDzLTEGRvjrGL8NqK
wUyWXK7bQU+Frps+RqqabG8bhmojazncAykpb7STEjfCx2tbOewat1AFkd+YxBvF
jNop+E4932oXk65sKh48gOBEBI53AL3IJQdMWQSS6LjRpH/QljMnikE1Z+s6mF0T
SgDAm/9RVf6evgPmSgiwaE8zKmwpVCTzBwXTC2tpTGvYGGU2zuOytBr1a8j6iWhJ
meCt+baDvm4pTreDm/95hoYt3tLnSFi8EE3xG2C+8m8/SIZIPlFzRIG9jYCVyggw
O1FZPpG/CZ7aqbMi7oZrWY9GKhC76Us0EjjxUdzsXVuoDm7ANu8W3kct9nQEyxe/
hHMDYBsysOWUDaCrmzCC9NFQFxyreIN5DeX2vHLcz4YDS/8NGrEJf7N/HI4lfkPi
g1/oS1A+8EncmnbzfjEPVQi/NIHuKgKQXfTEjSb+cYupas5Tw/13f9RuD4kl6qsp
Y39dKw1W+eD8rbHa/rxaWO6lY0k+YKMvz0DFy6zIik155o0TBmZi8OlmYTqqb5k6
3N9ClcWGzJ/eS1zZPTpRG1yFmTHc/nkpWtpC5yNIHAVjXHIjbpfRH5hDx2ZRbx2n
Hd1NH46aXAORZuPIFfywYE3ahfoVU0ewjjb16RyI5aDBqjl6su4Uq9YBBjj0cw0j
N/dziG+RRXX3ZsjlI8g4B/Vvv54dW0TLUvuqKjjLLCZBf3EwTfo+rdzW2Obwyfc0
gnwOjDV69nolHFmJ6yzDjxiyBn7k0VBa3JoCm6pm3au+E6PUPK1/ATgqnHSHwnW6
ijzdsAocy4OLZsa7a9Txw0La6jHVkxKtXnVDBIaWeJ+kQbAfKbstHkqfRMmvk4oQ
EsJAlarcPdOGoUympTR/L04HcBUe2vGRRH4sfwVxvJmbfqAp80TEINCYgWDhL0BM
KovD5eCI9dUbspCAerTUf+bMARWUl+wRdZOwKAWzXWXXYvxfvDs5pFIHsso0ILpk
6cdTkKH8rGaDrO/fyujFBhDU9lWw7XVQBD9z42MKhnBqnDupRQ6uQRZtDx8kQlEo
CZfE85Aco7wMyGQpFCYSVUW/L/lomNRgOZlkDrUatiGXTj5HIJzissR51Ku82Rf8
ZZxV3Q1weoRrxXRP60TjzHuI6vYtJ7j1J8DPa3MzF/AbCDt/JCWuluk1lQMPyYS/
8KF+ftlIrAmRUuL1apTQVKokdsQdcJcE4a6DACzv/6MWKrM+3zVhLz5CLBpPYCRH
VqXzECCwNO0XkA+MhT3/M73h+DowWOiMvRrL0JB4ShYOwq/468IaoDNDtmaEvx5h
RS20IB4cPl2NenQi1VR/lMbJHEBqjTlK87mB2Z7Z6UxlJe6NMfUEg/Ilu72X1w1v
dRqzZ8LqAU9ahrl+bmsvxDPzEX5we9jFNw5CjJu0z4idvTwLQBFUsBjxRtUsHaSK
sjvgPY81FNHG+3xvLI6x9uufHwkYVpAyzTFKZwRF/n4a9TqFKrIuKkQW0xextRYR
UWkFOb3x8fjU7NWrNBNPVMDWXQ/CUa4bCT742cONMhKZh0pbLGIqFXKD9fmgQ4E5
I6aO95XuZUHwjpXqpzYJouvNY6ujbDxoH3UVDca3ufa0U1dLc2OHVVvTZlE9AQUM
SGCMPvrzQ6B9J0pheXYi6UD4eZSU4zz54oRlCS87J5rSg5qtS67AdaLaQgzAEe58
Qq1uoiv7gcbTaR+U8+CxxchVD8NabXH0ynbFf1tAT3vhAGiAO9PYfa5SIHCpyCsK
Zlh5Wtr+CPgo46sx0xi78pwY0oPwCLBgRprRjd9KBiUcq8lVxPnJmobVeb5Yahzw
ztiAhCWCw03bMyIkFxAR6kDH6lDWf0yGh2IzAIrN1BSPygiE05csr13ypP6jEHxB
B3NmRyVEQGVquW/WYtFERhQK82mPRLXR/xB5DAQps7C7BGXyZnCxdA/0SZe3yJ55
h/MAFuoZCflEaZ/PLeevnisxKOO8lv66stQoaGlmeHfB6TlWo7ZsSQ/V6EfJm9Nx
xMbyM1BOSe/czUR182jpr2SKSpLboIZnQOR5DaLKamhM+6dhKREaLl55Hh6VLWlc
qlhJnG+oHuz2uOxyYQQiHQTQY8pNAjjPQpYEhhDpltUEpZEPTFUACfB4zQCsWMwI
/c2ypOZ9HiK7PsZr9kHJuieNGyht23C6BhJMGJgs1qFNqW4qhXo1rvgk8vidL9Q4
e6l66eTpWTId6UqJhsGsVCe8CMdNEyqrXCGKV9uT3FMHX1ozNapUQymzUJFWYPgh
/GRZaJ0eFpV1eFASSBaxrO+MFqVu8FCJ4reeC3jJcLhb6wkcrFxWSKojFNE7gvZ4
ApLLPt+RlyNzewipmYro7rJbwlBvc7Tpzwt5O1UYN7FR+XXrufEnWG/4NunNZ5yF
xuHZhddbBVq0DuazZNL1QperCEvw9MLk8pybDY+pMdob5Q1T8+InP7pIYFDsC0WV
AyjmSK5fLyoYNQOvK/Qn2Lz9PRYGJYgLsfvot/PqQlHoQgg6vnlFSsi1BOzo5wkN
nFLLJi5grnxu1D9C0YrkPK1THpta8ZEv8VuQk37b3HnKcKqaAbDf2E6ygKkKJA8Q
daJkbxkiGFI9DtdIJc+JwBaOW42X8blhfQh6colAWEt7M78/nlZSO6M6t3uWVleX
nRlNscTg+yHJwATxvslKD7VmL6yG7+j8/ehKwogmhNKbwkqvBOalaYIMAtcFRCAZ
XtM0SXRMBoR+oaDM1yyQD5vIY0aNLOx+5yCqNomyLiq/y39WfpFEKUHwA4aL1OBZ
fOJPL4Eu6xkIktr1H00hdIV3GOjOy+Ut4+W0QS3iSe8q7/Do02E+go8N39fF/e72
G9iDi+Fsf821w2e6jUCUhXk/SqfCwknq36r+mNL+2Rcjlbg5qXjmAEA3n6Vm1QHz
XXyz+Ev2BY6t63Bh4js9q7GNuatWH23hVKn2nH4x7l5EK43PauvGXlQfIAbIzp0L
qQrJQDeipd0pBDwGGIeM6N6UCMXOYqAyxaaKnlqHvyZv7l3oUL6tz9R4oeim+xbN
tqZCj/G1LKusQgHMvfRbqVJBXyduCAsNnpsJkSzmzdJge/6E9WDSkhp/SXfk2PxF
JqIs8NF7swhPPDulSI8eXM1XXxnqX8RQfVMoy5Y9sNfbs/jZLgnv7OyoFBn2ynbO
SP/ErBfuAVNfho1l7mEJu1vygLr1KitgMnK6W/my4a0+HsQBpvmZeyvdGxl1ytiM
WWNhe49n/ztbagQGqRRP4Uu3R/QRHPZoFKQqJ/ClPa26e/DhuDqvzuNNNvlnhnv6
sOjU6lqS7VyDwPeaG+3+/qqI3Xbt0c6GqKnZw79An5DxsVbZBO8ZR1xTEtY8YDvA
GmOVhqOR0JerPhOwzmnqsncdox0I4lCO4JpSW6atZNu/Auj2hFf8aX68xoag2Brl
jWDyDOyctPNiGjfJr3SpsFiwAdsJjuffyc8Kef6OhSUV+Z2QrJT8exHs/30TuItV
med1H6kmwvlrUi7Bf6s2bBUrSXg8hTlrbI4XbxijV/mgGjUoSadyO4OumALMOiA6
lLv2Hno1WCjDAeBjCHAzC8oNBxHWEwXJDgUqhX8EknI9AU5rIiiIXimSUXr7pL+c
UYpZQxs3041LAdqWTLgnrc32FnZvputcCRn5XgQuETa5KQVX6fBeDBSURGox1XMz
hTq7ynPiZpT65T53Jk4KHvNKztHQ2t8ZWEpK4NKRHq0nQZp+JehVUsrzFSg7MiXC
4I/RU7YwonuTQPJzduVmjTmAajbApXnOgyeEb6jZR6feLnsuCug/oDcvjXAWUPYk
w9JCy8ZmKiKJ+cTYruXFzx3BdUW6PPGZPbQ8MDmgF0CtG59sYF9MKFXWkfu6f8EH
eA/9fv8jGrVU5eIjG6clX3sQKFF9Ol0aeHnFfLWNwi76UBx3/DWjseGl+VZgJe9F
RGzxZqCNKEXF1w2BBZxa3P5O4hiqIQw+C8VFObSGOt1hj6SQLkgcfksHFNVpKGhd
6IY/9Gj6TVcQtaMQx+DPG9HhDoWj5QpDT93CRR2sHKgECBJH1WE22g0/o/VdX2cG
2cCdKKrxf/8M3uwDF8348YRW7dwIqzqSU3k40hk0ethS0qorAZUT4VRFZzGt/PIa
D1SMIAYUgN8LUkjTuWIoFUJiof0RfyzbJM17wZkkOsVnpT2uuI/8JO0USDfQ9/Oa
A7ombDHgHypb5mlb3auvn7ii/PYsOc/c/2aSEFTCqcNM4Uv3UAryAzkrpS1MsVX+
6jEx13evhFJJ2MWCe8vA2gk4zojzzbvoGG65A8hMHETAuKPTtWwbxvQWdLUVOBZq
FW9Grt/RquDKY915gimWgHotvMlTIWkpUCtAM9Sh51O4g+Imq/kybIlEw3lBQBg4
QwxxlDk29JI23xX0Nv4TpijS+cr7ePzqcH59Y5f/ITRPz2f7TXiRrD9apriAOFs5
dsFWqBjm0O5ansgaA2qWHAbBNKn2oDQ0oqXKZMZldmHLfAlQozWH8GWGPPVUW4KX
UFslT9vXip0H2oOD7jfOA28oF90/2jVqOTcSXzSoJ6GYloI0C9XpljSaDrrXqL+X
D1yJASU4ZHbfMYlXTx237aFjavki6jpwFSctCZCCmJNBHnbeVi62HXndaqy5eURl
abUBo+LhdZJTzBpWUhQiklI3MJIvwGq8H87XvzOgmQtaMa/TgERiji4K63Xud7+F
n9kF4UFAoxtKKWbNUXI0Qzo2F1rQkILVUwktDC8rnWwlZBgOKEZ1/pUKac1iPxnM
M/jtn1zgfkG9npZBEAePFf/h23K+6SRf3ITV3UpXqhyYmAMpoJmuBFNEb14uG3fO
3DhwmIFlVp8Ud9IO44O/cCRpiYCBoJSLARgMHMJqiW17hD5eQfjBXrMEXl0oOfdh
o98bAHW5/Ojs3xVk2vos4gl54UvPvzlwLuWfVwnKf9Cmk68Au6lWQtdIeJVlDfVV
gZ6/A0B6eoMdB21qeNS7kqr7l0uzD0zqzJPKD11G+WeJ5ZDRUg46LYS13qJYuCQJ
8U1zzFBlF3ug9MEEM590WatPpB2aPHEkDv2sZ9Fa/GC51Ztp05kF5eOhlM/VnaKh
NLTBOYT6zzMyYHg8LVi+j7Jy9BdtALFhArnd5lV3BgITC3WFMmZuDqt5XnmmLj/r
gQP9AG3urYKqVX/3z9iPc/0wJDLGa+AhnW1rpclQZG8JJplknNvKaySMUI1+OFNd
zeyIo4nXZicgCkNACqZQccYQ2uSS9NTysdhhfcwv1lxAm1GQlh839AfU07GDYJWW
8OmS1twKD+ozHQ+BuWVEVlT7+HgzZ/kpZlxmmdhMXVvLZBexJ4cB4r9Ar3woQ/US
2HE/EOjgsjfzRsaNgPDZqILIJ+a2cvF8uAmAhKQaMaVseEgN7Wg+RnB++CHQVv9y
Mm7AkidBy4+CqZbdAqsXhWME8fAnzznAgtzi7hJVCTO6dzajutlivYvg0OYUd1A7
q31tpPrbr3fLGJUKIIRrtO8Mojxv/GFazEuT2VN+AvIRv2sEghVvnT379QeNZv+6
ORs4xxUMf3WwgsO5+BEliBq6jQZyR0j6klHpoYKpa/A36TBWfrcKjYMoHhTCESyf
FunmXR5UuhxYalGajUh2Lywv3uMeAHPQ/TKsGI0BFYDKBcPL+h87EflaoaRDE1ga
xRh6P+kLk7yFqiLcizSvqgxTTC8ZTMtU50/F2rMPl7fiAKsWx2yVE6Gzo8JzJXsM
nQAIXWd5K80JKF7SiPPFffQPM8RmIKgzS6GyUV8GnmQ45Ydq/tjRj9rsJy7d23gj
RyUP3nEM37d7Zau7xaolSXdZ4i4Hdm4N/niduUs0x067PVatghtF0Q549QfHCKWs
LpPFBBlXHz+7sUsQs4qA03a++tOFWjoYo6Ko1jsX4BiA4tOnLDPL2yKvV9MMLdcM
c3/BYbkPCz8SvxrKjHWXn+ldWtN2Z14I8XmlRs16wJMlKt0HtleyH0EHvPFz4Hdn
CAI4zdqJV48na/ZFq75eyJb0sccTXh8m7RdUZ98MOEdQQj5uVBZ2ruHhr6hl21yq
ToXNuvhrhWSmQaPQQ+zdK1MoPYliO9Ab/APGnlLzhMsf7/Y3jI4dV+1KvuCGGUTv
NOVGyuOo92cIqEBF9hJokjMUUr3nVw+E/EvRJBQ4OgV31Z1RSkylp0b1MSFgzvYw
bYTVAeYJash1J9j8iIfzFLFKg0gF5wPU822QZeZrpsSSaQB6mzXXvtvmo27I4duN
lbZxj/VfvCXNS21OukLaI5/hmmTx4HiXpn6wuXxHv85XsNI4UM9XmyyAcZysB06H
6WujgZX/5vq21XsFSO4yfBkZ/beL3QO24C+BiTdKROV1ilHxn8hyvmknWoZH0gDl
ewxd0cVSwN+TXzKCMidzhIwk8p01nTLPGPbrYj3dfBMIB7oZpu6T8Ho46EsUzvN3
6M7WBb5GH6O1Q60Uwbb2zSJ151HNdowRyWdVYWbCesYccmLepBgDUdz6V5lf6LLq
/4z5pDmnhjpwdJYi14q3m/bdu83fZatZG+gt5Oyl+mWviBAQ4KAQB9u2cNK4b1Sx
x81wMAFVDHeMYpQDpIVGT3/xoCyT1mPTVeED+gfIMPqL5EOmtCoOunYp6RYZ+X2o
3/GpWef1p9vk2Re5rDfoXNAigpEd0F9FaaDc85uaeqJV1rPFEdB43KaxYaCvUWkG
9xv/UA4QDa4UU2ggE6EZ13D0OEVWlg9OQRPwq4gd/Cq9JYL8e5GXdHIyRyjpkawn
ydZqH+OTZe3XdXErGT9swkdJAhTePcWPuko7aYHL5nX0OHV1RZPGrigAztuF2/Tb
uEly+leTNURvp5uSNNTLjQwMeyiiSbCOhKxioIsIT0PYsqvJwZIQmuURKa6dpC4h
8Lvt0bQP2u+CUMJLUXv/aU1mW8KDtCDqtrPeSl0GsmTrXA1WEJAXNOmmN1fITbjP
y437KUCkzsge8l+XWR6YfAqqrfIJz43IIUKF3nk0Zj7115VuzGKczDtUGIHhmlnj
G0iugHFVwh+xZwmi3jXghebDTxMeljItOTc7XhZLhAwrJsWZ4+SKAAAxuPfvDihS
E2lD9Ur0zwDt9TidQTmvZRRXo7V6CtBqdGICJvn1hrDWdbSfEc1u1+b2BY9mBWEc
ha/ycTwuqMq9EneaD1pNX2O9bC4ezA4Y/aBKZ2CitT+ZhP6umHsYu9FoIwSRCD5s
Cs64Xi6g2Qu0l5RFNuj8inJLsN4wGNf5NEWEcE1tHHH1Tv6TSEkjS9DTcYiAwZle
7zjTuSnGDb3tvFWBpJLjMoVr6emFPVH/Ws+NDh6A0yIobqg37n1Xdjrfcj7siVy8
DkG1X3eINwAoNnInUB9RtG83QomBVcvTWRmV0qT98OCHiu/S0HiI3F/CUb92myKp
k3/XgljBvW/Qbb7VAwLWOQ/BOatdAg18Grv7gsMonhWLjRbbk7+Im1vue9cYObPY
ZIELt4aNAAqEMRxwsp9iyq1o0kTfXmqA+d+94ytM3LPcZ1Gy+2OSjW+I/Qbghu7G
p6s+taHl1fPndM0dxSuSeTQQDpwZLTEFYTeDm87WusFmx6JeKjPQl5rXWWDxa6Zb
VjuiwDAmUYFSzOUBo0t10RfDLQWc2cxtYGCxifg0C0QZc+txGGs3ZgkDGiRDN/sX
oQ6AwL1gPzJgvYhb0u5RFavT4jMzhEmDfTMKl5y/Nb15rMHQowXGOCJlvKMbqudP
c3KMrNrwiW5DrRSY6XfrDjhAdnddHAVyt2QtOJLPVG10zD4ybGXYygD433irV+6C
c9p9IV5y2wo2RJidgdzKUd4EidOlN3iIha/G6UJrARlEJxlfVjWdtHCtCETFslmg
la12gTo/Qp55oreC9whBje+KadIm1L/5uhEbwPioVVgRs/9QNH1Rhd3Nov3PQuv/
ApWxJHZ0bkOAPk2Ds8ufPTkN6w366gjGMwA9RL9KkU5roFsaY7Tt4UkM+8oUuMrZ
nJqPRVRYzXiEBTF7xqoI3MaRvYvKA01eP3B/HeWwt+dthhSFVyeBGVGMMmQvsoY8
T8hPdiH7BJ4galGte2D5ko6Qs12gUIJOM01+ef4n6fxVYqyJz+xOeYrtsYtINFLy
2uNS/eLJow5xb43CvkhBI0B1cwm/sa/tA0axXLKi4RrPg8/HPvQIp7PCDR1VJEiR
FPERMOW7yvNx/wuutcLorh1o1KIpQaF6yrKOMbduQp5dUiQ/VEt0Z3S16KNq+huv
x378EMV3PeumIzoNDkuYGxgfa6T3RIeCAMdtA16l1qDkKVWsJqnY+iqbh1S1NFRH
+YEUO+XUzyOrZqWSv1Tme/nHooigt9YruepUiHUtj7E785OspNK4Sgag1guX01Ab
wXh1Ac5eT3z+pyzFKqln2lcvOmebALijWzQTuyphxazhSHIN4m8sWal2a3Zk9sdd
J+X9Y0pyBRAW1q/6TgdDH/yl0UU5MTkwXpaW1s15nEho4eFJlMTLOexqW+G5l5RP
u6Nrn/apbbe6eSUrIWxKcXBsCxO16dn+wQkQYvjrfy+eQCeTestT+PZixEQYDQIX
tcDO9S29UiW3YZd162sb8iUeVvmh8BqblLquVLXS59EB44H4LEPmoIGwN7dfsYNL
TMM3XPy3Qn4aBVGRn3dY68nwLj/202YZgwwAtyb//8Qejf6sftofKZLn7R4avlBn
owRkKtOQtH+rZwa+Swjt86YhB+K5HVV9pXQKcFqxNdERZT8Y3na5hvh06E37uejm
AxTNgidnBAq1Nl1fesSrUXTcWALxca8702w/HClZjtie1PYnMCNFsHTGjgrV1ik8
EW3mjUFo2NEL6at84oXlM3aornDwtTxAD1bIMfvxLARrLrdBo/bYrfLmoiHQGdcb
lhQpURImnmyrT/9uah3VP3IH6lfIE3smpH1vTmTznd9rK/4I3hZ1uHh2zjly+y+D
6g40l4yZhPdV2qQbK+tUWRwTr69EcK0CwA1eik7r7GDYNgow+0uCCaNFlVShVnL8
NSc7klmzvxdvkmD2Is8oyys4XEcmi8P0IKUYTGbAXSncZGoObvqazIjWd9DR2xfF
2opkpPwa/Z+XzXpEWjkDtuICVJxuUGhGCgyFrpMxLbJKGcXHieSG90QYounMFjnM
FHC3+lTzb83v3IF4QPsvBBtnl+IntUg57ueDHdQUToDCQLL3CRzBdmjN7w8wqmYr
E/ZkJUd3lYTzrm7YabCy7wDUNdHgI2phPQf+/f3zJPQz3URMGTRCELgqoFajEQi2
fWQrcsnS8itprxe6Q+gPOD2VmIO65DCVPSM6sxlhws+bbJFF2C3GaLhh1Hqpjtit
UlRbg7PZn8IOFWTOS3I8vWmLLBT5/9oiuFQWZMkDL1Es+oMsdKx4v3UYXn38K9lM
e2V9tBOkF7Ohoxu2Ym/73mJSApX3xsX8da/V5vvU6dIsSqEgxxavn/otC0tkPS/c
ePloAF7G9RX3O0rwMC47BN5+A8JaJTRC+UFIYor4RjIGUl6zpBPbt1UrErwNGPxU
2bn72ekiG/EDGvWBUSXkgUc8Wx8t0UeBomw3N+0Fg7FuWuF5/M45lnaxQxl8F8x+
s7vzBtzCe02czWldOzWmQyFBK28OCNq0RDVf3Pq+QOBnfd5QMnLJ6nz8gasHFbWk
gl4Ew0Z6yo/FI1qqAEk7aGOpswszYA5FvAONdxsPQ/VRQxMvRi2jIiOtC8bH6d9d
JCL7uzxzd3Ia9tZBE4wEqZoHuEwJb0PbcmQpewKMW8yHPByOcxM9bSz6ko7m+ZRY
0mRdaESMqNEFTv8ZQk6P2uQSybAxlHifz6HgnLvGUzopKr0jLrqqW6SzgNZGSLvE
Z6F4TXfCdB5tIkDurnJV3ANlDzQT28OCf79kSr/NmyWU2fCoAOBvDxWFCY7QyVVl
SGMBLh22l6TGy5V/fy9DtROY6fdSOlDQrU/R+zfXw6NJ7OjoS322ACHwoL1teril
QJ7W6Cl8cBUVUXbxKHRYn2fR0q9+MFdQ23KxAyI90tS/h9oO1Q50GKV1p+A6LcPy
+WTOSpjAAt+PJxbZTamzpSZik5PeaV9AMnp9L2Z4VSoSO5gGDQlDxV0USbPz5ktj
/1uQD7mhLC1q5D3ogGpPMr2OpGrVqnK3oKyZ8mpcO3d5RLx32wI1ByW7o9fwuy24
GXe0sOi4Nf6CSt+oVuYLOANLXxM6upgTY9RiTfKdiZ1xuBN0IVReJyMjOOER77vu
haYD7gQQPpy0r5zCmQfPilwsoA6viF9bfQjrDYS2W/v+ViSOXxjd07TRtSEi/E1b
ZYuApPPKL5a8HgqWRTIImhBRRMNwDo01JL2SarGAemP7kJN29itxgJQU0xuMgMxT
B5H5ywbLDQcUuyQjsuVk3XF1KnnjGavoxzPHWRHinc4KWCEKuhW19yi9AB0h5A6l
P0Dbf2HmD6ndiSx/kgLyqgoyxCGUXol93l5w8MGlIK2aaQTwl5kGEj7kjXsiARvh
GQGKVXd0y4uxAfash+cV+g6+5l4a/Css5/P2SD1sCwdwabLBTrd6PQWLp1S5FM3p
pPH6tqJvN7cckwMRLqqzMf6xQwv9/+FizycJMrzsce51lCfiu8CD4XZ3oqydoru3
jYY9JPivU8dhroEHhkdrdtj3BYbTgimZGVB0HPiLnKinbUsV08pyqb0wFj/GYt5I
pomIJ4+/G+Exixk/14ksudZK6m+KnhVU3Q5BJk2M+G4qAH4EKsjvXj+iAEoVNwL7
4UtXSsIVwhflgLDgoIrSxswqCc8wxRbOIShLNnot0uZ5611QGbOib9trQQVmfRFo
tmMYGgtuX6bxkDLXDb2aDIeJR6ziMFV8Y/O7SNnCNsxzvltjab24o4zYF1XW3yKm
OAuGOV35q518LBmw9ckaYmYP/SfdQXvxDV4UlRl9Ar/8eh0LaL1bzDKH9LhChCAQ
ae/4xZ4viT+TWuoz4NBPvcILudfQHvCJjRtEMqXbuX9qHe4oXlSOMP3RCvRff3Kc
wcOHvJMfrhByHtpbQyKsLLcvgrXTxq2UWqHk9dK2OVjfccFz2or1di3LmkggCjm6
dDKAzxvpHF74xtWNNgL8WH9MoNEADsbvpULmn3P2/ibph9P5CKxsqf+Lz9J5lCW3
SLssfJnURaOYShOVTyzgkxPxnWd88zepfmboZquCJUhiHR5A86AMdG0Yl1Wsp4pG
c+PZIP9U+qGpLRDB7h7ilEDZyji8cL/1TRn++pU4Ly66pMwyjHv6l0sbxoMLsRTW
eNWQO5qa7hVdNAt+tn7TkjQmqow5Db/KtdgN/i0zS/MNjqc49x5PtxFkXEFnD2d/
6uVmSzGRRlwGypve9CawKtISzBei5jT+Advy5IVXm0QBVn4QI5wvuNuSeo4GNYeV
fFLH1R5djvz04swlxWiZ3f4p5J+a81/UdBRDCrBYfAGbJcl6v2WEPSTh6uj7CfOV
nrWXFEZsPrM/icLlBgA7q+VX/Yz008hNFfbMNfW7rHUUPhpRLvEWTEjRhUzejt8X
h0fum/4Ul3q0fL9WTsbDH1MA6fdwoi/+jjqLGjgZZlOTm8s5P4JUvAxxbwVhmFqG
5PByH3yT0DNzS3yc8TK4hn1VtU4mK80atAqXb1h8a/heHgxzfMUnXaRH7D5/Q5+E
kU4ymB+gOoPJL7Dmhy+hPj8agw8wFHBQeK19bx5rF46r3h4fN75W2JNy8U90CgEp
1K3ipeinidKqc5kJPCbVBQ0LmFMLhT2VcqbRR7gYMRsi2t8xJROumm7e/6sWMDz1
ZeVLWRmVbK0vVqJTs7t5VQEWkIDRCRaH76T3GggAfAQMnzNDtZ10EcQtSdxA5uoX
9QU0teSeSkAvqPHYixpDSMbgOvbWtYkq+isS0RB7s3JsilwiZRKbjUpMQO2p3ZkW
s84Whqu6X4PMqbeqDZFDiZe79nqpX4j3NV3Ki+Zh+A0ioMh9t2BpIhc+HjtP0gTZ
/1xpaKYZqnqBOyFudeT1yK0RqEWKDq68bF7QomEBNLOZOiUG9UHN6ZQY8w91CccA
ejb7thqbldGtiL+UZKsCUrOmFZd0PQ3+IxmsIjeI/vRkEawOaP9pHH3h3mO17vjf
OnjVc+IRpHwu/PAWZSt88wE2Li8YpKYhbt3uWDiRHpzAxmFXgg3DeNFGa/cP7Iiv
EbgeKVkFvNkujVJ7tckpn/0ZGmebCsIsMnkrR5jZYj8J2bvx132+zSlekHyCpVQh
nS1vbHTSCVddsZYBEg8a0uO1wmJmQ8Np72qONxHSK3evImCADSXOn4WHZjtPT742
ZFVFXo+q9+GxmRHV4ERuNgd81r4WLrvDkj/WQtSDGDRRMhhNnot1ptQjub5vRyX6
ABTtEcBLLmWB3cibjghbTPK2LHGTcA4Uwq7wP94KSfC7Pr9gCJ+W660aFH6+WvB8
SB7gbJg5d6Q6Eta1MiKv/y+Hus2edKqXA54OHd7tBi3o4hyMpq2urZCiDGiHZB9e
tjlRas5l5N8kaOiUp0i5w1aCUCt6setup39+UkdTfbaX+wPy7Mkj9hHKBUhLQJwS
bBLGnSAzDWEqoNGFApo8hXClHCpnOUZibTlT7nlN/pXsCW7O1ZCwiBBbmB5q/iua
8ThHMZ5jGh4wujj7BgNCcUODJlQ7STaQT2GRS8yU7amoSMYRVkauoovnXctNxxUh
R+il+wPJ5rW1g0tzdeLru2sGcmGzBl9tHBzY7bttuDGZAk0VbCphQWPcXb6e9VYF
KOSPSB3OYSmNZ7GqjU/jGLNKzQC5bjugT8VILcm1oDS8tR46Yv9eybUdN81T9Si/
5L4EPLBM17KGT0/Qxpi2bzq1zTvaUACCX5ly9HmKgHD/hWcID25Q4Fcf+uM8mhYT
fXIdVBSTlXZvICsKmN6+0P016j+NgVN//Cg5d3niu2UHN0ineQSPh1oPD2qcHCoS
Ymgo4ybwhQ/TGZWh8tbEpLU8iudaySM715la8wxaHty0SW8mOi9QstvzPnNkjK/7
5WPSgXzyebmRyEKupKsN9vy6h45KQARXLLPpnRH0v/yeWgMLuExDTQoBzhp+l6u6
t+2tF+2UvFFcQAxDT8bdwZjfWBQFyaTdUc3nEMpfkxPP9xh76o6JKZ4CSgyUEUDY
n4Jxp4GnlEXKznKal6woXq0NxkfOIlo9nhJQVzHNYhw0BcWLO/5km7EFJ0YLRz/e
FEAC46If8/LgynbXkSCeQIx9UXfHWVw1hGXMKj6jDBN8I69nk7HVMsha8MvH88vH
kC4uhMDTYnzgdDwAq2Dx8PueK0VPZyeEfGXCQ0g3HC48kgQbZEs6vcToT7GMZVs2
qRS37mIuLLKOvU0Y9zkeoVHI3K58ggkXk3tLKO9Z7GdeCSRndQSz66lwde6d9jRD
vNQV784qMCiSh+LFQnUxFmaSw2p/VHiIDjW9/MQjw69QtdH49XxnbKtikP/lD34/
KVbOzi7m0QMJHU1XDcpqtaUOO12qp2G0EgDiFs7D6c4UoCggxmjP+zrf+vLaQTwi
aIscD4O4jfk3AU3yC99vI10Qlj1i3YXk6LxCQtFN7HpvoNiZ4jA9J/sljNDk0mJm
Lr7xo+XuwWKIuhtXefxkaJkEt6b30YINClL5Ypg55Votbp3BOAuI9sZDWUWFZNN5
aamDSo3GyQ4s4Clj3xA1dMBkbmyhjHvanl2miRNJnQTt9HoYnaOrJ/bEo4495Z+V
5QMHEWZrvy3JI12HcHFKb4ryTb9h90s7QhDdf0ABYDuU3wJzqt4kSd6MWNFMRXyE
D8/DLzGt2Ct5D5SLx+U52bd7R8pHtIDgqqA2QxVtJKZDltBc7YxxblNGH4eGjdcK
OV4rMPg8xPnTX3Sqquigu2oMzUi8S5KrWZoFK/SvcmGVLgIKxy2vJGOkGEJFm5Kk
jqck0BkWtwqemIYxpfbEELpmDJH6m9RV1NXxoeDyKqUF7bx5HR/SpHmljhXda4mU
L2JzxCOuqXw+rLPttA206gt97zP5rRc3dHhIVSL5gL6O2zOtYnZB1n9TpnUBLfS9
Q86X52YQFg9YDkUV4JbmhxE70dUchFK3bjECG9Rvd88dfeQcH9ab9+3oisiDsmRL
FimpzB1u03+mxa56bgd2N0xysRgYtv+7gShPq3E0nZhL+xAM4/fMb7IS6EW4ZO1e
rv68ymv98UUej3gytHqKlkQuYVN5gINrkntw3zyE4s6ZYyipA5z/562f2jENLFYQ
K1PHiVIoaJmbjPAkJdC7Bpt6MV4V58scxN0Yf2vvBY1Dta4cLnpj492EVA1VCys+
r1BmYoLbTFNB4Xkmvq4V4DdN/U9zM6W/EyktWzVaFto1XC4chypdqbTf2wTw1nkI
w9YF+PyvN5EPfLyRO6ceS8fWpcKSmUj6IzSM6cwBfbSxJmzC4YTkvFLelBPSwmY2
gvyewoEXYhkoZb7a8jvTpWS8ejEpMfN7YGBfko7De83IoQEbHZuTvgi0ih/gxZ9G
FNujfh6cPVd/bqQ+VrhV3jVNMwvl6I2+5nygUkNrkM/7WfdrGqWIDEvnXm/FFQSE
soGUZlKkTR3u8COTmfsleYVKe5vA3YC4PkfWKJmlu+qwByaHUXHohgMx/LzLbL6d
/1lpH1CB2juBbj1Skgaq2DZM7sIWHfBF5L+JBmogck/aHQ3VKs3x9ayhb+XAsyp0
Qn7ZzXj/lSMKvnVUpndHkSKZcHFuu3A7YavVqKw2YEYhVtvIRYwxhnGjQJh4RVRK
Cv19XFs0GqXKq3kDe+02ufxL6nynUS8UF2meraD/4kFMjE/kcgl7aBUhkgXS1g/K
UKHheYsIZd9ShwU+nY2qH3edLNh/rqIyTsboszCL0r2v7NeAVjlF/Spehf2tiw6K
LwFn1ceubVNNjeYKUNpF3iZeQGTS28x/5Ay2StTZdvyTZCXCzUDDnJmmZGgz4tUw
ntUx2LJiYWvfZtVajEid8ielGi+ykxyb0SFz/0IH1Ggr31HqceuUrtBdUXKIvO48
rOT6pZN65U6OguD3HZ1tTSTVHHTVKG2ZMtvpWpVh3aDMJM+RhtbQqTaIVepuoo1D
uXv+yawjenPUTuHn619BV+WGqRqv5L57fVHgHgfCLyy1nYqoGlpFUCJpzbS2Fpnx
USfOfZ7gbMGwjjJ5zuSyduw0RweQenFVNRSX/ibGgreG/FZcNvpYFDUX6qCIjf/T
N/oTTH3N1+r7vhlcU+0QlKZ/wEGzRUPTPjLowK8P0aQfs8GVgka6erCnUBEYzUwZ
2v3oDuc9eg0TT9BjVlQsWsYfjTP1JkKub7wZnszDdM1D/YqGf/VreArtG+TdkKps
rOB+RotW118BoAZwiu2rVuqfojghU5KFW9MJ6oeOmwZ4zVen/EI/EQs9JVx4SQk2
+YVgqSz7kij5kwNWLS4+KFiXMJzu81rREfl0Z80yBeaAF/TWmccAEB8ahAUyLhCx
LFEwW4XHSJlGAO8LiFbdQClr8bxD3WYZf7RhqUqo+J2plwLor3JzqrHtYjDgPCy1
zg2sC1AdnNDenz5OZgRaLvXYt/9bM7CIAmjfe0A58QC4IeOjMDeDYxMVkMKawFTO
onRDYJoBrqXa/zvtucWVGYBS+5jn8ghzkv/iWLs02fDDQynQaFk3/J5/PpOScd1T
QzK/5u8vJ0EF/aGmqq1gSULDyQbqrjs5Z4aeayF8KFbPbCdcGmvJRxK2y6KgzmqH
ytsNbN1GanL77iN1y7HPLEKgTfn7ptcx9p6EtnLsu1laM8FVKV5G/PLcfH0zFI2r
MWtD9xPeGwRGNGjED4u1Pisb05Rr3MSq5H6YFJj7vZnjqD9ye475/tY0vbW5/gHo
tWyK9Kg4/CDNGoKsfzdHUnE9b6M4Kdk6cKg0lVTWMy8aUARtuzUisQ+xRGjYorpf
uUTiHTJbYUlA7N27m2yKv73TDnG/CLvUxCUdFGzVo2fo9N/mjpN0P/YEcwqsanMK
4KEHl8CueLcHqqlnT7gdBclYKesOerqm1Lp7hu4fT2D0Gmkq1vGCxclKBK7aHs/+
qy4QApUh6OJLDkHkSPzorByDrnu4fQgoKirL+g4UPrTdr4zGXckGWhubQAGaf0uD
czPrifTezKAcit2wgiqN40xTsWj4Mh35b+X7h9EgCOeRdEFU/EbCDxh8Bug2jKcS
zoADzi5Evz7vYCKk8xyvm/RWm0hx6khOWsKtvIysYA374HuY8R8LvTqCVsEb4V2J
Vgb8vniGnu05libCoDMBPUqO7sR6FWk49xLqx0PjdoyblrXo9U5SXhCxHfoR1XTk
lN0MuzHZA/9N2qTqt0f7tkjuEfaQycqSabMjqs0aDAr71wlvTXMzcTJHhEm8H5oA
jpN6qz/fk8+r5u8aXGtAhhqtQbJ09RBef5F0M0ZXPlrI+dBTjiGW+93GvpcZsUqq
1jR9Zc1hVidUf6JOCvtX1ZihiZVtbrOnxFBMx9miO41Kfqm9LUrQnPuLN2FjMMc/
fvnxJEWeEKUB6+1cGRcA5SECHcE7jRspbbZpiiJA6gnlgWBTPr/FoSHi+QSGRntt
CcqQVRiufxXSTDDi0cBIO+PDoNDEG0do8ZkTQNYC04xg1ZeUCWztFbiyqHSA/dfk
iehohdQykkRzKP6bi2m/SuI6+QrXyND8Uo3SDTz3nSndMne0+Mw3j8KhcEHyJqlo
6XUlks+tY4JdTP2mnOIicSbV5JhtlYl/UcqM4rrAlvnBWoPxcDPHpIw8gPsqSE75
QqYT8x1eyG0DFF1gj7b+Ww8spYULk6BcVe0Edm/joMcZ9nunbofmHLAsdxJFS/dJ
UWvjRtKwhLJv4gyftPTmcupUEkiJgnPqBThbe3KXbFl0JgacVuJAK+EuSInqmV9A
kRcm2TNkeJx+GTegGdT35ZKaWVY4OP6y+TRvVrPgeHZulcgcIS9UpuNdF7yak5+o
dqqqDuZE2QvfSZWp89jB7bzqPQT9Nr57AINxYEAYrNV5guf0EuQ4aFP3vdLQnX8a
CtBjBoMiArteG7BT9AAbSlyHZgZEhLGoiVSWQhr6jgq8ZE4u769/TJeWAkzPFMVU
8Vucu5tmZMHIlWH4IVbXGSV8XCA+kHSIKt6oNsL+hs8I1i4ciCcc6/8qBTIAOgyA
RJc6M0RdSvIyhKcADsjoCsC1o9CldX6NH+Rx1jgs1zLFieUp+MZcY+F+0Fh8o0mX
I6hng/m61F/YGy+EIyL285raN3YYZKXA0hnEQrr58FYSJB1R1nSAaBF1nHhEAcpp
QSX6gw3Kuo1ndkTyZwyHxlzaZFKMOT5g0xgG+YfqBYqgcA1ce5ZJ3zbCdPKUzSfS
CML8QdyPN8KJpuI+crbKlPLQja/9FGepwDDHywDGe0LlR1mWWznmXHhp5LQJZL/6
dkgPXiUcKpm90zRWSWTwFXGrH6d0XWZGSLyJgfZCej2trStsqXWX01FTO/ThFzai
ksR//AeAfRT0yv5xRxXq/2GAaCAwZqyqT9gdn7VF6qomuc5SqiwXwnJf6pYq6/DP
+wIfrphu7ydAtlBmU7+aaSxOvT+YCoZQ9ooHwQCQ8mAj7MopI89+nq+0phobRefA
IROZhyiU73FUjENIqCxUYFD56IKAWNiPIK5MI7/WF3w+mnCl4C5ZfJ/5ClcnvD/L
rrJnwIq6fQIPme2ZK3Ed48CyeQQ3YNybc3sRHZ49Ju4oXjeZdo+os3/cXyRGQFCV
Y6C2WIiQctEf2j5ICJ/ZBjvlpbGrKuERpZB/ZBw0Od9wXsnkuj9sKlWcV+TtdS9z
+/GxPao9HY53oI2+KC/LnEF6bJm3Pk5/krhl1gpqNf7E7g6WnyBYLw5o1f+2rap/
y3aRMvUuRg0zNw2MEVya8Y8GaSbGJXl5v2rZQfPNUTkq+eScCip7ip733Wg6zlgE
gAqud0SeemS16SbTZOpnxFd3hUCtsHiyPDZ/9hbMoEBzyinyO34AxSYTjjeczMUx
bZsu+V1enR94+z2YapWAKOzjn5f3tNhTU2kWkU/2tyT91czRRvqYBBk1c0byRBB5
hfIq1TnyTWQNXIIfLpat436hoxqnLkHFiMMWS2+VloYngtHI5zgs78z8MXyqRjag
Rpbqv7zV+EQPu9w5bwrSLgc54k+c0Sc5WdBK6oOvqe0+bjws6ZSlXaIwVBTE9A7s
i75U+BNsEyAxa3v8Yu/qENxO4Dt9DyLbpnQmBe+voxWEwNWB1LTLi4/K+8Ajsntr
kdkyemZGQE/BGgH3kqz/hOt8THnqLddcjSn8FEk2ZtjiovylprgUQ94nwClpTONq
PC7yk9lakyIKUgibtBfKKXlCuFaANKzSotOhTRm2jZMOC1K6BL8jvIpWpELgHuC5
OVlEKVsSIJE+Gb8n0f5v5OhJ7u/Ae6KLvCqVmsUQXQBSaPYec8E1unr8kK79qZ4R
e1CUsK72+X4Blq8Ph+4AyRDh3252JwkZzZSkweNibxYrnieVtQOK7qWRxVP4DR3H
04gxwma2ts93VWmd9cQHhSg074UQ8fU5VaNLM/zr8QkVc/ylQmOM91aISkhdqyLr
tp3UuyxzGFV7Qbtys/pxToZ5GKNhx5+npxR6YVQcMMM85xM1guoZ14A+jdMA/199
LFg+1i+8+3zkRwAc2v4mACPJmPiuhJ68L2e7/84CfXfwHUgyMq9y+cBATXd0CRBO
SqRfl/4ehPc50dRQ/nocs1mwo68H0rpQayFXc4HbIpANgY4m5LI26WlUyVQ2Vun7
mVkpzTABsyi7wjPwWUJ6ZitJdlGIJmH8Jg8QbgU+H1ULSTBvzZLBScWqpWjM9kHm
jjd/2r/+Y1zj3Celh+c9WGhA60rnqyCADHnj1jKk7pTaSBKkntHqXdC/bWd+FoX6
fP8Mjp5ddDZ7R3KrfG5h7aXGIDCqCxN5lbFCIqOCxddPG+aC/WNyN9gjk/4d5JZ7
cBKE989TxjNkMF2KCMgyMKvBtKHY3hwMpBD5QkcURBxyy9VrvMZJX8L2JTaZfTSr
+aMatIPZwmt6tpfTt06nmbnvIt069hwfPqHH6flTqoEIHtWxpugPEGLudEYtqKeh
DO8+ZDtiZRLvdkAJemUb/y9d3q8Y7qiJ5fK0F4vCLsCQbXTI+LP3hLZCE7hGOAZ2
FEcwPzy1k6zTvUMLBRHqHEw+c69oZl9qtuG+XtXWEGNCUfZIQaYKmfk5YLHqzkAY
7OfVMtpgElfYLbBBQza7VzbtW7utlNUOZ8GrGqessmMtkkSOd3VTcL9q4WaUQa4G
OzAZ5UKUrksoz53UK2hwk4k7qVGWt+iRlxP/awtMAiOEXL77xuzcJ7IM5Cc8k9uf
MJ9Bdn5dEPh9/ckptZrU2Eiva1D2uf6url9CM3S1IbTvMWUZfu+KPg7Kha3zi5F2
zO5twxaRGbKuvMFxZEfjnvT0CBRfhvCl/Q77rO4Xm3w6duZ+D9v1gD/7JyAHwqxE
eOwxrZT5OO2lB0NpVhtncLa+vEJ8YQcvAytG5XSd0CzDX1NwJM39ZK0XxX1R6RLP
Gsg/Vtoe0xMEymDInqgkxA0CNtoDFRu/zjS8irE3V8u8ZzuD8xeIoO1oOngoHivv
Hex34U/Xj0+Bw+HN5vljtBiNZahYR8Jcvd4tpLe2NkPUxoSs66vb8qXi8M/t2+cH
x4HptIcVdY1zV0+gYOBo62mE1MZO6dinO3KV75mAkWEbsiA7ddv06eNIZg0VrKc8
i7aZIc3m0WsKQGDbZv0460M49uboseOeMIlHxk5UricCwB9s5K/wREiYW0E0M3Au
c9XzrsYwjorCUymPjUqVnZrolWLRiTSSfedF8QTr4Yvdevp2UzfwOgK8ZRL9K4Rz
sh2LCOvGPWi7L8qW7WVY1jYHkLqXaF1WNiEkQNIzTtra0PfUpOuC8m0lQ98nG5+E
8uFS8Ks/ac+u/4rvUHYsaM2pSKKSo6DwfqkuBPxgMt+ttngJXQKyvo5vM1mFTCQZ
QHSo4ZM2rgymUhtGGpn9tYumTcUtQQ++gjyrZcysYC/Zf4vj4Y6cjdQkbadNv1vd
zjinz61LPzZn5F8EQG9d9359wxXQ2rYxeQFP7Jdljh0kGKrE4E0Ja52eG9n0gKMm
cQf7jf7qrTdp9l7rOQPQ0TOOg+2HAVWAUAKK+DSp+gfFmKakeIfncdQ0tnsZSBtJ
lfNCJNnlDGIrMwZ0wP/90LunLwtXvn1bAOtsc5WQNxc4KHcDBJjHI6cRVFWG1/BD
sYuuELWPM0B50aXp+4sjTX+TF6svETPNujX38aMkpt7qOK7HJ4FwW9CLOhlTF32B
xDjVaenU9XWnANuHVrQ8vf++zSPLiaDZM1SbxKLXTy/520GlMdisGW1NSRG2S6X9
rFploiS1KodOBUSt4NjdCbyyTfVk6BX+FXopTMAWON2/EzfLnNKC0MGrrYIwjwvO
205yLnHlTVuZ5YsjaC40Lwrdv9NW+Cg+jVCgJjrff7FFhDQPEr8M0FiOCy00vbwL
VP+x+X6uy59NdE/17A+0aqYJwxuYqdddyBPc0+Yjph67TpZEgeTvGoT4rXhfjTBA
PSwZVIv5YEpUnamQuuLEuJ8GIZKFQcSIrzIkegva03CQdMQtb8N5WKOb5MzTN8Jn
elAozcAaEPUGtKRozogneE8QT3ID2v50tvLKDWjcIqZVjtvN+daB2OkyfEZx6UmG
NtWxa373xaQ/vTt+ZVME8FvsK6BUWnTafUy+yipqy3rygqN6vtzge4x06bIw3Zn/
ASk4kpM4nJxBxdOwJ/iWAkvBpzE9j0rPaIrJmEkWGMlYiQKgS39SGktiNyHDelmq
ymmOfcyEZIhlEAVbEeNlxlkJrEsTZYGLNzURwYGrm7LeKKLv4pNqvOYfpDhi7RLA
hFHI/eesbtCIubELPSnV7enqXl48b2tp3kVjX7rZUSiMBikUz56GF9QJx5vWGuqo
VvWoEMkZ2zlUJsNaoSSD141N5oXZzV4olbt+N6kBXE4Ct7Y/HoOB/l9aoDFLk1gj
g7G/vCz+kWrv1s6pixYGuBhy6Rb44Mje/aif+XlsUBoOl1OWL1OgIQL5SaZ+e+z7
bvu0dzM0Z01E3tDRALFk7o1SliRgM1sxYF7ealqdFpFTEEjhxKCy+4AZuXS7qw5u
hKPzNB3FNnOsOv1r7YtgaaGAErrOf83EVfiZkyjo2NKJHToSZKT9nQw4/OW2TCLl
KTyK1Lz7pOkn94us+k2nooTS/ybrcr3LkkMoqgE8tMEXfvf6aQix2mfnqLFqGPfd
U0EoMBMvjLaIqRs/TSHWbR1crlSAFbzwEFRvKidoTk3KDIpatLDviC1wtky110zq
Z5O60m9fi1RsTlRjcxxjCib3nIs5karCbPzP1NBn1RpycOLvVlFaqO8MzzniKSoQ
NNG0yx7uGlqTKnNGoly5+hbYfkABU9I//VPxNiQ/lFr/+xRjAag7FnNEG26SxIj/
E6qiI7+Ekj+wM6fQUHfJIk5Lzw3oc5Ij4a7C6FrAAUD6Yt5aMLFMI8S6viK2CM+Y
w2GqayI7M4l5rJOt9Ahe8ImmW+ug6QEsmqLsjPhBudOPpGpFhXeu7I3a6WAH41Qq
mEJBkUKdbtGj4tDqyluKDmqC1MYCiW1WZ/moDdj5lkCylVVBYiy997FoZttehper
+SPWqtFP9Ke0jcAUQebOmRap+ub59ia8YwCaw58hPR9Hr6i9h/bvhigkArmFubYg
nIPd+jkrmNDuCUm00UBhnUEfDfbHiLX+4GdkGNmorbgqHE3f79r2AMdW4M0GY+G5
omcVU4PbndRBoXgXRnJ1ztG1qdsvVFe9NrPjr1WTMXiaFc2ecqY3sao4a+igOUPo
X28XgFh37Ldo7r4eFyaYFvT4r1k/LfppoJxntc+Kl9gUdVlx5uysXazRFC1XqQKF
Seak6XA9gaddq62/UQHP719Q+F8nM1Ht1kOWHs9VUvsqgZELdydCLOqF6V5OrZ1j
mkCXZJjTOBE/4eOytZwD36uot5F/eird8Qzi91imqv7nmRlL+bfw6wPlOYCWwdkR
eMLissSMFFAeYcBzAmKXsJy2vOLnHFrRhpr+A9IRjaD0puDj6bovt4yxOMkSK3AQ
+o558hCsa1uOwW2k2qFcmzEmZYIoBKRnhotXsJQqVuhJ2PitoClKFtWaWAnQv0EK
81J17+2wSnq+b3CYczC+7lhf8tw8Gi1Y3zqkQOESwTKH6zVCIeI9lkLKV+BdvKKR
r87RpJw+pwiIv93FCtVA9l/vFTxc+WoQXH5FdymXlitU73azbSsWyEAx0NroS+u7
vv90NnLhCfwtrGVEdM71ZASyJ62XsqIPtU5Nl8jpFoeUPLtQtXWTpwRKZ/VC4FQB
wP/n3qx6xKO0Ph44/SZ/QiXnYfHcuABzgY948O0hqSOedqEPzhJE/M8yzeg3abmc
EblitZPBq50wt1x4Ia7Uq8/jCiDQ7+0uy+gL2UsvXXNi2lm5BoIRGV071NCdTQ7T
OkTsc81mppkbtUKY1E3EZnwSVAQ9KKAQc+mUK5t/WuCJIaN31XBEFNe0QhOrBgmC
H/8h4+6MafBN7iBhEB60xcFRjr/ah4sySRbxqbNeMAmJrJ+o8bYFzyCtBgCuPbpJ
+OAjU7eZQkNpRbYzOVEv+gz4EHBv3bdqBWopdBsCAFnq/30u15s5RnMeUajeBV9U
7wGsAYt45lfNJkL3wDxLFtpebdLVS7ebxJe2WJ/bj2I34dTtoPecZGrvIkBZtZPh
Op+M8AyUlYmvrvQ6+AD146Vhog0MBkqN5d0j9nRiWSSDMenmHvEXRcO9XyoxpacI
5uUIhsUv2slv7pgrAD5DxWQzyIIGXzvRaSYB/d2t3mNQtrhFxD7/YCzQ4rEwzec2
UDwuww8cchN8SOBg53kP12d+/pBuEM5Omz7tHEDgVqPbV/VjkiMWKuzclOu1tePs
FUD89JGOpUQjkNVbOVU/pqyBtNEjLIWxgOX+NSfQ05JGqmukr6mc7+tKcX/ZSrG4
VJfu/Xwy+ba+stqAhfrNJN/2b0W1noYg5rZDe/EkhutFmR7GWc2YA64YSHD129Zg
9lcIUoC1AjGOX9c4CrdxK/jiGpcTucqrC6+UGgFNNkjGkBoOEo5V/XPWJiKbPl8N
FzdIm6AmwlGeymEKmLwRYyRcJO7c0veA8KCAVTKXspZUC8w7k3Y5jccgcr5uJpVi
K/o8/y++1oOpxJxMu3VAQrh4QAa3dZyH5ESCauln0Uex7jkhVjnVTlbPNGUcrvzY
OTX7Nr05zt31GJbuVc2xS10IFqQL/nA4PgEkM0z1lafWxsVcXu3LX6BYIXcNCgaN
Ps8iI6y5KNgPUJvjNB8rziDvUR9YhPkWxwWhWZ6kLf/kiMo8xla0BP/F7ZMMW/l6
c+HGTvTPI17OEcRCN+0b/erb0nsnFuYrhtcsG6Z4fgPj6lvw+ooEvu0HAiHZT6kQ
CzXtoVat6DwfpUwlDSji99coKd7+8W8MqwTKeKFsPIRXrf60SPD6kUNWVWjo5bKz
r7/KhnSWMlgRgpjFlA/hPnO4I29Xq30qf3Yds1CrDVFXcUSWe1+TmGCn+tHkA4pz
9AQHdIOH0TCI1H57iTKbDYSHQhDJ8HQzw8kjzq+UDJw0CyVnONSqQCAa4ZvwRTZ1
osX4dorg0Fz9PiTKdTQusTpX/borgBqR8dZ0aA0F3wHU1H70NhUciHu2bc1PW/0m
TE+qs3cFyr2/83vkfFdFSZ1eEhnKgS12jErCM/FFW8+eIzFOloCqm4opAN7V4h2e
Kf66PaL+Pnxz5KpKVpDOtZ+1yn8eH+3ECNhow5Um7VniV/iFN3x2nViYVvcEN5Da
C8SAWNeBf54qxNpe3R4AZLNHAM441TCHiMUFO7XjVtqUJQeSG2lCyP67yE9n3rbv
wo5vZe877MeKbWkmjtur+eQHHPaSsCkpXdNXNmbHNs/0kfA1EV3X/T7enMGJKQfs
YX9XrrvGhgBh3eaCbl7mgdVMphJ6F4lAm8+h2u0b0586L9v0E5OuEcYt0sD+agIn
Sud9Dm1TF8U49LWQPiD4vQ07RQXf1g1oEwWKTVW5juzYlKVWHez8RQxMByvzDIDi
KKndvs/vbPqPq6HUWoUH7m+LO3yfUKevxWRsTIRUeI2g2zpDkWKuVDWsh2xuFZ35
RtikiCuXXRUNM/mNzuGHy1WqyiNP9BhQGugKLQCmoSJSw0wFYMEWoO/AtfBlvSTV
L/VYaK1smlvzX9qXXEUwl/RVwf9+eIVZ5ApQdUcQBKrATlLoIj6nWGjyYe6XaxTw
ylBtZ+Bp0JffYNNxdxe9vxhnHm4K7RsXBH2tOHwbmIN+Qry18vF2XKiRFRKsIjjg
8YiieHq/htfNY+89N1cSUvtMbp1kV/ahhJa0HLGQbtJWmu77TMPBDFvWECT42PVv
iYv3Sm5zTfWno3Qgph/lVIQOBe6jll6Irg3tqsQ4O3atxUb3MQAQc6Fv/GihsE+E
vwcDRPxoJZ7dIXMhXnb7TSkG5657Jc8y0Qik1PPMH3yk/RCLUdgslJ3bAZ8GZTEK
8TyLEl27RIxvE6dHaxdWXkSHr3jAqVDHNdks6Pg8/3YTiZ1ZhGREfMKZfIBfZnhc
4dYi9J2nMBS0Gix1coxIRjLIiq2mSn7bibQvdDZNb12uHJp4/j3LDEm0/twN0ahx
L3rwvrHhsKLmzf+t56R/AyWqSeXKEOAaGqJEwvlfoUIKbJq2/VdPJ7ul8dCVuAHK
8FSDGFZRCX+F3nXp3vV3hLahBanjBLeKHTg5vCnDxMlL8t3qvRGkv9yJnXvJURGP
doSiED5tqi3rdta1dt/YIXefKxj6wxABrr054c+m36XvQCKcRh3Rc25YByClwjg0
Ogk89RIfbW9bjw12PtC8YVxRRGPKWSLw3KRMeBiDg4L+rX1zOFfkJ0kumEvExOML
QgiyIyy7TuE1p1HbBtsXfXmoubVCO6ySWWcRyr+U84Zg3jbcgCvAT7amEL1ahbzZ
Dgr1tPriXygJMDAzruYLU9ZiEbi9bWvL6TO1KlQgYK045InuTDmC3RcSEcBvexr2
OlELbUfzKDA1Gi6dddbwpaOxJXeF6PxKf5pvoEenk3ifuXOKLLkGm0b+7IDPU5gI
pSb7L1P/cdMzO+2hxb8fzkmoXCaQ/O4lW9WV/zBab8r5JXO4AW8TnVV2+6lVAjTF
ox724NDsWZU1nTOheJmoCmIOyLHp6AxP6J/EFrRWDtUgTbdBdfcUucQHQFEcEYpY
Fz3GK6w4V3tozIa/nkdohXRL4HASssXgKWq23l7u3WSatYUhIUSeR0M4WRXCHk+4
5mah8cE0KiHaML3CEfuKPOiCKrg3rKLNd7rIu5E4WURkEt0+aOcDTxz9LIx6zhuS
6c6nWhtJ/YPWR6Tf5Z+p8l9cxrQdDentp3/9Y7Vvb9l02DjJlZrOlmEUgXpnILOs
XbLgT0dlS6skDxdfGUOut+6kPJln15eH86WrCvHf8bZguIBhVufjxjoHmdBXCzUz
Gej4rdke0Opxu0lx0ifNQy8bu/1vXLPpBb/4PrPZltZljkVrFl3vPvplS4uguWY2
j56nfTLFVoeLnDD4H9PygNnU9iVFcqXn8dduaTt0DMq+kCS/bUieoYY2/8kWNskv
rEvujFB4aFsq6clo2X5ovAKFJ/DORGNTMw2CZ+E2j4QD96tMBDeHlXAUp7jRFpuT
FqGKBguCqGXnJqIkc6503++BEOFJKFomJt91yWkUFcTli9opkNvMDF24MLhA5hCn
EGK/qa8cfz+2gByQJpREbQuvysj8QJ62ug+L7eBIdwRzkuMIck7YqvJCP54M4Usq
1ym/R5vVjLPhHMGWAMNxE84i43OlT7gqcEK1us1LsTfBPWjVsMOVbGpaMC9+7BDX
5yfxzoFzQhbL9hFHa1iQUStcIrEj2E1hBOHxu59cIgtKmTxPN7xFISuGHhtm1POC
ciBjSbMiqEtM5BqLtoGFndPPubYQKd1vHQj4rGkLX1fTL/Jm3Pk8TlG5CXIy5b5C
FzI1cOtXjzb9UI3KhUC+vmPvIrxlz9YXJrWvPv3VbLbI0brL2nm9fIqzdj0VT8Fy
Ph/dXW57EzNvkQZ4OawPeOvpme1b2xZ3H8lYl/lLItpbydLpztwZWzMnxUBU0SWQ
hTRvh3g9dzRhkAD63HJ0t3QLI7sLyvl2HjJJOgmwA2qg0LkK7JMzqgnhj0S6AWJc
LHVLYBqggNt9MkSOxPFoEY6x/qi2uOXxVuZFfcGKBtSKZ+89aBwKYWvffdsSO9r/
n5+SKjlTeA2dndcpTZTTQZRrf+j3+kQuhwve0qL0EqbbeTzlNfsaIS8FGZoZGkZx
IWJJ9epv1L9kY62MSi5roBWOZLx8qNgKaKqGBEscE2NlO2PuvYRGNJsK3HbPrmPL
Yhdxr5HebQWp3JTAchxZBzyy087EKQLebj9z3drVn8qfOuny40/6Bu8f2M/EyqJr
suxWdlq0LwZI5tdlNqVZiIH22tzb1VuyOID8LQhf+1gfNLB8qgSstv0suF6/SBFR
2mt6kEvhCvpeW0BxDik4rT1T6MR7GM1kkrafs+q7pOoe4VeKlF9Nng1APhe/zU3a
DBiW2jpZO7tls/iAnojWZB+AA/B1oRH4C8ZEvu7l16uG3jkbFQYskNqjkOMrZUDr
cnw43zsAFGGcyCpUO6xuHNNsrnr7Xa6Relng7wQhqYfln4PzOHnBqBRLB469VWus
au552V292LtEMk5h5riY2Qv0nYy6Rz57yn+zd3IZMw2I4r6G8KHyeYRZ5AZMFhHe
kDakaIkjxHb0cwNCIu09dAhEECURVVwOlmxzIzdhvQk8WusXH6TNP3ElPD3tJb/S
RmWEAq3w9+bIEvXwaOwTBxnTGFyYwqmtRHyabxvTvMaaE6XLns2o335oYuIEkc0R
2IquTeUMF44EHmPV29Ww8g8bQhnlyo758XiJfJ6dWDe4Db/+F7EIolH0kH6vup7n
+VDBS3Pom2KTl9CaUkYRb7TkZ5r11LUbnM9KOBe/628dTZYDxXpLmwDGeDupXpph
tSpYuxM1BbZjjxe5du7BkRa2ftXuhNy4lZygdlrQdgsYUcNAgfM4qpwyQ2K3b/I6
gUnlz/P66Y7/NjrIQoWC97mFhMxL0sy8KZbVEdr9nuf+zSAI/3UJNJgYdmyTZia+
i07A7ScUU8bZRoM1GC5f3edxsWtvgz9tPJnKEQ/zSYX7qEEMB3RTpc4Q3Q/AGzmq
nAipGHKUUCwfyyWw5dfpRGKtaLU5Fd1Sf08t0rYzGlsZdPk0p0bnRteR0ypj5bO6
bADCv6qJT3+BW36W3MpEMEEvy5gElCO+URaUzLQzFkQ6VgaPtKzE9KM0T2C5iweQ
StcbU+7chNrZX+ci+AgGKQtpbnaj24WP6XuLBYNDxksMR9NfHfKS4quclVi0nGiS
aM9ZsCgnY4EUnmxYrMU8Fxb54UWzHCQovYLxzlOx7inhf+VIwkcq6oj/Lt+4AQ+b
oJZKu+tVLHDKx6iBOihjtAUX54lxR63h7Df0/cEOzDY/DcNgxOJM2mMB/K/yqM69
r5rOjk8SpzmI+Ma+r0yrQVUHy8LKxSdqcrEVxMMMLzY+JRDwxR2AtMpE6rlAaOJc
AV0CRV2wy+FhJ8pvQc5NVVaibWnflLUXoRz+J2cLMRjMiOZ175UTmo/F6O1pfRxl
9cRL4d05fUYBAYEec+Js/uy4wasmjX8uPugSQHY6AORk3Gh0lvPS+ke3h3FmvMLM
UvEEoBhppPlbsBcAv2MgQo/abtb4A7jYTl0LBawCPrxmSgDnh0+G+D4SnfKvjvPw
Y7lhV7pjxtVIyNx4frpjm1CIN+k3Is+zFt/PkHX74slpRQvjuE54XIfQS+vvybvh
g2cWu8pai2EVLSlybV0NmqKFzEf63juCWH93cEktfgzvXvgvLTxJeRknaBBAdZJL
RdDxMEmPEDK+NmjZulzI5FRezeKPVcicgMA8zquf4pr3bVKaGw91eGMr+XWnxiPk
TaI9L0jPx21EAeKqDrnFhNi/cJAhaRjavi948dmlT5jzxRNcahol8SxhxIgK2rht
3jUSv/bNv9+h39imbGEQEQuAuQfHxRRJWO9W27iAeQU5NYCs8GY/+wmoAk0ugIa2
JPC8WD6YVns745vPYfVTEpkD4B3OyA623Pp8j0q5Svkjh6aVMzsM+oeyW06MNwtZ
zb8f0nXYl2Ep2OeXae1n1D30wb5xqN8oC+ohCkwp8nETJHZlGYMotwAQQJ4v194S
u10sS5z/SEQ//VqPFSrdzNArWKQcTxfn4f2hQfaOa8S03qVtrgledz67bK9s6Wec
PGlMxRkL9aUNNrd6L8Zv3yPbJBW+ZVwNhyGiaNpOd70qpY/hY+In8mcw+ezMp97E
mmUxv/FRJb6a09TKIPucVB/OX6QBgkmpDoXuoHPWMMMDmRQDFn5jfmSqIMQwJV9N
XF2ktz3OkQEZzjkT1jw8wfoJgoqKUhy5WTvF6L/+rlJsFNgKZ5003ch5u5ByfaZB
zkwV+M8ACHNCd8AwSFT7enn/g4yU1bcMm52Fv/zRdr384iGMQNIOhpVJ+oHlZ6vu
fvFsd8NDpIDOF97zZ01LCn4UjTrPYdv7pGx8o4YA4krQdzCSkm1l7Ii7rkV9MjT6
1MJ3otPnznmTKu4YF3rsHkKnzdfhHKwlHyJyfBIR6T8gAG8TcLZlSw/IIfgqEBjq
j2FaEGK4/gEHIUBnfrQABoRbhhQxoO6xTJ232dGFJfSgn9LODoSM+SbOOrebL9ZX
HnWIei54LX1sEMOtKOi6mZkKInFTsHw7+idha6cDJmrRfj8u7Gg20IpsQtNK/Vt7
v7nZrXwtjYuTF9KLgIxmEOYitI86xYFPsLeehjCRKAUPZJjjvHI/9zisGXbAmCl/
cIOxumNgzBCa8xF8HIVeIxVVRGZMk9K/IFqmUj5wZT4d88sXVx4uh6Kpx2p5pK2Z
bVnL6WOPJCojOduIDEDtb1QiM9BMWMEFc6aanJlNp4pXvdqW/G0MVLqKAATMv9F/
AFt/1/w94uusHpBVFLVx/7HIavkC5lV38tLn5YORinMVGYpy4E6eMwreBCuXrNUt
YPvstRb5sQqYauvPGsUov6sy33+LV4CPPRqHJ+YrkiZ3JHrp+wbLm7bV+Jb1y4U4
BJlPYI2ROPf8IF8LzJmtq/4e4euQASNUQ+ZTtZw/UEBBrB2mbwSqYtT21cYkCPpQ
PgFww7R0BKkCjhikoUzbQ6t432d1T+GLCHCe6wcvomfM9ItISuBhYP5d0dGonPYp
pLdceXWEa2bhuUDBOlRJpDO8j+/V18hoiPDIp5x5O9m/qCyubIkkVViu/Vp5Iz3y
hhrCGhpE66IVhxM0rNjNXh9JuELUFWg3v7Ip2m9D6lnXo85KTksJBHa/7PT+F35L
97KmAfyVHz5QrsmJL+4aoGsU0N84l7jIrrKAA70RTgJT6QJByPzF3qUSDvpfTmEu
C/JiIcohU2IqQ8h2atk4h6Kpd5ynfF2kJq3fAlfUyZYOyXdT37ErHyVwGjHAp4Q8
/wcftMAoMJCR3zv35ZGk82+L1E16FnafBXxDEBz7hG7IWnotuORdPCserjgRt21A
7FdOvXCN4HLpEPid05GTZXQ1nU84lJ3upoIMTKUYt976wW2azepUNAZy0Lp15VoJ
Cm/wxwjNm9/puXEL02mFGm8XVGHF+OVhUG4YfFF3BCjL0wHY3bdeLx4/h+K7uXGy
ynQuOu5JdmGma5XmCAC16CcWrnsWc7zZzE1pFMXxnSpQTuixAVbKS+P3UfxqC3Wz
cKBklXWXPQYmusCf5qZRVp25wGMSQ6/tav1S0afFbakp5kaX3rdLyJM6T9yxhzoS
rzbKeSen6j+3S1A21O5uQGMQ82WL3qBntHl3qqQjlPNU/b3CUbgcj2SdtZJb18g3
oj8NWlKSi6pnetuXphd2sd+BRUpXTTEIQd2SYytb5/Gqv+i+hFB2Z1zJz3VCF67r
dg9Tj3KCNkFnIjPiMwxeb27jJUlVGcToACzCkBpNWu1JiPtZHE8ilvdiBSuIoWyi
MSytbv9bF6HiJJMMvX5Ppl48uJdtI9IhuIoIvgRvrvv6U+IMQzYKMOwLyS+/tr8u
aJepxuSPRXc9EhnY5nE4IgEY1iGumo50NFFo8NhtIH09VX/cIP99Qa3IB4elgkOJ
5vjlUrwV9UR5qhDm4QCI10y/fihUf3nW9VH3VIBIcHCkcGi4ydCDt5gduLRld1JS
VurvP7oXB9MU34DuKigS0oLtt6DhWi6yaT6w98iar+ZyoUiZMWle1DdMSMxfu10+
SyP3B/sHQzMgU4OIOjbhSPOLRYOZetw80/xGrWV+wn6th6KTnCn3Q4OoYyxDnxo2
Hi1Y+R1aHmf2Ioooi1B6/yCz56+dFIybQLid7/z71RzgWxRhNyynO5U5K7Wm0dFF
M/rP90+FsoKfs3q3tLn2MlGuN5HmRWe3NUqC9Mpp8VWgCFKplcKI/QxlcDNr8+Vh
2pQuH7ZKlexYujsZsKBwCWwJQuZ5cD553wkdOXjunNh+0w82T6BmDNtLWJZ9gaLC
UDp+Wft/1O80ONbbE9YXFjOtC07FofP4JqoNrqnDbMFrQJKqomr5/lrkBIh94RP3
aIGzNiXL3ONzXNfCc1h/okGixPASaOob6wgHwSQMsnEllc8h43qAMaTzlhPhzwqy
LFiJxSEw9Vtw8T2wlqpMAj0QtNx/PquCKO8fVHRe+AbDC24hy2EaFp9altqKL8bp
NPmMqgmJ+FPxuThmHSGKE7g5i576rcaDIoxVSzWvQj/PiUQe9D+/iiEujuuKgaB2
sK4jRxPtRfaojHTPHM06Mc4UDDCfYqFJZtDGPD5koLdsmIUvHLfTA+NfWbXJ/sED
IbSjP5ukNayseTOKMA2gkDq8mqeHiz9y5Gg1k3tDtZ+cx+ISPkxVCJuxko4BOtlN
ZyXRyEO6S2gok/eEinKvj92POcBoeNdTHu/FNVUTqIJop+YCgl+fN8B66xjLhpHe
rgpa1Dlp3cQU3r8R/7+KzEBr8FFfDbJlxr3dALqqAWrX4wHWZdP++zHDotSZpND2
OvatZ8m8JSFy1PRQ75mm/e/5yAu/Hzok0F6xjWZhKUizjMmkyXQMS/Pt1ZrESVFE
q3x2GSt9yjU7RD0kcmJntmpAdUtQbNknqKVnv3mxAn+tctmb8/2h1BDvFYRWrm8r
u3Ph27mVN/VSPBhoWq+0oU7UrzBW1mfSu9lH8uMc+3COLYbmaZR+LxiNvG+naKbx
6Ild9Behp/srUeet/DYW3WApacU7G0jHrNF0VXQIZ8jBi7GUGKtI6kLk3IDrNHO4
uGuNfs3fW2WwTBgJX3YhkLbvy++WW+iYd92CiBiiZZTU7QsfJeAowHfyg0vPCMVx
0IuB/spCfjKE9ZXog8Mzyr6HxrLmPmV7Aexc44Yo90NSM0+amNsi8X/kIrVa73ys
ZBc13LlHn4AZzMs7YTPlGoxZb3Q+kSXc6cjaTlnPXph12cRVXrpK2vNVvYhxfZVf
Hr4HgnQL9gNYsWok+XJPgssziOrOE51zrK2x68EFZMSFj3QhwZAG9OJmFIzjvMUV
PjvRQHt4LniZI7bUwvjx0DYicmSfeKnZi6k5mlPWHKVAMahmLjG4ULZ8ExUVL08e
YAuwjyjTAn3WkPCehOLSbq9wpTXpSg1nJ45sok7LRPSuEyDYD1di2W5Qwry7kKL6
4z50obmUu2NBLHXJYoUKOzkEeXHFFOQD/IAdxZvMmsaX2RkvXeFVh6JpAiNgUVDP
BgEvI7e/+aU+1fIy5FjGJEwIUnzcLLlgKeLMtvXk82VBaRmfucKKQO4LMmgMr4yf
gD5gm9q5zBX5ZgLnVOKzb1E9XATziysRcKtekNSpD3lETukkdaEJGwuVDy/1bwIY
ULY7UsqgqGysuXIAOGq38/8sIV5V7BHxSMnG9yBF6QKZZIpnmCk98GTwo72bR/Wt
AG/1O1jSJF8hLza5Aq4LlEa8WsMZZo31qWDfyvYST5o4J1xNeIsNLGZYorSw0asJ
daDg74hL7E+U1iNTUq2uCKRdM8y91eJ+ixtbtZolZTNAZq/8NAdm/6GPlllluCsq
t4n0MF9VYE6/n0diOXYCLxS0hhQOZyQjLo9jUfQTAbY6hdTnUsEb7FxV5ZWsd0He
OXu3/Z2jBOSugC37YsXiNbBGzpKNDgteUP72C4F0bHKoubMiu+oZUbRCkikcMwsW
mAFOuDaOnHLVvU6CEoQqDEvMRWV1Ll3lH6BSaJIfxRBSE+etdpBfReuFafEJED7+
Rch9X+c4cJviYyj1cDwIB1eMGm6DDh5Y5q7h+gc2bkfid/MTQDrGEJsxOeQvVgCS
JneftTsCTfzC3nCQfFosEmqirO4l3C1p+UDvfQrI5V5IntlvzABEKrbcP11qzLHl
2mp3XHn7t7FfaZi5JJIcXgU/D3YwSjTxTLpAz6x5fXJaQATT5XdAfYblvssW7t8R
yWVK/d2XH9mGRb1f9c6wrZha6dgqCC6H6yr5xxMLr+9Qy4YsSnva7IA/aV8iisSi
7r+rpkOoWiJzlVvpmQfqeDR8RBsKPBiJeOWXkXQYeimPH3723qXe2vooWHeD71Mv
T56Sqo0h7CL3OO6rWz343/mwjUfb6U2KmI4sx4/D7Ilike3SW9BL5Q5q4lJc4i/O
xL6rpd2ZHf8rm1RuX+SjWtF/mngh+WH8GPs5H2ywiamrvP7thoAHjGkh1ZBkHCWc
oLyDBJh5jz84xvMXI7gSlMQoQkNL+24CtbNjQctirBdgF7V3Hous22ave5o5uZeV
s1dC021mIrEqf5TX8szGH9loXZimIRLupGpGB8IdxgXCQnsA1ijZ47B2IyHSzDiA
gySXec02ylckooJvcuGp8XavREUYsOMhmTAHqWolEirzDHISw7DiQ+62f7/kpBN2
O/WUnzDjWOV68uLRMatYyaY+M5SpZgO+6diRSOagvbC2RRY9P+/sike765ABC5yc
7KUMyE0hpcNJpEbOjLjr0ZX/LssRdUOn4xVoEZbNAh5yXPV64MDIfo7JGmIUjZJ2
GrkDWkQKk/R1ICpLaDiixu31Uc2jZ1f1xAnzQQMK7M6ooQWBn7iQepWPcsO3sZU7
UcskHfO6KvypUiloITskYlIVT1S9TfA8RxzqO9iOYttxvb5MA5SMynpDnDl4ohz2
RTVGN4GZjavDcCrkWkoBYtzl71Tb/hIuYRG53yiiQaBJckONJUywbL9Jhlhe6pPe
vzK447Iytz1h8t8bZK8sSuqPWKHs/4gUAVzKrtBQ3CIDh99VJfW9lz4tOLyKuaZH
OiHSAWLJuEFY5s5VK4eGZX/FZtMZjvbYsgqEv6Jp58ehXNcdLMNovvYZR1J8ypOS
f/MPEFKtqLq+sN6XGB2ba+sWJjq5lMJtw2FyoLETZL/iexcoI9AVFWzrxR1RK9LL
sh6pJc4mdN2u9JsiJ8km9H57uOBFVMnM/4gXL+vFuxP9U2nJws6/ZqApGyaFIp9T
S9Plwx7BXbI4YZVuN7g4HFwrppss4YuGM9mnJFBn7E9VnEg6IdMvRj8QI7mnSm/b
zMnEzz460Gxv9N+QZhLBqnnXuHR+WBb4MYFcSg+6kfoHrPCOi4vtnRJL0w40Oziv
RNxOzk/uDYe0v/8dId0Itewa0WW61VYZlu/Q32XHQSp4awwM3/B4pDTVPcVW6BdC
bVrGdQBz5h4Btlk3kaUron+2AJoSVt+TjFOsp18TYw9nI8Ube2FA/Lqr+bkf3de+
y46qD8S5ce1ePZKVAg81gMSNMTQtPZAB90bn7bZPZYcUzEJ8s6wsvXdB8EFmmpnS
gdptxyr2xLvEk84Qy7pntQyogAqJfYkjEC3U4twh8DNzHvDzLBGbltOGMgT5ecH8
0iQOn8HmexcyEYxLxlgfQ4wNRLG1iEQbdgPr6jibK8UwlHYMR9R4piByDHwtMunt
3j8M7VkHyCfswO+ZQK2FWoWEbBKOVGk2sH0mLSv7yOkfx2yKKDFwTlOgDwcLNSkJ
yB0QQyYjavxj7nOJOM2OIDZlS69q1EDzy+vR3tbs5s6cgCy2bhAJgyjGxeXh37pA
ccIdrwDoMklIQzUWMxX/WskEScQxW1rxGZF81yIgHy+yorO6RZPMI8WOrzS3k6ex
KVXUWYgJCtASr+sl8qkIJtVk4pGMtczy5SrmNbl8KvflIZVFNDgsflTNk9G1KYVj
SBrCF6Tc57FiRYfgyZcxL5GDaXvA/vdDDGq0iZ819IjpTfUf8xy0eWncPjLtyVqH
pp9JuQJk0qwvEK9z9JVlPTRkQhECnrEZAPLIynRvxWfv5NcwTWiXw0O2+0a1dlEf
FJ//xVVZfumPYPlwXMvW6au2fKs1tFJHJrosmWugXYRAKAXmytAOmxc6MojHuCuc
aAvggPU2OS1GC2TZr/1nGEBHxnMwE1qMcxS6CuKRmYb/lI/tK7v0JsEZ4kjDRvds
bZ2hNfU2VK7ZWHd2Xglrm9nkHTf3p3HIL6Uh8RKSHyR2KYXNH1mU2AzQ/20rp5HE
BKr7CjyTq9uHYvnRhbp6/a1umvDlRelLpTaJkXZ9AIKVwTbw9gkw8wTHY7AsKGIv
8s4vQbc57Df3Qk8iBeylXnAk/YAtbx0dBzJMZYi3z//zxMt/jhOr2mac2Gj58kVk
D4Bk7ixGmo3Jl8m57r/Tm16zhEyyL/RLvBEwoM5WEj4gN1nJZ/HKHcGW4eF0M23Y
eQw2MOLdNa2VynFsZxbSNH9I0qhTTye2kCiXmjpGnT8Uc0cDx1GbSXPkwIewQr7X
j7rFQ5rXe8vWVSmJ4BJ5UyQZ5VCcH1YD6HGVYTi5L+iXJTvyqfypTwInrKxSPMh0
Go7jprrHc4mdIMPY7rGue1DeXDheLbD60LlwEZ4fkats/8Q/cJrCB8ZXjWT9C6Cz
llUsCO9fp5VX+SBHOjBdDJ5YJMnsG3T2RVZEENwS3mitAbBhUK6HQ4B373GhO+OX
oBu6pivOvzHTqSYnOSNKL0KEJYOn+henRbcUNk0KWdlgb67ANU4gBGuK6Lqo9zAk
+QMuPui4LLlERGWdalcafeL4+SRMzaZjzw9JJG8kuB31jFK3GIJFJnv+tujRMaby
s7r9iKDhOy0uUcEfWzRGhjMhn2dvYI8E1NNsyrUHHZ6zpyjZd6xaDFV41eOOhXjB
ZnlZQN2exWqpeo7CockShCmnegpIAJPGxsu9ev4V/hI+iiVtx2M2J6V/1c6K3B00
jYGFjh2zuWzwy+5UT6QvLFFT84NC/qo4GcznAw21gzWcJXsyrYIALD1mqhFLToiT
rgpr5spUfICwutk6Ml8xsS1H/LdabuAfk0T3JcUWKISnJK2oztBRZhTY98AinDAi
gppilet7QHC+yKqIDAfmyl4RodU+G5wmZOCXSP39w1dr1FphAXnnzpYYCjyqF9MP
IrRrcozP9QiHkivtxytOCKj8Es1F4E2x00M4K+3r2tiM30SxftrprE7r0xqk/xGI
8osn5ldJtjQa7AH3l+Uk9MCXJD8WEcQj4fhKk4uqyI8Y63+5bjV8Xy57ZLjxUhTa
aQyprtN8q7jg5XfUzdI298HUloiWmmBjwfuepknTBwXagJ8YzIBYsJwGzmbRkOJh
W+VaEObDBQqIKuVyius9EPB+5SElJVDI+d7F+iR9BU6dzX3iSLaBtspDfT10mRi1
Q7A14doV0whHHGua1oELgbNoEV+Xc8KWGsdOqo64PuqIDhXLFRcnuhXYBDvsFdnH
XWTEJQmATbJDnchyWJfGq3QcTO0PzmmcJ8bj9PHETH4lvMZCjKx5KM8XDvVjNszS
3Y0f9+2ZUnsLrA/7HAcnc+wH/YOcS2STJsLY3iAPPq54q/HsChtrYpf91qOj+ZpE
bhLDrcXC9wSf5C9LFq7Jktx906CYMe1WED7zUisucBHzAHrnlBQzKsMtagvXXWj3
K+F7HazckRcq4XTr7FNwWC2atgIvEK6aeuj8xnSI1BHoCGSMB8PhC/cnW1Eqfhhp
fDU/QLlWhkKwIAq+fZkX22B6zGqT+ghrwoxUT0TU9tS8qwPpoanjbbw0795nmDoJ
rCLPagRB+wi10PZQNN8waWVVDo51xbdi0SS6gA2qQqcNvEKzJG/IIHp6AFFiga4N
T8Z35Kk8kO4wpYwU8lpneia9PN03F8H07EVassVXE7t3KxDA5AjnDxHz2X1ftiX7
QHHck14kBGKKBWLu0k4/pKwv/GgDAfW7zhk07pEQIQXOghHa1UBxwaONPdPgND5N
44mX9K894TKhy5HG6mtnI02DGNHN7a4Rf+EOBv0IDcDCZJAFEZCHfncSD4/xEkYg
PaINFn+SLwFz8yZhn6+F5LoL/hNItF+cRsNS3UqXdhrWDKEYgNrNdI1duV6UEjIX
v6sNQZW66PzdHfhSff0Sx8WhoHAgHC1w0Gyp/fYvgA/dy98UCDquw142ktOzt5FI
i20r/q8DDmVZDHKEo1rUEmx/lvGVpYBvUzIhiDl8hT+ble/pIAVpmiLWOgXMIjvJ
s5trAEVYK0k+7SxOPwOCj4E4GPphMskK/eLV4NacL8arLjOHvWukrPv/lXmrfe/e
q0jJr8hY1H5xtzPsGHCwJMfpNG0mnMUHZMo0Ra4Ri07EjMDIXM2EPEewX+3qDzuI
pneVhO5arqHWzYq8cB+7+fiEYJdn0NIpnckEuhllkL5k71uva3QPB4ztpyvk0aqr
02fSRANQkuQ0qaKcFW98DS2fmoiVzkNiC2VE1tDLo+qq3YT7nJaOsPclUwhN7V7z
waXmbkHkUzU5oFHZgaktaexOzRWyGUqcPsm+Ye3bwmB9y0yTn2hdQgjGOMvQg8XL
4h5CNQi1gF7/STv+mmL5vQlduYMm6Q0w58eKjN02Hh8vMFwSw8xLFio7gy0/5W1X
VVd0DToyhtLlh9p6gFpB3A93ARbjyaUDJbOWRGo+vuINQo3tKFHleApxV9/IwbZj
Ebr/66H5N9iS+M33C7M66pSrc50iE3ZLr3ACP9Jpt/gMP305tuWq5d2HfPCdT0AL
ilMxpGkoHqmIYZVUww18HjAHaZLwg4KAvk8hehOK5BJMZh5qA0XfZYqv9kC5Ryf6
VuezwgQSNqrrXF7qpDLjqSOXRXzTsEMIOLRW3sv+qalAmLFlsCE4wWfoVUvaOFkS
ip2ZWnpYpNRLLoLFJ5dhvCU56n9TFtKXM+IytqbMvhsZ3WqqTwaMig06QvBvumpM
SxBdVFhnp9zepGWsppoWQeA8J/RNR0gTtZAHgBpb8HzfZo0eb/5e041C7O6jALvL
jOlKGtyCFXHhaE0HPsaSAIYGd1TocEalldVerzDTqT3CKFGeQq+7Y3CNChAcWgSn
CdqT/WBR6S6QoDLa3FT2QaZGzuajcX73gNyY6n6CRUEqTAvUYpGx9EuUFTVyAqYW
vy8vD3xTv0D320ubSoWDQvPnXEPm+ZGvr+esQYH7e/9PAnWD4wgvYMGscV+19l5z
xO2vaUBGlmnJSmg67S3CZugJdYB0BB43FJKJ0EzXLx1dxXDtzVw7UbqZr88hnCSY
oli1XsJI9BitDzvFbxKHaCaMSpl0Dz/abA/2T64heytIx5Xdc47zp9zqdqf1iPHk
yOCqijs9r5UyR7GxzWVsbhUnHVUBeNSDow8x+L0T7DJVxPkHNNd58IX7FmzrdfUE
EBnggMNeIlg2i1reV7DdTwx4zpQ+8k4kifiTeOHoXQaC5RR0rQECrhzYk8xM0ZAd
JZyia8xZlNBhYVE4thIsc4FCceEAlzdwmmWUn8GKeXu9a/Cn7ZEQ2kjK5S53Q6wv
tNxFLFlIvrPswbcHuC3htqLvrdFqiiir9aYVqXvlDmPy1mtveLvHgjHKPhhyHPXK
hdsLKpTI7ymLAngHTSI6uZnK+F5J9YBeH1UAJz4czzMO79U+sGl86H4iqxWfx9h3
pNkrf/tJ5cXZIGdhiooneeQIs2T/lxw4gQCsv85w3Ufw9A1813z1J9pkgmqXQrmN
6ygLWxjbtCAmO6bJIP0nXWD+/hcPkfxC4CvP/6mGke85OVt4+Fp6QrkVAoCWGDq/
CKedrpPLXpSp/0QIQpi0XNh1hzPTrU+ilCoEBpVN7ZWJLlM4r6Hs4BvjC3fx52FD
O0TD3sqFft746wZRhuuwz/eeg4FBSd2wO9wQCl6CNRPiTvD1nWAhbQQonemVTTKu
Du3iKCq4u1xqgf8LucZQRA84SpCWTsfMHSqMtkMyPKsoFi6qec+Z3oSuHK1tPInm
FpbOPOUtwmj9UIhyUBDU3T/mA3evM7oecCa+ytUJPh0mz+E0deq4o3EkV7M4fDrH
CBAI0EMqv0B74yBXnvHG/+Er2hMbNCcEMDnK+A/uBi+Ph0NU9zkWnTqgFNg7Sq7I
tm8QYdiup9pt0TmCKJi4V7i2/TExUkOz12EC8+8jmhW8AiR3jQybtU0Gg8f+N7he
csk0wRuKEnsledG7VgcNJp+6vbqQHn3MhSJ+jBIyMYK2RtEypzmWIplZa2Xeip+H
2G5BKeTlcToFQPHq0QUNCCmFBMev2bldj/QUdz7K77lY3rzKj5jhRwFBu6X4axlj
MlW2Ir67D2FYeZTwDYQtQXrKPIToy2F6jXfUHABAnsALIIEZ5PybI4a6Hx46ZeI7
GkzIXZIWL7YJiGHTstfITUtozdBIxsIq0dGsXedXj7YfCOn+gpjX2N/OKdf6OXzu
GYd+JgW1aY0iTPv+yWLiVowUoh7bT/8/gUuaSJ/jhWgFY8H3Z9X1Dyda+mp9DBVT
dvMV6BsWsQwGJSgUtdAg1fIz6mPg9MYvCLzDfUfl24Fe5HOq7r+Jw3CfL7uQfzII
VrvdhWnAlIXlNjoOJdwSAtrWxRPZhy2xZCg7ULAeqZFhqW0fGroQr4r/BaN7M6on
JY2X7zI7230ziXYn9spqGKKm18KPjcSGFC2lrMBBNRZLR3cR/WOAoW1hVGydF+Ta
FK25/oYtsXYXTE9EmbEzi89EJTWcN71uDhLTCWINNp9bibfgN36QwTrUukcaK1dc
2t3SdvkZaXHP+d5rF6mxsSuIqe/H5+uoXwqc4Q/Vc5BqpKj76pauzZ2/pLxbzjHG
jf8qMBaR1qSV4j57OumEqTRTw3my+DJ5nOxegwiE9yDlAOPjbs3lHXSIG3lmBs9s
DG8WzEIZkeCE+ImETOIOUaHqnu2XdS3SN7C66CLq7agn2ZV4Xb0QrooNbh4MlLsM
uPCIPIawL2vHvXtoqKxoPDIHvYI/dsZG4t/32iINgegJVhQP7sgVMm4BA7wW7bCG
2mhVVWkotlhWx2bwTXnxccD8ivNzzQqP+xWQEZ4wTS42igs0sP05/T3b3mqDqsLg
KH56lf/gJzZ02cf4dGGHkbrfjrqcltRa8X5dEmp38buFHDJPB04GRnW4cF5EqZIV
RQ4ESnA9FI7rw0/BOVzZHTvsNIFz6+YaI9k8Boi7LSwqCS1SNfjH4Gir/434lck4
XDlmwW4g8mSGYkyX+M6bfXyC7k5XYJqd1V7VSZgRm9D6O8Dn9K9uXdR4dV0/Tob6
xsh+obTCEpmIeJAuuWAPtJ80T4JEAe/O3Y3QltiFB9qXO5fBrLzWOFaCIQcnuhQZ
Mm+95p9oQdUf8lvzrLZ3oZYhEzUw+vLTjU7Q/X5owq0vxSgVFE4J9I13/hsiMXHl
SPwDSPFwzu/wls4YRrj2dF59OU5e0O7bW/GEre+ZDhOTMeVopsQ0OvyIMNpSh0Mv
SFS+/JA/Kjr4B53Tdzf8rwGmKKgLuNTAbFBarCpE+GSfZAG3yjasyQQtNT0i/d5f
BWXXpE2AZ9++YGhiyO2ciJuEZPx03S1+f1sgPhy8DDX1l1nchXVWYBpqAxgwDNxs
HENB+cLDEyAVBswaEPGnVi4CnO9iw9tFLbY1/Nh/Bd5bAcNQak4sCrKaq4VgWRk3
d4jyfe1/QKA+QNhLJp3DYkCtM7lvb2LAoqM7XisnlABBXab7fCOQIFMpRM+hIy2u
pGTl9v8j3k1FnaEtQ2mXx8Jem5EoveUWLzy6dFQPuRJtqI+sKB927OdmZO10ofU5
o9sDdDl6FtIma6/lvVGAsiNvjcN8b/jeQnVzTGOJ2il28uKG4qaapjzRxDi6kDSY
is98aqZWED1FCsQncJtM+uc5cqWDH88E2ZvBQZILOsc5OWZp7o9vSoh7qJkXC5wB
fTrYtCdXvLkb91R4dbtFj3wwmFQVbWuLo/RsWiukRcSKAjHzKUllSFe/XnRQIjeA
vxKlahaW4Kmwl0Baf2mg1EmVxe8WiVBbS6owF4r2m5H/z3uSNaldfX3aDdSRHMsM
C+gb36/kJISJaOGr+0X9j0XalkRZY5K49CPcHeKnSWiTp/N+GO7zmwxZNhZfNTar
jRysJbH4cWgjRGw9I6g1UOIBEE70jZj3wE0yu8b6bknxCmMHXmtY4kFXIayxx2s+
CjCMO2fT78YoCi4XFd97iDSrPGU7saZBGbDMlcyur3TD5ao5u7sKDtl8ko17bAYa
w8WoGotyLjfRux+K6nJ8kC0mDdyPjeebtIWHUdBkvB/NSjJOIlubDKkh7Ey0024K
yZ5UtzWLNPfAveRb98MeNdEEW0MJ/o6sKY9voAWFREnV2TE1l+i8+IvMZuXhJLH5
rH1t/Ogr6ppaho0XlE5mNUL46autJz5CBoQt/WO7wVMpIIAxcvU6wfCpA32fZ2qm
JhXai8DFm9jHvAlJkiQULxDoHNjZV7rg3Tws2m3CU7EDmj0cy/YK6eQ6VrNJ1rfq
Ip1XLkSRm2/BMc9rov1V5ERus+3iUucQMfp+OGlG67MIQpDfonZvc5cotGwXqkfc
igphfO2VypC63bqNu/3FqgDQjdxz7tUfjguQP/QwzxGoZ2RDPbhPv/BPGE+rTP1w
GX661HbmDytOBGHpqBhxd39uc0YjkDZIgM6y38MS7MXTFvldAtCL7pxrSnZxoWdm
62234fcpX1Xp7gJoo4brCcOWv39KYVBc7cxJJX5T/L/fF37HfHEYamErEhogilbb
CDYow1zTMV6C+pRfAcI3cNRPoE0FccsnuPLjtQko6z/nESevcghahVVGiiRjlqPb
wwItcG89SYEFdRi6//0iitKWJc2KKqPYa7xzSrxfr0abqPuYtoywKbPRG+jgyFto
aKdbJIjOQFSD9H5n57DGaqnyT8jr9SFN6U/8YJzSUz5IaDXJ1jXf09mYkNUyva7J
xbUXcydQ52ISmcH9WhSdXfR4Wht+PB46sPYkFy76t5ISwyKimcRVt5ZPjW+8xXWq
rdpSJsAaIG66+elPE3qKWS7Fvb4aciAtpKboyWS6r0Fltwr8GDe3pZRlmNkuhn6J
wYNA3yAy1PrlFOlOdaXDUeTHqb30ZfnSE4hbee8QZebcHgDcVgdqusfcJMqEywyT
ga8sbUw7MuV4WuUspUqPu448ftfECYGLuHw3W36H9tQe80EeYGx+2unggEfekodw
Ff20QNg95/1VCL0128QPz0aolzh53G0pbhKuBcLGeTpDbSd6zuJIn7zD7zV8mSiG
8mDeEg1OLVUbiNyU517LgMZmSmVVS55UB9+W4t5ZHzeSmXWonDjpYGak+p4Ssim8
Hlfy2P4Vgq5S5LGDXRDhMX3cWwV4Kpae2jjRME4+au+Z2nQEngXT2+riUWCigCPj
LWCaZeuLCQ1IXcxXwBfByK5T9qiEiQSeJM9ZDd6j1MZc1oXrX3fuWKtgNAbd4Ah8
aO5bOP+aO2WRNpfVgHu6sBFcPNRRBKA1vWIqeocHPiU3O6+3Ftb9GM5k5fjl5LXS
cUYAGIg4AN7WUY4vj3jNjg93uy3consxrcMkWP6NdMeDc7N7uDem9PUeSm9wrrBm
7bK1VG3JFbpNxPlmY0pHSTZQTYCXe3FlP+05CASGNrCjFGvEYAd2cuPW6Uj+xly2
gwPo5u9dtZAaAoZROL5W8+rOhRx2m4YDQ7q4v7AJkOuVsDaGuBQ7AncZ7PROuJbo
iFQjuvlQ46TzVytsKdwu7O1tl80+bUUTtcYbcrxqRzljIVP90KBBTAg5/thDD3Rp
j0vQnyn0C2IAuY4zFSgCEJJ3nXl0hB7Ki8sjGcX962pWJIvPuYRSh/Ol7oEnsiaC
uIKMLEOUzQjyNORlk2aGAJwhjhkFJ8BZuxzn8PcHCUnGRr1Ejvn64v94H1QffJKy
DfugqAaCnwKA4pDS8MFKMDTfnuc0FgXLmm6jrA4jYBmA7inZqeiRgC/nMaU72e4L
ERZ4RLdmkAkv5UEn6TZfV8+CAUY0/1spK9A7r+aPSL9yfmg/6lUfIDoqY6sLlP48
OyLtdXA2Jcgs3IeRhpIxA7Djc1leGPDPhkNUnLr4s0um/vR9uJW8XJTkUgmVCOBA
0gfiSoIZKaKSU35eq4omgKIqJMh7EQ3EHXxT6l8ApL5VdEp8Vjkn+AABGq5mGPer
Tt7SpE4reum6bonDbBz6tLDKevp6Y7Rp/P6w6SgqrpQ7DWtUzLvVTV1umejd1nwO
enRsWRiEANyDAIvNCVQgIXPn/syoOPb/nImC+YZZMdAGAKBPW5vvnb+wFsjfnIvf
cE4IcPiE13p2IxWseevjCeHR1fJcioGJsJW2jjNWZCfZvU756eVUOODT4li88oAs
ejo+oki5jFuusAC44nFP5iD5colEoAyCWlQTp3lAMpWAy0h3eJ7MiLa5TgGVvh5r
uznLECnNhurk2wuIIO1AQosYpOss5toCURxP573fx1yeeXuYJgkUL3JxScyY1XvW
g8C9zyyquq2O9BL0EePuOOB35GtTWNN+HXVZh8nUne09+yqOLMRoyD4HCxGL5nGw
m7FLVQxJ2wUSKqJ28wAUPcwnj+FqA9MQYLS7AVv+eiF3THkMCdCEagMuQDtKrlok
4N3b0/lZhacK5tBsa/Sa1mrPSXBAPvlzIXRKNO+NDzY1dVQSzWiHlHmh3uPjge32
wsDYL8Ub+yexBNZ4Hof+k3lo3sBaLpY2Gjz0CISFq6hLv32PHg1Ruzri6MjCdl9B
xxpMLzFNtsnb0pwYW8Ort7TxQNTrYfWhlf+xuI+jc4arRCFizZ87D1H1b94kxgIh
CjE7f5gIJ/vM4hOZEugGiQyPOnh1u3ujCnguj57ySUYYTS401BIdySKLGKxbMuI+
0XBocnSnZ+h/qW0H60zjZLuRNNPiqn1GkiTh5ek52VXcQ7U3Kvqz+Urk3KTqLCe6
RuwfBRuzdkULt+RokNokZ5JyZ1DUvSdXEemIoAFrCvNIYlnU4CocUjCBQcrLRg6w
P0BBT00HEBHXwj9eFCrwbRmPq4gBVOfg/pkvNVSXLyrrM6CrOxldTmtMwRE1gzX3
4cwn3iK7v4olCwaaz2Z3xHcor5A+t+ErIzMtLeI/uVLKZl5qeThfvfv01Oh7AcyN
braozt9D09+CCZBPypTcI/KTUb/YViNC97Liz5G5zXdR0wncvwyQygpgBsfLkKdC
cNao9B8FIn97K9BZcsq4cjDxvqenqJ+MgYVdOf/u2CS0jId7NkSX+qVDI9kkW8k3
2mt3KHOX/AaPWa0GK6/nw0nFxMBYlRv/bOBDdKPRwKFr6xg8V40DW6CiXHHfjpB/
R8VFx5pmcKklxykWlT+k6hFpGj6G1GKVMMHsx4N3dY9EQ0CMWffmjQV/RGN+yDUH
w6wt+Zo98qJoGBIovmJ2ZhRhMjvd/BjuIy4c/7HTd9d6RxQmNzENK11hcyN3i0q5
tSfOeDxb8o3lWIvz56RDJxhDnEiSVoLpw4oFx6Ld0dyccBw6K+TE2hUuiSUWfqwW
mBL33PAzABL4XmVn7o1afVY8xu6BMlz9CuSf0tu+2iN83N1ud+WskTVRWkTA4u+H
kWoSHZY1uAtwOCV3couRJkLYgELaIIrMpf8Af4yuDjR3c9dvE5Og7/0rG12cBqyM
OiPYXiKUmVe+1HQFYPvTWWKUQjiHfLo3JB+YYsEyE9WmNmtb/7ilwf+8hrgnT52S
rbbf/d/uUgCxWnWO75GRcwHV+K6B/Ijye891zCp/qOqSL3jtUnQMWc6cw+BLigED
oiG6oOTA85hro/RcrmXBaZiQ1AkM11LBy2t3CMwg2RFNgIoO6ln7OSXzej+pOgVo
+JUhmldfgAqq1jqCq5u6tFUFcpBspn9FEF6CEmLNHec9aZeplzb1roLuj1WNmGji
0FuBGWlfON6O51GJweRc4ZBNQyn+QdwuMyjaqhI+G+zYxmNHBerKL/nukWI/cvK1
Y+sDFk2kjDBFpfr531NXtyjZA63b92GNroH2Y+AZQy3Fuyef4j9//WdV2y6R+Cny
/Bu98Qqr6sUHo7c01fhhxa10TZzhLnofdg1CqI84P5DBxShI1Kcjb3vDTQF1442l
hLFX9WAkNELkpvBcWMCxrLDtPNd3Sckdly4MeKZ8fnl1wM418ZE0oU5Wu8cATWTj
Ahg3HMjAn2WadHM6RBxCm5qnyeF2drvO7ka3hxzOelKTLvPwCBOSioJmZSWs4aiH
Jw/QkTRPpeM6WlkTy5l5a1HL4uZroXeoWzGQWs8fXdwP2nUh400RovayE3UjROF1
fDkWNoSlkZ9VIFCoIeT8ArFz2mF2CktfeJESBKd9fla/vyu6vZljjSyHxokt0PUQ
npAcncgHMkeQHT3qDrVw1EkA+8pqtZ044v7EPG0z6fTpwnloftKkfnJBL3JkVOXY
2zwKKXGWBN5ZdE35wQmRq8/lFCtKEshXfZz55LaNP3Ob4r35CMtLfZi0QlWaxI+v
8+7iiHI15ZQnYjorALDCJ6uynjf8Ks1NfIMPYYrtmSEkNp6ll9Zta57dJjtptEfM
0xpRBQEe5d3PK7nZoVEjbmC0wIphJCvOILZ+uHYheBoOtFyXoFgIMSvHJBIop+GX
rsctnAjq0v+CnXXltwIZZMRmWFvkj3f+RSwot003kKzUP92U/FrlIEuNYfN81UdJ
dB/zGvZ01mJyoS3BNm52nUVT6giGk13RHCFJGyZzwJnGwLINv68xUDz0KXxo94Xi
Lot/8UsQqX19nDkZtqr6p5T+mriIlGX1cL12EO2KnAwbnPaKYzwnqhJdQGjMPEBj
6lsfSGaiFwTnTIC3poVnBpJoSKwc4PTP5a77eP4i8RutwO3qxyygJKhlIypjnTvS
RmYAGr6uazBFTdLHkoZtjRj4a9NOuiGRdXUOBg4alm4aYSmb7cviWF3xHrYwBKb7
MF/6nF7rnf5UWnzIunmnaVOEwrdXuBfvRMjbzXeVmG4XcvoyoiHKaeDq+l5CT9mw
WTSpLXnwmjyfDc7cSdIEk+whCYOuHLwauTApC2jwcxApXpf4FvNaUIY5PAXSC/+j
cHbTqh75LmS+PM3zMd7wwkmxG8vAJTLwtEX5hLNJv3DGUahTQAPtUxtu0I+Rj6w1
V/5bAvrP/UVZFiDigKkfGvZgi4r50zH0JEPdbuz9lC60PBxuWWJ5cWuyz/aVx/Zs
65c0UOQ7rheYPkIjiPf24yh1ylq5RFyj4PxIxRecDZxunIc25lN+7BRGOcL+1a//
lJRGKtlCMim1I7EMtKw6vDc/q8FK8H5EOb+5amduK/5VFKCwt7VGD0+kYC6iU44v
wxy8yL6vwDDcUeRVyIJRGKhNMU0v8RVbaUf8Nr6ZafEiN1SbrN61Mv+BCEJYHj8o
PciQYm8AYPDnHs0DAWv/XXl19YXCy1Y1TyEQhwqiuPAVZPd/c9XzBBNZlzUOiBaR
KrxZ0qwxtxb1muRlpav9/URCkE+E2nVMasZ/VBlAzB9u7VHrOF1fdR9ggpPAyuAj
dfZWDR3ZtoKo8GrmdOiMADY9K1RdTzQh4lsP0UbOG9yG2LdsyARdDvvu3FZWbniu
tXkF2sUI3nKMJBiYU0vo0AYp8grZuJYPehuxJgHQddp6MuLBTQFekY3SoQWVkIbo
7dxJ40IRNPrneS3bIIlOUhEAqhwwdwHOr2lC1IDO/kNS+eJWct7lD1uOccV8Sscq
KVGxNI+WLB37a5R591kva+FSDfZOZcBDG9IAbWZ2L0oVALR0dQ2FAlgRsxOP4FNT
rHedhEVPJ0eOwO2OeQfXQnj10AVhlDCpDOU9tOBErKPWJdZYxb6KcPxU9sWUD/2g
cbl3uyni5P++Ba15vkmeslKBvjh9BsDI8jBl3skVMrgz7aFndJJy9Q2jr4aDUCXX
dTYqeCADmvIYvtgsXkOMarbsQmkHojP+AqLoYH2fqzDferMZztPJSDOkvyq5USaZ
W35+PZHCtvSECboh0UIGe3wCbb7BZzbD+1C+vgG/jYeclTBrM4uGszdsMghQ3ihQ
v5ljF0Xgs3XW+K9bc3O8J+tImO82rAFuT+2QKaNlTOZ1/+jLFJfuNkxHYe3IMd7c
6ySUrMES83OqK+eNFaPvJJJYjZ2m5YVFbkVmCW4N6aQ0ipmrkga7gp95nAxySH9j
313EF/i7jkcSo5TtdWx4u04mAkjFZKXKfj5pmcrtIIDdLJlnFMj7Q+dariheqYue
9u75L95yY6fZcQqrdRnQfIIi05O3Okjn3jrYzJ9UNTaLNPciae9EBN3IPI8J6SsL
dULE6YClrSQDlSdXI2DRkK/yIRrRCWqAbGK15icsEy0a3XBiZLldxooFaXhqHuLf
zd7NN1n6Bx+rti+UwzEMQ1gkrBL4vFNTIS/mYRjj3NP0FLV6bqZvP5HzB2FXc1CX
ODE/Q3zrJY8LL/EgGNc6BpimXVAJtPpjvc+R7b1wB6BLFbT0riGxMFBtHvGWdasU
4OlAHi8QldYd17QPYbClCL9pY5GBVjtB0QyOeOor4wUNbqwQtuhHDzWdf/QuDYDy
UarzXGyO3Nsvdg9cI/lB3pFARrVWKZG5txrZeZ5Y0p9ub5WF11ET5cFdFTVKLxqI
woKSN15t3vlyvTYyhzGn5HPGWv1UI7N2Dejw7buLj/udZCMf5gKeP4NdGGdBN8sv
Sp1CKyzuy28LWSdaspiWyW+as5gJ3n33j3zq2N8kMv49rKAtVmuh1NfNYzRBc4Dy
ASxLSv6jJdvmOiXnfr5hNLM7WwjOCal4g+CNrduDqbkfJy5OtQ73HeRw4cBU7kZQ
qfGdYDZDRVvn1ca65H2MpVK2jRU4A3G1wxUte5e6Cgdy7ux5QvGzRPgp+z93695t
HxMaFu6UOoqBAECNljvCifRa7M1eOVH8SN3fh0Tuf2HwZq2M65orXzkjfRbVgVYB
JwficG28uQe8HLReWYjkO3n0TLlqVbK2vqRTeVQPThfEw29hhVjHkU40ayVS4EyW
O9hp5jxmVCSoVhe8J6PVriq28Cggw2y3zVPa2wH554h5AhCovF9g9Ly3h1B2PH2d
fQJHZNFjVkmae2JNSRI6PaknTJGV6P8rMjpKPH3CD4uLGvkcoXOJjjxRQSArQOgG
Ibz+VfNm5X5FruEru2zV2hkOBNgU1QYIsx/0rbNdm6J/z5WsDjeCD5bF66FkI54Q
5eOWUNMQeino6uHDc9bdpElTlgze9EWpiUw93Qz6YpAcS09wh2EwXDyahQJtnbs9
QtX792FCbvYgEh5TrPL+pn+EcBKQLHLGIg5I7RFMQQPBMVXRN8oqa8a1cj53uLk/
rsHt+rXsuPX+HhTbAUOyPFn0o4f8FjuInNCSbSsQ3ox2XW245U0+OKi1/KS5Gzfh
sO69PvQPvw+HDLn4OcZ3t4ERnze8oAV2HQWLa+AuqMLpJnqvBPW0MR7JrWxLN51g
XvIY4uWbzXzlpPhasW3yn31E6hWlndAjEn44V+7qNWf6lnrTBJhMa1M471Sy2DXd
/nD/s8TZ8jL7L4Gq/xzIpiOP6SEEbyy3j3/aESpj7e4jTBncOKad3NFEvqIJmHUG
o6bUuQLMzGxQvE+igQlRwtdyl+wjLwLE/e3cCLHuggWeigm2YXfCXiI3nohrYt+5
9bd29HK9A5Qci/5mHG8td09nflcBM+qAJLMddoxO6vY21dEY9GMmkl3iDe6hvSXz
DVvdH1poglTTK+dfWTeXmn0MPKVDoHi9NPGIpdUkqx1zqZAJ5/o8kyafgk9UzfF2
Aj1VoFuVyTYRC+PNBYoopLLm05XrfHUOzK/1249IUrIrVSYx9XTf692BwZmwomH/
d3FCTuCKM9etnTYOP8WMUQtYhnQoQ9Hv131m9jmS5R13FC1UWg80zl0PsCfRYM8B
GdWkVvEiYEtRoGgkssNNgGAeKEOua9r+Xwlq6JPaxDgEWYQ9rQxsr4b0vQRvPOVL
Yo4Ln0gCr6shxl7TlOy+Rg3pBUTSuHMeyG0Tk7v3jAjOprPfnlMyEjX2jXPodwLZ
HVWJQQ6pPyPI4mWpD5uKT7CSCoo4+JSA0WMEvDjtmnSPGAmBG0M0AN6bFzG88z+S
sIrAJi1DuVRxjWs5yJZq3D6rg3OvDkBgZDpj9PpKXbDeOw6wHOWyt0C6bphcwYhJ
FApMG9qE8IS2Jt8awBaG9JjSnIeFD84DW0jDQz9ADMvbKkkeIq0jcEEv9n7I0OCZ
ri/L2NkSsxj02VNkFdJQJm2hWAB/J54koNiYDMWgOTSXZ53jqITCslsWHqe8b+0i
PerlJAAuu4L54k4BevwCLZYpxHPBwpKOmepkKWoJ0IjrS2rIP8iiY4fr4JxhKcs0
USfNfwUvK7IN1aLuNDQdo2WJYXW9DSIyucJVSgFNoQJBUSNKg1vgEM/lldBUzZC5
Vr/SJPAF6U3Kmx26IchJgpxZeT5+IbTJ1CBn9nuUpHSF03c7+hbQMf/mcMigBddZ
/qNPYSFPL3aVFi5weMj/xE/Le7Z49mkSmH3k0GUvJK6PvghsVJJ6qtskXCabOFRs
LwyTuvteusX73zJXyU75BQy6tI2WRjIno8LEQ2qXxz6FA5E/lHAFtSlBzx46tjrr
TmKvyp/cxuS/NmdFEmc17AVFJFf5YGGIcilg1SMNYVN2zw2zdfeIVKJPK8ANeQYM
EqK0YTG1R3JTJSd/ClLWcrSrCVVFTtFitz2cnQ3m+0405Gi9q9uwxyqj4H90ejxL
q87milv6/HVXm0cSsprOP8T0c6WlIgY3L+OF9a4KHO788dRMlPnpYPrsoTAKwcdC
CrEs7TyHwYLMeXkZdlycQoJFY9nY3pWN2cIepDPQFk64fuWqWMQCZnln2c88uWmc
9Yo1hEAzcW022P5aEfhcBAVTAT4AXS2s4S1lPWU0ePIEMEPDKQqrE1GbrBpYiuYI
CjwRwTfmdRRWL5b5Nmm6hiHFz2NF9bRC+FanqFh+1uiCJSSLBRXW1RyfJC5k2UG3
0UeMJ8JM7uQCD26TOXbKKV0ulQVxKkiCFNRETTuLCOjlejyVDD7VviFjk8WdYLBr
4i5H3yTJipZ+ycrtaVwVSPFw5/iXeAD0t+JxMGPZiLfN/QbSj0xz1vmy2qgslKpG
CFW1Sh+EeNu4b/LY1VSpT9giOrlbDvAaQMt2Zg8xx36yHRwRCUqyl3CgFiQuttyC
d4n7GLbvxLGbTLv+X2i5OM1mkbfAS1eONiAWpvNtenDuxQ5U9AxkEEBcBmzT4A9N
23IbtQI9Yf2AWWyoKG+nyJ7kTp8TSzsVdOWguxPbp0r57qmro9/qzdoh9+nFDtkc
hp5YuYtRi5C58kQnnl/h927li1RV2zX5QX62LTZ/Os/yPz6KzeONgENO76jSnlRD
PsiccBygGvNfSkNJ0mRPCSG7tpv0vpSZY4+1YXRuHHtKeqx9Nec2CIJw1LKtOooa
cNCeqYbDmcaxn0ukUsnb7SMdl4EnofWj/R796PK7VNU1RmOlr23Vm7PpgcBh9gb5
s+Z4h2hAwNHGBobnERMaAS5DGSIyLK/d3hhq47qSd6Ygngt5ZM7ncCGo+NaVvNik
slSWyQW9yYmXSkdaPkGJff2HLgb0r5CAP2zaVSVcQdVTc5x61fIEH6N3S+OkhDOw
pfe4u38Q9WDZSF8y6h+yRskpmMzoKb3dITbPwpdrRaUOxGZ/Xj/hfS5JHmr+Fd7d
EWoXtQT1gj5ix0OPdl3nz2YYXOjGmXP7DDH1Bq9Pon7MmVpP55XOtdW8eyCStWWC
PcYaARfZkLLeakHJ/XqLVd0ddHZ4Tut59f81eJpfc33Wuf4PXUtltIJDCryuP8Cl
FeOQcELLv4q2b7tMCtqbH9nfgebJ8BID1Mb21DgRc2YcFu2Ti6pbAMLi0UqsYwWd
+fPWmjB/L535QZPhObUmMWZM+xyUEVG1OArbXkwd6VSafISGA401JeEREvqJBnpM
ryGdZr6soBaPY3lxusjMaFDalHGdL+PDAjAQknZ4uedxOt7glS7rK7MfvWYVLQMP
hSAXV+fOPHaZfSbK8+JzE6aceHoWLaLFCMKPtb4UFxa8n+mQpOReONhXMlLbW/6z
kyasdD9SXgOhf/KWlLfO8rKHnbx/LFONHhpYNp/DaKxuYOPdONa2RZUv9LS6lLVt
c32MgO8jSqroCA7hjM36mKga1qOwa3UqvgMhxeUk1uvQrldLsJ2jTyM0/0nwpbPj
zgN9vJRQ/2kU2GKJ5WwqJAN3Adr3ZJ8Y/5re5y/t0EHf/mtR9dL5y5zWQKRbyuWb
ZE4C2vI2cKfXSZlrISNQiu9lFDSkOIYcAbkYNNEAPboJasKgAkgFxg+ESeddpfh0
cbCJF886UjAKHGga/4mRgQU3lrsrDWTLMABCIMsVkxCTosx8sEheW/W0CMFMbvZq
tRvwgb1GKu+YAbIcn1Hz78UpDAcC1/og5b3LgFvfy+3JeE+15CsGNu/gv6Ss065M
u11dgXGIiBYAfAwBMiJLXyYeBNFU3EZB0KYSLHguVki5cT4C7ErTsW7zCk3nL7wG
TeKVM4dx03ksj4yUl+y1RE/OxGoWGM9DBbuZ+oLOLYMSCDDTVWEnIKFc1tQCsVxN
u9mp4YwN74fXN2L5johVYBlFFO19jB/1FbVT7gAQ5fIM9Am5vD6ACU5N6303Awd1
XC0hlop+7yQNPdN0Hae20vXfOa0Zkh3uwsghx6PEeIbVkQkKPFrqM5YeJgc1wPA2
5G6txItu1VLBTInBXKToDz+1t4KOnPyR70N2FMHiV1iJ9XKQHOVjbugu+G1ddy/j
ShlgYWZwDKIbxc3cPoXifcnKvz0NKKB+xDkdrJec+N6staE1pBjoPQt8vOdiuvlV
wPyQ61rvGo3GL9r4xuynYCe3JD8WybsFmKEEVcFY70plWvL8Jg/22WczNHefVRq2
jvaU+x3H0rg9ZXuQAx51ig3gzMNY0WGjAsv7qVtMrQRE63DV/EAF+WdF3lGJCvtB
5s+arwws8XWp67hdGTTuWFbrlXlFIEw/RefFfK/KTRB+MyMnzLzs5dJmSw1oglIC
wGsuHgg6CoxMCZ39+Zr2gQGqrjPMzVxhXBACZAKdq6BbottvX/pq75NNHGK1yw5+
mjuRcT2QcKSkWEgpyDfqQKNCskB5olpAWlKCKHpquTylOeOmFjX58owfl6F0BdI6
TSh+df8KVIdt52i2aj1Dow9D2JRG/HQ4FDcStgH2zrhiu+GFD1vliKbvS1uCb7XV
3z+YA8n9r2zsF1rPIeKCTsSpWy367o9xFb7PYYG6kENj11YKVYICc9spJzoDnCgc
gIciOjJGCoCFf+iyvdOECKaR87vEYnB5BjZy38aJ6rmBMWLFBJeRjzYPAyJDNOEp
HgLJX+stSPWP2XI0C9TZU8fMMqjj40flrSeH5u1ZyCjcLw3/tOcj3I9lGRe+76Yp
1KHPatWzl4ZkZ3vBeSe6QwZVrDNyalZPThRm9hLO9ueLoxh/+EwQRlDHxl+GaHg1
3XUQbmk4MJ+F8B+P6t3Ft0y8Z9FbmYCS1Z8WMQDwcPXTVxylXYt/wqPBuj1jflJY
jK2DO+U5bFvAssL3IqLXgWPkYvftRov8pGcUhPq552rzxnQNk0iolgf2IBMEwr4n
RCKYG3c5cIsgW2zChEjM/fzM38kGI5C9PRIZLM3Bh3sxJkvZvjXgJzX+dK4USKUw
XQOTnLfiL8bJiogYLO0yhl/1HL8RR9bssmU11ekm7XXJn8jLvMoZntgvV20JSsnc
NsjOUX3hQqmj2M2qFv2Q8ecVc9RO5qbLblhEvWlY6S1yvN2azm4N3EcVJGeBsPYz
BSmDyHPJAlAEVPhYTk0xxsoCZasieuhis/tqtmwJ4vpufCWJt47VkQNjAxRLoAsj
Gkcge8ilqxymmYcVMvIcuL5zpYRKodQu08F3LwJQfNdaZPVWtC0qhDqSUV5z6Ozo
2R91B4k3PCqD9sUIseA8IFyWoKQjBJtcMqhVWOelYD1vuzLcBSrV6AGd4ZdTyOYI
pu1D4P3cLRDEIWjcnzhTvzfv+ie7BFUoX6nJCLTdFcQ23LEcJzraOuGdb9lIYv4u
GcfBSYvpDmNeKjZOZehV5yyGSV4C2s+SlHPb04BKxm8cR0fPcWp5sNUod3KiZk2H
2nzUCFjkXhwJXkqCHczepUEcpb6aItKPoG8shkwZGezsQFbRT7yT6hORdiVv1V/A
Pd1/2sFoD9Tjssj1QgjZJD8F9akVHBg/Z+PwrT0Wb7U9DMcALDzGFb38rx9+m7Iw
Uutnuek8ZBCe6yNt+0ZOuK9rfeg+waiaic4DCLtRyqjvlVUxqBbjY6b/pFUyeO8o
K5XqwJMw9sdmV5ZJlzbC5nG4Vukt/OF9HSJSS/QaqKaWPC2+IkvWrqmhV7WPGKth
l8sAs1lnq3IwYeA/GkWSWmBiTEhTT/GBfiukHfE0PEtY4RQU1G7W5ZLsD8g5h2T2
Rp3GySr7cBZWj5F2cUmXWBClWchxFfIUuKJXh2avUdMKgBt1lC0JHN3/Jr3E/p+J
aKICy5lYWbj3ij4F7Me/qyJjta6z+NidJ5FutVM/w59w3Dx99nQqApizbqlfd5j2
m6rRNlZNZH8v5TPrryBRdln5Hk2hZim30mYfHpEkkEnHVYSAfwHbuKaqtSeBjtvO
beNKD7oRe+MbeRz1pT53qvIv1p1/+jp1r6xS65ozvkVzCc/VSby3Qh7CHo9W37S5
lmMfzb5Uui885D5qLgP0OGTqWs8q905m5nfm89LeHlLOqkMJjscimQ/pmpQlDjBU
KRX7GWxRgnGleLhewNusY41etppGvWMLsSF+wql5+hMyIFtbU02yweI9n/L8FfXO
WPqfYetxZ7Q4nSUZ1oQqqKmjk5CYVgWpS68b9Pfpd6iNhDlihUyx9w02des5kS/b
JTN0RJpOKUtgVb/iOQEqnTawbNeD1SJHrtS+WKUdA3JswGO+IqykQckD4tCknh6w
qLgNLS0TxYyhGTAnwU716yo2SdL1FkDvwdnN/gA0x4eao3NWBVOqCXp9OwIDV0r4
jI5PsiJgYhTY73nOysirzZWLzklzxCI7SS5lObALDQefKklZ9uCo59D9xySbcyLj
2Vwl4Jqk+JzQ1pu7po4dOzKp2UWkm8IjmduaqWei6LHTPioB/HC4J8T1GQHnzix+
oy0/IhFrgFbAWy+befwkguFPZW7IWTj4x1jJ9T3cvXpzh20TdZDjcnjkfOrcsxb0
H424M9c3qGFYDW+aus28z29Q53mK1SHAHRa1ZVRJZMaWpWP8ssjhE2kpbIvG1sWO
Z2X2er9XVCSLSexQoodQQDkkX7P1jY7nvugifCzIFE5AxHoRuNXAsDNrmXqKPEKq
bOy036mA4He4sZGbIawiKK8wGDtPlx8KpKt5mtZud/8oQk6zh/vvW6Z4vIYsFlPw
zs0/v3Dt38z65M73qdOPbAewHbr//J+kSi1FdgI2opKhAzncCNRVtGiABqJmi4Eq
wgt+xh0M6bIPn4SZGP+rkbbT+TzjyprFHMhXZpCsjqNYqLB3ZuVu5LAeXJ34WDLg
6yWe/EOEhsyj8QXsTh2XToemMLGTihFBygRR3U16uok4npQKNOnvm9umiix8Ocmb
88gjeuxjbbBFyJJF5/ToruW0ZY3xs+LjMYzymN4AKMe2iKWYcVQlnHoeGs1BhoGc
6KMi1Lr9G7jn72D4tPNHr6qu7HTopQS3ANAVIWXpGlejkcZfQ/O64e2zhUbR3lri
VAv/fID09abb4RMoOoa0twLTzR7MOrfBi3b7UtaEtEUhOmWvaEW1ELCZ8TJjH1Cl
wRtuRlbszAvFDrd3NP+iztlNU5bVrX0OaFCr37OeVFOU+8Vwl6OY03Bbq0qRH4uv
wn49QXvGIYQkVwSUC3pykUuwQe7Ip1TwQm/to6GLIHQ3PM0Rmz8n8ePTbbeJS6My
nwWuB3flq2DKxoBxc3p+BqgdtsQGR6zFfuVkaBBUPTKv0p/H+8ciPVMnaZfqNyLg
7PkphkwU115lpU+Rb6LdgVCtInNsqVguhCyrnJydVZ9RXVD0pCh9bNpuTT+d2bES
Q2tZZmoaOiPF62wprJm2ivgVKROx+fiug6boIUmx2rh606veV8m4Q/zR2GoNupLl
q1FJ9IdCTJEXlzYRek+0cZGAYvrpfF/rb7WfE2tDrXGkv+3m5SgmeZ02qbQ835uo
70SWLGqI5+6pWjr1hkmz2re4HYgc4dq1rh0zC5RWxFiiy6VauHT1YVLFV+QNHRqq
fTmob//Z8Xc6lieykeWaMQsWAgiJ3YlZqtF6NuwvmRK9jPeSRiqLZoADmrpzjEsz
2HH/qit5735VQNmuBbPvOvxv8UpN9xL9CGpU0ROI0jKIL8/mYwvyQa8I9sQJXmMz
6lCeP44i+mHT+hEBnw3yXUGsJMbDtIy8a0TvzlofttfMloz+W85CpVjGndMdK7UX
xzHYdgfhYK8THGR7pXL4mO/f32p/khJC1wkPCa6neOK2GrWkwLB+zRwp2zrzLY6z
YCsQ1pHWgcXkVcoYvGzFHB6GpnRABc5MiQHK64BWDdYVhLBboVa5G+ZYPCbshqf/
Y1U221KVQ3hag6soPhULPt82DQRit6p7j6YHWch6069UHYsr8qlYngHPkZC4TPgh
8W6+kAaA1HrnlPAOh9FoeEIWC/ICpeOupq6D0ISLU4UH/5fncmSLZ5oHsvY/HsJX
T9Mole0GRqhI0Az3ZnGeyRhWMjXSVA9e6zPAiEVmKfh1CycO9eNesv2OmShuf1pH
MJhIkzzqyKShKvG9WiQTvBZ/jH8ArQ7h8RR93XvCTANcscby4VPGkW6dSI1CmjUG
LY0bhpca4K9RjoWHiXSLlv4cCcwVS0bmAI+ESHO7V2UEqbP8paTrkSlvY4NIcGeU
r16NcDSomLiFm5oRfMwZOLHgcj6soo73fV3uEOnGRUVfFsTtjJd/gyGmvzR/gu/H
A4SXmUG5Qw3G7I0DcgRUlsbjlQjNPPMHxXDw3avyt3dtXS7vofG0upJOpu4YNqLV
AAWP5wd0cmcfdm+K83tK76aa5Upa7+S85FUuhScZhznoa6MSUiVGt4qCY5DsEU3I
pJnr+hgyfGZiVhMJjhis00QOzvAzY/SZ+8ToDmbjEJvCLZGY8HKV5Ry3a9N3GhSC
zNqO7EJCYs7Bxf6Sfo9pOin2yLImCOCDl7d8m6Y0Hz7l55j1UBb0E1UT1ukmt/wU
eui78GwtdQnnCw98K+1uvShpZYJWeOX9XGAypgOtSZhVggN5sG7l+YoqVMOlOaVi
fD9kWWS7f0caHvSmMTpiVPcRpeWxigrbUHB4xALhh2N4CwSyPnPgfoeAMmOjLzeK
4uz0/9tfRYTtTRuBrLhcXxIqi8Bj8nY7MH0H7K5bLlJ6KH5ar0svPS1WCVXZdlOn
WbgEBbs34zIawmiJuwymcAFCJm2bi7quL3xoTi+3/Co7cY0nm3gZmdwAzwek5Kc8
Tdq8MwU1M3ylBFnObbeKF02zHVtkW5BhP8vOq9AiD2iO6/w39p+JYPtBY27yiF7c
fcCG9XBVcMusRJ1IVeXlkeQac8IZXtDxSeJ3fZ28JcaCfAStWiheBO2YEYeaKiwV
YfDxT8VfIkHmoATf+siUAsTCd2RxdOLw99EvGifffGgYc8wAs+rU+eDZVIvlg1wU
o8BY4Y6KTKdbvVNhFHJbncp+armyXoevdkFvq1N2y7JAc9ulPGvT9w4uotNBH+0y
P1j3MAkkqgxwOY2l+lzFhemQMKIJ2tW+dbcyQ4IaOHygxVz5z81U2Fso0gA3pWES
OtplqyY/5iNNcdCqLYMn2Ixln+4mitD748v3A9sYOPN76HOao91VIL7nUEjnT3la
EIgEP8ASHFon8/wHlw680+nJriqC9NJwEx4yBi7llmQlwlQGXFH0rUuJQrVvAxCy
0yEQEul3A0vx7yFWjIQ/Sdeq7dZfQyBPH6vcoDQVJr0W2yunB9ZZPTG2Jxrdqiai
dPJ8PWwHh57S1TyXZFUXwUf6lBaNa8D3XOlxFabw3Ii29uhCm8rv1X7Z37yZbwbf
yncf0R9vLjtOo0gbpXkX5YOJhvuSiJ1Y9Ikucv7amZObEHTQpHCCK/bC7VXcgPgz
GauT9Y6lUsTzMuyzZMpdp9cBdRX9fDasdQnTiimKM7PQ123Sfwv3/Z/3y/n7Tytm
V2+pRiCty9Y7Lv6DhkZsWLPsrk0hexSNAoVMYiYaA24tHFkU+RD/5i/AnMh4Wr7D
0I0fGZyX2D3qaq6vp92O5RHem7/U6TUcKH6Sz0PCjVNRlxfIVxnEMcxim5HiIqCK
VfE1I7kda+zeyDR5wd5YbKMjxH2IAJ+bCYw2qGYdTgAPyql+lSQB7wgYjiq+e2+h
cy5MWG4p6Ssh9ON95DigeJYXn4zInJNjeDp2geLQIkCjnX3Ux6WecGgT+h9915xj
IPw++P39bZ5h0+lHyUnxgCiQnNRa9h5Tb2GCXCGiAJKlWyV7v5LgRVGpO9sCouSE
cmmvKEoSAJnXhPE8Cuh4w32WMv40s+d75RUejfq4td+NH1bZOk4ZdCE/rxPmQcKl
NLV1nnVok6qahBknZcx+uDDtu2/K2VW4yWB132e2Wn+sE8WBMgCnA3SSlg8l87lC
lXw6KfqMJ8Fzi2kRQZJxA6ua13yYHRXUq4FXrxaXiZC/oIoThI0dtbD+785mP8+y
iFBtGXPViknjcIXEfukHdSUSFAJPqTTuzRp0TI9RyMBHHc+TL1JcRgKCQzkw3E5a
HINYG6WPnpVNCQv/dSam+SKKWfp08CLb+AaTFkKuycOeqJpTzvaJt8OB98KVc1wC
SBedXJtt2cPDuXaRA/eBxPzJmmTFH0358XqBStpWsPaqWkkBZIoe8iZ1mCLzzZop
d2Hc/CmWnFBX23S71/UeJVckuKUnQ/Zid5PgCPTK9evvG3FXySzKh8lCbnYUgxqm
nTFMqrRSsaWGHSLMXbC6HTSYNdQDYs2gv0TZZW60xfuaRwfmfueod7hkQwixMpBn
RgiJ8xztYm4emLVLrXzA2DVpsEH4fCxbb0JliVtkp1vaAwm39MCVLfdy6CeyulbT
WLnp0FxVAcwFtWLZ9bwowmUAbdcmVpXOCwAv+RuhAq3sq8COjBSKwh8iqQsmrFEQ
TdPECDGmbN79BmLO9UJR2bgdZCdDqzzlHFwAHyr/0B9Cpmkj3/s+5RXygYncP0LL
EPA7MTP1Nwq8Is3I/u4B5jHbeOrQ0K0J2FoQaPImHxCSAFL4/bezhM04AB9eugyI
afKYXd7srECqwSNDMKJj874+kjQhbjFgqqX63WJhIrUGWsw+ubn4tUKrmD8ulDVz
SUqFPE7LOk3qBRbw+pHQHeGCnpbjQ+pq4tfqOdpdIFaK+H4jkisyBwTOd87o6bZV
ejS07WKNSBKJxwouoNVAdLfP7g7zMLEda/6VgWEHAihlDVmqdibmkho4AHWT9kCb
hqdEax7ztPX7gqKrZ1yYRGQbSBRa3gIcBhfIDfpjdG8V5LIKGv8NNGaw4+baO1yc
QmJtNpCcQyaFWuJkPqdsr64HQ/6PeQCLO/8sF1F2EkGGpWE1NVZmT8DeXDI/vnul
uEdaD/RdtqoN3ArNHvqPoK8HGAD+jPwlZL0AT0JOCNyS4UpD4FqbpHIAJYKopwOB
MpP3Dn1eOZaqA6F0kS+d6C3erM3pyVdvORoRPSNNoquPHHNkx1zoujJWSiq2r1nU
UGdFAZeMFthbTDEnppO5IUpsNCR93Eevnoci9xks/cBgniiByrtMYKP6UVrbltX2
OVOA2p9x1v9h0FDz3/ZIGHH5VDeDNawEBMbXvc1Tpx/jk+anGPrAC8xEtkBVGTNZ
zRM3U//Eq8Fg9+JyEty+eABu1Du58GZn3qsvW1yIdP6te3Ckk0SCliH7dWWdDyXK
bfs3f7k6kyNjGZ2qA3NAY+hkTB53KprR2l3bAneVxFXz13xZcNaKJoZobUHGfBog
Gqktm8VpKPrDz2Iw65SizrP1uHgLLrKAT7ybCipiB/6cnqUYlfc5OoBeirRRqMrT
wVSAuBtKzALVCC0Fi61QBefOvtEVr5c33m0zIcZ2R2uIhneaSIEghApH78ZUAhG2
M3ZGe8gwlCmScsjKGxrab+eStxoFW9aTpSjYemrUE7YSf0DlfbZjHjxdVryQpmWP
ZNSy2WDEkYepCSHpNl+qnPYkNQUGS7tH0CcSlTQeFNrNis/jHJcXfalldAo0x5GY
dKt1s7kcFuuc788WsMpG0hQcxJW5WRloRedjMte+np54sexquJDN1SlxvfQp5f36
n2/Jq+z4XMZ1X+NUhy5F0KXVHOSTh9vNScaYub50oOg2kUbpI+5txOf9cMuIZauR
6DUDqdloTY5TVdY7jhc/YtZ+iRjV8MO0HJ754c4UTryVY9G8lDCkowrzDvMyaKe9
2LrxftqvPasQ4njcwhiCkmoekCZ8z95ooJiA6imCaRMC4kh4p2UeKGd8jckPlu7E
ZrYiaDA4bX/hGchlxEHsrve5etXs8rv6PYzn6Z76Gipla8U/sZuS5iQm3CdHbXdI
SyeKtzS240hxmGaOfgJDmYio7rqq58sg2nmxWYrAPW3ZIvxo4R/mQBv1IruHo3re
/wM1MpfQc9Aj38ejMefDAiO4YJSm/2Z2NedtePtpmliGBlDwazc4ukFxWZRzVHsj
qhKUJTOIzDPjKFOVNBepqsEZ1yAwcRg+xec1RR1v1Paq9el0nLikaWg6oBq8HQPV
NHThbXmZhAw+uqCC6/nUUITqpjgzcI5rdyzSF0ZHZd1KRPxHnkeUcMLbijGHwEP7
fR4vKqh9MnnJJqJSRcJtEMttLs/wjwuudMnqmhK3dxbAEf2cmUXSbjX/DkQL+F/G
WWQSoCfCOtvsN6q0qGuccKAY3wGQcoPnkM/8RcAmwdDA+XdEOUxC+fleoXVY15zv
E3zXL3ox01FlJVJqfEwsrGw3sKLHGWd8FLRjbeTuLAOi5z8TQpvjeMdtTlvP4A4l
J2p8ojkp4nD+dQh7bJbSOgD54VqIwt+mo+wDjvLPPfnwgOzZY2LWInEbdQ2Z+RGE
mAHll/BnYVOiHYCa80htCVT8453p1QADhfkVKMx2bH+Gogp2pXYMuEF3NeQD5qZ8
+l1AU4cjrfihk3Kh5XSx/FEYJN75kRx6vIgQLSKD+fWvfIZArz4t+hIn14HzoEer
ARN+YlRizB4QvG+IpLvA9mul6NU+fOJZKu9z8jivrWHijthzlYciV4mOgWXK9KCY
WD3jK1Fedg492M8fUWAI8pPWjJFYJAwrcwi9AyNhvlAQoS9pFWxHEng8CPffeOa4
afZ569PGaF09WT8vvU+c7qc5co67ffGd98YYR1zltihNzuGt0WM0WY+3jMuv9Szh
7RD7lW0P/r0m+fpC9bHkbYXpyHgzejC7sw9LTRSTFTspvHtPgGSD33xxLOmQg6N1
/gNPgQuZ2fyV1+amK5aCsrionP14zunOEYdplsMa3WdQPDg0BlaoJpx7JxdQDtKC
Lsd64Yl+hAUnB3VkDXyfbFgPYEeK99J+Zz04uJE3GtTxXl5+0ePOJ+9b4yZdUBJH
1bGPXqQHQLOwTrJcdj/2vUljRdS5SvHaWsQCkA+ccKT+zUV6B4JrWPzCF7EtTb3z
evNNfcxJ70G1LBGzHFkluIMp2prHoGVBf9oF/ZN6OP8ah0hjAvmGiiJp3JQc0rva
sibCJSvNwOPIOZyh0bIB1bundDFCJb3DcxeN7TDaQZJMd1Pz4uqDjYYCXKeY4pCK
FjYpa0RkNLnYSJyfl2d0Eht5yKY8wLK60Ja8hjaCpyhJdqO7bkI3ivDmraZTc6m/
joeeYFkGgohgLvSqNe8H5scMO7YmqXoPVjc3uM8FpSZ+hEsQEz0lZlpWd6xNR0me
/NUiNdTz5IcjaxR+pZjSRpunAFbsRlkOCeslM0fZKZAtnIw775k90BRLPAGMrp/5
Jyybbh6a9cOLF/PgTePhMk+TU9Hl+WJEYbiSDAppOrTu+ywIAQNzw+fNuoVtvvqE
McYKd5ruIf/hBoUfCzeCJHgfomZyZFcJEA8KDbtExAXPjbGGY6FSetbtjdac40Rn
uo9tax8UaHCKOOOmd3P+sA2jIr5e3IisuFOdxURHn4Gme0cnGHkI3bD4QJle7anb
r8VTlp71E1vE6h5LC3uuocPQ+8CCD66t4bFPUcAIkfJN7a5r14B8T1Ha1Fz001in
bUi8g/IC17HKR8kErkeGQyw1R5NrFUHjWsNb3cPJC0L1SmpEDkIn/FE4GPzOUWVO
GbY0E/LpW7NlcF9U41zeyOmoluZA8AJPkQlMIj+R0fEEFjjIhGWVpc3Zxp/JRMGn
aje1C6bXAThT4z+7eunNH4GC4TY6+UK9LMnmHGYVZm3KMiUn3sq9fLk3++xNGg/Y
sw+itRiJqSWpDsfVa8HsmNwDMGikRZ6pZqzSY/FVImCcnt++Rpp0p5ksoi82tH4D
sJNhIYA48/Rryy4qOQnSKTJRh9gcokaTp8XBS4g8dMGZtCtk7NqZmtdTrZNAsOJ9
e15hufs8tyx7dsWKfXS8IOYK9rKnyBDSGXcaF5bF3Yx7D65gWBRoTUevtoSot+T4
pt/HV/gfUBQOppNt2rR7A5tWDxzHWcjDypxaFYGmA5Hif8hciKtnWlGhYfq1Vsib
6I2cv9Q/wvvxsIsCuGxjUhVlONOjEasGoZ/NWjcjoxpYgCIYEUjjYCUTG0kV1md2
UHr0HrKF2j0KcTINB8ey5F/XBoB5WKB1ag+meBVYeOB8ZGGi148x8Lw9tFMBahH4
TW11AS5lJupz3ce+A07pSzhLFAvX22ndTHeAFo5UkwCnjMz5wcJ/yeU5Ttf9EacT
DwZ2RPri6f2/RRw4CEutDiStF7EOcVEs4dMbLxo0qhcfJvPE42LI0tH7F2y5s+sm
m00FYGdVx9hOY5UG8CV7xT54htifvP9240zNhtnn1zbH4PHmYrDDBT9vuDfd+06y
NVihHO/AJdn+IiEF7JO5crJxs33dvJmd0K+gPc9MdD35qZDY8mcDlOVX9dIek8CC
TN3YwhSfwIvTiPOfaAWJfhZjcdZYwixugoT03jh1PduwNzrXvOxP5U1zZ79dcTQt
S7fRJHjuL9061QCXhANgpqJJ9cyE/oRwsaKQ81sqOz2qy755g3C+RgOhK751Iym3
xoML2MJA9cTfVicDdYVnJOdtyZ4XQItTSjMdZzns0UGPzAW6RCkb3zRMus8ToA+w
0lYJ7Ktwhln4AyE0fX0RKi7+zwthRvOTUtJnj59JoPqWN75h524F6Xn8rIwFBV58
tmIUAdWHCtfbfETVV02DGMisJmqjxe8a7l59oyZVlmxNRg41YyJLOiOzFWnDonM9
aoDvBUR1IuZXSvEnhTl9CD/SRSrOAH3xg9eMlXzFw/wT9q0RXuagl8+NGNS0vpzK
/KxUZVg60Fj1fCkj9+FToejOiqZWpldr/1KtD1mqqBCPOVTiXEuDBZoh6sx2KmIN
IZMIFSSEE8EVnmKAmoW9CFDforgoWCW3ix5oRAJ3q0PZKoIs29MfQSDk9E4mMBss
xPmuDDzxiGhjbGkEZ7uvTpVWpLUU5/u0zpJ0K8pouX6dTll+os85wpCTApiENsbs
0o3TB6qgzCp+9nSAWCDKxDibm8t35khSkOIq4HkwNLOxP4tUpVzmrs8NjlPWNjAT
Sd2KFF37X+L7Boo7Ua2w3+RBFp46kiiKpPG+5IEtUlpsuFkqzmGzz2kVjPxGMrYv
twrhoZJa0y7yVp0MkY1xdkuramubKnHNtt/HSvReTwwoqDmO8Ko6GhxVqfxhsnma
nPLt5NFu7lzfvDjephiGC35ZzJz89+9I39zzRy+S9r5n09Xy5xwJ7eQiHgowz+R6
7fnSLSuu7CHkQ/FGfdhWoNokHAZL1caIZdxjSzKFJLF6Okl3RP61gG+IJmYzZsWI
GNlfpV6waditf3iUWazn953KcTNepq1NUEVWx3/NeJPm7aMMs2+9kfxoihDG9GFX
JfD8suytKRdGYtPQfm3X37lsD9KveRaaOJLZKeJtq9c7jIDmJbRhMV6dr7CNX8AR
odxWiR7qt6EXojgXGXxNsv2tr/rOC4ZcVepn5UDjmHO44WBFj0I7lF4eHXgXHFQx
BCsGomGB1+B1hMXWEtM0CTWrYualciGJKkDm9VuXxF0GcWrwk3bkpMmkostid2Mu
oBOZTpu7aGPriZKazzeJ64aRbRcxT2Ts8CWZOm8JRjcwZgIxXW01TlL9IHftDQnl
VwMgusahVahlb7sJYiQ+sTBUlBoT3iGO7DTmu9u/RgbM6pdojPEafD8/4yNU2z3K
HM0eYNmrTDEY/JXUT4CbatmKWD1AUy4vEoziRyhzDzaDORxfbkHBal6zBMnwaTUx
DFKiKsupQYIcSUD+j6hostjjOpa8ruk16OdKacj1R+GQ5shvSP7S9S2ctNBxU+lq
XGw9kJWnroHKBw4W2oqztwQ6Uw44Xneehat21yLCBKHID2D9A+uohbE3YjHIpNXh
O/T9Y1K+bmGcgY5FZv7uKpoJ0r4Uc5wWDoX+tJgGOWAKa+7qcGsYWBIwO4wHHjWY
8kZFnPSghLzZQHuIxxTPzOiVDIuKcAfI+7Bk9KBOsLz0piGe1+uHfQI1QN+F5CoN
VBXrfdrZDG+sIE7BO/hDEf/i2S/H3055mcEaeXtgSjdGgHYJQ7NdBGhq2Zpy1wGN
/owukDGcBwNiOsOIhXuhjgwNnWVQuU4J6vliVtNfGwR9f8nfcTZeEGhnAJBRZ/5T
z3bxHSAe9P6+DgPjj0ErzYudt1kiy1INUhtmkRB72yVT8AJ9fZfC3E25oS/8n6E4
5IR9JrSLYoN/RcROsYecUwF6JqQqdhhkuJztPnIMgzP3Dsc5p2U3XnhMpD65X9h8
5JFhKCcEP4HHkyAp1wpSDlQpUITqx7mXqw/3cHLlZBxcKuXbdQ3RmCNX1+vW+pSt
Soiy6I/RX8wbjh/91gr3m8Q1vJHIYsfx3Ag8WgBRQfx5TPpiY5oZqhCfcGG/IkfR
NP5sJUNZ5Rr+A7Qnz39cPWtUOHDnvzRVTjeYys93DthVRcGOP2lPS4VRz8V4+9TJ
VC11wlFKMgAXw3wNT/cZj5akfS0VQbD5Gvn5RTQCIOxze6IPpN/RXLDwyELXuIwT
+KXLAvKMWOSq3ZSWFTQm9Tac6bwhM862LyEucVeue/W3s3+KL9jcrYbKX9gAuIqV
k6FsApyO4NXBl5TmQN8cxeo5dagn6/e4JMO1+Q9tPIYoejgxmVKt5u/rU2aBe3kG
sGiZs0fWjOw7U5O4WL1UM6vuAsGn4ajkXznu7VQR18sM/E9S2q7uWWBDoYQcLkRN
oQ7MqeSu8On63kwQExDIDsL8fkf6yq+ykuywnWuesORXaTvKXdCMn4cbaojQyG/A
abVyLF5kMYfIvioYunuC/DNd2SH9YMk4vOc5uLuSx2NvUpckzL+zPG2yyqfftGsn
kwt9Dtci1RlCmLBM6/TQGQOEGST6mvZ6PVa+bL17LWO/AmUswXlPg6EOXwWOkXiR
NUNXu2NF9tmhQh96A7QygifWnDPFgbleL8uBT9kyuaNw+OaIP1DVSK8krCYVeoII
9ml945UlEbUJKbUGvIWlVLJbtEEuflGJmFw4t7aFqMraSJ/cxbkIJ0ZYdGg3zzoA
m2x21tVnyVODG14qmJQVAte72JuIMpN9lvvjgHdr4O8Jl3PMlxPujI8iXzL++O9t
dX6nGjb8HGnoYvfZ5JvsNQ7AGVK8lIcqxORc2GRIaWSEprqoICvZv9Z+Brlf4VJC
leHIfWXzPnMn75p2fObfNObMk3W+ORmwqQ36dqVSW1QBP4jJiyHN4hkQhInRjs66
U3hincyf6GDf9y2gdorTwASPSsqTTNRx7YLNViguvdJ0A1ue1KGQYhe6U4CgSyHB
sQICZDoM3EB3oPMCWmD61cVb6NRb1IFUgAMUVt52E5ci5rgTSdofb/ktCiKtehXw
BJUtBy8t38D9GjLNGicgoZzROCdDopUoyb2vS6I6AnsseA21IEkYKD/7nzq71JOV
VbDg8o9Z9Xbjoy1Cw+cth9yrBh45fsnc2s6HI/xZVT44fOVmBD1wkNDSkgUBDuNP
xB2CwfNAUxZBjNvKC3+lWwyeTdS6kRnSCgFuEdlaED4PUD2MA9R1Lluvybjsv3eX
vUVU2sMnQr0x1Pbl1Dvxu33yzUD8kKUEnhHbE7Kngya/l0aiyeek4GjBGHalfDPy
5i2/97vD27B9HCMQKN4BBqFKRhZuUowuY/Y2tc2I28sl7jVh/EPNIlsg2mIxJXc1
mnS0BwoulEpZwKqfig3HAc8IVLMJjQkyzxNEjX6Lp6mjtU7XPfYfj6aSMPnIoLaz
buLSF9Vj13HOvuS0gKoyU0a9TJkJvtoz/zZ/K14B6IEHG3KRuxa8g0qayr5F4QHK
bdIP2V7Wh2trUl5FEAq7MLjd3YH557ec0BOx/WK7Ab3wyzqoUpkfEjG9Kc4Jn2p6
QPsLYgz3pXNpY9UXuxsxm4RXEedQi1VyZsV5CtyvMpb3pZj3Hl3f+XrvJ/kaijdJ
l213rUFRCINh30d2OFl5LTWupQyAhjmEVQooILQch6CKrWjADCmfqYoql/ciRa8s
o4sJ8czRSZQIWKTb7KOuNtViGvSFR2yTJLhHiYvNyy6RgyNpfmUEt4MJbSi6eBvo
CiW+ZIipBFyJ8o0pTjCn6OoNkxJLwqO5eawp8nSv9+wLIYK4FHLayXXku+wbGj4n
ky3PsWuhawlf25ZmVTFbuAxYXGPwt9N26bUk2HnaG6qxAHXgNDCghXzBieTOI6fJ
LKBMLRHnZAvXxD6znXETyvMC0Jp81maDQiDVUJ74RoR/opjXntqGAP19S7KkAsRW
0rGiuii2JNkqI1gLZNYYrQltSuz4zXlSW8ayIbpWmgd/BsWsbJ+EaUEyFMTVrEZc
eBBKFxAjw/D7MrhJ/pJHYmr/viHVw79qoH3U4gRpOtRFepHEqP+7cqaciGDqJBiM
wMCPTmqQAteDaSH9cgNYDZajvkH76+d/nOTaRdJNETvLvGH5kaN1dvIYDo9z3bmn
P0pRnd4bvcRdxk3N2AuQVJ/k4dkuYASRcq4rNkCzzlNTnRB0MjZ9LGY0ftyGZ0xd
HKVzIforyFwlnE7Ge0X1Pozn0PTSALi4UXdmHiCH+Ntj6IUnEPiMHstGIXk7xhjp
2f/IQ7WmLZsHBZY9jWcEh5QtkT91eTiIooJw//Iz3I9y9QJo25YdFmnr4gopEfL8
8AXFphDx5Bvug5AeHUAUcs3BJ1h11JVOSj4GqgMHmgiHllJIk9mILAfwZj2EHMLV
RBO3mfmNN7GMlZPU8gqz8bd6/ZQbsJjezln555s0BaNsP5gYXlyWIK+0IhZCAj8I
/sqg+br4/Ho90ixHhFaHWkL6xHLnhVpInbSskv3jDZfMiePXtS0SxNWszbLIpnos
BjpWn+aH6Md4yUUMXiwsMNjgpEUo0NvyKMWSH26Or0TqxXf23sNCHiPrQPkTr6Bs
EyxzHvpTSE30AMz9MGdBemLhUkjBpYfKqFvDjjQbIpWUg0qKVciOHIps9zOvHsGj
JHh+LAoH/wSpmTnV+skPDFRJZhg+WE25Jsc8tgSz2idBLGWXYtz1+KAeyruFPm4a
bvZKgw5q73Hrvu4pJpubdugTdDtzNkQ92VvNDavtkgRko1yVRfT+IYjxdGLNN1Oi
y8FNG0O5d5AaxNPQ2wQ9jSrzW/4/1FQ8uU2NGPZFxA+1iPOkpIf5fn+rd7HE0A/M
vThyd0ailXdZEZURVdzuTLrEu9Yy2BXEkof4QfmK0NMq1+keCgvxjizh24zkfFpd
TMgD7HvodHyoq+Ryxonb/TnzPe6xFbWBJt9I0JTMJ6rSyKjxNUA2KlV0qCEdVIaB
+Jfge21qHRKEPo/H8pGndSQQsLCCjzRL7uTmrq3vT+3bSC+Z6hqjmMyCHfTnwjzU
kgEvkOrYvnbUtfNf5oJS7K1y7zygkapHacm8hg0u/5p+1Hr8sM+Y/gJZUNtoJ1KV
5NDVzSnuSjFtzFkrCSj9W4wyEGf7+RxzJiEqj+QppIQJKNtyo7Jm7i/bFQFwUV4l
Qeek83L/7vU/LrCA77fMEhEr+ATJ3plB59BwwBKiuyAHq+BOg2n8Djj1bgNP6RA2
5vezs17rLt3kIG9rC2F54lMB26ild6M8j+PJQt2HGbWAbuR5pxbJYDf+bQwO58JI
Hl7xd2l12zX7lsLHx7wAiaHJOkHfQK8sRpIQK34f4nhPVmf+mH777IVpXqz3iTVp
lPJoZRFXKCy+p3m+sAk1v8+u4gELQoXxL8N7vzbY01YTQRdIcYHkVxObrbvAgJHP
uCVKPvsSi5v0uTvz647mBUlIKhbvIpzXLSMjUsCL5HSu2MUkFcpENctWaQRAouzO
DMeHruskSdGNugcSa7sIblRLYhbexqUlpXGZsH5Cwoz72+ehjgsIXV7lUE/ZYx5Z
a9kK+eKhjkjrhepakclYP3peQah5w3KVU+kAXR/tRGrn3Arb/hrHspmrH0YB917I
JxTqkMSp3lF2Zjoi0jktnwJi0sqYbvA31o6TWjynmg/lnVnydNQ8tKcUiixknMae
crITBdYvYydhwBJUwOLZPxgEVoZTksrPGsB79t2nkMQjoSuJEFq9mliOO/CcWYud
MzwKZIDLiqEGns4EpHT65P2udN34NEgDCl0Bvb7NYVR+NK4sYImz1VKxDD7WY8kD
M2E/NhZrWXUKXwnKnDI/OEkfZbf0dGBlac7YuOmNspE+Gfe7fL60tinzQiSoD3fH
Sa1AtP1/s1kSWvA3IOs1skphhWVinuQWrd5LGcAZN8mfLFSkduQSuZtbElEilNhK
4ubdHbgcDw6mB61f4kSTXrGufdv3fwO429LGmQa7zefGESE9Z0VQKw66yeNlnNmS
5hILVp9AKunCFaHGJBYdgl2cLyVHBDT7JnuJeyyrTX/aMyYmlP0n/F4oCo6gdnh4
oWGuggnOgWRYqhIpZIbgnIroS0CFbYQAIrH4UUWXmW/Ci6lc7kYfDcee2kmCLNpl
6DIWPPd9RKw/W84qkrvupfkpo5drbG+IaI6nijKUrSyG7U413fwJjHjxF/1BK8rY
F4/6CSC7MNAQTn6lUaSs9RIMiUO1y4eLxNYdMNKKmu7V//B0MZelyW3DwCHdkP/S
ju2I8qTWdGyxGPoBFB0bU+O12P5N4u8XI5notP6nSnDcrhGvGBFmrpnAwMWUlvte
bLDr5yJFLMMCVCTu9g+rZx8VCsqQ5d0wgbJFp2ULF7hhLEzwxaxICby+++77WTMr
EZNYUocl5sDooSUe8vL6XEx+rYStTEWsgzVJjURmU0FUQkdPM/3CtqLLR9YJeQBi
cNJij0SBNZ1HgwrG43T8Y0/USSmLjontcsA/ZkGeoB71iwy8Z2QEhQ0vR/VsWxwG
l0F4k7oPCrYvZMh8RM2t/bIv1Xh4/sWzC453aC1jEbkzek+R3B1eRmfnX8YjwcsV
/GyaCD8KrYfRoopARC2wXsfCuvkPpXMmo4C3/qdKRg1kbUjiE2TXtbIw6tmTQ/Z7
lzVrD453EV1hMLCTyw/pI5q1F/1I1e6zKJppXtoMKJLGVJfdeedEDmR587VycRp8
A/7WDZa5pgGHnv0H4YdWuYaXFtEHgymMvuESAF0igrk7VFuqfVNeupePR80jj8MA
BsgdEGAygqz5lbx/DnWGMCM9x2TdAONEF2/Yx8QHyGWDf+oXs1qaazWush/rX0Wq
S7b/htsKbRuB6zg3rLbOSaOnkfQlW1kP6PRZOrXSUoq+0A18M7g83NLiRQS9ru6y
HZxUAxrkhzsDK9XwtkirgSq18ROn6a9vNcY8JwkiMen436GUrO0nKlfhnt6NGL+v
TLGn43lybVrqw9JtRSYx6AXTG6/4A/7sLDWJoTl30xzs6olzlzcOc2c4GPmXspSu
3ueuQPXVmv/itqYQD2qQFITk2i0XKKoq3aHIM5yfs7fAlNXwsEifaYoJ4jIHo7R2
nQ7XSBmfQaqrXDotJmm/K6VN9nn6BL3qdE9fy4Qo0e2QW6v5uiu5cctjuwk7cQ5h
ncy2TR9G319g6xmeM/7wVU+lE0Sn/hjfIzViBkdyqZ6fFPDTlhaxR06aXxEmHAqS
qhB+9hPeqEEWlrytJQMhkw9J6cqB5idfwnho2FoWgmnMiCQwBZq/ZhtDLp3kxHcQ
Vh5tW62Ly/sK6+XUM20aTjZa3e/goS0MPSNKSyir+cYRbHXuBtdE1NEUqxjffhrD
yJGrPBqz1ITmwq2S7A27jNbaQJLhBK1kpOcO0eprZsfjBsL/xVTiNbM9Lrllm1m8
Qe64mLJmypMskx3+5yFmas7TUYopEDi6tvGvJuHeaivwwjLO1m54uqCDRQXRd6oo
lPLcfXLbPzk0d36i5pHx47XGlrvXcvbjmxeRhdPqY+SH+vuRe5kAX719cNKu8sSC
+xEsv9spVHabgA7XDqNX4lxjCTlycbJQQ9iIpJvXGDEVaYis/CBhvX5v+tq6X5f3
MST98/q+1e3UGpOznOZGWhWQfb4NgTNpj3HGw6y6WG/t255ODXx6Twf3QbqudDWo
RG7/Dcx+wQ0Nv1Bs3AEmZnMc3pNMwDBQyFr2/rcXYFReXrrKmLsVOoRI/EADcDmb
9RVg+UrAUtJuZKa80XwBIZyY46uQ5jHdJ7JkcJ0K4xHcdqloNphHTIctS6xHWsMc
ogotLjWWqgYI+IuGBqWPRCjW0AiDKaYtN+ogXag80Rc30Gzo1EYDLrQbfFU3ijEn
+wdoe2Y2zAwvRnhVXC8UjaWpEyLGS+RCqYI1YNcPIYLYXBRnSVGh8RAhJqHUDJY8
cdYdK7FuMnrh3od3ch+gui7vdFMkCzhoB8e0EkBYyOrIFJ81tParaAQyNthhLJEd
BMNarkElo67pYHFXatFZEdcw5cPiNmgeY4fQSyfkjHgD90Yb8F9ujuP5rkiPE/Z7
3Ndz1dNY2nPd7TZSFwuJ33oeFBuCMSUqZKmw0woW52AX5VgjdDWqAdfUPwYJKeTB
kXpwtJUBaCNIH76SKXRXmclpb+nEZlLDoALRCdVP++xod0J9KMkvU7TeKfXM2ZeF
zz1nj2Js0PrlumUh1RwjzIeXblzwcI++BYYKYYbn35YrsjVTaSQ1MlD534O6Lspn
RLKAu1Fm7K2h0IPhZ0ZEf66Gl8vIKn7/zybfJbMMg0SshjypaKGCyBPhy0VTbzP1
LZ2vCAE4QUhSKZcM39t0NI0NO0n5DurLHEKI4fQd6OMU/ZT3ObxROAHuvMwC8D/W
5nXbUYkR5PMq58pmmWvlid/4y4pebkc1uz4EcsspXEBJFEUxzRNAXzZvOf2nbpfY
Rm36XaShbT9GzoOqjeDa9mW/nKhf45GFmRoVpCD01BY+0qnttCLJmvflMKhtoikz
RK10zal/XlwLs+LD1NFBnUV7sMrj99if3x1NzgTY/ayVGLMZnWfJxWy9R9lVwovO
TeMDI7km8Nm0iZR7OMhmxtDjAh6kZnDBCH57iRNNyf5LpFlZsZlIx6+/DYgDO14Q
WK/vfzOpSigwRxfZlxmem5VQ9QdicfBPhBNKCimaN386gwnckbh0YqRkc25fPks9
C+leeVDTN/LIvu8y5u9WbJRei/8tIytCwz6/xEyohrj9EIWzkDu9KURiqoT4B6Lr
f2Uy1QMAGfJQ6j3ErUwAgxCLK6M1TvtA3lRkSCVPZ1nZg03SEsksWLCix8oJM/VK
IWvHIwqYGB9fiJx6IuQ4OQQBEwEhTI3ftZt5H0SoC/Mau27XTu9KzbTBycE5rfu9
PkIwqhWisZg0AMz/0pAUb+3Q+RmqTg7lJ+EMbNLBBcAVXS+6sQnL1WFCAc6/LDjJ
8IsUpv6QnNmJi3gPKyF6PKaEHSNb2OiruOjCPEb4BjSE9sjIaycB+z22EFmHUdT+
yhFgJLOaRdDSqrdrwGqltmGB7T3tskdn70E5JtRhYI6IoQwVpH2YeVg4sOWRCOQZ
uZFEAu/jsBGFNtx7DI1hkQq4k6DS7J6GXqXFDiwGcOK7jT/bnrMdgR/hklIKQ/Oa
woTLNUAnhsf00dfKjiMm0x2+BInpnlTIf/UAb/miZpntFGENFbZDDYHyqN06PADz
uBkgra+QB7U4bsy5IHvAUJuAoC7VyJuVtxENDLT3aqKuue9Ql5BeQ2zYhSum9Qu1
BT1YQJ/RAnzpu+JJY5ohfRsVEiGlPCNXOkOFRFxGAmqdC+WOeAdTMX+3Sd9+0viz
vGhhXuRd7hU5IG6e1X4SYhxKD2iaRWyMRsGgCuER8cV5Hw/FLk2QtSVzwVfAZD3v
PCXbO2Aph5B6FIfR4ghtIqBTr6bqNs3C7PsBIF8BowG0flNrLhOTX9fPY7QHDEQp
f7HAucBjcsjLGn7EQXFW464KUoDJmPM3XISYTomf3U0u/Epa/ikwA9TI5DjRFlYp
LOaCqCOL2znYvLbXV4eUmavD/Za/fsaBYgoJ0u/aENLRttDAULRRM8735g/zGnze
cfPkXt4i4gCIz7M49YF7CeAm5IFqPeeFKiLlPUTXNZtWnWXgqfRHRZRKaN2z7G7Q
dbi9GYC8fQxr1K1N25COJ0007sEySjwyqOu5C3ccN9H8+AkupUMjC73PqZvOIpmI
U4UO2xfa87+qLGrB+kuK/vMUsUhVEygnnuSOPYGMiuEeIJMZSXjmduh0LQcTIjc0
wyhokU34iyMujo9KyaHI6X4vPTJhq5Oq+oUcSKKbS7jZ0KSEQXawOHW+P/iRNvGS
7sQ6p4SyKmvNvrB8wK5uvtFHAtki8y3kVXtJ3j372h9o1/kwM91IvNe1l114Zmea
HpxpwyDyAxyEBF5f9OI1coJA0mMvoLSjScN6yLgHy0uv0vLi00rL+Y86HrcjYrpa
7WB9EY3wODZGTHR4NXABG/rNF9opqvVOTjiKLIr4PtfjY0eCHR4DqtZ+z/sQvpN6
3igMHKRYM4yg1vwuQm5TH1WriKjoAcQcsQdt4AQkVWwSsJNHm1wreVb6fiKoWoVv
qZ5Qa5chj8XKHkVf771D/zWqpV2R6tet8tZbbJwHwC8nIKXTdVZKZnmorENar1Uo
XTd3bT3cxQ1NpSxVLHUdE2KZDvwouDAimKu5Xvd6dGQ0ipv07nr9oH/MHCQu05Rk
3ggyxMDwfgYVMGpt3SckH59vvRoxPyoHia0W3/B1Za55WszuVLCol2W6H0xyCxK5
yBL+38CN+ooYc1Gvsuv8DzRn3AF6LZcrzqeusiMMWPYsTJU/7z5Jj4QWPz5pf1GZ
6GRzpUcqag5PTlHWo8ZdFQw9suWwPAsIZNPzLsOY724e/OqUHmL36uFrrz2KXy34
WYCOJV7KRVYR+9bOCPUqC1t30EyeVYh3qpKjK5eEN1lf5i7cTukO97OJjwXhUM7O
eZlS8JK1moghvtizLyQYP84q482rlfCsY4WhbaWwxzWV7ZQURL/Zz2bKRtJiMxoZ
pIkvGd88qOmSr0j4fkzydsHAUMACZ5sKBvBoZV/QxjK3rPMXvffjD8vPgMB/5Yv9
/yBcVjNMrz2UwEzcdPn0ByrRCYDCpDw9z0ptuqIDCn7/BVn4fq0cgt/X+byQhCIX
+0yiOfHmohWxZ4XdR2BbXppKpzmEWwh3kqYmjzbaax7GtqSIn3ra1lffsTpHvWcO
yrHOThAXVMwyFUp4CBCIGKJSfi8WhsJuqiePsZhWxqIQFDW+CGoQ8pWsSFL3FGrH
tpzkrhFDDiuISTeU1W1dc8HToL9BQwOOB5fY+xp6F1WTFg/cZy29TLeObgbyVHn0
oMCZ9KmXY/vNsSlT3j9gWzQRquBuH/PBUs5Bm0ZAdREc+zlO9zv+sWoXjplzw11S
vv59iWHiw3VVQorneOGPG9BNdQAKHYxanu5AoTXIRQLODgmF8Qj7v31i/OgyadDw
CO5wcZlj/reUen4/I5ZG4staJrApLbPBnkTWJtZLacec3rDu/Q0PhJIEHVrHse/k
hBfSqqcg5VJ7ySq6Q1duZq+wuioaRj1xhPPbrBbn6xpSG472lEEkE3vDetsAoT2Z
N8W6StBdvScQ9mboQMi9cHM9Mvy56FC5GEMxcV7wFIy6EApKEWv7UTZHKDrSlV8y
jYXTZAEOKRQcslhKey02OEgRhzewjOkMuPVw0HSRxP/25qtneeK6fWZyMLAVU8y9
gyZyc68/vQMuEvadC9kQ5qmQ5YqkjW0a/aKyQuKkNme3fGEnIka6XeLyEKVp9QI2
PzUQVz55Qn7rxfKEae7pEQrrPNqUOM+YnY6EkjVXPeJk2QiCYhPFkCgSxT4O8MsF
2Yyc3qYazaZtNIQIBJ9rsfrs6/VKtR36qxGAMTrxaLzqXlCNXYRFJHG8762cinzi
jhnkmRFPMhE1SHm4tKDCCc87C1JsJc5M98AmgyPiBJDh3P7oDxaBeSxXW3R98N3b
gc3oloQbyLegOK3qEkrf3WqzQmHeipmuYeWxdVZTPDCFkI5OXBey2XMSk5Co7YQ4
rQIhcI91db+RIk66L/OQC3fsSbcR+8T/Yqx+1ZmY7NBFQXoq7xRj6/KSxYX4ZPLX
eviol2RlO1N09ZSoNmsI03a1ZL6bnHDcJoef+RMTmRgP+28VIYB3+2s635mlDRwO
Z4fUblo2Mif8URadTyxY3xUHpomvW/gzuZDxHfaM51FCktHq0lcedwAAb2/OmoHU
0YDGqLBnEwXmBPSoNawOq4HoQMsj4V2CJ9H01YC5+ZczCW3Tk9gm6GabSoG9YpC3
9qEqANqC4i1Y1idtoZbN+hOXc4yOAjl9HengZtlpuoudr62ujMNcgJuGYuqAwMhF
ailG04Nk0sCOhDRLrYOWY0h/YYA2g98pNIsp1VP0aac6ndjBMLcKoZ7+K4kOm8y5
mIFXRhOfSzWN9K375kgl0kfP0MrMzVl/bfCAUOuP6llAOoJ/qUW/l7htRoiDsjhA
a/mJgsFcxIDTNkYnmXtKyZmK2sBWH3PzRitZpdEI9z1AT8xH4JnLRWNDHOCBs5+E
0z9pAkcZfMK9FWTBwJN6/sNLldEaaFlS65D2ZeiEFFqh41xPEkgkKEMeYUEhwgg7
hktAIU47fqViWpKtJ5bRhl0k+i5p8wf3XhSGV5n8kqsw+r2ICG4+Z6EQZMdnw8tf
tr2xvvvFMXPlIFEgj46TVgJP8BlpueVkBdckOJEqYJf/6t2Kzh8FmKNQMR11hlCV
xCZGkpzjqBGLdm8UNr0BL58tTcTrp6HTcKwd76gPfasoRn35xQ1jNuuuNhBFGOyB
tDOxSgyIxHHz+YGsZHsicJmO7shim7H0V8VcY9kS6w1dxyWbTRF/MoZhJ0cD4e1c
trr1+UrXGEiewwjjx7JMpLpyXlNtKB6L/7NL0eAKzLUrmmNr2gmDo9c7/fh4PMbT
H4+P6N9n0RRuG4qRV/sz5I5dknlbQhYcV+L4BK0YtLSPe0IR/2bMfP13Wb55iiqD
H5lG2ZnGEHaYsJJa4IDDZ7Su0FOgAkA9qNOtt2KZME1188fdl/qZMHlxWhpXBOKd
MiAy5OX9UsKUQhcgZ2P41PyMDxHn0j666tIGMe9ohj962fErc2CHd9+Z4lSzezr1
rRiZI9cQIdcDhbVZzZpC+NIxyY+fpbjABSmKRShBI5O/31h3pSfbkJBANsQP09Xd
MsD5N96b0Ab6waAFWedbWKNexI/nDxofoZVSshKc/OwODdJCapSv7sKk6cKLObOE
FgrRFjejftO6dYRf1md7m5bM0mHk41hPc17SUNrN5LxmRqoHWfQuoq94lwfBa2eb
H8CoetKylB45hrH9NUn/DqYXnES8t7Vunr+MQhGlpimCDqKwpayjkiaFuR1LaJrw
5qetFz8hEYV++zk1jrlD7peeBz1FUCbJ2hFksR75+efiXeCkja9Qy94A0nsbhjbb
2pocUSZ7PKJSXvxCv1jz86eq6TwLLPO0hUnqyYfd72jVaMMXTp1prPPr41Accw97
iRPp9yr2tmQINAa1OwtI0NJl3oV6iHTGaV6ndNdZQT6BVLpNwISyZQ/aWdpr9r+H
cNa02RMTbaxge4aP47MtZfCV2pKu9CNO/zYglm0+QJIDHK846hS6fT+h2BbnEI3i
9+Zk0R5WE4s/EL75JhK8Oa1TZ7X0uLcXwAfL/UaWcxL5sNqUdSFQrJvXnb+yTVt7
LI+4nVyFXhcJ89FaWXi4C52CHT04+9mlDe3ru1ellEsZhaviARJSz4H8WWpkeiKY
W2TDRIriIZP4TmkvBcGE3RvPCpV5nkQXeLSIzRzHqeUa1rswv1P/rcmvJRND3DKI
7pattj/eqNQMEP7b3lyxX3Oa8BVLkDRmBW1LE4WCheJsjpD+91iPHkVhZorxRTl+
ppUwzflZLSVDfOOuGvadrwXWCPKjxmM0ebCOl/Xt4/HfpwYN2UhEI+QujBxx/2A0
H2d5O+J0A6xfUwbHyi9gpDUP+KjmuR8YLm/b53zqww5kaet6jm/20C12AgYDliJP
AOx2FYyeIcBXY2JxJALv5AMYMv3po1odk/XihTnDgfqIQHGGvOaO5rfGCg97kkCw
P/lvYCx7riIbLLydI9aqfoIcBLyfqwDdjix67wj0/hBvjLdpJqfpy28Jbvl/Do1C
PqPLJ0lJQDNtiw+Q+WUP/U24CTp9L8uUPG1ffksHnj2wEYRMQZN2GFxLYusWnQ17
BkFBYuKxv4qOC5FNTHzph+PrFmWPRBaLZ5BhRWa0K3CNn/H9lTPy/QxTr9QdPcb+
rd4EebxM0lVSwyWpJ0Y2t1HV6EV0SZj/xUG1y2iPpVSzm09HwoWRVYOBwWtKY7oF
0kWNY6n89GPPnfRtEj01Bzp76PwwkoJtSZ7758uXvuIkGY0nqhGjQ5OlGwtfs8P9
kkyb5/rLIAbwWPADLZYFCIOxYzag5sOoE4sQq+CREse2eOKL6dSX71TbkcMEeCyN
7uBWvKP5y0erM2JsSJbtEFXLct1aKWLEd/r6kU4IEYBb4fXMOc3XqH5dDTJ2l5yL
h+9HjUwjrTywZV/jUf9AD+lHmP1XLrkqM5uehA0w7KNbqtwEc1OEuTH5TXGi4GoB
zb3TXq3GBwO6Pe8zNCpkbEexts2G4csGEKWjqmNyfodALnxUbMleI5gmQ2WGnPFZ
T6IDXpyWlT/vIgvpalgUiau7c2dLZ+Z/mBy6bnuEhX6yxbOdfQb+knnJYVMPp743
x9zgy8CTaGgS/cPLXoZ/1QtI11aOCwPk653b3ZSz85CnqqIEsS0IS29twEpp1lyb
wrxomoxB7NR6cXD/1LrU386nXTBkbrKxUlMVMOHTzf3wikxl6D7OqiBncuuT4aJd
OFf8Y28dAq3GATXaT3/2/ZOk8OouyG3y5acCeB7N6cTM8ETRspgzZm/5Ptk0AbFo
miXBQrBEH0oWMf65O0KwpwmErQsZAEPBbItfoH+8VmAfTu16o2m8IQ37w/x1giFL
kRJ9q0zuvbpJCp20UjE8x0N07bXQDple2LgLp1IJk91cJ6VzTykwSGmcqcICDBJB
5Uw4HUD0hFFFdqNzOi/biT/UV0YLO+KEtBJY1/RMyE2v8aMkChTeHGQu5mMdVint
yOpRBKnJFlOddY8Cd3UicyTUk2EvcfNXMd4ivfsNjCQTe5TRCGEkY8UaS+grCZxw
JX7gMuiUWcMgbbwiX7X3JMljLZPCWXWOVa8OTCg3bMK1F0ckVnMBKhenXR0rjv+N
FzfTmqHbxgDGpFK+NQA9dKK71zTbZtUbpToZmshV9rSbBFSmsNJ8s8Taawx4TjGv
xb51riGrlgYgtADGrc8NXMrCiILIgZ3SSqlI1OoGiUGM9tyW8bRcEprlzkJ9LFHr
ywXfio3KEPbOSRUOFZyNqgkiikJIRABxPzEkRKJDFq9dIUWAmhjfw/UrONrLRdq7
OSSt/9sH2/4W3AUpAPySIPrEOXZAXZWQW+9yBp3mGtGAD8qgEfxJkxXgcttSmYtZ
j24nmJP0qh6hE3Ow6vNmwBtMGkErYK+vJqpNPu6PWGTBgeFFbemQCUc4rUNRujJf
4mO+meuL8bSVhtMvHqgo7edrBJGQgDrnLiXBv0eD6jqqu/CFApKpvnVtwqQ/u4WF
NqPZ6/FX6km0Z5TecDpX5KkTkS3yOuHuZZSHmC0ydWmmAVwjfZrYU4fVGzfNFIff
gtiutacJaPIZTMwlfoF/5DSVQCpnOmyf+VvOOATTJecYfketASEflqM1RoNuzk38
BThiut2UKdjJxo3BiDTvDPwoaP8fV6E0ZCbm/L7Bf9b+L1RjPiIXhlit20fYVOA9
1AQKEQtN7DOSPK+1jlppMwnq/TtTwdaCMngFZV3D/hHZdhGeIJ7IZuniIlna9FWk
n3YaQBVtGCgG/xarzHDGK/F7PShsVmGtWbHwByccpdBEVLGgQ3s7ilJxhkiINgaa
3yoGMiLMFun1qMmhl88V0F4JtNmh+AUkHY/j684dVs+y68Hizi3oMjvlWxB1hTbo
SoqyMd+vWWkpFrAFZ+TAlDb2ts2zgXBzIHR7roq9GckKK5DoR64imKeGNUq2sG3X
j9nnUcNXC8D3UtBdUvZCOhKDX1jdzqQk0Apkdr6W4Pcqa8Rb4VRTna57+iru0gkl
wc+42vwc7+2NjElMxiMevCAMMiCuCOps8FdWR6yktSNCTiZl7xOUPzyefDHNR3h1
IeqJbm0V7ljV1OyLxncjnx6aRyyOrrGoplqj9S0WKdmQKxjAhSB8MIFsutk+xMG9
AisMbLKCmyfdhtZEDxV/fWEx8d1wGb2tiw1Ejj1gfqiLn9TzXdBt55Rfa4j5quun
g0tHX/zOYFhQ2FnILHd0RbnN0NaY71PCV6wlQmDddmseXDW4bp6nojW3NEOx/p/9
XJ02gnQC3Dabv5HC8EJ00umd3Qwo6gw4UYH+X6YDn5mLwK9kZ8g/vGdrCWeLdBob
NG4EhBush4LK7Yg0yQiZGgsaj1p7A/Vc4vVBYzI1U1uBlfqXvoj3e2W+5N1KzuuI
rpPDn61DMduITZm4xMvzEXDFIuU02nL/XNRCqN/iXVDkMb9Mj3zeg49kZauXpUhz
8/C5x6opOHXvF0ockPrt/B9KgkUNp2vVJPIEjv12y/M8i+EtN1pk8AF08i1JyxCz
ybdrGJJ8d620YVERu+hZ0DBlnffR9dbFGHA8AeROKt3c7v+hxLuIOrN6bWGqZpEp
xy+siK9JeqezMTOaTeGA0KWMdPw3ja5zIhNN5305Ph/LIz9bTI1oxKLRyUU8p2bx
zoz1iu9Xxicvn3gNZu6x3SaALqs0Q7RvwwUOU3phZB1RPhzCkvd9AhVFbvMTOK6I
VYE7Vcd3lLR3qmnBTxfcoWWJ2lK4ZQbHiX/iFOopx2wwsS5Qk+fWswCK6yS6YpT7
ezw5gidiUWcltSExq/YqfKAKjBGx4OGuW95XG6bl5DFolSMXbDlWFtOLfxJM1wuR
UkGre8gpb/0fldg7HnnV1GbjH85uoxPgzP9Aj9yUElV40Zbw9NlyM7pavAKiCrw3
wsB1pdPZwD6oMt+zG9Djm3EPbSi7g3AdrQWRRjmgLS7hVZuqiYbuWJcOArsbNxfC
EWwXWta3odX8uj4ADAwll/Ae72+UC4YQGRyP8U/+9cqxmbUyj51/UEBaWRgZKhp/
T2fyxApHUZokfedtSyguLsp8LEp52SZIUGUMtkh2k5QxnzPgJY6Pm/SQz2USoniu
krzVoSV+BT1VahyrceqyFn5+hj8Kq2ZwM/GxO1bPjlcAOCPQsdxf4r4DumxlQmk8
nhfXo/Pa6nipWAKna0eRkdAom1+QzjrJLWfB8IAYXbHgFVXhOAqnD8VHs+miUhon
p5WVy7EK0Jsf3FrrENXySnYR6YCH20TDZCsKTikooGF18Cl45MjP/iR16b3ZwLdP
JwHNpoyyIYm0lzXZRWc7YfHvedblji41J5REXUNEfGczcCwBMfTnwOBAUM2T8b66
5LRgwzXME6FvrTUvP5ehbwgocka+7MxrdqJ6caiIaSCTpYG+gW/JTzZq+U9JbvD5
42WNdHETSFDdCy6O5qxaTKeGpjk2RtyL+G0LNjAxlAsjOpViwzeahxNYImooy7kB
6c4V/vWXXEpue3Gy9JvSAKKjHQl7ggwp7lULz5B7MmBbYa1O+N7wo8TY/HIxY1tg
CqnetkEYCod9L5qZTgVeLklY86SeOYVXPFyNKyeKAO7Zvq0//rZEoKW6n/2LZrMK
aZDigct3RMbeAwjiFjgEtHR3XY/eJOKMyEanW54bcOfpPaQTuZWStJZBlNhtU4LY
1VQSAcpN+evS0DZ8KWR2/zbHw5nhVv/c/mqq+0zMu33VFzBK11GZQksgzwnMMKZN
sM2jnZF1hzs8IME3xbwscqztM8jjHW1Gsqt/mgLyzKkoXNzTW5Ff0QlqGKwYIy29
SCl/CH2PB+lbdB8QiafOFyZEdkClyW0gCzvXUCEgIjo5Gu/swIh9y663mNIxUZjC
dNr+2qgoSc/ztR4rd7ip471pAWtUeyLiSKwnb+BQsty3vfO5J19sojyA34EMu7mK
riL89pxCjchaXzYFraksjp5osz99B61L1Nn4HpkkLs9M+0zskBn7ViNDa7SSd9Xy
vGtj8NqtfpSXUGfJqHAjEknap62PjGgy72kRm3INcp3cYnYMurLD4KDAZtQDkF7w
QrtN4vfDtsSJWbhcjZqpZa05vusSNv0GIlG6eNPizsvmZNi70F0bnD2fdoH+qsbN
Aqkwt7FU5haI5qWd4AEKDnB/XXFGxN2gnmEwM0irlJHEbTBM5MpR8zQOt2OfuMCO
K32gIsZYnxS0fTPvESHiEjllFXbuLMv/GZUjdyES6GW2JT7tLqX49rMTkha1eo1A
cqq3NZApqfcrv7O8HjmJJiEV8XTr8oAZUe7Bf1ImIT8Z3kobjcGYDF3VmLPtIdc7
ST7buPydx//YVGc2r683GEkmjadVDSAmrstbyEwCJVY4z5ArhvjKR+agHbL7q5Pc
QWVkZI533bcROBKpgiC+LJkL2gCCPbeaDZ7N+/qsOdMlMz9Dl06+rJsXmGj0ZrmE
Fmx+qbhXeanSOq6TfW/7ctqE2RpC43QeVLTXqBJDN2iVlBQZuQ0b25mUXstZOj2e
wiUDNYqtv0fDOKNKw8IsUcw0GlvOskxRLVwfwKCiHg5tonvPlm0pOmewyMTLLSfV
rOmoEE1k6hB9wQ8qZfA/+keGmVehaaEVy53oMgiDwvkOwRGbc31FfSe58aH5vAsi
OaxGn64jiZJSxFQKbKA2Rd5IPf/vAZGqiyDgIGSQEYmeLCc4CpZcwEBB6NYkbvCd
8w5vYN+xhi+SZBbfgAqn6uPdlu0xl20d6kZfb9V/mF/4FwOC+JyxM/ATq1PFQkkO
uCZ0/h0P8zw2aDbL90cvf6FuN9FvKyVzOJabiFax80DvkMKiD4ijLhW3hzwvwcne
6swDmareGpvGSAqSuNHCBNtErHd1GTwlFjJ13nkoPPo3VHsRck8E/uXKChvaaJRL
tii8qupcjToro1ez8EdT9+2TE1ZZMMtT9LqrKEWLHfCIZs2tfdWSYlralqzr/gUO
Z2FGPXNH+ng9OG6k4hhwFUpVYzSiKCpQkFSLfagc6zhUOXDyNfFvdw5JlW9ZRlNP
2OvQu+P1R38ZpScUDgaQXwFySbuhvym2g6HwHRKiUmlEK9tEWdvkJsKTCZLADjL+
3jkbOEOTuHNhIYxHdu7Yl99iFgPRYxw6Oc/DXfHZd/Dry1jS6NbvX341qQVbl0hd
ELxZ818QbImzi1cUBjosuSj32m41YlaEj31eTu2q9+fDblprkA6CFIsAjxoddfCs
OUg/exGsK4nXFdMpCh1gWwo3CqsUAkySoHcISFRf2kxRZqKurGsGfTFMTFdWr+l6
3QBNmwmLVMDPCphAuPhkECNLfftg8r00T/rR/jYZP89dlKVmtHmAjFhqeiCtgsnK
W+XvFOHt2Mc16imX5PADGNXTC2vOSnqCt5gcbo6ql2h3xajYnYr591U5lfIydBWL
89HBkH56EHAnOHpXe9VdwVjLJAdOGuKOhZUdwm8OVZa8G72Lf6iht3TH9QSEmAj1
qgD+zkx2pnI4W6px6/7siEFZUCVs5knBYmSogWe6P2ITHyNScp1PyL53viW12T0f
x4qyjJfkljMwOAlzkOHvFTFqCYAWdqT0zkLy68No0JQoZZqeluZVSQeKf+GVgxWp
JHGqFkQRf117Y0UtDm5WkWEmGGzyJRBJBSWjhRTdqsN+iljTJ/trvtqPdELRE0Fk
fS4uW2x3p3cZrc8DOov0YoUeX/eeX0DJbLR1IVs5GeRswAt672mA/H4zIXT3fzkF
54RSNhg+ojPH1SvFeZghGWbZaoWMzvt3ntFjKvHtvPDV3SrGupIqzJb6Zlpon3ml
dytClGw43pQosJRo1PTDAUftCv2exQnlrAJe9c2tdpVVIrsaXPUy5m3u0A9ftLjX
rn6WqFIMPOBIqJHlPuLRhqF2PcjqpWXgl+6GrUHBreF3EkkFtNaDiq9YzVOA+QP0
ZisDjksYlHnXT/fXTJsueLnZ/MGkkIBooCrdXendPHGN9MCjXOqWr3U4xMIPoJhc
2hSvEykezssIaPUVl92DqfuWSvikBUZWyH4j4k2xLMgBl8Bj6sBRPb71ZFSy48M7
aoR3JNu10x1K6wCsFvr4Zq9eC1/pUv+F6Khd+JoFyp3h3vJs7rGAcHhy14+VvQOj
MKHEa4J4jfk71HMjr00uMB5nI3uSXtuZN9Cj7msOAR6CkxT7T5AbJ2k5osHkGq6e
SEX9VAgyvg94fP7e9yUILbSWeNJUT+iv09GDI1WXjVdzKvkjBWfqG3gCpStCfD/Y
E5bR0qV4osIDXE5491OBcfiD82epOdNPqOMiTdSlmibK9G/uuHJaKkUn3PLrTCA4
kEiSDP1hHA1NfJvkloxnzsUWNLiELAztU1h4zXrkvogtpl8qOarwBauvc0Q7UcBu
zwp686tE3slQhRdZLzjBoQtwHqkD9BcfykkGdqPstL2e6tY7G79XaqcwlRkCXahf
Abq1cQetfUaJFSYsOgEZYfsCYXbOtan2JW+CCYyFo1YeGkh5kDZQhQ8frBXMDr4A
YWd7j1ASyCHpj4QmcjbrwdOR0R6MbS1vte0vZ9Ip33ui11NuSVx1xpsbbx1YNty5
xIipc44kl8OvsnDNgFnxn8aBgb4WJLRr29WN71giz9mj3wESnVhAZPHDYp10ez/6
pnCmpY9O+LiW8ukyNXjN5WG4d9QfeuIMlbZHCeapzqF2lul1V473+ftza0akjCdT
lvGCHFb4oQE+30UotOTElP2rNlMtBLMbz3RQl79tjDXAkE4b2maAAC+5lCdkbr31
s5yaDy36UjD8KrDoZdfnJDkupJkC6sNvDqcoIj42GvWYOy2ckJqoARNuwjM8NjKy
66QhUGuwRw1mkOatWRpF/4Oyk6QFtf74VTza6xc1DfKmtyd6afYLpatR3x3HTYgU
kDaOCfhgF6d3klpbXScDfr8aPdNNPMpjzkY6KvZlp1bjDA9iH/uU5ZYOgyK/3xcs
yiYeTfXPw37yhTprnSM5nYFyEB+8y6jQt8dx2fh7QJED0j4SU6Ot1EN518Z1NtHK
ncS+L8cVooIVVV13kQ7HClV+blA5pu3pAjzSkH/eTO79dZRDNpOwWdkdGs7YjHaI
VVdwcvdsswMwmbUwbMQwE6ix/F1/NTVgKYxHkpQ5Dbg+awxYBK8YrO98/V3JS+to
`pragma protect end_protected
