// megafunction wizard: %Audio Embed v13.1%
// GENERATION: XML
// audio_embed_top.v

// Generated using ACDS version 13.0 156 at 2013.07.31.16:42:38

`timescale 1 ps / 1 ps
module audio_embed_top (
		input  wire        reg_clk,           //       register_clock.clk
		input  wire        reg_reset,         // register_clock_reset.reset
		input  wire        fix_clk,           //        conduit_video.export
		input  wire        vid_clk,           //                     .export
		input  wire        reset,             //                     .export
		input  wire [1:0]  vid_std,           //                     .export
		input  wire        vid_datavalid,     //                     .export
		input  wire [19:0] vid_data,          //                     .export
		input  wire        vid_std_rate,      //                     .export
		output wire        vid_clk48,         //       conduit_output.export
		output wire        vid_out_datavalid, //                     .export
		output wire [19:0] vid_out_data,      //                     .export
		output wire [10:0] vid_out_ln,        //                     .export
		output wire        vid_out_trs,       //                     .export
		input  wire [7:0]  aud_clk,           //        conduit_audio.export
		input  wire [7:0]  aud_de,            //                     .export
		input  wire [7:0]  aud_ws,            //                     .export
		input  wire [7:0]  aud_data,          //                     .export
		input  wire [5:0]  reg_base_addr,     // avalon_slave_control.address
		input  wire [5:0]  reg_burstcount,    //                     .burstcount
		output wire        reg_waitrequest,   //                     .waitrequest
		input  wire        reg_write,         //                     .write
		input  wire [7:0]  reg_writedata,     //                     .writedata
		input  wire        reg_read,          //                     .read
		output wire        reg_readdatavalid, //                     .readdatavalid
		output wire [7:0]  reg_readdata       //                     .readdata
	);

	audio_embed #(
		.G_AUDEMB_NUM_GROUPS        (4),
		.G_AUDEMB_INPUT_ASYNC       (1),
		.G_AUDEMB_FREQ_FIXCLK       (50),
		.G_AUDEMB_INCLUDE_SD_EDP    (1),
		.G_AUDEMB_INCLUDE_STRIP     (2),
		.G_AUDEMB_INCLUDE_CSRAM     (1),
		.G_AUDEMB_INCLUDE_SINE      (1),
		.G_AUDEMB_INCLUDE_CLOCK     (1),
		.G_AUDEMB_INCLUDE_AVALON_ST (0),
		.G_AUDEMB_INCLUDE_CTRL_REG  (1)
	) audio_embed_top_inst (
		.reg_clk           (reg_clk),           //       register_clock.clk
		.reg_reset         (reg_reset),         // register_clock_reset.reset
		.fix_clk           (fix_clk),           //        conduit_video.export
		.vid_clk           (vid_clk),           //                     .export
		.reset             (reset),             //                     .export
		.vid_std           (vid_std),           //                     .export
		.vid_datavalid     (vid_datavalid),     //                     .export
		.vid_data          (vid_data),          //                     .export
		.vid_std_rate      (vid_std_rate),      //                     .export
		.vid_clk48         (vid_clk48),         //       conduit_output.export
		.vid_out_datavalid (vid_out_datavalid), //                     .export
		.vid_out_data      (vid_out_data),      //                     .export
		.vid_out_ln        (vid_out_ln),        //                     .export
		.vid_out_trs       (vid_out_trs),       //                     .export
		.aud_clk           (aud_clk),           //        conduit_audio.export
		.aud_de            (aud_de),            //                     .export
		.aud_ws            (aud_ws),            //                     .export
		.aud_data          (aud_data),          //                     .export
		.reg_base_addr     (reg_base_addr),     // avalon_slave_control.address
		.reg_burstcount    (reg_burstcount),    //                     .burstcount
		.reg_waitrequest   (reg_waitrequest),   //                     .waitrequest
		.reg_write         (reg_write),         //                     .write
		.reg_writedata     (reg_writedata),     //                     .writedata
		.reg_read          (reg_read),          //                     .read
		.reg_readdatavalid (reg_readdatavalid), //                     .readdatavalid
		.reg_readdata      (reg_readdata)       //                     .readdata
	);

endmodule
// Retrieval info: <?xml version="1.0"?>
//<!--
//	Generated by Altera MegaWizard Launcher Utility version 1.0
//	************************************************************
//	THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
//	************************************************************
//	Copyright (C) 1991-2013 Altera Corporation
//	Any megafunction design, and related net list (encrypted or decrypted),
//	support information, device programming or simulation file, and any other
//	associated documentation or information provided by Altera or a partner
//	under Altera's Megafunction Partnership Program may be used only to
//	program PLD devices (but not masked PLD devices) from Altera.  Any other
//	use of such megafunction design, net list, support information, device
//	programming or simulation file, or any other related documentation or
//	information is prohibited for any other purpose, including, but not
//	limited to modification, reverse engineering, de-compiling, or use with
//	any other silicon devices, unless such use is explicitly licensed under
//	a separate agreement with Altera or a megafunction partner.  Title to
//	the intellectual property, including patents, copyrights, trademarks,
//	trade secrets, or maskworks, embodied in any such megafunction design,
//	net list, support information, device programming or simulation file, or
//	any other related documentation or information provided by Altera or a
//	megafunction partner, remains with Altera, the megafunction partner, or
//	their respective licensors.  No other licenses, including any licenses
//	needed under any third party's intellectual property, are provided herein.
//-->
// Retrieval info: <instance entity-name="audio_embed" version="13.1" >
// Retrieval info: 	<generic name="FAMILY" value="Stratix" />
// Retrieval info: 	<generic name="G_AUDEMB_NUM_GROUPS" value="4" />
// Retrieval info: 	<generic name="G_AUDEMB_INPUT_ASYNC" value="1" />
// Retrieval info: 	<generic name="G_AUDEMB_FREQ_FIXCLK" value="50" />
// Retrieval info: 	<generic name="G_AUDEMB_INCLUDE_SD_EDP" value="1" />
// Retrieval info: 	<generic name="G_AUDEMB_INCLUDE_STRIP" value="2" />
// Retrieval info: 	<generic name="G_AUDEMB_INCLUDE_CSRAM" value="1" />
// Retrieval info: 	<generic name="G_AUDEMB_INCLUDE_SINE" value="1" />
// Retrieval info: 	<generic name="G_AUDEMB_INCLUDE_CLOCK" value="1" />
// Retrieval info: 	<generic name="G_AUDEMB_INCLUDE_AVALON_ST" value="0" />
// Retrieval info: 	<generic name="G_AUDEMB_INCLUDE_CTRL_REG" value="1" />
// Retrieval info: 	<generic name="AUTO_REGISTER_CLOCK_CLOCK_RATE" value="-1" />
// Retrieval info: </instance>
// IPFS_FILES : audio_embed_top.vo
// RELATED_FILES: audio_embed_top.v, audio_embed_cs_insert.v, audio_embed_frame_seq.v, audio_embed_sine_clock.v, audio_embed_sine_gen.v, audio_embed_sine_lut.v, audio_embed_sine_ram.v, audio_embed_input_fifo.v, audio_embed_hd_packet.v, audio_embed_sd_packet.v, audio_embed_strip.v, audio_embed_control_packet.v, audio_embed_video_input.v, audio_embed_core.v, audio_embed_registers.v, altera_audemb_reset_synchronizer.v, audio_embed.v, cao_fifo.v, cao_merge.v, cao_avalon.v
