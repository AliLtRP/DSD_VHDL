// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
eE3PoT9jElGNjUQNLuBzJUKGYlP/puUGQSwDza44Wci5LxQ2Cu0Hz/+DtIAoH2CX+kzznSRsgWyR
fmJnrZXfOHOoyjKgvMYQKXfzuadwi0eMAn+CbV722+6Wy4A62XXI2Yk0uNvCa4gEswhOHeSlIF5m
L+0FIJSVVJyfUmZYiBeSd03yIJJ5o40bAPFlaug9ueUssYNinfXcDXKmH3COph6UDm1oIg/cap+A
zONYzUwRqf02WQvrrsyEVpkCGLZeUl6wHvekw5pJeOjVFb2/CzdEqxqhd0JKyh+RQuK/jB42WqPv
6HPmlj6aVBKsdea6pnt2LweeRX5/0kwZJ5xrxA==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
tuRp7A0qFVa5hKt5xId8FJz2xrO4m9Lk9BN4Ml+7fOotNtVUnPn3Bd8YTk0K39Xedr/8NbxK8azy
7M+MNu7rQgocmcVnsS41QwmzJoM/rAV3RZpUoaFrn+0xfDSOtR1zeeXWe1779JoONkucwIcG5/3r
IYCOUTJHpVnXp0WePK0u2yvFXugvPFWo5Qe9wPguAjpKRMzgAQTSs99zl8mUMTOBJqPNfWdXCf4S
8NdLngCHd+6ttKL/fAfH5iZItU7s0Zqaar1yRhdukfquAeOifm2GLu8o4FdZ0MhM49JeSiQ3TbMt
3S0nzuFjK++lxa5eGhDuedDr4ObwWUJA9pdQ7qWObrkqQfA0Sr4bmH4W4uUoGlZ3kDcC2f80ojdq
x7kZPT4IXCBPg16kI0THSQ7t8zpQFWGonyDN7ADewviMI3WpjGbY5ZV8bxtN9IPRae2Jf/aXMJ3i
yPEchmxhPIzCL/YdY1oy54TXoZrA9jE4RoikvWTtcjkb2GaFHd5uTnECivSqhezoKumoUvoWGd0T
ikj2Bhu76Lz0X32mRsFvjlXA+2m5MwHElPhXxyXgfWV2GVkySyFnM81l1ix3Cg2zSs7AlJJ0H8yZ
RH2OnndYUp90VAbzeT1X6dGxd1/hkMjd3yyx7gLpBeNrf3h6CRhUTnL/+ntm+mzpeQNn7A3qYtXl
i0m+ll/uYQwYaFkw+S13SL9MBV4sToFstRIJyM897btc76FCL2DHNjUuomkczpPRtoeTCXalwXPN
FdBtRSiZpbIaVdKcUsfgm7Z17EGTqqVLtg1NXzipiCn34qtuJ74n0tk8G8pKaiADAwJ8kFxSdgXm
20Q63oe+Pv7JQtsDko458qSt65+6VfJbDMC+914Hqj+D1Rt9Zu7WdmyAJrkx25vnQ/r8XOC5/aMd
4jboL6CmCzLwtlUb1JLjtq0UoBrWNjWZMkVSisxgukuLWrFsbhfUQn6g+q6dIx0C3UAc0/oiL5vA
sn9MWPCvn15E1VqP0qSg+lOZexL+zl+oftK5t3DNHZ30MUagqYmFJmDJjz90Nt4/RibyL1jKZbK0
ZagbKXLRdCXTAMqlF4g4Rn6DbxYax4Tu/1ZXgWB7HEI/YbLJHZrTeryyXXyPuGIwaWjd9GSt6B82
eDbcg87cxA7JJQ0W5fAcJ2L76Wymacjb12Ammd7SKGTxyveqJi2tahj1pJU1hgLF82o6n7pXT+NT
L3VRA0mLcjJrAQeISNB2KCMC1Kq1/35XxRJBBefBSyyUTXGBTgO8ZJz90wDWslYyfvixzeYNcV3t
q72JEHvYMXp0mfo3YrUPDsx1/GnWNf3v9fYMouh/cSz7hnJZaUWBf3DUVouWzlmce5k+1njfbQkw
M5jQVuBwxYQJ2web0/dpo5s5Asi+7GZpExRl485juj0w9STq9zFwkcALpMYwzqP54uHGBqsQOsYF
DYbK9jj55DE5pdd2Zm3MNVI+oOT7JBA3yZcT7LgDOUU4EHoevUa8zhVeIrQ6lF6Va8bThv1fET8V
kUX/RYeFI075bOZ9c/FpZukXQc4d4jlRDrrUv9M1HLjGxChZjbhxh3X4Xu4kVVQ4W+R5xDWvXglT
dfrEkgFZa3FBghbis2uPqlgQjM4UUKz0cQ8zI7U+CKEOaxCRmllXxQXaB0HIxWSN+EO1lj4fajry
8A0ObPeHUAvxmYT4BOGbFXY280X6dCm5Gn8mM8sju30oQ5PtbpfDTOEbEsrOqHTwVnxSkQ+S+6Io
bAEEaN5SsF/n6uDfvPv/VLGN89BiyhxAXvLasqCYt2O5KIPbWG+gokmH0M7JgSvZMXRlNdaKl6Td
BauZ3zOqAo84bgaeeH7JSQjamTwQM/YlUkX/5S9LhdX0lAFUgTLvQB9ztvBbAhAKU3CqNvLX2tVR
lnDcO4f1rjXe+xnSxUk7tm7gMJ2dWCeucIg754OKgEWBTlxZjLB4FXBOiPHQw2/5MFGoVwGMsfW1
+AZJvbhRE+0ze41/kXf1RC/Fa9Ndy3SY/R9/BNiUhLCqp7g33CuGxy3YBrdSmtjn0ihZHGoFeZXt
9HVVzdSd5etakr0TN8mnbdW4yFFboHirVhx5EfPBV6+AF9o0GmJ/AE9KmglLb4yNw2eLvzOPgiRo
X14PuSmuWbsmFek3/YvlFJTe4J0OiCFJ+2sRiK0Bezpx1N7TdIK4Hyngor5iMutBJvh52xWJs9Ld
tZQoESlGQZalvF8m+lD+nWRliSzuioYi88XJ0IhDQz3s/WAWPRJg/Epfgys+Wnp0UnX2BnyqKdtZ
VPWzhXPEXHywFU5oDywIDfkdc0yk0uRiXHSo1bUTB40sofgkyleyKMeHX36XmsF1U9rLUIVN5VQl
MNEllxMjx39QtsGunDxQdnLLPmgTqIpTd3/SRKWatxPY7To2STLmaoLuUJ2WwhcpwOHrIKP+xzsZ
wz7edQK1O7dcoyvU/kJ0INefjf0+UbxFf4/LzM/2jdlbjFRBa4bCH9wGNAGmy8Z5Hn+oLucLnzoj
GcEx8d2sFWkgALd9gmpErT0ggAWBKxQMwlnl/kM3hfPaPUvzp5vmxRq1+LgkRWnjYrMiAS6Jg9nH
oKKocEvo2AbX7G9WvgiG/kFGXeBk0u9sksqLzc+dZp81Dpcu/2cVEGmYU6WfBBbWpPZvmf3MfQQo
20YJL5kWQC9emGVNv116nn/1sVBLjX3iXg/z/XJhzykru7eUuN2IScvdvZlQ7osPkSbGTS0Qv7Xo
EQDY3O97zttgIhYLoKoQ0GxnruYwvxeWItXPtfH71dVeG2Fp3SKWzrj8pNDw0QsMA/X/2th0L4vy
jT+H0+HehV26ue00BUWtu0M+Yjl0yjsyvYt5kq0/tUtVJkionbNc9a2SLdjb3sQyx07js7irHtkZ
Zc822ODf2MAVZPqFFzs8SzbMgPH6h1/bKF9JXBAqTe5/xpj2NzRHxbOF8lGyL6kYPAUqsrj9cXER
g6eWFn0VAI2dOQCch9lwBXOcOFvru1h9ehsPaIZlDsWeD+5/Xp6wyWj6Zwm412arLc6VhfuJPBSb
70twPZ0P5cvKz5iDAxqxrlZivFu/e07iPrfFognNLFLePo//MR8RSgf93nelYtdC1wy+54Kansse
FgcHjw+AeB7ySZwGPKOyNQJWbTwPWo+deEu6+GL+8JrV3dyFiyUGaRNF4h/k16ILaRNY1KCGDVYN
4SczXRppu0D0wurjNVHJopBWJ/hXWHTFZlpLquQVFled4BpcWIrGRhY8ZngWsghR7FfHFnca4bK5
9r+sIPx/33jmuUMn5B373XOaacdDAZTZ8zkMvc5naacwk0minX2bEnkWNjT1heQHPbqKB63sNj0d
cv+4z+Nl2Z9NaIAaAFMKEqO5j3taZi6rayvUhlXbBaWMwc90ErQs2xumb9yUbnvIwhTjEdA51zFu
DhtzVCfdWHcuj1vMUppPMskuNPUwIoQWwmqf/jghANx96XqwnNIvHLzK7nAy43nTV4NJO9/BEHji
3osR4EL0t9ISFtkHsW8dROH5IQgL7ByHIPSMEhvDNHemehN3Ke88dvzK/trgdXWOwKKveMGbZI10
Ez74ZU9UurRJqaNMKyz95NPApTJgqpvxoAJ95kATOJqpFWb4PCtfQZi7Lr98MwloeTY/kqiCBJ4e
Y3ksPBZfOpsoXZYZlf5zpdSu1zGkiSiLx94Z5px+mGj3ztot/aaPBGAJxpKbU2SAmgcENCMOFvF3
+ujZLsOrQ4kVNNX4wW19EoEwTCoPtds61JVkkaBvWx4xx6ZooiUGKBIU0f/7GR7WUAlYMQhp0mzk
Els0glzan7I2paYpNQMC6AhHrKsezhEKmLqwCtrPPyi1eMAv4KOlgUsy/kXZQULItVXn++PfAgLq
PQpML6eNuvxJB7Uggc6QFMTY2nR024uX1Y8z+muWT85fDsZtJf6bwrLDJILKp09Vwe3v6x6HZVQy
351yE1Mtk6jxi2drn2L22DWCMlmJObnvPQIKqb+WqRZuWInxjilkoJxZbhipGgGfpgWvYwvhYU8E
y9GbnS2tl0NSo/s+nD3IHLQ6Kp9x0c6dAHmb65AdPTIr1iATQyAtD8CPkFs7WgpEOZD6AjBaYpNf
fkPUO/mJ6HMTlVHePC6mFPOs3uSEqqCgtw71Sq0dEmcohKNkkndwA/twK7bpGZ2ty7wLs/F6r0OK
nmVNYNJKyCLFDmPBY0kfCE5ndb3UipfEqVyq2W8cAVQ9FNe1Pym6BQi0P2lLQ5pDHiA3Zcb/+elb
lN05qikAZXxaKyKAbTDGJ4dsMfevbhGUzjwWepXQw8ElRzwEmSKwxtXwCo8NT1xk3QGgyDsOxtJl
c2IycFhAOlMflM8UrkiKp5z+KaLVu6hAQBspwjusdcjE9YXSr2R80czhHBnOvjYEpcK8mjPKyee5
psv81WrrNthJd2MAyxPF00tqmUZECxLpYY/SVEm+QP3JYeyKi+re9jlVDP3LWTMzaSuqNCyoH9eW
ZC8+4FTkCBEEwCBQTWgWLPgXSsYttPZ4D/O3w/+bjdjrMDdoleAhfrvRt0ejoD4ECv87VuRlzI/S
TyD6WQvkmekpW2eHhM41o3/zd+qR8Tg7XsW5Uq5FwW2qZlhRI+cCKXQBr7We6056LBS2mkc7vKVs
Lyea7hkAS++dx/OmSp/Kge4//7nT0ONmygUBB/dyR4KoYvpPIg79KlzoxN+pfVgeLR87/w96+PFs
2i5V9Pv6lxevbI1f+7JEZe4a6NWuefTMJ8UqbsMcITpAuFqQawoz2EKyXoU0ZV9Z1OCOxYob3cTk
rK4iru//7UZJeCWD7xRGDzn9luKu90/jZEZ5ebrqP8jLu0E+kfA7Oj49urhbxad0vztRLnccbgJH
eJmDdwUTWJ4wUarEl1njmetPGvrLEZ0mqRGbTsMVDtcbVxUhe5Y9igCHRs59bTD/rcnI9MBMPsJQ
hkhawMC5LB6V04JwfmmHkopdnXdPyOzO2YJ6kOvQHSy5Sa/uDQBoE3kAcKLlNkaC91XpyONjb4UY
inSfkiBQgDc0/Qlc+6u46WdwW3SoKD+02Gd5RHC5j+uNaazP3i+WvcF1GSBCOlJw5zoAMwcG4L3C
IZctShkvJL5ZKMx2lgzfoGnXZ8LhMNY0RXp66fTRz8BNi2MpS5eq0kcYyZ/bzLUJuFrRkEm0zzLi
osNgYqPv5qxYvMvRHz13+TQn731XNXCuuaiTUGh+PKvFpOTMq/aINA51D3rnvecbu/JuVjNN5t+h
IrCO5ZL8cHagcgc2zKo5wecPCKpuV1GN504e5TYkqOvvqAyiKT9Qc9kHGni5r4l1Psy/WIrUB3DY
zjDtwcCLd+DgEmSTl7tmorOwA/bOhyVLXnhm+P1tIL2WcjVTsy6es6G0mNKWPyIgYolsUbLN7kHc
54sOEI3e6zBbv1l83xd/floVp1kD8gaLwSJpT8wnHVgYQVyhjEBPxbMAJE5twFnfKsXI9caHODZg
Rk6qoEXSqMe9lFiyBKFKXvrziAjxPY8p2BO5vQ7dxcwNExytHY14MwZOLfVl2CxzcwOEw/TRN7Md
OHn8PUJg2y34Dlg+TCTIk0tIGTCBkwrTsnls9liFyahzu4QqPn3IsfzFscURIQGm1IPrjwFp6y9f
/I/2Y1l0SuPsu8IErSWxvi8of0mr/yfU+WzxkDOCiXvffTavhXfRG9m66x1QxdgWejz7T8JwTXjy
uPdx1GV1Ih06K6AeWhUITWNmju314zBVDY/8CApeWt/DeK7H6DBuRW3sTDy7UGvIqw0xfzcUjE2n
RxRXjlp3CWd6RQZEpPLKoTkIQGPXNMyiG9Z59HtBGpTb9hbfAnBAP29isv/Z7h0RjGGVSCuwpdkI
7eos4FNwhQIT7TZsUQMSxf6WGqD8wgTq8gI+g2hSc7XRRZ9Pzr2Gz1cJwvJx5EV5oQE0QBy2ZNY3
6GnlvjE/GN0eJrxLQwcicP+w0gVdyhzgY45CW9D2EdBUwFi4YBwEvGKAZ0VfjZfNRk/+n1nShu2+
sphUKpb6HO17tmYD3duz4cjQ/Tp5zAXWtRKGZs4BEGf57vDa/emhGNJbW+/lHyKjzXR3BJhQOaO+
4+Fra+gUUwwcQy1/5zZvo/ABtQesujbNj6TX7xW1O3YLWO78V8xwYGtkkOozDZ2/fzgZcZng+wnK
vWST4wbxRmO+9nxLW9XY79z4w5qPpiFpIV3b+PijZjoyED+Z4tc3TEZ2x+lV74s02n/JOSVqpOi2
5wdWSu/Wwf+3DvDyOvh/dD8NcixwGnd2h2txMLbcY9kN0N6D13yuxyhDDYjuRm7z8PsrV95Emi1y
8vsG+OUMIOAPqSELNvR5ugs6NO8h+Kc/viqgoMRVvP2/JIn4dWV4wMfRh3ituGPiJhKHK6LzPZ7W
F/XInvGUuIZJKGf11NDR8tA2ocH4Nw4vwxebyIRuhqiZQEMWOUR0jFvkFth8MbNYZjwuKeQrBlMR
N0BiTO6EeCfk65Aa8L0EKRjwAsZas/KZutcFagQ06P4rgKM+A7XYjLzMjBl5werNE+5hqpZ8OJvX
z/KDwYjnGQM1iP6sT4NjaLANVWkT4+SXeAu8hGbDCzDCkGxMZN4Qm9A3OxI4lgA/6CqgywPCHj7b
TkEq7GpocG9hvs7MCsBCBv2DUhUy3sXp1qV1M9fTF/LByaTG3TEynk0lxeAB8boFDOe0yUUYD+bv
VdK/25f5Y3/+qgumIPBPR9IXO2Stb2A9FAJLz1bYy6DwlQ0qQMRI53INIMO/YcSEcgppNcBV2hVJ
q9hTvjz8Cz3Y3MlLV8GyiMCQ0gY0JaU1eEf8dzq8+kMo5+7VvH7s1n67ZFi7RC/Ehpap441R3Jto
Ji7fGF1LmbPGD9bO+AfKW5BO82VBbGdmeFMqGk91vVDvvDLHTE1R+pWa54pEGvtbO0N3W+e9INqC
6fvoXTTDnRkvcAN90aBzss0oB5U2gOZZLswHku1DZxX2zPG66IqzdaRzxAXdNzseSIOeVmBdKpAM
g5a1X2m+pvsranpk7X+cLaB/ffGUSwkcllQRDORz1VZPLIG5aGSGwbxSoTRv6QSVhmFLphBqw3h7
+bvcrG687V5inX2s7dNHf5iZLHJ8vdjvY13RaApJmTWnw1oekv1Y9gkg/KyTZXtbeCN38x1UTAAi
lkuWSin+yaMsCxYjk8HID4HBK4yN/I83ffF3JZZ7rZGY7afsnBc27bFIKbcir2Wb+rSkyTTP0rSz
dZx2Qb0utu3xQ76Yqfz2n4fxlPZkeuI5rHnTnF4Nuet9UweRKx9kZcLsG1ID93sEBGHkl7LaDoT9
+0ivuXbgdcLrDlDshv7P9YI5xSe4ZwYueRC3TU9AI6OUpWGBUeS7HgRqJBq4cjV9rB3ySSsjzzaT
6RCNpDhCHzE0eweAGPkq02E8WB15SRu8Z4P9lCy8gMQj5DRBFr/yq8REPlrC+Wa1mXXEr1WiwkTK
90miIRB8XIxMx+dYB4Lbzsvawr/JV6MPQNmyuf0ZJc5lxINaZgdFCJQwazyoevf7aBJYUTDorxXZ
+FezxDLAyy5Y02P8hGgbYs9pdEWRpb/ldGONJfMv9AFpgxEKyaZL56ucD8hFS24+wEQAYf4MRyRf
0msG6/kZM1DBMFrFxwGiu58JjOweTTwZdNSOyCsRzNyAUcpNzz63bt5eI3Xm+vGKFT/4M4/j4gr+
GvuAMlxtoYr30X5wO84/RiG2rA==
`pragma protect end_protected
