// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:31:47 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
mfFigyVmFlWKeUFCZAQmahTAG1RocJolQT38JSB5tXUiR1YEZ/yTeaGpaeBXOZJV
aXtya7+VFze3fnG9Srs6hqRu9REVw9e+hUMWc6RH0seHcfNPuy6M/f1KHzDZII5A
y/i+KndpJTB1bygZZmyGM+aerYo9qeZlnXS3sIWkhJI=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 37632)
p5jTBmdpN3Isc6tqxs5CffJXpx4uMoA+9+Hf5NI0L4iTqGefyn0NsLdTNxudEWu9
f9VwmKfF6/LETZAdluYABYzawVT6Rw4W0Cc3mowzeMYymmuHOkVuNTm01KIIEu0n
xuCkndGpMMLta+R9X02HE5az91bFr8irUDPiwoh4dkjNt93A+P7enQIJAhFp+KAT
Zx61ncdyb5QOxnO0BTbd9tlcXQASNTTDmP/QLDo5Xyk/u5GVa2qzh0+E2xbzwDkk
sWiUuA3MaYapvy7bL/5NDyi6D4ONINxHZWz2wmn9g8Mp3PmhBbVtfe2cfGOgWFYA
vVaAPRcXRlgemN5wLmxPuNc5NufEkGTVdHyB1DYqlkpsO6bw2RTGYLrJGD2Htoj1
1CTOGdNWyDbDXIsH2F/XhLgFtHEIWzQT0rnvdDPNRPlj4SPwxWhbGkigL8SSw/wj
6lHmwLphKaQPfnC3F9VF3QY3ApnY0SKRZevzOOzfNVWoo+PM7s+YSOeFv30eLN9i
WHfH1x5EiuXdOPLxRDvKNgKNPwPcgNBafa+OS86guBsp8pw+ZCnyQ8/TWjiLuOta
WdNaj1d0wfJJIjxqbP/raWrsKJdrpymCVpNAy0XIUOnzOVUOgKSCSykvXxoEHTRS
u9+A971R2Zb7ASml8MUtlVLOYpqC6iVnLEtlWXoYcIdU7BLrvQok1MDBrIJXqxIq
gc8wOY1NcH9q1PnqUnTVLyJMHFe5Y9saidZnUVN6NXQ3YPfIolmWcohkPDI9MNqL
ttkGpLsU1W0paMtpsUJVmG3xZCy+iS/aa9tRzRkdzrap+FqhoemHtj6NvTisBf7Z
AxGXBOc4I7j7Jf70ODfkPWcdNXmT2x3BkaWSm1dPynunSgnXcVu25Hz+rM1UrUKh
P0UcVLC2kOZj0a3tfYngNUIVO1k15uyiUNXw+/ywbqJQlRSc/SCHxZE+YsHzTWaV
LC6/0gYlPgTFUd4Skhp1+M39VTCXJYb8yrfRycMsV1EFSSapS/O1wWxc20Osw13H
p3EO52jxLGVWgopRH71uPPobGJDZD8U0daQUhQ3DteCdIltilGYr5erm7mICbRrN
DWzUy4b9do0JEOdOGDJ5OmjIG4pqYlDQqE1S/mKUe/+5tYA9KcGdC2a2z53ni5u8
3JEZA74iKgW1Y29vE+PC+X6Jal5Y5XlPTebAlwjjhIkYF2mUD4nirh4BqddmDUkz
alQmtwdffHV60PlIF2dSmcydAQMUov0Z9sAoI9XxXhTC9JDbRahSPTMwg9rAYXA3
3Fi6cRAPYwCc+opoBoEsgw8nG49G+0sNaIg2aHus8uq4EIa2ztVEmxshNZVAvzvE
auxQvF2w1h+/XNIxSSDpCl4YYmMYugHvfa27I76rgG5ddc5JNsYOYGXrMOq9537f
97rFDj1rmQg32QxpZ54Fy4ywG2vKMzXG47BVuE0Pmlkns+BpV2DPS68ySNfi0noX
nG+lbqYc3WXwWkJCktO8EqTjoKD5VhvlqhD2Zwifks6R6QsjmSBWiSx6IE0u9yB9
V8IwHhYPqVMbcudV1sjG4yqdCGxzJhJz6vffgbBa1F8HLgnP5Hs8v/XFlxDPvpU9
vv7ePLB2xUv6FIErEmW3j6frlBxPrjbZCVBvX4sGuQ+Kckl0yi3mhoU4FVDybtqn
WmuLwaN6K+hK97U5VXC7esE3oHM1hv77ab+3p1z3owDBtCYbGD+GMjjJ2BAm0QAV
O07ywPk8Tr81n3NjQ0wO12uFG0IgL5MsdTWXhPb48+Ly4+O1R5IoJYicrgDGhsio
gBYr2kzDc2pa+UU/vq8W+0pq7w239IWPsEPdaQ7aYInmmnzd+6kRPUUuw6U0vYjt
eUFnBiN+94saZEAaIa2acrp6znez8LRyQNAIgzciR0yRERF367+M7MeBjJ4ayDtJ
QdVSfsdoCPuHp3Dy6r5xyfd+/PY7uPK7JMJxTshFBh007g6yzpTmBk+qCVBy4DGv
hyXfHEh+R+Rjwp5wVOby1bKE33vt/lAxJ6og/W+Vy8F9LB4ZemoUFB8wG2Ndewna
8Wqn1cVOhFJudv3tl9M5QeS94gC2f+0zdVsrQQ/8MdwksMv5fwc+XSGIKiiqewTe
0ecIDgtlaC/PdEgtxn2isIZD2TO/fVig6OCPC5m3k/ifEumidwgk+Ozpx8Fuggct
owaGUFgGolrmCAqMjmFKFM23V9gxGoBa7b+l8hN+CFV/4CyfCyj+pSDM/JQYThE3
zbXhZnKS3uWlACZ0KyatnOWXCVECoqK4p3NzFRX+iGDzcU1abVz9/FX6m6Yasl0s
OMyD3Sv5KxPC7h5Yy4Kkk1osO4tYdenMTQG+zfKgmYmF1Rbl1dYUCYqP1L3QI5/L
YLBm+xvnc5F+NN8LxbWLhBP30+gUtbd6JiUNyS/crYRONoNBA+AopuJzRTpdoeRJ
couvVE7lhFDw5a9bGycO8OiZZtKsyrOULawqJyFBGvq61EJgxVqJaN2Ba+qmRTpR
WSdBNOBQdYXIpf6V7velND67vorWzZYtKSBCO3JlOwcHaeNxP03wXOv4TORExVAg
S6LIWGyVE0IFQ7bvljSlgXUzEs1ZamfN2fmznXcqsYbWptgKdyQynIx1GScR3nTH
UIfGSKL6f0cuUEDYb/7zlG8P+Nbm4l/jGM5M2j9wdmeAp2++u+ta96jkdwCm+ucL
7btB6GoOf3WOGaJr/dG1uC/gdaSF5VhjTO6UldPii1ipeLZh68pkQPPxwwBSGKCV
wdvCFQ0bcMnT1ABpwPc5ZaItCHXEVnV9VlMkj5obvuaehYm8j7tntuo181UaHBcR
jUl15udokeZqkdgnTJPLGRXHbvYYvqlOJXOoY9LgU0yQnYrTn3HHqbPU+8jzx/4E
+zknzxzgsfkwlR/Awn4cgprtwJfei0DzSbZvu5V3kBvsW+kCDocCipm7LPm/87Aw
9a47zu/AYsyThTKnVBwroJ4u9Otoof85Y9e5TXJEW9hIcBlJOanXcSCplAq2QB2k
Lb9WpCql2Us1iPtDKXpZGrUAUJrdIV5zVDQ1NaMbpPj9f8L0ZxrzovVxCKICfsZ2
/QGOAksVxc7dU3yWuyta1Fd9evXm7VZIfOhh4AtwVvXFLMDFf/5rjkYiiIWdgfkG
KDye58tOQ9m22bUoRENmh0iuZ+Mq2nASR+b3irY328ftKHKs0E4wvqG25ZpALhyq
ZUjMZI2Lhiucgmyx4D+faeIzRrW9lP0IEk4U799bM7KKj/knodZ6WqrNaI98OuCr
TUpbGLA7Nm+ZbV3ivlKKPQx3AzS6Okpwqbh4NZfGv9YaoRvPbL2pCGt5E8JlR1lg
yhGSTYetZbJzfSHWivtDCbQdPSMWWdrwWmZGHiWTy8MG65GCwdxykRYQNwFceegV
d3nNPx+APmb4sacgOYUigxSp5kENQpdC7mUuORYEDxJgL58CZgp5bvFZICRCOWPn
KN8XBReqoqBXKNC92ILuWJKGHBUJbg6zqhNkHhEgDbrbM+NTJ/AzF3Da8+EE7v/z
Ryp1uusiOFiouh0bR0AI5aRSOxpQYHW2mPlVywsDiRxVvOGsAraHwJdiOy8w6VEY
/15oR5NZTds3RSmn4QOMp/dvnMbjl18mpsbg7XZxZ4GgRgVTHgLGoga4M5tQ65iN
JBXnogba+bjWuAscxlV1IC4SZLX+vXTbcTJzAjJXo4R1xDGfAGJ1d99BTRKK4LvY
1nMcaoOGR3mQVT0bzNIORcmz+FW2a8wDTB+lp8Fj07/WBU9HXGgtv3VJVBCMJYsb
H8B23Fe1GVF+II2nCXAO2ySjHSeQl9nNX4x5vzkzLAwqYR8H/P9T0cDLLR+KRCxg
qlsXIGnYHsdvgSvlBI7rj8somBeorFDEi6L/jnXrlSPxNRC+qdbh6TvvTeHRhT5B
uO2ZOMPOMSXV3kPDo0ddvo4UYnqZ3/Ps3XYPWP3mxxQGj03Wyj+ubJdNrqn3ZkWT
+pHAPkqOo/tEPKh8Hw69Oh7ygcwtTIPc0Ap2a6sIexItpQR5sMGYmVl8otwmRokF
YY/dDSf/MInPMjwVrhkgs32W/XPH8C37EZXDSx39DGu/tqYbbvQYGvpv+FqwEghC
wAEdLd7kAuPEeOPeclVEJgOR/9UgTwx5vcozfPBkor+gh9/jthS1Ww23xZJCEfxa
BWN4sVPNPsQpJEtLhCnYhbc7Hxfm7nnv3/g9GM8u0k8tt/Ucc7zC+fPT1P7KfviC
qhD/kqRLdayL4itZTkSw1c98+6kAfvrFF19R8nWamHPGPCiVNHEs7YKlmMh/G3r9
Myq5P+eAOtD7BOD3Qnx0rRI7djNbuu0uoxSHtIB9H3z92rpE1xTTIMeaq3Ggz9u1
wbzksqRTpWhL8y3Ky1ivpGA1TMKTFrG40eU4CM+rq+ivn98kP3kWDhhhz4SZBeo6
lQlIiuJMIzppqG1uOITI+YsXZaRs8xcx/G2Fe/Omv6DG+xN3Yn3ZMGFqUlfWKrGK
VyrvG62w/IAwInXuwXAWsFntVzq80IJXx1SNXBBt39JbQ32c8Jv/S3yhZWyo166/
elQjrnPqZVdd3jV5xYvMHtNvIBbuwx0jeocUe2KfgR+q+cucuh+s2DbhoPp4pp5B
jJKohs3A6OSNhNu6GUqm6CV7TEh+NINfSjMje1ZHySzKaDRLtFmp3gVqoi0l3ZY2
zwcsR0GMgvJpVqzkK/OSRRbebMOixJSPu6J4pdnHmVfLEOkCp94bcfoPF61S0gfW
cChdwXpbtEtS+8GsFHCwi75Yp2J0YJ91jvD/fHkl9litR32HoOWXjg15W/+3UuMf
fGn4ogcDVDdONseIw8QuYXEPDOjK9h1X7x9kcOWz1w3kdxn4AAPVcqNsBsKUSjb9
VUDG9NILpyVYKZI9tHdP/OPCxDzgPVTj8wBR9b+p0BNu2zTLGIqp6jBIw2v5jhIh
OpyAdT0bxwkS/0tiD6mHdJsP5uW+LAASI9mv4mz2oDfzO6EiP0R+esOtkxk2Rbfp
sZShZaONBjBCiehpniOsBzNb3fcymXUAg94I3gxk/og9w709kZsgTM7e2kH8mg++
O6sjqgCu6GJIAj3FeVjQuw8CYup+yY4YzwbMfKUP1sf299OguW5Hj9gyCsLqnwx7
TIaOA60SQdqbzqkZLTaS4psTXdzjB74ONe4KgRkvTeaWBRRDNhsFP6hv3sv/8IjL
i0tUg9PajJqKir9DmX63vf5bBIwL+zdA4VQU/cWVrtSRNxxSj0CVMNo36j1i8HKU
tRnPNfm9eNCk1lPadhWgYpMbFqtYdfy0hgEiHnWgmApy+5zF06rV+QWDQj+eogOq
eNkgXHtRw57pefquWU/5I/Zuyxs4FFicZd0oaUy++kYZhAG8Qldv+b/Eoq714bys
Tf62dX5cm42Euv2kGSvQI4Fne3+Rsiwu6QHYLd2gKLVGHb1vYkQOn3GHrY8q8S0E
IPmhsOCrgGn3gdmCG9ppZlHKikGCPtChvr5dXIGjBn+6KDuQmWcM8YvBB8UGjwvk
t1wP+kJzLVfJB2NdwAHvkiIfW/ctE+o+AffN1A2fCIaw+1Auw8kgX4fqDprPvoR+
5mzygF3JBw4Qw4gvIGaczC/Vw/XIkEF7dUfvUliUckJc66ROGE4FxWR222L6E3WY
8lhB8xHhM8Xc0fiKnm0xagsy/ptev/SBGdobgtzIkJiIynFmF2DTKsWN1pwCsMwz
2jKbyl1+e3bBy9+ea7xUNpBhfIx5tuQTPC/U1+hoeGWUhncow3uZ4xnL2oq6WT+h
YD0h+PK91y6NbcH4gFakABRrxhb74Qdpa2ORn5PPcewqV/wuUXuOIzOAIAz0g2d0
b2Gjn0PHK1cj5KmSjbI6Ze76dBKokhuZ3u920LWJBZViNqYxJDQEn7VpkT9Z774l
V8bncwtIXBKDvbG/SWDK6Z4nXljy87ywiDTMFqSBDCTPWwnkmDeIgxj/B5hdwqvI
GFRNLssGi42KjqhUsBosuK2++T6zn6HgfNA12WrqdVS0tJ2ZXtVaysTzr6DTygfx
Evb14nUOgvRf+q019Pu5nQVN1TKWYYUU8+HssQxZ9EyezkKTi2CVXZwPLgjpTTMc
owvtc/iJlwWlP/b2qRzn4kulCCRdiXmlnkFJpfF7A9HlGEsE/vOFXtggawmlAcpW
an5qxnYbi3FHI/wBnPThhyIcOn/XM91FRWeKjP/NG4Nbox/lg8fdYf/7sxCle9dv
pAPLj0M1+oZvV9wqpfYpAs6ejL+KMCgBsSIAzXrC2jIbytMLtb/85Z5HYoZw7GMh
VY55+KvXFOldcWRyUfM8CE8WI+ZM/+ruNw3H3r4/4fMFWJv9CaVCHo8WXDrPYBT/
FLOU7hKI6PsPTqQWr+a4tl6MAXgmNFRf8FAHpfFOVmo6mGhMMJ+yd1W8c3aqjmD+
Z/DjIrTGnR1bEY3RJUyzLdbxCV1ELijbuzazgu0mJ49Uq11YrnR7fyKslrzU62pC
KbvhLvxvK3/qvVTB7YtbEknqkyGp0eLWjgXoYpgkoCwJVFzfj8K34stbsc5no9MG
/OsE4wHo5jCSULZQRdhWOuBj/95w6pEo8llq865hEh/kB4eFlVfMN6t0szyXMOe6
wGiBq/+Flsa4wwsximudSiIuPMgYe/tYQ8eW8XWwTD6CAErOEvngVooJ3olm9D4R
Iq2EQGfLQs9zy2umXET9zLHhIckx2JV3paChG3CDPhb9FyzzPwaNPSCq7g6/Xo+O
zPLSDkafPBLQ47hAUnINrnm+ILXSPMwGOTE5ARrMfPMTlk2MVnvhKDc5P+daSuUE
NwkHghrL2xnL+LouA0AVVCa7/KJ1hpixluNQdYZiUj+fDemTp6cPYVtisfewaSTM
3HtrOFNt7BELWwToutDBDA19zdOpveyAJZ24XW/fLRLaCbflcbGKbEeJPEoYRlbC
UElrQTuoUL8IHQ5Dg9Yyu7DUz5La54x7Dda0bnD3XD8+cQ8bo9rtU4kTfC5WoQVg
lXk40/zGLW5iz/C7b1/SBvA9TF/a7CclZqC6muL3gpdSZIMaWXON5pWlnj21uBKS
zr76tLHkfZs0UICp1cYpjGjQegEQSC9O901ZmDgUEQH7qN4dLg2Z9JPmkXix6It7
wMu/jkkKz4cK0IiERAj+7O1n3s//zRXRAi5rR5yN0UccfUvszYJhhDfY3OIWhgOM
/LC9a/sR1PPRLEPVQQMHtiY7k+Td7q9GvJ131V77Z/cMxHVujrx4VPTzXVNcaZOr
n+fNmqdWevgWY8sE31IjYLxdNsyh5QISpthPKkuy8TXroi4+1rKPd/jWJ2n4UL8V
fUyEjNjsCh5BwMynz6vk/cjdmjwZ9/NwltHgC5U4OXTJknj8iYjpZG7dDM8lyimT
TDsAW0coQU65rK6wPYBQIhuhh5wKhITpCb7Z6SVmz1gu1yETMvs5fqptZ5GvmG+N
Semnq63EEQZxgMWXH8EU/aTrIp4jFLAIm3LTa3KPyOVZGZTY6D9FUyePDseJMej6
bARNMsgOtjncjfiVWmF19UsGXUhXaXhTwMNieYEnhnZRz+Kpnqpc+MdBm/9m8EXb
9/mg58kPjhYXgm2NctKje9f64epGZoZbvGWEz+fvzePwfdKuNpiM4w+EH78Dg1yY
4jwt8A0AGfM6shRJ5E5CXYb4oNojlyFmMdAvRY01pedRTpvV4ocW5wIg3TgcUZzj
QGd2vwy6sz89ybx6CjGXpSv9Ugnwt9uMXXQ9UeIKP2bIlIbebLhveFx6r3Oqnhsi
h5ykwAEStY9iWBcKXBf/oQou4hOKf3hZaD2N90i8rCUJuOPIhPIq6qXdJCZ/ayxO
E7+tYQh7RUbXtZkh0WORXJKvBU78LHxrVUloXqq8jB0bF9PIHIA6NqX/oLvXhvoV
anHG63NUOE+0auyNalvMdF1hjQlabECxSkP+5GvS+PHIHdmLoKCsXIMTSDWmbm+K
bBfdEIgYMKELb0o3VoaoASTykl1XDUaoGzHbgCzpt5IvtsnmTOe7utR3TqYbPznc
HJzD0WfwKURIbh6UGgF3FtPfnwoJmWMSY0UGdgb4D8SxSqaMPcP5lgyScxUO/xAs
bu/UGPjxIn9WLoobsDSNayvfzXjPMrULKGBcCugTCR/3NvO7USx3noEsDLYozdEB
44Rdgdfy5kOdqrfLtvvicJVG6LI5d3dTxQF8PGbfaGC4RWbD9Zzg90SSTVB2Cmfn
YPthuO7LvKpqkYRz7q5C6L1O2+QeuEkwjgZ6Ingwk8f2FOQLYOiVvb++k9o56sv8
xnd+AJFZEMNpvHRtIX0CpvtMszo0lXDoPyeYewzG/BHH5fuI6ppTWQLUV6tQ1MRi
q07x7MOEtdPos1nRg9VMGQZFEQJ0+l/JLILY1cTdGaj+uJ0zvsONUkPSRg4di/SO
Tqs8GOL7BT7Hn2GlEv2q+Nq9QfP6YMlgadXjPEIwDtKeOC7q1dEJMBdyqwTNFb5o
vmw3iDbheaOC6hvHRMhEdJUx6gahx5BCbJWMLvfJ0n5XcglOF+C3TMLyMxY68Zoe
WxhJwUE5M6Fsx0hxJ97TGqeVDeDsjPOV6c60NkMRXFNTRHCMml3Qs8ko4+L3gW2a
Yt/0KTuujanfuKRNGnAJ2hXgZvFib52ZDda2gXTrW4lR6JFyFbLv8lq6VmQPPH78
yZ/mKO83aUF+PKzpqrdUbIEgMQ5Mm7hOvyNUkl3pnCtfWFucwQYaRol5MjVDFJyN
rASk1viF/Oyb8rozOBD6hBWqCk99ESXDmL/DF+NzCAGFeVvkQNGAuLmEfdCjCslP
C9o2fQ01CrEdxLK++2O9A6coYG4nbnibfenwoew3XJiCKBCIgp5+AcDIiywgReeO
RixgXqRx192E0sI4QbsCP01DUGWR9wWAvY/QeLBztlm5hJgJpKEILCT6Xa3ZLTz8
8Ygkko/tkW4ZmWnDbD7jVIsqbG1YBm9S0PmLL0CSGSpe/Ck3KzSTCrNzztFp9UMM
WCSIwhoAqe0GP48be/FuTJRI9U9vRlJCWTh0nX5BiY1a4EbouUeP4TwLj7O5PiH0
o+hnxyaw55VKdYiQe9imPo9JNM90zSKd+FcY4rwpr2M0leSyArhQP9+iDCC5Io/c
h2qWgwj1fcjeyHEyx4oEYLVepbnZhPCYfv1W7X0BQAhT3LAdae0budAzB8Dfj0wl
L5xqrZkLnePEKw+SD+x/IjVYU9iiJ386PNcBkAwh0hA7I2CiGX9yDs4jv+Eu0E5q
CY6e7UKXRBwzX/4+dLrO7KzTLnHTg5WE9fURhsnCA4obxXF2yHLsxvqgN93G88Sr
XKIm3W9XfxFcMbp/P8zrM6xaRWyzo770l7Qja3BckdPS70d1wJ6I+vJlYXlLZBJV
Im+EMEpUB2btcLR7QALRxkeMZGKXIAa8nxTvVYAfm4mcxcatJmrKtXiHqfeLL8s+
gUClLf1Oo5Mcaaf9ZB4sFUjRq6eKU6PtdBjVPA1DT0Z0rJmyqDWF71trkrb5B0GX
XeeIsvg7OeR++uIXNk5HoeCtlJkBnETcFmlGfxADXbtrNL0OMAv1lmsfcnGaEOGq
MSwtemJZROXDG2bgUwxWSCPJX9v2caI4Z2ylfkCWzrq1TnvSgqHUijFW3s4+CY6r
sSX+u6ruzh/zsYwRKff1uNrFWNskOTyVgyq905a1fTaw2v+ZgGNuGFbRagNqaAvH
qavB3IOSSrCzuZOs5Wzj3r4i4vXz8bx59PRKvQ8iMFPw8TwHf7NFuLgHndvgRgQr
jB1RVp4S2+JoM2xAPbl/m5SCmQRImV1ByaShA/2+swQ3rjstPisLtkjbSAjyYvq6
zJvkECOsQCqL5MeSvzttyRQlskD6zZcFo3Z9vsEHeMJ0zqKbY66fP5gAiQne22iP
6rGn6ljHEHHkMZJFAryfo4YLiuZv/jaczX3Z3F0/wBrx+/ZhcHYaNYOJ/lJUTbY1
HP/tXAs4qOIPpI3favIErQLzMvstbyx05wO36TUoZo2wfAejBauYpwoUhFcmOJTL
XAgVTiwKPD13yr4NZkYoAiw4/i2FYCOU0Y4e13l1XLf/qV5xzL3zYoAKmH8ZKg9x
V0hEqAkv5MZHBAWykGt9b89nQzClj66Cn06BWUoiK40k2ZPG2B7LkkPKO7BJsPOs
svVCDmf6cPtoXhs97OZUFFC1sd9PZMKOKAFoep8Ae6XsVUQ4BOmr1+POMVvuSL3V
oom4orjwLhiJPlX4xZliH1eVG0E4HJW89AYWvWz5PAtArLc5av4PUgDAY2gng1aT
n7LPn3vgSuI3wKiPkc/xhry4avLAoRbE00meHoh8BANlQ2CCwxuz6+47YJOnuAHP
GdX0HXQHothDyzRRN+ewbiRD2ouH0gHdAionSG88ajqrMLtbp1VA0V3ew5Sppl02
+nXlwMvkNfsO+jI9M0W2WK8tIj5LKXKXv47gF5GefFUd5TmlSYcAWIkggc5ZGwTX
G+mCJN3lHreGrjeo0XvVv9aFO7Pz8kLXUyZYGOm9BCz3YvHobeD/0QLxRon7LiK5
FGcJCFLhRy1gYLrh9xkvCMMCHpdatwelmpMj3eTfHu9hzVp1+Zwqvr3un5Siq7Y5
gVRg/e9yh/JuyJx0AT0B//Jrok095BquxA+HbdBMJjGncYwbZzVJNovqxPVu5ELt
ahJzW/HZDKwctAeHk7SVZglNTF5HA5JOfvcQ8/v2xr2rrSLaOlAgB9vGFe5Ij+qp
Vf+XxNv18wlv9Nk36oj5Pb5/YGgEI7quxfnTHFJ6dBHYl77dxr28SP0NYlx7pVmd
EKgo3R8xmFy3cWXtIg83P3BJnTAuouaydbNwARM6P4EDw+ZVtD3Xwov9Uxbiu3ko
ZEvKWF4qDnewdAUgcaKsHmGrdZjJlTPsBLD/VUm4T5HDYBoZ13hx1YWrqG9PNwRJ
6AOkR0igXJ4Llfn6oH5OkW9FVEserPPSLNnLatzQoDWzHlcv2m3XEsjek8snoDIG
bFQiPUWgMLHoZPIF8g/m+jZ+rLNgelhVr0ZEZ/m0z/C7D52MOlckWCRyKYbw2C50
Gate8BPdz1u9ykzj6WgX9a6Uxv5biwCObRHjhZ7J/4WzNVrFqp46H50/ZBxI7sxq
dxJZGL101MjPow+Vbt2vP9az9qbCX1+pRP7QL8qWgKlNgZNkWiU7ZINwNogBCaEl
XvFsqC3qOzKJH9Q846uabhipGt1uh29dELUG8veCyBDu3afeKIBNejynfxNulaWp
NhnaIN8B84ScOYz9iIXdxKhU4oapUpBKKpk+oRQ67oR5Te7y0VtlcQ4sgh3Ran+Z
CKkumDrCIFrAx5TtQAjkTG16SG9upDsGgY0dRU5fcMMcl53QlyYIZobs9VvHMGYv
SyHlgl+vSSaQh5KXbtEzfZDYxm7sAphJDoOuBCt5G04MbOsAQxfL7kzm0+/nWFI6
vO7F5Gnxfo0cjYM0/a0V1k8MTWF82g2tEX4DbXvHuiJilkZC03WsGVew5BWnpfcO
B8ZbivZNbqvyQvMa8RLTt6395Zy/+rNGPG6wecGzpCbA1tHoSQv4mzxNkBA6EQTB
mgytU2eTRZQQe8rPRLPDamaSKZULNEVaGmCBZCJpqkRQP+vsa8jZwR2eMeC7c+vU
ixfNYbbKqUuk+ycTQoki8apaHwuEPa5pHaM233ERId/kPuw8VGTKlQyP3LgG6Th7
+sAuDGhQ+xnywYj0/UeTCIPjv2kxe9H5jmvg6rIDZ+eaA1Ar5+XFCh/oviSuJCab
QCxTDauIe5XjNGpa2cmMP+3K/Z62JEWS4rx/xzw2sFS9BXbrNGef5xmsX0ytjLzb
pTKATUnI6W5vqVrAxB5ic2w9YV875G76wZquU2z0duvGPhSvHYkXXDrYeMyp1H4g
h9M9PMV/GFxXbBaxaAXpuQnbZ7BDe9ddjeFZn1nTkaxIbYubtafsdOS7Ba1AFpdO
aRRhu/rtlMmEdp9a5/QbD/U/4IDUKUD1nPYwe/T74FR23gzsssa/ZsNKYwnQUA2i
l1U9khxuCJ9KT2gM0u64bqdLAu7fRfdRNAyC8iDs7lVM4HSmbm16bCGYxkOyMXdo
sYt6irg+JghJUodQm2zAvpT2dgLr/jj0AEfL8RhgPdsY70wd5ki3egOBb99apHOz
8HcSmCdAtDsg+jdEQrhvV/LAlKlLFMJo+mBP6C3N0vfzFgEo0MnjtbJ8i3tYNYVK
63PmjVtcVU7Sb4EkS6RKxOFZQp8h+ZXlnm6L57uq+p+2UBibD5H3cGgKTC97DG5d
Tjf3CrFGiT6hT/a+uR5fCRLYXt7Qdmu361IDyr4u0cpV6AB49mw55MK/IE3Loxur
vgB327PYUxOl0tC/d35xSVmdrJ0ufUM2pgSUuyyvZXcNK57fy3WvyEF4x1vDV+X+
pdXW6+zi/KRC9Xc6z2xRhonOJlaVrOnJA+SCQBJBfaUtsOGKSWFKSGEpS984Z2tJ
ftDxFNb1jWrZ0QVSgpj4pGPht928wWHrtCgeZC7syDq7pm8qWTqrnEAZCiigpJeX
MLxIgCzpcYVQn+Ebz9oGM0DtY3tauphmARv/zpMc5ZI49dUABIeWem5yunr/KwaB
GR5I4BqChwfcawFelQhS3kK/aSQW8kbnui6OXVMwkv+nETPTo67CygA8UuvJEVps
vECbyvGqN4NtutIXjctidH8AEfHuoaarMreJgRHbmQHSYFVLmwJedZFtf7oS+BG9
KDfuDVet6cp+92kVn7TCEzayInGpifuX1ZXCG6SiK/hJjD+RvonlDX+MlbUNa/TT
VthrRbpASghtuIbAWnm4ZeGa2wx0uYnlCvVqZhJw37LYVWWIjFkIkYS5JPgc2+vN
jmwcPzcK4NTX2BJ4SibpOBNQQN+uS/W9Df4qsHDc0ibaWz1zUhbmR02xZFxD68W/
LB/FoLqKPNtk4kQTQN1dh3fEh3gY3ZHo430TqtEh1D/6nxqGzXz2Hz2t2DcDHsoI
8Sk8l3zjtnE6ADccOJMdfQ5gXICrRW4eDYp/XWTk9IDmhORIGTTlQ6t77tcf59mL
8HJKbLw96ox48LdiRzp9v2a9PJZfwz7RDt6H3EIfKTfZHZBRX6hWEwyFPHfDNwIq
MHpgKVvhLJDIwi7ZlnSAyZqEU90Y++Zkch03U5tUpdZ9upLlnANapvCVRXWDiXHx
RWbdLJgwofhD59U3BgM2ZnnG3VS7rY/rADXFfIYitLsc7dNnsdnqU3FyOnunY1x3
a4hKOMfNHEb08yzzadCWEATwUdSSHUhuaX/z7y6TzYKHdUEtrA0KDGHkNS7GwS/d
nYj8T3JzN959hLFHsTNpqH3oNOE686bu4eInars7BbuQ7YQf9YgTPJWRuPQH1Gco
3EUyuMhERxRzVa9/RvaouW6FEZFrC/5fWtuy/6pPrQ/TklBtfR9xFGtKS97cysWa
P7MLehYbAYJMTGxxPdSLF6A+63QLxhmoEpDWrNYn+NbNwEPZzYDN1ETE1G8g9KYM
tEqkzrZKwQF75VkotY/y+r9bKYIA72RRPYYouZ1XcNIPgRzWThSkjBNQvQR7br8z
PX0MHXG2zrsxKwmcWceLL3eivMTSWhzJr4KBxIYV82mYYezxKdNZsPQg21y6O/tO
DJWKuV3dqfPg3tNyhaTrQXrS0/wI8ALlKe9ClksT4Fjng6qmFC2wHplanhZOEvje
GDewMWyfNWMM94dVcHD0GDHbeuUJ3ieT0gZsvufk2NsXT0euiyogfoT5zRBxxA7T
T8OOVMrzY/a6fd6oKJZY1V4B+fKq6pRQIrfPqgP3cz9OyYP/5CfWYLg5s0srpr7y
2ssGB5g6709smZQVVfD+sKSstJvJVaBl8+eYWoqurEuteSg/++vHkIZ+9d0RU0Sk
eytqBsYslOkJhfy6bFcsZQIH4lzmqhmT/GYZJ6LUIYnV+UIizEJVgbSdQacvBDHM
GXEXe8cIEOmRGT7WItP+8sIlmpGeGOLe4CLGywExe+dbkhnRKPvwolLS7Tq2UgXW
Rw1gARv/Zj/bX+QD5fC3n4/4Q6CFwv2eF5GSo+lyWa2rPIPkHO8Wcb5toEXg5RqE
o+Uw4Mw40McxSp/24dA9XVIOSnAI1vDJOMke1sbscPQDVFqTK5UCMZ690A5PuF+n
LYO+sro4lzYhqjgIPwvTUwLeCrhkfDi1NGdMhFf1tfabhGFuCwLRTQQ2mfCB6sgW
capIUBjbO9FDz0/DoHI6Z9XGIqzqylyxidhxTcEOlzggsdqXz3/YyGA2I5biKEAg
mqMH4zi3mmreapKVo9nRT9VIzxaLl1eiNOyIiA3c4lrtqxlfVv1a1EFll6/X0Oqx
e01V+yfkOBwU5xtbPO1IJwt/pESikV/Xh9W8UiGIfHJACHlZOquqBJ0PIDvO9qVL
arf5DjYcu2swtARQB43vIKa4NoiuJ+Ko2k1EIxIzr48vGTHQHvJvdetLXN6APx6d
RUIjfj+UmJQ+PIn+BHtFnUxiW5rmuW2rDdD0/8lgcw73A39/AMvNkYFCp9cy3QNL
e53S96ryJROekSQLWe1ZBHu8tfE7IQgqKyeYp6hbXd+DvIg1u9f55pIfEICPjvIK
a3gkvglsZcDI7fDhF9LdFwRCry/FEwaIqqPZNfwfnMCxbijGeApC3BufHl5KHpsX
FubFmWGG4tk4/DBUL81Q1yN+bo88xsvfRR3kX3I6LTx18k7ZxpKteZ7fk68WhBPq
XAZ1a5hoZzG25Lv4JiQP7uoU0wXPAGAnBb2TSPJ1UO0MDga7iNyVVVFRXZFRtD2u
7GQNJomBoZbKEOydio4k7bhJn9PcfNslt8vrO1N91tQMNPPotPk8x7zY+7gZi+W8
2vAlNwt4yQzADOxe//Iol3ht+wBmHSLlItBDwDKKAQGtes4FBSBoOVAVIZlsAu3u
2GkURoNBODG6znkL/K8GR5CGU7eUOTRJCC600etjUpQpypCZ2TBqpO3/0SBpHJFo
J85nXr8qnKAya2zuX2Esxtzt8i02FiJQ4kZsJbKoKXeDxnjY//0Z8JQpwJWFncOL
gLRj0cp/iwFDQym3SQDOLdPgg8Fi5tFHGfBqSYP5rcOq749k92vFJIJZZr1T9fMq
6azSGtEGT+JUn52z1PFWvb/U9dUwOTPR6JL0Hj3g0ho/HRziXWICWDEPmqm0Dguz
p93mPGVc0N6398I8dMCcJ70urbPmF6Xl98V0L2nhc6xdri4cUEL3w4EknLbD50L2
ws9Ur4W0nAV5kKbOaPSh074CJI5lVTd9zQxmaUf3aZQU5GKuddNMwTYsTEPTdqPr
9cLwSVyH5LJaZKoB5BefoPJQj5BYd/zDwWvNOQnVyir5Zz1pFP8OpsRhGKrO0kRm
tN+lG2itLdAIe060+fnkTW7BmzResOaEaml3Lopi/xGH2UV8SX+19z8ZJm5Vnxcy
a8TJ3wf+Ijek2AworWsnfeaoMBGnbaNg2lAdiivyltGUIdchBQPsk2q4EP6O51MT
4WQAZyudQiSTNNDZIBRZF0dHENWnTZYIhuJ9FdTWFvrOWTZmGKGw5rxd7ujQ6EVF
Ft7R9KSRIfI8GQCTx3znYHsJ4AUFc3R8bgyRAv1r1MAdkEWQtV29iTGVtxsIFcvn
GNyLZWm+Xqn+ledbP51aCssCKun0JYcN0zfIPR1WAbnvOlMJqTDLoZWg9limjMTc
xMhkeYMIsLtfd2/wBOcm1uxj283BwUhCt7n7pdYainpq0zAlmoSTHxg3YjqOIDGX
9bi03IufEXUilKeRKu3q8//Q5NJTys0z9hPIdzwmK5ndBHZnzFfJmEsIG2pZNNdZ
jNgihQB49smxXI2hqoy7Nn3jSzTWO0ZMD5DlR7eWtNPh1wnKWFhuZvNk2MSg6nIs
fIR5XQxcK2hRARRhhocCuv0H5p5EUipwxK8JPOuqmvpJWE9pAxWqyHEmTBaTAIhj
EUtuGdg/7nAeCc2X2s46/nlJBUNx81Y5wCKXlN6JGNf+wtPNGObUsko81K8U/FZz
E8XJuT/ZGyJUEg3vjXzBXuTTb1hjCW4BfLS/Ss2iqzTC/a1HDnt7toFFn+I2dbdR
ysAj0a8RS1/ZJMD9o2ezRvp+WNKlmp3CK++ZklBtQJEDq2Grssa61I0h61dazpGr
cWWp8doJumFajCj8MYv90Ytto6f5JDew/c1WNqMRy2jfI2RTzCJZnbnrHIod9cm7
5E8CWyjmfhSJH536uk8zNRwgKzKFTi7PD/8k4nlQQ6FedCtCd02Fxkn2nY+pUNCx
usxxE7By9W/EwFSLBHDNMKX0VqZ8eWWgFoYJrgxZMt0w/WMsoIAVyKhWBs5JCOr0
vkkF0l5OKLxlWJQa/3OM/owXDBqKGywkdvmbPX+znx0oELDogvs6O11IwRsVlONI
0AxcS9jFGECp3j0C+3yCPqKYsM/nalhyBmNbs2JNFw8QDl8qJIOnR+ffARYsLW20
s2ztwXkWToD5ccQuiioTZ5Hi31RfltQfHN1+frDjnhY+488gTrBbdcy0qJ5Pxe8x
ibg3aw3SZee6Pd1REGyRhQC5AZoD0p1aMMIKuc/gFDLDMLvFS96IijrFRgKmX6PX
l3O/0EgvcZ5Jr7aFu7autI/X5lQ2BgFYLcbs3sQZb4ppeMWIVwQ9BV25aKH+OFoJ
cOin9/65t/vNRIPmgJO4/cViW9mQ7sEHhq9d/FmlGyp56UCdVnTnH9mcBox6CQID
tw9dmYXs6cdezUxsxLbgO3dI1QbAkIIwkDDGy/I0LwXUuWdAkZdHmV46PNY/pcYu
VnRi4h7Q00usxE9e6v1cK0a+sUu4gHu0RHHqkn7+hJPiRRltMPKcbUbXuQr/I0gg
rBSz3ZTqnU+Q+MtIGSYDIzDZmyN0fQUSIfXIbijMWni6MMTvHjo6t4PyWMOFTWof
YAa1ibhzbeUN8J7y6JWFZQpuf9Q606hjb/nRL3wA1B7dkUTXuxSBPjFyl6D860kQ
ee6UR9diQJ7UXPVdFCvhtidYq6ycy8drB6vWa79CgJzAfUrsPMJmGcFGPcHfeI23
qarOpD8DJrDpzO4LuJI2YcQnDrsVZTa71iHNQf9wJP86kynMeKb2qTcmwupPEyxl
UsYJijyNBhJ/+HGL4/FEcgbvIf/ssuXC/W6WUdTrZFNmtKnXEyX6LHd4UCtqgNd2
d2wbpV/htaHTo6ZgYVfl1R9ciUawAUlSZEd/eqNYCi7DC+bPc1wifIRvlhO1QhdG
4Bztf+xyy+NqLFOFlzxcbymz/qYFYUs9pzVDt4vEQUDotYVE69oFrsaq3UunG8Al
lXEVKgLJMLkyMWjkvJEY30HjemiXCK8EBl3kE6qDquFlht9VMXTejxObAh4L/riE
xFj+FYV3v2JLgxG7DE3UibRhtcRcuyTxxbgCsUUE7ex7Kgrre4DrgMtM5B4POeEm
Kw3c8f5Vbv8b7hMTCObqO3g85uHSbRh3XmkMy6ejCHQVSGTNeb98aiJIwloyMZQv
1KoO4iVGzpA5rs5QZg0ZtaZxN2nvij7Yz8x2IYYJONCAiLSZi3YtoxBz5FSZqHNF
wrOetw4PzyZiRwFupF2gnZPu8otrkotW7bLyiS5Y7eDSUYTYdS3aTHBsTwxGnnb8
q6XMNbVE5n1vPK30A/WshC344NzsLHiCGAt9ojYX0pod8owGh6EOLcOa/J5o1jsP
teDl+7lxPyVrP6TOVDjPGuQjUIoWjNMGgyKXv9i71gQvPT8zubbx6XoAn3MS51hu
CFJ1pDeBauO6JRLWt67NxeNC1u8k579qQcb9e3VjS8s3eR/iD4a4iiVbG0v7pY0h
dKT+tX3FL6Se6HLcMmPjMLBozrbGBtYvtb7jV7rQNioJXVhts7nlTFUP0S4JGbB0
Hk9zOUjr52q4xFE8Ho//UuigBTJZ9fyaQNycxEPnCbYGgW1cm0yomhfxFxibYf2b
T4+7OsljKZBXS6wLr0Nj8/bAl6US1sEI5uUKuhhtzDP0EecRwh2uYcMILT1Qu/1y
YzktRIYTB+238os4jy3FrOmVKrQTWRG6QzkfuvwW3k9A6MR3ItL/G8QBBpHqdCKC
hwm3KIxe/TH5/Tlv3JLuuMD221kWT/g6CxYmMFnAJJfb9QkV9ZyhXl+F0bnjhDzZ
QSk6EjzzyNQEpyxCF4cwzM8Pl4Ukj4FZcl3XDvdeDTqwucKvA4Sajn2RjuZuhkCV
YcOMh81+MKni2CWgHve5XPanOwXQuDXBJjNYRNCQXT9ne4O4pvE3ynSFm5I0L+eH
Okj9IOiyBUf79lwY41u3uyj1TUDNoNRlpBiLo9XytKc9udswU82fIO7c7VrJgrcl
1wB2Be72bZjwZ3MKK6DqZsWyu8ntac8oaXc44GJT5hXxJxvWwaazm7HxsXUQ9Sf5
ifSh1BFgloc9geDnu7/IvAdiBWH2P1RuVPu173pBAJrRGDn0Qr596eq+GkA4HExy
vW6PKnphlOJ+sBqEDWvqralibKeCcXvT9kosCt13UDuAw4nIiGRii1wy9yYdJ6Hl
o5OPhgg/plrCop/j7JezwD+gOIPuL/PsyRdi3+XR58xrMp74keFvE2RGdCz7CqsO
YjocH+pDgaQauKJULx/vCqrfJewzTbRhJHWWeUKZj+6/gPvNck3+SkQWUkkp1aNj
R4YfFaAqWHuHzvrV/DHJY2bA5ANfxLruwNF5py+Lvl0uxppjgo1YjpgHUGUYqroP
XFhrGOEH8QiA1m6RuIOK2KTe2U8RYrfCg/0/PhoynBT9+Rc7kzmmuaMvo1Pxqnjq
XWn48Gv45vwlflvaHZdrhfAjTv0NbB5qZ2g5Xv6tq41xhJRI3N5oz+PNXkXNqU0l
AQsuClLVObl09UdFrUzloUz9mAQ5pCHRWBXAw3yQFnaLoilAelbrDBtb144K/qae
UXUN4nDtk7a+Ia/QRu9xdKjeLi4Z+p2OWcxriwSsRP/q8IquC9d1dPtOIqcNPZDI
N+CI4r7euJoFpEjrBWbGrk7tQ8/5AEMYptpcMBuBuVvtvtdnqeX8N4qZhhTAbSXa
wIIlI3XKCOVM8qyKcZdCDJnlFe7wlvWWQgafbeOWJdHflRCO42TCXVnmuKVmvPVb
973kjI/Ykv3mWX2j9W4eJ0q7qeL3rAm9mILsAPWu5C3SM5yQzVVYcMsaHIOnyp6E
RP/z+GHf4e8EdnSPuGqtmLb+RUMamqU79oFDx4abTqTFcUBWPKY7/DB4ZAbwJ2t9
2KB333p7k56IndSPhPGPq/TYRK8+5cwjG0qjxwQdHXqoBputaR4fs8Q8SwxC41Oi
induOvibyAfSseTkwEWMx59OVO3q8X/kDbbKD/7gDDOxVr6bNXoD3Sk/74YSd2SW
nSsqsJ7n7Nezf/7VcozV56YUDvz5fl5Yh11+bm6mfsqBJ+V6lUpGyxvPXRX/FqbM
SRY0cQPhujLaXxwww21FiGgmfn3ZZzDIU/Ygx4aX3qH/xW7Wq+3AYG9c7TV953kA
+vBhPZ8lEC84N8El3fXNzizwTBkx8RxPI3fEWPuPnL/NQTnJZutWgm/MGPSU7tqs
daVj6Njcco/PXVtEPc2Z+2cSludlLAMKoYZOs5aWuRIRXjmTCSgQ5jlm3x+JUHl6
atVxQKCbKuLW0SIExgjcsV3sh4GDtxqMt1gm+p8E8Y4rHFwV6yFIDKtpESfXcZ4z
jY8gwSexG8nMlVFCYE7ENqX5q55Io7fPveIgnOJhBNwV1JKe2lJH1XIpx4kVlFzG
/NaGuUQ+VyDEIUspiw0/HDu8VtokqPFNtiRfFTmyAZpCSQ3BrrQZy55JeLY2ipBN
/bR6o0mpKYQV105rj68UvU7L9RU6NnXL+gJYY8KlUzvGR33uCTRZ09IHIjBQJm7J
pADCN6SsWwXk8MY44Qk7MsMs5yG/smFv7+BBb14Q+dWyP0QwCPptJ8yo9h7Os0i+
VFrrsed1RxLkPaxCZDTMNb6Ttlztfciupg5tL1hVvsBcKHYofwYbdulwUoFGnspY
Qcb/QYwLUa0uP56yQIqdWE92ZtPX7rS9DXC+YWi8rIpQX6x8lFGviegPMIGfQVCd
Mig4Rv2+h4Fi6aTjgQXl119uvibi0OFTe4UYxWbiaq0eD35vyUPz0qrLHK1LWbrU
mm/9Q4Kr8eWeC5Zk0nCwJB6shuLcjqYpljguQLgT8jz8S2sFijSBPVq9eGgNelXj
ADA+NDZ8MIH/Yqf/iiXCoedR+j5vpXjX8A3u8DSCbGWN2yeyUFTqUuF6LIxD8saW
JfHTTKnF9PYzaXqA2f6GMDn3IvuqOqX4S6AfJuJWkft23HRtigM87+UpNkE5kxw9
QnmEWqZ3TRk4vI3w8w9vr8SxUwxfBu8IT2gOQHkMcLSwq+nLEHnp9DWHbGjmHF1h
/3AEkQNX/pGl8ujPcGPAbQsTD7yctq+ENW0BUvrVcON9UcNYGZwTtRole0Bw4m1j
c29WuT2mUTiGWKwVnOOxRB+bPGeLLyjpw7yjVDYFSpm7K9FDln1VVP18etC1/RfD
XjIFt+dwpIA4agBEmRP6jbxzM4OVUZtKVIlblhydS7W9A50HxjmDuEqovA4HATNC
zagvG352dOdGuhkDKe/gCHxsw9LUBziDltXpyLk7wsb/Av8g5yqPQ+czo7vkLoZ3
2Tw0o7JuKas1aCaz4IZKAbP0jiP23JWCy0U5iE6LvSnXtBBAdbCkKLedP96Wlpn7
4Q4/amCMhFQcRddkG9vnch2uhgAZMmpB05io1K6lmL4Tf30sIWI8pWRnxfTAELAU
g/+KVOqMJ49ww2gUyxIrUpyGWAfH1L/xba/ATIXIPBEtgiFkHZFSRuJk8Nbf6lnS
mlZfMLY+Q9SL6/PsLV6uw/J6pRpPccgj4m2T2GICGzhCFHsbr9SgK3UsSWZb08Va
MjfhB6WD9BtLP0NeEo1SuoAWXDEf5yH/Y7xDFDiiKUHGQXVy0lNKfbcQwR0PeePi
pafPnON9xDgvHJs9IyWnJ5tqN7C0ggygxQ4ATASMbELT4Rugaf5UGbfiSWMFItGa
qECrhPEgq2L7EB2gZD0YUP/axlOcykf/WudOTrexvSKHXnXtiC/4jd+3Ouvy0bKF
cBNKsQaKGc0S06lOEi61PZrFM4deor2EMHOFvia5aPcr/iH5hS/dd5QHL0HsaLZr
pZIPxOburP6uqphuZdrZYhW6QqpxMnquD+MqjZtWOamk02KwzIHXOMDn+VZroaa7
1l+yE4EfWjsw6Cr1ob2OwsuaCI4mESsPhm524JYB/fR4RiHfDJdssbMSrEr1yIH1
+YWWXkMjxC/PiJj4XPWTQV2eMHrjr8Tj3ORn7o71MPc/+DCe1VscmnawUmy8yP86
Z+qBG+4qce/X02sp7dBcRcbEPfv73R+at0skUpwdDqC6jyInfOBWI1tIGiY493cC
Jy5Y60hBvzbZ/oEvvUn4/+ETHiKdoj3evKGBOEDFDRA+xOxearDJR+aM8FxXrJ5I
sjO2rEJbmj9pWgV7al5aXD4/32bXAzjp9tV8Dn9WiJ/xAe8d/YFWTYVvZhLQTO/y
1lpTGGxv9w12HR/cUXFpCfbaEnMV1XHrDNo+HXmrXuU6rajMQASNVG+Z8mzCJqSp
P9XAgxbc/S83sQPFJ1wd7ksa4ADMD85pqg6ZzT40VyjYpTWmLyBbYkZZWpzoXa45
UsB8GCEf5E11stlT5WlCk3YE4hmfzD4qyuR7hWdRZ9EGELRvGNokYkXG6Deaip2o
dWrJ4Rk6hHD0gtRK5ulbvxRFBShyyjzVh6eTSevKsMgl9J4EGZqup8K8ei/WVm3k
1mdlh3w2t58oHTWVyo3FhVI2ChRwJP+YoVvcH922O3r/3/qQK9BzwINymu4W9Czw
aB7bOEqwCJ/4RtkLk+GW0oLyRxJUkvmtFElCcmSx6KQeUg8z9rQ+4BtudTZxQHrM
Q7tnxSpIxB2gGzkXNSVH4Ao68e9MiH4zEAXIXB6LdyiljurBTGtrmBJ6gzvOfe5j
flrTDGWf7tPfisV0AIG0mJS0YpuJCWL0U0bPEC4vx+d0Z2sDScfJosPBJCd2dABD
+cQc1eoFUfxzoMIzhB3+UoYlkm2emHGgeUUVOBdf9krrDR+EXSGoqwA3+tFsoSQr
xEISeQy5sBqTv0/gHtdLezyHGcZfZThTpLDbNniiGj+JJhq3P27KyDjvPD+pTw6g
LvpqzW9HwxWPGM2xh7eAfZulysFJC/H+qxce0couNgrZCWeF9zezpe+YY4dAB9ag
xlU4qaGwyWtTaml3P48KVHSEuw38UK2+sQtFcDi8f96wLT3ApVTqpamF1xY31CFI
Qw6WvokclgvCJWazPjJ3VgneDXV3oOXPVqBF1SQE5YX2/i7VqrkV2onVkY1usVtd
4pkCx9BP61HGqtSpF48/+SBmJ6bnqnbLtYnVZaS+vXMB3dT6rxfPeFORCfpwE2BE
uikY64/GLhumH+hxyyQ389qh80qmuvD1uEDKmwCDE3kb0h3nhXIoiWRFjFscm0gV
Wi+h4GvQe0o2V0hd1PmG29GdimENMVe1XwMRN9MMgd7wwUaiIAFW4Ed0TENIovrN
8QASq4d1fWlH+/+yl8SeB5vMwgM0I4xVyn41/4xezXBbGMJwxjUlqJ60JMqbHrZ2
RN6jEe3i9D0BxOXoFlIOl4SyrTS9bmes++Oidfh886Y5yXfGMtiClNiUnEev+QL6
WEkMve3rEU7HBM+9MkIzgijIXP1bn8XcdQjrLf4Oolaqb9172VJuTwbt96EZFSiF
BsKNscOM2RouLmpPvUVWfEkR1WV0mu75sddJjTvZko1Cqp6LxRug+XSbHWJhSfUy
MDjM/HTC9QsIObVOWST81YEel1cjTD1SSggBSxXyIqqIEoDkg2ARON4KnaFgfv6j
fxYYPKmKwcHuIv5uBIo4/NJBuT/NiDJjoOs1BeUixJMuqLecmz5pt4oA4vGbPN0U
8Jm4Nz4SIv7ufw2Ji4NqLeaKA0ZA5Olz7QTIMvlmnCrtDz4KG71V75tRAgl6ce64
NvRFs4mYgMFAHeK4b8QCtVemm71IMpG3bHBrF9IwbadQwEaglz+1AABoUqJd4M5G
2XXvix2cNWTLaOC40bac3V/sJkQEw2lVhulXtpcCZK6vAYABZf5FdpQvyaY9BvAS
5tT5e3yTzD3Ft5XMlPCrZWCrKKGIjf8KrpyEuaPLXUaVwemzVYfYF3dtymHM7lfQ
UbB9JJSb2rE1d8E8yg+jAMlPB4Bk3KGHrKORyqdP4yZCt7HIL7zc1b19vr4VtSi1
dWX/RsZrKnpVv6UQnzScXYo0peqQSYBqFrN+0/3y0C4s2Kp/hwg70wDn4Fz4B53t
EBm3tf+JFNbdmGD1J+7LS9rsnF0hH4/ItWWAAIpK8b9RhUCVdP3quCv4+1cU5/mq
BiQCDJBnMd9nOAMbSyaGTDTNKsx3kUfw/AVZ7HG3Qg3VzL58/1AZwfkXeYEsOjua
/5AALxByUt8wDdJyn0uA40Fas2kuyzlqcmbCoJwEZBDxV91qICwNlS4jXdme9OOE
xK+oRdF8xetToMJ6jzHW7RWxU0cLc1wJILIiKbpRpfmCTPsMsh7LKgnBsLVOExiO
ORjztXi9hz4rJZ66MYySxfcANXZkoEEcH2EmTTuHaMpCh2xhMdkvNJp+mY2Fwnm/
UNoMEEWxVdiuPoNb04Yxxp1ai50driM+l+7EYZxOlKQppovaxni/s08neP8N7b3V
O/BVWaVT33Bj0wNuiT8q2quLYPGKjxYLg/Dp9yJI+fcoasazoQ811TFiUm8Usjl2
qr4J9dZmMzQR/uT+WxAUfPfY2N31b0jaHDEv10YSSuKo5gCtBODGGY7kqCziT3hk
9UYaVpyjbrF5ubc3Dkg2Ap+GDo++eTJF0MM/WnZkTbHS2XeFAVTabps9Rlx4kVgv
BYbPpPDK7Gti0nrzFVnhA+2lr+5bPpOx3KcRM2MSNykoOPbTwQ9ChnI2oJtLedbr
aGB/Bn2T8dKtYStW1IFZM3cTBJgVJ+BpRsbWZ6ceOcx/7VcFowoDGXaYTNnR6oVg
7w/oyZST1QcNy1TgBNLYWYa7LYJVpd6B0NTqsUHzuv1tejbH6qMtSWPxGesYP/w3
Nn+5khvPBoUvraGBM3irEzePFPsGjmeW+SAnG9kQDde89bzoZUvo4ibLPoaE/09u
C5OqIKbYBL5Pxskvq2gfUWwJva6eBNzxuGHfL4xcRQ3euloZUUgOfCuTrtmKf7Gn
jIYSNyDhmcmo8kz84+VmdlQ2YHIyY6fOHz18lG/g7/i8zoKNpvjcig9q42EtqEIZ
iWAeQBtpdnBuSKkpLaSHHBh8jIAhbuCuj/TyJi5QyMF0fk+jLJiK4+OQmTdOaVFQ
qWb6MGoxRU6c8xsiC3WQ5aTqjrnM6qmevMQgjUJUtYieMyBoaa8Y6IppMXNThylQ
eFOaR7pgh7FiFpwl6qsh98dmLk5GIeDJtSbX16eC+iFKYPSIgsNk5Ax27YzKcbvt
65ReCWBHpKyc5yXZWnX4eTzaS8oYviIdUOhAGd425ritp9cHSlQ91XCbNL61ReO2
PXh9j2HmYslg/W2Sgw0zWPQX6SvyrZkOTsvlxmrPvRfL/fdQABs2RAEjnHJFLtZh
WUqvM51spz2tf5iPopOaTbEQtMaPFJ7TObKVfxaZPJFO9y+Jf/E+FxCVBzJeZfvk
LoSOtXhcPGNNLZkkCu+FmzYmacY0d3lYIxAZpmdUxDdAsb9I3T7W2MioLsbmE+kA
Cw4ZczPiEPK4txHbuBA5V/SxaZn1Yaj53Gkp+/mQTONdnMjYSvTrAOJ908FWXDui
wpIvgRC9nLp/glAzb4uWAu84GTQEbgSgbygkhWXFsdf7lLAUd0366WnTm2ZXeAU3
8xcEt97HP4p7ajL2MvrrccwQZY6KDu6RyDXPa7efaV+n8WnvTFYv06e8S+Z51Fre
YfTdtEgXT6b2uVkyT7Ez8VFacMvrPXEc7RyTxJG6ZsksCLyvQSgYaFB432ki5u1K
lIMHoghTyPNnLb5LtTLy6uW3/HlAuP8ssoz/zcKC8O3+uD7l383U5IXG1mfmiiJU
XrEPxWtfUxw90h7FXEUA7USOg5gcswtMvHzcaUWVtt3FS8GPQj/8uUO1xRimj/FB
au9KxyedS2+SqKLpRdXcy/0n9xuw3icNBXyxrseeGuL2Io4kNULpGXmNFF/LMhN2
vhTqpmvW2KfGuHCTGKFKQ037IDmNSuVp2Cj8xdPOKmA+d19S7Rx1EE7vbpkC/ZAJ
SpmQgNrzdPqXZNuS0HFxhxBseO4jd4Tn+QvDHlMB0AL5NIdwjKiJvI5mMzLJSe51
Evk/0t9SUWqTMJ6nW7nucXpmDkSrtufX9E483KbUDUn8UFb8e4buGTaTBODiH6ES
VlVQIANTi5VRgbJPYEEEfrFx8p/oP7HMy+c+sSVz3ur8e/i5MvRgtxSjWyTL9+Yq
S3LFyt7Y6Qbnm5f1CW6da7eNH7jZloco9c7m/aqxDc2Z0NFbP3nSR+lT0RE4ak6A
eXkVbfnsb04qRBDuUi3sWjdTaafA5qMhnA6LuCk+ndqQ/ovdJP4fr5GqFxBlkvyd
9eGAyDd3lkgV9Tz9CLIxf4onl92gk5mQ7tNfz0I0ZdSp+8WMAU8D+G2bQNH7j43O
dskc0a9ik9P6PBVbCWTJg2FykO7JNqAekDmqEdl3poB3EULZFwa+1VztFlcl8tL9
hbf6OAc+9jnCH1+XY9v8oAZGi5PUbKIJhSY6snybreAYne+rGjXxHQqFNoLuqcIG
bfFQz5XH0A43xfg0RDcA6c6Cehym9G5Ard9ePcDO/c/nSg73jX4QvtDSCC0zsXB1
STZ5BtHw3rJInWQd1cbtnu/UY8L/0GSD0nTu2bOqziBfxwyYaUDgF7F2rHR0syYr
nATLJJKlsNot+AKTM+i7RjAXApB3T1Q6l2n+EkFSnPiC5L6fhN8UpAD2FdjxddZp
gUkrP+qCTRsb6tuOdu0FwB3Dq4xb8syfxYi+1OPnCyYELl4ezQtHT3k42dABYgBG
T81br1cuBk3nJOdgGVweErCJQFljSgOOeq1b7aZ2sj8z4hWF8SLyh+yTJkUCfeJ0
yYw2xSwieY863h38ARU2BMc6jUISIMv7xEzhaM1E1o+xK6Y7GbdjfUSWd/X8zSx7
Fef3pww3OijbEPY+JsFR1SDNOdVyWbVwaFI3XZUtuhtGzaglbn66AGaxMSGjAnBr
RiEI4l2/St68C59z/oRql/GfLY+Q92WZ9ijyXW3l3oZVAygPT62GnhBPHjeupPY9
iFKrHTiAISlAJ7OjUYyMQGh5kWwhMLhKUejEmG+rLsKmSeh4TIXP/VQdnuk3YJmZ
h9a+XiQ0IWZBS00U+1FJ9NBc6KOZxbpSX6tl0hrCn5DEfxJH5zbnPeDizou5ieZ8
Y0o1AsnX+Gt9kGnrEzbY2nCAEzCYbBtz7FLE5G+j8fF2O591B63vkUKejSuMlDui
lyCxGKsA2DKk79A+OQ9x9G6oZt609FHdBf/1gAoXHUKzE3CARehDIkEHqiFbTGc2
WN2w09itFz46FuapfBtj1R6aq3i+0IQhe7tr/xj53QA2YnncmrJZASWYzPFlH9zc
eGRiO0xCXU57eE3SEY3j6ddzggtF4tpa550eAAKEBEExy55igG723rjWxKevucSz
D760catJIe1x/ymrSKewQrQaRF1UXOd6to0RlSfUhwkmK7h+uIWXnL5gYmbEn8Dv
U100lchZEoD6VHoAQWOCp4oI3p6iUdcm/png6Z9JR9LffwWbeoQK2A5rwLhhKGAy
gDEfLWzIVSMJn0jdVhHTAz5g5XqjugJ4qyiLMN72pq6nrig6lHkR+OpSzh109oht
u8Hh7rw3Gz1AYR/dxoyZWbkJM2vtal7Y+5Ew9wnqZHLyHL+hA3QQnIynORLp9zwt
XlBwFWwS0pGvz3rgnlYyGvfWYELedaNko3Cby5tB6IA++xOTvG6F9uPsiCoOMxfb
/Caydl11BcL4DKywX2k4N29G/5a1Csh1bRF6TL6PZhQIhmuE5EUOKCNR+cfrSq2z
hr9IogPCJjx8+AgAnmCyCERp2pgc+fL0KK+uqiqwND2gsRpH58FOmwLS+y1zKGHl
H+/E32QyVsomh027eyxCCiFdDzJFLEd2PIuBjeqwznz0kqquKCHJQDv6Kbj3ewoO
Mer4Ghs/0QVHYvhEAbWZpsMH7G9JZfwaIaPI3MaHkJ/aZZRONSv5JVKYiPPfr34R
g+ZS+2O9qtuPjZKSBkKWuqro5q+i/sDuSxfoZH5Rd2mwhcKWl80p/ef3fwBX46Sk
OdSjiKj4oxpEdxcmy+l2AQzwWa3iQeEifLCimcJLxRW5YUesK36/wH+aHygialdx
Bp6Y0YLoYfPygpsNNWhPeA8U+BAc/02vqzNudHRIqaAd/AQH9cZRguWceykEr6RQ
euwlQB9n6Ug62DyDeP4AGLaYV8Y8s7dErmyejrcjSPcm/lg4krjkTzpU0RtE/ZZc
KzE276cgmt/ytsGhpmH8Kj5PtpvxapDTJAFgU4hKcNizI3WFa31LxgXhjgM15OOv
E49/8HCtw+nYwhGkeMxmTBvK7SnqGDouLkubbGYonDlhOxak4H6YxKLfakOsBcly
77/Dk+SsRaWcmy8dgJvG4TdeaXeq1FbTzOrUmLrRpgtBNSBzpVm5+S5HvPV9K/79
n7KKoZM3PSLTVH2AxMIO9SrvHsn7vP8Q9Cz3N2vOyAVbH9iiW6PcqDJ932UFIDlW
nHGyOt/efigW9axJckR3GpZLx84fPoA587mS9CxzpYX3wAjR5YipMDo7TMVR1tsZ
cYB01Fjx0+mBd2KKoWalM41Dm2fOebCkJ/EmnDng1IdVWtRfd7Y13Tq0hBZOPPF/
+V4wsj8CSLqtwVGlWYgUa+AplJ+Xeplm/kiwyToZMZkTjRFzcZJYnVLj0lZe/sUk
EWCEy4cHV3h0hkg4rGfs46iAZxRJc5Kul5wMysyj83Q2u40OdVlgYMykFt7ekheo
bgMMuPGHQ3CzJ/XgjX3jLyJoY9K1GJGzofx3uLUJJXjU2KvV5Url8CoOEWgE2VbF
lGrxdrW5e1PxE8THTSN9cVsIzPcXG+HSwVPP+fwJj/ww4mJLMb4T9GJTd8MkSk/g
rnQ+6HbzftSVwbm++0aMnEyvbV2kGidTXer6Yl12cPOLNJUuyhTpT7ioCUDirhBY
+jD3o8DYfhWm6aHKpmVq5GJYNpJGgxNE/Q/sonU8SgS191StnUdT/OUjv8yh1qFM
TKUbqCtLXENcGJSefyGYlYIKO9Iwdf5RsX4Nayao2Y3OE+WJVRACWK32ID4FxgCk
AxRMJTALdGrIfZUeiDIwsqONek+8gZ5QqsyCnE0f4i/x0FbGeR/j4RoBx5Wtc3sA
DYZK9l6e9EIysRMAOEnkKEMkr8fZU+R6MmQOCzVYOdUo4QqxhLiPCjj6KaJJf9RZ
cKl334qhikAfpyQAy1MUg4i5n3+P7QF6FDg1Rf6ucdwKfmkizyHLzccNt5nK5Iw5
E8lYWDCMbLM/q6EdgABqM5aIGqXq1C37wDgidW/X52vjXelVE+Nmd5HbA6uM6u4B
472MkmSVVJ96ApPv4k6RcuLZQ0THdrShvOXrERfHMDNFkDvMmt/c5G6RM9dnJZDX
7CSOaSWeOrXHIxD52qV4C9Yfw4Qx+Rtyd3wHrbSXr6XmUvKe1fvuYrWcEo151Vx2
wsMIXUEhDpfC5uAk+XSOyqdj47u7KXK8BF0qOD5tBCQetIwWm3YyN8iQepqg4eNK
gNASb+koVR3wFauENlPGE8CHmhMoBncVX5QcgC5FKZp8ihwCY3cbdueRUJ6VTlEl
+P2K1dLIaBItjqbtl2MsJ0uc6Qwz7G+Mp3DQw2Gg2rBB/80oy32TK5UepjqDAHot
3YYQp+n75kWid3gHPBrxjGUD4wxJ0yV7PbOxWErfRZfgysXU4YIyM5kIvrc8mabi
TV36Q8/XES6rR+dPMEjsJ5ZUE3B6NK7nTpx+iS4mVfX58TGGDm/Y6imKEdNkB7WS
CigSMKIQnLXrwGZ16cWtqKUousjY9VpD+dV109AvcSdA9qtoM8aeAFB1orjQYPSC
9Jj5t2yX9iqb2Z0g40NcGDNPR+AhiqxE0erZlyIXtirMn0OTGIjpvOubHHr5hIdm
ctIrmQQc5yw8o+1K1kbQ95coQVCHoSYA3QGoEOQKDDMkdax227adAo+3JBg8hP8R
/XnN1StX2i8nG26xLvy5obhpfqyvRVb1sG0hYUhq89NLOmI6TRGasbekFMna1eum
GmCj4UEldssRlsansAfqpWdK3d9CT49VBIfXWlyilAzZZEFmCQ7ByF27F8DRAAkv
cw5UVoA/wVwaqcj/7gWFFg1/kkKLGnNzpJL9S5YO8E49R7rkoz8vc4rd7bokz6Ie
0gndmfvYKdBftnW1HsccBJq0F1WdshGKfggbhCWV+quaLhEEU505Hurs7WrYis1C
5i9BXe7RnpbnqSDW6vGU8yUJMntqHTVoewLcbg1ZWbm9PVYU+47bHzN9l2bmB9zh
Jsmup1a7bYqOk9Iz6XTtQU7zRQv7mujer5bMPAGyUz/6KaGtpQERm8a9oqxsBq2M
1H3TrvydgeDp/Xlx+ep/wMIRJbcIo3JhJsg26aNozov3IE4FpJ4npILJg4uLmJNn
qwYo9ZGLQZEcwKNdEu36cY6v6dX6MNv2hf+LBeM+e+e564lo9+YUkvvO6XEk+ZfC
vKGuq2eKCvuDNrL1vOcV+yf0HAU4eCFPKNK+kaKCmHCOwURuVP4VSjk8rrz9/o0u
Rz8cryzaeSxcl9a34oaA+EpNNpjhKuGpN+QNuAl7KPV+zZgUiozGrR1MEXTGq7jT
6tj/txAbyhL6qM2vLcjCYOUb5Pc5zI2BOReJrcfRQh9LvPTC1R7CqfgN/pibWbW+
rB+jozABMGx1c1LwEPTnSemMT5BxJaYe0O7qsSNJff5ElcF2pemEqlZD/Faese9n
9PFxTxRIfUwAthIZ30RobDNYchrG8MjOdZDBnNjYBmfnq6MP9uXRVq46v2aAr2xp
jTrzKcRo5WVreRoKh7mni5Sa2dhpfAWztjIAY6eK0OO4IvkTr4Mmoc+RH5G8Y8cF
GOujM3Uai8rsx1ERNqDCmaDbSMMwv0Xg3sXrfXol7izqNbsRyUjN+FOKr6LCAnat
gEAOg5HQuygxkCaX7G6mFHPjhbFgsuKMsGBy7jNH8zpQZAGhKuNxlYB1ZIFNUVJo
y1SlBbuvyRpehi/mXmZ+6MtEBCeOMkVI0Jv/hKvvy1jxDjLvuZDWFRhkLduIlaFX
2jRT6qZZel1/r5OwILN2FLMKV/siIkdGfIl5RsRihMzY+q97umpQR1uC4eoCkTG2
BiT+vQRgtlI3uL1bvoZ63p8gzm0ypQHyk2gH5gCqY3Cn0q+3KNpnjsH5DPgevBDZ
gnjGGFCPFMjvifKRHmyqa+hRfTj1vKGj8HDwfKfb9lrS57MBqFRJuKqntbywMH8u
q7z4r+dGi0IK4yzQq/8B6NTdVlUu7vaU+nC2DCOy5bwRCKq+nq+Tx6EyagzRfjLw
OfrXGhQ2KhHKb8KhKaOCFCp2lXQPFAubZdXwQSblBIWX9kQJebbyTsMpPGva+hWM
gTQBwZcA9JV4l2hpxeQErLPMOmcxjiGPLetsFl24e+IOln9AnvhSjTrC5Nd0tudm
OgDso3N4nLyWW0yM75ISvkuuwlxnN3klgw7l9u2E/lsphA4PtNtGK8f5sF/4NTN2
l80rrv7EKgZT+gTWllXtbN0gvCjDRE4+ecUZMNlQ5J6F5nKR5hDfhVjq7Iyaw44K
OLC8mVXLTOVqnJAYNHTRPVx642VwnLWQSuI5Ac6UDldaJBq9YuYnGI24+imb9tvZ
FgY1UP54Dh71zB4LYTVC18HehzkqXeVUwBcsiHJ2AK96kMnS9Vpjrl9NibgwPWXC
ZcHXYbic9D7RJEJNfrm38qNessiFWUfrT5LpTPGV2ZOQ5vqvvTNAwH39M1W9mFoj
qbbPOYxk70UmuN2EdRYyozD5K38PeB3W2hykDT/C+SOayRipNFAfeEm0/I8ejdrg
iM6z/aBFCQZze4G8NYW5GjzUDuKGI5W8IMF3pdnPETxiWVCDD+X+V7LovEMUaMze
1JRa/2JmyTB5eTlr1KWytJy+c1SlvLz4FO+Rm45qFwNX33kJi+xIeDga5NuKdd1G
V//5TH7BuvIrjjU7O3i8LXhj9AaudWSzrY7eaSdcwGQKUyLcvwqx7BmUKxKD5Rp2
lAzfuNn3cm5jpCZeUGdHHYeDjXvdxR0sS+hbyEXmIFBQxoafdnlV22PST6haf/zh
mvzbpQ+WM1kjW52bc+lmqrLHNrJIBQnRvbRw9/T0vn6aVC+7Y2Q1qkTfB92AekcS
xIqO4Q4GUffR148N9OQ30VxNLD//ge+wz4GQVN4TjI5/r8YLb62j5NKj4YktSJEY
usADWXVLk9Ub/v0VCbUu4N9YeMDFbuhP7oxPZ18hpx9nJO8O96xzfl9Dd/DLVgEn
LQpJNZfT1fMlbTnw0CjKnR7SWlRSN0xB7/TsedWPCFKW6/JPQJeU2Tgqfed4UpGq
bh+8QfZozEhRa8/CnJDDHp0wrTShhrVNeAVd3oFizRDOSjYqRjiKwaNzUMI7jOb0
J2YUWN5eKB97DlpSquXVBLXAWB8i0SHnAUrLlsrWhnzaXRV2fgGL1+WutOiSLukf
7RwrUVx4Ilr6o8749I9AeCnTb8THX2CMIjnB5Ubu2uYuadgV+UVZzJ+GGfIOQcid
/b9BbZHr7kiGbKcq4rhYWzN/KT6aIb3hQKm/c4VInw3m/7jTa7N1BSsUxSQtB9v2
qFzNZvO0qQTy/oKynfFzh1EbN6iUR1Bv4Wd9DjJRBLJO34mh+0GRYwYnCQeE191N
tX5Q5GYqdn6J+qgpP2/JH0Tc2jrwYKDLRy18M9fmo3Xf88trRfa+n6P2UzcrEf9T
0Mhl3NGHTEYKAEhRJEFLeI2ruGMaO0yuMckNgRYU9r4MwJMZ8C97UFkVHPc9BZSW
EG3B2Z37NkR97e2sPW9whkkn0PPu5NUzcvP3XLb7ZWxMB9ATc75zLbXKBqaNe3hm
2e6lkHxMIms98GH3pT2wDnL1s8voINFzjB1YjuhofTqAtOme9TOuT0/+Z2WdU6r7
DfwXIuDzbi1CAGmKBKfPsK7pOfxsjY0l6lftbdRYW7nS3giVILzC1iY9nF9abPuv
kFa+AAGid9hjdg/Wc+wVexDJgTQ8xfDvdiXZxwyQARf6rRiqOoolR7LCGS+etZLH
4IgMmzuG8ftZ7o4tcMQOSf1P6uYS1aHWzmsU4vr3xi1m8fO7f/ohugRgx5jYrfZj
8I5f25n88DD5ZcNu7q/3OIKwSLuUIWyUVqU5rBzultWW/ZJ7oOuZdkpg89+7n2aU
NUqwjVNk1g/ANZGn/2kaEXBO9I4ZJoA3kPQqmo13THbqVW73AX0S4T2LjquvhpwC
sK/50nlZi08mDlfLNmcmWWYlFgXpvEear0Aos3gtaeesVgVqLHbjoO6+oSqA5dx4
sJw0zN+N0N2+xxoibfFYH9jQrbiRvlBKKUZElCIYvViKdx1UqoxFNixsqyuOpa/g
s24NLa5VPyA3aHVZxXnTWn1HDsFCRlyh7Th9tRf3iy9XJh4c8wifDDwsnh/LlkI+
+nCviXVDOzDIRixElWVdAWfD5PKWV+1zRcVWXTl0sAdj0Z8STuTN9kUaGKuZHrRf
VSOTLG301BXnSBdIo6jnZ2OjY9AXqfCxD/N3aioHL6Uo1AgYz4cOYfKJ3fRnOrBu
bZbK4qLnqcunegL2ncAHiR16e+7ruTDYbaHrHtzMWz/vx7SqfhFIkoC5HNl/WEcN
1qeHwxSTuLERGlu3mRFspWcvKErjew0WIO3+a+sScr69fgNfaSROWnMqdMe19LMs
/jVz2A4G/IR3yfCaTDwsTLGFCJN3XHVCB5OdLSuOKpT8+wq4xPQPAxbcnRpJoRfH
pAScmCV1dQAtJV0SvS25osecEILsuR8+Byn+rmxQBFTXKq6WA9N3gGkKPhaObnO0
hxfT/NnPepuYHBTUM3MKmWr0B2jMH0cimg2ZCel5Bnte1Cawima9c804cxxWx7TI
hqsr3hVQYHEDk3hUhWoLdu3tEYi1uf9Qkt9+HADC2R2adeidLhNbFFi5uHeK8a7v
19kR5yyfXvWq5gnW9nuhQA84l8ouuQu90bUpDWJbmgYU02QJfvpSEj/C7aMtgvpU
jkI00WH94K7OWicnkFiJHb0dEcmU3dalHOZsRgT4t5stS/TPMY3kKDPPayfCOcbI
wjT5kOKGMzZ78weF03IDNM8iGlsYFdoflpMJNxaCcXm/NYMiXnp+5U1X/BUowOSc
8HjKoY9fFwUqVwP/xmN73zlgt44SGJSfufU5vQGIt/6DL8+/74Yo/7kPuVJa0b/l
3AkN8mumGejg3kG+cEhFPN/WFT5UsqHcKqIMmb+Bgvxx65KDH7NZ/RwCWeJllgkR
pwRHb4S3XKQqJv9QhqfSQPVRbDol5aCk0lBb7tzyTP0urJ+psHmgqOMjO5toL9f5
B3FY6COqsg2PMxxbjURDbJb1eOwhSlQlIG7lDLLcOlC5HA5cL8srOXfgF27677T+
Swz3AEVpCid2JxKFJMFOZamLfYii2fv7s4kjk7cN2tkNkTMo+rIAtoEeCSEViE66
8rd4+2ui8iMjEEUnI+n4j9MgppW2OV7fl6P7/2FsyAlDiu+oO1RzrZEAKxM6FggB
bbvxt3/1ZUi9TlbhJixdettoFlbxtp3q4+mRL3dk81e51qm8en27mKpM7a20ljTU
+piDM9jcnmm4xmmSO7k2Ps16Tir2p2jC7ACmvMFWkDiwhIhhEOK43rI5Mt2UHefN
QwQh1uFWIYeGD4/P4zv/jn8A8uTKMb0dJsCIYzg4dhg4viXTdyph6q3B5ch9MzQZ
1IWUkZWYyEGQ7TZ6YH/a+phcepBHVI2A96t5bpHdt05h6QknGagwrYKp2c87UyDw
OJKVjc5f1YXR/AUxP1hAZ+PEiflh+zJhe84BrzT/3BRXJR/cj8yV4KvBRMnydcey
HEDkR4iJtYvxKsqmC9+QXLAjiyNTBqm3rLOugXZ5Zxp3iMbaydff7A55v+u/xnzk
CQD0o7ZU/QgumHnBT3svsaGisOFnnuAoIgYZ4L6/fZp2+7Kim8WI2Yhf3vyelHDI
0sPsHO+2SaLmkENcBHPtE789JQPpAasQUlG4Eby0k8ZILG8H4Rude+81OaznphY/
GnaH+aG9O0FGIHXVj6PbOpm6WJr0c0gYW4/ONXAZmXuWLf2PAXFYVJx/4l99BhDd
LpqqPIh146JKkSeZ88EaKE8c4bkLgQ1AcxLScjJRlRSYTCN+oo6Ufh4rAew0GQZz
h/Yfn7JLZkvxAOamWbLVNuUuFTLJVoicSGqg/XyyPTKOZR72yVXwsRWr/RUu/bcN
eH9kB6iUDyKGHRcVg1PCNRyHuJAK4xF1+VLZS39ERXkxyzAkorWcE0XRYe1B5evv
tJa3C780vEkc/0y4G7l6kBuAX1RldmmG2jJRrYjE6GQrrxfzzXkGnKHp8eTaE+Hr
Hr6EC77YixdbC6wznEZtEQ8ZAneuMtYF/npAwFL38ZueEF03xDamSq6ya+Vzijzg
7X7FQ63lzTqrMeTJga/nkx1rnZjxrLyGe9Axrl3z2lnEhPmZYH3CtXEa2a5v+rUb
7r5m3fHXQsOv6Pt3VdWIU1MUh58NdSj1Rp6kcY97J3rt8OpqBzDyKMDoYO6rim8K
l2eU4pLkhLlByz7saQm78YtENjmhMR/HACT2LMm2n6cKz0tdodOSAVYGs5Gj5uTU
4Msr/XN8A2MNNqq3KTapGg1PWnG27OlGvyurkgUrMK+uLZJbRbEO5xy6eZ85UN1k
gNeli/QHoVnQbMVYXGruAolNnbk/sicGFJtut+JGqTpdg/8+EEfC5HIGssVYs2nt
UVwtQjn3xVgpqUD9QHcV+vOPueDfW8QRFyApXUFVIqjI00VLahC//drVSwgNJfTf
9EFQ2lAxqC8GKTBf8NiYiJ5ndUnOLWOEt8XENWhNrpk1FlPz/0FURkQ9+AcMXNI3
clFXXud+ri8atuNKuWtD79UT+2hep9wMM3twVp7HC4jGSFVkg93+YNEpx/vm8jRz
W7OTQwSs9PU8fiFBpNEvYo89+vMHW0mGUTWiieiSifaJFbTJkHEAigaZHgNetZ1D
j4dCC94qYk4B5KolptpW/KQJLsXxcb/mRsC6XuoRxYGVX3kXGtU5rpgmOS6CIUmg
ygxCFRQJz3JCH+EhtokP+pMP9Ou5oR6J9XDGTlpWzHBIMxEvm1ObWlrkUyIXEX19
mBJxNOUSoCZ3Ldm1dsWY3DQzYOLoxgJ2SrbpxvNmf0vlYxcRuIwdwdqgzPsqEa6+
UAFVW+8mVyEJ4nC2GYKZ1zcGMCrBPiZpm3dEGy9A+Dzo9Fi2Tz0CZYLh588IZZke
+sC6wNU2XA3yQNDBTjssUwFCMFoEDLheZTGMOXukIzYXORox1TRJ1SZkVPQMg5av
Qu4Zppc5WJitM8u/3qYMJMCcSUapMToA9X1l5zMM2wVH3vEXOvsYl74yeOhvXzNA
OK6rrW03VOqsA3+h9kXaaGmw16p82Q644l5Th4QzbGk6d6+rOfSpQx7I68m2VuwR
06sINYZ4UIq7AVBKdbH7xYfyDckUCFndj56XRIUWkpco6uDbT9/hC7AUCaEmegGC
/QScTEsUcZFMvNSk34iQUX7fHzxxMH35b6GavtrmUZ/YtPNB/VQL+WkN7n0sAqOO
FLdFrciej0Uld7xiRjeqFrIHNEEH5oSDkaAhzGSBVvgc3cng45N6BvxTviS5CZRe
ANXliOLAPsoUqS/2/N4vbPEgrcxY+CqNFp7LtHzN29Yo006fvhWf/kin8nN2l4Iq
sLzXr8wZHVDWVASR56cMV4CKcMWqcWheqSPHFkkqk1XHtF/bu3cuR5CzTq0Z9h2d
lEm7P7pGZLDIPsrLLB6qWDUafLxyjbGLd71GbYGa4H9Gna+79hqeI+61L8I6MEoo
WyJUuD088NV7S2tU8GGj6nQqKc744j7BheNi4N8Zx9WeUxZeB19yoFY9rgNDMhLV
gtF+JBPpb+YLWKpFZiZWzsSsqq6lEJDiJnhD+9ubEz4ES0zzSKttVWZN7qSILL0i
7N0BU1HZr56h9KkjmxdWk4xRY4cQjWJsnd1b/WM0K2RxbUK/zd9TdNLMOUEQbITJ
0dw28gntOGam1bsLcnmVakEbFSgCWJqkEpLYr972lUWufCviQBrofYDyDO8bIse8
RflVJwoALoSsPhVw42kIFV/m2jLKSCAzBAeu6oyF/yfaSj7kvIwAOR+8J+9DJ6my
iur/WM8VYn6M10TJ8O5IzFT/qORl8+62BUX06NPq0mXJsiPvucS6F/UYGVxaRXVU
YX9zNkAgpwx6+xc+/gGQYqEPaLTKcGdFi14QgduSLpUzEZmyD2AC742EJ/lf8fMs
sFcOo6wb5bsZL8Otg2v+mYRyBoA9SUTVu82tktKy9FTC2phYGTXVjZx0JpJulFme
zNAMuMNR3ik/wgok2UP3ADkFSOlqW93yKbdEwLTEm2sRqUoXp8KANNJukdxwimIz
VWFBASSdF7Py1/WKjLEXJ4A2HKWC7W0VYEVeHZSBFpUnzn8VUh4BXUwDpzjWbPP8
WRQg03cR4IX8QtYVD2cVcpaipkQAWy+PHxnTFkT5Sc30EyHonXAdPW0urbgQVRc7
qRg/85jLMX4Yw/4qrqb1H1v7duq/SH5stlTQV8xfGTaJi8qEloLMl1LVNJMdbpKi
WatFh1SFqtDdXQHH8wEwIBrrGb1nYVwA0AJijShTm+1PvAwQH/TrAReCrG6h53dh
3LPUMY3o/DrKBC9ofpJ2CDcNrLVpyvPvWDUFkeZbnv4VsY+OPg+uiICAt+YZb2M5
ovVveeYbCFZrvEmQ41sy2p2349+U8TDjs+ZpT87qoytphyad1m+dN1fhEh8MW8ot
javUNdAH/kzInpUiyd/7uMhWOszXdNm2Jrjx6u+ujEe3PXHz31LcZWVu8+0kFFoJ
0AKQ2vVVyIoq2q33G4TiT/RuQXQEx18EsRRijAE57CdnA5Dt3m0XwEDpTpr+aGgT
76h6n3Ih0dgmVulhj0JcMLK1MpGfp87mXf3Mrw7jXzJMe1Bs17YEBvTN459auK/B
xah5r9ifRh/Obc/yxjVlUE1lJTACojz4EohV+sy/l6HpR3hHO1qB/RtCSNYkT2jJ
W29T7yTPJe6Qms8zGEDo6o6n5sRyhxqKr/p10loIInQutFadDTeyj4Sx3/y7hAXf
2IqFkeyF5sSwBagD51WuxF0y6okJ9znUdLzFa4aj/hdcXeAUdN31hLeV5Oj+eRY5
LoMzfXPUskvA2U/JHPI1DFHIjsqTdud8bLBZZGTgmtP5pnr6gRMx6l0M3Hvuy77f
97bSeg1vTE25wDpcSRBBX3rM/UYCPCkZw/yEER2Gc2hCaAq/YvdB3HQxP9vsf0xk
lVCpBiWeVidZbwlvnsawP+gAQxgenA67Qe2w+ifoxORh0cDCcm06Ml55siv5lknu
yi0SY31ZcgyhmIrIrl0olliRxxoKKruJG0N5ocyDG9rSoRuahHScvPgCxi6tdZJU
x0Oi8b+IfTMgZhW0qrZvKFrs0+x9kfbhHOnarOx0vn2eaq19JWYsp4UC2MkCJglq
a8zeA87/co8E9M/cK3OxbLZ9Z2NuFxlI/q7D99+4TKRpz+AsQ+y2VHUM/lDH+hk1
KIczI2MyB/YNfIP7bbiO4m+CIDkyNNwDUq3+1Tmd9ixk9yQWmeeGKJyr1ESPQUZM
IDKss1MJzRCpPv2HVc+3kKCJ9Uuut5ioB6BmVESejO1UlyiB8mFueDTMRZjRpqKz
xX9t3aeMzydy93avFxPbTOwiEBeF7O030xLTCA6hxUqgW+9rLdM/NVPuX6Dn0uDK
FREwrl4wX2zEp4Yr9X4N6ViJ2/Jq8uoj2QntuS+E0dgRNWd0IPxd5nP/qghpIHyj
C3c2n2t20TfQilIXY7V+7uvlGjLhll2dndxfpoqG4a87Q1AWztGD/hgGtY3Hr05P
e/wFBCEYQ6JHaltiVCWq2ty5F0Uh1sc3f98YvLDEuVSVZ9GwXu28zAQIL4esalxW
ngkgW9KzZDeF7On7ibs90+O+J4gHifof1U91ZRK3NB6OhmlbuNNDtZlLi39QjItd
4jfkafgYqnuDUdN6glWgrHfzb6G9bkfBPTLabfjg024VrIaioA80TunyFpe3AZ6+
7f55t5wFoB3NkoWgGuwqQIaupnKaOTXXPeETSnbCi2oiW2kZ5pJnJ76A1mNesoWl
PF8pj6xZDICnSOEVGAxqk4L9ocwZ/6BNvSP2ovBn9t+ztOSLqRSf13qu+BrXseaV
v9bdSBYkJLHXco26auO6H1GZDv6niZytG1jjDH/tEf3v4t5v9x3Wp2tvQZBoyO//
Y3M/+7QO81stgpHCylEzDXXY5Wtxo/o3mZeqCc9+RdplqN7/Jts3LJy9VYADWZYx
Sj3xwVRDy1biVEcefK0AS62P3S/nIyf0TTLLBYdLTacQ9P51qz1dfKz8IdwPGl5f
ucMJbuk3bG80i+ThZ2hdz6DPIkMkjOb+EwbqOlioi972RqijMjwDDA+vgsHau17c
+GhN4qCM0m3UWdkI/+zToOElsNVUDmN9HFWe66L+H7xD2MB2AfeFSUPbGFfl6UwG
mCB/R+WqR1+kuY3tjvg4hKNRbLVrasauPROsoWEb6Ixk8jVxBY32JOSRbuLT1dg8
jnJFGzqZPIBhPt6a2dksPP1OblWUzVkxTNY0z7cirDb8F6NMB9Dt/c+TyhiE2Mxr
67EGkLqx+8UVu4neiNbflQoSYeiF3dBqMI5z7sPGXvkYuUzLV/bNdmAYYRw+Eua8
T57nuY4nXUMJDfTCDDjsIsVi3gDDAmu4fE1g+KbB5D8uVl5Kgsdr4Anv6VCp/qZ9
wNo2J3XT2IuDA7KHWfJBd9l30jGsLKrlJeztaAaYOqwIopuKxvVznP66kSGhMDBQ
zlpd/X3PSIryviiTLV8KlYEapUxvtM9RM8anLCNKGaQc2bqWTO6TCvCWX3i4S3eY
lsED7qn4Er6tHX11yvsp5PsNKBESk8lGHtTZ8x5gG2ldVqza6Zfg1EsX8xSHmtsV
GqJ3BQqZO/TWpN0kPgqq+Mv+ROfo6PYVSXTcRZNlNEIckfDaHQWwhbmNEcpbsCsW
tnKQfDXGWUO6Qtq6J2w3BRrSOpgVdz+THTb4jxidEfiz7RvOOZ+wl9KLe+nvseZy
Kf+FAJ4aX635LvUfCf7/25fT2rnOmeZYwSglyYXh1GxtyX2ryZoud+OH9eliaGlz
cFpKmVIf1u4FtTOanHi6ewqtElMSnD+1GiyitJMApZAKbA+bHzgNj7aA56TGSp5z
lJi6NyJ3+5e9ruCE4Ep4Hw/bNz2SkZ5FlkCgl7zhZtuCLtIww6MZGJQ070YeHaRB
eHJJn4plyBEHJUXQ7kTM+Af2OBxYZYJx1fNt+AkqlcN4YmmaTHgTRZQAU3xyw5p3
ey/M8WibHJvQqGR1w6eZPfzeWI2A9tyfZb/Ul83I6P1789za3ZyukLXrskee5Tt0
V4jWLD5C8E5GgE06DkN5BRv4fvLe0B85TJKUSIhnlDmGjNiY6IkHB1nfsMcjnjrY
dfFd92KO38V9wwFigK3wJZBIytZ9HkEo6d90S3qcVgg5rgMcAmqSFzNTj42rxrJ/
Ga3SKcahLIpXuKKr8ofedRVOXS51CA7sYUp7/7eZZc3aeRPk2DSb4so+9an6+rag
qQJ3kJLpmLmyOlAuiW2VDvHsk6dpbxEFZO7UWX7adnCOCRO0fW9etgVUJpB87c/+
WA+he53AhiHMgOKdnOrrgu6Pm9CL5m0yVidFF9P9593cu17pE9Yoqeh/321cqm06
SW1xb4IBewvvbj3GrxBxveAiYysP/Q8uqK5nMkpZM0b0BL72t799qsJJGsd8TrSO
ZqEwwmwut8EDNZ1n77EWxw1CWLu3YiINBBaqzfqHLgcd20yekd9FZL814mR0snw1
7JnNaov3HEYjH7Vy0jdOD2oD4DQ4OgD3kbPLa8MebF5J698P709jmWQLCPJG5z6e
0DR5gEaQe+QZZyuBfRgy+qVQMLlntuyrFJY08ft1tMxpBhCLkXgaxafix2cou849
yJ9AKxPHrAIy9TKDTsVUrwm4Y5OBXfbSKJnhi6kyDmGTlOLA1f5MgT0dT98mF60z
+uloxoYV/l43YVEWlZl1kxfH4qnoX5mb9pT4UMXtPxtWxpqN17cBe1OvSS++t1oQ
IAE1T7O9U9hVdna6geysGXLF6Qt5l4NMcVddUhyTa1vvaqstYrjM4cPt6C39gYJ3
25O5gy3XQ3zgNSA3OGV3PxYqr8KY3wx8S/0Wbbp/e5dJuM816iy1uI9S+upva3Jb
T8krtoN8iNB9tgYKAoTsK2mMqjk0flUnb5Sn1K8vh4wzPFq+3fqBvTeQqvyw0wJ1
z8+EXA0R+Xs1jR2NYkGraUkp8DNQX/eQ3eXzqJktD9O6ZX+37vVxaD4Ngw3/P+Fb
/+EmTNmNR+2VAMU4cwmSl5hxujDD4MHapl9PENecPZi2hQkoNmIbb729gxJRUtGs
ObgaYuI6hfY+bkV23VGehUQMgmdXWYhWHs63q1vPe9hDc44aLct9U7C3sqEOAIXf
IVtEFxRIR+DG5pdatKVZRCYVsUbzBy2q4CNvND7cW4Yiszo2Do/8XSAcUM6X52sY
QUjFW9WEWdxYEJXbyxl7DuRBwvtIxVpGJiMYLUvoyePubqR61Ji8e0XsYzHygw/U
TxpbtXK8OHXX/GbTVK1DTooQNwFzI6I+GGhSTWhPJ3ZKnuSRxpWUUXgLYCk2YsVf
gs9o8D1RIaigwqWP/Qf11xsJdH2dA/zAlovMDxaPu/UJeDdspQemI62qGfg+F5IR
qhq2fh+GxxbJ3rnxixAmNlWTKfQpC1vClElT7IlhSpHzvsj+xbYNqbB0WDm6YuNw
7N5fOJgiylhvKQ4OIhJWWFzaQy7WWUn7UYRCWBMhinXycF1z20NVg1lKNmTVB972
lfI6YhiXEbCnq1ImnWe9i4z2kQE7+WZAyg3OEFo3651w5SQVrB8tH13YmnYTNHNq
dftxYYbsl1hEAh6lSG+ThypB1DcF4aO2VCPotCiCBgzNCJD1JWHkFxy3cn6Es86g
4R5+1b0lPl3R8/m9Gy0Ue0SiIV1YXM9KtIHbtsQoxYh57PtrtTFF3KX1fJi+9i1N
Gs7kcHfzkiq0KemtraZ9maVsBZNq9bmWZQOVmKX/k0V/08XDlWgRIkBovuADadSB
laLMes4wyRtkgPiyIslg1g8CZGfTayOT9lCNFNuqiByOTiej1D3VjDWY/INX9Jd7
23uQ/T3ucGHY3xIkQ4jXNmyhXvmA/tJPn+gtaC+vrHwIGCZFiSzyIav2pOiWBb+5
3Bg6sirXCUQnGZtduesIQhassI8T6yyXmKuVvZsNI0t/NEMJv3EFobRqhHR/OT6T
i3hnT+04qxpEvo6BCocUwDYob0Noo8rH/D9Qv+TUiH7k14JMGszl2YTJg3YQtWDx
4UiYYsKczPXFRDzKCd5yoEcxFB+CMKE7waUb6QjysU41xpVzVNF9Bym7z87QQeCR
CcnUP6J/wXEIOhg94xZI+IPmygmPE+u+wJb9aWyE78PF5nmAvcCJXPqWCs/s8f3C
xsTzW9WMrKGQQZbZ62H630545QyC4t22tCfeFsEHgZ8Qynlyzf22HBaL2P+giLKi
cOWOozMrcwG64bz8NvvpU43N0SRA0BQEGWpA3FH/m2d641zvtdpUWmVd3WdBBkUN
1vZcszTlzH5zq9m+YtBMY8wdYANc9W7P+ZNB7vgyin6VOe4MAN84+owYSX8b9JVK
2cNQsm6GAjYMAroOlplKnfzrvdrZDQCzEa2eOQR5ahSM13dBQps/qxSWpPMSmEjH
Wex7wBdr51yP4b/krnF2qFNNf7XyY7B/+42TkujRsRlOUa2So6YKSSk4irn7Ymp1
2sEeGUzF3JdN/fC2ku+IYTYI9OjynndXOjEQSNpRmRZMCvz6UPke5PtvfRaDg5Hn
oRBnXZzKybgtQHUfbJXWwN2dn6b4wC4vkXkz0k3kEcsxusJBctPX8zU0jnDM9HSe
nPbfNKuD9LSJ8GCJdbSJCJwEdXwHkL3vQW98d67EJhD8boGfwL5oGzDrSheSVNoZ
KotzdWIl0+9GSK/dE3W0FkwcGpgnCZ5tyzjmotdeepRkKaR+IpbIUsxEFrkaYBNn
XQoLmj0QKxhpej10+jOxXVJaHRQZcmQM1dD3sa90pq5+w7OxZ3oehSbf7y7tMq0P
KkBjr0MkqIH3QE12L4pSmEhR1IxylI9qN9ujA56XbwUEbdOB5C3u7DVmgAgrSPpv
sAFoKzOE8EN8vVnQutsbsoJKsmlu+QV5QHCSe65wMrYX6Nqp50Md1t/s3/aXz42r
wENjL4a3ybbdpX82mq8+tY/eZHRRkN6L/M8vVvyoHJSOBo+ZhBDskonhCHcKEJDt
8ENiwRUSYsEMPjQM/gVRbVY7PAUaEzj4adYeChs1s5zzU54kaX/Z0RFEaK2WXz0J
/Pqc0XQjrFdI5WYBqT/z4GlIWSI/1HzeUdqBFvdagqrZ2dKUzkaFIKUlBEuuv6fW
eLgt4u74KNPbrfpcv8G1F3Eh9u60s/CwtFn5SXwsnMqAx3xi1s0B7CltbYui+mif
BiOROaK9QGXLlO75Uv0gXjNMrxeoGDJhBNqg0BTPjD16BRZDBWd21A0XTiu5lR/p
0wH5qfhZAiIp5zCjqNBGroJxEbf45aqfvI18KdX2fCkqz6VtRDOwyXGSzjENpc1U
+EeqhHqtiLkJB+IOyUa4epAd+VerFh+QMbDb5AZ8BYcWMjBgTW0Z9NwhoAUC34jC
1nIj1dV43XVUjmmga+BLzRozAS4ZzWXypbh0chKtEdzEuUfPxRsleDQtiKyNtOUS
sPkregUHX3zbrXKapFM11C3moDeYrl8Rs+z9ZoVGvHJl078LjAVWUbyFCssR5OIs
sAyKbt6/P9HdvU8YgMc/QjRPqHl7KgH3T0M8H6V64MOkE06fN2Qysh0IORhAG9OS
ifdYz7uUvtVL4STdReox9SB2e73CWjeQeAneLJZkRkvYtVitpUC94ze2NDJzQzVR
UN9xanJammgiqQg/vLj+xzUsaIfoSa2nXFOyrcpq2LTHGTGRvRsK9mFa6xVNvJK4
St/fh6BUfAUcm/Jd45GnZ1jAAjPTpvXIE3vdVt7N7GV9PTMIe2kBAdsyir19L6W0
6CLPcAfODYRNKJMHsLBJaOJtOHQoimNNbSdggv0OvMThQaYFI8lGmVXCvmG5+zMz
kmkMALY6DPq/A+OoxKxbo/IdNedTFLTrGal5VVo19fBq7WABxJOgdJsS1HGa8ZVF
0aeaPyjQKyCLEq2qR2O9okXjnA0+LjtwOevDylzkkETDylqiqwV/REcAdGk3pIb+
TwuL4E0dfrczx7x2wAuS5FNcJEwFVvC0G/x5eSN6OXscM5tCBqeV8dUmfScYZSMO
FuPDNOwRZvRIYbtl4nEf5SM0fwqIE/fqWTtFEv3gBbCBo+vBFSLeSvqU5zy+lBdK
NbPJp4Ifm+EAY9JydQye1PBxc2BdpDFeRmNNjS5hSRKkXVR5+0dKBKJsANZfR7Fp
5eRERR/zlv9OwWaemADYpDHGiXjgTXzqdfUtSWlkFAHcGNHTN1dJPsEJ+hfihsHD
z6yzgKbUmp5o/5LTc9oELycLpm3W4vg8oLpCSNXkPoje0E6VdwyIq6iO5NV4YMau
KeOeUcjm9dE4RFcT7BVdcFh38XlmdXcD6Gkeh3paemSudFzJHNZKJF38j2nLqoH3
CLrVIbBvdFHB/QtBkVtBQnfm+ZzNno+J3R4wu1mIpzU8UyFXTcpog/KA8rFrSfc7
O3qnvRwZS9nuFxHB01P1I5mrDxRd7dcRGZ+ZExN/fG6Gle98jbpWGjsL5M/5W19n
Z9DBPlAwaBa6YmAK4Xtcc+OZu3DQ1FinSFkvR3nMzzI3Ll9+LFFrJ6uk3B8ceFyZ
+7neT+glmykmlN/FlEP2IRIno6HPSXu6pJfXF8FNVvnWFAT85EgDEaYHR3dyNptZ
ebpNXrK2TuH+2q0sM1qKS0okPPeBTWaXocq7luEGrDHutGQdhSHujC294WMIZfEQ
minQitJi+LdPsft6N/3q4yokhF1X7Aj0ktAcAwwUUG7dALVyGYde0RDO8Ljio+e9
qZT8r3Hd08KTzPK6e+82hFDjnA7yeqLtFDAlN2x6sUEitZj4DRk/GKZUtqsNJxzT
2hiSj+yX4zQqrzGA9LDVDUNqAGw2mEWwxwxciAG1G0N5391ceVE9CPt/zlAl2KgD
zXLbF3P83eh0OU3YR6gfalC5JitMuKTZcziKkMj2+XMishUUCmI8sNZ6022QG4ZZ
Ozgkjl5cFB/tfg2wwTecs4VpniC18swnEzh7+7dxVE+NSFezIsKfJgxxHiPNdxYH
+BvLnUxj2d87oQ4HmP+lsnm+4hPkWmX44q3U34Q3DTJ8mYu1WI3tB85ewKzM9qp3
hfmgQgbUunPTp9Z2EGvnzAFBn7hR0526dCOCJFAGLnZ5FxN+E6F+P+lnrdh1PeZj
Qm8BxR/+RRh2RyCvKh23ee/5ITKt91weAU7RUbV0Sqminwmp2KKCFO5cnzSWl4Oq
FFeX4fd6uLUBzpqVDdg+G4wYjbF3t4v/mdnRtFgtYA0RVk/p21kcPcH26xJsdNan
JqL2Ei4WacJP8DoUc5W2lFaFc6wJzA3x+UufFsWvKnAIVmlNigVGizPhn5HfgC8m
Zzn2EKlJzBk3JfpJgZhFxK0DlU5AGFx5cFG/4+dLuojry1TnO7xEqZVSgUr8sUIG
GVrwZDcdgUUoOM3vpMZKt7ppCN72e/cKO4P7MI1L1iXIq1R1IeU2D6sjIW7K0SIM
tZHG5MGoIhNbBsal/0G62Uks15X57Hd/NjYel2FAXfdBuG8TX2qc3cQf0dSgrGZi
QDNV/NlHrExiCCKMc3H7TGQtgwrMpJu9anoRs1HpSFoj8Lx1ZEiy7meaKRj9BKLD
CgQPwI/7hCDOwVeCXe/KbqQiyBrk9UPAbJNMlI24E0sQRW5jAkkpadam7Ck5K5nI
cZPlM/9+PGjkcJYH5qxTbnP73x0jSs4XBxffG31w8fPDZoiCy+77QsEvSp2j6E7D
AHD12w2B/mvYP47CC/qWtehEFG7yqbGSgHJAStw0gZKxz3hNM9uXjU8fYOugF4e/
QVGNnb355YEwDccmpPkpQMycca8JdrBkUZIqDMje/2JVSy89jgRZOHM3e+t4oMIj
mngqtfYK7lqHAn9/3dwqk6Sq/++9bi6rKWu5diX5dy11j0xxhySNBEmdtzD2C+6P
ENXja/j4jhuEJJFwvuFSHjDzonEhSNupbb46zYc8wbiizGS0oz13nUzlofJffKxA
Df50Ci+f6odk8yle4mM5KxD5l3g+qskr4tiJqXt2uVSm3PjxSfzBgOYVyBiQ1NxD
lWqtjYDzabQ2kvvAnJ6RMnsMuojfpo+FseZJQ4GitBuxcn0m1IIAvKqxcJexUF6k
W7uZmHI6BBZtzN9C8LURU5uLB4D7IALowBqNzQht9K8glaIBQAQvAsFxSTpWBooT
4FHRdAaDT3J7jeJxhnz4OCEiotmMM/ZUTryE85/EAsiusWZ4ziyCK/ZAP09UGlEC
AEq1nl8m7j6BtBmYXr/A8Npeo7KcCDyph3zc5ApOCrfAUPtWOavaOhh9p/qOQr3v
eRJyeEudS7dYm+ahRGmhPvo6jvBoihm7ReyXp2sV1JcXNnfN5vxo7gWAMJA1gC3N
n/CwPo+NyEXaqJ/BOdgAZohXNBhH28RPqJNzymoTr1/qxKYBHGfOEx7T6sEGPPlr
altbRgSE1ncxt/47rGkWzCSYrw0iSlaao0ZcTjElG9u6ZGpqdaIgyktSZ4xpK8e3
878T6bs3IDO/xxv3LWvTCgfVMePwj9dYhs9Q0g3vhNp50dBZdxDEs3A+pddH9uhL
X58hwWSfG8KATl5FpAbmeoXJucn7GSBwThnbE5oSZ74GCizbpXEFzRc9GehgdgOi
K/BUyIBbz8C7FDtMCp4qowlV1PVqWtod1WzBEXyGmsNCIlafJaRgh+IyzyNSxAEn
w6nqihZLXoPM/8PRy9mW82bT6jYaRQ+cEGGGgeptHZvnjlDj89H1vd3WXWnq7B4W
zYnHnlLgIJSHXgiHuMkBiawOCoOA9+pIl0PMRuxObYD1/ym0VDdWlkKU7072hUVa
/DvGuJ+AkbYY/QqNz2mE16RyhZGEIigCy/h1nhkUcZZNeGxgKl6EJZm7W0Ms1GAg
sQ5AE/9w3ck/f5nlgJBYle5z5wEeEUNN31ohnE4siyQNxxMRpnIethuwC8kmKOgu
NHopLE/3tGiB+rSwOZ+CQXFZDxG4NDoBD0Edng1Ei2u/Px6tR2UyuQnLl/hafeGg
LfzmyPXOPTK/lt5UrhiIraKGUtdipJmzHZkqd80BGff7EwJiXJSwfK9JXWHPLIWH
GMwmYD52ffxAOHVAmcAWzgPECUay8Ga52Bmmf1WeEZilpOXTiMGfuFPMFwHsqtBe
cGMu1744QB05pPRgczYgWZkWellS/0EuWLb7TE5b7RZY/d5eK221EsQlcNaxj3PG
b1/mRGX4oV1SY/xwSrh70l0/LeC4mDQjrQ4w/JpaIxdPuzqVQbBI3+ECvbWVoSvz
9CginCQUE/XODu3Q7Sd2+eeG32MDZrg+Viy3Wk5ScSomgrQOi17555FZGcUagrlA
dE6hc2RAUxjuo23iqETiLnCnmXxA6YyPiq+BIQ9D54rfSJQK9h5G96iYckvk3x5a
nZnLUB8SSm3I8Ys44tNPUX4TFnpnHxAANBX8xWkUBvhZjLTFdBwaIJYRSNJVsUOJ
SS6QdpbMvBPJG02+XoC1Afk+++QgAPueokVj579+YJ1DweQvI0jT1jmLqVmXnykV
rBVLkQX69BPm+WePhHGRVN39LZHhHjDyBDDGcg5E/43mbcrWIsWnuQBBjkzW71Y/
HRAL/lm/0wTbv6BE2v2p4juCUqijx2KwjKwb/Rt9rlJCV/rRqnYXmZ5iVJBplIp+
y383VwglyE3DyQeiff8rYgTuViDJ/rbocFedH0kbZeL2uMntBxZnUtOgLc+pQyWV
C7jLoE5izRlDOdf0uObjeoYleATInWFpW3VYBS9/RaZGtgYNAnWF45r25+kCpdYQ
4W9gMhUzZz76d9v+B0xfldtCKhDKwDhA1QASuwe2zppGMd0INu7koXJb4MEMEOFE
fw3CL6GJyXt1T3CPGW4PwZj9xhk7hJ0YLnyxix2MRW9ZnDZT+E+nN73cKbq+P9Wi
azF734pNLX85hwqLZ9nET+SpEcYR2fwkHKrMaV4a5+sxilSlyIbDJpeS/B3QdFSd
vk4vsH6GP89p6CJ9AKFKvlGpcU4Grx7rqhFy8oDXDI/T/wlOk7BLfyCaKiLpGFIJ
6vc1iBHLVKYlzvoEYL79yE1i/LbNG/D9oe7xM8LhUA6vgMyA3o8F/DYSaDPcNW5k
D3ucv+P5pluIPwPsC+actV+o1mPNw/e4zj2lpTDtqxDV4ngRbIFNKn4VJyvATB2H
g1MvUlyn0iU9gyKif13Q+wqj0bA5YsnlFj3vZeqjtdzJI/vg5UdQQl3mlu3UJBzv
HXbnmFafwgUj6rs2qtMZr0+OiSLlktnYzRrJGE+Q4aSkOzCuWR1Nt4mPzUvUK3Lj
NYimo/XNBV3Cx7WiW3NTGFnRbaT07KMiCpXJbafsJeE/QARkTHiZ3jYEdGcaW9Ry
cVUp3MmxZDYy3gsvEQIDW7z4ghDM4aRihdXMObC17Rn5g73s09K2BfjCw2LtV5VF
8I7mgHSu1UMxzBTQSvdgTvum73+2unmTwJPzyW5JYKnk3h0oALzYYbQETU6pYYgB
pEzCiDfnMInHy1aIEn+9mQEN9CrPTJ3s+XvKhfSLaZxz+Y0lDeLxehm/Tx27wSg+
V7K/psHh9ng9dTPobfg4g+yhDlemC+FDCbXG/5JTrWsFZxej5OcPX0f02vH2h0Kt
hqos7AGly/pLHP97000HehkEfk/YB0Ljk+lW/4dJcKL540Ch71PBfzCMax1eS4iu
PLKclSgLQFRBspauhfsDdis+H2OCvcx3DQplgU3dMCRmIhLr1R3mKdevyFhvyobQ
R8XAl4IsKcuRxhrWNkfiTFDOwLHM4JIecG/ARsP42WKEfXrxeXv/AVv+rvztqGgh
xJLS2rhrMmDQGoSz/pclHMwEce59+F1r1i5prekGoNhj+IwAPNAPec8pmLM5h1Xu
F9MAvmeLWPzGLiCYn6jF3VPSw7+UYusKk/khwmtj+Z78r4vlQnfTPCzdSIMNfV8X
p4NhYlnNdlSz6kTgQ/gT6BCLxt6ju97RW7J2B4asdTeUUTwMKB0gkoTC7YmsYgXq
X9rKNsIZBc/iz8ZOM0MxcD05+eHnLVFaMFvKu6IfoiU9Uxg4Y6mHf1/GTj3qMYPJ
EOkN0mL7/56JcczQz58cq7nkT+AsH7H9qWyOHd95/SwkyhQ/518WA1fZEqYWA32O
ezo9s/mYv75KAzYKHTlUkDU7PZLKo7ldUh0nxl/5JObisMsJB/MPNMHIfRo9Kdkc
4k8NDrCm/l9wdWIhJqyK3FtSKEZOMJEEreTzTssimvKeg3xToYhNfstxTNYiMNx6
fOMlOsTcmLnt4e3KPclcb3b3YdPgO4kHPQd7RUqPBr9VrtsNEnbnKaCjQHq6XXpj
vEasF6vDCCWHhMsxuvMdRYk/+zsF8PLcwKKkyXlEtc6CTMRns3/f7m7FKdR6jwUd
o/aer6URU7rSYAl7TIWZ4wK9uOut0b7l/B7YeWYeRzxgex6ddx9jhmkWxhb68fWn
ROcvCMRfHhEE8wR6dk8uNVxwy10rAJI0aVBQhIOk47RfzyjKTX0PfyPF5Jlxg29C
XtCrSrj+6zmXVFFXxT40lF8tj4HMSarGsC5xoAljRtpqee8qd9Qs0U+LLgjEUPTX
tqeghdSpWD5BGMEOS8o2jj2K66AWupA6wTcv+Q5Ozg4h0hMk+fAtakEQsS01gs1+
6EKkTQVTXmy5KgEHSI25vVN+zPPu9le5Vbwo9AAviN60kr9cKKqSNmxq5CBGF3Xd
bTEPfbOrPtAVmeXaQUxYolq/LFb1fXy7dA2JFWOlMNv2lS0nal8g3jvX3WryHS0Q
PoEuPjaCcR9QAwTe/ac35uQFkgIAoGaBEJB4X6u8j1PLYAS7KF7Jc5bdblI6Op4X
+q6ruodd4F9l4oE4gErfFO19wmz6N2MDRkYohToU+ol4ZxfEQd3bjlKm/ayAnOKB
dFh+WBRt9g/E6JsCsV21swPu2FqkWjhaWscdtZ4+uF2kkfL+jg1OZIPV0yJVNpWc
xJWyOXzCKSFoi0qaZQBOQ+YZHIC988Pg6zs9NFgjBn3tHdIx29fov0LokLvROlks
08wVXmSLfzzO+GkmWa1jXYYs6rUYTAQ9oZIIsgwJYFWgc/fHHsoEeRRDshMqVlKY
+jnUZjzk1lp62OhqGfkv3+YJSZ6zKUx96aaqDoGIriay2vU8tEBZKjoNsWUwa+7G
CuDBbjOWf1aWCBMfR0cxqlKldSL23Fd+yY89Kko6hENDgxwBF+Gwyi3IUd6mlIQC
OiOb7A7DpQ0ykMBiRqlGkkQsCJ0Td1mZZb8g98Q/hE4Ml8Kb+lttzV3xsYQu8/j6
XSLNdnYde7J7zyDqYLIHS990E6KciGrvw+hrp4m3T8qb347vn46I9OuPiwCTBbuL
+DBqADqaPW4NesjONVttvJAVEHN0nY0YwegEZlb6xOWGxyReulUgY9HrqecZV4xD
go75nBLDSdujQleCu53Bi4yQ26UgCUUBDvKr+pbcNgZDgSaGp+2GBsZR//Xqc92D
LXCDMKdmOL/qqlZudIj5koL0MAwAHt25toiIQpFiel1CaTp0C/cO/HaTmYjoE+1f
MVwizY2liv4/3EmqvUwuNsAdLpbNLTbzaBdbmhFaETJPZHnKCXw9diSGo5Xv3VUO
oWmSP3jsvICWCKufxxR72Af2Uk0iZav3iqNyopsP+rI1brxEGQ+riTkaR8wbBQD0
w3S1ogV4uwIIJdazTldHIucOTZW5eUcm+GPgm4EnYF4dq1ilrIcrc485xeicNyT+
`pragma protect end_protected
