// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
pPCdT5JSK5q4RZfI6PViTtjjcEIMZ50nX//OW9VIMVyR5+vSzNnKT/3H1a9kERqZspSq3iWkpi62
Km3WpAqdJaYhvwiY+F3rilpNSXzUaTldGkbYchvifCLgULHC4r+3hGpVR7SRsdb/Z5Tr6+/atg9n
Ac17XovYoDdN0Pgl/qjcZ+Ny2fEKmXl7jqkIkIv8i1M+FswlK4qKulbdqCXQXYI9Xb4zZlKAEg1c
yeniVBRHK1xieKUqZkBpi/PxuHbMI2oegAQi5D0qcGirie50VlK7ILRyOGnQMJb+uQisUQLGTY0V
bQvfnMWp3iaeluT9X3Lo4kPKFAAOsF9nJX7W+w==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
/yWl7nK6liDok9geCiXFjBr5jxfkpVcTOMxgRP2gDyS0F8ct6QGDXtADP666tjwWACUrSi14aoRl
LFLaM5m+B/tnF6o59cfBzH/wcSAxk0UJ/8DteIH6d+dohzUjYhmZ0rRhzLqlKheP8V8/SK+BiAym
EQ8t8Szt+9Yiqj4JuVZat7cOg3QMZX2oMNPJWgY8lMtA18EQ8YJiIreEcYTKtftfpTDl70lu2w6W
mW/RpCN0RiSsgMUjaMIcQHvesqWwFCje2VoGEY9JJaTs7jDBCscvrZ7d9Fsuk+B+OvXzfvqSkdh6
VipqTYQsvnaqSNEDAIZtZo/HjQviZwp01WiaDhPWev3XxnaTg5A10mjoR7ehXVNDAE4+B9tatyTf
G1RL1BGJ9JMa1ecy+39F3EiepAICbIda5A+z4MC4CPVkXUAnX36OWdNrdplMoK6hNrsi43cAmra+
RZgXFWtTDv7Eg+gDNzgqG8ydqWR00y16kfTHwcaXXSZIsMWhpkQNrgBiGRQW4F/u5KEA1hCwkNC1
Bm+FQf6KIoRG20AK2G4gwIr2yR5/VfBmgmVC7JrFV+b5NxkqXYIR1oSc3s+Z7S3F8SPwTv925sRh
JAHZk37sxZxexVmwZP3ef1godghm1s+CTSClbc+hND0dJiNEzZIGmThzPKBmiKicmMHvUJnlSpga
f0uvq22nZOkLOiybDJ4f3bV7DnlTnInfXnVL+suvjCJiVKVYoRHgmXtYM3DK09cf0hMH463s+wwj
ldD+R25xRORAziE+mbcl6+z7r7EZj3JYCQc5+s3YYZKifkbK3vAWmCzRsbyrXpp42qaPHTVvmARE
qhfUd3/TJUZTeIiNz8miXCgXsvHMO4nE3gT6KQ63c7YwcibkCR+uQ4r/4tOXUmheM+Y73IOxW1e4
vMkuCYI//cAlWc0dy4UyW2mg/5S+wxrVwPcgrnde3nzfDHsQrviMOhuzge+GoxBRnyBGLr71ZXOI
NGYxxBVUrewkgdevNEWEJ1LbBXTWc6ZBMvhUot912YuMx1WXnSXGE062p4HW5Lp1KsEztp9SxzSc
z/Md5AMbW6T8ktZgmqXL4vM5xmTCjNN8SCIeOQ4aUXwykRvudWTToLg+DbmxCwb+NxyidrL2e2sm
pqqqcTW9M5ghmiaM9/ny4g7s0yz8yGM2l0unFIFXakCLiFRp5w9B/kIHuktjeCd+UgQxRs10+r2E
vLop7UuXBfIXF//25h1lQkdZddfsGd3HFFH1qgtogxFoYn7cPCKO7WXMdE/9eooXMPWaMUudsZNm
M7V0arp5dWHqCFtEl6cWAy7s1+AK1QAEI2EvAAch5jlMf8LaWi+FXQWyqrXW0vySoH6V24eTwOc8
zExfjKlQ2+2ZSz7EPBLiTcfiJJ9Rox6b+h8hzvM+OszzmXxHIIbZQ+Zp0eAP3qTsY/lfh6sZOOjX
3ziRmhSyx3OcHZ3o/csdLkOOV9UwH8mZ4KYbtdLddZFW2jexYsgrN2w6vOuLgHR3gBCRg5YCA3U7
gc4jx7yVArYD2iGG8NkPWgR6MHjzpv2Q1JlpJ1QcQNmoZJyJTIctWua6PDeh1hWF17PoBmVXAR29
L73E/qTBvrt26hLjeq98bWOTje6iXOIYtHgZnDEKAtNJpiwtKESRcmmOTECGOt/sOGakGEzHlBSm
omT4VzsKMBB5tKh9KHHUdbmm6/JYGr9SKkMjKLHhs6uPnlUtXLiaIc9sH2gUap9v4HIbPVYiwl5z
memOypKjiBAhCSE9UMVO2Xtnyu0W2tYsZ/B13l+5Lbe7bOwkxO06H1AVv0H3FNEEJiYLmS2wjAO9
Db6DdGFFQjCaOnnvYlpoLAvwocLyopY6yUWecJDwyN2AEhM89Uwb6dU5t025pu+Akog1DwBXdPHN
s1CL8r+Mix+mzSgrdekCGM8kt3vHG5PQxuv0D8iCQa+NdprynbHXb/M3SkdiN2LXNLMwQ0qa8P2i
wlBxmgi3x8VhHIvYgvLvy2KTVDvtxOWxxzwHs5XuKn/O2zsSZ7+87379CBQu8jjGa+phIyH0//W3
lazhhJIolLivGZ68Vt6uncmv5CfrUxMzrq2GeXPFasUMIwg4nT8SM53+mqgpAPU3yly98Yov8RJM
xKct9PnNL1oMP6LrD7uW3NxBH+KYKyuqLQapwDcOOPqik4WKyqF/g9Pgcui/NSUssdlBHtGCx3F9
t58rd7cJQe0hN7X+5tTwnOMDOncNbyCJt+aKHp45cbh7xYYCMQxSXbRxYfD7qWvxT0czu4ZxMV1m
IRM7veeLj+/f7h1tKan04KwEEHEjK7TypAQ9+gJC8Ew01Vj7GMvHfVak6Tq92egmgSBK32/h1RQP
cE48EcKYpKvVkhfVlwv0nxZIyNnaewuKJOrwMCqPaNFosxADxDO0Iw6FzgZl4aSdwIuOszH06Ocs
Nzjvw4+1UkTpRcIZSOErzSDS8J6loRWQU7ClK8c4F50/VOAh7ST6k6ykr0uoBn+0wGfoCX8AdNv7
qfxOjjZcXjCyIjB6bfYagajyN8lJStyzM3TRK7A855EiYFCdhXXFKNLp/JfIj7l9FWR71DSfAK+c
b0Wc4qusMLnx4zHzyx5JHjEfXR6g8QbNZ2QjIzp5zZ49AW7uj/uFGwVx0dzomUR3eOnOzMZdcwmb
ykgrk71cFmlaX+fqoAJkIy3KXikm3z9t3aV4OqyrfykrdSQ4xPhcE1R5XL0wkJijTl4cg4QRPDA6
ccKpDQRRFJJf5JwOtkXYvTE3iFrIWe9EGKjjpykDPyYZN4O8c3tpArsmElvA4n+UOpib+lCghtmp
bJEqMkSRxAFiVqy+991Eu/ZuNR5U9UWDoQLNfw8pc+WGKiOspQLibhH25GkCS/vvMRaNcmAxoCDT
hJ1atJlYxEbbRlC6ThMBD7yqGB6zax8LkjT53fOaSdIT5lekTDRcA4EtV57qCR5UsJiXsutxPkTH
9KV9nh4LEFC2svTzOqt8W1yDIw6NSPZ1v0l7RYL+AbGv1SgThewF0MAuR5+/Y/BDkNzBeEYulXeV
x0BjfRoTwj+LVkWwKtInOEMT+qNG50KrH+IOcoh1dpyBW99MnTJ5AdnkFM8RTY/Gknc+tV0xyxcx
2qbLH0QZIv8VQ9HDRP+6+qdSWaoDEgRlvKGQFXE2WOfxoiLl14VJvlEm3AOhI6x/dxz/fjJ7WDS+
jpPXWdm1+b9/mjmw6N1VUB3XVxnc9kpBILkkBX8cf2GLE5V1vbsfh5DexXTZ8H6G/YJGnjL1Osvp
qR98eAvO4EZ85+Z4CZHMsymZzYL6f/MhSS9PTH68HkDms6Kevy5maHiYOn3BvMndjDpfQSuGhnmu
/V8nE3JT205rSfD8p2qhuPjzYFVg167AtaIkTgUUjA0XTdYgN2y+hnjeBPmaHTgFS7GigPHxjFVV
Iyi3uI2Ra5AI4dsZgKj2xxKn5Mjsu1qiuTsmWOuPUvz63eG8vDpLxEpRfsrXi31ZNLgVeaopyCFs
N6eU3NBCQuHq8guLSgR6ZinJboMiAHdqBmTjDlHZ2+sGeuFOkqmMJVxt4H+TpgQf8XR5usO3w93q
+cThosYrbBiEvPq/luhVChbyJO2NwiNHDoBDPZhZ5YAND1CLj7cokkwUaD/87XKtHBiwbJCgBVEB
tzdS2lYiuJQC5EHM6my6u6OuXvyggX7E9kCv1NVuPj1CVq+T3RxD+egWzv/rrVT0DvD1caopl+YG
JkDq2MPs0/HGUaOw1bOYvKX/b36PzhbUg4Cgl2+mH9dytefiBPpm+VxA5ihJLLU/aqu7pIjcWmOc
1h8oxg4fFU5qdBwr1/5WD88COrJ7xEVLT9hC5RLQDV3fl1iiup0NHXEiU/nPWIR20WmvsYrAneIN
VtqGmW6Qd4Ta452pAeQsN3NHO993/BmffywnQH5d3pP7vwY++wIzYvtXX0NrLPIOIup07vfaBwbz
XAOX2OG39gSJdzEFrWq2l1ZBdarIKtf6/Exn81E5bWbp086/LhX0WLABsEnejoMSsj5GuP2g+WZS
v7344b61l9Huridvidb4gRZ1aj7C0WlncoVWYlfGuZRaXYcwoKzdGoZBcx8Np+lsfIxrmkRQs1BH
mdRWCIM2BA304VMwNe28Ql4H6xGQhuyalzSFl0oRWqjK08+b0Qq+rnhCd2NKN1GpB1yDHPR5iO1v
7NLTLCoBWnCGWcwr8uCXoC9kq6NbHmFGPbnbqt8OBIj2czBJt7HidGqZCCYZNlKedIwRFqsyja+K
IpusrCy//qvd0G1Da0zwq9/p7hXhva8oigvWrOl+99kJL0EVSFNIBOQh11ERJbctDf7Kqzmu7Zex
FudxAIkcICCmFWSUdIVLCn0dUTeYQJY46UOZi2eL+IRMv5nfzjfK9SKiyr8wvOb1ebSCOtCRcsp8
m1x58udEaapMcEN2Pncd3V97GtlpVfjgO7OxOy9PDTqCRvDRVvBSD+DK5DgDHrRS9ab2Um7a0Y0J
C5y/ra86gKwHZy9V5zigFoqTmuWouQH0C1GrrDkNMAwEkeuVtobaBHD7YMaTqtOk0GFNs+f7nefx
/ft/yXBrRyfqllyYeL3nRISehVHgaVu7C1Ojoiw0N/cEIitEiVoYLNgAEx+qNoCOAEInWpq20WGM
PcHo4T434zNJjtNYPb5fGb/ybpRMtBySV96CjQRiZsE7sQz/j7sSyA/OABd81jRi8RlcS5VDsWCS
UKKHFbg5Rr2DEOE2tDjjlp4YGzQLYrnQl8Wj4rOlcxM9smFPQcucdmXeUNTch/kXbqoCWdGP5krF
P1SkcFBQ2oI/C2PlCmg3hYlPoPUMfD3ADbTkmD1Rzrp2AYlritptcd5FFIPB3n5BApzZTLP9fMM3
hv40ZUI4o4HkmyH2eoxaN2yXeo4HL/DVEGQq/qMDOOtX4RbVRqN7ykLbJr0MPOc+WX5GgPQi6wg8
bh+xmdYIqOhtBY6NVCO+h+cHC8yFxTS9lmjIlHU8bVDmyaCvpYT/fRvLcqfF+0yzhfq71RAz2e3k
PD8xUyqEaCam8Fr33Er6LFaqm6CHZCTN3U/4NAExJydEkjikTsaG6u/ds8JhF8AcEw75jHTpMSa3
/RwNdeA4Mhqje0pJQ5XywxXJOclFpSMDihgOnhV3/a/TzyqXCkLoVs5dy1lZxsVCFcaEjxLT2Sqh
/E2ReFVvw3Lbtah1qtCD0GHdLTYZIJxr2ymSyW/Ww872MkXPzxBYRJvijW/8k3KWdDfjJT2wWJ7Y
67ZkT7oThG3bgWqPr62pWYOqwN30JOIUZ7REiv+B+hMjmWjpxlY2qwlQvvSkXmDo0WnMn34IpU2g
IiPVSSIMfPh2MV4wUZgguBpIsRqntTYOQbJyZbSRRuezs3L9RKz38xhsotM7yobYX8ldCl16pLFc
o66Nm0IAr3zZZiiep5cM4QndtJ0V0dKvudUziVuilAydwg8VgyQaEvvTYIUAwCqQq5Xz8Y4aRUER
bHX4IgDbAY4+ucMk/8dk0LyGLmWOTDnhF/dQn6jpqMgHfGgDn9fTqgEUP0lqTMtL03szImB4cq05
2cHmMsZSeVMeHMTqpZ6KXft8ItdYfu4bGYdh8t8ZIcwjgRRvGyAGcjgAhDMhMigPJVM7j2rcR2EY
UpIRYLcbymuQYuPYTmhHeZWNmeMIVmSzPv1FVJg8PKfm4yAnIacXoTE4dAFCXrW2W0WiSO8mwjXU
RH0QbJ0l4zAGFUWJy9YzO6sDQhm4zKWrsQ/OyBsp94PciHxba6rns1KlbSv/Xi7lF3wJwGTelXCr
FH5KTcF7ssFF6EWOJrIbZIJt6pq63nXbp/3vdSlCt8TLmivCxYqWW4k1n2YLwDAqjW2Fbh8mJJfD
7V52tqFd8DW0zQmHSCCakwI1ZK6Jeb+yKNFVzfUKYzAUlHUSZFJMt0jAosXse/Vxc3t+Mn22HvCL
F7O0PRI4zGIvIYysgADM+ZlBFKh0cuIMgsjXh6nUO0kDqw0KZrCCkRPCd/6I71XEw2P9SdE90DHC
xAinCJHa4+CyeoxqMQ0QP36NuXoRyJGEoiRGYSiVhsvXIhMcYKeE/tN7aOu5/u3WGbLCmBHPmbJ9
PJD5jWij1qL2A/RtGWH/63hq8qMpQnQ/6yofnKTICUId/lUk+MyJ6MwTDMdkwWcDQqbvF9TKKC7Z
k6V8ZXypWK+sBOryMs5zwjcwOYx8u/48HMjYm24PSzHrsCSFRWKTVon2BrVIbeus9VM6x1MaOIu/
KA6WpHttx8XtNdvXaNMzQh4Lj3mGnyGFiG1unVlPRejMBAgc3Act1/RmXkGJ+Z4ub46OvNPoGGRD
4d9ldacdFF5RQN6ZFXdRmBW5ZDjHzcxjDzVtQ4FV830NfEDPM5ybTlcsw7lsqvfRMYFsPyQnNX2p
XHG9+OfNxBvZ/cqRNU8wWwhzTt5Kpl/H/8lq7EkkktouDoqtnVmhUmN2BY90YSeLVT54mX3B9reg
LgWwVzUguKuoHjmcfFq0hCBY4RMK/9naQTFIdfyJ7ZXfP8f8jyihZ0EdowrNglxktGxK/iinnm77
2L+61ifRS8OhuWjY/bQOd1/KB1ln/c+dYB6XpPQXq59iPn2e2Y8KgyY2GHlwc8LjqUfrPyZeT27r
50LrAac8tE3A8p2Z5FGxVcOACOXbd2L+tKGaR06RyN+CitVwS0YYaOU6r3FIoFPJuIQODfnJt3p0
gZFqCpPBqTYfO/LbKpU00urKjBHnapGTfjaj2H1HMU0h0bW1RVodgBgZQSWMb6y6JptiUpRhewkf
+Sij8/XQnOYh+vATHMTkLcGkU2S9W+QavypeYKvEzl9/hws2X21qHGytMP98ShWrKR6uDAp6i7GE
+DKgr/G5tbzKyTbH9q7z5LRaBG8sRkjlgp1HIVCxp3wIFfjz+20kg44gI34F7MrLtNUKvYNs3gtX
z5wUQG+Iv0TAczEenkKp52KUEeubHjqk5TFkxgA7HPA5Seux9EGyaj4NmlnArY9QvpsyE8LZLWQJ
AictIezlb5zBpv559OWVjB61XvN8CFV+uP+o/wv+tkEhNizQDE9eO1NcNyzDJnJX5QsUIHmyipLl
1Wg0jjPPpRh7Eb+GLY2+mLkeqeHYMxkvDhoIHGSdbv8z5mHFQBzDBs4gsDtKJARZIunNGNIUJ8EY
Uh8fZPdPHajW6U6maTGEVAzf7anyccElwcbv7E6C6C0hIGAppAKBt3X6r4uDZYxNhqf3Oz8rUejP
GsyNH9yP+Ud28pi4a75ePcWhgs581jVwYUwR3hDf/teUc89G0iocAYsEzNSy+Dl2j7958wr7WEqc
tLDCZnsUhvjo/apS7hKBCo17caZLjW2DQLCCWL3JArDOS5+TgDD0nF341taNArRhmXn5JHLAhLSR
IPMhYvAYkLn7CnDQ2DzmJxh83wbVldnCs/d73Orl+O8HfyRqFiIop51jcDEPqZSNiB1QXmovFs9M
y64kh0mXq1H2Woa7K0PSTqB6V+l1Po89STzjBV2+AppvRrxwgKN6BxFsE9VZyoBfJNvYoKDtS3JD
fOXmDhovnMmYC9jeDPU+fCP3DNxTM56o5ikZNpZ8j+i5sOjiJntG9jZxyTQd9zFrtD7JlI7Kngl9
5GIgAWdEZG29gv44bWop1047G42/jG2s1J9bUgP/dmNvtxTyr/f2x1TX4wTfmukn79Q9D4qrvdoc
u6VmM64SE0bnLG11TbdWcy2nI2u/0aMcZG44/UdhXSgwCgQq2UFaQOo4DZdFAAp6bUI6xwccYvjR
6ULQzuedOAR361knstyNBUWWZkYSy9+XNjy22DfRbYFlDBnhbIhCRbzI5YrPUT+5hFmVPx/Z/xSW
DshL5XHcwUHKAmspbZfuro4GJGo2CWIhcbXxQSUyDrhg7ewU1U1AExYY53aT3HaNXRJkboTJUzIh
qrvjQI5Xmu62tc58pVVXBgDydxdhk0J9PYDeGp4oy8H2pk7Lhz+q2h4Div/CwwjfmKleq9m3MlOq
D6lGNx8N2dDWl5S0SyRg0L50Ox+foGkkOC5ugGTHB75cBfTjdLjbWZYdLypDZhH3o0f7RjU57DGL
9TueeLFBUdf2nxWJG6DDoqEFGQCJdXENsmxcRHiKmhtvycCIHG6+fFaGJXFvV0ngSHsiTBRBfM5O
DuyiCzARZJfjN1Qcw1mySBG/sSdw8mccQJqTuQOVo7Om0Te4Sg+ibeVFTNslhvOtvHNRytU0aE1w
SwGoWIB2h6pnfTui3hDpavUUoM4NkJqdb9YEHY85Rb1NGwePdeNqg4RcSuDoQK//p5c1Jd9326OR
thm1cKl2dDpAzBqguRwSIFxvgguMooNTdwTTHP3NIgJeZcXaMWOZkHU/LRyEdLtHR7s2vt/laP1z
jeI9LjFZrZlq6xe4uP85KqSZjfAG+Pz86yvUu6FDnC25nV08aUhW/8+OgPlVwfkaC7E1niLrYtMl
+wfXXsWy1GTUa0jaFSy4wfDOD1IoFwC+6VZrQkR/5iwQgVY+Cvc1DQytMxDZJ2mHoYWjGDB1ouuw
k5AoJggjc69mppc/BI655tjqJR9J5t8vSyb/MgW/qxccmnadobSpRkb7sDXiqmXBOnAgcoIIQtJJ
13RHhEm0zzTYtVPnCIOvNoTPAAtCP0o8EpINfFULCxIQX/iv9tp6J2HeEOtjlJ0T+ncm93FT4Dl1
0nlVCmlhrerfUUgiKdZvDkaZF7VAQ6b/NssdbEpqHILLJxPR6af3BkFJQE/dI3u28imsa4K3vm8V
4ECyZOR6wyhr6loWPgLmOWrKjWdvpObjApWkATCjvTWZWV3WeaTDq+TLCfX+qM5Vl+9E79FFjC1C
4kWKUHuIPt4TpLD40myHVB8nnznz5BRdcWlvzMvZ7Ef1FGEiyzacnEb4pg7/fia4zKwrSRW8L5Ri
3FmpMaNcm5dMW7p/F7xgsd7Rp8X+URkqKyeIqnEEXsdhczWSJMWGfcL3WA3HogK5D0yvrHq4V3Hl
efMTiPTLhLBLeRyjHu3SWu+CHO7U+4vyfeC6gMNTuGGAepD54I0sX3mYbhSU8JfkU2THpAWHw+lz
QiFfoQUbswCfnhaA4E44mPhipJc1vT95hDivWKXIQtAzM9/q/Gk7iR43MpxeKeoDG4tmV2DQ5x/i
JIWfP5wF0tsTNpc13kdr6QqMNkS55sPh4R/KqfgJ1nh2ENPamNePX9bm9a/FHcywGZDrYG/DrW/O
lyXdg/oLoqloN7HoztU9Ficp5yigbhZOVP3eFOlJdBc/1RPUzxxKl9BXN+Ib3Wy+rPTPXR7om25f
KfLwOuu4nobC0YsppsDDFrw0yX78KDqXuTpka65QeiTRMvpYrdhS5dYZ8ZGei+Yk1F07ZEkctHVE
Aq+VV3J0N6aVZ236nadBRbqmPqpzFqRBC7ttI+3Nbt2aqmb2zv2vLrTuPpHwY4WZnsaocQx08fwy
TaBNONHSVgmtP+QNP45Dy5Fc4qNPp2qK9jGhAmHQEcwnXocuN4pD0fBz63FpQpe9QLO1hlmmBK7T
g7eKIjE/75pvqzqguT7UQNqThtoXbPhNfoetphRd/qHr7R3slgh1jDtHAiCqS3cAysBP+pAuI5uw
8c8TvZO0ZzZ1KtUbtd9ndYN9j1KdeEsVOSSUvECjDsLB+Vlwhs/WEVSPJumZVk7uyl8d8cURUELv
rCz/3ake3SCCvxxXafx24wAeFt7xCoYTKzbvgLiJr3flcw4jPwmBxzUtOe/CY9BsmrABvVHRMiFK
vbl8WlLEior1MRQr6B1DW8nLJLCLCbs/4ZtYsj5d5IpF/kTKA98ZmFTacqUYTH5OVM61FQwzwPHi
F1H01aV2benUsmDKfYvvfDqUVfx7fox3i2lOyOB/lVS0Pdzk6a/GIFJKjIlZl96zy8vQJmf9ll/r
Ing85gmvgYXm+UNCh0t7GfJULSqU1XDb8FWllhgsFz08WTFDotL2y0LcH0oiZPrRCr5I21EfMoQX
oTUztY3lY5LOrqHLuVhZNfJYJC5jOhpJOSk+uj6VGcVP+xjwyDS3K6KW+aZXaBWWaS5WfIA66iNs
CHIG8b5GFyJzMby1GfSx1fzkxHyWGY3enULIYQu0tx6KQuDoNJXg9a9xHVxhBn2TSzSjUvIJsPgR
QL0tMWXWOQQaCCHRpJY7t3ha07sA6zilOkJx6q59F3ZtTBm5k75Ztcd40FhnIT4pO6Nv8f/WbITi
C/No4h2mydb2v8vsNdjkmIotVtuix/WwA3vYYgxV6jCpGgGwWwM7TM2rjBdgEmx5qMpJ3TFCjRlw
i/xBR1ai/mhr+Sxty6uQXNctlV5XTSAv6wshnOswXBIoNTeyG3POo+2cgjAFj6CqwzLVSmZbrYvl
b9y1t3q50V/gk/nYZw0zluihxxT0de8H69RFk68622nf2m72p6OvwEP1TYIBU5eIFbXg/vVaPYOz
H0NmtAr4JfdiMFjnnk+wkeFxgklcXyX2wQvR0t1G8LQ1xKPZr+KjWFmIZpLYlKa51/r2lILpGgMq
rYQ+/7BLN+MZ0IIGb2SfFl6hRL+OqkSpkIDSP9TkPoUWAUCWG7VLNzyvKqHrxRBFNd5THAcB0WWZ
aa0nTWYcjb5wvh6pUCS2PZbldUjbjkUFXPitlH8rzloggghp3KrRNNEv6bHdGIl7YQrSPg9x5NoS
Yw7pI133e/miaF6ULyLjhcRnKHh75eE4d0ri7Ae5Q3krI/d80CZfmkeE0X2LhqUr7KEXq9MLoBa4
VB4ui65g4mLVT1LyvqpZH4bAhTkGjuXEJwmTiU/iEMG07/3c0cCxPobmDOUlQqW8mGmXoHQN86CP
0UOtyMrCbKwBmNV1v5shOKenHbCaObfXq2Yq8jmxuxUX/OaEPSTHtU0edZW5q7ncRXXjYgwt9VjS
QluQzUjWE4UDb1A5ytGGtekwjniV6xt7ncz6o51peu6bOljrPCd9+2IxYUPuD00Ryop6xjAAhUjS
iD1M9p1H0GL6CmTx7CVGwfK7fWyrSFzyD5B/Ei3E8zGRl0D0Z2R9CO9ueeVG48F9iElIC1l1itZp
zSCS4O+ZiupncBKlPS76gW4FCTcTTix6FZ0aTqwqwbWPpMDupoo7QjUyDFmEZ7HAI+XM5qjVDDmh
zO/goBBcnlSB0Fq+BZfV5C4/j0ONTTaaSl5vPOMc2hRYHK0oz8f0PZba8V5f9IfZyVoqDciEVJZA
29gTHzqCgMmNGAltoAJJQU6VqycUpdpZjQp4rtaX7DeFj+tQFThzZtgVT9MtWPj1Jg1wuIQ1pWef
3jAqFDr26Vf21W4lklOAc9QLpqIToAMWBpUOXUIB/s/irQ5x1onaWUIZ9m/KsDdmun1p9kTUmvmf
BVOZhOWan7ij1FfD5kfHLJSpbIv55cYBdCNeRMK6foPsH11zXgr6lsOdXrS7uJdykScQjrwPDPAa
jVJfZ+emkOOeULxGugaSsumOpdWxJ8+MyJ2gdZip/xGzjfOnQQqgWMsM9jJuwIhLjOjuVFJLnRbR
z1T1TeACiueNRAU/IuSTwg6Jx3tMRgY59L1KmSByJYsmCUWqELInW6L1fHPK3dIXYDa/+PA9Cj6t
nHyt2smlm3XcIHOczlDAk8ehZv5w18xDdVMKusW2yA2Z/zVqJ6hCyUI+QjOF216GJN4r5/4MnLRm
EaOUzGYALcpt1hlhQ8CNpXmPTz16v2ZJMABQ77fsBPQ9RS9FJgc51ikZtm3oMPybnP2bX9RfE8a3
GW9CEVDf2Tsxwn148juEYk1XZkZj7cTb3+aF+gEqKfAgtM8OBOpFgdt9ipvGC0dBA1/a+67FsBHm
BhlPeGQwZUkxJdkeaBJk43ppWw5CT98I45U0BO7ceGBgwPhPnfBvu+hq9mHSX+tkHQf91DydOpZ/
pOdSNWCyzWLl0Sk6cXMSLlq3H5QaZ2FVVk46vc+IM/CgCIKroUdt597RyJouR0iE/R14Zkj49uWi
cHjaA0XcloHrcVTcp+63TCJkdL3bH2IaWJut142w6OZFZA6b1nk342QzuPdOWrz2qZuXvwJrfywi
HoY2WRlU/SAGlp0tJmbYcjidrOTpgC8shu7crg1pThIHtgAhgeFFfZO6tYGKId8ViELwHFWFL11z
8ELVToiX/wVN5pJKY+H6vkFt5F4Uu/feUtArthkdCmWvC6XM9846KgcJJsCOtgMx/EsvEsfeYxhv
BAJMACxQaaOdhVmIl+NsqV1oQOWBc+FYbnLHLi7WkeH9HxDMCuASTCuuKLuI5Dp6Y4tkILNr8MvC
CJ62qFNcFqZBdwr3h90fjCr+LcZiIHb+9HQV02cZ79ACztMN0swStxYQzWUNJhWuIkEh88O2iKxI
SZz6/o3TH1BVj2dy4nKziyGPF+2XfnOLe8+vZDCHWN6xGzZK6au//uyFl9tXaX/BGXeFNk/v8cvB
Lm711gU7PtDXFq6/EpTDZ4o92opxJHBQfyUnt0LzaWS7W6qAwjn6HpX8GyLWs/MsOrn8BGnEWTJR
8+A5vKwoEubdZL30udVWI+LpDf8YDW+JiIILbMiUeo5NA0UXdYhnRZR5AAfCsX35J7uTyA/F9Kdt
wU0NqR/1TMMji/3258Hy+Svo7rXKUpmaDQmIqMJq3CEm/9Gdu7+MP2gxKx+58amZwccYXt15aeZT
frmN9fjzBbuYZXmFXFJEhzYJFgeaIDZOMmMv+WIKRJ0sjRdGYADdYOIZbaSm1acFlAK8P4IlNLEW
NQUysjzXnIBftDTYGFcbtYxCn3nDOpCeCGUyuPR7Bm2dNYngniSaDI1fXQBI4C8F2BKo/j9ikm83
BYa43FM9C0dN+vDD8caoxC37YPxiWT0ew3Wwz0t8wV+9Nz3hw77on6c0z2ooza24zpW8VC8uuSbj
VJeUEvoFxRONMPLXIA3t/7Bm0+taBMhKaaNmxZ/6pfaMloo80PAPQQu1/TftHxVzCiaKQhCfsG4F
nhduHod60sViioiQWzat1YrZeXBrn2cVqEsYFRvIEigotEe5suC4367TqToSrZxHtPHpHG4ezw+X
nOXNDVUZwYk9FLFSn4cgQnfHUrhTqn9oXITEl9HRcQ3wioSUSgHHcJ63Zd8HkN1tdBVqhnSsVNl1
0r6TymaKU0Ix7pJVZwYliqvifI2cXZojnJx9rgU4zRwtsZ0TCdzoUWKgp4mm2xVZLHAxe6fdxZ2j
X+4v/6wqrFOD5fCW3ciMrDuJwkzSmmrWs9ae24R/MHRL3s/ZkUFPWsZOCCFhbBKRHfyM/2DFBW5C
kELVtovsu8rfpQKC68N4A2e3Pt0ypq96ZHJSS63i911vTrdjYHz/yQxV7kmohj7dQEPjU9+T6FQZ
jfgAwxhWXrjP2ztaEoOHwZjD6rUJb5EJIfKAlrZYbmnUcShGgZ4i4QjaBmyrTPZ9ERT6vTNqSvNJ
s99DY5V1HcJmnqzC8Isaia+iPMWhGS0nUSb0fMd6FS+RafDfXbLqIyvZ2YGWs2gGcnfW9tA16hnM
YtAu2gAOWRAg+sjhj4tFD2D2B71CAEpbGQrgBEqGKQ96cWdDidblzUljzVUWU5g91trMPEVvjYBT
71iIv5HAfoFp6jh09yucZS5izzpta24u+aJwjYe21ZmzagT3XHmRYseGxmlAiOS6iC1AvZVu7Lc2
mlkuFAFJ54CXcNZWMQO3f47AzPYo9UVb+WVby1ygMk+QfGUS1efSYdJ0uthZwLbbIwel2BVixmXZ
QUthYuFDL3CRAC6DHBgki4Hw3cRxRhu/pnMCtcqVKYFdxNu8lwLUcFwPJEtDMnEuv6VigX06Mkrs
p5mkW9R9ZLpJtQgyjl4oMOYD4TErSHlZ3PQgUoE88FpqnezScZCgDpRFUhuaRFEgVMs6VrsPDDK8
qCc/kuTpbcmzrFuzEBpk7YN9JUIAITxYtsQhpquRdExjplhr88JGVWnnJU82mpIe7yMrOw7KvVvG
uiQn7ggpCnb2f1uyCVXSlRe5St7ly+z0Pz3ltCcvVp7YH2qmt3XO2p3d1yEyvPGffhdMNhfs+Hnh
u0MN6ruXJFb5EYeQcxLqw7JF6YpaS/C3typBT6UB6XyXCDrTmRGt8nM5HINV4tlS4Zz6ODTKgOBB
+LfEnBy5RW1xWyq+EgIIVrjRa5HIWxrkBh6pZhkmFdDScX7gk4THv9KfK9gjZrTiwH3fDLhQPPul
lPu4nE5iyZoAxgdmR951wyrcIouU3hYrUvgIBseMU6P2oRNNCTxcSvnrOu1eKJtKKDzxDh8eimCY
qIt4ijgJQiEIQVFE9HNcwC1HhVoUo8jcLSZStRhRLlTX2xSJqL/6zWHVt7p2NxDKiQuvf58V3gqs
U7ElARR4ocrtMalJ1M49uKMihl1T8PgXpbmtrviN8juM6ffQafiQaTrHTReknJtKmZszzXqRpY3l
D1Db39pKeNWoBcxoQQxNx504cgt83hRuuAm9dMFYUuZMeBUEdKzlHmK1K3aaagOnnyL4tDgw0g80
jnFtbqDt2dNd4einIeKAJubzWcUYdayAZfDHgHSFuLscjyjWca/b4mp1+DUNpYfAKWUJJuNzapLI
kNO3MvJu8lCydkS1Op809DeEjZcLWSm/uFAdndiUGZZS/rC0I9J1dRYMBbxn+fsdctbVa04E4t7A
BftsY06o3q+usrkimtoHMI/ZyBJKsrcVRUx3MGNedCtoaEOEr6xD/6iFUlBfRJifY5hn3NfpI1X1
/IkLZXnyoEG9Y9BHUakFn5+fRPbNlrc2KAqxocwTeThw7Gz0GEcGOOvYauu5UeiJI24QOWLrSUro
eWuX9rbMNWApEk4i6IFdAn9VL2+xQs6u177wi8Ii5oUpFsdHlyyBmmKmUeByW+g08CeWPIrbGa+F
mGhpcWID6HXuY/VlWi52sjzzw4tEM2CLbMUFdZhRmBao3PaSKV+CdxEPkes76q45PXSgWXVT7SJV
LlNOYCbW6E1BtzJi2+wuhqmj1YuaHzNd0l5tjc1bVBG44RaPNoYnkJsqV/6wH39Lw0SQYEvXOwXe
592ju+hsceV0HBUfKVE7cVQZX6wk7IvAWzcvfAugMMDt7LcbbZ57v5FnUvw8Z6/zoA1fHq9FSWlA
wlwoBr6bWncs3adGIbugPKhzuhaxQZU3Zv9crYs3CelqzW7uxP7bMpW8vZiJ8EAbhLtyYdOm7wRg
ueVmlxap1GMTFi9CUafLmKRu+23ba2meHFIVbnJwdECVaRuZrXc7lmibbVHAm+7vLVkujVZHVqJl
M4SqefPb5CZCzMMwgNcotDeW++uvpw5Pn6az1g9mFpCnGJKzD5OjPZqyAYlcGSLDGM/tTBTQ1Kwk
Ye61ds2iYBYdEeSxMR7qbOYyLPmIeP9zGU83wNDQCUtmIQCSxwZdZ+li3NMCx/y05C2sRu1MOyTt
k1IV5Dg8m1lU/S4QDcPQbb+O08qYboI0JCqHr3QsVzqNFPlKziTYJbhZW5Dq2TuieoLIz3J7haR9
t/0JB7C84fpEAgr7yJGaxrGQ5aZSx8MfPOdgYmF2TZuYvU+yUG4xYOAyPnRwZLmb5qHz3Si3Aro6
IeeI2qmQD9ntatR1gZTxqP1vKk/sUpRNtTFHzmesTusw8CsL0ouav4YpXNuv5lvXJYVP5I5Ek1Xz
MLZLkpGTpF9MKOykNTPP/b7lJLsF9tYk51qovz/grOkAhhOMdgdBJ36fCPxLXh4J9f0+Uh6lUn6N
KGpfpSURgopJh+ayxOoq/7LeVN2HzCUmV6FOBHVRiaAHRiTXcKNqaCJ5r4d0YPMLWy+piUf/n3Kh
lsr9aNqHPxW8cHcEbi0yygv+0hkAsnQLASC3PYpbTJcp3n8UoCUfPGiAGW33x+CfuAqm8pY9i0BK
wAmZCzpv6RiS3EvNsozhCCJ9aGLBfKW8HpKOHJvr0LbOfF+nsq4lUVZg+l23543vJy3ufvbpAjN7
LxIMgO9sjtr7h0NxMH5sjEuQwmWIYBokSfp4pzYl3rgZtlW/c2R8dwJJUzlnHYvKOAtzTLqFM1eu
MB8pjABCWbZfwd1RNWLQ3u/kvc+jHYsC/XWcH1rMyZzIV/VyB+nGqIxeVu0IehlciQiRHMK9Yruy
qMg9TNoIy2yTs+pjR3Ge2y2y87DLEF3Xlnv4+nNoW8AiruCURbRIclKb1jdVCvscxeGty96sQE3o
pPQRjdPxwBH0yjRu5YrVCDigbGtwTq4GizpPz0P345cns1BASJFkgYxy6ntIRXxUm9jiMqgRr3AS
62ZdIMut1NSuSViO+MitFEcqVpjYum8gWTwvLgGs5hAoxteBry8b8SNPKt5Daz9aRIzNO8jXRmLu
+5xcU7d/wDuvmYkTbeAMBmNlcl7Y6mfVU/FYwcszezXrswUx/S5RVQIYne4iWuwwgE5nAOZodz1W
g6mqB7K1+YoLWki4TGihxujnCoyUuEvgxu7QVbEL4Etzq4svUZDauFke1kC85Nx2ETOKVPbrqeGx
yzzt9yWX3nztJvX7BFhtxz4BTVcGIy/OTxrmGbgnW3yLVLRvy+zOVHnVhDlyHlLQ778uwA5qeipc
f97FdzCn13Q3TTa1p6hEmsyQPpmh61muKPKTSZoWspAbpBlnBrn37AMEjv6q8k0=
`pragma protect end_protected
