// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:27 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
VKLbunfcFE9aoheMtIINSuAE/ajVIAIeL7n01QKv1gr9T5pVkSkP5OozaUgXO37g
qpZ1xkEEP+65kJaeoesQeA04JW4FY3G56RXgrpAwbdKHWlHGb3x/yEnHN/tLwK4N
/57GVkuilrO4bXmOfI9VgUb5Efdn7Cirxmt5N2nPKyA=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 9312)
t/HiZsfh/DWK/KZLIoOtwu60vPi9ZDXR7fcAxPq+bv8F12ayCP2iRsoUAdq7oHRc
jEgkc3kxOPnXvGRCRsaXZ9evsnpOoKDPGEEqUVBXaMBJ+B1p2ImBrPpayoGUlWyf
Fez1kpQ/ZARVnrWvXdkiv6oUaUncmlUOdLytBM01KxoU98ICmxpranpUcA3UGduX
jMT/166jpWTZSjUpcYUHT7MEcTYEGE5r2NbfG+b3GLw3d7th2fKf7XGGp1J7sXJB
6uRwA3rHBMmPFa6i0zQM3+vHydZU2Mb/UC9tLoOBK4LijvJ12ha2w4rdI37R/DdN
6ufUjd5bAGOlZx/xS+t5CSKrNtkatEthUUbSH5Vrj42N3PxDCr0Px0LgfyBESrNw
+A6mkR1l5Vu8s5HPtBxNyABqLf8tEhxj0jIYP257MsolpVAzgJt3SvbiaaS5YVQm
epgOy/0v//pyTbppLcsGBYe8hMoapZXO8u3qFSkawmMZ72LWQEk6WJo0w6lpCg+G
K8/Lgers8j4tdjfafn0W+hAJuv9z5Mpo7dNLYzlyNPlCrVlZ1AOPtVG09oAyn3x8
VnnatSvCv/x995AIJsEfpkBEnKvcyMamak6b/Jw16At3OX0yLLutJNettaGbWrXJ
AMaU2o6KVVR+VxLMh7k2sn5uY2i242g55aWTnTEbWL5eAdVX8pPxbdy5k6gngbTA
l+19JdRLUtyWUpVppwzXMc6T5bhm0PzlbW9UBt4Z6s+IotQtPNv18Zd5b4FrAHca
M9dAFK8zTiPsXuiqt2AHjtB0m3A5h3DHVyfyfYd5MieQ+RdUdYJKILF5pfwFKkiS
EWQW+hR+6rwP0oofbzG5z5AL5fM2clPkvaI26INydQGe3yruldyBh6LzNi/6/Wep
Ge94TumXoEYSVh66rqeZFamhX7AQmepTaMeCbOdFy+RGWAhTayLHgc6Zh0XH2A8K
+dJ2gGGo0cDzhK7/iJtI0tlzO0ObXpi35z0u/TFnv+Ax6Wqi6p7iQ6NyzjsKvN9Q
qwMdgq4e2rKtWHmKouLESjF0NIrKz0laLO+Hpf7lOfHty+Exz7HUhmWxPzbC39YB
C8zhC+gV05eTAAnqU78ym4Higy/NHErF2cBdj1hja7qaMuP/wvTBuWeOrSjX/oYY
Bj7Oe4tU1Jy00tBxHbthMPYnnEjrWkm6wOpTUZxjsYCAe3+kRTc33NaYwpVNlaBp
gqgURkWokG8bgVowqNFc+3NaHCtH3/Wn70PoJIHXSZD+1hHWQSb3+6DIPYCOZrBV
oNXO88VBMAgrtlm1e2/I8Wnj/folUHrj3/QPFw0AE0EtIY6SMwI0EoCEbc0F96V1
YvNyeMF0ni61B89DMlQUZ/+Ch3LATYOg1jK8gVc9FZ6XhLVZNewWPJ52dTtVvN+Q
i15vM6J182GhvyybrysohSV6R+dTBuPgkYQ0gUKOyS1AvjXXUF8GYyHHfxsjsm01
8gFQxegthkP20tj5Sux32SslJFpECSYfbcCkFh9nrEWkeGSmbf9GN2NoaGo4T8Au
g8WgYIl9zPuY6ZM5we3uI2mrvhmZlvgg46X2mYQ7cXu9y7q/uBJG//JeEJKjEv9c
MvpR06rd2Yqm/r6FZ1Rc4cZx78Wfy0ooziJNNO37TcihkilkiZmexrvHi5iOfB/1
ndEp04ap3Upds5Ex4kDlofvZ7uJguWn8RsfiLe0ZVNPyd7m5UUSdcaagujXshe5D
Qb2rfvaWlOpXgj3tmF6BDpyC0fJPRfP81Ete3QV1FMefjj+Zh2vehPc76Bkr6t0m
rZ7MBgmm1htRNk16Kz1cja8d5DMQGS/4znhbnQAlJ+mBBDXbzr7eEnLqHOPY8tPq
lRhWkJPWu7EPEHfzKzvzgbgO6X8XK4EIkEeT68ceesp9jy/V4eNJ2QR4psMtFnSg
Np8eI1PqKU98x2PqJ1rtJ0dOoObTAJUajBz7Lk2/DT0xy7jlFm1zx64gkVtzISbC
rwaY8Qebf6tzgiaPsI4Kedasx9uPA+z/FTZSdZn4jfsz3cU9bvA//KXWyx692GQ+
8e24NdivYagjlPqZ0c1kVkR0+fZdgD63WnBnYKldiZLqMG4OvHoWmDvNqyKzcP3U
PR1Lp3lo3uzcxR832eyIjblImcGK12qm85upehB7YIZMH3ErAkpt9LIKsZagsCXb
6LwOqaNUp0pTFDzKxsJqflCYJ3sbOf6kC0hVC0i6/VbKy2Iif8uLG8iHwe5xraRd
Hn1duSDjSDzzWsieLSJtCtNsa0+F7kfnP03IxIyZ3TMeNYq1onk2GGubLG0JUClN
PkfozNxxJNxgWLvGzT4WAbMrszOG7qQJQzthGV8PH8cMR9HGpVOgFpacNcpSIPZf
9ZW28Eo3dM3goKNfGsYg7Aj1yNZR9jJ6hQhGfoSsv7J7HjNrenTZEVZePnahp2b5
anG23fJjuXbh2SoHeBGXna0e2covCUYbrl6hBr9J/wxmbE2mwMdZZjkgw72uxJhf
cu7z46M7zEd43c45xHrLvZ6rUW70Q/tQrIKW2W66axJ/xHPnKIFCHJd13NKuRBkE
9SLCmn+Czd6Uq1JmT8EPOyzYj5aSA2de+E2ilPogmX+29plBr+GU/6XMHJ7W7aEI
3V8GoVQ1FWN8iJLmOBgsJHxAaANDaZEz8ed+96YIUWeF6Gtqpj9VWKrfAAmqKkBj
IkXhnF8fXOpW7AIvnpk9x39vP8TuQxgf956O9lfzOVF9ZrxpOPRtTWY38qbp/c8J
e9r75TxfXAjlW1u2/TVmHKMjLS2pTjLXDnOgCcwoohHsMNWbd4OZzzdmhFp6S+u6
7prdB3VzCAvX5Z4tlq1EWyHiHvGLEb2qqHAE2BmKWoLuSadREZ/ng51pHg5ZUcP3
D1E6SviRaVoPKbFPlqRupmRLRRVwXWdnqBTu1ivuvI5CjeT+mAIyRmNe6b5xTa2n
2nTpJiivUbMOCTL1ZaV+bwKm171WON8bhk9d7Xvigr09FosJmk4kAFr3p3Jk9yFR
Zc/33cgJ6RKDRRk5WG0ZQjiR3nbj7HCM720aEV0QGqn2x/fTlcOZSuhYmn9JfmJ6
eb+QJv4pOa0gphYa1YkolMhIYjAKSCjSKoAGveFwb/D87P+c0XNxFQdH4JcUwNfe
ETDiFfYAOuabAAsS1/pT85PYeXgc1qjw5aJrgJyRBFtBgqbqmpUI5HAv4iPdjGWY
M6Ed5qT4SSZk/9YL1q80KiGMyPzCY6ovB5MQ+JG3RGyHPLW+1U4nE9a+FOxLj9bg
kz5qre2JP0iSeDjB+fUdWauS2FBZCn2XZhYDXbZFH54OJq+z6nII0Pk3es8lgPKn
prJ4a/n6L6TGfDLQiksMNEgy9H8ifizMWABx+hSUKLlEvdz9risqhCzEGG19bJ1z
t78Fs6AGyG8l14dkTIgqafeZHjH8Oa6WQ3ahm1HJbIwfHmCYDkv2rJlTwGZsYbC6
NFuD35qXkcApmROZWHhkHhmL9oNF6PphQj/hxeS2g1ZG8oW2rBwm6Bi9Bjhsyquc
RQ9qA+VuUk0GpWaPLfg5VFYGc1/DMunkXb7cthkdlZnep96hxRoTft/CKsR/91Uy
RBd8C2LNthM/c5i8eKeKkvhg1IBftuNrwUntCcBY+qbRltvJioZu0LSyzI0qm/+S
lWRa60/JCp+EDCQ843IIxr/46kS78ZqR1rivggq7AAegF7+ye6UaZvqRI+4zqwbq
rFmB3wJew2fOPtkSg4ZolKtCaHAecJpjLePexFE+0/MUnxO6AdU9zYQ7bCpZ2RlE
RAnUTZInNCyG8+3r69B7kG5O3JTExi4O5xkaPHPm9h/WpAfdrq0zOd5xR621cNKH
4JaqfBPX4D1f+jbUJJDcJKLRa/NLKpTzk7QU6kP8u2zaSLaZWPBn5XvWOMAM0E9H
263hi4Zok8FPiu3rZUb5rr8IFgtY1vyctnSivvEQ3QHQpT6ipG/pO7ZD/cqm6Tll
E7XiyAnj7sdOVPqok6iYa2vDrMoNQ0Y8Qw6pxC9/YqqeZDE8JDEGWTpffJlcZcwQ
6KLpw2Z7Tj9YIiS9iJz7iXPlHQUdrHjrKpDYo9viBwLEJtIEUt9THC2TSHiaUlC9
OkFoXQ1UQmg/FIqPLfRmICMi7JStu4YVvNcoLfjxWxWCXR/GgdzfrQ2HRCCI715D
U4xCUdjcaudznR9F1Fqh1jzzrFcI3uNO/sMM193lXoMwFT+WUhaoYw1h7TN1KT/r
dZITW1+1qUueVivRY75g4Ap690kPamlKu/4Das9rTIhGVX5Jsc+h1WXa5POTEma0
ePRQWGicxq6Swhxo1BWZcbzGOBA5UcGqNEe6CpYUO9RkYH+tY5zN8ruDKV6gUJTh
Dq5ByMILdsiZEq1Ng6/yXzZDTtN+QS6bpTViKZZzjJRfBCTclDHKRVNaYONB/j43
RSGEmnTd3N+IvQKWKtD18RW5h/BEAJN75XSrB+EUUjVOA9CmOrafIRn5CeA0D18f
3Znf8v6oAvl+bR5ODXMy+EfuZ9jug1tObZYl0cKXQBeZ1lwM2dHVK8azNs5YMoWr
MRyWpSUncEtYNfK8GknnqJLAvi1sHSnpdcaRS0Z6G3cc5hvppUsvdagAroRGpGUP
yJfAwdVpkVL7BLG5L9Dhq1UN/4i+Yk9SwEl9qO0FJqKRR/xwdBBK6gb1Jx+66avU
UTsrQbvGV38SHNNYCGIxRlT+rbS6vsBsiMvGIESq+I8vbwah3R/1HIpSBC0N+mDl
A1L/SGORjh3FAZBFENZQbrxMttcmQRM7Jnn9laVcWYPFVKmEO5nhswyRIwJcWyy7
dy467fa9nhVdOcbvimOOL4Oy67qwgh65Giwk8cKw9zdp/0kbsGFyGjNxKxiQ0QfY
jceEYASVg1yeeqjceV0awPaGs++xJTyJmhE1iLDxuAGHbj6GVfezLvM5gB1DglY4
dxm27O5PfXrvf9cnUmXd2iLKRwBa7U8kT26yp+ZwNfdXSgQ9R1sXLqerTlEyeZE+
CrljGX2iGRY4G9ME7RGVhJD+vxLw7JTnQ3PPJyeY7gPuOkg3Txus0Bcv9WAa5vtB
3vpqPlYwq0HOkYlyFXJ+9dZdQgg5OCw8L8rZTwlDxUiCcx5v2t0PFh+vIZ3YcgWM
x3mY7DdTVpn86lIQTvhS6x7Ui5s3lPmFjksB/NooYpraRxu0zn9AVZO7t2taztJY
u4MAUN+Lfy6mQ0TdP3fMKmgihoF1B2pUsAz8fYCtZTrGwm17gvK1NOD3ae2qhVgr
ORLWFwYPlJcua/quVRZxuQJDwZoH7iMvVIclhqQ8nhXWJ+SIuNXEWldcPFsK094n
qpnppf3u+C24jnIGMF6+eBJGWjTc9g30jYclvFXfDgD3Z5Ig7X1VP1zHCnWFqUun
cyp0VzkLEu3cEOYQSFZ5RJd42fYfLd9ow6yvKSqi1G2fCG4P/EZgyOb0CwMxzn0u
pUXODkPGpSHY/5Jifs5zbwFNngyN9asQcoDycvXcwMdixbKBgW7Ay4mLgQvtd2pn
EgiPtaM0Yi2CTlkCr/fb2W2hsa6pPW/qxGk/8W5dCKqYhRsHd7q5HIbEmuM8+pnR
e7Prjb8hnM4WaDvmzObvI1goMGu2kRIdd8w7GK9oJLBnuggTEyw6R8mUC/+fdED5
waAxA7M8gn6gFhyTN7I7noQS2TqShS6sByBteFtnh0JZcHSSs5dLp6yQouF/F0vZ
OvmhhB+2znWpFK6NnZr8l3NRgDg5+eCnNa4+SwYzgQh50gLmXekbUUzV+jyYQ7U6
q1BWRbvX+WYZu9IOpR+HVJfVDqtPTlrpSpr1JBXZVyadXNO4Ax9gnYHgqOcwYWx3
1rCY8vf4+UrtQsyLY7V3s86nI6TLNgF6LYoruRuvROlxP4Y2rk0f3nxjpJquvHE7
nZQ7jTFz7p7uhJu0nTinSYXHgB3xT+DTxwqqOONSiGySrw7TGTvGtE7DNLwYvhDh
wkHOK1Wvbg3sckZm6BrMjh9H+kuo4ibr+HqBW/bky8B1qYQf5Zt8TTFsFDRvNKgO
YtxOEi0Yy8hiUYPjUZckTBgia05OCHmqBAAv5ueJa17KHTDfQmWbCXfZV3OuCsNu
1KkvK9cQlIzHKUD9eXpNTvjq+WkRS1kYgAZQ6zGswKMaiWrlHgZUI8GYGBxxkITQ
Z7kzgyydjhNieixo8Imce5J7Eg6utET7nIL5OMysAlDBT6e2KduXcpRMAgFf0BRx
Xbrji45L4GTmbXU3osh4Wx5+tZ6vcWfZSWl0w42Pb/ZE+0sEv3PQn2EJvXA62Rfd
2yavpO8bl7QjslCrDwBoin5hXkom5BRzBTfbYTpbkv0fBcKuW9YzyIlRpkpb6i0Z
JjSEdyFQ/+jYNZbrCitWkqvIQj24rb2radSfS430s4ARoAQzZPfdQSWd/aV4W5Wa
4WHgLSZjtd1EBoTD/1RPxTcz6RnM9NdAtRQfringKcHNHZMPGy/UiH1/hWcC8ybs
9JgogxxOcdbiQsrlJQ5dCKiZkhqFazyaU2fRdyaUijQvoKfV4aUtZw4XstuI+enJ
EKbRrAYCRsrmpemVXXIpuHF3y39MyObAcEvBfHTuFsP7N3WQl3JHQNCWDiTX/lQF
UJTVOemxwp6jyHEqpn9bA8JHgJ1kGzAjIdpXD8tNsGqRHJDjc99qKF0KPlYaVFgI
h/UJEWoNoJTADlWo0IFGOCaBTjFxFTVQv/0u0h/jsniOHOS3zxSP8LhU0xPQTe+r
2niSnheQGLaxd805MmvwkhH/m4ro8B/oxl+NIkcXyC9Sj8ieiqlQOORgw4+k7/3C
709Wi45rV+qSx5zdIp1SnsZHoiRlKQI4XG2pM1uNJlonHe8AHJzHlw/CBdEZziyf
0e3RAux9oFJTEIv3OoDGZ4rFkFdBa89wc8K4KjYAmLtpf+qw/hNcP3Phr3yY/lLB
dcOahrarGFbp5zFpIY4px9ezLNCPqXPnNkSK/m6qrUrFUVgtR/m6L1e0vvIwcGxm
XULgbaTaQAjD91I/97znxVyaPU0UsqEbyWzXA5jOd27YUTmp5jMhsqldBIBL+joQ
QNYYzZJL9fPEfyLyP/B9H8e/IlKZGWlXHIc36tD2kcYW99xfnnapcb2gEGStdsM8
SUNNpwS4SPCNz1FCyBZbIcnxO5o2L77YdMJRpaqsadYs3WyqJyXCNLxRzDGYWWp3
x73AYuDl5m+dy4MGFwYhYRYQouN7AI55MuIvUwpNE/E6iRlE1ERbNYy9hwVglr1n
vblaMn6IEBS9iOpC5m7QOhONN8hsp0U2CxzmtcyKipkyXQd0fJHurlFhXaB4Lo7P
sFGFDy/lCBMlWNvKIiIyrvfGzeb3KP3g6qDYzUmQ/aYzZCfK+zp6S8tIwDY+GyXs
FjmrCXNil/0NoO4xHZy9hoXt3t2bfrlPYNnb/dV/rtIDeoKV3o9Mkf3DCzgrGNLi
GkoBitDzLYp3c1URffElVrsh1VG2z3pJ6FNUdXOGXve89Zp+OnFlJnSzp4fyCION
3FQhffupIjJU1sd0/zvu2S2lZsdYw9ZXw1CanMvmmXD1OQ66FENowIPXUEfSFLkd
RHXI+b8+QxIuKVDpupjMC1d1dz3wtg6lv0+SyKaEw2XiYkPEZzvSccQUEOX1PBCB
pMw7dCtH3nNCiGqyZolfcgvn4twtRUSB7dlT82OQURLDmUkhSS8nYEVqiTAPszPi
ZWTgWun7lL9m12bfkftA2p1KG+3THFcL2GTf/XdCHu3x3w1K3c6l81xHJ7MZInGQ
1Vwok8RoP1oEMXBw3vTnexXRW+XHmZ7gds15rUrnKbRjiqXSSu1zt1hFIkyuik7w
f/739JfQQ/xaxIbEZk7qobJvMbN6xglwJIiiDu5yghGYYJgwlMIS9i9RVw8ke0jI
0cMV9gN1xh5GbDvLqePgpYv3eA3zgYQCRO7MxVNM/SqOfQgTjNapuyINvlpauqAq
5bx628EAkPfWAcZzDUfqqowa/TfS/HC/3cKUatE4GKwnhRruXBqo/5f9nBGYrJa0
A+s9w7aZKueN4+y2jlUD56WJWLR+P6mcJOX758nz0kA7/pg7RryXgtM4WCy5t0sY
ZHf4ILB7VA2nt9BjX9Ihj2/OImRy6Jh473OXhv8sO2ibW3jAW1mnlQ5evZ0CBIlf
d3xS3w7VwpK7VoSMKyFmBLtS/yRxj05xShTHkAV2EWUxf9xqN1g346j0JNsd2YGE
CwZwUb7rWFiShH8pVkNcvfRDz1DAs8RS3wEIbXrGgwC9LciIfgnAQ3mtMUWthxDh
5O7wA7fbsmLos/d9YzWH8AzyzfVmW4iWhufFUxaMT3Swrper2QMSopEuxV9OKu3+
03IV/V3xU9ZTU0hxg2X90rkgLkbXlY3/k+XqppM15fc+vXwPYGkJx7MpQrIb5Oeo
ZjX07bD0yy698QnJqEjqSVC38Zb7d0XUMrpWhwcG6XAyJMCVjy4uePfyGLsLvsv+
WKvVAJ8ElSt55K/0ck9Nnp8oEH+GBLY0OZ4ELgpNkT43+CLCK28gHWw7rXMg9cbD
UP5B+L5+pNXjIyYmK0AgdRTTGdV+ZvKGGqQV16tfe2bvQpq9ihyjA/ekSeizqgOy
B3hMc3l88hek5CtNr4KfE3FLHq0NtEvoYZ0ythA5LQ1smTt3qOUIX1wXmZvfqqT0
/1M8H76eGF39KYkADRj3vECt5IjyekvqoXDZJiKYhRCEl8NhHqJ42f8edhn0jeoS
DYIVr8Ng/wOe+25p9DMvp8iqgSziKDRO8aJkyBrgOKxE3WPT5ok3kqLKIsXYFodU
6v1XaNqpZ7ar0oZOXH4pug9EuHtg+F5m48FCcpC24bHPEbagrniR+r/cdNWx1ZuN
6+WQbvXeBqIGbQacpKqwP/IJJuJgGYfKD0g2E1OK2AKTcH7u4u7q1NR0lmmSpNr+
z1PhO3JoYAE+jWbLXnspXpIbqXGQUU9S61UJZ7Yw46QfJ9pN+RSL5QqZS/YtexBR
rK5bPWvM7jWfupWc2wjtlxfmbz7qKHVkW96gKOmoRUikKupM8Sxi7XYvgtgAoMQ6
yad3lU+SMu0pSw6JwX25ot6/QEb3Zbiw5+HnRMZ3WrLuMYh8zwbtBwn2waYN4Atr
tSK/wPjlxdqDJJlNvMFmIl3cKftmLlQknrJmAlqn9NJ2vowiJ7oxLO4NJ+b/ADgT
GtoNepRZuKeAg784Y5+8l3x4/RtP7DcPm4dkjtGOLoqRUWybyG2HXUBFIrFuV8QG
k93IK0KdlEGxgVVxCd1hfl8+d9Ve4d494izormtWflkwsWapOZHYFLCrAZkLZdqV
l4sw9ZcQg2AnLacUh9AW2umsNbUnSgu9vtWEzzI8W6yQPGXc3z6d6e4hMXGJcKVM
qBIcbV9l/hCOGOND1Qgk1mWC4yNtQbL6bmfqI6eqJ2S5NEr3CmocZ3aC5tM2avm0
BxA69fqr762KX6Agens3VG78kDE+4NeCWQF9LhMZXzYqePvrWzG5B0P2bEVJbpYr
d1JKk+t5QE2R+QIfS7K18Gdo0OdGCUUzUqvOtb+lHtSEqSEPo4PbxsOp9cRilq96
MlYvoUE8D6xf7hoeKQElMwy5dVGZhwMxi6fF6wcKITtSZaw2eMJkM8I+yDUg5DVY
6xqgCk79ZLtFkEOTftyWlKveoy4Vw4OeDR6rZGwlP06vzv7UXBoZ/k7nhwnn8Avl
izRlc8/33DqaT46L/7tuamkTgPiG9o5YztxiVkpq2mcO6u9+lOfsl8fOdby8aYz2
mGAtkuJWoHOvP+Lmh8CAEqf8UHpbXClVf+Kr9l2wwlffWWjfB4OjfT/tv0jYvOii
2NsWmSh4YqZbOpP1lfjbTC6raQk4l7WUv53ygOdVoKtU0I8+lMsTFfmRklEYTGJ6
1DMLU9C1frIjUFOZLK1fkrfnAeBwJYdGa+krWQn8ZSwVIWCGNTKdJ2V7nzqy2Idq
v2Y+dpDH9W4DN+MCcgFTNSepFQrrxcPoeMfYTZlbu5CrvSwn7LAEXeeIeTx4jeDF
d+naUJpcAKDWb1CE2LC5sl4p77HCJLYb79dhNDyda0tVZdXkHnYZQph5PX1ZcD92
naYEUpLr4NW4DvvzDJvlmfYHuNq1HHVlivziWbg1CFadLxy8Co3sHGomivvTF2qN
UGzNVHQtd0o5tvB2DdFJ6+Yb3S6K2m3LfRLzJyge7uZ0lfL5Ipdl6J9EdEhSlmS4
NEsnUeKg35I9BR1AVP99ox9gLXj37M2ZTwR5G85M7HsN2KzIhfEohDZ7HSSJJMeM
Ob0aRKmvnEV97cY5mhk0ho2LVQervXsThZ2FqX8sJaAqi9AWwdk70O0w2JwWX7it
bsGtHFh1gkso4oQOoKqpU84wggyLIjmkToJmwTjw3l0/V/4flDhCjfMoS+/gaGBU
5UC5mqRZAkgl1rhNfUTWnMbeQk36taOgaHi5ef6hDlctZFFSAFReChfZETjF0aqm
pJhvFUhagGuaOUdU7By//+MFCgpz+SpplyPjowDBxaPFVo1uvzv216eI19eYTAcV
V25W/Klg8p9GJ91Z4NdKcEbTrFxImEO3kwFHgNCL89js/70cAk3vU9EcHI4NQPqE
KfaP39MfkkztibQHRk8rfXaMefXsj+oUyRjxZHXAOGpT0yRye4zPw9EgigZtjxlK
2bIczmNmBLzqaUAtCsQaGQ3Hf5HPmz1qfLYcgjhCqA29XsWX9eOyy6I8II+Ud6bD
B2vhDzqPFrEHp6YUSNOQj8DQ5EEIZdrQyFRvqanUqLAvbLQbdrRfHgows8YQTbd2
5u18jf/fCMmzUxxu2AxaOb3fmWt2bI2B6FjAovszBwqzWF6OY6fJEfZX6RLNXsJo
53p94nLpiFdw31/ld1MsHBxsNvD841oiolEEgximZIbYlrK5/jx1i3nvJjVFSBt0
4U3TCCEGXDg2mD+m6xNxd75Sa/bofoklm1VNifRg8p92+GkSQ005R80YEK0jWB90
37eVKw12j2JFEbi8WX9cbeUF4NyhB1TERc7fgCEdenG/tE7v9WlPLM13kQ776AMx
igTLYAlkhCSm75rbwENsc1Bd477IkxSSPVj9nQzn7eKv2+6sH6FAsILYEtR8sNf5
pSHKcr1slPsig40lZw7gBKykgAOWi/oo97qdqxt1Xa8n7wTD4zy0OU385EZiFo6b
pSwIdXiOvcpgqoMuxiiKI3AL3i9QKrjK9gRRZJ4PGF2KNk8BsnhbzIOL2PO2mIVC
mEIK3H/3ZKyr1NwA0HeHtNkyqVBrAXz+KQap6Eir3iy8uFk65PQqrL2TVNuOZzta
dxSrQb24LELgteNdCekMSuB2LGXLQpk2hg8Bj4g8NhQ4CZQqDfWtPFi+2soDiobi
67K7lc/hJQFbuwNuGOdyNQAOn9LRQdGIZCnogwwlA2ltkRpESZE5PVvoSVF9xpEj
UYaqw2oxx09rdUoG9iLO+1877zAbn1e11mqxsmOggfMJo+QLmQ2t6DfKzuIDzKUW
9fRk2ycw4v3SOIl2fTX0iDRwJxE4UcejvKEvPEFfpeVL1Bglu7i3tbDoi1I8jn1L
jmfI77x4kq2NKVYDFnVXh2xyxmdSAYj7vljPpbyLVXQep2oxwQ3CB+5ymvAb50Le
4X0bwy4Fcv1vNVijPyL6o7oT8R70A5dJ0mBGoB84nlBhZ5zHsPaK8z7vz3oHG9Ja
arqRZ+0MPWaBj2elQBS36gt8oGA8a0VZY9D5Uta2uCXAYfasukc/IZNQEcW2Irgq
U/96CU87L8GH5RvsfLZSa1RuXrWLnckFo5WieQNRPU7i7tuS0Mb7RHuPWiuWBeRh
vjJPA+jgK+gNDUmbjia7dzTkC08jjLR/oN25GzZdx5N48epkteIRH8bRFoPS7/8h
aEfZAX+ZyTery3d/L1jvdqBKCotMxDlsCDjRps5dnz9XC9NwJZpYCnPLyKnqd0is
pYNsE0/t48tJlfPQa4RV/4ZTlvgK7ZHXofrtUYhY4j8TqvPeVc5bNLYNDRmdztwD
//CpCxJ3dHyn0CevA1PEQRiQBEd3Dqujs6rDa1ESNPj2eBOi0lgo+4CI2s43XwUS
5c/5EdPbSWwkSuNgwd3qesHaJTJGEbki4H4pk0Tzc1p2qce3QOf6Bip/KckA4pOK
8JqGgHjemMZsFsGrp9tvU+/ThgiCg7mZET9Lb9LKN5sq8t4yBXXSDABycMCSveYq
0KgiRt29wpo8rE2soY34fFzweL/EyIRf7mrg673ghSHwKxU53qHeDNmw/6PJKL7V
JlJGv8i3jKW5JeCPqLcKgZlbzMh1EPU8UD45U5wm34rGvohEY/mkWBAxJ2vOVz20
+YINoy99T7Wh00c4zvF3Rm1eiDpCZwHWsXZ4eMv7Ln/4fhQKVWANs3u+k8NeMXae
27oS/FW08F1ROSF8N/Qyu6yodTnslNilDbQBRxQK/lM7lHs+PzLYCLZzWz6ZFzZy
`pragma protect end_protected
