// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:45 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
A00ovTfBVaiMGQVQnbc/mQ1AhZwWIUt9CscyAi4OxE9LFbHanJCTRjKewVU2mwZP
Ixbyr36MKvVawJr6KYQa38V9hmvTe+UzURUHrj6DOzW/Hsr14GxEYWoZZ88/9V2d
CenTYvKgCvMKy+iNGhRDdsJ7XXbsnuizZHukIamc/WU=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 105440)
ppfbjgPq4oKe9C6/SbQ5bxarwWiCPDNUmsWnm+pp25s3QD9WadNQ4LyyGHgm6d22
yhCcOoNOeca3y0+j5S56U+N2jwO7xqXC0g0aoaxebD0ybONPZbFaNzvqj21xm3MY
rmPbZW/UMrbCtko2UilHN05juatIiHe26FdxqYCqlHj3H8zRq2qe2dJqRipq6c6i
wWgRO3kvZeFff6hXiJM5eX2+9vCaAvLDN5o2hpDAIKWSDHvJE7YGtaB9toGg8IxF
ZUgS4bt0XSyeb5iyJNXRSGa0Sk3I7EyfBfx6ccsPWphHYQezr/9c//x/IQ+RzGge
IOj4n0aiJxvhSuSsuXistFHBATe1NfidwNPRBAV787IZQKmcAFtsjpMT/NldOBhD
U+Y0t6ae9M+5fQ4laSUT1q4UIP7mi/OgSaK8cyXol9nTZKStUd479cwMyDmdIbjq
b30NrJBB9Xv1Uwoilc1m3vjV7oZuxHV+mqzoplHUpMdApN8S/vZhgTBEAfX1cxFu
lBllBddtLBZJALsrMIxmfu/LbrgPHfglD8SYUtGP0+xqty+quK+VnmcaW4qb0xVe
Mm8vrbzLrZHPE28mFq0U6iQxKnJAMbIYRFQ5+BTHh9Riobh2vLL3Ddmfs68DPLr8
MSMu19/u1dbxF4Ytpde263mMPjVQe6K0rmXXhTV1WSuRxMzXwih4r5jxDgdi7w8X
PY76rupVIHvxGwDqo9d8KnphEzTefwF+UbXFci+KaJMt6C63l2YisgzbD42HBrLa
hcuCrUEaaOc9CK/RwVX9p2FgqUhO1BA1kq4DK75C6Y96n+juU+Ql6trYJSsfzFLt
ndDqdhVSsWGzPvuJOHO+6Gu+dSOEh9mYc2G6nqehGWIAa0UJOhN9eVNoS41vCIVq
uCfu8xsyDRi1wU1RqlVvxdxIFodQ+ewoL+bkKrrwmycUp76qqluqku/eiCcETvBl
sdj3vaz22ulgGxfL+NSIADYTdpX7RrttlxELAghhdOb1GO0Jd2eBS6hiFRGaYYNX
RNE8r6Mc/Di7GiC0/fvX4ZxLjJ13ArZtxWAGxhpP3ATXMozwuXb45xvfx/vY6re+
1bd1GYw8rMXVCG5JgLQKxAozGRoL5gigzGo1W3UKwZDC9u9O09nGzoQzARLviCfC
Im+6vPQHDKTIwDiRI6D/uwFwBZ2YWeEYeFmimVvpoK4FXnvu4gdGEQZRdlkniKn5
qw1kitWPV10l2xIJO7dZ/dwYDf36iiRUkj9JeklhxZCbc0FNYqB759l+Cy9PaZXi
c6h6gPXaIrTYfq/3qOTsrxl2p2A+Jx/V/vaxfVxph3JhUyRRg22ZbpQlxgZGo2tV
ObQHyUWaZrLZ83ZPV72YiHvoZ75yseDNapq7S6nquH4xzCRQFqF1OZ7+Qff7pI+1
+puwcOQrcsuywR1U49VULzcif/8Zw48sklntVjqA6kuSG79+zZWQmTTGOP+x7MO3
BlVfHFQhovNRZH+VAPhN0Yx8hn+aMcQnce0DiaZOjLqYW8Hi+4Lb4nGpYeq2keoO
iw9f5SutOiRPNs1EscB1qvvzt4sKoPAv7BlqwKt4GCsLzt/TjMFs/CJ+vFV4whm2
pDXplrzOkDk0KC9CzCY4jySkyDu1R+ZH511ko/VD8xVS+ylIuhcvAieIwcxKwnfk
+oKemzWS1gVUsX95kK+3BE0HdoHWQ7t5oCxFuEjbcPUAMft9/Ju6u0mF7VfLM5GW
qTxHo7GYgugIzuYpPD40HlBQ2khz0kSLu1VUazOcSD6sAAGkCVyPB1AXQ8oze94o
65+j27Wv3AR3MtTgJElGca05Gvuzokk23QpsGbFpMA9w1PiwsfR8WbUfbiwmYhRC
RNawMxGhHOqCIYEH1AUpAhYnfNYVjUkkUHTjEGw8vwcVTfK9H51W+Hc7E4L0ABHG
/yxfzz13tbtuuHWdwPsfG2oTl3rFhLV0APrhWkdPJCQXNb8liOfTuzvvEPj6KDZy
rVtMvu912g5DTkdTWuHS1Vp3hckUJorBPcKJsaP1DAx4WlNGvfp/Y3QM5X4Jfnqc
msfGQl38C4ttX9aWLdmanJiDhB5F5zuxxALA3zWQ5coPUE2CsndOHWE6nyL0/LFa
rxrySBW4weg9XaQT67iWI+T3FT+J8t50omvq7rGoidmP8WtAVUdjbcBjo1C5BRWd
exGFeDOT38sbIh0YhLUDkoVFlfS+GNDWZBYsgUcc8CJhc4Wo1JTZoeuElxaoB9kF
sHmqNE+EtFkV4GZfRvqUXfDFdWa4IBK4OK6UpZiDEQas8fAlrRe/LEvid456nqUP
3eoPCmzG2EEGhi59gO3I9jp7DCLwLWdut/MYWXZZBcTqQuZYOtyNpz/eR0ax8cK4
6qnZv+pBNi6SQQVVjjR5ctBfZBOxoIWd7hB6Ur8t4c1Dv6R2Wfr7t2nwYxU4YVQe
UDqiwjWAKXklCtTMGMTG9ICyjvpu0xLyhoMBem3Dsq65YnNVYjsGi0j0SclXluUf
vMGIiKUeffARQiw83UNitdboFd6lLiHeSPM4PuA5KcKEdoEjQ6poW4uv/3BbHdHw
/DsrZl3If1tg9Rp7/gWW4ATxEmzXWjvl+OkXdoXRjcBiI+FZScoa+IYzU+LQF70Z
MfTET4ddFiJ4/S15yPsevjrnZmYoFy1KVvIHPv3IuWL8tfbZYqirch2i9RaGknln
qdSGDIoKWx8OYFAKsXHZUvrib4LGJKoU6EaE8nO8rlJmISo93EqD5SLXe6offgND
RG/PQ+NT/4ryLWYZZb+HM+yv276+JNAWgJg7UrWMePg59QSoWh11idu1cFTmChwc
OxBKGX67gVj4jgkzIimxLNrZMyXIhw5/Io9BAqvXwvlCkUAJW03iKjdXwyB4nH+h
+14Nsn9U4tmW6Y/dkubCWGpZ2428ENEnJB/TGILhoEoWnfMFy+IPcZlQRrkMjZKt
IrN8WcsouJt2nS1Jk3ISn3VqHEmQCmojDxmXP6fdPODD6bT2O801H9AusxTEZeQ3
FKazPNouMsEe8ZG3aXJTo/d+hsb4+dtv2FqJdVMHh6XR4ZCjqel/pr+3YRBvjjwq
O/fK1AJqI/FlALQ8EKkIyizN6fRz0O23w4gVNA2QuhwYJyEGEKwvMBLcirJdayRI
Cmgey4QFTIs4yhYu4S0E5Vs7c5EBO04ynVRy8jEz+mFL+5/3gMiE1YVgdx/cfKmr
tA+U+bhaDdsoQPuq6oM5KvEjEgGPplEo2WCsDmc/bfPGATl4kHVYgeQniP/b3UXh
3VWIWKoploqV3+Q3zE5iExgnPMrfuKD6bkorD5zREqcEaA/eeVb+R4vuKmPmasYR
+WAZ2DvCeaqTOtX0noUba93arUGudYIGHCx2BkX77wlCXI0eelBOIZzGHpxt40V7
D6hoSL36jTVWOneTJC3PGiBTp7Myz/PxgdtnK3WwamXMdgcCVjokHxQT2QTp9sd2
J8OxpYllVzebvO3EooJDEbs5JfolqixMSx+s0vfeD+djWCffQ0TG0q+tzPeURGHo
kM1k87BVVnzBbQ0wmAmB9P/7mQqe61Gu1SH9/ztEdRln5u51/EOXquLunEMBp4lC
HOCIOlv7csyo+reFEKGuBg3Qjc41ib+O8kaz5FtfjC2+LZaI8KKzC9Pvjvw+lM91
rtnfFyz9d7UGyIJU7KKgZdpTsW0nR/4aZK9zAof32EBJLhCWuvoVlRY6rfQlQk0/
vkI3uQINFG8Kz6BODTHxpqO99kfh4/WGYIjGEACSQuL6tDkAZwcLqDuqdkxGBgcA
bWiG3WJnIyWwYncZ1nrsI9EIxA+zzqRessnpe1zgP/xCWYZ3FuZkGwn3w+Z91Z9S
PV8BISrg80h5uv18m3c8YXhX/CNkPXBU2a4I7kcQ+bGZIbDs3luDNgFJz5go6oh8
QOnKAnPrUHzgAaYku4xZTms4LavVirlx9LS/9+7yq0n9FIzY8CDGDTI0Q2sKhUR+
2DKWDVgipJ9lFqOqE+yrzwFjJYUFo5MF7JH8uTFsjz7xgpjF7vwcVLPxNyenbFrT
ENZME9vpAT1b4UtS3Ld+ChOsYlHE79I27ITEckNIfByh/lqKTPj11ad/VdWX7J9e
LIqCOtWFqVF4tWFXqbZJFUljqF6enmJaGN+41FOiTl0rlsBdRD6RZH54m5K1I42u
RQGt4Mha+ZL3Vwyr9eaGSU4fvULEwu2zcsS0/PS/c7w0EIODt7IuPbNU13AdOLl/
N01RRMuAgEhV6yxGrLVGUD3qrR7zpXsm7GRuLok4wp9+pJjkKiWLwmbp+Iyxix4a
lpwHE4zn60W/ijcGAD3PB2VZdtPBe08VEG/mAZzpcF4IYa5+h0TCT/r/C6XC4WJH
576TQBobf5tsI9IBX7r4DuRwpojPBRShH7ZPrFxA84rQAOS9nxxgUNLPqIzp81op
vs0XIPLYAECJ2QAX4TbEs26WxcHhw5muF/pp3DRFPaRn5gPLrvJ0EWyo15RUKtGP
npiQbYjbsoz7124QlvfklQn44TcxZ8yn3Ibo60KdIq1a1/TgNZikMccKACCGyE0G
5Q+zHOtctBbZo2Wv9Xzjyn5If8tICgQG1VzpJhJ6PBT9xg3dH5QXIa2HEw31IF67
GoxRrAqIPYU25f/hXP2/gv5VCRkke4e8fDDTvSjIwyVtKBKSw/EX0DceHFz5PhLO
WcKlxeQud/lt6r9/CU9Wf29qPQOt2cV2ACFQcFW/pnzF/jKmhg5gFNJ+HS2XcGZA
rVRAbG8yUix2Q8Q9BcyNHkNi5kr3LdJhB7I6fUM//diCJawfv66TuHTYd9OpcLBH
rjjkfB3nS9VA/PfhONBkX+Nz9f26gSTkUKKxFxsSFCY9mnEoi27n0Ero/GtVRu/f
KvVAHbJbj1bTUTv4Gzb2ISOuymqUJvzqIc4dN4dkQ82sNpb+58MIPTOog+5Mc+BK
xXk9nZRdOkW8jEgjWL21WFNRRFO7gBDjUleJIJu822SQBVqGIzIDF3syBdcokiIZ
mdrD87ZkLbBxhE2g+CFndtqjDAY4Dja0pUTQ18R+FhXhzCgiv8oTOjwISp/mO2FX
Ijb3yE/2YN5yU8DLw5QLsONbepR0kRjb9q78JPXH+i+7xmoFXcu0ibLNteGjDx6S
XrPUz++ThSSMz95th/1c9JO/VOLDO4d6ZnILaT7OWpM3/a/eRA3FQNo9QlxBoYOQ
a1yxXQhdQo+y3qFEDRsUSp6nZHOaoQnqKJCAGNuBNTnnUEzJFr75iUPGHhUS6Ze1
ZMqyEjJ4oBRbZf4znc3+vQD49tX2C/XlJ3+VD9BkLd+K7aQNIJRwR8IcjE32QK9u
FK04dyXB0BO58/XOw8xt7KLizzNLvcIUGxz/rzqkqSLpLo9nFXTImeMPsmRWATDz
tV0NxU+ATNaoHkxU0DtWET12dWYvL8ZagZYG+dVUkEDrf6RnyNPw+C6TXs3Orq5K
+CfeXEUHNBvKth9Ucd5WYRkTYbL+N1mB9LklAHVwZaLBF4ZxHM1dhi2M7XUItQfY
0ePyFoaEzHoAlGmWQOtffzA6yJZQsenl1XJZbLijXIFwUsycq0TgrjVwpUZcFdIz
B4OLCXsDf+/FYNpXs1dHNRqLFuuatUnZhUb9yr2UGywDdcHi78k3kJpmanFchdGu
xh6xLGZAg+HSDP1jwE+lxlvpIDp0h/IAXheeqYcjy9NtPIFFIgt89Macfb6xDSuu
FJ3vlWTFP+E3vGkjBIENWVvBIf+a3/ifyLj+QvmVJ0dYJYWt9x1GsjM6krvU26Bw
+PGB24zQSCKzrXYVzlE4O+idFYhb7GNTPN8U22A1mypV0nPqsx/tT7IL9ZK/EYRZ
RDD2UVnhnEI1hxhgvB6PlgYH4ff+bslMM0Gnhh18NjKauLXv9xg4bOmLfrcRdwQZ
7i7SqdiG9Yi/peAbZFFLNeBzKzyDrTBo7hlp17IYx1m79kXh6jzFeWUeWsXob0rD
niGxavWKIfQ10DluR3MnJUlXQg3gwMG4PEizxui+iwj3b6jw52dvRO0uu/hdcqkj
LfNzDlb0VBo9cjMEkdh9o5woq5lpvXnggNuiKaqXBq5R0zIAbCifpjBJKGfqUwxG
2zLhWNJpMOI9N4HYOGc9mpQwJWG5U74QsYKFamRPZtV2Vlm3SUpJTKulqiBP7DCK
7J5BKj055+DbV4ErjCtMxA/G4MTNMFDkXcEJirONlT1Wfb2K1GztbBDxKvBqIpEm
N9Z9M01b6Xz1FD3G7LeDIiFkwDn+8Ba1bJ//ppOCZxD1+Knz6Anc9LnXPjva8g0J
tLU4E7RtEBP3bM3qcyTSpifxyoskxBFlEi+HdRCmYiTjYg1PkurCcNJ316LvhwtM
BvjOOFpBqh15oI440RAq96tGobXO2Rmc2+xsEaq7I8ZeqR/VDBN5I40ur56vqlkm
w6oVWdTbkXaAE201Z9AeCG1cEY0Tv4hiU3dNbzE1bjpj82Fyx75p/kcK6WrPL+vh
U8EtwbS1h9q1Z37nh7BeQjH8L+fIbdaAhcaQB9MTUGT+3js2UR6EFuBW4bvj27UO
IKgG3dG8i6oLspCnkjMOggg3WRNfMADL2qyd2bSDx9NNvnlCkneZaiiYTcHkIkBJ
mPxuP6jQqbfYOGI/g/Lbyluxvdu/JfxCKO+G9dgdTo1tkASESVK8XMH0Rcxo9q2y
bJ2JmHWbnVZZpk3tQRKthN5TaK9g3g/BOnAc0m8Llm3UNN3piwblE5YnDPrjofv5
OwOTGNo5HYJ2lv8YFP6ipT1pm2tAXCdvhPQVSx7chGx8hnsuYYjLujG7z2ZFunJK
vqSW/Q6VjumWqcFEBK3o44quETnGxy00rgbQLAz40fTjh5v3yfvtmbXNQpTk4fJz
UVW3ayqf27XtZfccZHeui7X3J1aAy7LLYv1mGaFloQ01GK0nFh+vmlJTRXS1vp9Z
8ejni010HJm5CPKYgc6Cru7hAde3QhRXc9B+E/dHPh/OXenEzQHughPkR+Pl2S5L
EnkgFlITJlAgQwX9X9LidyaHxNoEdBNoakKcEPVYKXMcP3gD91HX7QxIFk6s/twp
tWxJoonS100gBDnyfCjlT4cs/J7u6V8r1BFVUnxkDk0Fat6pMNnfrGtKXUUDYcN2
cXzd7cMYXUMwyzmuFjlgmEGK68Cty7PFaMwx/9bjME/1oj2kylHK9i5WZXfOhTkH
SXVC8lsk+cnLaKlMugGq0nQ7Kwh8bBGrawBMJ3L+W6IgQvlGPWeoFCB7+V9nWXXf
tg9aie2AzCSSTrSy9Cyj/AzqwHSd2DscVwykXXYuu1qmIpKPY0U7l8p3N/62VGZ9
61ZZXYUTxD0Y/WDJPJd5MCaJH6MeZ2bdOjDg8+5P/jIXOJAnBjhxvkwrFF39AaMO
4z04mqX8M7kcNn5hc28ARn7W/yhrtgnnNilZ6lnlvaqN0GEPMOUy7p55wIO+4ybQ
K5UMgg5UfiJgrdTiE5dw1SW+JpZunCdIriAcquw52U/Nr9M4Xpo1Cn+aqEW3oOXH
9q1ghtS/2XsHzzNWa9xrJ2ALNEce7PHaIYy+Zm58bk3+GmwdIhkDhiY+MDPOJFDO
G5MgRbBX0RJI226YuRG9zQOQBqj/azqZaqf8Z/0NSsyOWoypOg57ynxRYS3zfV73
UqkfUOavQAOw4rtQEo4iPZSokp6S8aBrQZO234UGHHTb1X/nLMJz7Wiwq+4xD/AS
9YbcdbugOw9VDDX18VbZC14nSb9A9mlYBCud73kj6ZnILqUd/weHU+Lr6w2pMZ07
ntXRbQjei23BKYFkKZ1EJitKBBkYSowDJwVFPLAg+qdlFKjhuix1hfY3Cijd8C1k
1cap5mjP2hABPhYteMZNjEUpttR5PL7YfAEiTU/XRcEK9DtVw/GfEFrCfJl430DS
K/wdcnrCqgVtVs5lNEWHE95tXZBg+zggSgRduxFY8n5mFK/wlQKmswzKTZrxJ6oQ
oxeANzdZs2fejAIQy/ynaBtHYAd5CSOdjqWEegxWxckcZtHuXW1/jdqHC9hSXOjf
yfOoeg3eck/SfQWTgEvs4re4+t4CyqtCxe+9GoWtS92fwB1Gzj4ltWiJ8raIUJ8k
UyoOlvCx02HgwQTdK1aGSrJEIftzxZtIBxsJRDeHdReEJWZSykeueMBCMk9D9Wjc
MBjSAqsnFHkDarZKXR2g+bLigaGn9oTgWxkEyhQcL2JPMcRucOr22xNf8DAIkcLG
ahFNI9347OucyIIWD9Bl0IZCpm/diaXtF8gdrP+oaoqSKTtcg31iXzxMIKsfXyFc
cAFkIoI2/OFw1u1DANZBH6SkUY2i69VReC4Gp2c36aKQZzd/iOz6IuxrxramiWfu
EXT2LFK2cVRtpWksNvJeM3IhqB7ztYLbMOmYWMZY4LoYsR9kwPJxwgQp+Hd5c8r3
BmeOdHrCoPpo4OLtskGkCxItv/BDlFrf2RfvRrPDC2dhP9F2pvLV4kaBbO7hVHpy
AXABMP3hCSpjoM2sehKOUS4c0PCFa50d8ZC/Q9UAJsmewKsKqMRTyyxNMOevFltp
U4qkCBShumbO0/J/XJ+ziyUJZa1PiFfgNRlKDzZUnvj9w4kqesW7Rs56y1Jbra+d
39qGvMzN1ha3Lj6/8AGnkz906D6g5n80oqFOmjDPFarD3rF4Fdqs679n9wpw79d/
Sz/EI8AviatiD7gCdSLWEtQK5ozZ4XtrGWZkr7BCdPnB7s/CS8a5D3H5RWBnZScl
O0xcCkzgQ5WLa5UYr8QE242ZHvYyA1H7/RIzen8Cv2PI0f0I4ShHagrTc/1/3sBJ
4q0qtiUCiEHqs29r5dCEHZlXC+DzZFVVRknGn/Kvi/HxNzQMM1PFu2YmX4OiZ/RQ
Fg3GVOz83c4B0IwuB60rRxztQBpTqoFn5gYJqhU/hORnQ5bAboY2qzniUpUh3xrH
YaczExFtY6Q6VC1OY5bRlXAbAcMqNb+GBfTkiqyXhD76vdLdYBMz1FfKH2fi6RWM
slE3ME2KZ1O7I1ZGBRlhfYZq/a+bO69XdTFcRYlTAJOmmdN9BZwVMun9cMRTnZV6
vbnAgamCOwYZHoWyGNIJvisJQ5g0gjrFY91T14AUdt/H1QFXjOiI37rEoYuzdP4D
mkvnBoI5GIu8Oekel3ZbCB7CbrxjMVk10FLQGT6I2reS/zv5iOOyqeI2OG5bOANm
p6ogo1AwhwpxpAulXgdE4XztbRqrqr+W8V6m06yGXmEUdKg79kdAw27kbdhRtsNx
om23a8eIUQS/o5o5b5ZI958AoYwb8kk99pNUBC04kOICuskwuaBaUzxvFY8J7JUO
5kOvE/XgX4Fj3TL6NlGa5F5j90ocHgKQFtORWqfQcxwgb/UVMe1upmqmizaZ9g3+
P96mBxnQtRvx8mTJAB4fqYLyEb6socn/Gfu92u1Zill8XccZ2gYhZ8apbXSV+Kac
Mf0hm/+3aFXcPMuwLREOKz8WTlHtro0w7UFT0RcD6gHzXk+M/RYXobl7U90KayI7
1EiAoNEzBLvyNUTVYDHuCWKFu6AEwhZsUmJ1JMRPO0SG1Zvtu2U0aq6HWZFXY0fq
2CXXDKUvQvHORDr8X0sfhu23sGqKvwrgZr/vsWSIDgXcholbaw/jyC100DVfrNFL
v49gRYv7MQ7k+S9/w9xJ9Lox8TJ+KSQdxsnIAIoZDbklZtgkCVhOTwu4/JpDjhue
6IJ57c+hWn29nUxF/O3i8TBBs2md1xOC095NhgpOxp5mm+3CTrBQZdd7LilDqs0/
oq0IWC+gIUTAEtl3EKPi58Xz8uSORINB/sIoAsXRBYcysUXFv4oLw6hY2zYXz9sU
LK3o0Zj5+CzPCPirHRMbhze8kxpahxJ4blaA5IJ7zrcAkp1kEle6iXVJSJcUf1lG
GV5GCLHBrHyowVihAOun8t3NCllaPM9DxYU+MRiP3c9VSom1JYtSDUuCciRuWQt+
CvTFKhY/TnNO8z3qWpp3rVoISEIJOEAAvr1ARHQvQ1awO60D3YoyJb1oze2fE6bC
jjdd8QijW/+aggqM+f2CgGDAEHeEr7uc5s9n1evclhmhWnM5MEwaCX9DA6pclWlS
/1EZkm7lCUs1mVSFq0leDyzlVKZ25H3OQbyQsNs69M4FRjTzF9CScMdIpWjSrUq0
E+2CYm9Cv7N0tzzL+A66JCdHpryN16oV+QEVKVny6lXaEWk54KbJcLkFTaqVglNo
lfVjY98kd1nF8fu3aUZ6oCd+BVg8Ya7eu/KQ2Jz96FmQQx/tzDsYI0Z3FzvPSksW
iGgdAv92EtAjim56yrTLUoqj1oxUEfbWG850BoiwcrqX04bvUa4J3yl8GeT6a++V
YnLPclLqoutFvvRKEei/Km6DL86HSO18dhqogR+oeSMuoXPrckK2Cm183uF2eqNu
Y6xZu9BkTVrRarjE+yL7pkKOEGO+CeaepbgLB9sELs+znti2Gfcfzy9Z//seViOt
LSzZuSdvRwhlKeFFVuS8mUuGficnXdhNMLP6zGlGMwW2ZHu7yzZeoNdSp2eG9r45
V892yJbWAUZzaoQQU+qYm0HxxDQHzl4Jt5VMJS1JgJsHhAZq6vtojKF6QR8yyOOp
l6BKiJRSErBUFF23o4nO1LSue0rqQo8dGYORnb6c8urMTgV2m5Lta6m7h2KzjpfE
iEyLUdIZpNpGu6acS1ZmSilofRlg4yrp/rIHwV2xbcFX4LxmOb/NkUtVn8LMnpv+
JKKOfS+/qjWu5CIrgtauOeGQ40e1HmOLgstEUDO0VNp5JVu5jy3As8ybYVdixPfG
8YFWO2qs5oFy2xyeF1BE5oFr+GmFlZo4nFvWofZyILUlWv+0gjyr8l4beIOnSYnt
1cAikzmakJbf7tykxkrkb8MwWox0AwYOOQh8hSUCeLgHdFJW3dDmg7RIUEBtlLdI
i1vdYlpTX6qZBQXjidYgesoX+eAE6PIi/QlK3Gc0gYuHPtCmrHFRfahFhwufhMoJ
0NB5gjfI7yrxz57/CtC48DBjor/2DBgwLpcZe3QoP2yCJhDngEGYdRrbGUj7okYr
+pfafqFrHfT+GAPsbJbw+VI//c9URSXMbY0c938M9tYZXOIXgUYsfTNX71rMlQBY
MW6SVSat4caxeUOSa2ECMka9UhsmzedwzIyup5kwzPHPYWWc/8hU+/mPZUSmhpBh
wlKsmAqXEySxFuuvsI8obf+0D+V8mMBWvZOnJFuMJqnQdGEDON0Vt3qbIWUFQEVj
wMVwKb4En9jkfGlSq8erfzW6GEKsHXau+xkq86+EMZ8HyUpE73k9GiCUSY+lULQO
FjxuH+RdDlKaCj8NkaJm6H1wEm5qrMROBfN76ca9iVqzE0gl24ChM2aRXw9wxnxL
Cq6nf9dmeS62L5RnrGmmlIbj9E/trKIECBv2HydI7BgNrCOErkVmzJtw1t6tmATd
s6s841UUOT8W8ODc85jovMMcZfriwLUVTGUoGoOa9PVCMyvmGzhDhH+V7wwRD1mB
RyQPrzir4M5m+faEXqYIwLRoOR8K/vVJODI1CXvzcBaBzeXhzTwq4W/i9MqqXKHw
MM6REvAvQDXZkvg3tGwLFKTO+0nxUSByT2x8Ji22+f8Pue8mesclWYf02m04SUVw
YSRPOebsy4l0V9doQfT+SMOFEmbfUyGv6/wj56rWdy7WTe2bDSVJiBX0KraxHr6P
dLX4zl+cGg3UqIfbuhgfdLOFu1CsxJJ1ZqJ4ZzogMT77aQexXxKW19PdU0CvdAcC
L0WQ+2LerEw1yOTBXwwEFQUVWpc2iTwCJbf+wHZh02wqGk7kAhZaKK5Qmc9cUTvz
ZcenZV3RJrbuwLtQH8EmPifFLJJwsFTXBP0oVisAWV6m8UujuWtcG0cK45EiaEgP
HKRD2pZOxj4kzicKAaJ42SD6NkzhDKhx2TqoO69/xcUlnKYR9TMOPS/+AAf4G10i
huk3p3SObQgGeW/rc1seR+gquCgUe87vbfJSHMuX5sSp4+JVmHLHoiLfLZrcKJ+8
lgD/K9NO4/hLgq3vtRAJHs0BvsjpqViBuc19syASyGyw0AeaA/WmB/UtbET2Qiyt
RgnnUBPFjsxiYD72g+OVwWqmlaVG8g8yLDHTVVduTLeKW0O09GU0K9A212h+oWgh
AjeuqP7ohUlBPRM/0+aAB000zSbimTVDrm4Mrt4qoJ/9WBQXdCsyMQNRijy/mm5k
ojNO/mHaGx7MjKW2wJXpaJCb6nwY6LX/2s1XvkUUay3ZZjNtAWpqFWHlYY8KhbEg
HBZFmTJ8yDzGRnf1aZ+tGZg/9ZI2IMomTWjHwkOVFNP2Dax4joqzKjBaYSKCWFdo
BbqvHUdtwnwMfx/a3Rt+zaF6czP+YULU1kINcMYAmFgPyj7ba1DdOopaY7CzatAn
kELJDREu/mO3shin1gRowbOFB3lA8riUmrr/UoUFvUHsy95l3p7g8dUo5GTw2gYR
7YQRpQt9XoIKDmIxUTOGicg8zvftC7PbRzB3iYdF6ARcofRMqD1brIqywwdji2ZD
1+KnKYNiQL7UQUUK2X8n7QqHZfi2B+LKWB6CYbJF2LysU9yTqfCk0QavD/wlsfPc
jN7es2YJWo3DoI+6rVsGRIKIaFvu9GdCgeFVCeBTWP5vkbTX94V6wziAYi2ZPkNx
ccoqj/lO/z+LZxJjBe7QiACcViZo/YZAJOhK/E4T7kCI8Vwd7HVSNIgBgqLISlbB
a8izqhwhA34DY6XMIG7LIocL67YG9AmRXmKFGCjolwFWB58zbiNIS7CX18JHNJMu
jVjYgq7PnxZCT603wnzWqIckH/v9FYOBmGiLbzM/NulFCFJust9TxqkgfWurG5Za
BVKbNCpNGITrJqqhgyhtVb3PzO68laHVlqu523DiyasA//JMK5z9bxsFxOA/EIJ+
ryF6/onTbXytfvjANab+KTDQeTd3STV4oyn82rWCgQpL0DQHvvN1tskcKdJFztID
HgqnpD+jVQY2H46x3EQW421EsBcRigl7n8z5iCeGnbv3Ca33QM1wNe5WnXJSNko2
hs+kLZ2h5yAnkpikeancgkMFfqfkV+kOLJmvxgdYENxqQ6EcX+5RSctZRZR1U6Lw
7XcuZ1mnbFVlu6gP2NnInTfpZlwxEmFXbCrs2p6VCG3e+r6UDKHjIv6wQ7eRxAuB
W/pD2VC5+LuY++gsoGpWL89Es/+6EbWbn0ou73N7r0bEm4xjcZq563bVxOrV9INl
F26U5k91bwAwRkAkfA0WSi5e2KXHkHCbxUV3Kw+xutctKV7SnnMjG0/p9vPoIg3g
H1HxCg8ZQ+XUkcoqiBK55vnSTLQDRHmXhzj7fBPKldo0CTpoMOlu/D66i5+8q6vj
srSc5oehY6dIobmzUZH3DPLK+p+P3eJH4TA5hoeznF613FU5UzIKFsRs04zd7PrM
uMIGNfdz9GmzN61e0znGeydm6AD4rWr8a1XMIKC/WgMYC+E2f3mSpJaC5GlFBr+G
gymnxdnFBsMB3poHJK6CbmGg6casgl+XbagomRuQUBeTpby/zlT/vI2iqh2xr1ZP
i8EoWkVMs5p5znUG6xZTRfjvO/8T7I8bcvVJpZlmgcc45iVN81rhaTKUq7ACQ9FD
iJRhUrfP0+PzF51UW1TtisRxOZWBYfTzyfOFHAdE8bAhDqLgeSZ7fr9sLoOGpbVz
BvuLyUThr4C8g1FfZShd1XxB8moQ6lQ7r49LRIRp52/67TNwXj/e5TIrm3mN7/io
Cxu33Upyl1cNu1ozU8qG/wf2lRo6FCk3fuycgcZCs3NApbH2jrZJe3xIJ6/RT/fl
MRZ9P8q6FvnBlrmuw+9WgTVcLc7ML7+i2zH6UAZjXTzFvZDjPrDRZ696PpPD0075
2QonXrhurVaccO90W3cNYvyT3nz0Be7ZBOeqBgGlwu0rLHpT7AF0c/1k+67FYI7O
ZrU+XrK87wMAj/pLoBDWkW+L4m7rFnh4ZteAI6ZxuzcXcg97mP02DUzYdjBtyg+8
4/ViRzjMYMy+zsq4Vgvk/hc3er+1VaCgblat22wVn7D/48I3F6mx2rUFZref4EjC
FfpMp/ilFqPUdSBiDSrDQWmffI8g/095gqo5Wngm73w+2fGDc+/wcIkr/A34YdlN
3kjAuc/JVVyIJ4pTULrad4CRdpY7mTgGmlfhR/EY3S+H8lZMXCuvSY3QlmFr3L3T
vfn2xiNE81N4YgfmxQGvz8ksakWLkeMJnpIXiGmmThGLjs0kLYZ7BBuNyLoCl4Yg
UJfEol4QzC3FeGxjudy/Sf+UTiPEZzoDLH8lv+HKO4ShcmsDUl2ZB6WcFb3t4CqK
qaXoDBg96BBpolfZKL8GBDYWo22RukCUa924JmydW5bxfOnSmbC5cI7ZZfhU2+1a
WHlYCNkPxTvX6mCx1vR2EDD23ZERgs+L5OVBpAyqp2XiwAWrute9ho1uIGg0j6vT
Jt3PCYwqNG9PNM+AKNoMSYAG8Wq2zOd8hDgpmrQwqAuFHqYxzNYLt797grJWHi2A
4T/dHWHRqDiGiPA/hIXQyQU5aDYaFCSs21tSSRynt1erGX/OkAbVDLDbg5RFZfgH
vHYSdGvDW0ZIBvHjNtH+s079kI77BftK/GcWfIaXXcAGO/bceVJagE/aMg2bSVg1
MLAEBSUrg+ZMvceX8NZg4ZvJiVwDA2Th4aDGW/sgATBXtDKWfboXTcgBlWuYRRj9
dam6DlLuEo04d+OH3F+MQcdgF1QqYvqQ+swDv4fmKvqRtbbeiggoKKaBoFSF70oY
yFATGISMK/bs7/F+ksyZM5TW+UXE4ZDLHsq/JCGgwU9miE/H1H4PpkYIuZfGI4VF
fzHsoQuX5eejW1CuFGKXenj2oCc5QxF24CNEftXexFaRYA4sHdLpUDWCVIYjFTZt
pSitbKwv9/fraIBTA0YssRoxDb6jRHLIEilFUpQWJsDLuWHUzotNqT9cYc5M8c3f
l1dNbrQmR3b27fszgtd1CKBHS9Hbc28hH8l78ecccciXgGgpK9NbuAkT0EpGAvEO
S8/uxseIx0ALP7gs4/50s4cJpIbv4FbOSe0fdTUihU8AMeIMq/ByJk41ptEUqGVJ
pyOJjvpPYg4i9J2KqvCi50etQvrOnTfARcq5vaehZYFD/DlpUVooZlrlPqXRXAXg
24Kzxd7cZouWWSPYPEzpf8C5y1Fm6cFVOlhaLot8RoC3zNgFSmMDcTUZWOZTlCsf
qpSphVizFv8CQWcJIHpTmEi8SCWoLegDVP2BN2P3L8NY68Y67dDmR+kfprnFfP4k
vw9Bakd43evQ8hoaJdkV3yGcgtM/aUc5JOokByjCz6TMqNady/2fNOOpUR4TDeDL
Og2Gix2IyqkH3x0COvura7Hy6Z/szlkbMEOmA62fU6ur/nZCXMXZJGdmo2RhTcNS
Ux9BlOfzn7npVuZEW+eGdbHoYkO2r4hbUKWfHkfhLZc9NQr+gA1edkcDj4Md6YAP
EY+duR9ZUYMciolzf+SIa5wZjcY6o0BFmSwfEX/W+SxV7XFYE0KvKVTUEYoMy6/W
lthg0AopS2PoBWgvvXVs8q0iUByKUiVMcZeW2EEWO12iVNe//TqIAP48sow/pFQS
+FHwGiwpYbHoWYIoPqdRAzO/UHBTmnlFEYEqI0pw5MytpRBlc7mmomLbzsL0PI7r
iAHP7ZaUXiNTeHMz89toI/eky+nEvLMzkKKSEKf8Sd8PYzC7ocFk39AK/cVbb3i6
wjznyQ1t6KRZm1lo3NvJXN6UNionsCjMMQwbTv2GfDc0sLzMN1elP86xQHznOS/4
wIdjs+H3mFF5YQyafp5REgmX8WP+MPMxRHjAaxn9KwMQTg9zfkINozbJA09qPGqS
y4moCTUZLYQ4zpFGK2t/rnyjL8s+OaPF5QxXQxLS4L6sw/SeW1mbVmsNdiOoSVgr
luRYS8QKS2/LYj1TdtpADkNv1yehv7aZGximFw+Wt9X073cOk9Mnw+6DgjnYz0mF
Dr15z58jSoDUZp5szLS5hp7yoAAMWfYOuIVt0dFPmcABXy7F8nkO/h3jqkfh0wVA
sD0DuBUSdrJ7lDX9+SG8ey2Kcc5gKlXZkJGwj6nK0IzSfzkb5DGRmU9b7JmSU54G
RzhfS3JmbBqUCXRpZp81Qw+tqegYOjbdNKB2GD2uCH47MZjNJ/jvilhOvhmCFWuZ
NJrGDHhzOpe8/vOQ29d9QbNDFkq4J2RJohLXzt8zVi9QfiE/VCFK8+40JCFndSz7
XXypqV1iO9TmurcpWyj0fJRWMhQw0QODGLeFM6Kl7tOkmZ/6EAiAaGfzDvAI06lp
kn8IR77ZARqzx554DOId6t6HawQuvWpbksCtAmh+c/WHdFZlMqrGMhHsggYya2+J
vuH6cS/FexOIfj+sNSXD5LRzmyNQ++G8NL3QB4oWE+VxtTnQTglwarUMZOtdZ67B
wwCo2yFVBfYpaq2PLD9Y1cyX4aDA0aQY54AB5r4+pKgtNHXcQOK2VlNkthjY6uQi
+QBNyY9bGaMKbG7dWbo9tzQ08adCJYpMiyP40NzCIM1LlDibim6koJQcVv92tZKr
UHoP00NvBNTFnTNmKbSzpQI6DZe+/IggOOpqkHk6PiR/pdfHp6LT7Nm+8LqE+9Ne
Cqmnd4QOvwE/pAtSmDJKIVNlmPSzMbdK0pF20spYdFQUcLTYJjI7aUaNre5quKJ0
YUTCAKcTWEpCkuWXSXtJF5wzmepER3WEG8qfd+q9p76fMFFwloFDFDJM3zLdDE6y
pp8lJ2O3uIAKX7ce/Fy5LM5jKtyRmBryOYd0jVTgKa5nUYomvRCkMFlemCyR6T1P
t/G/3SYqvWHxZJa+AfnsXdz+qf3hEyvrkFFEztE7d1hdKemDW0qrBc31usU3WFlU
rJRBqOtqpnx9dbIsEMouE2bR95VBKPZoqeh8Dfoml34pVodazISr5W2PuQpfj9BZ
N4EuMUlsIsKKcJDrckaiW+ZVFxt8Du8qUiQSbL4OHifo8jE+2r9wOR/eEAqqhWA8
Myeta9KAiJp6LJmIBQlVtRWj2ybS9EhAgm+OjE1LW2TaGklePAKqGJqKzS18wD8z
lJ4Fy2vVo57ROaGJHBCOtQrOAXlRJz6k8/vCpd32jahDAmFsYW8jCXDPPbMSeRcf
mKz/P+Za3hK2w4iXGpZDTmxk3dCq0akEB+wgRKFflybYMUAVhUQhhN8YVtawTvA/
Jcug7UOf0u2XzICe+ETDBxDreNFMTzpHlWQXXyAfhNxVLym2xMhJLAmn7955dmji
OS2KNolN9AmI5Sh2QP5snveIJc5Is+OOZjU8shKD5t8/JUaPsD3lwD4VzlSaybxn
HTOUzgKaxnlPgqnZRsV82/9bSh2hHR1jSVFOWzrKAqLpOmBfpFnRFuB1eUQAzS9P
+Q9TrcmEFn9f4HV9Sjvg1/YKjAnUNPEjwD7AX2KkmarzC+Vkvjmr0jVXj6pN3Kj0
mPFixLOxSQ7KdWJzdlgkmnrPIubGss/5eBrQVeqD15N6yWryoPua3/1kV8Iiym3f
PBwIF4oSNMDMHF9aCbpYdP/EPOw7ljfeF/O2E6unX1bCvr4dwWxg0sNcPjJWSCEy
7j2fQuYLKsbOK6SqASEwCEyGGKNl7MzMRicOxK5AlmXf9LEMaQ1UPS1z5tC/IB75
llLTi4txlykXosND9uxdEZXDeLD+/9yH1OeHoCO4a4LJtDMjlOxEVBfiyPzBpfaz
owuD87vwJ00Ghnz2zQf8bD4xfK6IjVe5+9EB56X/wKcgtYwEw/TdRjWr50a6ZcC5
cPbIxzajg/msgBODHP05GzYPeJy5elhaT7ISVMydOkT4u2/icxQQ/hl1U4yGm8V6
TwdSCDhd/JhyGseBtguEBbji9pPy+0pVjI5U7GK3STmH+cpCf7/y/Da7SegQL1jH
C3usqRA8BF0zdAj02XCiBYO6QijSfujpBEHgQNNWGe69d1MDzPx8dp7rkL3bdxyD
530slJwXKFXyEJABzZzoIwp7uqkqyxNZmjcYKchHyqz5gXDw+ZwcGZ9a3hHjjHGi
PqbE8SXCuK5u2nVib0HvtF2sDn/UfHbNwtTIw/g7mjO8cMKxMWGfruXWMrTA5r0q
JsRZIvSjpFbu7WWRX2SkOF2PIh3C7+WHGFFzWUxR9K2ASTMTCuJRn57czdztAJN3
fzqYSFjbzb3kshk1RxgaBdFe6OxzMy1ueaJVqyeIdQJVPmAqg4ohwadcPx2qHGBw
OXyGOwmUbpeZiiu9oq03RvkmoEysUmCwyS43skzzj5y6t3uZx7J7Y51oyeCgHbHm
p+TUI8DZUgEEI0eD0kU8nuamBI1uyupRQ/++PBA8MRIlb8IHQYGtAXpNYFXwaF1X
iGYGjYLOt2yHeCs/2VAdnUnPo88MRdM3K/5Y23rJA5gpI0f6VuGS2Zl4fPP/HAB5
fguyA8SvyFZk224MOSIN6sJFIMma3ieQJzlIziK+bPBbQzCtP5QTQ/V9zVB87EA2
HKdzO4nt+29liA3qPCmGwIVMkjYhvYTuBtPyxXnC0YnG+IJX5VbnYMXfoAZ+lI8f
Y7+pMpMLGbZh5CmvFKECnCvj3CsmfAFiJT3EF5essFR9RKYh6KwkktiZHWmKSq/q
x3BQsgEA09BgK2qq/ozBn2mxzaZoIb6ifT5PuSMScMGVxPX29fJB6aBkQZ76Bpuz
/LPUBAgnD8YXTYvm/ADp5gJR32A8KSvqxh2z8KfrsljtRt+6Ek3mT4GApaOgcdCW
tEgQi28OPaYVNZuFMxclKcB0maQ7C0J3fQuOVfvYZbEtobOyCootcn5r9m4vhuK9
F5PaNpywtoteV5ypFJ0dfo55xQLuhBU8zwu8PNYl8/0MMbbvZ5RFvKkroZNX/eb0
yV/cLCbk9wj+o+8inALWQoXMG+tiR/Qs12H4N5ouZ9bZx7xfTAL7f+RjIoLyWTin
OUtHdm4fMWfynGZylW0uKTSkcIGH7QYJINhmjzrFmawNP3oMLqelQmFQxJmYUr3n
mD6EhO+JUreneLZdlVWDnvVdbzKheNNZp2CJyPKXZ9Wq9erugLgcgnwWnw1sc1uF
nsK54MKoGnnMkfZnJmQTo8hUAQxBODMNUyxAo2wOJqztAqKjQLiG7U64RuHEm6a0
oHPZAqwkJOY8Mk7jUul4UlDeMLyB6fe9wGAN+lbbYpFUZsze08aWa0yyjPg6FWNi
UD05y1xPrFVMCotDHDOJHRuYsp68CaDld24WOlNffqPh+5WGKe1bkGGsd+J7IKVv
Z62ikQ9+8Qqmy/bSiqawz5fQZUm+RT1KkVf6mK5U4coT5HR8JOz/ekm7ovt4jLiJ
TtVi8WGNgKt5Z887LH5LIaa0y+MuzsP1rrATp4v+jIwKvRW+c8L+IZevVSZqjK9u
bkvldxP7JNu5RpBT/HAbUgf7DtWj8Fm8+aON6+/jCIWnv6tGWFTg3mrAvihGW/ha
l1t3FAumjgKikpzc2L9p1sl568gCS92VXQplq4MEPGAzhZKXaLcynBfrlunoU/s2
XSBn4f+INSIaLP4mM+RDYEUiEsOFASz0OJ/hk6Fj+JQaQ0w3Y5aL4mbLaSio+SCx
isGYs6vMH38W2HdqdJ0KqrLoT/SwbrDTzE1sxBRA8cPyHEv781UC7UIrjOHFHHbc
xHvg57XN6i41DWnCdbXIN7M4ob8yGUq5k6CObnQVDOwJK+s2zRbvObUQPyB4Rsvv
Fvc9V1erPl0L9n4bQqBQQxyMIjUNM4mnbDASQAETixYQJ28K6NwQks+XSWI8Ov6s
D6UNjRKQf334mOkyIMMZjdRwIB4kCdlRSon1xjgnuVvHlIFRaxSoqR1/cAxh+7Z0
mAXwSxPhciG0WLr64C/8JxWL+kJlHDv/FKdECyXXHSzCriPWNIxKZXsxvkiRZSWY
qtU5Skg8R1WpxBJPq2lMR9lC0NtTeYUySRDzlryBoYLoBIaPsKcvVlqVzv1c6WuZ
1r/4j64nzLOD8fAUHkHCsK/6F54u3NVTfqts8ohCQpX0jXQ39HYguJ1Rk0cmMpIr
RnYk51iI5OuIV5vb19lIfVgaDZj9TjQpG/FFiRb0UTFsVho8cAxmeFFYcGhsra9a
bwY4VolY/T1qm5NfpUFtkGp2FqjaBCj59U96MFeuojef/JmD1R6mfWvH8fo6imfK
NNxUsgeM93IKYPO4kzioBZmUsoVUTmzv4/pLYU+oGq/1tb4o8vBJDBLHKoS5RBqc
DnWB2J/m40H8RbPAAkdQjlm+B4WPxzcoiE1V7GEduOrIdFpOXKh/PgIPoI4LQwQG
aYLkdShso1U9Bkb2jsfTOevuOi81z3CBlQ5CpyTYFLslKUltNMANYWutNdzs8wi1
slMvCIqfeVx63iicIa0jTq3uIwg/RliNYjpE1Q1muveNkxd+gYU9rvsrKp2k5MwQ
k7tHRvtVtNm26OYKMJFr483TmLjheIr/oWQmw5w7WMO8rCBxedlhVCr5W0B9lyya
jyHSfykKplVU4QwtF1cqHViZJ66jf27ueEBhGbVtA8r1EIeoY4gVowrLFbG63jk0
p17Rtklo/06MpQ4i0bFEkmvgZP2Se9auJd45Fa4LB64bXRTuCqHe4f5qc1I1EyvZ
XIsjxeyL/9YbcL2V9lHd5whSnsFTHCwGLDSsOxlOY8F/YgD1X/GZc3/eZ+b6gzUO
ixbGyGSphSFota+dvAFyrvxmLaPgNm4cKBz3vpvbumrnJjBKC1da3iyPe2iO0NSe
NUdH2FXvdiYEMRkF3EsUUAokus7upUszh+rIIh/fxTfd2PDE5lWvDUi5YcyWoR3P
cBt831kgSltWCcPvp98dSmC+B2mi0wrRALpGO/OS7u9fPqZd6D1jJmaBb6qoZ+Vw
kp0pde//+BLh4jCcQdx0oGB3q9NUgNMsxksW4+w1nTnUTEQpNrYld2OU7yWJctjO
Z2JE47bzsSfANVlT9FTrINwvggWcHg4vBARUTWg95pUUUbep5mmvFLEe1dDaTTvD
q4t38PSQAZd2kjVDWUBHxPAdZKue88+Q7N0lwH1w/OZJbdsiwaRLwPChbXzG3ul0
Xy9VmQnFxt5cBEUKsBnyY+7pnJXCFrZpA8wYDVjbAGfENTN7C7EMImNs7gsUsl5o
iQxgS3MtekMU+FnXmA8X/E4nYzgbCjvvYarWjeq1iY8gDR6RB4VVBiyTfenpZ9ll
nJk0xc/5na6gTqiRWmqSdVwRpdZ8l2dr3bF6+k8+DHleU44hsEwOnRSmjnrw+Xra
7b84pL2kX/w9zDTg46OUXMN/+lZIVw/BtnsMOVstVSLh1fImwS3M5WEbWeO6nqhw
Cb4fofbBZZgxv8r5lKFZt9uFu2dKLRpvNONzqXt1y1oHgWvav5Mcj/1MCZNt7vrA
495Bsuob+sGNakvghyAU7tw4pcAk9xyoBNxAVtiJwuOqHGLfqnSab3Idi1nyOFLr
NHq+JDkL7dFwK6nNaxTy676O/svmAbV+Le7edivxzKhg1+BqyjAFVfA5nRc8meBN
67+k0PTQmbcsVKxGKnknvBb7QYtjm/ocq/uJbBWx8TukqmCJGK27nb+XCoRSAncN
OwjSQgkt7mVarH0qcO1fT4AE2jB7tR13CETPu4gUL/ouI04oRP6+Xst+GOaxLWLL
cmSxTipCOIWmdrT5CXnQiMrdDPD8y0fyl+Cm/1Y717vCiKRoSnGpEfMnj3QHGif6
QB2CuQC61YCwzlylkhbf86UEE1JuNEpXw2rWKA/8jqi7kfO+xJdnP7Jc/vXDPNbF
T8Z1T3ogSB34RXkk18wzvYWeqBgjg9ry7h6nfXGfWy3HWxiF4L1cnL7OY/cUU+OP
Zw3fG9sitaF85GGxPtYeFCtOij+otoeGUslL67viZrNVqvEJtekmFPnauXjoAOIm
MNW9TdIZ4STRB4coA6T7X/z6O0KDb92fcPBzSaPlwlZB4ItMebjbjK87Ys0Q05yX
FtMZE7qfE54UpBiNvng95obQsMHwVvIJretia23GLhuGtXg7Wi3hG6ZOsG2YUeE3
B/TfoiboF5ZawQVLM90xJWZsKzzqspupE1Z63fFvaDPxVgSaLI41fdJQO2uS0qU7
RV+Jdk/QUE0TtLvka4C08hgTH89wMDSU/7BTNtWpAZPLUzq/b68Rgi8eZDkNwe0Y
e5hC6yVUdhqS3K024Cgq/HYomc2/XJAwwPQzaWQ9qU9cKTpXokmvVeYn83vFjShq
7356Nussk/0t68S0xNNRz/NVI+3ihwUbcSIJLUvXLxET4jkZIYQgMgzWza/ZlV4X
Li2PH9rd3i5kmlAOl1XSI4n3U/QQpQnTamVpwaOrVgxfrGG1JU8HdCH+Lbe5dYYE
M4L14HnjkCLgRZPbGTQIAdQe+RDTuwGdE0EN0DIvZ8doH8m6spLldSiDLWcKMxMw
/xCTLnQu/AZW2AtlUjHcnHWlKOQDSdOYLIJm9cm7AkAMPeJXBl1xMDy768OqDYB3
cf834iesglxLJB2U/0kGDEKUBfx5N/q+Fkw4/cl+wIaP4DEv7YT/3FKP1bWzTrwZ
AalhAxIi4Ehx0kqQdee5hSuIV/uy10tieYEUxx0gD71DlUJUdZES6tn7VaDiWpG9
lYulguSr0e8fd+UCtn7yig4jUsN+CFFMYP4g4Yty+IVsEiRTdpetbfRCBqO8yqp0
qHngbbjM3mtkq7EyjF7ny4wJCP3ZZdCjKkWRo/J+NIuBqtQ+TZSBqCVFYdPhqxsj
lqp2CXBJhptSEqoSiDS7p/nZEBleaPfObPGMp+2ko7pmPmZDCkW6/mNsbApCj6EV
jjoaEyTrzyG5EJh5i/LbbbFEXFTwBNwdL1lCZnfldta79r7z5DFjNPGtF9LSimwK
Bc/hi+Td3h5T0jNaq1nsMnAJgPEhA0ULA6XCFOTj0DqK4nlCo5rGusGbGF677oe0
QNjImT/gQQHyofHvQof2qB0GYWFuqL6GtlwjcoEvdwwG6e/Ooo1wT0Le7IjtSQRO
+4WrwArfEmUF0NUD4YyBA4a3oUe3UkESSZ8Gr/oevPCvBSNx+3LsB03Ijd/9Wm7X
reQF1bEI8y65yPOahwh7muKTbc8Fht778GSsO6OQkqh8GS0kPW8ShhVsVlnDEHvq
kVNQrr6APa2/TBSBMLgygUYtVxI/DPfBL1t5iFNa7oD0PI9nBx6AeQ2MZ9KZLeXc
R1xDilT9c8AzsJMbsFQETnU43RUNnYhIY3XAEsgxwr/uHiQh1Jtie+L78OiGGjoi
c7fPHmKpAy3y7C+1F07lDApXOJFl6PQX0iJQImQWnHZ53x3tclYJD9EImXqcDMqH
dDjci/pgXE2+vkapCi34w5V8lggkJ9LXmM4x5KwCreqNkd2vPRlkdV8Ny2VQbqJU
E6cHD+l1EREvrkCum/ZXbFwDAaJrFDEdBElbEFpiex5Pc8bB+GlP/KgYAo9yA2MK
GaONzgreA9cOXLHRZCZ9Lk5LHQuKsUMjMFTJqleiLo8jQ55ICL3TDtN1UxbnRtJ2
Rc4HoZSVfkXoobc4FRcNpXGP+Qb0jzuyLM91hicZh37Sfdm192r3caks9MWEuYBx
e72KO6Tu1Q05SYA47o+BLc68caTzLPJJmSisydcvxd7G1eVYZ98X41EiLmzPyUCd
D54xEBzymzRg/NKH3JOHNvDgdIyVVdZZqdPOqGfhH2WzUp7L4ZYfZ2vP5MBHmTKg
LiU7YUIXDcmmP+dpfM7umfhOpBtggBANuGTzEeNn5mRl8fgyInBf6Ta2VM4RAfX0
jejYkpxJfShn+sJwZfRcFM0qM6uSWax2DqoDPPmV6uUkRLyb5T8h4/wWt/1BxRHW
YOnAVxMOrleAEnceBURFn7pQQmrIoXsAGyZU4iMW1hL7BBn9Wb7XH5T4F/DR/wRs
dhcPQ+7+nvf7J/Zx1cEYAx7zFkO4dtuDVEvHR1QrxGTKU6tun0ikyTANk2d0jXqZ
ZOV07iFwOYnehvGr0n4gpmij9G5wpOo+INRtQ8Q0Mim8w9PaW485aFxOKr/7EsPb
BfLmByRIL6b6lwB0K7uoWqzMLH2hzyl5XbgiobciJXydA5qXPdAvTIZSBhvp+Xi3
UQvYu0TLMCnN5CXu2OGuyEI02h3W8evRy8CEj+H8G4L+oXgU3EzVq011bqrjr8hY
W7SMn8f4B9Br9Bp4/+hnbpCw6uHC3/u+TpdYtM4cdE2wO4LL9D/FTzoNUfvsVrxN
PzsbeqjzBjtD+RbtRGL7QVH2GTW7Tcq8klWe8P4+xtZr3GkUmV+jUvVOQWqm47bD
z7ofdRqaq7Vp2p5JVTjCq/NcwDoqV6vqOUeJ46D3831BD5Us/8YIgm22ki+KWyOh
q5WYB8ZXcZrbiu7/6Hzgq0tdR6hk8JxCfLLJnp6Io+pkN+vfU51ViAg1J1IsSXrd
83AQAlgZzjxjl0YPKNDT3oKGbRjJ3F5nrlcBq4hhYtVmBX2mBnpG/HUFphe7Qd4Y
CDZ0CT6GwbkLiEpi1VxQlPe6cz58+xVLtIfev0Yrh/f0sFM3XA6oOLCUiwzKYum2
Cg2tNh8Y9z2w8Y3uRYWgOm18C6UgJ8+3TRPjqvrPeKqRZRNlq0dg1QaRl5x2gQ4F
rcqImSqidvcqZZH1GXkskTGR7XmEvhNYEQXNJ0fTyU489AkhBltZ0FncTTmmyKig
+9uriNJnFQvv9z20gdaF/ksC6tEKlsXQbn/rg4XY6LypKsJCz8K8XUf7d7K2SKbA
mM0SWCLsHMG2NMRnAoc1rz+Ur/QBYHChm6DJvx1ABhz/XUVu6NfDKdG7vmzHUBUl
/HVJ8TzX1ERmmXuYmFWq//c0FrOf8B/fCLT8S2nqzx+YAX6O6J7X5vvjfb2vyb2c
Gw9ZsSRzu7bQ0wzMfcbX/u9j2OYROBharlButOupuPRiLm0uOg1J5u3x+drnXD/L
dGs4b4+zcChMKxmVXPSph5r0QoCPRXnIW9IWVEk0QsC8FKcaxnMSpJp3Jg0oUlQp
m5i0lY5i99Rpm+JIxU3qHGc+8PaD1h4FhrmBexK6z3hvkCapi9dX2DC50D018lIU
Qv+FTlcmDXdRElqcCFYx8YcTY0ExE1XBHY8d+i9bh7ZSOy4vJmTrBqfyj5SuSxZ4
nLVEQxwmUFIRNfdpKEqWQcghIx8jJtX1Vp0yk/WNHsx02CqckI4hoL0FPSkdLsbR
M+d6Dn42L6IZRqJLND8NaWFmSePMDvCkxw+M1u3gZE0yzdI/HlQhjAZe3EoI18nu
kqcNvUbHkuE53aOdmveKwDzG0un9wWtBHf9nSZyssa8g2vHqAo45YirhuV9tYcrw
5/a3Wl8X68QYo3+LTwOLJvXTs3fGf9bE6AmGROF2xhIEpodonKEhvWtHyrBoldqm
j2C5f6UaNRFN4DLzcTsPwsJO/0LFTy08G+OtzF4qtC47JewYRLrqf5ylcvJ/VG88
kugPLNFJbgvkn2svV0ai390d1gpTi0qstQ8l5EVi2EvfWEKUAhQuklH02Ezel87m
S8CWQtQCf8xzw1/LIU17C5w2hT6D+My/jaCZwjrPfCvLXISTkylrYb9LErI7/2v1
vKSSaZDAtXF1vJOMykktisqPUz07prS+Jrqeb13hoN72fJXaaoii4aWGytTZM4si
QtN6fp33zxckwaBRtWMZz/KfZUFAN6riQkFKc6p0nzyXykOjK7XsbjUenf8uTPcI
SPJLQnD4ynKZIF3WljAy+U+1UZvEB4VkiZnhpISK0rcg3R3iPb1RnGsAMVF2UwJP
XqGiZ5DzIyDJEZ3Z+fLGr2KHFL9i5I9IQQVn4Z74oOlVGgE5C4OcyKBj+SMxn1BR
cpjYU1+KWDy9Eo2KaYgz4Pd30uoYNGxyjIaoGG+8GLp1b4xGHywAoHXB2bChTbdS
h3WsZMSMdDY7NLcYbPnAx8ZcWQD31bazU/lD0GnM5W9xvVj9RJzIe+V4TbIjxEU7
qxjw3+t19sLvsZhHmytF2IDZLWyCL5qpLwXlAyko4GshieLTDfNmbCahFZb3f+L8
8KE9w8FN05Z/d7mevr98L5cAHqCQqSpNT8QemQRUCHeF8Budq2sIEukska28eQTI
M9LHALC/0XzHC+tI153viHPnoqIa9c8aGNEbMrQP9vCc9c+vl1TZee3iZjZ7InDJ
6wrKvhwZvCyDQte0Jq26H9haBQAI7e06GJ9bgFceFCLgrZ2rGlVSgo2gfSgJXbUa
jOzZ2I2ra7/NzuPWt0AyVZIzsgzkc1QrgV211kGiv6OH51F5GrMQLJgzWKLRjWbQ
43H6TrYqZ4P/QMtmpI8faTh3vhBrs8/ROimyvCQLo6JgHreMK3EW14KzEziQWiPj
utDZPPi1QvQgc30RQBYbWB53uILtsT6F/Qb2gZ1YLH+xK+Q4MH578pJeKDdtjkl4
UZcyUhZEOEWFmnrVegiORzms04G5pqqf3/b0LDNGghXQbAaMKjhphAb6igQ5bcd8
8nou0MGHWaxCYnhBqAVjoZbWSLFULV+Jw5f7w7PfWa9gmKc8vNo7h1tIbJNPqelF
SJjYab5wkf6sLUwFt749ly/Zc0SVa8R8Af/16uzgl9uwKD9TzVPG5I0bK+1Vq0/Z
Hqz89zNy3VwnlbxTF3jGC4kmYDFiD8I8G+gVcMbRAO3xaJqwHCBGMFAHliOLbij0
wc13Ox5S8ktHttNUSLPGMsaMzIVaY8ygOz5AMdVhHnzF08XEILek3wOU01QmVmM0
yhXU4cPXOrNtpPN+AdFNcqL4mBSTN41W4ZRIDxhCvMsmXxntXBZrrioKbFlee5gM
IQ8rojNRfl7ff5iRBKrl17TIr1a1kZvaHOGJrys+wjZTZG+/7oSAvyYM7I7vMg4m
evZs4ATDcdJwMTRr3X6DKUBFNAbmlzLBkcjCi8HZLW5NWCAFLKOS4zIWeU0OAT9J
yLlX9IA5pyo0MIg8iRrPp+0XJLUZOyp6IkJbp6m0if49VpnvOIdBTTHJ4Ahw9MzR
fNuD7TmVZhjHwym59Aae4O6dKGgjq/LvStq+zTy4GXT/o2fmOJieOVtmD/xgIiuC
+6MkEwKhWu87UlPfMHvqPzr2UZwd3K2S707ovCMPjwKvsdZKtwR6hJK3JQDiEdxt
tsiETQ/1nWtHF1ixOm4NmhP5nrVOvmCObsNgQAziSVSSTcOp+pOd6hdQWT4wvMx8
F+TOGxGDvKJh/U81L0uXc6Hy8RY/S+ozNEiX9SXQL1+Hxz8hoFCUqo4V2UEjEMRm
VoEWmmer9f4cQ4paPs5Otiu2NBrkEzwBlC3h2+v6vHKa0FzBHlL947vL9g4scpuR
HQi4LZ129WRy2z/SuL660xuSXSurmTDdRjk1LJWRgtn1OD4Ky/W5hVSxW4bL6BzQ
UCIfjuG3YsMMyMHZlRwzUkJIgmrFlrIDzojIEykltPXMRptgpdRzcXHji8kjvRKo
qJ6FkdBa71IIae29SdEkaEJL9wefCatPsoqZb5wCWBCQTkDQqJNoOuQ6S6+syi1X
ig2emgPSw5S9W5L23MbnVnHpd6zHRK2dL7Hk2f91ag+hjbiQKmnD3xlpmoFrl3kL
QISLX68wXsp+6V0xgXEFUrrglFQ8GW40I5/fukUdj1WSkGuBMhwlfRxXcsshxBB3
a2UXhYlEk0+QoMdH2zFS5/VyYa6oBOGuFB5rzZvTwfU14gtk1Hrcqm8wr5cY2meH
IJYXprRMSckAIPPtWlxc9WW1RHDsmTOy8j6JOJzjMBMf/vCblbvqkrydu/hDteup
rLkW9mbY5LUxRGGVmxpHGf+EJScB2SyWHCcYuxcxS5Jn0LimrIdeVG1s2sAORfSt
iZVlnLfnQTVFTsVn/zJM+wF4k8mQL/Mx3oJEfUyXOYpKundbhaclGEgWpKRNnUOt
GvDgKEx3JI4uufNW7kd1s6+5YjpPGNr6P/BT9TteJV0F+WxDRneN92OSlakY56Rq
FCFioU6cSInkxIwzu3ufIRo97F90urxziJPg392WQ1Pn34Ro0sI+OvmUfJuMqmhU
M6PbLT5mMFa/cFBUeqjjY5lsND4NeIVDZm9JSmatYnGle5u0FLRDBHtNB+UznGRu
43g6wsj+1M8YgQc7CGs7W+d2rN74IeW7Kx8j5l0HSSz/6WbxMhhIm7eB5KYKP7Cq
IBeGnyyKwDgJbKFNwJiZPXWYh6BITNWpzoxv6zSBHTkTtSW3310Y8TMjdmRGy0rx
NipdlTDoEl7DRAh2shGPwL82rx8BkX9L6M85VX69bG24krU+1/vN/FphJ/xpr2qe
fK2pHtdRhjUgJuAzdn+JRlVH8tvRA9uLXHJfjZeNkdtXIVCLVJ4QE7SIEJgJo5HD
fC6uEwWGhOBvMTuOzfspIifHx1hxPfkBMDjxdpvrlbEcALLMqzpl+2Pl1bCOnVXa
hOt6yY5mBW6gW1d86GasQciVe0sLBlmKtmr9Arbu3DzGL3qAlXo82GeymJ1IIhUK
5YguEYivzN/y0oa+VK3QOK0HAfPIjeR01uoIoF7xAJ7VMhs6vHUzD3nAOMomQyWM
RTqFCAI3TAWLUwUK8UJnROLJe+9xun5cSub0UvWmXCCgxMDfDRcD0BB7MZnqtyzZ
eEokJEs3ay4vCVxSINzsYciR8PgRVVXl9cwnTCzejLddYJNYRQHWwqiebX8wYUUs
6nrrHg6dP4FAp1497N4awebyKJGaGAUQAfR+qhzTB4Na3QFtQkSwcclCHa6WwCtd
AzQlyOxN7WTTq/eyNtRT97kB2MOqoPeRGunJ5GQ88/NTHMpCJz3KVEbZjvS6GjSu
P/DetqeRiXfFyfpluylUDwsjLlDb6atcgKDHaWDMN+MnT2MZqiKn/sL8pql29/7S
cpmrN8rgmIu2lSq6M7QkdAEU2XF+w0hjTNKKwj5h4GoMtfoiPDjL6R+TxUVoJ+6x
MHEeK/LlE+SEvcalFOItyzj1PSuIC+k8wul9z+C1PUhkYiGuqSvNpuIVCVQj2cig
sc17pIqbCQmdU7Rcn+KjAzaEhqC0n4z4ABmUd7Ase5po9HnCRKf2OYyVo36UWGcv
0ALe5Mmn707QAIihTyMIHMV19HerXu+cR5XSU6HN4G+2t5EPk+CC8akqE1Amzd1v
sElY7tpMmmyNfaOw2NyizRvk1Q8kWXDaSWMXZg3oD1AlDITBuVsyOO1hIQx2uWjp
Enrff0GN4uPGGKrP8BUBrbnXWBobgOZljq8Jd+RocWUELFymtoYW89GKp/vZSBVn
RAD/Mp3MAX/kH44M0m3nzL5r9hAjv6W07OpUyBpJ4AHecdicD0kuFjkKIN1y05T8
A8uj7qiTXwU+wnGfE0TiLse3vuo1E7+/4hwMBgkv/0P9nX8ltdFuyYnNbMHS6PTs
T/h8XI9wi0P1YRKlUGdhEvaSBOUuvvJMvTzM5XlteTSMQ75XBOKMt7WDW0AUr/nh
KcL/pUm9yMZeR+SU+8ICkuztHwtXQJh6qHhdA1eQ6rY/udRxo8YvqviksP9dug+t
OPf+ZjXZtBJs7WhGdPDRwFjcwwFJstSR4Anl5UG8uVeC636M/nYmtTI89XL69j/S
YyrSQLoiz8dTZNldQS1kdH6snQdNd2Q7l6dkJ2r0uEgjI8zMOmDek904jnZwPbZJ
/p0kQNF+rncbFsEyWah+xV/yvUGSP5R+vA1LaT5BefUPmyMu/+HKgDP79d5srSj9
wUZZejnIS3VU3wfrM+fY8RG8f4MTKc2lPdGwJV8SOINRsEvBoG5z7MvMnkBl3jmk
IeE4BY09XaEyjho2bT0xZvLBn7zlwEgJ4xhsXIv46zzEMc/dbCn49R59OyRaRaeB
ecnz4BAWdg7PdrRAWwontTBUYCK7FMbSsrNcnoVwwHDrLo+wqB77GvqWH+PkgLBY
5RoDhZBDAizTlFVuXH0gZOJ6HDMNsJbGKZz0dr8pVNNaD4E3ilY7pMusFyicSz8g
y2LHEnAK4bVEy3KNNudJbjtFolvHKLB3qWgsvcUuwcG9k4/E9/unCw0i3jH6SuSG
Ot9oQFoIJI2wHtQfbNbgY4qhvvZQvY0K/PzHQe24zOQrY7CINfr8yrVbfPNj9RH5
hHWRDH1N/0GxhPrIvr++c7d7Gk9cQJnAU+fnO+GlTi7D30xajoVdiqfX5ymui4Ru
Ze7KfaY3Yx6/1TaCfrMpMKJ98x+yHRbkdS2T1VNIla+osw4jQVFV6H3Mpcm849h3
BHY9rrXDf4OtdIBfHGSWLAd1oZIKvMZWD57RVtuHck78sF6k/it+ty+n6OFVw2t0
Z9AqIgcrIzfdnMB75q/YaRMFNNdRCHQj4a14WLLV91z0gdZyWaGpDK6qNpahnfzu
Z9dR8tYSOQeZtFTareVr53fWUyS5ykqC9mPCPdwxWJ4fFPx5UOudVdbVwUc4TV0H
OGjl7dn5HZ19oNCrrEqPcF5QHsebvbj08NEgJpCwU5s3RqIaV79n5/Jy7NottEpi
g/D98g0xdNFha9PEiCYPY+HB3hHSgrHRaCBzc0C/FFHjq8+huDKMjZeLYB0Jvvk0
rzwfTJOuE9Z5fP33zlG00hs3yMi9QjblrhDSMqVk76NFsvm3xCDx1hTqNgLfE5FY
+rTaRXfEGS0DnziBGRhAfaZmTqlqers9oeKky7UvzWB8TD3cUZFaoUroq/VM/XzU
4zdsySui3xKxv1Y9F8ndNY95LA3Oz5n8l+idtef5jiTYWT3s7DEPk0Il18iUjXTE
Svahu98CEB6YUs1m36eu90nG3TwXb0ORgIt/wF7hssvQgLVkKldZRoN3GjQYLGHS
o0EoksBGejIgWNzz1gmniL2lOGYtLsXDjD3dFasJU8RdgZzdC/Z6ehiJX3lt40xk
G7C1wceI3s737iWSqSNpeoQMe0w0wWhkdMCwVYUdPK/HbVtmjfSbNEIwRHp2DXZ3
Nm+cPU5Nd26gPE4GTg7nRCg6MzlT0KLxV0vQcjzJBQtEqZmNgFE5IX8O7toaJ4VU
Nm60iwjTDTS3ATxFqk9A+HNgWim8wH2/8CX0mFz8YUHhkDJEjSGu2DMtWiV1clIA
xNAr6Nx3Re1mtsl84XHPAaEd6d7jd5L4Rz+9MEQ5o11bLXOrSAAbY+yzDdMkSQmY
UvdqXRMI7qMpSi95r5R0ANgmSfjwsxLWWZ7OXShwkGDbIHA843Wiz2TJuLrp0klr
lDRVTQad+EzG1jZ9nzZtawlEa7E/tO/VUjOczCNiIZwGMsTVugtxKlnwZ5UiArJ2
mghf/TW5lO3/s2cgYtDHImm3c/umVzShwIHfdByTzV/+HOeWFJRLrZXPyqSO2iVa
OVOCOJ/2p480uXxqfUZYzd0sxyiW7YLouEpznsiffgiLxLlDaOsCuTvWHbmvWnYV
96RwGOjRcedBwIss/mL+/LmEPdHfLSBvEkz16+3jiucnNkhpO3J8Q3+HGhvL/76n
paSH2lEixrsNqVfez9+YPuCPCT+Em0UwYqV9ka/ploI4hcHI1rZ6viNWpGbBvKJv
OZWsjLAAs41LW5AnyUgswI3HV+vPDFgl1RrYT95GkR2nwdBztPsnmhGl5j44uW5Y
K11hnqFy7E6g42C9oYUoUcbMLVJvg2YEoNKTOZ6HB7yzSdszGLF8coP5QhqGOSrx
Kv2ABd+3IZWViYHrybygy+GmRWbzrzO3RZakcuKDqoZQcHIaIEEi7WUaT16e0orA
/A0Nb0HpaIxzkfnd/qa0+v6EB2c96KNCdKndin/xsB9njcbKS2ffD9jXYoKL7u8K
Nv6NEBvVf9dhynm/XftEgc7Z+MDh8MtTqlbPrRJKoSHJuMijqqZ1ZNC6+q090jz7
Hv9/ikC8Pj/mGnSnXlKatnqpa0LW/qfUJhCQrHJbg5GnFrcVVTBgXqJ3Hsoo9mrH
NeamWUcaG77HwjKil1uSLyhbwYh7vyU/wd27gzBbjBlXqTzXP+yw7g2Ls7ndsutW
r2AXy/zdpjE0wBrMibH5TqzX0SmI9facf36lmnxOzxNnhLzg0ex5RUV0L9hhwOmT
9ZRe6ey5OUnQ/adDO6yxjVAtVcVm0j35AAOhTVaeuh2BnxyRT9P6pV4i9GG8U5ea
HRTwUtm1/tZz/xUj/SogmMd1vS/UYresaZTGcfd66nm1K8WgIjLva5sLLWxvjXnG
STEKKxTBoXGjCWyNhVbAEh4RUNUDSugfsLJEMFKe8X1VCeYTMqQydVeTd+dOn0kX
QcLQk7oHvYqdr02jIwDk5wSBp0a3ejHxwxXaGWINr4uDRyV7aLG85Kwvf6eRRTbq
223nW6oJrRzTeVQFok6jZqIexEnHwNia40yKiqi8oGYro3XWUM0FE9zFZ8E5Yds8
4jTKFkROhARtJvd3cuRWdwu2fWEyubBueSj5Rf+E0ENHNSZ1CphMZRHpOHDcQB/t
c4DONm2YdapseBBm9f7csvVsz6OKLhvVhxGNS6CM2MLdvMdzHoJQ5xGNzjWXVBFZ
zv9nUgqqhPwgfsVXYymGmamzgh9etQg7+SjqtZxqmL7JEpjX9OVhjHbQkuK2OAhb
gTEzXaDv95BGf2MR57N0KSQP3CN/6Oqc6hwpyEBw7fAf6w/QQ9+zVF2mkaAwZ/FI
ai/fYnY2NGbLJ+bk3xS9/VhFkhuWy9BA7IFDNvOt4mUsiORCdTuFWIh8Sqr1dWpT
6o/D6x8szXbqQu6DIeOAA9hvrp3ELwgOoQzCMqhg2PA5tiflfrr3Su815sKMzomM
BCSXeM2ivtly1AHBDig+wHw8FXR8P5Jmu/i0meAOkRo04ksA7QiNLfG89CIvPxT6
veMV4NZptVwILZWw/AhmiHS3cvJtT0Af6LxAbURBjay2f3d9mpOZhabrpuiddp/E
nQX+zomDP9yAc3Wf6Eb1gS72ZYEBBLUe7PDODk+bP7ZWeoNbCpHoA9/5qAqhKzrU
gcXGiT3LO8EeLpfMRg1+1UXA7ujWM9rmAF+SSpg3u7vTvLuijUNBHr76tObaZedO
vihcJpk8endA6k3uDb6Iv7jNYxjG3zpy3DRHzVQSZ26Z7AOy/L2OGV4K4HAGJvx6
iONYR5b1aGcquxcUMYdewbYk6BCixUu0hJRVeg3P7qCHQLWFhJcv8Oxh4i4IpFdm
y7EANKRQjPzVuLaHGbc25E6IArWDShHtxtaT3znRvo1zwNV1lLr9z1ssArkVG7uJ
AXmj5BKMt8nCJAFCoiOO2pBNOqvHHluuCPFYrJgiVKkc0GQyUtnx12wOnheXX74k
QqIdAI8wwo09XUXCXkLli9fMHrUHzoATQqc5EpsCFw/NVRWTFWCza41DT1+Oo0vC
0oPxgBL6sFTE21MIiWpA1ZKGDnI+WyTTbQwhQ5a8TxBihA4Mtw/OdR1W98UY498p
w/r1AtUuIJUbSV8CdXlHXsxxpg0GQoZ6D2xeGc91zHOM98VciomaaUoQhGgkUF+d
jTn+CNIMLqVGg+hqZAA65Se1WoTgPJT3wbjZKLcE0inkVebt4jwV9peILtOS6DAC
+TEk/j5lwOQI/fPHaNa1Vv2Oxf/wIUT74WgwrPHuBImMX9pRMW0vwIKMvO+zyDYd
wKd1/VEZdZ6QCbamM2fHCPRSsXxQLplOq9yqleT0T2RRfxFSBmL9bCaAp4fSruE5
p10nRBDjP7khRh4VofEZuq5uMzmozFtAydBnJ/yCgvCtAd01BT3Bf0qJ+qyF4rhj
1Tgw098xvDs3HXIf5bdhHVJMww5Oyq2lVGV4gdFBHGqPzATEZ6lffN09mObaWy0p
u7f9cv1qMFT/sCh2zCnZTbWkv099GlzbeqJvBLwwwixczfR+GKvpeH6rVHHzx9Vu
hEenUbg3mhwLMsiK+R09jSyZjOqUd0Jzp8OWpRmcYAZQr53IWbuHVTZE+CAlQaGs
l2ZP5GsNHAYMgSAXDoUk48p7MhqaTrqVS4S4KNGCOJMtZbvwcaioJw4YcH1V7WIF
cfjonXg8RUO6vxTFmjteXzeeHyalxTLVYR3uTnSRHwyx1I4pNGv6yaffq8U+/paP
twinbdun5Tq25xtBGyVG2obIFj3achkqRF0ohYDSZ0KezexvHotBbKEZ3xzN3kPM
s1zNA/M6mSv1DnjpxChQ8BvT0mPv5eUdZIocufXDIdi1GW/jS1luvPsLZdGZB5e4
PVAm78vp9pe7UJ3YjI4AcpBXvjIePcknCVZEeXenQJ56HmjiYfhLpboFKNdoxYy3
qpBJF7leaMDyQh3GR2DiQ578rgVXaSLZ2Sx1Lcnf1O66QrYADIdXjS23ppqttgNf
Yst0dAoebxk/2GeRrIOiFcPgCsi0f1GATiKC4RnI4XOz/9NcObOnocuYIFRQU5rF
G1cBxAsyj0R3S1Z1FspDyZCVfR9/iY2vnZoMBqfHDF/817Nh8BjxpC3174jg1yr/
YhIZzEhKeIVv3Wnwq7/O6FUKKhfvFEdIOyLcP9S1dUTtJlBlwk9R6MBLweeYaVRi
wtTEfFqhn3IVijSpLq59QHy113LGMzb1yXA3uxoq3h5mYXKhiUi8tbFlv1AyymZ+
JnFhERUzPVcLCSvHkfY/aVyAaMZl7vmtXsiOUtV1SwgXLDUxhJib5m3uRcg/gDsV
wZuq0g6NAZZ7kooxqefohmOXCq5QK5yN3olL57kZRbiEiX41Mm3FzgdwFR6RoUOr
fNb3YXgE2k0ZtfpqzTgnJWQaxwl8MjOk/vJGr8+VzpFNiXxjjuvwUhUiLIHsgW9U
x/8lEUnGlnS3hQfU/U3oUluUmVzU3IlK5YEqnw9vZIulPH6N8F9Mn4/cob/Lmfa1
5JoD34xXGLssAd7hkhEh2jNpkeKU+zPLZQ0DgP+ck1m1Ky3I11oVME9W7tuChKKT
aJSHVFtK3LKirBmuX/X7zp/E7QmhCDH+qLlq4AD8Io2BphXIAiYsQJGsCRtsGQ7K
3eNJi+QhqQ+PM3Kowkgkw75Ma9Yx2w6trozfLhTAJYdc6cxRbrhmmPs/oJpkmCxg
/2wQyxuVM4OPazisVTW/8khTHs9uLZx9tJtk2u/hYdfIyFm+N5eAJiAOXP/lshwX
ouPdVXL0DKgW/2ON/vQctadGG8WBGlv/UApx3aTywE+Xo+HKMurt7n0NbpcXgsZa
k25hreLsu6BP8kgbv6736Su5fajCYNfFKymJnik491zZRkhrry/tu8b25Xinmmlv
1qOlhal8FlIMLTMHjsYoiabqo2KDFVkf1jY1TmjX1C8QpWEoIexTCSPzSMyh3NTp
CWRdO6B7dunlOknTXFYdzoOrJ8An+r8ciZu2BlrtAJImCCfCFyzCRA9jdOcAY27e
Qkh7he/CuqsSBSWXWOui9XVZE4O4FqqRV131937DgcK7yseyyq1V1ZwtX0ummjd4
YxzIFtgp7yND/Hp9AAcAi1vJJ9wAAnFDIZmzij21XUzn+Y3gzRALyFBipwxhs+Dq
BIWUCCGaD1mAkZThkVJE+C0I4GgGwg2qTY0SY3j51NHSRaDbxhDkCizNe+/bgdYM
UJ11AYIUEBiJ9ATAREbM3r3PS1/fWiyXPWQdnzfFcltIn6CyfgBt5rAZAV9Fuaya
DM72cnb7qv4n4YHBMhZnwzUdj/KehJXB6b3tZtbDM2iSudqbeGOPLlW/3TAWC8ul
BdV0wgAGsfa+K5tD5gd1PoyrOCHB2WvZNE/ZBRT+oFj6ezsPamW/Sx82Sc+kWet7
1tyi9hK6pdD/JPPBxpUAvGN21KJoD+lyh6uQLSV06PGIUU8q+T+CzESW6Z+/yL1Q
g9jVwLIZ8kwFm+4lDYmYBuepVC/iMdiyfT6fcPLJkqz+7ppZlYihfbSGCXnt0czR
UnfU0Jh1IALh1U5rl6Wws1F3UbtLSrzU4OFXS0fyjV0dKnpeHTti9gONvYv4yUY4
Zmau6mAhOVsXwF0cwOgDCEeVSD8WyiWrcAm0PznrARHNBqCaddxfdNAzdHuog2ro
P6dv/5pWhnas3yDmnE7KEXxsinj4j0rAVbu0noMyMQIpao8qJK/D7m+zSpIVjH7M
PxxlMCYOP9KpxaNbekEx1ix8tsu+1o2+8oDV4XIoU5qWXGmVooU9BR7Lxa22GmSN
xhukw46dUwH3GMipS6ZTvk20xNAjnhOiJwceCFnJQVvZw7fwCT7V+eyXjp0Hqem3
dNyvq3Wh+VJrNwQj9nOj6scLNWhOXGWqWuwuw6RisXm9zoe/FrBH7cer40jAKgcV
4XIt/O+uVcemygLjiRgqienY0QFRjdJPxEXexlCTvPQdOvoBA1Tmmq7pIU2/C4JG
uHgAFlj732lbomjc5uA6sr64K7QlXfwGkLLF+W4mroWTH+bdmsO0S+ehhrq9WVpz
sx+2tOtqEBC+Et1udM1NuEZYJvke+ejTpf9kjxHK7/++NT/At/gYOEBfJFBArz0m
5tt6AumFbh44VRrypN6oKZIMZmeqAhKPZYynx4LRFmQ5w70qry+lDtUEkHV4qe/r
zR3BfqzCRBvJPQormGZlD62Sq0uVCqo15orHRgMGrfL3fC5B7QpkD43Z/ru6qLmd
5wxzguvBUj/t8cr0CTnHBtzvvVzARA/cFY5hmtkpUzTujWn4fDBKu9S/QB+QGo9r
UMaGn8BVJo8PqhY4V7jTi8yzl8JT3CULJmtxxpYQkJQXHRM4h/2LUB1W84pEQnV7
Vtlml0ft0u2M4RE94p2Nf8blhsYccRuCSLCS7BpB5PVf9RyyyyKwdwxW/j2EjwfL
vKKrHMxxO3qPdOJU5NtQtGwo4Gj1NSo+2h/qQTmVwrgn8igDZeplOgPWTMzX/Pee
NZ5g2gzeXEuH91oK0kEDV+kwia4kfVNMCReGjoPFb/eV5Us3ZgXrhaZknnEFohYk
gHjBJeknzd4BCZr0j7kVAWZspHDyDO36RZMwybO26qeauM34z8Wnh7UtYuMrzVCZ
T5VuHf6Xfbqhu0+YL5LsIk40QjtDN9dPJmbSRzgtTvQRrUYiOc+9LDrnKdzYc1i4
qHL6mvTQk4UQuHDiTD/linUc9MxNq8Ye9AW2hbgVaYZ9DNd2/DZEFnzjgPXt0JwC
YptKYYhlfvdGTWWRX7+2HIxV7GGL8NaQrq382iO1XqmhJuCg04gOJm0G3NBD91pI
O3p+Mt8QV71pU8bwZzb+syhRV0OxtFkAGBZ2f73+0FezLS0RhnAFLM9YpTE4mX3F
uJ2RNvlGcc1EfG03tJZWyFGSg+qdLdEwAKEJc8V5MTqdMB6Mpm9dKXKd/GjwL5p3
pvog8pO8MRpaijO/qdgHEgaA9PmV+i7M6VKs7vtTpmNWc9nwHSeHmvwZ4GdEZayO
LPkkpbWJxRh1xxI6P7IPFhI7SRjyrXcXBYeXQNMG2tRahmnUdrlOrrSs2sQIkrv5
TGsYLxXa9vqCMFTwOlYWIwYd0eo2A0ufxekIPIytFuPL6HozaRTdIitycwVDhB+1
Pll4Gq/45r6YAjL5sR62NVzKsNDfYT/QBTSjKXZbjNzVCUr/DssQsfzoAqgZOJ5L
w4d33ptD2ItuHngh2sub7WtBGSage40AK6rcryyjOFjz+EUVTuE0JDm73lSU2RuQ
Wf+JfFiFz7/cp9werXr+8zlQX4HoB2/RLCBIcXYAJbwL48g2LuyFs9YJxBxct7oU
e4uZCAsigl8s+zsRhL3RW8l58NBQNZoANATY9XgkKQseeHwewBcQNRRFOmq+xUiJ
wtD1KyaLntuOa370RTH9bQhc0V7dEnjHzQ0QaB0QFgafLdSRkwGWEXoKzu69jzYt
ofT6zimMWzb/k0qQR9idAu3tibW87bZCvUNnD1EHVdC2iFtm7Qa/cKIpkwPCfNRq
YGnlzVp+YDzfDwslpq+AeZi8+2b4FgfFzPo0hnPHhtxYlm4M66p5+EbHbUNOnvJ3
ghmHg0rHI2Q2o6Xx8JDJ2bQuPbbf+3elBofuDnAvNSZMHf/bfbg+jVM5zMtiNv4n
SBDYrzMBsDiqwjBKgg54NkuyOtwQdLPAPc2mL0E3/vO6ZpXC46TRwvZ26GVdIYHG
eI8zgy8FasHp5OpgGngCzMlp2hHO03pHA3M/uoZpbr71t5Z31ctxKE+t9i0FRDYS
pJN91IV6x4zCqGITahZGNg2nQjWI1BVvf3vtgtO2a+15Z/Sk1x7la2qbjuHsjmMV
2v2d86AGw0X1gN9BQbbmwN05NLejN7zAuaLt5uYsyXh40rOKQbHuKMk8PyO92Iy7
2x3Ys2b1wJivsCkI05kXyvQbzmdXrLFR5muCo9ctmI40XDfPidouDh2rU3IDGw9O
OaoKC5qGCqSQYl2W9AJ1XkcCUn9r8SncJoCpFEMW3o9TPQWD30QDsqpL/qJoNzG0
aRNImPtSM+vQrLgLoF7EzqrbDJh/XST7VauIeOHnK7qTwuLaYpFrE1kL+uz+UrrD
ziwH8dT1EVyPBnHJJj44p7EwE+p4iMepP+dn5sd5I1jv60wgGzEL2R4Psa+tp5so
UByjX9XlzBNpxmgWdiGo1PbxAsxDCwEpMN8p0+bfUNzHtJSR7UUC2ofxwITZrj4w
ipCMmUrXcxlm4Cennu04F0P3lNXp/i7Tk41LqhZR0L22wnbeYwane1Q9PjsW5Tgj
CoOV174b9/K7AgtW10+MJhGHhEg3BVtIqIRJHDYkGPoW/8ONRakNDmqskm7blvpC
YZ7e7jA56fgdcC7ehBsWC/ewxYGZgT6Nh4lWr+hCef40NqkPt/hjCGjTLkuJ6AR4
wJ3kBUyoCdPv+h5GSCNVlL3pnvwNJ3bPU0mPgXA6yMrEe0Qfnjr69jrh5lT2z1oa
8XDRevFb7sK59+9dAeOgZy4z5wh5eTP3TRaL1rF/gzPXcReoAx7MhtIerUhJD9CC
dPEJsjTLG8xD3ItX59i/mGqByR5DqTULlVFnWh72Htp9jBNfRUTg8NB0NaYr6AET
hi9oZvqxxN7I+VILRktt3tNrOIkacpv8MYtECMY3BWY6o16cf/jyjt6CKif/0L4d
4Dg/UNQIHC5/2jqVWrDSswC01z8yNyeGA24GDn0Q6Rqw0V7yStc9/kvD6rKlI5Xa
zK8So2wZVFCT2JJJ+UY6NHkRAziAEON03UiD37jjaN/I9gcpQFWXjXRuRyZU9z6j
pRXyur6ql2mLEkLbzI8HvE55a58oBpsVlYbTenQ66kPn7K6jrNlKvD//I80BLDSa
9Di+80uv2i4Ln/rsn46ZcU+J7A2w6u+Cwrp34rgaFkAUfhdrnwqzL5jcTT0mtHqb
mArkThuSc1Aa0diuJL1IN4GlJeWtRrGa3fJDXnZ6hIE4grOWOxW1p85oiC1estGp
1R0tNmTqisMhUyo/hSgBacRDulhMYaOk1uvcWYmRc2XiU5+aUHL6O/J8NLwyNMh2
QmJm4AQ4QP33H9iLRlBWtifiqpvdt5WWrWa0gQlZwO51fiqKUt4sATlAW8vkKrZe
EgUru7SKcc7wOKR5b+nGIeeR7P+tzFvVTFpSKIRD9ra8T8pQNuDmcooy0jI2n2YL
YUTUihons8zk6wIZ6rQqg1j6rj7fNYb4oE7epHjplkc2ryM03I6gsqTiAnUXtI19
UFXxZsWnFeuIhaf8M4sPeGy5bkJaZwy5aNi5URf9zqOvyA8QYpZgj6/EM477KSvo
bKETmJQevnE8w/trQQkitUBmTSo9UjFraxAoYP6KV1sYwfG1KF3sqrFdQKTKLGIg
6rL25qMJZL1HLuy14CExTN/NbW9Cu93AfnslCDK4k5oGUkQxrBX2yntSUNJdkclx
BSV6DrqUEs1TbG6iOpb45DaA/7QpzBm3OZkxl3w31rEvjGASSueIH3JY1cxCVw9V
LLZjwZgAgjTgaVmilLt7hv/+0LWCr8UCJW96PCBsSy02fijZTio8adRRYV3je++l
SGKQDIpGQ6jvI6ET83SHHgGSTadPCWRMWtDnHp6VBa+5BvcMUSmM7kMqfL1kx6lu
N1kfx2eYFGUFSHzy9o8zOU/vKjlLZ1xL7xKL70dngncsm7YpSkrsWMoCKez33YAo
9q6uCWxjYuTYEKyuLYMlhWmez/2DsSh5P0DCNdGDofoqZZLmY5FMgkWKfWE55zci
XHjIF6WKngtzWO1VzOgb8/INRENbSug6az0Ce3AVWyz2GL+s/e2+jMhrMBDPDM5y
CI0jOaULcxVBxooK/k80s/hml/5GoFDddH7GZMu94I4c1rNYMxM9OJolNelq8AzY
UJAXeG2qGxouFByarSqO7qlaNBxzxMFGy0hnzn05ROws6o4aFqesSLpaiYRPEqV7
dGrKHwG9JSnr/6B5vzY9yiQBN6ZHjRcj1ZxOkkAexiN7vETv7IO4KXo4CRXtGUo8
Nnwa6SkI2RkoQ54JX0S58iNkGM+/9lFqD7izhO2EWRT0QR9M/gqoe9Lw62jBl0bM
yvK6QXMZO5o7Cv1BzFnbhecxp8iTiZsa7GrH5pjH17veAlhTDR2qwOKVj2QN4Id/
UrE5l4IHynf0cPo0WBKpkcJ+493plgV/K4BwWGXiCRLMqQIsy3oekja/p/2tZn5V
Py3/9Vr0VW3IDmmooUgwG70lhuWtlLRV6kg0Y5CY2odU2RXYuX9qZNMcybgk3gIE
X5NT5SmTZ6mZpqL1YBPW7O+8sDuZvKImf3H+URlVnFxwXtKjbcXAbVkrqJq5TVd2
e7WPHrsAhlwjytOSepl2OYt8X7cBbDSeZXq8mbBcvEKEK1vslP7zysi+N1mud/dA
GHD7diW2znHYVpm0UF6HCWQoEGD9BMqIMPD9U98hBk7t6cqi1WiV9zJGccqdx8kB
O4+WSL1h5IleB6qXjSzxY8fWev+pByK7BJECVW+Jfu4oolZr6Yy0vq5t/OeOsqVr
vMboJzddTZlkEpDRfV3bMaTj6A9R1HIojeavEdXA5QXLzQHZ60qjq9lIykgnbYVo
HOm6wSdTd4688iptQlYbODEBvgmTxPutO7OJUboNOKrz4VuuuNp4jxJLJsCccTjj
wbXlc+uCN4W21bLWiJ5zxoMVLTW5g2JEIbNc4eOeR0/DoNpxElkrY4hiPDMXqFYW
rbQ65BwCh8wW4QzbsIoHQ0xhvbvUyvWH6eQSFlLfEBLTbMrttQPfx7LwEwm514uQ
90Psh9OGb+u7kEtZ1Y5N+9F4Yow014H5ubeMhrQ4mNhH98+iPDkK3cMtNUa3wMxP
zNGTxZUku2gp3mWZ0O54i/lsXvR/C1OsiImEFPgVA8eSeoZhcLkaR4JAFx0najoS
pWUK5soz+xVLgmAUtKXYbvKmWVVn96DPgfLRdvd6ghutBpriUYoPaIIH8XE7o2wx
BIth9Pmb/V2L383MdlGI97gBPIOpxcthR0Ha3kMO8XHZntrOaRYhml6/BYXZIqNz
xTMNhPwManaBLde7EJcuhwdLnJxRQhRE1VF7F5UqOGwmqsg8x+SY3esYohwHcabN
2f3S5zuyP9oTUaeeVHPWM/+Y6tolYHiifmh0I0WE+4hDdkkS0YRg1XoWibFXYZBC
PHLGPeTl4ElVZTqWN39icpp2/5JRwOm9AlU5cDm9ORBaFRG6fRH6AAuwXrjeTgDh
NAFHD+uZbNFxbpTaIfkT3KiwAqL+gHsniZKLaRND1IDx8AAxlpGTOrG2w7w9bePL
jTS41BO6T3O+lUHK8vgwcW9JQoUG4TyecV7RxmWylaMDMIwnYbPfM/FJ89P6Gdcv
28m+kvKB9gv+iI9ud6gmkPFgJdA4k/2T+/JFQhs/jAuC+Ga6oB04xs6NOdWl5/13
mjhX2b+ry9fRp7jDqGHP+AxfcJU6SYFvpuOGfsd6ZFq4vWTyUElzZISOuHl9KHd0
xZQsGpK4DtkHzoANKJJnI+n+8YoYDr3siFBK8jnR/8W6y8+3T05hT4wnD890wv3s
X9B/2EBP/CEfixO2d2B481YyEGncrEXitQpmqbGsufSTGFiYx4FQRWRwQt9iOmOo
R81TtcDW5itdnDPvbG6ySe00SaFa+HQTHGbhA2WdSA50vIm1Hx9Yf0Y15fDQLNOK
1JwZ8UWnQRMWc4wAEWrN38rzcopu+y8wuUsFmmWDUayVQpGhVX7/JNT93ibjsmE6
NwKL7TR82BaK2fhq2PT4Wq25RAAougIk+h0LUoD5jZDbWj5VKUbNdazzg2YVWoEj
E38jqQARWKatgB4f19ZJ6UI8aUfcyk77dYViwwjQNssoKJ9FWJQvWw/GqR/Si90C
WC/3HUZKh5ioInko7Tp6nImnotKPFMOCHAtqUK9Or1X88sfer6Yx7XqnpCy+Abvs
3I7m5lncLPD2kfdkKK6HuegmmtS2/J6/VaNB7dmzSDX490GcVS0DnqlgviZhoRH+
Ddms+iYp+Z0mhypbUgVzsQzlaoKIRAPddes0s99pdhK8YColxbTwu3T3tEkbW9yj
bk19K8QAC7dqkQy9U4KF7WLWIQGge5pydTb/XugH66QrLnCNTALNuWPvUMzxu0DL
OYqq0/HATos6XBQ0pp1VZEfjzGcmgNyXQ1HM8D8XFUvX7MJFun9XvsilpI2cROD5
gizUvnkGpocououPv1hM8BaLs+myOU749UbkDljawFS/X4MnXmFMkH+7sTr0Vq7S
DulTFEFQIey+CfCTyB6+881SoZjC8U7USaSF/HWSetQZKESBpdbis5VceCgTG/lU
gXyptzBGjoBHVUEqb8V9IuzAAP+ioBEph9Srtbjwrl2rkHm+KrWXNxMz/uIeitsu
mHd1rnXGAA0rmSpGeUMc7RIEdBp89feVAwcKgGsSS6Lf1rProBC5gTbB3/RlMQ6x
pPwsBEFRfW6eWoP53+EvawfOnnk5/FQf81mPcM/wE6KS38y+Z+dOc6PY1+V81apA
0wVA6WSDqY58kgHzz1YhzwSGg+qYfHWTx+Oze6QqCoxRIOj4jEB2Q1up+VVaIor3
7eObDnXHNtAHCThLu8u3t+15DeeKhK2QHI43OrXWJqABgWFiwvQJ5qlVRLzFR1Uh
6tpdv6l1uqerH/X+8Z/zdmWuPRXhzc+Kni1DhbbbuOTvcYXslc674/D6T5t1YBxc
T17cay201BqD9D3eK1g2WzEFaNTNqHsX0RN/0WrmgK4OBPXw+++0VQ1oU2ElWtQ6
5njZDQjaOVO0VCpWXfOQUR7Oua4COR4QxKskFD+F5btfF2hVCJquDalQTVM24jg4
O+PxI4AXuywyhNeaQewFJzq7yTaKWz7cn23WWLXNh46hvN6/WPfVNmbh6IrrpvyD
Vo27kHF5z2vNUfjWC1LWvRzS8s8u3XRThGnEEyS7OHVF033igBiRz2cUTwdRjLXW
PZ4UCg7/EX4S60JGKNRDj1GSPqtZprDsx8PIEdRdghLN3LLiaKCzIVlxQ2mQute7
hzukqeqQMDIeFKdDOReCFdmgFKUOLoLgCdKSaS+ndW46FRFvxkXZ+Y0AXuPUBVaV
PAVyRODhINnwI43bhkun9mGv07DFQZJ9NEly4w7ApWUDmRHtbk11phQppfWXGG3Q
P/MExcOvmKffZpGVaxAIZdYKnLWzjYUkJb+zG0+p+kAoJOHadvcFuzluAFXFg5b8
nbH8e+uE/dr+wrPaTWQm073PZToR7XgSSCxuNFN9cr+5MF+FwRCvvCVCIn+0zcBM
onloqc6jfZW3KTCeZQx4ReYkfNOcry9Ay6jQ8VGJIJvUINkbkf2df0gVoxqxxCJo
qrTOVioV3ZGIwlt/Zfi133vpyGQIO3qJ+kAwJUFpvypRqd+qRQn+JFFs/jDY5nOo
aK4UA6dGrowA6fDVPLXue9mmGh6FGLj4/zIK0RC2WH+/cEqz9dKWoFr9MFQpP/0w
ZQPGNx+PaQNX7+a0DwGmlA95PY/WyHpTBou2lpRpgsJr9E+z54zDH+BSClBLHtpE
rkGc56j9zSRrQ8NHLETPEFtHVWrn1pVm/2V5wBLgfDY7cyU8UpkkPsi2voirrWzs
EiiQnThhXAUcTwjMpZHZEbaXpCvwdcLaRg/uBJNk1KBIrRnXkrR2IsxOwEtpWSBy
bpVwY4dMCJdzWbcSrekBjMf8oIYQlUxdD5pdkQHrcG0cxJSEBdLbf/hV6BmpgQbh
OC6Ta2ydazFYa6uUF4aYjvv5n3IUrCymRWxDZanXv9u+5kG6Q6lCi03ZMp5VAyu6
wMu/xDb9e6xHHWp97zkoQnig/yBxdjO0pB5/r6hHYMYbzZzyjz/EMxqNJoaTsMZ5
AQOEH+M1yuahtVrqt9YBiXDM0aHwJcdbSYigQXgZFCDWxfkKLViZOqYgk6YRNWJM
uUXpUJsrbBBKc9rnk+ohWbyp/zAqP4zKGxdZvZ6R3aIWA3hvZINng/f3CePGbwhN
h6Ft4yJc/qw8XmXw5QJ/WUa5Q6zGPxngU96/AxmmcmHp8VnaGvmwFlVa0zU+4Mzf
7ki9taXHmVFYVysHebYAsflGrIrpUqGfbM+ZNPfKKP6/PaQ/P2MViXrXxF2xqO/W
VfuGUPfBvwcJNalDxYqQJnNqunYmRVUJQSC7K70tIKWwPBRp3mX7tJGNOBqOI9Cb
5rjGHstfb0rZs2IjoiZhvWzuubehB+MVX0QtDJJ01sJP/78is/yCyAgol106jZqE
dtjwGOnyt0HWvbqCXPPCKtHhY3uIST/LVbsD1W4zErE+0GASc+OyiaBaCstwK3Oz
DwxPXtrhVwU1h3V4vEBegASGmhHhmVKdgVi35dCBIjw3Nd2vgRqjhn9ZPLERsZqy
jVDZ6UXDwIBKpr7FlrPWaHiS4rmOJQzBOfAXj+E83Tm/EC2mGtnDW1nlsoIFQraT
xBhZbt87ETSEMsLvA/jRz0HLDVOW/WUOVEbRWb3vKEglWxeDGMiKCgqn/sTTRrPK
+lySMplP5p0bcpqH0U20CsxF01+7XMIPkhQ/sXL8eQZHQXJSepfPiFR1QdKmqSvf
15ovJJnUWrXxb4R+tHFlS1Le8Xd7raybc0dkeRMwk9AD9ZNcU9B3Xr5cWWFOyv0D
fnlPbl5FKRpXyQEx+352iVw4MiKJFi65RYCe47iEvPufmdCjdxvCv/gHvkjsp7X8
ONZBKsdofqMMui+bbR4qiOltbokwsSNe2h1vUsM6Wc+4yKcgFaQ1Jk76QOKnZACZ
ccoBSuqD+xOircoQNGMZGqZbUgGFuughtjyvP+gEwK7oSqu5+H5wv9fDT/sKmC+8
RIcLyDfy1+vBxE+eKhTqprXhMi6sHhSVr2cC3l96T4kttrvE6vCAF0KOwzk1mZZk
VBNrSCu9uq3S7/orcPP7KCVejOxnYpqYnyACu1K6RF5bAC60zYGYilHHGMUdasFB
r7ek5tTphQcF+Xn6ERhUsSEsJ4YOujkcq/Zu63muKuRLOFceAzrJNB+uLOzZfzzM
W4zufXKemhOIwvnWFc2/73BRWzdp1yLYb2L1dpFasnG8/aphFBdtlMzew8qn2x1I
p+NPpMHmOvVJb5XrZtsoWKr1r9h2twjXevpvVUxiXp7bt7Y5T6WdHTWcqHrg+zxu
C/fbIe8EfgQaUF4Z56iFmvIzi8d7yiQlebCb5b9emKV586G+apxacdvQgRtVwtCY
vABVsaogL8hGvK56NjhBJ5EgLz3jAmZdY/i8csEmLGjlClcBzqGRmk1T0axasE1J
nIjwORp+imFz6xNbj/Do/OVJgb8AhtNxwXFEVrtWo15aLZWzzdlWOymDfdbuHCbp
cQ79WT6TaPMFpL5UmDzsbOXk68KTMHt2Px6TtIlE2QF8wQrV/15YoOmKHzWi8QZC
otvGJNeQIZoX2GFQrP41AtjCN6QF9MDv7hgdnjf59nQyWHvqLamPI6YrSYgSyQ5c
uNdqYkWlBsnwNOEqmMjlXwG15t/d33doHaJVaVyh6EcuHOPgal7ReCYbDwxke0sa
35gLL6zls5AbY3qZx2FAuWar/ND+k+nv4GpyLXbmkdYi6CF6p8ugZNtKKEVhSOuo
kQs8rBTn9zC7TM/djTI3zHo08gHrFDxeSmHCfu2Bsu/ikvqAwqYZOEFLIlvVWg+h
47uh8JFnIt58lCTEQE7cGoPi2c5xmMxc0GNGPLhi6a6V/OapfAiYMV4/c9u9cM40
luIDnF5ZdPWt6jRjbSW5qwekJsYKEBBMP4NJooaGwieTLODsZaGPabvQpP2fYeDo
LoKnWrYPzP6iWph4Eaeg+/X5tCatlMaifu/PeYxlSBXR8iCszOX7YfPjcaB4q7zx
8V33UnlZ1SERg1+voOMWgIsmBJtiy+TVm6JSVWEUefJqrk38oPMyUiR2WX6hQhYm
JfZLJAQMAuDAMeY2X9o/+QzC3lqzWnOQlOxix86Ytk2G/3N3nOOTKQnVh3E5ZU4a
0L06Kqy0D4fQ+OuIKyF8DpPyw389Po49vCyvuVjPNn5HXef2TVuc0O0cdlg2/zaC
kAJdqgeasVL1eafNhkxFsNH+NQaHM8SaW9xoVFPHJzBGi6yowy3clymoElKcCYAW
2zxaht9dNkX0Y5nnslGi2qmCvrZGD92+cmywJZ6xbbI4ewGpYqaOqw59UFKQz257
nu60X1hB2Qq4lUqAEmOFUZ259mlH2xI6d+PfevX1Rf62HhqufQne1UHdyywo9Nau
o1z/22bRHMz+J+PLiiJ1fT9luclPq0LgXwExhgXhw/bm9T7x4iaAMYGneQnGOep6
f8vxTG0XW1Q1mnqR1QY4M4GWdB7q3X8MQH0JcUcG+T1STd5G5BVU0J2J/4b6j8fR
3lDvT0spPDmD7vElFJHGKH/S97T0w8nMimXQt+Ck5a7Y8GjGOh53SpEXl7p7/6qc
i1Bogn5zUh3XNZ7g5FimYefYbFX6iGWyjiXGT1hv11AeDfJVuW/3UUpRAm75P/XF
ijfjAl6Ot9f7RkJ8e2hGsWlPpQz7sqI5zQf06zRdULpOBLFLtO204sPA8xz+eWM0
yGZnX4rH0wOPROpaJS//T4VwkelUU5SljfZsWZ7ZpYGVXExAifx7KoEJNrRl8wCA
FFXmn89aHFGiWgEc2eFfHDX7hBzyYyKIDMMZbhJdsRVe3shNzvP9RwXPt1KzNEuu
vXiP8DJu3XpIqUtF5HbXwmPRvOcLxWdeWwVrmdPXjC8yb8kYC4oBSW565ao4B6wC
jH+huIzPt22fzBzz7/wlPt/gqkG+ZX6VDW/7EReUYJbmbq4yKqeoADeSMT+hURMQ
K9p7VB2Qrd3b9qFE79xwQWNW7dv4uvrGE+wpiBZ94u0ybrryVzr8vK2551hI/Vj/
LVRBurQmgFdGnrYjaAs1hlKwa6vW/VPbjh0rhje9h8tFpEGCQDqKOAuc0IPORUrJ
+0h1nJlPIh1YjrYKttf5CVy7rjyKL34276t85ROeNq7s8CPXfJWBYSWc8OotgGvo
YsXT2tDMgUPJ2v5Ogqm4E+y0LTWUUZ6v7UAXewUYLlrWot7h7hjRbuY0vBd0q6D5
Ofo5hH/fkIaXcKPaQcOpWi2puRL6nyPl4YgqOSDbGsZ9px+JUFFtr+6Sq2MPnYEn
C4yvj1R/P34bdFUStlhHMZVGoJE7Av9c8waH/BtCneDhIFRPxrCwxOVZj5CN84CD
FBt3EWFQwA6Y7q2b1BSqDYZTjw7UrWbe6qubn6G43UiWkzsAtelHyR0YYmlxgrLo
wxbIIUwqHHjCuBmbrLcRwZnZe3oTqYJkzvAHOO8mHSXOw1MTn5v7ev0xUn5GumvG
TMf/pilR9IaW03ap50rfzBOQHHU6f7xdzveX6yxcHiRxdv8AQpzR61bp1txtyrV2
qCjTUDlPGinULxLIpyT2HexSwxVJIgVZl5ojKtrhqChtX7qyv+SqT0y6TqcHC98C
kmlr7y7s3NGN3th9dLvEyOyrAABFecP4Eyz/Q5Xop8hNwbWPDqz1Rw/m/K/EuiQl
V8ghvdLSPkGVYu4TUPM3CMM2gLpESJQDUpB78S1WxdYJMXqkTSPk7weyHK3BQAuh
TVDKDw7VpmVMo0IC5ugkPnSdOPniPXKNEoXR620MkGCcdpVV1vgpiYJLwhwCW4mc
rridBKCnArlihrhChgIA83MrO/uTThmFhOILSque1bhaHgOqesKCrnaWpRme8MIw
AKrJ1v1M/syaFSMkYJ9io25c2KS7Zl8wmOFRbBYxquQA63u0C9+FvDUzOJBJ6WIL
uL8C0TZUn1BW3M2zVPd+yi5wQcYbGTn3CrphmmVTLxFs1uhOhsHz0i9KCO3bc5cn
R4RLPikXorCC4iTE/06u1c92RB32X/o3AvHdAjgBfzfDbqUkRvmZWBwX9kAs4/5N
k+pm7iUaqyaUCeUbUXfjgq/zFp0pIWRCcVFy65wykcL8TqnPPjBnaG+T/53F3w2o
875ym7nXCg4Z6cxjKZM/SEdZK5MTTKmAWbqHGSfo+aN1HzTSyEjaVBampPri5T1K
yN3vM7upb8n4xKOp1ROgYMZhbfDyIDG4dCI0otdkb9Wu7gK7TJRNqiLkaE1tEt+V
GgMx/SsP98hf0OURYrPoS7gtdrJuLhRjCVVNWi9wRLBXTsddemSkbLtyFJ1mJNFc
2JgWXAZHkNn3BEzZzryWq7shau0Qj5PYYA+vr6JxNF987T1bZiPSq5mtpz2aJHDP
3QngjS97oWUGkUUqGARVJOhlSbP7H98xbmv3BkxUf6zjm+0+pYZWn6h88VsqDmfz
2zIxvMT7696PrNBBdaTEFlxgsG9Q46bBD6MZDcWuHLdlPPyWrdfupXZqIKpVxR8r
aQhm3h8hsTWDYd+a0NI1s5uvP/XIZUY1xg2lvzIMyJao0hJsDBZRYYuoN547z3w+
QdmLLyAXlLEQK4X3Dv4arYT2lcX5ZjTuwhiAFNbHPcNrM9lb87d7ij4TWj3p2YXG
etREN4fEDxnyxGBThzFu1vVmpB4tCXvwSLOQv4O5zu6iEC4w3duB+LKvyLSoRxGR
JqJE/nhXYObrK3iNUiep8k34xURalJM1ufyeJBYY2cIVKZ1USl9jfKZKTp6pIYVK
SxnOV48ske8LKzSt3W1+fymSUx8wXvBRdywnlK1EnnF8ZnGfRz9m4oaAeg7MH46/
bfTZ4AkHP44Bxka/SCv0i/Kzq1c886bpU32ImETFPOSJGWIFvN3B8CQDzSyDjTR6
EQrswW+/+dcIM27/brGfBAS1r9yGuCN6RdYDkq6qUNdIy/jmr5ltd3NOb75EFN06
gtV1AO8im6wAUgpdBJyclprki7MdnRg3zZyhDj5Yd5Hopjp40OYRURTf+doU5QzJ
rwcvErxThLFwRL00ySvN0yh0FxozVrrUtsYiqyoVoWoH7DTuMz77A4oehjiVCUgR
iDk4yUMWmLpvVxtMIxfTPT/3v6Y2I66e1km3Tttfi/tQWbgsMNgq2CdJpptSejEW
FbxD3anhptOrLMdWQit1egYDKS0PzK9LeS2+nzBEmocAe8mVUPluvjw8ajJoBBmE
ziWGFNXM43cXjmNU787Y6cbApGIeYKNQAMR5IRuNOz9K122retJN11ciw+fjdQ/U
m0ONnUL4j7eXO0jfkgoaDXXrzwJVrCzTLeRpMaTXAFBRTfe49xueL3cTyqyq7fKK
GLH9kf19huVS61TU1mCEgfUZjR+BwBTb0RTGkm52dpglGoCUPi5gXtWJIwl7Dzj/
uws+krMKWEw3wDnEq9TAxzrpu2fGR908VWxqI8Xi/tHeaxBewjbugKh9Mjf0/tf8
acrPtcbCYk0eu8Z38p43IgdM8dF/rhvyRPvkUOtTkTc3Mn4BGGQpIuOXux0f5dda
LUZ2QUD9qhxZzYr+FS5Z/mAuIlvYJFSI/I0lRvHJaAM+G6SqBKtwc07+8TYMRmcw
C5JBG55SdMjLQGjdKxl8fWKJ54GELQPM7YHjOHQ/q9d2fFIVHWjMn6YLzhys36iC
9QFTuCMUreC2g2swqhycK+0QEzdfUU0B5WTdXTp0EuKWOjrx7lPyyRJL4gwesryt
k18Xc1U4S+dsgrU0SCSOIaQBcgQVs20oX94qnhETn8qGzATydzpDP18NDuhW8rKm
MnSrPdSyM74p5MlKL+863awk6raJ4T8kAjpO18OYJx4pQvp+rvLlfjQamGZNFuuK
btvZO2LlhN1CBTzl2YSt77Z1JQntiqZpBtX22Cat5wP9rW7WMrnS4X2kWBjlMa2z
UnAle0jG5mp215kjs4/asU9gn8Xd/VmPPBbA9Umnhdhwfib8gTtQSv43QUdcUzUD
zpF6fF3e112RZa8YexJPBa+z5XvXgWblEaRCqUuVarHp5kTTUK3cnsvoYWXaH0Tv
UcIbS0VdApviGKgQo0TL6O7Jc+KaFIbjKksXm2hE62mnI/X8p42eu6/o7/BLMRSc
c5L9X/mxKnY6VPONi624rl9KsN5yNEOP9OwqPEoHDLGG9G/7maR4pPAKjAE9Xz5d
NnjRd6d2mcP6U4uQHq73UhQ0q9TtY15mHQHHkDMXCHWP+VCqti1RXd/iBIEOq/G9
o+zTYbkgbilGAkckrHgAAITv3B9IkTnasn+ruQTKxjFNZwyiQtXVBAqbR178M328
asH4IWsKuhZnYyVk6o0sqe4Tnmmj0qn9xJxYEt1xYrTTFNDlQO8KohOZRSwUDaIT
VgnZz2Us7rT3Nr1NFcbtf2xkCQDfS4LKD/hPKRwoi/H/5xvXMOkyjVYNITPCqyeG
ao0FyQhE4RvCTU1Yo4QZdJkvNPDckfYLvcOg47QQHIycG2Q9lcWc0sN7lRdAca/i
RUwaW3301SXbyv0cQ4yV/brjP3H2jsSt7FgZFdNC4KDv+PFWVXik6SvdkAgpS8hT
vZvegKAnJhXBuJp9aIQhZ7tz09CLWn8200i5yCCb2AEfl+noQq6OlxIK0jvbC0jL
KtDdBcUolW1EgmgbEHZHblJ5k17MRMNHbrAReALByq6wjmO1qmJ5s9K2wxtFqe2x
xYE4fwTGK/Eo+S9s0tEmtUdE94q+FYB2uoW+39i7vISLA49iCFm+i9uZVgoUodhG
JJkUD4avjI5/FI6S6FTqlQ84I9uV11oVf5YZiv0XZAdKkBsaw32jdL5HOAA6uBDb
+9F8Xz5OTrng2dwp11qpwWUMm0mk519tMlxDQ8j5FBFDOymbyZ0kJqsPSTCDZMRq
QiCuBs8XZdqLqKrc6D2c8fwPeejWB9L1Sx6RjZHV4jzxsmmx7lKaROBaQw4DyB9O
UBt84Ie+jZ+msv2f1JcuiLzlTtLi06KfMoI4SKIwZSt3Xg83PH2sCk2wwZ33T0ut
3Ig9qERFHXRU0chvJNeJj+3QVfmN0i05mkyPlZ9T6ieXLm4s/QIh9yGSUhFMp9R+
gW3Q9M72xuQDMI6q4a0GCY86XNINctiTj5EwI28Brh6orJEKNNVR+EMZsZ86736E
pUsR0QFdwFBVoVKV1QEAXAbfDhr8p91v6jBNkRyzcWj7sEiJZWn6B53VVBgOIaox
AhosU9PA3hA6+ftchyHNCkWMkOR1NWvIHJAtwiMmrvoQxKAsGlNn/Qh0u4qZNef5
QcgndOEkz1Ntc8av+luHLCFvmPXBpXKTFahbV5O7noCLOgb0rL1pEk8ZVFzpj8gQ
K7FnXATRirAtUlZnegwteo/fLjVWxmsV+Rfi5nivZNuyUCIfE6GeR9FaQG/4UpaO
Uwc7jrEcgW2phJA9PqcZ0HkUtB3LL4Gn1v3y8Uc1PoTWoHYEbXbnGctsvlOd36W4
P8sFd3FwNr473W/ESx5NdTTBX3FfNAWxO517E+TjGAeDJwyf01huYPO9ieAYK7td
b8zmQel12uCSKRLA2zIUwpGZyVN49TYkMeVVB19JdeTwqoRgWYCWTor7Qucv3WRU
25FNLMGlCW+x+AmcRjt5zdK36O36MDUmXNrfyrSi5mBMm1dt0T8yXB3X+jU4DB5D
2rqmhon6O/3O/ANy4mkl3JFK6Q23KCRkhgTcLAb4hS14FcMM6hy/Ng2jRfspHcXv
znq7HcDhY1f+LK+uy26EvvGXQM2Uzp0BQIf3GWR4svSCncVu6AHN9CXFvfg7KMZr
3H39q/Fo+zanez/DfLtDospek8xUeLfMblbO3oare4irBynDdzCvzoAlmAlgIbsU
seijswp67ZznlsjnuV1de+nw3k6F5mMj6gWxf55QmyR99/RG7S6mBu31X4CyFL2H
fcaL65PO3tYP0LdFgCqfC6tfPElh/qtP35vCv7w7kLVtJTAb82SZXLMX2EZ9BeHH
gGGsEv/TxLc2VC48zlM0QYZKp7hZrJ/5/6t+gdCyhGVIZ7swwUboMnF6RH3xOv7W
i2XhS47uUU5bvoNG0PGQ8YLyltYTUilGcVaclnRelCJu8eE6PGYBpiQ2GFJws1dZ
sehnZLL31u6Q43AzX8vWCNqzT3p2x6Rn4q5oIDQaDsScvb3A5xfKTJ9Z89ef76Ed
26dDp+yZ58wlCriweqnfIimh3L2jz9BLq8Fx67469VANJ2ASwjgjgE8XZXVrDAue
nfIKCNnngnj0ahnpCh3dLbpkw88EhMYQDukttzBcVZKYVLL8wqT4D8bR/G38iReP
ECDFjgjfUySQDjI/cj5U2i8vxsl3irHbXToTZ9b8fLuI8+GXv9hVg45nh0hnQeVR
1UVS9sGNtuUGKu7/QrrBWtIvX0cs1N75vMdgDN63TPanEC3FC/LzY2M9i3lh/DUx
jT72czjeAP0r9GtHhbFRPzaKNd+PVz3lPMMT7uWUX/IOnHZtpsSqs+3MU5pHBOzH
3M7nyOwaWQIZRn1E21Z/Lkx6TT/tRqFm7/oUMTnOCLccHbW6l7Jz0Nxs1VWSs88I
w7ixrnfbcv5Thp2epwJXfTw2E2GHFOuftHmTBAMGfDZPqDXpOdK5rTrW4MT4u/RN
BjTA5GzINmvPwit2b2oPiC8n0IkEwN0Z2XYT3sGyYL/p80xta+wqoYpcLpS2n+fD
xFKAdMC6Hf20FgjSFnqJKXJRnhdsvSjiIj8812E264gyIJvY5Bwun7b8oEDk+5+f
jZdPJrh0IvjtIWVXZ1fcqbhzND3psKHYPMwesffv/OGh2AX2hnUEyCFPW1hLboOB
BMbEjCaHA2qTvUFgyiB8YpvmIcOHcywRT6SvzJAGyoJ8UC7pvfenPsRz5tRZtscJ
2TbWol1Kq+vHek7ws56wWmqOqI3VeleIGipTGz9cWhr/rhj+APvWl4iC3G44uy91
LIqmzrLMxo1UhaDCZOz1al0T8vRpZmZ7RURKvS4LXZLTPybqmpCZt+kDIOXxXphl
5W+xTxb9sB7SWO0iF7u/WUKaxrsu6tfeIPScZp+qbbT2JvmM18YJQHSHkUf0oPfl
pJTP2xIjYc5J6R8ToDjRkOzwES1C0kYlw4E4n5uPqLVDmxYhV69PcZxZBgqrmH2v
XFWAozn7XW5qYH4g8UUF7I6VUWVl2MtE1dTw7kMg0xKgnJDkhqwgZGTEbZI9pTXJ
cn8BYJoB4TgMuWPCJiH8VbPRGI2DoIkpaxCHcHmOzYQHdRhTMgrJaXrZHvALAx24
ntYgFLul2HeP7f4oTmkSAew5safLdVtxZE5dYaQ4AXNF5x7DYWxvELhublHfIpOH
YN024Gnh2C3r+F7hh0SMFY+dNKu4CvXSv1l06FyunzDcHlLnXmr577B+R8MLaRmf
vYnUJoRJrHmTqnT3M0f94qSfnQW4rnuVbV01BI8aNDPfVF8mdvOGeJaaizRBkKZb
MefQ/RoVnQDw7q+TOFqnsJ3KGIBP+V2GOUT7oDm3m/eVbFpZDH5Ehsq3sn7yEOYn
hBqINbIP2kFuNHFl9b0oYIF+L2tLGddNuWBX4Af5GbaYhj47cYwfQx+vBtREQb34
2tyveqeFKa740wOxIYO08ZM78NQ6FqtmCNqyN5O0wvY+ry/Sh4xeCwEF4vdwBM3Z
en7tEI5rzUEZL9QDAwCZwBuuGFMKXii6570RT/cx9FcIEOYT/yM8MJX1hhUO0+mR
4/LggxalX/Wo8aM7KPpqm6tSGJgo4mFYAGXoAwwJntLT3vvV5v1C7wXQyTrMYLmy
Mjyp602WAa6W5CZofEvp/0MSLd8oiHqJsL+lXFfnzFHMg9mIJMQGPOyze4AzgJXr
ZfvSSL9oypm0uIb/4wX25pj5u2hs2MYSO1Adkn2drwvk0XH6e5uKmkpjxa+d96ps
j/RdsqzYPSnWw4SzI5coQxmZ6FMdS84Wh7J/wjHmLledhzO9QeQ2tDi6mIAIg4Fx
843NvsqX7CP7OX3eaBJh9zBs0vOHJkXKbcrSna5pih7fzfGMgDzCEJsdCJWlY6rX
hO+oJrT1hi3oT8/14KapZ/2KSMQDEqwt9ip4iUUsE0VUZXWD5iyv13/ORPmBnL36
w4NZmzEgz8FMWZsQKPGgd9ZPx9GD1947gSH4NqWTbXUbc8XG4AialLD7/c174u6T
Himox3VcnpwQ2svG7UloZ7s+ELh8gQl1TykKg1wg5MpoU+7a0zxzyYqZ8t7OkSSS
1o0yd//KBBSii0FOsxVSDQmN/zoIw3lANTmKs71o4CEYG7whXNo3XbA0WG2i1TmN
kU4iWnUqv/cm09nr82YqA5xo6m1neu5fpMxriReEYmmCsWuZCSORU1DyUsEydmTp
BgrQMgnbAv2HgqFX3pb4q1Tzq4JgREgy9BQHZIuLncWmc8Hsed7NOSpE0QVOIVdr
ieJuywO3itlmZ7VwuJVuiIKRJqlcBaqz/wU/YyL2RVIGZ9Sp8+XI56QrPfpY0ayU
aSX8qGoliNc5XPBSjlwcwYWI2RnIckTwKuQjl8dodfkfpjXbmkblyxbfjl2wZrY9
35YU7G3Bou0dNTiFpC66Oo9H6JTnu7B1NyCksTmY3Pz21iNvwlkFagSGCQYgViwI
ahAfE2GZAjoztpqutZv3iEmFvyfp6a9CEcI6g5CktjY8x/FyPq2aMJ0mHgbeURap
g8MiaclXgLVC7T+1drFtq7GrOtwAxHrUvWAEjDBJR4rv7WQ55l7T/INKcRLB+uhI
0K5U79AytglN7nWhNVdWyk6HYgbWUjI2dV+bbo2Al8ZzEAqxGvjrlb+fM4+o+cvI
9OBjIDtb28NnedVDqndTsve2IP1haQUhsEak7+5BLZxBBubgi9z7QANRhG8k0lFO
oZqbC0s1LvPittWNB6IOKjITiKso1AktctxNfKQKPeSqmDiRqEKCUq4ojWgInCMb
q0JELgJeejaTVQPgaQvNcq2gPaogEWCxVXcQ/EGvFQ23CUFqL9JD6aiGTW4imQX7
4MM7YUMs6VUTD4gupekfyak9jLwJsormA13wA88tYlAqGCNtLLipIVRMPqT2ek3A
Vnwf+oezXpv7o46mE0LmbiyzdRHzpwuIAEHbXF6g1NE5+Lk6XF8lOIP50W8aUz3T
BEpmTLdDScpmOEN5ygNh15Moz0xFnOHGr0ogN+mkd2SllLjpWr2pNIZDZQlKPjii
XLQjF1rx6BRWfi2vk6/7UL0CKhHG320aYiMA+u6CZ8t5OnmGTIO4FIWnBJEcPnoH
rOp0WyVtJrj8PQiTQs9x6u86RD67v4P0+WQAxRTq7QnvRzCh9kmWYI85sEllPsKy
9MP3fMyMmkIHk9GHwc7ITIgGUH3yzv/CQfzK5hUjefZiozo92PbD5SwmSetrAzGH
YIpzHVKoigqRe7hNTAT740zdu+epKOOihJXvM7tdYNwQNa5ABV43HcQzJn0nS8vj
LIEsIu8/xroRDcH8GsIQU+REudkzT0FRsSPvV6OAy4rVgEkd6/aeMkhJ6hSqSaG3
VRdSW+55Cacv9YVRUhmWrycsv+Hb/r7Ht2e/R0XEfqCsi/l8woRqbT0uSZyhJ+Py
uDuoqJtJ5LfKmwacBwODEhpix6VUwFGIemeHkwSIgK1JK3GkEm5Aiancnn0GHRvk
7cOCb678qlinsFYOvXD4zpm6KKlFfZtNX5F8IAq70Gtl/karmTFfWQlWyJEP/vTr
4Enp67MlceJVcgywadalZ/vy3nvO6poaiW6m7zEHBs1Z/2HKxSgzDCjzRPAZyiDc
IAtF98U0yNSmP9sA8+czdPsIDs0tRefUyo9b85bkNi4eLV+uYog7DSSZsYnmA99U
o2Wwm2fjwoX282s7BfmJz6V9jSjTZsGhfHYRplG4notfr9huagSAVqXNf4Kruz84
SJuGTMYUXo/HPbh6EsbQ74H1YOzuscXOUdI2RE7cBnN3IcS5nXiA1i1r1ndiJ0dJ
ZYhV8q70dawnv2X09Lw2BJu0QOeYWgUGYtLAMs7xAYxMdQSdqKAfEY9HhKRJiWFk
5YyBgB9oZJnCVnj5oThhnA/6hysltZnO5mj7ulnab+K0TlJldfMxkhQTpEc+g7pU
yfqnEEeO4ggrYKfYctOSdgtQ+HpAitFKJP7yol4GSZ3uNTNFeStkdBIzKvw3fhQA
DCeWlD89LDHJec2jo/V7SLR7N2NNBvb59mkjCRbbxw6Me4sW0TPFOiI8+QAjhKKA
dHcR91nxmoSlg0jlLKPdMZcMOk+anyH4Q0vl98wEk9QU5jTgUmACsdN5K2Ti9S+R
rk0MUc5bC7rwJRby5OdqcuL/I2mjh3b7+WtmH823NNqTyNGaBkQEVk4TRCtpevk7
Ic2iQIc07/nIivTSoxy2eflPNf8h3HMY1CcdwH9f1M9YfVJshPW+QK2bI6xmBjxm
yF+PhKIqQkmU1A76zVO08+rgM+lJVwGM6ScAa1wUqAr8oHwI9DBA6LqmYegkUCju
4xbeluqYtjtG3xplVKzZoMhW5tho3bSd7pJtMUW4NVPR0Fh4FDirjkXO7aqKIswj
Zz6IaPT3pAL8UBCE2kJDK55j52uzV2Iv/R1WM8Chrdab7lMTfTVuOSJOH/dr5q/v
LVEmd3+aLgnJQrqqa3m4YA6kTxglmBEplW+qlX7YGPRtANaqFjhrUpVZaZ+nUSzK
VjU8GDSC8SnB300TdEJsE1V17bRMTIUZqWhGPLTeGvNvvv8QYv1cfJZIgfHYTxuj
IiQ+K+URc7cqvVikEv2Vjyb7006zPgw/mMnS7m31dJymbQ39m6dS69C7G1dmB71L
uVAQcvNKM+z/E9+EXXe4FgzHX7wC4elWnw1/gv+ASKsufqrtdPfnVZMf5r2o8M45
0/SN+qCg8qbyWPPSz2jbtvOtm/6G+58pD/ADT2kNaTjx3tbB/SOVWZY/G1uDu0vM
hFc42MtxMFy0dEadHrqCenHUaA0MsuUUhTLOP7sCHM19EH+U05fR4kU9HpFT4Oh1
P2VXKaqVcw8RL7Bv6Vhp5knwF/RwNis1GkqEtsZrLDdcgBLzZrHLUr9RqmZD8TvX
dMrH9UpikSlryDvtiU99O0yEW3i2wQgD8Y3foadBLYsZyJjY+z42cWcjGqWs78ej
rRvx1g3fvEteU1htAEGK8gLYURSJxcZXqNS5CsKCBE7kkwp1CPx/gxMzl+uyck+L
iMGyrbFaKsdvMGsDj9lC5JPgE/RoKZwDp4QmuuNzUIoxt2t7gPqwLT+vmEgJKIIh
Xh2HWM7pzUCqZqkmBl6dlb/u3LgZg8t8M4nY+TbVF5IU+HwznVEaZlrn5eJHT8qP
losXCZFgyhdd4fxVTC69PPzhlAwwXBH5Lh3Me9AaVgEQj/bKS/CiYl8rdzeL4wIa
0V6ue6IZgoE9TE9BUV/d+7Gom06M5PgltDkuEV1p4i+saNubJR489sr+D+LzrkpE
c1P2x0Hzk3Nu/f5Pk00k84e6Ylups3PDkEJUqMLJWJpo7C4oj/TaYFatdhClgJIt
o5Oo2kWvrOMNKwVq+C78ElVNXfjt1AZfZx1EGMwuC5+DlSJnxN8Vcr9iOANhwVm7
xftvLTqtu3FK24280mq9d9kYpVTcD5KliAMePrMABi9PD0X5LAPgD41pszNPDZ4g
V1uPzEchlnnIuktoYsTbDr4UI52186tOrgS7wzhdCFkAxo9A5yHsyeDskLY4mpBU
BmQiboatkVfbHpmDCOZDSg1SnNe4LLMMGCwKVizmCBBU66UAdqJ55+B2yEwmv4s2
hGc29yEq6CI41h2BUEKdD5O3U5bUr0CFlPtlu9rfRlTS7p625F6ACsofk8WLgr34
BxKJfd+u9fUgEzprmxkYB8Pueni5tdz7caB47RKJtmcC5h4fzNYNtBxX23ELiffo
yQpWj/7EPrnIG12bqPSj5naCCg8zHU2Haa/A2W9DvMQq5d8dbPKq/IOw1AYPCvR7
8PZ4vJqLokVYJM6bZD/gM8EB471t32njpD1LeXGe+L2FCqNSWBaXopDbbkrnySJ9
sw/GJQUvGZ4falNRo9cSCzad7yK3AU/0EOkHdkh8xXktOHvL/k0ASXbztwc2m6W6
cdBo5bz9D8kfcFjKnyYhuceOH2oAspOOnYHOxSP63DwJfV6rvTYrAfOT+Wz5AVcv
QpQpTgoE6Nd/Y0ofmy/gCgTK4PNDq0Q5Nppx4T4pX7xmdZEg/gl5PKg5zmE8TDvx
Q6WIJRXHBbXGH8A0b0qo0495URBeT1TMh4eemy8dHUxfwof8TgHEj4sHtDuH4Jnl
rUXc4srGr+vt7RP92lGTaP7fU+HZVcvYJp9fBAUqyPOFC6sEtPCnHloYp8iLAp+8
PETJi+RyPtRudn5hbIbToM1m7oT8FxW1codA43/A0Ydn8gAX5Hov7HyOW/oNKDqo
/fDiwpAC2y0B+UR4wo9B6n5N08FGYo/VpdfwUNsv316wvta5gCPeLFxr4CnWeTHD
XG9LmPYgVMzklX3IFvBuxSSWFWSuNsNNAACZ4ocyQQ/FeEIqwld9/+4vZrykdlUA
Eusw4tkUGtE4S/T+W4JfGte3ex/Yf8B5bQQuDe+66QJ5/bkFmcxjtX8WbEPezlDo
26AX5eJM39OevZbbfo5qsb8UKWHhBhKrmYqUtNwUaPnolETaMVhXHeoERC4kMEHN
aiipBCUZ2U9xO7eiRZKuWdR594/4u/C0OPmtOclviTyIXCO6zJIx1ufsNMHC0x6G
TNBzgszx20xMelwhzk/Z2bTTRM+a4BpfDA/76OGHXQkvdTJk4oitnRvSi9sK8Y96
paq68+Lyrn6zSvd/3wvQvQQJyLIadACfIXlb8OnLjYHRLe0G2o+yk76sizRFu1/U
pS0iAgzuUC1Jc8Dc8lfElH317LGdh6Un5Jl3qnEM7GXrxqWd+yClI4MohkDEUKpU
wrLsS32R4+3qzFOs4qAu8IT9zVB29yObxnWrs6PkI5TdNZlsxNjpUm44GhsUNn7E
7gCUU75EY3E5v1Dc8peu30ZFcS86DNUvMSA62y71yU51C7u5/o05scbKIbjSQaJh
6qYyzh0UqMNp4IJE7hcBKEOGnB9PoShBamX9CFxstI+5O45P9/KXsEpcQ/qROtEZ
nMZxLZP7/9etCLCRiGV+nU4eckbxaJY8J5/p68JILebXwvUFMTyvbq2qUzcW1Ucp
7001SM9NZ7HtrAfuEIeUZtRaK0iStPRpiRb/TAZRukrW40WOslXnzUwIWrGP1GUh
DoLncFmXg8XSoejdnS7cVKllAjFJGoQ+oMa/bnM5olsFwAZFAtzBkARjIAA8U/pU
pB1cYnxPAC+LhqdU5ZMBxATmvQfULopwaV8lWfFan8wYYoR1lCG1ocWJd2zNaU0I
RXIOVk74Xkq7FIE3np+eHLHdvXUr7um5P4vNGOZYNSzzL0zUo53TK390XaoxtN4K
N91THS2vU1JBXBywkeUwNMqfgCKi69hRcmkT4hPi3ya24520UUOYDU4iI+ts91aY
1i9B/9sIWn3etOoS3788fsBP+xSXzk0QsiWJH+5N4eHAJgZrl+93svcCXMlt7d+7
ecuvAvUNFANgKMzJQtLOOjR4nokXLhuXw4B55rOa6pQKhUK9l60msjPg8Ve7pbHP
XbEuz5SakPPkrtyw385RhBE7GhUaEULjz/VIY26wIq1Aq/eUXFhjRnV0WV4/5mDO
POX6FusNPAQwTQvAcX9wQ9gOLfi1H+EfIBCm8TNLPQyyIFuqOL1u5Tt8JvqQYqtc
nZ/RbHaEhXl1NqNyGzjkLEqx+ECFo+lHk7lNxCtuHsNA4o7ojUvfNL/V6P30TS2D
RSS+vkj9pn4zi4nW9bVD5fsuN11ALtvTDmE4cCcL3gQkRJyEpRMyI79cR/SXnadi
9my23lERJSlWYyRUZfZJFLOt2sBwDmAC5zpDYwDzWKw1dgcpekLXf41GnDsJFbDp
uoYER6JzTkMUPtqMqE2rsNuUTim+Y2An7dOmOoTvPVHwsK0S0cu55E2dsWRMq2Vj
TUY/xxfjNOC702kkd3lAiBzLW6hLnBRU6ZmSMOPBYrFYRTMfDbI4hKOxq4NHg2Sc
VOa8MwWyQaZAaspVwW5Dv401p3DRs5hirADQE+ggY9ApTmrEsH87/q4QVxo47anN
HtTJoBlHki1SPrjE35kmTvckzVBLXfyVTrGUWlGNSl9Yv6j1qxVB7FrSzn/vYQ3w
uXD8l5ZMHEx9IO0ntUDfMdu8UD6ZY3UYxq6p7rh92hL08OJUWMAbi34KmaDD77fN
/yz3wyWMo7iPXVUaIbTzzGWAu5bo8WWTd+kxBO6hpst6vuaqgOhwTvdk0/MY3XNC
1Etd/oZIcKtJrqq3DfMfvaZ7SEVNqAy0pLX4g+ZLkShD1C+gCw0cAWxqDqg7hmOl
rpxJcSJGnnA8yDN43fVnwFxXXs8bvLYUmppVngqcKxjrj6sqtAtFkZgcZY07Zx4U
ZxNkBZ8kZnguS09OOXk5WXgp3CZ8IDY2+2dg6J+ACG3j0WSXDQk+9LJgqCrbt0l8
DPALwdj46BMfI4irB/rkVj7eGX4sq4dinzJYPKPPu7iPGkvQnyxtvujmUb1rdXxE
xTBHt8EiXqELQroB2HqBpfM6IcZ/Qp05KqJSbb1h7bNhpU20ZsEsXmj/lji0nOzK
eu8z6fo5DoR6bGZUXpPrZl+jj+jlfIA4k7BghfM+TyA8JCKR1zTeCsZGxWtBsOM9
W7pqsaa0+LUtN+EUPj/YuvQkn19TVc5M68bLECh1oYA4Nr85jf4ck3nF1wwxm6jL
WJhRpqDwJl17AY547DY+azqz2/YIWeewMk7+KUFAzN0Px0NDgfg8BKEf1Ohkmrn+
EESz6DLm47xjUfUXPtX1zqwz92kmxAiKQBG06w8J9LE+KMxnN2lwydIy5ljp9bcP
0WLoA0rNmxgBWqsuo3ulCBcwXOt1kr13upfQFp3KmXMdv6AFX9pu6gQNtB+8lpoB
WWdVwwfrmAO4EaXw59x0KxCUWo9FDUu4c7DPqPeTtJytGaQ0MWx9801mc6T/8UT9
/Ndg2X5PT8yUcftqZJXlEpdybP8wmA+W7osWrWU3xRu7YvZdUui3HwulUNwJXjNf
MVjo+nGhL5A4f/TvcZ5o5Sl1KtG4H/KFCeQK8RqhULB6GGAoo45mGth2ZoCDl+hU
57Ta0q5aX0Cqw5568smr6mkXCMWe0cI4dnlHk2+UY6gxGbz5ZvNu1cFJ0YIBP1NJ
xiexS0YJfjFeixetG42vwHz5BHaHmntUFu7AQIXGuvbenWYMtm+MVb3y0iEoi3fH
TUeLl2y20aGOwFY37Jc+DdnQr11Ki2UKRk+Ag3dyhkTyYhE+AcIddTlrkWVPUG7h
Vq5sdYLDZaBIZMbR1qEi9CWMII4/thMPDjghwC/UTl8pSBuUeuw/cCxFZq8U2B0s
hlQGxMAkgEvyvI4hqf4iDufBEt41mOQTguLhD+eBB0pLqx/mIJFXwsIIbyu0lXPG
dFcGdF/TtJreVJyZmfU2MfTssyje2zGqD5ptmYja1/BQy8obwMZAVYaon+NID1Za
1HFZR979Nn/O2Yp+35wIeJ7xv91spnvmb8XYQxLGCrA+CyXjreLFq7B2fLX8cLkg
IGngnz2jjlhJY9JF8InfuMbQMxsCpNSwIfqjBz1GZ0bQ80oiO4dAA9C7Mp7lTyRu
T3BQjX+sgH/g/Opzdu48wp7UbTY/8TvaytbPsCEcWZcwBdoJQlzgJlEl92y0gNsh
VxwWpR7YzAy41LyzOTjyH15dFevKAlNqgQzLl9GXaZEhqL1JR+xEV68+afqPqIXf
k43qhQ6FQYfp1Hk24xbYYYMzgQQs1Vux88TisqV/5CEzmtRieAZiBOv0SCldGp5N
UDBOcmSODbTavGCuDhVMivmk9uUGylCVCdWMcXRXqwpvlnr77cmxo7T1u4n/cxJn
zyMk88ktCEZ3ZV9IBvhHpNLADC1wdHn2yT8xTC3aAX3fWpky6ZMu1qkbUbY/gcKR
3GKSJV0wAzwEoc6Fy+5AjNzOp2/WC/N7Y/M3snjK/CcaxpV6Gg7gGUenRMBhr+WF
FXblu8qIK+S6gWbW9DI27mKm0vqEARqRo9KN7U+cA8vCwj/d6rsvcX74nyDIGp9m
kb3ijvSwj6ST6F8zpi2Uycw2gJIsZOxvvcMLbD7z/2r+IvjZ8eOYafsHI80vrX4o
sVBPR6bK29M1ljLj1wTUKFQTpItvTevmyT7McULz/iLHo37Q9rp41rysAMRI6TPj
NgISakIUNdYyV9AlN4phMrrp375vdGR4L0FssCvgW9pgEOZJHsX5EE625hMkvIEo
5Y0ZoSENOkV4KsBy1UPOwU87ZcGX+rQjeyNBvZ0Ic487xBLGKMWeQzn0H6Q1FKSU
/i3ijXiprpV33Z7OuJfOI6g8DcT/AwRNhahYdKH0PoDHn3GZLo3nZR3abwJ6XiFL
BAuipZfTpTdb2v7FBTdlm6ZPx5EVigjy4CpYK2d9sjrmFgreCzjh2hlKUzeQimHa
WX+8a0DFQF04cxeOR6KDfddYbH6X57lBgigUkIsVY7EBASOA6eeyE9c/te5AGxoE
t43QKd/flpPaCL3FaFLSsrZ5JHNP/dC+H/LK2p82NvzgFjFhd7bnb4l5oHkjzSbl
RwHfLTH3IAvfMXRZaiJNwU6N3+JXboIQWKdT9noMJ7InMlMESAvYhg+Rh/BZHeFB
tbNeueFCnKtwfMF26ivXI1t94s9REqHECTdk0bMA54Lae3Lm9nijGZAhrJwz+oxs
+Wo7w0Qk8Kyr/d1maxB9evnqHrC40YTIKpmkP4he5SiyR9tZOnQ1Z74rWAjUxV3q
sahRDgbS6e2MseV/ZRX4a3PyTChsWSbAvuWNeWQc9f5FmxE9a43SSKZ7cgxhkG6a
7FDw39un3DJgwXSqBSQbz51oACA2ascLmcw3HqdHEAgIkn6NJ7J0CrzCaCcBRKja
rxFZl6bFnMvIbinvS9TvakosMhIV/4G0Lkvo5xlz/JUXxosfu4E4bgZ0jh+nxF/v
OuSmETF4DsZ9zMDy1Z0Wgb7oju/5UpN+aSvDnS+IAj31BjekpQXGM9LOtVNE+rxF
oK47jmk/vsTseyR8O/x+k7lZcga10IMuygWTKnsD2sgoeBWcgn5DuNVZbF3GHCkw
MOMrl1Jzt3FBnwSQiaTwu6CikaPKTFDMLYcgTeh4e0OSX4GGO6AlECOkLMTllc6m
Do9R/+mzJ+tvoJO+zGdKJIE2ipX4NKI/xlLp5I0j4dlFhMJqFJ+OG6alaS3qXUTR
eOj/cu8v1PPCRliFSWuKTHDpKf8k6t1a/h2RMpR2Yx8AGxXqPFnTbHI+ZxpJ+hWV
aKAx0GraKOZgCp8ttyKejn65qhw8XDFc7CweC+LdaB6X9aFYzfolpJZs6/yaDgHI
2MmF4T5XNqkkpHUDdSnL55fu4j7ij/X2yzsUXGu3GBhzsGu9++fxOJqK26dKT9z3
VfBSjATelIwNywGwz0PpmFDwA8YjCkD31Du4j3wdXNlrqVv7CuIDd8WRnd13jBdc
wj2ZfInf7FkahtAn+ANU0d/Xum4zMPhnvtmzMFP3GQZE41d1hhMsDDnvAS4T1UEr
JTcwe+kB229gh7aPdMeU754Lqs3/YFpLmzkyIIkZu395yx8LGLLLO9Dm18Yn+rtq
AIkVcMqhGTAPe6myLfSD5ohexq6t2Ybs1ec797aCYJ71yMXWfG8c9fc/EeKswcrv
sePhmXi6X70MuPhsaBu5+CGT2mZssbczUmpajIRq7fG39bcnmhbxCnZRSl0onuqL
o9/XSH3g/PE4oA/ibemx5sKVDvxfhTvOyQiiHayj8oPImdSG3oF2bPK8FWsbUKWl
E0Nya6B2j81RDuZsddR/xW6DRc+HRC3Dcq7MmLB+fRV51XK9CiUV076L4rVLvyYv
qqhSh2htiQLGcYGWw57h6Mqf6VqQuB4louSwkkbKWa7Ss8a0U5yXMKKWEfgP1mMA
4ATAKXfgagjLJrMgvH36oYwKx4qmnQ5G7r6ue+fBVD+/k1KEjDmV7/Ak3G0Ne5UV
SxoRs3tLnyH9nolfuq2uX4Zl3Wyu/oPwtPOnubHVOnihsqPclJYOE1qJXB7rDJyw
YwD7dM9kuJgwWXp9pwhKKVd0BXLybUQfoWFXuqMCvdZIvTV5efSL8beivb++4Uhw
qW+EMP/DY07m8sJoEVj3ky4KagiX2ch1aTcQFweJuDPvSqfFEtOqtkqXUs4NtVOf
vMwGQ7LT9gwi2zSvxRiCMyOMO9I88EE4dYILbF0Ve0aPHC/9eGqR8Q1FqLRde47K
dEG0lXPiPsZYLc+Dhu/k9pdMmx8gE/tJMIuFXoflsLm4im7F2FyJIY7iWfe4kwio
LZdEH8q/HKCnEg8AfqDZiOX0scTCc80t39IFgqJYqXTozSCn0NzvyRGsQ74v6SDM
OSgf9Dm05BTfBuN/akQFS1LhoylxuC03Gg5pBD4oSRjnqV4VtmW8G+wet+mjKB2G
qXETNmiqUsrCy6KJdcu5MPrc0kuj4WOjmANj5LrxF/echdI9AYJ/m2iHE4jnIv+Z
9LyyN3YelhMHvdIUZZgzP3ehh0ADoAY2JlhxEpCi8QZYwXZ+BvjpU9WJlloXr7Y8
5rsO6l6xul/coux/9hFcn3JtELoGrNKaK6MJo8CcYiyoPiP3rsTaGNpBXsFjVIBC
EwwN8pBhp8hT5QzVYB3M7EWkiJ5D/lvhFFfieS88RvwYxtpKt8NMJvl8HyiSnyc3
lqB6I25IQodpXDkS7fcukBQ6+K6cksnuoMkmG4pabPah4oudWJ/XAbkFZzVKYPUf
pVWaVC17wLxx6N+uDT/ljyPDosdRD7fJ+rvi+TagQqmwy8Rq4wYhZrK83WbKhYPy
XNhfS6P+9tp7d5KOPXm029pUkt9eDLHvqgS+FU4pRkXNApSY2QakRv/ISD9Y5uzW
rs2yZ6x+y8DCKC2sG5Ev/vpS+nmaxVZl/JfzWB5TnYu+nscKvwd6TTmgwZ05XJCd
TEYP/t3ZxzzzB9i8Cc6dfYnsY+5QzTJETFQOWmJB3t35tp8gfz2VgVBZCs1FsNaL
6Pq8K1trAH6DfbQfSRxTuRpHHkux9tlnQM3yX/ZHDtmSOhgkNQkKnhR1oq5vnJhK
44vSyBjYz0RE2NIFuribeRwgJkUqzkQIf8OWsWIPPjdnH95d22S2TIzkGdEHXPVp
wTbjTuwRKIPTt9MC4lKpIZEojLelyXiMFv7au1G4pthQjznED4E1iKB56Iak3IFz
O5CQhSMFB5wmnxxQ6QJ9qCoAClxooGo7tr2O8MBv0aLNw51u3ysAf3SRsYJLRQ2Y
4oJ5eIZFRpDD8YiBYXpwZ7l2RbeCskkgEUHxJUQf02+a71ZeW1I5vYDnPfNbS39w
JhdegcX9pt/FVkTFJCg7wL4O2Mulhd52j7r8jstBbdbEDF1hPIaNqUBUveTHRAAA
EbNNcOlNml/eSlpCV+dstdF6WIPVmZs8Wl9tRTb0KD5isxm8geUeK2AyhvSNjHC/
Ps4yhmzP6Caht6GgS6lQsUzfN2lcwn2+x/8bI/PCAelbXGycj+8gMdxRk5IkVO8a
3nUe/yuyPUzKyARk2dQJEG04Afyjt98TyNT2yuhT2KfKxocl1ZYgzvoOhamWg6qr
6uSdSfm8tTKjmhd3kOW/e5H7dyz8KCL+SBuN4Su4BdEcmdsobf+gNNzzpdqzdFeO
wKSecPd6TpvA+T9T2XaUgB7dDgLoqqNF9ncc6tv5cu6mOnNzsQRukkEkVA5nA4mR
JEC++gstKCcg6aHYPInf9OO6eT3OGVYkw4ZxZG7k6hShjW1PrSEx3AvLnH0gLXE8
e2dlB5WigvnPlZa6ETihIUEefPb1Di4EADCeRTUn3XYkdRqP2naYNQDeNT6F55Jo
Kfb6MIkHU9uPXzfV4jmiRvU+bAelXs/jniCgVeQYgZpkqCPo/CkPRaChFlfunIrz
0i2pAL8ReaTwxkVAdxtBwZYmZ30VgzBk19SvkIJZeA1LRcxVkIZsYim9NMaGDeAK
HYvB6p0O9mDP0tXBqb/xsh0ocwgNdjg2rsYJ/KECnIzvnl/QTdZAyNDKjW0PbZ7o
T3QWjWf+N3+EJXsPzmEDfYuiJoR55+paNr4h4UEc8AmzC6vKKtiXgvpEOD3p+Lxh
Vje4/wpLfNm0j4PWupkueQSk3JJLMElah9EXaFcbAwDX73bPq8ZpHYG459Jawx6/
ZNzXAR38VPOCnBhq4WhBSP+Zobuq3NH8c2B1VRpbbK5fOcz4oH9YJSRIqrMxeHj5
UyZ0/iVms4GuawLIVsr+z9nQCCafTILpt+x1L+7xtPKtIPjA3WubE7g0Hq0XldgC
qtj5S74myLnwkrBpj1tT5/dkc3+v96v7fVkYfGNtBUf/MfxVjFLniLMCEMKEVsOp
iQ9whBsWxI8fYxq6OF6HnJsRKckdg41WfPjDekyfc5PkmRVAappq+FoUjBPi9uYL
FCmsZcnVs1hqWt+D4uFDqVaPDMKKALT9UH53qK/0fk8oW1cRlBOR3DgnfhXbADAR
CNMWoCDLuU/rUW48wcA18PK/MMOab+Yxu5DqVBamtL6YAOuxGNwP4JzZvEiSnbjE
nuudbtsWfJuA8tOkjE2SXCP4DXRBUxMqF7zfBJ8NiisovzOQBmbAmJW4KxV560K0
zRQYM4HrMSDw9pHy5VLqYUT8j+y81ydt8bRWpHK3V4RwKYOHBr4Ncty4U7Vs4c/C
4e+NSG57PfC21qQEVubOHIzsppRM1fMArLhHZvdqkuibYH/WDOIXvPM56BsnUTZi
dNmtERARMmLeIB7/2lBGky4ha1Q4WBhT35P/c75MzhoSF7vZheBbQq4sN0eikMDS
X+5h/6c7+/b1sMxWsqvZGyXIvpCODJ4on6/01ZJ03HBAMQ/EJoyqGF3IOpUnWdyA
A87abHWUl9VfOXu0VKoK6hcbEP1/orOrNbdjpWt2dpbNie0QkxYTECH/TtqCTqnf
unCirrakfhY1c6mG99dBrgXsXC3rCvOtvLhHxk6QQSisWkJNfz2JmuxNZwwIqKbu
Z+dJDcR+AKvjv7XduGg9elhRddAm9vcxY1/u/tMHFhwNb5WGV6atQipslewK/oGM
o7tY5UTyDG+qfmqMkVx7yzXIoD0jSussWveu5tuNWdOR+8Qkgf+B3iCGb+kyNGKu
r71IpTikDVTdB919JavZyMadb71FLigCyVNhCg9ShKZA1toMJ5BeeBbVvmAc+snj
CiDsJ7W6j9guMJkRmwEkRqdQfa0dfHSgvEbsT9/UMo6fD8iTKWoizOSEDd8zYKF1
lk8lGte9NflC+spzSitcj81kuImSEMIzBTgeG2HeVYMP+5zKPFuSlgHWSAniyjpw
YJmLhYaph4+8dp7yFelJe6jHS5omio33gwX8YjvikqEy+X6mdaMGJzS49qL4IgrJ
WoN2n6FwPF/2jy9doojHslj8VrOU8F+MFquuDsiJ/PnzxxY/zyuKYkOu77FZefm0
xmdd0LKinbVgCjwj1OcDBkuUWxGF//yRZAWFcGEcMx7QAX2WmUxDZH+fvguwyFWj
k+tiQhI4k5jRKc1NkEAnS0XP3EBlYiHiFg96J08Q2YVh6qAutI6x1+jKnPCjPooV
I8XFak5hljzqk+c+R7iJ32VEnI2AfiwdLRJT/a/ShHLv3tZDmcvZLKau6qhTbun0
RSNz0kT73xUS8EqtBCVrXZbm264xmYpLBnhCuJFAfBx+NwZ+ovUZ9X7IHVGr42xT
l4Pz3N1cdHFSoO11fk3RJe4o3It402LNPOVeLy8cHd0KxxEmUT/fAyPxNKtabrXW
0y1tvGycpU6IBIpdUlZO1PqBfdbQYoo36qsjw/p0X86ehaqtC5MXnrR8i5gJGi9z
tfdikqRnFzgb0SPe3X3yESg+yaPERsH9zqgYwjRd64bBLEZL9cXD52XoPDXx/jOd
jT7Ht/xQ5Is4pF2UIyjt2vo4pLJL3ELcZgglWmoBBTD9DIKMHMPYwBl4WBbP5/+x
36gHZvjMz/i/lcWwGZqxbFy4OA4Fe+GwD/YrdBeiks8j0cM04eWlV1R/XewjH3FR
tLYJAaxrcU33MBhCuNAMadcVBmmzqWhk7z0XMxUHtLrMri0M2EQjDohaLPAYb7BR
u2k+5DyCXBGp9TpU5QGhiuad03ntYdhhSbOgJBYnRCCrhfNxVQlSY4rRRo0GULfc
RXLYp1LFmDqQzeoUM8cg2iWB2+ZZNa6FX7YJ2+/yNOrbZftMSKm9frMUgbGFmc7N
gjEdf7C+VQeMocgZxvR68PW+xNgtLd6vtqWAW1fNYSn3JQ22I8o+uhXz4F078rby
QAyLiDU+8dLpHH2inXs9XUdGWP3hyHwwbQLJNng8gcsp1lkMWADcYvCRbxno23c5
FtVfVq4th1ItyG68uHHTIPl5dxu4z8M/TYSPpAkWzS3h5s5WdkWiUYJs74J62D9A
04wKxJ7q2+aGYGH46RoA5txX3yTllp5DNXLrSa5jK2rzAJKaG7Zlq80PIkXb8kLV
NZlRt2JY4isz9HE7h/St6vZhrAH813Kq/ZaldnK2ZDAfJadwqd/X+35bSdCanXg5
i4OApVnnDBQ3m300FsN/qZM5lvIJ602GPMslepVSTciwxvf2JTWFUMxyvChELw4U
7r/SMWormVprSHYJI+6gxe8xl32n09StDcfhB41MpFX95nxloNq+Md3MtRUAYoM2
LImMFJi33hySNwmGBy8pfORM7ppHojtA90j7f3davaIZdlMp7cFfbp7v8KbgzRWX
GjESy3C93cp6HzxZDg/g01BDqfBIF2aG1sk9Zil0cc1p5lTX080KhRoHmmXPI8sX
NaxTthgpZrhbEXrLsdE+KkRfUWImTGRAKqqQH+hPXiweIJEVkEvEX3roGcNFrLFY
b0mQV0ZK08+URqKzm5YJjc6BW5MAUoBSnY1BjcTSBGDxy+jZQnPGwvZ00TBIlE5b
m/qjyKLiNo57V9/wFNkuKf0UWw16Gcwbz9PEsnuWLe7zUDcbj1GW8XQSgr4BzRRR
4BDo/YyeFgaGDgGEGDc8shKFbX+gST+YXXzRyiCCe8kpGUsRK1Efwn+ErBOdRI4B
VmIPraay/pCydUq8rTI4mIadi+vznU5rbh/loYrPXJ/uIk6ldKVrxLc5eICd4JR9
JnZ6ihP6VI0ONqNM3YCuwiWvFyZPk08a2ht32wSaETchEo4D8PACH63DbFbB2dzq
lGoXOrSYXSStgFzQPjSbHs3B/5f0qynO6vPMyJD7B/ycQsPNsDOcXWieKkrACPAk
rhrOmdEFaTmb5ZtRzS1mg1xA4yoXr0HPxyerQxEpunvCBxJseFZoyN3q6f3FYedM
sQLDWApfEclWh7pA19G2/q1OU/NMIEkI8rCx2g2mjXtwTxk5BAw5BIOsk1auCScH
IBkMbt+KqF+JLGhBf9FHk5MaeFVJ1A6p1/w40FpdH2nYGbGx/4NifxvGWUpqH/aX
FX8J7vvAkVcByqKk6L54jBc0rLgEehEJdLw+Tk6d/iN7Jfa/2rZ/VGA52UnQ+pHe
WxVR5n+LaR8j+ZaiBN4B3Zt/kEtpVncOjJafjWnGtl9rTxCb0a/LivskmM6BNfmC
klV/yt4bIVd9/1nXI1mFLO+1Y3kk2NygOOMV/Cpj9IvfGQ3lld24OVKcYadjjnt1
6rm1knEoNyqcoFpqhXtawc0hY2KN2FtbhRx+tJ5jpOAIttX/AjPiAv9JQkq6PuTk
ulO7Rmh2NtpP230gFOJAMWUzPV32e8K7PQmnEeRlzTc/rtoyADFft9BSP22V6pWq
vZu+Y8xctAElV54JmW4jD9VG6quM4OOMRgwFjjdKSVxLBccjpjYT/ap7pdcxAxNW
+IXtr1E1xECV1QM3jNpGu/qFbgbeadrnNeqbMOaIBhHa9IDBRr1TykEKN3gvvCFH
yNYeNwgcOueD27iLWSVYL5ulgOYJhprK5kj9gMg+SaM2MTAdVZi3nV0RC8HAguIu
YDzmScbg16ED3pLjlzI1p35dnBE045dSqm/oAsXyqGBiEAeBeCA8M+j0qnJng/Cq
HairOARc2eI1revHBNWgTKxYCX+gjAqGi1QiOca3ced9qpx8Lhb18B05Sw9WL17h
VOPUsCGqjJcAjXq66bBzh4MnOfmGjS9ESK46qsMvAQsXEnM6BK57bAAcj+t3fy5E
jGamaOP1jUCB2adDtVf/deBM2BMC0jU2VNFnripd9hx/Utit1uuAT1hY1Swi/n1W
QBygb9t2IPJ18XQEzvo6nl509KRl8GL5R97KTtArzYrf6bVkCayLD2eeRHU5+VEi
YeKJ7pd93O6mOc4uOgeeJgruDnvSaGJPVg0ydUOc7B8mPfaL6frJE3dHG9VpfBw+
OF1eUhKC2FC8HGnK1R6+xx1nIxjMUmenkyJdzewdVAml+WdLHJREtcs/YZCixjkT
gVK9fAnvDMJW8Rpu6/a9gHuUOeCEPxReybBuHrvSXOWd9zjVJ4hCkh++KpQkBZhO
precIrZpSJzjDUVo/QIJOKT0IofEbKP9FR+HWTmQXVV+I0/Y+LQg4XI7aBi8QMqB
vEuKhQoQBy2eI1ptHjZMoCYO/8EIMjePiKW2/ub7RwaflC7MqldI6Cl20JsLyZyk
YqyfJX8P4EGeBIJDCoOzJav4JEFOJbPXZ97vsbUFMMfiWNou4A1nrQI/RxocOzGm
cG6JPQcyY0QQSb/aAShgn05ZD9xdkUuLIEeEdXEUhWosAJE/hwG+r2Uy2/oFRz8P
Jgehy9O9Efuk2p36weEIUcj+0sC0HPcN67SOwleFbnApiQfGlqWe29mrXvN7NI8u
dsXhnTJOFu2pqjL79ggR1GB9F0qEBT+LdMK7Avwf7jRPeH7N1uWUrKyHBgqsduvK
xj98N2MbrcMYEFW8JasWm1tTlogNp3c0CwVTMsDM8wbb6AJgqH6Ow77oS8fmaCYI
W7k5tE+3ux+UP+V6G8j5mKrlfEuUKOpb6l6r/GDAACTHRzmHx7ixTus0QvVInpUA
6Wn3uGq1s++5GAy5VY9sDDz8xQ/hGNqUJVMSc/djsdfCVLnkeASo/PYC/JJEbApv
L9ji3YrsHjNCDPZkRbE20Q5tb7CrkLDY6xXhB/DSCrlDGu1BWQhdPpTdOVqwnS07
w6ksBd5vozHo5wb3iAZ2sNZEaZW4l5PIRypPli6e3FYUuveGcugjlxljAF9CUwd7
6q9XftcmQIBRTNmP2mcNGnsuF1nN5CoAhk/mpiPTgkiiuCO/MxS7eAeSZsgnFiQE
3QW7i4XHL0avuzJG+aLyBNZ85NQqXUOH9MmT6ozkZIUH2wjgA+EVjT+zqtqKnZws
QHrkqdkQyB5pO095ZxfV5YhH8tEZAVyVCHQDhnSUWuTb/Byvu9NFVjyP2Ps+xtQJ
Pg4aGKfWXpfTulD0835C4DusDwpI7t9yEb95Iqxwr6z2p2R32iA59KVtF7nwHenr
x9O2TwLklBviMJ3DhO1H/FyFoPH9t3pCkaoE65JQJ5AJzKaRvede1BSgkfna8A79
PLsZdUl5TDIPngmHbN0Y0/jFLMRusj7OAu5SNkuFO2eGxOP20dXidco39Xv+Jn+q
MT4I9VCj5I1MgRWLomLEJEaMYG7eeeIvrRVfbkwgp3Ph/QxtRZ9Qm0tqQT/TGVIY
LfVBp4JBnqFurDOtKFRpyn0oOXT2XUPpp1KPNemv2HAH5PY58n/4jL67X1jkh/Gf
kGq7pLPv05Fh+vPMQFJ6VHOp5kwkXDg3BTn3fYdCKUp73wooNFMt5rLZQ2NnmNgK
tiVuWU1v8kFf0wXedFJ8/NouK8cGCOvEyJJPtwLHG/6Df5V9ov/+kVHRa3qmZMsN
NHHeDnD+8EHjc8OVKKqYH7kiFmG9fKcvMxzg1ye3Qn83wv9Pg12PG12crt9zFw9e
casvb+6soQAllDD8Kaoa5kn8CUOmc4g/JIrNSPyVJgeYJgFuhy952wcYVH+JCiod
idnqkrC4z57VQGWUcFAdenvqe/og+8D5NqBbmkjiyDOINmIaQZVBeuTPMV/pUKXq
afCHvWSiM4XrWp/UwEMpVGuymposzLuhLFxOA5PGBfK6jaB0BDuU1VeHDHItCKHL
IzrjLzGdd9eVHqvC0ozgPf/DlbVVaTxbC33BzVVnpbxNlsZn2zxxCmL9wkTi6k0u
skPtEUa+VQt6cd7/EH4K6FbOvo9GGSaz9SRsidrHh7RQWQMr/4mhzyWZyNHTTiXZ
FqwIW1lJI5XtGu1Y528iAzjOMpB8gpJ3YdkWGFfGzf1IqjQNqi7uRKzLOipIZ8Ja
yx8AewXKc70qX/Vzdp359c8PCfcf1VdGAdwy9mYFU+10HFzbT/NrmzOH7ovFYL3I
VH2PxuppwspTrRCNDyfh9BLJT450ar6/piZ8DiiII+53c/0SR7rtrMcZKAw05aRH
ubvHT1UQUX7zi1kG6dk1VD+HjB+peOXdFRPYdB2a3qb+eV3yQcwCHROjE1Wbhs+X
AH/BzSK33MWgapG2pbPuxkvLGrTKPe4ryfjU5a6enV8Zotbxgfeb2UXFw4bglnGh
xkJR5Nu2udpBQpELFQ4EGLOrMnIdZBRRtFjvZW/GQq9Ixw4HYijSv4t0tAP+rH0J
P+uVZDucmMYNaWfQoGQb2ja5PKEIc7kYs14ZTiWpNgxiGY+MlV0vGT86fR9cwMFZ
M3TgcWAb5M03iMbeWhgf+zYpeuSAxrH1afCebIXmQ7N5CZP2q1SFKHZT+p746EDY
6M64x9V3OEHXcouYdTFJPIeugoHsn1rJHLGXF8SG0cLYGHrPTmaVclILBizv72pk
i5pUE6GMBV7KRlJS5fsnFk4SKi3i4DEPzjL4JhB5KqDveBa+Gse8cq0LcBHZ1MJK
TKvqfGOY4P67smDfRisB5k/RtjQxHI8OfbdyMMgyR+nh4bg3lg0H0vue61BvDkN6
PKaMwFMylwpjGuZZeaLdqHWo7/dXaAreZPYTT9I4vCPyHo7P0nY/wFzHWLGn2Zhw
U+2N6PVM+a2AUdHUlFc1xOgZwmk/xdza/E7p6IWB7mWB7hEvQitOyPoOkBgH5AdN
KauFCJA90HUIos7+4/HVQzBPpyWS3gBdu1yafiMN/KRKiu7PUSyY6ejylgZcXDmQ
DzPXny24ojN/no82YOwI9Xj3ZXawjTnDeot6FwWPZTgtDd0dUgf6m4768k4EFqfC
HL8HvHJijTpCxKR5y/qAXW2Pj01er0KwznSJIe3gh/YY8kVwuOXPv+Z7q+bPBsrm
VhVV/yCAI3fif0Jc7odpiWVYdSnSKD7Ao0h5CkQWsUbtaeilSxqu5iMPBIBhgBKc
BVtcu/F38rJVLCX/jJSa8pUFpCCH0H7xX8kdwA4NnVDZJVeE1otgGwOWmxIQPk9t
CdU3AXskHdbtbwXc07wKdMwtKcXOk1+2h8254b5Sj724Sz8G7ND0+35X1kUNJpfn
HkkdqqxdjeZsDIx5B5867DDHbSrj7XlhYK5WoIwg+D6mXS8ZHirtD06EKgF4u3JH
bgcMfEDofPtc7lDsxX4rZNIkTY8mmqDWvY70KAceU/+/Bl1st3fBSvl6wL+Pojf8
HLgCi7JHthxagAfrbdUwoJVlYMop45lHo5vjfMDcCg2hGF/PTRjYAKOtcjOoQ8g8
HFhFt8ge0Dw1gXqAju/O/ks3+39znYQySgtSwr5LjuwkWbt4/VybgEqEJ0a7+R22
fNflCEkARDxBBBw8SQMdbqoIvrzclFqV/yOh17lfbb1ukbpaKSEDN+1TEhEbVMk6
xUBZcc5KQyiZm1Pw/1aDIF8lEux7JEKw81PQvyjd355k+P8CrjBP9/EaQo9R8xKm
1hpSUmnP8zUpsdlDUAxy3bK5KOvbvgzWSm4sOCvTzUWwNF71rLgjYx5INnzcuAFP
qc0KF9UR9ZHiBlOvDnhUClBWsCOIVdanmBwAkPUrImgz4FJxK9CnXdsM3PXHxWnE
VBqJsLBaAcTIknKaenma/JDV6G9D75m1sddhUrb7zpkQ+1DUBYpju7Awmuxtl8a2
4PLOC9UHnVHnCvwb1sxN2wGG9W1mZJmrOSqYgwlbnU63cX+oD59AsyUV4tgNPOi0
gqzmyJvkUWUAJuVx2KptjU+aZKM4uOstWQPgtu5tUc1GNBRsWjdyK6oTA1jyvjiv
qIOFF4+U83n/fr7dKx+Kx0w+ddFqZmfRyeY+ACo3YmcF5F0o6sXLRs8ILkXqxQcQ
NWRtIETRRBMUNZs89cxgAfDbgTLdGNZhgQ2jMpPciN+/Ux6NMPPUTMUJKIHAV2aB
jpB8mPOkZppwVC7+1Zx2v1aOo4C8lbSvtWuEZJ1oHpCI00hp2y0xKDOS4Ua311/t
5FgC+3qXiD8ak5mttfc1+IK/1HjIVdcMBwsqsF1uKlJSzwGTKBt7uIhDC3ozJX4f
qCHjYl2owlr11DKdx2iPDkynI78nxCFhEfaZq/w8ukOnGSJeVZgECknrEQBXOFi0
pt7tvZtnKPT0YH4qAmvT6l9DRsWb24adBGZYpzKoJzdSj/6IuHAOFH4cOttnFnNd
nk8AanoK39ro/8QvBTp2coG9xw17r1LAZLwpYiUJm5RZxoA0CUn1BCOH0+C27q+q
DCpnZaXWm8EzO4HXhbX/Ee76fLp2CZK0RpcfUycAkLKT5sKk9l5vF4xk2rz+EEO3
lrHu+EO6lpNUlKPWGiA3KxvyDgwv0gsZeq7azKX7WrKgvVXJSovbQS+Up8R+0IRi
r2NtXa7FCtRraWHS8NWct+OWVlbbMZ8wwAKRFeNLo6AhXs+w6LQewG6NJnhPjmTd
PFZ4VY6bzaHddyIIsh8d0TZC9V1K+XAFJx703E2sO1Dh8FZfspPItSGtdR/DKbmD
9f3RtwkAyYFKWI31bGUKuXFs0/nd6ZcsQl62N/b7l5w0UJL1X7KSL0F1XloMwsu/
Ox18kD2AGnQRPZaMNovFhtxlYi5fN4g5kH3EYnc+dydg125ZRWsGU5Tqjfp5HwEu
lgBrPtpKwladZ/eN8JAirDHAh6lox6CwkSfkpPfi953Z1NeC29WW8RMD1QwqfQz8
6pHz9NtbTWc8Sfq5ZXcwdfAqs1OFVJu1IaWJsIdlFFk6yBweGrZAemA0uF1Yeq8u
GIOTaUMOw1u56rCLNWvECEXoY0iIRp0fJFHXrr+bnWCyw87G+w4i7IcFAK6SDWTM
TFDVTn3Qux8dB/g+1DklxGwEoPOCU7YbGF2pzU0N47M8Yp7Bdu1KylCaEz81pB3t
1zgR67cwsDUFR9hA3oSk1doItInpGkLCTojHL6cc0XampuUBrkq6t8GZw5yT/9J0
ijeKUV6AmwXuAFaMovhXsXErSkzuFq2Pf2TY4NGuI0LhtNoFrILqVt3WgslcfRFO
SbwA05aWMwzE3JNM4O+mw/SUKsjiKKjRFSCwi+cPGkcQyzXeN1yPlw2zuYBDFtSG
fLP2tyDQ7LGyOA0kEDq6QepU3jWlYfojR2g678KyNq3NCpOyT/33MQmVmJ004GCM
8j3g55OPdgpKgkIHSpc8Qlnhh+OtEHuGnCFNAverkniSoc43m+1fe720X/dxCKb3
giKquw3TkznXbbPBZbBBGqgnE0hIpouId4ldIEMEyq2b7jFi9GVoViavX3u2oH3H
ItjgpUvJcDoRmcx6FFwENhfpUXwhnpQWoADRwHMGtL8AkMiY+bCCJeOAtzTvV77D
JWq1FzqxDgoZt4mA0d6Nf2RBpkZuFBm2sUdDIE/pRzOu/RpLlo509zCB6yTN+wN+
cc5HlI6SELKUxl5U5Ecl5LbLcMQsHBueKMzVVqA4uWdIczT+OQtubYyWwKwMxYNs
+11bgu6BWqPg//Tr8NGvCn7tL/vZ+DKzTWeJbo6KDMSxJPpcgXha8byfNgMfwuLA
PuSzy3D9N7iem9wP8g4fn0zv4Z0g/KlMCGHTxym1QEdNWWSkvDCGs8873RgC0Sb2
oTDu0RKmFaNvHC8fZsMZXvFBKNty7ZCLNdEsX8YV+ZDBYn48ntTuI4xXS+6Dr8Ds
zNz2C0GI3g0UyW1P3kE81abFez4OtxO2lgZg/1tc+xr6zZ3Evu+c+KdNOxpuhvzN
006tFJmwc7ZcV2tEBwD2R80PnEQNzhqWWwIpNrsfWM3odkvNxDbRrVNk2Z0PCmyh
ISa4etl9midwfSjUVplWy6UvoxVQ2vSHU/GAFuR5isX5WnOS/ZSpWGc47YunVcJ4
Nab/PBa0r5OzhjFuMpYz4eT/mEewdnVo4Bux5UDG8T+xtm4oL7W018hhigC49U7J
cBY42ZryYsTPLgf+LbH7Va4uMP3XNy68Z3DpntO1BACpkeox0gA//mOgPBTnhvZZ
hp3ydYXKzb5mg8n4F3K0ufPi8Q8PECxgOML3RZM73UdiEL3w4GMzLcDAt30thThm
gC7Jtg/jVySAJhxSo5D8PWQKtouioqVYMeKjGOOmfMj1lkVmymnrQRDtQPX7c2H4
bgoBAjB95lIenfhV9ZL8rQuQ6HBLip8n9/w1TR7uusOrp0bRBQ0BoL3197YsT+ya
Y5ip9DcKMcRFDwnWqlee9oh8K9xb7tV51yzGfLofeaAK6LCuURu1kfeAM70jLS6S
hM/vT1bknXP8jWNWPFYOeEo9q0iidfQBjQIqahXWPuz8ky1L/+0QgNqoWqD12/U8
wvNWVjEJH/QOu0Mveqkt51lpWRBcy+jTtBrPu6U86aBRnx+b4ioPH6yKFO6AfZ+S
vOUXbn2BG2WPXmNN6WkPDCY4ft5hxC2XNrkRgW2LLJSeK4OsNJWjCu/GmvUaIqvI
s3JoLb+ZXNV1TrGj3F5WzeHtWuc8GLTAh8uHPY9UXN3Tjw6e42zBYaK80b9FcNC/
GQDofqNRLX1jWXfyYAvgV69epEu8Ol6+fXLADdzl8F4AnGarLKa5hMls2U+xu7np
QmqlTa89yn2G6T4+1lYOMqCpnKcfd+rKpdg7ejnJyhZbZYvjIIahgOnW8oSwpgXt
Jo7he0nmEXaIqya+rH85LUppXKI4ZgnTwGvdIkiAmsALu8McO/yNULoepOhwrCH/
R1eI2/kkGUwXWtv+sW/R4W4KdHUyMzg3FVMdCUbzP/pPln3TABo7gihW9qtuO1u0
O4UyA41HUzYveFjM6uZY99hbdp+0ft5OIazXqGygFWwC6JNNGrOBOxU4mh82Vr4k
bGBFndHAAP7eNO4vOdJvfTJUpXwoe709g8SstQsLaF7bDQua9VFQIZ5z8//VtpRu
gPp80KTl87Of0CxBwrzgoI/Q8uE67Uig0HfiVj2FZIQNlpcHzeSUqHY2xw2gGK7/
FDmiE3N2+ypgRGuVFhLkX+fOmpelYHf+rKvIZ/PnmEnFs1PmtIWEX5+MBLenfoRu
qEN865IgMG7RodcZCVrWj2G+Ih3jkNpmR3mMuwxzcWdka15GxrAETmqkNiWv1CF+
HFrCW4lYVVh7Vu9eHC7waLtkV1/rlWvo0bPisrhXhzDVT47unh/ktw/7t32/gP22
F0RwJgm8cGyQTWhS5+pHFXQeip/08psX/AIut7Ph9BFcC/40cPIfiQNxcwvwfqYV
ZRdKSKESfSINUCst5KlOoFBa2QbDCZS3wMV79bOwHGigys9fRIwjtT3SZ5lvT8RK
BhgeCKFxGrD8gybK/26f0T6xmuJrlD+IUFASD0NWpkJXI7MsCcU7aAhBkFw+u3IH
BQu3vUd11/3MtINmM/iJmsc9jLEuUpdDt1U94QCRtSfipwgtPfWliil/VxomhGlk
LrPW/o+aAUsyk7CEwoECNa2488hy7v6NszD58j7JtKKjZWTmrs8DOWwXVl5h8+aA
YaPFUpr1qibq5B5hF9I4zajim62MQuO5XCb1/c/km6iG9zhi2TseChi4TcqFyjdR
usHvLAOIx7PWyuKg9bpeGKkf/PvL55GL7dn4XyRsED10CrXJxKyNDeKkIatQSeXn
kgby85Qjahjjwcwfs8xQf+VUodIDxv5m20YCBBWoRztuGA4asXORHRybyjADyvHh
OjADrC9BZPTp5wVHkTfNkjDhfWTcpxFykiHeY9KaCsck3u7hjHm5hQiUf7aJeEQ0
MKIWr3Vp6t5eJfoE5nNnGvO0KB1ZI2nvskvfedMIarp8rPwLkKL6/qMZvtKY2nIO
GCxei2kwWKtqZOPL051uDZ7Nq23l5Ctswpcujn9b52vc5s9k97Wu53xd+e0CTdg3
2+XWBMitUs68neo5sPADcBmfdvKi+QxnZn7FNdUPLf/iPyG42Y7JffeFAxVeDdRV
fn1eh0OrfmEvQu6fVDgb3yaxI2peLxGc2LHSJkUxve+iMIpXzw6WLDzp+t+hqNc0
vW4BMCZMiWtiiaYXOZCEOOzYtWPA3Cn+RzGV0ARJtsm1e2RK4IejMOaA3w+HqeCH
xGWPokbRN5RXbMpNb2sAbU5bTaYMB8P+UsBVSCP6yRPl5MF7C3YgP+JvF+KEVlin
goVBTLnor6ZvlAGYVKVOnU5rUPDVzKXj4TgbODS+vKdxG9U9OfAer17mteR6MfX5
8WsJCzf13blTI1YjxLh1sRZrWU/LsKaLbhvNXln2thaMZjqkozp74mh5qGVhdH0B
YTOfqzX2PPz2btd/QGF8WasBVT+vzT1wAsimjj3JzkuB1T8g9vwpKeCHtKRNrLnA
5znpfvStaSu25DzhuSLVEVvP3lqnTb5SjIV4aBMX70VHIuINhv6BBkhphpsR/l9T
savq4JgePe6yt1JIbkjkWGFI4ikRaxxEul1WWBJ2qjlgOWL4P23tJC/T8Ql9DEmu
yc1VOvOqhxBOFuzy0rb7i5v1qemBkFBepcmAL0uc8ykBALPOeMRg5rTXtwRjBHef
a8MYaMVNIrILQcchgsiHlMvslBhfYAH3r1Cgl4EdR/T4YKJPvqw8GUlYd94vAVrU
F7zqDMAHMlJ3gc5F8X1uO2ULikHmbzqBQI9EwkOy7tOVqbyo9exSP79ZxL4mMMZU
M32RBvLC8Ka2QrZEBStyUvA4V0K3cGM3rkgJWvuqjjHqkMrWzna89u/q3hXYmI3j
kcSJdS74/pXimtg4sI4dNqNBGQqyZFJ9PM+7EC6l/CM+Qaf7uYwzuMqXLkm3szsC
7sggS13xXib5lxqs08P4s3LieRwRIuztpainfS5yzNBU2hzonYiuHdAZoReA0Txn
FLeJ3n+wcdkxbVuzsv/4jF+ZJXqeppiW3okdFvkGl6g+o5l5WyE3nBHzS7VZ3KrO
VVUeNad6xhOBTvJgjGPyxbaNCPJVpnASSC95HfRYJ9FOEs+w4r2omVGE0ROYxJRu
oVUwWBmnWqu/DfIFMc+ZANqdBMemOZBR1XSOw8VrPNiLsi+g2/bwT3eiZiC8miiY
eykhzxivtuGLuVDTNYkl4ARVP7U9CZcEHfvu0NF9SqlFXq9TCd7tBCmcgqAmdfFE
UTo5041nWjv6CmPGKdYVEL2n+7O2aqynrQ+WfTg+3+0kjUPU8uRbVvILpzJLohHK
f2fseEfd7MhkP5OTjERoobb/muy2JtLFIHPf0aumcGMeUcR1IkWy7t/NzM7RqxPT
rzuvPUCgB25pWoV57yV0b0EagHLyMV6OcwLDERkcw6UMN1PSr1p9J9nnRr83rpPz
0aR6M0sx2RDaMCWe+gKBB8kH+q7QhjqjFfrJRyZfSH7326Yr8nCwawoHrCLeg3Bj
vXtWrVzIqqRPF4pBJ+jSXIossLR45khYLXCO2GFStVAJZRNbnRBSu0KQbfjWTTiU
uVstXFyfXGwh1gPPwLn/SOcMAxrO7POCp/8lAaJSu/V8uTEhxUPRyZQaxXOb1hVB
eTYHgkfZwl6Vt5gSD24BxPtP50P2XgEvuaoBkm6w5cBYZRXKyBsC8EEAx/B7K8yF
EyO98Lov7Lhj2ySm+wAb/noqsDAti99ig+y7ADQPAU9L/6d4U6r8o/KPw2rOXFKB
w3D6IHHtH6Ls/+zR8zoMPfhB7zl/hFbSJcyHIQWIZldQQcDrwq7z3lZuQmq4kFK1
gPjBXMdyKemPQt0ZuRIDFXquA33C+VqSkjneefFFzi44ci/jCqi5/ZY6p5WOuHGG
0ZM/W3cyULnyXOmY6y1LpC0ddmcbTdnFtfV6vFEtW0SfZMBVM2pIII6uVpw8H1pg
j2dEAS2Cc34Z2feTmT3U4vZjZvlkgbDRJCyrJ0vh7IM0pWP06e/WGgfKqb4vapza
mQwMlamB3Fpc8D2KTsli/utxmUXaUzru8LZ0qg7X7NcsMcnsjrRLfJosYNp99Amu
ZtgoU/txNrMCEgvHCQWHdZayk5iUyst86BKdBVJ3mLr7vOZw1xFnCVvCmdbqWBIg
h0MMvAZ4gxe47Hh4nxPxfPSkamA+Y3tS7UHxZp/SSejcYwFvynbnTkTLMXuRhZrO
ASjIkXhyboE3Ojk9pIW3BUyrGdV5rZKx9VJkkMhbtwyw7B38SfPyftI/ZZCHpfTZ
Lae/c9bdozAhdWYqlLwTCefllkVirdyJinHLkfwSVB++N0mqkqStwYxk0iSEleuN
SMxWYipwnFI7FDHF+fHzlVoXh2THAbP93dJT27IZmA63lLneY8UffkBqibjwcWDa
IpMdKLRvuF1DfM+qcc+EbLsaKkb3T4r7tD3FgAEl4sIJkzjH5ZHYDrIXCASptmuO
oif+YM1+tOjBLEeEmvJcIXHYyZnIjjfZ7Is+30t66zLvukal6GkQanFq8U8UGBJH
TkWtkxI+ANqiWXxAvOzqO50ex9vsZxuWqF0+nNLoNsWF0uzThtgn1u2njl9z2gZK
3SIlffm5ph8naj+nlDNQzoQoz/MqM1viMyxKL/bzxXGsfRdleg9I82dtc6f0QBJw
eVL98ZnXvKfMG9Q3Eg2yqB4BvPryBCQLHaUnkE3z3EsdgRYUXw5WDg1/LjWbGerm
x+UBGXF616PB5fGvYPraeKb0CS2PwG0EV2df0DNDHhc7JQo3oKqFlaAyDfOCwPyA
nvwntJU53HoOXupM6YF0jQttc/WfsYJAWtRD6h9vqTMgGSmkGU0HyydCTrQ1wZSi
wLBUI6+PPnic3K/jnvc6fVsRsPrZrT43P8LrHu6l29Lxr5TTN/DvA27nyYA1OnQt
E7NnL49YEMLTAKYz3XLnmhnSd3N9MKxJJ0cR0HdsFt3CKV/CzvuK+DJddTvPNq8y
UssqAKZvzkbZI4++TzqfGt4Z2JsHPDb/mfldgr7zALDEHzBMejFFvmXSzIu1ctRA
zJYA8yyEFdxDCRxOoIS2dvZRnHi2XMMF1IpNbbEs1AKmexf9w39d+AWhBMKQytsV
M0yLMMrzYeOMtphfbQ4Zp3NvQ/8LdqGzIgRhVJQqxk+0TRreOORaHDfY7N1+kaIy
ZKM+gq4Lf+6j+3o9qJWyWD29wsAqs/c+H1Z2Yk43E98lauxOMcHsS8uXdJx4Wbu1
1AJ1Gvnptvu56M3ZJ6/S3aQOZYcVi1MafC+j13363OeSzvJjvU+MColXD7Vp6Zyt
5j8nUpprrgnSygRNm2rwJcLFd7IwGJZMowcHdjqaMXqJUFbGAMJ2uKzLIzemQgDG
T3yP7QpQb8RMD5OX5w49ZTxrSTi7WGht3Z2B1wjPviuOtoeRH29INuZFbfA4G8xV
okPtt2Yr2Za65iziAWkIk97FC1y9zM+IJsGTBRLeha4lZvpJbOk83Nvhri0RJFgQ
0VP+mYKa7MQTEACKsxi6/afOA1apY8MMmbqmFAjTIvTyHmWf0DBdpPaSY4Mdblbc
HKON+vyUI4zrx59vtXz4l7+W1jrIwfnU2IxO64jrhvTMGR0Bi5wWObh686zVRdlR
wwYDyRh68SWNdaKNvamns9RmRmXeb8elxBceIEGo1m9eAKbDOdFCCguuueI2DlAc
851j2kCUiMKLV/S/7GAK/rwadIZg11wLdfJjZeuxzH01yuD0c9qiQ97pvLIloJ1s
//vAjx15LmAV6eA931XOs67+66B6l8ofGcGEnqD2nYBiptMi15mMXvPrRKTecGgL
gRYo0d2WDL9kgBvyWDJJ5vjXj7H316CmuYnZg2De2iG4nvX5GXjBSO0mX0wdJe4L
0N0H7D9Tmr+lGkksCerBAOVCA6KmJvNPLrGkHqvQ91kWtYn8yvcLHBDrN5E7CvaJ
fcpkZFfP/K66iGn+zylIjSkpma7kJyHjUuGppTd0b4zoUPiP6UG2Vf92DMASkOST
IW6egDpp502uMLnNcPlESOHUiN2t7IlnW1s582KaPgh5yDSIxGiruaQ6uHMTRfiL
7iUMcFUmhrCDZtJlg73F2zIYh6qE6lAfsjWHjQeR3VUuLGPT5xWU9ip8W4O5UYFK
FFewPvOcytyic6J62WDJdXjnnakc/YcK2wLw1NeTMtQxoFw8QPAOqrVm6bf/oxvE
7QSkkJf0c5KwGmmIaVoFJcZphTlOtwIHhIG6wWkuUFVLVf/P/ilsaOoREquipuVe
LRHbT1oDWHHkEJHIxwqtdvIRdqHIVugbcVB951V58GC2kV/R1s7IqEMJYL3Vcd8o
wdYoDQ2NVBPGjCvILG2ZCTt9g+BzOVAruA9KNcUMrFfH0zqgmQLjTwLc/rp9cFb0
J38h2YCVaT6/V58RyjetVY85Pp0E/m6ggjNtdLqzuBTATBgPvTiyVhzXvTKKVicp
vvzfGD43EkmIGJaHY/PaliSFMyU2zSrND/tgPWCM85LQBtUAnwBvS8BnQprvUnTQ
qycMFCVpDpHRyW9smi5UexHLh0QuUJUJi3AzljFU6z7TOlhGDT4vq3TjuK5kX6tg
oMnmpaDWLq5Tzo2//9B8cOedxRsqRoi4G66+Di4QEXZ2ABfB5SAgQTnY2VcpnrUC
5CTZ0rxkdTgujLZTSFn+Kttkoy/g3AEwEf6pRfhagaDgtwYOQS6M1oBWWraCagsb
HscK5OeCmM3572NJ0KyFcSdP+sjUHYAsHpQshvX392DEDf93WqEUvvrh9r3MsZ4y
W1SiPA+VntY7I8gtB5GOl13bU0sv0/L0MlPlIMAcVN86EuagAqeAOjH0qrCGVlO3
l7xsuomPFwhZ9l/d5y5oOQ+xqKuJsb1RyFx0gktcyYhHsV5YlDEy0P4+TdDm2UA7
XESbVJ0dgIn9RqU+lLqOBrFsXQUrf0aFV823k/TtIQt9y3tzggTpMmfDIL5xKP0B
AKPLYGsuMN+pGsJ6tedln+PcY37k/ggU9OVKEinaukZbVJABHv0s2drmCktqypML
TRph/8kRroEQa+LVSMkm3lthXrUQqO4kGjJcebS+/rVBX74CP3DsNeCDI06VKjr5
i7qPL3xvM7webvxZMwmyWt8k1IiYxxO57Q2Is2MzRJB1coc+MfbcllwCQwrsd+SZ
8HO0bKao2sDh2AR3FVAVJaW56alHjqOt96x9aCvIOqVTfAHzh4EeefoiOzEGv9PQ
1v4YneGrSZCT2D9t4xS/MMs8V8Bph4oj4JU+R43rlLqcvVWrwi8e75b7j3PYoggp
Z/FuLSiijUOq5XE+pecYyYumoHcv7l+8gkMNeE4ZYqIhCPcg73/1J/rmPuyf9vRz
lijx2UCJ5UVyy6+s3DVG5wkac1bmDevk2KmaLC0iamIC8/b4SeXMMHzEFbDW1NTf
o8O7ep94uX97aCGeOkIriJ+2kh5VG94oChCvDUfqSNuCX0CtVrkQUhTJUt7WzBYF
6g2avcqrWmRM7eyB4LSDIq76/mIBseW/RDx66aA6EBeEXdn8SFqM+22QtkMBzhC0
VK70M8mKgGSSEcQ5XUPy94n4ygjBMOpINUCd+v3T4ivylvRKMaNQ6KOE2z0rCu8Y
w9l/TRuarKthMtehzWXzIpRyolCaWIY2pALgr9HD+Ai6p9PXjHjMQRGmJimFFIJa
/go5rnsDuewrKmZ6P2XNr1o1j9EcsgSk6jgyqWDzy32WzWpjdEPCR4NKkKagxNWH
mApFVBZhOA4S/xhMSqlxeKkVH3/jogMPqigQpoDKj4k7jsbWXYpdGMuzv4RoGkh+
Tv18YzrQm9I2mHbROpLTZL+naR+oNWXZyfOQ+Twz9YsuE2cnQB/oYbpmkXFocKV8
O38u8tz021v2Q1snU0dVJj1YE9jcXlMFpxPBMtgKSE+6OQrKRUSYxTzkPtApOkgb
W8Xq3OdGRYe6VUFGzDseuxGhsHunPfsKbxI95N0GrkpjQEQJ8RXlaFr1+mH/h8i5
O28HlLMnPozIbX7aOCniAdbPYEdr0a2vwjo5O3gZJFbqCNY/b9F9DP6QQiDgU+8+
4Kwz4NGH60FTZ20UmJLdSKAvUKAksYEFzBhpbaEn69+3ybgL1hYzvjRzUXv3lpOB
raFXKc0k5Qwwkpu2yrTHXi+BNKEAuSy/wfoBZoOWEhK/TMBOCAHc4wufD+CdKpri
dI4qwFhM8ov2O4LYOQrt57fAT0oh/lz8pmmC3m6vcrMQrD+/o/KLS36pgt/RmSMO
CgurypxyB1fwv/GOqys/bhsNOrD9Gk/8gTi1j5dDe8gpKVUnFsclTN68B+yXqk7I
TMfz9YNTnij8pCoZLKs7f7D7/zZ84v0CSMZ8uQrWUHpvnSNTPotCf9lrQJgkVxcZ
6iPExapeKpipZb21UfRwcbMQYvDjoo+ICo5yvlzqS+fDxwn465iQ+IRim3n82RTD
LCHcyFG/ZYZOuz3pjBMpvHuUsBKDb0gJPyHhH/GIXQW0rS/mNQtgFjGSwfCXvyNj
RWnHUYmf16T+rzsjqOa0An4B4XfRj9wYo7ExRxt5uvdfro6zDH20V7Bdsba4GIdw
zpUCozjZ+y2eDVzWEcEZx5ouIr5gfEkvh0VKHgfwNDfRZjCvm+BWaXnDR9mI6sBP
ZJoGrF4G6DdUUrWpQxW5Y8AXK2APw72Slpx71tjr6fbl6ShzOxHPmvMQ4dyyYYz+
Y+ryH3iffll7Il8ZDjUbfG7Qeq0vEHG0nLNnnUgJwhH7N6Vcb4DPbdQYm0uldwL2
hpNXDPe0/ghTgRw4/pp9ZbVeaAuyS31gX2xG8NYvn5RLTzDmJgi7dHrfHLk+ZZuB
JUHaLZs8CtnMyIH2pLmfG0yZUAgq2sGLDD81Mu2dBGYqqBltQxfOEEr8L65S3nNk
MESJWegBG4ogtm21Wj4BvBFkVYagi+JyNozDbwowjw2Td+45GmO9htLgvWq4myOW
PaI1XklrMvKR5zPu4Y7eePwPqVaz33Hg3HBIhkNVvbpad5OvfkxkhPRS+wHQw32m
QGNA9HGjQMet4kMFtz/YivRodUUitAfVWlJ+tmzzDCJNBMuKae2z1jLzonAwv0zm
rul0eQpKBHkcDzb2QoVjPAJb73JXj0GW7jWi3Tsqg0dtqY+QBm/C5jV5YAW0da6M
9Y4tfMX3z7Wy6DN/Tzs7gmZAuIesW78tM6dZ2XuLdcEBu/xBpNGf+o3YqiAv8BnX
rAiWOhQ/+n+f9Fe55NixospW4EL/h/krGzpdYK7r/MiyYe+kzlU81PmtBJTUfjQx
uqS+Ggts8z9vq1vPx+JZfU7Q3NbMyIUelG9rVRRYY6H0dkYjow3oJb1vVnlyy5rE
x8hhaGZjCyJZl3G1zULOhzHmg32utHD/nD4/dmIF/3c1a5PsG10vpZvDxgnQbH1Z
BCLLBunqnjZ+Ii6mhybsGqIF0INGoB0JZY9BHZ53PC7yAfDBoRXv+M5CdgCp9WfW
znhxtSWhARFJeOiConMfkyPVG+ziVeThXdqFU3VX9n3qrht5yE/uZ83s5EFxYpwK
d24pEHilP1qo6liYOmBkNQTGrlShohjciozDejfPp3HPF/01QiAmtWISzEd67kvm
m3wZZ8vvl3VbWWh2WYgGMrRaHBGkHmzBNbcfgD0kEQM9yCBfMMutC+Lqts8qO+t4
gDiU67xRHxOXdrZn6TBe5PzP8CPtgoy92Q2zjCfBA2ThInObjvtuNENEsOukWgn0
7rKCxLlNkD47SJrkneX8kwMYE0FlQedzGQlH/HhXwgN9k0ydXS950vn8eyjX6ggy
Qk4bnNMNdM2fZi0Yo3bEmx4aIOI6XrVVXFQlVYrvtYMs+IcSYrY2R9elONYn4Viw
YsrPUGw0GbRZNgAh2BdUAwO4dWIrf5sv+ZxbTP95HD1ibfCnnGZP9hxtuh9kUsd6
WBGG0WNgLJA/AEYghRiydJ3SzL9T83y3M0DDNZoU3RL6OEuyjWTEujSIRJtfX83Y
AyTQyEyQW/1qp2zivDWVzVfrh/hD4Cvosu0/AOKrbKy1iekvGsEBePsG1Nr1SnJQ
fHJCyxfAv0idMFXZRuKqKYETivyMNhh1b+b8P5eIKXQ8HhyZI4uOCFmUnrce/XZx
PwwwHtjiKkxohrSvogGT4scfvddx6Xko4mswyWrZKpdo7CmGyM0s34bADlzw2Pbf
YJ9gbB4uWZL3kZO97VqVDfN6ZTagoWgDrl0iY2v1dBT/cH1kNJCCpS/Oheum1he1
iJobZMPvBUGui7ZGsBz9K7GHVkSzN5Ei1HJ1yc0ctUimxxMn/2VGLPDEOkfE+PYH
4WEzlJ1YJUY+3YUz+Dtz6UsYqtHqFQDYC7STloNTx6ouzTEc/ekltoDZRUUNJwaS
3B+BdFtSkaMGccLlVC21n2FkJs3vZQPghyslzHtEjywDDFdd5cVvuUPpQGdHxHKh
63glgwM5ODueWdfn/EiD7+oa2IC07dcIW51oP5VVRkxoOast7luiqM1zAPLvvhhx
PvVy56JV8jddY5y52fSWIFWXRl0v1GvnrMRSmTcI7oSH47xgbnrsfIiBSRlodCr0
/CYL/lzG5rT1rgeItz4uNjs4UwIIDzT9NASVkl4MRNU4gOk4DJ8BgHocDdd0HWpI
naWZCLb+pfZvRs0rHUEwzYFXFekTZyHMnD4a4zMPzoHOhWo7gtzE18g3SMzblljx
JxdhcdKTB84/GUl4+ygoC9lS3xya1IWrvtb4qzybeGXY2WPGgEzPh3sPd6ek8fEV
GLKvCx03R3U9GGuTpBioRilL4kVR0xEHYqIyckfFOzdFxtA0ckUTw4/wCh0zFIaH
pmV8bzSs81W/QU2F5o8qj2HOxGnVFWvgQS7Fxx90aMPf9j6O/02CZ/5HYtENLM7M
gevY15Bl05CbXY1wAUc7Skg1HCqOULvCaunSkaOHqCGdVlMhF3eDEwYLnaCOgjzh
KOU+tAIQdKN6AuOPO6CiWxpPDSoFV1FFyf6fGcnJ9RUzQsQoMy75qgfkmjYcQE2Z
zY6zxOqyblSFgP8ugRlJkrpmzOnuIAcKfEi58ujVJHL9uLuwRpBXwi3OHA1o3zCz
PQeLZAVCsV6cEaZK0a2gvs/WShLmRqqMNwTB/g8YjlAlBLl/kl9noyG9dIPmsjvc
nzkhNaUd2egvPLSEbOPWzUxqH2enaP71yFJXGlQ+WFmdCPYQNY9OFfbAKEAZemh2
ltTcguJ7pILQNnN6AV1Wu/xqVam5MreGKAIqewnipVbz5vypr34CrEI70vxwPJMw
nUDgZJK+rIM9hJVHsizxACvh4gMpQAnKYCFUjqs2Cn5WiBHY/AthaZf43TtN0+OD
NMxeKD70iYk/ScDVJpnspYQ+JZXLfaZ58YhcxeCSaTEwfz/hFSos6W4E8biCwrmO
wOIq4EA8hWzTHaL96mqq79vs4JGKDWAJXC5RRStVW64TQCwU6jzX3rsa9+Co73yN
r0Vvg58gr1A1iMnZ2o328sOdnVQGz9U46XrXN40mAQ4J/wL9wgAaIf6sejCMnKvj
+h6/8FD+BZIdkgk4G2vRA0yqqFMvv/0ozWeoMp8jC05+qHbObbGJNYnUmsEXLtSK
qk+AehvLFSXaLCZlzF6HKsKgliEdEhwouFH7jM7uNB2970yADzp63LSSqiPr06m6
zQ8ShF/PTy+Tz2ydMt2gxoy+V98v+q0yu/rYJkoo5OpxI80bvjGfZlpR7A+tprTA
LRMDIKGQg9C8eahuwVeQnqI+lqgrBz7KghiSvWl5oXEPTBlbbjCDNiVHsT6jbgGM
YtUEAfMg5NG/E6yLymarP8Eac5mBPqbzrDZglt1QGhU5ZK2roL3VbyUoXNOQbKv7
xDXrM2hqiBm6qiFks3gXUAzalE1ITer78BsdX4hnunYxVVmXCzN+JChn0n55vVTj
eR8Va4MwyT4qIDhwuD/UKBgNX1OT8R0m19c5pQGYfLhfeSNJOFXQrxW0ZminffbH
Xn2CjHvCcPqKYIUjkykdVxtdN0tza/miKZ/3YnUiAw9ucVmisydn7FQ7rJG2Av2i
M/9oPJ3jzdeMmioI3jLbNl4/L1RKz77Ts8IOLg5tTwG7lP2V3yjZfB87G+wXS8Jo
ICAGvHBFN396HPtjbZIbgj/FpLAG67Dzd6hF4OY/IXIVvpKXYQb0QEOYuTDDj1S5
l40kf5I2P5ZW7WwfiuR8NLQ+4jd2fvXCDeMKFOk1P5Ty6FySa8ebAmYFNfIPO4i0
I/9xPeAJOm8volfZvupeVhPYCr0DwKn96z/c0agF6T+h+UAUu4UYHMKNaGuZdONc
8Ezuen92aAJdmXo3yz2rzOlVlHtoAOWtIlBmSqiwXPzOYWtRjtXfUa5BFi3Z0N/S
A0yVoXytnqVGAVOi9jBW6BA4E2oCbUyacaLSIgZmKkyi19TEXlwQpY+k1ufh8Avs
7JhHWIB6ECR3Gm1gBmn/SLKSrIOWdh1HIKpAXZhHdhh61aN+A10/Ja5Ogxr82rKQ
rjtXZ3/rwO5Kab6kHbKm1cxAIafsPQdABAiVmLYG4o128ulTLq8Vmls/xhnZlmP3
k3ddu57SJaY5fLjQySMUjx+7BiVk7s4y1w2nccwOrx61vQC+NgFaa/3dScqILEwT
P7XjZRUJQr00PXnX4zGOi1HDQq8ESDatg9pZEmQr6NlNbWm85tvFkB78wmNLb951
3jKapK8keNIlLE0CXVsWEbu15VzEYKBog0eW0hgvGIAjOOQwTDuCEFTGSuGS4I9+
PhLMzPE4Yzq44MhrG/ikE9S2ASYSZKVzFKa+Adaq3D70ykU+YGjjrwbuJGZKkCR9
2GXY65r2OffCoLFfi03Ux+R/5vzvuBjamfblY1T9uVeET/jrGwGn3lCMPaKYEM15
il4AEO0+EWqMaQ3cgZFgsRXHkSQ49VujTsQ3zGRWtyqjAvppXw9+v9RKxMhraxfm
R2iKpHpjjTU4BBZB7x3SqkDbf/r68OD6Ohs7fTs5QgfAscOlushbZSrzSuWpFzeE
orUw2+/3p/I5jxj9QiMFamVOqROouxvn4OS9E5JmSPZ7yviRtI2KnD1LlnVPwX7U
Vts4KPJuC/usVvipB3yskmQHRdL+nDm2qqQgPs0x3v76gsa/G8kzNaPOzibQeg9i
FGGSFx+HdtEw2PRzqyh2alOJxTz97TS7kmlVfzy3RVRYwX8IALbgj0YETIOpkypb
x7u2rsAqcze4Lnuu7w+mzY+HpplBPB7DUjZbt/i8sYEQB56aM54nlrvRTiKZVm+I
z8Y2JfrkPvOFlyspKKAfM6c/p66DYWYmZkAPErdVKnDz9oSABrHUkreLrdTunr1j
F+V5kryQHG4Jtu95smwcdMdDdmgBbMUS5UbTREQqes/oBTvu4QftKIgsNZBNt/Vq
YpxWZvkaL0UOyWNrz1kMvcKg3cwSJ3qRTL9BzNLKakRbAtnAbvDbK4c6kAzV75Dp
pmYHbRTAmgjhWV/5LAQasglssme/LRddo5goOkDfUOy82XSp+7OZUV32a2GbswYT
INEeFo/phrB9GFryuOMwbutjlQEI8JdTUHArFEAB11+2+IaW8EdYpPUUqaJ1qVCX
nHr9XodBR0TTPvdZ/1u0lyxTT6nR0QPKU9cRS5OA6lobvFbvmiiScwA7qizJnR7q
+XLUJv5D0YEhpk4CjI1q8pK+eQRW4w2gwDBMkgeCwUb3uRsOA/VATwCOB/uw1nFk
7EYa4nm1DZc+695aj7tPwZTlcReVH12/LTsuNWlrjvtvDTp+kiIj/dQFJDo/s0/7
PeTn5Bp9hAelCw+VWvTSVyRGXVSFJc8Ml9iPTAAyY2OPXLP7zwcQNFZ9q5O5w75C
Csa5ZzrIfARxFTX2cndtXXIrySzDYj+BauKaRXLT/dFMaYW5J/3S+G9bcKLAECMR
0xPGvtktekDiXkIXhcPaqxdEqlp4+iogBmoCane7fNhjDtuNA4o5qpu+6bdoAR2+
0F2/gih+2+d7VK7PqPINkCsrig5dCk1kUxLN/qzUqsM+hzVHqca+Rz3MBKXInyEG
Arodn7vi2SNQvv+RfR8J/JAuULKEaxpvQdOOgzUvIuAiSAethd5NlBUQnCneIFxN
28W4iBc4B1C+U7RAb9aqe1OrgVU6gGxRt9i+7BA6FwT7B4mj9RInWT/mfWlJfzlw
eIt7OgReccgIVDrN7fNUw7T6o+W1eUD4nf8OFiynnXJ/z9PEvBMTny9P3v++VxzV
FzMfpaiLaK3ydWJ/1H2cIRE+0NojZfW1TcvG/qcyNj6uYGXHqhnfJZQ3RZPIrZmf
PNf3MCuRi8kZozwhZVw0NbyKnBFne8AOUmI74xlRJrwA1wO+hExPrC3HQAsix1Rs
qBpu8KR4OLHnuc6cQNqAHJ2e8s1Uj4uB3uETCVFOCgAOingPdsdAGGuTImn+j5Cs
cPzhSATeLYyNHSf7+HUn7k1An2eSbsIevAyaF6/GH5DytoFrZhUSEIYGrSBgH5YY
EDFQ0cCBfmFnv3s+b4wmqivGrefyfkpr73U7M3jOI9wRVLUeUnPWzfSuGQ72Tvoa
SmFLgtmjBhvTp1cZXzzKuNIoFipKbtWmjVYPoKVbqW5uNsG/Xo8z9JktTunY2WI5
nxA8d5CdlGgDC8SQOXjk++3TZ7f0NiE9m+aRRRn5vShFzYPVSrrJdSvZaOAXsNFa
B7Mp0scQY6cBHXE/imidCPmK+hF/oYQE1qwyVrUWWJpihNmW6ez4rYxujaacMdBM
VrB32CvrYKRZeiCx6AzX9nhOGkeC6dU3fnpvgPqb/o2SCTCyNF6PIz9k7ofLPVUY
3p6GydaYye4LQiwIF8eU+0b3RYduGp60+MwkpMZuL0gqcaf2SylQOrBYF5xjhIFA
D2rPGl+kNNB3l2WKbF5o7ohIyr5rdpxbj7CMp+6zs7tREvX/0ijc993VQzFZ+hTZ
KGGxKV5+Uu7V1QgIWfEad90Jifj1IQfL03VgJMoU3M25TFct4UDRc/YiyUJQNHhK
J7Txzf4hB+RWUb/CCA+9CcFfjJxZ+oOHBirzslQq6V+2nvEz//ptMbXD4VUNKRr2
XRdpO8nXzPBeh0H0VJ2N/JH+OU74MasyoDDGMFbUEjRHLetnZYwchchNrzUSpIAr
JVrl9T3ZnG2Ev5yB6BRNpTGLmIeplA8mQz9XFlKln0CL3v2U0b5Y7+gYqkt3ZJ3/
rV10c6pw9G19br7ytl1DyF2BqH9oAS6K9mS+pQJU97XGZc+8GLtksr83ZeAtwOuk
GAUQYhrn+9z701GJSOWNHa2Go9DU+aAPFaEySwFFyWwrCR3dV6BKRDaiSJp6LHhJ
zy+s3P72Mh668FtPixkI/NKOAbSNbxzNQDimLbPZVu6OadmEhAU6wOWEUwc9LUJ4
alYIlGnzbTDDOKpqiXEGcAQtxnX8O1ySarTB2hRUm71u/kKuqYY+Z27J+QO4+jVb
FccjmHk5Iku6hVcSLdr74faL8jNscsfqSZtBJqZYLUGQpj4EIicHbqZtSpSqpu1J
6Fhey96UwbmFgBTSx3vg3vbJpe7OoNqEUpEZVSw+peXAp8v0R5BrcfvbwLu9MjNB
+2lu9VLy8gubPU6u3Feua2suA5Yqi+rjQsDvQnI1FCzXIfLUImA13HEhsKCxtUQj
Dx5lj68DCMXHn/A0hSZcP/9Y8Gv4kf2F6g6opKe2dsg7b12r0ih9sVPXKx8KzYX0
z2Gs7g64Pi4s+1edWznYVF7e1tPxqDK6pFOzGqTltmQnZmwddAaptUohWqdVCBJP
/Ei9tF/zdFXM+7zVMEzgvZhL+qdngnd8joczwWjt3TQyiSscC6ZHvblXUxYqspzZ
0MoCdi1S7rtvVoHN9UKuoNOxwWCLZkQXSh9StZ4u5QF68F55uyfq65ep0P9l25Nx
SQ+/wH9J+k2NxO4LPfzebMGkIU+tB7fJVaN+L+wo1/MLVYiCw+eVBZgZl/aFXayV
4131gPoJZo1qix2Xw+6Lz5iBGoCh16Z7+IZZgWE+Radn0hL5/bqA3+JhK6keRl3O
ln+65b5VHyxk+KqnvU2LDNFxqLDKNSf9ZSphRK7fuzKYak4nIUrnQvqys8Q1TWet
SXa/KeDQF9LxMFJWB8QHMpQpPQ0bTcliQyQLNuguaJugUSTqdUYpGYmjNxXzGaxx
v+6S5WAuI17fB+hT6GO7kuvSK2jKNfaCCODm+M9ueQV2CG99AxEJlF3gXs+RUXR4
2EE9/Cp7SI5fSAKM5BuLVYUJYOazwsQ/s8bBC78ayyzLFLS2dc661xrRgpzjjKVR
ap4Fo3y3PXBOWfBtnF1Zr7kQQQcW8Q2+bhyMO25XlkdGY8jmI/rpy7ysWdxk6mNV
W+3ZFN3Gm8F6eGY2oIsZJIvOygfQXFqXf9BRvJDfZnYObr1nnDse6NHIrXqn0f7E
wurnT4p6uolVyTVmYMF0xeaqrQgOaKiPUZHQVMKPjyVGy4+0F46VMmAoh5U5r1O8
zToC8gydLXEs2Ruf7RcGisXxtGLQu3UXFTtxSnrkoTAYT8wsMmNfKte7eQ1pLXPE
kri8oIk04A07uEBG1+YG8bPp3ZxArAUeW/qoSfhLq7HIHwIvikXhOe3PJ1hrlG+q
mvjCwXs7MiNl4ba+ZpzuPUuPBwLihQE65qvMiIK/bKEL0LOmK6u5V2vPwGzDm1ue
F6tBq7DNbWoqB4dAqT21t3c7EFaXpa7g3qRw64hyMa7FAGL2HvheWEn/myQ1ENgB
J5SG1zJ6jmGVxEpHZJb4z0/MMamVAyMdH2bNWYB2Vnb+VknH/8velpKqUEwAmf3Z
eGiJ6CXBRjxRfNcAasLFtJVHX/nvUhNqTJcJxPVWb5hBL0wfF6Ec2xLFaiJGvJBD
qowIiuulgnRwr3uvEMOSuGQ3jNiYnpFgUcUoXkkrQQggV81+LUQIFjhb+xV9DYNB
WRH+XL7TFLKJS6Fk4PjeecUs9kLk/NNnf40fU2oCJCw1/zMHMKgOQEeFesObbyfu
6cFedJxM8AUHfnQQB4++w65B7NPHhSdqws9l1bMcHcOFt6bUIooTA0LzwThyX1x8
0QJXnm0936dlT83aZfJ2oILjEvMEqGpJ46V80Wb0VSdq5vEvsc50XmTPlHlV9UrM
nLpFyt4J/JHcAbeka0vtYHEfcLJvLDMYxmuD5MfVCRZLnvZ/vZooMEl00ElPVEZ5
vCsjrHp6gRAxYlPy0gT/dZBvYw2nAhSgxCAi8fvgPPBcuanpdvKvukXvddkr9Vdq
YcxmmChtn/rHXeYy5YJjP9O6LaEQTPnNBsXREeY5euFjlH2iStuPDipm+HXwx+QL
qgOP6wCV8NckP7I3mybiOqVLaisptTLNkmX5N/g9oUzPNI+bRm4N0MEV1apaZbH+
7gUgxrBk1oh29jxEYanZDKnJDkoEbRII4VeSQxB+nGkp5LAiDZXI4zs+XniNMTNv
G4dt/qGfMb2kaJ1KYr6Alx26MBjrHhiCB2VnD/SmWKba1c8sAqwvB/KmpVZtuGlv
P5PxCBP7lvePuyQ8dHmxAhxRSMWG2x/dsc7afksCT2cAGHyqD5xpSKbYTOgFzKWJ
MA4veGiGwXiFkG/eQnIO+0EBoqZR110Ym+wZFATgoYyLPhR4xMYOnzs5pXEK2xg7
px1W/8asGuBT6D3WbqTk6KjaMxOHLyb3geYK3AwI8YIP4AHoQhtNtLz5GMW+t4tz
k56rmDBHUhqwu3ls4DVbQbQWbAieusGpozo5plrEY4Xb0W7pdQzAcUGRbX1sEXbB
TdaQqJiWcKpRFDgllVxezF4cuOmFwT0p4q6RpzFxGsHdBIj3NWC4GsCpySoHLSFH
ICjLNis8PZ/h5KadXM8FSdEuYsrif6FoyaiZcPyagcWznJ1CzGWUqeCn4Yq4JOgI
3REozQ28BWmIIzlIpltt0xKZuCBife6++97Fc7OVB7ckw13ZK/VKSxsvnEtjMJbo
7Mwup9k4/SMEfx63LwFN4DpBVG5PoCb6P4KlpI7UjwI85sukysX/XaFP7cAfmuAw
lpaNbNxhxBKYvjvhS0ueBZuxm+GNDDVw1BFU1BTLvlbcmsXZ81JrRqqCH+fJIdJU
u9LddYP7gx9S2AKbKsEkT+X0kA7OoiOkFRiMDR0uT5cOY2YfqF2q4lzyBCPndxM2
OIltWUT9I7xdFrL7ex3SqSW1aUJwCUZLU5K0CVbs0PXjM/wPJpB2DFZmA92y8qjy
68kn6du3hdYz9mrWvL2vtvIC8hrlLBuW5iMl80WNXReQ0A+k2Gu3sX/oa8m2QLLp
ikxMRxAqx2KdZg/8kxw5ekIHHQebDXJLSLWJBTY3Btuxnq8pSu99RnAlm+0E8sId
gHUV2G6QvKx8MI2webpVM8LHnRUEPW1FjNkYlFDOIg90XkGgDgi2SZVMJgoNMLj5
gBR0SNr/PN5RHVUkmYsYzIk3NPRpb5LjDdIfcbhuQMFk9YMPKH1rykFbo3aph6et
Ng288SE9jb1BcZVydaVbrSsYOwub36Yv4xlD83VLO7YH0E6COghrYBBt04Dgbac5
ljxHhDodcXYQq3i8Wb4KnZ8Ro2rrn+B4mSAnyE8zeQzge4J3ErjobKE7a1J9OEyd
4vgWZiGjsbtPvJ/8Y6aHnQPbt8rTV6FID+Hxpn9tqocpa1dM/xj5szOz9k/Deb5u
n6nnI9lgzV68x5mDBlzxCIV/GPwcy4ygYxlcy3Lmu8T2k1rI6M5jVKXNVKke/ssa
DDB9bRh0SM0afgGs30s3YHdlZbPR5nDlzCsZ7rxDnvtmIud7hyoi76N2BKBRj8Qh
VJoMo7jhdGdybngpfUbC2y6UW7jo22ZsHmSmbtXHPa2eX5f0QdJ0GUV1vYPeKzIf
S4Y+Q5C0oRQNAC1rAz+6059PgHEWDR69EW8W+BRtBNpHd+5UsZ7PFnAUsClOBWfM
ZVvG+qsTn616c2gsXXh1ZuxYFGYesG2mw0upodAMPu4wpOFFnSBTvwyHrni0iZAx
nAtA414V4cJTBCRbBZrqMJnbvMqB7SnrBXhAbn/1dL/T7vsM/terygkvvAgtg0g/
40LX+w8mdbm2sLysLUpSMXfTcNOjWptQZWLervL0LF595TmJ0oWqdruvG8SjSWB6
SuuJ15g8qcDTIFOuvzr9hCLJHNBYovGQEmNzejp6jUCar7PC1ZS6lehGyl9c+Y3I
K8x/6IUlnYM1zlcZ++Sfgqz7PjYmBri/Bw3TZS5hmkq231FdlODk2ZHTUEjzXDgf
VDHempE2bkPUdsfc/xVR5YzTosPRoo906aqSrsg37mI3Z3JrEapzdYpv56cJGohv
Gergvdfxc8QQ+rLQUkC4Q3Lszr4QWphper0mQen8RBel8fyRCyFt2wvvHO6iYR52
FtqOc66KkcOKcVF6OK5dPiGioI8eEvizKNDalOroIH59mMBaCBKiwokMScfpP7xp
131kCRq868DUKtRdQUnKaAFGdxfS51ykhY/ed7ZNpZSXBCBxouyN7pxQzflesIaZ
k2Jaho0c84nO7BrrJR4Iw6nPIXAl11GZ+ZyIxFcTJ6GdCTz2JABPXxdGubMS8swJ
6t5tQ7oj2rxfLdi+5wpEhs9iB5T3/iRUDDJcHKdnb6Dj0Jjqbr4MdS+FvmeXnjSW
Jk7llVMaMEFd/dF0YlZaKjDE9G19X65VndQHGE8dBWagk7DRo0UAbnpsbcM3tm3K
JpIvRmNFVlRVCsKLJj0BRxQWW/STFEcRxXng78lRfvhzTP4KxISf0F+3nBlUIUrw
MWWC41mYEba7Ee1sWcixxA7aY9Oe8Uq3XVynl2nBCWB61l1zVafLl9gPIEDEOvXf
ZvZJu1GBJlkSEDO+3RrwPmlMabMNqKGW18mqWdvVer16OqgKYvvTsL560SHsAAU8
Pgl/ghapfnxMHMV/aATYORuBzKry368+E42raxXFYe9/mnM27mTeF3AIRIoVvKlO
AtavDD6zhkFpxG5B4lAWNq636jNhWYwMT1BhDLPD8RF09HHCYb3Fk1JcWexcy9Yr
k9zDUnKQJBbsbiBX0WEN3S2NTX1/Hlu21zkQOdkwIYXtHSNhv59VJGbELUOxrFMQ
Rx4A2gdU5oqNvSNyR52apKQiQao4TCohX14wGS7LGRzqa6XYkmEowrDhoOeaNUMs
x1Nbj5dzCvhW3a89ALwOiERaT5gU4nh4gHPpFrwgA+XGxGHd9dBsnbfviL5UjMwy
W3czLvqakvuToYnpLt6eAnzcYNx2ieLaC68zCFzKVpM6dIR7XwZcuRwg3DWKLB8M
OffC+P88xXlbbM6ufc9rvTiAuRu6fSHO4hhVQ3XWrkwcnTabhs7iJ801V63alwms
DvHzktV+CYKG1H4dPDmmxnChnUGvmf8keMFF86oZq26As3n+Ert8+ArWVjKnjDmA
5jVdRETS1Z52iYAcX8qJ0qJeiVao7mSHozZvmOGQrqPtl31IWbe86oChvEXe24Hx
cExDnjf4zQM2pKXvLOYQBX/n2Rby9MJu7Hq/pt08Tq6gz8sfkU3shDuPozOW1p3m
eULCJahhOdZBYjZWikeTSPjYgPYCCzeppuEYW578BVULRc7E8+n0e7Lb6jt7aJlV
0dCiLimqg6JGp6wyz4+L3Iya/KdSTmHlVEzVJo7dEfaPKB8cTsJlbFQksGzcp0/l
5w3pKOrHmNACBpKx10UeMuMWkGDLkBsDMO9DIu4+vQu2GoynXJwwZjLWvIg9MwYI
M1oFSdDZgAsdd0cdJrh7piH3ErhCb/MsHnvTS55RbFqbjh5YvtJc3B1Tq3Nch8BN
vZKUsl1vWT5eukJwhuuu33NSE9cmGF45GmkuI67uHDXQhP//b2tgl1Nloz23e7G7
E0kPSqqP6C2uPKrgtsq/j+MW7NFONcTUyalFeyul+fC5ft0iZvRzendENDZMJsLX
/wekhGpQzI2uQMlbUyeaDZ7Bbc5rhxivwoRA/06iNEP25tUciGSdtUJulEnlVspp
eHsgRISVc8U4ly70T45/Ovscc6djW+BfYnp3mjJDul33eaGheSJN23+Asn4LnNDD
KU8vvGHmv4/8rAUStQeHwFXXq8Lsr8ft+5o0LOlQXDkADi424gvPTOPOlPOXUEWx
zQBf5n+jNNGw8/lqIt3KBGEh4muEnB3NoU2yCIPknKFUfHW5J//etx0Batksx6NS
egC6yxEANcmQGQaiEF4S2UL3DN0ahKeNXu5/0RS5O1PExwxlwotoi+06h1DvOyOa
3NNDCpOInrmsXVVyx8CIAa8RckHQ8hndV+b8nvcLfKjrFVQWfCDJGsLJd5cOwOhq
CUnCT+5rAAJQ9In1IdDLBjG5pYuafShNrN3cO/96utbfAGnawVZNp2crCRRZBkkj
s3/SDbfsOod/aPKIoDXTZ5KQ/AIszNWAQJBq8+CYz+3surHpSGQTtrTq22CYO2Zh
0SBX1lVCmuk2dkTHks6T/GNCUaDyQPKp9F6LyuJlV+ZMdIK5+pVRtaBGp7JDsIXA
nIsT8/1R4RF1OeiVz3a6VBMI+wDppmqqZ0MeFQmDtSJa7K24QDuRcFDXCVLFbPcX
Nftlr9l0jfg/tQFlSuLQ5QaDhFgouLwqp2Eu5lVPfUJcUb5ZTRibnpKxNP1AGSNa
lqYtzGjF7BJ+9kWV11i6DhaFzk5lHnwADnQ0c9KB6s4puZailQe2avc+OBxa/Ygp
i23FkFYD45TudMZTFED3bwR94ffWHpu1J5XLnTQp2QRfr1J0CKMJ3rYZUH98waUq
4O/52StblM6invBjWgejtWIPiXjB4QrvQ48FOAgTO9tMc+VSivd1EhhXaLKzwpQ3
IR7KZY3iPdNFOXQHTzWMs+6i9XrBdn6rS88ifMEPp95eWAEFVOSmP/gLQdAncrfp
rgtK6dyONr7eHrdBYgY6tYKYUcbYQJwu+LrlI5jCG61QVeyB0JTx8efiqXZ813bt
lxCHyJvbJelVjEwirwqbM+zvwrzgKCkN8wAIoAidqhHP67ErTomRMhUbxJx9PZw4
H/h/sXS28uHFPqcjcyi+drq9Ks6ARnkLiK27DwTSgyFzEy0nd0D/OkbJlg0Olst3
yfPkWP/Z+8Viv5Std+AS9S73WjlyRfAPrs5/uoDjC5Nm+BAjdZRbBzX4z3+Y6Bko
BPzaZi/d9VQnAV+AEn2sD0aN5TMWUVbzzqVont5K704aePGL7CneUB5/p855XikH
ZzC0gaRXCsZT3ahQPSaE85mXftfegkiPEyQoZQJgsHOLKSjuNH3jEDnVmSRY43Nq
7hg/CGGqRu3kD5dRGmUYRvdyaLiQMEuoCbD6QrYIX517ER43BjKVcuJcvJztbkF3
U1Zpm/oOH5T/ip6I73Im/qPh1RNAyDvE40hPYrssVWUO2OAOUa+ecmYXGom8CSwQ
Pf9wGK2de9cd5+A4LkKix5enHWHaLr39a4EXR5/usR2g6wTgsOUnN6uQEyYdba9o
Cm/9PB90sR4+h7HIuRQcJhe1+F3kNHyqQmepP5qG9xlFeafEsgoQLEnERZW4txvf
i9eRDKRl0vzUIT4BPRJH1gSlyuESuS7drZlFuy7iA7KB+8sIaF/oa/oWniH8v6IQ
+pFgNVWy5gjOCppyAK2n2+tlL2EVXCHl16PQ/t/UYIiJdDTZT5REDwYShNU++gIx
f6UalMDBn6Senl0LWmscu43elGod9MYj6zjtmSQyg+vJniit2Hwb3A/RFT6dy4kr
idD7NibhtzSTAR/sAhTiDD1oiBVci0Hgt5vB6tJkhBjR+io2ZsSKS89HIUpgmKJt
umXiJoEFl6KegDMpvpCDB/mpPFeqy0tGVhPBZKNamINNyLPGdRPPvn/nWlwE9AN7
H35kXV9QdjcTvopJMDYe3zhux/UtLw/NLkJ4R3om2Nc3ZLmhTU+JSZo9ocSsT60e
9vz0e7btYJIWo4/wIT7W7GLxkp0Npz6HvF7109arot36cQINL6Xta1JpIsrhQfw5
DnbcAkEXztsicB2t34hRJJcot0Ef0CMFdVaH/X0w1Dnh8bxXudtzjACS2zFRggFH
HaVUknmzJ3bP8sGPZ1C5jXWmCTWUAvhGJ0Bm/8RC3WkNZ57GUV7/qZ1W6CpCV141
Xmw8fKoSaCgr9GU5CAMIz7YnalMbKKTHB0WVLBPgCEi4lyXZolYwrbSoXYB3uXG3
dH8xUBZ8FtY1CSXsEvOLYETUUlRJwHjM0lxM4Ul8YS0NFxvmF/qGAD4tYEJz3QKQ
qsreEvzGQ0oHrGD3n1DqsLEDdbXboVvdBkOKl+j3d0FylsaXIrHsgv+Y6T4PAMa+
xiorGXxHHxnnzSqRIaUD3nZEj0fj9J4BeX1EQG63vXMW3CzXArhcKnt5DCWkTil3
xF6NDUYpzYsASfKc+9TxWpsJ9hghITvmsUYWdlpOE2LPK5+bYgqGpV+kzuX41s1N
eVGQzVBQLV0UnrEGO55UP6RxRJJiFgaxz/Lx+51B4xomvbyjsvg90YMZns9e7Fys
V1oBJ61sOWnae9K3m+Z9YFcZJrvuK5HwXEUCmyJ2sY4io/SUj5Z4+ZhDEoqpf0/8
Kegg0q/vUhChP/CjpUR4/eUufYwg/vJmU4Dun9h7j4myQhfEV1NtPz/ihU+wkLln
0BPvNiRaxptqspMhpl8KrnKoqvgQCeEX9IM4uzJGY+S2hGvw8rt7B+JojnSxF0I6
7nXqk3qxsu2sow0CrbqH46RcRlmSk8ofEJSpEYyMSICFNX0pcc9Itc1EeNh5stDs
NiWfw8ePnYSoe2zoyE0TO8N/JTklWmlUx9xd1XB+POUZrev4YF+tkeP9KYHlajGl
p8qXMHQcbKKQCM0Y9KKFIw7MH8RkqkFxNsFYdgP0s5l+SZX8+a+pWF80kjjAI9ke
vCpYOdiN+l2g7yOXYTLGOeYTv0hJnKE2LnQptBn9b8eRgmauNULXvUqXTiKqdjck
nHG2dm9u88lXSXIyll2dIAaqDR22L3szOhzMzThZYNOFITShvhI9vs6kedumxrYo
2coxO3YW21I/IG++AuXaDxsT3HMgbx9WnLTRYiakDtjpHrs0aBJJAYYQdkRl1juD
Wl2vOigtz5lbVpD64JbRNUWsZL4tnuLbumilDX+pWmm9BrYe9CMuokfNWQkPZ20P
0XopZTkMz6g0jUfVVtimAGPGwYi9D1QiMGpQWY5iEGk9Rg0qxCmumfWVCXHipSGP
BgTBAO3H5+wwOxO1PV8Zl06aZFSRAAkBziIQU7Fln9EgUVHbUvZJnJEpGLeFrXh7
I/7nSSCT5kcxtSepPRfSe5nIqt7tE8FgCCiKdaoMLk5VyL8aS03FJWZOMj581TdI
u7YWcyzPuzWZDuti8178WrblNX1cz2HKpRG1s3T6Ff99J1iQBFk6gPTgcWygRIDf
bvf5oxliTO8HMFuQYFytoSVw2jvMrTwPz+i1QDYQaXbZ7+1QRw5TFtbPAy7dBWI/
hPIimMB3PwFOXsj955eal5tU+1ZejksKo9MTRv/oPDbctU0YY6JITfI7I6yhoagG
pLHh8/YZy4kjpZ232ilgdSrlGvKHFG5m2Lfz9ffsk3Tg86k+qVlqZvU93lo2dKdZ
jmyxhHCsZ7R05taX3SakMK8idXi3yvxiUf9zcP+xcnmfBzBD+1+SI91Fi2yvSLMX
U3vjKt4QjzQw4XwAFyxXSPkiXPTmYQBFlK3dKUTifd/AgGoQtTnB/ut6tRIvHKme
NrIgDukHOj4ADce3iIVuTW+Ru+sxgXBv5tBA3NPQjPOc6PFm0WRX9gq/smo9ot85
nxp/o1Ni9Mrz3c6JOHUZGOqedJf/oUv8PNiTWs0KsB34e+ae7BwBR5f9IBRjdlJb
CQiCC2MWCbQMYvSUl5+TfF6Vco66pk2TQOTO4tbX+3twT5GZzDcD5c1MuCCcl+of
CUBTIS5jzg/kPmYVIrbOoqMyLOiEGGe9X/UlzRszO8CN3sQSnJjzPZ8Us3qhNnez
4o88Ou4nnDonFIGQlCnHnEJYnVCsrBtjL96JEbDMajpF+MRMtW+mCGMwPFmax0kQ
wo8t8sfRoI8piPdl4ILUWMyq2pbMwZt0czwAgq+8bSo3sR3kYJ2jruNzcIArPyQy
wwUeLozVZDaGsiv4eUk+Z1bpmvub94rOyAmTq5Q6a/t/a3ttMy0BnSQQkr62DgTd
tLfTRxDqHVpJtI5mZFQKlz7FguotvI8Cm4PGOEZhTk1bMsXaL5Sm+VwaGfz3JZUZ
jkPv12bjC6cq1bi2dCcP2A+U2z2pEapduEJ8tmEG7moWoF9ScGZhd6lpIzjTLAHC
yFsdx0kk3tSQeX4aMUXLIjH/2qXCy9uTEqBHGc8sdUtowTL2QJX3arZB+8ia9XjS
54LwnfbbB+I90ROFONA4cLN6tuBzV0w7gfL88AHJeYMUY4dagSOUenurIMHDJP0J
qaICl0CHzaicxtM2tmJOMEOhbIjxBCURCe6iqbW9x01QDUkxxarItwdM8FaAjpR8
WtqnOZWKX1Lsgr3ntwyaco1GdAXwHHIeqz+msMf7ym8o3fWFBv1moqcKVOl1CLSi
loIYukklYRkh6xSqHcIFnDvLBiSCOwO1dPSCnUAdWSwiPcalAiLDJjoRa9QQW7Ky
2Jsm8L2dUuBq7ZRX7buJGNCBtpZsjn+J1Xh2N0dErpfWl90aT4+IwOQdNWIFNZXe
AOT0R33g66my49uFq7OEV5xh4nFzwxKHnivOBZ1W+QmlBFSqbvWv3T6IVFZUNLlj
FDsKvZPtSoqLHPtvQ3ruvkeGdAEg0qfQbMPtPBz4Unvuq/jufzMbfm9MCODbOevL
Wlgmv/wwUMp3t0uo68sZWJOZk7y6RAmKQtkZFfjbIrJhGFEh97nt4DCqhYh5O+of
f2VJ0xL19PYg9f7ziwA8GD0f6jXQO+NMSwyJiN0heASgEtxufCDV4Qov8+EntIp4
C7Ffh2CI8WHCVqrxfosESISB5jOvxc7PNzI+8VCUpl8b2Zw4TjNkycA9zWjAQRg3
IyEM70VQJYe8iQBdsxnNLJChfjnnxubkvWaRYlhOzGZuxUzRg0/c+xGqOgvR+QKl
2dSRl1eEWCHzZ10m4bQuCbAAiXNo27NzyFgBboIWm4QtHoCEGV15h6UX4x+tN+8S
cVSWTqrX1/ZkvHL2jM/oh+NsWFuyFtXBvUiesB5LvgTrcbwgh6iZbbEuhcRuQDYX
CvI1b7QroaRcusSPEYCJDV0T+WW8REAxZvvt4bLv6ZW9jpex9JUn3jmIOv75CAO4
1WVoX96LlG2FKniUXtoojKzHI3p40jowZiOH9LRuPfwp62/o8ADFZC+IR1HnbdIG
I9ecEtoBZy8HxqIgruSpwnEtk4xvV8G3P2cAex97Ef9HDEKHIP+SCqyIRKevCcRd
RYUrvMBCm8DIKUoYrH2q1JUIGZ6z/oTpPxL+klVZe6+DV9MEZA2fhbXLfGJueBuG
8qsI0C8Od1V7LfOHgURaQdJBC0kSk4DzpjBiRzwEe6m7oP2CY08K8fwJpf/E7/aQ
TGhZUiK/9KLs6ZYUy5FJsclIns6QfBYgQEx6KwxZZG3gk8VSa4Y2yfLVst2JI+AA
FwsYIIxFaaieyTR0IOB+nsKcvBUS73zybedMx5gBVrJij5tFNuBhpHK5ci3wfZKN
t/O0D73R75AnlNkyYGhAMS5XaC+TBWGuCdMkHpfmzEfvo6aa+AfPcif4bETi/h0A
inZZbHr8ROzyEPIwn6Zf7bT/CayPamu4IgA3yWjjl9SbT/yxIaLrR2FMMewRDmk8
01irHcch4yIIRMKjfyDkQihLiJdFV58B2u2TykcZ87DqtLdNK0ZV7RHY0DOflIa+
Uq4y2kBCd5Rv2+p2H0Gi83gBst522hvLqXi1NceucdQ/AlR6YkC+ua8d4gwozPMm
ajLbk3pHQTjM62kJoRKqsMQuZiPenULPCYjlyj6AMVqVEadYhnqKyHhwchHTN15A
chC8nMRlJiN1Zy5M1ez/35OaG7ZobXcyXn9OTHzlwn+bXSzQHK4IcreT7P3PPXjq
e7XNOIZYm8hvfdP15EPdcFMhSvCJ+XKk+4dx90hJzP03909cm8h+PnpOfiWKmZ1v
pco1WXdaWvoWOZ5PDdWKsuLfJ5Kw4FFNQ073o4DruUaBDV1BPmXV/Wjq4+aoYxg4
nH8TEBKdNn5eeG094NSlasB89+Oq0fQjKewZAnCsHbR7+g2+V8lSrisNLx1fbU8Y
c4toZl3/5X/lGFtt8u2NLY+fLISiygTnF85qifa3SHlnWabXZNfS5yn5uZpu0Qn8
Wh9Q7KwnfEDKKnpnRXI/mGMRe4r5Y5maIxefNWGOWY28yGGcj5DomGN7uILxB8Bw
yL4Qy5O5Oxp4kJYwpILe8UBKfGvQGuzDgzeCN1VpWgr94lqTsG4sRPxBIadrYr0m
Vw10juYr9/deja7MFxrFtM5aCwFO/nBiZyrBnEVVo8MAjB5QLidja31Q4mHBp0eC
/CHvH/QAgnRRl2qAnqc0CPTm4dcg96Tua6T4XHwuCAku0BuMHNVwSo//v+clNseN
JVsO+Y1XXqPYMATjT7RD88QE/V+hRPGzkKKuI88e2iJlzyP+t5zpqurf7MtnwSIA
nEhQco23+im6SOEQ1OCBGdtLSBW9S/1kYcN5hhVx5ItQv76Umin8+FMtY4r8bktp
QZsuxa7cFQlakPOa321O8OIiENxgyalJVaTO4/wdKgWow2Qp/ngyrVhOiZfES/xv
Ao34+m24QnMUcGvX1Ei5RxO/ku9oRjIcP4KffB+1wJi2fHQtc01QrONhxbqOnkqp
e32d1IzzPwpY4EH/HH2D4ENV38qYoJlfBa+i9Sft7rElQnCUGpS9SvCFocvGXG8/
3xe3r3vx1iGmA+bUe1CUyr4p+2ShhtmruVuusephj2BstwWe7dnnbJBa6m64QSz6
6m+GkkEwbxvb8JqSgLYbwZWLquMOWYXntSobPNbnmAAx2mKpPrNZsVGbjCsVBgfa
RXr5LarXSQGtzuLnkHxo9abFP8q9wb3s9uMOe7GdAVUUT6fsFA/AQbJYv6aOXShU
OCTWFO+tJTpitb8T8cB8sEkIcwWm6pk3qcj86hZc9H3W9G3xCWART5KeuEAU6avt
KjZ/02g1cffmJPc2z2G7YrBPEsTKPXaaash4rkwYAcXZwIpeg8HpBSkSzaZDzbtm
3DmNFuGkaI2Gy8iNkjxz1xfgMTOBpw78sIh0rIe7ZZ7Lqy1bfy1xuyOqfJ+m7cNC
CJUBOFyyjp7CCuDMYbJbeYuD/V4ei0Wq/bs/uAiDPJjOvyUfsbKwbFcQXU1SwDdU
ZMnBxcqbaZfqMYZkrBjGn8yDxsJlDWn964DGG+eyGoaKqjZUqTGx4kWYO6csIHEn
qRfrt8KcEK5r0JmnQ4gitOf7Njl2WoQQmDwMoDZSXP289ZLoDSwMvmWNr3CeQpOI
34aViwNKSwq+dOlj2nx/wc7e7k2w5wN0yIvd3v3QP6ep2gDvBbdr1HdfAR4I6DWb
yCNs8F0fIb/ZJonKzh+8h8VtW1/h2WqeFg8dfKdzoAdtjjsXV8sqnj3MAz3xAUVh
lL1FvRXO2LOYbxXd5I2/FBW8Q6hs3re+wGdy8vD2b/+A4mMqA+rN+nuWn1ZxdNNY
4KIM5jw7l/M13CDzVsBr9pt1s1SU4rIY6j/xfjsUexGWq8ocl0e8j3bu3t9BzJ74
GF8PIQXipOHfqVF7V3rTUL6UCWFLhyoJ16oLQHn+GO646BEJw8YkOmPHQDE+ayy4
H5M0CoDc8qwPliJZ72zU8JqmVV9sLAdRMaQ4Bd9cbqAa5xg1JJ5XqkhuVE42cOLV
kcuWJ7JDrkhkrYIYqNTi/LA6rDJz3UCp+OjZwR9TN/tHKw8RH3TybY+rZrrPsluA
OObcotNx1XcYVsJjm9cEg5LuLHEhKVcN8AgbzxKib3j5ovI0/VLqjA09klO7BIol
4cUDg/eu23FR5cM7WvZpcYQ7Sr59JXMFVgdZJ3tQ/gJPQtGZ49PFa/qcWarXe5nX
K22zbivgou8a7feP9oTyNhuirWquTkhzaKFS6xDWjpD+p9c8nKBDNgWtEV7LxNmT
Q2WDHAD5ysC4E+xXEFGFumZTG+vWKF/5/RKpWdeQr+VUFjHs/4Z3h+qRU9dPmkNT
bXQltL3v/sYjTG9M0s/pOa6Ljdg8mkYIq5do6+0Hau4awsOFG6atPBmSXLZ6fyGc
K/hULS+jyQwxg0m2NtV73TESXc0DdpD0JSwcF4bhta1kCZtnmQJYxtSVfK+NgBvu
9iP7AY1382g2wZE5NepTtMp5L+mnA9bXkxGtApOFo5458sG3pDgNOs85YH9XuAve
zZrhpL4bjtYiBOa68pvR5aNFe8QoFAlifLWN2f4zqoglsF8M6lITYQDhdpwvhw0S
InN3ASoSY9EiccGuSRrdsInk0Q6+JJDcrRZfCN91QDAYoegpzEWmx2nVOoAJIwPV
fsZGC/7Ob3uANJ4hwKjxARnx0w+7pbSkeim1vXoNFft66osaPlgJYRlGjwdoR0r8
WZUALfDg1/imZWIJXXukhqwhDE7ttyNUUlm8zppnMEKRFxfw+IPJuGsIQ3Im2aje
DEmnQNrz8EVZNOvySYf2TWCBBb0MT101qk49TPypiDB8gDsvSdVkuQ9PxFs0iMwA
bHFssZ0lSyyOmpbfyEmuHJEJkVEwAo+tZ/FG1LzNj934L+Xi92DIshu+t/kRshe4
0igjpnEwZEZpZ4iT8HQmdpCBFvShDYyRWntNjnBY4Pm3gZ9cctTopyLsupu+Rpsa
J/tUn8i5m7VU1j9R9GrUqXvMMrqQEhLSPVMyVC5vsyp7XMVtOxL98pzut30BGwFH
0bXnY1xIOn3f5LMy++f7Z2krTRJzW3LYVqV3TCfz5JuvQlbhlSDMpVM0/jJDlvU4
CkMqQ+nGNByz/h+ZrnIwHgqIrFs2YWJI9MsLuqqCFTkFsTNoFd2h46jc5mTUTtZg
OaD+Qff+2rbYLxfk5948QxfL0NdGXDrUBrs7hT1OZm4Kbotcw39C8UmiH3QBU+9f
TCbnOeVp4GKdz40hGzBi1Utavk+ds+JCNZc/Bz2BWg+UwWfFyLn4oHLdiypzyRWH
/Phak3Mgx5FEDUE7PPiOROGyrTaDMahjsQgshmeTttLiy3bhQCAlvqTNOFGg2wRo
mauSIMMTkItyYJiXt8bIXS2ugh2S51+dnXcJ5e1OsULu0sFQjvcJ+mV0WOwINCgz
eyxPn5xKdgyzUE+cypWirICOViqTH7TSZ+K/9VXamjACXNmjv/LBOuvaFXCOCIDf
lP4g/tg9nncn1vOrj5Og7tTCZTwf8vqSdc1owvjQmaHcvkryhbzCBvZj8CiIx4qi
qVztIiTojCL6ZCVjf8D/x+uTfFY9xqlR+AhSjqOY1OihBBHwV0y837NgXBw/6zxo
iq4DvsAFIBvWh+m0FWul+LNsvQ182QCURRwbE9qPHHeqsmCSxHVrML9Hdyn1NIQD
rXGN4IuzpOPy7OsneatmX266yqMzM7INodYv85VlemURAIdRiZ7t9Yk6751nTV3M
2dOvcArwblVqDFHkxERpjGkIMwm9jhA9NLJnTRT+LNHkx51Bw5hUvZEO0yEj9lnf
3EcktNGngIwlylcEqgBjBc11RGEC4XtEdFJAWajhOQVEgXZkMj0eI3m/sbaOKZTv
3pZ4qmxnYxZzrzxuTpJ5952Ws4MLs7JESnsFoDxgy/keiEf93TGG5mq4CNrolG1Y
ku1BYLuDH9bNV2gpS6oLOSsI2giynXmNd6Tv6AAleTDKXvnJ8s4Blain5a1Q21ZK
QH0nQ83wt6rGYPQk5v0uGwGqAeN7O2pjLDY3u+cfrAYPsxzwXH3ILgj5T8tK6IUq
WVy0eE1+cazj1yedD33oVv4oJdorr3fDmW/WJ3n4wxJBgtqq7spbfGCfErU9oLzg
iejFkt0hYr4823WN7DQGlulAL7TN5TZX142t/Ga8XYrdWRQ9wW6xQbCACdLmUYPX
citabh86pp7XEs8qTsiR51D6vI8hRlVytfhH4W2+2D8ALDBFifVdwpdWnFq2OPEM
M5sDAfw/wWctBlQafc93laoOSUtOgad260OoKnw0kDQ4K6qGtyh5xXM8vZp/xhtj
7yxP+WiOSIHpD7Phj5spWxnf9JJ8yo5oaV/nBzE9d/b8r2tUdC0wMme2P8CLDgaA
JpXmReaKUV6kBzfb5xhq1XLPqzHPQrCy3/VsW3DWZC+JqZV5ESKyUYbIG0+U6XUi
0XapmkUh2bCxse9STa20dHLlIFev1kuDlW7A67GJgFvDJ/ZereJN0e9cjDUc4F9b
6hR1UewZQ9rCYkbqcHh7HDY9nrTrT5tlr8VvKiskZRSUSSXZUEwKhEnSnmWAgTfo
ahC149467my0GoR24pt0khlivOtvTQgoAeQsh7fwoJwX4Ig8z0+7FUsKmkIkvvWe
eUGRkmqvhVocQv9JaioWem+cLtMzwIhwsizJIKS/euY3LXgaVVBON623/kRIfdwe
F2YooCT1pqrpYSM5ZZfm4ttLQLjMT2dVO2HO7gfKwgt/MSuEKME7lSf3p7IucNt4
YPWzBhSq1jWVKctQRpWXDnvJculWhBaDQ5zYnSmBNz0WYKzkMErXO/MqhAyvgL+X
RE1mKKF5efHK2mMr/BsSP+0ApimE5lDeo1dj9U1OfDKvYbfZkjrQJJ0pe5eurv87
Lha4PHAyD5F8sskxkKgeyDRz+R5Eb+LtG4QRtiNCgVzUiDFG8JiBBA4MeK4T787U
txYKhxloKYvr50jUI++uAZ4vYK2uGh2CLdvJGS64UDVazul5Tou8XRd25s9IiLMM
9TlHKShVETwRE9HiSk9pXyk4u9GKsLAKBOcFDVpiIqiuwOGmZ1Muq2/BKYmrl5I7
vyuYctiKVu2nhsCkTY+0fb0Lv6eFr6KC/Jd1TfvD03z4N2qo27MznpOMSd9aVAZY
qPzfslOtEktUgeWRufgCwrK+bN5CCC/f/pJpHW3Jphs9EfFbL2KVaP5NX33HV8+C
96h72HvqJybS57lA4u/c1LMEJZmGweAyYYHYxx72tskUHyjUhpoIAefj5r+MYtCY
ISfCi5Sm7ukawP/I/mZskQpvkQXGYpl36PFg+SX3Z1AZIO1taiZclu/+bG4AyLwn
HAQ28JVKEgdOyb5cMsrrcBQ4NR3HEXhKcui9WhqVnm8oLerz/y4/WcBdLDBUhv+8
F0+lBWWnnSk8i//l6CCkGviSgC3ibsQhI3d3oqtvteqfO4UzYkqTjaIiTOupvkmu
5kLIm6E33RDSctscuZW3S0M9aAMQxR+m4wxecHUebI3av10tZ01k+o55Q/uNj7Zg
FBb2I8rehRn3F1a6QbTxI+6mQ7T4M7InON89lcIcO3p4efz5G+mTKHrMKhwiNiYV
W3dPxo7IpRViwp4iyvN54wPcIP0T88PlcVCIH7KU2D8jTfP3h56BGMaiZYm0w78A
vUkVvjR2sfhBjSowZd5A+Bl2hk5/+qCpzm47g72UWyzw0+dk+0VlyWzi9VFhHxzA
NtMBGic0hzt1oK1s7KUPiVhI7xGQBkxDM4uXq2KGuEp8goIgODP09wJJPNWW3PQo
5yRYIuA1SD+1FeI41mCBui0B/Qex294B0KMCSQk4En1HGumXdO/vBPDBGbqKQlQq
PoI/ovjiefQwPupV2dMHc3zmuEiU9aEWAEqaspc9FHnJvrGoogRaVKHSv5orJgIt
sI7Dkjqk8Um5bnyv3vo6HCjqeRE9vjfFhjSJdBiTOgvFHhHw59hO8HbZ035r2yzA
SG4s3ig48PwhfXqAv3L8l8YbthLWhxo8/RaUOjKmRSoWCVGWr7qC6OVvv3QH6jef
Z0NRfAJczK1iU2uEkW3mJshbd6+kMHRz2DPZTK9+qOhGDdRejsOCeCUCKWUV/AJn
8Kphnw+cqAedzLXOfAD3qzC4vQvEWnaxrZNLg/yI9xfaEaMHen/Nd5i31yv5BdsK
RiK8ltFCjUTnPBGqWdfV6DWGQtO0Ls7MP8x7fjSEZ9FqDOe3Eku2h/iik+Nu0lmq
Kqv0xy2JlJVYsu+qVvBxcqvbIrQ6bDIbkPPz8XV53vBsyWbPoowOp/q/CP9+XFeo
eR+HDjPXfxFPG67XAxlU4gL2++zcc2YqWbGL/5+TLP06As62gx5memMB3WBSDPPg
Fa+/9PosUId+aHLzMtR50NgUK3qtdvMyBfexPz19cw3Uc6HHUbtnDMd90ZeSmJ4M
vY7OC7jhUA0Wa7ZA23UEMNThjKNjg5TeQBf4fRjdClhzjE8iOMj8QpkAodedM14+
Y203mI3lSGBE62fWbMKlN/GaU9ohfm903KYvH882zBkzZh82IdkBdE8Joo7X09eX
UmXZpDgxiQL8brqqeaN4166BZG2JeduuIx4Vm7X4IbawnDgqbvfuJH/7mDl+xduI
IOb9YlUgWLRdpIuPb4nQY9tdKi0ZyOOPMa/y+J144NQN3XScG5apzK0cDPhQUXNy
/X9zPkjm8/p2f0jdUOl5/dOVJcGi5DDO/oYI8LxLVnhQRZOpygjTxfI0mTLu132d
3TS5WUJKq9BvmRL4qDItly7dWYkzfZ93VNnGNBmbIj7VIlduH9sd611/PRCe7Z4C
rEocMThNtqvqi9jRiGVjX1sFD4W0w9ad/wkDQo/CBPMR9SXO4v/7S5CkQM50Cx0E
KQKaYw2jtZGEE/pmnzbJiFin1fQsp6wlcCvqb0EfdZWQqZlE03flZYGgU9JdyIqH
8Prs1zZKhlE0L137IKQuKGFQChW5cVgpUYLFhHp0BtUSgKaIxL737AHfu14x4GoU
IXSV1uh6jUa0T5M8PXzzpNmRvmMvuITOvksvquxW159ePLu4hjD/7FugXM0HFBD6
8kuIfObXk85qypoSz+0zhFjRZGDF7RHxl8jUhFqZWwMJYyEjx6jhtWMGiLvc5rCh
UUNHM/qBUBh7VkKDYoRhPlbAp8ZQXpqXr1w6/GNGDjf/GjU/twsMtlF9RXdBUT6U
1AJ+2JwxrunRvJA3UcuRv7M9MJdZVptcgHLRuSFxeRqLaP1nOPU8smDYbEVQs9re
IeoP8gwZZyLcXHEd7ouE/x3H3TvdhB5GmMLGJtsjVzOZxcJim7GUYl6cWrVyiJN1
5InhrRcklJeG1OE+sS4a9ghWyoeDR7Y2YxCRS766TKxxsxtLNqSLDhK2VJx9e8Xt
r8mGQUHlxFlxsTEZy8VV/QB7QaiirJrFe82Y55uxYyNruVGt5w9Fv0ZwNZxJ8mxP
OhprQxlBxmRzi+uBHD1Y8XVQryhZo7fk/EFYOMEvV81pNpQVUVyO1sMCyQBtfxJb
eDG9B7uf+/JZlGvqxw4PhW3DU6GPUS1x8Idf1X72qgeuU3COprIEtMCulYUC1ca7
0S575QYGneo4puN3cLMvC0DiOu9CJM5kuevBToAXgVIXORhGqWAfSo751is5a9n8
/E7tdaIkUKl4EXN57yiRfUYmRAJt98sTPkC+ZfAjJJD3RrMDuJ+xPCWm3fk6z3Zd
bUwX8BSHx7nCHhQaUeAAQPEmKQRs3N6HaRZldgTS4D60eOA9PyXAOYopfMp7iSF8
2gydmNKX4B3KOO3ZzmhTF7Go3ygoAmEhOoccr+rItxvawBqY99+5lllBrq2iFA9h
9Fkue86YeM8Cscoe+3H+MRRWLHzEE2qbM/j5ZHMO/uItpQrUoazSaqWNlOc1WaYk
P/XfHj1QSB400XWMEEZ30GekdFtDWuVC637SXu6jjAD6G8MRSD2qzi64qtITrbwo
L3HGY4Wet58N1Zn8pqlonRmW4gFx/SyfXk1P0bnTo5ypvLgbadyir1gOFC8YIebK
BYGdis2gegIjzEvv98mKQ3mThgxBlcXtBPMtxvmRsufry/KGqtOchYKUbdzCXunO
YoYd7jZ5q7n93rbcuFLMMMTczzfij8ob8tNzwnVdqf9X1SyssLt1dwVHBrvKA9PS
2/6+AWFuO4u10esUU0f8z7qf6LBau2g22oKBlRwWvDGoDLqS65p5DeRwkioagogX
ABnNgU6Pnc2PmvERM6M901uCJgXs3IKAkbMTSjWdjYU1kCWbr1BagT0hoRkQ1zTf
n+q2Ta8uMkYlNT8Ur29S4iUiqfLZm3gQd0Y7R4k/qriz/nRMCgy9TFWi4TS5SZvv
w5+4AzPo8yxBZyAKM24QSdThY3oHk/xQPbAXUbkoMfOPCy4DDUG8IKIGxQThiTFi
ibd6MZWUdwup+luV/F1IgrahQuONpI1fSAOFEUyV7czRGd2twS29tlBaBslCrfIs
XWSPdfgyt2yIDlwMqKejHUyfB8VheeXOQfsVSGNiVhmjnTltM+b72fed1PgnHBvS
6FNevvChmVRu/IkFNu3M9bPudlXgDn2B6fPXRKw0OJRdS5iwQFKN5ocNigiSfSZ+
iB+u6syROirpTNVHQINCSndF3rp4+AuaplpuwmdWgbacG1qXN5dJglS6jkI5uvbL
i6cZisvyIsbd6yrOAghTUoiWoGZy0YAkNCz9K3LM4cDahvTmtXg51TQVvCBjkaff
/fegvcumue1tEt69O1ms28DW9cPBC1wO9xDf5jEe5IHElNX+BZxDs2E+9sMA8Ucj
rZ39mGDZP8WlNT+iNYVSloHJWOYwbl0r64dHQX4lO8n3E5cLfmEugw/JYtVGSD7h
f6xwPR1iKUf1nbVvd2Ihkc6St3LvIjy3UogSoXd2XF97nzgEuAOpoEE5v93OSziJ
hfdqPiW2zP84z/c68wvK2Hn7sZOqfEMaac0eVzXE/1BQYD7eIXGteFkXcQ6VADfy
n/fG1kq3RmELu4Gc4ZsgwUSBUNvXi15VZfBHDll/285oukhTNSrApgaE7wDKObNb
vnDk8Ic+jYbOkaW0ASa16ZrDMJelLlEuHYpK6JnLgGCgALn+rB47Kb8jcil0tph9
P19xbc4Cws9/Ex69kYujX/PsH3bpeYLdAmxEU3HxKOq3ekxYOjUVrcpreJXrv87w
H6bm2xkLGBUw2caYwVf17oHC/VZdxCvr+h1kGi/vJw+gPIABhFV3eiRuQj45MNkt
1/7+odKB5X7IGdxEe569YJAPZ0n5pJMTkjFYl5tpDfp1LDJ5oDAqYU+373GeURRG
Xhjw+mf2FDwqRliAHkbMC22OYK+ntrvC3mpBBWCVZXg87xneqLtIFRhQttPmxfT+
CLB947gyi/XT32L0rxu5hw7AZhS5WDkn1VjUawokGRQNL4V0lsEs1mxgd2XJYj20
KfF8/cvvvNdglHeZnMy/1LX7oVhX971eg6BNlgsIamc34tB0ao02/cVx7dEW4WRg
kTA2wbxg88/4t+p8exRg8aAZNJr5kQlOLWKyXiQZGLhrMaLJHd33FRuc3Gp8cB5B
FIPmb7g+BqLV3ay6+0L+dsfp6QHoYi50reWRTu07Y2qweUi//KhgvoGrjQ3pgFOV
dKCPx+pUH87iPDPC0F2XDwVgqAiWM33vj6CeWIKx8vQyT28y/CMiJG7M6u+Nic/y
rQ10DjeX2vbx9sdERNHgUkmxrMI09VJfBEeS1Wd+s2rJiOo+4YSdMNgPbAjrG2gy
YoHS11r120UB2TWfANBfMRIsBQdRe2nUCSy2Oj4rIY97hJ1cMpUbnm4q0+mMXMvm
rA1E+saOAkJyWnbTK+MiY8x+7n/ei+m/XRarpIpagd3eKuUTUnDzVNNijV8+jnR1
cDQ54EVs1PmhpYMbMS/25xqvUAAwstubpZC0rTYv2Y9KlzqX+p3wIfLG9vOPtL6n
jkJHBvm4ntglYNoEGhao1FGaLU5HGQ8MjWlxAj8yEKPmrKXyqKuOYr+cpfoNwJFx
ntxdY6XHZ9+1wyp1voSHMXdE4lmez71D8SKW0KDwmsxdSGWNJ76lgBpLf7uladOj
OO2H+XOlhSqlgYxAp433LVyLe5Ybj2ZWk486twQNjWTAAxEdECOd+7VsZy6fFpZN
o+RDdeHXRMNlOlU+GKr051ffq/n6Lj6HZAFk6/NNoylV/ZJDF04dJKFwkGUPN6pt
7VCnbUD9DtW7ifMsNkVZzwFfvTKYB+oF2uK6GDTWXJJKT2NAJDtAXTCFZLQhyJwO
SM9A3VR3pR9qxo/mKUXZzNbNpa3ybur1sFsL43f7jiK40tfmrWyw11WvuXUf95rd
8Vutyydum5932h2LtKzPnqiYUBXMbE65iNCqus7ES/HIauLmmWZblxuSdGgj2cBz
QzTSnJPCoPOClQLq7HUwyJYfgi4Xxyb5qKJqBxlBcpODRix2xRDeSjBeupcS0PB4
BPe7yEV5jX9aJ+YSDUpsEeHr1/plGjr/KvBFuIsa/57zhK0i34TOC3kMlGoNzTjg
MQsZkmxlQHA9kvJ/s1CmD9pGef//f0wxHRKZBNahUDNggLm/I6Bwhw2cqzCY3zji
Zlrjqx5JkxqrcBHS7rnkgNwkBJwQDtlqjWFoA0ydYfSXlefL2OKIRlzx6ChUgtXf
K8K5+BiiW5CU31r1UcP+OzId5k/sCuTjikYtUDhpN5D7XeRNmQM0V08y/q9hB3o6
eqf77e9ZTYK/rZy8lPCxf2HIxRyfO0/kkO5o+mQeGVXhLvux55MHvIazYIMpC+pb
WGnjBdqwGMlI1RMiiHXYvYsJgOY5BfSS4wsORqgGxUi7fKsLMqTwlc0wrKV8n4+l
HgUUtkjP+Nob6hvnP0M0CDSSOHJRFKmDfq7xnXI15v/tJyHL5xrS91VjIyVU5EEX
QYwnglBdO8NE5XMevlVX5i8aqAqvR7DRUuIS65fOJELLn8XKBUtoclhNIiP5sb72
g+YRaADGZ1JLNwQsM7humwBhdPbrA5JXjaT/U91I6kML2x0DhpvRos3hIhclL1Ji
Jq8I7Xv1EatZInn1w8GruvzO3cPvEP+ugVDwwVrBybwX+IEUL3ndHmNK1gHmsYOJ
IhdSZj3ml/KMaU03wMYoV+LU8Ji6Gwaa3JBBCeKWTHxMTVncYx7pGHUuP/zSr48H
N23ZG7I8N1uAfhx5Ihoxt8U7/OyFOYrXt1H32D/7KyeWondXxs2mtoG/ANZwCGRa
eK69n0FHMhDbsZNT8k3WKRVLYqIwstQoTQXxkfIsO8uPcXurBqm1SkFWjlGbHW4m
obUJcnEkOPAhv9EYC6BSmgSHT8hri+nSMQKqkus0pjoprC2jg3ITqx1R3q++6EkP
Imh/CsgNxd3dFlhOagJ52/f3Vfnr0JX7Po1fviXCYfM7wGI0EZ5Zx0RGKlWnmBM5
ATArLeBOPyWOexj79dSPEwUy7zrT8wv6lSkSPIEZ+2l2+A5EKQ75yhbxeUjNg3XV
KGFg+fvTbsB+xFCiEuG+Z1W9STTxjNyjOAON5kGFk7ISjtsCHKdZQNKG4SD6qV1N
IvfwmzzwhcwbIX3fLd7FxkzNCKiEKwMjbpDrgaTfK3Ulo8B1Wf3vgjnwWld/lgRG
3+J0ufAQ09bD6QK4s2pzTcPOvFqFKmAI7lsApdMH/VtgQNI4hyCIvHgBdzcWX+F7
SNLpAw/LgY+4HUm7a/UxM8k3AcBy5z4MVQhjj2s3Bz8mPuhpF8V7++dYx/CF6WFx
t7SbjNDgQmXESk5geI36keV57t0PRia4+1hOEv8qsZ5XiM3qnRzbZXDMfrbxUn1d
XAL1qaKJy6/0pp9TVNhVR2Eo6KBM9eAbPCDyG3yRvpsRuEgSOpW2QRVliYx6NK4R
3A98aRA1xOuw2DfcCM+GeBKgWM86+Sr3dPN14wKQZAuS38c3tNg5hyKXJIgT48pE
h/ts+PZc48W7SHVM6QoCfRV9FPfNUTov59OF4IQpA49qvyJ18KJL50hGX+CnzFbP
Epsm64mSInY33RK5kHM+H/57sgVPuCfwjomRU7jmFhLhu42cvDfihjF/yV0vRWU1
nBcmSnVghDShm/6EfnvBux9hl+83ARO+Sq5VQKuqv2HVMFqglNrC+7BmugL+ylXg
zwwZ73agckq2mgVi0c+PCpTGLOuH/us4TqUkJWgOsSBEhtxHNVbLPPwhKX4/s3T3
fnVynjdyGhr94oYJlXnlJ9eXJzs26z51Qkztn33VFsp0559vrdQEco9b7URArX4a
nV6QjzRB58PGxjbXxftkT4+wly0HHi0wxx0/inhV91j8m//r8X8T/V8nTTXkeiIH
mXv9VARsWKuBi5fiGMhqwOtsyls8CbtkNXG1othnen0IisgA265zZcVEK5/CJoFL
THfV3HlPfF/9kWCzA78bQg/1iSF6B63IFrz79mWEnGMiwglY6A9zhH3NdmvD2yxk
u++goD0psPDfFQh6sBsYREuMIc2OBi8gomXwjitlQHiV9SF8Fh3IToxsEw1TOeVy
9Gl5ynMK/PXtvWxDCkgYRribyUO/ePsFunGyoBU9ECanqpMUOuv3JViyHGoDZVHY
o6rLjLDYvwoLLWhg0BCQgjpuP3rA8awi6JbonY6Ee855tr0CETAc5ci6z25GlBca
w6y5uPWjET54g22EL14/KBB8d+ivWn/EmVT9SyHwx+fMiAfzQVxt7C2KR4+NCoLq
Df7JhY+vTFTVYWs0JhtpL1inAkV08NqTLtVzJGlGXliOv1aPqVvB7RcyFWSqDZzb
vP+qg5wCVZUJ6sprQG7TAQKmaeGqYVsshDC+N9UJ6eo6B8p7ZwWJWe3a3szcjb4P
oHilrDkF7AiimcrWKkV4F2NBipBOYfV5W/UF6LJS2Fp0kRnFmcvud8r6TewLlhcj
GrUztdb0lLKeHxv6mjookXvpWC3kPoiNIrl3/emVVGl2jdwBkAlCaEmoVtzwGz80
l1q/v8bjSAX+XcWEmV3K333bgcCKjizl2HoxMoDLWqDbVwZw0uY9Zoh4GIPEKqRI
7nNjVGNnGsZ7hfAeXVEKdltvDa3PSvyU8DxE15jWhSFSGqBI+idMyifpo2X4GIFi
936rcNNre/RpQFmJlUJaqtYfgFi1LzxNdS+FGsnqyQYFntSZZg+JQTEY6+JzQ6Vw
GtM67DYwQomxi7JXEZN912FXezqTOvuElL2ohZ4chzb6/izv4o/TIgAx+6NENgVd
ekC+w2k6xV+kXAaoW2BHkBGYc12g28zYS4592KjxkHQq7sM80DowPA4H4Xn7DsII
sOcvrghYVAVXc6VavRi7tPAbTb6iQwW8LIMaj7QqNRsqM7Kojwu/LMTpnk8ga3LW
o6PYyYAUdSj7/7aUCKn31qA5+t0zymwI/Kha8e/mdoZgocvgwq0GsdcfT44PYqUM
QbFZz+IhWcmfZ+hWsk+PrTQq09XKnlx1q/mKQUo/m72bGfaWKv7IW2tXS0cdThRJ
vlQjTAz+1tPcHb1LATCcVo89SuVrc4ZUgu8y2VwsxkDh0BM3V6U/LKUYUXokeXUG
vxhbDH/1l8pN1WRnKWrb0MGO0biZ2aJHA1q5D9eOpXbwum1iMCCH4t0Ofil40bP5
CkmnqXi2cd0HD87oyps9GcBATE7psclbrExCuaAvEcXUlD9+56iLVjhIX3gDsLRH
lcRFkLXfk6wQ56cnFZaJcGNceNPcNynlSSoDzX3zx8ttqzQ47+9U6IFdjC5WfNxm
nV4dVU+DXwTkNdDFAX3Xf06n9Bm0EYKfOfNDYUVTL0gfxiI9JT+USuBEluqGwVI9
OzPICVyoxBmg308hE1KCkic0xGwxm9WH6nBwOyelm7omVsD0zo4SJLjeulJL9iXj
QPiKLnOgq8EVI++WcjD7IlhlNr2j89QwtEBixlNkf57n/K4BWstqTIXcXRqKjlYJ
X4Vcmc6ha3aFjHeEb4ne1ZlsPHUb207fdKgJoM7HGxJURJIFLN3CK/7vInAP/Akv
JDj8yoZcnSZAaQISjPVv68y6OkO68qKnDZPrTRc2dI7Jk+OR9EqlYe0sBg7Dgbu5
RefMurajOiiOrliCNsmCm6YlqNLH8bdIxSAe2nheTlI3EQdoOao/U7dfIkDys1Ib
ZMlrMmOcWDXJACmPdmtZfd6bF2W9ZOGXqiQRtj+PsJXzpc3xcqjd42SdABS2LF0K
a0Us0IzUHIzlj/LNJSKkvEilOsVMusf+KR1shn8Zjq1dBkcR/XaPNGd7pCmKp3AQ
S/m2SGg8co21gPBmoGZZIq+0ll0IORzA8/3WhJQoS+q5zD2nCkwdVuKVWUxbu6H3
XKMYsrwy233FlheuEhj8TBh1URpBZQeJHKJgv+8uhqtHLEogGw+39t9CxtEkTg2e
CLgWrAX1T7ScSd1v1pXJwy4k/W8bhBcU359MxdKGW4KA+RuQilriqrUK39nKiD6n
KKKiTJSNx/pdTE5Uro20H23bp43D+8m/N9PmHAdN3WQGu1Z02/q25nKOKHquxUAX
uc50/SgeZWEuZz5qFljZLPqMG0+iqaQa441c3H/a8N+XscEUN0mHza47PV0UzOvt
c4K3vFCZ1zm5enc3WcsB3LtdA6Kx/qhIOxvUCspwsWlO/5hLs8PszuQ4PZifDT/c
waFS+YcTqQDBpnxD3/IoldvXv6piSLDRJOaNMjRE/5BYgfMdXepqEjZvOD6ve4IN
f8wSJvSvoW1LUIEXn2mrJM2vXWlUtRWxTcMtbRTMLPBZLGCJ1OTI0z8JS+IP0pGe
fi2ruvnK87Z5R3OCfEavEeadxvPwJpLS9G4vULbs5VqorXg0+JaKUQ4J5pNKGrSz
xbs4VAE/fB52fdByvTzxVItHjJjFNmxo7VnAzp4ol7UhGjLbVxzlAbB8PAe3SUvF
6pq8vQgDnMbkNCQ3RqvEJ7mwhRHQRwIQq8Xlo7YQ1aqlSOX+9gkGOvgAwyeqsjsH
iwhGQILAhlnZNa2HfR7vY/Gcvd/CVo9H6qdS0FqLcQblRTSHjj+dg7bMLaHaRNvZ
GXIrNfxACl4t6K31JRSiLporY3NvY9L0rcRHtfLzUMCLkXj3z7cRYpD986VVMDRV
H1ZxDg3RY3UjISTQE0KvGvDviyxbKarKGAXx2WOEeZDuVyRkwdtemOtHXB0LnqBF
MTg3cGjsgF91YuEAfpnZDqTuvBbZwVvt7rs5M2dt/NeWZcQ8e7q0Jjcys5kfRDkK
G8adgaqDTl4ZgCUQBOhNEteS7HI9Eq15TO6EgH86J+aEWl12a++P+NvXyigy0/mp
w+2SbJY1QjAENpO7o8G0EuOJo5e5ZKrXXx6xHMOdpPqt9IeUoAw02qwhtMfu293E
qpJgqoQM/vX1myoTJWD6hrAp6I6bwisdMxDZEiJdLDXzhEN2Kb+nM29niT3BQzlj
/fGCALTcgzGZQ8DeCf8NT7qNehBgUF8kF7OVTYeX2SucGnK3BdGEzuw81qflqfZx
LK1Kz2lhB94zjwrwqcD3Y/TofvlOK0GlOjzvQSnYi4gUn2xdGte5azi5O1rNgmpn
ouNJCBqxemY7oJIiCyAi31kMHFVxbimvt2GfYY202ZdJm1q1bLA1+ib6fOTMYB0S
TumGO2+8Umz+qrcJkMfZQd1THXfgWjs1iOp6APfy/3QyhCIrGMezL5aVZf8N9W4S
jUQWiF8wM3FG6QRwslaJnWmV5CLameCiSlk3QZx5BSNhkuFGlK16wNLp7tPwyqP6
D+06mVSUh6ubT45sNfZrlmXO1ztXJHCQeSSw9Hm31f5Sn4D4j3Fp174K/5OIDWvn
IZJ7jlg/Ooefxi3tXqUZEsc15CacNlbsG0zzNiEzerthwPnU8ynmGTB7Sq6u7gyn
vfd+7SFqp67/ZX9w8Flt7RzEiEtdYs0yAkkf0yEZsrjUQ2ht4QcGE2jSuEn06pXM
89BsM7+Pe3am7xUCzm99j1f4jCE66oWuLXytz+mmOVVI4Nax65zA4qurSd7FHV/0
Zm5GK8JqyirPZQqWRa8nXtbUx2pJhYFtbetniCq50ZKELVtovNSr8zt8DEAkYLdD
Zmi4o4H2GGf7/2Yn7jELX+/4XI8rH23RUju2JMx6CIJBdzo8Wfibx0B/MhTVZDgJ
vKLAWs3Lmf4it9PM5y2le/v6xFyAsH2rMRFq8ROptYrnLegiKgIXgAPxxfFoFkQu
hIaFSI+fuh3m/lWU68/oBtgDy1dWjgLaXSWePslgCq4R/A/i9j98Ru3KorN1NtMm
25ul2bWMVAYz8ygyK4Ec0PYTXMz6DklbPdxZ9AN9ICfaWjO6NrylS+WhOfVPaDBD
YihiW6hPUbqcAnK3UwR7hET130jJswoFtlMalTQjR59wC2qc+UUay8D5NT+suOnL
B3mzLgT93NdXq+v6GnOc/o2vSTZQTGUt9lhsWYCYAEWWEajvYTOZYfpPkXhaXsrL
2HioJvfPGfsfPoC963yRyf9sFxmfdUd4WxBqX5PCiZm9aR9Hd1wtcw7jRGIgceef
A07zos+SD2RTNPxiPeW4oc3WJM6UkN99jSPloxmwvkr467hdsVxu4aUaIZrvZzB/
NiChjjUWZiPQ72dz6FnEsJI74ng/ZNZUZs8OIkOlVKAI0HJO4HYlByJZMHLAxCa6
vQ7x+1GMjbxf8kF13+pkD7WH5+dV0GwJhsR1dC6p2I3aejyrEmcypt6r2rvY8s4O
RqfGbqdAD6Fvj2rQhJ+hsatoOM4vLbHdnPsdknrJ0Wk/HKmhNpoN81gBoFwX3OQu
pst7yPNaA29gFaryUZgPE+nHQlmrh7QTN9UsiN3Doq5PfBlNFC1x0166TTRtFPVK
X7TrCJGgjZYGy96PVWHnDhG7TMROt/Vu1a/fOTTMhifMMIPjaJYxsf4y6DAhlgfF
xPAlMUto8Pza3lk5h5BUyJRZKJvg7IRLHZihU29/VE7Uf13TRvYOg7azkH+H62IF
mflZ28iYZXSTkHI52aYhLU0+JuxtAg8LO8XCTtloA6e+SOxFu2B4xdtb+LNSern1
J7achv8X0WC2IPqQd3/2Dd0mJQH/1SXwEEmNgpshqRpSIi/H7AS8yyMnhYsrjX8r
2hiCySJYzxMcbihjdIaCcuUzUbWdMUrUuH9P1shxAERhScxbiPHwyCqS3/MuLJUT
l7zMynmbSE+boW+S7gfX4F5zuydzz3Aga+pSXZgdCiiDR4Tlkh+8CIzrToLJ3iYe
BFSND790h1tNvp+NW2aL9xutoMlvjSrVq6juHJmWj+fN9gL2HG7EdjRK6kItDLzb
G36HpgE/ZOkt55hNYOsvBAHbPQD3LXseelzDt2X6G032MmW4For3ZOk0zXJkFJe+
0BorM+AbdJB5Y4wHB71vp/lle1o5UbgT9XlJa2crw9J2PrAqPy9XmmmXICmSL1wc
6ectCroGR9ZyILF05aX9m8cY70rHDjHWVFeXLivoCtSUU7XdzCuKnsyNdXy1J39r
OWIIxfqElX4Z6Q4TNBXXBjVdkThBZfYb15c0wrFegIacgc48tiFqGqxOuNb+1XYb
nzWfWIYzFFE1Zk6kvSUZzrolmPFLl0QpQ7JdqJCA07Y/ikHtODT3hTp9wwoF/8FR
Rd3kfYsqHGF1p8VZQ/p37KvSVDnqJotAs5qJ0jkoeTf0SiApVQlcRw+qTjSAvYXr
brcHYyiIhuyEFXL/v6a0qqXtTMsFfLin735Y7NtfkWHRkRn1bNx5tnQs1HnyXF5k
q9scPGU2cf8cWt2mN9yo7Rrvk2BHvttukmju5U9vcEQko49u6LOWkjZfH+UrwZ02
LwvDMxMM6FPnyICqpaJIdxF7wnAryUFiDGTa4VD0B1UCsl6nNOEuSS/lblY0EDUh
J4WdTmqyKdMZVCrHQ4kNh1pYKw10HKaSByVEjocgo7NX7x25xbLKJ4Jsn3zphFK4
1zpWtcqkmVrgXrRVFMg4cOQX36vL8l707RK60z6/mKz+wIiBVebwDufI2/PfJcqk
vMzS215vbphVFe37bZ7qvE27Eo6F/UbH8IooZj+zkvCOm2BTY1+y9OCBZfKD+af5
FX8kMSykf9VX7EA+EAKST7gNI9dP4hrJKQM0uPv48NNevUsnpizIxhWGtXDDjKkp
qgREsQFGntIIj+nNYEZIKjkpVKIgfKAUC07R7B6trPf195s4YQ8fyOhaQMWb9K/p
ys6JM64U2zhmZu2E47do4gHf/PuA7WrP6pbvEj81izIJYyxC3WL/sZXOLjzsCXU0
t3Zh5eoouu9ABBrXi8YqXQUdWfB2KFlkcF6pCy0v1idW9gFCgxtHznK8P6DlYW+c
5b0iWwVZDfgfDrG6L9DjuXMlBDjpW/VwkR1b4fyTQ/p3KTyxFxtnDYMXQ3gi4lrM
wC0c+XhfIsHxG+4w3KgE3pkJIBD2XLgR+TRalDLz1c3+58rBXYG+yMXjWW8EU2ep
HY9BW0DwwPXpjownfp+6xZrUaahwnnhRIzV8JWTJVUhXmuADxJAkeZEJMSLmbFQQ
8EkgcpnUMJH8OuPsaZpc3PgH04I06+ao1YjOR7kz1lgZHo1bLpqIWlgjMfstPCIw
vertRptbcPImUNcXsuh/pSwjR+RAARDCsmg2IHuNcSHFfMCYyfNkR2tN3WQuFQvf
8/tpVEc7sfYUTJvR2JelhVkjKV5toNbzg01J392+ZTSeobGxBqf6+oI9vmQwaX7p
P5He4Kpq77ZbRSi6Eqp8K+2FkomdROWBhzaZaevnHAEG3w2gdCictl79BB7grgMB
IBkPiulXTPteOZ1U1KGBa2gQzG2t8mw/rBLww/ogr9NOEu5WTx+1RE23NL4gZ+x8
nAS+IXGyu2rDmsFnFyeWS6pwq6WdNTDdLpkpk5d5kjFHuo74OXnfO+JvW5Xhqayl
sbWyb8bQgSLzTTJ46gWaDItNblKBf5mjPSlSahbp0CDUb1it8OzkGNprinap9KlV
V9l7/jY/M8g1j+rmtYK3Rb0W0dz+f9XgTTs/o7Kvj9o1uOuDanW/CRceYHihKUkp
0xTF8N6fJlk5GTURSDkT2Chd9A50jbTTvFMoBG3EkRY/GxXfV7IIfI+eN2GGbiHB
Oe4hK4n9tfVVSMCnXBbqFLtuANR6LdbozQYt3VT4xY+xkXEDIwIJfsKV1y15N+kZ
zatQomLkF+eKZYPQ5SGWU+Ac9tITlTeAzeL71bZQfiad7kNjs53bOu7oTG7t1wMD
61513C2bxkC0c1KsmMh0Gm/LNJurA/2m3qxC0NYohcnCgt1d2h9Yzte3UUvVj2Xr
Zmzh019NPBLtw6ofPU8SNkwERAEBCIsjatVym+vBkWGDlvx76KIJr5WU/NCKY/lh
XkS/z3KyC0lkwvQ5auuLqeqWzhHoJ6CTY4CAUeKKJLwey3kB7Nu6hGGgGSZr9dxM
9rG7dJvLHC9WFnq4I1pIAHb4FADJVBz+TQZ63140ncWYqAupghduP8lNQvDcQe+J
N8q45RpUfCSvMhVJeeW7UNCCKZrDXd1EjetFOz+PAYLtJMm/k90zuwAy4GUmYP0V
wd08R81Rbd7esvqpwan0dypJBM6DO3wUj4IGi/wqmfuq/SSvcOpQM6IHWQO9VmkC
F/Be11Z4Wc9s/unAEGR7FcyMAundUEa4RvRk02a1nvnYVEb61j1FSxTEgzrbOf3Y
FL9hpsJjrlvRYQgwxB5bIo2WupBUz3Dx3Rj5o8EM5FU/OXMgHhPZOc57LJBRjrpc
vdGFzoN7jJtDcgskctVKvn//pTAD/F3KfPRqbtoPWl8jms0y6BxVxdkBTVNQJY/e
FlztjbQkK5YYpzVqZOYuzB5vtM+Uzi6GpbZo5TGzqEtuAzJAmKZM6xElJcBVpR6D
ecY6eDdjWUsrwurPe967FyRj2gEs1bPojxUFrauDGlcqI99WPLRJpv7k+9W3CqOV
spxfk1vD34lq6Vm65umpjWR9oYqFdEnhfS47nf9kfpczDi6dhzLOOvQBsReobsil
AUbTZX9cE/ii8Qj4hhW0N9Cz9farBVfs6Q6rWvAEx+qaXNRkgJvoy6JozX8BICcW
ROZMbKJ8GlDsRvB2PZ9jM06OOD9wdNmNM9+e2i3WCA29K4KYb8+gxw7LYWWa1twU
sUJXHI8XVlKul06DA4+XZ3yg/njUhWgcZmrvblVAC1KKyeg/c3sRUuEKPT1eGCCS
6Xo2jyk7DMEVDsC21wcomtaal1vKnmlyDis7Fvs+5+nsTBXmK+40/HD/k38ydhGR
/qxr0N1Yj9DI72EOAnrQtFMDCoWHOWTs1wO73vuws5bCaIwOlIuL7uqDrsuef0YH
aDZ9iXj8N8ytbTcGu3v22362vdEuWXzh725wAVwdxvhOhB2wJ0XblbM9bCENo3W7
FWq6p6IfFaftR1rSMpzeZ18XcOCc/MdnXARSN2g5B/lAm51y3liH5E0kIXLywsNd
hz6u2fvy5dvquNALXEaPiDr4w8mNFTalur7SP/81mF8EM3+xHhpFvcYBXO4UQgVF
etVegckyrRpViOsouSl0Jj60YxjJKDT+m8ScRFh80xJXMRrkQQ7+yyVLIhf8YwWM
HctXS8jMqd39j3bqfaBp+i8UHEuAtVoo5uCZYQjipvY9hVKbLA+xePspJVwfncUl
6Ww+3pcfkPjUAaobMyaEvHVvqwOtInZRXIY26S6J21Bxp/A5fqhzgDtfUcQe5jLF
59p/TxuN6xW/1tyl4WNChDw7YnOAHt9iGG2klETrNIDMMgDBp08zW4YpYc3VPP87
w+NryuAU3z9d8Wv/cBC6f3vI1cVJXbDw7iaVr6oldVr2Nbg8Ev1/AI0LGQ5ojcJ8
bPh4owr3uobRNXRFYQAETdXyYqrnf5/D1aNJ1UWF8blGvgedsM0FOooqfe5cEN2F
zoeh+idGMWaFhpQsPy80kx+KtC7hak7lB9PM16Eu0WWX/yk98e6h8VlA6bWV+TB1
uvBJay9EVd9y6SmWb3phutbktzO83mdvGhrDVRknctXz8Y6hDHTOfN5wrwe1i09X
ffwwDKZvys7tuRjMsBjMxB40jXqhLalqTMZpvAHnT1JSUeZ0JFtybaO6FQsSK4S1
wO/ZjfHMOXq9c6cojXXLcWcXKugxysXZa6JTl7J/zB7POIN4wR6Ttx3lJ1lpaTjl
Br9Ivvx8CuxTFDiclSVKXAOUfCEf9CFuIMiJa8XLZyrJYMpn/lxyJ4nInyyacOTC
UN/rdxmMj+kx6EQPiPvOjwVPpu/aSB4BFpaAoBddc0b9TTTv3uXHmBc1ykhOsv9J
9s0IveCyzKcfi0M5G2TNWEN0x9YXU+JyDZnf2E6iEt+fnpSrObeH5N8b6gaH4cfl
0tS3ay/n2UX4syYl1CwrTsh3jfbjyDs+fn6Y/XRIxTPjz7wVXe/+f1TfPBPQ6pBf
guM3UqxetzzxzbK5UTQs22gdQtCBE1gx4YcYXU8JVzutwm1E5QPHtYk2UoGexjlW
ubqeu8qodmIw5+jsqQZzgptiprezMcB89l5AfgU6cKKkV2M5Wk0ovu+GHr0E8NET
kkmCxgiyAp5t1bs7jCMlFELznlYDwVIeMpeabJDDEgoRiSDVR82uEgI4J2A9U9Kd
F727CMkDOHy8eRqwtsfmnY8nN5UDISjWrNvbzNAdVrQXbE6+4/NLmMjZN3vezhh5
/Wzwq9qhAwraSyMBr0bncaW8o9zgTkGHX71DllpTP6b49flAzZ/4OByJZU+9uAR/
g7ChGixneJ8QO4EZOkd67bId/A8Bp08j/30fias2inS8CrXqiOxPxHEz9oTi17E6
dzg/m46kepAMnrWS09/IhuPYRhHSuY4XgV2982VS9R75XZsAZuN534EDL7hNTbOP
7LzeJmHEGCPvSb6pTlzgqXInv/okdVRou98j85GW/l0uRnZQw4UAntkIqUw9/dBE
+rZH9WgYysidLFyIvinKIOtk4P+SKnNLegTZRdxo+EjBOYsW70SNV1+bOqZ/gdQq
0biomAMqaGzCw6GT3iDRGwBfQpScq9/bGwuYboS/6d+O/JpAN9IkeZQVRrxT6no/
EJtgqfU9aYSdYL4zcIPDjE7OjKd0Pyfe2mBt48jLG2yq0U2ROWw+bdrmU7TsEK7z
gmRma5qDUbGANr5D/11thPq9DHhpXS62st01KfkKZViVAkNkaiIac8lLEm6bRyA7
q3l5TFm9e05XpYLIFhs1qgNMyC8C3xENiPg9s4PuZaODE6y26q2X2amZOTo5shI5
7inn9iEZgjFsL1d2jHfFm4hJ2re9DLgHfwx3Wtf552ebPQlmy15A68CDv3suSYg3
ipWnuSzTCnkqVhYoclXD7dG9wwZNwzWJK2FtYlsulcAgIXTa6g88pgi6y+annhQX
wHX4MJeuIb2HgdB6X5x1qL7J14dpUAgaet87Da/RX4Gn2Ns7NwzoLY2Z5LL9XIkf
Etjxo7ensMhabQtF4OWCo3xrTLGEvmffVfQ5DNQLfMxtjcYDxmC4tJopfeRgF1JN
HFgLM0z0K/5SbbaJkJGTZQ0N7frzj/saKK4Hc0pQz5Da4FxVk3v95R2VPyOh/YlN
nTIFMGTzPOypCGHWRmTIaw6YovBu+3Q6m209svqRmKx9xg+ONnIYG4T2YJlGFPpW
o1B5XSj6YFSgs4/xrKbjxNE2RN7uttzmUbjQUCIqIeWpeusFjfn3T4fs3NTB309c
UBEDcvJDzpUupNGV3/pSkTVUl2RboWq7+BEs8m3MmgkVrJ67wFiKo+BoqBTdbvQx
a6TouTbpV+1utMo4yNp1TVyWZeQk8oV9XwaMOrgBIS0AvxUtaWWF7opL3yudz4Lk
CPS3U1J0kRMKUuhXxjpl7LexaYv7NXcW5ObBHmFR63Vf6h3rxi9nueA1k8jmI3dw
c/A2kWQ+aoHfXLWmD1brkTwh1fuSc2GXHvAHSup1KkvXH28avSNpYfOR3FkN1FjS
SY9UaDDYfjfYyar66OjvPO5bgyhcmPbk0UU137r+/68ndg5JOD64QBxlDOQ+POKF
R7CiUgCLfxso/T1LXe7WuvyHvL662X0Avi+WKnDYRZD8KoU/B2B2+6y6iRN8bet6
ZL0VZ8+CW9vpFsNGPBYrwfPyqwFSFkfsLU/mys0cRLAYFreaNl5QvQuDE/jNlm7Q
GuY0nyuFlX3X5db/jm0rfDQROX4M0Bl08r4CVpRt7/o4E3zd9hRdMldh2FkA/fBb
w59qv7uoY4ZES/U5vnyxKadYTQXT9EhtmfESQ8hAt730Yla2RWjWOLtGwaYlRbNK
8AGNlgxZinAYx2JAV+JGJ/Ym57v9Szg6skWK1nIv6D8rSBlkOpwKPRRnQ/JLaPV3
R5UBvOu0DzbyG33RV2JsqaiCOtSL3Phnw9GhDjRuGsfDKRb7dt6dPn/MMqXeaANr
NRPZ3zC11+53OQT9kUK9HhuiZiqhWUvwRtFrehYq6Zq4hIyA8P2eP/VmPxugbpKI
s9oiSKw3uxulcQxT82pqkpfKDCYCVCEEcL3/Oh9M1I5UCcoGlZ3hCToJqbhlh2ut
ERUTv6rJiBqSNqRPA2mW1g3MbJvXCGJlCPyds7zyfVcRXC/sOwiVyn+vI7goyhLb
Z7v5O2B7LMGp3Ouwh7rzXtevdJ06wZNQQWSGTGRljr7IqK8WXfDYb3oP/UC89vng
e7DH9aK3ZS9NFtHhE7Lyespl5VDNNFg3rBakzct8wuPNACuq4/PHeLJOXJXl5JYc
CK/5ReWowBGA/qo2XPFNnm/JPt4jBg7k2aBLcCe1eZek0wf05MOKLM+GUhRskQXR
qtb1EHZSQk51gqfj69PU1dTtSslAq64bYzwJ/tFVLAZVTMVzSk7/mGPa/Yj5ubd9
rtIWv0rVsbiy+kbKy2oRZlc/CEERLkF7ukfY58FWOTNrj3qrr5OIK3ARYNN2vtHf
AZ3NZ6Mesj1/ICgto6gow6D9ELn+TpaTwCKRWCGECvleFBTxxXsJ6ymSIIsW1zaI
VvbrvAqu2Sq5H2bqpaKbr+yZfaalG5crntGIiSiDGyqaO+nMBWCFQr6p6YoJoQlr
bitVl1Fp1yDr7nHV/a3jY2CVk/zTtnK3qvjaa3KDCl8SeB4HtTd41UyTF2W59kFh
cTmpYCKGEG5w54BcqppD30Q8cHUfPzmClSq7tbNlghu+QoTEcCd/mXdEZ3yS7cHU
OFYDw0jLisGwYQmr321kmK+740PC7FKGWL3y8kVxoRevOI43eupZJe5dKYDjnbd5
B9Kv8LpL0sdBYxS5AZwGvNTcWCBlKwOR3DXKQ2ajaX/ttdmtFTJ6b5QJg6x0tLRH
6bebJKqJydOX7g5eVTE8XcPV+xxjy5XJQelu5mHF3INACtmYPoQtqWklGpdKolsf
CAFYY6DBsmW7M2LsEXWn3C+OeWDU9StpL4ZEcO1kSO9SUn6oP2XGOuPMtw307z6p
oVSBKGxpaxA5WdCBOizrWKtSgfTpnBfNcxc1y4FPOlxZF8vzQyn6V44PwamCmraI
8YiMn2iAUnRxAwW098sgKs8STltgdHbJr0XSFT6KmpUHiHr8MVaPRhDjqagqiPRI
X6jP2E3o9hDO3cej3GZjtvy2vyDHfRBQGr/E0GninVuMl6IylNQ1PiC727XhQQhx
Dlwx6nbCYCCeIAkKLZVlYU0RN5bF5YGyE20RnConInrpU9ONjrUkhsEWH+lszqJk
lXEvVyI8bl5SBh25AokrBKNVAVN16hh1MvZOlFbdNUH5bTrzGTxOLJj/TxJ7HF/r
ALngnPbYdOAUhys2yq+EFyg11k2eOb3hjcYE2ri3JhghZN6uyUKqpokoyzhGSSVL
6XCmrY19QeMHBz7SvFN6EW8QS7+vitqfAX+LgB9QreRYhQGz2yKta1aEIPepTTrR
MxWDDEMPDUzW7NLSsUoasiZ/+0AdWjNUrhW2+/TUptaaF/Ios2FmqDrzAdPpXb2u
pNK3mGspv7LuauyXPXK2SfiTI05DVjxcQH1Z9QbLtFvHDwsluUE+/Wcv2CxkLbOI
LlcynJdYSdlj2NQIkQZUSAtSM679h/FB32QYVt9AIKt2F/MyCW9UamAgGhOnLUzb
LP7RM5LImLyo5gjjhmxuMOTLZa3VaVgUInmnJZHzlpI+4Gy7FrXaRaUeXA/nnPxi
NLEBZaKkQt3wwvqv5lWoMKslKXDmk+t/clV7CL68WG/IPYkjHTjjByYkoPusom+W
8uZfKKSHPPnLi2qaym3REYTgmJxbgGdrdAq6ib9OZP+sqqhnF2jpJsAikyYEerJl
eKf3gkOsx4cs9IKZGMO5iFGuQIwHDhBh2wpnbSTqZlVhL5prBVlq+Ps6Ncjxh5Ou
3Drh3FaDDYz1WknBvdzDtAp/rtvdEsxAx+3n11jtXEmVpkU2S+gGIwxQvmdXm0ys
GM8z7YgyLjD04mKUGm+kBeTls/hsVX4w/c/K03+nL1ruioOO0+ao4x45iuQiUbc1
6Yqrz02eDPmb5MSmSbA9zasCQuwSNDtYsuPH+D6qmZI/1/P4yzBuZKEBURWVbbKS
qPtlBhG28Q+VF2NXHG/7CvbELOiXI6iOsUTWsJNfMF8EDhSWPUesh5FH9lqc1Dzy
mJd5VWFzi6SFA8jFznIhpC5lWD7C/F3Pu9+q3kDdJ/0AWjQejYf6gbaQ7EXLzKr4
m4Kc4AOyjefgqW34PfNpq59HUck+mVoIVoBKgDga1MQfl5Yzr6rCgU0r6l7it83o
VXTJ6305Axf6FRxR5VSvB05SPXHdpmQdNzh5Rfz4/ccvBq8JLEVTs59tv+ypJ997
WozTIom554pCh00doZZH2VYU25OQYwrs7vXhCBFojD9I54nL0ElcyAabY+EfNPxr
QJDQNgvwx9bdSCy5RlpepKwwFpied/ri1Z/+3vZJ22SayrdtKChJw7105a0LdUT6
p4+NtIMYAo+xj6mF6DSCHYsejnzdiLG2nT1U+K7XjpBocDcpEz8oR+rIpjg3ZjKi
QHHsgROM7N/xfC8wKbF59eD1VNYtD8XmFKVyBXVFo2oaqTHjFqR3rUjlb9zohcpC
Lfb40LCr72HrQvFMAtGPpE3f+9fKiaZnH6t0tF21O+sPzYh8D+w8pPVDQKfI2t6D
M3Q4HhTJBn56I0jU88+hubzCyX0C4MWSi/mGI5e9jhO6whKTvNr2WgvJyCFrCmZM
ZTgBG1PffUT7pcLonBpswUSCUum0Eyr5C5mJ6SnyxZ70iif6TPMqO+6VY7XHIyR5
hT4qtM0XpAIEV8EiFowUQlTeAihIXwS90IwPTfq+G3Paaq/NzuiKY9QKobBzBiWW
MbijmtUvMVEAaAJQlxeyBESOEsEDCDWKaeWFYE4b4DFUnJ96FZCNRuO+SvqAuV/W
bMmre5Z8RskWGv8cMIsMlu32NtAsplmI4i99Pi5ikHKwIyqksA4a9dssNNXDHj2Q
1/ymgA5Kwx9/QvZpE3+3tpM97XfKOAQyRNcYnWnrIDyS3W5N8qPssuHz3c2Jpiqa
r7nnlrcuzdU29Qun7eS9q9CgcmRy6JtnkiG1PHr33tUyl7anUNkGpFRdsOic7gXV
PbV2l3z6cMviXKWEsPRCWP26inpZYbY9tRJ8LgzPsMuXTMIXwMOE4ZORmCL73Lso
nBPPaLpdq/e/nmsjfiM0Vmv3ZsPY1/zX6RvhqO4gny/Np83MM3TojH3vZYESlIKJ
4yzfBxmlGvnVAbJMbuRiiXVvV/xRbu6OMk9rM2RzlkRT/hy9AnrNFq256jFUYimW
QoFxbdj8SHy4VEwEZ0nvldNILEg9h66tmCQ2LATkadYVnRblXtk2prJAPiRJDzAh
c8K054sF66p2gX7dOaE7c2F1QubG1vZQLBNyv/NCSwKXki6yWE7p/MECfCz3BUrK
HnOZc9C3UquXeIxWi27Ux6xoWceoRVWNlW+u8I/gYKpJS8FHc+Ug0wDQAfb2PmZU
5d3FKBz7ldarEikEVJqLN3VmK6zOHAdiKLYpOzAHFR82jItdD+4mzhTiD9cfNlCK
OjvduMcZeHkP8GpkJNCUhAPOiwqI5nOQ81BE4CGP/rU9YOEVXK4lpnOhRMg+Wsy5
vKjPGEHFKbICywz6HvG6QFfZfuPAZ5QFlCuRSOtRDsMVHONKRz6Y/TTTMdXOQZ0C
ojKF5Gdb3bewhine9SVbjYNKMCWOQtWG6GfAv7Vh+bqa/6/9h9TfTu4Qj6rxmxB5
lkxaaoJbXlBJVOXuc59l3sR3YLbI9v9y/twctopycX3dqbvcIMLkOVsNNh2GdYVj
OCHD5Hswci+fyUSgC3CFEtELaOrAd3d0BVnxEwfR4HyhDe10BwqCbj8TD3+f5MLx
Y1GcnpjxDilHdNEbJURiNVha7Wg9n5F7sh2z+lMy229tulDN7qYIUaE+KwsALzLO
Q3qjWaFFw1OZ8XsHiWa2KnaSx4JlBlY+6ZhBnwHCa98yEiJ2uvbNC1txSktuWXnq
4LgO6lXsHImWznq10ODdxxN8BAjwajSuk0crEubHFwktDAhOeHTo5XL0up1EVtzq
QrlqeOjNUiLeUPzntd7Sdimy/0iDESijefQ6YbBZ068scf1o3Gmq0IZVfrfUDPl4
UJQwJzGTMklbIOIFpzQ1b4YW4Bje5JoJ6dwRJRQaFeUix0Cu9FMCnRbEvUqJ7buL
wg19w6ne6MYWgCtejCdqUKzaqtzZpLhviV82ijZ8cSJ6lECUUzzNcvt1JUfl7xyd
T5vDcp/66QQCVFkFndhsj1j7ygm4o6vXKIuxQEU10f+KAno40FZejZW9rk6QNqWW
9WFVlMqrOERRdPQDfjtR8tGJe0JcWzWbXQKr5Z3IUGglKJgPytFjPDwzFEHYuhHy
Hw8dBGAJG2AB7k42pr3N7xzkEtqLdQpQ0eroCi7I08jxnH9MFdwDxYuMEpE9CwX1
obbviLUgbrutp7aY6UHvXJWtkh+rM9IGiXqwzidrpD/fsG69m+IG1vt3ToB22Zkl
U2S1CmfxFhWZUOlPq4H95+Hgt0GaoByZrul3UK342BPJLPjIftm9QYXNd7EEM/Dm
79Z+zMSsHN4enxyVoE2wPvLFSxJ5Vsz8q/8u/BIIs2AvEk/Dze27PKfBcny9u6ER
hGyrSWc+b/UQFakE4rZbQhuraa4O1GrZ44x7I/3E6NQSb8QP8S+7WUAS3jub4Lxw
5LDKNSJ3RMmafZ1eDd8gGUMUiLbA0FVsokVMho1wB6kLQtYF50Ua5ugfP6H80ubW
RfDiq1K9Biw7H3RRzFJAVsGbNGNWWkL8u52kLpDnwa5wtmCI6lqvkOTnJwfYb1gk
nz9dinTOR9KdJtoJSTYf+lQ+1fh7PnFmSs7PeD8aV1IBrXynykyGU8IEuizqHMKh
60AcvmgYWbIGFG+gyZqnwcNFgj21jn6D4iDeMIXWgoaTwpTgcaSW2mjnUo9lSIsD
mriaxjd63vstOofMqiVIcf0d8tdT48noIfWR9s5Prmh73Y1VumdakJSCM25DHm3y
hj11fK6pWuoO3gTYCmNLDu9YvHcOOlEYSNRHZY8/GpPCFYxJ8r3Jl3EFn1oddVoV
Y1hEp9r+HNVX+CYbsV0HHGh8UFdlA1JhZi1fn9VTAkUodM0XJ2bpeetMXbNc97tC
V+hf9xMLFlVHGhULjQz5XJvKXuJdybaZymYrntxi8WGZ+GBrD1+E51rjzMc6xaZA
nrC1L/V569yqtpNDVt6lV7P+wROnJuRRJgaVnRvKcTcD0IKeRTZMd4XHPO5Kn7tm
djc/YFXNS99vBIc7LPB9v70ztRaZ/Pgtbz5RiNMzjQtKGNq0qg0I4UnznZKihJ/H
0Z1E2bvAzhiYAxYE01qhvn/a0vFHpFEeEDDcRXQPPDJTijGePV70TM4VEHYkximY
O+G0TiroslyChShDK0kGdM+uYnz63ooKh2HyNw8bso0GeZN9GE/wa2lO3Zhlew3S
L6sHimgEg3NnvGlehFeF8ZXcSiguq9QDAIERFYbt+fsKuZAtupE7P9AuI4ScaDRC
5L+bLwQ5DDOdECcAo5fyRhitJOR7SpmGMsy1ZGJXbWlXMOxQ2baLbCXslsJ1/b8L
2C0n1leWfPfIF+NLg4XoNU6hKkmZ3MTyCbvTZeKBgbIvoqVsMqFObNH3WKCtFuBN
hnweDit24SP4LkpHqoRipEvNmSgx9XVM/IbF9uNicFPVTm4TDaz2C6yJ0TqmcijU
ggUjWu12WALKKTphjC+cEAAK+epvOucVTCgZx8DUq/85zR7r6TenVGJF1OyEZTl7
yP2WVyqAoVMfwZaHnpw5GjI6Duyf9hFqYNUP0IRshdNg9sOHRP7NKhZ29sRvo5bv
7BD/6Va8/6kGxYfyTaqN+vA+EVnWgnWYpEJFTuBpIXAvnBd3tA35epJ7BCltVLJi
Oau+633+R7HwidhGoNmeJ8NPDTlu7uQanl2E6r8Xmevt4SbhK6Suibu728ooLt8C
+INBd5eOZkmh/P4L0Yak2Z2oZRvk28ZqhEa2xQtOa2hx8L1nbEtL5ceI0Eh/2zS6
6yqzdOeeTAWyuDBdo9boVC5LqXRy398l6LXFRyDmfAz1VoQx0joljNISLdegJcX3
ykGwZonHmrOMsJP6TjbQRKTfVd8BBuszhG1pDXa7zpoxX+osZBRLw+VXyHgZC58v
nXnN4Qq3Ks1hvij23nejzoYdkIyXnFftwkp2KysMGgNGJQjz6M36+jQZrgFEIpo6
IKtG7l5a53OCfkIw/is27XpbJxjG47x7OxZXKdzK4eHneZ0ERTqiwePk1suHk+GT
uOIgHtnUkPhO0rXJyiSbwOPRkh7BNYTscAVzihipAI6Cpe4OLhJVvBc/Rvrz3a2A
0l5ZpdKL1sMO2MOE1eZojPi9nYoBjGv+mgGGDJnx0aZmPQZLw5YE8W9vEObJ+FEa
kpC7T5LGwdJMSX/WFb2GBq0TDUZ8TZ2x9BEHpAUfySTrxifyJdvvDquNaDERQd8N
XLNWCbpqU8WOHHXhAOZ/aHE+oeEusj29Ro6MGmz7/vc3LH8KzoeaK6Cyfp80bhG8
kekuH0unYjbz8BFGTt3pWmv8y0aiZe2DowFlKrkT+pt5jX10SutVWsorWMM/WERl
wn5qp3NethKRVv3sX1ZrvQ3r+gN63TO+vEaBgu8LeIZyFwleTPf19FODHOGNOIne
z53nqA4U2d2IpYEf3avOW5ByzLuGO1Lmvi9o5DsSZVsrcPeMpuQWZaGqSFTG0ZGr
whwJ+fcFHwdAsc5FOtx++01GGxqSKgeSE77g5ofSJHL0KINODSl0d2IGyCcYm5ar
CSmLU2+tZOAnQ0RYCvwVocYrd0b7IOf9pau0QYuaoXKmAYYkaAiOgYib9LnLOTkl
joXwIYbHBZUETJKMhS2HSAr6NnlpBqBwT5mvaunqntT+/5VeWILkYIUw+ML1vpsu
96KCqR0f0OEcr9LBmkJ9cM+SmM/jdGVY03NW1CtIuCzpU04EngQnQDrnXB7uwDKh
MOy0wCwPSEaW3rOgdRAWaQWI5wINvFQ5psbrhYdn0H/fMJQq7plKNP5h+BEwiKCm
8ab8EJXEPxU7lrar+rvTNSZDqHp10WtT1LZme0MbW+tvGiTA+eOJw2lllITCAEh7
Bu5ZsU0Dl7Kw/nFgE7maG6IzqoctdcD024jWokGtx0Bd+Tcmd/d9jWf5V04lT1cG
8+pIZ34sdp3RxE6KyZdMo09MRzgoHq3C9bCS4jh51n2e7IzA7oMr5CcoNF8SZTQT
DU9vG12jt/ye8upeAfZLx4bkYBovUQncPOJqXlMKwMCDw4zdX5whY/HoixpB1kLC
vT4RHVcFQfWICpze2Ts/GoEIXdDFYt2KiY5av9JJ0N4ma7+8MkXwHfYWOAACnDkw
Yg3fiGqprnH4F/02VBuxp0CGtqMtxAEhJ48C2B0RcUJRXIztAaTb+ZOWNx3czyXX
mOmTSc3upbzy3e6SAxOJF8iAz1iuEIBk4T6n1RGbh6b9EfV46/T/nY1gthv7DaaK
b/v5a4KBuLbW50/fAGBmiq1IWmE15k5Q8hMqC35xKh4tjeyGQAgOF2Ck7kXaCzkZ
9DvUks/6QqRXU0+0JDOB69HeAZMxaU5ebhuf4y+Vc/TKH8+kXsAPe8DGUZg6kEmF
O393DZS5DahAEnfzaSt4TfL2kgqh2HJbAl+2R9/wrDHuIZDHvmoT5sMvtqaepKyt
IqjstigulAnDghY8Y8PsFvNIaaFQWt2RgCCiNQectu1bjmSNArD0U5irpLS2HQ4m
rq9oUts45YFHsuhyNR7WgbpdoMlGI3smwmBlUbtV0tlBjDzkm/O6DEq0KZ1atM6E
3YRrapFlrkLe+Ec/Jp/De6AMPJGDj53Xn4PGErtH/ZKivPG4Wa57Vjpwnx+SBze/
jPNfQzmmdQxGh5+fD8ZZ2fD1vuInMAR/uRovS35KzzJOYWWhsZbT4rbpGybWT8Fc
ojeBPwizoMKpAdmEOh9rcDKvVaADiFq/WbYHBaC9ZENSM7j5sSew0OAaK2jWGM/O
sYrxiQenhTVf8KJYwih/YRo2mrfyRhLCwEPjyZPfbZBhGdnJ3dXq0xXDN1wwWK6T
d6bxBVuUBkKe4ODe82gSzf8sI/G0hzHZ1s8jOxPYth8XBdirZRc5o3fTzq6JclNZ
Cs8sPW1XKNjIIMRNpO+Rp3/WIg2S+zS3NwxGiXIIZWNSq/ZeCH1FykurSeM7pv9/
zzKyM+NWTGrPOPlE5XYw1CDbm/zAoI/TayBpk0hx0yxYbLff2I/K9nGjzNyPjKb2
NUG57UO28lfVSqjtddGaPiVaqIu6KMmsBgCEjsfzyw+VYX3BCTNVt0EKXVhEVAUj
qQkna/nuti6tiesU14UcXMkN48oLJX4c0D01As9o3eeRuccoSCSkpUXbW3UnO9/l
s4vfx4PUo9MnGiG3bm+QkhuRyRYAeWTyAO4ZDGM8+1Qfpue0jIp2NyvkAV1maPox
+d5joeKtu5ks5Y8f77+2HW5gkKCMJXt1cwSEEW/2vNinneirVZ5LUjTnmP4azSfp
CYh5FA3dkIsDUKQOqWk8yFMJ2+Y2din8nv0l4JIYvoDvur/5XKLnIhhR7iBMIxRM
4pcQCocaQf89MyIFETJ95jBoeiJf7qs6aM1NE/g/0RqhEYs219vttS1dq4lojijA
AthnGSyaPATiybQtBtpmvCelXVS7BKmPywzs9rY7PQmixt62k4t4nAB8UoRSRZ1s
k5ig1hcWWeeXVbw1flYsyoZuO6tGQDhOdBo8BqHOaFBR2ecbyRMcDe082swQcSUH
xsIpGVjnuYtqatCHcj5lwyog5Z8+zlX8Hzuvyq6zjDnlZb3/xPUM5FWInVnSL7t5
rOvpQbieNsdbbvDHp0yLTVqslye3emQAQqGNQ7s7lIcMwh0isrklblsOx4DOJ3mO
ndO8cNtIH0vjLTfcAztRByLFkv+59iXzVD49knoE+c3JE+BB71RBJaxbE6dqGYac
ONQayOKQkmjmpK1JXy9DA1OM7kQno+9JrEAkom42ae5NBWvqJAEUX8MqwwAMYRR8
+2kezzlaeAKeLdMtgjlXc+cQ2nE/qNQrtkBQIaDhUnDbpzNV4ZJL1Q3cVuB+Nu4w
AgNK4sSaNUkZoEL7OqQFr5DRiEWo0cSlf0Gc57v1dTkvzdGwo6OkE8vcnLKomkQ8
x4IgxwkS3b5D7PjQ6s/s2oIwW4n/DHEgJFiwMvjtfmyhGxbSHEi+s7ENN+7792bH
2O8GuZb12eUx5j8M0A1qSzkwApTfzvXe/yatlpF1xpMi09SWS4QS89Pq8LIAa3OV
KIyGMF8MOGWwZu2/gPRnmDEPsh6Eowbb63NT+bpjsFpsV2Ot6wXK404rBgkZ2Cuq
aZd8xuHv5J7xL5Iu6UEuDN0jwYsmTTHyxizFFwh+ejiNxzkFQlib/CN00Y5jWb57
lOmHgbaFqADsOXMjZeuk2r4eA1FxCH5DlwF7hBmqBnKHtB4zwJGyaBycrs5Uor4i
7sdlDgM5WrqkdhkoATLVRhEwD6KJiV2u9+b8wAHGSx/ctDoOoE6N8+xgZZtU71v2
7O3XdEQrLfuR/AXPq8Rj0rOVb9v9N2MGIQZEWDw850jXFqJVMCa7yi3B6IXRJzGP
ExGvIFZ/3JQjQRcFVgyp3/b48HBWj2J0caT7r6RWdtr4sod3OSNVfwJKKnSLm5kg
yEqTJ2xifH23pSTGGkErnYn9Ni0CtV7Bs63IauOF6NRMWUMoj6DxMw/vXX6qs2U9
9fInLJlcrpD5ouHJGtTBWuVq/YLOpLFSuwI6AZfweZuT4jQhK6T98zabPpX2+zo4
N6wJz/JYc7ZSstPcCgQnhSf/3CCgykAa6KdBYAfilLCMuPfqMp8yowhy9yZVb11e
QhskAFoQgZe3zSXznOAgkycYLXg/yhdjlOSCxUbWDU2risP/ncTf3kg5O5jnLL+u
usktGBnICKGnqBpIKa7403zBdo4g8lTsxzXHedwT+XMOrUid1jZH92O/DJptJG9d
vPFZyjoctLZSu3y9y0EH5PHN4j0Urs49F7jKdeVy3Z25mZxUjtq3AFGNKBonJqUH
ew4Bp4ylIyDKZ20ujQVHXrTsJRDxqrPvAoTIqsxsyaz8sZFFBMmA8UtOaWTjDY+L
tfeB6FNNfsowNtRc9Gd4JZv/xKWDcre2HO4Jcn6Kmavb4zT7CRTw4buOWTetVMiM
gw9yG9mrmJRYbIy4MEAO5BauM6THMfGi6yponc9p/HsWHWiemZDGahxPxQ8lD6jw
9bC3hevXYGJ4bp4GwI6/NzAjtmYOBcZlyTm3Nf6bMeXQZJKl496/rPmKjIyAEUxU
Cgps7zLCMcgVkyclW31uHv2QaDhBqyeJD/dNsAM8srpcro2ENA/OKcFC7XZh4BLy
nEvg3JoBdH0l+H/i0/sQT79Ul6irom4goxQ9jNe2vJzf15Sp51FqUBGZXVEBk8hs
15/BbYSbLyiWXOeFqRxhWTGTRwiqXdlFVZyB2O7ihyGePP/glHi/CDNgWaVJ54+6
4crjyqFfkiF7RhGN+eI+UMZnKg74EgoCvlFmp2vgEN9ogp/Oae98vDg5NEx4wwc2
+fp7hfWB2WyM/krp3RKyfuEg1hI7vof8CEBSUuJ5RhCC7YIzLZI2aZnnakABNGCD
m/V1/qdo5WlPbdQtIfnyJ6By7VFcmM48exHa3X6H84Unw1PAXQzqnIGBKHldaHDz
QcYsqaM+wj3OAJU6Mf+zmB/B3cgcjsdnRpUVpvlXhn0TiHbrTAAWB+coUWPgC4cv
1DLfh+fCXHkQUQcIo5oxgur27nGziRKztWBVErW6hgTrs2T1HDQh57IvKz9p1s54
8nUrZxC9sDHJFm8VCllxADZsxwVxrjLh1FhVUh1b8N3XhcHXBD+YzkxeSxzOIadO
wqjoP025DdZymX1360ZgHclSa69CX3KHZ6s8ZqSrhrbBRrlODRE1aRNT4zRKUvfZ
n1J2uMXUSwsRLf6oWvklGDOlilTtPfYBnHvyMaosAOoBN8aDRo1le1beC7kZXn2n
MTftRHOL9egHIAAGmpwIERM3tMWFjVGpKNCesG3ZuLgFirLLA9huxPcbOLfKId8m
5WVaWytCng/RApMvD4JDXKF9uU65oLFZv3xR02xJhuKeMFQ2kMXYaWqU+lQH+E13
69crbBxutK8PCgaTpjQVNqNvCaFlySTtHEx+O+1DcoDhpING+sYU6L+Ae3NC66Xx
TK1gasw/yoNdAmS3DUNgJgYuGPN0OlpIjE2rKMScr+FRFVVYSse4H8NPskShgGJz
Ig9ah8DbdSpnE+kkkP8ZHkoYhepmRwK82satPRLJ4C3R4VtIfhJ27dvy1YbnynfY
BAM37zlQjHfjCOthY5zRxfO9oLEqHYlNolC7OMhGI9Gn6fWGadnkur5y3yvb2cIS
AB2olXLmSdlrKYc3tKIKmZLHZp2w5r5qcinicW978W+1V1+7/vWWidjZtbsOYutd
3iT9uLu8JKCun4zaXvySFGzUYvC5qJF9QC0Z/Ijoq7DfR5lZF9oHhJKSUvrNa/Yi
G8AVxVcxii3Bc54kM7khEZCeHrGb7BRMW8K+g5UGb2ykkLtUQjb/Pony8NH0L9MU
TJfpeTEDZ5EM2x1oPfLG/6P7dZj7s9uk6KLvAfU6R/hetpvd4kLuBsfEY3AV3Xl0
TlYceAUtknvR8eK+daSC2sRKOLj2jlHvtvo3uurl2+dRpENDUR+CGR6AD0K1gHwS
fk+/a3EMesTsSg9PSjmqgWegU96UZOVTc4paaVNjNw/qMfkt+LT25YREFqph4CVd
Om1VYrOsDbogMvITYSJ0bTepKPJRoPfJfIthSeqMJo14+DxKUODPYpKoAujwuMNL
pk9465f9Vvegl1olajGxFjUkQ+R4ks6svQXV1nqqn2CNrNoRxtx6hdkmDL1V7/p5
jQypMqeS5YLR4c4+zZ3bVHy4ZWl2YU28d1xR7nG4Z6TUA6zKph+nI+gy2lJYRL7t
aYxpA1h0tJfCKw4bpQUuayiUQceXYIm5P7QJTDCygk2ZvCEMf0eycsPdRpHfpDPs
HiFBfT06G2HWBwZiBr/V/r3pEtt/gAs4RTBIaXMKWQhr5RJaeM88N0GliYiWhJMV
TPJuZ8GsSclVqFsmk4pRtE0Oj9cNGbS16mreun5ytTWz5bYQksHSXwfaDsrxhQpE
cNSDdWA5yVCwpK8l22s/+5dIjVHW+VTnDPFv8uv0e7PhVtBOAOCC9S8efTOlDGEo
lRHaYcvPyFfPEYJyN9V/3gdYfA2aT1KVzUThIKIQ4HYoyQbuaQDWbPd/pDpklsgn
MTuelS+RzKTQ9JFw8BePRu2T1cuJiSyUQ363BnYPnkDDdqRaAo+rx1jiKp27X8ZE
0cIp9HBxuYQmtxS37h6qhnYFObdk0ptgJQSObgGrwQmhSJ+vQpHmdCFYbQz+e/wG
/dEjf8JFrjeuA6W/cxGb+RPE+kB5plKDKcrnru8wptwT2ZgDdaU6O1WOYXIM+nqw
zCNeaRRS0tx6Q03E4t0s1P9to8UjmpZ2Zw+28uEVAUq8rtLSXnXATA9Fu0WIC+7q
weGqaByBqbZYmg9n+SaAPbHxKPBaDMpCptJI6dwL8+52c9qhEE7PIIqd32FHcVQ+
JF4hJaeex6IxAjUNdpDTKVc/9cvb3ZARSmckQvMaxZFUdu0vpMgr2hSt9e7LTWhl
+qfuiBl2rNY9z1YwgB8N8OOJGHF55eZVLkAn5MA5zTT5dhgfO9KeG4W6il/SZhR7
SCmCb0/HqqZbzsQRkw7BCTcSN86TQEuq58dEf4Znlm3cCxX4wyz05MR8DJLgyRRT
lsAmwdRsEHea9k9ey6oT74XlrBkXgFhr5/OJ7dTXr1q08lK1GyqnzBCAR2hb/emb
ovWJsWb/MyI8nnGX9y6VpeLZwEd0V31AwalI60L4/hlrobdGz2dMd04KexRIAH8W
LriNqwJUIQG1XEnUpSlkwmX5Iz8jLuiCcgGbuM+uikmlOnfok/CwdyXqKVG9n+q5
g816qWjYzxpDdcSN8ibPz0El0jTjAeFAJ86Sk+W5oVN+2m1r0z+dbZWHTUUw8ya+
rSC1c015DQCIMWFsqpZK5jCPY5ilRXm4uTtbbHx915gOpwPwHccIcY/hLOrSnibp
z3Fb0jVhgGj1Gw682mDHsfojRxQcsRj/EjiELbxyXjvIm4shmEMDW8Wdv3jmXdrU
gJ8doMO0nnMO/VaJDQMI/SbPvqbGR970VIh8Ena5l4zGILzpwBwldjlc4EaZGgle
8Wt2UmN0MyXf204Dqk+UlWgsyjoU+eR4ePO4s6COqnpugTcyKMM2o23Z10bcOjRm
kxrJz9u3N6W1F/WV1FUSjoyEMFn378J4g0jM9buWPV4AnfpTGvcpNnNoeTDyvREf
HhAkP8gMaO6suaeWhvv+ZvDedwUwlS81x0dvMiACsQPnXlWInLN2e7h8JuHIzG6m
ndeiY91rJgypplWke7oONksFPg4qTCCNKgIV1yX716/Ai47Wy3N1yN7OCTNSUu2y
POwCBdYDSesW7fyST7HkVBvwKkZa0HfrEwtPg9DJAKxlBbk4V74Gm7kGsB+ZC7TG
sHfa6dw6wLBKLLHO/yWnF/26omHmbHijRGzrWj3XMPOX3mYh5GyFl4GRpmxHo7eR
0oj6SqzNiwoICnQWO/jK2i6U/9ljTQuH4S5FxANPy4SVDVpOSTvmMmoGvG7Cbi20
0an6VIWylFwxoV6XpaW8e0CZZ7x9sdgba4VlMU2+c5kSANnD5RxZTLwX+3kkBNU9
rSl85JM+b/XwTLDdd3mW1C8D13loeTw/XkpyoLaWjIez1hwNs/Hux78QhZaEJyf+
902cPozT3/8mYTQ5ulzMLkEBpqtmAPyikdbZsafi+QColJsL+GgXJTU2HsCPGj8X
LPtIpIg5VSV/+X2SJkeI0cZtgmUI1XFFun7yI5ok6g91kU/WPdxsQbZ/Asw1gUfL
80jLF1jivEAr+ZhwTB94H25TbyZC3DzY36G5anzbyVsmo5TQXIn06djbOoj0Sm3n
a6VSicnyCONdelHZr78KTTowayV0XpI46CWQCDnn4HQXxgTmV+HAT7lJ+PIk+nl2
xvBng92QwuSBLvQaitgu2YflsakvKafLY84MuXryOrDxeaEIRMth+sQzm4K7bAKE
twEjHOjST3JRK3oJaMPUploRYelp4aFcVQC6GT5mzBOODx/SCdfUmay+XLBdPNUv
ukM56kKgpQNIwyiitF586QlRlBpSSlyRbDDFGb13hO4eScM1aoynpznSDCy0fSo9
hGfTEYcHiPvlJV9+9MhY3O22enpOaN4O6dHYRedDtfvuCga2rEqh6MoNUUJWKbPm
9EKHcpZjz+cfzMnyqc4Ydq96gROCN7Hg8bqMqATHS8tyDxvbycIkjCj1kWw/4da2
yFfXhIR8+8GUyskhoV+xij4FxSiVSQc7h6QzrYO3DNE=
`pragma protect end_protected
