// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:35:36 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
PgMCqVjcYAaMn/Up4j4Y6MTVh9Cf0EAdhpii2InleQxVYEoPTb3SWRc27XoFcPK5
BiJL+o0IH2QQfEqMsHFm9Xm5ijPbr8OcH+0oWvQ9/denAhawAtg0uYcyu1Z3ZQm3
ZdL9U6JCEePcO3eZg4CjAxG0bWHddBTLVU+RujOKDYw=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 7568)
L3o96/ubsx2MHXO2v0q8pTgd9Ff7NEGoyS7P6sY047qMY5JpY95d7rksNpJHNGt0
M0mzgfPoRKg305bIFZhtROEeA38pieEKLATcJ2KD//vv8YAqts/HrKvKIwvLb9XG
4AGiuHKjNGFSlW09f8xys/PNMX+dE0O4nuZBrBZNca9HP7cifiRZBPKdWekugQx8
S5tITbHODvfWt8j1dyQ5yBKIcgjJUMbeH5JglWhHoxmygVx74jh7j8jgEEHTzaYI
5Vk+/bSoXxn1zGiT6zEKOTMaxrD0XcyIh51aojTC0ygNUJ8jmM+OuQv3v5Jhce2z
8OcXph7aygXfi+RwL6dTduy1te3XUxLhvMd05hy7jWVWAT+SpK+QbcBhSTYtxyL0
nZBiExp6S37ioruuJ2bvCoEjEJUfnBjlb5HT1peBteieZ0HGLvbP0hcfHstYX+n6
BPOMuyuEkQazE39qTReE0eoS3Mf64CrhhfutqxO0QBIttM5FjxpnLSvyACTInPMN
Hdgvca0ieXnFHr6Y1vNy72BDHLjL/e1/IW3PzOy7eg2+ilsAA/EezN4eNFjbXtmo
ukK4iq91xIljktXFPYoHMy2MoO60QC568uRr6V5Ks7h2KflgHGwvi4aWXGJ7ZI91
TbLOHgX91f0TJSK1wGw4etNEygRduGqHPlQv6hd+YA/o7XW5PcGTeRQfUq9yYqfn
UOOySGfPJlJ7xQEO5CSd1nUVrE8TTeruQ/3iULkLznF79lzxGzOC9SmGi5y19IFd
6ocj9hyRJp8g0v65CoKCBtvXIIU5hG+3EbnFogK78ZguQqgMP4jTjJIm4yPBqwDt
MbiTuVq78y+L9KZ/+H7/bB44Bz77QbgSEvLafJAeA8IYNk3+s1Q2z7UPY0uQoo4M
Pbs26v+uls3TBgCxPLyUCXB6GOhvSrIIu7l4qE5coJPIoEntJ9cTwZPLmmgglexF
IHuQv5ERZ0vqZLYcQDVK+iA/f4iUFx4Ex+74beAwBJKNeX/ng4eFRZqSMIb1/Jjp
/8HEWrILivynM6OSfdLODRQvp1NSlSuc6J9r10VQQ/XSL4jakOzPJ7Z5XOPIptex
nsy5a+7C8kCSRBXMTC1Ndtr0wUTXVcqbUjL2B5fW2VbtHQhTPCAwlNu9mtOdLmxd
95HmauHqQpizgRdZTMfyZh2ibsXTBwwGV7kcGZ6+bzUi93EVfJEQ0HOPCHcIyTXa
uCFZkZcNYYbKpIUb7JxVLWlyMG/i80raPriIhueJ87p/Xcnhh+ILz+1poOm9Z7kZ
BJe+7TkXU8fHfqZTh8kVMWJujZXHjMOsNmnJuugjnQ69rgDCs6scwNsaf7xKR9W9
0sp0gkXCjB7OIbs37Xa0y3yWQ5q737wBy08OXtr8tPI9Y55ZpDaM3f7Mog6E3FBR
3chwdQmtrPqHN3pDWsE8ozJOcr92E6IICENpYC0y7bXVpJ4ZpL+ukVBmh202uESp
2KaNTmoMU1GR5+4W8N8arSZ7jJwfKXKcVeiT1bP4orYykY7787AAHnODxbv54mH5
/84TbeNuSXlHToAnb5V8wMnhwcj+EjlVClV4w4xvKaeUn7E7eH/6Hm15pqSrFZ/7
Kiqp5sZ5hi5e6srzzPOUh5/9K6q5L95eYUgvEMKl08g6ijSWOBOOC720OjNJCDWe
oUhzZETrl/PV4gM+FCLKqA4Rr4t49ws5/MGhtbyij2PRvmNioTVuRsdShY0r+dVM
w1II9GAsZyxRei/uwR2UUAIUstqd6g/zwXac8o/q3kha9Uexc8h50QcCxR/LUQXc
DgWIzeegIMuW/mS7soJPQnMjiWOnGHo+WCQOSRCQjpjDs0gAAF/jn/wx/vXOYFX8
z1U9j2hP3u3eEfYS68ozvve/k8aj2layE+uf8zEBf35HwZkSeLIZLnYRQ16YLTnS
Q20ooM12Dn+hSA9Mr/fN2wYMNYq9PqMkG9NnZz5/4kDHEzhE6o03v5cpgxoNF9cD
eTr0Y09s+giEaItkQdX1znYOhlLRXFRtdnI/TpVi4Wg5rPR3fbU3za8gyWuAbX17
umcbfvw3KIquBFUqdzgF9lR2WWnf6MFScTh7h8rmkea1Fm8Q75TPN6APYyKaRBh6
McVRDd3HEtxnh4Nu3bm1sYCx7pBHpdLgrEr5i9hNjdJRZnYYSfyTAaDuXq1AzEVS
snUwCjYYSL3fFX31wyhnzvupoinfHKzJx1Fmw9rsSuyk7bvQG81ZyfmfS5JOwDwv
s+KM2EXHcy2BokrgxbKG2wiLREo3YofIdOu0lTFmCt6d5LFwdgfB2h1vuDsgrVf3
TWUtMOEy4mVKU1q+6py/mE/U3iCwIty13/nilKU0HWxn0+dGLWDgWVrdstjJJkms
DpXildO76b+E+2HO1w9HZq1NcISZ6JUIuGyoEOH+N4f2WfQuaYJyqZSz2EoPKHtZ
vAIKz6WTPkcZCU3VYJcaoEiue/yELP358KL6P2wh1vsdZ6T5oM1eV4cLFaR14x/c
AfTnqNPI/PTJ68MtEqFIn//k+NZ6spQ4T6fnihL2LtiSpxyzDrANzW0H0AZ9UbPc
2LW7tWIwlKCehad3Triy366gKinFKV7uqe1t/3qQHPV3QcobVHeBcnPtO73eAgU4
nXj5gtRG4Jk1QvxHvwdk5OqZlBSCUrpGdd6BYdC44E12ammwD0e3zmEfb1s2JjH6
ddRYXky5e7RY1Fc5dc0hVa8OKg12NkWNWngLpku+gMgknshMZwI4YzLmbadyMOHN
N++HAbpkrQCZagauSnd/Uuu0bepM7uQAqlkl/Ici42U2bjx0FWvliGB/ViPBK09G
bm6G/YzMQum9j1kcY5hcqN3tDIc3GinTmI2XYHHWOwfRthxQ7Nv0GsdNge3Dv9vm
t9A4F0KvpC2YGqbjzbc/ZMv78WKYgnIZel+pMMJlq6EuvmkwjsdTYpRCzv4+cDxU
hGb5/cEdUhrZheqjzYqxArSNpYaQ2IJaGM5c27F00apTDoQSSvSN7Kz3fBg62iiu
yk0P3M8jKiYAf6R7gQUq6tqqf+XK6i2JwZswP40edn8PG9e/A/VEhPpiH9EbT739
XvyW6XPwid5PHOIlPVeteeF+pvBKgRo8hzLDjI6q3fv+FCjYST2+2hFippLSWkl/
2EC3vZCY4Astjq5cbOhcDwo2S8fd4vlAhMpcuwXfxburnIFnKBPkZwUv5+0P0ypF
7NVPHIAI6NL0SniLuSycUCEZZ17bRXisN3K5MZJolWc7ZIj9Z7sZ9MC32pMWvqvu
qb1DlycEQ4oByZHeK1MRHGq3j7VVBWdicFHJ1fz/DEmd3hDOuZPX20SvM5iqvqnx
LjskingQf5lkcwrDUfpJZp9QrLrCCnDyFbwR0YWxAA8kAr68e8HjoJjK54so/P9o
uQM79VaBha6BXAvQhMG9Gvn320GTmMtY1PTmRUFdP+y+mPAUW3ftbBvA9Tu3+CWh
0EPB8oMWQGrhVqjWYh/vAIx6n9HuKbQCzDkNTmeokVnW/wvPZxvXLmpIqTGU6Zi0
KeemGG8Fl366+JMm7P+Ol0hYI9sauou5M8RlBvXZVtMhbCJ3H2ci+yW+1VMQVQce
pCIuR3AOuBj0smqyZkB+c8mfD2vAW1AAhiOYf+ZHXPN3KuAWn6FB4JMx7hAH5BdW
mwT7wBchrjATWvfk0ud/4DX0vHyBZJksn8IvQ5E3NHxkhaHQFTly5gAEh4nyAzu4
eXDY5Yog4PFZmVTb2YwI0KzFPEJ1IW0f+NDgxL4fw1wuJvcwYW6qtFrOEXiF9OZm
8wJ3sBDGRARC58epLAIb+0FCGZEcdIH85cMMoNFZWIvP5cLcSnvRyjvg8PPuLjCQ
adoQU72UDK7MZQHo05Yp01tfCaaQyKi7Iop2CnWeIxTFsfzjpwgs88aBdnM+LRiN
omRzdR7FMC3vvRv96rh8m8TFoeM50AjuC5G5q1Ve3wnl2ck32ddiD1gUUp1/GepU
Z89X5dVzf/o37b6gMMwt1AU/zofNCv0iDIt11pgbsPmVJMC5FoVMsmRaY2uMxOXl
L/FRO8EYxbGdDi5Zc6SUn2DvkX63Pu/7GswHhyeQQ5SN7Wr/Ak0Ob971zIONb1SK
WYKxiCvQelp/+WhCdAGzMQDyZgbmagFx7h3yrG2KWwRDbWad2XlGFdC+A5IhyoAm
8s6uDa9Roo97014Qy1C33i5xTOADr0MITEcNVCPDAF+tHC6gtqztIwIOiB2HnIjR
WhbroJDbr92m7VanHOSz5jP6A4hDjtBVWO35l2Ao7s0i8ANa6y0w7VL1BKNWLFcE
aV2rPTJ8w9bplQVkam/oZWxx8N40jfg7dETSFqc/9aDb/qyULc5y2UXBLqyD1EMK
TXqsZ+OjRpWvPdfffQ6aGQW9oESjLMUUHQx62HTK6e87u7K/ovm/cXrtTkMiGG9V
SaLiYZIYYMfNyzlOxoysXhWypQ/lQHTb8rUoYvZCWs8Pe7GxOUZS5JVBXIwcKf0z
8nXb6rhRVPdjx4i1cuOEd4VnFxrmAztEcLwQCxPavsMe5NsBpMidfGEduoOXROIp
4SGYWNJ3StdGLrWcUA/1Ub8JPyFWjev98PhzvUA0ng0dKfCyqRZOjrKDakuv3sd8
gxXsyPaliof+JqH3W4bbZsY2+mCdRchzZ9UdaMBtJYsaWxR+E/ZshgYPjxJ1NprT
rLxri+zqptnKIE8rdbx/KdJWZJE6esKCErIxRwROwJICglRyMO4GXin9rX/ZYWLa
vmmwVrkW+8jl/EB/SCSkmrcffC8aG/Gd6L1COXtlgtwvQz2XcA4KSBtRSehsFrqG
nsnYf8W33CqYwRTfE/zXWSedk1NwfrX7ybDETf2Zv+iXftGQxZ7tfUnH2EtlJXBq
qNz9ZqDJ006Qsg1BU0bAx+S+rX/J9hMoaaAIGNqCk52I5ut/oOkzsFvRVwuiGrDP
1h2vL5DiakvMHR9G8R5xOf5nJgnx0b9E3XAcQaZm9IcBNY2vpEkqKGM2jkpt2vNL
SwZuQ5c4bMWaIHt26se6OqnAaY4/41sJ3nioN+lAIeR4D6xuIdI2ljDGdBNNjUIE
pUaAWczSpBPJU9ZxYWfhDDOKCDolz98MkBs2JEqM6Sp+j+Bz3pCxN7WBO1ITPHWL
obA4+CDBenWKfD4EhNDvoqqsX4u0InER/9bRijXfbpWxQPAirVYumDmMizVephrG
RnHVOvF1T0zR3Np5AFi2PgHczGVek/JCT4mOh1AMFvjptEa9PilGG0uaJv8b0ilG
2o6LM5/t9itg1VzeE214amsIM0bSg9uUVAccAAqgfF1UDqLiPJ6OHYOcjuAL03tV
BpKcP5uTjaPriAUgEJusQ/DA1h3/6gb4n7DSkHa3AfaPaufWazwiCfrt6B9HWzca
X3cj8EvdVz2uxSjxQJuhJL71+3HBq/GBp16DY/YE704n82onOrYWZvKE0/DjirZy
hE07/X8cmX05uXQCMK/TSdJtygjmESez7F+Ue1jPlkn8vSJXtljb9kSFC2BaQHqF
qCD/RbDbNqejZoCsGWPG6EJn52RZ5EwNPw4tt2Y5/B8OZTZP18XnEVyPWftJ84g0
e28vLxaUS7pcEGke/ZtblOydlyhwQZhE7Jg3uEMbflT/ybo3iNezVB2IZWT2Auoz
b1MA2kIC8eUHRqbJEHtw+bTqdXYHBicGz14ZS9AXeP64lvKqXRCWJ7tqsSG1GmG7
If2bMgNO4pJYzh1hHX7tZotrkQ6vHVVZ7OoTytnuVLFUtYMGqGvDWyuAXhudpf15
fDvcNBfhUUmANW16f28z/tc9Cwsi63QWiVX5GMXY+JWLgKpChYV4sbU/zqpXfTFg
OvFNQrtONQmJki3VO2oKYdqPyeHnzfVFfLwK7Mes8BkAcLtbMil8n6AN2e7JniTZ
nVkc0nZkdgxs70RUvHT57A8z45TuQVnMNTtYX2oPdSl9AAZI5TNsoTu+0obd594X
RpbN+KIcpaLPqOAlrHs4S3gBlgd4KbGEQUnFtawGidxi+BoqwhZQc6f+gGdepS0a
OcOZPfNfleGb5VM5knQWn+d/JTaTmKzoGKbIF8FjRUsYI0HG9Gx5PVCaStqSSTRu
edBfQVFpyBcfTO/XG2FJ9Yc0IpRKOy4yUcCoDio2E2GZOCiMzGRJ23hdWqK1ssww
xy9YKkiff7cCBGjmkJyl306utjrQFgwhw5Njr/9CS5W+p1y6RkeIEkjxYyywHhCE
sbksVUJdwFzpZCVyqpIcso4uNhtCCm/TgPsyqJllXo9L5S+qffvYVif1Z5tf7pmw
xneJiFVrZHWJio2edV4GyVeOlDGxFaeclKgpnFY6LvPmranfQwwniTxy03u/sDW1
0cc1wqm9W6AdbhV4zUPvEs9XysK52w7JTk3vD/Vu3G2mTcK/WwGMyUR1fWwZBHu3
pVzca3uQBObl2oBK3gO9rV2eu6RRmR2y7B8leSWIs1WTNgIHxLRQW/Qbk4kX3z2z
aonhyfmwaUHfrKJPkpJmCOCzZTDAo0dA4Uya/goIP+eWLDF8XlxBW/S95TJP176R
xc2/GaDxfqATgHplz51dLJ1gfRwZvHqgTwt7FKLrLnyr/fUnBKE9hYXXdk0yZ+Eh
2O/Sw+nBdfxP/kDNuHJtreTWHr6tZ45DRugSZLSTt3p8z9JDiXblSDIqJJTmyFAa
WBq1WXqrTeeb17LICp0lVyR+4pAp520kbvVG784/lfkPZ5aLLvjoudeggCeJNA4y
q5b0X2iCrIQ84saJjFexZF0/+8cBvGCSF7EajT7M/EnU+yMfoIykbnLxsClLZtIk
x8PR2cX9u0KQr8ITAEIr5u2LbOMp6RJDNzUx80IWvGM10Q/mocA4mr9lQlO2vWnv
efefficDn6DpUpvYyUiHhcKSa57YVD4H/veqDCsYT7TVGNB0KVsbqf7b5bcbU+C4
KagX1GV5CCamm5XQkGFqddadVtp44BIu7Hk3Os+Fh1bztSMKoFO7EG/2uyzfKaz3
1n18kPP79e454NNl3uKLZth7feN4vE+eT9eN+sJscd/57D+w53Bca3X3xISeFimL
q2R9JrBLAJ1waVu5N2QVyU7lHJB1iodTMWab1XJngCdWf9w+FlSeKZOSonWWyY8C
ApiEaCBAPtSrmXxl1DcRaaL2ZOSMWX0SAGACuEcgLrTKDo5+CAy3DL6gShMH6t4v
LG4PyKQUloo8momCvZkunHvQBUTpYaQTjfDtZcK+Caql45ppGYyfW0vuLZbg/GyN
3VjXJSdF2su1G5VjIjDSsJSCtg4yAF6MMC2qsibam0pNJfPF6iIX+yaRZTKiJpUb
uWL3T+pzl5SvrCFgKLHxHpcyW96rtTuecyymC8hyVJvMnfR4Rg7shTMryWJdFGzh
eLkJH0iRzRiL5pYfdjryngLbGzKrC4hzg+dDiNRSKe2cM3Fl/xoh7CwxOdSdS8nf
LB8OaSL39wOkxYf+Pf/rzAUUL8vBLWt1a3qTgL6smUE+cNngUTI/ADJsfctwnG8Z
7AWphy8d8HHpWWQWR4VVsFrQzLdOaTsKEClAuorgLUWf75sLJoL4auBxMqujIQCI
FRuv6/Ib/pNLEUBwP3VcN39afR3U8pe5EcLxxsppwyMIixRlWWzoV4WbAYBmR4XZ
azQqGfoH0wZ7r3sd55rViC1cDr0uV7rWt5ecgGfLDZIWcS05zEIlVYCr1eQHImvR
D1gPHyKLDGjP4A8W18Wi2jC1/YhSIUqDoX1FH9sdi2fqGoSjsnC6yI984xJjZb7m
AmKvWlqQDhL/4YFMEzw9/UElZxZTARUujSp3biN40JC6Vw98XopYDbPnJY1OefY0
cgwtwxWs56GlJUD89LOphxIMwhr2jPc0YgthV/PPgj1Qna0wfgUgztcjDfO5VIt1
yZ5RThqIVQhN12LKi7v8LuChIfPD1j6YMXBDdWJOX4bAQCQQp/f/6PV4+eaVk+GT
Dvi7BGbh+PkSySOxH4GqRmi/63SNBYa7ptzBPMsT+o8MLTj5u+3i1JwOTSxsK1s7
TdwwPBpt7STp1HvMHNfNIE76WSuu+JnRkllM9QlM12zKiwU4c32JUfaoKlyzm+u7
MZvtQuxDswebJRUPnREFgeBa7q3xa5u2HfN2gawzw8U/691jcB+yMCcqV9A86X60
4I43OSMUH3JhDQkkbMVpVDw3b6n/8mc/6CaB9X0dDWq0vh1oHHUfoTFil6F4JjNC
Jc9nESmf3l03mpfv6h89BmloklrANCVd5i0bnHmkg6DSp45SvkqpyQwpc712LQ+G
IvrNYfC5MdQwteAd0KiNdLw1nPGKPxKBFrHHV1A0MWqAsndomDoW7rJe9fG0Zz0m
0QzQdkwlQO/UCtWUvbnqpErmABajU419cJANNE9KRQuIt9lA+PSk00scGPctaNUQ
8KGTM6hu0tpH4XC70qGkNjZSur/lIQd/Ce9DLNLJL6TIzGpOZaiwh7r9MBGDS0Wr
jGTT2JgBEWQPkgQ5ICNQs/fm4hjEcmepms/h2yUummuvZbUkdaULFMIIV8eGsrVy
zvHgxDJIK4gDu+CxXLb2p7MQFuzWOEYgdVw726lARvwj1NjGdjw0lOY6/TR/0qBC
E9Jf3GDEVDLW0ns77qY5TtdtO7bnp48rwR2z1WesTyS0HcSPMUQkzpQjZmVF6Dxg
w1f2V1+vghatdDLBAhnEuwxe6LmLcVhTgsrAjrFbHd63QGzHiTdNjFQpOaURaXbh
eB4nydMaonXa3kVsbfrpFiVEPDIyoSsnqbcLV/Msm/CT3XYwKc8rv7PK5f5Az7nV
OlYbst7USsc/CbAyyBocJJoc2zem4cfvlgz8xWL0YCYmM+XiZ4lsj4JgNTBMbHDz
uIYih9iHehtpbOQ/3PEHMMQMpIh3MQrua6I6ldBg48Ra2SoNB/KZ85crmTOuh1+7
hARpb7EMK77+WIcU83oGKnnVKY8fHSiCtnthYayJVqdzciXqWq4XJQMk7rTiW0mA
9TTcSM5jUpx/26s26Y7jHwcex8/F5qopANgWcX8St22efbrO5AOszq+W1snZmiiZ
hOsfmLFdwveqT8U2JEtnBa0gd1s7FN3IX2DCUEExb2O7gmDMjNFch6d4oobDg0K9
9OjdBxGX8JpidKg/HPVYtu+utUmHkRmzopNj9p4TYyvvbMz5u3o/n6UO+JBl7uyZ
keJV4h+2NB3esy2mVRVqHUBtrbTH3mll8uhpNq5lW3h/vb0sZIMaPfcE/DBzgfZe
WcgmLCfMp76iuDeuDw7Nhl9LK/g8LosPi1AYqb/Fop7ANC+YTrlzbBjWjLkzMn16
0WF2XzFjRQ5lKxVEUMsjnX6NQrwW6SvzbeYr5rgkoL5NnKORuIA5khyH6sWzIkMF
EZPlgBo7ma3En9T3zt2wpzGWbooi25JiwbdU5HCdzxgrmfym1IzMRMwCfbD1Shqz
fKjjeHmT5OBcQDjeiUdgFgJd0qBgovlGHRykFNBFP91BUdWr2fFJfY+FUY4eAaqp
AGlzdypxk++DTAtQXl/AhBIchD7bMtieg9A2Q7J99fvQ6ogZWQnesWelZYIiboBb
i84pFa8Hb6iatii8wTX3pb0Xj5ZbDjdB1vz76XF1XTWLosRKBs0prmjwJHt4Uj74
JLIEzyxdJJB3s9C3l+X47Rm6FybMPVkKBQrqswa3fg0jtizBCtZ89RyDsI2XzCcL
riFaFY162wueiZz6gernDaDhJz9p9FywTuWuhU6hbATSlEr5YXZiSB+l02XRbn+H
cp0HZyppu90yOtzBxvbSYUTEsVWBQpZ/G9sCAcOK4mpth0GWmajQ4yvc0sUp0VYu
JCQN21sz6ObO2oxFzLH8pHiBGijTcP85k2IXMd9haVSELci/Uc2SLwvuoAqhvGbj
ZrcTuQacsUUVqWQ9yrTPqGaay+e5d89kt7nIFni8fXXR7aTba39EbcIlB+O7TPAZ
y5foqkCw8a9c6L3hLfNlRdUyNQpTjNKw7vSSOyFC9wBuxaMUoAdi2a6ahOTDU8kS
2irxfUm1NPILOsXjG7+/i7KdOFYTTaxzj5RAOle094D0mkxVNSkwb9+4hkcPDd5F
5OA8kTTo4cS3/NRq3GFIW8OH0aDdui5Xk2nEqSBz9Iw=
`pragma protect end_protected
