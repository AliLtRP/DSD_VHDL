// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:23 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
cTTOuhhbp47SK+rAuWBrX3Yo6KCqVRLv/sKhrDcpA0qW/VEckJiCs8hjmmQpg6F/
2872YDWx8c0oAaVv1FLYoeeypEboRuyPdUkCa9dnEERjcRagOvhpWk1Sy6lOd0Me
VCjF9fSC4kUS0KPDuQxpviRh1peQqfoF6OtRCosKsZg=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 7376)
qg8glwRPvfQlkHJYSbAnci2HunPFH/YqkjrFnluCGRZp+9PU+1oL+uvFVVy56odr
4IEG1wreLklNq1GyPQdBCDEPoz/1mIWaJZNuA8TC0uZXbFDvvnZfiogPOyL7cHxB
4xRtwH4qdCUx29449RnBIezkPZPSN57+G/ZYEd1rj70EoHDvpGNRxe2MxgWGscA0
+GAu2pTiz0Lwu3IMh1tvyR2TJt0GQ2hpMsrgZP4/g5x+6q8dVzbCIF/gHHhsvbhE
P03/X36o2GkRruIRxvK844/QxxwHFK+VMfRvD7at3wbjdLnAWIISIvtljMQjs3iA
NzumjOepEP71+amUyuQtdzVksAVXRgwxQILqUL6s6GqMaQ3FjFn+Gli5lJoYTpQ2
A3vdrirU1ZiLu9BHr6XFjhIWi9XngphuslX8rkO9U85RwPWo4P48d9ahBZ3XiGM0
phOW8N7NSAAd5CRqLpMpJBSocGIaGgMdQPb8HMhQRvXMcCWEwnni6WpXO6JzqrnB
kKM8LWhtwnnuPJEo+oLN1JGSYm+gb9Bpk1YJl7x/HIiTA4wwEXDPfmpZmswOYRGB
PpTBJvwuPlJmYC7L4pBIrwwPZv8nyC38Yx+hIs46zWnbropIGWjKLrPArYba3Lgz
jUWuOowjFuEb22+ZScJhtp5MqSNEO8Y1YdAYTDjEMr7CBJZ3iqpiqOYj2BYNFf4M
Zl8MoBg+J0u8NrZQLD/FtK7c9RmUriE79L4W7hy4KCL+6gsDtge0V+GzFF5dDVT1
y5uBOuTHKj/5FUsJiOwIAA4vY8k7mpdeF+kMheXWcBs1Jg9KUMwWVk3LXv4PwL0U
D7vOPrIf4tyVy/uDvl85zt9Bi5lQQgua7CR3LE1Mcz0SNKyponIrtZLtmhTliJsz
+ajh4lVZV8M+tRb7n1tUgtlsjyGy7Id1pZ3eif9RPEK7ldQM2t56gfCDhE2yCHhC
r1MZzdf3nHumONkyGyvbjhu/z1aQYa9r9aQER5rAjESlCqp9MMkN6W3Fpq0ZFGqW
hndOOQmZb7TiDf65OlC8BAuSu8jOoUSHTsaUT8UISc3St6/ZpFx4i2thEZStEeUG
r3Ma5qf7MJSAa4x89AecDNaBOV3wJTbJoxRscsUTrdJvNYvHPd38zSlXcscZ/OWb
cOm+qOrrcKl9ILanKBgS84rwG3QbvR94+mGKNKhKqzdj/j2ng41AK5BAk/g+Lovt
eWE/K//GeYsz4BlQNbZzN4/Zyzq0u0h0f6BHBIube5ey0yI82dUiDP0VZ3lwCcCb
mIAnAV8ZoSThIkM0tB+FPdhWD2vYZNBxczMLRiwf4PcpYxsP4j0wW3oTa7Nsv53X
vP7Sd/fCHS0XeUHLvTnIIZyGg5I5g+BoMUAXsgk5wlEYiz+JUUAu9++UbDcWqXoW
3uLbAkodVFmGTGiiL5Y2XsKjcIwnvVkH398Xm575iPepzVqwF0DAaLGjtx3VvZP0
FPTBQO8uyVQYgdYvOUdAG68avmw+uw+e9QhWTBO7Hl+796crmVrLYVqOwVI2Z5A+
D210brn15wBTNFkfDF+yc3BhcRzW1Ixi7SlPPQh/WGKfNBXCOQi9bW/O8XyFbLbk
a9BS4EZ+3UzNlXfkREnjdoMMxA0eDHic4vDtoXc4f/r3Y4Y711cqU9U+qgkDgHc4
BrfIiyuoDqwUm3mhmyJUCQvIx7F64XZ8ds4qPqfqQjvwgWN/k1FKPV+fUHLtjqpv
GbVVhXtqqqHUmaFlycpvk2LWrrZGnQezzOUauYhouNam239sq1rF8dQpMMnBqu5B
u0CdeERYJTNPHDXQUBWrWYNOewxY2SPtuP+VIyFL1oYcGv7lHeZGNsiVF+1QCbiG
KOjWIWUJBzO82wMxRK8nv9KzTRYe9TR575+ym/b1lmfztG4Sm90sKAGnxzXYVRn1
FSFjKSQIbPeKrRJO9QpLP26rHhY13zq11HcC4P8tD8VZVCKSISvrEeG4fDwC3/ZJ
LZIQyTxI/3PP21CtJG0ZoZfasV0C8vq4xNuZVDUWoRgR5e0SmJq7FwOsvg3PuLVW
1OyyBRWPa01841FBgzhFlXAhUWp3jtF3slffVo4h4VQp01C1quBKHqC/ULYTE02J
CfArL54ahP8e8HpeTLqkskAO/bbpPj69JSbU8M2FoBl0jRXtMqrsodbxsekZdr6X
PJhPH1JDVLSQv4u/H/h4tbBTdZp7RJjOHWz8NPckxDxH7iaMk/iercalC6MJhUlY
6P9zhIAJe21d/5oWTSOsdQOOyolTDw9Zv/UvpPBonZVqX5uUMGdNMgonFLRXc3Qm
cjO3Wund8ZCQfhEbAYIQQlgFMwsz5kjpsDD/w/djdPzII21ZiMhpWLVD//GKuBNY
Sbo57aSP179CWGbVIHC27QyteZOSE/4cEzAhj1BK429ACr4g6xcrqXo3VvrSJoTo
qviajCk8I+H34yRg5kLpFOXPK5eaGf9Q2iZef9Lby3V4oviXxfPMmHU1GecPShZ3
Sp9d/CjNrnq4H+E75VbhGKNVWz2U7dQAwiNtoZfs/yoef065vyh/cVx3lTxfxuMw
yxNtawziXKq4/X0TDsOvlvKIDJ0EW42ux/gVqINJ0ZYB7TazSqALhnLknUOPslYU
AdnbzoTw7k8wgKpLd7UIOD9QEbK4liryvlN2AH8l/ppoB4sqSn+klrCfmgO24yqK
A5riyDaxVqtR4ydANAjeGbGSq0Uqj4ihsNrxqzDRAdPiMK+F3YgkW6gASdGhJUv2
IFEs1egFUj8nzMq5xgjvrZ7CfHbYp/iS+yXE847fNn+VppaMyTY9Ov9+DYtAtuCI
RVKGuAZXZ7115JzYqhv+LELodIX45YH95/ODh+gJVJ6zCZm6eVdJ+Cq2PgQ/hGFO
Ry3MOyBWfGzMqY/k6liXSm6Se4Ci52a+BF2YfduUbWXu6KS/oEmNhFWs/1T/mPVf
5sdf7JONp5xQj8w/4ptWAYjap3y0pnzHgMmZFwX/mZ7gBsh6dQJ+7gXCeFufmLYi
p6D8j6nTgHu3h4R8mC2OLCtXyC7SvWfIYHSTk8Pu5+5CeKF9qK4qfHE1c2pCMc+w
sWTKOneScZS8+0Cv54Cy2A81WqWTW97FMXpPqu7pBfnc+9BY4jlcfDIGcPycClVS
WnqVtN6CJIYtT6kG7htN0v6wVU9n5YDqGWn4zoFxNTxGs2g6eoyeMgodf7EQFiWl
O11DaBV0e7a6RqVd7TJJ2sU3mQEn/8jvbJqat7EVdtXfw/FqYEVOnfNpWPr8Jcv2
VgxnrWMGWlk8Mr4XXwSvnB1CqTw3UpuKHTvSwnFHhmk2Yhu2YK0W8UNl9kv8IYNw
rH9KNNosmLE1gevgIvTi71yJtSbKgcKpv7oa6ETEYUjt7Gek+9dt0CcWJQ5FfFYQ
kKDSKP1XPMQlXIFnFAHo+CKCadNs66/mfVIuGOwcPdrAeveSC5v2+bLruwlJM+Cw
v2DnzbHZ0SIyI+XrfVjJ2K4s/Sds8Y9jnMa+HJU/69WO4NCy8mttH5T7PdF/Byod
goTeh1S3pVywkQlkDjcVyi3b2+CNY5lGds0Xr6C3ffFA+lHUDgLodj0n6LbB79aA
ND98VgngQQww17Swt7FMXrkUezdx0dP9lUFv0Snq4G6nqTX4bkKOATsjRRkupOBV
G4JE5kX1LxAF8gei1oXWpiGXfEKeph1FP6f1pDlkm7bBotVB6m5jjuLWPOQEVmsM
5HE0GF4P7qlGDlkCSX5Dkc4sc6OVGgnLFp+mW6tLid8l9/UzCNwww9CLZZ29LUCJ
vVtnPkdl8XDxyPNxyyjZB1uGahLtl8Yrg7LjoKL4OzsFpxtri4yAhuP5wTvFOYoi
f5wO+Cwx7dur/Bf09Y/XBcAKmFFusytiP420bO9OgCFUQqnUANbbWKfXc9CET+Y5
3pyFDsUcrdNQ2CXRjERoN6HR93SqevAwJX3kH0PZzuSWNuWO5b2Wq3K61ACVkvu8
16OVxdanfwxFZvjg2+9x6wNHwmRtMmv12+Ru7J3JZlrfXbi1Eq293+x94fUxKqaT
RxkKT7jYCfiBefHZ+OrQc9ipku6KcGdlHKMrfSiHRBJZzf9+0ocU4hLuZjlRlHjq
vJv6FjIx5x8/Jz5AV49ojW5Y2o7SOZh6oyZwLmwmftXvZDK+kxXAq1eB4dmb2pc0
Y7v3qkIaF/hjXB1bvNIKm7DYd0lve4NM3vJ8NvtKWkG+u6fft3TQyu6zdpSPkoFf
ZKZ7QrPp4R7vGNXxLdQpRGKsx4fwFjWE5DMe6zMq8GDkpommAzuGaSA7D9SnyJsd
/bVY5nuqP5upk3fLGksdR8j+MACU+Z+A0s2xe7GThBZq/YiwmNoo3mkHGweKhdDq
69Sp9MFp39T4V9ZJtAn+Jk0vVhsLXCzfUTfpqyUW9Y6CTgkZWo4HYnQd+Gl5/6PI
5Kd9NAsQ+0dvPJDScEzRyGFJYjWJbaokYcthezGKhbL1nqP9cu0PTFhGXZbiXUVh
aABZqe7wKUMe8wHPvvNLyr5piD8lI2CwjGuGPJowZD/9D92Do90pcect4VvXtkux
2uikZK7Nzygyu3eqk01onijmhDxyjkoVibwfc9WI69HUunICxz3s4z0G/raxiHqI
YkQ7YLGJh58VlM24lM3wo3NdV5XsBqr1ch51hecmhupE+yw4KW4ztXVqivg4b9EY
EJACIcUDstEOYNOR9jSTnDs4M0AJqAEiFwrG8g8Fs6mPM+0eM941vAbWzZ9RDRk0
BGm7xPieEqJFnYRKRNWzbgS00+SEJfiediJw8DeaB3cE50idiYuXord/C8/q68Fx
jHRtceLUYTur3Wi+vx+79UCDb9u1YbKv3ZcbhIW5gLf/GcKzM91LR3ASkmSbKrn8
K9YoCJuVVa9EsikpcIKiGla48lwuZD2j/e0Bcb0eHguLj643YxPyUeJdyUMA0F5Q
q9amA0XdK8hRbda/nIvJfWuXIw+0/Sas2s2q7wShUb/Xs5Zor11E0Kgws5VCGrqf
tTsAy3aft/+ikk84ZrjTIosurJA7Wq/8GF/Euc+laQgZ8kF/wujGrDIClyIcSU0b
HUSJFKGHGJJBqzjYe88h3+LczkYvkGZemZikvot4jKWJ1kpPoiKpc0Y+4FKfcrTn
CKHVm7UhLCj/z7NuVjnRobvYqjGlDdQBFcQZpRVTvzaWsaridKMwghxOsSL7KWKP
iUmXZsvfUaI+FWGWJA94U80LZ7zWCmDa8OcHk/j9RGgDq4DUoKP5NCBxe9R1oLAB
mdqVUOkqEgRBE1ASycu63q0BYGY9raBsXnd87CWIG/nRFqnczaSAXAH3f3l9/Q7E
Z7waMxaJ00eev9FqI0tgDUhnsbesF8vF1+Rdj2PLbkes8HnMLnB+qKAF1cQjRuDs
7jiuoECagd1uCczlrY5HB5LD3KOiUULk4UiqE7UFpQwK9+1V+TywFt+0Scw72OVa
S2lBdOBU1MfXdA4IAKM2Hnqsn3LhLszn9KdPqvzq3j8URPUYDFP+etPFqxwiW5XE
5xo2xzMlGU7LlrT1iCQAWWaWqgU/0Wzn2mSEeTyPFUrhQnJzIUNSJIb8AHgibpQk
ZpzFlbZmVwPYGxkmM7aumLf4NLdMd60giZajwMuhLpPD9xG1spR4DRFCPJPSPA4D
F7Bt/g7qeSkLYN7BqkQ64HLEQv5EHklHwBZ3bPaKzfCH60ihuC5Vqn+bpzdAuOos
cLZWgl9n1l8P8N7ZXGcmq2TLqQM4f3NtnlYUBU0a4GIfn8++mtkrkhhbGVtqVa0H
l5Q5Z0tudFF0lcMfOgX7WLmUEkWpT6K86n6Qvfh6ZE0g+r6jc4mpLA8LoxPgjYFH
owfQNDQ27YQUM9Xdaj5TD9EW/jpQI7XbwNfbB437b3JgUDSJGY5IdnUElDKMcygu
vXMF2kYu7RxQu8nPGUeulpg5Uz4UV+6+XQCFUWUADgXY83krZ2b+A+xhjb9hJwq5
tUPWyw6UqMRY7+gh55QliLhaqGFbMR1OH+cc4D3+z/H6hz+37n86txD1jdFUh3C7
1ivXLqpZhS2Cls/V/R6sD4sYMoY4xPMPtCJFq7vXEcSQwO/pEiya9hUqs12uPGhj
UB61KQOaDEhlbA9QJxmW5XhDYeD9cfU0+5mmPShacBA3CFJAgHdVDE4mEeKLNjtM
yLLcpL6IAE/b9sSlTU+CWFIR7JSuHAwNMEVBi/gKU8W8l7e8ORy4vmBLnhYQCx8w
MMz0VIHNcECOjkEh5yBOX++FdJbDam0pxiHJ+F//ycKx779iDrtNoe6T3NIFHETy
YDHvVRja5eNrFzeS5J5mwobqbZSbzbpVqdfS+MSzBJyI7MI3Zy2kMtvjtEUQdvAr
5kxC/yDJIqthCDe8XyyEibDl+LVj/Yoc1IQ+Q4PuQC5RwP/BVFrYMPF50k5kOaos
wqHjzFbzYX47Akae2GmQFElqck7GkdCeSeY6yaBuTtAuF9cAe9/zuujjVj49of8L
r82Fdd6lq8cFykHsselV4peW7hTkgeUX5lkHoV59ACY585t1ihsonJPLhPxoycDQ
NU+7zKlzLI0wLtSlj/OvY61yNDEk2qI74qVbZ/3gA40RiNQEQQYnNYu02wdkaIhW
79NoK3udrhqzKPEZWX76fL+xY9aslobFodNWJfY+TjB8ZCiRgjCQGsAcULyJKR8E
Q9KDAhGAVDu9693kKCdx7GM/31UKvCmqB+2owr36K0xYccldX2oV+9T60n8zCZHq
t94EIz4K+j4K6dBN7Rkiw/wTDa4MSwAdg+a1DbhIGfiPIIodClwwSR8HIDZgzeoH
S/QzCqio48iz1JcfTylDy2WI2Hn0yAh6PFXP35o/YdNnOHmynnYp66u3z5Zq9nus
XP/lFcsADzzjNp6TGqqTjsOaMT4f7LcHlc8iB5dS0WZGnGrazf4koJEJGAG7G5Le
dQqMUznDNz8xztRZALriwoTpjN2fcdRmvrKwNsRSgkv2EL9yuUEVZBzNg6pJRdJH
6Ejlf19Z6uuIRMSDQ9eLhivVm8RpGH0oIIXP3gN4vq96Y3tcw3XxjDUGBTasp8+Y
i5tPUgumfoI0dJ/mh9UHhQNiUeng7wjY+HR3c2t0caI6K7hZzxoNW9NjWwjHjx9d
Lgp/Ol6Vd7BNi/7/wm3DSiD5bfbjSqlTh/HWAwNj2Q8XJPvveFUh1Ngq4sSpNI9G
p5YcwETKiCUjXuIoBnYmcnOcXy9ByvVlQ58NqRiEK6++px9OBwQLRw7VcSbTB7+O
pK+hZigcvucQWByDVMdx3Wi3SQYYx2y1PNabthmXgdzbgYkZb+EV4R+jh+b/MPHH
fyxFLqb5eQ943IW7cQNlOvPJFfyFaB1Kl767hsHAXxd1qZq9McOA8mEXiQrGEmFi
jofZJXIgvn1GZs2bZOV4qMefmPa0Fq95A3Yk46T4FXCuhBaotDrRcaTURjO7lN1m
P6eCdFJI3DO4j38hjffiW+MN0sD3BqyTls8hSdlW6ZsYHZCy9FpEq+EoCkASFFx4
d6w4yqh7ATSa1bBlBis4I+XNX9he7YVt/Tr+YfXxFeD+rGikwYnl14tUblcaH9bE
DTffolLFXqQ6Y08Of0USuCQ9iA/MEPo34ukARiZpWMgXLVKMcRVsTT9W1szhZJ6r
8I+YpwboP74qCyt95VTx1lcw4nyck+b/rd3MHgAJ6uYwJb9ex46N1KgKKzB6FLs3
HFU562wUBoxkXPSDr8NzVleWYPjFHsRmjHDoG3GJvXW3DuGIrysDpupRu2o9Veau
19N16toam9wOrf2a4MNmoFYeOYC+hfNG3uqmvLbXZuFPZ0hQfn0oCrbWq5RCXrit
lE+y/YOMIJ/FVEuk4gFzdjVYw1HgfFM5xYX0DsUWgc4ASfiHvbIYuwrACbfxgKmx
y/2Cl5qlBa1OPaqBcWyzS1Z5Ks5/T+5wNNNSxRnt2zF9mc2nFZffHtKOjEw0Dny/
oaypzL2Gxam2RQBjBpq29sJf9Vn3aDa4BnKZ+vLAqL7SWeSJQIwsaRkP90DTNVm4
Hw1G838w2aE6vd4jQVQeOHa2YdiblzNXBzrJDkOzYEl7V8fuwqKpkxdkbCLtdGxc
aVNg0HXRGD2suKaSfx9PfHAZvBXp7HO1HIjLZXOV1qDM4OYA4tTZ0LOYflQ+CfBX
YibcHLBgUb2MDHTnjPGHLQdtBw4wPSbLm09Z5LqY0xwiWbuoP38eDVjkSgQrJ9HX
BfB+jWCZQbEtfRdHAxXGapNYPGxIovrIjaAfY4SNgy4cg1KXxN92cAVp9cx8Wg1I
sr4lX7gpNMvv8/nfwWSA7A/kVSsnWuhxMN38HWnwVXrqnSg05QUFI6CSMuzTwpWL
uKBtXQTeqTnJlWYCMBg/WO4VN6fPPanwEb39/FTrcKDs2Ih+/XzDOCcCiFbFR7g1
O2iKB/e59Hi6QRBbRZYj0YLUAmCadzqsRj5YBSNJWEwbEnXQPVEAiZysV6qtvxC5
c05iWwp7lq773rmArAW+hJPq3crS/5Esl9FulouCG37zmXTV8YnKAfWlDRXpO1eG
cPPuD77OCLT3jFDLj+uO5IMNtCj6FxT62Unx+rsr/pzCYrJlhetA1HIAchVsZdtG
bNAGmm8sdudBvSLO9+gCPcccU8aTduituHKi+/8zS3bA5fOfkD+kpg4+9SeWCzwu
R0Y6120vQgvHzOSnztUUBsZiHs7GGuBzCUfdWrbHSw96jMA0j7zmVxzRr3lmUYUi
Z/CJrQfZscJ5De8O2HNOeWqA8EpyIW+740BUPnU+PS9D3uWh/N7bx3McjSWoW0z+
Ipvd0zF+ylFOksAIKtTO5DSyVhei/noGNL9yxgW/rpf2E9vekPIShNcDECz6f9Rv
FjVWXowNx32bfiFL/YGuezDtqQ0QY+KlUIC8VoDjhD4kYsREni1D/llGUj8TszMo
6ltXpCbpR6dB+oTqufhu0j8H+AzRpzbxiJRUtDbP2yaJDHC5Rtn8hTelcxlQBweS
ezleYP7SQiyAY7D857SXvwSIfvE5xqwgbqAmlLEysdwuRb9c5JZEl9nQHYYadsI4
iZNybp7c3RaipDzCklmeVHjH9LtVhH7FUuJvpkMTwk5QGhFgoPnVWcU2g9HBJGgL
Vd6LX7djs6tntH2nb+uGzyrR8F81ufFeKqt6e6wdcrPx7JJFcF4O/q8VrSlayEfk
0GBZweF5oe49K6wmI6yzrLZ0bcJ9n6Cil+tE0RMV8GUFEAqWfPOmpXrmR5jehDkN
W9uAofwUVHdjufHfKLDUpEGp4L6+pqS/+k+WkqP94O/aHzH+KhFUhH9jru6/mqKR
OVjZG6SJLxXaBTZ2EmrBLsw2x9MPij4bquzbtghaRDGXaQiSt/b+7lvPdFbs7NOd
mN38zDBIxvwwu2WSBzRVuqY1H+TxvQbN4Es88EtyyfP9baCXas82uY5of7D3sl1m
3g0oROiYDw9TyP5mPT08mpL7VfrvtS3MumdeAZ2WQlclxHTT5F8XYd0skFG4RQuf
ENK+guVsQAA1xw0Ny4nyHP0l2blCt79ID+OPIak0PTc9Rl1cCiruNBY1XLk1a9Ho
CYBTK5vEJCurtEAq/E1Ed+VQgZj0jUEBb6dmRqKqa+/zX9Q/IULVyG2dhdDhgZXi
MCZwuoj9p1x9t0kygZ6de6NiVS+C9FP5smXp7zJVfrLb8II7XgXneFC4tcdEy4OP
q4zH/1ykxeAlrp16QPd91WgFey1lWi4Jbvgqne9G4+g70Ygg7j6lI5KGKysbsLgh
dvrKLNqLqTcON2k8gCsCTqA6zsWsuDLer5zDqU8X2Ydd//iNiik84cxHMggJRVer
c9+XIDVRGFvQY70mFuvVXB3htVmBzP7FlmtR7mEymz4=
`pragma protect end_protected
