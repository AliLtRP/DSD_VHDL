// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:33:34 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
YGc5zSWfTwUj5UTAg3z71y89AxJiVwBg2pKxONLJ7TVyCcR/ZnfC9zSPoLyndk9m
bomdRsVDB5tJL+/ltyDbdMWNXxZA08GJ1+d5lYriXXabN5GPuSYaKrmkc5568odx
hQ3MeJGglG8dMxJ2ph7hDO70zNhC4P1geS7z3iXJf7g=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 9696)
SY56wJ0p67pY26jqEbDKflYszx9rfJegXldaQ3Tf1qjs9eZRsRKQ4Pm/ycZIsaAp
7CXDCWOIzRVaGEh9s9amWk7AWOBfncTWNq1Wudh4BFsjY/M0hACOQPE9YatoSlfY
PsRpF23+WlhSoiRz5WuGW3lkTAxc6YhFEXuSbwG/UFyE147WpNCbVFhuDXzVfOeR
l8kTaGSnafJcxuFjkSlFlDzhfwn+VDsABU6SwlWkmlZsHPXxNCvnsEXjdU+D4Qw3
4UcapYKxzSDIUs8k6r54JJqZj84rzT00YNIB/pofC9KhqI6QRlMSlMeEP3ItOgmg
Pbaf+lEP6W6Aynu2Kgun33bkZjLa+mZSA+EfupDALi/D90oMd3rU7pmM3X+fZHuX
6X5UHqI6h8d5oHyLCgcqeDVyRYl8lovCZGDqzdcOAoyKsgjUfiOO+ToEz8DpeCw0
dUuF5eJat2bbRrkff7MLgSFPI3ewkw/yUV52LIExH4gX5KAl3E9qImTXvOsNJkDR
sXN3af5THZ1gFLQSbTL+Wj9o19fkBSSMx5YBnvVgcC8pV4Vnc5n8Y6QOmpGXaicW
vSXJ+oIagIugV0jEabU8Bq+2pfi+gFfyqA2r80QQOs0mrtAXfTiNSnzuCB08sqPT
50FkmmxJ80qTzKNV/T83AUua3VKqsWjqfZjq44MhcvfXaE6o805F6FsZxBXwTlkF
iM7/DrePt9UQ5xY+d97Cfgofv66rYy4gLg7qJ9eLdm1tl+sGN8tFQcheYDnOQMwM
TnORoGCENRYJ43PnEB/9ve1hJ+hF1EPKEiiO0sYOZ6z8wsHMsswWQToS65ggRQNG
DohasenPW7581UiOMrzcXlhUbcocvzb/KGwBdSeloCmIiqEzidp3EUs/dXs87UAZ
rrS2qB1Mi9mlpWbWaSWDsK/AitIBHODqrOYrBkTkYCb4yZg0jK0AYlQ9fhDp4/Vx
HwMpf5BuvBuBna59pyes5WWUWmBRNqD+zoFvVnxgM11GkfYzMaVpBf6xuu4GbUPH
Ws4trdz6D+M7c2f9hhwHvWWcpNmm5BWx49K9QEXnTDnTr+Q5rUT5Cu8DFiEsCRaH
8l/aBnR7J9oJcfGR4TBZpnC10D+ry9AnbQbA/h2+9d2p0izAbIVBCmMh6c67Ud47
ZmXQVJ6DfIYP4NVKECiJM52xrJmN0c+7XNURUrJKfBICET0TsTrDAcp1sMnXCQSI
iZA45crYJOgmjqDRn+D2UNgrcpn5WAdKFVSTsRzlV+ph+KRROSdQW5IauGyaERkb
nsoUxNteRWJNl6kS/8LNBZ1lS+ShivSs16lxuOC70N3uiNY0I6/Ge+EV32CPkiF8
0M6DEs6wQ8Sc5Aqh9RfCrfkBeRajGPJG+H7NIJPDzRIbk95dVShuizwt4ZXEoLem
Tg6Chv3Tjc2kpdnzm9hrVJafZ6qCWVDZuDEaEeseLTGbABFGGWtpT6rrXJoSYMgD
sg4Vp2IaICywkAXQk9++y2QZ/10z9zFWGr2dIAyJDIpIEJhAx6vvx/EfpXCehyu8
yo585x0bs2jNmGH6om+XBqbZi5bTNr6v/3STW1oKRLA6cHstSKyBZADkcc6jj3Yb
qo5yx7xuIf2ojKl3Gly2BjJUFh9u0kZAssaEwzBF/xH1t+MzuZXxFtWej5R2BK7u
pI95Isbvg5ElJSkg+Dx5tugeEcEYQa1HEc2OH2YkoMFIYKBgFE23nh3k3G4XnL0Q
KGo7c6DflxTYdxy3Z3wWJBLylhWpJV1PB5JRMVaQ6eCdG63hi213qzSLweeVpcGz
e5k2aQKQoOfgEVXGOq1LULNz4MDdgp9jZltywKhD9PCU2q3dMhtcr6SwQ0ihmAy7
H+BRtj6zy/grk1Ydke45pFOK40zCeb0sSh6fKjSSBsSe2J1Vjl81tUh/AX0BXsFZ
1uaPDoZQQDOZJ4S18WHq0PKjPUcJOlvaup34dCEU7UiFNUU3JABE8pbBPtxX3OLL
0KX0Dn861GwRZKP01rr5isGB+BmZd64mEWWmzMntMJzi/i/9Cbb9EwPIEX4OG1+o
e3UL+Cie/f0vKK1zwIDC1iDee3DT/EfB3iBNLyqgK/Vu4i95XRO3AItDt2iE08F9
suaidHAhJyhVspWz87Q341Fy8h584Cr7Q6KegkFWUiobIrkoMH8gFFnCWFagoKzc
wdwGIG7udMpk1PdBhe82lWZjiTg5un6TGnIeNijh0C6H7d/lbjYuA+z/V0Nbjadp
Eveo4LmSqJM0jHpdjGBSHL4H4jwu95f9k7cCnq4kjmB4QsUgl2jQPF8IY/yOS7xl
VDMo9hFkwDgQf34e7A0zMAxnR+94KWL86hCVzHJ1dCXVfgoOvjzuKK4AIIqn8kSu
h5QFA3QnKbycaWH1l0AGhXST6hpDixeldfSC8aMiqdJGHVfhMPMme2kwll7Y0QVw
2+1uGyuuRSN8fxFpOzCJwkKEZbPylxxX6URmDD4c/lncDkwRuSQlnXxGjtioKtYc
n2KDL1ZB3qKXL1Ssyjil2Hl7nWGsEPSDLHktrcmdek25JewfOvY8EXkDkBviAGAK
wSJVlqPGIBgFWCrYcfxxHHaxLhJZONeSFXl+tVl1US4bnkFckxsYBiNVPjWBQGKv
sPLu9rvOlctBJjd9zlPBvGB+lQWl9fyYQEpKW5fWCNuUkcenYdBTnonYljYKItOI
TVV7V6dAGEgN0xVKVzH39LtqlaOonxD0mBY9wcRh36JqV6jMEukzYqtwofgPqKgb
fQ7EkHWuTkGR//T6bbd7UXslC9maIlp9wzzthTVpvAsB6gMPXvbGFxqInHriRb/E
4ynpzqIE5FrPmrGJz6pfRzaoafYdDD9bG46esyoQTbZDhsWrLOSVDDoKOQt4eVC3
OL4gSW/enlh8QiYbAdOI9EaWDGM3ANGmsANP+ILtt/iZL37VhHc1d7vXX4eKchUh
YezDQp/NP/I9Px0bi0XWi6niIPvuQ8SsatzN46hILVxXZxXqnnQ9EcDgT9+SpX0X
Amv2AY8fVn+8DZWMtjoygJrTOihZQxmp/KoyJVe9+21BdeLMY4Dj84SYMJ2E+/+V
zGPe7geehFPfT+XrQA3Jq8DMGRiueSsr6VVxEoqDbncy6cv4DrSu+PLmMHK6nRtQ
DULnKw8hlCP9L7mxM1A1a5kbYUkzc5LnJWqoBXF+iNNkVxapi7hUDZHhH1TrBLay
F0Iw4DmCgMdmUPIdisogECqodYn57/W3jzjqmgJFPBw+fcJzsfcBJx8cyC7Tp6Eh
+M6y2dgo/PtLLrwd6ayh0uIlMzIMJIZgSNbo/Qmpjhh2WFKq+WZI4QYsKDgJT3Ce
g9iBNm7iCqzUSHLXEqI68WumnmQospB+9U8c8a0JZLBd7sacnXYajyxz/FCa/o+h
LYvw86NjzBGNfi2IvMUqn2siqe8vnoN27ShbscxfwF4YdKm+Il63La+OphUduUK+
5qAhtau16dY+W1stO1eZQuxv8OBaDs3m4+WQkKiWo1GP8RtA2Av9+uCx0+f0tjvq
9ERNzve6MhrRjqksMN75c8afPE3bHoV0foC6XLowC0LIrH5KwrfgRotkaRuSc8Dj
k9toCkuWw/6iyg95XziqxAhwfqY2Q6XtWUPAkPjhHeq9zQKZlzHgVLtS0QHD+lFG
Mk2F38bzw1Rml1/Kk5q9kRV0auZ595mW9YDWXz5sxzIQGNtef/usXmmjaMJD5vJL
GbEw6jyH9bOc2WbbV62JtnqgwIkyNXRrYCAIIuwPm/H+SBCB8WLiY0ByYZ2VsjxP
fgyD5lVWtEO6tL+r/FXx1AdDD5b5DmUI/1+IBerm87X2BG/Srg9/5l8PwdfHAxIo
8F50/Q75gcw7Mu+6DoNbiJOcsYVw18CA+pe4vqiu+XXgyEOKjNWG1bB/e6laIIoh
IVTLSP5WweBm8HixmXfb2brNjSsbmuzn1go9hPk8wr23Tsff0PD42x/w5N0sqQHM
U/NS/fwbuAwKFJLj51bwFZneZK99jRXAsH9Y1kcQVDe9qk2Gy2+KHpN7ToQKyjL8
jWAW2JWMQ034P/OoldtSQoOjEnexgI3G33wvLt77fTswOPddHkjfvN/QAjBDPtGg
7b1jbP2ZqQX/KbU5BjLnNcZev9904M3ONW9hM1V9Uc5Gsz9jDkynorkFbZRLmQa8
ScHZ68Ds4FJThZ+MH9P8nLmqMFl8OyJWh7TM8iLo6xzrqyaEuXe8scLd/sBQKvwA
spFQ6maM+1BbU5yT3zjVNMrgJqKgV/M5SIgdEdrHf5vK2QFt1jl6l4nzMGn9Cddd
UmtRM4frOc76zm33duH9by/AdSRhd62Onbg7NoSKUHUc7uXt4nzivsX4iddfSKiu
ZGT7M2kIjIvViIKg5g6CXHhLdR2peg/Jqj3V0dyBRCuzysm3AmMr7piDvyExEyHv
7XdCfFv5iPXxQyCdY9tY6XbQfSTTFqFNyWgatKw0IX34NaOEHWYep42lIvwPCVX9
R7snfrtMNIOYFXwMJzrOqlkfVxB8xuwoNGh1hZ39N/brGYkPJGdJiVQ23FARagh2
6vYFUeIHKxVO2Ed/cZJmO6HuEel3nR87qh7/LJOM6K1ofs78i3ZnWEPiYBx+/4C1
IdSjGEGuL0TJntp4v5tPII870asF2ciEXkW62k+5pQZ85aamP9kp9htNiAue+Dgr
XRXDv8icddkv6vR1VP7N76h9z6+0+68wFZmY7J7kZq32dUtGBuxLHKo5vlHjtLrv
aJ5fyjuVw+WbDe4bQLuS26/wkqQwYtiM2+sTdQ3jEyN0bQAezWQkjgnmkDCfRTsG
BhtxmdiB6oYVCEMCtMlLO+6oDxmaQe/Ut+JQaMUvVX+OPN8AJBMASjCfE8kC20Md
gWxjlb/rI2x8jAjV/l0na6nVNjmX8cnABZMBteflgSFabc2KXimvCOGynNjvgHue
JlvqBN6kxEB2YODSrq8KRioO9IsEGWin5sEW342Cooi9YRzWCPoNQDG6WS2wJVA4
FhEMA+5jRaCz448vTtItJXvPFPgkQB6PzbVYGKAL5CzgStT3McI2RodbYqdGhKLN
OVBnuG1aoMcxKDyeZ0MJQb/poI3KOPXdFxZQHb4PHknYxsK3jQmbAlde0zhGBiFv
/YXgh3/1CMpyXgmlnzg8A13o5RZORsTB2L+oFHYIxmc7M2xqn+i5ReCpqsShtT0i
gloRI6d1Cpmb4LvAWxh3ydImGAjivv/UKrxgg/HlhRJgJPBEub8H3Xl8Gq2JhjCx
ggGfFNVTbEW3ZMQ7zH2K+Xv7RUtWxuwxZ6ZuOKNpyASXqtQYnyCyDNq91xNrOiPC
5qgB7OVi8qWXzb6Q3mJM+tPvXGF+XC1xLFhAVoaW/DIQwfZEfZHjFKs5lLIF9Hv6
JVfPooTjYHtwRdgQWHVwnCwHfe7KDKVfFVcEgr9pILlMtDtS1vv5JJ8m20aq5S8w
sg/0xgXX1cTWisg9kr0GZxmo7pFZxWFS70bHGvOz25DzN+r7S9oLRVG1FoNoc3AF
hfF+CqTZ3mArcyIovM2GCjDW8bDXrjrwyRTrfgt2+ciQ4irMFsDG75TLycJF25s1
1e2VEuNY2JDXPh3taFe+SIjz20CMZV12LSbtT0loiW8rjldWqeCFRTmEH/S4yAEq
BGkbgbUbKyOYTArvfceCe+07fPnUNQ+NBQPC5S1/HJZOgs4IVYPb1DAi46tFoa4J
KaQbp/Ndam69WM02uqBYlRbiPqVB8po9zNwJWH85R5mhhGGIVUuE7aXSDEKCV1+F
ONwFlwbdnKCJbfHHJ4npxWkar2Y8KXZnnQXJoqWhN1teut3/hmgrwqH7LMlpcE7t
67NvbANDOG4Fv2hKV/6FL+1vxck8KxBRmR7MkgODqW9+UK1PsP1+MNVUaardM9/S
JT+WxKxtGigSctX0Xg5Kiy8af4kky4PZuewkTGRrTNb7nl1/fPWYgo3Z0KIdyUxU
roLEAiIXqSt7Mi39eSxFyzhu6xI9+gm2t5smIXv2GgfnKcsJmu/gdR79Dk9IHMPn
xHszLJhFR61wjkBvi5sE/+dx625v996w2m5oIuAjnZ9KjXMSK8KmnFQV9arImQKF
hVAreZ8JjBuGRJaYewexnlWMP3hohiOhVxIT36PsxNeR6bScFtbhPuW0Ta1YhRUu
9FedeKjtJk9c4qV//iLG1QsyUIx5sTbKkC2Gk8jZEMmEXRD4+Ueb7ggaSyBAC4mH
W7WCjS/0oPIslnX5IJucbhNK7fO3FvJEYtlkup6er2sHsjR8jP7iu/ZbQcMpUlAG
WWzUAVlp0invbrmsPmLR8y++zCKzPKQGGTXbvmPRVZaI4Ao4ckJDv2YKYbV4cYMP
AKqiTWDFAmL+mEzgdnQcINnpBr3HNDpJWrG/a9/2ZkLV3OKWVns/4LUrl8KPDpEr
DsJxWQ16R/DhbxBZ6zCbguWm+FxKBIBR6MDnoOXVXerx2QQhx6Rkx9Dtye0xglkO
i6Umj7WqtlCSPV1fMq64w4ij0xOmY4jAYvTbSxYdaHGTsUlbftd3LpbFRfdMX6LC
Rd0vT1xeKaCHn58xUsnOeCrVqzNfI0HhuqvKxVSv9W4YvpGSIFnDrSsBkhjlegu7
Cfl/Vz/IZaNYzPDvpl5xHCrso4DgME1qWA8/U3k+WKnjLW9lbMX0WMjhKtgGLwCR
2Akva5StNYEstjcO0vctPxadai2656ZbY8gJDrtY5fHLCTszMMnTZz2SNAO5Fk1I
hW6wf/EIAWDM4fS4LD9XWriqZlaWEHVtDKs83YMCspnGvpxpH9PWtSKAMnQKAhFE
dgBJGOatkdpLTTCq6/p+3XmzMvTKOL0cwaVbC3Mtc7wWdgH8P5IjoE+TP9BQwU31
6KvrnaJU45Gr68aHgs0Wh4dMRx9alfB3s0xuNPoMlFKRzJVbVaVQyFWFAbWftcpY
Am8Z2XfCmVMOxw7GXKDJPAH0BJdjhbpSnDr5n8ibgU3SdJA6xK3ZdrfAwrSCSHbS
j6WoDMSPUZ/xvyq4yUJT9j/rvd9ui3AcQ2tQBG5Cnvsl5Eu4PazAb8LzMiYjJtxq
E8yGufxZAlsM8z3KtgVKxJz0uvkZ2xQjjHSFubb5MTv2xMKvcnfluUJCyQc+Sl7W
2dfCviTIkFPjkVRbo86bzIsl8EKoDfetnMIZfUMjlqtK3RSP8KhEgTt47WS2MOz2
XETnGKWz+bTITX0ALKXesWJLSm1R09LTq9c1CdAuVoviDNC9CnbGpRu0D6U7OI/h
h1G6QZ5GYdOlCP0hiUQ05sAQwOwS8ImwK53ubKMzfazkdOlxtL9SJQT9ixXYTvKm
EWX5IDkZRoNWUhS5Q6qe+X5U9ZVy/XJvsnHsVteDQZuouj+od0NGwK8GGjr+U7Cs
Si+w78WK5I3CV7ozbnFqTe0WbORJE8XqpAW77hkjzrPEhEmmolBx0XvMMFIGNcH4
LNFeQ5h+X2Iqb7UhBYKwN6e5OlxrwLP3SAsopebFvj+E1TDz4SRA444MS793VOcJ
ZRWdOA9FgoQxcmpkqIypwwLbukgNi9pu7QEqFjqVQnQMBD16fGG+zQrkGc4ASKo9
DQG3yGT6p7iw5jUolJazfua4lTnPVOlFAbi2DHC6x7zk11+NOLH4cp9Q6SQ3M1Oa
uSydOpz01v+PwCxh+Huy8JLW/5of7G6EckHrgBcwY30GJ7XeLN0fB0dieCuoOKo2
Znyw3qgMalqTs+e4NLfwY6aCqOmQ6OWX76MkXHusyXHHVaojFIgjifR3IeGST4LI
bl4ewFzb1RPjhLnoXDC4LPwXMsxhpGU6QrTmYqtPddNYmLTl0V/GHSGXeHVhk4om
usLkzbDa0sey5tc1MQfpjPmHaLeB65jYsxOiAXRgmfVSsWvJknUv2X8UKdjlMMqT
ZGtVK81qdqfTFAnL8fLgK+Q8TpR8yGjA5Q8qiw9v8xJW+3zpDB7LMQjK18A/7/91
y6dCPKs0KGhe6a5A7ZFi47UfmB7kUGbVrkkpOgDyFV4T1MgViFXDh+/JlP1a9TBU
giKdy24ZbesvYVeFqunuynIwvBY5sz9N9N9M7mb8CgipisC71mtNDhDDJubt1RBL
1lbQp9yv5zJatKmjE/sdeZUhvxMgSN/ZVeUxPXptq7IORkn57oUYJaoIoRarLSUO
vLdm1JPgiNCRWGtB0MYc8Wfa0ApzelKnaJbDbvTniwn99+XxmCjsvHEvuZgDBzr7
Att0GFzhTeWopHe3Rj69vyf3gA/rnz+6eQy8liDvIh/A285ViUSXKryFJ4VifICZ
ijYldx5XaLSJ0EP4enE3H/JtgEeHqrO74z1dgwvRIsnZh3cBNULkLIEJRQJFAbm3
7C43w40bN6HIXJo1OfuYoQLJioKukDnCjhC5HaF2omHYEvpQLDvJX9rJdBlySgW7
fOBx7kDeqMWxIVBFFyjhNZQEBlSTPydztAXtW2wMlIuHN4CHlj8cjtpyYSIrxX14
WfInbPCC3t0gpbMFe8hfDxwlavIRMZC1eeVKGlzYwfftLky4DqaZBI1MGMyeIBfS
eGX6XRY/frupzoM4vuPgOJK7f3b9wFofmT9qtOXg3oA/R1tNwGrfCLEb+MdWFvky
CeoPX6NBw3Tfv9p3y9imAr0jPv2PgxTJIkMgnSd3b6Yuxd2EgfH7AoabGdhh+KNh
RUEDqTRk+fDnyjPLAyB9khstHCtXE3wRsxdp8KmuHfgAS2jW7ddDIlEStn+zGYFS
viNrbIwjIJnqQFTitRZnb5mJL845G3EpO0k4C60v/Bl+KGGXomJVRaTXE0/Nqwoh
IVsD6FWzJmoHKjQ0fAGCLm4u9L4llU/UsT4ju35BjEAFLYOy1HiaQuO145zENfTY
HPZc8W06drgEtF+LG/lWZwOubdYr0LTB54JO5irTmSg/ZPG/g2Efco9sdEiyG6cu
J1AdjDbcaGOPGZYMt67e4D+51RyehkS+0UtPfU+E0wjih2D15SAQiza+V5AnqDAJ
N8/NXuT9hrH00O6cihpgrUTHSIi0t9KNFbm4BSf2CD2J0Y7qJ4xYfiCYa9QSWEti
6mZloVCr4BD4WLHJYaVcJbUw/x3DF/4m1pUVUOtuWOniGzvgecmUAwIuHW3P/8iG
QK9PFa34eW14Um2Vu2k8QgRF5qwqjR80ie6Xl1kojvuaA8TH4XS63UpmBLWQLXeQ
BESOgDBVLjnjCdfYnRJnrCRQcG1jnhVKlNlt0+j919cvIDWODMpVMp/aMi7Ke7Mr
d6RWhNFPbCg7omIMWWZdgRqX6K2HmYMyIREZ6bA6+vdymoUwvHSanleJMyjx1wms
Tc7bqjpDOHtBXhoXvnZUHdrQ+0IF+hN9edg6CY6es7iahBiw65DpAxrnrYzHZPqU
msRxCn7EepVsWa+7z9JmuYbOyhGVOJBv4LlZrR1Wa0xymWWSfia3QjlOjHsxQgtk
1vV5GEnK4Z1U8beCtnmtJ647ez9VJ1yEgB579pZF3xS0TgqSKMVCrttOcJqJfBWh
EMRUumFDU3erA3ugnJGCfk9KaiNd8cdxTuMtFx2szBhKUznlg+8Ywl4p42xyrYD6
BwPzez1YuMe1IApvyDZfMbZkKplZO2nXzdBCi1Ec0EE8aEoVwfoz1Q93KpmwOvig
DSYCfYhnqfHAvq5MjyqOXmqF1Kvu/6si7Q3zdnzVyzUfJaQC9BXohUp1GW+p5/67
fQ/iEy6SQEVH35h1JOvPfuNhgRQatO2sLdhCW2zpiw8wt9eYPDnyyy67WT/Ib61B
APYEqBkXkS9Rlu1fKi9pXyGfisI+GmOKzcmzJuxJhYIsONGCL18cupJNMm7lkvmY
7hovkLFtgpiw6f72dU1wGaTCH88VxSsvkTicUPbpwqfiKklG6xghPWxIIjv8v62A
PgDeTyspH+03igG4m94vXb4Sh761bGFbvS1MiwXaayz/YxdU4MmntNw4MnTk7Crl
3/lr8gGfumT6joWHeZkVBu7LCOL985z4S8+XtCnYulb1knogSRTImcRaTfCs+gLg
ouwiq9wPkveMVEhcRqjiXY5FxehuUJvniQ+a2oZOfc5rL4m3xu4hde255NYRhuAf
ZXg7xnddGR/JV73hwkN+kqt8DtCaa1yhNPyCHPM9jKFWPHGLFJcHT84uF2KuiDrX
G0q+nH77W6QBBCwuOYOwZ4kD8VWmqB0J7Gn2vzom4tGCiTHZG4zXypkCs+4J3ZTy
cG1Snvt99Llp8NBjMLyuq0Pb7r0ydL1nSkm3nJv64smpYyCik5DKmgaZueoz+BXq
BPjpycKKa6cKMw921/4sgalPKLBChmoiOU2FzpwUPyYExRNG9A+m8C511alYt9O+
r7niRHIVjgSv25rrw6uyojxz1WTOrm0wZihJKBRd3vvYuZQ50F5QuQjfuLzV7Mt8
cr72qVYGJ671Q+5Ej1m5gakfAy/XAZCGxxpANjHkFtsPrRTiVTWrFOdga+Z+lRSo
e7J2BDW1Na9RRE3aKVWPZey6wQjvyE0E1y+4jdLQEIyvFkFlhhUFt2FOUJkEsBZh
p3VnRBkm92tvWmm3jz952fBtcB7bhte6EH/AzLqVgprtOw6VSkzIbKcOUXPwWqvD
ESjOulBrnxaK5pe8yE+gI8MT6tJNONc4Aaotln3lDNtEBDRM6gNMVM6fXBVS5n2N
pf+3sZ4k9pQEjYaYZ6gwuzckpbFuxs0MfHBIbbcS4Aw1812SzV1HWREAkqMKH+ow
hac1bvhMiIBhK8yyWB6wRSfrySBhGOIXkRairN7yK0QAzCNlNmP/eC7VKvmts6oQ
EHqC1Z08dYXkfTC8VVUOhkpVP3ORUCMUMpLbS52dncsobHHKzOHlqCo5NVdPlcL5
KAuGPdk63/tLTRyyjWhoQffr4qnERGCNlV//WGAFVu2OzwwyF/OPGaKclv3sY7mx
8mSgsfiQIAaMREwDKvz1ZtZkutrZvqjHhP9JQwGb+USwxmnFBJVSWHIsl+SRJz+M
xte8kqVXdvFZGHdie2Do7b8x9zF61YsR+ejZ0FMgclHr5ShI7QoT4IRnDsIe2tEu
ppt5a8ye/vC5L8LZyaKC1U/UhcwfGI0SPj3Pj3FHJxVUAMBW5pUICHmhY9IcHr75
blZoHQVjUqC7W6g+clDayzd4/+j8x9gD3o/n3qrqL99azWS+VoE1/7o9xVcwb6Xu
chdYI1IiFmPwrQSyyJMzzM5jTmBTGt838OX4SQeKG4NUEqfIqErBtWc2jJjxs/LN
nBYcBDnbGchYoTGtIaLqaQu4cSF0DL7+vXTj0vmaBvK0giYzZYyupsV+D8930kd7
MZHzFKroXIHegv05H49a5tzs0kFeWre0+babbu08uPPvpxYtUExoCWVnWGjCBLEz
nBaj7hv+BQrrAJTyqJxTJ22/fSdO8iHDd198jkJqW9A3jPBR7C+PQ6JjDsZsF4gI
Lj1cAJP34TvKP6M4itEO2BTSztJsHP/ebCiBqf5nj79eQthhFNXQp3URV0n7+pXG
GezHgGcsWjND7Gs5O2NFo3/m2b4eCqqgw74I4MGy0r9wNjZj0Cnmtks2mMPqN+xa
IKui74U/HRd3hxoxVTaDtz8t119ZJoRRmZ0OIq+HKpfNoR/IwfciIKF2di+24Bth
JxLQhxD/GKsEXPtnJ/3oniE/SgiKcq8e5IZznr5m0RRKSD20NAbmsXTPmcxz6d9s
JzKNMS/M9nTjgr4Q5ajYLZPCfEM5ZqI+JQq/SrqRxNuRiHRtP1b9OB8XGph/ylx0
h7kH1fS4Ls/oM6Xw75BXEZRm8reopt9YcTt6x5yGZCtRvBpwm+HVWZ59354t6x04
/FjWQwaMLz8J0pV27OG4rTwTlvhtBrxl5RRTEtnJ9LU2dIfaE2c4yXNGev66HETP
JCiX8mF9TvdmeUwmU77mw5wTGLlvNIJxuL3VmFBqO3wQfmfxu+I4BUgIFNwZoOTN
zUMUqTWdc6G0Gx9hbg4g5UpNO0o6xttCkOMl9cNqnUxmB0j8ESvhplc6LWQcoROw
T1uyyDPFG6Tusqp1EeHTIXb5vfuVagsOp5pb+aF4Gf7z/U1uFrCahZij8FmwJYkA
zjbY1fkeUp+GyQswfOK0+AjrHF7zCZoflE2ast45FWA/Sr+p+AHHS0g8TsjuX+Ej
0Ovkax7K5K+B44g4gDHrf3IJecCPu76fEd3CQOISEvrMwWDeaaNXGsgiDpj8rBK8
fkukboKLDij4EI29FHZpj1jSA2RPiFBMXnboJcgj/quhNg9c+LCuCEFXj3dlVyv3
fOaK95ABB6yF2Pv9S5OOtw8EavANBdFgGIZUEB+cNEnYma64c5kfUNRu3pg7GhDZ
zTx6UmeJ6z72cMnOGaORXzhu4yzfNVwCvjZtPyOD0Ajh8sdZJ5cn3i7FkqiAB2dk
g67PbYzUJWj7sVngYx4m6V1bVF/zvvQzAXSIF1PHbnhpK0hnueE7CPGgOE4suDkN
3U5q+Zs8Qq6PwObKyhb5sFoA9G90z0Ez0gcLm1LLxSwSZrBpiHRY7M2ykm2Yumbn
x2uV4KEFUNigYNdxhexbtSHwMu0r5jQsvXP5v4arvQKakEKM8Oefuu8+Mm0AnlsE
WLYjOKK+CmPUSOcWup0gS4XKXVKH1Gw+i3tffC3gQ0Q0uRJDZuBmJae9Xd1R2urc
C8FGt8yLke+rQ6Q1YIDpj0ZbUbGcsnFLKl9uhe3uUHiov0o+vJGOscl0eQWT9cZA
N5IA6HgSH4FMCjXb8bqEC/z8Yx5ITh0IXmLaEf+AjSCw670CCjz/7Upre6svR+iQ
FJkJKzyx+KxWAY533IT2urJmNlnW0h7oQtWqayvk1ziIk/pBNdDBiYfQxqawDLSc
tTt4dljJqX1juBkJYzh80Bql7rnB0NHU0Aat7oZF59flYFfcr5ncOVRBrzpuz1Ew
Oqdx9nCV97gFY5orygLxvoeVZsxCAPmYMvxvY8XKluOoGF4WZyhhLZPHCIlUBoF9
`pragma protect end_protected
