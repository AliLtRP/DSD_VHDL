// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
tUiSAymOqRFgpRjK6YOSlfEwhzQU5py2Pu2jjTTemE1nfYkJgI2/MpAogTZJZnMfGJSdM4pC2fi5
2Re7dZNNn2lL7Nba918My2zobsdZKgUblam8GXGqN0H/hurfY2h7yELyOY49ZoWNTc1ZJjVp5qD/
vSpSBycd/HCur//pEVMwS/ldwO3OxI1dLKUwngvfbXjmqSU6l/py7UbsB31M2J9BGgwXanlDtuar
TNyPSWO23FGfowRRra+2a1obZFeN5CyeP+m2t0Q9V7fN29asK+8z0UcsQ0MAZ5R7DYajBfPYjvx4
NC/m4qcMcpCICFowGsmUQFtiYsAEYa9k7zwx8g==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
0Rtp+x5go5yvpMwV9x8Ma98q3/wMYByWqLkcxRWLw8o62o5Tl22kkKJWoN/eo9wabd1IGRwmYBGu
08F0tXkJNZHpKFnYdvq6ueI9VflhFXOev+2JXUMM45GKhFOORJtCvkTUqxWerWqUkzsGoh2ijGSG
yCjwgHIZKIIAtSyrUyn6ESwalPtstkoRK4DmLQXMUVPUwmRNRqP+aRH7SNsZvBMg2lK7CBlbU8HC
5CEQpcEqMrjTxviBAjGa1ORDpkkT2E+6uemokoeHqmGw9nmu8YSTzs/rrNCQYiAjeJzU0LFaUnNV
uoWUGe0blTJnUqimsUb5ShzMV6UuIhTI8zNMa2MHSQhSkYw87HaPq0gqdqvrtdnRiwZju1/5+5nO
9dZ/I76gCNs3OkfjaHh7Qo4FF8H/d4JuXVS/tR2Ngeivn/BQ3wa/AkNo0cS9rHvsn2kcPDv2QVe3
oVR+WD4iaBVq1UmJQOsyy6n8eUbUWrzP56wdL8jc6BUM1aM39Ll1GLCEc8TddRJXjWzNt729Rz27
WHRHOpJ9Rp8R/n3O8nXv+MnICVGo126kdMcRxLH/DZDlrhPJYJUzC2jOi78BWlLt/0MeZ2Q3Nvxc
6rPJMUpeLjiT0b1jhMR9lltwoe+FVQvlmNoy1VmBd3RJE71u5/aOq2OYGQML5H4wHA5fKnrPJ/h3
RVxGjlg0iazdB8PNvvdE8K/TAYhjMQ4UaPDM/Y18wfPaNy0GW6w8/m4xCeK1mZwJiiheX0c70Mbd
vV+62/wMgtJKz5QkAQvHhPW8KoIaNMuYo0UBpJ2BlOVmGx+v5ilWmmcqL2HRsGFqCmuW/OzSbve8
EjcQaQProD8QFScLYZbeMP8kk+CcekcPxDkry9rYhW5gSXtoLssOokPv3URkio2K6Bv5GLBRB5yZ
QCOo3z/totohfT0wBvcYLCIhhZQGN70IiwUyJWDXrAPhF1px8ehOLePUaQYmhlxcmkrCojvn/6Zn
1o57Hm8aMmmRJy0DcU6IvHJCV7h7o4eYjkqN5LDlpla0Wjw/KVJ/yQ5DfkTCfVOxx2PUMdZQZ1/G
us3H0CSGXqkJjQJww5iI13GEm0csd47/Saodpwf7qRcHtdT9ZVXon0GXXQKIFA8Xy2JKACbAmAnl
B0Z0uhl5LTYkspj4dm4xGqO9guwufjw6nRXucXIq1KSACTbQ+0X92rfCGHMsCwIfi/5zeFBnNzlf
V+VAJprXWb8mqYU4mlIesvvfrb1ajBicWZqVPuGAzaKw/pP2c+JjFSeTPob4319TiY7A2LExwNJH
ikrggLoZYdM51aY80o/lts9/qUc+QSevNrVBNq57SU+fqNhXFaZhk2zOgKzn7nwfsqC5RgKKiHdA
JAAch2ZLpjtyOWkCuy1bgq0WGpVoD9+ySVGllfhscRiLqwpqG+8t/NCriAR66zZyQZY//r2ZjdAA
ojL0mr/rijYR8+qv0axnAfafSvwov2peMle5jSk0Qzgi+/sbrYnhmhXkGDBAPcK5mIaV2EUzSWns
R+yiD65D1WjDiDy2PtET3CSNT/SRmQqjvt1embuldsegm/jSnC02Mh8FE765Z4EkOFeyUpBfpDXP
s5H7SNxbuUey/sOmbACzHBLcG0EVyjzdO7CSoxKI1oqlKUh+LnH26DLdZLOGc0j0prUWLVNcs73f
18vdg1B9+LfmBVXEcZMbURsWK9fQWzKojg7wZ+XpBopw5otWWpzz9UUdXwRw82+wEmI3iNRMELm8
sKhPWC+c1cJzX7vI676J5YqFuDXK3mRlRzE6LpA7FpaABWj4Ce62i7yCGJ1RccpMCdHgGSRoN+7u
OjAX5k642M2h5JbABIKsg+eg1V+mPlMr/SBq/VvirbjCAItQAjUuPaEvOBTVjaJy5oozL+EePxXa
f4S44y31mnjS0RhNsHBj4wwWUqw1HFNvuyrV5aJ/RgJoPRSY/hgheUfu2YiBxyN0TvvHPT2f5zPU
MPVzzjYDGZMKe7X2Y+7eVPmLpZg1aj+t+KrOsO5NIqqAY+pqkER8+RlLG1A80CjjQvhPip/wX6BA
zIuXShxx9omL5wNckyUXDn3F1MzyJDf6nGaNBTZO91QZNxE9td8oMhMhSHlTCIwkvmCnAopl2ZVf
Q+Tl/Sl6WkAcRHLCdaSiQbb3/1V7bofZIw8IWyO+xGDw9pnvnAMNHrfKdNGOe0Iwvj4NzLdJz8YJ
G61Bk3oIAEZRIff/ev/6q/KCChc6DqEiYoilWXd+XZwFEPSKsoLTIT3PedMHMc6tJHG8U3hGQKoU
dOGL9LgKm3s/XZxgVmJqqIcG+XUoFmCm0HcrsLEikRJWEV0JT2RKMDli7ONx8pVfSZ40GnITzyta
KQXz7BPT0WVnsgF7CS1M6yqX06nJCMSEZw4rUmTwl/PXq98ll4CHJqT6ulcchlZ/WJ1XGucBx2XL
BUOPSjXE3+xW5eKedVbzdXyDNWwAqzStxbz52uw7AKrU2fvsiy8k5kylY0gPkMClSF18RTfdTk+F
SsymX++/cbsq7njsjw/gIon5Mv+Cfp2ivdc1p0Jsfg8e6lkKGYP4KUBH1ls/v0L7IUTiD7+6FVR1
OYPE1xuI6iKCe0JWd2WsN6gt6eLu1LrgDeEhMklG2FOUptoZ9z3F1ZEFXn0Eu2MuRh4YhDC5T3JR
VxElL65W6PxvXlvpNyhLV5ZCk92f2EMw+i+LsbxZVBgtlu8OlXiiRKjrWnpyDZab/jScfgmA9MHR
1VBZEKJogZMigi79vOYimEru3DFBRZqiQvwnhvhS17JMiA0cMUon1CxlFeem10wO72+dIKMtVX5w
zVfDIqPe6uSQI0YIwRhSQjypw4gSer1rItUlpXUIEgwCOj/7kbESnF4/HW88zAmClnxz7UQmkU73
A56IaOBtosv/xLM5+464mkpLd1Z6MRe1yWHtf4EJNdgkBm2n52ltrEFO/6EqK6MxvV6BQLl/NWG6
EP7dFe3lwNmFcYkhTrq5bVRMdzVrKQs/aDEB+OGMnKGExK3ONx3WdduYHGJNqZU8hRr/s7HlN4U7
tQUGtHmW9UYzj8eygrAP+zqZC5xx4MUN3CjwOaA76DwS2IRijF8WHHZH0M3a+/P0GHO2eR/cJdEE
icj0ZB2DBEAFi3V+pr+blKfcdIDUzPxecE6x6JCtZCl7fKf+26lNk3bjncl4zXh5VbBcQJVnP1MK
DaBXvse3hrN6yfPmuiO0ILytVLYvDqpiN2Lr75h12KIBpfuGldRZdGgpfhyA6i4bb15Dk/WAWsJA
uPwmJg5rnPrAb6HxUxNg1EBuPJNFZHOI9IZoV1Md0DZex1cTnTGwVzpoa0fWJAX3O+nY+MwarkIi
tptWV1RadDkB7/WPKFmPXPp9mzuPEaefTzo/s4UJzG2Bhtd09WxadklUdtWzoKlSVqMl6aGdRKJN
hWQSr8wvQOo8NI4RmA2oXoL68sswBtvSBXBVYSVtLje7Hb3i/pIdiPYiJQb/fBiQpp12POJtweJO
caziir6djjF8QrHqubQai44UovGKhKSLvGJdRSvFUCiqgqMKQNfCwD/BzMfIirLx0x1yrsFOlp+H
cyrvw8gRjcZYi015PplaKyJrFCmDJT2vO7Pf1Prok+SchDq8FcPLCqL+ShpuYpe6HfDcG6rU8dcm
40JG825tXcq3dME98ohLM39ypaPCYd4HCW9PfHpZI111QB+SGO6aTaAIqeuhv6+HoDNyVXjzjU21
sSP2OU6BGRX1G82DaRUiFJdGGqcMVcQuhGaa1bRL1zTTihZUgTnRMiQb7i4IwjhvcHnsHy2Z2aaA
93/xt5sGRC21wqpXjXIuxdBb8XswO2B+WsTL/pDvLaQAXHjT4jw+ZZT6Sq01ZW9aRaU8oL0KtwCO
tCbjgb13F09pQuh+7fCxhv5agqkGP2bGgkrKcdq0N0Qm4SJZMFSjDdWH+2NPiDRPKZS2nkM0VTYt
VjG+TUlH20ETjqqFRYqFky1J0E71ctoGYA4v0jIGXAYQaFBUk8g8i2VvpcxLAG2ikFrqIkpl66yc
k4jP1ta/kwqxz1dUqPVmiwYHfCnu0su7yFikaqS3hT7Rbdn6oSPnQKZzXiLps+yE3S89oCq79fCW
YPNMW6TDLOEeowv7t3bMbp0OCw8kt2llzkyWJcN8y8vlrMi+M9R1YFUZ6VhC/R/77yx1uT/iqUmP
pi3Y0j4hO/pHINbjA1rLFEg1opiBYxQZquEjxxgad7fwJs+M8idM40k6NK9H6qehvSJMQYlRsTbo
uCrV9ABa39RT/Fjkn+zd6GSItIwgelJ2H2+cQ9mE8EtgajN/zX1ieuxZ0B3pa0VRewqJ1ZwvraLu
l+0GvCFwi0hiuNvCMn3gy5kqc7oU6ktoWGjvQkcbEPmnm+ZJ9SWi3ScItoMctRXaq0LQRpt5IaLB
IhGJXZOhg7su5OxZeuSUPx9mwVh06H6uY3xF2EKfyu16NaivbHMr3tHyCmgWj2Z19SR8yxb+kcJo
caBm5E1g/Z17xAZiPw0XN0+iv/lUHcgovRRTO0sm4ke8qqHA+ZTr9UTRCmpF6Xvjh2XhBq0bOrpt
GWY1GV4KLpqv1goPNaVySrANvAYWmUdHX7RLoFZAfSKgP8a0G/pjkSk5Kg5TouVHcOnnA5NXGV4/
NcoAT4rUWqh+KA5d5DdILz9Ux4mGuA8maRGnUULMLs6J0vAim+E3Go0AzgUxnlXFx6U5s/rEimgf
oSmvAaaPhde7YAEaQLMoR3flZkMvFmixuRmnlQLFGk1mCbRDiVAODY35HkuiRVax3z4KxZhrJCi3
2L7LSwDI/HRUqrB0sPjsb/EB7jVqCLtdJqBm/oGAgt2XK0Zl8QQTyvjvhPbkAGUS2v4+Fds8HnwE
2RozVwzMrVAqgDSfayNf7J3OlKeTZdKi8WWZCEHnDtIfOrBhE7/oVse0SaDTYHJKXryg0FfFNV+7
xIxrFhpOlk7SP4YaIDMEZZHjkHEfV1p0M7+fkM2HNroSUtr8f45xAikhIPQVZnRjzenxTA/tAehG
3O1d/dMtRoMEYw0VW9/wJ9GoKLwq87Dv9jbcTBGIGbbWz03tDPkifiTvFZlt+Xq1ah5ve0CVgJZf
ggbmDVNfP2B4ocILtrqUflH6xXwISJgMehtEd4OC1PDHH5diRABuklIMbBUywFagn3ZbEEJr0axT
Ua2lHtkuAtnCGj+KMRb1BC6/2eBjh6xAUUh7q6kVRLtZjKPVslkLbnk4smwJFJdrhNBdKYyHBy34
OyYsHZ7f8669a7x0KPwCjvulCOL06FT9S7eS2K1nKVPnyCxdkwAUQBAxqgL/8GX4dFAc0bNSFFSn
HSNK/xVYdsMt4EsD3W7CnKzS7VdY1GIUUV6oKTMX2XDAlw29suq3NA5fj95E4vcq/FAvh/kQ1fBQ
fx5C5twI7s/FzB4KweVpAyQhHDXPk477DYb44UO7GzYj5EtncWQ1HoTyzx2WmgO77DXgtHiWPowN
NJQVu5G7RaYMEw/Z/rppfw3OxB0tuDWJl8jJuz6H0ABiwpPDdRA8QbY9K8xopvzevNUQ+0ctqpxq
wn9LVnLJm0sqormw3hmEvBaqcYf8lM/RyZkip9DdRlOVYgL+xF8H1pPVohe/1AcLMG30rAlchG9H
eWhiEnLSZFyW897Qfp8p42l4+kSA4MM34hyfzjUyM77F9r8MmdBONeKhI44bU23crDmE+ydddcyV
RvLFreKb5mD2xDUdUTJ8nvC76aetxYl2QgTNkPZs1/IRlCc7A6S3aATjgihs/A9jbZSXBAk/1Ref
GDiX1dsO7+N1sNuTwyX99cF+kFUDuAZ5GQWBdvF8zZG5Nh9cnQuFoHCeppfdMd2DsgL18FMp+enh
VbnzRL5XJXH+SEL9xXNaunWtItlC5JSxUE5e0sXNwW7tDf+EX4+ED2TwYU4GuQ2WTvqpQ8to1xy9
nbfEZxpcHJhu54CPEpt+26w4XtNyerE9IDy/WLuZkMMhR43si/LkzVrMDWDB7X5TFc/ZAh0LZsEN
/A3RlPwY1JzKCpI7lx4Naym1yMkyyE3waAL2B3TM7EWbuHt27tcESc+5r2h32dmEEnfw/BODErN+
/YAiDMrlIMu7GEQjuacDM2RIaJny1jYxxYHUhp7j4XJ4Nzhgg9EYi+lWTsg/+/7iwViPL8lqKiVd
B/0UDfHG7+dychECTQVSlyErBFqYPoYZHiwgItNbd/OhWbH7RCqFSvFShzc7HcJ24dmZ2vE3Y9Pp
BOIoeIoFRy3weRGErkcZ04X6Y37PTpAYfxiofv5QQbWpoq6ntGbicpV442QCQY0zQuxN65zH3ito
s7etcrfeq5St/FKil4OlLiotJ9X8w4VYvo9eN1f/h5A802KHMhKVxT+lVdfL7rEBlEHhZBwe3cCr
FT2WbtDQDbZHFnXJc5wPpIKW9cJQIQ8fZrtBLPa+yGfiMf5G43hm6kdoJYzNlybzZOnbQtFsgZ+Q
3qHMhV1ikagkDZuvjBt2GdE9e00HAg9vpVi/qf9Ti8l+zkicYm9eKh6G4v06GgiI+w+a/LWqHqfA
bW4bijWS+Rg0FNkrwsdsWSm45YDuz5WkuxH7LpL+8rlHDtkEvTsHCubu5R+LpqCHmv1Q5x3OYD1E
yi1p/AnWb2fBS2tPL8VL6btTZUln3EAgndkS2xnQEjU/Lrz3nw9PvHsL3GwEQVjyvsOp8mlTfyDx
tQZr8+p103SFKXtpUm6FcEcTfbMPZr5PksP3hYkC70c1K6XZkDne+KZ6uNbt3BOjPAvcbNAnk+mQ
PksSSTkq75UkYWVH3XyUyW2eCQiOmNY/YSNq7sqWtjTT+Nw4Fi6uTwvl+Sfwwyj5OAZ2OSZ4GuNF
mx40QK9fDDCcfrRG0wKG/HGla0tYGsL/jOcvWGZVYH/Y6EWrnOt66RyTdCygaTrsqc1hkDueYhW5
+aQkwzNbj5Q1jZXdVpq5y2lzVwpkrnqLmTZPjpFzgwxFnTwb7223lT2VRCqj2hVBBI9SC5FW3obQ
tcIMNTMNzHosm5ujlkV8TDbFgMp3YoCCRIZDTBCtVKTh8W7cSkFaTGmEYhsoUfg3ZBswEjn+hlOI
pYYmvJylQwAvy9wjvQCtu/PzTpmL9UURH9l1s94K+LYUP1MtuHQD3ZyjUdPjzlb8oQD36f/fCBJd
KgjZzJ05zu0vIWI6WHyx/Ah9u7BAQgnrok7HPCl6YIguTLQfCiWcPCs9kEcqb7Qy0YGXENsiu/r9
nKgXsr90f/+0c/FJpiUl+XCmsWb/q0pf+5Bz5UzXMQuQhOBOiGniGp3ud9gLY0JQKHYQ/rPn8w4/
7y79exig90STQo2dQcYXak0u0/Y3nC6Sm41rOFtY/xDPG3ancC6RCukU9m1w2jmE7zqS0eBgcihq
UVTp4Vmqb/I3ttSwvZ5oVjHzBnoiZi2QD6/PsxzjyxwV1/KGQEyLcaQi6p1ulue9Wij6y++jytIM
3Ctc+cRrWR/z3oHLn6io1U6M+6dETTrMZ1io9eJz2KowD7dm9age7uNACDK9I20yo36lGmkAZZGA
D93RV0+fD1lU6x7VPZqH6LhtUZLZAkpc58ny2OWAt/0b9C5jZ+0hcg9+VPRJycejMBwjd/WHFL8P
VGt67ltmO4rCMX5vWPrqfuLnAuOaxUYeTsmcOoE4He3EyQfCXWALL1g3syiqs52/4vvZnSekEqeG
OUs1KDPkJfuJXMT+RHkAZyqc3sS+evbs2Ui27P2VY6h+BMaqFHlUd2xSQOy7s1BG3RTYM9ZMR1TX
9FQ/OqDDpAuCv/EzAA3kWwqJQLihqJ8O93Ra3ZB08TjXE+38vx8cF692Fs4ZCmV9+4CZ793zHvOf
8/YPXMCr/WQnvDwqxUi9eACRaOE6maj5SXdM6AUOG/d68kLtJwk06FdVUw5a6GM8t/vwG7J1xYs4
tUlQdk7Wq7Y20FTc67Vim+yE4lQ7XQZPq3Ee2UXDNH1chs6090csyDq5jQ4NUrl+vys6a6KxPdl3
GrF3qbH+WMxB+NuO5E8vV1WahjVzFrgIvr6387XzfXo1szbYqeAh8nVcRUcbku4pmI+TvF6/iXJA
ndYI6VQBZ4aHvsNNSsR8FTt1rngHgKVI/7pPqj7BA6O2+kq8xhjEVvPCaxosYQDEu7DCYtlEa3oh
K9Hcr4YS1qqGEBJLJwyPuFEyXrz06TWoDEFPzxHU/NMejTqsYf12oAAjIWMzsG+kKDdQCwx5N/wD
amveDHkMuVqluchs1+lQUpwPs5HymhckFagdMBo9GTPmDDZCL1rgm4QgoS/Y7qY5h9U+jKQNfNFI
JOmzZHLN7X9LdpoprKKoLP1lhVBPNpUiA4MydCxyfvEohyb9ZFEz8qrp4d/LWt0dqOx/0e488p1d
e6fPYdbLD9tbzZsy21TADUZmtIOYc+TrOmVHG2wYuZQe3+GLO3TfZOBhBRSQLZQgLFltSeit5p/8
b+/momcoUZ12wvy1wQJ02R9QNB/I9AAXi/LzlsiF0082wXtpkC0aQKGml+RMl5vGz4a+odlqPQ2f
JyWio0N+vTrL+M3UDIRbk3E0e5uqPt6+XEdLyfoJ4wUo5qHyZc4daWPWfMC92fHXmb3BDuEm5J1C
FuTiO8CIjreEQzNB7nAsFi0+8mw1VDVbBh8Z7ajtrnHdltncbHaipXWfrcdT1dqDdArwEwSWxHY5
CsdnrWa7idBu0x6iqrZnvWKAG46EH4VpXhBBcI+i8jkuMCOeI+kosW4ambSlpqn+4JaFKV7MADeF
CBf/SGDvvpoD7afl+AkzO8PEUXwPbWJuK6Ns7qNv19N0emqQqS0olLY6DR39Y1rG9woyewV5C+0Z
O7vJRnv1rzEp8gzGCyzCwhoi8j+nF2NXLaEDpb8Immxt09mmdJ5p2nSKvcgj/Z83aj3VAiG92xUn
AOIzVYC5O00811oOltpuKXBsyS7f8QmWxNLg97elnv/Z4rqi1CbyKNV1QTQWAgpXxMbQtiLbUc85
nhtCbJUjg6kZ4FUv+dQVDlu8pXl2GVuqJKoXVwmv4gB6bYJhHRZP+FYmMH+IDzzx9lNbSB/CZwI4
AGP82+HjFHhqidnXszKN/hbWen6RTgQDEx7Fc+SulYmyH5SgU1Ap7XtZc8YH7TxQKwVc5S8EmRSi
oSKk5XHWgeWVcz5m3bUKSOQq8VqD66h99Ugw7XALkVeARwGGZbkOmvKjWkUmD9lF35o5/HQ8nuHC
XpzHEz+QMW2It9CdWgfzclj4RUSL0UAWPXtOG7NcvfKoJQpEHnw1DAGzNfdAIJzp61jA/pfEZWQn
i9PLIZjMgqMFn+4Wn8mnN4RSqEycC1mbNjk7llCXkcXvXRPNfNAHjB/Q4sRdscDEarU+1FEmvIT3
IVWKlEdmMWJ+M4nB3lL82O7FV3Y5bwzQoFTK1ijos95aMQUllJ/miPAj+nB4zKDH+Dx5eSYSYBwq
fMGljwNUXuWjpTOg24l6fleYC9w8dAZDriz8Nkeg1aWpKUMqkXtVfM6e1LQJPn3JTDiAmzNs1oPQ
m24mSyD3Sf2BiLPXlELYx5Qo4vvuWIZGZpTOlNiUSCx0KC4F9IXP7HVcApxX8ZCZhb29GN2siKfK
JEYz0rla/CF/wxujrAW3Aqud0Lw0opF9ERRh7vvs1sm6jeCKFwFbxU4fpTlDq+Y+1s6UD3WK3E0z
G2PP5w8K/7wiQNmLksbT6ennXo9aj1JU+n8UddHk7XaBaRTGJwngBx89nS4LmmaH08PxqDfvIB0X
GU4wv9vAb4Jah8zhuIFgkFjQa/2bflBJDW5y/DXAnvP2wratVP671vRp2TlXeNF7WSq9v106GmI/
4pICVvTFhMXoVtvz8U2UBIO3K/RGiL9JQYzKRlvbs6pJTxkwjY03JG8revrKJ3lvtVccdb0Pyg5M
rgv6WKf1FvQ/EztBRsPC9WNi9FInj4w/ON7FC/8oHhX0ZqjuIV+ojWD7/4j2Mmk/aMi3YP9nxBy9
dxDE4hexHsVe57CJUMh4mTZJ8XCqMBKqkO1ixxaFHiThCivCuX+/GVHe9K97NktH7mtuQBs7lQq5
DS7Ge89GIIKzHhgqba7Byf8FQLouymDFKhQTy0k9omF2ojUqGS5Huy2aq5p6B6VQPXgH/LHUzip6
K5Woi3Iq4OGsxy5bp+YtT4iEc1qxvWY35HcDs87SqspI9YeP7KZhTZ/b2f7UCcX+Q9M/1ejIf1V/
PjcLU7q6/SivAVgxxpDYBQaPsvN5TyZr41qpf6BEWA1l2FAXPf50/8KW3qJIW13PHLw9yGdm/Wdt
t6P74fjKrAWYEMUZL4/YKlr5PJl/N++Xhf64JNBRdtwONN+FRj41tT8L/IZaAXH23IfR8yCG47EE
AULp20AwjnwxmLk4Qk+Xubp1ctCPMJWVIUM2RsvlYrpGuJdEAha4+/8XSU8Gw+9fRHJRKr6mknpx
oBBnk0QYfYliRMYmY33uah9pbFy4jjzYRblSFb7VTLMQfdOP901zqpdpSZ1j5+4puHXOyXQT8AI8
f3CTnNSqCJO4ufi5TFg2sx1NecemPWMWP0Vu9mUEEZqhZw/8Yn1US8vNj8kbN0WRCViuUsAxmmVj
iBjleDMHWWgYBGgOZNn8DwaDTLS94uRQ5yeyahVU5AhVFiIVJwd8EuweZGJN10Wmoj0ckmGR8MAH
FsMUIuStXhp+t3uA2IuyPTtuNyr2asprNUqhs34HBBUjK4614gWsKiddhuBfZTqr+9NNxS/57ycW
5A9A0ntkwXlyqr5jD7tVtGLqtzMIaHNkZydX4JF9LE8wzjCmlbp9kS7AKkVpYpGfpMEkxmhQsTNp
6FAS5e8XsuQvr24iawPdtxvyP8wBV9lA7hXsooM8iYZzX4khrE2DrxNY9Qhn1VXUJXx2DsuLQZ7D
2e38vlmtMKg6skpouTzJmCOP1rv018SmS2nQlNxzxxK7JjMPoj32XF/XVq5kpPH9AzV3gdK844H8
Jzp0v72Lv7k2xQyVCmBYQ2ABfxAR5VOFA55gP8xCZIG73nf+fGSInOFJxojDQIu0YlWmuhDHiKXy
Hhfuuxy/X/mJ4hpQvnkBCfFh8usKc2bspO3BGLzMCXojKtFkJM+tCm1A8YrddtASzR+124gVGU7X
FLQ5V7BwzL2oActk+1JSaVWXaMvoG4ev6YTA71vzc/bX4T1yN1Hrr1CScLkg8ENo+H9VlGcVFeCC
hl+OGGbWhdCSCvTSEWGOrbJWGIxd3JQi4zXqxzQ0yLtjOPAN4zlzkNWi/6U8Z3+eTu4Tx7UuSSVH
ueCotj6SgOahD3vulu/cFMzhmpJq2I1yo+F+jiMsUnV27nOJSu+JoZlVTNcj5/o0Y3h7ONo66mwT
d/sJLZr6U5vl+aBTpmiI26ATj5xgciQ+MyQlCcys0DiPGjt5md9sZ5AeHSmBnBZHty09W4+sY635
aeqkrkKaKerDMEMIWjWXKUhumgjk8Z7fAIL+BJ4rzmRuBLq3HwbaLkd2So2eIO7tgkRfHENQXWH4
4hT45YqRfcwPo0PRj3TelaKcLdOG3rg0jg55P4OydCg1Jeds+GmMbCmMSqcHSt88lcWSAZTkks0B
vOKW7zufRFPXfvuB2SoQiiaxvjtiVd3gPL17gId3cIFuTZhpTkvs7OLa2D9Ofj597L+VYfo85LRY
ZqsEYhgwT9WTV3I/sV5aSh3ic1OqZZL6qs3K7t/+AGVMCjEhLMGKSJJlsxPWP7W431MdQu/SRIe/
vFhPbW5z3ajyMECS3zHNuUsubWvkd59wuyYGG6VU+3yvWb8cq1HoSoL+JKHHH/eYX1b0RVJWqMxy
Qf7l+levNDFgTRn14gFBC1fc9qDM8qvOxEFPYfzYX9MBWpoxBjcAtDovnWOk9uI/plIvtu8Qh5s8
2zT1yOMowf0Y/iz630HOj2bS5rat5JM1Ik+WKjb6BwLfWMp5rc4pHjI4TlCTD7aoXXpYqrxTX8da
qrY913u9o3yKI109XVcLPtGqyfHbW8Mroh4A5K88Rk03uVzGSJgDs2ADLn/mZQ7HVyGI85NJlDo3
bUknXUkxQ/bBt/vBq6ILSf8KHcDGyqUNNIiKIauj/LuZkO4nhsejhL53PDrKXLTfon7m8M5urCNk
34ceN8Z8MxlRAAxummRsyXtbZ0i83wCbabrqD5TjOOzvGkHhIe2sapiv08HLO0MZ5ExBqys6fNTq
hxkKNpSezIH8iS4kBVnIudzS5fnr/MrIzbniwvw5T3N7ZGlgoF7++phhhCEjODNgst92yVsWQ63y
lCN1e1CBWHvqlyLgTFwh53CG0oIF4UaYwXPVkGIruKr/ZBiVvgFN7yhV7hiaMQXZCbY03x8Wn/0P
UFEMOrK0IMmrkVL5z2IlwiZewPYaA6eUq6mo/3ru1YLVr6a9ru855h6CioFpvdP9Vc7dikXXMjUM
C3ha+W7ONtAd+34ROIQ2D4l9It59imVVMo35rpRMnVhO6SKPFYMsegkylHd6SDwAp/Z4KPCUGSI9
Jy/ZrYx40wX9A6NSXjSCXgdyS2bC5bp2JjakJc683GlnseA9YLJgVILYdApCbrU+HjFtdwouOA8m
trvyhU/sJSJroRAwBaAa+fsXL81O7YmRRFyXMZ8t5gE2xYDR7zNEf3zwmHS2i/IrwpKYXgL1f/1y
fLfMLYOnVJhOdq79zbZ5Orv6PPsp/TKsGSpRqKDMqWXvuf0fRtu6cc6Lfq4bkEA5OfQAjg0y5xz/
mpLr4MaPpOMy2jZXReWcyW/8OH9IEZH9FN7YWUOwNs7e3TO/7mFffSI9PpTx6gPqFProb9IQaojC
j96cmlZfZ6XzuZdwESBOMF8B68uZVmH/RoSo8J//Yhvy/6aIoU4Nqqe6vn+y1J3dLOipVPJ1S9PK
EM64DLpaUnzN6Xt1OTzlsT2MGhG/jqRJ4m5tTQ1QsWiBDHLHxQVcujFSKfQJ5ZVww75FbanyWHBt
hJbj0anixLHiGAfmP23Fu1tVCMx8AYMV7FF6YSAfvccxoFSsjdYFhCeM3ASmLCuVzfj+3XbIgti2
gJYVnfwsjbmO3tsGf4qRgY94qBLhjr5Fp8s8CtSkfwXJRIC89fs/XEleQiDjogj/E47ofIhAhvlS
sMV7/i0sReqOrh8twoCW5MTkAwnEYAKLVXIS6E0XIq/BYHpAAN0u3iIQk7bo06dAfmhE1J4LX2Vz
oykNaK25u1TccvrjodndA61fWNsEBRDNAFgOGVf32vIy3noIZsvM66TnjBBFv4rUvWzzcKm+pW/d
C1ldY28v0aMDnbFaGRKZlKvgHNU+R0iCAgVHkacP/HuQdCiJCHLe5vypJx/loWPNy5lm44wKt4EO
3ufKBGRATDH3wYlkTyVaOAkDBOCLEl2lsHff2unN5qrmG29WQrnJ+iLKhDlrMVBgi1S6g1l6TOAm
To2dy+nwweC55rjwm2LOmTtOCapq6iLxa5Q2pnnjuxkJhdQ5onwpjSG1TKodrloAJ0V2l5Lorb0S
gOVVah10j2Nd5IS3slnVYbs0vIcs4PNtUpV4SRBqvYhNsnTsCH535pnDa+kVRGJkgMukquOZdk86
7IkgvaVJ6csA3fbeh1muB84ctmpC3UWc0FUsfDnRC5r5jWVa/H3JoFBu10pwGFA+aGwR4qjocafi
5dtcrP1sUOAEC6xEulvq35q70l+yfk/h2aAL0KiR52RfQvORml/HmVaIuB4/8tysLtWcMHg6QUFJ
zEllCqjMXbw4IQnLMK0RN1vr+ENUablotqum/mnQNVz0eMUjQoeNqPEkvX4LVR/QcCAuVSQKLyB/
gH4BX+giPgx99WIGl4hMoPjcG6oNRRKbaakEZveK3szNlNr8dI79aXiI6QAdwlUEIAGnp4IaEUHn
QqahogYXRWlwJPmKQ2sCmM2MUoubz748D8NL/dvJWVNRN4cRfYOy9iy/JfYOcYqdEfeepP7XJpZC
vDrJH02vJnXg18f65c1dFAgPYppqWaUf2sg1sb4SuFD1z4fZv06HIfTTqc/uYGwEzoXT7oFolgRT
/VgMt0qs5UG4O77naeMQOCoIyleD8ErSq1EAtWyZg2MNvLd9hDWheg5qLk6Z8eSufPd2oA/OPDm3
045jbVQIXoilNDbfI/SCU2s4TTmLNMmoz65kyngrzax7W/alB2G3As5ynwSl0qX0mumscYIveX2O
VvEa/vIwT+LCAtZf6YAPcnsaY35DnL5zZ5qwr32guCreYFmRCKZR6sM2k2mliBwkRfYkXP/odb6e
ppAP6bxxymXQ5DCmv7Ajwp2rEM0LNtbgArQmhQ2uGPTBCwrGLyTI9uawOkBoC+JMa7uaodesrjyc
Zr7zPkjDX29lJVo+M628bpaLldIs9lSvDTs3Yn1CiIC2hC01+umOrFGD59lwQKckr5vXAlXr1KtH
nfpJsFDX7e/xgiOdEwuyNynmushjQxLShZFSXrOfYd+WirxVkdfovW1fBNBPhlN73QHhnsGpb5Dv
bEf/9o9duSjZRCuCA3EGNQ5yWoGwBtdS0/I6OQ82zXUngTvfCUzJTVIffyA080CjlOOpEFBaFz5r
BRwWiQB095QaY7r9Ul0JsxZb+0idwuztiPmhQXnAjxeSxLV8T4vYoVoovqBzE9CnuLPEyxKFfhgq
nU+vJjc3Nm6oKOI3aPsbt7TXcKg11uq6Q1l3RGkpqaZgvKzZYJQHdVlykzkNVrmHWMLtQls+ZulF
gkWJEjznfQQ1udsi9jeVqPjHn/DIXM1xKkg1+QvHkPIfeG+ajJr/sNbPNpXkQ9jYYMGkLKLviY5b
fcZf8cWFum672fshgmAe5KfxLoiuMP2AKabGpxiFveCdBYhqDgRUkbtya1+6bVUEB/ehEOb4e5VX
PtSFeAt3icbKBxkqQRtTpwPdwMrUnSLbKJDOiEPd5k1EwXzg2Rbb3WWrU5OqYCA47YQnKbgKQV+w
7kAN4L6pRKzxxvkoQ+8nI6utgEB74t46vTObyuGbArIyDJ5u4GiJ+za400N/DpY1XekVzlU7jato
XFiSpJvxZryM1Wc9zwsbCs8WDYo0FRuN/Eq14xcy0MNwBySFexVhMgwm691qs0XLCj2aub5785XR
rzSweRV7Qwm70zif7/e1sdW52J8r8JxG2bZI6zBpYfAxs7oxkrLpWEZ4xQ/O1ULqJVK1XMU5jcxg
rqgyjDW0UZ8tamKbuQAQt5GCxJw8MawKsqHy6hBk44gFRJjt7PsxJnLRNyK0ingxVSxWXRX0b+/o
wDe/THqBFOBcV2zUm0C28pKpF5y4Cupvy5Kbg0X2kGAA6e7Sjb4293C2LgmHgE8pW31A3GrlP+l4
lIFzCWmVzxVRWxY16gg08zpviUMndHn2boPI1gvV8V8a+zshSD3WPGItEU57OgiQy5Rko6+hF3Qq
YdlSX/vyK/rPCjNi3OthttMma3Hri5W5VtL/uEew/qrKwy7tWQhXrpQzwpGiG9s+ssRzaT5Y+jB/
KjpWl9YTc3S5K0f4t1k1bKbSmVH83WIVjPsTHQaLanuc5jkRPZYqA/cxXY6BHCQY9DrcizZ8yqhU
SEhZM03htuT4tXiSDHqM9iYue0EgButlIC+vH2wuD5zFcLOjiWDSvt3BPH8U1OrGKn8Gjsq5zj2m
vIjCBkmuKoRL8Jo9ki2QlhjWsurNwmLfuC516o/rBebHf318DX/JnEQGHYFPx9FGW+ZXU6Z4e1eq
URgHbKYg/ivOoYU+MYgFUuYBOftIoXKAJMST4V3Yk6NABitgI34Q2k9MtUCsMKymt9m9t0ecRiel
2+5NXhyns7XYFGTNbEPcGhPtUvat3nUOrnzgJKYZ8so6wr6hFv/vpIwENLRTSTMTHUnjtDbTrC9y
XedoTJy0CT/LNsyhxdtGLQ/y3x5zJGpeZGMP5OvGpZuvGrlYFRIxGHs2M7h9Z/ReEHLfK8XvoLXT
K51UtcfKP/b53XMem05KDvwolp2UQOeTLMx2OzDqs4+06nKz45wtM2xRJKERCNAmU7sKVodID17s
D0I7l7owe6Bz72DGOIjtMXPtkAAjcZ2iPz9Egda16wThXBngioqrlJiWGxYTgD5M+nlYlYjqZWAa
5vP7yQoDeRckes11YEz3LLk6p33E7oCuCVpPcePWx1C1Jd85ItfaOcJIAaIBEXl0Hh6Mf1XEbzS7
35pxZ3bpyrbxYWI/uAD3legNlL0wgBS/GjWRZQxU/v28bBKgo6WRyIMMCRUiwyA6clQUwJWH5aRN
l9Nf+OmDeou9jY2hkVXR+CQPTE30NWOHxqZXudeWuGy2Wv6/3kpEgvcKSnToXjgCGcluW4UcdNPE
NcTCixwa5xsievCGwW021GPSfS3yHaE9q1wrBbELkHUmp43g7DMl3IfeAiFvoYmIKQftr9kVsR8j
+LSvsZ/ivI82ePmTAntqLYhD+mxk3CHENDFFn5rRg7mfX1fy8TMD94E1G+MwMjN4UscDWPiakaI2
JrH+NilFqNhwVDeHBnHg8yicL9F2Lb8YW/47jxviH/WAkcqWd21lBUpf0xi12Fbrzw6XgCPqi8cI
/kumfqM1DMjgydWSYI8HJnQrwTgj9xsHqWpE209wVJoTo0dexmMMcyyZ4WCTBQTlHjtmDHzVT64v
vA7osdpE7I4l6bSVPElk3OIfmKZyXf9E72edvFd5BUA+/KO8Od+F6HYsCqN8yAZcYLPRE1cv0qyM
7T5srAk5sopGpkvGd8PNy8O5of8z/oq+SI1501jOxqBnkrr1fWfoC4xbqs+2VT00t84L9OQVOKuN
D3o20h41EJL3JE2kh3A1a3xALQ3xaRtmLP09Z7q50LHbzZsyvBYvrAsziwnsL6IJuuQzgsYxZtaU
R93K4MOYv9Kzxwfm6ZtAcJz51Hums1OB8pFTBzdiIMGfkWCNc6Kna8ACFS3RBvOR5Klr5PM2lDRD
/9GvgU0NX2mONilc7u7ptVpfYO7DaOQDf92wNeeHOYvcrfWsKKN2BLV5mrAPCiQeHpXf/ZIKweIz
m9myM8mZZL4MpDt8r1A8j7FjhDV6Pgpzj86v8Be1GmH5szUVMfAdfWEKYK6mOgqjWLstEyoHwAKk
lLYPivWvdim8LUL2VyZBKcPd0IebhzffM04yuX5TKvxh4Ts4eXEH6UGRmS4ePU0rDQY28STbRd3p
r2KgBnvUQ3DHjyp8oFBeER0IcnTCrUWcokW5WNWaozr0OQgqWgcep/nlUe/b4t02ajxosTXe4ZDt
sVxBbV5rT+3X9jN5tNtqNwT9VxswTrBdDLkyrrDP9iAjjkVDlhi7WS5I6shyC7GzLnRH9kFmsOOh
1n1safv4Bww3/pmI7oSLBL4T0aDcYsXmkFwjeRoLvku5wGrmdllFKDNfFE6wqkUx+v4bwnfChNoK
VdNNkH+ZgZCVUMMYYOmqsEjxT5tY6T5lwvBGdJAUmPY15mAJP0nnbmbTges6iBERtUCwsdDfYjC8
wZ+DzvkAfvBe/JlgH0qHtX9wydWJ4jCMSjeqYT2fHWLaumLuDrinu82qyTEMmhfiEIxEIGNqSL5h
+zD5ARlIAxAfT453JMkKSVE11Rq5jbaqKDAOrYksHjAIhSJJ/JupiMH1M7MnNC9Eqjzdfu820DMw
MQ3Rwt/QPUkZvA75c7Dct5Y7uG9riD+CMWw/7VydLivhSSAkBHDxTX0f0zBUtxPHPYYZDsC5R78B
TQRqFLz4DDEYHgPOAcsLNWH3Wp+J2BdH/Kwpt1DbfMRNeDwPWLh1WnJHrj0mEjnJUpu0G+G3NM9e
8dNPzQIIlYrtPSCbGqJ1ekKqkvWZTPudCfrpomua5+Y1MnFXbn1zzuN+Q7rlU88RJKffP4y7kqWm
LzFEGv/ycyzAGdGzVvbYPIPDeEm9VnBo1JB+fqHMo2jKn4kj2aWSwCvdFw1SjnC1rwAG9F0ePfk4
U198ZL3dQORnD+kCcn480+iK8mKHBkxDGr8vVhUIJtGW9i97nBTMJtXMky0/vnfP8YRdYdkSfD3Z
JcpkWWSNBlMUpNWSSHIUuUaMmnR/eiTSW+0WHPbGIUv/TqokCcTHGvuMYxk1C+K4KIurApFTPLOd
blvgOIpI5RnZOt9XpX5+qHXIljRi9zj7pGYrgFjSuyxFin3FQeqgaJHxcz8ZTqyD/P8UERmbvzm2
PfA5tenMkX39u3yYEVBy7GQzKFgpDsNwLhCDFC5tUyA7jzqZXHPwI6AMQcI3sQ1oJFjuu2S871H5
eOBGQ5Jhnfc1ZyA+16gfPwvop6O4TNsNe+7/6adlSQMVUt88O19cO2lXDLwTsTD9OxFBRG2lEo6y
8L24x74zDd50/eL/nnzSm+rz8AOLGVzbgjPTUiF8/dJwhgC4mGiQlWsUEE1S9H1bLefnkmMkcanJ
ubvqIS1hfJI/TJ0o/c/NyMsWW8nXzXZhhJWX7F4x21VsTpidaBktPfDjBo+oVDilggFQymAMDo7N
DsTazlu0vqUQYJx0IVISLglKMXrfUkPOmdNfYqMDyQzY2QDTc2NP93DydvzethJcyQWPkqRH4XSj
Y1fqvu5baU4n3BZAay5J9HLn2IYxe4CHs/eAc62KRxGVqt8zSHK+bPa9ZG1KdaBZMLj4jEBjT1Cj
AF207B5fpvAiwd1yJqqDvoKIE/2TbnnlgcKmDqNbdThGvb6ABU0uMk4zEdPng90UANgnBu0Jk+ib
3IEoM/TOMe5EM4I27RaE98ZkdZms4WrupsQANBNj5uEzCdn1ns6hZXyCKZOp5lkQHQ52Ymxwl+Y7
VANouQ0bHOj8Cky0Lnebgo1yZAFZuB+YSspO39naErnmCVgH/2bWfi36qpFVlXUVNW4WY1IGW1yV
IzioDAr30VhrZSvnH6Lo3dBCOMEXCfLykRKH1ksP0iKvfBBal1ux1PVafR7cuUwKi2WGxIn/X9jJ
/CPHx/41MVVWIDmRotON61J+IGaUFQDq7yZ5N/xHHaW0g42SCPL8/zX98TwZjjQmya04fTPlNp2E
ZT7ooVk/D2tPTqIF6HjfcHymO478M1AoL1lJYtenNxmEiL8hg0E7N6uFUZlaLWUJQsMM41koIogH
8P29C1x3GfMRhJIVmjlRTzGWP1fptTbyJOtaJvroxuf+/c/YoyjjUC4NIZdaBCA7aG7Bn20SokMo
c8HOtRLmZrWByUOTxfTxeK9BRkVVGP0SStGnD8eQoW1rzZ/7gjLYos3W0VollpanKBFTpCWIQA1Y
CU8XGJJCS4bJnBBJZddednEkPZgIuGGyTPNzxdw7mBV7SNOd/jKz081xI+rW3wtB/fw/DukbFG7X
zZ9FYxKDkqMRRQBu9eUubdOkf/0jvI/9UiufSnhAbBIsEYoBdyV1Id03YtaBnuiT49H3X2cMAhlE
qDCbVrOdtKyhTpkko+/oAzqoECWkGu6zTe9YJRtnCc14UgXSJjgdoNGJ8i9tDJScMkr88pKuljZP
FAN9ailWBbTeZKXsQ2GdXJluDMfUBKie6yH6fEFbBJjzveLl8u4ABBHBStqzYDKq8r1lyOo4xRDK
sGNBy/QszNd47FzOAYKsP0DFB5Y41RhwpkNlVSMEU4Qj8PvLGc+TGrL4wrQTat6P0ADPZl6U0eiq
g/iYM/9O3rdSjKF6F7eR23oXN8PyNYbyE05UWUNsG0FQDziTwTLummqGrYLCYKgGi6WlLduqsQVI
R17oy8veQYYjQng0ouHTShQpaeRdeiZOjNJMQueH7w5POLW0ERMjG89ous+PcdEQNH0qW2cHIJpx
BwQayy6jOITMljLAXHsD35bXKbcZbhiLklwgJRXEQVIGFxV4wEbHWl+RKhOgn2kmHJDzHlYMuXI6
9u5fT/rjv4H6dcf3fomuEeH9xbBUYnKbeBKPsH8tL0RzP6RmCYLjE9p/KNkNc6Nd+E+LYSAzE4bs
5c9G947Rn8Kd4xtMjAF2vd+VNCC30XHMNh8DFCm+jUugH6Oyb0L7MktZTxJBEogo54V0jjR126Ez
wx+LsPCVby7bARJl4byCQRq3H8No4AJFtsgVDeAgOl2HCZiWvbRL/cmoaBNDoR05I24eiLmSiTtL
I6ldfOU8s5FY/zxMHwuNgYv7sE2ThZrxZkWDK7Ax2vhfyZZj54wbRS9Qhg07eYIVWocgcI1eoLai
YLs72gl1jasEmg07TDiOQx372UHqGo9I+O7I14vs85U2XbNi54vWGyhLPb9jcFZrDCaOAxjHm2/c
guFSZQsEPV5FoLF51hQTtYTN+GQ8iOdChbEWjiOBdGkmaSmF8PBWez/dAixTHd5tPLBeAOaWTv2M
5ZaHfWOvMOip9opNU++D/Yi+O2DpEkOovtkuMg76TFjzNhI83RrIouanH1bYQEtRg8bT/9rmPE9n
OMSP9Bcn/Ah/pTsfpFYSGvtq45pExAeIjXPoYvuSsIXzJ6uS+Hc3F+K48JUiU3FC2FsrtGWNF0sl
TrOd1st+FcL/nyNx2GNwjUkuuOECDRp5n9TRoEKIscy8QeNDn6OptWcfBv5hT+epnHXFcPLnuQd1
xbBaAyv2Ih/aMvBjNDLL2q+Vc6JeezmPdgpZ726EnMrxZgiKn0bChlZomSyoUDaTRMkFIcHJ2UnI
JiwJHYNjBzBoeIyFjPFbsq46mAgoTc+O+Sz51zc941ATD2vTO4PoBnkD1bj5uiWHNE46Qa2YOYKu
0WSw+6WLBUw2X/2AVoVFsTH5TA8BUnaieEcVODVSeuOAVFu+IrUufO/BhGNRNwwpQ/GI+ghLBrFn
LV44PGcoq3K6N8BLkSsNPx7dImSk61lqRXC5XinQ5RmfW9CenJIaOVElmEdvSgyDfB+WmNr8AMav
wupQSE+2tXaCRHT1/+UsCbV06oAwha6YbFswbH6VtuSsCiWBz7qMBVWMtqflq9BpyAgAeGk5Se8B
WGkEab+h4KFWpSJpOIoNd+xr9Bsu7ZbRNIkCnFpGQge38slPINAGKcQ/hbkjj4enk0y+ZP4x8F9f
jp3FG4sQKyf4rOUST5ubYSYPmgKmukRumNkVo4w7GNUtsi7ZeW95MSp6OWQxlpewIbxEc1Hm0lBy
sdSLMSq/l/oLKEIVOiwj6Gl7LwNVeMvVBOv7dNB4hkldJzNAqbgdHSV1IKIJaP2ARSAfZTkZd7Y9
3kZHSGQRvypHKfzCPPtvp3TtBRn/3paHahFcAAMRITTDX8hqRmIWJpeEp5hCsDVDwmvh0qtzrc1Y
i+BpGLhRytdM+FEVUClmHKz9iBiKugPtgnkDfPfQKPa7vZJgB9CNkddUbXuAhwIsvUvBJhuwqN04
9aZZecUwlTWX/I5iL01YBYR1TiKHNbqDSTeziX2Y1JUBVfoRuYHnmF9ULvhpmSmxxhbekNYVRFLE
VspgXDRO8vOrAo3pLLRQf40blDKWekkp3UAtgoXHbmSx3oZ8JlsaY/4GVnqTEcV1MMdwQEFGWQiU
7lgiIDHivsJ+RAxp5FfbvJTAanEuqXPGEo43s8uhoXFiE5eGlNR2VIsi/YbRXKcFZU/ab3YYIaXm
mEY8NVDOqK1pGAHuvq+F/bDwX0r7jSDWX6lInsPEiL8SWrFWKWEf1psjZ4zUtpt6vMnKbNwvLU/p
DGk/lsiYzfvGh2YprX+qdwcgKk50nG13nUnFTV5uz/RlLKwdPga+E8scd/Ia0Vts2sPV1gto5sXf
2GVIMonRmsfPIhox1TYFZwXFAkH1H6eEZTlTQLVKRFrLFnLY2T/RygIpAcP4e5Hwa8mVsw4JYzqm
VCyF+PPGrNlxqdOqyJ7FeJY5YH6HNMFOZzSZm9JiqTBvCw76YEiBJlMzCGP50Xh6zzPR5Hf7UKyM
K6La8tF9u5xkerXCDIss7OCjPLrBD9y+qBG/OB8tGCPU1V7Y4FUeJ5FQLhaueKESWOIWS9Z3ai4F
og+Thb4SJmd0ZAKaTGpGyCAibs9OziS2FYssFBCMQrQArho72grabn3eFFbHBGdJVS+++9+5fEP2
k1UVXVtuwhtAPUr9vVW1PFcv9ZH0bYAK388r3AIBkpYjtyhSAY1kBlEhOHcAMRc1iqlnVi8PJzaJ
17kH+qIdI7vstb0kUaRo+AdaQ8Oi2csQ0G7kbbDMmD/BU4non6rBONHh0UTsN70wm35u1iqsSG8C
ADXrUly292FbIjKb1B/OEZ/Td4x7BriVyBBmpgMJ6mNglAt9hAvmGtMiic7Q9bmg1ANRxI5FT3JL
LZDiDzaDtDJEhsoBMErT4DamoY7kaSQp0tTIr/FwwIFdI9JxCARpWNDGE7voxGas8W/0IHRgRwo8
WMioP97eG1nEB60odqgTBA4MMq1d6Y0BlhFN8qBb5m+X87yscu0ETHIj7/UWuwyZZ0wqPZOrdAla
UAWL7l8upViWJeO8nOKNnlqbTdvIsgavhWeS6GHWndUMJDSmhqlEaY+ykMp3LFHtXjbCwydC4c2c
Z4pF7dR9E967CFswV3kn5kYa6PWibpz00PCOvwsnwo1kmXE38c8ze9YOrVe48gcufLMHc20WT7q7
DsBADWytj1z6aoTRe6LhRz/eCJYR1Sf2eQfbcx7SBBfnorLSScoPCTKWu5tZa7PxC/tzBO0osB74
9CnBBirL5vofDmoiFdob5NV9628OqPWLUvby3njIvCF6eqrmvgX3kJ/K5YHDI18Bl4Yqy8cxNHYe
me4EhL9HRwIuqAZUcx1ZJJCzdgVT0Vq6Kv2W3eOxN/GdAkNNvZ5BARR3QacF83iaYFEvWSNa9ezo
jAWjrkuTMTGY6mtRjxJJl5gjI8D1BHOl3fRkEqGOFBdIKgy49Aq+729sQSw3JtTJbDSGf/2aK5fH
QHGUwb8CF+Uiu/j16StSCtSe14VNDrTiKawHJRwSjLL5seBTXTix3oMRmbVVGTSGeIg1Y8m2puiI
RJUm8fLuXpLM/PMlFJjssqN4M8YkMdIgleOfTDU+ugI29/s8KtpvhorNWGy5S7oH96iCUIBgoGXa
lYJ8Fi6bexLouO4uz4jEmqdmWvqbvyltDAFAgC4VPu1jZiTQCXJRtZ8ciXfw6YcJ7PRL+7gcz7Js
inPL682RiLF7uK5M9X75vNcqbiSQoo/T5p6sUIeZF0/bij1RqnR2Q6uKtjtvOjz5sZf0eawj4FI1
xi6C0emVZBpop7dSwExJd2Ts00P83NrKp5Do5Q+4z9uswd0p8BJS+pVdAsPrbNXkhi6YZRbSuD2v
6Mbc1lnDZS4rUqD0kK95TrxBbs/hgkOkBp5f4vTTv+31Nu565KrETirV8EIuojY/oO8K3M70jXsn
p3IEDz93eXjDupJ2lPK1doqRGO3sljMQGTk/cmCbKdIzq3/WPV8hiGzCtl57MRDgUkLn98dFMHNz
+erLnT2s1KK1PxTPKGpEJcOIWafPNbnAztKKjg65fxcASXVUDxY/rWbng0MN1DMFwMdtuA5RiTPR
8XfqT6M94Kcx2s4GTC+ZvCgfx7fxt6MlN4B619h3rA8Hj4LwyW/Rsqw2AtHGTJphxgW2gKVWY1mk
3+8y2GCbqEh6EPLz3AAnBKn/tUY1SfLlUYZAtRiSWNBLXz+Fsx4QATErU31CXgcvFthGXTDrXhWf
1Uv5/LwLWA/6hHu5Bqykew7Rv8Aqg2a9i5O/aUWUNlT7VzIM08ue0/+rtDmOSo+MePD2Jsmbo2K9
YJ9/sOXtSXzYw4dkVW4m0zSC/PBDj4QUMQXIF4R+NQxjkSpYnLlj7c/Eaw5IyoRgklqBeOMMgo1x
45JCBOj3cu98ixjZXQnIWxqqk6lGLmNkDeT/9BclobXKX/e1DIThiw2IWAbydLIaKUBgYSyOc/Hd
ZWhcrniLFoS6b0OwPcqhBMTxtk7+IXcJicHBUYfPdIBQC17gWsclMz8nytqQrhuux2yFF5ORt9YG
GddDFxHBP4RuG7ul5I8TB47HhnSDTdndLfwE+6zc8khqAH9rYMQKWL6lW6oCvWTV2iXEt92QFlqx
ClgZdEEnSTSjMUnCSlx25G265CcKVxxer4ZyGzzDnKGYzY4bqv4ZZitQCbDlwU5TUrNn7Evs6H0l
ZwwR9eVsXnrzaHNp+lm0lC0T7gylOyeXcbIaVlpJkCw1eI2ZQjn28EI+Gt53oabR2U30JTGETt/+
BnrxkrYDpJNXfxp/QZI40dwmMKk/kXfTSK2S39mSezTy38chj3Zz+do4Eyt3+j52cctJiZEG2kDK
ewbHTrgXfSF5+9R2KgUr/ey+T2juCXtL0+XSSDfcaKLaP+bjoWHjIenFreATHF/0q2H/KQf4LZP3
7UNxeB8XEVKTFfyeO8fa6T68san/9tOwCIBjDPx2ZGqR8vPqXzv6AmgJbFdptQ4b6tF8OKVfLYKF
5GNsR3IoFlnsNTr2/8BwMf0MQo1KFobHIkKUTTqfDrA/kbbnRBZXF1y47YG6oCsLVlSd2MBzdeFt
oQn1+UmJ1RQEnwSfTUWJ26GxlvnIYRgPwoMpU8o7RnlIVjxsq7Z9VptPlv/IBcQkhHPiF3L3rDK+
4eZ7lwAxT4ye2N5yyg/iV5MzPJMkedyHFSj+QXjPD+4+2eUtQjbBnYRArltPyWNP9WzyzSKTTACb
DUn2lCWlkY9VWrBmu9VBiNgmK1zUaOTTiDlccWrastAij9YeupR8mhAXUj7VabvWxryd/XrzHHFC
gdumqEWlqwp+4T6pf861luBUSQep7mVCya5Km9LhOkY8D5rf+WZZJrysAK0MA6+jNglpKIj8URqX
IKOmPCqp1AAurAYnGrYCUfQv3+rDNTBRn2WG9LANbICOCMwAR7T8SmMevSK4v1EF1EXGVosSW7Nl
FCrsUcbOCXO4xEoSmJLNtS15qm5RqHK2P+NC5vTTtxKaFi+ognQVx8UmRjY/gAP4jHoxVP34k3H3
Fsn/MxYbT0ukb8I9YzmZ62go5HtC6H0O0H1rT0f1j0qKY8TWkSBP6kOSEA7zodFmGOvJk4ScZw6H
In5YrMyWPH8Cn1MBGs8zj10U/bTbU9s5vrM37ouFnVb/OsJXqHtZRv5HhTdFkHNVTdpOvtEEF+GH
Johum+ii5WMeGgrVZ4EeiVw5/TtuW65HYli/OEvj5ScTTvICRFV7kkmWs/YyGiganff78uxtDs2F
RCgi1kGJgh2r8PvLyrX1/fCfmb+XT2OL/0c9MciyKsYxRSt/vVPGfDse7DMmEMe1mTiNHPCCbjh/
vxfBb9YpIYXK2CQXhvuVXw//3aNiQoXBQrwCYAlw/nrpnzd4+/gdYn75P5P58+pzsjGArcX5htce
RY+YnbEtZXz3loYTOiu1gFlYeO+ZfvX6K1R/HEuu0Ij8qMVSQ4rpe/04dV/8OY+pPIjnYKQGTg8u
qmcbs+OaAM98DsmgeoB0FGptOzs5+xwSWk9o/G+dmEs0l4cKbJH+9XltGpikJ33b0sz8u2LSv4Cu
aWO6wYKtFj46k7Poiul0ixJtaX5adaZw2PYFh9VqY3A3a/uE4D2AzFtif82o13uJPSB9t2AQugFW
0QC3nD8MdWbijF5LkySA9LLLdtpLZqLv8tWK1v8Q8dspo5kF1bsYIrw+jMUnZEouij2SWsclLtPI
1Eb+F0artNCtRwt9kIi67N51WoNA4OfuY5iFpLKAylNbySklrF9LLhTJjnY/7aQI+1NYm3IFgx92
udezcmWLlM3qffA3+/ornAAVo1X9lcNcXChmvkIV8BC1Da6EtnmH+Ci1hYe/Q1a828mpVXSKlc/u
nB+9AGtFa/hUyie7hGJCjxN8VB3kXUtG4DBKm1OY1en2lAHPIQxqRQvfyI7L5SRCrpvYWohc3+ov
kGNRgqm7358Hs8TKmAqRFeujalfIej0sze1/Ja2pC17jNV+THlRBdMAahwdR7CHoJEyEQSav9Y95
sqIoqp+L91wfWzNxmLq2qYkkgPmXbvFe/riG2QhAdSoCN187MMsfToCvBrc69qggVgirz9Y4h1zO
WEcSLfPLA86QDhIMORWUSNQ4AxiQl6zENrvzGJICPUrjtxydRo3mCjnjgXPHO3zX8oL+Hi45Cbnh
kGq9ZQYYFUcaHnRVQmYlD7cz0ajzh9X/oWNSxS9rG4QWQ4/CAhhXf9HxKKe/PE59yUgEF98lI4P6
Z3OIWOLgNo1W5GCUvsuvkHTmBMzRisCR8ZAdbxPeQbL9O6e4xoRJ1Ze4YUtEb++AlqRwJGJEiq5c
qINmpA0PtCAedX1NVYZxsO1/d48GyNsuCPVyMetDoRFblxwaunRHT4N4rhiyral9d7JgapihZKEy
2UWJoh7jTisSfvQPDAgz1KRz7l4ORAUstF3XYcLpNGKlprT+OS9vT0c+11unbjW41WUPjgxeImho
ffMxJsZNYt2KK/uwNv7E/oIuAbAkmYJ1y84I2DnZ8Ip0zv7SSea0jyJ74NzIg45fVDXhnHzakp26
7kCXU8CekoxWJaIrpiKRl22rIA/Hy0Jgdnjjdz6yDxC6DGC+B1Iprk8P0Psv5cR7E5mVxOUNmeKW
6DK3aNJsPLkLpoEN/TIj4mbiSNfNRH3iGFVbkDEo0JHJ6CtD/mUlsMVan15ZHypb7HhVyU7MPYSw
EPWOUVPvv/e5Oy1jT3IRzoctLFZgBGD/3rkMz2pnT3eFPkE92M13qfak0/Pv966h4NFm412agCzl
jdSxz8LSeweJzwlMIz8rZFSQUWvLVVU9zgbgj4ogComzaqNP+mNE7nQNEZsT7EhmoFdXEe9+six0
K5dnzQRj6+GbijlZ5/ibsDD8XQKUqfVjoT1pvEuv+9yK2VcVISJr1MiSPbz3ZeYGmKR5jcALvibp
lIkIg9rdknl6nGnkadlF35p/dpgqt2DipJzB5ui4PpU6XBbsSjzdkZhNrDp4WsvVd8WjCRt/fw1W
4oNwLyKYZ8A4lih5JanR7S49D6CrvY6tHjgSIfJvyAb9Wfph2u7gUClvscjTBeyIKhhlOe4JGwPN
b8SE4BnxTeOyZEdfeKe8aucC2XAsWAZmFwelwJKmgI2EC3W6az/5a4uHDSh3xfWFU5iNqlS23UBL
O1c8cWvdwDLxVPfWCz6V6UNLEG90mPSwk67+xLPX4X/4R02DhU3A16wadwFMh9eqMVOcu3E2DlAa
naToNcLLK08g+aJwohF5jTENlO01T8UY5xwEGAHrvkYe1cOfUHMIaF/hFDTsCi1iXFgMzTpwJ1i3
ESQYDdVvP9KWBHNOhd2W6moGKqx6epTR79SYtkKT3DKfTwhyDLNx0BoMb08vm1P1emViGbLwcZDI
j+PbkWtd7BiUvc8FlVmoEQyDpcqXS+VFxLOanCHvUGbzJ+4lF0/pZYa+rVHbNcb7uSC7Xg6Qy7rS
KVyVdVNiUGbPwBdKPaR2rwCAGAlm0F43AXAXgmEGHqvdH9gHkCZ0JdFShRcgWP32fnVYx3UKMptR
qzhNoNIQa39gMTX4WNx494GSN9PxM2C/ar0B6I1+QYsEcP3dlgoKcXYv3ODILTbdTg4MBvKIR3CQ
GkBUPSKBedh9ZF/pUR3LAD4jD6hmi5LV13Z/ffQe4NsrbJkJ8iZyufxYXHwgIK+lGnzb4xAIjztH
8RLNKGa+dCoK+n5Biiao3VhFYonHZb4gZPZenTB5+n8qMEz9Jo0J1pnl1/HUW96siETpUvvVk2Nq
R0kRS6mqXT8u8i3F9ZmQVB7ehwLyX/cHlwDwn0+OgZ6TO5xCmo6G+pU2zmavN41EyKRtMdI4svr2
qm3xoq7fOri9uhRAJO1W1748CBJhx6kDFI1UZc8GGpNDLEumrHwxbWhZLCpagxUrv2n/2FuBW5Ec
cA0JXHm+KwYHolHxIJHKS/Epg9LMS8mi1hgvNpKW61fz+z77MASjz1PVrxOVm3QNzTsNU7/8dudW
8rLFHhGEg1hubPkxmxj6FYhQYVbhooKXGMVtTcjxhaHNVLAD5NZeXO5kV4JqBg44HGmtG1TgIXSf
Qly8pclowhFQ1KQiODvlKYIEmOWsjrEiX8Deca6ks9kRW1TH6d1fai1i0ZC2CHipnIHD8TP2NCCh
qc5dZz4th6aEazcrs8f/ugNLdjNPITvVWYj6NrLIzta8lNPAmv27/kZp2m7flMgYSWVqhUR9GSQN
A6OLjUAN5pImNCJo5iD/ta4Rbb1R8xkGGnhfKx3lARlQdZkUD8eBzHYmp5cLObzEUQ1NRsoOnCtG
sIiEF5s85Sbv7KdQzRpelz34h5dWTaUEIoLB49JbPT7kpqyCWNnABgwD2+wPrLi+B5kFe78z4aG8
L0cZ0Z5xwQ6wS4TZJFV+Gj25Gyaogjaom+JYQdW3vxtYyT0hc/FfM4k8toP47X/zqvyFoJHixfMI
gw0TNVlB4Uq4xbdUMXGvxFcr+p8ER+ClU8VIauW7D9UNPbrZlXKWJAdkem9pmFMpTvnZHbSl/9yC
lR3mvw60aAteRAuJo4a16TEnhwk7O5EDTY0EnNEkyfyyiOW706P1ZRt8zUFvQqoaA1s9SjBFDhnc
2CK64pAkYeF5LdOdYeR0aO6Jq87tPogVp4dz7W6pQVILapmu9YZWYAxCPKfLNTomG8PfmvT4c6ty
FNykDoUtUydd8tMRzBBa1R9SbfYlhL1oF5MPyv2i3KU+CaQbjdBxeiyprAQ2EMtlzZ8OTe3o/oK4
VitYn3oINqNnQpB5G+iEA8n6c2Mahzkzo4BTfOKxwIQQmSs05A2B6jkfes/My/hNjmjK0hdBJGqj
oW0G0NuS8iROcI8j9vge+5imIkSlBx2JmxpcHhDvWdZLBDJKJhsAV0HBjEs5wjOHZ9iDsxNZFoB/
yLFB4VuLeZh3VRb4FopTkQbfRJOPyBTh+kgIchw7qBzylC62U40dcqkW2JCjK4leYsTG0k5LKNqN
uetTwtQj0vW9vd/XGg1irvfWuTxB6eE/jM1Lq8Lo2TtJDZpqYXA2UZS39c3X8SCPf1Sn4JsrAtQX
5qo/E0wrBcVrvIaRiGTauLn0X8U6Jx0Nxkx2WzVw4/X9iSSmrD4XFNt5bkx5ZLDlvXmagKNqrHHr
3BDc3kwXNFmu9oZrFHlPRBI8+zOie1avIM5WKqV1pkM1PThT4w6UBVbaIP/g400fPQuBmDvQl/kz
hnstWaFcVCzaw+2FRLHnJsSitU9Cnrd8tdT0bB4wveFPTroROHpHxW6meoMQoiouaSJ7FoLtnMdK
ujZtS7zf5FGm7A6aOgW+AvPoWQs6NBz9w1k/pd3D1ihNmCDcqzDSy21Oi7QSyMU0tpO4CD31yPo0
AX6l9XB2nl61GR5dv0dGmlHcWhp+K8Qz7oap8Pdex+v6XFQiwJqjGBwdh3GL8wlVHAUiQUagQbqE
Rq9j+mGh3Vc9V6E6IDrgdXCJuIOC20Tw81q4Jfk3NuiF6ukdcIW0cYyc0rFBlGwP9AeEDrKCUxTB
Us8pnlqBabVwfjW4bDiZyq1XeM+yX/PerP9XPV91aVaHhxINiv1n5Duryvmux8YE65g5ALjadiXe
T8uVlDIr8yj2uuoBacxXmvq1sN8JZhvRzQDRvssPdJnUgrWremCa4c9mYP8eL8CwJcKIwtS49gKq
SqOWT7Eq7USiO7yG4cJ1Y3M0AmRa8Ps/1yliW6dyfeFin0o+35k7cIv3G+97mXfw78fUXrhKtoff
MykQBPvH6StPcaN8viVQD2Ji9XK+y4k3/c/sNt1XFrTR3BE2epwyNhOOgcM+5eNQ7PPvCaNjpMNz
/ezK5JVqge1bW4gAadMaebbN8H3mw+jEMY8HN8qwLRYDdxKMJa5raVAvCSHOYxgGkygpiGY/dTXf
fqs/9X9lKjhtryA84+42ZTA/PyzXy7hJNMEykeWUSyxo5aDNTVq1Ziyq0y1sDeTinhQpkz7nNQco
eSH0fiNxTwc4pquXCU+HGCihzL2+BTwkBLVzT2kFsI2CqpJxcKmLs+YcLxPY6KLeocnYz40JGGhV
VPiO7shDJvwurfLmqF6Wgjk+eKwIyCqzEW3g6ZEsX1fjaOmK/+ADN5iWe7dgDZBcULrJ6F9tTRvs
YjWSE/whRldb4yAK+5w0tEgc7rEA+8dBatvA8VTSCCMquRmCDYHHzTqc4vRmGQifr0oqqIYY5Wy8
vgkpTKsOraS7qvu7GRQkSAONV9ogTf09TyjV7Y7frrI9O+hdsj8ZoShp1eaSAkatGce1Ox3AQtsr
iPAjAN5TwArGWW445L43vYfSAoZqu6p7YyvklOc3YBinekpbggQT7TGcbKFJKGrkiJDgXpyumNM1
JphHa5etpmxwnC1I9qV1bZ66NiFXAhH714duZumFdomPZz7cDmGQaLhpQPsATVJB0cCkTmvuv15C
J8/rTW04CdOkPV5WGSlKnSRUBTsaFY5Uwxc8I2qWma1XhpAmqx/4hB4McGMnE38NARAFC1bKE+sS
iQgjc4DJuaAieQsF19FQ3+ZTALxL4dlbgWGpq3UqKgMtQ9ea3HHfGnF5PLM7OWFLALQpV4SgFspT
kMfzDaZ9ZlTdq11GRqeauV2u/lpI/gUOYwvNxakxyo62pWyVjZOuHZCT46UA/wDfC8ZPz2MrSx6+
Jp2uWFwn9BXYNzU3Bj2hhjNSYNM70cE5zGpgCmQmpJy+gBbjzK9vejne6Fqwix71K8n/BGDti5A7
on5w+YDZoZ7XhqxnQmTl6vwbGY47Yexawt9fNQtFy030sbQwwwm6F/NYYvax7H7JynHDSPfxTy+R
k826p8MAd9osbCoGV4YVYjlSN+up6KZGSS4yR62qjNVk1dKTY/iKm/xDa/e6jOM76e6SVLOsEDxS
fey63SxMn2+Qk/njZIkBkR7VNHwNVuKhqMuXKl5BlzLbfw5Znoo2iI8i7FWwg3RzsrpWDcapnIkB
Fo3/Vuc1r7MCahTxDNMb/ZArnAebOM0Cac4P5knTKLpOOgZfDh3omOsM92SChGaeYu6X1ZWdfS7m
TMr/ZTnRfLjWYW+chARZFWLnXw4ZnJZ+LmuE+aBEIjG3xg/CJA7LR41mzlhaLLyHflVLwGcn+3PY
aPxYNuK0P2Kv5TUrnJWgzwColyM5iPliKshtVwI07/dc8lTKoKLAiq+9PbiH9GjuIGQhoCHNPf2h
w9FI331IPMrxBH+XoNmPF9ikL929Z2K+vL4eY/THkdXbaxSqXNqBlvZRrAA4OifR8aD/2dqN2Fuk
LznKXmWXuvhNyrCXg7uUJuSO+3RESfrvS95SQEaoGGYNAbLpHOFecSu/Jw6w0WBqxuCI44cNHTq4
p6qwtitWsw73tIl31o58xGbJNyniAf3atZBI9RV0uvQhlcGr9+1x5Qa49cNHmVAcoTCP0jScmvFN
NpwSdihqsx0nzLyU/4KSnhIx9C0VtfjMi2TUU2T9aET9GvyUjIcx/ueF3+BEFYVamWGng0FzbXM4
3vffZj0qUby/cIf63S42yBjfPCSaelS/Dp9/NJbvB+FKBQWfBEC3oxTXuNpIViPhosuTQRMlKImw
gnrjDqn+rCcDkWQ8Pxjpqly/cGOSbi+/d/UnhVx5hjjUZztj5JLFBnihO7SzxCzHFAMjmXOH97r4
f8TORw+o0yfVYusMQzzh8zviVYDqLazQtA8hyEx2BI3AwETvwDRM4aX5l/RyGZjOp9DI9l5S54Zw
cExxxVNd/NsUotXfH6MYUDJxxWXyeESNJgluWv9q41VKKe7MQaCmmaTt8WzTERbQaZl/1kT1l+7X
Jx8qTQ0c9n68PGr68DB9BtDhpzZNSi/7bh5jhoMSB3SeO0wqH0k2KKi53HybgvGNsL4H04HkBTJ7
dVvvIx2qKlgOhayFNYowko+58bfWItMyk+/nqvtFCEFF8UeOX7eJzw+5j8cZnlZ6lUosmXzBbMJv
zh9WMjKAFPuLfZqoxdZhpg527EYKfiUgXN7MBlOpR9bk/cs44UWzDNVNkf7JeC4Uo0NJGl5Pn3kI
Pu/jxH1ovHqfE7LRwC4HMPbSJAlDnullQu+tEURRZKx8xLyH3zfs2j4rj1H6mYFQ12r6JqHlMMRf
jn1Bpigww0NauEqQPypVRDiv/xYbhO8lKTgsVpF+IJAjNBPjSQYz3JGPD+EbOgVszIuwGhzu9q3D
NqKJk1DUtvOK183umidFif9Kx3AQ83qU+CVWT7jUfN/TaNqpPW6uu3NE2B0rAYtqMuAX6hSP2Q4c
vxHmJLLmoMkAGBFM0t5GiYsAUlFHpojS4OhHhzULVDWg27E+8gnZGCc0xqNFFmQ8rZfAnWeyfVfH
URbjGgfE0AKUc5pNaAxr6ufa9q3ONgT7EVGkI1PuVzOE56QLXYPVPyBEBu5fJzGw1x8dWGf+LNyR
W6ZFjroBPWHtQdkOmugPhQFIMMEZ2RWAmsdVMVYfWyDVNrGlL/CHKX4+dJuJsSWCCLq+CUVVcQ+A
uXyuywV6m83/pQpfveQhMIot8euvPBKnOklRPSPH+oGZU+J2Z0DabVBFaSVxNetIZFzN0Q9E4Lwm
Fn/QfDj62lyH/sUBnYyPqyZlWtTs4o4Go8bAiQ1X4q8XWG3yOrby4aSxLiVWU2iVfi415zoSpL63
uXkCE9OHqSAuC3aMtx+EznZqnXoTJ6xSXvYGUpKJdfEC6ciY6AceSqFPgQPAT4yNQeYq4TA2H8Cj
0Rm5Uq+WHjpCWyrvb0tVluxVLu/iz9U3yZiWP/C7cn4YdbIUW+BQPAfSL3DIj59EpsME2ZWoikA8
wLs0XEfRLfvsPQ5w7ktngx3uAUPTRx/k7zJqqmJ/dOvMscGuCIDe8Nk+tp0TsFMRKVHeDumVjoXk
udEPjcQNNFApnPmBQuoowjNAnrcvwKzM3WkX9wlqvESZ7o1Mq1T5cxJip1OT64ny/yLCEpmsSvCG
psHew4qOCtLUYfWWB0z6YFtJjuLPjpl7uusbhzhtdyGKo05mAB6p27RDacfSmO/qL/ztNN8jVjoK
fOwrBGEpQQFmJyWi7KNkXoGle4IeXPj8ThcKA3YBNo6533ArwJFQnh9wvS2JqZ34T2y3fQm7Nzl/
DTqv3KEdwWxfEHuWnc2X9eJ0hEHZ5vv4TlKTJlRjMXiX0L7XP99vRMOJo7thKokVtl2F4YwwQe+B
KOK0AHrZoIATfI6rH7F5k5L6Zh5/tMtSSOZ1F3IQ1k0CWyrzC2P1dtGzhhf7QunT7epkkXnjZvm6
0BTU1nEaKhVqxtOC8E6+NdXRKCYlQA61Oe0EzTRdgDM2itlrMRuWoK0x+e8yUM0PqXb2BS2+H8m0
NvisjTAGqYsOQ3BJKcZ1+c7LXubkDfAhfvCO1RojV6Cugm2ztRJrro7aJ18HMGvHfp6ppAWU9iaZ
V/ZBg5/fPBPv109cEehcJ9THtrFl670/VlHQOhnvsMVdATm91wLsv1FQxriBjKCxaI6wS/eM1BBI
aUj2pi3koNOGvfbL4O4Cc1SlROsRFqtHalNcws1nTWb46yplVlu4p7AF5s35FuCkQeLfw4dYcBIl
Bz6NUrAIsCFt27jLWzXTw1RC7HugrHNw3kQTBRhDZMtAZxezmZ41frLY3pNyKC0kbPLNOBTmhA01
0aLY08oUn6VwUG0LPQnLj90F8HZgKKiGZBYGX0JBPyHS1vgAG85nMkZCVe0TOh492CUL9q6jEM9Z
qFYRhgWuF+shuBPDOhzp+JNVRG3tRnFJByp6QzXFXzrQQ9eiYIMBLrXQypW2P0OMIKNWaK94gsxB
dlhRevXMJ2//Z/UBeEycaHqX32dZY9wCVxo6esbM+8SW8hInJk8MyRElCsNfyJrUs8W+ftX2Lb4l
y8FuAT4AOWCE52XNP8OfcjsB8NsdzLstz4yIul0xn+6p7SpKVcGuqGObOXSRIpyuKBil39sEXO9r
BnGW7NIPoPyZHaN/NsjFRED9UDzKdDSkDZIXjMnN0ImfUGquw09bmp1eMFrBfcudbBLiLx/z+O/Z
kkgi3taUH5hAXgXDNDYLvfaDE0czxt6fzdwJFVRQjcG/XUsS+tcnev7LhD/9HG2kDeCpqvkBYafm
f3bq6DO4KkGGBgYAUffmRSC1gfBpg0Oo63RBK4KXqeUvoO15IE62ATh5xfbDUzrFztbasyTZIaHR
yGu9YeiAwXY2yaTT4d/1fS9i74Y+nUnguPszOOJz8/jlma2KCrZy0VkeGnrxKIH3+hsXCTqcpHR9
mg20Ay/MVPHNOXhY5mZGGIaLND98/1cvs3y2mvou6LTo98OD9dKo8ugqKPIApObyfISsG00BSbHQ
drH5OUaQcIp1xgdwfMy0qtW5khR+de6ZvjzJ8umU9hFh97vepSqisH9mqr3dCvrTWZeYXlsEWX6V
mzd26rYNRl0j++zCg4t53EkPWEONX0ovhHOrG9VLIUVeP1JoF2BWIo/cANgImJAdilb85kDJJZtT
XoJMTsWtEqYgpPU3VbYK18f1Bm+FHAdWNsnD6VOt4ZszXI63XHHBODLatTEp4KjG7f9S6Gn02UFE
EvRlwPkbNvzspC5G6OLTXuwlJhDf+45sBEuSPV8sck7mrWVDO65vgdT0i8Y3po7l5CyaTxVRoiIz
IK7OH4N4n8g4d4pKBNZTem1CgdXMhqsDo8FMTr+xvWzAHxT4NXayFHf3/DNGSondd3mxNQdp6Kve
qZj6TBnZTmPpJNO7pmpQzhc3vjLJG9+97D9oQwaQIIbjv2LGpnaPAt1JqMaKAAsPd0oG+e8Jce0Z
WeqA778E4nB9RzYKmAnzFsJZQu8NitOCL5kXjppHwXfKVcOAK3FXB/8TqhHa2VkhZu214YBw5V4m
vu7om5ngm0TYndSVs269rYO9u83BeuNLIa4+MTuIp45g0u4MVxEOf0C3xrbLpQmWXNK3EojKmXcu
esjKCYrFOaTveo1RnK+ojCxkm9I1LRhYdm6+jofXDk3lQJeCI54wQLKfi7/EFPH6Oi1vkOHqBffe
Zmt+FiGjHMozzUUCiMbb1UDvUZ4g2NRvqUwNPrlFab7wep0Y3qKREr/eSu/EjSW7Kvu1vHTk9dTx
jxVCchoWvFqh+L4UJcATuvaowAPW+I46+sRxq8xdktyOi85pTfXg6wbtjm2Wy1z5olABjfVsodqa
RJHIwWr6hPotP+BUYmmw8gyroy8A/w6Y00yrEvSwFi689TrpOZdBvrROZbfde/TgSnjq8/tAS6BO
IbFUJg==
`pragma protect end_protected
