// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:39:12 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
nckDrfzL0DDIaqeITiQU83wfgqZa04k2b1MvP4mAH+fL7WM1sUx2HlINHw9LvKB+
WWPDp1+K23h/HnE6Qjg/rfQl77fhP6Q9H+IhsFrZrt/P+vX1gRHwbJaYlmqpG15d
GA77Sr6UumqOANUGw0bgDpsJWHrTVaduvqeaXTfsFKA=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 3056)
5Zl23mzKnLRh6TZ8QwBhEtDlbV5LIDLFutyr1L8tQc+cBrzK6mWRl8PDSriNdLDT
ER3JZC+Qo44EwYoiwxFMNTx/F3aYb0CBKz4PWwqYVrh5gdhd79YX7Wu2ayhMB+hC
kIolLKYPwEvV2PrQnFvEljHX8tLBCOkAyVjvpUkogiDVKUdbK1CgK9DTb3Eb1vnU
Zxe/ReH86deZjsxiCAUGZf83u7MCl4YmjFZEs1ILODdfJWHTPkrICZGYTx03Gy6R
GZfLugQfxdp1Cis0RpBwfKIt6edILAbompJeQWEXBVOOkDGy9UgtDOWP3JDlyJiY
xODZvuQ0pq0bzO3tv0a2nrYNrfdUfcxs6inzNqbq2o9VFhNGDtcx+a7830XKjy5u
czkmSPAutzlWvbUCfDxjK+uJYEKEfewvKYf74Ep7w7CU8ayK8k+YcwIUfr1lKJWj
zndkfgjtOh3VmZqViim05aNoo76Zj3fjwFJphCwhWOkIdOKjbvSbxebVN+pK24xm
Zz8wzskipZg3Fr5PiODkuDLI2vRYzFxNYbCjTC7+lYB/AzmQf8oSYBUMmrVKwmWj
lNvH7T3dRjx4Srqz4P40WBLNe85uSI0N8o8ZqnncMrq2/UXHVIWJduYn+uuBtrzK
FAxi0DIk3khizM6Arvu90ouL+TMS7iujQFyTBuO4/kZ6udclYTu5kCO+MUbqCLq1
VxpBHpEs8h42hNvjOwUwapAtqlI+p/3SVRKfLE28WcFWBMfr3ARN4LhDLrNqsHNB
dyRAle+e06piQ2nZfSzm+wAC+u4aMsOb30NclWYxRYIHpyXJ1+lce6L8/p/NDFxu
vXy6l1r/1nfKXxSJNvNu0Zsp/KM5dNPbUbswLEVTiZSTjQ3jk4NritxrB7Na93pO
q9tXVttk6JdzLz6+asCYyor47kA0pe0d4f2z0l+zVbXZIn/nI32qlt2psa7DsTbw
90vBEmIiXIUWU2MbdTt9ROOG/TW0oPlKZc6Im+7ChTkCaC+M3gJ4xtODly1YMcza
eVQPwIkW3NNVQPcM05g0KN6Cr6tfDjHPNVo2D1XyOuQ+ZxUxEleGy8HG4zkHDy4o
xra6QIOXoDg7T5RgQrf0P6rVvJ4GGgmwkKDq3EcEQHmjeVvEczdp1d7+nTRWIAtR
UJd+f7pPo55ZNaJ0drMyIA672Otf8zmgTaxpLFId0n3001Ch4jxNOrnJz9Z7PcVU
3XgYJJ804iKYosbzJIwOxPKND5xAayOOs1xayKs/t7mr09o0h9Ac7xkRQYBP1gz/
cw50KN9yAfxoZDkpscpGnmXRhCOpwxq9JVkAByjVhWPHjMgwol84A6CAYwtBwu/5
At1Kfu8TN/zuNWdV0pC/EBgjhhNY9a6Y4MsEYjVJJFuX1VDdS5NlSQOgdy4YKz8N
ru5aNa33FNHAFeMv/7qJccEyVW3wYyXDKe109bH9/6zHT8rCAGhzB7WtlpwuzXkK
K8hDVF+PMl8p02Wj33CvvDlNZCfaPCK7NhAXAGozGKWOCAF8q+6IyTqS+PacLT9A
PTnmSPNQ8ByvjTlfRBV4BuDhio+OGskTeLhovUgsWqazbffFAYozUxjUwn7LtNZf
VCxsrPncHqas6IDI9yXpDFZMmQ57/lVaJY7n9CqlxFesZiGEDs5xgeXR+h4UWiDp
whThwBPGE4zUBXYpNF9vvzoG4dtIo9RQE5opqOCMcdl/avmrMagqjjiPVp+ub7Go
4eSWS60ZE3qZp/YUiFD/kCzLHdtGf04iiwBdAgGXwJR5DUTQyL1DfAhRgXfrHhF/
2dOB1HVO6N6UBRttnJrgNKFYuunht9RN/19exuo7BL17eCGP4oncx0eFQ86VB0AC
GxhF9WWn6WoWg5xovRYUqZKjSXrEHSIBMaChQQDH3bex+WDYiUkqFriqVQt8q3X3
vyVFZmZ+/hLR8GeQLbMcPPIy2CUEJkWkcdO1Xcmd6ZZrQjF7VfUOsWXkBqHhpiaP
fpDr8U52djVoCI89wJTY7YxI/En/h5OLcr55Rxk5XXOW02lXKqeGKGioiGi41k6j
ZYOPjebG5ZpzfJCMo+sHcqUijvEY6kCC17kiZULlj/JzPxKPrqt0rWKe7pSN5f2q
EVds4FqhHmR7hqLjj6aLD9DdY6ruxdCJhC+Sq3foYGdqf+QobMByBGJvIE27SF+f
hBjljP8yYaJef3I11WPKWVz9jOXoGD4ky8KvuKQe8Sme5HyF2t5DV+PmWBm05W0M
Coo6d1H94WTmZ5Fs6/VAVf0MAvnqejYpiXZHL84p1D7mUNmWFS+kV0yO1fJP6ct0
sPuULHWe+GLzvn43fwWkB8tTQL+s1ojOoRCZP8ry0wie/lblY0ZOSs0TF7ITXCaw
8YTRX4bAIMfShtfn5yJPpMYPfq7pcbG6upzQhGR/sXfJ8lWAMTs0t8vLokqci4o5
ctxvzU5wpSPgpvlf+QDuhJtv7Uq0RVBIGNDo/MchK8pHISzvusmHRBuOVjCxowkC
epdAW0BwZO/HC8bC03lFMrZaU//MEAQFzggLi3kCtYElgGxIVLmSJkbXKBl1K9ZC
QQ/hgZ82TSnF+zs1ZUbHu0YW6GH9idxvWxwxA0BbUOLwnrvxumxkBIxnBhNKnGG4
+VlJochn7Nip8amu4SX0LZHjs8O4R5nmogI3ezLm5hrWK9kwxITqozjAPvFK08yn
EGw85S3zIU4LdnMZ5FzbQTvkB6XBmaCmkwoJwDw24RaEfwbNPBb3ryi/lZ8D43g8
7O76UU/lDqehrB2+U+pyfoB0jngGVl9jYyMziB+bBYwEjw65DVHkroVyjZNskUSF
ZNYMIJeTNzrIXt3mWvZamoLaslsINYicLHIDe+d+QxmPbF9juvlxbvZ8UiegqkUf
2uF/Lg0EHI7MegazHPy3XHlFWRfIInZy2t34N+mXCMBi33CngtCU3+FIW2fVlGwW
ghrJHMgemQYMpjPZnOFct12v/TzE9XegkMsknu93V2HXLWKkCIESHDAVh7EIOasO
cdIaaOYeY+2AI8bIXYAsX4W8ZBhcG8kQibMHjEtd4aIobqO8Oz/zH+r+cY31rc5N
23Etk+NoxC3HrfIvq1f7lG8LmRM9ACmRoO+dcVxgZTWeV9MSrWPoxWMizZ/6le5w
KjFHmfYI9tGUbn1l4cxR8PRQc3wwUfGGNNstTacttMkDvAucDfy0BFNvAq0LX7WI
w1PcWyRPbt3PA0EmKgnIi9iUyAOoDD2WMQb8gfezN1azaALEFc7bnxWP5mGKtTnB
5dUBrbg50fF3/m9Qi/Q8vPgdHKt2i9hPcO8SoANj9J7ROJCF3aqbSz0OJEtYhXm+
wd+C2Syb2MjxCUp3In5iPTBs+zcLOnEjrHhSPQ2hNm6m1XBXvsYE98L6twd/GoMP
fTLphjqbpsqKKD0xSwcPYRSYZ0klJY7E7Q2pjj7oPWPx0KFptMlM0FQXqXdM7aiJ
prCRTKKroAIb9Y3qO7EmokvtzlbDc/koSh6jx8a1kLpZrnDPR0OsGL7lFn3YfVGS
IdFA6TdfWLSqf5DRw5rUeAM02fVucJJhmmirSao98ha1hmb20I6guwpU41p5s8R6
8GIiRP0UDsQKIwFFAMRmY/njBXaiZFTNOkuXpa/NRfvWZwTaZfBEkbw+1J4CNdcQ
djkNlqoUOCcYtiUDMpyGgf6V8HMIT7u9+DjKnAHmJT+hjZd7wS0VuXEHLRg0S93A
6SqC5CWoAVrEY/OFsIcaQ1C7l6fBb1nfL9vgudTxoUx47vvqQxsuuPWQLetRmDEf
k3smI/MZNpV/P5fzbUxa5GHwC2cbE1HtowkGYCOU8hjQZnIdevn/7DVRoYsHhCG5
2YCbBzs/ZVZD8kX4RdmwmCvDa/a0/37KDDC6e6YeX8R8d3iPtKmXPkC5nzcsuctg
STSLlOTT6CEwt6fJnjkoMwUgRwL/SoB3OcpRUyuNh6Rw/n8XLpVu/KP5/cACcIbm
RdLL3U7WJYmoq3CCv1Ru2Bchj93qSyhLfCSylDlAqrbnNT/ESshIsK7BZgSG+sXO
ItB0Qj2mbLdvrgmaiQeXfx7p4oPXW2TlhszgAocUS7o=
`pragma protect end_protected
