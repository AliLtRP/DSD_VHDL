// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:35:41 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
DSFUOAeVnsLrGwthkaJq75IHaaJmtnmxeJzOffPx9AcHWkZnOt99nQqlclIKtDmj
lcR2r7i9LIZz+h3qTQvOZ1NOr7tov8YL30n4W0AkFga7+RwmqkUqjayntGtq5ho2
alQ0HN+vsrqRrW3hbbmqhinBgS44nr7iLkBQkkW/dew=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 8512)
o/j0TNjaii4egEK87qIBwrQ6N3bhQt9Lde89Ch5q3K9wiuPCFnlEFXHdUiCfOE4u
E5DGAlb9xGGQfjO8IUP1tR8vXD0ynlZE8z0mTOOyhGZEeK3Ml4WWEIccoVtUPMlL
kKBseaOY97t1/YqjvgKqCjF/ZiDpjWXOMwjKZjMYtAQpINzCVogzIabFPWsCVyYQ
X4MWoCeOWDZlEQOYWLw0SsGJDqW/pq/DvM9C9Qh/IZ4tz35env3Z62wufkjUiL0J
lOU29hV2WFE+SkZnK295CTnYg+NtoIaUwG1IGsmUQw5efEajG8V2APfscphZ/Hcd
4g3r4n703W2sXjypLIRVsSIuSRGfk3tqJcv2BXd/dm3MAWpIuaZTAYg1RTxd+c0l
pOMiXYgvzCS5LErZJ03imlzHY4xwvddnZjg0YWqI+KFEkTD4ShYT3qKb9mQcOBqG
VMCaZq/bh71nJS7T+bFK0CfU9HUBUwyJmazg7kFdddJdsJ3ECNMs1fywztshVmjE
9g4IS9Wt3HBsGsVRYj9lfToYTwJ1zmufbDl9XwlnDEz4KrqJjR4yRYivGUEn1z8I
StghhIMIs+psLw8UukMHC6QtmzNe5bZAcSdqRC6KsYVVCOcrQLNOACvFAwNi48f1
x/V9L5xk/OzaXaLpn/AFm79wCA9RzhoqLaiYli+UwUFZzHihdFFxZmoInOpqqLpk
nvvQ94nzbPR5IXYmQs5O9AejizKlkARFJP3vf7ie38Cq0s9psYOKNbQPsytLh71z
y+dMgiG/KJ5Cb2t5ZiFQehoZDDaXdCYykmw6vro0eNShVaDzbqpyhQr/dH0pvT8f
eXmFG3LPmd8SIGZKqXhmhMklRsv4kUILHhwOUC7WV/u8tSj35TAQAEVxx9nnEhZb
quHIXvc2gZC9o6il9thd6jjpteNK4oabc1ZCgsJ6fEDUrLYtNRG6vyQzqQYC6mnX
xQ7D5yNG8oJ3ETfkYd71CkpL/QsT13g5zRWyop4g5sF/HQzUWSrISh9BuP9Mg+ad
jJZW//ZXSGsHcWcxFNfCmrpkMjel8x6Cf+LUtP+U7CpxPqKt6Uu8TVFOcWjIG0kq
elgMEoBkltZSGHeZD1qpexB8MXw2VpzFsz5YCR+4j3YzTaW+AYG8pEIum2aBvHNG
RY3dgHPcnr+xsR/KchFuTEBGqU1yaDS31N0k8s5slnGveJg2tqvwMYTGo8zzRHe4
4xAK7T63Vv6NzyDvdtq5UJsJ99Knxf8Rgzzc1g9rRQCbXJ89XN4A+LS0qS1czQeT
dbQbaZKnFLNVS0T0x/hst63P4soj3HDAhlzd2coQBBEW2+SVKrVsOlHRCenl8iTZ
757+wgomk6WHNwBTVghFOG/VEG23ZE8KOVyu3o1IlNjzK8J4fX1KML9YBkBbfaiL
1WKSyqtuXpnwG6VbS8uoFue3o7iem/tOaOHF8X5Jk30URlcsGOdzfXLzX8F5a7xX
lWQ4LVeuD1MNfOWQgcsPxQ6iFuLVsuHyWLKBjjHXGBhoSM6fUHsZhLQ0+ez1ed/j
x1MnXRjNxL8bbTJfV5erzMUDxJmVOtVT90seIWNwua2C0PGD4QNLeW3p10km5rN7
vp7V+PFqttp1utSH5Uj9A6jdsNC9IbVIgVExfA62OxagxLG13S6+JcAmQwsijOff
iGRhLKiuiVzfExVSk3as/+49vQJh8c68HQ5H/u+o2fw1chDKZf5MBDdOTBXYj44V
/E8xYxeFnoFAIhO2XGQDZxagcMC64QC6mTyAiDobbJKrgzNuWOSlo3lkm97FNytI
JprSMoeC+tGveNRQsbEqQ0j7P26zIunKZWiZDRCnBO1lzztVA04wbYMVgOrrFxHV
wmRKxSRB3uhMVciVkxebXqxDabwENeBmOn33nPMoG/MyqNpddFTWLewQGqWEqCwh
20k/ODEfe02qB53HXvexKT1pPT+4CSY4/EuuCFnJ2F4yfLiSq7vYcMcbC/9VZdvE
ajoqkq82C+27uYSe86Nm0ho5MupZgBZt8coFIsYLdxLEPMgupVpgG+VIsKPw5IPm
U85kcOBzJSX5lO3PuEQxh9BYN+WSFOBlP/giegnBgX5rvUZjW8gXA7dd5RqdFoPC
SJLlaDNayagm78YTUEmTOEcGkjRbtUy0QuZovQOQvigv/6GPbnA3yV2Bwumrlxve
NLS6UtPAHOVb1s7osh0AjZ4mmr8tZTYEYOdA/tabtUASYCTN2aoQgyB1y6bWy+c3
tAH2tE4Mhtc0sCTXmwSld/m2CExS7byJZXGHBXpMcP8erGlgnY+3J17fqRzJmKXA
efXhxMLRCvoT28hE3c1mY3qkelE24l90G56AmoAd+aGYHCjgB/aCjv4SjzeOTNQD
+CsEhBI5k2cRfZxouL9Mn1F8I0stC68sqDTDjjdjSFZQYf6FBLQAht+qawq9gnkT
UsnmjSpjyzkmLVKM2tbqS5O2jPRpNh3O8kRzfvKETjRkj0aCSrGZToS9RKLtlmH3
p4qQrnaDJ/RTf+2ZzEaeMLlwoWvqBMSxGVWPtYkFUgTwGP0fzE5UCtuwluOCOPJ4
I8XcXZAE5UpLnXSgGSVrUkzKO4j4ZKfcit1es9FWzQhlZ40XCpijLMz/vRa2MfPS
rorL/BBKDJTOY4+p69D8M/XS9c/j8ycUV2BIUgQYBdPW0eWxQk0dDxGr2RNA8eKb
GqtVln416WQLY9g3cNS5iu85agvjee+xy/Z3fXikxP4dXBK9WQyaeL2SaxWh4olx
y/Hg0wl3TLmb6BVZia0kM4sfPs1nAWIOJ+Q7UF+ePMg+AMtfJ9jEL6hPBRDiVxin
RIny3hjAwqMzHNkaqfww8b9MKCoLuFvxD0/G4pVRFvdGUY2AA8eMh2iTlFuvDS5t
fIcRzEJ+okXXV34lkOrmmNP8wJNLG9GmkZAulWM5bgkxDq4gl2fKh/7CXdOwH5gL
D6jAVm7KvOgUh9kaLafxOaYlQN2dMXKCdWHa7+HNU2TvmLLmzteKF2FltAkTEIeE
dY8T8W9MGOXZrcJwFpTWAtZyAeQttWnu+BZpY6bqzFjZmunIipV/PsxVbBC6eMvX
Y3EC6ugHr9928iMH/FdwbaGuhfDV6f1+RQrGrXYu+a16eRJBAycw5il+pAL1BjB4
4ObJbG4llY3ksmHSkVsB5RzAgKn9Zhy0e1wPnYkj5Gh3nRRJQbtocvNhIp/+J8de
p/XKEl5qnD2xlXySWj6cR0Sj36avxVL8BOLULC+1/CggbK0C16P7RA++KvY6f0oC
UcEFOS2fPRHTkkowujUc37DOB6kuxvbQBtT+WV+zVlB30P/hX0MMxEFE/TyhNUeg
LKrtWbeUgcPGtfRKfHW510GIjXwcrZaQRweVcsABldtU2eVe4x0aOehBBX9Fh9yK
G9FXmffYBhxeo0DASJ84O6EzZ8qB48Tkdm9d2Ld44lb/bgnoyDc3eP5hoMzQnK5O
8GqEQeCS/nd+b3HFbbcFv6lcSCD0Ij7lyz57vHOP618poOOyXet8WVTXfBe2x2N3
6wlkO2zORND+HG7kAEWaQeInvXS9SWLOwinWQoS2DtZYN04QIZkgX8H3nscjExPJ
HEY2yM1LdsTY566mPhuVOTAed4IzYCEu50XrWmkBD5CTRrn2oGe0j4J8f3OjSMf4
6i7T48CX5BGbRMV5P8VKAcFiZmkCFVQlYfpNgX0SH0uvDrKgt06Sae4sXfP6+Mfx
XysuVPrZaTtD2ImpycQFoS4aEwld3TivMoU0x97IN7NXkXlhylD5PrdN5ZHalXrN
LfI8s+4ftpsxh9UJMWJH9HFHU+2oGg+zJQ2Fra1q+LKfhwzwS4Fu72+mJV4yN8iC
DDlmpTfDk6Rvm97K//5gVGKY+wHNq4GtwVvelaM8u3J7W6m1UoIKjlHEz8In/U65
Am0BZGvSKHy8F6+IiuFWSJ5TCGcpQxY67DPSwawekxtYAq3uSbZxMa+t3+up8w+U
gJn+h2YZpcffa/oIp1B3BRN9onJVvSxa2nqdw9tPcKeI03SjSEJ6frdS63XjaLur
/uTnTlAPtjj2CL+hD7zllkXqssFPy22UhT51WVmyvvBmIyNpdVsL+xRvvKF2z2kH
A1j7B2r646n/53Z42arOo+j2BCgYpnDA29pi79PP+dfP5ZdHR1RtjPu/shylARSy
rlpx91KVJdU+j1UKGhonjH1w08Sa6Lj+qBPKUMcVAJjSDWsz0f/kgJnMeoBTj2Zk
NFcvzsvHOkZFBRFgey0DpKpIdix7ouI0ZtSkbgF7NuKmAtF+lv9C45pD+TrjSJk3
pLUw4Rl2UZtGwqsb6g+QOvy0JyyB4SjA+cKVNIXmilgX5B3i7X5dPpn753rXs2Pw
H99og98CCLnAXksbvCyZP609n7HJjrVdw1NI6P6U+IjagjUmMwcrMprRIq0xXuNx
d7Eu4lHjcOUK/XgWLUC7yVlP7SIfMjkTBhhHlm3YpRkF7P1Vi8lslhtgiPF4dPK1
x/hkhUPO/xXECkmZRdtoJwCKIfNhVAV8JzPqnGM59RSNlIpkWAuWWQxHHp/J1jTN
FTg3PCclivM/qKFTDKtduu6qAtsa40rO7EFOgG4v7BIuEtvXZ+PwN4j4N5ULWUq7
pcNQWzWF5PR7Q5+W7bqzhSRvuQPv9GBKipX5s3W6Yu+OlCyoJQA+u7il+QC+Pq+W
a6ZyxqpPoQX5I6kaOTor3FPCavsjFkFYcFcndxl18c7o8gu+0X62wCjiXT9MxfDn
dSbPTpHMQ/bpbHAtBn4iwq5NSkd3ce+kQ/fLqj7e07TM+TzcIMYuAIbQdNLV6Pui
xw66xFHehALdyhWingo2BbEvHaJ7gGHYEiCB9I05GT6U6ILM6CyUSVznEXOFkljO
5SzxGjEQ7WhT+xSmNPINUCD16cJv2nM90UhUGV9rFh9MlZ/ja3jff1QTd5qkLHo7
y9vuVlJhLdSKp93CqT/Bf2S7sTrpp20yFw/7LPdO3XLUg5egcad5txqmzfUKrs+k
S2kgDASiKH7akcwW2gtdvySNWDTABdAA6MoUvJkPE1Ho4sZcq233rdcOkfUiPtWl
qKcwfXb4zBJP6nqiaUtEnHCOlByuLdXHoWDbPTsCohRD7Xr0S5K0mBaeXE0gqmJP
/IGlj1iDvXV3wTg3NlgazV+p1ehRq09BrhzoicWGDdW4M24Id7Ubt85rTLJrwlay
Hb8/tHYjWU6zQHHpLHdx/lJU+vOqhJP6RxRZL1CUQhF5FL+CDbUsLARyP+GtTkFo
o6Zmfq1AxiuaKFqavE+lWVEphNEvYdeIOAiL7xWwQQgpRc6f7ssYehkgcUcbLdEt
LrK/Y6kxCe0DtI7KjQVaoQsizGPdtXS7Q8pJd0gXO5aqicvauEF/TdVu3Li+1uVx
7ILIERhtMdGAubKQCS6wH8I8gGq1pEL4gXWHtOnPCroPLWYIWDsWxXW//A9xPF6v
Oz9LPYGTyosH4hoFolqAwjbA37NHAHUG7VPe7PCchqLpbt1fbIb3TcKKO7pN4sjH
AUWaXzAS0CcmlyOo56zAeTxDtbObZv69rRzx2VNMUEvJgMYmlmUyePH7UsJ0/BUr
egOTvTd8hQbVkz0W++Z7GhnMbfVqB6URPvz5k6L+eaz0hj3OfRqrlAmc4ww5JNSt
3ITwDpfJs+NsjKd3xZd/EfHDNovV9GZ2IXMrwDUbk+dZNisS2EMxfEnkoLbyjFS/
/BNFDTSX1zYScF3vK6UOmloe9SSXPJa+GMoAuNANa3sfGb++b7qh1e/OFCC+Ua0q
gtOdyxwawPFT3bGSRf9IHQNwIxXCU4ACNIOpswF7ProX1tzOKib9li6Zqj7hPNy1
JO5k8irCsRhNId3MVNtEKwlJNYZVQkZogOKHF7ug90ZfKhAYymQkb8722O17yIQ1
Ou38QckInHb1ZDA0BK3vC+AbAiscOOwWwzmOSt8s84sbyAwyCRNs+X3ka74p3Nfa
p+qB4phBGOcsnEcerfLtG2z4FOWfjqCYMPxd8m98jRehO9U10mYwfabjR6yIC3TZ
JxlJnZi3+Qgr1k7LzMDwzBaxV/teCo3JgHbZreiIiFEzIymGMk7vgaIjJoAXM1pr
2sbYu4UixTSB9usoL3HCpW1WNa1t0/ORwBc3P3IyBEAj6xWscU/5YelMMMAxjFxD
j41yVQSn4ej7AxMJfZEpFXkCrcjDhvm43W0QIDV+lsm+IEph/IclraYxzun3PFiH
PshSs5U4jtLsuGEvW1MoklQ6tzV5+dMdhsoCqxtL60nz4m+temnqhPAvm+huZEJx
XR5j0v8s35KeBXV1lzr1VEdtR/HV0sKE9RUenCDqXB2S/5Y66YAmTSRk3lfJZq0l
karP4zKYVQSxJ9mnEDJ+UlskfFaqddOAEH7WaMBbm2nma59/4wUTVBb0x13yUSjW
j+8YLDgm8CYKL7nQQ8PlXy95QTaFQNqJejRsXcMJ/t8qfdJ2Tdg2KM2+27bMdiGs
ZGTjy3dgrbzpxr2YAif0ngZpZCTppLMUTc/rjR0/KZA60MNI5fCkfOx8jzWV+gz8
wNnlx6m2f9dSNO7k/rOUStwhS4c9uEizAGkO68bHp/JEkhAXZLoJaMVb97DflBQ3
Am9DsP3zOnqslLjgvi+9czMQ0JBz58qSwxoggyLqTkrhNzOdFdfWxy+BzJYD7R+N
o+JlTC5rKkvrDKn3Ff3Ahrdq6dJUh8mU3oSCI2uX/RXuH/cEk6RGZ5BbeZpsjg73
Ydi7NQZi+qGZdLmQbXOGYGgaU/85KuFwfAmjOaFozCvjgyfAXAxRIgmI8oYBanLN
mUU6+kPle/WEloSBxcItpNyxinbrEYkmWqDVUukTr0M/l/oCzfOv50ScQjFxYH5m
oYf17Y4YhubyA25mRIgqjBZLPHZTu5FzlSBbGUHKrM439Lk+RlBfp8Hgq0vjDjt1
vT5ohFberWWGmIIzsJVdQOX2ak5dJI2jwYeKAIycUWcFKPX2EBMQmvR1/5Vic6LM
bbT7Se2pXRUuJAUMCqA7Z7W2OLzfT37o1CcKbtKm6zRCgnboX+J1jLMivuHpUxt2
hiyCVIYa9k+7a2st6Q/MkXccqcDyIlMm3XYPytbDoE8NZZ5+IaRRZkv5rvZQpeSd
STu/VFAOGjMVCh3q3L/l/yUA+4AtKEygxDu/4bEvn4Z1WwpM6rR2AqoAqTXqwjcq
V5nXzb9CPKNg5kcd3whpzk1WBE11d/hQc0JE17dDvLJkOH5HzihyhFdTXXjtiKx5
2guVB63p4Kh9vaBVCp0D8PgDgHfIqh0SgF93maVlaBJolKtZSBIBY38Hiy3n5NA1
QzXTWUrj/6flqWzdoNAac/C2XXELi4sEt/qS5m1x6LpXYm8//ixNB8jkBE09731N
ZTqxDHPxOxstQnECX2Q+q67avd991i60rrhvjNvEzdlm29XPTpsnU388129XvEP/
E46+YGf9RFrc3pAQFUBWj9mlA/K+X3PVBUo+tozQ/wPqmCUxH3/OkcMwDBor8yVm
NJYln+83H7giKBWsXlrCxwmYCWaPT/hPsEjPoyQek7rEAszcD6it1tVzIN/xwwut
7q1iXkfRIq4P37lkoSTx+WH7/4iNeQVvLCTQOJS00EKw2+f44BjX+US4vWUqEFvy
HnhjfCslwAMvWPtb/DoxhQBE+r2LefJOZjJ5MmSO/ZmbsOC9060f+yGT7Z7SdBd/
QrBEL4gCfY6nIHEfQO6CjuYT2cKcFaiwhBqDuGG/QqB/82bOLldvyEtOHT7e0c9r
yW+DP/qD+ZF55fai3irNDnJxqUia6fNOYpPRHdrts71e+8/QRNMAF0nJu6Ge70io
CdyAhBYo7JGL5NyrUKA2OCqYAkYbYMgtV7LA1FmVW03XVo+Gg7w9lYQnK2k4mnug
mI4GU5FonrlTitar4cHst7QFmN1EqYpg/bVIGlC0zP0/GL93ypwLigNJ9rJApqVZ
/UlyYGaGHaswiUo3kMtF07yf7OYi9QT1g3FVIQ1L8+NoDxEMUmrmwWPFb/Ls5hLO
Oi+ynyoiLaWbJ38FTR5zvGO+ql2nkwlUkC/AD/0X93VIsJ2eyTfatTdErUrCBzIj
wCttVoTTqU1Lcggk2peSI7Bd12rDJHdbDTd1TRpMbWyoqQUxRWXB+OxP6yfphxCe
GjoL8gk9if0DnGtFVeEgtH42l8nNDsEmHWt7JlSSTo3+/pciKao76lAV4qq2hIwK
ZkonrfL3VSpEa/1xeQX9AK+MtcFul/St3RiF7qe7hgd4ZWQQk4zdsdMUZuD6oGEg
WrCNRoaoXhtjdygvpWh79xLY0BZPhqUgkxT3sEc0Xgkoh26qX5b2BFr83uuOz3RV
A0wTGTgS0AraO1vFe8KhWRIm4pA8gJ7zzvtc7Ey9u4s39qdaAITGxlwQWft2gk4p
iByWOmXi6VX0jVsZX/HC5e9F/xbpvhsWcpGSOhtd5jLz52QP4Kw+CzIbS91cTfib
kTDZOeCMcOmq66/kDPBv1UM8r4smMy7AHpHuMvCUAkZeK+y7/OK4khxyOb03KBM6
vduODLmRCWXu1NxWqdmX694N1vYm8K5Q5dQf8elQihxke5zPylJTWlMToN17h5WX
webz1cEV9w1bfQMpVqApIgsdL9Dj2jbxqGy8Id4iZsFVabPXLj8555JfJn66/g6G
i95iCWBX7WobY4l+VyBK7yuRKRhjGBVbY9WHYM7b2dNG2mzf5N1EatMCYSckfLAY
TzIKL5kBdOtOKfKQelliG9yHsOSvs6jHHNAlDYXn7P76lrivM172AOUpELGCh4Uc
psxVkGAPt+fwwHmg/UIWcZIafCkAXRxSuaTEao3Nmdy/08dlu63fZ+niRvpehYDI
1mLHoia6r4vAq2OHjGYwsm0dm00VrP00Je9aHMo92YfKHUrSGGHNVqegq3C1bbya
HytcNAi0qLNnDnYjVvpWR5x/iN5akBsvUKIQvyLU+MouTNdV0EtLhcPbm8oPAWhM
AMqfPEQFtpJSlhTT+r6lbHoS3UCOWEi2dIeZDp5zU80xJwfv8sxGTUBJPpwLIm2r
O/4FtAXvPMuUXPphqzdjlJr1NvEU/fEbXMhXWbFqDVwgJbcUmIwDyveVfR/PTY/t
ZVR32C1PJEpwcvSxKxzW2rlcoPx8bgjJHIuUKuwnWu58NaBoVoYj5djzIqNNOFWz
gQaViRA3NqFu/hNnVL4YQXuH+IVOS6veH/fkhphIJT//oSqxJc2DmTq5NLJdGEnQ
ORW0FDDf0+UJpgAArtmJTz/24m9228nKoM/D9102ABbBn6Ofe7ThhzUK3B8C3wyK
U4q+T42V+5mKL73D8fsOUq8BEIH7D+F5FGjtBIIe8q2z35cUY9YTrYtX5qzsSHKi
z9ggLMKPeTy560jpnr0JcbN9/8uPwK0emx8y9lCxNqtgIvJlu9gZ6W+nGgrE3ull
kZ39/ijWWwzszDLZF4H6BULrG/sdQLMZFJQX5MN/sPPD8GJlwAqazm3LqgHPNOw9
tYNCN/PkyE5k/HmibI+cUpUDG7gMqPci77//nlBYlNIpa2akZpr298fYzvBgmwDI
FDKNzzpb4MWxmqDV3/eETgq3rz3Vp63zaIOu94uYJsjpB+YJ1sYvMwZHQoTAbS/R
KBbaz8icxbJz6BxSg5Tou67Vkobbw7JjwhZNMG6d+98AVjrc+qJLIHGbqb4eorXS
WIpbrg2mAKvl6vqJI1yDuwYBRz27vph5EPAbnyR8h+pc6ILv3Y2AR0Aw/MWqFVck
dVRruER8fuPRz0WIwOijQ25olZqdl+1/u4/ADTaBJW5hmtrU+xPPyrVDlj2VLA53
kNkRCt62DPzJX7MXKlTT4FN+Tb+WFx055T88D19etAAxtP736wwbe2L5NcDi/eoi
iao0w6JSOrqDJSz/f0lgKRZgtmqQzcUbBPCg7K5Dy3i2dMSVk//LMCp3vR/4ZZWz
mDUYnpnHKbcx3n9nHE895Dnj5+Py3odaiksYJYejPAk5KH1x5zXZ+HqqmR/yPtnv
eahR2sfyyyzqG8Eh59gHyr5U7py1Jj0phoptFAWhFOR9R+N6dLZOQCIRIqjpY+aj
lBGJ3bielVSdoDXoJjBCmRMAd3WptUEwtLDQW4mt1P9O0CC3Q3PODPlY+wiro3vM
3Z9SdSIGcM9giUKnnF3vNxOEKz+3mrubNUkkJYxNSkbt8tUd+wFSJErZJV5wWqn/
VdUuHbC7iqziSJxfTGLmrPnlnM5pg+jaJ5IuGBClfsf4ag6vgMjvDXWkPytZVFGp
B/IWj9uFGsLwDglaYcIckR/6WUFgGN8qHbwArHjZdN4CkqrtfqNJzdU0hA0NNOCH
kc/JxcLqF0FRvp2/mz3KW/MtBgJKDsF5KXtIUO5T/nZC6KqzCj0ZsNExoYd/ST5K
Z7Owkj9XkoZgZ4WlxsuOdrvGq4RozqaSZxUlVYCmxopOBbv/FQxp0UVwnszQDRIC
4RyAbEWdeBQHiRV+EoeSPfBAJ1zAxR7BPcNpKvyJtG82XILSDhQ308yJ0OnTXqyq
iTL6sQ9zTAbhJLbSeDfyAS0xhJLYAreC/CG5D2HSy6wNrPOZjXuzTNZIvPdtIBPn
WliVTFwJGcjN4t/8moMbDci9i83Hh4R3/V6dPQbUj2UybAkE7VWNuk3d1H/SmPz6
A6w+6ceoMSeQoIn7Ep1Rs98Fegv7FRY/HL3VNPrJd4D641u7uo3yHjjuYucFpOIf
y65BYt3Am8y3CR+/YR1zKenGSVUNjy/vHZvpIxZNKdARmZc/WGtAv6BH5vOnUwlw
7eWgt16lDDyGPe3qsliVeLSXAu8wZgGXL/8fUd1YaEZLHmYUQ9KscNWqK82qESD+
6SLtWfFMg+yLAlVxFaAlXWoqkqAWXGBJoMuPDRBupNH5PlT9W7joHJC78Ng7+ATf
kJjVGV8CGK7lLcZxe9+r3eW1wrN6qizBsoIFNWJjTb+hlJAKWuLYti1SF8FX8IbR
4ZHpZ0LAGFyeGOrVamVpMKKEJne5ub9r7Y5ZEgFc0ntDqFDa0LGDk+hd8+Afk+Wk
kUpTzS/J5UUWLi+yqaJQQAjUXuPk0+ttYiZg5rXxjINxs7oQIXv3EBdsTKAJqt9E
SJA2/5yZ7VFU11A414QNKGLfFys+y8R7ytYlUGGNbO5phXNJbPDVYXWSv3K4sqAB
L/jNmOkMqvSgKqelj1q7zz4i1BvaLujtj5MvAg250pv5DAEsqc54u9vLr1t26rZF
Zy7n4puuITNkt92+IdijFXQG3q4YydN0sYYz2iyPb+i1c476GWlWSviC4TdJf5Xn
P21R3wEeFME5ji4iqqMCL6bcLVbeOCNe0Zd9rqwIuXEph88PmGy+zdNNHWD5XTKZ
wI0qM7l6B6c3aimV6gjKHQ==
`pragma protect end_protected
