// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:35 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
r6JCi2X41YkWQHwWqOlIJyscVresruMnW3/Fnb3e50lvOLOI06qdAZrLg5VrpTOf
8nufz+o+bSeqAiuiddjW67NzE6lwiYY8KvtWh4Le0PVX7Utj/nB8ZFA1zB/h8j3x
AHsuQzcI9Sdoi0tGnbmFJ+sb/IjNah/K7tR8gKNGtBM=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 19104)
Ks3I7fP9GmRnqdzERBW2Z8/hh0YZDmm3waFXyQaGeSlcnJpfISFVzL6c7x9TAhUB
QM4rVrG0+oC0ib3guDEFkAoVb6VeijmTLjWgfmpyeORlY5pcIDsZicYigbuEg0Gx
R0AUuhB6+fk2FihPQ6ARn97ruI7oTafAEUKi4oDK+6AuB4gIAMvuVTJHulQ2uy3F
OOZoeZMxThDdoaJc35Uq2hso6UcC5t9qSA3NZGNC1bxcjqNx9xFoGg3KA5ITWiv+
yAUPeMHMQ8PFIne6i7CHhraRL4ZQ07YWwMDVY5/c3L5mij9zY0IcVFBe7s/bLWJp
rpIBIxL5mWPWXN+Jk+QJXc/FYSG5JwNnKad7S/BWFO2WAf++TKDWJ1P2jKQkYl/R
B1c5vm4iF+NWrB7E9pcskjvPRugKeATTYQzY/6srEcQhKCh5fXDaNmAYw5RZPz5N
jC2uZWGSyyjNUCAyp1PSkw9EyCpsgQOiIFZLd8TWj+Uc6Og7VsMUmLX+Nfzhg+pj
PK9vSiFzbQMCaqcPdVCB0hG4bQpnsPYZ6f2n7iUHkBRQQxErz293Uxx2jAUMrUMO
OOon/YHBXAdh8lYlO9DU5Yi6diE/TVUO+SGuTvI5wUUn4SmNxCdwSX4lLtpAzjEO
rOuffVkucpd2GkHDHO3ZjEkSZ50Aw9AzeRJki2+54ad7lmHt2m3jmnThtNgizD7O
J5HRfo4hOW4v0ZHOh1XiY8blh2Vw7jWkxvBHc6JRgy6C+4c81Mjmh7UzSIHxtj+/
BF2fbRvX5dtA8oBlGg0goG4i7LSTIGV8zChzMHxVHIYY9tPmbrAww/LFq9Hh1okW
QT7yRFGWQuDQk3eooygXQoRonKzEOAAolbfFXbFBXPKf+JbR4zqinnMqllq3bgmr
R89moWqCiuuNtLGy1vyJkNO4wOC6RuRKfNs4UHPpa+DNPKO50VBY6KvlqiBiyEcA
wYPvAxzG+r8LDMor+yjT5ZPdUG7RzTazI7P4N81OxXde10vmYZyY4C4oiTkY1Eg7
pp4dOG4JaVH5raf86ppDlzLu8JFpBWh5I4pLjuGgCnwKn0eqbJDqAF5nssnWRqbs
m9F3yKqKZhdy7yPCm8pftEtBn/xI1WvYOdICtgjEFj0uwpESubFWDy+zGcSmJYZS
K9LGgPqh68D2HKaooCB2WgZY7Sj2A+vrg1luKkPeiDWljtX63Gm4y8bTXZoRJP+0
3iNiaLXScr2ljg60x19GFR1yifMDBWN6ru/77yMG8ZNodbA9sTEp21SHpo1nOj0c
JdrUIUlqt4i9CzJjoJlbJPVwgzdx1SZocer990PYIumxgrgMZ5DX2KoewYKw9S2S
OFp4p6nuAs4CrQGbvPjwrPEXaS3UVOiffIuOFH59YpfmwYjBHsJ0IGFeqlK4mM/g
0OPU5gQXyoIdP4+9+jW048ckCVieDojiViZcXY4LDlCkZAju1NhbmIp7i2XB++zB
rBWM+z8uubwVFMdfbVi8btnTMe9hCbwbQCKrCgnkFF+tGCnQyRlb3r0h9a1e8wBd
i7N+1zjQ2+Rkt5YcW0gUm+lPCAvbriIJZzHDOPRdMn5gtpPHNPws4FB22UlKFNdC
eHFhPZqe+LJj94GiIux5aFK0MeSxZyJ+SblDQYlGMT1zVAuX/o3b/4Aj4hHqnKmn
jIiZlqah0pDrzjgJDplrbOwz0RbciW0OUJLny1TQoHpfD8T+Q0bLVxJUwJ4/rcP1
EmzZUTgwVE2O6ddUmHQgwXUc6A57xQxSjRXOVodvAsfwN2Ke6ALQXRD9AU52tBEl
e0z4gdZIemJv8WutHSPjv3Zi8a7IlAk3Gqgt61P5IGLBTlZO5bCrQ7kkjRAUqvAl
PJStauMkXEFHNhjeCU8bWfpOoQ7OrYXTKVSEq9ljq2BqOmGjqqCmQe5istqPFQPe
ygDeiD6Qgwqpjn2xO6FvpgV2yE9dnx7JhM9QGFFL3D+PhXwhswIMRoK+d8rult0n
OIT75okKpocEfMJ7GjEVU5eK1OjaLxXeqM2lrq9+xJb77eTD1r8vTbCjrLidcQEX
w0TUk+/GojUzeglTVjGQu9m4Al4Oo+dTIhhw4YRXW6MOz3k0EgOAfKiPx+seINvk
Fc2lwodu1fChh18XTXOYJBiO7xxWUnqI+hKy+YZ/Sk+oVAmWeql2dpF4/5Pdphcb
wV0Ho2KHWa3EX2H5ZBSMATsxAeQ/aEA7yICGCrHJfchc8DPFpiT346ChMvQfEYAu
QG7PJMeb9q30ITcHG+C6TLs9KNi83PRSbhJSUjzXTP1ezmn7VBYL2aCkun887blh
mDGxNJw5lkdqpVCE2B3B0hLxuLzHkvkmsue5MVKxMukO0Opg279SbIEbovcLL//F
5DjQ6rLtSyfJ1MR7o0YkR2KQUAI9pvc5I6YCDYsHS0gf7q+HuwrdPpKnYZWaMW6d
7l7OZssWY2xoFfwqIxROv8iMDStE7va1MQM2kx8obh55CjZlDK0USxX9i/esVHaF
BltGiEwHXabmXGnaYeSQO4KBpBSYTZinGrT2O9j9brMNRcr5mJQ6fbX1SX5NjBZg
+1nrlXqugjdVYv2nVcfkx4f+aFjIN483lFawcOxgwnp8Ezr3Ny7tqClmsHWYUomr
Z/2SvGyYQT8BnL6fkSDB2LG7N0y/JWXafkBpL46f5GbfGgMAmc4nPBWC+cUHXjBq
LnqFtuHXpokS2JgnYUDf0CXLVen13MfjZgG/yW6MQwiU1YceYytV1hBsKspHQ9u1
oC4AKB5JWqPaNLoVVGfb0frpmtHHRA2Jw6QnsqkMJqn37hWA4tm96sgALCjk3zAh
JgzR1+EkPeZl1b5E+OsDQ99uGWTwUsaRfYEIDUaoN+PZuZzd404W+oASvma1SDnh
x6XRiRHez6BkFTkcuuoSwbSVsIm0cYcNr5rdr9SWfarHXhkN0SPrDRC+Rfd6bg7d
NqDzQqBAjwTZ8WIPEv+twai7U9kau+YdhappOZvn3yuilL476vmUbN6AY1ZNpsuU
52jIO6oaEmp+HGdD40ERfahddLOdxI1uqGolkiS7nLmhfiz6H3o6GVCLbyzCJ5kO
D3jFpr/MqcIYcPFtV1xWMj889GaMcIgegczYXdOAfQi2HHem6mmTUWyWRMg/JO7Q
atIZneU+lvoJu8E857o43rRaiP4Fqmomja5HRwXZsKZAchTUE1eUTg9/iXvAyJIY
JEx/syVUJft2NzNv0m+GxD4TsLWUcxo7TrLNm5X+3PUKhLnea5nTNG9ejbOKbVVk
UMy/HBc1owxUtr2G2D9z4ZHLK8Ww6VMx3eQdbkwCuYKrXL4cYG7o+ljGM8X8Nkx3
KsiiJqwzFZpJlG3CaYl2EbfMn1TQUw4Hz9RE9UEsMWvrMjKX/KpJyg+uDfSrQepT
U+eeTJhzAbm9aV458Cy+KBzfpiVT0wzdwjVW5wT3ob3gEB8oVec65+sBcujTqHf6
b1zYSER1kPnqs4+PTx2+AzJkK9fb3jiP4UsJ3obL3fTKLNHxGvRVct74rsUvSjzE
h3X9PmIqnYU57+DWkZkZlIxyCy5M2EzXQSu9hfDIi1gU6DfVhjejvcwoQAlq5F5a
48WerUwAQEnedkkX6zwumCs9AhaPeVrqpsl61Bh73UconNfkst8eWkMYjOJTc7v1
pjL4rhsnlB2fIre88wA2bMk3udg3RSbl8qfzVsOTCAxmucAB8DEThh0dvP7JsbbI
o2f0L/GqtPpVhTFYeAb6W4JmXBtVRNu3TAT2q7sBhmSFvkJcW/3bvYdGUIfTmn7j
V+sqXQCsx3EGdDYy6OIJOxmonAMlB3OCqYE2b9CV9vZrRuelUSWepQQtm0mytbtJ
cDxTjeeD31eVZUnGc22YE2M/iishh80+3t0U/840K+W3qYKwmEBeSP5PmbaPxoqD
s70Mt5fUJrdvYsdYKvsHxKoLZ0LFldp6MKO2MGt6AX8Rta5UiS+zKmq3SNrNz9rF
Rky3gNYriO2kN5114OtYLTgXLAbzIuAkfKA6lyfTdRmu9wLPDrfoUA6tobH7szWb
/OL8E8Oah6Dx6u3/XNUI2N3G2mDRN3GNXeWuE1SG/C3A1iyftfs1GuqtcA0Rvwe2
/Nbd3vlLXAo6Op+i0cA7DH87T5Cx+GihUA56dc/7zL2GlQynRs23KaqTr9IG5O+W
3kK3dJm8MFZnLxUgD2/x53zczz8LjV7x6/+QJkqMZzC9AusNIJc9CvySPB4Jv+Mx
9uoB3uEiAFEIIZWR7GN0a6A7ARaReKyBeA4o3yYxOLYScWs0okA7fDUIAymxEfE/
3DHg1yyp5JNyjL2Y0gSurAqg8aogwqJ/u31LIFkbjd+eHvLtBJn/nleIkLTbPPs/
f+BE5bdmYljihYdbCXCAom+z/j3/gxInOE035MeQH8LBVkU/PdyA4pSMGJY09O/b
2OcMMslR7aBVbTmy1X/FImYRkDMj4toWhX/s+Gpnv9v7tNHKoCs/vMQpiRQvLQfS
glww0A13hz8UJOMPGIYUmJtVIYi0V7/3UTTV4VtMwjOWIoQZ81vzMRAxLpFnWihe
WAaD0je3IYLM2+kFp95PMiSpgcxXaBO2skLu6OX83si1xUsO3eG3GWTGldyox2Da
3Kxt0MG6gbsZPkgm8B7OhIk0ht5Sgl6mTwDND7Widq38Hao/+pBgUPmMs7KTsDH8
B+xXtHK7x3mtp8P4OV44FEgUlv9KbjfRpd6IJ1LG/L7DuMO61U1niqPQZpOuXEJ8
3R6rgdsw8Smb9R68lx4G7vKhSguFWKMfzuKhzTJ9TAWOdx6BrPdfro4+uLnJvnZo
3zzan1Rn2q5BaVZrFUC96s3ZXVL3kuh178BpSGaYiFhfh4rlmTy7YKPT/SBg90m+
tFgR+J6Ed8YA5iJ4AxcL4VbdrQrNX8yUc5QO2Jv9daRP0keIloy0Ay6kMclDzSpe
ZrKR61W3x4bw5ObJooJUWkP6g8kGBOz9Db65vffrOKUQWDG8FkXGij3gRimVZxZY
SyiTTRsRG/R9p6yMBVn690/4/G51zr4i/QIZrGKLT4zVGhv+1dWED7qEqD5DJRWu
d7po3eS3kjT0Ys/5FIwBoQd/NPthbbUXquQKZPJjSUye3VuCpdvEtStujM4AA5mV
+oA6I0dNnLZMUeGhezTG32MhpwZ6zQMdL2KcE+tKS97rGoepfdQBEJDrUr2O19Vp
paa7AduC83vTTivb3mWwsrkr4d335Z+Rg0oodzXfFpxtdioRq8cUCgPNUB/Id9gD
0xYitxQ2rjnvYTwzT811PB8F1RzR1Ngf6M1OOsgu4mR9/rFyFT1Xun5rC2OEssqP
8Fn2WQX3SimFkEYGpDxwHp/9Um07tLkzxRJPvvWAdB/rDZwNNKMrWrhqlFGUt/dr
k2f2T/DbvUZpX9DY+IzCZX3HZEAo8uquHpp1vAcObTSPNiSFVPH2wpHgF0mSb99C
68h7+zc9r6/mY4nGUs1I0VTfW9Qnw2GNOHNUMJ0PYyf21OhlCUEIGUn5Bamz48AP
TC2z7DxG3/w8/luHNv+ADafPvUgi6t/XihbT+lloCrGwdWQZzHCI4npkCPpjd4rb
v9bIUwX++zK5+HihSj7+wNoqeEIaWHTUsrUgKg1d1Gnbp1Ud+4C+FNi7ftenOfsX
B8rjatr3N6bMCfZ4wsoC2koW4qyWkNqwvuXwN7F/YLATPlbj2b+EWmJKaiKVP7uB
IoT7gHSb/RjmgcTA9Jlbag+KaCXJfBzGGu0sYHpzAgHebdbAeubDC84ctlfR5aRx
z4o4e5N8O1gvzwUL4wvbxrk6kOCfhP3x1BqubZMhhsHM3hpr1iVrYk+mRv8/NWUH
IfPGbnTK4YnSU6gBXtpjgKkJiOrP81cFyNy3TwhflpGHxtEMSRskyJ+qCx29mM69
L9ho3zOxtFQdIqdFd0nep/U1mICZl1S23OItTiGkzjns2ns9JXxW0nh73o32S7Qp
NsPO0GOswQlaTgZpqTCCqeUmaMPW3QtDm/pOwK3Irm5HN4B6Zefp/16L9JF2prKX
xkz+Ux6a2tyWHFh1mVzwn55BBwxshVv1ATUMJTd1GwJwriV3thYYGPOn1yD+eihN
NQAM0C7Tr/JpvF5OBH245Fi8O6Tn1iBxNTkVDzWiTF9mCjeWPYl0poKV1zUu593Z
gIBamKsBJ4s90hcKLFXhKznIi50l4ViEUwg5Lcie1SHRnlRwY4mmhqtLjbnWnLy7
T387HNzgwU2aTDyXQHU902TRrcr7Z0Ktw9k8je4iuPW5+DAX7ITZJqCNXeJGgnEI
ca2/L9siIYtD1G4Vc9GHq5TA/z2RLe9PLJwp+1vxjlk8QiVDGx5WJAUQN3jpztoa
ilLDlryUHO1WdQ3sioUx5uRzi55M+6tiDo3qgt+i1y1ksbrFkPr5307ysvMBFQzw
g08BFvN8P3PyRsmORRL6I/AzENdPzLW21K+/aSbnMhC/LjhexHgEGjQCDJMQZUZl
F9GcHU99cQJ1npInoq8a/ilYHFuyFDllXjn4/TUAcyVGHaFop/GidTiNUUaQyrAk
OyeYMdBNIYyyBaj7HvW+2LLK4XrjlY4d/1ATIwv0sqtfjF7ywVXoiZd2OCyNNFa+
0L3QHol4lrVjYS8GN5MfS4WAZo6nZ088uw5fhTXlvInV+E/29mtM7da8TK6H13MA
V3zsyEaZ1+sI3nT2mlm+ZoUwTYPQmwnBnp5Uvsv1jXCTC5HVp0jvuktZtv9/5bW/
22npRogX+y5btqmGw0TqW5ooQvzpNUy9jExSBue/W8dMiOzmc+oWxKmxgRwsDfVm
M0Xxt+vFn7hBj9S2WcJz4Z/5YD1juTGAKceJnEGxkjuHyYa+5ImDqwD7jZLHPCOD
JPJ9pGWfNvCxoM63ZP4xfgm/Z3/9uU13EDI2A8FUCKQxlmuMJpJbmjBeEjm/0PKU
Hbg9Lshiu13mZX8xCPIZ7Zf7klE4e+jk7Pra6QdSCNbHz9vuRq76MeNLFPAqUuOV
ENgwvJM+MhmBGvSOOoc2LywflzthLGcJIJKWRzygwJ/jrTdVfcbB+oi0NmLT+7Vt
M+qClPjeXQLYNINGK97kIlNPFtKh9Zd6OdjDeo1ciH7b1bwIM96/pyLzCwVIOMqF
5FGITFWlPNx7jzFgHmYEPLchzQnHq9jUpGynkebSBOTZahEH+2XwmL9N+uUoWwFy
BiYY1JbJIgW5oO3Oxpuet9yfZlQ5Jwg2OrQR2IZDqZwLeq8RBUgeeP+nkfDcj6RW
p1lu/G2VEjBra48IhKqSLZo0IR0OMJTahGGdMDORSfnC5CLTdwnSUkk3xuox3Tkt
pNPbo2RjS19EBUK+GXoaWWsUbmj8Q6YwMkchV3sMX9VDfHJVvpKSuWNHFeoQYdKi
+aStXpD4Argp27tHNjnqX8GmOySO9iE5GMV+3VbKovFAME94mdtTUXuhbOwkL3IJ
bbjEfEhvODI8nTVHytFCcoB55qmRq34uPu0vGj0lrhnfJdimv85vZSIAV1js8IXc
xrelEKZ62nmiTOFy5YeqqHIo3W5Mdx/R/aL7WD1EPSPl1xaEzILPdYCYqDdQZld2
Hv1nKfY++8fu02TtGJQn/gHwo/pa1p9LvTG1sJxEj+mXd6rf3vcIM5lvhKZwUQiZ
mIBX0cQarkExND6Jqt5akx6dxq4en2ZcDZkYXe74GPdj6lP3hIwiosDtkkggiw2q
HjoPMm2vMO56iMttD7Ia+Xih11hixbXeocvoD+zH4A9m+Vp1qp7/btyzS5wdjxG2
kxVBJuPVSRirWH6q4oQdi+MhUBVLVXZpGjz0b6/CelDtVqfUPt39VdA+mqzkj0hE
O9mexhkDb+2kRgOIo0o1nCs60eCSpMpMH5UhTHiPGvxRXNZDze/Al3Mff/zKvii2
mSeIUlu7JzCvgKTi5ZTkjPZGGOmlvLMRCNlFp9FAQd/7/MuNwUfnAMW6Fb05jLuP
OUTUMNHGzmgIrEi4+y2mTLmMGpFmIanGFPZu1+oIzLFJWuTDU1+KPBcE6Qb/7aFk
BBaP11soufDuT4riH9d51KRHM2MFCaM00RHUJWsEv4VZAOja46b+LtaHCFZDUMWh
DXm3ef10Rr9iuUMzrXCeVbzbDEDsXM9SQGclKW7Enom5pljhBhhtsSu+C4wJ/+/z
dCtRyB4/SDkp6J7GgH6ia6YWgXO6kuQhCXG1a8KPFTx9A2RU++yVt7IYj6UcpWDo
TW07j5Am/nwdD3JbJ4h89KRIUgBRC1td9y+Kb60QsorB7Do0rl2UgY4LVWUU1jRV
sqLSUzugdU7r24RCyjn6+Swy6pYs6NZPZ382INFWAYx34jOIvEjPzeLxYHCwf/Ih
lN7v637nCGKudqIZXWj9PLowTlOx9k30vL0fClDehijhxnxOPMow94jvT5g+qf6A
z/8jz3sFTIGcDj2hAu7UytdZy2l35wADr7/G91FE2VpNNQwuv+JEQKAYSdBkwPbL
QLCaNelL/ZiMDu/pzV1ikyE9ptdNRxXJ0gu6E5nsGzRwhC1ER0X5cBCftVMLC6Vc
xs9t5nAGDxNuEuQ4qU0jKZRCgknORt0HNgLovsilzB1Z6tuXjRvIPCAPZUmxQh8h
fKi1pCA+OMeO9CfIG2/5uIvvdQLV6NniFAiidOqti8J629GsJA/Ioc6WInKsvIpg
mpgpcp/1ZV513UnJkxLwKnH4uou8dSDnNGLpXPGiVDK52ASQGv7wqSLbc8rmDmyh
xoNXvwdUQDdgBZza93qNskwgsZA5oP7SSHEQVKHRUyIqI2sSVbYYNSCXQZ3mjaGm
ci4Pt8+Axv9+hpupAWf7/jCTDHwYY589UHraHF4ff6tXdCFH+qi/a1Hn3F9k41Oi
u0F1TwreYeknRhujnAbSjfNcVSgh4HLL3jTqQaS24hMt0/hNHc1UvDPJ8Yw8BbsB
S3fkY7C+aEB6B0lOQ+jN8D/+Ms2GvN+nElgvUygH/L4qg9p9zzTL9OFQcuNSnYdk
g0wiPBWRWYNOJm39QBt+fcQnknmIgShbJOMz/od84VHKRWr9bYfgILKo8wqQ9zQz
1jxeHXagifabgWlp47kRQm8Z5hsNjidYlD4Ataej69r6c2vytxQVQd4j44TSb+Wm
PCpTSppyO8eR+ddt8zbtc5p/CNp+6IRO0np8oDaRhfBYfxFAVEI3HUeVsfZ05fZg
hYgwBUcGO7pEA4+szUaWHiKWA9TuEXL+XFUf9A+bQeMeVKt07BnmKaOqmcxhSnnk
Ume0GwMHLJ6xsYu0O8vby2tA5UnhNxeA+jtQq1hlhHxrMuI0g54gkw1KVUniYj6m
fq4Vf3ZjsPGxF2PKDDew5tP6mN8BI0sB2JIakTjgNspc/nw6oUyVCpfOxP4senLm
2PGQ2UFiAggbahDXvIxQHftGEfU1KeuDxXqHXkYLD1g0EDAPKaOBR3dQNDuGu+dy
v7/380riy40QrN1Csa0G/gwstH1CeW6lzGO/uYRfVpscH8XVJOVQY8luQ+JHEnNb
OW1kl7kDnqhQH6R4DycrKZrhH/U8BpEL5Q0ylTGHg8ogQjCYowUOnXOtTWR663gI
hVMQacD7LhIP7xOxvpGCids+N2XCXkdW/Lk4vUtXNmA1dDDQiYlofGSXTXJ1sywf
iKa7eyCySCpYpcZMMFJ56UUY9y5mDWWyDyUCfGJVz0tfE0zKqHJHWFnt5xr5Mb1f
u36w1c9M18Gme09WJEa2BopQG6DwzjGaPnqyfnTY0G8g7HTXh5mlIMHaQ7kqxB2m
e/M4d6Vgalagj/cgWC80AlUar2kPjECHa8rPjeEvlZQBH36hVFHDTMfBEYRQO8XW
KwRK+H3ie9dpHR2HopZQ5ZCk8ncuY5pOhT7bL3qAkPZIzdT9jf0LRJXuLOHYcCko
TqC/tqTGGWaOs4nvlNEFAcWMisWajoJTdtOGYP+9cuMGgqRm/NwQaUmM0QPwDVtr
LsAkHxSsCjim3zAqO/bIQu8s1cXG0Qp6VAaVHr0dECUJGvoM1BhFT5sQV7lCQm3h
tcjn/SpU/xxaqo4YO7RnkhHNZc31YbYddgYvSXozxaSeFolQ6FlngwW3yyw743Os
8We1evZwnuGiheknJtWg+Yeg2PUKCYHSBzAPlhu5zwG2S8QFByChwmXNszY2ushu
yBWH7efeqEJNILTXjRdM4HFriktM3dVSDSbus201JTZbEUvKX4WY8PCYO5M0mAmP
MJhUqzGC5JQ/DYA0HCZSzGe9CR7yUSFStrnQaQWLxp3YuvhY77vqIiyCTrFgNeUq
0ea/gNNRmMp8UoRqI5FlNnzk/ayykjvtaEbDxx5z72lFnEoYgDitNZJhp2aU32fG
CkYzyDYrbtc34ut4LRj8W74X8uIHhuxGT0yw0qn+oY9RxDbujcIFEkkmC9OizW13
Z9PMo1tAFZxKqXm3gsIR++RU2qgKO4wpBGrxs9XqUqc2jwBiKPh1nilVf8C7DX9O
dCOlTtS1Uyd5Br9KDl39wtzRGRYYQeaIcnH0QH85B6gEwuwwDGkpWfEMeud/bIyK
WL02oBcVlUkiNTDFcxr7J5gZSNSt77SN6PpsnJ1PAiX/19ACAT+c4fHiUUxZM9ry
oclAjQ791ivMaSrWQkOR9DssjdkeiXdRbeyLFhMznMHQtq4e4hKCQ/3qKo56xO/A
6e937Bk+W7T9DRitMV/ap+zd0CA1jWbracwsS5p8watqKfQCFnDQjSXTcY8yApeW
l5BNhYYAAufySSl3BOSjrcZJms357liSymsBZ4nCASZZAkZULzLPXMhnJCr3IBgP
gAvxWgEzUUv0XWlHmDJXZpgpQ7wfUJVE/oVGgmXuiaECh2dk2foBpY53Ip40PP77
0M7cV0TBycPBnkQw26i3ffR6DCvq3m6hKdA0LtvE1va6npM+6h5JPL+uifZq7RTg
BcdFu23TasFige90VoFJ2W9hnQ7gjLTi+YiqP6hXAeC1Ox41W+XbRjgoVBTC+bmD
ESfAn3C3nhNmtwGtWmkiFQDKyneHTLrXjqWMFUIPF8C9forP6g1JUS8r/JKNt73L
sb2C6DnznWESvI49wfE3jOqg49BRI90D2NNyzAYllovP1l6+JVGyL/ZfoGisYiAK
Y17BTFEZrk07JLTWAawJKi3AfrdHyCjXRVkHFLu6zQa9KWdM1NG5qKmPh5Mv+YN/
YMMYgHvIw54JEEqJcxHZ5Xr/70dbB2emluTE9tghYf3L8jYz3fLSdE1Y4r1EPvXg
OnKsmsujS5rHT8STa2+6doieruHlV00LnP+WB89In1Irl10iifMzh3r9Az7IDY+p
08NRjNwfbBFCIJIEUyN9MN0gEAzi4WcZyzCD7R5Jmj31xnFBoqH2j8JsznQQ/RtM
v2+gVUb7zYQSCZJ+FSXU4JJi2iR/iFwG5CqhHl7R3n7ca0zGM4kNzGMJRCC9F3TI
sCKVfqxiiGREDqTvIno/zoEpwtCgI9w9fyg8ACDLoYPR2maOL45A7fZsEIAPquj/
/n3fC/5ovfPz7kiv/tnKbI8Pg+Vzunqy3METyhXH2a94oaDMB52JbW3aTHLY7+Mq
ImtnMxrVZ++CA4npnGSwKAEAylQ7X2y7/8mFz1adJHpy3m4czejBlIKAghseazkD
KjLgBKK+eXRUCT8vhBQM075Tm9Mec1JzLeWceDUBTZuL4QI8hr+LNNkpdoDvjEQT
lofJqfp9zETHf2C5pUDFDOVu4rRLAF435ZxYf9BD3U7BQCZhER2rKC7cgSwKwUaa
NeEhgCBIRLZAmD0UVRyyEBbxojuWVv0HQDe3pYGXndg9vsUfVQRNbYWqwaBPEjSm
KWPDZPhTe/TXZnTFnuFS89DG79HsefemXU3yinfJwScwEhyvhi5gPqItEAucWkWE
StuiTMFs05e9vqf1RXzLIPQnwDZkAMAMkIxNDpklwfjeOncPk1k8OesH/SrccDnP
9r0eQFb3FVfVk6wCY4JGDXGlwJe0uVECVFkpymTnIeA/vAaB5d19jh1uCPsn5Rb+
YEtzE9zfBa+w3IlGBxDKYR4qm/B8SEiHg9EaZzHn3L8nrSgvmzWBCLTtFdoGUKWa
VJvRKpgDbpukidWM4R5CL3FYNxVmq3QDBEFxgiph7pN18iUDmLexdKCKuYQ9LIm9
r2oxSWw+H/wIkyhaxpbb1E3EO4gVNsqwaWveR2gdS5NOE1HTCEhI7XP5Y55B+ICF
77LyodCsQp7Gq43LSMuFCVM74UHs94P0paUMsh4lcK+TZVqi5rmWaoLzbny2d75Z
uzcGFPblKttdUmjahYPHBdaqs+UlqcR2I/UiycRFp7yKQmwgyPIwRlMiSdCZtKpH
Xp4MDA8VesM0HBj/EyqHza6wwnrDrtJRLn68HPloPovtdWJBAHSDONx/FddPpTTa
/qrV4UHcbnY9Ki0dyN+WUeH1RfD3B1MUDr/TWmMGWfQYeCSScdL4j3ePbXl1th1F
+sQB1P9T51tMYncq4TBinaMIS9oP5phBh1BlnsRCpKQmUFwyuT69HgCj1tnub+rx
dN7T2+vhFJvyH2IHks2GQ3SzS+7lCds7QaVBW+hOjtRJT5IgWuyBY5KLEHmjFh0a
uLvmEQelaC+Uqh2V7em8t6bqqoKiG6skXxsGvUiTanCN8LBpU57vCOwoMOhJDlOi
x3sd04UJ34EOcJA781Kt4Aekrxc93VApmBpC/Hgg6JsKjoLIcpEuwhjwGg4jrxpN
fBwK/biXX2p0CDskcEkDiBnkK9T+umEwjHenhe8mtmxCgmPR2GosfSjANYUnUE8X
07T6Mm+GU6klaVjeE7imYwzbJwfmpxcPa6fkouJay8XFz3zDKryYVYV1uo0ky0KO
TQu27RBC4J9ihO3on80yYTcyoZ6drVT9jaZzCEf62ZRi0HHIgZ/Xk2/QUX1uRnDX
e2RwtWTVTP65GVtCpvxSbjPl2csFIRE664jz+G/7wTFqMfzk38Hb7wPG+8MEsM6H
vbfJZokdvNEE8oDPiVvXl6xdGze6xyWJ8lwI4DEeEQoda+uy6xr45dqMlAipLglx
4pwmMtkv+7A7oi4Q8q8XCHLEXYTMYmFgAB59ANRCs9ObayWJHrAKBx//I6y05kHg
R2XVBjqW3kg5V7OsH4a2jrnp90DIQsBYpwR7dBfjqN3MUOvX4/W5WXI/rmjWLULm
6AqrWQ9wX67+eCH5YKHngLQTK8HS1tCksZgj9nJKdD/ZKfFn6LDmsmegln/JzcWz
+ZJnu1o5jvtb1LXVcQWhUsdmof/DOxjLHAzRr+5FXsfjL8kD+UUGWxcFe+jnm3E8
WpuQmiNG65KQGywln1zVGNAJvTjC8gJ1R9/QCgAVh4AksOWkaOjW32uAMQDMIpL6
xq2B9VmNXyLQKgsZGoEecdMev8mpZ8wTE/h/gWK6z/i3QAi6a16dlLimVSyrFSRB
s/RNlzYEyXW8ScEGpU65Q/Hlub9bEkwBw9U4j8jhNqf9Hy/7jgZA1tQnGATK9xi2
K6uDKptdl74MPduCcis0Pbanjq2WKyGwfK5NWy8QFWf6ObqWCqaEWoQtrc9pNIzd
knQW/hgMM5h/MqEN8SWVisO+bNnExSjen57Q106vuc7H4XC/mSsiQ7jHcKIlWCwQ
KQT1sj8vRdPKucse3Ozd8d6FflLNrJ2tbXeOyOPEblrJX/rUziAre9nLAF5qV0N/
IObQ34vV9PuNvOclaucJh3mbn1Ybcnjuh8Jm8K/X5RznHAJwGmcUVKli/5EFzPkO
fsF2IIOb7r+jgCqBuqyWtb7UgeRJ6WE65eKqR3m/JaRKj5tkgkk/Vv8wRhe+CXsR
Xu5kabT8n9B05rNMsotBvLy3y/hs5I8Pwwshukqcpw1lT0m5RcvZTb+wgdHFYWGc
aERIc0Kiqw2qWLcE86Mre+FSpjNTbVKOJ2UVHn674EmN575xRsQaOoMbFG1BYW51
0GxeTOvUAzoKZ3XAwwFuv6Qw6JPC/BCtHvS6HmbMyavDV0mB53cs4fxIfeMPnM4y
s9xmxpuQOIQYEgNLYy4OBUgojgKtbSkdP4PIqHfBLzqjIXnEpMQqrqSf0dEnMk2C
pBZi35ecSHUUt9O6jkTuGOmZpNPKmcw/KqSExdWN6WmUturDm6nP+IYv9rOPVhLa
cMSOxP/h+JMmhLVYf6YlFYiIMDRG7p6nVlgkmvn6xUoo9m4CKwdsjp61nMdb6Nvv
W1wq4qDIkXhdEpqLR1Bf9FiMmMbux/1eFoas61vTnQe0YNzTNTYpq/HoxiO/KwjL
cPSSzVrHtHkiu1reotz759yHc56WoyikvpYy6XTTQw1GKv15yusqJp0aMOELXB8x
nqONVebykvkq1xr12UXV7ditqqdYTobWPvvVU2Dy3ssMUo0C67jvvLpXAygV7R2z
WxllZHuAG4pZKJcIB0aROJKXODDG+CzOAmBLhXZj4w90F9tAf/WTbFqenJB3SHeC
TSAe5I4kBjEaC+x8NtJTjYSkrqAEdoXqEmFrY9mAIpFfbqVsPnFlkNj+4lzF7G+L
P5pTav8Fj+9vKWj9JDAOIB0I+NimZYJOI3gFoTlU8RwWXED9IxtWemWPZXvsU07y
K424fuWAY8Lk68Zzl+L5N1hQVCb7k4A0XVAM+Omp8H4mOYZkxDjavPTKPIJQO5nV
Zre5XRVQ/Ux5gepdVZD4cwejYJZRP4065Pow+RDYETO2MkfZVB2dahdzVP3wL3pn
AnqmkevWT9TvqSEHVPyEahKXDfjPPddQyGnGMvUM0mPAbiqCqUUWbGVjKV/i1nbw
iGVlca9PZBRyelWX6lBuHMZIs0HFIjQ3P7Uy+GRS1M1yFRQHRnFzCr1MsvucCZAv
3P4OSueIg4q0LbZKvnkpfQAGW20HMo04k9iLXCuqCpkfBTDNSDzKw0Y7/sXXdq5s
LktYOvbYpWoY8U4Pik+VBwqYxevddRS2HK6CX5CgFn83agsGAIjp1n/knc8fDXHy
Cl7sAe+inKTfNlxUbPCKmO5TvPi57RUZ10z2ZpRTtajI7frTPLbfpjIDIHr0PP5n
1NWIfdMX4SeQ3pNBKTBPfvn7BCpV7DL0PzQEOZ3fdOagv1uvJPnsomwOkQfcMc22
8tjzNOFWTeCoP1FIUpWMMWn2shr9hwZEnMd34BeBaOEsghTqIihWIx4d3bqSdUWA
WzHmTFqDsBLk2u6GBRM+NxKR6CJDac9TZK6u8pmrNpbw8kR/3E9ZUlwG9Vc1HEHN
6oZbvhgk91oBWW3N491lJpMTZmqPldW8D7+HefFSF/UGYN8C+ckeo2gO5xvwsb8i
0WK62588rLecHZiz9LpbYUjoPPTdhSr7uZG6vRLtNszFmUjgheDMg8oDtTKxeQ3i
f9ZUWK0YPX72KP5uf+ZAK52ikb0sw/LM889Mmb6GkTHgk8NiTk4vStk7F2Qgsy6h
0Ph52QHH/omO/R4s9F+TTjA60F84ZWNxJmWUf3IVTrku+cfiWAHL/HzDL9Z9/3rV
G4pnb/o3vO2AR3s0XbfnjJ0qNUyT0Ws6f3uHIiMk3FPUlmTtR6BPC1H3EpITFi/7
PriVv8kOdIPPAx7yj0U3E/j76FbvlCmN3iRilgzi+Kod6e7J6LF0sqY+IQtbc0NS
0y9qDnzIya/5c2HjOnTnBDemXvjFo2JVdB88/ljzMwOxgU+GnTsr6xPVf9dMmKw+
0VojltdXVAdJn1WPxqZyjfUYQe2gi/4wnAbq5ySpo6LEDvszGcrmd7nneGogg+t2
wuktNVaz33kPqOQBqa+jg0eM9fJNRSVQx0qCOuNW+3kWPv3froaq6IDaEGXPNRIG
ZHxarnEdnRM7YkooEgvfhya+b95WoeImy1lJFr7Voab8pOxZqcIdvD5dvCV9fFpt
JBhJ6FA2fuT5yJW9MwSBvlNbt49qkAWIyGUj7opJF4CHg8Ch2zR+ZbIwkeKyNKn3
ItyyDEp68RZw3eg6tPbF4W9tmq3xTEKfNfpFeXizN62zQ0WBPglTKHXvfRIBQ6qs
RjtKSt/e2315yOrAuPLjTRxtrwPc/lbzHXL1aI4d/ohVwZY24IOqeamvXLhLu0UW
4ZQWh24CCKqWTY39RAp+FEbt7hY2ytq31KnpJoMrvwxdXYVE3bEN7CdCMLGkYzOi
/FUVypblaMG0bZJLpHZY/nb1nadg9vd+QUq9zB0NUZ31+2LCEy9MXPIOAcAyGNjX
UkJSdDnzdAEVkkRf+2V0NKPHs39+Auy8fx4/rmXGNioa1iKgIhZIbHkdLZEH/Ppq
uRk8xjtAJUryy0hOWuaSSNee/WQ48uAx+OeCaNjed9CaLofZ1JhmirNkTFH4V/7Z
96TXeWnE0Z7fL2zkjklmEra7uitK46ayoNXv97vBO0flGxM1y+bBv4vNwgziSDZe
Q8LFYfb9Sj/fwSc+yPKWipVaHpMV9tRT0gyS7vZ0XDzGN+UXgpa1u8At7BnQv5P/
SrM2OadBBhqfb1bAFp6fDta6HOaMOgRwu/oAZ3JEvnbuJc49Y7YiYTUngD1JAPpt
V1zvZR3xiTesnWFHKa+gyMFAnKMJrP+Aujge1EZc6DEeFT+BG32NADi+8+WCDLIX
H37LeSXH2Firsm//n6yhuZQ2RgJl6i8VLPMT0WsYgWmAJdbU5GfnUKC7XoXhUFRv
mm1iKi8UlYIP2bFGteVFnjuOCxE+ZmdCf39iKcCWkHLxcUb0Pt6x5QbKPK/JtaiY
RtxEUm0SeZEXoDcf2N/nHfspftPyOTImhjqQ3WfrH26rbKU4YaNF1BMCf3ztENOI
mNhiuy9r9/CiZIqj2t55nBLPE6CYXkhJC3ow1UGNjfe4Y/ZG+Is+rOU9oEJluh8T
gomq997VaJQ24DeWmpV35KkIlWAgEwRjEOxM9eIX8BAEPy3urZxXETNZUK92I46f
xzP8QAFj23MSPhjjk1RdnysqvGCJFoH3HxKZDfN64tscrX733K0AP7qcKkEwqYW0
4w7xsWuXGkahrrs1J5lYrgS6yUi6hu8iNev0SHXaLv7AFbIyerUkG+MuwOiRrRC3
XjIBX/sVnXASvrcyIyRdbzhq/nBPdyFyplcOJyQJSHyRR0P3iO5iBMrsv01npq6y
fBB6SKokmjy/0OqTyQb/kbEBQD+NVfm4Oo15I/QUlG65snT8hblHF7m19U/AuhNQ
+dIfXwZJskNaoq1N8rptudx+XxTqGb2prIm9ZVO96Uie3mVV59mtHSpnPSiUlXgT
9U381amLWsaXzwkFwwW3tes3pxE9mMwooyqtBZ8BFM81gNDnHmbUReydKy8hQ5FQ
6s61SJHf15ZlkIvbWzPDVW8cZ21jV0HR0oo1TQyOZWhB6YQ29jdHhOZIlD0EYXvw
TNGhaB/rQTV7xB04v87ai6FrCxD31bcrA4epUlvOezj2Ot1lbPXkMpY5n+9qZhv4
g0+zELr6kWMj+WawgnpkIG4hb+4t3pr4GY9KRiDp3JFRwUi3uCttNqoPps1yf/PI
6/7TmjELeXXROSmwKn4VZqGLpos4tJHBmXJGI7NpvC4YhIpMDrMkQBJ6Lylm3AiT
r6LZplNue8lE0BcZjaNVSb9HvoyBpg/lJeO6I4vWgZbrkbXV0VI5ij0YrqoJ+J8t
jZ8i99ZccxBxoeLSQCzBUy0hGcYGUJWyVGDZPIxSXknAw+IHWFjVHD46TkC2wMci
+wIO4Yx4shwGZJy/0XFeaSHLLPLh9BtxNx8Wg6DeE3QdVxncIInsZ7pewND2L34t
LFY4VICPkfzSliM2A9kNoT0Biev8it0fUBacPTU66TCyuCQL8oZk63gc4ZuMIakJ
GV5CfMrsM4L520E2vd5+UlCMu70x1FTEhHDshnkTcCTPfo0q//rMbUE/iUJ/cFv8
twSSBI7urXxWFFFyikQnB7LHJrG4/TfHmuJC+2AQjZm3u+n8C0psFX4YO/vqciqR
SsdLBYIMU88mkb9yf8NFORvHs7J039/91fBIGlwYR2rdjOn6jcs5Zza5ibXyekUY
6oE0kASd1gdX7VTflv81AQBFlzQp6DQkasyHY2R6OtSz3GR1KyXG87LcdUpSII35
UJsvruP0jlSfTUwOY/X2zk0+AC3Hwry0k9U08I8Ki1/GYYiLxg7H3dPqDLjgNRCq
8kGGkFyXljb97U6+xsvpBnJKe4AcpmiJWbVvoRRM3B37TTRaxwicqhtvjBAh6me9
3SktnteyC24SYRJFEFTQN4t6boa8zTQhVmV1enSbfR7Gv+OmePDNlh/7Hx3+LhlG
HTWkXgy2WIXtbz4cinfXKxvZCcySMk0L7mVVPr5+GXPmD2BGWy0PGjeV86ddAISU
2Uj48xlP0BGpbd7SRcalP4t6NoAEEOhwFiS9/T24Nj9cwThE367zCcVsk0q9yN+a
PNxHnhz5HV/NzFYowZROyqvVedRBSHq0cvv9vVo28tFHPghrRucVOc3BuVFnYCsa
mGX+doNsjh1UP8eP0sETCrBW8Sumn+qEFtKQz6epJHPZR9wZyelh2jdkxnrIjq9t
5KgjVRK5drIV+qOhBzTi78LYGQ112c6DNp8rW632fPgYEfOUiyhuf2TTzos4BQuz
wAyrgs4zpTnf80OKvgKs8qx/RRW96uh3iSU0KNLBNp5jW4YI3hv5znweSBhoL++l
qxVnjOGeF6NZOydsOwb8dDi1FVQOp//FwJv6eNwDKh8veK9lVqwuSRz9TMPa7AvR
PJvJU63Q6WxiHyjkqkmSXehavVQ3Z9wAiRGjdqt6F7DCLKUhfqt4SZ9AMW40df73
yKVHeuKDuoEmmerVwje+0s6sgas2EV0u/tVSYQVKmX6l3mYd0h6mev1+kd9/2DEA
A0zcxD98AyxMCI2vGSabeAY53ZD8aUAtVKUBLQDNbRCUGE8sjCf0TztAy2ljkvTF
DGK4iI8gyncTnj5HqIjzKp7nBKyHciXJBN2Lcn6yfI7a1fR/G4OaXSwVqFi9IHZa
b0CyIDc1CEZ7BLidlLgN2fUZ5ccaXOjHx6IIS5C7VVasxZbJkbH9nML4rAiHv9yl
YLdQSNHtM+Hw3yEBS0UEpCFEobrvqVBY6W01QatzIIlmQaTyBkxfRRwtascKcWpg
KZ2YbiQdWj49lrX8iH9K5y68r/nHygUCFUyZDQtskY7b33WfKOCIsQoTcSPQiFZg
KAVkHiZzL9+EeT1JCLD+Z5hMnkrmbIN2v3qI2BQf+OccVaU99vxaNtr3hTf1qIxq
hNEcPZSpjQJg3iBKXDX+/Gf4Ew0yYkO2JIwNnq0W2CMDobEAU1TEYeTK4aZZdsRG
RrMjtSY7FjGqWPwO0P6+R+lDDB5rRNqjG6WbQi+moUBd2thQicZS6A75ezaJ01QT
C1fHPav1yFsblqw57Pb1I3b+iXrc0sV/Rg6caVH6mQ8XxuWI4juSfW/zv8OUA8n0
OhghpuQozZe0lDcFOLVHCOCuqGinEu4cqvwKD0TcUWTuFgqVGsS/WBSNiZWEEdUB
7kkz/SHUncwo27yPNxgh3o5jOUbLhvtNXqFSeoPNENewMEK0ZPGVdG76m/CmAVxP
di//Bl0ksW4m0lTeCKeQGBFNjeXqFFPHJ90BHvK2Mf5ozncjokEsx5/FsE4PgblK
IOAoinRbx9FytkqZ2tt9De40oNyhscxD1bTlxyEM3DrJSJWkvxfcsyVBhiC15Kx3
m86o0l4cO19qyfN82vAc8ikPm9yqFiHgObVFfkMk6ibTXDjAtcNMysUl1/XKdfnk
PvBTpaBOcm0GO5GwUXj68dQ+/ZhGilY/XdIRVNmosmuD19V/YqDOVNH7NX+gtYdl
OVcTc5Eelzod7oIKjezrbJ9ZmByiU8ZcbSNyo8K4vgt1sa/dq+1uFVG8RSCLtp49
ZzHolDCu9iAiREUfiDTineIppVDMW/72/7fzyAzc5b4uhzWqIQvkqtGdTuhrOrB7
HKe94uhjUpmO8ibTgNi3xwPrguhaw9MhsVLl0RGsNL4Yp229CtUN6SdiSK2N8Uxk
eH6v6wXAYTvGpyqFuFweOK2SbbIFtjiK558Fitbhv3rFirskQSclrutuJjX8HX/e
dZpNJibtiz66ASJJsRK5ykpobXHyd3n5fMhRMOgDz2OTJ110GGJaERu3PZo7ML2n
zS28PVcIPGEuYptvtzyRy7aDnIfD3cUEvrvCVtWPyg1cZyPg0YR2pjL16JnWec51
x5GJBkxy2iHYjIlbQXN2yljCvIeabEibOlcIVBRZcdN39MNA+0nymDo8x+Lyf/7I
deWF6ZlL3p0l/MD0PBgta7Uu+DzkWxgF1PD8QOCiWh+PaWajYVDZf9iRA3ZGbtZb
o4NjqL/igYqcBG2HRsjoEQqc6ZkO8n9KNrvGhgUZpAIoFCb3ZaGllxGhoguguO5Q
POukcSB5FDo+6Gonyq7tU+3v/uTqrdFkzfUsI4pLXFrjgYulwII+Ffd5qE3GwFTc
PDES+nB7HubLZftosmrEyBvoK/4JGo5cDVjTQZGWyFCy5BR2fhk733I1a4Kxf1fr
+OcJrr8Se13K4sntbOH4BmdNkcEokl7BGZFEaQjkHltn2FbX1D23NJNLE7pFTFOT
FtjUZoZRw+i6ZKik6i8sZlWkWPvIYZTkIc4kFw9WG76RTokNmBOYv5Ote64aryk7
YlnPQ4c47y90ZExqASIQBI2KhVl1PH68iLm3mgVlHFRnvYZuVy9W4Sv07n17xEEO
HGpVQ6iQsDODdSAgaK7mFkson7ht7vAvhXSZnu/p7cny6Ybp80gVp3Xg3Zrz3Ylp
xQ66jrCQ/J+46lA7XWAP1wEVTlVCq4eLcC0LmE65dWm2e2pWtMNEQ1XHw95at49P
8dI+GRcODfJjSxChOHnHdlzTxajZGpZgY/hvOsMhq8yKDB4k8G9JiY+sKJP9GQcr
dpmv5s1XoJW4YUP6Zk7EZQwtaT38PQOZzj/0Fihjy029hGIDrvUPCmOf+5DPBWWe
VzOpuypOUXcyL1uxpBK1nd2wW/9NQmaxNwZehLHhrmxKHiZRWNngCScxPLk9Krz0
x70NCOkReWBTgucDuwdqlxK8K81+VNYb1w3QrOyy+fQD+dIusJiud4I5GM9ohPtK
7Y2s7FCPioGzwUcwl6KoE+fRKnM62X/WemSZ1TGxBjAP7JyBQmOh2NQYzG/LX9DR
rlffR5MsAX46mVtCEVCYpUfj2CkmDNB4JpL+xz66B7drSasiAskQoX/1NPxbeLbs
eXISGYOTbqsbZ8wwV0nAujvAC9Gh940VL7dYvtx/z++WLACk17y4kxvTUORnb8cf
a2L2OBLvDrWaci3iRE9Jkg68oIOjWsaFoGrsWtEWsF7gV6Wvp0Eauxi6to7jFCKH
Imb81R/BqfU4FUzB+xEmyPbr4kEJXpbFivuNI2wWCJcPHmCBYhdMOf0Eyg+E3ihF
63MElDWZNs+MlHFBq94mpPdlaHH5vh+y6MdmY0I5q43xXTikMoR2mHZPvi77ZzBi
uRe1yW/o0LM2CYfqFA9FIbTvkKxgdaNs1zB5J2MOPyALW6fPr2HhpS7tpfTGn8Dk
I4jdNyezBABdenkotUJbck7hjEoQmk9IXd5txYUxSCml4vLc50CoIxBkBvpLt2HS
p9vhTZDZlKobGfYJik45JES+HoIP6P7E9XvG4OyO7b+4AYB8WujZLJH1whGqLlsI
YlGGxRnT6wahBAcUdEK+mDh8djMtHHlQnsnWS08BGjvvGlaFXHGmfhWjmRhBZoRl
uKNeBlQCsoePDNk1+0jDR6sJQ24ouDesdl9C153+vM5XBtxyUry6uTo74gGmQ/JE
/8N/LpQWoTcK/+Lk20sPvBRaEl9QldVqXucUQyS4rfvH22IaPMuBJlYZKQ0SWnTv
NSKd+fKNju50+aMwZBnn2lUefbcAgdBGoMmlSxb3TPlAotHp+M9GiJxCxZK2PhKl
JTbemUKK5bT+FGQ+NbZgt9Dtq9arMkwSWfdaOKiG8t1MNZ9he0Q3stTEXxKMMMbQ
mIQq0Ffr700H0W5+4iGTnwyjZlGdNjqxx1z8De+kwZvKdaePVvZ6mxD9eBdcsiQW
vMYWSMNrZUm6slbKnUxMLgpzCJ/Pw6m3Ko641QHtTfUzYjA3Q/+P9CsP2H36R/VZ
ZykOpFb2Z4JSHtXrVdcWT8IZe31fsAqYLFC8oRF84RQwaSYwsxVvHhm4IaWDh7ds
vp8YCyr4s5ciXhXIn3vuBhKn8dU1n5aMuEhjYGrTETy8Zmby50IfdDcMb+Vd5duu
OO4bbr5yk62+t+cjBkKKvvZF/yxH6WsMSukEDiVZRUg3ezPFMXe33ilqhZB/z+JM
iWYzpiThCP5uymG1T5tr+HdgZ/hMqmrNqtlJ6B9i1kqw5ICx2F9eGCT0D88toV4s
ZUfOn1qn9mxMJEyy/LMt6Bzk63z4UZvudnn9toDtL0J5NlnAyRwxSpGU6rv1Ka0k
6QFIqAmX88Pi1WPR2+IdtKimogy7B1jcnJSlzD/rqJ8mr+j97OAVxKVRJgBofwq1
g4lCaYJfJ4UaFqd+KNiHMPJD/BgI2aFifDyFWoJU4jgfbAmSuKTsQk1U3BThU+KH
llR+1/IzpkasEnBZMvOIqzlUUVEbgwYjqa7i5oJqmB/JOpR7seO616ioJN0Nnm/k
z5bhki0t00WVSg3GFI9jY7zwcYlTc/Df768bTQcZgCSSwiRspwlBHp9WvgWGIA3f
ZKyrU1LibawvGbewl8hFj9YPF+qG0ZcxslJd1Xq6ti3espP9k1Q7vk3G7bZryPDq
1HzYQI7YbilRmG2YIuc+V3ZTJmm1aCC1J+FIQdNGcxid1gz6+92UNZHOYShHp+6U
cPycDiUdHS/gzXDIxda5F9sUnvm6Y6mjsSQntvQ9Z6iqGbnVSn3zxRajPLqXomf8
87oKwBQoc0dPn7OmVYipI3v3N62W7ViFQuzzqt7fr18yxGOgGlPAvWWMLkk63UzN
sBN87dWn5jvqI6FB0zA0XxB9WRLq1ZILZ5csKwZqqvJWsBM7bsUZLKkddzY1aVrC
iRix/EXz0IJtnLGuIT/JFd3SzNObvpTrQbXyXmzPgr9X3HOQDqN+8TuJwlnKbJHS
D+I7VxQde1aAYlbOcPX4FaPiLSqZ6V5xvMOqW0wKzSmMSxTOEHJm6WLlNBaQqQ14
rj39bMOmPCS0sdrbX2oNTa8i3mFBCm9HqG1IGAHDW4j7iOAMhQi4yTO8al6KjZu1
BVCW3h+i7vYDERed5G/wbHt21ghWBC24g8WMn9z8KRyO0PbSPaDIgf5rt2x5r9o/
nTeyGicU2ME5549Nruy0czNBu8zuqWhcio5lKlqslOaoqyAtZ39UdPqmHXUO0S+D
vSaFDVgWwOzJKycaWd1Kr3W4DCj5sG2YBsuzZdmJnHvl2HeKX+2KpSj/wckYqOTP
OMWudkDBahGJXExzLgnlfVGTimYf6Oeofw5gy8UGIoIqO0sV20Vcn5PfPoOnhsVP
cpd3bsheOsZexwTT6wy+ZFL1ZBVsmZB6G4JYKD5ZpyJwBD5f4n66r1tFBSdq5Hhu
6snFjAUvvPZ0SdhB64c830fVZKHB9pxObCbMzN+FUt5LwmFW1S8KmRCThDH4Zhr1
X0SkWjgAVlRmDme86/azoiIYFOgug+5gIHgnNf9XqGZkbewwJHprOiY8WmZ+z9h0
NvX3xjNANiiaM7C2yv0Re1MhYKcgWKMHyfSDUg/MmnFCeFMxLO8YBkpiVDMuIR5j
hdEnbVLndVm0JH/TOjDcisPo2ztfwYBtQTwSPRsys6gzHGs9xgKJZpy48Vf4gMh6
3NsFoXoivZHmtfSH+2+B6VY2xdrOBShCkPgMqQHjr8VSGnIrl6RiakQvIgW6anv0
w11fEmIXg6zhwBCHk6uK8W6wV3Cn0XvGFhylVHNLonFdem7WdrzFfPOhPZXLkqVZ
cJ9+VRtocnTj2fuCdsxkk7Qo3+iqgDE7xsg9F3xQLNYdw7NkNxbhON6kcV0rpTj+
986KPR3LfHMHdq2jrn68MomhJnl6VaomXDkmj7wuj4uEixnuWJXtZOwoukEtaVHK
kgF/Ow1NkIrrDpnVUkirxP7MMnALgrk2Uuhi7xb+KyU2iqJ7CqjQzs7gnGgtFLBc
qDkg8WyBVGQesNRHPhzRDaNltgn1VmvA3Vvx2Kj+m9civ0K70Dee0yirKFz2pDBQ
pFnTAVPXFUh3dzJgXdo4v0Tuk25MHXXsv53xsa9xTT61tHzGm5qZlEfZt7RuAG8b
jYqm0O9q+6Xed+lOSpgvz5fVKrPQJsWd4MeLMCAXj+gnj/7AOBHaXI6c3AgJFXy0
+831ztRXfLYb9GkLd76F4Nwr9CdltaD5CL9X4/A7jQDwb6M/tLLH9ilGpiDaXo42
SBCd+Q9rNr+ZkvA5hTUPQRlcsOVtHKbWk7xbrTUpFFU7DXH3RrnRjz92U8Phrfyl
3dGj58E6y5MRjEshFRB8uBgyjy4HR4TEoTsQKJFSD/02EaPLkdeJPVI3IXugNYU2
AMxmvyzHERCnDbOYd5a947S5mQ8H9fF7O8uXqzIW4CJuYztdOaCTBQPOaIgfZBNl
2SkvDFc+alRMkll62sDAW1KmDKusjZIOvo5JTu7Ke/F7vc3kn6TV207xSri+mum9
XBg4yz6BTU2zp9SVD7qYwNlkc6UGyo1NNW6eY1cZ7PfaGaYsqwu5DTQCf7DCWgVG
Fzc8ARu3ibx/hHF89b6TuvNmLPEnphxECzME5wXI0z1HywllPe4DBh3s98RUtlCd
4uG+6s5Qxd2hg5OiGs/0MnCD6qBMjfnN6kZ55cwMNP4rM+Kzsj5S+iNGcQTnfuPr
yq8J2wEseF792TgLS855ba+kRNtILgP9VqO8tuLLCWP68AwQxkOgzk0J3Se7ZMYX
dW9hkXMEc6s9p8ZbBa+8bQk/khjerebhk595Zs4VfnyU3Ly53KcUOH9c53AKQsHt
KmgDz3JRthJ63ppihzgDDfw0ivAOgyCleN7hoXks6tE3og44LAb73g642m4Y+XKJ
TuKiifKiMkNm3BUuKoiWptd64apcV3Jjw74+jlzdbtj3F2gvRzR1l85H0BDoYqnI
q+oBOwOOj6U/+UmZMvty6/6V1MgHXF9TL5hCE01u5LLlFVCjPlSryqTXNUFNvzMz
/Pg2+d15eNO/+FBdEAGYKfAxLjJ4rXFMdVI29EHYJ6JyGbhWYLCGfIBObTWZdhJf
sdE5qHgwU8WhW+4f6yyPd5cNusi1DSaLbfEJ30P7byIYU4aHWDZRm+cc4R6qqlP+
eveWDIvFTISeJsGBlcuJt60ydJgwN2uSCQyA+sZ+34rp1qo1dk1hUZfD8tcQ7Cvf
GTBGN+iUoBMe7SHJMVaz0yF1QS01NwcV2Te2sTon4QD9Jm3sS9zzaVsTdfzyfS38
LZ6hCWguR6rb5LjCQC2UpriewIX09xyqBZ+5Zip5EViRFG9xcf/S8EnuFaEkKwjs
a3BhExfTpXgvdNOYsmnQcHxvGTcpym2Xfn+QziYhqYQPUzBZo72rNBYXLplbhGAL
WI3g6nNLdtZ87FmM6h86YQOn/f76GvxIFASGMBR7cUAaAhLkwtzGOPHpsjHKb8+F
`pragma protect end_protected
