// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:35:51 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
hRJN4LKV6z3cxK5x3TK9HszJ21GKVXCazCXj19QYf77lkfoYUw8vsaCiKckElcsO
TLn6LBysGQR+vu0hi8stOfdpAQn6H0yf4pVEXP8JKGIX8OEm5WJmv+SqUJNpfoli
FmK7pdyO3jqJ2jiHKvsA90JDvnF8fHJmKMQ4ioyBNjA=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 4688)
aVmrqfNfKGco6ASBWrfLYyQTYInKkwLC4lDq2Kkk5yBm4nZtii5iwzhmXJLsHFol
t2Z7zWWSDLO4cgsc9DOswG6NyjEFXGIhl+z+ohnWJRvXfaJLutjtZFqE7blcqqtt
fncBo2H4E38oGk6pcBiIfeCKlxS1PhqNoWAGax5q8Zif7sihlb9+uQAo+KaSRZag
RWPNfAlgSYJKQBN/UmIOjXxj3GGVCHxR/NKXuJoCKVCyZD+et1epLcbjAfe5zAVI
6DVkUonrKNTHqPus1A2BCCfWX2VqsXHI71OFm/kgAG/bbmRA1MlJ/HL05XQ8CFKX
Wrsm00oeurIJvMBtiUU8HFASxz/QS4j7vmTf+vM/HIyBlK3vDvLapv8LK6FYlcSp
Pk8oxoG+cju6WdUhmXxwDe3ms7ooK5mQ/TEOtt8DLhu6mj1deUu6Iqj08yKa4lXW
5B3Ahl36n6KNArlYck7duCaJRHL63VWvr9omEoHJMKg8gWBroAYiO59SEw/SKxr4
UObND1bxH4j3ODghVPa/HWas2qtH3YJi/GDu2bGZ3ZhtxgrlIiVI2DWX8B3SksM2
4wStEOLMNmtvUMQIlr/TrwNKu31oH+pcjXP7jikg2YEk4FHXjQsRgAcqFD7NWHJI
u+KaXDcrg2l+sDeK+TruE87vHSFdJj3DH8k7aSDHipqjxIakHlkzkai7sTfEVrzh
Q7RekHy2kDdkByd1wtVLMo7JAt/0eG79oZSFA+jSHgXGbx4PXlw76gQ3rkVBmZUQ
tZ19Ny7BiZFWd13eIRnhW96KdZlrtXt4xRv0U8CSc2lj+6AX2xWYnGpS+iWIiS0u
CS8q2GxzT4AMolX9OkYnvN5hO6Ar+o60R3+5K+LnMFD+RE7F6wuAxPZR6otggZG7
JoSkMU0CqKATf9JzyQqtyPIkgqSz5vD4ilJMIO7PLrdmbOld/KDn/4AiK4dps+Ph
gNJeyEv8jUHQ7pns+iyLocwFVe3Ld0dUQwigc6IPXT9B7tWuRujJHbkTfpubvcWD
pqSYyDgpswt4dFomJ96cLenOmkTLzLUmj3+bKLnR4luP9SC5PzcaJZRZIW3LSr03
n65CsNHx7ph4+k+CHian9hcMjbC+wM3z4gPIjpYdfux9OyJqvJeYWg9I1bMDq4CQ
LCVnqzsd1UdT6w/wCwwLLfce2TzZsZ+KKtOmp9A6AikuyrqqkmgjH3AiINbUdlt+
5Pl+TzJj1O4TbgFp6jPeb15/IZaI+BE5j3SMxTiSMsokURWc6g8jFMq8/6KjWfgl
XypVTl0gmj5M8Pnjh/2m4RdqTdtOZTKIi+89FyLGgdK/87mAZAyGll30jA6I9pFB
fXyk3S8RlTsIZGYH6nQiwpDAZu30ZGvqVhD78UJ4wuRF8eswqBUJu6F7MDd0x/G4
rxl9e/SXpFgqnTCIeVp3YO3/bMNEoQtenT9+naoo0L4YwNrlyQ3B7Fsdr6HTEw9J
vEnsDyXwkPGREvunak3i0oQIOoGmSA3rpI+vpCW92ryj6k8MOJ/v+yc5AWLKtBG/
O3bYN43BJDbUmBdbCVAsyrv3fgMQtKMAgvWd1yCKH/HUKgnj/V1lsrHmh7zcj4xt
5B/rQ2pLQqo+DnlP/hmEXRWqNNehDPMA6/p83OIAWAqQgRB+7yGXDaBZ9qb3Nuso
kOSfFNfb7Zu4YuDK/K9YvZuUQJu/Kv8LDtmWM3dI1C0I++6rl8qkkH+VfCG5irN5
U8Kju+5rb8oBdKI1pw2Guc6QOntpj3peVm8bbXDQ9dmwWxJq72WbwqV3C5fxP3Ea
DMyp5oYwQv8xPCKrwu7F7RCMQ7Cvljkakm4X1+LHcRFn6Mh17q4QOpStH8DW8TS/
aVO4zje1u3J80gfYDY3K/RyOIVQPc8ZLnQ2M4lBT14fP6H+DmEuigBp9Krzhb1uF
Ia5OM6Lx3HY2kOP4Nyu7MSoiOGyo/YyDlDmX+FMBuQjIZxR6+dvhuGisk09vSJLF
I5dF82xLwEM8mN/gyMY8HeJVtlHRYTO0uSuBmxUYvCS1a0SCKE7fcXHndb5suMrn
7Hshe1dHf1RIiBLd5iSCf6WKP4dJQQ0o0jCs6xatoIktCS3iKOi7yKw2ygzAFOly
5H7f21h6IFi/ElXgMhIR0Y4g+5oXItaMZ216b3iQGcCjvcsa4I9pBpWvqWjgJWuL
qb695lNr0drhlvM+L3QFR71FlDRc5nj4CMtuo6ICZBFbUkTBIv/QhZM8iqIeI8/j
0XZi6z574JOy38IWCzfo+RB2das7sWghQFvy4fbpKNS6bMeZXtWyRnnRm8xThPfW
on36NFRA+T3rLFWIYwpFWWOsuzrITn75SdyjhoQb5ZZ8ubFRBiZs7Oq0eAZc0ohg
PSFcM8caTbCnLEuwdBMZMMhNbIgQWitcwjUwKymEln/kmj2249GNwL4mjtLeXrA7
qkMxhyag1KCMp4df91p0JplVzN3wDLkBGDxx/PZkzqlrBtfFgn2navc4pbzU/AiL
wazFbAdkY/3w3oI/wxpszoEG5VCSsc+Z9YDAORTptFptplb7yGJPM4kDHdZj0dYt
sjdbzmmFS9DL89IF9x7gPfag85dbfR07JWBSG2dirxXgK0ER5r8mY40Dj8CDDxdJ
fYR4vgM6UtBN1CkvnTJniGZVGTi3FQ9H0suJpHr3olqv2maJmi32ItQ34o01rtmg
Qp0NqNzl0l0UZyCtJXv4B5oHPau6SUEwv/dmrUZ6gp6TkZtag+0Ha2NH+J227JMN
QvKU0UkaB9yvr5ZkqkbB1nHp6m1h1zLI8xt/Xa+cDec1XetyEBuyZMDCWKbfspFH
gFo/VtlsSAwCHjtNUC4ipYSi8s08Tf+9V9mWDQpUE+CsNgeQfsZxFbzhqobs8p7G
oxTM2yjWPy7N6g8aLsFtsmjw+hiXlbfYwX38O9c+GX7+yJvMMoy91Cj3jPpAY9JZ
ZCdC15SSRG3ERkttws2QzZKXkGvu3aWEObScvmnTfoseg6UtKoCV0I34f93WN1/6
CGXo7M8yoiskcFm7eTE7c+GF83BcagsUa4+SkLgJX9CJnyjJA1ZoCz5xN0owInLx
g5++gE3uiboTSIcPfcKFqvy3GmEwqvc10KUv4J0t4siAg19G+2257uWI9iAKhGDd
rbNSAX4YId5yjb5bL36McjQk6h+eLZU+fuvGEvO0PIpAtgbTTxx7h90PsyYpkY98
pP1hwvIt2qEF3pnghvGE0vRyNzhVA8Smd0Iomv/DGLpPUzfVp8+H8U5amDDKPgpH
ki5HAXcwc+mTi8BhT/L2ll7UP8yZeGHBkD4+52jDn4/38hOymffM7Ksa2fF8lhSe
GSungJH2OIZKthiQ0Ql4S90uLKncFa2qylJ6TukkyryY/WtmSdn5NTpiqR9ndTzj
0jfUKtqjaMF1LR7CaVbDESRoVa4vHRVtAzNwb8xvaIEd4XNT95Fwr4YtZIQBT0pU
Gsiol/H7a0143WRJHvMJspFXL+sEXuJSdd+JwR1UGzbycLn/9p1gumJi+YEN3ged
5yvyLuVUCM19QrYBQNT1b+gmyAgj+MGBpE8/RO81Bw5VaXJ61O/UKbybUDVI+eSs
RJx/IEwrLvGh1aEdbjmlbNlZlleY+O3SOtjV8C0B3N3woV2mnrcjL5N1sR9YSjoh
O5WwX6rXLiND0sVxkmXHRsM09Y3+pZC3rn5j8VWjJW9Aa1q/voJgc43mr7TFbIBD
klRlHzLNly72l+fttzeGiCtnw4IguC4c3se6YUi7WIAFI742L7YTurQEsWHbwWyR
xJMBHix/92wt7wY4ZeuwuvSqXpf2I+qkHt2g/Z7BXs7ZXqs6Q6r/efz3qYTqdNlM
uSsDaC0nTnSVcB3KlBwbYVgJPbNDarg2g0zn7UxmcB3hgDOMFlJ6dOxaErVE1PKb
9Ksa1/KiddFmG+aUbEtCyJvjYKDjQocFEyXm8ByFNSz7SnIaN1AXbuLNv0r34949
FXswon1MTifilKf1B5OWopNbAd3wnD8T/PYsXQbyrq6jcMt8x54FElGHfKDwlTeg
Es5soxKIw82tejeV/NgL7Qn0aL6MP3mJkAtHWL0xpwkr/YkHzJ1y8harOcg0ge9t
Xdoxae8i7IYrChuT6gJqGW0/e1TVDz7zG/dFiqWCBDWomeMaRCnEN3AqUdFY6zSU
XlXJIUJUhtGWxuWGHockFgRiBJK6PR3BE9ShnDFAobdolfrZYvh/NBsJ+clyadlz
iziTABDCs3wCap9lwuYTFbC7djszyObmro7R0OhckrlJAlIXA3/Gwu7O+n6u7pP4
2M+SsKNqIL8ylGD2Di/ZeKrtbmROOFG8aXGGRv27BizjiP3iA+2xgXEn3c6vmOEQ
lk2VyOjxW4y/IBLvr2Si+uacm5woa5gPNY36x98L4maqyjdR8Mi3N7CXbxQ7i7Zv
72KwOyJxUZdyAPkLbxefvXpWgN2ILgdWTCIWdcBEs382xYfHdG2OVXObwB8VL7Nb
a1c32qsDyDF3wt+rlflPyH5kIDC3ikM8z02NDd28NwHERNPaenokqAKdWWr6dVnf
eo8pVmHT4PnkyfDo6wRd9YBnSojcDmD6Jgk+YeRQlQ+brVQ0hSKpmHVqF85C5Mru
UGpXcnnUawPTJkChFiQdajvvLZ8B0asw9dOe59ONiU37y0x5ZH4rDlgyXNHdDGoN
rpeovOnvM7FTCITd9QgznetKGygrEUIbpU6Wr13MTiATstvJM8ZTUC0GuA7a81ym
/7Y4y5xHaH5KAcg4bBOXHqSNZKlLadZ2bWfGe+lDteKDHdhSRJb36fvLB8ORcV+7
3bo9Bzp+Eb5F99zXWxyFXVaB+eEHosOxofm7tYYrhYZaHQfN0FYWEJvGm/x7i93I
qPN7WwQ08tRbgO+gYv19Z5zVp9BJKuxSYVGWdaAqcXRJyUZM7tc+ZKRh5Lj3LbfQ
8NSmuyKqTywknY3AR4heYrErQnU5cOrzEu8aoHI/2PccTaBzeMI02OiXUrwBk/3n
R/Qd9BzitrFJqDui/VMRg9VVPDWyi8EmghsyQ6AaGzads1RRDGl+hdm7jW/eqxn6
Kl4iwkAbMeKVKWHT+XTOlxHQKpkX+jCqMmQoI2QREvLekJOsRkFAOjOxlTZpkxYR
INN32jWev5eUITK0iBVZ0uW1I8vrCexqdOiQT10SeR6vUHsEOUsRAjAJL6JPZl6O
3wGUCinb/ot5FoMgMoDb0PbnbTi9T0iVMeelshfRjZV0bP4DWdTa8iaJJUlv8ISK
1VCKHLxcV6IrZuemCZsM0b1XdvFZwhUqc+xfESgD5aEs1m2tNUH92aefhtjOtcq5
k2Lxg8h0j22fPSUbZrnzNojDq90Q92mnIIJdE7hOTaE9R7rDyRepT1OultVd4JBD
Noq+8f1rBdnAqIuoWqd2ihvFwKQuELvjJQCH8BJ/FpWzoVDG9R0qn4s0ANs27t4t
0oHQvDFXQwXoHrl2YRSgDanADq4Nhvt965hdigOZawQSryJdDSblt/annJ0+2R86
Uzu3Pqcp5kKdjxzKYWSu1lHHVdDXxXacgphYYZF6qfmIXTVIlwZsr9XDVztZCdlL
PPGrfL50PELVOwpG8Hjuh2yU3nzYfOYn9Hc6eUMzhzSGspX4DGaw4pAosSfcKs92
xYWCarF0sYPtwwNp1GmBr9RWC6goS2/tNhp22xDvPXFsaZ7UFSdRlYIaI/Y45cZ4
fcv64Zn73WZy/6/uMF6QhrpZa2qibXyb20MOIXVfJpqOppe6Kk3fL5jWPP7AD1EP
i6p7I8fiTh9GKn+TiZ/4k+vw2FpTyRugq+OzD+rnhl6ssKqs81apLXjDRCIgWbbY
moy9EJwjoFeuim1CsbFJ11GA96jDWUyPV2d1eRMfqWRn0iHUO7aK3ERQEiaBxAjv
h4kHx3CpTUcBcaJcRuG+eawH1qNGqSjm6QWqkyMRGvXtoUQ8gjpLQ21XXOAUrfkq
GwxKkpRm3xsyBWWHwqSItl18dYv+DwjifGBby1DbofNW2HGL+PoS20Y3RvadY1rX
F6GBPt11hH7oqc0uwGMxbocVwMQv02zIfGDN6hu/X6bmR3AFhxGav/qlKnvHV6It
3izFS8RxzUpP8kAKm82psNQx1npwJ4NzY4o6+s7N7N7t/ApZyxxQk7Uqz+UJ1B9u
yFYkY577fqvh147+1AdpSfzS8pHTzrDa+g8Bhtks+Se/jyObdPid/gdvU4dt7AIs
VE94pr4JYxVDnb1l5tHes9y/s7q5GSbWrHetqk4X6CM=
`pragma protect end_protected
