// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:35:25 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
LVYPK3RviUEVYGVwLG39jay+vy49m1weOTVl+RrLJFZfZX9GR65fvTlFdplWkLc3
p4xZW6NzLiJU4COwzfCAl6YeC5DZ76mRpbpa898SvmaAD+fe3kd4Z4U+/xIjZUMu
Gp3mU6MnHFX/jReadM/xDzUDHuc8zZG+PUjVcyf4Di8=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 12560)
O0Zbxamzv6kQ1JSNJnCTPI6qzIL0p2TN0CUyLb0WzFcFq+yDBktjZLGnPGC4scmP
6VTFnZmvfogYyRJU57OTuKNPrvVVSU1tIyclv6y01guJc5cnDsWNVVzO907yxept
XIdQ4n26iNpVXay8rwwcCbIreVFs6xw5g8FeqFjjWiPM0KQMLDc2yrBJmuyjKvZu
qKXzmDEY6aD/3N6BNQyqo1HknPiU49CZICtBcRiSYIUTGbQVdHjIYS33OGAXouID
1IFiVsqkP/HV+Azvc1ZUTTUAl2jRMMmqiCdnXghOi5A/NR6Z24OvLZgQs3httEV6
lM+pamhzAoMHfi5fZxjknZhpsFFmxXCdrZH3A4CIzA/tXETAXp5JSXd8oKIQ/D7V
IdGybvWpxlVr3V+s4on9gV1bx4+1xY9fKaz/uOpunpvxyCjXADJm8BjRi3m+dFUh
EBFFsj1mLOB8w33hSuv8NXK8uo7jH/mSWXzpTTW5VGCYTmI/4HcPkz5TVARYRkSV
Le1y8LbIuOWlRtlTaM4miwlAm9iIsXbt48Ud+sH/4AtrgZAg659ULBd7LqwKzTkT
hTbL8RU+aoEL4NtNwI5YFdouX1gqkcmAJwewiNZ1wpnSYprmv8YzsgKM4ckLiIiS
bto/J+pB5/tSKFy7SE1aFzk/B3Zip8brrVp0bfH5Xtilt++ddvCpeh9kLL6JtBxx
IPnm9JkFpmiGt9/ekIEbF4TXNj/OkDBWVGw7LUSGUrbKu5SZg2oG+58yADat9LML
md8H0v0dyZIcl2o2eFT8Io3b3zKuAPi7CBiuRFOfLC1tcdmRWqHQ9APHws+ZRCrP
jrU8RpAxkaLATd57JsHqB2kK69Ejt4KzUQgvwsVWgj+ET+AFSrOldLdDciphJktF
8gbORpg33eHm35+m3TzIw3adCXPK7eknVYVJatKEYFJqPll6MUZJd6o3AWJ9U/zR
kF5iwjdOEL3U50ywTttxlEGqsGoVF6xTKP7r50cNX2erHUwjUnK22OnTvvsusZ+O
CcxrGyCPGGZJlHGz8jDB+W0PNrEQV0IsOjNNm8WH7Iu6YpDRKogKGs2VgfUvcKLQ
ZvmXpn38RzCOgGjFr2L3UiAkhPouTKTM9FH5W4WDVXskZCnjQk6QC/ssisekagHW
TFZ/cIJDmNDXB8dcUD0T4gepwGWm73G5cLnTlLhFV5cFyr9mpBL/2vw3uaeX5K95
PZkjGaiyTmBPaqs2kVg9iHpcQ2VfhU1UH3GNbw18OAJ4uXRMwK+NinDYeRfwQngd
87Ozdo9YnBrrHwmW8QzIKqYHxC7Yq38/0zU+y1SVqdB2bxuw94dOG7qMX0WYzkCa
mG0oJc3HWIMsvrCIe2jYQ97NaFN7NzsfZ5oR/zTia5Nu6ftpAC8SSb66Fv+P9KnP
BNLG+WoIQXgOsPF8v4N5qsW6fdXUs4JTCXVaoIl7VAUDVsPAh/prc5m41FYRQopG
ac/wnOWqM7G6fmZ4BBIi96lkf54f5Eubv5MH75K9GcH3AE0i755+KB/82DMv7W41
kRdeFFawoIR5Wpco+mL8iQTjIAfcTt5AMM5m+uzbDSIydGSVj4jvE0cKRORJcc50
jvEP9IWfuJBwqGgJzSfueswCMlcs90f/9bekEfBgwobW969gK3dPM/R4yNgtY3a8
a2nlagjJHRlDdEKpzsdRNaH6vrW2fnn3tAZ+dTxDOJiHKUJDcB2aNqvxwl7PpqzU
NEL+Was69M247E9T5hRdpwtvTV4AF0VJnhP5WBkXU9d95wv/S67qvoAQBu1dMz0G
gKD2wMaCo/lb+6Knc2Har5G/yLr8DQFmDb4fdri+g2QMiXyP5voAg/0uGTLavaNk
ahrA4q131zwXaeFg7aJzeOem/aORJwsJPfJFz6dwdHo/g2lU/Ij2nXWhyAsMiYIk
gCXK+P/6z1TNC7XeoXXFGqGcIOSOSn6avk9YxITGj7C9n48RUQ5Kk+sP0U0KobtI
zaY6xq8JvlBNg0/DbXyhzjGu6wFFFCkRvPQ2BgscCXZjhTp/cATQTz4jjf99jeZP
FTLf03cf8Gn+2W7imixK75TYyriFPIe3FRLeBmL1r/nmw1PsbRY0YKllI6SUjsOs
Uj5r8FhurhqitXLs31XZ/aN1x07zTlFlS5bKuADEIJFoJsnW9iEpAg9zoAcY1E5Q
2RniYpEloZx/lO/LbFZmlpMB0Ex6nn4z7dDUvoxW10cvH3dri+wVFsj5fb0A27sK
UoIVV/RVn4cIrM6zbgZCd8ckYrLVtiLKTnifUws7D4b8HIi0vzubsIFwvYsY/y0y
5stmOj7WbmiwzaS+D+tljgsVYy+USUCv9MVc9A/TViYe78gquUaA0xddrMF26E8o
pSZEuLa6yvVhjTWaTOgFLDUCtFEhbCac+CqTTva6zyU57ji56ccfBzipCO7f4I7G
fMlMbk7vWyOM470fTCY9bxtW1TuHnHn8wQ4aZUChxaUaILMvuf+gtIMJzGoa+FR9
ahOzLaPRBat0/X6f3+ZVQ7NFFU4xyWhkvRzqxVE+vbpP6a6ARznlXiKjEmN1gs5k
9NEt2BRXdfcfN1kFSTCu7PuKRowe1LAFTp9y2shU+bGpAgFIV4y+iYZLHinBwVI3
z4gPjguD3di+VFvvCsFJWGCA/dQo+Iexa4Q9+z7BAjRqWNkKoh49MFw+x/c+5HY+
HU6L8fM50Nfdb18U54/CmInLY6vHgb23+F7YdTUtvCfGmzjOZnq/QX4G04T8PRGC
aKk9h+jG2cqxKDyI0ziOkQ6CORsdWmp1CREtyij+tvNa9ZNXyIxEvptS6gkRNkb6
V+CwnfFdhlKH1eNzYaR90QbwIYyBN14gP3gLboP4Yj3EJP4h98woT4/4HF4e7/k4
76c8Zpcad58p4StY+A4h8d1vq78YJs7Ee07awyG2z6cGfDbjAAxepd2EC6kuRE4b
oSNomPN2Fn3ElkdLfGV97eqmm+xO1tEAqGAs3YKiKPTLh+kczhbWlgE7olYaxQmr
KDwpL2hXioj5T1V/OqDotzcLAko05PgcCbIxfCANWJPpAR4+kBi/szbs6yjUh9pb
reHawuGmhtm2qUdo7d07toqQSrf4H0JEorhE9bw5XQPUuTG0fA7DyW9FUQyMBXx6
TKXQsBvP8ZDsHxF5UmHhmpw5OObXCIArunHATSWvx1AH7GBaWKkzuqhzhf+dZIcS
6NYVxzL+0VNng2PoBAmWkJ8gsXH66GVRRPcTkpuSJELBt6mTpMlRCL38KGVEF6OL
CM/GTZ5Hp2g4jw8RJBeoRY601YLVCFXxwes1vwnFcMIPbAf/gOhQPvnny9IczVcK
YX/mUBhU6VdRCMC7jnAz4bb+aRhrEsRMQZM/6IjYnvuKr9A67/M9EsdqZrxaBHs+
81M65ybXcC810k7bB++YEBm9+vaDID91KVv1pPpqHnrri5CkNas1S/qcGGq/NxxW
jnPUTPtg3Smj7laspQyqlD77TLzsag7no7iOclGGI6HE3G/z+mLuLar8BQoPGO7h
34sW2O588VL3GhCqZrJCclzF/CMtomZBeyOGCxMwHEnbnbUatiGovxyMZqWivyf/
G1v3tO/N7O7pVhbWXIoUthZZQnIhQdzUducoX0EeLV3qEwOi94rlp8rCSNrix4lH
DdhppRRUC2htAs53kvI53wKB/4N9MMklvFsPTa08HGSQ0gXba6qEXD91R0pVwazJ
Ox1Jth3NPeuIx2GFVUJyP0W5F7Wg/7cPx64KhkmmvcT8sHaUyHQLZRnNldMsCpee
RBCSbjgfiHYOUu25aN4nYktla7hthsieT5V3kZVRkoSTiw4Ya/0BCXeHmsfo6K2V
Y24M4Bgx1lZUlwke9O/TFCz99eFXeyt0//HxVobKpwRtPDWjaM+iRqoJAx5qeG5e
DDiaD++1HK7aa7zF1zpURB7L3qaHJIT1ggEyhMDOTsTP7ny3Jk2ku/vFV4WnJKsm
Qq66377+cHiWxYqS7NCFh2v+B4SqDWonykvv9HSzsHKU0yPAPYmuAlDYrJhkybOK
vuh1EI44e7FSpCXWn5mHymVl6ivIqOeGoSzTEDduLS14Yym5tkuCGhTw+rITcMRL
iyTOpTd+RCpO2pEcQZy8jQY8xL7ip3gJTVS1s50P0sgrN5nz+uHw02QsIFjaektr
xCpFd9yL1962s/1nhEDrcdtdS+OUZWNuIZQSP9tCcXO2IF1WkuV2FW4Pn/aMJZju
Mv62cIfcveestNUaRrbNK4hkYgweWsIaP86KBwj8Swy6m1TDkRTUlrpnz5ALOcwU
4+BzfPSuAD0U9nbFmZQoT3QNo/kMFuvVS92zDnfAD0TztWbJidCkoSJcsCR3xhER
FhiRM/S9PA/9dOyKCwEirDHweFjtxBFmvasL6Q5SeJskLhomNcw388TsnVQTfEwh
wD0ezvvEd0rEVXQFVZnsFxiddyJQIUewLifP/ZX7XEUmbGbAcIYARvGGJkMgZkSP
xF9yyqdmu63yhBlxHgMqauFfAZrUqKpzMb6mWrML0bv4AXIcXEI/0wP/H9s3i7GL
oatsYSmTjmddMv2fWnMIx8YshYOkFlETJqpsa1eb46jSdVgpDIbQ+pMh+I9MOXeq
7799qKg3twEfizs3FVD2r4HR1d0vfTFtdX3SYztkch9h7p9CWQP01UvJOAyrFklO
9TFZSQrs/r+jOQl+qeqxLVkZps9gtQT7JzUJYVgfRdYP/2e0K6+ja3ERJawkNZ3q
6dHjopkLRnKqEcx+ZXMhG9/6bbhTtJJnxUJ9kQDrYJT7zGR3jxJokheS1AYoJyfl
3yJFo8Mio3Cy9UTs7P8Wqbs21Uwy/NH3oVaT4tzx3/MiycB47vrYM24qeYKnQThA
1RQ0a7CD+1JtxKOW10DpzV3woruOcSwP16RUFfyKzUcB1RvcUL+Ufjcu2JWokEJu
8F6EsnB5pM78Oz1Q7BNVj36vGh1KezGV6bcLSjsUKKkrD1TZ1Cmh9UMi7SAO2bNu
gvjXbU3vHidxp/zfXrdSPB2NcB3d+nWrfa7MrkCUPUa3WIiDjy/8wWapOObeIa2g
VzMyMdS/Z+Smm+tssi8baCo+GRsKWKRO3aVr9zY7C5dOSvh+3oJxaa9lLFUVFGnf
5CvLB7JQkj897MTM9j1r0AxAQdbu5hH93WNlL97Z6aiTQNquJrFgeCV6T5rgmCLr
48hdg5qhy4H4Rr77r0oiY435gMYRzQUE0jxlB+d8UQDtgKJCZIbWbY8C4giKG+88
GuOagcvoFQSBqealnu3u2L6z8xSI9gW5KRfVMM6QPj/S9XBjKF6Ya+PYvllVqSFC
T8J5gRk7f+wehhh4JbwXG8sKfNJzyVrdvlKiwOpmR5YBLmfVypU82HDCVFbLWXWO
9KvgdOgh4l5Z7F5mWlpFngdFm8vhAuORt6fZB1/f0RM7mV/qGi6dun4sj++PzdTf
OxLTQv4g3kCqPQSQ6nPbgW0LXS4pKjmwX/M0E0e2A0QiyS0IaRLF95Qz7Ovbk6P3
QK1XoMFx5/EPyvnA/LCVjDinV91n5qdJ2Ummg2vCE9fqYTtcoG6RgSZnAidgyO6U
KIUB3D7o0dkr+z/xv6waibH/+jte8cRtmMXewo9N2bGBN5+LxJdj3MJ5ZQuZn1Up
lflzbwTg7KU/W5PJ5brRtn+dwRtaHALobmmv/SnyN2+7BDMvJy+htwXlBpPQfkpn
mZUQNPERHk/2qjItqzwW+7Xeo0QaplF4+/oPAz2v08qVV2X/mD5TxDI4Tip3yBSb
6OSYIfUkNJnM5k8w2Wzf146FXgMs94ufC8C8RWGlzgYVZKmMfm2Zv3Ix1atIrBIN
bAo9bTx04PH60cbuIiFMgffk018ZuOM+Du1gmELWP9j3QYEBTPAVxvUPkcsC74Q7
uvOS8kij+Q0O2Nqvw+aVrXwmp+XgpsA1k6IooR+yzluay5WzNXUatUVYawbDn18H
vX0XzC3YGn04ymuJpOZek23L7TFJg1MTs5zCTjijKsR9Bf+xq0ocJpTQ5Hwpme1w
Z0qmmhIulDjqhw77CkXxf0QxIbG4tFOsRu+llQv0V7JtUBpqjXLfoGlgTUzjnVaA
s+e6V7TmiKWMN4uTpn6+m4qhl7IKqXUKgIZb+S+VAa1PzaFYlMkrl9fRLDXGWu7X
MrfiB/6oki2vAsjDZz5PUL+08dAitYorg9DVY5U2Vk7Z6gvpoaYIGCUN1WbR/avQ
xG+dRLqw9yXpJmhHLYd4XsBJG7LpJQapAexj50o7S/Fwo8Ed3Gystwfbcu659y/f
KKJmHJtCR/4tQKSjj5/7QK15IG9l1ze/aU8HZW+LDcWa3GE6y0uARKn+64EakMOh
oHs5dTfx21rsEFIOv+j4QpONcG+aPpXZQQXCUeMOjUDqB8kQ4tVO+5CMPRfNm8So
/sVKzVayz1frtsxJUEIjS71QhV0LkhR6FqVji5SRY8ToLoprn6lEvM66ka00/FAq
wPsibi9EHBW/9Re0OKnoCN09ega8QFJa/O9R6dco7lJE8GS/FlRsdUN4JmI953Mm
wH7cFB0DlP/IQkOjvF2xKSu/s0p3xfitEqN2Fd09YhWd3mtIYDDmS3UnGE2sdEqg
/hJRvZ3/L+SF0GQTUAKLImZQScsY3Z4miK4wqwM8CHe3a/rTNfWFDBtZODErdByu
QrLD8rXFXM8U8UzOnkCzGIzEWE5KdoanPtTVhrdUEDC9VJ3xf5iO7uN2LbUQYxUd
z/aqy84dcx07e909TVHdmwbvWJ3geib41dRIcib+ep39wcR8EYBbH/seiAiy1nGR
0NHr5pSVdtu0Bz7i3Zz07eOWxxvU+X06PXt7CdN8zNyYutgmRSiLCQP9E757mPeW
JFS9UoTiN41GePkK4T98Hxk8uQDErojNpoVsake5vjEYgJP/AfpLgyfNiYP7Xqxm
96ROj/8BU6gGPxkR0sNa39bzTXz0iogLyIUMQqDlYPheGY0WXROVYQqy0JT6IoaA
25eBxXv6RTO7qTT6Za1uTPpgtk/KsBbgo2NQHsPA9B7Z4evtAqXrTVNeDU8lUvm7
9EnpdN2D40Z2JqrjgM1vMN3ixjaS6JEP2TJR33a8Mo6ELgFh5MHI7nesKiRS8Icl
8dURa3DI7YSKulnWkjmFazoycziRvCvZOKqRqv05fZ1vO++2HXtvWk3rbqqzfCXq
dn46skd5uGzNN0+5pIx9iRYJaRrxW7NURv0dGl/vk1de10S14mllbBYEh+FL+5xR
1M7+RReQffCIi6LF9qloZnq8UXXW6WYHA7LqRbnFRw9ZupD4QQbJxRMcgGH0HqRa
/HfKeqvff/n10o6yLx6OQ519OV3UgqpQNGeKYu21Ek6JYr1r+ZqYUGHJKH+5ZmXN
Yzq0tms61bENtHgZ5TcegSVdk6cNHj5+7SwJNhB0yFmbh3ky++CUAs8JsmdrL/D5
2hYXwgMcmehtKOqJ0mSfddIlXAbwnoViSqklAy9KBMj6swVTWqVVEXdxMTNxv6wz
e9v7sOEbe30V5z58viASLjvuLTtEZC2eEL16YYGduoBK4DgQupqg86voVXGWZYQl
6HWF0SwBJldgEqXJWTZhaq0zDgaxRVydlLRkjGGNfyVoGO57STBAdhas+qgbxLAJ
6lAlSIry7ZFgbLFa75z0rEmPNbTUt41Nb0VFXouqriznn8i/V1/AX6aXFLcvTKR3
bviYj0X24MHKaTX2gtUA0AQPODajiyBkGFSBX0lq3aROm53JyYmpDLhUzZJ/E7oQ
hKJIsZNSwHbIdj4X0oEkTLJ43FnhAYsUZM1z9Ej4KzlQcbnR5M+LIp/vVM5D9MkR
3ySTNhswgofVXrexMBx68miEx44Dgtcb71yYJIC7c3SA+R/HLpWdudqE2RkkkfIi
oSg58SQ/fGVuY2uHZDejaek/THV5Uh2FFxP6BAUjpYU0b1KGQCsfFSq2guyHTTGZ
OOKK/2w+CQkCezrcQcxR9oea1jXHKnWQkEBRgZi6uTAAONyKs83ybVVzNPOVE08d
RYjV7pLxZ17vlFm1Otok9I3eBUeDyl/N8h6ATmmerqHs+0FNqlbhNGNo/Avz1x6u
Y/OwPzGniRixiJxDDeIWNYCm8rtUL5dzHF9+iZYYl3VJrsMMvCYOIlNR9Z6IB3k3
zM7HlmciPzpJEilIBLk+6lye8Ii2K80/pFhWjtFkHWCDkBmNXbVJCH5cdl5sWOJN
CCRLamAtcxGY5PGfnhg1IgD736e9FKFWJB2l256rx6jbJQ72+FyN1+z63WOlp6V+
eKCWBkju/EqCP5NoF9SrmGK9XYLC/whhMNfDJlnD2rSza2enltZPKLE9AIJZNBQW
QUbcjdUvH9u7Fz0Xk9LvoJnP9FQXeaN5h5wDnrpP5n4zhnm9ioUKEJ6g0wmwaOVV
ztH7LxHd23wzlRGayZOYNC6sv+ab913bS+jUBLKOQuO3cO+gSbTVYbOtEVWc5qy3
WK/4f28WJXcYUYg+s5sqcz9OUxA0cgteTriCNrHaY9vJBbWqPFfi9ajVBprRmSIL
L//vHVBNxD8ubjZZ8KH4aD0m88ZTTMKzdAoDjary/hs2zZXJw465hh382vFYs9QR
s9OUhrjgjkG03t/KoGoxdxQPnpS+9kZlm2IxKl3y1bp0l5jLnb1l+4xdkfCBTIgs
/Fa0RPAmIf5aOopfXJRFl8IfN3RoVnxAHJ/qBx1+FH+2HIJ3fgujwZou48BFUEEf
2PlI80cFNxVplNltZknU+AA8YRYiF4XaRELpy7rX8M/tt384dM3j9ftTSWLVPezj
lqjXGdIyCfn51qPLDuJmvse6+7uWHDVTRPoCjQAzQQ+DkHALkill7QyfqMyjpBRH
9M65xw4zgKFG0h6gr4KtLN8YG31RJE+nYtG8n2/OkH4NujyC8ZbGpgx60GQhQZsx
pJ9zSiLfdFq2YjT3q0grs945qOIqbjgvAXwdkYnhxxg/e2nGa+ceQ/952CeX8xXq
wY8kyp4pF8u9olsffaWboh1pmTW3RVIJo1hLpj2U5a2iKp7anGHRJDj0B/QuDbza
thjX1a5J2kKjvuiNMTVrDyPbTJxbJg81fw1t9AwHLm6ZC+FTBKK6J1RPCtIn9Wtm
MBJxgC9kP0ZONA8fc+cn+z6aLQHZ7cQWLwIoRdwJsqrtsOnUqmaDUTuUmOwKziSm
d/BWX961SzlLvqhqGN1B2RPiegh3Ys9f5AJDewHyN/qAv0j0irR4RBc/2k98kNcZ
UillDbHtZQ6YfZZxSz/zzh+bjC11U8QtuE95r194NIDDj6o4lAJQl7mp+xqowf7D
NABBmynqbcNeBUvct3XrXtSj7XlGPZGuUmmR/OwPW9APErZ6qpbA6KRe6Lk/ayU3
eATkElaiGzS6cE15tH2gjHEwF/E68xfaHc57RJqM7cGws7L9DgRiF3y0kD0UYAiy
bt16mdAZoYhV6wWwKSMZ7UHdHvsB/TdevIYKI5aYhfFZK2qyBTijPIoxzHhvzClZ
2MTy2a3jSQdkaNrRiV2OisyvQSFDpiy/otgeRDgwX/jqIekjvRFm7YYmy+d0V29l
gJd+Zi5E3D2pefw5RXd20EYzRKQxPPfk/3lC9vy+hhJCvP9bvaH9J+nzxqFXdpm3
QWrKRudDl2O5XMtHg6wYpaEIgQtjzB1YAWxMviNVsJTKwcQfscOzwsbNE+aaSA23
elpTArXswUcYYbmW8JWWsT+T5zxMfgyH26wTCioIERPsYqhxaa4wGM8IqY3/094Q
5SEzHO0M83hh1IfRi2GnlvNrJ9IADWFfTv7tV7JzNSHtCetE/ZU+iysBH26B9jkO
lvOIo8kXid+zlzkDkDFij7TzGLgbiOuWP01OlCRq1yxp1tv/x91m8hPEsH/bLY3l
bgkKTHs0drBZAUj3vx2KLJCgyjXDliqOhbw6NgZ1Dmum7Spoef9GC49OuWgGPlO7
Opqg/mEaKIKRNT23ob3WK965cTWNWWzGvISmtMyYzyg/h+RtAM/yiNdS857/uX4B
bYjM82gJNFYMhzY0Nh6w06mcap4vMeXEgFUHiXQqYXfWxA6RzionVB8MGnsWkp+3
dg5mA5w2Xeqw75aiS4txFP1JZsha5sWGCyeLuubolFvOF0r0Anfr76Z2n3UMAf+Q
uZEw1nwXj+MC1ssqPtFNgwfJdIDfJxztqMbvGy20DQaUKv8m+AR+1hKIKugsON6L
KLduRb7J5mVObV//9wx1ojQl+o9t2UOmch71WJ39rBFPIfPp7fzx9Rb3Op2Bt+W7
AnsAHSuj54IB2hjwvJxGErWGJ/kdgFC+ynqDSUJVexW6MkCAh0DAx/oGC4BypgOb
qgaOTWJhiuMhJmhWPFmbaLsEJktVac7vtfvPfaobbMQM9WadOtJwmYJTgthkj0WU
71IZ2bHrsnQ3Z76cxnk6cpeCLTfcne0gDfmTjjOj62G4duszAyrYkCs2t7BzjL1H
Ju2nvyR/BW/rKzzHbge+SqYkhtQPIHMWXPKU1KDkoYKb5Fl4jwU9fbcyUD+t8i1s
CmeFzGB8UYgx41QLuA8D9CePHKBqPmT4UC6W1a9YDj+FKuJRlrUsgkpso3pTo+/I
EG9z+gxkQsAxaaIlRmCG3HKiDLPDemTcLkWEtdv2l9lTbLb9HWmEq9DOE9RC5iDS
bskKe71r7YGYL949sWyD91RrY+L+ys5Qm4CdD7dx57M5e9vX/BkqvYyqbA0FGli+
tJ1wPoX/TN7UO2tvBRcOa9sYw2OFHk4NzR9H6/T2wSej2QRGhViC1SiGHFZKJtet
cRdHSA79aje8iETKVyMytF/hroyP/9KS2KZ3YyQO/gIWyflJcVC98BBP7DS7WVAk
iWFFEB+/EnR7SIRiBD6wuxFNVFuMf1mFzMDp/NbvldislPut7eAb2j2bfBNff7qy
yr7TzghPGWFZZ3TwRt1sjiqj7p1MuUZhYHmJUaol9JesUPS7aaMWy/b66oWpA+I/
nGVXM1PvCCYYKW2ekDoTSg+qNFFajqewTZJ5VOe+zXhJEJ17spcBif0xShRm4A3H
GUHpuhc0VZmQ9vEC4KanZvG9oTVWCd3/feD2JM2Slywt13JENquf8MMVe8J+8nLB
tPG5uIf1nj20nkcgD7FLk7SxhopkhUro6O3NnJJqnoVZMkBfqS+2uxPC/QwZovnl
roPWrtyXwyd+xx9UnxBWigt7Y5HvNNcStbpOMx8Jx3cfQF0pPcN50MpSFnm2C/V5
c+pJMOOl8IX1Li4+LKHwayTcqHVz+6UdfzXEtesGelRGOSyUJPJMZOI+5C29o2iG
GsuZ54Gj0guvrJA9PjPuBGsXdE8/0OsDtQDlNbVveCYcBhU7enIdiuV+WQmK/YWu
n76Y79G3EVmB8fSt1gCVbm/VZpRameeuny8SpVQdbu95vQ+8KhYGOTlZOoO862ds
/KVf5i3HprruEdY4HhngmXssl/tvFKE58/mDcca5k8Qb6SJCh+hpU0ccqQlRDK/I
jusIdL0uMylZ3PrLpa9q8YQaz2Peg5DaWjoBn9PqGPuBUH0E0LwtZOdEZuSWZI38
VRz4sFhq1lZvZLRkTSAZsPlPmqEB8f0R06A64cW5SJued0LUUUl1JxQQkezyaIKJ
msxnO2NLs5dP5Wsl5RnW8Vo3QZUUNTze5ZiX3qbZpo8cfm7ZxM7PfgL9JI6TcnBr
kKqyVfcWT8VvFhfdL8AXn2tkqPs6Zwkxg1n6v+yhIQDLuJ8067B7j9YRuw4WXwGn
8QDUcyZ4FwUcjNRObXk47E9swrBXwsQ7eecKcsfvv1FpSuH8fDwnkgVfSeDdtgi0
0HhvgoBtcJ8YVaPfGVN4OIwdsojwwhbgv+ShMhoRcCvqFekNyHyp6S43tw6Bo6Ie
MJWA5HE+Z/xH+hpG7AEgUo/99TitQpUGd3f7teQKsqBqS/bEzpBUN6lPeLHFSN71
3ZHOiG57pJY3ZHnZAfVXplgw1XQUO2aKIP+q+fhqnNB1z8xRTS9cCiWWUhcNNJcJ
JGAUztyjqHPXcWzIYEny+3qJTxhBRJkbcPw00v7zINrcaH99Zn6VzLBXy2kL9hIx
0NCRMMrTqYMtTu5V395wLDys8QatJvYbeuml8MU5Ez1Zd9I39380G64oWF9ZLWl6
BxWTqVmOtlhzeFSqvaahQ+D3b4CWHVg5LV9CZhuDJu3ZbDBegq7MEpfPaaRK1o7w
35mJEXHt6Ct90Qeq0nwUoonrhwg3RhPUwTiSpHpUjBCoNXOLF3vobmdiEhF0Zorx
gbiT4cuOM3SQbRGjKsbJSzaj2WiOsXS4OuGruOUbInDHhKrvtVJplP0JO0AZentM
rRZVOzytBc496nQgygeSiiP8XlE2eiHdbHTkxlOPlWH/wvS8JLRDztsuPYM3pmKB
fzBVYUBtQL80wYZ+DqXDr2ilrSw0DM1JrYKBs9QmDsn2mICQ/sgAcNslrKTxVkyv
Fb1lE18qhsFVbljEnBktoKm9RguHs5x7qgwUGk3GcBH3msJNWJvmZb0LCC2020rl
O1qRWQZMA0gz1UawYYefQ2GQ7JelLb7DMKGLBf9+8scrMdiZqaa83nvRfJqmZNEG
zIc7HcL7lIdK/VgpR6O62p00ZBJD7WKIjqemN6QboqIj1BaaE48rN7nQunoZpF8W
gC8Txn5Qap8wgyLxvRoEXUrJ63nf9y/LdLnKmWWSVpR8tG0UH4TtxYysR59YPkvD
DqLu0JN7pv9PQpC3aIX6mw9BqOixaWMhny11St18Y2yzupLADu7qax62cycolZkF
DyM4abxOsCswErbY3r/veDf2EN9DgR3JrPeRIZ3JaiO1y4p3eHwMEkPbJX8WZS7R
FOmPys027bS/gqLpBfzr9F4i731Pe1ezZ1J5rHGuqEL264MYEAAXYvE4I5YTEEqI
Qt868TS2d2UwZKA48TxQl1pjjOxIXqbUr9HZitn7q87CB+WWeFpXSA6cq35o9qLR
jObAo67wSBGkFSgOIrGEoeVLv41MbHkB8HduokhqYQwQeGm71nsYjTUxT0N/IqE3
kCOuXqZOXaZ6nYvojLHmweuYDrV2Oco4IRog0UkQVzPd2cnu78O5cSHxAKKrzqrc
taDmRm/Nf1MdAV623n3YPkx04H39M/IajbirZyPh/dqi01pTdkiiMXG1g2GBo5QA
ru4VP7qVwfi8KXS1YneauQgQz8hlmP28mJvSXROWFktCQYSJQr+LKqqplHQUQHFz
epq4J6+R76n11Ic2CAn13ddLZ7z/EVje4lgSy8npEVOcudJt8nVuE9sjpv02KMfC
q62NYSmQRRuAp5NlOoYT4g1HjoTSBCxv5EKKSR7CJSZnuqOtuiJtJ4X6dWT5+BM/
vkXeDIDEHoW0s4ugehUm+xi0Ztr1yfecO4rZ/s3yPXz/hJGQIehJdYhCxHfsynOR
V3irOgYQhuSTsWROGN1bGFri46+jiQcqnxwrpI3bfB6t/WjJb9luYlSCci7latLG
8u/IeFnPeT5spkXiuImiui98N+qopKOzT2JQzRz4sDYu6MmykY3x3EJYldB+XFSm
A0cC+Y/JEeJCA6D0CKrbvo4yERl+NICYDv2+jM1zr7ZisRRAjapQC04/BYnSfbKZ
RIQHLaxkof/LGAZx1CgkkNZJYQ+qEyx82pRFzwiVvJJ+N4wlHCX4u3CT8Q+XJWdY
v7jc8UymG0F8Y785QA4CPv2+30bbEIf6rSdtBJmvlyVif9P4cwFy9++orZzopvDB
mQTs7kDjXf6gZNHDydOl/kk57LyaUTGhw0j6weW5FYJ4IiD0EhE13KJql7x0Zld7
Y7DJtdXBl9vCu+VMantKWgIbCa/W8DcyBOIASNn9bVB57eXrIEyB0CadePSz+HDp
9MDkOq1n1/6q5EFXEKcv0bInFpJThS8WGRQLyDc7P5tN28sC3DZtjv9DOXlo6pHm
RWEZakhVcsQFjvWq8xrpBFSBsOg7XrmEtkrG0RFfnSn5VBw/JJNd5QBpQFZNEXxV
+smGKShqPMCxbXg35y6NSpGTxRRxXRHRnyAGrLsFwltdgKdSGOyC9/QwmZAFLhZU
ujE2sEEBvhjYw6siw5bFgccUTx0EnHdpOY+dmibCEDTH1tCcbBRqywguuiFmpxg+
oDoTvb7RZrd3DYMxeiLl6eobXfZ1NurIhGiYf5/pe9SDU4NgTjx2+1RiR2m+DLls
nh6Yx0HnMJ9LnlLOiTKwgMYk4+DvDfg+pGTeGRkr4fKL4uMKP3dclo3uoMyliJt8
14VfdxtUaIfAVoK+AIDGFaEILpwOPxiTiQZxmKdORrmL0cysqjx1TpN/Z/fNKJUl
BJC3LZ2DMSF6V8/2lhlf52Fu5T2y/qvkel28iH5T4ItGxe4NriWLjQCpYr4z8ZOY
T+fw5sLD2EOUBYtXuIV/MEf16LQR4vBB/Pdkrw8vXELmssVfxbFhxMO2kXp6uqq5
61XKr4yOHUViGh0JxC8UhNubC+8y24A0ckj0IhrKvJzhYhe40Bz2xcj3jBB0IuK3
TSeEN/dE0OF7/7n74u06GHyagoHnCjvWV3NvITnyPBlVIhwY8O3vcvi5Rs0Xe50K
5AFlXit6VDQ+qIG2i9UOXUUa2uyTk8E23AaYugkTFzHnIiq2l/FnsDVAg7+YeGoO
+rgEBs/R58BwfsuFnsS3IyvIgowoZCkbHgQOmp6fPTcTT7Jqs+MG9GSkuHH/S7Oc
jUpNTFJdpiA2Ll0sJ/9PnM1suRC784b7eNR2RU5reUrwYnpruNCSDai8KEDBJMnd
DRD4i6kSGiIVARVKdHTsz04zS6EY0oKeNVw1+s4hdgajqbl0ODH933fSlWwyIYGz
5rHiyKhcSyuY/3+73Pxxo2atIo8T/332gyhVare3eeyyXmZLojsco9evAvVxOlq4
curQjQBvSdrWvQnr53cxjtN3pNiLVO0JErRGiei3zcMcKRoVQA12VBq6z1HlD2KC
A9OG06Yf+HiebnqW9vF9HsCnjsDQRbeyf90xVtD30qfn588NajezjNEih2p+vGWM
fMHRBelMhjAwceEtxW1EqP+B2Wvw257Xm9kgWfxdheArOzVXQyAb4L+NBzJLS74o
1XDf7bNpR4qfi86aBvfRO1QcGX5vscCnBvyW2NxMY25+XrYWNqHWnSAKeCLSiQoE
8vMGuBgjHzNMUVROL0QLHSfVj6isZsiK6nzaGtFfs8E6aUElhEt7NXPxE6Ixo+57
L78gVqYkhGwkw2ETB0ZqVnRU3Mq5EsDNR311hjjyUCwDjC1VpevFIN+cf8+lFIuy
iihgTyzw5hG0wY7lrDh3483bRE4e64c3f/5dBnjRcwCgG5MFVuyghqAZo4XhhaU3
0sRgZjNP+99Bv+jlMRyzFgwU26CFaXGVgffhadN2Ka4RR9j9i9mVaKahELaEEhbL
PmkITk8x/rX8I9uvxJeblBZpQfHels35qFRH96H4TMw9fFGeSreFHvAWAHwKmECY
Zp9vASY4lHs1TqtifnR9TVvhanbi4OxQA0qRV7nCcgdW3sCq7Qt1QZ0z7auwGRr4
KptC6St3paSvZldSqpT0vYDY7sgOZrTJ92ZjoW8li2somykgCoyvoDQq9TtwA88Z
BF97CUYvHwhVdbyR3s4G3z9P6LxiKgek4JbeLN4nh0zla/R/HK74dUKuT5O/sPGk
+kZEppGFs0BKmC++hWoCSsT7IcaSBJW6n0znZZocgm5yfzrIH1QwC/YjKgRiDLWi
wOzU+HVEBy4rLQHqkyAVQyEXNUVqVJG/OLFBpJlhObR4Ca9Qojkjiby3zpHqcqPH
bf14jxSOk3uSbKWf6P8FTPoHOxJfAseW6TEn9d/DWozTTXoC4cBAAE2baKq3e3Hi
Gcfbk8EHYi443lMmUXx1o4XpY/Uy0XbviyNAN6ynN9tgEbJUsz1s9sHgxF5lOlmQ
MGXT/oaXRceQ4o4GsuZz3n+txrImfgJu4b6qaU0TlaSAk+aKP3r/akK29O9KrQkc
6gFwMv+211FT9ektR2JX67croLj+PJ30iJ+RmS1MGfpHz6JSFQYfMZg3zqliMTnb
6Uv6HHFcZSMWlUl/kXH4zT5nyCr3HQjm5RYxRcLZEo7erPFJDjhmlR1+LPBvIY/+
DAAm/qGUxjQx8f9hYmqEtpErTORZ7YIuWoXSXztuB2uIB0c4YWmR/IHTL+ZaRN7f
FM7y5u32zSOBI8JarRIaVSXFM6agmhziYEzW9Gf+/VLy3CLCOKm8rAd8XoslpuWn
YqxqLt5PfIdZGbjdL8a6sLhfCW4kVz7ztNN+Le4400qslPpR6GtQMKwEVZFkq+o+
eEygjJFWSfpSColeEJdfBZa1NVqjHdo8JPg8Ywv/IIwXr2KM4qtz2R3Zb9k3gfd2
oqDKbPjiyTPSozuAqwiGIo5ui61wPcjfdd95iqAQRa+Pq/a7K9hcpQmvm1DHUCuJ
ae67uO6dDTWyudAyggPtFVycNvIwPkrEDJXXdYX52+aNAIrsV6KFn3I0cQwfp6Gd
o8dnX0cf0ESzKVOFiMs6M0WsmiHlxr7gKwaIWCj1X8NVFvbjEwb/UQAuhkm5W73H
pYMyH/08mfNzvFzNO60W91nlNw9AQa5jdcK6VhpUyFAuwB+hrxxuEQb511dBW2KE
EY1D+M1dh6zPR+PBB9XzLjGByTTo5kIGqg34jaBVRePze3fXTmOap9Ere/7ayykt
Wyx9KIL2JPHac4BJWSvxkN6H8WSDVDx4SdyHiIcFETtKDxIqTLMPSJisIe43+d9R
CIzyxZWOZto37EQnb68OI3Vx7W9VWZ7dlednbiv2OaQ=
`pragma protect end_protected
