// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:33:06 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
aA1xbAB0kQ6LxZo4EkGODB7Uah755cA/+Ca4RA0umZ58WegJ9gQ/h6UyZvmx5nm/
7PVbvSrf2lk6wfikgsOYZ2AqonBpeusaGsQRP0LJfUuOT4rx7+WIFbpV2jp1srfw
9+YRIxmeptHwJ4uOImfIq4PoKRMi+VDzXy9pqc4oXL4=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 28880)
E5G4Ox8Znb8zNTAKEYh+sQtVCcdUH6YHw5ilMRBqZx+jCF92eovJWstZp/aFuRVP
m322ZI8Mkz4KbbgCoTQ0B/KGdmg6tP3heqXAda2yNHPhvA7H9cbl0pT4GBQ30Z2I
Az92kauVPBnDiwBl9Qci0y5GxVb/KepkPdJg/LOvp+R5EHtbQG6m+589IlCRfWKR
bj5QV5p7WuOYdfxWK4Dn/+xPr8HhGprBj1RdT6RsivqskZ92gleB5pBFK+POILZ4
oWSUc2vpyXIrYQOmL+ete9bn1WOVh1KwphZXSp9/pPXEPpvOz2njvMuIU8Ee36nJ
Uk7ZEcEo5CelN1wUa467ze2l3xcGJ5z1hywTXG12zMGJ0PorV4vsgBzi6oEbMVMg
+FDeiJSLdBVznZhiRTA2eQglOksGV22J+ehzHYvqX9Gy8JPMgsb/Z0whGWLDrKL4
5HSdL7H+tB2/zm2XWH05MU+k1B+eM1UihboguieT6Qjb00qgZVFbpuqrgNG7zZBi
rcv7lS1eSZcKU5pL0RKsVCAb5RtR7msp54tXG7D3UWgnbTZFct0Snxdwyx9tV2OP
moWgneissOp7TLvlmRa4gITbYStGjU83kijV3mUBG2hxc9OYj2WXlULeb96jm59I
+zu+d3zRLtF2SD94xL3B75QFoBsFj01bKlOTIIF5tZ6V2OrvvwCYLds3k/ybf4kg
JF/XGdgGzfVZmrHEybQb0HxcGiGBD6XCLdzwRqY7i3ccjrirjyQTqPlLakFHx1dp
+gq0Mof9H9qdWk9t/iyfGrdRq2vhDGleJXPiGvKqdmZ4CLYEIYskIOzVVaIFs/P/
H++yePKxLbHL6tFBqpUdVCZ52PqCeOAEVLxivXEWf2sFpMkAxEXvYPNNmdocZquC
Vfm40jNNgSyLJqNiL+W87z1EhywmBIeV2Wwo7FNwzvnv/3SqBJPefKhIiKj0CYS7
0C4AWWVTNMp8kdc2wi5SwZh0o5YFSXhcMsrhppeT7gaaYk3JhTp9t5ns9wiNWGEc
qbxCiITV7BMYBBl0IXud4lqniyuW5v8xoosctBG8HvtELC+4SfhrNonFPW2Zzcc9
yZEjbAeUB399HHoI24BbnMHPfQt2YKzpTm3RgvArLR0+8joVMmrJW6DBOHzLCbDi
aL1lxX/oqojveekyhqjS13ixA4tyTr/NwLiW2ymIAxRvQzWtjIr8S2HG92b2BbGv
Z7DUalBGE/S6//5vy5gr9Vxw1Wmzz4z1p+YujjtIAmhEpBH1RHSimgKx6hqsaPgz
7Kb/AV4wDa09ImuIWtykdfNMsDw7+y854SMHaO28A2KOvsDKWhLQ7Q0YTCW/gEPm
G7yl7u5oFRfUez7RUbaauZ9HA2e6Iu0o5RnvWoEX3ti6KKRRmYfFhtjJt3waE06h
BP88gPA+x0yvERUfIYyIAkC/mdcIW3JUSS/4JBrxvV0G1xJZaFBDAJesilxO66jZ
q0G45whyRO23sbOtBU8W3lganpnJ5ROc+oiuBS+/IIa/nKQ7QlDgdcJ5s9mA/TtC
NqoiEfFKH674Z3fa3SAK1wAZbHJkQOOxSR2joFwTVbrjur5HMJ2Xw87GJdZcMJsT
yS4PBXwpBB1tJLcX8ZP+NJS7051MlY5kfNehQa/l7zH42F4bztpyZdRt66vhJKLb
QLxZUW1AR2fPoUC4/UBaORIFDEQ+8H4wTFkZCVDUHucPtSl7yMPG/XuM0hfCzV/a
GHyjiO2DGW2to89wf39FaXbQmkJFfSc93ENhkLgpsxco5e/Udem6EqCbBeyPvVEj
YMoBJSvh+MFjTD3U7myGqrS4VrjKNKPH2MdVXY8AgwylMolwMuxDvDHYhdqk5gWg
tZtwhM1vz6BuLbvk/rFz9owPe8z5z1fZH4IHjy18JpRz0ak7hjwRUdW3O1DZ04qt
wDN0q+bBBsXqJAlWEuFlzGhCsPN/UHDCV+6s8U4XSxTATzIFbMSrzYU1toO/fxVw
CtK/93/EwihU6r1Qf2FiyOnmzzJvy0Jrn+ExMvnRrRim6B8G7VtAOd3EDFyCOGMZ
eaUT3apWa4ENNYuhvqC+lm94oVMDMPuFI3NlL6Axxb2x6tnkVgZLotk4iWCO/ijh
P6oJHvFCKbk/NVJoXR23DeKakt6+fL39UXfW8dQDDp7QUI/awAsVc1emJ+IPV4e4
m9yuPT2qU2g5/W/03bLRSpuGfqq2I4t9e0uI43+yQBnK3ijn7L/m7z3wYNCP1myZ
FR7lcwLTl+kBPWzhQJakNM8LsClyOPNlAejuwUJ874qbakahaIz4bqXlTDZBATPi
CWUQAa71bsqCtjk3/9g71tN8CjdLTKcPSTX66GeqI348r4rAyRmBQNlMknlqmvpj
t9HwJ1qslKobftMENBMVunZl2/Ou5iJlQhQsJVHbd1IGnlTbmDky53gaFQ81M0AT
zrALKG+uEjp2+bzk6+BhIU+TnY4S5tlj5wQ2hcD1w2QJKzhzdS83zJYjm4TtkaZv
8SXticcwi+PZfLQNw9hubXdNsX/qK9M+HilFljN/dEDLgzNFyrCq3CQC/lA2Jgox
4dLSxp2A1R1ezJCxf/dAMUVaSRjiAc5s/QtZxgeHKOkvSsMyCJcvHi6UVMujMubm
UqDfxZuMkdqWedg3DtTRD96y4XdMOwLGOutAWtrsqp71SLWd8hN218UOjQuVSLbA
BJoTWPJ8N30JPG7mikG9Zdvagcz0tm/y9J1s2HoQ0qqJj9fLjDzE3FwRxS+o42ZG
izw3xrhqasaDIz+vnYsriEfcAIL7KX6uw/hLj2Vilgio9n+4lMcuzRePmI7TMO12
LHho0+vNwG4cm4e++5CrVz/QBhqu+ulUHlhlRX4qJoMAdVhFFbf0WfqLDU2hTIYe
H7it1AcrWF2UxLbkpgXzeXEn9hQSY4UMKzP1zOLfdCOTsXpu1yxyDTbaxUda3rfq
XsZH5OIAY3DMKULfW14TyWNnP65KHh/9QI37UoTBeFmEZwCO8iHdzjwQjQXod4m/
7MnfLnnWT547Umi3v7RvMhJDmIJwhG+BeFTVZT82qrf+vRf42vMkYc97InBDnIoi
D4e+2XziZLBDlsNwoqkAO7O1JM0zzhQzK+yg96FzVuAdlCt8oWPUQiaPAURYpYbZ
gLKx/YodDG2yzGWZzKfssdqxpyFJIH2MsJkqPXNm1KoEJfpKM6vQcaQ1uouCKpDx
q0p+9ErZic/+nfCXshSgvJi2o2AVUFdh/ZjiQ1DEod/tvPdQGwrmzxsvLvlqzlpa
bFJ0Xnxa0Pxq/DyXa+88CJrlZvbKHbkiipgGHJadDOYgoTPvHzcBnoMuPEDnD1ot
DHOLmDaVJuyuUFoURK/yEXOz6Buq1rGSK2ij907Lu4Prgi4GV338rXNgSfLGl2mY
81GScOZEqkK0FreOV8iZESSe5NHcAQ0rtE8qCiUMvq3zVPwxqEFNBHW3xFnq5l2v
zGHXUnI14NjIBSKkt1C+0vFekID4r63wgaXugelCJbGibuGJWsn3MVPp9WdpKxg4
KQV0u2y58OXbtDvqvJMjfTaiEUiwK7LfVpnNqI6lAHpsctf/0cQeP54VMMnP7nR4
6mpMIO/ZJj1e4IHyFpkzHxDsHU5YH0FpKxebIN0XF4PGZKNj3JUdvlWF6vq2dRob
yEoZVxcX5mFIXHBgJt3Tn/7SAXt0Q+e7X0GgHxvkt0hNErooM0GRuCL710x2Ao3O
J7eDhU0TiRaqlvqP0XM+5DLHT4BgLlaJqilk+cBOm/JlxjrKKOD/J0O+ngQIl/OV
N3/xVwIJKDBWeq3IzvjjDpcVP8cFZnr5/IOvVQCQTCUg/bF6+uhHPdI1s7XEynct
eTn+p3MflL7SSeCbWcO0REZzxQO5JlbGlKpyBhvuW6eafxOGG8HWdKkJl8EzAWhz
4G1GO6CdWCeNYuCAHIbNxOSnm4g/urnXkGSeGgVNewToV+Ultg0GF4fq3xoWlmfx
yMEiGicHPSm0FcDWpxG5CSJKmJt6PlGnPaKu2DLpfhrjIizVu80jhDyOJwJtkgss
HzM+oPAjBE8/zd3RpDXYRUOfwXVVNGYWAlMQffhCX+AT4SNjyLSm6mbszOsEubkr
Pr9Sq08LmvZ+e2TIm5kkixeuXBuyzw5eK0EW7jS5Jr6iiWMuohoupZ+zJoiNvp4S
91e7o2oPi0FhH413LqfHxqOrsqzQEhOzWzF24xO/7PHUDdUanqCGt4Z+8Lcw4ow3
V0flGzYosIx709azbEbfr5WrSAQYUOp2+OXFyDqkUkHauN+ad8ZQHBsslUQFLWk0
7B9syctecLwce0Ixiqgb6Co4qf6tAco9W25lV17oL0On5HGz5p6gljOq9zrwexX7
qyH6TgkV0wceycFJspz4pNbU5aMdcI6TTD1ODeg7G4eNJCunzzuo1sqCi5dvVbTF
ITKdq0MsF32Il8ntnuT8OFvbhxZKcj1csRrqERXT14XF1uHsVpDirvAkexcvp1zX
gvUX4uny4O91UOihBaKMQC/LhjD4MCGLE/aMkQEgiG3LGaHyYnuT3ybN/9gfKOOg
rnu9EbXN679TJ5daOZ2Bc9jPiCBhvBBMd1Dp41nqthLJ7tQoZbVQmrhTYNnZjcjr
h8MOMHVuOkfXhBZzfpdsxslBhWM+XQeuzIdOWwSqiHn5FmxixV68OeyNZipZQLgh
neWVLL0/C7vh1sKy8sG1PRqFBd92THnmYbEih/WrScTo46h6Mb49B3TZnBzH2UfA
8TCFnK8ueea6ELUvzZBwCEkMhFgmmjx3xmJRwSQIE0d/8wEBatSibjQBJdm/Uhoh
PNUZcZzjTe+fH++we885JFOZie29gYEQ2zPDFCW83PVb2wXDTKEEAUOqgsMCahGq
hza5yi3Kmb0MTa0vnqOzJC5vOVNBrVW8jGUBsYhfQqs4C+ytdNpVk+3ma8UbRr5P
q/P/9mZ0llLwURAlOXzoXZBVGQUaMZzJekeiJAFrdyKAlo7htNR7HJi/bNTGUG0L
B1oMT3x1FOfhUkjd7gI8S8TDlxOa6X7owYJc/5+wJP1SmLw++9LaNWp396Y2MXTp
z5D8MqtRmHAexkuMNyqqjFKptqdOx4GsT5IiZaEcOr3cDKvdRuBbzRyI9DdMEa3E
jPm+wLVJJr4qg5Vc2bh8s2706W/95iagfN0pHjooJ4JKUdp2llAxsY+tHulneTog
B/B9gYYtrR6iSGF5h0FpVJOslIYeFEgY4wqzM2rBpwDIH156lcHdp1KfWGextbfd
vDGWlHPNUMcR9f3I5RGTYrmza7+k7UJKbGCA5m8kcQ3T0ryzvvm7IpM8wJnh2V/G
RmIZlSiF5xnBX6wZ2VACSHMtqVW+qzgdgtw1khfFgd7ukkNX1xUysM8yFR43EHsv
zumWEvWgab+gFf0THxV4oohO46YND1Psx15jO8gBOFv/j4YeP7jcyCFbqAEM0CbJ
TFcVoIUCY+RDrv3ZxiN+weJbrWFzf9C3lgoNa4xpoftujHiNM1B+qokb33bmykv8
sOlW44rOfteuYaF7m8zNdKAJ2jqXoF31ovL/yN+Bq0qu0rHXe+b5KvdEN+5cBKBJ
q5mRbSvh+meHVozDiTFNRqPlcfGZlS4qaZt8S5dA/vvRUjt/TmbGY9nVIfn31OAx
ILkA9XI7pGyNMZgMaQ4XB6cJKI4VNl4+W9hRWJOU+mybhzETTj+K0MokcOF1ULeP
Hvjk9JDlO2Uv7lnC7F203CAFWx21vhUPYR/KOcSsczpwg3QcBR3/bpJzJ8WWlwzG
COl511o7mR1Xsn2x5R+tX7E3pNrGthYCgkbP8icFprWmYokwFrtEMhA1KRhV5HqB
0S94BjuySdc2rKGsIWw5xFpsTChcwfBw2Gn7WsZXy6/mlJn/x0gPKrMgpwL0Yn/N
9CESh1lu5tN0FApHfhKTCGRmEPyU2umasB73artCyf++vxOWh+cft1QoQJwfYI20
Xmv1zvCZ5SCHoSApTeLRMhjpycGkt+BToX36X/9vaHwVlkQQ7JFZFHnpsjquRFtR
7Eq9SjXz+F986xmdkbv/cH45/TNcWI81m+o4LkjtNierpcGE7DrdlTv3lshrSV0D
//vlf+7DN6z1obZE1A/IQf1JlexZLmfWbSO66EXXYppmVR1egH/zWNrFh9JEbnLS
v466Ycz52q2nCvKSogiQ5wKtvkTJA3EwLUIqHc3dEozu2nY9f4QcgGt1wl4uPCqb
PWt1/PQBzRqscDljFt7WEHpII3PRL8F/D664Q+8qMWruvwzbIGwa8p1P+1NhGYf8
jHw9lcB7Sc4Iq9Kd1b9zqFy0X79479upvFPnoW288p8ug54ubUvBh6KxIpDLN9jU
dhbATPWGiyvYyvzL/4aVoiINgJurRPH2uYArwgqvjBeqbsV9Z48jMROCQhcVkDdl
EBdEgcgSTe7knpJNrbOp4RCIBHqHZK3sWec8pibJRWmR5/yREsZBM+QNZqOaiek/
FjZkX5vbhRNLFrbNKQ1uWASaqf9s77MVNmJlnuwEUUomG4q/TcLV5Nr+xjchC/yN
tF7hpCbQ1XvqtAZAt/BcTv5RhaRyALNy1dUbu0MDoUA2BfGiM/rGxqL95O1Naxfb
jHZVBI+A+FH/YNvl1vYLIapS3TPqGStmFHLUWhLFPJzkIb35auh9sw7NKsr+T/zD
8S+SHKYv8uYiOMn1840xg4Z/Cdp63PaB0J4+iVVpidXV1fDCTYnRdltSTg+1E9wi
l5z2b2bMmQv3SYjGvC7YAcgAy25KXzhNP83rwRAXV91s3iiAj+/cusrzr0n+32ex
Bj95nEPT8kt7leyG0MLmSMmQIrOyU5oIt2h8akjtjtbZlT/KKBnMGKssijI5nop3
1Vel2ganPe5A48VtdfwDh9bar3bFyBW8XA0oCMoOGPq2a/dkTfm0yLa5ZjTh9k3l
7H2axBinosUPXo8Vl19Uumdu0Yx9pfAs80E6Qbjn1qU1Fw4E7vPumqR7Aa+AE7Jc
Yn2PuqigDRM1yaGvffgvcFpdWCef8gjc0G0hrL/o8Yj/yrXMrYPQleDdRs2GDWw6
ZkYXLudZ+alFgup0XTXu7hXp270eWiUnIlkZTYIFp9+9yL97e3uIveiafuIHu3RU
voMWWZkbdtnHq8ehw6RLMdwoSwwTfUiYZBHoyUirKpyFzNlFwdv6V9AImXm8eynL
3wny2X5J183adJS+hxBVLNFBMEORqhIJG7+bCaz46cs9q7hIrdE1xWrV32RY82Sv
RGPEjObQUDGl7DYwF0haEDlNaIJ/6nwGgxsC1OaPJEGg9UO6/C6GjH/NMQY2N5Bw
st7ThgT7C3MijjL26bpXrOgg6agqge9oWN2bXayqxf8KYDkCKwc9Leplj4Tvj6IG
xuDEpBA8sSENmhJNzKkVWtgYlHqC6rS2GpCFihGZNrz7yhVbw2IiSz3hFSa2MBa8
sKyNDcuBfmpQhM+5/EOI9uJESnQtuI90zwKkvnw6+G4QPziwevGUPoKylYuejtcz
lKXgMbGrbiM4d4sO64GAtg8Ko3p9r6/4PiRdTjwpTxF//70NZOv/APx7UfwsjbH6
TR4zOh6dle2RLs/1+NZuFzapFjV6cth/+mPFegvEug7IWhl+erlgv6pr5y8iaRYB
gES7EV2Hv9rH+zU7pvx4mqImvZVMs1q66tdtbXh32jV8CNORcrz0IeNdkULKEIK8
LOauUq8NRdtjARktlX9mAiZnDiQ7aVUbuJeYruSfpfJZBJpLyofd7o9Tu3qM1sJ0
9kW/5DRWkMbjLa3PE48rVbPMKNaFTKVk8WHXtmAHDD1rrJCUzRKJRjK5fjkE+dk+
9UIqHXMSQajTf+bxKvqVUN8I4bX4Ym6GCLLBTRXcWUkqnHnMI259Co8CLSsJk79+
9O9NIpNQRZ/EwJ/YLmuAYAA9ljWt84YtAHMlD9mqIqXmc/JlmBA+mfTe+24SND98
x9AZzwTk2JyrEXLwBAcpTLzcLsBlvi45yLvAN+0YTL1ZeQez/4J/47mmzwnidhof
tlnCFpSZBlxmZkVfV9oxGNn0C9Adsv/5NjKZc6re3FdFj0kUPi3bPVabaOpyQ8tB
FNUQBcY7dNLNkH9I4Bv/UpraUIK3i1UW1dmcyhJYTeEfDtqDI7dgNlRSKpjyKIbl
yQk92m/CCprPoy+yk1kPHKruBK7XNm6ls5VlQs5hi+gJEugdL+NxfcvToXDwszwb
1DPhhgRfeOd3G+Wl22jSp/J+3pFaS1wz42CNbCzhMuwFUDy+Juz/2QPatLtKJdKh
utZzKevyp6o0D618eW9bed5xxjSYgrtdwotDVBx/n0dJ7ygOp3CBh2PNFaBsFtcf
d7jrNbk4d2s9QQgaYWqHQgqVF0cFW5Ox6O4+WytsWJXDWuJYJh/CiOeL96SA2Nbw
NO6uwZW2Ym4tmhTU08LTpNCTHedJ2kSPeBuzC/tcE2xfq+pFLNv9PjyRITg7bJUo
HV4q2oe+pmU11oxvMhFrCnXUZLJO7zTVimwRYQyBOn4ZmLqsbQYXJKUd6wg34ZAJ
v28afQJ3Vbkjry5GRcgtgrX7O89Xm2qi6jQf3+uDkUYDVJ/rCZBO1zguaDSvAn9n
I13G6RJbjGmxaxAIJPE/SRyu8Ti2mW4cTQ7XSV8gxyjDLR5n1i9xbliyqn2JXXBr
Z6svaO8oxLcJRCRzl+5BmyHKtHl48sVFc61ZT/Xe6d8vytl6d1BzARVRilQTXotB
3vA/94ZrknQ+Hb5DWv1f3eiDjcusN4FmLFNFEuYYRlmE051RxWUcl+4+t0lEqwsM
jp93zEh2G9L32s9+Y5jFWoMlmb9xe73AUt6es8CWFfMri+7yrc8s8Bd+oeA4zHpc
K8IKvdlEIfrK4o/NxJmlAVqBPfZ5/E9ohFTqkYjeL5dh9j3VxaabNHsevr3I/R9w
dtPtpdp/PyhyaHpnO4KIF/qjv7mcxwodwYyrEQnl+Pw47C3FaHIJnuvkqDPsJX3n
4CpAcNeetriPSocevn3pyX6SS+t5w+Voy6UsPqmg3XF0IpdqSyRVMpvVzJAuEUVM
dHhOUgHorQc62c3L04QjY0B28xDC0Qaef2ti1YBlh3vwdsXVAHloJwSbfpfIRjd5
6feYd1JXkIAl0E5Uw5XMEsC9KIVejtn+NnoBgKOtboA61NAIHpqP+9F279pTXKyh
rD/UY8yyoNKZMTddl6UUatG/8qRfGakp3ZbPymKszfCtDSD8HxEubreIv42Xq7xs
Chg+ISEqX8pcD1BoiqqvznLWFfzm3CrGIvEZQPFrqEyJawxOhodtiN+cM0Y0ZBI9
hTGyEu0Tjw8n1rJIjK5PVAe5Il4rSZB/e9N9UqxKi8wqLMQk3Qa9S//KL50Nbevl
+a4ajU61H1bx8d/MujiHO60Cf264gRBI9zbIqI9JfprMfACcIi+wChF6CSn+lZ4J
auesbu5sDblaCD5ED01lZ5fRkDG1d9h2wVIzu4WvF2rhI+VF6D1gdOtuelUI2MJc
mv4zUvE/MUMcj4IDzz5AcTuwyDws0ZZGAkkaO4WO7+a8af0unoKWk6tKmckXrL3p
6wvmPRgSOXjXYZHIFqq1ZayidEbsmkkEpFZY2pUgrZgz59BclUTnpEdvEUpjI4Ou
3IownMVEK++gfFhVuaX4LKovMLH8uNKm+RM/r+yAYrA0AjONkq/TD5LfzCZNBHNh
BvEKMz8BIibmfyNftjp1Hcks6wQQPSezXfaHlttfdsHzUI5XsP5SyOFzF9KcHMa6
HXloQFEa/Ni4542xF7fThenkZ1HPml5DT17RYcOevxpNjPRDzbVGTAwDtVOMq4rX
TtC7OKgt8DIFFIHCxiVq23CYS5MUheQlr4ZMv4l3fRMkJibT/j03IsXjO+VoenVR
GlvRvGfW3lKYHbHgwkYK6ahYRU67n6DjE+FZeeRyd664Rx5aK3l4K6aMnVEhVafN
tifAdmWSxi+ioflOEBFoKW13+NJiSSlTWrI/d+d44MACisZBK++7nwhWphys/NOq
GHHJUYg2uO+6r9j2HR7S9imGxIKqmK27r36H7A5jUO4QCk8JaB8BJNhVonvuLJEw
61UgdwRN/87jh7BnHRlpwuFnzZjDzEMD8gCQSJfGh1KDVlxGfV2So8u5H08qNUml
+AyVMJ5bL1RGp5lusMaqvCFHU+iuSqY9A5lyaFpiLcpQTw+VqnygmqkUkeNa2c/J
ODftHYs6kYNV8JUTYBEKTiGdek/7vSptddKsNZAfKJ9zXaPfq+JQxS3Khf5r7Eel
L7OKZolqe12aFotnQKUwVl7jOfm7gQZz8omSOJA4PsDdff2V3AgW9mrbvmQ2yP4w
EvTiNdJ9XOjJbMT1FF6spcJsl4z5uqtDLzOWs/Z8lbZuzGQ1XBYOr6dVrQ3nkIxd
5pBayT0smtzn0wjFu40ghf1SPHKgLmETNPJ1Uqo7BVpVeaIzrEtaMt1bef1Uyh+C
+YzJukR8EYvnj+si58i5X12sYFqW3IV10acQVRf9dN21rF76EZ9oobPyM+47Oy56
cAPE6l0tmREAKdI2NGJKBaBHk9Kp3cXS4h/vaoJQi6cZFUaLav5TW6v2n+jOrNxG
Xgm4yrZrFJTwCDe3RBqu82JL1j4Ov0/y/ozn92bzrpCMeNSu4oxGeHYkeHEVcVHU
n1AjKk7Iv0/NRObj3YwNZhcBenu/95M60/5+/8pnxGnQRfOZjteD21HcVBYm3nuZ
VPPmoOjZk+GqgpjbcKgkJw63PAvvk19U1Ru4vItYirzNNMuh9A3MHElnu1r4de7z
sJa7cB++AdM/WDDHC1I4TprPSc+5RjFtahG63TlOEYPao/rVTYSJ2sZk6QQSQvMm
twkF0prOman5AZp9jLCk5jZ1RxC49oU6OUBvwm3dKuNHSzvqDszpYiLLK5sa5TkO
tFVq3g2CmFE2eH6lThm0lEyqLrEPOATBIpp1afZlutY7SGHG6GiOpk9APLCJ5Tnf
wq6DOKNkoVJJgZSUG5sgEdgG4qyoQbb6jSUNVpq+sRSkFEvcZ1ymLi0/eZvGSEUJ
IvEJg8suMcQ8aa4/kRZO5drcKF51n4DYCqzu0DraX0P17rjlyjZxOq6fXW2/j3rh
Hhjij6Q2sxaQYXp9Mu3Af4LXJvXxCxz2UrIICmjULRm50SGa2bqort4gsnsgJwRw
x71mn+41c/chIc8f5bnaS8EwH2aaZGJREN3ecMCRMtfzNqo0jIZZv69bzdArQGTq
/J47CgHwYGOX4oFEMRe8cXHsOHPKl+acHjxw2z/TEuhzVxIvYwHw/trkjleQ9jD6
aMvid7F4EghFqUuzmSmwyq9vesO2/F2w/Y1EvrmJpaupMzrtHPMo6d0FoyJVHdmG
2s+u7kRujYn+VDwiHso7iGUtMxwWOH3zfNf8UAGIu+hnJY3hNFwNR1LWL3Yorzig
0pAu+sXKFji1d52nQ5XbymrYAeDDnUiKdqolXY+Db8MURBH3wtQPHej8yh+aT26p
1SCZMTSoY4yrbSw1WeUpuVY4esgIf4pBjCvy5iPBBoSB9uN6kUhAvoeqWDTDQi6i
vHHpELRTTlmtsOIJnUxwHa/p/78+UVnuDGD0t5/rIudPMR/EwsUjKLDUbwbRwlIO
PYtX+1WA7MoT+xa1hOP8DkqNl33wpVvvvpR17S35WUBra7Kebzqwz9j5ZS1j/+Sa
9eP9mrNHmwapNMxg/oX+yBs01jv0kAS5B4y9WAhjJFIx8AODLuzzGVHNph4g2TcB
E/WgfzMMnnw/9HPo6kXwSeuRcgQSoK8NmJ8HN0eqZRamyGKkmUowX0EV9SyWqrFo
d9jHP5LaGWUusm8XpWnbDtrMAi02YKSaErWZQ7pENgc+Q42alshLse8eZVr74usY
ELoF0npm1f5HEQoFm+q+PnimgUu/nNmOciBjj8R91gEyUTo3N6d0f1TQ6L7w0QIh
dbmp/1th7YBLq9yFPJ3VqBe18XFNCsx0AGlsZoC0CZlb6bQoAaPekkFDCULKvW+z
Djgvky19A18F08hDuh5HpqfNXZ3w5wHaQjSUPMkqsb02ErU+U12bFXryneSN867F
ALFmVGdKnLYSGXJNs9fNNDOxF4V+/cVEp8YXt2XRVNdlc7ohKKrHQmgNTrwbDgtS
P4OXX8eLOT98fDoN2W6Nk9aVF8IVWyViXrlOFTxns21pWdqOS6+w1DJ+LzybY+XI
uXGjHLLVNVaVO09eFEWCpwJVlD3CfyeCMN+l4WFpqhsjCw1GwyECF+3QfNvczxPM
SmSwHeoaypHPPFSq2FkOSQnjfd/BPJKCjw2r5EGHpEKq4JCYRyZ9O0/7QBbuPANd
SmiLzn0YFw5QE9FIdlxPJgtH3JdeCsIPC1Jf+6FvqfKgqGMe8FRcTPaezyXbKaxt
O19LPc8ZyW+CDm2PcFKK5Qu6Ypme7e6I92mi4FZbQglDc13sMtc0rIXucX7AcBwT
54JDUkvvJJxfdSgSEaBbUGghBr2o8crSbTzic9c9RL/PUSXsd2SgFW83e/kI63O2
QCx3CS3iQMDW4SK5qKOCaeNRLzgix8LzwgXx63rsDvjfEJt67LO3XmR7/U75UUjK
OcxaahXrQlH5TgwjpJOAMybFFw+HRVQS/gcCRkg04mV2TF5ak+PWn0DpTjSAtlZl
pIOmf1Wy/i0ODGgEsoYq6PVKafr6c6SEeotGW64YPu+ZwOwl4drN0WxGvKVb8PK1
y46psKOfwkc5AS/5pfUPMmXR/k0DDBhGNz+sS1bNYSilC7RHi7UJ6O8JLrka3rdg
jYfNipyyyWgVAxh3fx8by/b1l4jI5n8AY8eHpf7xM0mqxsDwd/Oee1hVhGHh5lh8
7sHpneFHz0G4NWmZzN0fNuwmtYwi9YBB3U/7Lzte442eF7t2BZNK07DHg5ZHhyo4
HgLGGmcuIQwgL1slbp1sDbsngCsDANH5FOb3JxUNCDD2A/cgua8HMgn6JQfIdVnB
VJFOly+Z1bvMVYOmaa634kNVsDLQzGUeHQpDd+cdJMHgsq+WGYabuVsrhV9YGGEF
ztBZN+fXFzNRFz7iwf81Zi8BcgLgy8JxCxrGJMUxk4BpZA9ZRNVbD6kelQBgx2ls
dqP66YTQk+JiNO9G527mjtlKYqYm+Lozh5uivaPqqFSzJ5jJ8wOfKJcU8TYkGP0I
pRzTImNlFjdg2cWYSTcy4KqqmenahSX5ceOoO9Rqfmny5W+ads7w5VWwsv7VCz8e
zTpClF0SRFmDhA92thTY/SnXEukbObSW15mNPojmQEmWNn0CMb2+s5tYdgYeWzJJ
ii6ImVBcTI2uMP5NAVPfNeQjacW6qzXc3bkF+/tbfTXtE2hdKlSNgplV1NL2ie2m
hpkhWLy8mHhpoL6UxlbiDEMg9a2RmdnecVabJgZSWHXNsWRwXrWelQg283mXhj4o
X804aFCDeascoIyXiGplkb8VSHkQ89Y1F2taWGRri9ylbnmLO3s7fFvQ/xlhh7ux
IrLP4FCZuqjzr0ND5Wxi9fZS3B4CkMyYjkor57fP3fgDqiS+EbwaGujR9lV8PFps
/qEIWe9Zi1LWSV0Aw/QhrTA3vFf4s5f+XJx0yz+tM3XHTnpQJbBqvaSQwdRBCQ+k
v3iKMJsmudWMA2/HiucEDEHJofGP+aqNM9aiB08onaqnaLeaHeE5jMgqWkYSlQVS
gqO0U1KMQWaqAIKZkcKMg+9xsR0G/nlE8Pi2+PkmWo1cWVe54L2IRyTytDoggUHP
wbQYONW1wvcJyhqtwVX8FTrvgDZz8Hj5K/+n0RL0e1eHnO0+c5opK8/fqG8iht80
geaR/TAU+vzsSNN3/clHSbwWv8ITqKeZLA79C03v3vzkl+Gzanz20GNbadxXdMD2
fbJLdvDbJpPf5o9wH/gqegmE7nKAXmzcHavq1l/reRTCeqFqe1Opg1ICL1/gGY1C
kiA/be9BW8kIysR8T2ezFIDF9z4lkbxCFUxE6cf+pGpmkFQ2f177QCWkM421L+t8
CA5MaNF2K/H6VDw5YwoKW3Q+APulAzZMe+vG69aOxGkcExs58G0l6iba2VEZISkK
vSPnK/YWScAne2cCEzykEaxZLPOnzPJj2I1i2wfnqfJMs9uS/7tkSHusiD/Op7qe
/tk2kLHU9XDK/gBR8Y9BL80S4pXsWamHavwyylyn9sq/fdP67r9G33Y5q+k/BlhV
j6yoVhdgeQk+zOUduN9ZqWMkgNrQw23Db7h8QgFoJ65TfcirGW2BFFzx19C6vP8m
zoX5+zUh0RbtEjlt4mfPk7yPzhqJ1fqMvgphiN7VZetgGZ00dY9c5lrX1mS38kbY
E3AbiKmSSbSdOg2GQQSrfa9Xn0LgZSKrYoHt+nUO1c0FBe1JbhC0Bc+Ubo5/XAwz
AlgwX9fWegMLoeg+et2BQMKU8hdinLbG32SZt+mysZSLz0K7Dy9+ZJaUQ7MPiT1Y
7IBN48YQ2Z2uXNqWi6NgY9l7HuDWl2vEEK0NEEiZ8xP/+e4xLUhVL5AAfSafSXTU
hw/Nf4HJL1tTLFEvUQf6CwnoJSfT/2xLNj0XJzx/peuUj1b3+FKH6ADiMFVrpuBH
9Gdeom9XkCRjwPP0XT4spSrCeKhiEHIHpYIx4FbEJ4BusMlJMApbwP6bT38B0mXN
akMSE0hIzZn0A/pNp2IrnX44/oJme4Hz+pQE60mEnFLkuIpiumNbxmZ8qD7INpss
RpOsKsxSNYxItZON7f3VgHz+H3pqAYINkj+mhpv4/XZ/QmVDQUWXEogTw1Z49gOo
5lnBtiEcimUNNqfX2oCGc7t0QIGxIZ9qfW51H910JH7gXIg3pkg2AiwpydVAeQ5U
kw+ZlMqYKCP8qT5n5dteAMMO+ljEd8ZgLmg66MmmPpuObppJsGpZ94Ja0hTrjyVX
L7t1DKRM+Pq/Hqlf+WWp/6qpi1773Z9jFb4TF26/fPAUZNMUJQotpAyDttCedCUp
uuN4Et/WqN3lkkrLsNBWvjMD221f3Eh7fWYvTni6BWs4LHQi0MvnmaQVVP8ylruJ
O/5MsC0nYGDTfgXBdsqLhxj8Z0eC+Qr3/iwjR+r2iHYqcXXxircQwnpAGEHFKdav
S6BQiOjjr4+XoBkfgoN1ENmCWpGjXkCgZFp73EK/iZYkA928T0mIijjt5jOd/lbX
EumiWu/bqUc9wuNM8Gbjls2cPlsZDxvHXqtkLA9XSUBSDilm6d4bhxZQXqdQSGig
VPsFQVnDIVaI/iktAMR31Z92MDYRXGlOhNpDhX6emx6TxNBQtnIiAacZvNKVvzt5
55Cg3OdalT77eRWTO/h6DjVJF5Es3wKs63H8dyueQRAV7vkuNEgQ4XBh1K6Q08AQ
Uq1cruISN7AYBhYQU/yPJa6nECSkPJAVQvXeyREFi4fxBTs/tLNqJZqowC5CrfaZ
0ldK5AMpDhPunTxX1S2mhsdE0CYwYbhlKdR7lJwJ2CA/Eua3LBT/ZRY+tpJiCsbC
EXJwTG8SlaOHhFPFDSXqSclUDvE6KdCt4/kOwBhIbhGKGdKyd0bPeSeWy/FZwqMf
nyqooQ3KfjmktbK/Touj4ztKX73bFZys0AQ+b8WD1MMQiENsrjss8hUeTPW14Jqa
F2LlT9mitk3mL3b6NDr+dwhAk4hp+FbARuBzOg5KI8J3sSSomGO1uA4B9e5aCMQ5
PK/eQwwXIXv76fo2KHIxeb9RlIIokJ+wh3uyLiF96IUgxisdFVlNBGTz809jkDE/
snOyIfVTdgMW7elnmDILZ1DcOeNTHWL/Co6c3Z5TOcubcIgaa/jQXESXO++A8LBu
+0IEcQpqDO+cgmZaga02YZlmTGD43g0lr1/OHQACvT0S1Vxd7bi3EIuOcvwxOrKx
1xu7JvgjFJd752i1T8+rDq5kX88ax8GNOtxj8L65J6UaRMkCe+fc5FUlMevf8Mnq
T6WAJE5vgWOmh4ePsA0VU2m/qKcqZvhElPb2cJ21fllgaO7JTsGL/BAkUi1Toyya
/oGJ9qxj55bZpN9KPXmtZsjRx8p6TtNyalLOlMkKZl3mvWQFUw+TyEkSwbc+cTbI
qdmytDQ6Hg+gFehnRLrUa6fDOdUels9uCReReodSew+PHOczPDquc4h6GLVJR71e
HSTBK60N8gAtbRx02W4xlWTsk7hZ0QWQIDpJf3Tab9cU8wPYpP5u/uQwVVupE+rF
b0imp4A/xl7YqUgMv9k2irp1Co8G2WM/e33MwKHXs2JygRNWMBX1L4ToHWlT59qY
1tZKJ0nMV+hvjQrWAR7kUb4fwbC/nnmPkHr+CdAEjmCgVs44Xz/gkECLLhgUhXsS
Fek+mqXe2kaN4MKzidW6gK9gRjrpmrLI+vPkMLftlLOkYkXQv3o12rGhX7sLtD/J
n4DnCPuJyWEVhfgFM1zhknPpTzzNCl+4S+eD8pLp0jbwySOy03pA4+biqhrfzdNc
QNpz1kPjuKBU3A/wZ4+SSio6hj/GUO+C9I2aPiwjoWuNM2P2h4VU89g4uAL29atO
E3yFTHdQc1f1GId8Pef+MK6Ma0Ot3Rj8EWvoO2w1O/tTUi5KX4bDRGeHGK40eUxn
UemCF4/Mi9BCFkWL+KWsA9bSs/XYRJqdNnQa33BTz9YAnPEHWrZ3xvbKq9Ok3N0n
mUBwSwaybKjXC5KLTMGhjkLqy7U8JNV/74y92XNHHE6Nv1m5SoPe4h0GH3TLjiol
MEZH/TUWAfo3WHsv3GRc4ZFt716BZprvlU0wNJRaM7U/t/8xGXRA3SquqVhx9rxM
OQsq6ETVC9idE+D37prxN7oLXFmsA/nlpGepk5BPh2BXoZCAJAWyVtdcGTUSNjUC
I2tjifUkrmuOzY4e3aIANTm35P+KZqM+mDTL2d1ELFxb6O6V2duoNkaYjbPgTZHi
JBJb1M7tVo2ynI8CwyemWzMC8eKSqmkeYAtb2ApGBPyCZjskpLYdAHPt2BKxoR34
ugtdQpCTFSaC8WnS/ngr8imIbJeO703KTCmQ9y4mm0qYU67qo494eyiVN9IdXBZv
SbikjD4MczyMoxJCY2YQvmvccbA1MLSiOwQYFVEBuSq8bCb8wrlI+ej/9Wz0cVaZ
MNXbsv69Y8BI2pPrpIdsIXu5wnCst05+5w+2aaAmM00spsx1JD+O66r15og2Iujd
KWB0xdcJR2BSh7JlAKYpFcRwaumt6dr/jEjs7VW9GArEkmA7VmVcaATGyKjs5dcd
ZWzdgyIMJKUb3rwb84Mte2nvieRPJbbMTOA/OiW42Ga7C7ZZEm2gcSjR3CNHyB7H
MSER/RcQQGNtDvpxEWlDvFORzv7hYX6OE5yshJLAWBe+77DYHqWN2FDiEBa2QVtl
/2kabIIo9BbYQDwSBk+lEZvytxTHFjJGXZlZVi3w8GCnqXZnZEgibWuOkdTI7PnD
sXTLkJjAQZ/TdL7tLSC2Ah5pXIgWaUP208KnGogIh7PY/hAZ6mAcGRNoTOl5BnR0
zltVeI2hqpjnEvTNJONfW7RdtEkXMjQikQ3fA2DYEZpA6JvOuYSUTnd71ngos/xg
182wF94HIa+vAYIbX8Z6qjxx9J2oENcCbiCKc3ToC3xHBIXOPNVmovzWRySnkBqu
Kit8fljZ6IPTh6hULRomwlkMdDrOoYCS+0HaNM71ncCn9p0Sr3evbV0bIA+4v6Md
Wp/X/hXzcycqi2n0PZWYqCCyzqMOcE37LYkt6SvJ4F0DiNfeIU3nIwJ/NCAE0I6v
tgJY36XTHh7e9L16BxAPVew8Rxpdnm+VRLmuUx41/HGSNkZGbdr4EmYB6vuFTIHB
XUa2/+q59083rykplxc5f3JG3BmAY32shDCSDhf//CjZ1tqtsqivf4m5pGo7CXhv
jpB64k3Tyw70CpipsW62ZCYQ4N9tzaWwVSezSc18eA8mbyiFmLd7KhOlp4MZ8Nrp
yBaERZtnw4qfVdYQ8+mPbVN8vHV4sM3ZCYAPF0zs+chCGMde+hyU7jpXG6fHUoDU
fz2OTHnXqdYrlUxaBJVJCA/W/n0TAUmkGRwJBpe83yEcJUKDRrE9YEZMKxTIOLoD
alNgA3B6nC/Lhqg+Nt4KVzpqM5bam/ZFt/JLkzCHGSrSquYX0vMQXok0Y6S20BzQ
YepI9/i1yH+3fje4vG4irQ6BjvFvUzGGvEiXaWG9jI4f6Mul2KM6ZiX6WVnFRodc
geYUwNX3mSI6Qabgtri4Do++chqaBeLbf1X3EzNQ2EcKkB962U3Lrn3NJ3K9U51P
+FXObEuTYdBA3jLSLcvYdu3tf7/5FtKJqkIx8TYaTrPYQ+v6H2yTJDTotzR7Yh86
MHCCP+TzcR+G3/ZQ+eZIMvbl5ihvanbRZvM+tF5cDGR4aEIYKrmLNjiVH2uWlRwu
v2nykldPevGAsn/y+JffHsLISUxcJrNh+iCFA/vaSAD5pbGQyDWo4gZ/eUtn6J8C
VuPcEVQ/aqVN+pAf1VKIl134HFAH4uRxiL7E7rICm3BT3fyoBFih9H2n8vOzT9bj
EKhy1pvAebFKmAE3lNPLiVGsdjcYor0wIz+IaQokiPmZ2lvzBi59fgtUa7CJtVw1
RSOJxct+o8vxkisyGA+OX3lz+fj8P//r31YiQtIDfOpzb11ptuNCmT+kH/VXea6P
pKXj4uwEmJ2uOOsvj5/bcIEUIgdf8klFQtLRhMeUy2BVvEfYp4OrAE4RJejYOkoR
1TeF2vzh99G9rYNuWvGeoOHOzzb1b6f6HgaGVR3EV/5hHRVGSflhq6Sy9/JTtTKs
WfEj8nghvOvIwlymnJL3aHYBLD0Vz0gW69yseBxfAumjdVEdNE6W3pSGKgkTa729
QFmoGQCcdIyiT82GBd6mGrS9B7rN/Kb3xzzTkRZqtnHrxS7KxcYU654U5BVwdtp3
y9QQ+GrurI8TyY9T+QnTAGL79iADPpZIsxTYaylHtBJkx2wKHoeK19ilNFZDk6+A
aEki20DXfB91hEX7D+oPmJ4wPiHzIR87vEN3Qy8ablB5Z9wEhkK0IjwFrcUKmito
9+fjgLypS/y0mpgh1Hn1a0W531cJB0GLvALf3CqbAKLgKRwXXDSMUtfVR9PMTQ1w
+xFHIichPRmv8GgUc+uUQJ6VOrPAPnu6kzk0SPDlp82btqLc/8riw6Xp22yRHJfB
8po9JT+KrZ0YgYY+vKtSHj6j+taYjD0j2Dh5x9qi46mJS6uO0d87Qw3ZpYW91NjE
bEFIqxVTdzmm9JItXIDnIV7lnEQysWOjCnY8o5NLmO9T8RJznYndkCo4kEibCSkF
7g2DsRuJ3UPWIyr+i9qqhaq1bpF5mZ1P430LcfvvjIOGmKqJYcHE5iGAem7no/qk
GGjuDIKf5O3Gld7m5kmCw/2ciJA/1VNQcoNKoxQ7sr+67oPRjit1r6EU/PpMNlJ3
QqnfXHzqeFaYWWVQGMriFco1JEiE8nMF+rcLLphjj9uwfrwaqz/KBRaWIRa72coD
9Auw2+pZ6Cp7swPJbQ8tKiEUCo+NkMkPk4CIn0YYG3QJVkdMiwBDjPwDmjhSetxm
GIXCjvGpeJaxAxBB5e/rTEa8A1nWWMmxGXKdebktVyzpPCEanprT5MMjK0glTcIq
ODIan0tzcXOQe7zoY+cU0sj+HSkV1LieI5hOhyRAiASs/ejxuKUKxyb64jHIHzAO
lT9M7s5t3QJYFqlEQbQ8fCBeiZu/g29leFKZmotsnVp4Tr+kajYtXbpHiJQC8fQi
IbOrqU39cOhvImSti3N1zSWxtMpNVf4km3Y7LSzwr28uKjGr+rLGhsfygKB/6Mv3
4WZG5qYhY3HpBpY1JWXZzLndFLs+LW6hcja17Oqis/fScRmyNplweIlAfMu2qbnN
4ce78WI5o0K4GSveFFeHF+eem/4w4Mf7ghJ5yhz+2tO8yGlgouAh7MR2LFZ1OoBZ
w7M3OIygrQf2GTHIB6vtuL+yqstzEEzMS1PXz6+A1HO5VelJBC3qy4/nx6IrnKPK
vQMAFRlsx9dAuo2r9dXxqSBpKTEhiq2CDB2mdZpw1W06q52zD5sn9Wj0H5UEFv0X
FoFiUn035Chd/D4rdWcXm3T/CNZvpbK8bVhvbap2RauC6qEQ1bC/8/TQtlgFC4me
QX+05/qFr5MsehfdD3w7LXglLE5y634jVLdvhoFWeo7kvY49Q59yYUgEFztKX/vk
tzpm5/2fN3kaBRgK8SDYj/rr/H15blNiZwZavKanIrcCOKV4wTOcsoahthdtMXNf
FMy7zRXrVRtw9ILSLVAcEwOaigM2i/Jf/YDkvBEHvf6/CXuuIPHZqGhh4Q77rn4r
hbSTr7P4La8/0Ea42dpb4NNO3iN4a7ObS3/iGaxKoYSI5uukjA4EeymdHbo9t3Zk
4Ggl47ZLEK3caVgFI9TsysmliIc0DaQ1kmrLQ/EuGp69M3Lyj1zoZqtnWM2Q5D0J
MI2jyTAn7hRF6NdXZbzwlzS1G7jdxO8arur1xmZLsTaSToGYUSkwDNdE8z7hxhe4
WgLUNW7qlGzFDxx3QplbOr+YG/bPw9TlNQ4KElVYusLGKak/IYzDcXkSiGQl+XyZ
qM77/l6FBRYMrobE6Z5liznTmt5nLRi66Rdz3O3Hf9ghbcHUy/AiBBmCGLxVOyl5
wbolNEcKtpho3jPHyZlnxOToL8mW7ESxYHz3T1m2lvJS8XtXcqnhsEtew8GIE33J
MZsBxevRVmt8dGtgqiQvQC3VtmmxEFe+1yN9N1wluNZAXwuyWftEs2os0kp8nipn
Q5rt/FpWYkiduwNRvSQKYKef6T9w/wtrSKlWnCPGDNiGX1oyfUnyjaFQ0B4yMg1W
M8a+oKcvcUQEO32SmSiFMDi6cJvE7ep/JJ1PDu3zSqncxxMvJfjrOXO36RHpCFSl
p/p1NJwlsw4B4pPyubanlJWlqXyDnQofLzMg2qnFL7Hgzqu8lcRRtI/VTSvEVEpJ
++GWU52gSXA0R8IUtbQPAnC0nxl/wVmtgGCfxowpxOFZG6JOuVrLZA8JwDXHvre+
JB2Xh2nlCm5LtMxF5VCOUZXj/VvFoGrq3a5BoGVFa7K7T08Swv9gTWXln7dtHRJe
3ETO4eKQpVegCZZ3FMj1mYsNnZaho3OuDW0XE3PbcfjweR0skkPZQnSBRPfBFF5G
i3IW14EktPemPOmtEr+6+r+0cUXbjLMQw9/qVqoIGSGzkwf5u9IJj0NtV+DsFNFn
WnWGANCwDP7lv3hZ8AiXtkQ1acoQeqlz5xwLrJQtwa7aOBiRESl+I/+Jk+lmCDSA
9G6ufSZIMCLJjr+cMpEqhhbzzzQhCFSnGwCykjsNHyMu2DtWxs95ftEWmlFp1lqm
RPtUdTDQkXs0xmTW+bYsrdPEvWCXCmOoHaqvfSfCydmD5JkSbq9vl3wrzGk410S3
zU1WE2fVuzlOzAfFYk/FVzOFW9BfHNFZvl8tYOnzTQAfteyfmBWEl91Lbjn2uWzj
tyeDmHw10s3+ADPIJ3EC5Ct0N3k0BPzXZPXIY88KvXWdLshDNwsemlRrOLNLtmrS
uzDug2zlOR+q8+9A//1OCaDkRC2MsjDLcHBctVjmyfYMzKAVyAStncEc6mvFeWFr
2+ddjB9CnL3+xJ1+ynqWs410e0IUaWAnxkkhQtmMjKx8vgPgko/roO0T5HTe5oZZ
KPf0g09hyvT80Np3+SvdQOo2IwyEwgcDAIhL26WoXKoIQtU6w9FTFY7r3uaYEt73
h5YnZ2obGv+OrfoVFW7c45u/OVirJxsUixoOweY9EF98OnZX5M3YoqPzPzBUT70i
fMexHYZ4DR0S8QqfUcyCmc4dji42ZDqCckj51v4orIePlofiHOGBKqtwVratFC+P
eLBBzqHJReLGLIxJs2KtKEcJzGFSvaVJhGOgsbJIRLGLY89p10yrIxZPyRvAPilJ
4vmIqd1qr+DSHtMIE5qFdPUN/GHKXB+klxWg9Kkgn/aLvQ879PmlO2Fv+OUY4mI3
cjGt4kPHYTUh96tmR5axk3qm2LR4QwD5IHjHkXAxuJGEDRxAWueaR+wQ7gTNlGKA
04UM8sZaveqdSjqBJv/qz5GMoJMY9P298Onc9xPDkXp2o4x1HVtJEQ720FAXONQn
KsnMfuEITxs4mJ5a0dQkMYWsLzdPmuwEJarTXmTP1uM+yB3AQ/7dvEvCZTc0R63K
8y1K4/v35zjeRI4UJy7p7fLQc1kJ0dwCnAE14RWR3FfeK/MH3un9kPfZjsiEaTju
JxnC3/JJi9qIp5H7nH/0KcHy6Nfmk/WK8hV5jPm9asmb8+GHg4vO4tOkeiNxHDbr
OPv2c2DXbnZn0uU57P1+jtHGAyttJULTh0uOaJor307Dgb+6auTJa/31Siy0uIfe
q9frs+ND19qA6J0co4wS08KnuF4XAwn1cl+w3Ghh1PBzu1A9/id7D3laBpqV+w4x
P8FhjcG2156qLwz23+eo2bJhncrfX99KGRibMgZxDcGXgzCbgUbLShCdyqoG4gjz
0DwS4zkRaRs08g0Fxcuqs8EdTI/Xd4XY6oc4UBKSPjPNZsKN+n2KtosIm8gcRvEG
7MRBGl79aizdCWxtYm7JaW8Q6PxAQRw0rrOfMiLmoymg8/OIf2BKKInv0KPNsdnL
n7Y42sdaIoTR5iLjposYS4kgvv1JUn6LNwbsC0k21pTEgVwzc4DHjbze4B9azVU0
17qQ1WK9Z6G+mV6XyeeMIoFPOe98qMwsyDknHUSTgN7PYKLwcEfYs57DxldYuSFg
HpbjCrr6ediqQ7wMloSMyGVRhhkIQRlJfBFlJWUCyIOm/6VNteoHvYZKTDIR5G8V
Uvi40USTg+yDB0wRQWm6Y1y44k3s0pcpQnM+UF5XaBASaUqqXSXLUwXrZd1gyNmR
jsdzR0eWmzAqQoOKq/hqw2eZ3DioxYTpUA7xUODfFTSUdcItSj9NG9WiUrT2O3U6
KrXL9KZ/lSUQ9Ve3zIF6zRFrasYP9l0GZAviCfHLiW4myiXmfHeNyEodDn5+PeOU
aP7x+vBFhyULXDITW6bgMkrN2VuQkP3a2swPk9CJJxrmAAZgBz+w5fZg+3eBS3vP
cUwGznXVvjK7Vgd7KHMn8Q86O8UTTVa9yRAa2eMdctEJo+IA6UXqz4KqX5y5ZQI8
VZHABxAi/rTn1IMyGQode83PcOwZGGUmgKemZn278ftUgCET2VcDU8aP53KWQqRj
BKvSv+ByE8RniDwKDnPO2ogqBx9uv5qITM80U/2Z2F2uqcvacKy1Ucu+Gwy2DCdy
zLe7cIz4vWKJ0BgBwknLyF7v6BLKUwG7GYpOiC1uumQAeSju71iahqfprmVWyRxl
XYagSQ545Ybg4BiiuMamfD5SLEIh5WYG2Lq5hwuPCWU6qhVHgOots0jPfhbWHi9i
n0nTJQXRpenFuEhteUiI5k3HSdYDdpcwoFKxXXAPgYZ4v5qmcGlP0ZleYhUhCMHg
7WlIf0n3d3EijWo1cqSZmR7wCobboZv675orJGcVFni6mRLg5ia+Ul5yFfZ9AOQM
QkvIPUUKU+eLiX9DxJ9eJqgtoFGrJb6DaDbtzWuKjstDZvblbk0HrjukE+1L2jOA
LxItfKtMeGH+Qyv7LTDQ60RMcGDUuksj2cPUucjJ5/LXti6SmJBTyySRlafatCF+
vltH93uAwluVj69XHVdYHaY6HfG8W0kLE8pTAwx5SOiKTKCWi/EB3T9baOKtSE4c
NzgKrmkHX7ZfOt0Ydg54crkW6BQfxcEzCYOQyzA0C5SHoyWOq624rEhdBlXhlzQA
KbfDgySX7BxRGblVzQiq/eLS6cALANvv28z/jblF3XHQGQMhh8IPuPrew1erLKHP
j60+RgDk/JMSmDny7cBXyY/MQAI0jjrc651aXl1gWZWfpRNP1LkGCMpsw/ra1Mhq
LhQgfmoPu/4BPiH+nggj6oE1YMvVnCNq7PlY26/is9DaTB11t/Rsp2nRBygtsi7b
qg/f5LQVbDmNcAIVlCcGABrDzKqJnSHK88cCYNByYKdPehZvDVeAPea0Hb7EnSVS
Eo8TUdiIVbIPjEUS43NU8AUX2iwVqKGh1gMks02BTa1ew/4MBUFJEIoV+TXFuPxO
S+UmQ+hQXY4Ms1zNECbR8MDJ5pDi4C2AsAfA5pocz5184YYvGiS58shT4v3XXcxt
Q+6kz3SL0jcTCunViJuzesqbnqPZIs4oOJd9dyyCB0jHCkfUfGjYigqCQ0+zp8M+
/clApeeNhY7MrqUfDzRzJ+vG7jr+gTSe67Uzm/pQMcJdkK2hnjQNqNyRfSOkU7jJ
EGqqz3d2WWFd8GZHyC4izADwzPLISYXmGrjSUuhOGEgOYLItiIu4TZV496Qy/gMv
sKOWilQKMCrEmS4S7cZGGFwwBrxlhS5cCqpRu5nXqgxAKLrBrPTQX3STZHJI7pD+
OpHsdUhdbD9uBl+XWpYOS/uGPoWad5I0EoS2v7HbXIwo4Yz9y3XijeMzkC4YclBp
dp0MWGzgQnYbSlFe1lHRfbDWapa1327lBBTS3Wuo5k1ogDOtnLhEKKvOUv/ZsHDX
1G+MKTlORqHd9tF0M+hU8iMDU/CooT0/1k16GTdipdabhu4iRqsejGZsR4C7iIPJ
pMJ/CAK+OY6W1yTzErNkxv3ldsmXZVisM6w1dk96Y3MnqHvQPRtoDWPDTpFKp1+Y
yO8zGV24Cz186G85ijRProLbZDDDhYoDaY1RrWV+7JTNYCCIC1ZwtWcuUw5ZuVjF
IRWl4wvdp/S2imFN7QTPpH2u8We/hFovGCKIyL7Te2HGhOPufUxoznTc5Pj8uWbX
8LYrfZi7nDI55NRgQYbn5/OilOGKR8J6Zzq/7R1EBLE5cbXG/b02LubeVJbsqO58
CqMYlEjxDSBMzC94MG+g2UH6yceU7K2PVPVwLdOIWWVFnX4vvUjzRD8JsYTUUDoL
pHmtb+GfRfSu3g6M+5M+V7WooI5All5CChfM/P0/gOD5pEkSMdAcizCgB3BGq0ue
4M7EP0D1yIpwDg4fwCnCny3iqOBUC+bzfj2Ef3YAZa4dr3Znxd98JvvH0J3DgU3a
ANv4mgKaix3FSIoS5hcezp/W1dOV5+zGVfP5ZFCXjS8DLr4gLdaU3OWHfPBrRxxP
emiaLKA7KWIT1EWhsPgTJo2zsmcfney1NdlanQzUZ+DHr59H+yYXAFXpV9fL65Bs
SJy0xrVs/UrhmA2EzLfBxSewHCeJcAD+6CbfGOMwWTTSPZo0XXmH3VjtXoEWo1r5
3CO7o3vHOeDgrIxGnH/Pge0sJzNrJ/6w3CgoItyRHA7jHyaPz9Ls0rQ3gSFVy60i
Qj0AQ9xaGL8cB1EIOTAHxq6lsXOrNwE/ykUloet97l6s0mIIQFQRQZnyV1H1QFZx
Gb6PYF/TdQtToLTsWDH/Y1rnvmq/s/fDk33533n4dQLadWY3++4/C5jeUNp2VhDZ
G+M3Ya44omgbOn0naTZpzvqpIDFLmra+z4bnmc6+TABPL08yOYMSnTV+sh6tI78o
llw3zEdVMFfd7vFUnlYBdyYwLomfcWpRq7f6do1dSgsyygk63TRJkNmr3L6ulpPW
eHNlLJzRMLmzIwP/hHNRuYCIQ56cHPDGMEjeMEk5FP0dTIrqLJQpYqfuwgN812gO
kAofZrVVfI1v2yg9U5+CVqbVzLFNpEY4Ma70ovbpwNaR0VpcENuk7m8yzXaY2yhr
JVpQPIPUKJTTO+MfJwit/RUoeYJax8bKD5MsTzsP2bPR1H0QyBp7+xXB/yXshUMI
aki2ID2CCoLDTEHWhNOnE6YIEiOwFTLDS0XD7bZ25QYWAXzScFLOAFp7jn37vEk1
b1xKF9Aof5KqnDFxVu+uONr+8vx+k0PT8vyS46boweaVPzIU5IB2tiUryAHNf4Sv
otzDczqiA7uYIwX8wjPIJy6uRAjx20FIQw7laIMQcXfT6Ah5FRa7j9oKs0ZmORi4
goK5proNOELd95trPSBGeRPyfRqLQOnnKdRuvVN9SOt8Hp17fvL8eH6goJyg71gL
eC1tFlvOt9cDd3FULhn4V0wh0Bi5LCVwlDbO47DmeHmgVsQ0Gh8ViHIIp72rOLeU
HNUTr5EPVP68oqBwGwh07SQ7NKhxr47EugudxN44zixbaR/eV8NV3ulf6cRdfDgB
Eyt+ein6flNf8PiOkbenkd8cxYQCIGx9cc9cTtKFMlFMnq7TwTRMmE607d9orYLP
m4sD5CZnzblh/BcNsopjzISotiC/LykW3rMXsp67dlzv4apmYdTF/BlaubtGR9KS
Fg0EOz0mqyt7WmCswRZDgQ7Ikf2MraHfiyBjQRRP0pxoSC5md0e2cFvNZcjpaXou
/aPZxtcRiAlIq8TbnRJkY1AhTcTliz9eAWlOqmlHcxTAqvgoPmq4H5FY3V/UhPU1
Npl04Zl3QdbRdPbSBQVbZLmZtcN1E7rMSEuWYaWVzSHO8Yp3n7NwFp0v/UW+jyxB
nEL8bU1HKC6p4/7FbwPWP8byahYQf4pWN5xtP7HSu0YFcbUILiyUc2bFcLpHjYi0
tBafzHnpF8gYjCVHrN8DRylSwBREOS3l0FxjpS+eG2St0YS4c5phNSkY+EvIw4nH
qp6YNUjIMf0HRrb/JKYDlbDfeHxZ+NEK3adzEH08jtL/+mgo8sdKv3NlEdfIzD0M
UoQdWTAKvx034yK7w+oTFvA+Zr+cl4vpqpa4MlAXWg+WWIz1DXMI5LvhWgcxqOOn
irSVU/R3pmzBH70Nf+K7Fk5J3RxwXZSlHJPgH+bM5Eg1TwARIYOsH200ljQEafKd
0KvlS7M5VwY4vcOdFbofggYyQIc6Sck2ZmB+P3khUtNVheHySM/ypRTgWKA4p6SC
j9gyt40fMSCogo5YSJYOCP8uzEiywONHPdigaHu+C11sXdjiuNrctcjpqzRkdPKo
fCZ2ulgJlYXPqV87aDNLDnOPvkwx/MdTiapcMar/x8yEyYER6lF95d1xePyouWUq
vWdmk8PA1KMMnfZ6WOPwCc0NNlyIyrPRK4E8XKxD/Iqk4mNogzwwUxNymJEwDMJF
N0DtEOj/e5pvUcU1viIjNbxfp4MPApijB7lLRspN4GP/pz/K+xz+bQcshYGBpulu
D/N3Tah9BtwHpx/hW1oyxAWgVBAaoSTGK0O4vQE+Bq+30/UzVuO3cUTiVRZFVpoX
kDaBrcbJqm4Nupew7lTCy32Nemr1hteXBQ4BdXBscIMhvLayKGHi+TxvhDPd3+j8
eKU9rMq3JTtzp2TFUFszw4/nmVnG1LlcluCoGoukErvtkTrU6z+Kra3HzqidIdZi
FODmi7o2G1P65ZbvlnzuZS+MZUnMIksLDr+npf7SxRx7HfOtbp1nbI05oY1mEyEC
Hd31DG+ENdKlFxM7GTnLmbpnJznBBZhln/W56DRuZS9OoSKp++jnjQeniMp7tr/9
8zqJpdSFsicXXBvqdkKgqtJow23e2nzB/idM/k2n15lqAlsgdfQquEk6h+4NXBMs
CwR2doOosaHQako1mgU4wnArlmgcNCKYY9CBVe/CCpCs4JMS1KTb83GP6R1CjYdf
QkoMenYMTh5ursCXGlSR+zPuqjCIGP2OMxfrebYGDyMEJ8xoouhhbhkqs6tlQWaS
sZslyYvnoGZxGHUL9wWlLzFwXc+WEbAYeXwnWB7srtYSLU0CSJBHdIUN9iU33Kvy
Um9qB5lPAzc8GT7lfV7xEmo4Xh6LcC3e0aRULF2KVwVcq0v89pexrDCCxq/YF/bk
bj8zdospcDAJVY6LAZUmuHOGYjLfuVCvd87Pu7ppAclkk3kpqsBTZUVfaNdN15z2
AwNmPz7z0hRgOixN76J6fWvDiaZRKohtAdAy50EPRqsJzD2TbEfEcQiFnUga1CeZ
FS/1hVp35/Ms+3M8dze+cPqOZCQpalal+KvI3b0QqhnZSiJCJ91Fheez1f8H8Mp2
3U2ue53seWPiEgCKOg18JizsVgGE1ZT3hcSMbiVAxXSP3vNNei+tMAldKva0dcTm
uWX6WIUAaAu04Ke7To0YBJBwrHYd/O+KjILoeZ/atJaxjY5k0BWhk5XvHKqwQQSu
lyIutwQV2Gzkk0Q4mwdbmk25KPnXsGNjE23/igmt86mHMSnHuiZWOzdK0nyO+eyW
wD0fTadIcZsYo6X6oDiODkLgQwHQHNf2Izj4i7nHOxsdXm0BkTL9rBo6FmHyr/0U
KnnQJzNaYx85l0Fr9yOWCTm6hLhugVf/FJfZhyvjp3Tc4Q0dj0mw8mm/8jafa5Tv
Tur5Kj40ueCKizMB28ZGVMoayFdj/U2FQ4M5izTtD6/EoF7jyLAQHRwg8o3TjfSK
clzC2IqZMaohiRIf8m9nnxk6EUmbN7aMBnnccz5BdY8YEw4909zy1ydOAFtybpgc
dLt6YqVixcIm6ztxfuTWotTkXMCm5hSpaMehd2oTjDivfnfaOaBbgM6117y6tbB1
BEOxHe4Y0NwJRtJ3B2YToXjl/LeEnZ4kBDoS4qoKrCnWhRXwUPvqmZRdYjNkprdR
5NyFtYRH7zxKGzrKN/XNF+jzVCf2RivVsbTLSsPzuOjZK6kUS3y5guJUJ54uDO0F
GVEUmQ2mQsgIQB8a9n1txVfKo3hmzBhO6/JabwFrC018cHf0qSEy8z9dZSzwSfjI
HkyU8eT2LQNxQQwiPYjPauH9w7PkLS8I0+8JfzUqBOMxgqor22q+eoCGBg7owlRO
eYkSeyRal5h0V9ThyIDUojwKRviutaCK5TeH1WfDmwnem/KC0q7VaBGzb7KWHjE8
xiPwlHhYZ9gIQzTmyqEOVHXvQ0K6NMw8FNXqX2rxyGyhC1j/v0QQjdKNqgolopsO
3tuOZ0V/f6vkBos/Qc5Hjyan/BDxKbOe+2a3ap6BXyK+B5PavhMmQ8RI52mq0Dq7
BuiwzW3ljksqObd/EaUFtu+qMucwXuF2NP1xApJC+PpjNUm38I6FZkfo2D0ACBg0
H4LVTuCOEc1y1AlodhG1N+v6poRVMcMewVtqwy20dKZnGHPifshpQGgbeqAG1+zj
+elh/pbc5hrAZYVKhNyBquN7YEvGZUmHE0/DB4cMtLDkzgfkwVRXfeJOLMLol2JO
Jvms51XwmPrcP2btz6Gfud6FVv4jyrbusjdfhzd9ci+QypDl+ciEim8dfTrkMlkL
9D4+74qyzbA9a0LY/RnC2UMKZrXp7uOj/das2TDXpRMmMiyE/9Nu6wAMPtBwYzo8
53HtaDfrdpeiTvmLZ30vr4OkXruQG9UnQggqeTTvOu2cVXglICLi54jhqX+WUxX5
iVyccLlK/oGp15lkzUkS7axq8ec8ORfRxwJO5cRpx7WiRd2WtreQzlgQMllrkMz0
w86ImLcHpgarXsZ2KjhMPhpEFWNBnyZLCptNBSdOyW//BNSeA2W4kb8r4/pygs5z
1XbA4CSjd8h53RK9WeOwcKxKVIeeC5u25d5mqd6sSn7TTg9vbcqtxWz7oLQvZ9sd
ZUOdewh9QV5PsDa1y0VVvTjxjncmmLv0AEJVM59kX9Bi295FjHHy5okFGCgt08Po
LwM49LFl6KXit22PklE7nx42W9W4w2qZ9py+z03ZWcUP3uV3rxkaOqREnF/f8BrC
bsypk2a7pLwvjtnTSj9oVLA3rYv22JxmuVRyNKeiLM0EvIrXN0wzaP9UbGzkibH8
j6VlwvvKl2OVGyjvJ/5vVdKF/Vf5ACFIYOTU+AqLJzcxjpzxWoEiecu3k/ui8PCc
DEok8xw8RTeHZyYwo8SkvMlTrfdA/hi8bLid53bMwDf6qovGOPOoYjn65keolQua
T50c+VJ/r7xHqH8T14dAcWFT1jLad81O3xlDou8oMRar2gDMiTBH3nbuAZzfnZAQ
mRomz7z+utnaQ6H8DTovfmA5uBwjQ4xnEgMF0peN+2236vo1wiVejM4rs8PbkYxE
y1maZqYaoVSLd7FcQxjuCbhXZrpsBGylVw/GUy9Urwcg3oL5C4/ZVZC5F4pOQih/
5TEJIQQvjwiqVlP7oFaWch5IZELlh2jYnyXobbpDDoKWz97msoO7ZgA34XLk4orf
CZKurBUw9Ys0VvEE7uKHU/OgWUlNU3tuplhNa+lx0BxLE5OcCjAw3+VddEy5TsJG
95iyv6UT/glD/hLt6z5qR+0hKZJ7AbB1sCd9agjNKniLHHWAtCOm4jXF7aMDRxsW
4kZTtzQRExh82O9LZCw76wnSTBVTWBFJgAzFHtMyzejL4A9kINR/HQdcdy1bn3XH
RdeeliPp75xYBqUFawSPiRetrsesNqajQQpavfGMY0wM8U+gFev4ggxc+9q+CqOi
j0rrKgxGDq5iiGGsLRAHYxlZmBjWhcfHgmfy5iox/APtwSW1WiKPoJ+923JnpPIT
PL6G7pyXdgGlmQkwS5Gs1ZNgPaJ6HPtvBnpI2WlEWvwsdtCcVrefqLQ3xH/RXYwY
4mc2S8plhMi9xGACJnHgur9QILLhKRnPz4nWoRe3VN2X4C5pFrN9Ls+ustolbHXI
+2X1DbnBUF+j7VtM4GUIz9WtGfYTjLUuXB0MCiXZ8vxMvtebVcn8tnGPfYbUbDx+
1+l/YGoGFtfRMQ/ezk+Z3E+ndLVC/6HUOdVgIERim6nwsAAFkEseu7IDSCuf7CK6
JHV763mgAlSqJ3XsMSUdl3Q98agCNzpR0NjJa5sN8DrCWXUQ3qropr2hA4a45uXW
AkSX3RM3wvq7KtzmCE+9+DDjU1XFhgptWMCa0KwE3NHE7FyRhcVvYgltROvj5bd6
zGakePTvR+ps+TGA/oOIeaD/4gSat75Ez6N2NTrg0pNx5/N4irroJBxJ9vPT6Cd9
UIU/j5i5JHs6FyKmFLJ1PKhNexLZ6eSqh1q6bXDdTkZ/L9O7qCovEv6paTI+kdhG
MffxoWojIIiu2XDL9MJ3zDMeNqeWblnrvLyFPCwSVncQ6Eec7Y89AxxKL01V4H8W
ytHIu3bNIG3bIXYPJf1yQYuaGmefSRgKbNN771nCha9TQgqbjvtjcolVoSM2EoI2
HViEIoyd9wmHBmPg1e5LAYA9nTF68uKwtyjZw2s1qnyungyB5nUQPYtK0LhhXZdi
7WIR7MMeV9fofErx+6EX0Qpdw6sblxA1UsgEWEpQtfEZNSWWf++L+kCXKnVz/Ftj
6gVP8oZ8xWl6CxWLLzAuPX7n2zAM+VKulGMtrGENFVvsHkWF2Ee98TJwyO05N8Tz
81iI/ZcI30pmVktsu6xjWRRwZ8Va2xR+ORgLIYuyyQKsYbAwsouN1+1hF5+AcsWa
qAS3jMpywwFGXuEIcvfQaJM75nnCSpDz4yyeIWiXAg46STpgeJFAy7qmhTl+DZlG
9H9OXlP6K0SJj9qj9SG7Kb8+PC186NUOgQ1S7XWjdAGdmFQovvxYfSmGTHhjQCA1
nkdFV41WJC4WUvvihkSOOdB7mBGoryQEDtfigQ0l2+adHuuBSg5pAKd3q/pS2j6H
pukiLfo7mGo2FeFxwi/S6naMOCjI5/LXgIoJP78bWxi1GUaERmUwga9EKIv1R04q
dHlsGJw6rLwoB+UrxxHPnlbBPhVGJCQ6I3ANR2MFE04Y913Qr7HM8nR5JDkFMcwT
NgCIRn3zNxz2ymqTkjhkZzqnxcu274FrWjXAoC3FynbIQwR1g2OHyT08D8yefcJm
duHfw+vr8ZudZ9IWM4IrfG/2yxU7aCQfvhHcmya9hfEKaUDD/v/Lm4UHpT/Ix5qo
DMgEW4qMzOxgXyhHfzSCN0aLt+KEcbGs7QHUOYzqFU7didfSbYqc85AMpI2hekgG
+w9IjeJRCnbUY3RDaZVPoccxTIbawTNjMtdT9uUZwQh//mi9TyAeyb/7b0Xsczil
Ov07Vdre0UWFwSjnNf7wfE5oLk07PusCg2tX7+dJhKr1QkijlLdYg2GHTNDNAYw4
lTcaWWMTk05bewWBXmWMYZ4qbrp01lxTt7MCvNt1BGevmFkCjSPEcX6slAoVvyLI
8p7ZvRty6QAcosjGUKChIDU9FPmG5dtpgnMUvGsZ9/GosJz5MF2ad1bFYZs7oh3z
uRCzUI0sDkaZuQWx1ZimN68zahuX/EdjgHqs/AiNJwun9WfwVUq2ge5c4oZN50AI
9CyP/NMnZYc0X7LoCEdrwJGd5dt5DAMR8CBBqoLocPQ6x7yjwnhO6zEzQA0DGPqq
Q0HULOpuwAEf0pC3Q0kqGCOfzyyEjmFaiKBN+AeeD9fBFKcmUim6XHO14T4NsajN
La4AHp3tIeKEb8YRasmYXblWZ7R17GAxu0ESVRGkJqt4IifAKNweeEYNN7VcTCg3
tFtJXf7LvZlTYvkYrKOoEri5as3R1+H9NfWjjaZMmVIpjMMCTXCS9U1a+ffMNlhA
yRXvKX6tI9NSZGyUoZx/xP1i3kL01qsdcdUAR1TnQb3x7eMIs/ARvAtDJ9MD459t
qjVhx3JMXdUOE0K4qVkoQqZc3j4ygTmLs0pmR6jToo8iPH7toZrMbUXgWiwIYPxp
AYpVtACdHv23EQ18YZi2biVPOjbIY7jkB4NNkF+55g8wh5fYugcjFXzYrZn/i2qy
Pmm16iTLcB9Q7UltyEEbGFqMVU4hleYozn+YoAqmI2qkE+Y+GeDBtDiDfTbNwauH
gt5Pu1Cqaonox2B69EdwUHb2+TxwwNp5dnmVLwvAStneCRZI7dxX2pkhROqhie1y
8mvwK5NemaIrkV7tSrWVOKe9HVCdDPAKHwZbwzDB++WWee7q97J56PibJ7GG8iUK
2Nix2FkW0LYwEb/LlQxUv5KIzE5aGrnFnt7sCpATXQgLVP1joODQlblc8m5h6tpw
ez3URHEaXJCQqrZSacJ8PJX28hioedcfY6gO3ibIRelJJV6cExtql/+t26ifRzdL
N9A/T0derG+QnS21ffph2GmPZ/EfJIcthPuSzuUf4Zjw0Dv5CWaqSyLBiKESBiBy
KeC6XMdvsUPNhA4OQVYT8A8yTATQZSP/Ig+XP1mPSPZtrl5MAw/ZRaHL9xa67rtX
Z1hembSkB9SMJ4hM7EfLD0CEjMgpi9PM/a0Ff7hF+lr9cwGUbQ81HYySt+EmZnf2
GOGuvBPlngDTvnie9bYreJez6dx/mHXrTV3EAwSABU2dandr63Eu6K8Ppsb1K94l
s+LdYUPTiTyseBEyFe7mjb+12GpRPX4/BnxoLTYr4pfW7VPMUTcb4EVY1KIB1aTd
SQzAWUNIGTZMbmf4ISdhZ+t6E4kUW+3w3C4iusa4l7a/sxOVzBopuNcmnxco+BuY
18KDaqJwzqgsA+gra+1sXU78GKyLVmDBqzRM1mBHIS0519cd1pgBjhnLPPK4jAeT
0AvcAdtapcUuy6rRqNFzHpj9X+as5/rdlPcKH4J4iMfSW9e7m+GY9GFbVrVP+teK
VhauzBibaJBth0oMSbRji+FDhrZss/gz/K7QYMuxg31kuszZVlXn6e5loISEg9/5
+g1yEy2ON+rXONsWa/7ABxR6GbaJjrov1IP83/Dra4Jb1/tmZ17e0aXOj1GZIW1v
QM+b77pVkCjWyCuvye5Rg8IB5O4aTEr/v70GRUvHr4eUr2AIHxeyhMSvdEbKSWjo
0ytk9PMxZJDhreDIc+lpa6pw8cUnw1qCGs6Pl4G2vsZ9L/wkouyNHA3MAUEamAYj
aYCNGuvIvd+xxCTRD7GSBue67oydO1LQGjvhbdlOYQodaAQc8booWH66Xd2/bBu4
nOFJ1op2RhenPT2QQLYrjieRe23H1RZZ6x7LhzOgjJ2g6+uMUE6zo4NelVWh3Zk/
cWTuonXv6deRtG6DoYDZpq6MxbmHbHaDzu++9LXUEbGNeo0huNXHiva5+K8sONZc
QdD3PU2o0tyJEnAnoKeUAKlGtOtufClAcQCgXFZn3Yc+57NV7QRPNR3d9tUZR+lY
flYpZGnl4iHFx5cPfHmWwgVMGps07QSijts70B+5AWhANKAOqpy8u4hacf2QHhny
bvwHJan63Kqg/bx9csYZ6iENLjW7/SCoO/dkTjINKQG57xTmS8OsMbe+p3x+Jhos
lzyZFpf87/flPChYMif413zwTr6/Y1l+3xmzIFkJyOdxD3H7lHa5FFtlw26K6/jM
Sb3/aLDUtOcoCi28kOCYGGv5TJfu5jJzBVgn7YW2CUCVIgeCUe0+inLQE+nTPnhH
6v6FYAU9W1aG51OCTdgFAZi+9fhMHqdYMVjl0Vv0kTitg1aTmmAbeanLqMCv3YrK
MVQttGzBHm8Ov/tqmkwChPJIyyjpHTFabPMoiPQkFUpJs6K8u5qMA1jSCFnmBPEf
6CSmATNP+CsqVrSEbIZhFrLqOUWJr74DVyDrG7PX9EUK1nACjvQ/xjpU6stgA2tn
1rRD4aAMwmDBQ5hB8c5Gpiv6IThoVOp4adRFcu7rFXR+bCCAcE4d/XoqhGkE6lmB
ov/BD1TxNQ1xJbA9YUWFLQkBTps/FrWRqGZjUCnYVvoNVbCzsdC19C8OD6abaKMu
8SbtCOLXD1yYu/ikV81+MviTNslroRskGzihZ9cT9LssjRiXaA3tj+cuBtlGqHat
duzGdOlhd2PypCxxJcD9LMqpZPdHEvTqIiJiR+S7ubpoKa8bY8Wqv8Ncz/TNAHc0
Tn0C+o5u2XYTEtQmkUuoNejeKEDeOUd1DoH7bkW6lUbaN4j6M45+GD6oY1gKIt0l
0QVPwO/NjumgZ6/Aetrtl8v6/2dw5tehY4xNhJn5PickQH+COMNarH77u/6qaz4J
q+Gmvu+kH2Vk50NRYopqUiEba7IKQQ0KSh+XcWc6nCcKOq5zGS9NbwPp9h/0VaBC
lcnNl4tbZN936sHESr1Q6l4zEo3/JIFCnQvQ3uY7HSzZHEccJ1C5Zc34VNIzkH7X
6uvEhc3Xdz66YKBvP700kCqVxUn6of4F1KHNJWVPS/o6M6Jfzedu30ql4ORQDdEv
vZZEQ1TKIfXBbqKG/FDVZEfmartPaftwsAvzOp627YxgJYmD2C+k97s3sj3Vwgsc
x/GfAIiIzgqE5hU2t3glS/91i+ryiGHycwfUhr8JVJi6pfuZjqGMGn/4VCkcZ2ez
in3IzC1pwmjcLNC+vtCwSkuLUxyBuoZoUDv8giiU1384hw1E9s2HK3MER7avA0/K
atc6nrik9ho2hPNR83tFVYn3v1IjyqJmdMvjYYHgmzZSj1kSoAWUIcR2pOnBrtrC
eZI/Z9dH91YTt0MrDDWQSEcKAgeNVqOIvaEzMhHtX89/6KW7Qz6i0kz8XyeGor+W
IUyl/8lUuzhe8MdJXtsEMWI8E4BdCjndzZSe+ZGmD/2nVso9vfA4/gn6Qs7QEaoO
VAtjHKeidtwJ/SYQPNcFNixmqQBsZiM4jdNgU7gEqhg2ZbEU4myzwJDvkehtqXy5
eAReCf4bq2Cyg0KTHmNEzx7rdneaR1aRKk1bamWpK3UkS6rkox6JVstzLXpzZ6p0
b13OGjMs/O2o39YByOTXM/yQ8X4xO81LuXK6ftEiV8dyMhlqj7JuqC8ipjKt91la
1x3UR2yhcuhvgv+c5w7HKm+vcRTNjLvW8xUadXU/4HGl7dHdaUc/ya8dJEMA0y6h
TmA1UqObyRI+zpxmEViK7ZLWbNa14ZNzAwMwCLCXiEQm+7qM+YP9cpg7LSl5BSi7
yeI70wfvrZMElEP/HghJkc6w1RvSJtxd189ml4K5V0reui3pB8CyN4vegqK+qw5F
/06o8wyLs+MEYMPWUt2weDBLfWRyvLYiZ6d/a3F28cGd8ML+yHs9M33GMIQIdP5J
WYrrLuI/T6CdZrgeXNOBfJTE5KCyuNIQ2LKZc9Bs/zhzBPKSFDGvsf7AKtgJtial
ANq0P6mC6xUrQLkt98wyxuyqjMdJbAgmZiMThLzjI5Bh1+iQEWAtRzMOg+zP2C1M
Nfn9VPAKJZWyho0Oy73cFN3PwnTmxJIQ86vU5zOSqYH1aZ28qiClQvALWvHFSqNf
GQPAg4CeFidEbHOBzWAzOVnFaSdPNmHm0W+6/pmUZTKWOmpIUa6id/cwhqpP6Kpd
CGxkaI9FmWvqMU3ngrEgcyMoi8JEzTnFzV7Fecq3H/GQtAxQ1soKeeJ+JobDDwhO
2yzXgBiEHDEwJf7++XrZbmPpVQC8GGqMAq6o+hLZsNDvt1O+bv1C+KuMoYBL0nze
WXobIpez7zJqljeebSzZqlpm4wIYNN5h/s8FIDwE166vJAbTADq4ZTzSUBqXsQwz
qOjTAgAy4eYady+hoG7f+nmoLYIt6ruVN4eiMP8HY1CXzbgh0KHxZj00Azi1vnZr
RPyht6eB5vWAPBurX8S68/b9I7RK5I16i0VOFz2eO6D5FYGHujlUhADy9WJ2/2O2
IXNZmQV0/nLWf72uwcMxwynrQyp8qJaIMUGHnu9GSXACFX6HIzWmQXR3uMj9FBIv
LVtBbq4ZNR30Nf+eXG/Y65MicSxHwbpYi8YsOIOmKveqJVOOn1X4VPpz04SihCl8
oXaWN6/uze79JiOCIB+TOgExW5DpgWRZOm3pLpDdoDAODj+iBzoRcYfgJ6abRciT
xB1fl/N90nncUAjVR3ZhpoyAaavQAlcptljkQq5rviwNuNVlGAgDZrdUbug0bkiq
DNpWt+74j8b/xmyz0fNiTFuTPqx6fPUyYGiOOooSyafDEhYF0kXbhHp2iYFpZkLa
S+lj3ZKNHQav6BE0ad5CFTXIgtF1VSyRbbWiezzEfsuPHex76p8k8Szfou/aOXUF
qSShOqV6aak1CkBBQCynV6tvx+jrxeA1plelhbk1iqZZpfosXH0NtoXc8hL78MSL
18hQBN64E6oFYlj0D46HI0a+4wZUuLbvu0LlcRp3th9kKMvqtiTZzurKiFGVmiow
AO3qSrwFin1y3CJHZqV7ws8AZ4FJa8Gsv8OszQV1phD0LpmcjMX5ZCS+qyhNKrd1
QKco2KAg8HqMfLgw6cU7jL3lN2uGu8mGvb5c1mTAJSTMzAI5bCbeIN/t8QPhRCa2
3Kh1tZoduCCz4NgDNoftu5iea7v9lpHyKXa6u8wZiDyvwGo9zlQftbYR0owNFsJf
70HuSNdO5XnWvRbPBmDv9YUii38Z4NIUhxE5PFVzw9PzMOfdpqRogF3+sQO/xtvz
SMwOgbTFUCPl//bhfoav5gwtUa8ArV/R7vnBJfatatHHgLgdJia9LZNzJddKSZiR
Rm0fiNoOOXRl8+QeGeu4YnqUKabmqAE01anLUCrO/SGKXccdluI0+FDMzKqWpkXg
chJxw9DkYTHqDD+XA5mFOYskFWOchVc8/wSHrHgoV1WVmyWh4McNJA2gEM9dk3MG
h195wHhcgLWcr8KEOclCTN0vlellt5KLh4Y1fxnWYwY0it5g/JxFGOlENYgblb7L
Lx4MCV2v5pQd8lPJzBsQkkv7Szu4Zqlj3jV6tf1xuwa4P+rzaJ0zIqG0mymNjzf5
Etmd7Pf4Zy5Pz+nxZgsmaMUnoV3mlha+LA0DnUM5/sFuFcv5Nc/d+YFR52xOk1rz
RTDKnb+PxJPjrnGT42Yveqr3VKDkeG2n+nU4+Hf+FOVhLXNk6Mmsyp+a+0TCxJ1T
xD9f0y+h8vIUgH1GTeL4DsGoIDpqQJpq59951gcNINhbxJiqr//n90zWvPXooKYx
e96sfvMOoZfcPnEbPnyH84tMpgjqfUht/zC1S5hXuMsmRc7ZdjvE4wxJz+LwpoE8
r8vdx+XLEEZFU77MvDPRrnOzm+ju5gOMY1HsI6jyJMED02U5XTg0UIiN/5ySRfOc
VJ5Z0YqrQJe0iS2AjG9Em0yDAGjNbsDJ6Dtuz/l71lUDBBn6Cf2w1wRqibsgjjEN
qZwCLIBQShmltTY5J1LuyJwPEQqaed7piQhN1EhQamcQarc08TfEfYDtQbQhIl7U
meEyygn+2TuseL+LqS+6PtA1toF8VWCRKBA4GYuvqK6KKRfeHnto+hY7lz9O9+sM
e6cKiMDPXP3XP44GFhnEkgAwrE9J/R6CTjgJeF/oMDLZwrYmCpxGaXyYj2kCGF7P
gTsW/3gIcq2xcl2cgNgVra8yzLtcinsmxIbEPHxytOTz0K+CbhMjVtAelF9P9ROm
WKnJJQ7j43xerNRFEhhQ63WkN1meNJZNJlWFQ7+SEB3ZLi4vfq28bU8zXIg2qGpm
RRurBWzIHizcCL+YQPbLeIc/8OOSOfu0wAqXspFZkFJTJxl8ANSlRInQHLoXYhi3
cKllO+Babalj2shWT5s6f8f0ff8T6nuptzbzAezrAyEASPA7PCoGWsMGTOX3E5Lh
IKMY57msxKkEjDHcw9ltuJaxL+KzG/493jf/uqxg/s22MJkfMlsnA10zIi9oOobv
OWiZWB1HNC04fNNobdpbXFDcNJaulfwV8ob0TePOJVAxclGqBIciWLZ75l5L7kRo
EfmXJX3HzpQcaqnoOVeeXfWuS1WDbNKuiU8k03brTmaEFrj6FXMkEDQBvW5tLtUi
JeiLVGO6ZwWt4qH5cZn8ciC7xXNWDz8GE3dNG0T9iYR8qUuzdFdWfikW1yxQOhg8
vBvEDn/VKdsMjy0BcPGzUsaA7W3Ds/ko4VZQ0sV/be+FBg0RKiArsCXu/SnQ1BG6
1HlN6vmp2+19+CSTJZ/MDMvx7SmWzaWNuv+1uOPU/5o=
`pragma protect end_protected
