// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:37:37 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
mUeRQVZ/SN5k5GkEQBkNzMpo1FDVD7MjKX9LJed4pkY312CQdFmvOreST5OCjs9E
itpXVarGFdBqDl7/o8HAizJNgXADmaILtdRT6YA8LbonEJThCxF6gMTKKuXNvwnl
HHELGCbFcd3zLBVVIsN1USeA1/RdzgJUZrSbDescz+g=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 25408)
2/2cK2olh2+qSTLZCfNvVZdUPHl6k0UvxIHqkQGZaLTYJ+NjHCMHKEcXkd0WcOHZ
fyN0jPlTBYVXoKBDrQ7Rh2xvSULSja6RKCCnZ0MhpqC/39yC0NLbYS7zt6mFZcWN
IOgsxzeZLT8XinAct9hiYqayMDawaE+oO2G/nsErCmIxxY1jvaAUK4BQM1RDn9Th
Vyx/qOLuZVGpW6d67kdG3DKwW9UeubbjqMU/2yaDxZd99i42A4dpE2p4vf7cfNq0
hOVBlcLNytYYoUrNzEcMQYL9vad56Gp0kXMOj5BReEH//4jefM1t4wIFTAstpmCK
PeKvfMKEW46LT03/FZrroKQPv0npWmZWJ0e7rNOZIwSnKDe9eI1J8fXHm4PV2Gt5
eOsQrjvjwokmWFcQzNyQSBMz1AQL2VitzIKAx8GHFPefYGk2kLop7ok/iS9OTvh8
igYxXTeA2UXdOLwy9a4WhHQx72X+FSxKe6PxdTFreI5ghLj6GPQBEBEAQ6CIT6XL
VzU6LYMk39v6Z288XuCzKU5UWNVRAqveESp1/xTdFdnrqkjPXMk2gIJ7Z0I4oH+d
rP2KhOkppqr1CIM+Wvuz+OJat3yQRD2rtMq/mhNCwpTJBU32TL41OBg2/ZFfXtgC
fNs6N1VgSZMFwAoCYNX82BuBEPtJZkVxuhR2Jl1UsTPM/11AJJMFx59uUrmvwxh9
6mWAsx3TNmgRjcBrfUAyfLwbVMIfJVysZ+ZgYJDf4hJuVdH8aVewxmwPHFr82HQx
x0f5thZiwCXdsutNgAePUJqbmlYg2eOsJctXUbCB5kVDJK6K9En9EJKZ4g2MIuRL
T39dVyfOORD2+CgXzfrGfLFyuZMdJJ4reh2wgfGVE+2LOz0SDs1wPU2jSxQ3uOe2
ppjfeQ8z2r96HwvjjWE8dz0B9053Inl8ejvWAYlx4ED42TP/kL4Dj23RQ/cUdP6V
KHqdheyzlBbdGcWROgv09I4kUJ2Gaf1oGS+BAOXz3+slOGXf6Bma4yO+Q6CDhPof
5JL8trur0oDJCSKjGw3puVSOAzk+tTRZqCG3ujJULL5dAkJ0B3UUXWNqy+QfiD/O
+YEX3mLNvbyQH+UdTnMnvbGDVnW0K9QjzX4RALQyc/O+a9SYZp51JqHoiu8xhUd4
wCgmdBo0zT1K0sMhs0D2nQXD3VseAIVFAOTzoBWDosPlEmCYBASybPkb78lkP0NY
BEWs2uP3oAUgCfgOw7pU24mHnpLYyPjoxBkAijqOfZlrR3KEzTll6mAnZ3BfkHJd
K1LSKFrQDBa1TqCODiawrrJEnEtwUFErMczjkwMOcWDdJFr+3iD7AseDRqJcA7sm
g2kxzcl8rDlC8wEIRC7Siru0bds/gGdERVnc7uckXHS31GBQnEoUGVuS50I57M0a
p30ctXLz0Rkchf+QCzJPhBtDflnZYYuY1upcZwS+bI2NekRqSs6WJBuBb9R1QWyB
WOGdEhWKTgMoke85/dmJdAAP++pwhU7KZxa6dX17Dr0eb7UBYi7cliBiEhCm5Xh6
PR/OMJsOsvEHAZ6XUq93dmdtaXr4loTfRd1l3ucPdSpus+DzsKEnqoEJoj9roL8N
z5KO82lSHRpggbbjzWDfNjgDOLDTMVxjuwN65i6wtf2BFNX5U7dhn0GgMaUlk6Mn
AIbXzJJRJP5YepYVONr8TEHqFoxe+hhWitdiu9u1o1FOytjvwZxxNL6ii8AsRC4B
mUsGeKUNWSFqVfcRmYwtyCV/YMQi6QcB9LOyN/ixNvPZfJKtdeJGaxcy8/DyVRZ4
K9tJlKyGQWkm8URjleGc7enjObvHzr+Y1C2dQMw8W9Csx9oCNDibXGVZ72FKa5y7
l5oYtLolCd2Jqy/1nOUBemnRJkMr/C2vpog6Mtz5P+e5VwRZg98QljoBIphFOfR1
3FheCjQEx+NX2dFLYzX5H8AcYGxR4l+CYRkcJ2xEboP7MWzWCMynBtAUPfQp1jp4
XQzgLu+RFOvLpzJruHPkGd7peFzBUB7otfetkauOAgNSt/Ob/LjQqeK0pcJCZm2C
q9CckPWNmJ3epHwan9xpHQYg7STrh0hor1/1+JtRYvNyet7dMBep3EHbBmvw6eVi
PCZXUs4+PsiWFjXAz/k2uK/bfxGmAJF3zXK2uPW+yESCcKhz6nZmq1OOYXE7Wyvk
M6mh13m4ccOgu6nQFC72GwhP1IZinyObBFQLE83Dh45LaN1+NuqdWiYujd0G7qCu
zbeFLK6irawpP+DVO7j/G0ze9kQxRfzrhpfnmCdwvw6hHMNKFG/HUzfJEMIZYjxn
A6AVSs2XMeyxVY3NoIYh7in+ppsp71QyB4k1gcUoEZ2+mlCIvx0PzUCvCaJEepgt
9XSM0WcG6+4lQK7vJzC8VtcSO+RNIF8aS8UL4mk4bJMBykVemXjFREHNvQM9djaV
hQZoiF6Ch1GQgVbx+JQ666qPz79vuGEOifqvqPU6cUywSBGlOPsQ/cQ+Qy1CdbVb
+7fBo3dfJKnb0pziG5aDL4MnjIwuTaRFERWGvmt5z2HVWtULDKYOxo0F3kGMFfL6
vNpk+Zz4HtDMy1p/nMUZz3/eITp0sRYcPdjLf2+xfnX7U9UaCVkbpdp5D7LnYQ1V
rHRnW5kjHpNk4osAXQHcMpf2NrBsEvdQqrk/bJsyckL1hh218BnxZvMmCZReHfOR
f+tJ7iSzlQAOdkx2GoBvWXbdapkhsjKg7qyhM2UNDVEhp2c2Q/Uxyl96nkegJtpG
L0W9W7hf9Vri68VvPEiQMm4nZqj7FBGtQoInPXMVwXODk6OFnRV51euc8Y1/75RT
VASpd9TDKNMsuu1WsSpJYCmyx2c/jMYMTjGxlc9kBse9Rzrrd77Hl/SWa+DUPKNh
Mf7g3h8VDKNJ0sf2NeWcsHH6LXp5YfEzHpQrw70q+UTnPAenvQ1f8X6kU9lFnZHv
iA+/CSFU/NJHcb3C5A76ld8eDSb7ygIDxNxuHAJdoEeTaSH7fSllSjFfG6egbaLB
PgxSyGuZRZeDbOjiKKr6sSN/HEzQgEd9hKbgCyqTDF6DYY2fvwN+Hn5fK8KIXleu
TCbwSgskUhLdHx58nvwn7viEMgA97mnX8Cf5FgszgsgkCtyuFYeLUZl8cVqn+nzX
8CE6V57faWTzUqK/SvQI1mLYVAVqUzzqH4A24DOFLYXxsrOf5ASd8tMd9fGeIRuc
iLEWI+MVdPoCxJMMipOuSrX7ytq5Iymzuh5i7ELI2eaebThR9sLw9jC4jXh8sOWb
1zDqkt5CE7g2cUVlnnEHEdwtlTtqlfcRQHuBWoLM+Qi/uVZtrBWLACmsbGs7p2Yq
zqk5+ttJuCgJCNnJMo/JiaQ8hVhPJroxgr8bZNfTsnrwgmvY5Q/ul33rYyjoZRWd
Phvirwt1vzhxJe1z27M9Wwuf+BXE5pLEGkyYdZ7a6PThLQ09GtiNVuhszFZldSIR
A2+SqDhYyhOVlAgorYWuQaTCXYtXwzlteh9wP2S7vVzxB4cLznAdzB1Kf4ZnRoVZ
BpRE9t8LZEZSTxqE6oyHO8/CRt9mvNJdeB0ELNDSG5j+lg8vhFAu3XtVuoIe54by
NZ9eTJPA4mck6k0EirMGgXnpSdGQIP/BatkorlSQ247ZUkWTKcVQJ7RCxnuqQI/s
+17/Tu42OaAp3mVdR5Ae+X7NtLm/4pvjtpo9mKxWFPb0wvcaNujNS+ZTDU2eu3Ix
1LQoPWXkUf7LXC0sACGMJ9W0gYGmSjUwz4aD483G7BQfhtaJYpiNxe0XqPI51tgo
RCggp5ktTEelmHNvmpnwLffUl9KjXcJo4oP9oCLNa4I0heemcLzi5sBNwUzGo31P
03aLW68r41NoWDttBuc1daZIyjR4nRJmzPf7BFLRIlK9odvgvkAQMleVAJoKpN7M
+1S1/ZxJoRB6ph8yPramYPHySn3xHOXkVnV57deWVsHemMCMQMS8jLd89FZTkbYy
ItYmFlPPW4/RnYw2TkmAP+Ed+4aDCV2/4ijO9VGaCp9HLneopGNDybm43BN994Af
1G3oIOReqc2a04iCudTxhbEdo4dg1ofoTcGQkqsI7hQWxlq69mmNpGxyGkgwF236
3/4l4yY6ghpWJhxa6Bs3RoBbLo76Fuk1jaS8A5u8B6DBN7ul6qmJcgi/wcY3wM3B
amIKq5aC8YA1o1o+380nDVyTueTM6+TDf9LhIzUWkNslIEU9Nm/kAqSR9Gqt9J6Y
oC3ZyzzDYaCb2fzNQjxC6qG1bED1pbTYbjUHSwqUR5s3RHjxI1e1kR25rMt4AELR
NiD0U3n4gZ/o5WgljY8g4lCpJ5jUzz7o/XgrrtqylAv6N5dxb3nNJXxNIXybiAci
cYSbdG35aL6k9YZiBBda1fg4o6mA36kRybvonJ+A4Ef7aR0Yg4I1PkXZvDhLoqG9
DBtp8jHt9Smn6ViSph5VDIureeXa31cV3ZbAxX9FZhNXnUNKnjAg2w7SaJ4LkM0L
04iPfzwyZfunH675QprCkhXfY23KNuodgTaEoJKh606uWEL2y24sdlkHtRxJqMn+
zt2rCmB4b+fQqO6mFzPvwM0y58Hr97am+HdIBnAAAGo+BPmiT1EbmvBTmcYZ1JDx
D5roaONDrSSPm8e/aSHG5nbNVc6SjAdpYw8yAs7dJRr+B2meDrQLXx3WoDHoAXs2
25j1Zxh1o0UB1CIgeIEZUYyae6wZB1/CmCMR6qahcXaMM7hGF1+5IDp/ioIVd1GP
c3a8xYpqtETDXLyeRqVevvwFqLIqRFOa9thFbMyQC96WncCYW1Q+nB8t0b007pVZ
5JK1GX3e4yxFXNXqr0guccPm5V7H8jEx3LXl6nVSKEfjNaqhmmGJ3Sril1D6wCWB
RP6O0o/+t+StyiSak+ITw0k3VqPJxEL7R7glYSfA2i9DXLvf6dWsQHWsWF34X/KJ
3LtCUwLlj72GKmJhyuALO3fSGgfBJP4BQhXe9uwiqnFBTcdUDgvesKA5+e8h0LPn
8RpfqoJHKvrfn0U9JCEPFds/8l05JZZqIOGW1z8xVy0afhkfJnWEx+ignzpVcTOM
jJxptsw0dJ9Xt6LJ5ftt1L7KQilHmQtDqk7iO3FSkWjzvUN3wm3ZuvWGqrSW5wex
Hqi9Dn8dTdoP7UQY2u094YxfIutY95I0NXHe8gybfIavbNHogrHCGMdX/ucwiext
vwEBbnIt3AZpMGQVD7UvZxZGIgJQMP82FTnHZHWMHuMoWa9IbW8mF5O1O9XIoStU
VH5m2rTAjj8TIL5st+ckFKUd+Ja26RVg02MTZxUsezWYJIpH5PEwmt+IFKo//njE
GMLMfJBuAg5gUbG6pT6SPDTA8c2USIV+jSxP6Elp4i3VFeWC/6291Ouvr9DoGrWb
q+jlzFyuFPVzdUG9HHAZ1Lm1lXXB30zitQLxuI9IiM6jfIA1H45yYiljkwMq7D0n
XFw6mMwMW8kUziIXa+faua1ayPmazz1KknxJZNp/fI9+e7s7zd5v2KjiB2zv7Awx
/en3Q6ReW1B5HG2wscvHg0iToABdvYb5xOWSTZe3Q4fXfpNbZ5/p2F22UU/D7HLP
+d6d6U6mLBIfUvTG8uAI7aldOnuNsj+vlpbAueWO8vVvTaV0ykN2SKKilT3d4lpC
OXPUnLLqYPVUhD8yjo5CY+Dt+f4PPNbg0HcAlpyQCGRSkJbCYWLsJvYWcf7wGR23
uS8UrRQaIoXDK/SKdbhtB55HW35yifWsfyBkHl9f6pAngUh//Nn8SWUvja45GdGV
9aH34twB79v4h+oKi0NH60PYGyUpgDF+0E1tmphpzMgbDko6aHKL61aIAKqXgDRc
81biSeSmvyeNyGH1yunY54g5VFcGx/n9UlAdxJFHvQADykAM1MZHcimQsmvruvt6
oK3F6WXJijloE5kpywt7106P5wRHPLH8MPpynFbYPBY67xx692nOta308NZovafC
ldy2ktuawNGUdJzvBDbJyKQMkdMOfjUYjD/mbyXvqOE90c9IBACfQaG6Qmi6UApe
r43vlUA+Y/x5sF/mnaz8gwoSvTj5hDozjIgqYv30VR65tqjPn5T+afUWqV1qIhFe
sxyz1ImMslKxhONY7BXZutdi/mmD+bfz4ehf1K1KMy4JUjft1wtn7dvH/QV7EWzy
FB8Q6VqIUkIpeqvyz9ypm+wVRp+Ppjzp5uRH/LJMifupXQ3PSyr94YChfSyqNlDb
VA0A4cif1BuDlbUFJ3PJPv3H3GfJ+lBZsKgxPNCkB2I9pdQ8fZQbPkuGAsW2SNjW
IpxlGsfsy802LCazaNHeBKqyffmBkhbSYGcwononpK3oXxT/V0bhp2nRVn5uYMZ8
ISOkn0E9Dq2dZ08TdxdpZMp9MvZhCMsfu+ptwWcZ+Rn6n6uxIhoQPdqtWru7IkNo
ZFcmDr8/m/kPldro2SdZ2O4H5uwsCTcIx+rfi4lOARxzj+iOF/CtIBP/jN9NA0It
cgRSgABmqqCxZ/wm9VmIueXoIIj7oq912C44gwgm6dqtcFUYOIjWp1mlcldJbeD5
Ze7xY8ZhQb3YnyL6KTYsBLmhgw5RUDpyxXADPSPlsN9iMqK9Ywh/rcQ75Fz3samB
M9moKYuWxEeWKUvQNed5uUNQEgGp1xzh4JTNdVoA6fIftMGsjArWxZcl/PbiUjVu
cQR4U05M3WlUlyeIc3RX3Ai28xVnWMsD84imrvThaK85IyBpXufuafnxQ1Vd6T+c
gfHs2779tZdEI98JhwcoZTiBaL4cb3WBrqh8UF5DWF3Z9RgFs/JFIt2iNwpbICCk
9ZmOnmGeqPzQL7gmmht2SVlVXPAVCiFq3TPLEjzFy/qk4IjK75VCBXl4H+gu5aRw
d2nf48nYRXBIxJZL5KW/vAeNWLsJv1K8+dWYNZK+sjuR51WOaBSkt9ygvtaFEJ9B
d38m7sbUS6lMyfX6MetPeIGtNquodJnZ4NpygOSSmsmcVAeVk+wBpKRcJQN+ASfY
YMcNwmkXZLjCih243TFo63wRuMH/FNZ3ao3h2pV+j/Y05X/FkmtQuaqKaltVDQVC
momUrubdSgVQGmFiEYMXLmjUZpW6cXDj0qy76iHH8UJpg3l1VMHu/CTructQ0Mpu
7qFf/Iil9Yc9yC2xGzs0+AvA9KKesXOX4rtEiOmNgXMuqBOtCAQmIIUYauAJjWEZ
TIAvLx0xcuLpWZTK7isin4Mwngl5N9d2ngVbuzgy46s5VD0xNLYb2kaMhP6xH64f
LqOA6H4zTrR5I2xrJO0CPFz673n+vdi4hIrblYKyLJUqiNPYP50imZovyP1wBoEA
95z8rU8d3DQBrsQGyLkLFlNllFFnve9iNdb+Q6necEyrKqN/Y0EdUT9cL9sA00ca
xoLWao8N873+MXounMc+TESkNuh53KvZFiGDZst70qhjasmaWtb4YMMBBoxaqvv4
QgcKPSl2kfJJwoezr8Zb1KGW9vELhlV4bX0fth5fS2pcmcxIKZ9jMteN7muTDL0i
LwhfTnAghLeQXyD3+pbKuoXshyj8yUnr0YfvAffvG9jLX/9rNEiWsYeuJyDg5G6u
pqeljs+JAC7AqTadxRyu8Fn0y3bbM2g5q5T6JZHbT6EdIpvWdsSDNjlp+1R5bIZ+
QTcsD9CjYfaNUyk5JM7t+/QDm2vz9RF1TIg4q7H64GrRDM/J7rKvDUy3rTGiQ84y
TNEzybEMiuLIRlYi4afVa30aoA1StKM5LDLdo4RJjAqWbnMq38+ypZlcYinvVBxH
XBoMTD0BQq0M25plHEkXOUvZKzEhCzRQSxCQCujzC6efrpH5qP230cy/OqLGBTIh
DhYby422PL8gAatCH9DvBgPNZgriqVxsYAPS0TLXvz30laewQLknUB6koVNtdPCl
ZCl4tDNz6vWcM5LmNh0qifAJcTDtj4Aatya+ogzFViTf+W6UFK+p6kIlWZnGI77S
O0Qo8kI+vjJdeb3QmEC8jpgPWCC9twFFsJJQnGOBcs92tziuwtf4RNO8zfpLTdNZ
rrOf7P6W7oBMvgFRj7iMceJ05xtpHosm6cfNegwtTT9q8yuQLXVUjH0u/XuSnMPH
uzJgQTpqdqZEeZzd2BovuktsKLFu8EIL72wdWU9+KarWgZ0xPkv7jmGTfllFQCzE
NUigHKFVnjc6ZCFRiydFmkI7Y803mpscA+gWeDdFcQolKH26NoQcRrDtNDyXF1qw
nTuZ4Z7XvIuDUoSS0XE8RklrkCD3QnpaBQ0kBOxY/5Yc8DtqgPyG5rJFQasjDwAS
QSRyQihk6C1ij9EBZdwh1lYDOc+Btzemj9zGJXbrabfo2Z8qabQMdd3yCbXzOsoa
MohQ0o9m3ptqFwLab60za6zvSzdb7HBcx4tK5PVaTO3dpetHu+4iymB1FOGI5ukF
xHgq2bLQxyNQt5Kmj86Ls1H27QHFb9Sg5BZqJpJUm0FhDDg3IFH5agQo2RpUV5JG
QqlQh7Zzjzowl14JfnyGQR3+cvaq2/wZCoo3JTPo/crWl9BBilSo2EfOeN+EM5m/
E8rv7EMRNsiryKIdkpWoHkIEsixHqbpxK3W165DQy3Mepug121PqgekNo8ZF7c0I
bU1FHsWiTSZ3ZZelJveCVy2KCxYO7W2WLSc4jlXIdR/CElmwWKgQ4rbN3ZqDcW/t
0fq4+T5G2bXyzk5hvzLybUwLN0zdYLJsI2UWhGWSkMuc+g+2cOORdVTYcJA5TunJ
bjhYwXcxgbJKizN48YdDkxB9U1UsXdyH3NTxts7lxcXdEZxeeKadV4knJYO0HVW7
bPRu3/CXgFTrSWAu63327CrPbulimPpOOvlgwrny3qn8bcOto+yrquLZJLiJ/CiF
oWI6twyeSIFODey2AcjJTpgkuzPx0uLdb/nYocFGpi59Pr9QOhZ3oog/V7fzBhki
yIIlipkFjwbDA0tekhJudvVjLzqfFMxC9z9yxs5gxedTZHajbRT5bMcLntWmgETb
jP4MFIbMq9+UteqarRGBUvZ4FAew8TXDTa+eVI72dwQDutYwq9ftEZgFeG+fielU
K8TNUrP7Lqxk1H0f5w2ZtFBXo0DPIxn+DzRCX4G5zcwXQaeeCWjcPJ/loJPUuhoM
eTGXmorWtK3uvVqAh9aR536GBzIhhg10w4N6v+HawrlRUQVpy2jCtxk4ViFvgCdS
NHLZ4oTcdbtFAPQO/OWIDHg3cYZOof2rGb3piq+4Nzz9rMmEK0NZ9oa0QNiNzPcD
8+RqB0ofkGWPDGQDVIxYwSsfYMnv79oRqoIY2gSUwN+HvUcJSV0JzwtRZ+Aoj20h
Azds6ya2WsId7mxGu6shdZFaXho7ZNARj+e5G7mrwSI1ZHZGObokoh5FdFOLpKEI
T1cB2n8C08ATZNR1js6OG+zezLF6XH+EDpFG/0TXSGl8eDAoUVDR4sjDTvh11x4m
qNwpGJR904dwR7Lv90oFTtaEZUBZMqZRJOa2/PCKVSgTht9WolrpRDM8T9TdY2lq
bvAz5pIcvInYFle3aqW/Xvy+LF6DukjX48oRQc1CxUMMfswbkEnn7CNvn7lJ76Pm
aBCIC22EostLzeAy3ClGr/8rZszJzEaju5bw+A8nflX7u/ND/BVSNzL90w0YOPQP
NuS0CaGmcaqPjgYTMM8v8Cidjt/vTgBWChHgNV5I8KICBXdxPGcSNkFEndf5Opt0
47h5tITqRyC9NpYfE2IFZjcvWGxftp3/uEuwpeE9eg0nZO3SyrOEjd2AvcW7UnY3
qBv4dXupFUTWhckufVcPpVJrF8sPFNKFcPBzGX+tbqbmmsaH8ANrZECu/rki3nAL
jkwyrlfpw43cbSZ8X4X/2tMEZmEoHflltAhMBujIGETsAMKODdXyJQFmMjMbE8b6
4OGO8V9c41B+M19OHOQKsBto/DbI6brw66bqN1EpMmFr83h0jcryBTEa5p1m6I9q
lE8Z3bEtxRRaha10Sts3YiLbIxw7vtRJXyLZvGF0jpi73+hcnIO3STUM1n6ELGj5
Jb58JjpGohlJ2v9oFaKlwfR5+Nn+5/5hQ462ej+SPBxLkPHdbzwOkTdeMeGJ2jwG
vYTDo5oBVvv3S54HVhkdE4gR1B99Xgd9+5a6W6BEyDleG+tweFmB9Jd4duN8x9Xz
7YMv5tDD6JpifeE86/E4xK2EdFqqxvl1s4RpAqZ0hOwxooBgJPJxJ0BnHxT9ujTu
4kBWCVDFykN2ia8e9qA5AShv09unw30qyUZmcn81iZeCzY9AnZogxyM/wXtilloH
hnXDQj/ywrhCjyVFaIIVEtSI0Y+AOTyGcj3Uc9AkMTmN8hfeCKH+2JvyqtJkgqlQ
IHwOxpPlznx1/shKB9H2z0sq5EoHYKmNATJE0JTXp7L2+mbmEYiiWCRbX7HVU6pF
dXobPpgP0fCs7xgpz+DOPF3SVwsBJTp6DamoMgUc4XTmgMjiA57nnEko1k8/H0gK
MlMQyydxebOJ0wHcFKvVd3n0SnaGXuqkv26rSl1feacZ3gyFdw9rOuzeseTNV1Wl
Q1sHeyMzivpj82yv3WZQnsN5i4O+VRJXSGt7a4Q/MtEHCzHzh2KZLEx3jEHPShzK
7WHEoqEwEiIe8CZnEU3nwhhVU/jjquXAGXjrW/fceaBJ5BF2KWUBOJHn3RTZ8EGD
+JlGFcydDXhSw09F2AorQu2vaeHggtRep5XB/xP94W1YueGKUQEmYEijFaRkG959
lOP3sJPzpnwMS6oDOTAn4EZZqrf9m2qv+AaGY4PGXwl40S2rI4THaCL8dnXvQ1i2
VxWY3jMCrqquWVLDY+3XSxNtsLzaaNE4JnjYgM+T48sZ46NozKlNE4GBMz47O+2G
aJbmF/wyG98HWI8v6ZbOc8eiicCmSqH07i5uRJTcDeGZ9itR/KHB/PTVJSQeMgBf
m89XFvRpjB+BbKosDe6hWLh6bDRgX+tMryvM14R/wOoXdUO/S1qrYul7eC1tnPiw
1coWIHcYSKTTd5NFIUUJJrjcWfSfloMJ3aZH3CvmUQP2b0EWqKfQJkkNh9Ebjh3I
Kmprh482OHkNtWaaxNAQ+YeupKzTT8maaqpHXzZM/YPgedLsxvyGmxrj3a/CPLHo
UYVV/gfRH31jzMDfhF3ZjVEiOMtJMMQa6aQlNBI6LDMepCGY2s/0ceoupSYxB0Ve
nknH3HELAWlHPB+0T872iAsWhZu6tlAmYUZoUuuI4c7nVE3j8xM1ULmPjb37CAwN
4PjP2G7GZHE+21yQNLCILR/lDIOtFHCaV4PWJx78703YvLvJyfOSqw7ZAcsMtdv9
pnVr+PD/9Nu9lYptCHQ2DEwl+FR/PccMojzqeSghn3D/p4PBTJ5/Aor8+bD2Zc7X
WA+bmyTpbT6H7svBaFBP6zSHGIziKhhYABcT6XsRh9eEsuhocb7xfs7SY/EPY4UB
LJftfUL8FCL1Y9LdqmJXZ7Zkyn/S+5zwcmc3LlW2IH7eD1IuX6dEyhSUHO6PqZKk
KvyFJcEi2vk4O0PjP/WT3xGwOYEN94RwA1RrgdN8ezfl8Gjvz2lotRoPdavDysAf
tHFEkQWLHLTv7MQ0oUSp/mcSqMEOhfXB4XeCmbPCt1AP5gb7y0rakhRMZinFAMi7
f7dacEhuQIm6vf2EYRBj6lPhxVtOg1XiB+yrMdUr8QXSoHZ2KL6NDVQu367W1wzZ
29ATkc0afZZcuTLsJxbnvzYHA1oieN+bK9WuV1sMvdslRu21+GAgdq/b6W2srOzy
USD3rfuSsq0X+abunIgLQAbNBBlAn4BIcHay5A2PpkG+Gd+Qrj81wGen+Y1HL1WE
4IMUCG8e2MX8r9+7VonkoRdVonFWiFQOMHNPsdFtALkJVYT23V++7eQy3ClFpCWn
6e4L4Z5JLNICNwcxf0z5RKGfpGOt93OfoWjgbvCgv1Nu+C7lkS7eCA857vPHFHKs
HT93TQue6It3wkl6hQPhZojljMr3D3wfekc/c0nAU6XxevQ219RbDygklCYqUJGk
ySEfH7iV1Fq+czWtBW8r3+SBEX1h1sSAgNgrSedc/qe4GWZ/pYzMcjQIEZL7SWHV
WF9goRwRLEFtVeUXgyMgPtpOfWxXzRi5LUG8kHITviPg0x9FgcQr4MIfOJYlctCq
Qo215OYiox8zJLMSM3hMgg1caqpP4h7Qy/r3ua8tTp6DM6JmCEKIqSwZaUDH20u9
pZaoU8F65+rfQ8hR7MpGpPuTEZ3EEiLEcDISdKGkS6XXV5SgMLFOgoW/+FLWgP+R
ZtDrhkMotKeeDJ3kePfnuXR9mqLN0pu4vHYLErkWfXf5pl+ZnImZd0EwL06M9him
/iV1GTkShARXKZ1Jm7dTreRULFNzyqdd5gWw0LwkXEnqnCcqYr51sVS/isP5J5Ya
O09DAIaJEXUy3TBOI4zBzuBuK5gGB9Vx+BDlk4kckncNkDCAJjZGUqAV1NzA8GW6
9Je+HNMhIafLllvfQZrwI/9078sF7or6GwkPSsVdje+NcxsvY3swsTDc1jnam6pd
MOLJgiqvz6mMFMDafTIfSCXNJ0m2Dl6pGgA0lHHDkDv26t4K165NjIjPQ74FVjHO
s4jvVyc6iu8GaTvP2UZ1/we+wsbrP8rPgIQbRj/pJ7Ge/4BhxDhJ2CXXwW/Aso2n
YpTHJJqPD7OyQqoL5DmTZLOQ/8XlJiegQrDTTriAC+jreOivH6AHRjI5FeDO+vTu
Wh/Ricdic52ED6JtSLJwdJ2V2Vd0YaOzPJn1qOSQxPHfG3XqVR+2yqhfAJFSdGTC
upiDF8tIgv0YXAyg6SkKfoIqkVKwNG0FCq3jvkA/0a4uT1wQCwU4uA8mYidnlKk1
f4+W0ujjQA9CJP+5gEEnhatNj4u1S2A/ggJKvtD9fkYiNb69b98s43Rn/jq3FqSa
AxRiP9zwMIZIVKk98f7tHM4E9GyYrviEEJy6X7jgCkok0RdW0YCN+eZqe61/FhO4
Eu3FoDWMuJ1w/o2kNepim91gOxf0JeVaqswoh0DQVsoa7dvZ6AIuSyZfID9Sgl0B
Y5TeEnixO5FyXw+x2sTSvh1wZ/sISQ6l4QwAZrweYWQQJCWFDPpOz/WV4GO/d2FF
voUAQ7JPH3LSPDZlBf/agWRZChuEVLfSCWDP8WH6+WrWzr6veo3Xn28SieKD1zlp
+AtUjPCfgzHr1v6Wvw9IAOFOsCGfrzAf3TwIZzyg2Qll8Azji06qQxqIfdgDObj7
Xpe16+rz50fYhEoasZ742NmRa0dSpCsbI9YIJKghnrVdoL7uVNkzt9wVBcNNI+av
0q6XcuS2bz6w2x99RFdiXlnQDztdBvw78HFl6ELnX/6AGBR2uj7t5g9zFYGqgQvg
gwAvyyHbM2UWSAPWUdEGKF+6nhJiTtweurRo3D3uz3cNruuK6Nbde5dSTFDzYU53
O52+iSvEP3gPD36ZaDIudC63k3YhtZwOUwCO2ZRrNSdgFVB7k4Jxh6H6giKv44mb
SWjzeNsJKU/5E1PSlpQI2yPdS3uVApV5pWpb0KQWHI8OTAfZRas4SObsTuSpSNLZ
nmJmAx/a0NCMRmMyySm2sl9tC1FZcmUTH+JoBXLMcCP5KVjdB5VxXCTQD+azgLiv
72z17c0RwE08IdCS61xRyPDSEm09O0X42RbBZTOsMNV4HfQtLFqOxyfjwXJrMSHW
buWN11fvP7pPzo+7IgKuvfS0YzAUQi8uvQJPqsyxFKlceUhy5Gdu24V36BR1THeF
qCphhrRtSejZRq6vvomAiuT+gTO6pCbfdZeYSEz9K7OnWQcFuYAEBCup0b8ocHzQ
iB6Emqh7GKVdZPt4rsmLJruykZhDhqVbuzLIPnTc5JleVllNSjlonhStXp2kK4N+
MfpaHp4t8Tzr/DwS/RnxSU9/OGXL/jjXeqF/IbKAnb+5azoAzam7Z4kgOMrXPeRq
bEANEx88QMbjVe944DbjS9BvxD/t9LTjOBjeJAiP6d+ocKskb6BKVCDp/HplJv+6
3x+iTSnZ2y7Epv6APIlRheJBwDmIgG07axKywnzDxACyRkWpuyShwP7yDG5II7xU
T1Xwnto3dLQkhGS84AMR0uPuIp1KTBcfZqgMhmKjOc7hH6s8nH4O/rYIRDSrMYXf
/Nny+cQSye3Iz2mmW/ZnQKLZ12lW1qQuK1OwG251GmLOtdmBEy4bLeOfi9nrCpBX
TIxro4D2cJ8Nvk0w+/rb7nr2m8UU7aXa/yJtKtadm64mpip0Xcxvwnb16gTskq1V
6tE0XMQBybVuYInOsNk+rWz0GZFeEYeyB/NM4sq1ka23ia+yN1Yf8OFlG1mPvC2s
r4fed277LA1jKG5DMpehsWW/QNGBLkM0Z9Tazb8Xgy7rznHvYNe16cgy5YkFiNnI
Q34FMCsYebwj3sspxNbLYW0TiYlyMHcSKwnHzmwiJWnfPnZUKAJ+34XrT9C5xMOd
fBs5D84EJOWoo+21Rpo5fhlgKqREE3e+RIfj9dIzuTqkHUxkfLqvMO8b+llgcWVv
TeBFTtkf/gwNiJXEHFwYCkIqm9JJBKz3QzHI7EnR4cck5935pZawh/pz3GJHTLIf
HuQhJMrbwDJWJ5noPBENYLv2ctykAwIsqTvrzbdVVHLmNfYg/4jseIso+kNlPrpe
Jw4Hn2qFyGhGco9GFFnhZHc0hakrXIufCBGFgj+mf8t4QwqXr2t/JgOMXx4dLWf2
moak2+r61yIO1EsUkZ8/pcbDY9y6ZRRIzoY/iMEhyQMc2fQ30UTSsBgLwNL+ruVe
UpsNGEAr2fOhpKX6ZH0Jss563nJTrljD9dHAYyG4nC7Vj2KNL3/p6I6wtAlpxjf8
f7jwUZvVvUbEj1h+U9u0hX2basiOrS5OFIOGb7RYL9Du/THPVDEx7QZVWkZljTQk
XTfqeh1rrb1yJcPibKbI/hhLiQQ+x70R13YzuSNIfcMlS31RfCZ6FdBqdx2SFNvp
4nccrlQuYaUB90kJ3qhqUqY/meh54N/aN7Vr+mkR9J+6ypWusUasGM6VyU3RGWy4
mUTCvwqtZ6Cl+fwMqgDmramCCIc/aT/P5Y4ZWOiz8d3rekZsJwnQQhtBsQG8Wn3W
TepxBxh/SapqQpxkMmIYm4KZB3e7xbGocwHv3H2QRF36G8LGpsk3zOqVzlooUT/S
cUVH2fhtlrIZ5eOhHAj/xusIlGV9/MFbTnfGXEtyC8PQDFmarYjS5KBkkZssQnot
tokUi66hTC4pMItxAHxC+iUO5NudOSX3M6fQFaEUXEFACnNmVIFTPUjVAQE20YIY
UW6MU1QCEUXjw0JKJ99OGyxnZcI4a/26ITp0OGkDOa5NsZO9Zj1hTNW4+j7Q1r1R
dhmKzBDQHR0Ngf9zvHgGaNHIEVFUfM66LO2sh9djIqejiymmNbhaI5YSIqnYyyJk
C+2ua1kPxT1syDdw5J6pJGPGN7fySFt0QcoJ5JcvI2RttjZDjfreqLj1gPQEZQIR
vqbdr2EPl3AM23LgGZnoFzoxP6c4baq+xk6wsX0V7AI/QHsjOZdGIe4xuExA12ZW
8fo/Q1yFgzrRkyIubueQJR2XutTRp5EgCGmtUBtwDF9xdhNpQ63zqNsLX8pXJIXS
taYlhXtcewe5gxwOJojf+yydVmljB0cGgVjS5V7Igvun6JrxoI+YE41Vhzo4f3/2
ZhEOdXJB1olkYek2Th9y8Kz+KP1S4XSeQ2cZEKE45d9Wrwh0j32lEXED+1hV0WAy
lR80gX77v8jHr/zUJtTPW3iUOmmxHXNX/26gf4vgAx/sVTAiDOiDWYQrlqm27VBI
utj/hf9gnRlIzjIspvAJ5pkZdvk3JDpQg9OA6bAYQODTGZjmQscbuLCYDWbFr7Ps
yc04rHaD7YZs+O6AXYS3gWfOflncjeYYWdhm/HgsNF1wfvQmYad1zBROPldqcaZF
EAFBXyDAgi6jCn+LRbXSzBTZHZ35kQH3lt2CQ6GAQx2zDDp/5fNQvL1/DiQ5iZaD
HDphHSntuF0ICOjWRBxNU/H/UdoUVRa1SnDEwJ52Dn3+IfF3m26pcQwmuQnWBtIV
+3aMvm/9D2YL6OHiJ7wuVpIMwHgMTf7YkUS8IRgiY0p1YJGxF4LUzjoDNcpWLMJz
H869IaKBVg70JJfT6f6CEZTUWlGR0wxICjExa1yBPPJ7IIeL/pvoQKQwyvyLu1EP
JPMeInUhSEcEbaAqBilPaONWKIoeVpll0FWLz8lGsz9iQtwsBVQuueI3Jcm5upXe
5ZlMDOfXuNtbE825qKYq9gEbt/Uhif4naSx4c3o93X8/nPUZexXCt/N104oS++AE
yJh5Cdz/3EFid2M8gTDGUZWR9oiA3ojUpZKGBGE1ty1iLuq/T3/haM6UHuan7ii2
IEBPnx9aRgZTZr22zNJl4+jgqNCIpSrmMFU+rNIeMQguMf88VopuByt+KjIozdOe
TCcbzh6EjDJhrQXSPnXnucWw6L5p+SUgM16B3i/PhOad4iQkTdZfhVtp6JlyOkj5
esJ5+4zmpSLsuOFIzunbA/ZTel9WJNCJIwSZm6aZpiqDndEjxH4o2yPnDNnPClbW
M+qfowZv5l1XjqhbLy0GTBcPmrcgjqXMjUwGOzdcP2cmCdlKZgQRft1CpZ9D1Edv
LMieZr/xE1YHFelbL18ewQGDcmhxqlnq275/eeGyV5gHbQbWTLMHFDfId5Vjxtal
yRix+4v2XE58WIBjGcQ5x2JfouqO8iQ7+6cMxSzepIecJawe+azY2JUMuy5YaMsw
OFXcnMZa/7dAAxvSDqMFdehc3heIcwyPpRw9mGDe8zdC8sl6v5tSD4cFMIan6aIB
vsPOUTqLdQ+8jHC0S42H1CbA9i7kP2U+5D8E9gLXcz6rrsSlFGTbnkWYYoLK+ipO
aYbQ1XCVh6+u9Qhzt4nMPeEVK1cUa2IO/P07gDbZEZpfFGyRReqR0ZxKHTAAHFb8
ej35TkBemm64hZoc9fb2NcOskeJ+hhADEVd8+/IXUfxa5xxW1ngMcffnZCKuu48k
2HyvOK3+2dNiwgfBSfSKct4MOAsceAA4qHE8FkJPTq4a+mLbbIC496A+mWZkWmKC
BCAZQMKylKXKlebyJsrgdOzbe1yrDnnNsFqDz8qZkxpYQ7cIRJxQSS+EsBVImtHU
4r4mJ5b1nd7FdchoJZF6URIHmaFoVVn/e3mw2oeTpdmKKkvGs6shkhIHP2fBssDH
vv9LnVonbbfdL0PGjyo8Um7daBQSqdWyHURLQMJ32WjKe8d4Oa4Pr/Gm2baw/tpL
JKu8kjSb1MoAJ9sDho9PmXZSN4NuI4Ddu3lOsCqHI8alDrwCTAVHtUkPLIKUqWnf
uGlINp/NFllBJ0CqtQxhXrud+2NBb+enqXtpR2qnxtYeViQc/O+vTa6s/73aepk4
Kibb/2Zj/olNtGN7+my0yn822e6jiatTV70hXWWIWK7vbALIscZ310HgbZ8lhgNA
zcHnoX2HExNsZ2BQqZgonbqtTsJjwbE9hwCALXf5nszNfSWqeO4fuzuG6ZmYmyoA
tudOSvQIqVsRcNA+kyarMlvpWM/naU34ZlGHJwX/mJlscR8/KdNn4Q3Ih+NUNSlF
9FSGAWeXNeWjMmmpm9vdjieU9xZCg1+EoX9Maeajn1TwBgBkA9YaeqZellMbcHXG
/f4Ve1d5YLK85FsFYvixTbCsLwS0aseFa+dDe9GLyNwN/K0B/wEP1K+31ernn2lS
TDTVUxKLfXYPxX2WbAs9L9LcPQaIWVYtQ9QlWoFfl/fcvGaEH676Kk+bilMvF3fa
PW+ksiUVxC1W1WAE6McyaUncYO0Hybe6S1wgYDY2DVIFgrMzDaHlomLiZd2K20Ok
qv+ysi41Bfls4tFS0kCWX3w9q9lui6vMoETBCNjQlSZMYsj8qgOwJU/CAIgDJn/r
AZCYB0TlEJAMGyzCflc5rlhxjSOBBUARghW22l1bTJGAYioQ4CqWL1CLtKZs5mIQ
Iwjcku2mE82o5406MtCme/oJvIc15pKYhT0QI9bExa1D/tWcnoNFn0CHqkVSUqCi
ftT+2DGnpoQBY+dc6YhfanQrPI+5tBvGjXO0v+CSsjaBrJehMD0xMZh9awGQGcEK
6jOyRXqP2asXVphg4N3epRsSk4Y5OAtHEge3xKDoANAbNVLP8zj6UFG3NvyXz8HM
k8vRV9v7lCehhWVvy4NGJKbf+e4Zn97kt9D7DpaP9CXF1L4UHkMWnrHfRkSRrB1S
wzl+EeuacBwTNpItmrQcxdMguLdAOmW5KjKpNuv78llBCFxEd+igVkC30C5Yd+vU
ZtGm6QR1wMlAO18cz8l7lUsCo3AYH1gTPYLMZhGzRjzV4Q8DDLY6ZSvHho7nnZB9
EW26TTZ6zFYnLStQBasO6pX2v2w1pJMxBE66HgGXZhMR1+S6uIvgD+YNVbD41HeZ
RED6yA4KCuNhap0arTn0WJ4x5BE62wITGyHqCZ67SUcW9p9aIWg0PqUF/qutzrq9
Bx0pXefc2QLXmheNuq+/NXkWpQE9Q1ofbBjCekUy8S6KqtVbhNB+WruQSIJ6MO1Z
X+64MBbeE0UW4lxJleaew4J86VuLkdPrF07r73b5EsP5DOVGJ5ZVKCqgckT+Jg53
OpA1YYMhULWA1wKgRV+3mBzbdHfbLaGTTnH16BjXrn0XVGUkpX5hSZ0gTPJOwW4s
pzKi/GCvVVonGh9+Eg/mFF/NTu1yJ4U7Uj6ejcgHx075ieUlBvJdUmiBb357vkZg
kdiUQFFrbCZ/oiIGmfXdf6nQ8d1svJ0U7qVxbdLxaFdTX+pqeiMk4NTE0OOgxaUf
pc5jUUWQI+HSDbtO9hmMtu8P5G9cEQriF1SBGl0trWW8dbE6uHL/TTYBRlf6WaVO
8ZCihl/xXid5xec5bJP3i9ETbUAE6zHWYnTFXpnd7feBW8C/DB0efbXYtBbjfFlA
JinVTl4Z/YKSPQG/pxo6iIOAQPZT5m8WPe2Djchb0YE1KBqpj9T1MXMur2drWk28
sqRDy0zraC0f3BuGeEFMUbzfJFNGMiul/9aMPf2+bogo2e61hKFjtSGLcQ2GywDR
oW4NqjwtT7VyUVWHM5Fhw3BsWCChM9NAaqoDsxSxet59YJJJDYfx/rjNr8TYhkKQ
O30asHp5k/sfpnMmmjV+2FcWLX0L9QjQisv7Id+Nz50n5OzUlB5FW9gJJJh2Oxej
JVxAWKXaKA/56OMhTLW1/LKgBE3Brwd8U8FizmDBPamgIjNyWK1N/bmqY3hQmcRa
oOA1zIWtS9IXvQd/txgIDVBZSYAoK/AR3iXWKYkkUQpjEDQN3rlidRR1wSUtyPl1
YF6q0SGGZmQZMb43E61Kf8HbCimzOLqbUbuz77YN4Dje1KhMOLobuf5oA48mXBXT
0vhbCinTKiGabNbk65awO+3Y75ynewQmr9rxyKWGnEeaHOgsvxumrsMHHk2RtGiN
JFlCAjLRZTNH4ZUJwSnnRZUxzbrKMlyrW8jRHNDO4jCV8luhQB+T2GFrhKG+0xzx
BfIz2oI+nVaQ+qdSdD3WEfSBiJ7miZQfXSdz+eVufXQRl1Eqxs3IU8WMWKJNnJWM
RK/QcApX2x/DYncWJp+4Bz7Z+XPGa/uKNiSlh4T0lfYwz04u+BwnfUF/Ux4+eyIT
ue/ZCnB62D6zb224AoMUrvz7xeXZrhGhM3lHg8ess1PMR3UMvKTBh8i7I3TTXyFN
p4SGshGoqdNuQjjv6r/678AbQrO7bY0DnVMzgQgwykQvXf6osOAvl+FOZEpBFLag
/QGXHCzOTahRe7TZNdx9G1vPub6lTyehff4ejr+zcXcNBvuprblrCERqf1vzi4tL
bE+xAbrFQ1/YzW5rs/v8tBUOnHCsOy+FlyoRtBkz9N7ObqntNC7eVX08im2exOWN
etlTcsSi1qaNrnT6iMf3Xk7k61syfqVltCXz5x7urTak2ZAgDtrfR/Jq5pKWfEQz
9t8asQz8mVmrieLQfGgbIBULqZF6gKUbGb8VkIA7kgSwv6JmTgf2bY5iz97HJX5Z
jDFvJ3y+0kCqPXdw2Dar3yRhSlMmoNJvfggFR1iWwol4K3tsBexqcLeBC/W8CIPK
Yptsuz0z/JpWoUG84AmnTBPs1Z+H3Q7VmpMVE89970H3DAyxiSAGkQLj2NUrvsv6
PmZebwaoFtyowZuvWO6WX6MITFSNamgHqk80hzUnSbPEf9Uvff84NsQDpZZFEcls
9tijF+4POJLiFl8GNWb4Zewum+6gT7QYIhwlEI6bn6GMaXQ4LMMx/u9XkxD/WM8C
5Fcy9dFHKVHkZLLflwi9PPf+NVLN7rvl+VgBfmZ+pd2pj3DA8UxvYovg6v1jFfBS
zX8auCFU6w2GNq4XdEEW0GIzPrAEnabr30dzqjh/MwYeS0jdomv1UBhjejn/P43D
LmcQTPwmZNg5yWkRyyjv2mFeCZ6+7Bz951LGBYxEmisVIMHypOS2vCu/932Mxfc2
dzqg5bAfR+clJeNOP/ZSij2yOw8iV0AwYftGPdtiK2UitPPgZx7+jW4mR6hrr4a3
6ODaJVKr2YXycOL/h5m/2laJQ/vSf+uImbuBUrYSU5c154hzuQO+I0mJKITQRDId
t4GflyFUSBL506+Qa/x+vJmTjEk5qziFxv6tDB4g606A5Pz0QsjmM7pPixV0r1z+
K4j9+g0TuQMdUIGsx/WSnhIWwTCq2honFI2/Z8TR0gotahVdspsSp1HU8QmXZqDr
030rZYOu0mUju0OnEiNYGYOJXRMr9Ad3C5TXJ5CtM8yX/+dnojtPLUyDu1cXJFbm
JAjX+A+R2NPweMA1r/PdJWugaAy8Q8VUSrhTGneOwBUCap/qzWr5UzeSxuOjxmhn
qcSB3ds58cHy88NjBa2Lmp7NtuF/1EUTMbTYLC0zQsIYbKgVg3FKhrtot7qexyhx
Z7mp7S2dVlZi1o8kzFeO2iGe+OwHv+n4OFLdmvKQo/Yr1VaahgRxMJAyGPWIrwaA
c31C6xpTbXlGz7mOwVfigquSakAPojvaAmFMemeQj6uKODjSVPZrZ5RgcLJxOIU/
pVfcOLBGBPJR/sCaC5hq4NAOpA5b0eYiuOB4uaVy+0Ix+gFwYoB47x7Oy49ORKlv
oLWMRUAtHmVgW8wsuEEIFPtW4Deh5lMSZnf9/T1ui4XbuIXL3Ssr0r65tRNybrjN
ktOooPB3bUj/PQabnL3sRsjCFOIq8NdkeI7O15EVpIrMLq6lOoHezKEliy8yaqm0
8ZPHI/9PIEAKdi2r3IvHkus4I2nyLooTY34OVyPusJ2R85NEhJtDuZKHeVBgMYIc
34zT8NfZ6x2mbO3FDbnh4ibnFL0Ow4yayhGQ49tluNgDH5tZP8K8KfdlOeJZ5BTf
zhO60jzwz23wRonbpi389Tz0mvmwTMCIoodFJCQDjCN6uNdB+7hdsGFSNMXMsOfg
Ty2Ub+W1Oq57EgZn2ZzHlGSioJi8eHsSjwyj7hJNmaEAZBWY+BN94IW4Mg8VJFXP
3R6t9NHLndzlLXKrmXg98y7iAtwmQ5Lim+zUyGJmfKTtWMe4DQg0Dl8fkGhm1i6r
3nqOWnsj7HRtGTIxiMi0uPteB54LUmQO8RcNUGNAEQw/uYtTWxa/e7/JdnNHrSfo
FdCI4N8+YDb9/bP9avFuVmYWiU44uJLZx3SMX9Vv0GmM/mQONAuWhZqaZKA3ozfJ
zGxYfklqqRWGU+DTg21ypYuP6E/HAK13lH/XRjJMs+a3CtaEfEbfm9e77T5QXRgt
MIEwETPV19UIs+BGW5pjSLgArcMZ9SQIhIvn2tkKUDITUreVmZNVrzGJjRtf4Dx/
UIxMO13XqwV1ELhJWZT3rr5jRS9ZlNxEi7hDcMjWHZPVbTdazSk4vO1R0tPUl+Qc
XVWank52B/RIpJp9I8/7CQNoOl8HS2vN7+El0dwUFrvrcjjxE9nu/62pTICntOQe
8SgIAVG65dq9Fb4Yg/+rV+LpKzfHXdFg762zp1g9G7bJCpF6mNwHjv4MrT8sqZ1f
ln1Jj9sYntcwh2YcgkdyVBfNOKehvol8GHiMbgVs7GE65euaGjj7UknQTvp8YGey
sSCDxeflVq17jHyCbDqbwokRHIX4O27pAwp0rmx+fd8ELOATa/4g/gZNdYQYzW7I
17YZP+QKaPn/uKAzRfQSExIUFOFUorP56htr5kb4tXS/5E1yf7oNw6iL9sDcPlWn
0XvVyTJby6fp7p+k8rMC3RUiHwEgschP5jfXakp8DJ9xGWmBiCdYOkl8KNbc2Rmx
RlMpNEVBD6FHz8Duvmx5e4S7mu7cWKx4j60T4LzCw153CwGkSGjIiEzBmjxYSSlV
6z17VI3vLf7SVY6yP2ulThCzWqXiNP7YZ+wSHxV4NRq5jYr/nx04lqaGLvKm3OHz
KdwFzAWlYYeoJ5sthJ7qOs0tYRrbvHrF0ROE+YQ0MTLkFRxQHPV0vKK190xzuQql
/winkB8W4HO0/DeMmLFaZEIcRUJMcdoPum1dGYcWKU/eyjPbBvnaC0qlE4+vnQ7r
KDBL0cMzc2ORLKnIfHAPIZc7EupMrLHiwmwqG6qX6jkPpsuNsNWn7vcRYMSQtubK
nvXN8CVkb/UkAeAfL1TFXb9kHEv/wwQVbjBHedokvDEbJdNmwjmNr80I+BuxP3IE
RNR07KYa6JiFQEBv8XVdDOY6Bqk89AUqTllRogaL83grkENhnuKS88z8nbWzSMyh
aA8jUGuiyyC9TdRfY0SccRCspbobOjrJcMANgzKRKVX6J+PwnpqvTzTO4EOz+gN1
muprmf+uvXNyRx/NVQcFTtTPNANtZWUWuIsdoynB0PEaXA3OFMUPYBtnRrphiYgd
v5ecEMdKqfHMBBDBVxULnJAlOHI/kMNOC9SyITwWcdCvp5PUoM9KjHY10CTU+qa+
8iFxqcN0Rb+BxH1pfiWvGUOoAbd6eV9TIUQ5+MM+AijQR59koUknPDjrMau96as7
nGaL4oHB287FdobAJwbIVHP77zwz2qwIcnv1R5YYfM8TzkGToams1QtoCh/nM/NY
tTd1+tn7fR9Jfa9+4d47Oa76KQWuNKYk8IcjMGR6dDA4W2NmcJk8idXuwxaBaPgo
nv394vOhYzCzux3igbuu7cUvYfwzTuSX55G6vnmaZwJc1gjPoV4I1uxRHfrLil0+
fUcQTNKLVta63QypIgichSKLvev9LgbfGBl1qe+Phiqof9ESXd2ISnI922mi1AEC
9jKdk2RrF3ZAeFmwDTwT/7fIbLSCoKxxH1EuvFuZX39VSCewwGDcndwsEKGJ+N5l
p1waiV+9kFCzDU5EcPPSvOXnrHoSlUg629x6cCa0sj1Vxd7x7D7h0P5+HCsrL0HS
bEMDvOVrTh381v6HaHGY18DKFFVmbwUb77xptxEdxdYnXXZZjZKYP9GTX6955FSN
HTdzvRpw9carRdbmidE4vJG4LaURPCKcBhOxZHAW9yZa3rMYuboBMPbv0H1+UXxt
JSJSY2JpoKplNm/AaVEbGgkC76NgZ0gc03ppxaThEJqtFYhVk+312eVMI//ZHwxc
7HxQgetEI1GMnCh7bxTO4VSYMgiG0HC8uasNH/1vJmzu8WIG1qnix1c5w7Z3xldB
BLAHA3pAETRomZDMAs+evPS7sB9BI4ekme5S3MsqyYLyZhW9gitqQd2o6yCMaglb
wLMDDSsnLz2DqAAxzZYF6sjGExy8t+947a33QCcRZMZgdh05j5+iaihkWXFf+HRn
Bag64BbVDleDzyiKDlTOojWuV4V4vVvPW1YERHCl4ytPnLPDnh77gD1WUDo4fYQO
o+6iRwbRgZ2p0G5d8b8p9I+ISMc9i9U08A4Q6BXtEx7QvEf6ohxwl9ILuzfUzJw9
EC+grYh6IrUqDkf5LFzmTdOLCaakXgZerviY5NcEsDByWWbKRTLMGxBNattq5ZAL
/ahPaWTgB0+lHn4ojZR+tvlLqFCvNEhoZupBu6Q4ImXYUf0pJhcj0dUQhxmf99V6
kvSc35/eLamKYEr77GdQIZDwwY8yd3YpBvkDi4rAFYo547JV0Pcqf8zap6DicJ8w
+/qgHu4K4yiG1q/MW1hsn5Lhl7ef6DRhYdqcXNvClnATAjVS8doeJmJvBsE5x+g3
/wcpFg98wSwaN1KTd9wOEAXC7bqgrc/M1i7h8xD8ycm5z8fEU5bsf37xV6J+Fu81
SovJtrmSTtbW+RBd4G57H8OvLxAr/2Laxd9NoUQtWcNgflNw5iZrPjWI8aFlr6wh
59r/La6G2IsVBiTB+/QTMW0WsB4F9q2Bcu9bUIRny6OY08IxmT9dg9E+v45Qq7Da
pufF/Pi/HUZgLUUWEMJRE6GqiomY/ZIqW0jhCY8b1zvbioy9uBQQwy2bxID9q6jf
a/iC700Oma+X17h4LcQ703w9xGCH2hzn6mtLFZkr/vTkYHxLNNEvLkOiCAI65XK2
KDDpWJM/d/YbOgVo/fXiZxLdz9TJksJ2xYyQAltJ8BaYD8I0h9Jxvm3ZzKTGjV4U
low0nE21SmgbH88m9vHTATwXbueIa5PPsjqc+TxcZZadf3oagu4RvZ+TbAYkF3O9
V+e7BrB7bCM9A6r/T6JC+5gCp0DcSTmHi8JNEu7wCrFck0Y/XS3NDGNx+ECiiI76
/RxQPJKgYPraIwhFvQ+IJaD+sJr0dZ38mLth38sxRsw8MJt+RnWPnNvSUqpsCq5T
WW3x+7sgmCTmEqySMYqbAYEnxmJ/RIhrv/cMs+WhE1AK+YORyULJn91hNghByr2s
JEVzwJX6pN4X3svzb+JxXb2hiYmhqHDZDz4CHrCz5irZqB6sm5eaxhCJSmGASEUr
j5U2OmMx4dsiIGBn5rMpcHnCUzL8snDeUnSqGyj4sPaXg/bzOtfj6mlFZEPm7AWO
B2bH5etRSFSrJemEvohnIhlyjb2ODeg0yq9Nif2uczWCqSBC4qlOEgR++4G4eim0
pkLhcS1J4lhz58h7PLdlbzQQ4lXpK0RO44Jfyz6ROd4tWWCR154l/131m9Lfj2ni
DHoYaOtdEk1bT/l0dsM1pEzMvIOrnzmzmqWsYA+WhEmVye1B4P9uvmq5fDgmGxSe
h6IqSp4cPAzY8vPPay79cZTLdJiz8QCoiBmJ0Xi1CXCGNfMZAigTNgyIdVLnLpkL
fejA2E365Se2Hj4tgLjSZV1IoaVYBB+wUCf4Ag1Rr2c8kqKRfsjJi8KDujX3tm/7
Cqyg4FuMoN4Bzap/Vrk4rb2D/4uOU8cQZJ3xq2EV4lgMG96hhi99sWrSwK7nFyVa
UILZO1f2FQx8RtVVoegmp9YUOTY3/r28Q/rCX25NVsn6inM/1aeXkFAFesi7+i7K
G2H9QDN4zPIx+pKQ/L5S6NjdBJCYQSqcnx67MAy4H6cStMH7Efwvr4JOnwssbSFs
czj5jFjWi/omJxq3qgySAySozBwj5cez+atsasp7OU2gKMOXS3TWuiG7IQo7Z9mF
WK8dzGipHy8PEb3Z8wedIzPGYX4knLPt9wDLytZHj1yeyK00EqZovucvlHsTIol/
4/S4QtKfFbLMxxF7MSKHRB0d0tuDn/JIMO7DcPVJX7JpgbxdHMkuI+L+C2lAW29K
1OG3CNMDCVaukknF5/P2p2kQuwWTq3BKHO6HRJUIMOloVIqbiQKVw1HFwZgZpLU+
W9SlU+aGMdkADpsvLU3jmlLt9Sk8rtOBWkKTn8ll8DkriRYNiYCSxFTB5IbiZzxR
86aKIWL8I4yXqnRAqwbZtFVg21XH4iP8xWvdPMYsPlhFAX1ViC7ybRqu78Om6qic
Klq6aBx6YmYIuR/bpYxsYRz+Rh1sjROaCSPDQmbbhmW3NqHHAlvpYe8Tp7ttU2rA
0YCLt7C351KchMQR4/tHSlM8aaOvy7+miX7BzP6hSM4CiWkBZFe90YHc6w94c5TW
K1KIwEPP78TYFSM31AXTOPK/lJI8xzEtgjeLbXS7NQl6pA/30/QkeCCncdDCbNPy
+4JsKi/avk6iuMoJOxJ6LhJ5/i/9y9LbJCXUPR31PThMFxXiHAcB30GK1uhRpygl
ZJIDJVASERl3El5AYKxC3AO8SwQ4LZK0QlcTwp8o1NP5ps0INuxbN3er0yJETTq0
q5wj+zBmqPJqjY/J5kwdoO8bHx7ObKTDdO9khl9gpY06PUqNjKEMDEt1tUq/Snur
esEjYbzTKYCncqqbJZVLyoyOBgWMhV03eR/QdnTjmk1NIpH9Q2RUx2Yw8EXQngLj
Mnaefha1Gycetrm4rIgZsNcvE+OYHspMvnOf3GbJNW1PQYiLhfaOMi5iKsg1fy3i
SzyS2vG/FeMRltzqsaiLRQo2CEZwLC5ZVzQIO+z7AP0c0xv0OcUbHj4aMecJ2c62
mab8fNvG//GHwOcRPyvbI+Wjmnpv6DboJ3kv7dPy6621Z9oh0Pu/bF7CURBBES2j
2dqYOZAe+ywVLtyP9kmUMXq7tZ0sfrUsEsf/CdgcFwxCNckCtkLKm+n55kAKR/DB
pk4a8ucXeg6k3MaJRMxaxvA8gdzydou8my5Qi/sFm/SvxLIbZO/te8DUDwdtYyFv
Ly9TfxCPHNsUwpEst9LxepGUDJf+8Yj7fN7HPLlLVEMX113lYiucDf7Cv6zcrcMf
kDFkeY59Rehh5qThrJD/cBJi43dHaFsRBtzkmBMXryQqpzhaki/a+bStJhF6X1o6
Q/toIJHSbB8BdwrnNBqPbRlWqxK3ijgIdqepRJUhRlpd7lmhJGAl9nIY9M2r1wb1
K5PyoCmoAQ8Gy69+YG7xOCMko/xIpUHPzxDfe98DVolW2YQmtaZ2UhPzNBeLcs8z
/14Yu+AmhW4792gMDXuaFUsWFrjQEqmLHUW9dhvxzU1bWCYv1OJSE3R1zKuKGYeO
v0wTbcaitgqbEVTvHSxgggzutH65PqILb++6sK8LqsOQg+wdwWTXHUCDex6wYtly
lPgZBmzt95lQe96XAyLodAZRUbB2GXI9fcDVeV/m6jnUGo1dbnTkpZhlMggW8AKm
Ja3bd2KV0/npeJs6f6ysxvlvbON8Fxjo0A/sDlvWk/sZAi/M6hzn+1WJUU2gAXLI
uETWg5hn5+4nNubdvy9mGbsZcFFxjW3RoAQDX6wSuywZe10nIOgfyuQvtt391BgO
7h4WLSB63Vwm2EVra6uwPyHfv3JEvEhdgyBoi9IAL349A4hSLZRzvCBNWaD9PEQF
xKZuaqsBgfdoWlmoqcb7AB8/TDyHIPMgyj4NppsNblac5ZcFv/7NrwWYjyBxlm4e
X/5ZlKu7e0DLeC/MMtr5taASkziBLcdaMOmPCgKW7DwksR2DHLlF/t1iGtfaGyhy
4vl/STiJXvMKcmCdv4jgFygX511AgeIJW8sq7cA79HHEzb70Iu9QeysPgNrPc9cs
1vGvO/IS3YIMNJyo5udrPs3rEzFlJLEwZUGGUNZPdppaYOmYz5sK09kpQQtuW6Pk
9RDcQF8SLftjsT0o7rcJnMRkyNONUQgOatA/+1V9Copg7YDWsMlcym4Br4AIbU3e
j3AHscK4huRe/+GDforbD+oZsAYRRhrhgjKumLqwLD0uSjSRWidCJwBvGz2PZjwH
pIk0s2pRMDo4j3Bw2ZxhsLiDR6fxL1N9lo0XTxK4rA4FIWi7225JeYBXllHBSkVn
lwaWHOS67kNuf/BbYuBP1p44kA6FRlLnAb8oYBY92fdcbAQOBKkN+z2sfWF6EmuB
qBHRGnVVgIpCUQptAuOJhi72DhzLpYepruh/J3auV/Pj8VkWBa+1ylClwOaVk35S
NxaYV7bGbwGe9jBoxDbiVziydsDIUIHKP6nJACmpLTpoZPrXlcbBJuDeAWyl5WxK
GRk8hrkdr2QE4mc+2Zht8BkUUiwPOIAWOqbpBOu5Jjp3jezVJj29p5NC4rQpH6eY
Vu5Uc/5b67L8TF+KxS4/LextO5xK5rq0BERTayYxPT2OlFyo0saaDia/mQdB9phw
qNNpHj4x0O61mTmWsWkcOiFjHXxGmJGworUZ0mDrLbP4CPm81+GjvqIeZw6sFKTV
Lsp8ja22zKDNAHG9ZpmagdULGG4Fo+RUj7IYF9hC7Trne6YHPa0Sw1p4W0xTmjJA
VRbmSPnnIpt65IoZ7A29jG7eBO3zpV4YUs9A1VRG3rcDt4RED5nx+ZHO0Ry4XtOC
hZU8mReCpXZ64Cq85JZPIJ1K1XFcYlRnZuLqcHNDplm1E7jh+HXKJlHBzwdFLXBw
dCPUg/2Axp8umS3HYWJ1HzFkCeLa6o8nOYcYUlNswQvrlADO1xyPZuMdxAu/c+Oi
bm59DAllnBZ5gKPacgjmBpF5u2sZTLUYfoXlfIE58MuKExVBwdlQ2lKIjMr1msri
PfVHiBNLvGv3d7UkDV5HXygSrLCWAxTm1MDk8ubfRyCdNmbmAQ1CPDLYTMk7/Ekj
pCRd8amEjS6vuzY6YPc4BopFNINZoa9N5MSCmmE0P88K27taURHth4teOZ8LCGb0
mq4jccuci+M3omOczckfUTkXroZ8dW2BlsPaOeRhuv8twykYQS7iy/1pCMhpBqfc
uKXH/NvB6lW7ui8v8KfSe1OEfO0OKOcgSZs6V58waYeb7W7MEH7AS1qzMQOja3j0
Xt2uppkzzLZMRGCCfhf2Ndg2VhumnJ8OJehGTnHbwbyKm2CBfT7UIfbdn126sFzP
IJFJkeYta8LdlvVgV4OB5hjLCcscOGYUHEa30aiv7HkhNAsU2NRTDTZLa/niAQj9
WbadOgkYZx6FwCukhf9nOQC4Q6nvZ0fTyyr0mCNU53zyPVomZ8MeXtFrJ723O/xz
mkyPZnkqwTXGl8hYGtQNe1RRYEqhoVRU9aNSwmKEGPt30FVhagGbgHSipAgO8/fP
LH+rh6WYE6RuEzdYdCGLEgAqe5ymjySD/QRJaiTWSAA2s9RKuX8Ia/MBfvk1o4mR
CZiSOaS0ycGq3+L7w75WrUjd1CLeGmQ2uc5DsEGfI2PxNqXi501oSmgXNuPBvVLm
0IPMkwGZXJtyXqmoHw1DpkOtH4S+6LhMBcRlkb/iKoozmDEGUFdsL8vT5DJB4lf2
Yt8QVVUbW/1NK0UPVq3tyhyOo6pImHWU6jmCYjXTo9JlYBNzz58nHRCossXMZHzU
OKOnUZBvPDJxTLsny6GNHskiyg6hhMUktvRWy9Eb6G0ikZogF2a5IiaKn4hdie3W
5B2MuYXJDiRli6nVYtDadHScnT+XgJ9Jj0VrM44xly3u5TFr+AovKfa47wqdkOeS
8rIsFWAKSbLvjul1df3WII5l7TMrqvqo+X3/44LDu3EE1Ky9+/4ozRlQyIzVuRuN
6DXmgoCCW3JFAU7Qi9aIQcOU8IUFkGcmLrjx/XcNBOzS6VniMNnfonSEjv3CxVUK
jJ7avOFt5vTsgL6qCc4GyJX/sk29h2Y+yfuzDzwJAda+2X7a/bm9pzSZeWzH2XeR
xs3ymWDgkgMfi+d3A/c5EwpdvFmDalIZZgdD8Ts7kCgOCBtkqM1A3bDoFRrq7A+i
fUo4z96ZazGuSkx6hl7Xw7wAYYcp2v7AI1JcO9jxm/697tMnifF4uLoqlqHhXc6q
3IbgpylhN2T1GchLm8uK5kryPtsxg3v+ORJxhzEPFwv/UVwH0TY2UxZGx+DZjWy7
MoW5v7GdQ5i0thDWUpQ1nkyNOHA6sZcI4BtVEodTX8+9caTI8A5CGFe3k+Lb8+ZJ
qstO1uimVvCfYf3MIeCqTeJOJnAfKvkNHdj8N3hULOGU+9fDKiLTeQszjuf0dt6W
OG1eA1LvfbL4mxgRY+Y02mG4e7d2ViicYxQQaSd4VImrAivyvtXhocyvTqKr5TRO
KQdlTZnCqwGtGS9MYM6qmtDQbMtIzwSmRevtEWc8DskW8EHFTXJHtq+eHck77eRc
jdtI8HqWhXsIAONRpM1Giv5lwzkiJNMQ+M9rgBw31CxqRrJ7+epxd79cx3dYkxWn
S/A4hOBlylL0N6tfN14HYitafy1QbN1UWELhlaHzGPpc+fSJJjhKrU4TBa8eCmAu
ESdv6cM6ne6QuXNTMPKn5X2VVA9C6SKKWk5N2VaAShJFfCmFq5MChZ7wkPUVVERT
7lOVTstbSOBOz8cmaWIBrbu0JXxUwmgZj8bnKhHuDrKq34WJU7Js/FuFjBPfmS3s
Y24tCzDChLlt3N1UFgqkXrvnfYbwybxGuhvVvs3uDteqcxl3ies+rNjtIev8rWov
JQI0Vk90Gby6Mcqy/76q+Yf394Bd2I95k6Cy1AJP/OKZIzCzLdsQq/nI1IChdBM+
bPFEfUSNbgn54F+4eDIisaTRA7rdpMTmqh7kpZslYoc3lwOmHUjWxy+GZGk16ugx
aTbSd002uemwnEmzTBCl8+SBqvLou6M/KNhZCQnKlJJVoEJfN8mj6PGLXcx7Lhdz
iXSLKQWUtlK99sNA0HBL0zVJBRqWtMh+XiV72RAY/XI6OHltOXlFhQajlRUx9e2Q
MZTCEWfnR5NsIjYv0tQBiKTu5x7gUrT06lcsKYXavzj4iSVu1hGiNxgZ3a2wuvpR
K5TILWWRXuG/vyDCqvB3AMsvQ2zBsUhZcbno9KrJXI38XUX/cIrH0wbEYJXlMU8l
iUgEebW9caeOZeO5yniE876tToUqSrPYhP1x1FVhXHdBupyjVzkhnEsqViDRAh/J
avGzPpCUVlrjmckbK7NtcJC1nqTVCGAdkIpfhtQGwx0g0096KXEeE2AmDNjqkEGC
syln5dKgMyJ+KRuWJQSyuqPSBFy0KHy0GKMH7yI9St4bQQIYq9WlaXrXZLDYJA5k
I37vl5Kjj+ySJ4uhNF7DBnKhA7kQzX2TUJn9GtNAZVLvLPHeSAu4PBQ4/RrqD+kS
/V6Mcm83dqcgi9h75Lk7w9bPuUzQvtNWeFYQ9/Di7HGVSYBIr5KaU9khzboqokN8
Z4tNJn59VWHDYNKk60GHI9FfSJfb9sO5P1wZLOKIrIPbt7DH4hFgZ2kezX5ldBcL
s9lyBCOYuJ7T9iNoiI3y+zRw1s3I6oBj2YpYEQEIt5flmVRhn8KM4kFty2emqM7C
rg2PeoP4vRSk/YUiY5hCI/gxxmG5QW8JJBAK8jYw4/eBDdu0KGCJF52TXImNMOlW
Cm0+5RpITPZHO3nShhReDkG3L/P1auD8umjuNjJCgPGVQ39qYT6agyFJZ4qyIFJy
T1njaH3IeJAD0NajVmdijmJmtR9poueBLj3PN81Eh7HPbmNr2gK4N1LQMHL2ZzWA
9O++kaNGd2ZT8bcPgm8DG9pg00n1rrUEwMESfsCcuI37/4e4KC2vqUWdVvUEZ1ih
nylZVxGIunGH7F2MidpdtztnC7vaAKd6/kD9tOjOrfP5+uqgfuqXZe4/q10w329b
jZx12HS8fzS1c6lFy1ecNHpqfO50W7nw89RbqBV8qbcL3yCjRpjPXArnBWvpIyTZ
Mz0gjCNOoFWMSbvrSMD7BC2R64lDIBrZzp7G1WZcWpiSj7vHbCPtxXIbSOE34Zy8
+FNW6cSKRWx1lEwxrxY05/dGTL8M/8yU78quGt8a5p22Bm/CLzLpLtz0TgAmtzCz
TW+3u2VevVqYD0pVbDJ+uTX+5PxEFYg4m5K3nNYifD5kqVUxXyKAjWVDBzJR5M59
DCHNjuRA5wWHVFUuZ+FLAxjiAp48Q2ijScW/3vkzYfYtRsngplzr7eOwbWwy5dzd
0c4dzEISmkmYDpGxGGg1/yTcOOAP3kRodcOfUNPCAbYM4YQkBSvm891WX+tg0EhC
teL7/8lNOYObVwgM/ULGZtwnv/RVXlUBzuSN11z/9fpAfHACuuGh4me/JIEgHAJw
+I2fUi/cxQd8+Q8gGMEcnGGLOP9i5DrIYEMjfiDHZgyOM91S8nUfe8M/Ba6V2aru
4CWycZdqiwKuxkPwf/j9kmRJNuHR3Sku+0vQIagZahot9H59I1fUnSIlvPLBFr77
IPqZb2GChYXITEPNcCUlnlOFKl+EnpXELK8Xa3BpKhZYBEmlxYsxIcAsEksJigBK
Ce+XsyXnMkYPl+jMfYJRXT0hGBYJIh+ylQYinmozdULvOPZfYCgoyT2e7kAO45sE
jLWg5uxQAXc3bxd3U7PZ73rw83lC/u/0g3JGAqdCfHOAzfZ1jRDgJz7OT3xL9Mnk
TtEuiqj9FNgLSLBjtX/Y9YjMGUiOlvV/mZpWjhpSwdICtiP5tn8mRN+sWH9PtJC4
qGKafvF15d5TfoDTAmh7b8q5seGdV619y5Wymyql9HaTmRKaomzeXq7z22wsfPNH
9ZUE1qp17pR112bXefuVKsp+h0inIa4m5lrV7pVmU1BzHsa4YU3nitdEU8ezZaJi
rQ5oS97FWQr7ReDEiACwaZbYaVPpdnWX02+AfvcxViWsYJqJnyL/1GYapJvP549Z
2g1Nw6loVZ49lM9Ki2kKMVkzx7MNhIAUmPYbwSVdJNYXIgU8HWdjJzDoDBOWA4S7
LH9RxWijWCk0+2mMQFh8VznEaSrSOTWfC15DfjxrY+Ae+9Ncl+Nn2pXQrkjnb0mL
Zkypm3xXVKxjFf1BEPWAV0gUnmSPK2Tr80m/ciEwdcAVfeg++XR6wQa4IEPYGloD
csFVnaZKXYFFRhOZyTsTMmJuUNs9WU5DcD/4cDZGrxheG6QXkM8WmsSFCHEgI+LH
4TD1vOTJBeE46c25cbvRET/dITzmKZrm0/gyGPRWgntV6IEfGYFJ2TUXvdXKFkfU
qBN/j4ywGx4n6dsIu+3M7libOkR33/cZKXU0a0IXGqmrUgppEGYzWsfAYBrb4Lv8
kBRsvCXcv+uTuPj6sFlWWjXCiY6yAEzGrOUFU534hVsnCH1O4C5sFMEP8Kb7axY0
nLjsHziWDwT9qbb2Cy2BGLIHeGXSmESyR1kYKlgN+/GsQw1H0Vy2OebpK6eEwBxT
Aip7jXOZgNv30yWQuuuAaiGZ6RDqHypG9FaDsTKKzuOwp9npyYU9Bevys7KdSjZ8
ryu4r04hjfep+eUVr5LkiROESUQOfPJDhji0xWMtBEAH++GuGrs+KKBXFKG1rRhk
WrhAlVcpSDOkWCr0k7shKxE2g0x4F4d1dB9bUO9MWV6X4AGI97yhwYmigsYELBtK
0BowTbkLPWpRBdkKFhfKAA4vk1t6yfx+LCSLuKnLzEc8VBrNTfcO06+tXhTJQY9f
jIA+IgWD+3G5VCvXQKJqfZenw8GoQdalmpeS7QO/3HAcBaUPskC5J/ypQxjybwFQ
lc06uC6YJCVpv8qTYPX7hv89Wd4BGE3UX21DvlvEWlZHF5nHhV0xCMIVMCaUwqvB
tqlRj4hN7rFDqts0s8spiAaTDVpEqi2JqgIqapn5wxWfZIxipq5xAm0jIVk01m6U
mvD3IyJ+wNmnUpi1itWCTnVlk9QsXxmzk++3lXUbUD2sKwFvsAramXfXxSJ//y8C
1MQ9nFNLWT9g6RE5XaOII+csZafSNgxIPq3ZIwAYJ+NEJ9dJLbdfddGQp7931tBR
5uLMbDYTJQ/9/0UCqTyvulr3YEiBzLOgc8V75gM9uZa3R65naDzaUMKfVaZv5nW3
HlTZ+wF/gWboCxMonhZPAejIL4WubjECKlvXs4LH3FZd4cs0Us1EfXcpvFFgffE5
+yd5LF6LZUZeFFvhTHKuNhqCekF016NWLVKUqWeUmF4g9yKBgCYx/OKCvannFVyE
x0G9ntvmRKS0+erP8tKhpaPdopHqd40fg4bqcBl09UmeXTj0XCPIwJ45iZww3mI5
lyUvalXkL82Xzh1XL8HW+YG0xzpWWkMW1j960hNDtcf85e7sxmXruuEojYvvhOlj
HOLqmtgDIQlBTXK6pwjpJKxdOzH1K3DF/o/LKZCkH7HVJ4E330Xv3j7A9x/HKa2O
hKLwdUvPXwmUdBDqbrlqmmgCtaRhkEnUe/kydHDbxdxcDGABYEuyOk3VLQDCOIgT
aZlp9XMpwcMdUtWwChZyEQ==
`pragma protect end_protected
