// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
RV4LcmooABJWqA2IrkkemH85bHJl6O+TO8pNwjhSfeGkvxxqkpFyCVIsq/8fCh+9qeceCnxFMM3n
mb97JSeNRhQ0FpLimPhMeHQdrL2o3hA2itK5LOA4rewHyMwkhbOLXYFUXCXhDArD+CIq3Y7hdpc/
f8tmuvsbPkJv4T91gLe1LM1qxOKcs13aewyylspYEvF9a8MlmXHft3Cm3ivoAho6PbSJPMkMhECj
gZXR0tfhaCcWCS+5N6ub3ZBmNVMveNleYndEuse6RxS0DXlH/PpjmMEeo/BiVJkLVP4NydhIFITR
n6NZJM81BNqabPMWZ50bciQA+tmAQYXJYG9EGg==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
sH8CFw/5fG2tlxRM/6wZwfOKSJ2A8qWr9BYP5YVm5RrdmiLrDJXi6b5TWM+3S/JaXTMpWEcP9IO9
zn9uLhFYHKPcxlq+8El5mTV31gQ+t79dybbEe4oz9GiFG1rfCqz2uVz/MOEOtnQ4AnzgzPZluTDE
BQR1IFcVXYUfY6VjwWktuOzdMmVAXR9Svrc7PZPiL2tKek/vEmnmoBJkUqSDY62vnxEOuP4S0/iH
j7wpbhdi0qE18xgbPmAGUWh2ZRPVCKZE0RXh1NgWNUSLj2GyLH0RjwVqScazPRainlRfZxCPuDUW
BGYirgEZdiZiaDLq6JTQbwcrbjMqTNuWVu0nlaB8896l34kYsx2X9c2vlnrYYClk9vmsEh7BNI+0
wLgaKxYIDjgpgSceZnKeBt5BfyPNnfAA5F+m1LnsmG24l30wPWJKTCVHOD4qG8slPevGwxD18vck
yMj9czfEufWuX/D8U8kuEfQxywNfAB9Gd9gkAq7TyTg1lwD4rX2VmwAulHaYhPk20WpdbEgX+0FE
rtuBHz5WMN5YflWDS2ziLXKeenTz3UkaNA8P/TmHZlqa2I4molGVSJsFH018+ItM83YNp7l2Pwx0
ra+SeWZKwIMDIV+7U7jUwguYCh0gMg7hBOIy3v7w276rmw8Tq2hsw3uu6oz1JuMNt7v6EtmFQwBP
azVPslThgGUA23dmWy5tvhnV9QD2xghnBOFm4xbFRE2Wk0TAzzOiRIW+axw/xp7+Iisf4OyoSYaQ
bWqWVKZjQ06ZJhL6UfREu4Fv3XDLlQVI+ERlofOxJuedPW8fUljIpsgPnBTO9uhqNZIC8Xry+oIP
i+dFpBAZ8BSjYrNX6K5fkzsYfokiKm1l6fZCA7tiWbuYpSSb/QjgNc3/xYIALw5MeER7BHdrqQAz
DwPF2wzj8qn/S5nEzJ8arEv6eg7RtNGXXgZQRBwSkjOuv/vlKL09nmh6v/ScoPiJYDHbsBBvNSKQ
zr5fZ7Z2b4EU3G7JDQZCBhF/qPeXd4Ji4vrfQuYknKJ9se9xURhVbg5RzvBDSen39FI2cae0S7zU
lbcCpVZsn4dJ3FJWljXLElrtrqLtxIVBjau/uSj6X6Ubir8E5SXP8OyWckgcLrvQMP/kB+sT2wbR
V/z/00Hesj2WDOu7+kYOChqeONGyJKpMV4MYs7bpzvusEsSEgo6qOyyGyqOf19fyqT3WbF98pfnQ
GJRt92qN0waRK6xDaxDqdqGC2Rng71bjtvzwlp/X1Jxz6RntJIASAbI/OyRh3OLoS5x7ViFvGLvK
JN/6XIsBE7TxbtvpSinWKRqoEKBfFhKTBIZEQtWBKaHcq4gdHYy+MCnd0Q9w9fB/9W1gFMpGD0zG
XKnY/b7+KjNKMQzQE8G/TMWKjk1rXu0O4YZTDmPCZbP7Sf8SvfOcj/ZqUaua1KlpXo5qCd5E8ja8
RUiqon92vvOCsefY7Q3WVf8qgAIz3TRRb38u2hBSJ0bfY9vC8CfgJLN2q763+V+UA55AIc9mku5G
USLZPQCwick7B+YqDBGG1scKeL40iiYJtn8pFbwcSAZe9YHL69lQ4R3w8Rlj8PAbk9vtXzbXqO2h
eDTg8ZigDbI0Ae9MeNDni+1GUcm/QS7hAeveuKROCAH5fl3ONJcHPVvc+hevroi3BA+ZyhDgIYYr
Deu1hoMr+sf4/BvbqFDY/s05qcbyVE2X6NPwFjYW7zwNBIoyQn3A385IQabeUBIzmU0R7XEB6Zcq
fJ3fROXRuqZAG9pPm23d0AISuGWxG6YTEG6SfUnM+CRH9oiiSJE7wNm/tydZpnKEX6NSJRbQAOkb
MZnRWSj/wrU8RdIlPublR60mIycyTplNTP2G2aoBLWvApsq/TiKANNq5Ce2OueXwfufsG4L1Fjyn
8DLgJc6RYySCzEucr3GZRRJCaAdlzrTZMYD6ry2QcNvGv+lBLgr63d9KjyLNLw0IHsSV9TxcLLSA
hZsq6+nD4RK2SRDDYQbE6wAJunJkHJC1FGZ5ZP/wfDN5aDs3rViKdh/1B4ENqX1/rYZi75jYg940
3A4vZ7qA31BJ/QCqtgn3Ewr3TY6wC/ydnIk/9+8xErEK6HfGj7dst99kObKkqklO/rKEGZ0mK6Pb
CtdPkOa+3yPZYiyPRqSS8Qytk4oWo6a/M95agcSwiJi80xFGLbmOnqRYgR9Mkw+Y5p0vhrKxASB/
yYhdy901QEICUXk0zJxyq44RPhG7HNO7J4MBTxgOE6GFI/wKdQg2FknqyK2iq1j6WxVO8/3btz00
Zq5cHVdA8v9pztz2/7c624v4wlQzm4t6Dn3ML7AIkfQkZtFwOrmZfSGqPEEGFeOlnKHu0UQWv0BR
+sZUvv4XRperSYWnQuD+yge+cYQ5cI1vxlNSrzPvus81LZMLN/StTCiZMmi+mMsrn3vD4yhKAQfS
LiMl+EO73whQWskqLXdj5ZCobm1ajpKrDhrNtO96kp+nnemcmnLApnulfQ3lWLvpRgRjpEF1djKX
UuepVT3nmXf0Pex83dKmwwAm1eonK4SnbEnWK1/C0NLNIlXN7iJXmoSomwU00Xp1gCW5ow4KjB80
dlJDg4D3AvOZI/qQ4N996aY1eMurmE6QIoMGAg/NH2MgQfiK9hveW0gNsub9IvrqpEXrc25RvIkt
uSryptIZy6q0LZ3ad6avLzjpLAnpvbGwK27Z2BpePid44Y7bwDUkLVbGAx9UnmCSvc313sIXns0K
zowOBIf2k1tEZAMFzgG8hLoiaaYPvO/BveV+LRlAbeI9EjKy/szEpKt9KW7swsRkuVI/QCvsIly6
lsfFlnsQE3jJgBGXINxFmkZtzl7BRQ7BU4aMZmfsYw0k95opdbuQd2SKSyJFPnWXZOmA9UZ2CBT9
FOd8JMHS6oGEJ02WtfYFi+nDtXS95pjjnSqc2a4BADRClosuIuU/Yu7mxYaRg0LsBJLAFD53pdlf
+CmOOiZpLX69QGo3SSgLqN92xYWEh41Mu3m0iam1CsW+hQESVE3oRP4IatvKfrsmUGMrOE245pCZ
8eB6al0Jge43nuziB77ua7TRIPjYeSq3lGItpk92SU+QFdKC/Z6J+Lhpwcg85np97clRu91RNA+T
y/ttZyLgjLqrmMRlw6TsxlXrOVwHxm2iufLiAiN9ZdKSPvyNHLUTOIeqDMbsBrAue6rORtB8zeOJ
xBd4Xp4oj98/OeS8mWDqQMDOZgYTvAazkNXdzbDMNCDCslkC+Rp4OSsOfsswKWy+0z3ASggx2duo
FnlIRGBNwrg/vxOASJY3HzGx2oQSyDndqy1IDO5Hl0JqU1iWy0707dzuhzrsVibwOQKgYlSWu+oi
RhF4e4bdHhWv4kq5GdUBUVh0oJpqCyej/GG2tOSq6OFltSUfFT2hUwz2Ts3FdD484mBx7WawhPpc
Hj+CBEE7wFfCY/I6dhMZ6EUFitZaEDgxPYqpPO2dZvTNVpuSa6QdHQCa3J0u6rWoV9eYno55i1Vo
lUGQ0ljBlhT1g2XX3t2XO/yjIs9nJLW/i/b1/wT97lSYOKvqA522eOeyEe25F5yKIQN+JAYiO0zr
2ryuQeoOfpwAQeSiFOA4ZMKTUikcMZBAS1cx9xGrThFwAI69zIAEPWOab++28Axs+r3w9l40d2N8
P4WF9HmKjoGG7XAgbqR79lgVd6GWFIhEdakgnEd5A0s1kLR/uPvAludcYts4sFXr3NVnja63r/3N
ItKgmtzEaUrdn00AaycFFeAo2fRQBPR/2k+GJIIpePO0qUYywKCGM/ANRjIk/lCU47v5cTFAN6MF
/UkyzcWxGxKg1DAM/34e9OY7Jw1ceJtFpZLhG4tGwD5+P35DGEvzLao54JdHwdJdU4L2fONyTNfI
kgov4I1e0Kt4AJeupYE3tBp3uU9xfc48NiRB2PxPwjO0jRjpY5agjW/2B4tiaCcbGBiG/nKr56Dv
QZCNasEXQ86xS+60BYbidogwLr5ZDYm0PwmbjLUUVajMnKpR05z3tQKUJ7iVXS3El2qWU0/6dL+W
E15jh9M73v4Hpme8WTDgYRUk+tQxP+UmLdM3XMkAbDc9dETYBo0ncfOpVPU3C+h9DiPB7LONKpH7
NvP/zOnsrVXov37mPFNj7VqYunSQrVuburKWUblzBod+TODC2+bLpHXG1mKiAt/FIacQPUtDX41q
7yOPDIu2zBExQGGCzsc6rVahdm4wFogJvu9b3iwXkDAngdtfGPjJ+3TcoJn+mYFf0QM0EwXTlCri
E1hUIE+blzm4LsNUjroxjY/SjGuPafAQ/5YYqFS768XV1kkBcN8feMFhqd0AhRuo3WPCFJkXfWxB
YKwzzKjHvGaN9Kt3BMIC1oIG8CQMwqCSTCFO+VqcQPsIn8QYBavvwKLCcHo1C2TJaguFiUG80JZ8
tXqQkzVaBSPS+uZVD2yHgayVdO2D6SVTVxt/tBFiosw4e936ifxKaZZ5q+hdPubwnNGzclsQ7qym
ljMEWNko+EyQE9X97GUKi7Wqp7I5U3zr3AEfJwkDvOL8dGrY1yAGjt95ToeeLNa4dmIXFclTVEJc
lUsRTmuZC6jcU0cCiORmfyiZtNR2KHO8okQlStBLFgajQgYdrJKHx5t5vqSdjd5XE0HWkeqne0eA
MxDTSIYneIQU4MQlDLoZAsnat2Mmyq6OrWFKT1zHWo9O1jvT9Vg1bVFps2kU/UehYFg98zNhNwLz
dZmbbSCWe1qChGIv5ENbYRXKT7vIQL66SNymTjvzX/mQK8juZ5Xw75MRFGqALsxshuHbcAcWuCgg
7c6dv6+b9toPqNwFCoXUrdRMEFLjD3/Y5KVamU6MX/b3pfDlGtDJIvMGO+lo9IOYLK2i7uigSVhY
we2A+ALS+ThXO4AgY8qiNGX7QviTv9sZzyUvQvqnEfQxbyHMVxa6JuS0bdvT+lvWVPVsXURrA567
9uJUDPPrL05fmtwtY7gzHmIgHLQOi9LKtTFq0fEi051B522ybWRbL4YCn5IS1bJHG4VkC+vhj4E1
bZUfUxy4V/hiDE2/k6XWuk86w8UgCF5rEssnF4iCOk4lTEwI+9CeiZ4TO8OytTOFNdpSitUA32lZ
hNTxcEv7IG3aewLUxRIxmlMAPz0ovjgco6DVh0Yj8zBDHjiMclvZ6ziuE9TGCStPfCis6BuS0XX9
TxSn1OHyKjxKo8ePYSCQNhAqfs1sm25/YarUvCNp4juzFsMvgxA15HVceZLHBRqE8fRQGL09D8GU
JjbJX/h1uRF0PU/jzRdPlEQA7LpYCKRamsz6tsfkcibRFcVRxlzQsc4jh2sNOTTPizEcWa+ACQHG
tyTg6rp9XcZcFgSzA9R7GHUre+371lIuE8CyRVw17QDDlTAhDmNGo3SsIx78fONeuhDY6NfkBePP
JyzLBSpbUbaWIIjqBMH7P5rek0dG0tsi5/lK6s3WkbZ1VuTTGiLl3CzKhZzAxnxnCt175fDV7hrw
Tjm5j5bDABrMV6SnF+ikbPCeWUiIbr5AyoNdCA8ZzcKI9CKghSL4+nUudKET36F2prDbEngEkbXp
Hbsn+m39+15AmDJo6XsF7PgBiIhACMA6H7HX2D85Q3E3B7wvZP80kemxgBaBWCaPbeplHTY8q8Jd
Hp5AEuzi5irzY3JTo39RlkA1YrPRG6S1mrGYNI8BpRk8HZfEv81AcdybZ17m+jBSBOVVagvoQXfb
u2iOme8Ot2RkIC7sHpph6vBD2fAtJGO3vwLJMeTTXhUhBCZWWhVxUFANkPLAYWOmoFs6PY1IYzFf
AK0YCVILx8kBYT5No8TpbOyU8x5hKuZ+hdJEeOmS7k7otwSm3oSoqTpCSh2usQ3r9IqtensWe+vt
x2G8LEhmsaT36OxtEIpv3rC9pzXGzywqbPc13Ep9sWVQOhSchd2VXP329IcWdpUQXWni4YEqjlR5
3n2+G/DXXlrZhacWnVwKxSl3x1y5PolJFY+80SnvqppkX2Ic+jF/kw9GWB5gc3AoZYWjqgNRjbmJ
TMx0SQz7Wu1sa3rvVJf6JGbw5biPwpE2gBmZXiHJddDQ9goGZU/ha/oBonHs3JpOOJMYbMzBo6vZ
2/BoED+bwUbe33WAlKh+So93MUzGyGsZesgybv9OiFvTR2pUXLlu2CoRy9HM5QC3EZLscajTJhrQ
T6H/Lz5o/1Ned3KrQc/hORZYcysRe2kXG4zkBMJU4yZmtDnVVETxUhKX4Qcat9dCUldEQLU1VUso
3WdLsQHWthVZH8SZVghJ1kpDFnJzS8Mm4BVWbWo3Cw/8ybEyeodGJdJSe97nVfPSdgEnEbIkvsFT
AY4HPBxTb9tnAm5R0ap/EXkx/z9o/0RBnrO5SfdrT9s05HZconlXxzlsK/tt3e8L6aQFOzLVPb9Z
6TXrQvdtG0Dox+1XG8bsH671+WV4h4xfmEkqOpx55FRXjh8kHj3eywzSRnYqIaauge350zQNf/Gt
WojrEuyI8Dcw11cguvV27KBeFaF9HbRgiDTKbNZRWjLLXIFHT3/4Z4yKt0b//YG+RK7CWReLO0GN
9hqoHouhcYqNfKELZvCQYf86W33V/cDdjkgUJCTvFeqY6HcyPM71A0WkrTvg8/corPoh+ZnXE4t5
82tcxaLH5LEYLjHLxzpMsQFwQyaHSI6yp4lc4GtBkvxblYrkSptGfg91+r8ivM/ml6FkCi/FY2G9
9xz5QJzWLr+GRI+6woDy8iJzgYSdJL9em3hHLmzF9sGF0xSPpLaDOY7MVrmJVgqHiKc58xCmMjgw
WkXJ40EzY5ElSRmlrN7H0bmATa8uERUVSjaKzdvpntkp+8pPGx4pF7rDbkj+osS6lCGti4nisv6W
cXlWItfxjdnO4/Ji38bRe81OaxyQJyMTUs6jxBExZfLrMs7Jqiug7FAFa6dPDxjsbvCkaxXDe/7w
4d1WK0Pak+5wIFIXxMUwa7+CT0elFpFNmDTFictFa0G3OG3jbFAc1cjccFfF396czh2fCZxGcJU1
OACLMlH3Hb1cRYOWhAkNPFU0CinYFGQP640GCqi7UB1fUn0+1NrfFn1fafr/KQbLT/x5EWnDmKz6
H+zTiQk4bwFtUeJ3a4QrrG8fhrbOE4zqKMUKGiHrem13UfCZoB8EAzouTCtbjvFe3ibu+EbOGfhk
wP1727y+osKBY3VFnLwj0iwiNHiK71zEdmkAHzOZlfj0lRwOVs6Rd+8jnIRAQsSfqR5ogSyvkgNL
lA7aJIqZ14nTxOlSgcW4FwkSdYrntOx3cOhiiSQZUTsDYWYIfZnWahZn7DmnVmgqOcjU9YFKga96
tDhLfkBzGLwUwzYRRi6U9wCWhmgsTJFYzdc87TPFMGi2fJWRRhMowIxEzujBldoxaGItQiJI9yxP
ZAY3GEYF6cJrVO7oE0BNUOmKHDGALv0LEeN+EvirJptbza6VkOEIBPm7lC6iI1ZeiJOeFTeaMz7v
EDMfl8MurxNaoj8DQ4IEb+pjZc4qYvWRJx3y4TCfRFSJEo3ZAK6NBE4eFcqH5l4VQYDPHfkmSw/z
dqq12v+16PpvYk9Xt9lORThUCWwI19TEojBL4zrdQdr7BjaT4R9O5sCBgNnefzhSxChrDQFpPLGF
Sfb6bnH1hsyB5UitSLeeFjcq4K9/YUXP4kovYsXS3sQzIJM8BhhAp6hbIA0OucitHtW/PF/Gpelm
wXL1zLdhulNpYFV23I0Ow1ssWlVNtO4UsDtQRhDgcNKwWoK6uRsfRh62M56HHiDl7ioTs8lI275f
9Avgud1GT2oFv0PrlCe4NsjsWHXWeFfwZ8ZbSkOcUyYpCgjvgGULRnaeSVyyzThGwJ9FfxP5lgpg
+G3y6tOTh744HG2sfpzKFgxN8IUpuusHqr/ur0aybmBEqqqFmeCvoiitsNGVft0E1RhatuIA3u8e
Uco3N4nhCH3cCX3trekWU5wUgrKpCigrUGOC2NgYxOai8SBFCqu2+RacDCMvUwGOzHfrRYQQDm0y
50RaPtnE8oKqDXlJhbbCbSpayTdqh2vZAR6aGZ/BVR6QajExDXiFpSKaHMzfKA7J7K+Revqhc/Cf
loT1KHZPb8GN61Mli9bNg19hJfp/gbaNmxXdtejNyqM7zAanLWdaJqWgDW6aGodrg+I6tjQymW3s
7FNHXhPKjcsD9hMiDOjAqqDVxWFNCU8kT4c+WWs0AgX/AXSAUkdawXd4ixOEIjBetY5QEKTRGC7f
XYGjao7Q5XKNiVZHy1eI0Of7GBSpdJKdKYtaDhQsRDoZ8uJrtjsk6Zr5qS2KeQbCPmycAqwLQTF4
vBEnI9eYKwjRLtgfGMvTmDgVyWQJ7MU9rK5GpHdHUOgLcT8YX4r8jmICKTuaRl9QPOl+9E/Rz/1E
TvIoLyZe7rf3Ry0zk9dLSec8/COk6PQGh4G04rymNBHVpYD9/z4hiRycSXZy/mlAaSwDBCSyqe9W
bHospO1lEYzaTdogoEFfdba7NKWtQuO07FH2e2scE24/Kzu4TAwHA8O4aADqdgYM97d3vZn6uB9U
/nrieqjqAfLv3vZmlAI4EdvfUcvMAOWCJPd4ZWwAS1PUP2mK1Jl8yHxVMlC/4fjg9NdHtRulRtQe
Wv39oTqxuSkzud92e2ScA7EKp5gx+JoZTMkxb4/132b/ZBrJcU8vLHfxMtwpFPCB8I0jjNGSopXP
deVsOhB9inqZ/OLXc7WMQzKD3zBQoUs9lhGZHd3JODVSY3IZJNtnpasAlAkkkYlLAw8HHp0ZaNWD
AfBb1xs9xYbJ7ypRNx1lQ4zSA9pkzucivz9+GESwfjFi9FXSDHIZTj9bSVZFVB+KsC58JTfMH/y6
vvFhCP68DPM0IIP06dbixzvs/WdUW/8rOX5WMqUyX9GqoxaVJwhl+xe34jon4Bvkfruadeq+1oyp
wNxWJ2XZtOQi47YulxRH1Oh2QX3eAJomVJVFiiwpCV5lqgVXA1n9yyUu2XN0yvvvaGpLl+piOoKf
WEXdlwG7nGcUMeqveJHPf9OI6urXetRS/iLQdcSDw7enFJgcI4dmIm1FJxjs3Tedq8vb2pn3kIeO
3xBS0uaRl53wxuQMwFJQpMbqdCucFK69JjBuY4LrTj3ZEiMGo+lRLclkY5vl20VnrFTSBO+R/vjo
vGrny6+f6vFuvfVvM2eqQmnbRlD3ZCGFcXw4/VTLwAZMga45VI1fYNz5flqiXvk7uLnDf7mvq50/
lWP1b+fSxEgXbbfaf5NlCdSm3mkzxhv5fHIW6c7j0ysFvzIydVqJYVcKAnnBT9zm/9YXGO/KFqvg
MGm3fWuKBChK1Nll1LrreIiMIHMRLeTm+lW6XzWM/eK1TmpNhqB4UpYjIFArjwVLGuO33NjeLLdE
FnBrKAbMCNzCCduFpBpuASIJf2dD/usOAnsV+6OxC37Psgb/oPiZ1K5gFIECCJoj6D6M6pSXZC0Z
jwdi0Yg/tFqBXXzgTL9FV0T2Z5w8vYQKYqCY3JnAt1qLoX3HNujYoFIhFpOTxRWjGaBhfAFccb4c
gt7vhTyGtot1d/5jF0+/Ri3SS2/EyH165igfOgYZ6ClgHS8hg08vWlPB+iL1XhebApgtMVMGPDa/
ZOFAnFsgFUbmRWN/U3KRZw5lwoNcQkZgoQIB9zprr9XYCz1Wk/Em1XhPGt5XVtO2jwCYXgkm+X4+
5qwdJMePSPJ3pBqWlw9rgXWYLT4V8IeqjF/gx+TfhUYoA+RLgQPWfTHt/r3BudlMIPBr5i91mQQ1
UYR4dL+VzJByoE0OVcFAy0DqUu+1KzdOrV/GX8rRiD1V5yH2YG6IOzK2Nen6qXNDbVg+UohOMGIp
hb1AUKZj+QJMrI3NIRj/bP6sOW+Z0f2rTEX/K9FgVJEhcdBux2+0Y9XHqUy8tQXRxxEEEX9tHOfx
w40P2ldyf6zuMvpTQPQptis8a6Q9MIZjBiti2FzQjVjA0cR+5GKXT85yWg2B4G1Ich2tgkLSbx5u
JJWRr5HxqrxGdjjmXFOnWuwNBKQniNFPxDsq39dqDEquKlxXNoovhiMXbBiZvXhfGgFWbly5TazO
ZR9oZkLQ35/qFBvmJJCwFEUjpepNLae2fh07fELnJRmE+1TXTfk9N1U8tQYr0x/Ef60UMPN/C5+7
9Pns7TcoGKw0LXNtyodAiT3Pab8dXlExQ4kYydZ1b3R1C5K3RvWQ7I4v1jlA+/eq7RsAahr9k4Ov
jiadKtUQWhBXgA==
`pragma protect end_protected
