// (C) 2001-2013 Altera Corporation. All rights reserved.
// Your use of Altera Corporation's design tools, logic functions and other 
// software and tools, and its AMPP partner logic functions, and any output 
// files any of the foregoing (including device programming or simulation 
// files), and any associated documentation or information are expressly subject 
// to the terms and conditions of the Altera Program License Subscription 
// Agreement, Altera MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your use is for the 
// sole purpose of programming logic devices manufactured by Altera and sold by 
// Altera or its authorized distributors.  Please refer to the applicable 
// agreement for further details.



`timescale 1 ps / 1 ps

module frb_timing_pattern_ram (
  CLK,
  SSR,
  ADDRA,
  EN,
  WEA,
  DIA,
  DIPA,
  DOA,
  DOPA,
  ADDRB,
  DOB,
  DOPB);

  parameter INIT_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INIT_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INIT_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INIT_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INIT_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INIT_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INIT_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INIT_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INIT_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INIT_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INIT_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INIT_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INIT_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INIT_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INIT_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INIT_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INIT_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INIT_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INIT_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INIT_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INIT_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INIT_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INIT_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INIT_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INIT_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INIT_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INIT_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INIT_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INIT_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INIT_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INIT_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INIT_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INIT_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INIT_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INIT_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INIT_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INIT_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INIT_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INIT_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INIT_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INITP_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INITP_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INITP_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INITP_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INITP_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INITP_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INITP_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  parameter INITP_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;

  input CLK;
  input SSR;
  input [8:0] ADDRA;
  input EN;
  input WEA;
  input [31:0] DIA;
  input [3:0] DIPA;
  output [31:0] DOA;
  wire [31:0] DOA;
  output [3:0] DOPA;
  wire [3:0] DOPA;
  input [8:0] ADDRB;
  output [31:0] DOB;
  wire [31:0] DOB;
  output [3:0] DOPB;
  wire [3:0] DOPB;

  reg [35:0] RAM [511:0];
  reg [35:0] RDATAA;
  reg [35:0] RDATAB;

//------------------------------------------------------------------------------
//MODULE BODY
//------------------------------------------------------------------------------

  initial
  begin
    RAM[0  ] <=  {INITP_00  [   3 :    0 ] , INIT_00 [ 31  :  0   ]};
    RAM[1  ] <=  {INITP_00  [   7 :    4 ] , INIT_00 [ 63  :  32  ]};
    RAM[2  ] <=  {INITP_00  [  11 :    8 ] , INIT_00 [ 95  :  64  ]};
    RAM[3  ] <=  {INITP_00  [  15 :   12 ] , INIT_00 [ 127 :  96  ]};
    RAM[4  ] <=  {INITP_00  [  19 :   16 ] , INIT_00 [ 159 :  128 ]};
    RAM[5  ] <=  {INITP_00  [  23 :   20 ] , INIT_00 [ 191 :  160 ]};
    RAM[6  ] <=  {INITP_00  [  27 :   24 ] , INIT_00 [ 223 :  192 ]};
    RAM[7  ] <=  {INITP_00  [  31 :   28 ] , INIT_00 [ 255 :  224 ]};
    RAM[8  ] <=  {INITP_00  [  35 :   32 ] , INIT_01 [ 31  :  0   ]};
    RAM[9  ] <=  {INITP_00  [  39 :   36 ] , INIT_01 [ 63  :  32  ]};
    RAM[10 ] <=  {INITP_00  [  43 :   40 ] , INIT_01 [ 95  :  64  ]};
    RAM[11 ] <=  {INITP_00  [  47 :   44 ] , INIT_01 [ 127 :  96  ]};
    RAM[12 ] <=  {INITP_00  [  51 :   48 ] , INIT_01 [ 159 :  128 ]};
    RAM[13 ] <=  {INITP_00  [  55 :   52 ] , INIT_01 [ 191 :  160 ]};
    RAM[14 ] <=  {INITP_00  [  59 :   56 ] , INIT_01 [ 223 :  192 ]};
    RAM[15 ] <=  {INITP_00  [  63 :   60 ] , INIT_01 [ 255 :  224 ]};
    RAM[16 ] <=  {INITP_00  [  67 :   64 ] , INIT_02 [ 31  :  0   ]};
    RAM[17 ] <=  {INITP_00  [  71 :   68 ] , INIT_02 [ 63  :  32  ]};
    RAM[18 ] <=  {INITP_00  [  75 :   72 ] , INIT_02 [ 95  :  64  ]};
    RAM[19 ] <=  {INITP_00  [  79 :   76 ] , INIT_02 [ 127 :  96  ]};
    RAM[20 ] <=  {INITP_00  [  83 :   80 ] , INIT_02 [ 159 :  128 ]};
    RAM[21 ] <=  {INITP_00  [  87 :   84 ] , INIT_02 [ 191 :  160 ]};
    RAM[22 ] <=  {INITP_00  [  91 :   88 ] , INIT_02 [ 223 :  192 ]};
    RAM[23 ] <=  {INITP_00  [  95 :   92 ] , INIT_02 [ 255 :  224 ]};
    RAM[24 ] <=  {INITP_00  [  99 :   96 ] , INIT_03 [ 31  :  0   ]};
    RAM[25 ] <=  {INITP_00  [ 103 :  100 ] , INIT_03 [ 63  :  32  ]};
    RAM[26 ] <=  {INITP_00  [ 107 :  104 ] , INIT_03 [ 95  :  64  ]};
    RAM[27 ] <=  {INITP_00  [ 111 :  108 ] , INIT_03 [ 127 :  96  ]};
    RAM[28 ] <=  {INITP_00  [ 115 :  112 ] , INIT_03 [ 159 :  128 ]};
    RAM[29 ] <=  {INITP_00  [ 119 :  116 ] , INIT_03 [ 191 :  160 ]};
    RAM[30 ] <=  {INITP_00  [ 123 :  120 ] , INIT_03 [ 223 :  192 ]};
    RAM[31 ] <=  {INITP_00  [ 127 :  124 ] , INIT_03 [ 255 :  224 ]};
    RAM[32 ] <=  {INITP_00  [ 131 :  128 ] , INIT_04 [ 31  :  0   ]};
    RAM[33 ] <=  {INITP_00  [ 135 :  132 ] , INIT_04 [ 63  :  32  ]};
    RAM[34 ] <=  {INITP_00  [ 139 :  136 ] , INIT_04 [ 95  :  64  ]};
    RAM[35 ] <=  {INITP_00  [ 143 :  140 ] , INIT_04 [ 127 :  96  ]};
    RAM[36 ] <=  {INITP_00  [ 147 :  144 ] , INIT_04 [ 159 :  128 ]};
    RAM[37 ] <=  {INITP_00  [ 151 :  148 ] , INIT_04 [ 191 :  160 ]};
    RAM[38 ] <=  {INITP_00  [ 155 :  152 ] , INIT_04 [ 223 :  192 ]};
    RAM[39 ] <=  {INITP_00  [ 159 :  156 ] , INIT_04 [ 255 :  224 ]};
    RAM[40 ] <=  {INITP_00  [ 163 :  160 ] , INIT_05 [ 31  :  0   ]};
    RAM[41 ] <=  {INITP_00  [ 167 :  164 ] , INIT_05 [ 63  :  32  ]};
    RAM[42 ] <=  {INITP_00  [ 171 :  168 ] , INIT_05 [ 95  :  64  ]};
    RAM[43 ] <=  {INITP_00  [ 175 :  172 ] , INIT_05 [ 127 :  96  ]};
    RAM[44 ] <=  {INITP_00  [ 179 :  176 ] , INIT_05 [ 159 :  128 ]};
    RAM[45 ] <=  {INITP_00  [ 183 :  180 ] , INIT_05 [ 191 :  160 ]};
    RAM[46 ] <=  {INITP_00  [ 187 :  184 ] , INIT_05 [ 223 :  192 ]};
    RAM[47 ] <=  {INITP_00  [ 191 :  188 ] , INIT_05 [ 255 :  224 ]};
    RAM[48 ] <=  {INITP_00  [ 195 :  192 ] , INIT_06 [ 31  :  0   ]};
    RAM[49 ] <=  {INITP_00  [ 199 :  196 ] , INIT_06 [ 63  :  32  ]};
    RAM[50 ] <=  {INITP_00  [ 203 :  200 ] , INIT_06 [ 95  :  64  ]};
    RAM[51 ] <=  {INITP_00  [ 207 :  204 ] , INIT_06 [ 127 :  96  ]};
    RAM[52 ] <=  {INITP_00  [ 211 :  208 ] , INIT_06 [ 159 :  128 ]};
    RAM[53 ] <=  {INITP_00  [ 215 :  212 ] , INIT_06 [ 191 :  160 ]};
    RAM[54 ] <=  {INITP_00  [ 219 :  216 ] , INIT_06 [ 223 :  192 ]};
    RAM[55 ] <=  {INITP_00  [ 223 :  220 ] , INIT_06 [ 255 :  224 ]};
    RAM[56 ] <=  {INITP_00  [ 227 :  224 ] , INIT_07 [ 31  :  0   ]};
    RAM[57 ] <=  {INITP_00  [ 231 :  228 ] , INIT_07 [ 63  :  32  ]};
    RAM[58 ] <=  {INITP_00  [ 235 :  232 ] , INIT_07 [ 95  :  64  ]};
    RAM[59 ] <=  {INITP_00  [ 239 :  236 ] , INIT_07 [ 127 :  96  ]};
    RAM[60 ] <=  {INITP_00  [ 243 :  240 ] , INIT_07 [ 159 :  128 ]};
    RAM[61 ] <=  {INITP_00  [ 247 :  244 ] , INIT_07 [ 191 :  160 ]};
    RAM[62 ] <=  {INITP_00  [ 251 :  248 ] , INIT_07 [ 223 :  192 ]};
    RAM[63 ] <=  {INITP_00  [ 255 :  252 ] , INIT_07 [ 255 :  224 ]};
    RAM[64 ] <=  {INITP_01  [   3 :    0 ] , INIT_08 [ 31  :  0   ]};
    RAM[65 ] <=  {INITP_01  [   7 :    4 ] , INIT_08 [ 63  :  32  ]};
    RAM[66 ] <=  {INITP_01  [  11  :   8 ] , INIT_08 [ 95  :  64  ]};
    RAM[67 ] <=  {INITP_01  [  15  :  12 ] , INIT_08 [ 127 :  96  ]};
    RAM[68 ] <=  {INITP_01  [  19  :  16 ] , INIT_08 [ 159 :  128 ]};
    RAM[69 ] <=  {INITP_01  [  23  :  20 ] , INIT_08 [ 191 :  160 ]};
    RAM[70 ] <=  {INITP_01  [  27  :  24 ] , INIT_08 [ 223 :  192 ]};
    RAM[71 ] <=  {INITP_01  [  31  :  28 ] , INIT_08 [ 255 :  224 ]};
    RAM[72 ] <=  {INITP_01  [  35  :  32 ] , INIT_09 [ 31  :  0   ]};
    RAM[73 ] <=  {INITP_01  [  39  :  36 ] , INIT_09 [ 63  :  32  ]};
    RAM[74 ] <=  {INITP_01  [  43  :  40 ] , INIT_09 [ 95  :  64  ]};
    RAM[75 ] <=  {INITP_01  [  47  :  44 ] , INIT_09 [ 127 :  96  ]};
    RAM[76 ] <=  {INITP_01  [  51  :  48 ] , INIT_09 [ 159 :  128 ]};
    RAM[77 ] <=  {INITP_01  [  55  :  52 ] , INIT_09 [ 191 :  160 ]};
    RAM[78 ] <=  {INITP_01  [  59  :  56 ] , INIT_09 [ 223 :  192 ]};
    RAM[79 ] <=  {INITP_01  [  63  :  60 ] , INIT_09 [ 255 :  224 ]};
    RAM[80 ] <=  {INITP_01  [  67  :  64 ] , INIT_0A [ 31  :  0   ]};
    RAM[81 ] <=  {INITP_01  [  71  :  68 ] , INIT_0A [ 63  :  32  ]};
    RAM[82 ] <=  {INITP_01  [  75  :  72 ] , INIT_0A [ 95  :  64  ]};
    RAM[83 ] <=  {INITP_01  [  79  :  76 ] , INIT_0A [ 127 :  96  ]};
    RAM[84 ] <=  {INITP_01  [  83  :  80 ] , INIT_0A [ 159 :  128 ]};
    RAM[85 ] <=  {INITP_01  [  87  :  84 ] , INIT_0A [ 191 :  160 ]};
    RAM[86 ] <=  {INITP_01  [  91  :  88 ] , INIT_0A [ 223 :  192 ]};
    RAM[87 ] <=  {INITP_01  [  95  :  92 ] , INIT_0A [ 255 :  224 ]};
    RAM[88 ] <=  {INITP_01  [  99  :  96 ] , INIT_0B [ 31  :  0   ]};
    RAM[89 ] <=  {INITP_01  [ 103 :  100 ] , INIT_0B [ 63  :  32  ]};
    RAM[90 ] <=  {INITP_01  [ 107 :  104 ] , INIT_0B [ 95  :  64  ]};
    RAM[91 ] <=  {INITP_01  [ 111 :  108 ] , INIT_0B [ 127 :  96  ]};
    RAM[92 ] <=  {INITP_01  [ 115 :  112 ] , INIT_0B [ 159 :  128 ]};
    RAM[93 ] <=  {INITP_01  [ 119 :  116 ] , INIT_0B [ 191 :  160 ]};
    RAM[94 ] <=  {INITP_01  [ 123 :  120 ] , INIT_0B [ 223 :  192 ]};
    RAM[95 ] <=  {INITP_01  [ 127 :  124 ] , INIT_0B [ 255 :  224 ]};
    RAM[96 ] <=  {INITP_01  [ 131 :  128 ] , INIT_0C [ 31  :  0   ]};
    RAM[97 ] <=  {INITP_01  [ 135 :  132 ] , INIT_0C [ 63  :  32  ]};
    RAM[98 ] <=  {INITP_01  [ 139 :  136 ] , INIT_0C [ 95  :  64  ]};
    RAM[99 ] <=  {INITP_01  [ 143 :  140 ] , INIT_0C [ 127 :  96  ]};
    RAM[100] <=  {INITP_01  [ 147 :  144 ] , INIT_0C [ 159 :  128 ]};
    RAM[101] <=  {INITP_01  [ 151 :  148 ] , INIT_0C [ 191 :  160 ]};
    RAM[102] <=  {INITP_01  [ 155 :  152 ] , INIT_0C [ 223 :  192 ]};
    RAM[103] <=  {INITP_01  [ 159 :  156 ] , INIT_0C [ 255 :  224 ]};
    RAM[104] <=  {INITP_01  [ 163 :  160 ] , INIT_0D [ 31  :  0   ]};
    RAM[105] <=  {INITP_01  [ 167 :  164 ] , INIT_0D [ 63  :  32  ]};
    RAM[106] <=  {INITP_01  [ 171 :  168 ] , INIT_0D [ 95  :  64  ]};
    RAM[107] <=  {INITP_01  [ 175 :  172 ] , INIT_0D [ 127 :  96  ]};
    RAM[108] <=  {INITP_01  [ 179 :  176 ] , INIT_0D [ 159 :  128 ]};
    RAM[109] <=  {INITP_01  [ 183 :  180 ] , INIT_0D [ 191 :  160 ]};
    RAM[110] <=  {INITP_01  [ 187 :  184 ] , INIT_0D [ 223 :  192 ]};
    RAM[111] <=  {INITP_01  [ 191 :  188 ] , INIT_0D [ 255 :  224 ]};
    RAM[112] <=  {INITP_01  [ 195 :  192 ] , INIT_0E [ 31  :  0   ]};
    RAM[113] <=  {INITP_01  [ 199 :  196 ] , INIT_0E [ 63  :  32  ]};
    RAM[114] <=  {INITP_01  [ 203 :  200 ] , INIT_0E [ 95  :  64  ]};
    RAM[115] <=  {INITP_01  [ 207 :  204 ] , INIT_0E [ 127 :  96  ]};
    RAM[116] <=  {INITP_01  [ 211 :  208 ] , INIT_0E [ 159 :  128 ]};
    RAM[117] <=  {INITP_01  [ 215 :  212 ] , INIT_0E [ 191 :  160 ]};
    RAM[118] <=  {INITP_01  [ 219 :  216 ] , INIT_0E [ 223 :  192 ]};
    RAM[119] <=  {INITP_01  [ 223 :  220 ] , INIT_0E [ 255 :  224 ]};
    RAM[120] <=  {INITP_01  [ 227 :  224 ] , INIT_0F [ 31  :  0   ]};
    RAM[121] <=  {INITP_01  [ 231 :  228 ] , INIT_0F [ 63  :  32  ]};
    RAM[122] <=  {INITP_01  [ 235 :  232 ] , INIT_0F [ 95  :  64  ]};
    RAM[123] <=  {INITP_01  [ 239 :  236 ] , INIT_0F [ 127 :  96  ]};
    RAM[124] <=  {INITP_01  [ 243 :  240 ] , INIT_0F [ 159 :  128 ]};
    RAM[125] <=  {INITP_01  [ 247 :  244 ] , INIT_0F [ 191 :  160 ]};
    RAM[126] <=  {INITP_01  [ 251 :  248 ] , INIT_0F [ 223 :  192 ]};
    RAM[127] <=  {INITP_01  [ 255 :  252 ] , INIT_0F [ 255 :  224 ]};
    RAM[128] <=  {INITP_02  [   3 :    0 ] , INIT_10 [ 31  :  0   ]};
    RAM[129] <=  {INITP_02  [   7 :    4 ] , INIT_10 [ 63  :  32  ]};
    RAM[130] <=  {INITP_02  [  11  :   8 ] , INIT_10 [ 95  :  64  ]};
    RAM[131] <=  {INITP_02  [  15  :  12 ] , INIT_10 [ 127 :  96  ]};
    RAM[132] <=  {INITP_02  [  19  :  16 ] , INIT_10 [ 159 :  128 ]};
    RAM[133] <=  {INITP_02  [  23  :  20 ] , INIT_10 [ 191 :  160 ]};
    RAM[134] <=  {INITP_02  [  27  :  24 ] , INIT_10 [ 223 :  192 ]};
    RAM[135] <=  {INITP_02  [  31  :  28 ] , INIT_10 [ 255 :  224 ]};
    RAM[136] <=  {INITP_02  [  35  :  32 ] , INIT_11 [ 31  :  0   ]};
    RAM[137] <=  {INITP_02  [  39  :  36 ] , INIT_11 [ 63  :  32  ]};
    RAM[138] <=  {INITP_02  [  43  :  40 ] , INIT_11 [ 95  :  64  ]};
    RAM[139] <=  {INITP_02  [  47  :  44 ] , INIT_11 [ 127 :  96  ]};
    RAM[140] <=  {INITP_02  [  51  :  48 ] , INIT_11 [ 159 :  128 ]};
    RAM[141] <=  {INITP_02  [  55  :  52 ] , INIT_11 [ 191 :  160 ]};
    RAM[142] <=  {INITP_02  [  59  :  56 ] , INIT_11 [ 223 :  192 ]};
    RAM[143] <=  {INITP_02  [  63  :  60 ] , INIT_11 [ 255 :  224 ]};
    RAM[144] <=  {INITP_02  [  67  :  64 ] , INIT_12 [ 31  :  0   ]};
    RAM[145] <=  {INITP_02  [  71  :  68 ] , INIT_12 [ 63  :  32  ]};
    RAM[146] <=  {INITP_02  [  75  :  72 ] , INIT_12 [ 95  :  64  ]};
    RAM[147] <=  {INITP_02  [  79  :  76 ] , INIT_12 [ 127 :  96  ]};
    RAM[148] <=  {INITP_02  [  83  :  80 ] , INIT_12 [ 159 :  128 ]};
    RAM[149] <=  {INITP_02  [  87  :  84 ] , INIT_12 [ 191 :  160 ]};
    RAM[150] <=  {INITP_02  [  91  :  88 ] , INIT_12 [ 223 :  192 ]};
    RAM[151] <=  {INITP_02  [  95  :  92 ] , INIT_12 [ 255 :  224 ]};
    RAM[152] <=  {INITP_02  [  99  :  96 ] , INIT_13 [ 31  :  0   ]};
    RAM[153] <=  {INITP_02  [ 103 :  100 ] , INIT_13 [ 63  :  32  ]};
    RAM[154] <=  {INITP_02  [ 107 :  104 ] , INIT_13 [ 95  :  64  ]};
    RAM[155] <=  {INITP_02  [ 111 :  108 ] , INIT_13 [ 127 :  96  ]};
    RAM[156] <=  {INITP_02  [ 115 :  112 ] , INIT_13 [ 159 :  128 ]};
    RAM[157] <=  {INITP_02  [ 119 :  116 ] , INIT_13 [ 191 :  160 ]};
    RAM[158] <=  {INITP_02  [ 123 :  120 ] , INIT_13 [ 223 :  192 ]};
    RAM[159] <=  {INITP_02  [ 127 :  124 ] , INIT_13 [ 255 :  224 ]};
    RAM[160] <=  {INITP_02  [ 131 :  128 ] , INIT_14 [ 31  :  0   ]};
    RAM[161] <=  {INITP_02  [ 135 :  132 ] , INIT_14 [ 63  :  32  ]};
    RAM[162] <=  {INITP_02  [ 139 :  136 ] , INIT_14 [ 95  :  64  ]};
    RAM[163] <=  {INITP_02  [ 143 :  140 ] , INIT_14 [ 127 :  96  ]};
    RAM[164] <=  {INITP_02  [ 147 :  144 ] , INIT_14 [ 159 :  128 ]};
    RAM[165] <=  {INITP_02  [ 151 :  148 ] , INIT_14 [ 191 :  160 ]};
    RAM[166] <=  {INITP_02  [ 155 :  152 ] , INIT_14 [ 223 :  192 ]};
    RAM[167] <=  {INITP_02  [ 159 :  156 ] , INIT_14 [ 255 :  224 ]};
    RAM[168] <=  {INITP_02  [ 163 :  160 ] , INIT_15 [ 31  :  0   ]};
    RAM[169] <=  {INITP_02  [ 167 :  164 ] , INIT_15 [ 63  :  32  ]};
    RAM[170] <=  {INITP_02  [ 171 :  168 ] , INIT_15 [ 95  :  64  ]};
    RAM[171] <=  {INITP_02  [ 175 :  172 ] , INIT_15 [ 127 :  96  ]};
    RAM[172] <=  {INITP_02  [ 179 :  176 ] , INIT_15 [ 159 :  128 ]};
    RAM[173] <=  {INITP_02  [ 183 :  180 ] , INIT_15 [ 191 :  160 ]};
    RAM[174] <=  {INITP_02  [ 187 :  184 ] , INIT_15 [ 223 :  192 ]};
    RAM[175] <=  {INITP_02  [ 191 :  188 ] , INIT_15 [ 255 :  224 ]};
    RAM[176] <=  {INITP_02  [ 195 :  192 ] , INIT_16 [ 31  :  0   ]};
    RAM[177] <=  {INITP_02  [ 199 :  196 ] , INIT_16 [ 63  :  32  ]};
    RAM[178] <=  {INITP_02  [ 203 :  200 ] , INIT_16 [ 95  :  64  ]};
    RAM[179] <=  {INITP_02  [ 207 :  204 ] , INIT_16 [ 127 :  96  ]};
    RAM[180] <=  {INITP_02  [ 211 :  208 ] , INIT_16 [ 159 :  128 ]};
    RAM[181] <=  {INITP_02  [ 215 :  212 ] , INIT_16 [ 191 :  160 ]};
    RAM[182] <=  {INITP_02  [ 219 :  216 ] , INIT_16 [ 223 :  192 ]};
    RAM[183] <=  {INITP_02  [ 223 :  220 ] , INIT_16 [ 255 :  224 ]};
    RAM[184] <=  {INITP_02  [ 227 :  224 ] , INIT_17 [ 31  :  0   ]};
    RAM[185] <=  {INITP_02  [ 231 :  228 ] , INIT_17 [ 63  :  32  ]};
    RAM[186] <=  {INITP_02  [ 235 :  232 ] , INIT_17 [ 95  :  64  ]};
    RAM[187] <=  {INITP_02  [ 239 :  236 ] , INIT_17 [ 127 :  96  ]};
    RAM[188] <=  {INITP_02  [ 243 :  240 ] , INIT_17 [ 159 :  128 ]};
    RAM[189] <=  {INITP_02  [ 247 :  244 ] , INIT_17 [ 191 :  160 ]};
    RAM[190] <=  {INITP_02  [ 251 :  248 ] , INIT_17 [ 223 :  192 ]};
    RAM[191] <=  {INITP_02  [ 255 :  252 ] , INIT_17 [ 255 :  224 ]};
    RAM[192] <=  {INITP_03  [   3 :    0 ] , INIT_18 [ 31  :  0   ]};
    RAM[193] <=  {INITP_03  [   7 :    4 ] , INIT_18 [ 63  :  32  ]};
    RAM[194] <=  {INITP_03  [  11  :   8 ] , INIT_18 [ 95  :  64  ]};
    RAM[195] <=  {INITP_03  [  15  :  12 ] , INIT_18 [ 127 :  96  ]};
    RAM[196] <=  {INITP_03  [  19  :  16 ] , INIT_18 [ 159 :  128 ]};
    RAM[197] <=  {INITP_03  [  23  :  20 ] , INIT_18 [ 191 :  160 ]};
    RAM[198] <=  {INITP_03  [  27  :  24 ] , INIT_18 [ 223 :  192 ]};
    RAM[199] <=  {INITP_03  [  31  :  28 ] , INIT_18 [ 255 :  224 ]};
    RAM[200] <=  {INITP_03  [  35  :  32 ] , INIT_19 [ 31  :  0   ]};
    RAM[201] <=  {INITP_03  [  39  :  36 ] , INIT_19 [ 63  :  32  ]};
    RAM[202] <=  {INITP_03  [  43  :  40 ] , INIT_19 [ 95  :  64  ]};
    RAM[203] <=  {INITP_03  [  47  :  44 ] , INIT_19 [ 127 :  96  ]};
    RAM[204] <=  {INITP_03  [  51  :  48 ] , INIT_19 [ 159 :  128 ]};
    RAM[205] <=  {INITP_03  [  55  :  52 ] , INIT_19 [ 191 :  160 ]};
    RAM[206] <=  {INITP_03  [  59  :  56 ] , INIT_19 [ 223 :  192 ]};
    RAM[207] <=  {INITP_03  [  63  :  60 ] , INIT_19 [ 255 :  224 ]};
    RAM[208] <=  {INITP_03  [  67  :  64 ] , INIT_1A [ 31  :  0   ]};
    RAM[209] <=  {INITP_03  [  71  :  68 ] , INIT_1A [ 63  :  32  ]};
    RAM[210] <=  {INITP_03  [  75  :  72 ] , INIT_1A [ 95  :  64  ]};
    RAM[211] <=  {INITP_03  [  79  :  76 ] , INIT_1A [ 127 :  96  ]};
    RAM[212] <=  {INITP_03  [  83  :  80 ] , INIT_1A [ 159 :  128 ]};
    RAM[213] <=  {INITP_03  [  87  :  84 ] , INIT_1A [ 191 :  160 ]};
    RAM[214] <=  {INITP_03  [  91  :  88 ] , INIT_1A [ 223 :  192 ]};
    RAM[215] <=  {INITP_03  [  95  :  92 ] , INIT_1A [ 255 :  224 ]};
    RAM[216] <=  {INITP_03  [  99  :  96 ] , INIT_1B [ 31  :  0   ]};
    RAM[217] <=  {INITP_03  [ 103 :  100 ] , INIT_1B [ 63  :  32  ]};
    RAM[218] <=  {INITP_03  [ 107 :  104 ] , INIT_1B [ 95  :  64  ]};
    RAM[219] <=  {INITP_03  [ 111 :  108 ] , INIT_1B [ 127 :  96  ]};
    RAM[220] <=  {INITP_03  [ 115 :  112 ] , INIT_1B [ 159 :  128 ]};
    RAM[221] <=  {INITP_03  [ 119 :  116 ] , INIT_1B [ 191 :  160 ]};
    RAM[222] <=  {INITP_03  [ 123 :  120 ] , INIT_1B [ 223 :  192 ]};
    RAM[223] <=  {INITP_03  [ 127 :  124 ] , INIT_1B [ 255 :  224 ]};
    RAM[224] <=  {INITP_03  [ 131 :  128 ] , INIT_1C [ 31  :  0   ]};
    RAM[225] <=  {INITP_03  [ 135 :  132 ] , INIT_1C [ 63  :  32  ]};
    RAM[226] <=  {INITP_03  [ 139 :  136 ] , INIT_1C [ 95  :  64  ]};
    RAM[227] <=  {INITP_03  [ 143 :  140 ] , INIT_1C [ 127 :  96  ]};
    RAM[228] <=  {INITP_03  [ 147 :  144 ] , INIT_1C [ 159 :  128 ]};
    RAM[229] <=  {INITP_03  [ 151 :  148 ] , INIT_1C [ 191 :  160 ]};
    RAM[230] <=  {INITP_03  [ 155 :  152 ] , INIT_1C [ 223 :  192 ]};
    RAM[231] <=  {INITP_03  [ 159 :  156 ] , INIT_1C [ 255 :  224 ]};
    RAM[232] <=  {INITP_03  [ 163 :  160 ] , INIT_1D [ 31  :  0   ]};
    RAM[233] <=  {INITP_03  [ 167 :  164 ] , INIT_1D [ 63  :  32  ]};
    RAM[234] <=  {INITP_03  [ 171 :  168 ] , INIT_1D [ 95  :  64  ]};
    RAM[235] <=  {INITP_03  [ 175 :  172 ] , INIT_1D [ 127 :  96  ]};
    RAM[236] <=  {INITP_03  [ 179 :  176 ] , INIT_1D [ 159 :  128 ]};
    RAM[237] <=  {INITP_03  [ 183 :  180 ] , INIT_1D [ 191 :  160 ]};
    RAM[238] <=  {INITP_03  [ 187 :  184 ] , INIT_1D [ 223 :  192 ]};
    RAM[239] <=  {INITP_03  [ 191 :  188 ] , INIT_1D [ 255 :  224 ]};
    RAM[240] <=  {INITP_03  [ 195 :  192 ] , INIT_1E [ 31  :  0   ]};
    RAM[241] <=  {INITP_03  [ 199 :  196 ] , INIT_1E [ 63  :  32  ]};
    RAM[242] <=  {INITP_03  [ 203 :  200 ] , INIT_1E [ 95  :  64  ]};
    RAM[243] <=  {INITP_03  [ 207 :  204 ] , INIT_1E [ 127 :  96  ]};
    RAM[244] <=  {INITP_03  [ 211 :  208 ] , INIT_1E [ 159 :  128 ]};
    RAM[245] <=  {INITP_03  [ 215 :  212 ] , INIT_1E [ 191 :  160 ]};
    RAM[246] <=  {INITP_03  [ 219 :  216 ] , INIT_1E [ 223 :  192 ]};
    RAM[247] <=  {INITP_03  [ 223 :  220 ] , INIT_1E [ 255 :  224 ]};
    RAM[248] <=  {INITP_03  [ 227 :  224 ] , INIT_1F [ 31  :  0   ]};
    RAM[249] <=  {INITP_03  [ 231 :  228 ] , INIT_1F [ 63  :  32  ]};
    RAM[250] <=  {INITP_03  [ 235 :  232 ] , INIT_1F [ 95  :  64  ]};
    RAM[251] <=  {INITP_03  [ 239 :  236 ] , INIT_1F [ 127 :  96  ]};
    RAM[252] <=  {INITP_03  [ 243 :  240 ] , INIT_1F [ 159 :  128 ]};
    RAM[253] <=  {INITP_03  [ 247 :  244 ] , INIT_1F [ 191 :  160 ]};
    RAM[254] <=  {INITP_03  [ 251 :  248 ] , INIT_1F [ 223 :  192 ]};
    RAM[255] <=  {INITP_03  [ 255 :  252 ] , INIT_1F [ 255 :  224 ]};
    RAM[256] <=  {INITP_04  [   3 :    0 ] , INIT_20 [ 31  :  0   ]};
    RAM[257] <=  {INITP_04  [   7 :    4 ] , INIT_20 [ 63  :  32  ]};
    RAM[258] <=  {INITP_04  [  11  :   8 ] , INIT_20 [ 95  :  64  ]};
    RAM[259] <=  {INITP_04  [  15  :  12 ] , INIT_20 [ 127 :  96  ]};
    RAM[260] <=  {INITP_04  [  19  :  16 ] , INIT_20 [ 159 :  128 ]};
    RAM[261] <=  {INITP_04  [  23  :  20 ] , INIT_20 [ 191 :  160 ]};
    RAM[262] <=  {INITP_04  [  27  :  24 ] , INIT_20 [ 223 :  192 ]};
    RAM[263] <=  {INITP_04  [  31  :  28 ] , INIT_20 [ 255 :  224 ]};
    RAM[264] <=  {INITP_04  [  35  :  32 ] , INIT_21 [ 31  :  0   ]};
    RAM[265] <=  {INITP_04  [  39  :  36 ] , INIT_21 [ 63  :  32  ]};
    RAM[266] <=  {INITP_04  [  43  :  40 ] , INIT_21 [ 95  :  64  ]};
    RAM[267] <=  {INITP_04  [  47  :  44 ] , INIT_21 [ 127 :  96  ]};
    RAM[268] <=  {INITP_04  [  51  :  48 ] , INIT_21 [ 159 :  128 ]};
    RAM[269] <=  {INITP_04  [  55  :  52 ] , INIT_21 [ 191 :  160 ]};
    RAM[270] <=  {INITP_04  [  59  :  56 ] , INIT_21 [ 223 :  192 ]};
    RAM[271] <=  {INITP_04  [  63  :  60 ] , INIT_21 [ 255 :  224 ]};
    RAM[272] <=  {INITP_04  [  67  :  64 ] , INIT_22 [ 31  :  0   ]};
    RAM[273] <=  {INITP_04  [  71  :  68 ] , INIT_22 [ 63  :  32  ]};
    RAM[274] <=  {INITP_04  [  75  :  72 ] , INIT_22 [ 95  :  64  ]};
    RAM[275] <=  {INITP_04  [  79  :  76 ] , INIT_22 [ 127 :  96  ]};
    RAM[276] <=  {INITP_04  [  83  :  80 ] , INIT_22 [ 159 :  128 ]};
    RAM[277] <=  {INITP_04  [  87  :  84 ] , INIT_22 [ 191 :  160 ]};
    RAM[278] <=  {INITP_04  [  91  :  88 ] , INIT_22 [ 223 :  192 ]};
    RAM[279] <=  {INITP_04  [  95  :  92 ] , INIT_22 [ 255 :  224 ]};
    RAM[280] <=  {INITP_04  [  99  :  96 ] , INIT_23 [ 31  :  0   ]};
    RAM[281] <=  {INITP_04  [ 103 :  100 ] , INIT_23 [ 63  :  32  ]};
    RAM[282] <=  {INITP_04  [ 107 :  104 ] , INIT_23 [ 95  :  64  ]};
    RAM[283] <=  {INITP_04  [ 111 :  108 ] , INIT_23 [ 127 :  96  ]};
    RAM[284] <=  {INITP_04  [ 115 :  112 ] , INIT_23 [ 159 :  128 ]};
    RAM[285] <=  {INITP_04  [ 119 :  116 ] , INIT_23 [ 191 :  160 ]};
    RAM[286] <=  {INITP_04  [ 123 :  120 ] , INIT_23 [ 223 :  192 ]};
    RAM[287] <=  {INITP_04  [ 127 :  124 ] , INIT_23 [ 255 :  224 ]};
    RAM[288] <=  {INITP_04  [ 131 :  128 ] , INIT_24 [ 31  :  0   ]};
    RAM[289] <=  {INITP_04  [ 135 :  132 ] , INIT_24 [ 63  :  32  ]};
    RAM[290] <=  {INITP_04  [ 139 :  136 ] , INIT_24 [ 95  :  64  ]};
    RAM[291] <=  {INITP_04  [ 143 :  140 ] , INIT_24 [ 127 :  96  ]};
    RAM[292] <=  {INITP_04  [ 147 :  144 ] , INIT_24 [ 159 :  128 ]};
    RAM[293] <=  {INITP_04  [ 151 :  148 ] , INIT_24 [ 191 :  160 ]};
    RAM[294] <=  {INITP_04  [ 155 :  152 ] , INIT_24 [ 223 :  192 ]};
    RAM[295] <=  {INITP_04  [ 159 :  156 ] , INIT_24 [ 255 :  224 ]};
    RAM[296] <=  {INITP_04  [ 163 :  160 ] , INIT_25 [ 31  :  0   ]};
    RAM[297] <=  {INITP_04  [ 167 :  164 ] , INIT_25 [ 63  :  32  ]};
    RAM[298] <=  {INITP_04  [ 171 :  168 ] , INIT_25 [ 95  :  64  ]};
    RAM[299] <=  {INITP_04  [ 175 :  172 ] , INIT_25 [ 127 :  96  ]};
    RAM[300] <=  {INITP_04  [ 179 :  176 ] , INIT_25 [ 159 :  128 ]};
    RAM[301] <=  {INITP_04  [ 183 :  180 ] , INIT_25 [ 191 :  160 ]};
    RAM[302] <=  {INITP_04  [ 187 :  184 ] , INIT_25 [ 223 :  192 ]};
    RAM[303] <=  {INITP_04  [ 191 :  188 ] , INIT_25 [ 255 :  224 ]};
    RAM[304] <=  {INITP_04  [ 195 :  192 ] , INIT_26 [ 31  :  0   ]};
    RAM[305] <=  {INITP_04  [ 199 :  196 ] , INIT_26 [ 63  :  32  ]};
    RAM[306] <=  {INITP_04  [ 203 :  200 ] , INIT_26 [ 95  :  64  ]};
    RAM[307] <=  {INITP_04  [ 207 :  204 ] , INIT_26 [ 127 :  96  ]};
    RAM[308] <=  {INITP_04  [ 211 :  208 ] , INIT_26 [ 159 :  128 ]};
    RAM[309] <=  {INITP_04  [ 215 :  212 ] , INIT_26 [ 191 :  160 ]};
    RAM[310] <=  {INITP_04  [ 219 :  216 ] , INIT_26 [ 223 :  192 ]};
    RAM[311] <=  {INITP_04  [ 223 :  220 ] , INIT_26 [ 255 :  224 ]};
    RAM[312] <=  {INITP_04  [ 227 :  224 ] , INIT_27 [ 31  :  0   ]};
    RAM[313] <=  {INITP_04  [ 231 :  228 ] , INIT_27 [ 63  :  32  ]};
    RAM[314] <=  {INITP_04  [ 235 :  232 ] , INIT_27 [ 95  :  64  ]};
    RAM[315] <=  {INITP_04  [ 239 :  236 ] , INIT_27 [ 127 :  96  ]};
    RAM[316] <=  {INITP_04  [ 243 :  240 ] , INIT_27 [ 159 :  128 ]};
    RAM[317] <=  {INITP_04  [ 247 :  244 ] , INIT_27 [ 191 :  160 ]};
    RAM[318] <=  {INITP_04  [ 251 :  248 ] , INIT_27 [ 223 :  192 ]};
    RAM[319] <=  {INITP_04  [ 255 :  252 ] , INIT_27 [ 255 :  224 ]};
    RAM[320] <=  {INITP_05  [   3 :    0 ] , INIT_28 [ 31  :  0   ]};
    RAM[321] <=  {INITP_05  [   7 :    4 ] , INIT_28 [ 63  :  32  ]};
    RAM[322] <=  {INITP_05  [  11  :   8 ] , INIT_28 [ 95  :  64  ]};
    RAM[323] <=  {INITP_05  [  15  :  12 ] , INIT_28 [ 127 :  96  ]};
    RAM[324] <=  {INITP_05  [  19  :  16 ] , INIT_28 [ 159 :  128 ]};
    RAM[325] <=  {INITP_05  [  23  :  20 ] , INIT_28 [ 191 :  160 ]};
    RAM[326] <=  {INITP_05  [  27  :  24 ] , INIT_28 [ 223 :  192 ]};
    RAM[327] <=  {INITP_05  [  31  :  28 ] , INIT_28 [ 255 :  224 ]};
    RAM[328] <=  {INITP_05  [  35  :  32 ] , INIT_29 [ 31  :  0   ]};
    RAM[329] <=  {INITP_05  [  39  :  36 ] , INIT_29 [ 63  :  32  ]};
    RAM[330] <=  {INITP_05  [  43  :  40 ] , INIT_29 [ 95  :  64  ]};
    RAM[331] <=  {INITP_05  [  47  :  44 ] , INIT_29 [ 127 :  96  ]};
    RAM[332] <=  {INITP_05  [  51  :  48 ] , INIT_29 [ 159 :  128 ]};
    RAM[333] <=  {INITP_05  [  55  :  52 ] , INIT_29 [ 191 :  160 ]};
    RAM[334] <=  {INITP_05  [  59  :  56 ] , INIT_29 [ 223 :  192 ]};
    RAM[335] <=  {INITP_05  [  63  :  60 ] , INIT_29 [ 255 :  224 ]};
    RAM[336] <=  {INITP_05  [  67  :  64 ] , INIT_2A [ 31  :  0   ]};
    RAM[337] <=  {INITP_05  [  71  :  68 ] , INIT_2A [ 63  :  32  ]};
    RAM[338] <=  {INITP_05  [  75  :  72 ] , INIT_2A [ 95  :  64  ]};
    RAM[339] <=  {INITP_05  [  79  :  76 ] , INIT_2A [ 127 :  96  ]};
    RAM[340] <=  {INITP_05  [  83  :  80 ] , INIT_2A [ 159 :  128 ]};
    RAM[341] <=  {INITP_05  [  87  :  84 ] , INIT_2A [ 191 :  160 ]};
    RAM[342] <=  {INITP_05  [  91  :  88 ] , INIT_2A [ 223 :  192 ]};
    RAM[343] <=  {INITP_05  [  95  :  92 ] , INIT_2A [ 255 :  224 ]};
    RAM[344] <=  {INITP_05  [  99  :  96 ] , INIT_2B [ 31  :  0   ]};
    RAM[345] <=  {INITP_05  [ 103 :  100 ] , INIT_2B [ 63  :  32  ]};
    RAM[346] <=  {INITP_05  [ 107 :  104 ] , INIT_2B [ 95  :  64  ]};
    RAM[347] <=  {INITP_05  [ 111 :  108 ] , INIT_2B [ 127 :  96  ]};
    RAM[348] <=  {INITP_05  [ 115 :  112 ] , INIT_2B [ 159 :  128 ]};
    RAM[349] <=  {INITP_05  [ 119 :  116 ] , INIT_2B [ 191 :  160 ]};
    RAM[350] <=  {INITP_05  [ 123 :  120 ] , INIT_2B [ 223 :  192 ]};
    RAM[351] <=  {INITP_05  [ 127 :  124 ] , INIT_2B [ 255 :  224 ]};
    RAM[352] <=  {INITP_05  [ 131 :  128 ] , INIT_2C [ 31  :  0   ]};
    RAM[353] <=  {INITP_05  [ 135 :  132 ] , INIT_2C [ 63  :  32  ]};
    RAM[354] <=  {INITP_05  [ 139 :  136 ] , INIT_2C [ 95  :  64  ]};
    RAM[355] <=  {INITP_05  [ 143 :  140 ] , INIT_2C [ 127 :  96  ]};
    RAM[356] <=  {INITP_05  [ 147 :  144 ] , INIT_2C [ 159 :  128 ]};
    RAM[357] <=  {INITP_05  [ 151 :  148 ] , INIT_2C [ 191 :  160 ]};
    RAM[358] <=  {INITP_05  [ 155 :  152 ] , INIT_2C [ 223 :  192 ]};
    RAM[359] <=  {INITP_05  [ 159 :  156 ] , INIT_2C [ 255 :  224 ]};
    RAM[360] <=  {INITP_05  [ 163 :  160 ] , INIT_2D [ 31  :  0   ]};
    RAM[361] <=  {INITP_05  [ 167 :  164 ] , INIT_2D [ 63  :  32  ]};
    RAM[362] <=  {INITP_05  [ 171 :  168 ] , INIT_2D [ 95  :  64  ]};
    RAM[363] <=  {INITP_05  [ 175 :  172 ] , INIT_2D [ 127 :  96  ]};
    RAM[364] <=  {INITP_05  [ 179 :  176 ] , INIT_2D [ 159 :  128 ]};
    RAM[365] <=  {INITP_05  [ 183 :  180 ] , INIT_2D [ 191 :  160 ]};
    RAM[366] <=  {INITP_05  [ 187 :  184 ] , INIT_2D [ 223 :  192 ]};
    RAM[367] <=  {INITP_05  [ 191 :  188 ] , INIT_2D [ 255 :  224 ]};
    RAM[368] <=  {INITP_05  [ 195 :  192 ] , INIT_2E [ 31  :  0   ]};
    RAM[369] <=  {INITP_05  [ 199 :  196 ] , INIT_2E [ 63  :  32  ]};
    RAM[370] <=  {INITP_05  [ 203 :  200 ] , INIT_2E [ 95  :  64  ]};
    RAM[371] <=  {INITP_05  [ 207 :  204 ] , INIT_2E [ 127 :  96  ]};
    RAM[372] <=  {INITP_05  [ 211 :  208 ] , INIT_2E [ 159 :  128 ]};
    RAM[373] <=  {INITP_05  [ 215 :  212 ] , INIT_2E [ 191 :  160 ]};
    RAM[374] <=  {INITP_05  [ 219 :  216 ] , INIT_2E [ 223 :  192 ]};
    RAM[375] <=  {INITP_05  [ 223 :  220 ] , INIT_2E [ 255 :  224 ]};
    RAM[376] <=  {INITP_05  [ 227 :  224 ] , INIT_2F [ 31  :  0   ]};
    RAM[377] <=  {INITP_05  [ 231 :  228 ] , INIT_2F [ 63  :  32  ]};
    RAM[378] <=  {INITP_05  [ 235 :  232 ] , INIT_2F [ 95  :  64  ]};
    RAM[379] <=  {INITP_05  [ 239 :  236 ] , INIT_2F [ 127 :  96  ]};
    RAM[380] <=  {INITP_05  [ 243 :  240 ] , INIT_2F [ 159 :  128 ]};
    RAM[381] <=  {INITP_05  [ 247 :  244 ] , INIT_2F [ 191 :  160 ]};
    RAM[382] <=  {INITP_05  [ 251 :  248 ] , INIT_2F [ 223 :  192 ]};
    RAM[383] <=  {INITP_05  [ 255 :  252 ] , INIT_2F [ 255 :  224 ]};
    RAM[384] <=  {INITP_06  [   3 :    0 ] , INIT_30 [ 31  :  0   ]};
    RAM[385] <=  {INITP_06  [   7 :    4 ] , INIT_30 [ 63  :  32  ]};
    RAM[386] <=  {INITP_06  [  11  :   8 ] , INIT_30 [ 95  :  64  ]};
    RAM[387] <=  {INITP_06  [  15  :  12 ] , INIT_30 [ 127 :  96  ]};
    RAM[388] <=  {INITP_06  [  19  :  16 ] , INIT_30 [ 159 :  128 ]};
    RAM[389] <=  {INITP_06  [  23  :  20 ] , INIT_30 [ 191 :  160 ]};
    RAM[390] <=  {INITP_06  [  27  :  24 ] , INIT_30 [ 223 :  192 ]};
    RAM[391] <=  {INITP_06  [  31  :  28 ] , INIT_30 [ 255 :  224 ]};
    RAM[392] <=  {INITP_06  [  35  :  32 ] , INIT_31 [ 31  :  0   ]};
    RAM[393] <=  {INITP_06  [  39  :  36 ] , INIT_31 [ 63  :  32  ]};
    RAM[394] <=  {INITP_06  [  43  :  40 ] , INIT_31 [ 95  :  64  ]};
    RAM[395] <=  {INITP_06  [  47  :  44 ] , INIT_31 [ 127 :  96  ]};
    RAM[396] <=  {INITP_06  [  51  :  48 ] , INIT_31 [ 159 :  128 ]};
    RAM[397] <=  {INITP_06  [  55  :  52 ] , INIT_31 [ 191 :  160 ]};
    RAM[398] <=  {INITP_06  [  59  :  56 ] , INIT_31 [ 223 :  192 ]};
    RAM[399] <=  {INITP_06  [  63  :  60 ] , INIT_31 [ 255 :  224 ]};
    RAM[400] <=  {INITP_06  [  67  :  64 ] , INIT_32 [ 31  :  0   ]};
    RAM[401] <=  {INITP_06  [  71  :  68 ] , INIT_32 [ 63  :  32  ]};
    RAM[402] <=  {INITP_06  [  75  :  72 ] , INIT_32 [ 95  :  64  ]};
    RAM[403] <=  {INITP_06  [  79  :  76 ] , INIT_32 [ 127 :  96  ]};
    RAM[404] <=  {INITP_06  [  83  :  80 ] , INIT_32 [ 159 :  128 ]};
    RAM[405] <=  {INITP_06  [  87  :  84 ] , INIT_32 [ 191 :  160 ]};
    RAM[406] <=  {INITP_06  [  91  :  88 ] , INIT_32 [ 223 :  192 ]};
    RAM[407] <=  {INITP_06  [  95  :  92 ] , INIT_32 [ 255 :  224 ]};
    RAM[408] <=  {INITP_06  [  99  :  96 ] , INIT_33 [ 31  :  0   ]};
    RAM[409] <=  {INITP_06  [ 103 :  100 ] , INIT_33 [ 63  :  32  ]};
    RAM[410] <=  {INITP_06  [ 107 :  104 ] , INIT_33 [ 95  :  64  ]};
    RAM[411] <=  {INITP_06  [ 111 :  108 ] , INIT_33 [ 127 :  96  ]};
    RAM[412] <=  {INITP_06  [ 115 :  112 ] , INIT_33 [ 159 :  128 ]};
    RAM[413] <=  {INITP_06  [ 119 :  116 ] , INIT_33 [ 191 :  160 ]};
    RAM[414] <=  {INITP_06  [ 123 :  120 ] , INIT_33 [ 223 :  192 ]};
    RAM[415] <=  {INITP_06  [ 127 :  124 ] , INIT_33 [ 255 :  224 ]};
    RAM[416] <=  {INITP_06  [ 131 :  128 ] , INIT_34 [ 31  :  0   ]};
    RAM[417] <=  {INITP_06  [ 135 :  132 ] , INIT_34 [ 63  :  32  ]};
    RAM[418] <=  {INITP_06  [ 139 :  136 ] , INIT_34 [ 95  :  64  ]};
    RAM[419] <=  {INITP_06  [ 143 :  140 ] , INIT_34 [ 127 :  96  ]};
    RAM[420] <=  {INITP_06  [ 147 :  144 ] , INIT_34 [ 159 :  128 ]};
    RAM[421] <=  {INITP_06  [ 151 :  148 ] , INIT_34 [ 191 :  160 ]};
    RAM[422] <=  {INITP_06  [ 155 :  152 ] , INIT_34 [ 223 :  192 ]};
    RAM[423] <=  {INITP_06  [ 159 :  156 ] , INIT_34 [ 255 :  224 ]};
    RAM[424] <=  {INITP_06  [ 163 :  160 ] , INIT_35 [ 31  :  0   ]};
    RAM[425] <=  {INITP_06  [ 167 :  164 ] , INIT_35 [ 63  :  32  ]};
    RAM[426] <=  {INITP_06  [ 171 :  168 ] , INIT_35 [ 95  :  64  ]};
    RAM[427] <=  {INITP_06  [ 175 :  172 ] , INIT_35 [ 127 :  96  ]};
    RAM[428] <=  {INITP_06  [ 179 :  176 ] , INIT_35 [ 159 :  128 ]};
    RAM[429] <=  {INITP_06  [ 183 :  180 ] , INIT_35 [ 191 :  160 ]};
    RAM[430] <=  {INITP_06  [ 187 :  184 ] , INIT_35 [ 223 :  192 ]};
    RAM[431] <=  {INITP_06  [ 191 :  188 ] , INIT_35 [ 255 :  224 ]};
    RAM[432] <=  {INITP_06  [ 195 :  192 ] , INIT_36 [ 31  :  0   ]};
    RAM[433] <=  {INITP_06  [ 199 :  196 ] , INIT_36 [ 63  :  32  ]};
    RAM[434] <=  {INITP_06  [ 203 :  200 ] , INIT_36 [ 95  :  64  ]};
    RAM[435] <=  {INITP_06  [ 207 :  204 ] , INIT_36 [ 127 :  96  ]};
    RAM[436] <=  {INITP_06  [ 211 :  208 ] , INIT_36 [ 159 :  128 ]};
    RAM[437] <=  {INITP_06  [ 215 :  212 ] , INIT_36 [ 191 :  160 ]};
    RAM[438] <=  {INITP_06  [ 219 :  216 ] , INIT_36 [ 223 :  192 ]};
    RAM[439] <=  {INITP_06  [ 223 :  220 ] , INIT_36 [ 255 :  224 ]};
    RAM[440] <=  {INITP_06  [ 227 :  224 ] , INIT_37 [ 31  :  0   ]};
    RAM[441] <=  {INITP_06  [ 231 :  228 ] , INIT_37 [ 63  :  32  ]};
    RAM[442] <=  {INITP_06  [ 235 :  232 ] , INIT_37 [ 95  :  64  ]};
    RAM[443] <=  {INITP_06  [ 239 :  236 ] , INIT_37 [ 127 :  96  ]};
    RAM[444] <=  {INITP_06  [ 243 :  240 ] , INIT_37 [ 159 :  128 ]};
    RAM[445] <=  {INITP_06  [ 247 :  244 ] , INIT_37 [ 191 :  160 ]};
    RAM[446] <=  {INITP_06  [ 251 :  248 ] , INIT_37 [ 223 :  192 ]};
    RAM[447] <=  {INITP_06  [ 255 :  252 ] , INIT_37 [ 255 :  224 ]};
    RAM[448] <=  {INITP_07  [   3 :    0 ] , INIT_38 [ 31  :  0   ]};
    RAM[449] <=  {INITP_07  [   7 :    4 ] , INIT_38 [ 63  :  32  ]};
    RAM[450] <=  {INITP_07  [  11  :   8 ] , INIT_38 [ 95  :  64  ]};
    RAM[451] <=  {INITP_07  [  15  :  12 ] , INIT_38 [ 127 :  96  ]};
    RAM[452] <=  {INITP_07  [  19  :  16 ] , INIT_38 [ 159 :  128 ]};
    RAM[453] <=  {INITP_07  [  23  :  20 ] , INIT_38 [ 191 :  160 ]};
    RAM[454] <=  {INITP_07  [  27  :  24 ] , INIT_38 [ 223 :  192 ]};
    RAM[455] <=  {INITP_07  [  31  :  28 ] , INIT_38 [ 255 :  224 ]};
    RAM[456] <=  {INITP_07  [  35  :  32 ] , INIT_39 [ 31  :  0   ]};
    RAM[457] <=  {INITP_07  [  39  :  36 ] , INIT_39 [ 63  :  32  ]};
    RAM[458] <=  {INITP_07  [  43  :  40 ] , INIT_39 [ 95  :  64  ]};
    RAM[459] <=  {INITP_07  [  47  :  44 ] , INIT_39 [ 127 :  96  ]};
    RAM[460] <=  {INITP_07  [  51  :  48 ] , INIT_39 [ 159 :  128 ]};
    RAM[461] <=  {INITP_07  [  55  :  52 ] , INIT_39 [ 191 :  160 ]};
    RAM[462] <=  {INITP_07  [  59  :  56 ] , INIT_39 [ 223 :  192 ]};
    RAM[463] <=  {INITP_07  [  63  :  60 ] , INIT_39 [ 255 :  224 ]};
    RAM[464] <=  {INITP_07  [  67  :  64 ] , INIT_3A [ 31  :  0   ]};
    RAM[465] <=  {INITP_07  [  71  :  68 ] , INIT_3A [ 63  :  32  ]};
    RAM[466] <=  {INITP_07  [  75  :  72 ] , INIT_3A [ 95  :  64  ]};
    RAM[467] <=  {INITP_07  [  79  :  76 ] , INIT_3A [ 127 :  96  ]};
    RAM[468] <=  {INITP_07  [  83  :  80 ] , INIT_3A [ 159 :  128 ]};
    RAM[469] <=  {INITP_07  [  87  :  84 ] , INIT_3A [ 191 :  160 ]};
    RAM[470] <=  {INITP_07  [  91  :  88 ] , INIT_3A [ 223 :  192 ]};
    RAM[471] <=  {INITP_07  [  95  :  92 ] , INIT_3A [ 255 :  224 ]};
    RAM[472] <=  {INITP_07  [  99  :  96 ] , INIT_3B [ 31  :  0   ]};
    RAM[473] <=  {INITP_07  [ 103 :  100 ] , INIT_3B [ 63  :  32  ]};
    RAM[474] <=  {INITP_07  [ 107 :  104 ] , INIT_3B [ 95  :  64  ]};
    RAM[475] <=  {INITP_07  [ 111 :  108 ] , INIT_3B [ 127 :  96  ]};
    RAM[476] <=  {INITP_07  [ 115 :  112 ] , INIT_3B [ 159 :  128 ]};
    RAM[477] <=  {INITP_07  [ 119 :  116 ] , INIT_3B [ 191 :  160 ]};
    RAM[478] <=  {INITP_07  [ 123 :  120 ] , INIT_3B [ 223 :  192 ]};
    RAM[479] <=  {INITP_07  [ 127 :  124 ] , INIT_3B [ 255 :  224 ]};
    RAM[480] <=  {INITP_07  [ 131 :  128 ] , INIT_3C [ 31  :  0   ]};
    RAM[481] <=  {INITP_07  [ 135 :  132 ] , INIT_3C [ 63  :  32  ]};
    RAM[482] <=  {INITP_07  [ 139 :  136 ] , INIT_3C [ 95  :  64  ]};
    RAM[483] <=  {INITP_07  [ 143 :  140 ] , INIT_3C [ 127 :  96  ]};
    RAM[484] <=  {INITP_07  [ 147 :  144 ] , INIT_3C [ 159 :  128 ]};
    RAM[485] <=  {INITP_07  [ 151 :  148 ] , INIT_3C [ 191 :  160 ]};
    RAM[486] <=  {INITP_07  [ 155 :  152 ] , INIT_3C [ 223 :  192 ]};
    RAM[487] <=  {INITP_07  [ 159 :  156 ] , INIT_3C [ 255 :  224 ]};
    RAM[488] <=  {INITP_07  [ 163 :  160 ] , INIT_3D [ 31  :  0   ]};
    RAM[489] <=  {INITP_07  [ 167 :  164 ] , INIT_3D [ 63  :  32  ]};
    RAM[490] <=  {INITP_07  [ 171 :  168 ] , INIT_3D [ 95  :  64  ]};
    RAM[491] <=  {INITP_07  [ 175 :  172 ] , INIT_3D [ 127 :  96  ]};
    RAM[492] <=  {INITP_07  [ 179 :  176 ] , INIT_3D [ 159 :  128 ]};
    RAM[493] <=  {INITP_07  [ 183 :  180 ] , INIT_3D [ 191 :  160 ]};
    RAM[494] <=  {INITP_07  [ 187 :  184 ] , INIT_3D [ 223 :  192 ]};
    RAM[495] <=  {INITP_07  [ 191 :  188 ] , INIT_3D [ 255 :  224 ]};
    RAM[496] <=  {INITP_07  [ 195 :  192 ] , INIT_3E [ 31  :  0   ]};
    RAM[497] <=  {INITP_07  [ 199 :  196 ] , INIT_3E [ 63  :  32  ]};
    RAM[498] <=  {INITP_07  [ 203 :  200 ] , INIT_3E [ 95  :  64  ]};
    RAM[499] <=  {INITP_07  [ 207 :  204 ] , INIT_3E [ 127 :  96  ]};
    RAM[500] <=  {INITP_07  [ 211 :  208 ] , INIT_3E [ 159 :  128 ]};
    RAM[501] <=  {INITP_07  [ 215 :  212 ] , INIT_3E [ 191 :  160 ]};
    RAM[502] <=  {INITP_07  [ 219 :  216 ] , INIT_3E [ 223 :  192 ]};
    RAM[503] <=  {INITP_07  [ 223 :  220 ] , INIT_3E [ 255 :  224 ]};
    RAM[504] <=  {INITP_07  [ 227 :  224 ] , INIT_3F [ 31  :  0   ]};
    RAM[505] <=  {INITP_07  [ 231 :  228 ] , INIT_3F [ 63  :  32  ]};
    RAM[506] <=  {INITP_07  [ 235 :  232 ] , INIT_3F [ 95  :  64  ]};
    RAM[507] <=  {INITP_07  [ 239 :  236 ] , INIT_3F [ 127 :  96  ]};
    RAM[508] <=  {INITP_07  [ 243 :  240 ] , INIT_3F [ 159 :  128 ]};
    RAM[509] <=  {INITP_07  [ 247 :  244 ] , INIT_3F [ 191 :  160 ]};
    RAM[510] <=  {INITP_07  [ 251 :  248 ] , INIT_3F [ 223 :  192 ]};
    RAM[511] <=  {INITP_07  [ 255 :  252 ] , INIT_3F [ 255 :  224 ]};
  end

  always @(posedge CLK)
  begin
    begin
      if (EN == 1'b1 && WEA == 1'b1) begin
        RAM[ADDRA] = {DIPA , DIA};
      end
    end
  end

  always @(posedge CLK)
  begin
    begin
      if (EN == 1'b1) begin
        RDATAA = RAM[ADDRA];
      end
    end
  end

  always @(posedge CLK)
  begin
    begin
      if (EN == 1'b1) begin
        RDATAB = RAM[ADDRB];
      end
    end
  end

  assign DOA = RDATAA[31:0];
  assign DOPA = RDATAA[35:32];
  assign DOB = RDATAB[31:0];
  assign DOPB = RDATAB[35:32];

endmodule
