// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:35:39 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
XyoQ9UV6hlsvqgPZw4Rjfx1FdUH3HxIdUqazdZC4aHCytQKDh+56H2eLUFelXNnW
8oEoxY0rrFYS0yUPjXETffHdWKRzZP5z4yZuRosCpLFwgQb67GY1Kou/Myz2nJAx
KlAOUjAt4H34Pvg1FudbJYuqQkSNwIlH+nLL/yYRuSc=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 4352)
Tym2RGOFAcqUxmPyhYyw+ESI+afVL/bSwu80aAdHBks12Kq3/ZhvmB7ZefMclMAo
ZKtDLwFJ4mCOURImLXB9/ne8GQOYCqmahl/NZZxeTcRCR3ZH+ikJ5nz3jfXzee8z
iQ68COxfrB8sWeGXiiDJ/1JH+HLama4S42+8SXfGutMylBkMgQ3TNMVCDfipovJc
aITMIWRsDEKsUp+4RIq8cD5pJZO4nobcaHxytSsCX1BkG633Izpw5Ff3XbhFx+bJ
Jzco4EX9bxrofo6ts/a7BU6bwGfxD928lqhrd5QYsS+d6NVL9/6QH/CE06Z8Qqtu
nAbLqmrFyaljvXhuME9LSyv9eP8/y75we/VUXUvy0FnVB+r7rhymwXnVHZYww6YL
13+xGohPkFQzVqfEw5U59z4AV6ooWRcOJes8wZRZp6t44/rT/ls35PAohwYQVviy
Rrsc5timyOkGmGSa3wE2pJ5qAyx7alq7+9KpHpLfw4fdHtI6IlaIYA0gMUmESPdQ
TVrutZ+joQJI6wxdpRzhjqOtc4fkF0TOpsXWqSfi94XdYSLUs4jLJD9dEjPL+PKj
Wf6t583iZZjATbwF8db8CNALiwuLYqDKvNfESVzrA2yp2FBvfL5z4/6FxwfpJmV3
hhY7QiD7CtWjw+/5HfUH3uXBYioiZvsJ20LExV1oKpM7PcKkhJmrJvqMHRPCXBfu
mEDG4g1J4iHpsvZyi1Ma/33IPswkTwrTZHBBs24JqG/fbupjYSqAiWwNccvEoBIF
MkU9rDsAL/ycppWD84VApOxHLdGD3ya7r+BLFfJfumhv6ALwP1o2L4+sidcHeuPo
/wtEj6ECeu8VBXPs5kiPtp9L3kREEsH8HYPpI7cZ414UsQ0ujsNc47hwUu1/c/ob
B0Igqrd27Na0Sgek8PRDHM1gLZpiJ3smB8rTy+cQNyJe5bh2XO1OHQWQf6Xk4H4P
6j0RreaRxVxT4LAj9SprVhbeLIAQRHZZYtK47q9yNiEaTAAbSPujg75OS30teLPx
Vi3+M66BbBfupQCVzhepJ/dhTztdjE/vcKOxoC+MFU8zyL5HMiD4kNQY5/K9VKxE
bw8eF/aUhMFJNtqxNDkCgr0zOdwKWfqDP9fiVQ+r7MjeK8M2u6HrP8hDdJmGMFW6
RYveaXhd8iPhigrVgCxkVL5iD/utBeJPsJa2MiqeM47BeXNEJgYA1JYjQjGL95AD
xJDokqaWUuxVUqV8dg3KTPO52Z199MeT1KJgyuxQ6ev8ezQFnGTEPx2GYQgwyoPX
m9wJHuAjLmD/kSAsBh793Uw7Eo7l2dzcXlkhlisvZ3GWU07KedkfvLBbfjuC4ZzJ
qCIlZuRFhztgKZCbXIRIyIG8d0XqhQE5E+pIbtgOODa4C6mOTolxd0w6RRtlo0gF
aRt3VquKrUS9o3XrOGrblsKmqm6xsRPFky5YN03zUFoN9eEThY+ZW5WX5/zM72Nc
1kCxzp5Vfy/xblBLPx9ruBWb53o8RG4hE/NxF+N+SbqQKH2peWKYfw1nNAbsNNYe
PJQzQEIKVL8et8dopunf6W4tRvA4FzfddItZrY0BeIpHuXxwhxIK+UU0FGtLT8Tl
QbNLXM4+7b6zcsDBcobQuarA0XjThZB2MVKAnY1JUtPKHd95U8Cm5UeZlf+ULXHq
XuultTknv0e7e/IRSkK/0401KwcF8I8lTgrrR60mw73FoZRjjEurH6yS7j41kAUX
n/jEcvs4gUbp93jBsiyDzjNVYqkL52kY1mNzRkkCRYYb5iwAdK+IqehDMaoyWMf6
TFYDiTBGwuuk/eXnv3Uow9GG2VEj9C0huFQycw9FmyEwc7se0/QURO2v3fulgx3T
1D0IbKmL8rOFrXcpn7lGRNjbtfV5LpOfZmK7cecWGQak1qo+lb+ovtpfxmn1biVB
E6t+S1sgWxx5QXOelyw56OMyGHcgM/c1xzv7GEXsm8TYKEkI/EPLLEymEqnMfhL5
9luWEWLpHAj6TIqrEv+9wJhRI6EBhlP2oB6SZWaKVMBnjgWjQql/avr6XF0v6TvV
219Ooi7+U0rAY1Ovy6hnZ7qjXJmVeBEkxzhzKM+4ETw1JiPSgZyAjd3w90zMCLCI
xC7TPImEBkriX2LxuWHrsU+xdE0/H4RWJy8QpdEoM9MLLx32FP6jHBjUFI9rpaT2
0aIje5Iub/IZg281zQDKpKthWQW44RsVEWORcAb6Jtf76llyUuuzqCDe9eT5X1tA
elElZixz6TcCCtkUVbkzW9gFOsleSxv/1jnCHLBppWeGGfxvqoLCechdjBv2vieU
3sg94rKUnaRCaoLAZeoJlwy329x/f3WQseqTaQQcZXOxjeWWugXe8UPS0cyaoQ5L
NfLrG5Ml6qylAMIaKw8jAqeivcoZXDJkTJ5JKcP2td4AVd4aUH32Q2bo2Q+OxCzh
eQIKyyI2ObDb/4VHcxyH7bKHHqjNVX/gn3MiO7RxFR8GQSkPX0E/C3cuKcnNeaRB
F47f2FUrL0bQ+qARnnqLj7hIkCbnxreAAhTZMoDN67JlRKF00x9gpspPXyV4SgYD
ttxcxG/eyQ3k8ITv0W+1vF2RBLNPckOZrIBYX/G1hxOJf5aV0z2Y7ZwCZ6yOdO0T
DLEWVQEzlSDjGeIpeXXLpluMmNYOfqFKJUWS+CvWvK2nSaz2fCp4qYv0M0QIBNlc
yAAh/Xs5l8PbBKrVx0AQH1ma5Rtc4+DvoLpjxG7CeAaG0PzkTSvWp/giQ3Q4cVdE
svDAtAf0e1E+JZwh/ehofPM2KmA3EwuP5/n8TOah08bZAQ34viX64hTevqYxcA51
UYCQ3wM7MoM2RgVc855MLlel0/cKTFSrGZ89x/J1QAIz9ElJzSNzZl6RihmRdoIf
vmhYtXRbp1v2bRC40+22UGzwz4ATSmi6VEYVgzl0iW0FDt0BWjbvABLFWOgZAA/W
Pah/JgD7Yn+pVtaiXeHyvky1IDA75MWAnroxOCRqW87SzidYdAGrbg51Len0v+Zd
0D0tthARMx2sHcLdb++mFtCSDrbsi6rN+T7tDabZsYYgdWRS/5m42RoIrjl28nvw
AL9NZ+A10n8lV1qugvRuVAoXMVORxSSVl2yFeOnrNY971B1jYT6H8uYJDPO4vcuS
rgW/hBjF9SDE2YUMrl+4drFdhcmsAfLF2TICnwDhS07OaHqzVy0lDmu0sTZRUqWW
gvjEZdIqk7A1TKElj+o6VEfPZmM8m5qv7gaRA4m/4Loi9XUcJFAXZJ5cDmj6fz6V
u5xeLNfnMvz29nsxLuD4xXc6IAlZ0P45Gg53ifqUbvdN2Vi1sgnytBS1fgG1dOsF
tFKtG11aZk96PsrXWwaee5ciI4eOn68TYcXxqTbryYSwOtz6fUfKO2QRSirC8KlH
T8WsnLwbEHi8eCkg07t1kO4Okzhc6Ue2QqtsKSGXQB2mZnpEBSexwZcOVHJMPkC0
f5uOhSCl3r3sw9ZrWsgXw9IkvRzK7bBSzGdK7ShNX9UjvBU9RWAhAylztnmGT8nG
KPwJXR3ezpD4fHs/KuDSAqApdWrTDbTj8ymXbpwzzYxBkIFQwk3JQqK7SEovAcA1
7LTgToFiUubuvRPtD+7/Xh4NOW+zX7U43vpz8RtYiLFE9acIRGHfQhRzjBzrRNWg
MWe5wOSXCX0okhvh+AX3XRWP2Jy0zTB+MPgkKQ5ZZI5LQVT61Hu4ks2kHiHAEVHQ
KlRq5Gt+fs2eVEbXC8auf7VCNWTLZEAOUfpbKeBjvs9uDlPlInZ6MGiwyChqb4Dy
9K8hWNHFk1HRWx5lKCbqAPaDmc6KSOF/K7V+EDzIrq337hYigFowlTJJVKM+yKAT
GxJIyzp6nHdUGqyRNDhswjNlRH8bFz89kto4bUHvtw8lecnix7cThBVhqhXLIe0Q
TtMMYaPnY2CybMen7ue8FSFuryddbPiza5RA0KJw4S0nnyMzAwPIpWHBeG5PAihQ
5XUMP41kW1bQoriqIvAPCxRXa9oqPXCNwF9s8UHL/V8iWZoXrEEtYJPk5EmuYH4K
B/fIQgPqXwHzTcEmjXLQuoQBCbZLCtvG/7s5L0dMR4SB+PUB36i3MyQ8NnnHwIgk
ppwMjmWTX5CdaT6z5IJFndgFQxcUKRfEMMXqJx0CqK752oyfYhVr9MekEzvqiaUD
946r6X/IU3Hu5eHVeQqNAGSyUV6U0/gLpjwLqtIT5coa/3TjAAdCLw6P4Z+veSb2
HH12F+hwyR8WcuDOpQ9NU9673UgRW9nk7UEomoqppkVX/I8kulFnzEgiHj2PiRVz
W8CFjhDB/mft5hhIfLvsQFjjbsUklbgE50nfxfuJr5vettRkaEVeuLZF/AYYT7HN
asbbJZg64a2uwWne/M/MuEjsRIG+NmmJto17d4k3xkzkZyKZ8ddy7o2iAm4kStcw
sBr9PyKeapn47WFqSuJHptiumcJtSfGGomGYbSvLF9v46mjES0/G/mdYuqRXZktj
UUiC0RSP77/AqUqfjyjIJbybJvqrxdR0FRWd90pYGxb0B2DN6VJKcBOuKsqDEjci
NzwZVJ7cZ5VEV5fBoMLS9XntrM2emaHis0wXhjRuDRGwOuxsLI0SGjIW1kpAauUR
rKp5XQoDmJb4IAQlUCgCdH8WuMjODStMy4crFrm4oH8X/9t7aD9mypYf3qr6cYnh
TGQj+xvQkaw/st6uyl+DEYXqss8r8UJLY64WkZW07GAcSBFF3hWeBVHsi92k9R9g
fJBrCBUawwhjL4JVC5cfO9pHHYSl/AF2KPcfBGU8HcVHDwEwNz8F0lPYRGqAX2yJ
Z3GqkLQ9DGuRBOPod8UsamThTsgfusw+ONX5xtnzotw7qe7FZFk/Rjwc/UeVCI7h
xrSVk/SyB/15/BTAZEwxWdvdp6JKVGNW/eTxm2TImjboX9J3Dxr+2F5yFgLADC6v
koUEPYQ2HncSGr7b1culpks87UausU2K9qKSpqP+byvaA36N+oELMIr8GG9Za0kx
yH310GpjK0imKb6X8AtXx3ZO/nEtkDJMpNh7nusPebNGIrordmPwzhxw7+l7FHGV
BNrYG4W6aJ28fRYQg9arrAgQUWD5o34N2czh62ogKsk8kmR2Z96Ibo/LiJxLdZaa
7Pv5MSPCgDqGNnN3aoYpEwr87TkkAh91z9Yb+NXo/htsr/1fle8cBRTcSjRIRS/L
3hTmunT3dhrcI93mcWddOYrKU94NYkBytzGj7B1LgcNP76P2m7svWgi+13vRjYH3
6zPLGzvQ7yxLGBbiZKGi8dvZJhrG6dH6jCbYit6GPH6Vby0KTnLSVQg5+p6RuKsL
SM4IxuY4BBZR17IAYwCJB5MlpnR1vennRB0KVUOjabdo8lGNicwgUYgyLBYbVwDi
ZBwVmF9XwDJeMPbhy8fle6eGDuy3OH2hnJdYMkSUdaP9Z4Hh2YvAKV8xkoZQ3hgr
8ky9+d6joPhkoQerWN/S3S07e/CPlGT9Pc/LbsudexoYFI/5GC1yCAv03OkAQVjz
GoJFG/Rt8TH/RL7O5pEi2CYv7zf24pmUMrDTkirkVGc1Ib0+0ooXLn8YnC3o5+LC
OEongYY41BAeBZxC4Ppj+vV6CSBDphB9sd6TIrFxYMYpuwSQ89rclth9rRJM8+Jk
BSpKOlhEabmhU+g+Nvwh+n/jSsORJaX2kA1T8WHt1McUOnKFri8K8mrXoBGnfmHT
KafkrVmb5MYKYiwWCxubr0vJDZOoB93XhjDXsw1Nqk3txEPT84ZPlW36GSCmpJoI
rBY/VuN/6k5vRU76275RzTqW64Xv3+o5/16i9BlXfvE=
`pragma protect end_protected
