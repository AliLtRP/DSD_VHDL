// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:24 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
hdzntQQCTH5MVSQjHAM+S1FW5pQMw9IZEzXoPAiquChoemssjrfvUPCWKNf6pAT9
bPm3a/2cQSNcEjaj1g5BGgZ9FxPLyG5wsO6kFmQxyY2ewESV/laGU3K2fzWRALUY
dQPJ1rx5oTy6XNTkrHEBWrQPzOq/83Lz6lV4CnaYkxw=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 7424)
HenWWKOm8yxWOTx3RUdHLbI+GNcuS1+JAyADzUMtyUaXn5Jmx4nHsAAMZoRE3TzG
oU+QfxPbNPl3GxDRBCBJb13lb50WkY+19sKBePDbaSKyz+ob1qc3SwXTJofiitH6
2TpmWb1fWk6redy4/BJe4Eax2SwcJ1QKm7YEwVFtH26CnI77g5WCqVo+uDmNItD1
W7lq7yAXQbNYXcxR8CukW3JivD3sqA4tYOM+iHP1CKkePiUksguYmiWj2368t5vX
ubffSkoKiSs3XfRk2z0Xu8JjtgOLVaISV5id1DlqleDBcZ9fuGOY0S6htVxm+skr
EFLlky+I67hpzSWpyTEN82Me2BSG3OwFApPFzZj/U7mWYvhFUL6WJCk11eBfDbfl
QamIqCQRywsqMLA1dLQkX+w1gK0gHQnOr24040/tvk88vbsNZkAAAJ/VPwk/Isto
BAH0MksFQ1L6sfOLapCvYydWwVS2355J/EVqnh657j/PhJhmMpxgo4hb3A9M7jwM
IWqN1EhxfoJY7g4ExHw0rzDbxTqFs1Rj5ZxaX+g0DyTAIKEL/XYGebiCS/hj8qi9
1hxUoiFwWFAgwD5txAgUhgjsYlg2Alqb5/mK94MQv99vL0sqfnRAw76QQsyjAlTm
018ftQb9D2h1ScoM5HTl2g8RAfXQ/+bTnRZhweniRrQnUjEnI2q6r16HNMWp/ex0
T3p6RiQ31SwW4K7peLIbctnLpk+I6+jXndlZU/IP5ZxOp2CPXKjyeler1QY1WvM8
3Yfe9xWPP5dxRF2skEolC/IoUSmShuhWZsfoZXnQDYYOIN+GmtfMZ6N6jhyRnEGD
u3asMI66NXIajD3AMcy6WvzC7hTkawnHAyIdVgxD3hDgjQLdWEKm7ALvNnlfcb9n
QFIAP0WBMqltmVYI0ulS0GgnAXGhe2wCekClrxtmk57a0sYQX2WRSYgGsjiu8gQL
QF+goZRYSqWhysACMshDMnv1viumOofRWQkRMhhErXeDG6zjyP+vSUmYRnojK+VU
LxzYy9Yz9v+B+iOO1SsyarUWQsjUC95NwUX1BbKOnupd4Q2+ncgoykbNxWTIkpT3
2tNZDSXr58blu4o43qvyHKRp+EmIaNNAeC40HSmzuozs9dWvMOgRwkswuv081J5z
dvd0HXTJ34oQ8bSd2tRiP/b971ygBhvm0/XMxxFtMDoDx+UqlAuixI0Ljb9x+1it
ipOtzyYOmAxnie1wT5Qho6xVH0AhTDRS+kEhVan9GaHUVLk1MufzymiovOnJGO7W
ULNtImOJ5sj5l+plA0B4cVq4OEqJrHSmcOsnoxIKUT5remM5/5u2zoLo/9z+0jK1
4TIMADByQgDQY8W1DbHYdeSWHSllSKqzEjTrSZVvIRAmf5v1CEPPKrJd27lnpxQP
DjnfkujOjAgSEete5RKIJjQ9I/Fd3Qo+VZvq6fC5FF5irt0Lli7D9USln9dPvoDZ
P7qN3u0jy+LHPrBQFoogDj/Pa1ezOqlU1z6COjisGiI+b4SWUTVhUkIXchEOljlz
TR7u963GKAxSwPc+f0BVWU3xtofSIHnZji1AY9Ij3c/8yKXyt9a9YTQiWxn/2aQU
kmsNj4X1bqCd21ktB4wh9Dclgd8S5MV4peBclp2aUucD2m+v9c6YXLvqb8t8TALF
uTleiPjL90zJ68Lb0kDjSYBdFXcS2a2hbA+ln3kSv2P7F3flO21WPOQXmoROn4gn
fz/eTE2zjwtKCjOjb33SaeZ3t/yFGt2Bey1Z5pkLykxyDZ9o1Kf6rd2iuK+K3Ke7
8HIxuD7Rzu6j0PI2sRXGa8rCCKMs53E3lJOsOLd8vkJG36Z7qmK0ULuZ0kpxKH/f
GHIiqQt2gcdQ/66SwtnO7qYBeeNs2KiOWD/n1Xuo2uaw3wEns30TVMd815MGrulI
WParV6EHlBCe8YqhOIIqeXaF1DZrbd9EtVpdZcIcny9WOZouMNRfmzrUacZYXhCj
/GT8dwnCzCuQYZMDS9BNt+JCDFX5+uqTmnqW657//TkhR3j8yIn8C6m5wlt2d3H6
r+nUauOU8zjReJVqBUAYaKILU+zoKDvdHQDhZn+YieXrz/O51Nul1Kx4YwKtgx0Y
exV32UyIhT9Av1dG8O/NQc7pimms9SAVrF5cilGeDvkJaalxTWGdJGlweLhbQV00
gQwkJIsL6v9qM9oeoEABaYJG/J4ITnoTNB1hkq1iLagRCxQonVkax0Nq09DDjhZ9
9k+FJbgGxqWyJX5RmcWrp/gzpGKDn/CS94yzeLNskJ1unuLP0CmJY4fBe3Bk2T3s
aapHxUqxX5QdjPCb4xJP69ts88ifOBx6PqSMB+cjUbEp3sFpbNv0Wwm0Xql5M9ye
K7238On66lmTH1gvyfAWYATeRq35L8m/p2RwmUGfwwP9t4qp6XUqsp6WQz0eP5xQ
9BtkzYxfwfIMwiXhgQqgUFQBgi6fC90UuCUOe+CRPxME0leOOCXuCcjJi3Az0rmk
iljHaIqJBHYyFSHLadPg29SBS5BsDJaU8KOxqxAMOm1YcgRlumeSRpyRZnKEEFQG
CTvMO8disBadel17KwZwLdj/+kviiUd9lSuARrmqodHtGBjmeyf1hqlwySWPSgmH
XgKdAXp0cvdLbUesUtp5mkkwORAw4jrCGe4jawRolaRntygLOn+M0l/kS1nWFZA+
h9Uv85Y7J0wEKjphV1zc38wwFlOmjWCjoTYgz2C9yeJ0D8DXFBpJfT1IVpiC7kYJ
xMFKGLyMMHfe6wjhUeLY2sWEUuBE1DzM8j/GOvRGg8l6wUy5V11YPgsCh2lGNxIa
QeS3SGfZQt8CfG4OZBmLNSLSxPRUfcUImd5zorn3lHg64QA0Jkm+hu7FjMbnJl5I
/5rpheFQzU83CZLs5+Tn+SktzIZkWWy9Az5pRdh8KhGLrnx1mfM2hFn5ZPC/HVtu
G8vuKyjZt0DgL4llscD0YbBLbYQfLiSlUllRmFXoef84nGTI98yfh4pNG490vkow
V2zB20uQf3gbM+/95FBe2Ghzo4RVhldK7EGur/NNnh9gTay6FVCEYKY9Xa9Bkbz9
8YdicdLBYyHaKWT5KimQGHlfeUeLSblfHic4Y/hSbs2IAWLjryb6DNp9LHK+OddR
1kXv56v8hGtGlsn1maoKWFOexF5nXnxS0GwymzWNsmOISRUKjbMUESJl+L66c6Xw
nEgqxL+NjAMg/gEczxHIQDHH3um41fkAowNfxZaMgaPhgVdiIgPhzAfWz1q9SMMp
t4NGI7oKmWREUV9g1vVuT7xLFlBu52PJ6v043e+2K0/IrW0de0oUqSrCqXw+mQmG
mBHl9b21NN1+mpCe6FKd4eWGYGQ49XpeCfSZb9MxxbNwQI/WcateGGwrmHbfb1mC
sgSf9Q7YUQ5Ui9aGZWvH+Flg+rPmYKcjK/kHVHLXdeGxei8uoOFTBg1VjU6SG2XH
oNxXS9A6fybfaM6P4TFeNiGx9NJdujw9yFZNTtVPjdu2M0f4Q2x3PPCUwxaCIyBT
sl9aaFNYMTfaR/q+gOY5h7OBTmPF9MQ6XcVfMlWtODsVGkmnbp5H5jAaOZj8EWiA
XpWLKhySgWcLD6uku5MGhS27Rtn2VFstb53sRvzRNqbIxJCJr25XOrcmFYzidUWP
0vA5A3q5hbAwj6bru9cPKARVE7qqj2FOfdvtBND2MnF/iTMEGk8Ii0MKhXh8QZsJ
L5AjKu9RIg7/kMiXvJkjkc/A2qOmsFPrf2VJQ1Zuhf6hknFPFt9sAahmPgAgv4/R
0N5WVkxnBIzkR9+J46slTqy1XQ62PprCfEFZUCJz9myd2+7sa/aVPbokOaiYADdt
YdTTNDe/YyDMh8tm8U/SV8F8lb6psZGlsGEEk7BDgSAXsp86Cd+zN9hTt3rNlBhc
ItNTX6PP/5MKNS3pibliBiaNPE38bU170YWUA0MSjLINNheaq1arO4MfVXMGhgPp
wd7PsdmU1cj1CIWUDe+z+vT+4luuehTrS1a68tI9Tr1/4obRWtOlqWIxhNFHh6pU
b2xuAHT9bRB2B6W0mDBRTkPGa99pdPj9CcSPtSawbVLVxFkl9NSllRkN7tJWPsRR
fy96rgwmEAmWc/rOMyvwOW7ywenpj069KMIy84V/dNQUhpJBPyzjPY28QkC6yqzH
Zaob8R+cbjucvj9rWOV8/EZWHN0oU/NEk6qvPdLbnk+Ytlm1wQ9VYgAj7fpQKo0+
BXlGQP00jGsgeVGSwtUYsVIOiF1MvFOdc0Q5tsd4fR71pf6AKgW7JNX7glgzM6ue
BbzfAtJeCaIMxCsFaKYjxBq+ReP/cdAsdoOMtF0/nzVRJp7t8oD7is/4WrQGHD74
1hSRRsZsozuINENkbtMBIVfSVS0kTzYuEvKNkg3R3Rol8gWmn39FfAv97TrvLPqK
I6YvtwjCHW+bkPrXHdbR7OzugBgY4+swpJIt0DdXhZSxubSpemgWbZjIjTXLm9c/
4xEXAVwSf3USofCiGyG5wKx5BsQv+OXnk29eW04e13c9CnPnQdIg6cOTdZWJqvM0
qyZsF41AbxCYTni21arG1EvCX56wqt0UAjqzGb0T/2rj96E2xZxHJaJ05wPrmv2R
T3GU92hhv7/W3ntvz7xPt3G/0cR755OI3jcN4PtuSNkfTNmKrVrJEQtU8mL6X/3C
3axyBURy2+buhlXf2Ts3VNgbmRFs1ezrvpLJiJRe759NjpURwy2usLv7hDTATGcg
Fw0ykbvNyplHQAVbRKGpqnhd+b4BRd/YOHxFeAKq/9/wRC2hLRbVeX05rsiI80jF
8kHbRh+CJvOB1oPdbiQmBM3zgm1TgOpFHAh7EMU/3clDNG8fe8XPjBKlscjjHVwP
GFJtUndD08fLoeSOJGQGM4NC90cwxjoFWsEy2g6S9WK7Ly60SVpaKrhJXq9/jWSc
sVjz6EUD05HUAsJM6DG7G68ujhETuQyKjX1IkOY15mmxY+EgSn3hbH9WMTktI6gw
l3ds/mxs6pNsn6yjV2kuUwX+kM7fF45QKmFpDJRtRp4l//ekdc6FXF3aX0hB5Db7
ZdiUF7EyT2MAcucIS15MBY42PguM/nAvfci1qXamuw8UKnJrrEWJARD5aYfq3RUn
PjCJhlqyrFVXmLCXJ/PJJi20s0djDLNnVN3aEA+UNpgkX0tETd4Uavsv+3IG/mNX
RwdmnSLH8+6GtVt/e31sL/Qhqh6D8a8Glnu9p8yld0UP0rzvDNE/CbBNvGTelrOS
KBtk3Fnhh++ca9xs4MT8QdiSs0FiwXMh9pNdwTepYGPUhB3zDvuoYy3P9PFhiDV7
EqQsMwf/WlIFN+761fU8JsUxjW+oKBjsZPn/tZU9e1DV/dOFXmJ377pTM/Lxah4w
CImk4OdlrpMs5wfBjVg538fjrRoDV8IaKAYNhL+5EfeXg826S08qhFnX62lWKpw6
axVVsgjGjSm1KjVv/epA6Wl01xNrkxJTGfeUb5/oBFV8QD1PeSaz1v4JL4miPPG0
7uzz5Azt4chGIgyTgqIEPgjfzXCzSSynmibVcZQgbEx3pu8b/mZWayHqeazqqd8M
Z+r1TB5Bi2wr4GAHuecehgPog9JLPCAFkfpqaI+fVAi+RLyuGjgmkgd2S2qs45G+
dfF8I9XifYSHUnCMk5KCe/ldF+viUYtXg3i+1yTLoz2oIO1aqEvsu/rd+U1LBBub
4iXQaLrIkjt3KHMNvJl9GahXX63XCrCxaSQTT4uWdXqFfOG5ypu/hnb08kHguZf+
7Oo0P7SlA0+sEjhkpEkuMC55FbfIbQRP2LjxCm0YRPi3xVY1+AmS1LkEVOpGdoOO
Dm9shkeA5MmvDkG6P0ZlRmR/Fsy/CdIyobcpo/Lrjey/nqfsWfS7OmV1cbURQo0p
GJHc0bcSiDrl/WbwWbIfYDaSfw7kfFg/DErARur8YE7PHbSON1e203QSkO9Kfjx8
1+FEY2WeDso8pl6fKolpQ539Y/4HBxAmm4BUH2gnjgiTwzBJVY0hctncHkaXjRYL
2wPUtmDhP7yTqJ2WvrTVZdL0zINXZYxXHPvoRjo1OdlPJ9wqXjDJiQn+yVviavCp
J2lN+BaR2TGaUcCe/5RIFOoMVKGiugnmhJusPBEjXXOUpKxQ7JV2rwPez4bfQmtP
bbOAWdD8y8OBmleQIM6PvjwezmwLMEFqhmR5o6DoPIAeHqsB8s1GG0W6hBt72qb4
cWeT8A1ovHYjCK7rX+bOx4N90jJi8aRsnr1j8DbEasfwmuTPZsTbmowfsDHpuHkQ
AWjL057eYDMxyifbM5reljRjiGH2y1b3D1b08BK9ZR/1JefakhicskE3A3mlEq0T
ChzFcjccT3n9Mnbum9YFFNAm55dmqaWRN8P/DYA8WO4hMtAaZWHrXQLhBg52qpHS
eRcAdgAn9PPhx7rMecl/icCPDRbbSb1Hyz0IphsHltFF0niBNvNxJLpfXk93Nsl7
RzLv/qEjDZhjP+1L6SJflLETUCaq81AzZxD2K7DvbyybxK4g12QF4C63VcNuXtBA
JS0m4HpMsxrzmI7sZ5joNbCZvl+cpeeUandEQav20fKsxL9d0W9RuFaTqsUCEo5p
KPK2Ws5nCBmFr0MceTuFmeOoHoY8bxQa9Ceyg+iJnhGhYpXoYqFg2ntUFmSiRG6M
LrOGBi2wcVut61NyAmmVo/khpcm0ELS4czy/iqfg7ztuz2HhgnJbX34lAOkBLY+W
ZT+WmpIT0MRITcoAOPbDSrPT20zqSjZatoIqFWQjIbqAhZV/pmoI3p2lIYV/W0AW
K9W+vMzbUgLvOJNg46k1DaHUsdD7nskLl801erBoMta5sEnDkTyzT2nEfNykfAh6
sE7P5dWGLp4q26GgqrEYBBPKsaBwAYOfwZMN89XcmrwBh9K0gTf8LV5wqiCxvuss
DzNSsZCPQciId10GNXEuxTiIeurGO/71eu6apQG4AHrz41mi26VBbVwpB+DXpAtS
92by9SuEsyDe99lxAy/nQX+Zq8/E7WUWeOH8dnnb4I8l8Axufgdd4HxHiTMvauTR
5vaah/uhZQIyXCYEUfupUllfOrzPUZdOEO5hqIqmme7O3IxnSoKy23QJyWfALdBb
OIvoQxyWGEhwoZt4MoLbBu8edLKz2/OPAA1UQayVkJmlmoFjfVrQmK3o5fBp7qyx
dpnBria9rnuT5wT0QZuheUT1/bn+GdtrtdhX+e+NEXmPpK8Hfjn7dn531nyc3yd0
ghvOzysSmayOzUwE0EzAuiwF8S1a13JwsPJwLshiXTNKv1KOQHTGNHcdCjWATaUR
M2JPtfT5k0IroHrOb9cUXIbhFTcF4g8CzIi85qz0wvtyw7UuUlJmJfJWl55hR7hf
mDZbjf7zc3/PzpkinBg2xxHBvp17lFYRydEDKtGVp2y16Qy0mSpKBu+4Ly46hki8
oMFuRNGFo4kdulj8/KJBh/dKvnIUYqY+56GNhW0wjUiJtamFJIBaRtzPZAiGtbPV
S2wPUuAqR4ZuMwrBeLf/z7UPdluDuiDPD1huV0taJTu6kSoKEFCOAS/WvqmnUwj5
MgsrPGuSWlGbM5ZI1ajyAeR7IX/X1nroJtIoSZG38KlE62DoS8s64ANh9C0hE6Kj
zm+oTJfVwqG+JUcauVD0S2UaXJjhzz7iyNg5WQ473ZNkdzvJvhCbDS0CJy96O57O
wrx6fV4ZphP+lSOZ/9ydxpDD9IShOQXjflaEq9gniihiowsOWdZulFun2wxfkeWV
nnFo1bCwbtagUjUBpOL8uo5ISfK8uav8vZwRKLGIQjOHfoc88UdIoqDJHGSpuhS5
6mDs3ZXY+0HhJO+WznCN999q3nod2CgzGREgnUGVbyLWXfvB1SOX+O6eH0K+AxYk
lX0VSUP4OimPDG0iOurGpR7/CY66BrAxTR7Vgm7qFAaUqLu2bGHJie4AuXB072U+
2QdvJA00RV/zX2E140OoNRWSPD3aFd6WuiI7v+D4tX3JzM0kF2tyUoS6hcyV/Dpx
FvSRMo/oSP/q6lWig8aMGNx+HHISPhXK1i+MgobjF+lge8G8Rb0kG7TzFk5FTHoY
K6zcS4wyfvXCWayvfD8NFtaRCvTe+Bzw8tg806GbES2rCoi6wll+f53K2vDTr1hE
0MMqffE/G9j2sVtS7AxoYYYdiL9AH9XTolvhRsqtJNNk7KPAfwk3hQRA41QK9mew
r9w/xDq15ww03kWK7FbPT8EMC49zaKZMDi+V1IDURYiBHAoY9Qbs1JnhRloBQ30F
keOClu9Xb3VFOjoeTpDbeywW34vcvO/ehEJScugYGpLGw/gsjty9FOyi+VCo8JLc
Hz5re7OWwRDiRrlEADUdO3O/PJhHeLTzmX662fGF5JQnSslvSFFmd9OpiGj4h1Rk
dBRy1kItF/mZrFoVpr1YYaN7AVB8WYny74gauDJB8C+jwQD7howuLhVLzq8L2yBR
WNcZ4IOIrwjuQgLXklCMjR6iAVB25QmQV3R+86JWiB2tyuIDey3ON/uo8c0pIBLT
pm90budIyv9cT4Ya8pLIA7EI3Ol63FO4iKkLMdskJUBqE3MGNP/AQAu1UUlZ4SAo
kKlxjXuQC0xEHo25KBazv/x4A7/af6x0OSodWmm+/iofcgUNzxvSVr6vyUxuqsvo
aQhEjPoc+TpDvFxEBsJRkAERj2MlTYHCkf66ZaCeTEaAT6AJWrUz/AULCbPbQmlQ
5+lDs80ucx2dfE6dfAfFf3UYB6xKaxugq7M7Zd3rTlJG8p/Fg6UWC+4E8H7cQrJI
UVtNtApoiLtpKGaPXCVL68sbz6yms5ba27+1WnDCQHMKKt7QgV1I0IAdRQ1Xwbk/
o8m+gvlHYGU4AMRWiV302w3S7SydNoEP2M8NX7n7BY7DRZTGB+yxuLsVpXuBPjf3
Ul6T6g0MWP+Gx6FToPDMciGnsQpF6Dmb1bl9grhtzcyOhPkPIU+VDM1SSWDZIegD
T1J9f0x+X8YTFju9ufzY7jFX1Mh0Xc7w+OE/9t6q7Hwzs1u+lGRCwFgab35U8m4x
AtMvA0M5YvXfoXntZUHB0ZztqAlztZOsjpu2Wiiw4qPrRJ1RYlKKZ1UPQGe6XIjm
GEdmvWdTuHa5ldc7865O8h+qs4ECiswUPdcykIdahuUxpg14GTOvZ0TmY+cYGE/4
GAKzLPjUgFUroJjPZ/gvIzUn/WMfWPsXq/Ny/g4PhGtkY7Lv0Pjyl+EzZ33LgNPq
eN4hsfqgIuRkiKuaEwMmw1wvcz7zL67Hnm6VZVFOyMH/cj7uNJRp7IjY0VSTCMf5
I2ChMhDKpWIOCV84OBoM2ESRWE0aWKGCE8Z/idt9giH6mhLkuAYSCp2fhcm9rIM0
Vz5MWv/3D3KHrtXlzDgbv9Mlo1nFVJXg6U2PAjmXGzl1uELqXl3IJqcR3T26Qtqf
7150DUYXZN/n7Qspx54B2xHhQkgMFZ1+JkvINJJqiw1SIEqVgxJyhjck9mRy9rlO
p81izzSacNV0MgwSoVjYi2SFUHjJZGJ3azEYkUgqOL1/6O+QvB0Dy+s0oaMtMESd
/GOHLVILl7WdQPVzB8BQ1AG4mYU7Hg4CEm/ZlaCrQBcUeHv+fqNCVHwrOi1GFAYd
B/pSw2dDN6bBkvFLSl/CZ/xveeLsEQCN9s+Dw8rp8jTkSXe31c+O1rvxSDLjV29x
Rjaz3d1j7lj7KIg5UEHQmUXTa2QQ2L+ID/4kvhtrjArurus/rM/p2eiyK9Hyknen
CJr2c5HJuxWxOiFI3xli4lhxug5JJXP5dGhLMCigiZrGqqsFCUzj7QynkHVeBT5N
bQDacuFLfieZtKX5XmAHOF/1AFuw1DSzP4UTN8W0O0/Bw7iZu+kHRkkAFd2nWvxV
7kjziZGuedkgQcnzSYE3NcD0arXlROSJpMyDx2QjO/k=
`pragma protect end_protected
