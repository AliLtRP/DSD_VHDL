// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
SXe/eevH4Nm7COkUpGKfZ4Sb3tFNOubdlqrDVIlDPFH9IN1Oi6Ixu3JyMomryk1voP58wODlWSNO
+DVe0iu0fr/Pg0kgxtpU8iKk1GIER7lansZv9PG3KqRgo8v/A6aNpII3GGKZd4ESEsKG87KjCAUC
/q3GwkNXdBKzkD9BGQhks5Q++kys2JQ8OMQ03vSKHRK8/eb55ekIqSvw5DexSj2sz1xf7UnBADCP
11KYZ69Q01xb1UCy4uX3VYrNhAH2Ioxo0t/QsWn0G0tQkGU+u9ZTtgxoY5v+K37H5fpbihsl12MR
2ACR1aAUzpnqpwvyDbYhPrGx4i9VyqIpF07B4w==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
+UEPM97OHLQ9s5iurE9MINyASxLn68DxIC0SCO3SfkkJZ3Vd2KmoH4x5xugr7chv6ONV8db6Njn+
Tjk/rx9c6iBo1mnoC2LBaYv8uQ9p/RbDvcgN67LpIpKJkrcTKBs7RhHIm7LZLZgwKwa32LWO1cid
5ziOT83XCj8iNR+D5y3mOk8Hpo47dgoWZ3yVoBwxDbk0DgkA1CHj+PGecdY+r0YEpcCOuf8uxvaf
qzPRUx699gHWAYl7QvvJDdRlCLKYacF5tjZszsqEl1mQgB5X1eIPH0cXIjNXndlFOJRUJ64ts03j
ZmPe7QQUXYHVbrewWgYfmAyoSOAmwK+psWtqn3anftqy0EtcHhVQ3ZEgvufzbtVBBGrQ9LvAJEfb
KCvON1qC08yLaOQTmTafyIqE+DP9TIMOrOw2dVmSQANuWwqbKw6d1i27LCTmVy8KquhvUdZ9Xj30
T5SUtcGoreDWlYG2YkrVZ8hrKOx7Sx2GiTGZeIddV4Ep8KtDr142NN0ZbljNsbuKEILGtM8Zsh9/
umqNxggzD5wfZxR7c67k7ZkgSoE9PGICwH9/6OIGv5BuT4p4cgFhUpj6Y7eu4ykiJdMzrWj3dr8c
RJrR1iYTKK/sYCILmyXqGhZmk1fOsk4f1FBMgvPWpT+W7Mk857SC/ff71viR+ld+MnODs+64Uzf5
xs4ER8gtM2FeM2VUgbyY2rAgWljN+m4JXtvLiClKjxIpEpJ2ceSEbA6ijTE8PcWCL2KOhmX4tqSA
Xbu55akf+PBZFy/DHrMEchwsxset4y2rNLEFmEcDaQBPsQ7DCy6jmT2rnN9XREkYHTL1iV3AiHSn
gTAhjbtBlms7fPHlJY2JrOXz8xgNr7dEIVxLDY002nFFl1mY/9n+lbH4pCNO0ul1Hk8e4lxQVlAA
D6eU5wC9BHCKXCikDm7GeWIQnJvOUR1Ubt69tFnrogAqVcJIsTUgMkPbWJO9OtPI0CxfuQvgIflL
vrp59gfLPGP1zru7imBY/PXbSmLrkBC1bL1qkXPM17ALNvfZ1JUTRj0L7poQ8p8Aie1dMcA4f57C
EMNTy20gIpd9Tb9Yn6fGAvhiqCBMJut+A/p3gyE43O5WSDvqijt5RQSN04I43e5+o331fnQOebj2
/UlUASMAJor4sKUgm5hWTqFTFr1IR8OPIQOP1qSXm/Pcu4GyJkddmU+y12aJz3WSHtOUXW1LljfL
cwziDL2Q5lo9ypoXKBNTYNmJ2K8HL/nzd4p2qEazYmf62XCwWajvHmMmEKBUEN2IfHRi4UrfiH/h
oynPRe1JWiAAby76M3DKdk9WaqXSNcJPH2V3cyQoeVyj0kYtdwVGbjPuDNpVnl5+GGdKh44m5jKv
LIvzBgnAdn/8unW3wTI1KsPe4fy6u7eA4bKYMRJ1REumZj6kxJEGWCtAM4uIenf67d6OALyyyNin
2RqYWiv4AANWjmgT+x4p/Dy+Krv0+NPYxFVOQc5s+NfJAp6qiXjJToJoQsn+5I1NWX6hY4+pfQOC
DrE76DPpyu+bzrk7gfvdgdoAtWvDr4yopSHnoud/cjlP5+NRh5jGU2cmBdMNf2UNegZmUqcHEFFl
sqwiTI0iChkbnagnZ5i8GnZ/cSGcdKJ1IFwJ8dUSUvOtnAdceT7WDgu8r65JpoyC8tmr+/WU3MvH
7O6qyWzBOSgoB+cLN8bb5E0eL/LGRRYj0cS/q3EQer3liC0XhpOLkWhXnCYFw8+LC73hRNlA8DQn
CTvklcMj1+OQNNdM1uPN1VrIlpQ/DvUgpRpwpqyhLmVvAb1uRFr59sZDRI55P1UWiola2ZndQG15
Foc3gExKg8xfaSZCTXifrPv1Hsnj+nmvT3+9UHVq45+Uufq3IbFyJf6b+uPygJ8USVKOc69ZxZBi
d92kQPXJ+iXumTV1k/wxWPHvfvnAhbDna+tB9vCVzmXYnbDk0BmW1xoKOKUG0jDyTucLdiREv7q7
pq2oTXGnwCTqRT85ecBSDZd4WNcAJ/JMKYxYc17dcSWZulx9BZhm5S6OHMjf/Ok/t9j0eKTd3oGs
lO5IP2oZ8schEUhCuRTeB4onyrBttbfxvFowBWLuiTRYQqVZmYYxmIAyILfDsjYMBNrwcQppVDPl
gBbaMNuogac7UkjQluXxBJauYkcqS4imJSLSULn3WrCIH3tiSxHkW/Dk9wax1Mn5YyFEfKl1YQX2
Jq+COwMhE49FYY5G7wscIVomQhLALdxrWpC03yYS8vKCx7yVlIdeAd+04TDcc9qjcTX77XTCBi3s
VVTyRm/i+/FVUTpey1t5sOWLWaXv4Socg24iNDbCRSYskt+O8CKE9O7+9sui7GfuaVVuK3tES3qD
eUl+pcqK/+v+TjnZdrAi/MdZ2WpWBBQjmWv+UzxZJ1Yw/vPsZqY0FzsBqmITY+16t+3NvJ4ucw6P
Q8lyAkGwA7GVUxLzl61drYvN9quqXK96mWBuDMgUVHPdhx+MvzX5dxjb/+UkdSEkiCsRNPxsYSuF
7L1LT6Rhl0TOn58UGGu2LubwmLFHY1PDzDXBQEH1f3j/s2qWzN2UypknnAo+C3gAKKneusiRhKO2
acrRPx9Znqn/X8/kmHJQu4a8qFJDY80xRsCXkpDO5bA/FvRXq4x3TP6QrnjnAe+EOHGgeMTAWLA2
Holo7uTEQl5NRrQzF9CdMXOce2ATX3NSxYJdlGeC7nlEMnUrYcGwigL0bxIWbmCXIrdzTgX1bP09
ME2hFd9GN36YDiU7JP79KutGH4eRjzIMscqQhz/oSQGzy5nYVbGowXvdWC0hPa4YMLvNZsM1wJbq
wilA618+UXAVJP6SzfVVcA5JuB39YBesl71WL13stAJfE0vPOnOQDt9duASEHyMso+vM5Z1HzCwH
j2qY326ir2/3U3rb/o6C9OzjAz0sAZe+znhZJwgDtkqKDUZSCGPAEr1Hku0V1i8OwUNczMSGDJfs
UrX1JAUBWRVRP+U+PzAd5DjNsXgG7DilKfklU9ZneCkwBUcjRS4zeaD3nKh2HebqMs8XxwCgxu6M
NlaNgAvwNCVw8arPJH2tjxUadw80keBzK2WO+rS2tlcyCu8eRypfUTaMJRmlnXJXI7z+JbD2G3br
v6btkwrroJ70peKyLN9ZVsiCEvSso1EHiVBKYLvP1IKfX28FpS9VeyNMC9B0md1QcITQhWYN8XCP
bwAa0+nVW1LfH4u0q6LSoJUnogCVbO+8qkIPQGhHIaTy9FbOOokmLL+iwkXGRN5UBuG4IFJaaH5h
tB/I+upd8Ok6IhvgUETzbN0S81x0gjSWIhhKMuPZM5PXeanYIchigK3YYUEW1oPiPIrNVwhabv0A
RChjTQ/IKrFrnBhRlHkLspSICowpKOBx31fy89KznUTLOMnDJdHXVm2LAWvLCpKstVVlBNiV2y18
TLTPBpkRVzOWHGoXBeNTouzvwm75+QlehT6bSLUzlJvnL2cNllNMV5N5ldLQV8Szf44omZYqlw9s
dEWQf1kGkmwIs7xQw+5p45TH0Taxs2B8oy9qwxoeZtNqllTVJIDWuDBfVd8wbc/sbjOXbekIni8T
CptO/fRRtCZg76V6rCAAS6kx/VNXy6gi8pZxQe/9/Tc4sPIFx2EYgzzEZ6cCCDxjejCnA/oXXhUH
9pBZsMBih+3L3NNMuhq0DqEFo/hsA2HIx/oCr6h6VxgUTMG24KIo4ZowsQWW3OxKTpVRyRxcjtNa
IieL11wjC9sFHfdP1n32wxvzVWIsNKspe2zpImm1pHM0izZ1yzg4bat9HjSiKzrBYRNZIFcYKq2x
dVRsSEnHdwZ6VYjDWhUROSR6rNfv/MutOyBFMKXwnGEedjedYaHZnaOTHJMvCeVBd6qPIHXQ8X33
AW59quDqu1iLgafTFtRzlFtCfmaD1P0Ht7x5xywcP7SsclWl15yaJUT4XWXGwsPaPBPZTy3Pmv6N
/TpVHwqmIsaEXlsvh8ZXBTQS6nlzhvpV1ffgIetC8LtFUItqZ/89E/07dCg6ZyH/wpGj0KUXGazR
fi6S6Ot6s7rUp7UJXg4prfzeT2VI5cAFTIeUP17kM977QTKTi0aT75MXfApA7s++0HGks5w9C4Li
BY7FUwSsZL67E6OV+bxosCvXXJ35FEbyy2RyyLYtTyW12kiANdsye6xfHOI/8Uw7V3N7iIdFGUSG
lWH0W83eb8JOGGS6zJPj7pYlnOGa5+Uv7o/jzfWw7WPAfGRT+Tpe1JN/RZiM7iemDaytCQQqtmyl
/DruPE3Df+vfwxnX1XQfz4OiOOm3ms/jL93SDxzws3lER8yHLUZq5fp817WtSKtrMsHnsz9OTRKA
J2OFiwLHl3TdFmF5J6oTmjU5vZubFdT9pb4+uW/6HJ2DqHE2g7d7B/cSBGnHEPZo99APSY6uwHFi
+gz6R5wyMqa1wR8HXF6RS0oXw2ihvpcOeuWOn2NWgyPDNIILFWwvjOtQMQ84cyVMBhKzBfuV2NcG
gOCIMChQISjbW7zeqL1wwWWKLcubMtYo2ReUOxV6vYg6TUA3uzFa4ibb9Th+2HWnZ6/7F3q5wqxF
MCSAKxCHWYbpf5n7ARykX/BimGWM3RNrARAjW9yyRp0tRFQA6/KjD8ieOF5WIs4oxEPH+urx4E2X
emi1nVkXshwwHvQbRorPgjQN7d4C7FfhmQxPMn/6YizMHK6xvS4rwhpJrxkePvF1eNv/WS9CS2iv
tpdF4d9jL0ZZJqCScr7oWMiy43z09vNnR2ux7FV0k788zaPv5719mgr0ZMOAawOj1Mrwru8HJN5h
iONuzANO6tsN9EHbyn4xXnEbs4mca6Y4gQv0otv32TzUAEa43ec7RsBBFbygPwdhW+ZsRgzuwgTN
lxgefsrkrQhXGbrSCAfznu4Mpx4sgbT74zvy9YXla3lhVePpRDObtFftHMYTvJtAhmsjEt613n3L
3dgas1PdrOCPeUCc0FHtYa5WySNiZ+C7lQpjOldgJRdJ/3lHPJYNP7k9D2j1p0hKCBhW+Qy/bOkc
SfvkC2PVG6sWoMq4CSGD5+9hVXifLNk0A6P+vrDILt+MRIjm4QmxXyBiVpdKR/RmQJG7iaEtSrJ7
AtFh+EErIG+zEVNvaHJfNODURDMMZ08h9YHbEQpJo6WhAjcofHLJbZ4KsRrwU+ByV21iR4Cz93kv
3vmDOHkgeAOZguvckK86TLHdJBN+pVaNFrlm6JQtxSP0JKi+KIsV+7yt7P8o5IHCwZKa0Hqoegdm
SYYI5uW7IxKlucASbnppCu3880InzVTiYbxX/nh5W1CLHNE/w4GHAit2bBfSvzqIN7q78U7HL7Ja
2hJ+48S3SrkHTLR2XXtZJMq3kTPFg05C0DLQR+jsj8i6aQzMZZ0ceXO0z3kCoioFfvVxSgpeGFdL
zPZPTCaIgpYvFTkNYjQl0RwIff2MxLO5kjABwbimup8zsq39zVH03w8nDCbz/4Oxn/xBrYc3w3sL
6tOpO7stCUcjcy5iz1GsggFjwPFj8ByEWj7yi2WLXookhetQ+oSc+l+CmDXZPcHKvuo/8I+GJ83g
DBqe/QDjLz2M/0QTbIlJ5syeo8ob1Y7yWiH/LYhZsd0XdtP7oY7CQO7GPhXeuOYgz/D0JrgDBbQt
NwyHB37UxCNfOkV8io00hm9rmftfz73Hv+NV9VhUdq9GZbirT9BQURo0DLEvGqfl1oYj+fZndksW
P59vRaAEvU2Jj69pfT0YRBCqV4lW0C9diEhQj8p5qyhglwa005dguI4Q9E0IsLXL95v6zETdZyMX
GJM2FwYda0FiWw5vIGUgPGN1NCGO/lX+7WkNyU7r1FlSNsfMOOoLJfZ9hLebra79LlJvEHxtIzPE
b6ciz+NXd9Uy7+9Fmadx3n3n1fOuevH18XGKIqJgUFENwdVQTRTqDDUPD4eG9cYmEah9lt6t4JBC
srF52/RiauYna99+7XF0ytCAtAnLbbEk9g6TFASG7vAITi491PfUZtIh3qYhuEbhby7N6QeacdsL
fRSDJnwq1ZlRPprRE52oETZdQrzG155VbDrHxSZyB4d1fGIuK69+w+k95/VkujhWMgHR9KFt9gPG
2ysA9lrmaQ8l5GDSh3bpMaEp9WDWyagJgOVPYAqexaTcvodXgPtdfDsaBmZ2+4cBjU8/gogdhsjQ
fuzGimS/wF6mBejqObKkE1Zcde/nY7xo3fj88teO1x6yFNi67nNdYP4J+fumL1LXabmzl3yM0+4J
EE5pZ0sFAwz2eXVb6PxQ1grQpeeJGoQJQmVayHd7t5GYoS0FWuivlQ7UhCSAoYKF6VIM5i9L4vPR
giUQlJuH8E2LjK6RjsbPdxLF6GpUWMqRtJF0fyhQhi6KngH1d0OurjJmHS29SE+m2SRJ+GPGOypS
a+FykVE05CDOKoQh4lD4fzpd27HBjrBN0m/pBA6vIznskhelIwXVY4y1mU81qhV6jDCJlNDRvjxT
qeVGzox8XopH5fwiGjPeYH3hZFscf+z0Ix9GemH5B6Uqv4rGqkn2J9E/M0n2LrvpGzsInZ65ekZz
P6A4kRaiEyIHIr0uz9HWaG6eLeL6+/TpNSKAFi1PfXK8e4ohES4rj4Tm+ERobYVwNd1I60givBuT
6WiYM1TmHq1eizC1fQQDbVVhdRMA1HHT74eM64WXRCD+LHqyrwJHwJSs1slEWcL4laMFrjSOvUsW
X3sE+j52WPrSUIbyJz6tYJRwe9NmKMK0PUjARqAddrjFgv6S4r1EJ6yIsJsHp5iq7aSO3B/aZkr7
PGlhWWMXGSicIKxTksDNkW2eCckuvqZSIg8oFSl9/Mj17cZCCrrXDYuu+Cc7/rmhl0oLmb7wl2CS
gCGW8UFXap0fo6IngC2wMb28FKL4MQe0ocplujbRT08dpkqAfLSxXYoWr6cXgV3vmxF0p2im8DG0
ZN/kYreCPuPrLQl1pmxIzMvRt6qowvWu9txv3tp1EmNb1ViGOLhjq/sNQl9mOXgZdxLscg19P+M4
fDDqv0YdLNb+wJanCGJEYkPKai2kyIVZhRQspbdzeoy8lBn8R4vwTVqXkb+cJacl7N2HvSC4dcZT
eOUY8fDgRdA1f4yPobtvIub0ccFguyZY8YCmdBZ2xoZQs9Gm3iH3TPcDnHzsgoPxMd59iRzwZOpe
BGaSSGqSyqB2mwFFbrAnr2h4Qy7tUuiu9b57kFnLQy37mU38lRU7H1IxEMVqVR0Z52fZsA92p5BX
tlxzeDdVs+Bw0AYAhXWc9DwkP4xo46iiKnUYZwxhsaHNsMG1w4qzrIV8buJ7Sa9ONUrHUkWb8TdW
euR17Lh6Oc6pCGLD+hbHa9nY6XhPZFfcbi+E/FKDLY6IyUE51FSvh/z6x6edByJwhBURchi+I1Y5
G5G6O2G2Goe6D5/6GTa+dNZvLVWPJaljk69pqEV4bAP76WmG5Jn2wxyP0jlMMM9FS+va8qwY96RI
9pOW37DRdKM0P3cSwZQtJUZNhgTu93WtMzROJnnUvz1mq8ea76S7E1bdXacFH/683aM5HF2Nj5oF
mF6lS6odn94R8Dqfr8CGFp6B2DKr0GXJbXjruh8anqn9uN5U0zB2y56Xu1AaD3Q+4IRUIXm0RPad
NyeDcVDvvs8mYpq7f7Hmv8Bfx/kTQZxDmI7R3tcCfhOxugAZbrT+bcGI7ltlEsOwAxIF6NGEanqB
NyCZ2tZc07DpcI6gkTe9YjFPyFU2x+dOaN679yq82hjZj3exPMR/vugilF+ZpgeDpOfiuZ1+kKh/
mkqRctY3snCwcY6fUOZIWCP/7DCMbTamt34CpYbxbAUx75qRv5ZIcm/WIpX3n3XB66lUZBrB7DRY
iPcap6u7d8Q579ddpEM/zf6xCReLjRpQPrL9CWL7TRCuPLVc/JjA50B1WXbBREel36OZXv60Ub3L
cxZQg1ca9/qQ5xML6BIb1/2/coAfSMtvfSrxPUo8Kr4+3jAdZRqOYbPqGYc5wxTMyvv7chZwlOQN
HuyEhvBSuR6GL6rVvzgJ4EV89kD4+bdnSkeAYjAAxD1+PylSSQSvikyRhMOAffhww3nHQCueCCqC
N8mXUtInndnmGOYYiVpU0dg/0btEQzys5eiPVJ4y1TeUat9VOppY03kFrPbz4IoCrqsAuXqYpoIM
bMo4WcGSF3EgHzIK4VTnnfkjcuYHC1AggXiR7xnfKQp2U9taIiZYfTzLKOS5+aA/yJ817YcWzZqS
Qzbz5IkO1KM0cCs50IjnvhsfI0K1aU56fh3Lkr3ug4B3OQbYnEFS4M75u/ZWlRbm9ixxtG7hvJRu
d1/p+m6WabJb2+MPYEAJDQQr1Ijus/u1mAFo2v1XE7S3fHpiudAUuXJ7YO+z/cBCC9Lnoz5gDeXB
EGK8pox7ShaLV8A0rYZYkUfznMoQQT0uFL7x0Ga80mF81pNX2dFW/d6KbVMqClVRg6foSg1uFI44
0wZsnfocO/QJmGZTboDDWZ7eJsJs+JcHyzn0HQBhHGV09/w6F2DcAECKVZIMUqQh1WnhEyqtW9Uw
1nKpsMsgDw9CsXfyoUYhIyHJWBhC7lGmvYS1E/q+xXaQcRqqKrbvTJpnGXTR1ILjOoYawt6DCRAz
po6EwTzLsLIIdMGY+7bm5QiP+s9/uFNXiTqi20CxAvFkKTlzSqPkSKALi5g/lz3K570w8zsF0xHS
Va8TD2+NHoGQjM9v2xVfKKHfp/eTQJnVswpBjbmHZp+LKzp+Jtv8Z5reZ7n+cqxJz9KWmh6FWTKN
YuxoSbNTEWjQX5DaIvSFmOtiMRGK/eGya9vzmgJ3wYwzEg64d9gFvQhD4AvDIH+8TpezfldeHNH1
Hus8xg5rIkABC+NC8EUUkusY4fgcZbZON+5dFa9wUOriDUzTxuTFx5S/P23FA5XWVvkgUB1i7ysR
dc1tvdsMzlHDmiKL/lH1embvJjBm0Tuv3sfgdWtyzoXLm4jduFT0Y6dR13kbNnx60c7gHGmVKw0z
MrNR2Ev8nqRyoDPq3MZ+wBw3J5Q/wiTbZlLje7QSyUnJ8NjYElPH8VVpLDLGyehQ4qcAXrtJiCO/
yQkGO8dkc/0HIsCD9Y3PodLupV5byDEMRPqyB7WGa+lE6D2F44FA4eU9agAKKAGggJiokemRrqpI
VVCaE+DeCnLLRWzMAdRLDdQdEtp+Rz6722jxj7TRg6A9YgPfmUnnrEsy75ESFSTv5Le8SoX4L7dx
v7hZExVA12BXhBzB/FztHyxCK9HlpZeCZ1luM7eNE/gv7kvnywDL+pkQn4FiCBFH4WeHf4uTCHas
X8wqSOcAsBbOUWeLzig3/m3NQ9g41GLUOacj1LsFBCuCyT0s7apXlnCMqj6GSlNP7xMAk8WvTaWd
MipWGw6xjCfliXX5CF8Ucq4cwtipLpEP9PJcLgTOd38oVka/Zio89KRuReR1Ov+s69E9pfMe8rnB
4WexZsT5GmRfTJx0DnNfl9xOPebkZCpl4XB8EYJgC3IqWnmDpIFLXsLN8QNTgRVHUn1dvF9pTyPg
UOfE/Wu8sGTtUZ/DaBdUI+whxnpUEE6JTeir8UTPrR7vbQ3n0f9yTTzDUBN38EsHwUPedcAUftxV
beLdgoXseZjn5qD7GlbJkCqCeHFOBH7wU2gtKPbNNPmZjk1OuOzL05mRLI/uddOkhMv32cKhZti7
gvrX5fAMrTpbeX25LOgIwFIijNzHWITIRkHrVI8L5USlyN/J2ktJYFlzkOUrd6F8tW9axcBpjlFh
cQDp45Oz5Lmx+pjsyhCoHW6I8VhKY/kcTtdLFo8XPc+DAXpz16B/n8aIU6pi9EXmyTHhbcXeQGsv
IsHoI+BRmP9lEt1MgvJd+xQZEL8o8RfKAuJWN84Mq07IHliLoedzqQVWPQW9d6fvhVoprqaF8g1y
VJRsrK98xOlQ6U86yIQ2OFAlFwZMoe0pfTd+tZptSiNYIWBAdpoOQKkwwf2QpQIznLr2diMXPS40
tlVHAJjjOrhyAvzGKgaOM9JEg2ge0H6e0QPhg3wtvpxFgcHoI2rD9cLmZeB3YCDVlTHsivKenX5F
jtTBfR5jnMh7jjcjx+ibF4idS9Nz97jN3DK9jojty6hHnPoTWUwUYd9XWyNAe/0RXnOB6F/Mrkj3
yEwWB2WwlFTz1yk0x3LASn4+InqCfzV04GcC+nERdj5973UoKpSNf+6Ry1t/cGsiTiXdK9F7wlZe
QTnrnSuNbLEsqArcM+p8Kx+rqIqqDCV/OsbwTjOzV9T6I31dLjIk7lpuczfz02TnhTIImVWbYe1W
wNRacOjvGtRclLbGBVd0tcGq+mGAkwdsmzUV7FF4uDoE2stlTiTlSQ2CyzFRvUZdQtBG5/kY9yzF
owvW17XLtzv8qr73tie9+ik3ap+XVM1ZTbeZB3JwdQRsQZtgt2dadSsaO1wQLMWj1ntsvZh2tmoj
70VZGI3k7wnDgGFwIv/vh8TPM8b1tNm5YG35WY3FfTJHbZQtxwQCq7anYVT5GAJbCBzdxeSR/Qbm
ytb4tTIMRR0aZzYp6j7d2XkQfp8lQHGgo9QxvYIwx/wd75rn18CEPyZxVGPXUAuzfJTb2jaD1pX8
jb39nvcofmK01CUOxaJfjplR8OW5hoIH2VREMKyjKhIT6fdOwScAVAf//peM58f6yLCRwtWLzOFY
OZXdb98rHO8wTT1ozx+u6vmT2RMdqH4C9GG3Yn0YpwlgX2qBhQpPFWq88csBiGjx2uA/GQzvsYGY
263HpvoZtD8wZFKu22VffQ38sW51tePx2Wf0Rp60Uh94QcSR99+AjWOFCSDzFzW610UoVJtEFLOe
axZP4Izs8nWEeMRe5hiC7pUB0t5kk85LbrATu7pnQLUtWoBaczP/lJlbtzAWudOJrRYsCqv2YSy+
0RXw6gHVmeMuInfVj0YPkJ7qndnlDrhiotRJUrbWRLlshmQVM3ZS/BJqYPfOZM5SdvVRtaQUQ7oB
Th0KveyNjbEQBQHlqw4tVXae910hpfjh3MLEzk2Xm1Sqgt5y11F6hdlnQRCvN+mXKwJIC4fPYj8a
eWJEWYOKmesopFrLW1G8Rzuo4E5FBjLYc7SgIetEMLLaoSq+bJGyniMCC8h+TWpIfBP795WybhsB
pql8RPO/lopJpMLvSz4C6vdd2x7JJByo8HVsFxDlnHGbNGqUObjhlJRmkmglnY7FOOSq0BdIC6rQ
eK4j/rkr6eechEbyhHEfws5J9EBO4thZTu8khMYFpAGF/4pNHQe6TKmYL/tYsex20IRsuTdKH3FK
/sPDa/UDAVuQFPWc8rKfzo26Wk8nIqrQH8jo1SwTfZoMNZbLR+oDZ+lGFn/fLiEvHibc8PtVdwpv
jo/MsuI+9R9+fAmA3mE9mPLwgGilj7Lji6k3yNlUvXmWCIKivCwXYUf5m12FLV6whYKaXxOibybP
0132197D3x655TOLzBPc+EGbgC+0YAOq0P1VLGn0r6KSZ4s9fqMHX4dTspEV0yDmFdoKD3ouzGpp
vViwdfeoRaWvuCKVC9t95CI1oT6IruedWiPnPI2adqE01uxwVBXkmiKxM4Nn4H09RhdS4XB3zNb7
VMnOHy9Pt1zBSgV6eUHWrNqAczRMFyvd+WXcNoLNMNHCZG7nBzeQpqIiN562HYcAIfffuJ3cCnmQ
8+MOa1TyrHejeFaCtg6a9EY6i7Zx+vZt/fVsxs78/sTIfsW4KE93oSIgvqQWiaLdTSUp4SQYfAVM
WSQ7Rga+SjfboNhY97yh5sUEtkEEh2SqH7EUHjW5ikR/rOuQyzm63l1J8cgVH+X9a9+QOQX6VnIu
Zixt8CP+IwG8dk7YFiDRwIW7Qt8Pso8hKWkWZLO/ZVVZcsyFhLjZZNvvbBOrVSuH6cwyaUUOvovv
vY/N2ms3vx1utYL2cfRxyATmSNIHttqiVZeKZh6DB6GdjqBIdwjPelDCVt6kK6py02Pf95ael32B
kAPdIG6zp3kezxa0YmRhkhAROL/l9woN7Ro4d1ivroaUVDzbpERjBmrsHFmPihg3BCrxVsbpCpD6
a3MCm8LFrX3JLbf5cFCDrGMhikHSzS3oJuyUCF1QY3lDlVSry7EgKj0dw/9xhqA0dkS8uwoXCGMQ
yUQd0qpOVjmTqlhbEXB3vloSIh7o48JzW0/jIespP2NIYEXYmbPaBjPjj5G6ZI31TA3ZGLE+RMJD
sGXP4K36pk1vaadw42awFFgqW9ybvrhrwyfkSEqW4hT9Vdle7m4l8GUA1X13vSu4RcWgWVVOjL/S
4N0iu4m8WnewStHWFa3EuoftA4doxjAYQ6gZQf/jg5qDwCI/WmeHauSA2Y7UrdbZj3+mjbqogbLn
oQFD4MOg4u5aVrSn3FYHrtZm2VRmHuu4/PwSJAeGCUkupLdhS3moR3MIPxfSP/D+1UEmkp33vGH0
/D3suAnL8wPh9IJP/feWMuYerK/SK+p/aZtdPIHvGmlh79J8epTlBv0piXf4cwBlocClGaeILa51
iiMLORn5pZhKrcY155FXzqaHGZEe0l0+NZCe/t6VFcmrHkHQOEr7xeez9VGrCxpsmVeSz4DjDn0F
fawsOGyyp33XQWHoFz2BO9x7ZA80eMvR7sYnMGYHbcARX3dbCTU4SucRi4CT+VDKyyuPHg5Ux3Lu
PaU0GJZ04a6FBSXid/3C1xPWuviCx5P1++U6sT6pAlE6LBmYiffGxMTyDlTZqOxaKensN3DP0i1w
K0YXU1HSj8Ul7RkMvWYeGdQ5Ko6X2UDz2OeUnI6QHUK/rwvlXS5eh64GHww8bx0QEQlu6N0vY/Zg
vVa8VWFZ/9woExJ4H+fJfJZrLUDA6U3/ztowFe8e83kKiggkfKL/sE/Tbvg9zOcPUuK4VVzLxfZp
aR27WwuJrV5DvsD9axd8koQc4Bx65yNva4+7op/SR9nwTGgP0k1g2jA8JPRTNc41xGPxoSyxULWd
nzmFmsY/LNjhZUPzWxgtfiWm2Tpi41Y8jYL1OZonaQ//QuoU9r0UQtvCAsirgRTLbcMJyY0KKycB
l0DAtTfrxqz+nLZ2HKEw93/fJrFhXc0GyG6WKOW8Wxc2ax5+FCJO67XYd1nPw4l8AfDT9s6dNwXZ
9RJdIxyDzU8qWLfDI6Hae/QeqY3z3WuM2JTGtEz0xjFNDENKNmjWadutJFtWGub6VudHCT1R9kMX
WNnQSH6gs6QKSrD8qEckUq8sPOKZ5AKe52Fl11Uv8BXnM+9fX8C/gLGWp1PndtiW2OByd/cQ2JUN
GNzg/sqCGnQ6GAP7rNyFYw5Av+3R0SThEbodeptbpUc+viGzTo1TxKAU4kd/T4LSaBFphHA8jDvZ
xTVHEUjexKEfDpkFliwELx0HhAYGhCPHlSj/r2hsfkqv4oN0h4lBrLjc4cz2ad8CEeocK+tJfRwK
uiLrhn5tWHF8ayHCLUlAGCl4t9qhDLo41V6TKctcTgsNsbtCP8Tqxh690q5tyjJ/En3ttkFLa6Kh
8l62SexpBlBP8OVp5lJ8eV0dGLSQZiiYXXoh0CxFDsTlDcwmOp3bHc5ePLER6S88pPyb5xvcpACz
jFtj5gCp/W5htoPyJnETFJ1mnEWqYjlanFpmOVoyj2wgfsj1AKJA+GAVAj26mu/mM8BOlV/qR4cR
yhd5i51pXIN/4n+HLursQShURNjnGx4vPIIPblGe0OcSPelGIbOomEiir5aABNSvTTTr/YNnLLn/
VyGshaTLt3qppfCdK1iyY8dpyWVvfMolbaJg/a4G/XwAQWKnYs+GweXcCd0MDwQZHEX9+HqzjKyp
YfwVABq9stwvsNv3SHaJB2PBzVv2yyVJYTfMtiTQ7l+IwEOfS5EQgzuOfD0w3CfIq99nhGY/ouGU
/9F6OWzmvr9f7HDhptLjWv7WDWXOk2YL3Jb+ZTBvz6alkSrQ4fE/jw6N2BBxKxwmxbQ5exepY9Zv
Pb9c1ACRT0eZMPtoh8w8jdFIQLpqZLsFTTUfMR4xTWGMdCuLoligaQTfF74sbkIJE+ufiW7RhJHh
0gIw0X4S6NHvMRfRyjZLbk1wjXw06LKj1S4PCkeqpsAVTO1m4z9GDMiPPLfnZshPjf6RAzbDazDf
kr0adC6BOOtgPbijUqZdKM9D09QljkeXSOjxUaeoyumH8+91FpDZqubJqJOE+QGhEczM6uQJ0Hot
kYSG/r1lVIxWN9X9QUKSvbwMbpiUpn0d7t/Imyixh6hbZBn+RqAsPlNX1bzn49j6/1vvP2qOdjKu
4Q/zLxDvJuJnFKT4MapJYGiaaTabOCF5+eixZ4snwikrTscqgRwPgJvuEJse0EBC8/yE7i/jSaRt
/dXMB0FW6Kp7uBXpOdov8UGjtlXmk32c+aZNSXdZfoUgEvDtp4Cl0f8hifgs6CtH7bUEUBWYfeD8
yKRzMI1aT13Ne9sPzrmOhJ3wqnFHSbrZ+5Q2TqI0cFYiDQ3uoI+2iI3Kto0ER+rsG6G2ewI+VrKS
3sbKMJfKoagSBoNJEdLgP+l7fXSiqs+x5leIpz29xMYW3DP9SXnCMvXXvNFafP0/qp3TVjkxKeu0
peICPRNGlcR13jjHCEhQSVbbPiS2AkyhPPXpsbF2eEpb4abcFlqFuTPLJHFFPekdXR6a1RET5DVa
vljywHHJ1EajyBN6tS6QdklqexYt1fL1f/1a29UR3c9tjZUXb4fu3YoSEQ4sj7/wil0swgjCn5Mb
oZw6l96aDWjuvwWabEQdR4Rilaij1AVgszcKa5gH62CLWQ9yf9GMMzJF+BNiFOV7up207irOn9D4
eOIftT4Dk/alpTtj5OHxel7zSdfoPd04kG2Sop0moBgEckMtLgO6/UNNqayvG/8o3RQskEnRxV/0
rKmVp/4HnXDawGXpB/VxFW2MdAXIue/dVOclxmfCgA9mMtWL1VKRGGw/8ZzAht+fmDe1UT5engu/
B6RqQ3M7b6KHalttzTS63TPkl3nMS24sHhpOhfvic2SlD2t7xexUjIuYr0r+Kq21CmnCfJ4F8Npt
sVZyO6VvdMbnRwHzRhEjVFawfs7qJPKEjZMEXgU8fqryYs33ok3JTQQntbVWjAIwrcJJrvG45fus
H+clCpCK/c3O+M3UQZF4cMK/rXjND5NsvyCHu2tfArdi/+OHaLLcCENg3GFd88i5SUrPA6zY0fit
CsEj+r4hTSyVma4urqkEdfwSWmgwFwvXfxY1ltgHZaskmHgcbDFzJ1uCfME87RmmVAJXQZYkIeOe
ywUVq2LhE4C4h3keTzBL338evXdG28wSu05Y3ACExk6Z84OHTSmFFcqSTlPcpAtU0NzCVAo8sZC1
gpEOSWLxQEa3xkhHa6t2HxmjWCxsOrP+WCg+c529gE8d6f2iELqVBaB7PlWBlxKQNUeiG/lkzE51
lu1+u4u5HZL/TdUBdXFXJCgRmlstTQ9IV6UKWQYqQN07xZUB3v51s5N93j9FNks2x3WRW44p4tF4
Ui4hdWS1k4oIF7vYCPUt3PduHcnlQaj2mzvLcQHGpMsZle0bJ7a6ukqeZUp88+POmngAydSbsLHF
YcJYxikWPbB5LRI8J8oq6K/YRg6TzOtTw9TYaOGhlQp0PCnmVjmHdpZKMx9HWUUqx9GtjSAaHkeW
YO8oyQ/jHXPBQY5YKjmACKYdFR+i7NBmQeJyKc8hHAwJZ9jC5w3AjW9EJPZveIvhTTaSc+sYqF6K
heCdva7gP4FuPbmGFlWgIDgf8U8f9/mH+Ixtp/2bN+zympjtqJCxp8FYD4bbOzTiayLQ0XQWIFu2
AJBFKiHdzf9eCn+cmXosHu3YK9I5cQ9AAHSQHKkQoneB0TqBmzKLrCuuwv3URUdPapHd8bfgvF97
0X5XaiKQtrnmftdYKVRvJz0dvoalMuKlt1oKSRhlLscpLeoD0NPD3fjfddC3Iu13ucXgBpsvwfmM
nGceEVSKBVg1sJ9eXepyeG14qTTJo53nCD/b8ON6refDRDjFJSU6r6D/c8YzjijojJHCmaBAVNkF
DYs99Re6Dq3cGyRLxKmBGKEnytl8648cNwgNyKBR2Nd/5ybSXgtge9Fho7IgCsvktvPPPd9aig87
F0OUiEcG/14abNm9+gDVzHr4+UOZ+nCjUYu2eFPo3MDahn58rLV9rQeE4x1VJJpevDtRD+C4wiTQ
mYMvjSTpgTWDUOMjySSHXv9KdHBO1l8bG2PyHNTqw39ptqhfpeF2/vAq4P5lbulrW/sfPPqSxbIQ
ZBkZ0l6CnQ742lEM9Wgm995yLk1WTUV/mRluYHjuRqOT6R5ucZldN24zjWy5gWX/JNgWpUQVjXOn
HPJ5DJePZRxfeNHYyk17A2u2LlDH/9umW+gN2enzp1bjM+iN+BvV4Aez14/rxALT4i5qJ3H6zyOh
GyVfpg2Oat1/msPaPKY+9vk5APMp5Aeg3YRT3eGU2ENnJSGeo8KpjEzMvSwyUu5Gfn1mro0ZKOup
H4+fjUsadD/XIDJiU3Zo11VLuKm7i2Utuoz63Sv8s9v7HemkhOqEuzROd5Nns69fzOVQ+SJSPnVp
4Wy3UKcNlceN4ImvVvgCoFfvkLgM0SUmUJJa1T445NHZfxehxyPlYc7auyVmyMQj2M+gRY0DEOj6
878naKmsX/qDtU3j5l407a4AdyUZ5fwMnTorYTiwWYiJ9FFjwn0uMKsfEGcvxcEUPDn8fLa785OP
S4kPZZmQD1EUWoYAwKOx+Jl8s1yes2RY9Wpi9UJh415Tubfd0efy0BivvfKXVuYabIYnJaKALVWa
fFCvHuuVlg/ndIWQw1CFtN4DEgbCFWqcVD1OPFgYsoGBxNRMwhkWNPzpQ5g9jL25mxiomcJz9VKq
gpB7Uixp/8zvZ1slGUXbnGd5P1Yavn25CiI6H7Xcjk8S/Po2J+RnGzcXPO13K90M0HLb/EdWOXHp
4/7gzMl87Hrvj0iIpsmjq2i3ujoR841n/pOQ3cVCiPRswXIRlX3U03ihUUXiqu5CQR3jgUGa1evK
aj77dBShV30h8kmBNFH++fykTsGgI8/+AN/3AUXgPEZpiXN7clahJaxeaPJgMTxUC7VdHDLYtQyu
RXwONEyXiqMCJbOdlF1NEE53WJOvuwp+/oXxgjrAzYylP9Fq+eP7nn/b1TJ8jnm/lliWhbp/gszo
2S2zJ73mVm0Evtq+zUvgkBTdlWe3/258YFERO2/oxtBnNX40hoMeH6y3cyS/DYl2KNRUKiRB4Y3Z
frJ/+OEh4CxAkVm2wewUWovDVN0nuHxZ4XddV6X5+aijBZZRuYNmNmxfEHz93gTvgfhvASsd/rTY
b4aSvf4rJbAqEfcZQ4i9454OJWBLsA2bE6Fx3j/AazvSLPiWVuYKSm2qiowcbEhFm37NWJfDglq2
ed6fhugjC2VzgJpwioLHj3HFly7FIu8N8B/t6sngoA4jR8/J0z9rB4XZx+l9miQf2xulOPJiwv1E
J/lpig/Vv8FthhqpQVCY5Zj+M2kuRTxUNYjlpvRt51eZhdtJmZUfbclD+aBNQYBkBi6gxfG6DsU6
95fVq5Ng9QLHzJEP8NQkYxhbWWaWCtcWczeHlH8EY/MPE4D8nQdrbDQMTVO8gUtyo9ZIhpPOsLNJ
CrKxAJgC9zL+bbrhkbInJ/CAf0jDhN+KbCyfKh/QEED02PH7drRTkeUWQHTtVX8KSJPZg1QlIvmN
DZL6emBIqSi8EdrPZsOqdHscG+dHgvWICz0EPfdf3CT6mS3wy6g/7yliemlXQ2eA8H7l+HMwjgtK
iHZcmcQWHG7W3WVpKRFnubkHJiKRiBqfd+SQym043epOALPA9nJgFegDe7cQhgIk6n/+1ofUmIxd
JJCYomxgt3ScVS8aPW0yzNF1WEVdPFNAsGr7MFMOqzKYlmpkTaYGqWrP+dXeQF5QQMTTPJVmOePV
Ab3KthSyY1S2B9SZz7bIOB5MOLuueMpv2V5Zaf4EVQYqIRoieWKcTYHj7+qiYat4rOxshHjNQWpc
cJo2QODtbyMAufxUsTdfGAzCAXEBMSUOr3+mW0MeSePHegm0QhirnsMKloAQY2jm591L5kA3eb1H
bPfAAuVilcxlQEIFRU1ISo1zK2L6veKK9PLwZSa8KduBLA5Set6NfCswOrqwrCvTwWLgGq2lqwQS
4br7oIQMUWrBaDFjhg+TevoDRWuRmsNJ6Weev8CHAikQuPsA7vLiMmBkUK3bxOIgzl0p/BEvPzEO
L/3A+KrGpbRasl+unw5tsE+6hbwHzSLslkZH/QB0aDARlSPlXOc5zXzI3S1cyeu1fIaRgJx4AgJo
XifU4Hw2JJZzkayoGUyFiJQ81Ix1pulewL2thuoy1XPgw1ddIFb6WK6QvkOonMeEpyLly+breWxG
m7iyI5QdjZHeQ4UTLCayYEyVk1t8ah257++zd2HE0ZmP9o5EyVWjDKeomdpiNnjxK83TvutWMfBx
TgiHkFP/DK0qHHJkV4cArlLKwQlIPi9zSp1ecP160SWnloE328+5YoF81/H+NNjB4dOmQFYLPcRA
RJKhHshuJ438RLrB+Pc+OelIP6Od4VFbX4QXw5Cpwkpz2fhWhlLMUqSB1Lua5BqyehX2QD5WDieD
8ReGQiUZ5uv4Ak64VIlEmIpw2CUiu7XEKtWoVrDd7myf1i+tSSYHtBuzZk9rarqFaJXyn1KZhlil
+0Cj62c9uFDF6EcrtyPfgeZYYn9cpfChLtdJQND8pbU5ZTzxBtHmf9t6skT/Nl8Mq78UNMHLeYOZ
MuTa4sL5wK2RPXKRvxngtvvK+vQbkb5l2vAsGZSWbCaX49JYPPPD3GNdPb8wqj7kGlRCQxb3YwZH
dFijna7yVes11vkk4UMCUxZZPAG5y2a1/heoOX01UnRT4KxfixrkqxOW5DjPhAd5qbfMHm14qhkG
Op/F8waBTu4h+15c7spZqdTiyOWmwd6X1oZA+azm5DMAUPukLEtuws3rHJ4qnfbnCN2tfR2wGFd/
enJOoy04EFscU3ZmTIjQoB6K8NuSnPULSbQSyLXjEd2yjj4Ku9JXEtxMGBlSmb/hjUjVBh0Wa0Qp
a90xfS384YBCYlTwZpm6o2RUA0KB6JStdeXus8iKPCmozMsTQi5x4vYaFc9zaw/b+MCLJ9dLrRXd
UKDmQR6PZOfyQT4S9ZEj7/r12Zo+ZjynM2WR5OKYvwtpRM/dq4o0bOO/FMHk/pIdRm8sjkscc/4X
BY5GOOmTBNJzA4xHBmI/AQcqfPPeCT8uoStjj5/Su5XnsIkc8WiDPzGY0Gclo/eVDXpWVTgUMtVz
cS9OBb+QHI6MbX5Otu8ZHhkMQa4cOVHGq3a3AxBq0gdStS9JfkeTBhemR2PM/kMxdQ4C3bD6fpUs
Ugk9lPEdagUldp3dGCvfb7vKm1hm/ay1xoUEh42A8qqSm2rpXCG0kZvIoe5UzrJ1HLb0Lbn0LR62
DQ5BJoGiseYpk9LjS2IaY/FQ/tu60L9ysYigg88wECW72kW/TbCl/A5qE9AmvtYgWEZ8nR+luX12
U+4KWMIqhml0Kq7/Ydwe0jVqVjXCLW3nHQ5jeIt/p5UfhEMVYaI0IUyb9EVs+vHnI1rbSiF1m7vN
EaJ82oK4rdAhtqaFiE6HjKoTYCP6DtUbe7ImDTkBoXPWu7DRZ3YjZ+OEtWeRcMvZVWe56TGIFEvM
pWIa1lR8qlBcYOKGAyZvI8zWZJsl47COWL4Hsp1ryfunhgZtzbwOZ/oTqoSCCBlNFzSZscgpjNdU
qMf/K5+KSXwHfHIxbQjOYU3CadJPohQsMKTdwmQSkemkBjkNtc2IBgbwedwi9oDvZD+1twJudhDL
Sd7gYW7hGPJ3TiXOT63OsvE8grvT5I+5/rXShKikwky18MQSMo/5nwtn44fdQg859Hrt0/eezH9t
oQt4MATi41tBggHpftDNrd/YFj5Xkp5MLWMfKYKHX9qoki+J5qZF0cL+oabTuX9P5QvP4ZcOesN5
iDqR2Bc6ViT9hxv/l/JRvxUQnIBYn8pCd7T3nk0OoiELuRYbR9nrPcacmUEgSixEEXQlOI/bL7Ps
tMmmDb44b7CdSRQxt9zhDQw0v3JltCWoWPBI87ms3v1zqLPEfMYXvcNOiqDI5Keqq/ljHlPbKlFy
fzEY6CyNUyY2TcYLZJGapNuO9DJs0cuDkV8IArJuW8lX7Rq33A8RzvtnGaOaq28u0YtGqh/t5Fnt
N0QeG2Qy5+eR+EEE8VmO6KJfUho9/1QR5S/LdjxSKe4iMzE4TrlOUsutE/RpPiyGUP3J2qTgUWkw
xNAZuCKAPK9XNm3l/TNJdkampQSqL0IvV5GmguKvnNwGjZoj9T7Mt6zvXm4rnMjnsuEzZPrUGpGo
oqWpsvHR4P/bbZXh2dRwlUr2oKKTaIBcrvgByZO9gCSKFBtg9MTT3ZP+X1KM+B+4Wh9MAu6ACNJ6
dD0RKeC2lQj/8AqJzYPqVcH+SCUfwtTvj3nUeeIldgAoCGoq8w6neqEHhDRXjznQ6f3m38tE6G2D
ajimDjbp7QGqbCItM5x8QbpJhhxav12cLFTJDU1wMjKXYVHkhduog0BbjPgvvmGGCceTAN+HKg0e
j6YC0VQVShGmM7Z25f65OMJC1USaXd+XROiflrPNUs1bCYx6pTdwj+1CuqLThZd+QOHLVm3t1x90
smsishkzf5d7v9cEzKt5SxTa1S3KkRqVdrc04msxgSjP7k+hFGOmAEMzhl9x1X5acekGrzMmvUjF
aCr7hJCWDyWaVymqeujDVW4D7YuHOnO7eNts2ne6zPekFYZlPXXvnwADnEwEzXSRRL+noZlsy3K2
dBwkqxxm94HsYzqyWQjnwyuGCfdnuNIpcCA1XyZ26t16U4CvYqiAyDJA0Ca5S17qzExoofBG20UF
fF7cpqHs8IrODb2pQWFIIZ7zLqXsnX9AmiKQ/0oZBMWoZNv4mK4V1S9hiWBbgShYHoubdH02iIkp
G4wayvAR6yUdVjN1/3rbdITbJSGqOzsMiYu08XXOCcjPXCvp4omiKxlu4XxlitnjM8N4Zrnxran1
ZHZrQx+CUv5CRMp+IU+wKh3geFdY4t4tlWZylgeiBfFlss2DUJGNEy9Y/RH3ajFKZ0BS4Y1OaWNw
berKfj9F4ymSn3rV4kdqwD3kxpF3nmPWl7SO44u5oX+020GsbGvsgM4L7r+yO02g+jK72iEWTwh2
uOIdBrWRxuiEr9qCyJAuZP3Z/PBFsip8z5ocuSXyApverBiWMspGThY8RhORyziwnap7VGLTbY8h
8qCH3w3Tg0xSFdSkoCfcnCKXGUm9abUBFtGHK+6hpwpJMnq96pFiJhMcibtvqmTzjMJSrhlK0dG2
DwybQs19HetAIzK+ctreegbf1GEWGKqFmZ/pCGwB3s1F+PWkJ9GdORzWrqQeS87CCp66QZxy2Epo
tRO/h5G8bNn9VM5ssv1g948gbxXUZb8OyPx12ALgfozed60UT15/bzByl/lI598nDWw2PCR4ou68
5nOa+cA0+5dqYQ74JpOsrZdRXqA2tZkpS4wLBkG74A/IuvwnbAeIbLD669+u1x2ivp48Np0CzFyw
H2qVUAaUvzy+QapBW9G2IBJmfBZ+CEX1BJPWy9MKjksug/LPmvz7/+Q6qFKIQteQBGB+kOeyCqzu
S9wStYFspSKPT5EiHp3Y++5KQF6Ghd+18uqxs3i2bvmCCT7+3XaANLOv5yi8RG7I6ZqaUV3MBw0H
k+z9d2+xsmDUZPdnFbvd8++gfcGgaVUPc97Sf5L7u3S32QEVFkX9nOojgkHAf6d+AH2rjINmXxp0
ZmfSJTw1wNAF77dXpGvy3K9pTw3A60vAEe8Xo/4AFsJFGV/BsArrvMRtSUK8dhUMN3ncDVkdN8wZ
RXd03JMQrF4csXJan0EGrdhjghsdMrz7oOJ8l8/nBBIRzK3X4t0A5HbpGXzPDBdG0uDn1XLn9xy5
DTSx38/1VwH2qD4grKlHqQwghMZTTtJoAETDR3+uX+erN77OM8gFMBaz1fruwrHegLd0TEvx6cFM
U71zfby6V+vGQsqVTkQjAACGW9vkrzVW9V0w2sbAmaHSlE/OZvJbuyJoOmf5IONdm8yOvI80qCB+
UcHlzUDoPy9XSt6DfJI3mcXkVc/JdQU45DQvnuMkEF1G6MqyUbhDH/9XJIrIbbk5BGvE0tClVjrP
l4zeVvHC10ypALTICYo5v7DhGifO9Zcz07aHIgrlhFBvVuhqA4gMIMW/M5G4mWuwAGGzcbo3Hlg0
WnxhlDAszdZDTJJGkZO4Y2j/JBg+s4ki2K2Mrav4jRkkNUl3/CUTCdqd2rraCzcvtGvTxomc0GMR
+NAOwApATwlvUZGvC3pq+nBv+rTDBg86ibRov4Wb/oiv1tgkW6bfY56zNx7wkmnGYgYaw/CYcOXH
0GNVAT3pBr5uGjcs2GWCjtqcSXV5+nRIQxvzn4XRy+y1/qYBSdiSStZiZ1oQ5rDEjlP9hYzMQEFN
7vDgs5em07OHnBpqwCm86I8ri3b8T+/A6GXeIVVR2/3it3Hnhzwa+eQDPcD19k+fWKRMMyIvHOUk
zCJc7W4zYU9MnKbLQng3f/vTWYnxwj2KA30AYcP0h6q5lkh5PNfmKlmmILT2jFv3/13+M97VTZtX
KibNLZDaRDSldh13FQ2QmvJKnah3gxoSoL8XqiWj+A5326AsPTqNL7eESIF1GB8ContAEldxQ91J
RE2XgJdNC0oBFrrwAmujOHbPDY3genPgWjytbhr5UOIQoyt+thC2+bTlHr7cinXHXVv+KsU+SbEg
R2XVAwgUfjrCT9NZ7VDMlLe62p8MDmuYK2Y0WL9FgPa6fOpOM2stWdG6dvhbLgPkHqGZ6aE0Y0YO
rNPn8bDkd9thQIt/OQNoKjTLA+GURoH3beLY4wZI9ntQQNX7ZY//i8dnRHgFwSamSkQn8MiwEGU7
Or7MT+bJP68rpZSjjqANB5kyr8CwNCOIgHVT99U4Tqi+UK6Rq8EuVSbUSD9KVSJltZNY6HAx4TjD
QNtKLQrxK9gdG/TFdJ3JKE/gQzdrrLi7Sse267v1xlzXhHg4m96hqVCz7yJGbg3C+DwFABhffQrg
vEXvZt2iLX67Lc4WWggOUN3NVzd1r0bn3UZksLH/YM7alCpVRyTcPYoEBBi+KciRgBzBD0ovIu2h
TTo0JxBNnh8BNd/5Kzgwo6K97bGLtS1FR5gEDgaCNKWzYGFCOrkv8B1jHN5kGRrWyu0Cev7obaDX
MHxbx5qrGbXaB7H+BhPUSekmo2BmdMxRaL/qJP7UThHJMt9PEqg61KaGk+NoDPx6wFf04sy0PUpP
zNiJtXJS4NxJll0JYeQ77bn7WcjypJ5gHQNqhCokhXtkBmlZkDH8sZHQyMtQTTXWyz+SU5Cw+GdM
Brqar6kwnKnMwanFfoVgTrVs0TQc1Hs/SqE2p3YHKSH0Yn/nuCbpzmHBmxHMOBa4j68jwHoyu2qW
1x3kzaAFJWC9d/jiaSiwRJUI7kKQHbacpdnJcf9lUti2CXY4dUQFScAUAehp7hiQ6DbfpIEHIhNW
K6DcLgPCNm4EOoDsAaXr7q/tFoVve+JuHkb4xC7ymAVQey3cEUxlnN6ykmo5Bpxj1zi837KM+oQ2
E2NsvFY2W8wIC/H4kyVcEc3w2ts+cCUdSr8pT64ql6dJIq+/0W90uMKS57iGB9FglNh0En8+StZX
VTHMKCeNooAoGhXd8UQkrE76GlpiKY8lxvMwVAXs1hVIxEeJZFNV3bdk7lQmi9O1sXWFhywBvphH
YPsRVK1HpBVNl7/rgrMG2MgEJn0i5MDOE2GvXp+lhP25hLZeyLBNvxKX8Z3C6VxCXz771hK1nsTM
xXbQju0NHtn7ecvJwOL61p4E2ZMA87elHCFaQxSOrrZuNxvCXmeDMY/6p3sPYvLSeZ75VnVzuUbY
Jimtj45YrFBPsYE1Bwyp6rM7/9THQVewPWysAEjd0YEx8Uk9shgdzPAB/Rt1UmgmMQCtftbdRPo/
zZ+vKS3mHF7G3S2RKo4FY5ND+vLh8A+j+LtbIVdBTeSzQxqODB4ehwtXSGFTwvR5cP0No1wXu1xF
9mKE7sUc9nBuD5VQ9mPdZJvivDIAAJ2XwyRFiazbeweM+o0zps9rpdTFLGdX0u0thf0JJoztZNPd
QaYhr2WhaK40aHURr89c+109TDk+GpCXZVCjUPXQ99c/v8szjDDW1orHukgnkhlnO35BtR5MrG/B
onWliaTI0B0yu4siGHYdONmeaKV3Ad02iqn/4DPy4XqTDCqgfbkopu1WwD/M0uVQnuKyjoHfJbS1
qkjiF1hQdEO0OBd7Z44fu18l+7YujvTFsdTZSTs0Hhh7RRpzsRW5vEwvSVswvBDkPOXWa4Yp/oyE
Ec+x9mO39kfagfWJHMMY5jzgOw1qqlnbw3mXTN6mfW+s8i1WW/HDdUAApedL/xANndjxtmVsjhvX
pHz4+TABHYyff2G02f065syN10XhJU2iG8ENxSZXlk5GArAOWWN1Dy72GYvWjNKXI1TdLPE11PMk
YQA/vcrzgwxki9nuQrlCIjqv4NuK2Z7OVsFd1dtCD30eoccOfzUy3FRCCpBa9gRciTBJOLHT5YC5
qD7hwuMnE3kvD5p77Lx5b6DRMB9FP5B9lvDR+p0ptMODRfFDND7P+sCm2DzaneZK8MNlkbyWByyc
Lpvo04d511IJZw84U3mETQwFlOAtPBHeJyQC8RemsmkeRvL2K3QWOyMoNvaFt94zAdVe/X5vqlcD
2EOQurcD4hxRdf3jBUfkGzdqqD0b0VnQ5vZaZzR1yU4r5Y0Ws+7WHRwjR6IbMY/oedu+rayxALKn
HqKfML2CylqZ7GohWf20XeTXp/igciK1uWvNB17Dw63iEJhw+YyCfokD2NFy9Q5rVpWhQLFfk0Nj
XkuGr1uw6nwAY2cI2yxvV5XlxvoI/lR1wYPq2t1TrrTilGu7IA3ZhDNEHcyYDKiBGuTqPkO2TWcg
9XXneEIxX7e9Ncc0KghCL+1IypSGfyNH/FvquOH593KG6nl2i6JkHfjrHhHJFjDngzlGCPiYQcoi
kZXm7rp4mNH+ZApSXKdevPq0ehJ/e8TukR1Y6HFH8CmfZA1AGK/saBGhFMYSFAE6L1xMroxBZYwR
agJPtmO3FcpF+AkbWmYj697vHMBcI6ZyMf5P31JNSeqpCKizOzMnGGGw9t5xdSdmpVfpNae3UhPo
qUvQeBxdiPiHZ+ctJZEWPe7s5KjkGJzsX5ggH3YA8whWOuEMmEQ9NIZYbrh6hjxc+ON0I1hLjsCq
FD1wpzB3h1pXz3TIfB1sLK0d9zK+O1sdSJLm38kgwpRj8tvLGoOzOGH1cYMqe6fD/NxL+ohVQCr2
VkTMzejrIk3mqYQVETgwoRNref5ueDL9UwtzqYHUfCuslifswXyLZdZq+70Pz7YxxUqjo/+g5a/S
aNhOAbn1lSW3PymLVYIvo4r7EXjbQfGemkxsL61WX1I8mmtUoQroL27Y6+4kBvijbyitLZYqWKB7
1z3gYCwmY54tnIuBz3cuVpYTTQ1LtOLnuMvk4R2YQ/yZf3D4jsjk0NWlTYutxSwonvDH5OZsK5yF
+SrpoZ1McG1HZkacuUHRI+7hYfXLkaIwNDSQm6FFCGND7jiOBaPAm1TCf05fJG695NOin5iTygHZ
Gl6tiWnLQuu9Mr81M5kWwYgPI1m4sBvMjaEajCkkoDauAmDjX1yH0BohwF8S8D9OOBOwMZCDS0t1
fjqEAFGcA84I1vJ91FDDcIgkHFHJF+LwnnYxR68kMGFmC9LV/xcwKnokmV+2LGa/zfzNbwR6OD5K
i4tt7XDYt6CWcmUJ7WtLy18dOPOT6d6JCx4boTEKjs1QrTYRgieJR0wuBLmwPKE2nPPNDYmvEihl
eWlgiQB134pEI8z75b5RO5OgDH5+dG32UwQJk9QILYVxsyw8jCJh+dj2t+o7ryHEL2bYT8l0iUPu
FalB/RMG2wQ767Z9QTkzv+HUbP9HCJRwn7XTKWWIFMrWbnlY8EW+jGtW//fUAQdLR9zKzaO6yrnz
af7hqYOYXqltwkTOkFXMxi99zDdjbnndksTL/vcs3q3T/xN0C0pEaPAsXF6uoDwTkez7kLo3YDj/
/P2hr6lrdXha7hyn9bnTcCoagBit+MGFKFsXYkhgC6rHp0NyVULLMJq5fE9npqTtBlrYQy9w1ppj
r1n9TLTRNmqe2eod24Upgw+4nvAaqZ/mtX3oPyG2NzlRtjK5ItVQONxCPyAZOW82PeniALqy5Buc
GIJkhpAbhEOOLm+Ktry9Fa379eSSfkZM27xZXluFog90embC0upDeTZKwFNGmZYPho+jcPJfsL7n
KT25XrrBm9ws4w3c0xEl+W5LYpxLbEt9MDl9BWU5PowTRknqZ+Z2q3whmoX6YKaZvwYd9uaXN8Bl
06itMK4vcaUQc7geaktAShH0YZp/rQLe6PfbaNPyUjJmbboAg4QJH1nYGBmsne00GleEYIW18UNT
LlRr2V6RwjFS4HFBWKk35XpXIgK3GwD9ONNyvXVhFq59SWNsaIeEBR1nX+QDOhdotPz+qUsAdyd6
9Tq0Br86OU/uul+QFh6IaaE8AXCyOmX99mV9iLndbMARR0srk4HE/2iLKNkIIeQiGodE4WNmbDjT
Tck4DWPhoPQkTm01N+TExZE12HNUN8pCLnBgXNhHrEQ+p3USc/tk+IcscM/wezqmGqv1stWWHByv
c6pivDO1cW0P6QvgzEg2+9cnCO3nCDdpOf6kcO+xbDvF9NlK7vILTYrt36vx0/JIXg3/DCvShWap
tuNTPvgTPIurO51rBCa5CEOcZc46edy9Hj4CbFZZEGN7gYhKy51WMJy5GKzzPGtJoPBkMgQ9Y8FO
gxJjw0S9bx1AJV+x/7L88AHjVJsYm5M16GFe/5qQld423l44ChVFFChW+p39kpS6g/RSvAGM8oHA
fo1yahcReh0LCAFapN5mi+z8x2jguv52Oc9mGxY8lqD67SxT6XCFovFF4a4wol2tY1kE/L04oj7P
24nI3Pg9/eXYMDBYjDjWLYXNVrnxbio1HcImtYcYqLoRv41zrlltzc/rVhj7tjXTXreMPMW9dSrX
5DmYhzJzsH/m2w1t4aZvVyTN3bDPEUDKeVHCByCiHowLhHzvNd0T9VAG5RiGvPZOXYBDtyujQ5SH
aBjO3DQMHB0dhDsMmJjGy8x/XTcrNwtS3GApq01cFKHOqVS5RC1QYOASTaSdw34nf+uDu58Ra2VV
isznIDRYMhZoLBngf4wvfHTWZd71GQIFvQ+s4ul+ar0+eK/4B26w+eFpNiK/cLLg6Ix3wFmF3QW3
CdmcBYpaE/O58tHE+Wz3TAFza5G4G4d8FC1ot8Ne0YGRV8UNVVX4QsU+ih98G6kvHpiJMMSDrgPc
6qoWt+8CxxEvwBgPjixeUTrrftHNv2pmpcbsA4ct65qL8XsUUDDDRYzmhGs6zO+vQdB3t3/qCy2c
Fh1K5ffLDyHj0YA/lOtOGD9BjRnO4+FoYW9QqLYDZL3ls6oX7ErGHLNwI4s2fxyXTHeLpEC5l0da
QtDz2UIAwj269g+wuuJYy0F5KSg63+bF4alAoS9kYjs+3GHKhWTyqR3aVkmzyv5YULU9RWwhFhPn
EvHQxklrQKewF59kLer+Kc0fBd2hygBpfa+CaJplXE4nf4jg6Orve7HnRZLMpKhhQSEhBFi4TVh7
aGA6Tu5oUn2am3F40wcNM0rGgnyXxV93Mqfr+SkgzA6vVg2d3BphlnqUD/awVa8MpXcm3Ka0CLzy
Q6z8h6K5mZI3YbIhM+/rDaKtTlgVM565mp3p0Ti1HrElbLOj+LC8ZUPI9CKoam600byWTMS9Y3nl
apgbHtlPnbi4Tro4Y3bIX0VPxWT5CrxsN/SAlQk/k4fsWjHREdxiQZMhHacUI2APeHpX6wL4sRFh
w4MyUqKPvwhZhaaUDKMbeoiC3+h6djIc7B0W2q+Ioe0aAAaE377pg8V5JSI/aXUcuSa3rpSiwuqI
ZBl8RgEiSqzwgM7vh1WBdDna5WL/EfKemggIiIm0ygrFz6KHYA48uKTBBGmdKmGUwKUx+UXmaLmM
XGzEdDFYApI8UFU04EnM6QhtvPzKub5D9v1tPg20YCpqBfKZ4RXHiZCe8spZUwLuffX/miV+5VtP
uH+0wJMHfe5KBVvrsoiKUw1mZ9WLScFZPhlNT2AqlkQR6H+MYz4zFuuy1zTAX+1hbJVelwJ4gIxm
KphPT/GmRh+5GOguEEH4/W0R2dZRAk2RURs/uTgtIQLyRLqOfl7GvsRUVyjDPpL3Jj0Day+Zs+Em
ttl423n/yk3xa7vXB8ubpTPrlROmji5y+wQIVBqaT8EU1A1HEO6+VXOtc/A7WkR9de25n3FDF70W
OWESMQUok0sepf0tGyzCjf0gv0xDjRzpGFlZ77a72gCfjvip/ss6m5m1SJUb87R5LjugMsCjLhFZ
YFfiEGEgZTx8ELJRJBeYhx0hZqIopisM86wCdwMQj5V6XoobJCdzcL1+8Fg9/RsaKjD36Y4BB2Bq
d+ao2vrrbOpTfVyAsBKccYTA/INpx8e+A/ghjbcu0GdyjHj9+7BWUcqx/sR7j8W8ldmg/dsgmVRt
72z8aR1ROwQVknMyqrSWCi5ZpqM8qr8k/E9JbUIpVhIHF2lK+Ul2IWF4u99fTnNck/zd5E4l8TPy
9ABEja/XTZR4vj93jABE0tFOYJ2d0ZzH6uKeRAJyA4cnnyPM572rYFDHze1X+WWesIke8u2JvKh/
VeLhczfGhRfjX34qWgXvbdcAZCZxqyxjHfnRQMlQdl39ibLWGSMl6Qa9YrwRhszgljwoLczb1XkJ
pV0o3+pOT01Cr1/EO/tZSBzQwasvvtivw1OP5WF3JIWxXNgUtt0Zz0C2wqMMzoL2/sSlBqyfTHwg
SxyMQlcvpBHTasVgI15V5U4Fkq791uuKamYMNTU2cz2qKVNAag9sjJEOqH+98Z40U+C3uOmSh2tq
P7gofL/GiZWVlXLBBAInjxVW+JrxDHgz62YCnJ0tkSlomzEpVJrQ4W7hAabLi82Om2tRqGqlTi9m
fcNBAtkxAbhMbs1LTUU+R0Oxt0wQzGc5lj7PjuhmG+CiatWymF9qwhijnE3ypyYpKL3YLXKzvH4x
lpwqoCvxCrREwEOAAEKgWjEtSI73ZY1tLCPB7fGvBWE7RaHSQsTc13q2XapXyeePjVsSpYNe57Bg
GC8mNwCYV7YFfPg1p9r0yhgvlAfSLkt0lRNcZkhwfNCEq/GtXRfJt9+vW/0M1cxSBJSv8vPt/HbZ
voU7UO0R6ZuNilBqaXaR4agI0HO8yzhKN7QdsQHMLxW38W8K3+mhIMZ9J0Vwqpkb6UK/nbKMiwzK
o3BxZqS+n8q9SO2PcwUS2WjFiS0uagyCyeA87e5dqkAn8pitPJTZwAa+5DBgq2csayg0nUASaC2x
K8z5BPVuobMagkquyJMO67jg3UAd8Epu2zBonjit1T+GddGGJENMIUlr7xcZvOzLb2wsyOttJnyK
iuZpAMQlkZYK+3UOHg0ZbFwB8ZU+JaY5UaGwvxiSoSoFVh4CUp4SkqwYO6xAO9sVg5UHrm0yQHFv
hRuFFK0VI9/dHjophNOmC4LVhxlma6KWvfS8YT8tRS2mGPnV4Y+oL0UU9/hm7rWOazZue8zBPv7u
5KHYtpNl8iRu3WQaorJOEqjLIlVyKz3zABLfv9/gxBJu+bMtimmIkkB6T/a0lhEVQC7KDrz8hV8y
i0Yfo141DYq1d+oYy6avzeqp7FdI553dhnMx0mQfqJ2ZMi3w/ZO9cdMHTnJDkIBHVGL6y5PZAZvr
1ALs0TN6eD6b6Og44B0wE9SIhxz40+pSa0PhuBtnPiZeU2hzJtKpqaZtE77DkmG2Zu47kMX1KuFp
x9YtTrMb82Dyy0mfHFdFvpr4+wsxbXb2zE1EWn6mTFZnvC3M5E2JggYPyQWOCl0TsansvWBR04Gf
0Dh2eS7vy4hIcD9Tol4ubL+NL5xO5CXJ3Z4Qfy1TgVzFmgJS/FHCfONUFhvs8djsKV81d0D3Sksj
pEOkKtoMGShPZGopwG2Xdu2wWPx3nvmaFCo6NyjJ9W0AyoamoWb8iQBaFOdrnh0wzvCB+iv00EoN
heig9WT7WaIq7T2IIO8PwBE/YTHiPPtaiKkacLq5jLfvQX6DJ477HnAV3Xo4xvoP4WAZR8L82ZMw
X/2Pxo97nu8oTIg4Uepps9BweX3UDrBb99vvAZ0wecMme7RBkl/Nza90OdzEKcBVwV0cu2uuBD8G
PU4waeevnoru6L++KOwIl1APEpR7EqPv/enYjiGz8xus1LA2gbLFlHQfwD30tE1Gp6/BcQuYDzF7
KjAc/Ovk3oRyhthuQYYpdVH0OSUIpdoslaKoPc+2kCVUn9PejOOdp7qYDbeMqoJgcwJYPZIw4Csq
odrWXbSsvfMlPH+CqBX51GfsDMnCBgkHImt8dye56RRQCDIpFZ20Z+e4R+1SgOJ4/jD+h1wJzyD8
yCzoztw+dKRqIkcTX2ZIockIsB96oONs27wkjon/If9gAt14ldoRGahBYowogq2jez8DE52S38OC
9GpIl/NB/qO4D689q42ZdzJVFbap08od4Ngp4N4lQVCQFIK11UTzqlkzIWsnJEtBb0Jy8Zk584cy
Il0aA6jI5BIWbZYeHcim+sWmM7MjBy+1sjbenzjQJ9wuQ+/JmTHTSpcS5ngM+bKOltMyIvpBVi3Y
yFZimlp6j3XfrASiB9dzd8OpxdfgGpWp6XxKKbMmamjc8kolQEQ3gUA/WN5cbqVNfbGBxhYwgB7K
XzdQnWbNunye3a/0N2YZhDwrf/LF2w62vHKNhXWP9tUB1KQhAZUxaehnnEiP8C+gH+820a4iYCGP
PZwZr8ufT9F2k5XuVKTceHJhnXfOpv8S+a7JHKTWScXIqaOoEyzqPUKUaEeQGqJMlA/YSjYsPDZ3
5CIzqVDavcpwUUxlFAoRC1GrVXrBtrM0ijKErgk3wBc3zE10SDdGbiT6JLRJuSZGh9T8vDJVGKLE
QQdKBKBL9RLgf4q9MrKV0MMPCpgmF4Ix2mz7T/vD2hILC2T8IGc/A9OIHQXyruBsv/m6ScIIHiFj
bs/mTfnz5BP2VSrOrw9BmqZYR6KpznII77lG3VsbKYd6jP8hjw0igFjI25VipLqPoNg3SIEjI0gd
JfXgWkjiA5QubrMpikFOEWyTA21+laP682XCq7X3GX+kmWIAjJ63uF5XFMCM+w0FzNijFWfaUASE
qU5iYI5e6XNfz+j/lgA3SKeEXCgZhUC4zedf1apFYlDjHTWIEXjDHXDDeB26+YYOoiDJt8bzQVRE
Ad+GhWu09r1xt5/ltYiqejErKN09/8OvnULxU5NTTmxo+WlGxfYn+HZUYiEWpfvC7t+VPQcVSF3M
8WnzI2bWuPGKfheVDGC7yQKtYndZ9wuLKm9oIHjOiVo4QzS4edywuJp7U+eNogB54VSlNkH2dwec
1IqOtlBmWgYSnYf70lleam2DOvS+E91tL294oToZCJXaPRRI4Bd4IpBOXgKjTDmL0VB0tZiO8hCI
LraPalDiA9gl2KCOU8JsuUEm5H3DWR+rxpUaHqonozJyzsWu2vbYlA7kc1QhjbI2rsNLJQxEy6/m
h3EeQrYUw/EWuzawtxKhZclyDLanRUWijkkVvydA5UJwFbEjIN8KCiYNDyG6UJYSFzlmHFFI1ptw
2kwVE5dU8XGpLmdmZUikd/lfxu6e60ODC4ATeG1AHl+8tIDmmtJ1VKOg1DdKYN52IkccHGcU8WOZ
3SVO1Xhtq+KToDcCS3vCRzE9f6zCXs4nXi+BmBbLIgYnLOUco3dGraxTdXrJxDi3PMVOoPX0Ia1Y
uUEz/XdRblIgvdaPiUvQFuUURtMfD+0FJ+KHDK5h5NTTP05a9ScUz7dxQLTTB4g7svzKwbo2xags
TLK3I85jr5Q54VU2SK4WdxBOqJssFzhNQ2xsNqe24gihLc1wfWKPIjO8Utn+bz4G8EG4NM2kGYZ/
AEjrJzVnacYAUovcsG/obZ31aSVVrktse3qtTPeZFbDIuTDfzhrKSdAXRUJi9ptD+b5rEdrxK0k+
EjtdCff9Bf+y9p9YS3WS8xL/BMKySmO2dwlQFOZWEJyLFQd9LFUlDRvF6u48LXS6KsfbgYdX05Dr
kpU7j9XuvY1VoGGHeSl/8Kr+80LcH9yDLpQdpXzh67rK/FBbHL7wZLylVYwwAytQryiMdPNekq1R
NNcKYNle3UG7/Sl2HmhwPSExDKPSdQ5ro5hjlpNDWPF6PYN7DM/O+z0X60zoe+rfW/QfmB8W2+f+
h7yyHwjl77+LjBJlpmmPNGvElpSkj6oBc8wofZod6QFrsIJvOqZe9Y9lYkgYYgcnvlLQXzrTLTzM
ROMN3ql4//tqlkJn03U4MConNoPznD9WKQnaV4lu+MOm6JaUUZ14nk8WcH0+Gb1v3XcKPDGfGpSN
yovxINE31u8DTOSj+OBqlNuAdBbBKR5Y4waGqOwPDJN8CUOj8zSArHnL+slK21auzjdhCM42//T1
WyVbj85LB4Z8oK0mpJkKrTQMyuoO+k+uJ2bs0edzyCKQLq/aWvwNvF+GW4yrHE10VgeixhIuhkea
ddMFg3TpW54GlXjtm1zDtgJ4JgtkB2/0PWCF97J0QXUp+ZX2DWUHRMxhd6RhgczlWIr781zf/CHd
eGO5EgL2AnTaDny2DLjSP+GVcAXb7GauqdNEG0IgGys2+wzORzm0gg3X3GnF8HqHgIoeBiLJZkaz
dzNf7HzxVOii3F/SUcPBOQkbLZW3jC/WyQdJ+tK3c1HxXLKyFPrY1YShH26M8N1/r00Bl/1LY8Yz
knamlptoTMjo4cBvHKYCsgStsUdpAVrjcqpHV9kanFuWTReAjzkHKHozWpXnEcNG712Y9VOYK0Ut
hI8YRvyFIG8OJGltykFtjgeJkhf2vGBp7py+XLqamik2X6PVDXToCDBXzI1qLyLXFhQp8NDOSqYd
UOylOdekVGvXixGF/FnU4bUMHVodlcCskc5Hoj4QnYlFGiS74mLwTPz1DDUsVdMDm0cbrFyD2Gxy
O1GzPuW6U8vHGMY8Ww/ZPLIB4X9RguyjLWb3hgUWWgtJM2JL/pYJtIPgPhqqqVh6O6VTPqQNIsZL
CjhY8YGQUOPhbBOaGLKtYQztg6KyJl2vTckTFSVDFTZ9GxKaO0PglnFI6GCacqTlELz+0byNupiz
pxpq3K8rcmnOvv1xn+xt6rT+IsoZm5Gzonwa9BFDGfRcGNFrIDT2bRMM6lR3sH9iPyDdQXxwrHz6
lHgR3DoyT9+P8rQbGOnF6wnM8yeOByWympk0/6sanKpBH0V8VDDs/yT4R6q4pXIllK8yfSNHISOD
aUTh6UGWTo8Kdtjg8JGKON5NydZkx+WaNDmmnkCLoJ6jI3TIK4L5vQz6qvsilegHAIhbD6Oo3hMp
4my8LWdJWEfOc3KJfTF09QvTX2Yo9abaLFtef8YND6+CPujZX+CXnwf1nBhd+3WUKBmxOf0TtoiQ
Z8ukPJC+e8mRFRzdu/bHSmBUU29rIOczZjtP1LXnlghNUudF6iN3DPNNc85EIVNrByXwnCaJvoMB
b3BH27u1X9M8uRYxwpiwwCC5SI1F7ZSqTpZvP5xMkS0KDGOlYfT6qrGzMTpFFCCTpO9CidOjvodB
0oX3VI2tJd09vRNmv0YJR83oS+HRCYWPENrYO/yD4P70saWcJB7w6DhdokHJA+r0q2pP45eDRnQn
2Oln3I7Rp+bUilM+GNbaa7jl8l4MViQDLs7BjpwcTLuSuqeeeE0UaykI3LlODFXobeY+KpjSGgk/
/prnZuxIhfCntpg6uKmYsbRGuvKFZV42L2v96hY4tJU/2GhlHoNNhP61KhJNBPDeT1EAom77i/Rp
Dg70kbTCMu09dC7DVW/mKA+SDb2G2OEqOR+2PwMW8JASPssRBCw9eMvk3NFACTcWhv0+HiZP88TL
+J+2zafOEXkINCvRawrI6lMHFG2Z8sqGu0SrQn+wAS3zZxlWNXVvDJDFv/j1kp5Wo/5IvLSsGqYf
qYqjBDZjlwmkclgMSWYZLrgC5Qm5fbW3ukXJCwOnnM7/ut1fgAMck/EOew8/v5Tu27a9Y+XZSKQW
zSFYeJd/WPTuV40j9oFlJ6/Jv8SJuOA4dOgHQozk0TZNWIOsCWJmj/qTpgCnDEaxqtXbmze3VGPq
qyZGYlIF7vfuLsSXj3rDYXza8Qi6OS8VTTtOCyknDC+NGi076rXSnKQi3bP/Cz92D9trb0UXCm/C
/uz4zFSBZPUeNNyciMr1/4uSCjs/Zibc/mnMaKQ7wlNTVMSR06T5WF0/Oo3nej660EQvLDqJ5i9p
6NPLMkUkZUjnFcCD2DwVPMqffjVAk8cPRoX5pdqP9vkD0KOtw/Und6ouPlqDZRFbyk04VBJTx4dN
8ND8ApBj8CM09a6r1Z9ICEdZctW69T8/CEJkJ55yDgGeLlOwObyTGJv0jfsPmAnNzjyV6FULC5MF
EvmvWEmwvGIv+D85hLOvp/RqX4/Xoz+kWxAx8XrkmwbOqSeYou5SKYygW4gL2WA0yu0ZxZZl2jCt
rnE3FO/sLudwQ8tLgU4X8FvMjsWINMe/Xbg/UXVmEu46rFP5f+5eU2hnBKv5+E3CcEfIzhdE2wgd
k2dX0dyv8e58Yp6qn4EfdBLpO/zspxtyG7V7gfLYWNsWYzwCF8rNkQqOjijN9/UFCkN7442vvcKt
9JL28p889nBrkxjjOJD37miBqcnNf7WDJW+oY26xAe/3i1tYhxW/6N/stWbYBQhoT93Y4ryHvNAr
ACpVf+p8UcKhDMQSK1IXYrMDvUUDywBlF+B01NCCXzRybGa67pTIVubQt60Du4sKH8aDrKswEZLp
DpGuNB3Ce/ArvqyuiJNyBoYpgk8IOmetdNyN/EKGo0uM0Ta+NIeXGU2x6348HtLadF/RVK0TmDpe
/2/Z3wJiwZvL5U6rxn2zvqk3McfD7KvgJfE2WMUKxAXmw32grTDZk4DqbbVJUC3p9ZA/1A4xGqux
cUhzCD92PF3+i5JXVYGacK9ewa19l7Hw7LJS/xgtByGw4qKA9N/Hm7Fu72d3w3cpOYQqRN9Ls2N8
9qWeGjLOsSJ1n8w7yHcdfOdjTKlsjGITyXFCfBCc7Zdg6xPdEeblTSuGO75UWhKY3qAbUwo4i6gV
atQAIAmL8eVH378diISg6F+xT+hXq/wmHKDhOT2s8B/rHTN6eXDEDZ2hQw0JVmLdF0PFTy3La5gY
9HiGYE5jF55/IW4LZPJd3TMZWkzGbvQvqPWACttnAFlryzq4TGpNh2ePB88sYYnT7YX3hdcwiVq1
FPuLXhGZdho7O4ncPjYbzOn8ZS6BKHbTF0zz2xUxdmWQ3IbFZzM4JfFZgYJ/nQ0Hy+YQu+r5dvwV
tQIhVcmPiI5eGsPPLT+OsXiynvp8YcK/WQEi2LwA6Q/S+Ksm2fbK9/Az0oJdumwf5XSYyi1W/KZJ
C0W63Vn/6bDC8NIjLidYIC1qjKgtm8cAPkhD3Qw6KxmLmLWL/GjVaWlaOQ5nvpkJQGnNxP+t39sW
ldshP97VynlL4jvecTSiQVHp+Q7Lk605CrJM9zp+hOm6xskoj9ELd669SZROvrJnp1oMhMQS/2ao
b2XKcjI9Xva4WkoQVAX5Ud/U3HyoNY8i2R+1oeidIENF1YgIqRYx/p68hEvzSXNrptzolWf8vwme
oXeix2sOAcNVEDfFfRNN/qsAIVnEqPlE4JJH6cqFdKB4zCBG14VKunGjoZ8TTgOZZSoG4/OhHvd2
/+x84YrOdEalDQL+aWfiULNrVYMOq1ln/etQAOtW3k5VV3nQrJUIKZWI5bBkdUZq8sjeDaToi08m
v443YRA9UT2e80RStj+qGandHXPyBwHqlR4Vgk5fyTN3a1TOXHo1cn0BKMzS79WhrBMBrQhrXssr
q/x20fJQkGYYcB4Nz+ZdL8dKK7rLalNvD++/AvUlgXFsAUn73W1q9FxD8bFBAtmex3o7WvxqA9qy
HK0DojclTjVcCexhYN+U/CfcL0n4PcOiFVIT7TXUM3iY7ie/Vnwn9L8guANOvaYnq2577NQD+ERp
39MZZcLSmpbYVFWYJq6munZq3DUnBsgcI9uA1i9NfVy525gS8RIS1Caq7QOVmsVjj/e6dXH2pfG3
zY0O1Y0Z4AWLOU6gmAeVJbPfINzkOHfFsY/1HrJNFVAmqe6+EC6G7f/1OBbYSoBeRTNmaK9YC9tq
xIJk5U2NJkB1WdayoLucIkadFRsG6gs5fOxyu4jQ6vBXRNe/n/IGi5+LMD037wnl43sosbkLq+hm
8ycNnlTz3Jm7+2jdfncQqZD5F4CII4Q+8U/zt3FQGdKs9jCka/4S/3UNAL7ARMfb8gu2CAO2PYuU
auYL5HOzZ21jg7dxx5voNOnhR3NPjC7E3ykh44//kcI1sEMETtBxnLxhxt93ttEgHjj8tLbS4bV1
92SZiZ38dwFqEmyBUi3fPA1CZwmsSNPN4X9l/OCG2geOFulrCNziLrvEezqCXgRB+ww8jk34pnkB
ZqN/5JBcPOZ1EQ3H/5P2Jvv/hlFbm12VOqrzW+QYKATmh615JtjiZuW8IzBRmYFAY/wD4UI1zALz
O9K+M8CSnbR0QtFl1LcdKo29MQhHmWDNG9GAp2OdY3aj9b/mXMeDYtIDgArJRQtZZuEp8vl+aWvx
LeH44tiHsNjsgB9NsZqtLGEPiM1OcV7d60JfvnQMymZ5wdaobUo+qTFY3dclCRG5HbC0Tqz4kbEm
clYhOsT8QbqoRhsrabboMJDURGPh6kZTgs+YPT6Ivk6E3NrqxDLf/Ufnmqonm+B5K7Y52h8f/YdP
4RiHw3Nda89vX5Oof+jJnNuGBFKi2FqbIvMcJkduDSWxgKpKVmabKElW92bUjJww1G64P4dyM7/N
WUtnIsRBW3g+SG8rHYTVeZUpmMwUuaWpb/kKKlHooMS4whjE52dE11rKD7u8vhHGfXPKnA8Su3V2
3RjeHt/HFxFa47cIwbbgYyQ/CKyTteGpVgcq2sHudJMY++buoX5CkTaTCWBTj08aXYwXECtbe91W
Nd5rg4qRxc8w2HGnld8Hp5Lj2qxtrgvD2YvrxxpOBoR0gKNzwcEyi3t7KO1TYkcJqly84PdPnmNo
AxMuiP4T8GeveXMLsNUz4crx0dqAR9l9oIC1vgCWkDf4VHGrE9sBvVyVNLpbTWHcaK61D+/xhXxO
V5C5xm+xpGCkCmjYEtZE2RWsLGpKfYb5+SHZNJeoL1E3dv0hX2M64AaYSgRiWaNActFYKrflUd7l
PkzCtBtiSyR1LAl+/Ktgembp2MNLODHN8DuJLeVyP1qedwsf++ZJ4NyTqfGB7nvJM8gwDkD2Ac4+
oZtWP1qW82hxSe+hYklYAJYQ9eu890LIs3CRFjt3IVUpRtM65pHbkx/t06D8zT/fquUNQ3mum9Jj
/9Cu95kecCGv8AEe6KAKmMD0HeeV7KNqhbpUzkPF004/8L15kHw4qaBAIklsoJuCNcf7fJC3mYhf
iP2BLG54jKob7WhBIFoQrqlHv2gQ7E038M9nrXhBkFGdBSj5tpDTHuJgWS4wUU4dypKiJ6yNDFqW
YE6CQS+09ngZnCEUO9nY0QT4/0Px7MYPvlV1LXa4oNCr505ScEmw0vA6EFU66EbT5n3kIS7R7i5C
HdGFloSOlUb1EP7MFYGt1g0N7YSkqYqcQr3+9xpcMHkgpaqgRN+5P5z/y9hXF4sGhviXkkWBGEcG
FqzgY0PUOvvYWGi27z2EPYB+61NdcMzLoR163OkvEEioEgIi283cQFqOKqoNBt9yYr+f/Fqs0JYl
McTB8SmRP407SJb4YarGX3pfzDaSlsp6iruAVOWOLV8Ti0oqwLS90o8QtWLrF7ipBpnXI/2BK6oK
qxGd72o9AW5V1ISwJWrHHW/T8ZX7+X8NAzDpjfIm7QV36WA0yX0N9lOAQsqpQSjCnO7qEXfK0PVe
OiNZ1V5tkvC17M/sAAbpzBQE0iqHgZXNxv/9TvFl9oPePM2FMkDBdDsIiIDI/nlg1w4k/QOBCd1B
x3XDiWr0TUP7volpqCjGiE7F9Km/HHTBCUU7aCAqopubQ4StpxhCfc03onhDlo9zH1N7RcZmdwqs
DDJFFQ/SuoEGr9h4iYnJY3C7XBHOI/3Uhw/tOraJD7jhawlHgFWqnISPZFb7aj7HwaMIPB8aR85Q
DilN+mVNtVw7KL5mumirHsjoGQiAYAKKPZAlKNhboXIdboxO7TUX/rANfitZm1O8bLOfbfKRNxaO
trp2HNJ96BAnvUiCM2xA5imymZQzSvdFPCcrrE4zUL2QNmQH179IRT60GDMMnXRDPzYQyXzGyZg5
WAo5xEXbENTVoWYa1BU2KluoqkpJ6FmpeRmJ0GFX1U1xP1Z/xNwj+wAgysPvZtGfrVtuPet+lCHr
yRUxvDbZC+w2wlk16CyBCLegu5g8IyFH1JhPnMPF2v8GsulcrXH6JKUeoV6KV6E8yqX8FPw0TwuV
tx+VVwWP23ASZ1HfZcI+o06JtHAy4gNAjTxXycoLhu6YBkCoBqJtPJh9AcK0ajV3LFAHcdD2oXVJ
cIbPjUY4UKdYprjfr9QGELivLh8apwHMV2IDn7gJA3yYqzvvPexBL7W4OsX9vAbx+URfkzTfsc76
mVa6qLc/DltyhqICS9SnEzav4j+kn+GgFKymiweqoHqGVema7/olU+r4ps8J5eeN4OdN5bHwq/E2
dFnpjr79acGI4zcfSC1SkQYobUQWMtRTWzgVpRWq9I7JGx//V/xorAEOgJPFCHgW/vw3MjziH+Nx
A2cn9CkN+dmT812HNopFrRftVUuJYgy8FrM57lZREKibBJZsFAnMaQ1ok6UDJkvfXrGlYXLTVJQq
X45NDeQ26v7qoQvu/NSDwWYVb/ll1tTXBspuSiGW05oHNa/ODWYJbA7hjF7c3JxlDOV0+77Iq2LZ
kAIGTrHDlVL2ps1f1qPszEOczAgKPcYAFgn32Y+VKn33n3kq4nlwZP1dRMeKSG5lSgNhqXJNdWjZ
p9Pa/IeKzFdfBudgItiWeK0ASLNQ6gx6JlVvfep+80Qmho5TC7thWe2EnExlCyaYi3ePDKxvTavt
LwMS3ivXk5DSqZ6VsCuET2fbGCK0G8rLHApILXhCoe+lf9RoQv9tmzNwaXldxMLvtqrh001NRL/K
x98q/cRllbPaVRRmYURraPZaYcXxIIK2dWEWr5C0v/6cVqbDOZZfJ52oA6JrJoSSZpYEEyfyzy7q
MDzatz7ca4PvZ02XPnhRJc7FwSGgZKLYBqMByPLBXECWSUlVgOQvzIg5DRVXPEMZViz/fOR7Ynnr
WK3hd5PoiTJ73EQnGDcOkfBHgGmjExI0VE3HBTPh0R3nxV8AmawZdc57/Uv4yztWfTPcRUkWFemW
MFEYY5DHdMr+RZxQzN0bdChiRsEv/HzHymNLZIMU6HD75UgvuQdzF/eddzT6Vw688bjPtoW7AYIK
/RXnl3zFPfnwgI5U8mnjQEJ3sxbaVXOkywuXOJzLFV0/eRDZet0E3y7RWuyLYQFPX5dCDL14lzuz
/ZvWV4LSOSLiMV29C3Uk1uk9gAiTKdt8pQV8XLkZob/w71KPU6pUCVlQJrvDfIm6vg3wWX7FmuUW
TF1Rt+j4VUoNGQCwx359fd2AmYickoeEAR/yiMM6nZEB91NHbER7fxH8rRtACI71QEcG58I31zi4
iXanioLNNWTLIXpxDKJxQi4cF7PuwA/1mB0zsGUtIBxrKen3cNMUbkLyJjW06akkYmGhwr0QFVIA
dHQCy3Od5lZhk4Xn365yUcczf32xwoC2c9UVwHM+KT71rZa3YPRSHSWbRx2trUROENFQDjzEkD0B
ySKREf6ubqD+IEusQG4byUWi0jkM2dYsRckIH4wi33ljlkSjjzSJg7ltEcAxXOpzmU8/G2CK3x+N
vrIr4ac0tM99sjuGuMhs2uXrl5CA4qhBKklWjgxykkbNJv3DofkJDeLiAWXKYPPjx/Dy3t0I8lFb
TXcV3VHjbfLVxC3K8mrybt+L4Mb46+wrwPQOkLJ8LbzVL6QX6eQefQkm2wcjd/82Svw+jaJXzQlk
wrHPYr8vyew1R4dob3JGJNbLqtu7I7jjwQws354ysvDOtgy2/CCZZ3rCB7H/WQsxmmjQ3ngi4RY7
GKwDl0fmPRwzPI+EGZ3vI6zg8MU7cYksARPjuZUaZd1f8Px07KuvowgTMIALR5NzQ60Ri7qOC8YJ
zHatiW2l9llQSZQhZSkSNofCNaxlBer+rRuH4hWMwnDggrgvxgmmq2s66QwituL+MnLBMTtyodEH
Wv3sD4/HCDhiO2TN2aT1wE3RbOcMy/z+hiEbGMXN+R6+yzCetC1/eeDROHRSZ8cfTznMEuao/CJA
U2um9D9zJe5OrMAPvJe3Z5uxQan65KfWZctwtjQ8PxJJyRKG/ZLgXTxtpbo3786WVEBp1DjrG0e7
SKS6VJEZXYVLtqBxsDEwRisCeNhohYObArHGMfYt2NjY2Oe+fTXBAEvIJ3Wn9WL/n61KSsTujvrT
tIlxEdIycp0PgrVJmDSLwuaOLk7tbFFU0mUJOz0PqsQgISJw1VuXqnPwFG2Z6lrr0u3WKl5aL+WM
G3y4jkhlAnRJjh104rJcqQhFL+c+p2GRJ1xEXbgolCx6YmTXREoUPRgkNcD+VN860YMrgweX19Hb
t0VFsLRaJpiG4UxEn4mduqrVwojHTDLRdTrvssMtM8lrOdpX/1cW9ShI5yrbHUeRbgRK7ufpMK8v
8VpfwkjeqVVxzTmtimhxICTxOWuMfqt2uHCR3ExKw9KWgBDZDpILTZQMizU/0vyXyPVmEjE6rCpZ
biN/x0kLw12yFQJCI6dANowWea7MpUeUD81y5qKFc4GoDJfQ+EjapYlkS27VU4LlQ0Se/eh6M6Pa
yXCDMM8ZC+BSxZdpPcSdey+TgXj+d2dshHb6Rt20UQgUNTaECgn8gVnAZqVfqsNP79lX6gWaaCNi
+SIjJHPpBUm9uofZmg1aHn0IDyePLI5TLbvMCm4fAyvCHZjwwe3UUxq6KVAtEmYHBlySfPBymeQK
rVEAYU0TD+yj1+extYkcz1WvhlH8XVzWxBSE0zB8tSc1nDJGHCpPQ32Mlz4BWrptHTFP6zHE6Edf
5Ng2rH+M2b2v0dRa9ceVYzTiUlqBq1hqcOlJ02kybyTkoyPA2V+VcpOHXhZzUbChjIdZqGi0+a7T
V1RVg1NZF9vo8egTTXFcpplaqBq95fieMVjGVB0v+rWyp7kGSwLEsAxtvRBBMkFn8XEBdO8HkEs1
Au58jI5hAVisMTWJWykfw0wZu9GOAXxSI/srhktNaVWY5LfbNfxS0SIOzAouSgVI69ekm7h1bxHd
OyH7Z2sAE2DHy8HcVbasDhzvbWS0N6k8vimU5vT6jkOCtoMigIQk5bVQwHSU8g4IQXpeoh/U1Xbw
JLtGvm97vqKw2dJ74pif3u7JTAExJ+X3xtFmcLTIk7AyGBGGNDtcS8UJkbBGbc33UfFTKnK2ago4
FPBJhkd0dQywX6jApSknDIrrJaEdsp/mRqQm7G5+5wQcKy/V2RLax71uGAtbAW21fvoMGRgIOAL0
pAVpAXV6Ibr2AhLOxx1biH3x2nf7Hbz2rXWquqHIXvcSSN0wPwbTo6qlHPBGwaCWjIz4PUn0GDkk
03kPb5/Z1FzUYgWPeduZrCivwe9slkxf5lmc9vAL+ecd+yExPbcL3Via6+zsH6Enyw0zW5jCEWWr
y1sP4bFqFsvlzs9Z1V8Rj2zkIrz3tPVydU1Etd1fmBe62983ryNqI36MmF+25mRauaWoRJQXdD2L
aOkN2f6FH2b+QRsPzUGjZffhqEFWAsy/Av+jijdAvJXyZbEy6bJPIwgJJS7vQvxSO8DPrpu+jx6z
JDQpwlQ4zcrPMqiyhKnMKPehJUg65kugjsAauIRxz95aXrGRwaI8RnljcRAO+D6O+IKs2rqoTRkl
flJUNSAM5xaV7ow3qoKLzSkdO0pp181L9d7frooHyfOl6cLuF/oZxoO8uVvvRmfbTw/7zIHNRIwu
D4O1A/ly9RXX9sTlOE8ATz5PLvIZtTTKwtMwFy1XikBWqIVMoYxpLe6xPaZK8iOM8nhXvMXfk38q
Rsd/K2Yka8MJJDNckF4Oyp96jNIBVEfW4WMsmXYj82ehr6YLnl/8MkFqZ/6jOFtrnrJ8y4/T1U+w
NHTjeLpkGh6eOY6XzDHO/LyHMto9O5p7qLFVU6ea8m9FwMgHZP+3IzBKXEkwa59JmCqyyzpOqjTn
NjU4Mu/ErNAY27DiPP0QwuHw1uhN5RsYDElxvcmlYhtizb+3rag3SOhSnp7HUtbP4lTexdoBV9Ol
o0oDDV+qjg5PEdcUrz78Cv3gNSDTeBCFAMa7PpgqOJAg8ZBhUr/b1tSIgiGJLovA5TmGB+pV33BW
Sl2h4n+kksp/rImv2XLthHTHBsrXutCoC8jwSCUDr6xWDZxbx2nwacRYkqNVrffDwazUlIOUOn/B
0DEPrPjhuqybve6hejvOwmCZWyIwTnZOQvNypNH/qLDw3u1TD82F3YhB+gVZRsiULl1jofgVaPWF
5UMR6Wjr8M0cDAGqDH4IJ4zqbIyiz1nqQas+seWiXGdlks7Ls+ejGeaSlrTROXZONtZ5lNymyyNv
SmAAwOWiU/dOmaYWYDBCGGW0+nM/EfGAnuwQCPAae1quOF8rcuaIWnkPeJC8injPfndbuF4ZrHvn
qPrk/F/h2J929ljhJVuJGx265gTjDF6BgoMJouXsbci7qKlEaIoB6Iqxmx2fXTiJt5SbNC9KFRVg
vQ3qzQLU+Jp0lzv699gutkHjsERz23LeQM+82PXOLoQfBcJEbTwoLuux5GPZfBk/UXhyPoeCatDH
33qaYgdQbDvs6HJhEfKpGEu+faamKKabYCh6Sy/98+9USNqzC59AP2rz64EqBf5Q+1ZabFBbdZHQ
TGihtUnuHYkwBKFWW+C0W0RddhB247h1F7ycq0IlDeLyvwmw5hhkxZURTXqY0I9U7StQLLYYTYUa
HdHhdZhjogWhZTFvANi5W6U7hR0oQEbZyzZlqBDgV7iCUXMPnIdHDPq20/TpZUNwl/6tYUcf+2Th
X85zhhfhJMxGoNC7aWByrTXX0i4q1PR/dmSQ2E8uxWzdLGYhFArwpOTLN/fAONSYVMeJCUpoGSL8
CLWs/NEoqSopWzzK4s2hyU3c8iTjr/RGUJEngRJANkC5x1sxFA+0ZngzR155ESlVhk1PTrrgv8h8
eBdjWH8xA513/JtbNnnz8gJKeK105GrFgk4MGeGAZUlq+rRwhPx8AJKVYUgMk7tm5SNyPFemuGuX
DHLD+7I0+tbrAniHA5G9X7KRSXwgjhe33pXXJQlzbpwcxl3fss2VTxKBYKFb6dNJa4zjqYT/KkYU
eAO/lxL2op39bOPsPX0vIs+q9RHq4C2qv6P42Xiqfkogn+UBzjLxBSHowvmZomeY90TEHhDk7TcU
Is+4tOg0z1R9REdMi2f/29BvuEcsnhmA1ZfjfokSl8zoG9HWY0jpELtFIM/pWWxNuLk1oFztVzPF
Sm9MINVG8MUZhox6SvjoN8HeAo4wDAKClH1vWJKlu2vFxsNe9ysSNRS03A8ythB/S3jXEiSo50mG
yBk2RjE59S7UW9YreldUJheVUUa0hFNgfLp9qTh6ULeezUu2rg3UEknVo3GQcU/D/2pPtAod3JEn
t26siZLZIkV9FYw5SFAIo2aRUViuN0JSWiQzs8KXV7aqCSAwy9TroxkGL9muNAeBA/bP6D3bGATz
qZkf3/Jun8DoPu3WFprlLpFvfyvS/IZeHBUS17YhAz2nl+nogSMkCELCrzAQ+MqfCSh4ppDMNm5z
D5kksqNNbs0ypwELeBZIY67+13WamrlJjWrhhMREd2INgkYTzaKnvhKo61rZzfkFIQxTLGrUne/a
Gh/+y86Js87CKYarm5ARbqyyrKxqW9nD5C5/eWv2NHSxjKnm6jBAYicoCC11vTG+GHExXGr5q4+1
AJkv8sPyNBjS2Lnr94em5IpMBb4qGkaJOn1RoeLyT1SQ7FkfbXu7HXI//CjANLvgH632ZJUuwxSR
l4TkES9FyjuzJTmjwy1UAS21V8kH3pDIQLSJoRttU4zEYojcUSofaHN3T80iqOR7bB/GVsQAhQZ0
Cr/EQl6rF76x5nciO6rfLr+NwkYzY4z0nCpuEgxOqGLfk8T2pVE6F8Hy0TQuH9I5U9LuZbPoPZCI
fuXpj+kRG7gtHpaU80fUdTYJt6iOZn6XywrqQ40HZDoEiXcOJ292sW525wsdu0pGc2m2y9dmqMQk
OFphVhSbuumxa5sc+2PBwpmcE6zJzq6XM/DxvOwPylvrWTq/qLXeDoz3gGmEz7RteHHU8eseenRT
DijlwfgFg9ke5EMQZWN3IKxBBhzrcHgBulE9nJzkk5HKoE3tHEWg3JUSqAc8xY0vn3h2oPK+qIzC
F/ZZ3oXMx9gqIKEW+bOoRYtnSeMG3Zsifl/EDqmhz3uytN5dqkzESq8/6IbzULwt/EUg42kPNbgD
Z27IbV9B/6Nppsj7P4Qc/sMaJl8HACSwWeFzcFioReVvM5LFkGTzNS+DIAzrgEQlXpk/NwG8pcxQ
SWkomNOIwl/YEaqj6yIT6SX7uXpAFkAboyv2JYaizVHfv7PIMFvSri10O//QCqwubeIvUYmadSnT
RFR/VE10FsT2nXrXhY75PuviwdNtOHQaWOSKVGxgtlMSen0XLcsWczMbLJ3k8KyGz7VWFmNv3QrJ
ypRacK3gNGOILyIGyMnAS8PGtxqujH96ByQWDUxfPQz2h5P6EdJqCpXP5tAl4zpJdglnyaNC5W/N
WnFWwSaO9GVxzCjTBKBvemAiTlhzokpzxK3L6iHdAwcjxlsjY3uCFMkBqLo40iLRo5ufXS+etUHS
QCN2/a7O9o8L8jfrU6idK0puujO9XWwhDzOV4rNXz8Dlserr4/ITEsy/PxHUxq6Mpg9o57aaZQVj
7SJv9Ytr9s7GQaW0U+rYVSKJxKw20/2HxrK96eWh+OS+UxlnS1ScR+KMnGTyfgIjqUFF89QKdZpc
pSSw3di+hW8JqNOSXHDy/LElehQdWVhQUUaOrKjO5MsTH2HoRPz9obiyNKEywDyvs9v72E2w6tFp
mEk4pTjsYlnfjoqoMmpPZ2WwCMuNbEzbsvVg2FB0b4wT2FpY0p4n4ZTZMYu1q/JpNgvlPMX8ry+4
IkqREA6wmvOv+bmjOvz+LdedFp/O2T5sss9bhjVjTrIacX1jVhpMK9100hToVE4kMi3AFWO65iX3
UVMo7sBZlS/bx33uHUw4/tdIXBNHfy7YRPa+/mtLah2viEGOSdu9KN+rlHeNzS32+8GbEtkKqf3K
PenU/AzNjxuacjWvhp+SAdOYuCmxf7ENXQn8lCfPSxL9dPt6aCy1Mda5zN1XdPuZjIA54IQ82IuT
ew2ibS+A/CwTtlQFaIydBAF/WcFqSX+8xe2Ryt2tvI4nMYT5dOtIVe81yTFbDDmLFp+24h/6DLvy
KInMXmipcctA+B/9faDxCHujxQEBMtz9fjYOWhrUkXoK1yUBY6pbmTq9In2mbULoF/hq+///Mexh
24U1or6ovEF6DsCWg4dBI03dxQOmZAF0FivxXHMKGz5E2f5S079hXbSy9N4E8gt0vd8fJBksFYED
001rwoWysOQUmVwPwL+RxGelqnbfJuTmpSLIUjtDPYzZnXRy8cVRHtd9GF2y6CG3/JlWoUpMDXHF
tsnFoVqdoEM83sLOWcNoCpOq9ypEc8yHvo3N225PqvAB2v1tASzDcOgznZhMlEDKB34Y34KFO3gX
EelnWpMoxMTPwiXHfM8w2I4S/OtZrx1cJmajkTtFGmavp20rZV9fz10vpK3fk0vLoOjpFSECEKi1
0qszLuKp3hFzi5q4OviQFQ/062vRQ1dcvvbnLVQ840+DIWqau4LyY6GfpM4EIsfXszn57h+aLA1y
0nQpHIHSF/o+oPRU3GXa3CRu3F621ZtG5JW2abZmUpFUGt0bI1KQ6meXvIBCGwpb8mCnv67BCsPw
aN/JENf2OGk1o3WgQIeaNjnsWgovhbj/wrx7PE7nz5OVRSwswlZSth0i2z/J9i/9zOG3LAW9hNsW
tCLn9R393vaefMBbzPCJlGDuKnLRYqHrEsSCdAY+27GAYAovycnkAhDr2WzSVuYU1E7csveejQhI
np0O9fv4pHz4bEvAt9/YD2flqi0PbRPdKXepZ9WUG4/M8XnMngigIEKq+TTwhVv9wJ+zheZSdvfi
BF6GbSBwnzFuXPI16iv4g7w5fdM95IChVVHDTLsyBRu5mISSUr9fI7NTWoBn0LoxtWhyaxjZ91Ti
LFnTRft6yqFqxYhIfgymB7FiJ39eNjJY1AGTOnnO68rUOBekWQtZwYVksQM4q3YDyy90FwKycA9J
/+Ui39hERnBEE/o/NjouBoiTw9zff/Z7FPqw4m6BImUKDbg5NO43UhQM8eterrdld6RndQo7r7sd
JzkU1P75j7TFla1wVczPzDdJC+GBWngw5Em3TlH6sGFYgHB0NM5Vd1xj5OmlcbBVsqw9//xyylcM
wfY8hOk9bIWt3guASxGF3Zfk4NJRMybxo+uxZ8Mk+j6CQoOClHkbdoC4CzNOMfO5vhv0Lj6XY/3J
jqCP2mEqV00o8zj9yLFWgJ/cHu76WktNhLxIa7lBS8fXK2YOniPtVK3STVcuKg61Gmz0ftFmBwn4
hELdRGeLXmJAs/A/vgoUY0U2oa0V1JvpQqAAPapD4ZsLCKIlg04UuEK4YCbbk/iX1jCfHUKcKUOG
oV4z40ChCPv0m7UFCZgN1psjm0l1iY/Hk4ehou3dRjgLNIAQj3kOKOgNWpPdE6/iGwZX4fGfrhzh
H93H4YWDTRJkomGHu72TYN0V2QhYZBLm+174fLPRhid6KcKm83jVBvJeI910zRY1QnqL/8G/gme4
kh7gNqII1mN/4WQBHyy7QmGNj8/8gHOa+0Xkpoo4aHw0dr5U9V54uLoWC4WMT/A8pRHb1oCl72u0
xws+of3lWE7EH01T7e48w+IUc8uWTcilfVTtrp87656S1qLAD4vRPv8Xs+6kdwtAGNcIbqKyVmPi
8R2tGtkhyTtqYJOqoShBYfRA+fHA1ojo3R9jwFv/7zjQtA2Q0Jsj9S2ZUXQF/34bI/kp6j5ttQoq
kHUJ4yRP7ptifBfqiKo48rwLI6qaacXgLktnlpI2o/HyDSgPfURnn+XWWLcII8an13GG1ZZI7+1G
KvAS60wgq1C5UuKww+hu/8dch5m62yjUx3SjpfNIP8BTlhFQNNpBWkILBevSDGhrQXjtMPa6N1o8
bNcsJMSN52jq6NhZ8HqfDvETZenRcI/55PmvE4o01vRYhcHY7RFPJoU3kiaYUXwRCpbZa53lvvrx
ARbyWO8KmEPdM5sLfS/bXW2n4MfTAn+1AfKM/rSkKlfAj+TZR85SHGqki4/9QTNBnJpbDe/GM9mh
VSHgXzuGr7TFNmgBIbMMz4Z9f+vhGmSwGEhGvOMT5Wlp3Iqg+88bFffaynGM0BRcG7FtetxbQINH
c2TLRNGh6Ps0tLCNSNenXsX2ZBni+v3+3RG7Lw87AZuYF9WTtK+71PBsIcK5LNcwVZYGV27acezc
WUEeviUehG3pGwIZ6VV4DHSZNkM43XojgrJNkLB9Y6V8dog7VCCUxRIUvjXS8CYmPWraZ8QyF2IL
wGcGaaidKIOSOqCxFEHQ2ZzRpuO2Qrl08ovqRchIWxicnq8lKHByTBJGu1HgGtrAxdq/R/GXLkRM
6uwSvTiP6c8iH6PceF5ZgUCy6ftM10VRlinJ8SToGG3EkjzlI5mTExrSOrHj2pg56uzDrk6kO7F3
tIF7Pge6v+KHtDvJqWmqGPg+pBN7/wS/1ZulKSvvPVL98V31wVNezCDxkjQhuEtr4A71SU2aCQxk
BOYWkiBAzbuwQjBkLCpZxplT5QV4ToxY75DRNjFUXTDk7x5qb2W9uTIxzVRPFJwBHWtlRFzPbFsi
TUjduPczToXb4B5GbQOuxeAgJHPAlWzJ7J5AuHfSmlJ4Gfw6gKc2jnwMN46cnjkVubLAwa6fk9cU
5N4FCZwfX7dwQjUa8pUv2mzZq458mKMWvbh1WklCu28j934GwDOYqW+P1HQzd3XRrTPRig9uvnuy
2BrYCDxOcPudIJaRO64xPe0O9lUlaL+jr7hOE6zRTkZqF0K7UcMEanWG5827i5O3d8Tu1L2HIQML
s7ekaJ0Q4zhocLNtnPcVAuRtF2JnbN5O5naPvq2xdYdkTGzhh9zwkWJioUE2C7sg9Alm4wJQ/qPy
EPYcTHSIMZMP3v9T65CzdtHVbZdAnLzbf5plorSZEqvjy07UBbJu/MMWxaZKiUBDA7t4XchxISRz
K0lI+F/QBwveqIf0dibNb4S968u5PGZ+hXtkTr6qp/KVweyYGsX6nr4KaUy0qr3/c7GuQBtWP83n
j/CtvkWtC61+9gULDRZTsNkcQaVYxpk9hKCMevmNrA7dMoqzqNNhxyGRa5zg30pg3qPbG8s9UdtE
iiFQR8IuPeYcx6b9C5INPAYbrRjmUn73r2mMZY0WQcDcoQuTvoFN5g9HSptX+w7zMtokYWbms86L
WAmbdMBne4T5JlZodsw8Uz2SSjOX+ZP2UBsuPjri8vObFSU/WW99piReGDXnEkwWH0Jslp8FeVHW
NbxyI8CR0WJvTwMOzd4SO+hnY9EVwHJqFmdCuiVh7FzeWBN2HRtf4P2H4hVnUNz2K3t/Er/7iPyQ
vE1TE+UBJQkLkbsMkDHU0mh3Mi+urlNyWg/FBK7qJd/MoH5wQVRE3Ru+8kED6gX2YFX4uANOoQFy
wPnN+Bl87zF08ADX9/rO/KWuN73A+jxXTUMwGXvRAokVZmd/QtnTKmSt2zg7m+TpkLOjUCWRsllO
1ySMn40jhXGdjuEsWTncbinst1FTzLtty1qMWqoMSOlbfrFu1M6suGPVCg+shPPEDyL5bjgQ1dBa
M1ZV5BRk2DOs0F0yIEjfohLmItw5k+pzY38s4qpG1RYP6AWryauPp4NAUlrPnQXZoMdRXrN5ikuy
3r2MYAQfVPjcyVsoigtICkHBugKV5Sep4/nSJmHvV6WZk2gekSl51mpipuLaJMxZ2Y/G/MY0mPDG
eDbyiQes8EyOakadV1Mc0rB6fiypQ8Gw8nWYBoykufJVnu87kp6kwmgkqAKonj1dyDnwHnqI4d2S
VwxhQhGfKLOhKi0iy1sClHtUWBZt8j6u66OXpaewvLerLhx94xx5elqJ8Z0bbEpm/lE/7GS1whYu
pR9rXnSf2n8cy+uqClRd3veFugZeGoccWW498sQjbzBskUH1ZpfCyL4L3l9zOW14IdZ3iQ+HAiwn
IZQ8zXBRImPjOaub2EyR7C5B4o4f1OkezLTzQ2h+4kmXkg/BAx2tsZbt3gLyNDa+y9VmgB8U7b8+
/1xE0KxdPnRzov7OlphxIJIujFEfbTm8UDELguVXuC6ZjQ3FsP0TtZlfDCLmzSuubUc0RE+jPOGI
yHF8g43oso8kdKodmOqkN3YtKjDv/DWIQ38n2+nu9KdGFKUpI8Cmq4QYMP/kCRrLbqvXIEcktXTH
VDiMtCZr2HFuGa7FrnY5aVLZfU1Qc/ThOGJhSjosFHnJJzP/1HcPycHZAIKz5K42PqtnnHbegjOc
xnbNY/l/ZElKsUEmE6EvNcHJL8guOn70FUu4tZBt7ErbUIfxjLAfN+7cgVaAohp/LXLQAwHdiDeY
7sZLCcA9aT6ZX5DVQtJDCQzK7NO9WcEmXkH2TkJ6sUNQhk7C820zTGq0wQSp/6K8shjX0mL91/8i
/ggbYb83LIvxfK5zewlMZnbBnaALeOD6IYlg4UzURPlkTTCRaGSxMWLjPCsYKCFCac4g7sQX0hyF
ihnwIj+leWwqvQnUVMqGg/QWU00Yu5MzIbGZJ/inoXC9iNu8pWsu3IpPLsdx0W7dWIbgvGXvQPxR
Sm0qfULrCX2yMzpBLoIZMi1s9LGB3ic6OanxhkqRNQ8O+hyLonrTJM76vTYLQyiahhHzO1GW/9Fa
hZMOtkQU07TRFlekyOxI3bezuFDNb0Yez4Hix1uM2k0nXf4UTZ2Wtc1EruYYEPxUr/S2MWp/bD7Z
sYRpymjI1BDIyqc6usyZFPiWDc+V2fU1LcN+eZcVH3PLwqx2mOR82uKQDnf9nxLhpKkdYEF0zH4e
LEYLUVGOacYxhOy2AxUz7Azh+B/TzsQJU8mpA4LTEJ3JvlRKEm7TTGmT21fcsavTPsXYRFxxlimc
sJWnlJ3/EcKZsQw+Zb6/Z3TugsmNHrlHipkB3+hozE7yQb2hj/+t+BB2osL4cVemoGuIW0EukHsH
zOjX+p1HzqHM4rJOLpKgnxYHXhGx6Qq98n65NzXzcqnrSP90T1UMn9eynU9A8Csu9n+ofDyRyIdb
EVPQ4xtSxexSNVamIi+Gc/8lka6jIhcy14scxM5+aaNJDuAOzSwPxDPTWt0rZq97aK8w5UmkxMt1
2kJWG4Oy8+eg1vf/7ASaxEl8wPpeVmaPbFhNqnnhYVhvlsSF1LiS9+Ik/XRKXOBBjmQtcjzmqN/1
tU9ryTiHCcpO7nEwQv6iVhUdWmRMYIZWZmOAtGFmMhEtpiokdUYiW0zg59qM3/SHQxFTbaL4RbKj
1fyPpPy3v6XTK5ZjGHYR+AN0YdyOWUfeUTSiqFMIWFaYEI71HVM1/bdkkQ4tzp8r+F6u6yJGpkf2
hhYvD10sMKpi9NkiEDi8UmNyGVtbIhlCPX2aKHvGYbVP4ikZxLiw6fcnMRDH/ztpubXBukxVGiHd
DktJGrz7/a5j2am2CFq3SssSI7e6ZbBcJs23DjNueNSbj/ABzVPRv60+2IG2FCcTF4cBCUbn+6Ts
ZJoKQmpAwSKYzj5UTp9AlF5FI717/4tJAB/mmcer2/vUXju7ZHrsv1Ip1/WdBIPlZa1ygf8yieOB
LVr6fYn/sgQfmWClYwFpRlioLlmryrHLTlAYFsjUU7lZt1IvbO/lBFpOSUzHYZUxiAgiFUZcFQSW
ROgXKj/NQkSi99JEEdk8e0rxXqE007FTYr3KStOrGfZHlq0Ha6C4s+XXBpHaZ8gwtvpWg9TFR9B2
O5p0J9ZwRGQT2sdPPNH3oKWkmN0lrw6kaT1qsnMiqVNhneWOko6NqP3+S0yxv7LA5i3MSEN1nJgs
oOs2gco3T3waeJQeLOMJRHjh2EJzBYjQTGKgfMK0ZJrR6DYws2UFcm0EDYy6rsE/QFHBxPgUSSTv
o8dckwRENnCmhuL7gbJdHUn92sVEShKtDaRnLkVXEeGcWYf9bKcFH5OpYFOZkyQbwMIfydQ+IPgb
AgMoPhjC9ENRvK04j80qrzW0VmBq1sTq7q3DYl3txvmungCdcXtHuWpJ42/RuVe0ftmSxHjv+jdS
OFQnmCFVqGL0p5IA3ytUfYcukVtjYL4OJVyHFMHKCNvnCkPfFB8tJE9nFmXg2bBMJCrqyp/hBWUg
hkIe2B8BNId2TrfGfX3G7uVFfxzdCc5hvt1OzNb38vt3kFTIwWv5TVsIq6O65slkJX8vcHFeE51v
YAn2/zxDb4m0cohV+toQqAXq8qxgEZ4aVFvoXz56nEtws/d76G9fWbbcQRUouUTimalx8zRv8viX
bPpl8zxd3hcyTkZBNk7/rVvkKVQhfJUfrzTC1BXHwrah0vKEep+3RXSxPgZ5cJgY6wUv58+zK9jT
g0xrykU3QYScjA44A1uXdalrNjV28av9IaMjjzXgKVCZm7wI3391ax/aAOi3UA79uDPlLYl8fnK2
XxaDOUnaT5xVk6n93CgaRSx7bLDF2kSCe0p5uTIptRtq78rm5jikKOxqnMv7bVxzg+WLXyiTcoAm
/dW86x6kI2xQptySk1HEiDtBZVZNO3KtkCxa6Ve9tDJjq8ErBpUMYjAajXfoplhONuZjS1xrfihZ
wZ6azwCYdLqENDV8N1t/rVArJikhB6TMEKvXrAgTcqRmvhOBz8D4QVx09lvLdetVjBAAPiuNv1X9
hRCexU3n2W2CMcQi5Zn3LTbR5gcpSaCFrdcvNWprrGGKqlUs6l0NlG6fhInE3ANj8kttWSXWHiNL
IDwxTyEgGsbNNj52jSQRtHAtRufWxN82gCbqXDK7IatWawhr4jVe8sfZEF45n297FBSaakmu7x/A
9q9+Mf8948anytDJpf80jyEklZLCaV0aE33oYp0v2BkpMhJxFazqHa5VPQX8FRtUudX0NvTvucfI
01qz5VJDd+RdrHMhyersrqD9IpRnFM7ntDd9NTKcsIwJJg6UOwBFJIlC6pCYBPvbOOgDDqB+KMP0
+DHZJs7kzA8vbS3iFCCViRYHrQTHrrTVAANAMlNoA5yN68jGNv1yerpSGzBO34nD27KdaD4NWaaB
rebvU5+nzmr6kQ7P8oKSyIZO50DAspxdFargI2hmsyrkNmO0cUwsESFi91P8j0DG4MOaIP4R/9ao
gV87AAfzRLwnBI/YVAbB5iLviIO/5bcPZLOjUmq/+s/JXrUA0qdC4fgeC6A/HtnbqDjs3cS3IzqL
lyFvJ74AILUgzp1OEqCjAPbzHJPy0I7qjyyaPL5gR3i0qTDu2TWbEmcMKy4esduPMfWZWkPrwRPV
kCxFQJy1H/SpGyvpmQd5XxZfnl5zKOwJNQI/eHyVONgrXr2JLfV5nRCk7AQa3iDc33dg6RlgQpAm
7ar1mH9MFfZqrAZELKJsLMk2aUvJxFDgZTzthtuJM5znt8xJlcXyYA9nzB5PLIVZhy4gdrM5ANrR
bJ51TAEqFUTY1MheYzA9LJXqtq/WYHs77M8gdwJf+Kn5NjS6Aj9gHXpihjxWQ57d1wtyje0pseSV
i0srq2MHvkvDwe65ZWifY8rvRAg1VWgxgy+St7xi2w9ft25aRDGrD+jI0kmNH2EcpRV93GWBblyD
wvztB7bzkbcibdGeue248AJaZqRPe4RlRP+rhi0cvuN2I3RZl7aRwN7kxatXaC9DJUPzsXNmeTjT
JVJh5oNXFtpNidX2qyyN7ezw/9uA7BYC+q/I6IDU4m0NWlXZvr9XDJtg7l8GqsxqfdCOKaKYoRFY
1L48YjF/7RMSoRSc4pz7pewSlC+SyK1nQITD0zbVLFzgnp4RTfGtS7rHprlu+iLQLIiF6NieQWn/
fUdBODWnE2XOdNeuVfyyQ0tGMPIfMa+5PQmI02f4AK/QOIOT+huUimxxNiDa4J8MiyMkWJ5/7hG3
JZ6FY8yI5i9QmUio8u6KN5culnBe1qRh+DncT4pnauyuccfCUUZNndWoT0681xGN0Xl1tGOr1qAs
dYq6Yh3itGORqg8RJwt9YHNPcNqEBUOSdpnkbHFzbZg3FNv4XbA7xG7MNQ8y9CPOFEIRD9ROeGpy
cH8juWHgeTJfj+Z/uIxnH/j9Vca++Mz313dZinSaHamSLF5+XqVxVTdJomsaAtkqIlnP1auFvBRh
Y6I7GqVyy6FAHtyquItXSpmfBzN3k6AHXamL2BKQzL2chH9G1dC7X+BBNCFfEAZ+29tkWrDbukGa
uLDG3J+lOIOsClmchMPXZKeUQjA9ht7prkibEA3wBl9FUQPayd54+QFPZVkb7kAcXR6I3CKKPdL9
EsPo6PGDL/UzobFCulJhBAuZj6syzqGQ5d94WkF/aOc+igs7VCVUVLHQpSzlRd0ysL254UT4gB0W
RPMchjzwvboLTXJTY57Cx+K+S/+MnRu0jdVH2NOHLH9J++AhQchH/TF4OuamKZL39/m1WZwfxk2j
qt9YXkNz41m/I4OOSwbef7ty2/4BV9HaJDeUM/on9FzCYrNeaeJ5XPenB0qKX8mwwRPBcwNeUPkY
acX6K8EHRKNkeiz6cxMU8zqMI8tVnvtT9jNuiHpEj/OdDrilYCAHL9k9ryO6UMTDlpbXHuSIvPPu
LY2NroGUg7ugwYgC53n+vkDkvpqxxoVWimjyM/Y8GkWit4bUIh2OORQN9gVvOytcODlPzFX3mDYT
aWq3suiv/kQrfYciRdgGzp56Drv0ISgw94VdZLmXBv4rDMVJQRQlSWK8XM1tXsT2Q6lBnlwtn40z
WIM2KaI22jSdclDu7CfFRmFOOqEp0kV7wTlQxIW0/4B9AT5Jwx934VSJ1NjFFLx+UkZdqH+Ks6aE
MslPtFCiYMLyBMaPtYYIl6XZ4Nv8zHUJ36SkGdkNZYf39OAOlI8kTB6+F7OenXVAPN5utN6J0uGV
3q0i0AetgqedIMVUsMSCWrb3T8S2Ea6UKbDQj1t5E2yDBrHZE4/CNgm6QgvTATuepqzTiKNCqvLo
UDu5X9kOVC41L71KjuR6Yf8wQ8pbmpfsvRHLPRTtkhwV7FU8XxHZauO8II0F/J1nGgPQEAq732oL
Y5ZFSjjeur1evA9xoy9By9fNwfvj4RrRRHL8YM4AssRTSUzh/8YJpeBqWY8DzHosYi79A66xseeL
sjGT68v95kBDmlff9AtanoEGFFjSw9JJugLwKDW2w/4EwYIOXzdhltyn6gPUUkI2OC4EsQkO/x0I
n+Wg6sQFfAd3t7KgMFm+9hs3SESVDiAFhiGYNp60DDrM0Wd0fK+s6IMuwDPnH0vQRVddJVZr1v23
w+SR/IDmo3RouLxMoL22MyxN3H30vt5Tp+3C6cxg2DHZzn/RHV+Fd1et6k+CO7t9AMpMaI5P07Bj
X2LRP/z+3f2KgX9G+v1o0gGeZKovpU3gJ2eRktZjm25k84eQmqJvcj1h8rs9K5Nd4siCC1YOzeib
iXknJ8HT4UiuBzw0/rOTfM3bCdbCSKmFG1KqjMdnCdf5yO1Ve//aQoKf1kj5Wt3WdfNEtS1rlcT1
BwhVmXQjmhFCJ+p1stJwa1lcEJ5Omawj7iIoNxzhtKrZDlY1UNR46IzyhQpt0AOhKU8DS3Yzi8Wi
mD+pNtghWi7Aq/sXy8PIZPjcz7KHWw+wokV6VLmZG87sQg6JxKHwR/pb5I5rlNGDhs6icf514dsl
CMUDJibVO54vg5zcgk+f4vmvz1tet2JPUb0t2DK7Anj290N/EgYz/eh6H4wBYm75JfjzEq0jgrvG
buz3c3Y7KJZpnaslXrW+SoktoM4eYIq8b4qnkBRnIYvfAbMvy2euTOCUspiGrzG4ggJ6rx+4z1xT
PyMC+7ibyOyFjEpx5UZM7vMbEscNhY0SkPF6PPOClb7iif3VBEwd1jHOIyZHZJTD0ga+20+i4vu7
9+obTTD5fPiTHKLBKkae+Uqk/NPVnZ8zaG74zCCw4is1YVxk5/9auuWZVrguWUFqfhixDmS75UW2
45HOlVnNL5NvOKckKd5z3JSqqwVlFAF3Pf7IP9eJSuPfcWMnUnHUEdgORzTQIwWhILbclJdrxZ/k
L6xWziqWsOg2PvPGm0AbYw+nYtHkDKb6o6+tSQ0HhB/suCVYVLbbydwv1ivLyTecMNB37cwrkRec
oG9FNmtyat+kvJS3F/FyD85Qd83ELdEgS3RAh5QrJ9KRyZTJAQ4id3YbtkMBWPGzlhFRmQJVoISV
5AG16yB/M+RbJqRVKNzlbqPo22LVkdUnooNXvI9gtOAenm+6bUQ23E5th9Gmh5rtBUgxs+AWFVi3
HpURm/63ky/3J0hGTeDySzwiwDB+bHNiNQFmz1A0lEYiq5dwkTcXNNHPn8OOjR44fNe8iL/aQhlg
rgQCihA3xEhHmE9xn6RNMp4RzpVDqoN7ikF8CSYzzOFT7DUGnf9LIr274Pqrzm8BkC5HAzh0i0At
rWWLfjv7s5lrzKCW07oMUQoqJrO3Z8Zpq2Gj7sGR+7+j9QD94u7jiKK8q7+yvRTzBmUrhic83hQO
O6fyRvnUjUsOY6TRpkPRgTjgI4Y56Gygo56Npo9YMI+hQxuMxT5QhY2NA+XsWL9HxKQrcrjKMj1p
jGfx5lm99e1ClRH/Rk464J9HNfA7T/mKRxu9agqXRZ6d7FuOT/4L73qCqVEScWtjo8P+sz15QadH
Akj7JRHTC6Rd9TBPbSnMLW3rx1bflFgp3TX9FALImGUR8rxr624ZLdOnNZMmRcH7ouTZlPjlzHjI
6ymMTvEqX9CqIH20p0Df5tChS4cv4VecmnAYs72dYDdUj85OoIxUFnOyW1JXWtfd/CtSMe5mDIe6
LdxVAgzR+7wDxSRYXChLJHd1T0Spl806PemTpajqDGdvma4FgXVxN5Zj1VVF1itGV25CAd+Aq/1u
PVOnVfNJkKB/8JXTo04arMWVVfVLzgSB9OaivHZ7UFYUJvvZn+QpDPLn2UrjNp7BpZsn2iNXd3oM
6hT1ErsFXRGqslRBfnjBZQ2TVnAneJgFK9AsJncPm9r1DeKjAnpW57GdyG/Q1P3yqztGo9LiR60U
lhaUnjQgUlHM5S8HcU+oP85ybrkevX9V9wMQb18ry5WaG8K6s1471rUKjGvD5LXI30qE+bKKxCg2
g7KjLzwZ1d3qane2sO0zmNJEtKuMTmdZI7e0nd5IVtgf7KxH+S2REgDNJYmco+X4Mqf1u7WO31yh
4l+Y3RvE0rGsjygCnkI1nzKM6LbziQ9234YI0GPX7dArZ2eJaZnErqvsHGKdt11BMsSJuC6Bih7r
sWSI815LYkO+v2Jz33ArsEaqgQlz+b6tC4HKeE9HpisdIaH0gOT3txzEWcl9Oz4sPsakhq24x3t2
UIMgIY0Y/xTw557WTER9L9bzkorGTPLbWUqk8p1+EvlwjC2F+1K7JRfBj4zvsznAV2m51LL+3ZhT
bg7EHPPe2Te+EEgSI9iOXE5r0gptyF7FAJt0o5zOP3iSOUVMtO8QbM9/rDXb9CD4L7TtWA+vmC2E
Z5lEvT8dIx/djE+zvrGPAQoXNPyfNH1o+OgBqRBrJj0/ibxuoSk8XEYoLe/M8HDdTPZvCZDDeazY
D9Lzpptr6tyZLx/ZtbOCWXHHjxPgWgQos/ajcN2rwJykkM7WpB3CfeCreuApy2Op4OAXVOhIPp0B
RhqmeVAE1QwPCshe3/xuc9+tck3Awv/SoA5ytlgvc4Zyi+EesnJk0eAit2RObGjj6ADIqwd14u19
SiK5xhVDL3UWxrB82uXSFOp01YROLKP40MMlnzi+gb9dyYmcUPYiLorIsspJ7oHX1I3TbnU9AI8j
y1sK2hqVZ8RLEeONszTjeUJgXYMcvynC694eYmo03vjAbRswK39BYNStITntFyGt2n8x7Clm+efa
1XnK+KmvTjzXe2Jj/MPJQ6C8HY/s6M/134AM7wrWlTWHV22ongcClJT/J+iY+vY87b7b4WgIX9Bx
w1qweFxPgzcWx3syTp8+Jq18pxl6LGj0SL9ePtpvNlic0xFqMk5S06KTeoSsD+4th9sfEdOOwuxj
rOjK5IkysE9IdBJ/lpf9fC15PqlIY/h9wH3eqfD7mIp2A4xPedDOdQ99iuZzIl5ziG5UYDY6fZfF
TGLDObH9Yp+HWdN0ZM55HkZggZ6G/Oz69yexw5Alh0+x0IBs0qzRE0MDPKWr2dxU7zzkffKUlvTv
qaNV9xrjfC6VU8f0G33n41OHCeV/Vq9V2RcLfmHOM+7uj/0pV/DMUSrod470E+N2wyZ6b+9vpXMc
jTyHa9SdWUGaf/V2z9buaZORb7Lkiv1UlYX3kOuEwOCibSVkIx24CbQ4LzHPV+aVQVMOKULUC4YH
tV6/c+R5U41Kn3vTkZW+JQNGHGdKy4x+mxOI2YiqIYa3diwBCceycng3pSAEYwgI5WpXuBvKvbCy
ZZEZUVBkbK41M6Mmg7MTpiJrQtH2UA2T05qDhTfO63m706WILIBUcmymaeUwp7J8jsvW3DR9w7Rf
x/zxOpRvNbty0A5d4DzR+kbjIS89IB4A3viSzFbY5hkl0+FgyLbMIasmnOZ69iTBZ2/vAqWoU6Oc
FxB+QnTpwDnkf3vFYTdgRnhXTkTYw54CrZQjmwSyA+2UBdAS9uAFV9/0k1EmcdiV8JsgwPJOxXjS
DIteZpIG78PWGlnpYKzT1/vNc33dZeGJlVr2uy0mua2OIUnIgnCmC8TUB1EXbo8DSKw+giHioHDa
oCqiXPx+kYGvJgv7WwAdUrsCNOfQqHkwPEFV4D30RwTOQ6zPw+clSuDM80KflzBLSLr2UG4O7Otc
FQ1KTUtAitYydcUNwRLZMIBpvNeAoVeiRyoqbpkqNGo/JS18PEVXxUyESctDC7EgL1dvrlT7dwIP
Y6Ci+S81LQ8paVCGzHm0fMmPjVdU8+wURXQ3n5Ddcg3m0Xy2+PRBJhOEsvopQIohAnzIIJZBtRBC
2dEJYouKa5zTJ+O5ECTET1LgSgXgb9lGmiR60K64x9R9yxD/QMMh+JPSYXwcFSbuXNrdB5CAViXk
0FiL6uzPHFlRWVFPenpdtBFzj+97SF4wrev5D4LYxmgHBZCQ5qUV77NwjmUkRCdhJG2++4jnm5l0
aqRoem6g4D6U7o1h3bcyTuHvlBc/n5t0OaUepE9Da41teq+h4GrpiHaA7QEJaeh9njnwRsoIJGBo
g3tS2an0UsR2cCuKfA3fhqrRPi9XIcjroQMZN+XnXNUp9Mf5sG+lJ1jitsjI8ZgnU0/wpaZtez8n
6zP2n5HLsZ1+mpP/HSji13QdBAljBnjeuJ6NKpXUj0vme4oKuhr6Kuv8zneuNydP07X7MQF42KGa
bGagcSsvSIwuBJbir04qMbmFfGAWkZ/wy7buirCKCDkVbo+CT7h2nIPrwNttTrWP9xZ3NKDc/v5T
nJxt/eQd/vMMD5Dba3tKUz6ZaZ5H9bYOcqSgPPxZ2JbuXEvRO51e1uY39kr+LIMNSh4JKFgvBUAa
239Rioq4rvsyCP18kw48GipXAWN4/PfSi1SfiS8lP1D4bB++bJgZgDzsQ9SzA4gvPISC2kjCjkCi
FlY8hLIlLYvFtXDdhJXoKigA6qTLjrrysUroQfQM9I2JQlLvjOYi9rMWAzAnkL4cTvNUC+ocNzxe
78LtkNUpHhermwsVfGfh1TNwbZ7djf4wNtFm6ktEU8ylLkb/j56LF+oA8AT9BVEoy/Bng1ylBU3u
S8WZyWbrKa7xxq/Iawh5DZiAyv2HiLMKzjzOgpZy6UmGcG8xI4aAEP9SunSLkeiAu3avNSFw6O+F
QdzflLtXcO6p2Wem+gR0mqaOEFa7GL5nEFiJ6SGEvwdHx2DIckjt3TJOFSYqXb7mvG6NIqc2kGsW
+qGOuPrLXGrYRVA7zrrhciUOqgpJMlUAWNxnnfbAksp7ZcMKzjT3LrMBo2FDr1dX6anrLUowtPAX
CEuyosgBit38SYCtyd+QrdSqEcMyUjcUE7yQpwVDAJ4l5jOI/CL/4hijQSXOgEKwYXv38fiBu6MM
HrqRwLofJZRJyFfUV7rBtYfG2su49nkFWbw3lURBw+zBM5tawjZYdfi3A50ZHiwz0Rwf8QPmnT/S
PW8vsQj9v/URSPXWQKybvz9YU8dOyPJbehyb4+NSoMMlDina8m+qvv7Sne/1Nb6fda4own4fXYEM
yzlXiSXpDJkmXcdNLoaXHsPHOhOMTgeIz6xN8Iy+zLozMwdhgLElJayPcn9XhwpSQHW/UZP7CoUs
zsPM7mT6IxSBvKDrxd5TW0bt6Ez9tlQy5GrjXzGcr/d4raRLfQfx/CrcJsLUJoAGSacmyQlUdiJV
eheeSNWFwjlC9bvRZupNLWGT+GNh+FvL6OPfFge0SSx+sPAy6nbHS03EShm9AgDDggGeuP9IrC4M
wsJH+8u4QeW7OJII9D2ThmqUl9NNlRqA6fbUx6+CwxdLmyvlF7nKdxNHBwmaWFfPQF5xd9Bl9YML
TmnyZnzyXbsgMtNeki2wh5gud/KuBx8ohZopF3G8s+iRraf1MNxa6eErSWuddIK5Ocb/rFY13SOu
qEEBZbP5H1yRjx587fLSf+20nqRTm8qBhZvfNUVGOh8l9Q1LnuXHw0F6eRX2QKJWDd9GElFbqi16
0fnab1/PG0k2lUBHXotn20Uqi8jouarihrHPPp0CNu5aSpvt+PUWhVFyk9wAJ+/DSGlGhLBM2mYK
vFmOPxiuhkQf/4OHABSq1e8eDcrl7VXV5eQDVP1E7r88ErMW6rCHo1ZIIO9vtwXEqaFLAw7XAKtV
JqwPch6A0R8NXseT1duJAAWafIWD6/UPeBQqLzEAVXeI/PSkqFcPlbp1MIlb60uVpFr6RActJgLH
1gxTPC/uwRDiuK31tw4/LsQMmpPICrxlGFe3lOsb7+3BGPoXYBNsaQ86E7Rm48gU7jutsxdprDWK
/EBlSTnoRRJDUXvdgZ509+Zp1VaSsn48dW0facdEXmM2dI/AHrvBYW+8eOmSPT8mPxvpjceL1S1b
WNiywhYGWKov0LhZMRdvnkShkCHEM1Ia8OACjc/Yk9ddJt1JV8kObRUtGiWJB1nx8keJABHcDAx+
ssnQ6CVax8rklKprVcRl1Kq8yrQr5YmzhxK1K6bpXXgcBI1i7hBfmL3WUwPR8AvlQ2FGw2Bm8ggV
lmHmPs/SqcTU+tg0hbPjqCRnc18iRrZhiDnKafm/O1TX8jAag9kD2dm8bYYqxdNf0fu2sb6NcIQj
VuaKrsFjcG8D9wlbrImNFxyzOVIl+GWse9Pph0/3b3xlu8lN8RghNXnhCxD2ikSv4GXd5lJMhUBi
06JzKG0jgDtF6SM8Pe9klVhVAhJj5yQ3JaKdrPJwPn9vI7DrSguCuQ8d+SSSQBNgkGKQbZSQmiQZ
mJzLWkBH/PjCmiPDDQCnHpXivaFgMFMSV+cIooo9LVIoYvd3tSmoBs1vPh8sA27SkJvyDLjiw2PZ
BeMBzIfHN7D04Ve8DmnzBokgelQZhm8f224xs+rJbYXWtKAN5OaFdOIxBoxap5R48BED+bb9lxQq
q2Mtj9HGVyhXzR1rNhZIhPbZUwa+EUhDcgwYpc7ti3g7X2wDFNxxexDYrmPPKq4Dq8i5T6hcsAvo
+JsYkGMeHZgOkEwsTDl8HjWmS/j7cJxEo6nDnSPqGnXXmpjfsErN4M+3D6oFjfGHcwVQ3svG9YiF
XMP3ldbUxJXLxQfm3EwiTKZGkZz1kb+JXA9WcyxBqzTQM7o4EJB4p8YFTmvKz+s2iwAKQGmzJmYZ
k1EyYXebRio19PqJTb/R+bRZGWgO3OQx943uzYYZnJLVp9LVsriNsNbK0WPM8LI2AFEuD51SnzEf
hQhEqkPV0czpRhhnB0juVlxJ6vPycGfdWe1cxhiB+9U8ljzOaEa8YnhWkn5A0elLovLl7Syb6yPX
qgTqIkW8DVwQlsp04QhI6IAYiMyXFw77jkyFgefXOHWug7032U6rqyMFpiUXHlc+Lizj2aaekEGH
7W9WLHJN/Kix9Kbdudoy3Tg9qVCfuBhKJIb+XjN/MwCG1fV8wGJi6xatrtYI11oS1qA072bgjEw1
+fNK+WfqKdZAPaCC+s1fyRGDUyh+MBE0BoZp/IVdim5TWzn6pEVINa//lfGIgZPE8+QamQdQbJNv
HwY2U3hKurbApd5VTp8DONU5DwO42XABeNrnH2Zyul5XeP4P2qULfKJkeUQB93L1tylVjySUVuVB
IfnfTwsgL/vKnCv5PW3qf07S8YJY64W9Ov1z4+tkyDqbpix3DZzxEFHN0OFc3ACATfMoDiVnCj9Q
wQs5mNBXk7iMdk87Q/ng+L1LOFiJeJh5II7w0TR644N/GtDZ8a+F6pq8zO/doqAKkojwZVzSrn4k
VzmK1uUjCL9n/DTNu54LE+mca9BXRoj0WUWWlwYak98nIhqly4uSRzaRBF3+vSfCcnNArFU4xBCh
+G7BhE+yG5cq5QMNE/cJp7FnEzKWue5kloIqfxel8quyHGNCCfoRDqTvxYYtY6+TN2Gf0oT0vSwb
pKdwXWAlpJ+mNWM2p+cU84T64dhj6+gsDozwMxTnD/lY4HJ4T+/PHygTjKZVLPYokaxax5MESnYc
tDibX77Y5SdrdNxVLHwbHF3OXWNbkPQs/8EHfZNM6/xbclCnEz6cYFx8Vj6Hhfg4XV7sAw+h2Eoe
31oVzX6L43Swk8jzNQQ3lNc8r2H/zqH506rr/vM5A/Y3jI1+x8vlbHVZTlmvvdHUZ9mXzKWhPeVL
aVtO9un2BItYKDB7Df96ZG5S3hWycdOZ/F0wt0v3nmvM/J9XLBw+HpBvjSncDlQitkdt4BlWd6vq
5ki2NDW8JB3vitasJ40TsI8J0Qkfod83hc+33vb9jYjXD4GU6QMFiphmpWnkR0GjkubydsveeS9O
iSywwR7eknIaQFjywPz/FKgysMd6ly4v3ODe7a0U5+boTnj4d9qrRVE2hxUQ2OBe/uYfUdvoV0Dm
7eA3X6Ot2na+4QiM8v0h84qmKWfWOYTKiCXjqSUJc88gsrYnrgn6VYoJXtxQ8/ySPowqAS/HJGae
j9tiVx4svTjrxS6UhVecudpWsnfqIxwYh0eDQl4f1FYMkoyM2CCiVh03SWmNLRF/e5xlA4LHUsFJ
dmeV+XMQiLW1OwPItOMFZSKpNQZcdeqliktbtkxXDD/mH62DE/FTgYQ0292ncplTOcSUaljcR/oi
Ogtzb3v3hsLpMhCcwe/d/AwanCdYtZHX5YUwqdOSvBD/9wD2Uguh8pnl6ZqAZXxnIyYnS/YwacXL
LLZEIP6uk2IL1POR825OKN9ugDo7uEbJH+WhxejNgkPy2G8jrIBFLcxX2DUx6AlbHlr5/d22pCYL
uVfakrRKOHPxsIcKkwSCuQiR8OSqpaEBc4ulJOW5zxrk6zkoSQ9vT+HOt4ZjReTeRFS6UsGaCqG4
xOcTTiXLX5F0joT2rru7l4xYN2W0hIBHWJHKZ07jUoitzMsHvP8DU/wouywTBUXP1F2nDy2+HZdF
FBsSQqQ61RCXoikGOOYm2BS0vOMKry7/c4ZqYauG4oA/oIIjb7sNh6VJhfIMaTv6R6+vXNyXI4Fj
iBU7p4l9lEyA8g9KT7DExaMwFhW4QQSet2BF35jF0/dKip9coA7SLWXy6KbTvu1tPj3dzylFUVUH
RglP0vJjRhr3RaYtboDeQ4KP4M8v9EaYG3qiWZJd1d+xWNmBKzsbCxgiA84DlLRnu11wrzAf4Svy
G/hxZ/KQxYzE91YPd+wDK7EtDDY/eSavUsUWP+VFYZtXHBmqWtNVAy5nuY9xaAtxq4iksHCm3gio
NLnDpYcpkV44RJvvlto3LnUjjpR4y7mAGr48Z7rlgEpTFAJNeQhHByBTjGcjJGoXYeGP57kx2HUH
Vn4lKlQ6xY0sHqnSz+STLuWBahX0wG1pr2qz9eB2eXkdr6mtmMvWOKMQMaeI1M8pvJ4UmUux/C1a
CQX+WoKdOKznaqXf7WqtLU1J7TtyAx7ZUGUZgPX0FcX6OBLTxXJfF9Q+gy6Q4eBnJjdHsURCHQoX
ZWTQLgiNtr6xOYl4ZL+zrd18diVCwWPuJgJZgf0B75dD6eQvETawbmkn7XuZ4J8bNReZC/HjW8Ky
lPyakqtLP9hg5lzOH0Oi+++oWSTzBPe1QAfDte9k1wNBhT8dH5mxTCJ8aAf+3MEHEr47rumyVMIX
vkYXbhGTgDI7RxQnEIdHW7OTurEOdPq7D43Gn297tTm8+MuRXjmGKYOqc0dZyc2t9Eu4qM5C7faF
6/M2l9AeaM9VTba+SvsohK8DvoNjX4nrzWT0D8N7EvUccjGE/da9aporbCGF8Ozw5t+j8889YTNV
qqEjRI/5aZ0220BaQukbt5bVfNAX2KLpl1mHbjLB+/qcVqggPyHscvxAPqvFwBVDfx6oNashiyHF
6MoieoogUIwKLvwKit6lOUk93gzPQ+Qffm2sjrWQyUELgq5fWJjML6GQpL9W6dI3MOCoTqcETxJB
MMzc+kp0PY1EPXzHGuCam04hMeywtM8ZacH/L5qGlA+itnFPsr0yzp0h4hMG+nOO58XYIRvMaGwu
HH6ZOeiGRLwzUh5DBpvDV/2FTq1jQX95daL3HASPrbeSjP5vIQJAUTMiEPyJZPREExatq2KkcYJd
ytidm4D9kuyxSaOcv+moJ2N48i9r+edaPDpD+9LAEtj2dnyl8CDUHN0JDWJOcdgHy7CENkTV3PzS
8k3DWgK6IyHLLeVBn5C1IN+x+rMdLZZgm5g0W2BuOja8wyPCKBIQtUJpzHPnJ9j53XlTP5wF4cGE
oqESSStT+1FtRqjoZoAgO9BvX93upAEMZyFNNx33DoHHoyD4pqN6vwzALP6H3jN2JF9osUKSgElL
b65u4L2JBfKQtWbC6HORqT3CNjYVtq6Pgmjt6A53fOhpP5mYxrFS9Mbi5trzHrcIEdrFRhxsqPKg
qfWjdWJ2Cynr6vEnTq81+j3+WGS1P0eJj2u1wAlSD3sVUaxu/Rn5cl8Ypn5VVWz9H9/4AkhGhZy1
gSi7bXFDFoRYifmKJzYNyJMsP51GXsPXkk7oSQ6ukPl817D3m1q69RFCMjVXg4TbEEwyqIP1RNuP
a1bBipY4JKXi8iFjHLlSCFyp07Jse0DY1fZHk6kelfTBcWd03qOQC/khY4ilN/N2y+qna017jrYb
Il027rQLxXb5NOzJvQEv05hkhsSFiIBbRog0srZq5nL3ptNmejio7LzkqC2SH3usPzbuyeoPKowx
nlIn2NbEZ3TpX9CRnQ65wNNPlPa69WdJHwpAlpUqTDS+aThyGPhGTFDGJmH/2A6BAS6xOzyWxV/E
5QNrDfnmZNyebLhnvhZOmB3OUp40avZ3pXWexQByh/wiVbObP0nkrOZZOSFqDmqfmnOadyVgBgUr
x5jL1ssGoSx7MLjuGw0ECq8qxOm/wQFpUWa3h6X4JEBrsWiNVA6QTSN/GpoXmYCcugAoMGWO+cIv
8z1Ga8pzJQ5vi2tlsrZ1YfrS1rF4r/ar6T7NQID60sC+kSSj4I3V1zj/MKdxfTJ7im616WBZt3lc
vvB6l/cA4rOGB8CG54Qt7jzK4HbIQsD1AI1Z8uEu1qx24E4837mH9jVzC8S2yROVPxO3Fgd7Wnov
aELDF+aLBF7io+3khsWDEhnJgr/6xWb2kivRMc3/YbvtYRyX/OUDc340RPKVhK+cp9o7ECJvARVO
xt888dOUT3s/A/LmGLS1rF/nZPpqsXDeQJImoq88aCECAinXyAee9qJeqKukLXRD1gXj2c7nxMNY
2iHFNzcHKIHxwc6NoRjW+xhDnZ7ehTXxdHTHBeXBitqDiKIMyzFnhNy6ulniZeHj7enpIapRQ46E
dd/99ARs9ucCCDJwEqUUI/p/6aKKGhvtOxBwGk8UsopMBqY9xIqv1jx0wRbnJZn1VEJYTs8+E7eX
SqVIfQGFuhhWEWcwf9jH2JX5n+59848l+09PwwnPvK7FUB3hJb3piGFa0xASZoAt+g+4eleIrvus
te6rPzAfLOKV0moaxbGaJA9btN/WvhiCRoajNxVR5/ndk7J8cEBKdGX8hIWtHatv+gfuttBvYYCw
WFQ7sVW5Mumfikq1+iBJq9qGmsCsLq1g+CAEoHoN3aOuUwL9x2SyMWtOeiERM4OyTJrGyzzLyfGA
8Awb5Xi/p/HMr8d/rXgzgcMxb2cSw4i+Go/YL90SzaAa2hlUkJrrcvw+AqQjqMN2ApgAVsub9f3E
jDtpxdhc2ajzaDKrSG4BKU3SXwSPF+E7R1HvSApq1cjRnVHnOyosqXRfCy3mBo59lnPxtSfjAmxe
2BaEIe5NMhVdaZTatNuBWruGrz+bTWbFRwU1LW72eDCgJn8S3PY/45VHuBTV/o4RQqGHou5pETxS
2yql5C8WEZr3gFPhI2zLqvgRPsQ1zNu9zQcYIHRHn3UmX9WHc6tyMjf63rNTx26hmMqFHJqHeX17
AIyUh9HsD8z6jtnmGOCEpQEc8x5HsAYHGEaNUXknPJEIHK+V2ZH/dLK9xb7vPGadTkjJBR3HdDiR
Hik7kj2kvLYVdQOGJHc7fVlyirLIWSMwttK+eHyjkkRwNq/Ynhib3omxAjEiDabupTUXiOSFyio9
wqkIR3tvf4UjgW+Q3615tFOVtYMf1Fy1YEXJc434sKnE2zSyW9mVPceKSkVKcdH3O5kGnm23T4Tm
K0g86yqS5E0l1jsuj9JjGzyfFV1Wrv/eoisj4eNRKPQlQ6NucOzf/wmFvK7k4F/TDSCfTobdjbfN
G/H+ZxjEqMaVYjrsB2Tg/YAQjPhPipzLpzvFkMNKoqzbYrdfD0OPr9Kfw7rQh4K+7W26OgZMHeQd
FAr6onliv9Ph2pITTLNIP65yfhFJHwwKtNfXeWP0LPihrNZrzQsEg5aql6JChmT5o+vlsTdOEMij
gRC2Y3fLa4rnIQYFUOSlx3e6RtLzFKuGCqSPbWQU8ne6UPQJbABjxl1gtyajrw4jJEusnU5nD6bg
Cv6AzeodN2axhQcaRWCxbuG3UtvNMetkRt72AcC09cJ5yQk6yhx7zvDLwh2oJxtfkvv0V2qZr5Sq
k/jL8vyrJ/48UoDYfmkkSvjAvu1OgjStplb/5l9xeJ1peWoHui/+SMSN/LWdA408QbkhDEiyC3X/
IiXgpOXQ6whUByC04NS3u6QMItd4gqegQx+mGNAO0M9FwGLdni+49iyYddOlPoViY4sFzIUlZZMe
32xgjCYszhuuTzPYk8kH9/M5+jO/bYCpYLe5eFQs44SGoHVDZZll39hAuN53g3MQGGWcZJfCWBdd
BLwOtvyjck0uMTXJ9QOhkJcVVlfL/CETypE3JBw2ndyHgY0ENMp39DXTFcFiLIO5RuxtAYa4wzDO
E/4X2zva+TIv/ZcZUHNNjniw59bp/RC2OM564lGyAhKQyI/2qXb7sHS82ZmbVJ3jBT4qBN0JIwnS
otZHU4Kj+prsxLd2G50tZovehG/2PDwXvLNJDjg/nw9xPAl8nOd9RHdpVHJflb22jwFi8N1W62+l
P2Jy8/aIQT8cR3eXjKXF253weB3BkVD8d1CNZaTlR4AEHTT8qxhcJMMI6DLRQFkDlV0PUAD8T/hV
AcUBD1C7Jd2aAu3Oks4vc5m1XYHrBenli3kU2icL00Ql83HZwruHjEhnqn2Rxyk0ij39F84+OZki
Yj6EDdyh1bOuLxRMu4nmvOA4pKOvMhhkEZ2L/CK2Vyel5ShNZ/W33gNPhnLzkp/Ng3IOalfaNchj
i9ia+EfRpQYr0rXkK+AOvOC6i2ckRJ5sazB7tsFrCbS13F3BYSQsp5z/gQJA7gIO4wBjjqv5q0oY
NrITrOO2GzT0QHBtRRROdA2DiAAY2JmRnyn/OYg65Xee89t0T6CzkSErtw4WUO2dGOLZbLJkm8HF
u8zA00j8vSGoolVwAg3eAzvJ9itOaq1rotvQy6yl6/ryub2q/ATBN43Dfnq3WQwuylQmtwV8TYEo
fwj+twy5H4swDl0D25uRYufwolSjYWStcWJhM49ekN37C2VU93ThpuUZEd95dAqcWU7StOIGFAwa
EXaZs0Lm8bpD8pkPp2dPhBg3XYDrc+mBu7STExkRccw4YkO3D4ofgSLwqcEn7MTdy+XTPmgEYbtS
tf1ZEYV1YXoPeIL0GfBSvYPr5hsxVVpwOTGnB0WLFVgN6gwFTl3t015Okxm0Bz0OnkYFDTDu8hxS
0d8wlXOkFXQYWZpdq9RNd1WCjvqtVeW0vKODM7l6+bYSOx4aH8iiHo5A084zvSjmvkI+zu/PaS5T
CO4ptzshoDEderJfvAqMEeFjGKI4GUDCRSPeIiMGekUoqG0L2beVlDfDvsZPeTtLv0iS/wvbr5NJ
Uv/sHImhRjBI2rf9ga+a9FH4phQ6DfXpnsMfHtWZykTpSv0WFsUGa1aBtFXHa7AITXwePlkH989Z
2QZkyUBOyngtjQkIltW0o5UqjWK71ip8ZrzTT59wCVVNEJiaFHIyvH3s1I7oWSKcYuZCZwunkyJI
TYcJIcx6YBDwJhnOYFM3nWeIr3ZQFCh+fZ+OV17r88J5Umd4cPQkxyYs0sfyqoRkx+D1CupbBrsU
jVI8fgfXwl7etweLNY+6tLvipiwJG/QnsPQSnp13Ods88UUkk6JVid5UEozMDAGa4TdG7ppsyYxT
eq4K5+4ZA0n2+eizJw/Q109syM7Lfwdpflus52MiHgWMGE7jDSJCcXV746D4erL2KeOjTpLIfk0n
GZ8Vvo+yWXrDZdB8CKV+s0Ngj7rdKRUTp9KyzeohBggxAzUEWjEvc0SmPdyfU5va5/GAukOqrK+0
LG4PmmI31Wxi/BDt4pSLVCxFS0+7vBawCqI7jWbS6NWoj85cUbb4F57OIvQcqDmFSKYc5syyUzeV
Lwbphqp9WTAnrrOjjsbU6Ai0eHFZ52NKSIC4hqeBF8ywsvh/DvNNcVI62mLPWQ5xiK7+xXnGnYo2
e0S/GelEUekNdzBkC4gfaZN7QhS62eykhBwS5GcgZ+ZSHm4nSiM5XPd9WZEC6FfsRE8o3/duymZB
XTi3uDdMF9JBaRzCV2Kz1oWL2TeoXLSjzDbDDcVvtidSDG7FJvlk6iI7sRib+Pd30KwO5y/bJqPU
oiM0Po5nrdtXEmfeBT2JFyEcikhl/aWrq/tsT00+u/pVyVKcAcjThECbayPkc5jDIcJH+jo3477X
S3rvbixxYVBEhpx093z9MLLoZ7k2OMBcmy/IYEL4lPpmb94L35rmGgS3yumvBVrjNx9mniqHI75v
lOlIybQtvMiPUd8PUvjovbGe4N2FJ+ox5BAPz0ixvFoay/ydGpojrnCQ0iMTS7IfbigYyxXOa+SS
XTVx1V/iXXzQh0yP3RdrnFZ8ZoDBkSrt/Xv5LEBlsu+tz+Z/89EU2zbSc5Q0485Yxx2LoakAp5TM
FaPXh+YJIl+osY6JmxSZOFi70tU46EJm83oAfoG+SK+K2GoCo86A8TO75fdfH/JE7ehkwKBU75Br
zo3HaXTWRLPMmlgSbzXLO14fr00UgOb4qVXXquCh+opzY9a0pIW5BmVCVROVyknnwvJ+D66ZzRIY
22Oatw3BX67I5wvWLEHOI+z7cYgahq76pzR8zWc3Uoko53KhKrrjxnJgyQEly4oFOQOi2oyMDXzD
ClbEhXlB0Wrtj2FhTH7Hd+VFgoSFrkke9812JSMi55QB/Z+uWZi/Mtzoax+oZhRZeDOjfwfgIAq0
YPkEsPSQr/KUkIDSHyk2huDsXM5KJS+OXeu0CQkQOLCTT7ZkxjTpIOPB4W20WN7+JoFBcMbn8N+W
yus78on+nTyqcDktcuWozC8Nkb/qLTVYFDZifWR3uUSGmJqnqM2OWPWRX7ZeBvicYbZuMKetIG+0
yose40EnPkmXAbt1AMlVASzYVz9/18S6BwgDEdRyvW80swLv2hN1qwPRAfZ+hnFDXUQgdJXDEe6/
Ak7evDY/3SAf68EPMOp9CfXehTSfQ/D/gXhVLazt0At3qX3llWIp6NhIsmUQ3yUX5l5wHRHkBqo4
/H6xT7hGXvdcyuDoN1M/6EgtQNjZ7RaWXMFqkfRuZ+0bGmS5b3AqBgRVAc+xW355TT9GMJB8wbzw
4pkV19IOskxcYCVgpWRNqXoGUWBrwYYuN+PnEHTSCZXOoXqJ5EnJHZHQIDp6Qjc+wMgKP2xK3Ccy
zNjo2CjQMrLDStcU3ZB1dJ88U2dMuzAKd2nruHTLf02/AHvLd/4RV3sgvIhPriXOxm1SWH8a6JjM
ahfw+OBFlQRYItt8zMypoD4HplegmuWTDHrtvPbiBFkQ/gGwlUsfHtj2U7z13xMIOXhw2Lh1qapJ
KvWMoZuoPmK8fCsEQp4DTZDxpJkm1t3Dg7yg8s8l/BzBCIfLoVv8JR9v/KEx4Y8gXkig9LgJHeca
r6MrpXKrl4VR6xYbJIRLERYbelINYGtsZB9VpZFU2QxQ2YM/ncBDsxTFb40bYlTkLBMlxPuQ5yKG
g3pUPGwSGyGE7pUEhK9nCRQsEG5Iovef297WAHkCj0PtMqM/udqpAwt7QXa6IjHohMDfP2398Eya
eE2XcnZWgrJhrtwO3jXsFI+6vbE7GCXPW+CYDHnIi6xEfMgc3wo1hsrxskCLATCKPhuGa2Zcp8E8
F40A6IJlwnGiHba9ffjUAffYwr+kdCrkd8YhZ+uo2r13KcoHO6COTBGaU4i+Hpj6UGEy79LBmGCw
lK6DGPlxGR425VApuGCS6B6xEmVSirVzFWFtmDrgoeDagR8V5+unjF+BT/qMvsRt2ha6ebdFjt6K
+wit9wy3TVDmJlspubueD0SLe+YGPy4Sh1vTI9xgmY9M2j/H0YhIRLu1Fbcw6d3aRwBlkZDwg1IP
wtgT8OETwjmyjrkIbK3HCEEPRbsbesPDxPBWuF8Of7Sp7mPMBRgdyZy+wM7w0P5wfwKP10Xwogzg
VeOvkM7+qWleVOj79eMkeIkXAxBxxXOaKi+70pczMVcciMXyk7ZWMXAqG4rMDXgqgmNiMoL+1pVk
OmTt/oysqzbYnxOJsNJQdVlJwEhMwe3ISATZi0QA+pJu5nL1wHGIyu8Dm+aMuZkXbSVdL1ukME7n
nt3L5Mq3WUFFJN8Q2wnnu3P8d0eTtf6FSEeYzdrP2Q0S8MU0xm+8VzqX7kN767y1Ef5qVd088xuz
EVLXou9j7rvdjJvOLq51QJGuam6WVZcEZOBlnijdLdM74HsKRRoB3IkwonLbzPlhelacYTtcMo6p
MqHkuPgQIfWyNwUTH4OR0RtGyr4pqr4iyRxKawzFsNRkxDiRjjwvhg48yqlH0o17EmDy5280vslh
Awk+00zrJbB9NzgslxrNl5aN4rZk5aVYZiZKfVLONIixI61NFzRK4XA51P+Zyhg3Q2XmysPeYMty
IJnmUwfq/f9CQ5cv4EjbYI1vzsy+wHLVXT9G778NMTJQUuY460HvmmNaO0hAQhiBNAjLjcJuHGuQ
hgKl0u8Y0Qf8tiK+2NV2EK3O+Opj8G0CaUoOzMJiqV7omfE+o/y8bS7AE7bdEeQikPrnP9yv3lLL
hYeeVhFpGiPrgkwwOkJFuy8cUsSXDWEtudEDbQswmdjgqsdeoB0CgEG4eF0Hu/9wj3Alf+2kOwk/
xEdv3L+niofN6YKCNRq+rlzFMOtjtx+3R8QdezizrY1zfWRSuCrq5PwTOJquuWYal7wivcreEvUj
o1HvXMgMLZbM9bc8qcBQwxT7EmTvh5sjMBJZm1++k8AlzeDC5OjUrFsF2VLONqe+Q+KoM2OCmCDv
tI09A6azXHZO9i+Tt4mSw9vTDTznpt7b+h4r3uw6DD4uoeoNObkC/I5SJabpB4z/T2UYVY49uUIx
hpohUh9Aq80T2/I4e6fqcyo7bhW+tGRc+xocgDzWBGwPwBLzArrcLrgGQGfxrvvV5T1dWK05ws4J
J1W3dFJiqpmYpUsRuVlldONh9IEKZZeByZ7pCVw2Bj6py5XfuVAMib1ldH7fDt0gN3+ne7GBSqv5
w8Or6QwGpbK07VC76Gn/aIeNsQQVMZSlqxh+RhFLqpeYMTvKmaSXbH/VNlbxnGD+7JqZyWGmBfPs
WL+MAl77bztExFEzT2m61mIWiOhSj44nlLq5eGdrJDbO9fYYzBzQ13iPrj3OtG2dX2ga6AlK0XcF
6u0yYxBISjhwlfpghT+Eu4Li3YNT7Ad9xH9kl7o/wOpmucavsqD7mTZy7oHh2Z3taW8lxgmw/Fme
syMLN4LIYIHte+cZKQdchmu593nndqna5A0q1w8an7/0fHWGuyoogRYBvMcHtWCZLQR6OCd6+CYl
ENmSYNbLLQs4y06DZgW/yceupuzqQurNHBqY9EArplExGv3rW01jGz0Vro4plbDtZZMo7vq+kkPg
lAnuOcJNOfu/KfAo3sT5bs8MFLS3QxApZUfgb4AWS2xvTPKLSOe/gWHgWPEgJu9ptlquqCcHBKYH
rfA5YRk6hcUmEDi6goZsvENT3uFAvQUoSsnuZdBOf5hLVXoOU6NPoRfnkGsLP76Q52LYh3AO7tI1
dz3bzHZ437yzgFOuptcX0xnon2ldshZcljJ98NwSShQxJYQB5I8OSYmj7CO7MKWf6k4U3dTEmXyc
LhSubPR+isbg0mqehLRSbib48/i6GdYzuVf7dds1akhxR2i9BbYZEtIM7wFzoZvrUlxtWqQUJfQW
agjKYf9Bqs5PzZ208FQxHljHbmRIVVQ5nFeUjKkQu53XdKRDuckmxLrKEt0K2wXuXZDqHCVapaEN
EUW8SSwuehE/gTcSlWbCZ8X0TrXRWUcWtBmfOIgQcHkTBXq8M+o6ySZREh+C3O1fdtuTA9ouWFIf
6dWKQ6GLaYdxviBpIJ9Fs7pvLbbBmfBRF6EKJzjJ48XMee16LyZqWLmTslQWNmewuQfchZGomuEe
PkDCv2SR6+LgxAxC/iTKFuN5V8eEEDOYp5EwwBaxE5YhNbSKErgd5xGj0YK2GkqErTCE31EtqrB0
WciQUAMxJc+8pXqoUIYFh7qck+ZlcydEKzsCizeUkGYMxkkj02vF5Gh9/ZPXXJis0MfATFs1iA2V
gCm6yL4s4Fj1Tqovy0hpJxKmKbb49jv9OwQCj3KIOeqS6Fi1wF640Gt0nEryMt4+OhpRQGiKt6Fm
0YxgMKpAd2nhYUcQj8Olo0smdypIUxLJ1UAMYVDVyojvCI1e9gC8pHJTX13+nPepR9v0Gqs2gz6u
/IwGRJ4P34DVZt3F65kRWSMQqG0EX9pzvm0Z9/VJXKWXnV786HdUW9Ay+Kqw7j9IK/IFWX+GZlsA
x84kBUsv3E2RfWPAAxPRO6TGP8TyUrELT8pxwP06lB10edC0IcdIELGHgmTijvUjW96Z049ockeM
aHq/qjtGmbsEctVc04GQP3/6XEJiNom7uwd6cs52bj1q9CxQHZZiv9vmuSXSZW3CUZ7wnpPKiahK
2M5kNfkG6ZVdXz9xB5V4tFtViHBAPmKMszebd6W0v6OPjdZPCi0p73P1U4I77KXhw27hGYKSQBnN
yxvNjkFlIhV4zPDuO40CsjKpW5PM2Y0BHIJuRFHGl+fmCgNCZWpUwdJoQic1kg8iFA7mAu9Xo+J8
YsZJNG5i5VE1q9b3Y/0W3bC/ej/5ZjnpTV1BE2tU1PxZE82yRGjGsp2g9g1WBxdyJhDapOakDuGv
/KBC34T3HKZKbnWfXqG6stUfblcpFE6Tpq+FkrGxS6XeK5/dG/40Y29q1SVE/bzZC4nbaWeeLv1e
2vt9v95ftkJhUie99qaZE4X/LgvZIDYKlumuNIYIFGj5VOL/60SLO17VAwi9Rlyt79C7cK0pbWA0
QdYyJcPpJ9GsEay0uMic85QWarrjKKuFl8/zZRMrwgHVc8D6K4ygMpTsy7WnaDJCgWsoDYCWYsAC
1FBa58m4RjZan3oIPPsSYNXubb54H1mQLmvjRwJSI4PuJoQwfsH+yOqRBxWmYNj2FEA6BTfNYfeg
oQy7mwQPw7xHzcKPejOcpzMMQScyOG31p84Jd8RSiG69bRcwegLFDljSIvtpo7oezdykD8pv3rUD
mKUrxFU8EZxl9AEBsvqlyEB9F9dRY57B7/vGwqGYvC/CVz1e7ExemHzvOR7i1VTqZhxZSrJ6Hd3C
2FDczqeJQ/EbIqkHEO+Yq83ro5vdCd3E2lXt4/n31fCw7V1kmLWYYGkmoT1UYb2JJsOjxYcSSc+b
8z7CroPr36ScP6/f7ET31fCb3D9mbzaZIE6SJMcV35L4C/2nR4IZZK0oMUq2DcndEgLH745bU/Sw
PyDzgDI9FGWWYpL+X5T6rEYPjThBPCug5MkNNjbuoZ+hMJWfw7tvZ80HmkPqp2Dg1F26Q9DuCVMe
F47UN56KlhHFgCbh9xpe3haoo5WzQKlRnk5FEl6jfAZvusEPJvDnDSPI+yUh3P7l3fovBhyJlPOA
xusYG0IPy8doDIDm6u70TqwnnEy2KBMjBz5rRCzYxqnrAwhQLBdbV52rhx3tKk3QcgCV9JhqDI14
JG50taJhBpBkGTYv8R3KKOT1zhPTCGUpKRT9sjDiT/Gz4gqZ6RsnABYbNOGB9ohLEiaw3CZCgx6Z
i1eLodcxsfnXCJjrH3MHpgM4bIjba5Qf0PniiznjsT9yfCtf90JkwxWXERpyDccC1qFGMfVB465M
H+YNNvYWduijX+oMhXfwzZNdzsMHyHcYepBY83KYqg7/0aJruzJ/Z1H0ORGZZHBBBXZ0oAlFC5dB
RYmruA7QGlcDjM4y7DCI916a4+qTwtLKvwshBCU5MMNrRXenEhrrd58llyOFR+H/+q9rLLCSQQvN
Tzrph63aCHDnsy/hBP1H1/nOG3anACjqGh0fPcLiuayrH/bCjoN7snqUMfj9jq0Saw+QR6rIgw5j
Pk8HqDsJp/RpZB++5d9/cnLEjUMjl4sh4L8FqeZcR60F9uuBXaDCwz8KF+Lz2bVOaCmTCceMP+l+
xAo9JTkbJr31RqDZ7d96yTUrVbxQ4/c1jO+sdOT6JdKAY3YGEa7Eof1hSCbipgvJMB0xxsiieGS0
iWYn6HOwk0qagFNeV0BTY5u9SDJunh7pcOvDsw36+HDE5ewZLnSJQieBO10knCuxN6donX5oErDg
kCq2w1rLYiDVBO2O/Ovw4RB0TvkdRYAEQDSogebWNeeVKuklVAc9sqnFn+E+j93LIyETI/JaJvSG
AwUusaU9sSL1xOzhz2d6Mj7pyb6czqakF3HWkAXSdBGpFhOdpsL3/xpdgphD5JyOADxHV6ZHZUNp
e97A4Rr52fUh7zCNYuC1hny1hzFga1pBM2LqK9ocfsU9n4hUV3vJoXxqtIyoXf73P5k7TbottFyD
PjV9PCFjIh8K0lTcmG//hCWn4Pr4trKu2LDE49frTva4U2iQrgyERPnguBptWA3auFY8Qw6z/gH3
BTPEK1u3aIU7g6WrWjJa6nzTduGdeY9h7hMmfJywLMcfzF6nlnlxgkN/vNwwuIbIXZdVbC9a93YI
6i2rY3stzgT0g0DcmicHq9CyapP8lTD8981U8DKW6laZ4ES2cu/XlowcxYJs71R3807mqVIUNJMg
gqGP1RtGNRYKnSEMv2mt8wFQXrAGAA27zpbwfNSvqW4Q95CkyWKaOyVdn9KPSBc+2U5vvhxWDxfL
eD2wnGHWOZW038h5aAdbkEV19lmakgTXFQ8yKrpyBZVwmXPcCdKib9CHGQrH/wlcfOAMX8SmkUgY
wnuB0oFizOPrqM54DF5NPbKcInaun8vRJYFPiKaqWcGknzuUNv1oYvOBXaoLaAkxOnArZJ5h+s5v
gq5iQ0LichaiG3JucMamw57wUITc7hBlWzKrSgfKP2qntUd2qn1DEE5F8Jp58BtWDRjXmogkcnJY
NAJefBB5uYcDrPymyuwVeNRygkPBebtWMrCU3BYxzLjnYcuC1k/EG6zyoZ/t9gUeqceW/52g6XaS
QstnnUZubTKnoDvBpwMV7D9IttiEJ7XsDw3Xv7+8hnpmWQGXvI4I42puGB0MWyNy8QTNV9B3YNf4
oql0BZRVN1wKEXV4DfiUYc1FVP+WitTX2SHIDBuXLapW9g/h+yVtYq3Ayh1Q1j7EH+G9vvXQ8r9/
IR2IHESHAR8FErZZD1Qzc7u3aREQXtWld1EImF8EPXecTfugmjBoN85ynYVCLKXxcn2bA0qel7nl
miuqWTw6T1o2RtEEfGteIKCWENb0FWeWdcFK5d/qP15mSEYVcpDQbZtgJITneNopIzMEWe1uXdWj
fr5KE2JGbyY03avGXE3kQlKcYw5gV/OD7av7uIHwzxZD/HOUmoWo3s8Ag3pgFBzUyQv+JsI0eNIb
+e1QcuUxbJfg/TDombzmexhVYpayrj6ZKwvEU6eCU3cWjRePMYfy9FC1plIM1Yp5mwH4r7TPpqxz
D3CS7G3XJGsAwahowbDCPhOlboyP/rH4ntbxzkXcuJYo46k1kbqyYRmHPOCH5UZBWo4zyvM21oQg
GGCBC5tNeXkG8cbVrMyq5DGp2xhF5mpxfQQscwunKAni314TMMwHmY2zPqaVQAnn+LdpQgA0eRNJ
VmmtYMTP8DHmoeyS1mySh1Lzrn/J6Ys0ue9qd9ygEWuZqxt5rRhxOGqVECwjPMc/DU3qvcoSQ+zs
rPsZEZAWsyC1XANgdslm5X75npUj38UnlcEhrH2cox+Wa5S24377tg+OzYMqNJrJDyD+DMi49e1W
mkKZwnt3zbdmSs9u5wbilv1pH6Vq+XMonfSGytLeuAJTLlCpotEgAhbFg1rnQp4wMKw1ueIU5Nhu
0dtvrJG5JDfZpppmylRJ3xXZ24dqnZhZKu9Vn5v9648j1fxkEQL3jTpiczK+yUcMjr8qmmM6ez9/
f6OEtIxIPVXD7cI/q3SMNXV+Y5tQD1hp8CRvHIXTLVW7km3HSRIx8zffHxU0oDrEHs77MgLIIezE
y86sApgC5vTxzN4KaoBDV7f/ZmAuiYii51Tk5PCy5K/71BS5Ag669o5VEeowg2C/7KvA2xW1bDIf
8WDPtZIWTuz8l4kA32/fpSL/5e/jyQ5hBLvjC+o3GwahOU6lGhI7h8ORo6ElOQmIU+z3KStXy+Dh
KKTtUaWFPMMhapvWwj3EsLJMqumGAgD/40Bzam5o7TdXlHavNJ0pDJ73uaLPmpAxYMpAEnCQN4LZ
WnF3Q8AD/tTcnU+MOoVYVJkkjP6MtNBwbcxeWbij70WsGgikBt0vxFxs/SQj/GoP7HjUDBdzfFpj
QIG81A3r45Id4j3ffuV72WIaB6kOc8I7z/0XccacKEX/RsLjVHu4bmmQ77TowT9Doa5bZVtfyj47
kZozqUT7OCQ3S1AF2G4EJ+9nuhAttK4+r8ty1SrErDD4xRC3zloZZKwEDPdqs+/mRHfeUcHQ6tsh
YMDvL/2nLGtVlFH5YY88hFBVCvH8GRci0s5jvkLa+jPnhAqqls+gYtED83FLK10iyvG0PG/yhI2r
Ny07/oJZ8UFaSC2nZkhrNMpEC4lhrHAZL4J/BJtGCUkeG0lTC8sSbFrQn1ACFt4p9uP/FXhMEEV8
eONneBgVAZURlpHWJT/KKMXLec9rVkyRLxvWFGQD77oGb/AxkQ7e1nXhYbUpkDQsynCGcreoWCls
vbFOLX5kaPBIWMjTfT4hHnba1IKZ6I/R4ONsOoDd0s5lTKgLpjThQdTbBBop1Pw5gmn1YNlMlFjz
TXRf0cEkFhm4Qmo6r33/jYdxf0kx5lFIHwtOZtJUnvw7+SzNIUAtMklj5WpSy1/ukPA0xWuvywEo
Sviu0Xpwodq+jDbSE00+HvsGQPB2i+UCYwnX+95JVGIVrvv+B2zHETC1N73i2suTeuswDyt1vHdZ
7EtW2+faelsaL2ppgUL4w5kWRrxFnmYfKTvDaw6J7/r7i7zFdSo1P69KvWDPl2VDGayAE8zrTRbn
ESHQCRIEgOk/INxzUJMKsRtB5HTVVT33XEZJN6yJUkBbAVTFUy+SeI0Rb4jxmjctMGeE/vI0dF7f
xgkfX1So21xJXUKCPPoqEGyrEjh73EbXCIGpUpIZLVT4GiNEYf87Kl7ykIn0YTQGDHH8HUlLTs1F
a5DIGNmsG9ynGNlamM1K5TNz8Gvu9C+LRXBL/aCBwF2q4VNQUQy26zkMQW7z+T9jWW+Ch2MPyA1o
Ps63tUTJ9+hBbT2HkZLrtSTvhBNgQ5mlApmprT0FUi7Wy/rQ9BAEW9sLvl2zi3KGRrSaxC6/yww8
mpuZ5ligRlvmYGEdvJHBoPycuee+q3dlIDxugFD0XKP4AgolJEoMMnG19p7LJSH2vyjw3SVD7w1P
Hk0VAzznRVSDditMJOkBzwSzV46sxQmRW8xGu9rSOy2vpaVlxCOUJQJn62DgbANPV0wR4dt2LFEd
6DCM3P+4ZX/XzRKr92hzp1RoBNjLoPTG/C8WZO86t8YfIY9iIevKQLxT7Q90Q7oVt2nfbJ6DvZHt
vuqcFdeaped3fB6ji1+ON0rTjUqabpUV3MDocdrItzlnmk2P0H5ixyGQQtxLoVlE9A8EOOSMStex
qT6X+I6ODdYwlGqCfEpYd531GnxJJdFpF18DmjcCauiL3fq03vmErD/SyKRcARjD6VYLF0UxgDfN
GoHMnlGrJHNei8wT3WTZvlwC03AQtlamO4LKpqOzMdvxMqNAT3da70HXZ2agP31veanzOtrG0z81
CtNz4qUg/FBhAdqpE9XYe2L6r4c3NYefWigyoHtcsJ3W3AGk7QyJtUQINrAkk6Yiw1Byzv87gY8+
BEHrjNw9zlfvpAtBAq3t78QPH4v87rpo69izwGaNEKX6YAuPtX1j0YTqU/MSNREKEceetyvV66yy
u1i8qJkenZQBpaab2NMy0p2oJa89A8o9cdLtUlSysNNnSnzwE0Joxj4OGZc3Ix4y9DQQusPoXJEe
IY2wat16WM8IocA4myfSXQj0k9H651y5R7DkK1pPaRK7OFbXF7eFwXBM07TE0I4FgQ4D/00qQJ6K
zH6+ZYP2bcLtMFPI+MW+kos9BMzsMRsMeuExElv/Lp17nTrg9l9HIBsfrYztIS9I7/J7xsOpr4aN
wiqXbU2kwdloV+igarM4vr/witgMxsgQcy+XfK86ujI5EGflD00ORCMIA7dDFluWWrl0QpsQ5S+E
qDgCA8RbyQzweVFO9JbTc3v0FBjb+9C611GalSikdwTvpSEJb4KbmtPKCGqid3tDl92Vwz6QpFlG
JT9+ZIJ/isngAHJhjq8y5Kn3TnRISwnMhDNiuOkDIL37UQNMXQOxnMXwtjUNKJrZvvG9VES6YxPC
qYrTJLhqiPLCvl+HQ+bmRLhMJv6j+2xB4xUBRUt+CyP1kep5P3FwjcQBjEVVRthHa/oeYfqLSkZe
FxJGk1gkYBwnDnGfBc96s9ct5hmq3nWzF3dpV2bb+9a7Vdneft6W4jA5DIMFgPnVhFazYEwZgvFU
Hk9OZA301vXzpF4iOV3RQhQK44xiokvRedPFM9JnZ4U7XXj6YTgfeWrm0/XCdPlZNLhNmZWZX1TS
FuiKFoa7eqeyqRplZ7CyCHZDe+JCyWny+4wE2QaEVJtxi3bPThE3bMhD4fTaMNVZ/+hL32kwdiL+
PHXq5aYnlmmKf741D6ys/x9Gv4fZ2FMBJ9ibCAJck9EepWsfsFWfTPzKLiW9au0JHjg0NPZqp5WB
CnFP6X7MYA==
`pragma protect end_protected
