// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:39:14 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
XE3+FErDj1nm13LCbd+za/o5FP4tj0JgcoaE18Y+NGTSSqImto72M65aaLrVmvRc
YIJKOYY9JGrYEF+6DqdyvRvAfbUayJ6Wzjyp9mExUpg3cclUMSr1szSrATMyTWXP
Tw2Tq+HuhF5JuqR1/KZW5MxEuad2tKkIwEa0Evq8p3c=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 58080)
zyUCyEGLdz9ORIeTuFUdkkUPbuYodYH9LHHWEU1q62oeOw6QWyFvzWk9Eg+9gBIA
TWHg7J9AlwkiYYKVmEvbyZWq9e6K40uEsVYvZeEy4SKRZfPtsHsIqJI5xxuddrnL
cgnbti2s5PfVr5SfIGXEZgItaAHwcakjc3o/VuDHe7I6o+KIZVBTauc0ba17cFl1
Gyntwck/xUQJwEykcX/mQuNsX979tHpW6BEMaS8ukzBnu6Y+iIiyeSfmkUEhcraF
1p15Bpz57vSoo6z6iZm+CXvOzLCCSMmED4x3AG3jWvwfeTEDQsO2zSkqZ2yTQ5AM
iVQEPeTFNLtg2FvqZF7v6MYegKNyljqLbD2y31tyvHVL8RkKi2gxTF0oxxDoRx6P
u8p0nHXLI+IlSZ4WWrqumGNBgPc8/ZvgC6VVRq5BuYx1uOA7AWw83mh2cfOX7TnE
ibJNKP26cXTVV4RNR+/7fGUUOEHmfg8Y5Hwt+XGkuZcpyWoWNzh+4wUQz3YI+K1a
fR2VMRZlCWofn50s93s12vTQAJq7StKZ9MOcyDdiuM42b1DTgEjBoqXysZPXW9XZ
FumSYvtGvxXvZzA1fMVy/cUxWsYPshGPqzhcp5mFzCmBeqLVrhOUAvmSE3R5ZHXY
mNvUa61YLLq8sWYtye3lkjy5TQe7AotIMsplRolMn08vvNDsbEt1F8YLN8qDKErR
uBgUqJy0lf3rrCSDk+COt24UmXzK481ftzvMt09WqraN29qmzK035HlACSZbIkf4
P5ks/eRljaMOwO9y51fnGzD2KvHmDL2WK7uuGPxoBEV1Gb/keZUE9epb1OytJQPl
aESCR+tR+QtnUwhszbaxW3oMy5gs3e1bhh8ZBYetG6gtTwYLvmJzEAaK72ve2yBj
IWVrJY2HxSJgJKgnzoaxerc5eShgHPZn2ptGXIlzfTxu4fK+1xgVDyPD7YTLAJPh
kuboi7077r4Y3XZ9OrFVtPllqTbG65nav9m0CvvowsAFBY8fRfDBYiERMILN8dYA
9mZ3bsMWCquuhe0r2WJWPDfLye7MHYNeG0wi6ZA/1bp2tMl4vCd7S7LOZjm3tCL9
vPs2vrKiGpnEhiD67S9zMPDmO+v51o/WO9mCUpZXCYQ/AGPzA00+8alwABkHeUtR
/03wpfNTU81XcNlx8bXWO/iVYGZPUgOmi40QwAfeIfzldJMdROq5x9qrQsQSI0O9
EzambK1RMjwvZ9fDntxFKtKK0+W/uobH9HKsOG3SZSImmAy5g7OwEybjPgMJJe/P
zKbrVePwe/yzsabjvprofhTyg+usSSmEXd5PFcVeE+aGPJbatZ3b7oSE94xTg1Jf
gqyHFRR8v8dno7FsZ7+tn7Sg1VHDdOQc+hrn5OXglsc/N+qmOpHQwcdDap0FNTGS
utu9KSYsauiyGm5LDuqMFVsBGw7TslHJXNaygDpo7duxRsp9arJAik4DMcp19Jeh
13wkhZy7xdruwXN6HVbLqdA6UMmel2ze1INEp8olJ62+tcZWevVJCXYkk+vJqURr
ps2hdTFaK1htb4+2tBOYb1D/ir00Dumbbgi0sxCzxc6BWA1xAQy0KINgZvx8aCIt
aeYOi/X3AaIr5XWWhMdibkFb83MHfYMXc6i5BIk6E398eYQIuvowtfmaawFRssa6
P754W5pHx2RP6VI1e4VGZX6TKmAih7RQ9ZqDVsdmrguTBYUZOoDLucZZ20f30Dom
W+hayVuOfJR4vNEgRbPAFpeyt3cxINYUJxEkjtmml9kM/PgLS0Uec9tljy1TP/TI
3tAQ6FLKgKdv6eb8vBzUf3IMO4S/UcLydawt5t/yJFO0i7Vt49C5iVjno6D6VKVA
i9PlMswteT9b/g3VwJigdD7nAVT901uy8aDplz8zQAZgYzdrTqmfhMIr2SIyIHkc
5gM6i+Bs7AdYESXS5VC6aPfJ6rCFPxK2gCCTHmGJInTszeBJzcyf9Ld7TS/exQ/K
jx+MDpfUlXX/xTaiNPjS534XnFVD0q2snkV18kRJ/XKaS3bxMAMDI+Tk5J340T90
5RWg1KQORM+SmKk//QwGv93R+JHIVinrmwmVWkwchd7IOH0CxWnhzAMYPnJ8t5VF
5KWBx1ZM3pKIvq4zYYLoOAOM3nXKfecdWdXtmyGNPAJvC9sF576ue6B7vxftJbg8
vVV879LzexZ7bZlJ03aO1UoM/lScNdhB69lQEOtDrHoWV3bHt3SWee2pQLZPop2K
Ls5EoWKsXskw153xtXF56jKlBRn2LVxrgKFjV5XeSwRYK8hzcYtnedsOdOHVcWi/
D/tTg6g7rJVLTwU+gpM3v6dU2klRvKYtXnR6gRTnCwOjX4++McDRZaNzlQmnQEGR
9LdyyXzmp0+CYZAslHj7qqdN5/BF0AVWqRlrB2tIL6Nc0XQClHbr7MIYJH74FVrR
8h05wzqtZ3KdZnJOKpgXynKRbPLmqd0BODe++sqLoNnDhe4Qxn0oouGIPE1iBpSM
1x+m9bxfnSJbEs5FUf6pMepUCTqLyr/U34u0ezMroZtFjITD9mhWpJda6LBbC/eh
KthD1AZELw9wMUfJAi3AnpDiEDtRJi6IhBl3rwOsO2uqfzmTyalXWC1KDIGL+ZJk
HatSJ9sjY5hYg10/mmEo0rQuHVMfzrw1zNhM1QSIbBHKCfTK7zUhJD9EpilYExoo
5v16iznUheaN1/Ds/5NE7aCt33eg8yfIsqlBunDOf0t2mRITUI8avtAoziETfypI
CrAEBlwOEFAPuwXo7ONfpM8ANNkoa1/hl8Y4fwETVXmX6Mz93asfnS2xUDirh1IW
zM/AQTQA2hd4gVKIa6kgutt33HToL3eAHpUw0ZIrjXpeodJdZ/BsFTqiXb/8w0Ak
LJyBBBxEKxV0OO4BFpicwdlY/PlxTvDfwxHC3cs0Ovup8jzbNnGuPpIrx6bi+z5x
75bthA3P2mu981cl9dhq5dwoQ231FKjpSxRj/FCGc+hFi+00sHaLHHN0YsVxHjeW
hsv37+xjgDRQJy2qOm2weAslCYsrwGZ4M55rnqd8Hyff4WGF6lVBHBxzM83hWVyi
u2x8Dl/yC0U/Uyu13huVY0zMDpGdqnWipEwoddmBSkIXqC4vVOYd4l/moZL2pPaT
88j6GQnXoXwWbHBs6QXIe/A9DRqwJVn//eC82dB/GdHFTQlikmHfIpGtnv+s1UJl
dn7BPM40KSTsc6mgNTzY5tbWtCjAP7cFTrqsCcrWpQLkmJY5fezu+HiM2qibSiOF
kgT0d1cVZXjuqbN3T7SZt3gEjrjRl8d4MbxdfCUV78h9iepqXAhXmAJ9+C0rvUmE
x6GYXbUL5yWVvMdEHE+No/rOserjQkghwVLEfglq6JB1NZKUMVnr3LlX3+vqBJvI
Nq5kvrucYLmh2UvjJoeJuCA987L2CYt6tvYZc4Wut9QHVE3GRungdD22zn6rluKR
zXJlcioCR+83vwPjFV7958IQ9cCaMKNGVmmvxMV0hucXOr41isU/ISqzWwmfcnic
wMBivPxLSU1er8AcfUDcFPoJLiS3bRYfxn5i734zvd0DUPSJ14qg3CahrN2xT0xO
x+/2hXpmogVkrOVo4OJd25miiA1aU+HWpexOJX7tvITmPSdegWPO2LegFjdr6O8M
y83SJmL1/OuZhQMr32P7KO+572VGhhHNzvvAGM8vCM/gdCshpmy+FXHbRRqQhTc4
QDMD/4u/FX6MWTJbSKQb85gFGMwyMYJIjTf+Sf+9nMrW9yh/MW0z9CvyGD7+GjGq
LmOa31YnXOFiZiU5v8i7AoZHJMuxu299EXwebGtjCQYayi7ebomGVIyTKjkA/i5h
8hc/MuC+yceXRGh0U30n35KaisjO+HVE2+V9uZcXG3GfYxApk06qksY2aBjb/EDY
V2gL2l54AwzrGIfll3n0qRMJ2H6gYiOMKeIZ8VJRhVQ0D5ITDWRXwM1uwV6Gam83
Xf1Yv8Mc8tVDMuzJkro8AOzpsMmU7V7LUPrRSblLfQ6WVco0k10bKLEI4LKUtpE8
pLCT/jLx3fXYLo23suBVBrBFrqkNA+JY5bJOpGXgeyJeMRGdUsa+C24yFyT2JlH/
bsnRIkwVoywCo71z/tbP+WjLPCoT+gyscMkelEXcTQMR5/aIOSSDgtHgOjpO6eMy
RQI1bD08x/7OCnHYxtLJsUXTO1wBkOTS6jBM+nkodBHZdckyjzaLQJnQpRII+phL
2lWm6SAmF4wIE5JvX0/3xdHMMiLGLXiEG+1yv1oVh8NGrTQR52H6pNzZV84ej/QG
25Jb6S7DR5jLusC9HMvE5JFwVNmJn35pQN21gGW8KpJNMQcAKrkZgnNQTZrQRT+S
8w205Nbn12LEkHaHDwWETh2ksGryqNuuER4VBzUu4Y2XiYvDhfvCPuBN98DfFSZc
hCAVJZZ7Pn0cpL+GYbbhOsGKN41XDN/7uEoL0upPgjCio1YuxgDpW5wsTJrbiuzo
4GoaAc7nsxM6JE4+Jn2Q09RmffDq8wrbL1v0/WEuExKG7mwoOnkg3+Lfi9fyTqm8
zTE0oXOysBkzBW61sPSrJzDuiChZpjlAD4qcnQAvGDhoOT0N/f16RJU6oImH5sYc
NLu5j7HsvwAZG2o8MfPS36nR0jwjwHxdRM93Pp5Q2MM0Bh9N2irUHA7nn6ErTI0x
ZFbsCsbh1a765NPcxb20gpnX1Yho2uRmrqM10LeZjfJX+ZLcxentC1WVFPVe6TH0
/MrbwOj/2sK4btIf5+SvAynbdhQ+qV6LsOpHakR7t17iOrJ/HuifAMWkmaef6Zyo
c33Um2+/Hym4J/37inohi1xdmWHwFuM6sb0f4WNeuPySoejPPRgsYSa2z8H2La03
4PGp/o8PR3/6IafGJTR3JAQn786r/lOQLYp8ZaGfYzdkSmvjWT0WHC5YdVTfB9p6
zCjbOrv5JCKzfESBN9N20Mop7wByhOoAN2ukjFq78QDgOJFks8D06IXv0rG2XIef
ye0t9SGJzh+uEr/GoNm975ygBn1HoeMnKrRa3Kpmq82Zq/nFHjWpjEDz9vYO5icq
lccZr+HIm8uEXo6BatiehCxL1bTzWWfXJhTgo2pNqHFHDHixFlIMzc+AMJ6tSlYl
k5KHim8hWIEAEkajq76UV9EHYqtplCvQUy/8e6qYx3PA2aGcTRrMjp3owzY/lBiT
OyhQo2sikk3miENZpoBRD8+CQB4+ubQcIUkgGlPTyq8LVDsiIsUonZHlz/LF7lAY
iCcQb2QyaHED+TrddRHr27iRbP1ResikiAp2nzF3S0ypV+THWpGPL6OvrYXIre8p
1li8jFHxn/x7XSlW+GrxEXD4CIt4qOtXIxObyLtGrzNkmIeqjVAoOEmNyBR9J5OW
1SI1VqjGWq6O4Zg6u3bdVtPgnL+z31JMkaqyy7ttSXNnJuUnqTZoAmuTTHhMT72d
RwrvJjJ76FnAtvav3yacfl1TvwxijKzyNmVLAx1G1z5f7tUx6DMtlyhqcYXl/G28
9Ly5hWl0cPe18ZsrA6u+5+XWEUe/pXQnmnb7zysvvXYl6j4RZ8SIJOlUdmEHjDl5
D2YyUkqg0sZqD8bjZ5VmP+nEdp+suy5TnUtIOWfe3bXJKhg3nU5m/sOPrCzMv6j4
rvgYtOzjrXu3do2sCwrp55gW+nCfAbApr1PM2CyPwF5sEoPbEcWtxfMTx7hHM+Wf
71WpVZ9zRAoEkk+V9yCngA8WYDd4uMg1T2MwCX42l2/5OPGhptIvXnv8X0LdlPTp
wRqCtCyKUwhcCZuevrq/y1itam17fTWYRugpVRn59nmmRKjphxS5Hzf0SsjAjXdQ
nNvqIXN4t611PAMbRd9MBrYnFSdD+fdgp45Tx4Fwk4wssRPrqp4TTMZJPSFkXQ7Z
2028YJ51uzvkpsX13VyySoHngjB5pyLoCr6VztTqW0SWf+FIRnYAEeYnl3UcWnnn
ddhg4Hw4O5YFMLdS2HoDr/dCAzUTNprfCH1Il/j/SGYGyWOFzEduhuB9Jjje/pxL
RwnAe1NUkYSQvE2JMkRX2zQiaCYuoEhmYBBvjYFya+BZZwziYefqiIVIPACYEwfK
h3YCO5u7YezTPsNJpNmpt4MC/W+CbQiAuCfq7JneRxUa9db82dlPT4LOn/9GSo4c
fs8lAuuCboHweIOS6mOmF4AX05WKWetZUanyOhsYfBuBGVvIk1vdxYrHMRrUzcwL
1zSUmPldtpVtOaDwXFmkIKiD4oAxfhoP7t25cDZz54NbcfTB1rJzzp6ugSW6e6ll
Sw7BI/8FpO/XC6S0m7+N/6SDdNymE4BK7Y2RhSEY+/wLvWeQHaiASME2FAowq7ug
YYyp/+sGdVGVNSN4q9xevWjfYJ+B2bFZqcU+PVnUmshspBaEsKBWHL64o88OG0sx
D9vOVxq/Y0YM1XFbYrayOycTeDsRxXFvzWilFVjFBKiZTyB0/iTwl25aA1mzDQql
TKOAvijsr6PXK9Bilk5XA2fwvVJ9SOjSTHUX51EKUAzY/Uk+GewoPEtHtKqiuj4Q
T+rMCBQN5FcP8O+lIP/tihHXO/mn60LZ57hPW11TCe1zk6FYKqzTqxuQ5jYdhjH4
jnPZ81A6vEMHLNZwW+0ePR/AQI6Ni6Zfte49QJ17Cp79Lmrl3rWOSrYB7kBGzHEF
QetzLEUXaU31s23u0kEZfD1do7s3uj/0jh609qV3Q3Bg1PSah5xFUYz7E4s6uuIp
rz9DYx8YA0fjr1VIUBjVZS3ptNRfEG8PvbbojADA3qFzCgsOnMTiCMuOnoCcT/ob
5oDkWFrUvF3mNNNem7gK5GiY/tMYQKSJcOMx1nho7GeztTOowFF8sn2hHajLfzK0
CGtV/XEUxQmRUccaOrRuYKuemyRdKg4DRg0yc3zfs3zVsK45flOwTQDqfAAuNy8E
IGx5TmSmSWAD4gjlSP2gJlcN0stEvWR2j4TM93WJepmKoDEvkytFNvBUnZak1BJU
GcFVgYnLLZF45JyFT8zxkFGrx1ts/DK2fl+aLHsOPYVkguXVhsOYEb5hs4M9oGIM
pic17zLsFf/LefqEipEapoQFGq6y2LvTXAqnkGHAJiK/FeR72hg00ATZmIUKazMJ
oy7Nvl/frWRTNWMRK9qns7ifOaM8IDNDVmuOmY83oYUmE+GUpt5DXt7rjJ34Omh+
8noLFu/mTA02dqDAcWE7ScrFiUZQGaR1PFmJ8Uj/PjMV4gYdmy4inQfeFchgg03t
Zgl4lP02OsJBAEP9QFUA5mJNw5PFTH90CFyO/xbQ5raO3TqpfEuZVWXxK7xXnJVK
LPrKdd+hI+agSEBL0W7xlf3vGMs6+0HnQAIDr/vYhuQOfP8ANDXkywp2g9NcWEX8
bquIObLVBBO7GVbtDljoZU5gqgBhETafIiiPxluApqE6zpevFpk+UOsTPijgfetv
QeeofZgq6p3/TZCh/wohR0ac10MCbCLZDVX4SwVMSCNwNvEXYiBRiKuZxzdsJhhz
MKzeijkECbwt1bJu2/9SJoQEciIPsZaw0FZqzK2C5N2U6QZXH9Q/vaZinXn06NUF
OS+hfW5YmsVnwwsCU7u2So8bXJTHDP8/Xe0MK5UrApzTznjOoFKnJAe0fdP1Fg1l
7t6nvGE3OhmXfI+9ysCaS3DpUjolkkNMUQQfD/Q3b8f/Aly1IEUuhrmcZHDoBvvm
60OKvnt0heVYWPG0xp/v45YHm0vd+pV3ajqOScX19CJTqEIQClNRxPMAUX/xPPV4
VWZrvKjpiBlgeGL0j9AH2VVzf3oCNveOQDa7qClE7rECwPDxPphSR4uJGrjabDqV
RuRcYf92612yBT/sDRJXRH5RKTwoJiQArnb06nl6Tegh+z9RhlbNdAtAQdzeyvZe
Qqi6n7TgC8ORStoEaIqly7t6l/jhfXB0aCvV0HE7hndY63WthwQb3nmpT8CYPm1m
u7oSdFK83AizLQA7l6vaC2HWK6+gmW9XVQZcFkZ14mYCSednTlAcX+VJyNscv1Ig
UPd7knyE+cx3jx2hw2YYnH2urpxdlZOLrGp9V2aS9Yqk1BRNAnQ6luHR3Jv471pq
eFHmWpWJpu6MvlylXOUdvTyKcqetyEaZFkHoAPQYWtlzakktpShbqpqHkuOKwA3d
KDdPZ+iPbGwOCUtqdWO5piOHfaFSNbA6lE8y2m5egcLMVVWubLTtx1yXpoTdJrqu
QQmZmd8PIdoWvbDIbESG5oeeKpr+w1VAjACj4Bi20AaIGSeSa3MsGiG+9sQNOEXz
ZnPQcZLlhlvyt0XGwfVhZYJniyTSkfaVdcK2UWEpkPRayEJEpCidm+vfBpeFZ4Qp
TRQKvo02+ZetjExdNwfU1Sr3aNGzMWlCLn6YBi9GIFWPF16GLRefLoQGXxTTRCgu
pzVdaro+icZBtrP4EAVb2slBlnzS41bH+oK7Hxdw36D2417JGdm2hWxJPghACife
oVF/Ic+tiqM1CQ8PqPww4lWZPBJCx+KRSt5TLdfB0jtGvc4c2MekQOVUOzAjQfrb
Nk2yUkAJLDjqAG8DRCVFqTuzAS8Io2xh4PGyYZL917RxCLkKhOgTV4zscQAPAOTr
RpPkpl1Fv6AkaTYC+AJzwxJ9y/XP4wpcZ/PIZ01FRUGwdHN89fO9jjfYr6rNupwr
XrkLFmnKNUT3P5H+I+dQmyQl4ekRUHqiO+xJaDZSo85zXVUgLk1Mso4qlzstbIuh
6nP8YptONW/LV1lkTQ2oSDb9CVa6NFePidUdfQKaxGTaN35eLEyLfP2xknka7inn
/ewwqylqNX9U8vz3PT/lPdYf36s4YINzr83npd2mMGUFgFlPuHP6fX5A1AmFy1up
LYb7l40HgNP9PNhWqpnn+7bQ2YKFMjvH4YkBOGspeRmtULR00k1So684VS8Lx3Fr
BpVc6LAYldqoVoELqQ8dYQvfSQIv5MkVBuYk/uQMTnnJIGwWUeFlzJ9TLke5YBDd
cJyT4eL8jJtWyhzPsCyzuqjNnzPcPe8I6Zkyz6ObzctgL3C7DtIdgPC1SKEbN2dv
vcXAXG758omrXT1Uq3KGoTi9olpUi/E/CywUXJVtxdcHtWaCU2uf5wGcLPvN1JXM
bVeXF76GP0aSPrg7CflHUAxp4g6OVLxr34nCLHifggVVFzJUd8Q0Sd0KiiSjWRbQ
MaVNsqTScgmK31S6pLhWLIGXUMNemiavm4xi5cinBJHyP1kMEmNDWnmc9J/cKmQC
kKK5TWhQL7dGPicQ1Z41y2UuXlTPDyiQMW6PJLtqyx72oX4aYLUdlOy37w+T1ywZ
xN8f2HPFEDLGlEEi5Sv65awGQq0DE8+Y8r8R52aSBons6on9zzQEs3plQEzkCrTk
dPjg4kO52NkLO3CKoftOHjicL28q7WNBYHf1d12NyRhoh38M5Oqdv3O8YsLJdZLH
pqLZIMSgGwRdbCVTbLcg2oLzoMSBrypiltabPYE//TLHanUn6GfN0nGnzwJk4QZd
VjpQJrj4wWHNNfMBUfYExjxx3iD4gBewMigqywRTAUQPo72+vLllYWGHpAatMhu9
TzhO1ASfVNaHPbkhCNcpYvakou4Mk4m9X05HK24eDtMzYqvdLYhgKrPQbBhnW8RH
rveZwyb2UDC58tfTsubSszLafB1fvgI+BOLIrJfxBS6nzXO8b7QzkerZgEFpydJk
FEPG+pNZI3ZqLhImOFSr/uPp2nx5PJoqxiVQjncKGSmP3nyb65TL78c1ZgV5l5ei
cT2nj+5mkKfouyLzaE2DbG8XAFrwTGnDlBJ+ao+ccImLR/oKewHUx3d1iRj8ghLK
7HitMf/dVahto+wfrR+irdz6leWu/SCV4oLtfzY4ZnLCv8z4kI4QrZCFnN6eCOJs
ll2raahTT6Ps/vnpJrXZzV2jMaSB6ifJRkaZQLFPCYYGTEnGfOLkNQNtlEEkHmwo
ACfR+WIsugLC8OFBvPV8nyhDzNYmFQRiq41+NUAZwfrVVIoXvVWz8bM+r4xO7NuH
p5i8kPr+6/Zz4Q0pO05jrxH2Ej8YSWlZ4Iq5G+dIDMVurKfvm7GIZ2qMroDboj1n
rJ8drYWlkQOlMyTuED7YRZ45gB66EsJujdd3IOsx2GUDn7uOvkBxqRNIeu9l6yLD
7EYAekkhyRXOuD9Dtb5AOj5JyxgslFbpEjlKHt1tckVw98lM7aCIZuxop2yC2Gdr
jpdTW4O7L8iVjyieqLhj8F6e0vcacM03CoNbfuXuARu2x1ztyfJeSaNnXhf0ymg/
ugMUhmxonJPQ1fPFnvihVi1LHRY3ure/Q+LMR9XQf5Ygg3M/ZJWt+haNMage9Fqy
MOAvjoO44kOQnJ/aXDcPZGV4HKsvQk4gyJdl3mdWAqlNhKlt2rVmmUIu9HaUomaw
jJE5Se0dy6rdvJOJH1uLab4Xm7K7cpQSju777dv16WnIbzHieliVRZDFvsu+5yLa
T2/zeYGizD9FjO2ocTmDXqqw9yxNNYYzi2Ijd80OCt5DfEcdk8MaR5snvbe2GNFy
a60t0wd0a6V2sq4BD/NbhWoqO5A6IFcF5WWG7DTE+gkti9Sm+0RzIgm8VqPjVtYn
WMg/PC9BNGHZaBAFUMXm6+P1agq7cH8dfVV8Rby+oAflCDyxw3unvD8ubtbdSyoe
MPzxuCSvFe/ge+9Zqnd1WpSL1N3KR5mvB/PX1YznvYXb5wnE9qTtYz5e3s2rupoC
odsshZJBcdtDurDkEZtF16JlL7k2IMYrnyKzgGycNdXZr/trGlMjEggxMcublm0R
yhyIKBwH7hnYCD2LYBRVdiGHBXSSfjlQg0VmRrEZBx6n+WrAvZREszk8aIdJA34D
wT57kw3dJU23GbHD0NLzUwdAjDKuluQFA6SLfzEYKsSk8I2FOJDhYIdM+v/nOOtd
vqeMBJ9MtSts4AS6K3RJX/c1cllquy3Ydn8iKJqsfhuZuNIlA09J7Y3lDjRDsQ2j
8L559hV290aIqOAtgDLMnowp2hEAXMMBbS3MX4rfABJ8OBEcFhPt7xycmjFJLMI9
lKVo3psFndUI+K13tMT5gB/sKh8krHeVqOTsQx0dVZ4hUnAon4k7+vopBufj0Q0w
HPNPrN2WBcNoL3kFeWwQ3Jy9uVKXIurcnKj6TPcgu63zh5cL5qKQLi+HMZEU0rwm
6rEI8jzUIntBLPeQCp7bhxJuQ0tmzVyWfvA5mY9vtuDpnxX9pFoIh1xKfqoKHeuf
4e/r5O/MSpE3E5YKo0QRt1p7h47NTRgqKXUr/tZQrW/nCEvExIshNFTHssEUQCw0
AWgQxfqe3KUcvWAdVGTev1zSZvO9r38zmOOmZSBekKAqAGn7j5BlyF44ygwDPPtL
liGlleWkHCD8m9JGKoIwwGiYrItx36zeN4GRnumUM8upBvR08y0pC1WhSTm7Upxy
p56TPsWqoiJ13Kxcz/SvldT9AJjAl42JGuXWBTA+QRyzod2cgMnku7J1JAvBHfLP
TH3kzbEhFY9LzF1BT06eHoE/KhfDW3HNb325xZEhXUVNxYndgy/ucLi+8O8QO3W7
4CQjq1XQ38yT+Zv5W90FV5wXVNXh7ypZZ3qYnNwJEsGNlP+T7sY4LqIba+PEXMXV
k+dokfCdeSm4xNQaVrJH7Yo17n6I9LI4KVIUZGMruFvRteTrYLps8exjAh3b+eDw
LHyhYRHEqm9VaEokZ1iA73daCdHTOxnxN944g+7rxIlyJlk8vKxaz59IlAAItsGF
CK4Dj/r51NWXjz9NWPpmNPHSy30W+hIviiwyq0rpwarrzZjKGi8XFNtbrev9MADi
v0QNlEqsZSqiYzC+xd3YoUwQQ6pAgDWXw5WR8fEyfalCDVEzqqp+aDXNY1ABSSkc
s77tHPExl3LoKOfik1iQNol46/oDOHtgVuNPB08dnsROI6G2u9Npb0dMb19HbcS+
/ZHwmj0GxzD4/yEvDSOcB7w1W+2frbFaM++dW4NUgrv0Ghg7RR5QVY+2MSK6mOZW
9o12WZFU6wzbydhFaeNRBb/wlxtHAw4+NK5DJG+kzieXAU4QfIG0iJbQN3hHE5Ql
adGm92YgQ2Y/GDfs2kxBprzvJczLMkj5qAabI8sH4HzPlNYiLbC/vhUG5yQJpJGZ
tPpdWUqRyibV52bPMeVpz1vWynfo6b+E7GsmQeyh4j38sY0QBup6O75ITsyTM47Y
l/FH/jXfQ10TJEbKNbaYVBs4SdRL6URN6FQP3U8lkfztB1TMS5TFgYLUHyHaO/1X
pz+vOWVR4oBY53rVYJ/eeOinMlRniB2zej/cvavkkhZM4gk/qboW7Q3i0gaQchEQ
55j3ihaxgNP17Lila4OJZDy33NhT147BYXH4CdlXkJ3dml04mL9oo0yE/r8BdvrO
2XuaR2mpg2g+hahHbV7ilvbtAi7STcRJYvSf1y/OJzLGXSifMhFaWVqQ2vf+aHrT
Q3VN3N1zcvDhhLhFvjlI58iDTy4z9DgJoWkOCr1Mq84ywyRhWzlIVeDiILIly6D+
a542ROHcYTw+dNrCs6vspdFaVj2SI2/ZE9WGT9wOprwd83EBGJBnFse2XU3PH61u
/nSaYE7t2vXm0vuXI1IzbE1x3ICNwa0tpWfEs7vcWK+wQ1h+VoTDoaWGICMuZ6iv
tU5BRsJeDP+M3zBJ5lJvhM3fpGM5npAz2STbS0tyEPCVoZlkoVGo+cUJ8F7iQGKa
i5aZymuPrsbJ8WoivzillnFTPiJ06b4qs6dZ3ojxB9L/2RsFn88E+xckjvaWA7qM
UT7Mz7qwWGwDtA9nBMj3BtZNE1EZw8iaDztDE+sl0JjVFjPMtys/Kn19wrZ1Nxqs
lQnDS4AYj6Fpa12eOh18L2/Tgi/EKC69J3BZ+BzmHsVTQa66lSJKHErRQPWXEKT4
AFoQBXhCwDHZh1/yu96/nFI32SkWUxQqVNm5UbD4Z9kHsNRi1X/u4r2BzbNETwi1
Qj918egySdjA3cSoHYb347pJx/Lxrwk13vxDj0uwuZ0Nn0SjaV21nhPAPJ7jebkY
ccd5FhYD7W7EzobtRPjMME3AdJSYk8gkW5XAKi7sU5G5qi5luQv8UJDhIVoOUIWF
Fh5RsBKwlVyJvJNAgMeeGOiV0ANetJE+e3CCXmCiiswMsl/xfqvdXXzN0RxwtzwI
UvRIvlsGPo3ly8qBBfBpwse7lClDVuk5pGnrWgsM2hjHTfQhi6dQxX0dw3IIy+nD
TLVBD0PNR0sguc2w/i3wg9jdIOFQ6dTFw+04QD9DPn7aJHQoJya6y7i+1ko7gSw3
cjaEgwzjLa0C6DwqLgPRHLxcPV8y6YtmbGSNpsqCvJjLzYv6R1E1uxWBNa5c6X7l
ah/wdNTIKWBuqel8MqSsBcfmxlJ0IXyoahoNFGoebVsb2AsCaAdJmNg1HnKyNQ5k
c6z5417XTYOVKPqB8g/xfOPrxzHBBFvRNolvJqIaMJq/P4ZDPY3XMG3/3CqqKGtG
yFAneMcCk6j7LANOu+EU6iSdQNA1JecoDzLGw7d7oK1pqr2sTq9fdznCqOTI3RuQ
boCqYeGtzxt28r0wcYVoTIRzQ57DM1R1eJxSBRjk998jZnoFUo0eoKM8jWVByx0Z
7iZCsqKGVfXF4CQHTaGcBCwpcbth/B9rIs8V/2UoCLfC9dLfwfPKS//QfPJDUfOF
NEvYoKxGXiA12gW0zzRE1gYTfHOCdcVsM57dyfMER+b9/dbCY1Bcxjs1hpe6iTRA
ZB6x7XK9s66cB6EbDaUa9BanOZfVR2bD/T0zJO1JbPj35bHoK7jZxV9e6u5sVf4k
fWNtdGn5BcONGGGT1SExhrDChD+/q1sriIvdVXJtTy7MT4yQoZo7npGrmAkHw3mw
PTCvnAj7WAi092Adoe/WVnTWFJCEJuXQWrmtH2Qj6Cs9VGEGOIokGhdwkaOSKlOL
pW8zMaxEuia6CCkDEc3WzqzeNzwkUQ6Rknbkqyl5tWyqlMbsOGw/UY1aUaZpn1z5
0vH+MKdM0IzxtPgazZl6ypYpkiiNMEl5+ou9+w6OLhJRZKJ9Ugzh6kbA0d241UCJ
3BcjsKOQoPxPWkpalUGMtYLbqqKTz+d41GysmIZPygoP1nWaqw5NdEUbnL9z17UA
pBfCiQlNbibXQvGI2qnjm7RnaeX6ch7hs+mV/+HXFQxKkFVDhCfQG4FacdX2W59c
I0q3fEGrjIBR7KjtNIthd+6tUq7qVw7xuyvgwNpn/x+4COduDIBkAh5IjzDm7Pxl
U1FyO4+HnQd4Qvop1BqzwQg4XQApH0OrmNDAs1D8y/cl1c0eDEjJqSfO6BQKCT1W
CcOwgaowCXUThVeHRWQxfFUmYXFV8o7cnTW4FA4s/7b9ytZrH7mJoIn6sa4Ar/b2
p2a/f3BjDaS0j2AINHrzMCnDzV2qkWW5ZlqZD6nsEah38mkJOYvQjaxfnOJ+hMmv
W5Wnfw0c/FrPk7HNZIv59f+J9NOiOOGIU0XgU8nsxQZS0ltVygf6prMGchREowzk
/Z+d2xvv/5oHVfg9z5Pg+74r6BhOlQtyWWgaoPwP46cQaWZokAlIfDR7/VkadrxF
k6jrCSRwzpc/IFhYzwRokLT5LdeaKFOxiHDg076pE1EENkab45cpqNXHu8dS7DvE
FjoPGtCEJnC1GYySwjoja71XVA7IyLh9d6FQfCAu0/lxxq1OuYfmyZi4wXrofbOz
HCrB1+kdEThFDoGK/ddxyFaeXHET/XZKovBoBJnfigRmQiTUKBZIsG97RQuFGsOs
CC0ZhJu7Qtchsj/xoVg8f8mYk0SUJXhd3FAUsT5uqUC2IJ738GifsRxtAHhI2PlJ
jDv99KUBdg3PQF8MTpncH/e4fhDu6gEsXcnEhPyU/aviT04U3X+KdBwQ4XRbCeDb
Pcf+vuQNkGnu2V9/ZtNfiJWVfig2pc35Cu1zGmL3e+dKIwxEJ+BXif1ZPTCuAkg/
NU99oQOE9vdb6goIX0ZQM1sARKZ2kw+iVZnuIJLgTM7DyUDb0OjZrmXbu9gzi0Lt
SJHvh1j3mcxnP+mwyPJNoEbtLp0lhL7N9kr+BP5aZEMEfXO+mhXAr0SHPm7BVCDj
lvoicMwP+/5VqwMcmbg3rdbLq3bhGPS7IgGCO9wPWojlX6nGi6n+HUKYcVPADmxT
wwi0J/fZbUOs88fG6Zb41RNN86/vxeZwf3DEenXpeiM7Xz9TUAH0l+HABLezy6iK
Dd2l16HYrwtTgsTXEzPXOHO3rd18iftmXPxDp9DGrgP3abRDfxVhemEVVkgoOal7
ww3P752wdRqb36AMsEWBA6HNLh75PQePt3WEpFqJpPPXYBadJwqeGA4Abr/3L6dB
aRAu6TOt4+SDC++7heh6x2xHJUukIYkRwd9evJpGwhIzB0de6rGEDMIjTO4VO6JS
z7G2YNsz2Odc2zDmbhCS7ZRjNHWdNvxuLNyLfRceMmYDn7vy8CRKG92umwfIpXp6
4uUfjeF2y/Pji1/CUwJTQba0lVoCgjqqaAQzEcpTQaH6PTs76Th2LfKDpdqjSfAm
60H/RSEvP2VvdtjBkFMCVktCoFB/Dy4WtdyS3InEaJQJUv2eKrQS9tPndEmHlHwE
0I/IWQzoC/kVP1gr9Z1etHlUAArseH4xT8FlgWET3J1T98gkQKEMQPGstsXB8XGq
gxZiVv7xvfdLOGZW4ffPd9R5UbxCYbDRjEoav5CnY2Ki8pwn4V4exqyI7U4NmhAi
NTyBKNxaPKPqi0s2Smk9y34YKoqinWW52If85fpY59/6sZXrYxk0bYEGYw9eaRfa
LCB383CVShTziO+rPZ9VmPx/o5ytcH6HuiVsFozozn2P9hblPwoo35gvuSZsrzVE
33PD+vhlihOqdir9Mr+lUxG71boN/4le8UlwBxm1L8zJ6isNpZ3M2f2I7gdQAm1w
M0dGuvBiEd/33iEu/y3kaiRyzt4FzMvVjwFHgfswH1FGsWUDtWClMhYTuYkeTI4W
wPL6QfCNfX0zndkdF+gXjUvyHRPi+x9L6IkHRJnfGuMDbk2WqyFZKZTm9DgrnyEd
6aDN25c1IaDnnkZnCV/wlxK2WAiY7NA62RPr8tcVjAbcWbJwPKRA0xuMpR20ukmm
NJUij1RAn/Wo4JL4sDuctuCcdjExb2ekpPrvz//PPlK/+LWaUb3tfLKTPs5JSMHB
PPiL0GJQRB2iQJnmvJsk9qNmnb9L4H7Hwe4ShJuX43OtBjwLI6+yRFLU1Zfw9C/d
frpGgwVoBVjZ4eBHfM9i0u4OU8ySZib59qV3sEIQ08pVtA6g6oiPAYnpHFkqNSy5
weWIv+IzCt03vS54Ma5NS429gVqZ9ZBqvRLCPXIa5gxISwo3FfGdyNzOvydZhczx
Ht3pBxLSgYeoTSJKsnIPA/SaQqDTGsELbLyKvh/4bBkMmV4m9x62HX0ryrDojkEa
b69+D+BhYIA9ys9Z0JvSTzp6xiNOCjWE9XW1raTo9MD5yfo0eyWj87MxppGtvAK4
d2jWjlNoGAh5QSbidTns14xddqKqEicDbAlkCEoScmZOQiR922aVidGfiCIragGN
ZcZBoe/MpH419Sd3fUyPeAJqJ/6tzjax86+fNRDUETRJOV6ygv6waVJE/CqT75Vy
IoFXPwpC+ibOUJUZ17O+xFQBMEfUktCS+z23ngUBMMFeHJuT73Kh7sVydM2+uds2
icGmJixJE8Ys3ay+TCQqK6Q5dciV86PczNYM4frHYnpE7VpIti+u4qZPDn3T64R8
5G1TMtbpD7HrTQ3aECde+B9d1ODJ810kms/V3CRz06zu7DAUX1MpXVLa31gzMSoh
6PLhJwrudPfwrf06SmKgbzTPD10oazRW+RgDdO4q2py2cajBQqVDBE2wLxq3NbSx
8A3FDULzh4YrIagUgA3vab4bPD5jlMCa9IKOIO7YdKTtsTEN9plL+bONFhx/xXga
ZBV2dYhOEbcnPileQEEPkgV6gB6cE3gjbgJZFG3z4wlMhX4KvWS69MsQgrHmGJWU
GD9+eYbv3R1+3nx1jtdb2Q7NMPivsB+o+QXztoGKlj+ntb45kB/xQx6SKFVFdl0d
S0lQTzxubNivb6vznQ2tTJtgY4KRxgLiocdvkrs1oJq4sgC+jWO9p7C5WmICsILm
l+KH5O6z+IYuxE/hNqV5qfRrU2QjEap451fAzkxqyyflvWpAB34DBTZSZhc4qvAK
ywkRQBqL2S/LbbAcHuj2YfD72nBgswmEogct3hnc5PP3HGRQzq5wFvz1L6o2v+ws
v/Ymghk5aKo2VR56Fyh8pkdlruRaLxBWWI1GJ+8XUclYFNCRLlAB4GGfI4WabRhy
eWyPBJ938gKtsy/cCaa0L1vwZLpmak7U/lmnjcEnsIpF+PFFQCurouJIxyCK3/7I
SjgqBzo3lsZd6F7qHlaP3u0d/IUOGAy2cakkp7a0qeuN3Bmm21blGtOIi0y+swze
UAC9M6OhOC4CaeJ+z6pAfdcLpkPGY6wlOmtF9cMnmomiHnvMfho8nIbFbn+wtuhd
Yu4kBL30wqmKnvmXFSnasdBrSE+9jvyx23WA80Hk8OuPjrqdROVB4p1cCqpidPCH
SHac9pUZpREp+KbS/7a9vj5BXgbQ5VBzgHvlGhkgDMHDb8CoZgYU1r78k3O/MToi
p2JkZr21jHUpr6OJrCfl2FigAs4hDGhBFo2xpDZrjUo7POT8HuGpbSS9Ii0fQ8dD
GDkEwjBvcx/2PslGTOY2WcQPdSHrkxkIm+8op64fJ2/RFBOnQQdB1ZtWkF3XUlbJ
XLoa3OuB+Q3jBIgpTZWqSJsSBy3/q1BEb/vjr2AXenSVGD/VVv1h2/LiOLkud3ye
42w6o6og0ms1DoxE+NvwbLjqYHYjvBaYwljiQLE67m4HCSXwvJClxNBrJ2b0le0Q
/QZawFPKTU4Vsgu1N69ozALRyz2G9LVmohQV0YSj5uhHdwueJUeJMRx0AaxLP33M
unb8dH5r4rso3ayh60azwULdmPNz9/8r5IOjmX4ZwTkqYnh4rQ6oMs0Rwu7HG+VX
f0Ly6cSm1wPhtIysQFHlDvX9zuirfC5pkQYxiDgmo1m8PmX+/6M1V4pDeKqYGGiD
awZmUPbVyLVCkHE6I3lBcJauf5UpPSoNtNJqmLqcsGAQPgV4ESBfhff4D6I/xze9
GD9ZqyGAWtxLTQ1dJWzLqq/c5/qRkiS5aMMA1t975LgVlhbdkDrsQU0q3PiJ0g9E
8/1vqa9Bx0F18IklhurW6juTOHpB/vXZlDPcOhA1yrNQXa1orb7bCuelqbkYg0W/
00FW11s5zkxmY8jJayAnkZAcq+A3a5nXgKWkWxce8NSKndgtCXV+kmttw8Lh70KG
iOgJ6j/0vbLy93O9JTo+lsqOyBhhlLgkDI4F3fCqMungicq/PpIjPVYIRdpvYqH7
RsgGvSVtJ4MtRsefjyS0+twdxWvvRItfO0oc0zhAKyfbHq6MJjhSdG97LptLff4k
SpHu/rYPFBOb1siIevioGNyL+sR9Ue3ND3KBtfGr5UOcL+s6yipqyZEt72R3C0sG
QJM4hv2SqotBxY7GB/k3qTRYtzy5Kr6Ov4Wz7j9DLgjqL6ksaQN4newbxqO+fCe7
ssxyHoFd6AV5WZ0vV8KWq1xmnJY9aTYe2o4ADjRo2ng3Do9CS0RmEFUpuxwWF4oY
+fPzVhzaIPZYhv5brjJPmEBXo+lG/yuuaY+OJrnkhNphdxKHPfHF7/qDsKGpsH/9
aRJgR/YDd1aCSY1SKjvmklQXQ4WS13hTDcid5xqYu08WAKZrL93XY/2c3ClzCYbM
cyohwaTV3cyMnkLb3eNJ/zqSu9GCEHSAhnzAUCNoxyIE3uwmuiJkOo0AUUINntET
E0yjDIivaswM96COn3GWNNY8zi3a9xQspMyeFFk9FXV/Ll8p1/6UN8hdgYaekTCQ
VHdw6COMUSnIYdgy4ekcfyFw2wz4UIHh+V8HLz5uURjp+2oFU12ue0JgtuoZF52A
Zw+fnNrXT+CuZwLrzNB1S+Yy6HRu6/mKa7khc8mZ3mk/TaOntPE+XKeIuDvIG9nO
7weo2O1XDtfHM6j8RVwCsG285a5/eMG0giLYdvvOcGNXVn/cpgLexjES+0iYULXx
RrlV1TQ8DBQeku4qWpb+EXGRz7D3rQWEt3jVZE/tgN5xdRu7mTDh7jN0XMU9v+vG
u8d6uMvDLza2CyC6J9yIeMJnPn/+iaC/h5U5cwn/n9h7XHNR0WGZD9Jjpxk44dma
WsYeQosSh2ADVvhepI0xu4ij7LwUWjjQWc/nQjmyToJ/uEoTL85vkgU3y+zzxK8C
/+MPqTbOnrMNoSUrsSIkz94zQO/urXV8YDoUgUqI1j+SP6putB9WkTKOe6YTx4Hr
EDWGh3hR79tb5ot2TUHeXJR8VLp8wq+YugnOspaqxs1b3FBuRQQrobntHH7VJfUn
QtL0lFhXStMBZzV7DAP7RfBpM7KMoBPGCIF08ZnloQXrSsVXTtNcZDA7JVmPAPf7
7wNbThl2rNPf2ennn6YIAsvfcmHtOTgRourja6EjwSBSN3YmwNDpdb/O69s3nwQP
onnr4Tqh0TzO/IWQ4d2uldprlYDMkJSDgrd3sqNAlmz34ZN6GUj5nWyYj+3bsBTa
xrzAFOq/8IztwQ8GDZp6wu7W8CssEDEZINJcxvpTFNkkNClT7K26tpoIW/Ov/sRh
eHoPdH2w4D9ow9WkKONsQYwbac8D4HsKg6EWUGVkSihKYmKsm10AHUTCaczC01YB
cGh9vPyPvmVyDusHjYzK3SxOOIJszOqbdxpe5H9SzPKWdyQf7q3fur0UHjp2sfYO
Fk+LQHbzzOW60TU+Dn9p3q5DPoxYO4P5XdjOuoqmNRkkn0U6mfrHybz3LR2fDr96
V1AdFT37+JvCSAp8U0ti0Mf5NKKxrI2osOVLmyGug4qQgielv7vJ7VHVpkMgci0j
pNWQxpQMRU4LyHRCT/9ww3T9rGB2Q6dEetK/pOm7sUfOTcchH6Xx7qRGiUj7a+TI
EmgD1twjXT85JaJj7wqJn8YDafhtRfkopDChmeDLeHb7lSKjYOQovKPehH990nEZ
Exwpe/1SV/+v5KdLAU1Db4u8IHikbzfuJueOmqcka1vRY0Zqp5FSX1I/+1zUoU5P
hqYSD7uFws8EfSdGncU9rz5b9EFnhizk/wc61+tHqkdkjB2zirn9n6P3dor8m8Nd
b43aABEOUdhdBTToteRwrzIMKz+D9ZTS2ID9xuOKJHtvzMlU5uLVkZXPdjIgw0y4
Ui0oLu/lhwVkVXYSrYWcK9/emcBMvAK9REpWqZjyptFgLhXMLKKfuN/8pfZfowDp
c9k+qPl9XsazySnk22wekQBopGH84rKFCeIbjTuL0MH7aNDbvyREo1max4RSLAjl
l53+eQdU9CDrUG3eXgAZT1w7i7fFo7dH+6XreDPiSo69FrR44jZSu8QN2X1ak+Ks
jtH5Z43nfZXWgKqPFWgAVJAei1USuLxSmE4c5z4r71gnaXoeUx47GKLYn/O3j/kP
1DchzEiKZRDOH/zA+BHisUjaNARJa0+LhbK9btyRS/0w3PFgW1EyIzMmquFv7bx4
gj3s89p477sZ9jtkEtetf++R7Xi8vAW+qCndf3jD5yW/ZDS33gNTPk/BgiOM7Lk8
LUEFppdLN9jefF+UbQXJtKqKtf9Zid4h+9KePZjr61tGWEwrKL5IZG2uXv+JAOD8
MCTI5QpwtvzAPugqQp7q15cDePa1u0VmtzdfTzHgJ/5MRUOZj4qjT5sM0OLw0vyS
TyRmNtJLRgMmJ1dFVzBwNeRLCq3AdOMaqiJgoXPtPudWg8TGELc2fJjkY3xtTABP
vAzGgumROzbqJnwDMy2pRgHPsQik9Zq/OTu+CJyctLa2PpElCQuZ7KiOYsIwdpsP
Ejcl2WfeYJ0rF4qtlwe1HP1xGnN9VlrLeYpB8bFfdMyVALqPq32cZp1HygWBmIE4
TQERQ5+xoi69j9Mi69WiNL5oqYpqBnaSdL1JvbzJaEEjUWkZB2a3YZ/Yu/XetBr7
rn3g/EFNm0Yr+EbtJr7wjhoLDkyLE1ZzJ5t/cf5myvLk0VIihkYja0Lkn/uTtFfi
j1PcBUCDOA0FDy2WKTZOj7O1A+BCYlDUwtIQEI6O4Yih1nKmUNJm6SoAOzB+h0YL
F2BO/sDYDttSUI1maWqI0nlbDfHHPJUudkjIiRWXWorIPM8Euiun+IC/T4dwc6mw
sNZEXb3WoSLT/yjdG1aALRy4PU0PgFH+Rsf6WeMea1WX4QKC7QCmBED32VWOeBKN
C+t2CqaAsusvR3ks5fbxzP1M36gCb7Rdj+UtbTeVrZAPTvvsMMLtTM1XM7ASB8qc
VnJASR0dLwgkUNu6YDCcKwcD4OCV6rjAAcvgntAvR1PlHXzrzNxq8tBMzmSyTFIH
w0WL6T1GqPu9Qd+Q3RHHUKr42VIWROw+mrI0j4pvxv4ZWPXjnjMywS9RXe3xg3Ex
xzJkorkweYtARiM5O3OJyLrPpWuGIfZDeSfBE7rZfy1JmB1gk8kQtK00ampz7af5
t2P1cMP0O4kl4CvvfdI4ZmtD/8adHWZS8IZaeziuIGNErpODepLGzMs/ayCq81NM
bwl7AvYR097Fwt1MDvq3BJFK+eUIEvqYzeZTE3LKYKuRyieyZLQKfv18b4ZSMvHH
ics/PUYyOeJTiZ57Lop0kZImw/Zlq1eIujD9VxKUX5BfEfA/5EkuB1xPeW+ICU0w
Y6+Zp4pDOlJns80dQzT97pxALs1RlQ5Rxujn+o0Higrerf8uwd7lr9OUbuPkBYXl
FjdmjQwy1LdyOS1Yr3yOQNUTUOONLBnutNNQ0dAI2XFNMqnILfvev6lD660uE1N9
nYsGhjtyBfE+mrgVWIxz0Ur/80c+l4to4LamLtogvEyJZkmQS3uEaXnU0uH4uOUt
V5tbsDMm29bTNQQ1ZM0hCe+L8qwV2L0SY2ZtsL3s6Wxzmc68IU0Tl0r1xIGNTXnv
XCLilpnRRLSARnMClW9C6i8YiEyTWwNrCE+11xuhuLaEqSG8AowSvJLk56NTxCiy
GK6pweH5YUfDeE8bFDvcbUPnGfxiZJzdK5BgXXWJzGUJYGmkIOS1LDBkWqMR1Wqd
Wl35Mo/7AmI8le9vUCDS4LsJ2g2cKYYbjW50f+wo7u7xaPhXg97bO+RehIMKvCR8
1qrDPLW1GXRx45XMwg32/+wb9jRaF7qoEsqkCa02vhAFG6Ua788XRNu+3Ge4RgSx
oqbocqpUOlWTeZEIsHay1PiT20vz+LmffyAOXP984EnIS+lxTa4FiRMFxSmLCgks
yOXDXH+n8VQLupSbXCMY6qeqVbmlM/dqyBXllwe5e5JNOou8r33cIjq1i3Oi2hQv
uXc3aw4MHeqNvvCRlpFLrPAyLF+tk4iwH/Jaq0TtKueAuw6iTCDlS97u/8efXcYA
leGQJkaYhPhW8PWDuLvfMCL2KKJaHLFffHcTvQYR28l3gMOFKM7YmjUrisq7VYGG
92rGixwxKQlXRK2519Lvw7NUWnKtB1/ifVPi422UlTRKecBdrcBMB0GQ8K5eVZ8r
+ZlVkfQTgQlxuWEXQcZj1uMCzQ8BKOdxX7MydjRgDH9DYD9wnYfgMeMY4BqqFnsL
cTU5VDAzG2dDgM+EmFFaCEXYDBihcKcB1K/C0zlxrvUPfijqFNYZ4Qd14aZFLveq
IpVhreoOPZQEQSlsOsGXIvRVpr7tC06gWPmSmH5ivcOUJ+cjaS/uO4G6Iet0wozZ
BB6u8MoezFA3I9MjeU11ltZnRGO6d5gI0UCoqyylOZU8WGTcgpdBkjOiMFgVXQa5
rxlUxTOnvU+S+iiCpiWSqsRl2fhpjjju+iaY25DJVOOWPnhv4Kc+JddX03+RrGrF
AFXt+eNXHjGklJ8sTBrTh/MyvRCourEh6Vmbi/JOYHHbQAYMuuN5xHFH+fbT1IRv
AGOy2c1Vd4iCp8s4MXhKV5K2hU+g4WiUv+4EVJX6WfCHILSTcxQOnWwrokFi3lGL
IFKui5EmJL6kAnKAtMsiIK2nUVU5EzDg5jryrxMpcXehRiXedgtz6piylFL0rb6e
wnGz7mo/4wq4T7xk2h8zdLgVHVcrMocS8YKz2jihtVjwkjcr62SMfYOs/fanu9bW
nKOwsCH1zF1THJnZUACc2V8cqIqkYjRqLZkZGZzUd0NqpralmmW9j8slLaWvtPV3
QmTmyOYoQNvnTQ8v+k0U2bt3+R66xSzuO2uBzRiwd7hZMBmeUP20MPBMpOZgxNv1
VBrYianR2Diha2M7mlYJiUhOQZUs6vk70tyuFRM8dv7uGIAUfA8EZ5ZJXbcANB97
mnPZr+/B0mcYUL4GWBWrAxEyelIBmcI0lqLkooWMxE0DGDS7uacxfDlKlsVgvott
17QwupEzmssCfnkCph9Xv9ks6vmX8O5f2UENMNacDfiBApX8IX5m4Zb6HD0oJjHH
iGNDrh67IJqLkPDh/BU6xsgauYD83CRnf22GxjB7othpdtXPObgJs8pWpE42U6Ms
DnevUNXW2DTaz8uhWuleFSjzwO1w4yK5gXv2fDc+71SBshFgLbOeGRyZxo20Hy+E
K8hRmRx9hmB5VN7zbhSL2JpARQvOyMop8wNXesT0ft3ZEUpWPGZ8n448WLt5G24P
p1wBT2hmxcCq1diobfshVzL2u/D7RqXngTwVY+mfuYvbuSb2tDbg2zF2kVkeSsdL
wRue60mJMBc/Mqqbx36irBjaIf8b8YbpefEIe4ogQehZnCa4+CIlr6vBj4P25lBV
g1FBvb668VgtFnzNtlJyLpkq3uoAIgmyFLBfSYjvysvy31xn7YlnX9x7lU4bmO9S
W8pNoUb0CyAl8gJPuoZ4oPFwKR5DdsLBO6OayfYl8hYX17iB5hgfMusDK6lqzMJJ
7MBTc5wnpFCW8n7HJ7IV2M1YaagxebxJnu5v2r2kictCcRrWOSsQfAZDkvOOo4TN
iHIbp2nZiyDZi2cgHKZCijA9GPMnMja8goYUdVA5+C1FMgKWwUaK/tL4I+ychw4X
WFULF1kVsguR7q3li+DLIV1ri5c2sPRPInGGJFncKMwNyi7nQ27Jl722+7AbChn6
UqjYOVVyC0ZWa7cUpLO/BxDF+27Tm8ygLONmkEWdhdhCVq0Mu2kD7EUPiC5Wus16
kS+w6czOnfhm5hnWWqFZJLHA9OIz5byu8pi0ZfaqT+40RZgE+0dZ0BO7hCbUBkLI
MvUR0kQ9upKdIbhByzpWYKjMriFN9tvTa56npRO3i3LyTkXCMlcQl6SX+Q65sVU2
P25mV1oBgoYGBZQjYHBuGLciSs25KkQmyJODh9YNkM1NA8X4RePFSUqvMHiWm1jC
Vdwzj1yJhAySMymYcU2KAV5NPvPD36IDHGRZ1uk275VZM1vcxO9hNF4SUPxZVdjR
nrAT8GFfG3QCyegO9QPBCkc9Dt3ycaHUhdzWZDtPDom606Qa1hA5gHAdqKFKLpj1
fNpFlCmpriM78Qk+tbSQ4bbDsZw8h/cID6yo+etbY5XYsJN6ykvb8CODGYo0uwz5
jRJGrYYs/HV5evE6y9YE07BQV9uYS4BMaKCi21TbwVIIOhZUpSh3Bn8McYpphxFF
V6ypR6TKXOs5VEhtdnQLqr/1gkqvuYaK+PtQ07nyXnkHDZE36katJXMDKbjZT1QS
3XhT32XnX/gt4ObZFukxfFVBERiYgxxcA4GnrnHQCWS32cmFkeWN74tom+ljbv6+
iLwcXaZXq6HWlXbi6z84K8iMAd7VjXuArwvZLZRBUQRbI9W8vDYUnFkZBn8bDJSO
UCRzuJezs6xkxgxgUfIUtEXCRG+khJjx9zxuHAwTaw2YlFVaZTIW/8uvuNTBa3TW
BtuIVYnpNMV1NBG9lpigpsloUlGdQ2hRu4ym2K2MbD3x4YCnDUkaUMvo1pBe+yJr
NB+GRX3f3TpPlHVaLGJxVziWllcnyV6T1EN8QZ30a7a5HvckaY/BY5isBb39q+F9
uD0R7TxoJAXGCg2uQ/uKR0AZ09IPGe3h3eUaTwl4qvr5TctBHfLwPyiBdA6AtkOz
QGSd4y18m7VQRNyHSG/kxgZS3z2Pv0MMeJWxi+B2Q/en/N6aTUPWO6Kre32mXaIh
H3spiTBUEeq0kEvhbK/7pnQeEBoe5q2iBNmSOyhlA/1QPsPfBRRJ11q3ewHvxWGL
wDABP+hx3alNgR2DxTDfUYTDv6clG0Fyowt7f30WG3zVCW23AjEj2zT2/DeFVJ+r
b+MoDb4T23YyOFzcp6RoY0uGFvIQMe2d4g2CwgY6kv9osm71/MitzSc35uLzTgHi
XNsN2lLzWP9zHnpxscBRJno61HFZ9iUAuOS/AooWAzaoAQ/D9572U4tMuFVNzUOY
vNtxCVmldYljK32vZ3dz6ZYgGY0M5nQIPhoxttg8n7nnYjA0ROiwkHgNlL3X2LuM
yXib3iok8xJ1IyhFaCYww7BEQ2laNh8Qbozr5j4a7ta+IzBLOeXfTLhX2YO6rauR
LfSsYF+hx97latUTnb/ZJjMgVPTacMmrOvjKYAaHMYrRjjOC1xPGE3LPyejLfzWA
IglBHMH8zjstnmWHevR+9n0fR8kKb3im6WTRDXgnVHHOBYdoWmQuXOnsTKkP7cB2
OTt0HsJDlY9P0ZdeZBn+yYE96tUTu/6jhAr2L7T2P6VYXU9eAqF89DapP3bytC1H
1Mz+HF9EhRg7CgceqjA7fddb0QK+EynTwoyFDlZ2yRa7hXEiv/9JKbFS50rz2zFs
m/erTXgsLOb3qv/iy7QA5O89z6u5JsWKH82hk2eUeIkawILa21RvFIvNNt8j90vR
DaWp5wGVFzlZ6mESnd6zU5pNqlEcNOLeLKEGSMKvr3Lg3eCmZOLcFxtIQMTFig2X
9er2+oAqxpshaJ6Jyku+zYHLRgCeYjDW1nZm41qUduTZP30Q1KxVjKayBA5rKdU5
tt/PlCJ91P0z5zdp/I6jrjzaq4rsJr2HvbOxGuCsp3NXWdB4CtGcCcuGlwQOsP7E
olGciAyBv+j4SZ3anvpX/dKlnsxf9BVenDSNC4HD2FfNbIXGKE98uyyJubWPiXzU
nc+6o9/jziZALdBdwbxjgP3wd8VV2xiv+Z/7C5fUh2tsesBUS1b36mpb29YnMsp1
4WQfGZLPWtjNvtqxL6Z+4qR4t5jfmwvowwFeuYnNNMzSmM1dSmHrQ0ifeIFvuwKD
/JW9bZi4CB4oX7ANvNccTYd+Gm4Ism3cNoVZSRA6a5fYPqlEZKq6MqfVxCZqkwUa
6VGOvAhP4pl8zfzBZIOKHdJK08Ma6ygXSrP4KHcBJtIUgrMbqFHov92IICAkkHjA
A4wc+IpTm7pOkWPmUIlTdA09kMdjkGm6b4UdEQOmwYzP3BNqCMXNFbJrTVDDSe3I
sVC0Jveal3yjOT7uX3KpCyEaHSykvXizeTNY70v6YqVHPRkra7rGhTHPJF2ug4Qn
NnztNIBQ8R+NibQPcNXRGoUgaHxJ03PlJbVHMNCVkNjwkHAVzVWu1YTo+9NIraSX
FquCCfcY/kzlGxf8qpNVJ6xqMb0logBQ42G5RceDlDhOzO78g+9nQrcyEnP+5Kb1
/rDPECiqGUkd1dqqPpWcm9etFF8UcagbEcweSsTNdD4v747jmO3bNpngLJJdhpUM
i02W8cjpjCh+zE2AE3pncTOEkeaxQjnly1y4IhZpzY5t/sOUE8iJT67MkT7HzWat
nhVfJvRnGeM2aJGxeof0raXaGZi6XdTgyGsMJ3a7BjONyup9VTYlsXSH06eXeWtS
69knJm0kjNXartCbOF35/9nMbPT3/BHrYks8QkEFDwlN27T0x+YDmyJJvZYK/bmF
fGhkBu9OkU46iEsAWPfgY2s9dybZNGq2UA66tQ7mz1GF3Oqs4sjBJOLeFS3zcCIE
FKnAEyJXEY+EnHhLsNDUqRXn8iB20COD1mDoK1AcCH5IK75n5UIhpkpQxj/MCOTO
pMGoHRlMjh4X3jCUPzNQUClthJyt7MvP4CjIYBYbLaoyv2QUyP24z9j0J02eDqCL
hK3chOyiGxlWqsRgbIzMpfRf6w98F2PgJUqjOwFPMb7JYzAP4gdw6nu17cZ3ty1r
XffS41XPMwpOdW3QaqwIesw2IyrufLCDOvd6BIXmfbqUnZZOaPQ2OC9/Z8TFvUta
ugxT8PJsJthUu6n+RAHIVGe8qygOTrpxMFbHFA0aJSiVKAMDroO6tKk7QgmvAGdV
aJQFTQAkUTojH3VInllpvPGm9FTjPQJYMv39a50L/uNsuFke13hQ1Y5gRrxGZgZ+
KOoWIBJZL/vbiPMK+jGeK1t8QbX1CIqb24cfxy8Xh3RWuKs/Qyx7o1mBmKK7lvut
2PR0niMyiOG/5ioAaYp40yRM9WdPo/bB3DrY4QgPqqd0by/etLr5X/L9w2xI5Nsp
BHQde/zkUc5M+8qfDewEq4ne3AfK//rwVtDY3Pya3jlcQ1I57rbOmWt5Na7JFkTt
RdE4670bnYBkoROlzRg+nyYcJ6I8EqHTzovKdHG0gqR/HBqhrSuBPcfPSTjGj4ZA
gTt8J3ZnMs1E52md5D2bFTTi0ZxXdny96/Ulwo7GLVwYsaZfO3wS3FuDD8e+XWun
2upqE+L/CXeBJzyYQgeZr/0995c7W04BgmDqoyxga0g1DZdcsgXSAbriRhxf+ptO
CAvwJmjlNWZvmTLm5sZu6KpFXjOsOhgeoHknbj6IQg1Lz4i3kDmBuKFr9Z5xto5C
UDlrDjdyG5c9mwMKiDUA4rnjVia1Ikzp55CbWJV0dPQfU/ybZEd7udgjTiUhozjk
l+SK5MUlXCIzie2Os5Bnd6uzEem+WN7vNEImnOl3ku3JL59Q15JqYh1kni1AHPLx
OGmwxo48crlq05KRV2u2/hqfo40MRVdp12Lk/a4tTfNXejRodUEUsUUODL1qywzm
vAUooNcV+EFCa406vjnQpNGjFm3WS0P26xW1TYj52O1W9ecNXdlxFvRpekKgvRMC
GSxLYmuCWDtQimEn/6vaRmhb64f+9wbIHHPBZ/MVY8gjNYONg6KGpQo2g+AcB5+l
Bc48CouXrWlW97yNEb/JuytceUwlRxcIS6lxl1hrCLFA9dYhk/sTzINaNOj4uaTK
Ze3bmOPKrMtadEnSGA3G1iP0rYo1VmN5ol2ET3PKHgRCam1EVwKzw2RwyzhFxJN7
AffcMoYqlzPZW1oy603sjfnL+GU7n3z+WylFi8Bq5Rie6VxfHW6VvuhSjuDwPVLR
BvmK+Uxi3yr6lc0sKaJY5j/987eFtNu4qGtg1LmwMbOcocNL7dXwbsS/7qtcDcam
FN0rbJKsM5Y4hNTkeSVzbE+1oiNiFFRW2QroZEimORvlY7zY/SzCBOGuoTwkhMCy
9q36mTCTSKre78CEKvjcpIRjSSoZlwZVyz0ndlTJ9zPEjyTL1BBHpgMzBIAfgjqW
ZgtQJzCzVbX4W3M1jrpx/m3P7AaKuXyvsuVg29abujhDfOMlqaa5fkFJEZPDeN0o
L7FVUpi2Uw/mlJMog1C+ByS3G2pyIU8d7dXlykwK79LUrqQ8R3eOsSZeJRwJaVY1
fCNkVgIDPSVmckO1QHsH3EPDl7+io+Fr48inRxW1wJqlPIc3773D4fEeFxgfHPns
Zb44UuZxE8EtsC3/SZ11DcyLm/ozENw76xxhNH0C9ylAhB+8an2cBo/zvW2BJ9Vb
o8GQt+hLXMt0kTUGN2ph9MLflb4jUHCSHk8KV8juh3H0I6bLIaorFyD6gmeQm/ad
o0I6/xiriEbtyFPBwe6IX8OTlU2tQzCMGI9oXqn05Sm6X6ZHnjNFbbvybIOCsxJC
ROETUajtoUr8gUhpj0rNn27IG7pPgQVE8fAmPPb2QJwXSXUTwg7/FhwKo1HedIF6
1HpMoHusZKOIFHluXqdV928usrEbAzIEnlq6QfjcWQZInzEW2iltQ1yNurYERXqB
VNTctWGeJBvNzhDlRkyXpCfy1Otf/WokOosdB7/IXG6GEV1KSzT4IQSkC+DlbHB5
2TMJ4dauRoRsv4a92Znc/IrhQy9x3N1Mrwlq0ANQR2DeKR51n2CE9zpyML3hQX6U
Q59aOoX+oFY+Yg4CmpBlXftsbKgT5sNmiVHrHLPk1htP6TiKDudB95OppgUnOr9j
oHSv+BWDyTRVdZUVPRvRKGQzFJkqH3PrRhOtsOTLP3VBWtkXb0xugZy/b6Wqcu5l
hA5TIYyZNQ5KyNybAHGioSDmf+1GIhouQLFyL+Z2BLlT7PGRU7RnET2W1F66sulC
4TJ1X6qpCmR1jxq7zZ69TQaGdjS3i4myDe7UNNMyUiVDS+Y9Uil/j8Iw6bEfdfWF
s9wtkLZUbBZUz5J46DB7LqFjwqGiHRMEcb9yeAbk4tvqQFT8kuhmPOzE4oTLxPdD
lQSY/3hOGH22HENdgxyrTr442ikyu26cYh5R/7uvYnAnSj6RGyDPH7DJK/pswY0G
O66P1cmell8reprl7ipsh+PBiAA4ldF1a95voFBemycucsrJtPiGbkz9L/PKUEty
t0n2PYzgM7QKAt0j8fIO9wTTxAgXhnnEoDG/B9GrLSg9qMYOUYIub/epmLH72S6X
IDVGG75yM09Q7zEPL1JX6i8MXNlPJpsV17n1rMj6mcWAqQw8Yjsbo448CV6u/sXM
2htp7Z6px/yBOKPApItIzYwFoTZJrdawOegNMYYF6Y1jiy/pMsN02XpQOUfupdw7
7K9oW84/zdoDRmh19ppDvGEqc2D3yHMtSXIV+wKmx2LBhzQ1O577Hcw95v4at4mI
t3qJ8cWZXmtOezs+IAhqeKHdg4TJfkjeIMtNCyfxy+CjcISUP3pg1qk+bsUMaYBJ
ytHsFXRnE8isi9diztpFI6KXfbAvVnitolMVG7kWQvjSIoLYK0GE3Ve00kS24ZtA
vXCmOmYXjxUHR/IIi8S2QiJtzqxgmDdlpNWZBZfnVpwiyrnlrxewd7Mx7XsEq7oP
twRQ10YayOqSVclii/+jbKHluKAzlaIpld8tmFGTGEkdIuUwNGLbpqoq23T3bjOC
VJZN2D0c8/4Gdh94g/e6VQQr23jsrLWe4URur1U1tni6XLHnnpl83ZovDzWg8xAi
Lu2tbxwvTqLxzgcH26MABp/jCBf7hAh9MTkOgN/Ng4aFe9wPFGjULNKm2oOII9Sg
mk/cHkyadlgH8JgtOLO7Bppn6P4Xvd6tiF+f9bAFY/MbGRH3ptM2wfpQwLHM4BK9
t8gu54cCi6AZ896BA0nuJQbGOAouLxNYB4fKQecbJM5byQmN+bz2NrjKM2E4JG8z
0QG6N4snrDm94/RSmNrDGs9hePMBeFTcAa8jIJDd3VXxMtkRhDhvZbDRTiMtKFjp
KxZC+Gmljq+TuA32XxB3jaWh4sYnnd5+PhMW0jZRGqeT9JMCEFzITRRmaryNP9wM
NtEf9bo8xCrRjKZWFhv3l/PWTG1wtSQ9269V8lUeSg7+rxO2shJErMRWQuwaOIFO
3l9wQfmCDlR8Vvrjna22pHo690otKECJU44Ri7Kp5tYV9FsvWHYujBxWfkEYyw9i
pFrDbILslVvrS0sLqjNB4Rl4d4XGhvzOoVExTcGTYLTMJsqbPijIEQIrGurVnBPe
1EWppdAib6zzVi7R4zaxCc3ZIZOiFh6vv2hSabYfmQo7at64yB9UJD1JedHj1+75
9EzikSwopy82HASC7FFRqv+UaEpGT2Tp4Rf2Bbb7LyVp+c51P3n4AkHMG+AjvJEV
84rShoGiNMipI7GIiZFqJEA6cbki0nwJASlmc6GwyGhzVY+syomxj7ywVOj/ZPlz
6FFMkrPeWJ1HFEqy940w9JlRWo1dAOUCZGDctn4hIuBi9Hlw4IgkAL7wV2KHIsdH
Xy0Lj/diyPrGy3Ikl2e45jZlgVMycbpI7SKs2sgaXY0F1JTNWHpvmWAt1yBtQ9E4
Vz7QU/QQAfSTV0mZgdA5yy3wCMAY/EuoaC7+Viu1lCuBbbWUAprXoOtd68su0z5T
T82fe1T98UTJKDW0w9ncF6DuPgFL6cfO9esoxjVGb4YbiOWoZYRcIYx6xS1TjI7w
8EgFXbJZZYA25kdYAZE6SDIy+7ZioquRtPdLPQr+X2yBjMoL2BExjQky3ccQ/7N0
wBNdbtCR++DFYWqqmurJDddh7YFORpr/pc44QSr63PhYFR3uzB/1xBsK/bIZabYI
v1+FAQQJDHE9BY0WfLdMDwRqqmLfut7y+6OUL+XWwrvYvfEBIm8G3JgCfZzs+2G4
oBU0lXu0ZScGLjAmzZ2YUIJpQcUvStNU2lRzyHTL2iN8eV0FDnbd2RNL/Fa6T8aR
lACNgvkwquPQr5bYvtRzzmO8oeHToWunBDLnmyARdTSX8/zPKknxmf24keeOGGUO
sdGcf5OTnmEG5XBfQLJorb9lM7h//E/3QzMQ+hZ0ZVVAdUgkb+dBsaVNwW2FbdLE
GvNOluKReYR7zSQtMGStIOPP9f6KPjFjby6zK5eA+1N6lrC0I22YMkPT+/bx1GFV
mySLVyFANjIQYiISPpP5OzX4/U3klkUVghTq2BB0cKvFhCQuWulwRQZ+U+kcv3wC
aMHZ8w8R09hr2cMhrocj6VlC94F+0PLCGHFVn4RiBbY1uyph4Hyyf3oF3RQqxHBE
vHE9gzl5Npqd5Aawo/yZdeuEwNqV7iIUz9hyniDKs0y8ZZn102t3c3eUs9YOWd47
y9lWu37wIUpEhJa7iMNLXlZWzUw0672BxuVPZicWiuEvn1eEkDbXJ3W4BYqaDvZY
jqlNxMAb+Lw+R7r1IJeyU5D5i+inleZh8UoQrQlCLaHkB2wQ9x67mh5/6MizCf/z
TZUqRNNXVQ4BTmlDEg6BlmdZUiOfqpf6pfPEXIVSjhNEaz8fGCPUktWbM472grAq
KynH2f0riIgkkIbIDdviNe3n3KLHWDbLLc4AeHeU0KvPsafcnWTBG1raWF+lERYW
RrerPKuanjPJ4+7EUCAGwcUm2nbGMj4mGqBDP1su2iosXK6h+arOCqpIRt+wVNqr
G4JCX9vycOmaK2OaDucui9w41M6YqndgSEq0eDAMFjiPxXnyKV2PlMMIpbQRnQPg
lzFyWAsEsAvwLWLMzp4OF2snyw12EdQlSqf/6DFlAVs0J236YFNIZVC6PVebN+6W
EK3zhVBo7OL2/fZCGSUlQoEwapJKifHW0Jtc1sbYVl7BlnP4srYmAn7w+qs9aIaE
v9RkfxWT1KX7aQOkefZcCj0l7CONKa3vclBzzDxnpZ/L844UcC+Zfe5g9Uq0WTQv
rEQFfangg5lT+oZmUX6LP8X5crw6Q+eAKhYBClhNk0xpqOohLTCOP+G3HUn4DjWd
lD57liuDOW8e1dzVr6Q171arH2BAp+HzMWND1zE3uaDKHl/KU+7AkqHFhPVcTUhC
PIdQm19dLAdgqFKFi+U3kGT1TyDrzXLrkzDixTAZNxNW4sbGPLTlvZxWJAM9N58b
v1WAw7ihoaC+u4QPIDNjIrNC8/nF8vq9+NM2IoFlNu65KojegGMuBwaeDdEdL4qU
HkRoo53u5cq3OnJMs7RSGbMWbgMKCfOqRcKKRFWRuxWg4HOE+URyDmoZB0eiiWtR
o+s8QgBmYp/4rN0Cz7kAiHkEe7RgLznxnawlk5kyaeVqMhMrdnRW/6O4S57e0rbg
jjfqiEr6aV+P0jwyJTVNfRVvQiqB0jZ+EXKv0TYCtfOueRzRTjoqhmpni2Z8g6le
a+HzxHnNJpRvRFmfn8xUoPrE9ZNsPyN/PkuLDWhsMEhOOIXGrjReGulExtPwudP9
2grcYqjX0Vfnqyn79KvHgNh2go9S9DIMiGrZ8djlWpgA1MM02IXJz+cQYIMsXn9l
cC/QemrSqMaFKCtvxmTgKtevOLhivy8iqhqOT5MIUWdhd1zIgH7w34IEdpZ8n8+R
poR3ZRS8oCeX4hVxOBkqDfeiEbV009UmGdkHDrjXsEZvzIKmu8W+BMc9Hz7BQSwK
DtDXzhC54PK/2q/8WZjeaTE5FuGO8QOpUq+tTZOuEvA3AU7swPd0ROLd1YGgy56P
+nPkzI70IAP0Gv4t/GCSR2BWx+Auth9oZy7YNCc9m0sj54dAeriVZ8/1W2Zux9mo
4LGXoGIsBkeMwBjekeIFkr+DRDCOcVGlQkpmn4fMs6IaPzC11TGjthdLnb+PXcdS
cZgnut0iTmCvDCXzrjBRrplSEEY04+Zg8Xd1hMoFnG/Gry/qsGzsXLTDz1FzKbva
amgOk00Mn0SD7hR15y63B8x+/O2pVqlb02VQCR/zjSWbVXxN4oDeEpwOWJokVeWK
TE+vcztL5y5GlNa9Y4BM42Hj30k6UFOk3xW9FtUbm3R27nS1Q9NTmn/kgjXWOVc4
lkJtBDnL8WveoMtFcgYTR12GveWcgWeddB5k/Y39uDWLmUh7CeyZ0BJD3vHx6QD4
I94w75NivhIYKkJB18aU3SNVoptqvhOGHXGgik7l6nyIz2e9zTi3lcUbZMmfT1If
E++z3qrjxiaS3V8Pm52xb41i079mUeUAJ2q3JL2TG+LRgE7ZjZHEnwen34tCRuDe
8R46/5E9Hvf/L4qeheRtsIJIaJxl3n03WvxZ78PrN+satLVIDpFQJb9jfA3FV5BB
Ez3SCfp/dzBlUmlQB0RmvgYqRIuNPw1ioQfTp4oYBHeLtH/Qr7laVm/iEkZcMNRo
ywjf3rL58c8/b6bjtS6gI9d1XjxzZhTMyIQqFSt7OU3Cg4ayNd2bmIslsxajyui4
CsvB859reKEltiX9tNDfK5de8VQkIxK67E76JDPHIHeao8qFeqMewG3RJD6YWYNH
jT/8gb3xjIeQr1j4GBYCOFcOd+dePPEFlWVLD3XtPRliUg8+CSxuurbfvMi9SqZ0
quUlfgrXjQOp/5JRAVQ6OGctItDW/yp/N2Br50mno/l3m4rxejz+QlB6ZYE4CyYK
OFnfcUgtUrQHdTVyBSXISSVF7dGKH7hF9TIYO92YOP1UIqevc6CuvoHmjb2uoP5E
dEa2jppEJyljIoTRRuLQAT3hA6VQmHcRT0AsNhEWGbnwKWDy3Ixnj+Yo+CRQEurO
mWR0apwenRHwhThk7Rkl/tOTl9lsVGk7pdU41zEX/9h+d/GGZ7owfQd0qW/bs+cv
iKIRZFdlgXYJxgi3LtA3JHuemuW/c31cllznqZpMMtvui7eQ8/TdCFIpq2MzKzZk
GA6hnGQBceuYBfi1R8vwep3SUuLDIXaQoWbVgnMaAnzvTFh2RzxSUuCZEeoKsfxx
GRe4p+y5weVAcfsAiQa72gsuRV2Tx9a1qgmFc7XIB3sdmPoKk07vpNZXxTHqUEnD
qBkR34sS5CUqXK2TWtPsJ8OdQ/ZnJylt/j+4W1o0X87h/5s98Xu1MoSaB6sA7awy
RYIQR86rqQ0C1ZaEJi/JZv5xefBqSo9WXnYsNMgGTAfELgg7fO5rcAbKNRVi5Ibd
o7AL+ovDd331jXA5tHGYbejnKDCCr1VkKqw/QvqC1lPEtlr6a0PD9et0APLEzUx2
XMYOyXN2W6GrgGUi5Ae61KBEVLXriU7mc1fqf0Q1HT8zKQZpDrDuJxTQ/W2u8WQJ
QzaAA7YAypjOvo2hNZfEWtE5I8yId4++jOTQSn3sZDYvcdSkXLUmJmAyOBDgVR8A
eRv34klK/+dbWeU4vFSFR1nLt5UZ1H2+7owXRobLsnAHZN1xhJXb+s9WvxhHHxPH
lfotA92WXyBzlxGExG+vsfciclYyyA6RhOuDoqyi7g5gOCAm3JZDWacPlBnj8R/i
ECr4Y9kt5KUhfIOOt07Ov5UDEf/YFnPsqcYeBBqrQb5nkrL7VvWndgHo7gyZ0Ime
G1q/zDss3Vhme+0Bnhqmp71d7dyjFPaEZ33hMnEe8JHS9E6PtY52ucI22SZwY0Mt
/bf+ZkgklMC8bNU8dxPzB2euhD13zWtjr/+g2r8Ip3UPW2OBglNL6qeIZNuUQhY+
ol78kBs7CUhcTgddfjU+dvA+GrYAROxQbJFAzUB+XE4LlPJju1NumKgDgE690QAz
DRdeVUo9zDkfypNGWzkzRE637++rUPn7m2iPZWLUQ4KtPtD418oXF0+MEsS83jAu
sYYndTWsRGGEM1hDFYbdWhuzF7sZ2rnfb5ysmJVMgGlBitAIZjtQD+fxK7GeIT1I
s1SCfIp+WdqPAxUy9+6KRo4XQ7dB0PtuCkAIysHG4DgeggUzAYd3T9IRXBEfa29/
ZMzigcAFjs3ewG36BbN20dz0MEdAQP2NqS5XMrrnELBFodZ06ds23UnfYo4Twkhh
YhPAqjjiIbl4IfZ909YfcCTbR4DxMol+uDFFOR1jvlA6YfdxQg2VcTQPKdfFjGMe
HZRyTHc2g+3vTz0pOlw7IcvvHDNFNvf7QYv6dlvR2IJunTobfokBUOep1on3ud4h
jz+z24RSvK3RGbHj0FqzLT7zrdv6H5WarcvYirijcRZX4w0oAcHPZnYGEiSOJQQm
vkVoBKnPT9gbI3lCwrhHpSu+HqBRc1pt7A/235Ajl23jJWYUg7ZSIUfEvKJxuhKp
xAb8evJdLz6VsUKBmuT1r57Ft8kPmIp6pYVPlXkB1KTqGrQETkNKqZz3DaZF44XX
LzDjgrJJoxf6YF7F870XFzonOx1tRHDr0nE4bYHNm0j8LstuVx1xPfRhXSKfI8AG
YkRPhjUUis5aIR1AIzoMT+qrfW1op0wYoI/fOipV110MsXq86v6yUkzvhJgt/FU/
UEoKOVknFniWWA+xxmox51NFR6GxgAymxRQpc1tG2kwIONkh+ZSpVIvataqDBRj1
tgA0A0kcNJJ1WPO3Miz9Z4vqn2mENE9z1f+dSzwkDwzJBA+QNgqFVOhfmiCIFSCM
j7D6P+gbObCHOZAriKR7dXgi12k5P2sNBPsr2O47WlktpGb/WOKXp4b7WNdnEo9b
R+HKyT59/lMNHk5EzQC5oX3OV36iJUjhOv0e6RkzbzB69aRPTbk04fSrA+I/M4Wh
NyKNRu9VNqXdJRjmsmQH+SfEEy3K2gACgv0FfmBBdmG31llj2ka/QR9MGdFKCX4e
m3cXJ54K947ZIwZ6DPIza0RMRp/SqPjXbqoDpZusDuWD7vc40aFf/HzUzkEa5EZ8
O/vt/lcBnxTaK+dsdDXilC4uGoFqaGS0TZieJGFnc2aG0q6HVdFQmVAWSMUNhUoc
lGf7hFGEkCj5ZN7B7e2RPRQjsZ/5eZypSpUBdf9Ixyyh48ySo+duuYPnKb93I+Kh
jThBB0yTnupzoaEjdyOfKU6t2SX80FBXunr6utVjZlcQMmXktDhoKnGTUUk0xfw0
A4mizWu7j1/diuzY5Yz/csUmDRngnd9XL/aOrqjJPClvSxzCbvlTFjLWMkIVY8sv
ws7eVpG1syDFAPJ6TWXjOsJCI3q12uOTBej2wCm18Z6VRFO/pWByKk2W6OF4guRh
1ZHgfxErH1Nnb6MSZkLMB5tdCC2Ghi/4qteB3yUgQdFua1I+WCJgP3jjgZb5QDSl
TaJoKCVt55FHcIaBpxE6rvV7jRO3yhf4K9kYHQ7s9IhTDK72uKd06zNqmYl5tv4U
RbJ2/5nVzAuUlD1TJjJoXV5HYGBWbnmexeNVkC6tdF55EzUDJuODB0il/3GyQQAk
ZSMwzU3o4+EJRlhLb09a65RZ7fZ1WzAOrkj5Jzc1RSfsiGzCabe4GgKpjUtfuw23
+O/vto+Up7hpkzmoH3I8eWXiAaN62dVHYJUH5TYtW8egyQJ86WTx/Hv/pULeU1dF
GhNGly+PgNpr08FdeMgHlKCVQuLIsOX11kZR2MekecN2lORbo3MArIBdeV0BbHPi
FOjOWAXm6CDCpn8vj75K3d6bUXVxTmpNwuA5Du+NXFC4o9pfTesGIokUpBiSCu0W
+3u5z7pTCawB6MlZgJVCjtU0HpFekyNgomYe7LDW0ouDGBY45rIPjAPksLfhLnXB
d+zQ8WA7/0fvMc1JGA4ixbKkgRySQ6VInZhP+G0GLv8qujfujssV6iuoZ5AFn5VL
vlcx85uwXQ6sHsy/bdzZdVr+Tv6ymWh1fhk+/A47jScNMzdVu+xfs40cIUJPxMjI
m5hZe2YJ2909DAyTkqmMl1roQQWMBCFqbc++hV4nxLF8sjww0/51PxawHFPjpRJj
XjafcwibF63w52NrYGXUJYZn179el7xljZWqzOyy8ynQsGMfPy7pfnPtkVr+J0+g
5Q2Jv6ZXm1hnTakcIlfg669EKzpmNNR2ZX1VUsNeKkppsAg7H35PWjdgNDDooTbx
ACI8ESYeQBiaN52MDTec7tKfKhODJ1adDa9CiKBECkF5B5t/HDDa12ylvxHfOQzS
AHhwSb6EgfKrY2+iq7bddIXoqFBkHEAFNmDazyV+UfYVYrOZPMfET/AnIVMnTi4O
/mfqjyTa/g/7VfE/U40LTYTVf7fFMm7ZuX7c4bZuMORpYIj+DiKEpUcNJfkxMrko
Ttyac7OZEjDVCW6Uqs7KxjV87fqNYkSVtj/66vUWFalDSnrNvB3gl4sTndcsmTk+
n4bC3cYscutJRwKk4hL7V4AZ+JBp4Vuh7T9W9rPbd5xtHMlfcEjeWAmLF9w22cCN
47PSw5hHrgcrtQu+y+qFzKg2GWU31FP5mToN7MWYI+emtpjjH13kh/AwJIXvNYWZ
7xB8MMEyFxu1RuPV4Fs9TY6sICCP24UyDOUGL9ElgbFMToHsDpBiMEzddCYbnD1M
4nVUem65/rzZrulxKNhkbweimV/W1/F8dDq5N8AJ1I+f+aAahltZdGCFo2gFIoxZ
CbA0OaPUrm3KUpgMQgs10+QzvSPne2Qsey3/XSE/VZegogzYptaCmMgiV7LD/lzW
fEJMCE+vUEf4IHdPkmT2/gAwmsiJx8FtbNy9tYdKz+jTNONN5rUsL3UccWo5uwCw
1dh1OpJKSTO8lgjosirVzQPoN/oIsb59/SWSRvqsRJd+m8UhY3BkCqbyK/+v3Igy
FeOfqemK8u0H9UIL+SD0LZOwxX4csNltc4tKuXWcXna5/xsZIaIzzRLYLjEnkvXQ
5kWsHcmGbqxGkoeRl1s6XzDWGMol2on9KohMT/NSCF2XPqYy7ScqyJwjOKqs3WcQ
1Aibls0DdRWZse2OjO3smaaeodoiZ0Mf/SOuRxHymFydNsP9HuXP40YBfe+wI5/9
kfba1xVmdORO5aCzNGdOVGFx+kQ/rJT7/oKzmPq96tEnrIvZwx/hRv3krhQjKLlC
d7OIRdVAl3qV67dBwkRROw85YnY6OYRscwe4SEhy3e+KtWaad8uchOzYy9AK9ssu
wkdbjfOk+MV7yzb4Thpm9jEj7vHIlfjGj8O01og81iJox8pYiI2natY1noOLYbnJ
67Fqb249mOCVIO6CX8l4K4bliElte104QG3cHstfPoXdBvibtdxs8bkKB7Wzua3p
exJ8Qy5p4bIbJZNvGQ2LIHnBkTldW7fZM01DrfSc70X1dXs3gcQtWcr4TQtvimTh
oWYK/EE1rqJePs1hrLYe5ZTtWITSP3eFTyOuPtcpQVWaSM5IdV2Y21oR36k+/a6S
F1htbdTW7EwJW4WHZvjlIWhjoVM3ga6sNHo8hwq9xdfE7/9RO0QssLmP2OatFSU3
QUapwMkUZfYs6T3XJYdtqs91n6j/Qo/UIy05yiqFWH+PmmNekvqdILsCzdXUkusy
oL5rGzeNABv4iRab8FXg3c+wn15eDs75EYH2AMWJ4yf+hnEb+2I7ljuCCpTtTS5b
W2j5XF+217yQdLatqF7iQOofHqiXkLLjqB2YDe7brz5Z5EWygwPRlk0aHGxPfAyE
V71pHTIfvwvqy8a6tZOwcfP92IbXdX6dDz3xGYPE5xtjvmeb+cEYAnswusVZfE7Z
Hf2Tvr7d08l9OTAVGord8dWhpFue4GXWWdB37rxGhJzlIPIXaTyf8wXdvSxX6Vhu
SigD/WmPyTKZMzGDf+se+O2IcOnM1KoY4hPwKquux6bIsnsOF1R9v5s+J/Pa51su
tlpJX/OUvyUYD6lZYfzI8PtA9kLxyqANXNuW6vcwwh3XQlePeXeu1bGvYRDSpVuz
5SWodjh5qMuWQJfWu3+YOtUnnlDpgQjfKvDxRC7zBAv6B5Hy6/gL9sFeEic/Gtfb
4cqIFkRf7+JpOiumA4YgbtSd0eu7TH/Vz/gOEuhKt61O5FY2ZH1jox6rihelLN4C
hMKJwLU9n5ffczeDjPeBPc0aYiCuoH0gk0nBHcVjZPbiIPNagZFYKf6Jua7eJ6i+
PDQsB4c+R8E8A6IWULot1JqfFki65vRCRR1deJJ7C+Kdh5MXGRw7ht/j/gsWMwv4
WELWyA2RhQNKXL1LwH+W3xEO6/BaAeCmZCDjUMQprljwqCK6SOaNtQYfojQlgKBs
rk9sOyppYupz8GupUto4Fx6D11yW4QR/rorp3nFVxcoZuZznoIX2mEXZoeonFqSK
W3Tgwrn42HMhF8mQZDNc7QW8ZSfbR7gd5v//XF4CY5aXyEQrzPspZVmJaITeL0/q
xrVk6EW5DXMkP5IMGBckH5IggeDcHu0U2Mn60BOyuYJxXFMhIcMza5E/a3e8Ye/u
nzRJG9fbnzQyQsgURJwI5t0ATGaeZoWiaP2hF7uFUPjzxtL8ev7YH3Yda/PEDLxz
IAoaIAfboNh5TizNtyWKPUHMA/5szNMfGn1crHIAFFE6UML9P4IoMgGZRNrBDVkX
Uqpy8PSELXSTDArewcyYV1R9cU6Eg1biJmTAleQKzysAVMj8rduC76k8COgvnGQA
4/6yu6XcexZEqjZ3yPtmd6tZ53MCGm/E18FuSBN9EeqV+8ljadc3k1TrihFI3G68
ENovFGhKmDrKpxVOYFPQk61XSkn7+HkeIIRz6RWkzVAdIZxvNVvgQnhRPHIkgrrJ
KdbDG0PvVAvV3oBTKkaUrJW7xkecMUHr22rnwtxGDKz14ErnchARlkMXIoLpODjP
J4CXhS66EzWH06OjgK3i8iYjVBc+LguKkh/0j1Wm5JzsBhyHImfd4WW3d5JJ0NdV
OaPXJNXHk6VxC03HrKg5CEIgd/NpUvnXedEwzKtm2FmzSmz0ZZGpwn76zdOaKbVf
GumRbGzKQ9QL9DGuaFXExKn28xNmqFxN9UpY2n3yiuN5TrcpjDZAX33u/YcSzHMN
OeuX9mL36kjjMtWV2w6iNYQPO2rFyxAkP7X94xzfdeynJpWGbLkCjHo8uzsk8y4M
qk0IfpURac/eg21id0Ht6sVI1Vvkn+sDx8WMc4cPIdlCjEgHW5GQkDpChF+T2LnK
rBg27to3GUXxSiB7asU1g/KHm/xxYD4TQ5+FVTvxV5dJnStxAl1A/zdJMD5C6qfq
psv0yWKvIWQMkv0zBrk/L+aimfWSAj7m3WqI3jKn/bf+DUOuv+odFwoKJEnyw+bk
DHH+2BOCIJ1q/G6kpkYCXf7vNRlLg1BZYajjJP3PFZY0yoCUUP4hZtTQr+eSB6FO
k00OrjJvtJ/lTxKOSh0/V6pb5a/eQzJa73a5ggGke9yP67V+9pIqIk1fNuRmB8r7
pwtCP8swrmKDCcOJCcb4DVdk2Jy7WV1hNH4bTC0Y7YGsKKQvdPLp1ghMWZ6LSeTI
Skjue4cI7hphO89SUAZXrhujZYKXsr0wZswqdSzFatiYXo1QuTmwRIN8HKmWa2/q
k1JbRZxQBFTCeSz/HdodAcvrc9NxKrRQoLBWeC8lmEaPnC+lNECXzQqM0hZySywH
hMZQS/RxM1/+n380mmdxDujohump5W6kGuDTwYwZlh3qL0zhWjpJQqjsteoU180p
TTzPLU9i1LMO00CirZABOruutQp8Q49pkQihywEGt87PY2kBesP9hGsJLvxfJMAe
xiGrWGPe31kEzsQPMFPlJkjhjo1QvX7+dJGarUjmOfD/Jp+W3xjuf6/BDOE6QbQQ
ovTFSOTx7kTD8i7ePkOc/HnRitRI4l+bDXs2WfBMS9GWjjJIi75jycuAPFt7wpw+
0bVJJ3RU74Lhx+m2WTmI35jNJT/BDCO9mvbcHm1B+sJP+wtPV1PFDHGIO+Hq0l9K
lY0V1kmbIDBHEJwzsNVlQe+3pkegh/4BaqtlwyUAxNSkTg3cMfDMNfgmmmF3Ktam
50v6n5XrCDdSD1wVgPi0B/LRAtAbMg2xzAOh0Dh2n0yZ102CS2euyL67vP3w0kJt
ROHk6t7XpJFsrDA8jWyK1mKG9JJTZL2p+eEuv+wILYUXqiyAVQz0ZaB+4lzUwqOi
8hXA4hnRGKg384/3TtWLecwGiUNuZLF2JZwDEqGQtNkii96Ap4AZRFnxt/CjJYnz
9bDrh1beP/RvfmSgS14rpd4L0jEb2F2GQIiiQfUEmoR6o2Ihgp6FYT9SGu/VQrFd
oXtttpVumV2NSCNpMeD4t1My/X/QVFlg58xQ01Vm2f0dFSBEJGYkruC5INT25+Lk
jq2rW0QkyPsO3HmxQm/BYbOlEpjMCm+C/Cxhn+lKjmFeBxSQseAaf3nAzS7YPkRA
NEtfOOnTpl8IwNMQ7X03mmylAalZcn9a1hdUj+C93lA7NkwCRfqrkfsS7vu3DbBo
z2u+Kppw5psoMsWIOLI2rZ0d3yive7WH5Nbr8V4Wupk8dD7RCe6eur7SfBcAsV7V
kgAD5mJ90XP2FJCpmnNZdk1ar5EwYKOOKJfQTpjcSYKDLs0GNh7/BPxY4xcnL+4h
QW8Py9mhJdJOjjq2QlMVGJb+AgdM2DDKCwgCQiHQzscfW3OERQL8t+89yDM1visX
kiQojA7OTzPfZt2kskvQCAYDdlDnZGRW5r9brINyTv1q6aVW5fG/tUscWCfJTIie
b5AHgOLq8Xgfm0UCrePaPuubnbdS/5E1IBNKxE+EkaL7QNaqXg600XYylZqT83gW
ChpyHNntgZI6XqZmM84hJnhI5fJ+0SOtbokacDAPdh/wxo3uB86LsWZOA7nqL3dN
iyG6FHr+BWokoSM0tJQslw43oFgUHV97+R7mqboA7liXAjbWNlkxMBYreZK+ZdmP
UkWn/sNeno72X7owa3xajwCc2BQLS3N21DdsZ064un36vCQrI1ew/gOeroVizRug
rDpoAibNLMUjeltcaNfDpwjq6VJLNsCmJejGj55N+NLaXsUG4ryKRlQSG7lb+IIs
fEt1Qunj65wXfgx+iFLLoirlzwuv0uH30hiaZVQ0JNq38NVGOXYhjtRGUq0vL4iS
H9+tLX+HPR3JLp8hFl344+pDJQ8heCuRUMArJaQUG05I8KuYJrpPtl5l6Qle/YiX
lxI0piQMWLtnL/Ztqv1gkO6hgia5Hid+sObhg5P8F+u7bxTflC+J2eMsDZ8DK+Qg
ryuMlB0eCqFVQdmHz5LusnFx5E93dd1IUkrRNHtSuOSZFMxMBzjUlyPU+UB5SqCD
7KF3ZAOaKfiaDVHZI3XRVq/FLCW7VlrJMzSyRFKIogE6XILaqfvKLGoPe9x2WCUW
A/sj1y9PCLKmWO9PF8n2RndLBDCNwKMbpA6M/S+Q2COtKJMK+xgc0xkPcX4hcnxw
cQOu6ljCYA+tBEe/eRqsMgAdLNVERqgn1q+8IZk0JQJLUNB0p+knETnucc6Dygwt
fmJw0uLz/NYsHcs0YrbqYF0PNWkxuCnqLdEQTUDtoY7U4tuZYRw3CBlkez0aZIa6
OjoqaF93/6tXDGY74u2Q9cVVv90AJW5XLBMJWK/BGuzuUX4AhayJMLUcHUCIWRSU
96cZ6L+raRY4sl8QC2Qvbq2w+FLARTISLuZPX+luOQmiSRbyy6iDkoJAbe7Kn+j5
pM8rlHVsv1r3uc6YvnQmoHcyH1ebkrBqJUq70Z+z8fi4v6SJbURQeAX8IAFQ3Gfv
6YUgxQAB331q9iIWixK+/iHACR0+m8bP78jHsgtejgfKEoQ8D3z+oOUcIJpqzs3/
UfLKc/pTwDFQq/nykodzUgo/mjSiWpUXY4QOdwVvj6f7XFzRVHX099E+/ogpLjkC
W0uvakCn2so2xUoexp+ea0gcyChs3hvh3w2HNbbKc/+Yn9rqKF9aIrpgClNBeiQd
yffiAThVDtoeDVRYfmxxolrF3y16uFRiHz8xUUMKN2Fas1W8Qz8EvIuc/QnYCRIH
yXSRwMeAcrdDJvoYGRfHlU764XivS9gqLUbFrvEHtytNg9Bg1mgFARR0O6M80t3I
XJFTnbznfF5Gnm9umHJ/qNvoNpsI1/abKb/vmFA9p7RihbZbMrRkhBpLC6GTf6gc
NcnJTHAubEYvr0sszTTMyjnNOt3EjsBKEcvbBtm4xItvkZoAMVPUHy8b4SkQFD8Y
Ulh0yQFn8Jg6j2DLI7L2a6FAmrf0Nq8ASRZyuil7dwmcHdcl5FDwCZLriFB3JhrU
lPPXEo+WvEMbR+aqqr5C5U/tiQv/NL+hArrecA+ss/6gtzv9KL8xLi64LXjiTeFH
DKPzE81uUTMi1GgAVDyb9ywQaaiEOGXptjzkskO21JyNECPPxSR68ud6/kEvcRhS
T2oZaLM3JxCPlj0ZAdcdPnc8ZwWTUomotnkXoryJhk7WT4u/CluIq5QEboUJ3pMc
vM7HoFIp0TYm+gj9zwlr6mrB7gj+BR65EEYcWGi0ZfELtSKsSmml1TeSEN5apbpo
6jCuHMsDDS8+v5BvQ81Dvl2wvnzUtcXOCLm0DDS9lz4/QaK/G5I3dMM+KIstha9j
TCyHtyou490dbTf42KMUj0kYdP8xsG3SZHglIW7QsMHTl6M+SPOmbSWhnv+siaFO
bkkxH4AqTJKUun8JfHd6snVrJ8Jn9ie9c5gQxiPkdInUtHvdNLsAqd+dTAAC1PjO
Qsj3w5CkE44eDvtUcJIL0JM1TgGUFiAOKMswdB6+msSaazqZ1I1bpshfq74PiEX9
B3hDWfXdcM4jL+xElqLrNLIs5zEVWngux9GjJWnnZZHsbwWQVPA0xkdOWpuUtPna
VlOG/Fqw8E2Qlo1XHW//fPMO+z8FneUtSToOgAHMTZy9z5cfgolAxmWaKoj3UcKi
Hxhvt1bzf1C/EoQKNHRZAgzoshPjxwohwHX7daFYYOjnv37CgC95ERAnVmKl6sfk
SsyWZ4TI4BfGxdNPusWwhDPhop4xuoDtyzAppBxLCe7G2mt6jFu945HuU57urWwU
CIZ/pHCIhlqJenDngMI8dh9FtQFZjvwh9YSYDW6Aq6Sx8CU/mR8XUizUeTjYmuYc
9yQWxQ0+vbSmNXmzCh+8JdCsTg1uV/xzexBQWywoQ32JXivvX1EMk/E2DDPHKdzQ
haJH3sh1Zd8sUhlXv6UdwGFJXpdVsULi5cmmIWJs1ND0318k09F3fWeftCXwKhMx
h4loF/ed0m8AXAQKeUleYLA5eYQCuc8fUnahMIadv4tLNs8w+2x7x5wkotYN55Ik
pzzx0CXsChC/PWucNlJ2xQeSNOZQKcoyQ5WsdU4//I+Gets50KplGM0XcSK5RkL7
cfUDQfq84+jNp56YJ9GtE38uNpksAHtyDN8EJDtjUL3XWi/XfXcKdEfUynQ/kwYP
uO+LvT2A4qfjP+nsG+3XY7pmp0f821lJ+xthvIJOiUC+w5Y/bfGGALIcfjvOa9a4
WR1EB6XNoNmgmmUMD7M8/hmCnAfdRXbHoniheL7RIBF/vJXwjk3ViC+8O8DFXCM8
qOkrvUcCb4VrSMBR9p8n1JUhW5H/NqDGDUEFdGA1izRnkoCfd+Ct7/v+f5Yl05n/
Bkk4JY56DenrmeUh05z5LUUV0xytyXE5HCplCje1KJG2kVDCI9MbGy3CHrAOvaUY
JUqIQvKd0P/siKb8tC7e7vAiKv8P5xr69jFIDX6lY3SdX5Dcowooj/8nvTlV13AD
v6AGz8ulnGAVlYyz7LXmtgrnVcF6bvihkkKU6ytu4ajI9wK0/VphVHznQTd8kHlQ
v+vZo0KhE1MSJ8BGqxdjqdKb7T+HP0khiVdGQWlxC+mK6e1LhoEzXfUu/lf2jLTw
HLn4q5zg2iGNEtvHbJNzjsRzov+DHMxZDninxpf6bd4oVJ+Qk3oZUMhiHFKS7ojb
gM4IKWiau+0sN8a5B57qhhIFWCVCEgIojjLFdRgq5/d+EmeswoWBGvH5GDJameIG
G1Vl4Dqe8RW5zM3OVvDtjQbsuPdVg98ULg3XoQGDBrqILe2qRmM94Mnhw6eLaNQo
BbmPpo/1B2NEyCku4IK4wgbtRPleAUavxtEgSNyUUKAD9sbgd8xfO2TKymrRcseK
VMLHj2/zBX/X4NKDM80D2T4kF0mdo193p8xJvdtqYnEeJEGDEjqv19eLDumpmdC5
5OhaHXi2Rtfw3Va3QmrsvPJvfLWFTqgU/XYEPP0AqzPy4d9SoilZqH7qUA+BOIjV
3J9rwKLyQZCEnwqx2dBi5OyS6B4Xg53u9iVvmtnVv4F6ZeEQFZMKG/PELBsUrSa4
61wFyuadL+RXd86Shz0DrfEwrZFd3H5IFr/G0EpgPMQTKJNXXCehFwM5T6wfUod+
rWZ+GFXhCD6z67VDKs4o49ZH4U/9xiE+b5Ha17QSIAurutRdnnSjIvCwikYLv+dV
MQGEU8vXOHPQXbIiXEYn24YZ/tJhhJnG5moHNo/equ7EYI+mTHsP+WyH75Jbf6+3
29TjNcAc+9Fn7cFZ2csRoS0ZivgrXFWuORQ19L8yHCIPKCBv2F8Snm3zMXehOUJ0
uACSBfk9LbCtueFm6u1nXPZ+6JLsRDeFeLrF7AKL01Vt9RY5aHWKRfte9a3iNZVj
eTu/zZ4A+LaevR8SZ3PzfWeHmfr0yIdFRjvA3rjYHyGo90ic7hp4iQxnXD0iCzlo
6OIlPpvGNJAqJn9na5PDJS11tvtI4OGjCcbuonhwWigu2XTiJi+oju8LT8Ne0CJE
G0+SZdzvvwdqhfN50ZaDnsH8rSy1AQZnvwmQBwLGZ76rowC7EAct/+v2Rzl5dlvV
6J/iQY3drpfx8OGXPxSmC5pxVrgx9TlFbBZf4RGbc+PhV8zZjrsR6gMqvc4mz/Vv
LQH/AO3VYAJvUSMD5AQ1CWPWC8ckrbtnWeQsEbIujOrfnrxBENKmNIz3Kq8Pi2ET
sRUsgA84gyfPDMmgl6LfKRsW4IQXg3iaX4Zt1QPggfQRdO77O7vBub8Wj/D/X/c8
RrYDClKFGKdlOmUvAEEUe3STIR5TBpD3b+MyWVBkqw6vyNetSsGKF8bTY/U+pvyp
qBw75DrXjXTsjI6Zdx6TowjzcEMiWNbNJjzY5b3DGPrTyWzCPFUmNuApBA3j/o4z
D810NMRZngdcts0hfQUGMt1jkaDSyZ55nEDB6g0XlHZAPsSgDQB/CdOuCYl1IrLP
VAgKSJT8PZJDycGSi57YEMC97TzrI1IUsEzt0uDoEe9wSdUseeVmTo4mwhriDa4H
xp5fYLaG/lo/V1SEWreXcQ/pjk2m1QY19Cl4HXhpR70KMMjLOVsYa+ggGgba6e2u
x7XwfIoSuTWli0/Ir/bAviNWrwqqVuL132tGclxH3VIDLXvXnzkmP/n0VlwMxnv2
hz/OdfBWh/FS14Z/sC+ODcRSw48fbYN0Mi7fSavB0padNvJNtxZ1lgPeQhZwkQpK
1Fzjk6L6tYVih1aeim6sD3Mo2u+sKh5dabuGPbVkYW7XttN6tLeADxh4aGTvXj46
1nOqtjfSQrylxZco5IdgQM6JjqEpQGfkujLDJFpofbCHXh7NyG72nUpkhFd3JTvS
0zz1CKb9gLHYuLrxfVPY8TFuPMaTqZ31EqxT1qbafXMNiQJicbvw/+dWtibinyqm
YQuJWhPYMzN+7Av5ILtCePNz2iOi0n67xmCW+3IuxC9pewrgQvqkbgKJ7H2YlE6P
G5rTXIUv2l8XPghm+7Fgu0qS0dFuHNjUFUNVQGRdTihEE2ga4mgUJQb/q55O+CC7
h0OEqtjT7CnxGHo+feVnEQwHxNRr5ROPZYsX+OM31P4STrFex9AbcSLBFQ5Dgz9T
M+lroMVG/MXBPyS8bzHhVGtOBR+fhcJQzz/g2v2jzZ+SwYmKdw+rEzwoQshoX2jZ
YJj4YR9h7Tf4kIAHuzHGJRD3E3Q5p/fqOxpFEsXZ/dmtKRnWDmfI1nZNhhUcjMFa
JxZ7MUqSNRcX3bBUuVTHhWvWgJvHmcfnevpXennymOaD24NG9zGmlXoS3/XFAs7F
fIs1hgxcItM4wiOPMUMQhPEVAOK7hTvMG7J+zxrHty6q2rmf/4t0K6hiB1BHf+iG
gqa3plEt1zlC+yMTOns/VE0AHb7lKB0+ojjdj5V6iXzFzX07wKbwy1w434/FctGz
C+U8N86wE/JIWoC7Mwpz1ETlpE9qo6wE3CNYl7PepKFbbw4mXAphENByPklnIEza
WCA7pwAYfR8LkgPHDvTymCMZgnVOo4MCaMHnhK4WC64PrjlP/W73IgnNBNjA150s
8Rzl2aA3h61wQ+10ocCP/XDpAT/jNaGROnlQKpR9+CqFhNkRrNhYEhX1vPUfEIHX
O8JIkTeeprqL47zUE5emm1jF6IV/4MrVYxCdf6PwKL/dHC8XFFgY7IBJ4mMXVi97
OygW0UEputm+OwWxwL0Hb1nJX9/R5S0K8kfrQoi8RjjHdqkECcpGdbinhNYw/e3i
g7dy/75tvoQkClZBg2zWKhckZ9D6fqlFkpxjo5jfb2Zw3bCwJoMlK8ZiwLm5q4bN
FaiK9hQggxqmHe1ZlyqXha8u3wPdBrvNGWUjqnTJ7g+Qwsz5h0k3ws7PD5tz6udO
gMPjwpClHjvsxhBQw/dQtYj0RosyEcwhC/dFqCytdMByWe3d1ju9G9DQqu2QdR5o
sDnPZCufUpBKW5tk/TViq70mJDqIzYYhDKK8pvg2i2V9+Bqpl+/EMAUhH36Xru+N
ArxcesqNBN7wkZIXw+cqYLdwdJEZRyIrtnQYdrDjPtOIXeToYxIQttzwI2NLMhKq
dblq+7OKIhKrPwaK3RanVsETFhOyodvLtQM2Tt5P++7cMqK5VL8er+pmsnqDeRht
ppdB9E+3UjEmI5vjqZoayJVT+WC5LnVYGH4LqaNau5wSQJ5h0EZzgax5mHww3a+j
7AaoXBQzDyFQvzKaMDVmYLNH/ztyPy8xrgjzRfrMYWmlAMVyUItT+Wp/251A/Bkf
r3Koe+l9eo9bXRSNIJf5yF6Ru2qUz5scVzrSUR9RoTI0/zzIM39AfWefyBXIC06B
ER6/lGw9n2EIAw/3VFQ19UnFv2bcIW+zQwydOPE+tHnsvFz2YEl+flAzZYUjST67
RRh3Xz7didaw82OGAna5MFdnXJZ7TfGoZbV7GMO/Pt7iruKo+AbYq+ijZMRk5Rwi
t/KPTAbiMcz+6htzOZoWqVB5zu//R7zx7lEGs3mbd3xTHQO6lout4sUsm9L+6zdZ
Ks7UT8dzQ71MCVICBO/EFGhTWU01Zk9M+sNXngt6F8fkKdf7Wc1eL2+2dHKjFVlW
2nt+E6wM70cXwubiIObwSp2FC59P3lWiZLNEN7pBkxQeKABZxfnLAMQ2IrjSgFZh
rXrGIMMBcxDQgg6yZbHcAeYl/efggy9ESfOoN/VmvU0tGGNcLExbzTeInxwOVPvt
wSti5Ykv86ScBX+tQ5g+2oUzqPDc6LRjTdAyFS05ntBAtH5qYiYt7iv+YSc5IUgW
s25yy4wFuTSpHnawQWLsNbWQXFJm8xsIxL7Omtk1NCxSEXLojVHWr6pSvyrfKFOH
0y8J9AiODvuKwIBAeATZJ/hnZLWPLq+9Q60gkfyRdvR5TaKetMNIlhwFuZIGwVRH
GnsMJtHXQGKpppR1G5VU0lCCZkfnzQ305Ch5uf9OrRiNkllHa6CjSFCWrJTCTGCG
I8T74GSJBmD+7O09oqPYct4tPH1u5s+Y3r/KcowOsRd31xRdDvzJ/P5fOccybwuO
BZnOYqfNNVEjj0PxElyz+8SPFIRuPk/Amsn4YTuaQ6VNPSB/QD5ufqIyaTWGT3Iw
T8gI/VXaFHtA0Ysmb3QtHSJsZbt0sGUrTIXN01x0cjEY4d2M+JCgjykmLLUI5RTl
YzLlzQa+7LgGYjCIZudRn14i7IT2y802NwmJUXVMUsPRtAHoPX4SSpGrjU6NyNWq
4KZp+9TTMGBVOKpqqLD4CMKD+7d3kT3hcINi8xkDwPL6jGgliT+h/7Njd9nM1i4y
JwaeaHXckj9e2G4/H8uAqpAIDe2BwPVSJs1pR6h9a3tDmJKtlWfl4g/pCjglzS+w
yRi2w5N093AYfJHMAWtOlqqrAx9JMa/cCi991QjOmJgbRMli1lD0CerulvK9dDgU
2eJ7cEU+sT62BYv5DjEpbS2SK9EIMxFqG0lovxdv/dFRSaUgS8cdCFQtynG1WMCj
H3QhJeb5040fCZevbtYIoNBe1dDbJZkLSgKAhK+eTh/MvxIMJ1wxmrfnxL3wd49C
BnmjMubqvdto+DVYf6BGK6/ENJOm5hs0aLDZH7tt3a18riBFRnqzd/iNwYyh36tl
v/nOzgI1I//0QByspODYwwgNaolzfUW8dhkCxz7HzU5N7fhuyHbjIevvBteWtnJl
6FdaYCR67TYbBuBpmVsKPd/FaNCireCs+c6qtjzWnSve775LFutYlM/oSYhHbvFQ
dELUzfdK/tyZkG3zFLHdnTzrBMk09BtZyIQTfGtlz6Ajf7zsB5/lLzPOz2UB5057
Y6MxoirHSRDUldCp0hgEBjunk9fbkoKGPvBrq6WonEUNtsUUzrhR5tnrbF1xkAzX
UlT2WWtbVJhqCWb/JxlGMxce1yt/au65MhpOQOGkyL3UF+3Hgm1Nv23m+11JrlKp
Jdl6Q0L7lR5+iYxeUyEzjGEJRd79HqOj3U0YLPpehvCwdG1GE0O89AjZD9RgKTIG
wfeEMDmZPsOiGnOUcnjQgqkbcgx4SmIhb4p9fHacO8AvIef6TYT9ek0seQtRVGor
CcbDcrra4BAJ7diTuSYgpWmys6xKjyc0puLfYjD+hM077MRPPc/ge6ILAvAkc7/d
LD1vq+CYgl+CiHBfoyEJG3Kv1WUcAI4tu/G8zc3KAc38+sb03CB6qs9Wn4S6XVay
FLeQEnEqgCgZcE5WpBJrdHMWWlnze8LN+MRJCJSgoRXSZ0g1jigv3k9N2FEvUyPk
diPPlwTMQ7oS1bVFPT0Jee4TZ0uwvk2+hWH4+evvwnaNNFgStxiyl4RGl/Ea0KuB
/Bs64Aw3izejimsiSGWKNsUwUpQ6JLvtilOA8W/0ZMNLEwTUKVcB7mSdFCrxJika
scULPYOrZX/iaN9UnP7neokuN//ur3+6Ic6CyRg4INR8dXA33KmSdRhx2+PhSUWm
X45PWIR5dzEQ/O6lndNBbSW8QMbft1VnbRZLGP8gNLnA5pvDg5+l6hRPcOfe+fW4
qSPKIqIFnqDtPqnhKcZAwLkRQCwHrUtqsHS+g+vAfhAnYJR/IAhP3G97S2OXfxvX
rc5B4U+q7v50ysu4gEDOGAuOoyIF8SD7h0EjOgZVlga8z/5iXzf4c339CUHkSXwq
8ARSNEHPsWr5Fjy7hGcFFr/s1mRfK4kDWdzpp5m1tGlgu7pGT4aiV1NlqdmYHJtZ
ZT025TNisciNVdVmxoG+M+AFAgKZLkWENpI8zCcjBS8omlLhL3X32/OHkrGAud2u
oZyflXR6QU34ePCmRMtqunu6mvhkggN0/cN+WZMeMwL5wEF4+9mYf1W4c8rnuKhk
eqd4zUn8ZUgK7Yw2hKfpIsUGO8JH1Al+gKPDZ+lq1g02qJYrfspjoJgSag0tMzUr
aYybhk36bOia9K8p6Oi2jl4i+HdAx2S4OCG88ybwURH1SFP5bmLWM8k5lkvYGVK4
G8OVkhl56o7+lmdvGeifEqjxMnvDCbMMWmEMjrPdWQ34PaaAvfCK3zwK6XO8dKIO
BE9++5Ojv2x9HZfKFUdCFWU5ErO4HVt3ndfdbMGMVPqRL0dkBwYFso4YkbocEBU0
EX37YGpEwByLRo1/9KwbWErGeI1Amz/RsbmCeAb3igzKP+6byJfh8/SytwJCwg0B
PGK1XbpDlaUMeIh2nwRsydLEo+CY9EkDdhWUs0/y4TMdvFqqj1m6NlroWAi/xWdI
lGGjnU3o3Js0DjN5grjd07uKbyQqiMIYgWsZKuDLF3VKS3LogsZW+BezQrXpltUO
U9hz0C/JSZEEZhCJGZ5zEI/q7PluJGUwxAUqElvcAsA9k0VCDgyZYDOiYaiRECxm
wDAfp0VTSC2aKNoPDDGagd8bFxB1saoIZ4LsT0VHtnXQ3F9MDg7vQ9kiaLBwBvIs
l/zLYQNvPLxsKflntJkBYAgnyAxons1sHBxY46MF6CjhHITw1kePOwJzkQrm2ZDC
dlMgDZFZMVRl4g3NOovWZzArpdK1dY7U+pRwKAchf5MA244Yp60ieTtyX5wwgRbG
UZx0bveZySrL80oqNI2KO4vDuu+2suT+Km9+gb9nlh0EzqJeCMXN3ZIQsCK0fC3I
8cDUbs4qRfvW32gQJbP8H96ScyQe5HLdhr1ps5M2iEFty0/fg2HcvFZht/HQP9cI
RHXiGrFktUrOByUAmhPCAv74gWPNDbEauHqk9734n03J+SLKa4oNf6cP8jJUizMr
LtDPS2hNBlM8Vh+Znwv3pMJMyWn5suZ4H02qOQBgUZf0yNHAHxJ+LLgimVgFZw9f
GeEGEzcpfCv3o/z8JKNEjIaZEXZCRLGys4LLEAMBCVpbxaOMk2bnNUhhbmstD9BD
FNJG745Tvs9iE+0PJIa91UJ3E8vtM5WPLY4VTqcgLpph8HjflnNOqTgGxC741+Ta
3OijroCTW5EKW9rVqv0czGcVjWSetbuAC30fL5Dg0+7GfmO+B9AkDk+TBsbOlvMw
FhLY1yzmqQcpHg/eMNKcPvtqTbNrgbUZWuVUxjfeUO6Xg7ddOnIYOhr7qtwCDGCR
nYh7kbsbhpDxMCEgvZRhAZowWoqq9zM2cEpRyKdNQdMR1sfIOW+YR76rrYBXmEDx
YQZlw7ktdfHBnGyh3dV+5j1jziLWYRbNQJyldJzC5Nlp8cGsEAAu8F5KhC8Hbtk5
EcxzpWcA9Kj65artNSdDZrPobic05qigqEhFTcmGlpzgAZYkXL3n9tNS50gMfYe/
mrXCrydGNEaannWBXhvUfVhoAgdLV86wylwtrrTMKq5GoCEEx5FBMpszmtjsHrA1
BoAZSpE2/woJk6PDVXTq2xrIn3lRFaE7/wTntUtazdQ7DVB9ORByN7mP6whTsaug
Z86hhspju0mB7EUuu4WeEcJh0LybFSih41Q+GOXegi6J7uLgoUDEyVPFy9G7RSgO
tFYRyIu+ADuuQiJHPBt372X+bFyuZsTEpuG5Eb1giBJfNe8nCA7ZKpB/rGqT1BqL
oNQKLGRxl8Y5LIcq9khwag25/Yz4w6eCYdukHUE/dwf6h3YItz4a1CGwq3Vfpneh
U8V3v8V9QstoQoeoffXksiavL4UQsjQUIZ/CRGqCi71UjTPHipkI6+kRfBpxglVr
gFr+CLFIibcY3t0ZELKSabIe62er1kA+DLxOdcwue5/nVU19TyfMyZlkiRuVr+lx
/KUv3s524MtgVQHz2hadPn7KAYAw4DSK0Sto7jkuPb8kk/m0N1moRA2pwFRyUpR4
tTxi4Q9w0nvxuCIR+R48MLgZcdGH4cUG2GLOQ5I0+0ZFxKn5hT2LAkNWvNx38BwX
cFNPYRNzPTzI6cj/ph5q2BySIH6KBZ3VJsnd4tYhL2hBexZbtWsKdkOO5cT6zsCF
sq8ohEZYGkL/DZK8LvCvxa/G6bB/VYQAsgoxYOQEu2mLYCTFzFPj/NeibR/XQ0bU
wdLKQMar0vpuhz4129+iJMPJku3eHZ/nals5E/DdzMfCIJruQ5GFJqgDjL+GGOhw
NkRUaHBofAEJ0DvJMzuK9HrN+Qgz8vd9RPy7K2vJqgcpHt7MBksLsjcgNrsTO1PD
se3+74q26TDqueWuv0wfo2otjj7+sPMB08m8jFA5RsQg8Om7dtjwKjDIOI/peuN2
RI3W2I1sVCWxlHP413TJMKYvoJSK1QYc1SWacBQUkypPOnq9q6Xe9a5y6PIojBlB
76j15R4EjgwK9rcv8TaxwWm5nlt7xn1nIhyrfYPDy+QJC6HUpjqYjGCx64I9Opc9
Jj5qsDhkKsS5LdheEVvrSChRYvyqIfKkQb8h+E78TRq6Y9oYKkrTSvQfiVZHMH3E
d1xgMZhBuBoSUR/YEIgUVhQv18265U8ib5YqHzPobbgG6xnp9q2eqCilF0o6ucB0
JHUbqum0MtmPMwxcDu9doS1zHnc+5DgmLzkOdpdU1WRDgd/Bs7UfzTNem/Wm95aA
N6mUmfs9EpMoJr4vqn+6GSSM47FdiHC85FsMTfuXUg4xJxlOutpsxsnFwPkxw3iw
hVsJDvJsQauHRu9HrTVp6jxB567dSp11bmTayUWZ67O8AXhoozojAQiKntQHSkcl
mOqKPGQRckyEW8l2HhQrFzIyHzoQ3SGYlQVUoLXoK0zsMSLxOu9FL1pzyTc5zZNU
Z84qh8xW/q7qF/jhxpJwWMzE7VFDvneueNBPAPn/rROK4lCKz+FA0PXEG8CAs94c
IeiRtQd2T9cM68u5YF/sJWOhb8hDWw2y0GofszCBIhT/yGgAlvc530uPyYMtof/7
JEaAMdjsvb1ScO2hHo1j9e7w+w/ul1GFhY3X3EF8SHxmKMcJ4/FH8fyJRL2lZt4/
qwES3xIcqkPaxvuauvr0LYo5q2Nux+LFqzj2mSz8xEFq4hTPgAcGhhbfy8ewquEP
NE7xEp9oFA6q8AaEhP96omhqaCVVtbthIacKLfB7GkfiPA6L4YIktpEFkolaXp+P
qlYUKEEKoE1g/njkClOw3z7dkw/34iC6TXmYTqDr+9APsRwlZteXrCCFJRsq8SIE
scBKO48Img+wBqLi/IhTsQjkWa8osK+Lqnb6ScYkfD2XWVDoMUonPJJd0BVLTZvx
a1NQ4EW7lUJEnZmDsjngtFtIqvQK7Bz8SEFN0C+X1mnaLkZ0BzoCF3nMn8Sm48Ta
9JqXEyUwCSKeVjkxcvCwQHTtCezJufcoMfR1lrw10Mr1y6T3rJfaGIEJWe5yxyA7
7D2M0m42hNZpQ4e+0hCJH4+mDefP4D4IkBHzzTIv79GXvyLSM4dRG0rt4GibPnzR
bgdWhzKDijgnU3YsTRGfViCvrvO709yiO1uj5WT7GzJhORTpVcmVCAzEU7Ewb8b/
jSE78p5IWDNviU4lmFDgrE3I5FGwCZRqHCEW82LREcBGDjCDDN1/7aTIdCLzlpSF
lwz/ft3rn64nfrmmB3puO1vLXwprKr9ksX9JV/QgB00ZvpAFzglTq598iv32Vj5Y
ejfetKBfQgSOxmcCWRwOi70DZcc69Bqh2Sx+LvsEmVGqhOebp8RoeeYxo6iAbdbb
QEyUSvicjUSAOnD7WrK7Ua++zsuVuvocS5so417KT9etzUJLmpxwlkxySMqHRjrZ
vCsWPBrB/mcQs+E0ey4PIanNDXbmFY4OY63H/ZaitYpePB4UkArY12uJFvwuDfGw
vIBsFtieJvXYEKnRlbGd2GhwnB8kcTeobsqXOIStrWSmzN2iR7kapDnJ1UomLkht
9NzEjzVWMkV1OaAvueh3vRTzhImJBdq7BZl18DjJbZl8s/JM5+O57unCzKei7gL+
aIIdzsBoystiwbLK/CFQLALfpOwAAAjMqHPVmf5L080hrpxU9rTGmi4akpw7DamJ
zfrQx9zgqO0IaHtAb+SVrrH/WCo2dZYJ+LqYv8CqjPIdEzDBnLM9kXibDMrlr7jT
Fp79P9ObDxkBp7ROYu80ZfdrMQQ3GQ9JP7Rx3JgWzr+qt2+U+AybpuYnYxGbb6mZ
PG3A9ZH8H6i0eKRkNeJYEZM4LnatDc40vUQLMjDk3sXoRtPyJ0Mq9HaeSENbtJj6
+9oB8UZvexbpn1y/FWmvjFTbEmekUQaf/WCIcKoS/dt9m81KfLdqX6NhCcsGcQtK
41hhwSj8jbEXQ9DueXcf3sEoAMGM8D1c36qZ+Yk4IVKI1LG3HsgiQpmN28C/XBPM
+fO+hVooVQWp/WdA3veuqk+OhbLnHX8TKEl6m9omX5cqj8gQ5gfJKkg0J/6LYbl3
cr8EbRL0pS0nTtzVB5VbSWrdqCfC5dR3aPkCjEPMGiotcPqrKHT1PXS5Ab2pA66n
o+0gFUXUPtTEhGBPbvIiSagvc99m5+4tR4juqzNgKUeuV8bNT0e04UguGb/3MBuR
1jb+/HGC6iG/QwpMgRg03d9TqtJ0JEV9OHSm5OF4pAuQfLTn6fqpoVHce02GP8gL
hCZRNHd7011r/wprDC1lpprqH4aVcuYWsZz3DLvOtkLTBJRSuDXaLEgm38bsJo8g
bQIAaY9W+KWjFAmYxTyz0rWSJ0x41FhGB4cnJiqlVGO65iMRuhK56EctTqFdBYvd
SRzzx4cQn4TLY306u2TWF392zmtGu/n2K0un4+CfQZHOccmjtGc8iEKarIZHrSZz
zmBeuU56X5J5+iE2nJgmbTLQMlDkrcAoKBSv1Uyu5uQDk+Hc27nQrLzSFk7k3rQt
J4QQyHqRKQuE3G5A9tLg1zE1yoiidgKLvn4F1STGN36vi6KMUuDaCOmRnVxKteHx
yCI7p+UjtNcF7MBtNjQbedSWGtvM/ICQ9qcJ1FxK/BmGuPqeUjjj49GZmSFvZNOw
ZxSJKhP+GQHCqwxaNiJLYTEIjk82miiWrgAAYvEGE5T1KBusQnBcPT0T57wTEyyU
U0TKXnqq5B95iU1wRu0wwtTaHcrlbrYm+hzpDVpYPNjaWN2n++CXgfHe1pRGL60S
LW51HPBXWvLSPy3D7A1e3HgLloEtvMrMQGn/fqdJshFBv15kVOO2+ol1kPsNVa2L
WMJSNr3584cREF44OS6iN1SNMSydtXJ20QQOKxgJcbT11iW5OVe/4ouad9Xq27F4
ffVooqdfMDe5lsafjF4PrdmmtqvJEaPaQVdkpVooKoJ/Cf4TCmyyqmAyvQ3GjzYk
Ym5sLuRkkTh0KD6wcoNQ5fAchp+mY2kvafl8XMp3/SGjLIzIuTYLZ9Lr2xbcQ8op
2bk5K4ZHM16Z1zYIz2cxNtxJ37FKkR45QcGRc++AluDl+qZLDrm1vJf0a8SKgMDx
wGb7NhpSMyNm9y8NVJbt2SWeOOm5ItF0yn80v9g4nliMzLSOG//Mmn+zD5EXZ+19
VHU6k0MW8E3EUbIL3ifUfgZUVIagRqenhuJevFjhnFKxFAWkPm9S5BKZNQwDvjtB
i6X2NbOXu+gLQpNDypWSE65xlfZ3AVRKmqdjxhZ0GyouHsVuqcpmcm4ZnEbZbv0O
+D/i1PuefTJGOd8AwZCAAsUzXIn4uOjMKjxtfYD3lINArgd//nb/piGOmSGLQPLV
Sy4vDvzD1TxYnMEAV5vhBL+4x1s3kSiFlz7Os+PGD2/rj04iUhP7V5pyAEcMo4F8
NXaBIWuikhqdTqpzs5Wc1ItFTRvlm4Lt1r51nru51xKKPRYf9yIw4h5U4MQ88nFE
ysTEW+yMbWHaRMioWQGxrmeWc2eWndnJ64MBEbSGsf/lR1R6hrNpGABUkiYnDVWd
4MWNRIVDIFaK8rrpKFutyz4jO3g35rFYTSoO5ZmZvWOAs3OZMpFOqOcBYuPWcVb3
ctWRnAlNzg2yrinbWl09pGQeasQDLRYW6Tt9kWhvIouNxr+gQAd7SH0hhj+Y7QZN
ytf2BMiAFTjAYZIVma291xHhwQD7oxabmN1pBgAwcj/uaxlFkCZCaA3tWgkChm67
2ow88uGermKyGY9Lyk3JA/MOvHdJ0znu4OmSnRKcMXr1OLDpOzHLBPjBYz1Fefv9
lfgwnE/nyj3yb8vgYYoEjtxgNkKVkzO7tac3BuCKBrc7zj9dH87GdldzQ/jNqury
7EodlCBgxhKeoC5Nk9zJWkSBJZ6VaTdWSNF+ZdpSNmMnD1caiHx10tux+GIFQ31K
8ogjsVHF5eMNKRBSBJ24mosHGWAG0YhvisQzK0xAPZPOHAsD6QNk81nDRlbalr+B
eqO6M54bBjlFZUluMWLzEIk3WsaT3pIXzEOlT30Lso/a6PhsD6rXukkSgvbVY4gG
DCyYoRUcq4xq6S/xvJiLuskCGCjOlrwso4L7tCscSRYWVdRIeewiK0mjLDlSbgSi
UABZXuubFuvEaCaikqmrpGQDeWLf3NV6DO+h5nfZRV/EEGiacokcESCYjrRZB50h
5eLQtRLPYURFASgkMpnH9Ne0BYMKaBJaifcewSAqgB/GbyAg4dRN19elb26D7IGB
ksdEd44VRqDIYTjsu+2K6wKadKHVQwgLfyWs8cIChnHB/GKOGQffqg77n7TP4fyf
IffXe1x6oAYBg2+VmQ4tzPjaJ8USa9yRC632y8rSX2a23mVmRfHKQ5l4nn1STA5C
rT+TFfXk6SdoGvWQgLbjgZ2OxUgtdgPwxLhfDMRM4qllWBNiu0CFQJ6tdliVeEdV
4UC7e6J+ssYNbkMIU3JeI4twPLo0tQJxBOa7SCrhQX7E/9dQEgJ5EY0+oj+YraWK
KhpjlmtB87uaOdtGwx7zs7zNoaZOBddL4hBWVxXHPx7f2Ak7TasvjSWj3wNHMUmN
U3BJT3vpuhgGungL5go+V2GDmdvM4UpM4ZDmFdF5gO3hDmS39grgHc3kNtBIYWHS
F93O7ErzLCo5WYFz3jlCPGipR/dBAYJ6DE4iwPCr/mPMGHIqjw91a+0S69tY5lTX
Ia00NAZ1kRhFX7zguxtv1UWUhB8zne3a6rqOwKlpAM7to+reILzJqexI9e/zO4lB
cyBO2JsfnoIyAji7OWwWzDHU3C5FExf0boTBeEgzJ5mHbrH8w+vHOPUHEGbEbvWW
ZEyCIcnYfLh+ff5+xnzvxJtpGHDc7RxyuUJG1BmDNfh3CeQoIk+sTWIJITU4ZRWF
manQ/J9uarr7yHXZiYVaney76boCZ6Xe0xZKqd0PQi+6dzs1ByfIUFbXeBvKu5wk
wGDMPsZR6jYVDRJVkSlIQ6qdf/UejHlMfBmOYepi2jCQO9YYanal8JDGXIt70upE
rJouppdV0Lw+p08kM4si9KjP8VkWgbD5te2d3h1giiZn81ublxSN2YNEbC9EBVF8
vf6US6dxVulPvFH8ItbZBZc6hBy9q9XN03V5OfzNFq+9LPgrxYqAKaIjXTua+cho
kbK5WoMQEsKpuGlW31JeS/mHp6LmxYtEg4IC67C2f+5/inHhCKV6kp5VyC95FClH
RpUDx7HqCzv0PjtIwny/B3Y4WenivM7Oh4gErntjLuqGwsrE/dDJv6T+4/ajAjd5
zq7F5NEzdlvOWIQ4QtLxJj43whQLuFBENgG3kQY703x97iIl8n1YMImZoQhEAMLw
tnViCOwdYVuZ9f6RH6uxLTHRxz1MAAZtujy5GkuD8YMPPkxJRB4WkqlkikvgIUBS
ToVBDh4kLia/Lx51eWXnXGwa/nbSvx903O5/SZISEcMK8FZjuuVuu9ya4whPIEB0
YQR2zftLGVlZB9YWsHSuQcHUgNYE6p5Sb/7ms6CDbfpaRYbtvmSRZN94B+m3x2df
VxMFNHI73xLoNEmk4LzPGn0zMEVoEZIlHIIb/wQIzVmifHP6RZ9yZuCXOywD/17N
AAwLLiIkuR7pjRSvBMF2hn/5TpjVzM4y7Cs4kz2RY/6OG5QTEpBikztQSee5MXK3
8QjNTCiNuedOYuL72Ll5/8RkSi8g9aK6Kp2NQgJ04mt8MwzHDw2UDLovAEs4yVDs
gXFNQLPOC7hZDQCurKoHXZyq0dNZ6M1mXoJVnyeXYPeAPFPnYpi1W8gVvNfoK/kC
JHfO14/LmteMeQT/gAlIgdVdkErcBa0/VB3qLJ7HaQoVILH8uBU7tBn12kgo0rBW
z/qCf9scnOr4bMzSC7Qx2RJxfeJyL8E75xeBSYsqsY8BCb0+4Q4YXhGOHfzZeUZc
p6uOxOKdKoQ5+a1WR866oCCUI/mAFMAzlXfu09Gm5stAZvDnD2smPTJZmMR4DcB9
GagExbZh5NW8mf383fkFBCqftW81zx/IEmXTrFz84Ihn9yUC+PdnKEqLBwhZ3sic
rl9vYQ9TpyXU/nVTHTfF2YPtNQ2pKq/R5krje41kSkOOwXnII4xYHtiq7+dnX4lq
i3L/3G03mdVh4Yaw5Yck6GxwSlTenb7BkULfd3MQsESJU24wmFjx3jm0dyimETuq
nMEbKiCJabBfbclAuo2RiDAP+j77suqY94yFv5mOvrWmGNrblqv7OZrL+XZS8Oy9
Iix1tI2XOKFCzNlupmT0Gbf+2rCiPAhkFCA6zcL65VSdnSxdP731pqNFZKBn8eh6
qdLE+zyDJKBH/ObrPYsnWNjGiTXMvJCTpoVbdfFP7aqBkV3gjWhA8HN6kymi5H6V
5eE7yi2BJEO8oByKzb87EdqZcKyzc9pe8621zvKyx8OyrhD++91HPk9KiqOugc0t
2eKVXcTi6v8aVDch/5mZlCFGXL/Hgxbw4izxad4Mq5QW7IKko9r5s4PEBSxw41AN
xL3p0hGtKBI72KExp0e/13rqca7O3zjDrcBmvDKH/qIoktMmjiAkF2i7Zh6Bj8/b
UuVDmQaE+huijiHOmXWdyy1Hd6grRos8jRMnLajQGkWO1PBK0PT+HWDSXWgw6yRY
Zq939eAllPgtjpKFKnl1r0l74CCA3A4+vZZxL9nrqDWIwkowgr69tGTbGbkGDdoZ
RF/s2fhq3Cow6sarDQfkSNuz+9XCcQmMaulH3YycTjMD5nONhTQiyi7w4Kr6Yein
C7kn93ImecmYT+9A014Gtyrdw0g1cCiznjsQfWmizNXgF7QuDrVaWUGCMeqC+FzS
j/JF5gmpHAoOQIBrWGQy2ekNgzVRM3jw5VR6yjlEkbxzBMOrSEx6DTAZBNF+7988
sMVBxd1zvx/GKUBFHDDbMy+iuCF37/h/nL7AqKZ7zUGlhO1PzAydbNxAJtuK7J6x
p3uALchUEX7HCPLu1YdhT7/QixsC8DaWa1N8ppbF1FilyFd1WOftf8FKzDB2QTOV
GsdN83vT5F9cjJwiUhF5ORfSErFaYerDDlpWZ7I/1TmEG6YTwVKFn/b+YlzGl2Ri
QVVpLTL47AxfnO5rYzbQSxwvYxjNLxXVhd4RSoxVciJVA/Y7/7zsHHrri8Y0OJtt
Mj1JEtbywTLLxuGPUl+/Hu78ia2X8nTOxxOYhXtiKZO2TKSFWcyNLJxBo4Hqpr59
UKUNB/h/9XZj+TlqtxTy9ObtOw25yo05NG4Z56DPyT+f86TSArOr1CCbr0Yi5Cb5
f8LKAqGp5xMCICyzvTT7b1/sQ+XHHj+PARVYZd8oCvIzZxjk+Bfy3WP18RSZzqy9
rM4bn+pTsKzqz+tKjvnc4yAo4b4A3G3pXiHWk1VT7Fhg7hzNkq6x4bjGNNVz+HYr
aXOsY6J6N5HOwolTwnRuJF8wKpFR30XlBpFWeANpidZLrwvz9DY3JeEhtWiop2dz
6hWY+WcXGBcBG4Gp2zSNySiE+LlOs0sfCu7u69EXcjz48nRlgLa3YJqSuuBHXbOw
UNV9khalINvD5JHK4rRD05glFFrWygvRn9wBEdsLA0Gx/yp9UZMLzmksv8tjUWkV
x4mNf50gJ6TqByodGpLLtI2w6cd274C3ZsddKgcMgSZ9kD18FEWcAHxr9/uKmA6s
6aYfDLDwDatWNztX9gjVnt7ODChXbT/90oB6rtxwOfgsRKcyoWerebpa6xgN9hDa
Aw1J0517+8Y4DoK8GZuE71XX8JuCWuUYtR3vFkWrD87x7JNtKiMcwe/1RkX34KaG
T2VFpaRhoNozblB1/9O11VbotyhoFhCXOLoi3KsuYitT1++0bLpSwi0U36VD0vl9
76Us4IkpWiagbYFu/VrZrAuM1lgVsWmd5Jc8jv2OzgNIrNH5T+63ElkTM14nNeN4
PA2UjTZoE33W2pXvaT79gO9DJ0e2/6lcQ9+pygpJg5G1a7y7bcrLr7XyxUKOei1W
FHs0DP6ad9kbWUF+9Wm6slwMcutmPF7jkrobFSgVseiPwFUO2dt4FkZPMLKaV+dB
PcS74pmE2luqKWNbWbqOcJ5Fu6zkoOGvzYICzWPG/mfAg+x7lvw1CBJ69YfXHg+V
2HF1Ny3t0VxPpsvnBG5b+jvlKU2npt/KFjcKyVVaDvw2Vk9q12uUGnOdk2MqtB7/
8xgKAbsHoVZcPK4JB1h5MKQZaXgqb7Dn2tFAHAt1Fi3iQnn46nZetRCpaqoQz04m
9es9oh/5UUbPUJsWV5IA3KAKxNQZzgksqOpir8BtVczYU/8zS2Zql3CTyVNrVozR
SMHDCv5LNL8mcmCCOPW618tLc2DOWmCAe5Sbnw9yw2O8bd8o9vfnfQ8hPMQwEJSl
iTHrCcAr9hQ4dIzRRZX2QpKfDLqFWKWxgwZoBiHuhDZ9lv5d4g3gvhmJ2zZ0svOm
ZLPteIi8Dgn8NAVwN80+5peY31f+3eWXS1PhjiC1Ocz8bS8Og1PkeDt7MorVxzpy
eWrLPePM4/WcZnHndnF50JVXfvuhuiim3m8deGqSwK/fK2Y8ToanBvIBix5oo34l
hfPAB7v52IAqv7hPedxq+dbuQ5Bb92b3/jl/3shBX8cp2I3JGwGbv+pWPHjrclh6
bQF3tB89iSJrHHiCk0qhjc3seCXyHIxuXJ+NT/Lz4tJF2tW7UjVb4SCFV1vIutoV
fmg5ut56VVP888IGc6UM2uftPDgrYzIjLAcJIGLoq2H/vJyh75STzggVyFgxdtWK
ZFCWGrkE71A8/1aoTYDKkqHGfF4LXv3vHybRcj7Q/Becqzdu2wasIPoPkA20mCKm
XEQJfB6I2Ep8CqSIj9hL6j6SaMoe0czrAbPV+sOqDT2IhRlJUxFZHXs2R8W4++sw
PkjYlyA+lgotqLsgaZQfQBuG/RJuCEyixqTrEmmFZHIDChAWnWnMQdq3mJ1oV9s3
ka6jC7Y+Aj8OFoC6buTiLQURk8AY0+N0WQ3/gsSD2TSOgrY+ZL/7XMLCmHWCJuhS
hUy+hnkf/yEikfN1ugZcHUAjWByalPUViTbD4LjBoiGanV8LF4aMEa+TBhS72OTu
hltou4ydJlhaU+UnRuTWDTAimMmOumZ/lXpdPEKtoSwH/C5zumDCg7ataZV0vWY0
Fd1R3sbeOsjyFSXGxgb3jYRJorMOxFrN/09CCvTxwisLoijKOk5q4eSSBwh/MGij
8+p9neipBa98IKjiLxoUs2pfNG4ezbN43sP3NtD3TBxANECEjS+7eafAcQxIqWjV
Z2I4U5Yb1PRgu065rqi0+Lkbuly6E7ou4l/pCnxzr5PfopxvIrkITzYf65R1SueO
7hjqVTeGicFVs+ulKe7IVjOHczjfFQCDBOv9G7RXg7Z9/z3qggxVtqvwGnpynipr
cYcVv/bgHlv4G9wNpAivPCGc64amQj1g3MNIiNkKll569p7Jm4WQCpduEkdOoE+X
hZzoLjNxF/2Q8swbEsa8vKm1xkw0jiZkJ3PhAVfUErlkZ8qutFjLv0ffrWpK6H0r
YB7tQDDxxclmRYRiqtQP1FnKUi7Im8eFlgGGeMzowl7vOUCvS6v7e6LmvciXFtcl
b1IOrkdvKRvnClMFTQK6VEZNfpKwdzi9arlx1mUzi+Vqme79qHor7P+AddIqnWD7
QUr2g95080CUgaSRnewYs0hSAcL57XYfJHTKoDfnhh+dEoCFngEiWQZhpKFqZr1L
AnDnTUjNdG/d4t8RqaaYU9X2NQpLLp+yXaeiLg7PZs76+p1RnUmdbcVrLym0a3iW
eeAMoaIvSQzWGZB+CCjf2wVthTjAMOYKgrPywaDP1fYamK5Hpcro3mvavfyGSbgn
x7r94QHiyAxoYVKhbHSmxPKWYi/fugI6ubd++bPNHHJm6nYyDkpWvyfeWmmZSq5d
kwEfsaHs0V8U4PVXuG194FsfR35z1Y+iyUHTSLIsU8eiGbZe5w1CIBg3HQ5jvUrV
a9fkd6uU7vTD8sujL5wKsb5fz9b3inncmy9Oe4y6GhwEk1cpD1h2LsWlMkOPdx4Q
sG3yiTcu/A8o3quB3aD97GzAPeu6NIFQK1dWuaVpr0hs47D3Re7oFP442Xc61QD6
HJThPuJ32/WpNBiL1pTyKpTCHFgn4i1VVqxMFB7NCrhXUyTp10ogEHnRFnRXtNC4
D3/9J6OxSNcpq5126X4fP7Bf2GMByHHUdMMVAxYRj+85j0gbjLu+zB2KO8l5jjdy
wEc5fQoLcgwQ4ArnqcYvO3rltQ2C+bF5YBufQIXprxivBTAeIwA8bo7WlJbCaI/H
pHCJv1J4gCEkDUddctiw/iAfyneTZ5fqVxFSVpWTSSOp+9MXIDuJg5ctls6B+x57
5Zba+LvEanV1IsWSefCPnerszt70E8FvacOHos6m15WqlUAnxWSpwCaXh1qW0tRn
IfbG9eDgsMmGddsSEBQ8rexFfh/8QTei10q3qsvDUFYTVsNckcBEnsh/evol35xU
LfQg6itRigirqyqjFS2+E4sNjKE6yKjH8JMvJ6KjT1raJ4NPkWRxZDDxp5vbAPat
6c0+KclpiTR6s7j0g1U86X05ZdYUfK3hFtn1sNgzRYLyp1/IDAsMp/n+dz3+7+IR
h1Rf7IH4+f8iQkz3vB2F+Sbp7eUOdjg71Cx+5r/pBPuGQLprnSqkY56XAjjpAcQr
ylOx/oiJF7ZERH5azL4OLomD+zblgfWwI0ofY4M8IKU6hgLua3c7WFfvOnCMq1Bc
FBMZSRQeSMvtLI4BXVAqijXtVYjtphBMaF6HMAvDeFeBzy/4BLl2X0zJR84TVsss
2JfAg5nfX6V8OyTbgK+S7BNsyz38jGCQgpn7l0XRZt473YWOdtgmf6QSVaECscTn
gej/I3bbrBrtRCsce+by4zzxEoKFH3d+Ypt6bD2/YivyzyxrAgxqdcccp2knpAPe
endi7KkqBRhvsRGleoebMl0hovjVEuzZm6ZL0TjY0CJtY5u8Hvm71wkq4zl6LvHF
CMmkBpdFOfqzsWgBOhIr18zkfQt6g0BstBp+VOkZ4LJzhYSB+cRNzBI/Ec0u4H/c
HrUGubNOru3jXJBQNJxczfCU0Q2TdNKQGzj1090GbVBmhnHg8pZfcpMHI6IwsyOn
xR3bLP2n5GoBKvMie86qQxssofGP+Cpx8E0gQpdCGMAbMp0NykBaWHkvWT7+5cKm
JuTBORsIBZbhpchNjiqu8vktFtrgBMvYn7cQ95ZbqBBckjeyWCBTqvlXJuoIRNsE
y3k53+Gk3yfhDKTu/278v9ixPOZYM5FwNyGSZ/fPIVALxDTbbUM4j56zk7JltJ4q
u8cGxiZnnTcStnossI/cr4uPecNqUbW69d2m7MJUOhUIasiIF+CugoWcswXWHnSd
Ynuhf8rCj9ab8adaFp5jUfDvs1lycRDFeR7j/MnFMNFs4P5KJQgeCEQ1HCaPb58M
V7Bsdzh303vgxSI2SLjMR111vb86H8fSV4KzZyPHWm/0x082+9FsOfX9XzUNpjxC
rjBtkjw0Psi1hcAuxHGq0fUw7EjINLtB/jnkcfn4mInOpM+RQLL5x3AtuBpacbyX
C8D+QocxziEHBTykwVJjAr6kD00yHjILoGMXakGu9Of+5R+YROppIDgIAwQUomMK
5xEUD9ZfeZKrIWdg+xZUc9P+c9ySNgFuaAZvO//q/JhOhdQKqayWUVg1i9whSjPG
DU3OIQJanv2okqAXHtA7lKl0ZLxxSqgsoeCttltTqEFRGizJuaZu8frN/JhhJQcO
X0ZRJI7whj9fy3NAW2wNfAHQk1fP4RGDJ0ZDTy7aXxAJNpHOdSzUYoWt1y3P1Z6L
Xe/c9Rys9TlaMzZTfS2NkXXto9ysbWqZ/iVcqs0FAJLFyEj0IDsvzT8SJ7qFki91
7McSRX9LGlkbHr0w3CVWzvSQZ9p7EC0fTZA9mksp81/BBAHKYuK4gpVpgwjcuc1u
DaVLsWe0xEH8YaKjSzyIEYYq4BDwM3f4E9/uEPILEzOwRSkYKMbzNfjL6v1rxUJS
NVH3p1P0eDi12gYvv/65B0XOsFOhsjjNpMyTyuoKab743MDG0RiHk5fUBLuW1n3J
If6bMmC2Isc11HT6uFC8A2hSf2qqoKP1TcdIoeHfX5EjbncNNZx/fDEOXHD7jBx9
nvCJVYCqZdU4rOzvJ7S14JsN288KINbf4RXoDRzOpinK91Kd1HM/1Ft44mNYLIOx
34OS9dDtF2dysT5jN/X0/GwFHY8cBJ4/sWle84wjoUM6ks1PuMuIFIi+eNRYRDk8
hf1DK8VvLbFFPD1Q2S1mIh0rAO4YhLEVdFYt9qLiOVb+oqrkhjZowiYlmF3NSIi1
KtloZLFcRb9VYm1OMmWe2CqfFzbzJtD6/QUVTVWAp5aAcFti7wz+hLS/VxJhtzAN
fqE8/AXwogIRXtBow/d6EY8FcvgoTlyq/MR5oVEYqm2um7Q52p1dadYxtgyP+me7
wOdYS/3e6k0CHsRmCYQv8IVxfpkH+23Wcip22u0KY8LoxfsYkJQM+L1F71X6eB/P
KtRB6stQXH93rGEEzm7GXnc0efLpzRV02A407FniXgwMdyyLA4KEpp7ncHaX0swP
cR/jQGEGE/+hUWf1Eg9ePS95v88nd1gujK/AlwnOSY80mvCpf6876NIiuHhbZgIr
QmYQslaUJR27QC23Ws8K6MWJnNDywFFfLzAmln5ZJ/ot2mJLB8l4Xn8/x6sYnxRD
OVh51NjJlCJindZ98gb/WH+vx6nIok4KDRHmeKyes56wAzef0Bvvou9SqBTI3shE
kCc6LnbxhAzvb18DdsaiQhyZ1xuk3EctUvRbSKs21H23S0gjctXyqm/gNOXOYVkP
yiiDw0oj5JtzxQZ9UmQpuEuJsuZhtGVwC94hZob04YCaCUBztw5VCjfz0YR+jIL3
QHTNuUWJrKlcTdNzobVzlj+dF8agI+EHuCDjBbq5j8bPatXPKOXWBTpuF+bB6Jgw
z8tYlRPof7AC4DsPTbEWBoVpzY5pyfhord5f3r0Erie93xy9fLKays/vQvsVXwBT
AdJocWNPwSpKZpG8IpI+rm4Sk41+tfRCm7lM4y9qJlh2AzG/tAa6+aAo2IPUyEO4
fOWTdQt6UE1065i/jDtH36SmoAHmJYMnpj+t2DkxzArKHsi/0bn+U8r1sA02FUbN
nJUo+5kSTwcuraxWvzZaeGrcrten8mbjJEHx25gtS7wnfHZIbARzVHPB4Nqpfl4J
+2+plcCOQsHdDA1jG+htqc3vH0+Lte1wGNasI/ce39i7rGwv9amP9ylZOtnJ/XEW
wIGu18AFKYIJdV8WLeVApT2n8wRGv0V9Qih815m2wxemQIcw4Y+Y55iOEqIeyOrd
py7gbJ+Fa098O1Mgiy8BHDMXoU5jNLarphiyVfgkP9WUHrHSCHvFZYNQNxc2yHuo
u+UyzByBjwWu5AhxNstMhoMZVT8AMDKuWvK+7ujS95V63ow50d1uIE7iT9U/smM0
AoCJLA61HBps1iiM7bd2WUlklufz5g7Zk0A7P+gD1kfJS1xz1yIUT7sDhBXm0D/O
CNAZsCGOr5/QX/5WnrPIjhFOT+2/NXT6FILevtJwa1cIWXEZ5J5LJfnsuqsGmlVT
wdcDMrbKtmyYGdKT1RlnfDy5q8n0whHt7szbCfmolvw8uBGR/38iVT17RgWfhh3a
7XXm5qr7RaVxQYqHfanYJTcgNHHPmrghoarS9BIPhg9GYf10mh4vISeCq/ZabGWL
z2LPtl9gbgKZSo/AGvsRg7zXW2b/jQmJJGS9d2P9aCZE/XQymfF+I+0id/KtNkTH
m+qpY7von1c7Ke6pBpuj1uKv7UCK+Vutzl+talmPB8KiQNPPXmB0tI2o3MaJC6T/
YlX7StmfaeUQOHQ/VaoXlvKoxm8u2auTjZakYNKYA1/Ls1wAcVymFdsvX4t8kOgp
aJbyxabILW6p5yzO5JjPBTew7KAJIPI9cgPCmhZRw5ljvaSdQ18YdZQPnNK9HxRK
X3ltrWe2lWpKtHuZ+ALjDMnJWAA4mVvs2ZI3hqRCkXKFQddiVIQUjBinZkDEiUn3
IRB0DoDchd5B1q9v9/P4bk8kvFWhOsjTA4P0ruE5mdSrK4i0WFjlsCRDLNpdLBbU
BFXMAgfmluk5pz6nofzhUgbOui9ocdsicPpl6tVwdSBasT3vqgPvVDavA5vTRN/H
aWO8/+zlC8OOUVgFAfPB5N79aH6VgwSSkRz7WE6xfgCKT3b7iB8rZ9R3ShOZFFWQ
zlM61UDoZibW7eJq+qovZi6ogFAqc24CrjMyQCPII1wSQY0pH5HINkrQjW/Cl+v7
MFDEnp/Ach7vYkrP69S/hGZ5jU5htEP3mxRwr4u2wYAT7c+k13Ojsqkx1e/+Rio9
xLJ0TcpmvgAuXtOYcH5TzVjMS08knJ9tZQFhdYG2I4aZQDNpYeXJMAu4Vz3EFdTS
vjbwS8EkMdSh0IsqRFfy94Ob0HxhTC6zGzahjJ4IZt+HPwEuDKSm3gYmBtoxKy6C
zfmEQuLleTP3RpE+B9siKkyzJ5aF/lYDAaG4Ys8ABkB74Q0fw4ahDWmlXwUKS+zQ
8SRZI/Sji/N4GwQGYfvndrO96LW4HfeA5KQwTVOwjKkOtI0otaTf7iqlrYLXnaQH
NbZ0gOz73gACItnfK8KpOQk48uOvQ+0cU1DQxjBJFA7PbwN7oVUtwnq4FpytVs6+
9iPAB2vuCPzav9Jcqa5aKvVqN+oPHmA3Tlz2YJdDAOeehJuzFw3cT8E7eWdMrvR4
ScmNJzC2QCmr3ftPHHVlAy1/v7pBQcMxiwTTLnr4Xfgo4IKtwK1T/PUb/piESs1G
MD/Thb0F0kA+8R5C/KcYEDuULysBKTbc8qdteXN9P6ajgWlA+oZaXl1MdnvPcfaE
AieyNR/dj3DKdfHNiyZxy05p+An7F8TfmoMoD/YSoAY1++CHwHKpMnxwpILmnaei
iItuCUkkBBVpAb9lLCPtQPVuwSorKzvCZ6qB7g72Ukybwz5Tb66I0Zq3ktckcc0H
3plBM7akioMxcM0y3f4pb8ch26RvTRJeHthZVzqOHRv+nIzyB08tDlSDlVzajLaq
Q0cx4ratXF/MsQjZbaX+HIwhDERoAt3o50SH+izIIy/TqvMK3BMAlm8G6Bal4tfT
xZUuebvatXrZEXx1kqX06XnDFCUizSoBPGl4Tco1ltdSdb2oLp5hzKSTLOf81Sv4
KYGr5wxu0+A6bL0hDtXvriQpYsig5QkPIxNDodGE2fIQ59KQSYZ/9xTDk15mR8xg
JxaY461wzxfZELDEMOdj2ZRJtkuDbdY9Ej+kocYcZcGm571uA5AYyjxfJylAQE94
ePn3zP0opxcsiRv7h2p+hWWpJdGNA35PwEhCj9KEwyjLC2hhIlpv/pbifRth4KsL
VBziEzs/DdPm/0CljOh7P0G5nOXhh5qsRZ6K1RmECpSvhWFzNuib1Ck0tuHae2bC
1cgct+Y1NgFIctfIcxE3W1Atki+m+R0bA8EjQGdsrZM7MRUNwhrCESqcYvT5kiAn
6A6x9hEqYtv3R/vgYIyINNk/j8Ew0iM9JqMDwqmYE4x62rdmRqOfyBMjlgd1qJ8f
JDq5k43Sk2XPGOnHJJykKBZQv3BS9cDlkygluIEZgPy3b5a4DxpgGTnLd5vN9AhP
BtDv0wWl0gNg8EhKiMmDC3unrcrFFogeZq4Eu7pLYolPmBhvsOD33m6vY85poU6R
aivwRF27hk7AM1bynkaZK09DrPUhcU7XSt3DwSz/4IsGzYSEGwLgjDsqrr2dwk3f
BQPodtyd3TfFM+CWitZ6SaurmtiLb6fYm4GSnEStpjNYT6ckcWtYl8QxlUxy9k+N
poXX+jJRl7xPHi1VyP/q6hSwgnlT6rAJsa6FBA6yAR4i1GgAI1F4pb69NzdXP+/l
m22kevN06FOLqzgld1Ja1Mr4rdyBDpeXSO3F88z5+lmtTfetYHfR1a5St8G2Szbg
9x3i5Q4LgEuAS6IrpUvbCJKi2KrWqgvwsxzssZYvXz9FJ2FzGrexZdyjiZy1vSLT
CyDb64KIiI17qP01iJa9PjHVYzuPffsGqhFHg9Duy94NerC2JQUbGTRfzoqBmN7r
JFEAZuWPW7XsAcHsuKxezzAljqC1/0C1YRxRFzHW9jt3FADG4tQGEHGerGlla3C6
aL+1Qsouyg/gi3IWwuKbk4VBVbCbZJv5WE84c3uj+FlCa8+eRXt7nN1IRUrwdohi
1lzfw+okRXfL09AF++LmVtYEiiyYdOoWadoxl04nXL4qNn7CcCbC8baFOegqqjLH
waY+TGzxbPAj6zwsnKAYOtFreb9Sxt3gNtPG7KoRKSn4ZX/3g1qp3LUU1u6yMAcD
6GJNw6oyl8pH86QcJWIbTDhLVnAap+1X8b+7EG7fu1nNjh61YzIjpCMtWllb2PFX
p4rKpBC4i+EcQsUv1lWkS79gxqJShuYS//vbLD5W4aRqp47MEmt+iVJ1BQI6B55s
f+Fd+Gd4PwJUAEtZTcB+jxIBkq/gCB/EvY+jpT0nDDYbEu5nZIPvZiSYtEGead1W
Jyy9UOcg2f8E4hv0OUUuuTxvSsP/sx/mMAiHppJ0QplBRKHKKGKx2Y2Hbf6J5yb4
1W5ybY2eLfJnmcCjBofw80kXTJd/ab39ta8PIotuDQs8S5AU6EA6kRhcpR9v+yr0
8cOKHWtKpwTJeHiGi66ZTAAD7m0bOmxXS+Z19pn31ElGTgPQLVgoOoKRrNnP2fOl
8QXzWDtQ1kH08r07iy6MM67myv+k1uRFy49cpu/7kqV+LirxxHyDqjkifYEeQaiK
KXmj34/bUGWZxUoYifM/N0vEd5rajAHgAGKSEGSXACmkFo1/CUalpZmOBgfkeNqY
K4On7MjR4n0bF2zS5qfjMJAMZgy1jD4R5XSzIzK8cs6vKO2SFn6NNhj3VXtdhVYd
c73vOdzJS5rwsbVMrlxc6RN0VohxklL7Q1Fj1xzemCzDqKc9teIXoYYUDmFadQX4
Eszo5v09sYC1dlpgPNNMWtsvxAeKQy1r0wa7Mo7+ouXvNjzuZqFmUSSDbsQVM2fc
wjks+WIl4Glj0fZGRU4o9bC6tXFK/a4YoXKxpgS3VlsebCmKuBLeKxdF7BkUHm/J
aaNgftgn098otI5NHelKHAGQNLM7ec47TerVzjg91AU6rWlkdov2Gg1kTu8L3ZQF
GATy5iiC4ZoqKsQoKb1BhQaS2AydYQp2s1TMKc6pLlAOjqpdhVnRfZGhn8159+hl
UPnHZgT9OQmCE4VNNNvrdaqhXYn4MGh7zULZpHph0GzDQvZ/8nMnCbeRvGTVlGBs
kTYjD1oOCUROK89dtP9Od6fUgZYf1zcL7ecFFlrqatT41MxCUuZcKIj7txrmgtG8
RUzfYfnAByJrDKM1KsC6EW6rJWunAypy/CxO3LN8e2Hx/XH5gyK78hbYyqNe0JHl
vKHrNzlPgPxhBwOfb3kiAtHCFO26raeBp+v64f7o175XRsrsj0blZ02R8fvJ1Lcb
HUKBOzbOUAK7yukWFJk3CJs0ic2/WIho6N14NlPLS7rm4ImZez9GsjOR35xWUaD4
9Dkf0zPje5swmtqlqbqr+3p2DNt1Kk/NYAFKvGpN5ZLI4cMJ9J2Y5SkO2H2AKY6a
eu6YkVDfm084cFtZUolpzmhJUSG0U1Fb7IkrlVAqVj8f1ZN/PaPWHQPZPdDp0qXB
A20z2bgBO3BYycGNXrV52mpbvox2Rw4LFhA/9b4iJP31hx1FGUoRBp5WrGmRMyj0
/UbPbfGswc4H4ImVAZND9dwnm1+QLBNpqmpGt0uX4+PcYMD72YTN4H4COQNHUawH
ne4ZDd6upguWQ003Jm/zX98NHRRkabF6rXRBc9KuohF+zeGwsMF902xARyoJbnhO
0h/gEIi/wniTeHOGtJn8BibAcAZ5b72InkXQKdfHyEGC1NCSbmQVRAkIrULJhx5m
o5ddTqN0BxhEgYUVmUETucijSpQMVUw8pDARioh26dZJ0O7WOYWvT5xoBqOtCQOe
6Gj4BzeFy/vrtYzCVaiZEv4gxJiwMJCU2mlazqUtOvZdYtBDeMXmm5Kzw2vQqsQ1
1Nqta7r7JHLW5I9zKYTb4Sh/6mXjXUOHx0dgL8VxxMfc6u2xeLhYyDS6ICPFQyeq
PtOsq0mKkIaZBGEi4Dbl/SjMOWI1CYEbwl2yFeRpbHuSJt0IkZmosEZIS5seaBzP
BIgNjtPtoWZHqAfkrmS2sB7eZha5Rze+8WVxK/KuCIKdpYb9D/rvUQrJ3/+R5cOb
T4a6KHyW8Q1zufl94e8Kndthg7nT6G4X88wkqPN2Tj+dHWsiq7BTF97M84V4S3lg
KcHytjcMQChJt/HPsDpSHZQe1qDW8MC3X5NSAoKoxW5k8V1AystP3lXYl/x1H6lK
IPk6TpFRcFry7wGT0M1yt6btq483Seee82rad1Fh4jPk/bRA0ttUDmXcUzXup8ii
2msAyQe/I7L432YemTaxmkpGsfwWkOasGfJXQazh+EJc/XCA31nF1qz+bC/Ljzxi
42azLfZmyzilqaWvmnP3pk1Kc6e1gkqDWUqNja4vO7sNw36y+U1rgnXP2LPIqFmt
bNlNyVjMA1h046+b/DfXT0e/dyWyNwMRa2Q1h16GU6X2xgB6wI0va7+cLnH060tJ
53LnD1ttSfejABhSpAfZoRjyDxl5a5ZMBzIL5EPgwFaEixr1hAbHpy6xK4y/tVHB
YnT84Lya5w8tCQn6VRzRDfHk+3HS+ZoWlQ2YSqsf/kPVCqNbgIUuDXo1Gn0WcE9B
rTevsy4j49cL5vPLDxVGEMmRO69yOaiAN5Sy+4oFUfJ92sckYJ1zQSFh1Lg4a4te
Qj1QpUENmn3AkhZ8dqDU72Ur4ES3gxJt4PCkn8qHOKlZzsxmw8DVsIMRkLKntqsH
+qKwF5joqPDfSsUD+uIiM0ip78nnAu4vr7ObANycySx+GbyUMcDZcVTv7moV0m3T
QdCnRMBXh1Pu48VRuOZYLw7tA/iwiU1/d6OGGsQ4PgfEdAecQaYhDHclNOwTZEtA
fv9ygG6/gUTwrmepA2jLzMoLuJBE95AV5RBsmqYEK/0JNUAKomXdDT8p0Q4Fpm6J
6RXgcqbzbBbze9CQdCGD7Rtv7Jo4tQRwPl0G+EQZnqf7TLv64XsbBjsx7NCaKoVm
mbTt3CSoTeJzbVR3cu3I6k8fy6wMI4JKhQoI/l1Y+fin3UGEVzRT/LiPy+WljbJh
HWw3HSJ2gBv7tFf9wTymyLozchPeFaayG1iNwcd2mB8zjUEuLG/CbiFKmYk8wIIE
QA/pWPgp8TCt6aIQd/Y93PfCEyhMbxu8Ab1VDIJm6zAgOZfmaRpsEbqjjykgMG5E
Zd39Q/BoI/M6FGytvX7caiwVh5t1IFVeveFDpDENswC8RskTQEEm5Gjzv6VqvEhH
ulIV9482VMnSxHgBILWePUZqM0YhDzbaKuIhCPJ6tYFnB4EWDEXVFjEAMzvTMAlO
aPf6pubQhUugYmLNUQVxL2UCNl2rPpEm5L7+SY8H+/dSNIi2OrxrdmNwC9BIvRSs
OFB8MxyAoU26zhmOvWXvwss0zGXQYD3VpQfKFAJyOjNtp1bPltTfeGz18+P9ivZa
8CnaHJv7HdoJ0G/1qwLE8UJsZgCOToZzRCS5FBA2Codl3h/vQQXlT2amIlqGYDgM
2kNB73EkFBZ0AJS1E4t03EZa7vg7/1jk04ffkmh2Q3h4dyyv0NbF1KaOnyXn8+Fk
y58olEDWjetme4clZjKvYTqpKcyIrvQPx3l9v1Dl/3PaVgQJ3qD3wwJ1UCMFR7HQ
8EncYiBxKKiexE/JraW0GW0udzUi96FXqa328DMW+IglNRBCQclUGwC7cURtBeWT
gruq8eXAbPICANl53UiaP21c6OMDtiBg/Q7eIaFDpP5ZgHmO80UnNdOCPWpdHOpW
1xUFGwDcGjv7DNkaxNThGkRUKbcZrf6itXtLw/Dt7xL5lHwKqFEisEcZ0DQd3g5O
iq5Baill7Y/EUC2DbieHRsGFhwBeG6rsVo0+CedEQD9LmQK4z6oX2RnloF1zw1DA
XdJ/d3hvBQEU3nO3PnDNvdkuDhRrMTQ7zaCnMKYrrQa5qApUZE0TXk5o9hK2jXk1
WGWTU4xQP6ZaH7ThyEtdjzYPOfiiCnDN6ft5UnMmIt+EgdqbQ6tOfHtX0ZExF1Ow
3Z9OXv+It/dbtDLQz8KPCLge4QLWCJlBLox85RH+SGZc7vaYDFZNKGrgMfK8jEWj
D7qFAVSv7zpV+R05+vJCUSADDEJzEgZ0lsDEWgkVzaTXLH8BAB8GzK3snrezXRRD
Xlk0Yh+lISt51Gb0kfR7o7CEHU9h48W4FZRVv/HHBog4Xw9un89m55ydqc15mGBf
9ZHwJyZyKOsjW6qKyFnchw9lerMzlnGiW3/rhEsAYdtqrCraXMkRPSEZvohpkBjJ
EaYuj0qYPn0IHvg9LSz7CmUJeU73gpxrlyKws9+2KDNiSmz6ZMHsgce3fu5XbO8w
vjDBvSQZb8UNH2XqMekCEAuhFZGIsLu+tabQ+4AqOHbfmpMKWDlobyOeJ1lvtRh4
+OSuxiTcvF3qmJAsoxmVP5EIjgTyjX8my4/CgRrXgVMqnBMY+2r1f247mO+8VRJy
tE2vh5+D57tEBIYqmgxbmLO9p5NCgYZ5Si6vzec8rCHt9U/CmgSCsFqYUlsnZwdn
QipaJKZUSE9Clk7kf+KhJr5NdMOL9o5HC58/VvuJ+EeSQc51jC4R2lRwzH57YKRA
+/u6uKYICNQ1IxXkhAj676EH67AVIbOFKCAot/8ZMnJ8TsCPonlnCbMTc8WDxsYx
H2PWYiAUeYsnj383elZvqesAShmynEz2SSlPMTjPw3pWrQYRfUNWcBdwhbkONUUz
V8qA6HWy5y8h1A3Jd7zfMTghjfXw9akvgrr1yKZxalJE8hdnl+8DDYZFpFAX/un8
ZIDZYVJ7i7RYzvvq1nZYqWY4/ezzID91vb8oCkBOOeIrrcAttypAzpNVT6EbQELo
Wd+TlPVCLHzVySC8eoSuNzybanrUyYGuxLyP0kSSwCkscQRz+tFPKJXBoTYKjJE6
WThBc30qC6DH9xz0tu2DrmXYNBKkdh+sRvquVeMCWjfFHPP89TCFTPJx7jMVcwe9
GG/4raTJpPZVGa62KFJc3mvpjC3oV95p3sO4y4GRAx7sws69UJ3le+9swuWonQAd
4WnByQm1iGmYgK/rU/Va6bhQQmjyMbHucHbltAPAbKZltynhXW6HGgUZIirK8SzE
ipbOTSeUO1KGlIsctvRRUCGLSfo9+f/xr67Ks/q3yq2cNz2zlFszmdrPs3nKj00f
wV/j3/90AyDd2SAmWplbqm4ZUl3sY9Y4NTcBSZ4n4gLrXRxPPStCnOoSh20vQtSi
3ngPckBKHMb/EiJJyWiff9FaxjtikYTEJ+Xqnrj/K9rPamBfyBxXHCIq8MHHOSK1
FZVlhro57CWk/miIg27X+l+SAQGJ/ds3yIRNZ0/eKFyZGnfreBN23ESOqgdGOSpR
hzirGgmGx3EQmRFtvy00tViB2tEN5md9/2VSAY9IJo20pvwgjGjr+5pqybzrXm8S
NnchvBMCJNW46HS1834+gJrGbYoQPcCA2LCJiEyUJ/4O7SMY3hKsHjCVf/tJLOnZ
zLuneUj8WwxVoJj08UI7IxRHpLobabo2MZAwExZkDtiibtPyv6dCvdlCcRFrd1dh
WcgkNXJoIRMzcxsrnL7lMH8UZIoegJqWcId3UorcPIpw1XZ9h25jwh9652p9jc2b
gB6aFIixUejTbLb6kB6WyBEZzVmc6gW9/tZj87qYYaJ7mjMM7Bw969VPoGeUCc0T
PqvNP44Ey720ELy0c9lepnkwu8QeXPD18LlL2oYCMTwTrODCsBHe2s8el1BDIBIg
KjW8rMVAPJPQv0Ix3U9kwcHn2T1HFnJN65JTcUr31QM3hIh/ZB3BM/fC0CmpuIGy
I/B3V2suc9u6SP+WMdNR8lQr7WODC12rLUS8jjyjVkivNExKfLr3HDQZpYqpTRJ1
S/B4Hu4KKUjV3sIlruw+WMlmZGJtycUdTPiehebESS0zitC5HqWOGJzZQddBfKAr
M9gIit8lYXt+fB+4txDiqCNGML6jAa/AhXHl5aqA7PN1N3Ou8UgXGNkf8pUzLyrQ
RQ2WrpTKQCXaPTsdQKMkCFoac/KK9TTl8fFyVzqJBfM2vyJU1B+haleGOzyofLpO
+LegEKF1xNiFLx+qpW35nbz+243Z6zn2ssQrBewaXa1cT2opNbaf6yz8uwwzGdJt
psYflzpUaiKf7agCQb/3ACtfH4tnhMqJTZ4O5nLmZbqvcxSDZpgaTTQgNKRn0tQj
E7IZMscOqwi3erfKrYLBO3BRQk0Kb6CHytj8ZSqnURbK0Taynv5PJO/p1YjgeFQZ
C9rZT41PcNXFrU0iTnb0O+3D/xuwxcXCoc38KCmcy+avZtTI4bPSbyuj107Tc/gF
Xdf/aMQKIbRuTg8rkUUFjNkWrii8zsiFGl/JI4ipg9JEUWb9UXbfY0JsMQ7rq6h+
dxlisSzRS6DHh5tJBex9HQgkRhb6E1k8fHHvF9RWlkskmJRZkoNpPG2tbGxnkXgf
iinANn2Q9m/EiQBeyKcW7OihjE6iJg3LJDODexirIuzeGKkCIP1KcpemZPslMCPg
9TGUONCCbkT1Nqgd8/qvsq4Cd0cSmhryniH5Wou3zdnuQy0MDvnywVS//Rbe3a54
NDM0F+NRBaIKl2c7doA/OF/cf4YLnwWWF9Bt6/aBmsDAR4GqfiwBPfWQX3uieSye
Luk4E45eFirYheMW0Uv7W0bNysr+Ysj0Fx19WJcVoU06da0P4gl/1ujsT+XIQZTE
4D+QOl2JT2rdCtNoi3KwZQfu3y5l7D0p463xKWCD+kqNg5amUgXfJOb20+xhqKJ7
2iIqHE+ffG5V474Uv3AYYQmt5i8Wxif9icvJwD0G3NxzxEFKibiZKxgvgYAhuCgx
5pjQ+yepAyB62BGSh4HtT4thIaar4ftCd7FZY8msYft8Qz90LfygDZx53+cCBdif
2L8/A22scBpT3JCRVS/d01VTpSuPuXa4/ChAWnq5pv0PZmCTatFX6XYaOYq73iiP
3Xoym7rNjcIdrbw0HE9pZdzH0plc2zA/6o3QUT39Z2ti53/DLij3mMh72IXn9oJN
7Euf+ZZoEmDuO5gvT5VljVfjvIzDaWSQOTOvWz+ljt2LYTgq8kiQQ2aRaZiqDRwl
Z24wZS0L4QnsrTsvQ0PzTr9Y9zzwEe8S4ymL27HvyHUK8X4aFb1o5ovNDSyJnVkR
rrHP3Z325QL8qRb95iXSI2qWTabwiNMeFBrc9Fnb4UkQyCD/oF/3TVEM0PxzOp1M
TSR/WZSECPqaT3/2mBO2mSNSjqbOqCZbSZrFPPyZsDHplzw/zs/rjceKmtmGR0p2
bQFcGt4bCEUaGG2AAzKKNxwtfUjQSccuEJUaCyxLqUyxuUnqjddrRZAXKJHw9wro
7Msy4x/pZWKRb5Lrc9bMjnEY+Kta1Y2xHALFP/CxI6/VYQN0Te0OM0elM9v5XKG8
N7K1jTSdSVLRnULdtfndL35Ylo3NL8Av7+TdTQDLWuE86XWmK/THY99/lwH+cMhx
1ciLKXBH5ck5FLqyK5zRPdnlZgAdXB+2hNFNcpTYoKG8poCcfacw+NT8mLCT9Z5q
dnkDKn1yz6huIIvCHkQjeQGTEN2Nqv7JSn1PMEaHuidxI0D6y2tUJx/GYHvuuRQR
a3YjDHkwVQhqzBN0M6UyAyAJON/ROA3LCrStIBhxHNvXOKOCd2n3yQxOZ5jikSac
1UmNkL0KQFFFNxOLfCtTAAZRcp1xytaE93HhQVfk7mferT4fDN/wYMMpDJxbKDL2
w22sBIabwjqgIOxF28yC34f4nGSK7meBF2WDufyDF8axxqLicdU65DGjfEl+1mWx
ts2YGmJNH2Mht16venwKsWpbi3Xu1JKP7xw7Q2Tw5nuOBG86vSMk5CDY7VqGUxBl
h1F8QZtEsrabW75UU9gx+1k4bdp0vgitDEsWmJ61kQQ7f9XriOph7ACY6nWAkoTc
dg8eYRezUE8a/kb3RpJCeX48RqRklyy8DSPcnzsw/YXvGH6jjIu3hhEKZSHE58Vv
pVmoJl2N5hhfMx/ajw0YM9UiDc1QgslUDmWPjtqyacSM2a7kNKAT49wNSp8wXhQ3
S4SJNd76qJmUtpSgIzFkq6mBF1OTJG7KUtaDgR+i/BUXgpgW1Kof8SCds3JUooJM
Oy4vioHUTuCIahmb6nMBCORWOMxDzzWIdoLbO0tnQ/FsfFPx2w7eLR5qnRvbadC/
dw/nW7cSWDI6tQ2KpUm8ikk4wDCO9Pu4H/bgdllvGcYbbxC2PBoFEZOX+P8C5fuq
N5OWM68CUMuRgVH05FHHPQ33Qj0reA3C2pefu+qv2aI6VYnp9LJR5v7BSIhqx97X
`pragma protect end_protected
