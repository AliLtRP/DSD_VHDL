// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
qOcPoWX0DTyofLcexladQ8D+CLIZ8yMlguZvyXqb0EO+nwp3sDlCeX+cgzEsUWqI1RKil4txpdy6
K8V1BEB3VfuqCrcrSSSWgQ8vHXPlzMt/WDjlihWSPeEGGGt1en69XR8NSS+TMetXX0I6fKiRwryb
WmCxlUSg8pQZedg68nGRUiouQ70x+TdyNBoLWkL2iHHAb8sgU3CFI6bpNx0VPpJiusYnd9RkcufC
sjkAA1I1pIVRe65BRE8etKJN+2eJEZGq9eajw+4foER9bgUx0UbJFVsUm/yrrVtRRPCL15d0tcKj
ug5TbKQnLEBNrb0dNdEPLkCzGBaEVrYAaFs7UA==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
/lREOkgiGRlyby9M97zawyvmic1EuDqEAke0mNMNsrhf3rUI4SRjnsBso8WP1YfKvJE8ggm2wMii
d8urMnRaBgODCUhN19qnXX1H1MmsaBwDGSKS3t6DX6jEm3yZZ6NRApt+6FjDhLHt9xojrnihY8V4
b9DeCEZhletAZiGrRmfnX8KVuUe/oRr78Z9/tghP5ICp/L7aepG+4rHnIuGNzgqknjqftv1gpal+
cEXiYjAlo0rJJdxJ/s9QMJYLjK794fSV1QkY2oisIiCGHiLAlWMS/naINTl9aQJttaHXuH056SvN
fMQEDOiIRpn5nuvGqfoghWFYwUe2kUWq2FXMUNyoGb5NOua2NBmaOWiWvbqmADivlaUZhlZ2k+vN
xRUg/1JGDRQ6XQjGa3Ov3wXMdjCfueGFDaUIPDxcNB1bXMe/CK8LaF6Kt++Dk3N06W5YU1ah6Jgr
XqvDzlget7KNvV9CXwp4AL+n88dA70+Z3E1LjZOx5CxAjP74MZGoXvJEoZ1TnSAGB73EO1Av7VVJ
xKEi0HtRupMS+QoX9p/2jaBLk3FK/xkK0mTXgrqsJY2WRdbmNsFrybR9AB7tvidPgVbCDzuu6lWB
54rMP5isG0GsOUgDxmpFAIRrZ8xLbE4PHUBe18GmwBl+LuhnONo1gDSThxzTRHnCVq4ad7eu9aix
+Cz5ItR7nLV2Yv7/XN0nfiq9pYCVvu67ybDq/A4dzBCzGy3JcZJMIAci33br3n6vH28tlzEWyH1D
qY8udbJGAXf7wDyykE/eGOD1jph9xqwn/6MFtmyuY4Ik5fJvb84o0TSilm7xAm9rG+jQYIgYNRjx
2Hbo7Wa288Bp1yj274YwvFYGJ49qDEFQdQs0O4HiXBFb3PNLHjxCFr8++kPKITi3OouuC07Cla7t
4Y8bTPNY6tDvL7pY5x2IFc/MpfHtboQY4Vwx4boxmewdwu+Op9JfZS39QXKg2nrJLOr6NxFP7SY3
m3MeHFuoG7uNO+Zwv/7xjugdCoW7XrcoStjfac4hStlmgzDdVFDnwZHs6201agAKDQ6VOEh8UCV/
oz3BDQnDjP0ZaUHN0jz1kcLYgHhTyyZ5ffL3LMz/La3aCEkJARymFMw17IVWwggf93IOHwpl9HcQ
z9NEDNg0UZKn/OtYEgAH20QEsxiT5RwygaXxYKK8l4j54TyqklBzb2hevmU5mFGzOdD71/Lsl2n6
QbehMOMzxKEw/gx89TQo7tXSMxyfEWNmWg6+p1IELsIMXJrOew7xOu2UNrdKP7yh8ZGCMrh9lv5Y
4t3m11RpTUwKXf3lvR7gdev5kLulVZCFUmkFC2XPCMMsUY0yD07BjZTqgoz1PUZowNfT+8/xKzBP
mGPNIRZtUgvH2H+xVHCf3WuE4mHMI8YEU+Dznf4zkJo7YMelEyHjoTIwgR3GqojpoN74UWw0FYmk
5LiJ5g62dL493YSmbRaklBLgU6AtVCFxQfz4T+LZ9e/Vn4fJWgyWCbBJPSR9WmkbY55uPbwG47Mh
B0xg7z9N3pTNgliVZA4++VIsDD1gyPH/mt/oW0GMMYtDdDcVFzrsWHBcaTcycGRb91YozOm7etHn
cn/D5yXv0XWpnjZQTjloq5FXrQtnHh/k3U5NcBAX8jxjwB98UFsaAIioCKGvj5IjODuWyugUt4QJ
OsEzQHPEw654TG3qtlgkoSXi2w2CNL8Jvjk4Z59mDe/3eB20BkgUJqtIvlRcmho8P+6KVNaEIk2x
LvJHMCSGbPtTLWlOP75ESLIFQ5sTS0r4as4cFANXjtrZO/HZhe+i9Jk9Y0ua57hhTIZ8k8IwNkAE
pgIn00wbO+1YRrstEr9o67IHYm3q5c4A3QuyhH4dva6CRKWogDJCG1ms1GShxcE/WPRvrm2fFZ+W
b7zQn78DODkoP3hJtB6b0ZLQPPxkJh+x5GOoFm4VgI3rtaCXVn+Shbpa1JjfoTCLFbx7uePbo8FG
2ztUkTK0grD1UtnEHqCpwGaAqbSmvBsyaWnGs5nsCq7Dr+l+ZUOfRlREfKjzdjKO5TzSgBXU+Hb0
/cAzF92m75/P4miIAq7bHt+3moJ5/VZ74qBarYWAakbdVA2KFXYq2Fi6yi7fzBms44WpJK/sQL07
B7NV0SG8tYIYfZcClyY37o+E5lXleJQNgvtFjBSxPxCddjwr8IwOwzY9/RraJ+HMs22Z6gVZUndn
sq3TeeyEKG8GHaGpmLj+XKFSBJ1DCsi2XiOsLrO8B+VQ7uIXKf30pBbUN0bUz3Nfg45Cba5Q1NPZ
MiKyOOB8oC3yE2UmBS3jqrKWDZsvWrgxTEA1GZ+tX8jO0amM3vD7HsywuzstCayn2uKa+eMSqVZj
MyRt34em93V7xqrScahiPFWLt2B4JrGY7+soQt8fuZ9oFnJlJrZuMjS0hVwyM+w1oepZMnDmE+Ss
NCSpjBI+N4aWIihl1g5uPD0chYzpRIMm6rYe3iCxiyYhLflIX+NTLHJojx5t0SQiz2DJuRP78jKg
cpVFbLtNUqW17xR9/jxymnMh/wuxxgWYzE8qawzzEslrhRbUQJwxhJOeuhfzvFYLYrrIdxm4BM6i
7vIR41YYr8eTL4m71af0tfHCMcgb6smGQVfz4o9OXpRLLbIJKQ9pRx7zOONcuW6kenNwnucfKR1u
4HTITKyVXun/4VU5XDcumtH7Ul22NYi++CyTWsqnzZBIN6VHaL0LISaHl/KDtN6P5WWCKsP/ylaR
9ohIhMafw67DjeL1XNdNKdORYgobqcPykzE8+7Fp+6DLnH4yGh1+zicSwuOifV2bxetoQFKxQHaW
VuDmJUV+sqmMEHSy9hFgwlP8YvSJAIWIWHArxwPvY5jlkYJzk7xZerlWZRcyULf4jFQWqYN8LS2x
Pmmouo8VdBTikp1yxJL6OqDOCQRcesM8q7EdP2R39x7NF3YUszBEt+TKlMqJEFouW1ucWq3KQE1D
rYskQCdaBJ0VkbCL4MsMpT9jhxH35GIpS8/A+puDj9cN6hYTG45o8I1cZkzPduLOLlwAb2oOhtPF
/ZoS63rpHTl3iApAEcAHUKE0JuvPDBHlRH59wM6Ea/HKkUGu7J4BOUuKMUyQE0YoS1RIsgpj7m5q
eF1RSgCE4j+dxnXuqmCJDzNcs6iYXOExU3DrOy/AMK3SFwmHkkZ/d+mL0iehTwd/AC9uMV7qo3I6
8VqrZ0eq74iIAJnShMXmrlMRVbq/x1oLPE6lFBo5A5Aup1tPYE0r3qFw2drphu0tYiAKcNjzHeaV
4dMgamYyBwZYMZajshgMqpaT4iPX8bqo716n/7MA6DJkXXW5ObJfHUMVYJMpsQx4k6Z+UfwwNm8h
gLoWNphD0VKimMccYopTMkREEL8YT0oAQIbpUbeBpVRA+Bz5tH6+kv/rDL/pb/iwi68w7rzTGmx0
KBG2dCUR//bE8HHeiw0JtFLk1IioegF8nQaGeGue+z5LD556mRy8IsQQoXx7L2+EApiQ8VYtrNaY
XiQpvpowbG48yZ9tkNlB2yyXvX1DzZQavu73ZQNyED94AwEuOXQqkSOVRbz/AWT9TfDU3OyBF9ni
9KkLyd/u+xBnKVc5yUwZWjwZOnA0JXumoDpmRpoPunOh/IvS+wNeBldt9vI9GoGa2VXsdjVpFESf
6PrQ84sqlJS6fze2Sm+nIOA7MqPvdg7xTpFDQMUkGEWEu2e+r3L7B0ReEsJFRXw3HQGF1x6i57Rh
Y4R/YAhxKrixi6cUztE7lUVsqQgWqwmgZilsirxaBzD6JHQmkeddREqf4CZ8zLDlZ2bkhnmKOwVg
XB06X1qdCz2nvSbKPMvUo9C6/0zG24zaHbFbdSiIYmmZTKS/2qGl/VxProf3PiwSixo2alZdTfzF
4ivNjx49QrK2xij1czYMy0O4Rja/lml5Wd5lYcj6q2PrVLjYvBG57tjyxW+1T/twKjc+w+LPxNgQ
zPN37mKMUHSrmN/SW34sgoJb8bgMfoGwNsIBZXso3SZm0N/dhI2xfOKyRoL6IJ+RlUVFB9O2uwDR
jmc8Jb4BdNal72hB5YwO3ldrpX8zkw0o1lnLQj51+NnrloKF67ofG0tW7sFtVXgna1i7Mbs5n5ML
KB9CPuPMxnFyMb7eS6biyXnXJ1lDuFsPDCZi4PwwPFvZJg4TF0ppdVc1BROm30vVrbnE8nSfLIga
ARZB7xuKJiO7GUtNAL3xcCm/o5oGWakFWidxpzotf4cIS1iov6+1kPNRYzcni0B3tSOkkB6id01v
qZRgIR/yqGBbJwSNMtDl+6pu47k33Tgp61b7Js5D+DwzANGod0K7SYJIzfOGRHQcXUjqmFSui98L
8fmbaE0jS1loPmUYojgbuS04oJrDJWI08dJUWNz4NkMNBvOQ/hrnl1G9E0OqBp2YB3QwBToFL6EA
5rHZPqguxgmvVnY1p/EiN0U+GBnTrtONMFLVOWnMNrpARMIfz5YcNapXL33cmCUKq06SXA/53jaL
NIvLgsfHf7leMnCgFiryDFve+LCShnofqvDD7WROVX3tWmbOPN+8qZo7AemhbY8FXDcujQIhloRk
KHwZXDWvo5ZKVR0YO7Q2a/1CIEBRi2yuN4tCA8Oben4UCCD65xMdUEO3xAbJmmcwg9GWXhrdWwWr
KoNfTD/xfgSphPgboI6GbFb/RM+b0mH3VN8ntxFZmjBLN3iIDyPwB90QzdCml1xbQhxj7egtBeOe
085RCoBDT2s3yHWiK/bqj5ml3Ks9Mi9pHTQF3YWDHAviHgstE6x2iwkDqHg/rhMEVcq1CuVYLbTW
/3yoJYr+Uy5D4jnlMHvR7cMyEeTVQwmtYV2vcVHu8cZjUzcNYuz1DJBgSRhKPVVgExgsUfTgkUPU
t75OYVofSffy0fGjCrjE4hEGiGEB+I3K0nAeDTqDHkT2WBGqisolL8Tdij/CrL3D6YBOaYRXWUcJ
PglEC8wNlNsGnyOt4EWkYb8oAVeQMxnEFQ4x8XwfLsyE0XMTpXS+/vqTiYyr8fegjTDK7hyEfMAX
G5RwaBoq8B0CMHJg2sZlxNrrC7b42U+eXhtst1f3XTRjq+eq8Vo1LWT0admKl1UTo+AHcjgbJdky
sDIaQBS5Ib8fv+IJTLwTcEirW1FJpW7q3CPfwggvFdfX+zJnJYHJU/MXItAQDy2jCRorz0km54Ei
xtYSto3DLTzoULDP9EsyNX2lwmaoPA8KDvNy6uKayW18jXre7MOxPo41a183GlIACIOA8SmtMLvk
trjBgLl3u1FWDU3O1RCSOyyzb0RprXAqxGsJAsRxmIYBlHzdzexUPmwG/J5Ny6Scr23N3WM42ffV
PmvZd431ddvB0TfiOQ39+9RtMEnfIZlGhOHoupLFsHcHNqpLaiYaUeNoTkHUOhP2ULa4LvwpujTL
ZfC385WtlfjFPN5WSfpH0/606xGjRB16XeS/6Lsr1LN7Dzm3akVwelVwihmEyLxp0/PQZHId6KGs
gX9J/mWCnjjxRNlhWoVSsHKTPk6rSG2HY2ZHtEWkS85vWrLuzjOWFf/xG9IXA4wMXxcmmBoSiYwJ
EI7OKPwZwf2kS/OHPfQR+7pQrrO0xC8DNdQVMPwmLgTm6m4V7Yb4k3403435NQkPejI/crgCqFkQ
DQmJUr4W5QNCe0ILne4Udy7kUCfXT4ylCwEAorAz0wPlW+aREpbIWC2jwvF029fD01NMaBgOly14
18zFUpT6WrOxBC7Kpeg+48R7aCWsjNaEaeuimhp5G+B3pHLEAX4AlCR4/YfE3p7kjngsZIc0N+n5
B+rENeqVaV0t0m1FdbgaZXWtz0Q/TPZ5O5Hrt0JIZlWRRedk6JrGHofGkAiZEauVKwonR5bD2US8
KHhJVibVp8mP9ppoTRyqogpZi8d2yLejSoUZEG6JjrgJwudNDYGrKpxHR7xHi9Q/7zc44+rnGLi1
ctEawGwzbShz6hwBO+CTVbUpK7x7DGGqpSzd+uO3sOE8bSAjAuctcVvAuwh1azbS5NuzQufHHbeK
2hFsmm/Fic2E9sImJq9LIkMW8o5Xd8q7NAY29AhOYYUKuhXeBP9ZQxFBPHhu6eM0kVAqOOAKXGWX
wY7Gxjxcy6TGyY2eHtIp5IXx5aey5TPT2b7xoIq9R7JciRl9m6X00H3lm7lhrno63vKHV6t4TmMv
pSklqTaUNnksp54k7z2wuTe/V+nFTwYnJR7M//cMuuPgG1OB83T66nkAR/FDWyz1j1ZRfftPiP9h
ZQoPqIGNNysjIQLpEsC04T8QIsgp6zTx9veKVZg3YNxIVEHc7iFWDRKQ/LlnztQTdBJpODfYpQh6
jjgv1FYLZbNVIau7LRa6qJyaRWIafHyQs99xqiFRE/gV++0CwHhtQxsOoif7lgGb3Zy/0U5cA2mI
rxdm3tw8ivxjMQ2+KFyYQHkau4RE4GEPkLi6wsN699lLA7+AKcklNtgeVh6pcbumyWrmY1JP0Zm3
rIEBUlCuCEDSZL4c2h0XVSK7ALRt9HF3KYh9mB6nlScJGQUlx2lJHkjYlDNiqbcWd+9IUqXxkIQX
x8Xt2LkfeHvYfbBRvrmmAHVH9TgX8SWOig7CvlGf8++z66seZO3lbioOH7c8rLLxrUDyXwc2KBHp
WPMwwHnMxZFNzdlForV25RZThE7Bsil/405SASoMJsmcyJh9sqxY2OroJ7smBrfW5mf9mxAhTogI
R7Dl5x99G1acyjJa2RN3tWf/CKqRpIVoz5jcNNPsbnHFgPlxJWlTSysLgDuLnnwELRukAaAkBAqL
5Zv346zMPjoYRfKKRPwQi0+Xrd7XgP3ENHuxP+zU1lw6JU/rvbz2vRNhgKHzj67BWkrL4FxCaBXk
PIVmAyJPUR2Gl3+T9zcGz5Mi5CTUW4zNzz62aDqKpqgdr+H7RQs4aB6BL2Y5bf31GzChWem1w2oC
CPN9bPPwFglmNXVD1dMJxTtBLRyvOwVu1/61/6K2evSJY1+3vCX6/yUmUTsIAo77mLXKoBYNo0P2
i40iRp7kh0YsCMtc1TrYoi7P14XpHRKapSFYE93gW1urALA7y5u4uoeRxXEJVbLkfwJXkAaHauaB
y5PWLPmEi3kcvxNbqp2MgMnHfHjf9cL7GldNLzkOQdlniciyfo9WoR2MlBLhTI6lcuLZfLsEBM58
Se5TV4F8yvcI58HpxbgjYvajfVR+yBaeTtJW6z8+bfsT1U9zA95CyP2zZ1R3DmmI0X2UokcHWghD
jcF3rpLt33pw4XKu0rxl05TX6/5yHTe7aSBzi9GpDVMHQLIk5Hls7lOlaRrSLZcxgSX+2CG/MBQG
499pLSdtRE0zrKRTAoBjYbU5pa8NhUcHjATj8vCl85OYjZCVORUF9mA4kT/Kl/35Xpx88SYP0E63
ukyPHSEfBr0wmX6Zh38Zh8FgsemKSjp5DycpgjBW7lLEVXwUrPSWym20kEEklDJ6YFsh03OySpDG
cXWW1wpkXAwySb5gmDgIGX2qEhoEuZ55BrzgJypdzbopdsTgSuGqOX/QwpHqs/kX5Uq14oingF2v
LIDYulJs3U04nMRGAzrDsRpszPVXL6lDksM1BDYL09QkSL+VVNt/jSqydfesoyJ5BxydWkobm4/y
1VFJBXslUwLnqSBWZR2/d5Sqrtc/1QZCPKx6HqEYkFRJeRXz8wBGQsQkhPrdpykePPRasD5QehTk
pRAeOKpLxpoJpoc6PaR/LdQbYsd2B80zEGnKWb3rjt8ByMHlCxfKIBKs9p64BweghDsELg6i1oQH
2CpOb+Yn5LNo2/DW5q4znxg7+hrYkFiERgLDN6c9EzmDW3G97TSZ3RFsurPeSIWb8NAsLR7eLXWy
+PWFLpS67HGGFeu2+ppWkcFvM3u0eqRohjCeAe142qxJNYrbDiVdS7KTHK0BZHhlzfM7T1/jt4j5
cD00HGivdnT0C8KR2fgumAqawJvj7Hv2j4qmbc3v5NArcS+XIv6jntaso7B6JKniNwphlVW4jIPd
9eCCG3zbhn9Eh64+iFhRk/SJdgVRfswfoOW2rUe7OMoLkayKApuGn39HkSMIM3RL2KJ3cO1nXOwe
ndeDQX/Xno/49Nc95eDl4/X4aZpIogY+hvAojfsLzOSAaC1Q7n8Y/9YfXD8pnuMi3b93eGfFrFEG
ncP3BCxY/G6X+Pss+wHgRNOM5z7KJcU0IEvFS0OG6fYmS8RoRdkNroWgdH13C5BCE6QlFag7kexA
7IT+bmk3/eaaOwsFGXRphh7Lv6mVqzJUHfyGfKvzeINZ8SjvYX0gEVTnIO7P2EYQF5ImDE9MjRWE
QAZ4d1ECN4G61NEEwUnc0X1oEzOK/iQs9W8LsnTnPvwcW/C8Abp9MZoaQd2QhCmW5uecXgj89afc
6ImpBJy0EIwbqbb+oK2/SxldCzP97zZ07jVB25uxUYy9Dm2YZ4Ejj/LgRqz5X0rdZ8lWo83e5kRO
o7T/5X7uCVy7yiiu7pLZM/wyHJ27LcZggbeBov9VOqa1NiU1DxrSgezXhoklbjY6NDsJDVPtV0o8
dWMYD75mm4JCu6IgDKXFrLewqMICf2hTh9M+sZjSahqy/JqBcKJ7Qh1PzeTbROmSPea9IMiM8hf3
Tp04PUXz7EPWj+m7amYJhVqr6DTpb0esjYSjzK5rkMFI+UWFT4rm5+LfjxrKMDJebky1wTWZ11cT
z3ml3jBDlaRFXylMo6YWqYFzas/h/Wx2YVcXvJonuOrDmIIheZWruSuZCPHa+A7KMa+F57INMmGS
sdkLP7XvOskjt/hkgcCZNptGdgAXYqKz41MwMtUWgoFuPidk4ner0EinjX7ojUkHeR2l8Efc0Z4I
LIzXAnUHLiFhL06ONGJWAIBp0YdrTThLkzmp1qPQGGf3Yg4G2F9eDKQTJNDoxhSgpVF5I1sTdgXA
LG+QDNxRg6CIEz2lx0r/m2r9MjaMhsGz65WkkFC8DnPQz+cXbVxglyQ0YTCbr3JHy3EEjTTCeQWQ
YgccPKzdchcEknDebPtxMKMLS2QwCZi2Dp6TN8bCwnXWVKlEtmziPRDC/F81gkmRxyTc/WekUDia
zv2IhgNP6eipWO2HfaTZirPgGxl0Sb2XK1W9Y4ITrxo6Q7mnX1MDpdKV1pG2utNYCqY7UkVV/Ifc
TXEZY7jQjE3SozglPTKqIlgsSGjaxJedyWwRwjBlFLs+h2+G92jTH8rl59zhC7ax/s7lK8sz65Xe
TXMwWwzlPLDFbnQAkrwnLKS4yoA5rqaLsAY58RRyJtH8jN34RZk4SL62SrZKG3+AHFGDjNm7vV0p
mCVzmfdsGm7E/q1MtCRVXyHitoVZUkwNSW0ykBxk7PK7pv/0TAj2OVoHcxsEWi2G2rG2PsEKwV8+
fWFQ3S9P1hM7mwf1nG6hB8Iaewlmwftzp6gsd3YlxBeJvgFZh72QUyMB/HOet6sHmED1gCvYvgYz
wrMRnPKClOMaOZenK1s2OTZDdN1EcNL1dywMOPvOKQ0MPJso3xRslcY4C4MCLVmA2fFRgn91IbzX
o67rTK65QmPZzoDCKH+75y8x/0kgWYJfWVOB+j0A+lC9vmLJ5rvSr5HJ+ESAL6VrwJ922lYK3fOq
X54l0BRniAnK6YwsAHawNc6thYMio2+kWnMLgIU5cj57Aj3UqvRAQTXd3UXUF+MA+2U4wrYGtZh6
igcEjefUtaZijKwuVOyjf9ILFw0m9IJLeXwLwbRjs/GvuSpboBakewmISx7lpa37FhCixjtOuKlk
EXxasvrMdDoPj+qKgeL2NUGHd/No3C/lNapAHNZvod9RtF353mF9Rji1og54o7y2ac+1NR1LhzMd
M/8mfKy2RwbMzYG+NKIrPzZEeHZ/st3vfpTDvIoQn4tj8qLHeCcAhcbwUwhCUdqCMw2c4QG+5fF3
eyqEp2MCIcjnlCInoiwjCl18g1nGld7DSdQ2wWgXC+n5Ioj4reol94GdK2aNShFM6Orgh7GaSbyp
p17mlVGqRNQHOCb31iu3jc5kvZDkHyE4ziK38jIHam9iWjfEOKJ+1yxM98G89mpg2AiO6j4lL4Og
ljdf1cYCrdth400usPsrI4zfcKtBvhCdTi7F9JQcaESpu2vzUftrO/01QLncm3CR8lAmqmcES6+u
cbZEGxM0LiOEhZEWPH6wjm1kqrlgmv+BVWeTSdDLIiMi0Nr2QG2/TqlGfOdbfctFYKjtSRtqYr27
4zUgD8f56V+JJbh+eT2M4dqGerwVL8Z77jLtATz9U290WCdHM2fUqHGTAKKREQwGbnZ+N/bTSzgn
CG2LmQVWbA3lKK/I8uCsVph1xW/t+AM4DTWhkSR5UyDF4qFL/ID0TgYNWNrcaqVsH0D9RRs2xuwu
KZ0GkLjThYfiC40rCPQEhtZv2y6c9Qd9vurIKyxEW0aezHAFeImz+PGLhbVNeJ0XRy9x6kcjauTL
G6F3fFjHwQRaLSRn3Nq1Qdxw4A+H1qMN4pMuy0qkBMJvk/qwO9VGaSbsLq2IgQn/QIHib9kPb6rz
DN/ND3DWgvbCkDi5UDJslvg2b52QUe1bAxQCgnidLwFlov3DNkvZy/9SKF3/MxUYoRKSExeYdWx4
c/sasasNpKvdRghZkQ==
`pragma protect end_protected
