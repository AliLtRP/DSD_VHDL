// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:37:18 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
D1nNO8W3aFI+PjlkWLYspSH6+GrtU8x2FG3pa22GwQTxciZan/cOUs7Iponw4eKp
nPZSBBNW5VydcRS8d0Ium98JFdSqAW+6H3RbPtQFJQ5900JM4KTXENi8GwFGfyV7
zvMFvuaQy/VbDKjKC9tXlYuXPrklG3+wHOF6esxRxmk=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 16560)
LBZnRonaXzcoSzVV6KsfMNWwVzq26eTvEBoyCBw0BUQsA6KlaXUPAFBqeZqnGBpl
GnyomWOQM4IvOe0B94kRxzhO6iARJuh6QZgRNKEP2lUwH/jxyy90ceQ7/kDhdWd5
QJd1dyaPBd87WVyMeh5CCAjLipSR2tC+AaZzumPDMK49jPJCkV4FRpRUbQuJlpE1
nnYsy92OuIbQcc/EGE6nK7R6TRwKUPaJdygxeOY6PqiwSTl77ERyX6JUqGkQ3lJn
8dfVGP9fnGpb9kw1KF4WyynpEX6jCBBgxY4FybyURhfxqnTUnNavvy6Wzr2Ai6uz
I5/cgmUoObDRTHt16/4ek/6si4WLYFXk8Tjxd+RIV+euvZLHKfS5f1CuyfxE7O6D
BSApCZ7k6MGxabP/QacyWMfhrc09+SV2vBjVuaW5MsW+SxV9sA3EV3aVxllUv5vK
gYsR3gwg78qXxMAsVlfUCDuXxx1D8ZBxiQ7oTwJVNQjhx96PSuS/avibAy/CO0pw
mG9mPo3zsObgM6V4c+uROMl8TUDVkQlJBNDOBoLy60WemtzZqjKQxGogmmrGF6oP
CM/mU8/xZw+QyWOElQv33w0dak59TgVaFVUjaDc/zq68+P+MZdwNvd552UzlmJZ9
6S0JGb1laCImsgfiWPAEx2ohBEg8TxmhsbNxLNPP3nodT64lYPybsc/Znq4f7pB4
2o6z2IfDm5RxOSOj8WnI+WoQNAIjBNmiVRni6YK0LwdNDJ7iri9YazWWKiw4oMIK
6GLYVq3sWXr8XFobF5o35nGpAJNN3hXeAYWm3KLD9fWZGjgtd+azHVp7dUsou9eW
F1J02X1rK3wTTMYbfpAFmEDc9aChycSEqvHtdniz0nH0l5dmAoK2Q/ouz8Ro5YSE
qMrmqyhlMGrsBJYUwaKBjcjj+L0Gf2halhSzNuI8aqUJWq2eSBSWbDycSqIFK09F
XgiQ7YlqSx3Cp0IJbQsM4C/ikiBap+7MrTjbaRr9D5t8GUmIwT0N/bp0cUYuCSrr
OSpXdHzWr5L2MGLUsCbxJz2FDOXmOZJhvjj5Pg8e+DO6q6HzcDWTKk/OArHKlS+C
gbc5jOmGNOBzLmTxV3QSJaCa3J1vfANRK505HPjxFGw4LxV/B+7qbksFqK47n5qR
QPQWqSwZ030LWm9S9yWh7BP580t/YBKMmg6+b8uevm+ulXQDkT2jAaHR0ILxx8nY
ViiyY0rRxSih29oURd3iZW5aSVGC1dh7RmDxhqg53DyB6NoPSTyzrx/8u72DodNS
CwG+9HCB4RcabcdfB56gNMpvbn+9lIMgIiRSEW9s1fjp6Cv+W4DcEQt0H2Zi1t0A
WR1tJjgmc6SAS225TzLWAqhejlCfszJxDupPfoK0shzTu0PClsCUMSyWWZRMysaZ
nD7nJ9SuGhhnLLlrvE9WKPVOB5YRhl5WUQNq4RZloE0BEQ7RaWQ0xZPSMkhdQRrm
anDJyqguRBGEkp08x8jSYBhvrQoDOSzONJXCnRi9KaGCnUjmj+S7z8iTmENK5Nzf
FloCtihNDmqcsWUb77eDARHTWfbvG2NAYRcMJICOp8h2awKWaHObfqh08fKwj1V4
1qqiRNn80Pw1U5TVOhf7MiqxdZrxwN5YZgrQUMq8/X9fZuFM8wKgkiMCXIp3jEy5
6Zzwr+vwh31Dzbv6ky2ibojZrBOeUubwKrn99F8nMwEVjEF1WqcWB1t+2pkgUDjc
S110mY5GTIsdwOF0eL45oSOUcxBltczQmISCWU0EtDoC7Z9BDfHf+iH2eU2/ebB1
/34OA+iIYZX2aDZ7h2YX/fJDNoiqn4qVSK5UUnxq7PbWWvqliyxixRCc4PlhiOuN
TZ5Yb/7cK8al4E86NyPQLsfTrAZtcHu0t+uzD47RVLZ6aztqz6w5GoZb9ITH53Bw
Qrcn7eB4ezzQ+L0sPWySYshIWM9X2OA8dPOqJYEytFiOD59MY0SM2NbO64wdB4UY
QZwqZhoFzWoSjFmbibA07U61YVd1H8ZTugr4qSbGtEdBMNyqh5Xl3JSZu9fXUIF6
BwANfmh99wHf/OXdseYkjjQb5KlgVHUuKCK1LrOTeNLLsZ619eaQXIx/tYQb321q
yEIueMtLNjw7/rhhRhRpU5WSY0Gp3zHOtuZRS71VIAYcwRpuMkyKYBnoZScp8+3R
BadavIPOQ1M6mAw+7Vql1av+HN4LrgOemysc8mt8+T/jIyLrduBvkVRkAIrBlABr
cX7arBVlZ+PN30d2M08R9lf+5Yo46qNEy0F66pPFY3pVLiB21Z1Mo0agBkODa98p
R2SZ6xZT2LsnFIcOG/v9lxPR9vwVdZ65/3P/DKz5Y/7PeGIlRsxjjw3niAsOnRu3
DGymD0KFzRFhUtlm6GsHTTIln17oKMmMF4GWz3V/yUOTx37EMKY8j1z+DcZUmZV1
Cd0IWXnaQo4wNb9uDOcoziXWKa+u7yeGh1hDVczcBs2QAG2RVWz5H1VkYcv2rJrt
XhG2Ad9xFBXsJdW94wS/1+pdiZ0I5+jeRpbFN8ysqU7mADXCUJQ16Op60UF5zZEc
FISbskDT2BL8DglsRU98CzGeQq1b//4ihZruBfSVvMezu4f9vlTv397ogOwNxwx5
N85f7KVyhN5ikRu9p7uM2cgOlQAUPc1xkzQa3EY7SJkpkMEGWWnCQGMe4AKDteNs
F69QyM3zb3KqPB9QXKNsirFRyo00nIvGw/94DEugTjVPZ8i89qOtOeC+Hyk7l2lT
bEH/WrlSYdX0e3slE/++gFSiXrubk5AuAPZfybklm4UXEfBSS/NJ30oLh3VNUixy
YkTtDOr3VRXfKiqGvjGwNxYCH6s6eel4hhIuEJEwovOr6ocshDLzS83L9uKVNrfc
Rm1v3UzltkG1tuXFSFORuAbtaeIS8I2xfcKGA8vuMC3P5k+AtyeBTp0taVVc6qc1
juOIBTKsYhdXupdog7Vj7VTsB4/WUKgRKyA5wRkl6+JOetM5qUHtUDUXwVy5MBi/
cpWX0DeTkLGV2tC1A0uHV1JHvb8jMhQxxAmmDtTzkYUmxWYHMJnl6clXqOqdeQV/
/I3yexdaU28y5Im62oWI4hLgaBkr1wzhHdvnwQ9jh1n8gLNMaH229jqA6wwL/2tZ
zyTSu037qkeByEu5kgmD4QobO1R5k/rigSMtxam1si7DdU7ktnV22BzSqCsM6DsI
QJ7DiNpPoJPoGj8w161sX6sokLf/GfwENP3ahqd4JD34p21P2XaYIrnsdB6Axask
zyQm8M6G7er/xh6UqED+sz8XiVlnz07u24J9uTTTaRfOcw/D9gltffUOaGKJWvb4
goV3CLCi3+aBrhSMVKdJtEnTi6SBZ6HUzfc7OQPHqx9x3FTJXy3BRNi5nmOq28Rv
pnGh66efbfV2y6H/nI2Oyq3r9qVfBww+ctNkV82NdZJMY0tWq8FkfWKUIKqH1gF1
LAyP5P5JA6tLIhqQGpuaIvrA3taNkDcSLcZkenXdsLHQm99P/1md7MFefAagZrI9
4TwlzUcu8uPGD/e6DsUNAwx/FzceH0WUIoTkQI2co7VCYN2qo9g8KbiX5/g9u+Tp
Q4HPU5UUooqZaYF9S0fzNcKxNO4+b+jRfkWm2L6h81MjSdfDWB2G3Fdxlowjwhtc
mB6Qyloi/ptlIQZgFXYGLXx77k0HMJhmPvTH7O71TCZLfhExIDyspefy0N2umtz/
bWDuW3tsQcWNUlaUdm7yy2uE/vAszSF1T0KjkAQTrQAOwe9TTP7jhSIEA2gUDil6
cRi5cmX5GaFMlNmaNPlAauSskJ2S9KMbL3TUHMnZtCEjSryiXziwfjtIljdvLAAn
LmZnPhcd1ZD20cemPrO83zxu6k3EvbLYLZlEXRPU8obEAqkald8a2EGZQad2cR/J
dC7RhpcLpeFpVbic7CC16YoeqWs2I9vGlsxCEja20mvV11kOJp+l4ZjrFtptxOnF
Nlj4lzTi5y6PUQQFevM0OkyEMt747khXkCP5w5mXOQssFNxIHhlHgDm93m73zrLE
/l9zNicXp5S17UxOLU7bU/Rn2OXddSf0x20qFhLwK88aL9hnVfz80K/ct1WjCjtd
rq4LC8wa5eoNPWTyE/GflG4RF++P8a20kYtRLijczrxgqrrpigU9HCRBGrYM72J0
oR6nzFOmf8/m3veq9YlwWi9e2b+RHmd49nTCHd1V1/oKBODFUJk3YIjEBWP2CPX6
Ek45cMkOZvTtovc7CvDhzpx6O+P+//FqvkXer5F8xVkYvgq8/M9VH7KArxuZe2bl
EhYBYSlcuf9KDCUBfLOMggGQ2XrUIAjnYGCLHiVmH+QiS9nrLZ16OeDD5hEZ6MFH
4t/RtRGVpKD7iNb81kZNrSuq1MHJ/WKojoNuSHQ8a+Opg/DQVNBfS4dLOsulo+IE
pMxr2eGcrTJGoUvxa5ykGhZ8pLtnEomnnHGJMaoNSqBobZIWpBZXUtFEn0b444OB
Sa41McuCSoE+rKd/TOnf6Wd783e+IbDLT3Nc1Qjv9/o2I2WYWyCr2FYuQHhuVdvD
RM7euX6WMqfNARdLi1VDpRcoA2k9nMajBNtkx5tidWwg0gNvWUteWLDNPPerHW43
5NY2MTIjB/g+tKC4fyb/WjyPo/e/iyPl4BUwZUCJPGxVmr30Rh3sG6R1VOJNqH8i
zfGmeIH8aEXD574MpOuhcoltxALo7E6+LGNrlA26emtmxHDx6hE2xM4AIp/HZZPU
9lQukSDs8XtEzkyPwM1Gs6YrEb8OlPWHHCRuPnk23d0upqrlZsWWpqrxrnK8smWa
kqi0CR75zu3/hG4THtVov7eO2uty+GcQW7c4802Od0HNXRM7CLfucu2MtepAG+3W
Q4EQtffoNjv1IfKPBwryPeNal6Cay3J0R0vng/Zf4GrR6qjn1bgYqQ5CSbawCKMr
BuW430Rs2lPTWc1YlqgyYmYAmVOd8X8LZLN4F1TjT6iKb1UkprbRIZyzIIsXLxpY
P/2yns4fmDkRwTFUO4j9MeuN8hp/MxOpgYjXKZBQ/kRpd+sjxxifQlhghtSVyLi3
AFJSCwT8jF6yplBVqiaBXNuXt6oRHjuZKglyRYA2J0M7oaToafS708/jpae/e4V1
GpxrhfPnK+ZIR4JFNzrVu5heXYYyq+Cg62LNZkId3BrKAf/cq6Ocd5EJDTFXcoss
XlBSxcn6esrbmzCFRpDgaZiSzfrEUjcqq28LdxVDJhaXwtN7+Z1+IBINjvUGfG9a
a6W8V9kxycj3qZH4rVJPpfHcjs8NYHeykRTa7LLx0I2Hm2C88c4awmO+gvNxU1nQ
OPDw31EFlgTheUeYdeSD9Y/6+mTEW1OxYXxLe/8uneNS2XY1rjJMMNL7W3V7857T
UWVVKchoUQ0InjeqRFIaXyie3WIDYw/VyrQHkVimixCRSpN8QkZs4CG3cnn9OI2s
ifT/YHkJ/Ni5wDdBZ8AasG8ThmYOC3I9ADtF0CZJYJ7eyPSoRqh+cVcD45r8ECjA
+vuV+w8Z3+A7LhF9+WrxgrKoACBGokw7FTB5w4PznRtKwDmHgckZoe/oU/+2gPWn
1HBk0HfSYtTSm6Z8e4FVNYFasrAssz85Ye57J4NV5kZauNxOILD5/nA0M7nxP6O0
glWje5xA6LUPh0aNE/Gegk4WG1kMo3CtTQeeosFZBCXgEGUVAAmh+s6c5K88TN53
jN0KiUUKYMkIWm8uUUp/w3KMXeP1eRgftW3y7C7rNaCPs5FMj5tf9an/AYu81Bez
LFLmxXAYrhmOOWxfOiapKfGruUCgm46Bu9xG8dhq4ANfXgTwGZdd+O44RR+429bd
l9Jy/uEjc+hjTE92rtvvZwtHq0abstSLLfPAty+BTs88QEWSeri0rrhsCKt/yfCq
MuzvgvHdNeQ339yZ1W/C+qZFK3B+XlXmWEnjKALYSn1Sgd8gMZVzFxO1NTBEDHkI
MnmrDBcmtqVFdMqr18je8BITb17gV7oz62sZMw1x6mTASTcBxHQej+PbFToZK759
/sr6wJ58mw3CKrcCYHxa0x9bOq4UbYgb6xpIhRatOfdU96nxbRmNCzCvRFDUEFEB
Qmti5gFNfZm6iSXLSamvdSitOV+gJ3AafEbPq5mkntE1mp0bi7tv0PRoninShTW6
xaUw0s1h0S6P1b1GhWX2u4O3EHoqe/gL5NHBJKtE4KuTq3RmMOlaJ1pOS2dy20ND
nZiZD0OaI0L8s+Fn41+7yTuX1IeDamd7LyJ4gr8NeUAAqYwmY/G/BrrL8yK3QvCU
yFgOrf+tmgbqYAQ3HjP0jQNl9zUH85C3sCh16oKmi8hPtW9XFHUT3EXRfMaTorTQ
i2zQidDAk8H515TTqHxnqZJO6vyw3J52cxo+QjMvAAGbToYpqiGlQzW9kS5ileNx
KY9IltvhdoGV6Ic32EgwFgbTsyFHV9GPycbB1SXXMMslwM5A7ZMgQy95xfO+zd16
qa//XeEQacbGKmrRFNgzOWybrE1/zDihe4UTDxegEW6z9rx690tZnwdtBwCZw5hb
bJRb21d7Oope+V3prOowDN6U2K1uoxjTEl7TXlGzlY/Y/v/Eh0hIzHTjNtxpjYOC
BZ6rTEYU4+0ZaiovI73khjfl/g5PsupppJSG/NfcbxJe0DxcvmE7vEwCZDrJVI/a
5V0vT77qnVe7aFJd5KiAT24Bz0/BLB/8hvpQtynT6MRIO72e+DpCTVyp21wBMymL
tha1cVdxB+tbQ73OU/jM21yMrJGSE84eKAAC0IBh7UHTzCWHkELuHrru69bDPYD5
i0svZzf8XvnRB1np9lwBhO5QVyatV3pz21yj8EmNzM3w1z5XwyFJ+I3TfC+NKrP7
vly0hV+WFjLBlMOFzvmgujOEkslFuGkug6DKcm1bS3w8yUQ5wFtjxBEKzZCP2TO6
WCXXUpZwNfX/2HCqqCu5b+47pPgsOv7/dAiU3SwzrjPEBAEgxEYWAkV7lY4HB4si
x1kwgOz34ZtwIom9AaKc9LbBgALXrj81aE482O3HjMmAh9No/zDx0KtBD8JtT7xF
nWZj/DUFvqJv1ZDF5etQXHsxOrRF1S+g2PJGvvmRCemGaRmHBX+OW13mqVIn4yXF
/u3jMUW2GayYIuTHPtBImLFVzm32ZNLvDUa0b9aFAPf2KWMXGTiAFBU9U6WrEK/i
/x9/TuULoBBdh+q4gaJz1ki78WuD+88Wskak1mEt5qpPNfvvwsTiQKDZsc6XJdGH
5I8dBOzw9qv9oJpioR9XJC8pDc0ga5Dkn0tApQaucD2We6oUjYk49Z8bZFWtKGS0
ugBzhtVU3tOeG3ST+g2qwD95seEalMV6otKaup3KiX/wJUWBhZEqGaommm8w2+OH
ErTh5+Xaj+gj3UVPIXo7oZTZIKp0wHs6S6mBIZ4Jj+ljMt7SYESvcRaiWNbAV5wu
O+inu0+LlA6uklcQ2ZhAouRQ01aFX2u8gK2+3D0vOo39pvMfZU35K+fb9tmwalD+
poJSMR7czj3hxjM0gQELmOMxuYiaM83PGXBqw4tGB5Q3pgC0hkwvkDCUomedQ888
d64dl+sxewfmDInBgOaaifCEWnRBQm/7Tkx2Z+8nk018FU3QU9phQ18cDlKQwris
5w9g4bp/rRz8pycud7uUBSAnGuduP6ggXxoDPSqzpdLg1xI8pwvo/04cp+fdmV2W
1CjxpvXeMGw+TXIQ0Fb/obz74KcHo5CTQ6a2JkYEuLMDLuz5cJQmmNvYwP/ylhNp
ex06tpzDVCjQLP84U+G8FvlBFSn/0mjL1fEFj/mJy1oZKwbOLWcns98YwGzHXRVL
e4+1QcUCob6eFBo/a3GZz6xotT21BqDACI61yP5IG+5ra37wW6UT3QJvqFAv5K2n
2pDhjhJNo/hrEVvwm+qfCkRKzvrbsPJzUl4/hjONX+PtddYHmaU065bcPKqIEwOB
WNQpWBsC6p9LnXymP2hIuRJSf1KmC73RiZzw8m1rTUaCSpEe06YtYHKX+sJ5g1sb
qVBhhuODt5i80l5GIGu6RTFvX+1hJ3Q4RDk55swC8hZ7Hup3WyKg5FCJPrZxf22E
5waCto+m/dD/Hk50YSTxx6F/PDx9t3FJtuxdZETzEAUbVld1VWly4lezVE02n6jW
+SGTzFev94ZEteVO+SwiVssXyXONGWyZrOgEuXyxHH8MileQvh/2m0tKLrUTpOBB
tJUK1EV/+36GbOOS6w1gm9vzGWtU9Dtb8cQBgMi3iCb8ltTzCictUUCzZX/Hz9es
uCshbAm/OQwoilpj95Rd0TYe8xnEx/exWTIchA/zCkEPgvlDtm6pBHxVY+qm+0cc
hn+2TKBIfr6H0mzi8MMrj/QyPMAVSxoqoGnivTLuoZh1TBX8oFkdmtfh6LfNmQ9T
CZbKMfDVMw+KItPSPt0F0L6GwlX+AKSSP8MCxuPyPy7maUU3nN+Y6B0LjfXxXPby
ZdHIKbCMwTaeAInTMzhEy1r6456MDkSJ47zVRQedJnb1XZKfDob2oV7hyh+FzD98
2Y1SGLgedGDJIv0UWGX21RO1ghpKx4l3vSYMi6gajP/QkS3kS9pDrU/IOeKwJMVd
dMelB1H6LCo7BcQSkQywpU9HC7XHOwIod0Cfj1xxrB1US7uk+ydj6jHcUqeQsVOO
dM32s09NWNA+SbwWym0tTjhVgVkAae6XIz9oGh63UDN6g4owI2z00EsGQKEFaMMp
wi0PjiM6QpxdlySLFyWiUU8Xm4n81cNPn3A6FyeL6zyvRykE0UNEauSfH8AWCEGw
QilLx8XFH0Gsi3xdyHAE1q8knze+Si/w8dEAjKKmmPYlmnIGGSxRcIQA5vn3Tycm
52p9KfnVtvW7ICEWlq51yi1Xwq9ZY+ZLNbjy6wuGoErmuNioFPwGlZmfJTLlgBYZ
JOM1La0ucxzQpx90MDg892RfNtNbcbIaUgdRkYax3nAmyQM/ou9PnJWnSlYkEBj7
PPsUQdDHrp/DzOOLsBzXcwUUgGixLw/VGCclu0uLMc9l8rHeZ0qLlSj7M5541URY
l9Ku1DnZANQld2vkvC+1zMmoexEAWBvreI4fFG5lA0SmgKpmhZDDomvx1fHQWr6d
UDsY8NgWUyQMfdygitSbsz8EAa1t+/D39UBGGdlv4Lk9An6OQH/Oppgv4mdaH+nY
4Oynr4anounZi+VcgG7ZHGMzFkfLMQSph8GKZ41js6E0aAMoxMNFlu0VqFuJ54zg
9SYSgk71vnLBnVrDSfMX4JLKT1Wvfas3ktHylFhx0iw4tT1guJgMk+V/h771QSfU
iE1orBDMmESGk+i5x8GtomEy/AenBgiVuE48bj6deGEQNL8DFMhgRF1w1mmQpsK8
J2kJ0f1uQfbKGhBU2oLtl4aNHiDcYJhMOy2ohhG1FWdn5faeBq6A6NqJquX9nfJ2
36M/BFS/tAL+oIrH+M4yxbPuxpALysEuY/mNPXf5ctxHELjy73hERuGoi8ZjPntA
6cmjxxtLUQCHZi02d3c7EGlCZlO1tvMqdQnrKXTRjmevfNZmKGXtm+iOQHXO599f
aUQ62VZ3yoWucH91lMu6yv/sQCHue0HKCfj5BBztnfOW/ZlJzXrz/ahJW/1T6Qde
DwKquWhtBjjK+EtXjBOGkWgHU1elUzWeoL6Iup+lSEzqQAHARlRz0m2fnqiz0R9Z
47j071azIQp8pBRAGO8UWWuZ2w0LJIKW18sW5DAlsWAmASKoOv9CSCAHmo5S9Jnq
sgq7D/Pwm9RScq0+ZzCwuriDJgcBwD4/fLg+CLA2uiSeuyW5tcC4gSupqq3YHoOy
J7frRmcbJwXQDgtxvKHhwWTISzYWlRLpLYP82oP/EhnhTgINmb/Yxjt/aZLC97WR
6zozpNVuNX6ujWlNL2U8kWell/QQls2RWyRXrTULWzqdth2p3Lia3I/vpTHDXZyi
K+uOhjuaHMZ4pZzVBCFwOenhNh7/ONC5K1Fu17TqUaSf8pt0wF0upf9yVt2KwIoi
BnKU3v8lZT7nLk+9PypKuxblkma+wyAJN0FvssnqGoUXMXpPFM904dB1MQ7/pty2
w3Kgl9uFTfI89EFDei3HsylpJH2CEFF3QJZuuLJmZCOIx4W7TgKCRiDEtBRwBefx
0vgnXCVR+7ce4i9lau7Coghk7/LcgNEjuVrvFlaL75eKuRqs5GRjBJlWD+DddVM1
D4iiK+siWqqSP5WuHqDOj7Sm27whj8dIiQ7HLoeX7pZqak+W03raI0bX9AB7NUG5
KksiAw7iA3c0Fb2y8CVREN9r4EA7auXbvByJxSgqnuyIrs/3mVCmo8EMaZ1dVZO+
B/wjcw9k49FI0NFFYw7uXi/a/7Yoq+74dVpI/jySPdU+m6GJAbyOMbOsrRu36tEJ
OMRnoCaRvhYrYIBJjpJ55byoFm8w+sqRmyorxEmKA7kiu9RHo2wkjPrMwdjhZ47B
vsABiXz8x0GaD4vtcpIoZxLZ+dWAsMFKw/DmiM4wDBhhSiLIGb/9vNotvF/nw40I
L3M5PAVlvRoSga+y65+IXe923bFXkK206JwxQjXb7zBquZGo0Yv/PAOGFUW3q5sC
Mm936gzAzO29XjOmfcisrp4F3gbcT70lj4FAdRyiTcNtEBdjd365Px5ke63Xfu1x
vl4Ij+PQULl8juKDjfwqzVK2T7xYya+cTUt7pgWzSo76IDMFfo1NhkV8Mgj7fbYq
43NqEm6rvZ6aBfqArk76rhdEVPelTuV2qnRU8H9ab/zfGnZb5AtqS0RB2Q/1FaJg
251JvtS0a0gWHbGo8SmRPLSO9cM37j5v6dAfTCRzLnz3KSob6FdXs/4c1n6wSrGG
9c5KqwJofpbvwYYuDiOmWWXtjLpj7SxR1pl8kMCvvIM+tjn18fvBrBBf+iJcK0RT
3daZYNXYryp4oKYluFcoEsIL6+xD0H9MEIZfXyRrCGxeVge4Gh8wOdW88kpU1zU7
Xo/pQfoLHHkUhJw17nEucyeEhWZHqDQ3dFxx+sTw7iW7O0XJs4reWxAF8HOdwnL+
gz/9trKz6HZlvVtBmTbGYB5P1e+1sVY9uOGM6a3Qw27FEAIxVi6otUgkjOWVFVOo
tCWHzEpo/X1VYKm0vgpv0uLo6+I0tx+wgpKhAFHVZrD6Sn4pT2hMkVhQgWOJtq09
mKqbBQ3iXgz7NtIi4lzm3anHUm9b5doEYGQoBdAC3A0T0OLNGJ2fA8+eE6zOAPDx
KcPyG00qUXCBix48ZxufJ/OUFctEprX9C4S0GMRcD8Efgi+hl6lByWPg3IWA/ZAG
d9bQg81vOQ/gN0WjtM49lnwSyMpeMbP6/qy1y58S50LF68zhOi26rSdoCfwKJzZB
JylB81h2Wtpe3thqVuXdU0cj8qBB4fcrPtEUej/CoHFxrBbaGMx4dXwCxsU9H0/u
tlFqAQWyAQKjbQcAK3gTt+UhZoYC8s5X10FsRrN1bP3Q+HVA8mvPvaJ+6vPFQAXD
ys+wzJ3P9mv9WqqX/vWWYwQAP83AZ91un64UAoqA/YOM30nGapCEOqDJQWPeL0De
HCSkV89DmMcOUhPOyO+7HG/NgQ5V6ZqQiolryydUCm4ivIXJDV2PUU9s+nas1vED
9AP5sSVEQwmkc0mI22qlej/VALPrq5DZjf8I1y9vpbLpQ/1b+zzVNbOXEoDO1Q2H
ZcsMYmWvtiivr4Nz0HOjexskCtFLrIfjDjIc7twIgp9M84OlyHbpJQJY7iDom5Ys
+H4aoi31G5ZqLCrzTXZaeas63sYTJIlh/hN4v0RSM4EFIwPdhh4bgcIL5dfmyp09
FnqZwu+UO99j1GXRoTzJDIbg3zSx0l7GGOZMJJi/6BfhZfI7aPgtfDMjr8uPWO6X
VdhdRHjrPy7XiSiM1gu2COi+06e+Q+vspsEenL/4z/7JvTLH26Lt5wCqFQxLsgZe
+4oDdx73Eps+scfgJYN2+QE319tIFaLtgqY5NVxKabmgFeBK2faKu1WuuxVYnGIR
qvNhgOcsrfilC2orCyUyz96/U3vJW8M/kS6lmvt6lObfhTC6Ia0CaPGBHk9CYF+B
ETP6e+lI5jXbBPwzN8brXdiFOmdaPPpBCe3d7R7h/S0LWrFhLFBD/wCfovmI4FvD
Qn9zs/ILKf5JMgBD30Q1PZ+hM7voIRUYz1S7ohVQcAhQ68TaRngcTbO4UwZs6m2/
D0+HEEroFBk5UFg4mk4feesh6F1yvcGWIbtLkpl/WJeAikob3LYTAqu46wLd2+Jt
YuPSQT3LS8ziZt8sXFU1YIaaZNlX5+nWyE6cmYbj+A2qOrvC4AexJ7LVftRkm3A+
S/bvakiE6SgeEUexbzDZhmkZ2NlOrt6cqnE/i8KpibAu3Qm/5wAZ5JWiHsLQgEcf
yfkZ/vDRuBIcfRNUySNzhx/hTcTbAHRXiWQc2DcfTPtj2WfjkH6g/4XaUPdnfv0M
0ZDv4oyCYFyl24wanuf/bMjYYIWx1SB0Pup9ZNbVFzW/XlqeADwy6spfq5wUO8mQ
fjZXrIp8a0/tvrCY83D0/SAB2qY2ptt/raACP/cvA3NEf4pjyT1ArOxxM5JMYVuL
l5Defut5f3T/SHvZcu23ouJEAd2VgwQffUC4fIwuwGx9MwJnYXCBg00AS7nQgPpa
H56YcBt3b6hgRiTBXNPqZPyn4f14ZUhPWFUE2ejSEq0A+i9cSIaC09T5M8PnWsq3
6iO5jsePTjPjgzAqfspM+rrnqP8D+aRZR9kspxRp4JRBGpZ8KtxGFu+vE8NeTHHJ
B3JMf+/iJmUy5Ak8dBA3myYV/cBV2NWWaA3YCchLAAyV2jVqOwG73lq1dmGEzW/A
QGfindq+nopRsimRhpe6/yzl+k1hmFYrH++Y7vJcjWyY8DfgOwCEZxnZ1Zs7LR7h
ctr6q1/OVseJKRhqWaiKwX2wcjJ6Gl3Fm+Ud1WKFNADtRx0SHcLVXIgs3E67TfnP
bWVJxrLv6stb8oX6hkxYBZVaQBJ9l4icwsGLHoFZXOy1ZXc+QZeC6LgtbG4KoF39
KLma4+sksuJaRkgJ/0QQMINWO27o3LkspALjnPVggfPyIctDGeEOmEGvtlyDiyP6
ogwx4PE8y24Me9mD2VRLPqnr47b01iITkxE8RYNNk8sWTxVf6jUnhPIzqqDExVAb
e0bZiLPSP5PAZDEPHLamEfH2CX2l1cwg3SyqnW74WRVJhk+BRb5HCd630oHuyGJR
ZHay5SBeY72C2joTe5Uxbg4uXRDMt4z8WFcMJFfvqQm9o6DrtwjtuwRHdEAh9sC1
jggE1fD4GDckb7iKUAKpevhs3kWp0jlxSMP8TyU+FLQN78gto3t58rxL43cb9Exj
OM8RQlqj4EJEBPdvPTfuK4wM0FdEd3y3OHSzsVbq79GbZlaA0H0Vo1FDBVIP2XBb
DE5ETiX55OBXMT07KywcCrCsEiCETH6UFGjTmpUGinx/RFE/iO2Nm3aOP30RXQaO
Qw/PuAyFuQSeElDjN7AW/nywYw0kJIRswxmP9cM+6zLjKugRtOs1hY+7Q865C4et
gPwGqLkLNlpmhH7H4CLMUeeicHissOFM1O6lo6ZcOdd81NWxUU8N70UHGfVafxc2
L+skdTg8EvuEhUAXtRiyf2GCkC5kjVckFRf80RA/pEgoHWUs7YU+gig3vgGLCMN7
1gvs/wviNqR7KUvrx0u5Dy/84tD6jyKSPQkVgIcFyZCFtwNPl1ryLxUG+O+pjYWn
z+NoL+dqhhEkg0sTnbXg+I58RjoJ2nokscgeUlbMA+Jova2au0XG88ut8T32xabY
bsRVoj++IVe+vSYgzerLvOwUkrdmuq3x2vgC1KY9cjkF/pjPZVQ9D0H06USDICRk
No2SO8IcC8JNXAgKI7xX++8hloqkwcM0cRcuEp5nbuI0d1sw9JViaXqx1o1vNC8O
mC41lCP0e/u6xMuJECXQbtHNi8RwBnhzdYaOedIQf0IJeZFFzpFkxAkLyFNu6xiZ
MCI7+Po9aMRhs14raqcomLGqZbhdxoXjDtMcYa2OmdfIQ2is5WKoRep3/Q83OhSX
RWE2+hEqgak0b6Utlgghre2ikAmUjUR08yEhdP4yoVJpFqGnouP1FuJN324/dtKl
70l/+sJFmSJL0lLbqGZy6oJdMTGZMpZ0liZU2ZSoi6ZE5J/x2YFHBIvh4u5W4zEO
GuPOCgBcStkF7P8fD/t5Yj67v8umEh0e+VvLYv7Unue9CjmBN12edRx6eMW3TVpn
gJtbG02YyFhez5hvPcsjtQnFSXnoieGJVa9QLfbL5BNZGYHNHCU+jt6COxWEfYgf
pwhCNreDY7gD6lzui9TIN7Fac6tALEiMlg3Ytmo1VIbgFYAjN/W9RcQwiBCJXfY3
9HoesX/S4bg2re4QQbBUTpiC9SJwDFqNDCNUHjWkPN7+SOsyscXOOGE4uc0UOoqF
dJDy5GeLkkhuvdhyuFpiJvO/WIfUHIkUAOBQPsIVql5pk5U3X2F3dHARXrHVLG+k
0HH18jEeRbbx4d+LEimNSpg41FLKHLQgGsoe8nSy1epXVRUCz3OP1aTE7UM91OGg
rKbg4wctNKq0YAR2xKBMVDSfpVstqc25OMDSwzJjKPjdJGGgvx5lJIKYvBPPnuqJ
GfEB6mmk+kMtbgiBuyjKs2Twt3XcqyVMNhtpXeQLjKuHcU2QW9ItKi8VecqNOsSA
0Y94yAqKRwUN/fMqm3uf2hX8fQ3IU8jIcF6q7tQpL+p3+oakAV2SdZ2I+VZrri2s
cI+Z2iISqA1R1W1cQgo7EDWw2DP5EgCTmTx7A2vSXopHbJrHmSzbIifPhk9KEC+C
uNJCbr66D68eAMOdJ37tHG8WrfgXNMe08xPcVKtTLJ400A72fHBMH4+iLq5SonQD
waRz6SC3TFFcXRynSVr69gMvPjVikykWAdcAkhoOfKpieud9pQjgBXbj+0kfdRht
7B7nI6CpOl/c04QqEURI8pukc3KvApoSX7s2l/Nen4AwgXTWFe69ePD31gn/kwsh
rUxNZr8KdLkFSbZ0z1QjqoCq1hzYosKawBmnhNhAKY4XOY8IyNsKHofuXbe38FE3
C07ayHg+sPlIUjaPErGqDEeGH+66mKEjy0AbC3gdQkVXyFFoCPHmtgAmcXtTBS4x
NrEliNLqe/A9kBseZc+5y66IZJanlJEMX20YjEiAJodRVfXDCyq5f8LzCrXRlSyp
71u6d+sVVo8goz8P3OgoGikcGP+Hrdl1Y6SfUUGD/NVQneADZ2iQcfXJQR3AUIho
kpIpOZccuAHCU0B87b46AaV2OexK36ESQxDBggx/WQJZHh6Ir9lwbbcXyPv0c2tZ
89XvnDnjVmHikBhJtjip/UacSzoI3SJnp7kB/XoFXXlUiij+VV+E2s2+UcvQbDTo
nIQtVWRJ27AW8oFY9zhlyj6ByigjsV8wIF5DYTF+zW/2/02f931FY3IcyfWfgV9f
HIZgJQ1QWUlcnDl44pq6fOo1t7BL3np4iEK8xRC/urIZZBaqq5kjwO9Uc2paUJ0q
D7q8cTbtNabO/U4+tK5hbupbQLuQ/nm5VLBzcI4uIgkW5VFC5wV+VerN1AzctQdh
Yqcs6F/qj9l0ymif9t/IrhhnsbQtwqznXSM8pGUt3FLKPi8Z8bKQUQVOgCm4U/Na
F60oT64prt8oc8RuGN63fVjhwfn50ivS1oRtGm+kNLxBhOBZuXqEzAZgo4FUqSJb
Kx0Mqlci2Mc6/Xv5f/8hjrrxCYfBgc0ASXjFVVHfoGN3iKLLFMZEyzfs4UZ2dVrA
bxKbDwITyFPKXl97UvNN0k1gYuZKk4tPCBGr0pvKpURNg6DUAAq2Fgeo4wPdiq30
g08K/xXBcT2NElIsrv8lW/RUrtm/iILsrGHJBkjMkHIm2+6WlEKWaGaI0DECLQEf
nY/oT2rfRcD3OVnpqJ4I90ZY00nwSg9YQ+Px6Bmxxe9MxVjeSXcHKyWC9VqKb9Vm
u80a6sbpd9KPBb+2TB9kkj/jYAGualyWnoNHBIxRtfMDJmuz2KTXVh8Fe9VY8OV7
9EF0m12IN66V9ZkyKAha/wWTzSx8/4BagRtb6w12ujkRA6bXB0xwo+7hmB5iHQsW
FgEg1rGG88oQ+gb75Xb4+nFAVIScnHVLQFCBivkYbX0GXtHyOYT3uu8ijvv4TREs
5eTrlkkJWWTpL+9+UxrdOyuczoG3B8GHMK/Wlj+o+LwzBVajYZZG+8OPUPCICsyT
UN9geFSz2BncRMRWQIOFdbWylacndNc6XHf/hRoxr9wCcLaGmAA5hlfmWfhtc4Sy
PCBPl7mmzdKXPE1kEvoq6ra5sJOsJ4MC4SY5elANNkHRW+jT035tu9PYte9gafNF
K4WFJCLdIaZQ/L3B8ZPhYFvNsRXy5J1bQlci1awWS5pY8fCcTHgdAKBWJFNT2v82
LrwSDg2jgTta9edsaayAoC1IYwvJvWIkQ/L/aY182ugC+Uq1OqxFWWFUvUcwQZVp
9+NrLHJmmZ1BNP/wyd3akRyofOs9Q7n7QbZmhNp2gNwXdHuCHQdg8H385m6dwzWI
mwG+hpoXD5rsC0kHPTBl7H1AJcLCid9BqTG0PTstPJPvxtpPBQfPmbZcD7A0GlK0
uydgAEsicdOkrF7Q5PmkCRmTMpVlgNaz8lwCnyO8VZfk4xcMtaSz1tuN5/VHKQOL
HmsJBUs3leGMN2CUkxYltLj5MeJFRThQSK4+YWdJ4yAeBTDJfzCAXbkfO+jkFwHC
cfxKe2t38AehM48kWGH3IU9sps2GyIR0/Yz8cWyBRcvDCQECGmpfBxleNl1egLCb
VmAEWglM1TywEmYFRZ3/eRVNf0q1WOgsf5eKH7QFXsKM1Nn10ZmZxyTgxwDzHNSB
2/jVYru8cMRUUQ2SwM3PrJQHmIzZEiQZU07QzNIXlSIc3d5cDb2fiBKHBQp9D9Ij
jfWWRQgDAJXRaGh40Bq1oExCM7mFQgHk7qRimfz3MOex3hXyeQLsJel9CHYJDDzn
xVaPYL4gR/ApIMpcaCWXNmYDk58n20vni1dASCW7r4p0BJDYH93q4vaxdvyHig+g
OH4SQCneX/cQqF6FViLTV3KWYWZECWLO+t/PZIJmylYmT7yGtRji2P694FqF5ca6
h4zi87tcKth0T6f0P/1NnF62GVPv9EX6StA8dIdgDqOq/Ay+7NNBSITd7ccoBwki
/ogniu+a/7YODuVUlGQI6WNKr9wPK/wT21XOxPGb7GuzKOMiPp9H+Kc1eiHMo7jx
GBE7+2eWNJ4N8C4FUCDzgewSKXWZOjNk+QjQZtcP5s+iPZSvRLcG9fQBeqXr3DRQ
ki81RflVG3+TmsG3Oux1Quhih13rITAZalwMPx9U0AJodznRFxgl22DShX6MVWcj
pHUlTtUMdY3jFDj8kreq3KRqfc28xJG6A0YqaV9lGO2UctZFQgr0LlynvFqn7TVQ
7lsLKDv/gpAb+fxcI+tDAMl+Lzrh2PABYztjzQ5qA0u6R2OtjLs5upVfxHl+jMKV
qTSZQaIxXaZk3sAtwHxJE/+aJTQwNvHervz56+bbLFm6MtTeC12ZUDw4Fuw4RT2v
tGv5+fF/oBNftIR7Y6Z4GaUVmipZuu0gZsSaSKqamSlzvLENZ0gYAVHzkbVWh2Gt
URJ96VK4bGK4xggJ19KE9zIRqbZaPrzLVlBQy3VImKDq7iyMe/jGmprwH8NctuQV
XPj4AKWRYatkdi1sZXiBL5yV1Lo9Yrbuwy1zML/Gq6gvuPX7hwTBRARXt8wSSZFX
lR6YhAZPUfj9LVtAHd3/9Nx5JI4Z79a07+V1TleAOOd9oagn+HSPyz3YeGk2P0LH
ObJ5NJaQcIRMe5OiiZKuL7bEovhgXjhwIfGQoIE/CHTSy8SSMelfbhW+NI0gzm8S
qE1hk4LUS5iRbGpRodjkr1JLdOHUu1GgZsyyjqQx6oDNFMg57Z4K9O4JjfCzekmu
Ni5rJJoKCUKBddslY0AGvivW5UzdXeDVdJRLa0fhxY25VQugJqIkXM6bXxTcfyO5
bL723UmnpLDtH8OjtyYl7aikvjzJDSHIvLk5I9IXIBp3tET+VJEHLx9AmuzfSppx
Of13TnFTPzYpBO+Et7g3xyw5+W8JCkn3fhNR7AvyW1eiqCHINyZnnm9K4YWliYHk
PYSBeEnsmy5Y+T94cvRxyMSWzUZeGIakxCBFnG9KT3zykk0Zr/RgSvOm64rpdC5S
8zUuNZ3XE7tvmS8XOz5k/i5i9saG9CRipZ/j5ZamjwUqbM6sGz07SdfvzK2+ecAk
B3ilWrGtqoe54f8gpnGInLxQLErR3NXeEHeUJFATkPHnv+HOa55by0IN/QqW2qaB
tXJ+xKy4puAHgRSnri5ekWySj+NBH1OtKQHL3RSx0tV+GGL3UeATQErVDcANJLHi
7/xPMC7/CFQrvMLW8qRessR6QFYNv9wgJ/qoQeZD0dGtDKOI8KppfkdPvV2y5o2m
69RdMJ2SmFQOUtxhWOLVN373raLyGFIFrokqM9F0sAuOC5Uyn2PgBGdIbCdJw7Z2
D8itHUA5P4IiD4GhXncGBMXdqMB/l5OumGDaf6+7ToBEgeB/GrE+2is1B4E38V1x
7p4YNyNr4sV79aBrL3i94swNZZCzgvBRJqHcH4J9O82FuurE4t/9d7mZr5m/ZTqq
rlvHpMBZhns7W5wJXBEjhH2YtEf3lWZqzBkeC4w4WbsLraejHvWNJh4+F3RAx57s
+w80Sk7pSd7CK3e4Cwrjez5CtRy2ldeVsPNVxCBmsQ6Aqle8i3TbXM6TUvJpIxG1
RhvmhApf88UL9zxjRWImbYmoiNMVE9yhh1RPyVoI8VBNIqbTwaeT3YBZ+b48aSNH
4AmAU6PyyLZMYWmQIk6sr5jAjfrcvIdBPTKiPRyVrqOlzy380UWysLQrNoZ/6/a2
ZsmlKjKM4pVIYEiTCK6/LUe1kEZ/OEsTxKnFqFvSCBoWNhO3kuU3DQdPz2EzKfRT
p/uiOUFCn+8HIiM3M+JJa/uKz0Y/nrxu/tgfe9X6WoMh9yJ5JFnQRUjs3Y4r7pk5
aZOBNwuCQBl7E+dEHFw+RfCHhDlronmrvNiNagNsXdWutvq4CrHCuXtqQn/aR8UM
HF73q73uHsBtdCt+7jO1R8DDnKlkC4JG8e17U6OTGCIa56KLr8GpuhmAQp5jy8u0
D0mIrIRpQ8SamAfWB5/ohy8pl2+oSar1NMAzBnqSj2ZguccoKk3bPQPXmMrsl2Ig
OMcfR5mrIBndy/vm+5mLw/7fbWcgc+/9D+5w4/wtX2t2FoWDQEXFGyuqE0V4Wzze
9di2W9SFpa0Cn5VZlv0QXK+3ry5X0Yt3dp1+fG2GbWpFagXh+vMM3vZ3GEr3pHUB
Q49wG1V7jHHuW9dc2VlVllxUSw405V6IjprY/sC6LYJGI1kLY0PLTGyuFv1NEz5l
0C1e9u3568z+/EQuW2hQMH8eQJ5oqIVE+ZvDD9+EapwvF1du9FjG9/p9i3Fgo7EC
rwNZdoalqr+e2hU4w4GqBQ1RvMQEj/og0wMeWIKWdfweZU5F7fMU706gZv+3BRUi
PGxWg0+ZocM5yZCJ7eGPArEzeYkVCV3nb0QOeC12kXDeXDAoxEf7pd/M0Z+dlCMG
8CUO+2L48vQ8qwVhTzNf/nioQEgTdhPJu6LrN/v33PzKzSQx2VFCbc8ivYkUnbZ4
T64SKuDqPDzHltgJ8ZfT4dXvh9JSxDPdH6I7r+O6K2RW4kkaJW2POI9uVxoC5Jm4
laR+hLMDFAWTMH4Cn/3buz3tyebdLIF8dLYqugIgX2cQBk/Um8/kE0ToF+3pwxY0
wHwnqlm4gJ01/mSTtLmVkqCSPzRG1ATdFeu8nSLDaKKdNSw8wi4id0/0PEoVt+am
OpIDGIflVPqLYucz8miJ3jCyT5c8uvwYgUCmGLNCYYn71QvrX2ImBayRRt6byWKR
gvm+YSNhzM+d1KdJmeydQ31EWYArXAOSa2M5F01KOmV4ExeVfQPr6LR0SY3QkMOB
haQMhZqDcZ8NNVBchUDEHNOa5IjmRutVVBMVDWn18x1f0EgH2khU1x0Df2xXxDoL
6Slcj8V0E+hH0ujFaLVqIG94GbQKssaRS6fPoj6gY+3iZab+fT/dS23cG/c3X/v3
1BNjXUUtPEMAETTDlSI3GazeYW0bRmeQWOGmz2/e0Z8RBmSfdB3hVTjVrrZGA/5x
IvGJLuD/d3MY/q5Rtyr9lR7xDsC23sdSDtu/yn1khtYGHJROvOwiMrUOgwHKYc1T
oWgfwyMqxt/fv8di30/zN/SjT8/XOtUH5xsTb9hJ4ZEOwgrc9gWRfnVAqMRjEW71
e622H/7qKjQvSYZlG+DObx1qXxyUyjqR9lV2O9dpZDxbbdpBRg9Zrt+edCTMUDQu
oNoCaxsL184j0bGVMZFi8J/SrYH5RpxIWML6e6KBjUAL8bvOjjNvKxKyRUoQwaIb
JdJnrAcTrUCSXsL6Lc9K6bDijvpYxSXNZrFhcsfVpgPgSxWwi8ApjuC3A9Bo67Rx
n13h0AvZm/ITGyN8K5f/lyT9Tz64U+psKc9aYSPxkPrZWzjC7/r9k4byaXnD3S6Y
k8lvjrjv5QqmLFrD6hyOxkJSqTxs3JzB3087zeQ0idbI4q9I8Lmw64x10Ba73evW
WnNHE0dFt3B0SKtO++7QZ9poO5Npc+j1kaAnMQip0lcKaGVOzY4qhsUo/ZCd7zMc
qf9vmmcMkHK575WskiyHwPLmK39O5mb5LhQQou27RCHM7AUG5JUlhLiwFwcTvRdd
wIRRM6Psp/58DB3rpYPyeRypuPUydufVxS0wyUSvwKVBPxxSfDK8+6vGarun6tP+
wjfRzsEyK+JjviORyexC+VouQKNExIObCUM9X+AOVDo1nJbWLnrGhaPnA2x7SWrE
fxzKwantc5N5rqYzupBe0M3r93GZtOp//t3DtW+rEOW2NFnXhqo3ydpQs3W1KfsU
E/GM1uA6SOjB9x+nE/+z3f9gwCQKKxEpH8etkRAht6ACF3PFOvNYy4j9OMTn9fxX
RZ5642HAFqDpGKzStdPBhRFitJ0mTj30/CFNsdaDFaJaPm5Bi5igaUb8EOU/HeMy
RU5BlT/rWSrSNBOMlxNseF7nyW48OyhtZ9+xXAp1Dv95k8LPpyTypP/VLCPGlzmG
ZHFUbRJFEfmlcONm0t/cBDrN0zqrJDjdP/aYwRX/nKi91zTwJiuPy5Zp3yts1q35
bW2RNberHcouaN0OjBkk3P7U62/VImixA4VoflW0olbgk3/hjoYLNwx4f82/iX6e
9eigqhaNMgWIrE0M0R9C2DM6WdfzqbMMefIY2NuwCOkpLFQQSveMk2LIWRG1EV2r
ybgwTeW81/oVZ9KWbFnHbESgCzShUOtunfDTd+5o29zI0nO9U7fqK9jydFDdeaQy
WT0eSr1DCG1v2Oze+JlvUV3skSl2OvK0KSVerpIPtCTLrp+Lsun/YN6j+PIqfBmU
n2qNd6lBNWZ4yodBshzqYpSNMDStXhK4deoCR1RvTgwze0f+MUN2NPHnsGdbpspy
WxQUCj+cDcImg9/IlY/oqBxiOpHJ8SpFdwdxLccmM6EFnjCndzXv/dYkvt2CLVuB
hWcGINw6vNAP0ApXLEhjLf7sD6voLfL9FgsDIK6Cjjj+NCMCHCoRLzfOXHuqQkDV
41f6B6vnzlH10QCcxMzJrIpdqidDe+by2J5nvz3VnSK2n4NOuqEGlUYmnFJLxXlS
j8dn6IqobSIREMx4YbO524ZnvfwBZ8lT9oAf6t8Tvqx84mpmmmjM9U2aG88dZxTy
PIazMVTAFS2bZthnXZB8SvSS3tZ5cWjckcvLRQn+Mc4B/eDU9E+ag6GmcHZHKopR
Vu7bOZxRy4hNt0ibS6D7YJufNOQMrognJs8qFxqXiSWILRYk0uHy6iYwYqIfGPTL
asL7U7zzgBFNtRNTrSu2FVBvEIna/WdLdVNcv9tmHYDIjPNDSpaiea8Eg7pbcwOb
REeKvbvd0cyNY8VRdTW6P1NC2CvyeYwDo103DUq4PPY60JXEG0sqjkSFiAWS7qEK
ALcnL14jKF94NAlN1mSJT9b1kjBZJxrIyOVeLfoixBYGsnlHAhqYTSWg2akY8OnW
`pragma protect end_protected
