// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:51 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
OONl26srovNZ9JcugrkknZYbikbprcWyCxZ0CEwMJTKGjvFSQmPbFa9lTAC5Bh7p
LmBPsc+/nWH0SV7fWEXCxI/VVgClZsZv+oiU7GdZrZHle0sOPvcsDS5WReKEKtld
XdD6mZtJRxpvpHzL0XYnnblJl1v+9IxeD5Ecu0QtqcE=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 3360)
BDaRw2hzcHUdcStuNWq+MWahYZvgIFZ+RB6t3VfIIzH5wHNWUexAFvuMi2EWx+os
EosYpUS7z1hmmbimsBKWtiMFMnBUQrjEm0rNUYCMdmo5QlcrVD7/AaJ5qjALoD9Q
U68OYXJZ2akJ5hCIHUt/369oxhxwZnjcEuOZ40m56PVZMIErTOivTSatqa/pRqO0
tOUK5orxMHDAjB84WvtPIVb4bLYP1CV0P/jZm4+RoTlW/jARawsG8qBG4ht4GvZ5
qylAE0ojKAci7OcK7fFzRk2XT1MS82sDnbof7xIFTD4TKrsNWqJc0QbqUD9hAOBT
lZ6ppGL6r5aqekhxYjO0vyLUBrs00Aig6SNRxCFYbKnxw+4pbDALwG3y9WIGWjSC
L7mLeMJCC5H2PuOmHGDZZJbQK67htPN4pyqsbOR28O0hqyhgPn322Xm8SgemMMY0
KA5DLVAObpHquxqu2P/9BG0Nfr+/pPqGeFYwe+zo4CZWjWaB2KFTNXExeQ5eAMBS
3eOsoYYbNTo1cEbY/ASkNes//Pd+Hlf1w+KI0nqbaZH7/nDmpaI3oov88IHfciR1
jVPqHgKSoGU+x3F1NK1tB7LkxkvSg/E33E1hL1+D65KkmbB/Q6lJBZkMDnPJ3dlj
Ru8oN+7P2uQzuxHq/r5dg3NVWV1wjlRGQFutPiqdYxaUWr+EPAaVQ/5RA/q6l4zk
4PyuWwFhSn+sG5h9DJyo5kHFsnK6V/JbmQc9sIIRO2q50aG5gUph4c1cKzowUFLg
Dp0kEWPRhgCiCKlJqSYrt4YINJ2s7dIWYBsvTgrfkbKK/WOxMREQxMi9ncfUsaWr
qwtgnVAZsKIdfCKrt/t8ot6WviHOgA+c5aZMnSoOVN+yRsjCYIeFqjhTCe/6AmCd
uHc0WOHk960s32za0K/o0+CZcospNzSFDK6ME04gjwp7KK8W+stmKQf7AsScehEm
apBTgo9KAr5fqOV4DIgsK4thHw0+0oHf5khYmwkG+OzNGD3Y3OTvUtgpAZfOXONI
lYgxrJPBUrsvjiuSYYFuzqWmD8JqryWEd3XiXHGVeUe2YQabbj3NHhjZYRlfP1Dz
sOQ9FXoDlWPUecKLz6/2NCJnhcaCtQNxb1HK6Sv9WR4i3A5iMokDkqlS1D+p+p6N
7Z+eFwilLZd8Y7rFz6XlTYptoSgkuRUQ5NXITH81khoCGBYCf4T64gkOitN0f9i8
j3//uwyfcgaBpFcFytA8oa6sCrARzJI9iUlh0rVDeGtoeOjVU7FRmiMCOclQqLUj
N9ZKfs6QnSrA/o+72tY0CaCmBgWSrc5woSm119owFuF2l5EzGqszpulm30lSw03t
hzVAmOWyaPHE4DxgC5uoGpPQ16oyTLhsKQCKu8jYA/fNTSMuNwXyLkTNdudlvOqD
lOJiXNsqXlA/W3zM7J/LlIE0qiAEc1O2b+kLcjDF9s4K0XCPnNdCW04gkN9tmH34
o3odycve2WYARGjrFyARMSt7xYLAY8YG38nz6+kuqXsjzejdiD9JU7Z1Z7LTFog9
+/Or3ZB4IsZYGiAvppsFJGDtFSeetMG9LyULJjHRtwGzNy9Gu1h/uENVkNjNMABL
K0dqBX1E8G4DhMRnV8bmPu8UiHvnwG8NktsUC1XLmdak0mq8XqZQNv9qbCieFFPz
kL40orY62/uoOzTBhL7CRNRWniqCUw604FQh098XhBFUKPlP9OQAHr8iaCwKlwz7
HxbAusq23kCZR8YIYJtQdDo48HAgCkGSBEiPZCetFvBMZuhsTN24tKUq5221kBR3
OOFa3OT0+3NV07edIvqrlX2xV6DMUK9hYbuoDs711BDzyAG+WZDNzbZFPZItGiGB
srNocx/ohlSzxbUpK++b6ZgFefBtAnQX9fAgM32EGgmTHmqgfBba2ibUmTiQtcEa
Vp/XF8fl8w+0K+iJr1VNjLbhMAtYXlcXv8d42z/A/FBlbO9/bSqb+p0nkKWD9y5U
JYQuxCd4cqMSxfYg5xedMjzm7zGzuOX/ncBcFbEn/eOIjkmZywRymp2AX7u+77T0
YjCaAaGQhGDNeGiDeYv05c/fywi6Ameft+snY0pgVQN1M4QbD3a92Y+90FVegVmU
KRaGjMDdAeVOUw+wwN/c5BAcCHXPSlzXXuW36Dggo28jO7r0LU+TOmyhdLktutfY
wEfgd4fIuhspLoZ4wG6XwYSL/GyUsWZtx91F561wFpghB5bvKfaKz68Gtby1E8XT
Cevpd58v2pr3lTv3FXard3na2cGOrV0KIPLVZwy96EO69LnoMycBEaXZlAHJX8eS
v9uMEWe/duW2v7gO4aqQVzgSkI4xFWbSAbklmSA68nsLMqX//mZ17BMsKphhofoE
nieNlCNQmr7W3w+sktc6/xmsRLR08/mkH9Gt6b0uotJJlPDJVfOyZ+cHt3ZUu8vY
V0o+1Ac6TciHNTaSygHceV++pnf378sQzGIsMSJ3FdfbgoFHcgV6eiD/BPJteBlU
BgnwayOFrJqiG6d5fZDbYj9nSDndUupgNlbCF5T5HsecHbdsHJMHznpEL00BDvTU
YlQu1Wso8ojgfBfX7jNu6vT7VzIHvkjF3QEGIqKB04JywOW6C6UHKXAsj5i9tAxy
8rqcEvuqElIKqNES9y0ook8Nz+xPKqrPLRw4FpaSMkpP1pC5bN9g7yoomrgDhiRf
8eW6Jxr5Vv1oNl60PFRu7HkPPabpgL0akMDFC/GcODy2qJxf4fl5iluYk4LQPBiV
5YQlzBz3kEBHoueSwNBJpiDhBH9JlVirLcP+he7vNsykbawrRss+A6g4dgDWrLGj
qNpr4HCu2h62gGRTCWqvIwZrlGtLZ78ggs6orynclOvfqth+qXEklyFUt6gkrDgP
HQ3dcPaCGseWr/zbxvwkwJPBVeNj0Kq4GkuFHblSgum2Q4hARSv80veuYoIoqQo4
GhJkB/QERUeX8IqmCuBqnbz0ZILVdUVdBxeTjVpor7oFbs087GAMxnJomx/h5LoI
KZb2jwr3f+EoghBJCyJMj7vYMEQPB+x0VLhH/IWg3RvjP4GQp77wJLhxM5GI7Izd
CzBtACJMHz3G+WloS3BxOpXz2fbkoRAy7yrsatMYP5o2kVdCBQ1h/wsgLcHJ+p0B
4fj3E3p7OsqQil5mu9gJgxA0yPFfd/HnO8KZ+uTQZ/GU5ZMeLGjHlIzH+AojMjI/
kpHazrldYvkK6UtfmNqHrHEaOTOEkWU2pKgbtzyzmw6yqg2Dzi1JXI+VZOaPfrYh
6veWXMpivSlw0wgniMnpl7h0t1DtaAWIIGEfsp95rQ6vxI14Jw4xtmUxYe8zbrBD
cnRlPQK8SAlJFJip04dWfeuGxd0omuD6u49X0whHkckFLmbRb5XRmoedxxDcDLrv
hSF6VmmJEcOkGPsxUf/98nUd0J/Oirxm5QI8kIr29OEAeJ59hd6sLGDo5aXKssyg
qJxrR35NJaEaEH4HX+Tasa1Hfa0XYJ3xm0tGmUdGQ96X0ZKdPK6PEjW6iSq3/vCI
miT7FcbLIyKwuflj1JMknK7enL+0wKkqb/+rZ4Fd02/7TZ+z73G6fg672r/I4HN/
u5rc3V50LQ9IHd8suMOpomTSfut3f++S1sSrclJNKP4Syg6yXQVBk+oOJd0uUZPf
SCvypbQdOKtUiXL7WFuruWtNeCHuOC2iAFWDGpmnJZt3NPuEpPHzi72qiuLNGDqA
Wdt/6/EY1QcgfmhqYlt39Jvzib/Ap58sxSZPUJBjXOwtnrc8dXkO8yuGIwGYa2Cx
m8hEibCUtTrWJzIYAdsr7hnKTVR07pBp1ieZjJ1c2rHhXyH3134pSilx9OZuC8uQ
z/M6LRtQ1+jZRlhMpFJ8pmJ8winQdzkOeYG04km88k+YQebjIWG3u75S8nNxBQZc
XWSRW8NFkmirKt7WcAnHePSHEs3tUBUFYawR+/Juoc3pldF84twO1fDY0K5KVst9
LGOAJ3OsJa8bPUKyZ6MOWDPfbbErsZ4THIs0sPb8sUL9fBVh+fvlEBKM3UvPgvld
nXRRCK7xIOC8Ham1u/YpEimcqbdM8MGP/WVJPNqEbryrzEWK5xUbGvFneUjygBGP
icLAxIAuDDDdQ5mzs0q1B/4pL3OPgzyqKKarbGtDso7UdXYC/HjNcQqEImiKQTmF
CwSjYPKhcLcS5wSiF7MSnQB0HIs2Dv6r0+h3qtpXX8SjFjNjScwsKduKlltqDg/5
0/RvX3GCx50khWuFZ9HvH69LjJ6S2g4yKKqP03wdnOMQj/fWWJsE6qe8QlKJTZHc
duswW8o+c7M3YEs7FLfXW4yWRhoz1z3ZZN4SvC1nQax8bcQt6WXCY5zbP8wudOrx
HsN2Z6DY/mf1FCd/EvjPbDFRWZj0v3HfRSKbeoophsgocHCS+zKm4Er/Vw2Agb1p
8KUrTScsSjjdFM9Ub09cu1JMOaez+CJ0QPi3Lnc89q3q7xS2BTmO64CIWomq1KcC
`pragma protect end_protected
