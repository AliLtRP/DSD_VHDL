// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:50 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
XaMOaRFZgk0Acy2FSrfFjV0nb5463ZT0AnQAuBTnPudRTgTRML59FgCHpr3GVcBP
6ngyCxgKstzLHCQamr98I5tETD1YefCPgsNV0rA/lWTsLovqYK/W/VJ3RLPUoXMu
hBEohcswKXI7VyFY/5p2z58RGpEM0606dtHnZS6tSZw=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 29040)
v5GJ4e4GNNxvcZYelyJc89ZfhxFtyaRTljW4Dy/c2j+Hlhlw7ICGN1lcdoJtJCs1
AFh1o0Y5rdseBkAgyAcAd6N/0NOprAZdMB/vyXo2nLuiIugCmG/edEhAnRB+PzZM
7ELW0lLWnn2pfvcLm3NYUEeywjupDi9CO5TzhMTsI4a7Vs0x5ytJygFbGpaDj9SI
KM3OixcVrJzti6Yb02iJHya4npuCnsKnnkw/eWPAKqttjZU8X7JF5V+cuQ6yH9qs
SR3Ns/U7c3OlaoNuD3WVNRyLYh3aBuhC3BWax3QPo/UEKxWcSDH5NGn7tuTSPwwm
qIZXAnO3gDaM5BJUnbl3VaDwV5lPnVbc4rzCKy/CyQ9NZi3l+8DEVZVXgPo9T6nQ
dzvx56WD/0wsdvu/IEykQRQ4VPd/r9S9S3aWk/FmFXmy3QKK9B2YWR44FBTXexxB
nVM7tjnB6UzCdhYwNXckOiMzEcwn+88CXC4MA7Al1XV+GWcf7rmBvDxoMicu+i3w
+fIvYgwL3MkMWSJ/gXS7gE0UiO4TmEpiHCLxwOHUmTPza9wEIZUSn/QOglcjnqsF
+ypPyWbOut5sJoWr0DIL1iWpTw3Xh/wNRdhFXMcNishFFad2FJjdFpwhtv196m2g
o24nUVWQNmq3j8lHzCqd0Jx3SnEVUPSXOeyExGZy9xg2YUOnIVENhw6MSqRu3TxL
7FmsXRAbH41SUre7VoX1qHxPliVtJb+B1WFqsOihUMEZKxf4g7feJvHj8LFH5qCu
mVGRkN6sYaIYXyWzUfAo8mkNocvnsSfztIorSrC5LWlpKtozldDVXZPd2wdoSeMZ
hWx5U4VtmJSz43yVYwzo35qvllSY35aM7uPI/4e9jowUwuCSMQQeBvaJzOEkHg+Q
xmzGK+lEuyBBBQ/vfd6HMKbnWrWVNh6CYhA60Wen5qTrsq4Jy7FvRh19vDa5PoVs
pC7S2Ruh4sFNFszcK2bJp0KKR0I65xMLV26VfdVxj0EixDzg/nwOYgAkNKmjFnhR
k5IgRQ1BETSRKL+9NnMDTBDvCr6uth0aEg6V3pZaWOhkcGW2hnvMqWadc996/No5
hhGI72lpuQNKIc9SYRPT8UUPBo1tgoid/UqcCqZEdHarpknQWhomeQD0JmPR79mj
vYzKXUdBVypSDNGyNrhFKlG50OI8BQeOGT+e7UFruyLrhhsZT976mEEvaKgbo85K
dZh053c2YIODqiZXXGvEKFxqsF5av+uz6BMrI/SqyW40dPrnw/LvgG493lwgQ51l
kb+r4ektQIJLtpcVA4ZsRybhLNIYSB0LWNCtc15O+UYwi0fmejDFj4A+7048n9ez
B6RbwYVD/I05rMl3RjPz9HLv7oTUqYlpDOaisKqdPQkRXxlp1/82eJZt8e0bvbzP
eAykjjAAaoXCimds6fkG8Q8rjcr7KaZ275wX2LtIwYr6/ygH2tor7+msmCXBp9WH
SfNyImNIfkL68BZRaUJObQHv+8c+kM47L0QnNAzdIbMzdPuftJHBPCyyuoiyOm8D
R59e4Xx3/iWlgROEaxkWS4bh5Byo3DENYRn3cBn2CdvIqF8I6PGzGbNt1p2rEMJN
jWC46EE7SwAIAmY/KbBuMlF8Wa4OJJW/ZRJO362EE3mrrRIIfHYfWIFKZeJN6fhc
0W7IXmX6MEqbaiQtLKoaVo0FGVDmUkKJShBQAx2qOCg2gFXbP6KMOUEtVVL/+e8t
4JZjlfNOLdriKEo7p367jSSuaYpWe9g7YqGLaIwOzKJAvaLAS36CboaJFfinZIHG
QYP2JdHRALfqvQT3PC5+R/1pX61BvTOU3MkVL/lmKSToRVh59StPNwV1b5kJwusn
tMm1DU+zN4+QroHNP9J384WsRnNS3Y1iUR1Bw8bDvkZrkVww6ef6aiz8Xj/YSs31
uFNZPZtYlRlgs5Uy7tm3g0O6oADIc2TIapBNklXCxb/AcyxOb7glQUVuvn1H3Phg
zgEJm36MaulHJgrJamERYOcyCcjHhPIHir7m6oe3TrT1AbvlJ+YxFJiQiQ9DGPb0
8q6ihplsCgYgAseJHfI/dGRuk2poAHfXW18xxNAuufzBMGcL/u47Zgexq7AHX4Zt
7guIw0E0G4kNQBKTTaiE8TSTjevoWI3MgHGFz7i5imJMVd4GW1RWD5CYzuuPfVNG
VvbFgLEZPbprc/5sZwKoOwRNP36gLHKHe4w6LcyiTayjF+H6qrulDzZFKnjsPE7U
0cp5wk8YMr/mK1BVOfG0GN/D+IP3IomHI/EDxDCVsV/n/P0nQDpzMq+hXMlHRLpq
eDIL9sjf7VB7x+1ToQlM3qrjV9iV96vhvQ/reEAmmTknW6uHB6LqGkmNS84Er6jn
BCBBW2v7fjd8IQTaYiKninzGOD/szKluPpeuU/gGWAiEJrFidoWlZSSHcR5PfpQ3
fmATod0JPipUoo8QhXYHEoeX8loFAJdjvsOkXWCGWWeItrIPfFXt+ReURh0gNNw4
+h1yQ4iVSHlhSAbYUfZmSXwbboXMnR+xX4D3zqg6y9iVwVpNSTemzKETBa/1e+P4
y4WwsxldbFA1C+pzxLtmggcGqBOPOYCsG9g4CHLenVcwPv2BhMX/oThGoiDqQZoW
coDcIYft+FLFMhnMqoZlGcGag3zaVINymBh3DssTmKT4kpDtBsYOeq6Uke199cMt
kGLRAJoMEcKLngE/zQzM3Y/96Z3JKD/xC+h7obruFd7B4HkLVOOb5dEDAUYxnTpR
hxs774Rf3qu9+illYuy38jjWh4mjAaVYYEYZHVZF9h2pdEIuFKNy0PSQSwZCw0qR
YMdiAVrNbVQtg1yBpp9jYXWY5gUNUCOKSpfQqArpITm2XvCI+opAW7e54Rn7ROzJ
+CcAe/Xr91bMu/bC+cGTQ5QhraUfrs4F9fMngxhjeY2MkrAHF0+7V8r00aGPFxxR
476qovhLSvLVMayRwtdRjqp41aO5vRYK6MiDmQXno9ffv6bWjQIfMmzoWn+5AROw
Lh9SxQ8R2t+Sy05v04FCc1vcycpTIBgQCCWFvdviZ3EfyEphTibXW7AKcktNzPOJ
59E/jMY7k0rkX4/eBXlSH3VMtM4nxGmdveMgC0FNv8hN8prKK3zKVWjLZQNFJE20
+WkzHCw0NDk3PoHA8JxPDM2NsEYgR59FIVFwKzEuaTIn8UEVlhlr6TambCtVlPWF
VnRgae4ufJnOaaWbnHLGacQ50pj7MoYeNrEkqmbzqjKDs/amM3ftB+WT6PFORQhv
kLd6ZuXPetI2XB8p8zVKdpvvRMifRlJoFAMpiRvAsbEA8YxggoXFS/RTqO4PI1lO
iD5zxSVzpQ9zMZ0TvEurbxFVbMNk2dfqPd/1iS4rSH3KaPPfqKVT0C90+HEAuX/R
3vb4k7raZDKOJ/J9FGhPFqfOoZJoMImmXiUBt4W8c2+Cw246BtUM5YWhBI9yxq/R
UT3Dk7MtjmtNudOKXQFwKqPIluDpxba+A9St15PJCqeA41mA+v/dNsLXRIalUapj
J+cpwtrNhruKIXNLJIsx7UeMmaInw7CkEaWF9RZxRuoeopT9JysvuE0siAvO0osT
FOAz++B6zgN9SB4xsWJq4Rxg2Xe7CZm1xWJcKmkgpCKu35BXWPsqE0jwuM4MCSCc
e0qSwvqDPLPhJ61BByxnjCdBS15KvLwl/pIImNvdl3AUs8eYdHWp4pG76ggpvTNh
VD/kKpbB/3irMjLqyLLqG2DbFck/hqouNSGObAlR0o6IIINL7+zrgDy4iN5V1FM/
vIih/YZ+OFKXJ+HXdEteoW0qDjYNNQXrgkkq80dradE+XK6r2I9x6py+nL3iflBe
C4pPbqmrrbd3ljN2np+iabUMpF5+8yr2bwai+mTzkeCVAr4/eGFPyMgIUf6F/Zk6
3dK2DJAAsmV0XwSuE/cAvwabXY7/spalXLAsRpVx3a5kbH5gBkc6mDGBdffCmyK5
w9+yIV6mkp9fEXhZ4Epx2c76fW9FE1t/M3SNejp+I1e4OrRsNwYQD6FmhnoLWCko
+0aWKhZSQfOfiznnleCbO+QLOKg9bfVv7k2nR2bJZhJDK4p03WQ/6Tfg/8+kuCvO
adhPkdlnvL7juSERb2DycqUBsCMiOUDq6Tz6i0ZAuQ8K4mcZpjaXT2YdWi3bgHUM
bNVl+x3S7Nx/+lffB5PXjWJMnaknq9MkwHiAyNSsnbfTPkC7LbggB2efhstNJJf0
gp+uVCr3yX4xIo7U7Vmz7z/NwoD2umvxtknAiKmtyHfwMA3l061kW2xXlpCwGkCF
atBsj6tvWxu9v13fkDwLKNoNn0r3EwYYZe3I/EerI/xZlGUFTCCkIjRMssByEkRb
S1XJdV29QNdWiZmYWMAAJCt4xxsRXUkgDJy5qwElb4mbqrqewVhcK83xeRRd9vQq
0KYscL78odBhClfv+PlER9Ko3t402ETMYLpgNXVQPDAUD0WoAwizq0QljiF6UhFL
a9A0/RJ/06pgyfDJdKu2xxXskSUBPFZzwm9chg/Docytwf2OS7GEu36jIu1S+dxE
rgA0uGqh30BXvEOkL3DrQH1oxrBp8QZ6YoKTkaRCLDhodYhPwNnrB7q2DPeu7YhY
8xZ9yd3oXqyNaE8dIHXYzvwrEjoWheUKlcb61TYoN6SAiLOFxgnpurMR9CngaGp+
TTsnxy9EHcjq9e02oJvi7tqgq6AfzdRvy8P1xZvuIdIQW1Bq3Eo0lfBEUuPp/EjL
BiRRDEPFGyXLLZJ/lykXH1egxk2bbNxNtKh7kHLG0hMK5DHYbKv5IclJ/+8hTzfu
AWUhl0f1V5rgur/hgyGF6Mkwd226oiLx4jIudOgv2Z2vuirLvx1qRkeF6KT9C7P+
GBzdMOmYBe/Bgl18Nwox44WUKL2RBTD9Z8YOmfjZjYawigiIF7nSwIyxtn5L3WOR
Q3U/Q/jkzIpauthpwzhj5sCYIOdQpntYKnB6lm0SVAfAV/mRpNFd513ral445D6g
L5nlOkuDwxplFtKJqhV01giNHNMt2CKgBFScaO1hBd2xPOZGtGxboO8B5z6f7fkP
tWzAvaJtz1+QUC03lcEMx/zuaBmCxpWvnzh+7zIfWe3sPEitln0d+J7uZdROfVwb
/avP6EVEAUQBEWuHVbchst4OziKhEaFyXozCjL6BJkuAiuleyCLiWauWUqEbPCL9
0naFid2OwUFHO0jceQuLSHFpQ4ke22WhEDfR2Ee038OWaqPyz8tzbQr9OTopxkK0
HgIrQ9XfXREQ3FdT7C6I3mdndAwhlvqgW5gaD7WELK/9QkyWdSxTkxj81IFHDyeV
rN37kV6xz+XlCpJQN25VfzyJ/QrOuuJkHan4g5RLgUNNVMRTzi8oV4F34A150IqO
VxvgsjMp5KEV93Q+5nf1CqDMkKU/sWGU/Vzb/O4yHC6Occ/qDu8OvFjk9vFQbpe0
iNdKyx65MAM0t6acoy9mikJxDy0MgSGiJVLsqcqzVIbAhD06GriIdzjKcGZ/NtnI
pssyNUt0bmRm37N5wF1ztD+eJDa6Jp4Q9RioQcgGxbTAveYGHuhVkNl3W6uAP0Z5
8i2Is6A46D3mdIdhFYhiQx0xQhhn/6lD/BCft+EMpYR1hKnJvJzzzChaEBswQZyG
qaK77j/KXDU4Lpg2qII0OLstWLKgL+nGBWYVXfHfGiibAl/fK09ewJfnDeUjpYJf
+tmFHccaUTZiqMqcxeV1l2oYl+ia24OKiF09uH4dO51Vhru37sYanrNfv5qjgzi+
sXNgDhooi0AX8qcucuF9gulybk1nGxtm0pSDNPIy1H1s+aQArA6GQX7xVkh6roYH
jH4VvhVUxodZX4PhcjzXkSe4AOzL+S7iXn8INCoTOJF+0nd5ZLO5qnPi1zHU6H78
CvPFW6SvC8CzO4FUnm2TQJ1dVdCCzWXjAr3t/MTDJ+gei1j/8aH7wKeQN8uZd70h
u4/Ns0Oz1wSo+vJSayNz1scxcd0Px51WWjOtYNP5Ki/MyUb2loDfQhxdLbECJZJM
vdjXlW6fTKFalv8aM4n1ANuKI8p3TFlEKZpXA7j7VMxnp3pLNbpp1CywUen/sIEq
9kSAhkF9+1IC27hFqBVxWXRPIlqaZlS+R4Pl1/ZividXUpNkZi17BmYMaSFplPNh
FUYBTTLi46FRdnf3zOuuE+9IKbCWmJ8K6VRSxDg1aZWRGEBkgh0kzqykX/87AZBy
v+Cy5/IL6JH6dxP3k3mjbpLN5w248YiIvDxcQsX8w3ryaaUhXRuLmET4a1Vjwr1v
0HEQmhSw9xfeL+bOqwv+rg3oBj0G8iCqvJDHTdh6nA/4GrZ10cTPK0QuxE+tcKgl
OXOoNdHeDtaD8977kVOtrphACj9rLIUIQUZRVhgPhBcvmjXNmccoYkPEJI4yVr7R
GvWTUSnKgeRrGkwOm/4WvCQE8VlbPZo0LVPW+RAzpQomBXumR53THye80BKIFN8T
TjnwTYIGZvlbJKxsngMYlrV9OPh6OOtiqickJND79/fUk8kz6SFKaM5tiqUa6jg1
C9QvZSUzwKdRkmwd9P2JLV8swDKEdc2kwxQUK9Ors8ssUKtaGfg4aX9J5utog2AX
XZaadsQo2r8Iv1zdDdQ+w0KXiKy2LJ3eDWvNrNRJPp851LV+Sk5KCizJbPTLDYqz
KhixIaaqIM6iGtKPdJ2uOP1hC2FBmJRqW/JwLWQk5hmQX7wTBFo+8Z9co7fmnSxz
n5C2WI7dAJbLfXupzQ+S60P6G7ZpfNhGircXZzJk169BEwG17rbwlw2jtKucjolV
i6hmzL8oCGhu9RX8U1fnCxD6KksH/Ctyo5ERGNgKHDnN8zwbggJFzHM0QMfsS4bB
km8/GyKjAHovJii28Qmd4oD6SyWm42O5fE/KWUYF4zUpZFhM0SudvUGNnsaTkh1X
PeMX8WW5Qt3QNdWXvoAO4wRGidbrdACrN5u9v3zOSt+lcpetqRwdApELx7DxdiZj
g4gl73fbhRcO89OOBCVgEhX//FGYeYWes7rVC4HyUjf0zyudvCofGPhPjmC75sBY
8qLcsbbN8mGT2nKwwPf6mMvW6S3zK2CHAyvuAfMjeBsXXascLAMQxHPCcmoLKqsw
ZjDDu7WObbDz8OqJBxUZP5VrmXayqFzdEH+g8Gs+OvIuEuVUcBcHoSNZbIf1MGNj
hqo8Aw3FP+xOLBjcsfgDXbJm6eSbSVG5HLaCooNivPQgrZD13sYaRCDMtp8xKvME
zcLMVWOsNVLI4RrMqWbufG3N9xjDF0DnFV6eM0jeL/5lxe00Re/c4jwMC0bya9hA
XMj5YvMRh7rDfjej4kl6RX73MuVfGdraSaKzAzokD75fiZ60fD1JJC3TaCguIUOC
GQZljkvmb1XnBrGwBiKJVLFuueHm2unpoYrc7vFozPKF0fefWgCEMORR7PePV82d
MQzAHqXtpNFUUDIDq0mPU3pwBianpgkaqjvcXrTWYJhop9fkun8CNfM9Omfd+Bvn
RV0T1CDfvja68llizbldINlBRSD5c/hSCx51gVhcjotM4MxrJpsc4qvE3rXmXLP+
1gyUpIDh86yaz5M+OFY3f37O6URBLzUcHwYwABy2NTMGS6Is03jClLuPwOtuMwYX
yESFdpv2eeigM0Db4beNQhFjMOTYODhzwtpnB+3aKyQ5TzXLigo8sV6NHAsLK8lq
lUQPMCAH2DKLJgT4NDBf6nQMd+y7H4AfbmqvMCNsIMHWeOcACgxfrhpRp40e9aTT
2vogQXwPU+fqsnqXET5pT1bRmcJcAvAffAaRCzPGK9/RG2BFvhU6EamtTz05yf7x
Vck3cRcIQuT5zwnWMGkQtQcMDN7dtjiE6w+V8o41yCas6vrTKe6faEzyJPBUXkV+
v/SttDtqfFZ+fnIWlFClf17ssUYPPmggm+/dBCRx3/zlS5QTwyImSuR9bnwUfRhn
8CRE068FsBhy5ljcVNAspvYBeBHr+Jtt0D6RrTZ0DbtoquYQkgFbDthUXgDkG76e
qZyJr7DfzQyaQuwo5jEFXIxkSFtGe76L/WMGab5JvQaoYgEcq3JArZSzKNqZWscJ
GItnp5YCqkr/HmAnbWB1wBSVn75nHBinrlZ6Yw72FUiQjlo3uhCA8+WpWel1PqHI
inc3D6xuf2SMgAXHiy3t18ir9KJ/cntwV2DacguLBWtVcNfwQnCYZ70H74YLfV9v
44GCM3WG6Zm7jpq4jnYoeolcysjRa4w9Q3FeAQDJ9C3zI7Bbr3OsFz5LmvA9q3nV
awoHI10XhB0WAow+zDYCE83aHAxVNxtdFSOIM6+zp6ahP8VGtkM0GuT8lGctXRBc
OFLHPBOLfBF038NWuU7yZfetfvq2P4dcqr/qcvlferIdYXgHWvTpCBuilJQGY/FS
sWSX2QrBLqFNeWUFSCbnL9QbWqY4pruzVgJzsLEHSGYSC3Dz/a0fBOy5b8HIpDT9
vECYeyL2SaGc+3dXK/qOJB0uJgs3po9uwTB4oR5N8a1n3d2sp8OneE/X0th4e1z3
ITifiGjvatJagnnR4HufXQOuStIxg3YHGEue1f9uqRhuZjhsG91yQ1RAikg5D9cl
EpKZ5ZaCCSDyMaA6/lFOlJLL33OrEeWRhu9RL6Apnf9jtTzh747p8xO1uxkMiD8w
G65T3X4oUQB40AWh1wXWlzux71OaCrYlsfi1sqQ44pr/geLcrHU3GYj2672JBjXI
mYspZqzG5FhMVJmIltXcSb+7CenqiB+UyoclcSZs8KXqR4ynBmytjp4s4KBccJ+/
HcY0HxVSNIXemJn+yOMwhFtWR6SqBHnKScrZyKK0CjkLXHSj3B2teV8d0wKWo7Px
Gy1I+82+v94QTrzKKzhrEu79kN36TP/OJVYSt92YAxED5PtCn/S/yQrRmJ2isWuP
Xt4zaTMiujFy2WKQdtbvd5th7eVXQ/6suaOH4B0+mKSQ+6MU494qoZXYAjUZ0t/a
0l04NOx77pySqmsv1nYqNDkRSi3rQtz2iDlnuxxueU4q98NzCcRC1BYSZc8oJKdW
Z+PhICZDm0IdI61r7DwuAfB8cNf6SPk3n61JZYiByngTRYGNkRrnglx6Snr7bGFO
v8IOFHWPayiTvqlmyPZT8fuwk/QDfiLiNrebGwRhuQ1+cYrUTEVVt9af4vqcbNdu
bJTwzYYcbEEj0Fd3H3tVbsgXcdkAYHYInpN815CJe25ueaMwCNDeNcvNW6LgNZ4z
KZ7M58eU2wS7jJTbjiDEzFeoWEQXjbNz09/6eOzkN3QCgFgOiI8A1IKOnhX8aD3F
R6fUnmlgvLZdFTS/891E05Kc1uww+t+FS+kfHA9Ak/XoTO08HJD43s+Mm98Vh1cv
V/+WoujyBDZaYNDwOtNuMiTRKV2ZkcZe76Lfnny+qzEUfmQ0TVFHHSr5r90W6WRF
ON3wx6jffi182CRyYJ9rf9rqaniMX6z2cK0cLdrHooaqq0bmhaa95wJ2QCPSJgV5
vkrwWc2X3s0ZXOiskMIWzxRLbT014o+BbP+OWYyDe2YqQ5ZVyDB7xTK/7FM3e/4o
s9Q2/cIZ3k8qaF1eZT+xnQenQtGAo6Ne/sGdkNR56DqL8XbfYmCYueDRFlqmoVbz
zlL+tNFuOYaUdMWwpO2ttPP8RVVU3U4r9W8jTjPfWur125riwK6nQVE6xLmrvsBp
QK1iFkv3nrwsO/01yZqmB8//wxqV8cxBVgCOVy6lncRdPAXPDyhVI8cgpSw+oiUl
HovqA/gD/VfUBu0UT1raC3AwGORq/ng0KBPEqPTM2XSrdXTkLSd9Pr+BQ9Y0oOu4
pGiuujYl5bSNoBSx0Oud2GxLGCsjECMNlkfAMPUoY1/vMm0dXlJOnbEOs6j2eYlh
kVTlvPR6qvJmr2RfRVeSbgehRDCmBS7RDpfWDOY3Rn9wYb63eIEZpletiwF2RjGy
nqObwMLh2EK3eKtA7ZwcButRpC3yRIuTlGSERjlFajeC7Y8HXRKeiZZ3atFfIlTs
LI8SI88C54AOcOIS/waeK3TMsxtWUHLIGxmThl32PwMrc9kFvHiBXOafyZWEgfZ0
bIpO/spXh7Xy2mwdUxnlY8myXdyyeUNVuBXN6Lf/EaDlmW9vZPXDf+xYXtJ5cfzx
yYKUugN+GAMnY4fiKBUPkYeOEXMqurvPc9hA7bOyRnH3tN52KKrhmTYMXx0QhN+8
fEUTGKNtUhQyXtV2StayrMuett+OJHO9AAHiQzHrNfy+Iipe4EuYWL4IrjyHIc2w
423Tvuq7pAffgL0PtPkTlySH/Tu4aeqgG2hTpdM7yCsGRWK5eYeXkRyzSOarci8s
yTwIJlwMOXN4Sjz6+ByyPyuZBY681QmOM842KF+yQb7IEKXrQHj+KDjNu3v0JvRf
WfF7+wIXJM9NC6mabHue/sKAqLIjRVpoteprapremzEsEfctfDYRxRjYf9jomZk1
aK/4tUpXwGQ0jFaCbmH8mqZ4sI4joEgHC37L4R0hwBhbHGyzlK/0REgAtUM094ck
XJFhMAWkCWLgsf2zHr1xN7juUyJ0PkOpwyaPwjC3UKXH10n/nfltqbW5jr3wfVhX
IvmuqIsU2t+8JkYACgH5evhy5brRqlAtjsAEt3VAzguOQq3zkpyXkkYO2MdhIFTT
8+Ll9TQvtqsl9gz8+wrukNSnL6w0Wc52D6epZ49plMlzDPdDbrMP6w7kLMGaN3VP
n47KzpWx5vJCkedZMcuI34tzh3QyD0FNOsdf3vg0EcJf2wM6HF7vPv5LgtOert7A
PwZkaYqrHPdmKPoJRrFCnC9ggeJG4HFnliFI+H5KXXsCAgLDJdc10hepvxniUUlR
C9CdhbsnsEZKcDQAFWqGJtSUJiHInmCFVkj6ekqjo2fb6B6DxKyK3mk+TPKYXxxU
KxiiZJRKXAdGg7rHAqxSwcS2+7o54t4nB8RczGtfUykPoQvRFBSbTGylHRg5k66H
goXm4kV4lSEgrlI664iBSdeSLGamT3VFYAkxbl4+2doRAWhitycwtX++JBZyYRpk
tiJP0OXS151D5+xAlb1KCKy+qG5OeVSzXykDSjfhdcN3evwIKCY54IKBoaaiTYSO
asXprBa4GHioG0uAvGY0yLqr+SDnSY8ASPfa0nn6Fstk3Jgl1Ub87cSHi0s9k2Ko
6uwIM9X9bxNIvI2nrisrB5al/2Jw9+LZfdYMpvBTydFW8xucLdPMIpvF8rdj84gR
lyIu2Cy1I9i97eZ776v1lxWihu/MgSXBSGfOW00pjniI5vsf8iLuyiLNGqzNwkYb
0/E+CcltpcO/amLpPuzrd1XeCfM0KiYNKgvjAs+Og4auUIoIs9qqManIrze77zSz
tjFZ0uOZmY5PjudW9lx8no/r0cYdT9RQzkctCxNUONkqCsHhCJ1cG7wB5vJtyND4
n8qob0cRA+lgu2T9vz/d3qCe+wWX56/+957p0u2xJCFSr7DOilVFa5Lkl/hFNU8u
mcktISYFlMmjjJQOrkrmVOci/mFWOBu+tFd7XDQ7LWZ7/+eHCa5KciOdOp53sSfc
+GvzT5cMbODZXYyqDjTJR+fdbcceJEENRF6BF/z+eaq2udQpSx+0q8JLUAEuxE74
SNhnKxm1gPEHU3crOE/rm4zQGvh8E1T4TTAeKTKaY/9zSUEPxsHy5qbp6CQZDpvP
JwgWPelbkpdp8mm/xkMb/QnQntqqKdYmJZz3M2hZ+4VdLH1DtyYG5VQwDXsfOffJ
RcUegkub4rHcuHOwQ0I5jsrIyC/Ho4dR5Q4n5g1EMZlC9U7vFT0CiIivpH9Zlrlu
vdwviEE6uoMVcBKx589hzUyC/hD3fSLLRWc7oUz5Mzwj9I6ZQK3/zwrorFd1G0bJ
lH+F5Z/GUsbtmbc+LIBe/LhVU3LhlXqk7W+WaR/d7+7qEI008NUUKysmGzGOw49c
TRdEDLEncwg2jAmKMkQqT35G2ASRDyh/Guh7OgABJLIGa+NopPb9Y/5wos4HH8JR
hrtrBjFgZxrxzgDGeVsgJx3WDuWHdjTeenlWjvVjJg4oUiDn9GcTJ+lgnB7ErpP3
Yae2oMKLI1Wmqc4MxaR+K+J3kcwnZ6DVgoNVGdzSxbGp32ji9Bw+EsStfRmrxhtv
AsPxu+7mySMcnskCFCRJWXDT9hxAxHAPloXXbSTmWMyiv4Yo7gKk6+5irMlQzdy9
qE8M2D3sVpWLBjSzPkBFXdBg0/gyI/cu2fBfeSIQnxblZT4nMB/Ac7tDDT+JOcO2
vIGkANpvwiui4n2QrpwmmUJNcqyw3m8U1C++2ZKBsTLQoVq7xhbvFvj2yeA9ZZFB
TKwKi8y80nCHQ2fdVfW0RcNJ1zo15MGUi6WzpkAzIjqXIEYfZIZdbf2PE5q8pAlC
i8YRc8yLz8iVd+iwXEQnI1bauZVUOhqLyDShdqd3IvYYvpZ05w2ih4wXeeiFTiTi
alAa6DQoFYqgiYSB7QKHg5XBOT9FmRVocxrXFrdI/p+aT1Tnb+xqbEU7tT63mZOs
Ht5AGDHyXvXNPCivyJk3vScgHl+tQ1aFvpm9gYoSvdnlL8kZLkiaXzgmmxaSOAXJ
etx3dCE7D6bxed+e7NcSLsBr7W3SB8oXbT7939ihC2DeKVBeUu309v/JrIipRcCa
mbVrZ/cBrBq/HKvh5gT/qrxE37qJduuaMOIgBpQ+4Z3F1mMxtDKu6NI7fZAj9bAH
Ya36tykRlJcMYpqYFPu8e2/i4H5FsdU++Cnwn0T3j6jlOPCUNlPKleNjwg58lonJ
/WwqAPhmeCxt7TJDRiJw83lMb2dQxYFH+p61KreTk6RGirgJgLCEebazqkqIAjcG
J5gvEC9Ki7F5zTBeKplvAAgvh/SmPuCCvDqJSs/H992Hxsg7Ic7a0H0EJfYXDarI
nUQq1IxWC1YPn6OGvTV9Cm2rYEdXzU7sYF9NGEwG07/eR+DHl9aEC6K8tnB28U/8
KvzNcxoyqmW6BAJMqwtIXwzy+ww1WZW92Cx1L9jSnW8+NgkxKQ9/Z647MAZ0UIy7
gP1lEKng0bi7Do5S5KN0dqyVvONejBn8EfcWIKnr4/pJOtnnHxwEGxWzgO5ewVbO
c/ZXYolaqX90FSwMO6OYAsEusrSrxKJ3rS1RZ+uXtJDp+HfUXSfCQ4RAHwS2YMdg
25hVQW6kyOn6WcE/2I0A9RbJMwJ+IddTzEr2c2AMDPg20y8zUHTiSkZEwunKAfO/
yND3uItWxAlrBKe3OFiGMR1dTS1mSGhj6UyLMcBYWj+ieXL5FvUXOvZrCZX4MyBR
7SvybvfqwaMM0Yt+LZofbHlKxLjAlfsNQ8F6v9VWrbnOLUCynbipe1Wbe27qm6e+
6ngQSH/OK8v93+8QcDt7jfYbhXEKJanEpvYaqe1pf1PKtcz0JK1VRoeZjhrtTqU/
VTZxOjGiwX+S3VKfboweMEfdmSYuIbuKG9VBlkjKIpjFKN7+2wjErfZmzcGmpu0f
W9rZVMPFce3TxGl7CyT7uUlgH08+Cqa2bfA+cGy8CWtuetn2o6K/DFLuaA3U1Y6H
ZkY3Yyuyj8+ceoLqMXft2eyVo1wmPzcHmjf86bOX667RQB8UE+Ds8e4b/ObdPEk4
lIL5S33IW10rokE1dQmJ6Jx3I1snfWwrAv9GS/fmNARrp5NHHcn/5eXHQCVOFYdc
vPx7c3wBhzAK3V+fq4i4S/SHxW1KO+/73pho0dHTbRVc8Z3Rhc7mD70/XpM9V4Tb
2PcLe4+a5SFWTTwD2En7AYVFWs5RslbIRMmTuTFtEHIgifOfJK2RYQh2IcA+LWAm
NDfYsDcI5jQzyJQVMA/GfHsmhgRA7BY3uOQhbrdnbVrwzNZkOxSvwPvDcifowtEp
5nTnIlCeUNYA0h1J8I2kCdFaSLefxNf+t+hupdBzI3dGH8Gx+AXP5Lcce+vsepls
UtVBnlCyN/279KTywzQOmtVMxhRadoq7rxQM3KpMlbICoMUjE/0Y4m0OrhwJssj7
KhB+wm4RD9/VFK19bn7dEWLpUwFA7xyRmQt+7xRSpvasCYLW/1gOTWZWi0Y8ZiTq
7zkbPEcy1FVU1xBM3cG/JJ2lnyDgiDC06XgKhu+E5i/ZlvPdRGm6Lmx9ddSG3Jog
YXNemkQ4Z55ds9vFaMoBuHDrXDEoOrC1om2u/pAR2IMtPXCjLSjZ6PV4qWKgUsz7
6YaM52lBIwWcgVX0qC9RSz7Bev/ZGzg+KSY5CwjRZt9TDbrT1fT2K4adGsdgUlf7
e1DQTkJ156OU+Bww/8a5losqxURET1tiba/04ss7OOigqDWDSmQ67hh98DewNPe4
XqmhxH7yr2+KYCySfemUcgB66ITaoeOnH6qlrXxRx99wFhDMqTCDYzycToLEPlqz
1UiW0HCx7hKTcG3rjwoK9jreO/H0mb2iT/ik/DHbS13a4fKbLOpp2t3urKeSW0Tq
1jN+KX3BKWL/n2N/uVHc8sa458U5dzynes4ifvxXs1MSLgMByGo4WJaHjuSzHqwB
tT6P7yJ7yjkHmh7VrZEOGK4CyCTxcNfeOc43w9LYOq9rSqiI+lU4suyX+vOTqD5s
PezSFIm4k+76UMBL2lwllzpllJoy8gHyvB0B37p0LfmdUcIiWg3MHTZ0AI4VraSp
1cCyvdi8zgqRIfcqlG6zae/8XH/3GkCQHe4dy2BR3bgUZIhfWoaqf2v2ySngUzaX
jWn2LE9v08o55UgMJy4PSPhgrNWqkQD9dcEZ6MPFQmkTQ2TdgIZbwJPvCYR/Elqa
UsgLdSHSwXzX6teyyxw0dFK1EP8GV04NM+eHcPaYY1ymQ/9Dler0yshcEywp8HWw
KtXwlvmUSLOXv64DtXAffam6GAop3uHSI4axMhyJTMhWI+rM6oHxbSJP82u27Nco
7kXIURS9fc94T7HaZu6PXi+3lzH4uMQXV7cJFdBj5/WFh3ajMrlRJT444+Z3itXJ
Ir1t/D38zkAJqQPbiaCgKvUdJKtQUrddMw+xqx+bngDf3LiYo0/QajGHju/agre0
oi+071B8UlkqUIP9etXro5E8WF1je8kxFvUB0nGS7E8p4mhVHBkUbapweCz8AHol
Wc8TO3/IlBDGcT/+W5w2DZ7roh1FZTzwMdC1rhB88/G8hOqGJSkFgRHX8NTk3I8H
KGjqZysYJ45aMZ0Zo3pgQXuzY3SUdRIfnXw91Iic7EYSGSTIJdb8aunSetriYZM5
EQP5C4/Z7P3lvorfLy5k+tTGXJtzflI6dI2o2KdUe1EGjmY2P+qRwiQR3bO2vdXJ
cvSRlJekHCMXhovd+SDe22sApCRN//s2frqmy0eyd2/48/zf1s+/YmEMbF1DKqri
C2/aaQon0JlU3Uqg5nHhkrxvYw7QpKiQfPBXwWYPicn7RKWRPbG83Propd0NBiYW
KO2D1+Bb+49KvEd09WTDPvSNrN3uptEe2dBXdrIZXwcm4rkTcDKkmywMRaLcHzNT
G5JgwTBnmcrra+esY+XnPB8BTBlyYQT44GJ2hZSdXUiFF3b7ZJUrCk/3ob/lAMip
YBtCXMhWrU95a3IyV/5aakm2TqlQcHl1WKOp1Yrg/wX7XB8mp+VZwU+FuTPBrw5R
2XDj/Pl6zhUJquqrIHMu3UN2pVElR/lqnDkvhSNmLvB3f9C7Mw8BRFomJqSX8M/7
WEbbRil8rDootp3hicO1RvKM44K88uaNzgUcpveTztddny8ftv6jtQMXv64I4hEh
rFbqhu5coNFXtWTfx71GppsSnjHowqheH7dO0LPY029an+JsNGzWBNFDfSFbW6KB
iYpV4QwWo1qcyvRrGQDxhWfv3OrlDSQHc5j/WzB4PPOgadwMRFrstXhxGkR04nBB
yMakeC5llRTrvxhcKJ53nhXlELt+/Gf1Rn1k2utBP5/sDEpzNvSeENk6w73b6HXs
abEmdNJOSGCQPhytSMeI3Den5HS0n8kbgom0MVUZtmjH9osx15WitO/zhECBm3yC
Hq7+aavUKjtaz5xIQ6RnsKRZoNzbWUwKZ88Zp3XB+76i1IRHXgR1ucptjpZedcDV
2pBh11K04VWhVfo3NmejGwgebQZ696V9m3QKycJvjB8mGGEPzyzH6krtRm/xCct8
wC5s/rH9+jiyJ8tRTNSLcseQ7UbgVcHVlVJmYlp5du8nojIHRw+DU+1rQ5uJ9qdi
yZc5zKt68T0ftrAw2s2ZiTAuQU2IRQJkad693qDT7LVi0luXVmkq1ApjZhIBPbOu
T7RbneWfY2eZ30KQTfAai9vB5sPB4A2Fh9WzuHZEJT7Q+JYy4zvj6+qTvIeXSsq6
1pvjTmYr0VNaWzKv+XVLR0/vDpfpRcnSGqRTTC+4igw4YUK0f92BRW6FuKvct+yg
xgwDIwWqHH5ZHRm+4iOk0462XLTrd0qFWntF9uujuEdVVJky43e29Jh3e9Um7oHY
tIOKsCLJelwfF4Jk01NioedlOWG5LdBlD5JJi43fy5yUZq8egB2bSC4rGza3nBfn
jdGFRcv0GeQeblwlbzp1oryAyCyh+NbCXJGyl7bKcZPbGkWYg3Fe8cDk2patbIIP
dkZlAakjmIoB/aZYc6eKXsG6M/vX++YZVEjNpXRqi4tYQxJRFT5YZUMKOXyGhzSJ
OsVheuZ6wOEX2UzhM9R2yzs1u59LjwgY4CBFlwgQE0Ip07bLLbnUdZ0sSngfkFX3
N3ug3kGSybLFG31TchPeg+sHuZqysNf6PJbcdxoE6w1Krf1u+CS+peEr8y1xSKoA
2PYJOZ3rfz+CAcOcnMcHw84d/8nxJQW2u9pE/Gdy6NH0UwAcPg4MQxgtnJjbfpaj
8l66Q6vd37x7kAxIyTCr6OCe5wW2TN5+1tN12oJIjJYSkiFSphSx4T0Lz26zZZfa
MUUhiQqYo74A2CTNq6BRDPNJDP3mkzi9Z0+phbgdTiRsL7B2tGS8JewmDhF2d3yC
3PX9aqquHoeiMTA2YW0TcZNFXsmYdC4kPw3bJ3CGOhMJE9rY3IEjoTEBKYPJBqAg
wFhjmkuFF77eFEO03C0vIvDqmI8W5gcgYuXTuuV2Pas19ijNvT7ooxNWelqzvLoU
O/1kU9SnY2ONikpkWwYQfLKr/WTHLMVroAfxijf4PBr6Yp+ZlbEF/xF7+z/g1QT4
t8UFGJXwvkcna2BKaTI48BkMt8jq7T6CAhTl8+kaBCGsKcvYjP1yZ36kTvnhcbBh
hs4ZS32lSdbTGFc2r3I1Csxdnq2qbEfEjNg8MgdNtvU91ilYd7owZNqaasFH+kuS
SfV47ZbyyrwuyigaGBcFWO4KwuD/m2fFeCem/huTq2KwpI2vhW0ZyxFI8yO2gR9c
eB5eNgl+Rz3Aou+qd9V22aXDKCHuWvN3mfZgLWbSmb/4vtNKksygZ6j1CQsCYdQw
dCL8YlJM6m2VyWEROUp6EHyoqPXAqpjlaj7u8bRr58Vxr88UVjWH6/iVTKwox0J3
/pE06vc2Rs1qWS7SkjHUNH+cv+I/YDYDyPpc6Mq85UO0Vlr6aMeyhXLhs9uY/ibm
gN6YOyLx1/28A4aFwWvGWpIatWvSnOcerdsrzuPJXzKP4RF9pYVc5tdt//e+/E54
GDfrFG9y1yeT2TbExYs2Cxubzw+1/4cMZDMQ75O3KnNghTwvdi/8OaQi74jXDygG
3ujKnrVTH/P4cQdgTO6UHj7QZEj5QjfSxJgpBh9X1BdK/NtGU7syzyrb7rtrGXd3
pSefwjmqcKML4IMUsg5JEeMkXDGGwDxkzzm9vUntkoAFlHAyAp5+jS5cX5gXFTku
G8nqd3x6uvyMFdCOnfZ0gPl4JzGK7r5v+aMP0QoqnXgJzucQ4FOT7Ma3Q8/J0Prn
snfdTRt76XIUfOqR0yuiguTtHKMWY3aFIn/HauS1QDqQLRGwY/PI4yEsCjUiBa3s
GXHlpbFSiRuuKgF0rurw9tFd/yPSOOtIezoknQo/F6YP2cPmaeOK9njY2Ljw8r9e
LT/EoWNy1GRu5HPAaegXt8dteA50TGtd+F3tlDsB1u68cmgc9n2HDDpnFh28nYC8
IgNlBuSlolGSHOLsBzy3IuumwERXWy3GBJZjyj7utkDj4l5swZyN/u+gIXJVV/TE
jGFmNznNoEqYlClcFl6MhUT6ZUpbuPEdgfNwjSPWctJTxrLOiwhhsxuOAgToW0+w
9Eu+l/p9XH7uvWwIJTkz+sd79UP9D/wTf5GSzTTAcGV5ClGPYz/8E4GHM3RCk4vp
Ww+lqW5EgUhKgN4DN8i+Uy2Cx1rYmZndauRRfkJnTBboyYJQr04CXke9jORGewQB
h2MqZdZgxVfNNlO8vhzyALmPLZkEctwORzc8w+csJ4/87ShU/LR0TJagX5a8JGSW
O5uSm+UyRW2w5m62ZSJbNUPS0E2ACwy2kY1sHRHGTbLG7HpnbIjc6agVZgKedPvK
+7Kxi4V33GCjHMl0fsZrbCPxlju+3OuCw1I+FucUm34FGPBwZn3E2ThQAlr8ybbT
lL4UUrwZaPzdugSOQwgFtm1X5kuetf++6L5wwZ8JzF8NXsjbuFo6xgB0OnoJbuJ7
qc1umu4+g0pL/XRJw4psttcwDMMIZx0V4Zo6PObYNt424MX5PJNbUKeONH2i4yGF
lXfXE6UUzH+yJsNX54dLWaE4sEYusxKvIOgk77ZTvAYVyi1AVdPCD7lhNJI5RkoU
cfTYKpJnEQakI0BpozQTV03ffUwWRXbJa/1vrT+TgHelr+SR1mhqRmp4p9lfHtZ6
09s9RO+NcTo/IgDH5TCBJkQVgo7kQ6TL9VMLuUGbjCu264ZIb7H4GTI6maI/mMlb
D/ZMYoii+J1P4OOby+OuTL8mPiVVCqfo7/UkM6B85PEq+bLimpuaeJRBqMAwR62E
G/RL+4CnojX4rBAH06xhGRCjisHzytinX8koiinFMxRFtdHDRP7E5dNCl8BeLs1f
ZVVqybpSaLr9UtDd2KzM87qC+9/cKOSpQeeZgtajf7LktIP63fJle4UZgLERYeJK
fbArYNiOr7aPddKtFUULbG9mhnY2GkbsfbxGyjcTqsSARZOCExTd+0LnIsy1ezDL
Q8FqvIzJ+XEc/q+gL5cCl2py26NvL106WYF6SZbRbJqlYTuBBfSsL5VpZD8HkZBN
BDgcW87/dX/6Ri2z/IIjJpM5d+UFjQHVOCX69AdTdhPftCyitLmKuB5B4ABTKuU+
APRTodEFSaqazmHS5lKsoDsoGPJ3AxxCyDREzKpv1lPvf2Uox1J/NfC45WHhIgZR
bNC9+94+7bbkA9bmSn32v4QSLhN4uPO7EI/Ubx1QGjN2FIsqKgla776tVdKAe7DW
Ht8hD4HBxQ8PigY/tKf/ZE/zLsqOcHbNNma1zOF1HYp+WjffB31UIvYh+m/8n1u9
gMbxduxQBOeGphuOZ50eNVbKEBVSAiQixhZM/yzsIcmO4h6Ld1Eo5QD+Ll7qetiR
kspptwt8bn1Bklzl2DHXoxiDP31m0Q3AqCOfWrPUQIpHJV9PQ27Gl2+fMx9ZWly3
s7fMIEmZlK260/LLMmG+ObMsJq7+4l03pdyzMA7anYIDrEOnMov8lhgNwEdYtIxC
C+VVnW7PpB2iD0ImH2IGHdqLG48RMY8y/4uFoEh/5K6pqgkL52AZSyDm7sRztaFK
Ofb8MUPkA5GN5WSEQ01mxDs4/KZ2s423jTBw5Q69b2xXXtg6xrd1AbFp81vm+MN+
EOGiHJ6djT6Qg1A7PMx4D1FZH/CHDbtaE6PMu6EsIk9dmeLV0QMY1FmRpKPH3Cs3
WmgkrZLRIqJDlJif7dydnvsuFOGZJL7egTgA6RS0SvI65Smt2VFsrY9TMwLkpEvp
JOvmrWxSeavUr8I65y4Aru8l2psmjjlGjkAFL+ZIWRdTvoHxPn8NOjgvrwdDwjrP
/Eol7c0ZE0ISew+++E9pc1GJlvrCXD0VXi89H7zc+BhQWt8hqTtWZ221Xg3pB1FM
OM3uRiRHhmUMm7g59sSffStUUFKOTP4Ge6O02bpwRwmFXZ3q/7S0Z1R9r68CNGqF
0EIxrs76wf+apWPQkWJKVMHjhZBxzd9ErCPhCfBaL3HSS3WE1xx8NsxUTIhihr3o
2xDU25NxAhEdHv6WZtffvxzown62RE4TW2sihf3INycisWPTee9+k3ITuIz0xoXv
JLi75SmH9ZP8L1kI+506VQ4fx+Ce/fXd8s2aGVcGM4WhgatrqXhXWGDZVyoFjiWK
Mz1PHGaVoSatT1AgylAKf6JfrSdv9KqHH8mXXzwpnljrE8/WAWBIuR+44Y2tLvzc
3ZPy53emq3cWbCd5N2ZUYefQ7dunOzhpgSmQRnJM+H8kQy1b11H8Rnzab0q7ipY0
P3hXodKEU3D61zud0P2aPaEligjSKRhOk3w3VxWgeJBIOdfHe6M+qneDY2s1ZvEY
HRxVkhS2eBs0GhnRZ3t83Y9f2AOlGrsHcF9xFuGB4E7p/drXfIE+0sqdvoqJEEmv
9syKe2V0pj59XzEiaLfOEugkrGaPTef16s8EhhSGbXd8bFwRL/xcbz7Pzw1FC2fX
oVeJyo3y3fN72zlDAAO2z5xIbdqA/4mcJFZQCXVFSWYn9yI7cz/ISO0Bw06Ixnsn
0xUFfChOeJfKHW8KLwMV8ZFlkBWRoCYMVGVJIl0o7YqAhTSJAcueTicpY9JJwMlX
7Ciqqa/a8ZZ8xoasJ0nxKqj5IT3hIaipfWgnUUP4ITbAhJ/CRl6JZOJU0dxoNbnu
rBo+QsfooWaTmemgD/2N6jiPka5sbxwBXotgQu2auSfEfPPiFRltlgs1CoaoZ6IN
e1UkfEtdwsRVeOXrbSUPUxmpV6qMu2ScDrUKSpsbXC80PGpcfygurg0hd2ECe8nN
AuaRgPDforippDpfMu09TviBZjpbBpFQxhqG0mEdXpTHjw3/6y5kR67UxHMeZCjY
/mf/xyxmK2ftZxFtphPY5XvVbem+lPOL2IGenCAlUdJIDqBSqZCsvDmuKjYdB8j+
TgAQLpl9FdR9nTfvZOLfaVrAxrmiekyfM5mVKwqnHHcoR1mEI1YQKpvQn+hYKHxL
loBrxDUzirSmR2oeoJQvK6Fe7xrw/T5j3KEzQG0Bt9zwUh5kpefa1AdBVC7Ex0v2
n7i1EvWo0Z4ru1SGzAShRGrr7wIZ0/OqVt0pQ06S5sGHRfEuA0B6NsFw5J4mEDGw
RppZuRiE4WIm9/XpbywBUkcH4FOyLDSb2S5o8wGqlfNoAiin1C0bA2BfI8mmWT1f
XxOu3Kfcb+0FFQTgIIMVCkIhSZylHcefx3SIhW+iF9Dt5txiQEnLQKPc3a6blZ1l
tINWQx2KIfmiBpq9l2aWC3prwRMAAOReOCAVZoK8d4zh9smgI+rb3zgWhEslArxi
Ubd1wWtS3VCD/jd24MRUoa/pAO4NuX/m3PTAupN8CZD2/CoS1kJDZVgIfMSsjzww
ru7ldjrDw5PrYXXvJjLZf3PoWfCJCwTDOhLTHwTFsUOKwdzaORznwkTUPP/reW2E
1Ubr03YtYtdsYSt+JR35XKHciHaYu6kOKyfMgpb2b3kPxtEiq62CiQHPuCgCO/y+
LO5AMrBZWGF+LYnNXVo++TEfPLdy/EMxiiSJv1NwJsME1b6Y61pi80PoeDBHQHDB
BvFilcylp8ZLpOgH27l2Jflrk159LciR5FpFMrqEFTSw7r/yYsMJBchta8/74jz+
y9eU2SSSHrfTICDQca3fspxORvR/FkTVxeb4guYy5/sGop9sf7gSRMtjG3M/Iqx2
xeOZdfnmZyZHg2PX3SDqBRhifar1V5UjTi3RjLw42aplNthbjSUpKFPmXbktXZrP
9wwvYmiaWLrdW724ok5QtCZhNxVz6DxpXyrFAEmh4dy5w3s7raU3wyrpOQPESg3Y
iE3O8RPyWKfczuAml8f4FXFI9ZLzBC6Hma1GORwJnsLIF8uwhnE1vexo6omGSEUU
n/Z1lCcc2OeIoW2FJAaAF+HEP5GPPAD5p+mlYEqiV5eK7NUuP5HZj3Yw+UVzqmHl
xHjt4mA0gam4p397CjYO0rfdxWhtR4Skas0LtX9dlEqobF6UerUWPnPPJRcnhGxq
NCOfpTugmG+Ef43W8PNgSJdi5jjRYs+X9WPIq0ywyjX67dXW074VsVH+lxyghEPT
Q0mPW17OhioeNzRD/7zGkrb/r1HbjgC6GRjwYUNnP6tv5RXOMVzSXheYWgbEfcQb
JnKrDD4O6T+dwDI0Y/7smzG07JTGRIYBrhP/vR1ceIk1I3A3MU9T91jPF0L17qeJ
+2nzA+mgG/uP1IeDXJ9F0S4nxteqSIruT+01423HRpGzD7mpjafFwk5H76rXm3qg
3BAid6Lj/HLk6J+RIj9Yvk1NwcWfA+DlR9LjnBh9WgtYcY4fjL7e+0hK3JPDsSPg
Z40GZ7U5VQ/kztPBmfP1/Cy8G/N6S1LIgQ3gkqLHtPLAU289FdzxOG0B/04UU0WB
qYzeAdLQ8G9p6jxElIIeOSIlD20SRgtXJnFjqcXln4xPRHCbLNIu5r1U2L6xjfP7
Pej/Cs8HbEQQY1Qp+YOnp6H4m2lf2WC0IDq9LfyTlCRS0eQm7ZN+scXcDNlSp1rs
bxa6HfP5Hh+hWfhL1b3f07roLkdgr6rHKd8phYvTZ68Nnj58OcIfFibPsOzApGh8
vyh4NcTFWA1KTbWm3UhHbYde3NAGvh+avj69aSCAYt56DJXl6iKaV6S0UXDF9WOw
1I4n6cCHVHrRiW8YSU2xpkinLAmjoxhKZBUd7+MtKqNd6IV/huEW40b5Kvx1et2Q
hQxxPjMI6gIfcyWPUkb9zoQKCxllVEMxGbtS17ayajtv4eQmh214/SJWYHkhT6J3
0AC2S/9fN+vm1NAJVvTFiazGVFPFNuYxaJqa1IDtky3YtVdi7YCdCI/EmkBD52hK
WDtawwzMds0icBvJP0NdhuJVfM4skC++Uy5Aybbd4trGAMJ2hI9NbpvjGTHiK39a
WXYxY6XSOfMW4mmh8tByPmqbJX9x8QBSaDwil52St+LVzJdew4S7eUHPiZvflUNL
ndLUsBCiK6w2vnqoUa6OnfVFyoWe0Aa8rfgYgbZN3D/GO6YRTUTBtHqHmo3+LWwP
ch9uG4vJ2pcH/zkroXg0L8D062boG2BvGIGCqoLxRFGqmLaDW770kRnKhCWzOOpE
df9nxgTyFK+WwDjllWcNWDX74Fd8aekuoUkETQk8wDxVYhHRMJxaum2nvLN6FuQI
SZNOTFjvbpV5LmU9AlGuZAzb+ycaD/sjpHVUe3isBgzcKIWWMiYET18W4WOOV05F
pwSo04/6q84c9iRqyq7Cj/Bby+bI41XLNbX/LBox05ckY/P05gxTKo6DFyqaAcwl
aVju5hcjRHHwbmjz7+8YNavF6i4SQZvfnVSGEouICMio6pDTlr252f6VANxpzQsj
flGNzbxjG/N8SpaNKzjHE4tuNQiWDwgcYcLqcO76EVorAOa9UlpwMsX06++8ZWZu
XQFyOLqtmSyGwxi+Pz/xUxnjKT3YAzbELF9gHiTrYJ51w1wqzz6a0oaYqm+WGVhP
X3m3BNvKVLeZKG8f5d4gh0Nu0bBilProJtyK0ZgALJ1cgUQbDAuYeFOqBuh8qcSl
Ljp4p9IY3iNeYnOxGUPDxz8ob5MVqbq45sTDdaC5FG9IGscdEo3qNAs+en0rChP4
1gMmbeDr2nkWlepouyJp+W0mc+MBTK68m+39vbTkTuXTWWazGpxJ6eVoaTJJH7SJ
3c8XLLnM5EcOwiq6HoOrGqEOJjJ3ukKc7gCgSp/1Eh9ZDq68ZLUF+SMcVmoGupgk
rvMuxi8UOnm9khGQ6hXMSuU9vRq+3zZFPoHjEMNxC/HEcHEjRVrnNY2PIVKdprrj
yb2BS8Il2psJV+9jjHlE195CR9G7qNjTUMOYRr4W/yIeKxCzeqPL8yWfcL9WvNFy
TZ7wQW7xhRGa4W0176KCfqOMmxfvko1clmMX5eV6IaAzl2ma//x/wD3YFlQHmpq4
suDLJdBf6dy2XIlgsAd24x4xj8eg2EEx3Gjj8Lps/SynU6R7ouTZ3hIMGI5FKw5J
o+YesgyrqRrDyGMpJj+D3Bw+eY99FO57lClgxC0HGCeokC4ElLjgE5PMmPVBINpx
xzfa+PdFI9An94ROlDmnD13S6LO/5TskTAKCnG61ORKNFgf+Vjl5FdOEIqWCuNVl
7h0jCz6imPP6pQMaLPkfKBjYAL0F50e9n5VSvrq7x0D6aWMATF7zJ0kmqWQnfVH0
vrJnWMDkC+KLq3cnPjcOhQOFfhcVair6pokK0IyXCqRrsko+Rj1qK+Mp+usbtf9T
WUOjKf/Xn++ugephUqVCMkA3L5BU7cOCUe6ggjsqAjr0CjVDMWn7vhkl1zre8O6E
Ocv9lyKVhbPyLo5jKhGuiX5K8XFiUXbs2TrFc1cNI09vCw8bBJ+QKhpoUFzm/Lv1
2RSJE3J3B6rCIEJxd+PvrbCu4oVvEGbCQzAVuSjdDoyt2SA/SeG/+He+VYI4YK0R
YCqKYQqQ+/clhhv2pbqHrAhHPn6kmWxZu4nTXuiauh2hvMNloDJPh97FLXrH7bOM
FITSWAiDRiVq8yqZZhw3qOSPHeFfEyZoep8/8ED3Axr3Gjfh0ptN9/rxGySq1TFp
RE0bg22nDol+fJAihCHu7OdjHgw6qxvP+IKtVSpJ456hFOZYjjqSSDu+YF+Thl8R
iVBaT+Zf1MCE06OtNYxFbHJB2oFloIKGikEGlENRwBUCenWkJtSVTR3UCkthK0Ag
rvjsyv3orO6hGzFZQoRFfw7uL9HkxM76EQAdY+PysOYbGrChmhgsS3HJDoYl2mSk
w+TVr+24lYVRPNimCE0ckpBw/u8xV3IewOljIfzabAh7Tor9wVjrjVljV3QXd55b
RPOM2UFAmuDRP4XYChPJ8g7vacOYqxbKrO5u98Z2+yFjd0T8vVlY3U8Z/Yqi9AjZ
USdrfCxuGI+gTYfIhQ7Kp4Z5PCA97RHOka57527Jq7KVECk7uyAAa2UaP5lQ+/MS
xqppqDOLgcUecHogXHFu6xChl7ZH4eJtxBWb5/mgE77hqHA7FuX0di2JhhqvYzhg
qB/ATox2Td/vn9fbgetnGnvWPS0yyqO5ZTsY2PZpZ3BbDEwIQhC7bxuZRDtECnD/
YKWEqBb6ldb0pPWAMMNqv/Vu46c82VkGU9gzBcHI7goxVw99VYJjK7EmzI34y1P3
JPKvo8ZOWb8Qi0QhJPyx1EeU3hL+rsK8KmMpsCBq3nhWpnsM1sEQlgF5cS84UhEg
N1ouBXFDoZi9ucxn+eeDc4AHPu/mC5SOZ9fu/Y/Z0q6KmGy0q4ddFPHx9xdXqnFU
1x7ujh7rRX/LYXT7XYfa0cblQPb9Pp7I/ekJH0F8MND9rBsO0RqYA54EEcjizc+8
Ijyp8KIayWQoJDhhc6d0exIhjuaFMdUd8ddbtHSusGL+E1AtXcKF3iTT/8aczfms
KnQe4ehSNByvch7ZLMxW9diAGAfFgQA642TJWFTH+cnGE21o3VwkCjjJFQgTivcT
kP7/dJFLxKUP73YvGJW/NUxJe8vGvnbfYz390y3gf5+sgOygwHEKIpa/Di7Z57dJ
ms1xAdU339ryMKHiCYSz0X1bKr+Xk2N9CZ7ZmF+o/IPyAyaVKMX3izLgV1UHMyGQ
VinFo9ULeS09QNgBClF4VNY7ipme4dHtRqWhJXvH9KMDVqWe5bta2HzaN0B8xCeU
HJ1lFAa/N0RCQB4uzt3ZeMb3ys4PEaB8Wpep+dQbVeU0WdJeaBPPC3X8OzDX0np7
d7hpeZtCioOF8YRq5xiQkpv8bxDXkQ+6HCxSmlcnDC6HTwplQ8OvPwFuQS3RscbF
hPXFyoMScHy/BOJ50BL6OCN5FS7VMz0ySZaD0JbiKXXOk5rTPpTZx0Glcsy3lu13
Ww+jBBP2vMznmh/V8nbctwmMIaFurtcFRp91OlJVXYfYEZubDEZU+7udVNrAz6gr
9mieQJ57ovhIHkfUt03T6l6Xj+yKuRkZ3U4XUl5TpAitBgfgn6gVrNRvV/0wov6J
EShcW06reJ2G6KrqUg+bNmKsKViUMKAUGs8mIGMIN0z5kKmH8VjbYeLZvHSDy2XI
RD3QO9viCD7H1T9H3A2DjUwF/LATbIynAabMG53e7UXhe8OFyw0r3Luw7yO3YpKE
KfzWKOKF/0T1jXMPRQC6W91NMEw7RWVofyJwx3CM6s7MSZ2LcLhhGY47SERlr/yZ
ciX+Hbfhim5NJHWY73xnTZ0SoBDDxUzoDpLtZ9+x8uK6SnOek9YErc9Ma5T0jcAO
LjTLe7RKNdwIT81lzbatqCLD6nDA8sHWVTf3Fx8MCwpCqiwYV5GZxng6dgAWG64I
t5L4mHlMahVNmskSqfygfxito74z2fIh0FzTYJ2SkkOVtv6nsf+fOKWGfY9gmx6v
yi+W8ukUiAojvbymcYjmwNQBEH5723eJa/RLGyaDS96ONANRjvRvYyT1H34BwYAb
dk5MqQBJcsPQmr/yUAxjyVk9gNX4d8k15G/PF8aAVofA4G5AP1WzhYKH8UN9LgBY
YjRCfM/Nsot/9Oji+IEOsoepw701l+PRDs/Evc8cCuMm7W3+bdRclUblz3Me85G0
82PE0O5uuK8r3RMUTOGq4qYoy75wcSw5hE8NWAwyWRhddYIe9yCMPDWxEc44FicA
h2C7m2BGPUUO91N8AgAfv4oLUN79mB1G+mOs9D7/XyyyY6r5rAybvBK6CYUGqi3G
GOnLqrDqY+rGP4BPheRrZWo1xHoQpjuErGhkNQRPLK9h9emT/MiawrAzsRVxTAb4
qTcqtYDfOmWnW4UOIsx63PC0nR0H+wpaM1oEEz1n3a86aQnJ4gZZsS2OvfYklSgO
cv6v+wO6Jl5ZhmyMkRXwMjvs83bKHuf0V1OdW2fcn2Wxirj+qjcmxz41AT0u9hyM
Hbo7zMcPii9csxHjbRwBRI5K+XgsZWYw3bZfh9U32wztbUeyGtIsiidQ6OGYHxNx
Z7RT6DXQLj5cOoavBtvAG7SmPPpBXFhF/A4ubdcyWKR/FanbwUnDeUMGtQhAbPiI
dm1gvoEzic51ZEHP8QNIgTI+N8CLwQWSr/KQgRGaSiSnDlWM4lMf48zPNKfsdzfH
bxY9GjOLYWJ8OAU6hP2+xTfmVOvA5myDcgE3D3jxH9TGThuc1rlK8/uK6zTzIn3z
562XUi0kyD8QxJ1PaQWm6nMItKXtrTaMbwdnOGbfHypHtt9ak1ZOLvWwifmgjkLk
DrQaJHVcYHFsbS/9WQ3vaOrBnkI03k5NkMn4x0e46vuxX5xYKsrnwylSn5GFMSve
HJn3UgNNh28ppy7IUjGvwRc9whsYxw6AyJm4eXX8Agvd/CQDdwd7YQniiVsK47Vg
cbQyh7w6B9AcYtYKhMPT7mqY0z68MLe5/V5IyDS+DxarKneutvzy9ZUOvIpfHPNQ
dw9OTypzR09tgpXnztPMpHnz4Ttn5qtHRwzSGnYOCOn66OfH6kPdwpa+03D8xPZr
vJ7WZqlEq0A+GGDfCm5SE2hgjavEVK++yq5uBcdmL7JMaLCKkPe4T8ufb0KaqfW4
h6qxDmGdpct50x83H27WWmci6W3LO+vjgprsSWmrpm2/lEPjYTlANP5ESjILcw/K
4mpOapoN+ILVpXArvSFMrf9cba94sonH2l6eJ8KxrcfHz8xTr+7cXaYOAZZ9yV/5
fNA3fO7rt2qxOi8QI0r4+SpqDqcJwIsb345B2M9hwYUKQWCRzEo2YmXWppbZu/ua
ph4crWGsVzzLva88IQidWbzeDgA5XPltTm2EubT8maGF4Dn/jR4MM9SCPSggK6rg
1Hm6WU0s5uhk+ZnsM4RwOiLC7Jlr0E1cACTPNC3zLQB1noxK85som8PZ28bJhgze
AHfzZE8JO3pJLWGQcJKKXG7mmWO/2sF7JpSufikl5tB0jeje73ZgAhAyJw316A+q
FYkVhy5IFYAX3eyV9aIueneS1N3kpENtOUP16RphVvwMfXoPoTir5VouDv7tQDyV
03XctJC4qUCK6DP06gFLfwYKkximPpARIAQtgORpf6T4+f5Z1TTYlzx4YEd4JQfJ
EVTZKTkHdJrE9THH1hG0RlY/0BbMbd5D9aJvJpImAUVhZlz64bxin0+UGTVa3ddq
L1IVp37UssLGIflt+Xl/Ll088d0u/UjAgZyjzR9o4O2B62yV5LkQ72GfSl7qFl6D
Kto7qO60N4kLdRL3auAheaavmy8rE5JELjyirB8my/D49i0XzLguZAzOlGI46Dtp
IKh41kKg2i3Rv79IOvjH2lI2iudyp4lsuOD9dWPIr4dzNRWynHb+fY0ZOaiXydBQ
9FIaZ1KAGhXZLUdO5/3vf7K5s7rRYlkDOGr/GK8VkKOdVCgZyZ+TPDPc9dHJ0O0I
tPW4cfk3cC6Ob2CrjMwIMCePaNPXfvtHBdBSglRESu2W6strrVmCFyg656IOmMD5
v4HLhzGSstG9WBMxxdqPKqTiUyJ29Z/AT68vyGYCMTSy2xzszjqBFYlFAkg8xkL+
Lup5UnFAaX9JyLtDfwyt+nHGAdtSTJHmo1cec8ZE0eX33+NaF4469wkBKNvzBDoB
t9MeMbBi1i0F1ZauVwE5mQfaNcpNvAFKY1bQAdqOEQI6jsSkQFttrEnoKDvlDIFj
9gYhTfEwT/hLLbiLWavqwE9RnXB4n9baiIOU8Zwowx7qsQjNQhljtFwysYtn2Mgg
RWuD+IO9MWQ6OvLxvuuImdERw0dGpeR0SfAIMg5r0s/YvXdRZpj+NAn3McFf9v47
icpXGQ4EH3KI0r7XgIOM+7P8bAd0Is9A7Tun2MzEoSPawCKWSRcuCpdz78U3EWne
44xwfDo+lz+2hAhLRTPETm56RU5K1sOV74TOkuj8yS+EZDxcyXFeqfHguD8klZkj
uOMPdLvy3Jw4spfbMyPYw6RyS7HDKVQD7bF37rwUG7zV/8vP6EVtGuzPTiJyMFAd
QIAfR8uzXkbWdh/hdI0vC1x93zVHozOgmUDM68YKbFyyLqLXlESiFES8e+V7c593
2bjKuHdRTq7QA+3wzawPsOXqviKFogJrGr81jTqGeGddrojz12q5lDoKyt4L4oqR
inurTnFacfdFd+GY1hHHbup8kyRk79UUYWsUymu+denA6g1Ssf57pWTqck9A3EUQ
xz2g6wQtEG7+TUxnNFhkejhE7Dzvldh8TktxfweVSNCV8DHgTamVOOiXjnKp+V5m
tnU5AoJqeaUm2THMS+ngySeeO2+nkM9DQngNoDU/iyod4UhWdoKmEPjUW+LMXZ86
qTGQypnD6vO9Oq0yPlf062HZXugWn1Bjm7oudKDYscFFftoQ3uKcFh9nxKbMLPOB
tPWHDSEHa2QxO3QuBfw8OdGMpeTqyfwMshaal+Dqjvw1CD+mNzyyqEA4Q9NiP5DF
IH5lY0yPYDbMpjDDkvhBFIQYwlr4TNri73bQ4FjMiEAZSK1l/VWoxLWEMbrGpU1v
XlzRliiH8sPrywWS76YAuEgxku8v7iWl4K5+11y8xR4Utq8mSFPYwleeGu3QTUkZ
N8xOahbUIKKdDdYfDxt2yfH2NIvXN5hikJDuRPt/23X8ut4WkwG6gSAuiqpFQwga
8IlsiqguglsAw1O57jWwYD/VBwJkLu1MA1B6vUgP9x6c6RqYbqld9QjJvW/K32+e
DYWi4fOXdh3geYiekMyq0WdEw7eLK//KOuWZKltRWmkG0Yh90GVlkxi3pZMJZCx4
JEJWDqVcdjd6RTlZl3koVc48S0uwR4UMVnX7A4CkzUU2c/S91+gK3T0OTUNsch5F
S0gJ4EI8eCPowCdlvID28WkQWwm2FzeQ0O/BWN1sWFhMPv92voAv/nS28tOSggjn
C1xVem9o9rxXY9XJ5y2mVZtMvRNq47DRujTdvNiAoHQfpXbzyYv7rNifNJGc32we
XMtR+TxU8pyT5musRn4o5VV2/DHM5ml84hQc7svcwBI4QfCPkkDTYx8u8AV0TMjT
Mg7eoDqVyjrwd/88uruWNkLkzuPxhmTj9xg0YRfl/hgZXSTgy+qg4PqHMcduToDU
Id8pJ6bIn5UKzZxVfWKZIqFx+qUnUPf97Q4CuAHLazcZT4HVbCKHtphwj49xKMlN
8/vHt39Bv+m4fVSKBVoSuuBYbCuG/NkA9/Svh1zMCjRxnAj9jAyy2ZMf/y+VcyU9
EXNugYx2Gk2Px/+KreCW+27Bc5E0MA0pS8l2v4Oae/Tr9a6zknNccK/rHEnhZQIL
V+1utNdiI5chjjGnPSU+OJ1NIECe4y7Te/ijr5EWyYKQtsQHIDsJvFRhLWGeOzwp
1ndA2REAh9i1X/Hf5Q+NwbiuEh1kXuI33+cN8dJsMXPMG//2wgrT/3Xaqx+uxAVU
YGXSdsCfeN1AHhhfgHVI3OSJPvtPISMKh5Z7z6icGoYiPGTBlbXGGYOOW07RRIyV
MLptTYPz+qj3FKjuQHEDuynvfwRel5b2Dyy6uszwO0yncYDG1iedPLdF6NTV7SvQ
g15epozocexOpFwJPljhPDpqGYXHLurhrvAWH459jKxidEeYI7u7qvtLN5jK9OOf
gb/gj6VN/WFw3LbYzbO9ByAci50eBuZ+K3u64nuUV2BPjjE0D2GwnUNPYumnZULQ
TWWLwx5/ZBXoK02mwV7LsMzYHIZGIVKiEmI7++vEKf3KfwO6eJazycX4GyS4+b/2
BhCul18p4fhyjHatKERYW55UOMMs1+pTpFMQ2FBiljgfMipi3eh7d+GZpiZUFACA
DID/e8t4DfmQUX9V3X11WNx4o02UT0s47sNb7Z5zZAwrWPiaupLH4hsV3dgk2tXo
FT1Jkx+XAOkrAzdgwbxT8LL1eXlPYNJ+VTkcMdYs6zK8FmGQwKkT/i6fRmUktfva
C44OuLjYm2qAKNVV35U0vgtYZNFb0gIddcCuZglTf/MeHRiCm4eNCZ3nUM9s4l7p
K7zDXl+9Z4+tbTzLkYzhDIHx27nrvW6lV30eGA7hpf8kjuwiWyHPSBcleNHWVZTR
wqvzHc51zlrhpeqFGUnR2G9nyGjLhFONAmlzCw6kwTyPzUBMLMh3Z15seRcANO48
H2EiYn09F8anJSjoA4O07QjKFqPDmIuNdYWCvixCDxuMn6jV2ozNc51/IdEezXeY
JqyHVSvqk2TJy7+yc0dhPC0U8xp1YHfjL3GMWghp4SokL+b25bGJIOR7hV3zL8nR
DNmOlzl77ZYaP8yUu1s50BXV+AR0DX/fCx/nPomxfJzwwsnotezu4YqbCWqcVztD
G9rgeU6GgG4IkB8wpBzfIiDpf9y0oHEl8LfqzmBfDGx5o/2fajfrSV719CCTtwfA
l26O4Kxed/Agmb05lqCqducxkZclBMqY7tpWOrRlNAvTYH8cev27uXlOL+lQbNEJ
9Hv75fJLPkI8ePcl64XgvpJBu80cEmB4ep5nt5K7loX4t8jESkDAbbjfg0ggWiJH
/Iy+4IvrIITpBzlWYNEvpyG+HJx2ruFU7324alMJhGgUgH4tmw+JqGhLcC1pFfqK
2FGJxVVWCQunS0nl87z+UtmqRr5uLxCwqPU5lXv3qz9+e/I7/6lHbD9nJlCvUUY3
AegSKUvZDX75HSJu3jvNFstzrC26c0KMshPUw8AwCXLP/H9ndEEFfIfDf1c0co+3
rTHkRHnDhoHMLfobh+eW67j8/NY0fAoL+kAZDnrzc8Om5DPoz9Y1dPhgAva1kdQK
/QGtXLMgjynC82919qZCiRp9IOlaikT4YsNdM94cMfT3eaBBcVOB/MmgQtNNqXOW
Y45aD+w6dSIMW6cPKTvz5is88x8GN42flAAsLMmVIf98m2vmUGVVYP37bxXdnIYx
T+lE3t9gfIZ0BxChf65ca8zJzxku/FlNGx+65vGfDe1NMDSLPE5x7AXBsaxyfx34
Gnx+7W8KM5ek3lNN43e12/MY3Fkspk8tulIKNvV+flpEzfdI0yvXSbk1/OEELkK1
ZOaw+3zcUiwTKXE0U3COQrBuxFKbNEvlePm02kYyHM+WDWlRrUDy4qeaxwR5tfB6
PKky+H83UQ8yL/mIWxwK+HNRGN/WE+HYAdgCk/UceyGAIsbuXGJ45D+U8b0dDM4F
5CzeWFJMCEVUMgBqc7JpHIj0VRoB1MU2mQ54SjDWb66aXAORauSb4dGN4IA1YWvS
DQ7gEf5iugv8T0tH9qYNbJ32S2JTMoiAPn51gWgmXWLZF/M7p1l4DB0f+IGv02a6
XNvixcLtizjmznftG5KI5g9pg4Q/NXqf4IpuodrNmuRt3OjXcK1GFIpSVXLlzCWX
UgrCvn6Cj2oRy7y7SNgxH/JlbI4PiQOZOYOvxoa/FN8WGIjbrKJw0RLwXouYYLcP
fOMOfWvIptHJ1ohy73fEWNUC5iVAeUq1e5co+kfl8ifXiRHwdFk8Ljfw2/r/be3F
diVxY25Bi3PV0pwQJa4L8Q8sgJ4gUcLoCR+sxoCKS/wvMsBqlz0bwCy6cImkWvbW
n7tXRWmlqtcggRZdV2eaDYEpLNvTp3WP3nJ55rkqKSogfNw9ZmyIh2EvXSrnwa0A
ZPbkcMQKsCv3Xz2uzpN/JK5b4Bf9H+aLiBr6/ICKdCj0MfY+6Ctx4lEFEiTMXo7y
xQ0jHLYa6CneCokRhUiXnFYFqzQUz3ZwekTHut5TceC9oXdbPFbghqPcx+P21Kiv
DZl1UXh0l/C1LDaVwpJbgc4k32Tw8Dm73kH8htKI02dp6FSKrghTc6BD5JUX1iqz
aHSEQZDhWiOMcYJfkFNHxfPwGz6Px4R15CD1/KIxsVQc/myv7MXzKECLoR6cgArE
KP6+ZbtsOXw4/6qTWmuehHa/0XEwnpOvFcYSqYcKoCUvHwrlmlxv1ra8zEwQvS/k
q+rNlD0uTzyxYdh1IdpZ+jN/c1Mz6UdZdrMQJpmsO2kW/RaWr3Rm4NL7LGPuZAfu
pbsHk9b+8ebTDIEy7DVgyKsBkn4rFE/eKkb3biRCVeX63S03bdhXNQCxbRWstfE9
8Bw7dmV1R3TBIiUDKDWPXHWjFX5KT8Dh6sq7oJy2mFRAS46wDfchHgBH1MRpw3PN
NiITuzjp3Q3VauJe4XDs7VZCGwFaU95ryWX2UOViCEs7GgG0pG4tUc5wrfJ+zI3o
XB7UtrqUbEqD0+plLWcRRquaFGzSqHo/IMzNdjAElwPt7GBSx5TDJynZjAJtBPaK
C3UK6JmeMvpH0JAY6QquuAPfXoh8PYs4Fvs10HSi92rN5MvLcNulFlaicNzyS2wJ
gvEvG8/c9t7QxZTB2iBX2hxr5kmjuxPi8xgmYPPquw0u4gR+oOUD9y0+7mcJmF5X
XBHM2gfIJCcIM5TDnyqxYSnRgU0H9xhTC+TGQzYJhjX1HnQB5zqrqfsWndZ9lPE+
OHYO7oleIQXqEOO7rFuhQEMxUn63fbbiXREZbUowhGE7f1eef2vyEi23xTSN3qq0
OhmWPVFnEGgHHNgIJGxtLQ5h0lQBCtYA5sq1/JiYgd/r5vuefXIFVteu3dd8BlXa
Fwu21Na2T+Bdp/xS/jwMYXgQi0rD6u/hEIDG5GOFK1jj422h5DMA4NbLcrr4namA
K/8dQ1lnwNaBIbTWsDCPa0+3EUFRZrgjEASgMhZ8kUqHMvFlxC73obHkGixcUaka
DfG01PvsVBsWGvcNTnOPweqEzY92NqiWCyiNwlHBA4Gs646iL4mI77OxRgXAaqLW
M77QPS5kkl4hxBHwx7Lh95sYbKSKOVT4Z9bOcnkmx8/+8MSY7+eJdP83+Mc31iWq
bN9RpHdJKoted9aCfTw+xmvRS7mgIHVLeUf+PWaHjD0d7mgChS0oFOkNqUTvXUnt
2eJfy3ku9mjtcVsW5MnLbeu1c8xkzYoWr7uS7UVR3A+JWU4mteIeATly4HK9URZf
hftUrfJObcRTzXV7seN/9QRNQGGBHFXnYVFAOIMXhEMbBgLJyvQZbFKLndCuwpUZ
3MntOvEBuFTBvN5sBM0Y/vJBAFPZtv2yXmnVwP4dGBAfkrbv6t7yC6p5SV4eD5Hb
9N2+SE443w/2L6bdPE0zhnhly/ddEBWlWcasPStm2tTutv2cDkjWCFjnmG/KOPRY
7YeM9J7sXwg+aRjCbryHjUUBc/yxM76lDbBPPd5tlSMEKM5Z8zXQoaZr0Cnmcpk6
+IaaL0idvGLFK/xwX9+DHk3P3xUj4vmdvllSGKU1LmKXyXyy/QsRcSzUMWxLhdHp
798F8rf9pLcLs9w+nWBbe47a/vU6/ltSSYklspouHep7SAv7yEKqSE1+qfyzUnbm
W0Sv3shUJD6hCC4E7kym4ROOqmqCAl4ApHiKpAVgNONJOtnqZ9WW1l5ujliU8RZ2
MBKU3OiVECHeo9rcbqmCd76puvkT2YZBpEs+1OEkWK0w9J9+hVq7qhg9zLnktXA9
89aLNQOqiISOVQ7br6iXvCdxqW+sjfNyVytRYK4cYFtUZULiibnbapx9ewc04cLI
zYhG23RnXcTSAZH7hQQ/NR+qRydrHpDIGNW8LtWqKTnd/3Xko/BvyliJ9+xa7da/
DumhBy5GWeC0LlDiXuKZ6Gdi+9gAOCSD5bL4+DxyATRWKNVA3jf3Mzc7Pv058TDt
f2qq7ODPaS6KH+UhbJaGQm8ZoDeQLn5ycdXgKCNTxOWQNd3ziDU3EsieB6LqCYla
OA9rj9Yl2y9SJeZQnDjtczrFMIfK+kuTnDeGWgaeum2ctmH8+YOgghS+Oug4P7Hr
eQEnSZ2qFKk7/w6AREJiqoND1XV9MAnMyJiSUqCLGDECVJSx4dm1nbAy0/f6VmrI
viu8ZwtsAzQYEIR4FgzQ20M7aQ1++2T1ZNcO0mFaDPpVD/JqXhKSoXc8PEpRZZYC
ZVonMCXgWeKmHXLd2HhEgXKtbzzYJINVm0it8ZIsZPonSYLCsnbZA9q1kHiWTR8u
pGcK/3QwFwCpaohQ8lTNVj3MbBJ/FYQcLg5/1cWFah7247qQBbu5XLcuroG96rB2
ABkH0JC048SycMepefuOLZk1Xt4vBwxy3SBFwq7BxYw3Ytq5B1aaHxp5hpZhV4oO
enNkUc4ngMBeLBVha06RfiejpFOdgg1AC2Vxlt7wztCN4GhkYYrmkndlKUY1UilC
wkgBDKdlWX+McV2c+lKiSoH66lN7tEYDvlQGmzNAtFVMW3nc2sTTgsoNjo4HJL2m
pqefiDtCnGRx3Rmc9MMuU+izgY8SFXDiH+9LV+Sk4/CkU67qQaPdINgZqrCYmN6U
oy51c3AtzQH1r6lU60eSA1B4ZhnhjR/LawPBk34ocbAmJIR8aASQTiMUNqh1u02a
UGhcJR4C1LiFjyu/iZtJwqBBgx2zFLJdXCdjwebMS8e+lp4P4qaK2BrqfvELNG8B
S4r/kfl0eHQ8Su8sqE4d+vAfIgV9rzbRjPx2vs1HzY4U0/vsl/nF9GMyijpeRmof
ms8n05bWyQOz9QPi/73zoP8savYIATrEi/cmQTy3+E7RQXYPmi7Q6IAPy2sPtecf
SpTwD89AIbNdvDkdVHDhLze38FAC0vyhaNW2fEgeZptY7EOVJdrbZ3RqJ98kSu5v
YrMv3lujdtb/c/x41PIWTfO6y/B1hhexEaZFMUog81EapsBpbHHZ6SXrMZZQqXU9
paD1Yi1RrS9gGAHDS6W11xI4jgtHcwMgGC0nWEaGGpCzIw90dm/urF/njUvcx6rG
FowST6m718dTbGa+ufL17ErzrE1XY2KVJ/IMOZs1+4vc2zKjxqp3327w+MgG9HvK
MxGfE+BSOfaNTkWR04ee7xd/dyDt31+JxhwzzJKwP9RtbB8nD0XynX0ZJ1EgCrnH
KmICFdknFdGjyhN03B2K9w2v28Dsg58HzThJ2SlTRPElbT0SMZe1BKbVZ0KMMybm
WQBe5EXcSGNuZ0kemDMi3WK67YdlKBIpEK/4yHoPxiVAxfcabVDkj3K7bZFmmLn6
o1BLzv92X8Hcgt+U8toWgkWNwm6eowbmFnQZtckZ8iXsG/JUXxnpIo+wXn3qVxb1
6T8JigFkQWr4XyXBRnmCkEwFSSiutHMI8plESnuDdttC/CzP7D66zB5Wr6dZKMi+
GpnYMDJz6SUik5ByIPdqAbmxTBpaSz1hga9+9MN0j2+wRCXMy80qbL/qmFnvAT1W
k05ZqS3h5MK8bJZ6Z6nrjtGjAFJ7EsykSJLeBfms24en9qG26oFiLxSyrtkdk7p0
hVke7uMwf5LqaFb4157voCadpFmPEZmlSDtQ+QFOJTCpLJRI7ZITJmHm8uHed7DI
0h5ThKuM222D8JDK8tyqSBL1fWDwfTqf9SGpyArUxUJbvWRuh9pnSG0avW68GEbv
6QELLCVYUEz/LrJoLrkMTKh2wFa0i+yyemvAXnMLbX6zVMLU+SpOh2zvHTOizTnr
vQz0VifChXQHVUs1Jp9c4Jti6zlD7rIuyWp8y+qxHDDtopa8K9lVrT5lnHUZSftW
VnR9bufAhbTLUJMVchetUR1WEBiqLekzeTYdSKCCPQjj6zzG0h0s0Am0INq5MH1a
zFNfKNSex1QOMOSL42+L6L3iHwp9ERN7hntrLi4/2eAJtKij/DnVLZ/gBYlYyIdL
7j/n2g1TKfodKP1DT1CE4Zizecury37t3xUdY4gMlQuKJTPeB+SISK5Yci69obY+
DVDc+LR6LEOQIktMBW/5x7PWWUFNYUTdkLijLYnHsUrSMJHJiHn4Qk729/7J5kCu
Ax+myhiLGUImbZpngLQFxpIkLxKydKz90yvBfkIgQowwY/4PJ2f7ywlkZfSCKR3p
Moz4oZYmVYLVSO4XrfnkPkP21/P4MiAkkDMPDl7R0JPP/Y+rlllFNQQdMgFcO3Wp
/S+COsv4Od3XWAfpBcgkcPBi7CCduQ+xFSzDNsoS9aj3OMHfguobxIh6xh9LkwNh
9HZ4gT6IOA/FCyMRunaOYL9N7ph8JGbaldLfODYwQZzWIJbyv0cbXESs5b16YNeb
0Qp9BHesuEk/3GyTSeLyAifW1L7JRoPG32E7X7UdiTJShi1CMC8NlibKlfddqtqQ
1OpiI4tZHupmdAA3T2ph2VAbuJbQyPBxJ+Slng7z3MMb1uXfe/egbc77sfTdE8db
rjZ9pfNTaJc70o8NFlkZOcZYRTXDLe2uW71syZXuvZprGYhBcHuJfzEFIPybdxp/
IXtbqqrPONve2HBzrsZb+7fcejf0oFMrv+zzhVVM6MhZSpKVAfLeHZYBzfY6JRoW
KCEewlu7x+X0r3PLUGGp3vV0nzoyTo/ctqoHtP8GskaPfuTgcetfli/rWudoerlf
jxkpx+SyJAKf4bl2/mJeOnTkK0gjFYG2IZjBL3ppEEWXKsgZiP1Q832u4Ko58cZi
Mj1LIxltdylg1P5/3jSMqZVBUu6fiVUQdHi/Jf0+W4vVkHxth60URPbr3Di1ySSu
S+QaFW/jcgeTEjj/oEdCFhYAItzgYNnmdrvo93gziKcWWSqqSMG6maZcdTU7X0Kj
Q2u/Gtb0xANxhW/Zp3ogSy0p4Ui/geGoZjMzsg8mhauY6M9AhUDvatOUCK4bMQal
7QOzofvsvQJ9iXfVlHWgUxMqHeYDW36YcMHy5L0mAJMtpmmhGOTbeYcTn02KeMyV
puYS8bEkyWbm4EzFrpgSPh7QEtjOF2cF6O7Mi9fDgJLO1ZkkS7Pk2XYFr4U5Dr1Q
pwy2u09fStO+qvq9B9sAyYjrTpiEDKNDXRG0GVsz+xdPMH7AvRJcZAbAKxDt30wQ
bRNFalTPxaSDvRgi/cCnKxYUw3adBQuRruTTW7ze9Peu6xfrq03ozoagWwJ8mLqM
V6vZlb2DTfpuIAepGSi/XIu90ba67AAcu7TOMUFmcZM0gsqCTXoP8aSUBhAjhcrr
s6WuNb0e6/z07fEIOM3iqABfZRxAdkyjs60ARmeLih7wE2c7Y1Gy6iEgi5kPeh0R
tY8Rabnwx6Wi0IjI5kGF/jnjxWHCLwxTnGw+3BGB1nB6iCweFoXYL/1/DwsC5wXr
Llq74sIjzAzpMvZT7HyU+29iIpIbhDlN4D3UCKQL3RsrcuvRkDbMzUfj3g5/rSt+
DQfNJBKNAYWtFL6M8E8BIuUInyOfgpXiAC2ErAmmkgbFbnonYTagibWKR4HFQWQA
aQem/nLXKx15zxbVhcO+VURropy1LsK+H+rJhMRym7GaBNeHMzd8TrQw0k1+q8wk
0YaD1lJA40v/omNZcKfUWPMT1gf5YwCZWDXsSBrOCi72fuO8x0mJ3gaCYr1mWZQk
XSUb+xNYsHJQ6i7T1pIwgWXz8sWEOke0yOQfSYNeZ7EeSKs+3EXh20hM+8d47LCM
4CKCAW+SM0omQ8Fs8+b5jM2ILF7g7JEPEHMnMW3ZTH+JH48lmKCYakBk+/EkkM5G
WXhyS6yZWqcsmuUqbG77ULBz8WWk8S7F2vwfyKF+kB6sEGn+gf0+DClwyZ3aCG2H
xnDDTnd59LtZzmtKe1aGjcHJNf/d5Nocv7eQYiEVv5LY7U7iOnj2GMJO6HXGELXh
JLxrNRmEZHR5wBLVjM3L4Ao+DNpafTyKjz/68Kd7erGjX418NCRAkzdE3stbxtBV
UkFpJXpoXi1ONxSIZMnTVPfArbl8gnmr1Qvnd6qm/s8xREG9OcaIa/4PTgCbpdNc
w4/Jhws7V7Lvnodcgb3q98qtpSmPAi2wZJZxLKhsZfDl3zRD1o9fIoB0o89jL7My
18dAVXs4oNJF3qLETfMf5/B7W0JlKhrH2IUfnLv9A77LzvWFcVUt2sNNIPyXnSO4
`pragma protect end_protected
