// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:31:33 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
ClA/IX7LFjTqGtl7Tg9LHOpCFCFmJYLV+VWRuRD2Dook0PedD/qMmeRK71RCfGpR
QqECzinEkQAtvLu5ZG09/ZkY4rRG9cUYysno2oWieUYuipupDDAv/LEtCHJdrI9q
0Mp2nEg0EQ0QfhEAKnoivAYKvDC0RkNNYiuoTfl+JN0=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 11792)
1wekg6qtn3cSzMjoRS1zzoPoJ6OmP9SWX2K496xYN7flgeokJYOiVExRwn9xKaR2
H8poNbzLMxZNecVOpWA/h5+MZXSJi7RrabToEUhpHHNmwdnD0umkRQ3Z++UZumm7
r7LaBsqL5sujMabCoJ12aUVGnIvHsnjHolM7XjYDF0xYiKGw3PO1yQF+wjAH7AE9
axfSTkNm5BIU7jxr9MVmcEx9iw23lADDHXRRF07OhRSR6dse7OfTTlVBAbgoQoQt
vKg+8OZJYDT0Fhc8DEsoX9cT61LLjI7OoO434RolHR0sHD5+AnkY4UzoS0tacDwU
t6YRnjGCdy4LXm48ruK76bSVe6rVt8Gg1NBiRbEDYiz12O9y5fnJ8rW9eBZK7l74
uUBDr1GC20dZUXGJQP9EfQo8ftXRClLCNciBwF+XhlhsCx/W6nTwvjqgs07vvVJ+
pQQFKdoME764tP9QKtnTklJf5ayZ+LaVxzAlDAZmB6GmZF4+HWP+Gwi/sjdJGgR/
DMKY8uiJ+gFQOeCkOZ3bH4+UU3nEXJy+qR0QVHX0dWtPUlOjPcgJZqY2I64rCkur
EKBLLK/b0OE5viRIn8q59vfsQKT93ynIZ9MKHLciQ7df7FxHyPUWD6xHk44Bzz2n
xB1s7vXuLbHgynSshkm9xkybxIYB5GBHIhvdw545sgqO7hMyX5Rzsot98sOC3sR/
5X9KyddbZGCYfUEfuEyfDmAQ8+xV5UeaBRHv2GueOoPgZEM95k/tkz/vjgPDLckq
8xS6a93ge/0cEvWPD2CrT/gZHcdWUNx8ozIu3C+P6syVdIEXSzqogt488O4njvEk
nfTs8bJhSx5UFp0GoctxCVj20MUOgjizapWqaPr8cZlEgMfdOkd0aVaTXFD/hg7a
wMd1FBjWEXJBSseFYQXt7tvarPVZ/hck/R5XkeDukOeJBc1apdSZrxn85dnEB2kL
0eW9O2HBarGOZEZ0LaexC1VE5XPvffDi4gFZ/trjDRB5tdY6eLYj5toWhHHggyR7
T0uN6o+sLJK1WD0HWpl2917bg9gWQGuAoASG3g/6kdTwSZv4ni8pbMjsfY9q9TTh
/H9jAjdHbbAPcSWl6pA49ISedsgElIj188BShT9xJ4EeetBecfOhhLeDgVj75PQ1
C/hqx+ShaXsNxKYonru/ZnUkVWGF0d9GS2dY0pBKvJtrR4uVwQiDX3i7A52UMcxH
o8c4d7W0BR5IQKfhY7idGq33IH38anypkLlKjgYkDeM8raBuehbNP/E8FApCzL6u
2zbLYxnrMLESQBg1qC7UthRjq9SR6+7XbJRGeLE5OZRu4wyT0EicUuR9G8F+7ZZ/
+Kz8/4HanvFs07xyHyqrCqMFSrIT7cuOeTa41lpK1Sma4SFi1Qsjkcs9FSx6I7Rk
sX+yfL5kYo3VNweVDdwCmxZX6t2S4FchTUIrEhZRxTHaThjKZuet/ReKOD5cfmy1
B6M7PCW3GWrRHjIXhzbjVUy0HIodjcH1BvwdHGz6ivuJaGdn2QMaNsgFP0EBjT22
6xPjjekRs88yodPGTvhEoXfkiTgUGVpNQEW77NSG0ZoL9V8u3dSybFS2kn13U9kQ
QKx/z3pdlLKSmCIhwhwWk8WYxXW+s2LJome5VZKeC4GiQn3NjTuuBheZSv119L+j
FOMoar/neHME1sE84oO/aRKNsQ9HGEpsa7BoCL3stO3BPHGbegm6S9H7UaOU5sWj
bi1N6/qAUWyVxiiGTqMUHqbE1O9/BWx9QVW5MjKWhlu1BMRDFd2eFawbG7Y5YV2e
LlMLiRoBd/Ao7HQyAAjOCS7VhTeyTmmNcxREe+W1nRVLK7SxkFnswCzNyvEjpR1X
ysMoxjhPgbGUziuPEu076T1djdWFG7D+DoYUiPT1uI8Tmmwfh0n5nFE4/V5CHJd8
jDq65iVA7r17WNKNqmdmfLh1NhrbLQRG8fgN/ji2PeBFQ9jq7IYb9tpYMqf2RKtk
xH2VySBo0jpTuOLgaGqXaiMqJYZoav+thvtFX1q+kVpu0x+d4dMokVMJgQtWQs9u
phLDw/uVpDDPCBWu5ZW7ey2IDuWeQsZPLKS8kvBlf7wQ7jGNTXnRvEtvwJf4+3v0
ZDnSqQ4Gf4f0WpvNFvxll7neXzmzJdxTh9i4xIfX5UK1fdSCjXA8EIilxODl6X4N
nFx4qqTHaJ7x28EemUat+onpkJsKI7yjx9BDohzEPq1X02gIM42U4pRLey21nVgw
7FA6PfU28ZbOsAQ0WaLEQVftxuFjr69tO+CX7AQE5ZR79PQsb/9FENIuFKhliI2A
o1vlNu6JsgEVx1bDtsmke+rFqpfr0NSmHtA+1tqAIK+bRbJ9T2xW2kXYn1PqKFVD
/gKDbPIwXI8MrEmqoJJXqYB9Q285X+iFnM2uZ1JQxOQm17rxtQpOPvqD+2T42BPB
9EtUB+RGkQTUcWhD6K+VoyDrnhEGQgFr6jpzxt57PzcW14oqSO1t3yWvYZZ7bXHc
OifRyiWp64g4NAK2yTfMmUVvDK0GfySMrMd2uMij/6D0lrvLg/vOa7s2OfSP6EqD
mQBoxg91GrycLHyudhsh8Z9Tv2bce8U8p7KRkqdwoQBzxYdfVz8CRHltHvakufdw
eYR3jLjaC5bYW1gqGI3k0iZjErfsijmN1z4rR8bB1tHrKy3bmFA9rxB2um6F+2Xc
NnlwXYopoMFl1tlIl5BkQxNFioIIgMjHQncf/48vUA3gowf45kW9QPJJneE1ODrx
BLVw886xzWhPb2gmxopB9ITRivkdKenkk0fh0OOVeBqPAJ0RLueRCCGkR2Wh6zfJ
qfKv1UTwdDinp/vlnDPeqWt3XD5nqpT1JzSq1rTo4VyddjApU1NskIIIt9foPVjy
2NVuup83VPgymoFLnvTbAK+YOiViIVQoGgbLHM+KJAYontcsd+OkWjFM6xO1iKrd
4IyIuTwRE5lFXoCZds3HuGkehBj8jsFr0j1O2aThqondZ6QR/giL9U39ZbJvVc9K
vvlwcoVEiKn1hbxnP4KuW05gcz8GOY+6gxU7kXSRDinqwCYfBqEp/LWgGLgN47tl
ORppvEl5BpARh/cAeCYaY27+JDAWPUh76HOAg6IYjTbwzdhZDCMq72RMQ0+zAKvp
+zrvRIi9ioHHS7J9a0OKdY3FdbMUUmC/Ji+wbxG4POgQHWQnuRcJJF00XGvFYz2L
zvbBupeC6BAJCyASXH6zUypbJmwiupN8yIzOXl3ij12AaCeZc47Lkdb8+4uFqFUy
85T83DTkpJbi6a5UvnmUkMolc0xErKgKd0DTny05wKYctwBqpo9C37SdZu0JS968
HkoUnNiD8gXCV024x8a0XStOzTjdEe5kmWlrNwDAJRTbpiC6WYzD0CbMy/A2ZE4+
vwpfPfgHw7Xy7CZdSSwDnL0fOrddzSRpH1Y+E4KOkzceqFvIk5EJ+IJI+mpTlhfn
EkEbRiiqfSu5GB9A6aX1b1RwKEs68dHNn4hlhxRgTdKlUQskC5tPhB+0Ufv/xi+b
e2olHWoUIe1UaE0Q5wHpq14d9XMux8DEYCDdq4xfa2Jeavw7PDhj/OObXRuj4+vS
QxSItRFEQI3bSdCvyBVKqEb04jcG5ab2RQ11Tw0ceWSH+rGGI1KKXDGTfRpZqeQq
p2ojk9GgBo6Q1e/eAWlMiBlYAzUOY5mKOAGHvPXJ76ilnivOGu47p8gt6E5HpSlT
ZklTfWhZOyQOqZwT/WmybT+PNct0YaEgpCL530qVm91HYTpCsdwSqcf1EyNqSixG
2Cf+Ao/Oyb6gIJ7C6CJyGQKuGwcEXJpr/1oKUQTDK/qoAXUj7JTGUW/85vcLVmjm
7d1v8TYDd26sz+zHhs8xDRWo//4Xw+TQjb7W1SJuFe1zmQ8Tuj+5CSfpDWQ1vX/B
xmP7BbPKORxsrQojYku6MtJ1urTBxDB9UPEOtCJZwbup6nYcszkg5ApwBE7cAmPy
DPWRuvr9Tol8QwgOtzfK/NfXEMtc8e3BqCLrCvFftm0nyA58QfzPmFXIzx+BIHhk
XDafPaAhdqSXUJo5s0TLlEUzv3QCxuDfPoqqwNrrRtlWv/FbJJa3Z4HGxtU4SpHk
2O6P3LkJCcaruRrU3/aJ9UnneM7VLk5JD2kaqjGRCP+vZ1o4zkaN1YEKdFZhC+bv
G79vLuNK4UhUQCr6zVYDBfrz46nN/ZGkHCknJuzANn3eHCawwohhGm/EzEGfRUqY
LKMticyq4fAJ+eK0z9Occyue9JCIzsQIuiJ+HuwhsmMTm2ZfU66FIY6/tIfIBN39
v8E0EX/a/W6tUv2U0wPCv9vWz9mfS2UQgbVXP2Y7M9wpBPmrgeUAROzvl/DckKe4
9Z0YrW/VOiGBWYGMEz9ZsOk76vtXULPmZbGv267+10cEUGii543RdkZ1rw0x5U1d
ZM3WGIHYbyaZAla6Rnu0v+CU9fvdDh/JiLT9PR8nJdTQsRJmFYO2RsbbSHo3PYbW
bGoYRkoGoO6D3p6ntheJOo1Q1q0uBOAtGchC8yo5YB6b/GzfoXmkUpe4+U3NBCL4
lDuOk9PKBUNoKUVGu98lbEqQtSnG4gvrVHTAW+zJr0C/Uts3bCzDfJwWPKKer+JE
P24JhCVCNmI4aIivHPzqqza7D0tmXkRPQhFlhEoFMTbBGHNBhtXqFQGIIrAkdaUD
DE+XR0yH64FTd3j6HoU1TEm8UT97pDqSeANyc2qbsPat55zjb1ifSAnuCbKq9UOs
EigQp3nda9fZPvd2hSLwApRzLs0Fkkv4/s8V+SaD/Ij2PCVi1nSKN7SYFrxpcKLP
iauQM80ud9ILNeJ5Pm/6hrG90+K2Hy3EG0FKAL1ofV855cAhMgjsZD9JMWmO4NKg
p01VkdPG6g+HoMgetanPcqQsfYYMR0jxpk9NoVHZ8gbvCpMvvcjNPi58KYhCvXPI
W9FCUg3iuBYIeDYSSQCMyOImdCZVlb4xqZ2WpPPptui4WKTUMu9f7IbZ6pkJv+K6
29zr9p8t3aoAp9+908NLwP+jFIRzYfm6awGtdPpwAbpgRT4KzZKVjcx1Hy4YIYlr
z5KnY5cIHIa67dnLfJ6aZW00ebhrICtVpNiyLxH7KjowFCe+g4in4fPjyHEhl934
N9ECAi/YlVXQaw0GHFOvhocqlfNZo1V6hLsKBtFIpyf39jkYR8bEmycLaKL8xujy
ar8CbhJPdrs4zHeSJwfOr+xeQky+v8+e4SsTz2QbbVe5wVuiqg2H5o0zN3Vo9c/E
3eDamobeJRUh9cL7KPEYytLxL46F3GxlxRgJKx2AP8sAyXwhxdKPQdVYvhkWGE4t
UvVUTG4FbMTCZo1+IS6LUriRGk9rHp/Ivxjz9eweufM9LUi1Lg1innLs2CQScuNr
DX6bJ4NniL/LyeB5tdEgKjEPPmVsVqEPHj6j9qeSNuXqlDCDX0VmHbcBCfZIIWQa
htRiYUTZ0PWw+7LZ3FWY42KNPghLZsfoLN/CiX8zc/PpDohHySd9dOxQiA2TGZ4e
AHfVkvWfhqeemEbbiMWz8/ejj2FSAaacXxmPEEzrOqj1vPHCx7o/eUtyLNdlsnAc
u4+qDJF0caNsKmgcF9GkiVL+9vK4IaJ25uSjiP2tuenA7yrjpf5hQRTi9u+OKxSt
s7ojiLg0YeqcoBfiB6EGyKYwEELfIW5yhAaTeAHaJdk2chxHTuKYiOa48+rXgppS
gsxkWanVFlulSNlnD8uaa3VRPDv3q7tAKlvxkKjvF+dzc24yrYSU6KZ/xWxk9A5X
OhN5qUUlLx+r5Apo6VVCIsMkDUoGXgf38HRlT8hW/uQYpAtVSOg95AAHnBehC9qy
zH6a7jTC+XHS8Q4cxvrVHxNupc4kecYxVlY/U7vzbV5b3RxL2Awz048CdyYEavfR
bAn/Dg6EAEmnRLsJvQUw2jbOJQfT8nN901P+/exhw1aujno12EPfFirI9igpumDm
bj6A2rIRynzgAfnq1AeX7VmndmJQ8pQKeebDcIF6qT4xTyqr2637zd3WBD7qYcQR
xGKr5VHS+rYIS4IUv8tvs9p7EH2Bguv+kzCD4uyjC5Xchqb/sK+P4z4QhkAsbzNe
gzo0tnH59XeSZmkfOZc7Sw50LtJORDDvighqHHv3eQTqjz0zyVfiNGG2uskyWr5S
fUuhM6PnQpX53Atw3+Tgqi5NxCIAXhj9h1S0DHgDc9+4zeBl3NqG//vsPkUAM9ni
lBVNvRT5bNlC1LPYMOR5rWyGCwm0WbfR/m2DXrbZvYWHgYx8VsNenVkXbfdSqXb6
oh2NaARynJxKm55AUryHa3i7I6gBN4PLx8NLBI5Xl4+irQfIZokLpfI4abKQ4eOQ
5A3x3l3QQZZu8ibvPxMTZpiiF+pg3wyaX/rPCKCnXzSe7HYsK0flRO8Sxjzz5N9B
LNtmnfMcdM7YsDAslwDpBpZC80nDD5yXWRQRufjVdbcaZKeAh5KopJUEPyXQVF7m
qJ8ZHMhtieaf4Esi/PVa9tATpp9h6e23lO02BPi8vThblyPI7kdi7V5/VhVwWitW
fLCfKRoAymjRd2Vu4Xa8Zj7BdP69WcUBLt4KvCXCiN/VXjev5KKrNeth5SpoVbuk
JPkWZJpweKS5Adv4M9gfs9jVWpZOpnC+nWmd8Wlh6wCg2RB/EjxBFctJ2X3Qs49Q
X7zqs3YJw/Bg/AJXfsdHBxJKQCowj8Fs+wXUPIedgO5h8RYLwhaSLksJIoEFn33X
WNXLSwwJXUGLiogJLHhRjf5aOzHm7+xcTa+XQn79GOwLTNbowbdpi+Q8kJOvSEZy
snbxPhktlXwRjJ0wB8tMU6YPgNwBEuU0EbS04iuLHMz2NSsDJ63+qKFoJn0tmNe/
bw2aWvtqZsHC29UzQIoglER/bORfQztwsXHTZ1f74WBUhd4wuJq6HLDgoBL91sae
cxwhMBfKhfzoUMBK38Eb3wtj+Cr12G5859XHplacLiGSjciVqmn2Bf25Oav0pdcr
C5pSYnmGH7FdAGcao4I/5fuBEf0HJ+ZHYUyPS9yNMbEVSRoJD6A/x2DZUFaaB/UA
JOzdBl7DjDCUs8AmdRbHN53V5kwitCzhjQ86x4C40RHdVZq3jJnIcpju6xqPdpyD
NvKXEUCO4yaDE60amfBwCc7TZhl2K+kWjIxb7aEGNtoWck5Qh7cPbgeOrSk0INdY
SwIMSF3Plo8DAhXFBOlQ89RbP8ee6BM5OeUpVBhJcFVgyGsTBHI9ddC3/ZqRNiZ7
ZBMY3pEVnor66ApmnnsOgsCdhnfxLzFr5UF2hBo5AQIhcUBWMfiwWgh38fMX4e2M
6HKXLLDBxvrjZB4n0r+prFMqZb9No3vYUJM+Uhj4yHH8zeRf6pSJH5BK/zPgtZdd
/cdUf+WujJRVP7kxZtmJLg5QwGjZ8El93GNPDZ0KnKgTFVK0XyruRiLXkb4nKW+Y
U4IKRxqP8Ao0vciCmU8Eq7G2uDGD5MsDrh426s2m0VAPUfrDtSQkpmw5HxVdjLCY
B8rZnKhbVgOFbRfvPC3QCDuMRhuON9Unvn/YuzMG1XBOVRa/5/larfDROFPvJur+
WNAeMVmuEGVlayIJn5cbkO1tsiKDi0w+s40yxLZHrMGv0PTMrUlxiDswzeXmtgiD
zZq/yNP4xH0/ezxkNDf3ZBFkDzlJtBJALSdL7WiUozEkfxGL56EGluDbJDSQinp2
6QXGtrzAxvQv/xJ0eGIY3m6147hgWPUP5Nff8F8llkxufU+tZqh6VgP3THzmjmao
WVDp4UOj9aVciTrR06entpkRtVhjIRuA2n4NRmoh6I9IB42dqhd5SCVPKpgeERsb
FrYztZWnrCk3PKOYbsFrIchbQqK98Fxj0Rd+UMHhPRgTgvPpwExjIqOeQc+o0akZ
bs3o67ICkjtcL2Us6R4UxfyP+QyGyLzOyQzQDst+lVBdXrCPw4aOneEgowTSIxHh
YHTJumTlrrDwzPc85bfRQQVydDpemffgm9E7JPbz/dVYaFPtwJG7c4dNT+ogBD/t
3jQbCVoixB7kMAXW0CyFdQ3kQWDO9xC0zw8LuAqmR4F3CmvfTftroBdfT91ayP6e
M/XekI5NQzrLuDevFBNt81gxebvtdE3f2pqCJfEB7lPtx7Lt6xVPVawQ1slGUMsr
LV01p9wnY044ZiaxUQEULtctXRbOjW+l4oj7vm6qEzq3tnW6utQuFz/VSnCwANqi
YAaUTfrjY6t5rVS377+eKu/yToWp3WNm6Oml0Bx7zSl4k5UiOyrYDcMrXF5HLl61
TY0x12kFn4ftV74Ng3bGHDb+Hd1ROt0iMdkR3JnRwyGO+yD9oaI0D5IuTrbaJzyc
zK2WdM2qS6y+uuH9IhzbhYGC6FE8e02660PLLY79GXzy07XK1yNLAWXRtfhBe+Pv
dgzfkdInvSx+II2tSRo0O4N6Quwxc7DCWb9Z3m0OzM9nW+ea1Q7QAoFT7g1T7+V4
a9ws3X7WTDycsRNetVtFMdMR3Iqdz5iEGl66She2HYf7NtYpG0c94pK/wOVZPy1r
nJIOgiyVfXKGX0BfowciCD7XdSvdIP991jPTLb9IvoLSlcmU8FIX65pYRTLWb44l
k3fwkc26HLL2HWmpOnydxkmKGf+A0koGyGDPfBB8IwMGyVnk2rAoQ5743qWe2hKj
Bt89sVvUvC8nLqi8e1nFjvMsIFtB3EWFxFp9vYsAFgE4oHB18maUGwRE2Q1ZSsbx
AgIYjBlmLEGny+HC4fVeClWXz4D3xBqyTto7vKIjYJmuY5buQFNY7dPeDnb6HGGB
yF0VgofXhTTLLEOrxe07jpvA9rvpuje9G5ycn3ozpZzhKQu9AQttRPLlOvUAXt0x
23hIduGQQe16dyxCIfP+t+TXeIz0/gKtgPJ0wfRF4A4dcgLMZaTUsM/ddQRvOXpu
YpfelQhZhzx0nS0mQPkB8nkvFNTOTO8sUtY01H3X/CnHbBSRyeGIPtnfAMJicEBV
A8T/0yaVwnkxVhOzLCKsYG9rIKiWJ2dGI5lBaDr1IHewFhC0zesVRD/PsXOlP0jx
bA6uPmJqls6K0Fry9cWYN/EAfXqH7/7lw/Lv2T5Sdis3h5oaIedk4iHNOroK8cud
9Ec2nt313/bro3Mlb75JYHFJ03Yb5589y0OKI+/w0xoX5tpWyV6i+rycQzRSEt1Y
GrePkfWd30ZcuThhL3DZSOkINWPynegRYQLv5Oj3SZbkZWVaWxT8Hwti7ilwOblI
UQbJwrQT+gPsBDEgv3MlzpF3rbKQMN7kIAgbeVgGXPwhhHmA8TKIiJ7nlj4xUm+g
UhrGDdAHyyQzXK24XJSvl7ZthG465y4gDKb5sHcuxkybNmOJ0KAumwLe68+MtCQT
Dr35WD/M9SGOB/IVi3VWGG9JMH0uVBqQmbWXGfos/xK9HZlzN0ICcewjqvUCIqqG
mtqxNivYoALHmaSsiwCKLGtS3+Ao7v55pvIux8XwzBzcSiqBeiNWi72V0UCLlCG+
obKuMn01W8y/EKzV92FA8omJ8YDivm//2aVP6Z9bfCSbC0IUZNfPu1CnIlilb2tC
ka2uAE2NfD2HjNDIwnkivvBThxL0LYcYFwvzBfKnRkx/Je6nd4n8coMCFEkoHVLH
zhJvS/+1iWR59scqLhh7BsBOJ+qnKFkHutWZENEJXFwOAuHoVJYLtEt/+/GOI/F0
2tVfVnBPgafhycgu47tyFBaqkEYEN+3+l2d3dJKWYwRf9GZNnLHkwvzEoMvcmwBp
WBPncNsJsxMwZ+QzvD7DBOL2SvRrp0Y6IiD0glAYkewjcIcoJZyDWD1fQc1CrQpW
hJyNricpfbMjFM1M1OT0dp4w8ZnVQtdPCGUxxp3siv0jZum/t4xEcawuyTFK92Mc
gKMTmfaRGzUknzpqu05vuxBbALWO6TIS7geZVd2D92nVb3QDm9FZTGudjV22YUrz
bEXiYTAbrreQ1fqMFLxIOWs4HNfksTjQSKTe2JDk3uIbncWlDjcg4rjrtGVyROML
7sodz7gdVPmlWil79TTiC+zNm5QFBkQEQP3TwLlY2P00kJUcIXndZK77LjgPZ/+k
slGuG14Bef9sBepIM27hypcrtgsz84W2GPZsoGFahnrAbEf9lwzkUUxuuiNnNfzY
x704aQCR4RVBC1T0eqHCrzA6dE3rs3OI8egaNBNSGszNSabWzvdAR27D1uytR71/
WKf4tvSy4dpb+bTwnvlRm66NeQch99ONMHjIMFkHRObEBHapaF4yhm6qpSXtGR+Z
oF5QTUS5MslFe28uf8XMOMDj7gjA02iRZQLKEuipjjIB19WM/zI0EOfzroDHX1He
nCquX++X9JCFzx0szqI6ykrXFn5Jx4qCigtSVJYaD1J3kbRFE406ZbKs3NwFm5vj
NpInH3fzBXFe7PQ+lj/vCleBldQRb8q+C0+ery4Rb+7xWLUhD0rDB+44vaY3ETeS
FaHS3Mc1kW7fTNRin5CJGEGOfjl2w4Vj0CR8XUEhvgMXnveAoEwTKLE2WsPT4k56
SOOqDYwBRyHzvoJlC729dHsM3RcGniNQpBaIImcnFjyWnEtcZsLDiJpp7eJMkIe4
POB/p/1TD4L6+Eq3yeTR0A2+4roLlLXZDGxJ2GuMoTFlJ1/bMyLQuQ5e2m5OLESD
rtOLIjPcj72GCE0wP4wUyCsvoH7ly6P2w8UGKClS66eEIlixGrT7IEa+2sRCkzIo
X0a5sOu6LUo4j/ZKdekU8NZJzuNseLKHBbU5RQxqUf3bxEtBiP32zSBvf8Wl645N
Afnw8P1/1AcW/+23WfoPHzv6y7yFossTBKshzev9Rk3xYHN92oNcwnvrd9KZF0L0
UJNJp7jN9qmNvKT9HyPXGo1R+OCCJjBOB3Qloww6oHxkFn6hXyF7niIspmg8uGdu
OyFkwNY+/xgO2u4p7j0MTSQ7nKkwSsrV83vXfUmNd96LMPQ8EUKTgpcYn28Q1wan
23DzPQck4fgPOJcGnFTxV9A0lsF7WzOldyZ180rXspqDGPqMGJ60jBX/vlaF+F+V
rp86/x+AbYDzk6Ska1FvnLyklzxyJYsL2J7t0j5iXwXlota6bu3y8aqEHtEoLTFj
/sbOeSXJ2T0vSepIfBneamLoTriiwYPpdlo9EDWZxM0ps4w9ft2B0vALr45CnkC8
cZQgVDUmxE1YrA4IzHnVH2wlPvhnPL+1tPemAdT+JPJ2wog98c2pGYVlBLuQWPGg
mHOravxUzQ/KCpMn1oVQHZwhRkGT8pBoVpQCGxZlh8OnxtSlbprj42ZXifUQiagH
LmSBKN0cK/EZxVKfRdHysbj/Xs+Cv4lARqU6UWkm/9xVRzBSIgTdFmfAQDGNb8n2
EG+hDL9igXXxk+h8i1tMKNe28w/k8LOWweH/dDo7njmPzQEBuiG5wCrROucs24OO
AMeq/4XOMkxlIh9ztIYH+ePvhsJnjd4PpbTzpDFGfJwt/WfuttyDnHsL1JpQWG0z
bPkSdfD81lRD1A6hCU+YpjKMYdjgtj6JZ0npvhkvSX1oVHrjowBarcUfBOMHq19L
x6RaK/AO3RYR/GAlUwyUcalKjrkyULmgJRTKQtrQAw5wMK2qrbtl4QgG9+4FfHmB
RCOZOBP02BTSVYtBXD2P2yv9Ae+Mi5UqeeheUlqxlc+JcJHCYiIMtetfrN3wa/55
xTl4ynqpVAmQ/ysqABjIyk4wpeiQuFdn1oW1Ijo0ivPpjtXMEndcx2ahAFXLbAOj
GRKUmbbRwdX8NRGczObTDT2f1eaJVR0vqXUlXxUVSmyD8uh+fib0Y/RmakbjipjX
TRpXYewg50oDqZgKzTWIHT0XT6XrACq3LlBQyFNfC3w8C6ACPbVTI2zMnHMbbGju
cwoym9r8j8mRjc6TDPJmm3ScXb8NuxngAQSty5bvppMzxrAAOBR+Pdb7c4WTRJh/
WvyiDcnXYSIoU2iTsO8C+Z54KfsN8LokSNnb20mwac7roNi6Ij5loWmb1pVZUMw8
O4ym2wLglmqVT5mX/Kmr2vdZbERPJRritwPBjQ98MA+5HNUgIYwmtASGEu2Wt7MK
1jJqUWuKDu/Le4wR3HGv08sFflR1cT0B/3H4Uk4kBKwoSUkwpEVfPB/t/aRz4hU1
NVTwUfrtH7+rwtjw57Yph1/h3sNSOWUndmwgys0SwtqYx2m2sO0TF6PsCznoO7sM
i7K8/+P4O5g8cFNXpQN2n1nysgSJIf5W1L+fIEF/MNLlWTGOef3xvk9929D7+WrQ
Zyry29ngoZTVAq891FWNjvFv7tmqRp8zWB0EJ2oLvKM1aELofXCYd2voES3lDGVi
8OYNrPEw4lNeuL2e6sXKmj371jK+SGetZikwRxXQo0EH5LsXSAca9ZxVfWORaCCJ
vVDpV4nD7x8biEzJf9jr4o6NTSsECatXGSlRukSwSw2ab2Ns2WlwwDEhdAsVFA3W
saKu7VRe8TL8jsVLYa6JpwmgnmrMG7uZijRwO6LZ/ragf4D39ZSKvneLVeYDhrfu
K9oHeS/yvgbQhmHsjQnk23nPWnLYipv4YXF5EYtC+0clqbAYewpH+QR1TGODKC4C
8dWi+q6BTi6atsuxLPayRtdL11Oh0+v9QvouX/UtTvEe2DTYdqLHs1md1M6JlK2V
pv+uuE7Xenc1ahjBm/y2jATcSse3pyJxjZWmBNv+GbOxIlsg9Xt7GeM4r8GeB/EG
vLTyApKCCR7b4JuJLsja9P19PgIfbP7R5zgt8ArDDciS48c1v2+HcdN89i1K/SDN
5ZEchT/MiKDWlfBhFndnct9NdBeae9CkM4cvYHlZeB0tzRkBogJF2PQ36oqMjYzZ
6E9sDLSwrEDjJLMX9uVJtdh4jFiS0uRNgmqWhJ7smV2jfthiGqYVqOAvlmgNQCaj
Ng2R1hA3t4xMypEAc2H+FRo40Fv5Ddop1+S5olnyfIDCs16y4OJxTKPnayCi3W+7
70Zs7kM3CbMdcvSYtbhgzLxx3g5ScLJOQZgRn/LgmYF/RqyLGkg0c/K9oXcMpXgm
Mhvhf6zPAn1Mw177qrkMyP4SIhMDsfa8BPNtkMm0D3XSwST907uYrbHISk9cLGaj
2vA+KTJX4+Waq/K9ouD6AGzaG8CmK34zO97og7OxE/k8qkVYhXoGY9EqOR0ZIJe4
MBC2IJ0qAEzDR2HNvKgr5VgJW2HbgWmcpeNIRGQWLWaU4cVifg2L6Jra27PEiwtK
6ybtt6TXKPJK7slkazKhUdN/3Bevkllt3yGbh2/3zYxsRC5q3mlN2W8NAYGqHC7k
zOjce1abW2gv8HZNZbf/HMS7KOLUviqNS0rmLJmwiVsuIm80DWWP5Dj2A8Gy6CXY
e8sZdsNMUrxMAk2Nnk01laxFBxvTtDtGmVqNLUtaxHgbjV+V65M9dVZtXV+sC1XX
dfic+C/wtPIb2sURt08AIJjDUhZnMWO+/WjzV8dzq3U30+HP46BnDeCXysZfM37k
89bfXycWDVNUu5o7l+INYFNd35cbA9EC4L4nKGJTufeCFiP5cIbrn4BuKgG07V7X
EVdWzfxLlJlG9a/PJKSb81hiQPD6Qo7JrrjDHZAg36rzstbJ6MrbZluFaOXebEoh
yo2dV9hEz7FEQPE3iPevMOuEUwn17akfWwiZC1gjPae7BPDj1QbQZ9ETCKdloJD2
iPwAs03lXbBiTRgWL1F5juUevZ3JiMjVRapu1nWmts0lOVZfLSHlIJ7CoJA79Msh
B02V8VB/7UtEhBZd0+8PZ+UIrXN1BIFRMQvx+kBOWFhTh4EJyko+aJUev/EoD/WM
UcbbxrcnRfA4C12/cm/k5mkdCnKjkg4OqrK+zVodRbAOJgPpS1zoQD9aRc0pPWWL
o9Q5bOEjA1+ZTa26izq308p04kk8S0SpuR3RVXQm/ZfY9AQ+MPUPOfs7MCBZEOkM
FayxmTm2oayJQhnNNqC+aH8Vrq26VNnh6ZIhgksZ2/SlJGqezEa6wspNkWq9IHNm
AyFvmN1zgNBOxAzdK2Pnu6zyr0TwaiIDd8JZiP6IvpxOU0aBgXk3JlV44hbkieuK
kIcPbHT7Unb4csXSXrmNKcGHux1/+wiIRx6LdOgOvDCyXH0oKw8pwC/I08KMlDLL
EQ1CzaPUMnOSDXGr3MBUzCrMXD2xy0B9Vq8mARQfnfOPO2JqgYhf5Z0gX6wwJy5x
RLLY5NL5fZkNtGBcLdJb1WyRmcHIyaD04+UBOJ/buuQvAW4ETRHbpEDObCulstkV
/gerk4n2nzdwoMwOUTzGkan56KqnFZACx+6mcs4hDQPUOP8v/R/gzHB2Zh1T32Su
2Ud6aXiWtP5ZOiRamGkWZMwDT8SlIC4L79F5TooDWVXUJLZMkG83Y5QDeH1zICl1
x/hQPZAm+3iTRkI+3aKXDloZjLlm5/HyS1Rgbl350dQMLhyq98rKfA8IWP9MGcVq
+IlrZI/TQUa9lYviLCUljlDfamTU/Q03JgeTaEd7tYcBEUMVITnLNOacthqqsMqV
loGun9QgBNNxmzqWODAkXyQIJBJBblRllFEujaaueJRJizVbRNXqgTYVEwibisWR
Y148p3hABsqFadfIqoyHl+UzFbCv5m9UCX6EF8OemYrPTD5awbxhslWsKx9alppL
Z1s2jZZA6jXLf3hXJvno4A0AYe8q8omV3DjA2vjV+mySng7vue/0kY1MAxlQ2I0/
beKPXumEmrGcKC7fkeKKeMCvruqbdAHRuKgmC4atwZtTwQJGiz1qq76tmdgLxpkF
/YncMJNM0w1G/3TEtHHfzU/msWArMVRQSxRTsRGZwGCOkERrgP6/g8eb+1J9bSP/
Ufb4JvCzK3F87cuq+nU1ctlgUS+EwvaZBcbMiwJ5NcKoCfqtbM/vuHC62+r0Fnz6
QdTG03umvlWWky0OQvgPBEm/ZySpk+XN5BYuCPMoouCA/LkZl/co+LxBTHibKUaZ
q7yvHJ5Fq+RGhTSKxIgMsltUexlwYZd39Eumh0YkQuOnX9z1+Udgt+XsP3skY7J5
J+WkxXXiudZ6TOZOARR4sk9oz3YETpw4oYT2pwp7ZGZjGmeSsBtbeMqrpL9LASAF
GW1rp16pUUkPjohK3e8hhSkwyG7Q+0cGB8K2mBwacDnxgoshbXX6RVOzU8HjiFmv
z7MRnP0Hso3eRdnWn5rDkqISANoXFgROMRr157OXr0EvqxSytCJCozgFzk4koUB4
KFoqN8k6t2Nh+ILgtD3+hxX/jtrN7oh8EZuW02ED/BfT8ILEXZFBFv9JoWSKDWri
qEFAkaRhXeZFGBDs9w+KqX9pt1IWkTikSQ3BBql8s5u8RZb8qp4JPgzIr4p2OifZ
57xIN4JbQE9JWjcZ3+2Q7kzeAOi5ZbHPraFT5FuZhcO7Xf+/XoNO1UU4LS3LtrYD
/d7gWeRpB2OcB1DHhAk5Qk9ihyJILn+GYHn6cTAFsNKvcd/cDOpVzCvRfTJ1V0wm
RiWMz3fnXT3ShLUtn7+NQHrWoSXGsO/a8/Be1vmA4AcSTlBfNLAofCtdnM+84fk9
s8ysySPOF5HEQ6qbBo+uJCt4hd+lR0rPEZHFojTZ/2UZgAw5k2q049LpBd3y3JOd
VFIFybWe6QaqpJM7bvNfqw4TvnmabB6Yvuz4plFVs2W++iSYVNMK7wVLwwZZmo7V
pBtcgcfKN9a7MFTVJt6vA+9sx9bxCVPOJZZzDQfYNov+ZRAODWQpCQJFvmb/uhgl
dBRtcIeqRrlVVRDzkqtkGW7yuM/+7yq9GyrZsg4Mij4=
`pragma protect end_protected
