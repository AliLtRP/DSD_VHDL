// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
gTPRtfAWCZBKSPNSGMrjn0ByYT49btmJOCpIUlvyY4yGt04Rq1+A60gsitqq2C4gMaCK2SOxiVGC
Bc6VvVPY3Q1j2g8n0wNCrmVmE2LCsCpZ8kN50OLKLlvQ2GfujW9QXinYAI4+p+wfifv0CzMCrjC8
bxHugwxYNuCIqtYhZjQ44nCcLHoI1ixWjs1/7XRE1HUeLHO2/vmMM3msIaEVNiML1eYfuKArlSeZ
ai5PCVB8xXONDhZv+ym1lKXaKxJ+ceVMcObBuo3/nBHKesATm2K0rxtWTFBB4EBR6RzYY3gKwljd
+fsBe5iuOa9o/83o8aMgq2qmXNPz2paeFsm56g==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
LEj4D3rgK2AUJz8kBtj1Ud1pjR1EXhJqQ9epIwSEdDXcCINsuxzYevLoSeB5n0ejtxXNuBsrM01m
LqbjjqQGD2ixKiFIt2Rx6y/yPkhZw5q4ZuTztPyIdUWCQfhGAPzqQJ4IRcu5q52tboMGy9g9MEx3
LEXd+MLK2o1YD7Rp0WondCtDvXYByGY2OuU81hu/zBXGW0ALJ2S9qvpDPc6IG1W+SYC4lnUsUeTC
RZhU+OQC4LhTjn+d5hKWJKLUQGawqf6lcCLVKawwr7BaVxXyw4To7HiEKYL+ga+KLbe7Xff3N047
xCd+2vLo8n8UUoqNxoMvAYS/11ympHyQOfn9C6ZpAWCEU/O7K0EVakw1w6MbkR1PnmR1VnWQx2uv
5/RP+wsrdj1AZ6C2yfYNqDGnDatXjICwmEn9+4ZpTjezj4QlzIzlzFp0mUf/paJHhpRph3RGTVq3
UdON0w65oAuyPFJ6pzOycHcOpdnapvYy5miz83vMlqryCExU7rh496mIcT8qrkev9N4tt2osxUpe
i3VeibKTgh3W4lWUbCjopWA2By+vclSP72fV9ix50Yro12bmNpTyUFHt9jHixeWZrwoJDamAnVkt
Bynx5mA+gUpugGhiLByyhWbbkpAUpCLfgrPpzK1I9AZ26qV0gfeGsKJzxMOOzbCHjLkc81e2GEDJ
dggnKR5FR1ntyxPBaR1Y+kzTF1oWnq8F6SjWvjfcsXv82noY3YvYSQ4D2GWKlFZB+I5RoH6yWRnb
t4dXg/YkhsZpJrsLUvjzijtRBWIroQT2yztq70fHpMD6CdT2vG3R3nUGoeR/QmtNx86ToYSup7oX
rntUmGP69tdWEGFpycN9h2h5z7P15CpB8+beXPVrSxuKeU7Qcdz9U6yDhFfOQ/FdnfW7UGkEdhBV
QkrdsD0Esgqo4XH7C/ECxmgt6r3KN0W52u4MHDJgvR9tuMbKJ2V605qvS+rbdZcTKf+6Hu2b7yP0
OkqaHdD3JpUFbQ+zZHm413I6y4cOtTZhxb1mgaZchf0ZoRyKU2ABzn6NqZVIJWu3tnPp96iNUzUM
9kZGNDwrOljR/f9aPkyi+eQIkJVjV3mP7NQUhipojJGRXZImMT8LM3Q7ZgxmNODeZ6CNB2pDF/rW
gAH7+KCPnDX+tH8iX2YRHcOyMGPMnjh4vMNAPsRAvgFuz5/hL29yQJMT2xPYuEIIiNRkPnd9g4Br
emxG21GIJvlNgM8VyeP03Mh7KIIlWj5FthIc3AlnBIo7GO7z18kXa5IbtU3kimqRR82a1RlE4uQY
xUYBt4qSa8yS9IbeK/r6ErWeZJX3wX7xGyDAnpRXjdTGOU/lwU+cfryyyNs/LhhdFuJaoDvDYCvr
Vp2gDTz4DG+/z/ra6MZf9HvUMH9LKqDzB4qVB2SFlL/UyU/s6kTy2e2Zmx+GzqgZjKYzMEqqTvZF
e/yvzjZ5iTnkstHpoQSX2SRQeRsvxTb6SrARWMJa23VsBkaKT2f8QyOlMgdciBpj+8cxvwDf5keX
fBJ7JAsh7gDaHrD3M0bf3aS0kdUxtTdgw4jnCQSbYh3ddXYfXEjdwjwf6xoMmVyePsKiclDqyHPO
gPfbTuQJoltcdPXUoDO9Y1SuHaR31yNMjY5fYZh6dQuE264+3aq4tAN/LzYxKlWWmiNIvoUFlkdL
JLVFWy8td5UsK8Pbz7+Ekp4Tz6Q2ogZFvbxxs+rW9A7D7bY2SxtcRWYd1qLjantMt2gD/Y7nR46s
habWvrdszdmqRuTu5+19g0JC7DfqmlGDbId5FiIpL40rkAWNZeucfmAmuQIf7f+RhrqgdvWaQm+4
Y/l//MDMSuU=
`pragma protect end_protected
