// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:31:40 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
ATpcsnCghtDzv1PrCLCF+3XncT5ux5aH9TtXNfw1R2f3KfLlhuGDnEhU1H50l2Pj
p55750455ndlb0RFZJpRYAeLrePBOAO1Cnd3Jxndk1oibTNC7F0e4Y304pIX8FmA
t2PUSRBQ85aatvfDwX8oTewXvxNL0722oZeVqA3cjl0=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 7200)
tA31WkPpI0yqc7kBE7eccOJp8+Ks3bxm1rm9/vQ499NpeC2Z/m2r77DDMrqJPX7Y
PZULF2OhcYwWg/nVn8R9r1+EDbW7tMGNjlgEOV1cBhMA7Ont3t56IiOxDdHNFxFT
zZA545pDtrPYuueHKJH4hJaT9XpmbBKhIbMtpDTcuBE5CgflrIyEBH6xUajUhiZE
5YmNYxDtYsmWcdndBLX5F+/qotaizhT8KBm86iS1ZPaifEgPN9T8l92KMVj8seWx
6whjwnRV8GMp7PW7pevKyg/p+xpMOrHMmIiscA2UETpU5l65Mbg6f8sU4A0UvXs1
K8CsxDiuo8ybbuv6++B4tBBb/prcY/XHgegxXmZaWU1A1wY+AHLL/rySeHbMY0dG
LmQIug9CXHGy87XKkhKx+/zJ9SCwJF+/Bf9LOXNx7Fpiy8YLKbphFoxZbdANtPAP
MGB2VYbIG+gw2UKHuRL9dBsg+1kbpiYHCBfSWPxgIaW/eaXJPQBc9agH8CBDrY3j
4N2lSBT+YHieMrinfbARiVuiMuxDqPuJkcnbf9S+KQvSkbOB5NX2RFKyb2+Gvib6
2xJkQQrgDX1FjLiRNG7SVaammjO/mRs65WY7ZFH/2TnXlAZ8LMbbN0ORice3fQn+
tQ5zyFldIaH2WHbZtD3PIqaoPd2HgDjJw6np8ordLIE4DJCk00XjF7FKiFnpyw96
0lWt9AagKNA/YKsm4cELgYhM+TZGT6esWwltpT2ZfJs4NxeJ6Q1JTDQzBTJEb8Np
yS7pjy7lg55nLCqMuT2cuOO7OS9gn+zKrD4hM/Sn0AuDnFIK0pud8Cn8kzm5Uu08
Di+sxGRg4XNTHubyVj7+ns3/+/zPznyfNQ/BHggtbsjb07Sbxd/HjvLcxC6S+IS5
wzOAgp8VY01O7vaSID1ER68/t/EnXu8dwQf+HAm5388iUwnmPSZEIlzV0LeaydWe
kPNlQDg9Uz3MibYIWzaAWgAd3wfF8F3eQHaVo0z7hlCXdFWlHJqdM24bYvLkQ8zd
J/d5QkB3b6ZELtB11durpZY1aLMG0YlVyeBe8NitARRUzsQ2gwihzLwUVnPVVcqW
xXUkF8EUVL0HYMcvmr80aLUkDJun8iRvnujjfiC5OZA/ByGUkfRjomIC56GLSXEx
25TMKLfALL1twhQu4T3ylRmqgwfOoer8OupMeVbRiVRoClr3E/GpSPZUO3ibRTO9
NMKG5Jwf3Hb83M8oD1Eb69Y/cyUzBvEioImsNjFNLnsWFe9axzIfS7XzjbQvB69P
paxd5CzmPZq0EtDxk0GapX1x7JEeHbarbX8UZmcybXvfaNgP67zkY0l4WG24847a
hjhSgD4REmDYoculCVOVwaQ+gG8qWropNbC1dx/4UbA0s+Un/HRRt9DjqflQM3ZX
4yybe0c+mW/4/uvV7XvOizDobBKHlA+oUo4SABxT07eutNyKglHvEeZtoRxAephx
34hfio4JFBYsNAmLa5zxPwDSQl5y3/wKuWvuT3YuMNA7/slg5ewvAyLYSR20SrW2
Twh2+WXrE04b89XtwjH1DiBbNnooTxIEnWPW5B+Z7NbbyLvyk8gv4UboV2yr184n
RkqdQlKjv95CiKq2sXERRsBCmoitTJF8kXCBO7U47kGzZ3SkdRGmmXoX01hot4AH
Oay63ZgIbqqNrgsZEFDu3DM9eS55OSd3DZwftpO57HrrlngVrzWyfIYQpgAp7spq
Ra2G9kU2g9QlY4Bq/Kv7agRqc9bKxYMUi6MTuBgGAeWZd6Tw4QonXlMu7cuZWdc6
t1xpSThAq59mDtohFJozNFXHFQw2tijIoiqyJf1sRFXXTY0w8InUXtKEJP7+9L/E
iSf5Rg1P49ShcrAE4xTiaKch6sTMytU1IFp6lZvwV9Uv14+AYuvie2CqYyDtmsmn
J5t5HmcXXLZkBiBflm47B4gKICb541WJwfXMTkY2i0r9NiFINnxjvPi0guw9w7Jf
NmrwxcnI/46ECevum2TOYb20SvUtSPzCfhkoVWEzAvyoKA7idqJh07jHKm99762l
jeFcDBjESDA9k5rZh7PGEmF7s24p9HtX+E0FXsgS24kU+usEh6tt0kTOOT0Q4KCl
KgwQJfqunl0314k1R5wAC2ObFJBJzRJMkcrvYvfDGIWfR64d9VtSeYmnQ/S/V67e
l/wlylFBU+t/BE+pWiJmeZ69tnO/x38IRHPkcgxO5TMcN8TtH8MMrq+PJrbc/n3u
jltzcNiH/QuY/FGzhRiDXeRy5BYhZ2lZbdRUkzX1Kv+cFmif0GjK0enQ7HQ34gzG
N/u38bOMAX7uh4ZjElZUXegR5dXZt5vyOti+6FZSTrteTm+yv7SbX1d1QueRBnPH
nxvkxb28N/ASnxe2+dQ/AzXX9ztSL8ehY7U+0LCRIF6hPHLTUNo7luaZFDwZfYiK
Jw1l1zq0IHg1YvZo9KnTcfTyLyMpo6cpF3uq0uidWNTnWbr4v8j5A0hhZ0QtPA1C
GAN7NSo1aSj7dxOW6H2Q/n+IkG5zE5O777ldsHbpHp6zURMsltbWLj9bbbdGQ6mD
Y4SlaHlNo2OnOScUfrdVyrhLUuR3sibSmI9WoMLrkSwlY96oMtt3H6gT5/jaS0tQ
smdRuY/F/0oGIMIQZ3oPdE0vraUIHQ/YFoJ0k1BgKWQco9Ry5r/WmDMhk8kXLw3P
+IDU0GPKLdWDVY7Z4IRUtRTog9WH45GTfY6HfQ4bx11FrbwoCllt3XTrOfDBttkj
IWdmFYmJOb58l+3v6/Hhn/ZnmbGDeaI8xTAW7/3BeAY9gHfU8acryomH0I5okdku
lzmdbRAficz1/kjMaZf6Ts5s5C6OhLE0LB81vLV0Z3j91KzSnA4qWbS/ZHRF7CWo
CAWaV9kelHY+GJB58e7Sv4JPSrWmnQ5Q0nEwMGveF1USoPQyYgQK+0FU9aJlrsTa
uNgSo9cKnrwfaxv4kAkbiqzY/GXHRKwqrSBST+bXyI1n8gv5fhQWNpC6aOMG1kCd
UClBogC+FjzAAOf8O9EyAGgtracQoqgSHCtKgxp9ufznS/z22Jq4eXZIMBYv6kOI
Y11BD+B0htDoZO5OatcFaJdjQxPXy8sQwp+HCPcRwTPCUugOL0E1aJk/vu0a2GXn
05OaGzCfxAdcqerHbx7V7sZGkpL5ComOpd+7F36xKr9/vL0wUhMD0KpfnUZ3yd/O
zeI8cpOT4ygEJXzVItxBJCbAe7akbsM60KHNPQ8HPaKmVHXlRI9QOnQ+bVtzN/Qy
mbRmxd6UwHmPoNI9A0grywMuPuqx3YjS02bMaKt+C1CVunY6LEPJmlU3QJ7bBHT1
GSxzx1UxyCSUVSIly3Qdo2HIq8w5gmLb2iH+s4BuMSE4qhQ4Ux+ztG/IO7hFib74
WoSDqWMygmVDL3brC91LhQiM3c3ti07eypEj4lua3VaCwV+YWyCjQaIK3/Vdh1Im
nirAj3zAV6zGcjzxa+14T8KJMYnnh4mlSWSTPgRIH23fBtNWOAX+gb4dqEYf4rg9
5hZdNQ/zp9wv/+L8RnfF4NSUhIwxD3YbmQrDRSFAKDMXFCXnPCW6NKNJ9c7r4Q2d
NbD6C8SGJs6MT6zJz1v1t9XrkVyJ9HsDxlwLPNtwwN8v868d5RU8d5yvABDCO1U+
yvl7YwHg3/g2bsKDzdrWt+/0GTUzSw+uMTyp2LJIs7HQpItIRBPt5USC50Xjo5Z1
DoYlM92TcCFr5F1MeP9p/SLsJ1D5MHmy7s6OlphN540+9bKxhz4waLhD1njiSYS/
Ea8xvKygFav0CYBImjb1ao3WdrFOk8xUhhXiN+P3llUmPP7CZJxzH6SOsYurMUHp
gZqYuTuKzWdYy+EDKhsK3YfkF7x/6gqxDKNuhYa+fb7oCA4CA2SFc4pThAoi6pdK
OD9GI1WMlrizNO67aV6q/3fultN527ZR4y7mITDKT6qWkIv5pz9KOijddk40dqct
zmaf8knSNOWTIJeCU3teemSDo0t6uBJPtJoE2vAJA6shIjQriKPD2Zt5sd9mRa7p
mK7SlcgIGBTcDC6D8T48ivoDB+YXcusp6UtbdSQBqswQIsEtOfEc9hXQvXjj8YRn
lLHwMzdfe9RTVjep0koeiK4bTMMU3JvJHah8RZ1lTw+SFf4VNmKLVFaeY/OLdYei
xfPIv3FbYw+lzRuRKAgEk7oLVFlaIaKGCBhoifTsDj3UcH7zwfZ39UbhzldEoNir
46bd6D58hyGQf3ZNfMNMzrweQCPeKSp7wl7g6vYlF3YR1Qc9fixOWD2wP4M7legB
/p7nWC+XKMg4mH6Idrnno2ZiICdCuxAWY2tqGnHh0KwyxFmCDuQpzGDVBBqbM2PO
KVJlolCtc7Y2AkEWrxsxChTP+yWSS/9QRJCzTX2uWy2BwB0sGtEYzhAUQ9LawafH
vTSdVI3SZ/X2So3Sqo2xR4MZMvuVKifMYkIitw9wWmjiKfTTKpjCWcC+Jy5HGSss
xOazCcpSZvP1RnLnQ7V1mThBEAgjOL873r1UXKx6fGUsOPAGgsq//jbkZOtYN2k3
U0nrYsqV4ZhLhlJcWP5xm8MApeX3X9YZKDotkJNM7EYPTwbF+7mjA5hrCE0yywpj
8W40AIB5TQEYAnv84mGjf0ehRTrkdDsgAsmWC2TbuSlxJo1V0qYQLd8vh/c9EBsn
QiXIFnqSNyWoGE4l9zSfwy253lFI1edRJnTsk3AkLQ4H3QSGlBap75//BV8GQ7aD
0Job9Hq0BGSx8RA1nu3qr5ceWiOFYMgYEGxPYk+o7s6XI7X8xJGH4zfp8Hy8Ln51
4M1BLyVleSbRbsLNMFHkhSXh7GOREN/GaDRTMx1vPs2HUfKYJez16p7cSHQJa+nY
I7PR/FWJHw0SFTPVQ6iBFNW6QYW6m0NjMO8ouQc2Weo4KLZe7i+q6tSOKDsEh/vG
jKA7/1z3d1md6BU2zGnt+h/cF0lsuv2257RI1xb30xscDEdD0zj9e0pK9quTG9xP
R2z8R7AKE2qlOa6CrodJ9wOKGz8Sf98NO61WscLlDJsQcL0L/xeKZF3RgMr+NFUm
MuczlayF/4a39YpbjT6srAT5TAe9bVGAMkFv5dpY2OyKWGpKZfO0D/uEoiRKtpuA
bsjx6Ui/ZvlJ/eTsJfoiBIiGPhMs0tUcKWwE5yME2eMeTH2XHwtlfMIkHojPxayX
/zQ3FI+adHrU1MRKULup6/jFZA/PYLcu+6zJQMwMl6Q8Eh7mFxUOnUowbAtMhNx0
z/9g75Na0z4r9zW1PsC/GaR74OXXiRwhPN1kscnPKzkQC0KdxnxnqZrrzAFBdP4S
0rG/lPISmwtL8/Eiz6fRW2jLTSkwXcfegnRqtcnvK9n2cw9d3oV42ExMhAc4xpCc
89jEBUn9atAPMcvhiGfIL27OFTElJvf0kBZq8w8memf2AQCpCPLNsqNEt7tSkhRh
+xQ+HVojKkeTxtdzL/BvvDmMvlORDdtXKw7sNVfGGY3g9spBhV+8rMtTsCrJI1/F
a1j4QtI6cSNostL2ddsKqXO3Jal2oJUmxEVl2R7vnL60hQhDuLWLoz2etSd09XpL
/OMAKv8akZpQftgEt29+JySGYebTgbnXksX8OfJFDyqf7c2Va6SbOXVk8etHOovq
6GDcWuSnRyMtto9SPzv43yLwWsg51R9TbCX2lzevNR1XM3QUL1DlIqCGtiW0bVZq
DG2jyp/Db6rJ0JUsB5Ynwk0Z19uSKlSZW9s12U+9oB4bPAHE37Ty6ifd3N9ATjR/
kLbfxCjYvRECysWLAh9xBnGwXAtMnPYKxbeq0shwWSS+/8tPUcyY356Nxh7O0/bS
ygC0ZK2EnA0KXJmaRMc8FzcYJG3+tpPqZkoWM26fhTnvZ3HFd4G5L/7b0rHWjtwH
4XppYWnWzP1Hv4F3xNCDN66xDAceeUCb5rp/LN+PycfOjBZW9dhKs2z85S0UYwew
mhB9MCAEKqyiPfYBTB+0N2oZmG8mK5v3Brw1e/cQzSWlsBsEFFQXZRLazihyVhLq
rGVW3cUmqAUs1u+1GWcnxYmycfwSRwgcEmpA7ynkqmbQcnX04fXevsGpOhdetv9a
z48QP91fWqQVkEg5cqGpOKyHtzbfch850W+qdorPxFPa+kaUoKrHTS98sDh+RiQL
q74SiAyQDii4vUByKVLkmHFb7f9yTILFW/bJsQ2UH7ERYMEOqDXCpcd5+/k+qB7p
Dr1sIB/Oof2p1tLY491mipAG2O1BewifTbEkSVbcmO9BJQhKtNEoziMldVql+rTG
FwjJBK7re0u61kMJmELt+4De8g5eWEJ2wvdzHdQYw1BB4ANsl6plVdfLzGIJ23NQ
jSs89GN3I8Tz3w1aIBTQDuPN/dDtqer302MnrTNOrCmbRHXJybjpVAcTnyYrHRPb
Qdrvt2I7S2cRYoU2LBv6JDDAXTg4KU9ZwoBfOhPRYVuw6V8Ps+WahJYgWa2ifKt6
xuW6f+ybawC1xCbuPZERX1R9bN3mO00nvPygLcDE2Novbd91IThuwi2+QZ4V361v
xJ30yREa5k4fJsZi0EpD24Q1tMohgJfDt7zr47r9LcGGlObL1H688rUyB5eqbiiB
0qT2JsfgnGRknS6ufivHmWmpgdzWUT71UTYwyg3DZZ+VfnZa2hY1t7WKR3KiViUy
/5BEgZqN2MAZS3sqU80rkLIuk0BiS5w16ZbBbi1rjH7vlb6n0Kli1TVQZuFJxXOG
2XpvhQrxlZWVMQjAqjT+GhDOci1QS0b8Do2h1q5IgG7P4bh/JY8FHlYSZD7vithy
cj6kX5cfq8dcW4TY22c964xhC5Kw5dLkNJmYHO9WRyX60jelCqOoDwwz30OvZEzC
Hs287dzmD6fmnMXEnBqJCpB8rt5wnNTljsUsSSLwgJYBcpgV6AGV5GSFYipKnNeo
EP85wTd4YqmIhIgcxOcxmLpDinF16eXTEc0di6pJwySjSFUpsolcnOuFq9prcZse
uazE+QuSfZiVqEWb7NGwVRDvnr2T3t7+UkbIe2jobWH7stmdBXxy9n7PSNaY9fya
4OpBS5WR7RcauibuM8qvCSaQPiyEIs/Q/DekSW1vbCEN4MMPjv9sNWtMXujMRa6K
Pl6kxBJn+ejSEPFhSBwMWWsi14NgMkUjPSDzw4TKovTJXxuOlaENp6F+XgLBSl3y
8gwk/KsOVT0RuaJfqQvv+wADJoAMTwXO1+iYEllm4cXnBReL8BomstDSS/6kTqcm
pcpS4yjop6JiNWT3c1id22NpiQ7kJxvh0qGXpRMsUdGQhcV8aAOpJc9iGFV9lsXv
W4PYF5jLpO6rC4CDw0vui/pYe5I1aQzX0eDxseq63aptzloCzt/szfOzpjGuNlJp
KS7n6n09/Eiw8NSRxDDyrA+TjqzNFl3HP214gU77ulHetCLVSSHyxhKfdDe2I42U
6xvCaWPfORc0dmSXzk/p8cVL13i+vg/J4pUCSagmr+KAzmH9A9dhNL4WW4EIYTfD
VTN7MMmYdoJFCKFKlrCqdyNivj5iVnNzKX+ruqIkELiFjOM366CqzZBDVH/dV4R4
xx2L0e38B+nuB7BjM3O89z0cxPXVbvALfnUyT+4HZI4p5MllVVRlvSPTeNUft0pv
bMdBCNq8qjPgkd47NAguEv4caw5V8DrCxmCThcrBLWXRnycUfZKpTlKDYAYc/afE
0l/OuQKMKQKc1lGIZJRgZyt8TrEMVvNwE3R0FXayfX9XPfOP5g73DEZXio3G6grD
WJvHLs9Be90MHUID0jCvyDd0L2fEelLX4b8CkVf7aTsiYVdX/0JZJswQwra4WIsT
t+EPhXax5q3H8WiaAqsG7YkRII4SrYHHc7lYXZ9eTHZ8erfWqIMlsvjmiRfAb5KP
J8ZwUKLQnyNfbOIIJ5am9ohymh/m810UEGXdIk45a/P3Fo+n6cL9b9N+QTb5UF+i
snTbjprUzQ4CxqqWKQCWSu2fELIKmoofX38oTQfxP1QDL5vwCuk8QCG0S6NBb0/j
md5G8rZP/vQY0XDfMUZIodW1hOMZjmSr9bXuuS4FjHlvtvoyMVzAX5Ge49yosb/a
rq7RyiiLh77Uoyeo9C0ag3z79NfkkKNiNbxSdpAc/j2mB2zM/CUY7RP3eZiD9NYd
345hrIBmkAwqg8l2kjljH2QH9i6R3yrCVgi4qiW/CdW0pzxsReZ2e6DxAHpCUR/b
Csu0IJp/LSYeLyAjx3cPqhA26pfveLJcp9r1Y75kxLX3X8WxmWoh3mQ6g7Bht1cW
WKX8JmUAQIATsatnJYH6Jvvm17OFUM3LfZ2jTvA4D0R5IYNpiIH4NCeWKotLks6u
Fh0NjpWGnC5el2dCXaTaYw9o/biTzYt0JnJN+h8GYezQe0A1+eLVksG+jHe7N/tb
aCBTJxeiSftBLlwbHz+XD+1YiQRtOksCONCf90RYOsjZ6lLVZtwNTCY3XrhZBd2m
2hkzjD3NF8UrUWrhDyuJ50Jy7y9tK7Y92avKAjR/x2xQPrEVMZAY9b5fLZAQr20L
EZlqItny4gAfiUHMLEht48kbCjN4T8EKDswlSn2j6/fE/HEp9zgmP9LBsEFOfik1
ei9XabtmxCbsC4zrpeUHraZz/mVNRi+lDkLKKg6eE7MZeI7jNP+/vnbE4MPL/SDS
DTK7KQ6Y8yQcCgtzpd5wDFgwZQGPExvz/XaJ5oVww6GJMHpju3VGi8QvHoftIO4V
Cz+lvNcbB10GYhFEmqdveLfrRFdgTjtZ4X61P1RlCXa/6mhP+DpVCS+W6IyExxii
OY3oJI//YAyFdWOJJzgtUTdPiF6Q4p+cbXmyxUyEowX52pHbtP9HtkeiyXL8zPot
2eqQPOJ/lUWkSSM93jKVhejsJ2iMFYGAJQUctvBeZDsV9RY0VK4t3Ir5Ebr6tpjy
gdt1jgh1tL4fjU8XaU0oOzLk3pbuDvZtfZg6rQ3nRvDwXwRHSiE2+IyGdfypmWYI
PcPjrC7yzeagkds8fBHXcKe7UnICsK2hFoHZ9f4tnQPaWyQL9ouy1LIHvhZ28xC5
J7GdTqIg1qkyFDTQxwpKAmaySSn/t7nvCNFkGCmysHd5WpMen/Bx/6fs4Q/7n81B
pVW0TV0AGj5wZ6wpF/aoHGhPWqriYdb3YHzw1vd/KX6T4F4jCXCTINIhQ7dRMtgX
OTdwrXOHnudSoW4GauUyEr/abpdJ6P7wDlHOaKgR/P6MCimeOtOsqlaplYMEsuPG
fOaP/4gpENqcnV8eFoWXJg1GGBQD76JljmPWXkBO8+i6BGXq2jMLAir48foUMyyg
bbMqK8SE9dZ10pj5lttQB8viLhEjwd4zkgM/lJj3AW9n97GyrSmFXxCMWTSsDMSF
Daj7g/CWxbTpJ2yrZnZ66ra+oCQJrFoKixrycFp6dqVqiAlWqoVksmtafaWLEwPg
gMJAv3kzGB9P7iwHcNXbBh6zinYR4vGtMj9a313wTpxo0Wnj+M1qPo4TBzvx9UMM
dYAx4WQeL0w+sxVDJHUJKL1fB5Z3xVJMDeyYVQ59xFjo5lP/SMgM0y4RO7T0vezj
qShRxdXlD2Npn6ZpnrAJ4CANltD5iXlXFShoTBvJKXHMdpBMDOVRxe4L3PCNMFz3
`pragma protect end_protected
