// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
LodrOyL9pbOG4UWTTkLHtGdmpoU2DYK4WpW7uXxKvpv3XXhdUxh9ERXwO9aBWwN3goTGGysTNmvb
Jpv+Pd8I6UrqWrPlIhE/Q/BI3pLyQV3MHfEjHwbFiBZxLaCzz2Zj+VbiOjJpqxvMCcpl9b+RgO+T
YHvyoBaxTNMHIdf9Yh8DmdbuLGB3mnS+VYYUU2dz+TBBXYGeVnrWK5nDVFtZ2GJKDZEMfZ8ufGsb
+8+A/eEI91WaYMu8i9Baax7OvJSq6xLqs+9IrJNK3WBf8nz5kQ/IkMl9nHcvzY/uh1S64liWSq04
7iuBbUAlXiBgrq8iS6RHs22ICktp7PauqfJ7Gg==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
W6XNn6Y1+InSwxf0Eek0V5J49AJR7VzpDRgD4mjRh5AzN16mWZSStoBv+2u+Xl5JYUapylObR8nT
Ohnn13cudv6Vz2agAVLK3Azr+pkTQX2XfIdrxA5TtfkxMMzgqCZ+Y17fsUhH4n8d6fbxenBrhw2q
1mCnbLUmIB2HXHvBpCQ+Z94u+6GsjksEd2DNIDYHXjua36edqZbw80YbJYgbvG0qO+Z2XR/n1eaz
tu3A5UPK2hSf47RTUKzlbZSmHZU5bnrEyMgYpYHUm/Sd75X2NU94gbK7Xyv9vv4Qf1n0/zf85PBO
03VXdPoRYXTIBkhk6KMadTuqkVlTYt/jAReYg/8OJ/vedO7kpAiuyDHuLASEPj+GxaOm0NbjcZUr
nwSm2XeRJfWPjaZPMYrEEJmX2y6vRuE7VyvWyf5Vfr1f9bf/ahZmUtZIn+y4rEknb2SOMfarNtQX
oSPRPq/MbFxvH3pAsxWjTMODlpbYsdpm++IoKLtGU2qJ4WVLKnaD88BnPchfZxBiTl74pE6bHdHM
wK4cxQdN4oK2eTMkC8q3Qixf0WDtCP/qgxw1E3j1AUeQEL3wmgzswhJVuoKPxMcLvyMTbTXBk9Jp
dmHlilYV6g8ZhefPqyyz/dMrjijiU+qur7G+Ifmw5dPgN5vX94RfOFtVEWRZWqfTzwWtJ46C4+r6
GHbq/2Q2ymm4iGzZtcyK3xpaAzvRJVfPKGYHElOL1WcEhn46qhfo5D0HyJ22db1YgSy4DZS71iLd
qnmxMlJhBPyS9yUgJhrgS12n6+j8osBFKJq8QGR0YyyOTQaRRX/yP0kNa3GF5JS0Gy5TeQKRzwrY
+upB2S8dEZfnrvmzC13OpItBnf/jzTKSx01dSRj/C6qn6V1sqeRyCwYDhDfm8tPX4Q90Kys556OE
Mc9rikRIL2u8hnzZJdDJqgJC1snNhWUY4r4QzhvjPZhNNKpzUOXA/sCMmSvt8ZxJvzj44TSSujUc
8e3ggh6kG5AruF2jb2cK+0JG9WTApl7/s/rdyrReucPD/NX5zA8hBRj+djU9O+HC+EJxwjJBsRa9
Xze30eQJtL5bjAuTkvD5DXMYQJMAh0JdDGiQi+LJ54Ntrmolh9otchi5oHWut/7gbULis4QpEP0q
CXT7FrXnxX+RMZWG0rkIhNUli8kjRWMdeqBZb4pbQEeFkc02GPi2H6RkoLfo7l9VjGMgdeIWJZmB
GwRPnxRYkDOil+tGPALQTmxojyUe3GCtgcRmM2PP0yquu20GyCV10FeYjWJ242B1dSTWpo+wkzxG
ThGQ/yMK1qYK0Y381dg4W6WNjzaxyixh/8QA9wS1hWgPiPbs9uGujGzbKw+8tYqXmhr8rEVHCcg1
OojRGKPS5RZyZ0/4bbv3taX2TKkPQ3rVBH3j5MsTtUqSjLrQrclla0GW/PVIKsf9kah2KlbDY831
1NUG90OhhGgpNV9CcZm7bsR7v1FCo17xuAeMxqLknwrXDv9Rdk3HSo18yoWnZ4a7nSFxDw0Wj6WQ
UWl2QyhjzDKsJtAJyGdr1q3ZTHUOxif/1GKDrRJlc+1zwUl6aBciiSKpL/xNDQ58FuWXAz2yKTnj
ueupDbwDP3Cxih4OH7s3aUJFRZD/iEXG042aXpcPc5ahGaqHsQLWn10/hVPKTO81AmmSp4eJ+NIV
gAzJQTqh4U2X9txHuMd7jK8JFZwDRFA/91FMbnFflPM0tAtg+x3vw73LxT4bwJ41sJ3i1AJI6b18
Q/44KyY3ACQbJ3rOJtOD4tvalvly3Dmgv83jDU6uFXSfB0B8PT3EKYetzFAvuc8GktMpgIqFVef1
sfBwWr8NJxx6/juuL+mgjGFQQKBCL+15VH0Rp3ABKmjhtGXnbANdBW+TPclu7MwALIalLghCKQpn
bHdUDuoJS8oqHbRRmFOkqCpt2/0jT9Cf4K1NEyKqEpc3E0CX3zQ/ZiM4NXCb3/yYMRcz/JgpgU6P
D4u+gZqEYpnntpuGql1Nxu68K2Sb/yCbF2fZtoEdSVGTVNXCnD+ExLDhtlWKpI8lbOIAuf5mT/E/
UI4VCjiuDwu1mtAs+f9t7hQEAryXtqohTNbzw5TqnmT3fmPSA4oLu7fGGIwD5c4QWZxUhKSqqdLM
kACxKAOkuG40My0bN+f7eyP3FNfQdB52OeiuOzO8hdj73tNQApcLH3tI7u7qEKxcAfTrDOFEWP0w
PAiP0JNGve380qzOHnkfURC0vfwfjEGE5HZtpxHfORhR9/cnEy3oglqzwy3x5jGbN1RJgAb5lZqy
TJxyWmRBk65mUCk7G1Up+pK4drxSuCBJDAkcncyQ1G94UbqwwNcVPL1p434l5KAgRb0gnBobsgRj
0obWkDT3gFtvb+HKMZJizxSLvA859fESpBZw9+6mses3D3TYnYJlJJJx9B+R1FPqfvkwvweTUL1W
LHhUBjPuANR87iZ+ZUdW0c2Cmc4fS/GwjHHZ+E7cMzMX2kQpZlRzPfyvk1BFKpPRZfd14+DgZTqM
3mQwiHQDQGWIvEj5EMd8bPsbUmqUlv+pEiKN95ZQQchiV0KRFF3JwfTWT3/2vYRbhnR5nANEzEys
4ITmbj75Q9Tj/sQ6L4BLbZFJY4dw03soxezOqN0YJh61uhM9exp018Ps+NEXMK5br4kLm4zBFv12
Ih0SoOmhi/GiLwygrLkh1jIMRA8Agbh9kxwcZ90IM47ERl9YtN1Z4jjcQ8DyzrcfkhMwg4cfWFAZ
0m6cAovICLVDcdMdlKtjcIXrEpKXG4xOz8vgpVrTmeqfBCM93wOo4vwiZ0ENhdeuPen7vcup4vxe
1F2hoJVx7gkv/eWaZzsKbezOESEVJU6PXpa78Weln4qo+0Su8BffHLBcVNkSdil7HCYPGExXlYPq
dLwPzI+2lFvyDJ574kN8Za+CoiMgjOKgXEBbFAgUaLgNeiuCIIy1dqdWIpDBexsbPsxL7AJMzDyW
KE5NIoNJa+eA9dqtgD3HByfwhu5CEHaXUWZwmFWH2+Tx1p+HtxL3W01WbRADRG9+K9DGb4cIVpjr
sEmQWIhd8hD0gLO5zm2TOubF+NOpky3M29pFr9yl8hskiws57OzXiLAgyWSb0od0DfG1BtIEHb7E
ssdr/0ukKsFZE/hFmrLfgO1u30sGjOtGBFtJrQuWSGu4Icq9jwZgVXemvdOPPnq96bx6YZYhjh2C
Z7fcs1A81GuisA4I4tYd/x94ZJpYEwH9yunp7Mb9v6p1+lkPu8iXF+xv91OG4dkK+qCi4Khq/yLk
MSInm1VisZzEPRRcmea4PTLjA1RCj1MPHHe76WKYG/ei76mmP3BP+r9KLt+2/Dd8foyzLjay93SE
4WXuBlbmIMEHFLYdsZt2Gi4PWmXO6OELoLQO3YuBHe3p8fwyx9gmJ1R/JjW2OXH1LU9Ea3HmdVHv
clfcRs+6858AhrUYK4DKWUF6VTpUPSqtDlC81vX8DOok3T8/IR9QQ8A6IgBG/LtUVysiIzNc0y1W
okUvQp1DD8z3cDO9HrTi5d+6wO2yav/fKAM0fTUFN9dGKJbfAGQMRwC3brX+fBq9aLLVajok+vsr
juiDRwS+Qoh2cQyA4kwk+0gbmC/H2gTVCLahnUAwixLx7p+6VYUWjQrB9rvtA5FH+aNF9+b5wNU9
iuyyk3N9g98StJx9g12707TVF6yDU3w5GsvKOjyeogYwX1GAJbo7xnpiOm8njMH9H3IrlY64vZ3l
rmyygbhphR299iKq6PRqObhFMewEWjx51dJuncCzDy0QAOquUW9y0EiYb5lnVdEDcmaG8hyEWXZF
MOq73AsZSYJIe9mDNDi2Ab952A+N5snvBLVRBrIWyxWtl9Rkc/VE49Edml6cHZllSS09E3ktSVm7
J3nn/q3gMW9kzfhnXt4v5f/mGxEpA9172vsC/b4ztYEHfWL5LBsGjlkQmKpwWMcbNVwO2MX4tsww
HQSMXGV8bD+hSsAmYYEQcUQkmkOhcKjT909auUDlkC5tcvOueNXpiA7doBF2gZC+YkCceWtswc7J
QhVgygR9xrZzQ6epYbHkPEgmvDorAt3QPqlQpNQycq9oZaou/lLATroG5+E/SkB2H6ozEUYft5eV
nU7qNJTRcqX73s3HG4CzO8ObBiyIl3kvtnKcR5qM5TwbFbxdYzI6zIh3+tb7W3PbA01/mfIrWArw
K50hMxdZjmoyAKLHEjQqHGmX9R7U5ICur4GqHtwS9Nu9HvIpKrsTkITGnoc+iwHkPqsbeLRXSE5U
BeRaHjXBBvwyjG5gff26InbnTAF82s58ZUeqt+RuzIw5EgutDwD8siSj+aUf60nLMb6DZB+IgNB8
A5MZgZeD+a5Fb2br8DcGSwsPMayNxba2Fwc07mMh5m/690/O8tayh2G7ckwYEkl2bKF+ErDMuJmj
ajEZurT0melDxvymEfQ5QP+iE1KPWuN5lE0htThBrV9hncVGZz/upBFAKcgBiT2LBGsLlsyeHXiH
PtNqIfKmGTv9IeK7L1lK7FYqkvxOHlmGPqXUeiFnK3yGvhsjMm8NLJ1Wg8BQMFvJgALAHmXWU0Ut
G6GUKxZUpWmO3srrCcuiGo4z6wFDBLscNvHXw8km5nECBapdPWl7nlDQfu2/BFBp4OHzooTNVDbD
rnPKko39gkNmGuvpNKkTzFR24zzehNDMi0JlNMLf1lw8Ss7w50bnyrnqx6Lvz1npvyEdGNmrykue
HtPD/g142ZwqGiFn1rMiKcpxhX3cKfEda78s/4TUNyPgLiisDFiZbknhdlTqR28FYYVbooOVtC52
fB1W+QQtQIRsTbkxaTlEnZgrVmhEv5QShdDsHwgeb+b4JHcaKpp+KeBUnBMkyd9tGpGFHmSIcvCd
XVLarmXXF4EuSQ/jq56sV9ipkIRpGLSVsgr79niuQdrdcxa62jNeBl25utLZuOi4ksmbzblPzdJN
kd4+2gJfSpNAiCXu5gUFB0zjij49CALtowGS0MP0tMu8YgCvJN9Lmkoh/OJRMy1BfIsO9LMyYPbv
VvRKDJYyZAEDD3MuPbbH2pnuuza50HIUa2aRTn4SNlfc1Sx82ImfgxVOGVK16cLVenueaUopCrJV
XNWmKkzPcjpKMHwegGsJrLH43htFp4Ui063b01NW7Vo+YSAYUVHPHgZz5lMDni3vD70bzg4cQtlU
XNNhFzwdVIzDS/NpSo0CTJanbEDghvqe1y3OC5ImKb5X5jWKfRgBDSoz+fRMYrwMK5+Ej+T3SzBF
DIObfpQc+SUFtYHs22GjxoVGzHli2vF4frfoNjE0MTQDmB41oP1FNhGqPX64kKP1I1QsScJhoD7I
bEbxeYlwKJU/p9BI5TvqV+qQPbBzAai2kRtj+p7clX3VsdSwf+m8CBak99LPEXVvF+uzA8EgUR4w
wrGwj0GWt63ytVMyvkHg0Yss8/cIVUwaKXIQeSSyUzulabJQvDCjhPwe7/VcnJ/OMx7Rj05zb9rK
5XmcrvCcaC6ZtD/PUziCTysB/5nlofE384rpcsDCj5fC0DzEqruvZ1bw8TrTU7gFYzsupTBt9KmK
HLrGtQBX3b7gTrbsvucNSR9ZOWwtqiaIBNRj0v3bEB9MVwEV5ES5APEMZvZQ0Q57kmBeEqi3RoIv
TePDhXot6ZX5FMrlCbYXM6oNlWRs/NokvXgQZmrv0KbvNgxnCzYy52dk1Yr2hBXz0S5pc8WITx3k
AGHh1T6wa0hzZueLq8teNgkBTm5se9zqAvuZy2sjHn6fAJw4T24d5z6uHWoUU9O7AdhUe/eTaCTB
AhP4kFlOM4pKXhlwmca1e29Rscwx1GhTTvoUTkZmPBlzOYpvLaD3+BgMxqYcr3Rqd8WlTvxH0ohE
jKJ0Z8pnnEVUSX4nHISQAHgfyyRG1OUyRtpRN+GIeChsVspzFyR0lnyNh1kTbroY0H/3g97AYzHw
l4k4ajsAdRizI7y+oWyndGRQhyJq4/pDfOXQqH/Z1V8Mr6+LcOM0MRXpqTFzqpLT1pW9B8qQp3Ij
mQRmoLI9ThTKaSKbDN1MR74PNhJ9SVBiXZzzn7tLl54hs5C/rwurL5iOn+CbMgOIaShJfhF5XQmT
inBxwIzBZ8AvY9Gw36n2gucDccuQZojX7+03wLFG+R8Xtwhdbej0/9ornP5imlQTgl87aVI0u3qc
5JQZx4fx3PCSe4sWU4VG78bNvtLvVpE6t6OSF4OERyQpqTnR1rsbSaJDF5I329T4o+2/3RtBisn5
oAuYzbvTzB7KAVxdXj7TOH04qUw4xJ6cFBfYKNVF3trXNIc9kcoge6w7pnA4uCzr4uJR+U2Z3Qw4
wTvMqt1q1OTerw2mbLpgcRE2Jr3QPDOiZj9WpSTKRbXzXsuoBfas1z6jMZE5NLDyWTWVOnrWvoD2
HNtBaC09RFpYE2gD7UzHJv4gjTm6+b819YW+kwN/Mn5ch7PoQn1zvuKWzJ8Dk1F3cAMXky/v/i3+
X6dYiDWQmwgnNd+snVM3hwbxUhecSVHh4RYPLIBkS/lv6pvpB9bJSWGSa0AvYFhX7NMxx9EZsVVJ
geDFy596AzVTF2EGR5Z8aEjtwsyx2DpEOnnolLoro+juC5gQgJ9FPsBN3KSiM+T9UvHmaatrbvy6
MTvbonWNNHtcGC0XmdZUBOoNIFNN/PpX2krEQtUg8z54ytKNmllszvXdPgNCASJVcRbyhLI7G8aT
JKG77rZTOIg04ALraliSMA38hXoUv6mfzY0RX7g0aYxzW9n4jD9g0vWm6hU1FZ7khEPn/dgc5BNk
uysiNHIfHMwZ3zMFyeB3r1TxaCkB7Q2MWRpHY96/riErNOTOoSdGm/RzsyH4OTGsVJSixoXdZhf/
o7j+9Ojb1noSnLIMHsbpCvIaEUR3mA9Ue6DL4zVtj2oMrfyxBNHvj6HHBigzqehzLN1EmVn/gJ79
os1zx0/j5JPWtq3BF4OFyH3Iyg5lMkiAdVzOf8tOgDdNQJptQYZg16wFSvPYq9PBzPFcQB2O91Cj
jA1Ln7/HnfilbSv/8fDkDUqffdEQ2/pkTBS5cWpEg1Mv39p02kWZwRnDJ+xI677V0Ca11UElo3nR
hc30XrivzcNs7spuTc42QCaATkMFFOnRJJ6sXtwxdrHu9ziMgZtiZc0EZeSmI29bR7Aix2fP0FRg
e1qSZW/3npDhdwu/ENuMoqY+Vsv/aSYOGVgUJO29hGM27a4lMgOyAp4GoYNTEv7g/KpeqyBQ8Chb
wLR0fafzzTBb9QYswCi3PTI3CR9ES5VKa/MHLMo9t4vDFR0WFmerCB/d8BsfHMJRvMs22cSJam/W
nnNq83rSRkRikJCe6zE/gEGgYqHEUVVxFiuysSp+Lpa/22baB7+uWoY8B7wOwZGxJdDiu/35LvN3
TG/IYwRWdrsfMgjzeDLSyxA1OAFuSE7yD9c2suVtj/wLZO+QEnew5qO7B676+hXag8dH+5SWIt9D
XKz2dSNSXiFrDX1n0RayrsQWw3VHgNO4din5d10cTvnqT90mS7rRDMT0GUKbwFtJTRH1mG/lku0E
NBkt+u9FREHSb2rE2nPO/DmaO5Imt5D4z2XWm7+lUi3pfzS4fpDg14eHilxcbDFdXxiR+ZvR/oQ1
glPoqQEHqEK6JKpiBAJVqN0GCcGK6sKQk/TiK4cyMKt2d/xOyWKMhdJuQU81EOhuzkBGq/vYwNph
g1lUytQYKty3uZg5GjjnsZts/1ZKmH4rQO9fsZeqSetvzryiSVmICEmuWMHAuAmXslItZqB0nZpT
WFaVHw1wC1vYyU2BMRYJA4LKm65hrfH92t1UOJCZpN5vknrARcWRhy+a8B+MxloV6R4tMnwubUKN
PBIJ18dQtubKo6yPcXyESgSHdMut7djOrfk/K80TxdsYx6f1se1pdR8f83dZCPg8sfw9jyWxN+Rx
yVi7mVACO3TyP7/i+lgu71Hb6fcmL1IpeF/x4R+s7dEXEpc34HS9tSzNxqGWOFQeof8l0rfdqqK6
b35S1dbCHFB7h6pcJXaA/kRWG0liJq30rtCm4MIyAwBKHAdvRPsyFneH/UrS3bNZDzGJUkoUVid7
GvodBvKaZNRGiJ17LRvMR4C/ADm3aQZUep8aH7JjnwFfK54qNP2wRWGwHTvCJBzF1NyBMC+nSGKv
1rZDlV6AL8I7xOt5rdtWzu6W+XO9NjjKvX6uPE4myw3x3Q9GPRQwVqzlLDWonKe74mBDK2hk6JkM
nxS6ca+yqtVlTuNdQiBiLLiSPVtGyLWhdcNjVc21ADb5GozF7tAawJ5+4ZJ0dVhQ4kNrp5P0U9O8
R5Z+JSwpvBsy1zooZIsrIZbtF/AI6fjwkFP42pKMugvV547LlhBAjlhFDUVl5ylB0Gpq/XTjlQbe
1ZdvpQyYPPoTdGkrn/EoRKistCBj63SyZjiu/JAVeTEYF/6wTqb8b5Un3Y3LqeMvmFggDkVBBFyc
kadVfbU87ZbZ7dKidlW7Z0OTlwLf4ll2ysJADJXf+IAxLW4XTH6y/iaqXFqpFuyptAvGDd4gnucQ
54bMvBkuanc3geQDp+WuB8S55nX0vtx0IZgNSvsdFCHdi18phpbj3ZmsyN9zoNGeIwOHL54nl73t
YNaZpmAjHn34FRjgo1CIz6nklsRKm6M/FuOfcepIuVNBCEHzdEyWY0uEbVqCqQ4o09CvI46FtxKx
O3OOrWmkUhlS6ObXRWPUc42EiVogbP01ayFQWbBJs4YYIl7euXwYHFix3xGIk01V/mVZ4OqseEhf
itotL1dDcPBacdjEzKRE0VKvYZ+HwQVa4GeHbX6i+lt7UKTDRGyiaXxs/xNSVUBdF9VzL1QM9w7o
gjfjPvvNnUZozRgrpBXzpTp7zd/y0Em5BXG1n/iTU4z5X2u93BbI61+jLP5FFjjCBWejueffovyk
hbtpd6VkyR7Ggshd4JAw0ilBznOjW7qpJUwFqnbs3yK2wR8fOzIB3X6XyXxKzTRV+N86p5MQTNme
N1Uvfiw/iIAOCMizgTiDeh7YhD6xJYG8KkfUzheci75ARmSdLAtkBnDOWgbYlKdVRP72Ffpz79hG
g2HEePKjtSd3vVf4iGPnntBx/jOjtAVgs1MgJcE8aFbaspwWz/umSyrFzrW/5IMJs8knvdxB5PGK
Ddr1xREpQaEptMctr7kipGLHEAWJ/eIlsUXeyLy+T/TwkQ1ULTrnsZjf+FoHMDxR9eyJdePgmsba
wrf7mx3d3Y82yFd9ENtjH32VIXLdVRexmLA+jW+vll5HWT0k3ncmBCilLp6ey0bkNWbZtz7w05br
QO2A4nkkdKq2oqpheW19pLiqzChTWxR+AzJ1hiFcQTR4MA9oXxqtjzV/9OECUETiC5gOs14QuMs/
QxrCA7mvBG34NPBNjzVemI6/3nViWqBhjDkBD3h+dc2RyN8NlaO+Wa6bD+fBvdd/pDx5y0HDsvfD
FNWmb3VA7+PV6ouDijhOWB+cMCtyTE5XC/FoMHP3o66RIe3tETKGPl2bkPIHae6p85LkqWBRsKvu
s09OE8z7/LJM0Ly7qKCFfigPkLunciCZIEWXm3thZAtvfbWtFdJlgi/CFnERzcK4M7qvnMI3aIPh
WfGu6HGvUDzgQ5TWvL4Qb+E6B/8DM0lWAS65zs1rF9OU5KdOA0ri7JJBgcBzBrWNCZGuOYK2VQR9
4rsbE5R5olEsmLW6j5MXXdrgjzATcg+6H5eMywt33G36B0Vyr4uzV68+QR4I/55ZyVQ7swMcf3nE
duHOPZuCRuSbSKOGF2kk1untbPzMjsrNTPS05e6OddQcHjIOwu8Cz0yBmtIEPGMTsIgLJwAfxO/u
Mgqx6/OGN450wTTW4ajOWkHp48Vb6cGRfW8R07lZO6RX8eVDYK4ArubYCf2IqAZKYe+jj0jCl15z
dF5HB73LDyDKdX95XbE9URYs0K5u68U4I1HdfQLCBwnNVogeGlSEQUi5sb7pPadjltlRIcwhodg4
IAA8/NZekCfFej6T49fJtiIhyZlW1t4qNuEvnz21VvU/JamW3UdKW+kCK7S3tPlM/LgOuNsbijy1
V4+B4bAl7ULVcdw+I3jj+8H3pH/OVIYTRofwr1huao9Fs1A0dY+cURNExs8miLrJG959HlYrUgI2
tTaRrh2lPfrtoT0GZ5qZdcuNiwbXTEV7+kytgGkKmez9YVmv2iSJM3bC9CkjS1gVdIoiSzFYIuDo
0u1VTfAycc6iLmoFf7s/a+d3B4i0wXUSLZugipULeNgrwpPDRmZg3nrrjjYRXyFeEST4OWOgqxoh
yULNsnpDkJjrBiekGB6WLe8FbHInfvFfo5iVVCFZ/4N+Ps/ak8Wx5w0kM5ONNq+dyD1KXLWqUTLQ
WF34bjaDwL5W2LNO2vtkZYoMujivetIL2FTkUdtAtBnZwPRBjAdp1NBoL3uJGNF3A7su35xMgf+0
B9Y81BGUJraGLdTu+wqX2skrUYsA3QMh5lZnOucNA/j05LSVyE78xJblYP6p8+6Rto2AyZzLXo2/
qoMBxxwAMQ7fDY79ZigtugzZ989v+iWrOKaLZZh8zj3WxsoP3cbqv7xvcqpXytosJG4Av2wB9KtY
/0QiepIEj5la4UPjAE6XlETZBOtwkdVqHW5gewm171/+AHMT3PWFnX43TlmQBIU3AYJJmgW/MIAW
IVGPsYW5A4WwKSSyA0t4MhDCZ1oj0eD8dTkcwQgOyaiejhVlJEVufXbvYeY2F9WRH2bzwAsn1zHF
SycazshZRBcuh7fNLONAxNywBkxyqANGjzBpdRTZiFTaaJ88ERbUp2NQ6cA4pKxtHsyl3IvfPdQd
kx3ap4qMtgYx/wLOYRfrjQ0WVCw2axuNh063VQMLXkaxCdupUgBcemLz8rC/mwSb5OQQQ8/Irx06
CtXXo4+M/ZlXWx976kc8DKwVr3IgqVxyWsqJiQTcda5IW/lhGAM32M/tfXd5/51LTZtV7ovvfrJT
UigqrkzvzRVtHzZKX0RvxsRPWSKv1+386ri5f/Tl15VFHyo7acPAQuL+yEwFTELsm0M++rdkIdhD
UF9jOs0nGR7F6is95Gw0cTnhvFCZ21ZsZcKL+6VUEXzrTGmlNVC2ZvU5u4yyMrKNUIRjyFhHAKSk
IT8mIBJDZWym3O81MjUNaUwY3Qjg7446Wj8wzCuHGwHiDYxCi0cbU1V3qib/JgyaVIUyzjlKX7XO
V+9Mp8N88zat9JcnTbWRVFF9d3steLbxRhhG77tNZ+6DL24DJAFLMdEE2PSa6q8YT11CWTWvi0H7
PnG605+6Xbc4Z+w+OUewoDWJD4tJJUaAxkBNIL/NzBRvNVBMuWhiKOOsGRsd1pQPWmy33jIDLetP
zTuiaAW1ROBUYBOpTz6zEPLoc+WS/oLNCGSTGTbVwFKvOqkHKMS8AWViovBYskcte2BregD8LDZf
bUG1zMxvS/MRHBLJfVtbUCpGeTNDsiOoxJaeLpy/lpDREvpE3BNoPw3cVEeto1Zjz4CkI42G0AYl
y5gLKapfXrAIYnz5HzNl7r7G7S+H9SvcxSXAsEtAJ9/N90ZCET38oK0/3C1B+WxNSOqaevNn6ChL
t5tLgr5JKsKTfuQIG6sm7fXivn2q6dUzqaymQ7eO6yD16t5xt1CR49C7lr+0jLnxyxicvB4SCMjS
wv+J8FrSIftR5Pee4ye4/Mpb/yaUvUpdH4WsiXSsVvOKI2FevlWyxVAkIjC0z+TFHVxDiGIHikFs
Exnt+nLw9HHNrxLUPD6gFzfpPwbfvD5FW+ysw4eXXEkzsTApHHzsvLLLcw4Ixy99/pWnzQOjZQ4D
v0FI+mU8UPOzB1M9c0hpUD+dU0J4Bg8+pbZqceOZbwhJs6pyV7o7XprAT1rz+bCAfnzjdNUnV9qT
tZTWUi57c2eTjznFcJyp8uDMF+XUUAaUv8GrHAAbbyg0czMvNMrpd2DmHAfbzeuJTIi46LmichCr
5mspOpGBaRFmisuGPiR7oam0UQvr1W49W5XlhgYCLHpQGXEVDCE7qyDdeJarxbEjwnW9enoKP9e0
50MyhCE7KHG/CU1w6egsSzwUm61OkSx7hHKmumtdv6U8Jd+P4WMd1opLJCUv+cQzVfCQQcoMRZQK
ZoIjOgagGBzKewgS8GYgAjyatiRefKQq88uFM4imDyeDPRi8NDtSzrbg1pmxMkHcUGeLUMdfHG91
Fmtwzuver0w09gmHlwuwP06F8Ko77Ca3QhVapYB3o+q6b9DfnhRt1RaDPgR7pKNlRHnoM/fmVQD+
BBKOajuUV35NnsBOXr+TONXuXqpQc8kjqyVwxAd5/MrSzkLzBLmlLfs6XGLkY6hRjvR9k+R5SreH
bgPizySe63qGsMk1Dm8dc+RS1P3fCe44M0G1w4xERhc7JkfoVcZEwAlKPlpT6BmVzI2Ke/wxHup4
0wAfyRia/DtkcLIQXKjFerFFSG3H7qEYm9j0K4KGys4CmvYKC3uLNV+fAWSRi8JV+miISxyL7U+D
iEuqixhBe4e73EB1Z+4GxS3A4DoJe5vJeRuhu/UcwFn5vk+YEGr4EwEUjmCI3WhP4+YBS86bcWPD
2AAlAVKDShW0+EiqH7kQjmXRapqVsfEnwdAGvRMj7ENiiop0XKMfrdT0Ck/ar4KIhFHRbTSztiZd
Oq0X70D8eXfbY9UzPv+g4zKC9M6TjrOMj6K4it5SB8g6A4HH+hvmMgqFdp/gg0iqubqFJmxWjxUU
X9sDrtgfo8C1OSb1DswrR3EauhHsNFrjf4KGQciGc7NvmOGfELodXr6u9eKPRyEtee28K2IWQECG
Gx0W80Wp8v+34XYr1/QlppF/xCRebQ9GOpc8x4O8mf+LGZp5Jb/YmUILjML2LXOtXZT3qKwnveHj
OO2NP/3jW2Pgq8VAdd2b14YNp0rDMrzfCpB6mcTvIyY6seKFcH34nbAfgobGuRQ3CUi4M6p26mr/
pCqz/5XzqnnBWtGiVjDsyvsqBZl2PXXoJDDmwanEWluZOhsGnp23jsKdUNDFG2sTwDUzf9T4y9mx
rfv4AgicZ+PsBuipMinhME6mjC30jBaaTAmeI3k8y1yD+fcLZL/o3P9X07yCabBV846Qax4ciFo6
UJYgVLdmQbovHOZG8z2OL5dn8oarF4YyqKe10Ag9t3DOV/azrzXdHTNQkpVm7rjp3iJ1uCFY0KYG
3w9h4VDJsD9KYaDFCP/Pi06BgBMORX/YexRrXUP5UA+SZYXlG5UHeYodRjxPf2wYgnerfOo44K/H
QQOTXisBLhVru/w4JZhIGvv7mqyhXOchKSy8UFHeSFE9fDjqs67wjIQlEa3mcKPg6qxHXP9LEGdT
7qhKdAIt/xUMemLSXNr2FdEOOvOnAgFfOnEwfouEvxi2oDQ4VxdwWvkWlmLJASo42WMHxIHc3yDE
mg9r2769pX/zykBfVW0SgJbCMrv+1Djv6KNguCqPIixLxSv3ychaLK3zlomZANBiu67ARALXfgma
VqTSkswJDSyenqCiVDpNcVSAZ0jXqTVLK2AukPgyjgqRSTuJvO0brTHLj8XAa9DhdcUqHoWnFJTU
eFs30VRY489KkyedkP2dYCzRf/49d12T41uGMxos7Z1IeHtF0kZ5jD2nSc7Vw9onbH7YvClo6tSj
4pUnlHul5dJK3yyNsST+9NaQq68Il9FSsJc1fnp0Oy4vco3KnHG2Pwh32yAzewe3lCJBX1zhhULi
nz7moL3juB2mfnO0SNVpXm9h0L2VcUEMWIi0cXY2WzQR4nT8rqhN/NZvv5BtCaThLtofRE4sr3bZ
XzYO5/IQHhNWqnWvAq+axdiuMWPysQftmUTtYfEe2OalJWUgtyGNOUDC2MRDVxeqU1V8u7cESSEG
Z8JP0U1Wbv83jj/VLZ1/DGOPAW9I3qqrMM+8ae7UDuCvlTf5F/Q8b/Z1Ed/NT6qdOaah0RAjLByQ
qpzdHm9eHTo10lk5mBvBG9t1S2k8o2zdNdStM6eAYmC2yxU5Gw/bi07XYO8wQGF6jneCgR2ETAtc
cxzUFkFfsgACrBzo2xDBLro7YHRTfCcZuU8s0MN6rf9su3ptDo0Zv6v5Q1E2nwk5kfaCM2NobtnZ
ZN/OdUH3VocDJD/2N5QRwDMY0HYR6SWnBB679iugdvlROuNnOehuP0WjXqYuYMiGO3vIYwgmNJxN
hukkSecH8qp0wzhOqS8XX23nUxhj07090MQ6DQ0geZ3FQsDMJdLmsy6Qo2yKbyI5utBFk7I3UuXN
HSTsuF22TQY1tzJAy6DhN0++q8t6tGjxcqanne7m2QJWiK/RHSyhzDZGM7SI3uNSsjkAZixHeceZ
aAeuyVx2P8AXzsCbxrXgBY1/O7UNUXMcmiYO2sOvP5Jw+vVBp/co0vwwNWYGWkSazgzwJadaMc3y
QpuhyB6dYnp3Ww5BSDytSsnfCphM/26eNmQmYG5VrgDjqQahCJ0F6x7rykYcUFVoid69gVfXNwVJ
W9xQ2xW/66qmegP/+GSj4mMoN8mn46nfwQdpQCeVkwCHUwFOaC7OaTg9ZcIeaK82knELC9qx65dX
5Kqx8RrZXks7c4yqbxqh7v4XanmDBpSAbNHrqjt+qwlZHRia7gTO65qkIkSBzfCQzEoBKSvHeLim
szlaUcyR6mXhAUnr5eO8zDxFcOiC/0/6Eshw2fg1m/GhLuK+hzXpjQvt9Rn9Tpz6Lx+LITUh2Wkh
HBuCwXhEBJpjO2wmwdgYStIY/ma7iyJrpWrZj1iO+76RPaBHYk75aZJIbj/MfaI5qjhDnbjYxB/O
j+d6FSX9yoOVv5g7soJXGo/+uc3fgZxk/ziMaSjGVGjXJF6zj3P3ih6bPNYTdwGvSD55vhXRCTbg
CMma1k0e73E6JeU3x+6Z1q68GAHW1oe01HcIi7RAtSIca8HdqQl6khRypsS36Zq4gHCXsqCRlk/O
CYMep7BH3lAsCz+q7pbyFEGu1ZyEyUps//2/U2vBumxbg5c+wun8qd6Y5FKTEYVrkXL9kg+98lIc
W0FO+iX7CwXN2W72H36ce3V5GZeBLAY9qnH8kXsPAxprza96kt8F8EPNNKkqWuJY7KEED1gbVyq9
s5qEh21nVNI96iZbzPoM1YZYZcyY+qJlk1n6x9YZ/+QINxFy9UmXSnkp1YwF9xxPbngALskJq13f
+OYJPIo2POIwWyG80W2JSWQJyolNzwoQNZXl6+JHLuWAn4LjiHivFiWhSw8rdxZEvQJWIv8WdJ5P
qcSPpH3ZtMI61Dqby/O9NuE4Hgh0XvzVMMqsx7jPBHQeumPYKW+rDQJXSEhlRwGuz2pGHBzpIoAt
KKq9g9bptmBUt+2TcmBmgm3ceYdqdqMJ2IeeOnZxnzOxn7iSfCx6qj09/N9NdOeLiXc3T9yEOw5S
C+9yCjtNwTpcvRQuLWrg5kNYAEJCHxL1F6mTPsiTSh5GsdourcgXf0EWAXxtaS9kjv9DQhiyR9py
W4O/H1p/amzJEqnNv52N0hinTlcRJ4aq8lk8S3Dj1xys+YZ+PdmEEr2TCjLhxvvtFg/5S6Xl8LIM
xAUkanDXdZmgRivfwzqMiL+p5ga39k6BQ17UcnoOG6PyxK7nxFN2sl3qYvp032SAuydWYqLcQr0b
pZK7OIMnH+QiCBnIFQqQMoNEZcaJB/qJN6rZEkx/FzbnCHFFJ92Ce7ZA7xTLwGAFQzbTW1Qk1aiG
/In/McGFKIwjtZXynt4uI4c2HPoE6zSDQxqZ6wV0X3HNS04N98xkS3OMSRFkpUkaF0yha1XehC+j
1kZGulqLKsACUVUdQZhWf6cGZweThM0HJ+2PdHp2uNJ/+B1NpFM1j8Xsc7cnjt1yPVa7sWFvdgPS
/dymMIO+NmJKKYM+dqwgVUmkpYpsCJC/EdiHS4GvwfF3A4HKCcOmBrm52SjIUipC9MzPj4j9675M
AGGhXochy8okh+fBE94kIp/7lZ+oOy0CdE05nakxgViUbBFPT6RAdw27cOnxitB/BThZY9V3cdG3
/JgNPsqjKbwrY0cEbteovGcgVkurt62ax9MnoerON4vuxLnPvO/yz7on7ho/Zke1RxT7EWNY/o0I
g5ylFaky/VYpj7sKDK7LNxQ7gXzGc1+RAXougU5y6COIzRcty72HeXVHurUsthcdNj8b9DTeWWak
z6MbSnHqnQwZoB9cRlg/heabfCCbXWrsDbqtnjo32SvNVtwTCpupLhpKKjCqD9dHcDO4x9Y0Tgpq
t/QSpOleIyznJ5JhEJtf2e1us87PSAuhiT0DE2q3NQPLKmVCjv+CdWogNiEB8j6C3cJAsHpPY8QH
dGFxjfG20kYFlBJMZhODMjcW41aYEryNq10gyXSqZTUzNRNMPGQb+EX0y4sCjI6MLiPWSVQp71nw
AF/lnIVivdYn008eDvpId6Uabdwf9pjrOJIXSxjQZ0OXSGcqz+vqFO5Hv18fT77CtG0xz4xAKCJf
qJa9X9q1d2fssPpqZDrO57vm1S1d7ftJ0QDSAA57P+d5a0Tp7uNRgGf3kL1fX+vFCXBfogbPUHUf
F97ccOdBW1Kh2y9tOGYYwF7J7y21WUNgT40pVEgPKSR4ihWQD5/HyvgfELer/zIkGjPE1+R3K1O1
OGG53gVhfqHB6ssOL/sR1tEHarkMPzk6nrFIKQsoDqRoqNAiarQITUM+0DdBMalWFUyxcfSvnb6/
zFEubP5tA9NFqy8ngSGfDXkULtqjBPoRKNMdP8nUs2wCyxE0Ywj1uxEQdys1kZYez+n7iLQnyR1G
KmEHwEASOkh1ImxzIurqD7GHJQ+JmS7cCrsxhhXeqDxj1t+LI8N/59sp+nch6wsKiIJHZN/oaHbI
Z7zZyTVmZWlWjhAsUIXPAvPPFGPVeYL1CeB4pWYo5+PciQurWsLYQ79JTrFlldmlgII/kC89Hh1B
1FaILb69trSSaT0hhd+xZ0mzjIu2tukQbT+f/14crnoMoxHK2b9ZAzjEmdATpk3WPI7s12Zz2U85
vrJ0bVEyMGp4SW1opIElnimOzgSOoASPg5N4AltHG7ILN9YKiXmIZqPq+lZ5+1kGF/Uaakz//QT6
NdWNfVW42flesPkt0fvSgiCa/tdN46QO6axpV5OCZUWgrJZhu8qMnWxYyuQh/JHC9NimQNgt6P8b
P+PRDzjcAUlYHuvkkILPhKURqiyCRqre3HWBNJ4yvv22jrIA0czcDqDmpZepuxCLbUi8RbTLxlnk
yWuhYQkeUbshNWNYa6D6Ebjf08G8rhDKAGVrnlb4q542PfV577LQ3InoG8DD545l3Ob5E3aDTO84
X6RwXW+27CaUBqmqAgq0wqWkd0HawnDpoLANMh7Re7eO7p4IiKK8uiQ4q16yMDrFnj4438tqqr58
2XI8EfGh5M3YzPStLOeRTorHpEzEP9ncqfN54X7TyBwIofWu5h/YRBtFUpapi8oRxjNF/3EBU5/C
+Y2D+0J+E5rkMoByblnQb9voKbWoddZDXSW+pv4PbDxaKvA70uTYUVsegz//3Vxv+QbNq8m5MhXm
JbwO1sP1OPDdIsIneWLLQpSrVuqGWAhUIrSLDMiq2ojQYFAG97g4eePBjt3piqXL7nX0Sm0LZc1B
HivcjEFvV4BeBvYmphNop2+FAbJ9yD6uPoLPFbpjnlyrY5TELr55FLUdCBxRmWHhxZyng8w2HqJP
64hK7D+R/1AG59cTkGartlAZIhOgr/spydGk8PJlEX3w4m9TntOG1cWmjV03qviCJ88WcsekZnuQ
4TZIBLytVT0ObU1PLrqQoD/pFsH8bTSQJ5+MXd6ySQJCtMX/7euhl4zjFW7zCpjtNGII28nssTKz
cfPaWhhHpgh/Ebvscg+XYCCTrASYFDeC5RkoNkcv6av52rGFN/kXd8HfPDhOefTHW1y/aqgvtYFu
7yr7pyj59ZgWT1vAQ6209DWp3HrudwZDnKX83ZRwEOV5vQYbobF9M7r6X6iol86ogUt205aFA/Fo
McXFBUF+wKTyzXgV5kNqikw6cjVBLezMTGjaoMeq9U/TFaLsNWIOYPeYiksgnaHBABzkIfBgJJrO
e9nrtsYBzvIiEtfizDrMxMFtmxC1yZEkWfWhDPFmaxt5jkTUc8hBArhp43oerHmsQFq2NO+JL8ZJ
gSAXoG6/NZr0aUZ3iguB70kI4FJ+6BtQIIv+2tFrUvzphhbu0yzSI98UjuErkHBf8TLC/7frtXM1
awglM7j7TxIRFefkqs40ZMYnF6Pa0cMZu2kBGaGqPEt/ihuLRmx52fAMavr5/qyxgea57A4i4Pkk
emwE9xzECgQ/SHUZcDFbYs6CrRrQxNIfeAHwbA6bi4T4WEooln22XY1n9ZkjhW/fpTsjFMyFJ0e8
uiBIQWK3jmVU0Oyqot2uiSy4Gh+m7PiJdGYl1OdFmAPdMibLesaj3x30dWJy/gCcBr7KVSXsi+9B
MX30w4amIJYoly5axPXcku1fP0sLO5OGOEYThR9ItdTpEInuaZqIY5bzVp9L9zOURJIBixQNpvEB
S/6x9vA9XR7oYOMCWA8EKhuiPiD21OqCFcvvAsuNMVz6aO/by6CLyP92QM9vaz41rLm5fc897klw
vdaqubuCfsaR4fFR6+8ShvurK64MpMCEh/W1TUWGWUmvARzsECjZ5zYagXAUufrhiUdvA+ev63ta
K71yo6g84vDhCmwgNdkSAqokZUl/3TJupeA4Fsrg29/8Ar04lt1nHnL6Nn7L4mglDWiKj18+5LN7
UZVBvjOjspbNnh8MaKyq8TEotcPbSZL4ijSv4CND2NmOfQi+VPDCzAtnbKuTQBgaRD8/2Cg9nloO
yTMs/e0X4MqcWzaULLcBn6MG4zOXa7FcCyZezrBRyxgAq6tLUTWCsPSs+ul6eX0xXAN6CQy04aU4
stAPDhNiD0TYwzz2Hfu6yMTvy2we9+WP8I21K/Z+iFR7PHsiSRkUpgrKeVY7F4gw0BUItI+RZDol
mW1q/i9JzY+uzR7a+5PRAW3DGqw+Ss8CyrKGkBGJHcgo+E3F5DATNXnEcIqH/sIC9oTxlkCCD49t
hdnVTbOVaWdXlq4+8RLEpH7ETUPJTxQlmOQw40moMMyGO6SmLA7+p/Jvy1/nfR6fPzgsXBFYsymo
aHz9pznJYVnQpnfSBpkwtFR5s+Wd3EOu0t6NSgTtqQrM8QisJyRFTqr8Nvl9BkhpMju4mECJNUAB
+HaOKwdnXUXB1bQ4zjpfJ8kYJ1rVGQDFBbOCqVnRfai+HAiY7cZIqdI2LW+vCyjNN646CZHe6q1A
NTkbvzW4MxAQW9KnL8ezmeZZlL7PUsnVjLer01huCt6gnNbSp8aITiuNrpluceun8wA52B5yveid
KAK2Ge65WqMwCPGPhDGlj9Jl1SewSmDwraB2y1HJyRQ03ULSJeDwRdZVwJ8i0OvYeh+iiwnUG6pR
48iS5DzEy6cJb73tFuVM/Dp3PyiwXEY5Ux+YoAMruIslqCXp7V+jQR2Em6O/5dZ80LqEOzRC79h2
ytCkI+S2CqawPhe/8XakaMK8HQCPumR7S9eMnBWKrmA/eI0dIgjQQ7GG+opsKiZqpQjMMAJuZc7w
idNUcpL9pavL00MiD9w+aME7LbyK7+OKi/pqVOiXsXECQKC78tRhgRy03vYOnQw2aJUBVT8KRziY
p47uk6R4dU+oAgj35H49UkRomdBwyz1MIfu7BXFyHktW/xenCpro9Sw7VWi+ywx1W5pzgnQRJ1jc
iVJEglofNsOh4S+7aakVlYXCRmLQqS5uoKsTDabr/a6XaVgMDIBItbAXEIlxhT8oLdpL0paMt9wp
RZvoA+srDPDnBGFl5lBk+p4U6ToNOAku5zAhlC5PF2kFGrdH99WGb1hiC2WwPvLpU1F+bBOPtjQs
N9AuopYDwalyymVG1H7UXOzorFyZtyLbUs86l3uXcMHoy6w0cIxhc4SuGfr55FIzTtjwYNX47zxV
VxoivFkQ7kPX8F0nIts6wg6DV+nC08VoDIMrZ9vWDKu1Y16MefkbvaBE6MRQ/qllGxRqOYpGrQGL
7Nrf0cdosYyoXCoKyUYMBnNjZwYEZ8bBAOCIOUe9kMWjA3DD1MGe/uh+rLofPGZlG+6Vh7EJQuDn
6uqBve4u8SHKGwY0i6ZHyL17T/HX61NI4t4+NAHaeFQ3O3p59AuJzP6JSwX7uGRwGWQW9QItOH1R
+FCdKW8U+KOQuLxP/vH/yJmyx+i7BmAtgEffZb1SPqKydJZwQ8d7bT79ll3f4K87JRxFHknGvW7n
z2s46k/huXAR4fMYNwDpDEZvgdvOWxhWMPTYkmURU5bsSiqYbva+jPUuwCqbxrtxziu4JilUYivF
dFHhKlaI01YIXPBx8VyV2EwOQsdIyC29oEEC+qYLtfiiIPWEHBeE/n13Vor9g2jEAic4aGA25vTF
oqFGoAgnJyTFIv/78oFM2CkFfcQWucyOozwnHxQrNuXVWwdDQV10xtOPa6p6aos9yYMfLnE2FILU
6LR1yE0N1HT2NqqTnOcKt15xrDMDjy9v9Ls882ObdIs5K1D2N62KZJbfu/qiuQs+FxkgjU5tSRXd
X4Vp6YFyGR1rZHCyO0G1xvzdGp/Tifg6YD/7lALHEsMLEyW7cTqOshjOPsqS0GxmzL05ME6cG3EF
R8fzroNHTEInzaJDqY8/HOi+cJtx/gslixP3jG691vqGjCyp6TkgBl947nAo4QpfjXIPVoiynVNm
zLfR+kyZJ0PhKJ7MouBsjaBYQcWuAXH6fbNlt0YWf9umiKBqtVKqedYE/NL7+b4s3GQ+1ISQkApn
vdRt0LbKXKDYZa4nD0i/NBHm90fORoWEVSyUyMZNXmQ/2P6+evsTEkt6bkiHh1dTZI/AVjC9bVTg
jt7QqP3OyD3CZknMEtX2MgcxAI0zwxMMezTKxq5uC+xYSGwSRRzxpZwx5p7pt7LG7SBUzDlqyNjg
Iu5SNAmgYJkm6b6HgrIC1itXnKG0eL/Mbjvb9S6uZVkOg4ZcaInA3L8IvOYw4Hxl9mgmtc6OMslU
EGhl3E/j6lbJLpK/ineenS1lj+f/gPCQWKLzWzslYFQxNZRG8vyz+LxBlSe2R/CLlqyeQzuxI/0c
w+UXKvt0t1TO2oFCPhjr5Xh/lUURMfqDA5d/yFv9AA+9MnKx12ByB0XrU0k6b+suQkhPBODkT8Py
ZQVBBvAGb2uY82BzG9ZG5YVOYnR+acb1hR0vhN/FrkAT7c5tA6l4+Zi0+wpTyt1ALpBbhdeRLzFq
D7+WsaRbl3N/IWQQS7UDXkE8rS50VqdISl/6LKQq2oogAmnTzQOJgfCTT7s9uku1pmEBCBdMbrW/
pbI49DrgJDnHxUZZgrGxoCUNjzo/19rMU3Dp+Tz4fUOB2q2HruzaPI+Uo5yPnKMcWCl+clTJD58Z
yYsx2lco1nzuzo+DGjkHgrvSlL3UTq3+QruLakOpy+IaduPe/UI5ZSZAfYb9sgZlNf0JN5B7LR/u
cwcEkApQf8zE5iA8D/PQ+PhvFRZCUmc8MCkWHBsnQGFESCBpRo+SQgzaXYCOrbOlejTYI744i8M9
gKjEtWdJTGU/k/w7QGs1gWOjKcDcMNrRIBX9pP8hCwc6ltfre8FsKyPqQFUdzzRUyWY8Q4XWl58O
GYYQV+EFC5fTcKDtqfcMbebsf3Kw7hmK7xbEZjuKhnNQI43JqT017iA1jK16WtqM+y+5G92vIsfy
7tYwL7f2fPRXQfPiawv5d/BuC1A4V0NZLvu9snxlAdKKwhAFCCJYP05D0Np1ZKPPtUWoiVn0yqBc
KvDTg2J50gxec7c1ADDGQRs4X8JsTzBin4K4f0DG4xKtwqxAGLZctXa5K1JK5P7FcjduBZQeaxpW
2ikU+GR6/CFpYncC3GGswXbXFmpAJm+JpanWLyJWztHUyHCeQSbgNOutMIVDC5O6tcJb1CpsO0pX
pHwVtyI66Pkn/vkBcWGel4umn9G5OxWjaOFiq9RtrkXBDI7ut97Ln7YahMKhQ2IQovweA+GW/HB2
zXRI1Hjz0y2VOYoCmPKyXOgDRZAMkYmRc8XctkkL55Bs7HUG6Ieg14STVvxYaDc3iTsgu/GZWSj6
UVRZTx7w9xsDGtG7sFajlHDMnVefJ7tI1wJMujDw1SUs/JWN+fqBkFJIRob0dIaNbNRH5gH6AxDv
3T7DPHDiTrd7Oc+sYt4K3NmcEIAJdUUBfzoiRZmEd9ZD6HrbG6ipwYWqkNwCVDSi662GMjZ/WQVR
MPf3q4MVeJkzcuaPzhMlilT3XWXcG0D9HpCYcmM4MY4OmZC/lB64XxhvuP1BqdYwvXXLfflPtA/L
1rjfV6Y7K9yPuZhubex3vG02wSScZUlZawAx1G+jdMrmw2H1ZpQkdZbOqoELGU7I8hYS4MDzFfIU
E0UYTMzxqK+ekuTiQ5+thjMe6Fjoyput7pcQtLK+B/Brr82nAkBPAjIE8MiGUqd+6a1/ije7sWlT
yRQ25aX/BrskmQSCYD5Q/APxM6nzmpToK3EtAyQh3ThoURkDngWBrEVO0E3l8ewNhBQmMIi4gcJA
Zn/B75x3wC+TIkkyljzhxOQNJJb03syupXKY15GCHCWwGvqXLlESJWVk/xe6dupYArE/J5DVrP1C
RsN2r2dJtKb0/plbaeQs6WqLE0rlR6lQ9d+ARWVvAOIv7mzAzSDDEuWxGnw1Xx9w/LDzCxSZkovf
hUeYQ4U/e5KMsOQVwNtXK0d+ZJtsyLJKiG3Xn+DjZA5g3mDidowtRwBYIHjJOr2vCKFgg5YB2SWR
gMzXWEn7+L8j1LYE3MYOIRc4rkeY1mo+qWFmMP0fv7rW7r8p3DXZ1TqxgnoJy/eqpQhbC1/z8QWH
yoZEj3LIpGMg4liwO2btekN26c2QKOr4vj3SnGVSwJd8EXk+jQjYLaoo9VSgb/2O0ue2E3CP9zag
N3uGeZ42hAxQ7sTsGMFnysmq8vlbr3ETrNt1ch3032eRa2+hNnPlmssYbDeGHTX5SUrbhDTkjA90
OfWohStw3dqOLgDoYOULvG5tfHdUhYZqiY1bd7SWGK7wjbXgwgOvpGQHV2Ca4bSI1pJw/qT5jpBP
sgB5vjXYtzVcNXRt05gkTpxh60JB0CSkXtB6S5AB52ygCjjXaVD1fD582DNY1Qf0WxXL6ru06pQg
5uMU+j5cBfG3xPD76RW9lZx2H1c/KDcRvCVUxh/sqfpcV9ESeISrAO6edZ+PBgVaz/h+lJBXNvpS
Rzb8nOmynCptxM78UlnV6sTkqq2OfZcsVwVWGj0vQWZc2qLsVA8n/cZSRs0bZ/zUCTHy4Bd7lDOM
Nx2A8BwtNekjoMfTD/3uWYdmEz86Sa8LoKOvPDh4/I58grvbKZEv58/6MqrxNT687bGqbN9QYIj2
xJfuJ3tkKqDbQT55jmaG3ed2PLHbnlnZnGW7QQKhfAd9DKEiLtOooHIFEhMTPbhRITdmTvstB9/t
L3h3BpzpTLZ5uwY217iatclJ/SaSlA/olJkdgLsh+KY1dMcKpMEz0NQh1NKr2ZPRxF5/1fW1KP9M
5XQ1n5tGn+JFZGvy+YuCFoZVb+WzhKWblD2aAzgtTa3/aTxA2EZEQQEm1LUQiC7J28P6e9LM4Cpx
2g0NGu+NFzIuiphDyR+0XT2EYAq0RLXvKbYRc8E1IBOZ7H5WqtwYRzxD7d6w5qn+hFI/AZwA0VFG
n9AWIJPrB9MGj1jxpBybGZL+/nqJiKuJw8eNd+u8QRczmZPbWzAqk/CANHs5h+sCWUOmTmIYtH8g
9OAnao23EiA4kbjKaeJo5t5CGLliVE1a70ayGlPqxDOC/Rem3OZP7RYbLV1obptHfsizFISjPWJ8
ue1SPjIq3UHKEzhZxVHfKaonxY+53iysgjJhSm+l8hPUceKB7ijJKwro5VGjOvOOUZuBe1c17Baq
82D8uROFGpeg0nxJLLwUyCmPm38MGe2AW0pc48r6ldHT4nGbXpRxUkB5uIkKC+N5ep1clYGS+S9G
1S3up0Od7qjqUjJdLhoRO+pXpaIUEYX0JMDQvvuu3VFEjhgilJCclehSztb4JNJy76tx2j9NnYrU
sM43Or1uxNh3n/3q4y+3gVGYLznOkq+IAEWrGBkLGCAoG0VilhlNCDnLYGn/sATmiwe+utX1+4sn
ZJGckesaE5tB9SgGV10Vqu3mz255C5mnatnqa6Iw9hEYs8qH4tj0OminEzPl5NtgqWfxsPICPEmo
cUJ4i/LAH5P12I3j/SW8MDhvpVvs1hsve2PLKt4kSz0YpUgIul18601ZnWrnv8xlcOV8jSrtORLA
t+AgQ6sTYtnbnxDzV34cUexuJ6Qnb+ntSRzmMm6Knxsf77yv7ArETBcGBdz6YoO/szEM1qW/gflB
Fz1WZjZ5WFMi0kBHLR248EDYm3i4DYQsh40W0RTC/YgZWckFatpNAT6KOGfbxEiAdj/GQezlCUEH
Bd/8ySv0/eGIQZvGq0UOA3ELLO8y8vIWD1suJ2PcVyYlEDIlsq0IaCfRLt6r0aTPj4ytKh0V4CSO
mJStgplUNWjkmCMm2MsoGsKXApZObfFLBSKRTeCKDVNjyVsfOYkxuo0Ob02RW7dyWZxqtrAqq9GN
J/w+AdA5ldoCbUjY/pnyBsceZOM/W1Oi3B/b9Hu+nUY0xTL9ABxOYPHWTbRY5a7pMr6qpaxANZZr
uMVRa4+u9xxLzheLb1OjPaI5e2ZM7/2zObaU/dSC9Rktq3YkSN3vy1TtwvnOz6F6uqQmhkEuLg2+
cTF/y0cEQ1NmqSf0GwvqX5oRH4powhPoDg19juYlB9yLCRvXAEjU8l2i7jfE48tf3U++SLbll0j3
/qMh4ppz5j7RMl1rb1TtVv7M6f+hHdiQUOUvxhjNxCwPH3nY3L2cZGMgBmLpqcadvYGQOe1GZdSg
xhQc1d7p9plgRO8QC6H+FJBU3x72iyC7G/sHZuGMNsP/IUUiYwujsUpIW8TOjmVuK/+tRLr4k16S
8R0KH8W1rL0V5V9tjTDRMMqbivSpSAj2xnNCf8kki55pVOojZ79rYbt+tPNZCZpgJ5qnh7W3JyKo
SkNJ/zN+nr820eclujXvHL1YjppNrW0C+OQfGlhxFA2vYHlXIf1TQF8nvsz+JIIvUaOqcU9hNqW4
iaIIGhv3rvU4NgVJ+GYfPMzvRxhuQFcV0eewZlHKAAxyVmZNQKAANAfeBcR35ipdwCdbGlLljK/B
c/xF5qSA2OgQejzGoE81e/5VTVzj4mi84NpKfez0FyCaXDsoXypHLZQ/6Mt6U7yBNWgQVoJzuMY0
jE2Nde7d4oWVNSaRf/cPnblmQSIWQkBUA6bXt+Ga0OqUL81izf4gB7wR4G1GAuA/hl1X13jUoiDD
nnZovz7Fd/IwazJtpg6ByarRNfNqFBWYMbdE87K0QPk6wb+KgZtkUepl7S/rW3Dwojay15g1L5vQ
69G97P/sF0Qy5Y7QYnWlLUUxV6OfVg5IlWcaDh3RI7INV61hJ331Vm+Vnk6CS88qHTOoezJfrC/y
MC6CPGPN0enfW4cG27H0CSXaGm6G1RcDrTq7o7QE0dDbFuCbD/558pBgEFucGQYx2aWcn4w3EnLo
3Gh3106VRjBmSEnnteUkbcFc/VDD92YQ81Lmkgx7qJAqnfIQnawcPNJm+ocRKCE/U71HpFsf0w7w
pPJUrEcI4WOGqWGR4F74uzdvyHYmCCRrEgtmAjqiPHvmKXeLOUK/rJ68DZFtTCuWNIo+R7nDPkEI
xZpyyWJSes2ANzCndLPkQmJb/eTpq/DZCtNzX429aa42tdvJ79MXATnSYuS7F+4VVHIlG+7p5Aux
TkKvXG+RpDuqLCWPrZ3Y2n/v2d4OTSRMIyXVURvq+GEtVNKKDwU3UTyNPnMt8obt5QP6QrRqqf2D
hNGCc2VhJDvJKIO4Mx5+21Yz+7VMF0gHHvu8UDAAYzVpLqb0HlD/tKuiI5x+gCHhXPwuG3IdqmED
YPPfz66TtIapTmHFn0C7dxOyE80XZpID3HhJU6pZywSIEsMi2E6gSocgdeCMPWGoKjYEcxu2BU3u
KKUyY2YmSa33TOmCBIWyy6CcpsCgMb9qdEO0Vf6HiWZkRUuH+imNn11evJTGf4HlUEZGFCMZJJog
rRUMj+8s62mQb0NIVZoThrWb42U64A3dmKA0wrEpiCTM1xF1VYTMfiPPSboqwhxbkVx7sd6ITyuE
/+QowP5Fi6rRIqRuJZhenI3BmZwlLLHxZTZ3OHNI7jEPm5g+ix6PGEgW7tD3QrXDCsWtR8Uoan9u
lJqp18J52vSo+ouBjEkZtkarx9TsQtucP36OXHiZlXtUO0t6N+8eLWChp7aRR9nbzTJ4H0tBtrxy
EbFbkdqXxO1FW/nIIANslCc1oCVqrq/PkiAQcdTIGuHXZGi7NZVDYNiKIEqoTeb2DTTI9DMPN7fv
OseLNwi4PzJolC0UgPYv2i2xYHA2pkAYGJiFArG+eyVgY+18QETWFROqZqfBqpObb/J4PlAqQLsK
uG3xDWP6sjUFmakazAG9FCv/v5ZGPPlF0EUATqb2ntPw+uCquOZ62+5/7P5ziIkiRSatt6xsc1gW
ouyqL4Kk1a+eqOkWMXsHrLnmaj60vFYSepxYNU6zXYz7w0mvNfgD3Ts/idtPbC7wEfuhYkez1Mib
46qc8QhI5Z7V8Y1+9b4qla7IhSKRqMuB7BjXTojn3NcFrwmoc/C/1lXKVyi0gKMkE7mJ+waNdUvb
noLYSnLx2LT5rVi0gcJ+xu8vUqx9mPmRZa7k/pQhLUD62sK1QYN6On/tjH1fpoQOL4sdInVe9xA3
2QMU8iV+HHcD++lOm3MFiuNUnQbLq+WzRqf484cdqJFRU6wiYbFFATak+DEoSrF8IbZWQhjUG8Cw
kL60f1HjIYndz8Hc85B3skJ91MK9pG8S32veq2K3b26F8f1rH9PPlaEbuWJG3z6lDBK+Q1XpmWQN
Wa3W2ojoTFp0LTzvYlXZKVQMVv3rIl47YUEb9tnvZbrbSVSTSD1ZH8AumYDuT6ZnAA+5mQkwOgF0
pynSEljHrVtNtf50FJdTeANZ4DFTbxNI2368SHyn/hsf0bThrMchnRLOR2kWhLFuayWTtJdJjrd9
TsjVbblZmqZ7PWGVys4o8pHcmWhd7VaIIias2KSB5U4QUl62eggUxX7YJBm2Hy621dRog2eoEAKt
/8DHwLHsUGW+7rQH2X4GHJhc1zGK0dGVdpqvX37QjR3wdr1sP9ow9qR2cUkONEmt7GnXPVJg2VAz
F7jr+kstp2tb2qDnjt8ODSLRwSJyVvD76nnUoY0ahcP9a3DlL5rHAYo1Ff7jpi5PfhJzpYEnNdGT
vAQldYn8p2TxA/xeht5UfhdYywbGTMvMoHNTVfsVx7YSD7OBkQiLjT2eSLSA8CTofT2m1eHlPS9y
xLW+lxHVQTu33i6uWrMdjhqnfIyNHyuJSTlvm8UAhSKghQMA/kIhwoWncSPz5/AYiYecJLU318Wa
Z447V96coC6/1GYcI3T50o4qjplkkJ2MYT5yo+ObcXFs+tHFgISpnnruFh3HC688Ct7CVrWymxUU
zf03aU1IHEsI1lV+W9aS2ezqHqgQExi3zUo5SjI0kVsYs7CglEInq5vSdiX8HLFDCzo80q1qorCm
9RdHe9+o+ZTinTXoI8mUuJ8VR43o0iunFWFuegegfGxMkBaahAUyKoA9yXipXr+ZBeLCE5db/XkL
fFEUCIhcLILt5f/70FtalLq5FIQz/XPsrVGu79ONltQHCJkoGPbybVVsay4o8fvUQXjvLqohmn1Z
v6RHoD5sl5pAQDHQ43sgItnd47o2IU1N+Vnm3sDbJtmKPDH793kPkGDqfFuR8MRH/lejWcp4vWNY
/C+eCMxv1kRzG9HwBNDhdSI7dJzAr/N4EGdgaY5bZQOwmgyGON8wMAC6zPyGDB5sMe/YUuQ/OBWo
8shCC/mJGDwitvFd8IqxGiDm700oeufVxq80Jtrrm0OwDJOy+sEHg4w0+y+OZxUm0Sp+HdczcIkw
XBx3M1bb1FlXsu0dVUoYLRmt7ZtGHwmWN2xwaNYHs8iK+SYHFI+hhZsbbeeHPZuPYJRzkUIoDKgf
mfz+9BxkqbiicvEEK4uZEm13sbda/v7ZkYOrR/k8V3yQEOXTvh22PRo4kPVNL88GBfmDz1gGRH4y
Tjkj3wV6qyCniJwOX0W8KiJ0wbKibO22XLiB/IGMS9nnQtBQxQgPb6yrABy2FAFzlLOzRdi1v5VR
clp8W9s2Tw2CssBtt9oZzw1ziJCyXrFgCny/i2WDDaQSo58kfIp9odDancxDeaJyCM9UyLg8yfaS
d2J4H6zMSQcj6AWNCUJ8nu713EVLzX1p3Jgu8u8XXF+CqCrC5J1WTAXzGTJ3YKksziTQr/es3Bgh
7h+57kkM9U75Iy2I78eiiRQ0WuTTLbPZl2SBByJ+kLd5LyQKrnDoxcZQ4gh+T5Ua+w4MQjo1Z2ZK
w7fH3r4j5YiDDr7FBsg4yVqER03Q4SNWW2DbhGJqeRq2DqD6LFkJDqkCM1aqjRIU9EAjAA1wLWeJ
wB5kG63iAshmseaIzpFyuidZCI5CqcA89d31rFEKVffgzshDZ1cmeR/oR/BoP6dkQtHuP6GpzA+m
dBHAVjmBXjeoNBRDAx1q1VS3RfOHohXn4GM5bKNWGSS9rEvFFqZE4KL4zcdz6OC6yJgIb6cxMRuL
zJ41bKTH1smml1iFZvcaDpCzHLjBNtJl2CxtduLp4ODBCrKJjjBLhlmve/9twyPP6UxqiAKo1Ndt
yX97yVwhKvXGoTtaU4x9ETOYsr1mYOt9PCkWvYDe1KwjUDftqJJBVtfO11IbigZkqPbzT9b09R2h
8U25iLRMrVeVq/fDznk0DEqGOqmPgnGDcUdtmF3qvSn+22kRSxJtw4k39JI7XU6btbEp/qPpqnzC
EQxtTHOnSgxfQFE25FHx/7VgHMdaqPqy5MK+CFZP2zwe+M4ABLRz2gWNV++p6NRE2Nf7CHbqadX/
rfKgjAM6ZtwpYC8iCyI3ekQ/RyJVy8SCDrE42Dra3v4ct39Es3LvTwZHGbQEsaWRGa9lGOhYy1rq
pf58YJUBfoBdacZKBKF8Y61PvFhulIJWUYy/BnsK2GF+CniKNM/0JhtFLIcFgnWCkz84lc7/vUqA
AHjlZdWOHoWvGbPfppsVkGc9jFS63MjYyKaF4i5lp3ZnXIuKOcvddSBYyvY3Si59cIXxQ9bx0dx9
aksvDUtB0lcFtkvzP9TUU3Mx32cyMzMIkv9F4/GOIgKnbcNeKJa1TKpU22n5QX90ECQscsbIln8W
ibZ9B7OJqaIjnlRBSVg8nQjKJSPmhDwn2of90kIo8uJAhzsAeRGyP8/o97qGafp+ZUVMCAx7FRpv
M9oRHBgQ2PYnGzVKwafe5G9ynzqmK1THjgYxVWeIKyqg30JLzEk6KSjk8F4Efy19k4v0Rpj1vpnH
32ppidEh+Z3C48yJHKMBLxF0MQUU2zR72AXETl8lIrynoC/C/Tu79e4ULg94SXEsQ9MWwz0EqiGK
VXj1CBnAx31BDQqy66lCI/UT9nmPPQn5ryRhnPQ6Z648IFqQZh0ckNVTkgp6wU/sfdShIr3iwswC
ylfDPkIEQwUQx4F0tdJNQuuO4xiN09Tq3NBKmAcHnjTrvDfDrf1s8hbgrdLj4YuIamyoxOF7nIsG
XYeX/cYhoEHZnY091jjP+TiKoavynKIhG0UteMcNLxe8CI7Tj0Yx/or3qQz1bXDsKGx/CJCRIbCH
dsl2PagCA/9sWhWCq8oY+AF1vRquLmh+WhEV0cgPeMnGf3fmU+tIQJ+NGyRaPEpYo9sQPuZq0BBQ
cn4IeVDqtYaboQd8qZ0+PNfrP1GkZTkjPrgU7kN7S+VdXy6CAIFfy7UmZ3lLzXB2CLcIvIqG09A/
+sPnnqPqd/204HUx8pwPLbLrFyTHM20H8PZsJmPAoB+7My7q3XyEe4HjC35sXLFHWYzuD2HgzRnb
OgucdT1a0visRtkZMN0LQgFPk+h5pT00EN9om2VlZINPNP5xt3/XL+2vcvAVNYVtz4hr41EgYMA7
xHFRJ+V9QMpuKdAQkBpmt+4wRiOmZMIYKWWXo8jo89cXDptcjPKSJb2V/1I9ZKOCInEKvUwY5+K2
P5rnH4YM1dl2YJV1JfRgZpePy8oRwdtdjqlydS+HLGvavm3ZUiCy/3WQFBa+OjV9Vdugjl31iNok
VAlgvDW1hWEgvsVztTAVQMBV29d5qcFzQyr0Izlua8DaW04IpoLWD1r7JMY9XZcAd5nif5Y9+a8F
JtRuhG0zbjj/Hq4m+DPPjKxCHR8mo/mE3+vsHhBvBFc1dVOL3s3dN79BNTl/nxG66z5cr7Wijehq
ESSr0Y+Fa+PJs4KuMQaTl2bca6C2uj4aULPm/wS7ufbXInkUYG1MSpgFJsfOjaw5f2zrPrHeZsLa
DqvF+DE3WBvu51B3flwuWNwEaR3ad1fKvCKI3LT3rWIhoTuwJIL44d9SlAzvq2PY1vQzRaZaHH9W
XoC0ExoRQxrpjESUY81F4EEFXLjAftrZVDP4d4GxAbmbGB1a1MNDpRLNnyGmy4QIoPpU//BxzSsd
DLgQScAQkuDYCD7+Z3J4n67fa6Ozy1FatPaIa0IPUOylcaTQNmAnOj5MJnZHJMB5ILTui0HALvu/
M3OpXvYPBdBqUOCDaawsPfOtwZQrKhjfzeOlwOtEpA33XCjKs3HVLsGurRWwqJzdtp3oNhfMzE+7
kisMFThxXV0bctMqUeSq6UzTX4NPwiaKLnJG6HZfgTD51XQDMiVSEf4oj8YbiS+4uEOC0GlPru3F
NKrm2WrZMCdJGEW1txhUSJnrY9p9NYxyBwkbabsobYTkloksBd1w/I+8lx+ep/F8fqQiMSi9evgi
k3ZdOOL7coFmO3jZxkNSLHM62wkZsua1rTMKgngQH/twS+1/QiYuWIbm3uaTWBXWGHRsdskq45Lr
w/Jb1UmPCY7nMCs8QnItbjL0KmSR5fV+jOlbx8CDIv6/1pKl1+rUHynMcptXKqGgBPnQVViXa+Le
ae+VeCw5y1qZDZYCLZEusT8vG6DHAyJ4+E/Y/tS+XMEMecAUngbbbyS0R2U1S9QxJD/yffV6gtJH
9+/QfJ+9nvaZeZruIC8GBViCxxH4S105Xws/aucF54e4mZiNq3b7G/zuXcskCVOojUqvX6rxbPdf
y5RWhfypmjjoiZ+PlEIXSr/5Zxir1tUqTjFBLBnteGPjBAv5nAFgb/5rrFe2SKGFfrZjfdmIBtnN
nuthZQ2bvmSVKFAv+x2EylarYtCc7MqivQ5FBrY6CVC3bgkpKy+f1ieirSwVQ7sVhoNgMss9bF1G
ojj+EX3FnDgrBVKmQwR4Qs+tSYw3jILXoKeUCi4FjyJJmdbsRpI+Zn4g5+YSny/xU/I5MuiWHuYM
Dmw7IepXWNRk9ezPAwxvXISYS4VwkF7/t03a+IZxszgrj2GwOrrisXR4tDW17MAFszhIaS1tBwfn
I6JKgbP8P+Kuv42rRZ/26gM+FTWRkhIug57R3yQHYwT03STQ5f9hJupqJDhASVgAE64JaiVkwuof
raYtEexxIZ6uvFD6c0XP6KWefMSSaAWZ0tEp+uDmbj8f1ZgoO1+h/eP3IhlJp4s02drlumdetwdk
G1YFUC/hLjn2DW1MEJ4V4nC9mY7/+kTrynHjOGEg5fHHH+yt7YtgfmUX9+lmPXsHUkN5RaN9M9Q+
gsJq8Ot1S2RS0tC6VA5bbDouvgRhXvzWNB+XWaPWEWeleP6sA0dTgQVOEY4dwR9hWbyX3Ou5ibx0
RCFZCibmtM0ay7f/wfa9rsLMQP+micKc+oKNUZVPT9PHCFPHBTl6hnIc8RK1RDnn4s7D+rYc//ln
GvMp8fWLqAGOgT0krHxND9m3qH6JGUtwj/DnlL4wk2m9ywNvyd/D7JJZ7G72Bl1blo5z3sxbUTxf
BPMDOfkJzmk2VIV/4mly0vrj3gfRXzXUdAHe87wM09+bf0AY14VyqD/exJoAv/bNml3IIXadca/h
D+m48ENJ52zU2VPpIcawOGo60kGUEvZqVQPPqUflV10QdVCsgFd4omVxv7ovLAmsBxhqjQgbQgV9
5exZmDD4vEZ5UTGW4fyTmcdr2iLlA6v7JpmIkelRtRCG1xkTwTh5iH3hAeXHdoUhBrsYIE18BiHH
rAMxZgmtxk1cjgrcbiAusSZ7JcpbPiZ4ADGFWYcCeewJyryaA1PuHpSivWIrBJnOIh3SCpXtOEr6
sw2FAQSGc1FGMt00gG8Y8fy63Ab3Z+ywdO8VtffICqevRo8iaT6uykrRv1C6vvoZDTf2lMedK23s
h/Y+qL1FBCSo/T/F2BrdPeNBH+8quluUw3eM8tOQHNRIcYhWjlkU410V/oHf/IY9IXs+Osrb8zx0
/tzWacyi7Ln9PDQ7JDfjvLtWB5y+ycDru2TCutePPrFTL6UwS5VSFEJcN9/7nZ2DAfl7RS43PjfW
JIfocxyCxcUmtYUwmTAiitBWKYFaJvZoF4s30ENW6739V/1JwW2OJPHAgGWPLCFe7VDTCapGatPZ
s365yPsGhjuA5wjO081mLIcj4UaabOPUVVq6b1TrtvcWMtrv+mBmvI2hoCKc6VuZL1iL0v96HCxg
12nwxayVmM8i1cnGqah60JITQQuwVny82CwltNFH+hcpGevaZCraZrb6LvJGGcFDUaWGzxKGY6kr
KpGBg10nEGDaGw4RPsWQNPr1b1k3JLXVnqCV+BoK+sCpLDEeZyOtXrNnStZ28lHnTNHRvWGbL7fh
AvXSt8M+Jej2NiZMY0OAJYYyIKBUREBn4sRSx1eSNyZMfdiMCe0qgkAtZF+LAMBOUyraJ+YY7Zrn
s73jEvsBZK8vgh5l/oFjnaDQnhO+OVzHSJq6RBcSLTZL2XvGKLs80RUAFSnPWXhqch81gG7m4LkT
vC69bwAxw6l1SeeGMiwVni+DGm2FcW3KfQyJcHZRKec/KHGDjOiBolvb0REEmpEkxhyaf5i06Pey
nF6mL2OgcqN1A4JsXVDPQBg9GDKrNZOtT0vKw5eWBGYpfKzMq3ZHLnlq9bWFkCo0lDi5BpbioWeg
5M274Fca77XHoXLjBtoUJk+81tpADR3euxoBdF9qUkwal8Pwiu5RhcVLn7bby0Bc0YEle7mYbU+1
9hPzgp4OQhzgPpdqlFKv3sDbdxg2Q+rg5KzgEbulOEYF2ukcdUtlhKAk39+SOeJY0Cpyuxce2MG4
W6dEItrazDBjtowLYOlHalf/8Kfd6EASLExuBusY/3YURAUmXGOg6i5FCLONN/tsSODdahbmXoM9
pHhOKD1q6vvmdRAgs0Z2ApLU72WvZ2YLHN7gdjnV1M4CvqJQU0bSNi5AAkcumjYryj/Fph5OYMEy
tYBocgJkWx9xDjmiUutEKd1VdQyJabSWSH9+tk5i8G4Z5hTpBMyQSxzM3NGqsDrjSI2Xq/8rdve0
9vLaERrWDkcMdL8BM6aLIIsABaNILACZt6hMohNZDOZL/dNTTeqzenhmbH00I5SVb7VIlI8uPpM6
a9gNt/isBa0ITLsqLYAdOvdU9YVH0OhOdIYm1/lhyn88yqaVC5yZkuhrDyIiP6LmsWLTYKeSXlSm
/qCyBsTDrpqTsU5cGM4xKLomfWn8jeUmTehV0i0qAopnutp/UtEYKWXirUOZNm2jBdFqMoD+smiA
XH+66VpwLuPGBGPyoooAZKhwNZ8LkZ9gpBKRHmp6kGg7fatEsAgiuONPoHcJkXSpQt7EIYdSZXYV
qDuvuTZo3X66PvcbT1UmGpv10lsQrTXLMKY2p5JqLXDigRtUUmFw0Bafxr6kZkgO2chtbD1NgSN4
9ujJe6+EnAWH8rDIVSfc4OWHo1KUzBlBhuJwLIt+VDo4W4n1Du9T+rA74jDojJVmKDybYOBrEUPd
AMOdSMu7wAoZn6bfzWnsu/TCCsTxJoWINUHzc3yMp0cgcaLPtsesOWhv+oWe99HXigYdKmtxO1q4
nvqYr+/xH44Ktf5EO7Qk9ZFMZ8+lstEDG7ERuNmQ+d0GwVXx7YUSv6pGR5y3YlVrmYnADyChXkKb
FMuVEMyoDF2547PkT+yOlEwuAcSls+KjmCF55Y0XqYQ3lOTVUuwHkYo6YGKuWGfhkQeSILe3pH3o
4dc5af8OKrTLaNgePnCvzfyEPhoYgkTNHPbHAVkUNEbg9P9fEqOhYY1HfZiEKtPmKVOLaOM831Rq
L8ispN0rfXttUZgsQa0GGrElxLi1tD9LXDFCsbO8/nYcV4JcwQCxs3AYD39oNCKFWHvWg0r38x8U
RepSOxUQ8fVV9BHG2sgvXlL5G0kGHCjJVbc89NAr4r9uLS0obFOvkVsMSQ9AGC0pDI8nABJPYiUH
6QiGDPgXTbzvtKy8M0n7zukXcJYAGVoYjwqqwauqxw8T1FXvN5kOH/LHcn1lQ1FjJqqAblPcttfD
LUo6dYoX+HQP3Hj0DOO6Ocu68SCY169pfHAFfEg/bholZyuDO2X/HlFXfRRwn9wXk4K3BQzo/hvG
8INOSeWNNlOJyOXXQ8VPulOrrewInZNt9i64HkaaROj45G3CS9gh/n+hUm3WYehBrY09cYeB3AWO
TCF9ArsClvKPD2EDEvEuPijRNNsChS11d+YoE5ptHmJg90Bbt+FmoHpIVHfNEr84ffCDcklN8l5P
U7/6DHk9bEt+1FxHRsYv/wbEDDom9GTDyV2BL4VYxMFCnzsxTOSdx7mdgIXLi2attbGOPUTX4iXf
NdeiJWoBo7iBU42zur3mSEBJ5R1nlXx9l0PjvmAKUR7lJcwMHJFj4L0rHCOjYlAQkfqLAW2GMLB6
llkqumMkcfnJd3ZXj05AnVRUWEfcqtlUIChPcJajepoartCPWbZhgcWy7g04wHOiyg4Pkqv4baKh
KCEBzc18GiTOYfeYjZchoDbnsuxfboLjcqJTA8zjP6TKjePrLQNBiLU4OztuQ7FjKDz57UR2sF7H
kzObteWxB0GdD7RSFzuTbI8oobIfvLJh/L0RWILwbHTw5u4rWzpqSIJgxYMYRoBx+85cRUGQQXKL
+G6Uad/aEy4j1ZzTtJoJn7UlUpGBmWl9nGiAJqo6C2T3koy3pgWh0YnAKSz5855MpWQnV4WcuoOj
+qWBH/KShOohYQG/9Tv0agRlbpVQviILrmghbD5+yMslmPmcM7cTvQOqVVemvWAysXdzpBd5h/oL
U0sOBPXhyP0kEUx/LEEQNQSq0XrHSRFTa8VIkg/HD8Ckwo1IgX5d0WT82lqy0lIbiJfJq+KfjWhk
mGOkM1TAcMtJ0OQXntRMdegLQNgqT02SJfQN4ER9R7kvgJ8h5L1B/Naeb2SFxNOftZExXXYMPZ/+
L7pshgeyJm4nDXxMEft5WoI+Mc7o/m7qwW98F8NK/ObhUEThEMyd970yQKFBhU06GJQantEmbf2o
aSSpDrNrKzGzJdDKtbdBWj7lpuS5Zve9dCjZPM2DQ0K6DO3y/jSDYQb6JOQVmy55esTz+6tOtV4V
/ny9pnLE60WqlD24G+v4EOyKn+X+4JEXVlcNtUCUOH3f6Cm5pJTu9q3QdyubkIP8yF8uoI1nkcCN
LCqZpN5zMHtdhaiceaFkIqm+da4Bts8XDt/wW0nawBe9aShNdZ/I6juqu3FqihV8GvyLjtvqs/W1
oCo3u2q8kAM26pQInAZCQ9NCVibY1/C3kiseyiOh3DKDutfCPUwISU9Z8Ccow7NCY8rQCOrxz9vf
KiZUyO7kPnlAk1I+tjCnzaEWSTrah3VMDMq+Cbx5zlgCYRYtOtmQhkSDa6NBR3jlO18KErsNxBZh
mhmVgiZmYYAFAWjpaGISXzOe3ghXkt2vJMIltHTTqD5pvtvUcZbFhp5Rp2qSZ5oEMbtOXjlV+Kz0
n6MlcYx/IY/WBBu03aXRZC8GR8KSsux3iXxX6gIgtgo2Se8E+wPHoU2JJCYB7nkmpv9scyFYbcIG
llOrC+H3jbzzrWpQDtuOnG5yWyOwfCaeLBjrGYL3ihb4P96LdYZJS729NAKfEdffLZxa4MGIu5hP
9loyPuidrGA09PosiopC2ZYFG44M31D/HHpYb2aBticfOPn616LxUO1GWXUIkdH1vfCSNGsb1nNh
v01ShQxfcO4/xjiw3zud2FW5qcQnjXwfAb17JB/lKOcC3AmGKxs3z9JW8UTAjx4J8gVlvYEIZLCq
tyHxvJc2hrFlCaszJxgKNawJXRYGWb6ZSxsRFkzDQMXvPE2Hki7Mtrq5davC+Q4LuudeyErYGXnR
TYcpHHRtHtvRNvr1/NqViByJNX9ulmiLiY+4NldzELKyJy4O5NaSpP7hCWBKqASoyzrMpJGqBUsH
f9wtZu3WiOWB8aVSRIKx/NMqH2bPOop3fBZS48gsM4jhbhbMahJ2retTerroshYeaoJlWc8LeJ8B
4sRcIftHmjkSttl/xQm0pdeHfzVVoBZq9HMsOn4RtIjX7Nr+vqwIiPFF91xBPVPx9hudsiXf0Y4D
Xafh48tEH5KRoCBK8PFN5dmjqWmEfHf5rbyPCYlctYN5dSXzCjavLX0AAXuidG6lsPjX8aZYYdkH
dwzG+sUv5y1fSnzuLRtUkAiK8yR/uMSkAKJEjfSQAsl/fN7/MbGvIK+g8IE3KEwhWLkvO8u829gf
PLlWi/kqZbPXblXmfjBfVj+y4qMPkl+YpRufTU5FQ8TL5UqL4bEVFMglajTI6t7IEOvFPdpNxZgY
InCTgO+VU++pW+G9JQE5vQ0BtqdqshY6J3YB1pfMCGHTD0cNEH9yTgX0e1SkfSREagwH1IzqI0O7
JwtW97aKpudllDyNQn7lyTd0WCPB2AK24E/K14vQ8MgIuMPwTgeXOQLYC37cPcEhhjqWU1YfkgRg
33sijHlhqeobgvbcwIrKb9x6VHyCa6Cga2pxLxCFZ0Zbdqbt6qmwaWsa9/loO9ArU4blUvioS66L
G2lGKPR/wUv+dfhXkFVjvGYObZ4E8A7pmy4pnzky5wVZAGCA6s+wYRPv4k6W9VE/5PFOQwC/TAxy
SWcC/assKLBlM+Ao14EcEl2+1Q9EFo0TFxo6iYC5RQjKdAmA1jPcdUTxx6CN9K70jF7I4goFB+eZ
049l7ZQIC09URwBYu5tBBEvlstSj7iqFTLdzIkUzm6ucBh9yrDmG8ptRU7XUHq993WMnu2cHmswn
0/O4KWMNNapdEeSYT/+EBt0j3DaKNzZ5WPu+bO3Co3GB8K6EuqaEIOvh8MTTSj7v2JADODEDrUxO
/CVULAMGuC7d63Bz5ZJFFWjx/Xa9eWTQuKw8eGVLb75ruCfvQE+6JUFzwaF14pLHNfQNbMOCAd7r
nVVARMWBbAbHNhh6D+iTYr1bEfpSVct6wHb+JhtosHmKI4P1GH+fUEWZLTeFJaipjh/CRvt1xMFa
1qalf2KfdGueuXBGTdYzwsGPnOqD9T3+74p6wQVFwqa/cKQzfIsoLrcatcwLlINJaS2BnPQo4Gi2
/TAH2hYGMGuNqLfnGFrIIaJ9uAx764tGkSqGIP95pF9X99BnPRao873xwF8kus9drzUdOmfiFZni
+61RI4OY9AX+qPFYD+EgVtbkQ+rYd4owY+AsXBxJBfuWVxyDzGJcPMB+2i5kMGZdsXb0jKbgFvaa
GFVWk9SdOtMxi4tTbjLR2zMzx5YbsDuiXnp3T6iIouMS/f5AD7ypHt7AyTIlK6czZjgkSjoMadYf
n/pMgg9q+SBRcuN1atadru3tH1aBYYLKSC5KlmuiDT7HdM6nzRF5aHe9xNF5NwRdWK/WJ7GPnlmm
ijdl/wUbQbtob/xkSR+6FcZzaJLUglKWSOX+s4P8dL/SX80QyqExMIAgZL4LEPzGZXexzRZfwFnO
3lCu/Sw/BS+4TIJ0zBrtQJmIup+L9o+c3KXgGpseN4+Xp3EBb2v6iLSVbTvzf/68uNHxpTk4G+Y6
yH2baWWkS+j6/ehBX+xnDeD0MWT37RvrBPjK3ZrnMx6SJrtfZ0ATHgXBSQd48EU/JzlYgNHntIeU
0XTGMdiaBgVpCCQcEZ+DX9ldOhB0HEOuPnEexN98l5dUpj7m6jCSoBW65pWYrj+w6JbHEetMdLoU
z8c14MrrmMdP/4Eb99C4/A+0bOvNm//PG22VJz1V8E4PoQNaD8ZSe6qWH42hwoL18KubJ0vSQgb1
3sCmTCJIcN0eAcz4rKOpKEC8hXCV75dOPu2Asd+Jl0yXDpt3LsZkYJPa32Shj/Vzqea7pFRqaASm
VtKJYbSG4SD8qjsN6tg8x+xCtPCW5XdmFyLs3YsILhq4eXPSbNp1YfM4iMqoERwzHBPyCx1kC8Sz
mULhhQqv0e3J9S2wf/QF4t6rTxrDpdobeywMCVxrmIMYbHMgF7vCxzwsmzT1TtH2RXgTdq3W0VJ5
P9NZXUvnatzekpnyW1sRC+uX00/MDhYvLVxTYAdDtQl2ychS2Bth3Zio1BBgkHIIKHP/gnAHS31N
UQjo8Uj4qgtOqwfrAKgh3ruxx+sMAU8t4Pw0R1wW0jV7LLyXBaYkf3gtlLUHTxAZs7yNYG5G5AVS
1AXIfh8VICNRUqhjsBEVq2QJk4hG3avk73BbJDWHf0Q1gHuWLr8U7eaEtKHFyywS6GSQaEKUGoOD
I4ihrktFa3AJPfbnbrTrxd6zYa6Fo+KK13a1QPk2hw4dUVpRHzNyMAyQ2wlMIz9gB5qgxtnKoE24
H5tqyfywwuXyhlLIlRTVPqAhykfFtSI63w1PPESHnRY77x9awVCyCL+uacPNNoGmVHb2/2/RzqRh
q1CRnMHi5qNZEU2ZaUBQwjU6fLgizhHQ5XZwYYr5YvcYoITqwtCSPKQb3JG/yq1F2uukSHOkui7X
pSF9DxhGgxIMKO+BBAprk9UfAj9aS7RXdrp6cNspef+LUeeQfBEitgoowtm1sprLvKOZ1I0vIfBQ
zp+vOCCZhOmca5xFJQ9XAnY5r1N7sb4L9BS6pzr91S+Lw4SYAaXtvHOLmc8BjVSGnNKJvpmBF9sm
wZ6eHaxBKcPjYM0M+P4ghxU++w0xeHBzkcn2pbXARcw6BTaotK4lhzixyzLV4k6835VC2ETUygFX
CjFRJpPVSWCxe5X3Nt+B93UlrJ45/Kwq75HzrGtL1qhmybWZJHIuTmcs1hv2d8/lBba0HmoS3WZx
mwQSo0jzLE+G04BaYKcRHuhgVkvCEOA5jvzdGMaj0va+O7Ip2PCaAHd+60RnGGStalg2lITCoEF1
PBD8S2PAuK/xc7W4D2bX4r0mpyrhh7PH4dv2Yhv+vyxacvIqmSZLvR+lcZayEjR8eizWkgVwAmZL
rv6PGG8BMwJ6Room57F2SoJ2NjPdoNRA5+8TEBNrDPv2f8vstDageP6ya1hl3VquEi8YqkKGndyY
nB/gX/S8XWtL73B8svb9cTVZeFjYQF/a0i2vWOl0Os0373pKRnmXnNOdEcQt1Hf/4tX9q8fIg9cg
y6l+0FUK3mVH8u78r5Buv+7Hcl/OXOAHMCGJlZINlvyN8BQfUOOguzuhO5749rfc3X6T/yV7nZ/x
5wpjciwMCcAO0GZisqywkgT3GpVQaT6bjgOQPDek5ws21VetrKchxbwtcWT/Vyo9wLoEBwhrOUYF
xtggyBOYZmbkc7F209Nr5LiojXKkkrRZxVW/zpmzZveR2UmsJDin/k2kwVdHaNsGqxtq/QB/67JA
oEaKX0KR9Ox3vLvIEvwXQWMKTmbdcNH/hMtdsTuEYrSV3Df0fAZ1w53/8foXTVAUaCdJg7CmxRNE
QdC+7KoPvYUGIygRJwEsU2YWkgVNR/4yiDG58CBKt5qWUpYdpbIDWh8jvGfbL7B9uHb81aQgQ9w6
e5fll+pfbFhgD7LfFz73y48xcQfkLTKL3W9gEeU48sx7CWBuMKyDOUB1owLapWczKWOL5heiqHzo
2f1xCMuYyXsgKk/cYvKBqISPzYzZhr6+0xmXkD4UDY1RMRorwYd/iyWRpSKYWVDr1bGybFoZCDhk
sB0L6G/T6Mq+5RGukw9Gs6itrtxkU2ObjTMNvsx85ep7z9sQ68I580eZgbJZgG+rCyP9u+9ST9Ht
2aVXpGoe9fKy4jJMY6NxuOm/8zKWlnYsiMNNna8+kwsSKffqw/WGRZ2xyUgQgfbVsrx/lqXpkkT7
JmB1PknklFzLN6OlrBZU07DF9De6906qjFsGhcpYlJtpRa/pv8rvO2nEHa3n+O/RZ57Hq1SW8MIL
B0TBtFRsgKKkFfTf6vpFPBxEF9PokS5ciQQ5OyyUqmm1DWSOPzQRK18wFludpYMRAhn2J0t22vcG
cEvtnUsHqm1gzv/Z6M1gpZiaebskc3GfXVdJm2DuW4qK1cOG4PTgLj2vxRiY3GgeL/0RIYqW3Sx8
KomcR8tj+DmgrMoZs8bN7exhgP5rYW9hAYBh0ENNpLXpm+pZxPqAMuwJZ6xKt0rmxhoTCImNV9RV
cQQPi4W80EQqX/JYi17H2ccdg/1NTxIuJO/yQ+SIFz9eNzJWtX2EhOszmz2K2jYL4DRd09IAznAR
uF5DADWmQhwHTupwq1+WOX8wF0uprajmMoILTwoKFCnuelUG65h3p7DLc62W+h3JngnFOVWkgU2m
rtc+WYvPd77vjpW1rMAM1w3xVNnCI2qYMOOTuVFIAgmWzclGWjNNIRNrlhy2bXYqtI7lefTTrbgJ
BinVY+g7o9s/MvWTkaYzhcg3cjMO9LwPX+v5BzhktFT16bZbglu9i66q/9823N8ouXW4AhTKw9dd
cQZ5QCmBqX2OthuKNB4BzhzdPuqQ4A36qysGDB6mCvvL8ebNdCSUVuxoISGZbPD6bEwXpqRUbVub
UuKsnggcaFx2gjOKhfhU9ee8AdZN/nhuQaNXrIANnIO7F5km6Vrf1hvedkZAh/jXUo+jy5X2nvD6
TMeM1LDme0SCbj0FxEfnJj0+czxtUne2FXoeuvixcxrljRl1xm4RWalfwnOMif0a4EiHzf4P8Nqc
mKjPrkkPxJYH1C8MInw6aAKzemRc2Gwvu+B5g+xfc+u1OG9yrr4wo7Sq4ZGxeDm0gybPq9hg5UwL
EcAx44LQgyUmO+NMpi2bbwsVDdAx2DkVVygp/YTujul1Z/aDohQk8l837jCYqWVqgsIjS+DmbcA8
v/jiTWtjABrlE5oOPC0XuvdyqxgfaPKTMKxDJKWFbz05l1hbb0LrgJNmV6O0ythJKjsnwzqQgNFQ
tS2fP2YdEfEyxfekSl37+y7TSn4AAL7TZTqkkUNsJvtAD1UFNUj1YSuoh7i6JmNXRS7vs0cmH+lD
0JH6lCEUcDWTtwp632bfJOO2Vs9o4lo1+3ak2pqzzo4XxoOFz9Kd3nJsYpGzh6iY2p0nuD/fS8DE
G5NFPVoQ+deNsQn9f+WLZFDvD4D8m/bmcWyEL/QzmDb+VXRVrnlF5k/WPq3GxcLJATw37iPhupO4
Km2Uso0ZFknURm7DZjVNZIUBGAsDMY+VIb2H3l8k0lwMQTtSyIwX5mOjZSRiM/BjUI0bAcFX69ih
XyuuQ3HE+okJCpcU0dSg98f2Xkw58IS+D2qCH8yg0Y1+Wx56k5HSOsSZ6+NfHNTe6hkWsst/xKXf
/F8xfILRkiOnJqK3QZSqLoyBzQjTj1K6b9z+yXTlkjCJwQLEfUzOcClPgvcotkwC/abJUP2cVtY3
LOvG8n0QKzF8tSlQJR/Ix2Ep+BXZRFe+SzbQUiF8dNAhg2kUl5jTnBycJ6txVhMG9RD8A7uR2CC3
3VKf9fm6vGatYR5C9cI2QWPjUnz1bSzGDVquXEOIo2fTjaGqmBtdDm2WMj1VUBq9jMFAYMilX+b5
xoAqQbRbDdo56OGej++qSlajt9//gplypLNuFn8sLDkF6QTlTyYQ11GYdPjfpADhZwG6H7Ffk2yD
nRlpNRyhOr6NmuVQ4FhFopnDjPO5rjBWPl5MxpuQ7h9CNvRe4Infy0mR0bS8AyUPBOvG9S1TnwLb
dPefLlN8H04/GAHjxylOooHOLAx62Y67WqQIC0N/zYuJsyb5KgKHUXfkqiiotzICpTUZKJLIjdEA
A6/Qd3Vsgpm/GO61uQcqQAy8skTKCV8YbAOAPZQMnjVAGyEYrqH440Cmhkd32z083Tpzt0jmQ5ka
ddUtee7zXc4lv4ajxC0QmQuhf/Sf5wrfV5AhTtS0BjolQ2D9U5dvtyQX/2hEEFkMeIdxNuYm4XR2
VCNmhHgf2/xWknn58mhdf9QqJcJtW1sURzvfCLiG+yWhQbmH8WhMSL2W8EuVII9WF4ggt4+gihEs
Ey/UxlbCKYapoqqKSh5EnxeIf4/Z47XNsP+eYGe4K8fuesk/DFOtyJTkOvClZ0CsBs03SsCeeEv4
fO1S8nCe5LyhLBeYS+qoIZnqurGoP0GX684A+Veo6M/cUob13PgBLKM3JIMudRNaUtJHTrgZWboD
PFak1say50ap6PwHJBbTq+yG9rvIANBYGhIaaHzI7utb5j+n6Y8L02MucVuNxbr2dTiEy/KuShRF
uBGpkULUNCNUbEACYpvEA3v0ZfeENkUMWxIT3a9P+yg6knGCuWj3bGlmDmzE98lbekPAbjyvOnRM
V4xnns1cUoxTIoNJm06/tf9SQagZSTqFktGDeoc0UIzpkc1UIslUJImTFQTBVpe5ydnN1lFQUZtU
tOGyZUhETRLQvXQyL9hjTlBFeIWGiwZZ4jlaoTbYqmxRMsmIRAxuZTgiuTRcFUuIRKZDX70bNvpS
mNsSGiLnXu/GGmsxSwISoCm/qxFP7XssDE44XG7ltJDVhkzHdnZPWrY6bh9+enMpeLZZ9//eoM+F
C4ToSNEActipLtQF9r7CjCsQv/5B76QIYDRCYhR5JUbLjalgCOwaO0G/4VnA+WdMFbbeWz13vAt2
OBgHmGJ/h+ocixYzaXALY+idZdjEGydy89WsmEITPnrPHN20z7KdFxs7YzGITfpntlR4GAaNwfux
kpjHPdgjqOAxYSRQ3DSN3exLvlbW5+FVvm/kUntj8CUA0F6i19eABz4gYlkCFhy7BAZxCFMKcTyx
aWjQO7zOiXwx/QGNl6WSlX9Jps5ejK0Hevmv4drSN9FqLqcEVVDKdyHigMr3ab700R0s8vIdX7U0
hHI6iHE9TNwXtNS0nQsQlrU19cYY6S8/hpNAmJgT5o8N2+QFBTBID1gnPkXPHOmVCk2MavPWl4Ww
r0o8EokTlymzlemre2VgIzcVpfcXxIio15hBVR1uo67KVPMOPhIIrDWQE+qqHld6WeyMScdLR2gI
obzjjPQgW63c13Lfc987
`pragma protect end_protected
