// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:55 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
QHiKt1+lTAtfj3Hsoej06381+fYOm6935aH4B8PLRsrzsU+1TBhGiW/M1eZEfe9v
5itlO1JYSFF64DH7iW8vmSMl/n0g/d/4E5wUYhPK27TlvtnYLa2V/CJpf9KZWr77
Pe5qEA7XxnnJ23R4+94LuV1479GkZhBNYiWfN59iiFE=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 21408)
pdJvdZgsnBO9K4TiBWDSfxuS5G2r73bb5YsNZ8uM+CoLZc41o6riyyvwe8eAS54M
VmUXgFEKyr2ZIzElWhh3VdNz3xZURGHlKdfTWyDeKLczNFZ07dF+h1NBOMBiDbRZ
czZbvMUTEuJWssHibIKNfpF2LxEumIZiiBMEfPmYT1HsZMrVkZGIw7+YQWydiyfn
18kLMfSyexVQHGfLPf2C76uMzcV/BkWfUeqHSZ6QAqjTTvsJwFBOwJG1RTZc44LG
vf1/3dAkKfEf+lrdxQiX746QtQMRyUJwwp1UlEcHKAyk1pB+0qBxhzZTJqZhe+KT
M2iqv9iFuas+AHTj0AcYMBAl7WT82nU4guuzDCbxTDUQlcBX5abSgA660IFDVNdc
N1lhYnuZgk3RGlGFd6heol/MpaegahpTk2aKXzxb/CLHvdLCdmyeagE8zMrt/oTP
AcqZttwcGSLBk3+FdyGgner9vzR7SXiv4swaXdAosoSijwdPKb4kM+M8W0fLMQEE
sU4zOfIyrD34WdH6yzPB3vKRvSfOTp6CX63sHL+ecvADC5Xus+af13ba9wPt4MCl
v5rK5zkpdja5BxGQepKTmqqunxhZwngZqgtnBZS7ab5l1nbmJx6GnpQVihzxJGkn
X4sRzl30FaJuMx2ql94UkMMz7fUe3UbYnrxJfOCih166EkcRSm3nGn9qIaQQL5cp
d9/IuPEPeXz8ddMbfJVFIjfmcEJNmFZbgIztUCQmJVXBijPVL+yy89BCr2yocGrw
RDOPcbPvMVwgaGlGhnEYP0YvAI3t4P5spYnRcn4WZdVL7ZkTqsl+zRgRPrlAPvpU
RBOrCNVJs8As5kTUe+SZkBeDOILOFoab008fov96e09bgOF07+jCS1XUd8qH3FLV
HsxxFtm0SlLnzWn5uTn+zcdv4qSaiuM4vIuHMKcd9MkJzwPJbt+jtlOCsYAe2USD
+TtwxGoW6gbVXZk3R7/l++FdG4eefme7thIYBQGPibUcgi0W1vG8Y9/MgqCZCl01
+GY2/gi1hNkFj661gPG1CsYzYkWuwBnJENXJdOzPgXUEHePm2ubVAwuNArRbHa0N
tAfHCqCQkg7yVtziJTDfZp5XlvWUruuveNBZe+OK6xbvayElRRQTdoH1zKi2wlTn
akvcFiVnfP1wekMLg2zFPaQz8Z/Qw27w/fR6UKmWiy7M0gKwNE4FzNpzVW7dp95g
DGWExbQdgomOJlU+JKIJysxRvvizOyIhKwHmktTV5XFKilkOEMKCjBL/AqPxf+lw
7GQAmaOXuD+DNhhi0FadZa7Si6MkDtzG87jyH5YdTzP9Pc8MmLgIQ2sTz11yzwc5
DPPbKZPOjVPdb4bx+YbxBzWvF3qa+KhXaECqsv8kh4lc7uQXHRa7Lt7tojvezl87
vPnppedZewyaE6uM7Dl0A+GriINdmTY6y65B1qDS8oy/WOZbDAlnkCEJaC8mgbF3
/fKgSvLtSsBhTTNY2a6j6tiy79zumRuSFZyTdjBLjxr9r2pEr06gkPI4y5OlR/Ns
PuMDmdbcnX4AJEy7X1JyIrr/cZSeqx6K3wMJFWkCIHRu4+nuXpYw4nwgRKSCLB2B
iltkUvXllAmOQY/tTW1NSHi+S8FPHT+RbDXWluzNeBM8YSu7B1MK/tcki0HWM1WW
7a1SLW9JoqB7wZIiprFpOhhApPAiJKwyW4TTLzkWSf3cSYVK0NXO1ISoJI4vfheO
43nfkCXpPPyeHVN5z+osV1B59Z6W8ll01viQqOi8Bt93G0nj9qXtjFE60L++05Ju
PIuxSVPnOxJicKWk+ht+mO3aISZrYLFJtFQpcao1B2MBZCsXOTziBDPJC3SBanQM
wJJEyWz2V1ebe5nuFVxf5uTzdlNMU8lN6kbWPXN5ublSqF8Ev/LpEgD5wzULjKqF
yMCnj7j0QsN8+ktpE2d5jhw4I51pbs462QVddOd/ir//SWeaMITb+NA1tF7lmzWH
JSp6x5Oku1sefyORbXt5r2B9GLXTgBu0zlbhvYwhB0l3mJXcd47PziWVlyAIzwJt
ii3JBhCrvNjqDmQL3UxaqzXYqhkOIU8dUJuiiEZOE/k5WrsEiSuKZZ3lsRt5sTIL
ESfWYGySZXOUHV3HKvLJb+0Rgv/thQTA7Mbs/z1cA8dx+BEy0tIVZTDj+Wq+LGpN
Y+ywr3R1ZjF9UwcgqXkfU5oW/BjGXMo0IgzQ0C5V2p9EmxMczaBirmROiUgVhCxP
vGpJEwDs5Ox04B/cJo5v+5hxl6YN5eF8tegRP+TBont+K7s/+vElUA9j4TLnVmBF
3zSm9OkU/q1TsI8jrQ0kpWOcJzg9wW0meqSFIUFppxDnTTZVLEq4GlX2XCvPbYTF
a6ylX2S1YYjZEvt3acuKc2rkxaBM47wsmCQ/i9ABpQwnVG+1DB+rBu/tl4Zc4LNX
drCKJVi6WM1zSHQjlSQ9YGjkOC8uLKpNOAJMFj29du79EyZ9qSPP3EC7NVED/378
HWJP8hMZ7OgXyj57VwJgfGBNBvrPnoR2Segitq0gMvU7EY6/jq9/5Yu5d7tDKhtM
VpFnIjXEm6Opk/S+acq0M77xgrorqYrDr8DA5xXbha6Nq7S6nGWFfkJsoGUsvCBr
B7m+dnuwRMR14uOy1RmxUaAQHUpXYSePbV8mYyM+O/1EFAnEQ1ayeaW8BpUIIgN6
3LMVP+Ckovs0Mgjehy9f1JFoLKTVrORQhma+RFGWXLIbsbS3XKs07wAMl9Vprt0D
UJNHMK4y3gFLh1c+mC4dwamF0vpes3fpRbG3PZQlsYZwotPqVhTJiA76RNOrUfZm
8W9Mkr23KPHH651XQm11qVG6a07oFK3xuOVE3AfuloE6ag1yYkja5zeWbJQtr+7k
gaNwavHJqCHKeOuXULDX3gSdpe6rDAWdr3vOQNXOajbQNrROTQzFlxqfEP2zxNXj
pXeXMsWffAfEVTBsnbvvbbrUz7glGZ7JyDLKBhOlnnnTD6JgP9oXcW2QKsMXbfa4
QYAL87ApADMpZO0GxKKYSwdwsxZJ1lQD0UHSsP/DEh1Yre390Yy4g9FHUr48JFli
pNVogLQqudtpq+x+UtCyIViCICYQp1YzpGvDlcDDG6U15G8Gm6r3KWTaFa4rtymT
Z7eLrlTQtBBS0Gn4EtDNQai5dcz7s6sIgATJCJkwre+A62XFE3l76aftij8RJXcP
w2dvCoAlSn1Pg90K8jaq6ZmPK2WxsjwTx75h4TK+6VWHlultiYtZxYOiKG9OGNAF
VVgrQvqh1ld0sPNtOq1n7gt3wRZ4YWIdnsNd1jM+iUcMP7VMVs4zrMnHodKF/MYe
+7SO7FaGsm6MP6K817xoc3Ot632/RQzYTvRY4dmh2p0pB+I7Gg68OlCuTq8FxV0G
YECLNNwAOVnJ/GXLnDG86toSgoiVC40rWAifr5N3iBlt8UMDnd0lflKDzvpsp2sx
If21tXrvbCLCr83xVIxktX/yqbeLUhmC6galSPQAGLzxMHaKU6YIHKTCgN+aepJB
yj3mZ+TMBEA5uUJizxGuF9XdMSHtdlUxE2+aVyxXVCC7g5VQ1puv1JBibHlgPIZo
OqaxuALsT4o4hWDc7SZubsAjHkQQuhmjK+PONiFvLsBtCKn5U0pwqCc+WW5oNTrc
8ENBHPaW9hbP4WP3q9OcEdSIx/mastOmUhfexjPQ0BQQJDYA6PcrVXWt101KMpqF
OMNGSt2MTL69QRNY6k7DIvvuaXHZWeVeJvTA2NzA7ClxeM4QB0ZTcmxA4FX8OTLM
DwzpUJpOe9+RUAy4WpKZUcR/shkpGjKkNqlsO7lv477+V2ge8B9E7bCTcpal4dJg
Houc5Tvx7sPJI4qEPezLteD+FTbGLr0+n4YXxZw9FcTqRBk56Buiug0iRXYrpZz5
V1zAx3O30k3k6Yw5ESg8DeUpiYdLI5o2GRfT9NHVb3o20DNg1DM4dejdDPoX3fUj
z2t8/CTGuWJ/Ld976xUOLdjOED+SaOUMKCrGVj/mROttp1jd/WyYmwn30ll1UM47
9dLOoCW9aIoH08euY72H3/MCnrr/yCksHqHeey4Jeww1ZrdIwEME/I8tbdmjdtMn
cdRF/u8FjDjqFOGr/kKFX9KKsy5N3HzJU1nnloOwvJUy3kkO0tfQ5LNUTSQMPFsS
O4b0Dyw0xpWTZyF8i3UMeRTa466jVg8orhMEENuWDEe8NZ1mVTJz1WEe1OSS5Ldd
W1gKGLuLdPPuGpMHWUmoRkQSl5eDTSxiZLVdF2cbPoDYqyGRQ3rzpynsH2MW3cOX
QSOXB9hlMLjofJiWisYvfVOyYHU84teFWvYV5IGjWWp4n//J/xXJ5IaWkGAFgZQe
N+AvRCFDPNuc/fan/DyKolzqs+y+JRTVELXuluWotn0Rzj3o/oY3LW811Ry/Tpdm
3xFN4KhL6d83Hk6QbKKdUBZpmuUmYDNzSLbO2U+aCm5e6rjpGRw6fgyqtb+0XSZz
aKSuy+UOwJ7/StJ2qlP2f222nR92l3Tijym/vVaaOfysq216hm6R+k2mICrlPqN6
CdfRe0cqZa0yenYkdl5khpe5FIyxcWyW81DBFYBqLEdLNwnJfxOMRzgg59lFQh4h
goNsktOD5NCpr1AsH5s0Fng5BXiUtU5QKZz5l1JUfDkfCpx0rEkQMYXGuj8K8yii
fFMwOfc/gqWbrwlIYy8I9W45KgZoMUCghL1QM5x3tOwVwCZyv/2oSOtIbkQXxwEi
jFgbwHPK07tTn5O58E1qYb34ZKbym+gbPiXlElFf/8mLeUm9dLfUrWn+Ui2ofIhY
+DK+sL/UTx3q/E83xn8mmwNAniCgOKML+tUsPbr6P3Fxjj0zhlpLCnaL7scB6Wkj
P5iKLhC1Zz8oM3JJGsnMLyq2i+4JjtwyidqzUnuGFFue5plFPGdTi6CqY+v1KHxa
qyCXxLkFSVPzjRKLo1FUjmO52dCJGLrwieW3juKwr7xjrLGJu0mEV8eZ8NTW+zHx
vK+q9nJ7hy77+lQt1Uuztlne3uoOfCH5nl1V2pm3rlEtNiPpzOq6eqLR6f1x4Wqq
jekW1tOMJn4exqcEwRdPOpKD48LelYDXW4GtrHPHaGSeGNz0aa7Gmh18gy3b5nwE
ONJ8g+p/cUBEBj/1mMzFNaEsnkOCxT/DdGks1SEBRWfbr5Z1u1746+v+om48gMkW
iSs5d6fktFU9p0kUamZk7Is4oK/qIvfPM5BWQqNO1DTRPv7MltgdaLazgEFRBxD/
YYf0Kbu9Va63CrJ6yC+jibOW5EhlscJGxTflcuVlwoafJaD3tJ8Mo0UHGHK3DGso
PIsP4jfmwS/lQfVp5fhrsf7tUjseZpV3b7S25kc+0Hv9J5KOXXMFfeis+pBAoDND
djMTeMLTdBkRfK6JC6Qi00kVxfJpBg9coW05xq+adcoeVhcxpTj2cWE6+wNIBfh/
2q4FhPfCyyL7TP579rTLPLrFSQY0nppUtVXRFuO/iS+LGy4YTpuGgrfAB5U8Ha4a
exdy8s9z8h/pwCjx4vmN+IEnJz72bejDQ79hkI/E3X7A68AQYr+DCgIuni+jfWbn
2j2xrNPjikiGgnYyEZC/uc/s0WUXsgg1U5AzVnOtYvd+KGxkyNNhxG1lVcHV1uDu
CK6qfdCq3VPAgopyceB1hbJUdMvBMQLyFRlpxEtZlYcc/CC7jaQgVsEzzj9Bkvtp
ZYAKD6w1diqojoSDbqIepEDgn9KhXD6aVQKyR1LYTIgb4YVdOnwYWgtpFKioFHu7
3JqKgYRqTnQVPzrcXDKL/aM+oWvMBo6gAHD4UhYT3XJCBe1cshev1d3Ws/Y9SQ7g
/N6SZedfN8RSy9F0lQMOj4VGnwYiJndHW6QRdEhf3iP+k8Fz09Zz/CkhIjHWQVMh
PzVaZO//v+wf8KOiaSVDGY9dWH4144AplB+18RqimF+LtDhqTkxHuGSuW24Br+t7
AIbNMQDpYOWvkOURwNrANmknrk9N+zH1fdfVGUozvWQXUAXjDj0DqY2vvGeRaMUi
NzuMeszhQQVAlnstq3c7X/iFF6cpMKsss91RhS4XTTGg+yxPabISQPvRAovGQ7+M
/+vf+87XVQAOOsEsyMiuK6yPu2l3lUjXV5uzDhtooMqH1nBin3MMlx4zwq1jao3y
wJqOgtB1Xl6sWhUN7MlvIuQBa1astQ4NJpTl2TYreSdZB/fgrf81xktxnMuW9off
KSzpusMXKLvvyVP5pTib/6qbIxyfa7T5nRDwTZjd8YUy5XFKFHaxrhd38wwTquj5
Ovs3w0TuGdHqt9pgSoKybrQZ2p7LwBvRrBHkN7gbZ+40q5Rva0FoS8xHG0iHodD7
qh+g0/l+00CNoHFY8OQjpVNPn8F4oMtVCq+qovCto5/jo5mcs5JBc+i35i2DjgVa
o202x3tcGAPy0i3ofC5Ssv9VvBFbuqHFYtzSkiiOEKxseKyuwEsG+ydgPodtX8eG
N7Mc2TXyuglx5d37B90qbc61XghP3JgwRoK6Pbd/g4zXBZ4Hajg0+JboUg4SsxYN
F9IxVip+tT2Stu8cwwtErO6JD2QXEtGgTvW3jqXAAerF7zneFj+0EPOV67pn+YVV
iGpX/TW24g1xLBJ1VKJ8B3YuwepyKaOr4wBUYAnIeRVlY7wOwJ30hvm/RjqOYzoV
5TRv4jNWOeJkUIP4eclaW/o+rtCXE/6RrczZASxFFrV17KEJQza+rhBVdGYESzZC
5FE62p3dVUfFjLbgcWjNSSoY8uITtahxyFQmXVZZ1X3jh5TgxF1OHbwMmRVBE5Ro
Rzu58+pvQyphjqWpl0xQrs5HhjUqZu6v2HxUUr76kiatrlwolnWHcGBKgM+bUsIK
4LjagQOUsdvuzqkrxbP81hzoniNgfmmsx9qEHn44YL7GM03CymJeIW9fZrabWiS/
Tvr/UYF22d2xprD5Nj9CiEYXDVNwRLIO2LWrHPSQMdfGUZa/LAi29Oo79B5shXCU
4HZrb6oDD9mz4mEhNKAkAVoqF89yv6qljDmASyA4Q9CqOqERdfNa29dV0avLNsBM
iUDfyX3sDhp3Kl+Vz4jXqWOqJQHPnCeJnFv3yewoS3us5wkj76f40+9ilLWvOwqU
TR1IMMNVqPyOyJmk+7GdXggVhW23+4ZGqcCy8WpCcLJ0hTdm9td7/Y8Yy21Y4knM
DvBk9jBgbH2YHdhePGJxNs0AddfT+5g+ljrIbpgcl6AzbU1Yst1vcgx5PWOMNj5p
57xvibtPqkLteBTPz4ro2LyvQ8xMBKGMp+HwqxhSEEd+nCl2ap6a2lkK+oaknk+O
yTjs4vWQYqonxsWend+5KLp4CXK8ivTrhp9Rhj/msCLTbEFWajdJyqbIYzxAf9if
Qlxv73HZMb4ApcWoH05xX2VVKjOfTuU3elbM3cHQomXUlPzji353A4O3pvpjzhcz
VARXvLNR2fqSIlSwI00e7PZEATTr+ERpRdUfy65f7eOCE7qTvArj3tHwPjgEg31g
OeZ8OviEwhIbH0cs4EMSM7b9WZPCSc5I3/RIQD7EXqigVnz6VOFiBGYwertdr9d8
c0VboxJq+rsKnmPqIKUpbChDqqDmsot2CxgDHzFuX2ff7GEGpFGZbJNKFGo/9AJi
f76eW5JgHQHvmaW4jXj6a8kX1Z3TjOg8AS9Vect35X4wrHATokx+8G7BORfFBQfe
FMXQAZ8MBVTZ52wtB3DhgeWNsyhovu5yhHHjYPrL9wJ6dZM0VhLhrNJIkfoaqTfn
b5sgrINDyOu14e4NZpO1weQEpclGA7SZ7dxlGef45i6QdleH2Ce+zv4Q9lW9tvI7
7xodvbv9WWZmdFuDrYLQyt4MAt4eLK8Fqkyzd68couUMDxGWsJBGGtQ1Y1yHhw/+
3V0dzxNuuvNkiXs9/9oc1uGlXJKrFr7nXB2DMChgKE5wLYyj8KOK9OQMbiFul+59
+QeyKXLZiYIEjjyvzZbWqsYhlXSQZW0bWUSD8nXo/zlfpAxiuxf8yoKEXA20Qt9F
NEp4Lw0Bxduefxysd8mBRrH45nw/leOlfXOGqR5oUjMdfMlSBZTZlBCI3JwvN+Q8
feZrAY46gImIypI1c1Mpu7/FJtHHjJhSpLlYIFyf4h0ii2TzAn6MFA8TLuX7zgMc
a+M+vKqA6/QzSm29c6GyPg+bTAJ1K7dV34Gu4ZqlCIDGd5ZkPlxbQ1dIkfXt+ved
/qrEC8fgV2Y+UkrxNhCoq/PD3jReGfZKwxOGYLAawXj34uysJBEgyNFmeH4730AG
JrPVGXkuGfA4uVgR1v6vxWd+aZJv91HcHpzlbLuV378/V8T8B5DjFlBplZsvWPEk
6IVNiwUETq0ckBGuk3cVG2Mw1nwmp/7ij+mjLe6pZzsO/Dg37N4wxihJ/kcN7AVY
n8TNiY7udH9qF0M7crsOZKmJcBUj9zMtdVfmfJVXgR5fU3SlTVkOEFSYQWL8yNgW
hWMd7xBhy6sJzI9MoIw7cb9uURlXCkKtc9eob2rVP+G0NcU9oXvn4uNNIcxzTHgF
BKoD31Q2nJfl9Jsz+ugcbSVXqKQX/OPGLCfmvDltP/HmBMTFHfdHYIy35bpPVFY3
Myb7CvY/f+V0gbZAfKLqVhGH3mPUseoT4AL58bXvhynk0TTpEmyU0UXkX/b24LuW
oCfZzKdKG1Qh7FXLaHhMEX3h1aFk0XWJ0plxNxZgVsACX3BMbC7YTB4Hqq/GRbc7
h+NYGoJxN/mTHjoZ9lC51aFu/CnR6YEOsf+/a28Bnemd+3jv2UqO1qGyoWu11vbZ
0RaJQgq8O3EYhyDqaQ9t56ZnspLuMQY5oF9CI58eIjjKluYIKDaf63TbVl3GPimK
Hlvt7yDzIydQnagrOpcvgDseQojlgHpoCtX6vtiCYkZ6MnNzie13Rg6FrOofmcDc
7bStLZI+I3D4686gGgnarVXXSnTkbXPRbHgexuIjDVXVFIUnQMu7JCtzBIaTWxGP
CMbXPUgsZU9JMozjJEBqhU92yRjZ4T8fjvmdQa4Krl+jmQsACD7/bVA4ix2axINA
ynlFe9apCPf+i5PJWo+fQ9YgunLP9qb7UC1H9JiMI2+mdflK8nlGmV3lmXAJWUaB
KASzCK2zzWZ1/3ElcOhMWlmmjI4hzUToUYiaZdMMMMyT9cFNaV9imvsVc9skULdo
/gtPKd8qjLCvAKbEISDIYU+gmzK6YJ+poItGJ3KO328f2OZASyCoeUKRsp02Qxto
N23PMh+WXVDcrsOWLrEMIRMqeF4Y4MEhG4qCV0aca0exxa+8nTFGr5OwYDdF7pa8
BUtDnyhNbt5kRG8TXK0fPuOAM5uJ1zbDWEDIm2jglrvtA0fhbJ+FyIvjA+5vnCVR
nprWM6E94iEjBaKWIZHQ2WiMy4/f/gtLXWB4CXSly6nrqOg70gSoZ6DIJSsWKbmW
/tdfopzzU9VvtfhhxrYiFlVuenhN9e4+wMHfo+N5Sw70Eta5gANRj0oRJC0cvgoR
eHPs558Ze37mbnKpysW3Wb/xO5xFunr2qN9m/adMM6PuMtlWGlZ5DLJCVRlCYmhb
wJbcJs/aybgKPcob5Y3CjiEj3Ynu9CZHexm2kQM+ewnanaY+Im84ZA1EzWT623B8
3Ri48zOzi7wMqPeoGK2Ptd5z0RlJqcpLtn7EQM7krRmhFAofzaD5XLHs0eCCOnsc
ORZWvYEEawp+Z8xl0Sbfy5OListjMpJpBBLbE29rk0n2AVuhawmo6sQZCRnTDKGD
Fzqu4hY9FFVGCWFwPN8sote2MR5NPkbQyrvECpzDewk7NtpXlMGN7uLMVb+1CVoO
CyEiX0aKvASBAhUarzlAxm4HInYBGMiaScF6dLe/99U9wsRdMg2RURpIOAB0XP1v
DyQc/VE/0vt8F7rhE73lD+H0F3AmG1QioXUPPM60/vMf0iO0p5uvv8sH4Y7hGfMK
EsFNx9TiEUKdk1A9Hv/HU2fGEgbNWxr4i0QHoGfChVGnQORZVvQfGPhEfgY3kjN+
P32sSnvmM+WMjp10UltbYnLgBtdCGEdHIR5URnB+DY50QasrGmq54VOESRzGVDHd
bWYoQdYY1wgczo1m449buuRl0WwttR3MmEkmJ0rPmSBLQJ3bopEr8IPTRjk8UrHs
1SXkB9hawrIktwOg4iI/yGHdy1BuSrYAehU2OUcJkJAeywjheAEPVT6eSDy7X62m
AlhsA+curHK/imDTHt8/ZNSJFwfPzW9uA5dOiJNLW8M2tGZHfMr3GWM8E8vPEWWK
oPf4WL9Pu2l8wQ2p1XjcD7HIIOKLF1yfBvAcmaT2UBBccnSCpVOEcAu85ltdN7bh
c9w+faKdsLv0/uTq/AiHjaLAlNK3JKUW94olz38nNq4jp8coMzvXaPIQ2Fdo7Q30
Kbdi+TItVCqqvFxk9BjccRM5mxR7wlFGZY23kVmcA/FQz5j9+vnqChyYVsTENvK8
gnzrjkIbgPfEAtaAaX/hMvg1PNP6sGnKi4SsPadkPD4nNeMnzMfXbn2sROHfO/FQ
Jy5PvJ9jp4aJBhPe9n34gDftkKTxLTO3zd4rAEdXfRE0JXzPzTqyNTOsj4DBHxun
K3pSZdQvDouB+vcFnrxGxjuh3zCqtqbEVzyntuUU2OGcv1duoGbeyvIPAbjzaJV0
+6wBl/TKYWuYB4NatuM2By5mnmo7v/p//TDtg5rfWpYyT43Ma8ACwcxkLhv7+I40
aNchpTcOh5GJBsR6NqMy43hi3kisJ0mMXCKGatS6DAE6JXH4xFisrB/DiwWOU1k2
gHPiozPSr3J0lO7V1zlHDYRMJchU0scx+rj70vYdkph8gi3jv6DF3MHkVLOjBLO5
jYDlHNJw44/8KZSAUlEZw6RObClaEVofWsULJBBdQuPkSCnOkag+gEc1TvVBMWk4
6rxkHKTiQGqdHdjSVkEugb7rCXh2FNUmYw8tvnV2fp5we+vCf4N6eYXcyrfKHJ0a
aa8REXNkqByiK1F9/Dz3JjP7HDLFkRwolba3SVxg63d+0z8oE8LWCxxFK2HHB9Fd
SGYgyHn9LFMoFfnP3RxxteJhNGTxidD+Xd8WzzeyDDhcwK39y5K590HtEa/aY+eb
vJKyDdHVDGOTLegg724KYRlQPoBRtEoiY6nuEoxixVHHR+fD5aZL+9pYgNR6ZeiW
xrI3ZaUxdVJJqlSFnIv3KgpnlglOlMEx07PZ0dRsZxOnfIqwnXRW3Oth9jnCcRPq
ZOkoHD+gRggDYSZxByIXey75iv3cqOzEhByyJx0OOYVpiTUdwRNWFypMM5YwgU3n
4KTwKKRU267JhSg5cM9Jqz9NBTdToNIZ1lI55Az71kYvGKBQC7DWLQuxh7nU1pZM
xBQq4pkJGv/rzPPCffCs7b6yOwW+RTqNgMLLIHkBlaZ/QdcVjtqLiQ3PlSAMZHea
bfdvg7ZoNt1r/kFsq58YYMqNdRtTf4MnuBbFjsBJpytdCrjHgt4VnqR2nbiz49/r
/bDXnfAmzxRL3C1rj/ZACUz4l3QYfNSGzDzk8HCu+b7reAv+cz793B1hMPTOabe0
bDvn3RXw08+NavzolMl2GIN5g2Jy/siu3vjKRmpUWH7f86zSQm24c//eKveOfpOe
BsN5NGQKhex+NwLGbQ5g1I1aH+BZLikUrqzkEMlHKHH73LvsO/PwexHyqvDwAXvm
AJkJtynRPRveiZWvuW0BcBoBb35FSU6U02TAOup9UI25OlNnJ4mJA0mV+lRaVgRZ
hK+3ZlPKWqsn2uP6OCPorncVhAnmB1G32QYArGZZYGYW+uypHbUqgITxW0GYxlPY
m+k5WnwU0nnNXVlWPkUXh2X6HtBdZ+rF76aoFhvblcEQbRwpMbHvOpVO/+HruWrf
WollJ3vSwrej4JKOTXaMXzjQx2Tcs2dRJ+5opqPliihxILMgtiKuC9JnO3VqYETz
lvL7uABibCO03C3Zy+9qDp2zFeKLNM7vVP2Qq2U69lX3jzoUL1tUHUI6beFZxDtB
JhEqNLAQ6OjvHRPIQ8vcPQYQFknQzS1FJb4kCe3cBI9BT1X6G/owLtKkgtc+pdEc
jAtUcNgfcQhRlEBD45mgJaSjyyGc1Q2ewvOJJquzH0sBIxtVV4x1dG3HhDX8/uSU
/rx9cdV2B45apc3J5Ia5kj6eb63JCZdfBz8euXQ9zDaa3oG5PC3eqSyGmhSa9WJa
v7lVslvfLrVqfVVSeiawmu0s8Ey6HI68QODSi7G8mlwgkuFZebvwmjKo6tGSIX8N
uUc6m5rD78GM+dshgLa3G1x+PqJ5f9OFahaX6MSfPPhkBR5bP4HRt8F+9Qag/5A0
UYbIzWZrzly6T6v/ibcTgEpZmbbhdN1cbcs1DYQoUpx7cdoSXMHYKYQ6UtofIpLJ
rp3kfmWM7U7kBF6MuLV64Vf7zUvMuAFr63sZNKNlNFPYw3YUAll73/1m9/Fj7LWj
7V3K85nHVEnKqMKfM8fyyQ2yW8zpDQ8r9OaTgfEFekMLQVHPOIZfagKjAAE0FMZc
8jPkrC3ofNyg08SjAgS1xdSxI038r+tW4JSgk4EwU6ruCs+T/PlVyTAbrCyd09CA
bIDkYyXzqgTEPzWY42noWpyXtYNW71HLIqbnDlngxVwWdWWcp6pSzefj+rF9S+zV
HP8EPj5pYo6Cm54G6+nAdLvtAHCjKukgVY7Pu0dEmvQ8qNnTMHWtLCKcvrLhkzSn
/nBVmPv4WIAvp6rwngeWofPc8Vq4U+cGDxHTlXI3IVlGrEGaKr/mArdQCYYuzC+/
iJGRnnuqJQMiaJ408bHFcbF+nALKgAmqx7A89RCRD0/799KGYS92PvTphzBFoz1X
brKDhLV6n1yODg8lxSgCxxvav1u1a7ELlWOTt00e/d91fBsP4ImgNGwRr7R5jbPJ
mco4dot74JxRGveMnaqCeDpdRcvkdXBpFDUpkBUdwYnusvBfG46An9dLGDZf6dSR
TT8pKxXWmaDSMDqqSnpHxNZ8m+qIfNSh9Ux+fSCSwKPwo4fdd+grlamVoi6q1/Jy
m/NChGcztJmpJaOfkyFJzRrRPhXwTwbJeo+7ovoFk7jw7CGPD07CjesHLcE0hrOa
i5V2g5WvBgjm+8oEwrnJd6DGwWml/7ViPMEedQ5lKqN0jL752CUJn6GGgaZUjtTg
7UpTSngmfGUFLQKcsswj3DbKdsS2+mwNBajSfGJDG7wj6DhW/V2klBtTMYOU5OLu
v7AI/OTl4BpzPakD70+dTfsobncu0O1ON1RlhEy6GEV5ayp4WtM97V+DP5YqM+k2
mDzVL6XprVlWIABsf6rSKC8pCsrgMGPxFyjaucuLlLiABWqh9XGToIzvgwCy+mpf
6tAtW4x8G10MHVSsw1qqgs2Y5dfuCcM0wCGsY9RkPL8qx4hZzcqbyCymGUGEM4R2
U+ahFJ14sq78HUPueVo/bBesRY/adWUA8x/KGm+uPIWWQjAup2wOeS/lpfrEi5+9
byezAjNITdF0PuL/EIG7VgLniAhnpe5HGJG0MKDE9yTD8M3pNGuOzK49ZluKSIUx
nNTUaRR8ry4P7xRGNr88JvsCApmSJmvjfN73cjb4D5iolXY8C5YAb2SA628zwkii
KOPYmpxHnoye9FHBr6BDOq0NEUXLt3R9K9ZpSJxjfwm/31Lp3rPAZqCD4NPdhdEp
sw0YZMRvTEAn1ra+KfRl8shVjx0MCulyjWAp3jKu+dqrwzQFyETH+ULLoyH9a6s7
o3tB0ZmtFBn+9c5fT88YUcpRKLt+NdvoStT3o3DAJqvo2q5tU7AF7SN9CvkXMHiH
PbtRZ8rKy7rw9Nqq7tFX6lsG3/5ZdaSnYJj5WRrXL/f6hw6dWeTeJw4u5fjt1REw
IU6ribPPfYQgAz+lqZcMYGfACDRN20mvZFm2TaAfJ8YUSxf87NqO4SKYfttOVhqr
OP5HTAVhwsaNn40DiVrtPpFQs6zcdGY6HSlCoLuXjbugWeO/e1PLl71NbW4sw/yl
bSLC2vWvgeEacd7xQqTqsq+eHRsGnMil5pWs6qAwAjp/aqeNdKmCLcQyKNAiWW5T
EE0TYyo8xgk3AT8k6PDJ0Z22QLIymHbCfylBsWlylwwku95229aTf1DOp3tBphea
HMvvlFLAFMreTDOxPerxAI3OvyMcS+WUZDSVu1kddwAR56Ob1vpVhifePGW59eJn
pFnpkBt4oiedvFcYkErHlZ+6C/iEyerYx7RjXNlB+2sViQvOgOs5N9IWjqN8HsZF
nrKPbeUvA4g8o0GQ7oIEDS0sCMra1lGVVmq+RW4fXrDQOGJkxx4ke9sJNaBkEpHz
cEQb2ITmu1+A9CZqO4ijkl3aDLAMRkt2FtWxjG0tvD+J/LCGaW/ClnSXwbxo4H9A
0kdNKlZJCuhcb2x06JWsjjTY5vIkEAjoazV0y6roqndJEY02eUjGXeMOUjKAA13S
QZFQAy24CTdwHIMUbM1Ci6yk8Vwzn/pPz9kjtUJGB9+5oAEY4sbSt162IHI8PVvB
SVQPhwGoxzzEEPHAqNrgvWIGKOLcWe8V+/JAwMOmmdj2NVQT4yVB9YuwlCSBlVgt
rcoM0B8KiDHchrFNspqiSWPrxHfdXoQRs/OqsoNzAi86x4YVkfwZluc5P4AXgWTk
2wrMWjS1hdcRK9JzD/759CyOUuUCGWZqFZ2kO/JYJMlj+oY42r2zerellwjky7uS
RBVzaBblK1BJtCEvB3P/6H80i0psu8wxCI2W5GVfJJcMIZSa4JEDFTjAIOgkS1+v
oxGd86YPGnUtoPSJF/bzoMxBZJ8YRTbWelUVnbAz39OGg2kqtrzy1/PENsY03x4i
XV4RBaoLHWyuj3vC+Lzs/0Ridt1T8vq3u4pwr9J5D0IYVLXyQrw8jq4rSdU8Otay
uVY2s4fJ3lFZIBW0LLSVQIRvETnzlU1IlNyh+mQKPcRXyXoHMTQB3rGx/dAnztRU
n9tIv0gmi+tjzgtwJyj/odGuSYciAZYUQ5fD3PrpmX7NXisu53AsHRKJfshz16/S
zAD3E9NB84LOc9+Lu8jxHX4EpVVK+0qJovOCUHkZdiNC/Bj2O9mWhnyzp1xSTw8W
ppdDOT6mjmkA/NWqri71V5M6ZlI0p+2AFyI1T7WOgrF5rYmqWQMY5xF7gpMd0qEy
6wwdxdZEKyNT+8RBGv1gD85DVUGZ9JIFkQEQy9MSMK+XKUbjY6LxcqCwO8a67Q1U
LWdEfdnCSLr+ueM1jPrWLF/9Z5o0UtLEZf4J35jm9w2xVCgSYxqcPFDYyMy5Vwyx
MGl5BaFL2DJSZ0eHXZppvf7RGna6HT1RxEWDmzdNwc+ZhsM6NrWxJjQDx8GTgsch
WJe9AvxtEP4gRIoYNyGchG5WkU1F4PB+1LiCBKoUxtUswNFPhXIBPbLq1hYA5+2t
3lpQHcTxXhCNLcotr0HsjenF583yD8uDZT/LdJNQJSxf+sa7y3S08JXw2sKkaFn5
b0Q6nN39cUka1xMfOB9rPteuL9r2b5QRv1Mhl65t/mZVHICNTE2MnLxMazCQL3CW
nn/wfPTgt2EXQUviS+8S9A7dUY+2i9tsKmfwTQgxNKI+Lx9T+17NqlwbpRL47iPa
jI4tJh0AY2W6dIyRNvXGOzyCoCsYyTN069QFHDkuBFXBFRf1quGarnW9mIQxdRzn
9egjPNLup2rdD2OgNeCtsc9I7el206d7KQHRzdSxYYwlrw6YsB+1dbrei5oJPhLQ
CInfUkDqGvl6jbh6ucj8jmmo2//NnSWOBgu2pr0TPVdXkGWMtXcI2F2OBn77fkIF
feS0ZrOyXcBnuTt5YYiRs3DDrewm//NwQiJ13DxeajhOc1eT3HinxzlZ2upGaGtu
lNntw37gdDivS1k020kA9mopcnn2e9UhEdqbO/DxLfXZzxCoCNCq8KLGpWznslHi
d0zBC2huxfgNDKwhGmKAlGDh1W7SkxE8Mn1/0TjFMMbyqUfXiJCUr2GwUJp+H95J
i2RhDMsoQpHsk22ACz8cHjoHLNum+sasZmqhDZF95JIgrYehfIZ4oo55yk9142+h
8ec2rSG3LXS53B1P/cXgY5uOD1ExjU+ly4H+D8eE1UQOvHt70dQZij4W/sXwT1mC
FJ7sIRncGGKw9aMUiD81eGbm4E0fXcDnn05vdbIfBiI3EqpP4C4BjGnv6y6LN/Q3
rSL0lnUJwL2KooGQ+5sVRoObmegAJebiAMV/hQ2N4vv6INOmE5YoZVpCXSd3Abul
EK469xoLfeBvPtfCBpJk7idCjDyRvE9DM96tJe6tQG0W0S1ECVcJBxQdGRTIhVny
A2p/OJGQCAUkYUsdvWeY696N2lqyPPqu4KradqJXC82kI9+siEA4fZ5MjwDTMU6C
v13hZHRI7/cVAi+PwREA4EKSRB0ar7c4r81pAy22dx2674fxFosmaipP3qGTOKNR
nFGs1H+OTtZ6bRFz8bCfpvdNqfGgcxWtmQnLzSoYsOt5GgDveRi4eUxgIMErwYYQ
QES9U4s4SO+xxZv2iks/NYKY837HL/9UuDekUQyYfLTr3Zc1977OY5+l0dJhktdM
FKC5xHvLLSeK98E9GwvlqvJfaJcDL4Q4lOLoX+4x3xWHRrpjpo/mtQtmUnUAbgEy
PjXoSc+fazoRqPKtFzZighboIELfrt7Z86UJBBWgMv6Cj3SUp0X0qwo+n7E0Ooh1
3s9w78+5BqieuI23QAx8C0Rbf+RtuWHnxtNiK+fYFoXrusuxSOCSb9xSQd5qP2rq
GtzAU3Yduuz2qOpy7vLXJkSOXJrDH4f2aA9SmZT//tppogXFyRhTasYGuyW9pVXy
M5zlFi46DkxgGT/6iRqsIhlqhlXxw33fIriv6rqrNBaQvrSHmhm6z6gGwfDVAnqx
ozPWHp2KJ2IfAZb7afXyUoOu1cJxaTVRzBCqFVkqy771l5KyOdJ7Cr4CV0Jrw6wC
deWxADEba78nnQeSMB5T7IoftyzHQgWilwVVHAk8ql7M1q+8Gf7UDvv29SEpV3r4
KdR9mfGmjSX+JvmZ6QYfdrRbK+BAboacoxwJ3kepuC8sj6yAUHDrdp+yUk/WgCEX
s4yxp2yrznM4n6ncBzqEyGuNXcVKBjpW8VG5Ye5uQfZWWLOSf9gWxOd+CTO0wT5w
e0Nw1tW7tiaqyuNsJQoBxp68i/TNNGkk47UuwTlg5ZXkZFc6kC6cx+4RBE4fmucN
MlIGhnrik3ti9gTRCLW4xfuOuDydrK+lt3hiDk8K+nIid76RArMspwVmT7bjDNZ5
OrAE1sRHU4B+vT9pJ8NT2mk4xbGcqyB8oA3Gn21kYNWNXvsffwOUoy59Jkn6hceQ
2QMsGtYPDyuB3QZs3/6mui+VYGV8lnWyHeUqjdt96F3LuXC02DKfptN53/bmJIVO
f0gq8YGm6zq4bJQI2fJYdIi7+ASEfYTfqK2D8wmKqP/zOARDzWpRj8nurfYDZfHT
aI7DQ6GyQtwKE5AsG7IJmPcUiAdEWTpKkQVlQt+aH+/5YpElcxVMPa4We0gSXYux
zZh7ZyFBQZO8sgjPx5VKr/HcKT4vlaaEzqmLhMFjbBRAZqbPyGYhBjRHTGGgILOP
1CUiHpMXRxQJrqK72VlT60a1fo/jOrVS78hEIF6rKWFTV1ny98AAiRJPd/ND/YVq
W7v01r9XnPAmO1fZcD25u8PWuRcJ5lqQgyZSEqUM6aKVQUibxlphoMd7Qva2AYxB
CLa5SncmCv3RyvMrO+3kljITaCoPQ4Lz1DuYyzmdk7SsZauISD6YliMQy5EDMtVc
WKCS1QlURAM+2dhMSIEFn73LUSbmOkukx84rdVTauifctH6dSFnuqdhPouA2ELA1
n6End3r1mYvDiwLAAkUIV32w/3q+IkkGe/PbxvwOM/16Kvt7mJS+PdUVYfTW2QHv
5GbH6GuLiZM0mxcsWJiZEIHeGCak7DkEEUrI6B2qrhlcewclsyzALhMeuc+7tcrm
drR//TYa2gndGXMympwPNoo/0kaIe+aEVDNPAfhQAxxE28YkoQ6RoZxYakrXEadD
SZIFLrkp88fEoazAuppUKC0kyL50lE6pn/7AVYvqMqllqZRVM8frpgaiwqijzQRY
STdNOxB5UZuJSf2rWhDRvXWIKo6qgFmPkb4zMoRMelrPMAqiDdnb6noGhFwiiGrV
rGn5/3rXvskJCn/jSY3AdNXd0afUj0bVe0getLyUu+1y0d8l4gFgDuwT47FHI93q
2fI1y0TQHrYDXbRNiS6I1aBR0dIdeTCyhPIqnZBjVJkObeYPtppg3nIR2EbMOj9W
+xmMlPEUdtfL+oNqR3dh9u3S2wqJA7/o80DxA5qyJgOTA3Y8XzBZNrg7S6NwcLkw
oV5eTpWg37DTCnKn7jqb7IySTYWirqyxwmdS6Pfzl8HBSWQZ0qM910roClwH7wZa
UNOIdA5dKj6xM4SgPDLbLxG8SHSEQ29o/PgtF8e0gRR4tJGWVz3pfXh/ZwRpVsxq
e/z1ANf+k7Pz+YcrIgQlk3gIJnDceBWPIc487c/rxFpwDZLrq7rv3+WqW1Vo70ff
HmPEzOMnpkdMeqAuBqJgxKxx3rLXOXNbVXzPzK3EflyQGLvl70OUH9rjd+gwJPu7
2k8MILmOJYGN57dwx2WCYC11Rdgnyyi0crPdThgzl5+4vUalPZKvsuMbRLSD3ny+
MnGDov+vcputk0dQU7KKbh8dwZ2nkZcaSg6sDf3iUA12sLI9J4GXJbVwNGLjWfuO
YcisdP+B+wEovQZlYEofn9OpvgMm6Uvo51vQYarko3ZEQBdEgcvXSFQz8QKeipIh
Sbd2LFSXmAo5BMvgqDbJNcO2eGtg6ogZNzOpsgunV5TNnxRskBhQmEKB54WXq9u4
DHNnkgl/j9IwHDoYim+b7NLREuS4vZ//+tqUQkHtPOdbH3ns9bFLa7CH9FrtyiXU
+72pryhPfOwsrfyMQ4htORbvQiLmhHqZrmqSj4lkoCeMNjhNyYE2HjjPu1oIIgJg
Ph+1ZjQ2IWoDuvKWjPUhFRGA241QIVc1eKzdJMzIGZxoX5RrFdxBE9Q+OirBmtP4
qrnXXw/c+q8JhVHktItZQQCbCFpCE2qRIBHExaQCzZqJQA6G6vPSe9Wa08COTrAO
s96JKrZ1V15lke5/+0afqPkICHpNetIEuXaRMUImbhv3qrcJLkEwGnsglAEHXjDs
iIxVxTDd1mXy52+i9ZGH5UmaFloFvWcokakdWih7S1hFno5B63fr3eQCYnWGyQgg
s5wIuG1VI9cvu9Nm4cQqWl3Ts9UJF5mvJBC4tYZ98KhMjG7uOJtbJzLorWocjxAZ
H4NuVsLkQK+htIEE4ott/j8mH3IarbTJgQOyeVplyxNHliR0upL+AP4kzQAqqeGn
+Ai9KzBTuAGYOsu+tTm13CPMk6siB3A7mDrIYTJVcHQi5l+KwVJRLeo0BxSYXgFU
n5bB4kEcDO65WOypoy3CwA8VYvXP53Afv6ISbA5X9W7w73al8djhvsxcXthcJFa7
A0aj291+IRwQZshGlYv8TZh2il8oIs5toISJw2DZYv1f8V71/+4JYw1I7gVLkbZm
cFkoNh+UlfEvOxOMpGHIiYoCpwC8AOuobW4N7p4L6y/x9WdKn+08ctFaasEYFnwI
nN1jz4kMbFbM/IuQzCYyToFud96cNCcO+ggW9SS3yfqvM+OfsPHre7AJSoW22Tz4
QRjgqIvWZHa4Xn1whq1QfZiSuCisiw0dRSmb3tXucMkptS9q+c6yHzjbcwzwwUZ1
CDKa5jGmZ0KF5uzdKvuYL2JePqBn6Gte3zD1bTN55CZC/gaBs5+bFx+2cGZKhHAw
NgRo1Uq+2la5WuG+0CPA7QgspoKQvJAqZxcVUxUQjXWyUcqhzoOhkVXXkBWVPEEM
83HytNTRF2UhgqhlzC+zIeOTRxpEvn7XFMf7IPcrC4QDYg6YHi2GAfwKNOS+6PJf
9yT3JNPgT9kwYmmIX1VHYgGuCtGOv5FvTzt4tnmSxEFbyTl3sErYR+4VMaACBHeM
A7bUrda5z3Lp6ZE9TFsniO/875Zh7aXbh0XFcMk+GMfAxJSLrCfY1DDPh+XM703N
LWEHfO2ypR86mtZslQSV0xDjrbQtHoS2hjAMr8WqxmQFc5Mhi4Ur/qqxmn7RweTD
6lxjNhcc935S4VZ4SQjJsXAJZdqb1qhnsa8qV4k7J3c6TV1cq6JtghBmLIJHNDX/
Z+IBR39fNh03cwfTWKnD4/5e/E0VLEozgeBuWoJZpCggx6p/9C0IvzeoOmiyrR4m
LPYErF0i8yaRFSvQYRBBsp75uVLKZ89dCd4Xwm7fiK3w5rVCPhFvCSXf+XvHMjmy
Tl4iJ2jljBvoHCaQEDFXpC4nEGKOy32h9yum4MR6q045pjb4wWvZwQoofAk0s3f5
QwEAc57eythEw8v3eFXTdaSgqKhI95yOz6FFL4+KyvuSLZ3jjhJVGLPZ68Ksx6Bl
V4EVVFEmIeql2aSaAzGDrc19912IcqagOyshiIkbbXouhP8+G4FHNbo0tUsqW5Pg
eUT//qIM/id73doi1oqHKivD3jcE2mOrxzd9a2wK71072j3PDWzgfmN1viABFHTN
Ah1VW+Zi0xEOEKy9tyfByY4jATo1rplL+V+YCevZL0VDAscM9TwxBsTVVB9YlHw4
Cspjzp1JAYgjPabh6xNmyst9qalhbvlGi3ucefoPgZBC1rYGCV408eJDgVI5uUIz
n9tytlIQCDQ46l2/ka514wsZ//CJtpLEB+6Y9eaqNtrlUwEzDVZGIYk65AgJznZK
OAgBWuoDHHwj5dJ5QxG7M9R9623N/NJXG0qr7kgwSG/xb9MarE0jN2iC7g1USdjG
nAk6fODa8JvBA3u8I3n2IdEDzy1+gPyEYWPXPZksunV6HU8NOjC4dDQu2lxyUi1Q
Tn8en4oV2ae31xLwluudqtRvooZIr2QeXc5UdZltjkX8E9yTODUaNCXc8T8wT30U
Tf7QD53RDPPF2R1J+NDU0Vsk08bmtOsDO9vN1AqNcZ0znKNgJDyHUIazh6zr04e2
9aIoZNog3cCnREP0nkFDqByGHpI4vGh8e2I+w9AcYHM5Dx0gAUROs8llJolDuvgu
tuL235FrdvHNEiIxhlFVE97wD0q8x5shnza9ZrklaUV6wlE3ZnwzwjHBjdh3Czuj
u/+RfYZwO13SaYAGInhSq4SJWF87FLPb0+KtdDvSLakvY7voRdtOaLb/IDRBi3MQ
ZpPDqzoXdgUOR1+lowauyPD5JMDkP/JwGuDkL28rdq1XdiRTmZsyb3Ejza24MI4m
gKI7yvadethB2sDOoQKfetAPGDVrlnCR6Zpd2FslLHc0x4zPUzIIuOdK+b6gttbq
LihvVjxBO9v5ErV5EyS5CAhHjjvUzU8CEPGxnS8nYzatILQhYqWmT5/84Nsq7jac
/+qWrZdQ5hCkBqxz+ntUZOhqOm6NaovWcDsUQpZ7GTDou+19PmqaaldIcdsUjHvP
KqGH+6P3M4ObhyOi3K6r1Xauz5LGSfpiNelZkj4VzsGXXuvB27gDev2o/Ouc/+M4
wspTc29AuKm0jDUBdVr51EoIoCa8YbGdjv0K9IVHAY81PmeP/kS5xukiVbGlcM11
gjBCOmdtXA3KLTtPvHwRJDCMrJW+mAdTwKLpV35evkwZB/QkGbV8ntWKEZD9fRq2
TyR4bDbA/FzmWKAs9/sQAUqVrNLdWkHCcqzkNoNKUheU4H2+GIOtkgbNOVgJl/K8
MAyQQy+cb+aBECWu/URjCpYM2LJWJA8/gMrVlzFe+Qn9rUg1kNRhXyvwXX3g05m7
DsGnlcCSRK+hn0TYZ8067bl5adJ/D9+l1bIlYPCEhzaqXjMiWyoiJtzop1cC8pFX
mIzYmu6gY3ePN2CQY7LZrYsAe+YZHjicDgN2Le4WT4x6rYnQGI8VuT7J+jsgME9W
TZiiNEJVOlCAYLApyg2dSg9r/sZJq4jJwV95ePHhzkF1cSNVl5H++YMJF6SYUmwS
Y3YEpiOf68nalFNkAuE82P7JflMtREQWncBw0bLDEIvGA9SEsE14i9PMsQ8qXqox
eC/+CWXGMXDe0CazfkKbf1W2qN19C+x6ffBvpQ9zdUhs8snahY/Y1VH6dEpvgNmJ
+gfJ3olj6gS2Bq28YzXgWBEOuajZqnb7YfL9xHHywNMf/5pUA50Z3UuQG8wLjzaG
qg3Wx/beaGttFe9C2kyTA+ngquSE2fBelhh5+E1tjRMA379FjARnVlyBMiYS7m+F
r3xSjf1J7qYXZOkL0UCwEF25KM12sCtPLHBJjMCdGKoMSVxKfpVIovJqOUClxG3M
ZrJgK3mVneqbyy9R9CcX0V1jlRWncofIXXnhi8HYyOZTh84nCidFvJC2Euigcvrl
QtV05b0aPIpMCeICDCEXBmqES160g8sPWGpHgg0WghhxbLxV0i3WkZMqx4GgCPAv
NXYGkIPeI0UHJdmjWeKIA228gbNEuXnsKQF3/jBBovXGqX9fal+s17BzkqON6idg
fy+4Oe8I08TM1xQJmMlQ/Y8lKdzS3NPbLiWk4laTK8pChbMRD8wDMIlBpq5Inunc
Q8Te0jPGPhUPbUluaiMI3Dcw09RCPj55Ifqc6Y9jmmru8r+7r0J5spI91f+xMFqT
E3Mng+GPdND6OOWu+pAhK0UFdn/Qv3BrF9pROwyIFVQELwPNJLaA8YJQLO6Zhh7y
y65Ynq3T1CTLsD30sk+egH58utGxhYy7/3P2cenkOAS2m2ieVW4O2dEHX4Frrptt
C87nPwnDb7GWzjkLC2Z9cu88HRpUQMdq310WPBy7UnQMZsDxC3xsTj+cUJXIUOtM
0NFqdKQT9cJZlFRnnP257ilcwykjyrfDhZlJJ/1bDeRPQ051sqfqvVNDEvNHsfC2
THJrxo568zuFeoJsKKSaDx0yCMQsYx3VOk9zpQvNqoY0M0Qb0s7R660LJ4QE7bz+
GnpC9Sw36z9W9jZrVlgvi1rMZUI2Wh0WJs4pnhRAQs6+1YJQ8YiLcigXfnH7T982
mhWzGqpWdh5csMNJyyCD6Zww2rmBh7Mk0umWi9HuZNBJRaas2SgSYuW0bHQs6Osi
Zn+3GBJtwJcK3CjgjEF/wiW9wDWoH3GWTTbivHaiq/pb6GieQDKttzONoj7d2tRb
Kr2NlDwT5l1ZUMIbcw1DEyxP+1AtXHc0zFB17uscqB7NnmFqIhSv4bQWc8+dE3BE
gfqwMxFSAcZabpUVxQQ6piW9YCmTRrKrzVvPBkwr0AGy304cCCfWynFYQssbsnCO
lWAM0VVyEC6uLGKFvzyen5UcZOX6DmmllMBePD4cJ13r3MgmEsfUFG/j4gYybq2k
JnNV5sb5Sap5DpyEycQelT/PudeDzpCaO4GvN8sVvJtFKQ+h6G6/MIRpPRlvDc9z
AoMBLt7C5XWwNFoB2RzNoVuQMM0Q13T0WvOThNePvi8nLtFRlOtAc4fFfvWGXPlW
ojuvQONTN1Obe2GVHZ+YEg9QNlX+Nd1CDb3lkuEZDV20h43L8nBmO/OY7y5pG1Rx
+NCq+MtCX8Q6C/nu/Q5UykeAsKqcrN3vGv876ZoCX6OCym+2fkW+SnvicTn3JGlN
vC/NdkaOqMhbvoByjGRV+EpAyuM4mBiUC3Yi5KAKs4sos6ptkV0rJF2PXzKGH9tg
Iki2d35RY1c3bA5h2peAW28NYNZd3tg9U0qPvWPqFteYT/dkY8josQeH15c08MYz
S9ft7T6zzLrQOxzKTyarlRe0DECKXC1C8KJDvk1QYapUC7y6QC6D/mPBaocrvska
DUAiiIyVyU/w11xdcl043OJT5g0bgsJzuctgDPkGQEqCiiu1/3x1/h5ih/iIG5ri
+KR97FvwxSj6ULrleo0IRNvVH1sU4/mpZMbqgsdbSmYCeeMUAmyKegaw1c+kCna3
9DL9Z3ud85BkgdoLSBapNvwNVAAHL/rHNqjIUcSMqG4a3nW3PJfPR7O1Iydr38Lk
fKaMO6tsPGVAVcR0f/aSofePKvO7Kf9DGq2lEpqg7itqM/VsupMNh6RKBpq/r7BI
c6ePNs0yNhx1ausYgAmZDm1XGObyoRkxH7ZoiM8uwvLW48jJIbOQOJ9B5K8YhVVS
qnOU14+RwfNCjHXiAq3iTcATc/3cWpWM4LlcIcACKAwR5Bdq64uNuZsIRSFutSl/
D45GklQXPjHgx4YVFCJjgcg2g6eiotpup/y0D2unoqwVyN9xQSG4k73Dzfk0rYHg
U1lEPRgvhhTfMMZB4/5tOYIAAArFvTjL79CiIIRAgeHYp98XlcLCUikISgoosl6S
CDabNy9/k9LbqmT1D2Dns74WYD3eoYJZxJNNArDZfu3+Zt0ieI3+MHV8qW6cxfuC
xxgizJW8yfsYPEs+xkBpoAmTur2j2XhKcdlRXIApikVGGwH8RVQgTnQqr9FAx8oq
Xwn7eaWnDzMjmrujTzvD/UKhOYdrVESQzSz8WujRFlXgHnv2+QuIyUH8ccYaHodn
WKCZ8LrpN5rSIltOlfGJ5RsOBSE2+W2Dh1KsLYVYzR5Zjvj3eR8lslOxLjx12G2M
VI7FxHwOvo0GJlhouVO3Va7jGGbKZ9meY5KBjvZ36BMN/RiyAuyfEGR3vIBOPdWZ
tgtYNrYx4gvUfp5gY5QcrhzArvE/BrqgYa3Hip0kEyaU8c5MUCVfZZgkNe1ikjkL
pmqxlQlwE6G/5PSJPuzavSN5wMbUfupC7r7bq32Jr7vzDMuFn9AmPWXc90LKK6zE
1+SR+aB0WwHWUAkr397KGA3ho4Hm8SFw88VPoKDHMxPL1gzG1/809+GDbzLME5x7
sm4po2//lNk35cVeOaxMeNUA27w+r/jivjp8fRZ9G7kjdx5I3eQnfqnibqFDsiEJ
25Vgs1SiM2/p9oVHVoCVWnuMCqiDkLt3zpO/8FJ7ql4MSTsM/zMzxtc7Y3/ZHrlp
VfMfkG69uCjyGPmriv0h1dtB7+CR85+LwMcijb70eCtq9pqyixfCJnSHvrrZHIGY
BNJb/fr0DrrqpL7DL5xTTo/lW4clvAPB4vTjC0CjGCc/5sT6RxNMRb24U96KmIMV
YElKduHc/Jwv9tYI/hRvclU54BgSbjz94WEvqI9p6SKoi9xRit4nQBoP6EV+T+zq
6ZPxPSauyDem0PoRs7GtIQNYf5g+Zdyp9XaAnYsnYBgG4q4TvYbdWBzuya9kMVTm
aRafTKu0KtPS89xI25xULC9QRPqoIanAZ3IZCI21MmAHj2mBrLGxd6ZZDrB+NxcD
0DDhEd1AFJpBKosdQYVVPZCKbkQnZgtTV1l0t9LYIxNbUlYKKJILLNYz2DKoKIVI
2xGhAZvVDEeh+yAPmx1igX6v3Nkv9zmij+Nbc6W+vESoC/B8aEUvNHJvDYFZZbqS
PXjN2ZckVYPQ8IcgK6PihqW2UqVJmCO9aXyKglBhLh8iC0KRkUsgQ6JhDbkS8rEB
QPqZoB0KlQPns/2VtQVoMKNSlirlrAXHIgpX3R7PcgW2nU0TNeexQzCRZEhRKot1
fSeM5F3DpH3FlOrpY+YCY3m/fMXFEc2XDgSOchDktx8M8KKGiZhDmVTO95cJkMcW
weqtWrs6CjpB9FxccXVH8Vc/h9FhqpImCdHG1gm309Xl8BqTIDy5lYgGbHhoKFlT
AO/WoIiHygfp190ahEvwkMebsMhu13F/FVF3O8nj3WGd5WKrK+xTcr4uqkfD6llR
XfGVKNycwUin8EbmdcBQZ5ECntILrizq60rRphviaE6xJCDPtBBT6to5gHrZNLML
EUZ+ZBzt8upkqrIGC0azj3lxRJ42YuhURYHyjEmgBFSUFlpYw7tM4KUnykxvlv1T
Y32wo0BzdOkxX36cJ4TcBuE79f4KQAE9bFHFLrqDGT05NO1uSsddkhqMxm4qsqUG
B089EMPQtBLH3267BvXsMJYzsOK5yG6l6ULYQ7VBKIAPh2Y4lJeySd6i0oDjLCg6
rTA6u9rkY8CmFuZFkd7wLn8OCgwjUJcYLWeoe16GcuDntu3Qj/vq3lw1CEEf8T2r
Oju5N/GS8NP5UuyU1bb2O5YDXa+7z4JO42MGtuW5O2rJMoHQjkjvSKQbksq/gFLW
91Tqasx7dIj6OitGxh9jZjQkAhYeN5l6HBa7pteC86gYb6rF1c6SiqfvgjARLL4u
4uoS+iJB/X8sX1VZ0Dyh1E87jmeOPZopr1EPmfLez3dgVo5RaurDaNb+s1pxDdZ/
oXAjK8L16j/bmqHhNSRBByuKaHskub8q1efV6AEO7h06n+e0N6RZNa9sN7rF4bvq
Cq2EMqJZw/uPofOaWI2/aBaj3snQCc43o1klh/bx9UbcPCzxs7uS8O2NrRnyRBMg
wbAgwapAgWB/G8IdJVInwraRAfhJMeuCXrvGU43wPahfLBfH68c38wKKYUp/gi23
e/+4T8SGtXd0/ebdow0gNtYQpZLAAG7Xy0NWQLTY+QIbm7TJTDTp09Tb3WxgpU7k
HO06XxszXFtarxjOaQHf2biFRwVSRjNxSCVdN4vczCrDIpNWYHqzSIiUHIlQTaOs
t+Ytj5UoT3voqKpEnJto6y7hiUlsLkPJifutLHT3AnIwBS6SFQDB14iorNiSgIBz
4yW5O68ld62/yZdMpQ192969LQxouvGwt7clT0aqiKQ6VfLzvfG7q68J36erQug5
oQ7JMM7YOUmQJpUstPDlVSZ5a11GnFBnQ18u6biOtSdiJHphYZXXTGNuT2THarNB
61Eby26FtCPU7mR1CRiav5M6PwfpA4yALnLqB4D7jJHCUv3JwQZiOvv5FUOsYrPW
F+TxLk4L6Zjs64C2Ry4+mnm9+rZsvxIjoHL6k6/NmbUiVb9IBWGWq1bCtdkwrlzq
k2uNHjP6oJVAv4+lGs1SDMOSsymJdKFFTFYQ9mToF2Q+q0qaEwpWKjDv8aO9JLJH
rrgFha9LAkbmw/Nq7EQwuA3HjWe7suSIGFMuHvhIoNBIJ5Qrtb2d7CRSSOkr8bYm
VVhrcoovzfWpM1Rk3Gj3rHKYnELLwMf6Va2YBSJviungQyu2h6EBHiuIX4OcQ/if
avrVKQkrI5nmqqdzid7WzSJCJugtU7iBeMNpIWDm/xk/HVVTV/Dj2N9NLzC81a+r
41hacS1SkjO/PHY7HzRUeZhqIM0llM8J19rZ8zGYVmkQe4+p0UhBZ6yL62dWwQtb
/7zjdSj9fHquIXwQ9tasUoR14t1/ri6xGNRixWaHgDMRH3OZZ2TiYtin4F+ejEOf
dIoAUmIDbZ0Z1vm6v4Qpbyw1HqtyLpNqTr2iYZhLnUPywPdM3k83g+ZQ1pMmQyIN
VhJNgYZXlpex0N9TFvP6ee0IH24WxjqiXYR3e2R24pDwGCa3HPQgB5T4R5sCFD1t
R1jmMwmgXxqEj73LadboAnac4n4i4bBdk/7qv8hwN69EQ/fYRxoldUfm1ekuv7nE
7WwOnXDtoO/SHWk69DSh4nUF6RDSxga9dWInocI/VvBA+Y+x/9AjvjIPVFhmaaWp
o2O6E8NO0wbdw/EqAQnsi+hiCygcE7yS9mdgxNZiN9k1RSAlzkJL0LLAx9srDp0f
+n/9mMgvJwzZPdgmmnxQGnArpL0hKbBAz/4Iynjf4jmg9CvUFHV+Mu1lxhqvhdPI
Lahuelt8dpbo8nI7bGxKP+MIg8PGWf/+loHhKHww2vLCVv5MBWF+4X+Fp4qJf522
PGB9stSvICFVybK9IqF7bqRtqmm2Du4p35vT6szcwx00BOT3imfGNRkFAZ1KVEvv
hBCNLb+iBz2fM00DZ8QuTXi4bNudnaWkYhg+L3of9YiAY6SvbRHF7/T8kZcKL8xE
Id37miN3HvEX5eUdR289E3vpEYtZ/My/E2e3Z0ZhhT01STMasiFdeKEONu6sScjY
9yrn62Ln76bcOb6HLI+r04RRGJx5UrtfEiKdli0JIOxi+fqMlo/MzJhJjL95xRWV
eGS0ORH5kkrNo2Q7vrk+fJG5B04tcyQFJzNukJImy0hYT95lB8ya7mDAYLZiNpkT
1njcLyu9VqXgV9MxQl8KBouEA83BhVvhRCMQcyfAiCD98wzjgAH8J4a9u2oWZ3R9
0TD9SL3T00+PfABB7fMKQB5ZOeoQu9+TCn9HPCz4PgsqTBcO10z0vmFh3lp2dyPO
XNA51BVafzFbJl0o3aKI1SaMljW3dXACyRc5mREtSWiKR5v4iHbQyE6/7tIEwHE9
vspcS3xwP90nZoi6aDL0tAyE9pF4Jf2eqnjmx8WtcsTVBo6E/NyYePMs1vtod2Hw
Dtt2R6WiBpVAmqipY30rS5L8SzwUzMIELVtTevgdEXGlhpL+OSKn9i6Ir3Z65D4G
w5P/HpkK3hORKR7+lsAbhnueREMG6xhMhYvnYsU+1zhSGxSNg6EhOUWZ1E2mva4l
M5uYkyw3N591D1BB0Pg51qn4JSDNDPFn1U1STt+ywUJTC/ECSS1rDuAZtMmHtl4w
UZiozyD8HUfgs/k5U+PTRRQ7rdnONt7UKyAxEGhPHWqMimD96kbTU6ItBc+Y0bjp
Vnsgohgj4PKwjEoG+4kQmPuagXZs5U+cg9jOSOQe8VEqiQkjmoH05xGHNFjlbflX
`pragma protect end_protected
