// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:50 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Z+Mi1/mqHTdtanagCSRk+kAJAYiQWNEhEkYJII3z6WMbpn7IfkJoq1WJlozt1Z/p
OcASSTN9AAGLB5vaxyfkoQmrclj0F0QxG+7X7hu6wQT5zpzVVXkhTY2kQPtbsU0n
ucaQa8Nsrs0AvSFG2VE6/dE45W0nFKQgSAl/zMTMcFo=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 2576)
pLIX5K9GMAEKUU6oa18h0wfqSJQnglajXKuuvKyxFxDQMucegecBE1cd9jXlaEPh
77+eDKr6fp7XCgD8zjZChj8CsBFE7J5VTOBHdZ7ZOwvT9RD2/izZqDLOyfe1y4kU
0OR19R9bqpBpwareZ6K2lIKvgk5AOJtg9mcYjTPjrFm2Ud4clJ9WfhsGUesYw9MU
wpy21drU1RPODYKLPhKmcP9fQ+KM83mtgaQDNvKb9hD018zbk4dYwF56tca2IVdT
W3ru4DsHrGN08x7kkO+FQcAwuZpXDAMEdzhPkxZM9EcYrIMH0FlLgjUhSi9KKdiF
u33C28U3fGUU9kNELRhuvggaAPk6muHvAn9TXfyf9agyKvxqU09T2xJnNwBcWZNm
8uUeIMKs2Gw3gZA/rzJo4Gw5Fch2ldqWnTgSg+wWaQbDuDMifJbuo5oszESglK3D
+wx4COHGIvqTB5QOIDF1VjgcISCkCI/Xxp70FTWnOCmxvF6Prh3RBa4yxxV7ajVR
0ngc9n0bdDOyidSSp4aq2Mdisy4FCBCIFbyiBa600S1uqDkIYxKOlRm9h0O93tpr
vtNoHUdNDS+uYzqgaHDkb5et33rSruuthfAuu3K+W8tVk9pkOVlSHcIwH8GJCgj7
YoCLoZpywE4NqL9BBz1jBWn+D91cmaoaa/PMN+BgWKCyA3p09WFWwqAts2bvjTjV
b5E5xXKfyjBemD1w7UB12uJwwtAXJrSCYjCOgUR6B+6y0EGx8N67Z1aMAYv2j39p
tmFssEjHfU4Urr2ItW3tq2+oxE8dq5in+pxhhcp7DJ3DljP1fVzMN9psL70EN0LF
Hw2cKYXxxheV3yRYWn50NILNnw7xQNo8wmph1URW4l2H3m/JU7Z73FTerRbRk0UR
MwU6lzW6PEyCqc+uhdn2aQxmM/mWrrdbJmZKYi2/KpKS8n5kmPL9IPuaconlW0Al
FSQnsxsqVq6QI5nG9qQJVwC5d8i55GbqCmieOvSGeKHpWUWl4i8c7pCCMijqyAgC
sfpDEFsiD3R9yVHou8m1wkm5DtJXcFM9C30h9rRHSxBvOykOl0Qvt2vn/7lZoAzG
RyXs5g6H3JW++87dUNhc92EpVwa51qjWVMClKE+PtUgI3bmsCOO1zsFucBlOYQn/
kgL6i6biyhqx5ZThALRJr1yPLLPX7dB/B9caG5CKHosaZicTou7HJnj+KUrkWKwb
LBPbvJpnPjiZy+XB+qfMMub6kHo7MMWFt9WzYWiW1YJDJ8F+h6FAFV4buJ4DyFAu
NLlvia6Tjdkit+jobDNUPqBw82Rss+l/IyILDbR13nc5nBqVXxcqbvYvmcTseBWN
AlwK9h/tGRtang5h0qxKmLXg+G9Bkvhhl33rtH/KM0Jg2leQ4LHzaTQrALgr0yEs
q752wDbwwHV9XNcQOp8R62pFwODwex+8Y9qBMy1qpFqZaPFJjoPrmXDxq5z6u6my
UzlWuJ39GMHqbSNAqOFBQSBq19FjhlpZkEcwVnsSnDQbnMMBJ+3urxR1AvkKtC09
xoZ6byDiwF7f2VOZ2Q15Gije/2bLrhU91UM36B/lYDZlh8PGgP24/8zPv/ZCaieq
mbxDQBKDgD0Blgr7Zqtqf9GMEvHR5YFwufywx45fFv/eQM2S9jEZRuralCu0llR/
pYdM81Z4WzF0+M3LTUC8yK+nOjFNOCgNC3+EjqZ70msqnqEw0Ix8BLwLBCqgA5ep
CnfqrnBpHbNdlUat3UqwrZ3DR3kFw03pOAJjDD01oa1RmuwIB113RnRCAWCryfUO
r4eMC4G5IQu9T8WaaaDudAhmNLKgEZLLZhWhTAyWlIbp6qfoV9kOi28S5RS2wZY0
Zfj+IJE37OtJagzO8WAv7HrqnDuoB+PHWuceK/BGOw0eMXenBoTliRVcQvXLL3eq
305K/ZnMoQC1Idi/sehT2Ri+JMf2wZv2pO8jqRsy9167S9Plbx0pbTfsjUna54ti
jHG/EgRfeEPXtNdcWxH1BCHWwx0jyWNNZmjwacedr5QdcGIUg1MSyyxe0nEJIbf9
VB41xHUFQ3at938I1YcOu2eQXI1tNrmJZhD+/t8EjxnmjUbIHaJESDrKZ2Up7LVb
KKpN6nm05nurQSwoQQG37/0lOMZy0pJ4ZHmQR6PyUjRQKvzr00Y/RQM+MXn46Vb7
plxD+YDNI6iIVexdqBmQZxdXvQYxKAN/aTRYP55v82gE67fB1KOBdQrKlm6TgLY7
J5TowJfSY41NujsVDL0EcSvEATApGcQxmvSp89tndqdKC9w1aXjZ43n3QvO9LzKF
VOwmp1JTuzcnVj2L20zDwX4uk/TBYIj1LEWs01PbyBPoTLwHx+oKlaj5BFaBrHRU
JhPOjobuUM4p5+tXdYt4h67kAmL14qh1bEzbDZadDoSi97XE0wPGR12HG4w/f2xi
+wFRsjuRj9Rrpvun3hIGkBpMqt9uKluGKIc/CUqgSIElLkaWrrnrYenRdcgC+lOn
NgqO1Fm+OP87Kz8HIlqFkLItUkc3VntfuOoULBOzyoBoMEmbtmuA7QONCZBskVxt
CN+geMAymFb7cQFoIJRDHifXsSb3diFVzbN5DVd/ZbHkzpUSv0uPbhZREIthroNb
64y0xPkymVs1rEVpq8hGYFkE7U+5JUWT/wjOeJsLysdvs73CVYL6ogSUuv7BGOdk
nM+bxhjMWb4U+bEUmgNancVylqBTII2PFmw1/dWWZXL3vI9HjST5Srn5pWkLBldY
MJRjbIcfyLMlvBafnaIag2Ic1LgL6z4dzs1V3j+t7YwXB7FxINBjQ++lKpD3T3E7
QO5C5IgiEJLzSX0VKqm0c689uVGkojGg1DZ0kXaxYCtraXgM8XwUY5RyBHOLjX43
z5TsQJPALTnKY1rkzytYGtdWKOPd74p3f99xKeESn4aFXmQxl59/fJm+BE3SJr/K
rDyheLfer7qvmIaztP5BTcaHjC5RG1kGaL5+1oS/r9W8z1lu4crz5l1vMPYwa+D8
Nd5y/xcy9n1xrh133kh7gwkFa/7kZkMBsrE8JSSfPT9PKvat0dh9yG+pLMEZ87vn
n/1L5Ce+rjibtMR1RJTk+Uos404jhswbU7rH2cPCzseELcR2I+NrDkdJTrS6u7WI
SoqChHdeYqp+sxIworJYye2ld5DI1Yf5d1u6gKOIYCU5B8fZtdqcYi6ovf6yAb5+
1Fm2NR4BLEdfrsPmJJJbVbrqZ+iyhb45an+YaxBWziycAESrBpHOpzopLaPdQQUu
5qsjDShifeqiHIGP+fvW7ZqEjBbibBc0ucTuXZwZbOCDL1IkqITulNHs5iI/Byio
CFxu1VamjsOnqg7h4dyY+AfVyAx8GTlh30MB/aGguNblm3JujVSelHR7p2SbyhtX
Ko8pOsefovkW5sWxRxwv0Bof4k+N5Iqaofyw0L7TLjo=
`pragma protect end_protected
