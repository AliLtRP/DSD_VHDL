// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:38 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
SmE/xgD8SJ7gzGBqSOFRe4jjUTFSCEtG/7jDQzlULb9BqeGG2R9E2e/pQ9QT3gR9
sHsHaOzdfT9hgNdTcUxMfAw8XzPEXhG4PS3AGpL8dGziDyI5h58tpLS0Mwc1ZpL5
4U4+mNHEfIB6cP15exZzUx44RHv27My4Xhix5VdrKG8=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 13056)
MwvMzTvN6iNczA+4CbEmi4InJUmeOk9F5d1nypIKVV56PmBufCL1WLifhSr+YoSX
0oD/lmbT+MpIapqyThVZ1hbgQ0THRCytFp858B56G611TwqkyBVb7p8QrRr0KzMR
iEE0pf6kcd1W86mc0xckUGmKP7CzKjxxCbUMl9zprKxd1VBLa3OBlVC/U8D1M7sa
Vu2EAybWHHRp+mZD8oz3gZBKqNw0bgZti8mgG/FlpOfPHATFDT0aVLUPJPP7Nk3K
lqJeuGCyBvI7x7p/al0B6D00vf/mOrBlJ2QdQmmw01sMJFbzaPBVOTf+/UO6tbq/
Q733ef42gAOqRwRff7v1Kz/Vu22GkvqDiv80MoICVRtkx/Z5ca5Ci2eDvzB/sKan
Hi58n1Gz4K2xZDfyZ8e/La1o+qBZOx67RQmG4yxfVEYteqpa9SjZfL9MLVW8UnAP
i4RK65c65W1QqQZx6To45TNuv/8ALeS7SmUSjke7O1k/mS49x7JZPDwUM8rZt94O
5AvShHvGnyrJQjJnkM+c7ry9Eol4rkM/FIcK9hpfrhHAtDqfqX4D1RnnlFNCHBjr
GMoXa5NYDQwFZRSX5Or0TSTQ1sdOqwPIKF7vA9iqchiouTzptUYIFmzPsY80AJ95
Q1PqLDgJPdeUYRWAYda9oBd11CV77G/Yp4qyGC/OA30T4ws8TXOoKfkKdR78WIwU
oSj38QLqct1hhGE1Gj8BypGFwYhiqnDKAaKNDj5Du4QQnDVVprtnMac0c2JwMPTX
iirhWrgEES9RZKeTrzLRVS4GVq1vEPO5+hhehMtutM+mWFN/sb8HzunkuvQ8PX6O
/+QAOetd+g1LhaVhndjqjPQqIczIoV7RV86/s8OpRgnOSPXnsPMxOvQ7iuuQs4e5
rT3nnpHJRqqCJiEj3KflNVBzzMUXRCadHAaLxzSySFAQGhgnQokqew5k3saKwlrL
cFL30/Kv9GDynfQFnZaIvUP1p6AOpafLsl/SyWTsm243TGOhyeHMNn0RwfsXLYMh
y7XM79O7/QD7nX4y09wBCyCtg9lr3E5LJs5Josh8UVnI3/BlYW3VBUbqPq0+vrFV
JO2gOLk7iAZIOfE3C51VqFvirY8SZrnFv+dkMTqAKR5kPrM1LWeXeX5GW95LAPvZ
9DUrBKhQpft1dUZDpPOyN2/Zg7VmIIvvZzoqcgw4sW7G/5NX+8mthSjWuhuQva/u
oIyf9i+VKHaYJ8RgVicxfPmv0PxSK7oje0IFD8duffr3+kM/17bUpq3U12dkLVSz
U7l3kraHOzNCtD9tQ1ARUwgNbxbvTeq+BEeyWXeHsFfn/5/iD1CStA7PhpUbEynd
UQ14gOyfKtBtGZzv20gG8oJNko5R2bo0DFQGYT0aiSSeEXnjIHMhpb2OgbzUP2fs
E2eHS5TmxANe6XptFclUf+Wpa9PBl/vCC21j//kCFs7ppapC4w7j28N9Ct2wJlom
MMyf4DvV171im1KhtLFnKG2a6acPQ7EyibqXTzBT41pvAwzQnggbjVFzcS8fFOHP
TugUaVV8Rj3v67ZlywunlNEHy//2Tfqm7H2+9v+y5pTDdlmlc+CumTiY8NUgznv2
GXaYydiwCaXfR+dYyP7euI/3K5AJg9sCFU41hChTYiXuuvenMmMJyBP1QU/wXcKw
YNvYMes8gh5GZSW2mrNPxIjfXa7sGSLqIL/0rN0BnI1lufExw/iGjTHsGgwnEy40
Z1YVdAyA345d4VgHT0inuUFUU0W574uU6sKAa6zJiqNfpQA7jw582JTIXQ1+cc9x
zdqTD7zr340qRm9Mif6ZCyT6wTKwy9bE+SK5qGE2JEztFHkohNbhS0Vp5HkagpmX
Chf3le/3xD8gZlvV+ANvzZNFheeZAmtZEr7WVJn8wNZSgLiu+XuRkGT7+e0m9P+O
rxPB8K4UDIh5ZBFaAzA/oI3iKgCNDsiXgcmdIbHUv3RlJXbcE0Xf+PV7n80UGrCP
okB5lwKGttxYFbrHaJflMdoMCzhWGwgJrouauH1FfopG+XZ5SbTsC0QX/8jQ6Uxq
TgJ7c8/pyFeodCEJoiEFd1sy+tIgcNvx1h0VYCpGyzahlH5zuNZOpx58RrNx9pkr
pWYmPSrSCB/upX8eehJAdE/gHH0GZ0mCu3+CJa44YhZ567Bs1//S71ONo1R9Njre
w9X8wI6aFMurLNkNLDi4DGfu0jLbP2IN5zw+qSI8Fi8NUKY88m0rHHXZl0+ZBK8c
BeoSEp7zA3jWhTx9FUai9iadxmsL5jzWMD/mE527Ex0p3Vioyi6h/jS8fKTiQYcW
D3PTJ9/q334I22WV1lhBzwNY3fdSVqSf6ftDxmXbrNIZzy6tshVSdEcCqCyM01J5
DdLq5DMVpS4zvIIMeQBK8FK9BsWyRK4RklWrn5jW/DUy/WiJq1AE2706riaFv6kB
a/fpI5c9QD1L1hj4w6d9rBvZsA3kAEcJlFB2WoxhTFtq5hCka0p9bEeJ++QCsICi
M43r8NQ+6aS5vl4SYpmdJretyrei+F8ZbrXDEXW+H+kW6URJogtwkBnpXTz6xONq
EX5tqonwkr67rvnTGTISg6iHheN7QOzAiCQW+jDVWlIgeG3pX2bzapV46cu+MEMz
9mXiWTrs5fIJ/8MZq0gwvHuLdAIfet7BIxcbyHwYH0FsSKPPdt4TNbdqrMMcZmkP
eM5EP3NzS6wELrpCspk00+hSkSDxMRLQhSH32u3evjyMwbXqqz8OgPVUt75Moguo
ldpa098ucaOZE1SlweSYc/6yJ6iLEQUCbD60+lHvdvi9EYVlxWa8DZC7Bn71BhcZ
OOTbmRkBmkigzNl2dRx/H1Ea7S5rjgMA5JarphrJjjYnhUlRVnD40laWOvR+FvOg
DF3PHijEqiMQZ1tQjiDuie+0AThyxQ/2plLuqFh8qG8JcpM3WmbGcya2rCdoWCB3
cjb80TXu/d87e1c8IRyzYyzDZqkleJNT849xJWbPIFb6yprXMsC9bbgPakTWmEWO
jPVIqIQ9Q/ISlRRmqLY+3ixG7sEp651JcgKzu2dLNRQ4yLgnT69sMilGaLAwduqn
H1+LEHgkx/GBJFvI9XgmEiKWKZOdhDCDMpQWc+v3wzHeXZ0UvtEkFB/yhllPKPxF
1s50z66AHX/x26iQRpgah+HNPY+suWIXgFWJ5LTiuOfWEO31zNsARR8E7YrYAPwL
IxGYL79+DDBnSNZkZobRbY5ZSeG1WHmYmPOSbwxLouHx5SIuCrU2vL46OmjVPfzH
iue57cj6LNvF+1v753Ghx5T5V1qAHSwjEJ7jh4vGNninDaR/MYmtaVDb7UUHytKI
yWMvaQUPR2+v/+y+jFG7m3vFd4J5HBGqTXoXWCKU+9299In7svQcOYJv6hqHf0I1
aXz7Oc04++zU9kWyGBFzNIeyNyspTT5/wVYDqsXkDMnt0NzeEjW5bhWaugx8OaaX
kSvfNKHHKhZdOfUL0naUyn0SGCLj4DI1+C1SmghI9Pmc4HJW2UJtQztRXp45CRSO
8k5v7zXrGWYm0l7OdySPJxbaOXRljGD/JyfeCdmIOLENijLo/JS/mWuPuqgJ1ooE
UHGSulyewLqxCh9a3lcDqcm4BtgdK7EqYy+ftl6WvefarUhncgfTW3PnxTdFyZ7b
Nz9I2g2jaj02l1JAK94suekFDBU5eAsnrZFTuJU9O/OefWrK+8bMIlqTSb2FAfUP
PRcrwjYdnSzJRYiFicp7aPKdflsthIeni27ThDsPZlYk3QTzPYP4SM4cRuqR1u50
JRNoJ4PYV+Yt48uRSIwpQizjpeLH2bxP9MwJ8p8nxl42y4Gf5mYTLnX33iFPwsj8
0+C8rZiWQ9FH1u24MjUERMNM04DFUKtNAViIwwteQP1djVoaNBLDaRba27Pi2Urr
yxv2aTZk/OawByv1iDdebH+/D7W+GJbrTJh53MsIeBnFuh9a/yF/53cMfvB5VX0T
EwC9KImj4/qL5m7E2RTGH3ONs44qlhUBi/av9ajxc2WfHE6G8FSfs6R7DgIN/LBZ
j8VTN/G1PpcSH9sEJWm5GfBY0SskKQTpnMDuk4ClhMiD/XKnc2eYJ7fUHt0F1qfC
B6TdIXhIVyA4W6qC7b4I78xzYzaTXMZjOOal2H1RGw00cHHPdf/KPiZSdQ+0xAFr
TtMMSxrc9TWGpfhkLJqhzQw0mE5dEoOfkpRuoMzwk6UjpXgHkGzjDknxkMPKMCsp
3cCclBYOURjeVRyrUUp/L1zVufTwaxjqLBgCpD/cNH19noDYPIgn1wykFKupMlcd
BbwLSSyaR4I6kxLOqQ+nNDu3/fhGN8M04nUutcnOBhUFSxnv8EWokiRVt1qQw1f7
5YBBcu68spwHClYj+MdkI/T8w4UMHiUcLkwUs/NKqUcOS9J6JZ2sgYssxqWGqwzn
haAHFtArFkOqBCfEDyYDFVll3Mixr7Tjj6tTL5wUVHZfswPr/3ZnweJZEEzoc1C4
XOWeIR6+ZXtyotQ7C9PmJ9AyyU/V1FI6U+K65mJ54BZTVgI5bOA9EbEc+F//dsRy
N1ezIDLCEg1zZF9c7jx5aCVbGWp47dSN/EL+S1CFRBjfyC6id+dq/VJndwed2QGj
DEv10hvwFaTeBaaIfjyir/iCdEiDQvMal4zhW2670IkgxeKdN7lrjP9LN2YYJXSe
ty683+D/NZ8C8kmpAYPf6x4ePxXL1VnmDGXs+z5nnalwWBFCRdQ+W+Y3i72Jmdpk
sRddWHeG0TnzF0K9CirWsKqDBYPUbWKUFfEwUt0nTjRvM8ugR+shZmjNO/caexa7
NY67mN19dy1Ec9P4GMVwCkR5JBMEkZ5XcRHicflHccPtbr2xkpM05evN2GAboVZE
0xHL1bvlaqcwTw8qMioAAQZTcnIFSH3/9+UupA+/k/ttrmX7f26qOEAAxZByQTIH
ov2EP0AZacBSGiXEtWpEg3k9p0YVtIUx3nzas0XKFpOXuBaGSodKTTarEsSbizp1
xnXLC2xyfAYyhhWfAhbYXtKuki/Dwp9AttAG6iEpc/bXkwABaVzq7vnuQz8g7PWI
4GVCSv8hpXXf5NyBM9Jqx0znkYFMnvQEKPzCHer/GSBc7KDS85C1mv1OPsgS0ToO
ppH20gl9hiBZpHOwFV25cuAwentervU7z+Zt42Ys0fPawTIwLulUSvpB7hfTit8V
Gi+ej3gr8fUSCI8ClDg34qHZ0ha+bz3mnG1o595VMmLLjFGmI0M1Eje6PNpaikXa
84nI/PYTEO9fx/+LINCfirLuUeP8iFOUFa9YhMePNfxoxu1XMZ5R14j8aFDXoj16
Vhkmlk/OGDLy4ezJvY2c6t8OCy3F5aD+Yqm/D+hqKMXu6oLA4dyrABuB6HKo4crS
vK38M1i8EQLCMj4qxY0c9XhUNgFox27M/q35SRK8jE4cz4uAelhwDlrDAZe9Mqwr
L6px+pdjX4AR0bfObL98+EGwqUEu6RfU028B7ukn6Qua/j103JkdiXz2gA+6SWkl
G0YCH3anPU7jETSOyUCirbC0ea1ljSKuTrSKVNUM9J5KsOmd7UgpIy1ecx0xOyLy
BAbAG9octLjIBQNGhOn27w2lMKmD90DqnaQONpJpiI1xx5atJTllPLEUfVOnQEkU
uhOLla4nLhSpVOP6oruq+6u/En/qmfsG9B3eiSEcexJf9/KOMFmopu+0vcNmjw/Z
T7yaCGnWHe6/p9QQ0SLyX1P5Dd90bfPrVbA5QjoxJ0WW5vcYRDq0+dz/C7vX0Pfr
sekExarm+RShFr93YJTBCP+RwDecraRkxhO9FLUtcB3n8Gw8Bx/x97AZTsd6CP/7
RBHGCGfV50Hvl2Veb5LVUDQe5XYKNA8mDap7Vx/w2ZGzm6ItELfPSoLOwoWoj2ny
uyQrroswGJ39O71Z+g+u9lualOPnK8M0+4fTYYdYAzNcIdKSPnOp1Qm2vZwVq0L0
k1s9Al0IeKxn5FnTyEwevs5ZoahqyX4hAtGXylInvKzVadClcdEl3lfv5vflDYv0
SFb+9fG/awydVAMRntGdOaF0iOBOvK7vHkurt41mA1zVmPbK/mSPVmuAL46Rqk+K
IR04qxjW4BAYP8Jidm39JXojR2T6l/K8vQpC8bwgVHJwJ5iI7c3MCjWjwfUl63P/
eIIBiw+ESV6LheMR+wIwZsdduktc91dE01ww5wrGfhoI/zvqgsBaTB+g3OgbJJ+E
hE8JQDw7nFPobqARpowrtPSAxc8uoKC+upYB6tjwOZ1kY7kMTYiQAokzkkc+/Ge3
1LJ4DwxCCldMgF9pp2ufET3XW7BfKHZSvyPvr+AJ5nuZyIXKFJ6FCj3nbL5G8mUq
EdbfYBsY9DkYdxLwRNcy6R5FpjDYpSQIKH1KBej7TeIjTlSOQVwrhoQB0L2n8yXW
tV1UdE/KV47Mq3CCCs6B9hnzdepnNL8TnF9MJ5EyKyFKLU9t+XTavp+fOzKae3XY
AfyJPrptD4gwvoieKsPNQVfeUxI84H5T4v5OlUrWo3b9RmfaZuMu1PSkkKpF7/d0
eqcLzDUhPCFCd1JCRmKtxnrunpoVe1UkvDm7WscUYRr9cG5tObxwQCYV+yqDg71k
7D8YbhOS1vAmuu2nMUY35XeYMop+3OgEY39gx6RqjUsHlTL7K0E6UrJCZIJv8Svp
8ddPFmYbSdDacF+3M+D8eo/edSnyfclcc5eH5Q6e0dnI4tWUM90PNe3GDEGlfxHa
t1Lfboe82qgnd+7I0qV5Vyhz4rpuZi3c+7UKaCZfKD8JoyRxUN3dyn5G5YKy+P0E
3vgdJiTrNqVX1Uc4zN7Xpyrc53Hmq1m/bm7hQDj43HBaeM/dfA2Y8RnF/6AJxdV4
Hl5ZC7c7Et64GYc731XtkM29ylUuu03RmnSRVUN03svVd18B/bA+IMnT4dPXmo7t
NdWvpgINtig5CE54Kp6C69wMLitdag+AZ4/WhR96TS/TF1qdvAwjt/zSxHVUxZ4j
HWwpqNiJ/foUHdyTPYOcb/C/4zPoCKXxiBcxGpc6GKv0QMcdvsf1ukvwUCWCuWqF
Hh10yCzNmktg07v3c3KXuvNfQ8XqbinVybXaaWUVslhTBYDN58AYahS79iFVvyfM
uysg7RxTmhkq8iYI98M9o/ktp5WTSOiSio8985NTxju63nHIV8LHD1WbpTNeRuFN
8121PhLN/DlvMcR2SY5Rt79Tn4sabj54crcQ2/0RCaZuX3LJv8rIwkjMSfznhJfc
Zv5h6beNXshb2chsiow+AzCV2yU/rrJltr8Z1XXnbrmRBrO2wFhXUjBNEPTUIXlt
DHH3WBVSbTZod+Je/6tZJ2RaoBLrL8tG1Xt9H/toDtlkkSkXfls9+CzwMdNu8BRY
G1JSc6T2QBDqEHE7yaXFMJC/ia+UxltDnJPS7XuC4kLzqoF2BJotStqugVCH7byc
cBtmo5X99Q0LX+XkVe2WRrnbJYbR+VWOwFx67qomaSuntgHmJ9dV269w0lfA9mcJ
REEEXkaiUeeOCJmx7lVTPnCSsVSsPAxKSxPmK3PbdtSOE1+bK6wcRopGMgK8whj5
r5V/6e9ap1mVN3BZY3SrdW4/WQpdCDLcUFwZnbdp06VtmPzkiaNv0nmGb1Ru90XD
u4SSxXU59EExmLQaLNFjKiLtbZcjWadN1KZKMF6tb7PmN5lepWqfDcVbIp+ZbfvA
BIvIWz3HFeMY4QtEmYeNP670MjRrUEbxdYiA6S6+5Ngv9NMrgt4D6QI6h7dWVNVz
IBEDBk3lyPHClkWl9YlP4fqDxksDuU9mqiZvzsr0EdTdLBbupNEwSUNcMtG45F5z
pEvcoZa0EA4uNZmMDdj5nSIJ1uXLKvm8WaW0CfieWQjjcX4pawlV9sDsB0DuSFiY
27U0hUulg8NTiBpZvHRXCxaHj/gisoN8scyMyl6fPzIqGfFucJjVji+4QC/cYidt
9cXsJt9OBmmQoyWjdm82kuceftRM7VKzZXd30ibPlsZstiAOnrWkKSpnATMKjjk8
yWLQVnTbY9WsVKS+Rt7SnNYttwKHu3iwUI2QXT7Y+sGYz3KzYc+j3wLnEAVEUNTz
L2XjRyegWECYoX5/h/gjPUFz99fb0E1AVRGvH5EHxQji7Z+s2nWj5hugjcS06TyD
vriG/Kh0jBX7dqzK0DkWAswxgHRwd8GhnglFmpC9AUOH+Gp+LQ6QkhKQeYqlFnjF
nJwHIhDzZyOY7DFykaHtu2cVkY2lE0CGeZ7EKPmfyPVx7G4NDJ1oAYz1LW1bf7yR
I+gsDjnDXCsnDlPDDSz4+8pqN0NIP1cnLOsnib2c2OsyBAuwKvpn07fWj+K2XYFA
E6FJjRuk7tOalYVqtFfX4IWrXK94KsMlAavE18lTLDG2cRHGogo6DeTw31lAn315
UU4fpEeifmBPK6PxJRNVck1KNuQRBRg5DaXZk46pbAOzq16l5HeRFK8KwnlTkOdM
UkAxIGUBsNw6JbJ7HjfLfsTBHKCOPXz8KmsFMbZGvd2BmPCsTEGXzsALW/Qj7H6p
NGH3KeFZ8JkTusFGLvnjvQRuCgsutTUnzj6j0zs18jmgLxDjSSjQT5lN3K6gQW4H
/foA2fwagU+R0psh+cUBhVvtSPEiAxz0jVQ2moGhF2SqNM/LUO2bdw3VCUbKs2/2
DyXhiKM7vPOLxhumn7o/nk+frY/7hGM/bBx7zL7AAlvqSWwpiVqKNNKnkj49MZSg
Yp7dI79HTnLWhfFyO7dWpJk5fsmRwfB/ik+R/uWZiaKLDIsfO02pqn3DYhdo4S3X
vyAER8WC5yxUrkT6LsOYMwLcqoED9quaf2EczqWQKWsibh8CYvimKuG5L9neJ3x4
7gz8EfdzwMryLWNp+jqibj6zJs6fMOXG2VxCi13X2CTkgRbeLaW8bKWNGRA34Oev
Yq91hqtbojfApLC81RMIsVKw5gAP83ws2yMD3J9fwloe4Ux77THA664vJ+h1NKD9
aNE6qkRssvEUrWNcY2l6GDZNT80VcDak6sQTTvRfT066h9iJvScZ7KWs4o76zo5h
s1f+Nf3Y2c9vq5yQW7YKzHtkT/5hi2OofQFqwk+gggMadvimovfAu9JP5zJE/fAL
/cWLg7fR1NKqrp1UKHRPOJy2L/7LT1pC56O1oo6sLQM9sp2Asa5VQK06GPVAL1yh
OPCtTAljWB2uR8tnkQMxF1mH4X5SggRP8A09YWGA8PwdhtEAxpdd2axC1i/vxoUs
9QKdPiZWUbgS7gf4ptZMn+0SeF3lyFEn2F31uoC/L9u9s5/ML8/GSZ/glvaNQNlR
uQSVu6G3VtA0zepzgVygkflBJ2SabZ2PDiUyCpesHMaRtW7saj74xcVOZZOLoLl5
T5ylBK2CPbUwLUO2N+aSw1u7+cwOhwU94L9s/NTJr9ZHZRNabDk97YXLtfjK1uKI
GFLH1uL8KJqVeqS6pHUwYIBpuNVOqESylc7E8A28i5jpPjRaJVNppaBAjZHJjf9k
wj8jSaCLNwRj7ZW4iKOaJmzGnKZnBFtZku/P/ppyThbAuj1dgto9zFdIPB6Zz7QE
4dnxdSqE3mNEcnizajSdJwpQg/CeHm7JmsCZvys5neG03ohqOao0Gy8rkIwMrZhG
5Ol69mq+dZvDMxZUpIM8TDVGiypXXSmzt+tXJSOk8tJYNNFy7juaIJybR65YraFX
cFT+V2UoE8zLj7Z4cb9xubsfVFAUhf88A5Oym2QylPZ3B9uzZmPgs2wdXTHPh3k8
Ps16dfly1nrQ3T06sxeTDk1VRIg7rdXfb8IOA5vWyVDd08OjPl6BmdV7fYkDwjlp
jW+RpEKJbMgvht65BBNjOJRls8HyzgWCgVwK9hilxQ1K1xByflccrvBgLsdM0+4N
h79am0x9LaPkObiY1I4BqHbaO4xESDrk1IGS5kAxI3KvuOOvRc7q4P3Ky8YGs59d
GkpqpqaZ7fRF6z+Vo0cXR5VW/uWvkVYbGbFlyHNn/SxBQZl8vr+ON1YM4FJkSxNr
zutbi+PLnA4aBlSbb70V/4TbUxLgWIxmhIM28J74jyUO37UYvj5z8nhx5MNwRBid
9CN3opdCgNp+h2TRItL17AyJBWW8mZTNMC3KNpMS59rBYI2NNreUY3LEYObXmLvx
C013XFRRCAlae/kkzueEEfirIvhK7orxpVQxDI+3+mKpKTJlfu6LzSYsx3rqqfOr
VwZ94Fo1QTwK7lGfkkuN2NlraYK/+WZW8IeBZhKuMaD5IKK3mbKeMPoV1oDQ4bhV
9NIiU4mYRIyV/O6P4N67cY6W1gsdIUybLwWPKFcDYNbxnkP98a8q4stSxzw/k9SU
cCEJ05dHcQjy9/glW6GoIVwMfNRPeRuKAJdNyI/Phvg3xraeSGceyXgqFGyrL4Bb
PN9YU1eqCmuz1xdQTqseTYZWyZV1lQ0MTTg8BqqU2gSy0hK1p+AePBmg46cAeCAl
C09sKeRWHQsC62ow+R8FPGVYmDDC6kZkwl0tcVzRnHBa+43eAoqAUG6CjP7Xhp7R
Mu8uJBdOpI4MPWxfH6A5k8+V/zMMfvB/BLA+Z+Y7r8k0Dy/KSGbmF0MPftHiADKE
k1iLf/Xyuo4ogTnt2j3tQH6fYZbmep1x6O7LFmfLDlqqtFI/9Ry+obCOiDg+95VR
PcFl6P8pUm7LZNLEbG2SA9NFR7G4QGGfFC7dLA2MV+VgB1McrfOS5I0ccIfKZWky
kCSpDjK1PYcjTIRCpH5oCUFs2nhD/Xm2sPO3dsG0eBbELARBQxoRjc9bJq8BcuYJ
Wt1I6AfEIkc38HEEF7pRN9u33sPuL+Q5LI0KOWmp3v2uT0Yaf87TD4OPJe4LwdiP
TGkdNOgMH8miNYNOBCbnaUFY5tBEpqeIL5mRPDNc00I/ArTP07NwSxnHDpo4EJUU
6kij1VvMlbcqrmWbjXogyBGmcpWpiFS8yAnhMAdP90dsckR/9yAl4cUbvwQoBSeA
yc6g3Na+oPGhoGa5yH1VCUwyAeOG0gU2hTKFY8NqBxWrwUsoSS1v+kq+Qd4tYUt3
AwvjWSFRxygzXN2TbHx1FIJaoc5RNxtDMH7PgqsV+hbNR8Ku46NtVNidc5sRv5eX
0xqNLYUG6RKnobq054IlZhIKLC3K0I8MYIc8ltPrP/QHjojvlNhUKfvtg4av28PD
R2p0K/DQayIyPbZW/QkgNLPyb3AT+PXYVR3HixUimkWWr9NvqZQyvJ0txwLSOOye
3vX28vU7+Y4MM9jhLHx/ORacEbJoEWtQ4YLcytUNiH1tGfDC9yz7b+8c8yyEvjn6
+2p+Ej/8AoIIjxdoLzZ+P40E+mpcO3Og15z9ORe3/zTGrLEIzO9iCHWQN/akzzTP
95X7X0BvQJr5KGNtBRRsG1+3AQopViEoq3jXpvZva7rtkrRctjId1d7VMP96IsTD
v0F0Xqzpa8Mj+Xy+6Kwxg4/sAMWJR9bBHp7FWIKKUt+aTWMBlTresaN21OY9YXd3
o9aOwJddwUmsKvfIsNdFfetKcjIueatimbox+fvNPdrcVDlyffz4MZ/cn0RwA7LI
XCMZrM/ggQWXYxacMAr9r6QgunN9/AIoJb+PRZau69SZ4nbuMx3SvDz7eI9y4Iie
cJC/NIOV/JBy7LcaZu2qV6yZ3SoiI/DsMrH0/DT0b6T/CtRxl4BC6dV3fiW6FWHK
XaGvQnY8ofAZoVB46HodNPr3+IWp4uULbUUpSWeEL3Twmld8mOYoiOzJe097r+go
TjVh1LjH5wc9Rhxw3DOOvuk/8fNfU2I26At29S++hy8lVuEZA6V8dYxNoerMQjI2
EaALwZW06WyfQIzJL0uS7jObTCn6dOmLiwEWY31Fz8KByq1Nphb0vQajAoo8tpDO
FTJTiqkAlqSNJgye6ES394NPtvmJCrilj8KyyKwBJRkLbX6uv0zU4qH0xfbnutBs
ZI85DazyQQRf2efFAj1QiQV8YiXKWI7DhIUwi+YKXYGB4M+juujEPXbzlg71W4Ix
hhEGIYp52qDHSKyIpIVhXDzSLUdytB3gTjqlXcNrsL9uMH4Gx5ZWZQw4WdouRi0G
qyF0Q2pTXi/fVncpFXgGqdTZ1mbIriNmkMY3W7VaVByZ9blpsUsGyfqGamdzH7LX
a6ANj99/XSeOD61M1RZNJ8SDx5vdhPYjTL2ZmF8CaJIpl90MbaewcMTl+R7V/Q8j
UxaGlwd1l5ZeIw5YIHy4DhhigzdbvMfEsTQQ+0TXwrBQXTvrsiRmr7Q2k9hf609w
gVS66wqYUhiKFrDbGbVRjXxXwgTorFSlOrLUYTzHX9Ts7fUpcKB+A249HDv406cj
zUX0Ysrl4OjSFWkD5JnEYq4HU68NC7UwXcUSruL4r2QemMBdwIpaNhsafvSFBeC3
zhtwPe306n/qjGfvWiqPFWqEQjDIrKjx0JcYRWBP+LhQutc3YyNSUk8GNPsvTt/Z
pIi9OKt/02yW8ex/JFqpZSKcfRsNa627mSgftDfcv3x0p+2xwHs06aEJ+McDIh/j
4cIggibWFoKTL1Cs9jVbOyN9lnMJ3J/kf9LKZKKihLlJjL7CcvIYSebewAHw7Vq2
CNq7doJSnnBCkn92wQXCG1NOAwqaAKtL8E1mBDr6Tw2sUQXw+PPsnqr5SN6nngbY
YJieew58BtwRykTfl6Cw3O+QK/dGPakKrST0BJqCGQB5SFnCEhMfF9LBlidcr5j9
tOsOQpAMp4JXQRG4MQIdREk4kBFmJA0tmIoebwLEXEaiMAXgun4ecfw85cDhRVxN
FpDksU8879QfgqqBlhvn2a+TL6xsCOczsbSo+Cd7Ps0cLRlX/R8oBrHNZAMNoii1
ZwdTSIpvZ81jgQoo4bZzuvZVWrkrD/YggSTPLibO9muu/1dpIumraooOl0BhBTY8
+q9S1H0tF5BxJG7nNASss/Y2He1M0gHLRHJ1I6WpwhT50qI2v22EPPs8aWSWWtgm
kV/g35dBNCQLJ7jitbqi7WFHZcyQ0xtYNpkT8RcMEIMDXCWbu0MTrWKHjMpxYpA1
3HCJurK0QPXf6ra31CbmxkAg28TKEzVdUyG53O5q/9lIqsZjQ4N7yBM4zw751tXh
1sWGfznBnduipYLLf+Re9I5FYLJ+JsuRY5j3yuUWZu82wmz+EWfgy2kvDMQf44c/
WUYLWBao8rQg4cXIE5o6o5Db937HC7Bmbhc/CJjv23YjOoSbnshaEf3qqAZSKm6P
vSO+iUyggJr+WEjwefWdNZj1b/qq7CFKoA5c4ytgxYlcHVo3l5unHpDyndhVBN7t
69kdY1mOCImeuO5mn7tVN2I1d2jysPTqxY/R2JM4USycYs6NFHix2F/yif7RaeTV
Vu0zG4mWg47gsZzLigGOwunzNcG1jQ9OZuFl+kK0FFpouz1ykul5ggEnN8nMLPFy
v/Gx0gGWCNkgaNNe0PBrxx2RS6IZekR0Mm7nsjaozDdEb2X6GwrtifpIme4tWmxC
J1ayYhqF9V7aRYPKQQ2gDuzPYcF7InQjz8PlilndxiQXoE52ljE0KqPwSkLq1BUh
n5AHmZdF0MTVma3vC5aDMiMj1H8s5ken0iCoXRSHDX+wuMffZH/pcgtgDIOFqvfg
1EC0xSRBuU2TBu+EDeiecJ81eBZIcNIt82DCj+HZiPEMJxDIyyNW+Ahp9RTw+QKO
OC4Lu7sdjvcPpKQKe6BQwbZw1BSE+ygyHo4k2lc48I/ivb1d93L9o2nym/QDhijx
ktOBl7hAt4nfuqfYUmyP78yRgPZf3aU9mcTNSwgn94II630hyZF+kp8rk+DuYBvG
u3B0ShZlX62GVp15+tzv8chaKl2UnCdM8/kCBdH4J6um0NnYS6H2MKuZY0S+dHaP
wdXtfjqGZbcv/SXg16EzPmmfa4K1DBPj9mfl0OK+YrPi1q7pgWHX9RU6ORVs0Fg3
OpWEzBfutXu3s35d2suyWImhf5Jindd9nauO0xHYf5fp18BZtuw4oPtFCfcfJKx2
KwrHr8yddDvDQtpOmb8IugpeawiZt0sQayBuYWQbYYdG1i1Mvs/tZRG1NjTwfVrx
RREQ/4SzQbxHPDmfGBgIrbza+VJnol8RXiN0FUIkkluYsS8MB9wwI2dEyOcGb1PU
TwYrMjmLE6eZnE4Gs74SvSlSM0iKepZyRpKju5BPx5NZnK6EVyYnImWY05WVXaI0
OIFQ1VDIEplcNKgf3jcrnqphtCDm5EhF/t5RQqTxfuInfaxyoHlxAc44MqU3YiJQ
qpjjoLES55ARfej0XGYiXNC4yYBCcEJ0VVKQhUA8WEuB0hvbjLDDccNes5wwPE1V
5dlmHXqGzqeCGDh6Qhj1DFmZdzAj7Vc6mFLLny9vqYfC+B3dOBCEtyuPWV3x3sdr
AcstufU2hS2v0Puadk4nYGi9eClgzQpVDvTGxll5R3kehmFqp5si8Azhe2UfZLQK
ilQINHfGN4nyk7AhCiPoHPIMvb8Rua73uCl5PACcPh/LCANip4SsyNJIwEcK6vwM
uNan3/FKErlh1lv1AKx94su5xb9vGLtXgyOSY2Fzko7z2EmWogfa5JnDAAsll712
C9oI9VuEmMTt15fHu4Ov0L6SjpFtJGo9GcUBlUo3sgEHwwgXwxTz8AquTTB1Hf5S
ofsANWZ91bipygbtaQg0q97b0YgItbT8SHfZcb56BbNVDirXcVzM6rY9axz2DLlB
UmvXlanq9pXG+crFg8+VEywJy4DC1Gq0LWbQoYArRe6UASFVzy2wRKM5cQr7Swb4
Xcy17Q9Qvzxe5IHHJxNVWY5wKwDJpGk2vZl5jdbpogy0GFGaDB0HIYI92ajX4P03
OdJ+5MWYoscVo+iIRlpOAxarPPG+UfWQdm6oeeOmF58jf74CY+OmYW6QuzjXidvx
gZwszZDyRV5XBn/0Q0gSrabjiDyRMJNqBfQUA7AoMWV2/zPmgO14XlwCP/PMmkBA
bOE8TAEXAaVcI4LQXI3euki8O2GrYSh0mCUUwPbCYI0f7X2PtVCtv/Z+OOWXHrk+
zA24Tt0zhnuqsFyHgruYhLe0Cvs1351ajZ4yRsqG19rd2leQ5ngUV/a2LLjoYu/C
tH5iz+3u/Khr+1r7AnNYUaxZ5xLS4vvW/bwmuthpfQjAaZJClr/JsLNQpYjDs17j
iBghTqr0adY5pnne7mGyOJcLebqqdpHK3M+hdCZEazMfnPMfVJctm8BI4NiC0oUj
Jir91S6mpBvxChLCj2khsnSj6pKbYN29LWMIdFxNjbezRIsdDe2/Ac5POu0UXMUk
TTdXE++ZqlDQQB1xMDsdGZx37tOB3T9s3KHTTVxdNq91/8OzJTROujuEMroUaSVt
03qpnGmNVv55Ot8iZTKz6JoLNFrfUyDZbCtIt8H14sYAN2ocsuaHErZsQF6EgHBi
VObm3kpToOT1+Gsy+5zK4JOOQbAeDs7aJEyPHFIQUSRKX8qWP9QZPEzrfe/yGko7
ZwvJLq8co3t+vzikIIXU5E6sJK4PW6XlWUHve3jV4E4zrrH4LLWu88BJv4zFfU9o
ZduwzUb0sZgC4fuq5kvlDVQoK+fgUxdYhKnbcrV/BNBbtVInvXP4jkTbr+fUuhup
tMZwnsnf2sJOMlvhS3u3a01zC1CXo/Q9F+n6F80LECdH5Y6ex8Dqgu9TtarFPcd5
uBTtSyB9pwb6VHYF/KYeL8dMadQG+stHxDOB6U1F2zOrXHrOqeBxymNqh7+0XFSG
cf82Z7++mNMfj5IPWCQf/SK9tERQ/NYZFnT/m1iw5JlRO9ntU8aJTaUwuthRtRCn
2WqAZSnpXRjyCRLk+GSTpxKR4+a+mA7tw2iURKrMx2WZosaQTf54tkNGsbM5nLQS
NJ3ehaqrsUbirsWN35pte27ZHxlE2qeo1flPJiMDtZTbc9Bafx+A1iPzZw49t3NH
C1dScioZ7K5/6pO08RzXvtEH8MzYHuq7ZFUsjE3YRh9xr092GTNjMtsadyFQqenn
mORuyIKnsORFpIWBErTFiYm1Uj0t68X1c+Z3sBEH2Kasr4bar6gc72RFEzw+Sq1v
UoMV2NAkb7KngfOF4PcWqUfE4bwG/AWDuZO3DjWyk/SZdO6f9tJwJLGLpcDim6hy
5X2r7WxsAUJKmrkGKj5fvhMH0MEsUfdhAh6MMAfpXUwayuPt8DbiyJHMerl1UJrS
PJZUFhXsal8i1hHEnYp8L6zBN+qXO0scQHR5N3xD1fzFcnftKy8d3+2NgRyQOe2a
qm+BMj/Y8NaTRItZuT0lqaZ/aM7H5Dt+7eD8axFRjoLoGjEEo4T3gp5GPlc/l0Kj
YeWri+dqDq5IQdu2CME3N3xSExAhSvbAxtJXgv0Jv4n5zcjtztR03SJO/o9uEfaL
/HV0QgqEdFTrzRPqHo3+AefvAuKFwhUTQMWqT0ux5pYuCrocNtn33lfaBaw0kjDs
31wAi/Hb6an4DZ048lChWAe4GOsY95Q68/WnX9TBxgEpNSqr92ozhgR3bCa0h3P7
Amt1/bp774DvgHYIDJErxeVhrKATpJbxalEHw9uHVFa0ej0IwjlMi7QmVkZ1w005
o+fCytGao9If+UiUHUH3z5PLcn0sgjxhb9JTQMvzMh2l3TKkXAbMrKGPZskL+1sK
uDTLQzMxwE4SmMK2E8Lo2UzBx7gNogtfnZE2LkdW9KCdnLE/LXTxf7yF0LPPwsve
3cZ7dauIrHGoFmiL8MrpMDClTvWwzQm7+tVOpYpr5DRR5VJHtcqkiANNcUcONR6E
FrCf7C1b+z+YeX4lh6nzviOft8reD+D7rXuuZ8cW2NJF1ird9N5+cvOnJNYXeRvl
OIa06v/B/fe84aLzLg4XFDtu4cI9JoodWGTCXJlYgmOn7SNrtcfoz40evLuJNow8
KEa9ILDC21sncmPKL99a3ZAJJiBG1Mr0VGGDdR9Pt5nHLUKvJjHoGyeCTuzAgfeB
0SR89TQP3QQscK10M+gIuOqYV+Twib4An19huVE89tLMawxpZNos/jIGDMd6QyRc
NT5crOKvEdteP0WBvmiuedJdigEQbvuc0jyUgJrn9VedyeQKqtomuJeDTamkqej0
UcUcSUcep4geYvZGtNF6FRWvkimy+p4YousrJU+TRiPzvNDkv5H1h1rOFfJHOlW0
AhvF92lfoOMU7twYVWfx7hfixCwOQgkdFFBYJYdAvZvvDWvXyhAKfS+Xnyp20fyV
nbl++N9RBqloGz86ldjGdw5zlEwLI2zPlsIAjLoOyDf6LVd5z8K3Jcr4lB7vxM6r
ufTHQts8jZgjQ36TM1fzCBjx4/GCJjE9RwmDDDZ3BgV+VdI0MH+Qkm1T76IJzIQ7
og9ZdLOML59PZCyo7HFa4Fyr1FuylD7NqyOlQC0ykC6V3oQhjUY3CADU/L1R5bTl
teoqf9xqoTlhE2Mh7i8Os4KP1EuxitBar0Cjzrj67hiOddgNl3v0NQpvxusGMqHX
`pragma protect end_protected
