// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:35:23 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
C258Jvcur8IoGsK6quyknXLXAqN7gUbihappfiHFxh5JVNPrpkAMzitxFHrCo6sy
NPfsQ+pPlECTzH+jbFBRIytnRmGve0nNSBicFrvQcV7CILpDxLFZpL8R8w2FVEnf
fOgePUFpSyLYP3NXVRWq8IiZz4Q19IFWJsq9LY/MYO8=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 8800)
3T6vMdbqnb+2y/NIfp+wAGg1U8fIkc+mfIEbxNvFzF248DAMdh4C6tNCwXr3qrf9
oM2rx/MmIWDRvvTlcBvcj156IYu7sfWKPvr1NDlZlT5Iax2FpPicMq715DdlCdFL
KoS4A0MIne8h9sqPffgHbeZTExfs6fSLb8Yep2I/AJiNUevU00H6Fre0YiH2vtfr
w+SPYioXCmnHLx90VFdZlhjycdydzqVPKH4umcrPh1xpZe8cBJyGX0Wxn+bjd5w5
lYyW5iQYfKA0L/yHHmZCE6dXbK81B1VRU26QtGiAR4eGxJ9a9ILalsQxhRRqtOKb
po5gStiEjxaLVfq/O15dyVQzbVE4/ongYBSp0WsD2L/LFnHNV0pEd29MKlSsN/hi
JJ73u+8lr70wiK4M//WUDHMvus0hEQ/JVnZPmGTcqYyu3VhmFwMc+RgAG4jn+QSo
/tG6qPGwt89TjooWDSaROL+r1uUywCZZ8F7x6eROw2N4bk8zCntDJ6Plca55exJ+
yR/gJKZbF8iqw4/5dXVIVIGJ+TmqZqyuB7LdQlJz5/3q/wPq5MFo0oSGVjGbfO/K
1LoygLAXAPGjLA/Pk/AOBrRTEPqLZbals18HNDZH5luy0t5mHERyobsDDFGxKILU
GmFzsOg13ntC0uAMOjsVyjSAbRODogMS98m7i0S2NZaX7rCffZKhTowlH5BIbqa3
lbaviU9zBm4d54asZ5yX0YPnru/khGRV5hmoHFzzm2U5sQZsbzIFDU5uJQXRFajC
3p2Rbj9Xyj3FKvOtTDZ8sBd3C7aElVSkJLF6M1XVdx1JAOqv504LRE4aZN1ae5qI
2+n0nXdN91aae+CRR/QgZ3DbwEh4l/5cgvOqoPM5hjHcsAkB9ORKkbBY1MLPtjTH
BrAAJpVIZMS99+khoAqnhR+3tiTqXd1S0GdnPezwSGVV2fkzuJBkUcWlOQqIgmSV
0BxrS1jC+fO2JbIyQlzdpVyla0yiuIQbTs8aYr/HaXnU/uSAmt8RS8PpWurRMQ2P
+l7qs4DSAIbuHwth7L5NE/hJHaQVbt+7Y5TqEUUQ/bEXJe/MPVrzlkaTPtZYNY19
tBLhuUB7aWAxNCcMuKn/2ZP5zffjJihcBvJiveTDa8ftgZN2BhvOhq+6drlfksyH
O4qulsIiQZHGGUVTA2eXEOCq7VvOE63rKLcZVD+cfPPUqe27UW6VJfBa8ZYN0F6h
3S5OlGGfEVboUtQFo+YTG37Yjq7yyNyEZjHbTSbsSWJCVox0AAsSAz4EF2abjVew
wPo61RZ4J5OX19D66aQVy/1bQTFLHC12C4/JVNDAUjdGOx57bdJJdxz4Ghtkb3tU
CnANKYQhb1/te8DVuj7KIQ9w5doHDDgDyIl5FdTnCSMriAKGPflj5pIRGj2DPGGe
u8Kc2L8vgN5/0ov/GdJIMntlGUCcGyxl/oVKBORPqgwrOg/Dz60xLRcfDpMEMWYW
Tw+aNTLze4XFdBwDWPfRVpiMgzj6eve6T7ZPbQNnF9BHJC2AVwexxH1eTbBCwxE4
3HeUsnrLWYLER8ChrYsmnp2FvjRg8HaCnbDgrt65PGGKerVyYJn8F9Dj1Mr29XoV
3PrU3+BQAZPPSXDRzaWRz/SCWhTv0VL8y4Ftdl351BvtUr9poNxOFlr6f3K2nWhu
e9UzkI2MaALwr3gCXf142VIyNEIl63KGA+3j3dbATANVnMARXQVi13zNZbHwCoLb
lX6u9PAZJBhQCufPwdAM5qgX0CpGZaZCiY1wnj4ymdCF+E7nzbXvto9BR7IRddgb
TD5JrZTg9qtzPo/DPscxq+XmED+OgZPqXZogpcfY/tT4zocywGO6vSVPiajYy+cV
6aJWmmEI6CFmGOqcNncLLuOhY7YqE05SBgffyjsboeoM0mnF1dxM6+IdAPfuu16C
COFPeTX7Pxq4VDDh0QbXHx9YIbng602Df83PGovMgYD/24SRhVC1XF0tjYqbsXsH
S/DPQkgHRVJQ136kp5bVWUTg007EGkT4DHp5SO0JQ0uUoBULfqmmVbR4p8UadM6D
rLJBeY1/a/V6iwxF3UOk9/p9pgsCVzMWypxAq4PsUIwWsw4ncqkJr4B5829CIJRx
9mhyUBZPDZaeCpUw07rtsZ3pG4uEE+pA2Im7mH8fsWlqKKyD1t8AK5iNRnY6Baui
RU/n6AGJK3rMLFAQxC6cslk/ZyTjxGCRuHar5i2y5oe9K8VNhx/shsKfqXdobShs
p9DywYZ4ZDQ6VrY22pGEOgMTol0TNfWegjTptUvHVmlxNrUTYxvdEKmw5WzAjYOn
/o5RPBIoyZGdGgN7Rw3jRxW8uCXOrhCcdERvaeWKnIhZmUVR+Pj07rMwoWGIEgl9
5p7FOeCDbW/TkltkVFZmJ5dDjYPtxbN6JfJ6w80MN5pZuN5EFhwVrVSzGSH7wk9u
CO+VASE4Z0XVtDVcFYvBa8n4YBsIlcPgHwjRY/vHVybSzGcmlheNHzro+muFQnVG
sj/C1zb50+HSxZ0ItM4hQJfF7cP+llSIS0+of/69MFuqGk+FjtYpJIx1uNvdNi++
0XXyjiRa9X2RwIGKNIlLxgm/8B4QuloSPzazYgpDIyYQRgLqJf6qOa2SErDpJ12E
ba845HfE+Bj/J7pVfGNIAZtlH9spyYTNQqHg55dC+5eLULdCuzgulfUW2Aw8Rw9L
9x+5WbzfqRuKBqIhD+IKtVRy7+J1+bIquC3b3Ow0a3IAvvEuGXWNccNYH+qP89jQ
uGdCPm5OzznaatfrLDlDGURBYydNePk2K2V5Z8WVb0b6Sf7drAwO4y08aIokviC1
5qjsaN9GeY/dhZplWLRYZr9sV1EitEskPPq0aPHmZjDCACVtpc05pOdxrA/HyorM
p4Y5YOgnca5V7Lgdrwv6UpXKhqklpC46wD/0L1Pqdb0rdCdd838A8OV1c56ipBLd
cu0J6COZxiqEmVxWPgnSb+8xA8/9aYIsj7x+BTKqBK/Bd3+jYqPIy5nsLKeKuIEh
JbLJRJLpo0hu+INzC7Et5vRSMtUKI92E+fHkUtI/XKoe7ggG/YvtW2LNF7rtjQMI
omrPpTUi/FSxktVF+jAnirFuzqVirxYSy/Jm4TDXK7XXXPCXpepUTpeMzzbhxCse
cmsr/fSb7gGFJw32jZXtQ36f7jU0xC/r5O9dWNlbbRuNEk/7s7M5lJV/IhHMRqfh
H1xN6k4jfruaSXby+65yIypRrJOmzgepJDvQF39I/NtnZN6LG6tKE3WW40JM82r4
s3mK+WXoPVAbFLMXN7JWlHNuNxXK1yvArHFbXZHQSwbWfofWGHXP1QWvyfFfYy0P
dNEmQh9CXQN/HJO/+FOT6pA8Ln8Xvjg1IsoANPT8om0LXMvq6kzaLeNizBLBWqML
/VGw6FUmmCfzUPeYhelKIaovX54hX/JK0SmTluLxk1Rq9MjfVmT25qY4OhvunUNc
9Q4Fs7JH8Rj/kDKBwWbroRs9gSwkN8JsKzqtvPh2XtAO2WmMdmHhUBR9O/UPCDnu
jVUjYJvkeRkUg145uAj1CRbKc+cwW6lbb9XpKwlIVKBWyhMZfJshZevVEhX+x5b/
6NyNUHlB4o/2PxGLkNiNP2YclfteTyGZev+6Jp2BKBwQw2ex5FLZ055/vbiE+t53
fnGO3924UASdUf9EMyoRRdNMphCAmsHn/R4lBCS9PdqyHr5sYw2Mz1MVxwBTE1pu
qLYpBeTKdpOVKmQ2vaNA4ylIBvRRWp1GS4eiGkH6mZuMeVinpeP3fqsLlggcJHxk
6xHgOQ3qfeQJiPZgwnm5E7rHbNGteCsMIuqoDOThnibVGIcc+KsSdCQqCrwcFVpz
AfCyRNZ8ut4k8Yz51xPTMv0rEQNbdRLaqVYsJCxZ1uMe3kUD773Wqj81076OaQeu
h5a82wzJQ1YGy/ZgIY7+31a4+hUe7PKtCbin2PzcSHHcJPsD8j2eez4yX63T/+0x
bFU8lJGYoFaGsVt6dgcJh6xpX5FoMsyNOFJiTC0DXyHgB9AICKRZVew+hIk76ujf
8R+LcXpNMDMIpNcR8eMI3rhTzrALhOkEBz0p55RXx2UEUPqBPrctr8+JHe+83KI+
2bsYvKlDOSxLhk0z1a/ELoArl4wyvAyh12ITRkzTjASINxacOja+4Ivov3wNK4cK
K5JQbOXqtSif2Tt4FqB6/ZxmcJtFOUujyLhbrgBs1yz6O/7Ujeqx3X2R2NhAlB3g
CwIxIETl+fBculZfQjCG5JJeUrBROe6wAt3LKb7puDTMtUagp77psFwwrF3qRFOv
fBlT10ww+3dYBAvs44PhNAgFuQR9EQExUHRQ5YtdpRtY5ZkUkb2+mPIjkhy08tba
GAkZP+1avc2EpwPMW5lyOHCu2iv+0Th3oY8IBiTbCh57umbJ+hRWForGCD6yXzCU
wZmm6+112IxOZl/amDVA2YROstpBUEbmAVvdUEnUKH9JKoYg0VVWpXB99ftdnc9g
9LAthC1z7XXV0TsOa8iivGC+hgwEK72y7fd3rJr+tVIMW3zsy2bY63z3KhbghrEe
DWNoTn9kYHdPW21MMXzsH/NSfRSdcxnPpKMNFbt/VHtOG3cFadKjdzkFy3JVi7C2
3MTC0qZgsGOrGwrMnbjaKxhqGXx1WDhAVU/pejQThH0D5vx6ensfmBfwvun0Jv4j
JvxwSMtDWYMgnjaAoaq0QqJdhh6hLaZV0NDbFoT0muwIrQ5+3+Pk9e1VCYjkaHmX
ujSw06RYdMYKxKRDXh1z43I54vFeX7xaJYlLNOSgcnl3u5dbJkpVUqGmo1qaftUU
eF5VYY4pA3tQgrXb36fV6s9NmpVgnIq4SIikz09YlaiJmkQZPCjA++iUk7w0yBQC
yzMERN+XGQ3utd29lsdfHAgEZIkja9tGGoaHhgn5S4SD/upMiZfE2Q+YGDiROsK8
6Nmysiw9WwNMLjJkb21ZbhBqmcrgjsOjFgYWmAdj/PPQ/urD+BsV/D+jhOCKdY5R
CmX9XriNgRGY9VVlXUHj+nKGGq/MfVQeec0RYX4belt/2ue8cvtJBczkBrir5laR
Kb/5AsPDMJmXMWppvoUAwqmeORlJGg3R8B8VYuAkd5l438o1KuCHmmlhL/Ov9e4B
9popvHjXh/dofziesirT4w545CRR3jItmHAGt4HzRJOFCjFtsCXfUVqX8U12tfAX
96GEw3/SFQLRJ61uumF7S7+p/iHo4OOwsE9Rj5w/zdA37sMDWsgGxXLNBRdGb94h
gpBffJkT2a9henpixDllIrqTM2sq0+6mHl763RxMIMgXhgpZ9h5nZGxXSWIycdB0
yXXdqM+u2JsrBJPQPyEL2dujBSEx+kyuN3TkOBb6Td7FHIBt2E2fi6eTLyvATy2Q
c3/g6dZRUnPfvtV4hUckgwqsN9O+0sCfttTd4mJbadAhEHM4+IoLJ0VUpeF2j1oS
iltZPuDZt4RPvxZ6yzc7jS9SKoQ7XtRcaV5Ukssy167EZRZNouNW3eREiREi1xOl
u8g5hgF826XQZuMTAlNdX2hPMK5g50H47O+F8IJ7vJ7rz4XrHgIO5RAJUo7Xze9T
QP4yXSWxBlwSEgC+pXWUb3JqqDFrsVeTFEPLwxz0N98U8qS/3ha8G7bMQOnnGpNd
xllJYilrRIZQjdbfUE7dUBTim5lGSCkUPMLluPHbRjr+r6aRAWyIh855pzjUH4gH
Q89aD7W4olMUAOIiI2P9cseVLgPBINBut3mC84MNoAUhBLRnc8hvq90pyH7jrPIR
bN+57dPZ9DGy4afQDXsDgXOj/5gGewKAC3WzxYEsQQR8Vh5atXeNI+FSaVTuFEDU
JH2SojEA567qn2/hFtYD0KAs0paaKUGBw/DiZLIAaYtLt4HdxnJ8IdrjAyd8WzZl
coYhyrAfvVbOUaBHmtaO7g47ygIyUElxXGWt7XzKbG+K62+uCv/KifOr2/6vd09q
Reduho/+fXbjXYNQLaMc5SHYs4NX/EEGF1ZY0dA4yB3wtAgHPuz9F6vM60JJ81vF
pyPqDgk0QbGMn3V/Ep75aAw9E12puqetrgVvs10mQy+xGe7uqjyi8KSOLo8xTtnr
4Rra3CO8Qs6kwbjiwZyMr3xnVKHZ9CmODKyL2o6r7uPznSDgrDl+01bWvvEY2EJM
dt5Fvo/4nfUviDclhSnAx7Y5dHQWSH2qmLIXdKSQmHCNIA+XTl8rWJjP4xKccs4c
X9IGrJQNzYBVgFHZDBGgSCduMYo+blISLDqmfVtESNbm7AO3bXKP4BWBtA7EZaXa
/GRSSMS5GADdKPeGL0IwNERmlgeoOkvdMPyja32RFdSL0m0qZpofPHWijwcnpklw
bCUZipuk/78PED/1+TqjLU47cpUcM/MPF7h5t0+daYHO+L+HfBemn243OA8FdvR1
V0AVOPfVtU3665nKT2KHmHoxVfNva7VgTJrPe+LhZHA0JsiumGlsqDc4GdAB35nH
8H1WReXEtxkM5bE5FXqSALucvGO5vdpHYussFs7+rzSJBGy15jj8bGWc+AU/U/L5
yQhB7ndoswvP5AbDY6uHCHMCsp1yy7rgEiRMeMbtFpNUOwBtAYkFeqVpl5lwe7f2
62xSsQRWIf+yU7luwb9wiGt4i/Q5pkGApEio6rf0mtyrrvv1Z3uq9kdlFUZcthYz
tGo0ceJSGDAfMQDTKOqpZeEUYwJP669LdkVbP50O8buWgooO42IspH2jBulgdOrB
GWTeeEUS8rKXYfKs1d494GXjmL2tg2qqL75/ACdhtisvscE8OAN2h4UYrshmhuXl
5p7zYeEZ7J31aKGEZLfk6/SoP+cCqd122EwL91/Aa9AbaSrODaL5yyItbHgDsWM/
md5hvxjhalybdaHI6qL412WxzK8YrlO/Qj9Ti1ZTxmGuZz23Vt5VVegLP59ar5XK
GwizskOGiNgAGgzQdmU+2goD0vnKZaueaW1GkYtKy4+/doKbYPTqGz36zH/wKvBk
T7ghHy/AEz9HBDSyeNTPKJjkuTRA1XAa1rPR2TofTeqV73pyqF/06kUpWKeDewu+
J9Nh98rn4qEPUA1WgzCg5HsZt+LpG7nhbw9y3jUqUv8ZH6oKBmlbdzNvmrSQBiKi
eU+rKBvGMID0tMaaXDtr4k+I/NKZbnvMh8UPth7pvRvlOqGIMLYXp8kej4UThpg1
oTvoSWUVfaxiUX8jx5PslEoYjBGLtUhxLtBrZRJgL1dZikFLTrXBhhuTHxF6BOF3
OV3/i/5fXZjyPKEXava8hnwatB3kEUBqSspzMovgqUcXxmgECDUax17B7hE1h2xH
J02tkRWOPRUA7FQVD+mvI9igtcwxPnsonjvJjn4svscpKI8IJbp/hH4Pl/5o2Mhs
aMzEOvJB+DmIW8Eis7k8mq3CAVblLINo31JVpfpEAVTN94C9810WXcaNmraHAGwn
NiJ2kfiHKQ2nkTgtdMPJ+nZUsfmCRnbGtt+KZpLgXJYr5gLpqrQXvI9jlN+pB3DU
dv21/nMMNdTsw8JVeEZhdr6xsMZ7KUG9GP841VTgUiB3r+RRH5W9LW3z5/b4uvLs
OrTurvrgFyob+wIlWB2Wsw6j3zS+x6PW0WATLSf7kQgBsWP8EnvHLJrpn5Kt1OSt
tuh0fNXxRch1eCqsc18osjRB82rfawa65r5mr+2DEtsNmb1P1eFBlb+GjJ5nULGa
Lt6NEaWOUHBQ9ES/p8wjgYIgNGQ1Z/JVNaXJwwCuS67nBbQqqn0ThAyydXeiG8i7
ikeTCoHC7c+vO1fc9k0AE5sl5MLfgRBqQJflEdrSHXA6TRqJfjsWuj9/QUs5w0mc
nnJLauZdJ9rSAx8DXiRCrNfsOL/96JXyTnCyU8rUoDGEWuOLnp92bVHRlJfJHktC
PCon3PCVoGG6VkE150lZhgccJRybwdb3p6UPIZhVgH6Haop48A0AjjOkEkwDSZXO
6RVUrHoBacDhTai4UQ2oYZYdSiQ99XUMT3Q21o/RAg94JZ+kEbUg/MTroQkbfwEr
5fp1EMwy4T9L+w6WzSB+xNlDHToNRPwsD+o0SxxF1OkkVq90Crj+7VBfZbDQAYZy
F8B0F63aCtoR15JKZ8rBKp3AjV9RCoGZPGLZvKCXl16eWZYM8+49OXGGgz65emyC
rZDN/shoou3csKfOlsBy06ID+bwg/wQu2yl7g25lAVvY+clKBw6rOHke/e7TmA2N
yHFGY4dzvRimPNSgR7VwxnPO1v1ytoOt1WS4987XuJz5d2JKBfGSuepjIKyoPtVu
7AyzWoRpHP7jFSY7WOJlgKxy6C5Okv4aSdha85Zu7vKvWjLYdwGiKePOlH+qbn/I
kJThTOdRXi+52aRsdBg2Kz8mspkcX4zYPhY/LgLyT7tj5qexz9/DtUwYsqDyQwL3
9XPEBt6mUzeR7uolNuSusajxci1m1jZmA80glvs6WYdkX1hHJ87EmUIs0fOsQYZa
xJZRfb+edb50027YW/rhSJD4DFEMK08CEg3CLWwFh9aTd0uWLbJ6TThO15hN2Q0L
TAPE73HBMS6DnbrL9UzIlDnXkl9P/Bor5jbxWbWjFTUCrSW4VbyGBqrLrvqXVdY9
LlWFsZ97MRQLnEEawW8/0rXEGe4LloqN+Yf+9duD1ZI1tQA0wMoloHsYwzLyOiDa
3Ny0li4WZI6WYatNXIRRLPAPyTg8erMFYS0c4u6MU2NUM2KOyk6YBr/oZueNZJqK
GCtTaCT4b71UWXP5TiL2qIKT1BQfjN0fDcY7TcyPnHcyA+4UysMqW8Z7ikXIVebd
zypJlybzSbyw4EAxn63u7Y/LImbxaDrG/kJRooCVNjTb7joVvV9pY2eSKBrEs9he
cgvNa676bFjm0dBB0GVB7LQqT12q1iYjc03mGFL5kuNuYCsEUy99qOMKOq7kwwAI
2IbgpSXU/7s7PPRO5m2dQkT5nHU9ahAruY7xmkrXLFTZfEHopPUFpksfqOkXmw9p
Mym1xVQfLc3OA2Xy2VPtj5iRKd/tyq38gemspR2l+cK0hfgbaB4vcci6IAgFqDEw
DaYabn+AYfIT9oZGnLMZZNZ6x+hZfLG5Gl5RBMtpTrTYbBpzWjW6EY71wcl17BiB
WeVY9SFwCHfnY4YdX1gj0QzKNG2+u8AxpQjZhnxmMls20Igx7t2X8aLqVUmk+tu0
vFcIXBbVHtP6Chpg0nUhlBYB2Ribi/maWwjGddXXPPJ23JFmaHvoJ3382Ie1d03h
xl/OYUmCaCUF72GF8H+2EwAMrrYb3tv/xSN66zqiuFfnPGV6s41Xb85tiPSgEUTA
Wgd6KVQZNBhOsTQJ8M6BQvTSuTkBOJHPz5ZQ/7dHNwxJ+VbaP5fUSkJhh3htphdm
W6frYJWAjrzkswfoOmQQRZVKwyKhZOP1Nm2VbOnn1Bv904hPx1fqGOXTMNxsQCqf
r42zmXJsCoOSxkSy2E8CkbyzN4KoZ8MNfPtSzInkJvN5mTvSxpJ2kUlUruqS4k3a
bpwFdblweC7tuoDojmwafcmcvBF0qDYwT9frXMOchhskojwaMCZdFAPOPsroUYYU
+9kX8BbmVPB+VNl+pVNIYnntOJbKff1LegIjAC0bPtxTr0J5k/yy9uxjKTxuNus6
BZZyH3YZPfrkBIUhPtDPBvdgUAyLCyRNuBNeJa75z4V9/GYxMhDOZUycBIRNbqag
ft7WN+zEcTtWbviUfW+mRrI+FxCtZ5m0qAwkWlopGEbgz2pRosqUJyMrmq6Rg8+y
Y1vQuuvPKSURewYWRTLfinin0uyDe6L1RlhbM3rdwyb6pBABOfdUtewN7VOBTCH+
xxe2s42LG1JwyiwiE3ApunXrv2g2v17Ur2xEhtqdcjWfmBMJG4AzEV/phcGbpsGl
03HNI6X/7sR6ueci4W3rgqDCuTJYZaagOdZkwr1f0Fua126nB4qSoi1lKQRpVCFI
IvfQmOla0gC3ydv4vv3yQVnretSGmr6NBl2yfwp6Q2UYjOMkfRRqWrYnp5SaH88p
1FP/5SlGwL5bnNpDWtNjT8Tz0mMbT0x23LCncRzT5p3+LVVYjK8B/raxjJ3YHgYH
SaxL5CdmmB19eTNJJlTDV+FM5wcz1Qz0tuR+SOV3AJSCUTF9BOEipd4ZemP1+UHy
wvN7MZSn9052n3PQtPIjUrbk6E5rZ0jIGXzlSXpdHpM7PE2AmRPoCk3eYeQ3eUdr
QWPxarEVrSNoMA2TUfahSF/Spg/Sc7Zw+iK3+6FKoHGXYm7OsNDT/9CxvQ5RlKUF
VtBXQcovFkZP9PFBUVK/RN93Ozi8YKsv2sn1rWOWlwBprGPwBMaP6Ca63ahR1xEy
GT1zTxniXeMeoDY2+WSnEV26951W6hd5EKqySJKuqfrbGQe4JFI+1YJwzM0E/sx4
BsadILSw1z4m5LE8vflPHSxSCU8L/ywsBe6baOx1DYrs9JjgLpog7wj4bTC2u1rX
fG8bDLlK+IFRVVaAZdSDA6skRm50NY2eOC5IkJYvfSu1lOiwpQ0ki+M8GaMzxEZf
s1jQNaXnpUkADM4dA9Q7GSBrggPbo/6Q+MUxYzKiB8jWy5joai0iQZAC1nK9OD+z
f9SD2XN2A8bErMgG21En8EUz8jqcculfQ6aYhYQRjTg1fA9WfEA2yLEWQyGu7XH6
3c/TuvxaxhQpSyugEDIxt2d1cyZiSJjBBc6318bmXPMXEP3CzKl5v/LjfzalAeV8
rs87Hbk612dFTiXL3vBZOLc9GbGFnRZwEy7BAnUUODnTSvJht4h7vhS/okqTwhBo
mpPPGBS7qwkQ26W3owDhHXctn/U+jPP+hYF6KuH3X3qVeVyahG6oZYgRDLIY1AGt
35lvlzaVdlw3ZDa4OGuXhMRS663wVIRzT+MhEkqQ195URnkW+SlbL9SMmzJXuv5n
jxjxEro1e/CjniQUuz0gpOqbI+IhQtezoeH+J3WbKTPUM5l4rrLQMaiI2kiMkD1H
kyaJh4WPGyDENSPpxryJqmktYvUOnHyQtzvkII8Wc+5TFlwuHFrY2ZnVChd+YO8n
TZD9qPeF+Ete+hYhcR8u3R8VbSKwIFLxPvsZhaFXRXBJXlMREFWElYqTM54lpDId
gvtQDCNLtxdhTrjH5gLbkJwVdj5BoyfRZ1pFDhs4K9saiGYckLM3GrkpLsZDU4Ot
RQAW0M38LMofxxIyPg/tBV6mET30FinQaTS8s+wAHeqqmTJRXGrqv57LshSzDvqo
5mX1PZ5mMFNxKjEAnzcxK7CRAJu9M9g/ZWwtmySMvtiX/YK2HnoW1pkS3EpppQLl
dCGngl4sa2ipumlmilqgpmXK1bvbT2BlcNUGvM95AMRbHjAmi55Lhy+e2nmYzgDQ
Bva6gQmCX3FyMFpUGHoD4Q1pRitpTS9xouIXGCDbwd2IY6oHzfqjXRXMTJUZ+gga
o8863tHgXm7IKYRFLAnOlSmCs6fAjrcUBDAENL7ALrHsJs6+pwHX66qUy3Fs/NMW
slmKitp2g7yGHlVWqfZ0ztEWxNK/7YWLgOnoKrfdBKm7LUj5b8j7dXURs+0+u0yI
FoOq09ljZbvUDNkYTk9mRoSwYdtYV65kzNZi6U5Cy9K0mmK63qlMfLDs9kww3iqM
3aD2vRitEMCjCsc0IpJ9/yoYHNCeHj8xY2Lj9bmvneXXzIWqQgfQMo5gqkMrXN+l
gDMPzr28NVoTeYQ7P+eSY/JgS/M2VwlwcCpAWCRNGyFG+zGL+BbizpIHorjBLmvc
8YPxT1fqmehT7t0Vexs3Cg==
`pragma protect end_protected
