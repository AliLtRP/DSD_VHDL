// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:37:38 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
i6qI3G6gNfU2/S90HgrZIHeNp/FOj3eOvf5AbjOkOcmKlLlgP43t+uUutySuEb0y
JTp7VbPedgcNQGsMZGqzgC9wW9DjALwSNy7ba4Cbblw6WwiAE84+Ze402G4TzUhG
uSWEl589UVlM8/co3vU98XnisLxx/zunfvyMr+x6Cn0=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 72832)
fJADmsHMmOEVLJa0zLtBm0krkQWCiElXCfB04y88Cwwd36MHeKuTQi5x7hZ/GLlB
kFcm0D5ZusG1HzI0SkqlCPHy+wC1Ha16Ucl/Zgrw0gXwGMVvYkUylhH76y33cd09
NLx/3cF5bsKn3fyt1R/mDrVpIJrsjRl5PzLnQnY7nbYgQ/65IQ21FsMCIAYogaZc
PhZj3lRxTVG31c04xayovpEJZqLHQiogjroOOx0KwpR2FU9VQ2FG/kpS7PTDv/SQ
be21bf5W+gJYq6mlNxqb+o1dEkEchWDn3bakB9qwgIGu82Btb0R+RVkjP4/H4VCk
+fIczfuMGItBw/8ZrlxyLqJsQ0za5b8gQPp2bi4BuHsIkriIbiTwm1ubpFE6Q/Jo
bDP12eq0qsPVb0L/+RA1bngUte2RjmwynM4/NOoq0Y7EEG6v2PsJtCi+PtIXKnQF
frRLW+LBLaAnIo+EAMJTaBUnaSqg/wugRx8D1godCc3qxZMsDqP0nG/mHzh/YgG7
b5V1osHwVpIf3UmkcLknUQcmM+WXgczFY66XiOduyyZ5j0PhqXd4SuzNrSjJC2hd
0OxOt1b9X9lE/YPcN/kcRA4SAZl149E1yB9fQ/C0loSpO7If4blBf3XNk2TAs7l0
VdL/DOEJyWHQ7Rqx+KDkfWGknUzg4nBC6gmEwGK88/vwW4wKaBS438pwRAwoO3M+
vZc4eFp7sctRocCSKMH0BHnnnRAM9k9bjniiuGIFy3Z3giOHZytK3dO8c7RnYqpy
oChMIpIk/C42BFvooLBws1b5wwq33shMUojrJjkRjhw4/awSiAgpYs86UBUut1JB
vxW52838DPiImJBEgReF6Fr7vSj1A6+ar/28d+jJ7H3w6MSAC0O55I46oIPBheK+
gLJoF5eUyllNzvivcI06KegX3deAFqxDyejdWSvWfY5iXHz9ivFvhuyu/mI2r/IW
/7UjGffQ4jnGbss5jEDiAGQL15vMSTzDO/b8UA0lYWi8kMUjJV0UkLjbSEQjyiw5
LvfAVWINWy3yOZIgY+CTqeZA7TCubCKNhaTUr58hJJIqFV42C0y4XpIfoa/90ftk
MBlRdtxOFKNgIX07rG94aSV2QN3VZyfQmYZx6nIol+f2u273/Nh+PPiCLUXfSxt7
Qv2kN8/WDUnNHSrz9ZjIpI2mNV2mGrSZ+u8KYDOlAqKnbK1ZDCwJp8p68oOp4yCj
vmX/gJ+J3xm5nuI7dzOGCepw2lwZRtImunLxDE4KWWbkD6VErXxn28o7jCR2t1wI
j2k1BflE8wzN+1VcWNszAnFUjGGpSoBfM6jEV1Va84P7PDGbYhOI8MvQjqKG8wtN
/xTsibW+QeyvCC0J22Clb8k7tXOZPsD+mFir8Ef6/MW6nO+/vsF7fCnGm16BaTnR
bmOm9lao9glT3EAIJ5xaAXfM6vKiZoEGxYT+hhRDGIQz+v4IHMHNLtXUvpk/BDhm
a7rvbDCfvbMVyzPJvA5kx9BH16jE6jt7Vs21IRTRcH5Xxu5lJ0CR5DvebDIGvwnO
z+vA3il53It8z+AyjXpQytJ25oZ3Y5/xGERDkgXpNx4dugZHLUuYtKmGNuRAeU3r
2bPcAyokXV8kYNJ2/sA9veQWbje6ZMh+w5aSx7bEnhWtcrjZJ6qS5ogONTLN+vIw
pRTHr3FK8x0aDLwBw2XXF8WA3ZfnoMSt3tpTzshbrM89qVjk4k/X+JFD6jJ+c6rn
XIEpDlLw8UZAsEkp8eKUviy3Iu0psXvUDWHeQ63GdPjaKCJEoyi7qRuBipETx8hR
C31xvnkqKQSAytGvF8tepeUHNSVWL96rXITyMHTtjplowanb+zXT9cCnQ+AKwSMC
H/WV4QwHxZsGChsrIsVT0NArslwZld1PC5dOvpwu/ZkU7JNGhdT1LZ0SsHVchnF7
cxL78u9gH1uwc053c5+kq51+PGpJEXCyvHmL75vISilU6hCpWbOsB08azrxSwBhC
9CH0aWxwCKrjRPG03prAhy6MEKbXWmLqSKLgo9YfmpkYOS522BtZS6IMTzAAV4Fd
lNfhqRVGovr8aRfLRkw/b/nveL163rt3pK6CGk4TWyb8HNQ5+UhV5Z9qc840e1/s
R4tPNGQrAF+A12A3IiKa7KU7z2nCorkn4ta8kwV8ptWXSrxzqB9PDDl1IBkWvG5a
zWmIscJ/CsahuEuCWKgAMawu7RL8UjBOkkr9/lo/v0r1zBZNag3uRfJcRGcXaDGO
TZJW+G5AXbWmzuE9TTz2JbN1ATGOJqpPCyLmfO8MZ2jO4aqAMoK6orILnjBc3E7k
BQ2Gtxm8LPHNZotweVgGg2QPPe122byU7nI6iALW0u9sh3yXWCpRmLEVgb4cMaCI
Bnp619pvAtt/cuFcm7WwLEF9afNUaaWkU0IptDKZK6mjaODzNYk1DabhFGzkyif+
/cAxaGKHsuoKayhvKPR0yrko9NrKJPn09sWHWDEi8K5HaqSJavk/36zOD4qAM+n/
fh7gHHsv1kDWWEEJ46g0N5CitO+GryPs9tzKBb2VyNg2UjPDiukMwLp4jARaItlT
xoT5pwRJooW0cjslX9TVWy+I9vQNaEec+/34TqwjnevwosJI4qjXPl/KDs1GE45q
Kt4zoxh5vPT2+WFI55zDu2cxvRSlMoG0VP8hZQKeOAc9+bTws8f2VM0g1vEyzPmP
j3x7B2FwwDk2aiu8GDfG7p9TY/vlAryZbgBs4yywZ8EwX/GSCKGAlJRgictHoWKO
YhdSm9BmS97is52VCQaJVq0K2e43rxjAqHYmbBTfSz9lYHuvEvQuIkxdY0KD0gfp
1g6iKzThIzfOuRQT4MFew0Mm5ZcxDHkP2TmeGZyYKRGwA02aoj6HrHuglNFv+h7N
ofFIW7G8jGC2N/DAuoRbMBX2O3Zie77aD9j1S5NbbHx1AiBnv8qSOzBWWQJZ864p
PDqcEgKySNE6IgLqq9k5Hho0ptB/KE0RIzriqJyaQOapR1M0JRqJxalZju6X6hfP
wSNQKin3IHtLETC3e2JaITXlRXQkmzNat9WHr76c73z7aQFvKq+se/pD+deVz3BZ
n2xF6gsEirh6+56JUiHWswlRjY4D3eAmz+r7UzoR6cBOqW1L0c0Zku+2WYBZeiHW
zZ+eyhx7DP1Sc3/CjnX8AsfFchKzR13wTkDeBhI7bNhb5R+K0wHYqBJ9M0I8Jm8i
Wy5nCb7w93WiQBFU1gOHyaUNBweG0SF5DzKJnZn2TRT2xj96aU03zu+MSDsNi6lA
c4qy1kwoKe0gXIsBXPI4bGuzwUEVLb38uevriCU12Qb/WF5dFA+QXXgpKDIjH8qU
CHeUNwfmeXzmiMJBBTfpHt7OYeIjh9BazyzrB0O+PT2O7nqpS3657U6dQQ1b8t91
ydPda5IIk2fRkJdU3eeA8CvWgBZLO/8xNEaGntbMoXp9J0CrVF1UbTnNskVA1hog
vmKuN0Q0fIpqZ9zQ144ZstEzNToxx7fWa5TtoLuB1hZNRbfmfgnTu7xxRFopcMFg
qYVUFTa8nVXp+xzFTkAPQJCqOszM/GY+0tYIKfghaCrbGotcv28mY2LOVNISF6r7
68ETLQHxtDfU4Da8KmqO1KePVXBO6st3QAlC5VHldsypff2V9Bf34R17088xxB/t
OzcNOCWFZtvK+BPVAXVXmEBVVZo8H/6NY4fKGBE+t8bZkHVDsUdW0pCuOSjq0ur3
G9IeEZtiQg2QBZQOnMWvHCSIRnxe7VyxY/7NkZ2FT4AEufzyDWKxDFu55JGQwKK5
qXkLNvBngYqLFxDpeU4ujlWQ1/C1V3HelHbwjLQWxhXp85UmlWor1/SE5KgI5RhS
Qb767FI0wuupYoAA3Sze0P5IN9nRNgt+55Hn65xR5UdkvvPyx53m0Ggkn+j2p4D2
N+qa70hFpypSZ7Zd9TtERIcfnkCc72ttqgWBDmj83HzsL1+KD6tvhFsgFv+/N8Hb
4ihpCwF2c6jHUskGIpPW72j6bOIFRCARo971CuqCvid0GEzDB02OJPSJ5dw63keG
tsHaLhq4zkzHrZytcSk+gdy5Tc3dpbVdZsH3wiwPQuKSOwuCa4u8uwuU0f7t35D9
Hi++eBmZTM01y6TGpafkDIl9Gin1c10UklG6GueNPL0HCwiFoQGLM4VEs93jR6+6
MAjg4JEfhJKFo0Z3ugNrp4gNO5yzR75rcPxGuueIaHMph3Pxzd9P8o3XpDmApgS8
AXn8bhyHc3t9AXiEzqtxoOj8kn0Kzy+8SrF+HL5juEtngjX8dTUvdY3Q/m6xaR3i
mx1/+CogFkVgLXGDZbN4acYqV+6cxx1HgUvckswBdBJ9HD5DSN882GDcyJKAvkRB
Zkk/FiryCzXlstzrZD1MPZVUcoxUIgnJlGctmoDDbUfYtT9ZVThYTBXeZsMaq6FW
pE8aFPei+VjuSnktx8cfKJc9deZIvQzR7cdPqak22ercuGvNp7eya+x/qPXK63/F
dFJiCHRy8xavvoKFDTN1TRKYoi2B91pnGJh/0i9MmdDG48XKg3/i8sfVfHQmtY+y
bdrL6df3ycSLOzuAlmKejzDUAJyXiYM45IIn+Xmg6j2vwFlpOYGUVJESqFwlhG5C
vpX5q6KYCmJ4TnKFTHegkucph5BmOAcqS5hRcmo9LjOSO8gvRZ3tTuwQurd/k1pM
eijVwrR0tk95PN6i3s9OCLv5rCyXRgyXaiMfb6iPhBXBH7Nl+aQq5FlGGHdeZ3yP
QeQq0Xd+ofHrodvgAiR1/vgmsf5mhVBdomu9hkOw8JAAwxCOWMtBMMP/aJ3cxAsI
p352xqBSpdP4e0x8LfynYTvi8cX/5K1OgiQv9XZCNOH50iZ2WeG72jEekhxjyEbn
hkoLtfuU7JxMKsJaHMSodm0z525WPFjncaWHYle7mEaI3OIfgc7hkMqJfvjOAzQ+
pDQbgAk9ujIo2sRAZWpEvwDPGREXB9cfXJwhk07Z6oh1pW14s5wj24pPc8XguZaL
tdq+jotmhafyy3i2+Cgg8UKrTEWZfpogIl/YyR8yY9Ztp0xnry8GYONe5u/2qw6X
rXjxNlOVmjC/Fwt4n2W/9g+/hllhMmM88P+58YEIZU3zP8urAARyrHFgNz6p0j5N
+P91/1PcX0J9GTRtDuz1zro8+qrktwA4G+EDnvBc6mzm2/viJHGTqSN82zOrb8KC
Ws3N/sM6REk4YuoFS3Nm0bLn1rDC6YCha6Bw6iC+ZNPi1md8uYZv60p3bo2dU4I4
XAovQ9CtV3N4XjgoMdZvHdXeiHW3Eaqh/dLGb4F1J1Wk8hPy4OywVe84veRSB6jR
+tI7onmptqdrqGC21gX5frTJEMIl/j1/FvHg6XWU5DyTDvxpW423imCaFGS9eqen
WBF2CChTK6HE91+QIeK2Vtd44E4CaDCCzWLW3WVDJ3WZ9khzd2L79j08uSGnZ8Qj
OmxLkIV546WgjsExr1gzg8IUSPJBvuLqV6jm834GvFuONSon+XT3RQ6VG9Tre+HB
3Jz81yNuwK9ORcbAPQJf19LhwsFCL6JqgI47f8WzWNokwh9Bqc4jShjCitU+xVPu
RUzyl3ZiqFkWgb8cVHUGksZr/DedGGzrSVieEPDFS+/rf4RcpxXaw8HOVTmmQLGQ
c7miICoskAtWOrt/HR4q9vm+XjJnaLSe85VzX0xDjFKT0rie1LnlzRJ2R2hfeJsn
P5aPBRQL8NkgA51o+ad5XyGFQNZ8n57NAyByD+u/SCKs/dbV8Ih67v1cokI7AWg1
4apemTaR9y/POq52utC0dVQ/LIO2tsQ93sv2Z+tflSDV62CqTzl4ZyeQP0A5Xgxm
xRp7KQW849PNpgYn+6/gAfCeT1v16pNvbV+q+PjVmq2paD2UjpaWnRgDgHpMZ5vR
bHew7Y/HVdo474YthcenzagWlAHx1DYfeo3CTdNWbVAqlaK0TbBXMeP+zTZmmPym
xleSRM2Hi1qFwRgDGpVAzclcIxrz6w/O+lrQuySO2RFwGYZj42hy53M8dmJNQ8dY
2Z9Y+i66Bx7nipW7aN6K6AqP9IXlokaJI0+aEINwNfiBXF66phf1ppNUuWQWyYIa
1/kQCEJFX+mA3VTO+PG3PCMwUGxba1qcaHDAp+vRGh1hwziHN2ViPhLsXiTl4nE2
Ke7qeYpssmHYue9JuW6eF0geyJFAfwvhVKL8fAAGyV0NHUJ61xtccI3pb8KIEFaH
lMDI9QMdG/E3VMIfQZ8Zr2Kwxzy0f0ERwahwPd7r5Qmq7Hs21Pt6MQxDGelRpXOP
maELCNtcAggbVkHP5yv8f7mbIU/f/5b8KtBex6bJHYN92QagWXpgumTWyIpR13Cf
bj4VvZHqZAcbHljFxMKVr8x9fDpXd8q67omKiOGJvq4C1ozwMYz7WJ5q8kfnzXXQ
5GK6pVW5/U59UoZe5R2f7+C7NtXOoBvMtqtnslbPJi2LQ2o1DzS5WlFjH+7eK+o8
Z9Tf3DMBygrD7XkYn5hd2V2p8ftLY49H5z1Nn525QTVzINX5TetJGvckWZHVB94B
TLi51OE3Y28dD64B7n1LYw8234B1o3lnTPAoUMCRMhRj93mrd9E1dWz0L69g6smk
/4EWO3p9yF/JO4oOi9wIbi1mGaSVUsprG8veDHL6NFj9+oudqmeZ9ZOFI726EwHr
Br+aMRWFOCZcQJt5FcyFS0XuZFSMessCzAwlDSE01V+SVCHytFtKImRW9vOriZzV
d6ASJtDxGubrM2RmKu+3Stc7kUUjM9rBCEVIwxFNkM+Bi+Lh3rxvEJVPYimb9eIX
MjL8v9t4tDsOD4MXbOcbTnViOrrS7us/QVPZWI8EzZn2WGDP3B5kx7Zla7l/kMfa
juJaElI/6Si13CR7Ev4CM7dzBk9CgV2r8QI2odxLeyut7IBm+0241SKPojFDtSn9
nXKspPbVp5MZMkk1UVIxUOtDc44Y2XtzlFgSYqTvDLVqglFqdrobZdyZYYmc7lJ7
bKiIhTQC8n/zLdjdy7sDKoNms8l7BaDFIWEk2O+eLTkqdXVI6RZiVPTfup8dTpq3
jrhx9scRmXJlYzlhbWpQve6CCcIrACiaTkzT1pmHIf7xYdU7zVpz2gQA1Wdqj8fK
DwiJZMGtzP9U5Z4AyytddF6xWYkgMkQ+WmbcGTxH0vhDA/21T31DKCIqHl9pmLBC
KBxWG5qRBOeIeNllYuP/WJbbJy5mzuFToSTsH+tcJBvOb1I4VRLVraUt+gH2l8UH
UcP8zw47l2UjcIz9qZc19kQGK7QeK4DcZuVDJ4DQ1zLDoLGAG7tTKic/bskegxZf
Hb/GYH5FsZEcs/uCx0cmJhJJD1i2ZbsL9yjkzskgJ43ezuo9c/1IKX3bS9xFNGSr
XS96juYhg6L8kZ8Bj7phEsEEjfWS2Moql49M9WdcSwHrOoZYhY1uJBQexUvCY83o
nzQ0QYcTEY8zCk7524MZNhKFTj2smSWM4QaBQ+WLFEWVwGFca6Z02OwngvC0M/ue
P8f0TABFJ1u2DddzFwxWICp7RVUH83+5SigV7QwFu5YKsggdyYPdkttJ21pw4xoq
S+u8ihmGC/NF9/46qbIYmjPr68C/062XMJiH8VPviAsYsnUpXK0B3nVw9/NHfjty
mXXLS+B7JdUxXsgxIShO1x2+j82Wa0L2XryTL+R8XnMMV99uUIqIBGXZKEBJKlGn
WTMZsNc/c57ZLOf93H/WJVMlGpAd3F2vZ4Vtd4RLbthGQuYB35qjiDbJzH3x0tZX
v4zVkoORUjxGnxxd/PlFPNFhErBWSPKnJ1vl24Ds8x74IqgRFgnVFnQJFAE8mxLs
7d1wKDGrs9XV9H9dh5OFZEKGopfePlbqL+Yj6MVPipC94UX2AC2/JAHJ8wtYRDoG
CphMIn67+3brUBpoXzb7JGPrWZF2zCCw799rFSFCP0HHCvNdXIKuaKsSZWjulQDC
APjxVrM+IG+T2AJfvAbLdDXj/b0g7L1FQs+4T7e9vXoY4JW6msBIItGjYdKLamVs
qKKx9TBC9vMXFbi2Ydg2MP2eIBRyDUaaDK26b8G8r0JkfZPmxqO+WMh7kuHfZ+68
yB7Z1aURax8aUL1H1GU6XIOayMAImBSEeZNvNsX3sgmbnbyjchLNZIbpj4kQBHgk
48/x2Ec9jK6JOarAlv80AoAz9OCUU5i/jqZAQuq0sp3NNKhKkSa3XtcCD7u//yfS
8W/uAXsL8uc/XXuhUheFmPI1doA6jneQG0tVoeBD/bBGrtrF93nLfQTi0htbgVn7
XUCTXvJ3763s1cHQGJOAzRwaJ4p/HDkA3epzhus9mv4K4rP8gi1IA+y6PqJwGc70
XnlguidLtE6FqgC78a/2T9dYtMYC5CVccL6QE6V/EixtmYv4puTxixykkOMdUeQj
RnP/IjIhTK2P5CY9s82LSr0VRiz2tDEgozeflyXGoQck8x4U1GfphbrgwT+CzagH
9KZ+O3UEsWbUnEu+5GVy3Z/SczRDaXz0i1X7SHko8j2A3CXZ4L6VhnLLHJWrrY45
vlHJ1OxlGxgeKoU2tpd+aEJKg9MswirH3oQoYFZkAPsLqIEA/v8WXShKptcvEgjI
KF48SkZywY6Qn3XN/TKvxFSvZyephxnqUGvtHllL3cd6IR5CaAmC83KHVio1xEAL
kowzi2vE6TtOH3IyagFFlpbT4qHPUssztwfW4dCjxtJXF/3nJVlRefBJs8L4TZ4I
dznOSFlE/fcKc172jDSS88W85C44YlaL/liE3QxYvYHvbDdC/PE97EqLOFNStnbe
RNGFizzqZbgVdMrUhirz2JC6L7fY2+DvWY6ZuGbbI1JXrxdAFrd+Bhpghm09MKs+
DBSXelXarLyDarXRn2XdDo4jde+F/OONxUTKdnf1DMXTyWH1ipRto7RvsQ361AgW
X4uoiEnbSwZnshfkkxppO2Jwo/JSJ5cn6n/Ouj+7zidqTYkZsXgg1U+ClIss4vfC
toRTR37CCuQ+goDfsEbRo12LcTmWMdnudb/aq7JLJWI1zUN52CGWXQ4ZaAccpG+V
Upl6Ao/Mm/L62MIqbbVvoq5WP79JpPbEaCDHf/Zn8hM9yKVeVwmBKnTpB3P1fhpI
aWBZrb3j5Lu/giB2aoPISKldUYmf/Nixj2roRq/PWCmbrNcTvwCQ/M9TszSkAk5P
+bvtHrIwLBxz2eTVyKlJb5z1tIOdYLUS9Y8kRnYZjjfubOSGaQQA7NH0lKeCUOix
CPDI5vIgt5xvPDpNRjsxhBe2Nhq3ck3tINk4b1ugXf3JCmBTNrUVZ/rZSRc+PDKg
7EDzNI9Rwl/84UcQSbvtNa2jUeTjnXjBbDH7nx85FJaYq4mhk46Fl0eGXTCcSHGG
S0khAfviDqles7O3XxaxYUyNX2/Ja0bMGwmOj1kE1o9wfZLZ1BQ14TpE/1dtUODw
QmQLuBBbL9k0rUmVUADHp+heU27bhUh1b/Di3N/qFvZ9iTInJV9CNJzXgH+bKfLf
GtEREWy2vogTCm4HqU6SKN8qDNhMSP45yBBOQRRlHggj+dzpB2dwYSHHobwht4LM
daHh5EKptnlY04eV7V1YxxGfkYeCJxBY3U/t1ZcxVsQU1poqZdLbmAuUsbI2yWWD
bwwy8hblYdbHu4f6SPZlwg8MAfU63oRn+o0R+5D0fuzQlcoa41YGnOUVm96sGJlO
2ZaQ4EihjbO7Wp3uIzOshiFkEbwk/2LQ+ZbT/Hn3beW5CIhR1+TY1lfaolA8JS2C
Ah6c/KKkjce9C3E1aXIaY7ye8rRk8b1d2kA1nnkEIfojM2hHxztdLcFWeIwVzeKm
0AE56jvQIcFlE1Kd7SnR80bmolAqPrFOnTRI42s+SDq/lgJZba5L9M6HnmuLg+YD
pBYuxaDrtvZVP3EAi6omWutOzuqg21YJEixT2G4HR+hV5SGk3CiJIVVg8Qg15LRx
wMA+6sc9XfnuBlHJGZ92y3UDCtESK2X089GcK8iFFCL2vGmyVsvzbLI4GAioGLdD
cVjHW6s9WJjUT9aTC3BQYJUXmDv5E06aus4ZUOAgicasWTxE7gaIVwt88frI+/De
8bF4jxHyxutDUfAxhRgjsHtUgFbrqCgo3yqhRBwDhVSiQTCQpzayC+Om+xUgXMEP
m4oLNxAj/xNnvyUuYBppnieDsUZ9fF6Jy2BKDKf8k6TxusTsIetH6YezFsQL5tpv
an73mJOVd/sXFN90cR9ii9w4htfTdUetag7XEhs6qy/TYIoOGnEmrQLI9Qe/Zn1H
l5DHK2GLgm7cnhQ2mQIGIQjlrCB2jUPuwSFDtgQMq1VZ3liISeDlYQHoXi9jrpWb
k8qLgsTD6+AdMzRIvmlQFoobY3CUm31LrEMVlTP0M46B+i9ZUzKDEokzViUu7Q+e
DGUAySFlxtYCBjnUERFU/QnLLdoebvNRniNAWLz8ZiTdGgFw4FfIaUFRDyqMzggE
CPzzAWy9mIdsSZa5rFin3cVwYezedi7/ENwVzF0Cw8wQ78FVTLipGXpTR9rTdjGw
WvayohMakjReP65qNoQ4tKiD0qHPUx32QTJLKO76N8rQIhBus/gOlLLqZI4Fbz1R
5gJCZoJ6C45p26sEoLgDaaxt3V6Z7EYU9u7EzLKvGxfXyVPs2MoM3iPt+NO1GNLj
jtIbV1uFhe07KSss9lEHS2IrV3WHL0J+choskutFkUN/9Pzx2wuRmBPUMTVX3Kx5
+eZTLd1YX7wmPrLQENnZo8ZlQpBWirvnWHSpWgapvSMrVd2F4dr5mYy7gi86LYYr
G9VrO/cAUu3yLMHuuZwGhTK/1LaoljtDwquVPq3tpReMkwe8/SClYn3lrCP1SE/t
flHgPVge7iI7Jz3vD4GmjdhsosVd9cbPXZ5PPkNz+WZrkdFoe/6qJbRjKKFT2xVH
Fe8F/vCeqycX/dF+7vG972tOVcaCkmm83RYl7nWymeJeN4zxzrsaw+xIxRvYdUMM
UlcaKlDxbcMw3cyUXq9uNCi8k2hfS47Zf41AGRZ58OR4uOunKCyLEpPvhW42rhsk
B/aj/UOYuPUIq/y+1rzMO9AWaq49TbC7pCjndt5NMCN3ptNOduQE02hOUj0GawJF
ILOjCONV9jr12t876BLNSTic/33QoDOVpu2PBITkJxyHO/bJ2RzCR1RnEuuwegtl
tqlz1esTX9LUCxU6/RKHinoAdOBfVeiU19gc4bXBYSbNJmr4j4J8g0lD0ljMMHF1
6ITDpz9JUbvNpIVqEcYi8tdARDoSNsZNxextD8ed9mzDW6fRY39LS+XGHCmz5tqC
HDKgJMvqCZ5gqX+/d8voNCaktbZc9WeYNbku3R9KBHtjYA2oZKsbXpGZfa2UsrcE
lVzJBaptQk2KBqXDPhxOFhkFw6SwWkK6BFnNpeu3MirkIshT3K9vb9PxU1FQjOEn
wgrK4AtHtvZbZK5eSrMe312v3zr0uyq66quZR0Os65YIBdaHJaxRRXcsY4YAHK7t
BMtv1Gv7J7VPlk1DlfaY9prEMQIdraKMF9q81Dcg90nPH/AkKIz9Idvmekc0zmNm
fPBlLCwusgeiXekgocJhnfjbWpuisSSm7dNuBVjtIQxzcnVbvKa1L1E5m/hZTX/y
AwEPeq3MXpkIZzbRK0wugkwS+veYEl2kCy0Gz4IpPHkiGtpuV1oJwyVGFTkNdFyn
aYM5HMktsnh+Bqc6UofDg+swXXrilDnlcmt9kDrSS5UtLR2ZtuIigoAzOKJjrhrs
zHpItawI9UU698fm0ZZdDYlxKPxsxGKv6ZyEXmpHUHyg0g1ogTHW1yRSpuFMOZRD
UveumuF86StjhqhJBdn2JSEhhBpCK4SGZeWVsH3nZBAl6/mCPJrMQtR77BCX/TdS
8dvrAdkNC6ZbpdOTR5gZ+Ul5NPoKMfWqG1D+7AuT/pkjNJtxyr9653m3egEdpUKL
+7wTUyRc5RfiCphdtZpzXmXBG6vZa8MTlcSFWxZ0kDg+uT3DqcoXNuwuybNOLhkv
IFvJCRi8/dTchY2vPX5j4+jYNrDCaFXZ7WWeBMro2bUEFB1aPDnl23InoC0i+rVI
bvUss44pH9bOog9a7DOw2m4vT+uHIeY06K7PiIQxHqoj4981cSiBtxdAC9BlRQQj
kDVyUqg1YIeB5zdyBfY3By5ttukky/KWSfGaVVMxj0no7uVWYvn17BhpKd91WxKr
/81dEs9UE+7outrYZTyfVxMSqNVOsAeGejGdKmwQiDb3LKb2juvCwxLWx82/fsBS
dDNaunmNnZ1rUzLJVTfbuWpPqN5I7feIIM3A47PdiNBr03BMAoIxDy3F1Ofp2U30
0yhy4+PbvqaPCRgQGyic7bTnSLii1J4rp5yxqwZObHRbRdl5ZmJpjrfHlI+oUZ97
/iBm13IT/nkxGHSMDnKTapQQbbIJHRy9tqEtfEievXfKwbAMWjDadycUpgmwPSUm
6Svy3f3Mw4X8FN4pwjTfX3aywFKXQ+1rMPAPE2Pitd2uJCyfE7xudigYAAKYbQtL
fs/Vzgse/MhN25A77vA6R1teut4fJD7khPrVzxgGIeBzUEtEj3nCNeuaSjzCVDBb
2Kq3bm2qg630TK4tgjA6HC9p9eum7kgRcnzAK12aS9llwRszzZ43Gye488DFwwBc
/Fv6a5m9FMdVx37KY/fAaSu+NJeXzl6o8J5SaEH/xMGt1653D39RJYGMPknSykZC
CIoPHZzFPSj4tmWAQ+0rPO06dB4NSVPWHcE8763cxzong0VZ2tCoZ+oc0oTEZn4w
+npWpOC96O7AXm5AKVsG3QUCVWyVLqXxqf6eBC3Cg9AO1tKf9BNQDd6P55cjCz3l
Zgd7NYloKhW8c5Wb1vLPbPNeWRxqEchAmw5RzxjnwNffCLvxavbwpAO+DZJfXZtG
A8BMGYNwD8KMJpgOOYPul+s3opi8JAac+yKeISsdpHyGb8u5yEz64Rxr4NE+it1u
o3TKvVVojMSr/WyLtYmkoZzoeypU4+MCOB8dyd4aFp/weg3BHb9ABrYJ3BX0btVT
d77AA9k0zqagFW1gG6aQl053+wkZ88NtTME16T1N11neC0auK08AwuZ4Le2ylZr1
hfJZLX8CX4kkLcS1gFtQli/re6ujjz1N/Fd/egoSMPqt5pZ4jGlg2EixPY1BZN0D
3y6LdccYciC/+AK9PPVXvXc1kTC4l8i+QBNQS3QwnX5oXPSBRQqQZoPW3wGjp9t5
RVrds0w9ElfTmlqq1h7O2sOcNzwlDCal44zumfXhqxL6ea8C5FLyYjiBxndLQj+d
LpTMDSkZRgNuiRyAYMT1lWxWyyvFLX+jc2nRe1a9EzTaAZl1n6VbZn+8jMn6IaA2
vVrPQu9WNUWmac1f5wUtCm0pMQ5lUHHYajSeni+isIifDa5oP/YpjdQttlAh4mRh
cYhod8xfJwPS8/cIq+dFCCDZOp07KM5WRBNkZA3C7A8IXvKeUa1ooSGkcmoTinDZ
m1UptH3sWuRfh4jmI8uOxgHi1F8reDu5CbqNW8Bg7JWGqJLPUqP6W6mVJ0XnSoGY
JFl+I4k895LSESFo2Rx+/e/fEt0Xwb3o5mbUwYdSdoGYubzWKuqcnP84CVtlYzN2
ac01X61MdKahf5FhoE3qqVNOYRXDSJ3YaCd/vj5mA61YEuY/7sBvzmzuqpztWZG+
Scd1hUOcZY3/uIzXLhCvKvgMa+VWCrS25hz9N8CJc9x/1anKuU57moEn4lczMAeI
Tw0Fehl054GgZtvIOPtOIn4mNgRGbrQEPVHjiBI4zJx6wgjO6GIvevJMBTsrL00w
91TYYiw7+0OrEM3xzUS3ek70+SKzCMGci33ERZeTBxImSFkz7em368UJmZ8i3QaS
0gX/LeduetVsxsV1XTOhT0crXcvzQoCwJ6SvaFyCXvoq3+x7rWAO9DeTgMkHz8YV
rImXPNptHWMxfLZC5jZRzsO+QbeLXQKXaCbhJcIYa7gqCUNJYzfv15aVeJ/Wg0Q2
9HqHtr9BcEaVnBftHrlZqItLyBlpXrYSzCRzIfL7B5nO2LhHjY7YetrwPd+IskpN
JopbzjiprJ15iPEJ+4Opfnu7EaG0T4AyqBfEji7oEZAopQyV1Ed8DeAGTxg7n3sC
3Gjmq5yoJmmL5E1noei3UxCeAa6/9LUQTdQDrjicu2hD47QaKRCM8VIdjiLKmfO1
s57Tdf0fgFA9i76FuKUAM0mazUpw6OWDrIyIqC3+JxbjTMFLG/IbPZSTJE2IJ+Lk
NRQNpgROp7dccIqL3Tw2SPEQKd24qGhocji+rZpMeOG2LRTBiRbjVKrN4Y4aRiGt
KznMiX4oyUcAifs2wB6OnS6ybwir+HmUdeqR5aKVBraEb2bwldBYFkrZRZrgwyEL
AUYdeY04rHEy06OZrWnjYs4ETlU/e2OFXodO8YUWqF3IfX9AqaXxBLKBn7qOSbOo
0AScb9VDDdPL35Owi2SQ2fcx++FHrH21RWmkKzSMbUwLJQpQQqUu2WumL2SwHe3O
DD9hI4xC2RTNhVPKxFjVo6mi6fQu3C3mw4ux62zAhmrEuO44w/mcdeUo4sZjkqEh
dXq2TWPKrF58il3LwOYcYeGKgF3nHWlrRbUacyellxqLSBqkwBmKS8iXS6rHYYOs
38D9JT/CLRQaMPy0nMx1piVWfbOU2NTh6N2r5swmgLUGb5KmmKxXBtJc8JrIAOKE
uAAohPtqGET767v0usbfgr6Vs4W2OozMX9U+84jMPQ/2hJZmlzvCd/xnwc+j9w32
FSI2eFymsOqgF9/exWlUwM+A3BEVAzToh9QHfemUaCgBeR4uAARskyOFflsza+XV
TgLEsxMO0wl/RC96FYXH9es0FI4bfelSYzgwkfileCexr7SXrp2ysAwfIRREMtYB
Wom8i5KftFA0Hvnd+aCJ5TDwXrHNLedSeTeEPPBLmvmm05jhmeU1QBHu8dLv4wME
3x0CvyqgsxsbF9TOZ3CMXvZsse0SQi3hhsBvqvPdcLdR6qm7D95wMgiMSSh9S5xO
B9sVHbHOSEa6eIiag2UY1UK+ctLf63Ap6Y6x+iny1Enup/LaJ1zPcVoDR1zeL+HM
FME0iNbzjhu50Va004ICWXYE3QLXDDeg5P1Yl88VjzinMPIXYjTVoaZsiVFzkDjj
07S0dIxF7wNS+POzsRqcbffO1yOo9grOO/O5rx4K7bsnGr3gabeyP1ONg20+n6P/
N46rFzCxjWZe+Xj8YBIpFnTH7rbOsoPZcaja2pvf3pQkQoAvqpz3+hi9wZ2di029
X4qVTNKmJMN1Ik334xYwH7l5vcmhz8v8OobiNfJQTqQSjR8HhofTDUEltjsZtEoN
oFTQwSzjTBQzcdfuRuzG5jcAyaTo/Y6D04IAqEpnESVqmvjpCBrUEae6o9UtOFZP
CUgO7c6qIPo2A1W3HoKjEc07cDsquRAbl2nQbbvSLPTZIDE15XpwAMy8kjHjwDd/
Zh5eirZkZ1NLd0WaVobaRnxSeLE9JFBqBL/ySleBBoOrpWnS96U4bgK2PpsJRqlK
mF7MA3hf2s51HzzoFUd8B+L/6FMaOf0kxyFKtqi3vtGDF5/zGLIYX9pcg1sZjKrg
dxpoJsosHtL0H81qHHoBw4b8Y7Ev9PlT3ILI92eqdM6+v8lNR4PbnKk8m4tXqnCw
B95CcLuM/ayQor+Uy0qoKZFJattwGRdLXHycVrMlW04jVUotCztKQNRms6JzTPo9
dipNWQ1xDrTtlsSAD+CW18JiZRZKXhDaSUFot5HF/gewQEYo5aUAEG1bU7n3DWIJ
bWiKeCPUS0dtc448t+O1G1xx5McWvm2oKALh2x7NPxOiV/4lavOWy/OLx10QHzXa
Z3IFiGGCiNndYAlZHG5B92CUOTgVlt+Q2qxSsUqt0sJVkfEn/4rjM8gSACRKpz+M
X8dLR+nZoEExxepiCDitP+J+vfIIbQzrR2T1xqRKmv5UeUy6eg2GtQbJEyX9OjED
qaHdwNRCSxnlntq3QzHIrzINU796mcGJ/cpNUh+0OqglJDetWFDGvgI+EVMKYNXY
ge5Pau2RTGIL1g+4fUS4Kj8NVAlvqcjUvLyiJTriylLlGIZCs4aZjulCNgB6F0SY
KN63TTLrpFgcc0Edcs//MWqQHjc9TFQABbSDEy/XsW16qWINfWKb4qG2+JC2AlNx
j5lNJCcC1ItUifQG7rTwlinCLeFh/b7S77dVYyhnAuLdUmIWnID//cDaUdqf52E7
/pEYkhswKwshNy9RUNcJStKqvcP0tf9R/QDSG8OslsPRSU+UL1y/piOUp4cac8xI
+XgAiMHFcW2mxiqk8iSDxNm7SBuB+YuVq3i1lHLTZoXBfTvGC2R0KLuP+qHA4sXA
IzGJ08cmkO1VP2uEGSV4Gn5T9hQ1IstOstRK/tqoczts0KJqJhRBDG8pJtjzY28G
f9h/YbTZz2I1y3x65v2aLefCdIKBt2QXd5/6yrngAWIP+Yk2WFJMQ1g9P2L/rQY0
7uU8BT+r2crQqT8t0ZlS5y918ylYDjrxAcXGj0wPX9+hCXUVCS/Vf/L7a85gxhDB
5b5Od/0iNNcppAJQFgwuTyCVkO3JnzVG+Av5QNCiWjJ3SHJCDWpUTuJZQ6+RQQn5
FzSE1aqIUMp0vlCy+BIMyeKrhu43on45UAhgY1FxPy0h7iY8EeoJXJNHtfZ0ErSo
AwMNSbMITwSCyDkbfKVTsJnLByZHbweqZwJYfki8Dtd10PxlOAq5DPPBrm0XTBRa
krzFa7fugqlusKkYLSYPW8EioBU1N8Yh/lY/nXlPPTrPSolLF/1oVVwJffe0K4jx
HOXcDnLZH3oUR7X/KUSBFdsAQEpc81C8ar92YDH1TESFlHe2S1E1r/dc/W7xYkCx
oS8Sreo6wXNw4ngM9vUQ0A1TSVxGR8iHDabOFil6MTj2xC7TkoYDoCxCdpCowJOA
6jlfhBxndoxlwUGYXV+wAm38amM9M4uY0gnjQGagH9t+Ft0YYyu0fwK4Md0Uw5Y0
303ykJw8mxARh25kl1xba2DRIScE46GyanZ0R99008ReB6TQ5ONDpCV4UkG1CXlf
lK4V5im+peBP1r14ho4W2BOKFQ83Di+24GCHcmDQRVTLv5cjqvFoIV1z19lE9rR5
Wim1LNspDWhHjxiHix2vIDo+WVtUypREYbGpONQLd0ZoIptkmcIiKUAsmGr92UcF
FIvWWEHawpvdSQ40ek7SU/EUgmRSyPf176cjPfT3fVYRmjmGrXahV7pmK9UIahsz
D9EbPy2UhjonN9PRgzeXB82P3wAjoo5H0kmz967zu5ql0RrnGBccYlRYRul/2kz3
XtmG036Q05EW2vYSQhEACO6dLmfJzzhhkmw1XLuRfgWGz+x8GJKeMIOg/JoS+n3c
J/jZHMd+CnpIQysgv0jwuMcPwGDWcBcNDIkmZRwveIFAw9N7+0CClMPq09+8iZKX
M/r39mZTRonb8gk6S/1C4wmEau8q3+RjtTXLc9WqOgtnCsPm6c44CStpqJz24oQC
UP7rd24UQiEF09ewfDeUx7guTRVuLlWAF07mmjDXRIg1sJhnu280wobPgLrY9q5P
vBeOL3XmJv6WjroYwPgc7Ke7p7ytsMsTc8qRpIHTVWdOhXrQ2j2iGfSxawnibBrC
OpjHehMr8+iqoxMy9d95RWEjclNFRFheDrItfgQBepa/fvKPDYU+jx5uWAXpPPnC
q5Azc5hz3zZUkRBADHpQmNV26k9ZCa58mLm0IZbqPvOVkE6smsDbsInK+jtvefBq
IrP7A9QqIsi4EYY7qYCjMM72lroDWNHXR09XHQq/JqxCiNKDEMtyv/YMUpEsupD6
CBiCxI/5Ue+rlkQ+5eMglFl9mdpzU4+wPKFGjLsEG0Vvfq5sCOcju3sTJSRoTa9g
RsPubz5J37d2Lgzs/9CT/1lpy/L4Y3wQiDziry5qiYePNI74OVn9SHchGLNPeLkm
8A3fTJKRQfCsECXwo6YrbjUBlHAXtjqyeW1i+AcbSQcZvmu/SkC70lqXJkMmXUT6
sTiV+8ed8p8Lu+wjpxSSMKXUEUj39LrUtiUFJpK5BDaOhw0AXMkzxuZXQdiCT9KG
VnSkYzc5oHxNsxzFsd9w5h4honeeCF3VJxm5q7k62wlZtT8HlkQ6nCgFmyk+W1mM
vY/ESQdWUUH7SNnQ/4CjKTTBa/doMM21RPK1rZ5yLiLXisZKR10xiTcKeWRWgvru
li4RJPjjvS3Y4OIzzdQ0Bt2thH+qp9qjeuczEpEsbeN9qfua8bEqjoeW0R/K6xb2
jyYLH6zgk/b+x/Xp8bVFQurm190AdIKaqc00etFGDzGfx634VxIXcricsN7G2IDX
BAbP8FSDdkifixdMWbsnF00JFKZJ4V94IHltmkNkucKLnaJtaHUT4gsuABN8gj17
BrD69Y+spuFor/svkMNtRcSTTIEy0dGBPnD0KDzPrpiR8QPX/zdopOlA8iCn3Lfa
SgpRMS+TKYwCBdhIa/sGXnJf/kG8GGKussirdcezWLz8i5z31qBPDUTulDCIlubn
fcuXCE3qXQOPCkHxBPjF6HWIc7LkiSju4EiynRHKkUccOLKajrSBZ5Jo7GljH8oL
+Zld6GhqjwMqdLdpihasFF05nBTFum4JI0+xJ4yFD2bdwYXHN1JvtXLmB3i/ipvy
RBvMRuAJ/6Ltj2I9fKJzcRXdeUA+aohiNCbNQG83sZzxzL2v8iZgWs6+XBHl/Aao
Z6oIsO9mkI0KPcL0ZKf63lqzSGT7P0t6428esUcAGa5imuP78ehNMHYRgu/m4CCh
l2h5yLggltYTZpRjzA+qKzdfIDRLwkO0jwZEN/rtUSmC7e3llffYnJilqGu4v0Kw
+Q+9Sq/p215Pp/fKZiY3LGrUQM95btvkx6/kCsbf0MWllS24DC/T81GJskUxdbLj
Ner5/LheCzi/Z86C9psb3cf9m+dfO0z8/voWVtoZmHfMLdATMDeY9eX3p3DPIvKt
kXr3zZSPwmfsdccLtveKFOhiF49ZlQL1pTe5BcuR5qXAX89lN9+rP41yIBxbbikR
aKqxOhOmcvEjJxOn98w0HZ6HgoSVUyax05OuXZy+4bRkV6qw23MmF7vzV7M9qxwo
RoHKNgSlAp1nW3eWpNvB6QFSLlZyp0Qz1Otzag/a84B3cH5PGtaQMsHtOa31Md1S
g2vRN21NepW4E3uPeQ7rLUN0JxlYld+5zMqI2T1jlJsEjvktHu2hvwWEwLLHBeS0
/S19zXN4pZgurXw9/xw1bTwTxw1EJ2Q5BaU6xU/x/LtYFFYEkxbM0kC6reqXVaLB
4Apwyrz6sO3UbvQBM6YFLN3ylBZg+hrHMYpiJUjTsnEu9sg7wRJIZwsgjsN7lHKF
waQOOLJN/SS8NOxGTwiSPiUQl0stde+GVqT4ni3jSRU7HGfkY+qMAMHCbI886s6z
ekX6SNUfzvdQY0CojzvgTQoKTNNHn6hgxsXknIr+hUWuIWo7ncA618c8QwfEDUGM
5S9BfboqXhoKk6SzyXAwLlJc6BhCyEq/ztG/tL6vq7qHwcSkmp8SdP/x1O1P3Fwb
CRWEVrPgyHi9qL1VVScCz+HZp4+a9ZSrJivIp+Q7Vp5QjyoUkTeHKRpTzi5lOsP+
1oFY3zYV71pVxJhaTlDETBTNsl7QQZmifn4L5mmsmwWzn2YEdSL8gHNRCE/EprzX
LFVKyjOsAkCoCCQV/6X+XQOxk7pyrSDU9XuPyYldpKkkB6IHNMmLjGPN7JQiA3xO
sH6l7LZP/9A8bUYbrw1OAG7R+mE/zEWFudyN67Y5oJNI8WOaqm2/nPd3eUYuwCqf
uS7RNDDs2hvGSHLSXCaIUC59Q4QnsBnivXV1keJ81WAuEiaDsgfwqtoVZ7Lu+LMc
/FJvkDTvhplQ9Ps2bJQzEB2TZPSgXR7dTEbbHeZt6tApTwj0F4cYKtWzlZ6qr5rk
ugcyiwj5es3/elMwusDw6esZVrUAgpVAAzYTCEvb/ROA+kpXARC6Ot+5T2K1Wdit
TpRBWwZqYOSqbM5hhV801SCkD2Yksvv+hKSwFOzYKkVvvyhRV1MdBlCFfQn8zt/H
xHhpQvnNsiLoeFDtPvHUNeUoJxLExYcTSoVQYGnV5zMnCq/I5hqAc+xEk2tgIyGN
61kse7BTkY79dR6Dv0tZL7bMWjP6szflcriKtgAVzeWzmJFlMwU2wbIqcvXplTO3
1Yl3E66bVWNkTethHu39Em484eDnQACzr6Y+S1DgdxmqveVRqTMjh/ysA1ODP7xH
9BkkVkmtaqZgjX7TLmkHMrdylLKWfNPjQ7ao6z0BwR+Q7VrS9ZM25jetM3Ce+FDm
H4K/tri4EO2pN3ENR9o4s2kgN3oltP8zmdrvONjlbo8bZ0+EQk+hJ0o3+Eq6yhrl
XHEAkac2cpAMamysbbPD8iWciujuNjQu4IG9nb2gVvuwSteqNKsBTCRBPEE03ykS
zS6g3h1STpjieJJnMuq3qiRC3dkyDYALzADdP3CLD9r0PgDhdY3bc7TmBpL50UMG
ppzdCsHye9dfhYeFFscmIWoJ2oLfDjwD9JcKMkQDPkAOyAz6T/Z7e3+gc6zTTnuZ
OLH2sb+Nly5c7VV1mHodS9gTcYFps9BPFC1JfDMFbesgWGoQ1ByD3LzqRCrWqSN+
YzIFSfHquMOKt7qYvRUwtIbQfEHJk2j/z5NgWEy64oYym32ZjLRF1IKtllbFNWtW
jtKG8X4LYhRfyjyXHZNi4KLa7/jKtUqepbvXBk/zkuvfbD7d++OYVaFxJJDqmTUI
XEm38jn1pHZTSPwE0LSpQP4cCCs5nHZwMoFRWbKLFGy2HD+zlAepI9Tfnj8gcTuD
hhw2WjA0lEYLoQ8K9dqheE5o1bNIGM++yKWqz4HI9YdfvZkAbMiT0U4QkpWEgXyz
mNuie1WjzLraIDz3GbsUbe3o7e1skm8HNhBRBIytYp0oU86d469MjPYjhYsWzXSn
oAYBDXM7dM08ZoNVwBoXeDutcw/TmGL3vuuua7nGt9KyqXW3uENQD6X+9w4ODUDV
CdpVtgkZsjhGwCyIfsw591Y3/VBbOalwhnMDrJqsC1Vza2824rxc7yVhOKB6rR4e
XM9g1f6Soz7964iMiudiT71pqfouDKHv9OEyVxrWLx4QKSnzgCsbuoYtrSn3ghoR
SU5Yi1wAGtWM5lNXRjy3e2j8W1JsgmWpWr8FNFoox12FKX1KMPqSiDlMGz44TQYL
jPywK6E/nhdq96hoRUqUqQ7TfLCf4TvwNylqIyKkVxTDqkgm27X9GTLIc+FIwhXA
rRs967zaxtxzLzWLrrRHxHr8/kO8Yj7VingQgepqogJb8lSUcVR/yeTDHrqgd+7e
d1pmoZG9aOjAFmhafKg5XJqkAaD1Adem97HuV5hP+d8NQIv/uSVa7V9gylC6fQT+
6k/vNYrSXHxs/bm1l0yC61tpL2iTs6nNztgvFOx9Xu1Aty9Nnyv+xb/JhOxrG/Oa
YwIgqg+lq0dxYzTHGi4wGzLhw7z/sU8LdsVeKaAIJWid/IgB3MnTurRNUn3ukgOe
OBGjx5j4uWr/tHegGHYZzsIB4mEQWJhDQeOjPobdO4W751D7TXyVCTSMNyAP6SsH
F/75o+WoJqW0UvIm5yo+AFE6UyJMVyB1sr/paxa3PaeW0PJValaAnJQMKtkgsEXJ
z5gBRienfKrguCbzH674gXqifbirifd+QPP+UJEkBa8Wrfm9ta94RsHX2dqJ5Npq
e2PVBhN9wK8nKo0lc79/FW1ZhTzmqf2hN+3sCpWE1i4JnQrs0XTlLSErWQ2F7wHK
D+8qsGHXke1U8Diy82okLDAAuQQkZ4CIdFmgGr21u1s+eGJKD6aKH6/h2bUhYkLg
ZvgSWQnkTAgfquELQW4NSQ/ua2iLgATBotypxHblN1cAOTvLLXq9Z3Do9Ctdjwdi
Lw1xgo/GT+PDnP5betFlJ0EZImysgK2osAZ6x939+4DvDBrOneqhUSOHU8dVu8qr
Q0UVOprq4Tj1ihtZwd5LRCQJfo1v7VzkH7APKemDRFdfFVdPkNaneXXdvMM8hZQs
1T7izl8MUEROw2RE0qpCySjKLuuN1V7P6XB6pcvRLmjwv77nQlSXAWxrjehpKsxH
7/Snj4e4IWqGeE2gkM4kS+7gdMuc4S0DoQ/BTQ2dTT3CfNlzmyQ11UXz/dit5iAs
OlObWuflLw9Wx6ewl6wb+MfiULj0XcRPoyblRt+6j3c8sX0ZYYeGXpwWs+Z4txsv
Ng90fRaOS/34JyKxap8no5bBJrxbyqeZHIGzK4FwzH/x0HaHji3urLQUIWT0W/E0
w967GuKu/7wZkBavodQjFoWDfD3pJ/65FSi8qp9PDyQuUAE9+yXJFQqRwGV1QEg1
A6JEiqsLM8FW8Xm1P1vBO9RKD9bs04Y5W8yk91aUQWfazgQW+kFiphg84YIx5Fri
8zWLtxcIvjZ50uVHiJvuRJslEsze/1ozA52lMOtSGb1mw3o7VndbOeh+bPPoSrnb
+LuwHK6FI8cSz3ElDPv6W76gKzG2tsRVs048rAnxBp/DDGNrapq8Qtwo8ZJy7ir3
NRsyL6C/0GVNTHdedDgJ8lh8fftyyO1dX2j4B7LtYWv6NW3i+YnuzfqJGqzi1TGf
PXlfubJntpolXobDIjnVCrh0Q+Xe+Q7BLHLXVYSEuhA0O0A3P+oHyBm+iTMfxWj9
zyg38EbQdr8FpJGWim+iLCnaXAdL62j2U44XxSkfObmZ+/PIpEj30bws1HZHLhbp
0LOdpMMK8VJyQjqgzDOuvmi+/8LqebWq6bKNclvWiqNtSTpHl/S33qsO9QjCPmfm
loIR36tpVrl5/G4HPikshN0Ky1/jgtH6BdrTdhCCQEPD0IxTTyWfmE204dSijarr
dErISpT4TNM4QyrREi+cVdoxsJH4ycqL43iZZ8gGxMs4svumz/5Y20wyUQdBMpkK
w4YCQ6qz4vn+dGxjiWUI+kZlgbnD8vf+cWQFuTBQDndhkBOcZIlMffmXZun0pFNU
oiq+sJ1QZETbanJsjXYk64HPRFITWbGIe54667dScxKlzgUh6UpWKVXcCrOfXBx6
aXTmXU7J5FYWfWh1uqFPhlZakEm1gAQxBFmQgu6pQG1ku6kC3HkEC4eHprCRnjKd
PyXw3kwsIaxnwEaLfKVrnjyz39YSiUEhv9/os5zBwfvc3ueLbCnJ3BCwjEIT4EJJ
t3Qf6/yvPhlVXJCY9yRdnBkBDdsypmzUX2meg9h7PDlLYYXmW4hKBvqxiN4Jj4/C
7gai0XLixRMLK5tbrrlWZsNxUNlWXtAP4f74FgJUjS+R8FtaPTAuCW3d2LETe+wr
Oi+/nc2Js5YYzYcjUKe69Nqas2Bo59qX11lWnSOdqErJRE7uT2MjI5mpWM+ryN4s
Ys/OEANUA+JZPXeieNX2l6cemiT1O1iswyE9i9aQBT2hgSUQJ+RtT619MvYsOETY
En2cvyMG/BJxpf9mvj/sRR5JmvvpdidQl5L/RcpgLt2etRDVa/hFupaGM8Z0EiIY
SgReDt61od4eSBPTycA/8YYhLJVwmb3G3tYVoJBcrKCk5i+85YQJ7LpykZp8ERcR
UCH20k2Kal8s0rxtt5sWu7WrBr71+lgyb5JS5b2yx7a1mUpibcM02igLJvN1nK/l
H4Cb2U/cOcOrsHW3vcdY8HyR9mlZypL5H2jRiZ0nXjeG96uhYsWtJmP9SnjF0ZNp
+8EFcMTF1qMjYbKPyJGMKiv2emZH+Lf6UhknRqULozIGUOpxkTKAmNK3PAfDqycT
+fIqKgKLQvto8u/l6ThfPoUJ7wqoQmMaWRXj4oNHWlrAOECL1FMPi8tYUBlmzz6z
K79eMkUb3GM0IPmACdD/NvOlTIk4d5x8jT6GWzs0u5KfDYs18YsIlfDwGUOxi/8q
AhPF9rtDAMWOrR5R/M5qHTijp5Q7Tah/x7AJK234jjRrPRDjluGmAGBIL8cJ1hR7
KN5RBjBqIiNfTxiO+JflxfwN+vaPMjseyrcsQqIf/fLLU/VBBtm9KRdLazkjjwnW
yzFTpoA2gjrwGgT1wGZGA3SIMwD18REm5LrUuG0TKcxKG65QvWSmT5j7aHLhC1zz
pGkwyUfvgA1eO6iA9Bmz4IAhbzvoRiNRt0P/adTJFES48dziMwgLnqz7x+748gbU
m7Zcz8BxByd5GMJXZ5g05aKCm+ol6LORIJJdpEcluN+H9Bq/k16pqQ5/I21dRBVc
eXnDwlE48AwZ4kb16fg/4kIWuyWBM1We5z6hcT0+q59l42FJvZcp+CZl+3U/vxHE
t+WkmQzpXvyBhIfG3WYNszsa6QdWiy7uuaIeiCeOtGcipKCCAsEIl4YRwXn6EalZ
fazG6viPz77dyzexOjJEuyIP/e1RvaPXt75LeYoGLOkr5yllhLA8tS0fGAPRc7d9
n2R3QC55uzCwuMDt2bhMflkqIZqwKK6Z1F1DOkdRiJFZzECHk8MXK0NAgmkKXcj5
NJPMJwksYur2DKV7xqQ5hJaohse6KwS16urpsbiFj35D5dGRDaNEKemvTZGyfxL2
UJtLdNhaZ4QjXFirUE7CHiNyopk9kj52LqLw4sFvbU/i5oQGlPHZrVZJJo1tIJ77
S1NgQtFF4Li+a3B1Ip/maLXzsEzVlki6Y+Wcz/QXW5lyH0KyYsbI51yNEHAS9xm9
qSuwiP+6rS25fFyXMjpRLFbyyfPPNJPOI1/FUbwbWR+Lj7lHhF55DHmbDr5nvn5Q
Gs6CI+zAtPB06Nr7SW6okDer+lzpiK7J2gTGmyykcByHXUXFgPl1lu+Z5rzfE9Up
9YzWExp03NhAShbh9v8dWwo5QpiYA3N4Jt5AAJn8j3GDDQDCpPfbgsPybbt/jh+R
O936gOZHNc2BJw2vOaFvNN0nej96yDGuDgc25b8wpEHHrodXw+PyAm9yWrt3ANMt
8TKrcaorivZdC5rJbwdxCNAdxXOUUqhbrHjzWLCJ1aZeOiuRx+AjAKZ5cyv4j5Jz
jQMhLWCQXUnJEWB7WBq/2k+5Z9Y9PscTb2Vl+koLiz/3A/LJTf0ELpb5GBp6NX7f
gvc5x0AWQBiqm982yaFUdn+ljaN2n2fWUvo/MFnJfQ8JWUfmU1xsbuafhbnLeQNp
6EqGZ4VgyrXKcIMiKQSY9Y3YJr4gM+artRThj3LTmMIYFkcVI1709/397j/bL6L8
YTBGJngxcAky8jZXjzWGE8ZaDF5/Plb+3cA1u9eY4yI7n9pDG/HkBKjtO1mEK++Y
71rKsNXQUyS6QOuXHHeaw7/6VvxuHlaHHU4EPQPijBtk6cmdzSL0v80U/umguvi4
bnAnA+exbmvv3DWoFPQTerHd3QWfXVgW2hNzAy5jn/Ipcofgrm1rOESJng1ll8kN
2j9aTHzj//w0R0fezhhmQpC5zHFCIH8Ogc2hvqrneVP8KEpeQKHkyu9JgeVu+zcb
WyEH1HQrD0OnjUEUg6vxYCx9U5BMMaID6AI2j6XYlFtPfnOGo5GVGugD3LYXQh/2
K0zyhaNtk1M+HoiGhUyuMLMw30HfZEHOebXJkyFEG9SH/M30WN2kaQow6GTmiBYN
xpVMpy9r8tIKqxsO/8gH5xHsNc5ABx72kq0JXEHWHWwCjxDBR4ZEtg4BajHmvqTO
4c9ZIxESsdmhxWO2X26q13/Xio/ongLbkTwlsrwGxh02NlW1G27Fjh3RqAreqs2F
TGFFWrtS2r97xM8sy9GQEi3gAEQ7Ly48RFn31Kx+ZXKSgfbakcGc6tPMs7DogLN6
ppHb6M+vr/bXpfp4Ke9mmVllhgeZs7Glvr/nRWqVbRTg/jzgVXSVVMUWspK+Uje0
lXaKUE72VhIIINPQBUmlTSPLZdwV5BQYK6b7gGu8HzpxaXrIbkixsUnQjQ3oHiRm
CQxzpb+de1HSDLlkmRh0TCkB97sJ5kO5qNorE1jZr07WGVD3j/ABzJJHHngnisKN
2Bucij76HCEnrs/2qXzdjKRbAAUfJtUrO+7bx5jvctQkz8RuSLlS3atFHqQ9C8qL
Br40mxNjVmCoitmYAZ2ZEv+typ47c/rUXIX/WYRLUrZqbjWvgINUmFrEmAFYYEd6
5ifzHZ5/SMFcUd9MSWyc4zA5lRm1HmulIjaQsnv9kYisHZIqmylwyfJ8B06b9EYd
FcMUmbjzmVlTgV0ZqeC4m24QhQn41i1IUrhO1a9GMy22M9ZVNLMV1Yxh/6EsXlJZ
NekOUxuEmrHnHLKnQ90BejLVvotEz++RwJpgf+ZVxQ9ogCoSWgsRUN7dstznOO64
sfuvwoPC/re6rfQ3aqWf+Gd8ktd/5Lxc+Icyk/cuVXdoMquNqdsMddOVE7YtaAJD
5YCmP3kpv5i765rWc9r7T49Jxi9bFW0EtezHLE0W1HNZN23/kNVYipycPEYejFSd
4REJ4AlWOL74CrWuQGb6Zgm8BdPXspf0IAHFnCYh6i/1jfNcJKLrEsIvIDPswFNr
sjuvcTMnlsBeN74RQ+JWaFnHe7jR3LXC28pKAveQNz4eYoqQQg5povK4ykZRSPgj
1PbMxmm8xQ16VplTU5yGct27ffzfj6TAZ1aY3WUE0r2yz5gpqC05oQsZSEj1uen6
SP0ngLtqQLzWu9EKZ/KmWR82IHo5uhMvDnEidzBMJ1ONGbYtRcPgODe85hux60PS
vEhlNpjrP8V4k663zVkuMX5w1Fx9t8DvsAIjFJAyV2YPQ/+OEng9Bp7uzg3R59jZ
honioEOh0glnrkWCChNeg5288/HbTlx9y+GzcmFh8pEU4FEu5KF8U1VCfCb08O3C
yMpHGZGIESa471EDoQSeMrf/A5f3mXTEjM12PZWAC3AWb4ygQH9E3LVqZ6Brg7qG
WWBTYBPp99oXOJklVbB/haGOrIlewIwHP7l9K8WcIlAUstnYGpiahmcH+pha43Fr
tsMnoK0dqELImG5H54eb0hzj2CXDn4Z4VcuADL1G7jNYHeTCKVyDf9Nt2Ruo5omX
kDIgWEqMPP7m9tHQwriHtfaAbCDsHdE+VJVNkY4TdMerTl4DRKiaXhLTJatc7xmi
VvTjyps7CKhiSGT7VMOulEUnkMakNufN0D53ht4r7YB5itOpEvi4WxDuwxJNuiZV
gymbrjmjRFB+xYradfVLdVM5G0qWITiut7METCVDj1Z1bLH+uhx5bF7e4Z4+lunf
MsW6YpSbo6g6VvupBGp0PHtmDX5C9EuLSgMs6TdOymCN8SwjA20bfOAeZWns05TF
G6VSMU0qp5kECzlPJdOH8jv/rC8Ve3c8q5CDDq0NDc4+Rgdm8it7Gc/LWtOXewbw
4BydzIJkm7pJVokZUUsG1+IBkuzobVDbKGDzG8ZycUkJYtY6KFbU3xWj3rCWydp2
udp4ASg2H94ssV9FHD/zg9kSea419kVoIEMdEmtKB9F5cu/BUR3IV3baZWRlKyHm
uKCFPhnXrTIrnS/HBjUP6SKVRwRQLxiRHUkEA0FNrjrkivwA7bf/BZ0jsFR8P7MJ
EzSkjrBHlqnzNKaDCHTU4Z+sy3RvPk8GbfOcmTYx8M17zo9SU1Cqc14R8Ho+y+yw
Fa7g0IfgGC3YXgx+L0wUxH1EqBL7BddUjyVNpUdiRAsWInXIA0TtfCjy4T+gwC+E
quEYEPj95SDN+tpSYuNWxGprnz+dHQkczASeojKyqpcGXOfExTnSkSJc6+wtGCas
giCB/W/MZd4WVEw/7VPp4h59L/vaT3J1i9Ov++8EZxBHbiZan5ull8Ee0fTwdcO8
8RgSmuZtPiAaf0vnuT6DVk0Kekev25fhOl0ddSL9eYzgm9Sc5U6qq4NkfrTNi7ne
JoC0qR6TQ0A3gXE2a2oXuXAd6axOL9LD4XJrVRaT1rzDWGrjJSJym/o6Pm0gpV8f
ZvtDEggmUznUQ8jGcM9tfddKdyjixbQGcnBJu81/tA1HZFG6dqXxrLM2835ykH8U
3BHZN4nnRLG8lbb8msQBrS16jdM0PFT3QSLOsJCwthX8Z/1GgeZTUP9OJ/CPB49Y
wcz8ig/wzAuh8B23pVt13bAWV4I3W2ZSpaIod23JFtbi0bgUBltYBq5XBYXcv8G6
d/iC0BFPDUNN7pY+mZmn8r0nD9XA2fFaTPUvyI9xkKK/Nj8sV4R4QkW9M8ZRwi/n
ibk8+Y97Lqs2fAMmr6WYcrRd01fdKzU5WY4TdQc86FiWKIgv4/HwTPAoF61okVg4
T4EuXPCrh1UnPD/17Y4Y46dU11sSncxK9uAZnTFgMGWrnFInbee4D+mrTrOwoQa6
18HAJ81E/VTdTDSP5wWWeTL9IdR3YQrMNZn15+ahynOd0lZ/vZrRTMqa4qELVDAI
VIBWQnF4mIIvRBFHqkW/FXtASnihyEnYnA2jVS7384K3FCYYyCCP2aFEvPZxtf06
f3INwbkA/AA+VVQHtOrSO1zv02HaOGojyEhagpf6P9LyNuTjpS9eurOX8Z4K0L5Q
fqZ+t6HzMTQ+T7wazuFm39VRv1rWKmE9x/V/Nhx8wtBp/lglJSXBfdzVI4QStPQl
QSOHZl83oHSC8jJZxN5u/oCmI8a4fgL8OlAUbwiB+DCnLASzLnLCW9cefa+FmEbS
gqc54HvvaRG8t4XCy0gqjLOSnZq3A7HBIePEI+iIjv+jaclhtSkqDCDhDn7mXzay
nJj7MqnUQi5LJkQHhxgQbe4T2Z73eXG5isWpoYi5zIyDRLpCmyYJgvjGqR8i2Ehu
AQUIPLP1QdRROjEJ3xx8OnEI+oXdM1rfvP/nGzgeeL82gWmFGwe7JCRcfj2SfR+s
EIfZx5Eo1DLM3HyZOpfUJDx/ODSaN32bh50SvCZ/aqXXLDOXIVnkecxfj88Te8NY
EAlWlmENQfNB7Ty3tjH53Pcjs/FtKAlbVtEkn83gy2QgKKK5fXVE/cqWRDDdIuxE
z9IdFS+iN9R2BUHhzK3gQtBF/20c/cLMX8nJAF1qWFuano8sVOlPqWbUKdzyzmdX
cvbCUrSy1MY0OftRRxT/7GCIBdjGLSa0gvjoOw1e7/+ZUr/GLkpfNWMl7NAygB0z
bjkl8geifewSgzT6MnPF2YpA1dWGPoGqXGLVF6LKCktnb+e0GQ6npiBl9UDl4LRt
nFFfFMaTMWdt7SI8Z5Zc3cdvOcnPedurztb412a4a5nkD3G3/WKGsYuQszElGRE/
5wyiuTnkV0XY8X4UeqEJ6anQz/G0dy/s89wvji8RYiAP62Yuv/3e1Dag8wPo5RFr
AAKK8QhC+pXTyewozR7umwHq+f7fKpoICclksSi94FbpwSvTTjfWUA1XBZXU1WcV
2dM+9FxYTMTAfuUZ62py0G8TdzcT5zS7MMZZW0vV2+CRQQij4AIFtBK3kDZPQefk
cnCgIN/fNYN4RFIf8ELqKDyFaLFk42y7rDi9P2BoCpclexw2iYP4XQb0drBFuNbY
PIognsXA3RxixiynGHg+lXvpciWlxm4kIASpjVJvntNOgkY6LWx75DM1jDnDA6oe
hhpMTIt9nUwTofk0jV3FdY/xUhX+bCE76Bgp+ho/yJax0cRyfK9P1sVExiEgigcm
o3XdiUC2J87rWNlwNzF/H2G/GN1GobmGVzAex+gD1Yy1e/FZNraDlZWFZLgr+DKF
8JBCReV22QN54uqfKC6xLxaOVrq7elzG9l85IBcRz/XDGZEukBqJ5+CrsUyjHyJ1
LUL3RrnC2A+IznSx2QBOaLKVsezEbFMP/eu0+Ikj5VlHCAct+zBbkATB21kT4lYX
146Eu4NyD9y35aJP7haADilXK5oupXpLVjrmDM31R1sja/amFKG7O/12ypHC/16E
blYClsq99X/W26PerFg5ux6SM5OP1OO6djG7YUA+U5DRSh93xA6LLWaN0bxRudZ8
gRDBI5xiL4eZ9DfrUV73/5s+/RHGPr1W8JBrxNWnnX4BPwxQe71gSMdtFGhe4rs/
I3AMErg5wCVpUziE64ifxN4YGdZQ/rAQrYz4j4FcG8JNp9jULvB3HUb6UlGghuAB
mW1/YbkpHqQz30WoyXT7xGUrwhJDWQKIXHL1rrg9W8S08fsNcnpzCbTiIXOeSVAY
DJLhBozi9+zr6VpbB7N+FvNu133l549Z+Tw8YEqhEcF7uROxpB/qsqSpxFn5RUdI
WPwxn5qvE8t3Bkxls71PARKr1X69hU6uMS+R5OdHeK0cAbgns3a1woNUQFbvNkw8
71MNpJb4YDVfvgz1zFAcw8vlIx/lENXXSV5r1pxwjbwV9IGxyZcgUkweBO84FaKk
74R4CxZo7TExeyOzjdHNhqg4TZg6iHIdM3dDwui4oByoOSSV7cRkXLQ6mPiilCdc
deoJEWobtFBTFwCNbTZ6ciqACvIhBeSBU8pTlOLU6TJMophMQUHbALzpfNNAte16
TRoBzjYKa0RkPjQlcvuQqYfIHiDm9mn1fcZRptQ1/H4rfODa74lNuIp3TXIeL0Oe
bRxT7Om9bxRMtC8EMZqjxCB18ve/2xVn/kSDOMUFjU6Ik//EVlSdYb9vQBx7zv8+
FqJLXj/gCRLPDB8x4vRrKsymJl56vGnT7I5DtUZpKgVa2ikicBgWnG/yiizK4qdQ
bwNZmjUdHFwtSrtQqAWG+jDtuxfd5D1cG4InsbLOnbkNjOYazPTtnfe2Jwf+2iyo
TySnFi0+hIlOgkfAN+k89HWbkmTOUrYYaf5skB68/fr+cYOzqLSbOkkTYLcriHWy
DK3XENUboEBMMg8ySV2hgbNhXBde1NPxT6vB9SOWeWZHscIX1VvIoEX5EZlOIWTd
KVMP7q/7oJJzT1yZYESE86QfOaBSY6kwNXZm3YcL4Xe7lYlLghrbCVuwRotRscjm
wjJuVLIEorHoqeVyEXuZoA2FJ35GcUODNf0q2mhlOZnQhdZ4UsUGdbMcDMxLn0sG
xEeubyn/q4/9fO64bd9kNFp9fxjTYC2tDIUaXAzRkwNeaf7pkysl+o1MqcCxhevS
u2LWAdIukXqQaxcb+hZJhGmAoap3gbPzTHkiog8V9idtW+AobXN9qVD1JY0avnbx
Fpo6IzZVinzYOPkTxyZlXxcMChd5bLfpLOxL9SVWmAgqOygJq94sDuqXpmfqoZCn
BzqLNHVCsyONA0x+5TFJ8whC1+Awt/3tWTIseI+l74SM5ucjBm++4HfbpjohmLWx
1IiyjHury3qXcUtY+bSZZ6P+tcKUm/FN/VPeozY3dBAy4qFEaGNqaCe803FopUC0
0iBvOoWIQoZMgyi43FGlAzT1NanxIppbmRFwE4BZSGJuavH7NJzjRk47IGAkh1QZ
6SYHoivxX6AayGbv1gW1OPAuMZpXDxZRKVQ8d0a6JP8UqPmHDrMyJXiPGEmNNXHH
ClPXsEyg4lb3siug2ReXcQPEYdO+8lxbnw9Gy8v7DMbYrPupRNfgr3Jwt+m4uN0Z
7hCLV9bcGIq4hohmppYsY10t9JM0CShmTBMIbE4UoSyKiiLhfKiuU79YCy6MP6RD
9W4jTFS3eFnyCGs9MZdffs4faDiYGUVcyndbFCFu6bWx2zmYhHMcWAdyQY4RAznq
P0vPbgrzSEORg1kqEn5/3FnXWDRRbWdf1eNLvEWeuOsSBfiOv/G1XHXOez2oTnT6
qKlAxdIsC10Y90PyOgpPqNAAq9Q5HqGxfqnqYCndWO5uQsGgKlAF1+NnkusIfWQZ
1hwG+DlL53K8mDCyjOseJ8bLJnUAMScfagS4BfgqJ63DmYLYJ/LaEeU2mCZpSEdG
03MQQDAU67TbKl6cuyWwy9tviheMKZuxOM2ZcnXKrD5zBipvVpmsADmvd2lXH7ER
GkD8g7KwPEsjnJNgWanD4GAeXUOHSUBCAF8GqyziOQOeHi2hhMAcxYjK0sxqStlv
TAXXtf8vSdvM7KiZswc8L51b6wpVxc2oVH0g82oUwiwjmkCX67pZU9WkKNMUv69B
1Wtg7jlXKbYk8lchWXv7b4NfoD4IXhh6Y/7Ro85lU2cb34cxg9SrkAIW84suSkBi
ak0rI5FKPkLBCiymGkb+7rS5TY+PFYTsXs8X3su2yqWtWItUb5dbBUMJfgxAvPIh
tPLSj2JV9xbmNebsj/uhAmft2hvJ4bMf8Spu666U+/nTed10+DfoYdv1PZ84d2xC
BsaPQsnMZqjfgYeG+tPNZgpNWVKHA12drcwctsr3iDsht9JWLXn5WpyEyJnW+SK2
O8VnF+XWMXvH2/GMO8C7c/utsvryoVddRBHGd4nMzFkoenZvuOct0mL2yyFM0MSk
cFIm3sJoyVbOneKxWCbFxJylsczoSS0s1yINAKNJoi99R5okQRoNGwDulAGrz/pr
jEa5H6HoCWagdBVVLNOIpDiWTbOw2+78nNWNhaU+Rrp5mlj/Oxh+GEFeUDd9BwLz
KOAXLZcc591wkwyruWRbY1x5GKKV2OCUexhyIuIRqdH7S3mYf69eFE8etfuOEH5P
5YqLXTi78xFBPK6nBqCxUmYRZrkUp22hk9dlywlsnc3UJb6qi7tw2SfmfpeCWvZi
h2OZ8oF8xbcvW04lqo5Hqtqy6RSqitUM3BmUjM4fK0b7HHW1jsx4Mh79onrns5AN
DoGqqu+gpvAMxrpbNisGkcq5StijGsVWlqX3OTEq9+w4WpQHZTyxZaYg4MDYjPtZ
nau03sNKFSAGDRokguGSQkcBdu/7nq1Y5JItciUrooSN2SuEmcQN8J8kZFaskUvP
/bZkJTRXpEbLo/5DkXBKYBlVADCZPAhufojxr9Dx5E5iGZHDaoCwWkxUg3dTTKD5
AByN0smnxOBepKUZ5eAeXEUGjcCWEd31yg62NR7xVr5jZRZ7FAo0USrgyy1Nttqt
mmXoZBIXkAr6MMp+n+Mhhomuoc5M6wwGjz0UCCrkb6rnQmmPPUuFD+ZA+2PMVbrT
fuxf4SgaX5oO6zGbzdDixuPZEZBWz4Y4IgsH0DpxL3Zubwr1IYN574WuN9CbG79h
ZGAVuulpeWaoDdcA4SMtEao3x5NskyWpaC5X5Ohvxq65OLunq3thK3Cek9N2LPLk
GCvaPHVcyQv4ijP1WA9NifZyGle9afu+bVXTMEFDSNw3K5GkhpIxtX8Ie5RBBY69
2m5tRDALgMVFWwJxjG90dLIb6fQrCL6Pcrf5FDY5Apy7JY+3/pLdMeSnBceQ+SMz
kiLN+4hCDhCo1YwP3ceVo5yylkvJt6jQO5U9PIaLlgBtlPQYi8Zv564mezmykOPy
7cBEYyF+4Pag1Z1TyiVIE7YAg5hMKbNH5a5XokL2VwE4fFICZzuqlprMfJMhec7s
KuNftDTxD4PK37RXLZSR4433BphqTWlUUWyAq9CLpMJ/jrm5WWq9qPa5DoLXDU6u
H8W+GlICVAj0iIHj1DcEucSnmsaGu+ckm+oaFEIgDhtv/JVdBrrrKtfLFaHGkwp2
ZusZYrYHWCKGZfv7/J8GK0WBA+ysi7DaFZd24CDpZ/M/YEOVXLTzE2BwIJBlbZHo
FHGuoMENrz3ootqDkwRQgK7DMDkW8GWWt9OxWx9saLRwUfZ9jTwe+nLTEB+kibLa
FkqTIDLq7cc1xZj84oU/6HUBb7c8IS5GKLob/WazeQgWzgfR7p4Uh2IbL7G878oY
SjnjkLdIw/IZ8k4sIDyVCcCxPCIKkBorocUJjKJwIV5X3mQUjAARC+vOm1rMvTX8
UwwX/isxVVTIoXIoXrrtWPoePxQeZmpaBMyzwcl8TFT8xmyXmaDfDUiwIn52u0Bm
CNFABc9ZhxyokAM+dyxq2yBdxbQn51ByEt0eAmgr0BGpTjpx/+ayccl3VJ9LAILW
Wgf98MrDZXHPBtr8V8j+ZbA/ejRWBcSeaeoPyM1yLIAzljslsT3gl8xHWcmKCyCJ
I8iJDuR50uk2Y3Fc1j8rtr5CsLCeXSUxN39wNYCOTTD81aIAtKff0ejPX34rl60e
YH9cEqNLeAR1v5vRYqPV9jfc+vHcaPnBBFj7q2yvFZsuVr60XKKGSTn2ThnHqPu7
D8l8OIbVQT2G9Hpjce4qNq73pCeCTyUIFEgcVBPELxui1Bc4u2J69RnF4Xgr3arB
ngJc8ATyosIiesvqmNki1fdsE1jpwTE7HDVob3YX9Y36RFfTvgblTLVxiSezvAsT
oXcLGdHouHlD+DJQKC4Ry3ul295HuiHeCRI7x/zPCYFxSeR9oFDMofvtJyGlRd43
Z2DGnD123Qvp6KzVkZKlG0ioo/uWEdu7r7Jlbfd/A/nIVevdugv7FCxd2n+E/4Z8
weKb+l/ndW1jQtMZXJrAtjHmkVQNmpEN/2uDufukBiLn18HRTgg8WN0msFS34b7C
/PkWhyUVpEXze4/YlY6GIO0XV7/KfoaeOqBj9zO4+Ua7RFlbXC/ZOydydXAhcEA3
X2sKrmrYqLRrBEiobzEswXlrFxKm8v0UyzwJt5D/1Mp1HdJmQFtOegfpjS94ssOV
1F7dnqAP0L91yERpRrhDfUW6nBxA9RimzUYpZgiFfbG7Ht6iM+PLZLlivJ9BMEu2
fPQBVmw/Yo+eAE7YoCrQRRE9vBMpU7avIpBGj5MW63MkXl/wlR4f6QVEDFXnA9Xo
D+syxQfy9fbFW0NGA3Hms+yQ9JSm3Nmzh8GycS4OggRUS4yo9U6TNbscQKvaKUd9
esBsQvdq9/E596sIKLR1gdFDHNI3ODeSDs4GnFsK0SfowebxjEWor6mHtqKFwmFS
Jn6DvPFVJxJfOwQC+W3iPQZzlL8bLFjVA65RGkS4Axa2zNf0A4ZmyuOB+r49Gq/8
0yx+If678AmA7wl+tG3d5XQ4NGuk+ysPdTdNd+KqfjANbEHCDUNYN6jNO4Z/AeVs
SyfclXBB2TE2uqLYD6yOHRTaE5A1WRrCFXmbC9x3mMHHU1N0J7Lc3mNlGknkjYrC
cvm4jT99+szToOngErC8HdwI2N3QMfzKyP79kMUaRzO6QW8nsacKc5iZpAomWeG9
Ge6TlenJZ+99CC1CE4hHxTkzoaW8uRRoS+P5wGm76ti6rLPYMEbUEbolEUgpKQk7
q85WJFnL6OhGYhnC9tBS44xTT05bKJyi4GsYJG71TTFuXhXhEzcIpdone/PRfRwM
e9T0/beVgsp7pUGfMDlq4mUeR4SHLy0SMnueRpdi8VMQQRBX91iSgcKM5HjSq7vb
5hU1ZWYqwcEVi+XrPSmp837bH09FeTCc9GQw4QpybGsBvD4y3k3vj31HrjNgE8+g
jKJRN+Zq24/JXjSep7iu0JlojItNZ1PGyxFS87ij2vTwMS/NRezAk50oXM/HGWyk
CX/iXGXCKKDj14ukvboLSjBolE5nwIZddm2zin1TSgSVVwxYKyce2yEIXUw6/KoX
vCx3YGUJKm9ImKuuB/aLdVqvnRJSm+EMKd/I4RijhY4O+r2AA3GDzpzqIrUO13w6
epCSKoAONErgeuD30i5eiwozNULYcfcwdhQflQYTGmeePmeJTVSqmAzbOUIl6KEB
6ByejaRfBjkmEHLuJ6WPAzQvS7TFV2JGD7LDp3449NBgfalUQKPwPZ7G+tBUi64R
X3/YGkcQMSkgaaSyxf2BscXK8mqQ5XWQuuGKoTICc8Z74f1MhL1/BtesST3w0NM2
O7ma5IHbryq2K+kBe45OaYdvCSW5bl+MiWLkkCtLCSx3sjKhzUDNekmGsa0VQcld
HQspE9FAIOfNHdEyUWW4kFSRGsrtfOHSUXtJXYV9+BzHvQGmVMnAVKnNniRd2x4x
nymHDatovQRFD70m1YUveLF0C3Svbcfid7jMhWDmA7ZJq7N4zGkLetJyiT9Mhpl5
OIKpiN+dC5MpC9cB248ev2IQ1+Mp0CZM6oipl1pBA2n5otcN4/2BFm7zJwPMSIdy
GYS3AXn7GXwAQ5dwOgmBuHg/j3YgiX/DM/5XFCrs9hT+/+1PypLqDnW4koBjwSl4
ulhL0lpEdBNHvVyjRCglzHGB3VlDEAb8u4TjOWxaAnCbcFm+LFMXFah5++GW5963
L3IyNfA0mVwosykFPwgpscDcMo5Un2HinMucPx+dmJ681niY76hVj895CpOJh9RS
xGp5/pfrNdDEE06jBhkHBUdu3+z8PeXWkakADqn+H3RzwG5n8j6KvEgnJvOEoJdk
8dyQKEHLlB/L5kfMzX/Dmjse5O5FDi8AMd08kw5LKeKVS71AG3IwVZar0hdw0uEZ
qwijmFt6fqcpz54RpcLmBPSS9xlb+qiRkh9r5/ItC2ov42hZKhtWk+OV+EaWaZ7f
92QV5pUWqFJi3VsD2wT4m35MF405qPbrqFuY3/aJMMdHk6TEoXiKORHii3txUcD6
2OCAsS7jQqMwJoDi3nmR4Na6WBsTwOCm5S+qXmTGO6gDCQVqAuZtpIKoSbpJZnfc
B5djFfjZMWuVGhdX6hrUiR0Yzrpbv7dCLx+8HmXyM9nlAfJUDbKrtmPcrZnNUpjK
ZB9+6tcsKvfjd524ZVEsZrYQHX+6gM1Qn2jaWiMuc7/srtO8bmJnnF7ldzSyWYur
zUSOsZgU2eIX7nXxc8h63F4DTcF+T0J+1pbv34Kn/6RqOZFRBDfSfVblbnhDCwg2
sTkINz/ZyQzZNJtOqKEbR4uyaQ/H9WW1uSoAn0sP980uo58dRk85MJrpVIG9ZOy+
dSOPoObYYhHUDnZ2DgNpxNamR2mb85dQnbaj5YobsGZHKh6dSn0ZhgHR+UjZhdIX
+DJFk+81V9xaPtfNF5lxtymi6ykdHOsOIRP7q3BjvRDZCuxsPWa9z6cZEU4FVzKg
O5Veyt3dtN0FBoaD4jnCM4oJ44AWLT0np6eSgProg2RQnAcjiOz5NSQ472TAD/9D
xEPF7VaGBvCgBq59j7jvuVbs2pzidX0S1dilXVxOTmrmt5qoSpfKSSG7lRQUDsXG
0WqJbVazK0mL1qH1z9XYQD9d+jxoijhLLwokE+dE4FPYLznySbSYhotgpgVk1Zmq
Oa7g2Kbi5f50s3w+uN7UH4TWLXQ4I4EGe30nndeDPAkzxj0LcvAcKypIjhJxfy5F
S8Cmc+9uEOVeAfD5QSMRx/Z40icmWTuoDdQTXNicFGWlVVHKW3vhS4B/xETFcnAO
SIR2Z7jdciCenuE/KkXRQoWwcIT9ykpacJmYg6345YOd18TBPzUPSrPpxtsnugP9
JOoBbcRXUqjSHcKetTV0GJdwkqtZZQZzGnomglicM61I3uM7ZTqdhEcD0eUvT9ax
tChoLvCQ0CvAz88qkuj3xXL/B0DKTtHH64imBZvRY3raJMd/lhTg8WkTXLosCK12
BMWkIso8ob4ZmN79kGuXdLqrsZ8zfXNM6gzfIUNyRX9ZQ0gMSkXNYwzr66iJuIXn
lyS0o0UUeaA62bAztY+7temPgtv6STVaWSUruIjDLZDydvAsqVT2oGvc934LmoeE
QxJ1EE1X3v/EHo+vlx6ir3VDePfFcxB0i/DztGMrRfC/nyJpV5DdHOUxyOJI4EJ+
/NdLUO4sdZRzlWFjCcjBj1PWdb/IXcIHL833Os54z8/DMBJXsspjJe4MTZtt++qW
0Yumz8C4xCq4IeMCQHrpiydbWiTuplK9Z872zQ/VLAK53mP2VY4GTq1vcZMhG44Q
uvBt8U+bFyxTQhMo1GWRLpJEf075Z95P7c1y8nXGeC4UlV27C1cdcp9Os9xJF/0H
pb01EyVJKvoSfEua2cOgII6dB37Bwsx1uMtmY3UqvSwUAfmAve7Djdu2C3UzbIxm
4qprdlMG2OSyXrAUvwRlyybuQzAP8G6qVxXBSrA8YcqzRTzCN0lhDNi+Klof32Vx
KmQzqKkdvNunScA3CR4cuZsRJ+Z9tX2NbSwOuT7+xv0bIM2HpYx8BcYT4AY66TBn
oJyWY0EvMTvcW3H5DJhYWgaC79oW6Xbj2fVkYmNIV7yUJWZh2oYgZZMOT/pV203N
Bl1dxd1jgJ3mFwX4Jm6symnEJcSTvkS65/EnyZ6oSIscBXCfhqgm3Tcn/80hMhZB
pxRCu+vGJe6B4esk6Q0vD3wfMVqixZ6sz1rKaGSDs5f7uGzUrDiXH5wNRqAKatl8
9eScpPA+m7ViBv7u/ylk3fxpaCum682evL8A4nKH+SxEPXPjN7q6IMW8zDYf54F8
84AROUCYSOX6MrYELsotiDmcs1PZsm1B6xIMrUDRmgQLOfERLPAvC5ASeWeDQ/fw
1y1sB7Y2UvfgOkLHpZmZ/l0GAFsXTkqIjiE+PF+M6WXPPqx5soEXYuOeHBFL3ECy
X6VsCT+R1CmlJvDrUFoPl0GO2KJodQt1G2dN+Riz+yESlzscORCj/uxtBXmq0FkG
vYWP7U91dIpbzyBeGjK2UiWq6C72MfgqO0uQF/8zP0g5WAjQTm36KUJ8ZC4bT14a
FqoujrQsAVU+Q5OhCNxLkLM3ZBrbnyk9/G6H/Pi4s5NS9Vq88e4QConEGmr7i8cW
nfC6ZjZqjweCgssJB+u1YN2WLWEDjpfe/T9zPz8SEjehhUpLW8FWUoigYnBS+rUM
R4E/8IWBAU5y0/VJw+2g11fk6bH70H67XK8RrF+/3hBhooxvDdiQJaoZts8EUqf+
SzH6ZsXi/bIHGfxsLWEXk0pCklxieAoSVPbRCoV6/EDvftlAAvafjt0qUX+pjPlc
7863kdmtDryJvzpPZFmKgEiHEnirDm1AyaJV/YbaovpGpBwq03dorRLxAKbWOpoZ
9RPSUU0wvZgl3QXEVe/KV9fX2mpvuj5B33bLH2/ddHB8+VXwUC70jUmMM/7DhRNM
48fKvPxuub3xLVn5aeVnlK6HxzbzH84RuoYnPuzZ39aJT41nNloZOGYEWzwVJi8a
kuT5t/VN3XtErzU787Vqz+LmssTFpRUen/8TbsWnUDC9ZTFCcdarLYjS4p0IPYNi
qYE60Q3d0tNPO4rbH0TuCGLK/DmCp4sCUn2v0zRk0nJMhA4n8CVwbSyPZEZi1frN
Y4Bcwm6zoix2RpvsxgleIF2vLh6YLya5BPEWBsJCykMrUE5vQgmTVlvwv8nYajgJ
g/pyXaANeDH8DdRznuqahSEaitAzBggA9oUtGpyOTaQHj4bgYZLolS/zk6ziHbXN
ac1F8vUsdZrqaL1fl0UmyXFIRPXlRZnhcIMl5bNPmJwE2uEhn+VmgKmHrBmB7yeo
qKHYbKFxL/7Jv2lzhSg5lbvCqi4QG40g4o28Bs0HLx/m97+ALNv9sgOJvXnj59dt
At0ze9tomcmwfPQplRfD+3Pv+AJtwHDFnPDtz0lQE1O0qmFdVln/u7skMND7VdX1
FPOuDuFyxRgImkrhWjgY2WzkKMHfYmnuXW/12vup9Dnk1mOGK+vs/G6i+Ku54Phd
fWmux7lBTSm1TINFYQH84HYlBt62tKCfkih0B1+MSr9dYUL+fo3+Vjd6lDGgvtZR
k6PY2oNqvzm81EtdCe/b8UhQKcEMDbUkZ1SzXz2oJ5jjn3s4a5js97Swmxk7TNAY
jBXDnk0AKHofn6EoLOunhR7oBfHPV5xhe34SeQqwnKzU5N012+O3mQ4JyE30pM6i
GIvLMa79Np/aD0oh0s5WLO9jAIqphhLxiiKMSKrVnrXKlTRmPgFPPR62AxBib0NL
syKiE78DSBl6w4ifzJDLP463YIlFExvOJzgRTH5wVVdGBHyO+bkgLA5MlGZ96Vpq
UVUhKdMtRBUjPm/rhmHdRyc2wzKEoACPU1L15EHtrq35ZlvC/ap0mwL61cIIOnVw
6IaNJkDsHPKAdu6FdD+3+nacihM8sta5wfftqMJoeaul9Is/s5EkU7Kt3OX8OQix
RMw3q/YHm6JHkjgDaOHRlx1Uk3FZr2HhH92oEgNooZMPrQEoz/ywlpc0ORBi2q8S
BVqKTSj5URNc2t+al2ubs3pZB/JONckWIvWIo/wNYYPvZUxCk14FCvJtRai9rilD
j4ISNwQgGPQLOHjTfJqqkLzVZnvtvERHWOfAaGBehSvG1HAPvVnv+vzb2I0GBGIA
zZ1zFls6wGoFCBV9lg5Cm1lPFk/SiJePbC0hLd9SHoo3W5CNhlUy6n3s1vfs9fxP
YD5cyIbMSSdAYKkVLoYr5ROihnVZGQ5UJU7VWR7etdaFetK+PXoRnTJbMqWg3BQZ
wwsC4KavDim5Tp9iRi8PPEwILkw6NYoSGxKFmFrvzCNsKOMKHK5uC/rXrtZJ7Ead
Zm8uQJ2u15NJoQeJ4GEToszCLVBlfo17W89kC97N2HwWwql33HI8vWAD6+uuTLR5
830WhwQ73YuQTj6VJTDENlDDWdwUEv3tXNWaFOs2tIb4WvFQB4XgqMHhOkor5OlQ
DVLIVMpoqCDMF3pYB3yqv1GrR4OWBrgnRfX/xd3dGyz2tvxH2tQfx9VTZK36zAgU
VrH2jyTyfhatRAPjVA3wzMJei/6ROjrEspKSAOMD9kWrZo55sWtiCfAgMtB8cKH9
S1JD83NtSaGvGOy5X7X9+oFyRLzLIhyfEt1kIcy9n+977/2xYgo3lc7WOHJ7gu5b
47ogONypsN3TxWgz8OGdTV0GPnD7lgrj/pBaKirwJEaq3JuU4maPfX+Ma9q3HzN4
U2A7a/UASQJvoP9Kw/ABkuR8XB7dKwDuXeTXW4L5sA015Nn9hQCEMcouc03RbnSy
fpfKq7zVNRVpvTAsKZCWIkNyWZaAfFx5gg37crU2Njp8lQC3R5xJ3D7lkQ3/xMoh
Yv7NDPg9mR1mHBDp0bN1UItKnEVwukoDGqyAGG0fE9lHCtnOxeTFXsbILHUxZovd
ZzXcUz63EpHZVQ7DoY1utAQ4otc/fNeWwzZxdn04n3DYO4WIoX3fDQOGNqbuAUh1
ARYI9WyvslwcSgA9cQ5nHyv8MN5UnF/X0nLDKzzbUeqYGj1jq7+DQ84lMooSv2IM
vKOTsNSTxcrJBfT7f59o6Lay1Pt+JK1/fcrPTs0XCgqhkqX/Pa2zq3JAMt/er/zY
DGzFuzGAjar5WWmMXvPWydSAi5S5pRSWJLpVeWKFVFYkZ8zLxIrOK/cnV8J/5kwm
dzGyC6Xv7nVNaKt8bgbsKOfixNu+kJWscFA3So0o8Iss9/GANWNlUgLOlqfgAojy
XHOM+XStxWTxLH14ujF/X4m5ZwfB9J7AlrlZ5QzCTHNBc0DAQCW6AcVJI6+wOtEf
6oU1dOq78Nw4rCEVE8NQenyl9cEr9vmJv4JOCIndKB4likvRV4cul7y2R0pcR36+
gvq2PFn0LqjxHjwO3ICEaLPEEps8awSwRRHp/zJq9ZmNM8EPXzP8QP2fA1m1/DXG
Xlf+Fhmdsy0wQkjOZqrqxfRW8Lk8qJh0u3ze30JBd3+UKhqdGGgYeAaTVGsuaVMa
Dd3tQrzIj9NsLVzSFnWBZrEyfoByZHEtSpzyVWNE0Y0HfD0uUbjLv0wVxiyy6Ytf
XT9rfwrwz+L4rLs5pDs87NPZeHh35+SSjKPovGdEZSxWNIKskKApfiGD4zozAD+s
e29vspKAiyLaFEB9mys9vtg22GvKHLfu6nPU3B5GknKxkFH5fMmoXHFYjlwNX8y6
VDaAROY44OuoIhXgONiPFnPPuQ6gk4uynXn2xFUJJIgihouaF2huAvRRXwYvgJLL
pxzkJupNy3Ic+wPncdPWofaBp1wE2/60kN9s/9MKkZvWXxZKKPfqGWglAJwwOBhT
KnxDijRgHv7ZFS/XV38RYuFFt7ykvjcmkRFZDAn/9x1vX1yYp1Pa1xFsfGMlWdWM
I/+47SdQSPlpE4+S1DMcbd2U+4bn0FtYyJfG5nv37bZhIffnRWM8eYFFwB1KzlAS
GJ+QDvNJbDiUdwOclDtRjQKhC1O3T6j2wT1tuc2HUm7AWk5hb1GeEJPHZPA3NDUb
WKD6aoAM32j9wlQ0BK1+WocsPCbgq5HxhIpdDgvV8DynuhXkyxECFlHkjD3FalrK
hnteNHW2k+pjUzgYDzG1Ro9LK638bOHyDVRXj3usqL6LPbVKi31jwIJEttdNkonp
WIABRV4iuVC2Cx1LMpn29lgz0l6uv4wD3/casA73JX9N+YT9yCUJ1bsmkGPk8NNr
qFsRkRbuID9nf1qEqnFNz6jIU5zwbGbmodGhiniwV7+zCPjugYBhTwskcTRgzuaJ
K7NbfSfFhhQbU5LWpjZ2b4ySenzuIG1aM+PbPt3ehkjJEEDOEzKIP27yC4Z22BBH
KCNLLVjvlrYB7bLXM8o1X4E+78hsIfTLzLlvMrLAUEuO8CgDSJqlYBdKdKnMnGiR
8waOaMyNHHU79BRKqPsI08dGPyEY27uDUrUItG9L/U7a/gtuVtg+bwSG4lJnmKTB
xO2gPRp2EptkkYaIsVx0xP6t8QFD55Irbl8RJKQyNpk1lD81KWiLS+PL6I10njxT
bkI2inFugCCTHmFYGZpMO9Be8AxgDijdrEa/QkGWVVuQThygpkNe7vnq0qxxWACF
iceaL7pjQ+FDjHZnl0kFnJZjBJduSqp+8AikUqb32jpjCnvZUEY7Comdt1yvK1bc
k/TqSNFqDl4k90xY3MyNs19v0myqUVp3eoNa+SiGJ1L840qW6gNJvrljsLjMu8Uq
66yQ5rjCZbQ3BxlvJZm5QEh6XJ3GDjeKKQ2Nc4XguUuVv2dXpp2pQcWd/D1lE78N
a/qhGpRvi0krfIut0eMfx1YR9Vz6PJt/xOI20dcjJgbrT9emp0n7nzSY/5t7narq
OzLX6m8LUSL7QJEQca2vgS0nvMToLG1KqpEe7VjGtR/8c8N/H40V/xH2dTEsuaKt
4N26d7dTeY5Xv3XnjQG+MNiveCOd4udnmEe0p5VJW3Fdx3pcIVimkdPc4zcCuq3c
+ywno/uHht4aiCvV0Jm3Psvfmo+efN+qGTo19Dwb1bZ6xiz7jeJIhh4U4uOKZj1T
5paaZcZM2qBBSlw7xrdhdFmz2Gqe90SaT1MdFEenIwyZBOaCVIDtXPds18mxvrbC
W/e/9/yZO8RlAJZlMcIEkrG7iACF5Tvq8f3QQFnw7yPL7Hu+Rk2dKuRHz/ngZOv6
IB7GmZyT4l7JVsmrji4R0qCF4ivaFcrUhRaPtJwzilYMAfmVR31V0tpFdz3qbooD
8pu8/C9WTx7Mfcc9n2Cx4Io0jmIW5UJNJIvGGQdjE5bX7Bwc7RXqX67AoE2cye5e
vl9NBfLwEs2MIhUbW/HchL1oUtMEu1I7vZ1y8s5D+LbsoqWtO2tlXFMqGujcHa3z
d8VgFoXa+4xS2ilqxzmtTIzOS8FBF/9GCz1xjrnQPwuhdhObQ9KvWj+/EYpeuLvZ
mB1Ipcmt+wPwJJE6H93h4bXv9Gvq9Wrwxxtr6GQVbs3njXNnr+vx8eEur4RF9+O/
Rj1aTqz7a9QUnjvFf1r6L9fT5S6FA6PKALyRTZzwHiPbNg7nBpjCvG5DPG69eVB6
dCMxvFKl8slohK+ZV/ypWWTvTspwhvDDq1fpqFnDL4/exugmNqEiYGQDsC/7e2Dm
16HdvXUavbATpw+RholTvS2x4SLUNokEAtfq3/k1Gk2vgGEGv3p8W5LuqIYimu64
9iXfXM15tlFsB+dXI/Y7aXXPa0MBQtblgeoNWe3SudpYGOD+tj+URb9Id/2Vpz7o
o7b+OK0392icBCq+tGNxRsjo011amueRzv6rMm59UFNZpCfLNg1TP6lHzobzhKc7
wVZ06SPLdO4rlkq7jEfeKoOEeiKelZg14LJh/lYqHI2pcGZAgV7S1/9EEZvjUa3Z
U0MPyjGKPD03zVz20nFmbZGjKAvPmn3CcKoJaLwyuzAz8DQ8SvVsmrIqtHQf6zCy
FJ0W77sn2VIBFob8/wEEJz4ZNSkDi4FM97NvZJmjxH9iilQeR1eaPlbHghdR4Urn
JfjG36/QmhxZiO330j84Dgg0/hzZewnglatME/vzM+vEYHvSmzLIEYnRm7+3Y681
pnzEFVMuhIczvr6ansgSN2/CMbJtZx82wxRS9opRuSw1BcaZOp39ERjSU3pIELpo
b4t7oh8Q4mxpY9rGYVJAixxwQf2AciFnzwszFb5xpmJC/SEjflqVrc7+DLI70xLH
l32u3Pg1K5tiKKTgwYpdeuHlwoPxecewziGbdNDcKtlWIqez6YMLfQ9bhmGKbQGS
2N9HBtEJ39wIrNmp4HHAZ6gxCH1rXrZKxGXmErWKrxL/iLuZ+yQZfGzqJ93Ed2PQ
IlYhkimbFpmid39UJtBHTearpBwKxeqRBkcMw2E99VFNXc8wPib7MwMUxNy7onEb
Zeg9IGiIcIUpRs9+R25UmoRBPWtepSVQ+69mDcYzX8AfD9w2Za0tZnU/o8GeQs00
2z6RVx7TuYZO7W3Z6wuU/UkHWIZJNZqmCz7IxiSMohQTlLO2wZk+0AiuXlfKo0+a
CfmigQwL/7fJfwiGlx/gGH9qHJLioDIXeKY6OtiHwqBMa4yMppWYTihbMYbF9BA4
Nxul5mi7BZR5TqjqYFZ8/UMjdjJjo7vPBAertesA0yII3e9kRF8FbaGomSLbjnCL
6NtjwZkkCcrlG1Ap1ykds2+P5OnXcZ05zin7+AwSikQEubbzHXZNQjRegMRVoAwi
7m3svXQwXhuH0PVLH+nkYoyIYOClXuPBiZ3S2irqyYW9Fp3T96y/caHlaXRoMO0n
dKKSqJ4sFynqWz6U0cUYLFv3/h8VJH968EzbRBeHuQrwzEnOqGWMXg/VJ/4ITHJD
B/Ts8Z5Os8yJLab8wr7wHS3KKbZMAHfCpL76TqF0SDLnfxnmMKArnp34JdenR3/m
gMNcAsSUjTNKmpg34GU23OyO8woJQO4MdjnGFG8hMp3BHc6MRo7QeZywkDsSg/1v
RLbzfjlElu3+0LmU/oa3i0xka4sLornUqUrUdnMm3CVFGS6c8erv94nGqtOIeUA5
nZzxj+Pf02GRnpEU2uA8Sq2H4EbGFB6aWNdPHums7nC4KVhfOd79/CaiwUFoP7u8
yyBAPbtlzPZgNhuQGST1f0nCHfIj2SS6dyf9xS6cE5K4OR1VY0n4Xt/QPpDzqwh4
hYkTqVZ6g5PLEyl9o4XypROzJzoKtfNOaG2aMQrpi688vYsT5a6/4guuXBBJgPBL
P0NUxQUCpXy7T2k75l+aZb8rXeN2gtbXhpzVcsInLhJTK31QwtXr5G1Nwdgutxbi
JE5t3QbDEKdCFM7YGqvFUcmy+gBheRzbJSrgI4lPn4p3EpKuQSkG6F8huqxMJGc2
Q0hjZhhQ68QCPM9LzR2lyFkZ5iA8zggybLvMimB2fGRmkZ3QdNkOH+EktfvaVuXm
Kw92/bKxGcL9ufJWTRzvzqpeDpVRVy9n92ru1tZdLXvqMGyjFfS3X8abLNDcZNuR
OGG6TIb2OrvTCeIbI5Jn9rV6nsCUzoq5/nIASXWBbWzV31HtrEyUkFbu5scZPPqS
PNy5mtY2kYGNPGkecIOQZFghkTpA1D8glCiPQXTavYxrHb+nCCsQxhRm4WUJqpGU
YnPoBW4grLGwgW+A2zjHAGdio3/FtzRu3W/zgIx9TXL7ccNhz+q7yMTak5zgQBGn
5O17AYnfV4muumT1MydQVAKM077HA21jlzqdKoDg6Q80D0ShQ16/QDWlX0eGnGap
wS/OKoxLE9HgZOfnacmYIBOqFJ8JxSWfapcMaRv9VVgVswFj9QL4bJBD7hN9En1O
Nqc4weQebWpTsdqlFAvJ+wDDa4VuB6juPMwrlYFt8axUcO8Mq9zzA9JduLTt20Ko
C7RjrjQzolpnxcVcgGPYSZM6dIwqXpX5O3W5gDpPM95/VXB/rKns/1UlO/vjEL+B
Vc9xoalWDSCH4MVBBYrtE5Wqzx+rFdq6D5K/yHk+hUe0lkcLCr8oN2Yi4w+R6ASj
LRJtQvWelauRSFIgsySWoUNTCkSxJm/GDKf6ogVDbcPYqZ3r5dUQXDGHBDcS7BzK
L0pOobc0s+UJw6DMGTA2sON9wzNHC7h8otOAZjL3oEzljTY59sNFQNePeu1t7/cv
s8kWQmdC1rcVpVKnxgEP81+9KYROWaNuPm8B2r/kx9sxgAmk7KoYUcZEJzt4N8lT
Iy0DPORbZKIUAa7fggos+Vttdo4ooUpFjOzDFVTIErQmWjwpqahBJ1mlOqN+eh1R
gp/wRI93j1UnNAYpivNg1Xjnjc/0X9QitPiAL2qcdRQqhcRxs3dWngyYpN+pReWn
Pj27p01QdenjvvTbAq4c7LZGsMC4x/b/ZEeaZeR7vAm0Ibsq/jeKVZy8C8aocm0I
AOCKHoNeR8hy1ABVB8zFj/FYn7ZoqxuoPMhaRh+ytwljwmjWxEF/vsPP5YF31sp1
D9MYYYnZrXrJw3EbJ15ZE2ozifl6Jg9ukeZOWjUkCgwTdHB0pvp24rIw5j/RKLGx
D+YUjdhmIAa331EfJaqCyI4xWyyOmtWl/6q0vlwz2gZfWXfoikgiSNR2gapjwVzR
GYPFALEuhMidCyER0Rkb526heAk6dAY2O+ayFaZAjP717icrd5NHqjpA/FNe0tK4
k53/ebFaOwZO44RwZgh5APF36ZONCLUJvHsda5yFIJIYlYTAs/VBFI4oUqq6FEma
XLp7s+uwhv592E/TA/T5L0gviDvRhpHqoT5ypiSYuqK06FxTWetHJQl5el5wCnFb
YBt5HEO9iGcYejgL7vE9+7vX9nrSL2lclVgPJQugFiI1WSTg4B9xClFSmJQEddyy
YbPOf+ktaLAMc3R+xUR2dzxvHuuDh/FpXvJ7b+3wmYwAPGGWNIJnJnfcwO+jDlGe
nJBPy2PhN13kYjjcqpe6gHJTtnm+S+SDWIRE4eMrH6SsSZw9iouy8FMupMtr1Zrf
nxfFeNrPZp61vexv8tCfDF7ly8JGSmA9OQkUKCGYiCJao2t2XrFKE/KZUk3hO4qJ
6NBt3ByCQHuBSslP5fYjPT8FZSESrccxp/R5y/PdWZdlBYga/W8OQheMgHwgj6SH
VwU56PeCqnRGlPLRgQQ56jPCoJ1iRBdwhBSVyJ9ScQTe2Qe+ORmzVQhbs/0rc4MS
xuJsxnXuP9KEsASn/iIzbaBpl5vlG9oU6h2f4WuSys5/tP5uZ3Wxi8xBvNVui/u1
QSFjqDT7bj4lowWtvG5LYd/ZTzn32i40tBaEtt9ouQ0+tYswHSjbNwST6CJzIZWm
MVyIYBFO4W0NZk4g9xhogiNwdRdpoyEhNm2qoz9l/cSVdga0rjHvlagcJSXaqWhU
DlIUVl+h7hT0aPd0O+0QwrL69VLWSvOohoUtSaTE4zhfe6lD2w8a/itoxyKjGJvR
0/iuI2Y1hY2MfvSeggTnv6hMQcdqkPKdW1B3njdOq+VZp3QlgzObuksHv+uHW9Et
vlQsBI3d/+FXQlYDwAt9Rkxe+itdH28Tr3KMnFuYAiqZ0u5XXUJv1JyjTU9F0VqC
cMQ6IUhfj2n4+aW2Gd/UNJBpQzoKdMFvZjtjNjyMW/jice1w2r/CD8n6/MRyagvx
ff9lwCJxk+4/oLAxB4a5N0o7THeqaxDhLUySsLwsedsY5LdW03DN06khZjfUL5FU
/dUoV24hp6TI+OdELQIw3nK1E4UlmqRK+VhkV3iysBf+nmM5p7DKd2GgSHAjA+F+
IQEjU0p+Jjk8Y9QRs84+mzqiNQ3GymhFwTpJwV9xo9CzQEKzU1Cd2ezaozMyU2bG
/Cqjfc+91oNgRynrtKMicKsUjl2StCKi7meGLT/HYp5GOGeUZCn2FMmvNzJGVxay
fDiCGO/K3yCc0Z8syebSOWX7YmcFHECJVHXxMgvIWNYMVIGo7lJVMLSa6RkDulsF
svC1jGUbNmGelcnqvOQMwnWWu52tMhkif/rWvaPLiDavhilxMV8pquweLeR4lx77
TIWvp0T8ZoyIEINr+RwtNwQSe8mQAenVUaZ4QaPSFnkCK2uFaaqBQv+6Sdac1o/R
A3UNgUgYLLETYGHDe94b+EzX5zYTX4hp2lOmAKQ/sQQWNrMosdfTGrl3S2C+D84Z
lG4mbQAOsQ10h89+tcsCCVRxxmlDW1wuIAtYyuSJf56c+CnDkP/zyYci2UaVHZUT
5vylBQCznItIsgnPgdnD18C0fpHpeATmOBfq/b1iZbs/9AES6oDAIqnDHKzO/Cgn
OR1GERb8jrkWopaYb/wRWUijwz27xvrIZYjDJ24GVlheDKLR3fnvze5/OXiGjGlz
MltoMpQ0UHxV85O8Uz2jUrq6bHrT9CQaecEB8caoaHcj1m0gRcCk+jK2tF57iYEG
LKPUsF4FRHpI5qm8I5Sraz0BrNj4RWWz6l4MpG1Hvt/VMjZg/5gYwh3eDgIkuPqk
nVPwtaIPk2AQuFKcU8dOYtX3P+QhKj64KMVWx8qejqoTsufCz65pPyy1xaxcJnBs
2wyF2DCbJeEMph02QbBhsfLRqeLG+k7LO67T7XGUA2h3OPXsXA+RPTUoyogAcwIY
0Y5uOBe3j64HPReqP+AdmW3mzHhI2gHZ4BA/zdcX65bsp2Lx6zJNnzm0s6VvLru+
PRA2mna+uAFD8lDoAhIM8MH+1o4oT3ls88J4V+kPYMUvEaSrUG4Z01GZyRZbndwW
E1u9lcMDmzUtx9xeNyBxMSA70v4IV0lIyN2DmkTqZBmXu1Ep90oyPro2eogaNcTk
ZLjCB+fOibZ6f5XPCjODGTCEZXShJiaXXLf7WjcAm05eLwKjvtSeVH8WEatw73rB
AEC2uqxCcd2G8SwiE82mZSrpeFScDGI8/Wl1w7ziThsM5q+/6vlY+tEJzgaOg65l
TmavJHHCy+rRa81OhVkvzarMQ5tx+zmUrP+gYRB3Drhqi70gecamXMeC4fR8ZkzG
ppPijuKNVyEuX1ZXmBe+EFaS8xXy9aBf9YylBhP9wWGL0twfthKZZRE4LgRXZp6J
vcOYzUUg7r7L2+8vQFTKIDOqqjzyS0apuRRZO+bNdeB88vcJdKv91yNEL4t2TVDq
7rbqdEu0GOfaKXoNHLCBz+kv64tn3taesgRpOD0k14c6pS67FsUxGclqEVHHrfrM
EC5OCMWwPm3d8WYAL4JUxZU73DAsI/lKEqBQxr3KuKlcZLpIJpNeE8A/aVDV7Bx9
uFNndpfm0L4St2RhpffHf3v/w/jDYCovuuIBkV8ipnJwvzEbuKUByNci/b+XMqqX
d9b8Tm2s5JvlPQO6Yu6vm7oYjRZJEED+Wzs1gdvyzZaenls4uwhXhHRSul4U8rhF
z8aFhloVpWOdZNe3nkeRNSofM8hfwN4i1XOl+a4gOP4fW9VvTRJgDB7NbczReUYj
psaEBQKJ0AB0mnjfzwtX0bGRB+pRWzXaUkfCDMitqgMO9Igswm0d+Is/2khLKXxV
cbdxJpPdTfsLtOO0qplG0NW4DLEpx5y4uDaaEKGHLP9NaNxkBENqJplKU7b0cmz+
hIPSy8pXN7BkiaPdrayZz53LCFejE2EFl5ik3RQS9LMT27siVNnIkoTeunwxGBi7
M/FY1UOzegTXbBYhi9rhrSiZgAhHgINq0jLRaSFZyy1bSLnoSZutCSSuAQN5zeRd
0pxA3IEjoPXxXiZ1aMZ1BAQD6E4iNJMu5zb8f4SxPYQjkPWsoKhTj/UuOES+jStm
NQp5B1XJRyLth7Zz0kYT9SokoO80p3uMHtS6a5404B05zZ3K+mX1uUnq4OnX9e1u
ecKT5+HimlZjE/0UNG++uN3wwpxPs7vFGH/fCAhF4Xa/UsYKDEVa3ywhBVo1axB7
mJ62n7dTY82uk7ZE12znHjbSb+3paj/pOHDzJOJ5MS522GCUeSQBIklFX2D1hbEc
eCRQvcNzANpNgNNTuGteDMblk3lfbQcUkTi5Cj+7GCJgWUxtalvDzJVSnc7W1ueK
UiUlZWtQ0qS6+h45EhPUl5a8FN+8BMNDTfuds/aLaaZnEP+7FGY1DQjr3ic9MoAy
JG2Np62/EKFYN0dnQmAVRKdvjsFkA93M5H+uvMf3PRhXTpeZVxg+RB4AjB9DprUw
11XS3KNUEho5Nj7qTCWlIYh3mglH8jSsEAaFEPZeIvibJXyjuz4Z20Gy+sLnmxTx
7YLQq4oexNu+03TBanx0FPNEITO5cx0OphuzhY7JH5jw1bguryhpx0iRm6cnvoRC
ZLnYMpmTf16h6JhWl7AXVa6oTLtcQeR2ojYGbcfdaGnoxA7MN12xB7FJAPQ6Lfsl
iB4elRjWNWo6O+4o1nyVni9oMfqprGR0xp0OnJ0OBdJ3q+JjiAkyHuaRLuW7A1Zb
84Coqu1mJRpiUochzXan0u6N2XGB9eWhuV8KmYXY80WExtr3KZBpQClNpu+/RaIb
BzWwTXsEWi/ST7ACgnM09fHZX7+0WwHZ+ffRmfgnwkBZ54P/GPWUqUkShq61Hjkl
xRBDuzZKbjfaU4dr+6mQpTry7hREs7zPndm5HmipPJUnxHLRB6R90QOHQ9r78koj
FpIJTB3l5jMMuF6OPhV8OprV6iHYpkJnB2U5gWnjU3bp7Fd9f2nxOiLjyEq+VRkE
fVpEMqXMNs8y9h3Vjnmhm6KjzOr5glnu2j6D8E2z3VUoniYFrWrvcu712EUGhbqr
QnomCXN/pTOeWGTiXCLhfJLaPoqNSN4XYwwKmTZZQuBOoJVv6ZyAQJEvZDicumVY
ZNfi33AzfdqaczCKoAh5iSUyvq1D10JUUCJK0IfocxVayMVNgUwgWaTbBlKrgq3a
x4NnECGbF4fdZI36sq/vBAoqVlNmWhHvAsFP4jP5/mQt1iKN0dKpR9/ZR+FyZDB4
DBoOG5X1H83wAkQ3mwOrdMguavLyUypbzpEm2apj8X0wBXP0khEThSfOslW1ofjq
nm2UH8my6sfPAX+myLy2SQ1RHYuV6iKXjgH7mzYs2QhOhtgiTJa93wiLrST3yncU
gD44BFeIHD7QjzPkrvthGOR1MxbQdpAAFGi41lPPoUyk2PoM5gAqFIU2F8+h0se2
+HHV9Y90zSMuTUBZ29+p3EOy7a7cjPs49XrXH3Mh48oKPhr0DX8u0qpIFP+d5UWj
rJHj+Hw0B2/OqtGtOFB+QVWg09BHf8jat9h6p8xi1vHgl4GoVRIurxCR+oslVKe1
+Rahpa0TUuKUS7r4gVlUDc2+1UrQHw+IG3NaG0VeNIFp5sHhlPo/Ko2HkiOlfjlR
coZqE1AmY0woAbfvmTVw33ZMsQt/kSDzJz2/ZxeiFP/RyC9M+oQMOJEa50Kv0UZl
9Mo9yX9acSdCz6BnAzNB6FXCAApvn0hKojXWq4oNxnxnBx+SAa7L1l1JtkDr79FI
bjPG7FiyoKDnCmNF6//OhnnbzZH2pVxImDxDtl7nhQ7oqndXtWVmY+nqTDO7zYhO
2JCQDGQnvPXE8UFciL/lAIgQoYHy7c2gdR2qJ6zdCoCF1lPbClrddTdXpkA1lOkY
M5tTWbU0V0BICBJNCvfPtaaC01JamesfvacyWIEEGNoQtsJfo5gX3QhztVVMDlfn
Xjhwv0oNWbItlfy6g7kciUsb8IZCXRrqDogu2fi1A5QAXoh492TVbTEDv/y8YkIn
0cl5B/XKZ5XXqWx/5omu2uT5903bXehZ6UeWZTe/dniR7VhytxD1jArH7ZRh03rl
WCbBWy7AOvRb3AfszAKIbZ0phXUmIqq66pjcGexf3g5UcqrRZLspmupyNMZRAw3M
1NTw0sQy7ayodEyA7fIMK8q8hHVjsF8E5udu2woBaEcxU+pGSCspAnOXsakFFPyb
qaWY8CGDtM6pmK3igfAqu3kaKke+wvLHCM3SPfbWVkLpPQqea1+dJhBTl5CQPwCT
tz98dd8PvkBpxkJyoZFsQybvueNwMsFhRHBrEMKa5bE0Vc+S/FZq3Gs+v5f4nW0H
K+ByiqvkbQmikuv3kiVyIthQzrK7I4bzoIcxUGp/zpwEQCmGaYL//312lEmcStYM
t/DzvttLwlT69ol2jqkbHadrcOFxtHlEtXGaboQ/8Ant/YPHcFZ0tBLWua5Az82h
1jjAyGphNFrOPgrvDC/HmpTyjufBgPwQWt6QZnonPBaRS5FLpFkvclJYw3Tjl9o5
oNZn9J7cy3yd+8BXGOoFDC7C1XjwQ+t0NVVHU0O862bCIpDiwSCCWMiKwlsys6ie
1MFq34rJox7DeSpvDn8u9EvW+YBl7eA1L9AFp7YhWiaDvu+YoTMaypUYkzaf6T6W
w0+lHOcTLxpd9bewSGwmYfU9lvfRo+BM2Zjw2ux48hoKhphxab/FikaM4gZAePOg
X14XxV4jK75Oks0ESyfgpwYwHU+Tey3rhK+mdlOvngRdKbWiA6aptzN3KFQ05Cg7
zzau5FFtdnQGYhG4i5BTxl6WtHY75OrOo3IGvOq3fP7QxjZ2LniY2AlENpnW2EAT
AQpr7nuwOWngDISZAONzE80S5VjwYdADsAt8NbQO7k4Wa1S4/WKfQgmk4KjwuM4q
9PMJrSNMzTMdqd7b1uFv/EcpWVLuxDkbhMI4270Gd6J2Wwr6w0YXamAUg8j1f6fm
eaDqzdAL17j2vcvU2R4kQH2Kgl+TSbi5IUJ7Og5he3TEmrHALsovevilP+BUou0j
rVpN0OQoEcee9K+PM2A7p+xuZE+yDRevAxsRi5e0S+e1cKFYj4PYtUFNFlEzqHTZ
BNpe9/5/Vblv2C1O6n3gUKuCvqeISzljQ0SE6J5S9vkYL+CYxhmaOgO+yEvDhfRW
QI8WtITkfeOVzKozkKyz1WZnfmQWpNWQ67YyEgXYszZe2k0Mz69rsadZ7u3xcbkK
ZkfIDOp7YZXD5fdap2bsGiAozRgIvK06Rr9pvbTJMTWLjl3EEhk0kKhpzABApzzX
6JSZoxdSl/2EjJ1mH1+DCLFV8GGMcCai4OsZMXysGGBaTQEI1+Xn1MRFGyLv7VC9
VNEgQ4dmDpQs1K4PPSs745AfH1hU1j6BvLEVH/dd9fHaUW7veQWKGtPgITIv1zWE
7V0NCHT0edT4EvVC4ei6MZD1D5uhdHq6g+G7e1Hm7wUy/VHzbmPxtnN4mUW50cI1
PkO57F1ZaA4AiAu2fdGm/8DolTp6HhcdOIxc61M36koyRoAa0H5Gpsibq95ddOlK
uTzyxa9PtY/NG2HTP1G5cU4n8LuuLfWH80nNa6RAnc0hbE8CWDR6aBhF8k1uNfiy
INstXAspMvWnJKU8CsenoacjRVC+aIP5JYoT3WKNJ6yB5tc7cmVtpf9zRt5FXAw3
wlnWWwFGheVTKUUMEqYtWBq2WkUaV0OXIdRBW2xW+mJv5V/5ISN4rfXUegDTL+b3
zRIMs7+B+6Cxeath6/gK79kFuSmaC7+40p7w5lVa8P47f6o+ZHxGQsQvmOpU4qUs
9eqfm34z33oVZWFqhWj/rgT63if77lnzqEzI15yIyoPhNbY9etGYarj6Vy41gDv8
CSW2UD0Vz69a1Q/nGOBVvC4ZzdJ0uy+vUjEVdL9NP2hQRczFXnpShDISw0EncF2s
rebrWPC4fuV5hb4WcCyP+NRAIS1rt/DeZt0oI9lm+JBbQ+N62yQ4UBSZdVeraZ0Q
x2xQQu9C34YDpNycN5oCaYaOFU5bo4kPzmJWMZeUyhuNQAZQvtwNIafXojZJO1UG
gkrWJzRjO4uZtP5TeePVUV4M3RcGmUW/YxkTKYP8bdQ8mMAQf6eKoq5g3z6Ng9q8
vCBe0pA0Bf+SouKtHwlNEOEpmAgVoExZoghXeSa+6TlYLwaryol7CHRonPDPV/Y+
3e+esxg08Z1z5ILOSHjAAlxV4bZdTuApxy1ITMGT6e7X/hIAeO0SXy+/x2AOJdcn
64JiudCFAFUJB036sRd6/YZFWyfLzlYWO8zLPT7wdv2WGNmqVxCdRvvB4Ql7OKpN
drIN5VakAdN6Cmn0dvOysTYgp2vU6e4ZdpvH6kJShif7n4F1yeMXnT0cOMM8RwLw
C0oueKlvofUV5p/5xBoqWvYKWPb6CcmE2zaHV8Pb80pYLVGdUchK1rsIh6fG7Elq
zyGW78Wi6jIzXvtaXsfcSbtPKxLH5DhqtdZIoLQxm6GF2nEXSDZK/ITWQ8fBFouj
5kXE/Xsg/+jyWHcAAszrjhn66PBUORF1MEPX6rjq7pI/EZzvfkpP3qbF+1N4KbTc
vcFL87wf9C0GiiLfXuLGXxgm3oXPgiqDwErZj0dOfje9/ZI/iuBbrmuZIVlFX7/5
aboev2PnVg8pNAwo9jZ5/X9b1e+HY2vYhTl0uzorOY2wtf6ltCajiTWcaOqeVLQS
g8iaG/wwjOkOM+sV0pVy/oxdNL5Rmc/8zz1meP+eHnP7gKPnEd/XVHlyq6jmMGj0
Xh2wO7wKtrtGBHhmfjuU0pcMHMUMdB00jZIK/Mam0Zy1cIhNA57GGEBJQ9/XRxy1
lwZ7x7NGfVQvj6NLbaR1roLqIADnCse36nIJ2rb6VHx1NROoIoL9DW85Kze7IU/W
yr82tX8xpPsJkgS6unQUKiHoGqZMsQhazgp1sjJz48mUEIKKegNmqFYOXwkdJgfu
hWtOoDI7UJukfLQPXVdfI6cagvnKMygIO2RQaqXZEUA1o7j11TJcrSBBpmU855Hk
LeL7dxpco4MteTa58fQpbHn9rcFkojEUWUdFLt5yLum6JWFOkOJGq2P7xv+r7CAj
1rkaxInrYCTCkhq5eKJWkgO5YBUPw1G9Pj6uXM0K0IA2NH3pTg8q0rl45Su581fy
5NMRoATB0bmSVoQ3IUIgi/NtLuhTErh5XmLQmNNzXLHezWbZQEUUkz57Ps1tQJNY
F2Kfvol01eLMgri5BGGFsmgjvXxDa6cV7sIZVO2xLwepDS98IZID40ULYyeu3v36
iKLEoPn0pmgCfLb9RSrXOJ1U4m9Dx21nbcopY9vGqP3zfzYiPSaVHqJ+KL3HzUyx
qOSQO48CNwlL9xD2csnOpSvdLU44Bj0oe95P2mDGLAHAsNvLgHzet2JFuSv375OO
pBrqfG4qxGb6ppE67s9Lb4ZHrFM3WOvV3ZWFTvvM60OOB5teZP4UOzjFfRylZAFy
0etwXYOmy8cN0pFJUrK7aj3aP6vqjk+pdtD6JdV7HMfWu41knpO6khrpuwgPhGpw
J1I1ATzsL1Hy3+LxNtNkSWzrcKW/VqJHDWG1Y9MfKI0TR0NyRYqRwLTx3SyNGzGO
BoOAHPSJw7/k/t2j1Qvz4DfRh9baLKwGyBEKvykCkHJO505Al3NooglJQvgnzOup
no+H4XI8NiNvkY1pCdOk+BGeTi0+OkD9h0H8yx2G0ugOG9uv+acu7gZvr/l/aoJm
o8I1Xb2yt9ebI/w4hXGare7obGFXCzXS6oVGQs/kZjlpgzWidAOieHHpafC+CXsH
y4obTvY2YBQIU390Epbb+IoTD/JgQiNtOa38zZlGyGvfpI0E7FL4UOhZtP68bgI5
och+g0ItwPhmAma/kJ98t5ktMb2OIAJ2UHBvmojmXDStTyApm5kOHz2jG7+PxueQ
9Sl+FcAHeHDxZ5BreL+a3VfMR2mlcR3zVPm+9h0ZQGAIfhsBku3bQUFzzE55S+dT
BV6x7jkZyKaAgemHwMPBV+wtnvHEWbcIEfbvjtl/LPXA0HOq0LnSE0pCQXl64azJ
1Tki99XbtnWwcGGtDKJjDYLBh7n/Ka2yVlge2CNihIWCF+aBOsVUN7sDrLrpHT0r
x2hz5Ud+TH8P7nqG6xzv9hHjTQ0dLwnF0ntfu9LcUZFb3fZxDV1D7x6KZAG0yA1Z
ELUxnKK8tnkRGBI0PLpw7qJnRQSFq6DhmYYBfd6MW1rfhRJF7ntjyXZ7KgCqas0u
N8nnOh4fYTtuqWrAAm17mPJH9+1Ea6JpHHGitRFn6zOna1ORUd/VTThqPqbwuLRp
Ju2FwOozibwI5Ec6T+dYGcPMi1rbxefMoPGnpMfjgLrGTKAgOjF4HWBAZJjOwVFv
fUgY8eUp8IbOo+ArwNH6hFTMkg1ZtXntRYxxzH+QauSAZ/2dPgQBsU9RzQfAMH+E
/k38z/a/mStPa7YfJ5+fboo6+5gKVe07WayFJ2BsuWCfmU0nv0c94cmn7lGDuHNH
lu+NeJN5Uhqt35Xo6vq60nNOFUpQIPsT0meTYFU/UNWnWqCiYh+tmxMC67cq6Ki9
bTIb7xnS2z1kCwrYobkJG5NcnMgcKKv+MFwd6xXJNctOpR9t0Nk9COSROU9hENJH
cI/eBlVtqakcK9UH9P8wmpXRet6en11DQGea/r+ks6BvAxuSWQqknlvCSoVfil1L
FHNo9hc2FZCUe6t1rQIQLb96W1mPKuFiDu97DoO3Mgl0mdFKOtTqN92C2CQ5LIWZ
jWa83CIA9xo1cdwnjy1MAQPLSYf2MkX3lQNTjq1mQazCwcdVUA3GypOF4duSyTQj
hyusHGevhcm5B+v9flq33KLpu238o705/pEVHtmM86gQXioiexHOs0XXYLPwvBKK
BSE/MYX10lmNEpFAnZOtOm1lhMAJ5lU/cRNNESiC9dywLyIJHYzFhXcrIWtAdG+c
KHOzRZnN8PH6gt52rixrGof0QPWNNYtTkWhFkzdhKMtsIkhz8XafNTdFxke3DQvc
fnR1a4zojBDKtFbIRTj2PJQLzsybopJC4Rh7K/W8CeTbSAN4h8t+on1pYZFPLG8q
TByV60E9kezJ+k4nSL2SWp5sNNI8T5r5mAvU9Z77vI1SBJpCtUESDgMSKY0V9mDI
hHmI5JdLmtLsbSAYXI6WuGFFyqDkAmgXrIXH3XAdWwzvi6Uwymb6DUlqzBrbNeUB
cWJULmqjCNg7ZAHY/i5PsHU+0NET06hVUErWqzJOzgEPvv6tfK01LVpvrEJ+NwTV
Pjoz/iU3HDnVMc2o5NU6JSOJ9EF7AaxkgIodQTy2tieqtLhAuDRbXnG1iEGGifoq
DXcDfPROZVmMlDL0K2aKgGn21KTGHPQh8eqalUADGYq4nquKR/fvrDA51YYgORCp
l3KvybP2XxlU52vRQHYZb8PkaMAxWzM7c1jksHgyhax0w8HqwKbogoIpL/3Gd+Po
X2LuyEz/3rPSkWKSAEoHwWY6QKoj0KZXSeyQ5rTKKtyojuLwbzhL5GI6wSxzvNI2
V3UN38GBXfLIEKi9DqOZ3ivJk+vFYnflQwNK1CzBWixyHbsI1PbCMuzexdvRQbhP
8IyZXWzste877oTdR1KOdFnam6nObmLchbgKJ2ugghj5MBL1rPvyAympiyZ+RrEq
AJDT31SPtxCfvrgV0ruNX0eG6JAmPVmoeXfWIxrzj/FG2rGuCLzwYE8R+yIBk2rY
Wzo8b7/VCzyRaVik+kbJjPpCJw1UAKrdKiHkprtShmXK1KdYURxd5fwCsxfYOJVN
4Xb77vpHwkm4HUcCTdZOHg5XHVD8+wm3Rd7ZjOXfrCQuwgxLp2DD7Dq8/WXhDbGq
b4ZUBlI+EPCoZZoGdhhVbIXrDOkiI6pDvpuDgiLivvAp/fEVgMN6wAzhVan+pZFe
qBJVWGmgsKHcWdIso+Um0b2k1K+6Du0ri+hwSPlPtrV1jCeu0Tr5+jk6z+2+h/S3
ApLaiuKW8xmvb2UGmMVG4PMiGxuzTIWFgvtHtHDg8L4V+uXQ5T8ZzoadJhFD5vHn
flQg2T9iw3dlJfFzqGF/pfZrBQYcbCrmAxYjSGPXP4JEaLZsYwKCKcH/d9sBqAki
yR3OykwiE52T9lu/6uPM7DPaaQY4eSq2hF1WHltHT0S1mMjE2ynFZc57/ic0W+ow
T4We0OeRg45CBhsJ7GWjqgNne5a11T48uP67oykZ8GVMkiXWrFU3vNUhxk4smwnv
brJ5iuoincdfcldeiPTnLFDtmzCM48XhupO47nfHcG8O7I62bD8BV0Lv2WzxiX0P
fLFJtDRNhtNRlbhRsiX4sfD1lK/1s2YCnkt+o/vRgJCFh7QW1WIS0caZe3BK7QGX
JIZdeGJS6O4GOGfdwERVeByUWEx3YmM/BerdTIBZjR47mfFquCoFSBi/iDhx4B9w
v6iOl+O88JEdAMTODkLIy4vw5/jLfgOcxVzwCU+4WzvV4RtOf+0udH1huOUBs+Xi
HwKP7ubJaFk+Cf35Ztx4cr7JWfafX5xu4UJIt8Kif7FpsqeqQnYbyeMeRuG+p4zU
9Z2C/NV96Q+wtt+HNLdB+yvzF4UvhwuOxTlrBdP2J9hgPNrVjOW4cL0ReP/Wt4DJ
FGwv7VnORO3h78OeIE20iIECiEOrjnwXali9fSefmM1XsAXrT/3rG2JvMznbQWYX
5UxhnKouca3M6IvcOlvyBm/5xcIY7nBx/dxIix4DLIUFi2mJG2EzXjzGkBn5IQWm
5WZ/OzVawNgByHey1cZ3qofnJgxWv6UxyUSTIgGNG/9fn8MGe4F5bMY8NP9OS1m1
nqR0edXAnS9g2dZoal2Jvy7GLeu3maEatA/Eic0ljG7Mn8UGVXqW1u/uc71gKA27
SllpyAkMLWqCNfnnrtWDFIyo9MP30VdzRe3eKBvjSbaY7R20h074He3Uz0QaZPpD
1xMha5oCWNU13vTTW0kdTUXfQUnbFHaJj5sny/ucvf/hP03a6qQxPQgNcuSrKbxl
NyP7itdL9Aa95HwY3nI52zKFeTs9SVI3w7ivr/tQtCXO/64YvmN6E4SJC0VIA0qF
sfx6zBIOewxQ/Lna9uyorDPHLit3dKyjhX7GaiqQHz42n6krmb1z0UEh4/e1zjtq
eGSgB0groD51V8C+nFedXn/uvbQpTz5VQd3HcZFory8Ndo5BezodIKoYWMFhn7GK
vJfey5sWYm8OXQs6B6Udqvwka/7JY/5YsUYnRD6nYXaQoiMW65XcILvV08H8oQig
b6JxRQNez4BOBfmlOD1JXCvke9uICOUexx/jBEeLa2WdUaIaEC82B7QJWkMESjyf
wfptOlx2rUxeCxxh6ArhugzNRPwhVUSiYSAM0AyZgh4nWgatVZpKxle8RvrexZYF
I8/b27Rsgt/ZRyfaO1/6MqfsY85U6avyriPkrK0xKDbP/Kj2yq2cow3vgigBiyvK
ivSyzx9TA2uAf/KNTuB63vQtbJZGeiAa5FF2uvYGMQALSa9fiMehNTNtv6CPkMrg
+F6AEGTYxjYlRMK+pacoIeOPpUaDtTyyx4aCPJfjAeLO+u5eKQt7cmYp4ImyOKxW
6ARJJ796T/yXnZOf/UBq1+oiSljySLP382RwFWKd+bspJMsb7F7Rbgh3JTwJRvE6
dVqRmG2Av7cn4ys+5zi3F/RzbUq/PDQUyKw2+YM6bzy8Eww9xSnt12mqoANI/PoB
1j5SX0lJOmn1WocyBwGNI6qGoXHS5vMQ3R3m0oAHRLKmcGa5AXxpd8QVgJ/J6nJ2
gTiFFiNwL6wZcb/l9LXnSxiKvtIpk3rpwwvUaDuT7DNy3z+xN4NkbrwxuR8mExD4
jzgPD+kyIaDyUPUC2JbaRK9a4q/xk82CrHe+SH4zrbosOd3xGm99VSd3w4YHb1z+
8wrmZnvz6RdD7ztIjncc6aFXSn3Hy4gCNF/HFe7yPfDTlEvCsq93frS8028A1vuH
wmYGvnzRKZBF6K/RmpKNMusy6NtXTwCTWfLzofnoNuJuhoYPrMUckS9i1jOu+wlf
fqTZ7tXRR+BA7GmUCzpCr+siaR6QL3ag0M+SW76vxZ1i5x/1DIhTq9UD4nl0nld4
6+UKK/cHiJ6JKIKHO/P1wNawqkmN3ITqIFbPEuKYiZvjcV8l8s9uKNamAuPcmRnr
fO+x4M2X3bePIxkqnGFM2Sve72fTZrpjNK7Ol5vQOn59aJ65fjdsWXph5U5CTbT+
QkidVlF9YrDDbyZqPqWGXlPIjhs4bV7ybFDIBDcfg+BFFI34bgSRaU6niKfg6X13
mESgg1M/mHvLobOJlBMVpQsd0GCPs0vkVCLJyIe7P2x6rl7IBVrEHDNbZ+20P3GT
fs/D+hBnxUYn25sHtzv678gi2rtjDXctYMiBav7mg+QN7m7L6hpyYWTmo5653a9Z
ZZ8G+Dbs9JMlKy7+x+W/9/JmnX66Blhe7Pdg7eOo86P72hjT75mtikXFtu9tmEe+
+4VfE+VK/DCt1WdzKmFz2SACYotVOBNwGzv6li8Fh4XWaRUtb0kxKwi02se0inzE
ZT0frMJvT7/71HP+MZFQ9rgIcr/1ev/iRAr7TOmOcnF+I/KqqUIEAC8xm0EIRE2I
Etkd3EKtA4sV1A/53ykr2DVHDbPp5DB47RCKjIZ3704LzukQIZAYRlxgmoPYUbVv
g9n7rQYi18ybixp6e8Ty6inGDRmyviw3F74QnmYQlTNfSY6iT33pUtYkOpTw4333
sUAhpUWqKAbVFkD4BTqYzxPzxm3lZOBEf/43o23636D2ouG/r2mP+aT/DOk+8JIB
BHmQPTK1sb5AqWOfhM71LoPIaNEOKFjFMkxUN+3a0imPIruBCJLWiJCaDgxGDNI3
LGHXHo/MyikvfFVD4lbD1nqcJ5t0nAAWXzVm+QsPppLxqn7mgoi1Szi7YPwpvDQl
JOqH3kxbrRBqRIBgo2Oett6E6v00Nt4rehI+upFFwS1/PDMvSRA+ty+ljRZq2okF
3le41ukzya7Gjo5PspClv32nTR1oTNY0hq7QEO/yhSA4slMYfILpylRrKTsV9opH
4lhp2AqczjoP7+nuPkxxzkU3whPFRaIlsnHXz6GvQHznKikx1veA1ilxq81A+QoG
8eC2uJwx/zpuYHLweL81p5Hy2lKhRSPT+r2QYJ1yCb+kFRQRYGyxSFxNEBqtrgom
9dRpF8hRC31JmsX+q01zIHgs+rgDtf7DHPAn8G7nmgR93qIhUzw+KR4ds5Rb2KAI
KqA9ISE3pY2LRkXj20+H8Im6+fG99RRaHS/UHORnMFigzoj5/pOeKPyFizjYVxMd
iPmoiEEsGKZ+tyRDsCyG83mcuoIAe3SmZuzijgtveI5IG2fU20TPm7/8fn+xWwoS
Uj9GL4LlWoie7F81rg54cWgE+rOyqih5V9HkLy4+Ek2dxkKvouVLX0kheLmTTgUr
k4sTZ1O8hiuNmsZBfqg/ER+HGdSeeR762I4RYXRVGFEbAgaW/HnON9nNssSDLdjK
McW6oxB5xZmkyzV9W2+bp7IJyhrYHrpnFxVZaXGaLNoJ0OhK9xuEP7/rvS3kp5LM
Hum7n1mr6QTQpviUB9WNm+a2WD56xcHaKyonWxp9aO47Gkj0QP5FJHhG6uQXZ1tx
L12lCNNBasKglPUZN/8qVK24umZxgSRVV070B4OMjKIRfE9f7jUKdFIrXgxdGc+b
xWnaGjrpGjoZs2GkA5U+TSevKuK4822DkDCkTD+S2avxWDVF1CGciv5OQDWh1Lqm
99Wa7d+TR62k+0FlomwxGU3kI22W0wzBjCvVwItkxTjpLjO4D+XmGRsGI+/TEOWe
PPC0l+XghRbea7iGXSGDZykx/Sr8vbjMuNSbnOE6mX0w/yOW7loiUejW85ErwcNO
cmHIl/uholWBN08MRZf7+ChMiWqd4tea2plZL3Oa/7psg35hwYciwlX9JUoMJQuw
YbS4KAzil0Z5FUncZo1IO8PexxbbHKDDbuOhH0CIS8NPLdT1DaeOs3eLfD2JDMmw
Nti8h/K01a7AOZp5i1nGK39m/ca5G1OWINIBKVFNjYR85L16SA+oUMioM9L+p7at
ct3eVUyMucgMonOyXUBsyND3xlQweFV+z+6hs2pDsRCYW8OXJzGPmxYhJqOgSPwC
ZZASLbCCCoIKkvb7CeqVtJMKxwk+bvI0V8bUf2BPh89AjTcH9tV/r8t729BCvRMd
7SbWj2VumdhKwkKe+1Aox2eek7XGuLrN+EZw2GgMBLl5UKqjTVY+yzjEWscJFkb9
rcTXqKLbW3ztS27mYtw8+0VBAoXeFyBH293E1MBVTA5+ccQr1DeiFyPuxIOarFsR
AQgfs8afe44/zv+uMNdIM34BUhAPRbXotGK4WUy/Zalery1ozQGg3h0RPdsEKgG9
pkLN9iJVDraQNB0ecOJq4zE3TUTisIUOVgi1ERBujRrSyxIWm3+nG+rn70H+nOB1
OJazfn+FN+1TpOPWY88DTYoVY4map/mjFHgwdiG/YtTrqPOHsgsjVq/FnY3GKkio
RIcj4PUULlrzyIj9vl8C5G7uE57r38pO8Hx9rtxWWbnFPGeQDvdm6H1gfjvAUy6Q
/7e7fC3TWkSCEZHhYsP5H9SeLAtNDlNA/82Bgi1WcuCgnTSa6ipYA5Omi9gd1x3B
qRQVCEVp+Pw6/kV+zyFE03G9BjIMXz9Wi/8oyMA5rpduVeS4aRVnDPC083EKumcD
exOhAwRAX4lUV+WuD0RFjFRrfdmDivUIHXAU2/cvI8N1YE3ujKjyzvDeawRHdo0Z
OwlvjBbMivDM8z+IhBl+jE7p9HeAfkBcuS0JVoRDAI5ndKvh4KTQLSodMJmimn8r
lo2VS2RxBk8OJhvawk1GMdKeZMctLyHa4ENQZC4bpfrYZPXitLLshaf3wb+iTlw/
Xu2sziEe5zEaDkuoNJfYyyyU6/9SVV4mgU2TR3z+c8TopEr5QJvaLGTKmKCVZnEX
9CXxh5Iix1rL5ClLeREPtncE9EMVYT9UrCQlToL9/FJyNDETbW5uEP9ioihiHkOT
I4kAnTTWPpzP3tYqEgieA85iWY7CPsQosoD0Ho/GUBkNSG3A1EVbSOxAKnEY3q8f
OC8za39+EmOOnmi0GC868EfSKo+Rqy5pvOg64MKC68HFX2Wr5Mm6BBzFWO0zYsc5
H2h9KKL+W7Fs7UVj9K0c5xqw4n+kT/37Sm52RNCUbrmhREEboRaIw/MuH5TN2/Q4
Pywo6FDwSQQDcMgEgKxwC4IUyUweAOvkDDVFfIIqr9//Gy2ieSfzGI2rhwPlXUBX
ZAqER+PIxvOiugyfzOcThxaq5S9vHPwC8vmQu6gQ/HPuvUcuWs2TuNHWEtAQ+Fk7
XHbFSdjKhIyjQ9R4xYpm7UL6a+8dag2dJaMMKuMbPpiwlLWqC/YFmuCmBOAi8a7o
+1lM30obMQtCYw8kD4DOiAuxo+wXILfjp6mMwRuiETZIv6ODhKscSEHXg7l1AS/o
oGtPzn1IGy/o8MTqY7D53QQcnMXsJLzbVLhHZPEYvKXGBAQlLEJk9vXpYlVs7yEk
8DNaSNxIrPJ6QtB6D2pEUCnQYV6GbivlSx8mayqWkzVlrcjqFq4SUtVw+vNkGZWV
TVf7ApI86gw0HMiMkyOCFKcZVEcQ6nxLeqxeefiw0TQMFxv7zVhVL7arSSd2mFz8
CRWVNHrmAnih51erW2cHuCS8kYNbEHjDDIIA90I3/ktLnaragTTeD3y1+8OGQ+xG
/FuDW8mylFyCqDBfkaXBMQ0DaAPoMfsq2IZr/T9nvZu8tOiukbwReb3O+r5mvlFD
RJSxQGSefFWbnuZcOseA1cj+tjs+ORHxQJWylSatFKW0GAnSY0h6LBhnhfMZOGRT
X54Cp6QWV1f3Pk/GXVPYBTGazpK+H6XGYAS2nznVK1KNvqlqGP9n3mTWBUcqJD8J
aG/kqlDK3QRqvZwSPPz0fc1Adbf+qqPtPfvvAzZGS48fV5egO/471Ln2fuEzi2Zh
DFuIV9YdcV322sY35dNr0PbB16SJSHsPEXPoVIgJknBB0ParrMjbkBAyDgwec7lY
FmrQhwmF+p74A3sMzSjz3upik+SigHoNgpbmy43OWDSDO1Z5UHONW/zatYlKhlPu
ZyDKy8u6MSs/jsokichbdnG0byPdyEeQkerPVjoPtjjAwWVxcEr/WS8rmnE+a6ot
7f33suCfGPaAv6oPrhxA8K/eqOdTnej+EFWvPf/CxBVDxoyJ9v1mb3O/0h6J27K8
biNUQJ999UJNegORxQZyn5TgbCKdcQN5gjx77Kc9OlNXECwvEXeUyWNHc6fDnYGx
2VRHhasjpvowYMrX66HX4IPTH5HY+kdv5y1kPq0i2sCXUk78COpVbXK/uOloJBzs
MXkZnqzml0e9RuX8BbWJpVkjMgo5hVQKBChOYn/fo+OYWZRdir0KoiHsvzFXbY85
OdNYTyf4AgKlhytwRS1wxAEwXRxedU55+g4P0pf7F0OwMh9toHi5d/BuAjDNyoke
f7WX3L9/7ddX2iJbGGHqDJCuoOa34mNHggpBWVpFr2IbDhbPXNADmRqC7JFLLkhJ
W68y3iTvBK5Jg4KyJzmpmbAGSf5cU/OeOqHpXYDPGcAMEt1Gnj6PZx+deSiewxzK
92xYdLbdkNgWGSAKY18yjv9dbGAdguz9ptZrx7+Q12S7YfrLnZTmsMaj+PazKzVj
C8p3SnftVcXbk3Zn2OdWGAYg3iSgn2FKXFid+t3fRySClLBhAKn9CcWt4931VQXG
CVnXAwat1yvv3dUGZzkxhLc3wodvKqARg4x/uBAZoFwRts38lZMY4PEa0Cdt6vQ2
aX79RmoM7JHWBtk1m1WREUOEHxFSIThlLftZJgcPmMKItJNAQ9thvt6FEMv96AWl
UgGP2IZWy6O90HmB/v1+DYLVQTHtMa4sPlFaYSR+/3gVBL++yREuNczHpAGW6Zuk
fqjqRWIpK/pq10EMrJ7JwVFzWfYclQoKsd0LvQAnlKEsHg9zWF85GNac5yyH+rC+
CSHjHClwZBdp5UXD/bOJj1w+fGW4Fd9bCqWpV2chTiOHHnW2JqLUJg5Fs6iINRkM
PNl22ovp4mlt9TRm49CqPj2dP2Jq9i7MXbPwGY7O/TbeHcRcu1KBadSCgcDwP+TC
S95esk0FBQRvfjg7hWgZS1LDvLP2yznGyjUmX4HKFJazNypHVnbHSt0WaE1cWoaZ
76yxXwlQedVf8MbYCLqAYmnWZQKLXsLYYAaQls82p31h4yzXkq8RaDqM9oI0lwha
uHw0i0mxKbPVRDC6Rp4zIMYuBbirtTw8lil+cnFpuW4kZLq3VhogivGWnu2RoO9G
XH2HEYrYTn/O3oU6VOr/c/WJRNeLnr1z2Ivz7hyhQh0bjVSLfeTKayUF/gEcwt6j
rJ96V3Lw+AxajUtSkd9gniyfD41sj5ghZo+9p+M/FwqCDyy8Sg6A7N05Nvkaevpo
+kc+1zf9eU+EGaynmwW0IroEXe4oLzbh5l0kPfcwZXeMYcsJl81JJ1TlbUByYduv
5cE00SZ3oKkcJHOQImLn/ZLZIxSlP4A+BADJJMC0yAGtoR89cRM5RJeMYsjMRA7C
/izmZUeYi5HLvKpfR7vSPLVYby6PWU+DYZYbVWLfdSv1MPaaCLnpmWw+nyxJ8uq6
K2h7wlVtT9nnOGXstlH7Z3rviPXzIuo5+IJkGkbW1XKU5Bhtz9qiPwurDHNaYTYI
DzBg5lSywez7gs1bCQHvGinJC2S9kCBrJ7TXrZK12uFrxAZd5nnvQtaRhW18bKnP
tEdVoj5A7Q9YKEVAfN9TauBZr0RcCJwurjaf+/l2aaEvdjyCeQzPgZzvcW1kdXOS
yQZPbb96yNzzmE8c1XHPnistllxHFemOaQ9kwCa/SYSr86FetVv5c5kTFgaNjzDp
IkPM6uO63UVPzrxSKz9ukFn72GtuG37TUaMMdFpSe3VSYHL5Aus1sILYrmyOovDY
eoTCIfRkNzLR0hZAQKc+Bxc6RB8HldGOoLnYhcYtb3bUWW419oiqHj/QqefbiFg0
a50wp4J1oE0woRsWurcRbK+JIkTaNGi+7uzTX1zpqfStvfwczOU5bfE7eLdF+Ouo
9CDzWX4tAmzae/N4x7AxOBnl25xjzvQ3ZMsfifkR4jpJY0I6uF54v5+/S25TKHmC
M0WYWbU9774uQZET7GzW/H7PLXBxIoid1pgjAQGe2pn7IQ8K8IIyOEn4Zmu2Fhth
RDlwTEsdWzp1WlmHGRzQJ2uSBowGSDUkTkPg+pEhVOs613CX1hwDV8m/kANcTAjm
10gbhM1XB2fYMUQgY9WbWp0dcaOL09MHZu6BFiZQ92LsuyryeKma2UY52CDYlfwN
SA5wiCVYe2Bt9geATNL9vuMC85P6XEcDjPjn3ZllCLylefrxh2SMTJ49nLLyrsPq
Bb8IGEH6hwd3vuMTkzEiSwOCMFW3aW9qdADm/PjPqa25xnVGfsUduuH2pEAeKMwJ
Rn9/u8zZKQ12UonljNrbLiWhpnyhEQyxMJlU3MrIYcAhxvikOnud1SDt/8m20p83
Nm2jwdoP/KPNGvup8J5ADz4fy21fXC5yOwCmLX9TL/zc6D20K8b0PfQTOBwQAJNG
MxWjhomxj+zVVGpx8KU1dD7DQw8aSRQWV1mkObAYtaL1qr0V/Bdc7+S5Zy8bywbS
fSY6FLL1DtgW0fm8x7YubOfqsf+YQkq4AjxUuyKCiejUyJKKWMhgISCgCZeadf3e
pBLJf4tOd95OcazmTo3tpaEB6Sq4mT+XiPR8xbQBSysad81L4DZYMSyrfukZahcu
oku64X56mGa0W42AXhELgU5FHcWpSrt8llpEEJz7CCyLG1XzwpZ3d2PwHhJjNP8J
s2Ocu7VS7TLW6ccIrM07amiMyQvCOS3nXIbdxe4/ZW10kT3jVISSQMTD5CWRqIb/
+ClpNOHtV3YYEF15zXGpurgNJehkqYRYM2g2Iy6uLEfMtjbhfw7kDDudOCsDTGMF
AEW4zYQEsMV4NCcjgRqWEIMBneO8WHhqKPr7jnEP+mvhTETpb+tnRJ+OJrT0Z3ma
RqJbdetIdei51xMnOmLtXJnRRbuPryl+g1YhqluNh/t4sxBFlO7DrI0CIt6yhMrM
vIgYJNQ3St9QzcECGiQ8T0vybdedwGiJvnYrzdFIvNFMTlw2DNfHMw2q1y9T9905
WiVG+hpRKmITzPYJ/Mxb8bg02hoZ1v07UZtoeqfjJ/3tExOm0P1TxEBoMTUWu91K
mKU6dremGHygY65aPqjuq3ZPJPGBK9DcHBZ+dkSg5UPIa6yQqD8PT7l9ld1yVxlQ
wZjAku5wXz234nqW5hmmsIBj/N0GedrWt3G7g4QtDT7fDfE3f4OXsvhxgUhttWYi
7r2pagXMkoT/Tt2OYegvOvcNGA6EE5PifzpK12FMLwohbf0Fy5wxBljm4XKrvjvP
GxBEtC76cSyEGpSJ1qmB5ki18QSHnnv7pUdSaouCoh0sXfVUL/EBuWu7+HskF/yv
uJXM3cfn5izpeGG5jsIn6ed0XMXqKirfPO5psgRdWbBtuQl1uLEAGTSptOKRwPai
G0JDmZ96dCPH8wsLg7ueGgWtr0wP6zubNV69OHMnhb4RmgdelwbDhEZDYBMsmw2E
ODrTLXy7nbkxug4si7XV0coVTuKwviffVQr9lsQUKnE8k8aCLfb7J6gZOLoTuyj7
pVRTSnp8qQC6UqLGgmJfFQjuNdcswq/ijVowLG7l2y8ERWNcSQmr2z4HoTwDwtva
QMbzQ2Akm4sf3UsVsMV1D9MQbhNltx9vd8Ix/XDMFpHlpmudqr2az7o+JWIpD41k
rbp83q7kksc2J2praXkk4LkO9mMutWrmWwV5j16wwDGpsJZHQ7ZqC27vsRq/B+cx
6vLTPNtn1SmU4+DNF76Iw/ytJ5sMPhGnZAYxQEe9Dyc6+ncyJ/3dFhju3Mdm4hAf
XvWRY21hFGVQL8BUft/Wqt6m9I6IwtTIu5EFWaVsrxrQ1q5NdxlHW/aBpQtJcdIB
Kbpzm9o4PJSiTd/yDTi5UUwKCNwIYP3UnFnKpSjvvVzZ6n1zLMTN+xnh4kF9DGA8
eg2t8QnOpbzaMWck2giwpgNrU2g2SPwRlZS1uE0xEBLcFDGXm37YJDEOxL3K1wlI
R1oioxvs1KbB/WF7r+b1CI7RohxXxxDLrKGdemQciScQl5xSdy9xVe1zVeMv6v8F
jNnsvqufxydFhnzobUFMPfIHMZWb3A3Z3zufnhkLRjFDA5Ypx4JCb3Nnv9UAW8h1
kpUCAamyNifDh2hathln1tUCSrUeeMGh0MzsATcDqnvZPg/3CnGPmAiCUTC9lBPL
xjtgc5SrNspIuDv05gk9jrnXWfn3qvLYoF0ukEccDcleJBvXHihOBb81446guGqt
hbBBc6CQNxpzoonYONeFii5+9PJJ3D7s/WNZ2wJ5OPG96Dt11u3KEGbj3cjEZC3b
joxKcHj+bHsx1M6OeUYdFdiqZf9Qis8RGaztmNHQBKiGkuR1lCGvbc15Pn4CxlmC
pK8nOnNz4Y9jX8RIDZOz4b3bsp/xxou6HLZ3UsyMcZ2L51MYfXGbHT4XeenkUMKl
XEfGUbw4ABOkeLGp/qkLW0R5lNF5FpJY7vE8AxS+QIB+wqcWkSAZLgVNmmZ8cLxK
iLwvXzX90MoZsf/kIujEjWPs2xX/GRmxQxuGBcLAYqKc6KYNZfXRcKdRElqB6Uo2
Akzd/yG9mb+9VfyTRHjnph+cIFS1JsY36OGCfbciWlq9q0WLb7E1HSk9+UDvKpQu
HDIQJU/+5rs+tGoOGphzM0YE78gKw04VxeAhR/by/4xPAOuguqgMq0xqBF8dKqfJ
rEM4CatCCTzK47e49QBGbDVH1HPuUv0pu73TLuPzrqiVw93rDXqwx80+FcUtdGcT
H0bucYYNRhQT+vXWVqSGzBqogR9P42naFSlk16IdEeMHvWaEexU601LIwoUYdKw5
IdtyluhyVO3oI7krZ64VUycouGOZUY348bV0yN2dPHphkQQEhGxJF+mm2DFAIqYQ
Gq9tuTmJvcqr4HOGFH/opnCdsghjeXMADttiZ7L8fJXAW7c1yjv7AXU4qW/YrEPt
LuDsS+PJYX2vZXq471KsHRH1X/sKBdp1pjeijmraZDY1cw8FaA7ZMZrQApx3nIyu
kfyzE5q5LEiUuY2kwEbiljqhqUXtnpRr0GzIDcyggkosbJ0k7sFROt5F/VYfMWyv
XBr09F9b24iHeNJUq5SKDm5ONajDyuIPvo7KpkxMnySiOpmP6jCO4Rg424ogCypK
65bxJktD952BzICrYJaxYqSKYa3y8lzIYnzr0qz2bGqQEmze4/PhQMt7SQ/Hcsog
Nm87uWxTfYgp5DQKKSKz2QcJf3PJQZZG2fr2dIEwMa1CnSPFn/7myvGZxdohIjUz
214xAICB27GwZ+1TmzgC/ESIBskqXCvPSxW5gddsVVRhxLqWzSKvwnDwipJmt1RZ
U3MnCaCDxWD9eTgxNfvi6B3Ke12gl43wemHVx4g9LGSt+JlBWvmHTp1RqHx+7EtB
fdd73Q0nIJqxa0V3NcxbvMFyXjUtQd40XguVnCtZ8CjBk0K3aar6rcQdx8rxT/md
zNHbbyKnE2b1RzVstzGeGwGpbpHam2BrwmGKx+xX7U7YRT+2n/JktpaYA2UreZkf
BzHdAuhdTASuUUIVBqtJXP7b2Ln2XwtKNn2Um0xcwy5I5MCliqaYFrrYkY4rhlfI
WAJm4E73Zh34SymT5AzxczDX3kffMC6jbU65h/iIx6H22v3YV8LEUMn7rAETEfec
04xaAsL4uuTMdQY1MmPfBIf+DGj2otfQRn9y0wdhU0rDHbgviYDWxN9xZJ5/aGV4
2FUj3BqhVx1ZCxfiSq6GzM2JCrufIK2b4H6snZtlRzO80ERVTmk+tv+Xr3KFnYRe
vT3NXNKEjoO3gvspf9FKDVgcWiGjCZr/gwFrNSBqr5rlgGhkQnkPDW1dtKw7bKIq
9xepcWeHySmakYyQ3UcXJwwvm6posAksfHqDGjyQFQ3b3vdRFPXWaYD2knY1bX6Y
DYRTp+uCr1thykaSk7Z3wUxzan9LOflG1lxqPHXjQGLbjRjJInKiop9nI9xFla4J
tWSd5GI4v59FgrwLcMqqFet+shISgPwMA5hPryCN8meD1P8+wpZtbuJsrskuS6Sn
EuK1PSaKdvBX9S8yY0o7f8jdxs/qN9/o6I72EPup8cThbxsram5s9TwKlvgbhFUU
SsBxkWGA6+42hSFRG2Hl5sNNF3GfbpoYcmBHd/A9LZpKDwIU3IgcoX6AtkLCQlyT
K50BYRSsNTVbVVo/CPoMqHdkgHGeo7NInEZIebkj1mjhtmuDtYd2OClJGK5m5fMX
feFYtoPIcrZwEk9mqOcewqyNvIBNup6Mz7tZTLZD01Ggjm/4pG4jC2hr9Ijf2TZM
rAepeUXIBrpJtT7ovoPhUqniROOcStklTtNi08IoVEOlsoA4ANuu8m8jORQEXCOT
lprGZjGxfWxMQi0VrZr+uY81ZCcvqqKBhcWXkX3kg8ZghY1N2yaJhsxYQwwJBrzh
tqDwyFzhEDLzIgsrt3XJUtQz66kxtJqYQXARviSJ3iRPKkAXC7J89/AxBeQgOhZR
K5g89jN439pxz7NMOLzpjv6aBA/OFOt5epOzYoBm3XisIZ7H1O5alig62a8jk1GK
B1FbjXfLmUhAuaEI6w9aHDDKeKntHuZKdyiHs5Bt7KXN43TU8PYFDlgRJlKErCua
fBddxWGQyN47ICBQu34x7/LJFBMOWYIA4P1ai38Cj/66kJDgpk0062VVy6oSzbBK
4mwLpbm1qk7XtXCqyCRbvEoxuE2uj3SREoASP9tlKZ7W2Y5cXL7PeTkVPl+oGhh6
mz2SEEZKqvNQg9igWoGwi6NRYMYfoyw4iIBgEgZ2/MNJcH2OlPLQFpiVHKBDpR5q
7PiS28apHmSLZQKk6VX5pRLyYfeCnOIEDs22YOIQw8TcknmUvgLJyO+9nVaAs5TW
J3NT5puKfALBOemnDHJiUvQheTkveb+kZ+g8KQGmOAySUxb/y8WvrRIzudLw3scj
r7QWix/EmlmQR1ImBPIhj09BepnEgox18AqXAwRHdu0QwAKI4Fk0UOfZWhVYPNjv
Nbn+yDJakkVMBdlYd8J/raZd0Vwtk4eU9IFH5akEZ+6aozDnvHgQEDjpOufhezOp
eqePb0YbOPbInYrwkMf+DMXbofYePnPZM/P0tFlMcbeeTklCkJu7/khwoTsDlhgZ
oMTMd/b7D0niB86j+qJboe3ny/gT5+eRsULzAGn1pMO2Jm5f4tSbc5jtKznr1pU+
7R5GeNdWZQDjfSbReiVkzdKyKI5rIxMV79cUg0fgxpq6ic74LNUUeSRk1vYCGXu6
VfQxNAa/Nn5ezPlWobRNhjTubTHyJlEUWy9Cdvcu69Hk43RIq9S8y0QCPDO0McQT
fFnL57WTIdoV7K99KyTSd5a0B+DubCcBOMcNSXzOoKQORhZGNFef2JhbMdk6zwWm
veZ+EG53CpwqQ6FDwmuXBH+m28cUHULHiE7mhcPb9r+1Fi7If08vNyZf08/evG9r
65LJw/NDTbBwhmc/McVHyJhUHQDw8+ab+Jtd07amPPo+wcZ+P196m969sxUq/oJZ
SfuUJIgsgajZGDxvGbExSibvj3nalIX0ijx2Wqg90Jil4xS3EHiK39dLud8u1FN7
LZQd7aQp0HdaKRO8ed6/8ZucWyuXn8K0hOHzxsj4SLOUnFG4qev5rJdvsFPOpvqH
ozyeEvJoHPjGZlWk5oe5ErHrZ/FLuyVfSeoUOitqgKJ5GobUPqSfLGkoiNMArPWn
7FcQFhNJYeKHY9FZfeInJE1VnUxHTiXvY5gyzAvDg4y3aQgDamkhHFNXd4J3zpRC
tJNHcuEqpFrSX8Z1ClYNPVxpNp7nVixkqaQhPxJ7UxFeL5tk2wDE3VPlwuZLaAPE
AC4iJ7O9EvRKBe8UoRR4DB2/ZOzGdwkvtSra3dt6pItwK6+QTIAdIpPZzSymDHyT
EgSufm6g4FVwOgI630Pyei/ZjU4FiSbJsK99tFvWK6C64RBhuewHwhzvliQU8auH
APDOHgZdYEC2w3/gz1OnzIV7wu8aC36wdcVgP11qKlfPC1bM1C/x82RUFNGFpGo0
tZeG8JLuuorymARkvY1uUAMoaO1uLG01xgiZusEw06iXJPW1YBfg7wrUVfoMl8Sx
daF+Bt30v/nGamYI/vlyrw2r9alRcapA+G65U+kMuPOEZB/NqQWKywXh5/ryBemy
MBIH/JPv7NdIyHWIsElNsv/3sYqFVwR1Nmy4PZ9/9WopQ1v+5qJq2W7P2i20c9+S
tKY5HqAFwaDmVbgZwNacWAHvjwvweByGZ1GY28t5tJlbJSXb6/I0sU7KPnhSBGV7
l+HXatssTbs7EWl37G2A1pzApgkbFXjAuv7Vh3heWCUPrqRw2IuVS6GCZVWOS8TT
VDjUe7e3FXIb8/RFWVxRCM5lb5dWzEq550+aawjsYJ+QjkeL5KuchIAguXwLUAgE
vgHKpnJlsY+YYaBLjwmd+4auBucOhhNHFgk6El4JXsKoXirVL9Cttss1u0qFOSWd
pWtT5ciNVF7fLBwMNyiRkzL1lgjZy2LK5+ZVdDjekqmAHRrTzx56xxti9sOB3rad
cNixxaa1ds/soFQ8zH0JG9TdplBYquOTnUMEQ2HD0AkZPGgROvnc59VqYOKeht2z
VyUUTFngd5p69yziOqWc8PvnjWfm21rm8yUBLVlvICyylz/cDk7HE9US4lw+tkXa
5Jq6tDGqlDse42r6xeJ7f2aTFfRqpmY7MRCVdGRZJCu2u6HufBkm5Ez+kK7++E9x
WUCzFrZoyt08j8eGJt5Xh5N8ht5mAqnCbLLYZq9PBukDfs4x5OYbvGVrIKc3cmXL
fmymYcyUD2X0Tt8pycoRIoeHOZ6wJWEk3Qm9mjkkVMJoIh6YbQIQCJqNjDxgYgmG
Ya1aXPXheQju+eJXUWxUiKiH3NHbnbEQm3NCBtQ+z1+f5RH/HoRdpK5BnHaP5hZH
3n2GH1U+vCCoBu5wMNFAghmv3fkRalruZgqZG/7sEh+rXXhy5kaGRMBp85DhJSVm
UtBI2hyk36onQL6tVeOgVSRN2Mno0juPzRHuLmrSUkcjgx2HmkOqcCQvkKY8SuOT
W7YBh8VZZCIqYp+KRgaKVvGKbh8dIgEkXgI6Dxihmc6TRqTq5WX2S5eyEcINjDON
tqIRmeGnLmmzZfd9gJiNOd/ieEDt7dv4IVOcm4FvfwRaypsue+yOij1mUjDs+2qU
7xaHnVTcuhbi2A4zoDuvOGGHu58BmGd7oS1WyaM7VAzrIrf4kIhKUxwL137XeAU1
q2llkn2Id/xh2RacoPEmxVqpiD7jBlh/nPCpxMxZ6U/e76ouFs1AxeUzExi4Tt+E
oQ42gTVFJhqql44jXJANCo1zF1xOHyiW9odP2gl6UlKe38zB7DwMFTVgegOA2XgX
wnrrT5wQ+m59hKN9KH4fsCHqpVpxNSF3mGH8S0TaloW4P7caR8+TGmR4dRHhXWkM
IDHvb50iHuslvTmfkpSws+TzjAWNOAMnT8yjXLWSoHx33HZRkVlck6BoeS7E2gCU
bBuMU9MbKJfY76gfkc5eho9V+7QCsbhQy7OHyOcWx3r0HNHSWMLv+t7ieo7ZD4/z
DCUBaCQWmN7RDQ563uQ0Qiu0jSgroT91iloUo4+5/P0O7Cv19UPv6ByEOTK9jwix
PNMgcndtnTR4X+GxrFqsxswnZ+/l6Oy5EUjSkVnIavxrF7Au+y2tI2sEr9HjWfko
FmYIoh3wgCgDXZG4XKBvIqsUT9oWc2mO8QyZNK7sy7e2/kjptB49aZHF63HH8PIB
KoS20sfYbh3BIv41GfvYy2/qD0I/WPAnAVhARbuGXwzt9kEA2K6bimjN/cioLWMG
E4Lg2J5de6rjfdbN25dPl4Ro30SK417Xw0Li1W73RDU9PZiSIVZdWUGyxiHK2YMV
5Ss3JczGxFAwm5GB5X+dWTyVtNTp8hb/NpHGHte8vfAFsxwdy+DfByanFEBv8iD9
PJyW/cM2Yvh2F43OiVb5IsPxItwFmwIfoPcIfBXLu7ibheNbeDxsnGaU5TwCZFqB
G8tLV35pIKpUfFIzZabTFtNK0N+lXiNKd90g+e+UG3CSYc2jClcLodxcL2pfWxcZ
JfMkif41HpkCEzO7C4Zb8SNDwZVSElSSRb1ReD/SD/KGdxY1u7DbK3L/pAEPvA7A
hEfTlPSDa/9hTRtOaedM2t1Qh/g6uIQtfO3Kb1LMSAMNak8Lms1XptduQ0u94FT3
sFl98f+SyhRAvoeqKI5tayNym0G+MY+NVBqmfD6v454m2Dsfena3l8eUDbU5m8gX
z+Pf+iN8Bf0IP8HcaF2lCuycumV7WDP4Sqi0WMbUYkyiWUrFeKIGGpNKJ1fylonO
w4mfgHA6TjWI8jk8CXKPda1/4IjGpQx72UccYNBQDKxH4hafXMHGvKosrdZQmtAa
Mn5hzB5i1Br4n8O5wlWINwGuxpjrgVghx8HtPlsb7N4sqpgo0BuT/FaSczByeu/S
lndbx60N15mmYfFFO86sNJGnU3T4+0S6uz4vYmd36ka8Eu3EbezLpFLb2rqTeAdf
wpUGQmmnv2lHVfwQwU0jUQNFP85wUuqVCKCjK/G7xE8iCVV5VEjm5n30oTw/HQRA
WOrmXyahVFSvRVpHXiUr1+ncsTUnXQW8fGVIvScGde6a5plRePmxtHkWAvl3SQjP
3RR8gqKu1tMBNTWiwwFimbMHsv8ZJ35W3p+o8c29RF8XoYn0egrydA+qBrEfI2yR
RLFM0m7k/tqTjHTw0xL2sPJ6DGrrgWO4YE9CqRRJ0LPijuZJeDPRWfQqbSpYPrBQ
/s2FNYkBqpWmCjjaJMnk0y1HdggSmJbrZ1BX06e20qpOGMSC033rH/Id1E+1eAlf
aJt2YP89TpFI7jjNt4ULgn694jKrnqkerXLT5g56KqgcTRJCVwiH+Q3vgerH6ff3
HVtfsD+/k+/Xjtxcm9m6lP7EbzX1yei9sBqCdzZgeJoGCBIk5byqY4PIV8Dvi7py
wlT0fZqGIBad2k8K1SYCSUiSuamvULfP/CxdJlfNPCXuG+18LsNMcRcceqYJFggG
pa3/6Ge0nxQJ5iOfwVRzbAMDMldKx5usSTpsgAQ+3fg/7H+RKOuN5P0WPe6ocuph
n2dVYmfrHpKfFkAwvJ5FiXanHabJvjBDLJ3K9dFNJ1Zkmqz+fxv5WUOAy2y9Ttxt
tG3MdufEF7Lu/HlNeEIWcqlbFmeAwOOWwOiekEBwB6UGYGE4lAXMMAD0x6ukaRDv
Fw1QTekEdp/OJnKsJlr9yvEHb3USrMX7WwR4VIGPMwfxHSJ0sVIWZPbiia6pS2kh
0Gdc3ffWn3ey+kmzAyP4jaV5QDjboUZnZlZM9iETR6m76nLvI7MpbR131TYtmrhG
MEOiCZwpkcI1ZTqWEcVUHJJw31cjakTmQh5ksp0/SgDeNjUPP+gbcEedH+nvd/V5
8g8XbwHbdfqSNaGvUXy3OegTtgGfCX4Ztc5VhsxxoTUczA0qQpK8pP3BOwlVrFSC
dDxdfBhgAEsBvIBF3M0GitxzqMPc/192gIQsrcWGRlFpcYua3nJJ4wShJLy1cb4V
ex0GVmUnYWwUA1TNPv6ElBYavd7eKsg+WWf6HMgTm9gIFley3QJMX9WEjXRNEfcL
qkFoa4S9EqT5MuNd06MIshDukxMf18X97is3lJnNDl58pHFFjWuIt7rWcLLH8oj1
YHhJh1pPLdEPvgVs+SethY9g/M/9N6Sk7Qgcu2lN5nZrTe+zeaqrNKZ3a2/bwEaH
FgroqqHXhI2LfP1XD4F/NiHia9ekcTKn9RBswkQvM3eiSp1Z2VVD6idM5bpitWQb
XG31PF9+dGuUPBSbySWkUmPVbB3uGZxWK5GUruGEE+p86yMeh6mczJ76n6JNaHP4
0t8KS1Sj5G+m61YTWehIraW4mllP2ll8KPY7xXS7T7Cw3F3lX/NvVv03yK7C6N6y
Fp2YPg++h8gGOfU6vu2sX2We3L7/Y2ho3jELW3tRHaaeSPUVeOZzBwJcCVPXmrm7
0fZXMNjtzKgkDZH1f+Ep41g0XLpzt8z4Mf+LHuouPjTTtdltI9n4etjz+D7eLoKQ
I56hS6dOfGCcxUUIqyNM1rrb9kfYyT8zkNT5cRzUfYt3oJgrgqzLt+3wt/MZ71m6
gXGok3NYvPY/8d9seNHNX3ZO8Eud3N/CH/spLVpwGt2PVIYRZX5Uqn6mRIbdbtWu
8ADYV8sFitrQampJNexgIcRt9ezcjz2a/10FQoLA/Xa/ltBB0mxVQkU4Aqzo4Mq/
G4Zh2Q0HDko6n6TM81ktbfQyMayDlCQYjnKetr4yiJj5PBdII8dsT3b+REsMxsYt
6e1rsSXOe+na1K8Fy+R3k8TAZlcZjPhL811hj3FL+grPGM/uV+yEHMVumzJ3z6ob
5NDKRfxfzLvr7Gint15LNKPZpB/e4rihqbG+wv1Ub/3g6YkeCM7s6OUq+9tfGhvl
vQPYswoHk80O2Hrs5r0cXRVT28hFZzKJTcJYZUKdd9Op46RvLJjKvIXXvHyZ654n
p7N5wsbJi16dzbWcSqV3nWW3+TkUDMM6WNU5kpyOPbGjzMvMCzryhyjG7/bcHmaQ
LifbHJEw+OVPHMwk+udmiWekJUJI8GUlu5MmxqgjbI5j/GLWlsGsioOH0Zy9jrrS
qLdCaG3FhpFntXWuKcBgduleWORnoP9i6xnVGnfYRxZ14pPtz7VUTyNEhf+aRc7o
zRlynLQRn7+udulSXi7WtLHo0vfuYnozN/q30CqRMRRJu7WGWmysYX/eOPFw64Cu
BaH7wnCzZdZQo4hLyfPVyF68Fh3uMOIws3LtK2s1uJaRO8J9kLrLeUODjWMfAJ2l
P2HoM4jqtcSd+9bhGoCwYhB1ig1bBVZGLXaboW2PlU3hmtBzJOXTdsmySnTojk97
e7RBxla/XCBLIOz8vT5BmHf2DuvnajvaSuriKmcAS75aZ2d/imi9ilS/nKYQWuO3
xKCnFGCBduVAhsonONcSxfZl2mRsGlODCunEVKGdAwPH3QCTWWI+wfL9VintIxge
oWW1+0TXOcaEP4qmMjovehXbYI5z8a5CodQi/SAurEEXy3Z37tvGiTmy6B6dJLLj
dd1wWmjtizMNSMMU0dmNdMC8t2rq1cl+usZbX3ux+c23GBEB9NJxqU6A6usSYP4W
IBlQy5XIwXZQEkNN6EGBTNKEHP4dePH1860ISbIcOzESeNdq48hbfwcTbtqVubSq
4ghV26tS/NtSIgciNsAnoOogR+Svynd5LL4d9607Bz/p6Hs3wzzc7YhvtFi8OcJ6
snKN0/nYaOIJhfTOsNQbpZxnvWR3mh1j5VQs8C9JzmTYiIOlUGSGu/zlc86SYv8a
Epmq2fiyzUdBg62643BZYmx7eZ2Lc++m/Xavr/dJRwc5OuOsE2THPXT+VCoJGTRZ
R25DMgx8AZbgCFxp0OQEYlRcOjkalTQdj/4j+unA3D3uZFRKQSTpKH+RzMYCEapP
hvrrH+JJE3YFSMDXcdn5TzHdfztZA4MMO+VBbh5t8tVOKLcA3WneR+TfkV1u7gU7
kyczC0LIORBmHx23dbxyQcrKJKrU3JZuVBZtuyEgI1AAI1BvfsE7R3iNNTc0KH+W
W3+7uzX75WkHUBmFXRFJVt5s1UBsRQ9TfUHwHBwOJnP9xTA0UFnuIXSIF+dPKl8M
ggx0kRg30KgTowQDSNODicXhNzCJhUz57Z2x7dJEsLN38hnvZjinBGdYjXA8LTuC
FKMM9WuCiZXgXmIRObXUigxOkL1f1PiS6XazChBRFO09/NFCijhS7T7QszvuwjQ0
yeKstEzM/E6+WyO/9zStjCvgCfwkjcXVslC46FwERtVw3YrSqzLGUupBnf3ZbHhB
sZ57BFVUeDuxhKQ08dBg/wV+VYWcsYiEF7a7F7c+Sbmf694hYOGSe2ysasW2wBZb
vtczGBIf1AAo5Tu8VV3asoRDTxgQ18RNnAWNASpqmgrLOgw1ZbJN7Avsb7Q1gDbf
vTmt/ZR1PkVeaK4JkRCP0Bpm1eRJNX+xxqQ+zKc5+8BVZN0noOTLc19F/4REejuM
nKgAo/HtUG7UdG++FXzuteibkr6uHtMP31E8A3reXIG+zFif9KxQtRZe0wkZIBlq
R2OsnN0LYF+dg2XES52GvFRtme38LFioLevHttqXimNbqDHzwSIrGpKCPI1Bs9R5
S6huDqrkxnIn6cxShkOBl/If9Wx/HEEcGKSH12/oEapN8hEbr5AMvDaKAPYGzoS/
dWSVPf/nO7V4qm7FObGAO79SGg6hSgx03LQqmYA03YYsZucpcTPzeCImdTb4QPDE
76qrnrdfVXxpjE0Emfxrz2FtjL+aV+qqoHz98Gp+KOy0NIxqJPdJhmJBEkp1+X8W
wB6Hrs4QuL5lJxI7ARIfjASBB1H0JCkO3+OIK8coTnGw70cNJm3lLrDhWA6I0mL4
3QzdWGy/Yl4BXtJUGejI5UcUSeGoT3j52gks0z84XZaZG7MSFWJYdwbW4JMCqG0Q
XB2OQ54NXVBwQPqVW4N4cfBXqbCYYqvG4Vt4VTT93zylyoxUEnhmlmfP/JYs+KJ9
x35VXQPt3OyZPa5J5pFyxfswiKHxjbnIBc7qTivIleCeLy2OW0eljqoNIyeh+DW5
9MWgCJgW++e5U/NSL08d33t9QkBbA0Ueo7Y5D9EfwmQT4RjQkI/jE5Ku0fmEyheP
nchwEvwgef3VDGlexSHBYOF04xvQDfMatYrFCfSn4gz5ib8nLe4yVgA1FbCfJPjU
DTbXNcCW+CRSMkeuaHZ1W1d/UWGnYugsKNGd91z2H/rsC2AOC+mys/Fsfsl9SVrw
otWWe32sjJ4qPaznT1HTFngXWznowl2AdS+tY84AUhvtD0rZOUtL+K+sVR58zHJP
rQfAj8Gh0F3G9/J2HoLisPmt6WrxQ4GYyQHpp2D7WhEI60S8qWKsJIletUCU3VyU
SkrX5BEe7MiXWDENuPOSvuB5IEWPMt4UZfQpvY6DmX+LAjO4QxiwXy4dmKSA/8/T
x+Ah64TBweMDlerA9e0xtAPM/P/7DuCuU9vN5cQIg6fBQN0O2dqmriiQX4FE3k6k
lk6ZmNsCGOLbof1MyG0m10EqKmMpv8qHB/V+HtEUTWCxTCTYuydcGtgsDPoTQhK7
UVlLQDt5vdZUt6MRAHS9KRr4pkb5AXW3tKwTVvBt44OkYTeMKo5weP9l4Ws/14sz
mJDpOdTEpBHfxKkgIgJkDnE0KGhJhyvNyt2B4gil4mRBRYwEcARveiylAjMg4hfq
LPUYAeFV20UkqfKYT+M2RXqO+zUUAYKUJMQJ2a+aK8RQfQSlILhGo07P69o22Kn3
pzZhnBUFMoQ65OZ6lWjZP4OIPDnf2rO/GLHJ8+5SHz2u8SVxDQoINSMHJqFbL3r7
Zn/n6RFaCzY34eMyte2pnArUbsQNQ6JRSMWyout2lhJotDiIq3pGs2gv7I8bmS8+
DextGDmOvQkJeHvytbTh4ROfSorzFmCx8wDB2lqkTjxV7AtUHts24Y7CrGSZ59ue
ZgDu/JL/E+ZumXlw3Lfq1Rs5BBstzHtf2e4I7b73t+1NjAFo4Rq58l+HInF/6qrg
M1HyDjfrZT/d3CHb+ccLGJiZmqY5W6T7IrFwfnGdVQ/wljE9oREZIn4DKsDq+WZS
1sARr1sAw6sHQNBIejHb59Cwns6752GIoQmlCaMKof3noro0aa8Fns/3GwTkoJUd
/8t6MG65pUkg++iEjRmHsWjYiNy6u77eqP1VWopI0PmPSmPXui7kbymrBjqV3AQ/
L0Sq2rHh2uR3v0Hm0+gQFrxGVaP/Gzx+SqJuROhJZZ3JUvGZ94+3QH6bBqGRZy1o
sZ2PrXH+fVt6Ntl6slz+q74HfLEsAXk7JGsP0sGTiHxwkifhqJ+RjiGoCA/5shur
jbDlLoBXqMrms3+kgMvKT3ZLU8jk03LAE03D122TksmOS8JRDrx7GmGRVGAatVaO
JTh/i71OTbU2viBs3L7lM8XZK4p1l3AXBDfPsZDJiNyElEVqNOvbMka6mtVkpVl8
XD+MKQjfTgCCopplvhT+1rjPU9Pn5PnkUwNU8leRo6dy80FlO5OB7Vy+8dh6Coai
b0l7IDu68/eaxZbGFIvDcWyzAbmxEr7ML7XAMvYWA4w9eORFP5W9JtO9wkCa2kce
c7FwPLLTPcvgTN1gCziuRBKsF6r/IVbuGQeUcc4gew+pnJLPF7ZwthUtWlKuiA5Q
HbtBgUxZN9gaA4lkQ5Mn9HqgeO7U/vbUVQyZFq0VzNUeKWHRfbvw/c1n093Iwi/Y
BYxQrC7GVQr6IMaXaZEVbXKGycWNx8jsb1KpMQV9rt7cS0aNjHKdVDGvj1L+QOGT
bt7HYjUQXTmiGVoLkHgnOzXXkhfw1qsiqJtK0M5D3XeavjP2u4zd4RtZf62fZN//
9/Gxpf476JWf8CJxKrtwS0VDbqADToGfkJxxeoVi57yuiZTkPI9bnZtohnnXAEtk
+3XWn221PV+5WfGmzivWfUBVH+lC3XSUJUp9Q4EeO5oKXCp3etwaRo2VmjDbxp6S
GM8q1oxbkP6/y4rtbl5WBEGYMJO7wVRumT9RMhWzaI43DGeAMPQk+nm0bmP0l7po
xtm49XzOlML6fvOse0pWVYKW+NAx6fPyOrSmJmx2BS4pQDKivZdO0bRd6poWlCAh
fJfa6T4zTgqy858je5i96JQ4658eH+4thLOyyfA81NhUWsQs42OpgXmcUm1VDbt6
rxwWl9AXx+WIIeuE4wWjsUBmsjvK+kfC6xVdDyvbbXEeouO1o8sp9CckELpk0WCb
Q5hNq7RrrTclJj1FV4kiL0NFZIxXePNDXCsxH/8jwpnuorZfhUHPSlT1d8+nv6TT
05kce5ToJBJ2vNOQWNZR2XgjKx9EZwnTo4Nes0NaZQzPw8rFM3FYmu0KGAI8H13n
dcJF1N0NnZrJWVjuu/SeItv0RaiM1DBkFTfyzQucsc0fC9EjaSnrfiDKhtOiJPLO
F5myXbcOdgptLw89OWLclpndLYrHyoKu6QtYmwEHBJqDDz7z2T4uSTLFmfuL9XpN
mrymxigHk8yLdrGNKhkKYzWkDIKyAUDlOR01zJKhJSRHqWJlruGgBdAekGtCjr5H
Wb8eRppto4mdPkl4kbu4r/PEUFIrihpzkY5R5qc0RuuKrcbhpWuDR2OFrvRqKxbw
Wp5+OCUWVRwvdtwkDkqsLaqxyg+Km5c3BULkAmbBXFW161hWR/Nx7zSvRZRTmDJf
w7XxeFgFBUmJBHTlFNwYzIpBKfQi84tAxl2C6f5FIm09vy0F6I7wpEWhjnBfO01p
WLjMionGrARA796HPNU1yg/4yD80Jabw9bQegCfj9u7ApTLEWFhr3BqwntyRCE7y
qL8YqqNeTbNNMSSY/wzAyNxWqJ0ask1mNoyr9tV+4YfR2ZlwtB/WZ7nt/qNc33do
lV96rfrvyQSmhBjmkhXYPUq6TliGSDrqTTTrTmtNruOytwDqzPptqyVNjf0epxrN
7Cfo//jX3l6b4OCFreVMbJmWOwsxe2F7I5LoXrUfvlY2PwxUtLg64bzeeu4wqoZ5
Tl3LEAMWujdWuLSbhgSHMuHJ+OiEr7vN7be2Ihv4RNEjflP7OAEwbwztgWxn7NRB
FwGL0Yj2J4wzn5NouLGIRkOB7IIV9grqZskHUzgSIrKW8qlzE/0kCsyqGnYu9dCn
ApsJ+rrSoeognWmzPES2cRGXMYD9jDD1YV0iYx53ZKsH9cwCsphaKk3PqAJTBPEj
zsckl+pyNv/KaOm5hRzrfIx0fqQlfYZuOq9nAtQxq6CfGaWhuFDlW0TWGKyou6GQ
tccKsfEe6ymsdr/OaYnl5Psi5R18zmQ2utEqOzeDHo8kopiew3260tgIwAatlWNT
PjTD1Dp5BuY8JYSIYBRE4dKUsc4mSQooXIqJlTkJZqJpy8Otz6Y+Gthhae4P2Ztx
59APdsNU8amP4GHSjn1GQ8Oeh7ja340eKUzuZ+pAe5t+IehIKXt2ga3j0Ari+DyJ
GInQssYYPYHj+jHqm1fHGX8I1Wum/iGWMIoFIJ77tMuNl46Hf9lRNjNAg07fYqkM
MH9tX569PqhPZZtpSthWcyZWTBcUjCkrkmnKDIvo4K2QwMSEM9Z6scjl0aqMpl+E
crq3EG4vUaPNUtnnj50JPSlAJBm9gHUxzjQwXp1vrg5Fet7mViDLUuHC0UfAnvoi
jGFPC0f53EufMSevP4xjO3s5iS36B2mC/HEfmr1iIvIAekDO+M9PMNlAUcj5YQvF
0ad2OuAsRqRbUGcyC398AQ/bepFTdW4BP3LD1Ua7Xu6hxFnZECmYtJbxtT+o94gE
kfGBdEO3UJfXy7wyfLC3FKc7hrrHAfXuWkpNS8u7bmmaaBZUxMgYfBdT3ag0y6kS
PJ/G/l1PCOlTJc3BNiQrnIpuEElUicHuHS4aiRl1YSGYF2Yg1OK57//PsSlMUAvw
I3sdLw5fo9FNvdLiDcBm0LbFePT69pIbzsPqBqNm2xIry3HDDw8HbiQBkRip78HP
TmTAKPjVjU8E86/7o6S4oHcXnF3K3e9mQ5VSbNYjSBwvOMn88DX3H9i2UtOutPm2
+/l1Sz7/Y/zf3ZqCFrSRYgqHpYMS+t787WsgoopAvl/icn+I9hzX8iU2G2fsSeUY
pKth/m9mRkDuMxsRKQYopqdIZAcigNDaeJTqNJ1YwilWDy/ggrjeK55UCpIBND35
gPxD6RLmjEUku6L8m1+c4/+0d8tmJeourU6b6tevXiX4Jh6GS1Q8ZTsDfra/EdJG
MI5IOgt2xfNphY9v9BftIoScB51rTlqGjjo08FaeZrB3kEM2x4WBB7KQBxThiMBr
pmB0YCnPRPU0oIr6QEia+S5KnveWUS3siCYDpRAdtSMbNbaDDqeEvTvxmrG76SKc
I3ZMvVZnZVRr+gotlAdMw/4z1ZH2L05zX8G8BmPNgdCGH/CLljJkYc26OlkEdRtp
syvCfPKAEMpCDcmczS/uizFoHGpuY5ReVnWCBSOvITog217+JQ4VpuRYWskXDYIF
6fElB8kKaIZlZ26RpR5WyphbrWfb2dgJC6caGJ9W/CW0pPfe2RL+SiQGAPhVRZMW
bAZb/iTndRMzEfUIB5ZmgKF2dgGt9QsAeReyGYPJf7aQi/nt0Am8PmFIFg9JXpq3
MbqCaDPPRBqqfrCfPs/hI0KkcFkLHux1dEb1iu7DVGBVZivbWLWdR6VYHJq+luKB
VGqMpKIzKABruRhqVhiM9/XHERb1q2E5svWrn9MZsuWlB7NzQiwnDoZ1J1flXBuY
9wKKqOD3Lj+sbib1CB1u07MUPmvcv47qxKERR1VO4YxGhMTj6hhIUCSkEt+AKsSU
QdbgsM/Fo6ZvY+TUa6Wu/HGlQulPXo34LrrhfgiXjT1BQ/7vOKS08bpbdrC4ZWli
NM49gLOuLL4TqUpMlDMBrzLCA+HcjjKywyP+AEreXLpiLH5ssVaKcBVnI2oqS++g
C+IAXNd6E3xtocY8yPq21EIm3/ycBBMsEKl5QPgk9vwtXsHaPV4WE+2eI/MqatHH
zgV61cGqdnvnfkucZpyD1Nk9oxao36UtkJFvJTqqZMJT48Mz6dyDUKscTOuuz6cJ
ajCvO9s/z03S3GagcjSsi62n00G1YKmRuZB7TimLlkDn1K4RDRKkEzU8CNKZbfDB
Zgxrc4C7v15+X97+9oOZi8kcS4HlFgZFKbtKzN1apRDf7WT7S00IoKb2yNyIO9fe
XJ4cILkBUtEerwr59olji5VkDE3ivTkrSr//O5CkMODL0QPwFjkIPZJtwaW15SiU
ONYbyyhZfOMwXliQAM++HI59E07sPKrV4UXsPFB23Jhz8g//rxXhtBxH2mI/huOq
kBCExo6EI9PJ9jQzIOhbwwUw7uX+9uEXopy5hSeHzvx6Y0uQXS8IZhb2TCv5GkAJ
6EskeySIxvGXMx9jXaBW+RF29aeCtL3C57SFKk/nEW+qAlL9xYSUSlZDvryDtLY0
mjM9mga05+OrNbYfqfLK2A8fxpHUzNq9sukU3T+Frdr8R42f9TcqDw0g50up8egX
IR+UHGaHVrlbdAukNWUCU8tyj2wfpCk+H+cKtuCAJFuQJDQUQoRUHRQJUj/42IWx
O0ST8ebx93H5pm4EXAYJ7aJqFsMn++lWUjmePKY0EFIRqxhBIVi0zFprB/O143IJ
snpWTOScBSH8AbS35QdMO6NQYwnbDjeCxvgSl69/UI9P4SbJ9edoM1gOQvBxfcUv
CqXW2LjZmbS+fBIzuJDncx+ZAPmrdFKr5LmJgQqk+yySFFJnY/gRtpOQOIYkH0JS
eguxlw101xEQ3Xwzmbm2zwcgHPyqD5jjOgP8kW202DRH5cb5Kl3TmRbYszbF4W6h
JW5fZIdxk2IYimkSX1P22chFBPmOuC6HSOZbsi4G7Qg4lJ/cdh4nxdUHMbKlFpae
9bRMRSmxdBp+hPNKJ4QyFZ7P+C+iZUhkqQWSdxUmV1FWbIcpzPbMYAd8DNu9ReKT
rHi6N7BXOJInJwku1L6pW3jTJvPGGUbePQvakLUxww/heBIC4uCJoDZ9n0s/TsaU
8ll1Fj/DFhM2BVXIfS3Ol4TopFW5+RizKdo4dhDR+elmVl6S259AiUAX4uoz+byo
L+fTQ6Ec5kTsg8dK7W2NJKfOVauQbCSHguAC638/05+GLdVv2ZFMmsFL9pp9nYse
EQEJWTadHemiL/3lBFaWryLgrjWvwe8b1HYXHINz/zKnKRXusu7P3WMSm9XvR6V9
oJHW+y5lIIS8A8irTbd+l80Q5RRjPC954liVwrahoy30tmY6SEYYuQGRFdXbjID6
eb1XuPFKG/iRJzNfzuTKQuBeufeb6jcFmy8fJVdNkap3I+QU+8nKpuBaFKKAVxE4
4MEBwReyXyYS/auvqYUvBgbBySfFceKhydFG+ndL4yXNh0p/iA32ibIN+ln9YT0t
YLOsg/v7pN8CxTBIbGkG7lI6y7IVw+vQ2t4+Slxw9iS+264CORm0oMHjpsVBLQzp
bMZJSxlWcuoAk+x2kSaw9eX1BIQAKWddMZZfAd5x9lNtBpWjIIbCSatQMt4LzBTV
hQTIOVu29AtXy5/yrzTNqn6fas8YRLKJU4+W+S6CZOqBxjIq9Nvo2pmcpp+SEolN
dCORHjbFwkDIcn36zmM8ixAgHvdEB0budVavXjhaJzg5pGBK8A4elLri7jaCsMNy
Cj742zmPIGn4JEAy5FAhB2eJOE/8a5Lb5u3yLRs+BIj+vtO6OdD8lOlu9bU0KcUO
XKGaPDrHQ1WvX4aTJ/YTg+F3lqtJX6jWA2i0ocqSyPOGD5ld3woF6Tmf9KLwyALh
eSt8cSJL85jp01aB0vFCRCoeKTu4M2ppcZ+FSihYCklSBDCeGCmXTEQW5MEZfUpY
YDlaSQYvf6kGYZAnXtjJ4TA+01+pP4WZLnTqerxqVCSH1alqdi66eW3d87y+27rZ
AvOdu10MwaZY7+LnjaN2rOiMB0Yblpx2qX3x+IDEEjwnuS4fv3xQ2UvBPzJbeswQ
LgFnVg/JOwBE/zzdWgXkobfPysm/ZVCjHUHNTrhmh5/wnvbIkB6RjMbgRbnDnnc/
qi5xYShckB4tzQbSiKfVRiSi+K85dbKyanmOUmROOarfGFW1vo7qmM7AJou1OHFa
6ttUE85mEfSaG5TZORvRBC9tiQ1mtHXauymDGF6mSE9IMTXGQH/yA+XaLbW1Bkxb
hUQEFaTiroOn3d0wX5PAsuD7kkzD2Fh4hgogOf+mTb5svv52wfLTzX4YTn1mQQXw
1WqB9aI98VopId7+CgYCpKMwn13TnCbBt20T8C+Y296vZDBcFLSFdXLEnyTaG60G
+g4TheqFTcB4yRRA1/nanmHxlhHJS5LO31vAmwqVfMWVE/Deb169o0glma8CqvXP
8X7dmx6/aDAYdGk9hba09Nb3HpbvC39v61ECLwkuVWtDSz1wE7KHOh+KQxbFInMM
9r4u/DKEEtKTDSNXyK8McGAH5vrJGhHI/YcL3gLhw1j2tcat1GMRAxTnEz0ym6a7
2Q5Js+vo4KzndqI8PUyWg9q7cDtxEs6u6jMv5DKl485m04PpQ0C2+OEl0TQ8/3iv
t0/oyUmp6x3l3I4P2ok1UiRZ0WsrxRlrCSxMQCxPyO/fjOThkmHf50QdEP/dLEA9
qJf3+0pUHMYcMEp0o32Zah+PmPEO7CYInVh8OjbjVLcnUhGThaeaaxIMTpgF1Sdi
l5PAibJdBjikOd5mUlRMF4IbGNBqTaN/7tImGrxYbWjiBU9mM/mP+4Y1gM9OPzU5
Se2YNFWDVuGsskh5ZmkiKJ81/lPhf6ptxYQJLEo258dG02timaRrMLW23olJtHG9
INQUVZ14yk2p1BlCCDFUMeHKp+DKI+8WhYa4vgkKhaBq8FVGDp/K2SMaDlkGEwDr
RXVy6PILW6EewRahp7SDhFuTNS+qCuy3DaLpG+N0CAWfZwTvb6M7S72SEgoHzv1i
4pE3o1qmtA+FcAQiH2afFw/K9jyPBvsZjDVANjVvW3LjFGqwHawe+pMs8cCDugTr
YDT8p4ukaa5OH4n69BPTYUiVAynpwEYR++BIj/mz9bFF+Mlbf4LMASMC61/hLk6A
ZU1/dPKg+roYCdfOyXttp5Xs4AHfEAgOdKUvEqRx+4rC3yx9joDDYk1s90k/Mi4i
8kpx3F8ahC0BlKY3sLF7FNb1dWXDNRoMvj7Ou6H8UynQzmgqDasfrMk5mzHnCzue
rlDmFOajOmBrgszrz7elV2saUskp4X/3WME6E84eBWWXmD3WrmLdX9poi02OyiK4
/PrYoWygZvJbiyi7WNTbcm9Ey81KimRhEOotWQydoTtPvlkhWyzSieD+0o35f9dY
R0fKl5V5D8zRVQK448SpO2hcgPmYEJo6wW/BxQ/gkhA+25SBsGHbzAU3PkUD+0kb
EAehrp0chU111SViad8NnodddafTgegP+fnd7k/rW2XwXFFfZRWd1DU+00Jlj/X8
fSemkjx51IiGg0rhNGX0jD80Pc+fzm2IbNVwehmyO7FefKu/+RQkLQ3K41EFyb2y
TDxnTk0hVwxo2RpU3qiTj4o5J8UvfukVh/OdccbjXxGnvr9gRQ5J7w22lZ6tCzVt
pyz6ZJBeKsjYVDa/5rF1Onih8MZezrFB9uuTTIg5keUaGmHXNn7ColKjo7YPFGr1
TDOeaFhatva4DGn7OYEcEEoLe6ek4J/D5t22vBBXCdRgbWdgDNnDwtWvr+1C3hPJ
GnqLK0zSsr4IJLNrmqA6XSC8PPe/karijpzYIx08KJftcpkeD9/3OsXT3ux345G1
pOGM3uPl6m+ALnLVNNubH9zhTOWU58Mj3feSQaraJAtg+SJURoTpVQg0HWca781u
uTRU9ewrYtkltY1fTfTpWAzs7+nQwk67oM53S2Agyn53YcnBh6dtB4XfYuj5EuyH
ce9591odhLLkZ+o25ZsMUB37ldbvUEhYJjvpbgc36E5jVkTenvUqh7z7y0u2Ouz6
9ok6qL2Ol2iZug7KIVNr2U1fs+bBO7dr6nRc9jpp+K7ra2A90kdi38UpVXP/e2Ka
7M26s7MIr04y2nw8NaqOLaXFMc8wz4sI6VsHBxCYVHrnM0XujVtEyYNBMcyNmQAm
m9P/2KvxuVK46PREDVJw5afxSl71jOl9ZodMnS3J0xY5hbB5zTYwUwDm+UaGdPTk
2MsUqvmOog77Fjwrwe9xHPmcANq4OFc3aaHHszVlAEWN9462Xu263gxjmCv6gp4f
nOf3TkdsmIf4TDo7U511wPu1hhU1sHL91Dy4hJTi6QTzi4CPfq5HeqofkfIMFmR7
6tQVb27GPFOIDfdKqWhtd2E7bjA97aQy+e4J7pX9gG//PzTU5Nlzhw7q5kgT+b4b
UxF+C709thSzIHp3C757EI5iOFA/Fo0R6M91Gs+lVVVUixvo+CfnoGWfNVBL5iSj
P4FYKgBjLa0Eq7bIs16hNWwD7GCc+eTAbzy80+rsyusR5q5cXG3u08GfW9Kc0yjd
aBRImqwjS+U9A8jDRUMciYy76dZVF1W8/UGSE8RfhCn7RTGb6bOvH7nYgAKw+79k
SG7dV0SiD9nu7l/berTsfOMtNjWAfetvq9COnIKlVYH1ufxEd8bIOmlrguY4jZLW
qd7J/cTz+YhkjGiQmyqiskcvh7sHgpglU+7CD3rl2lmNflz2g76gCwLIA5XUJXyP
68U+yKgDG8Xj1KndIzRGnxH2X2RPvq0+TdVpko5v23Fl/jqRB97E58DAmYchBtef
N7phIEDhry0zBREXfhaoj+ZO1POkmaxGu6MbuEEicdlZ0R2SZxli9nJ+P0XGxufZ
LCdQojBEQFYAmoJhWKgXrDKGVQVkSssDZqcYuibzf71hF0Rv1D/xbcZrfbuVVp17
NUmLQrmJnLgpMgy7VknuqWRWhFvUth5yp80Wy82oPSEf42SUslwhA4Y4AyrLH0ZO
TO1FeegjOjv/wybx9wH6VplBtEXbwpHB5LK3iBWm4wCY9YSG7ZdLK32n38E4DCF9
y0VsqWcayWDTahgT2GEHDo0vzqhIyz8OuA0wPmVZo9mcDpiNxVgxOCh3CZ4glVyG
CBhFk2ee3u6pb4q7WQfTRsj9veHN3M/jr40njkhGKMQtpOkoy5UrglNb3pn1NKpk
fWZzklhzR9BqL9lB3S2YI0w3ucndWoMNRBoacW0+FeieOOo6ZzBcQoEimZFeYc31
TFmtK7GH0I3z5EyjRbFi3AiLQJnq4eptVbj8UWv4xqffFF+7eF20Bi+E6zTDV6Cx
6OUSFhH8Rg2TXUBAMMP+u1DdCf2LCaNndWs0iO0k0zVWQ2jRv+M6eDzDA7lE8U02
5FSFOSe6ICfWlMKMGuytkxtajWQ3WKkjM27lrgY2NZN1qQReer6hVlCVhtdKrJfB
RIzWr8zAuj0/zA+L6eA68z6he1MY6DwK2NiQwjtwKonxxR7tMG9fz1xg2nl20e0x
f1T9gsO8CRIyMtYoam1Q6mQRBcf0sEJMhu//lS+YUrpsz3m1kDy34fn+dhWpKZ01
zFwrEB7hJG0UCGuThEMzXAhTSTTSirQewj5HihDE4ZlW7got9YCOFk97AtgYsKcs
fNcilPWJ5kTyKSQVoD+WD5JMb1DhdouJS/ubP0ETclE0SUJ7KCBZ4Fw8oB6UvFvn
cPTiDICOp4TS5bnxwy0QfGQ3m+BX2evVVSEucJhbGyjMMgQw/N1T70QTaFLI1AIi
MZg4Wq+Th92YM5Ai0WsvvhkKIi1euKakizWNrxIoYqomMb6Croq0g+SXIf+IuE7S
j8tWfyxlJd9aZ7ZIQ6BO8DbQMovQP5w+7Sp2IEWUGMF7Ol5zlTqM3cVAlAlpXD8Q
mcWJpHFKkJ5m41blM218kTvVLmazxhBk1Qi9SBGn9LHXqm7iS2nZk8I9l5SLRqKq
D3amsZPDX3qPc1nm0HG5D/X5Q9meAX0gFugx77z8/4pSIYiS987LzpaBXHLuRlxn
G0AkQGydmY2Y0UcxB/9HPPskDOG5ekpjIY2q1LNkjFGg+5w4lwIo07q0kAICDeUy
wfY9XPdVbgGK7nh+93I8leZquJWkNpU/KK82HINIj7TppsyVwKfFO4gpJqUwlaPK
tPVnY8P5awRUqyry4ezOBibXdHqoY9/2H7pFfGs8zk5EJUn0q04cPwUIZrvdS0OO
yqNvDsJMXDd4il2pu11E3MEXOVQYBQ+GaF+YYk5Eega+8+AqfPOneDUG6OtyBGRA
fVS18pFW82+YdQHLc3hzcPdpb9pj6RKj2d9GMGoUvf7ljjfWszJgJmhsHna7PeGE
d43SIQVw9r9qFluyjwcNpR43qUg4PeRxqIPKBktG4p6SUXKMvwNVSn66xrOwr+3+
v9D4l+fGHur1ngaMx4+KlUVoVgsGupwomAwKsXkYhF/EkqVlVi0z8AxztY7VycoV
XYLXTJSF23Q5bet+5SddiBUVQ+ydm6GMCxqOonPC6hGUBUultc71R3eDz6uYAafJ
TLlQ4WWKpLJ7wwbGD/l3lfMofEQmYl/LvgVlq7OHZIaRiV4ieP/HRdWdiBrvuLbo
hE/BCl+HbrM/gZeBZjB2bYC2n2jDD0SRbmTx/LvRsj8XBzJkBxKza51JiMlvYKjw
iDb5akch6X9l6eJth20gktNm2C4H2HDlGnEa+zsZWySXQ2P+Iu5IB0HafIDfdrby
ECcv5eP4Q3Pet2pzJVxX51d+PaJ8+sp3r11EMt3W60MycDtnSJHsAzLaHD9rPwzm
5LZauizTmoyXnEdtShoABb/PcKCu1Ep/Iqqk+FAZchKvEOkv+nJ65TGZdObRliac
smFqIcrbp4kLizyKcSKDRagCGYOiFCOfeXHy4EmaSOn6zG65oD/QoQomFGS8iJSq
uAnXRMba6E2xQHWgBlsP3g92g0pX2wlsnJGmi0a21DH3q4tvYpRltbcDN+I15Sr5
c9HkJdFMSSmG2EarswfvTz11QPVjBnqYkNNX7qT0vwNy/A9Kh8dbkGZt3Nt/I4wl
WWexh25OtUo7tcmvp6XeSQkZ3TiqapeIrKbJDd8PJxAifEbfq2IwunO/TCMhWdlS
1msJ/XEijr2vbMxEQx1nzRHkIBRGytwRV5TrgZF7p0D90+hQLVrgfaJll/ujwjfW
jPv3yUh8VZggK0UZf0pg3J0V+lMCkDI3mxXdJo3T+WTUb4AgOkWaFZAwaTUlRFi3
YCvK5q/75Cy9ayOQXH+osW6ADQR81TZmbt5rGxmgK7lOBFUat8+VKsuKUtnKuc+v
XPphYrB9LsQgAf6kbwAHvzzxUDGmlyQP0fnCwt6DTP928SRBF+nlASWGo1N8ewKR
rwGhN/94ODLvW/KjGFGOk0TWK6sceCLZWpoXOzMq+TMIKzRGi6vvNZl+UIE3mDpR
be3H3+wOOvW3n/rjhD+tldrdsV2xduXybpTOi0gUKSff6pick4WTxYE6gQQysguT
PTUZpof5ObdfYgHHN3jfdAVulkzsKiaThhpIXMusuk4Vax6WJBJpoafw2LznIdcP
uQv1Io7fvdMsczbnLpTOpum+L/LXjGK3Has21IATgRV/a5C/+Wa4Rv+DoAXOfKLW
gKrcpWAdEjeLpo0yWJxbiT6l+MkyRTMkOj6q1mZCBzQ31o9R5JjzRuhIal7wIAHj
JzugvBHqwyKFdxMsyuadphAX8YUzVMK1nzKesVv1ZkeYQocnwdZ/jIsf2s0fAFnV
iUdeeOaIOu7tfZRFqBUj/hloFAjMBHMl6932rofB2k20PuveDWOQUu8kA9UF/nnv
F85JROyU9vFQ3xonjMX7flj+z6A+0TxaCYdHR81gehenAVPmgLRR961+YgY9icsN
sfGsCVfLajW5zT+6wQ/x1DyzLkw2GbBQx1WVrp9oRvB2LKCJcdeK1yE6ElbyK9KX
zyX4t8sh1Pey+/GjFXWlO3oOL97o7ONmiFtbG2EMuFlepa8BEsW981g7sY6/5SLm
+xPXztKnn5H3WJOohIaJ9D2y/0pZtSRuYARC1zkCHvmS8VSmFyGhZXo1WRcdNPJB
+T9teO8vxssWR0DdCrnSTFJEY+d5mo0QOaSIQgO+hJxd+LXQZNW7NwhllaJ+2ws7
QNrvU+Tk9c+ch60+9r8rNwaHPkeBmf6j3cewsKbEqGwk5MlcH/LM6ECOIIGoFx/M
OrSycjt/evZPx24XZviBWmdhVUORW5iTnTc9avzEHlzHK+HcB1r+STWK9PVMsx1o
0jq/dU9cJkey/4gj7zGU6TqhISAm7MgNTRjUZmp0jkEYks35ezjcmxcRXLxbNWVw
pkSqZX+rXte+JO65i5FqVW1yiJ5CCjLNn6KV6pRkVPJhO0xSxM168GymO81bTGTg
Z/pBXRTYiXfRrmqNSJC/+TKrrq1JHlCwnCLpoUyuJjNwvPxlTX2DHsUBC7qw336l
7Xn8HxXQzfcJ4Jyh5Ny9t3mT8ir7mxM24moZAZyF8oqBtYYstgy9xx7ERcEmDBIj
UF2vIP6RINgQ4gCbp5ZCneY4ZKXnTkaBSjUYaq1wAW0lQGDxvv7BTjznSJm0zE/S
ABLhGPw3Gf1JQUp3PDsdw8lEpIgHaNdyA7YiVymg+YdNY9FpRiomSRl+G8n/en9v
X624nobdgzQ0x4U4V9CEUb17Ae7cYEZskV0ke+E5qw4THN+rKh2q1zdMLuFqVUaU
iIae7taIqq2rJFIu/DtidVspgIv151XlYkTIcIMhi0CgNDyRYMMhmq4tHCiOuHZS
wJsam2lT5PjKyhzcJezVdQxrE0FehS8By9hdZMZymbRwRls4k/tlL1TonzUPNGoP
7uItR5Jsklkoh4PHOW5edTmvQm3kWJa7ygm8UNI0KKpt7JmIeReA72ye6TatAPFf
sF9EPwnYSfNSfkEMUR09WXq+CnDrqDFyk200D1csZyXZoM/gm7z34iP7+zvLNwEW
NVmDQGjAeBEkCzTDgvaD+lo/A+ydoMFL6f1lpVZ1DfSOSeRx0qWpp96/T74hPi8e
PnZFPG/HRq9yzAIG0iLGJ9cftkpK4QbbDaLw1/AVfdOpFs/ckeIhu77kImrJcMmV
TLJvKuCkUgjIZOLxdqMCBIQ7R3zF3olUZ3TRavkPe0pIY4KXhGOdUg4u44U8j6g9
xVietYq84oosXqRJK3oIZyMXOku9o9h0ZiDaN2uDy3JAEsCzrh1KntDk4PWfKItb
9uO5uO288c6iB655elTnmVl9LcsGl7KKBM+7wEbKwwTAhEBJyEfOZV5IB3VwG5xp
D8RyycgnHMfPuSJZ5GmJqztIJs7NBBvvltwaOAunzgfGJv0wrGuwXZCagMiDza+8
H/wHBqLUqCuWBGrnt8Xt5poT/CXO/RGOnc9m4HG0rW1mAQmF4ZKoUCgsAOhdTEaT
ByXMu8xKs9cSp/KVpXUTQ1ticrCTc0iF+XfwNn6V9TfzK0P5eRPQEkoEEw4njRg0
Cv07Nerb6ZY/UfspxVYgyb70wOWClSh5yC1Kb+aQMenkoCmxRxWNOf5Q0LmysmgO
IMk62gUQ6U5ojUyfWjV1E0zCDy1zslSSoHR5fTTl32NODINkUB2fjRFHsRytuKv9
g8vnNbYwf/iW44kYmKG5MTjp8zH9L0wtDcukFJNL8j6gnksFXfmTfRYIOZZjraL1
ZhVyuAZbg8RgtgcQ9IT8TcNmYnQsOVmnn9iwCzG0Z1g+0A4CmIdQKh+ZBJ5KVAy+
Hn1AQ6FxavZ50gbbmd6aZUwBmM2xxRiQnxZKLA7Ing8mHWxm64RV3dXbzBbDo5M4
NVUg8v6BGLE8ewAiBhusGILUYYNc1jgK9tKHdWQd5J1X8Ff4XGHbwPYp3jZZBpOu
/EZSdJ7/OarAzGJdtbY5ugoqhjlDAFew1iqoT69in3wjhzeJdekdr6BuZaibNIRl
rdZeSBHB8oy9znoxIfLtw5jxGlM3zS9DYUUAC8uDiAmEe0Gomq/eTNUwK9OPq8Jp
kgvW+BPJEHEwRvizjRSvuCe1hGB2xDDRnC84OPB4PpU9OZIxnZtCUmeaFiTtw/de
jHnn12QaWQHMZzde7O5Esu2SHgifyag94E4T+0q5C9lY4Rghbn66npZ9LwdRKJSr
cBK5yAu8xJngmxjAmwG8XXRiJRu51K/8c0zE3xKMhUfYfOSZMlnjYhZfdQ7n7Vfa
txOqWJRoOugwjaexhYB0oiNKbj0882NwC59N6Uoic4cuza/csHlqUCMiR3vXVIUz
xmY7uVn9qsIOfiKojN1stZ5yWLsB94RKVG3WWaVgK8x4Q6GSrCCjpmqagiTcLbc9
lom5wO9G12uzodjBdAzDBEyaVzPl4LN3zstqinKIRpX7YaiTNOyNTlufTkKXPIgh
RAx0IS9aPp8PIlpmbW3NEhwXA97Mi3gXZhF/fHpdJX8eZPX1hJBY/Lw5QuOl0LSo
lL3KZdQUfdJDYDK3DYi0FqvDcWd7teX783kiGXZlgOBoHJ91u8mqUzFZRid2xSCg
Xsn8MwoRcx2n9Yo0SNJlJ/wliFk1o3Zo4PteAGu4n+HooQHEo2O2Kdldr32yKg6C
cYy1In+mOxRC0o40CxucdpQ8y+j56yhS6PcyUQFPocC6u8+L9aNJghbdziqWEk40
BhlXtOTVMOoJZSjdUViNwHammwkBAwXLbkUuCthtt5+6vZms/U/2P/ezX2zSGo4s
OeWBxXbvcgJeov65ugWwx9CaeHg4BymD1BGGAZ8MEaw0LjFJRGdpwCV9eCWFX9Pj
N1uIwEJCioDqBptpESnuU99H1sNl1x3KpMxqHLnFS3ZGBZkNEzQfh/KTC6XoBUt+
YZTuhnxZ2e4R4uCtMUbdXMWBEMKMkQLGa8Qqn5lQ6VlYndHI4dtoc9Za5Db2FlGB
+haVEJpEljjfNRGgSR9pR+uW9qnJBXOYhy4/fMmrrMyZ3MzjBdtAqSCxPsaoC/Ms
7285qlxeN19V2HyugLG/I4tbqQJJGd1wqYIwuq2IBHHubQ6wDd2NXhh/vzfWmPqd
Nxll92XJvahrRqe4QbHs61944OzHEg9xlnhRMoj9r9vAipziL1w37TwRoY7hH3WV
etFrUPjYil06owUbF8BiKXkN5e0JoQDxcMyIdyGXFwc+W5Qzi+bugYtAQLApo6qZ
Paw688RQcISySTGGCH3c07Ese/uyRXEpLGdVSz/ZYOvChJkaEJMz3AVXIdQlcjx7
7REBedUzNPjDqR2ltUcJ8S3LSYBVEDaQwhBbA3EdeRurvIwFW/ADtKl7kBMp475r
H5SyhHuT1DURRE+NzIwH+RugIFpCwyDXMHfvAiqkwrMPePhV2ojcL4GMY/7/GW7X
iTSuDgY6UUH5Ge4zh7f7E+DHVErWAog33QmMlJUERCDXfv6/KRhjCZX0Ma7PLLIM
Z/m4RlYzSuzfsCkYvDTrlTTzsBvBTVlblHrFfoYirQgsCFOgfrUgnS5oSVcctR2u
6IfX0JKR0Zg/BtTIiE34c3ztcUQH5PMvP/uP6lomvbfPMjkS8sQ3DkVX5k8m5VeX
iOeMkYR6r+6Or54RUuCEf8NMCqaTMTLFRGRulntqeUwjXNoe4HYsOnO13XG+4N2d
ikPJlcKA/G5sE0KVa6eOo34zeO0jru0Tl8Sz0Zovg4O19DuJcohHzJXXjEO7WVx7
k5SsKATf/hlqRrsi2PeRbeGSYhGhIah4FnVYo6glhYjQ6mgJr0/YwmlZ3tdJxSxt
UOWWiFE4o+vbcj44Zxz8dnWATuduXeBrv0GU2tOIGCmKQezpCwYdvs+nlZvaSbz7
PiFH3pTXtGphHDS9oVjaSlYdzFUImT7VomYEx4jzF1WZKv7sALhfHvB0wphS34CM
MZ3NVIENxQ0BqqTQSVV8P12Q+UimhMzlELOWKeoJ4QeKHYzBrV6CG0SR9bCkpKKN
RiRiwplgxw5/08/TLsHkQUjyIizETJOQ/AtXlST0kIZM1leEWFsgdFxPeBlkfHfN
2HKp0GEvZ0D9ovCaLo/U2/6Y0qaHnyltMC2BtYem4jVDrt1iJZoxKervYCwDQRw0
rYBxmFI4hYNHOiah6PTnFla2YCf3GTQeTDtmP+eUNjL0DSHKqfFKLWeAnQDaw8Qu
tNkHJDFqEea75FyE0CTaCmGSo63p8ahzfYto0o4GpncxIu4Maqxr/2/bgezuVbFL
k/FY0/feZttS/QmgkrEcC/ocZCoE2PRFrLkGTqfI9GW5o8bFr4ylAL3F3XQW5dEr
Z9NYTfB+2ECa2wcf+ix4BZu0FBf9lMN54BbVIUR1Esw0BbbEpLCXSPvChiUdkbOS
f5x3oqIm0J7QdA8piYur4VoK0RMyMHhd74bWHsXYXOItMbGcwKZbIG9Dhwg1Drt4
htWJEINv3cUPz5wauxeEd1/BzNPbXZHDzz+QdEYGn9HmltTuZIeOMmrW0lz0/QC2
84Z1V2qxpHC3uYWwoez3S7EgtqLee8dlWByFgZ0GCs1DxJg5/CrO31QDtwiscxD6
cgy6eLnhCXChdx7oj52yP92RWyQz1rZsrFnFxW9OVQ0KX5XjJW3hNEaYO+tVbTfG
P9h2+B3kLY/Uwu0ROqTY63vwHHhMpMe98jiD49kS4Vg/Tl1r6Wbsx1lAFxqhjUZW
niU9CBx41fqUPnc1vtQr8onLbhLToHtl+S/Rlvbozr6lLgLoZ08S//6h8qhco5Dw
vyXehI3ZNt4B0CHlYQY9d59TLwQzGLuUTEhXH3vYnz2lr1RRBb9s6aKchtnAixF7
GsHeykdiVJHvYqb6/ptXXz2i3fHfKrscyw2jB01j+0YbQUwM+Bya4o/lv5F9L8Xn
5QuYaEiPMIZVwOOJTfl6+QXVmEXY1YiRGrO3sCwunAvHidL4ooWydaeXNC4u6cvm
G/lxelCSHI3lBM+g7thGGI/NtT94GR1O6Hj64MWMYtLDyFygS1vObqlFIkfclnFK
o/C+K0TxpREmLEHfFn/skR+LIh4JeCRyxoPnXhiI7L/F17PPuRnG5LgcGKEDozyM
9dRCwySArbM5JlIX2wAC4eNc1EVoNV2UKF1n0OcKVvcR1hn0/QAzfwC8hkDo+thr
qG7OUONgvbeFuP3QaOVlOZ12UdKTOBe3OQxgwU9TeWOp0cbM1KSnHxAjmy7oip1u
hYLtE3RK9xnAEmqSWqGXIBr7D+uwf3YVf1BWo3llL4YN8blP8nT7MWHvVIed93sH
K92B0GY6BaVVO3VIEK6PnOKnK55JOBk4FsNKaULEdYwKwWoaVOeFkZKphXoAXuT7
VkvIxkjDMTRdzLY32MgHgS5LSS1S7T7S33tqnTMwwhAFrSJVRF50GtdThIqncHMU
KIX/vbEJy5OIw9qdjpXlIpI/GdTQ6VNr71XKUZXZk7QvMut3hR+sN7wPkCyCV6fs
czC6uMTSAA44RTIZhOdmSsDuxi7lwIDdUnjcFXz49Lh3B6rH1Qf9p+ayncDxwBjv
ZC2Wvkim2dXGY6X/CpluYU/wdE2Mijlb6r564s6df5Y0NxEELADcKNR5naYoaMsv
ROXn3AMmjuGFSPNHv9ltM3WTEsJDQN+jK1SO77Kh2f3SXRnDO/BfYjOgtPf3HmHM
wfiT3DdTtPsxP/n3ieExmT9LbLBU1TofWEK1h9WkXi3mhzBSv28cvv+z87p6v1gR
g4rHpKz5ON4CVI8W3YB/zeKQ0BjNcektEtHMGSdBYmTbFuirn01U/gE2emJq+89S
UAxJtbkT/KwOKDXF5F+0PFnFqxO60jgPdl7SYl75C0HT0E40y8ohf1BvnEZihklR
8Ha1ICuNdKdReq8zr9gn+X253LOHmcdjrY0h8B64227cVjd8kmZfeg0M/oFE+LGS
f/YXU5793UoioRJPXcwSbBoBs9VlXLH2hGBlnbRZujZP4ar/XaSdFPkpmEsTMSsQ
RikuUnFT/t+V7PxnVMexDdfBWZX7oy+hkgAvCygdMdIFF364FbYLPExOcNf0TreI
4antX+/gvVU2phZ77UFmxoyJAJQ3EjkPFQSNv3jWfPkz2IIDmSiORx3suiZUfgNs
Y/P+w73X21dvdGdCwuqh6extssbSwdMZTTc4JOvtLLL8csjE6FxOVpyBK/hdvQRf
wdqgCrcXGFpAGvbnHmBUwUwgfwMSYzNLEAJSW6nI6fjEgl1eZpfQbC+EEVy8CEqb
OMDUbLmmIMKH2PkxR0Yifw==
`pragma protect end_protected
