// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
bfXVEI/nX8Mo3oA1NYQQ5AJ5beAkfaq04/GZqyX5nhmz3Z/SOgCxiLM2/GopTVTAH6lb4eTT5cAH
yDosdv80IMTe8OZDtPVyAWCJhU2H+6RZYfr6PU/kSrkehgz9L0YtMiNEKObz463blwJhcfwG14t2
+gJQlRj90PZ4/5j6NfkuXPQBCKWedY3lBEG3m8cM5Msw4UXKboANGDDSqwWM2cXth5LA8Het8aK7
/S39AryR9bXzzNchChtKMamKDl50ebi9MWrQudXGVz79SYq5rMcckd3PlEb3+8qSxwTboNEGHwZb
ATbReEIA5ejSN1i659EXzav514CqNanqOy4kKA==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
dnhrVfhr6V/ZyAP9x4TCGOJtzaNpZ6kk7jPZHQi8jUzoAFZtjRWSSbK9fOohmYitHwGJVV6ksKBX
aAAgUxdy3Yp5v1y/yRZCBG3cBGb08agPqWc0zvlfoU+Nj8BFMQshOuYXyW5Hs++qtoIcvsO7OvpS
rin5gcIbVV36sVtyUn3STp3czjPmXPYuj2gLgLqPWZFZcv9P3IuIwzFiOrj+4VI4pk2yuW2lnghz
n5QmNHEFEXiy0x2N7ucTKZsUfXZ19RvQzTobT+UEXjoDq+Ar0DgN+Oy8IYGZZIzgB6VDqE2WqFsN
FALmJQsZRR4gRhAUV98LxpAIhMaI/tv1Q2wsgNwaevGUkbGeZo9I62ZXSA47tHhZFb1nTVi+PT/4
yDiNY6wUouyhpWp0pSnXnA6sWGH6voM0IzgcTNmsaJPOZAQNIdz0mi3IJM6DYexdztHdPlI6Hgzf
XDqSjRTA2+OW0j4sC0k/IX8yKa8BDjRi8pfxKENf+Dp2dbwHKIjbqghBk0vbZKF4miQlCn5+VAch
GelItea645TFkC2+/tvH2Zok5RVx4ydUsfUljxUpEIvXSuU8PskchDmKTtf9dN1Jxx+VNTEaIA59
tFCQPE3XFgMRnBTPmWWOv6wev4pGspxY+X5mbc0ri96n5PxSeBFCBI4YJn8uKEmfSRXrHOZ9PkTs
bA/Mcio/xLmn1gRuSbyzwXiRUnlbO97zisZ+iJYT7D8po02GK+AW5w+GO0b6S5ifFiw62cAUODGL
x/waffdDrBZnm8Jrmg1EpxVhslwx4zvHOEHvmOnNNsJZbD8GLRH3AWVUBG6INAqpcAVtQU5KCAg9
J2vVqQPnWVraVva/mSArPA7E/vaCK+G8oSt3InPbkHIkGjp0ODJHBpZp4xNgEEd+CMx09EIfJtf6
kaJPjFyX+1aJ7wdq8MxX9HXmV3GKcLhT1gMcCNzKUTlcoV3r6Q4nu89zlCKJsTpxEBSMSqwk1fFX
Rs9t9sm2beMrqujgIRJvDo/o9GgxYRbUECPRdSl56rD0Fott1C/Wk9mhbruDCJTMkTdV180rf/zc
Nv4EpyPKlIqvTl431bQNuGiCsp7i/bq6bAnGeVz3Hp7vm6fdj8XiwRznx6X3UDuxz19uIh0xsJd1
P3Z6p07HdgUEtR/IKTcoMJGKJY2Jx2SHuNldpcnbZW9PUa93AwACnhEI8ewpjWuR2dm0eML3VOds
hK8kYG5pg8++MbpzRs7D4jFssGV5Qym+m1iWgNKxgGlTNKFDPqDwYS+gg+pSIR2LFNBmK51AstN0
4MmNlwIEgNj2fvagoKl/ul/dso8dhHRqhr2qBahz97wUZrDbtTdXprxs4hoixe0eced2RZ83WosZ
Sm9JIKFaJjWG9sOGasanxOthdz20AO9FgL9ZtGoNNXY9K1BPXAAmmILA67Y6BgrNRFfe/gcNe5sE
nsrkK5lpYNmgqzzqS219R7sYYO0HuL8QXfDA2WDXVJK0LWOId52cToSmhOOPmDvZSRKOT/4L8d5q
l7moa3iveOSM4ZwSzhHZkByJ5lbgXGQeyCGYe8FSmhZfVl3n9Lg0JziAKEQNPs6Kt5ZxnP7l6ty5
MO0AP+pWgTSPeHuMai6MB4J+EWSyrmCCO9QCK4Ot5CRtHKnkDBnRvvzmQkb6Cj40cwrLhE4Ufen7
baUkYjXRBt8QFBng3p7kgKRTRo266LdegDmlAwJlYVLJqJK0CZKdOM+yhEa+caq6Trca+tRh2/lJ
FOu07ex2mY7xqYFEbyL8iKmxL4U3+x36F2gm5MsS4FeerSBGXxZCwhAmOCsI2QdKeENZtltIxAb2
kghGkiEFa6lZF2RdBH5UsHUX/dzPGigk/UJXbDQFgQu4DB1IyDrOFhHObWgoOSQuSMiJqtOyMQI5
3iCn63DCIGvwJx2NIjlW+f0I+4uZ3cJR0MppVL1C0w8l1KuAk0Aciu9ip+gIiapN/6I+9KlMLLzt
WuU/63adsSomfPdbKeI/47y8nlAO5Efw8Zp8yHBI1MfHTNofqwPdgaW9OBR4nvt64bauP/E7AALC
7N6xSgH/OS6yBiheMdChZ1TH9cN4EbFfGSkFwyyww/5iZfxPLn8TbNa2Ox21XWclW5pzRZzhUgbY
wlR2umlCiIdwI3Dm288+o1p8DhB3EwPhUTCvRuz0nUSDpSTP62JUdxwMC30WdW/RKZVvlwdOf9aL
Nq+/ua67YgA5U/sVM+EEArhPVnWNKIYJJOKaVLPaQ/fLAj1WM1Pc/7uPSjmrLG+6FV2AzseTpozT
l5D3+gNp2G6YKLm/QA/8rgH3TYwoU/qrhsvU/3tYushtUp0/UHZLTBFSaZAB5S5xTkDv0jBxuxvm
ml/qGzLhGnQVE4QLC7pkW/odRsW6WQVwx/SD7/UhBaS/6BjL80sTLoHtzfGY9IDCHVl4cuaiVhzQ
OokYdGWkZZXIRMg/Fm+U2OyNM01L7OKRHrVBSIVa7HU2zf4pl9irqFgekhQiQSWRYi89VHiiJ62z
Rk6IncyGoENgYU3F6y1IH5v77fYfmoeuLyL7Sdup+EJu2XDTpx3XPPQzgst5fl58MLiNDdFWeHci
1W9A9sKi91yheu4Tw1x/fBSmpa3OEta4jPe43CqcX+DOJHZCZ9JCKIg2LMl2Udzjz9h5SG2BkCND
KLbgmLZ1ppHVLgBqHgcBXerhaQd1z6Su9r6Ao04dAf0PRbL5binR7b/nY9CZp2AX/GlYXA4FL2sp
ukqv+lAKE8fzmOTDMrFScBJGh+qqMeIOWbBpbXshTnIGCapQI0JTH5YPMxveQMHeCvMfFmZ0PUdI
6TmzLeV2Vnm8su/LSkkDWCuzBwcHXf7JdvfAmDjOXUZgdhInEtX8GWbnBmriUZd3sbfqEXzMJXdS
PZMLiCzGr0VjD+LNGO/J60NkZXsRKKQGem84HYZPiAoY0/ecnxUVoeDtE3JzQAZwrosj0za4kAj4
O9AB+uLDy+IgDfUGCWHV3lZ9u5IZrxcSkgnXh8U2d7h5rfO7/u8uHBsSoAK/iqhc7bDDO3cshLDb
hdW1j+HAnpZQYl9b3l788CanzsH7Nd7xkJ9Jsp1xq2In31sEzDBgc6oklCl3LIPSutg851pTeIMC
m+4nOrt7kUj57o7X68FhCe85YuOMoELb5y9OEfFX7UH8a+drTuAhBUlamxJq6y6t6Ozj8ZoZEYhp
+AHOSzSay6ll55bXdAmNYYQXR/yNyBfqxgf06U2wqg/93YfOB+4Nu0glcY+cNLMcfzS0BQKVmr2F
uqoonSJWjCclcXNCKfZb4tL+8AjY4JmDp0str12qH6tOPsWy0ZTNmaCcKdMdh8Ek0is3DCtfa5p3
k1CNQ1xIBtpzA4Si+Xy7nG5sE0U3U3x/XSSoJzxdazUGGEzYgc8Vwq3alYikEspzu6dwEcE4LgV0
8SwySR3yVkVgS6VBlbz6nSxBYYU8pTsQNuwyi4ByTY3ZaN1Srm8r00/zJdjaE9hezWVaBX75XIUm
mpgsCjXGRHjIDYIu3gjFSMGLRrl1oFJ6aOVCFZDBHFwqSRfSOo/at1E+K84ZCNEeu4eYA7TjH6Gf
a9twkdKn+OKWtUU/h7XyCZryRyx9SF0ba6q+sMBaBAHK3BIEmgjIs3kZzS/FzdfB8JitGYy4TVX1
0XBRs/3Kj19N1gi/mI6bN3HPls2mX1WDEGHnNfXL9ejAryJqixLZ0J/6+or6k6ilWWgmAOw57+RP
2OAsEY+dDm8D/U8kgQ1/QU8qZUOVOWoFW2JYgo4dDt1LqNema3CSnFn208uGone1BlWFHJkiiQOA
VoXczxhpgSRSBn799PbqeoosO6yAwSLaIxNKfi3dB/HmekdpLjJqjRSQvoaAwNM5CJM+J3j1Vm+E
J5wfi407Nco7fBM13c0Raad6gHFOKolLRFttUVxwD9aHsFZ6jCAXV2x2leMxAmm7n5qpt33tfFKp
44mGCmM4M8HuHPWJgokvP5jRj9Le5g5zcKryzvaLDNEWs/3HmGAUIXK8b33/ubH6lzXCVZeb+jfd
ZCAPOQej4MbAjBD9VvPL27/uTnbaKnsDHU8SEB9KKo/JNS2GMvgY2NgifPdvW9J+knK54OOF1LNz
xfP/ekQHdRaWL0Ze4ElR91E7xGxaUCL0iInpzIqIU6U2NkACZHRbv9xbdUmsVdtxLtefuMHJmPn+
wj2tytdvm2+snKaKCxRhhm45QgFpA2qqr3dD2svFNkye6jJ/Wvz9e/idms6tvRoRCyb2Eu72CYds
NfWn/I+/+KSY5bXxCVwt9j6jlRJGm4BIyD4oSHHhZ8cUL5rthLTlQOHwjUpcZs/QYU7XlXqGVrXQ
GKjuHt9O/KNp2Y47ya/pnsqGn6vDqK2+PFBxSSwoZgWYiX8FuyP7KQ4QygG3KAkq6yfJzTfVdy3I
F9hHzOxB4Z8pnroQzckXAlCx0s++j5YUk3ZHGqsVAY+md1tlGix968nqp6TTGwGnR8Wr+MUoABnm
OrvWWWbp3HCpC+9GNcVc/C16bjPx7LDN/4spZUtFz2riO/XSD/NsRq6661sINI9rjv3bIgJiPGeM
+6gZTaMm7+Kxh1j0cMhWn3BRi9JDuG7Uv7v/ugwLD/efwOYNx+wqov8J+ZZj6Ne3xlGy/XYeGCJV
oXhGJa8WqvLU6EXaVJN9Zyi87bboqJqtQhNHrSPM1VWFZZ8C5MWmvvZCQHkibAey5Q/klai1+WnA
XPFz/Aby7Hjy83VgwPEr1onPNbTBSuKq+/Q/n1zhueniwlZ5ARuMzdheWsgcRroilcrJs9d+s/ZJ
ZX0R8pIBiWAK75F/tNwrwXa7i9CbzpaNeQsgcKav8MvoS+NNhH7SVtNnyMi2k5H80UujfoSFBeZd
54EeCyn7bhUs07lh3Owo+2rJCXqNZtLHIwtz5eoRX010TGsGP8dNjKv9S2rlJT/khUEG8Jsnqeqo
bp70KEO/5S/om+5ba0EBJ/f0ETOPOm3tXzXzo7No8e+94jjKuwRZlS2CXhBc/+EkD5e02N/fqMyw
Zhe3r4Rf+lOBMNLaa0AsRmBOADTXqqGYy8Q/tHaTgJayT3+NeaitjADLnP98IWVT9tUpWqWXNb/V
m3pWC/P8hNzHGAdiZf8s5YiUGheqsabnRVHDsPdwkeIgDUgah0e6SXgz6fUFKihtocp5FHeLzCyN
G7LBBKvufVM+RGhsqHu2eC9F5DajtwRTEw2JH2lzRaQD5rvEupJ+/2cQfzQ2Dr2862ePCT/UhxmI
H74wDhard2DCGZErZYiEjs1sEH8XPJlT6OJ+NRlVwCiuwbsMg6265LEXrXgd5AL4sM9mVgjx285W
o6RSYvZ1GW9pzdsKVim0NSMNMxUzHeLvVDvx9N83G9wx89yJsUoycsjJsIZeqgxpGI3U+laNw3x6
O/p5p3/3SoTCMoEnFxi47PLcf4iSFsPOoYEGKrvFGHPo9r2FdGv5FnzAHmXOiPEsJkoM3zdBhW2v
Jkkj4CfdDkujQp6Jkuhi6vEkVsjXjn2EnxBeMtK7/PKUk5Ogc5onGSBYCyZ9/0ausHNCLGP25j70
J0BBaC6v1bIVXDDJdGR+WQfysWIPolzweYqK4RRPAI1ML5N32oKYvyI81LqSTCJKsIUExvNcCeCd
5ph4cFwcgHQYNF9Y0SE8qcu4zLKFn/rKvepriBjGLsKRLUgf1/GrNbmkXNrjA1YZLR6+XH92nl1g
/CVGTaWVG52bP7mcqA5awhnoM1tngVFtUaGipa/xRIMqKAZzvRXxkVMFGdtcusnSOqjDmWHe/sha
j9LwvhibQzcfw1E/U8s57gye/HZNv2ZHlGdXvOUoL2Y/HFUxjHiwDsA5VnbmGD7tVD+WEqpMPHVQ
jhKv1SJ6nWUgAuDmjAcJ7t9EKJWpasPyoIKhLllffdKTKCxF/g3JrvOu7dut4HKFwrygSVvUpFT2
Qq7HjZGLu0mnGbtmEnfB8RliPoxcBXDW16WiMv0JvKxKPDGqyf/U1QWSgjkH7JK1LnWKgMaCO3xp
KhThEH3dC2PV2qnuPT0KRJv9gzkBGb//7qMuPqXnEPQvtQBXmLQQTWe4S2JelXq1VN1E+vrxy0i5
RW5M5LaJOuo2lYJBrRr9rMcuTgJL/bO2FVJ+GT0/bQFyR+nePS+CnR9XiyTFhTKKSMA3Ov54ECvA
JOL7tG4qeunvWeIgQPxzOVhnw+W/hr8C4q4Vbe3EybiZLHG543K4mvTMRuRBkb97OxRDCPDi7E//
OcUMNGbmQDjfhBU8VMKslsCUKGS2wvz2FVjxEI5CD/cayANiznsQqZYYbzP0dfNd/OBkOIozVDMz
qaPIkbadhfz3WUEamkpUY3jIAq2o8wOsWUsS2Ebz5cVjbeD+lKa+lT0ZiBwVsCynzeoqnAbDFtuB
QHo/QJKRc+qXfnjiW7vS1l50uMAInBwVGeolVCXqX88aZ7WVCQr9E1fOaI0nVM/v3ucZddHuhEqP
qsVbePMtx1FlEcPJKhu/wjV1WoUP+fQ1j0/blT3vjlLjxaL5yvsQB6XHvB+Lv1yu7DNyfFBNoLu5
QCPgGd3Xds7x/JizpQ0fh/AxY0xcgH65PbiMZvaMIJK8ZxCNl/7QpsA1KUvvDcoxcBDdE09T4/tV
zaDJDSPbktZIlk68/4wnBITqDL73ccR6AxBNJwtmHDUV1LPvEFpEU7VSgAm9YQGTw032+4kt0rJL
w5liZkstTWog4xdSBzmHmRIZgKFZFpdJq+mRt/e0EURtomhOkfdyBvwQXrcHGtnfDIMCbw75dpCi
nlWWDAC8oXR3k0zkEYDXGVaszawJMB81ZjC5s21hujYx8FeAPLkJJ5LxlhboGVrTJiz35DmTIKDr
9drG+SdHHlq06Tsa/E/L5tdiHtKGGDpo0xuJw6e8PamrCuKo6nLs5XKdtb58PHIr3oD9+eE2uO7I
OjfXcORfGsvU3mYyw0hj9ZbZdtpDKja4qsYvxFeafaLBc1uz+2nsh0giFACgmTDTavBPiQE81rde
scLIYR4o2LzqoceIr+PANYBl0ZgDZuUB9AwE4sVjw6KXIoWrWU6tT5pnztLhaRAh/PA3YpxXutdD
yhf/1N5vISGR0ZWWzEVvg00GMGT9rhfNfjxRqveE3CYcUSW4iuSMNGeO2oNAAQXpObaI/j04ylJW
yRaP7S1o2JE9jfQmt3hruVEPLIYNVYDb4CAmXtxlbYkjVEEsWCzqeG1UE/67bd76/Ofev0U0ZzKp
AlGBWViPTF7U0JkSDaLUK1uR7G8gK9d/esi88zM7nd7HWBTEmd4qT1T7wMbiI8MznAHgIFK5OX2n
Uf+D339Uhf51j06iRjluzqCOJ4yD6i4sQcBojy5lm+hAeqzxzEo8GS47nmgMIUnIQeyPX01bvqEy
/P8MLNbtknDqqmCr1XwNGob7eqebPbP4BnWJz6/4vSs9iYLlqCcKG/VaenJ4v/yqbnybzXDJjAhv
cAWyz5KQL4JQydBMSnAa8BXb53vgePrI4Uw2uc7txzYnszyGT7FDKpuddOujyqLOWIfhtxIxpp8u
fImGUdxFHkbD8eJxY5hiEhVZUqtVBsMHTqNhQYIlLjwsl6D8fK8eV5BjuGG4lgtzeJ+X3w97Vgdp
p6B6xvgtouEOSkhN3HPQ74mLZn2/OnlBo4DQxt/yaIH1E4T0T8g0dGgkGnhq3Lqi12jE+uzSaGQS
NEG1J5I/sluGY9csko40Ealtfp771BmgSq+t5umHf6TRxWhkxrYGy+5nynzuc9ROtUZh6Z+XszJf
aob2SWGg32w+d4+z+x1bwI5KemgBwnegUDoTKcAT9MaoHh8DM7xLVULcJNvSlCiMXerRYCJz2Le7
veIujfazMliv9Z1DgXbYYZjr8U5fpN+I9gflywmx6C0ysPWtZKmUD8tvpnGODfxkZaccTfbVajYT
Cnw3qQzkWJvQfoFzlvPAuZXZvkB7Y3NyWnvTVfbz6pGIsjjAoIZvDBoP4J94mm27K46huXDB/ItJ
25zP55S8yH/kpFo1GGTrbPGHhsj4puwrB6FS2I75s2ogXYUfHZX+/z+4XhVIHHiu683bWpBzCtNK
YRv+1HIWI4/cU/dVXH64vDNcypWLiVIkNlUeioyyG/spstLYK0A3OcNh4GmTnhXXIBrDkFzvOClP
L2HGU9kgU+Ag/ErvnmPHXrJFAO90OnrWexQbDvMmIF948EJ4dyvF4SOh0gP4nzwDnnS3a00qBTfd
OmAXY4O1INWWAOqOPBFMWvTwNRxSbD0D5eSCK7p9yZX9q/CFqMRudUqg/sNn0BDqigEsswfQEsGX
4pXQytesbYRpcJ1FXnXQg0XU0WkfdSQHDwa4NNWaben+SOyS4iQpAbNPmTTpq15x/QBkPtl2f6K7
C0KPQZdf7GVLg7hv1eCwf+wmYZax84PwAKzPoc2bi1vzs7nffhLdkyu7N/wyE4f+2tq6f50P/gU2
DjadQlNe5nSHDJqexF0qIcDxQiYfLchgOff2YERwUrFcRRZQBcM+LNTXeFK6L4PI3o0XI/Jb5vVA
L1nxdWozf+vKHnHVzvW//CrdZSYgIQom08MkG7HqV3McacRPV6mqi4FfJnBir5Bn2NSAeeHV2yQ4
3P41cS4uIDcf07u7W2E394M9I6b93TXK59RdcJQRJ4tOQsM+IbL9Odkf6JIsxKiNFjrVASK33ys5
YTTvE2dpeyNuEKnrGD3El2OeAq/99zP4m/4s0O9egiIYoVGeL/RdtsfnppSNQYOkI7aFheMPqOIX
n/ib0k3t0o9MtcsT3PqKwIRnK9y4ByUnTAyej9DAtE4Zht8guLSQaLLksJgon49pCQgJHJD2RP7B
YrEPG+Y3spFAcLdUE54duEW8WFTWEb/mUiqBWEk0Rg5hIK8otXPNKIGGHDjmuGSS2s49+mKmSHgf
DgDeRN0drPa6uE3X91BCw5jLzrKoicRhhMMllp11lIoPi9Do12/xHKGQr94P+fybBrDTFfgdswUB
Zt3awBHY93biLkNU9FDkprJF7CTF0OuKDTmSXiPO75h51KZDYVjgQauMmWmvk6EXnX7AI/DPidH0
rPZV5ECpnpJy8OCvM8+P2Td/MJP13Y6ZcVxmIVAGtiu8yuLIRsngaTjZRf5Io6FLV0BV/4htvbPR
81FsHF7oEpCjTe3Ub4SPDVYM/02M9mUm+fF4u7/E8xzLeOA24nCeYZu84gsZDvR9u8kBFg3HPB0q
+AQ4PN4pUKp+Xjj9uU5dMpBJ5hH4Q3JthExwtpGma5DdLDCVsOvdsLsJQxc0kiJTT3lTw4bqL4yh
ZzoEP+d3ASmUcfi11AaTLg/ZW+pQf/hSGtpbZ0b3IsP1sjAPtlbR4rLEXw0tfbZZYicdQ3+5HWEj
xXpNnTpAbsR/g2G3r3QqP9gBfYP1hRWWZKCx79k07Xpapi3EkNabaKMTFijIyRm+OjMeH0xC7ouy
hF8G0qy6oqSu9/1s4xvj1/9H8/R5BzQPpgxRl2X3ZSzN0ID0S2D8h5qtm3fDryA7Q+X8m+j2/h01
wvGKOu2PvR3k8liR1v/szPYGsTmNAeDf2eHUQ2B0kw1Ckojqi++x4AfKk1C+lcJ4ynRbkJoHPbLV
BI0/WXGJUXq9+iNvSy1z+zRiVwuRBOOVil9DZpRo0P2WS97aUK1mfLgNowjDYRtOPXGZIe63GZcH
pt959vz+SP2GTq5YtPiSMPM7NAjJsyZeD8tUW68R25u6Dtu0mF6QjpRCRZYf47W6sQ3EV4e5iAEq
vORFpZO7kCclkOHbluCDXWqRmGVicPN+K5lHwUINKoECrNe+Tht6IyqODk0ijcX2M1SH6EwpD72G
PS3kgdHsXEaIQ1lpRJFq6xVN6z8DJQpTuaHV3JbUg3GUKjN1jltJpuNHq7w5ctGP9PZqkJJojhFX
i96RhLrDibWQ+ubLYdpQ92dFmnfhyUxA9I+iesCvjnSv4wx5QztLjkq13MJebqH2gQd+XCKK43Yx
lU0+SOGo2epnWaQ151XvklN1Irs80FrWVF5CwOUw26JWMR9Ubo44yg7XN3U6wGz9+vQy59kzg38E
Qf+U9jpFM/kH2aS6I59KZtOkk4OLZKLNbo3IxCeFbt9fa8TWZ2WNbSWwfGdoQ7Tl3VSuA766Q4Hl
kkYXRo0XEsqWiVg04bzUkwfEOJ6oxi7BIxHjehkUDVS6oicESxtjlM8CwWqvTDcVFIzHMrXx2ooe
N9TXg43tSbhxfSRTw438cxOTwd8Y0ifjsepFAj3LrSeAKFe3haTxvRqUgIAUvWJxnb7fXKmsiEb4
RegBzMxEdTfwQacpWe6xlKIikABx5g2g6Mwy9EwI007RzdDNP4rojUnn/80YHzMNBFjFBW+1OJ5u
qpJWSTQ00vufO0gNan8gB8PTYnK803LwAHtcDoisGudOqPBRH5bDdeQMVphm9XuCthxzGxj+vIP3
AR4ybOXlUQ65+YxNIWc1N7vhZCGEx2I2bO/Jc59IhSOuGKhP2eGGVTtcV2lVAOAMA0a9v0EvK6Wg
vM4dJ3/3r2fE91XwNriJPXF8NlNmnsZgdwIFqZqm2mPWjb2rMhA2p0WgbV+o+W4Sh5euWnMlhQiR
5aCj2whGfkx5b6viUyyQfWZES/oatjlQG6x+oOhHOUAeYs3iWp2zJQl5vbcO6R5XaozVmLo8GJRZ
4PLfmuNvIONy4MnGdauzfQGtYXiUhfuEttG8pRvtJgM6Ycun8XDVqJNBKazskgjD5hl3kcqrCtsJ
8cHAmYeNuxZdJmbXpHTivdpeBC8XHu9+XGF/zliar2WSX4QRw3MnGcNLV9hW/gMlECEoTAOPDszn
ZjE8y/ctweWswh6k+3Osb0pkEgXrAZOpilWD0xzuHD4ySBx3EtVo/dCHn5sDvNbbNXQx6BGGRTNS
w263cBNv2jeRcc9ztbr3TZGfgUtFWBQtNfH8CTYHLIUpLVbfXhZMwm0hbK05G3ZuPo6fyMXgmVZ4
YTdFLrpg6cGTZwmosw7UI0pSQkaQ4GJ97v1Kql5JtI8V2HixmKqqgQrV5y7Bvmy+xQL53p8vIRf9
F2+qT7nWx8C2r4e2KtVPN7qxYC3c2vWywAku6M0QMLocCv/GTl1JUBWE/inqgtCEEoZYFBkMvh9z
XUEiK9qkfHLkdAEcwekv6xIi+YjCmtGM04Q9JQThCPX4AzJ8afs0a4MYZfl5K5pKwb7FZmNOUshk
qsayP5Ew902Fh1UmIYvfOkdHXla+wdbtZxZINAWlroqhTWIqNEtY+2Jlp5oP5S9yDURf//RMbIfL
xIKNHp927eku6FZQiWis0uQWvUfJcW+QNIHBH9cCntmkxeE1+145MPSQ2mPsS7/sq/3Q6+Li7k0z
hC7wTWwQer9U8ZMnUfSaVOkV2xXRFDrLjnxEL4NA7kXcnmWZF4wu9uKHjAZR4m1W3rqvpTSVDYPs
KW35b2ro+77IhVSy6dCP8O2caLh2cy1oHzpUE4ldkG8k3ZqE1EEveeHBv94RTaufAPjiyB5vUltP
UAaPMflpLb4wS/6mHs/L0k+vgvkEmWJ8U7KOZ4xVTarhV0yPYchD6wEx69cy7pSgpER+54o8jCRQ
cG2+lMIJnerCRMgHeBhbXGQizartcnekirXkiiJGX2jks7RIR5mtkBoG5Lvvsvjdlcb5/DDU79zR
8PDhFugKdRw0+xmS5d4VUB0N4dFHCITcUoIhrn2alHbea9u7mwpRqqVZ34PUsEjkjYLOr8IsXIxo
2T8ORFX31J3akNMhCEUhKc+rO63AKge5EYTFjClEcNt94BhEej4p/pH4W3NXPGccriB+WQl8NRgB
arPU3CtNz/TU6cPWIJufGcXMlsGTWaE0rSRuRuwQMrkcb/rHEDnDMLmRFoyA4Ojgwru9MUg9veDc
qf5rfM+n1jN+Flyxdeo7oUxwbn945M8C7Hyqo6IVZ5+aN3xP6Yj61+/X4ruh9i1VMuiB4rgeD5O0
nj8Yfl7T/lBiqBSdGN3sgvwMhBMr2zg/2O4bbeeEubeF4d+krKvH0RuZtIe9dSmdXKwgyJ04RAlT
291oqTROXSB+qi/6CYAxiLlRClyB0lYo5dYK/S/eCNVtmFUyGhIScgECy5C4Q3rG5uRecaA+mWFb
ipslQlcJERYJtazDGdrMWdMwzu0k+QgrQZACciMyG/4Nqw0iueWSzf76VPBsCAcf5eKy10r2J9pO
afPN4ykwnjuRNel7kPoVU7DdNlDW9pOoi3NKBDHB20xSZkt3JNr27bvx8q6Mm9aeMUc8jUzkYa+t
L/D1h6pKp81BVJZE6pnZobMbuBtiX5S860eB1b/svVZiki81hXEBtx5TuC/O0fLmPlssy9ahSS3q
87w7y0fqOQkK+wClKWo6GSSrbfkmSrZW/YsX2EomdI+/emXAOGEh09jKfEe77457OQv7ELBwdAcF
dMc0/gx1NX3UcRvmJAFtMtM5fVexzNck2ZyCic/4rOfyrpUkxatQ3aItDtC2CPbhU34kQRzx97TK
82Qd6Ti/qWJ5tgL0s3slIuYkM10Rn0hhUGOSsmG/bJQZ2J0dgeWLX22XrDAg3cAor61DSgoe2PmB
QkMg4StPv+P7NR9PyohY9UtCGBxl76vB8Zhe0TefV/84837JkOanGZcZFyFEvVxDJw6C9g8FjJgW
BzE1ZXYKs+bEBql4lFH5dyWL8xKOFxHi8QHHUKC8cC/Dek7b8ih8AkFv9yUotib+sayCO05PDhop
yV8YW/w6FiJhegQysScAlOLTE42uT7uGY+45Gm3odsPS4nKWQAW+V4GW9UQ1Hioyk+UsBUEj1UrQ
H+kcnbsBLNX3zZuuFpuQ5EwpxLDkYLCdMISsTf5vn0sbLi98+AO52l0S4rltDzFrhzbb/x3vGD/P
5pl5CJhAnnduGzzPBQyEblpVwLvNbwohsUcIL5ObS9s+jGhmJnd8mxUvQEd5DSQ4h/ie6lXjh5zX
+Hm0Mk/Arg9NIoCheaNjcWZOkVFwHpR+iuCzhjl4XrN3kXjaqmmkoR28gEOsYhvz58gjYozISEWQ
1HsMyisSaulNQBhexug8Q16S/iW69u9RUt2XqJaiwQshKs4vXoVXh44qsVErxJmnP7BSfARuzTvh
D48TdXIE6kyV3r3V3zg5vjVJS/Dr2ic/cj9+dBk0uhIM2oilOC6OgmraNvvfm88fNfNoeteZc5bm
fWuan+TSEOF/R9GQRSYl5c+QZW6jSnSMDn7tWjmhzhG+cLRYpLXqx+bE+bs2nYy/JqStLEYe/oOy
UoA5Lm3UEe2/a0uO/yeAD4erGCxrMHAq+aPVE8maZv4q8jTSLAZTdqtYq07by/Namt5ssBog5quX
gDYS50BM8RKKnd1VQbdDD2CW634cr1miNOSN6IRyh4YxmDAtgWLvyFKJLlrrVAPCDd10ChIev6Y9
kB0F1GUu40GpPrB2waJlB9A9vsSdhPgFzzyBA1Vfmqi6sPWvfzfIT9x8q6QmwqplL1Kp2KV/Lv8i
VmvUZK6cIsfkBeUPI5mMCFu6a42845kGqv2TdFSRr/9I7vniJCVmsGHG2Ya73sA+0rDI0tccbULf
pyDUjCv/9jC+ofwtrlZ2KOc+PsoFUuF9GIIIGlmAC2CzWq5usMLO3yJTD1TniruDhzdxnZnVPlGO
lY5o7BvLdmCQljZ8Rgzaad73pdKYJrw6N/tPwX/WxDv2a3xf/h43Ixokpygs1WnD7+YyvCD6z0Eg
S5DmDSnSnMH+GCFfpP+7gTNAFzW/sbG3l7eq3g+gYZRVkbzJEPg+Mxj5YYqJwHUqV38h9bIvpy5Q
Y6KPzbMP7ly3MbwCPG8EsiR2CzYSOMRQ6siUHX7zKQYBkiuaMnA4skfNPF6N5BbSlOLOYC9ZBX0P
QfyDYRgCK9+PWuF11eGfycNMjt/8CgdjNej3AjYfUFK2PYniECpNt2ksAb88d09itNsOcqJTo+88
mRaYcdpnUc3z1YSoSVvN+m/2GkIhcmqbD+zC6yKVQYP1m2ubSu9TygVF2Roc75KQ2Ph48QRuNzTB
zcFaayriCpk8ujAkIjlJ2YJsDYXZw+fahOs66tkUVCD1H1SsFj9XXFw5EnxuZIkSCrL4AaluVcGh
GXHdqmylB12xSNOni/d2S9WFdittvj5faHGIqI9U07KtcZVtDdkFZZku/0MTuBgZTDM63kwxzqjZ
/hEx9UWpNyCMJm6cQa3O+4fk5RMPwBeNCPkONRp3nxC8VPd+nzzvCo4ei+sqEzZ61k5cQoM/2Qzx
9R6kYLLkc/ltriBb/5cfZ4As2oLkfnBu5+pT5v8WCSyWUne7kS3K408q2J9aSr/WUqZ2A/VB6kgp
KZf+R0gtb+i7HB6jx8SOlSnegR2yQPKAlO84gpnh8PjCSkA2eDv+sZhK0ig8BZIq7/VgQCLqjyWZ
XxS03mhSqOMG9vLvPuHjmsnWhBhoEQ/XJaed8Vjf2KguBr6tf9iuwMebsHOvnVVlpRgBMxrSLzHD
rjGUzTL9xWb7l/xDO9IoUIdJgRwDRpPgNxAlxl9HDMgX6sLBVC61AkSMPxQPlBfKyddscNS+AeFG
0KuHQrPv+u7UZBjZS1sJX7YveMpjdcq7NGlWg+M5COZwPRm8GA5Nf8uqwmLyN1bNQOtT8dCBzR84
JMYsxLst1d/coWeGf9so6+UGmOrKRSY+dpeyUr+e5cosaCSwpQEdj/JhWfDfmTeNR452840aiQ6t
kZopk4KL+6XpqEQcGtUZdoxauuP8qFI6NeQ1WeeWBIMOeG7P10kqTf2yIC3OlGgHCi39IRPpJWkf
QASkTjeUuE7qPz2EI/jDS8NwM7DyDeAYgF7ggM2HiZjeGAnBxjiRbyJb/44ZxnyzuVTNgiAQLfCP
hbvoQUdgwZh/5HNckbSQiZNX1nFDDYmtjFiUmKtlDoKa63udPuAEkRd6Crcf7X5nrFdLX6b0x0QZ
0990Vgnnmtz6LvagWlUACvNz+rqcbLRRGympk43dmRYUkkj5GlREMbc71UCFx5lGURTF0PTiWl1Y
GyOQBrySDq7A1aFjC0tZvVHLSaoNCinpCegh3/Um3q2Jn1TJ/AE1yWn8QIsQGrFnsa6W5fKXAVyf
bVvWVX9XpyAgcooWgeJDOGkA4lRfnlaKliHX0L6sOzpi8ti2jrJiup7TlmbqtCzdnry2o0JLQ/e5
fHgi95QLpFF8jRwRy7fPNs8zHIrn1UYW1EnyPerlo4zDH0ZtBwAaKFvmE5GFO/IhO7PGQZoSmSJd
CmO5EgsoqV+GiFmVUwMClBAHvM0+8Gd2ibMKxx6+f1aL00nLfCeub64QhtGP/1f0lCT9/bHX46MD
iJycKUkAIVs/CRmy4HzdjHQ7ilP+Ng0gIPubxkNvWMB42LZJ6ED3VlrQAjtTDMZbejHFjtyFuKXF
qYg/PfUvnqxjTs5UUA5sDw/T6cf48IwdFtF6z6regF12gnRbwsaulhKUhbrfpyAloQaxCLXACXby
F5tov9RRG+W/vSnLg+ctWXXe+YTgzWGmk7QL6/NpVnXyRYDnZTGelWimRDW+AfCJtHKF8ZAKv3FN
PJq6vhc5yFXunA0NMlYZ06TRxEcGE5I/bPP2Nz4S1XPEnfaQsFMF42gjry7rik3W/xeSnBz2zlEi
LDZ5L6oApJ+++1ZpSGr3dPnvcMMl+kAlcRozxo+jhKqRkFuTNoooVFSFbqInV02sPiH+gHhyhUQj
nCQfmXlYg5ib1/mnjIEH7pgc7C+W2xM1dcM+UHjN7P87H2HUELaEwq17s1PD3L3lbdU0xlzSnfXq
10upVgNXEXbHnKC+cXoqyib3JMTuuePi7Ei3RnYQeRJQkMi9A1mpdKHuLl0Q6Rg1AMMYQOP+t/9Q
9rqWKf+zFkG8EoWgZXA7CuL0X6nCy+N2qlQaGUo7lkS5PRCOrFLTnM9qNCtpYkG6B1YMm3f/MxBJ
daA5p9D1VsBAEFLcttMWT6cxYOxJXTTDJi7nq2leJf0/seXiU2l0QZTx3Cm5h9EsxZ08V0in5a/7
hKVmVndKxYm+Pv40lFSu0Hi4f1F9meNrdDqqEClnUpUhgBbTfVeQPEa8vrQplXuVGD2adhfmxIEw
cUYF3CWRweehDwfiAK3oz3V2TU/z7NTuKghqjCFaNxCgjoFRGndKgSufLtjuAcTxiPKb2f35KBEi
Uf1ButdG7BlcHbkRBeI6qj8okVOo9xqnY2hYAgzLDyTECpSudaEvAU1AJUe6UI9m/uKgjvsBf94X
OY++j8OPEj+0DjAMcg9uLhPI6O86vR1XV5GfD9UjIAa5CIYwn5iFghm5NNTMrxNuWDMWC8LBRoCB
mxfhTpV9qhMezjRSBJ+iVOeer3/UXxgofNw7chmI9zIDgfVAn8hawSwp//yt35Bd3QWn+UxUMADj
YtWTLhFa4T0lRehplzd0dKU/wp0nVH1bnCO3BDu3HDUvkttBCmMJ1SzqwMuhMkHEjRyozwShYPLY
KbX5Ssd3itX3oU0H3tsz9ah6TwaLCu4IgTNez5MWI3EdAFkNNY/xAdyMCiced2wBJnGHqbKRm095
P9kmfzLblKDs+YuMu5/a+In0CkLS9cCbyceYcXfS2KD7mCzYq+iN6QgC5lkysjKtS4xGEmE7WoxN
v3Cc06WmjMP2YySd2b6CT3LkSIH2CxaDAzouzKydiFsjmO7sgdG7jcQ/whIXcQUJTjUDZyOD7zYm
XJCifEzYI4dbnNz6W1Ea/habat43cztrlhuVg0nYjJKCl+xZc3ZAs7+2pW17CYWXSZYhCfW0gNpw
BQ0vS6kFksrjkyLcK4S4wTm2FufpvCL9XRPYRodcG4CyUNFvHYHG21MahBdAu2us8+NlfKMhcKjY
avvMb47N2VbpFLhknHQwKN2ItjS+nN3MKpKx6pzaylVr7RvFqPdX3mHkgVzmjuL9xoGZ9XUfikqs
7oHG1sSyqUbzRb4x/2PlpYCshlX0PBiiQzV9EuUcrmLdf6oth+wGpm9JGrwEqbrNsHORbWGORxsL
6bMM83IsusaVOV/jPtxx01ifUvOL37xiYY2wUfg6FrS4e55Gr448ETK7PdWv+ugMKzqKZx8dmeFE
DJ2/EtqZEm58kymRPlB23TMnYPEoXh+5SgyL48WvqRjyOt56S8pHpVkrrHVVbl+Alq2S1vjlQK7l
53h4xwawFBpcfVMCmE8GDxzteWa0I+Jzl4Orp2aVO92T5YC7P2ZGiUp5/ADKOhEFfHhCA1H1BxCF
vvpjEaxDexr0vK9fr/y1B398NOIl1zc3zCNtL72cJSwv0l1iixI4ZwYO0R/3l/xqIicdwhQ0Aid+
MJJuUjfGwbkWgRDWTqwFbnsm+nUMn2frkS7olbl9SH47BUX8yFmFZxADN8eec9leZSM9uItX6qzb
lqaotGwKAlRaP/B/RskjTVhNK5Heqd6ibnni8sTuGa7HIYeCwnPCu1sREExLZXFQn/hLVAlGkyws
gaA7JhFKjoHYWsRq8jR/k88aNeTJFcko+Bf1vryyv8TkYbdnZX7Oh64G3y4pDVN1KrsvzIjmk71p
rMPVTzvMN3bhEjyp9Q8YlZR/KddVOohTZrkuli3qSoHinp17F4OSvBdgdMLMTcbr3zo09t56Q1wh
Lr5ZTnoRrmfB6Mu2FCkEjfjoOK/YtM9VNpsIdwbpx4yK9IIVbHA6R/UY6cORGxR3e9ao87Ri+A+5
bInV5SheVuYRveJgP+Nwt4Sb9ryDzSBldmdEviTCEup0fOqeyQRTuqHcr4JytdZSu3u6OrX7Ic5N
PeKD+Xet9lit4XD47lBrf2ONW3DVo+luxFumrd+6IXD/VKMLP9DtI0SpPDZcz3dZh9Bb4M0Piooz
ynrLOonGyc12e14xtZMBa6UKZ+nbx3uGcE9JGwA3b6bgAT/x5av+ErKMSchxrY6vC5syNC8K1wLa
VpgZBoc8mxg7f4IC8mE+4lDRKt+l6u1fO/gtxrGOHAMK8kAI5u8r6SpIwWfDnnolGmIUzD2SP7JJ
Erjz5QgYGV4hZejttzg3U5BdROxLSi8l+QxILwEvZ0H4l/b76xlggWUbGUiRDxdFcWJ1tYDroOaj
0xoawZcBzP1b34ADUfTCmdCyrkwac/djw1ckpe4bregrVCaz3uzrb/TyY1O6wL+s1fuRzhAMmqWH
OSlX519pt2jppmyj2IPiEJ/hYbF1bCv/aqMiUHNGehKwVjTiIH3D9WDwFCaXFWeIsAUuB/A7J4Ks
5hAwdmCEI8P2lrVRocit7qP0IOvmxMK5VYohaN+mp93UcvTyrbCZyI5EYfy0QXaP/AtNe2tgrXbR
ZSpyGa8KDP9ZqoSRtyayIhcEtvPalA31H5hQYAGEm2FMLtOeCaVTB+M6OpVnPSftSHU9vpI+BdXl
kWI/KiOKCAtR/A5KM4qS8jObjyq+myJs+ELDi+KUZR4YWwrKtjmti51+88qjkzdF1QDqI+nezyQE
KuHnM+leUQ5zmFm9gcZDqvCbvj5sGCOf/prGKhaiYJMUc3d9UZctqAaRRqommqgFE71cz2bmIVsH
7PeBGqcICw16yeUrpijANtuvrK/3yy3MlKn7UKI7MUb6hWdFImVMR9WshugdtIVIw92bmDRukNIX
miD9uKzs055wIHgKwNl0Uu5E+RGojcCnOXeU39sF/Xa6sYpQ9ifSowUZdUgzKmuaJq8Rd3JzpBLc
OPsr639LeYWwTE8Cei7J9g5sAT7xOF5jtQ/O0o+xjbDLX3B5npHzs6/uzbOu77o5oJsAq3jvKifz
VEorm06UWjM32Crh+3um1umQZSVKSm1Fw9H5OHiU96UzPgpWbz+pDeB9ZuwR8fAu7E85vXNK/xgr
qm/tstJ1kqEGwOacVVkA9PgmZeyFQP+AQiU4Cb+fI5Obk5QWDU9N4XjQqcn/KL9RxAy9jXrB1n7N
t2svNJGzqzjAv9RH+5fj0N4xCTDlJHWKtiElw/JVfp8A66sAXNfXDL3hhUKQy2+qqGYsaovo8sM9
Snn49GeOgBVYTQkJzeWoNnLLpaXvzj0xLFNZTmgdk+1SEAeNR2vCb4mZIJRVOAb2+JRl5giPwmlF
CUExYDdrP5d8nEm7/B/3HbUDJnwpkRr5BudO5WMDdhG5vvjFUiE/eWQvn5p39FFHiWfNgu5tddW6
0QRiZBd9HtHq+fLejDVtsi9dIv6WEvOz9bDfgWiaFWMLFWEsCB2CiG8N3vQ8vH2BYgKztheSFDES
luNiwClC2H65xiv3f4DiBTN49CL0/5m8tjxMs3LgpPqWqNrjof68zvvuGXhpgfNrEzCiFX0h1xUs
JgYWcinJTeKCBD1GoBhaCcvO3vrILO9kKp/vMtrJ7NVaEkju4HyIStle9ijcGXLu8COQGi/uyuq4
OkgW2mNd6roB/DG9NYbuFWNYMJaIUx2QGa7AXArnuveSvbH+ApEzSozCMpTlKBWgjxFTJtLUhJ0Y
EQm363Wh2jUMudwX/EH5Ddk93MpOnz0wBjr1AZ8RPvi3dRKApHpDFE64HCGGuxSNdVfQMJgzhPJa
nJoMbvwTwkBo2M2YJY4k7g/u1aV59lAT2E3MLKH3HvdzpYFmNJIiYKqqwIjUbYLvbAGJkVrlpGmO
HdFDf7fRxy/kY6Cd+FX44EkAAx1drA2RGfrVZylpkB/SQQwvElUfpM7d2lF19op736KVyXiur2bt
ZJG0NVL6DibX7kr7VS8NNeluPlSn0ySI2kmmDZfRCT/L+IFJzgiLAATpnEgkWrAAnYnJs5JF/g6M
xxZqDLUrfqT2+B5QQUbsmurK5MNRIzgyDV5fBBm8cubGoXLs+sSEe+iYgNMY4EOfw7YMXxWGqRWp
T6Ncd9kowGiYElbuZmcEJiLMoLyGkYHmw4f8PcA4YvrQFn4Cq7Q9AGqw+IBZkNF+wzwEy0hmznDr
+pi6LiOySP/E7raFpyK3M1zANY5i0xaHGKHaEvKUPqWYaIsxi5Z9uv/mxaES6sggls/Cwnnz2pYv
ElYkz7zUgKbXuaX2ljjSBv4exjoOU8XOxEfvCYVKE+NHBL1MC9BYkgQEDGcV76xJcD7Z9gA+Sng9
ENOm32bBfsSqGVC9+q45o7QxEB5p4hgqKBnJCGaQudUe0Gq05qtiykKGRSitdnZ1WLo3wwqJt/Jl
PJeb0hMleeEjE2HdtV/CN8P+9Pwbx0647tUTibHptyjqxFSwzmuKRWb8Iqo2u41ADPESIeJWKWVG
cIZGlGo6CzFwWIsvDkcBhkZW+OgsQ1c/p545vAKxMC4D7frRwDNFiVX9J+BNnBG7v6iVn4lIM1h2
tlMYoDTJLdDwo1pM0o/LTi3V5RHUGS8TK8OCP8uC+MG2M65UBFEOOCIZX9NrAmJaGl2Veu0VdQ+9
GqInJW1ftOio0VqBv9OSkGjnB+W6n4LF7WcbJybQNh/yKucF27Dx137p7F/BqDfpX2yFQt830PJm
dwV2UFxqpr7Nd85hMf1JLqMWCIYMHS5sTVYrxWjI0lHH+Kl/Gl3zWTSOJihxwNSPIzkftp/42zJ9
ADX5A2b2RgsXx+iEFnMWSc3NHN61aGgDf+RFuTEGtBnANkAXZnd1piqsbXMgyMAo/Ax+Fneeil+/
E+yXVZu2bdYb6jRp+26evPtLnHhF9X80t/Nnae9qA/b8xUCducBDtRXMYT91o/DvBvIdqa8RqqRT
SejnbMZxP6VO6k5/xxHyFfzJHCrkWY+OoeL/MYyojiNjWvDpqkzQaHDqQL36Ww0QZFXiyhj4g7t1
tLnKw1f0FuwsUYuUVZaLsAUNs2yUDx5xGmtqUq2xzIobkMYfOKw90q7Xjm8oZY2Vy9r580ziWYZz
1KIMmSMnXlSr1G8nTmk4ZZE8hjL5o3lIdzdFyhxjZAOpSwQD9+P0edkhWzoJakIONveOGvHNrfYE
uxdV/tM0lXPfEe0nc8RkOlS98My5bItI3uWcPj4wZnKTxsqtheKZB6dtB6RDPwutvp48HIHks1Vf
LVqKQbjJMwWjOAe7uth2b6ibE6ITHmvUjpLt8XWRlikdbC6o5R4gVqhbL3bwFv81DAfobY+771lb
sGZxHKMe2Z3WsOUzd1QyiLEgpkbCmW/AyCKUp6WuoWdYjpBwQspq7u94ID2i5pva+36/DDvirIPJ
BR4Z0k0gzDdjDWgIS1PdHsW85rIGlmqLncdspS7x2Ef0gptw8lh6yPomYYxj4NUoe3D+68ELKi9K
7AnZRroUzXsx1zl6l0j+pU3rKiaYg4+l11nVbOU15zfD2RfkU4mYAz/YQuLmrcHqwVDZhChtsBHE
sNY8AzK0TXR+GinHx1PY3pVWJpKIJYxRXfEKi1EALeYhZd/8RmKPRsWQ/W5uKGzFH4a81FOcK3i7
sBLUqOtROyIAzocRfyga0PLj11Ivj7VpH5kahPlGqzjhq5p+TuVuwcKra1zwkiGm6hVGcJJfeHMd
PZHBiiFx/T9UKQytzv+VGfBZjNOyMihCrCf9jPR7mrV7SZTGS3dw/k3VRNiJELrY5JQc0kAkwjub
pYVP3lKq8KgYRpQUjcDAOR3u+TdGHWZ2Env/aUhtNsR3lQIc19SH7vvRVS0169WgkUKysjlWYgN7
NJe1cIMHI+mop+d8Hm47PZ1mB0BTh8Ivym5ceCbUvTqYxjy7jStb3xRjJLuGr7uxR3vKqjwggIM9
eLCatmmR6ut3Hh2nbuB2w1z9M17rdhx5ZcitRO+AY2h/oGEGR0GLnVXMKDtgnIilhMPM8PsmLm+W
OxneGlZKRVMLnLKiwh/qTMsmqgiyJPDPix9C5UR9Nm9tluj5fRyL4zQd2bmn2Zg9678kTdw5xUVZ
n4SJHxgJfgMgTBSODdE4pmFQDltx/qZYshPe9DlSgIoLJ+HZ1HPiQP0IWzwZvIvC7Lflvk3kA5qs
G3GoptxXkH77X8m4/lCtcEHKz9LFF9z+EoKgSzAmfYG/u1K1kP34Z3KqXCS/L3By5cJz8HA1lLOJ
I1cmBBJfjW6uLnc163A2azRuivX7N0ZQQBdbGKBhWI8jvbcDDn6pyU2QTLqclM10P4YK2j/yVDVl
PitEyZvRni3/t0UDYniDTOHmEXnIgtxhht+pTveHgUxC/QKOLbVc9EJTsuvMe8tHKSzAnt3mwU98
Za+AAQ4FmfbafGCi+1JhAd/81hWL6Xma4OlPnIo4l2MHhwunOyrR2UgQQ1VhSrXWDXVRI/v4JQin
SqYDOjQLzM/0qQi4ciMu3G+2D8P3KeK1LL9TsazZLvtg3khiXvrUkqqV2CkT/EnwyYfxHEr2AhP7
a4JU7h0KxShx9rzrcilfnfzv0sYnXZOO4gIMaSre+8W71RSrwYnFQWJcHSv1ti3485VEvNIEo6oT
mup7FBj3EUI3lWuLVD/Ptl1mXQEWrJNjpUSu0mh+ifzUCn8QbPUKkZshFRLJPGsZ2KCfd6A/k8Cw
2wVHs1Ilb1C3j8ZgJd48BYB1DaRz+7qUyZdWK+We4CAmSaCQq2qHh1EajwPq07lL8eT4GOVxLFiD
Te4njuqph+ArIKre+F6DiCGI6Ng61M4GNCDlZJIav6om9l30ddy+5Y2E4lxVgtqhDVf0UQvCaFWp
cJxj1Y1fI5FaaZB1alo7O0fTrqLwoakMh2G2/M1+/k3qsoJ7RWWGF15xtJ1S2i34Ms4MBzJX9u6T
YQTIbcrgibiUT6zKLBmfp0U6zQ//SQANGIbmHXTiHxFCyu+Gwz+kq/FzGVT/D4IwhU6inVPWtUfI
pebe8umaYudujDHf3BG92Npvwmh6/ZRs2O7MhRWWQUVrt2eEzeS43sQTTMwkR2TW/zEZep2Pyb8f
8g6ukG3d3UW2+k6fZdiWm4Lb+4p+amPWYWv/qPcM9SJSk3qTSmhWHn6MWDrO5MPXOnFl2kuT8f7Z
vnTKEXD9ecqPxhdxBzBbvLlQBrBpS6ROEMD0nCYLtRuruBsOmVyokO5Zm9wJvHobtf+vAPJtFCJw
DDVzZ5qMK9fUu9JLuCU6bVq+PHyMSOFDWW9BtrHFMrsIWxSZ3CykAULY2TxyW1Y0zpd2kJv/L1sD
FaPA05ieEuQ7D12O4CiiplU61xvkzbNawTmU6RIvaXm97H+bdeI91zYVCgyucz9vxTI9TQWt8PYs
7WNcmIUsnYlUJavCMpC5e/iJ49XBBipw8VoPhC+GJLWX9YQ3XYekdX1i7kEI38/7U767o83zqqEr
iO5lLiL8JFiCkjUXMDimYVFjDiWLjJfvJXzOuc3kSyFw1s8PuvpjVoYBYU4pMxBnHg+SET16Duij
/lN+Ak4/lkhgBt70ICoZp0b5cQpjjcY/fSzVp2aPFXVSnbv+ugoZUZHcJH7jB0S3eJS3INOcLsth
5yXWlz3NEBvFwnBZBhV1nxkh8cAP/k+sa2J8giztZdEt/3a125cNlF/wuLVovR0SpNfnlXrnbTHD
6+iHdlXGeuRvsz7ktXV5Pg4JYR5kcR+Ow3wfeOGekO/+spMiSvFjY8T58oE9G/TocioZFPrv7upL
bux0lWm4GSjNnJWVDRMLbOnV4GkHhq+FgowGXtR+eyY7kHKA1gZDZ/y4xEauKyHoGHx0d4wDSuRI
LRjZUDeEvZTgm1sUoSlWfTD1AVjrE51mMbkoxfQLY9TMcW53jF+gTtZJtFJ2Ii+LaRYr7ygnnZPe
YdGnyWJX1emNLIEF565JDWVnO+mbe9cgynW1v9dOhjkHDh8+lKTyezoi/2uiEB7K/nDbANTFxvun
4z93p5JDWyBSp6UeLSnr3MGL0S6yPsplWuVTMvIpPISbTFb/qKo/cRzLEEonQ+rBufjMPckj8TM+
+wnun6BPst+7vHEppmloTsIXEf06h1dtWDH1VtNPB+05af1SOf8Bo4a9uKTMOhyCqUm/Y1flFoxK
tzY9AgRYFkYdfs9cCyeaAaErv7h4cUt53Wuq5wCxrbTYQYD2Zf5qD71xf6g43MEcpn6CThOR8MgG
cmmA9SxZGAaoEX5j8cSOknABiTkmd1uHf7sFLdrX+LZ9+dEZtg5t/zsPoRVTQ58orV03qIIgSNPK
9ESfJ7F5V6Pt3YC6jGew+s/TovIdxF6E5R5PPUpw6q0eh8Ye0CvEYPp45lub6Ly2+WqQYNp/Kr5u
emjz3CkChP9TIJxOWN/aS9TS2GgahTqd4mZS2bXiEmXw5NN8Ka85ZraakLZzB8Ijka+JkJpdBPgd
Jb/S8BWjTMVq2n1/4Mw13zgU+dqSWEO+Z1jeCmlC5fUoZp0BqybrCzNSHEvLzZ3AseqlECFvXCu4
tzvLayK32OPe7UzjQoenqxtT30YX9LaGvoIDbaPo4gMbo6z7NnMDzt7lBoevEyKUa20+F5mAy256
7QgxHN4ptuyl5Q8AVociQSPgMAH0eYTAOiQkWI5fkdFYf8zPX2REkMe4z2fhlLLPJzD+JJtRY2Ga
is/uRSaTQ3+GMR9YttGe2ecU9bKp98QWBlQsL4sl6AyoV4tEqtRruFzmbqhm/9rQ/AFItkTQ511e
aslTey4bPNkAh70jNQ/h7h4xg5ayyX8ghHxm+fVwE8FLGxaB5lTZTBeKRfTfh5S8IQz1Dte44cP1
2Sf4hh5FJiRnx1/BAbAriQnFG2cTmYIB8TQSxX5dQ8km/6lXSrrkfoKNPKtU546eUuBESgm6oyt6
FuPBcS2gNHbEVQmQ+F4g1/0wHmRh9UaSWt69uEq8NLqQ6MYvAy2JEh7545EZWCfT/sM+RpJiJY+B
6mNLkQ9n3iejdcT2kLTRIPZfHJGqtckWMrJhIiXsoFBMZZJb0znk+15jKHri+VbhJIYcEn4WVhMv
Zdtp+sISBqs6rN+dTY8DHxFA16MEoP5JtBQ0fVvyKdryhrXlEIOa/87zMfbqUt8T/0N9pCMxBoUC
0rLXpY8qjuwRDBq2kt/cQOVhngdSRaFWaznmEHHnq2SsVwgCW7Up23+kwjXqN9L+FwR1Lrdm7FhT
bzd4ksHLflmI7e5kjxEp44aYKMpYgBFTzI1s/dNDTxw/+lxxmRAgYVlcjm3uZ/VdPzQumtpaRNC+
T7147D8KSZsSC/UGjKZOUwJCo9dfDiI1VHVprhVtBzc7sQDVdQJE7DahoKnBb5nzGCksXlNGFJAN
TTLe4wh8wKyvYPRoxfa60XtU7tjoMzYsI3Rvy9FFBvUgFVB39LVZ55w1kaExa0IV06+JNsxMhQgk
4OKdImsGD81B+tCsCNoo/CqEo4FfVLxwbMeGqwX2K0cje0K+wmsdk0TaLsb4V356iUrmWB/2A8lj
mXnxKAnmV83s11S1bOa3rL+Fhj6w2mTPhGnE5Qoz02iV52n8hxBxx8ZgK4DSHmezgj6Mt37IfuE1
kJ1gAxeSBIP5NoSnS+TCBTfdLDVJV2bFGBnCn1tK2rz4ugB3uhtMTE8D6aSGn+DrjPZUXApy8Z4s
jsUtzA3QZ0LvbfGronOY9H0eAOJ7PKi+oJUbRksiU7kr2KmSCE9k0aDDie5/yw75e8h9JBF6ZHSz
Vh3v3FVGwFtVWLh/o0NpWkZuShSnPKjyDjNRjBic1PJwhKjQ9quVngCYtRv2e1T8TCiv97+uslJS
VY97gsfBdEWUMQ9Umyips9BhiZ1kj2IwSfiQfPJKVtJiv2FnAslp4ugKvez3k3YMAjPslry3fMhi
IgqS8y82jP/mYD4nHzFyF2B0AXjJ4oo/NT7g9tuT/k5lwb3wbMhZsS7OnqDcOqI4xqi4HoCs8IkR
AbjyzNUSXApdIh4yzvNDZ4uuByyeeSPc3efV/joBz5s3EGiaowq2fUZCPAmCpmEQR3il2pBqPYkL
iJ7a9DxZjJCXuMA6yoAoSMTTfny/Q9mOseCepFmCCZ2YUMGCZ9LTTkL47il9zPHJKdBMvrraCW/H
jxAHimUys15br0MiP1LwqctSCvK6yy8PFxnOftNa9z02sk+hQhO0Zb9sA+cP5/IghxJiZPs9NaYC
EYkLvCy8zu3y/TBDX4f+yhhzJi6PBuklOyIgLYIse0fX6pYw1ocMl5s3DDdBByDiHpF0gw/R97Hm
f+41hyONXg49tYv21W7q2FmSEATZwauSOvDlIo0EHzl6qjilNXWxjVHvKQGXccYFDE9GFGBxd+VY
gjYoSYQWlTDxVxjySaqnlJpeP9rcGdGdc9UWEEiA9ba4T7Yf5FcOZ0ZbjO7XPRsSj8YhfNBGpads
tz6Feev/QuNYzHqiz7N+b1RcI65HR3bvOjTY6yy06v5XWV5jzcEV3HSSbv6Xi/RD+mKUEFl/GAxm
7iVXIMQfgvXf3dS70hyC78LO1ozXGKOw/FnAjKh3Nqo8pK8wMDyuiu+uuQJOHF3CQQjnrcpG3q52
xIpE6uL+3h930PcwBVvgnhRvZa0fRDlI8svJpSQfmPcRBh7573GCkLx46/G6LBcT1mM76WwRvcFw
P7P3mx61RwUvttJZ6y/xdqFtzY7fvEEScpSguttg6rnA/pW24tW4zdUiJykPA4gtV3wjKxi8tDDd
439VeN6VmpUirrOlZO+6XgC3SSsvWEFsC3fuo4y4LfxvEAEWo9JzJAcN3uaWKgnmgIh3PXBiiRIA
TdEORzRKqZ4zxS60UtnvOSR1sDKlZAvkXBp0WDlC4YwMyJIrc5HBLeJeAF7SGlYlS25CoQN3EEnf
uYjiSjxU5vZ5fXucul5ZqwL2i3fYcjMdmRCPvOrywMOXCvSZ6vYdK2Jo03j+g89afU7knUk44A2s
h0JeYt3NlFjbPrEjGVpjhuCbUjSHXN31N0FvNOcv2a6sLFFaL4DpULxC9aOtTTcvtpMiqkiTKhDZ
FxxCfnebsTD+1BiKChFQwAxCaMB4Tbev92tPFdLp/KxFRxQnujygI8kv4fUxUuDj07Wk+K2xasiy
TEp7JwuLEyzWEZqX+aXLvHFZugu9v4R0azPMoU1NDF6THR0hSbdlcy3xcHLA21xEQX1jgaJ5QkUO
jv3S9YATvKD7KBezmdU7fo65RxTpdEc0PYDV/yAn2WqU6rSkAuLF2TLQrZA1kaEVvhG14gZNRPro
4Y6xVVQuaSNB2Wqd9dQvP9Awh9ZBtH+78Ul0Lc4dYsjxtL8ujYUob+Yy1+rTWRVqbmWOR6UURvFI
WNfjV8VjSGdkD7v7A7ky/dAq0gqN4zwVG+HI8ThUhXBDIa0tOAokYSzwFWcnKQYd0T8uHtXWOOjk
TyMXsx6ZdvpwPoNemML125p4Lqe6m24IuXFX6cWB5aXy5J/u8V0yg0G4bATallx/QitqcaayROZt
We/r8Ecaat2Sq2G2aj+GdPkEx57duJWf9NnxnSgsFXfulPCq42FxPV/G+FrnaK5M+QkYrxVMO8Q6
hMEPyr7voz6+q4x9+mUBYJXz34SDeBzhJaL7a7sJCtHPI9GoG0TPhKTYtZJyXQ6+mdCpdVPtQCnM
mWDFk5x/AtKSIdoI6njZumkW64OZSy/Uz2Mg7ZuaYsREhlP0mEBkS85JFBaFECHibH3bQYF9XHPL
1xP9tudc9GDtvTbJWAEfcLf6a/y/qK7+iQCi3YzD+EXHsOHnUKozMgNEXl58Xif3rhEqPXVDeDpG
pXE8yvCOmQjCO6q5C26donxJFpYwyV/z3d6TuYTlSgdqKQwjE4rBwaCOwhSl0xoeGamV2uaGSdz0
/4CVSo/C6SL4+4j9TuvWudcdXFd8BnBbfXPwjj9vN2bm1HgMEGxXy6mErGlBDXvSgaWF8HIaCZsK
8wnFABoYMcoMKKfWpUc9lpuMxDoIiw6BF8Ow08tWjqCFFPZDz+dKj92r/+BuKMa/JGRuEUwaCCti
5S5IF31iGc65dEcK9DKTZ8rDWNzkAANfldlwz7BqJojNrK6m8c9wUF7yhdV/vPvniJgoQhEntWQK
9Nb7GV5gwdnyiZ6UsfnDDoyKPE8+dUfJAVoyLKqoGAfnr8Nf9qhJAnw413pM4UieoF+/9NjPTtsI
S6WAN1WwbCZrvNYrkeOSFrnCWYFZIoQjOE2vcRS9OHETOFwBdLWEI/kuNrftYZZOSdwuFB27biM4
1t3WVQA8bFtZs2LNfuN8vpJLKLrafEHsIr/5nT2fg5z+18qwZAnEIPu7pDFiCx5LjwD9OuSBpXo7
MqprNw2fgJK3IIghDUDuBUomKXfY4i7LXirFQBBgcSfb43kiMdxLOsLohYeJiaVo0Bcr8kiNOoJt
XRQcpZ3bPUMN4m8tC283FP1OEpTFf2/rFx3npCHCwIV3BHGc1VGLHSKB5dW/zRJKdLxUZ6ANKWNw
f80lFufxAwiyNvtCQqL8rUin0DUXUT5n11s8U4ZrU6+Am42k5KCY8ELNqxTX3EfqH3NaLryO2o0/
x/9ri67avpCdJffwCyKS9VBT4afPmLRTu5NDSXEJqr+E5WhE1XcUMbqWXljqmp1BmmymhOffB8EJ
D9jh6TcXekOwIONl+Yo3CBNcswNdcfsdTdcOtBiaPHMpEifgon058RQDumv+sKps6M4r+QU8zlVP
i5fbHmv7fe+P+BsxFuzS3sIHxJ7Y2teQ79tw15IIUuslvlz8aqJprJNINLtk6jq+5dTJB9XeekNl
eu3yPekbD6/W6EYjOrYVehHreTjMbSrspNqqCnye5TWSiGUAkGnhcTN2gJbXZTb4MBCHC8C2MWAi
N0giLFinB3/IxbLvHHqrdAIzfljS2g67qumPE8ykaOK683W402qfnLkNehYfcroiZf9d52j3Y4B5
3QFCr7X+JZcVBwhgAWw5DsGL/iLpgDEQQ/5m+ZoEWuR4KbV5WP0szdKRrzXDkz6Iajnq4F3N5H8F
a1686evzFMG0LoTd64g2ReJBLvCohQHBYXOyMstdop+i21n1yMouFbX20lbE4Eqep/T3VU2bwC3G
HCLyISMGxBSRLsO9G6j0MX6mrFaoQCn2jTOCk0ARtHw4gPsC3+PNOHEKy+8rQBMf1rNGz1b4gVVX
ojr0C5FvmZkVtDF8+aBdgQf6HgT0714S03e1hvyPp7EK2XGuJCp9Ml/S2hH0zA7p6xJpozTNgXD2
q5WejMvbHzEezzk1JShg8d3+/xKCFBfAp0iF2o86ovL+NywxdMI+OKW6Rx6ac2U3nXOhMwXCHN01
HY4o3HM00L4hWPuNIvon/LtRbTFr455ZjMNfCHDlAm2mNLXIsCVRyIlmtOz3TCG+rPfkfsH9f5Fr
iJd/myElrTpLqUgDz7SXyEMruuqqBSETsGwp8+82gSxbky/iBUY6zqVM9NTiXV73AqKDMMVl1KWn
3AU82ptc1Qkbs55gtsoH8ZIiFJJM0m+9VTDXNt4ndNUj7abrgGpAO4491u9MTIOXPDfhGD0wjQko
0/cr7nK7uvElu/7dCUFPrElJ+gQcF/psfXN2McjA6uiGcAL0UsBLHA4++D88z5meDht/F1cEFmkO
7k3+t5QsSJFdpY9r7vhsoRXvWBMhYQPqFT7vTQ/DCbQjhvarJqcAufEbS6o+6Cnvj4EAzeoBNmYU
aIcmMQvjtqeR188GsjWiQwFGu2dfzrJKeYR+vm4W7fMWH68rYNRHmtngn5+pasWxK9hO/YMPi8tU
YXPSbVTDQ9Xo/wloTZnCDQL++FmH5CljrsTH4jETyZ5MgIeDGXLg5vYKCMEH4tnJ+ZdAdp78QwUG
qUhyhh3Gfn7xCs98ZFn8XfZMqcm9jjhgOPgt/dEY4w1MTjedQQnxOOBgPEc6ufIGpJu5he3rmObB
LG6nCcSH2ZGZ5NgUX/1JAx5DBWTpqZc3LhhXWgZPCkFVVk5pIvWVEVrhJnPv0dZhzxYUIGxaAD8H
nqEaQqYySYFG3RssEAo9B8bAYh+U0TEnAHnZspVr8wdLxvKlywqPANNgUutiw8FRwPu1xp+/SEZX
zfjIHiGIUIBNV5gwi4l7OudcIw9PdnCN2KbVRfnZEipJfc6tSyyfY++nNYBmicArCpON1z0tMx6t
6IuDURAv88SDgoKM/6FaOZ0la3dGyQv0v5kkip7bK8DpsfhjIo6WCjYXy5LMjAkv2OwFCdGDy/v4
pq4IoQ8RyziNgVlrc8cQpRWdzKhrD+eBlf8ws/EUPO85F+9HDZ1X71AJvNc3HTxoBYF9HYgkEnRI
qUPnpT+Zqrv1jEGlGlZTIZKbVRf/WmbcfxRNVCKZCc5riRVWjJhjLjWjMl5GpRbzaEG/r4R1tY8C
+j6rooSCwRTHHeORFgLBevcqrau35+WFZi8gTCx0uJ3EFMv1v015PAK4vhRRFECyq2L+ya8Mb1Ji
d2C3Eb7A+6Me8bkeZa2AbLWUB/Gi7V8P5FdkyFIBMIlz4x1KgpfLbjVl0T440XmvilZ5CEZWEUPA
S2nKtxsNSdOCQjUoVa/p/pQ8f8LE2nM5ZUxJ/qteaQxqe2mmghaTJNLqnTRPsyppQmNAqLCW3/NY
9kMxkFFYO2gELoI+ibA1vUZS81yHt+sPLI8A+P2FYOcd6qPVyEcyrS22ZeSgqVZmGqS/2DBwVPno
2iq7gjwnIwhQFCTWyPvBjci7Mb7GNZDaEXac7xiAm7iMHtUaNO88/h+/w5Sw7EFmTnK6mNywIDnO
kDH6hiZscL7cv/dWKXc/YsIh+8eJ3fTDJlKFYV1/NHFPeP3w7Dofqzl0GdNtASQG0oexgdDN/SXX
TlEUqCXkjfRaL9tqWQCIVGlFXzsDT1f7pO6Tki6+e+RVBt9OQQ1jz6YFAxBWSiBHRrRQfPe0zulZ
lMCu1r6GLPQJFxNf90KaENbL7clH+URTRZPN+fVNIeQnT9f1jknGX2hvHopL51WzaDsfau3/460I
R8WjLbXwyXZUTON1bmEKnbL8dl3MO4GyM1yJ6ULXtr+UM9/H61IeeuDgCmTEjCNXw3ujcU4jAaJS
/jnqTF0dDUGwCYX3Ab/LogJQKMvGwyFci6OTLI7mGSNqpq1hBlpihhzz6wHsW+GOF5aQIioafuqZ
S4dEbtm/7ztxshr0HpNGDpOnzVwnLe3F2lsHLEKF606mo41Srarz467UY9/DM+/p0TKYwl7oTMRc
iX3hVRiVs3Ir2nQnAeWg+YpW7yowYkw3NuHOlaVRCPaD+qd84VVCC62Rq7a7f2tnrC5HwQM4A1VC
16TVEJkcuWk1Mo86VLRq6CxcsiW5iTpsrFv14ZWPYVUknu3OP6mrB1hz6IjUe0+siFtsQD8wy0z6
JtfFgAQCPnvOVjapAvf7LrviIS1ctRlxdg6EdpxyHpIMPfNPq/YlCuxyAOyHSg2t6zn1w+rnBqy1
vZanZS0A2eh1uC76i+SSkMuvule52lajExV9KudTHrwr76eaw8Cig0CjkOJ1wIo2bQhotf4UrDOC
5aLSHpB7/MqVzwt2auWpNUNUeHFuV0mo/4e0xXxPWyeh/45xN/Mc9DEC7+A7UpTiwJlgQ5zdSpZ6
AT8utuJeyyCoTsepjifZ3bwecMXGhAhGeri9t/et8bUyOo+XZNYi1JBI/hj8cOYBdpAft7SjBtlF
jMcOuCNTZ7SjDyGPIZ63ddmF/f7NzXHPfWNO/AmGO8Qkb/Obarp2QeqknndCbqqxGewWul8uY7y5
1oZFNPOpONMW8x2JsJmrIjd5Jeop/oYTuPdERu7dJHGmfGNv9sy4zMzL7wrE1EFW34CrHFqtlr3T
XlCrgYLAQAVrCZKnKapQrmQOMDYjuj03SHQwGsBer36NdL+Mepx5WRE6pty8rWvaUjbCarV/s8Pt
Cp0dFjWCuVw65E+ppdHK5/pLh5bQJdviYVHwVbHJcd0vB89Yw7wWKOTNYFVm8VLk+/k7GZiQS92c
3dq/o4tqt2TtLwQbglFn886UiKr8zybIz7BHldPo0XN/DJUq0GwjztXxDtZzfgJEOXf4YNzicWL6
UYr4bL/nFC1q8ScrvjlCRLDRFh5c0Gw4FAoXhudmmRXUQGj3+ZxtPK3zWBETxHzN/HVnOU1YNuv5
NnIFUTHs43/GPuTk8xPf1BLQynA9BhIzsnJn2C936Uzz0y7BCNEzUOjkIefqzcsBp9RkplBINcR5
W3sIGBAqQz+EOWiHmgaESvwM0GNAn50j82uh+ljfPcb+s0J9p7EjlQAEFGyv5G0ggSYtP4I5hDlH
5dRKgKncSukSNUlqaVJh2C4tzrMBbmEv89ZnGLZSM5YkVfCxmVU1Yp8bJ1y4lHk+1ym0+lsqC3Dz
eNEjO/qBQuSNuUyZLH3z0Or/rBhnsz7+GquCCajAswYXV1iQY4Zax4Arat9vNiGMeYEqmN+sb49h
PDe3XbIbmMlEk2w/vU7OcRwjkABAIcCA0faK8UWRIBC4CKrtmaYrlRiecr5Qh/b8MmAh936JHI/j
rlx+v5HKs74XX0WqmiFUTwKE9h+ZdKurpPUc79UHcMerU6vNiPneSxVB6VRYdD5Cork1cRimF5ir
aO4h9BPYv7qQU39IBDXp0caCKHkTzQDkjgGAhf5hE2Tjy5MwgcJRoMVZhyxAuTldpZhOTQ2H/kjg
laiSM09xJ6hJjZn3zcsiW2EyXuWJ0SFu9iGBOK2+vWL86vlrP+Kh+FIRioU/UVb/KEOQQ/3bzBd0
NBORF3KNMeJ5F9r0uEdhMy39OmkUBRdS76s/rgGXZ1gZxjHkfv9goJbAaSbstfkL1WkSQ/9NQz+o
XR+IrewG1A39qkXlnRqITvLI3AWe3gAUSOZZQC0HLaK2XikKSQT3luIUFvlhXSMezhB/IzkmP38v
DVy1bt2136Xe+qXZaKLPGzOMK5lvl7+cxyoCTF/51cJoGKyt992T2rVVEW9CCPpWD54+vnfZ0GHh
bwG+fDnha5k6cZ2HnNYeQgJurKrURBoO9plepPZRO+jBpdlpAw5RoK+/9JjSQWjC0dJf693EtF8w
xatEpMCE50dPjTozLLyzqWQBtYJrYLtb0CNT1NykVJQFzqIz/FGBSP24LTBtzuTZ8fGyEBq/OxVb
UJSf6h8vMIE1YCeY6wTAE9mJ7dvrCsPjjm8rr9omC6TctK/12rLJQpNd0glxqifu8phbTjP58FfM
hybl1r/HS70jF2SOD7VJX+5RpsOzMVSIHqquHalKgDyg0knuxYZlA6LHsoKYQKxjbWM7Ezc3Knrm
/pt3kRCqeufVifxyPqA5oUfKJ+l2FR2PiKWqCmBRXXgXPvxbsSxqhbWNfhBcDsDP+vz33iNiNqob
fgAbCSdA/1is00aunksc9iu5MaoWnDMMYo7JqGDDyCC/NXYJrNpBjjl+f1ALTaLrxw3apRMhoP4O
DRMerm1phCIjt9ao6anRHGJuXuGQ6kHRxtVRBVdg/HKhfz7xiMpQqM9u1EAUj6NE3/XtJMF7p7ap
2Mt+M5+Eg/Wk53DaCrwDsljqMmicGZz5tDAbTy6hCvymDN80NLWSTjIQMpFOIdYq0nfRrs24xdgz
a3nBbKZsib8NZGii64oL9C02MUfcF4LGpRkYwJQ0ibzsElgvKwQkITOO5KtmbPNNDmcG9HutrJIT
j0beSRpEvJUwl/EbRylSXj7F/Nho/0S+xbXRs6Kd37uCND/OeFa3znkfTdcsMQXegd6uCRsvVlkb
WGzBG94AO0YyiEt3RigJ2cPrmHHBQO+BxtDtcxGNRestpJEkUhy8KZShjR13nvKnAT7HsIK8fYXf
WNvHdfL4h52CACyI7KGZCFLY2YXagOhLEMgPO5qEeLXYJHOGMAPa7TK7O1HYXlwCk77PNkKN+Nof
t/rRRo+v4S5aLxpsvnxecqRbVPQ/E483zwML2Vjcl/YVqdI9nauxApbH8oioSuzHMq+qGOnzC/Dj
Ga1ehXDDZh54qoyqRulQ9yGJwnHMjVcKw8aSQ/TVFo5OquMpsDBRflM/RKmsXoqy6h6WJK0S4it2
kL2Z7YysMjWT/nwA06CDr8KcZ28NLkIzN3rRZBvo9eMvZspQkvKd0dd5Yx9X5mZgAZ63uHsMNrQZ
Nt8IBgKA1Zrg2nvsKAM352nGkDer7r1QOSZ3Tcd9ThHvw6GXWeJ2+yIuZeQ3UOVsERWyTwaVMsPF
avZ1mHRs+TEQsOfeddrGWanUmh/oE3+Hr64kEHJXIbFbX666cGA6EdBBJkTc5OjbgjF0mg0F+U9K
s5rinxnJo3rDzTo+fhdNS0leNvMrm+ehltrKWzGkwlZU28o/R3XVpq+5KaPblfqaOhZJ8z+XDn+H
mzTvlZCEc78S9olJbf+0jhuWE9Ul3kkUoXb7puMocUB/moIW2dBVHuJ+OTT7XClAiQbXX0U5Qe7e
ijrbtGK4laL8LUhFtFzwzPOnn4CORCfaNzlOdcDS80q8gFRlYDSRUfjOv10JJJOR6NB2ZjwekkQW
wl1qrO5fZRJdqQD6qaWAevW3GGQzX6KMWQUEzwPrLO+kYgAAMZwSDSm+J40Mu/6sp8wEDdBz7nGA
d2VvjJlPDVCH/mLKcjDgJjreAH60fwgqPcf6ga/7QSXJCgWNKN6QGvifSnh+ei2Yvc5qY75egwhZ
KzO+WXIbyDErWK1nxUwup8Lx1dm8202R11vhnwLCWv22oZODrmOE3rNuIG2ldJbNIIP4+bA0YGXt
iQ+MPqFoEwN7qPCQYy248+M+hiJ3HzsTYaSgczRpYRw8MzzPs3mzVpOtUdJt4rDbw0gT1TO8T1FW
0KsKWINHEqRqcS3FnfQsb6ygikfrY4FU+DRz4Gqo0bkWQBYvbWnIdyHtwogI77lWrusEdURfTzz5
Io+paJ87166OpfI2lWNJj7Jl9jDIp05pVboMD7AentlaqSY/MDUQhxt0WJLACNJFvAZNixIipIt4
8lyzWnHg4TTHiB29FXs14dZ9YmZh5pda+foCKPfLYWhjC67THUHD+nRQmcDMNKLP1a9WkFcE1RXQ
GM5e9gq6GBirCdPlyjDaNTXMY5VDPb3UDbX47fyOBz0pX5v8RvLxWtghSCKidUj2eWKYvYEgbjtO
QfJQKxJoJiItifMRtNPLL/zqGEhsiM2TB2PRpdcAYPxFqU3rrG9SbGyMJZLjFTDL3a5jZf+Z1u9u
pfOTWrRAC1XKI/2/cf9x/q6BuPaAA4/K3qUfeTRbJQ5tbmjbcO0+32CSamM4snpyngbFdJz6FIFf
Qd99fl3P0E+wE9LokwQjkt+mzZt7eIorH5Xndp4OHr4CmSqBE+x06jWd4hzamnmJ3oFaMcwWZy2Z
fN2LpdXH1uH+a6VEBQ36ctz3IFsgudyDCjEOA/f7NLXAQjj3q/AATWhJGYjGUAM1pIn9JV0fbdRj
5MYotTKQsamFEzjD4t7m2uljFF1wZiyoH4YJciua7NUxmukVFIYSE4A51HKCLHmcz1cDzg4Bxcl7
eAcWjOgyc1DTSOvZ6zM1ExvkfDFUFmcAeevRQugC9s4I7U9tmOPV8rhiE1s8cx5L+kA788VcpiCI
GauZvBif2Z4rHe3tkTaYLBR3mCT2+lEHgSz+YEp+UoiOtQXaYFI6SjEgkUk3anBaPQO5oqlLh+lC
FJuYFHaf81cjnzwhj+SFXfwtc4BGES4DYjwVRSluT+egegAYxfDCxGdCRwgnuXHDO/VmGsZfyimU
WSo+1RcpdZs6+vnnY9coWb71Mf3bHpxJoJSoVzb4rWszfhVuJC9sfpDUZ3NfmGJlUubxuZkLCTdR
hvdNnnWvx31R+yEdsBTDUgEHJXF2616dVrWMMeNCDUnVtjRxWsQ0uIigKkeUvFT2pvohPv5mReW8
3RHbwCnwjQkJuMR7OYrLf9zedUMdf1SKQ4Ovge+gcLC55yXmfJ5Cj3x0Z+pXpE9+YQVeeUiu6NPo
jcikxDjA/MO9Tjk5w5X5DpFz6epG58T2HLS23qYuIIIeq426R25wbWB5sBikDezPCipOrD63VoAL
tStM8SwDhp5ZL5f7WrmV+LUqzSSjAz1jTzxemjeNMtoT+5dbl2xFu1dVpJwLpGnKx9DreoTy91BF
uW9jv7l+Xt9eISQlPH4fwPMgrqsT+l8b0zkHKtj1bA8nN7dVXabcANBx4bMElJedy9W5xBi+/Wgz
3uEpz4BfOC5qQ3deG0MuhaFbkzoTAgCn6Q3FhyzqjV55xMFtKQ0fNUUbhBRSoGzaVECpwpPex4nH
yoMb6oP2dxz6Jn6ZW886H6xtlTyT2P+1pUhCf/M+n+sNT7+A2pq40Xr57oENvVqqeomAKJ0c9TOs
9XdcdjvFVUDUxS4QlPprxN+VqPI728Ofu+6IkXw05AsFrm6szQAjup5mFJFANIGH9UGP4aaNFGur
b0VVyNS0SGcTJK5L4z8yI8+5uevRSF9obe3xIfOEunf+Ker7PypM/ddO0h+AjWsAhO9ufPAVjEJi
SexsPRaHtQAplFeiahTXDcAUD33/lrm8pDBES4xpUO8rXX3VdXJ0sE0Tzd6BdwtZawJXTx/wgQ94
ZOscduMLGJ9YWPYtt94LkYVkh0X4VuGYXcZ/MrwkZzNIXAmoOO8OnAumZD59c0rQxUi+AxhS8j1F
iTFs4dHOQNB6xxh3w70rMRb8Xb04y2ebgHK3TIiHuJFO2L/juiIffJ+AcXx8VguJ5lbSuoC19u25
WiFp8f4Syh043oJhY2AyeKGdoyroAaTSVKCpjPDm83dVmVjMl03GxazjkUEG2vBjO36TAM8EQSlY
WPTOH86umAMVDJXSw0HvMHyfXkQEoSDSUImccwgP5FVIJ33R0TuvmMJCsk8fOxXoKcHRkTYV3hSl
w1T4wxrDVCYoKG7R/dROCAI1Xy7nCaaQm3O2BZLyWA4I0uZNIvB44JCWoRp8VS+epbwJchCqHNGV
kIjiYOz2L/cG1BZ/hU+tO1xc/revVjeqy9t0gEXwmofx6uQCLzAy+UCFgobo+0oES3xxo77m/J5S
wCBtJLPac+gD8w1HpS9mGA5qqZUmeH7W9SamzGkkMTWYvNvXt8ym15ahHGoDh+KinrVVrLSacKCY
T4n9Jsd9lZI8nz0TRpHfwioRZ26OfVGWRk6cgVzjZ2WcCkScrbqfIVMHkI9RSXf/HkQFxG2ZL5wP
MDAzx3QCvT1upsNUI+C6d6n/wKLgEpzVN0M4KQeYiDuev2NhoDrQNDFwVcjcKPfnS+2frwtYgCUg
WAWMiY+FnUlzAcNF2Ql5spSzGF2kcS6YmU+MFGeLYtfrav7+5MfF9EpuKpy7jsRo1c/qYB7L7yU6
4vzJMqzDxfpbqAFTM93jtjioFIGkkxa6hGILPnZUZ+UJhG6p4ttCzSSUHN5sJrmXcCBp6xs8NDV3
eUIm8Ecrz3+nhr74IrDYjBgJ2CoZYWz3HwpjkOmPwEPO0h0DDH3Jyv2qEDvecxgCO8Pc46pBZBOS
jmC4i7V7Znrw7HKLNe9dcM6qPfUqOV+aZYvF4Ypy52RwDaS2vTuk5r0HhJ+CyCH+ncP5TacuZ/BB
8EW0pzSJ7woS8JBwHt5FIk5oyrHF18ogElehpBuYptHGtJEVNyq1Gvmz7tEY73OB7jLzPfTT1pNc
hNHvmM/VrIRrbjGLr2BeZ2R9lz/6KnBzMW41XC/qhVzb76QSJiJYYnlV6Abd+ml93tYMeJ4qco6W
hA0GkhHPyHR4VqBqu50u6V2iTBj8tinWlqPKyElIKjmD7YdXKGDNLOtUdRDMxy5pS+L3X+Vm0jz9
A0VmTkGEHKm4BaptNTXaGo/OGnRNSLiDJAN8pgFURhI18CttDhAgpeBC9dQ8+DRoMDNvdMou2vN2
dk0iGlnUXHuFi3aqbwjTCLqC97uZYO/BKYXapLyqP1Q+3ceOoEltjMhYDArKZOJoL7OzUGsXQIbH
yDnHEjruapjBL/tJDXY9H3idRe9Rd4EpoEIL10LShsKApvK76G9FdPiZKEOL4tAak88iQbdc9Flm
LcFuCY5jq8CDvf59Jm7KO4LuvU7QjIcA1uCx11hlmgcl/W3Hi0wmxnhAN0tufG8AQXciGzLPazgU
cieCJuJ96I0Rws1hiAVzpgRQ6pcpGVhFGkcx+v+HIq6biYarNMQ8CvZJsOqQB7L7L57ruiUX2gFt
eGzj8c5sbTzbwQMJuK3T75wb/iL4+vCFPpCDnSJ7chF7BiRKJ3m0oe1zmqG7NCaBAPKaOadU0cEi
ST8MMxyo1D4XWaN7jRyAGP+YymNzApvkN962k/ohyBd53mQWrv99DJQMcNh4Y6dA8kFS5bH2Ugyl
MoniwmYbDMNWA/8F13eXr0WFDnaYrY1q+AUVyYVj+sBc5eUjY+yOxdvmZGklpCh/6OQauLaeDVBl
Sa0LWELtrQL2pz5Qj+cKBfKJCKN17LfvjhsMli2boVg9D6uXDFjZC+GfiQHpjG2WwCGfpwXP7pI/
PniLv0Jg9ANu/HhdHVg5UccPUt1X+TUyAMUkVlu39wOqT8nDnMkkrM/SEzuBZ1Luify3rZdM6dBG
OSm2m0t01LwWtoXVNSAVwitQsaZn/wnePW9jNyHGL/56wTFH48VVxsDC24gSNDqF0XUJVFFfB+bM
XzrNYUPBzOGMDFfAn9Jz1UrLtdxryHZOsKF9Cnij5MUOkods5BWqpyKcpIkGpTkeUDp08981GvZa
f/xQEKEXDsiz4fxpEO/dH/TBZrX14g55rRE50LQeTJ/B/A9UJ5iE5yVgqGwBEaqEbiX9h1XASoMD
OxsVSqA2wjMFkXsDg9D5Pcjhz5B9Qmw5YE8fUcTnQUWEZ6j6HiKFzn9zOkZDYSItGrXaV6WKvVjo
MZZDOCNcxIGBeOIWDBL+YEMlya0dGZxyB3rd3PB85DIbFW890vx0zbZ7XFZU/CMkP0OIgINgJZyE
xStALIbiau0KlYcmjc2f+KH1cxbTARX6eb4Z5yu8eM2PhIzoyRE+kn1rdij0H6NZ4rEVU+12Wt48
Xb2l//njC1xT+yh4j6yj9PXAiO06bGcgHNdWS+VovINaFgCudO8aZ6nJGs9FzuRf3fSCayeExeTv
6mno5kYPp0sYs7NH0Yov71vLF3vOwYL5PuafQHIwLsNQOPyp2h5KLUeoRXku1/EpVIMK24UuOii5
z1PaG/L3a9Uxkm+A7RkhFMQ0oxGvHEN2w6VYOkBE4fLOHMHX8llO+EaVgUFgUT73pY1LbZ2z7O5r
Ns1byR3tJ8iasghwj/vPgQT6MN6JKEjAwhbfslXVt17ARj/bXyv29HG++9P6wenAbKGFG9R2fP2V
rV0ANRde1tzSbLY0VYPP0TMvtFMldmjfgdEtdT+R0VfsK/l1x+juCENx6pkHDe2I6jnE4jco+172
RAPY8QxBLCK6ZVVv0YfLoQCjcdl1Tf8erwkmHw+XOadRJqmLHu3j+ayn70N+17eHBbJ7OD11Zbg/
6eik1ffnt5labkI7R/UxwwPxpWLUHV6VbRhnnxNzge0y7VKFHjcCelOyRSd57s+T8lp7W9ld6j6T
Q7xU/Sr1quqqkUfPx2rzDLiZJ0FwBgQPUbjcIhWD7bjFc01LPqecsXJsU2VG5WlLJeGbig0WoJKn
XZ5gtwbAJwCVl3n42LEt3e+5KfxN9KPMcsfnGXrYggF+4E4MultMH4y55ooWBhVVXnAhWEnx9BCS
slXzVxC/PFCQZksLWqJAD1pGnBzsSvt7wmYGjvLlma5WSBXih9aQahZmvWy3C2CXmXflFad1Swkl
BiF7aSJ+UJarxRQvWHATDgLM/YQy/rBV801Pg4UfBhP4bNHIzjKl+Id4akcP02MAXyq7T8RQSVQw
cUn7RofSGNGV0FQ4XkYLeIhKNgK1o8ftkFZRHU3O2g1AdlhkFEbswwZk/ugIjfFBeeUXEh9uYooX
DyEL5nSCjnXlSBjT3p8TSqzmohfi8CRt7uIpNWRlJNZ+Ezy29x0vTzcsdJT2CuJksFyQPttcyHMk
H7K2n0m9byaOsGF4hqFf18R7Hu3+u27zpOPzUaMH35uBbBMHU/iNY1o/ZXySHXVtTHHr58021Cfq
T2Xf3zVA7w18JYf1QF16fEc30mguIINTXVp3YMhP6t6N+Zj3+BNiL9CCTRvgWdh5rRwglw4VXPun
wZEYmNnI0lx588mXeWY0vprB5mLuOyhn2XYqtdHLry45iB4gbrF8io337lu1sQNQDFWct36QZXSH
DZhvdHQgWgTvM2d14fcu/doXJM1NzTIDTWbVFDM82EL8xgSD0y3znV8GOMHL2zaGnQAajSU5wYMQ
Ca6Jc3YIOzh7A5mTM8pMZvBcfnmlM6oaKyqoRPW9E0V9NuVHAVxwDqeObRYFgHodPqabKj1QhHD0
anlaMvIqs7vFFzJ0imG5tlWtwPNy/PAVCGj5wPwRb9Uv4Cv9FRRldgnDQYAr+vFfSV0VUgRSYGSj
6sI9l1lrBUcb1uyrCgYVp48LOfr2YsYPnVwcdoY5oI5DZ7YpIUo4PsDjwMaoqVt2bMJ+B46e567O
N9d4uxUFMs119O/rtQYGfefiempUzirrZirHgQAfs8eJSAgKCrLR0MvTNJg3akCG/cTPXlx0Mpdb
bTXvXEcoZXikneVCrsofSRiQSYebg5L2Mpj3IMGRi3eLVHzcy/12T2LISTPLprwACmqS8YUBZS+9
IGxV2NdZuvsenIoR0LHl7WUTU9Ps4Ds5K3LVCHioK7UuKZnlmapn2PFlGRwzEWByBor9knTLGHBN
SFplSqffQCIVXiRCAfU0Lv1SgjN62AnjiaSXwc2LLHcCjVHt0QzEvWNgYyq1f1h7xERQlZBU8/o7
3g6/rFwkoj6YHu78yjly+/wBz4SVnP6DFu4DxcxHdL+d5iR+WHmqo3m6xIivrNTA1UBhYe5CpA6m
LGJt+55zbuZrgj1PjwODrSynS1uNawGKD8t/VZYOZz+a354iXCWKwdIu0IfrJ/8NiRlBPK0Q+gOb
EPgEaDK04XKddTkM3J/A1L2haCmERVnZhOa9yKif9fm59SVilQG0HjmMTdlpCpHNOwgjlzN/D/uK
iqFKt0xlBesV1BYfow137RBXsP6/f6MmLIaTInjzIt4Fm8jGJeODKR3747SZe9uy5wrX+2YM4BpI
SajHvSaJqYl+6oQqy6gfRCcd07zWdfuLpva2pwXJH8Vmpxig+TK/Cfh0ewr+gTqOBM0rjSN5uMOr
s5P0bIum7diRDO2m55dYKxT3fq/COMn0OIyeO0VYypptcwK3+94qIhh9hjFdgM1UsaruyAZ8apb2
Crt+TV9DpPWbnu91PSJFjTE5vtpD8LGzOO9DmScSiz8iRh/B8B4Exl5DT3ZJISZGKF9edIHfn7BS
BvDF30xmjQOgTefkKHcesT66d3lCKZRvHcW1pAkRYucmPQDUXdKi45A/7nMxcb+/N9i7bSI3dpv8
+E7WxZ08Rx5mVC3D3hYxS/lf/n9T1PmP9PQBYwKWcGv+J23DoKMB+MRi0oxaImRXEO2Bcrv0P0r1
lw69w1Q4eSyNNpYiwJYWkonHhj3vhmPSbDlRGb6fDqMlH9uqYCZP2qA3hEgLO3Hno2pIljzJK2xn
iuywKgEZdWrHE8lP4zUveAtWbEEi0MRlmwK/jGLmWrfS8uN9LEGwIq1DjlmXeyLXCx8e5Mc7KBpD
h9zDUyfu5hbiTYXUw0mrjGmjgSD8xAwoBYhC7SZrchtJblGajTO/lFlYYpCrCNKVT2VY8Cm+Cx0l
tw4TqgHGw8ATSXvEPJjnnPBGWAGajvr6H6nlwZDWY307j7mXmPB2jdMnli2Pw79N9VRHJfX5Qc2X
nereiY4ERoxanB/7e9dfeIyxAPR319D9Ag+77cPg7kqa3efeH38q9g5ItQOOy4DXPn/7+8UjYFBF
v30Jmv4qCH8NtpdlJzPdPyr8Pbi8xQ/eKvjY/0uH8hdSLAKQ01Baq2XXgDfHrVupQuDl5dsmEAFR
Jgqi+i074C7DmXJpnT4qkaWRFs6/uJ+zKxZloj3rlohhXmyRwyLY+Bu5sh1ah4xhXUuNMJnfktxu
bpIb4rYt2o1PM6G5zuLENa6OBE22Q7Zb2CEneT/ECJcpPIni0qQi7C12IJbtGXrO0PFR5+23BV89
YdwTV7uczMzRjKM8+Pu9cghPN5VbSO4T+sunlW7ANGdL7jQJt64OABP/d6kdJ0gf3a4QQN2kXzqw
NB8s72SwBAduZdZtjol0h/lIb5R2juBgKRN8wrDmCwrJwcY6xkSn77CTNDE/vT9HlDjp85kxnsnU
MIeRbxQGboQZ/zmoX7cG5LYx9QY8vdwcNXsb4KHUJPEAlOZ+WzSNOym8e189S4m+UfhNyGPQG7uF
UVnUZQCDAoKAXTD3+/Jc4Fn3mshYZTjz2vl+q579wUBy9Bze1Olt6TNEwLnvXCSXstTAiskiI1lH
H9Wf+RvcHN8q6w/ZS66TAz5bt25N5tjuhhWPjCKVm69oBHHrWeLfy+IU/oYWDWHsHqWb8SCK/85n
f+8fPOzq61j3K78707yVgB54wxIR/RnVML+m7mmm20/1W8LttY7YRCCibfg3QFUYtQbX8VnmkYpz
Chd/ZpmtNnwjsKiBeRRyn6707CLu55G7cS6dQETdQn0MyIckPYZAu4WfgblvzM5w0TWtgHEu4sO3
yvO895PqDBKb/wSVUK+3nbYuBtfCaqS9pfaFuQGdSSLKfqfll/QqJNZWFuGqqT/QhxK6yBzzt0Z9
/1WAo+lz4GqiX3QdfFMazI5kpq1k+BLC7n0A0s4mWASG7rEnAWbUBXVyRL4+MpguWDg4cQrP8Y/9
wSrrQJXFZ1RlT39J8fy2PkzdWmKrRwkK6gP9g3kmtSj9pFfYvsZ3rG1oaCqa7Yr/hOaL4VAiXOle
yczcwdiT/Y9KuiQ6IHUxXYjef32P5mJPjnF+2rlbsYUQxSFgKV615JZbmwNt2gTt69xHYLf4keDO
jbpMkbVIl9GNIYWG//18j+nE+aeyR+GKeQ+f+ueYUtBWU33w5Q/mIKJSlDAc2ultlsVbt8w1SGvX
QqKdN3jX0ASbigO4kyxsnKW7zdfK13I5sMUkTjSqqEbrBvkXM+exUMtS/bNwaSOeicCN0tSN0p/1
+6CmSYJ3kUcLLBdWJo8L6OB4C0Ykb7pzg+1n+BSvPm8cCvkkBaTvg50FGT4o63mujzaQX+NZhUnB
bWr0KM306LRIHRwfSC+nvkgiSOLW5VG4baOQ4tGz/0ajpPZJw1abhtY/TjoHH2IlEJjhyaOcoBc0
8xSoKwm45ZwgKd9Ke3209qQH2LTnn29Roj4GKVZ3VXQ5lURc2ypPnebfm8JorV9J6j7a3Di2craG
OIbCQfDsCE2Wtpbt/k/dqojxRorw7mpNIrB5HELM2uUDK4zQzGaFA9UVZ62XvZnPem+ds2HlMfoz
cPbh47siCdFnhBRSTEu5aXlhlsARxveOO1sYwfu9Qq4xTF6pz0VNJhQ3BbrwNWDQD0Oi6jHmZqQj
mKImb+L5R1gG0cJZaHe8IAdFJN+Dq0ako9CsScW/NmH0IvotHAfu+dIP39eo7vgeJBE3oqonsRSz
zLPtcO16HtJLAEBAGf617lY3aS5eRLUsRN9S3PM9OhTNaTxD6mXoHWTUlc2xeHgSYKHWZrPPTkJV
kZ9YMLpneSgJJ7kQltNZNxiSPDUFRTjcV8AwaFOdYSIJ8AWOVxVZPbQZ99m1xAk=
`pragma protect end_protected
