// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
MVy1LlfBwsWuh5akEm9excqjw5ZWKZvqynF4PxMcBK5bjxv3q2uNK1N6wskArKJ5IgiZqx4F6kEa
SOwYNIEIth0DBeFuhqgZTnAyB38cjrtDJJqkNITP3L7VMNHUaYDFj/KYHY5QFbHNnHaic4Kqikjx
PKZEMqQJYp+ivfP9ctTh+PV0IhbbjLJZnqCNtq79OUVREPLZrNSEzNgHU0GREBYUNm+/J7s5ozBp
S8Y0HBRccz/WHNrdeb6QY5CHThUL3edfDSKpr/nR/7NuRuaj9KV2xEuG5pVRkm80APk4L6pbopiZ
1/vWnirKpNt7ngsQiLBT/QxxUAhhdVekXFrevQ==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
cXY+D/ckP/yNOorhAhK0FmF66iaEjQJOMe5J2FDqxxpiNFrjtP2tqwhzzh2ch/yWxvTAPMIMZovx
GHGU1x0oLZA3mMXifHxxt1vk9MYNn1M+NzupWKsVW8r/ErzpTkvBw9PzMoo1MBNyNZvL/1w1dg0p
X+puDLn3m09eRM/38CrzVhQsqlT+pliDePFuaVvlL4wqAEUIMinUhw2w2NmnNF6n6rnYiuR9THuS
k5DM868sSrpN12SOX7fFuCyoRT3NiZapyj8VmozkMaK5OH1haOMM9Cam8gOJgHU14CG+AT1Wyba5
IeRcIJap33uW0S8buFE7MGx/LjCLy+tbwN2B7EpSaKitP6glKqtRWIc9fTIFNB+4Xx+pwqCHRtH2
X55K53bxIGunEDj9blVGyG87hEnTTcsemyVGPrXHpJc0UknjYwtEb+BkbYEglaP40Gifu6nJ2+am
qwtfGEeBmWH74N9w6jPVyJ9L60PrHFQop7oEG656PCB4G5lwLL/SOyYh3xDoJRw2zcGneL9H8bXy
rBaExRJWSMQMzwIqDwXeQ+VEGIDTKStAEKNVqsaN9nt3lxlD67iq8PIYV6Uq9+x0jhzLXlLblSI6
QMhzA/ubNPIeu3JcXR88ayeCtrsQ2HKo0rrliyQql/F4pLyqvKVumbckJy9W04vhV9SbgFB9vHCg
YTYD8Hr/CV7GF5BUHIq2yExflKuu8c++OyBZ+DOc+HB6MHsPf+wUJKzqEhJPB/bVt2tuqQLD1HVj
a15W88VMk06FSdUVNO5PcKI1OgrOjxxZliekprQQe3CRJXniem0xv5wSh1vK4lRGKC/UrSq6M4Zm
6qeHAZx5IntLz9bW2Z4/CRb/ciy0kpDOC+6h/OO2qmwFgybjBT2JaTLNYiQRkSpaZYJ3ucS6fdRH
HQ1v5SEmyTbEWgEgAF4IEaDBFQb3PVwgTImbhOexchSeYVbmsGsDLJ7cfiFQmexVzJO8ZhIUIxWA
ODAR4ZGXmuPcHfH+53mr43/xbMCjxD07FdDhQ/Zi53k5qFwBUu8QGJYtw9OweHT7+ztAt/fBrVul
W2zR4+NkEd7zn4Cn5AkqPEUeIhilgPpd86CwedyFqb7Qv7xCUwk7bt+XA/yXp3ae2ULLUwm1/QyZ
Qb+eWk37896dSCv4S8CEDZBua/45F7uEiP3IMjRUtvgRLqQnBkvxskLtauzJG8HRMxlX3bmGQ+b5
wXQptkoQTDee71/uR8sw5DIp2379QXrkV0ZTLUBDc3F8AFZ5JdLzYHftKxTM7dgzvUuZktLkAohF
CJvC2laQadjNypmqY9U6mHIJYNiVxKzKxy+y4ZJOdBEjsHBbH9NT/EqOKj1t28yEDAYdLK8RT6CF
+0g8PJCgDaTA9mYiBsguFM29tDWxeHJMPgVyIBYbucHlZ8RlwvaTERHUzZFNuVCPkiYvrC1BB3G8
GAtMJg2ncxFZ9lMqjpStAI16Jv5o0VM1N83vjJvJv2ncOSLPUTZANsPE+GciK/0U/7OJqZDX+8Xg
vPmEX5DReQSLwc5QvSQB57jOYX8YPHxpL40zYRwPlNmRyI8haTB2UIY5AUGrPjsk09RoGTnfg5ry
AJEbYjb/T0VwB9iITVDdhMm1Qvzm7VShH8XWYhZeZ/EsXGEUxQWcy3wjtGDPQrJ7/L+uqYmc1U8B
d9HzvuzDXmSZ2Cf3tgQhnxrHmzkbZnSrx7/TT7moOgc/xkFWtIm+pzeGEEV+f/M6QwroRPV0yBlU
ErXPuzBw6m0WlHSSvrgH44OcV3deWL/QfmubM42xDsoe1rPT3yqsKerYodxPVZBWNWdQ035t3KLP
5LfKGj3HgXsLHCqTbPRyNJkJq0EctlpJCkre5OyWsXVYh/LIQvm44I8NuCp3YvDEFkvIucsDLndq
xK6yS7ZJo3y11ZNHbSVZw/LAnPk9bys6CZT31hhsQx1yQrPfCOe9+zE7XR4gIWQN0Gf8sDyf/0aF
OBhInUqHYHbbk69BeYTh7otceLqg+grBxJ+BV2FkfVLoARfziu7uSjm3TJmjW6ddJtVb2pQCP+oX
OOvf6PQin80Pr4+ZZDakkkTS9H2jrkeZpuovGA8lUemdkS/iPvofnOxZUaC0BwJDDaG2Gp9yeRks
ZDnn5Ld7edesNWrtNcXsJxmMo5XnAsahn9IyAa+9EhGYaZPPcmgMDRlUbnkAzP3qd1I+ry6RJRxj
RIc0TtLt5gE11ld6m8o+aeEftWF4vCuNSAe1uHk+1MqlERnbwKGNAasNmz2rtpJz060TWf5LFZL1
0TejgO1D0afIAXF209+GsqRIJlz087mKr1HjeGn/qGTyDne8K6wfo/nF+HN79KxVhNArj+PPhtKt
VfabiNRdU6aM3L4ukc+hGHOc295B2NPF0L8lpCftDwJNURXH6YaL40I2NG5wvtQ2Mo++Kpw8XxjU
xcgvIwj2+QgDWBAo8urHmffzVnXOr5mn98wUA2+H4i1aNUqrVazHRDM82+kslfthBOn7ahGJcqGO
vBembe9SWJDdAktzXinfzbvAlwCutuBITUskOVlkH8vypxkTYfKa7XUC8qI2wGxpjnsCr502WDEX
upULDat5Nrh9y5iq4KynFn2Ksr39u5L8jcCnAwjiaq/CYoRg0JbPhblOEWYVQS1rOW2bw1KZP4a7
PiMuGJERZpLsI+bCsLKBay42MhIiAoN1zNSJaQVVg9Y/bH4CbLbl71iTPK6OoHQ4TpSqnE5pnpsd
GbevPKb+CN2vku+6n7rC/6N4v+vg38Bb20bS5PFy1K09zl46TwKiuGhRRFSecTBfi10t23WVPYc7
SAS9OsRPE9RM+7oxc68dkOehZAUVczxAwJfelaGVGhZCHAKiAjiYDIVVFm4LyJ8kI8IE3tPRVt8C
k/Pnb6RxBe7DrOQj6+1Ax1v5R/IYsJSDSnzmwWAIenLZ3kF5BuHYBG688/hwUUKeDrAzjBfA6VAN
YB9IRpz0iPGKYUnCv0wjAdUGvPB6m6UydqKdSop+jVKt2ntGZQ4TTXxoL7mZibIWBz1rv0Tw7K2O
+BEYwMzF1ip42/pCsKbRI+ezNzMfPVXcI5ZsofQAmqYh449pDSryETG572tOqvE3n+mVvofSIXK3
JxTv3jRE2ShO7TfZIzsOs2wh0erf4wiQlLcJfeLeF0pWFkYG1PYS3dUV8YPY0Zu9JTHs5eMSSKGS
3HDk5+qCLFlPM7H3muxv2lN9nmX2qRz2qBPj/mZ3NcgsbMhUXdffRXnjnFW1zHCkXdypzrv4MgHO
D6oVsYazQhXHbakFTrTBhme8ccBplFwWMt8uWFGf1WyrP9RuC9PdnCWWcsossA1Vc8kmGNKVJbB3
urhpUpsv31csTx3TxEjLgeVKC4eIZxV3dsfG2jBxHPEu9Tg6oiNmy8AJZkXjSUKL0UYKl9ioo71v
uYsyN1hk/2hws//X6VxCLqN/lF70xUfuY0w4K7SLF/5uGWhkvcSProIX0UTgr5kTECHBQsFkW+Fa
PBVf0+3K8a0/CgMJHbJeQS/0A/HMW6dobxUaCpJUKMeFiiuvsJi8+zaF8V38NO2JARfg4K36ch4B
hW+auLKtWXlR7HsiV0NtxUcbBL7K8oySHILJgGFdNVh3D8Su8eUIAd8ggpKU/3Gfmq22vxYbjOpK
L7eYQ3rA2Q4eAdutawBzNRseAon/oUNblNsI69UjG3eOOXwBaDIKWDqL3j3NrsZPseJqvrVAyI3b
Usozdgrvs7oSUqOFmabGgyeaoVvdAmxsyo+VbxcQ4G3DW+jjvODyel5t1T6eiMZsdgMWtuqwkXoa
Nn/UA1vPiPkjIbNnMKX03+JacA7d8+VUz9sVDZRIJWbWu9rPmNFMBmTF/3SPaG75KKpIEhNMENoM
hQ4kiwCrw6FgiJnVWP1UwEG8L8V1z0hSFp7cAuRG65+lta3Jldt8/EiYh2cmrmcFv96okr6O3xPL
a/+vi6NhEjxC6qcu1jz/VwU50DDNPrJcF6qYUp8tu0n0WyOg2uW/XRCK7sHXgN4S5D0Tk6hNIZ9H
WZz+oN5Vv4aaYGgp0CqV3BNgJ/SsofYmX2gL7Xz5wESgnSP3MDmwhAtpvOQfoW9KvWzkgog3bCcB
Tzsmu4Sv/7kfgLQVb+/ImzU608+KHyyBAKzw8k+pLRKmaTtYESHfALwuUorwapLASL9o98YIZBDB
7t333sYb1KvSp/REtZ6jFpWfmB3CgNkkj0cwIE8BSHUQVsbxA9BWd6Gk7mfhXwrsONYg30OinvBM
8zvNNKOlLMRfCzimT+oSlp8Umkj/x0n8FAss0RkilgFqUfmBHA3xuEEVOIPnpR+TnOZv9SfJ9vWv
ZYLR6wvMbszrShmJTKs5a1w/8373D8XQYWTKjVvPh2/PtDylizdeE6h43zD2dIIi2BSb7aZdsv9N
NfbNyRUaVSOdlSwxLOuKTtyGejw5phVfqzd0R4DXF0+9YKMQ0QKZMnw8HCcuoUMTUPBX6D5/G96a
85/0SQZuw7X2YJ4ZmrRZGbTbh90EvmkP9k67E2Gk2o9/Bd1Q5XFv2iyoyR3xhQp6H+U2/STlis4t
Heildc6p/x3Rd/aC62CD5bNg1x3R9XVXxabccVXVcr9KqqS1At+eWMq+VcC4n9Wqg/6j2j7Wr3PR
NGjSbWCh73pkL962kGBXudSiv/WeJlo+kwyKpnwhnb3dVgm9mjMENBGM3xtGSybuJsjPJHeZn4vc
bDF03vr4o8Bnbi7fxMI6V2wCSTTFcVzn+VcOcYR58Ch5VMjs+d9Rt3f437EsNvShCF2MLjU7ZM6k
CUwFKc+e/UD5Qaw5vjiH+vdWR8zvj5myLAWqEQn36DqEuuqnV7Qx/Qmjox6Bu3aHxWnbokg2tKFV
FIZ8itKfHP196iiE16H7iWCvPrTufjMZA3WJUDzifbdMcXziDoZrZQq5KIPqDfG32yl8LF8njlFR
eQTk4FN5ApUfGvhpkVV56MlmFcSiXPbBVpQt1AQNE+vMgb5L+z7BmZl6w0QrEE+gbOlR3h6DINVQ
xwVqDlC1eCL6TUx3ySkrkfqzJNH4zb8TLYusn9SKf3hTyB5MZiLSx2D8kJps8Z5RN1rsUxZknNms
tOkGkPnjVCjO15lVuLVbn17kjPvHUWentLhR3ZNLgORfDZ8cUhrFLx6CQtUW7tq/2XjrAZnY52FU
UzRD20hKfsCgkrROBAop37uLdxLYUogXqxQV0sIAgjLaPh24HgK1cWTv7sysPYrC7t/Ef9pecdgi
mAcpdiN+vBdjj+d2zazO5UR49vs4HXcABGwhJ1szzGRr0oDzktlK5rPJd9zZKBqFCOOqoRsg2uIy
H2uJ/8Bu1V422OvYQNpvm+THlD19QtNu4cce/yT6MTKkB88OpeyQ9FXG01JdL1OMnC7LZrZO2/11
bkIdre07fDhAY4uvlLvMO+NCFlj7rcwt9coEYx4pN0nhjzkqPEfcwPsRLWpEwlYgHY7YSzigQaRR
k3ZtAIvIktEwdn2xHyF8o0EO70E6tPHDeu9l22XvCtL6cKb+0ybxVeagJsIIatORuFSqeXJ3fGkS
ZQ7U4DfjBNmsdPUavNC3lcIzP4V9U0R2MShVh9e0my4zN8kNyWrk4KX1sp4f6CWGqj+SJGmW8f8K
VIurO0Z0XBElFKIJ3molcQvBCobcS2w7293HWjPyJOFy5vEuXlsVh53Rrw6MmxCGB3+Wdu7HiP9D
tL3xjCHt7jntbsbLjIRjdDWchRU+gjfmdd8OWGIUi6QUFcEDTfU58rpEZGNjpmiRv/nTuZrI4rUm
+4ZKag1sHsSvn0WtuBAzPtpP3bSNrci8zZFUqTDu8/vjHzFPhS7buivK3+eWmR/WoUB3Z++cYCIk
tsG4mhAVcOhu+2+cFHNFHjlijU+E3ifdeBumyAE915dTsjASy/AXgAHL1qT77QbHlBW/AcAN7crv
8dLqlM8rX2aw9KciwXxqnWV6iVS3T/Wi7Fg/ekpSkH7yTtixh3Fv2ZVV9j1J6lr+5yLz9YVVOqVk
/oaYzazAEilyW05xh1jRrbMBpN9ncsO7HY+rs+Bq1CuyHt5ChjRgEPDcoXzk2mGTw0PZtNyYWzEK
MnGhDyDm44vezXdLA+zCcSIe+tcs4HupHbigcSustPqUEJVbsFS7+wtZsJHZWE7KC5giytq9bsyx
hVF/dqvYBXaAbus9Hf10lglU4T0QzFL8/OffjSTMIiZ3+/tvxbK0grq8jG0qQ2C+AEtgBrGS+8KL
M/SRPcVLRIXmm4CgecBjj4FNUN4DLJO0L8Dlv0onVeEicM217fNE2n53ixB71TTTtRxmcfI0C2xC
w6WuB5SYREorvtYldXW5JCpqEKdDfpAswXBZfXXTQZqhNmwK8e7kBYikGrjvMQc4sBOMGhBZFed1
mlvrYGD8MA2L9UTA+y9ikMkXT/v9WN/fsagtIhsdvRThuaa3bhrSmOJOsoqvxpVEls5uhzi6S03L
kL31agvcMYpZydNDtZWZh9QmLzuLxnhZIDuG4QeK63D5xZ/UyTJz2G3lPn3GdlsRA2T/CAlfMbvs
cjvLZCtONop4MENEdazsNbux1OxOWaPZ2t9lHSelMld14CbLeT+SGN/j4WjDFXEJvD+PG1juoXZy
Hbeg1L9RGClTZZf1DFxOSI2aC47tU8WFbeI9QO9Reh63Z4pYNeqzM1/6rk8IcOBoqYYBoNT4H48p
S6hubsEcPRUTnH+dRsBr0Me12eEi8u7Txsokqlk9f4mvGjRZLp5Frz7pSk99QrTteJ9csl1vYmg/
4T9W3d/sJg8iyxv6KDjpI6bbUP+/72k62UG4uWisC6alW9235Y0a34bTvaJul0h7UMWkVGV6rTDR
/CChSrVzdGD7xj4xZ1ve9s9bydZAz1e62vuNLsbgZ4uEaeisS5LZYeY1HqAyrW4AAgJw+Db5Ei6B
OKr0AF65YKmq9tQyHhzRS1rwiaStUM2hKnlg4htXNQTaOdOc+1S7F46UvfRLsYjxBeyu44UpesbC
b9QaZYxb9O7z3Z83tsxD4k3gQvScsR63fMpSb78DpYNq25MSlRq8f+nDIkG9putecohCCJwlntxm
MEJc+ec/FZTw2upkt7b9EzxyKl8Qd1zIYYxSul7xzXts+yeqgQ1K7p88tELU2FIAXbOXGgXJHbKT
QVgBidfP0K9SUIZkKOwTxbKXxWzmheB1yz2y+9CpqvzwMeNlD6/KbMtrR56rcTLzT7pUeXazC9/u
pfhGTNDoVAwXHbrGocoWCLNyrZiq84DMBpkbGw/QPKR8lMOzKUogsKu6GisvdBTMuukWrnvklcWP
pSD+mlJtvJ/XN+s8bBQD36UjuLsCg22bC/+LhprIYw3B7dN9XWgLtQW7ZkB4C+FXDeD4RnF0FJuF
08hfvVRF0nf3jUcMUxehLZiOgyN9fnUoccQ/ioWSLTHyJ2up8afArPfNKvxvV+kau1fBDOZWuGGH
0RsvnaHEekQFKpKfaZrnZwSpbKOWlaig+f+PEjF3qji+Gb4EO7VathCiH2VoMLQl+Ic8UdEcu0+r
aVxhn2A46Kf3YA1OzCHqa88rIAb3jWDF+RIXGoqsI94NWGC22yp1frMEYJ7i7vD36GiOlIV6naAg
nA0eJ+tMwEa5KKVD19h57t1emxJkB436dNL816yHSL7WETB5fVrv+AHjMIMYf83PgVpeuqMIGoB7
A89Gs1Bl9H/aYNrwXJTTPvw9IfdEXLyg37hQGF2eS05iSiq0GdrXVlgAYw0xdDrh8ncNtApaQW5T
FnjEcyRnTIIxgBrrq3m7sCQOpS29MZQT6UEDVdRkrh8JJryNH61tLZ5XOHHo4HYgdMeS8vxn4e1S
+CS5YvvGsqtSkcZ8y4uWOZW1CzQ2wVXpBkPNwIx4Mjz51c7ATbNtSAG7NYL5Ydi2oAkQBSValxAC
6y2H2Jl60GaiwWc9s+swPHEyisgMX1wtdVXCb10kvDqoEKWoNbmd99RpobxuJbQb65wnA6MzzLPx
i6mqmr+nREPZJXcaVuOnDDJNW97ziEV9L63M0Vt2jg+BHRK+vVlOnOlvEYTXJZY9C774PdtVKT7E
b1hwlFshnAKUUIo0Um6yKxSxCd+7WaEcX6XMO9LsD2slu0KLIyYiqhEXGbGrPk819REg8KkSQWvR
ayBjl8aHr2y7brNHwNfZIrdWZ6iQJ5SmiQS4Iz/wqcvi+UpF8ztUSmnAzA0c+JXwtv0Pz2c95e0l
nk7YS58xBT0WkKDrBqH0mHqwBRMxff/5Y9l27Z8RgEHmkHjhICtrbXz/D0T5H+CzBsfAHgpp9WjH
GeOSvf9H+yr+OAMe21WVlzITpbZ4+rez4OxU2FgDen34iWPIXkSNTe70aXr0lxnPxJog9fNWfjZJ
DOno3tD42su4b95Vh0sd0c13daseVf4sHMYpzWNq4zQRBw7osZcy9s2YbQ/OIcbx3b7GDy554ZHR
KZyuHQwzmZievk8cnFGbMsW3z56mtsTnRhc7a+sbvJ3lMpDKmJwhl0m1Y92Rpby5Y6UYlrXyobhW
1gD//Md5bKNaqRakfCFmM9GJsUiqJ8BfW5S/jedejMw3/7LmaFO8VfLwpZ3HaHXcpk+ezw/GOL1p
TsjtIXaT67+PuHZ+UAwmRrvVdRIZwd75ERFQVPX2q+vh/BXaLAcagr/Bwp0/QM0B+lQn2v1bqsXz
RyqX+l7TKJJesAXLZxJKO5Lim7f2IRq5a4AdveQ7FjZS0B8n6sBpiP8vxSJqnX5NbaRloBlJ0r8c
B5tsl7g2HUfSXclO1jMHtQGv13Hddoye8r2x1CxkNIbbGzgHNHJ+Dt10L5GgPi//YhM0+7fH+yAA
eKnOZrOqe5iH1+zYey9ZNNEBy5dnydM393+uJhkkSHBQTDYVyOoNTEDT+9Jy8tSBmDLQZAHOppLV
U+QVRRz3CdSIGivUldxeDM/m50OLFEjwW5PJuPwtWRb4LnHEl++vhd7POR/hCdnxDh03j479a+oR
nXnUMgbKfPeGec/pnL3xDtoItJ0jeHNUW9FJsjf3wxHQdM14EmHd8pgbX+Ekf3QtDcyFOAKvZuAK
dhDZwx+ugLiETIuFPQjKvFxynBbduecA0LvI0trWTh3fqyqfxyWARuwHTwO1rKZqCxAMK2daTz+F
iFuCf/jYEAYVpKNaRqqJst6BjL2hF7CTFnLEeBwtF3ZLWE/netHaBbuB/sV04S4GPS9/hJcg/2qn
XBf9+0/EApEN3G3KvcvqFpO9PeRDe2Qzc2SBCVmBUWESVL0ZI+hWlUBaVhw/RYQ47KNJP3Py760B
XqJATeJqhPwSAuD7fAfw9zotv26bv9NRq3oiqTEK1Oy2WmHIR2sogKH5r1Xw0NmRfQ8DXsU/Kpnp
ZkDAHnGULnrn/Wird8MmJ0Qc1qB1UZj6m6BwhGj7zvfj6tMerUI68GZIrXlyuF150RG5m89xkPpq
uwFg2hdNyPiXO58D9HdbDvWPtk32saDQte8c7ynj/qd1vIxiy1G0jBfSu81p5qDh8e2sFoaqBCw0
W8O7GOwyyWuQRg+CrU1vm0j/xsYw6j1zslGLk0aK61ODXtEzFUm1mQijA+xjv9piRVkt9L2pD+Pi
61bM7SjB0X+/Fw3odo3Va+xHRYYzlDP4gfOFrmLMgEkV41KIKc/DEPccGAiRag7LGihiBVD9FJx3
h8nBsDqj82Sxgp5Z5++uNWjpLrUc7JyMSvT9ewZnP2tIjrbHJiotFOkWI1nwGPCvgCUpqVFYc0lu
PAU7H/dURMf4JrST9L9RzTToCuxQrU7XMsN/5/cVx339XNgnOihjK7TEmW7xMPhyincdNiHm5UJn
gyhmAOdA3Wkp0LbJ34uwjuqmwsjAtvDoVe7j8IdubP+OPyZ4eblbW7Z5zIBNQjlCb3/BsvugleA7
vpTmYG2Tj3Wgj9U/rQ6tHuppPL53DQozXzTsEm5+HotdQi92uxKYt8ITs9nw+g9poHknSZKQzC2k
u514LkVjf2+U25D1u6E6Krgid9yT08DTq14rXwLWzJu99IFBhDGib7N1vjgIt+XXoNlESmfdvPJ1
K3GEDbdBUUJ2gA3VcjQLPGAcpK/SmIeC6rBr5MyGl9XXAqRN8uYEca159kO/m/EbUlMhOkfCXUba
M1UWyQExcJnHsua1AnhioKepSofXFmNlHDzNCx7ucPkIKksjwcbnMv+IBF+ovlkBcWYXo4sArYLA
VjKluTfNkWJk6+MpiMv5A7GVBqD/FVFyO7u5B+pfB/KSzf12+5JfqA48QcIIYBwimp3Pt1d7qntL
drPqnZjquiU35hn1bhswTFflSTPBYTcBJ+MzyxmqpwXIFVoelW0Vb/TnT+PMAPOpvUDwoj+AH1PA
1vFzHw2mahxwO/pyaw4jhfTNAxQpHQneoYQXn/X15rMfLAXjkdJYs8XVo68g5GOh4ICT93syn25L
JN2QM15Kj8L8zXFUW4BeK5qkgTCQYdjVeObVKLpC9a9p6P0eQ0mCNTVjgf2cOsTzfjZMfkHI+XdS
6x8/KqrXgiT/cxBNnmTe2W7jV2S2LhyFRXTQQGCr1fnFsjN5rRmDkjiPY+C7YRHRwmt/V0YthhWE
uzThI9mRupBud07s8hQnxk+ctKA1Aec2+Vz0YIWciF6JJr6g/emX+VQ/E5yUXXSnj/KdHurCEAfo
MAE0mbVIW72JOiM191/XDmZhIDQJe2LzmQ3T79P2MyM/RskO3IRnirvO3JnVqNrQB6k9wDOCdWmt
SJCBRZp3FkuW97mKEywAUi9Zx29xQBiOmusQeasCAMx1kOrHcnbqWzduHV6YMxe6p9S8Ixz64GVI
WBPjlT1XJaQlUHzo2fqI44DyfV7SxAAvGlNLenvHWjk+gB439Sy58ue+Ak86xa/2g8tKr/C7fl1B
8tK1QJgsD0D6yXdFZUE+YpaYxIlVwK55DtCY2Ng50Pi7dfElJq3wRX7q3lvlMQ7GyCZZ6K3ePLFV
B3yeg670yae3Pgt7tlr5u3vKjFoPb7vVszIZ9PmOJiOW/R4siZo5nujttypbpSYYYc7ZAD4Yjh5y
4QZB2Elp7pl57ri1I2mlHrGUAT4uJkNfM29kodWbNgIPiSnJkZ5wWTabMMPv1q6bDpHQD7KuJt6P
DkYJznBUlUhgGUK9N/ESZnfifvNVL1rQQsbjHDM0xS8szzkKFlIxvhARZtQmGoubGQ06f4RvHl96
lo5wclyEn/7nGP4j3AAdL/ztbp69aFyONZFjqdElfRf49EVrAGd1NTY1T+PVg6xrqO/hxXNpAqz4
rroAPTbEDBi+8NYKoTgb5nxR42b+Wr59ZinI+mHJDedpPi5mnsqQsshXVgZK9KvjrlHw7Hv0w2l6
qezMwLzCIZcVqQiH5wR5zPrLWNjfGWR2hof6W5bLf9yi6LYSNeGM4oJSjVS/pKLjfP/U4EKVFRKK
0SSt8IUp9SeJrhd8dkExuwKFGRN+lwQXqnVp/Ykd9A7h+O3SCWqAT3/DLxumbCbYbAdz814Ndj3S
Jf63UoQYMsoEdGLJrURC8sewOKcdry6lqk/EhomZIdZUs4QTMZDqA4b8zWDnGu5IfhqAvBV3eSUB
x0bNeL6lLC95Fw6b6PfwvQTbOWxlYH9RZd1eUT8LkQcUiJg342GIPweK4b1R3bQxoWQPQsO4zbsS
chxMXUYpvovhTVIQLBxab8Dze31tvsnLOB0IyHF4C5JrQpoMDq7bu9O0Bi6G5iNRwqaLdwMZb3Hi
j1/Yf1TrYyzZTytUXk+d8DwODLP3IGc1vl8LuZ/dYqMStsvXtpMQ4iAY3sdVW7sGPa6r8qX5wYfR
5Y7VNg6PCs7l0yQdHEQceLgOBKBxtMCY7FNO6YFMfNxbSD1wTUBYIOvof7edVoc3QpEmwbcfE6nT
xjzMaviaxnMKO7o1inDzYGUfFnknHJvdMyrCZFrA9UFhdpIXs8Nto1wEvpATdSf5cJwiX4+Zm0fr
DVd6LpiwhRyxluIBVFn+THNwP9J2jKMRXc9Lwq36Q/zzdD6ONtSmkYt0bFvClAE95MOhTgIcM/z3
sd03Dgw5R8nc/IT+BXTtJEHYCD82umSqBRVmw7b33Cq2CRkWEXWM2CslTOP+utjODFJvDx7utKQl
M2/dD59KOPk2W4dWqu/BVASR/NPVrDPX4UcZg6OibEuZ6M3vFklwbObynNqh9mlaTirMovkhOFfj
150k6PatT66McO3kzfXC4lfzNI0TGkupVvoP01DoVFl/vVDwDHsNcCBBY2d37TCIR+MdNmqXIC/C
tjbMQ9ACHq2qZ+J3nmO1S84WlhwnRFkCj6C52Hm+3rlDLRpbCimtOxWyyV2dNbYwr8rpIBgyMg39
5YsNbpMp9dhYYpX8wQSlHNmA9okEYLs/qNSxMmeDcrj5rjTNbFfg4g+GmTz9WJnGydBOLJDWg2nf
IfZ6GG5EZqfXvcOM/bUTam4zj3bLizHF7mA+XBpgBDP3CidJ9Ik5+XmnG3DtAjs2xXV+hnZtf2eB
wSeiFMbjEdcnEoHeq3Bi9p8ybLaBMLQ24qScApSy265USXZBnRaj1uCL1pXvji2zXPsySSowBSsc
KkYX9ytlm9F55cs0IfSyRzLU6yKvUPDC6U6oD9LBpgW54emdecztXlC0chvUcq19oIBd5zehJSuE
RHLDVEKWs38zUvUxogMORQHnVy+eBe4CcO6Fwg+C5LOPopYd3cQ3PE8dRLOFLiG2wp3X6Jo8mXjs
3H9Zv7hIpGSuGWPtw5mEI5NDH+5SJJU+/kApAWy7Rtz/PcsGr76kE+/arh4jROhtAy8VuVRb0HSt
bMxqY9nbk3r4VAQu83DMct+qwsQo3Pe5+CEDJ8RUwxxsoJTqJHFMRofmmp7X+NyiYGnO4KbcXYP3
llfW+VjQIhTn2W2mL29FFIVqxgiPeUVsgacV3ha/ok6rQ3he1UbugHXKPIjNF11xyUSQbJT5hLTb
fgHcUeFfvLWl6oRjlRnh6T5ozUYpw38FpZEv9xlyp0YDjibA+6obEUXPLqEdznqKg0fC0G/T31rx
UrQHXmdjAyy2Qs8flb9KDtZ/s/TSofYPyh67xZLx5sFrMFooeYhqIagzfIi2Sw6CfnwxH/0qOnmt
cB99z8mP4GlxQMZJPj6ROqS02DJNnHlIgxZBI6emFWnWH/sbP77geByVm+iW2iQU8Cmia8HVoG3k
0qPJISRC7qI1nKEIL4bV3C3q14W3gHhW/KPPH6KEVwEQz1t511Vi23XNnIy4bLuMdIGmWan/WSzq
mIG6Yo7hCCqh5xpyGY7cppCqq2TllaToJSpG0YMfDnGzB7tfR13ku+JiPLlSBReTD6H57Kibo4+B
ZZC0bRowvRNqqgzcX2esuleVASVTt5iPy09diS5D+XWfDmU3bDtvxRtr4V5JP0zAus9ABNkuxAaM
OWRJMfRL/QvSnaFhGuNpHROWOfrGSLmI3CeT4EaPJGO4KzNnzVPUn0KXt89iGdIRF1vi5PLXl+9B
B0h748zG1xDxomA60RgA8q42X+T+PclWtmkmGihMNIX/Gl7aAdjTXW5RX6f+MYwecyQRVrUZJcdr
6mDsGYyGzUvlZs36e4ZG3L2YHr9AKAP2tnZ9xAD1BSYjYlGzPQMZZ4FnWbOR8qcy+JZD7rg/DWZN
ePlijzdvzEwxqloOivRDMhvFpVspraHmw6/FjuV2s6N76sKMvhOlI/GjgcnJv3UM8k5qOMuU2m7A
NDVyTFFAq8sPLwpJZVtDTXSYNdWHuk/MMVSBOepoNQV3fzuPfgSnlIrQDDJ3/sMBKZ9feFQSbODD
iDMdkreGc4mjhJOeraveDQW9vybetL4r4Ej5jZEEsS1MIPgqSD/QJJpy7bfW01zRY0aWke2jbtkF
x68j4srUx8IhFGrj3h+aHn/TOBvJHlykWch+izbidtZjvfgSpDA6y1Wx8ffgVMaMxiR7kBqPh+tt
ZMBWthWYTorapXGJnfjWFaDHXaLVRtyzKA/2ugjwoMxyYkSSr3NPw3A2u8W/A1S97dXPoUyrsFm6
BxuzLxB4EXAPotorFnIcibjhVaH6genYLZO3PEaSbD957pCXqDbt6xc7TMHoo+4ebiBFUpzo7zD8
xrYvxb4XWUhqp2WNSNQ40/KHbXloP5JnDrXqONAYblpZPtH7ZYj5OeVC7xBHpIX2BSbHOByVl7sR
R9wsNo1g0W/rT19xh5hOGlRO6+OMi71yss3tVN2TGYCSEbeBByq8R/JcoixmZQAguMwTXAYbBrvR
0xtQaTezgULyXRTvIpn5w6QHPvBegmwLWGnpiry0HaaXrbtR2QN8gpiLMdxByNNsaptt8BLTXMo+
z4m92Pn+EVlp7Yjgmh0R3RJ/jNHOhLLqxJtRrU1rmfIiZI4Jd0eP6kKu13CLj1ch8Sjj+HSjIUCA
kheuKGzSMfWBY5m7UjLCIHhsDorLOiuVwUhRKQ3jaaqn74f3hS7P5LKUyuO6kfdU2sE/KGuvQEoD
v7cJt+k0v+RovHeQfavqDxINEHPQXIkF9wav3J6GK/MgXKNsyXC2gXl3qLcatGjrbuspp+LQJ18/
DDKdYlde2RxkCug4eCCaHS0Fy2qQQ+l7XzAjh4HQFOxOI7UpTVMzEYS0sD6afGNCTGfeQ4eb8a1E
2EnZrg2m+wB8mLtsBi1e62TBvreFsxbJQf9N/GFNGJ/0OwbC+6u5BoMaCZBvwMCksadrNklHOCsU
02xVCak5jyJnYbKuw2wL2JnIRfFyattYayvUfOKLRQ2+CVq0XKG0OeX9Pn76CxV3CJCjlquoO8/u
LTw+sqNw9tLIx7bZyJVUoQwfAbKYpqwK+afOWXVEC7G2BohCBBzeX0rvgiL6QcW0k9nPN7C2/SiG
n9KLlHAy9CZ7kpYSnPO/+oQkP2/y9wFnS71DWbBy7yQhmjnyPDVOzByi6q5ZySfmMy8nIR/cQXIU
X+hoismCnt6NPAcIzsXIb68tzja8ompLxDzkimLhCMa4W4e2ZcMnKeG7llQvcC1dLthceSPzzEcR
NW2wPPo4RGOlupZUz80DeBGeBmanh4agFEFpoVBq8o67OTM+Hltz3n3/64dIUefIPW8LjTttQNZ7
EygEnnvRkRKtxVSTVeLeqP2GETtUZJEyIyKA/vuE8fYDX6j6DgYXFqZxLCBSeS3reMmkuXYm7ult
9SEybU1ElIrDB1oknDWrJ659OQjc+cayIv4v45zXSWGaPG3EaS3Q0lVFrC1DfK5Ifw2Rd9RfzRmX
uci7ZF+hqb4Yxu5DGJFq6ndRXg2nbeDOzqQ8ZsbfPvsINd3A9Fy9Runy1kxR4alUW1y9EOAS2wUp
UtKT8v7fs2uRnI7PjAh+XvCMm937hJ7jwTEIjs2rX33cOJA5PHKE7I2F2RpmuW8xINy+w4RRcCNN
K/qsBKncMIANYgzPTs27A/3lwnoAd6wIfQgxQW5URMNtXxU19a6VNRtbJt6lAUDYpCotlKYScGTZ
wpkpUHDNN9OZYO8K5T91nMRToLbGFJfc+EEZUzdiPBfut63FnAkFWDsNfxht9Nq3a/s31zKirXMJ
rpfgkxaOYASk9fO8Oq1Sc24YtHMTD1uKRNT0LnWLzkhcN9FnyScGR+WHuslISQi/l0B96xWRY1eo
2fG+vdix8z3heOBBqjXUL50TUXhulr1BkhmJfhad8oI/BUpa39hPCCzWUZnj6Nd6gB+2iEm1zlB4
kCeAVbHzZYFP6C92qjbWAmFSNMFTylsgy8jyddU4XKc3SWnn/ikA6l0OBQQDCEx0ywqccFM1Smtf
44rYtKdnc9JwE6zePU4ZF8Vet7IFkteXIM5qnrQ2DNeefV4rJRM8V9bsEuFmN5ko93xQ3JxRSPom
fGRtTqFh8KU+XlJJoFGbqi38Gasmz0hthJzkxQoJH5G4mfNKRBE2tgGQ7qPob3GPm4iBG88zJb7O
xAaA+gxo8RKCJ6ytsNfb8roHH+tdHEqqEmZVwxYeCkzlAIwBnqrBK7aM5rZWvuacDnwi32x8l3m5
iYgQ3a97+I5o+Oj8iKRctrpehubFVGMleLPD8OQWI5HlZ2yRo5TeqAhwtbIeTCshzRzIgu4+jpMO
3WmnJ/QeL0IDc9UU5CGigGI9aACBgnNu6YuXDfGMQrWrMu7T/pLua4ovStzDxGSoR1bpdMQNpRq8
AyLCqLoQikSNtmyjgOGOspeyLd4zsE+CA8Id2s4MAcccp3SEAw3cdQhJKsJqUfcxZ17pOduYc9Pq
ooxZTc+z8ehy49Gzjr/ZGgpJWC+Q7XRX1mP/FU+yv+OoK+4JLKLAtdDSnu3u4l2Hkc/ZsQM9a9Ep
ooxVdaV/QO4cjkCl5B+oeGADn0aXyayWl0M7R9yf8mEXiA6jEOJYsZAXPNxCkZWQ9SFGmJYhrKCf
bSP90ky34tC5vwc/ekxvKN2/5dmP41R8qjRb0LuXXrV5ObbqKkSMn6oKv3ImDaZtpo2Rgc7iOs7A
BGDcB0HujM/DE8Ldu2OmZIEjqUP6b9MKRuJ2OODgIlaVb0yV3kbNtODkd+d6qmF3GsoUxCyg0wqm
Z2gl+WLFh5UTF1Q/ckDR8rOijA1PZaXAA0IIrU/eBjX5ZtT1WaFko84icU+Yv2EFNrhh3M8QXBMS
UJs97VN5icrdR/6htCCxBdZwTwVE5cgeyo0X+xYyhB743VrPuti6rniDAFQbRGqrwmojv+Gm/U/4
HWitfYpW4Qs553kKU/QELkJoYxHHWmStan6KEUrxKR+2zvcowVab94ARjqgMYCkBXuw0p6V1dK+g
dCv3Fz3Xg0jJNwymMyD9iDG/JIXQpkX6am1IoX9WF5ASEGm0rsDu/quWZ48/Yeho5GgKAu8Vmo2H
X4rYZjgb/1CqlcaCwfmo0LL9VAanIH+wRzTnIiLV7/c/IC/yd++6DB+Hxnr0W7FPbbTTae6ECQTo
XjDnCt24WdT2VOFTEI9oMy/fyBKyPtGf8W0sJEicJuKDarstOHeqRp8FXRofXJ9hmvm6+2F5wdeJ
QHSpmSPiQ8sqEd4nUM25ACRcR8brs+VTmjbHO0pUgyKNKLj36ZCMjLyOl9L8hpjhu4tvUG227usx
6ogFh0om8iQPjoVorzbW5GC1PUUQng63IQOYShCbCreY0LZFeWhR29U5JnpmNFTKGyn7B4/L8RKI
GRQA43WFo5PZiuTHHIraeJqOsEV9LFKyWbDD6kDKbJJif6rGuaPaqiBx9sD/iJEVRHvzuppSpo84
hx1XdvoSLnBRo/2M/a1Rxc8PHmZFoJbG9QtuXWX5DJxNXFgs0d2Sg/0R6odYzknAon1IkF9eODUG
OwRJw1UTlWx8uyxna3Wu3F4V28RvM1D2duoRr2jElFzXduSQy3iW95ZCJp6rBwkuhN8ifLiGwPGW
6a4UG1vNwMunYVumeErOEKhUM2wsdrbN/ZPdMQnaSxd2xL1bauvyg/1Fbqz6fu7vVr0JcvF2n5H7
aIDpbSatSGlX/WHBSPxBecqDiDWloN8jbJ5B/P0PFuAdjsBdxbQBDScCDf+GeFQq9QR7lFbLe3UG
SSkhMIYwo3DtBegrF3uCtIRpByIfsAIQFJfNxrr7s4iP2j1BT5BYVosMQgGrEXaSsavN7QZKIal8
xCl7WsNvuRohOpEv+mn8onRxamLxd5MykVmdeqSWBD8Lwi4hbvJWQBCENs047jgr4O8HoeQ44Yps
OB7xqJRIV/d39xrD55r2x9z2r478AtclFcJ11jO8l2wB70DGJ2CEY2P/udEKMr7drbQMhMjsJ+Ki
rrov6lzkfFWNLaheVuo5o1geWNIuyigRHpS9t1K8iCDPN0OcMWI5wKgA/GIODpOdMTSc9aZ9kbmZ
ftiOJbo1urXVUoeXUvAypq7yfNX9FUxEuv7HtxPZz6xvUT1GTpSMx5zrmr+mHD55G+J4EXF2YM3D
8bfMiHRqiomUPSsMrRHgZ8kqmUZDfS1ErXVTJ0nCQ8lWzwX9Vn1wsVu8BrOoL4EM22bpnlwtPIXv
rM0PvXRaL7BaxBoEdn4P82yurW9xXzUsKayLsjqJRGd8r5SUrlJnjgRVYX/3H3GPUtOjHWDB++7U
SZvEmEn2xpasLAQbUeS1BmmVQQTV6ZtfzRYSmxIo8hJxxZmRdanfVEUpQFsTEzxCQvqr86Rnospk
0W66+FTRHIhvljrEAuKbplntA2G7aBnf7ocU/t25arOENOPs3/Cse4V2iU2u695MHqCPtPtVYFZK
ZUwRNnGA414kEDEpPqVUcX2AlBk//PJ+gVZdQCyq6vVoPhDGguL/hEFfnOU8bowVBHycKvVM2Z1B
ZTzcksN0+zyqg+5B+B6FH58EvwXrRKNlfMm7Me0BeVwt3A3Q8ZcnS2E/rxrW0rfgCG1C3GTBqgb+
PVaxWjpbMU7/PzXaJLf3T01SJW7QQVh9e8weqkfoUB6bc1cXI9X+DssHbE1kd/t8jFNgyNzZmQ6Q
fCFfq6dClKRHrY6NY1nT5kgiZvq6X3xd5e+pHiRWIYSLKslqwUeQYia3qejJeG35C57Cbvc0gQWn
4e+7vEWrDhVSl9K14i4dyHeKZUNPucmLBfkxV8dMRg3fZWvQGM3KlhgE7PWkVKn7RnI/oNpJ0Sdo
he4+dnmZ7S8CspAo95CWirlS9loXZwq9mjS8Mtb4pBsenwJhGs98NQgDqvfQdc+LM7nRlzupsrXW
XujToECP/qCX0/eQTEVkYLRvnPBlxF+oCUPpSiS6l8Udws680CiQ7jIuctQ6iWc5eeamh8SBZcKP
6vfQxCeOBhwkgYcO+U/HMGHGYdz+N64YKiT/VxVFbe2HNBGhtnC3Q7w6uxp1mhjMl+9cSouccV1K
JFY1YBJjgWjkmFRKsnTBMcYqSbQ8qy8REup6D339Zngvl53jyV6jxshL4et0C7PQUXMNzc6lbIEi
y+0J31ZbdivSTrxOd1c1M/aEjg02Owtyii8PW9g01/c5x2+j2RDtnPhZjppauZO/1UdklZ8hjGyK
e5jHO/u6djpyIy8TgLITRnzFxCZFlTg1EPyAl2K/zgKq6IRBpo7IZUaInfz7WesEtJngSJ42tLyp
OIIXAfsf/tnE5uKRfYRJN1wiYjyg5DrFluKLc48S+IlM8+aG/aUEpTAh1jvX68QMWKycG0WcsYLI
FiU3IDPek9qWWJJ1A1/M7SKS+YF5Hc2qukLAMVK7aExiT/TKMezDoCg+Zu+nYpcXbGYcFQaWhS1v
kMHa/G4y46F2ftpwE4Dt2DPk4BMGLiUaImYdoZFtPtKBlVIyHdrHHF1iOmA6K4y+b4/HqIcpE9vB
DRr5rmfv4lz1woXNCZIZu3+NzzaoOYvoio1DWej28VUA62dIWd/XSfHgzrWCbyH7mm3agfYSyvdh
Rh2s/rNqnCW+CS7CWbziilkvtKFFEAYSoWDktMWMh03mGqe5f7NqCHbv1Uy9y8H+nbAwDcqZeBst
QsY8C48J1QcBnYjx3EwPNbwgS8HWuFndutetp4sivY1Ombcvp7AQ8rXBVPVP4FjBvQDQAIV5Bvv1
ZSXhXXGys0mbCweIYKc66SINy/GXr+5B75975vhqSiI2JMQjXMjuLeq9w/hb2DqK0YpientXLjDT
q5i2pCKWaiVBQ8hpcsbgyvDrlmcgBGcRSIr4yRMQOgfFuowfs+Apy0SIACf4aaxYyDPXfyeOjFrP
Mklc7Tnn8vSG7KjegEe30JRN3QshxT85PFmV8MNENMt4jz9FCb/sOXgBXfKQh6T2n4XK3ejPyHy+
i4XSMMN1Z1ZkRZzfYPct1+D7KTCkbRfzfcYtdiXT/LaAlcmFCkxvYBRIsePynN91YOMrQS6OMKWD
YVmvWH42sfUFTArMnr0YskhhXR1rw1fHjTrcrZ65KKouwKtTRENLu6/g2nFaJMq1s57bFew7DVjc
6a7j3ulYdFYl6HNSsClms2qO4lOF9BKNLgDIxCmfMAyrYWWRX5ryl84nIoAIJY1tFuXb5fScy68V
r6wS7g6hBWlaqi+fAr60cglgpvvOYImT+UZ/zC9nvuPGnLK4bNq26AS7kQReHZqm0r8UXdEvzC/6
qWUoWK1TEmCWZUxHrhM/mRnkaXA9Sw1UuRM85kF2z99vPkNQ7gJPzDW66QGnDMMo2eLHfiXhIqdm
qIbd+kKX3bQMmEhfLj8U/jWwaAZYyhy7bHS8bpL4CxuUqcq1XyMTdMeZjvH5aQKLCPJpfvDNAUxz
G/eStgiJuhCcx2ihtByaczBbP5TYgoeFE3/gGp1NJLOzxORewXhZClp3FVONj0M5b8wih+D6PoiX
XqcGJ/Yl08jRrL7ps74dog+GN1rLS7vcw6Wl/32V5kc9cVcmNtycyCpFNIDp7ESOxyCxZbLjy4Vh
SlSIEeKvLTr4mZeB7T/L8j38zY7YAqnSu6d3xSKW4oo8JZA3E6ad2gIFWRldJcC22+8L/kgitafh
kgPKRbXPzoZymWah4qlo0whGn9bTKTgJEu5iVoES4a0dTn/fJcDzr0XBm1rQbxlAd/rjUkHMuo4u
SDZob9q+Pe9os+bGhdeQ3ylgJwsr2cCtopNvirG1LMoMxqAh38vVFQsK5uhKHO7gioVZNNOAR+EE
ahyYGWJTSrAHVcPXnsZTwIUa9JLcsbOcre/iSde1+GwGjSVfs4/4ytr+MIZneTGO5aHdYujJqFnX
4t+GVocZI5Ify5tG7+KPj1v2GJnfABwfOfRB9ypHwjqTYrFfnaY2JuAHtESYk0Hn5ts/eWxhYBXL
kxHDLFgr1fxL9WDTBCXT9QPQ/zhhQ9g5GE/LYPJNCOaZ0paucdG2QJzozpUJVe7HYRi10rPHp6Nq
Nr7Wlc7HI83LnAd88x1bX4KkUEtmbARG+rvSppNAnrnPF0USyQoeWtaynEJZhrmfHK8EnlBSePEI
FpXrDdZsSkXQ4aiiIgfH1PzpVIUjrzX6BAUUJIk8GvY0F/S1XhUwNq/oD0HLQobAI3qjVirI7Pc6
NY6zgPkMWvps5u4KYvsZ1HoGpeTBh+WLP78zeRuk10pfHPbI+yllVJ0c434ky0COTaSVyR7c67aK
NCdksfo27WlXLk/tnl76H0qjKsHs80FFRpMCTWcnoHJZ3JqFsYx2ZMMc/IKhCpRPJz9IE2Iwv34k
sK8l8z6az0XNs0TBsSIwqvxPEmdK5nKYwRU42xPVErC9em2O7PfYL7FB7LDIRS0gCLj516Lgdu7n
GXG5/UkLAXhGtoXKztfkN2XyxyVJh8ykfeQziX4mnkfHsSz4a2TQM75zIdIvDcx8zFDMPFWqUmpv
rwr8hbQb5oGX3hW1PLtNyteqiEaYM13Fc9Bn6wSukjtzkHOqG2ddBOazbs6ohmyayfbeaU8CgVYy
mAnS3r4eKV7EFm3mu/YqpfJZNGte6+Ak8ozOOo1V2rOyQ0PQnl8LjpjjIksavNVOpyCom+5/zIcW
UgUSU91VqrXS3ZGL2N+9Bj1v+o72+JHPE5SVxCLfwCz0UvLJdAPgOd5xBcUzgLIqKpflbzC9OU7z
xxW78UZMHokqgLWkT24QykqnGWSS/lE6YBTchEkqtqv2YV6vaOj7pozG809tYWR0OHCnzCOQ6EuS
O1phexhdGQggrZVUu8n2K6EPNsFqP6hYm/szxu0bwQQB4XC4sbXTtmW+VJ3mF+3Z65E5wiU1TzlQ
KZ3ulyu7WlUYfUYsfVeZssY/qKvr0vNq1GcEipskC3Sf/HFStws7riqTUDp1GoxuNAlv/J+/+bDb
jrRmBTvPBl70YpxRbX8YMc/li/6fXnAIXjAz74rCjC4FwLusV9LRf+RG0Kn0DCD9ClMAqlh3z0Hk
BWmCWwe4+rtFgnTxfQenOPuAQH0v0eM877/TSyTuIkuYFVNUiaVTvr4qd+IQC0NnaFfX5cKsbqTy
lfOgNCkx8ifNFnOOMsc5yQXBsz3890ggYD9ipABI7nlODr3LvmM75ccKe/0FZq46+3yB2rWmWAvG
QBl6shGro1QBIolT4rOhf631OtL3ev6D1qQ8oBgzcc60E7txbhsGrRJto/8thQduYh/7jVtvnVLa
ciDdDZDDbFqMrnKwvAyjAWAmLRpf96gmInjdPmcre+3O/73CxT+qg1Svuf5g0oDI/KCiitb6D6yP
HUSv/JcaA0FjwdhmvPI1zCmwaBRiA+5rQRDtjwxM63LKBGc3cm7VMyj10LauPmKTBWUc1pOTg1JT
eBOTg7DwXsPKxRvcf2BsIE/FHSCtMgp7chbN1T84av1kkpW/NgwwF2JrFNi/ENF3ZPUs76bWoWhk
z66L2NjTkFE18TX0LOJiDm3FnaPLohN2Wam9aGHrKIxMLI3jQGEf323l5Dsd0uG4B02CAf2f/3DV
nVqQwgGe3QGQ7kP7jTLusVtipVYNgyDf66NCdtm+nkWaTpK1z9dqMTS3GNWmKe1CZ0yWriCuEiB3
gnVjlMGMBS3yMXhND+UKhOvvnBV3ygxQglCS2rMM6M+d6tfMJkOwk3qX6bcOaobGoaOahelV0GNX
WRBDZH+L1LTSYrsIixqH18liEm2qSxjf+njDUwoVCPdZlMGYfZDZIG+5a1MRjHRyWvGS1UO0atEi
GxDEYJAHOVMSy39rYur+DjCTEeWqycx461/0cA1KN3+31o6z7RhSA4BSwN6ZPK7ktYOyFmnJP5hs
OmOj7o1PMlSuQIvn0k2MPWHRY/gs8c0kzBaF96iMdiCdf0bEGjmFHDCllhfL/l6gNcvlMymI6wib
jZJe37eRL+E/S8JfttIBtg/QBogxRhz0FOiiXYqqGQX9T5wCoA0N3EnCTVn2t+hFJE/SgiLkzZQ0
LH1voMEpnTtp7JFQscxTDUK4aJ1itsRMC6RAl2a/XAVkxOrZFnrbyhmTqih+wXWz1RWtbNpFnO2+
UR7FJekCcX1NGiZtjNoENCpEWFf5bU/KXX5sl8xsS9Lu+Mb8l3M1SiXT7N2nDSI2aqt6TrdDCJMe
RLMTmPd/2vzOMaXYw2URg9JHzZR4RVn6stExmY1OyktwDc7qNIuRo2mXkYaPRT5UhGFR9B0XUzJ4
MOH3AnuzSbhLJ8Uz6+MK50z0UXp7fFJfrpEDv5vKEnjvVGCCbes+LrVjoU8B4aoLaNo8jWjDatYb
8Mdve9aSYmt9Bb/kc1K5uSOzAolKi9UtkxYrrg3yhOF1+0MUhMuoRh78FOiUF/BjmVy/DYaMwfMJ
8QjINSTykXJnvYDEx7HC6nsdMR8A4bC9hEZWy+v11C84SUNxzWnFijhu0GUN4RIOlPvIvfgg2DU6
nQ2KwK6RZuqq7wbYwX1iNHyjLZsmC1XJlptUFreH4WjE8ihI785mMWXrpvXG3Gb99PKymAGSo1IA
Zc10KCOQAqPbWzkfk/Z/zarDNrARAD6Bsf8XGPPvlEAZZoSw0Nsi4BW+mwVu6vwlZWYzZawwdq24
oUTpqru6EMOeezR01sq0PCXIbK5wb29x+qyM8AaGxFoCpS/k4Ht8DA9pgAlgXVgPgXQ3zjbSadTO
kwire88d0mNL6/aLs/ey3ATBJjoaLOmTm78AD9ivPBsO0SRRNEWZ6Mcz2UYTxHwjISnARF6cbzZX
5UatKwB6+GCQQv/WXDqLZnw9S6aurkdK7qvUqlbfM+K8NULO3bgMegYL8TEkqsPceKjfXdEATa1J
JO1klEmTKGusrmLDIx9GdV4NmemRMlEs0YfPhgmu8SpyXxlsxAy/oXcRwKuDRwjgtMYIXqCrN3ps
dc9CxWIyBcZ2Rg1pnKE6TrQeYaN604KH+iYAQxIb2d9rcQHihJ3nuviUptmAJPDgFPo58v4ANHLR
gXvtCl6N8kN+E+MwkApzF7ks81DyC7c26hX+Ozg3uP5LlcHyeTmkvSek/eOlNc2sdjNzq2imf9Zc
Y+yCSsNncAJ0NebTnAXgBtqN/0/dGMx4EHF2tEeXTbLnsjQx8ekf18DIl9/7Uc8SZg3o+85+LfKh
+We5AU4keUkHcPZ7TkG6NSWFnCNCeh5YlhZ2WxoiJ+D2qKgL04POC+Zl6gIkB0MuQxuLFP9T5Lw9
7kqXM5Geg9Pl4SMrLyAbWSCoiySAbuAvugKGutisXnLqaDC9c670CvMded3mjOL9zuVVowE9M8BR
N42qLP673K8yvuVMkuhS11HCv2yNBoKfcyle3lH1sHzVtaqZceseH8q+oE0eWKDdh/KjAW3PTuuX
eSaMKVxaF6w65tRmAMlo3F02we8s6peD7h5k/GhnO+zl7wDtWrzXXSslxNFWnxB/QfTf0VB8HGju
eAitRHRuVkPPo0CW8t94EOBr4XaOuePCEPdqYqARNyoE2Il6ia79gyOs+Ix1qhHzAssA3qr0fuoZ
xRD08bme4HITT5A5DRMOw7MVacGV4r8lho4GVAWSHy06EU9VqaoZI4e8cxh+46bRTj/OuSeR6NX9
QmxCpI03Muq1zKmq4Mo4V2BszNu/dSQNZSYoSg3IUQxlAkoe3YDoXtzxx54amYSE7BJiZh83cflB
2Che9GaYt2+mFSmV1suLYhHEz7ALqp4BzKAVm+jRDg3u8lLFqw8K/oy8KBoJN0ipKmXW03poAw4h
fzoKia0PjA4Fu52KdS/QGtuo7QqBWeLm3Qd8pksBnwf+VN+NvgDww3Np2DROq2z4G+QkXCSHWauq
ORg3SoJ+CfnrRQpmZ0Q7tV+b0zvTKMhg241eIn4U1e9HUm+wgnKi4zoAY3YcNeYKqfwvmxhVBsMp
L2fwMiFVLFSCPBD+2rEY8+d8IrkvcqSGT0TBB1Vw8aLNDM3xQVJCk335NbSBBSetkU6X+hqrXVHr
Kgq+VjKcqAy0+7dj5yfnz4ccq8xspf7tw3NijSAMnjY29cpP6l4XXwa8qxZPGXXOXrp+bIJW1yc4
ATgjGhCdyy7tdJCoFgfR1BorcrTcprQNw4sJyBeO6eR5hkUHT/h/EU0Bx7VH5gnvvCNH8cRlWY7T
3zbGUg0bJFN/Zae5oMgCtp2UqsdCqCa2ZM8PZfo60cYa+tTKsJxaDFRPGuISoEYGZnKOrGnh4P1S
nqF4/vf/gNQmLFZQCKEcq9JW6SZYqQtCFQZ30w8Jg3Oju6V4KTcHGxaqPfAZQZEdoLZdjpLzrZYR
x6pwgTnUfFwX0zrKh+8jK5O0JPNGKbQDgzos/HLEh6FSfePQU9+gh3gORQZUkQdbb4jZaZJnOfT0
KJ05wvr+gM/SjXTJkeTAeunWfH7tPF0+YFQrjYa1inz1CaP1Hhq6adiLuNuCg8JY7M1+JwQNfF9H
90qfItACDMjPLJKFPxX3H/UQvvTP5l6C4MAdduZ+fZTn7TphpZqVBTdSfi+bpx5bQ3nK7OU5p7NS
JIEj+QCWMt47MxIoChkSH+ui5aCzyFeaenUTyRk5QS3vNARUWMXYBNuaf9StRlkGNoje8uynX9JR
+z4MjlU8Fti923yfPjxxByMiinArOc0TRKxsU0CpOPOJcN7KPforrkIdJ72cbYGbszy0ru5/eJCm
KX2QvHKTRdfOr0Jh/B3RvoMZem5nmZu5p5sful2fOMFAlWUJGOH/mHsbtXjh238wk0XXNvCH5Exr
Xn+6YgvhEUDEiW3ouU7RJ12tXkJa5TzPG0ZCtqWpArL1dflWFYiSNJakbEhszZQXlq5q5Kp/9Nqi
g8r+3Gll53veNt/tJM2RQQv0rcBf42fK5AvoWTYvVKzpx+4X5pqiAGtgX5LCw33o/J6gD8BhKUxj
fioWCRPNi6ovPfilPWmXWQhhT1euVBuouQA8NgzTxXjpGvXNCXKS+QREiqoHoMYo+koMXg+irXFn
lbMl6myeU2hrgfi0oJLMesa+dCcKxGMBNUer7fhb0bVLLIDPuNTeSIdSdieBky5rnaw0GhyxM9uO
wtlV3Nz/69lhwHgMy5IhhvmCFnmEOvBJLZ8dvkkQ36MDb+ggY2tR+HYMxYKiCx8aLUHVPCtc8FN6
iIV5eIweo8kfA11jHpE60E37qtyi0pauli0Vu1shnkWOUsAYGJok84P9vmLsdR87J7SMkikzOAvC
R8WeAgktfdecH75kguQMrpYFmHlvyLM4eZ8dY1pe8L7Bt9F2YKl8jHEDYNnjVOSe0O1zcka0gmoN
M6AXfsLz9BQMfqtaAI3/WeM5fU+pydcOzMG2uk0mCByUvW5rU65B/gTI6S+NFSwKK488pm/9yMf+
0jIbHS9SjamG+Tmmr68lKk/Zw7RS2cFSzOfE7Q5A8aDKbrgxcLtT+rjH8hhFH14anJWVDs0LVL0P
za8er7GSSqj7k+boEGdYTFscD7oiAvXwqv+sVDJ4J/QDe1hHvbryRyF1VCQe+YMYi4eyXg7cwSHS
EkmU+ymBSTxUTLYX0VKw0sKOddHDX1rpacxIM/hpgAkPODyT/WqLiByV4qHafScdon8/vM86V6+0
neUnldpKoprV2Y56KfDA8DLjj4XoBc6lUfan0ncK0t7bXnL5jmdr2C7KmBd6lPA0Sx04I3MOBa8M
YqopB/WHd/5tMy4UXHLC9zhGYfq0q67RhDI7mieXnM/UlOlsI5nzLZOMAePso+aoYS77vLaG+zkz
/t9YzBvBfJgnxmQsbdUnJWluL52tyzQ3g/awE0i4a1HlQy3Sq3o3la5rPeiiPLyXzWxlEqNHzi6D
rRCgaKxy8zln9WFzCFWLeyIcLQhUS5iv1HDRJZ3f+3TwPHjeyvEN5S0Yr6cjDiptBG/Y12Osnl5Y
Qnyuy1Atkmtrp7bDXf+KjMzY64N+rjozUshowtjbp4FtlenpiqGJFBAwX+JQFO4bvBT9MswtfaYc
ImlUVbjivKbSHf1y0xR7thDjHAiM7pwQrGjwMt+64xiFoNcTs5ee2ZjynDHytX2mSuSuolSsmyOW
A75IgpalsKY7bDNb6KlcJvaG3UTtFSAiT5R4xnTIaa4DaDQ/T9qfhfyGEzY+0oR8cAo2xvnnVpPn
ERd/T0TRJwMjwJXNLTINFzTqFUgjZkwkXZJHAFYsz3aiTKV7Zg7XhDaP7SXqrp1hesmnRayQvkb2
dsxY/0vT+bcpd1nMhNEg2uF7C1JMuHcpIKeWMGziyHsfq1nYZzxmtlAOVHSpUXFTGTUf76GjgNlf
VzNIs9Kw86p7pHYOFkRAbgQyw+Mh9DaNPvkb+4xdGcZicjARBRT0mciXoyNM5FOarP3cYf+9exQG
6nDd/pq3YJ2kn3GP291LqeSZBEKpPGH2Ms8yyzHeBxkz2/fLrUPNYeOdIY/i4ip3R4/xObPPEH3l
Z1Gg3AYHAt61kC4grseTO1XKweCjPSPjvQ8EfsqfxOYOwSvrnpBeWIVhy5KtbcC2MOZjosjH7M/I
JxTVo/1W7nercpiOs3HoaOKrBKG3NOCEmOD9uGhUl87D8yQ0ktwc36I9Uzd4rzUq08lKNpPyGZbE
kR3MhW82R1jH7Mwxm1UjEGqbSVVOoekN25eQ4MHtrpDgDCjMo4H53Uqd1D+O957HruouF+8WZKhG
+vz7kcbDDntlXeKapYCBOBFqrBcJRU3rwGFHKPNGhGdIARP7k6DCLFN9o3kjksj0BtGiRgCTRbVR
uRW/GF+uCr1r7OoBwcZvr0Dll2SmUpJyj5a+LC7q6LfHxthaPDH6a0JznvI9IGMUz0PNFLU7dc5v
M+jsjnwt8OBH60nh+jiGti+soI4Lam3QBxQ+4Tw8YX7fbEd6G5dYj4+Fkk/b3ZKUCTb/RTUJQFfV
YqZZRP39DkXfY6ELkSnPy59gfYQdJsbjpxWt42fcAIt/qJVlunQbt7uPTkrzR4gUYrOO2doTLZvC
LMkvib5wmhX2AjVpAPzQSTglosARcebLrMC2rFtblk761+TL+jWdal/FB20Q7G8Cbi/HtUjXuS8s
RjRDoUpXsM/O+wv0F3XeztV6tMVmifk6AfTZdGXZZnfGPyJtep/Eh2XFILCujvU3nq3l+U1AToUp
JwKjG90ylMdLm489mXWONUKMJdcBq4oa8tZKyjyXe3UAJ3+DGAbsvRIKntTOzdD8JA6Nqq2CHfs1
6lIPFSbXuO7NsR2O2n7xexAcOO4ypx7VjS2nVa7uP0xBR12E1Ql4TLlrPVo7fQ6IEi7qlRAdip0J
B0KCiPqA3QZ6EDLSGXTg8JIuZwQBrxxBrUsC39NwjUsciIZvnqNT1NDjW8YoMFlzdf+l90smR2zN
ddikwNfuwFex8Ug6jM3Vyol4BphAqiWwDMe3lLYUbdqaRP2MLLo0R0F54WzTQ4k8axYVufsVBxVH
zKjc0aZnTtoFaM6IItNYe/x0OhHfqGmpJI7GdeZgsXzMHNIWX9NFq8Zd/vGP/2ZX+N838cDDS2th
rdK8DOpLlk+kthVyOUwwFlkl1+kmcrM8V0RvDmGvQn6C77VBAVOkn+aLSfb+jxibuFbwcw6Ja4Lj
j+ZRKrDITQzj+hC+HhSZTq/6RGbRja8N9Og1ahubR904YF2cJFDzkkH/gCL+TKtbgfEKAgcqoDKb
TB0+dplr8GImX01XzvwlAOEW609I5lPRCvWL15LTZUZdWiBbeeaHjByMaMeAcI3/NCb01xCiJzU3
k58LzUen8gOYhWyZWJBgNmN446TdQhWEbchHT97ppSnOxv6KUEVP6kZw/mAy6Hphr8FO0BDfBsVt
fCAtnTMP5JbEX3TRNPYDUCcjOvixGCaSn8DVCOQgRKm/pYbllTnZhzxRMPhbzE7nH5o6FTPQ+t2Z
Pc0lNRbD5wqut5hNmOCXZm9F1RMGUvuFTdw3QY6VSwy5+z/9BmYHRTs/ih60SrmAYZiRyiENhTqW
i0v6/fTw/42Uv4yc4ygPiDGssx+yw3HqYwcSre4Rixqxs5jKXUBRugS7tjS3EXO1MxINFv3VU2vm
ZmQvcHWpfXsHUeM5u3MgjlcWL2x/QDw5Xt+x7v4YBOguN/ChX55hJ9tavch//d6pd8Hr9CnM+pxd
bfStJPPQgUyGWaLEuVPM78/gLmmZ2gtpRXveps0M41xog2tV25vw370iuhufqiqhmJ+E3xcGfBeu
STBMw+lg8YkZzkNlIt0taHAEgeJX6aSjKdEHJ0YUjTfP2kTRG5vhJp6fTx+Cd1TyHVBZRFH1LdYz
UaatGdV8AHSGs6ApFITSElVhWLa551EhuqbpZhLi4EEpuSXhK6F+IxKdD5cwx6r8ph8WNOWm5tJm
h3GUXF1dfAmyz/u79oK5X+Njhu/kOL52WisESk0KGDaVeqprRU4yAQvERxaNrmd5QpZvAb/g4Of8
0f5++bRfuKUFXSPkuLeGsZM6gHMKbls0V1WY+/R0ebaH4H2TXGwiB9lgkAUcZjNEJPqReSQktqAx
wkVGZkxcohZA1iMLKFwvLFN4vbZEoFBcHiPSygX6QzysE/mIgl3QChgmQsrltcomsThoP+hmOmwZ
wGTAJ5VjuG180zkYIdJ6k3GPI6zz4XiJF5u+H5Nsa8vUcZDuUYELP06AR5OMJHuyKV2ruadBwpAg
85Egahkn6nEJ0AThDIHLuBnJiV0kl8iptlO9ZUaPJOyCve3jWpSodVvrn4qc4DntuiwVoueaFniW
XHMSC1I4N7eHdFwXRWe2lN2jtf34m23s7UhaYr/v0VSdB4twCKKTi2jNSbmTO+xnd5GFZI+PvfqL
br84k/XP29riQj6J2V0rP8+PfEYwFe0UIDfv/8Y12Xb0RMpMyBzVQvi88LXa9+woQ9yLREcQ5vH4
hkj6k6cKKCkHveE/wRLj9CM7lNXtvrFned4IaegVTM7fqIzJI6Oq6oPugjcOZlaKOy3F2UYjtjHz
LHdO9K4q6es2er/prhWJbstQm0lyWo+aihdpEGWSQiczovpt/OMJZF04fawt/mFUYWwU1eNhAi3t
WUsfQ+Fq/0B5OEOXmC+o20l33fErxtoQZGFxd5BmWoL9UurZtDwu1Z8GXhBPXA4vzWYEMsAR70o8
+A9IB/EFLPUR+JZ9Qyfq9MjvvQ/QWPn/Rn6vWndxBkJ857No5vcK5lKDIrwi8m89W6wYZQ3B6wnV
a56qlqd0ZvONkZO3ER0s6lh213TnoFPUJxsVrY6NIzIJcMRqtASpKZBiXwC0J33/ZeSSUCjtpfDW
q3+f/mbV1kikfMCF2llw70UC3KSdCiqZ1K8ZLzoPISNTI/J1cD4y67saVeHqsCFrNlSQAP7PrIYR
eFMT8lAz64ICO3Ifp70qGHZYaJF+8YNIjT+6L0cMyN7yAIBtFPIbSJ1Jsh4eI6X3pFkFdqI1sJYX
YzplZJrH7d7Q3hU67yr4K9/9cvB7f665ZmqMvoI9E8NHTJ/aKH0tcWWlGtmsxrdzSyz+Mrxbm3Av
/C+fAbOPl3OG5wf9XlOZ95qjC1pZ4klLA7MrXkF2KpVg71QFeQrvUn3/TxW9m3x4U57ug90Mi1go
/u3RsOn66BKccUWLiZibiES9JK3Ty6XSe7YdPI+10o4ZHAqAjiYYpyp1DIn+/uRfdhDeMJX2oT+4
5EU8swXJsRekkdgRapEptI7uJ9aNTZCjuA+v0hweBZY5FDEGZ/la/YpeGUfeGQgcwnq5xt3+abb3
39L1PH9bVDhLU81cleQ6tkDnEhDuJ42jE9jOTguaotzo5/qgJBkiA+DGNhLfJev8NNAELeZ4zTMV
eCcRMwvMVWK2deovOMOEPXtSQujxEx49ZVCQso7iP0qgTISFF8cG6G5jL+J4Ugj5E7jQ5nDZIyNR
MlRzpOkaW8d/7V4IxCrLS5QitqohFggBGMAvXelj85jn0S4oh2smhqaMaHhfavSgkqBUL2buo5s4
ju0bkvu8q2PzvQ+3T0PBYZKN7kMmsl7+vpKViqcAOaPAEUHEqBy/zC27vGtSDpW/oeJ5QpfpHtrG
mnSvzNM27zQD/W4Rtmo0xwj86Sn/AfmJbMSHz0BZxAHvYouM/deSRldA0LgS05xu7rUSv3CWCL1L
IhM5rfeKfMpOzFrRBM/W+oAW4aB5lYOdyA4DY84pCIz6VesjP3EqYrZKkwWEbkDMxShziZNBR6s2
/uaFBBtLNt0mmE85ATlIhr5+CFk1955xaHbLSXsHJgeZSo7jsninBcovgOf8KaSnlhuxAGcVpgAq
RFxB3QCHdaGtB898LL43/A9CSCKq7voBSPKmXuq+uuexlM/dWaYfVrnDcUJexYvJlxjyBxzq/po2
itDXWlXWAISsajE4A3CoZPmDO1Pk5fGzouGm7j5ElYgVFz7SC+dHbUdZxYaXYO+hp4R6hfII7Zj4
7e0lcj7Zn1Z3BMRgaiNt5tksbmRJ/7VOeZjCQ9k0eXeQNDFaoQcOSE980qOmGmXcyCecURBjKDS9
o/cOP9E+6pGLN9xucikNhFxI/9RkV/MBkx/Vin8b6qOSDdazDpRn8lwxniNwDjQHLl7UrjAFHkwr
7q5T0oy/XuCzRyIrkHsfV6M0a9DWe9c4rwhtbarD6AmixSQRpvNcI+TA3k9rQrTAR4Vi4pibzOy/
27xBDwV1adPu9Ts1DKYk4ZSJbYe/wIQ/BFKF6ke8OHQcCcDgep77bNd5JDuFIQHoMsP0ljcWmXM6
79mJAjJHmMQ3omFNecKFX5MfqglVcYr6xxB9/wWJfMroJLaWsNJV1sMCewR27/3ig73AC0FUk6H+
w7aAieCPq8RPfZ6sKdEViLPkYOEmNlmkgN0HmA8GtN22L9OYLbe0+37BgGRiWwVDtvBcCAY82jGk
9A+BYDfLIGMpUwum/bIPQyfLZbYDWk1lfBFXmJ8KAlvK3kPk1QC3rB8pGQJ5XfwmgqI45LV9o+7K
BPytSDwDq81R5DGICXgierUe3HvkCVCO3sE0MbUs5qu3NIx0F2K2J5+vahRkPzwxC5s9++bHZhvb
YGBealOVVgCQ2ZXjOa5Jbm5TqB8KoIf22y62OikwtbSiniIq8HUNuga4Yxpn8fVm1/2s+i09JZa2
b9ELHzPDJH107vBCVaz+xHsQJZdvGfAppg8PNyZLjoZVsBO9UDAsVZ3ihXdDVovSyhWTlvAc+j5Z
FuId1VEbGWmAOdt5v8VljrRs0vwTCXhiNOaC7nJpjwLho8xqapLHCGlm3s5t0havjAUn/kgpegrw
GUFxcXBfXLTjNsYK13WgaiGp+EVn5PEPT5ZWglxgoa+vhwhPqPk4xVZkAa/f+IKCZ6hMPQKLSiH0
a2EUSa+S8yblbEPqpU+PTGfHiOe8pzol9YCmcCdKRcACuRgUBe+xrP/wO9zSaF83kX62bBYWks6x
Lr91w+oyvVLrQr1nj0BkrLrip1hVf8wA9DtgMIJq+DZhmP4mmJk1FMW3XLa2fRfTu2M9Pf8Ck3pQ
n8RE1Wd3t0yCEyftnSRa+Sgn9E4LIWRPobB5P50LHZ/iqzy8Jmr/P3bHwjaJHu3TIMu7YSg6CnGV
KvpNR451HRPqqmuW7MX3WlbLyhjoq41+HC90sHjb8CnN9b3tX+sfAjTud8Z0cMdJjVNgBZjOEcox
0GfQRYxFqKU9fxGJONTdHS72qh5dQcS/9n3D4xSMrJHdmoHgZ8I7X/VesvuQ5YtdcmStvYXhTw+o
POv+JJQFNFl5JD4eSF573R4qPGElubGgYX2yIE0Xmc++iomyG0mIFgmWpz4+RKJAIrftiObZuBsY
gq/hibBc3/BdBPTcxMxlRh5jZaFFIdk7mE57Q31T8GkrBKwf72pbLad2tDpmvti9uIEM9pdpi/TC
Y8EYH76Dd03RoFHNbzKbY/Ye+Q4FZ6qentmMEM4fvJAtqipUpT0Aa4cHQ18lAWaMIz6lDs5lz/Ut
6T6yRwc6qQmwFlrle5q/up+hlj0DmqoznwIRh5nb8M8kWzEhRbRIC8lG8pmgXDUP2DK5fy1w2b2x
5gM+aFARUGwomykImane6qcAntaYfBp47aNtuCoGrdi5fOuTaj/FMUsG82VZh9FV8bWWE2rlaPBs
b+76veQucU3KMgEUUQNtwqZl+BAUL8G9KU+RVa1yEjkVYB2FfWpmQCYc8cWdj5hwFRSlZ25Vatqh
TtKKWUBQNN4hSNPSkEYcqrYOKLgL4VPL+qk7qhsEmykmCVvhfi+hq3WxHQ+aj8v+9IujuN5q0GxV
Rzt9ERES2BKnyXwDPB/eoh30V7xpthw0sdXUdTm0V1qkP56bfBkKRPbLNE6KnUD7QNG8du+inRMU
KsW7QeAuBnYrdf1amRaI2FLDbH6vSU4z4iOThDLH+IL4Pe4UwlMqUmzUly4HAxEZKnUox7amLC5J
ynvLcEKQG6ytPbajUmuJRuPyPrFaA/fBWlV6lnWB5x8zvmA53bpq0es42fU/SSPiAi0ELxpSsv/7
FEIIZYhxR28Nig+UnAnyZxqKgIFTgJfzat+xlkn9vYpO/Udcg4RVayJ1l6RZ7jYD4M6bAblQauEB
vicxcvLYDTC2wdsbJnyB+BbWS1J97NK3uzxnwKbjhnJ1D0q9oz6Efbv83DLDVTmkPM50syhzO0wG
b67szpdZrzYY/FKWn4Ucq0cXMxmo9qsEkipW+MPEc3niOolc7grvGFIxxYNt3QAKdHsoDJD5Qed7
TbGNHkAvbpijxo7WgIwIFhViZ9hbCiHQ3bRrkjSvEhR3JcdzcsUlhsFBywuTT8ahzvEzdFdzeVFX
gDp9+cG881G1nLZyPy/JFU0To4G1p5BRuFrnhWSWv3CQmp82Nli5iawyS9KkBOsbGTEAhubX8ZjC
qbMF2tIGuv99KP6QZWoIEZFfE8zvjW2i5a21TDLjhowfazi25ihVpGGur7+v9Rs+0fUw6avRtQ/r
s56X4QRjUf0uNDfq/ThyzaWRMnPjxXaGo0F3PCWIA0pnmLRbCAxsJa/vuTbJWIiGTAPlTAFQRhDc
LjNG/wFxrNZrceJQy2pijTzuMCdXHkjvwgIbrmTpGEu3PvYuxujM777WmpRMrijtaM5ea8oHVa31
/6QA2A==
`pragma protect end_protected
