// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
lpVdpFIPuy+UnIWQ4WdCd3J2v0XRsYCQt4K+DAr9tEnwyp28cVJ8CkszWlExPLz7sM+Kheq18mBc
QLrP/oZWwhaYcDH1NFwjwdsIDvG5ObkIi/fwemSbOG8412QFfrlKAl3/X/z5eeQyo8cYLmt5md7D
deXt3ZNb86c0Ba6lQWQ8jjezC+wAjUE22Vuyk0PQKO8orNqjyAAbv6+YGJoAYJUdmN+zgLSNvIzN
W8LCouYHxCyEfidZ0Zb+b31BvDHuOA05Ver+IkFwZRE478ULnG/l0paiRnoJaC4VAwuzXWriBbAy
u46Uum1S1sADjFv/chTQq0FglEx59GXdQIfPIw==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
Z8IcIqa6M1/do6ZUM0KTU46xexwVn+OL0xQEz2PdH1ORttEVYc9GA6g2UOXnSXX3lCXNaCrwwkoS
HOLqu7sRO8n5jJ1mOvdoTbnWxXu9I6LG3SKke6RU7lVYfITKAhCuflWmBPxdirW6ktAvS4kp8HdL
kuyq4EEr/NLRr+qowrT7NgsCYjuEJsh/mbfetbBofPL5ch0hL7fKPA4SpE49i6m/RnqD9q+epOXb
DCmbSEJ6W/FFTMBhfGkeVCHw1vNuZzHYNdGLKMBWDeWblRyPO7+Qkw20V6Utc3z5Lq0Jxhcgxh3j
XhZMd7br7AGmua2fEMzAkzytyQCPcvLv0Xi7kTRzf8b90eyKNFGLTO5OqJsVPfEQj/bfR2/xUFBF
MGykBfC7AesisaE/yvP+mrOxcQfIWFVspw9bw8SG9jyRTg4okBAeGhuPU4h2whtNuilEeIR4cTsr
1cjXCYw2J0qwDZ2xIgUDoncILnuZ9xv3qe2Vsa2s3b9TvzfD5vV3ooseQfVI58HkzPTXDwYG7aNm
u2U38RD52kN/80ACPMg+UG7AL5e2USqawOVVlcn6F8slHf1egmGcJU6jtpMUJp4OjlEcNmrVy/Vk
2Ez0cI/Ttz5zxggNXl+JGeHvdL87KoQGmMAcJNRUJNKp7oGmePP0rCQq6oWbTPHLWwj0fD58I5Fj
JqGZ887jwIIAMyystGBF73F7Nys6IT+A5bfPzYNGiS0H4X1ZkOJz53oOi8QrUJAcDuQjWRzc6awc
N2VxHbL02LUu5VvSpE8pweY13RqvyFGoVZ3AQ1UDpvwL3bvEYU4d/JuoShmDg0pitCo0XcN9TRBq
L361FVIz4SZxU0lUCJwN6B+i/kfwwhr26ehWuwOaPaW/HwNwg15d3Xoic9kTj/5dy5AOwwJlBZ/e
aARfApIuujlvynAqZwPDgcLgCAZZTv819GR3Lfwk66zxifEf4rMTVbimbVfiHLyhKPq11uB5Pc+k
1nV4afeMNMptk4EELt0pXaIqxYbj4DdeHly9YAHmbGQ06Sjj/SOil6VEpTPuRryWq/g7bOFGboSb
Z5MwoyKff/k0dpjoTZG5nwXJ3iinriB3zujG5P9wJYfBT+ypNm4DbvoeXslC6oblGFwgQlnwuJIX
YXF/S/5IruRT8edQZ0JHJVuhSYZTkUN/0DHQDYjXtV1EgKhbDm3UqgwDAIkx0qGcQ5d2IC8jbOk5
j2a23FMd/8BQ3mvuSprVwki7sqUnS2jW4GBLmJxfs539A/YyqE+xpgSfWQn4Kevbyb5SMAdhQzM8
s40PphsLUZT9l9Q8Vv6pFdqnR1x42ycR/aM7wXb9YNJsAnoAdMvXb6VX/gOga168VMyRmNW+rs2I
xEEHJNVeAio0nzZeFkF5Omxb5OLLUZGK+2kTw7liafU4i4OdsH2aU2IwDcRIWGwiSEw3Z1/G8saF
KbW8+/lJn/CDgomkC98JaUlJWXIu7lbO+RiHSM34dgM1+wiHbexOrzMBeuJ1x8pbh8RhE2Ke5kUz
zYRImN9X27qJ6R0TZ3KW2RJ5vrt7IrxDH0cCJyQMBMjQfMAVBJi9puoFgNR/V+MsicMgtEjs8bZA
SWw4gxEFLhjMEycOPi7vJ9+BhDSARQCNq1qtKUXibuYhUrGmkHTOLvlRxE+jTUBqWBn4gvvjUghq
cvg9j1PrVZbzE8iUsJYXhrMzZR/sdhCKU85ipSKd+v41ro+pD+XJvTaqnt082wDqRX3B2gXhO8qF
zgr1UOQfBnCSfB3IlNKFp0xEN7K6dKixP/SlAvJodD1JQjBwqaJXc4KaUkXMVfxauNFZrvIeBgME
QCb1AntQfCt69XzZARdx/r5u8UrFa0lcdr0zBVKVYgIkcodZmLPRd+Q5txmxOmWIKgabiYAIVWj0
EibmeE/Zw6Qv7VyiKNMv9GMvbLJGrlJ9sBgWLF2+RpPQ0FU7+iPiU/TQUu3e6X0+ogtsO0bBcPjK
9W5rhwah+wi0cbuwvLtJDbbiAiPWGd7sQUrynLhs0aVtOZi/WBvE11zRZ7S8bv+vx+qvgYbOo932
hmii8FfMQdV+p5+TLokRjvHXQPEn8Tq1r8VljuZThbLkTGy5RL+HVUzWKCJj5YLOyj+8DS6Qdf0q
GbOHiZdFPrViFmRyhTNX0JE69WzIpLuLuA3J6Dwli/YyrxtVxb0p2ak3JGXaEd9cVX4593rTik1o
zTn3vZry9ldo37wi1zMg5/o1GRssUsh6PToeHS5zoRunNGTW34nisW/y9q/sQxxtCqj960hSCjEW
edgo6hF8PixdEh+KlVQocXATmifAs6xVS5XM+ZUTWzS0fxr7O8TOHsEdmpRG99823uLJGZ7scxyZ
Hjk3AjYK3cMboaEwjERpHJQ5Hz9dkazqsKmwkMXwQRttAavRnmBf0zaUTuAxpA4ffH/riJ/an2ff
jJVfZ8j4K2rJO/ICgJRBKI9JnZSTmzOVSFz3pDH8E7XWztFVzAjT86pBf4dt29r9hSBR/8d7kssc
RonQJRg4RU2+lCkmacDiGLKHomUUDXuZHL2JT7R0LqdNrLT92jfg/cSSXAjtQOEEsrc2TbBgtgLh
K7npRlqx2KEWolORlJcW4Ao2gUgD+0xqfZAuACS4Qc/3bwA64bSomE7A/shahJvUt7WhVEUqyhOJ
GnIeswgvXQrZUJvjHuV4T30xK6Kup8gQItNYYVu9yv/+kQkq2GBa6WhX92LRmU/4HmOW3AAhYie9
/b5oKzLOF3W17D9sHXb8Y0ZuyTaEIhtP1NnCDiR/cH2z/JmrkySru5ndvRew8jp62be57SKKJ8iV
MChLlzj8DbhRH4mPP1WYBAwMhqETx7Qhi57lIUk2imehRAjIEfD6m7QZTjw+bIlQH59aVmFZgIcJ
NQe/QFkiKeB7K+acaMSooWgeCJSTIpWZUEdCmuEbON52C71D/3eBaeyRpiPMRqQGZo3IVk1tuRlG
df7QgpNRtp6jfMXT2WrZtFayAsuE2ASRzmXEGJrfM/dlQk2oX3/74TQAGWKh0uFMMbcs/TQ7f4Dg
dHbFT3J5qjJAflWaGgEqEeONS+muMUp2sxdFZDFzGEdid/25ztmX/8kINB8cfeCBv1PEw3xqPAkL
oQukJd/nU7a0G4VO/B9KCLHE7hdCf34Zza5g8QxbzrIe6RiVq/3gAiJR5fES67+6aAcg0BOAbQot
cGjrx7ZDBgal4kPxb7nWJZq35KoG1sOm0ky0VxIrnOP7SUX1MdXfFlN7AmHqDnmZF/vqjTvSoeVU
BbcUwH7zauEGHvy9oSoX44jK1DGXhlGDmo7yIu9LDqvBRxnow6ThQuT0pKvKYRnmnmYrC/Yb+LR0
od+2eIRAifI6n6m0f9+OMDDtA6mBgsQeHDWFyUuRrGNQRGAfwMCpeaeZElSb8JNWW/XipqhhLpST
B5/6MqbjZpPLAfAYt0jwnDNKt9vPjF3vAVeXslx9zi8WRuC1hDe9tfgXv4klSW92LnI6nwvlA3qZ
gLg2nZMER/dzWiS7CwjPwlgGtkRe7ykJ+qZ+MtVTs8ILhqDAmVzWIGGWYdn2vjdaI+aE+zNXmwMQ
kPTXB8330bqOLrzaBrsK3g2yaFeCkdjl22AcbPK8jXnf/FGjpQANgxD/vR1Xxh6nZv9jIPB/TTzI
y7GMtLUKyCUmBqGs1mT9HppbMabdUxF0tCCJL23kkAdmwnfr4Bbt7+QjnHqyFvoawkXtBbu3zb0p
GPUvynSNDLH0mBT1qRIEPSxq0nn8wfCJttkBBUIm5b1ISI51lwh7Gt8WL3eEW7aUobb2o/MNzGC1
UnIysai5XnSPSe1cB8JT/ljwWm8gBg9T0GBxGnAKztDL7fME8ZSQngrSwGjdLP412zQ/XIGNkN9H
WcNJVlV28yEgZjMcbcobt2E9hRK4+6bKjlxfgdPaDZmHm4S8xt4T3ccljou1GUQGYD37jr7TJT5M
bsVLRy6kxRqsC7qky4HnNQThaojf1wpR1B6diWX3dlQRFi605o8esZv4INy0gNeYYJauOfqR8OJu
Y4MZmhx24Oh4Mpu5az2R/cf5gPoruNtJKIm0gMXlBY5YjMqSTP4fhLZibOibfiu4Ndkr+VB73k0i
nPUczez2MLkMwEPtxmXGVvRpotxqHBC2mZNfE7ItPgywFZtEkYqz72S1MJay+JijaMvexDET2HAW
chvLmfpMUiG5gM4IfPZ6/NoYeJL0wtbQNpTzcj9cPb5Z6bGtYnAA0kWdY1gbYe8i8+jF4qVDxjkj
y9wZTgXKmSxH994l2Snjnq4oUsY4cuVvUHzSiQpk2zuU9BVs9hnQolwiX8x8jMDcv/KZn1e2rCXN
VNg9kY2J73LWQSTSJJ/HBR++IGrVzSkmkbsbuXt91iwXbPMRhEf407z9+WI5wsbQ75tt4aFPsR1a
epapxbkzuUNiQ4Dz/6/+vRwog5vSUWtklxFQ9E8Ay0AwPg4viKEUVgGkTG9DO8UP1VIifeR2cqmS
B/NJE1u0/LCgRQsovxTJL7BD1nFMg4FvLnD3VugLdsp76NZ35o8wPcV1b8f1USjwAQR2R6QahJAi
rhmbqmGysnFY70Adz2AE8/Dvy8JTBztsBX4QlbhgxTczfx/C6WuZdS4p3QHHzNuXPvInG39rn4ct
pAgdvlz0rFdwaK30qJgF+lrxUkX6BuA9O3iUKZT1L+2GcnOUMwLrRMPyOPDqMyTTx1ihV2tB6jio
d0hPZTbgifi751QRUzsfL7PkR4eCfJ7pAi9VDDyubYfAYHK1v9KrK5thhNEDgCy8mX+V3ipWyGJq
HSLvg2h7o0L2nbSt1FDuIHPm7OllR7KoJDeN4QCxWaS5HHPxJU2YqtYCwSQzGniLK5aj9fVntmgy
EnIk5Kv9Gl10lu5kMN3MUpyEVQdVihR1lmXQnEwPvf8SGLiYJF/jy3qUesWtJOBD64TZf7e5jcHD
RJM64whM5ASMUb9AmIc5KoZKNG0lZWOeQks9tFdG39D5FmLpA42Dwi5qA3Gvx6vVRh4QG6UO4Ctc
YOxUpI1xRMlBsoZZB1vr5OWnZZsl5nM1+XQOpA/HfIvNQJJaA+/UK1mZNiXLu7MEANmsXARkuQVG
AvAkkynV87ogJtOGchZbC5gbszDU9sjg503DGt+/HXu+ezkojzo9JojXf1KZzDdD+RZx9p/fc69l
CIoXsawOfSSobNP/g/FNcFTsqq9BdJaSmRlE4T3IM/ioBaJ11Wh/Qzus2xyfdiNtpxxW0ZOX3oLn
o33J+OzVKA/Gpj1OQjTbdcWxd6q6yuxfSq569558EPKMDR229pcUttoN9OTGDuKYKUB1iNm8uGLg
Q3r01Lq/NoUN9d7oPBOtACNRcLE3v2ZP2mbQ4VVsNNooavaoDsE10OWAYGfHhT93XV0Un1UvqQdE
lqfOn6sF/Xff+u1JiIv3jFFj7qwEdf6+4Qcz3R1e3FlcYg2sIT1RRMCcJBpDTCLNIjYE629MjnfN
WZ3VSI3fc6FFJbIzWwsdyi8yeD5hi/r2T1C9K1tKRdFAdrCbr2t56am5ZzbhoprFBnkQo0ytTK8/
nWX1m/BXMJnosYq2rhR86yZuZgfQ0IeLYMBaA/fruONslHqxCWOpZIT/Cdvd2m0KK5xfQhXZpHkj
HF6qkG7rnCOkc7eeHi3CtJc2PL4x8qnUMT98SA26ADTLsyiIXh4+mc5M1kC5gNyWKZgP/0qBBha7
zlatqv4LpLUeCKqPXO4Xi2gNDoN9IzamMCapyTRm5tVqVM3crA0iI9TnXvFjjFNy/zPHc6Pzntbd
oPGfyg==
`pragma protect end_protected
