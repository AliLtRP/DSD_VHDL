// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:24 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
IJTNPk9zi8Pt0sn5Zc/ibwa9VwOk2jkXGZzCgiqChnN+mLzwUP2P94BVtc7pLplj
DpjcSMqWKA8BkaOUZiJjeGwR9esZ5LBcFC9qHQlpAJwYMwL0tT+wN0tSpycLYANj
zHPy5NKwCbm2xaeuQB52NR+Ex/G3qrXRj5ppJk3vSiY=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 6816)
k4+Sa1MQg3AGbNrX6YiuzVowvuhGSWmrqJGvcq28R6Hn29m7BXiRgBWNIqevjBez
bFtE6St4VdqtFHWek/tnzSOZm5+lpKEtQiWUVKWLiA3qpXzrjE0JLHab6smdNxdB
PVAMmOtYcx5oCCLsPHXZ8M2O9ZGIa3oKIeIWgMaFgy+yUpLUjWSfL6QAEKJVeG98
522eRnV8kdkAy+4Z9qn+WZ2FmrABhVXCVoMKaBKyzZJBAsjyGwJy0MaRkWfAuJyb
JtCuWuMXAYWAdTCyfkqn3ZfQofj9y4jTyxKyzAUKlDGm3RFyqqnuUHuKugARFu01
215xU+GrTILz1yZUq6KMj8FM+mr7P4GTcygHUztiAAYalDhAhMInZsNnuj3NdXew
iDKCF44NdmT9SZw86fOeOzxhPAsxOghSjua09nWwRH612dpB7POD6KqSJaCZcOqB
omaiAtB+vEIlnoK3icA5NlgRXMmKrF2erIEhMnviKO9R4tcaxTpFTP/CfMNu7Vy3
dNVn2zLqf7cFoMKpvEkuxbfRUgBfRouAEHgJv27Dl7YTrJjtTQDrwvgh7954RzrO
syS9JLFAHYkS2hBBvtSugIa1w9mFCZn/UmFM8slUIrlapUMp+OVUmlKj48nkEq2l
3oPc/FFSblQ+Wd2q7ZbOt4gGWcpdCuyFIbKiDO4Cxh8uZUXoObsrsfTX+UbfrKfr
PdNnCnQcVcBYBcAXHXdOvniuWNu1UTuq39lz+UH0++Ze2kwxkFB54KOY2tDuSFaw
GpNTSu9R6vjdcV6W8dD+cyhFuQTC9rBgHNCKCr1yIWHIEfX9X1fuxklLWP6Ko7kV
ETyqY6QneNjUItRs78wcNY02ZV4lgwWxTCrjwIJjDSJ15uzq7XB74xyYn6g2usAS
RHinOpxh5hOt9V9X4MXCcfzFhjWq8iuYOmUmDq5LHAj3WthAVQCVEorkUZszcV8G
pgk+eRyqOqp6ChX2tNjOqSzRsEj7oUuo4L44cyEKlkUij000gR75NbzeLQKdJ5jH
t7sOHzk8lqUwJzIzMKKo17l3qSMA02IiABdp7ecc/9wOMHb+6XZmkrpXtndEoDME
HuN9bOGN/6JPj7+ih9T2pAmFr5/OM94InM47DJ5TLHzxagnzguKuML3J/VeR9s1l
ybqFDBOVUwYlGlPkskI3tJNCSlK7g8WHpXtFlVIJTtVKctUZ20NqetgEYh4T0QCt
2SIHhZeOcOYVaV4+WoSKwShQiNLlsxww7BdpR0LX3kDHFeM51yy4/W9pP6ByZpmU
aCV0f6DSrAIJkemi+/Tlb+gnn15DY5etJShQrjop5sq0WT27Kxxg5C/tDVtFSqIK
KvbrCN9wp4UWGBgBfY7CGYej8ZxLXqBxcHRESwjbvanGQPkWvNZ161LCMNwJPHqF
QRpUtKNgj+wNsdqrYP+pGtCqFUIakKP6VSIFZtLxTVuuv7hPoizbw431q9EI8QfV
IHv7N0FWuc/BYkCFckAVrnCfPQMCgEwkJEIcECe17G3C/ZByrlLrbWNU2B8m7Yfv
d8ejCf1IDwy7Yqe3qVWl9L8YtpcMToR5yL+KoXqcaAwT5Wg1aZ3dyF4ZL0N1S9FF
RJDjCNLofSBWW6YaX+436j4GuHZSVxrUPHQxBYoKwbF6TiUO4wxSf3L7Y9wPZLfn
LUPBaKDiZqA/ZHE04B831EYvcOkOBFhAnJMqSvanuU37TORvTQpVO/YBytpCVZnF
l2EkrCGO/joKt5unWNPrw/2Fz2WVCUO5eVri0mpdonjfsSD6Rd3HNRXF8hyTQ6bu
lXk5boPpPK2DKtikGf0KgzIWm5uEkvula8SVO5/Re174z4fiAUXwW7lgAUxYfFUG
uXKTHWF2pu86tOxdtnt0qFklKxyQGHY3jeTey1Lty8CfQCLpvCHKce1nsuj1YJXq
dZnGjQ3Mc/3gdzOsgJ8TEzyyOZYNWRNDb8vTC832pthczFIBLuyqgVBIml3+v8Hd
f0wvWrKIFz6+MuZJl/kjo8rlehl6aw0ePVkiTlWknHrM3LSxDUncXG3Q/tyihcQq
Vm+D+xQ5yhS7XH8fHOmGsGldpnW7xXSKiEXeWjFb7NpELLu5lmt+X/bWg3qNAWzr
BHgPmJHl1RIHxVxqDQI7L/owiESW+/fifcSt41UVZ4jXKzRUJbSu3tC+rPuo1Sq2
dFPyCY/CUDQcpwvdfCut5fvwRvcZ4+eCXX/EiuLFDQSzgPMZsF/J4SxnxbJg0+wG
RHCv1R9bepG8Tc3fbdU6L7/MPCp4rJncdu0pgxSS+ldPLvMmMyqzCnSovBU4xz97
UBKyyGjusC0rO7SSB5qwcYRP1+2SKUqGGACu2VTFgRJy7EbdmLroXtI9njQXruAE
VKSqAO8RoNzkJqLpOYvkWL7sa1qOBCzWiuMzq6sDaujpxvc7DbJy5xu2uC+gFg1r
kHW3kJ7LsuV5+VH73lva9iT+5A/BOuCq8MfAjJQd1JA9PBcaixgGsjsNIqTyQvX3
9YbCvbzkgo9PEy5S7z3/TFJBkLrsL50GHaDLxCJMp3zu8F0kgEZkwi6kIgwDUpUl
Fe2N8Jwb1FwgHYMwj1RE3OOyY+rKXlGCWfe1zEts/ooVyY+QNV2+smZBtKULwTFv
y/K22jDEP5fjbiA3t56nsnc5ASbh/+IwXjNQFIJpPBvZrMBMAtzdtor5ghgl62/R
slaks9zo0yzIjOkDTg2qYuSBPJNG6eYYSFac3DNFojTL/UCBeY1vRx79E6s+jQoO
3rcitiyO5x8iT/+gcuzrkkYdkwaQJEDaAcutGPrff9b+sgS4otvrwiGV70Cq/lpg
3xADAl+Suo3m9dRcUHsWLR0uUJ8zswtJUJw7x+ECaKG2B+lwXDYll9wZ2V+1abtv
bw61mzUzufZywXu9DwYibTrI9ymhhyZNYKJObqq6j03oEF0MGKXv6g8I1ESKMb+z
xtv9RWEfMMWVyB3rqbnM/9Jh6ou1GZOYlPLkr3Eq71Dua/LuTA76bux4QqAWog5Q
Vwu/rF+crZfjnkABckR47k5vuN62J6YJc+6GwCV42n8OmpS3/1bIowOIJfdctLHb
apVZx+jUYcFg44tsqwdWVHn55M6rWCsW3DcFgANlnSPdtsznXIYhPoc0vG0DqT+E
NI5EsUQikCif6/f5wT3scwRIjPxj2y9dlPpworNraaNFj27W+ajIORmLoBepX4/X
V/K/S+Ct176Z2dtNAdffteTljgmpXWUI3JeVYxK+kGfaS9LXMD00/SB9SH20qf1Y
5Cy8BFKcVJwc3e7koENFgJqv5lm1qrmFWsG8sYl9xQHD2jZzGOZz/wJw6jUuFByD
foZgsNUSekUPgCKmGc8+Xecu0m6N7gOwnWW/atlw5At6lG5XH4Oo1foqsFcb+KyK
knuTqmP71FrzhB7b7+pKCwS7dezcU78Vr5zdeg+GEhv0enPkF6NQ/l0aa6543A5N
wKJodbh29BEiLJwdPN3qqeIRFx8VAmNafARxq46DJdwLrryOxlOdWMYtaYqj23Wm
eYtiH8dX5LJw0s7VDElq6NISDvhyEM5Evaf4RvonWMFf/HTCL2jMp3F0g/qPGdyT
sZXuciIlrQANYtcLLZo6utvO3bO2cVzE1uA0NheHeDjqAGrBr9dtsJTdzbw6VHBP
I2eosy0V/wuZpioyKir/7JgMI6RmsY1v4085Glx7DTPl/tyv9JSrMPGPno8XIdHG
GdfnKd8iXcNhBxcz5oDWgcR8tKZFFmnozLp937vKsN2W3NyVdSqd88FdCHPWPQNm
unaNHqFIVo3icgFrBmEgfNc3KS4Nr4i1W2Ivv6DLosv5ExYGEPPrErFCWrOGl5tP
vnmO0SFxFkUnca092y/NUE6ppWO2XQz0e7rIVbegB7UM0mjImq28dGZV+lTJzim/
NufhKefXAEWEH1fl8pGW3BMvWX01QqBVU3shgHa6FVtnZ3/FhftC0NVkKPHr6g6P
mmsW58yRu25cQHw2af1G1kF92BmKE2kKpE6d4KGeCwWpFZn13oCm1VhnWS7eZ6l9
2cI9EHzlGnvBTUXgOtA6Ocy2DD4DYU1+a7WB32l8XmbpDJI4hgijcOHJV+5RPOlO
W2m8HPBXL8zrCRnjSpI27iUQTNU2e4D56bBjnFb/ZEZEq3h06DmEIQtL/wYSwnyx
T6jNivguzpDeO5l9SbBhw32YKkNHEVYz3M9LvyhNx5r/18LxVwh1LKP8iRmeo8UO
lmJvXCQyBh5ACLZnSJbX4FXn7j4UqzI5iCi9ryFc+q/Py8kFjLReWxYY5PPfEjzs
yErNQgTdNRoDSVf7oNtuyVRUxVbjzqwz+Pqc3KmXyRR2ggJY2h4iI3QiMVHSVOZo
AqGkJ+oHgXt9n5QcZ7UvEe+jnkPOnlP30uKQKLYjN5pcUOH4pa8POoxfJe3kJNWA
0jqPvglOkv/ItQPqg4Fe9S6/FjXlNlC86o79SE8HioAAHvIMoJPb8lwtp6lQFSBD
SUPlbWCA05d3n5HB3xtf5ZX7NoPIIYgVKUTuMJ4NHhaengzdHUpHjEf85htcGMTQ
ZJ7yQdkCQF0AU5wOoqStU7oiX8CEat9rMrZlIN7D81qViM12UCdkfbHaeAbBFZMj
O1ZL3pz09RXnY/9Mse8Kf+B+uf7rrea83fnDdcmUuvs1GMID400dmBiSFM//9TfL
VVMhmm2pY2qXj8YMOp0K4SIWGKTAbfQqtEbHNKWAnZ5kl85SJYmehnQKyx9l3MoC
eV1oJmM8Cv3Wv88/qo3lT3JBrHttNrWTMM6aLHtfCDnFX2PwmwCgGBe28XPVoe85
a+iCKmMk4/fznV2rhjnqqAB5Yx/TSkCGbK5uiSYOwRHGdWi/GZav7+W07p1ww8iJ
lUUtgVal9qqrneIQ9iZseNuSwZwO+mvcqKPORqveNkTuiRrstt08bYrGWDamkNpI
HcflpisCryzH2t66YJnuyAmsLYD5dWLlqtF/JsUppZvmxTAxJ9KTfMeFErc53U4G
/yIotpTKFDDdxGJuqKHUco92vJ8iuaAEVH0ychNZiDDnQ3zwxWFavXRFYr13+AuU
/9shxECsK2mT6HkVeFHuW32BLRZB260LQ8cGFCl473K+HWxjUwxcYR9zs2sO/Dqd
bphyiW+P9ZR+RVfyf2Z1lEB6s4hoVRUR1UXB/5EB79UPnWAvlhi3GtdZ3YWjT1QA
00OQyLNVOxEwnaXgWQ+0fwGePI3Xtir0DsZgWd6oy1XgY0N+cpP6kiz8ZS/fHqoJ
dgS/3JYoKw17rtQOqztfxm3sxZFc/+ffgexhqYsTWHVn9VPldygc43ZiJsgbb0LQ
+8QcMYb3bzE9IqHyEtwHmMIzAaZ7tETtjXVNU0zxg6lPYUzmTam7+oCr4TLvpC9M
DCNiIGClpTWbikeoIet12PgeO0/gpRBHcQJPGzwn/sn/mBurfGl0dFREM+PIV2y1
cS9C4MteH6yCxthCwVgX+a4/aaMcnysdvhe18ayih0QH6nGagg73XxhhqQQikC1Y
LX6A8ZDbD4gWTwN3TmYzs+He5woYQHTZvsFyD24uoNvYAumY8syS7zNWP68+xG0E
qCgHhOPhuLzMhdoA8atVD0BytrV88u0fX3Y1hCqJ31DTSLbtNpnkLPYsC+4yBAqy
XyL6I8iYOe43uY61n33igD58GRy9W7L81ciDOcP4P45XLW2Q9lC0xlcjwzvJ62+P
7SnqVib4A/m53TIWEI0RC3xsS3DSJ3DrjKAgYOf6QkVU1AWKcT0Rs34Dd7lMgRrf
kdjKU1lnvuRfzVZlPrMrQ+708hxLF3ddpqOJVd/KvP2DNCA12s5BaNHbc5keoCPw
IB+AqhBYSsJqN4ZHX2k4SdvIL9EIkRZdxZCr2kWIAuFGiD26InFPhmMa7URymjqs
Mgof2LxKfaZoshz27gPbsnkLJyM+YKhtCaezF+qCm4ckowz2Sqki2Ap/OvzTvnBF
vpMGYYO9MKCZWabeZBeKMgtKLtiGJVx2FGJvM0+dlOVcH+/z4c8g0wHnutBFoTHO
bZCWa+2UoxkAWvWsEY6Elk/qynx4VUlBzrlFytIZNo0LiKytdgy7SCnZ3gJEg1D9
L++DPR8Cg5st5cYXs0hJdYpsNiuA+Htogd/FCm7GuNHYoizVLF1SUygR+buIVrZ5
h32mQXbLIKYeMFT2bm9Pf+jLgc1JwBZUq28/0k+wFagtKRxbyuQbn4Rv3Vb7JKDG
uZ5FsBLgpydacOS04fi97H5RBPYUGmLdlyD/pzl7YK1SfypZ1j45gwJLP7Ssr+Gb
3pWD/Z/CIFJN0ab5uP8AbAQRSSm7R4dOJN+C1iwU2F5QL2jubws8fpBhEufPlg7n
7w2Afkb2zGeXVlPaSv0PFtQCJzfmWFVQjITsRsaAg9PGYbnrXfdAAtk/DAVNLTFd
0zmhNnCFqafr4clo/+Rpu+aoSqq4x1w+IHCfGP743mcdJVojucUUZo03TU7oXebd
KKYHfTJP5aXfaMMOeJZpibXEiJ8m4WbTkeof9sHvWjsGmwVfc29albYjp1LMQ1w2
fh41R8mkQa8utJm7fiseC7YVnOigC4z42s4X9oQvxza70VKmXKBvNEdandFZ//VR
WK8LNHA2HiPVzIQreYApu3UzwWFNztFnIEY00oROTnbCdOkrV94we1j3DRnldtUZ
TjjLaeYZShaQuG3y3wFcNaM48+4xT4OD3PyRkvNqfcqOSfg6bxiQgmcwKJWmPOKQ
wt4h0JEih5rs2JbU87sysu/nAqkqxVZOGb1tjmur94VU6CChQYd8i2p1h8rPEX+3
zzj50ut6P1y06x5J2BFz6j3aSTW/1EcxGlAIh+JsC0nRmniUzd2POVqhJxfo6Yy5
Re9M16+yCe5DjRuOPn4WfPIQ9cKI5rOGeroUVpvCzIBLq9qS8gYMyjqMWxzV8TwG
rHQx9T9GEMzM4Q0iOIIRHYAC1UJnxQUn/ej4hqvk5K1I7zmiT4J2erZD1wEU1l9Z
vEiyzPDdiLN5pta+gIVkH0lNCg5E59UwcJNM/WmVO8s8kP4xnvfEEf7sLwI8gucT
imUa7GSvK6uvgvmtFKSa7YJF1LQobSqkLNsmYAM0iSSHsoB6xUFwAFDiRTTwB1MB
eDvSViUlYXxOrLc2G/LTMAGAh+5y5iHHIcyA8RtAcFxFSijs295REe70sJnxk8so
tLQ3ia+c8qhRpGkzo0f9tcT7IUvQ8hpmeqdD6qZY8q2xRqvXoPOJvSyZ1vCtN/KT
dGyKbZsWy2iNytBrp+dHzEUSAfp9qHhg0i0lsMOzWixEuzCWhMLDlh144ZM1YuES
1zb4I5DffhF43QqqKjTzxcg7boBD9s5i++NSeRssq/LIV4ZeevCswnX/bspzqSmP
+Ao9JarwkE2CUYb7crn/Md+6gwS9DRaHvMYCpF3co3uUN5hGedpVZGzj+eE8TmYS
xiQ0t+S+8ireAhhNq1xXoljrOjNq0ekGBj80KYwlMFRVDWXQ4ka1DBpSNjmw4mXY
us+/LpYOTwrVfoDuJVsFVLSosYPuEPVQsHCsV0FWEYys/2e5PE5nWDxQ4aqSPox7
mMgCsRWU1PXnZaClcxLqY7m+ywQTp1NmLxGLDJGXb0NPHMxhUr77uY3Q9tzNMPy2
gWXdbgxeaLPFVrwkKVplSz2OYBDYp/PYnSok0oZBW1aBDT/D6p74VMefSLcZ+Yf1
KhDa7ktsn9WWxOgA5LA+o0DVo8SxQToTUj9/NF6swQwlVDyp+MCnsgSNTCchm8Er
YVqCMtHNYVWHGeJiBMoD4tXtadMiUW1X9goi1b34/YM7AOhH1/ViGLL/2MV1T77X
lleJ2te8TjfaEez/q6qBIvrKqhwhSuPP/ftZ/0WMcFLmZLc8ig2ZuoNVpb4ODLew
WvjCgAnHX1i01jEClByJ/86VJoHdlFrb+8fvmjus80ljIpuvr7ZXpZRik7gNVv6G
V3oTer8Z0x62hfTgP/ygqIcCxtzV6iNdwWAcjlNP0afXb//TYxaSzc0kDo7J2Ckx
u1mMQEJcOEkAc3xu2AzTuBrrLEXr0Jm2d6S5goIc4gtqVPx9ylxDVuHrhOGTiPG5
p+nlja46CnmwK6bOto0ZwoReegLBHdFEuISBLME1cR8QBOxkX7zb7jA4fL0f3Dn8
uzC1/TqpFk8v7+99xWUN9aX6xP/qGyfaEP2bL91q3PXdHxUw8Z4oxh2ZJgzAvJhG
c8G05n1iZAYwFl9o6pkMWK119pW1xokBqgblkKVuHgdbidk8ltRD4rOjCnJfTnBr
/B/MXjVlSRIYk0QqSPJWyhS6tF5NG8/Pdg2FAeZPiInTND6OYKcI/Li6scr6mdQh
JyEmscMeocoEQd4uYDEnRL9ix4hLYX9/eYMm4a+/IGAThZ6fkJx2/G48+pBAe0nj
ENwaeVO26DZwX9Ht8JkCdBr5w+J60Q7VDiajFntld4QC5tQpI4fGvLS3mF2XIlNo
dy/bBgeqjXonVsMvQMtdKq6IZ8Y918WvzP9mHO/Raf4YU5JXIeyNfF5dnc0XGfHu
tWcnh1JUN+MUgeWCRc7PVgI/veqK4i+umnvOt6ImWXfOg5Mw/a4jblrNU3eQwI8S
O0gFobTBa7HmxXLtgx5WFw/GdmL3X9NRkYRz4+2LSpQU1h6ZYnLKncx3q5Hxx+OJ
UwC3yXR8TaVId+4wXIVObebLeEPCGHB3Ue48Y6/RyisKlre00dLZHDUnYnRYxLnY
PU61bbP0EgSkHZcAz+2abI2emYvnTg/l+QBOTrGrN2BPEfujl0yl32FciOxsN/KX
iDgAmZ0wEgC7sRztg3+A3CGTjM3b95IaETrh8/E1RHnisN7RQ54T8op3uEvAo7nw
U3zUILNwooxRiP/EY5/4LWHK4MIPz7jArT9qA/mQhNlHgXNdtxGtcOrZISS8RUYX
4HIemMxp8FSf1qvbzm0ycfFEo80jVJUiifYGK0FkrQZ681KDas1v1I6DXc32UsB6
aJXlsYUMubT34JdWO5WKeYg/MsK1x/zKpkmzL6qJNGIaH9ZvQvKlweeIXo+BmHNR
Ttk6q/2bmReFT6UVEDlIEejTRhxD2MehcnKvRylMjKlFoEPha4QAb3eZWAfrXngr
`pragma protect end_protected
