// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:33:01 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
eDZBXzLOeSDPvRCNaYPkSDTYf5hOWezYQ7WudvhyACEo2ZT8ZK8bY7j9mx+G4I7l
KfC/IfrrCpRun/pjmd2BXJIJHj7jaxABJiGe0oKZu1I7ndiuVOYNRn1UKVCMO3Qz
6JfV+BkbHHaFtp5/3H3+16wQhPlbXLyEIR64O8NkN3A=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 16576)
Z3cJNkKHHNkg+18vQrussaB0L7PgIhjboyGYEfILcwc7PzvXj2JKEnd66Uy2a4F8
x1EHs9JLIa5ROYkVZJSEFDcg7TXozQx1wSlLtZHdBUHLd4Y8N8JMZ+JbPkPlR44y
mqovu1vl9KG3b+N7aPWbNmXA4zpEdq8MGgUipx7V6Ujldbl2M68dyQ433qZ4bAhO
mDqlDKV+7xswueM+/K57KFOcckmCxNSVAPwTDsv9hEOmJTLNLggIq7cOJgHTrrn5
gVBOoNqr8hGWqNJcdghyBxcJpFSbCQtErJywU7Ok2bbv3F3WgMms5LYWW3vsRpKk
bGnnyAYTseHQejOpQnh2H/m2CxMUVEYGc7RHIUg5VKNQtGtYRUzG6pDRBGOJKG+y
Hto3Mpx+rPINlIKXTu2I4M+LFpObRV9xX2rfxAbu4C16/V5GRsdVgn7cSJhdi1gi
3+F18BPxm89E+06mAdXBbBtYtjVPaQrv7uQkl//pOqhQ0HQ3aA01XMWAd5LigzlN
1+v9/N8ktdxO5mhSYYJbh+Lvz9hUMIcFgIwmL1+OxIJwbBn5ZKPrbQuXq4cAHFWB
gW6gkf/PP7yN2FsXuzvk3RzWC/ez8TBZyeIkvp3Q5dIzf7QldSY20EK+ziDoT+T7
NRu2GgBuaokuM/CCx29Bm7BMLSmdkL9Yj8uCr5U8L4kFRhzBWrPa5qoYYeF5iStG
J0bVzWJR8N+bWv5GgM9m4xySL09Sv5zcFk/Opf/beE1vkGa59jQuOEE1huCDyDb2
kQ7ZlMJaT86VoCL9GmbYbEMyj5pdSa91u+RnMIKQ9BI5mH1jG3rVM1OQSo9CeVQP
kd+IDS40BzGITTJyHGIF3RmHoYzjswmmBLU+mJH3m/Lsl61FMKtFvtw8n77jEdP3
vHSwlAiCxuJoI8ryE0HoxrpU7khFeYXcqsbOdaHXrp+d22AdWJtmS+wygEi6aPPz
f0Ih3bYi06WebgOUQHzAEn60cJRWwlcSShUPsSJFuVf47yB+34kVMkyDUYnBKW4Z
N1U4pf5bbFSeeTzVnRSGn2b0cONq4X4JtugIxy8WHhMMRZdAfOuri+YzMjqwLW6W
bznqKi1MPZKR5uCV+ef8MMLClVBYBpVUg44T5k/OXvj6R3JSbHYTw27La94WKqh+
rDPgryHDP3m+ElMvSKMFScfrowmuRm5A7jUQKnupigrhXmTPCxRWOyg6GEnZufb+
uhjo0uFBPjWTl/mUwm+9ro7zd0S8il8Fy9dWJLJrnrn7DxU2Fn5WnMRJ+5ydkN6+
EdAySwlajoLaNsZixcxjz7ieFXOvUwd3eDzkCI++tv/Ym52sLtWotgiKBDcthRYz
1PLnuBVYyS/4gu0yVihL5Ga+RKoj2R9ZpVznb5nKTJpmtmGAAif9YUDApfkkdQn9
ZR8EFzgyFajTGpt/L6rovHZhQ1QW9fc9rhwbKoQCpq1YUGqlL/YAgB3oSfPesCDe
CNCcKPb9N2/xs2Hbn6mnnrFR5a38skol1ea1LzVBJV4P8rmB1NMVH2kZmaCnLyAL
ngPiJhuCLMfNtvcovXVkiZ8VEI1SzlsB77krJXRMPwyJdLva3ElH97Z0D7uaYEGo
x2ItPYjXfMp1F1ZVdFYamZsazBlkGQDHjYnUnYFCMZwGDvL0Z5ioGl801WX7+/PZ
O1xS8QiwkrfSi68/2pu+0TFKuEppvKv8N1Vd5tBi8sYW1wUOVlDvSoDX+NDsP21H
ti6d3Rf/6wZqN6VogDlEwDxabedQlZwmYKdKqdlz+PriG0hK0nAjFa5Efov8Dfgy
0eVrVHKPQf+oaFpSNGoRKC/4Ff+pvYgXNofeThGeACsBin7LsFrX9aA8HDTLXelF
Qck/Tk/UXwGlJcfFgODJmHTBETgw1DkLdpMGy0Jw6BnhxSWI+R7a2TftoKo1aUKc
j9bHxANsWmIzTXsg8ZTpJdL25BC3MgUsV5Zc0NdZTkcPRUk/oXv6TgKsvDAxxoGh
iHvhw+UDr7i8q5CFwNipliWMzySROlmiquMP9YMRHBGvEetIzQRVcXtL+TrBGF2l
+zyzXJWUjydlsRlr1yVi9JV4lV6UpqCJ+LPudiheHuFaxT7Y48SGz2aX9CpyT2US
JdYt5pZDm4BYdDWiQ6gz7rQxNtUEsxqVZXIblb5h1LUJnjZpJMtt/PWDgwygCOUx
aO1POlmFuA01DDuYPJ7aGlQljTL8aFNfAV20PVD0jsbVxqt/wvJPmHOlmatBtm6T
TgDl7/LmGVfCpKk1CieAaAtrJn6emJYcPfcPjweObSqHc+QwADbKh8B4JE7CbTHp
QhfwyU2FZlJN3NNM69Wnn+9nDQrDlYMrbNH/Ma+P6vIuEMlta0TT9eUg6g/SgI71
3O7I9KCCpu4TJ1SNaTLr3rDcxujYoD7F3D7zzzDxbWe4oF4Cg4/LT+q3eCE4oqPK
8NHXengOHr3Li1YbxbOVt8RTyoKR6J0RRUz3MMRKCq0MWZXEwwadzgMM0p8FfmaN
NroaqLgvKe8336ulUm3KYXWQxVTLut42Wbo7Fdlvls9xB+GV7Yyy4RRm04HnHh3g
VQTRzti57FyS2tz98/BTetRmXCSLdA5O8BUWyhR9bVwG5lH258+B7wW9VbXO/zYk
QjWuWrcI0Tuu2QgH91bL/00wZxx8kblrbBN751Kl17qcL4JvYLiB0tWx8CEWMzk8
9k9hL72bzzzRwKgOhh9oTKyPf2Vi2BZl2IOEshgN/lHljzvWA6eKRzfylBGY+ehA
LC23fctzoZz9MmXr9GYYHaa8+Ajt3t5Dk+OgfLcHqlEB6HcKg/m8kxL4w2v3Fgq6
oXpBOHZzj6aWOTa6rIc4xFCWjEWtq1Tl2JZDJc04c/CntPRst+eTE40jHV9Y5LWU
KMY8lUjL9tE6K/gYmYkz2rXZKerBsLP3L9gCmYDSes4Mmh3X74Ean515nPyhFDLB
XnIwoOrDFU2AzShLiAaTTf7Zs/4oLxRKlIx3oxhevCx0Z2Q3EJPaEbZW8bWvXv4F
hVMV+9Lgt8aZgu2o59/GrfKqhIzHDBzh9LurhpIrGaiqwZ6mF0YJmeBTPlNlilj2
PI8ccgEYhuWRGSl7g9u9nGTlTujm2K8nGvNOSjLrT6u6eO0dlVfuCXRuGcxiBR1w
Bk8W7jAdRX7rucqPf6RNjrlzIjh+J+zr5IG4xz7WFuC+ED43JYQ36lIjC+EIMZ9a
XtTpiN1F3nSajQqfA6xj7ZcyJM2Y6asReJGxYDbWNiV4h8MnD1yXPNgryQsG/Hx7
SxVkCsloCRIc8S6IN7bMbTO1+n1QNJIYD78hgeYsKewYLkCoaqzLKTmWGwqevFT+
qzG2Hcf6Tv3JT5BQjLtFvM9ONsDdvFttcdtgtElzY5vcCCJrpJUkGd3KYdfLyzzS
9bZ7Ptyw86FrQsuYaJ0zAxAez343u/qe+TiWMc5Balrscs1zKrZVvFLJ9reBom8h
S+H4F4T7OQxMbyTOcPxiPW/RZZ38osuP78tporVraNkqdrSo9GYAgZ4je/BGEmvD
sk/sZ/lniv1/EaH3TXLafBFS8QVmQAs350Wd8iWu97V3ZsFWu/TwJw5EXns+1/Nc
pHeiBLrSIIZKjqgxUulMTnD1u38fxP5hqL8uqhGedeu/JmbUahzsmKl0hmn90rMT
ProMsHJAgyXwzwyo2te1Ef+/l418Wr/TRNGHY/JOSZq/GxaAshwIYzjcJL/DvDjs
FDT63lrLASxKA7CpZv/pOhx6f+F3LzmI3EssSYHdUW56/tw09zOXR4/n+1aaFyy9
tE0WPVkN7Jhko+sJdM3He80iw+0Zyi+YKJSMnLv+bBx3x8JSGer0U4LXTvOK+OQ/
o5d+wcaWGFL7fZ4hD0JdJ5eJjJumF91D/mRael2wmrgnF8m6wapCwo8S9XMKM63M
rr2BpN82yhn6InLH3COsc7HZQESGfiztnXmYnjFeTlTZq1VS0LUz+2YwiRE0QM2E
5+Z4Ape44jIpmUmWpWJf1IL4tIARa0dG7/4q01ZWhCJpnlBywXvoRPi5gQzjZWtn
4k5t9KfCiwzEvk6lpj8i1s79tBBIEQlr8XIx8XO1Ro/RS+vgxadwUsZLmqvRgC92
tisxvPB5LFY41qDKqQJ37FISl6K0RTUJ8jivufT+TuxFtwv3eejaTyydPx2FiUfB
SQJCdLzcXodrH/gAvrbctudfzjQ/dCpypR8d0kHhl18WJmHyvn7jBS5D0+lwfCu+
KODbIQp8mB9JKB9c8U6GtzSLZHff3w6LZcJv0Usy1SGZO+oprW2PZLfi/MBHADTe
Pdte0kF5yZKH+S1PkHwGsrvoKEJ7b3H7X5OMYI7g24q7byHCI7H4LMRdHgOJAEtu
Uwv6hhl2+CJga2HT3IhLgVpuOD5ERWN3WB6Uk2QXuj+Aqp//e0MzPWT47ffNGsrj
nvPnZnqFMaMFebx2SEAa1n0vI2/frtAvTnBkKPuLoqwk6zZZmzE+BlGmQTEDPgn0
85Mf6MLSqqhvcCUxDtUluMz6UYetONc6xtEy13EqOa7YB4SSOLmnOqQ5bt0wnk6o
tKvi5CvG4WmDndv4YBq2F4SIVm7x6rJDG6FahhJ89XC627bkwGegOTglee3RrWZa
Y4fAJeeei2ztBNs36YOELihLOIC4gxHVH82vx4g96O4vAgC4b6R1vooRlgIAAThq
b5KmeOpK9+y/lP9AXtwIyY/OUbR9YyX2wGhaSBiVYM7PFT+b6W0oytX4mfDgFrpT
8VeXc5hzvTf35jtf2O2eX1qFX7QF0kgpfe2kjM6qhV5XbWapcmz2dOEzs2Y7kD8/
2Sc4ZA+LzZeFK5Q9gPqkFNYwQJPmuHzHEH8yyuxcP85O1ZYrQWVCWUAadPGZMGnw
rBtaWeEHZsY37t88Yd1cPE89wDRFXXvZTn0Zsm+v6GejqdYr9wVeMtZ+aCk22niL
hhop8OCMB8BjYBejRo9RV0uH+HibUDh4QXqsFoIn632UaJO8qOlrdY/73/EmQhAa
oTEJwjxCZx9z1Y2gv3Nj4Hcn2CKCZXy4noHkVtu6cSUAcW+Gt4GKmMBeCwLao6Ym
tUnV9iUSejxL9vd0hmg4vT+jZqbgcAWsa3xi6X+vY1cQds2ajb0CZzy/6a8bJleU
ej8QNKZP6801wchjclGQQPTcY6lYqySzYCKiY5yJM/8HtdToVQp5BZHn3qfqGrhR
yUZ0U725ppqVcdUp04HIJ0TDoSEjwrgYf8YnQ37204yUvvme+TaN5jLjhdFbnPvh
uqOL2G2cM1a16o763B9e0vGA3z0fSxhS3COy5EjppuJbu0hl2FtS2LXxE6sa51P1
OYa13loZgCU1KGRXnGb3NZ3C4sWc5wRCAzrTukcuP6t7XrZF1T6+xUTzffluqCU+
318twoIPCY/3XYzk4Ahju8BeFT9Ty+yFCiBVN11FVxRWEuveWzTAjpyc+9HE396I
xDlwxh8GXPA2P8NqgK5BpuZiqm8jvmYcmjCwCRZzZRRXiLLpJYYbCEsWqz+ZW+EO
djl9HvvYh7tn6U9zvaemSFrO62uFlyXYAREPAH36duh9CYUgmEC+FxiFtpqPZ6a/
PluIYTfRN/y8InBxks+9kvURL40a8iCq+PXDjUaRF9i7XjwxqlAOV6VWeRAULPGE
c+5L34nwfbsqi+UmLMO9De6lVJnVrrg/GdDP75tyEah9R3DrGnkVW7S+WdbP9ftJ
3OeZP+0Zxo7BsVgsWYrPccqVroALjBqXYQ8CL4eFGsBVIgInE03lCwHeysT22AkS
sNcLQBvjRKWW00PESkeyIYxqD3v1i+ZcvBsBy38djds0OdX3D9GuhtSgCavC71DY
Cp/EeMJ6tQplUYXqONvXmS7dSo7obZrnNg4jKPAxiRByF6erZeDi25ipsdckntal
JphoXKhigb99Rt1nvSpNSO0grpsWXLZYD2Ei8IbdZ3rT6M6+TwZmhdFFxvlZek4T
/f28zlhdRuNCHYIOq6ZJ07v0OIPEjWo99JeWhIC0MQIN4bI+Rzq1IDTClt2YDbBY
FGurcZW1SibiH4KWJr+5Ap9B/c270TLDxID/Ct5zJnpnW41f/EtJgGvfDUKS69dq
w5c6BbGUqvAaBpjY4ksyhzCHib+3JgJfIoQ/NdPyj4rHzEY2AqXXuub96g+u98AV
UBNK78i/KA04nx0yYe3Lh0aiO66uYBilymLaYlPzZZaqtskOd1yB1AapJx1szuBr
6UU+KUgfjjif9iFLmfO5efq6Lpx0KD5yYqIPTZMH1zv9+cGP6BdTGYosHF0D5h4I
gZ4JYqTCOihDheTqDUJBAhINhEIqvzjhIi5Zfl5sOSg3xy0P9tL1z8V7/TpdVkFs
wZogh0+kXikizNgfOSO+vcFkGw5+s7bgyu5VicKR/5Xvk4mtAFUDqjAE+anUi5u/
WCymW9FGwa/2Up8LWH0+9uL2V0SKCHX9cA4K1tRm9MLF6L6eHa7G80yFhE/aLe4+
W50oOZq5I8e0Qz+5OaXUrtD/6xOM7wlH9PgaXbKD3+k+3zrC1jPuHT0bqhcTy/UD
8cB3/hIMjnf0cbLMQ1Mo6UENweLpd9PN7lh3ptzckbrCEjMjAfc4Bfe7cyBNv4+K
skAt67XpgPxIH/RAYJAQ3VD/4GnP88FVmYUrjbKH/ur+fdLfAqROgh32SsFfVc/0
JWkSqPRkPTILX2A1N82hEM9cGVryzFgQLqHIgQRpv5AH+AKUGEppvEQYV/1Mfjat
72XiQfUJ4wzyofUN+iA+6F/EYYh0v9LM4+cbxcMP0glyjXDNdwmf1uEe+AovPEYN
Y0Z/3lJiLnEAS5LK++Bg40nhiN6YagKfaCBBpA+qi6Ljbi+jhpwvVovKp3kwrznN
Rnu/bgZDjRRfMOtTgVoZFF1LkzP9E7X90lg7nitsZqoUmKYU1dCHEGIWF4Dsj4g9
68GqvSQvJGdEkDJdir+whHOJKUfjMa6ZcstyW5blEXa8E2Lc4bI1YThCbEAkrZbe
oo/kdmSidhmQBJ7jwc7c0P4sEkbVDUT6InJB6MrbhVNyTxuDXhAEdZ5Ska99tqks
RE3HaUFVsCB+fVgspOkss9futgSkvVmuF5oH6eRxfRU0hn/D9XWXcfOJPGqCRuMb
OoybA9siPLvqkpvsbp97TDKwzveTvfPJ9SNLvJHVxDPRupjjxZ69LzH3R4rh71UM
PCJWvKF/hsA30c9pFt+VljWsxp2+EXIJajFTYRxdd7wKxKCqWJwDBEQ8vyklSnzp
GN4ifOk5YW2trzg5FIa3yxazPz+0515vCHTbXdX1QcUq1TE7IPqkx81thyKhi6Vn
fIvimJqrkeRO4pGjOcNKSmRBfxtgfc56d8BHjTZ7XKTP8wmAe9z/tXpy7rM+hM4q
J3SK848wb7d6YtQvt5jwREWu0B2I5wHEhCoUr50r297Lv9Gmvu7nfguxK91Dgo+J
5rC5TDC51IR4NOvl5TsHwrSXQXW4Kqk6dRNrmW7D0TMbF8xj+QjjlJgeTZvV9xTj
KvnfMBhgyeAoDdL09MfXIoDdGuEjt6SSvIW5zMNGoaREGRqIYeaSZ7/nIlMLkqlA
5r/oULHES0/8yOrvPyGkeNcJoGcnxzwiMajS4ld6MegIRUjQH8Ubqhlvt6Ae+uQS
7IpVI5tjIvpL9ZjE5aCZ8GB/h3JMahl07bqL0mPzLrCQmfd1h/yHpzLYclOkIUwS
/khGupzma24L0a5jzDuDN4QeVKZKMu2PqY9ncRA2RtCEWtOFpUGqx+sGi67N04Og
T2aJLbd7zwavSXzqsTSI0VkoCHG5r+TWhQ8gAXfp3UD7Q7r3zBVWyJkSrN+89v8o
WlGtdrrSetYPLGresrtG2OBb6B5h92uFsgTG/K55ts2GE2p55T/XModDI408evo4
gHsWt0vYRsZRiFZS0mnv7zjmcWobOfCU8jKb/86k5OhG38mWJXWYx7EUPNoFtFlu
DDFB97PxSMgiEFcuJNkYl9anLE4PL8pqtOAp3W0FSSejcFfn8vA61msA/9sV87oj
kvSIFUIGd91VnBV5U10cRMZS5zH59KKavDol9Yulxm7uRnrbuMv0s3qmDC3VGvGn
9FXB8Mc1EaXyj30OJJpUgFVDSBvmbVLQEa50IWvT7FXgEAqarZtN9gU136l7qOmp
IMr/OyHB2Q79DnYOYJWW4byhl/yE/d6Tsqj3u3VmTgIq1r2OLnp8QVan2KxnfoI5
M4QP35tYtBoKJqIfw8c1nmeCrV7r2dh/gJ43RYtiG9gklpp7j5NCWvwilGWyl91O
VyxBneg69QI1fTpiUXarE0aRToz/yb3yL03b0vFUDysbQ4sE3q3tIMJiICOqBqBV
4YdkaKb/kt0mzmTfHZ/sRCRKQQw75ehKYLTdGDKEltDBKlBE0c/UaO9NEdA8uAxK
97FOZ6QJrj2unxr82PVBIgFuT7Dyd6KH2rm/TMzmVOZPuFgXKa2BeubKsLQqr7Pu
103cJAQ2vx/XZnoErH/UPY1vRQ2DTVpSCSkMgsMjBU/dczedS/0ZsD8GKOcTJLFY
pi7ZF0TCVRZMp1sijmAYfQgk5gHU1nriuu2x0XbYKsD4ImK99/WawiTchqrEC3up
7IjQABazO88oUmGYqMWkDUrYlYCXjczoRz+5W+XTdkeZaYU4kQDmy26eUxDR2Rql
Bvsk0bMp68FgXTAJUtjScIUsrUinv6w/o+joDTd885q9l5HQvSJ3wTRDc/QBL0Kh
fjYBoRmrHVnxexFwifjI9PQ10fqbzot3eqB85/YSyq04ivVP6DlNJDYOfTzzMKgj
kY9xwKFRe3bEm+q0Qm6Q4j/V88OOhCPk5Z1e5JGHuSrflCHkxqJyeaYBhGm+dVaG
RiAe8lRuiGDrbReVHG7eT3nMe0y0t8myAJfECoBFzRqJYH85h1s3/wVi5WuS146B
Cr4a70DUIsQdZJjE8khJP85X8JXRsLaokAliHmh3/HAFp4P5AzsKzsz643VUgiXl
gH3Xk70iNEahYffHSKhHK8Lz7gsaWKTxjlXqJIVHzZFqNwOR90UBpOErvT3v62/r
cRYtkjNnCMwgpK+qBXbTkwdlm/m136+0L4qlFmHQAqBEoujWLu9RSbULZ5rKTzn6
2AjuO4N2opPhdvDmi0/4y4YEgbrmt6RMih7yCY2aaUsTPfW1pTUcbjFic7Zh1zGt
C2j1HlUD/W7776VGPCIUBX7qg+cmHJQXEd6QISHKT4rc2TaYjor4axEqJWdt+uKv
IeKAqeH09ESONnftmvWn2AR5i7eMrkFmSDuq446opip6oi5jBV2WVhXwufnf4D4X
PNQnnpUkbH+lYaZkYss0MniqZDRj3qzsQhNsSaJvXXYdxfKNzyOsuRe9NHbBATJN
C0SWoN1iC97MPAShfuuAoudCYyTkt8nH4sGtonUwbLA38yYu9rjUHQ7739uyhxhz
jGcJl45Fr84y4XeeBq6HntwrwzBhKtK/zDNF35LUrAI4NazAZAX4FSn83XMeMJHa
8AxglRmIyRmSlT5JgnNybe6Q6ouQifq9MPCiF30utwyNb44BcEpN5619E8Foq4Gm
eGJP4umrl6M1vetfEw1Qs5ln/cVr4bEVKHoSg5hVwuktzNLW5jnaBRlM2lo71rrC
oGr29i+tXzyX8tzSKFzipAAQHSv/QmXbw10pbbUd63m9fqe7G0VsZfSF7WiIoC2H
b5xpXUGl/gcHygUjttQUPmfkoOngjLw9YTavp/Hki/gHN3edCwBZS8lp0fzLDKTK
hGnQNU26Bd0UvmGxbjsOYteHv+SS8xS6ds/7MxU6fKxJPKAibXgNO70y7QNyc7Er
1t/WxRFtrFIwhH50oQbzXisR5f7pJ/P3ZwL5UPH9997snDcu/rvQ+zPjBdrd395h
xKDJ4ulJxoxyGoQe7OFaujIfpcC9obO3s81DzAdzXySn8rO5shaFNeQE3ucPAaSB
qzBsWDEKA0ex6XM0kj+878xATQ+2wD7PhTJ1kXaOq2k+2TtCa5T8CMIRRhemXR1d
2KFUbPpijmVFLWtiLORFAF3V1baEJHoh+wmcGZPy5hy1hrpXndkXU3bVOCaaud4Q
PT5xyNuIcflKWR8XMKRSACujfrxxV1RztZTSRaXHpPow+pBq38lp4ZLC4swwesh4
IBRv53wXf/Xddv9TOFBO0Od3JnvFaE5mjoQ5KtJKNT+Tuz4E7+60vq41az28DuXf
ocWgezdWeUC4WtvT46G1JBZ8WkI7LvdNOkjsxygHYfhrQkBP+1CsYLRwSqK1XpXN
jtaxznNt3tGaD0fFQ/frcxtVKRA7h4x27f/JcTDtf5pnl2coVr6NHWYlAE9euMXm
CCS6W3+Wbm1/IuyuU+IW2TNnEzY4eXCMdb4/DeUUQuYrTHqccA18+NJf5k0OPd+D
D03ps6DIOjSuTo1Utwrh02Y6Mk3SNWANRSphoWxSGyxc94zZydNkR83qyJyi5mWI
PnLHph4PC4GNRPOeTgzi1YhXwbrs03alrdbg6A2Zsj5wtDWnev4ZQrfp9Q9LTKhg
lK6F25o2naY1jCyma9MFTZnOPtpLbZunXp7JuJb9EWQt+NekQXVLYDxeqsqYyN1E
mfx0nbZrDam5PIZ98QCriw4Ds4q47KPRyFuQYUe69VwvC2lmb+WBv4oQHQy2wMCy
UW3ETLW1GBGtEiHYprwzEPoT8m3HC9m8Rl6dcREyljUEK7zBmNGUnMu46tqAJ0m5
1qqY9mdiw8RYoulj11FGfkedjKNk3QFRA6XBEFO/yHSG7XO20VcVHsMoArIzoj3X
hI/dmeb27ATCcb2lFleDJo9wq4rsEVOh30XmYrktvjiOhUSxN55j9kX0tqGr+5UA
/8aDm6rvCY9NXAI5y7780SlBbzDI/WdyaJo7A7aLcg5vTQidfJX9akmxG6I7e3DD
9O9Gge4c+HYX9RkOqz5tsh02cuNn3CeNeJPbPwfwL0SeQu5HYk/pj6kFXQSV+0eD
FbTY1lA3Z6bsIjxB9zNztWnlSz30lhL9cCPKx5XdSo9FMmQpeAgzuhRHYgLp1YY9
vw46CHTd1k7JsdPDi7uJITM+q/a3k/Ka/JtoSU9htEFY3aU1tDWpM8pOugvW6WJR
LJp39dir05pBmCgW5KHtxcdD964ooNOTZcQLlNihvdIVscheAu4pwAutCjkbS9tZ
e/NP+GPd02s9FS9jjlS1xfAuiPa+pBVfjW3nzujejULKQTRDShCJAx3c0p9THiZC
8lmDvCZpMZIK8QkhHTq3CQHoJ5ZKxKOhST85WmnWr1SfuUu3+3jtNZPd1T1kp1dF
kPwH8ILGmCxw1e2cczmfYp9beGRBCwDwMf/vQYZIuTmihapyQ+jcbQjxySwcPdvY
E/NnZnEtDN0m2YKMTb3x4cJDfPml04QYx3elmPI6tK2GEo7xnkwJxu6dxtiCnozy
Pc/uI1DHVysmm7gnheAWZZAC6ZVXbnzHgXwmXCNieTkLNlcGRPeHu7Y4G2kPJ4Es
c/Fon8Nvl1GEwU0RL0QnUiDhSSdHid+afHQOjnVwmL2Ac3KipwPXNsUlc0Abb6RG
88hBt5spDho3KobnZTSp3Zf9/3JKlCherB9/Xna4BCpwib7Y3t0RoiYEFunqUF9L
xxa2pN2R4P4qm/l6wPk26FIdnwvk4wRzbcLFHZXVrmPMXyi5xEaww5QSgIRbpMol
BgxZKIhmEjoUEdO2HIcm4GncB3l41H3vYExnWkQjfNNlqP0hmWw9hZ3Ro2EyEQlb
59hYPkpMDQXyTyPsB/DtJJZkRIjghzcmUtC3OmR+FtqMpDNM4kDYjA2rc0V2EAlT
TEUSAlqjKI2+EPCh2Bp8FOAoJUPyz4RYuD+I5gkiRRsqty5FO33GAIb/IKY6I+Hi
B34y3dHBr6fzDTRkE7SGyBxg2wuiq6EtdytvNn3mi088IofyEXVVeroWwJaJpdZf
kg/tCMme0wgGCcdDpoGb7KcykreI7+hZeeIE09b1Xk47hy/MXvwEvcc318jI6h4W
wUsv1CtN1miPIX4w2FnFuNpuroZBx25aGpWt0A59nmWuq/UiqXGZ78w3qYeR1DQv
9KkN+nxsbqnnU5GCdpc3/hJ9apohSc/c8TlGicdsu12oSiX0abLnrdn7zwbIwoYz
KAsbQhE1SaCvHAu8s3geAHBYm7mvw9Ph/73S/WXoaM26ve6fj5ePNYWnOLHvgpP7
iWID0/TelmKtIgTtQwbjaaiBdTYHuYrYnD0afLPMu1M2ktmiBwyDmmO4Da8/yGyV
EUCLEDtg37463moduoZXTx/spmbtuBaiy57J6TX9aIap4gY71OAGZmNLHINT80wP
zzRAnLQSy6ZdsY4ggDlGyxI/+ZjIxhbajacTexyLjpH3bHhcZbXxOn4yRY1dXqH1
CEyWlekOug5rjgnc8ij1YGYT+gAdqcFu/c9fvAWqSSvIvOEJSOhngNYWcMds8uSX
poWgVvZZO8z0rgLUPFvrkJfRQaxhhfOeWTFF8swXM851xTRtoLv8hFrVxpiUK+0I
e5BMbJ4U7qpRlMcfQmO+fOc5KPyxkkZivXbeJ5lvlfHXZ5M5lMa6puwPwzuLLsfP
oUtBup15a8zwE//hqFLawpu6N2/QO+FZiI8GgfN+ZY74M/KcJHgrx3ocDKVdClXk
+eNxtXfwkvH8IWLJs01lrvIOBRPut/13FIHyueorTLKhZUhT/ZuN5WClS9gS7N1C
3kjjsEEel3Al5rwvpXEG4yENmUlSQWHjrvsHrJUA7MzeTF2R4IOrA/Vz3j6R2YtB
YqsIm85jAjIt/9UASjWSddtSWJJVgTlEiouwc+KlR3qlOuAFSV5clbTt3Emf5fcc
SMCL7n6E+HNXh/6eQW0iP0RPBqcK0pJdwe9N1R5yBWtmp6p8FJ2GC5fjFquN4NyB
1cHYcRY9/rWN+S2omwHXHo5r951MDOiTUNZJPVW3MiVys/WysU3I/IRuinmabBY6
aQgvUtIspwRiVcR3q0FFBHo4DPrnnMVG8PGy6vB+g801uz6M/M/RPXsWL7WVyIVl
ZwrXhMtCKVYKaHlb1/R3ymoLTkRR53UbyQQA2lti2aK78PjmCFf6pAJJM4S+AcOZ
8ao2/sniYgksYs5mJFOqvseSu+whI4Ny6Dk7qQst7lWeosUlHE/AjnPE9nO3bmiO
kWCtpExub1dUZACCcDs2BnxFTsw96LHkRgFUa2NVQFsy91f5WDguTA4UdvnHbPY2
sB0AowXWEH5wmn+mEqs5TP6Jqd1kBetnZbOEcFrDk17fNuPDltg8uhcjZmkdR1EF
EblMIST4V/d4zdWjZcVE13ATIiZEPgvPxIIwuarMReFB4Fmdqoh3pHwz4aWyceYH
+qvy3wbePwQADavZ4EytruTzxYkuVvjM6EnOYdmdOeETSMGqxuVTPgoZpvrwGNMd
ePY9LCd3FgStmFhNvxjtivfi6un4Ng74uelvOxk4yQtTP66V+6t1IHMfHxAhRqp/
Jw71Js08mmgDggVkuxtPLoIg2brLQn/wBX+oKpIegSIGVC4s0C/IdfV1rEKZ48Yy
f3YrUiSvvV6XNvYjQVLDp5orHiFOmyyNbRfBYSUDxVPdgOIqSzXjhITttktf4OlL
PK9xkYyBRzfSkv0LDXCowYheIywK+Xoy4hJgh5fszGreqRrVgelX1JWm1LcETOp4
6c/iAYJFrxmfkNdUKM6De0oKAqtmYGv6Su75YAs9rf5KLORNYfuMy9yvTADyvg+J
236j+o2lnUxudSz6KyJ8RFDneS8GYO/cWHzxOE8cl0pfe2LxsK8ZYXIkOgXHsLos
/UPKuLQlciW3HLLVihqT0YdnAA95m5dTK6JpablZwsDNq+vrIq/3lSd5yLQEyZYw
ygRpu0u9NuchsJR6miPoEvJfYtjoBM6X7FxtBXaPB8gS735wdM6JKnn83A5jZs7L
QTip82lD1UQvoorTwe6kK4LCdxFNpIHQ2HQN6vuxQSNGecdNhh9gLeVscfiizGDD
DfsK7UYd3qGs2j4YEY83sr/+O2zZ0j6EdhaxVw0++mh/A0K+vwFyQw+w6nwLNvDm
OpacJPKPlT34wa88GpuO2YL1U7ksf9fML77Z82iSzCPZ/K6yphFi7syTERHDGy5X
jDYwqGdYZ66ayokXYjqgheHLxBtIZpxptMr9pIQGPmWg7kkdL2ZV/BeY8rXqO/aX
Bp0BRqmDAwunkNNzkM32hBmPusMgA77TYKeBcfGBHbENYxEXx4C2KzBeNm8Gz9oN
kWFFaWDLn33sSzMsID30kNOVP5L+7u+7kMAbD016XxCCchEm6RHr2yFpjq3cuHQ1
bb3WbLQjBjYY2N3q1cCjqJ7sDz5Bh5/Tfus6C2ZALFPwCTqe+JtvxbnnJ0bSw0wH
lR4zbnvmLiKwCeeqnCqbovS89+HuZWrPm1wVIroTOzxPiTccgG/P4edaMHuHJbkI
VFGskvuJ4d2KZXVAW+1Lu+Cw5x9l3Dec1akwbb1Lowpw2uiHvZIpMeygdOB0QUPc
ry9EoXs9Kev1HZ5UxJtD381TyRlZ5iGQimxYbdtFNK9OJy1OBvhJiIjQYP+AAeqq
TtL6BMFRcAtaErpREFvYRO+yT3YoVcp6au61edLiy1elwjAj6QgXyeid/PySJ31b
dS526eyczEOkQt8aULlLSNpRNzPr7YADCcWjOmpCALqrlP0BKy7lKaFWCSnUXoH0
9tlCNMH6hwFs58rNjPz78jhoTSOgHIk9liG0auPQb9/5o0us4tvt7IJrCWJn1y/T
nCGBQYWZF1+q3lFiX45+YRIoE7Gjr5d2FEd2q/cVYTgmfl5/JR+m8yiCj7Odzjs2
VgJyG4OngRetLjk5GooezGyk8W58wEJQiMCYBAgZjQCzm9hIq+wvdqAXRFQamUOJ
nwSMq9cQIenASosT/GGRiAYJeKsVbSnItYMeM/w9TSSMmRZUZzwXjiX8sx3yXSml
PRio1LcO8cp5jMzvJK/lzGcE9iTQt0CUAA8wES3vQ7PcT0WZ4tAHPJNEmXyYJOoT
RXy8h0wIFtLpISsKkzOAMPLfF2KC/khYjaAxzl2K88BypQDRnxcTAVOPbDB+35R8
2TGOu2JtAlb9md1mQgDYg030L5x6uvxU+LxkNjLJTsbw0Dgwu5tTMe4SSIQGZ5cg
+DfeGYuXicyVv/ZaltIbK4poclO6kvZklm9D4bDpL4Be0YHUQoJBVAvRgkEKeoZ7
xpjZ+X4vb+fu08czU3ilkZ6B6AJjp2eapoGaCJ873/i0UOrWsp+CLylyc1v2oo1p
HMTsKjMLPCmsYYIYfQ+f1wkJYZ6RaNxtSxtiOCEEW2UgStP9YEEVzqK3DJ7atgH0
0tKMWVTlqJikD12BcfYJ49wJSwJiM+MQpbqg60ITFfH8jQVc+9/7ljWDiJAQSJTc
PCjbQamNwdVYRK7fL+RL040eDVoMQHnNChnmjF3lMOeah6LaUtyrYeOQSzTEbkZt
/IpsydOgGz+n1/NuSyw5MZpQe9I4ANnO7ZjjVFSS26/G51UAxAD4ezcyQUbCTImj
W7amorYSEZ6LNVz+3Dthix0Mfh2G6vgGwjC1Oeer1OedLEmMu5QhPrDEd7Pc3bA+
mBKg3FIF+mL8INEAMKwVUG1DacYHwxTAdb+d7NwA4X2zQ07qR+NVFiH4JOxzBDYn
dsP/EB8NTe7DlgXInLNMdmQOsvP+0acKh5UfTA2zsePYXs4c/9mPwSJwS7KGPXn3
cNjY6knay/9DhS2wT8Iqu0N8N/4qxX0yNa3rUniBYqZsBCZyF4adx8X8/e78NPSC
eN7+Zy3ItCthJldkV5Z/wFi2qSogr2U5tqPlcoqQCwvk5Re7fvYY5VsNjmakImRb
E0Wo1KusfHA3AAUhogU4tiMTdpNVdxz3Bv7N2ZB1U4UXVoXRzywW9edqV/W+DMCC
ZFObue5qRX+XsTemmbbS5DcGavIbSvOmhFO6Zsz36v1NlYee8dTrhhzfqLt3P39b
wWB7ZSUZ3CuMwvqp6EyFUAIVZGGwfN/VlKEWiwXPG0tNgqMliCyT/O+si1kEltc+
8yAGSwlgwXsp4ea4tmRm8occkTfENOe/Pj1Zz+7qd3kJR57VO1Lucd2jMsZcKM+B
RlVYr4GuBoXpYHJ3tvI0BhPqujl8OO5SuLXRkEyglbPh/o44cV9Xve0mJ/EipJp+
prKSHQKQ1CQ7GiDy88TMyOPEUayBla0iBHclPgue1qFWgBvwJT7eP+XDjKAMINXL
XvSBQm7QP8Gs8tIfyjhpwbG7emqEn3DWmgpmCnNO95qAi3wjg901Cls0Ug8+XDwY
gMav9sjprgIh1TxC+ZMxmQH0pi/fvA32R3GdOuqvAjbEkLbcSo3mAk8sCZEzn4A9
ETqoK5jc64eHeTdlt4W48saSf5SLdqGJCkB7LfP3DR5TXjzSrWCE1kQoBHIIqIoq
KpUE9R+4I3xlkH6HX5pZY0NnjHaDyQVEYMPviRNaadx6k2LkVJthor+7udLpQKe+
m6olhkrZrnVQHmXQkmzv8cEZN63eO6hmHCdOeS2rSIlidmBw/fnOuPcYh1tYkwcS
DtGiCgZ3CkTQjiJQHYC6Wj/1Lg8+aCwr3yFnUDXbp1W1wZKX0MJ1d22nGJjWSH7E
NGjCkXo6zcE20GdRMVpLV7f7BkLqk1wVap5AQdJ1i2wl7wpn4NNZ7GGwmC0PvCu0
xh8Coi9uKxwzlFEVOLyMVc8lIZeig/Q2jo5g3du++3lqMXIJ+VARfyqYgFDhCi1V
C4WJDZS6SOpegLe+vk8S45ggmMk9Wf/KCQp5CQb00yjQrv8O2SU39YUUCzPH90GH
Wvj8UlZUhOiQV1an6rbcn/ARkPeFqXY5LcZXIeMwkHVKhY8gNCFrkcYLwxiT/Z0W
ycPVosSn6mLGDhgcQFh0wOWK6jm9mHrq14F7quuOYxSC8cChqJQMOwdxTmhoY+Fh
TLdbBuJAawuj4NRPWQA/6t4DtgnIzl9GNN/Osm45QUohffdrSRJZe28ZkgaKTZHF
1x3c6KsNxOAxIBrB5CE0A1z0WDdbEICA253LIN75uXpan6wcSPR6Bqf0eNehw04a
n7yQn6HqOTGgnKBONmvWZLTntAzGa7HYzEsCpL7obBpuYoVwQG5o7YTfLv0ha7Mc
aHC4G2A3/0N9Z9Cxk/LTDAUrUiW2cmocT7bZ7QTLv50eIo0gsbtlI+LHuAPyAnFg
PEK4/FKecu0jpnMAVJAGXILYxwhf62m/Sm6DglMXQM/0vMndBFVBX31cGvHhRk4g
996O2gDEFoC0uHuhZgIeJCnEU0pOkd1cz/UQKQVDMP4EVj/oNpTeQDOxIr1L0mTm
VksgMVbuID09smHnt+l0SBBaYeIupkJy/nm7E/FnIohG+6ZvA9P0CGIUtgm+NMEQ
q1XubE048pNNdQiBEiuxAlWZ1VdSk6JSTKW6mUvoDoQWjpRM5I0N5rmZYCsmXvnS
M4zkDgxuQ7CdCDnHo0XW9gSNTVH/23iFL7F0tWwnRTN+6yfwwe3Mr8NcI0fGsuX0
1RZhgrZg/YnT11S4up0xfK42QbgzHtyvs44TsJcYS9O7SRCFT5ZB16XgiTEvLz9h
z6jRXJpQktEuAWHbTpGIh0Yt+M5kE/Unak7P4fEmWLDbzqE1DKt3arWcEj1uc8q6
cVP5HRJzSGkPjJWrNc9VR2PWMxupkxi9D+Y+qA4Gb3Qh56ilURasfcBAVNC+DnTC
csWHFBxBIR8JimCtx9C5il0Ys6yhGy12aXmdLSbefY4GNS7Ct72bXbHeJPbS74id
oNinBAABZkiW39z/O36kUW2ja/bP4QvgtJvlDerGic6W+AeS4FYBIzuaq2zOtM42
5uqnRJDUYQLEnOcNZvTwnw4GMpQgHmYmNmE7U4WImTR1CXUVvZVzrLe7FW2tiHkU
fBh7/B3gvcKjxiqZ22+kjOKSnHtu/nGnK10TJIZjFCle4uAtaVGWmp0b9waTYQC5
GS2UDsjdNO2UdJw0VMnK8be4t9j+jQNlwS4c8FaDimEP0vDdO2atXRf7hqI68Dfl
4NfJnOy24qZl6NuW5sEHIViRLNaYKsTjFG9eeU6uQZwxiG274aqrOlzNNsVrsEpK
7ytWFMskzXS2dUgwkpIXbXAY2AgY2hU6O3kDF8gMEe70WVPj1IzhDmgr4HJ9/wGx
imrVO0FVhSS3y79WjHOgUEKSsNroBNn+JB8GIJugXs0/Ptm/4qq9qByY7UAZo/r7
7pySbNaYMFrm0A5mTiXHXQnDzfz5jzoZzPSKUdMRb1E8mjSfShkujp7dUoMhVAjq
9hQBriOAQq9kGdd5APtck7aFVmSXgHmuNr8Yz4MtXk0ZADdc+NZsNVBXf3xtXWxm
MjuzpTx1qd3SmcsZOs5A5b5f9Iwp9iIol6QWNKB9tEQ1fAIIv1YcM96d0tt8N1XU
Awnp5N6aPn3fN48jLz33dSdAuH4f7uWmL9SUy3AIQppzjLiXJuvmbr1cQ7Ap1HUf
Iq6PLnf1LPnnFH8OS9P3fM14k12WgAWJzDQFQtDu7JMENpRvcb1GnLfuIUxW3WrU
L1p5N29os0Bs5imipGYJOw7kBYLHJsjU2GaC5rCl0YkoVRplIEvs9jHzAg99yiE1
uPwgzhAuf4CKIx3noCAo/aaQru/OvwwN4Bm0Ydtn2uigW15jE586Z/6DBaOJY03x
QCCGvV9qICpM84kqQlJrJKCaUDN8txZTAKGA3LMRf2XnIWP/fbmCbzRKMJknRfJS
+sjUsrQ+7kcu8c+3o1jgUALrpkIXLroErZFjkEmuE2br4gNv81iKe7Rjemz+srWs
J2muWqcVj7aKHZ/xneSXRZI2hJkPnD9ptHE0oD7UhKB7wuH4bY5rpI/ckuvoRGtj
Ir28thGWC64FtWld8LIvU0rd0a4Y2t9JOHReKdYA1zMCQD9DfzVnhnLHIcy7KZP1
RNvzzN7C6k5xPdtO5oeWZwz1+E5WTXg6mtnfDg4PGE73F8NDHDAWu2JaUrz3L5Qk
dFg8B2Osiu/QyBhwLxXvCouTBMdedHRABbIcZyY5P+aOzfl3jC6URmZZJUv6Zd6F
Z8cFPa+uHZcVqS0LtP77ARzXLhdEqeXRZXp1L9dDvq2hSwSztXGrcR5xiGKxogZS
5/ox0Q7gZGQ1ODqg5z9pvuhfXlLLHok1yQtOhvYgLTJOlgkF08Wo/7Vl7ffSS9Xh
D8t3/klUwZetLb/eIIKVxNkJnvzBEP1SGa01HM3zSD09hbgm7xYgQXhJgGB+2uTb
drz3DKA5J3VBg/Ej8doMaj2sJdk6K2H6TI9/nvJOgA8WyEiJXCrIsvWAU0bJU9b3
etCHsA0QTrTRISV73m8n1lCHhfwDuWX8Htsf8VOeFJWhkzUG6z/uuyGzlG7quqzp
0yaN7HSb8wwfqeM0L//AnqIEXgSah3luDAS8l6C635L+L4+sx7bq3rJySI7qtw58
cmYjd+f39ZCDCj9QpJgP2MEKgcneOjyorc/KhV2DbzoewXaFLnlfK9dmbNopZl9X
/1m9F9VG0i4peicfGElrHiwwu/ggQbTeEHICW7NJmj1keugFWjRYdQm0HCCjwGE4
VQCd+bHpuGq2s/p99Z6dtYd9JN4BPWwGUrH8tZqwHMNAY5GCYdTKYgj9Iqru0Fky
0IB/Q9M3ql+x1Nx7Tqs+da9bH3WU8KsBqF/q0dK/rcKwcMvLB7p0Ld8yigChmyHd
bP5wl9FCsl+qrXifY4wfJKuN4LvF2295zGYnHpIjl9wRnFz08tc5S/VPPOjuvpYL
axoR3GZdm3eZylx6Z/dSmZDkt27olekuqB+fvQqqEqeTwIyU4i6oDyShbwI/eqrP
veuHKYLBezMycBZN0NjfDNYwOULaDS8r++M3S5yvnjldkWfF0jximf74foXtAh4i
InsrRu3/9/dQnhAhgOJI63pG1S07CpmrNqnpUQGcCp8Pury+UK7cpVyLrT5FwgDA
osIDG0oUevqrra39AmZ5Vn3dCFf3Ys0RwwAfJ8RjOn/0dxIkIcfiaUatzK5CE+Db
II+6I5gtczE36WYqhhS+EkQXS16/bsiwybu+ZSr7pCgOT/FMLYc+fqdMSO6K77ec
x+fOQO/ysrwOLslIjamjjjM+m1uwO9PVQd5s/zjOyJiVRfI/wgGpu1V7/1KRNnO1
D+7v77pkPlPsisLkd9dSwQnm8awtO4HXpsj9Bb0y96/JZbMNOS+mWugZDvBB1pHG
7kxk3EUoCh4lXbw0DEkEci2N0DKHUlKvxtq5zzLa4ADCP9sYa367RjNTesJvXPSo
kx345dUrWgjPTV4KJF8V296Rzt9zZhRkuDtlpzYiwRlIL6jtix4kPUsl2KwVkohF
vD4PZm/yvzNKBGCrcEx1uoYHFa/tz4yw5UquB5w5L4n7PfY41GqEAR8FHTgBnWse
gHeCf46MG9j0EhPvZf039gOXmy/Hrfa6szESHB6J2n9lqpOvlIVX7vRDUWuBmqR7
v441eVYVRWDYiNorvlteJlfxxERxkeAYhXXS9IFsI63pzjp4R3VRRyRVBZQKKaWn
1YDm3RThPsFBQLB7Y+SJV5R2qXlahXIptC16+A3Ego7BqrNqD3QRBqg0STSYT5Jw
pxWIbX0FBM5eLzoYMylrp7cvgc+NYBB3s9x4hHrATa+jA+i28h4LZoU8LNLaapWP
fBFHvB44mjizrkV2IET9c67cjnay/DffHuPg6xGnsZE/PS1i7s85eVVcagqPljwU
GfiFjSrve5oIIQbCjpqyWGaTvwK5i05pQ34VLcNc3MUn5T9xkjmIK4B7cbin3CDZ
EffA6hEiqYndeZh1aTlCYS2WTKQr79uXL+xZKjb8C5x5wdhAmxE29CNPVHopTC3x
1MN60Zs2wHC07rzKPXVIG1Yy0uFo6mVbDFHFSqCsHFa2QKPibdfuqJ1tfdmHqq3u
jKxX920d3xjowklGiH2hFbbo8PPNIpgFUOCWZbm7yYk6NQZnXPgIVOqp80ntYrx/
fhg0jCka0ecwXBViVdMHML6ef91WPN9JUtpCsAnKvzMwyDBMDuN4IGduyD94jx+E
YUe0IAJSIDT59DAJ+m5TRIvT8Zh5dvBwP+BO1Upy1RHNbOEk0n4CqLSUMxS3cQ2x
zH3rkP2p3udVI6ekPvmHKL/h0KPLLbY1nW4ETXtSN9z+vKEIRLwGVaUdpZ92A1pZ
dtATo1KhkLbZ3y4UdfPgfE6A34RY6q5RrA81xAPlw+B72tbR5eKNahq38aXKcKZT
/wk61wHvslvODFS5YdU2LCJXiORoH5wwu4ELOw7VInKv/MWY020Y7Qz6r2WpOj7a
TB9TEQWz7AT9T/Is8G2dwnQSFGhlIa5zzacqj+rpEVkriuOcTNGziVwerV61kZKu
G+KzmV0rhEb0LUJAqIUxK3+9HhmYeV1kd59/MvgE6qRgs+hdpDBwrnyGYKdzoGF6
9wbcvXVzFMXu3sz574Xa6rpRoFhYFfZavlTQo2nS5xmfchKM6Tq9vcV/c/9IqsEI
EJp700/YY7qdKhwENO+zBwXabwB9EsuHKpQc7ezLnYHo/H1DfkTYmyZ0JAPuz6Y2
LgM5aeeIfI9ZooKRhEA8KYwwVFZvu+IkxJY3CsBwJOvZ0yXFMKDkeFrQkG9wm9aU
XLuCUmjdsC8DsqN57Hh2Eqa91/tepxa63oc90uu9nrIa9wbWDyq1qVUaA4owOo/J
tWwjMWgHh3dycLjHuPG5rH5YvBn6u2HjbNLeSKeQaOUrknWIQiFg1SSmYWng4HRm
bI6YkwiZF5jsCCP+a/XW0yXpM5jiqK80aqQcXyyBC6Gao1t4SPvcvgLG06y1Sy5D
4fsuccJPvQEzh2rWEXg+Q9L4VmY8/jn4GHKH518hYtvchsvW7FuuTm7HtA5K3sie
FB6y4qrpxuTKugrANXkdIrOC/S+4lcH8kZUZNGSY/Oz07ITS2CDsUbplcY+wM5Ip
NEUsJemz/8SEqWul0nK+gcxBSgg1rz3XwBV4wEGrfbpcAyH2EFBCfU50lCBt3fpH
8MLfim0mPGjAUgqJ6VPm0nlLVJHbx2xxwFfT8oeD+M06S2Hn4HH5ROPsbzWxhGkt
ACfID6EEVAs2v+OX0QYo31QTOWVxBtN+Xwr6Dh0aGQs2yLkvQ0Kt5hR/Rgre7nM/
MpDzaM0V/Ya0/xNICvDUwA==
`pragma protect end_protected
