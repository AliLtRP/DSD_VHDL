// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:25 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
fWJ46/pY17K+r7pxH2G4E9pWCpheRSI8pVjXejx0gL6xe7zd3VWHh0y2m5urnl1p
n5v2VIvl3yN+AIu8VHS1LTi6BcP/5cxVR+W23cKNZFNmc+RsD0UwaY3qf4qBfuu+
ncTaRjWFNaB/KPnv33UdWYVyYg47I/mEGX3dWDngd2U=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 24304)
drr6Y/OezlgoRqzGNO7p71pabl8RP+edD795Gw8JMN/Jpj91JKhOyx9vOSuB672e
5yAeqjGbGuNgg+bCgO8/WwZu5zMzKBB8cZqmqGJ6+efjLG03qOltvdwqS6sTIMP1
DopvwUrNXDPNUaZ5lQ6JtCyTSX/CTNhHXJwOkRgT/JTBG9nphSwUX+ZvBd4GD860
heD3Z0ta9Dgl6ZG09Ljv9RNIKpjrZqKlFeAsUTfymcQpz/I9i2tIGk1aJXthFZIB
x3OAQy6jn1FegAi9l2ZC5faA4wJLSua/FPgP/+OZXGeS33GrAV9dsx6hb2/gLzCv
XsDMMDJZyv4/rxXWi+OhMzMGgyxHwwpbWvGRxo3l8ZObaSO1aRuV/E37l7uwby4R
lV6168oJpx1XCBuAANzOxAnCdR1d1LZR65RLHqXzcF/s4r+Bu6jn8lV6d37hkqJp
MlASv3imRnT6uKKEmEe8gwompiUEbewAgHfjLjErXuyHwbkTRHfRiY73rb7JJe/c
3OEldERhYPpB2MxLW/OdiPcNWrD0jO80HMIh5NAsTJge+rF3PYlpCvKqY1loLWTo
Jt39NVuqcx5AQrny/CQUvOjkgkn2uceJSZi1Yc/+iF+I6ITOAadTSTLEtGXm9+Yr
UBngiY7l3GQuOI7FpolcYULmmMbwI9lbWLeb+1Bhua30c3+UXEHodtrV8J20fIQf
j7F3I51ytJt3dhE0jU4PLai3NjdGk+kWY49cBn61burt/tLjA0HOKSDNj7h4S9Yk
4NKQk0m5G9aR72NYRK+6FSa4AOSbHMgMvsP+g+zVf1PzTPGg9uN2+0ZEELa4DP2q
fDAwW9QZ1o84Qx97PySjbcUud4/z91WCFQ/Xao+1kXYFvYFFNjCAAjKlwQir/Vmj
lACrldVN8s5okwXZ0bM39KjwCWfdmJGSsWdBKXF8Cbqik4dC/FaybAarY+UrKsAl
PWFNRWpYEHzI/W+rFkWRnx13YB6bkWk3wdPz6LXQdyQ+mbgJVipnpVroKONetZqD
meR9KdmRvAEx8mko7H4t116QJVTMLfvNmlGTwl5QayrFNIiCpkMBfs9hHOiy8AAA
JapO34DskQRXYb2CR3IwxCHZtV715AE+xh5odb//q/QVA9MNORuOaUdbw6lGmwnA
OsbaVDLhxxx5YV+MtN99YbZfMAiRfw02670abikqnTXQ0x7+dpdQSHaTxuT5D1Qa
kGdL5t3t7UHwHZr/gGqOxebr4Gs9sOF7Hsi6i+D7YXdWoqiPM11eKMAS6w3qkoob
ytRUKawG0Ic/w+UL/uLRLnvhmtfGx5ETzFfdteEk0GCoXQBs7q4dq9e9WkS+BqhY
UEY2twKQ+1mcjbhKq4LX9MfbW2+tXs+Hj1INameGVjYUO+v3ByDv+fCFCmaHeB66
/FILwQAVcCXDoThwhqIDs+ngS4Y7Ii2X1uyd4SUnhpje7tQNydeSzfoancLG6wvk
tYOhB3LoQY5oxRwU+EWsrLz0PmFl9KhQDBDdoYgNQFgu+nM4nkmylmYcW8pZafkZ
AjMzrVbadaxsYoQbF8A+YBmH2rpKOQKxtFQOcgBtvmrryyAMoJ0FJ65754swOxwW
Cg9LYV1nEN4ZN2F9UgKLM/RBwP7LwV6za4NUwQyHxu1wQm8N+8OCi8WYp3Mbo1Hy
0xh7l2K0CfVVYA3DvHUH18fqlne7kI30D848A9dHHr++Iodgui8FgDp0JrNcoC4w
D6B02Ln/kNxjZX8FWkhYfzopbuZe5RS+Zy0KL2hMRFoWBRYNZgfl0tdaNAUKIvQT
/IDI6wLowWLTPvI9m9XAnucScaiOkfEzhePlG9mCDYeYcW10WCH30XaIF7r2SpGZ
uxuUM7Zl64XKOcfy8KqNd01B9d8y0li/fJJpbYCLhyRhoDlFoAeZOcNdNp7M7haZ
ukxyz+HpB7J/7xdplw4y3Gy1V8O/Jh+DFMcNCYjcuZuv9Ic1sPFIvL7/D3XpPteH
L4pNvcSbZD9GvIwoohbohrF4Z3R7Kk5npSFuyhSwuoOxKtcc0CRKI/s4u16q69AL
nGuer44/dVXUegqxr17URFlLP+IGusC6x+dosd6mH18I0eyaoO6mcQBlU9P9LYkI
e4cQLxcxV2lgyiiK5Y768iPGSRfn1KS98VpcH8TvGiDYDJMR6eY5HQGtdRfKTtgY
CdLaVeFM0f+b6ivckngl5xUzsSab8Ny6Ta27vavKP+JxN9ZuahIAfIjZ27tktB+g
AchKBkB0Qdim7RvjYK17CUrJdR5cWIm/B7AYegDlRMHVALxO4bHx+PpGcxTdisNG
m1Ws5G1lVHpJbuUrdHG1rRo3ONrQnc9Fw6zWr09o1NtlVoIFHNDjKx6W6HxYZxpn
4a9SGXDTNJxAK9YdHz+uOKev4Ldpb6393tNIKv3jfxC3svTtLSG2PIhYLvDwqefC
C+SSSsCpzrQXvGCuLgaHo9DaLEQi+X9wzXMWQW7nuD6snTEyhJOieEwT7aNQycZE
VdMSasOhM33mmThAdCj8aZGww0qdoAAm5KjARrACmM8+RS5J1FNoZKmGed40RVIf
4Fx06R2rGcUwVMv/HOyqAFcv2uDujhn7hUEgNDrQaYPAOI9hFyZYtjn58gblMRKG
uwbNEjNdMFmzXmNLu/DrBMT2+dx4gFw/xoREZXaO2PNgr7PFLdCK3fls5gqxVBb7
UOKjpVUOaHouTG680t7+zrcLmLSmXwjgfDluOqPS63+mr40owyXrV476BGBMm3zc
inAkcBI4bt+/tpRpwRinSmLBvbA2Kj7OzxWpi6D3R//+pnhdTr/JotgRcS4DrATn
xxiQVRBw2SYFqjEgrdCM5ZhUe02TcqL3rYbRApUHHRG3IzREkocHaLO5syJceY1U
PvKuseiCtrL5Seh+Fjl1XWBaDdTk8YXNvGudhiGqEbLKcbxJUGVQraEZaRxMYTcZ
hbWGVKvbwpuhTZ6Ehczkk//zdKGhU0dOGI5W0mmnKTRbJK+xpge7Dk8WNgj2KvM0
kTRqs9w0eWI0Xc/hVcayHLQx/xdHqRI7K1Q5fnYyCQc16xgF/HNbEHmO9m2qLgH/
ZudeXjUbp655scrvij8AkMEfvl+RtXENbbEkLcy97OHGYNCyQZ3tzSQPWtg61nGt
SbSHKUmKJkrHXOvxQAc84RCPeBm8+P3O2VNlLU91LcD0gVGkakyvdOtEvN8jhmUZ
OcBmuD9+8pw2mlrSyfmepuQXO/0lNdGHPdUI7rm1qEPl9QoYGhMIBsVC4dbro5KN
ukOatstQHBrIHQYBGBZbJ7P/pj8CguSKv+MdlsGelqyx9eeab6h3Y12i8xLDMC95
h87BVUa8agfHoJsIJmHwlZMp/nZ288CIaaooWVr2cWMU/cq67kgIQ3r/u0TvcG04
RJQQ8H1Yh5BKgoaDILkBc/L8pA8CMPgkNKhS94ti2ow/aPNknVmSE9FzfVTISh3q
7tiAtvxeZhVsT31JfdtHKYkaEjnHjNjr+aAG97tJcxasyIf/stYMJv1VzNUv+JhJ
OeXrgm2r9Ju+cnBfqlOw95itde1a3nla6MXRcTpbeG6KZQUKIjrAIWLI9RHbCmq/
ldvHHZMzSQEZGdfEtlkEaCRY6t3PiZ3yCSa55zOg0d1NPgdZVge4/FkolCSdjDtz
4nNKy/xmWbPJ6Uo8jhufp8I5APiKPJuI31hRJZFdUA2T5HFM/v18y+jMaiNjfvKx
Iyd7NXaQhsZ5pDHDhaU04oqLVTFPcf/q546Q5xU739V88ykSmzG+EvBSBALfQD6Z
oiBjvYheBq+H3SyfGrfMnbEZCY8p5LckjR4IUK0QP2QoneREOcLeML8zKy5B4xMe
arP1HLbdP7LsRS5pMB2y3BhY7Zh+AdHN+c3PnnGcN0J0FCNPpplDQfCQLyfnDaFo
LawJopLB9sANiyH/HXHpg7XH6Yg2E7o2Dh3CrIp4YRQw3ZwPAvaPxQRuDBQxLt1h
L6jTvd4Q9oE13pdX/qfpLte+moqSLw1Zjll91JOyvOLhccrrTF9uAAa2SRbi4/WG
IaSIpOjaKCs95JmF0Pxzfq+0NBOhNmK7EsisYf2Wtgq4X05LJlODbI+sytBcZc1a
mAImtjU4OCjOykMPkaoM3cv7nyE6Rwln78e8IRsotIjvyrFp+n+mxGG5/yqF2qQ9
nRMAMzYhRK6TC8S7SG2kAmk7P4r1pUcdCEW/ZitLTd4SJogCQlLTUBkTmKRxVJ4V
NI4i7QWnB0uC8WANE6L+KQSps2BVBKKibjDeoWL7qqaoeMPfWJRHTjGXAQYcMWuH
lA4f8ktMqGqM0DKZluORL1VZG5XS65wJLQwVYtLdC6HNtAqO8daswaiRlADUnFwo
upSKAdvHPZfDoAhGQTv7HeevH2wX1Thi264NTfjXJiaXxW+WVm/TFftEVCQzSM7b
BGslqK12Gkja/GqHiN6ZLjn1NEK5RbHuaLdCiLoNz4v+SiHmomH6IbTyfHfVr2oR
9bKJvDQdTyNRWYF0BtGoiAkTA9rh8QC3IDIL1Hn+9SDz5hBEZhIyVDKKnaO1M7wo
gZ6SlDeWeR+Yq26DbPbTmNt/5o4bIR4yFBbIg5QetS7Xw35VFaeuW1IyXu8PdvQF
YgUtWD3waaFqTd+zSi/D7Zcp21EnbJLMZQHLxRlJoho5gdZDWPvILgXJsEnAUYjr
bDp7E57e5UQVOoq4MloSMDzvYX59RlR8iqBJKiMDtTfRLUTvTSnW2mTh37MEd4fB
+XabThFVjFgZBTOr/7cbHE8AIfgzPDeMHZJ/CpvAR2bpSB5nZY4n1UwMz1SB7/aw
Lt8VtnXWZsckEBbKuntfuEIe7jpq6BXIUg6v9JQ1wdch/AAHwG78WblmyaqiXlo3
43WWnpqoNgDsmZd9ZZda5fdEhGVuAGYhZ2MPFAkV5k7VwK6N6ThnhNSZBqLY6tk8
tSjCuCavKMr2ZGwny7t4sJWVFLUBZzGySwFrsPIYMkLW7Ncg4xqjiGnfjDDYZ/aQ
/Y/1X7TkiVloy3X37AahJDeGPGHOxVgKAA1GJBgulyydr6Y2E0vrBr33k18F6FxH
AwrK3W4yUcKDzvkM86htRtqNLkiviTa3htsMSRfB2S+Z+JKXw4a5dIVMT6S10yfO
PRnWA9cSc+qBJUjyLOfroCoifJweRpk0Sv7oHno0+wmvmcA49D2h2JVNNK17Fqyd
2f4wdp8akMbwZbrysefzErKx6Z0jwID0bdbrvLVzJVFN2vF0DR19l7qECSpsr7aw
XZn5pTp52Zl12kFsIPWjsxOMiDBbkYW2suTZr1JyzbsQg1Qu8jtXO5xe5kAiDYjV
x39Pn4fGGSgJNu05ymbilkNF6sPK6pe4p50pCYabSuXqdN8oFzbOHf0y+xS9870u
SQJ2xXNLVIvI0WX6WfhsB3ijsHj01P4K83PLHc0OtUcZ7MTj7vIy1ZnWwJ2gZijl
wDt1I4wS54MWFrxWmf7N0kR1N9XqpJXesG8XBWJ6PZisp4P3tkTKqLpdp5RVc9TM
w1Jzd09uZffDDphKBFev656GkvfD0CTMgCa7NWsRum/yzmAPRosfGuPz2kkcDnMO
39MIacC9UkVofKcxrsxUIZwuI2Yzmynnn9s25tRAJaf16Ae2TRxGtY3aoC91g1ut
QsDiZm1PzD3snHMJc5+JQS2KVKO3FQ7MSrFlx7zB6NwvXu/ao0gM1BF5rUMYoNfG
wDzNCpSzBWv/v72Sw2aEFeshRIpwILz0kL39fImF8Z9aKU1SJjWiHFJiGHK86XQq
3IEMjQQOFyJwm+CctN8yOqhi8lZX1sFVLSbvSPdRg8AaRcdl81t0YCSvffzQElln
EpQxQw34V09Qg71MKG3FyYDd+WhMSy/ujiraULIFUoTZwVN8329MgJRWhi5v+A2J
YqO4gXur4XNy8VdViAJI9YDc6d9duq5cYT0huTSTE+fjRBDKYYP1P9OwRGW/QsaW
Ba1G3AMNvmOcodHVZ+mIFPC+KrI7EsfFUCPZ5d9saY6vr/IePjuNE7LCrGlX8vRq
5DQ582VZVL1QJrAHzlT96BvdC4dZBkUH2I1pM02R/mfppaZdaha3BnG2VOREtaAA
oJPMs6PA4UdfSbIsDsF2y+0lBxItbwSK8gTIzJzFSxhq2mvmNd3WcJnYFgrPGoqz
Kc7hGNsoSLekV+4SI2WXWweNAPV9w0253pTri7PuDYJCYYdNhl70eK0VV9DFJzQk
qDw1tpMmfJKUJr6ZOgZo7OBQJRrXtr5ZitS6frRArr0zmP6GyCBvE43hvAwVfbD6
4/PFjjMfUrPhSREsMHP5Kk0Y0e2bQBjLhlJI2iHBFbo3lFkAEe8cHIPtmBhjm2FT
L0szNwPIikdZ3SUAQS0iiWS4CeSVCtQ9BUZ8zoTlUK8d74rSU0VsT2uJPLvEo10p
vxJRlj5lnfzgku3L+s5ursRugYgVhR9dRTnhVNQOa66WXWmUWon/FTfMdSBGhdKo
iHZZyTzCLHYMxa50PM3G8bpVazV5F9iWSSHQl5jKk5nYxD91LNDzHaYXGSPVPQMC
+syipES3YYmFqNytyZlWU6PzuB0doKLiA913rot6oadrwzmtoFyR50SsRGckCgBz
TIRnpsuDu254Ov9jrOhEqkQMvo3xvEJ4ZLcrvvbAz6RYlmTNuzZGAPdPO5PKKkpW
N/QhvgG2cidGSrwXgzy7rNXfvw5rjvKgKsg+Nkywr19lJ/J5suGMnn6gPhcAblcw
M1HQwVlKb6rXjnZy7GgoZ2bmYAlsjBp/NjPa3awY4fi3AqJ9XHlyEH/epHVfCzdB
dvYVE89xNp0FGsYG39C3XXtvYNBlJ7ZxjAu3ztqidj5LgECODUTs9JCHS3GJYrev
zP1w7gGmEREo56k2WfUywswBhvHZJ84gSimQ7yPd0UYpDOw1dRbMY4lkvFn8jUBS
mEtXMk/dgPIHFXSDtjHo+cszxWgfk9ZzyJ8QU3KWe+kNxpbw5pRPI4CkG6c1ZC/k
qEUWrQL5NEj5I8hfq/8eycDwrbLEm4CgDRKyBUXQyKsGPXACIaYRkqY4D2wcCwNh
xgpIBJnHqhDvXibqEjcKE/btJIimPpNgcni9nglSynZRyckOcZ2RpEDD3PGT93TR
8X3lSaobeWNL3tkHVS3Er5hdLyPBuka6JOY+Hro+mccGZNUWFZu9NbIl2g+DS3ZE
o9AUzJEo068ygJuRBJNUJECnGOOuuwhEwMUaA85WDz5czc3kgOOFNxALYmglEZgE
mfYn4cxq9ZQ5GzPQTS1S3rw+9zQHSqYG83Ehva8MaJWhoHzLcSmzC5B9zKGjxa6J
oIKnpayKXz36uVP28CECLUEJaHrdF6aw3JiwFlKPYDnuATzjZz2rKQsCtCorhZ65
J8UDnZfJnOkPYPN7UvCWcTeCy+Hgroa6Bvfs0mYv9L/eWvfYvGwR8DgVx643m3cZ
duhONwiMgRw+YIoXEbduIV6Yi1bMdmAvVeUV9bhPGVhL9YoW9/ucMIdz0fPaj0Cy
8XRFu7joROjFT8Om+ejf8KAwtorXdnQKBV/fq+sO622+rhzvoVvrrxrKWwgKT+L4
F3Qq2GWTE0lL8ZtNX/TicEzAySe5HUa+MlxIWjz/F/ZFOC80tRGNkEybRdV6doY3
1NNC5QpgNn3oRFm7pVTceamweTzJcxEdxvwvjf7cB9+9ddpFGSruFa1XrpcrvW5F
J/n1q41e19E/iJHp2qNwa6VDbZxVZ9shGoRim68q2fu13K4IWl8lYv2D/7fuee1e
wSkzZfLpdiNFxZuZZGJh/SkfjJRbD33b72Xnm6+8YvXMt6nQiI2dGcbezNVxjJjZ
fwA4hh3FKi5DG8m39lpCXeY/oQpPysdohdtybzU70zV491e38x1mkyHYPZpjeWLK
TENC8blnV2VIs60ZiroYfTbSq1IfElJJysSXdVrzR76aXDOdVZT2ZqcQSgzgNzuX
bKkG4sxRKcYDrHSb8DHH48a7LbzN0OBExKCtQB/ml8RC2LdAnYnGFX79hcPIOmt3
xzSSssQouVWa2BN6PG3M5rhlYdIyLuNcilcnyDt353qox04u9BBuY6xYpjs3lu0w
WKiLjt4J1k8cFp3o0Tf7KoJK6r0THgtVOh+GMr0zWaQeiW/R7CyfaHEBVaL/HjCJ
EwSD3DqcE+uM6UmPRSXveA7xl+4CFrs1kjrK74foe9yoED4Uv3TrdyhANADL8NFH
HFkK9rX6MlOENUGhSy22KnhgBrdk5paKa8nqJjUVdfTthbc/K3C1bB/SF0sgA6VL
bApoKot+zSV/fxOH18q78q9UZK7DhI29lL7xxrA5Le51yO2iu6Jfg83qu3KD7VGx
LdMZe9JATfprzI1G7sQ27/wv8EvuHajdmGo67xessngv72Xr1pr/GNjRSuG1NUDZ
7PNsf2OjlkToB2Sabc67HKRQWl8CxU1NCb2QwYdzKSl58qC51oapXWtmBt2hZZ5/
brqNj5HysDV2CXrtE0QfTTC+dhsiNIZw7emxeBC48uOT0eN8eh1JEH7qNVzDbHma
5dmRW/omxVh8hf4MSUm/Kt4+mfnMoFyY9EH9GlBHA7Vv2i0V3byQGzbB1gIM31XY
xtCL6D9UAOLYVzgUBXptolatMSNiEwxP11I2fspT4lnKEpaCz06vnYUzKbjcB9ic
TuBnR75ZU57CivNCcq7rGhvU6+XhoqZAVB6vrd8QKU4n09BEObu14yiCIH1kSb0Q
XY4lRSnPRhofuw5joDXiGy7MjhVEeIZTJskXquNrv/HHaBJDjuFyUJsSeF+CKrFq
so2W4bAR/5TQsra6DagIJQzJ12zLD3BerZtVpvhaLVvUpWk5yHzhD0+eOuIvNxO8
+5L9ILGzv5mWT0wU/eE52u7mta5Foy9aoTRcPuaq2gYbpb5RqmfsvR2pCda/fjhe
pKpE9RPUIfOMGvISZDJx5pp4kmZBuytemExk4Odvd2DALfeowb86ZO1Dh1tnRreY
oKBIYxL+OOrU4WonRCeo+m8KT4lb7LteaxLW70gkNZMIEgKwZPWIGDFHPAc5Yh4k
FJNp5y1txUgWQtFInef10WvU92j9cRxrIGVJjr/3moaclkn5tGkkNuH3joB3RNDg
/E82lZQRUbyCGCBXUI/0PzMAQ48b3FcY3TRGAwyzde3JzRdZpr2fzRfFBSuBzvtf
3437h8E19OLdDke2/CtqqIG3x8yeMbKXOC0pqXppg5k8ijTKAIcklyOJqPXj+V8M
udEMvKR/S13/WpY1o3s+SpVir8dgxizvENy7cnYrN8vG/gbAkN6Mcb+7Sac61miG
Aa1n/svAZ2a+TC/L6NMW+1IiRbHYycyHH+GvT3dDcOc9e66+kIgyZyqOdXIJnasV
hOgAefvC3zfgNH6TpYGREXbJbPzGn57eogGlXWr0ltAFKjrU/vSoYeGnuUfsY7s2
rjTzUSLN4nAB9R3a8UVu2OBK5MBFKrQ2Ikm1yUggUxgPsrM4UocnSMuZ0I9nki/W
S5RCv5xx4hiurj+MvLq8O8JsTdDVVSgoQ/1Gk2pyLhGBeehpfyBm732nPFCn7a7J
TvG+TpU583VtxWSs5r0gKMF0MUYy2yfldhfXAKOG9RdpP81ynml7omtTkY9aGWp1
nceumw9P8NkXjiXbVxqNy7L6q64yHzdYDwgDfYQFxGI3tCZGF4/Axr4pc3dXHQ0p
5DS0BH1cMc1T6ZhcjLrpbT0q8qsUdQmdhNIp8IL2zRBHWfVin2CQr/qVvaW9fBjf
dK6fryKDIJnk0VZnjW6ScDsFqbEyr7jUlQDIQw0430LAUcCQKWNCRTGw78hdVPEm
0lwnuLxdqvJfyPtqS8Y7cpmDf3l8S4KH/h2vtV5TSW9KHdONiUC18Smd2lA75RMe
6DHMixHZgaW6MN8FBFEau+f9pkcpieovJk5x7Tcg9C7u5CYxBUBlD9rqhENeDlxw
cAlkmbR5RINtst5kXuBA54Rqb5iD42/hWuiidB2Ox82BPujCmz9IkQfBBZAO9dBV
ifyZqnSzeZ+wKNxSyA1wP5vYSrGtHxBWgepnqp5dq4W+RX1RH0c161hGtNBpAnHb
/0kZ5PMYn2jzYhzUTzLw4bTbHsq4WysYddnobNQ4hoJm42crADFnNY9E7AQmhrnR
drXsLCCppQEzqWQeiRehY5GT3vUaEEbvSLBT2pQwBM8qSeZwtbc2shpCmpF2H0g8
Bl1DskjentNz5V3v1MvrjkGhB28lYo73V7E9C07D6g2lzPMoND9wV82urlcBh7s9
FDx718N2Eh62ofBiKEQ1At5J/dpUBl8tES9XUIbhkbjV3vYkswK2q3x95iiSosZz
dxrRlTnFGbnyyCQR6AKcf29eNxrUd2TQYfchSYls2oi3/MH16crTioM7MM0cuS3q
bJAbSEyiUZXQJ9ydhmv2N0GE0vpU5ylhc6X4nWUU91o8TTRke77M4D6iqjOBcLTt
Jy3x7GSyHT+18dSJfnqyMF6EoxtGNDtgHKZDUCLW3u8uSQLSq5l83Hk9MT+m5UCc
S9vZSxvVptHus3OSH+rNVOCaD+hHbsfrQXw9KR5J9K3JQiciXv32FIwjWhU2HBdm
F13dW4jGYVBfZQH8sPiT1T83z6WyUP5k87vVj84w31IW06IMrzye/M+MXOQl2KjT
HRNqB0weRswpzSu3cdpQ9sMsObeFdMNlxHthsaIDLjwGyARZ1zJIaFTnGxkFnC2n
EsX7YhNYFwFu6fbAjjT0j5yHbT70lx0Y+KvYbBCD9kAien3LeDtbc+de9q9ubOzK
x0EXN6uYQbexGwt/oIQEAnOajfCsv8nJfmRJyFJaN+YlGUWyMFZ1kMjZT6GveSok
GDU2xqq6ZFI0CD03p2jjgSriw9mU5TsBTIJ2gj7tTtEbKUpyxkm0WKahf+7Njd+v
LHVBeed1+dBGFHqs7GzB0jkYOh5diMN6oif2fm5TmzQdLrhQ1BCj9yK/si7J6E49
HR4Pf1DJ4orfz7IX19ukLEAqbv/z7ueK/HgISD9yY2P1XalcHkvEgpljaygTPQWT
dnaZuKBunB68mAz3bZ/MQttbJC9BeRUQHTGQS8Sx0xlUxSRvDGwnWRzN5Xw4RfBm
yJWjDfLt8MuDmA2qdUmIK+fMAsrzrEzURaP134Zs8zVh/mLUdyrcXx3Ulb/Kf1oC
uVTy9GmXXyq4/JiAECUx0mgnaRtPQGIPb/KzyRmUjST+cORfko+HA86pXxXG0DNc
EQsVSyxvJL8AaTyZr9YBgFvNaJCXwTs1THXmuRAR3JNXSsrQvNL9V9Nez9T3m/S0
UAz1BT87ybSOL6gwaB5iKB1RpvFXh+CR1nqH4mpU6oFXGkb9yUKGy83ShW9Y3rT3
nQfrdM6lAuwQMdwk2OBOOvPtsG0Smt8nE2IIO0DlD6tTL43smDQoBRmwCW4aEqhq
iMAxNS7y4+dI29ZhC34aXpXMGbv6JcrhYzuGl6KINv/UY7GpjyZBijD68vdKN8gB
CW8b+oEGBQD7vn7TA0y5wgHRLEa8y9PKCAMZYHCNAU+eAhkpV171X0Hs0o7XkHq9
bIHYEe7K6/ubTciL0HBgznnOJ+75oOBAMJ+OHvpdHA4XOwTo6BO5HChHPuiOJFHv
1BNiVJWjZAqrIUMfLqS8Nc+EG2+n/S7fry+t1AYZcnhWPR1rNq07JzqBPYaNFrfV
lYuSfXsknFwN/n5MWxZUHplf77tybPjxok2c0+ZJDGWgZHpzrBVgCY23XsI61poq
6dU/3Vi5Qs5undRRh+zReGsZ8XLPxeUQWnspVss/1oiH79IeEf1LNL36+du9uf+q
cuKCUNZoG0UwXGzuSWUU239CfFu/nYC99P8tfQfHM159gI1zGjdiImMeWJTjE5LN
XPjmXx0eLgpb+RTOz/tauO8C2Ns2WGvAwLOaB564pRXM5MOzSOzW2IKy22ETmm2Q
BSKq9fJaeQwGJFshEWK7orBcElyTyuxmBaj2det4/vqUYb2AvPAVl7mubHLYfhCi
xZ2h8jus5XbufazgYkCAXXci2FU8W33IHr80qNk9EGZcpq7HTOk+D6pPz2RfVwcq
rZWpE5xGh+my4X3NQiPc7k/2DcEOli6MhgmVznmCK03FXqseh3ENhM6/wo6BSEln
HawiVcCf5h0ToxI2cfp0mbi2MIf9mkJAgNQI1d2OsPl3U8/Rp7pB83ab76MtMjPa
qqb1uCfGOlP3b4b/cZVlnpK4sjXq5lyY6RFQAB83cbEXpakMSDsMH9t3FtJg+2pn
Pq3G3sU5oryMAHk4k3tKOuEBy83hafjUrstg/BYCYefnk1sLP4ETJZBlLM8biyaK
EzXlMhU1lJjiAu8JOuJNnYg2896xgcy/9thde4io1teVK5keEq5VAY09/LfkNcCh
QUK6d0nq6Kt9txLmkldmQNUwFVlgbXcg7ygZB0yawLoz+CtWHSizx6GsvveYkFlq
yo5IJesZSgU001H3BqV9a6BNt3wdaKlL9TmOVeq5pimjqUB88QnxuDTc3mc0psTY
KIgBfgaXnUv3BdpwmBepu2/s3aR8wMS6Xnyl/OBDrmI9/nEmNPQLhX+anJ46NX7h
ZN8EPGNHJZGvYZYkzpF919pSqiYJPyFY3HAwhH+HS3V+irSfAVGLVcNgTl8SSNPu
OtIV50Cq0E/vRX4MV06zpiQoWZpjNr8pCLoElkQWY7Z6FVsyXCBkNX+V0z9xkjVV
UFEiMdhrbmqbpqLReizNZPhVGqCxpLDt7ESxsOb/ZSMR6xTs9VDqFdagx6Pk0RIu
6pOZlD2QV6mCXdrzEhStUtfwkBaY5MIxql7N0eUNK3ga0eYUSY9NeEAylCFxay0o
dSHO0sygsVetfZUJrvTsYjyk/Ys+aN5sIiXAEBidgEExlJLisgCsr+GX3ZWLwEgx
Qu0Fmr+9q4MMfyefc9sbA8jlIDSOWAInOALkhtaVw6nJ1+WDor9IBM5GVm9wNtPA
Wsy/w3KD8u6ThmzcpNv1uuvI8AMepbWfTZBtrwcs0o2uWS7d46rpeOkCazuXCh6f
za9JjU//FAkuZrfopPAalsraYJIfOFsxFnkYJSjE+ZjVLZlMDrPC1dUwJfnp3vnP
h2i6Es8H5lCBtkh7x6Q8hfUSOh618RhAUGS9+fLOghnn7iK0/1yvaydTbeenh1Ac
9zjW6wo6zbIGvvN1TtPQ2cV1OyO8Gq7M4pf+ia6JBXBv5ybeb8aBGmBeuCokXA0b
TAQxpZoLhQ0z5aRLP64KE68wPinB25aNDuxFRDCwrnYNVs83jWNr8AP9Qo4tQSwn
vucqFHq1QmOK5jeHVGhbmP4EcE2gxevHRbavmP2dC1sU8PgrvRB2t/Xs4f7xLMYJ
gR978ZrZbbsSy9h25WVokW5hBBHJdlGFUKlSVS2bJwJ0sFlym/+/vzh7Z+avqWxg
Y2DbkGyaP4pz9+D7C+eWnjSjZ4rnPvwOMEr2MmjMS5qet2wS/7/L4WvvaRQebiZo
w0Zfoq+DJS0VerDbDdyAmSmNAy3ZFC2n1z/RxfJxcn19WNRviwKErDxvKFY6n39h
mijC0lF3NEiUAGW++8KaWJjLYJJ9YEcP0B5dEc4AlKjwTyCZdrhFPNAiq6890tww
6XdDxtvrkh1156b0UWsfnV+nORbUHeo7JYAPvd2uvir/CGuWbCMRi/LJbIu9RLyQ
cfOTPPypNHYRchU13089/qWEMP3DNKZoxmp3oIL8rkd05x8Gfjh+MlmqmXi34TtO
najW90yptMFyui8qtrVA78EqAwe3jHvJF1aSPe/or3E0GndtiOClr6nXTqRg+iA6
cXq2irqULnwwmgrgb461NVIYzirh1h5CJMiPcaLUedcOC2UGL0jYA1j/nX2ICDIj
LTw4tIy0wi4tR3dJMV/PLED58HD6IIqjRjCEhu9LDgzV2KGn+AafXdhTIUuT1Ft5
01VhAcKi+07X8PSQtxXfpU7G+a1AAIwFRJYRWJnDNRfII0lUA+7vhPzZqGyMIDQC
dJOpdZnSkrAUIiZZm2hjLYjE0AzInSJE5cFVH+i99aKYDQZVzJSko0vF2CA7ngOW
4R0DalRd5Y7fYK18Zw1jSSIE4KIBJC4VcPVu5vKpeBDr9xiSXzeG4NY5aZNsSvrT
ov9LN/CVbsiC5onC8pwgdcnc+rSOhS/TwMAx41rfp4r/g1EA2y0CTLqNArTMyr6D
OEDaDdI6fIbJ/MQqU/3eSmvsmLUq2gC9l4eXtJF1l6LKwOSzugcu01Pil/IrsrbB
wNiZVQr/pyJyWXqrRsq4jccfb16jAg8xAVDW3Pm/zvgebklIcnRZRIcP0Yf1CS3Z
GW/rLVQ3h67HibjFCoKBr5WveglIDQ6L9TkIJRvlms4qCk0JdoTuxmfk/wFuGcg0
67kII3vKm/j8KzVpJ20R3VnSRWs4wE9AVm2yEX5LbmjwCtNxr5c8YUpkkDfu+fFo
xZxf+xTPKE8JE87AmdQW7NwP4j0xoPaHpuW8dpUH5Pp3gLNEofzMyxsQMgk2KAgL
1+IbT/fCzf+BnMu+m6prwKY6bXudPMWX1VuNXo+8qVrE7aKCBFCNVhq/VrlaE3WU
7fZtCVdl0EEGkb2PsUpVcHbHdt6TToHIiusgYpVS52zQ+IoJd/bkQ6i7ebFypsjw
5DqNDbTxXLWThqO05MJmepXu9/vo/lW/mSEg5qywxWCeX3+WCy5vCrpcyNREzQbA
6FIiREY79uR3dAbyidamoZLzVRIm9lXC8GTAHJxgpxp8RyAVoY4rOfanUr+r6Lz3
aRbb76c5VkhlgtcOtsyUbMHo6FhisiVQKwLntx9JaCTomPvy0+oyKRlzEm0VbsBm
jnEBl5CWvZo6HDP7JNvsx3RoSXc/y5Na6sYtuVxGbu2Lw8tA9V8zc/6yIeaJ5Trf
lQpv3PHi4Y021FWf6NlBl30VoMuR4qtC4hqrccf6v4dzjMWtjYRYgWqDIgPCaN6/
5SwWA1NifXwY063ILNU0/Ga7CrVQjtank9y39HlSJvqfZ0t6k2/4p2t9QjGqDy1l
A5rqMy1p7FvoO7+v4qw8iri3V8LIBOpVEgH0zmixpZxUNCSj0cn38amaitVzKiAD
/fK4/6bIwTCD+zYaouGDcvPKdodc+XF1xREX2u7SHii+Nl/VG7A6ga+RQJyKjjSq
PlCi+6DkfMmrNtI1NFuVYNTLtuA2DBbkjl+YmSPiwKFGcgxk0LGYe9fjB2KlgzZ1
2iTGpGGqXbmG3sBDMUzNFImXCnrcu69WqU7xaHwY62M6fSBvZebppvn5ZeWLlHkE
0qJChUxB92gK0Pph2Gh+X4YJl+g5/A/85PGVKdlNEvVlYRZ5DhzjHaYzUQcl4NVH
9k5TZUkg4ehxL7cJegPZEOxI3pWpLDJ6LAKIUyVt+LUvPXll2w5K4hL/MllrEHPY
Yje2ErhiZZNTOT2hkHTJE0dkvSC5LNU/uUu/XC2pZfThnQEFqNAffm+VI4CKY1ku
9tOTYt0pKwF9Ia2XpqK9cO2omAntmHFl3rIGYQrPDq8sCOvalkGGVdW+IfzMtS6T
wMCKp2T8KUZWRK0BKQBFvjbAH6ZwzcHAoFApA4vsoYZUl3znKGPqxv9apK7FC3hu
hSk271ptGPIt9YtnVhTRuUI+tTldBog87PUWRnbINsY93CtR6TYTrsIQvGdqkW0+
QbsXhnt95MdS2R3foaEGkGZ28la4JDGmJ3aSChfAeo3//L9SDvTedDfe/oqdqo3C
IwmlEPU9YDRKUZ5SmGjB6rOrAj10eEZKvoE1xtbP+RtRWJTXa3Ugjl4ySZWwgy3s
iLEb5HIJif+XuoooRtYARexDA4fO0NhAr1fGeqm2l1Jm+wtY8RH+sqCt2lL7noIh
hztMSfGBDFnawaFwqBzvV7FNyGYTOv7t1KBmdTIK8RPAmneKwQ4Nqb934HrZSKUm
IgZ1u9hQfYTgeMjSwTpmd6A1ioRutmFyRLL6dQP60fz35M0sIfVzEz/6Bq6Y7LoJ
1UlH3Nc9Mj+RVhJxquKuY9yBEh9aHbUKv+ybGAmSTLJs2Vs2Xb+w4J8e5/2FVWHu
6n213MgldRCz/GeINHe8Px8gTDWRhTty/xGNh5pmMmSQC/8OEDIx8c2Elfx6E6oC
ZS5/rzAV7kCQzU2DZk1wctJzqi2zbzmmLw2xgRJ90DIAE3oaNKtQ9JMP0RW4ienY
+uUpeFWiEwLs4h0LxpGvYmIk8goGgUUwzcy8TUyvjOdUCGWnv2LlwzuefTgMXNd6
rKhBCkX1WZOYzBUolmTyrAPA+H+S6bBZHusQ8IpbQbVX0sPbKnsZldp9fy2nEJXN
o02Yqm88fVWFZaBeWqvbEAc5bTcGrpyvYy33ykUZ78zWjiVoL8mi+0IBQ9n+B27F
4sGAVaGc34qO/ZaooVUblQ07TcE3xSiBrGiDvKhun2q9uroM8Jk+QFTIrynDo2TG
eZ/KrcYeZOzZQUv/cWm6PRbzCs9e8Ll/tHM2v90dVBtQ9gI4cUbL+4Tlqv49F5cN
ryN+EW5UieuX//Uu4pGqHZpHzPZ30v1cOp94YZzmdPKXeVyfQtCZr9kKO6q8XP1t
I/yAxf8AYJXx86aNJPfQ9QYjlhWeDi4j4sicCYHX4yP8OZ+UB2l4gyWRpl0gAD2D
TQkSYsmaag6jOdXALYXZED7awip6GLSr/lJRihih4TGKEOK/ya+vBtcYtGL92q9H
9MnqrAByhLeNLIf0gR780ykjHPkDKb7v0WCep1vDExWszkc2vQI5zWsQ9qabcTlu
EpZhEGeO+QwnbZPYD65it2Cotom9sQutzh9OL1clGPjiiWbRt+4kGUouY8LXrTJs
zKHsLtYaN+R1onLvcM9ezXE6TbUokBfADB95AuaKIsNz9wQju1sZ8f7ZGnMJfZl/
xDZfyHrbZSVD8N1eiBUdO4r4hoioOwFL4zOqr9Fs7yKi/5ddihJMDa4xGt1g1kSr
+0eLgmnRxhiJtOr9dHs6G1yTR+txyRG9/+Hvh8HBB82nHkw62jHxo6mmCN2Ej4YH
NIcZyqOr0IXH3I/KPE0ZnhbdOXeE32jbe6pTpt2swQ/19h8ybX5kngOAB38wqVwB
rc4RL+BPmBdBN+g3a2567FmdaABqLPLmDb6dC4YZdwdeO58L3meF5Nd1PEFuBzZU
3+aBzpLNNeGg72vrYUqnqiBZPUDy3Uaq4y7GMUQdVANUXDcQpDKLuGM9GTfrRIYO
5w36QKdAAdTqwgz9fLwh1cp09uW7rFshbQZBt3DhqP2bOC+/hWIxaj3bBlp0Sn/h
AmYwkF7DjQCtkTauXIbuU3//U1L5IJG+Rq8NVlQr7KUUrMYn4IUdOKQElMYFZIL1
7tTtwNWCL+TVSZcvfkce2rxcg3bzHvLN0N00BaSJIohHTJ6ixdO1ZRYEzVN4copm
sMLFaWWiLk1bVX4MPkDITI+qOxcEI7UVUHR2YOwRUzMZ/j7jJ8exB9sOJIiA+gRn
aQ648+cErifTVhYbki7XN/nV1LjcTdJVuAjVQWMiYn0jiYFoX9ZEHsAKExPcJP0D
GmUlpAp71wPGdNcCj75RaEQjUKXVU/9Hnm9GYC12Zs2NFx0nAk8LO415+XPNmnTq
BSnLkIxRbiuOrkrcJpw1aSBP7hd0cbeNYBSxiU8x1HFOXF2LI7INWhYfvE3Q+u3P
sD8+bMmYQ1EMPjacHGAgrcVy2ciya2heuCrGW6pvCBasBwYwO0+CITPlsmhtCiqm
3vpG6T7uLBPRtklmak9PuzrXxuc6suWjSbKT7bgr/oRD3EF7SgQ5GSFJ+6vhBP33
sCs6a7zIc7Elk5EI3d0rgLx5McShb8Aq3QWjSrPacXxH79+ggELX5TF6+un1Rad4
50jEfuCD4qQDwGluCNxPPnXUq5MMo53U0H5OoBl64mLuXR9v9YjWmhLboXLPy+a0
noxSf9SUF3LcjXpdMgh0r6BaRw1WJt1IDgM/v6hy2fnWbfcgM0by6H38rJDoP3Un
vEtvMOzoxBe0+jTcqxZ+dtjjdlSWaY3oF/lx2rmxFAB8fhLKAb72nezVB/IFuD40
kTulf99Zcg01YGR5F7UrMY59vLudYOJbn/aM/aEAz/tIgIN1dwLCKKnkInohsGOZ
AQuJ0A/HSSvwTRWyOdkRV1trmjZIF+MBUz3e+zYfRd9na7Kk1LplBTW2IsyPKQOd
tikYTd0oQLNXY5ylL1ZuMyPNV5r2ZR9c9ZYL5Irud/SBu0dNH9GCW3e57FGTcuZb
b/QabMQ2tGq5BRtveXYGhjnSoEJWVyAAINrvzKzqcDYevP2nLnx9tV4QGFXF4aPn
Ghc7bYJP1wnwyoSHrYWTbvBGxVRNy/gH1WKi+ed0gGP9Xz1DpOlIG/xE2FJPX5fL
48uye4LZEkck0Ivj1SeG2iRoIgdkuAsONn0Xmd6t6YuTNHVXy6ahF1XT6/bZwjvR
s2LMIHgMyrVajlcnAvVwCLxoO6rqBrTY944KYq+DlMuZODfU78FGibZubjn2WQFU
dHYP/GRHeoc3I9GnCTUZxf1Q5n1ryVBJaokkrGV7CHsXSMHYahJzkGGkChiSYPxu
1+8Vu6gHCWcxPPpsCc42oa6ftRS910cQMkgR9OXB5LgxJHOYhF6ncz16jAbH2jdR
qic2vICb/+A+X5ENJj9qy0x3NYfGa7yKR3s9RLuRV1xuH0r229ey/gQWWaWzN650
Aq37HodJIF9g3F65LnOOj0OvHp8ASZpv03MOfkzraWkynxcfdItS6kEms1ElyLK3
p/YqFe09CAYVPJ6lqEpdJhFElO6J3NEOkzuvu8TLUQd0G/TUo8x+fX6NbQLRJeFu
y/kcF04tHezCnqXmW7UzzhcSciHHrWyC6U0ax7E2OkL+rfs3jzFz4WjsyE+EWxWA
6jo5498bVCgSjIhOdoCHIegU5FNgRh19DnGVeR2doDz1+UBe1OpQfZY+It90qOXy
4VsEnhF7umEfozYgHYqNoMytB1yilf/BttIL/epXz1u8v2jXTELGLT4uPpcJfm39
fkrHrkgo4KuoKbMHMkwM43KQ5iY2ceU+0DfzMfqsvL/ZPfU0rPt3hnAmDuB9douT
YHlAAfoJbkpS1m2hzKre58kZ8aVyY1I2TsmRKlbxOfw0DqySetxaH0566Chv6y8V
iphemQaVRft8u1o7nLB0m8AfDUrCywBiPT8nex/U8iXXFhEgo61RFTIeQiUFUc8q
AT17qevvZG6lIPhbXQ2mV5xUQumXSZCczwE9L8F72WP//pXJEzVGRT96Cht1SyNE
WidMA3DgQG5Vet4CWwnyD6iY8xJVtgSTMzVWLyNk+EuxCb+Gu2UeE++anxNDgTSE
clU/446bC5km5vVfLW02aXzPe1z5z3f5W4VHkekilbaZGcSyyKKKJ94KLS+TkJz/
Sc0eeCqSsveDttc1XkemMOrnlEZe0GmqI6uWJfse+8TX9Ot93V0HbAhlz7U/wDBf
5z2eS3gbE5O7LSxDDFQgjDClFgUrZA3ps/Le+WefLAR4wiW/PsWcGjGhRsjSO7t6
FXhsRGVj6cO3T1eHjETG3dAKIuCdfCbL6NlVNVJLaCZF2d0Mge+LYH4+BWDH73Ah
U1pxd0IM+wY2rCBgZl6l57hlLS77+R7Vrp6Ojgc/fOkGqlCpZ8YsXueGKwQkvFaS
HAzWECApGVB7c6gDbgRIHozfzZO0s9EOpPaJR/yGLiUGqyjiBr9Zq+eQbzMs5RQy
WFhQ1bCt3oKR/26+AD9TjCOlmxq7QR5c7Xy81qyKdiNAaxGuc4i9yjNrzH1bk5Ug
kMIxpp2qTkJSKCjE8mipL1lIXgTsW/CxnCd1Pd8Kthf74WsbBeMxKHOTo+yniH5z
BtQbETO9rIjxakjAD8CiGAPmpvv5mjS21K2tKyyy+/OGl7dR4sV1hqy+IV5mPQyD
ZcO7LE1DSVDslmTvu6CZVGcBbfLn+HpBNlHpyOtkd8tI/NKJVMzWbR7f4JPK66iG
/e7Ebg729BJyOoHFO2/L8JZfmXzVfQhTsGF/dAPMVSPXqG04+8W4pYq3hb6U+JW1
FplfsS+BZRUkvH2odByHMc2qmW2ci3Ua+gkOU3mjkxAH/Gzal+6cUroCTPBfpBi1
ZR5hxUKi1CBnuoMVqltotcXBJAPD9b37MXJAIk9Qn1NgCFcJvyb4pekf26eNDB6v
BtdgxjKqHzPKHSBOrRxxX4gdWdeT11tsNRac/l+dVQLmthdvBCkQax8Kz86DBRbR
uPi4HvoA0HaK3TsoodI3Ezc86GMXaFm9ujcwdaJbdJf+J6s6iidnVDLSemPTKy1Q
Idtj1zop67aeSkFRkouBNdshKBJPM5R6W0hPfhQMNkAOw6OpOOb9bHqGbHDyLp1K
0wVSiK08Fzh76LAousA5tq5fYSZwtVuAw6NXALbpPW5vt1TRPP2qMSJ5COds+FXB
vOgxSKPXoO7zLqHTPk3sOAg+K7ErDqAPLNWmysiXwyQehEOm3Qw244YN/NY3WS0i
60DdVFkxwfsNs6FULUStL235ybPPVnTI69Q8FzgLUNnrtHoPfps1QuSxZ5KcaRYa
UyrZwDPsORxKrShh4fq1gz44osz7wc+ikqsvUojCJX3/VEaUQ2L32MmKhLG/09Oz
VEip3uyQh5aWp0zoYiowtDD/xFTGtlrMoHC7X78Tn0sJF8OBguO919ERfpzb9+i1
cgpxCGuja6jT8cZMr2uSoDjcAtyiAKYmpp+RbC+R1649P+TmaPKfz924/VcBPeJm
ForzjLm+3t9YaZH6apv8H4sbXAkVwD/St7Ir+ITs65WehgUWlInhPqtaaepIzDgy
xJRUtTIYRaAdBhPAMGJiq9zkn1qXE/KhGHLovt0ApPtfZcMnZ9aBlz6nJbOTu+aC
4nkfPEjGJkBKNVpD4vqcc57NyleqJM+c5kTn/3Mi/m1SsoWH99SlCg5udc50kals
X5cmm1+ngBYGBv/UcJbIXrNT6tKC8OtAFj7BwETo2MEoh9V2G5uNzBTEG0Tf6J4B
F0Hj4zZVEHLYDq+pxIz1emrS2omBdb/wtJLN2CdhlZsZSqyZ/CaORqZpQUMLhFDT
7e57/SyajslkTdOXxwlxmzd0ong6V+S85oCIZpmWRhPQ965lX/ZfWqJeNdjFrKJd
h7oOlYXMOv40DuiUqVY5OnItIj13FUpNIAlmBem3dsAopI0nXZhlTfrnPU4sf7+O
Ehh/x0cmtKjpqDKeh0yVcd3ZgNWmuCpW+8NDiZwhfEjdurdtFntLdYegO1h9ewGt
ss38ikWFsVpUzpmBQA5Yvc+8yRuMOqykjp7BXZaYlFpTkwkIobRiPhTWiiOjDF0Z
67OrfiIhz+evICghELEY5eKE0suJZoce6CX3ygPJI/WJbZ7erboY/nIw3cO0Sc26
xQQI85Cs4FS9Sw7Ove12SHGw5dtSOUNW9uQKaDGNKBISipUCmqft7H195k5EvYs6
UBdQoeUR5Fi5Lo03afJUnOkjAV6ygc1aPgnMkoGZ/ERxEycEHc1du0j12qZqt+jQ
+KwiZ2slZ2F2pbQyWZHXNLQOEuA9s7XVyGBrg2ZmEMpMsPiScqjO0o4mKFfavLlP
u9j6XLHOf91jBWFTPxjjx0siq518SNxotnLIIhMi2V6tJkfJ+nDpnCUPq5Qkxenh
I5NG26NGxXHrjFXNOEzHZpf8cj3e3FjzNIL9K9Z0MF0YchTnILo5IICzpSO8AxRu
C6IeQ5BUH4D7dGCEatOXQVKmoMY5+BBomg9xv0NxdHyDuiXP8zBgaDaaaMsEFQl9
t4H/+v8lAVv1D69OuiliEtqiwDgaTIRQeVnch9fe6a284Hl5RCORUn2HkHjZ1C3h
0h01nLh53pDQu5P5s8OFUP9+uL6kL33kv+7dh0IZDGmYNTHU83Ura/kZ98/aNITG
s3+9B37U4Oh2cqPJh8UhdIkYMj1mEyI8pSvuxJ6ypGPblJC8/+THACFFGZMVtdRG
empAwAjA4rdZfYAjpxa/eWdJ1ekioGbmp2dF5We1YLim31SPzQSUNxGvUlSZrK7C
iVeRFqpXFiFgoakMk2UPkziHTNV7EsTUfcCwF1tN+1iuU7lNCje8rG3n2DUz6HDR
/RyIDwMZL+hVq53nzYjR32qYtWCsCFRAflpld3rms/R7tecOsrIgmAODUyAvBYoT
5YdobmzD/ISGUcuFMXX3/wLWwY9OyJbcOO2Vy6sVhILq87SKZ7s5YBdzUxmEFYkm
XIaPhvAuox5CGQujY88k4/JxPhzuy2KN/HQ1Xj6dCYuYwlqaR16tTClNo0nZikzP
SG1z/kJaqWeuY6U6fNo1+0dxmIAa4A8D6Uo1+jkfsSup4ZMyFShxeuVwfJ+HhHJY
jQ/U+UrefCWKuyr7vlIlq5z71pI1ImUSwivU5O733tyyNCY8rlz5SW5XgA62oJab
Amqfu/yrFcFg0l+t1fQ3PhHOBd/vVoLFbcnDpKaeaiZqiHoHpavzz6cPq7FAPAZR
xF65TQ45F0W+hC/KxOPeNOs1FGG1weJpl6la0IhhQkbS6uUdy4sN8/P7P+lj1ye6
MwJZSmCEJiWnd7sU5zQqjHHfJgFsQsJeKNJV4Z3fJdCtD2M1wa6KurP87Sv3Fl7g
n2s03tKX0LVuarawRa0y2ecjmbGe0IkX3Tbv4imVLVJTYcTZr9AGv7vAm55cWqHs
RXTsyqQP/QsLH21iezaYOm2XwmMjYqwBxXOe6LruTN8Qjtgy7N7wJb2ktwG2VNYL
jvuI4/PtJRdapG5y/W8dwNYFVqDnSMlYvbVpndzmBLtBTKomby2Mk0SNeUYnTqed
/83d+Q1zot622hH9U05QAHtRlm99E+eSB7Vk6DdrZCWZn9CYB2IIgjCpG37DvhVd
4Gfm8ZzhQBf40rp4jyELlor3+WVsEBAzFRa55H2EXAe/I+OZ3w/pnHuTFF5SIc8q
alKD07y8UlhR8AmhBgyeg1O3ZJrtszLTM68LHK4k6kev9XxArfHY2FNREVfX36V9
mMI2vXhNcEB+DrGBCijkdY+10LUjut23piPm+Gs+XA1y1+hfnIZW4IG3eU+cRBTV
y0CBxaGeFVDktF6uweObhdpX5J2qTrLdXUjibSQiHHhgmHwvga+Mbc8JcoGs2VBK
vnYOsn0de81uFqD3/5luyidi65Wbqepmlf8j8W9qwBCo7CngiwFen31MLOrJwxTG
3oLQYYY4nDmFgyek28vnME/By7ffnGc4Cjvq8Rw4EUhlN1we+SwZoZ4IJaDF8fuP
3W3tPt6JZOOq6LEFC8DTryKmLmAyMWtihBYnK3FUPFy5u9dN8xxpnKHPq+8XjJJK
d3PA1f46qQJkZnBQ3Yf4ihI477tdGfsboIaHHn8/REa0fx0gHVW2oQ8UK41narOU
C/+pxISqaBgWckfheBPIs4oxttyArwr3XDUb5oqyz0dfY8nRF+xNLR/jG3b/9qGb
7Qr4zfQjn90i2B7MRo9r987++F+17Mn7WdkeNRzNAWwBsew4q/g0MoArOzzYbxkN
OF/iB1w31lH2sMzYJvygEAKvfXQg8Bi8bZ5GJypPszXyf4jSsf0lwWM2PKwp6CMu
y5FJ+6YA1gA70YBBdDSmC8vn3K9x+LlCYuzcKRf/5JOpzmONFzCuMlwLcBtGIpJF
Ay9sg3cGW5M3tHiDYkQneBpCzNcj9n6JTkiOmFGWtcU1sBLo1e04Np+oHAdVh6Z0
SHzjyaTVMDt67uI2gm8oa/mJtj6nUgrmfjrZn04s8VTE2swC0Ax9yKgDwY+nN3zu
58WnGfaoQByvHHtn72CTlKOrQzZ90a1a30N7Bcz0GPurXEWy9eAl4K6BV8TMpcso
ggs9+C2U2vrNRpzTFXijN05UxZuexiICBAG8O7EZ7+lIWW1u8846Duol0Nnsm3F2
6HUWsvkSdJmAvrKUXFrJxVhjQe89HqdBikEdpvI3tQESImAmXijfYsNYW/vgsv1u
cVsuR9VnL3LeI/oi+7EkO1UmrCb1mne61j7rVxJS/wPeH+d7TNbWmdeaaVQH8Skh
dUvLPU2fVHS9+vb5S1G6BrRRrgcoEKJwwP/+Pd0+QsZhh+u4HT9/K0jU9iuk8jih
xl0ab3+9JdQY1xiraExj/IoNgEzDvr492lJlmuywYiMeeLG1NWtKClsJkk6o1hD0
0QRMf0a83PjVh1Mwtz971j4PxGoJkS/G8AzZLptHNe8TRDQaNkWWxQ8MxoK4j0Gy
PUOb7P5Rl/uFjZDXfoxXUGdu74quoJp8vVzecdhvjXuh48lQ/5hCUagMAlsbhSjz
KNjhdBdcOCHvlbHLw5ioDZw/g4hpJT3HZFGaJt35TtSI+bKebK0vvn4ygqZAnQTG
4JHaMD+FX2lKrtXxGQs1yoqU+V+EEeYHoTDOBLJkY7grzsh5hFBUpRYYvAbOeUtc
4b+FXRqFCGH4YzCOtZ+zBawM/fy5mq2JMsCtqK18P7UsZaqvYtRi8bBN4c+sa9lu
oD4u+ffKy2CI4NPC7nR9e+VRDujB64p1+U7OAvyYGjqgXFDPfFpN5RwsmAVQkOTA
n7o1BTr8y154OqXP53vHG2DuLyoJNOvZGoQZJB0nEUtLibHOGqmTHa1fEeWj1JAl
oFyBjYWLmWpUR6vJ1/c1aiAIplfDcAxq9W3qNqV60DL994OSeDHpLgzOmyViiUCj
k/4ZpED0Rb5vVbI1lGeTxhdZh1GTDwDgB56M1fd9r97zL47gYpMlIU7G1qHDRrEP
0oy9nW5X4edF9hqHCCrebfgdLA/+OYBA+qbXGirDflD7mijwLJw7LeuGZ+U/kBPs
aiq4f3+NxPXzPtaFUUCoSHwB2JxWa3FNzNQaAdbuTdraWzkho5EQ1WUTWqkZdu3X
Sn/sOfH9rFMKGkBVzuBJoOYAcEa/qLzMfRvmYivUo5ebZC2/AtMfMKOIDL1nrQVo
rOmeMjWrTPWGKv+zcsCbmtvGFYym6u8pYd0DSuyuLCXHx5sNwWv2X2DtJUWQ35E1
UprZsMNQDXoWcsog+QiU0b4WpBnOGeKBKoDE/NOka0lIhMW4FoPsg0l0YItZ2+n5
vuAEH10Db2h/Q00qoZ2cb+ONQ1Z7x+Vr9XRmvGIRAAZ/E/3EPxkol5f3rX9MH79+
i9W4InpSq/GMaaFNgJWaQjTwboAcqY/ZmVJjRKEZ1hU3beOM3AkniNqCI7RJTeDS
cbMH1Nf2kjjT3y/7+eoOsBZEAsHd/qdaFhiNcpLE5U/CxnLPGlNRS4sZ2s3wzrkG
w6q7qDms8vq1dLFkFlMcZKV5SgHjCh/R1aThO5f2gPh2EubP90EcBe3vR+lSM6k8
DgAYN4M5W/EN1fxVrkIWZixwUIrB0TJrmHLa5rUrcRlZuTReNBnaQoA+6fnkjzWS
fb4WAHtjjYIwCCtLAU1PbFhQl2BkcvsnjA5LL0BSVLoGozL6rnPzUyTmg5hjqBhH
0x1xcjVVm2UAjMOksfJnSOx4fm7SC28s3CFHMr5h8/Qyc/wYk7cQohANyg7XVb1n
kGGw3C13RWamdQf76pq/M1ZGjuetQ87bUM8BFGiwtrLyx3gc2LzogBrwxC0aX8c3
2cs3GhrMTGy+33lLUEEzAjzpXgsUPY344LyovGoK0vUV5m7ret+EPDKmO3YeHZcL
/oQXF43QkGXg+vjT34fuQCOAbv+0PA3TR8mBQ3M4X+QXmC1oUaOa4N4rhaRCX0E6
IL9OJlFpZRzvyuXW9c/oQlfmZzCE1m2hLm2rZpRWoOlpHuMBqFoZZN81ZkynI5/O
8cBZri+ob5bi0e8JSPLjPeClO1VEBDEIY8iPpkaHi0mGOy50SEbQu1rUAwP+S+M+
y1tZul80Mj0vYMkE7zjj0Fd6FEqiUycKn5HsgarMXeqz+4kTJ/Gq1iQa+FBWEV+c
/jxXIR67CuBDwxfLDseyKVW9HO9K7Ymj/QHZdFW2YxmT1SwJPevE/elVHlVfvdMV
A39h0pZnxHxFRG509U/CNtmbQKnv4DPPHxwdLP+eXSRtCGEV5Lo0ErV83r8J69pY
m4kMUxKhm84KlXYzLlbGsN/fCcZOVN5fL6WNo7qfK2S+EL3mtUSSzKUhvpxyy29g
aLHx/zju6eb3KZ684D0OdiEfEcjJudsjUdKjxecAdiGSLPOwtnTo3NqV+Oj4yFNq
I9rhBoNi+53sBBK+f8M7gB0X2Ine2Xn4BPb/qPY1pGs2t1m4ePNzeL28IJoGapPA
9ZhvICR1UfetrOghfB44BUbFpFl3ZZB6g/XjW2mBHlwXniQhtCKxKueG0Yk1eUD3
1ewkRhpG+ZMD1fmwMMDD/qHH+od/NH/YuZv0Vlcd7sD1vop3BuYO55JP/xQrG5bW
RmBaK3swcJRCitQ7B+yq1PBHdAoymIDyPucLalyu4mcjyeg2qasIaKquYpLtaWwF
0AnjKjkwEm8wfShvffCiChI/hqp/NubcV+Yxp/Ewu6dGdaLV14GuiGVorrrpNgFa
vjKzXaJf6OrFoHKV01dFCRO46A36F4hpjD9hyn2wkH0OWq4YKRv4FAUbr1JRzFI4
2oxwlk5ofWVVXmgFGpun+4VO6VODpAD17IY/FTJrdnEbeVTBeMFWFmDxzU/YkB5s
MtThBf9D4fiqI5uWoPjggw+cEkwHSiUhFM6aPM/NXxl+rR/OS5kjhKkbaiZ7G3PW
ef9FRC8djwdHnYSYXokASjJBnDf8oebBS+fjUZlctBX0/kbkgRRwTlLyyuu2QjHC
Sd2K0hc2b7uCpkNfvTALrWtAi4zFbX/BinLe8ZEQ0QSRaHYvMPH5koY2vZ77NwEb
9vfEcVcPlB322EGsXOC28joANOcXXZ5+ULcOZ4Aoc6C2GFf+8lyxjE3j5ZPDTSVM
GePUqNXbNYtlLf5k55hcG77duQG4VGuJsKvVCUxQMhxL/N0Hsk1OlRnuyQqGvciT
iSryEfLugo2Fb6mzxTif7h2TrJfvW3ykr1AxsZsl5HavWzdsVNaZhWQinHmERqWJ
t/Jc4ylRG8tVHIWXfJJzUu9P3stQXrA5rBwOrj4wmI6m8UlIyRHIGXcmGN7K6hnG
9SJBP8nluRDPd+Ebd6Cy39p6dEp9SN3l7G63z/g4KGGsyTCcb91NlARyb5hQtQO1
dCxbG3Fi8eVswSu5QjJnxjJ0yidBYFqA32LZxhQcUCjlkDbpbWQSXZOLLtTVq3GU
n6aaCOFwUcX/XJkAQF6OosgNuTzi3uiAfUscItDRgCStnWHGKKWZP1oh64LdPlZ8
lhjOwLTbn8b8SKSuEUlJZmN7UL92WzmjWx5Uva3XPFjEU7qo18KxcHN2zaZRXzsc
+Tvc+vK/lSCA73ygXZr9VfElelipYxXENWV4A7i0QNGRTasD81G2a33d4/agrz8p
hbDf5VxnZPYLuL7OGzzRf9PBUWremBVtdQAyHkDo/gNklPj+jHH47Ejm+1M20tWX
oeHOcZVFAHCcRIuerodFqla9Z9YUhn7XjvQTYuZcrxk/KpO0qTJ8dwqt+ge1+vR6
AgdkgtG1cOSQbte2PfQmWeygB8et+OouALvQd2udG7YlG9pNZcoFizL8jonNw1VK
49Nr1xzRx+HKNJhnObQqTFPwLqQruWMeTokJHjbyDpa6uzGyct0qNNrphSNVOQ5/
G9p1axe+1TyHjDHB7Tgf3CqhCv/0GsGDbJTzAOL8boSz1K+zWzszP7ZnOtEG7qJ5
IVoASXLi6hdTRRCVrHaWe+eva95Vmu9nK9SKCb/C/8ezBy+lOAXTArnnhgwHLvN/
McdNF/AVsJnZSV8ATqj+ybha7cyR6JUBMZY0NWgLSEqqif+7N3RP27dDPxkjNwKK
AK7+2VI8Ccjp+PqsP6NwRFp3XaLCJDZwlIo5GE6tazkCBiRx/6+1pmJ/iSS2CIbu
R6Bl4jZmR8vvBy8CkfhTGpN6PEa3YTf3VkcUjH2GKtKJ86ERKmH12UPqfIoI+57K
VdDAIn6TgqiuuMrn+c2oqQBZrc/9/fUr/P+FmtgEwiEWw0Q9jFCg0pdXcJyXgOaR
j/H9YNDk581n21X0YW2bUrIRCHRxAMx5d0ABB7TEHbpfinbyb2abyPq/zbleFpaQ
CWUewD/u7lIMk+I9XR3qVUomjSmc3okqiPR1X3pukNIrSgoeuOUzaVhnx0k1AijO
E4gs+SJn3t+GO5M+AlNsjp/xRiwJlXkBpWlr3bFST8QDOYnAzpQ1/i/yjxZ1+Cop
Cqp6j1qhid1Npa5coOFv//IvucuD/G4Gud4htyHE2Ta1IyF2LoP8siKNIUtWl88H
11bwebbqbX80sstNfGBs9gtih8J0F6FJp8jddoVE2/jgaqjtRM/NNZ2HyMQpOnaz
9q7eESF5bnY/Tzkw1/lsjp3qGT7x42hQNigWTOyEE7CCTAb+ZOaa9LkTLoK5lg6h
lohIkr7FKvksXwMEmSZlhDsmuIzrgXvK4kg/+9yqaoz8iCCEo8PGUkj4MnUpZ1tj
zfvSphgd2h7ATjzYCQlbTq/1sYC+7OoOb+wLKJAGJSJFOL7IxYjco66fXv5bFVhj
SFgjfd6mYxNOI+/ykpKHkYBEzifAHrlgbOU8pcB9+nFVpW/U2fGQT34+vCHB+SsE
tp9E6yuRPZGr4VCSKV0TLN9QXe5GYYVa/eEEZifxEa1OI8DBZM20FCjz7N2P4FRB
UKa7OobbVdJHVWvvXchip0ChXqNAd4M6dg7Fb7tINKOTmu5HuaCIf3kmR8TqOkbR
Wh2szc3wUpodmscz+16Td7mpKk+bi7FawYo8mFMHIdPAa/kc2wDaPO3LtE/08XDV
dLPi+Z+iGvyQ0zdLza70Bu06ky4gOOTfpvKDA+4vRq1wA/SSKMwrej/1aJhEymzp
Ygc7got/yifBuGr+c8XZCel65fjOKBs31gCwCx8eR9s0W7mgbmXsalfI7XPdq3dy
ib7C6F2bc2mbGY2iFj1JxvE5IiBNtfRj6l6P/h61fi+IbHNyukQ6GtkM7KxWhTeM
jTOH5PLWzjc9ZwMDO2o/3FMFXhZetqgtjT+YEz/UGsolVxWJmbvi+9Lxy8PW0swD
kZADmLTDjM7dYimRVQ0iAK98rbUyezq+A+EeAVTl2jDhj787fLIQisXfaWKdUGNl
TNXQPSD3YxpCYXt7Xl+nYyH4HqEefVR7Ye+ySmJ+c4hPj+yqcdfms8QfsaRttbtn
YzeY0QEiYjVUNsKHhIASk9vfgHXgVc8l/CEb1+pGs2BHc+JmwBbp/M0JBxYcsy4+
5pyiu59muJS6LP6lKg7xXOBUd6xo4faaKxPckyT6ZHagewt1CwcetB/p+wNPSesZ
+pt8bolpyHs32Yxiih6pUA1FeTVMGB3fzhutOz5AVaqUfuGVnA3KieMcl7Y1yVU5
Mi908bgSawcxg4MAO3B0p2lGIC1AzRmiU7hDQMQ2SDYA/b49cZp0iSZ3A2pOrxQI
io4vOIUaH6bzgjQUl4+q3HImo1LKIOILZN2BrZ/5gUrdCYz6v4ZsLwo979q+JcQ5
+gApoqKLYB7XMIXYulgFpPtVITBDVYSkkArnJumOxBVnQLcBQ+lfkx2nkDNnZyhu
ndmLJeGFTF6OCcqOEP5uSef+YCihvju/XZ2R6NLedQ+dsGCuW6+dR6FgW/R/8QDv
u1JoKfIlqGGq57YGJuv05TSuE4nn6JxLhh76P7kh9ye357M76fg0RwIsLQcQlpPh
gzb+I7JcKToUZOQPp6FB0CSpQA2eZFitMnMEZXq52tSiKu/UwQrBekOTizSw0IsO
Um13NasaEpnAyWbmrw7nVxhQIzPMe6N18yNeZXH3/pYPdHGqSQ8p1q3Q98W2SYYt
rAJBqMvlva4PB8fhiD0mJwJsG+5l+giYHHeiXBXx0jbAM4n3ErYnij+5rv0uIRBU
DiJmHlYDUETT4Hz2H5idwFXlMNyZ+Gp+cBggwPZQpnezbe/dzDP3inTD5FufMPDt
VLGcDFjbkzUCMO27xDUviXoPH5zNUobnSo452d2I19UlmpyMSKm+V1msvWm/1ux6
vwTX1wuM7NzLz5if9nDB7qhvaSz6uczA7a36vh21os1B3WIV0iTLg/xGJXGVpCaf
fFTufhntyCw+drhkcHG5dKXqB2yiSJXx72nHJgTYMecNM+TZlX7iFjt8bgYKRh9s
Rk9q0MPUkTg+48V57ZfIgKzW7aZVNibTrs3ntHyR4k9L2o5I9G+TLm1PnKkNtqa5
TRxYdqluuzhuJKijIADCg4m/SenUOmKFnyTAy5giMl1CzQLL679NBiwjkHeYifKy
8PQC2pnt9K2h8xugDgPct1WPJUnpiJW0ccLhi25bL8ZoQxkCfnm/g+NPlvr8Y/QH
h/ko6AYxtsPU1WZpk8oIPpe+jfwTvLkxKvf2xjXBEuYedr/k33U/zTtF90mlMK8b
wdOC5Jy8imIox1RVICOkLuiwCr2zCSUK8wRkg4Poi8M76HoNnmuIQ00PiDiHQKF4
IFjBuHzB0N6f5EOzAXV5NWQ0wKA9JrPUC4bZiq4CTAVee3kmKsQ0cYeOMDqAbQVp
UVN09G5CPOw7GCvPZFOMnrIY+2fE1hP6cXVJsvFBcqcKQvGYE4/ikwT9iQ3rFNeO
1duc5WE18dJZZpnB3yrEl66OfZtaUMdtXoNKRo0ra4Kb9X2q6YWr2eHaGeXOeWag
WPuFAWVO6v6dzDra/tbA5UWzpi+tWRVWCy6IlaUsLXsCb1AZZlDUDq/6M4p9EiUj
Y1o9wCunqF3jfBeZXULdu04JGB8m2LQI1tLIRhB3Zk6qVPweoU+xJ0AHOSVY4zZ6
MdX2nSpaKAzgua2g53YoI1/4GVqhCEVFWfTNeD7ecDutLMpV8Y7gVqTrrRlAE5uV
F7t1ZbijksL5dioGCdl7D4OcEoN47w8DDv/FzzzqO8QgRl36m6atzlC/nGa+GvFk
UYPfw7Rfwaw2kwiPuE5GX/HJtRS4mKA9wd545dvooptbJd0/Q51vMpFtxiNTETwg
8U0Sx+OFixnhH4OK0DMKS1dR/c+8BS0jn+BQAZHu6Chtr8NyOQ3jzLMNBgUzbIni
iIW4nHRADflIWfOBOReFD4kuZBhipv/0cXclSNPeYb9RW+fJGNLnrhEpb4y7ph+q
KQo65SxMHJ+V/z/plaGI/Qbvm4e8uIg0eV28LOFiTBEg0mP4om4PZM0lKXhXvwHB
iTmX0cLR4RUVWYzjfEo7XaOsRWCd2GNJmteDkgpOp+yJQL/kafNZ1rCyy5RhD32J
283pHYAhQmGEHGo/9ogNQHv069EECKzPOCKKi6CffSzgxyQq/a6ZBCJwJXoJXWVH
bwRFUh/MYD0ZZKz17i6rKpmw69SM5M0R4uOcb9Hg2hrthxJoRWgv5/gtqcw7wBT1
aR7gMBwzaJozVXYr0ILsyN0ElkSCfPQcIe/DiNFmdEk3kWCRn/0ri61LvTc6RBru
CfKf0SE4/hykCDR4W+eS/Tme6BOKthMLRZEMQimIITupYDrr/L24R1DO87Dy8rwV
N6XxnNqKRpSbtUZ6iHZQXgxcBWLw1lz1TpygldIDPBwySGQclcAKsdP+xo/w6Eua
Sv09YC69N7cOEw/+19WL22FoyKyq1mA6SD3QTZg4qmCAouar/sxK7f9RhELxkbIG
8Adbbh2xvCpOrUA1rh6sfNxXOpzAl9/0xHBxSfeh/vnnKsNSptZOiQ7nE+1IRE9a
tniGTfHJnaxhSsCn3iko9RfyewrE7ssilwZ5Lp/uPt6sGgMSEHsHET0ZXnzfz7hR
u8MnqhWxRKY+nBuXQ1IuYEP+uSrajb+Mx8iXMtsF2YwOIdAO6vYuFSeFlJB7s9hP
JcImcWUkipykCXcg5mIRlfpGPJ1fimBvp2t6oRUV7XgsES1xEfy1OXKXa88wQ8f5
La2UFWweDQX170Y45uL580thErhw1S0KAnyyVgZKPR9mrNuR4f2EDcY0330R5zq9
67C5BJlbREIRXlWUk/6sCosu3xgjUGo17YZdnkhVzVdSy+ElZYp7bBF4G3olMLLg
okl67ocEETYrGm0awi4Ih58pMTaIzk7T28IlDiqHA84onjhVFAYSH4iSkHdUMJ/5
y+IKP+RXgYlpJrqLgwsTP9cN1cBefkqXIItC8glJt8jnZD2IotYhbZWgA45AuNEn
D+3Q82w+Unn9b0AHnBHu/xyQJTPHYwyQz9u+j8YEdK0S7XTExeer2fqGR3RFGIcw
4a3RRPd6e607WhkgBLhIrz49KxDZsF9CMKlNGM41L0e9DZudH3NFGY29MtX7a+wy
h4ISXRlpPp7VvHiUcMZ+21lGi5zlksFyLwFBSzSJcvOJlCpM48rCSj76/2hgRAMc
1MysQbjoyyALJqN0HlGA783GihSM++D+YO9VCAUBliI6kf8drdQesP6mLOy4gtRE
H+38NijoMDdRLJmp6leI8iQgnkcvmSO8K9IIUZyzZYnugpcrPRyPi0JzLSKCD62X
dvxkQ6jcgRrfE8iUwmAUKNtYP4TWBJsRSbx2iwXPQvj3AsKyKsQA0yN0DPjlC+ui
ByvvOGgd1xeQ2Ny7h2Np1w==
`pragma protect end_protected
