// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
cN8iaaD62ANq5SJ+0W0Fq57sVgI0mMLObCviFUCUzdNhw4DJccobkgc7f5MCzJgu565fGlrcTfdt
5udLmo6yu06n2AZFCUF6gRZZIg/MrQ9leFCWcdNW8hfYOA9IV4tFht5LabmFxSd5hNhA+Rp3fPDY
E9aasm2B09eKnNSTKHBGih9dBbUt/PP+IRnb9wJPFaPqTe1AV7EGDKgKOWbImnRLQsqx8ifXfwY8
svT1VPG68C215JmMqRnJ4enskHaaNJzv+QvAHTbdE40a43p/XUkLKJ7pUxbXgFMe2ycbZzMoHivK
hk7uoex0nVbOPkMr+B73V1qSlAkd/DmTTEZ5OA==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
KogOOEV2NbxBEDVKiRhnlbq/Gci7wl/t6DWaXphYZGHZbwWlco2XHKubSZ5DCUvnX8m6iYBbPGee
6TQUzWiIc+Cj5cAMGONvw9OXJZg2cHCLFEJb+IH01WpW1s026VXxSJ/InbAZVG315+xUe68Fer5l
7RGkMK5A7Yz6ElzzM6RcJg+0CBSdX2qDkrRe9812Up3rqtALb2J4o1NEIrEH3KdNhZdCRLaRGzDy
FecYN2re0nboEuP5oCiU/eo1NgDlDneqqwYotevbD1lY2QiQwtAj50eTKwZFkjaGl8JQENtOti8y
l+n5y4KMOz9LLkUlfquyLc4HGMD+VqPz75TueMqpYqj4MaxRDpbdCCSdVw1seoxski3If6p5rQBz
JfzAGD7FAqcBnPbVK+hmuh5iCmWyUMxs3uwJCxdbhx5FhrsOH4bpbCMxUyHlripSVZ4p1qwn5BiG
Doead36yM1/IuDaP/+SfAw3f5MIpXVp1rxmDu+GKuviFqven9HCiHFzVz2QgAHJeU4suxgISXdNd
O9VIoQQWFkUlVpG/JyGfJ3GTkC7nt3XwLBFTF+ub+n5S5q/hlEnibIO0ViLJfaSrSvKSp33V3t24
+bYRN/ZfgE3GBO/QyXMfjw0AkLwlg4Ap6uaAfXojCalTj9sDLiHWLH1zYSy+QbRGCeEnNl5nAQx7
0NS91hDR4ck6fMt51H+SBK2agaNNQK9YKU3VmTCjFLT2mKfj8+vHIK69zWaT041uf49RFzNdZrE1
58Erss+gPoyz5iXj32ihWlz4axGwm9AzdbFKxPdfpkIBqzbZRQonWF3pJBlaHFUzYcbIWIs2kqmj
Qty8Pm4ynmo0qhkEKKmdQX0Y1si/cctB6JEkmwz6xrYQFLIIfeymy3KWXC1wK4GLL+jL9739bYi/
h9dMhwMb5lg4aUiASZXel3X+arV3f3PcWQvUfjr52lZNugYy+zvJzL+2EDynuMPf2KIowYsa/CKI
A5duFkZYVGrTPMvECkSDbd2VCAP09myNONUY+DY8drXJ00EE0/jaVdUzpYDQ/5c1Oy6XJ7ODBSC1
mqzfvwc+AA+AMO7ZgsNho2ovK+y3MD+XUjtxZQMsHVA4XIwB4SZt9TnPfKzO7IkhTPZJWL2U3zPt
qgxo81ysAsl397z5WxdoJTwHLJsPVsi7ySCogmZETmCe6U7inmxbu+XpMG8tzCWZMGwfdEQk2A6M
zDhuWWOZrZn55vdR1cjnAlPoKpVn5o0CBRDVrXw7Y8uNfHY09TbD6Vlk7GL4ip8EDbCm41zYVpsd
kOZZNjErSPK8c1ncf05SSPHvaGKo8pMb+nODoUSXHlkoWXq9iTRiD1L9ArClPgHzCsnwe8QtwzNM
CFK0VQ/wawXAJuGYNNpw4VnXln0TvR+oxTRnsWNUvbTbUqT9qOTYxszDkRWoRJOYWvGbN4az7V7u
4t0Q7lz4EM6ywOwbMNHkN3tagm01AgCZk2Elqikm2sKcY7snusiTvBXpKRstbRgrRWbtx8ydjR9n
A6xRZ4WlBskTYVYFc30KDbkXl86NAwRlIhZVVA+sI6b7XwSoJnw9lypsP+oS41kepAB6H/OK+G97
wkqNnWK39E79TV49YHg3yU3+DKN6OVxchw1DqF9U0NHf0/FI2WhuSZ+bsoetoqijU3q68eKwuzsr
q3pZs/mjqSizyMozCkAmMBYQ/a/9ySjvrnWSXbeVGjqT42lkR2b6ANfroJYntJR0piATMeRgTx5r
7qQ8YODe3uLwgFMz4tttLA4QhvhdNMZMLziiW59IS7vt8cOw1sKKpcuIKS5BV5SaoFcXVC/1i7Du
Mm8CROh26qWhkeNWFcQDqsMcyay6hafMKNh/3BhXg6cbVKD9T24/Xix3ZIcxUAZ/FKCuww6kKCvU
Pl218741nLU3kZjd5NA1hDCelFFyMJAINQIoG1U5kAkDeivx1B6ywDQV8jp9vB0/q1IwM6DPdxiX
KQIZw8F+R3iocABVpLOcbPbGt0GljrnZB2Jc2/0mp53W0wg04k4ZhY0stJzZpqSpBj/uejBF9u1M
B1W6q/q1YnTxmVu5+oPE0UDIPrZ2Ed6o1apa+eTIO2UdQi5kvnCx113A6lfA9ch9AbjVlbz8TX/w
GPZSU7KQmP6hyoqSqziIWn7ykUEPQTGAmJBNyZUiKAyjuS60W+ysSM5C4842iOqqPrfsppcnls9D
YidVDynN5bTO1JRpbJFwJ1NmYybzjgsk12NwclJPGo+doRCg+MnIGtRjcd01fxcsfxocMcciPyG7
FWUO9llZRfA//SC0wJYCazlVX7HD6Kdhe7nt7O2RrEce5eM1wet/F0z6S/MY78VJWYcNcYdeJLVf
XBsTHsmOZxVc7D2bt+kOdAdfbtKW9Xfnz85iwWeLrz1ZJxr63XU/16JVutBaZOIPeILTT6rymMK+
y9BHlT57ASy38CeQpwrB9tGO90WrrcyfeAAK2nzmvlkhqyEsOdsizSkLlTrKeHDCfd1An5VudwuG
vbdVrVbV2HBPeU2m0g/g5DI9V81q5obhZVl/Ojdx3GsunUdKTwhXGAiRJNvp9bXlFJAROwB5FRoa
RrEmFdiC8hf7ZzugI9QHm9nqIY7MY7UFFk5WuIP3e0wb66UHSJ4kQCmrhn228uhnMKn1TXyKir1Q
JrEab05cBiX1ihc/2rewFsdrgMi5ATgrhMDJdl+rkDn3pBpV8iQShBwSNxKy7oTH8+6h2JPAu41j
62qrvUIoNlfmvZ8QwImwoNxqoNMhh+HwHdHe7ufC5V3A0ZJNunsTMg03Ql2XJQmoj/trFT4gHy2H
nsE6BoPV2IoBQ113T8nDbKIpnsvtS5qUCWCEyaC9g+CbS7zzRa5EsUQBD/VtI/zFj/K45DFDTmcW
1yD4b+k4/EafSxuWAk1mmzS9GcHv282jKuVbd4BhuoS9XFJ9zHqekYf8FTYbRig1WORN9foj3oUR
bI9fAso7Mg0vbp7xRy4G6v4zUmNvtc6JhrVpa+q3rKPEmgtxeNS9V+bpHW/5+4+2ykEev00P7wNe
SgBqw91Q+FYVb/JQvKy7zPsdjgCzP3E9xrNkTvqQCUIgPJbjtz/WwChju9xO+2Xj44xgII2jz1zT
mC2o2SGI9VyIniGlEFKxerHTHjUYn3MuvTl9Zu1lEMitbCnwFgbmvzcvBT5639IVA2gE5num40rp
AlU1t5m4O6wEnIrKkBUBLd+mL6i7p7U2yaPpESuvloROjYP4A3ZklOfuvyiU+ndWBpSDKUXLxtF6
t+0R0NKsPpP3Oj5WtiXLvs3rOra8iDZLDwIeVlsv+QBqGMqUG77BSSrKp5mnrgIGmR9k2l2yK4tm
UVbBbxK29OksaCErIMVssZbNYrKL+yCvNM4PZsF8JcoRQ0DRBIy+nSECCZ9iKj2woctnsJHja2+s
QQXBPEpV0v6bkqIlDkp7ljQhKX17ocA9xA7nK7lzJd3NgbLHLhkLaD8/AokhK7HZOY96WgXbc+Uh
QlW3qLBjsG2I91GxEsIaUPpYks2iU6knDTmQwkFKnNENYYYNLcoSZcGh4Skny5IVRrFYnKgA7tA8
oAkhdgxKEMubhTeTi7ygatGghHttftv9BAZn5BgAmlBnrTn25n68jq1pkWtMPviU8/iOdKqxW1P9
jlu0ZSfeEt9Q8pFYkKCckTdV1WlnnsWXmfK07IIWaWE/J9X3inQSFaydMbuu9gfY24VNbQCXszCH
EfvuFUX5Q+whBwnsj7DhklIcWOOE1XrRL0b2NXqLxfkXPtLdLM3UjuUY7l/ZOwXtcDU9RmUQJ/pG
Tm18qycMCKFVEXwQNdktkNnC6GHnhOQhBzF9D8ntEJuTuIHAqnFcUFKSa7DU5AqtVfh0z95Hgdgd
yK9woA3tDu8vDwifnj6C+6dcWASKfTWI8Co61MvRlQhNIW2AodbM3/j8NOsA/bvbqwp5yt/kWVqt
f1yfh4wjqrgeZEVbCAobdealUkXH9IRuiEu4cdriV++y5N71opODIORoDznRKG9NASBoH1YPKi4H
6UkA9ZZC/rXtvOhxtO5ytNTZXOfESkJ5rxauUK64GU6n9XuwljvUveQAuq8jQnF84JxRCVQsF3i6
J5pCQYrWCzRWTdQTsRbECzBuFnHa4IUE7+6PUOeleH7/3YdBwKgZlL2fjy5O+bCA153cs73QmyQ6
4SVdoZ7KFhPs+FWtQgywk2HO2gSaR1f5eHNyzj2vb7I4LF1rw4oq1gYo87RCapKO93d6lGKyxkry
Y8osJQDFoF4xG/GLL1Xl69JhWQ9wbD8Htf0x5YVxXVgLf6O0COt9c+Am+oYtqhXQHMRIsUyjA8zk
F3aBBIgvuhm/zY/MkIwrjhfc5Mqs6NKojR41B0V5BYkkZjHQ2FypmJKs6Bh3w/O65dyjt9GLaDOo
ObbkXKDoTZ+9RoiKO6BPbSJ4416nywpH/+hD7XQKTOZk1lVZ4SiOInXrgQ980IalzpSSrNDLLNNx
KY1dOY8dnY0bZAuEszAsza8Eo+fn7/di9BuOjHlBmItVln8b8Qdjvtumlr6ZDd1vhYIcjHy4hujo
c5bN8rustNgq3m9wA+ORTheIfvTA/LccTrDUKZCoFrVUUweIEmmbhQFAWrxzgRAS0wM7kTUAB810
PnKhJV+dFwmSxx+6f+yvsCG1fh+gLtpRkcIY0VTQQ+6y14BMBLN1XBGZqsCHY+F3UPjTMfqngHud
P8p8RZSP6mri7X2JfOpHHngYliKxMDMOY6BWvOogHXMJ/duQ69Zt5KjUUi8AhqbXjwtthNxjDKTA
B6mYsny9cV0FjBFinqmw9OiEVVb2daimHM9tOnYXYdEM1Je/0luPkuJN366g/V0gbskSZY7AkdQv
3BSv4KJoe+/YlXqgR4/mKIzj/9PeQwEe2Pg7IgctprxH+g0i8Wk0WO2eHe2KBMEv+8GjyS+omLWU
BHNp7QK/e72qD/2V4N/ox1snPYPZvFAoQP7zwWqllnqJVcmEYhkdSlfIKWl2ACzKWkWjbp32jcAI
lTqjTgOVIWXLvA9Wb1j6BXVMc+vCxzGi7qOeOlRPfIBYz2v6pxT0F1CAFbx0TTaDvth+qxU4sB36
zWXwanwq7OE+e544iAQr0lZmGqRj09aiy1ZRQ1YLjiPx9+WdV9uDlPfnhg2EsF9genFNyxKFkpsi
TGKkTwzvTYWApn7z2dj4IROsWG0WOkJ7iGYtBAt2MB+0lLNSYpTIOyK5MmUd6DbH8PJEX0UubUty
rVHPqlFtgykM61HZUWugZhZ+yN6rTpVY8n6O41Nikc08LGq+W8qg1bFVWy9Ay1olrMHy02jWH0qZ
KQ4vXL++oo5/rdWjBcnw8z6ke756wTQ2SoZ2QuvJ0bFUJE1Tahhq7J6ffQqp8+uIO9hsr8eWoH0f
S1AqvbP3fOQRKfO8KeQEYT4h5FiC7KEB7W7lxwzuU4pXfH+GHUcpXHXQHN+vjF+BhwMmjnv91+sI
CTbyN/08hFC5gAzaotTXTpfvWDjAiEbD20RxXx81pIB5vWnd5iH1jWIxVXzmE4oh/ZkgaseWUn9J
mIrxnOADU1nUNLNt+Xcz0t65+tBBbtDyMcbL32JWtF8WWVQjPHderqhQq/tt4RCn271DmPDno+B5
TTSfm8/fr7yfse9qYS63TZm/NlXI5IuLcuCjyfnrVwVBe2UvWucG9kUbPLyzUEl/FhAI/cHtwm6p
a/9pw3GWRBwzgNMDLrIN+1/F9JW5Fwq5/Ktzq572ooabUa15bDJuhHGzVf1mnDQPECbhvz7u1N+R
eby9GRzeHsTik/kECrh2tjRK8tQstYwaYgCmI/+E256jXugTQhoN9UPrDkBXwKfhopV7JduBie19
LIW8OpMSzI67KDBR61B6qTLp2VKSov0WDWyAR/H5pTCiTy/HsC3nQaoLTghj4hJe7vNfPiky0HvO
JNquW9fbVY8cb2B5v2r9TxXZGOxAyOeHkef+2xI8OFmkCLORIHBWoxomIeG3gCWbj+kzeukw+1tf
8Qq5y8lgm9vh+9etzt7U4vxz1jPFPOFTRRywZW+HUFM0RhitjHaMMbXlLAic1bH6IysymsogQ44m
35z6RYkseBy/2JqErWotMc1S9gcjiXAV1fPiAT8XmGe1P944ZJrH6B932OHl62sQu0dak0zgPkMt
GB/PnTB1v6YNuR10ZgJH7G9sCLhu2KEBoZdcXsvQrjy+N7TlO2Y0+YfexQLuAWTdcH8nN0YNq7Hx
oJmVHGx0qJ1Wu1ZG8D0oW/eYYWApAX5g7Tynw8IyJ/YEzN2xrbW6g0WvBhFQN3oTJgLrvmHwAxlm
LJqyVAGCu4aJ4eaIeloq5kuy9okbFD/z6qQ8ng/UMWOngE+ql6/WPtYB0x/wOCVuN1XKs0q3ACQe
5CP7nlplg6hqmkSxEU/i72lfAhpbnZIjsbK1S+FKpMvNeo3WQ+5qgdHwrHhJYiFayGXnvPZu6xwB
4G2bQChKVNk/b0D65HKUQDIA37hkdBVCD/KVznTeSMRR+DTrq9HPeKV3gnsglhztI9MqlXpVtdTp
78MvGqkVx1Bt4PSf9de2epZsoUe0DdEMNoIrKy9OzLB6Dzy25nZ7NChxyXgGUqzP+tuL4u8klYLl
K0BLylK0firwrbQ5HQicg1t13+5fZyPHvkJ4TtTsAXdyHfGQsrRNC5yxf3xu/zqMhk5H4fEkvUyA
yXmVaBgea/ILnLCh30me2TYSLVaQhKYkmObVy9rr6MrOGXeJQTfBybanfmSgS0Ciq91wTcCkbwVI
gOwKX7LOAQIpVJ8PNiifzYzQ/8OusrZqx6fJdlTYlKQxHIsG3iT3/5tb1AS/jtrxfVu5x5nTIatW
Tu+z7GcbjeiztXtWOmHR9uqbrA0wkqx6+m0t4WEYJ6rx+grHlNSNREDj27Oq10kO0zF7mfN6E7SQ
3l7hnLx3AZLyovqGx5QWU789uRzlGyP0Zr6ajvHBrDLbtkdvF4EQgwom8FW8YLUCVkAZDGz/KGGb
MIHfsjFK01Qksy70c2I153aSLW9d6dqt4GqHNUxICyGjxOzRFv+0uH3aA3naijX/4qPNkTBGRhsb
Z1c5RNg8q1/xvuqAp1K+DQJdzc3+CZivtpBp7z3f/476KbeCaGem2FEZKeOgmDZtU1OPy6Y/Igpt
PJGDKbS808okvsT2fOjz7HTuTvN6Doew2GmPr+yULOsXKlYCdii2029xzjNC8i/3gRXddIzTDAnb
gF9xE0bir+F6y262e/+CsRSNti9eq0bUymh4JiQAaGjJpQp2IY737TQIo2lPbWyc4KN4GULa6ZBX
jvVCaY1bkyv2fJXHlR6r7qaGEVDtPzCe/mYEtqaVccJHJBfqHMi5MYACldYvv5B/muk10vGIZSsy
kGt+GksU+xGcwP3FaRYdCNEdz76OmTn7y7tkA7SPC7lQ4/m9Qn718amKY8iDsrjoesp7NS8qG8US
uy5khsFDDimDKUPwkfC0o8xRhM+6WkZBfVTfUu0FcfDOJ93NNnq3A97ISkIXhDMlVDsLYe9Bz0Ge
swlZbGGuz8wwg+KkI7tNj+UHrJa6cWU4+WCq55+xOQXnv9oRNStkgctfKBf5Do4SCUJ/I9cD6l26
qlFJcHObsYWQ8YDVT5Jusj69Ml48gCnrtOqtumvEh1OIzdI0bN6j0HRVbH77ifjo5qsCvXiwIvb2
oQZN/5Qi5U/YPjB2gatdzA8c9elJY4i81aV1DBJ9fN8Q3pXfbjhvT9hnXMJETVXd3uyQo4rjTLbA
4L2JmbJxIb1SkHhZ7Jkopsrd69PZ/rFh7GhljJj0ZVp6IpkikaNvn9wa3hz8CjoeQ0f+Cyw7dPvk
74dR+vCpBfoXeD5sLoeq1gbKKzrcwzWOLrWz1PFSgAeBju0wrQvQF6Y8dYyYmF8eurqxAuIb4Pgl
mb4Y8mgmzA+xSCvNH+K7q4OM+sNG1VH9LARmqP3Dt/PyJl8TjJdge8ARQL5DwCuSsAeS3uP5w4R2
vdKhC+vhdgyLrg+poJznzt1NEW9MsILlB9DlECGeZzJZiv3pdbwe3aviFEwL06s8eLrJQw9uOSWd
N7JbJSGGQgRF2ED8ZAut/s83bLITdI379ylmLJ82EbFKN/ChmPNSBabcdEKcvISFbI7S5B9beNa0
aWeq3XNxuHo0WwTjeT993d9T7YjBHA8HibTPY9K9NhM5rCVU+3tuXDt/19YHJTSmoR7vNxAkdLnE
fFyqs7fc8y77ZdNDAiUonLy+S+2q8wnZ1G59y9xeiqRMmXK095D4UMfLmhEyb30ES2257nFzcoLc
aOELUKXrY6weYDdzepYtp0z8OoxACzuO6RcygRyrJXx1hF62XY+8+M69UtzF6Qf/TOIxoTG1V3F+
cgxo4dAUZQeBkHylIMZILqZYpa8buAv6OrcHk718kh7qba2sRho1BY79h1nEFbJpJa4t/dR/wnvV
0hh7KNAB/NOhtImUx03RTCsC9UXaYZLRcKKTg+gABXX4G+s09UUJUGfbvG0oKaUOWhH6UwPZxkd9
ofYQeuyySr6HhThQrYDfH8cu+/+4izdlEcwl2EeVMlEF3hCyA5266DAL24aqpFVxN3cWjE2zA/o8
pj5jhj8GyZ+09XqUm1aCCfEKjIAGCbTVvvhwg1c3Fefj+9/tP6/tuG11O9cgncVD2zQtpSdBvELj
vWKMJJ7+tOla9iVP2bGDajCC4skm1AASxwLnsrv6VC0B+T720lGaMrf2PfWu73wRbbgS4B3y5W4f
wiMl6PM94+0veTE21H/4QjizMyg6uKQHXWKIqZpeC8zsjxMxm3C4LD2JQun/WhS/MsqdhMf0cMlE
m27z7ni6g9GwV69whDsNiIFr4GSjUms5XHAsbFx7WNAElER8l4Tq08YE7Xp+4Q/CNUuUfJm1QMK2
+lPCQIemjriSDj6EufDa9NXTLJcxc+keWkpBLCRUtfF1iv481lZsoc3OHrvss7x7nXE/ccVQbnjy
hso/HR/nZXeu+MVtPj7dYQ2SCWMCt4+54337fxbMQ3ho7w8ud7dsNlj7qjs6u9sJgzyFmi5x7SsE
S4K6iV4IB/jKQgP2bnNZgvciEvICMAFfMkOnfZigEkJ9JDxEfeKLdn0m7sLxmTWkoOl7L+EGCpG3
iM9ThsQBZ3zocdgT/xFWmR7mVStrH1rYD5gMM9saB/dk/0mX7znBWeGUIc2cyupHl0HWvhbCqKe1
QSkXRa6oRbJk3vbJAHV82fTnp2kmUkM3esf6zpaofw15+BKSTdHDWMpSDaOsDYXmHwPqlRyMy+Ok
hpNNFzQOJp/Q8wmUEpjduVB74WmYby8+xz9oP9fqkOJNui8XHVOx43fg3cS/lsqVn+zUTWKGO/su
ELhk4CP3UYvhlH5DyUBdPxQa0hBZr9T6kZWKRoDWsWudTJO7mz51Ny29gSAVoBavkxWjkzgS7Gz7
rx6meE9pdyxg2x5c+2BG0DDQSi/kqk74MoOhzehNgdz6vY/6YlCwZrJHK/ynDTMqgC0gwcqKjRTa
dOL5LkSVoU0i8afw6sKV99hTnM4zSsAPqkwT9J54Hb5yDoy95jhGwJJMgZg+gh64sXh50ppmuIHJ
ef9AJA8ID7Dr2AIu9CRrpk3dvWgKIVryqXepuak1AxjjHnihgYeYM/OrceyN+bxUigA+v9m56hru
jsrNCkD8dup0XwUeXe+SdUPnXgJmmBCd/UAOcMZiEPRqbxB5qlwHbuoDq2V/+oJ593lo7BBMXhAE
+32KcC0lQZ/SNd46v9o1A6E8gc5n49j3WohnSJlEKrPHqngIka9xJGU+8UwsJim/AyWCzUX/gzK0
o3hvhtfsrgmd8kg8wjHraAZmhP3kFX8ITTJY0DWHrvQ4c73W6Jh/ZsBen1tiZw20wMdXuQtS/oLA
4KqZFZVBqni5KzJTat8hLtV8y5Mx0Nxw9i0M0hrATZyrnV6LgajJc3qhYs6IDYnotNqkY2aVO1KD
LVJpUEw/7PLE/F6Kb7NDqKFS56ZbmN05Z4msye60dePMNHnFZtr2RqIyXz2OmEnHWDabxK4SDRol
N63UjpqsZqG3ZttOlcpn5UDVk/FFYFD6rtQo4yxhOlkXlrEsRsBYBQeunE7QBqOzHSg2SiMnhK+B
wAB6hQLkLaJn6Lf+MXx8EteQM3fRpbN45luKIaN41xBJNXOY42BxwBUsJx+/oFI29U2IGmP6F2kc
4Hz1vJ4wNsllkL5h8MFT60AR1+LMooNMWYU1Boi4wR7NANce6SmnevyJoj7s8kUsvgkSb1/Va+zv
04eLRCZmmr6w+IpAhodCyaG7mFt/baBkNRCTuwHkyRDwKBdAewflUCJUTQt15At2+Ilz1DpyVZDK
cUj0pnYTt/x3NK+TY6pR4V0s54LeNu7B6JVMe0ydu1YkzSwVijuuyGMGfVEE+x0OtayMcSnSL0Mi
BmPYJ7W8q9JOahuXtJMKD0q6etKtnAfuQ8QyI6ZPG+JztbZjyivijlGvpyf9BlMqMvJ5PIWOC0BJ
6fiVbYnH8c5vlSNYTi3sezMb0dgNGxq3SnRPwLCmhFtqySbjRAjTbo/Aela8m03J1cXap5u/+nmZ
7ipH620r7OeNil5WVvZ7EfpkjtqimjekLF8CY4kL+KO3mQBb//8Lx05QNpD1jRaTtnt2eTX2PAck
LGuz1ngNks1T2w8OOk1XVgfNyiiHZjjtaAaMZ+fGoQ31gTWqeAqeNVYZ1pt05ROISOaad5mOpa6a
J7/gI2dV/F8g3SY0wa5mG53Mqbb38XLW74C4C1JvIU2T0H5M6uCk2igejCBM29jr+LCfi+UmOqzd
Pg3q6Zrn/DRnD+6YASTc7r/CJANw/KShZF8VI7Q8K2Mip/qcxcq63RAu/q67Xf85hnMQLkNGDQmA
cRH2ThWJX+dGO9/e/r+kwQT1oxttQ30h/szMmWre9iJr7vgRlWucU2/BVmI+WN8lhQjhZ0MV9CWy
PD4VLJfc6LO5IFGWlLp/6kWIqSgfD0fyvWISjykyIECQ6NkCQ5tOqQYuuStASk1pQHGGsJpliR3c
ukqziTfsZg1Kn1AwMAvYsdVaHjh3Yykpx8gEbWrMtYDppFqHzZpYgWleUeBpgJKN79IyyABdRbnm
oqxtJ18krS2ykWRmsnomr6yV7g0oCUWf4XimahXWSJ1q76yYCC0ItRifM+6FYGdEvVsw41WgnAl8
JNZ5FKgDCZauSP7H7Bc8b0G24g7sTV2UV8OcK9L2ZS4AuZAGbO21PKyLKg4ZBLWkYIZf7ug6fhP4
+qtuk119EKgoPkTVet5anrEXljGJhNnJqj493hNd7y3p2PUH493tTHzPwuD6FFGRtzBgBfgJ/sMb
wGCk5oIbL/wHFNb3HeVAZ2KLoL2LueL67x3hX4H4UGsFP6Pa4nEA1a0ZpBnBeh6z7tmQKLv4PuET
BNgI4MmnmVsi8wXdgnlk4xcfRn1Q49Lh+RGhBSSajPOEoYDiEhzVzx8DlhIA/OWU+8n+M6Mgtnfb
cGDy84UEDtUm+q76kU+Jdz63OY8NhzllptBGwefmnLOMd3UDGs1Rl/Nmcmwvi1DBphX30dBiRTk2
6kqfqxmcIPrr4WifCpfHSf5dd0PwW1/GS76xOd2KifSAD6EBw4ATP7Oavn4Z86mtZbITAB6VBkGS
aSzmD6MRMs2RKqCUmOqbAbPvuSxfvOhrP0wge+Jbk2jOke4JS0UkMBowfDRtZFSHiPbe2eacsZF4
br4OD6rQIHc/IpIjTmPVylz9ohfbFhNafbUfLC/DkZb2Tc+03CzJB9debXWY1oW6CQBoiTrIxzt6
c/PwCkJ2BS9KOOcS07UeyMip9w0QdcDba8K1tQgqE//8Mo6ngiOt0qhbb7GGAWwsEAATR1EODHuw
i/5ri1Flyta7QjYwHJppIW75O8R1aLF/1F7UF8ZNKtSkYuzagXQ+/MT2rjpfKU+fD+IxoT1joLIP
JrsMw4Y+tgh795awvbd+Tj2b1oQGFa0JmcimeeaMgqsFs4T0YVi6xZz6tWcXWIpXJTAi/C2VSBuL
E7Zp6rViTB2D6yT3oJnoNEL5oS0H35KSj4qeBiwMsXwzXViM9T4TlwY7hD8XkEB1qeeK4iE1Bhyj
WPWNIauDXt9fqTDsoP6SJBIocXGI67O8aiFPjpChFdkBDxwEN/z2hBuxKeVXbIym81oKrhT4nHtn
P/B1APQmJWKtAmkukziooXK2GPfg2zCm3GAnsQiZLX+Gcf5lgeBAiYTHEOAls8BXbf1iSbj5x8RO
Pk/eVOTaE9XXA4WwWf+ggrD6ezlUwvKStD2FaJqa4UuMbkPF/gdiajGHocWj30znW/DZzKhdvGWo
RWMdy9YxVbJA+mnDmT6FoKtciOnt2tOEkRg7asHBNLlmemA3GVT4D23Kp9+qI3VScp1beQRBcTdi
/EdY2vY+8WogfDxZCI1CTJ+UuAceAeZssPdNDIDGIInSC3GBVc17X8GrCvhrWTxdmEDmTQFsMeJG
DCtiHl7jGI+X5wnhdvLZvSils2sWAlUQlgIT9IsFM96BosAmTbCIMXKug2IAKmk2xk12dPtuC/8m
L7Pc49qrVzX0ztVjogmF4IFDKjevXZBkRrgxdhCgrLIZnspcWBRokPz8pKerEUxRq3HG9vDsiehI
S1jmtU3j6ZFzuXaLOznTp2IU7ITs5s6+vSca0swA+hvEICKsrVajCTAsh6LEAlYvUKuJoDCl3vmz
5YqR3OwaaG00wQbwMCpTe4WL9YMdcD2zioHU2WxfzL5mIEgPwK3Z2tv0RS8eQ5BxreVifSCxDRlp
hURyp/t0/E6D2WrU2YHg6t5aQj1hVgyjWtGdQc8ZmG06JtNDfM/b5g6F+WVHoHvtbzoZEdwKwfD6
FOW2C2bzl9ucGZf/cyQw7Lk53QG3BTUCGPJjmkr1DsBg+y72oaVbQLVIXG7+g+4L7ibJVBZDEd5D
Tzi0S/6HokUJ19pOq0YxiEiRJNDjbND3mQW8C7rROPI9EKpX3BhjJX+df/oBybWrC/sglzp6pLis
UYOVY+MCjQt1V8eHHY4bpIOUoKaVbIs2fRCwq9TWNWkaGzgtw0nrmUJmiSIcyIyFEFCXGqWTXzbv
s+LqPYus0PS5i2uSwnoK0/dnKPi/Gny2rKy2LAjbR9NgPlW3eXu7FxNGVCHfgnerWqHsZWc9X2lj
oZF/KRQLLDMznaOwhwOqK7umIbsCMm0qXOJyal07L2bBQNat14x9VcGTDQmPk/QhuqqNteY3RTaY
f2dwbTxK1lRxTvrjNoAgkLcmwX0rVJq4Ywcap8LJSYBQAftzzIjhDulZtupLbkrqS0QpeBNlhTg0
pxOvvtIrjoptn9kYFnZS55o8DXZSqm8hRnxGDw1CuUPssDhukZMIg96zcGQ0s/uGsxyPK9eZ+AGi
RSm+GgFWZCtNOhoGaOXcH3JoMrtAcFR192KxS065AW4Lu+MQBuFnBdQBh/GrSZEo/E/TDI5kzKZa
4/66EIbxU+mrgkMGntPdZDAgE8PQBINWnmf++o73w9Nw5ASfhiDX4GRkpv+V1T3m8TS/N2qQeMC7
9EPpbxua2xMX23i/EEtiBiwXSHPlCnCetaiGIpg6Nb4tpqLNQ0uuHSl36qru0C48GKFnrHQEPv2U
cBuZT97uQu/nSEE7x/Wcqh2MxS2D/8UkqcE913YxfdfbUCd8Cf61ZJe3Uo3sWociljrCTTPRixbH
vQMxNq5aaOcchO1N3mCfPpOloS6cjTsqXRzgNV/VAO/6XL+dEXazgzWErqgLiYbVzF2/Pl1kCIWw
Bx3TGgTeGDg7I7LQVZdXf7KJTdh+UQkSk+sRMfQmPolCFVqfU5GY4+8cePkKYbZ+OOEASQPSNhd6
CWwndepZp8GC5mSGSjZlA9oUIT7Nk8BTh1LhazEIVwQTnQJLOncpSSXvS2wMODdURWcExMMDLa7O
dNm5A+0SWA9OWHihQhO2nTIaI569MO47LPFIY6/VDWtZOeASI7G/IU1FcnovTa2oClivLho3UFPh
DWs7uyfPADBBQEbz37Rzz2HghezufW8m0ZqUYUKUEgMU9I2nDnbP2vo3MoZI7Mud1QZNe9JyOy4N
GQ9xypvuUI7akINodQDikpCoLHHzmY7YfQRjq9cGmdBl+EK+RVfenqDSRX63q9eWiCzdakfXtWyX
FHkP+rqEhIuvV28/xuYMhklB6atyhNubWc76uVgFw69s8zX9NDAZYzWh7BA9clggAeYWzI5ve3nT
v8XbVGIxyNDWaF0HC5jYYrqfZtanCo1HEA9uw0vFK0KKPSvr1AboBc4Eh3/K+9vz5KwuW4dyELHW
CTIcOPwOZf92wmKyWgXuewX5+ysUp7th0A/QEABCKTTZYIq70IYppYaCWKDiRQqnaua1/K1Qd0DE
CJ5+PI4B6Kgvf6pkhIVA0x10XkJHmhS06BQtAeIVCXVCQvWmGDNWOSBQ2vVMecHYwl5r+o3SRCRt
J1iUnaAvllV8CveWBafcWyLkbsp7eGQJEFN3z2gYXcmt1hK46dYUPtwqT+UbCFT7bW3DkEQBvbEn
YGFWDqAbdaWFT60G21EAlI02ZYFVabk/26U7zDwkM5E7XBOi/zGEfqk/4vrZuwFZpnQeWrVgX13D
6xj1kIcS0Jt0vYD1N9kmYWvaZWi5OfrqYNYX8lpKoS0N/JzMWFwIGjhg32BuVN075A0+N0CBnZBd
tXhuv/p/34kmkuiAv7M2d0Yr8Zuk76FPwvexSLU0WB3yTGS4uHWyL9gBGKHJR0Eo9w1Dk2AySGbz
CFMNoJOS2Xc8qvivgQ2xG8ZZsLgxnNKhBKpGfKgFe/kkiZW1xztl6jlHNNi5HZ6+pRAMtgMp+bsM
jaHdVRQPxlKk4zgJlQoh0TuYsiUkwkhfybd7WcgIVxzv0rydHdWbnr/YfBkEVOh9ceoBe9rWah29
kFE8GP0duyhmXyEGcAp25yRZ9FFuUo/iuU+foAIDsRELP+Vgh9PG9jJ8jt+w//nKP9uXHVNZJi/m
0It2eTQpU1vIXTqf9Xy7ajcdL437i3m2O2t6pfEwb3HHZFLZFiXPHQ5uiPkEllXGVAcX3FseWIIa
7bW+z5tV1PBenH1T8kX2G6KGrT82m+9Ibkyt3zqmU6SAmxmEbdl2ououuSAbzE/yXTwMXiNZOTjB
vilpqSZ/A7UdaBHrXwYd8wpjtx2SVogothR4Q7A9zG9YpydH9Afr8kXbnZPAnT+EVH7ksY/rmnv1
qsvP84Hmc/rNvT6QhFLYx53xMxdwXiVwmppiFn4FEKYfflL46hzIsoT2GtmeSt2Wvw5cXP2ZnYhn
td0GAH6RUBQdNM1S4wKnR1en0YFz6bKqTtZN1tjr2CDpO1X5IB9pY1RXOwaXwi6ZvHKOojytfxUo
tBe0TUBgPsGGz2ar4GXo4sGqRe8oqdMl/6DoYGInHqW+UxTPJa6lVOaw4kp5O5E9ENIMYR+xMMe6
S+H2otvthp4+8XN47lZnO+7FSwNQ9laIIoo0cmDOXFKt/6Jv4Xi6JPpKcX+gnlC31XqwFIgnpYcA
nmD7AwecbksC4hjH04/2A2Q5QI5fOWwjsQ5pT+e5dkHM07vIBc1eVtdo3S3DwlU2xPxxBNR72QYG
8bmF9Ij2VycJVUjRpjphng/yvVeFA0+909UmAgBIShDRd2zT6+hVrWKVqDKdbmQXEss4s+4doY4B
7v59iz998MNY1kCsWueHeWZYviTItojeZdF/Pb0N48cVPPh3uipNHIrGPuaz2dOTOD0qo5wfzvcA
CvX9MthBwqrFF4r0T/uzTOWKvfPNykqQG+Pk4HljmT6MoRyBTY9Czo/oyMpO9QNqC2cY0pFaPpW5
T++Us/MaB1EfI6rbRaUs3lNKIh5wOm+3S9KYXBq31hOeFvt0XvaKeLixoi7ijDFTv8d3dzfyo+tn
7BTO0/9IhOMm0PMZpFGFkKbaUkaI+Ei4O1xISWWl1v1K56t6GvOwma3HS6Nisi90xw0iRZJkKMdZ
ltfQ+MLQ6sOd3vmCIpWkH4MyvkDnYgU2U6Nbwuz1JaKNRUbc8fmhnANng3Zu6jho1s94PkxHYhSJ
cL12SRZrAxFdltGe6Z0aqrELETsGs64rflt95ZbqPOYFEZxnD0rHq0IaM2vWxYwxx3lsamQY/H+g
LbGlLH2Ii/Bul/KZMcjkR5kc7Ue3JZNuWQQ5JeSjnpYn2L8kr/45LPjzRi57K+UMg/Gp1lTAn45o
FMpc2nGfTinHwnF0bO3UPiYQypd+J2KgoV1uWTp4QcJtgdFRaZ6A2jMgZJtRrCl5Y16S/oX88z+J
lZtCcUo41zg28QM/J+Cts/04+h7m/GQ9TtYcSL4MKDqXwUhruyH+NYHEx3vHJGXOE27wC2PFD6Kr
WuowWlnSuUJ4MoIp175rBWQ/4naeTzaje/eKh2Vhrmh3SJCTSMflX7P3dduz/VO0GTAwfQx7vUBF
FI282oprNQqnj3E/14/uw1O+bb65SOS8OjS424kx1f8TiWE0mBDHWAiCi19+o68aieFYC5dQvWj6
UCZmjaW8/1jJhGwV70iffVovb5mK9O3zJ9aZhMInEiM8TBu8fr8yTNs2iq22BZny0FyZCF8TLbIq
KOt8jRal1TQK11xb9nHATTBsF5I/ZVnMvSl6Y0wmoTXCg47IJtTbQY9qlaY8ZTzTOR37GEzny7eX
/vM0E/xNc8E1T9uQA3tolFo+he1FgJRaL07Irqshn+i/bC9vZYYluK1xoHu73XDnhrUesu3rkrXx
lsFoNllGOCLhZThAULvgc/X/9aBIqRtc/lRuX3RKBgC5AiSb+ukGj4zTESTYjK01MNMZOoD8hlqQ
z8RRg2byr4d0nsJMj74UWTfX6NMmpSP5xbyQ3HmOLsOFQc9AvAiQtUOB/mZ85wm3uveIj+ixerRT
fZ2bloU1sWzuM+5xgHqNGH2G0SNl1U6dbve65Lxc+frNRKrOYaKafzADu6WpNp9tT21O+7mZbSH9
DyR+2U3bAPfVJ9XnB4ZLQNo2uYgrPmodx7pVQAHfGa3y6xzF/u4WhkJJSWdX3e/Wjqyugn5Yxcj6
HxT9aviBbfT5FnF3DkU7EudP+Y4i1ySGyfzqzqaQA0AkqrnnSXswv/3yv0uh8BoprBtRx/46xH9g
Qy70zCMBRuDsDMwJQBp25lKu5O/9oGDc2iS6a/NR0+zCYjHJhHF+0JFJwWrrFC7aOgLsLXqq7nVa
t3fc/xmMaY3fYJV0sxMQXzxzi1Sj9wVG+XgD4BNA+LfM5DE68EafNelT2edaFn4EsfIGuKCtDLa/
cJQY+uClZOj45FjvtmSAWYELVTBEjRVaP/XIlli3TuIyjugedFS+LL+V17PEREvkms1UoQIaUsUF
onUDqMTX8Yl4thiSx3KFB9d2B07lD+faUxoiUaYV1/7hbHV358OukahejWd9unJzFLu1mgcmC1Ia
g/r8xRRXWZpFxLKzrARPzUMo/7Ucb0KUV0rhgznW8rnP8HEF6AJ7aIUxglYrEC+3Kms7WUpI6IqE
8xnBH6JVcBUvxl+tG6ldBBPF+hVvAVejI89lKmRrzkRoJaA6VWe3uHXyrohWsEg7TRMdPTCe1gQm
M+oq2pR7pEbC+hj6qzCaJMIxOrARqZSy5FGZFzV/5mwNbNRibdwYqOzQ4/XcZEvjUxkw36LSgje5
0puxVICOwPYThmEoa6V9bVIch+P7lEG9wB1P5PmDUksznYYFJEliSo8FKR46VKNywW/U78E/d+tg
1m0vYD1rcOtr6ScfrFqSeXf49qzlZtKBQNuSvIvvH2S8GD40vYt6S4CqV/oHhjtlhibbynT8t7Dk
IXi6gFVcs0NJ9ErtPgSYqSSGljHsnr2WdWrn9mTONNEg7qA43avqrV3jLU+cOdSE1rn7Yzv3Ov55
xshd6I/whVXLh/RWNOpL/mmNSp6gEDHq3JdzLSaCuYwpMVrmeDXRil08X9SuMU9iomzuqRlcw+IG
JQ1yz4ei+Kp1GMJt/VWmNyEZ7St3IhwtoBt7PZKwzqNs3k5/ZJYsObPiN8vfvkj3ECOAwrOJFiYj
RZTIEpeyrU/EmnlMUhOVAqwiaCYsIKYfhrVlGXuwE6PyNdyTc+l5+UnUcMpZhLiut8kDjtjsmfyp
mXsuj4SdG6VV1xvT2mEqj4YOmvHbJN1ODoZZDCAr+pbOKpk2jq97eb4MfgVK1ojl8DKVC+eNdv6P
TG6beNOw2vlDEKn0Ene8fn/owLE36vv0+fiiz/ioZ+8b38DeTGyedI3AGFZTXOAiFJrQbh7j+j2H
pOoqv+IzP40XJmbSfie/403q6Ezowq2phv5HRlUbr7JWay4SK8ymwuc777dxsB2pnd5yPf6hUf+g
uc2Puu6DhndZikti2GMPUtk2RLNxeUD2hYhJz0JmkEtP+1yLcuu1sO6B+Pi4V0/JgR84yZVVpHub
i3gaDTxoVFEd4RXi4/lZBebg6IokAemwbT/SH92MN5zcfcia45luXm9T5R3s8AcoozktJm1UyTNU
uE7U0nI2LDs82GGICHb8X/YVaAq1+qysL30NypFPmTs0vGTgmGTpPp2alnC/SOVPOPyC+brrAFDU
ghTjve52B/HPNzmUHeAIhVTwd2lPv+atDDKqPVxcc3E3r0nODI5AlbkkCYFc+uq9B3B3d9zwFZUG
0IG4GALi2LF7pfGpmhSMcgENsQIFrijxbJXjWZMeG6CcyURulZVd6z04r1BwEWKQDi7Nb3GLLAXA
7FuslB+b2cihJ+OaiK1uCjw7H11BF9rOuMeS1uWGCNFe7twymxV8l2fsi0QcXKeKDL6Jc1toACwY
kdQ8fatY2bp/kkEHgyv+F67V8VGiIn7VcMFQW3gq6pGGPibECqHzC8h2mvIVvQJkiGR3Afj2RjBX
Pd9JIgSFWLaDaWYg+EbPmVQiKg+vPPurOHrRLAKPJ2+cNjyxopyWGYvdxYX7vLEHXqQfB+9+1f5d
OeSv5/WL6y8Kj++tqXUaa7jETRf4lIrqsyG2UmToJerK7qfStPYmINWi/YdS1hipykRsgsPnMVcF
vFXkR50imS/CEPg3mXYF2udYYAMhNifE0D6DYvyyOZ4Sxdfrt2fHtVx5x8GFfjxJ+ubPFK3apYsb
JVAhVRUOvL1CUaMaVmGvofQ6SnG8t5532A+TrZD6PvNENl5vASyQ/3jwH9yS5AddBOzF7uebKKGe
YAHGTovjTUEI1dSrrm5uh7bVS5X3RRXf2A2KSViV04IIuM8UY0+8PXrBZVTkaCTDCiAqn734pYQC
8sjwRJiZmik/uDy+5il6WAmZrplo0xC4+pdegrWxCeQ670iZEJs6MzKPzgSjnJ6cLpkjEaQO+MLO
qHWCC1lXWPJtHm6u5WfRDMFDb9j1jMg0JsccbuETyMW1vREYRBf9CxAW9RC4qivOlyK2ATgyf28h
K5kbTb8gI+vUWXBjsUtCMVGmR/iIG9ZTd5HO0K/LYXDT3iSt0qvqVEM8FSop4jxuUYuJHTt6X5hU
JM2C9gI5kknDIg0mh8fpiBIyGQvL40Bf1xYgO3qZKbTm38r/mPSR+VsxuyRPFc/97EcmV4ZfBUyA
ZLSqvHp9YZrHxdm3s+rnonDhn0DqtuiXAOeDF6hPOr1/KXCVBXmGkxi59BcosrW8KvGGtQ5D2iQB
q8C4e9scNenoaNID22KdNh6u+D2KZI9RfLg2Xi7CrOMQa766/pkzNb1fhchhyD5mAV0d6HRT4pcN
aZCxxoEOPNorBuXifO+CmABHUE5Q5A/aJN+NpI7ZQannLUcHgouAP0COM9Q4bwCtqGuKlpgdN1ce
WrgNVwdOrKaGhNteaotd51VKJfoHPaULd0pikwVIuoLhnpeu2zpOebIGBnwSwS90gyrpd+fBpSAj
rYnT0Svo5NDcQ9J3Ffo4PCk5MRaV9+CzokVIoNKQIJGGLPLvTCxR95sWoz64cQnavI95H2RfTzsn
4eVsgb0jrkdKejz27HAQzhHakdnzyalPGzlpCzEiVZ2dQrLuNGiAPMlHCsVV9fuxa5PVYDPkibWf
1ffe5RjxxD6uIs81dXZklQQYPSbwjqz3txzewzWL1mmDYHJpEby1xfAGvxebwYSs9LZm0Hn62vHp
Kg5zUqx8msFcSjjUX4eS3A8W8ruMeel1w1NgHWRDyRwZ5mzWWQJq7DgT9gNvHQ6QtRGXw0aZ9KkB
Za9ljJ6O+JVUFviGBKgmqNjqMeP+zXmfPMMJqaRRKL7r22u17E3KP9nuv9ouzMUuGZLcO/YKlpy8
35dqrWizRxCzCppFHj8lLA4SqL2uK6qkliPnSDAKjLXyaRkFKA1nIdzrVpCtFbYSphq/dqNIAq2g
YVaPZgfbitXQr8143MTQnipmMa8KPBF7FhdATEORb07XIlGy0CiMuBoRZFUZRyB7dAsSek/L97Xy
B3MC5VkMIqsuKyBQkO6L8tUi3nXolSrn1GG/09x0VorMW5Apq8Zkk3MkXA0QmWX6HEdC0pcrFhk/
L1jg3viuWiT4g4hK++FgascswdhjruS6GYcWzcz4M7NFADpmmPqdL3dK55pcDIvWcWIBBm//T2ZD
nr2jN9OvKQQURQlLg5DUQ+4S2V7Xx7SQC/+lPS2B3Nj/1mfpL/AApcdzLVtthrcjHSgmf/iw6d/8
H8QjHPixm5FC0stYXldRczG6Go9RU6zC14KE65hGYYTad8wE5upkFXDPP7pLrHE7mW01SNCB0n9+
x6h4uqG+wEUpxDvgACr0l978745NDvh2zl0zX2nBetrwoC8BR682ub6xR0dCj0F0G++6uWg5gJRJ
+ZRp6zAYX1wjUbdk5DIX8n0DcPJDY5zs3E+pwNttAXvrTc2gcp9Fob42Ymbtdq+fx/ODFx/gpUGW
xgN8HjIyjnsUvj8qo4MvROQU9X+7gYYpifqpvBlfh1axoCXWROm37a+EIXHltSrFicFFCrpQEwXR
gg7iTTeMRtVu/goMz4fJSv/OBrnKoP5A8bkJDWEj9FPqLrkzpz8KpflmKLIb1CDmxxs3/Q/nfYUc
nV1Yl2wRQCS1/64okxHWZvPf4Sbygu8Nn4QaQvHGzkF1+IXXg2YhY1Tp6C4Q7Dt2BTIz3gr2aUaC
y+oAkkLLwIYW3/w5vNND2P35WBSHwJkQ6MW9tFj9zSJF6Sx0kB5ezeq/MVEjJWi3tpLZzqY80Vue
pSVDDZr7A8NwzNRAePcxLJeHUHcETYw6ju9TbHi66ru1MynWCjl9Z/dG7xaLw9YcGB9Or7ekwN74
FQO59naqb0Jnphy6CyW646t9zd337klfWuwGFwda0wvNvRNviyUggr7XERMexPWlPkQ2+8ArfI2m
pz+xCcX5R3gbDGZUfkpIS/ZJ+63BkNMB4EiOQP5ryel/DvZzDdSHsxXNl2UpWwf0F0ODCxhz16Ks
sYHq/pELkez7in+w7sHH36x9wV41Z8fa3t9iMqIp4kgBuz2AQK7wL5XbjvPs8AZD/B8AJlip+uvi
8XCtKXX1W7eD+O0Fql9sAZMYfKAmXooO2OvTOuFTk0Z1gWvpSKJaxgugc27ph6sWtiOOYNWaNnV7
tWTUtTW2z6khNuSufscvTwVdubAVIhqiFXm+sSYDQRF6sbuoW58WjofOYfbPgNHwbhYKm4+jDu4E
s+Tu0Q9NuHhXda8Y5mAMImTTkfmTGT5PbCI5JAK9HV2n3hBc+MI+qc4LfvLfKlnFcO/PmO2Ki9yh
UQMc6FJKopzGrKpOXF09qrvTtgcZbWGO+QOEvQTorT4rFoSVV9rxTF3MdO/LRLyT1/Jh70NBxBsw
tveO2atGeFjkx+pJp0195XFAaiPnf9kA0ATuYcFwlMjN3ckELA1PE/ehDrA4imqOhHODLFZrtzKd
bxCiSS7GJeWV5pOiWpRlK8WeeA4VhhiPVAHj7H6H9rHGTObR1fB8Yqbmhh6zEa4yygXHkCUy0WhO
IGUtHva/GkqnkSl4ATKnU8zudQ6U6p1vOFeKQQKfdV9A11zEoQtMKb5n8qoEQGx2u15tYXuJjDPY
O9h3Adt0AkcdkSiXWznFpEZnTZfwn8XU0I2162s8jNBdrb8aYuKggMSsoEdv7hs0IxNBWys1B1Ik
DntQ4KlPVE1XU2g1MB7f2WhK8BTiHQS/ubZl8gBT82mRs6ko1EDJqoV2Dg9ngW3/KDLkp9EvRPzj
h3MEc6CxPpKn8FlJE7PipKnPcWVTBceFVAHHBkKPBnvgIXHpxY5Ui8gNz6GmC8UVQJubQe5+8kls
XJl9aMkT2iiRBiQ2rLkCH4wJn6NR92jJ6NEYN1Y5PwPGVhwsgWbk4sGrPtfjJ6eyj2nCFmAhDYe7
B+yDpMx2j78SyHIbz9Cxdu9Mi6rSRil3j7nemnXx6GtX2uyggfmX94Vgx0Vezjcv+/yCJl5NlJr8
Gmnj3cVWVhPy1JOZSBi9aULBthNBpSfbZm6E0PwsspQ/3MAWEWx8S8TUfVz2r8tCOAhxPCWR6524
xZP4p0atsOa5A4DjPlKVg0EA1QLijbOBlulTSJ8EzxJMvWRZhSvgpzwh54qvDo0Qcd9+jd7RJK5L
G8TThUBAqIaxX9PjTSIGN+iHD3MDqY5yAyysb7Zlgc5/bJfG5YpRWzMZE6pfanUmlePkBsEQVEip
2P64VVFVT9RQen9tU6uQTAk5ey4DcoTwwuj4U6PQI6LAk38t58jtoXEZd9Mm7OFXfI4wna2sbt+E
7EKEJsnrB1whyVcnnoqS3X8Jh48GPDGNsZxFWU03s0vuGXVzU5XwuNoqvkPGLQV3m/WqfcLTE82K
pq4+8HjrncPDH8NlU2jKUWCE5Yb4srTtSG8XEH8hSwPqENJDUTqbKAv93rGenZ4iQicD7Lh2sBCN
0mtGMMyAG8+H2Fw9xiq1aCxmKZH2DvhARjMZ72YB0EU/jT/BRGgwT855z2OluhyaDEwrCaIglVXn
w7aRXttW8iYv9N6qw1KaKNiL90ZSUyxiHqPGwCliKCz8RHXzrGGYzr+Q+OmDUYlQ9ESKeXhM6cxh
E/5s/xAQJbCviRM7vlOXXP+im5j5CU1yK8Y/4MNx01EFJeJDXAWMMGHPmSu/rIPBoyaxHfg2GbwL
+qyUY3K1WaZm1BFF7RoYZG/FqhrnDrv4R9aw/AwqOSfidNtlgH5CprgBXIRRDD2d/NXMzk6mELP9
vkRjnApaoTei1Ec7I1NDFc59SvfYeq7qfXDLYLGkrjhTlONdOgLU9ltmBZdtnJEibhrhgS8FrjK6
DDAZa0pF/6aDPQ1jxzD9wTjxoOfh/kmWngYj1xkVEvNQ4DroQZlC82BsCHw7Q2ebaQ7MDImYO89x
MrCcEhvYDQwNgi2BF8Ysc4J6x8bH7VMTN/zJeZbfOdWl6D75v494OShJNKV4j9pB+j9r/qr/hTXi
AR94fkEksqN20DHSwjthyn8jbN1USuKm50D18fGsFEly75LMspXt6902LaFubsSpH4WU/UV3eRcG
uHp9ZuMLCZUWlR0c9l3bnXVWW+ZcIYoOeDB6BKNrf2qR7XBADl0Px87OCH+anVl2gAKp4ykqttxl
BjWqnkJEFwamtNPNb9GCimUwuyq3L0ZML03yaFG+zA5lGOZDOsMKd3UcpEtQsdUWxmX6v5i1cHJz
F3G4M1IGSxIR8WUVSVSNFOr830ucjMXvoL9teLYKGvAm3pjoTVUSt8pS0o2Js53q7vibVFv8bcS+
r1C1namdoZP7O5eSMGftduAkqMpNuK3qaPE7FF41qaH5gWOE+ZdhgWy208RIy5dfIk2Xc4nvrcS9
krXh9H8N0Js/wjiixGDnQx0kgP8hxieAEBFZqHADIxzl7US4IBjPBSooRsGrg53KHofDPdorl43m
EVHI+/wJIBdWsIixls0OnKnDPTzSQda8rj/2vdNsNpLHaCYOuU7qpfLZbXnVmp3DuHy7v2gWKRDp
q9opGTfFgzT4yBhUCywLH7yxuxImGbJoz85JucBpWzJgdeh8jwcubHUGLHqMtJ1p0Z4uyPOcfUq5
KgylOWhnnNU1XdVijSGKh78JpC/gFZZqeDXiwE/40LKpGdrEQ+sVVihfODwBi7XoXHyFpDNxTtWm
4GcvrRmdQqPbPauqkoyfaHeEe6BSnna4H1hFH9G6lKp7Ui9r6gInK7iJmTl9qfxqLVAmpI0BlYbp
3Qz5lmKWk+FfHI2oJDbeclYDMF6VocyiG06ZLVw8il5WSREnqdSKmfTFjqXuXYej6d3nnaSyGZXc
LlARpssFpqPhOUf+RcFB/nmItPSIGhr24KGt5mKd+97QevLoLN3RwNCuixBMojRrcf+gzgJ/Qnno
3lD5gootgk2RSpESEUPricY4b9JDH+pvtjd4BmMgZPtH0R9PfPZouiJl+LDb/3Dd9a0qDoMsKlfr
/JMCuRaoSAfaJtOOPg+xIe4VVXY4FMs4isugv52fLG5EWMDXN+Ss56BnVL9cMs7Ws7URnyAfFhcU
IYQbvAc67h4qwmA26bIWV+lY7UTE1rI8AGaB9yCBL9GZ1Mrc0Djx34azt+77eKlmXGqNBnIfD6Zm
LW5ZFps896zYZPklxRvHrITnpiFuKdd6z5ly6cMsOeFXVrDdme025we/ujwW3Q==
`pragma protect end_protected
