// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:27 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
AsxX1qJ2RCO5MxY7fYtkZQ0VCz0+8M+Z4EGrIrJCR1nLWQra5sFIF9VXUuhjOJEz
+LGlVUjMK8rKZJ6/Trl5/u5vrWucB/HdGOBf/ypEexnaVeDvnpacbNAQN+cId8Ul
8EddkF4oFQWmFeK6Sma2e9P0dOHRC8TgmE6Yygbp6Pk=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 9328)
GGjOC0NSk2gAAzGGGLMiXNLGq0rX8P+HukUxe6OEAj6Kv04fbddOeZDECIn1NhwV
K2i/aklD9sGSsGb2rCI5bNcxgsJmoWtwJAmDsd7ZpnhClaTirplzk/oGvcJHbACI
Ve3nUx6Q6WJzU2VJgYm958TNBf2MgpnU2eEz70ILXkJxlWUjCvhqse2dlKNZi4Mo
XQnRkWj1c0BIC4ZP1MDGqNwBk9tEi1QbfoLe7J7AaVA1c4psfnnpxO8HyIrXULhI
oqVkUYsnZ5lx3C7PYYncXWKKhbKBKY0izPNqxyp0FD93f8d7Olg364bsoZYAr+EC
npc3qAAgzNuyfJoIWtbq1LqmEDgkLqA/e1d6uYeYr2SwL+/aARQIw1P6I0/89iDo
wJRaNSdkDhVL+oud19eljC4TM7+v0rbDtGkvwWkC6ezWtcBL8sw1ZryHhVAsvJlJ
/7NpjwJpQxzrWolr2D42FgCnaJK8N8QoBof0FmgxdNHYJnNOhzMAcBLJjPo++dhI
Er4gUMka2tPblehLd+EaVO5EfVZon3kcOWJ+KNWW84WQSrmdZanCcp8SX2ZbxlJH
7iHOm7T9bUPsvE8hUDiQI/czkvWJSkVnPkwLbJ31bg5e6b4xld6SjCyZkOxd/Z6z
oVIxIAzQqTsCzYkNEBGrvld1hbB2Pa5RYGs8Pa6isMGN4bmocEhPeui+tg6zNg0y
4dWjLsld/cTHwUsaUbLWcxJUi9OvOS3Owe3+hqiLXjfl7YrRJvDPKCqoU37FdiA0
2RLGtqENQUhuEM43pyWvCYdtcF+uNyKZ1KZWfqwNusEALd7pt7/DnLXlTkQQhDOO
8SVpmqW/mGcc2AmWJQnc5mAFCzphmLFJvrLukuaQ++Xprvj3bwBVtLFSErTJASLa
zaqA7gp2IgdZQWK7O2R9F1MD09z27JSqhLfnI2Ax2BOnGnWQ/7vntp1QYnoSFtXn
Ly7p1u35uumuajJb63hoJM8c1otluDq8VtSkzTauYE5OYk0h5jUb2dvm/9vwOWM1
azBR1GizjuJJR07L8br3EC6oY23s0SuvrDcg3d4d6lQcZNB2jU/FBObtFQ/4Jjqv
hXd/NKaam1b4mfxIwbe9rsJjsvizeNxOwJi2IpfroTwM6n1QzV2SpKxsSXp8THCA
JM0eF5nSoyosM+Sw7lUw3+VfapgUGKKm714oqF+whXxX7gQD6fOOu64Fd5qtWN/S
uGqGmkaB294hYyHLykWDXF0G2d/gU5gziX4289tn6RIDGB82qhnlRP7DE65K7ybh
TBBMxKMUP4TnmXqwdAVBerR4Nf95nxa6hFTt5T7mw3wZt+fwus6BhDFLFT0O9o01
o15s+sbVQWwuRsTBXUC3rm+Hl+BTLaDw0HO9rMbfIby3DiMAcuru5wQfZgDMeMQy
ABVV/zTal1yfp5yllvz6Ug+Pz0F3Pq6fScSgmYedUsTL7tiE1Zymjjp6ppW/oj56
isLW1ZGvORRVzuHLvwO/rebyjbzwhnUIVhvXbzzQDF1DIdjlAOQp5TamRRsSmBI7
Qdp0EpREu/SZQS8zNhEY7dcpKy6L19jT64Zx44We4rATxiZ5dLySwVoLrvueXfHq
k7ztO4dk6CsZmM0UaST5jmwyMLo3NzuAVZS+DVKFX12CY4+FwU00OZBFW2Fwo/67
R77d0UCV8Eq+klo8WpuiCU9ezz69UpZWg+z/dfDOjK3eM8tYU+kQ4CygS9dvbiyu
bsM2Nqe3m7052lYt60H8wgKfeK48UWAi+1AJPt8wHqkrzEn68zg+MFIbDxHO/BQE
Mn091ZSzSSVKniDQ6BipVcVKbqXysb7ezRmBsLdaMyRtH9dIdyZIbajQ3UNQBbMZ
TD/037bWUN0y3cypXLUBBFDrTQq7oSpm2JJj7eATj6drE6JY66TsfzMRT5Hps0na
qRyGlY91ZxK2c76Yx84EWQI874SElSaa4M5qn02h3tJocJSdgw0lB1/SiMBL+8dd
0yXMamYI5HNZUxy1lmNURs2Xhea/kcJGeeYBTl6TT2cLTcVLCCFKpN3F6FOdU2Vh
pEfkLXvca7sL6oON/847A5rF3+Wc/FN98Yd6ent89vgMhOdui1xLIwRWGyq2E6No
bmxmPTNi/LEk2t0TFxyUxoOj1cAeeVBnEI5eGoyGRNa4VgnO13jeyauFlBhZFQon
jYb+/xlpvZZwZR2LL1t2MfjAlmgZIVpHwCqDZs+34D7lbEMgg7JnXpG2nKzMRAhr
PW5WrCn/bE4dxS3FJ5g+YYyglld17bXJVNbSHSD+3uZ7QbbrjOvjwBU3VGEB41JI
puISmWuldTBTLqoM6+zBt/vSEI5/x5ZWwx9oqXFPTJ2OQRXv+TAPi7/IcGQDlZTB
TR5DOm0Bu8mFTbCtXjCylE5JQToW59BaJyNId074bLa3svHueZoxUJmZXraub82f
AnSNz5AfHeU/8seVXxM8Hqct7t0uDx+VLWl/k+yb1X+AFWUnP7vAeQl2C6ou/tBv
NtCmjrlul25xY3YmJ0biwC2Q3uP6E7v8ZIYipUdvkYKFYnaXtcgzv1XUd40Ztpxa
ctZjPTQO5l6rUhQLTDzLkRqMfq4tbruXdU3+pHsY4Vq+TmEj+/1XkB8V06oRRMjB
HigX8Hh+BU+Z5e2jwLuP9zugfQquwyr7WDRrsxl/vSY1boPHShs9ZjCW2F1qutuk
W8d9n19KIvzKFbqIIDVNL28+XfNnDZKdVryoO1/jOra96eVH6tI/HO2Q+hoNXttk
o5+vLj6eyNessXrx2hY93J6D1f0yyzB2RcmUzrQbVoSmICMJtyRR40spKctywuNu
LjnCz7G2Z6wzBdHfvhQ4qm05kqrEC3GNbMf+9MRufBVqlmwH+F+PpOtv6XFqIeV4
Ny6j4q0Ms6lo52qw+W8e4OlNwYKmj40IVNmlM12+DvFBbD12lLdK3e9lKSeW0xOt
mcS+mhaRxmf8m/Z48pB0L648O+4edyFuqI2nrNdZyIPD+WJMBdS0677b26Hf+6U1
yCtWf90GEj+sFuBNtZ41XkF4xkf22O/FRiaEqx3iidF2v3MaG5ILgF6yf0BsRdtu
otzTQ8gjkogrxG9iPWmsW4JrmD/civdmNtyaaCfSXkKhlSNGpTtZRkSVVt9F2dEr
WqNKk+8fIxXL9csYF89wIZzs10KyKhBcxJptAQcqEJBuxR6KgD3X3CaOrspB25f9
xXCBb6uM6Api0XU0mHvvOH3fvqtJ3m1nfhz9fWOfWt+NaLCJoN0BMffcJj6Dcx3T
0/YWOIkay3jAPxA9/3F8IK46JYy5JyuSY8DSC3Ajn90QdbRfPif2h27ot6zQLOzg
XMm7wjrkbkgKH0xSfAhZNBOE1Sv56XyDyj9dWeQA0g1EobsvP5DGvwCxmzssTnGF
D+He6ra1+5f8cQQdaI4AmpVQm2oKG4BIc2Ah4hXe8wP1yY4Q1lPe+L8NTlyJOJpX
NyQNbeR+gYKN9pJ/fs9MxWuELNk6Vuen5lM/asXrXKwV2N+E/FX9ZbijJXeCU/m9
x8Jyh2fS3N2nM6dFBlUutkHMhqMGVFFDCygwg2YVJJOPK/pks0V8D39RZ2+DrKti
YaaXEKOoC27H7GmWhXR+hNURxqEJRRMammSNRlBjFUbPxpDQMcC5OirACulAqUal
ikvoT4ZiGaaXh1laOt5g6RtcKMFP7cL/GOX3LSTo+hcGwc9HKNKD/ztaAog19GwH
boYp8a0vbzOb286WvCiFt/Yc8adCAv3Uv178vWnhXpkNdrDXzYU8I20vl7C2E9I1
ZJ1cenLyLzpPFLN8g4Ejhr+dV7xUWe168U2ah6Wi3yWijv6PnSdg056RGrWlY7I7
nKDXywDkzII+TgtXjbuvTqV7WhQG9TT4Wxb4V3lSWF96wCXbejW3zg1Z/0bDzKy+
g0C52ALe87h6Fo7pzflGWXq8KECSBEaJdCwL8I8i6ogdzxIF1MfTol/ZyjPNycIq
e1imVyake64Zn//Zt4WxKfQcN/MwqQNxPkrCbpBABvtEE8FL3A4RyfMthIq35Xzo
60pr1gY762HR5Qh6fB8F6DmKLjikzHTixAmEj86TDcLovLn0e61yts12+OlyWXqE
rUdjJkjknworGhNKXYlXactmQjJiHprogoFkOaf1e0m/1N0mjvCpjsfRgu5P5MA4
obi9UG2w+HGiCbVqNQXBnXLC0G82+ydn3MURxeleKA38QYJw0ODaHNF4tBadx6fh
z8Sayy5b+u46oHDzCTpDuVjRSh0PbdvftGQnMSDSpAN4Wrr4BynAoD9iwHDltR2z
D3V1kkyq+OK//79Pmv7cUkeVjcmqZykzp9xS2bX7mSYp05gatnKad4w1Wqy2dkXM
WcXYxa0RnBJy+vYogp3AMcs/vIMduDcDmzYE3vXa1Qq+mJrJSMgUqqRnN4m3GDpd
aR7OXONhaaYUcfnFUrOkEERuLHM7sBZ0IuDD/LQkD01YAFFhrIMycY8ItxfDJbVR
jTeaViccaGI64hZHnuHk2P9y6FWpopGRunaHixomZnNfi0uJwVyUi/UG2M0eGFAs
9J3fgOcELaA3toGXq68smDhzGATTzNPx0G4/yUwFzuVc8Y3kEkuMhHVGSEuunJLT
Y/nZwN1UgpUtIoMebdPmG/7tX26vmWBkJ1L047JqQYuucsYcmnrscQLDTfyLsssD
G8sDsOIKH+Mh++TYTJxM03PMENu74heyYfOoZ6UMfrVtDoBMK4LVuKE+yCCAomWE
CoPLcl+WfKtsRsQW2c9OiO9cj+R8SF50wz580JuQdN6jFytNXP9GZWZWuqWD6dIC
CklXF+sdg0uG+Yk/hEoVgiNnUZwtJ13ZKWKIUgGG61kKgwszgThZSKTe0rUlwMHS
xVLz4PJO6F679XfdZc0e0p154irbHho6fw+/gIGaRtRaV3hRzPovKRAtSuymRv7O
Tva5g6CoItJzQQCVopStudFnUlDum2f9mGrwVJ7mAc1Jwtd0A+H3d2Crn0vmA9ZV
ED4yByB6t7/eWKseoyfW7czzjgmA1f9mtUWCc8qrHGJz1Rz5wS0KvQz10sj+wY3W
vf/YFPusZFl5e5efYPe48ztjoRhKCquyKXPQ2aEDKxlwaz+tYJVKwluIrYKkg9ax
dqI4uQTSqI2abJRT27MUo0lR7emh53r0l8lbalofKwCdhbRGr9P0gLBvB6/MIwdp
6Kmn1Pp2yoG4Td0Tq9NfAhjzuT8HhoNktvWphCKG2Z1loxeV9fC/2YgmhXaZK/hK
+LxKB4An051hl1bDN4BGUSPWE7V+D23eDJaI9VrGSt2eM0T99dnRy5LexN88tCxa
YPuB82kgyxOOrw44URIwAIUnT9nZzL/hn9g4ef9sh5bzYlRqsa4zsSkvgIwEsKjQ
fnstYfDX0FqPqPUgTicQRKXyzkPnxND7mXObOProgJlBnu8YaBDoDvXzY9j+i9wi
Nbt9ttVs6rHcBk+NSyPnocGX7pPDtQyqkIywtwkhejsOWzgTUPGuoSsMlDNO8JSd
BoKjmjwKcV/uIUYq1xecW3fjEJiDWtfn3fRWYEIXd2f/FTnEgmpJx80mVjNtH5Mp
41Iy78qFpNqttr6s6afec9wZ6wNHQRzk16KBg96dqQnoN+3E6gFeMQqikgaFNTd2
5PwzRLrEuAQUQeQCiPwb1jBOEsf9zIdpUMU7GDnpZfD3BGhmB5MLvnrVoBKrLKDQ
p+9lPEnMTpUpVJUwLpGWAdGR8DygBdYledfPeCl+Y2wG0G7iTk5f5PVws315ZNQo
E1V6n8vyYfkNImLUiW4gOK1d3dI842lphh74rQjWXNRWRA2gicd+KTgq4vlJAcEg
xwtkUC/jo1I+FiaHKTD93dpjQVwPtJOI6jTEP0wQUISNslrcXUZtl0e6sNIM/++t
IyWW4kylokV6H/gd4D0nGfu1sq4rkiA4tIc6lToTm+y9lo1bjfSkB4WoAGUFM1wZ
WjHwGk4xlhlzEK8nl+xMnwEJaVyqVMJJAtmDyAnvWK3ii3Okof3UC7OVBa69LLa5
n467S2YchgzqiJXxw+C+fDZG4BB/iubNq9KSqd9XcNSsVYx4fbBEGL8b9VSOHoIk
Uji4sBTCEcty6/99dpBvFUMocj2Uuo0U8XP+9cd1mj0qIouvLWa4lZbXl1GIRcpp
Q5QPnKyV/Pp7HIBL0jS0bpSdipCdREJYcm2GsoCst72DRBqJmpA+PL61lvUpV/aU
cV8AbI95iHzc39wU+aRMznBYoCiPsAKXGL9haSIehpuNZST1JLNBoGjZd3M7xxHN
gLQMoyTlSksPWV908sGc8FIOdtP+99sUHyCR9mZuFG0xlMXeA5vEYLrt+DS8D7aY
E4msvY+DIZVGzPun6uN3Gj9/Mz3X8yiSizLVx53hllNn3mfOyPL6r6+pYn+VQnEv
a/JDXZHvAKGFyIsqT6h83YRb9PJdX7k66vhsThNbJabfLgrCqAdQ2f6aKpNTOf2c
VZHl6HOLmc9n6g3k2fAgN8Iumym/8seHTroA4D4eM7cLISZxOUGjMPB+VqBHrFDE
FPXEF68j/ZHhdFiSF/XbD9fRQxxk7qhsgqZiff2S7gBcVyefUlNataJh8is0ZCEm
CobvcHvfaK4deCmpSwjyf3W8/atgK4QHUSelLjf9GKXmvAesmb6blcbvndzlFwJD
cFsXUAr8tCdfsq0jLZYubsFuTPXs3JkDKxda4+/v6hzaCXsx72Vu9uZeLzL9+Yqb
gSB3GG3ix/ooPOrGMreN7X/+FDTBkjiktE4BsFEtUD36RY/yfNHSm00CJ3fgBYg5
Se1LMN5nmqSBVkVi6VKIMCHXa+n9pnxjNMLPIG+kkgPhGmQZxG3E6yKFo1TRw+ts
iaRCWXeI4yoO4qngcz+kRK3n9AfimPh96E/qBvuBfZ4WQEIZIz2CotcWgesnkMGv
x6ts8VqAEz7+42ewkBvJmczC2t+u6VfDmu+kCoXU3xuXExLLXRIWmeuBquzTyaWv
cG42Y/j4MBjBuSn9CuaWftfUPlx95uTYpL0jewGK21kpfOeILykrpP+SJk0gGHZo
F/G64tElagrhqpfp+AWYdHNgrtb66pRniuJjsAofAfXIINH127UqiR7UK6JRMHlM
cP35if6U66WBAiDfQWIsMS/YKx2yVNhmcb/7EftbH7eeO879RqE7yIGYRK0uj3pI
GQ+963ghmw03kEshxFr5rxuON2RpI2H6uFFcGuHihIg6dlmbQu/myjKgCQcyXEPy
dVGy3FYR6Vk8GWldWiiJD9IoJE/c/tSW9YKvX4oEaPYbK4+O3CdpQ10hWD3fy9sZ
pjVrFrweYDyWxssCNsJh8tw2YM4U8hSGK/eIAN/lnROoo6Yai13mhCM11QeN2Hfe
gwxkfzmaHZgPsPv8ergWT0VbECCXBXQspD9+1XS1y6ewnYvOQP12WJFP8ylj3bxg
xwO012K3w25QjhmVF9PBtqsEK+vIMEzEJr1UGTzkljU1xT/0KhbxWttbmNemQlbl
Cj/FIDDtvqeDqionvYHgoz2QmHoEE9p6s4mY028o6Cz5UqyXrAiUuYUYr6rBi1rR
+B2XUsIr73vXL4ukAcU/5SbyXeX3mpSFbHxtDQ0l38yQO4eAWMvBz1QJDmNk7Obq
LhLilK/ZQSOBgxh+x56Mnb8QgRBQJq3HApp92BnSgeVbrUB3VdFtJ1A76DZW+K/T
EtfIWQdSBjFIiUO7HwD69dJvdjvw/UDLFsZ2jyzM4Ksa1UX6njO+y9b7MO3MmqAc
yT0R/gpUzWtYXUIsD0bX1czR/nKmhutX529yYq3NJ4atfWP958E/eNvQbnVF80Uw
yyYOO//TGqEDly/JVTDh7k0k4QfDv6O8TWckSq+EJF8b0Jp3N+Llb4AIgDV1jANl
mgHfDtvpd4YGLV3QXnX4eTnqe/hmX66AnY7YGQHqRCwMtKFxHNATEhlzBR+uE4hu
TV3H95ErsyxWRHAYnWor4RJ6TdcD+bsrzMzF6B8Qwswfhx27Qvhlcvd5jzyD1ek8
L7IN1SHHyLWWGttie4t+J8KalhfgK1NpNvhyfeejpD2Iu7i4l5Gbw0mITTfUD80C
e5ZGfTM4PAqoJYQaRo14HT4LEoeKwzjUj/SaUwcejSJZVeBSQPOhBWoGa8x7ZkqA
hKl+YrOM9BiYqt1GovUFqxJeXPCivc9vUt6t3TS60WE/sqvBecHr4HIm2BJfKxYK
fa+duE7fZgZS3QEDZ07RQ4bwnohyWY8aDYG49vsUlfiaxHoc9WaouoOQGOqGrq4M
VbekhSNE0QBw8zVY52Z3i28yKmWEmG5RZGyiW2FeSCQljlfIoZysqb0iUK5pC/XB
OjswSfOx3qWM8Uk28RAGgpcAPrZSknoUdhLoGg54GaWt+cwBG4XYlTWJ4XMfshq7
Gy6J0EfOtMebzk1rPIr0LeN+7T67+6DQSwMYgjqEBDO3FL0ZZensBLBzuB6LG4xj
J1GhI/azYqDlvXsGQqXQMj4gHpPrwj/eKdbcRTuBBOuMP/r8wxkNbxfHek9FAsdF
ZukhfKyUcIC7ZN4vqVnlxxUuCbkf0ENf5NkrHA4OyCHH3yTPilIrSh+jGdVlhCv+
nbZMDU29g7lzBYU0bZf2IJXLykp05xN6bdWQpAh7A7wV+2kzalDgupUw0lxXgkKb
eGTQejWKHGZHBZT7CeOKBYhAs+N15KWcEZb/4/HY5L5GerttzQVAt14gMscjp0bl
HJy0zXe6mm8Wp17llIhVKBbNNiUpqlw+GFucd1D13ztytsjkWuiJs490zGLIrlFy
q4BKNusUbJ7tQkze2PaaEVX//VMPWjpP54EgOrzOhh/77xo3lvMeBF69Ht9QFsdg
en6/RtUuaoD7oAyNv2UgtdlJmAMoa6S6uDTm9Mpkf/Oimvszg+iPkhTkYlXAV2D5
WgHiWh1kDF0EJda+E5djGvWKeh2Klclo7XMs0pGBvCTdqqVkw/kxaASGDCYvk0Qc
GqN+l2O8NAHTQrLjJkSxWNFr6306vW7pDbhwiZyoVcGk3qv4W17fxUo5mlig2+mQ
QiYku66wRScKsIp+5+Zyf7GCZzrviQ+IRginJBtf/lSUmufNtH5tFE92fY8K/WhR
ahqLkqAKGMFIHQpcZECm0PikSwW3f5qEQ6Td9XPGUEonIpNa3gONM29Cu+i0Zq0A
Nkex7XOxLyNY4kr8N2nizX/orSvBI+eddT/+SI1dOL2mUArKmPF40mX736lHpU2J
NyZPE/yPg1xINndbXgpaRn1uTuffASGyvVmj8AZ+dXDywNc9sji1CXwOGW2s7z+u
U7oXqi8OrfQFFHri0DE6K1zxOjX7JMTRuL70J22bGdVqyw947Euvv280hwmwjqEP
ximrRyTaqctKi681xG2Lasw2mYf6SseQ2VPm9xyLkitzXfeEIfBYzI1AUBSqIQpq
qESgva5zWRP08dxYsJ6zBDk5Xh8hEAd63pjAS/E7RWyf+AoTDSa9DhqcKwKr93YH
5QXyZg1cL3dUxNl1m0zdphLg7KsUdxsBb21SPf/WL70q7oPkaCdEziOqVvw/gxz3
vg6CCR7uOr4NhQ54UVvZd0GK0zVaStZBs+IDZqjahxmazFdCO6NBMZIbFy1sucHn
cJ2crcvdARbVV5oSDfcD7lvzLqz9VAf+qpiNyHdL57XzKoBUYw2Md3mZ9qKV5SmZ
VFWKwxeoIIQHd8G978Ir3lpH6Ag4dIoPerD2nvygK21XqqooDG6Zx3QfdMolyYFd
FAa2wi+3vrSx3sPMp174i0THQsUdVu3IE8ZSlrdFRSbc9si7Dev+m1y/3MofiSfb
Zi+xDWmmxaPjPdloLA/A8G2aITlZ8d1r2Ba7cqeCr5mx/vvHVXY9SJ5SKqpHch7j
RvilOSGbC1dDjGleHfE45vvXg6cGGkfPfCQNjaqy8ig3cNmrlFCdN0Q4fMNIURi7
y+2OkHWLEqrAfZ5y9sEBr88FpJlqtKszwxilHJOmxHmfnDK3WfKhhFOgro1SXEIr
g4K8RgwZ9E4Vk8M8vit6L3Bm5EHofuNcSrKkaC42/oyiloVXhiZdAM+O6PhVtEjj
5IFcnWkwXKj/tQujzUfGIYzTQt/OHMwYvAwbheiom3N59dMemiHEfOTWxzNlbUL6
nfkVgXvKX3QrN7lmOe8DvuJl5pEZSzWrlFUECQnP9Ibv+nhRT7akmzg1HZ1ibYH8
AcyUSMbLO7HvItY7nCt+nnWFjxarpKJxwZ5MoOTy5bKxm1EF5k/ocU0+Lglw2iDP
o3MrS+2QgewTO+hfxDfUpSNZDOe6uYuthVomyO8pxcvuXkVlYp3hsSjdQSfYjfNF
WxOupLJB+lgTARBkTixkl89RRFJYIN6mOvkWNua3IREblmsumerMWUuioM2qMZY/
59/vJd+WIiSGTmMAOaY04PdnAODMhZddBUX42IovU/o9hWTsxEKDo+cHnn3gCc/j
aNqOgwwh9xtrXn2JsOPHAgdM9Vxiwz6cx3oe63SlwqaYVBfCBWSekZoUtxUT7qWl
P3eGQ+ejKt97iprOcPGQGvBad9U0r274Z50gvre93uWlSlqUpYApwbDwquEmDHRL
BVgpD3FN5BNH4aCpfooC38Ba9axqLu+sUxlfE82NEhpX7Ojq+Np1D11iQk+n/Yl5
YCIW3uzO//Tn9bSTjCPEXGwW+bvh/C+jPT+pEH3Ok8mM46op9BAEc+z9C8st+CSD
8cN9bNQYpPkAh8dRiS9/PAmLDKsoJn7ct0vNk0J7BGrjj2V5qGCejN+0VzL+F8/e
QRB0DAS0FT0RdJT3d1h5Lvt9MrzyDE/UT/Pm17+p10730Q9lc26xbdaA1rad47u6
sUF/GktU6CMQF/0HZr9XCBFJSra0Nstkxw0j7MzReFChNqYM5MLjGXRVSy7hsHtW
sy5B+ujEyRiRDu0Bayp1G6KPMTqGYr5zBexLD831OtlUJ2EVm/Ck6OvCtWkIkwct
z5CFSl4AEXhz4rsGKMZAW2JHFRjacWyOzJE/sAfUNBEG1lfVmaYaQr4oseZsleF6
pZPOTyJvihPanip4yelaJMeY7MgKPcSNx8Aa6Fsi839rxBe//pT450hGPcyxpyip
fA4tVDYkIO1M86jw6NVjzubdTImgole9xC6lSx0iXzK4BLcA3UAq5TpBTOzOd7iJ
4N31U7op2Rvbz97SlfJvMIh55jw8zUFzj/WhIwNhtPF5FD2Qr7c0Si2644isPUIR
zGVnnzvIgUxVFS02bFvZnlvR3fvqg59smEcv0v5fibVcgjL1WUom0q+7VnJmnmDT
AHS0ETURBP6xeBMUxTVhVIF5k9lgAgRY1zCvQ1gUwkOm366QuvB4hFSKyldUiwIU
QQX3gC0j1GvWYSoB/OXSFnOrdNvYYeqGhUq2uduaeN3/lju/jG4jL5iHVC24ucBz
s9wJdiTSBC7lKn7/EBx3pks+Gv0BMlPgTU/+xNqlRYtR2At/iwEhfXG9BqnrtYeM
G76o5S3W4etJ+N1bc8Slk8XOvs9AQBH5EwfaHhwMmylONqD6qiWuN7Lnc4e2yVYz
HZGZcQtoI55Qe7pQoh1CXmj3OAeky7vzW+NtySw2xDYyrQiPK/MhBHjwuOs466qx
EF0DCCh0JSQ9PYKVM7H+tuhWLevoYmPQUokFXk76MfRleJJrVL32ZAo5UXDaX1LH
TJPUznAGAlLfUHoHPNV69avWgMzt+J8vmxNTZW2NRILz3+oYUU0hp0YMV1xAjOOH
IfOEqcdKer4DwF4LKbjugnJDyBMmcXPmdPKGNwD7pleOdfWOHWZH3EhblwXEymTd
bZyYv1n4/8zR86oeX6jYjtuZMceQDQOTyM9XNd6kIQzs5pdeZ38Aaq+adOPpbRmJ
qKze1vkPzJwgk3LyaW2V/09Ipz4Gk6p8l69QkWldz4IncPlBndXAKM0A2D5wGDN/
aVZT1V2Tq9wqsqGdk/4qTKa2e09yhZhwzAkoDojojDUphn3Y8nA6kQH3BQmHto3Y
sY1p1Z8G83LGKF2MOEe/LUFrdmeQB8+6yp4lmhstqMp3RD4ITOVyZUOKjQnqWy08
/MsyBC6/GfVIC3w1CWSHwm1z4i19ni1w5rcrcSYfn6JScvvEt0VgKLJLjpbX9BSa
92RyotDhVTI62KNc4+iKK5/lbVrPbFjLWqCZbw+Ik/zwZypJeZK1sUb9EHDYipCB
2wbEr07LtUnCXJq1nhnd7yYYnosZwB86xjPDYhksOW9YdxBxd1X/tHlIJR3kCWse
uB+8WBrTMnI+6cCdsa8Cx3qmhJeMpLNIGQmdjhNc7hrSQC87bjfvJCSmtz1cn3+D
oHoHOK23peBkXIHrGlgPttF1YUB30IpqtJReiqUM3VuTQLBkJGcOq2Kxsb3t8biL
n/TqeHHqcCSXwLKjEAhZfG+oKwzs846Ij009ytivFgRPEvuwk5Y/AJCABAz2TRwU
YZHcoFv6jW29Z0uFEBMmdQ==
`pragma protect end_protected
