// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:29 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
WdoL+w1NCGl1RTk+iJEywBY+rkRmma+Q9s02gYwpqXFSGXWpS9RBwZSKcC8mMNH5
xmuFQNVHDY+lpwhR1kMLXoDL56pCFpJNibigGFrPpOxJ4naDXkUIxpouhFCwlL/Z
kWiQbOyDoaRDVhtI08OF2rWa2CQYQ/LvmD0UrPY0KeU=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5600)
uPiQEg7Ro3SCpaS8fHYXBIbnQO1ODFUWH1drpx/yeZ4zyAet87osxnU+WX2eYZqw
wrTnGSEIj2G+3i8ZvWdHX3pOoLXq1AzhL5sn2py1DHsBMgQnI7Dc8Q/60YNNqSBK
ZHTfa8vinvtd1YMVoqGUgFoWbJvVjjyIyMWnuWO/0gFe23OHfa2je1YEKbkuCA/e
0XOJ8FFmoIwMgWf3qQqVXY8XgnDl6SC6pJjjDlslsnDEOEVN2duVoXn8DhJwDPWX
1LS4ezDBIqsaCLMUtaiqL+0X0XPH0cwEdZihrDNp02Mlhdqhvi8zMdK4lxir/Z+s
Yme4dP374jQpT6keo5sMj0uIx4w38r3xBwWvdadj6TqtyTKRwNjGjpqFquVwtpz6
7PUfRWys4dxON4AeUVXXo9Eclj5QWrb7kg7x7j1EUT+kfQWGhff+vA1BNijEjSmY
+fyfU7H1l+Eid2Z/PosNGNcDVEVamgIAizqErCIkSzs5oSGGxy61qE+5KKMXDyKi
HZYP/iiAmQ7WwzVKcvMtdzVAvt8O4AfIBbmX8fTwBhrYSrhCMfDINDuE2JxjpoXW
yfClJMshPP4ARkhFy7yh0tYKsAluHm4gVhTzxzNp0Rc1lAvDcRg/b1eu6IHCieRi
s7rP9AV643bvT1wcovyLthx+UFT7JI6tc933P+bx3kNyXCQCvb/jfmaIUDseXEZv
NbSE9s/1CYY1cFw+X9f3FZcdTXfDLogBOx36Dz6gjkIvNMFuOVGWcfj8/rG67yMA
anVqBtAaNiKTC9SvxhrNWzoqwBVZKstQqHjJ9R54cz19D+O+WEPBTnsOk7oL3WB0
EUgqd3/5EfhFMjjRnzXgLu/mxxuhpionF+Sa8W1jC1Ji3dlSkvzrL+Xt0zi+E1g6
vUxx83fONxy8i0MT/WkNzaV4jMvhGxRZORa2VY6a1V1HoqGWam6LB57ck7sEXnLU
/wnbGnSqKzens9rs0QihNs1BwcLF6ZtTxIiCpHn/VqmqRgJA70tqreJKGNDQn2dR
oer6haIBJIQM+849j4gcXmtCQTgk7qwXDkSe368+BQJ01+TdCX6AWo46hHzc/Lx7
3lWBq1m/bHvQ9M5wTGJGvHjwZONyzWN/tTohgUGN80EnQIw+l3oRdzLjvmrzl4QG
1ENViIMUWIS99DB1UDV6JynK2qf3z1bC0A5w50TvVVnr++umeDucjtUJFDpQVD7K
Ad+Wpe+JLRU6frKX97ut72iGENRfARJsLygQ36wlBEtt8k/07muNdP7WGJ9wS8B5
4lz8paJ8Sz9CSux69xOItjFj/iHTAyZ8mWu3MJ67Pezt20zyC0qQLQBaq0YoaUPF
aYO0ciebJWhg1Z4nvCOUo/rE9WnfJzKq4p5v2oBs0sKb6cLDg+VRHvBLx29F9Kae
x02Thy2OTy1ls70/nQtJeVcVIR2zV3n5+//OR0Q65fh/AUYelWAbkmv6wf4DiD1g
1XgcvwIlkPXX8RaWtWuDdXZPrgBv+M68nIjKQ+eliRahQ4mqtlW6ecLkLhZjudlR
0A4RF3c0gNiWAjaIN8CkFzGuiGwYCrhWjRuIez33VpU7uUao83FFwS/DkcQn9Phv
IjHmvyAG33j5kT0+aTMbx5qJ945txHHOnKHjZqhFrgbGOEnVC8Gc3EKl4gjlm7fS
RP7HwO//5W2e5wJMlbEoDvzNqWs6q+wawSj3u4tsvhOcgX0JNoDkp6CDHfvkOmJ0
f0LXDR1YN4ie717jS7I38LRwPs345NQ2CJ/znAGulCSpqpHbWHtVb1b38zUcoCmu
iO+4edqiFSMLMB8dlF+8jFh+14DM0KzuGr+3Cw2KHJhIyWiA/cPtABtYK87ZPb4P
xvc/hUlWEne07bRSrfMCRyd2A/MFmWyyybpa33OT40S2KWxBupEnfyjFawM6984x
TJf3a6QBVXcb20mFPWvooFr8uigPDBIEEqSVBghkhAHWQd7HjeJmV8cvUCoHqWKM
oCdqsGSbKM48j6itlM7dpFNJA/o/g7b2LBQKdtvM/iggmiWniIkyE8A4ixtQC5Xa
2nnPfOMIDwmBXMXNSsXra+E1koIVzFUz51qfXDTHWPIB7lAvg0wOzWVyu4d9zWRQ
ze7SjM2ZdRFOo/AGRQAGfUh4JqhjwMIsu5GlsJhWojrIiZ38aPEDUd/YLNU1jrko
O6tvOrmLZBTkk1b8ZoKr6ehqK8Lbt1Th86qYyKyBbBq4iFk0bfQEBHa73K2wbFGD
R8NBDbkB9XF0DYw0FG18Q1RLxAsnHUP8i/gp9/1R/JOefaUntaN72Kl+OmWnVxpH
AjaXhdaacUytbV12coDF35+MDKJkpi6FJYNgJu9QHj05rKLT8v5lZ4nNyp26U8nS
kM2sST4/g+ZEhuPDlj2rjgT5glXSdQsnCArNKYp3BXpb0/HMXLBoSRUzJGlmhgaz
X1VfQ8G8n1PSLlIa2z019WikuBOuN8KAgvrTXiFTLEcp03nxtvN6Ud+Ugs2Neg9Y
eqOs246JLzkExSHts7aHQIeRHNOegQq7ai34HgpU8Wf79AHmTk5kanG5TzUMGg+z
NxpxygT2jHpVIx1DzdQf26lsIYrO1Vp0Gs4EU49ODlrQGKWFkTSwfRyTk9N0lDBg
jprlUfLNGN2gYa5eOx0rKHWSuh1h865TqWd80sOXCgH3Q4f5TfPNgOmErN3Fr5Vu
qtdSNeznRPWLKDYBflC9MoBy6dZkjKS9lrVETIfzVG6ZplLZdPwihk5mc+LF9VYK
4rDkX9qGBZwH2H5SDSXBYs15UoPIOmugPcXTpDxwXs7Vq4rqdzhQYEtgznycBa11
M5qC/VuNRp1JmH7n/wVWfPmR+krle312YPqawi/tIvzQnur5YXZPfcZ6xzsthOuA
Q94VeiRPw3QoV7lRXZHfkDXmFiwk8KFvaiTWQujyZbQAiZKcrgPr3r8MOPee1zEk
mGFC7/RvpaV2mIh8Wy2VgqHvkv5IzFEnbyn9E1//gdVpRghTT8IikzVDSYHqGtMI
49kopzY0HT8bYaBkTdyAFAm8dlgbcdkfA4KGsA7SR8WX+YhNvPgYNUNYg23o+rr0
wbktYfL3MYJnYeGWWEJZYjw9AmH5SfrlE7jko6VYEJ0Kn/kYP30+5W8rwb1PAiD5
vVTtO0wc8K0KrEbuYvUdlKNjW8TCEy7oid1Z3NhK/Fl8tAhdxFQkcLz1n27tYqqp
xDJkblv/VWqsF60XxRQaOm/56v0gsSaFk7ZgDrmnrlkn/sKpRXZvXYF9xyVCDSHl
1jdvIh5rW1NIKRoDP6dsqtXjypbyLefLimofjZWPF9z/r1PeZJr6epXBlYPivBfP
uj61EsuY2ZjGZKhhKiOp7ppaxF3hxl5n0qGNGDJKw3uar1qrObyI6LG3xbZlBGTy
1bnKmpTXFEycEgb8ZZ/3KaqPPvXQBKi2F8LAy+F1VqKjH7r8VVjbyybcNoqKrj1r
f/GYEWmMrGYMeSedeQCmmMzpSBrX5r6nmRBN7CQMYQWNN7+3/BLK0ZHZ9i3nvNbo
a+JpU8SQAnwTeFuFuqu6M/NLeGUdMyx92TfWI8nH+p3i4NALrUWO0vxlDP+kClM5
t5HEFjyhpiMXXDFemp4qdGiWfUOgO2ITZLr9jMT/9vm3LN28IiscRp3VxFQxXRXk
LhXRNvmoMCPc+fOAv79sjbdVNFTWavFsYiFNkV4E0I7Ix+wz68Lic0d1wonBFRA6
MB71Ys/SVhe6F0/MFm2xgqnivEptPQgRZhdlV0sauNJGGoRvABHshJ/Z/NeZEpbf
eCgFjQpDSMg0WY92S759LXUx0PdhOjCa/Pq5G97DZv+xFy0V9AIL514GAWT1kRac
TCyNQZT2WJL9XK6LD1vSpNXBQ3tmywWK4V/RqLgBE3gFC4ILLtT0MworwiBZEqxD
H0lJgKAqzQ9bbDxHNzzf2CpCuFMiVU8PeaDdrY4jkr5qPT8TiKS9t4GnX2A3qX2j
PF1QLKCcEWx5KeLAIwUiWr21JBsc1hgHOFgSNGnnaNfcX+SxO20JVRjvax//PqVH
HO0SvIL5Q2P/s7syHjmDk9lul/Kvqb1z7yYcI5ccTT3Cv5dJAw0e1RWk1Xvw7cU0
pvyyxW+eO24W4qk6tEKG1ekce0/o8LmPXIPPpSnQoTnkaWoEgY8sbhANjdcghnZb
1tDevyNgURrWNxqhYxKdsqSyBosVoXC+xihdUasMdsuuDRscqs9zhenqaracLRNv
U/Euvj+2AGfcQvYbZmIWUxJGeW5eXpa45LHQOjeuvb7e0yNFkTzAjuA1I3lUhnmz
AuBNsZWUFgm/h7WdnxEBqp1cteWPn3UP1ndN3I9+63m2kepn7ddsr5+++R+rjWpv
bmyz7PMRyrUe08F7NjTdD/WqnrxF4XJvo+C5k+A0gSlktLU6JnTqHZP9tbVxfiNd
FF7OOLegex5ORuRwl3C7st2RweGCLwQFzE8Vs6V/gO5QcsC3x8km8Za7GUvjUeCd
PlQc00UGQMUauRvJFJhMnTW8bOaY4/p3DX6sT2Gax7eE8zcP3JkZus7tBcD6z2C+
avB/FfYd0UF/356QJ3F4T5N/y2nvUMyids5GmTHcsMnlsSshJ1OmP1hOyRYHXdcI
8PHFzLVX6y6MVVx++XMDZcyFdpeSrpNzaxvvemkLkckdutVllbHwngfKV9A7a1ql
I5Pu+lPO6grfYgw+5vm5yN5xLzL0Wgm6L7nCi42XXHI8oIyu27+YjoeYhzT+tZgs
5qlezTPryQQqq//PcmcGO3PY05lHxIdpV91fAQw6ijQMJYRlG9IEjH1p1usp/j1w
DZGY3/5XJDKDOtpD+HVwMArUdEwiDzhJI0UqQJ9VXISzQf8P/s/C2VFArxw3AlqU
/Z/eXy7oiLmhO+BGdWsjbxnlKODkJWB+wV+fHhsM0BYXlQxoWWW2IcEs4yEqBIA1
xPEnUaSvMSfJO8GuwVSRR1jU5El5zUwZW9VvKqCECIktBPvbjYw9ZWJGATVriARm
O3ZwhlvnTVy8mFVD3LO/TyIWi9vhRukoxrXdpH8BzAKTqLIglCTYXEeF573OFclt
R9+BWvlQDwIdfv8NF8grusq+nfFe7OrnacolvgEnU+J7qGsNkVvubvlOEZC2SpRC
1L3xyuyszrFPPAnqXeQAvwpDPSjdteKyiyqcOeJ1ghZ1lKUfuLHRDwuRlR+vuiN6
86/xRnRwIONAyRuHgWDHK3wRZa08iYalRffLvtvB2R2Pf27R/oz5Ld9aQAl4cPXZ
/m0U7RL5xoDZDE9F6qMWsTSGLqyNVgSFZKHbUC1B0ePSvBLIXHk42TESHdmk5fQU
K1XbMd65HIkv3apRjVxLLHHEmQqfvROR0WXxbtSGvdu+QbZNlbmS4oi9yMA81E4F
eW128L8uvuMemwkpfwiHjvRD8kZU7baq8AA53Xj34KXKBG6kfa8xokTLjcsMtVtu
XoTPIOik3S1hTPNkHmbti2hBYzoTn2kWOOakNYSLCQCT6nYVIUk0taF5XJZDvAhK
7MNTxrnjiYBj6bWyd4u900eHHFypA3i3pTFff+Egjownk1SWKQIARMNHKkkdHA0u
U/Nan706WnVRBE1Xuu79ZsX3ptYN6tjJZ6rWf4pAOquNT9EHHh8rVwIVZCcfTKyR
jgCiQddDvBpMx8qsfnBji0tKfIFtTIiYJIwchYSotoM66z4h1JwQts8Cg/8yJ90n
uvJnjbV8TPgePGs/5eWq31gMSawoBl0LdHIXTocNC5xrc6fkClU2aGGJCuo8BN1Y
TypZHNI53ynq+jIvGGs2fPs41Ry9CTfbUEqhiUsPFXVhjTIa+L8P6/dICZTqHQ6U
s0ck03ukFt29kPXAAHJW4gLp0ZoWLA1koqNRS4LU97+8rOAIs4n8HQKRV6w8gjs+
7V5gsdLJciQGYkL7UxSUEa1Sry0LVv3IYkKs9iuJlRij8jEvyw1gZRY59k8OEsGX
Ug3MLSa/H3osEAXlNEeG2bHTV9J8Hg/TaYc06D77Rva1zEsQ+Uo8Agr7WKWaLWtA
JZqvhs27MPwFljPpg8xv0BrqV6R5Q7fJNJsffL0WHwnwpwkspoasrZt+vaPZYzYv
0j3ylIb9KhRFwQM0LMhXXJRhE+q0HknVMHyQzUx/qC1bpT5pevnQpWXDhwjtHzZN
ws+wB9uMFH9zWrTPgqU4s3ukDrCRLj68odG+O/IQunKrwsRZGBIQrJWeRBEx0lIz
OabSCWwN+Bmj6RWIDiBAUAQs2HMYZjAsBS37II43hTc5p8JEcszXwpmLLomfLLM9
id4KJsbE8hWIWOs71K9Hoc2xRBDdIshs3KU0eFSVqsfF897xKNmoJK4QprVo9/Ni
4/dQuGedfJEusqz65Oz1O1pHAAfWR9C2bBAbYwmDEfQHYnZo8HSTEPk7gPbsETlh
Sg9l5D/eEWoGEPshuNg4MZ1os7oaQ3IZm0rbkUpDH7WZwktwybmIdNlLItn4Kk/O
RgyA3g7NPeel8l7uaNzh5JCcmAXW62VoS8Ms0xff44wfEDpC8lkgbLF6Sr12PYCD
LhADXEn26sjAba3WAsun4z2JHeSTIA9/lZ3bODZDT1pjPX3+GE+ZNu9JxbmSluC/
gtbfL6NVOH3rZrXPiJz2BlbK3Y0FkybHpu3+QOAwJA3oe7LAjMp8RWVP/dfnRStz
fhIGkvBszAabsRRdkBdV6ikCpaSwFIEaN2wsD701l7RomAOeaewxXfU2DrTUjZs5
T/DD3DACoww47YM7KLgtGJEY/cs6qt3GHhG+6ZdTAZ86sygFfODitRGBwQopkWl1
Gnhjw5RyiBl4I+LcjvF6qWhUR8uNuYADbBYMyZ+kYlgeo9EFc5LLk97XNXv8jVDO
2Z07tDoZVxwQuxWnbdyvFcVbsArpyHXJDtK84OdaB5tukcsNNG3FXNJPusf67pwa
JT+F6+Wc5LLhf3e1DbeMnFj3EA+ykzoiAknc6mmRHvCYIcPRECMFToxyxNpVpGeZ
oDktC8/hSLEFra+Nb8r+gJeZf1L3mclDyXHCMmTlBg3o7BR1olMuuDR6EbBDjjEZ
TiDpuLT4w4N3L06QH2Gsf6l2KbhseTgh7GS73nhq4AabKmvupH5NrDpx/ras6DlC
kGTSHI85zVddwFWESZpflfUmJa1qzh1mcEroE+3yho62Tc/YvIk3Q+gMwDQLB3tw
bd2H/iy5PPFzJuEQGYJoUpbDSMFULw9tvGwWAiGf5ine2rEDCBl5HDFEpxi5TXdy
4uocslBiV7rL/felbc7spKxWq3V+ikU/1ZlIxXJj7SXAiADtMVmPPVo9IRDafPcq
YuMlqaSCFiipRsWp92j3rb++hhPpYbC5IM8/AoxRYzlR7bP4lo42msb3z5INKPZ9
1txT2NxXKLhP1RpYTc8I2+rF1z368kIZn4GNILY9AD35KM4CMGIU4hEfy5FGPGv6
taXhbHnPw/hSEjqX4QpdsS+Ldo7zqW+NTeWa0qWOXZ0=
`pragma protect end_protected
