// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:35:26 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
tASFtch2kf+9ze7Bmovw89ggCCHKds7Ke9uTCbFjMnauACQhcZeAq+dJUiKch5zh
nRqWzBl5c5TS9nMv+M9VigTsX+Eg3QrQgUWxPajl/C+sa6NwcCObHDwrgin0R8HT
esQj8TteKQJUr+ZromNOXy7mCw4bNY6Mh3VYUoKL+Ps=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 7376)
TJlfKRyhBQW0aKDFNw5dhTee1YwR17Z/bE6+KqlsXYXRTWvZZRw+UqfOAQ72PkRC
Mr2gfhlpqjLMu4C/hRDymCSB2XTWPUdCwU9Oj7h8caeDcaciWNWEmCy1ei8QwXnn
fR4NwCobB1sVdi6w8g+rjDVRfabhv4nxaolgHYERXxMEaEXdxQEImoziN/QtGE2x
i/kurQSbK3ke5YEIU95G76jjv6aJvC2f2mwqoMaXYI9wlcuO5w4dHNoMPhQPM7PM
l6YZMQ7UZcsCXqFxpBc2tOde8cjJnSBxOgAU6vgejUMnl6wNZlL/15FOcMhvhLH2
KgTXK+g2q7dO/hZoaReH022Ld0+kDy59yJSqlSBtkQLtCnpCaLuxtNMslkJ2j+UF
4yucvHBL+Vt7EqJpBgAQcxhKZcQRSHwtEO8zwvgrDd0LOwK/yV/nAfxfO9AWH+ar
o4Rk3sEtgzbGjtArsRTVmmH765k3eRBrCjxD5yarMQH7hiqf4BUIAdya1lXXGqeE
U9HX0RtHcINT6I10ltbkPa8vVQkJ1Ny2uWRjefwAJ/QPqb7aWd04tUAiQA4AzL6K
rIxK+FceHydEM44zjVfCnpRcnnTsOhvvRA0BgIkzXuTh0E9RbbFNifAPDGJnzC75
Y8nC1bt/uqcyvFQ/foEQrNqLY+AYu61F40fZfPTXE1jisoeoI0UXcf/PaE4sP82J
ABeqqdmJ5GmF7RiZpe/yviRKhj+kJHzjJ0t2MoAhFnfohekg1EGYHW/6EtDSg8FU
QtfU4b+1Ic+YCl3HvW+TTsEWJTdiET5+2f8UK7vrtsmNmsD6fgyi1wWQYTa4A1LC
FlCEJfhTfsW+IVRxOowkmt3AqZY3obitUGpQjhSZG27s0iBMd/toN2i5rShcG/Qx
ABtiHUmUqMVm/MXddyPQ38noj8/pOVK7eUrYJfbbXqa3y47oWSmyFcI8JuAB3Imd
VaI07s3ioGG6qnPHniAloqCbCOFRvoUcdHGMlk4lhV6kGxyGHjxuraDpAWW4DDYY
A1pqiynfM8nSqASe+BNsijK3GIxir/9csJmzH+ekL74VpVfdUmxe1XZcUP/wZ1Xw
Gu2m5i1tkZRspZ+8qqV3ji0Gh++145cWGRoGXZU8mGmJ4+SCmkgU8H17fwDmKsA1
KBGVsYqxZL+98mrZ8Wz/z3ugPWVAyJg5hFH3DH0v+mp+Nxl9koDRt775998S8cEH
Dggr2oeJXfLk2P1ovtFonjMs7w8KOB6pyNhlgIa2YM9EMGaeAbYtcetgjNKb3KLW
pTwuf1ho//kRPv02A8eimwKTbnwPioZ41alCXHV34/m1wIahncsadmEyq8Qnwanl
29XsSRmuWdfBJbtwzXoF7UYKo+mnyROCrAYMZZn55s9yXBSF1JrrHVNUGiFSYumf
gzQaQe9mzSk4HFS+LTB5+O8CQClsMcNGiRvQTsvsVJgautLf7l5yJjr6+3nz76UH
VWA3ideVQvzzKwTw/gSjr/2iNEVk+VdZ2bb2FIXctKJ5TIQtFuhqhKef5yj7Pibg
LWYrUrPn15pZM7dUCeAzsJhlSbFkpbpSvPW30qZEvvLdruH50bzrPKeNvAt585gA
eXrR/PiTwsosfpSXr1LKOItCbkQSMFhiJRXee+zqi5qkL7qlAosT4fVwHMO9pv0e
2bU9+WQMXfN63OqeOh4MK1BfjcgGESG+F1ZIzm1TOOIjoWw+gD5Fw6V2jnTZNnZb
ynG5QnOCkdDmVUjNGEB8QSAEfIigVDEz3OhI9dvsU9/SpmEsBiVrCS46M8dFlvhB
/EOjvlvZ37HsK+oe7IjQLZFfvP8RwPUorbA1bGSSecaEHm+cfvFyiYgF7sGaZBhB
eqChDfmIlbw7yT1+8i7XoRg5SzGWYdb2o2BJ3n8sluKeqZMjK+ROQvnXacsGkEAf
XvM5F1j/qe1XjfQpRSSpTF9EhBzYlYDP+9UXWhAwrCYE3nBjM0laGSkwbA1Obj41
mTLUM9+3U//upI7ZPEnhvsgLDCkm1jcNPgfv76UZUHaWr6zZyQDLAu4qR69af2ZX
tzXWJMz62yEzufuvSvsDPY1ODxonxC0C4s1W9ehZIIeCPTdmDl3xUzfdxyiJnHm5
l5OJbEZ4mvovVfw55wkxnJ21aYMVOdCfPAvxkZbHH0ZcS4yzXQRIu4TnQhrFSDig
V87rgm8q1wmv+Sm6ZeSfW341il+XFaBTULhi0BzYfyj+7MWmesPxxNbZA7OVbpn0
9u88ytsoSpgywsu2f8wxMqMXINoua/PItwk65I7h1mVRyGoMuNawLLAeIbqdvhkK
oQbwa8u0Z1y9gv9NLcoBTg/UsTB3AHj8vPsft1mYpWZO/SNGQ2IcXJqmq5yQk4fN
rIrqay5JIvNyKtEEBeOUTwVO9GlgpOuA2fwrvYo0Mpcb4jMr5cSVXS4FOqFGnE4z
zX+5bAsy6DK67jhuWHCZMTFhWhvfe/XSGkt8HYQAoA8+NmzxprnQBxxfn6YmwVS0
J1ryA5amHLGo1K0GZEK//8SRKiDAXIJgArQaC4eLDerPsIOqX5gHNNY3ZUm2B+Gp
mRBrdZvW1XolI957hm5o/4gJXLgw118xAEuky8fFqa+5vOImhYm5MMGP1xfdbN7p
tv0i7JbsIlpiH5FlA2j6P6HAc6DCYzchG4cfWomsdwhH7sCKewNs8ohyx6gnfFFA
rPdvwlQCFPpHeK8Yct8zLHe2b7U63OrpDLvK1fuYfrZ6mlkFmAWduZWdzvzMfpiS
MvUlcmo04AOX2S2Rj/PfO01lUlYXT0MsYlG6yCmMPzuUuQR70uCeHvFBqZVF68rA
+2DV4bpUPTRKYZhknEPcBTI+iZTT4LUxQmNYWwJVNqNpdFMvtG3aY9m5za/WKlVp
QfWt4L7OzmXjCytdu7iIZyK178puHfe4RTsTetbZX9/xCePpXYbSHQ/OU9YbFLsa
c/LvwrnVmYydISU84b54kcBSQlsjtEm2140z0JKLH1cGKdc01mKRhe+hMV37mtnZ
4NmyB5NYmokgxQE4bq2MOkaqIFN8Pcd+DLOycfu0wntN4u4NKC8yawys2p4Ly/7C
H1jJHFGh0noJM2dqWa1w1LbPq4U4Xt5lEL8rKDyiRu8NMZe26EvWqkz49htBr1MR
aQf+bZOVm2AU4s89U1mlbiXvSFUAE+uCUbZHIGnUJemk6nX2wDL2KnK+VD6ENzGk
S/g1rWmOqXcSKBR6FHDXr38H7ResJIj5g0+U4jO/WzWPG3wev5eKuFcBM/3jKco+
Hz/YHxXJfXVIpFA8DxQR5IACUI3GM3rZvbpkRMtxOkW8fI2MBfrWKDndoBMtdXdN
s/NSfiLZ4a5S5jYX+SKqj7Z7KA160fcgEO1agYZLyMRFqtWWUjB3iIX0M7m7G4AT
kjLfSW+iZqop73M2uqHG8OPtRwYnFkCBw2TwYkX8ecarjbZ38vJyXCPsJ0aHK9Jh
8SZaqWotDeoREGQRxEEWP4ruGW3zsmb+NxqIQBYdwdJUxL726WuwlUGyIzN1m9Fa
pkPF02uQIigm6i7oCT2ehVWjdy7qmw9LbwT82k7R0nrW5SWw9cYrtCXfAEGLooHy
icZv/f5op6I79PV5BZ7+tjBPIOF3ccDuacn02zS89b26xNgvJXYb4IhgjH/8n9v7
2w8RRnf8iOjw5l3JH2slgHTFlmwNmCK86IqczzaFcsoWus6qu7L49F9HUuObU64Z
evplGd6wt2oUDVnXv7jnD7lr/KhPheAU8PDhowx14IF0Wd3SkwMHxgouYcAORhYD
3tsSBIu3qfAr2LBHcsunUuArP8q25RQ0dTN+gAyJSM8w6SPrM2R0tYiSUliVhVD9
4LE0wOmAZkCbb0KWluRRzLXY1jYs5Jh+UxymDj3rODuWS61TblTgzufcChKBcHzt
5V9MsQosd1i2+71/DB5KM8IDC0+dgRXtTD5sS600ZHrpJonB+XXwvnWeJhAdSLOH
Glm1YIN5uIiLmde1AibcCXVVs1+tHui/W1MimqX5zc4R+CJidDygyhuZCVuhvzyj
iOvc3ZgSfWO9CihnjdRD+mg8212TbFyKanQq6keVsy51bzIEHWAFpx6kNaNP1f1d
9ZwPY9L2tAGBr0M6Eox0mF+2O6IyYyqdkg/01HIsLGK5wfOgBFP6bdUoTquU/xwc
Z3WJyjA/gxI568SxPyD0i/ngNVYkmKC8/BEKHEAeb1gi6xGeobgXhw/h1BlHs8KE
yic0gSNCC9VJ1ajKURBahJC1SiireT/oksxMDzW1O4WJ5aYNx8NEOPL8Q6fM9AXi
UjEmg31L9feErfsffbn8t0sAEMvE7jkJhzmRPWiXUh5pttp3XWsEVdsdc7Di5dFb
mhGVKfbqEvlda3h+aQ6rdxWxn6AZ4adyxPEGkBqNv0BuuZtWaiaxyV7mtwUSvomL
DwUOqgdwAaACfVf7XfoE26YtI5UbMH/5H5mFdUH5BWCLnYugFQkCqzFseIBZ4BfE
p/gWBOfveyI50Ciowyzt1ORMvJXKhtLBW3gGBHxF49C26RL6wKkuyTXG0QJNpM9D
IrPTywQ1YckKtdYTtShxy+5JMEUslIRMffc/YMAbVQz29ncNieN1YaydOEG2knAj
SGQ9iwtr7bdnkyYZcTDVDTmB4IiOkgSWOXhOnv5xnrBYiatsF5rKnYA4GdG3Nffw
RFJIZQpEL/vFQ6hV2LZZHuriHYSVLF6XfTNv/0gDMOOiq241aGkqP5Zc/s1jdeGi
JQax83o+9LWUYXDyBp7dtw9Mz4f9NHvnLn/hU9WOijmvm1SJI14rAlay1yC9iQPM
hh8IWnDfMBc7URtmE4PcOyaoMFRTGezgr4LEb9/7ZAJK5CGyuYl7mSIz+4Gd0xX5
8jwd80x4E3wDEU/PKgz8aDhoiw+AtLVwCJgfHbHM86PidrqrUEL7w52iO/vK2eIw
f2k/AwQhJzi51JYsd/oiKCNBdfRuaaZawGVS3P/SzUA3gALSKSDoeVkgB5JgEmEx
kY2lRvD+6oPHNI0YCHrFybl+JLfxLXCMCgAUCjZUuDUrzaD0dOjj9PUaRw/zYprs
NqipTpUeAO/GEurwLuSB534IHUjytOzK3s+GXixTGPkB1SQXT8wk1d31Um16gsFb
qBhFn5VKrCV6BpH4tsiKPXLY0E/xXW9+dB48q0VMy0CtoaR3sdZ5EoTV6yT8NLXs
od0WMUSaK4LuLaNngW0LtdmK1RnmRUh4hQUUOz/XVZiogEDAdPHpv9xwoBEBgcLo
zYmBGvh1mXZLJGMOJZkcNSJE4RcXLnkrW6sDNBMeC5JxfyakcD2QVYURvCsFOTix
CFmZnlzuVF6360B+l60I7MADXd8RSP/CtALfDn6smT/45g9cU0+m/rA4oU3xdpUG
6izqt3Xs1pfRsYhMe9AkjrjgSCloNIyf6I41hRXhe94iLcrdOUsVsNS0cKqV4jU9
CfmelD90TIUiaJb8li89OKmxWBBUjreP+4IG25X+iHoRoTlGSIWP8+wUXRAWoItd
ny6VH13qNQYBtzKokKNS1Kfqzm488/JAwQRCXI12LZu61QDe9wtJbW9Cn/V2lNWW
DCcgiIziqgu3JdLIKS/xsGX8oAcX1m4dWeTHOeBMpDO/ekh3TK2alX5787QqNgWl
eRhkWSSjsCsV/xFcn85TAi91vAPo1bXxPY1n+7NApl0pzwVyuxnpTCRCNoWvKH6p
J0Xn8aV8NBu8ASPWUcB/uGV7sUa+ItfllGwzXLn1HQcAR1bs913GabzylfKZwXQm
AJv04uwOM8jIKM2vWZy4auz/oy4DWrWkwdy13CbsBgKaZFAXPA6G0bCq+YN1dMp0
JRmWLIO1aTLbHTOImgUCexfdQ8VGuz6qW2PYKzWrcrc888pbTCUbEXVEIv162/Ew
3jQSKUAmI2ZxmRqq70TE9N7D3tKzxzFmG4WBP2URs7/91liMaYAsQUBiKieltdRo
TK8u7qnsBSM042FBa2FsugaLlmxpI6bOuZR00x6MoagPHQxUcrh1YNa7f1M/y1nH
O7th7j2gseBjk2Jyy2NF8s6a0ZfoZYCZXyKNbzQmqMZyFYTlWKE97wf9AdfsGB8k
vt9gx0onhGBd0X2hKkyYYsmhiaKBMyFgggVpAWBpW0woUC35iZiQM7aK6kDuhHaV
xtRzRBf/FlP4cMHDq5UTPGpLYBb7j8MWgvaQWFaAmH8GBjReORPSL05Qw/FdKoaC
z8YMTT8le5x905sW/kMIOC3+HC6hD3NfbsSqBMoOCg6UniM6UyX0d82gOtPLFCiq
bYnCrxAA1efHENWGgPVslHiKFp/Bi3JyKGg5H+JFgHOIulFWnHISoqecqqClhpXQ
RPSgc0S9BibH/Iiulst0HPPN9frCGUuZ5JYL25gyEEe1vkWvlMgg0OszA6T41AA5
vGcclVGNE0yufzqJ8p3hiP3Esr21cFeXCmsjlDV1HKjb9x3+eaaJoxg2bFZolzQ5
TeZVBhmfbHkWFFS3Uf56hHDfFRoRt853S+eMMVEFDeyAaZSWKv7IP+xEHKI/e40x
IFfxfGTLu6SAyAM+J10VlJNc0lylZZhF+fVm4KprM+fW55MXgO4guddKm8srMG7j
8MBwZL1hm96YC91E5EnPU/4Lgg3owq1c+bScw8jYaoDqoTBxChsjLz+RwhY3tpWz
hfhJJUGsUxLGqbOJ4WMEibwHXQHCjzONRuYu2fT+nd7xRYIuMQyoFA1FepJEGiYG
zX6pfKynIXYTfMxPAptooc/Ego59YitcugMr/nZRqN+gMSPamagB5MrglzvUz0Qn
++06TmxpOD5OLDcW/9j40Wr22dYj4HaVEX71YNHFfXpFTLxhaWqm5VGQX52X+bxE
b1SuHb1Pyel0YovCl/SZ8PeLJGUUCT1pAuyANOBDErDBZ0XHLwKc/TU5j+hlOpf1
Y52xR/LvoXnW/n4fYz8uJBaa8a/IlRV0emoIp7JlZ1gbIE3bjEdNrpZQuKi2gqPH
nKmvHr1u0mkBSbreTv+Ol9lZSRTlc0gaQj1Vyru79Qdnww4OTb7kxuIAY2qgbDBT
H9+sQ1UiIUUmS7L3Bw2XYfeAYxyjzIjx9faTeX0L08F83QS5NkU0iKE8zQ6Q8OXi
O9Ahep43GFvK6iXjETez3dpB0ZWGL3eMtuxsWd95n+tvU96MQMR0y0IqPARGIeay
/9Azipf0jrkkTqdqQNWo1wGEPk2auSf+biuURNmUV7Hrr9FOEF+dGCnCcZwJR2Md
sioI/KVmAtzcwHlSTL6HMEqBYOW+UEWLYzsFmv8QInv5GELBt3EK2gfZPAWtA9FZ
0jqs88EMD8jy/PtbBrJjU2YvJz8h+aEaPbvtnutQoCPQglF1Bmv11zAMDuua4TMF
tKuuJjvuLUT04e3vzfuzAzz1HLuazeRsEuYeM9lo9L1rHFqz9cyDR+QLqcVADZhS
M9jfNrl0GCsYNsgrxz47egfA+rJjZC9ttHTmktStUu0Jq5DhUw5w2wMjZuSYAoNY
c6LnFNGX+Y/LrMgZgyknGczduyKgCO3wvPXWf9gwCijIpDcsS9zpPhAnEjeIoVkb
+ShKFptFZ10f1mMPNPEbAJBccZfAbDrKHYqVaOdfO/v1YyE9RUD8+1kuk8q8LNl3
VCogZR3Mncxv7i55fUdhkGsAygtmTke0+yUMmXvOD3jaMlqDtxx6jiUbXEJHJIlK
G4qoLRcaMX9qW5tccKEjtuWokrUPZkGCVq+mxEJGowRFB94t+mvtuHc74Lr7Qz3m
Wdy05uDEHvSqvSWpOEkaqxgB53rYArSD6Pi3eKHxoL2SP98RQHYH2kyJRhzz4yFw
pbuN+ObdhhwGe6iTY3sjX8PVuqKpauSol14gfZQT/nJWZdTiyGFdGehE9tcZJRpr
hcuwN+BGWIrP0N6X5vKdQWreCHH70gZDbLZ4hhP46/jrRfv79sjFG2LWMbGTgyeH
caXfyB0D7BXrIWqBgGzVVNVQSk95yskoYrhtcTit52JQ0d8dhnkQjyir7ZSgxCCu
ebTMn7HfR55A01Gd1ZtY5T0TILtCwwRLZIu1JMqMR6j8csaEa4RO/wkh9jnkCXo7
2qkKA8Xp7PSD6/I0d8x2LGcwYgzQQE5/lfsUuWjguVO05w8x9sS8LeZXNsZibR0L
tnetdKE0R6jecRYjKyv+gluCTxJ97crgvCMrrGg+bC9mBSgKYAEyczLUpB1AhYX/
/+lgjX/pAGhp62XLkBGHRAep7/XJE/4sTmlzldPXpPfXWKWiKHXd63CD6pAzKMd4
bSxbSEg8BdB6tqnAgrD0IyfMHRKp0HGipURo/yEXM7X1oBVpLoJDWtfCG7MXC7Kf
ihM/8kPBGemPOyLU7vZmFQpOMwfa1nDBdJ+lWwFy1aLAWDxr2CTS6y+n1v7BfeDv
WZps1i/ih5umZ/Ud5muQQn3X8H1vTbJ1fT52WfLTL7g6Idn2ZkgEnlhYE7smaXXM
wZCYRzHrB5Dbcqvd75myxSKR/+NavrCnxT+fOOEezr4uv9VlOzIEYqKXOIarM6+M
F6XxJ+gFwYlRKA1VaAb1ivage/hjTsUQV1BhLDPfNIQxY0mLds+foTt8sFBWbsBK
WVPJ9iS3MMuuBCQIly5Re+FpXs+D6S2aHpDRWnt5WS2cq+xdaKJp4ES5qwmFKWBE
HvyvIi4O9Hlz7aLkCooeikv4Xc9IX7El7qDyGmpj28mr1XjwGuF9aPjqIL7mnNvZ
x3q9qu3TxiAM0xTWZA6ZTSf7XjIiY/EMLqb6kFCVhNCB1QEriXzI9ScUuxjK3R+T
F+wcsH+xJTKZYsmMRM6rI9zQwH4kt4+6Fv1rMoFzQs8aXiBVDLjbEQ2nRX5rTAi7
ufqrOLHdWI59kbCA1xzg2YEI04WdXWtENOiuzNEnzjwukG/uyogTu9plUX/k4voV
9URhZW8lCORxzbKaRgDbr3ZilL68KJ6EfyqRG2ncg7H4ceu+8mRnP3Pgkz/BJw/U
mAmWyRi1V0mePV4iOuCAvdaAjWsECJXocaJzsJQoX/s5JZkgwA/DYp+CDhllLH+J
5hoBCiGWGSRAoknzLkierX/xZjq7Wq5Hjxtjmo6/KIYAll2Q2Ee0//ZB0NnQg+4O
4zxU/puozXntDcsiJOdWvgl78z1icM/Hs4Nx9Nmesi5s9vxfBCnK/FPWUIcazDdz
lx01F55rC2mPBFLPP1hEE6EhixSvBCVdS+BTdI/KexF7+Dph3laZFv3UqeGSP4hU
LeHM7VMtwtUzV2KlEW8BF7TFkfB8ApJtnp7H7tWI+gAz8ifBm5LMX36OFf5RwmFt
u4qaabcAVeuBSTV9gEYTAW3eRDQvP9z4If5zf288L4JcC0MFlTc7w06Sk5hT2nFe
+j+y1Rd9Srnp3mJ2eQE4JLDTWQkDIn6QPojbmUoOYESMAlmh62cA89oeLYVjrnxO
xO6y6rBWKrDsJ9n9WZ+ofYKgMCUvjaE58AL3nqXcgcGoXQgxe89UNSLr4coV349j
47a/xjQwhTxxnxEjMWa3Q7LowM+bR7rcmH1pZ+kyz0QInoMbKeKzIQoWxXKjMP5m
nOgS+Dm3E30qaN5p+t5gOmNHRvpt/RRwCTvDGlz7wdbJ69nAzC5Eg0xs8nmyMiev
y9Ui3D526Hsl/jcs0oMr1RumdrQRKY6yhBcsnG73jPTVRoemxnmKb9+tjSp0DOEq
y2j2zoEa2LHaZxHscpetU/qik0FRmnDZenFOSrvTDvCkmt0+0gbmAVARJCvS1R16
5oDM14NIcyr4Pq6QfOHRWJU/2YXqn0+FzXtuDsnLvUjrIm1sOvEDa8FGHb2/qtr9
rcLQEvIi2uZKeHzSBJiGd1HQgcw6fyRcr8HOgmCDdQc=
`pragma protect end_protected
