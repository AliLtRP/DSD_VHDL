// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:35:29 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
kYd2ZsQuZqI8DOZ7rvjXd6jMYQEdRycOzL06nIbgxS8G4eEhDiaJfKMV8SImeDJ2
RsayBYthFdO6w/gJqmLPEFH1CqdiKmPeswxLPc/ccTBWuK0ZKGlj0YpWLzXxaZk/
X2lWE/EawBesTgbuQ99AAXsH0lElV5faywLDgbUGq/4=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 10304)
pGoud8jpg34jclhb0ZdcS/UZsZjdneRwrrAkCHZ1RxSYhw1BPk17TY2URuN9gXn1
kwUv/EfhyqBo6mEhqZZJ83X/Uq0b+2HKqZDAHbvmxbjC99GVJv+FwO5aB0GfAG5N
k6T/h6yJuxWTzXk6Hfp9qF5pnEYZYxI36090ehxDBJJPk+9/ISG2vM2lRviODRwC
GdvteQIhHpS+U0fxjfYnbdZZ4wHtikXKw2kvNeu20kqorup6wibba3oyPn0NhqWL
n082tOwzX6YKuUeRlPOthpC3oHuIvsJgKCDYUHehl63Sn0YUcXj2CwK4ZumJ0+dC
bO01CMqre+4UCIY6EulZm6OqqrdxKEIg3jPw+F/wKVTAxRsvR+MYRAlkRALKIBYO
/+N3pFdCOBKzJA974tndhu4vAmZRyXlcLFcELRUudayUEIyrBAGqqyDtX4U0QX0z
kmOUiXH7kieviaO5I4+mNxbUYl3J8ZHFfC1mazJZ56pbMUhuAEMXppFOwoE3LHul
jeOgJxaUCUFhN2krRO6bCuhBQFMYhYnkWEdVyYDVo1EzOJ6bIDlFkFpurYW/4DdV
0krzap6v8bacjB1XrU5in+ecCKSaweeP8cLb2GFuW3SxghGnCcKpitCcpqFsQiR+
s4GgaC+oILIqNhVi8wTuPcTa59x8OutAzc0TMA/8T13x5VSz68WKIjANVO/+7bcO
xY9mgW3KbDTvEy7/awFDuooqI5BHQYxvid//QKJH0xa5jpOHPPWQAlakjNI9CbR1
Gc8QcvvCHPC4LuaTwScVyIJaVcCWjEsTbHZ05A8P65zYIcuLH44fQCKjpYMqvEZ6
ImCZLE5sc1FGt5CxXvj+jR5VQh3r1zSLkzuzda8qG07QlA4NpefF+irv9Lsrh5Wv
fi/g+kY+Me6yU9JyVu33SQbHFaXb+ys3Lnm2GNaqMTylSQWBOfPB85tGcjwEisdi
/B9Hs6p0c8AUvaOXVPrjvhz7bWpnm+RmPnR6+nVjGXFso9nH5MOyXAXwZ2ewOyiy
movjazctB7TIYCSMoyuG67LuOvmAvExXWhlh0kshLdZTXXc240ilD2V1d4s/IIOr
nHrrYIpW6tnQ0W/sV+tBwuudEKTukn19zvMA1TUn1Pc2eEPc2rBnMkntN+37h5Ux
htK43GJ+MC/6yVMSz8KG4GHU4dpE71QmrKB7FbtxvcXIAEajft3Ym5tq/z1jwaKH
h1PpAYLd+32eadwOjW/aQoyJ8tRtYl1rdBDx7hxiNzlHVEjNoy6xeog9S19Po8C6
H6bnCGlh73u2MozulEvq/wjlRCLJnVE/ZhvCsznLLO6ixkwHmNM9p8pt6X52zZzU
9mktDSXkooW+I0cbx7Uo99gqVDZmb43smJ2Jl0JpEYuymZQyZH48iK9DJypmBeCO
FlhdChcnrR2EZSrsnIqTARKru1I1Ba4V6dPhh867NsZLSRbMUZswnHb0Y3t5bZiA
zTUAPARDxXbMMD8TE/nEXDZnzzMqTJFgdi+LjqFY4bIAg9x1vuwdyUri/DkZMkOF
hqemUKvOZS/xmIajmwBX28GTRgZV/C9tZMqokbLT4v/1boBy3c4pJS/kyVMSd9C8
ucD2NUXjjrT9mQyxHRepN6Yfg6lCO13CDG55sQKUBYmbizS7uE9Q08AIjxBFApFn
pcIyTcn/NkzQoifwRziM7CIyx3SGgZxCVhSO2FSAeSaIYz+fGuLq0+BhzHoT/MUv
MtbaRImfqLvga/uHByQ7/uFb/js9B7JFAZIVacZaDp0KrkjGj7EVOrxa9dG1V6hW
3TbuOvMlOyXrT5Q54shWhL8Ca0DyUWyAUlMe3KZ2LF4iXGBI6uhXBmO00CYRkKpM
p6LlBx8aoQcGQcsg2XxsCFtzZwIhXOgrRVJdK4Mg9g03MA+BGrPSE5+MnKoAqy+0
zUDWprdkb2x8MJKdbnohg33yYMSBlHvonsEJo/Cj4kAWmiLMGSYwqJoAlU12WEzr
FO2WymjNvSozhGcRSht8PKcalBF8hwjlY+yM2NsyhrrIIk+Gbb3xAoy72eXkl1lh
A4FsndrGUZ9pzMK7qWadT9fNx5rlfAxCQr/166PZvOHmu1AtLlwWYh4lav3Y2Jyk
BwoPGn1KNESfVGmS9L4eTU7zC4Mnx+xb4BjM7vYjgbP9Dyg/1anMeA8JiugVNDH8
ucj/nQ3/LRGouQ3hhdWen+aCHTooUfrt6ufgzIN4NuPWaktp8m3Q/EmXpHUIRSdk
X6WlYMONR/nnzRwQlIIwbggGxEyIj95KqQHQj0yCw7kUBEoLMLsdfohme+GEUNr9
YekV0NmEWJC9X4c3end2w1EiBzMR9DIAw/B5HvWyv8psHS3qBn0NjcQdgqQ0sNN3
TovByL/++ABef2Q1uYoFQRGD+EbugP9UKSq3QoG5bL2wmnvyx5TkhhKSeuxNL7G0
qqpK1QD58bMhhp9R3ArGhpjmE0Y5VSxuxqxP4ntim211YwzacFO4Ne9Y0dzf4BwA
ndXaYljop23gHYtWl1zEYxKD4Hz4Kt0ETRH3Ali/6pT4OEhqp3muhgFTfcR46yHY
T7fqOrplDNdYKvyS9skt+UqaWPp5k9WVhq/WBnHXOS6wd5DSV9foy9CV4dLmQj9X
LjSMZC3yPgT3Yl2mQeWM66ZrNngPj6C4Op1HvEhjnY5vEhYQoSToyC409Bsa6z5F
7GrJ8QnbHOBIy5yDUO0+mdtKeoXZP0NToXL5S1ZT9KoKi5ChlQUuKalvUcjBvMzY
2h6N0alYDnOK3humwKMVIIVsSbgWt7eT4m3bT3ZHWgUGLY79q1oR2jdEgobuV+s/
hNgbsCM9qRj6nzudMS5dirGprNmGAHEJX3e4DFPn+sd9RGMgCZfvhfxQ7tfeGeo0
ZM3yBLpN4qEUxUGpuzvbcwycg/7gvyOFVxc/0aI6mVRQ/IB/cb7yDdEckfQLXpGg
n3bvmgvwGUqNUGtv8u9mlmgyl+NxtnC1cYxa85xS+5QiP4E4TTQo67881gz6R9xW
jo0TE+Uetr1dWlGY7KEE8HOXkiF7Sy4M5jeLtnjgRWCRTgGMJnnIHdJkH+MO3EBD
apLvZYFShbVAOYarf+qI5KzRTHc04V9F6KrAtqJAzcWX7PQls1j4N5nHxusTZP7C
l/c3ga6zB4C7y1oWUsamnDfY+BBXWciJwgpWWsW3wPXHzZXg2d0MP+NALafPIEiQ
S3CVDiHYrFpZpiU7EiL/dLpkLzo2buXAI4DvoASfs4/pWnfOqUSC+g7a+Be99LEX
kic3E7WAr9M7H/6XgvCBHvh0+r9V+EpE+3Nmtd+1orc52q3Sx9TBdWKrjrde4Cch
Sb3Jesq9wZkk8QqAYOMkygpfTkuz8JV9qz1g88s491w15tql1TSnsz9Z1EwyDqA2
Z71aAu6k+vaM7Ph6+/tJB1DWNaOw3Ho+1s6Co/91W9whDUGNrICAhZAr+gxevv9i
ZAAAS8CtJQ/EuudfaYf+h4aW6K+sKLgK1nKgsw4SLzSD/IE3wycrZ/A40SNK5Thl
EVwmwrQFA7u0zi6/8WvO3vsINTFd+EFXiChSJ+wCJ9Z7UpRrj50j6pio8M++hp/u
YGLzpolXF4EGvAR3BDDJ3QSDKESv96ovDmeE9oo9F+6fAafLt/8A1fYnbhBVLbRx
mPaxI5OyV7cyRam64ZCh6axaGFvEEotJf/L5HtpH1BBZu7EAKuNTPuIM9Jx3+q4Y
FbmpKdUHF0tB7vOs1Wm5lWMob60Orszpn79jjW4P/Wr26eeFwGTRP01Lnfg8ux+V
O0anK1mRVdWh7hdtU9zdDFzFbEe7blqfxWg3mReEhYax1yvoZoDoNWGL5EcTGQTt
gfDsErrOlp1BNnXaL2+FIEyuLTTNJgKWdASkO6Fp04LQAQcfi/PBgAvg6SGW58wq
X3NjpmKf+Mpnyiu6KC0I/ok5xKxUv18VZBlYa0grH4SAXnglmNe3dOz2nK43q7hV
H3gDEbAc3if0Iappkwmde1eNp9U32JNHuB5IVkvSLkh4aHDmO6jHCYg6u0iBFCww
eXNiZ9v+Te4NzOAX01dYaA1xTk5xkteLGgMnOz3AN/8I6MmzD6uIEg+qh8C2OF4R
F1LNaW1W1pQkJbLuxpKWbUZZaWtcUdW2LlZgSb0ZC+59dyms/p4qjl9d63/XdUAQ
hq63xdWi011JwZA/zNexSNj3Uifm/2/Fog8BN/5fk4KC6rbN2tDHmcvhmdWpvSwh
p3Dg+8MKl26/G6zR/r90tLzV2yBh8gk2nKiwes6YsF0yjkOWof9thd/cO2ucjesR
2QWwEg4Q6uXuxFyID+U97JhNx9xY/EWpdEUzT3y442sFwA5boXJ5rK+2AqWoW8+D
G7PevFeUARNZW3SrFmHUsrCHfzQoq3QEGSEJpWhQpdhvlqsVjHVEY06NZn/yzHua
4AE957K965zziN8DD+LdbKfVX3jKT8/Ftgtrhl/oVeLgTqH95HiQo6SsSNIbMe+O
LIwKN9c0zyhOQi1LRPZaIIG28VM5sQsMYPfdc+yrPRi69ZWySkYn1MCBNKrALHIw
h8EHBzNPUFadokQxRAgAXqGK+5w3B+YWsKWzyDB1OkVndKThSEfNG/rxGTKcCHVH
ibVuclvD4qVWlyVdYbNYQ+gtKAMx8EPa715sXCrimcvajk3f6K/j+INffH9WdiXZ
2dGOd0o5WlhpMhgQwhemnF0+dV+63rJbx5n59A//M4bP/Ork4xtQSftkcyKBq5J0
RTLawiz97rY1UbVNd/jVtTobWdnrEe7Gcn8r8qymrB3UWpq8VXDBTIGXlSxemBtB
tTK5xBf8Z/vbyQxISFYXY3uDD5HYfnlmDtzP23YJJuQZMf9FXOG1XvKNIwu4gWxy
/0+Zj5qwwYZQFz9CvjvzTznHx3fToAtiJYmS+n48Kaz+RIm34MHvNJBs1pYeOAf1
+pKDsNehJqMLb3kwIpLVvnnWsTPG/FJoxGzVzKI9iRUTCa+EJ5uClq2ZiPDsCCB/
5pJuM4iFNqxg6qkKuzJEU394/nqMda2z2nuRHvQDXyStJ387CUoBezusd9QpE9E2
YUxek3KBDihXJ1MMYPYLPc+nkW+5+H46N/lYMyUij3PhWKgbPQX7cwg4EPLyoyqc
PSY3xMiIwhrBXpLrEB4E6ZmFPdNigH2K3UTMs6flgmCkPzhHMpiFVijSP4Yffcmf
pw5yFkWqbokAyXldyN3HngTr/AgikCt0yRqne3x8FjAnVUk1NRWwGB0JzDykdZgi
aiCEbEbJmJfkoQU4bXEWm2JL64MshAyx945IX2kxOCClfPJnqTGRHZ4A3gJK8vu4
cw6+zcBcpGcgqB/AQtvC5DrMmoXPk1bDf0RbYKFZd6tbchFs4XbO8Rh1JyPt3Vgl
OjjwBSamCexexftr/hAUkK7AUDZ7KJf4BAty2D6SKtGGLBfv+A77lguQpf1fMPlA
yeQflAC478vMZwe6jCo+5jUmWW93AoDKxKQ6KtSKbQ7Nt8a9VzQGItYOZVaLgbgk
IDLl2wEtZwFOHqDdPcUS9CKpyecYLfFjSlAb9ok/C6uFIlkDC7VAYTZf4lAMb/YH
pfCkO7Um9lkPRpNArRsUEbFxiPR0nIeDkyE0zFLMRsXUHV+zsCjYkqCzUQnjnhKl
10/zwQpjYmUMi6w7NZHZuli2so++GKRe5+8gI7GxtZW8m56jiZklYB6A3Wr0l0On
CmAdVR7M01lp6a3ViBe21InVBUJ3npFet5JOf1i+98P4EC5au8+HCgg+vlrLoS5L
jYP3Oqw0p6v/+1nYwcEq5I0+D9SE3m/LPY5qvx329cegyo0lfmFKgPQtGbaLJ8Ks
rp7boeVs4I5iyptfoKi0O4stB4HEz9aaP4scg1HcGULzZzjzpt2/Vu2UZPzhNmUM
TEXtqMcJ+L5Ac9oMAspxCLwtxyizYnN9fr70pKZL9I+vzZ0s8dXgrshpBlp1MiqB
95ffurK9wVG0QDXNRuXKlEen61uU5yORTaiw7mQxzl1mLMMCFtv8BapFUVCs1Xh+
mvYeecs1pG0h9LayfCoFx4LTaVS8NxIvK7towaQR7thx/xwZAX5prbypH8zEtU9c
X5uOXlx3gawZr/u6xUKi21jbX4AXfOwB5fCt1552760XmLIcCvqESOUW14+NvlDM
GQbKJVTUKXNFy5RY2w+SVvOLpzlkaagJ9LAbJFC7M+G6sC4xeihoODmMzztvAkZm
S8htGNRJ56qcX4fOMRVSgmsXdT3MHRCe+WDc4KfBsfE7FcdmMQS6nZStP6AhU4en
uUQNCIUsoFFQaH5VeafDErecT33RZhhguwJvydR1HfkjmtcOaxQn/hapRb7Ar1AX
HWeUNvf2qUWtsE5kHHGYDeRI3Q+JfgClqrEIqzTmAiPHkvCfTJOxJVNm4XP8VsVQ
OKbbPPdb/0tqhlrLlmprLnArsFOpWwuTk1OGuPzVstf7WPm6DO30gC+9vVOn7ve7
uiiGb6Qg/oLTLrObrTiFUIqQpOLBPOo0jneaGF6RdL329hoeQNefAeUiUITfxVjo
q/EajUQlR9shtnhKQGPoUQqHcxzo7x39+Yffc1c88bxGc4riWXO5SrvADoq7IRdM
XBREG24Q8tH4FvYJ8XzgMuoKKgSSILJMsODGj8vFNqn4y5bKkrK7JgzS1ygwhK2k
hvICx6M1PO24+oGb1wUh19AS7uKVnuRVF1Mkh7R4HscfBngFNG/fbi3jf9uis0bY
Ffn7GKG9i03Te32jiwHJN9A4QU+3LiZ5k3+PPFF8wipGxGVPSEIcb/1jymIx7vzE
WJTK+mAAkwyMoepqZJn1SiFPHgkTwRW0YYelsnzTGZFXvk4G6TlTzHez3JtmpsMB
eFZVFYaIp1or/VDBdHYh2/z7XkWgyJJ9stX6kLQBQCegr2PZ/hDtWWc/kwjSFUwc
lIFpQX3n9KGvcsIGtDr5Sb1jtBvLRdYwNd5IuCVc5R8AbycCH1nGUCRcOkZRjhKh
+YuXXJzRKmaR9YuTEwQuj+giqSHvGiaYw0Re07WRzMSmxNwJnoR9LJqAgyWBH3UG
1XgE9gMcfDPzu++VnjZTFyuKkg4RlZM2E2pwBX8USmzuzdL3n+FDK65EcsPcRL4F
cr0oUbUoh+2T3ayR471ClKObsE9YleSB/JmQ9xNEvX64XfZuYy7RS8Lb/8mZGb2A
zE81N0qOQVjq2O/21KT3EWP7zEI2U1bIy+YKlbf0xZ/K9iQ6aeH3meSVf43Guv7b
70eZTQwMh1VviMDj8O5ixEOVnpxyDcXoJHH/KcfFMBtzP08qDSUblJrFBcnbsw14
CT9X8p/Tf9ExYbwmKNnhORoKxO8SGaNNKHhAuhuCHQuoa6B12Bhkl8vrviWclU+s
tfxNFHEZFc69NLRfp+7QA6/7wlX45ffrws8Qa/pb507msvrjGqPPHU2Ttxnuf47I
iI5Z5eqAGhk2MXa9iakcOxmVyd6brQZd/wpaPP9PNrWVn6jWtpct3gO1TxF8Hul5
rhjouHv3N7l9UHH97dRJYx1G1e2iO3D4GoQZhm7dk7fhmUhWUSI959xZhWT5YVys
swNUavk8ktg42NV+8KYhRPbqv2FUcK7dt59KTYQEcjTBUJiQqhYHM1GsbcqHNisX
6iqJ81hTfe/qqM+shslp0cTEhfDcZeM/Zm44c1x5mnh/vsyTMW89t9OJBIDBxDzO
57XzY90pBz3MFNpCEIr4+kf+UoN455yQZPNoIzeuLT2WzxFNfgGpkDmHdBno4dcW
vI4k/U3bk3qTvAGGfqh7yAE+AMPgfeDDAqQs+LmSyk2wiHhuyLvaBFSAh8Vf1p6+
oBONnhBrGPlr0iBvybVqSq4S1RGnhF1dD1LEkDZ618JVZOK5jffbOqHUaAK1XfE+
A5oRjWLkiB9D9RQf9kWXmHsTaDJ2aQTr3oY5CsGiQvzN7Y5p+73t4N3oZyv2XpO1
EFO5/PX+UTsJof4VG0HcD5siZef3IDgkZ0EaCv+7rcZeyMcABT/NkUEfxUqTBUEK
cieGXPyc4Eccdhy2iuYQT2KoNSqbp8ACksCqWysXrvMAq1ivAcDI8pI3ObfWS8fM
qa5oiiRb5um9ZH8TQSrgeReI31niSrqz7c2N5yLQfz315e1cik8uLr1GG2Ba0O6E
BZ2Hljh/iW2brbzdRVWtngWEtVv5ckotlevO9erj2ms6y+g9IBbBarrp9B4J8xxU
u5kA8owt0NjtMXeUfgJLWvDQIdk3ILO3LqPZjzmEeUxfxk2GS5DKH7wSMTSQisWl
priSwMVn46attKnHHvbdrEliGGWQNjMW4egt+EdkjdVH7b+Ivt8KO/HuwjxtM6JP
WD44kx7A4ZlwBqP5uTK27EGRPmRNecRRdLxIQNJTqMsHHiXN3QKuJhleMKzKisSH
NsVtEdalmgdpW6hJA/bEiQu3xusMxSE506a00IdwtHF6Z1guTJmY8/rtwvupYBTx
99ui9nU0znBq1NHldr5m4o/a7RRBJmVB9jhoVRFkkxzHkCgucvRMCfX/3vYnSTla
LM20KCSDvJI8+ikCjOLrRQUMzU/sKwJz/5km0eCX8+ErKUd3r2c+740L8Zy5HAf7
gz/B6RlipUpeXdFYRnqS0lLSWK6t3JWJlojYFLNxmDW0fCmqofeUebrbOCrZjch8
Xnh0HXgL6kOWze/sNjIxy5lnpFS5BFt5zl9Ay3znjW9re9WeE6BvKKoIGiEp0LrN
F0UJgPM5YbejI5dh6JP4ln45H3T546/OISyqBKRJqbgMJrhNOs1+MykCC7YTd+jV
kGXfwPlk4tP4JhW+KIX/g7OpqT+UgN6xz7dkUXg5YGMaBZhHfRYWYYHOOAT9wpW6
usH8KfxNJvILbwttE8fZAenUJ1Y0pqIfupdNQIvA726NKrGX6OOmxPy1rtzbYhJN
NW/dwdjx1xNQnfltDHVXgkFMXDvbljTsy+A7xjpqyPekDfkw0tJTWWtj986SECTC
tGPf+xoklafXiNArRLDcOskmqCLfPLBBPR/x6IfnaXXO4oNXe0ARS/o3IWzxi1TQ
smNpgogWKnAuLyPmoz0p3k5ErumGDkYMygD5MYI2kg3N1mQG4Q1EOUF4k1Ex2NTg
iZtLyd0fW+rtECpJthEQgohqK/W8Ehd3fly4cSfq/HOSwFS69MEbwWq/R3Eficql
IQbdvZnjWPv+eS+2alNYJX2gdiAGRNoiuUEbIs6xchCpIV6+bp82CBWyEmYp7t9w
WDlfoc3p1dDz3uKhn+buh7W5moRzA76ZGZsk1oTJKlxLIIp8nR+4iuzZkiH8PxfF
DdoERrC8mBcAMUSIdshfPjSnlnGeCkZiuQcxaRRBTh5Vt3ZbpPJvlnmgniPfEvy3
ZLumVwcOINwwCvqhN6PpOHDi7UdI3PNAGr6dxCz6P5IlRO4cYQzZWG33RGHsybq3
lnY8Us7CLKMhTd7MMHY55XGOUyBq82MJSd9Dh/p4vv4XojsatJSEBIUHb3SFk3+g
GyOMJ1YW+2si+QU5NyLS0PdZ9jaDc5ZaW6Z+ONfVCjx4zUXY+QzHXuon3RMgI1yb
JeNvtypQDjj7TgEPfVh0JeJYQypBbGLUhYCRSB+k/5qdapMOLydMdzdHaOUgEf9O
vK6pHESAY//4n4x8wHG78DxJRIgMPI+Ntwc88ODENO4/ykkuIoXvyz1VN/qZzksA
aHuvK8/xNLM4lWXIgPRDnCwPISuNIclo/C3J9L2XSyWeBWyppxIYncmhhbnDtBTK
Juis7yD9PGprJ/YTrrVLVwn+dT9g5Fe3GHI3B2pIJjmkwFAfv5e2XUTouPCzg8Pu
T7j01LyMIWx+PrGbN9ikTt1LMyR3IcjQFqfkN7fBmJf+3d8g7J3KBo/IG6O3F03z
0CEh8Tx2opD9VdsapLvdbagmMIyC4DzPy5aouuPLMn0DnxQ7+w4UfM5E+jJtpAvk
uIir+d1bFp4M9dmqM5qTPCPWZrJQXW/m7TKHJMXjF7/Cu/yDSrV7Jy4UQTi7IMGD
TXvKm/Rd4HSOUFK2DxDF1a/bbNU7X2tHBeYUCrjkBAWTlFif1TulsrhJAgLF0tbc
epaP+JcR5wWOc9gRW8mM/+MbH2L7QHR+V+yUOzdMsIr0cR8iRPmhdcsUS1G4QFv9
umx2yo2qBH4s7zx3W/Ly+7IXDYwv91J2cvHqvJbXSIYI6jgzbVMIGDJpWzePG5QZ
gTRfpVkkcLx7YnSPK6ao24hOrSQIHjjFjWhgU6bKG9wzVbTVL6OR8/leHbnHROTq
rFo0MxZ62uEwVkiDZz5s8mrnhlUFSqg0TEelFZuhJ1Xh7h4vG24n27bkFcNWhJBE
VcOyuIvXybPugDweNvs/1vw3xvzA2OIcQX44uz8YHyLkFhHX3M4a23HZB5XCZyLB
baq/aSi/CBpiC7etxvdB+q/7JnfGPH2q51MCGmSu//VkJQ4I8p/7LjtoqUXTFPGw
yQfn2qUQDme4Aekh/2dlLROvJfM95E4XqevS8wY6yEj6gKK5GvBAGtILlCmAbdef
YWLwfU1EwGFNVuRqIfqYLIRcUJMeoHr9U7+5o/oUODoo6208YZ0o56yc+HIWZE+B
2243nkj3gZybowVHAnPA1X6GCdn/OxgRtzZd+No4UQPHQFGarY4q8ScTMt93Znio
oVrQgEzKWKhEnPzH97jTlJagQYv37EZu8xQngugmzsv++kg7DUlmsMdUac9AnSig
NcPfSQHq/9lWuu12QnElEKoaVBp445LdOrxD04qAg8SwyT0rk07WOveC65mNP7vA
9j0GFTzwnNexyzchRM3dRMNmiJH/+7GkpO1rCQfKKWta2eis6mfDxVgGqvFItABz
ry1Oph1VioorFg9hlkJdHQTvInW/jy5PjbZwA9JZbYNvL1b9l3tInchrypsYhN1v
zOXOW0MiuzhO2AQNPi83BFvvdW7PGEnq4MeCjDLz+vfRco/glfl/ZoOATa+vW5Fh
dgiW7nkqA7Rx0jnhct5JriAmlSWZnRb79Z7lN6qA5KnP2vdVvLaZKynkiaqneFnS
BrXqlYJSIMoRNXCRyqvKtx9i+US5uDUSgavk+D1b6T/7qAcc+xBI034pVEJf5tTf
0meK9ra+rqRmOUqlZP3DL//xwwgUr0KKOWtx9wQQgGZQPXvKsE8KHgDfK2IkP8ZZ
tHTBuJwJnS9hbzmNlg312vGd8OUdSAQNzZ0J5dMuo5tVurSrcPNXEvjE5AXMPz2r
RI9V+8enz3WDUNy1K8BBz+nGE/PsKWvzh3FQUoTIB1KmhgFcmlcJVj2PeroCrwlQ
jVDshKw/BPmQFwGYBB5LUkbyXMyjAAzbKdf0RGeGvRG6XlAVhOofjWDpnXBufqb/
3ROSwOf0x3jVxpe1MdjAMgiW646XnPnDal3cG8ezcpx7cp3aa+MemJY5OGxdu96O
8E9iJXLVsYDJMo6L/eolcOiRzwtx+XQ7yaQNQ6BcHtgl4dA23KczfygmjR1E+Z4M
N1ABbB5Ogw+lyWQtVR89cc9nWMx5GEIrFAhgJQC050Jy9ATV3th79YafYpt8g7uM
hrO60yuo+XwLLPekHiEKivfj7yJS4syEsOSuoSzZ+2kR69dSRADpVdFJuWX7cl1X
vPak+lsT8zB5GRnGTLm/xRqBVht+McLMpKV5m8sWePd1f68xE36WdOFjb28WzmV6
LDP+7ZdTBgasCnC9dv+BYLQ41n3fH2y1jccpaHT5ET3CSNvLuLA7HAPm7YbwCBNw
2vcIu69hV56XJT94IOQgZvtDNVxpgbj7EgH16TQRGdHWuBwJlfJsXyFwcH49ACPW
UCJm+ehcflZIbUWKZs5MfYK8TbMBm+x5A2Xf0g43qDIXliDjRGiZL91413m3IY2W
WPuSD8qDgq7O/2gVFKhDI1UzLtI4AkrSed7pJLzE+hU2pKqwduXSGA590E2lI9qx
cUb3wd/WhUkEwtXhKgn8cRAvTZ1tbXQMjc/HVN6GqW2MRgtzNbLDg4P5IFm8jgBC
lFhRmVpO4RK1mWjS+wYqF7qR9uxhE6YOcfheW5Dx1HbGyyYejjIpqbbVfsFgiSnW
IjuKSu9KvFY4f1gUiipdnOf9vBtSmaCSU+kzyJ1SiaABQnzJTF92U9Y2vbFziO8T
dl4nSbbZwLhfJ27hcBUqIKPYDanm2dOpbA5GUhBtL1ntJj0dLF067hW5L2hIZE3R
M1PP6mjUQCD/cGRf7irdKe/D9itVZs4D3ZZBlgogBKEN1Dlgj6zCJsQIy9DPz0d4
OMO2EBmrrHJsjlhgm9YKR/wVO6gU7Q+f8V2GyED6r4/YoKrfL11GhhuIk5Jo2PrA
EYE8g19jd/eFoKDJQTOoAeCsw+0ORWF2zKI4jJ+lvI0zNQdkiLQmhxgiIZorKjqM
Dl/9cYJ71XGNeF0FHK/NCeZ0mVohjcpdN/4jgnJ2aukK6zgU9nxe0/jpOsilQDc2
wExWzFUiO4VN2iR3gPGLjhsMu5VJh2RTP1RDhyd4E4J544YhTOtDlHCy4uVrdRqi
tGadNICEbfTDeiptqJnocXmmZR3WA62wp1L40/RQWUoU6npn2GUzf2iLrEPOS7ge
RNijGWVeeVm8Yo01mGsKU21SPHnihsOQC67WaBS9NPlQqPRdPG51OM3mTsu/iyyV
3VS+aVG4jcXrjpOpkL3WSRHSWHgdwRDblt8n/eX/K1PNK+6UsogzXbCCEY4BpLQn
U8p07rUcCAfcVKHT6JLvF4ajxOMBnJaPK1uTKugTw1ETJwif2hQ0hw9x5hDFcaZ9
ssAURejAhibKq45HvsZYfsrXK88OFgcTX83YSrvLmYcfrdzoR7p68MR4Acg5Kei4
M99nw+WQVr1rHdaYNm1LMZ+8sUmtjrJ4HbhTd5Hj7wQ42+uVCQLpnfZQaOw797y8
VH+/J7IQPrqNvovpchrVHyxl3F+qxdHrqk0FCxmJlhzqwdPzERfqb4Jq3wzbNW7p
SFHpF8VNuVEfqikxpjvDg6m+QdkTc9/TvRJ/A1KF+jUhNVXIf92MR1HLFkH/y9gt
dWvGlQ3lh8dRly/KxT0hS3w1Ydy3yRYRMmtefPOQve/mi3uxluZPs729mHyZhBe6
Bgi3YG0EK+1dwI4kFLaPde4bl1Z3zItN0KIgL8/3wKwWi8aU2SuAHDYCPtZKHaZU
FuXTzVLQDkmD94gScJFPCvg6vRjqvC47zyAweJiWWwM7WqpQM3TeU0+kaAH0nqr6
08DcZqvP0cXYRB69nklv1mHz9BOeP2MEKBUycUw+15BPeUdllEvj2pOnTMAY3ncT
G/wgT8yay9Zz+V3Ac+QshpQ64sXmTgCRzJ4RRGcb3PyuPZkDEptSBKxqnqtOo2e6
xI2PswR28LilPnfkJs+QmBOIVsDX31YHricLIQQlwB37I3N2LVRCkutps1LRygMv
xpFxC/OnjJt1HaT4Jf6VxN8wD6m7agNdtdyxnAqS65oQv91IK6+AbQk3DZWPXlUr
CSRwJ5rx0+g7vCob6gZ1d5A9y224BMsUFROeNpTZLZaFoqZcjkRLGA5tudCotzxL
tjD0DsfI5oIgJ3ATGFoxk0z32XQX8rHa0wXEn8f6ZMqhFLYTTjnz7pAjXrLfUERA
4fRY3cqvSxOmTt6/7Glw153bvvr8NxD94aoNvN91G0SQhaouV6+2nZGaPHUWImKZ
J1yiVLea1956GRjxCZgpgHsVRwVAtTw1yrxkfs4uNiKDHUJiNR6MR4sCK6hMH6D7
r+XEOKhIxYvFqYZLSnKQMrkQUKmDg3v8XLJDFxdGJww=
`pragma protect end_protected
