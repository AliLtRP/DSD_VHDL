// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
WWjjcjM2CVTBDxTEk5Ac/uNXv2ecQABtlgbKW+IL5mkf57okZnEJTAUCplYb8fw8xxt5ffLyT6Yw
RQk8P9MsDCo8HrCGC0v+Unee65dU6Gy4x/EyrwQYsiX0dsbkHz9jOVC4l6N6X4ArRCX2M7D5e3vX
gh7uGDdJ4e+f4nFlEP4bCiND0vFyshKxIccX7X8O0RlxxpoRl1IXVm9WeE7xRKUFd8bI5K+zBi5u
SiWSmdOY5RWgBDv8ppwcyUzYp9DJS/2ZT21rNOuiP+JaVXk1/SujvR0q2+uKDgjWGYfd6UZL+m2y
feHQK/utKeS5ghbWu0utsq4A8on0YQcmintOHQ==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
cHmIfMa+2LUd+Q4NvgVq/PEuTrbrqcza6S8zAww22SqSMOcbzzDc0WlrdOyOdXye3FL9bIs7lSFT
7yAYLXim0g1l4NuS6rtIp8K2zZqeC3gYdjgQmRVaFIbGUKfZd/pAOFYmZ0qyl+6oCRmUjv9wLCWw
lg89rz8+UMVABFpC1kBhYEdD6gZu7GTaY960KZJwNU29yc6/VNyF0NbThmATCpqwCjkCNELsS8wG
f7IvXZuQ1uDE6hRbVNdH3H99BF2HUNUHIvbGT227uk0ZlgqozTjvsWTKdAi3wydpiQs8vSUZKTmH
Q4o4LgHS9apRJw/y9atcu6/xz3TrqH6XFIUjFCzFwOeGIOSphxaNsI4T2hiyyfkI2zV20D2eTMR3
IuNmrF5bycZf3RQEo0q+8kgvO4CfwKIfIPpw1vJROHEzgGOIb6pX+/1r5W1dxB6qS/fWg0ybAR0M
QL7CvryHtibUbZbCX3NzrDFjBASXH034Nrqao0UT0fRK6ePiAA+kR4HeEYUzgjEvvNqLcy/iRA1J
I3pCzUQ3rCLvdCknusn6ToP+9jusnbxg3F0YMdWotiqnBUowj2h01TLT7VU9x5FRGoUjEm56gTMX
qiZXsCuYyHkK+YFAysJTHXu6c2CSkFbOFb9h8o3/pS4UPFBfVR4z3sKjnAgWHDY9Je3qz39G7hOr
vTdw9SQuq2vNNOSVF9KZbRXKdF99upl/Op9OIPW8kEyRomFEoDoQonTrv+heggH9c6cdpBOJlEnT
GW9frbb5qeJDgFLX+0KzR5uoYQa8yCjq1s4AHP60JkR4/UpBi5WlvGjIX+QAui7p6rfZRJT7YkAg
WlkJaUKiEq5rriOuvgQ+zNnNpXD/uY0hXMT1JHbhOTG7Dr6y1O7aeq/D2A1exZfk0ZIRD6+MkOEW
vZ8MuXn7+B1ydSWP6Bw2R5KRVfeV6FMF5Q0wASqu1YDq37m4coVeAcIrjZFSy3vq0J8xQtKTUXcx
1LQCZUjV7DdKc9PX4I+lgkq62MXL5kXIwlMIacMu46vSDEfbH8rjHT+zfR9CZuC1ACNQgj0zx8R5
rEXnqSsiFMMWc61818s5VMfQunNbIoppFY+txo0XNb5EBpg14R4+ArtZAYBHbJeTMuWRr/lRvfK2
MSWsocUE/xOcvR5LGWSUeV+fhBPtQB4/Ulwrg8PoL2wTMQPgS514d/fxS0q7OQPhD4W7q6JdBFsO
buOiyi7vNT8dyAMxXIht/T/9gsUHtSQPwmLnmz6yd/DKoeag9xLoAEUEb+wF3nriAWngcSrV6F7p
cLBGtKYUzTzQ/f8DpTT+Hc8+EauDYkpn0KeVmTSdPWewhB+n4ccFfRDdc18oKy8iWTM2I3Aojkr2
iV0ZcAyLE6HUM/t+ls72THSuL90BkaCuHikwlqkHxazu6l3xFpBZuncl4EDlWTcqeorO4c3yjtmp
/VCc0WXJb4+7yHNRFZmENraK7G1OUYIxfpitzMtb2QYDOkfZHAKle+oWV5/7mzuL1OKQIauao93F
kcatn/N0DitPaWTfX9aBrig0RoNnyxxjumP/9Ek+4R+MX4KH9vZHhzFF1sarho6cbjxNsBbz10Kd
6ETInE2uScdPKFuI9n0CJih9XDFPY1WLZ/mvy15YV66XpI2f6GX9R9TBRyvGK7mjiM1MqLQJv/ui
OvZqObm8xEZOKHLX+YbBdcZuI/5kWQQICt3uCDE85jOjht940jyST00JtMlQrozwul3MnPeeb62R
rsxLB5MWe48M+Yq6Rr0TO2/d6Uxa378WGIrlo8r0SD6czN3UXnMSjspKvAS+dcw2rLsXCkkyI23Y
RXxwJ0y8BdUsOYqligryoBrqHm8xmCD8ipDen2jPMD4pUy+AX4KtI8F+MHGpZeVEATBUe5D6MUv0
/XX2S5socRF49UO+tMjWqM/4L0P1CPFBKNAnD1sxte2G0TOCtqpsFQIqjofYoCp4n4iG6mtPh9yS
Oy9UUNuQFa4jYZFqEz4NihwDdyxXC1WUTBCfqSN2R62t8Zw5eSwnNrKpzE/bh4f1ycryb7ILq5u4
2w2j8wYN7To4j2+cRIQA9m8+yzOUqIoArlXYLJVbMyMvk4AqiVTPSAGaydksVmldMO2uyjB/T6yH
Eqz7JtkMYH3M2xiaXS+wZrOSAHfGzJsLOkMMipa8jjVn1GqaBiGhOwbatc53cgTm72H7gTMca5zf
D8g00izsl1QbemiPyrsXbwoHr0gMzjJGHsQKYhJ7jARd4ZE0+CAbygwQxqdD1U0T0f9l9hzWiSTx
QVTfsH+FgAZSZLVCo+hQ0UN/BLuT9AFNWBYL2J4llRVs0Qen9RAGgCrvQVWEcrOmxDGEf1XY3rf2
AAKppV/mfv4i1e7EXssPaTvHlAwr9zj29mWhO8B/5wpFTPE+uIPUn2citKyKI8Y46URObSqOEwO3
xLKfZ1oUkcIifVXvGAg6ZQvaKH6x2d7Tx+Hx0KDORZ552+i8XeGL8JYfOYOaonjEezwxDwMz4T5B
P6CemjwZgR56R9LRMCpajsIBPgLNKZF5dkNiMdr0hhvkCvIZTGWZJ+fn6ZLiySsM+HAA5jbQRP5k
ALavTV++kI2UiJOg9nxL+QWdLTSMCPi3m6QnhifBnoEKL7P+chbW14kwfjgaTdyzo8IGwccZEr1j
4Wdqtj6+Sgzaxca3agTUxbnImEzNsdOnPmzPPlXD/494chaKMACJl6gyMtEV81CAXvXhgkHBRcRS
si2YeBFo+kXnDp0n1kSNLauDQSBBLlgyU3SrnWbThPLVjImvWHgI5B6NnH5cwWCuQ/iR2GWp+XbM
68Nx7LmbFrWh/avZVy1D9URYoC38YNQvmETjO2en5rpRKSTrE1gjO+15EEKU3WPWKNsArdNg7Xtf
qUSAPNhAgyTSlln1Jmjz6WRFqbzSSCWXF2qy1CvV1ZHqVzC8vwZMt/zsy5BVY2dyGqaQ8tmf9KQp
eU/VvOiqNoChXVPR7SV/vshDyElV9ZYexJjaE0UN4RK1kAfd6pGYzPws26fVKwyTlNweyataRB7z
XCjSLvD4lJvBag6beIH7khNf9ITGQA/+yBBNkdbiFxPdo9rYCOYv69uZPoSNq2QvajP5tcFdSpnY
MDG67VRL5FN1m/XSxC9xCEByXbjKKBaCDe1EcFnSUWFMc0mMTpBX3RkrU2PPUeuP2A5SwlA2w7vR
DZHYrYDpfLk+hG+3bfaUfozHlPbhaY8dSR8Nq0S8AKHRMwtwTiDMCIOoeseB+jrqA/VRTa4iD5Oi
/3CC0HgKMF7wZ67fSzx/bKkdRfwSJSQo96r1sstW2REyCq2SG2befaZ/NQa3Rop//CrOVWRh6QNi
P6r2i/CBMxl2PTK6GxR+IvmB16nZ9nw6YwmgfyJZgyF9BLbjWGBPzl3t5aWdCSFvnecM7CWUpDJT
EMKBMkjIWiyTIVsZ8mfbzSkhY7Q+ArWxNiShChAqE4ctEsg0hWlX3GArqOjp2H6OPqZ7WJIsnLWD
vMJwYWNumFw1wlY7v2EDmeQjiBhA5Ojgs7kkY6Wj8He8+9rnRUmW+RI30mSQuf7w9VAI6LpTL1El
GzlbmpQw3XoOj6BRP5sQMvxBeZ0P5q9iQXQMoq9c2lj0XEv0YkpbwFRgR2ly7CCOVx3+WukCju0x
ybtzq5Eghg4Xp/T2J2+Zft4FO6LlGfqenPXoXCL1MtCBPFXUJPvy5QV3h/QgFshfP3Kd/MkbJoTG
WM6i1QouJhjDavKqJUfacy+ueMQjAKDvWy4SJGQcKiYKDmCV5t2e2m6OHwyLrTz+C57fNDYqZDJK
fY56DL8w6yIsp1a9ZpPrpvHKy6BUtEb0t0oIr27uN3NoraBvYD+MnuSlAjtlXn1CZejstsIePl4r
Gb9kIdltj0kRcA86q4ybjuAaP1DIR+T4aSRdbkdaKwCCVXNg6mT1EEdppHWG1yhW8crM4HiR0usq
IeD4tKuIcgXz4eJ6IpgeafQqrHvwEy+84DPGtOmPfYNjUqt+UVQNK381ahu7sP1m0oNeNFjwsXfc
yHMay3xKx6uFirEehFD8VTub1Vzp1StcTyZIkQAkc80KyDgUV0XLD8NwQrqgnagiVNiSV4yYmHbQ
Mn8cpgerSrpWuv95jGPpYH7/sbmeCiYQA3VDv6OLRKJKZBIsGsM27jqLrDtWl0oEfYL1C1uGEhdf
sp/dFJ945sYzrLTc1b2eo33CtcGFlnYHAWzOCQzFt9pgf/Du1efpZ1nufKFxyE61w1yCPKKHy2AV
XPOasQNTnV6ZTLqWdOXi0s6n2l66DD3eHPKzORC7k9XhUHUuTIAUT7Kur93yPZhNStFr4sB9Y3z+
EJO6Ok8g85JdMpi46U8CEfKb5s97JP0TCGnCgwCE2Hlc0610NLhbwNu8J5yACLgU1tgv5xgha5CU
5aZaYiiNaChwaBkA0/eFDlUICoQ+YzmFcY5LJK+HPJAMb/hJJSzicysXWS4AdXlpxFOB3hSJWv7D
KqE/o5lJh9zOFbYlqwBJ7X2W6Gx7WGfixdvq11wqzdUqV/XU0oy+8idWaPXeP0DoEsAbvebj8t8s
l1qFRrq+XYZGAoNnSfUm1P9xwbEGHsTAIfEPHb+ChNgmzqGcYvWn7Gf5a2a64DnCEburPT3hRe8R
igZrCaewTa7B/pF7LCVjTChMu6qOtMTickHnCDT76I+ygXHBuTLIZDQ//tUUGS08ejtvBA9bcbb4
cWOFC90geY+NahUDECXmiYXn9nmG8EH0eJyOnCRs6UlySPj7blofBMtJ4f8fWUN0j+ypjKez/0rY
4lhSzv95cKGi9vuihPq4Nv0kn5OJLY8xTFLL4WrNQbP6RX68xYbBzmqLUfeON9dNgB+lNK777hk1
YN2fCILr/O+IpRJlvKGiSdBEw68epXw69aj3vMvN4xb3RRV7Oqyy0CYzy/L5dsnhW3M6uYDgKFZX
ZwrwZ4dSqISn8q5AvrjEzPJS5XXT1I1UG/S3Ii7+s90H7BqBvOc7O2LODFkg2w6iVuu1KXjMYHyQ
KLxMle9Tf2FVyPBLKAf4hbj1F++Ewb6fUJo/C7SEKqd2h8afRlx80iFZjDa8ZitX3rycZushDiAC
FpYNkkr+n1OjQpYFmdOjDY+a0YSmjhX/xlplAImG4MBH1GdjuVI/oIYqv5Mn8gULk4oIWWeipBzm
pxglUwPW6RZUSX0yto6WyKCJjhSyn0cWMQXN4UT0Se/lEvNyVaWdSxEgPtiMOhI5YeCzqnDciwQu
CTR0Tr8lxWVV2QhGgSzKME/gp1PfvnvyisgMUVZqtTIN2D9TJ+maYgOxHujyGBsz364eDlfMYEui
fkN1BgA8cyCeupafA3BkaTNDDWTeJByWgB3ETGdfURNbvL3vByguhm+sjgCPz3eAoRn3Nbm/SB1n
q7ulodZKcAYIbzCIgyxRWaExHt4YAZl2YD8maqq1hmyP8lEi5CUZ+enKuvalJhZvxtQ7Ogg4R3DC
dfWmLJs6niJy9rdjG8FSqF8MRSJi2phj4IyOmKClQr2Q2kCeMa6FzNzHp4BbRL/1yi+ky4zVDR3d
QahrygjvE34Fm090qPYrtwp37pIqzTpkRKcbI+Z1yMviixtInn8GpxoqxCbc6OoJR8LnLM0bT4WB
lmpQFPDV2ewtW7o9mc/folsGXtrrdVB0k3oDMXeEgB+6koaUzMnd13G6GZlhleXTH/pN8fLK1QAf
6HvdzGxvEhOHO9jfRv0qWiAjvZpZgeNGwBXGij6DDi91QAvuWIHLDROuYgXk2GHojQtGFcBmMvVv
nRxFIEm9+4OwXh0zVzTdDwKGGcW4eUmbYbmQtcSl0jCNDJZ6I/3OUjBwp6L9aqwdhbzBDEhKGjyj
B4mvpc2zhzhGXRPNL8YTAnM+YTNQRGZsfHuCKZDBoVYm+0L00pUoVbdHwfIzp+qBo4K3e4I3V0uB
wpQRubWSWhWjhUADfygGnyL+K6E0ttaMVbWpiWpZnvpA99cSfhQ3QGdtu9cRUr5YUjWaDAMVQZpc
q0gNvyA75UwVy/3VOfPFMFk6VpKskE/JmTIYXX61Bzk5Dp+2+1W3d5dX7ouP1q/NhqhhNpydEa7a
2eMOSzo92nKP4BNnVUo3tPNR8htKZFBQw0b6U33ozVzL6L7svrE6TL3DXplDoDEMMaeKBtZMfQxt
MnDb1TilEiHmrmXNO3dXWxUqi9fGpiOzXMbm7PeAt3wSHQ3N1mx2/s7didDZs78s0cs47lZueCv+
7Ty5Pd2qWMbtjiOYuqUA2ov6ypopBysLW4lR9mocx95cUeGBq/lpp1iFPOOSBS6Y1yLkHKMd45xI
Z9lPG6sNBJ3fgbE6Y/NGVHB5yBdV5LgTi/qkA4RWi+xKQy2Do8+cIs/DfSpnW70oBGHP5E9BH1ks
PLodvUXvqkn2LZ6bXiyTMJoKLn/Sl9m09vdo9EOlSNU8uQAb6vN1wD/sWFzCFvWqYmRI+yWAziQR
u50albaI2fgPFgUplYktS22uNA478tZvo2/aydhB0ELhRxlou132GbFMLO5GD6AafyP+7Qg9B9rg
yJaI75wr2dZJ3btTVkBPJvoOvzjw+Fp96r5FtRJzkWJKzPkeVkSlIqjqOaDkE8gQE1heTaa6dW/w
x+ER5clOvHMhyNpLVDdd35lYI9wwpzOXOfw3oufNCY2FeFs7X3/4BEmpxgDQlsx9udxauOlH9DHz
Ed4aAsg4iY0+O4hkeiSRnuKgf830dEfGS1KpnQIMZ1+rIRIPkXmQprXjHfUTnF8kkdPuvFwZ+h2Q
AdkPoHUr80Yb8htGyKMGSNpf/HjOEfkJxguC1sqq5+hPG5q5YXmxyUeixxWm0z9DCL+dgApKMC79
TqKlcsKdFHkqBDghdub4heS5YKti5tCwE3L7LVYuBIZpqT0H4BZPqg+5IESz9B3v3MYxIOyW5gsT
ggbLoM69IHdtf2jHlrzDqkjWj9jNJLF/6a5cPW8OtqA9yVdxMM0+Mg6+N1IQkD330VsUqLw6FsYd
PfPtrlo+vFDJmDi50SZIrISZTSbFlveTpPF1qUIVQ/4G9LJ2i8BnZKuNdRpy7/oChGtRnUA+LxQj
KBqCCNybvcjCMULglJyvkkpVbnotJ6RCWr20XdLoZAWR9YgHz88AiwGfR6r29sV9TJVK+F3J/uC3
31h+heboGFuPayQUY1AI6B/0tBwWrhzm15d430w5w6itW5cP3J8w08WXoZnvHrkRMCBCl/9RSA+z
6XKcaKWqGztGbGRLjlmGw+eSQXM5b8SQa7pThOrpQn4efKP9yKS7BId1S+NiOHo/RXGoi6M7AsWk
5yTU7RfSwcyUFH4L2YFxJNz4lg0IDNwmVetT9Nu3crW9NgDqmHGy2ytANsGOGdsvUmLhaoMMSX2s
6B5PQsTXVn0AL4Ct24jwFIY3DtJXK3sJzhixgCGhX3f8E/v0odSm7u+EhziXWybvw2EFOrNLndRo
R7JGKKrwu5RMbIxnuINNtuCdJCEAtr6k7PadFIAs5NCSSLd+tEjN6XCef6OcGUrnR73qstG36OOI
fDGwUX42USVWkoRQJfSNS0mh7pDGx2z6Og0fDg2qU2CWfcaitmAnEeK5VsCspw0/3RbtWMC4Xo0f
8YFb99Uw5URk3Ex6zlUfaMdUu/RxoRVIJpRuDKOxeyGfKJCYw2cOkNkbLhoIcdyMyKrS9qx/ij/1
pvFUtvktOVAxj4hwwbbz+rFj/rHb5fqMajCJEzGvpvTEhRb9DhH6JPVmLW56eHAuGInM3xYFp6D2
N18AysunQA19pXbcnmQa9/mDZWwF19xLIKOcRSoVRHE488D5TEWUOxwoxbMxDcm2EyDy647hWiQe
3qXprXZS1Lomggbb+1LX/ZlZkYMx3TmWhfSYOrs584OhmGMUcCpmewPpok7L5txf7i6WwO50+yh9
oHgCH5xBheFo9Af5UVCQ4cdUR6YEkLoNPrAcHDRBchvvO+hKdi3mIq+0w9WnqhMT0PenLFjO5eXL
LMuqFRTeP69K0DHCn8VWtxer8yWW/WgvUgGfMTIe8me7cdrVm94VuYmpsASvTccKr1L8g31iM0z9
+FAc+z2CxxKPrVH+3qcgl/0r+lICtiuByuJu9GjAND+flsjLlmVNzoTQ0LRFMz8LcDHa68VDKQqm
AAeec0T2AZY6CSk2DolcEhhQtSHTO0XBm5equluEG83d0QaGDF/2doEn42yqIt9UDXustNUxnBCk
wPdWH8ylZDRFriUs1kklH7HG5N43nh7ZUpioo0cZDmvnma5UrD0LfPlF8SyQIzsf/O8mNJjnIMTO
dG198A+8+SbWH2RL6Hsh+u2Opo3FT8Kx0yzevAED1V1qmusyLLnLCq+s49StY6wDAfhzJtGmtl08
SFyclXafJAtAdMmVWe628rA+xjkk+yAISUEgMywJjgfl80MyurKsXKbFFdDi7GjPMqOa2iz58jYO
zmI9Ln9HTg5uYaC8+OLSLkibTF79m+eq9R1xMS94xRK30szQNt5cCRNlJStKSMIlvoSVzKuI9P1u
t1YYJAPFt5MMN/K3WWGmNLA0mpoaIwf3mEfnLNxz/ojl1nfSOf4YKvolZ5lW9+9ma1a6gLs8Yqc/
ut6xqtfo1SW/QeYZ4aKnM8eYi1EodmGG8/8jAqAQtB1eUoX5XfAIjosu6Wyq3Ki0VLJLRQde+z3P
+ov804U7Xn7zLEjduqpFKdOfaHYafcvJ1E9qkJQoe/LmjeEjHtFyuMPekhwP+SN7cPmhdOYjNXhL
jhwUEKfGUJVfPE6bbwvsYipELNsihyhVucXrogvACdHoJg5mIlNSSsI1UrrC1DspXKTQw3fguL2x
emGxN6uOepkyX6fRan/apQ8qu+PI48YTgla2SDNobM9YwGNuP0OPxKXrDgiJRgaz2RoW3HSuCiK4
fxt7+Ipog9CgkRc1JlAMjJeCmpvKf7upVKKvKQkO88Szq/XEkk1GTA78dD5GWM9nsa2bdaVtnAqT
ZV9Z4u8Y7mRydk1lKXtpTWLElewcLwJD3kFsqjYgmcUFM0jz/fcLql81tLqAjrpHlR1dNlLUp5/E
FyS6uIkEdLLkr4s2iu3KZgwa+HKqhdd4awGe+pWsRdFHwyh/XJbRXArkHTLrnl9iIOp4C4bgssA/
j+BA5sfiBC8pKVmf4qiRrxKCDNpUdLrgCtLhncmBXZLnhqXC71BCHGghxhGmp3RPnnfXqWWT/jC3
wXrapO3LQrS+5JLryhfAtU96+IcykWUKUop3wfLywfo2ts2JE32Rz4JyUbDDeYPPdDXwFWQKD3mS
fiU2X2AmrLgsi0GZedy0i8KmOudgzA3qnbx5gL5+ZqQuloh8cbPUOzkRuEUeLAoA7TzES4mSgBMA
dTxsQZE4y0/oFcrl5+LcWxuOYyxK+q5Rpg0PCw8uu94o6cg0okF824mq2cigAYeNP+y/zx/r8SXo
mOa998rPyr5oWoI6yub1CX0haWKBAn6tcpl5tNlRa96B4JSiOT2MJH9BdNXIj/i1H0m8agnYgiMA
BuSalzDs+eHS6e3HrcYHkPPo26BkdZDcGiXo+MS1QLlzDTkpnROgINn6R5V3DRLbtNJgWD7jHgqt
yVki1c4mZrPvKh7iRk3/HBkQXs3pNpkraiuOVzXB/wM6aa/DuJ3+bvWHGL0dVr3lkYV/pC1FJipm
vdeGG7Qwvuu2HzALzmVD+ao0sSuXhJB24A6XPqJizKo+fqf2qBUKrfyyn8CWmPkp/vOTNvj+KXxJ
CtlUFBH6OLjKihnjajorEFKy/shzcChzdYu/mEvfIlBLFUEI+fT2/j3irzwueSTQ26G44MNkUUdt
Vc+LwWjVY//razX33O+idMkWtxWPhaTOivto7AuupnQ72DKfawrVCaKoY13fSzF8XseANSUTClQu
QrRxzCvvotzK7gHZqXEVyO+an5YeCfwtBG4DK9vhpWcFw+FRrbNw1RwVZgmNAth3Ee1nZQl9eoP/
ymmWla0dXF/RAJHx/zZ4UzlfqDVsrerqXlEhxXjqryrxVa8d7LdEBVRr8Nfo3tquCFQSNptKOina
JVwRBKysALFE/L2ddgApTmm/D/Pj7uVA+tlvQNeO0XK3I7tsoukM9ABC1DIaYtjJmyXjqInrQg2+
0g1Jjt4xaqX6W9lcZTSVhP0dN8x1KUyHSmFogxhp6+8usiEMutbuiF0J9siel6Upb0xk4rtx7OA3
wbYwslPXqiYlXMqW8q6LrqGiqiPlqLholnn6EKzQHYqXh4NDw563CQlhHgY5LYBe1ARQWviatb0Z
+0sSTKG/TkvnFm8/olJaIMa1oWCBpLTKywTd3IKDi7ur/a/XbiAT1PMRdRjtv7dOH9kHrzOn2och
lFdogox8gcGP0UTw0T6WQBjkygSS3xQsjkdUv9x6H7aRQJNcbiagEL2TmOHZGgUa1m3jI02WGZtG
avJiA71jokUAiwMasAtlaJBxv/q70rjEV9+W4cp6ump1cRJvIUS202oL0JXFqHpLEwRkFSXYQ8pj
gFAuMOHkvQxMK2tnj4CH0adVUluAIS1qMg3hR+udVBAlG2g2VrfA6MXJCxyffjW2/yRAK1X5zJk8
mF7fggC8icDgtlYTzNQRrDZZk6j0eYm9hLWItK7VhPi/0ssIzjbqgclJNDqKjg/Xc3Y0Nrias+Lg
UvOrKLb9v+sCVyjtd6m65GnvtvnhDnIWTNo3dWv/t9BTioel1eJ4Vc7K+1xq5OPXIGOQFaVX4m7Q
4ULta/aVyAqypAHdxssTLoUj/L+E1ZsFYnXzJtEdPaQ/2spAO6Av1z9955qX3K/G1cLY9g+sB2I7
+9xxUn0w7V82TT8RIKnHf4auTGAUvtVlhMuROrdVbSDjtAyvpbqug/4FlcoGeHaRV56oMj41XJVq
hskmZC9wiLLo7JpDZltKj5OxkSs7XKN5M3PKLXxglHN7UkMbR99VmJBHHu3hxGufoR9hUUulDnXW
EYhUgQq0OA/M5f8y5gHlMr+o64HWhh1+CeFVv+b6nVNbhl08OEZNPYq4+F/hnpgTEGWgjn1VkQxb
+E/xzwSTFlGhPFcJqKnZdEZE7uU4/I60U5WXVPEava7lrR7uo6z0P7fQuQzxz1dlySpI9n+cRiW4
2tgcFKtpkf0N+SL9e0qyOG3yxXbsTb+DWF+ZOsW8U6aloz10tbgxdt3L+Y4TCcsi3380eZcbk3pW
krQ5sguZeJUSOQrg8HSISN7R9rgpIQPX0dCyxnnQwcvPfaa8oplIKFjlZWCSC3HCmbBEET8PrA3b
Mhlq0cGWmHwT60t6vIwqGu2av0Do/qP71db5o9pw3EFennnFjdiafgjWU5bM/bX0hNGZltnz8jz9
XqhuHPJN+DedczoqDxspTfQIOjoICAjedXI9Jqt3jQYWNceQHTCRIvoUhB8/VSJSYbt1G76zbX1h
gVBaSpeCOTseXK8bqvCheL3BKLiR4LLMCYFbWNp0/PGufZls/Tl4+gmPLmZKno9K66e1CpK16i5y
NB4tsbPUqgbWJEWJQMe5stSbJ8srd5jevcRJ0UYH/gS7jBFVUQL850rHkuqUHbxro6c5FO+qQVR6
onfWVSvGvV9hWLFG+NVhh24fp4aJ3g5z6GXy8pROt5NvL2NAl0apiaDzt8hBryUR+GkrukPR/quv
LMMIxiutiOlkRhhGYS4FGnZLJh//h+5ktGphjJk0VKmLMnxz1c72/1Lg6xV0SV8USzmFL6+wjsMi
/2EOPOWtmPAhIUrpMVEipPYi0lzkiI0pS+eY7lhqCQBSbO4mfqVa9QYNhm6+4P7QZLuAPVsUYtgH
CTr4900pG/XSMPgFs+37a6uLAcP6bRx9Mn1uucP1TwxIb+C2Nwd9tjGHfIxmY5tToqCr6U4YAYXq
qT0/ImQSlJKcZFkow97zpDGdxxoEvi3Ua3vo2CjOfuEwaeK1ytLqD+cA3pj29q6ArF6Wlmh1ssy+
EkdyRFG4guMKZt71b0xfLnkxMSYD88r6X2/0VNillzqjgafwLGGdIdTOYbfhsSpvDWg1COQ8sT+N
T8W8W+zkAYNky7n8SHruJqWyFKp7LCXsR0DLYyflW4r0We40kAfImGGJPhExm2o4qXn4jBaYO/Ql
1Umqa1W2g8oXeD6qED7mVDxxWGnl6ADHqwFSGbDQ5TLODAv11m0LrnyRU7wxblH531xJ/e7tAp2j
wHMjkjnmUBiWNZMV04VdB4ea7mKZZ49jl1TuJkltC0Vr3UXe8urm1Sh1B72nNftOE2UQZIOSV78v
rSmkBugL6JmytAZN9UJ/7gSYu3S9/SUkB6mZxYUQRq3hfYh0MNDNeDSuOuudc6bWlYzauUSlHBwF
nhbo2b/xbQT3ncl0eTqyw3MV9DmWk1s3fbCL1K7i5S4ewF8QgW01EVCihWAt4IhN349OPklMppMp
fPcqSgtG9MFMvevUawCv8XM+WDBBy3Swrm2r8MbjeMeNivLhAlQW1bbJ9DI6pnhhpkTBNS7xh65B
Z5iEQ18d0sga39TXj0zRXquh4NGF/XHPb275YDpPHG+CgXeSZQXTHKxauR+8LF5ehgZTl+DehBQH
pw8M43UjrpXBjC4IU3VfPVsmWreM0eBIFkXjEEQ5duUk68hrwVGVXZtf6OGwG7ALr4jxRDfuHCEl
efgKlExEJn4I9DIAsoaNGXK+k9GIO/VbbI1qzt6NsHB0P6qYvSfojNZbuew82S/yO/lRE0rsApGF
TZpixnXwAN9xI4cbLT+0969Yv6GamrG0KkRoZ6rHnX6uZdOGSY4b5tO5gKle+/LHRy/uE4UzCozh
FHjdP6gV3eAdM0ckKp3YxzzfhLfFEl7vPMfOScaU/ocuvIBV/YSgwTKKoBwQE2mvWYJ2rByCr0Ji
99Ck4hPT38AoyhYMFDG5ESMynURppwvMa3ZLHwxZwQgtaW7kUP3/k1g3s4n2fmht/6KhsCbbnY8H
mYPS3t00e1NzAY5Y0+nEOy97XT5MP2eMlBTas7WZyLxXsWsdCuMh0541MdwFrqjFVMBYQZViFI7m
T+BeRgFiyPGPygEthuXXXQ7MY5HGGlikdll4Iy/iFOpub3Pyzgh8iO30Wiz6X0fBuuP0wJQYkbL5
PpcW6Y2T5GlJcHYkbm6dXNusX7QaqV5mHf1pc09Hz0jdcLFqBAxb6LiojpQwu41nZHXrQFoQUABr
2Q/esa4sqlduerMVeC0N/IwHp9aS0EqpUTOAwomm7OtMeA1ipsnI1KahAqHITHNF4tx+0cONvubu
5Wt06nR2Sf3rnBder5Cqgz/Kvg3fJXpA6W8tV3+E5mNR1RmOmFc/cwqqIJg78F6iDkq9a4hEAMXh
+haFUojdeRDkYjUKUWWOcdwtllz7OwN0BKUWFuGc0gtC1IG0kfQPrb2B5JMl7enlts7QBZ//W41r
hz9pE8YcKhYZOHX0Hi/vo0lvttfpZyN/A0qB55deqG4nLd6/Q8DXBLNjpzXwzpp2E+QjnOayKg6m
77ni7YOhniT++c4ylkvOwBZcdiKbr/zuSqi9QyFEKITYr8z8N9XJB2amwXW62jrLS79JCzD6urgw
Fh2aw0lWrl4p7CLDGuWYy5d7tcYJ92J5S3sexOHtvjN9FxrIfgMoa0IdgwKr2QMzhGeMeiMv8/+d
b81Z3xbUbG1/l01JBpygEo0So7DkOBDnDIydd8l70pghHS57looGYuboLrL8mzmtPDyyAewMLbzs
skHzwM2iJ7EcD/jS8KPGqHly7z2P0CNaGTwxpug4U+vXTtL0KGdcoVrPyx7CYGjombNMwkAhVe6q
iKmilMmmtyPC6ZCFujo0Mu6U7pErZBmu/sbOQTUdRg6lqIYMK51a881urMjb5b45B0SQCn1hRRBf
nypdI4gmVGW12aa120YrVpMOfiREenZRR78okOal8RO9NHjRPDSIWXSMcygAVBaZeSefB/lcUpXU
mAArQYYWHKiqtwfhHybNnjbbV+bgayZXB7uhdoAMjrSlovVJHzff54Iw3xLJgBUW1I/RP8Py0r6P
Z893JS1oZGBxdyUElmFDEEyPvU4+F5KkvM7GkAgvmGacIfWTNSTCO2vsrNcuoR6+V/F3guyLD8os
hFWyqQtHFsVRm+bgMJuoHJShMAe01TMwEm9EWLgI2XD0wvaLYOjUZUAVEjmsoHqlps9OvAhPVcEJ
6Klt3xI1c4LiDMVKxLzaBmvpLkDUzYsiG+xHDtOAdu4DTF6sHtblyWVVwi88liJ/Y4BWKAMzqKdm
3/mrkQCf6l5KG39XeVlHhPRWzpL2dIiBsQieHvTDrPr6vqXlwe8JoyVC/yDeIucBiNDnfPhhMiYE
EfPbBqV/KWkVuoU2HKQyj4JLFuR2SBVnRk6XL5o1fALiTN0ZFjTb+cc0YmdddHzOa+HFRHPChOKa
duYNdf/f/jHc3m86Nmxsvknpe5a+99ZIf7P6Jj3kjGi5rZV37y7gCk75ig8baMTjH6AJzJgKLcpv
/HvKhCsuq1pa7K2UhuznERMyyrpTzvq0bKFuDKUW9xpEME9mcT8Lh3lMEUNE44cmANkKlrfBoE+5
jdNtCxuoWz10S5I5q0IWk3Xx39qiQDWHZg7m2lXQOOVt3L5hLf81gJhGa7BXdl/2EEOyEJk8No8N
6G2MIskUKzRUK5Jg2CYW2m7qq6nlHAXyCmkMgbLcHdeafebEcbVj9jkagL2phDewr/S/+fSM1Qgn
udttPBBOtalUFij0FuiS+ErJ0b1huPlV9gGYHRLxjN/UujMixXanuVcmEjqrgihMlfN9HoEwhMkM
lXJiDFPQ6vHm477R8D59NdMHV9iQHzMwOVCOummhN07QDPiGP9Llr+In+hF05gdN72YwQiGGlCZf
tZYmmzuzDZ3DkgDZhqI/NIA94jb3m9KxDEUwK2cbyjB7jlby5H0IiCFYoJXlPHBO74z57Q3/P4Fn
eBrrZQEhmZ1jnlqA8PSTG+66s7bGyaYbFPJTnQvlxC5DldaJctKI+g85QSIoHR0atPjpyHv6fdpu
XRdB/U83T35tcfV4wXqGILlLwilOrUaqdBgwgFNFr7PRtlMI2BsctNmFidahtDFpVsdBPhX3BpPi
X/oiWb2TQd5oLD4tA44WIJiZ64AJp/yaH9JdPh9nm/4bBLZ61UP/XB7KQhR1bpi2EcqejH9iRTLZ
GmYeWOwIhpNElsaJ733pQBFsFLdMpxi5h+CCobNtObBgU3QJcnKIVd72f9RfZU1zcv+jRTSYHhDG
mYxc2AZbXJ5GkIaQVTKw+Yx0mLZWQlQ02ga77KMRgA+NO++KpJZdShs4uu9pLVV4+GEZqdQcJLgg
MUFyzqtkd3rJHdkDTBRC30hnEPr7Rv7M6dVaXI046dQN+ojP8UgH0SOcQqXA1WfQtRWSOo2yDvt+
mXjOUNSPWE2PgrGl9J4zfzUx1XNzwWca/Gzaeq8sf4YoAskzTMsdkMDJRkTGpD34NFRbmGNMe4hg
c7NvSifKO11zH/422bu6/+2+qcbwRWqWXSZSST0bKjST3XcFpXBhzN7XIp6RnmjoXYzcQ9w8dabE
SGzDltyO8sBBpHbSiB5yc65jNqd4NfglVEd+2++ZkoVdgu91CY4EgwJT43sWpSOk9rCXoo+fBLuy
iByJCbvB863+Ca5KwFr5USKLLq1s0pbLoOy4/iNYSQPjTxnH95b7Dx9v4tSumjdFOXC7nAlk22E2
wXZT81XG9IsjkB/1+zHV+nZJPG6JVhNCAOZfEUWQSnms/sXBlx65dgQMCloY6KxtZ10aU6XOIa2k
Ro9yNd/plRzLYZDl8pksChtZAClE1IojzzvA4N0RjmJXm56s7XSEyd1tA/trvgFrtLWq7ReuOIF9
wh6N2wJR2f89vmWUb7skS8mxI46QS1IomkcMMnIz7WqQfxjg5ltHW3NPfR98dO/diJjm5GNSDSkA
L6E13N+FoExugHo1FMuJU1kdw9n8ZmrgzQAihFnJgGsRYOisQms2KtrQ6k292fBI3IFgPn5xBdco
fOc1eaEG4YE8+BGntse3LYd5XWXWWzrMmpF3AeQzmoUtX9pPKl8jjt0gleoEWK7rRfUm3YLEqV1I
zEKc+4vurB3OYuxB5PyBFKHNIhozyb1HRVHVtpyX6IJ5XXvPcZ7S8kq1GOZVEdErqzy8xxQfO+tu
k0mE3g5SUdqF1cqXGThK3AooFNG5eG8tUmgCFX/kLfG1kFvqNRQFj2Cb26Fc01MMQHwiFhCpCwD+
5RO1QVo4pLWFOGA+1b6wN0x2wfoessw9FZWNHkHgx6twiXpTvSunGPuCg6RugiATPKnQokswdyed
JeOZKMdK3DYrAX1974hhr0kFLcidWUk7KIoywhpKQtDX7KzzTFbPqWApxnsx6CAAIAybcPtbHRxf
9gHeyUfs1fbkoxFLkXu1eIM2YvWy+wUf4RNoadXWe2WaDaeWM0txzjpWOr5z4PqbiYI7oFxWXqsP
QJ9k52nOiRy0C0FrkIbh8E2bTYK/qG4vy0GxTOX0UI6g2YeHmebYo9CHp8LRRm7HJ85HJzlhEO60
XXzQbXIWf+KBgxkJs/d1rB3ABRV3+KEBz1c1VatGuTZmWXyw4IF5zp4t2lZDprDIriGdQ08mO9aK
+1xuDmNiqHwSkiCvQzZoOpTrrNSWVfL0Lt9S7nTYOyqKXyUV+toqqegEaWJ5LsNwjeWOELW7zVtZ
QszXdd5AwtBwHiKHrv2w4f3dCA/hBXIVeCoP4zxepAons7g2a7mDnI4IztNOl7WamD8bNUNgPyE6
kcgHckyGTvA3muIjUcuQ3L+EmRjEaiOhJ+YBwO3Zlu2Au2HStfJjC1oEDKGxGNbDX/QQ4OAHqhk3
StCwqBJ0t4VBc+bYdNOmuJf5vqmu1svrkxQQE+ZgxdUJQ0P5kTP878bjffJlO1rCQOCG32T60Yvs
Y66cWbbVOcbP8DGeb4QHX8SOyZKgPO/c8b6HoAX0jxdO3lCaEoq7Sh7U20rwd/vJyX/OKUVI4RVj
xH236eWygl56OiFIKJHQVrn1meuGcu1RyFSQ1vVwQzkaY+yGrIY/okNUZTxCPzxKR691VLnNexMz
bZJX6kS2gbSw61ZRuy3OHAIFdjdbSw3/zvTKpcRiiKeY8IV85WqpzYueSTz3bedA6HZOooEj0WvQ
kVMtugwa4rUHZTo4ECJg4H3b8TLgBXhbmcOi1NYH/9uhmXc+hhgxU5tIJ6CynRKiR2TCjGaGEEWT
HZdaYuWMGc3oCtEObDcYk/RHkhSYdax1nD/mp0xkDqTQnMxQukfDqZtVf+fjoUoG7oZaY2VBdcg/
Du9+0YzwwN8zW/BR0WdhwPZ1pYB8087wc6DfL6BLEqUIa52KK5s1WD3je1ZtBP+rukICuBV5j0gs
RTYFOZAPaBeD9etXsL6OkHuSx+IguwL/yASMoAFYyx5IWr/BFcDIJGMJdK1lgarTXhyApzXP1piM
7HwmUQkNGhYqxjLxwxwddxXeCxvotS8liLz6FOdDQWF5PnRm6/6IZ02bl+ncbOh9/UfE96xtnXPz
5UVQJJJ2+Aw+Yi23cwx1dTr/+SAVY/UTmf5jZCLAje9TyB/TpoM17aPucR8L0cEzMWaJNw4DL+PM
nWj/mRsmNDH7rR2362jYO9c1OwCiR1kug4R06zCeNSb4/KghNaXYgnJ3edHqAgXzbMOIMhlViKOK
ZA9Wc164h3ZfMMGXfNATsEKjWfHFCwti2MiUEW3TqHVZb7FXYnmenfdhBFuBfkzkUcxotsiwg+Qn
o/sB/uOifUJqXbNjj7wQ1xFkVlLLm7s88najOJJHIFKXfhmof9Dh50mRom0jyKnljEMzMyU2iYTD
5rLK30vVLEcvvrr4b6IHhE55uQellOpm4Ot9XytGtuN0OFQRoBdAtYX2IFaD/0i+8x5EeB81cAUI
mu/1bh0dkk0G353bL8JPYI+u7tLd10jVeTiViVPDQZ6GLm04T/cEoS/4COqVsnaqdqA3y6jm7KIp
l4VyR+F8m+bKlc7rx+DnfOlJBu4B232izml4nkRqjn+XoEOc+PWUYHHGC41Pie+DlED6EntoApnT
ieCnzV8n0jj74TY+6f66co2Fksf81IhJFR+PnaVc/rPmbH8dKTyea7/PzJTcDzF8nU3grppNUQOa
r4xvmujbHtzbGgkaeCwa2SP9Y5/ttKl19WM/qgaJFn0EzHNNaeQ3jPbEcmEZxX8EBlChaLiE2K+S
oUpAPn6p/Bgbq0fAEevEzHeiMw1343LXTHLia2HXPEntg4PuYTLLZ2VXCBUQxrA1AXfyt3fEZmTI
d3gFu8afshMmxwH2ObYSGu1IHgVN60tg+tFMBnQmctJk7a/sxZsh/dMVMOjBl0AlTIUsGPjsHjMw
oD/iUzvTL5J823UJLjBgGHUk7UGSnQArGNjFO9fBBFeibgYQ1Gy2Qq3V7Ye4m8DJHZcID3LEMJR6
M0BKd4G5CcJ1K8XL1NEe8JJblZmkXhmCHaQTZfzLQafAH8eNIQ0v3dADbvsxp5WJl7gGVl+axX9a
emw8P05muwkFcTPH6cLBUZirIlN0ujfP6OMEsWqA8dMcSoiTsOSHHGxaZO4VyG90RKL1sPZfk1vq
NUfpiB0KVdsYtgXXUwj8SuBR6fwZRF4onTJoceAyk1wfVvqOjBA1ZeES7Jh2tGRBAKfxdzi7BsIT
ENTorTwzi8f+hWena6KxLjFS7tXHBsLtj2fpgGxFoPDkJybe7mP6UAGyENpNAavDrnWQLijhO/SK
yBYABeW+94eBtxojXWziH8DGCRD+M4A3qhihRevJYs7aL6tNoWuVHVFM3ZIsmsTI+8bBNL5dMG3Z
iHXigV+JwS82IvjmzWvjvVJk2+WkKFOpB3ZJ+RIn5sWnePtUbSHDm2BHoSf7Vdgj3TRHl1aY87Ug
c8Oj858TUWvTQGhDCWUKoWS6GCXX0u/n42foBY78pBcJ9GV2AQmObVR9pHR3MPh6I4WVkaRZ0vTM
1N9RWYNKQGHTVZiwvoGoz8CuZQq2iZw1Em2ZQViho7l2OAU4GtasDYS6qDJ2KDaD/zpRUkL7wSUe
ci9c7w3HREKryC6qfLfcfKyh8MkxIypwdGAVUjusCFKcF0vZSJkC6etsTz+3Lvy6klVwwgIaCl96
tnpMqnUHplFSkvfNQ/8Sg/hqfHSWLRG+sUDpjrCj81b3wu0Pg283NJZIiD1yFdFL9iDvGl6isSRx
WhtAD4UYY9wZqQEujl5rA8SgBKLAWB3A93aDoH+tF1CBbBg/usMznv/aAo5cAzD4QiOvIr7FrmJE
KwFL0/UrzrBcHRX5Jn7pBncWfN9BW/+v0bx4EZoi6ItMAF3GBFgRhLloJp8RdnzFu9AocRjpniNH
ZFgoZ5i6GSc5fjrNVYGu7B/znF4kpo5yGKbH8H5dlAihIHd/YsaRJJ1MhTdtfceulTf5llfA6Qnm
40Y56PbBzau4J9CpLvyxIubOrCzplD4xE+Yn/DKU0p1lhsLq/qp2Img8zaeFB6kR83QHcOtVyn6N
Wmrex1m8A+FyjTvglGTA/y3YM8YRuFPJg0k8yVGta3YPM4UPKi+YCeE7GHjoFYy2agOArX7J0PA+
e5iGX+y9xBM1CWzoCo6sOgHimDUwF8cbiEhNlHpG9m/QAhTDOckI03wyCNuA3U6WfdvALUQ6Y2A/
bJzrQGXw5Fn7d0rXCZKQL844tCkJvHdaoGrF75mmEfBO72k4blLHVMpSUTzJcaVNDe48ZFDITUwh
zwngdErgvp0qbGNJ3hGN0LX0kY3nFB2Cqs+AKV0Bf/NffvKxGjmeu9c+o4UE8ctonaAyZve667nC
ICw/oW41zxgBBJXQWSLgt6mpM7tmRzRhNBQkHb/eubnC2N2KrrxeBG3IW6+RnWc9ZP2UmswCtSc2
Zfd/pxlmWy8DDRV291AiNlPIgUU8jv0Pp4J/uQOBAZBlbyt8F8ek9+HcVvaYre9FpYWd9GwfENpF
6LqiHlqkJ4wytGFurtKRJkqXZicXcZ08UyYjR0Hb9V8gYgh9zmJSn6gWBl3yTQJ+OqiJBEIPvUz4
brUvN69MwAp/lWCnwKO1tXI6k9c9Fbfc8XTIwAdAEtLiM8RK9QXys5ejy9DnDv+M0YgIaG53T6Tf
gRXedj1+13UXfrB/7yVzH71zw4FynGrZMT3BCmU0LrFnG13F+h0+1zm9D1MDf0L4fo2f6UsRAUwI
A+PxzALAa2DCH2a9sMrqHSj0EVpZjbPLMufBVpVjIeI8Qm7mzbnbIwBVfceAMbX8uCf9S7cgiJK+
Kr8yYJCZo2q58OYAtikCp26FOgBZosCFPMXpJ+J7meg2b/rei1qQ60/1WGSVRll1I2TCGxuxw35M
6WZx+Mr6+O28M/MHD2xuKY9fKSghClhNAYstOlPv9Sj5k+gi2jgcHea/AX/ruJw9Hyogao6EfZfG
RYax23W2JxavMlWp9RJ2VaisJm3s6iNRFLcmboRlAnRL/dbRAQrd4sRQhfKa6DMB0dAjj1OMk3X5
JZHjQfFVdwsQcy4ZtopZ9ohsXGxvausYVjLtOeCoi//UJsIXGBb2zdzsa2kmMdU1KyYUNtihPOCt
JefmdL5lrOIWYNSt6ujnvDeIGhhnNAnqa4SiVnM7v6XiO7psQOwdfaEDFcH9DJc6JZvb/WEbZxan
bTdB/2Dhcwk/spXJd7P9eK017Bnc5FXzLkUsMWCLE66CwSKi6MHfP5sbCarEftz2zs6/IJeGYa1j
zkkbRwRW7jx595dxoTo7dT11DG8m1vZtvB1gTKH2CHfeKd9DVu1BR/yghyBBA+PZAwD3M9O+JVzW
rMNc7n7RaQLPIoJKp6U0gJIQ8Rd+ftV/ijU+xmO4Q5DRMPjzMWJcgEIvmR+u/0nGH5YtMpbBAW+R
+Psw29AriGGQ24RXFjnSdlVwCkT2utraNqIpAQvgh7UdykizHkAUOdyGvpT2LpO3cHBEGBZPoaEl
6hyV5wBi6uocPflbEy5fWJEu/OV1bhMBuxu1aueobCL0uZRcT9Z0XvBhx4n1+k+hxcpJBqwLnB7F
isw99SDvhvOT9QRGA4uNX6ENDpXWIjxf5aELQN5WsMPgpkJFTGPQ+J5729a7l/N99OZu9UnBIxo7
3PhpMpWa+Vmgnxylb2e0lm7SEPejOw6tcd237mczP7bIOPrOQUzzuMBc9ToMoFhJZ/oT8JRdslZ3
2YRV10kv4ER92f62gEmWGbVQKV6OfC2o1YQdKbYGVIu/fyMZxfkgNusj2HG2FkzQakzg5E8RJrrK
a9lTkgifC8MTZzS6m9YEmiVacBA2gYx44NHlUzq6XitLBp9yaONxngDHc6fhkSZtdtCIKcAIuu2W
CrVvRqiNJgL5bWqAOek9Iyu46bqvJsYp/bcJDf2FYFizCNYBlCRxUNapFgW8N7FSrFvU30tVti3t
gtrHFXU0sR7N51Eiah6Vgn4KaEPpIRm6Ci0Pw1sEJ/t0SPOdoNZQKe4ZHyTHAaC7iVc0zyDcZszG
WKMHO9DuI7R//4QK2AScoySaLmkyODH+eN/QS9zEAD96KdR9/g8x2WuXx10XLbYUjQBA7tKEQKQI
scL5y/YBim96HEHQSxrTqqCPRK+/rvYYNf0rHYKKDMcboaCOTCVdEGNfMJhrdgXIkcS1KeviBVgm
/Epyj5YV+pfxqSzK3TBIxcEQIFGhI+BtJ2/FK/MgN2X0H50oxdVJNYthhI8ddDaFll8hQF6Usdm0
Jtl462Jx6jFYT0RPhaNOQArj6Z3h+6lwtYAsc9iL4Jt13B6GY2fBUFpq/GEsMdRbB9gDoojdvx+4
HrPmklo76g+3Czyc09GXdsqoPz/N+VlCwQdz/B0pNeZ8e4wlSevq0h9veIkm8ay8sHp8mEEE/iPd
CZH7/yiqrb0qZFXmvNpXshdaj9pz2IHV5ql63eK3j376azKqW32w3cmBRyDz0ITGqIZ85eCz6pRQ
bWdzLqvlFlMrTmqSSmVRnehLcjLc6WqezP//s/zU7P97jtMDzja6Enl+E4/1IdlucThKOTDWGtNR
fbAt16Zbs42uCncO9PHtjcDAWpysYLwGsGqZjN7xNQFM2Ola+QmkRlNRHbFb6MVu+X2oGuhJeWmW
XxSXcuPFcKKFtj0LWfxG44WIsuLI15GS16jtWwEBi/TBXABysNGJ85zqONni28D8es94LKbbJCWk
ePKO2wCbqdd/g1DmsnKvzNYsfgkri3CDMU5UwbKAC9NY1GQ/0gfDbF5ZaP8Ql82CtKzBj7kZoEpF
2OEkId2qKzL7oatu0717fm7UxHjGL2fO3u7/NGnZMfg20ElXRvmcFDjR0oV22fu+iOB8+MQP/Tzv
AmQYzMTNyV7sulXitUpAeKn84PnxLK2LCV6GL99JVYGV5ADM9rYFzYSg3RwUdhMlFt760ZFuMg6h
vlUk47SWJxf8ea1SlFHG2Wez/hinUNgUOjrOEw22sctdAnvi739M3PvZucVn67Q8Kj+dpJBPQl2g
XqsovcsCz0t9ZDz4/XTWRp61UPJDVdPh8JJDanEKSWly9LgnQGyusvNhS1DzeCRNYbirbjvkrD/A
CDduE/oyZfBG6njzjfUaP/64gHQjFmK8trv/50V1lHo1G2fraqNkTSqv7VN/kvSYKp13/bz1NPuH
75LYHVbkNPfYwQQivcDXj+qs9jmNiI8XU/sYJseJaZAXZ7q59yEiIqvvEIuyvnVUwQQ0DatdFkrd
Qo1RE6lDKvM+Iwk92/0CBZwOnUZzfNKGHwyPKbzg1ksPtlNutLeNxgtIIBRy9dQnfF9r6Ub43n+n
9rDjrBff+un/wUPNzN5/tdFzCKbkrBcQSyYRkIpZhgHrgv7XxZr295wdDs7oPkFsrBUd/9eGT13j
3xGlzpacEHcehXQ8Iurf8wqYFvnpPh+c4RFS3yl/1sNwGaizEFzO+Q64m1z+QunLX8N+ZCwYk2r7
nMaCtg+iRm/2kmufo36nxP2uq/Z5N/3KkaMhEiUJ3pG3yfqgtqYTqjin7NeZrjPEk0hUl4DC16hK
JL7GKqahgePGsEwVo6wiPxd40JgFZwYSiHqT7Q4Os6n8kLPJ/74m+yxCXa5qPSDzGe+CbbVTKAh8
7TM4+QpRetqpK1tmBbE8P2wPPj7jn8wiukXUQlSAGg31VKAy/NxTCz8CxkrIhy0AgLHOmgmds+xB
AubqTFUfdIgZpTEdSMvGhoftSUu6svkIIKjUamVv2nqi8aLByJQvjfVjazKl9cC3o0H3twl6Rsr1
EZ3Uhjdk2ZDj/5arm2r/nG9/hTa1NqARL5mZGNSogB02bHNwJIYDlfKniuJDFW/rx3ZGIX5kQXLy
bOXceOvRF1oqpDxZfxaTqHLoO84GC02dET+cQ5s5Ay2zAVIRELG/bUc+x1ByQJ0sBLeDWAfu294c
saYnffIjKvsUzFt/VZ/U8TnzSUoUWgaCMuacZalGbWKEKOHe9v4YOZmFrRN5KuGBfrYNhwQ9wdbH
5l8V0+UXL/yyK7LN6604pFS34qvnXAowKW4K56163rmb7I+CwpMSuAclsPNZAIwkX/TT9oJnEQAz
4nucUx+eIRiHccs8t0b1s7nAQQiWVg7h1sgoumiewpf/287uC1RcUOnXHO7RQz/lTHPg+vwdCe0P
Jdnq7gEiNvVB5SfDBO/iu8Kk5MEQJrrdXfv2Jg9Z0aNk50rCh4RCF5OCDscyiho6RcI+tStjcFdC
PYZLiPtx8NJ1o3+etXPLzUIKuvJIc/G05jlkAJK6fihnk0Dzr0zhtzOzE2dIDiE0thFAWHs9JPAj
gSBbMUlAxKtetdlwxwx5PZ9qKUtm6Iy2j5tRwSUHfU9iOx1stR8Ly03orMNd9Q+E6pcxqzVi0y93
4nu/i5RQkf/AbMVZWzHiaLlOBqgzzIUz8+1GPiEf1WdK2PbBaK0+8GXWs5OG1kVWPpXHX9YfmXdK
bku0545EFLxJlDnffvJ9RWHR0Dr5pNJukaiZkAXujz4APrFEOfEKBiEoQeOGtCbbwTsJlhAWQ65K
BzHxuyrO0f56DxLbkYcESwOYVZ2RDoG1Ctx+Bv9MgtG7xv943Z+AdY+jRoU44jiXQssOFw/lMj/+
xwKmvdH1GrgM25e5tgO6ifcgZfjPiEvUr5xw5nBCqlWcxX6M87vHUbZWPzh1FbaKxMNLMval2NRf
L3gU89GQwuySUDupVQl0s66Nn7JDaFCYCar7rtQTqQswdeaJPPkdcbGJde/Cr121oukLVrHDRTN5
YHQ5LHJFs0CouotJ9Sx0+xj5iEG1bNu5pUeFkJqU3egICjBioDMXBaPehfxhoSoYnWvRH0U6OKlu
WYEawZjLKDvtAGbKQ7RjWiXmYzByhbCrXCBM6lX9a2zitzU+esVNQOas7l5mE5wUemcWaCti3YmQ
BtUZV7GtKOuAZHdPXZkQgD1imvOtmXAKbixXj+KQV4xCFWHsuF9rgvOhtD+DAcPlNXntTwh46Uvm
LM3l4BezXmGpShE7pNczLHjp+u7V4VJgb/rvOpjg3LMghsE3of8BvTMCexsJ9/phJTo/yLof45N/
wQYK7nxIYCnpfdt33431wVm25rIgKn3T5ZqFmi/4waXAkJ7ON6J/2TPAVuufUONVF5c2/Chg3WxY
hXygJLaA/dXPJe6oZwCxAamfZruUa5siemsNATTJ7hOFwBceye7IQYKcr5+dTthrW2WZdZ7l5aCq
OQVz//0LkeTU1AT+mAk67WNTk+/tE/55BZyzVf883tLZIngZ+6QTN/fdx29LdbwaL67L2kef2MNK
LHq9SMfISZ4n4eBruJmYvteqdbhd1Qtwd7DmEM2TAS6JoIAhXBXIf4CCErWGhmv+FTqPst5uvtDX
dq2cXYM3zubg9uyhoCGzrSRw8i0BJKl9pJZ1Za4RzewVF3LzBADyyAcPCmsQ1s6OqzucJEmFIvxw
E/E6umuobA8B6zSC/ArxCsIfWzcr0UnEgaIYEtBpQvgF3uCyNMZ6FuDqvF70g8bBkK6qmfx4MBNG
M7fXeWLtBaRuqnGIHk9wHSv1edm88jaoob7I2ku8kL0WFW+/m2QoTJLZ+XgQagr36cm6Z+bqNXus
gfgwcs7qGtuuVjPrF4mA3H3LDmbf/y9QUe1hAhZcZIzCea4n+j7nvi/so6wWJicHcIXZIOEaQRIG
RA2nUl6ktA1IXqTHPiy7Jn11PW9mUHf6Zfc4H3f3zLOKnwW5u6+FLsVqYZMX/PYlPufmH4uLDWHZ
HcpNZL6a6Opq3yh5dQsPiSzq4gePdpIo9pfUf/eGtf2VK88Qv/X9FGmdsb/5wodZKGSOlQL/MWmj
zzkz//+Ar533ntRioKDkZXUxtoO4ahPkJO7MgjtvgtFD6FtA7bpzgdA5InG2I9nk5LaL74hdkMFe
X6QOQro6/wjulNNljaeiHmYLtxgf4iNvPD7O+D7QNDNPlXjPOQvapq3/QQsj6U0NGZPTETj8IuoO
ODvrg+45BVBLVA/w6/YVVgT4/CG8/k5B5xQG4rXlGZlP2oT+5+86qyNHZoBwMw+FCvtUfzjB7lth
aDDrw53oBHGF+RsjStYaUZTBCVPSf6O6s/RoQTbNZoM6R8R2i/JxRWTMJJwd/IJkYx2TXZpzIYUt
HM3Xo4g7cdbrVgxJFb2t3x6g8AJznnk9hInmhWjpr26zsoZpEB77RLmg7VA/AQkaGjCJaiodk0ZG
8djWYLVjOadMEWiyUIY/eNsjt31NOIC26DIdiSLwe+6IHR3zEObV65UMTANw56Fz8aJqzH3NcknJ
meAx6cMK6XsOqa9vEtD572Oc8SfGRjc0KsZxhl924VyM9Mh0/KJ9N8sQ/sviJze7EdIzKCZn3IZo
JzkRiNcXwE69QgApNl2T0j3HRIf8kmQWWVkUXICrND08E3QdxGnUCrjDhgO3rNZ6KpM5gltZZQsZ
fsJKoqOjtD/60beeXdjLLXxyRAnffdedXR77kCdY6oS6c+NjieIYF79KfLLIomFWdTlEXtec3U/Q
yhbe2oio9iSCuoK5qakY17U6tq03CLr/8BEvKIFunDsdcRX1eTmK2YjMdnqcf98ug12NQWY/hbQx
FSoc7WJDCvFu+mffWKV+QHRJH/dcNQTpMwyNRtglRwxFqRbuF6TYkOrqkYt3ARO122p7gPPYbhl2
pvTpOQMboY1UPkiHJzuE8tGRLw0ALqxbbf8cNW/GAeHCHNXu07cf3mpAI11wgark0C1/PvL1FQO+
Ed0yStuX3rdHlBF9qovezdvDDhJuhghgOIfiFbSNsUSQ004emoOW6gsotV4Fqx6TSby2Zva3BSix
SUSn0PBUknfOTcQxSopyURjgZc+8LPFVvtRMt5ipJHXGnnP6HTjl6S59+OzNoYFU2dUqV3d72Bpa
SZy01nqxF+6k+tIS7pKjD2BnfhTXBu7wKeDobBr9rwZJYp5QQXi9l7V1F5XA6/wwj6HGhCLeKpIB
/3wnbPUsl6pGV3dff01COLes02Ka5NSIhdTYnmY0Z/q7pYJKbV8+rRMlS8BZ8MdtXnyR2I0h+GBW
hbBO7YZpUGC7SvJ8vzQJL2guyBMR10GnmV1t5CicYWnhFgj5/q2K+pNPZr68772+rsh8yMR1B1yL
rE4UCp0lt7OwUBOelbl2OZJhYs7nLkFxj5BAQBCF3urbiFBBq73K8r7WpOC/7M0XJnvDYYbXfi5h
tpaTbH4nnaec/pgSpnfKFOg8eHYOH5F8Z4GXS+v6Zu0LGdDSeHxOENIM1Vh/hzzQWp92mAoWuRSQ
cF9sQih6sgDKjvFyvKieuafe/s+3r/lqqLbO3HsgKhHx+nj+sw2jy0m/F/DbKdoX9Z+Qscss5eGz
o03PBraI1+coU89wU74KDRSdsNAkM3JryExsg1s6XfCFv9kaYT9yfBsrRip1lEkLciuaaccU2ROz
zVAmySYsDtMnLsLnZ+MlC8lQmc3zPUELh4DPfUWLojt5Hz7se1lo1gUN10gy80nXdOFXwL+QLV1p
U7y4Bfa5P33FK4qUvPDd/1NODrmhNMmJoLKeg2cIZFNfhKZaNy8ekWOX0zP714LKwhD+kFFDRPJt
Tx6RB6DZfwR+fxPD8GxxZmXolLKFnjrbETffyRANJzAYe01XaGJ+VuDQSXEc6XUxf+qgp/kZebpj
UNUZmpCtnBi2U7CudlHC08Ky+59jpJGRCQ0dp+z8B2a8HHUbr4GzTnOmHzdAi0BhrugBCl41iF15
ZYV1zlIifMEG9N7VhpkbjAIAA0jfAFqzVRgJiYGcgXHsc1EmSRmcehFIynksOaON9shssSybqS6+
p7QrXAInPt2THzecf+SQm+oCiYulsXlshI6xrRWGBLQ9hbj1int/GyuTCpCaJRbI+eKiLUqalj9U
vWJH0EMnPh02rnjvwY4xQPsCDqyjo0Q36kyjaw6XTPbCLtqDRQ8PvblGyayIfxJUWv3kUExsgNPg
5p4JGL7C0Ab76Qcf3+BJACG8HHaEcY5IJZDbQ6m4Jz9K25QNzmS581GfPVimaDgrtEXJrKHw8Q9Y
lKYKJWgFP1f+NAI+D5P+fZ6EuY67hPstvX78Xa+Xqw0LQdD3JOsfbKLXG+aUByYJEL2C6EicTFTY
np/QqKyHWqa46U/6TN6bF/h49c3Hyfe6Q8lnrlZ+qOIAeBQ1yYk/mNUUE4M6KDNejaBtIUBo2Wu2
OLjdwvw7Ouwz7c00NEdv+88kTw7bUMCCC8EF26skbCFBYHlHTs3ioNNPMzRihNsMkk1HXwCcjhGP
lH6nEHmb8yK0DaTo1aoz3c7kgNA0u2JOAB/zyPFOz69Uw3MnrYrIh6X9NKyCCLzZKk+5u63q9/yL
Nt/yE+vxcZzafgPEcMaKUrmvOMWP95mU9h+GjRAoVyY0I5ekdpjx3lEwma1gegK8PvYCuOVPEq6i
4/wE0GlKCSgiGWedOOZTdh6dexcSfmLomWmFAQ3yufYPAa4ZJPRtmBJSZqvDv8oUJIJMSQBvkBfL
kusxdwT49+sxoU4QzjDvVKOhNLg/IMBdDAIl/RaOiVt52W9XBPYbHojdInPTHDERmfG8TMwIdXdx
kuLCeIx3QD6SlZN9wPsH53h1tuASqhyWLwI2fw4q+4790Mle6dOAHoDlDFdV1N2ZD3nRmbFVxhQ1
y+8L2D6mmA6SoMpeZkKRoAHvYbPNeL9jiokvypGz/MnWZjfUEG1JPr+/02GMDnr8YxM4eg5IUM4v
n9tJZmc8KynHh/OIp+Oo8Lx3VQN3Eo1+BEVwTiYLVhB8yLLMjf6z2l3oU5CA3mS/wwks/eskKa8n
ss3HLuBN/vRTCfGZp5YlyXH6fCqpIBJ6iOecdbOXz/0+AzyMn6zNZLMSQbPK1SiaseSxGsCRrwVq
uBlpZNegUiUT6iTTkYJWu4O+yNEHtpShVkpr58y6GsWXbbtRZhnhFOw+Ig9RqrnI0DLWpIyiZSyS
vj6yHjq1S2XvllriC3WYXFsr9yVySfziEkROZubVRSCK3scVTglgg4vqM3Q/2vWSyPlCvxfqmkrp
ShXE4DWED5HVU4lwKybPWsgJdA52j37wDr3eQ2BBxbnyq/UNbguooR4jQE1FTpUMc6tdZpLSg0/R
A77fjom+rWBib3xswEwKyaEoLIWH1zXYE1kq0bupz4DZ3MMbP4KuaK1daToYOo16li1pX+wxydgU
tdn4vhbj/3Y6IqPwjBDmCm+R3FWQcrBIH8S/RDnQGMloaskpn0Qpk61/AyJggoqRtx1AZ/RmjeAW
aYqcDsLq7fzvoDvZ70Yev+g4wXYuGAaguSkREjRYEjp/IKbzy7VV6T4ibyokm0rAuQVU4BKc3l8Z
QqGnFCoTy9+694VOvIuzP7jg0HcRFfUedna92Qp5n+QDZFKhD7arF6byZ7xsSSXVF4eX+Oi5PcR/
3YB59CZltmrM4Y8snOO0fdrM32Km94+7BPSlUuafD7s0g3ioJLTBXMnpyRu3B4v7/YYfYxmLUIYc
5GU76h32XKaX0aAmXeSTXiDjy64KQjp2wCvWSs6qQUMj/kPb+5fdEfS+S4+ydrAqrJwF+0CBK6l2
m6kiEer/1QommlCdV+t9eylJCrQtIqdTJpFlxFggoFDyM+io37ViDBa4khLpEk7BhkijDgEWp57H
B/z7Dhjt/RGuoQwwAsJ1hpTwGBlHm1errE/cVYA9QVDfcdcNi9GZHFz9N4/zhm8axOrHNQimcAXs
synTVJg5TVodw07Iga7aDL8mqgqQKE/xlMfb71rQEIOjcke7sUw5na4qaMQnHHSLSb5OYrAmwOpY
rJWSV+X6+A+Q7jyIWuktIXvS9eyGLnZVUqggNM0Dp9X1dA6D/FIBdTXuuBvP1pJ242b9IutWvgHB
F5jTwfT5LwZ6AAFMY/WZTonSN3wyctEIE4G8Nn2DzzK15jtEIEhSYXMR7wEgj6jVj+RsAMxK+/b+
WxffGqLZ9EKLYyKOiIWos5PNG98Dz0gsKSYohPfLwg8yqbJ0ox8LYYqPfRynwwKm4u6MWyrtVutr
KFViqEpiR4e+qqGxXA92rDa89EZSGPxFb1xhk2lZdrI5NKXC4aQZR8O7y7LFF5pt8ejmzIHgzhjy
6poikZmXsN9F8KrsgUwaqkHD892/Pg4hRd2JWzowraZB1XWiHVIlohYf2AsNqFJRLkVDL+A0Ejm7
ng07nfUPnUTZ8t3K37nK0k4XvbZ+Af7RM8bno8IFTp9S5Z2134Ul9sbrOuYEGQcPi9sZRuqetFZn
eIcZbYVF8ewUOgh8Qpm/b5GU0jpPuBpaF1i7VJQfsQjY495RogyoiPJVci11UDH/LjuplTxgw8EE
uHL8KILJ+9Av74T9Ouha2FMep0ysuo2eESkQzp1H+S8yL/I0DdV9pMYggVVR6vXpd2YYSiUOcUKI
cbxyK2IGlystn6ORD5oL4gnMJMkc13qlBStPe36n6ooLPR03VuC9XQgZjaeiNFHVKzWXPppoYSJ/
n4QZStDtyb0M6RNW9l3MC2RxpwJszSYm8sEGFyHHQ99L2kn1F1RUNOxmr0X4xHaZlBXR0WrMRuxy
2r9GYeO7yKDGOctBOg9+KvJGyiJB7qSFMROf3vJBiMKkdPT6wfkPsL9jYhxn3X1hQwON4+4M4WO2
RPfMz/Xtga9VeFaM+/rKdNDFjGf+n1cMmF7YSYugXksy5EfS12JumuBukHdZOiTPcxfcqZuDGDvT
kBA0D/j3m9tGr50YjsK5TRIN0ncBsaSMHWGWRNXYGE8Mx+WyyOXBgacGoi8kgWLlmuoxME5fAW52
8R+RlrNOcDpTsqEDdfnZJD99zqwx4cHevGPXpsMpbOxMTXfHDTXFel7fcuUxnHxkSyFlJOdsQamK
vgdD0qNC55bGZY+GajdNGQshZhtJ6N5i/9mtGkliFQOQJGWaPl9OhbU3XS8S0+barErm8FG9WaUJ
q/7a5asSJLZXvOWcu1Dvn8KIpzRlFwWfc0ZXwtK2Nn4gMEvXx7WyykuRqojtf5/9ssztLnQSotUQ
Mb6rEnGcY8eR4FBEuvrf6LQZ+pWfFNKeDzm826gFisUN0nN9VSbnJv7o7fRxLzHKR2RNTOXQCmgK
zGzJeDFD/rR3J34S8GdEN7i+XFCugtNN8DS4LCVl204+c4ANinaRBNyYDc/Nq9BFZV+i4vUzi3kw
S563hy60QC30fGNAyyECqWc2KGcwSUb+yx6Ehxb7swDHJdGqexGn+83pRBfp/DaGUvWFTBSbsKY2
MkGZs1omD5leemU5vEGgeG29eqA6fpiGjqD7O01FQngnX07UCgbGj9z/eBGiOVCNRc1Uav2uEUC8
RlUhMBZ07tTBZXNL1Ob5uyDLcp0d1zQt0vnXG7Wt6YZYuCGV8hj5mSWDcZulnwaQqZ0WxcHVJzAO
wEJt/xPkPOiWMPGMu+mDNdOaAVrYo1qu+lW16ffjxN5SBIHIFreZaJtU8GF5L2oUkXW0nRHgWknv
j4YyV7oBF2tJXe4uYsX2L/8YG6Oc9Mbl6R6UtrHmxu/+9irlwzBtJKA1YOVDfymJjMYf7uzPXtuv
AciarxmrgIXQ94+ohxE+xgYfvyY24jKvybHFzyI/xmRhEbYzuv+4gT8Ct7uq9X9PEtMyQNkz0Czg
2bDyDe0mFd3uNVgI7gkQEY1LwjedYJG6k6t/4aIpGmt9fqzinrobfyQhmsv2Z9H7cM9zRz3Ow7bl
XeodZsX7etd709pInMoC2uZ5iSaaai3UisV/x7yJjhOvAyMTSZAdiKcb2drQUrLUwEGwTR0HgDOk
ApVBXBYAk46+Sb4dOmQ5364SXrmJnpvnbVi6DcQektLdSYAXAiuiPQCU/0fzKNpiVQLcb3PHfpfu
W4lRJINexEIaIWPwSjQjJasEtHNXkOJsJJZCVKT7Ir/p6N43qVlokl+kDIFlJETdNKYc/rKVC/ub
GN+lmc1R/qLm4zW0v2MurFo9uqdf91a+KLkV90qDHSuIO+KzS4iXgYY+Jt0KN+nVpoXQ1VJrWzK3
vOOtwHJmHWkJKphZu40R/Vl8E2fwsXBa0xLr1Kdzd+e1jzGCSrio9DXvkXwqN5NFy4qbACAb81UO
bCD/r59SwEXsxl2JpmOqD1uDhHbdiJ5y+z+H1+xQErZQBVcLj4TTAfGRe/4OSMxN1TPSaDIpRIOo
HaFNrY8v967h0dmqNUtJZkf693HhSZb1ZKdeHx84ZzdHsQS9nnKIQmRqMz4/WndExtEr4HwvslCG
D5zcql4hYldH/BnmSChHx4d5i08Oyd2rsuW9U8ED86QwEoRhBzuear9wUVAVBggXqwFq2j0X26Ix
cyh9BbeJLKJQp20dbDXiylczU6PNjlXmq8Uew53tjCty9ubA0lQ1KEdJj0Z7MGVvNzH3ioHyJrAi
1VkKBSBGGtuPoG6xljVV5LgV1sB6VCXMMEYZpICZfMZd7XXtivXzYFFNriGm1N6DvtQbJduvZ3XI
VavptfKMhSsJNeXOGG5qHS7l/yNnCZgwdJF16erQHw8kZSiMPbdAUFnbecg3pBZ9rtZiudczu81B
By2npj4GdE2wnkuOzojvkJO2jC6WUVxvZ+KwgkSOSF4QQ9zIYYGyxl7gIJTHq4YgqjUpT5fOQLZj
p5IC/1xxPNPRsjTBWQ8JYVT5NGjAUxBn3RTZsxbv8wRtpC9UBedxrkQEWYLSmb0eM9sAedIARm5x
citf6/qsHuQDyqXmBRclNB3NMOewSEs+Kp76M+lJe9G3EogOX2eZXI1YkjvCyOIaMv0DxRhn9Qr9
DvlOh32RvvU6NY/3hheotMLI0P/Fb6iF/cYbfWNkUJpb9Tf6SMImyOrTrKrt3u7wWH5EY9jxcpzM
CgjehW9+g8V1s5vX7om5H9jV3g/tuEwDoJ2IvZUhNF5izXl3vqGAE0hlIzjzNfmgcRC/Q7DA9HZK
MG2ohW2t6mecn6kXwZmdTqGeY27j/8Eb/997nvK61IgU8q5lCr3/KSzlORFDFkwj7Ms23z2r41bK
jgf8SZry3Wpepau36G9o6kcVdj6e7nqEMZHgIDeoQPtwVSTdK+EjYFWr1T/swRkByNQwVQoHgTTH
j0p5i49TIF6xsBY8g0ezQUx+Xz7OGh4LMoEcqDcMrkYAuylkSiDuyLWqyGr8zu5Am5vw2HvnqeVb
6Pafc06Qw6n1IBtiPhVvzntNx9z06wyTQPKm97kXL+LirjPfuYZzDQz4cyZ56IY74yzBTAR4m2ZV
2KeQQ5qT4edXacmIyGkkMUA4p5A9K2OZiOKywOzXxzJUOO2DaBMxosDtrzUE5/c7SwOG4GTwWorX
aIovd6MnrnbXp64zSyGjSomuBNhfBkOBvM5REcq1cGq3wSOrVv/QisHYsVjbcv2eQmP8FTzAgtfL
C4e91Sq65dhPADWjzEY1UwPmNvRldLEVaO+o56PzWGa5OKsR4PBTRvhjfWrSsRuVfMgwAjC4w00Z
LBLUKKvU+jdjTUG0XHoyycYWBfvqEXY92sUT1Vg/iM6XVvqCoHfsPFPWZs17okQrFBXgIxHEyFpV
0yVo6Q1IPo219va3R9xw7VozO26j8fp+N7zs+lkrYJbAvqRolDEz/JA1dMGenIr9BM9n0t1Ao6pg
RbFH/NOA+vwuUCQ/sjvAahLQrm99V2SxvaArrD9cB3SWDaAIhKox6P5gYTJKJN7RqMpDIcsTTiad
+XquAIR+Smhy6RLdC1MGPVAPQ+kL0739eme+zDsJOHeSxQ/ah0HS8v9DHKqbrhBfk6oneBWxG+3/
dF21VpZpTKajk8iFBRQLj5D4lAlgPQfGWNO/RuyNgwkY6AP1WbbXidtuLfw60a6AsuBv3r9x3iei
QJNEpVPN313Zt20ss5LqcfnIBQG0dUTeMDf0GKU/zQHXL0lqYrQdXyfGkxLpEfgiJKA+WIzFSN33
SiAw/zS9a+c76wQG/e4pdr0N2T7PTXAH/+Fh/jOaynC5PQIOiyBTlpi7Y4aKZVBsG5K2z3PFeq79
dh1uw4OtGFdArplOO5799ofJ/ow05tP5kl+Sb29PGYjI4ycwuGD+/2g+fnlEn5V5V3XGVthF+kyC
k66+tSjuNOovvw9DZjdaySTfFZoJDrBWjjcAF7TFA1EYsFr7jKvcc+fwpFcoXGkOC0zpJJIUxqBn
2Sm/JqdCRsR2jWd4EoIX8NY6JHg8Fy/S5+qgFDB1R1+uhGNgZ6yRA+e8A4jDAS3aFkIygYjPphJ6
IDrot0PgXY9g1RwUOD7EXktVAgyyESCCfdYMRtyD5R7DQuvZbpP+pxnJXtoj9zVFqHlnh6mCUNhY
ak8VaHVNFsWOxE9Pq2kIYMIFvmweoCvO2XYeDwfCaUerMvmKbeDGB9rzKPu26kblMZby7NvHqXnY
UNhq9RUqVfBOOJO3HXGiuPxBkVMAYULgRcgLc8G8/ZqJ4bSeUeVlsnSbVh0aQs3c7iwxZX1vn6YZ
JMixNxhNJPrXlbpG8UX4qF9leE54FapeePltEg8TWwPoLoOQREZiJMCB2pMccoMtJXmmVEGJaWdp
EvZhIOl+QflbSs9L8zU0ja658gL9H+Jh9zj+kYEXyP03B+RkM+aZPRMALXvc03CU4tn0tmFn40Jl
RPG1hJySLBreXXEAYAEz19VKo8QpRhL6RoMADabDRwYE9fFO0cPri0KujR+sUldEEHeb4K29+wvc
yywN4juHuHIKJ7X0zVPllvFM8LT9wxtPCw1nlhbqImWihPF4pFqKGWs4j0GVthx3iynLNCeYEaa4
Hqc4xVcRQOshfNO9phW2jVbV7aMhNDSPm5pK1xBMMcEt0gybXwyculyukOcIUth6IRpJAaX6GCvp
xP7kd8RZgpdmqmbNWMJqgRXXtGnKu3cuPyCszyEp8hXqmjKh3dLzIdi2R4JaSANjtilGaRPL8tAK
OtUZbB0KWddK2HoA+kslNNHCYUvJaVkGUmhiALc6XCEiWEYXCNaMgfW31IgGTj+x25ev/w9pwRNv
VON5vgjja3B9+KoAsjH3zF7tlY0f2RAWeVLRXV9JriC4n58ky+UWCn2pgeKHBc6GQMnSR6Yt6Mn+
VdHPPCvHmRG+/Ztz8h9pVakoiWFvEWdDsmkGU2Q9XCH5uWoUTEAwkW3gG7zlakJZVgArZYsiRq/Y
JkuvSHDrXvw7sHX8JNDH7AKvoCfG7SJAJKx5V6iEDtdd94NHWeyzCK3lA/DpqeWfBPgWXKeCkFB6
d+CxILrLCSWpMPIsjARLcAq3enG+vUEcrRjjN+lXjlYx/WEJcASzc4MJWJL5hAV95t1hxc438peU
tjPMZpXAiPNdtgKQJODdSEK1henBkJMRtcCdPHZJWEO5KCL1/ogLej511xRbKhQEfTP74Avo6fml
Z0pjGMSpq2gXayxUQA3anvOg1ldsOk8h+I34KsuffKBxN8cqssAmjDJbHAQXBIJHxNfeqPPoOlYr
n8HxG3e2Bbjkj4/dZ/NpkX8WY7VtZL/bAph5rhl/56D3wEvNSg88e1+gT5Ub5dV9e1rAmDYH4dfu
U8QnZAodG9aFIaKShY+7MyFtJRO/slRbCtDaaXm5H+EYhUrItHA2mXYr7aEAwPG0igkIVbc0bVEm
zkvat3Xxb3GME8roTSjR7cLzOFvBuH0jKWfCL4xo6b6DYXFiPxP09CHcBBjg1mA6Yyd0DcA/ww38
ZvTX1c4YoxrbcGdQ9I1bAEC+37OJOEmM7mr7jk2vug82RH3JS0xmBKDXcY81H9SFkCi835r6Aa7+
MlgRQXLryZQNCeYDd0Iai2Ft6tqYve+ocDs+OeTDjgWX1mTnMagFEL8o+grG3TT5YeWGFh3HH7oZ
G31T0MNxG5ly08Ue/Na9JSEW4ALIzMd1ReiHOVhmDhe1UtGpipv0OdD47nvANlYK1w/c+0mpDdxV
BHww+IrkWFCtcl3H3I7Vi08I3U4JWcFizpKw0q7w292n4VOuCOGuq4mWMc3k5WCtKJfVaEas8XUZ
y7C0JOaIGlFk6DE2Ct7MlA+TZOeNMrS/Rhu4hrVKGNAeUlC8cCftno774FltzyVyay64zy4VBwut
elv/eY3PfXL8ILGnd4pOy7DmvKNsTqp7EjoIzW64OWiEJoc7GiSE1TwgsC5pLzs+3IJmYcG5RtI0
7vKJ7E/tOb1ow27ZQj7yEAcaarQg1B3XnCAnW/mOMX6XMpyRQRpGQ4jpqJ87UYSMkRMKyCEVAwds
Qj6Lk3qU6RPfIVclv9Aiyln+uyzkBsPjJS2n4lZMzKzLokJcu5/RAFSCLZ7/5PCQ20CCQ8q65Y/D
YDWy0LbFzrULSwfKXLbxdkTFZ2l+ogNFTUwNr1kdKxlGrqdzXelVWXsh5Vhh6vuVULPG8OYCzYsa
uaOn3uDR50BFfW6neJcKHQISWNJcEHvB6pqYc9RqnctCvSpBEm1EiCh04/6LYDgOmF+d00TUoVcj
QdHzGMJ2dz93sRpt5TwzYZlsBYnPoa7mHATGvcRsP4aXxKp3sVUlAaXGdLMuGWd1ZA0PJIUdO14N
vpNpcx1aCGSRiVlwiBRz/tmDQaHk/6neQXxdYFzmZ7i/qan2OxQyGKnhWQgGq2Xn09lpTEg+RJO7
spBVOcPqoT6E/OnbDaCsHMYreuHllRqDMD8i4oL+sVqdTbILvWVAWcIqo2J9H6vzz+aDAQior67D
KXob9hyls1vo97zbbwvfHqL73/qZ5f2xRBouflknMSFVA9Ug8JJ2l2JHK8yUFWdg+lIEl70o12AI
Iw+2nvL8EKKQb3T/KMeSj+gQ+OUCWazQtC/3x3Jy1mC/CjgD4gT8MnhBjgHxOkg+6fxAxLkqOw1X
IvCXL4mQrj5ACRamq7woUhOcpXJToYMwLuXd8pQB89TmjDS8BgqyK2/5t2u48HgMAFNXD5hzXL8g
ReCEftngUF4f6anTM2CabPPWerot9VazuDMTQAOCi/bGtSRmIuS2LPOaa6DvKRUrLvEUB8Dtlliu
vTvyfuPm2TAtDokOntkk5rh5r7AysCvm4ay9UMl9XxwmdPs7qPM7TENnLvAzsaPHRMgwxnNXtUgM
1vHaiTMFnQ3OuaFkS6BjbytWase0TokoR9/QEgOE9TxZirEIDTqDRwayhBBn3IdjHDamPXaHkm1V
xo4pioJoX3oNvpCiX4HRlO47GVtEqhHVDid+UrdmcYnmZpEO9dNOO+minfdN0SumOROaDzAT2OK2
S7gRbJyRSFkpcStrtIO6RabaS5nmlT2y3sAYPCoR2dfVmZBsMigjzeJV4s9JgeFeki72q+FFRrqM
kKVEkg8KpnTxCfpRaDJ5zh5CH/Y3kbUOLWpbn01HzV8dG04D0DAQRVn8PHZbGyWaPB/fss7g/hoK
NUMD+8LavEKfpAqSt7GRKta3ULPHId13YIAKx9eV0N4OG/ZRxSwspqVnkImwPoIogMj5usGZplqc
ti2O2+TpiVY4/RKM14iXMLnqG6tH7hY6acfXGyfDUnFlIAcc6Y2PZ78ahuCZG+YG5oVsYcu7DjBM
m26z//Gnq9WrG709t26wNNNv3cxf4vet3dNMQd0P/5tlonmHagB6GJnJx6ab9fQUy0pBf5GG4o7G
UlGxtY7FdameCFlsPltkxR4Jv6HWYWs7tdmv9E6PSi0YNOaWL5TUFJoZnNXr7w4vCCmMJJtgy3of
V7fBL9CCNsgdEGxaVi2drbI/57nwmvFDZUbgS5mu52YT2/bLOEm0e5xnVyRlVhLnaRrut989RK7+
RbR+Uoq1yLLVPF8YH7QdJuVDuAaCD0E7/PXESMegvs1RMeQoNTjknz7yn2qQwEvWil7ePepBSX6I
srhYJCzcBptPr82ItFAMZ2QYz3ZGKtrkQHqmAMDKjQZNokmdwTZrEZVaR6568ePtPk8yMHaAmQNJ
vgqLpixmZ8re9xc8Vfx2X1DO5C8k/t/3V8tuHRN9Z6AZg9k3KF8CTXCpWnLoT3XVnuLBXSF092Rk
CpgChec5xGkMAXU5rsGJ9L/bjxGFbvQHN+QiHgZShry9qG2TqCBSgY4fDVFwB16T/1xXplesCA2f
XsL4lzL8qW+csASR1oDlH1OyWsFBnEr6oM7+I4Y+2eL8QpG2084VAq1RwCVzyasIGKuJG5OV5jj3
2I2QGmXNNUf7L1ZlpX82NBiDyu3fY5C2+usLMouX7y/7wMfzHzDltMXw5nFQ4Y3Gqy2aoFMKWbuH
94vnsLoSzNw1lAtqgNkT48QBmNrvZlX65JYpbbNlPb4XLYTDi+kF+sTX+98qkWbcc0NLqHqFcsnK
YCtB3neZzNmix8J+7dZz6uM7f23ceNzaTpcV4eBF2kQ7cwM/ZLPf5gEdPnvt4z+NfkNjsfGncoA+
VHF+KIQtiopyGKbE+VLg9/+XlfAXYB2e0dDfjbtGbO7ppjJOmJS2zvywA3S7CNuZNMZp3oXv/j33
Xfj1iSft/LkBox3/NLrmZcvzgvjaiUhHIO15zamLJae1eeou3Mtb0yuYakv9i4kmPLL4F7RCSDu8
pGrVM01oEq1SERYA3o+xGFbQdFOCx7tzfuAySofcTLxiZUskSy77ydkuQsev/fPa+2SvaVOdiAR8
q43H2u7xaTQoePUo9bbaqjUUmtkZvJ7WSKB2+DVdw4IHxG5ytYhtEgs2q2+mMOZN+cgcpyHKa/zp
8gDTPNr3Y/BW9XD/uQ9ktdTzZmv6aZZgKz+6nDo1fI0NOhZOBAIgJMhPW8BtNQfZUaPxOFE9XUIA
QNS2FvpXFu9kfQYqXB2AHgBJoRCRfeFiiSX1+HTw0KHDGkRktD0MvQhE3lWTAegbUMTXczhbukRo
V93kEAYbud8whpE8jQZa5EpGMoXIZX+5VZCQa94r1iLKCqLvwSWRSFO5YemWPYldOuPRlZ0YDLVu
AAvZpDOPMvVusSaF65TJIVynLt1RzOnD3GmykIZpWhy9c0RIifdWvcqxHOPEsF7XzR8V5KrG3Rfa
cT7pr6jU0SlXInN1mW5yEXdTqaYO8yUStoNz1JGcgJOX7xUeQRtm/QNSka5jqaWsSFe0aAngvUAx
9gy0oBiV+FTyGLVBRT/DTytNiDj6E+2FzI3qxm1Cg1Xr9CGGVCBhyK1w93CdqMX1DZUrFq1tW3NQ
/dEy8j3q
`pragma protect end_protected
