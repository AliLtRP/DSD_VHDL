// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
aq86JRUS0cw1/q2dkRtBlBf0EIsy1ML9c+zuY5ec/lOm4q9d9/C3AAlrOx1yZGMXm1eC0M5pA1VZ
NP9lATAfPR1anADUOW+zFrtBKSk+wUPFjX3TQuVl4zqcW53p+PxmpAzwcNq7trvHNgdgi/e0u1ay
W4wgVmRG5sKZZdKUz3RL8IQ9TWGHu9gQIWCX/qcVRdtP1NgSS3Vsf60Kw6YJo0nv5Ac92bV7ngny
q+Jjh2nL5EEExUMzqvITDEza33thapjxrBgOoPNppfYOo/MaF+dYj57B2VFg1MNRFt7PUu3bdFuQ
Jpc/Osp4sN3mRUtRvFtsQHRVHY55fU88fiWRww==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
3mO8A1+MZC2ufW8vTsgKJF67/0pPRvlHvlzmT4tLjWQNEEbuZAkzRFJrXOfHbJ+w2TURip6QsuBb
J8J72X9TC0BUx40cKJLLV3tnbwhcpA7CF8qslYvr0/wJC1/K3zSw6EUyelEGX9A7wNNKCYUzfr+B
tRPQGfpiRK6l+5P4zXDzymliMZRhb5WMpSCMVlLT9xC7VSMW8CzgqrmWD72iHAEXE7mFbrFwiuL7
U85pqWCZrGB/kiwC7FnGe/728S7aeN9WBqNGjqlAF18OEbbMjnnh71SfZS7ej8JRUT/QrCaYUbn+
zFovIev7rnZPAdUxBlwl/ZrJN+SlRocx5msqTPHAonJXLlqtPR92WXcqOIhU6Pg8FESc8sH8li/H
sChrC9Xr5YTCJad6RfStBE+7Ia8SuIWpAhjG2UHSQNkuzoR4akc4nEK9odko862PZfUsR4p9angE
17omesr3/mwdyU570aNgi4LTHb5OpW7cHSzZpEV6Rc10UNVrpH7g7+6Gyz6tPnI5sN7km024owPi
T+2bgZxch8ZPMB4ho4yYG1uWEMpuYrvTIl+C0Iq17Z5OvTF5H+dqTZ/Q2W99fGsisyiJIqtxyJTb
yhyQWHuHK4byCxWIKrvqZ0Cy1KOTIJIVa8lA+UbfW62HQv3L753RYCAvetJbP+o7ZPrkZPvpFeVl
P3QzVm5R4UY233ghKEWFn9JHgoFK9cX7WX8lZL3Q7zMbsaeAl/ccv98cnrBGS59AXzfWSlvJ8/4e
imCLtKV/acufMsrCFzMimtN4Yuq3YSyCRCDgckesKgOJhqhRCOjEyTQCpjIGLh4tduV+/lzc/4V9
yPDpRujzQB5cOPhD7oKs1hXN9yYRzURPP85uYmy7BekVkA0HTSGtvbrNxyDcg5Q0Deddw0QjcJXT
FL7v7YncPvBh0Ro1ObbHALLjoXN8TGMSpEP7Dfmw46HOCVBSpO/xzK6ZrjpIzYoaqjfMYNDfKhgz
Ht9KQ50YSREhjOxYm+N3qqWh+eqE3gH9yTVtQq0Jlww6CR3h6RTf7qcjzMwmoBFrvUrK7G4wLK9g
LMoXVFdNVz62EbVEpDtkvPl1tCxM/TX8dRf4usdgm3WOQHrjr4kipZv04uChUTx9OPzkWim6MYpC
yxWjGwP/i6x2J1rHpKUSaHQI2xMr9cL2o3SmqhOg308fefCIOe/1dUb2y2yFgWHFHX5F2cOGXKUg
ltfNAFygDhyRQA/15gsdVBOIORqx07dYVc+XGhEWaxXVHZQD+9IC/jILuYIVuBk6Iq0bGClAvVgh
h70Axixy1WmkwY5qGYbBbBpD+xd42PU81z8GxeAEE3GzFbaeSG/WFrIB3IC570OCEw/uBTpdfckg
PB6bCLKhJbtkwVDuCSlR/R6AoDAxI+7QYd+TITv61Mo/RPFDBBYfHWtAPknDC8gtWo2GuJ1ItDK8
5r1heSfHTre9ffnALDf3GTaCXYCWhSb4DeHiy4Pmd182e/UOVKj16cKMkYsnmISGeG0UujVDbk6m
j+BU28XWGzRzlfeIrOxHVxDiPL/VDLhQ2bqzsXYYFDhtZciphDLNyumnjZAoaF4VByEpHMfRZxSR
u1WLf4QxWoYtOf+rrdjNEQx9JTGfwEfb5s/ErYWbQP0kZNj4c9geLqlTJaJXVWoiy7WsrozwVeet
/OxUmWrZkFfXiQY7tfe6oS6XWjmr38WHQXDVyc6JA0DsgMPRGs0q2ydaZBAef3JkEUf1e9S+UfT4
VQbCR92qiyjB1vaHsckrrmK0B2bFJXsfRvEQ29K4J96J4gxcJ3DJT9c4E4lfalRJXgyFMWVsm0+D
cmoZRQ5haNbtqGigmLbWnXr+9Zm6M/xJSGm9uT/Pzb+GUFzKs1nC+i6pWuJFEpvL+PYvyH7TmKF4
ymnlBz5VQkdTS2s0HsJi+XzndIsrSTMtGbJVcczUx+uK07OO0kz1peSwwHBa0WoSvO3XT5yL+n6z
bsCUJBY0OEdWTGyzNlo31B7i/ZoxOau13RAOOtWwhlzTHw/70sd75H0HGKOKgjgJ4y4RR6U2mrHG
ztXusVejhA0DpKRuXUB4ofXZVTkNboH4SFL/WoS/7NyS3aFt83+lXIVLbak3D/blwSVpiOYWJ4OR
s/bC7iWX76IArVx1sreUwBYs04/AspoproenXzv3fWU37GEOep89Q7urcSSE1tW73p2a7z1c7m85
O050/+yM/mc5wjjUlV7uh+kuZLzCCBx5JEpLXPqTFqDRipOnRe1M4IbMfHBegQbus6wQB6P2x0l+
/2n9Z6BATJLyqqRAviOoNjF3d1nMoNOu8boMgt5nlREWrIaYPEX3cl5a77AFUmaKoI8raWntCyaF
V8LN0tb20lei6SYqhBxQSQkUuuepzGvw9o8JfCiPyniMYB8asU9BgM7l6Te+ektQN3z4dJD4fv/H
Z66c7Bj8lefgzJoFvgo3vLzMo8q4aA1YZkA7JFKOIbfls36kVYTES8uRybRe3vDvS/xE/OFZDdbL
qKdbgROJv9tPRnpkecmKviqal9XEBQTmpZVD0j5Mh9n6EXf9iVPvcQnXFGtyv7wCOTVUwhBzWgBi
eXxFe1qd7DMofuaDrgimc9Zb6Z3FqPdjGKi2d2fFRaQkUNScQb6hkaej9yiG8X7Ct73qWayFP1oE
6vrjLYnV6Rkj1ZVltHXQkTycyDuAW7LlWe1AOcrthZckzqQcTkruDKgqb4BD+NziwO2wc/kO84Bg
0za3Mj9glfcXcetLdsHV/OIsx/qRVGpze6EMsWqxRu+lu6gUF6K61/jy5kaRQYwCNxX4kB2MjUup
xhowA9lATgF67SC/VBvMN4eWq585ucjFZnFIRF2vSxLOgTk2L0R2U2aO3uWwk7INHxI8ZH+JJTJT
vChfu8WLQmbwspg81A8cGC81R0o3Ymh6KHZIAmSEUn8YgTUdzLxFCdOBOTOs+8pAAVW4urR2TXJ4
k1py7RhQfYRd80bff2EbNoR50zVF69meQj6d8KNVlSBNMHg6ZJxfkD4uZd7upEhdbZfqwHK7kE6c
WQpB/Yk5j7rC5I51FR010ruGPxQxVkpVlanfB4a1Nf0hxyiltmtWO7lc9+UeWEihgzwgQkD1xDZ6
Se9O1SVCsYkl74m4HxiEcxZnyY3V6o5cO5NjBqmp3u724HEV7xNAMajIUxkdgZp0qL9ZScEfd0ZM
koGkhvgqclwUnoNk8xeEcaH2wfAb7GhZHFbzImoLxAf6C0iPmJzjxh8dthZaUFfEW5Nd2JGtj5nE
3GTnvpekcqtGa4Rbg8kCkVPdNupQxowF65KWWTVuIJt0OPWI9JDY31K5aH8oIFfCYTU8KoWGyYOx
7tjDGuP/eB6lDcPtoXsPVljXD00sYc2knKa2yDYOl5d5wp1uROxJXocW8NWEafSkIApdY/JZltPD
I2QHwoU20lr1lvoKBJpItnOxI6YzTwqDU1IWUADP4ccq7IICsAUwEc4h8oiGt1/Y4R5oKet/7jas
Hd4RQNLdOMRmOy6cvqOKAPNMN5TaRk+08bwIkmN4Qj2P5ezbISPAJED2uHmXDb0h8Z0me/+oN1tV
mUFtXR+5Dpae8pAADfaNsshhDbPNe+VdwA/OyL+buZNqRdu/Vhes4Zs4OkswJka5Nvl09ARNcqDt
MTTKJ8BI3ACkdcrsW1lMjljNUn9H7OGAHLtDwi8SLlckcgTFKFEXIkgghxN/P8od6Ua7K8TFbY0q
4qq5h4qUEYAfCO9eOKGJ+mc/zq8LdcFOaFT6pFL8wdcy1Q3iCUqKTLEIH0K7+x8J6i4L/iPZIjn/
9JfEK9BK9mBf1idIHNkflzXdS/Dfd5JVMFjEjBf2c0w4NIMfKJkg+CcmNdUin9x2kt5KjFodgQLB
8YrAgVLJCZFVjq63S1vZxKxY7q3OI8An+XpAEiqHAERoOdJAPMrrVG06siC+35iJ+mLHaDKLb0R/
uU1XwqRf5mXML5Jsm9jGshbHaT6SLBH7iMhJfMldU1RKhvqfhRM8eMjefcoBame2gqsQcjgRz9JL
UqG1YWd/Qc9X+t3b9w3uqu74HyZyzXLVCjJFf9/ps+1Q+rXiWBvAzK7GxfkT/3Iq4k8W1f263+xd
zguBz/k/bcTsMeB2FFJ85yKfSnb30lzegp5pl5epnnK2XkNGnHdn/l9YMAJlYEetBP3pl40Ze7z0
OvxatJ9ASoDb6Lb/bKIOuRnmGWSCq1pUhqLWo4yxyRo7E+xhP+RCLYEkphNiglFGqul0cG41dMZb
ViLStSmaqS4M70XZGEpb2HHkftiNrC1i+SKkrP3O/OB7DF/HYNZv6yNXp4SWD1NDU3PVbtGUdgXj
LkIWgPTIBV9+kA/yFIySyBAG91l1JiN1ANr3WfRmdMrkzG0PomKYU7606kwg5p/weU5CD0lNTfN0
gF1uIlPNW/hODfo38iB+c6eyCZ25HJfOjZLo/dvkI5hMRYHXZmytgvIZMUgsNgGoJorR5tMSYcNU
SUmUV1va3Zk4VdsSDNDfjufg3Yfq/HvcS1hdhr83i8bznRBWTA8ZV7pWPFI6k6UG0Y3QKTqZxYfy
oZZlRfdhovvyv5c2tWfYnQNrKpNS0B9PEotSotpxiu06eARfM0hsqXshJg+AmdrefhaQuB7A9Ye0
qPiT2Us/X67462tfBxeHSgsheC5eDhyG4ihYQSqxn2Ig3i+Q/NXNLKXnjI8lPxlm4doSibkqvkXU
F0m9gLQxdqr+e5W93GrKJ3Wr66bzh2RLtPi//E7lPGTIOmS5764K3hvHhxgNDgsSQkCgcLVXsFYQ
9xXsXp9gsFg30Lbz+itUh8RxWcQlN5xsYX9nhp4nVkW50ot+ZrrkjCvYZ0Gnp8SieyTHGcSjRsjs
hhtOeHS4rlm+gAgDLEUMElkdS6NySYAXVNWtsjPJqrqLrfGIdQraBRPRVlUBDs6lSWVcrFDLMPB7
yy4zJM2EqDHaTHb5weyuw/+9HgWr2fk7NNFtSXe0Q7bTkhUB1qnOQzQ12njmPTVxBfoqMaWCm2gl
a+4jfUbXywYQ9mCwejgsUDCJWrYwtMFa7xTGxqyWRp9tcGA7RFlLVXqdwT0mFbxJ7EEwjKzykxNP
NkfVlBa7poKeQhayTYtCihpko8hX7bG3lYqigg82PuiHFb9JJqIPpzEpICQp5Tc2GU+QZ+u1bf16
7VWkhPJeGZFnTkrwmoVgOJiRhQ8c7M1J6SAS7Gl+A46Yw/F29IsGjkUE5bIOlH/q5lpvehd57XXT
V6SVmD25GNKn+fWaUrntZfl6FlfcYS89aBjDTJ4Z9BqUX8CIZ9N7lbhvpUg7ejfpqcPDbNHs0aMj
lq6w91l0Nl57uXzQLzix0mfsZbvmUyQvIGuW9LoeelOybVkgRtvM5RebayR9WQdptp/AHAlUdOW7
5vsdJx9A4+P32x4/FYq5QTohG2c//g2VzyEySQOsYpEn8VwrO5H2lFSEAZ0AVf7B3dqSop4m4L1u
q/d/s85RU+xa5+8Oy+ogpG9Y2WnhIQCLRtqY6Gxj0gVwy3uPZzwNSuURanAZOfw14RDspQeTwAuB
ob+k8PtX8WNofrpKdJbtQftrk7qHntgdJHs4Ef832oEFK4noZDUoGV7mszDy1/pfzrCbXH2XH/rZ
vgYerOBNn4koCnEBHzYWIOvVL6S9Dqht7CsmuCNOUz0pPOVWbzeyZuRtmNq8FQQ2sY8GGiZ3/XDg
PTY3EtlbzbDJyokINEio9PmDPZy5m1bqOb0HWi7yEERRkIyBgy884xvPLbrzsNhON1VNs6cdT4+T
+j7rNDwiHggXgSKcfC1iBEHNrx/5My+bVbRzv7QnjnjoGryt5+Wd7CtVmGkUq7wpQdmCz/VO/JxT
6CoG/OqjI/Bg9FZO5tVFXyTdMGedw9rx458+JDxbDK82otES32Dzs677lhp0wBbqPiMQZQYLyZMt
AnUJEPCDT1vMoOJeAOxVL9mIAbiB5ANqlzVXVGQhtPBskJNx1GnWdZvk0g15pz0yrYiTdIWcfFZb
xg5qO0Md9UmcXMOmHjeqWHMHYHiJDojIfGksPxPhBzMPWUp+hbVk6TdzqyxjAL4BSl01gd/f/ihC
fZc4WiXG3LZ9fKT9z8R+99ucHsoGEm3JmgGPEms1bppxlRoiEJcX1TEZEj7nNmVoJSSQ1bf3hl7o
qEHIHL5CTxILU7pa5iJTFusSVD2dNNGGcCywGXuXHvSFZnBVze9AUQDBg0325f0Ol3LUy8/2JqXs
0MDuoYzQq9oTYDoQ2uVqFUu4PS+RHvSG0eO263b0gylg9CqVRj7HThw6mynrEQf7lvQM96dbxPic
KXTOMGbMEzwZBhFkpsk+B0p0OMk7tNje2QP/tOA3DuARnmZb/OIICo/ML5jyv7BMU7osxpLFkSLV
G7/vDTjHKFxT18oMYFfdGt3xa741q+ykz5KEyBHOX0dLvSlqDKpulublxzCJ0deD7XmP/8S4zQF9
pHGnh9jmcYexsz1Gd3WXBXDx+OG3k7KUntRUOIeSJOTckDKRfCF1yCs5joi4jvqdyfXlvxwj7Gab
n6gSYFGfG8AQH011jf6NjWbBFCmt+jSTs3cIPu9QHdo0hv3MCwUDfYvgWZUdT9YS3zBXt91+bP3X
ZlGvITZn91aXd4YZQEGCPrU4Cq9wFpkS1OwAZfbUM1r3jinAzzsNfIC/r+t7fX7I7ri5lxC1q26d
zz99nnPw79pVa1pcmcnp8x2sfdqLfAX7aHRSEN6asQnCTAuFWJjBMB3qAY080anO09JOqlpOkJks
Br2A0GmF2eU9URqMxX5++NeHGtptnjYFhn4ski8y6OEXzgagPUZScEvA9IwDYuzZRpnt8615F0eL
FTs2Q/T1MEMoSbTsoQEnfhHECq10xh5Q7DNziVYsKZxkthneLfI3EuU6D6rXBKC7VvaWZcoDQ9ml
snBnl2Xhh+77FSSfaRvCFHL0CGjS18WjFNO3jSAyXe/Pw51zlWKhZ351sT0EkEDiCFrpGj6gRGzA
r/WCyOnsgz5IPoxzjE0PAH7Pyyi0vIUFAW95B3J3bvmlrl6kmpS3wOTuvU8JEMr7Bq8RnodS0yDe
YPZSzZxG1ZwBhWFW7lxBmdZxPewUg0kH7zbbIjZncx09LVUd0lP/+mCSUoOxB8uGCsnTc1C7PaFa
vsmDxgSJqve0HTgKNi161DxLjUC7VX8efkII7tz5StGo+FcJk6OfbZ1m9YJcTwip3PcxO/aZO71o
iH4yuK1fOC3QBAo5QwToVtYbZKb8MY0wXpgyP2COkERGE+ZzHTGkL+NlcFDjuAgmbUxluOfh1sT8
a7ITx/HYnCsSDsTwQtXz7k69+ZZsLcGTaozpRTR3XTMvSh/VikwkHlwGxawtpqAEPv1kRbfFODH+
4kpw4glt4jRZrv6tdJhPAh/F0v5/rZOZp2UG4iaJ6xsMx1Xd3Rmzm4aUgNQq714dwVubDpPyaKt9
Bs9ZRRcRnqz4YPYkU6QJPimcSsWGllXRZHGZ3i81s2eOS96RN0CoLuT0QmtGfkgsl0sO54/SkzuI
yTlhhhHZn/l77GIvrBI1Rq0vjR7WvgeNixpYgrRPdgI3ar0/2YJH814Cn2/nuktM7TL9QCcL5ejG
ea5awRXG4s84XjIoDCXOZdBauGt6g37Lgrx2AIzEco6xLhCpnU5dfuTCSAnVTdZy1QD5Y0yheslg
cMSLMDbjlLZmMLhi+3Cmnvc3NgDUq2teNqLHwMcLkXzIA5nRwlT7QLRtL5t1Jk4dWSZT1LimvTQc
b0rtMqscGzp/XYugeolilWT6U+krErHodzcJDuZnlfasKhSAxS60X81zoqkJ8flUeqkNj2hsU5F0
eEckBmO44Ue7BaM5gfwIPLl625lsoQPyDvaWifuVuIgMruiGxfcSZf3N7GmwLsDNUptoyGyViokk
Xa9rI9Eq1YeCpmR9Z1qMNWrkl3zjhEv9
`pragma protect end_protected
