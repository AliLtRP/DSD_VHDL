// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:43 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
SLOsbBBgW7lUxX4Y/f8Rtkl8gFX6LEMTlfPnnduyJ9fhsYthf3sgihN7W+fZSDlf
2K+1KGWs3rqpgtbGBD4EwzIElgRQJkmHocPTloJvz2HrRXX6I3pfwzB/OKBPKpnB
5U1M0aSVn+yijzz+0ZX6U7e/IVth3KpoKxzQWIvSQms=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5392)
+D4LcwQ8LNd4uBb0HrVMEqXMKl+gAElLT5B/MiiMDXxX5R7LwD3VYHsGGsYCC0vx
9/1ZnhpYVYthseqMPk4mGjZW8YQ+VzTTRcterSaOJhJu9hbP4coMaRHY9fcy0+tt
AFyAo1cup7Z2pRVSiD8a1ji/2LDSE67Dgnc4plyliI9oIveCgICN45lhHJZcyihE
UdGzV77tt95UVSfYMNzaD9oZ2Yf1+IGPWntdr+kIgMQvWdWbpqHsPl82pDTUFVx6
kgeEEzwI7ikY3gK9dGuSjQHpZJlMAANyYWc1BQwO9Epo6r2GkZwDhBqr+4AYNL4D
LNPKYmjdJY6Hd7A4votVp5cDePa/22Z3y8sOKQsZuKw23WUrI+6v4jgbZGp50FF7
t9CNiFoohI9FabY3aw2GsHzwlzyO0EoEbRsne2ZvQG6AV30optUlj/IZ4FLIhTYg
nc24E2rxK+188F1jAHm9Q06GMnsvaTsRKpFZdG6qcey3wmlWvnmvyZDVmIUBjqn6
3Z/11al2L4kTERSW0e5/M9R99sJlDs23EOlToQeS4fTtLfjHwezBofvI4rZOFEQe
KdRwoJMiQdzTWl9l+IDmkElh1gCqfYLo2GrQ/3dGCBbxfhbr5RIAuaZ7lIfLKXIu
TXU2lSR53zUjVhtxX3Kqtni10Svc7r6HydMhQ26f1OTKl2Tn9bv+RVCt3bkKWZOa
DEDs5dIUXR3r2XcJK6yPgRfxnbL5tQsRwUQrLC9v+cyp2fWeOewTkqa9EGgtCudT
/bb/ZSNDnkKimE1Y2L/K+m1gFQvtJpX13JDWBmhINfkNgMQlIkiaXOE/Skro96Zi
8qilP/ToWo6n1N1ouUPHGHYlB47gpoMoVXmla/QoSNg/HMlmiqr6Ttxcc0cQX9u/
ccraUWF4N97qFUR7TN+S++u+bQ+9h6VBItT9Z/LvCTKWgc6hIjasyeyEqgqHEHyw
ibLJlqexI8Sx5fZeT1QyMhFPwNkVMI88BoFjEdl/v25/6VCLeSCm0pApclXuxRGb
ipgi0I+5YFkd6M4wNOGP6Zm0beFR067BAW9ggADrlBzO5zlOf5d3BicUElhMW+nx
jrYCXk/UA0cv/7UGGkZga3xnH6w6y8NpJYOfjoksPvMNS6a799f7i9CYA5BRJ41p
gGbl0VyvOw+0OjtMlmkI7EJaRkrBC1ZPK033wyeGHT2D3F9Py8ZjyaZ4J5PyAnAd
1Vs9Zy/i0PFGFtXWG1NZBOSl7XemnzdKakY/u5/UQ93e/wRvQRVkWVv4icqG7YSE
OKVgqDlEmYjRaB+OasoXPCT2Yf8twkH9yGbpPDm4EFv4pC2gokA6NqwUDXUkI2k+
Mf9TSosfmycZU18pGWmL28TAc5xFOsaGTLUe5ncPphI0izpcCZcqWGNTWPQgsmbA
PPPvMCt3QG/uPw0B0Jq7vf5YSPDYtJ7o+Uptrk+Kt/B/2lkev1RFnQnR1y6Xn3yH
jvPF3PJ4CMVvo9fbQeUaVOGFEoO8cngfLWr5BKkb2KRUu5/6Hz4f/37QkITRCN65
8KvKXbfI2d8y4RHqBieVrmBYmF1o4o7Pt/h4bx4hKkiGL0NJedeN0+Xltg9PYYTR
LJHNb3WmidcKlWUnNCOCHbcSEmJp/t/Xfy6lrW5RHIDLsiijdA2j0dyJLEOk13Ja
XL1ewm6pypwucr4QSF+FYU+ViUxi60pC2m3P53pGdt54cdoXroD4TrcKFyvw1dMB
E/YvpZh4AKXovtIZL+I676/rj/WdseX3E6rVxq/QPdsASV2M8HcLLauE5yTPgk9V
coCDloWyq2h89NPD7/17si2Vm7tgcrCSWXt6bLh9X/E143ZdLuRoBujOmVTqG1sf
R8+zTd/4PqKhVPskIqTAOH4f5r3FiRv0l1/VNl9nWWQhfD3iKiKsOEdFbn0lxucs
6wemu2HOjgjrxD2rk2YG5tY4PNlwmwAYo2/mmSO5olWJBakZe/wN/ERiN9smTrmc
dNqJ5Euj4FW6rOClfoObkYVAxQLMFST8m9UWES0ah/vL9S1Y6hHJC/Yx6OwMK0td
kpmInTeONNEaYy1eubdb0N9yfjXXF39H0iwRbuUQHlOKeStLPCk+2g1Ml4IYbHl4
vFWSC4AjaePg2oe1rlVwMQc03V28rxy864HMCuy/5/r39EX9tQ/Z/+FmXSvNF141
y2So1ZMvUdRbpQnaDd49N30cZfJRQlZTzN2EpcNeIUpYmxiM0uQS/kFmJbb2nuF7
Mwcs47LmT65v3C1D4SaGl9ZWnLUAAiZ5+r9W3oGommVFf2I2QcQ79BMnfgV8hyPu
vcXzip9CPd/eGFWc5C23365X+annih++OvFF9A00sO+1Yg+lm4leZLmZMt/8Fw7t
r8/zJ1f6cQeZ5WnmrbQFIgWORV7Um+ij0eFAjyaUzP3V57tOyfwNgPpfiKKCdgHK
X8ECrQ+JalPnf05uog3w+28plasW/C5wbXPQ71JY4+bnvFEewK9fEzvZ1FK/mE0l
lEhtI92kyMd++hOL2ttRspgbc67gaGqvf8nZetJjSAh4433fBCMRKn/3E8y0AiqY
vl+ps6a0nr2tfdojH9XjmA2fDtc1XrpNHlEAyHpA4vXqp0Rkfkpp/rGSwGojb5gl
6evx4CxlcmhdTD5QuotXtXCl9KantA7R5VDvI3eHItJtCCpVcBTEQ0VOUZE44Fis
nf/KusL13y1ND5P3J87K7MQHg2PuE432DwNVODBUnWr87pj1UVMTfGC65QfpYGXx
G/1EXQ0PbnAwLMNjG1bzifH6gXHQvyu8DR75f0ANRk5GFAtlZ9cOSL0d8JB5klmR
1eAS3DFhAxTdVmJL1GXtwThRiCD+zk12JaK/QfeuHAq5f9li/M7/Q68sYT6N01kg
q/jD4MxBwMlRTT0oBjWEPfleekDBSKrJmKykqmNzaCrS+UpJjN1FItLeQlXajD83
beOQhRI46EwE20NhUAsJ25mUlNkUAEYilPyf14waRVDhYuhXMv7mocLZl7OcTMZR
3LkqJhGci1EgYI42xPf8/tprPGB3kk9MtkljlcJfZt2QEJLCbWJNLewmPzJXwyJ5
Jiy75pnxr5KWg3PqaFFkzsLA/qRmfT59OMuNZC7PEqlMSSgTqQDoMjDDYK9oiAgj
4teo1HoBHGWJGBdc0wmlUSVZQD+oD/BfuYNKYncw+c7G3HD7ncW2abtPL3IRoO+h
uKkLQsW/7HsqHxmjIagR/Vx7+vaZgYsCj4/8NZez47UDnT+hWuQ4O7IkcWqyYBQm
7zB+d45A4w/nAdNeXJuE3YboQFp76cXkzgn+EWAvHVGlvqo21kPNJ1wEmZA0Oq4q
ZfuJ2oFWsDBnYO8jbjko8U2T7CzAXfGU43jjt2Y7QNNqkKJymjUThbjvUj7Qb0sn
VNYWmHuTMUIGC1pah8O2sVdPe0Pdw3KV6ZaW9pIauAEMewSmBzCC0i/R7Gy3oDcm
bLmkaEoWhsY/qE4XUeSK+LBfr8zf8/EOII2cG7JEoXdrlHQQa5nYMlYewXwyeSiR
QDf6RQ+Iy+OmwDOgnmBvA28a8YHhfpVfM+SumNQzzgafl1/pocAyWqvOxHk+HgLR
TdETCmZQCcfLzci3k1sNsZDZdXzmb5UtKcYIAweCI7w+SgOlkD7Qf4cDH1K8QU57
Lk+TNwyGpJmMXNb+oG7hq11xMNTzQbiQGYNpf67/POQ6iPjmj6/su3yLrTCU2Sg5
naIOb9pj1t0Kty5HOR/22nICAonQI4giNps4ISxTEZyd2ROjtnq/tYi6zyUbqlSM
hN4t2uWAIDw3x6c6bdbfe6y3hAM9OuAtc16ANEthRDyX4QT1ASYpslUkmj4wGOMW
iaacEr/oEmXmEMK6Ht/AcTwBgi20gVWHGqyFmdtVz3pAUWPQYq+L9OAd+l10HLRN
iIwl2Ui9hmDXGGwaqYtCWA5qLhVcRqHSgwMYDfbER/3az+7FFLCqlgtAIxN8DP8z
fRZyo2ohNu9HgYUvZWry1eEKiFyFmiA1E81DZEqO1tcsegkq0C6AtwuuLtWM2at1
FxBwV0KIcL/hCfTnH0qfYKIht/LrN5JTq/p29GkVclX4W84gS3pG3bpQZ1IOvUX+
/vy7O3IghMZdD9YXMoxHBs+eY3moDuWzCCxtSbzzUZ9hJDyItdL+VaK7pWjew01O
G6uswEAbMQgaMa6A5jN8JRZ7TMFYBI5vRDkuzuZci1eVJvK07MJALYmAN+zbkP0S
kYD72UJgmIWy1hNF/1UDtJAhF4FUbwPJrb3bhixjrX2jxvXiD6clObbZ0nz4+deP
kyNwt5yGsxJut5JAlAlrr/14HVfLsLXP0TvR63BQesRWR+vyGFXPfCBTyMti3Oir
68N8I2lZ7WNSKEwut54a/wMA4ERTOWvqOqio0dm+sML6PyuOglXd/YCe5AC1tEot
QHuQN8Vzn1Qg8+7EhoyVYP+t7Rf1xPXoGOx/3FfSumURSxnfz3FgaDb16QmVYGV4
mcyYsR5EB0fllblkySOf6JsaE4fkFroT7DbTxnPY3gITXPiENRDbr5KolVIfhb9K
WanIOpb0Dx20ds5/lPCrhxnMn5JKA+kn6xpfw33l4xU706ddKMWuqNGaCdpB4V4W
jpZ/KNwvjzWY54FkpJMJhQsP941nuw/11FfbOaMs9jblD0J9yjchg16tQQM+pZD7
GAyuJ4XdyD+iKI4R2Xv5oJTjNh55BBcOC8nZtms6OpWV4ZR9QMeSWWWN0GBx3Lmt
E1ntjALzlPEXDPIgE8F+kZ1pr0YyZ6XA94X5RLoRpsx8w0iNOIr6jfWV1XkA/x4w
px6NUXz/51zGqvRX3uIJNOvmRUMQRIq4W3yfZx8C+oScsUAKnXArLcXMfPgDpu3K
kibv6qWkdwPhSbI1lY4uMc0FeQcqA4FmcO14cUtJj+Ug0GKh5xmRU2HQul4A8Jp3
1V55oRbjx0Nh8JH1bEUPWTrxlOyJfvGD9OHVPaUvyFYZ88nuf4jEPQu1H/Zo4ob+
GGzBTQGhq3672QBkBl4uCLLDO/t5silSJJ9Ts51fmJgsEu4J2ePzQ24DaiClMQKr
On7wFDpw2HK0gGHeaydLc34DzJtDHM2odWqekSQqKT+vc+qdAP4XE4hNOtiZTJmw
Ghk5AGM4H5QntsK/rM5Svu+27F4bxwIXKeN8D7+N4D6meCuwxtAZvVC1uNmGvLqb
2oqf7s7IJUsFuCCCk3fhuBawPw99PeeGfNJkMIbVQLim19wZCV2cxcsIsVqVnOyA
9hjeMmgnpv6bRqthf96DUVplYX0kNb6UrLDytkKZ4A3gxAw0t7f36E2hSWV5wLUQ
OGmw8D6T8a/LLwGEqw0NYHSZD3svOc1OoSQJl+CT26S2Mkp+YS+VBMFsONc4BYdd
xcW3rIw4v96jMKFwAcTeK6D9+FhqEXiaTlB2BUtX1p1tww6jHdVR7mtknrtl0QJw
dVyiNkUzm3Ax/tKdBs3DjMRCYTjzN+bs15jxDR8A3P4/1RNdhInvyH5bGAlObOPN
c5DCOt790iHOqvUytjNeAKZ6xAB+h9jk6NFhMTdqjAPXFH//ULVEuMEvD2ngviwC
aJFRDcDwznQl8YxNC3GXKasDVpN6PO5kgEfG493ZQXIK0/BaW1DDkNZokXpT9DcX
2yLvu4X1XyIlfvq5W0Xe+9NxBL/9B0iO2LCymiofKGOWiwcYR5oQhzSrRjEwKNNQ
5DbtHTSa7vFLOc00vChS53d9kpSFBzC4YpKWLxBme1tPjgfA9sWDT2gVeYLakFla
gjvIvSsWQs/k1mJlXnqEH7QESPCBjjvFIG9RjN1FQYXPGCb44uKbkwjgaYxaxChQ
ueUKx4w5MXZAPRfeWSiq685Lxd2O294zvoXEEwTtEEQnBJ3lzZ6YPlEO3ZTbYIIn
xeMvxBPgAXjlmDwgKoTLQRqwzQ9U65IWjqKsz1TvmZgqXQfvqqJf3oH17Hajb3jW
s6RBl291TZquEERooy8a1gOV1rombIXa2p66Cy+wjTyLFN67DlHkTXCq4aYz7QqS
JJlDttVXeI+nr6UNOYOi9LibQxHUEnlda6vTuhUWpARxDe4p/crxy3RJg/wR9ZCL
yxfjt1S/+MT66G1djWvL/14Ksk4h+Gt9fFwHKk2dmvI/tDZDJBU821f3+vSlzY2D
IZUF2hPDRs7AOGEetC+WEfoDV/ySL0Xa/9ea8oz2/6jFcex44hvwBYiNurAEwFp5
Kg+NPcsffAoNDUJevndgEYLkPeMznGwydSMEV6yd61U5jqzIXlVeHx+RPjZVd/4W
g84ZVa24WlN+JHX5v8TfgtdbZ7bxshzbPBQ4RL9musSl9iiVrOLjrr5RhR4fhXAR
8W1zTZMtCqy5db8gi1/EzF/F2ixqmFnmJPV1NncSI45eHL6spoDh2NYSShoIDhus
hO6EpFeY9M/oYdi6TiXesjVEYGXOv4SfxJXs/DtGYntFwRrDumJUT3/s46zp+Zqk
39zjRHgn2Pb8NH3AKrOpRZ2mdEZKPdShdjskirxiZiMz+vF/LbVqX7mCaPWYAbM0
GL6IPD2y4qvKfRPKM4m3qDhyUj+zrfSuDhsRu3mzSgNUmtkLRuC+EOapa7aVtHzO
jz3Ip8IonIr4/C0N4RxfLJoeltro8zKsN4fxSQtmei3uSYW38jrF5UWioNeAeRld
3GTprBWfKsVa3HK2XH3cX5hbF0wW3Xi7hRXsve4trGKCEAQi56TQQanpNHhzyBaf
saxbd4EEAnJF/FyMkLDcWiUQv8FN/FahKqzOBo9st6XHth1mNWHzZx5Ouaz5hlmZ
jGkUuyJtNfYllsfnrt7F44jtLe7QxFoWzfW9bCOkMw6PSAzQCTELbZUhxVM5p23x
Sf3Iumjc9CHnfZw6FKp5Ssx8Jv1eKn7+0hauLR+Z6Qhf7mPjElaTxOH0X+E8HLC5
xNScLatyZi3GEGagAnabdHnarv2ELEy5/qNnQK9pGgtGtbi/h1xaScCIRhJLi4Au
GCf6xVNreMOTmcC0ex152Mxsrho441Q3diOAF89K53qL+jeOWvyl1WTDGf6oB5Cd
JcVVMfDsaP9MlvXWjHHdSkJpHhSZIidjMXjjCO6piH74YF1T24MJw7xc/i65dFv6
3UIPl6IDD3Fe/gaauSvwRxw9eJ9a/MSP+RTcTuz0TUlC1VWFiuZ2FiSGfnxeFWD2
qOL3eJ1ofQvTXmdmTFDsvw==
`pragma protect end_protected
