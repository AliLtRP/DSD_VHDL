// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:35:52 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Gorno/qOANHKBwTuIiKYq1T6lBdgOPDFCqmSdSvWmfjbcOyxhLSP5+nCw/hQZ8p4
v8v+YJ+8DSUcxfZvDNhIP3lJTfF1Et7bakv/b+YCS+Tdbl6b6V3oRxFcVwSL8h0t
ZK8aAVw+EbeJRaept3+7qINHIpgxiZkkXTRhr2yzpus=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 7584)
DNnu04zTBJSbwhminbG7EfwceZTlVTR3iSlqOXeDSquIjSge3NN+LfFXxVMEmW4b
YzyvZoXcUyBYy1gCptTwu98WXceOA/puH5AyqVHmXJfH77FlqfCdmbqBRL210LHO
f+LsRQ9H9I7Hs7n9lJL5HBg2DthZVsJKobyjS7lFUT+F7K11hktyKZiVZoxfTpZR
ljjMqwzsGnxxi1Ut94j7lT5eLYVZ1Vpsa/JEgUlQJWdTHDVbUQD5gcFU8njd5ODD
BdOjpgzG1cgLzuIHlL1zwJJf7UdXP2aOPl7S1KjJwu8z8OKGD78CXfqxTcgb2C11
7puFfKZvVwR5TjQzI9f5O6N05G03aXL2N5rvHKobflfIeoJUufDspmqsw66bT6jT
C3xjvpvO5EgEpEfDvwMUmsL/pZnTUDBfCljn5EZY2ZZEJbbwvEaiCd7l8XAx9w97
U8DsmOgoxIgx2Ar11k+8NjbTQ1H3NW4dNP5kkAfqGPkrCfnfh1RzdDunAia7nlId
+OqzWJuEnK2ihAQDKTe3rxa7s+hSFeRMPks6m6zAvcRoVsoTsd3ESxzFqZRY8e56
KR+UY15/inEUwwYUu5eMDrepTzn71XSryR8Z/YjNwGui7mrmU/ufK+11w9o6R+wu
RKewnXg7/F5Q+TvX27+jKYXbeIUaYPsuSsRaPLCI2cJtzvkqCBJ+NQI+950ss+Ay
KmF1BjzdXAH7W5LOR6RoKYAm7JdOBs1XRJuSMxqfK+s0gJtPeLI6V/FjvOgeKgbB
Jblc9o/jP+0bd7FV6ZoLHbODJA0JkDnAM6VSRpqdWyr5wC2UrSLd8KErW1bBmiPk
WSjF0FZOzFfySnpEfP1wezPvbMgUMKLc+FIeVSzrXH885L2Px4EP0BgW03p4M44Z
8+Hle04YgirBLd7O+wDXDU+6HXHBGLyewq/JKs0K92AbNDj8c6uYq7m9K/0GzUGo
nN425TeeNuVtL2tmOLvUNPoRkds9VfS3Ni2ZnH6TD2uKniaSBuOb79svfSvnJjeJ
QB8VFnKF1TNgBGcK77jIscrfVUNk/DKwKhmFv9SHrUetYXOSYc59u2njG0RF1Sdx
3qfH0t0iuxh9nUUbuF6BmQ4bisM/YJnlHyDht5SaYZeokFfVPitY3JBpFrgV8j0C
F2H+I34SiBiMybRFmIkRw4jzKjQj7mh500FdnydqVrs1/eAEpENzNCsRjRhK59Td
g6JDKvspBv2SBfyFV2Bnjd1j8Cg+19GAg+MsONuGPBntBn3SazFhZL+y+LdM9i5q
tBM1sloYyBGz6ejiifJGiM5V4zV3tjFy+RvSk15WsfFiCR2qUj2lJf2t6iFJ9aVG
YTNOQ2IBE+Aujy3qOihtH92qHqcuwJ4QGlOL/ZIBeIHsZBgwaOEcwh5EeeQR2j9f
MrzgPTrSROdJxDuFkkniPaKE5T39ekfjfN2HP+jCH0CPed7canIOD4psHbnx1jtx
cE7fzvDPr+LNmnlihiF4Zmik/XYn5QyLeXs6GM2McZJfhfVBbtZXmuu/j8sYK8wL
AJ/+ELAE0Icg/H3WCiiLaCGlhl5aCsuE1+lah1bMhg+fgnA1SuMfxOP5TbZF1rNH
/e+6CCmTRG7j+/Hc1zaeiFsRHw7Lb8FP0jAjRu5tPuDmSDbETHsE7LP5eEP21DCp
OKOOB014rAL5HUu7VP3AwlJOegHnTaPAxvJrqWO2LGjB6HrxzdQ7fJfuKaO5H7Un
iO82bpzJeValTwyEfJpmMbovf10qT4tGG/zlaYESWaLsMywf75S70Rt4et/z+lf2
LIp5N2HDvMWQNUkdbc1SgAzJSS9+p3IwQ2Q2D01PKA61lCMHexi09OxKlRZD4S3G
0dzC88qFIGZBOkmaI7C4sTPpLhWBaIeA7DIYUyv8/zB53GhsTrrpkyjlPBbvfLlg
yqysLRIEgiAVMKPhhfgEMuNAPuVoRySwZrBC393u1O03ddUkqi0lLLTAOqA/P+Bk
pIgm2trUkHfxWRwOM3n97XyZQ9hc1JGfR6sfONoV6NQq4gCuzAAeNoyipAtGmSlb
PCrCSeMSPeHHyBP3Snnx3bLQTR+Ca7ddVmo/K8jaz4tFdHqMQo+9C3iu5Qzj7VtR
DqQm0hpXv4/Vjnn3XK2ZuOWZ1DgB827wCztlyxPWND7QPKWSo+ImLT1TaGKAWYI4
9VAY9Z0oZ2car9UJamSRE8vC5SZrVwdiJQCk4i44C4HdPltEfX0emFsq1x1vcc+g
WRKyfBZ5W55+HdxdWTNLk4mi8kuTI/Q8/7ghhnlkCFhmQYUQ1RC1oenFSsnHLr84
dYCFS2NixWuDVG5uCxTFTrYK/1DWYz/91SFkhQFahZ+XE1hd6R2Kg8D+N1ux2KDM
Y3kGbRII4aCRwt/AJVSsi2vaxGx4aebxJy9uEGnACKLZEZj/dWRoO1/VolgZsnVp
5emZbrFN1xejVN6yfFOA8FGkPG1iWzt5y84d3Z+1AN+DkwyBrX1MEr9y1RNSc1G1
RKinRQl3sHjc2xmkRGTPcPVum8GOsQ8JoslNtVRNPfRTJuzn5lYw9suX5AXJ1aEn
NCPHmFks32xtIJCrC/YKRgOzmFzkDssQ8kq6PBX9zuisU4FR9/WZV9wGVnoyAdJ9
oEQ0LPpqpV2Qnme1Qpcgzkj9wBwBUfK9R3fpTzn1Fqsk7ziFeQlj+58O5LDX4k3o
gvu6yY5dP0GS9jZW1NOVvlcTmuRrqO0K2D5ttgqGLdxtsnhYx5petoHXeGb+1sU/
Y8t5VT80IvxhFU5X3tGaHAuloYJaECE9RZzinLaduRa2LnL+xRMb/NqYgvBpxm6Z
1IFO4nMhPFtev3im7VoeL+0tMCC380QVUp6JV29YKCNdaDURYpLwOwuqpWwegqTZ
D165VzHWDbyeDN56T9y5rPrZQf4rktzaXNdJx5K3My7x3IF9QWQ0OHE85r1Lhxcm
zNOTcTeu7hWvMxcJuKbFk5oIC5jMUTjjrfKn4o+gACdLX4uG/fQ0TWj/wE8UobP7
71FYl0zJHIcfniUV7zyC8k5t4Mzdon5Al9bP2lETPzRncU37OZ5P7QMseYAn2q7f
S5UEfAH2zXvXnGHFkh5l1GomTcOih4nkynqaUvvUQ1LIflCkN0deLSHYvQD3rdNU
aJUr3ubUhkFPYrSZ6uTJGMzwJ2oW967qrmtNGLV3O9BDrrWjGjqu3MF1fj0exW9F
t5TqS9jS14H8/138EB3GpKnsK235PEmdA3wsehyG0UfiIdlF+vw20mUbtZkRNT7c
WroDveBxsPoAlezPKmenvsela7OhkHRfq1JiIQAkuqKsCuaTcF5N+TN/ehjyqVqN
wU7cf4QMSmmg/ab77LzKRpMFK4vqeM5GXoj2ZS1sNAK1WIHpewG3yMkQy73nnfw0
MBZsuIaWaJvPYUaX+a8zp7N5MyGLo8Bn1UXldmLJkLNXP4+420XqmR3kEws/LdDL
bKpz1VZaCQ488+LXXTviU0yOV1X+0RBE19cRogofTX3d7LSK+O8hAfbYpzoFnRnT
SUqYBHWYfPSH+8kzdYuFWJVzhBP3+R6WkNIE2JHP6qx3/MT9F8XpxqOqDdwjtDg1
aEXOQbRRRPqHcg50+54VHeV10F2McWxrCr0AFxYrNAywnCfwRcaetiP/xB5z402s
GsSje477NOPeQRTGjI7b3pqZutGxohltzenFU6mYNicbn4QY6hteIHf0f4N3aeQe
ZJqXdEkHXRE3kubZxA2WKEk3THGr4DkgRfclcDUyDSzJ8Hbsr4hx+k496VLiRF+C
wS9Y+449EP/xALK30z4XoXclnl96mq5Z6YA+Gr4/K8y5AuwHeoM4tQvH2kEZ2Cx8
9VtensYow/I40h3hCw+TTFjUT+RonA5HhTmIOEN4qHNCxwqf/rhN0GpkexD+3yJj
INBk23HXkIERI+WxiEOKK8cNbMaai077UPhKP1lh/vMsEiCEi05Z3jS9jcHf+BFX
7zxBsPxsfEc7z7Kh1WvjnznbgYEW5s167yEUPFeuBkLFwxX5uB1TssAzzh7YRZX7
kn220hDw1zYmdtmffi/KZIN1ai6pvYfVQyZYVXJKeHpvOSNHioGUI2HBYaj8is32
EUtktMse6h0BmiAXLzVvgHqez1XpaT7sBqdupw29M3OJYaDpPcjHL17wQmWydCS6
spii34HN/hYBhUkp8iowIYjhvL3kNJsuIT5Hi9qGPmImjHyX8BfGiAl6b+94SATQ
CzA0Qq5ZapVj8iFgplX6SKoKQ9B/RF2sK4O8ZpXWYhYb/xhLtyeDXfMbJ+Y1kxz3
F9cO3dbd8xaolEGa4HGlngyefd8bh75sZKP1zYmqAAp8poiN/PNklxLdPe4A/wj+
eqey5OTuaj2qVNtuB5/i66luU3HP0dUf574+OTQ6UgJxKz+oIksp+oBn54etl5iM
RIADWWU9UmHr8D7qmfka5TkuF1NDW5IzD2MZv8NgROHdH3moxVu8wX7rRUuaeSNY
rsocK5xRt5sdqnL/FcmSIMppIEtJqVBLFgDqhcWmbPmqFVlArrMJ/xYy/CetextK
n8cwGa1wy2m47d+vT86INYpeJuJQ3XEhVeHA+xzAXGYAojWEHTf68nhjrtpwgC4/
jUMCu21r6210KYR6hSdObkEEngDcDLJTMdpVUKz3hSeXa0xzYt3za22gjcxTExt0
N5RSPk87zP7rIiw49FyyY4mBVS2jWelew+oCzQSC6wBVPwfvzZzmVphIdAIxr4Fh
pc6hol9YXFj7w8eBRFSphgWQ9PHgolS5nLo9YOlFWNEtUdpBl2Ki6x9hptTwD4oZ
sJOYzyYbQbCWkfawd0EWXqeuoJ2hbY1ELktT5NQAJ/I09rSwHRnuY2PtM/QRRC7S
O3JzQyF9dFsmAUDUbZDhtexZhvbQdtjcHDnJW1MgkOOLdUHiFgnpC/MxUMy5qY2r
p+nL66I95RH5HPlZF0/C9jIs0QbT/4qTvKtY/FlwRNvXuwBODKWTu1KXiIz8JiIV
ZGwciou2T+ngR80OLzgRUI8BXYEhjSyJ9vOgsTSY3IV0Zks8G0djorhEVK7pXTr2
HkCNLthnshgaTKSjgaJi02q1agPHBsxwLO0AcH7hJ9KOAKknl7KHtMn6ZSBFlhpJ
nTZeq8O4mbIOFikGv7FNeaLGEyHd5MNrL2mBXcnEos9e1CgLZWb+MFPXTq5JSNFf
44j4A2gVLIbiazFYvWWO8H7ri5y6gDcDY5mlGxyndoEWYvw1CF4pnHKH3TkxX3Lb
Ue0ciPGsXXoxuZp2reXOmpKmj1b70KJE0+0YD4nilfiFOUZgNq2igXm1eHQEUGMJ
tglAOHxpzSQoLZ3xdAzrklqMAddBnnKe8bSxw4vsN0kr1JolK+TpvvmQQebdyAou
v9tclWHF3RSb6hk6SMMidOrbOtdowMVwjTBLGrSsHPwvn0qm08S4RVQG+wEHOMq8
0FO3PfKQFPIXHYmlhocVFG2/RMpEsBfQJQ6tuRTXvttdMTwFlwQcWkr/zPVcvKKM
XZdW1FXOq8naYUD7zJm7HgxDiLBe8dU+xSQyoCRFgf3lwCkBS5sRBmBBaqvxBxDg
KCKtwdyHiA3TPv2YfULd1Je7cQWRAjeF+Rni73RTxQ2XY9VmYjX5W/TW/7Q5chAO
l0MD/v25E9OAzfmeXe+9uNzH1U6uJsEQNvVvuEhplmFvQ+UrM6aMiQKR0B5PNirD
oUvLnsSjNoZJQIpTNWeoCX9mQgMutmRnBXCMa7kyGWtV6/m5YZEg8fOj0ue4HsU/
r00fLzlsVcVUOVAC6yH22fMgkXTgpk6OgtQppfbXgUo4qI7YAKwIYgmCesyoBGgN
M2utlJbTu5lmp+GgCcUEmXMDkuQAyrDbWP/SIQ6iGd+wzTgW6mcg2FMw0AYnT8PS
tHy6SZkg0tlKL0aQtkhJEbJT34IU12ZJIU6Z1m/AWKdPdbu/twR8Ow8QuVgUuupi
4g1UuMo3IPKqcBbBmP7cant8bPGUVJi1nr42YW04OaOJuxKUorCWtHeYduYW6Bs1
CL3g7M26haToNarRh9hws3Z4674L1uwVf9q1qEnq8zglt5vMhnkSHfD1OYyQQNtG
mKsBS3oNByVUHYAtml/1XZSFCJfBJK2VA0DJlTfvRDQMtZxxYS0seusNwS0ixL31
9TmLz2GB3gbBETQ1UyjiyalUezORWXn3GmY5o9XKgcbHuymgR/gXmL1uQOZ9s6nA
QuzaT59LUey8jJjp2eMMj2+mbRRnvg0V70/wDhJsuIE1lBI4RKRnJal5gRJ+PIZZ
yO4dTs5hoFOoOFZlPNgxruj0q40QiDMtYej/GD5i43UbV1AbYo6x1bnfgPqk4Fd0
ZQlgm64Kia0EdhpcqFvZ25ZKM1uKQglOKLeWGgVn2hAsXxP8b5RgevPgLQ2IIxqh
xX8T+0SZzTahgpB8Ph42C3Ncc2HqtVsCQR07Glu/iTcLUd0N1IVNi7FeEY6mi3li
MUuOT08LYFDys36MPWYd0iV6BQspSXn6d+9NQDQqOxPAQvcrr3WuGi+xVOBJ8Jx0
GRsovnkxdgfQR51dV6y+Pxm9tobzjGRq1/TUJgjpeI5vjq4Q78UqecwBacY322Wt
WKBtTcpru7Q6wN+Sr/Yz+G85/zSj9aoor/0St2Bi+TO8WF7t2tJbiEZoxC/Mp/gv
unQ8k+wVYjaKPKKpThF0l1jnJThffCemdYS+uUb7xGJRWaIBqhZqvahT+6n/w8xO
xv5xQkGehsJDOHJi872MLGha9BUaUE8hb4URaUEAOScm1hvxv2L3wB0fsu5SI0bF
lVOe6lUbK9kHFF6rzHxBfoaEGAsEdHgaUrD1NZ2E6JrPg0FVLjdymb60s5kRNZda
1OwBD23Xcysw3HkAZmk8C+GsGj1+uspLnSpWK+zjKvO/UvoBDirE7RRsHkPoFIyQ
zQTV4XIEi8BbAOncEZ6buVpFlJhoHc/W23kv50/h/qDG6EqrOdWW0yC0fBzYUyT3
uH9O+PAblI+PVw308T8QQAj4qBH8VB3O0frSO3y+kOq1W+TcJBmSQuN+jcrdTBJm
+1elmiOcn+4mHC7UBIA+Q10wjGxNZbkLXr5hidY5rvB7NiQXsEACEtjvhtC/wc7h
FyjWAw6mQMI0IMe58+8Opq3rki0n7EuiH9j3x/DIQk3EGDYJZM6cFDfzsY9yCcGS
gUaa/sYrZRbeUmWwYhClEKT78mIWoNOZdqXuFMqE7yisVewr9ob9Bypl8wz7Vk6L
U3hl86a1EXyac1+2gSRYeWgs6ukN1H57XEc6Mrv5Y6D1v5geVBsokb+QVFpr3Ts1
RWmdsewsmi8JuZs/VJPPsGE2xYBYSK3xYPQoIIQ121/xgYBgXYwnhgLnvr/hBWpP
X0DqGRqsNJUq5FA2ZoClFlqyDTeYBa0egcHfu9XSvBWCExLjwnCvDZpQKNKRw/Vv
GZUsOTXNbjh9tcZNGSKUqpOqDFNogyq06ro7RfA2p9oKJTXGsXG3Xiuka4UujKg1
qFQQRs2d2cTyEZMPcjCMNnTlMNAhvBaVhIaqxNG9qQQyxdCfML6M7o9fGkwRjcaF
m/3Q+ZETAXwAQyBymjJQr4LIZmsBbldGrnVj0KRSye7VsNx/WXi8LWOaXqpXQFyG
aPzgUhHWaRD5uOyry5EYmcp/4TZm7miPs0QtUSeDptK5JhtdfYYkOe/tSgE+r6gg
Je1bGRs/FH9LclgVbGbAxhtzp8PVplVeAIVen2RRP4RKqv0QjxDSEuP9swZH2VbC
iFbIQdrshUvOZS/HZ+gNUMH9f3wAASZ+FTZhhAIjNHIx02sLRn7XIKjiO5LKFqJE
uv8ZHv1+ChxAmg6xdQ/08F/afe4oGn5MTYSOsjiE5c4p37qJmeI/sejHGNRq0Mn4
myWtrwqFV4qdVx8PZCObHVxX6rNM4giiiqwehfzoc2PIjVhSaMIourT8mecA0dYt
Y3LVE9Pr6uf2L1IicmDKPLfx1uNE9mXGf6PH415FcfsUnO/sZpyjw+HOz+IBf450
/lWPmk9pcmfNPgOMgiT7dnshB/1PNiPEmI725s9TRQFpg0xvuGV4BsAaJwp0tcUI
pguRghIn0HCVKQIlzSkb3hTFEJ0FbrmD+4ZMsXM0bG6KGeQBCfm99yqfNsJYgNLX
xx9SY10lZh1dHYVld8pvw3UPmOipeijsKK0YLOoUSkEWMaxrDSHG+MVJKAT2MG4e
qDanOcCYd7DHlRLilnkmekI9bk6xuxPCPhIWx7rfFhX/vAqu04fT0i0nsIXTc+pe
JD+If9Y+xxeorjfXGAUPsuP34YUDTJiPsB+r7gf7ZcqKvQdh/y3a4pPK0dU5aOpk
wQv55lptsDZBf128mzzEaY+Jczp2hgFilcxl9h+plyvFgIECWpuJNbAqIbQwreSx
cnq/d/qpcNJymQR7+mF2OqFEi50MdR+JurWZEkt8P2rHB3kP2y182RLIeSywrEiq
5FxY7dvYRqsi9NhWnIL8OQfm2lwcVsQIaAK3ixf4pfrvjjoxGfH9wCM0RUhjbWkp
vSlevjcP/RbMlZoK5kPHA+UEBpXWaxwnIs2D2xy9K9eH3JEUoiYee02I/STKcf8K
7LetzWwx3wcBLj1m+pADBumXSlWLZsZssGjrZBM4oiwhb9xZNg6dz1I5V+jt9zIf
NHOC40LlVvPuA1bGuvSm7gNcmgQ+4gdns7fbIgwUMWp4n8RfAACOHOCP+Dzhrs3+
RRhbqFXyDI899kC0MyqGf4wXNvsVHMCqoDYXwPQvfxHRWiFd6QQP9OgS20TlvNpM
uZYpsxK21KrktiXPgwBk5oboAby/kmwSaOi+VeYRTXAXCR6F7NXOMvsgf020e9Gx
n645eczlceaV0vUgj6AU74h+oWcV59yf916C9bTAcNvD6qINqusgKBweAOPRZMMG
lO0Pmw3mZYcWvfoWAaM8EwOARWijOSYOUDow/T4HBo47An7XLiwlIZqU3d3WBI4b
1G3oLTnu5B6BCQffGCJjFXkgrpSZG1ioqLpA3etteUDwrJWYFPzUQW4/Hn/Y6vIm
bfqGWQzh3u7HO5I3DvZ21Qp04HK3KMhc0HsXFB5TOnD7Rb0RM/nMFG6VgkT9d0BU
y1FjqUa73J/5/JUgwhaOV3v8/tBDcb8O8D09bE5aWu5neOOr3JvCF/AbBm+F1FDF
qRBzI/GVBlIjsaxDR3hFU8j3E/ebb99dgbeHYnCZ5HhOnce52UL6l894KNhGHn7E
O+xdZ2gK9/prfpW9qf213Ia+PgtAm6ex1/LASFWN3y0XN2DW8KXql3Cd2QPnW0/d
e+fxq3WCEhXknlFhOZheyx60r07gxcbTV10tYjIXtOT3MW4Bcc924MmvbH1Nq3lb
0T83pJQQDTY0jFlrxEzVF4NmLhAH+F042c6tS2/a9Hkzp2DHaHYu2oa/xq+fYFI3
4q9wFf22zxRRoNAKAtivMWUgXcZVr2VaRhQu/TIQQe2Ma4vgwuCeUnQRCNDKSdQO
mNd1SenOoR8UWHgyCipLM1HXYgVNHsYYRI5XEghY76aVpGAIWFs1HibYS0Bi0D8U
rcTDGZfPhyR9wcFtWlK25jwbDKxnr6VLvtax+4QloZ+eAPMhwQQRpP6TM1ABF1bD
xLxxGJxAmxOoGXzi6JX+ZblzQ+TJgykNDrZQ1jLcwl1dKFzsZ18w9PIu19epQfwd
56QOPJt6pYNQnys7Vta8fvyqjLGxY6Spu5nWda6O3j5K1RkqBnsJWryioX+i+E4k
moWuECzj7fgESRTd1PDkJFLqWD7ucgCsGsEHTdxlZExG4bu9TJ/MLcU4M/0E8y8t
URY1bukII7DGpzWmleTc4WYiHN+i89yS7nDUGlZdvkV5l/cIB/PGacW312a7JnGS
utpsIoKHaDcYcc4vZJlThzoMUgc7YAk6DSEptunKFfROcCW+uVS2xOrPqoUaPPY4
l6aurcPlJfbVh1L4eHAdEHn2NAGfGHTJt8NnEC3SVPCYv4Psqm1ioNIGbWT8y3u6
Dwp0mv7RlFXrt1guxDZCEoecX7iHWOpbtofJ7pkanMigW212g+CTcWwo9b0qu9Na
d/eAVzo9ZK51OrspcwMgA7TGtMsJrqTO72YzYDqgkQDz3m1zQ4kB9dvfVztRsQyC
`pragma protect end_protected
