// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
sVm6hDwk0AN1m1h5uLljIU2Y14xcHL1pP8derSsNtPCtfBVZPk6wX/5zQi5Vzc/3JA2jah5sY2Ym
K2LzyKUKOBK/Uvo3OMgX0CX3isucU6U0UGz2K/Chk+y68sovYzGkqWLva+9rxl5eFTAhrgUQ+oPR
YBPYPvJj4UAn360SdkEnTVSLkh2oqRrkBfD12guXXX2LiDS66M9j2bBN+tKw1IFUB6gp5LnTAOLD
PRBG/6cxhpV05h9+it6/cT4+EjRDqiISn+dRmZhC25LYeRFA7AOmPwbed48R43IhJ3NMKE3sMhmY
qrv4BzXAPZtC+/vpwZdfIgq9fGEN3Qc7kZMDOw==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
/rmzGmbzfapcNkNQPIk+gZ4Rdr1oM+SQqg7BnWjYSWxChZbYPPOysZEu8J/1b7dlMP8aNkXJxt5a
8RViIWs20mztJjSvSx5IXSzTggkCbRa//VqvYvDxdbQ8Pnj/mnSZ9Sn3JdyCDryh4AsK4Y/RgHnV
GMYa89kkk2KLJYRlgRmQlenxUIHzavhtWRUtg9x9bUcM1+jPnjjs8ai8YnSoHJfEVOSF2Gai4SB6
z6VTF5G3++VJiGM2H/POckdU68rm5jGpMWrjRhEA9hCM6pUVjq8h7e9C4G0LcYLfD4xUsCRXvI4k
Fr2Zw17NS9ThkEJZSDg1/cFgB1WgRZZs4YrIpkWCmd5v6KjgUGVIQ9KgyJvIIAv7hHKhbX1MAZUq
er6u2Xj/hjdg+84X5jaVEHJtUZpDF/ndyi6R/rjeR179q3FfZk1TcgujwmI3wYMzdJdxfC2ChYS3
pZ3uZchGe+ruoNnpVkfWwJhYRKmUHqB5ibFWVu+HePLHjIW5PFOHsMcqNiiHoN0JioUE3TP7rrc1
LZyHEvnaPbNwQxR9ccrLZICMLXQR1SNz/vyvB12JaozGRNC05ci1c/5Ld6c0kGbG5Qk7o092vCVk
7aJVM2pAzXZwfLdWaFgAo9IDfLhuZPsI7N/W+7vRaFLLNBIUx96AnX2N7h1cMHa19YViwll1J5xX
76d0fA+zyBKfsqODdzBUJ2OGLXXPsxMdEWkI59kGj+ev82sy8nvwRfrMGCfWm40pdOp5I+SHCVU/
I+f2VavnU7GKjRn79D9wz35vxlhrloo4dkLZisks+QDUgFJlNvSzdu0w8/ecyQptpKXOlv2VJiLJ
gnuXJ5armFIHkUAVvU8pYrV8mda18h5OvCsP9FwB3rs4dLzJX4A5RZzlx4HNU5s//AW1bWEEaK4o
vod7pNVBWK2XZb/4yplYVk+Wzff6LcJLqh97Xg6FoB5kae297URkXwdo1VxM1+8J8tL778PUH9lg
CtHao3bGesUjZKdvQwe8us+lOh6WVG8hYr6hViATfCYKJXioyC/ShvwrThfCpvkPX7GB6Yne8cPy
/ab/dLPHmMgxl8mNmVNaJUmnhNJDzDxtmPhrtRmyLtjRMsNoOvmi1t7jr38C7eWkwVHOwP/Dr1I8
+AjvRbF+5IJSMYZf+trBBd7cmtVNqBZ7f9k7SK09CvVRcI05o8OzwQd5Hfh8AC6CkC48LPGpcR0r
86V+Fw1NevB8wKic8QVdsAYBiwTCzw6yRkmT4KLVtR6iWns/cR2d/eQOmxnXjgSuwmGqn63KOCR7
0qBon8udBq+hEM2pFOKxpIFfCDmMOW88VvSqq64Vnx7G0tkCm3/muk/whl+GEoHSVFzlAGkPqVdz
LL5+bstcUhRaeXRxHz9dUPxwcHGaTE3U07GQRlGh4gU6TMxm1pkmAqCaRTwuti3Rrs6QhxuO0JKb
qLHTJye+dfZHrGXcyysrOrC4XodMs90U9IBfLX1bZ32Y8Fx45SckwP+GLVl2IcpuUoX34KT/m7rs
oSCmi4+cZkS/ZaAALl9ca2Za67aMu/5b4Zg8CuxFisV0JAv+PQghpkK9u9ScYljhtl7G/cw0cwRE
vRPuI39ROP5j9smEpC2noUawaOQ28aTmwk8NWFgdzfximqXJMtQWaftTLCU1dzF6z3CS37azubKZ
K5KKn4qvTO3UliHboKUufBiMkul7ljWFqk2f7atSv8sknEhtGG6Wq6dzL4Gv9T2sbYvZMClsl3/K
timcji5q0MxaRw63Lozrohltm88Bq7vrnEs0ndGjn2/yK0l9oSi7pENMfFrwvm3vfQtRJWTAg7f9
w83LmrsvFsZEve7sYO3NA5jNA6jaOnEycTJD7W0tMMF0ta/CuyT6ywnwWPYeZLPn+u40BNq6QNL4
tGtUk4gOcgF2Rn32aW2jthUKVixOiSCRxkZwZ1YEd56JTu1G3sc5zZgM/CS6J1w2dIXU6wAIedgy
6SQZm9sb3+PdQjd6o7sNppeLDv0TY7wEBWOKjNjSREvhnlbqHDMPX7PrDyAFfw6SKVYo576Rx/IE
cvH/KEzu0lAcrv2pUFiU5xGHu937oiUf8M9KNUH5NRW0BTqZLlOsh+ctiT6KLGVEk8lOZWCl7oJW
ZydpyRr8mOEe7TJeLPNE80P9aXbtPRGTfE4f7LYcHDSXK3DeevGvOtz9DAyBOH1hJPK9U42ixBKG
/2oFM9Mxdn0CcFUcDLGru4MY04Oiqc42xKkXaPmuHz8eOZnlwFZheF1RHlYgQy6fxDj94Ev3cEwH
juwSmHGLv6gMDhQ6KRLyiUV+zSS4he0M0Da+ind3t5o7HCb+7XpLEW9rcxWtZY4knOGezMyCsKYk
Aetbweld86NmKu755y6QWjZttXFEV61v6EAGnKJFo5DmArWKS44kEGLGdxevWwLQLbOGXaMD8Ler
ojree2ZtBMwGoxIg86vwCfWGWWam4QKM9FRun7KQDKjScFz2i+FotQy5gx62MbRMop6LXoybMTzM
m5nAOhSxb7+ymvFsT0MLr787EhS3wA2+4EhyAMtK+3xfGpYZKyOM75kvidbeSDV/BRd3ZyfScX2b
rxIbya6xYqRxWKSIv3pkOFSuViaUXSMOiEfv7ab4oneeW6zI31VkHbrs+cBT1ttcrAl/IP9OGHi0
RW0Fi/gL+jxRUO2UPsOtKrRslNi9Fr2XGfynMMSVRYkL59kk2DOqQ6PwpNw0kJ1478w4bBi8PI1G
frZzhL46sgR0KNEtzZqHvELwxVjDbS9nXH1KCbyjH6vzhgSDIb00TrtYBUa+5pwC8QyMLrzrxoeJ
kLf/2l1xN3AvOaA1PiX33PZ2ZiEOBJXDB1HSkyQh4XOt7w6efDHEY2rNT/slx3MzqF3WlPCv5mLf
0owCoM+9evzVmtrAEuARRUNgdCzsJCfmKyD6nzX82jLqvrzJMRqKlJ6WckSwyzSaFqfrEsFp20/u
fCj0+p9+VI8X3/ES4B/oZQgChOWxPGUR2kFYBQOpGLSlT+cgsAFtov0ztqm1UGlQuefrVxruVvsC
JUKzg+ANp+FbW2Ih29YalldoGrXtEAn1RNrYGyuuq0SvgwxyzfaqTfOXe/lwp69vCghE2dTbe7dZ
cw7x/ChkiSoZBPEo7tKirbyQS8DLGuzivulm5UEOguqe2whZWYb9/JlYoXxXYjTsYhR86yAA7pk7
EU7EyXFW5NYxmylQpzrv+eaVxxNCsW5cMrymUA7UStg6iU5sLJVNrHbYfDqEeRs7zWAmH6+Yzbkb
VzIpOWWPgBrZS/KKV64s1mysLB2FsR/UJnctcWwL+stAJmlpmeoUQET96PzE3xbfuvo5U5cegJSe
FBfTnPaNFcBmNAhRcC3ysvEo+XTSvKQrKrIMjKpp1fGNCchd2jUbCMp3xYmLTmEXyF3BGveGGDtR
Q7NpyPTKMV+vgvxMMWbTTDHvsbbIZ6jd0EpeHOpT1SpKemQcUhChquSLqCVSLKB4tzYfoS5s9iHN
4vpHMrWUiEfKT3lgw9p8i6J8y36ZywVzTDhIk8kee0D/ofyaz85zhCgbyUB7kMIQVYylQOHUUMsj
GGKHslP/mgfyZyfOqkioVhd+M2RdR71Lepjak8Nr8L04weAF2jpiHR9mL1WAkVQmjF73UhqX1E44
PCLXOGhdMBh6qlg1JXI25ZmqSZ1sT/6vAJjNBdtPvNQdLQx2lTq5BUejJwRsmrIF5BlRUQ/mgMPU
PdDakE/b9sj05gADFi0KNiHtVf2UatO5x3gXqCX6HDyGQhlVUdtFchFu34v8lcykic3G7mvJnopz
LJDRWhQDb5TThCuuDUS0Y6aSneDUcGDAsY6HiXIOYXZlbnxh+D3vPLhB9QeZp2CafWh434pc5s+f
9Wc7YRu/yD15eLMfxwxHq2Uhz0bY7W7EVJPGIwLL9o67yczTL0t83VqyXCG4tvBXwACRFa+ouHo3
r2c4qlKjhsi9XxJTZf0mEiW/goyAfe/p8BGZ4A18Ojx0dnbGSS51zjxT+KFIDJ0MMyryaNw5A3q6
gK3lbW2NDHpyhkrU74YX+JSxN0wZLj1rvff/+T4qDof8G4MwBeFCgaNITqiCFgv/D+geqJKhKk6K
lt5imOxaI+XO8+qQQIZ0wst1cXLtR8IVuzSOuXTCIkP4oRznajseba1IES1gtXr6pFQ58P23pd5e
OW5gLZ0PFzZbJlSJWmoHhczHtLOoyxRmUOqALa/7d73uh4fUd8QEbMTJ1XHstFLjX4Jq8R32wons
NzoQpn3GFUIwGCZ4Le2n8k1PWO9KeESjKtBdDKeQ3lyUYrxh0lqUhG5WUTh62FnYGirxnC1WsBDc
/ABF2GoU16y3Er/u1E9Qny2HxdIR5jFa1wSYO34Gkf8XS9lfFEvmL3jbkNY66iboYlMk4AI4RMqK
RlFoZg4GNR0C6aOUEGXEGS13w+EmUAUtiO4dYfbdRojsgsCXyAmiO+dd+SIJraoRmkdZUeu4yqxD
jkJaI8T1CJ11zHiSXflreqzz4l9dI4AToPYdY7oe0+8OZJp+KiW2GPrsNi+bPXr/u89Lgcr7AQiX
EfXr9+i/6ct7fdyXgA9HqZSZ2mQdom1S+L/N/TmYpNnPKM8fQZi48YcNyOpdUKcOW5tKQTTEBASL
NMODwBvHNizBoMktfhNktGiAXwSIlWuG1I1kWFM5+CAwPdfm/NWzvICoa4Wr/L9qHFKTx47YTw51
kHk9BPh5IFcwaHxVf0Jhr0w+TE3E8r+NF30J1GEpFr8tX48TZ6HKfpcr6psgXsJabo96C3xMSlUr
sGgEZgUXrtcMGWMb8wBDwY8ClVoK+F0zNi33ZZ3k3eSeetrvjm+fm4nTI2/KPbHXHF0+h/oONsPt
7UPbjn8BAbWMexNq4sxvHqSSNRFnWIUgw1/CLoEUSKOhObkljDP9IENTpANaHRjzfQS1RQWV9VIk
o88eMBUwWD41fua/PpNqLP0VUYiPaUsvyl/2mlkpNxXPEzNa/8YKFIpBXtZBgX62mxuN+zQi96Tb
qEwwclW5imLRvrUMX53yaVFyIN1TkVcRRSxDhWLWEy5U45J1jN+oXS5SHoeYcpLbBz+GClu5sWzC
1mDUIu5hVyGtJ0wItNrBXNV8ZCVpsrBUJtFbGoURwTNtYjoUo7UoNeYUMvm0wFkQQ2Z096KcBr7/
n/ZsPzTOkbgm1hrf0P3iYBSOFmxDAGmQveU9mSAX5SFvEdh6Or+5r6k6SvQAlGLl+w/JHg9ZWuft
i4by0cydCgAgQvgMl6AkMJgRtWrBSwW3sqct9PkY80UuKBDdv1n7uZ49rTHyT+O7MtozaKQ+OivO
f7vTUoVVHfoTCwvza5GLQAI5PaoOY4f2V4aRX8C2uuc6CxglQtnN/G+qJfX8ODSyPbbLjcI3ruH6
v2oVlL0pL3cEVZLEg974YWTLh4S+7ZDlvQakAzcp5lGwhRH8dBMx/nVGg5bJqoArXSYRNIzELVea
7SgFBQ2FBnncPQE1l0DAdi6w/ckkboUalh07aFTTW4jV9KwPmqUXqKwr2akS+aDc5SobolOgfYEw
JIFNdxUKECf3Nr8Tfhikx6MCflDoQyRRjbzl4Lnv7dfvRgUSfLmudglWbTVLioQJkgdxD0V//t9O
maWKveLgPKg7SwbK5yypxuAraVyI+0JSliG7cTBMvryfeqLGj7bZppTmFyXq3lcqWIsvXRGyAfuK
oTueimYFnTw6DcclmCXwrPiCbub/LrLjhgEYmIefNMxzG6MQPav9XJlt96vQeZEKZTZH+Sw80JRu
3dSZL2HPkuVxqI8MqjxlSuoIumMN4l8+gq0/n6pFumzSw/m8VGrtv8W8FiA9fhWiwiwvDM+tx330
1yN1BxrItackGf6W09LtoPmQHRImKHKLmO5Y+wbh7yGxlY4ngwsiCbIH8+ulJoVwRG2uZeuAAR0o
CrQ2q4N0k9Uf+L7keLH/81c9VNJbp95XZIzCmt5V2A55e3oPTibjtTAxqaTWTIwn0CiAU/k4+pVE
Xo4xq6gvPFzWCt++M5rGKDNf6c6MTxQxMcSGYJS3WRZtVtdlyYZZ3NajgeC28jRK5fwoB5lELgLZ
qxTtD6TqH54qjuwFtKVXrO69LV941OC1gL2VIGtJC++wmQ+wcLbaE9T0J8FByR0yDUm93wl12aBN
lHaFgSmBp15d0h2OR05W6XNRWxLnH4DXZ7ggtXaqoxrXulho+qxz4DKJYBQtESK2bW0hoHFQ3mlT
j9QjKPNQzPbrIrtrEPNO5MLxG6lnSAodD0Iadsp/YNYI2EQb4GDWqOF1R3tqr0LaIFcEVSgTXeeZ
0DABai/dwmp8xhghm12NugO5ytLcAfRk8tGNKdgjM+Z/FAuLyHuy/fXIrIAHx395WvLyzbtkfWMa
tRuOTTN9pk/6NX66Xvq5n74kXGKaU+Rjjy/aHW9vvT+0HsZJVagvH1BErkVkWuGxASwrykEyDfjv
vy3OHaNa9tbCnAr8QPu09Yuqle4sCH4klIDO95HvYscopvuff4E7hkfr15kkZW65Kli5Zbk2zSzt
WXG+m365ifGqjx3J9B552GF2T/xnIQt74mSA06FQcpglRs3mCMS5Cd+9aBdAhEDT+eS+27VoKRiq
ztGL2aikZG/7itLluGMYwAnj0A1xKux6fv5aJE20uOcAJPrlMRShltX4cqIaTl0LwROzMzrtl0ke
gmbFdJ8sDZkqdsl/IxlRgjSgWwroWHIv1ms6nYiYVAXhWWT1jSLfNuA0MwoQ7irWGJIr8gKYiCdQ
AGUA3iTm+ryIIndhqo+Pog+00GBOxfDcRU3L/DG5PoD2Nvg3jMtZSmsSempTPTqBbZPjkWs29cAC
WIdEplzGAvRQDOirm2jTva0R/ld3Q+LZXPDp/ErSQEm6US6TAsgiIrAc/kycOsMvSh1vopZ/N5Sg
wCRRjVajxEpXKmiMLNi8f9nqJ4mTKYjof1L1t2D+dv8F29ioc6G4/Xx3qwXX2bWfa5J21rEAYDqZ
fQL3hy4GTh9AbS3R6kQqfjF/A3hQJhB1qeDo2PlI9/TLSRQ52ubSpQxwfeRwKLESCcEKFBR+SzoV
RzPwJel7O4+kRW6CUHPkP0aYQnLQPbwutCThzumda9aEwm0luYlGp4QK0lAGFVcQ9pA/HM165OVJ
EHjQ9Cy0iKY1zyNxmXbA1Ce1+QA4HU3luwOC8vbHmzyqhA3RHtz0h9v1NxNM1OzhMa1qweF69mGH
u+WrOLmbMLJP8GA+asN9i4dQ5MEFGxUX8RR2dQP7tCpyItDHCyZARW1h8od/0pBv5W9WvlmcnOif
onOqjt5+1ihps8GOJ83eC6FFXNA2oyIJ+kVV/3U2rJBrqiHBIhOTvwfYFOsgc7KRNRD8EKYQqIzU
EgaxId8zvk4/6PMeSxEDAZBdXEd32S6c1yc8rtrg4t+WM75LNdkkmh53XMqqjyFMFvvQEudSDPYF
6k3NKDIsGvARe2m7LUNbssIMSRIujStxKBQaYU4UAoJHu4Z3PssdJbmAnSVVvlbdrMBKyRFEKqcD
XBpWt53CRjTH5JNU1Tb1mxvzUd19k/8yil/FTf7fDGPCv+4rzZZZLivZkp7IPgREUIOGAcvjPaZb
MhtXWxt3LjS6gr6C6+PDLzz5DB8yruZxtm6G913w2hcmFX+km1r/uvkoNlMBPJR378AymSvABY9a
iYPFUdOAQlDXaERAYzhqp7G4WUPfWVp7vmxwOsPEBca/1kfAsVxCH01fY/6cjVnp1AsheY47g+rT
StwMFst0ooccI53Qm6dP2dpTGZrAWHCdTLuTVaajC/M1xp2GhtCYFEz1j2iJ7sWpXizZ2O0g3Q42
YLfpK2eDAAtHqCr3op/IrP+0mE0qYKIoaqQathgk25PT7fTEkB2dO2VA3scrKctIuEtEnTHKNlEm
WAMnTPIkd4OZfr8c3RItyHCsr7HOrq1orpCdQpqpOeQlv2V2OfpKrtFg3tQkOp4EeYiTuRluj7JS
WlTKq4k+i7y9J4IDr6DCQbYB/LEErMVCGa/aXFsHtYb6Tt4k2kpOfwmFfIrRu3gPvgSneRa6g+6A
UueLVCc8fQyqld5iCktuNes3DjpxX6AqFxGiIg9p5lFe5hMGgqJESwc8cdBaTSHjcZ/qy7qq2PNL
GYXP30zRiwCjmuGuU1T1ATaHoLi0LIsvxuj0ymwATX1yKQY9oQJy9vpmzbO6mpMqDazPdRNIRO4o
b10QP/a2NIEgZ9O63ooS2Inhd3GzSXc6GCnpbpwPVD8aDL5URzc3m/TMVjbtqjMg8e0wGLy2YYCz
Z6uugnvZ43d0q+HZk/RjpCnU4t/pURFlTvA7YviGSh3kC5UJ69hIpJsILhMb5zn7sZRmkoPekaCt
Wme7xvlTIlb14zhSJmKz2ENlWnOBp367ztw97LESGr8Em8qrVFgcBfCcsnxwy4ButGQM5jJ4PN9V
1MAaRk0Hom047b3laDNL2TFUf3WGvMpMLeWpuSdFmeifzVid62l+Hx1BSlj/T6+qF1QD2cL/WEU6
R6bYw2DOfQAYy4Uqm4Qpl5Ir15dA3NGkbZ3ByI++FtUfnrVGgUWyrpo9R1ZW+6BZYQroN/La1VL5
PSeXI6rnzp1ZmyapEKV7DWOh6UeVSh5uAPougV8/FhtiypBGAuDFXoh+7bP1+K3jFI8Ribp3UXfp
lksflpBP0DzxFjF6UBC23T3hN17cwyiuPp1rmj4X0VoE9QYednYW9iCzXNbL6h/m3TLKoLf96htI
8yXDiWBxGM53sBwD0LlansaixtsjnMo+lhIUMXlokDAox/qBTSmWm9B9cvrbdFRK2WRgU9/bScjK
p19Q2h9WCNaLnJCa+Kf5FCcTZ1nLTQZtuKbZ9c86QH+muCyhy/6r9EqFGBylBMyani8zqzfJXTlY
orXtEUy4KkV6r+DO4bYQonw9esm0/YsHK5rMDoHnVdoNMgEOTyEFFSrTqQ+K/2CveJIJTCuLBakP
GlLyZD4xldpVMImmAjYkOv7pUd4z3Xm7TWCQ0QKOBSV+76tywWhOOBVCfJhEhrkSdjoiFs+hB2q8
hMTdaC9TMUwyEYjCCzwI5O160B/aU1TKx28xivR3L1FJjj68FDY1mp1eaKUnnCrpjstobQ4pCc2f
UTJRrBTRI9AiDSiA140bwDajA1MkzhBkULOz1LsHkPgZ09JinuO6RDukjqN93s+XeboLpMRUB9KS
Ja4jIqAnZngJzbfvwji9/YD7mpaNIhdYnKAzEgJpnwjZ7YJQ+e8vBGcrHM9Uo92mxI1FOTbqPwZm
FxjuKo1UlRHUg/cbvIACHdfI83gTNgCUeaHVH6oIfI2qBllAacBGxUU2SJ68ew9cqXZYdnqDUQLI
TX+ZMwXvvqq4PXvuQqIr0SamFERVPwjJV7wrDrjZuOmqT7bGC0NZQvOPIM2XYNeVlqegKKch5/uf
kK3e4Ccsls3GoFnAm+tpbSQXgOZsyuGNIsdpJzIx/hFkH2d6PolQl6ASK3icSQXyxELIaZkesvFe
s6La1IQlwynsYyWJB4o9clJAHaKCGQ9GDs02GiwtCK/9v2wpeT7pXpTtPGBQyLdpcXCoE9uQzuVQ
ne/U+i1dnNbLJiX0ZCFaewPAv5f8X6ctQwT2ibzHfKE6+S99nmUoQSwxPUAxhYlI/XysxIltuXma
8jQaq6308O9T3o62OrmCUy8Zil2eQWyeDbmiBpb6RK5lK1V6PxYlLrvgo9gBV/7hqeFtSItR2mVh
Bma1RLBBGd65+64OKbTfsHfScpjty4E/5LBksokBGwpnspTWWnQxBYqOMcGIUJ8ilKMoQ0FAQdt5
avZ2CDJxgaQpGLrXpyBD8QFSOqGVJUwoCNEmPOAGHeLcHItiR8xGryNy5TOZi6YcJ5jkF5VCyC+d
gAp0kzEZz/VuTI/x91CD3Bcq+6bN5J8C4TChKdz8ic9FnYzNTzEm618unAt2eXcehhIaLRG3rJBe
hIxiKSGFdnHW9wPHpJv0WeQcc/+zA9TOZF5nKsISTDzVbJUcYe2T58SjulS7pMgxpJzPi37irSXX
f3tciUZNFKago0pgNyU/c1lo/qspiptrcGlJUyEisRUH3Ed5WGCicL5PjM+c1bRmfPmzBeYtDscV
Eyt9e8KzSmItq+zNBjccykqjK4k4JisK4KTTq4Iu0zzj/36oLIPuv2qrtF6gelYAXaHJQvLtwlFw
6EOo8UOuyxwegrbOc0TrBhLi6pQ2l9l24RYN+05bVaakaNkMpJyVl8rzGUBs47AM7xb/OVBdRLpa
lmP0Fvd8SJEu5NaxD+q7VWdHTk0okQM+yGWyd87ustaUuxpHAAd3wAjMBi2AE91EiMg8eFp7fz7P
kNxQA2gZQ+5w/YjHY71ZNUHcv6tTFeAWDWUZe+5Jk93olT8M0/b8OCiF/BnxtPuNzcSQ8k0FWiDc
3ekCsfmiZSeBdkFR8Y/Lu+Znavy1uTJ7Hs3qdIDeJQHXhIaXOAfV3F20us/RK6zwKpUAHv2TLR6d
q8LrR2D6z5TuzHTLP7xf1tH1VNObNDdQH+4JtzQXLpCqBnZ2uyO7KI1T4rDKeojEsLeY4A02Vzjg
Jl3H/vDDZGK+nuMFazmpDDhKtZXLi74SNzVWmABy8NhrxPY63yMQS/HT+mp2I/Vtox+ySkde27H+
Pjn4ohBMI9pI+sv1nh61Z8kAhOCJjhuKopBjSPSywbhWHN45oVC5Xzve06lRL8x7uGlPdsapcOt9
1zrXsWdgb9VjSW05uwLklsUn1crbw2Xry0qld0+eV3oL/cAd6bWq0RdQd8wFmqu7K7Gj/DlgnNQW
7t1HhvnFfEj+CDv+ls/Ufre7bUio7nrWPiu+39S+HDSAzpx/J5dkahkdk1kMcct8vIT2M4MXdrIf
QxoWxtk08O5jalEiDimhMM5lMzCxwQqtNcf1w8AfUi/24rMhr0McChfFJScNX2uC0tI773I+y8wW
MuReIa1ZFMnTo2FXcFwo5BJftOTXpDpY1mhQP5rbCSuFfaBGa3Is/OX6/Ck5KCk0Tp1AkPu0GmBB
nP8xdVLkON0bkrgoUYlRFWvmLLZP3UCZPmH0TSM+15dDAkHLtGKTHC/kSUvH7Bv912UraOLHkndH
tzrfxPIREKjphOwy4qswS3iwBZ6bLdfl2cQScA3ylsh58vcU+HMwI9rLU5P59UTntn+tmmsvuB08
vR8Xkxp4bOcThcBTlJO05UJzV4SwYFYcvM1zLMCzs75rgl2ECOrOsWPuKOeFG45rif/sAHkWzQFv
3hT4n6SpsGv6/wooxZhOdH+LTYFSSZ5O2f4cMJ2Eh6x+C5BtCirp5CrfYIyjgIPWJxqRsnOIBaVw
N+26GDceJJp5yrNEW4MBZbyOtmjYkAwkzhU4daNP//4mvjNqeCq2C14SAl4toNzhXuUmnPjnBXr7
An8phx7vE3AvYUXFJR63iJILTmqOqDLk3sRnPx8RNFjJ/l4IKChQhDYXluvLbR4DqsfZ7J98ZNyJ
Q3hGD1YNQRa/oAU9ZUB5wAw7FW9hZGJJKH7FTBoGy50Wu3fBGprpOk9PiJb+d5lxtQiZYtwf1C27
NZSmQz5ptpeLPOXziDIGKK5pwlNVUoMkr5MdNPakTuTu2pnqnP1AYLD5mKk2z54X3VkOrRk+OQSU
mtOS+p6wAy38xHoO/48T/p8U6jgFy+hrRYWUpvb/vialuvXckvg50PLrYBn9Kum1kEIWNPTTKzkk
70/x1LcuXjHkcNl9I91uOvF4dzKvoMAqU7vxP9xFPZ7m2BtLxHYpylwCDmVXR943TMAVFukXGEda
CrIW1dWpo59Z1EbXGL54qDKkbVfTKHEsH48UdOG56fCsyidGMWBWmncLIdW7IlwTS6DUSFRSugDh
NJYUBHyhIsRpfcRi+Y+ZSjUHpoAMLCcYiDqzDtQeTTECOObzB0CyQKxIHzmJLS6PKV2csIGbbNHg
5dxKWv/pitX0bkgKsdvSvgf/Q/spcPIViFunvLYkC8fg1ogTusdFc+R7IwzdBBktG6xwKA+dY/Ga
bfD5CQjblfN9b4LEokHjgGxJLNfLU1XtViIi2aXmj/o0YBFRCj+b+eJcSg1s2YbX/iIxb60ol3Gw
w4/esbNWYdcvpOkh7mw7ibXuX/5HvLK6nE1TM+0gUmMM684T6wdznDugMYS2aqyhaEtazHUOOmUa
j8UcLpkyxP9G6y2m1gBSoCB9cim6898CVY2WE99frY0x3C4iiNIyHXJ+hJ92KVrsLqr4Is1M9tZJ
xcB9N86ffAcZpvs31fUYUU1rmOBtFZsRnI3XapYjfKrzrGYz+cvXTRvXtfkOsF9+EkRAGewLMFwP
L3qDPBhgoMPmsGUju1KpmpArP4m/Yso/DuC8IzjIPnmGbyJB43cbIXJBsD87ahGBPyR3n9HjPgva
x/LuuDdJzoKO5/X6p2tocrf4ThGXXo568YwICzxObdraAoubjEO9XkhSIivcokR5MNjnyS39h6cY
e1IrM5TRBeD0AbsP+jdlj+kMjt1cEA+uhHkAFwm60ghgrgjU9vCSNJsyYySmiOMBFk/6Lc1d10ks
jjlgKE+fqgArxN76PwwPowHhVAik6uXcFflAZ3oia4QDBvNlOvY0aJqJeUoZCSbBtgAyPiPix9sz
mB5T4MCW47cAdY1bMW3atzQQh1Q3cIhCUL0iAxrB3VSvBedCbH9uuc9xbvvQpxJdZAYHbbrX1BVJ
UWBDXD2ZnoVu0pr97Qp6L7oQjOKNdwy9WK4pM6yRBJRGjk1iL3nhXB8l7shnRBy/nor4SedwTAfG
Ll/SK14t+omB0/CHaFd/P/4eh/xWVFwoEwDQZ+uKBM9VT5mOR/8uVZ8ct3GsECrAxlFNvC8gzjI0
zPTbssCzIsxU7DSe5ix/LO2VQjbFapKB1EZMKT3S7WHDROCQc8DNvRBRNZfZBw3dODngyJMFS69j
1g6Auk1B8JBhS9hvCPEXV0irGeL6Mq4H1i/hgMh7bVOkmVpAE/tVnBpEMXGjERG8UbbYmsSwBZ37
JCyfXsQk8t/6d36PBr1pN/NQVR0Veh5LXSzJ8ShjHr9wPHVH1Zy5Owi0I5LnSlzBocml7p4Y/qgf
mJi9Izii6iM+Khg9LPeLOuxO0wWQ9FVqAHmsjS8U6l7Zep3fkH39jIr7ww3t6aSBDZzfmP5F3Tir
6e29dAAtUt8y71juo+/IQwwKmhLqJx1abATuTYoLxTJzifQB+lhLSb6JFOReg9ssLjgVKLGYBAuR
4qubGRAExJqt3cee4huCNXP3qbmSii/ysKbjIqs+pAhdg6w/HoO4gmP2H37rKhG9JX+uFDIAijMg
LTcD44IHdx1QPcP/CJLvdotdeHyycK1XT5j3nZfaltw0bgcXhe+HouHOBbm1SVLZHe5GUjxkzqmR
F2flH5ZEv4BgLRsyRcBJC+5A64xes9YsTttx7O8KG60fSmF3ib8Mej1wKmfSziK2pCdIsMlGKNoy
Bv9li3wKsqCSP6HcPqBpU4H4+Dd8v5YENo2gr2Dkr6AmaLEmhgWunizHHoj/ewgy4/Vj6QCW0KJR
8NPe+7FpgtNDu69kvcXbTfP78eK21m5P5goA55BsCXGv8ufYRaH5S1aeSDl1VYPsLZu2YDX+NaWT
sqFDqWwQbWkTQ2sWFlgTPP8f3bTwgoXBd6mNg3h5J2+3lZsyG3fVgd1BXMjQXSG1v8DbpEW6B9Ev
a/f8nbkk5VxsMNO0/ZaZ/lrIuwi6U/F+REpc9A7PSquqDPUSsR42QSzRDpd053scCu0gxKs7g/S1
OIxN+7mZ/IaQ5FxS+KhoevwqrPj7sht49s5jAIPuLWjHCROGuJGcQKP9cjyNa5eq646Ft69qwLxp
r2IW9irUUGRrkoRyBDmu5LtwkLBwpbncd/6E7+1NmvW60ZQ2nNiDy865Y8MrsJadU+34f4lWL7LT
euSFgLtVVpS4U6zawm9WdWDEPMAQiGzJzWg6cysO10vOy+rZSz/XggPWl/8hz2EJ0wexhexEMSRI
cBQEcXEzNDf8H8HnbsLBCMd96uDBSLBn0hLHWN7zFCK76JNKbxaClhAfio67A0RotbavYI+0wVoh
+JCh/hzCz6cd6uYNfplTczFBjFawit4iFcAVw0Sg6iqVyD0JxEcKWzQf7InBGGAPj3Z44IP4b30z
bpdw7Srue9IaD2V+va3LRY/NE6kIgDa+WWhK4mBl7VjPiCNrNxRq+9ELuMargEw36/wAzYCtBgrY
TG7Ote/DraCxOVJicOd4CWN59D19nh9qW3hsWbLGobq+lyEPJqTN8X0ggI0GdA98N2dlIs+2yl49
OSu4pd99ARmdGoCPS/Vzh5stDy9kqE71rqY8BK0BZ/RQeW3OidqC6PWMokVm54NGm38iJk2wCVe2
eWopf+DN2Z+2B9bLF1OADiPy6tTXjaMc6XiYlSVg6pF6jjsVnFltYRIx2bWUNGfzlY1WcjPXESi5
tbU3zA6sCnIDquU9ub8x8s2XyywOJiryo3hfnFn0dpieRZw14UgMbHQDRYzPmInWO6YEVAWe0foC
0GbevUpwQarmNXTnRuX6Y7bkKYL8wE0Wa2I8V7HYtxp1FYBXwcIAEacC99mxFm26DkcK3CUfsOuP
WjH/DC/zcoXYsCLw6KlQ3zbYjuZ/+Krx7kptP4Jt2pGRktHA7QSQ53k+nl16iNn/+/CIXxaB8Hdh
BEtYWG4TswVmt4qDyOeJOtr977hmlFnSBQLmtwVXFDR0cNSTQf0XzIAlaBOWCjLStoGVCUe0xCtN
sQxNSbCtw3NVYmFCgsCMoUT0w1wsFlbpVYESLemDMjOqLu9fft+ILxWafCzJGhoMF2P0J+eiJthr
H7Fk44e5F3Ltp6L2VG4IhpH2TM1hQHhjTMl00XbJvlufYT/rWoL0njKulzPyb+THnggekGA5gZdb
/8DuA5t1X5Mnn9NUjjUgZhWwRg4JJRfCL/zy1bdZ/8eooS9NAiNyN/m02JmLbBxfzT7/dw3ZA9kn
0Qh5j34gKTliW9jwWqAYkX+vQOtDL3rpPYY/ik1K6rck+kqr9oSBA6xAgQirRntUTs236xI4NcKA
Ze3aA9InotgDuv5TEHfQjBSMqHtvc63V5DlRUNO711v54S6BZFNDaVMQvbN6qTkUxcjslfxuqlVI
NcH/bG1uE6+cGKKT8FHlqPcXmvwc40tQAWTWAg7TJEzmH+P0vc9Dc9B0z/zrQcPr8J3BAVYlPH5o
BEvb6+tVofDrEcxGXkreClAejsXvbrxA3T/3CllxdtgnEOu+0k10KSm40Wf4noDmYHhEw6KM6ptv
qlbuUi5RbF35MxL/zALvdUiGKstnZ16gzLboND0wQzulfmSisLX/9LbqH2mxR1t7vNVh21YHmTQQ
xZUgm+DtSNX0dfQzbDFko8+BgTOhMPMMezCAwlR3R7NtBdx1VfzI/Y6dZ0OgfBMcn0zyQxCXrjjj
UekOvvXv4M3CzaDGSzFs5PgmJ6vIs+4HIJORBJ4WTFTmKa7ows7WNNG54bm+CSXd1GppKutieQmB
KM43jc/nxAH+N3mtXkty0lGJxiLUehr9eRvWLk5qEQLwGbPLQE6Qy/VM6Lwk2O3Vy3KBPkzQNGSC
zwA3gekrGoXpGezI//3e8ksqvGoAMACysEVDMoYBAHwbftZqlO5WoaFkNRp9M/6f9zFVkGt+VOaC
8aj960tYDNQByp76jAyUyIKoZ/HKhZw+JXvYpVAbGrlpFAJuWidE2zpst+FEdG330ylgxBUeR7gL
egpVsKg/Eb3+OcNy2EIYRXOCZvR7lZv6Jnh+4RZSdgO9CZrPl5xW3+ajQJHvlup3/z0BsgrW4xh7
JSUFmKjBlVzFIYmGIs37TS1cHpPRg9MjNwiRrjIUYObZ37oVxmmJuNowmMO6L6CJU7OESCRMWKBD
XFifeSAezIiK3/Tu7eLyM56GsoSB9ZeaDZsNO5eYthQCdF8zoMt4TuBba6jruWBEJBGEtrPeFzbx
h9dmCEd+KdoJMQSDzKH+A4In1dGfkqQu5CadvxN19mQc7mDB5SLAGYNxDjwh+l4xIrHYFftNbc10
HGUd98ehTSVWq0BI8kPVk14++Th+UzcRX3aH+VziucEbRdWTOtUHP+gtsthq+UMZ3yPtfgOOLU8h
7sF65+eWAn8LeDqiOIdFv5FVYC3NPKD6rGBRaw3X481MapVRpVwPSXJ7Ik+GooIM1VFnUxDaJhmo
t+HeY1V27qtMYmsIFx7vOrfRsX9rQZTGbH5Uo4VuF92kCcgpx+w//my8OAh9Vap6x00ae9z4Lcds
/ojYObsp0/Euf0M+cK0xxl7ycCKHLuPfO85ukD1zFqNXVPr5wKMdThhm4s3+zeRk02glPkTxrwUd
lGOx6+2Z1wyEarwavkk05XwR7o4Rdo9hKh6sQhTEaAQ++Qc+fs2yzuZKFxHPpqa8yvDepw5xDBbA
m9SJi0dxhES5wsIM3yNUK9AZ2v/yYySEEvyDOoW4/h/pKrpcVAP3OwdEE5DppeBVAyMmlKWNvnU+
24wus4+wnQDMzAQFsJJIxDSJGoEqtRZS1VlMC4eGEkqaShErk89S+aFbMJdYrRmKejsSByNZKxB3
rA/4W94FKQ5q2cud+2LWBlgmwRJ+b7UFOdRRpSAqLUyFK8mBlFaW9ATOd9NiiB9C8i3FdI8colAR
Eh3hHS7rrb1GQjd/c9bsN7bli3rIyYF4ZfRM5I8Kd9RPcfphxSjKWijO3H0Xc1e8KXZgrYD3+lzJ
xZH+qZO63+AzBDBXfqs70ohUAX9AEcv3iGqlWLrPHllg2ci0qn87PpVrvMQMAgraePOi5NN8p28l
nqVKXpl/6wtxOkFhzNBkZaR+uPkUh01aygmL+jAN9nnsnhCIRYRcfpiub7/kl3x+aNaRZYcqdl5B
gSGDbIKt1zNgW8LpTyWSKObAVpkBdh0siF/3E3cz1zJFxLVPjbJ8P/V8zPmDyyNr0yoxS8HkYdDz
KtQ0rpWb45iEMKMtJdjyTlENTUTbTGeqUpBVJSAWTjao83311lQJtosdXfVtHeMjHTIGrcfVQfeG
B9D/ydGV8yTI6YuhlXKva6v5S05C+/FOVI7NJFvM4bpgTAxb3nlqg9G3AFdsy3aWuAopqVM9WMq2
STUyQS4ZD453p8mcjqGFX2fzhX/rMn66QmRAAuLf2UVupc9c3ZbbLP+LqlfDR/fuIqQKLicU4wIl
E/eaGUx+kjg/MecpChCHuNXEu3+2cxtqe9k87XfA26w9GxAJtmuNcncgyEAi+gJz/0DjkqNWzZPE
cbvFyGTvPQpGh/sK8HGNjMF5F3OfVbCPEIRgbIxQDv/Ep0myuo/DFvZ/KxJwFRIcWlmr8CQrDMzi
8sGmqV4EkWXwixVvVf/o9FKr45xS3cLp92Fku0OzuAXkl+r83bO8gusagnZa2nM5XqVzlcQUw4g/
7UDkwLw4M2ok7XtKlZv65SOk8h9gtRZzaMzAsw6TAWMwXmIT577EMLPPoU3aOV9hosD1YMENqsSE
sEHRlEVMuEn6jJzxALGi/1JTL0tB6Bqy8zRBXG762xUZh4AXAgHX/oUVZidD3QRNMBBM5yNoA5ag
uwfwOaYsZN4RkYAjVHeaoqFkBsKxGPOBM2PY7Jx7elfE7vxGqZ8xe5QFx0GeG6UxvDdaOSIuGy3r
F2PJCv5piD2sJVD3gnsCeVFB5nTOr+GEiYUiQpImShcTEuNRDVYnuGaP0PtSpg5CgXApLWqTM/9P
TNA5BCqvbVSwRm1sYhSI9qWqehYScACtZSkSwfv99mSfq3AongaMENAoWPVfQzokHtUBxU2AQr2X
Bu1z4H29pi48MYXBDPL5ZI9fj2AZMWWbPuLZT+h7Pj2D6KP+vyxnWBOorLNxBaTxAnh/opk4Ou6Z
F2yO4ohikS3pxOGPWhbd/nUQbOneJUMyk4RielwVVtcDMA2M7pOZAxaB15hCgNXG9L++RHa5K7NR
C+ei4Q7hGTR1SJMzH1btGs8Mt/9BMycM7NWU0gWM2siKgqjuWqmaPVN5shcsh5WjKT3fJbpivJOd
J2LNIFtQKG2APVwSroA1IkkLF99ixnujDHPp1v8Qvmaynnd6wVk5ybSs9ZZJ5J3Po+CR0bb/eK4h
4c6lp0ptzrV2+WjlTu06sDs10LbxXb6Z632OKabSmjLszdFKfN5fMsSZ0VelJPTLHY38lYKB8IQ8
Z7Jx9PphEMzXwOtN5BvofSif4JjTU40L0w/zKFYhVFdxgUPnNqeWkxekNYLIGfsQfcPcoUKsXdDx
VtATCDHkPK7TTPkA9vc1TkfhSqpiwS0nMtnJCSoVfBsnj08W6RmKlvNLRw7GFrQPtKzN2afX9vId
IfdmYlSsTHtGFCvoICF7ERsxu0KIYJDEFBzqPsgvokGuKxZCNVn4d+uLSgXgv99dFxsePwWeCC3Q
Z88ZdrvZ48jAvRXvpYUSw+yEbHBHw1X7kKA1o3hEwfvKkXiQ5XZg+TAlKrACZJVKrBzXYUovzvB8
Cka+bXUQaT9ISv7H3idE4JI6IdP5MRJzb1ctQ3APZc/+cVyyHD7z2EhFrs8/tRGIEIK3OLHlLAsp
T32db8cQonqiL7Zk26a9v0IjIQlJetN4sY8CHtW8V19y45ujr/6VfctEqvx2yetSxS9aex0bkU4c
EBXw/joLMdcnFwkwqMyJnPvmeL5ynjxWx6966G3mHO2PDCz3pr9wxnEnkAuDvRORmEUQ0OpQ8f5y
KgcO9hxA58WjtUNGP0EBb1WrL5nDjmTob5HOexxOWPkq3tNig1mzwFqQ0KGveZPgRDJpkq9PQP/F
8tUinRghGWRhnSjD3rxa13VGVsYxXzBCcTI1Qfp/wkPYtlj/WoVtKr93+syOa+s9bLDLkRI3gWh9
N7FGH4NIBtwFw1DQaLmGAMeM1++/AcJDN38BjQXvTOnnH+YL/saUehBTzfSAnl5kZe2tuKpaRy7O
YuEOysrAZDZ0JZy32wzjYHOOeUp2WAJZyCNE7qNiw2sJN+Ft6Dmu5B1oRDahIn2CAZCiGPoUAA0E
DqJwEGBFkvgUV4SqlySd92YFAK+3R33T6aRC89EyULKdegp4VFHFgRbSiZWPUMgLaDVnSAc1GlK2
quTYNu867mPuA+tcu6rl0o+7nNpJEMGhItX2vasoZQymqttmXTszMhah+G/4ojWW8Oslc1wqwpr5
zjgIAfSPFugXvnoMIIpJIL27lx7vIC8RzapqTajRyVLqTwm+QGUA+jb7dmiLlbfCchLojQko2p3H
Q1aFxUGRQ0mNLX/C1wVYUHI30At8pjOFU5EnbVr208It4Co5nT2c4LztjxE3TKT8Of+itzR/h5uo
PjFCFpyN0S6gPmWOrCSvA9UKL7LYXd1YFb1F6d4lfu4WOoqT6PBCbkAz1MMh1hum164vxxj3fNaV
r26gojb3Uy2FBL0XTNyHzYgZ9x4TyoB2Omh2EtABn1ZrNovxaC7Sn34m/w9seZyYM5WPABfBaUpT
WgOgfMPLMlcD9A+MTbMHUCEKAXSPYJEdGKoh3wG2BtoHol47wwIDNQJ+MsMmVJgjcKOtMvQUBfaq
kkfGSbXRssqaqQ9EDhPivuQletGaWJj2fGBjjfmIA28sBpszsUKvJPiPmSgtikti7gLjJWqjC3Uf
uFhgtqVQJ0/2rF/Sttdsl8nQMilKkRixbHCwUp3dq+8e5n9smIGKwKV8KhwEJtse0tetn29qzY8u
oF4o14gyx1nhPPr3CGkfN6bWGAWVldB8JVtfwFzJwZG9QMsSAk6pUjy5K6h+OYGwoo1ml+CF2ul4
KFWJ0eQJemDrinyi/jfl5IQVd8NkReCTPHe3Y3dAGnjQ50TqnZUbPJpqhItN4kxmS/Lg9mImhQf4
MZjJc67RfjJ8m4S7eLc/4pgcovzPvfzKdHpiVFCIqQFynxBuJdRUVo739hHzA4QZIw4xpk1AAD+7
WzQLeWhrEv8S/pPTujK4xAJDZU9WENiyDAQR+IzLyOWUZjKo9THfT+HGESlHAumMVola9oucYjAY
liqVEdQRVLcBArqHFfn9jDLD7xKU1CiLyAuanCRKChF13cucphth2h9PT9sGsGeOL0/1EpvYqVxR
r7fT4YFspCo7x03MoJrEjh5M/T8xkbY2uAsKGfdKQkcnQsAUFikUrXjXH1F4hYf4G59uYrkzgBfH
/BOu6xSN6C7l4DcbgjLtlM/LzOWK0nZVZeZWAyFd/XEjkVzR7s8IksN45b116ke0y8tPMtcqYwnz
qa2EvJkS0KH/N/VaT82adahRvS8jh2ip6HuJtVXoNasnvxd2Jo+HhQKq9Xb7vuZnwrgZmklqMJBb
C6bd0WpWoKH+qpQKSVN4erDDNIMfPN1TcJiE9x2/ffQdjki3krpdrJIzw4VcOm7BOBbd8fvNaZW/
MbDJ1mGcRw9CKgl8vrt45rPrAyxFny/ZQ9WxKvLVQlDQPbwySF7U4N0tj4UxOfsNXkgJeYb6eoNj
GI+sg2h9IkYJH5DKYB6d+6qg1I0aUV4Mk0XUMBw2tF0ZQzljZYnXtfYoAx3rcY4/iivNt8TFpVdG
9wNyhHpFikdBRRtYA3Bpe/6PjzBcxgXwoXc/D7lrjPkOy89J7wnbDyfxdgfW8rZE8eyzWcmqlutG
pITeBjO+dvBIh+GLkTHR5io6IJFnlKc/kEE8xl6AG6BAJuTq0RnqhHuRU7heX1Xa8Qgfvo4BnwK+
yNMY8Bx3XnlpF0jCVRyLHMstMB0+9uRuXubV8wTVUP/+h45gOcEn9jUWqRWJTQShgEYu0CdHxJRp
x4K5mBKV/qf0NTpHTWCR4020tsC9NESBSOrbg2q7RLkzINB1BQQn8UaJyp5kS9rRXBWnx4BPA3La
3L6XcIiWENpJ9c8XodhMyuXvz8js8cVAEiFJvznKRUVxMlHx7qUXHAmBRGJA/eKFK1a5vc9PNH8X
yahVvSusyol4xlQQBjTLRh9G2NUpIPLN40oC0wR24K2Ui1lZudZqGHES+YoLQR0ULTWD8FtbiMgM
z4J7e3vbJQwoFKuSLHDaEDNLw+++lnkAtSVYs2+61CWjDjSF5boueyatHye+CD3RzmEufypc9VUn
b0cBjSkla+D/UboiVI4T0W3ZyzfXZZR4p8Z2yFVPbfXJkCKhs3NNDCsm9eNI1SXHOc/jLP1T+CUB
+FSgWQY3Sg7FWid+F1EtPLVXTUGD0Wdbg+RI34PIjSYOQFQZkiLgbf4inZT+SRvRgBe3+O7mlVr9
M37+mpEj7OlT5IN+WThwudXRdwnYOvizsH07fYLa8c/wkr/23/RzrFbZPcqR0a4uIaRLDftFnFnU
ZG5Ghgy2h/8gsR5OpGGNg7aPllFZwAs1A5ULorNlQgsecTnE+rwhSvDkpnJCdyCUeKtueYPlto13
kIOV1ou0CoLX+8rCxS6+rf0l7ENzPHb0cp8kDbNxVhEkSyxsWH10Vbx8Ay8PcqTfxSKxdybwPff0
GMm+/mj18UTN6vhizqJS9ouen5qyotOjxrBHx/THpjQRjrnoZxBaL3AV29ZMFLY4zOtml+PcwbJp
9g9sRnQQfTx8WmYDFW5cowuN5KfCJY6M2jHkV/NaxW1weTzu8heD5XHNg/MaTnrBphLt9LbqJOZ1
ajXSAFZ3Jdkl3Nl1T3xyLrD809Jhn+5ytYpHYZR1/vFocGXWZgCD1jN7hM8Zm/nR3bYdMScrXoDq
VOHz33kM4jz9zupNR3nyFrDbZ3yysBTpwhiI5ZTmd61oZ/JdNKz+OrCwXv4H+vU4eLOEustCPd5V
oqFbcSaLqYMxQFLtJRP4aSRTztEqSt97ML2pg8gwI01VlRjcDBk2IwTH4QyCUMVyZuUcovqOeDqW
jLXKV8vOlXfP1H0920htiC8DK3AR/ls07wXFzVDC0rSrKShQbxQN/EPjRereEKn/C5WeE++haT7z
3vlI8EDdwrdmbazbBnaig6NUBhSJWE2Y7mMLxm/QCSBxbYJVCJipbi6Z74NCLmkNAoQCkLc5Qzl9
S2XgpS4Hjaw0XJa3CkiBrxyklqmAEih7E51TFEFqnqDcBmDHdQvLIFQh7/Gvko7FGcZVPMqTXgmx
FfIVc1/44AX0lyN+8GXhdg14IPhWOsbBx44RT49p//jJ5v0tBRWFLpIPl8RlYaYyhTW8o1zGD/h0
+GUaY0pCHRRZMz45siSIGPagpQIKRE4ZyGBHhpZxlBWuUemue118vzpfmHnWzAN3F3Omx6+czhNm
7Of69dF7xa2aItY84vQuhj5oqf7aUbzSYXJQ7GZbNX6cZibQgOWkL3lS2MasCCgq5MSOuAPL7iRA
/b4RfCDGS/44DbA3SUSc4HExIxl8HDxj7As0PvzsXH5W3AAmXZuvtFSPHx40Yz32FoPsddphkdah
MLGPxPjPn2gKOozNVIulaqa62NMti/ajqsQbRYDmzVCZlpzQxocdfG1wu5X5c0dNG1ifSnEbdMUv
zIfzxHwHNGwNWVitj+2vVq7SgSKu1ezAQHNmUSqulWXMzA6k1WTxMfqEAmVOScWuCeSPHcUwloKL
85LWCOtRVz8vqaeDqWtQFBwMqqBUc+oSlz8HWaHi8U7gqZlSuc22T2lX1CFRqUh5+jHlDDqtlK40
5m9VIORkGTDwYNi5YQuyFh6qmsss04QA7JahRB948m/39N+VCIT+vIDD5cwJzS9lu1akqmXqn2Xz
sB9NZKS40oMEvECe9eNymt1cqa5V9rLfWcOVmxCnRq75n7Dng2NZ9IXjUAygldDRfkhJad+tDyk5
oeG62SItusDvDPCSmlR6HbjsEJnvnRs4WXY+dLPdJt0Zw8FQ0iiqmoKiiknj0TdqzLeR06gyCNAT
xhD4UzBKyoo0aTk75fbjzCnb4PCX+YD1Rhuer5dd9EQaGETO7oB+YeVtWJC6EfErVRCWpyZ/Za5q
a8esUg2k2AvJ+Xn1Aca3cwszmLiNIa93HmOkEvbZaAkoAl1i3YXM1i/Nbl/980hPJTD67a0ZDx+x
fJ29dm7gfMy5JVP8GYbdq8EGAtHnQ0+2AkLeI4pSGahImxTZ/iR1mi+H761XnkNXGcHs1Q+Il2cU
umDnV8y9f7cescR0rAi45sDlR147zsciS9yV2hJL8+bvtUgBgNJHa3hN8X/WTa6f4KKu9Jkd0MwK
tC/xj/BBl3YApx5ZrJ1oYFMz6flpQUVMovt/Dr8lqAThl38tzBFRQhAPhtZfOda5Js1VnDGC6mn9
Rb4emqpsA92RR3Otldr+ec4A2usc0sOwKvAU16rcxTJZN87kMiSGd8dqGjwozi+njFO7X09oPFHc
bhWDqwQCY++Kkxs0R+l2H1z63OJQonS6Cj4fqW7uGDYckESBoj8kMIWQkzQhzxd2TuSBkFFKWSyi
f7y33oN1zs5ab1NYSCvIyHmDntCHU3Hye4WtVjzuDSaX3485OTj7Cy2zOPVjxwv5wAn4hxdpM8op
FHZYvEYjWs+o2xcEQAJzY713ZwjK8mnzSmgjVmgu13EcOwdHTQCIKUUxWud3GlXJLhYH5BibL4rI
598mqr8UkCnlO9uppIQXMWjQS+/1FA9ofwntPdnxYRwaXOsdVk1bfbqrKz9hAjsKSZK8FxPuvgxs
kl5pDomzKHroX8fe6lvD2fqk6Pu9kfN5srPt/8BDmcGzcRV3EGteBrkBtqB+lesbZlcy+AEec/0Q
fY95C2MA3OTTQivTwyz83O6SASV/Wm/j2iW7zy4Oh8ga3iqLM8rZoULiTCGwE8b2uVh9jNqxckZs
R1FeLR2/ds1e74xT1F6202+EpNmM5MFw2jv1uBr3ART0IzITQaeJvYUrsCzHu4tMByG4m6GA8dGt
R8CrfrzVrLl7FJ3qkEEauq1VNTJXkPvE1THfk1Yxga/qEtfYBaQJ5MSwRP1wFzYATSkVApTTPtLM
5HD8ytZmW/3GkunA19pk/8rBM4cvc+EAgRm1C5ZtVY84Um7ckKzKhI7BAiPz8E1CmufHhbko9wtG
eFoxUR+9HihjUyGxDiRjIJF3qlFSdoIx5PM2lB1rf/Mtju839EbhR89Bf/2aoaRhnfr9BFBibdUK
s+jMEUA0kwd/yb0z9Rh2FCyEcy9T0F0lFvrTu3k5yV8CioqOC0REOffUw13PIqpC3cs/DT5pkX5t
8aCwj6OOpNQ6So+HLrYobEXZuSuphfzr9sihn1PPqDyJ4qSqcJFMnkdUqCpx3SBCU66aRZOuQtHg
ZB3Z47p5nQF3CMDmBqPUym9EilPabhJcggDDpCbcm5qdTDiCEGEF7WLii4fA2qd1YdpVORYC07Np
1Ze02nn3Y46iAQ6mBfTg7fpFrzuI7xBdBfOp+U3aHBkgRojs5fMIyN+mUxesWM+o2NKSJ6Uf+URS
jERBUK0n6AggmApOMmTW2xPLhsKIdElpyD89+MgksRbQFggnuEZBvCwNTZm0m39rT9p+xkDk9KSB
64rjYF9m7yYiNusc5xdgn6Pgz0YiNKMxgmr37vkDWCY9r8atC7rYVIOaK3o65IiGiJTNj6g+ThUb
T75ntqf9JECy2/Ple+aPb2YMWbyt+9iWEha0tkKn/YjgtPVMH/SaOE40kY6BCsFThzVWfGTxMxiB
JBgQBnPsYxbaKf2lPNHa0MAJCrUB4ETP53oZbSQ+GziSYUwV8M8/cDMCtcbVIbJNZWzgMAigqDHm
hxh+W9clkJdhzWZ0tW5YhUNibWoRC3OdRxBPA7r/rKpBkFGDsaonQNq8lxxjmUuCZYBfDIaBuJd1
aZXHjE5orgWbdDZONH3eAxWCUkylQcSJkZqNb7vDDo1aY8575B/HV5Y/TX9GgtbbG5QatA573k1z
pWqiDyUcxcrlAdjKrYbZiZLozd87yi/cw11Q86cJItjBH8ObbHeVSHq/TT5WtTF5sxjPvYkYNnHz
WGxTaU4LUN17Obg2lfCNICHDzVdhUUjJxXu9s2D5va290lxoNS9TNh3d3B4D6FmWWn2TAYLCAouy
81BJc8d0B7nI23rnfGaJ0Gvv46EvFBPE8CIRr8ilYISNaCAfnLZPtLtZQarnfz1iQl6f5WthaNMB
Rw/WVEQelQ6jexQidjSjyRL075X9LO5vXj3bCqWQ87U52zw93lYbLKzro7+khOAlwDtjj9Ng3Nu6
EIuFnQLHiytEVTNX1fXujsv7WlJXNi0zsVew65UT+VdfS/k0fGcM4TVXbWYPnOS1jdrluAR4f/Qy
iNRRf88BTHPdUJaVUI6x8moHCTkhI1ohkxrmAoWTO63xSVakR/zLtOmEcUliDdBXdSF4qUHobEEc
jMQa4beRBjMgxemDpa7szxmjYTc8bVWGA/jIsKb4P/UoUNeBq9lfX08Hr7QoyG0YA2+Is6ysTgIj
5fjYwglgv2aIUknuNAHhY0ultvcZfjOzTLMnRymWPH9kabAlc2neFyIsJADp8vLEOAmIaoG6OpDA
kTZmDB2rlz17QcQhxFfxUtFiEbXeaoMdlUDEpuX4QIjXCGCraN386YhHVF23ClEoCtt68HkTaa9p
Xq0LnaMsjFeyi8SiTG1nlFJxzZUvIkSuGPEnfa9hCtxKP2VaS0rSi924GPrkrr2NF5nTuIuer1B7
lJT8v7478awAlkKav8OzMmKvq0n51NnD7hEBIBXIKJflZMxz1MWB+4MZD8NSuyIwUvw73VWv81sY
vbgUHE1XkIMawhZAH2JeUlWc1V7wr32k14JFKbPS4BIdCgMs9Y/bNP3tA/5MrYLXfMVyxDGPmd0P
Mxf0D1r+Bg9TOtLl7tMHqF7kQvrVyFroouT7E3R0vpsfiTvZfJC2FrO2982qInJIsu2pd/AiaLMd
81OF2K+phFYSN0F/IhJszNV4hVDe8x9U4gCTYJbGGXldyGahOBGp/eKAJkna6YW9YXlcUfmMcTlA
u3VqbXIlcNXCrU8s3v6EASl5724cwSPTM+BrklZsFS4HaTSA0pyNPOjtCV7UGejOknSpZ+3U/Wqk
9jlcNZv4Q3/lM+f9rZwmdzQMnKxeaxMpyCTimjAo4/HtsOEvfkOs0aSIzXW+6sRyftSeW1JEepP+
dKQzeZ9jJfDFqgZp7PAV7H9oGR9LjZOi0XP41+4g+jtYD76r6jvY9nPUjOIXvbHfWiVN9oUBQsFP
czkoyUeZlJlnV4aelFm3+sp0HQ/cIrag3z/T6/190wBLYi/Ak7cs2va+QsUxA7duzxMd8NVYo8h4
liUSD1e13ARN+dQRlvZB6BUGC90laiDpz2pdK5ZFmbik+DmtptBSE20D2vk53DZeCctgtVour9oq
Tqu+qM7iVzpLgLx58sARcu4H8vlryBWaI3NbXd2CtXD3hB1iA80D7SqOT0H+nFsxZbDaz5HaW3vo
OqQQLtuea/qvis9hp/afI45ihxd3X03fu1EEiOjrQWoObLhQXlYOz7fLoGoXtTqPM8p4EUHazU1D
QqeDhiuwHuJMQkV46DMn2fEPGKO1B2ipCx0VTgsQUwi0ckDXe9OEkC1Xwx4/U3Z20mSSUPyqja0H
nztqhWCIbcYy54dM/NznBtjjCFrsHjtDCj+rRufzTIQ/HEoUGcELHhSc+hiAPeD/QctSZoW31MKJ
S5ezwDIcFV5PlCYxMo/fswZPKxmTjRStDO7yq5+62avFDPWvlmqQNHEF+3JeJ4G2e0JHPANnk3S8
Gm8ATkmWZAs0gvMdkA53TWqNb+hXq91t09DjqjJw8KqR8ZrVGMlhCEdEuRSJoBypz8uKcmFT0rhQ
F0uSBHT8BlttkUU8zXv8wNpqATSmKPiVc2XZeR8CSZiZCZvItA9E7g7/YrAMK1l2YT/faBb9xnz1
HaJ0M2XEVKhZp+61x5TeH/1MNOJt29/KQbbcLELxmSPFsUZR8pxBkevbja+4pIT8j4ecvxNLTdbm
P1LcaiSfkQqFKIVCk58jh/bm2x3ndxKAGdWCLYVStWt9z8HiHlZidXoKkLeuQNu6fTvFE02/uDL1
YzY3lKvySeeRG0lBnFbKxy+U/HyYc5EKY/AUUbSi476clB/oV3Wxw7wggVORhm811NFt6QYPdy9D
0h6+PBGvdH1NVKF1L8tiseUwPVL7XxRXB2SwIwu68YFokOZgB+7ikDxJSK9QP5XW/fuYqhCYoNhI
LRImV5bKwVn7KXFuNDfAbPfeimsatCpBmAMdYzxW+AKg+ZAAXQZf0u5HTwBzscYraV/Zgy9/Ti2Y
2Lipc4TRRZ1k0hAiRAmVTnM32YVJAAUlWvvYiJNu8Z10gPrfYewsuFtwk7ID5UtXPmEkJBLOWYbe
F8FdzHgOL79MlIsoFxKwEUST+EDmXiXwEeuog9fE3MpLMf5zLlNxiqNqaUg5Uw2XOQs+x53YC9m1
L8pB3FaLfrhCs0phko/Ju0aFXoXrl9fMtFwGFJHcE+J0wijMfI26IPWF/4e+n13sj4dpKw7izuYY
v2LXg4gXKJBqX+hi4HSbWk3oAj4IdLtdrExSD1WlE6a3fckUMS60Fv77RVNwatGNJ7ovHWt5lgb5
KKwMzubOq1ZzJZbnJkuMWPuZkZ9k09lgsaQyJ7+cDYwcOEJpAkj40e4OYDTcDf7O5GvEIxARzWRU
LP8O/aTps4VWFP2veCkpy51/J73TplNfC/hGYYWyG+aQtoSdloORPDEyzmRQlKKcWOpf1IMnS0sa
eEBSiYtevI5AdNHri9Ds+pGrBxuf5chFONNEpMaaxbdq+OWw4UCjtOFhraXG4By6j1FzzsaTl6br
EatWux6SvCDOQM/vjrVb7DMM8H5D6spWmtjzZfQ01MLy6H5sQgEbGaYMTxi6yCRPpnQocOE/bJho
d4N4NZu+jNWYga0CbTg8Zto6BlYFpOWdbK0VQQ3YLOes7+yDDjtyGOo04tmz80ukiDuW658IKkIB
9Ts2c78cDHtnwy20V5CeZrkCyG8pMirJ2x65Uv1wJsn0dFzvu34c/6cnOXuimkMvwnoJc85sxAB9
YteF1fltU6LvUTCU1xVCne/SGVe46ziipoe4CbMrOpmSAqFZi+TKDMkRlZgkBUAY2W1cA3MMSE8e
+wSkM0BuIqy+WZ4a+qbYa6Wv2dN+MtPVGc1bVRPivDOqCoNM7OsnaqWsMQbnkssqrIxSwlcn1V5p
ueJq/LqBFaX5zw08DZdMkr3oj5L1BDkWHZ+h0A8Z7XBuH4e0ewSbFyew22070G0enCJwtObwSVdP
T3duhVUhAnHlfv3qlT2f6pDa7iggzYnVSbEhdN0owqc6uWWpPFU4Xta4DjZgsZgF03anwEKpxsSP
LbVi8niPdCLK8E+z/yNYGRzNqNa6gQKxcsTgTqqYvA3sfA2Cvtfh40yhwtUFDtG5arFOG3Z26qB6
mDgBPq82jclh4E9evBZUfNHIVigglXa5iudeEPPM2ceN3SvK4x3Npl56LKp64c6sC8lCUU82NyfO
eGM/rGbxn40EcD/JgPhidHZryYLigaAhzImUSW6fFqvKib5m8ervv8gK17puxcXBSiHzfoPITrEI
6QWkVzwFcaisZCqTDBt3rKbP2Gql48aLm8KP3Yz18hkedcWU6KxLxw8mPi/YjfEBT/V7cSNYVEYc
j9jcetMXv8XvbmhnBZ2KBzGhzigtmciRHap3MZvgJtAOicLHK8iYcoHW7p0go1xsuBjzl3I0JN00
20sZTd0aRJr4s5LZ686+EMU2t/g6abEg6yy7GyRKjq+y4hgGMPnPm5WWMkNf/8lpUpylJn1u0JVy
6SphERwh3pfoPwNmyoSqqBDBZhwxH2PjPuEnbXKnibMpCM2LvFGjQ9Zzx0/5hOVG8EMYk52e30q8
4jpJu9CZVCK6LR3Fui9RFDu7JJs0yOT7+Dzn/5tSjv7PK66yz2KXBvPRavfchWoHqhACChx2RI+f
PZqeP1jz7z0gE5br+mrQLIflIWj1smZ8B0iFnM47UJarGYsGfyVWrSbgi6+kLtr713z0eaAbc4wy
iV1CjhWXWQht15qWgveiHYRedSnZ0znY/mX2wcEmo/2dLovQ0viQpffaU+1DKtOFN9EmHqZWZJRi
H+KXxNVYaxLFeXE6Dfteuf5CVXjojphvc7DhNG1wplph5Zk4cLmUUHps41VzJKagVp7AaV2+rc9Z
gGB0r8sE5A/Cm6XglkIfzFZ0OOrdABiKfnhICRCyv9ZjO/wThdxz6Gv9DJkX7OG5dS1PT/bFgfei
VMdiEgpJKtIXKncX/RCqbLXU1NwlOAHPzDOj2o1TfojVDZgQaVf84AXo65lHP9RmENq3wWpYqOBJ
wVjrkkVF/JRdAGGAQxW9Hq5hiG+YvWEGondbM+FybgKPtao62APzFtzCDA8F6ZWJh429R+ZsHBt3
P8DPKb++N9gzg205yDA9Z1KUW9dnBvWuvvkKLwDnRHe6EB4UjfB9PG9cDLWq9exkCoyEuYUjCUzI
UdR/JmVePd61F21Qhz30yB/iHtGALNVn4d81o5RXV0EkQd+rZxNhvNBtwlQlPOMu4H4p9s2FrUn1
KmUTmS5DcpaaHhFiDEoYqvugAulm144Tt4B+gdAW/qE2Cl42KR03q7yhMsHc8+4wy/9uzG5u/Qhm
PsPmmaro0/aM5STobhqC8KLpWcwNDwScG8UvwwmKtZTEMyCGbHggnf6eS8+ix/2DEoRgwEXdJmCD
KJf8HglKRyzDSdfiYe7I13IDnVYdi4QO/AMAjD+KUnZ/j7U9DfHEkp6+DFuYHaM/mHhOAl/Wy3CE
usUfPOrGeYlcjMiknxDz613htMK3Y+26LF5HWiscxGiYZ7PH2p+Qbr4I6GYb7mVtUaDKPJgoaaLo
P1s7ff5+7YLcTHHUphTK+xX2P8PL6rabEwNuqT3Y1pS4BbDOYdYth0l7nhFS65+kBRRAEa1GhDsx
TAcYnXxlwqF22YvjE9PUcJPDdKXsEdpJHA3IlR85jgClndtiXF4PhGhdGuwDCD+9YNOJJbeUE9gL
A8wm/vgEnHZ4FDbI5qv8VVMaU4umo9vN1H5FqVxX93IApuCthT4DTWSvfFyIqrtKG+Z7y9hg300M
ezu5FSsKmVkCtN9PeWwarqZ5HUz8b2nHLlC3qE4MNeXaHNfztWUO9YtAu6JXiK7g0q3GzqZg35ZG
uYW/wfcqR42AHpTpfZj4dY4fcRH0NCbTJ9iC/jw+otzxUnAxYHVPuP4HcbWafj4FZIq3d5GkK5oN
+vBg/MY/r7BVebx7gaHNnlc7Und+Au2R6B8/TJwWBJOlsjYDVEgGL8eLCL9KAmwSmsny7hUA5Buk
IJ06s6nTprOKtUC4urThdWKB3mnV3cEdrJGU8FW9oQkasfULj5F3msQHn4utx4o43t3nZmMtH9sY
btroWAkfFhPFf0KnMHDa++gQ8FTYY4FUD5Wc4myV/2xfsn/qGKJU/AWd7tydmoFYwTRkLtklk7hW
npTrFZUU+FrffEyfq1xWfeDa5jxRmiNzuDmfEH4bcEKZHwnkjYuVb7+HRwYklvmjyiJc7qeLLEzX
7QP2RoqFbKoiPbibkgE5qhjWtcPlkXv4AYCVOetbK0VROFEInwEg2iPkkLdGUXzAUz0eDAdYFN+g
Lt9Vow9BcKjH4j6YhruFvQ+GlgYl/z4Lc0L59CDR54OhvpsSQhZWUyroqOqOoczBt+EjwdfayWxa
BUbEVUBqkDJcMwPNe+cUKSu5AItVOlGnPCjw2fyN3g9RqMmYrZB3axdtf30gAftWEdr40JFEjAB9
Ibde6AZCZuTJZLuaACIv7nwHKyemRp+10Wiq3mF0LYFjA1QLZIgU2fjiLei3hutaJ50+Z1oHtTSx
+PjYS8i3oXpJHGG2M1Zc036d0Fq5nEjf7umOwwKK9Uauai9ryVkgm+hLTB08/Alnoe8Cr1gcsV6K
UoVXdzPmH3hB69Y9tOzxMozaLtAWS3rwjSldCcNkEg7KCOjhm1yDZaywQ7kY+X4bf4/pq64gCL62
zOI4x59IkmdXJpfyQ4zNrHmpyBg7WvYwXLS2uATBgj/THQnAqjDbf7xGc02VuaOgx0wewFr3chzq
OJQTC7CEWAcj0EOd8Bh6IQ3s+0QnLctYPnMJF2qVEkVFsy+L+BWKqy8TGhZliwcU1lQMm1gNC9HU
KSlM/6+6rM6bpAn4Tc9qvoLlH46BNXOwi+vPj3Ptv32jFKyRu+raTsbWm8an0SJjq/uk9k+EEKD6
vyVa1jG6AHL7Tji3UcNP6eKkikVxM0QUzRMmy3QtNCkmoKtYM6jZ6TMFlhLsADwz+BY1xP7MUetQ
lZISLOsu/NnH4Db945FsQypatM3ofdCpKXzU94MsZ5QyJnbSPJ1a4UOf835rGqMvyMglFEGSO7RN
jHjkbrS8zdXVLaN2fpiycVlslqsggjWd8WEvSKV93FmIuqJiT1qNYgpbBIjwtvPzXMHeJDHcLLaO
ozNzFvPmOIqdugzLVPrDzsY+tsdHMULdClpgmAjgooT1gVJMEYYUqKAq9dTSem5wsVsSm2is6zwz
Ze42DxqiIwQtLDLl9JvMtrVAZEdDWo9xqQSsMODSwRHrSIqhjyYMyXDsIpThktHpvM900FLZvtRq
dRWe/3HdpffGztxTddAGV7HYZmrRWOElHPxaByflz0G0e1vlVhFI4/NeFXC+ibYZa2V9629mZxLX
ohDf9wuF6IAhkVMG5aqDYk3DLw5nkAdxrpTQJJi3yF36LGo/s6dUpHjkxvdz8yOm4B8ov9L9GoVq
3r+Pal8OAL/0E/BuKz0gQJ0yJM/SldoZdYIfwz85HuQFNL2HxYjMagMA0WMPib3fLtI6OY4FLiqg
pJ5Wgug6escxIS/y0Mi7l3gXe1B5cZQRjMXtW9kqZfjaCB2ioOuo
`pragma protect end_protected
