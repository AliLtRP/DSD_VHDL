// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:38 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
kpYzrb+zr0ZnBR6AmHUusn5XkUMGCe46kRnQpM+zG9xHy1S1gVG4wRX2xIvy37tN
4V+iNosxZrB1r9QIjnaec7aXgn6dYyUH5r6LU7B5HQHutQas/DIa/iN/va93hJKT
At9uYoK9o1oRSFMH1XmrzCDHoda0psXQT5+SDFMVqkk=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 16240)
it+cJTBaoRLGaOxowpdXhHGfCVUKb0sOqdxmbvOCmmx5UfbPkT1XYj7Er3PD9GIG
s+xfjj0SaSBIb4w+GvOitvgeQ7WjQ0aDpu+c9s6+Q5iqfRr/ggw4zwJThwM7+9Le
1PdFknCzvso4e1+WfPkf+/cip01/HaofQIPHLNcVUNV1ybTHIkwqvWsobgqkEctK
c2tnADsESifuGs2eQm5BmRBQIYePfE3D32jmMo+V6qvSPDg3Ex3lKPOMWkvqV8iT
0Jjy0Dcs3MKMVSWx1Vc4CM744gurnIh2/YwkWsGlWnJMHsQo/6QMi9uUD7eYqKIb
WiFwKrCQ/Myw+vKfYQyJFrpc9mQDF/NEE8qh9x3h3rolq8sQERgNsWPLqCYkfuRp
KOWiAdkDWgx20HBiMX/dinz0YXTaSh9+Fl1B5LUPbQFw8kglY4g3ETqek8VUXr0S
86h2OUUjqf4CZI5foMP+5/ZJGSky64MMX4oKVukw7n8QAjEF90CY26JUdrIWgjxX
xwGqRuYBKThXZH3o8MtwriXhGvz56uYbuQ6in1mYKiD8c2wkM9sgYnIxN9eP55Fe
CWnyxHgBHXFZh8WyBB9cSKM/Xu4Wzy6XectSG1PqENansbM9d0L0Kh3ro/NR4H2P
9bHr/71+mVa42oxLOiIvO2eaB3OZiTgNphWnBbJz5f+fcosIvyjxtXkXXoI8x31j
13ZuidYTj0XQnrToRUsyIUissl0t/ZobZRwTUpu9E6l5Fla0bDc4e6pMz8oPSz/a
G47yTeG90CMOZvyzRNCEWiQr/u8g2G6sBHUjThXzi/7Ri5P40R+LRnOIbaawXTTb
QODQbf/MV4gBtjFqO/dRcZZHZoXi6yVYJl13mQ8gzUArD6cX9aePZEL8sanPnGQ9
F+QuPLhdTcNcx8KJUSWxjI3A1ps/GN+2IMFXt8omCtNwjtyudxtZGysu1SM6KD0m
HId/n7X3SCQY3Vq3EmYyt3lUNQwq7DuLvqQu6aZiFn07OO0J00jHNEb3b3qpB8kf
7aOD2L/DS15mF805gmld49th61NLlj6hoAz9OJ3IKAqaNQSlH2LW3ytOLV4CMAmT
5co7/Q5sZzhmTVrk1G00PCKg1/nbK4Daos4GSUb+bwurOn0z87K254ErVAYsmhko
RdUWwk/fCOS+lnudY21Q8lixZkzjEGJHzDYzTtAU1AldhB1xoORfghWpgD8+i/C+
ecuiEbQ+zUTueFiW+hL7LNypXS0dySVs6LW8uwBq5206+zzfb3AGQGNOQiSvFstw
6vtP1+PTjgv6fUVzXaVsBfvbYP88khS97KoB0eXLhRMT80MFacDKXAiIoN3LpcnX
Ax1ffHIcX8x7X1AsKvvqiauq+7Vn2freJVAlLCwAMmEmu2Nfh7i24ESz/NAJYvVx
KSZ/EtxEbWN0oxit4jhHzNeWcWL96GtehGfNTXNHpnByjsei6b41XI7GO/XqBo9J
tNFsMUxDwvyUFQxi3/vwtgUKVcDHW3JtDARUdZrdSfnOtKLS6OxQExAo0kKgSdqP
mBwYL8AuDDo8hue14kDHNjPy9hGxS384ATLkBPezC3y35x25vmTbSD39IzGtY4Vz
h9cE7m0v33x6d/a4lY66uZUF44blajIqCOP+AFyrVr3W964NxlOX2NEZs+FvM8Vn
RE4ffL/zxTBTtd76YINyJ9pzdyZReixVLqys521R8xGkEYt55my9s6+0haS6J+tB
PHYRKBVjZWsxTJ8TMY8m+1YGY6bOqUhrvYpBmr0N+t+MNShKHagG3FFDdGF+La5c
qFGgqRBMk6e9VHohUoxmjtPgcH+eQQy8xYXguZex7Up1FZpE3R74i/XVqIoYA/RJ
hlmLNYzADd5o36YP23bLXZ1FdobqToHI7oFBKcbTYXWxYClOvbEQSqhhkiX/nIHA
fIEcEE24tk4eLjldun9G5Ry36JIQHg/PafWycZxouX+Mwmz2rZqBfIgWNqNLlYRx
EZKf2Qyt+1RzQTacyHMTQcCHB8AtPjfAJfIWS7bZ8vGwHnS19hhZWKnGuSO5Expp
QL8T0V25w8KtbCoFZ+S50DWgol/K5jKNeDj2/Mwxaj+AAmp97JsaHeoqePE9FoXW
wsVwFfT5I5b0+H6zpEIbOuFeN2gBw1gxzgpMk/MmqbSGWiH53YBlUOGcQoBrIVTt
EdYdYZ7psSw0UOQCHZDvJQGzlm/oVgyCKxBlDJo9eaYFEBuiNGF566PfByJKKJjn
UKfF0ZwnsQnP04rTslW7H2T4MBFtMjgKxmFTwXvIMNHd7bBUVIG1ahDiswdARW+R
ytKhJXDB5oroPygeBbDR8wYLxb6zp/xVSJYM08M1YUkTkKWx5ejV9ouYhQRQZ0xM
IO7X6hkf5YuPAwlzQjgN5NCduSc4Gc8Jfytgzd+XptN1XCQXrf4nhz4R/sB4ts6O
mJZTvNyLi9wc6C8Sgz0NXmSOvm5FAHXGYMD3k+/i6aTdZxBnh6m4U/RxMprpzSMW
UKAhFJO4QOGx3HQRoFo0DEsDRToSqaonLv6R+jsTrA8ODB3OkTmj/d5KaU6YGvdG
Y/nHdtTikd9XYldgvyUE2rdR2JHxJ7Ia5G9qlyOa0sdxxiNZwYnn+y4824vfXjsD
A3JqqaA8JrgmUvD2uX0jfk6r2WIxjN622jNrz7GQe1xSTLMmHaLQy/gcG7NX6B+k
WIpKlrokaXap8yrIcL5a8zd2KIyr0j2Zb9iwRri1sAUvn6UMjsvyAHjLgcRB0DRT
Ptxj4Btze/m9OD4O3XsntSiDl+8zNKUWPcRmHVEVpR3vmqb4+muBxNZwSZSvLGCm
06kWY57idYUQBcWRB497FJ8YzptjHgktocYAl28I9Ar/B2nP/Rvifc6elx2m+HT7
Kzfw0FcH3fP0py+CfLGi70dJGUu86nyI2Xmg9FChKzL8+MGSHjNtkASMbzZ2lvKf
0pPLG74LOnAZSEfQTK/fU8ntcubVCqcfWaX29hePOD0hH8CpD5wACAxIVyO/ZsCM
2LPGWdeu353h4qdCAcHvFx37F0xfOjmRu1+YXhhLyz/PN2zNFZbsWL28ZAxD75sA
ElwWquxiPdrKBUfAOxoMrObXdjnnxY2k+L8zhY4YdoeL8BGf7BtwLlyi9j5rSCjX
/IZcmKN86nw3DutGfqt6XD+Sw8/lLa2jxKsvXvORINnMDmA3YLIwXffmEGg275tK
qeNmpMcsZtaF4waToZeRisjhqsoIxP64zxG40znQbeG/WxiTrEEbj2BzNwKlRvbg
lLEeVaCyPQSNL2KBW927hfVpHlb6r/aaiwQghvPA03bRt4Nx/AB75UkiFS2eAi6V
KofDwgd6doaQ5edo0zrNDGAh+9CwEeYltNMw0s7dYDeU9r3zVX6lTP2fpox72wuT
Pi5UgRJmuiFtF62487eX+jzHeZY5hYhW8SqSBiZeLrGLTf5Bivn7jn1BMY6KENIW
FmIgvTjQz/Xx4DEZvgZPx3ZHwrQcF7Qaj8fsyakx5oI0TLidKjfdrlSEwbyaQfVX
guA/bF5wKw/fg6/HjClApEpfHAiv+ryDE8MnnqCDnQmV5a4cGgWPjVjnsy28Bees
eBa8NrjMosa78WSLQjrkNVIoYnwgEdpi7qV4oW1xqlmB8m6dLlxX5s5I9gRbN/2m
OwrJ8Y+UVisnxcS0kP38FhtPhmNTelYoVdr21vH/W3MBmnD3Coq8AhuQaBvZkH0U
DLvrotS2rM87oD4aSV+650Z33Md4DazixaJUIsrcN0sUwxhRG+8e3BhlDUZIcFKE
THJYgwyb3cJdHP7OAeSBEN/YP55ZwXKBm2PB81S9WiPdNrsScqHOb3iUHeNaECPA
GPcxDShfN7+P14SSRcMJJgMpYAg1SIK1yq+wcdOAzLGsSe5/qLvQMkMjOPMBJRQf
KD1mNeukR4Sk+xzclzPTpqGMa9lxBCNiK1URrotDuHG5k5gfXT30eTIEmf8h3W6x
Ox5j2Nxc+05O4a4g/TdE+WnbK0US5bq2U11ib1fYyJCw2DUcVmyKx5lAiL2fM2ec
8f4J1UaWjf97xGxRCo2+NkRD5WbM8gaXY6cTWG/lmJYue6QLlskht2biXayR48Df
qEpFw4QKIuH9c94fX94pxKyedJf8259MrjYTBagA5L6Wubo9TP/YuJs2iZtmEXuy
dZm4Khv4OZtrwrEcySV70CBQbAuUiBzwR/0SAZmTvByMjPIu3OcwFIPo/qIQRkMx
s2dZoEz69f309p0iYDE7mDonN7HCqMh5wJUZ6K6bsNLXIyauI9KecTbrBdgEMCvE
pMcDz0Lkkn2sDFHGMrcY7TKixe3O0P4T/OQS8/vBdNUpMJYflXPVxEZDqneQ6G9+
DXZpJZPAkPfF9DasxiiGh9CwHJAe0ckbwxA96Yi3NVmmlpoXjfr1GGuOLeZTHkEl
XdvL3HZcKRjwxxecUSwARneODTjzzM4tzC777YQ5ygfrKmnlDKEuin9K/LhgIQrm
8RryPrrpu48AGAubv/WQHlJrImq5yBLxL2ApnlaIv3HKtM9s0iZdhF+juv0lzsrk
4u7MWpuZn3NDAzyj+ovfmBeZflDBJwxCYRriKPCTtv1urZolqluDrKWOf738b68E
Vaa1s4AtyJlnI8ZTmO6cW3xGto2fHENj2cu3Ueabv/eE0EEDXPLqtIU5AJtjiBaD
2YNls3nEV4Pr+jhnUr0bbr5lJSquIyEO+/gi1JX2t9I/gPthGDqvKrWgwN3Vq2h8
6Yc3wVESfz0V3TKou7QCxudAmzGje+Nep6Wh/nmqnOky++ADEtppilwPw8cTSD6u
XMT7gebSIyfG/5zTVw/EVSjkNy8Cgm4CiNxQXn7/SwgBqa8jsnn2PMMrEjEUTMuY
XwEESlGJmBd1zTevQsOpP/hYgcKxE9x4eLEE2EjEx0BvnZYepXvEPCjoyTdB+3Bx
QBYv/jWAxtXElDa8DvaXqKowqguPaHYAKMqMEbEdoaL/BGre3XC2lszinz4IHPNU
9Z2Ak78TuocHx6DE7hkLLvQpm93mtykwzCAb6r6iX26jiVBmO2/EE8rVF0aPj2iR
ZcM6MZh/lMUIbBVqHqDfbja9DvKj8wb9YI7ujQdVw5cqwH/aSWQfkIW7DDAHs6ki
vIKMbP1503hH/Nq85CUs4/0SB2xpS0CQN2FvwgXtwE6XfIhB1ADA4uPFx+/Ufzgr
63WFLOWOuI6S/v1SVpeatcv1i8zxIb54m9c1gDVcVrlTH1o0zFb574PlQIyM0bcm
mDPnK4GBdsdevQr656NQhTKuF5czSit6rSBaUOjOOqMHCGeSLQ3pd5AtQI78lBp8
CBYDy0vGaicmmnvybst8nVMbCBUjn0sKDoQrJgZyKGnqk21D2F9faRdFRMiiUiWz
o0By1lXr5tVcWhap5KrQLvBAxKKkgsI0zYaOT0mXT1Ps34i78CXNCwRd94luY3E1
VrAyItkHS+txzsDqTfsefIyJed2CUBQFRjZjrpL7qORdYlkW7DiFsV8O/7RzHr8S
k9Z9WyreWzJvltbsLG+bBYMzxR6yYYKqTPyOXNeo6HxYzFEfoMGp92vt+oNRbC5x
qdl20eD8EoOuOwa3/jR/ZwcXjk8sSyMHZOALSaK+ysmTv7KfLVajFZiX5iNbh1dh
zBZunq7MI88DcJfsVBN3dgvuf+OBPhZtB10jkEA6fb6zHlPTRIR0gbzWrBurzmBX
vlwicp2tgxI2VYLolO8weFzQdHQnSxTaPSQD/26sVd/H7GwdEfz0nieQ2aoMaCj1
24lUuXitD8PupuS+VCzCRfSHOygbrzPrLyn/Iorpy5jsXtTZjYPzip02gykpwu7l
Mm9xwFfYunfJkydKQT8SI1Jimdu/Bnec3LpGczO2XKREtb+GWj3ZDU3NSKZAHS/x
klm/L95Z1pXVHj17EVxv+MtSulTe6M83aF2B0ZLi9c+KnyGf2ys/2DPXY5pbeldC
QPRjNaPh0V35G6EyGGYj4H9I7AE9nhrxMPVmomWzV6KWw3FJ5RxEcaSwwZQbopWY
bWi+PKdzErMkaMekdwauiRhncngx42HIORH2BghLPzw9XhYYYmGjPo8UsRE0te8+
iriowGwXek8ysOlTZp4GtqMn535uthP8jSaEUj2RhiwTVW+gsmo1OgPoy97UEm9c
yAC1d1cpc28vSoRZI6XI6YARLKo3T3Ktg6jBmnw+44pQIXI3GFhfKKPGCBeKpX7S
prLntQHPtisd3+JgoGb9fXI9P6/BompWA/peE7qVy84y65v2qpShAMtJHnzYu/Ca
MhIL4hHbQQgfYWQwyfYEbce1JbjO0ddbi1Eaii6d63gpY440/yxhblmFQn+mOexB
bI+SxWNEpvmJLfxj+YPmJHg9/mZi8BDzqup+9iQvcDFs8uGIsjJswNxy8A0m59lD
8CgY8zlmLYKsREwK95HwdS4cCQqRYyfXO7Ku9jUavxYYpCTMTFh3mI2OrRNS0Iwu
eWxWCcA4ApwCYvuV4xGyYIfB0E9asaAv3rLP6XZ4GYdYH2ItRX9XCGvSyTAr4UYA
1qywsaYZ1rHwh3SRznEaxtlwLf3LJPcSKbysWPnxlmblBtz7i8a0re6ct+PJ8f4S
Ksg/FICzvjLebxMZsVdbwa6oHzY6l9iZwN+ogKE3Vhlzv2rCSIpwN9Or2xtnQDWM
mZ9+oaFxbHR4gh/DiWX5mLX+QnJcCk2IoivFoKD7DujmU/PWPqkWxlxkPaJdGLO6
wE5pTLJ1L+7CgGJ/vO2WStKqzcUd8CXwsWro5W52ynX5wYFYRBIapujpRPs0a3g9
ioZ4RZmP0cWNmiLFgbLuFRMRwHoXjFX4vYleaH1tGIKjMdNH6hR3GyuiDy1Pq08P
fF8imaaCKSXlnhv3KoJmtieIJAhLwbf4/WJoUuMn2tVSnENSoXTqy3EsbYYTVZOB
2IN6sx++JhMH+he27/ZlNCeZO1ByAu7elycRBS6lM5ORYTXSjEWjX6LDnIbnRJLj
lcPZU5pQvxH9gfwwLIoUpMTcodO/Dy+G32LI3zSxzZjxILczW17fCFVHUkh3hjXW
oM5Qwxb2j4wJ4B3hlhHGBRXYlTlM77V//0cZxXGgzPiIIrUQQ3xbwMSK1ii/tAc9
HnAkPOTxHkz2GEkaMYssp5sf6sq3KXdSxBSe1XZtrB4ir4ox4tgM6Ts9Wcke+aby
xZQh0PGErpwLI4bdRqrp0cjegUpAs/p6KhFFqkcQeTci35sjC08Ze2cECP39NPCw
24pJyRw6x94obNnsH7kjRMO8Kv3hKuX1u1LmeC2hh8j9biCMSNF0gCxt1oAbjL0Y
U1r9F39QFA43hO1kG6ByW9Rh+iHbRh1Lgh/vbJG7rv4okH6AsrfV3vqLL9t1hJf8
APuQAHqenJOib9IevEjHs6/LriZVKObOihKyj1EY7SgjekQ2ZEsbkFEwMcwLf31O
xjI8AgeD2HtuDsZeq58mJpUTR0Hs/cd86ZXMRWjaJo1uOyO46WN8RMV2a7sH6bTf
Gj9OooadIh+8DIuaa0M+grVA+erTaJNJVUFUUUkN70nN6synsexrlMYDbREklF9/
8bo9vnNVi5/KTiLoHZenrLaj63kVDuqUy4Z3XfeAideO4DQ38CMCNBbiIjKzVZ65
2GbXuN2n4Ls/uUrYtpcWQA6edKVRSD0N4BmQ4ipSHhusQ1eubd+gjC9qar1A13CX
nqj79Z8n0gfsw7om/5w1kTWKuhztEzI8vuiD1S2k7BQbFMGLZsImTeHangXvw2QM
NYf8hH9LmUpGuXkRWqyHpyOa9/N6D1+gwV19YQ170+JZ04dYhD3CzTxlRC3zk3JC
qRdM+hsAGUMi/Ushl2Ltvy397eqVpOq/Y4DNdjppZff6UULsIXOzfRgbCK+owaqQ
0tjBGCAISziz9UGHeGBPJ5U5dTVizQ3wEkX3xmkX8UbAHXRRuHPvWSnOS4vG7vnu
5UfzbnC3btF3DhApxg5cMMGgp82cmXvgqrBEx93HTyTv9ixPEoaPwmNEDumsm6+Q
0sqeDUn8R73fjnSmiGwVebPxdWZTZRLPMcvtiLgpkWW9aB+SRrqn3NsAcvdpUTw9
+FLzFPr7FtTnFnpHJ9Y0TqyyNgXHeMTZr9wv5Pghj9LENiR5RgTGp3sjwMhKuwoT
jXcmgp6tkXcDr1Qvu3B5AID2AL8UJ5pFCjxl6fxp51TQvi81uYlDXCzynrUHTJtf
zNNdAVblTwZAnBHXBWWfDOaChi8imsuS0Ozvov8PM/17VjQXCUQ7eAOcEl17AYuq
tCUJSCvu15htgnjzNnjVVjAgTK2hugjvQCn073VmR1eH6MjdB313nQpL+CHwC2J0
KqI/6dxGdYxp/G7JNeyrQw55C+lDwVoosSCkxT2N/5m4abKES33CTROoI7x6KtjW
c9RAktHWYBN4x2K8lo71DyHvzOfCIJZ484ZLvjcMkdfpGUf3/KtE1iEmn1BVTF1z
pij+My+ieF4Ny1a+1u07cK5Uh30sIkMx1Aatip8iZ+qWIZO/+r1QHRjowz6zOFzK
zjW4VXzh/oqIuHVi78weIezdGh09hDKf/zvCMnVs8APsK6HqMbmppEcKXq00kdua
osk7T1hZm/qxcoaNIy6AL2acMBci3Fjrb2LAnH/3PtspgAlLsbLRCks8qVePsCB8
2VCBKiEwdTlT1c5dvTVIR2jrkacUxgcDC0Nz2fUSPW6CTt3y0j9qs7KS7HuPwocw
ziQFNBEmQX+wNMkxXbUgQ8RpUNeUBrZkqwyVQBLV2QCrw4YqWQ+Xgw0fPtM5G9oZ
Gp/CBW8FzcprJLRaY57ekW9CzqW4qkBfhDyUE7aZyt9tF+XQV2ZAkPcWd8IRrskV
vN4VAZGZtSujLzUI4RxDgcFCICKDYe3QSvO0FBUtzA+WA/hRzw4NExNm7rLHPOXk
G/NKqRQt2DysVSQEING4viXDB/qAtcj5aHwDUmyvGbwHvaU5dN9yunNsjeQF7Th2
CboN/biMD+HCOqyWmT8FoIU2thq7vEL2XimNoIYQ6wf1K0GnHIEkfMIfRwHmm6Gl
mA2hePbEwQ0KQvMqlcI9mFexgeosETMAucZWcye13/tAQ6ha0k5hgw+kKktMub5Y
qa+hptRZAQSBCIQEkQGOUIkglHU0SOU2fpupq6+++8cf7QVxim94zu9C38JTAxeZ
mW4gj1wSd/L/8TGhTimu0YvdW1jSlUpNhXeV+Qvb8g6NNqjr3qb/en9R+FQ+TKpe
TtBu4Wgea74IUJNoLwW4QtTkKJVnGhhv93yZzUSVBQwjF1dfV9Z/S+g7GTwtLs6v
QpgzCMxa8U31sA8lDS6aTCYeSUOG2IxAi3qIO44qy6D/b2SAUU+XFxo2xt6dmbLA
u/VxAc4Sff5FXPKJTQEmMbOjEYGC2j0EpCfB6+1lIZccxPNapl98D1QdwquPpz3R
UGfKrUh3xs4ql82PeA/NHrKc0+pBu93iDof2q5a3GV10/4mH+9VijqAZsoJsO2Wp
JBI+HJr0T0sz2xiIhnDwADeO4T8kk9PJxI3PD6kQkboBElG8AWO3pd9eobEK89sh
QI16rb2SWSmmxHVY2V/NgDoFOULWEYvYTfevX5iz/isqaTUFvidqgoDLbXPXQfBX
W2/u3E7F3UfQmyOLxJk+WAx8i4RlLcUHiCHCqBV33YX3B/bIKe5cxR/t65SFB79J
U8LvwP087ndjmSecjqkUTdgvXTZoUaJJFT7D81WRYHLVdQ551y4mDFf6NywOqOAf
CUP/kzOFatcPzzwXSVUwv9uplfam7xo7hhQmJYkvmfjaiwsRGnRNyfzhMKXEpwLP
nVylDVrtPaFkBlX+ex/1hwHkoLYo0Q2H3K3vdm3euixUirfcAz2Mo05aG9GIfOk8
0sZGLz+62OcQ4ZMdsU4couk6hAFs2zhlmEtJw8xypIoq7k5EAjfy4Oc5puTn4RyR
2n8b4gvtrbhLc0dHo/S+EZlwfmiAwuPaIMfXTJJOkU4ucw8EszXXXuWKmN7OM0UP
X7EZKL6gxxqvHsPpeQopHJbHFMfql52LK6n+tVkrT/cEHBQCyTMXCTkI0Sh/Mzv4
ydPd1MtbIADY7rMlu72UxZMjCQTsSpau7ywuNUM2CLTNRyRjv2oNOXWcTkeo7P3t
mgyNgh6pT2R0mZUAeuvkHQRy0GXax3bB4mfgGzb1Me30x7K5Ofq+V7/qUJeYbedH
35q+TTsx/nDmckhVhNHpCeSrm30rgWoYxD75ytpaV9nqIHUQshlcA+UwNz0B65JB
r7MI+JYR9jH/wx5PsYa6z6KukZkP3LttpFXCyadQwmy0qBYISYBfzlSYftawr+vO
khVqLA0UiLzrFSF/trWot/anlk4aQNgFl6powGuopvyO9qr8ZOeev9KGRxlMdZaU
h4+g01cUYd6EH0GxFXpmX0ziApzpaEXdYu0eyJTYavG2QEATU7Lsg8kv8jLDUlU7
LIQabL6yia6Mioh64TZgcTPw0mLNvpTkca59FIAG49+kTqF12V4y6GzAHUgxQDi9
VL838aI+o6ksLHyi9tdKZH0q/00wUzqMdGZbVemgpXiaQiRVsS3kPEkY//VHF95z
6O1alt4Y9467nzYMsjqmsV70ClO34iE7cLqokX/b7WMtuhAJVSnkNHUqdIFsvkyk
82Mb25tbLL3WkImTg+m3SVec6aVQY8+wlTDMjXo1cKAynOK9XjDRz3QdvG6+FgE+
mu6mEzLi5Uc1dj3AXCyPrznIepm+JE/5V5xSgSp8hPFgI46yUvmSpoDmiwcM+wZa
xeS+5cwiGb3IogkSfkQKIKI5BgYEqjJVQoj5A1/MlmIhSgf592RUTjJVb8fVKfww
jOFb9lvw5PxbagSb3CVNx1mwmN04ht7PH5BloosAbU9KjcMZ2TkQTHvTqsURjm/H
5LbbvRwH5WZ2OWtX5VyupnNqt5/5MvtXFiV/gm8+/5l5ToB6i/QnmuQOHc4F8fXC
DJVW7GnvCERXMjYPCkIcYiGNPoLCVmZuoq5leBLGhB6dmNdQfbYWfOHLRG1rQnCr
xRFlVcVjkjOksT63Ioc3TsQzgWvF6dAmDYdmrZ2qXy8fO9a5jcD++SmBL4k4oJgB
3TU6jXUegHsv0rmnZt6u3E9+I5PRz3JQaGOzD0YfhUypwbdC8fCsQHorkCnk3RJG
Tr4BNsqFC9YHuOdhiJ9ziRsNOdOuDmO605yZjtcYew5flzxOg3HqlhBW0WEOJUdH
CFHN9ALAU9Q5mouYInnVtaExLStq46mSwuWaaVoC6Hk504Y3lrO+2BXsir5aILhc
MSBoMGBI6la4pXoOQNR0pp5uWWuJgGUvxC8tjdFdP5+rHUOUq8Rw1sotvlmE9QyJ
hrZNi8XuIY7z9mZ2tiDdLDqJ4W2jmQvgLLSyyXhNqTA1DUT5bfEPPKAcW/8zJ8B9
3+ZGNbnpBpFov20HkAKrwmw/nAOJSd3e9xaX1wPH7jnDuGN4KRrzoZGdYaWASCr1
NCFxyGbQNKxDCd7GyIuOpU1HxuFE9VTH8woclxXFTXUJD/B5LX0jTrQCSJearkj3
oG0rsswDnhyrzhD2ihOR5khneKgU8wzaNsLIb1tFNcMioRaZCx0QLDXe7wj8WmqM
dgrTJJNsWIoT39yQIThBqxqwx0P2fgjo3D7ZBOGYTMhIRr903S0nqjhFXPZETQBV
mnUgD9rHNG2Tur6fo7k3MLLVT2KG95H9WKT/RlmNvziqdoOYlxhR/VmQW5EgShmb
D+l3yKF7pChmT+vpdsronaELkzUsFRsaRRwFOGtDbmsFLCa2C6z/T6gwf9I8nxR+
0BA+J2jY0ud56w64PxCVqNSqbdjldByUWLWAApgMt5N/xmoN15+YGA0WFmeeGHkO
5/rnCjVWt4bZ+dxw7RHqsoOBHfhAdX1XIn74pRPFT+v+Fs9o863EfcGdj+FTl0xs
CADYTwfspVNep7LIgRyQAb2dtNAaowV7H7zYeFU/Ds0C3RWt837rL9lFBvhq1LaN
E5Vzdzzpmt54WjLweJZ0elf75Vq0gH4CpaO0pjjRjquhXeXxaYeHmkBuXYPPYx+j
KfdFZocS9khRqepq1wK3HQun/gZ2Ua/FX1c3OYbeUxnZ66tai/2tKMdO0/kDVaGu
z8GyDYO6wmTGKiBmBRe9SCICAFIu6fyC8bcln49CfQ5pV3BdCxoR5fMwWkJN4IWp
AO2VpTWX//Yw+5/nOQWhukXLPlePqIQTNN+ZGZU+YkyKZ7C73fjk1+jmYgkUVng3
LLuiOVW9BjZ76QyWXhn7v5uvUZrqVg7RF+xOQGe1LhwkV5OqR8INuxYPDWKXTAsx
i/lqbuWYs5IrlxzA9NaN94RyXYEwXgmTfTcum0NrVxH+k349CqVbUJBoUXySOGDL
zCvG8FJlhenRG4hBBYpw7bKrJUBksvF1kYrV3Ru0NP8tcikJgwQtmm+b9y6NqGXO
msQC8QlaT8zg4dqVl0r/U3b+ErIFBSSCnfl/0Hxc0Ne7XL2kGODH6XqVFbq2k6XK
pPMrdEbw+JVfNuGvlwngNI73ta0ArdijRrpLsMFbH2kk0oIPVh433/ylWddjJQ6r
vJ5qYj5lhlI2cPcH4UWMZvYie2I+iUh7vZpTKx4VkQ4im4p25qq3vt3OM470DjIt
xWyyVF5M/smLVaJ8wGUJTdlNwQmxU56F5yIe0+hbhciXmfDbpEj/C8BeyKm8iIFb
X/UvV2WFLOINHbKjrQd5EU1pfI7PbC6UUyOqrouZmwdh/WmOz7lOw2EqWsjx48sS
dHBaY0kqQvcHtyP5D/hBU8lYT6rvqTLYfAYaVmOICOqNcgbaHNtTGYgCDg1881Wi
jGWo/VhyuVyYFQOYuvnKu8NUAMZUYF2HHaS9yI8lsEPfHZ1EQjuYjpaFScbbEGBI
q3dGgRFeE/XZgyFG2ih/NCRt6WnCopu9OKdmrLk7k0tJ6rccaGDROxywOWzoH2Se
3HdhC1L302IOs2CJVAtzjX7Iovs5T1V+bHBCkxaVQHbqh+RnjaMvBtYamuRbSosA
j3B3IK5CqOz9qu5m8WGklgB3arfVMd5NzToOfl+uTOuyGB+5uDL7zzmSXuZsWgKD
LXqcJhy9Ge5VNTT5nMlqpTzhikrVqSumMe+L0p42Xi4iTSUj5GZlAk2tVPTcDJRt
9HiCA3w3cgkyskPRSyD6VbSJ1Ox9DutKlerkCQyVTNS1UbelR5HG3Tzddj/Y0bXV
AJ4bp8wAaZurpngbxwzVQUHDe0bvLcYT9guPm/vkQ0i+BZBlpKkz1Nhvu88mrmdo
lQX3Orem8RPSOASrscZs1eb2ZeLzSy2KZgXRTwO9v68/aBIShiYyEaLxKp9N4e6g
2Jg4deO0DCqCTrkljR05Hq/lbAuJXd1j54reQuFZ65bZAsl4xUTYoYzqcrKgyU0M
OlOpRSYLG746kD8P4WZ4gBumHpLClAh1fp8mrT6rcfj0xdY20L0LALiSgO32xVTa
RZHGCPg25Rb+5+AG/ZD2OXNVuLyG7zqHo0QPYQMe/qzm/ogl2YMize8vXdags0wC
7i5uVx3pcO4fEARL3RalnAP+eDcCnBSlyC1BTBv+3KnLSy9fCXBNBeUW4CJFN2Q1
i7apYvhYEPf7/yjOz87pV0gIAhrXNCkqOfhRwtd4e8IyNKAE3IHot8ri0lELBJjl
T158Ve7uV4o3RGWUzyU26Tolki1vLqR/YPpGqMNayugpCsX1dHvUm03iIiOchNTz
yJjRfO0Vi6VWcfIDSosVqSH4Fi7zMiumunoXpe0HNTh2xqw1vBUVRiALDs3gtaeE
j6qLmOFbeuw1Ag6xLW/yz8XTUaEmYoo8RWX3qOYZVknF57Jw4j872JTGeb+GGod+
aanrVZKpA+4snLyUWkmOltTUUcRcW5xvnQAGMTao9j5RzINaQvguJPJoTmDDO+Gf
dx2PD/7zdoC5R5g15dpDKRXLJtXbCd3hnKnfJZSBnS6ROerWaDqxDdwUnZOBuY8D
0tEiapuz7pOJ98/7mLyxB8AT+eJLPvmrj3BgTL3xtkC4/TMPICyzltDIwUUUBoP7
P8jcGqAkAosWzv5j4tRzq0Lg3fxCTzh+UHONUdRA0diFWMLYLaG0tMZDlAt3zZtf
QPnAXFGnxjylnC1OhK845ugBTSaQpXscDicEGsHqC/XOMwjnLJMdzNs6CPmv7q86
jsfy3ZitvUPvXK2xC8Hym0Hm31G2cva2MxwM6ehdx4YOmBnaoOM8MdoEahFIMAso
MrriovojIW20wyQAhN87N/qnAw9QA8ppX6GlFNAhGdh0xUQFLoa33dShDC1CNn0J
l20v0VpamBtbsMk039Bj3btOcVQ8KzXELdv4LC3uof97RnQSplFW985xd3SjpTOP
fBGba3o0wruW8QHsP31gcRUtMMRHr0/LdJGmRmLxUCT3YZCp/sPrJazk/zXBA/LP
2Q+jTjbKsmxt6gYU4A1jlqgzQQOPWjb3rfJHq+IyXDSEZAFMdvYCfymNA9gI/2oK
Zsqg8W5aM0wWKBwAWy6goGqgn4dF/LWLqDFKKfEN94a5bKq6ZaZTsIFpI76waHFM
pvv2jbxRpnCcqvrjQE+I6SqKnPDfDOteBqQObV6sBCRMSntYVM22fGNYc528DTHM
qmf+/nJyoOLKhuPUKHOn/KVbx1EcpQi76AjEwp5hjIzyT4ZFYQIWbIsjJiz7jH5g
/TnMKS7PZJvbcgnrgFxIo2IE+l5hExIuK6P8begWIxDceyC2S+OKavvldJNbaXS3
L02cMbbFYFRhVPfpJzHhA9VPNkUASlr6Wc4TMqFQGJ121xtHitnGHW5ncxhcmXdA
nfNAANTeo/t0uPLR1qFlyw7NEmq2WYceZh3n04CtUHe+NQGoT4xmmB7stgMqNxNc
ORTe5qgNQXl0k4dhxTXlPfXBFlOgkBty9gayrzOwC7h+/sBOKX0uYA9z9JGr6olT
W70uWaPA3CFY7JMzicbnaL3kWTlI5OMzntwg9+V5YCLK1cJeV/lEvkhWjse6eVq7
0d/yI5k2spovhLv169sWKCks06j2yii0Ofl07H3s29oMyw2sAsyONMdtW0qNMlB1
QtYo4eH0B1mVHWHWmbmPxVAHwa303otudICF1fhGaC93f8uJ66KtK1Tn+DFN5XNi
kSto/dpQxCfp1vLfwfgIxFpZHzJOddWbmHvbFykgTveqGsY2z7Sh9m5U1wT/rQuI
qsEAxXkoSx62xleFg4nD8B6VHGaEh2fe5G7uP27iX5ZtlIZVJunmcnkW4f8KzFo1
O0P7sP43ZZjxwXJ9oaKTHOCB40AGSPkA4+x9EGTD+tH1of+tBso3IkToKF/F7h5F
j6pOG1umn65y4jAb4KHOYI7/gyO00SQmojJbW//aGow9VOjGJO+YoLwe0yphpmYy
+JOCgs8/rvwTJwKXu6DMMYTjUIzdxCtLZ6rPINIj43AIeffDpWeQLqNbCLQplaS7
NqJWehbbZxuMTmcYcpFKp72ahug+Yf6GkTIJAulvxQlWJ6F/kAIHF81o/n6avIjO
boqDjo0fDcznRnv8jaDdJaKeFHnRZkI6fZwOtXnpFTAE+oI2qSg4NFbO+bEQoZBF
dIE8cPGEdqeg/WkJQ67tHeFvLCgU9ZwqiDkDEk+ocs/1HXnOTUymnPUgtGihsYie
99JBZnH+Caw+gUm4xIjTRWN2T+TAdDVYvGniFr6gFZprC4hOFgozmEiEYlrjpkY6
l1EstqpiUaBY9avzKk2BlPTbMb2L0kehKOes1gC1+fTtrWPRsFBwErhbul17ubgK
knOQy65YrIMAeHfrFxdGYZo2dcGHzielPdmssp2FEQbW+Pyl/mllJ5P3iX4YxkEa
oxzcVavjxW7Aj/fq3G37kbvbLvkpn8DvI7AhAghRU7fBhgROz8JW6xJXPGjwOLhu
V0bSSnkFEi9vQH2qa+F88XDFd3C1ImSGRGUuzHMVSOj2mlZfaHYdWk8xZCEfXQKP
YYehG7s1QykD+d81fRB9/r0cAy8w1eilT2pPqDoOdz/xWTBTm58CNA3klplMSajt
au2/zBjYhndNO9KVabcQL2/GyM4jjWh+acigK2SnTpfCl6nhln3GXw59JKNEi4ra
OSk6Xn/pDlwZaW6AYvclKyP4qKHI4QjqlWiwZu6UfawtYPRc7YRZzG67TsF7TuG+
M+fFPVUMcxrDY9WWGd3jupYx07+2GWe9vjJGq66UQ8Pb4+LirDvNFsMM2goNHhz2
NDSaZKiIzGDydbIu3h6O/q8oYSOiQYe+b3wWtPDIC7f3KGc2ZV57t4RFkDWwoH2R
fZdFn5xC+5/V9z1AypKuzWJX1QdinRuiR1O+YRg6GQYetQwyWa/uMt1Cy8h4QjUI
12K/V6ET1yluFFwbHJ9gEbaNzaZQigywA1WZhq2weYDl1bwDZXWZy5WohXibBDnE
hEbU2VD87gywEnKSbbwa16Fpew25tS18Ga7okmGQDuOs7dWJuOprSVNnJ4n7ygxv
Zyp2Bb1nKDKssRrYoy8IbbCksC+sJeAHqqdP8tQU4QG1Vz8QvxMbsebLLFxKmzje
p5TExwN6KHSXrP8p69mfVrJSkX1oEXobMnoOUYTA9Fk86+auTYdHXxJ7WSloyF3r
p+e/CTlQuwZ/OUCwkdSlxf7kbLVfZvK/s+v8GEAIfH4rm2uJWbmP/MS692VuYEUo
dxS2EBaqy/xOVfWLuustk/x7l2uY0IHC5BvanhrgTnqU369zSyMD5ybTUt/cgIeB
ampExdFysvoZy3+MSm+7ctCu8MCuAV22FTTRS0Xr8uSt05kTVR9tnX+mVIcWMvgu
F+25KQw56IB9YkV4fX907QLFsLNF6XZU8KYMEDsqKdjmthnB6ZGmdhWG1ynobG9r
gJJcT0gWQ3+c296yRh3RSBDYFk484jxzQdMAvpjzBzVLkBsNCBsfxFWXMszY7+sV
Hse+d3p/NyK//6QSYm0JO0YDvmeGhiqehI+FHCIgbmFo/iuaYoYZfPjKlSwlG721
OFnUyuvIcvhbsbjKyzgDdAk110FkbbB29I6MXZCPBSwlc1z8QRjQzRoXyjoI5e0v
LAF+McxfEmVDlUododS8/AN8PpKQWkmXXT9V2trO2po600zxZoksKBD8FwjqfVfk
ojbUF0hfHwlVkAfdhd8Z4Wvekz9UBrSGcpjL4LMWKkzEXv7+8ovBn/XO5eZzHnnG
08htCuM/B5UAB2Gp1DL8UYJ6g9FVirzogpYoDYk7f00pASmhDU6yq+T3//uIO9Nz
gY53PmOyj+kLvESSJlUfawaKDjZxpnN8agJqx2fA45hyPN39p+9zd9xfhTQDSkHq
bRI5u+08HfJuYjbHWVh5nuJX3V8HFYnlisZXXswHRl4MoJxLSG1smqVPNrnDDpj7
2L/bwJJeYHa8WcWNp9vR5MJu/GdQ9DfA8wetYgSIGrugeuhUDKVbOs0cucsljnlK
K0yW7U0GhNNnnrqlq+0AnLgaokC4yU7r+UxDGYKO3TOXIct+Rnd7rK2d4ruad0oQ
a5s9SX0M3LDjT6BlRQqIaL+Pm5gqd16SnHbsn3/AHbe5FG8I3nNLmyULxVURtvgU
ooo6yfXzfE5x5juj74eGfPlzWkd+so2aZeWE5++n55irHW/cAHR4nng6rFA9zRIq
Un8VpGgdntBx4AGnq4On4ro1P4o1zhtAIPYfRVjy5+ezoA14VBiPLkiUiLm4zNew
ZI8MzqjkSYpf0ysZgX2GnprrAqj02kJd9GT4sRKHG7yRFmUmal6T8w9lqLNDPPSo
1McPqAfDUsPG1HOcb90X6hMpIHKC7vx8RS98gnz1nxwh/7BMp4p1VSK4iyUY/MmD
gPhvwLM+BpMCLfgSPhIYrYXvOyZGDCtj4OmWiipqipAZ+1QIJX3T2xjWTmcf9nTd
ILaBOt3nW/85F3TiVMda6rvRtKM6RwT9j3xh2Lir3b7UyCclpKoYzzJNX+MWMLZ0
sEzGk+Q5HlqGo2ZELBCj/aSWNHoi+3ZugqEIJXpIPSPvXRnYe11cHmtJsxNQRzuL
bp6WQXZKhWIRy1wR7DwNWdUubhHn7OlGol5z/f9x9vZXJY8lTSKCXK86nLA0D3km
JZM0QCruof/iK6m6rsEg86K4dsZpXtDA/j6KzsmwWo5qdisRATe/czYjXl9PzH5p
SW2nzuK4HqHWHhx2EqOpHPxsXA3YSLONUqK5nHK3yEBbbN85Bvwo1oDjd01NR1Oi
ab72fbnfRVQwB7hUUaWGbS4PfGV96o1MOblsZr2NDka3Pa9YHtjnu4Lc6MqxEcgG
aNLys0Wc9JzQnXmshSyNLFXAaWGs5sv6gRcwlsP9jgJ8PJIQwcsMpc+zvOaZ/bAz
bY/dgLEcRaYHSu/JoShBon7mSgxWxtS9sw0DsQPjVYWVfS6Uy2tkpJbFReExIeii
lPrIOFIeko4G7tOPOqGbEN76YKtuioBC0tJbXPlH45U1o+QLZH9ywbDfEAzBsu9+
3YsFoWB1vjcFeaDJZmIikRZonkxQv9uiqg0YeMCTxas4d7QRNVjt4VC+8kqTsrJG
y1cqVABOg3f2ZELPyS/vw58pETeY0TGsUa5wmeRoTg/NxX+dL5W+V9itfmrw/8aW
auyaQHk8ETEtIu6G9acr3T2iWNKIvnrh8+6uU5Nz0ZMfBEU2tqcZsh1cS3rfMkIN
7xgf/Ymj2bNTiQBMVWxr4otQF8t3KiwEJ7x+hGmloRsHtPv0XPNn09UsvPt5Q/bz
l+Rmw4TOgkyhxMyFxDMiGC701uGT3Yxhb2uKjUmhJEDhzgdf7fthqn1L1tb4SW/b
q0BXIsIc4fY9jjVmdX3apNFvx+sztGydZg9e0QpPB+EkGYxGY8XIMOsdHhyUuOVU
5DPh9NDjIvsFIFx/xEgZPl4MBJt66aSgaG09m3BPvL1rXFRNEGSh738PlACTU/oz
fzA+MxkskPFNhb3xIePg6Obsxj+NcyyT6eDsfhKYH9C7bltrnCc0gzDwGcVFkd/0
Vf3vgClgzWIk2CNvZ95txLQ07a2GaCpwSh8TwD079wrY/UNfnwcd/beNfqQvEzSf
bjrCqD/8XIs7wcOSw0ZJ2jOTLwgbX+HJKP9tn0n6RfzAfcAHRYB4lXYj4o5hoii8
94NNZxlnuVwOkM0aSCxp+uEMey+Js2wMp1zJAgtUFzNlI0EzsZO5rNFr7B9OFF68
+BNij26TbFL3NM+EiXkmSpbJXBwSysnnXMRI9U2WCyllkjMDTO7pLoJD3lqbT0bg
JidFbdcKDmm3mo65/8hvMKQO1F6jSrPumwCRMXGt6tOlOlgpdnpAKrplEqG2amxb
66tLq94Rx3uqX1JUYDjy963P7qpQED/OD/yqzfBhElwGUBr2Au8BzCLocuUahly4
Woc4qwky/MQ0DAhqABl6jzH9sEddhlNigOrCDkbpBWSXgSzbAzY8r45B/XWdjzVD
iKq3VXvwKWiI2R+0qni7+8ZU7KOMHXLtlfXHYTkY+36IbcKZWorD57k7TKos5cPf
BRvBtMXw+AIT+Hs3MkDm9yvP+OG9doljF2h5cOg5vKG4ClF6UiuPF8YVCS/rZsc9
NpmMec0kEJJJPSpzXmwmWpTNcEkA9+Yzg0bJ33mNbnswQukSzvtJvYgkK6H/Hwj9
ntMoRkxZ8cepv4JVenrk3cYAmLaaM8hvwhz8Ecg8UphR5cyuvLN3qSCW7yBWagU2
j24RjIsmAW7EnAPHZViXJ9iok74KBNTcMeObMVJkoiHepnOSgx0UruT/oWyhV21S
FPH+rsqrOv9v9OVB5bhM+bLOyxAIe08WIZKnnsmYdwR7KjQ6n8Iu7giZGGnpXcNz
Ljfe6qv95FztAojIGG+8aehm1eKdUKs8MnUGqaeNM0OrqHF0X0UTNUemEo60jbuG
Go/if+B/6HcccnmHUVxSVqcD1vrJ1oFqRWYPHnEOymQv0gWdpJvfxF//pZWLTDKI
NZgAacfc6WYQXh84YizXePM8I52bC9i+6dME6ZdkGJjWhbQGF5m3I8J4DEbQARkR
H5yUfQD6pJ2S9aXXhox48Y+z6GA8AM2DVjrYXy0Zn3rLy2OKe/nhaluwXtBfV1G6
ZYjW3/vpXhpCVsTktm/qcLOajpz/tZPC5qvGNIKdbloes87fjy/98aVgeqKNzMX1
iPS+gBFlgqQR4GMFtBQ32Bax0Mpped50rV0M8OHyNIbDbjtMOKpRjKCRXbJY0FGh
FEVyQyW9f1kS+76UBFZgF92eSfVvS7aocNF02RxARdBYPD/erRoyPvvXghl08RTa
XTdbnnnb/JD+tvzDXph9J8kJNhLd/5UOi846LOFWrAEdzkkSA6PLTrS7qPHbL8Or
P+OkzL93K/7THrfB3yNxk4SQOHVMMM+AacjiXPePmgkY6/iAUULe5t49QQMlDpMp
BcztiEoYKwsY0B/+QfHdGLQ33b3/97+1rohNj1OuT3Wu4iNQyOyTgTg4hj5kZeqP
LGajqcAuiCh4bT0bpfiTaKBPGuBTHiouFiaWAg+CzUlP/y5iqVXjk/n8bw58RGU0
MWWo1gtJo3t+/odr6H9b5viZrYwwLRHqLR21EGmMbjzP+gyzv3k5uxrNAinem9r0
TjQkdcfjEvD/HqApHU8ku6ZcQfGFuaI1Lxi4ggxMUhIFwIEoX7tCFi7yrreNbUmP
NqTExNDCiOnjQSybQuNlqSjgqzfBFWvvaIouYDyvdUk9z4NATLNQAlnFVPa0EeUi
CgcX355Uvu00tRx+mZ0U1jFqwbNrKQol0dqkfthfmDN+oa/AF+PFit8C53rx90Wn
bOalhSJUiI9Oe+fFbaV8hWam7OFsvl44W4ZLF8EaugeukRIPSI3jdKu8wgv4tfdh
HEkjKPGo2MV+oeatGILNTq3watG3lE9qgxJ4mXnaWyfK2k2yRswUtq3dCz7oqjb+
9sMLFFfrWugauYhyQCQNA3tMKWDA3Thm0iHgfn+78uWsf8Cxo/hPMPng3olapbcs
ARPNF9N60whdwKWlb+m4fM1rT5EMOrlkaMkkbUr5TpxDD/oUs62FhvIjzLZmSI4v
eqxLl9HsaAurYfngls9wWmOyM5IVvzwD1pNsfKXoL2FSt3yUCc2qCuMZ193rhWsO
Xpht3w2D5HPSrcU7WxadfMNDoWpJSCA0Ud0zbQxJex6AwVa73PanfAfCwcurEpZs
OvK6Zl1WS4wTG0SdE4pP7oodhh4ZEM26lAFlCbz49c1JQbCOI6DkyF6bmsTmdBcP
ubp8g2VEgV4LfJ+KHz9hmW3L0qcTvyT50B7wuVNSI5bgeArkuwwHHz92WwW9oKmt
+BnrJRS1gpV47XL3bhAQgjsDwrUzXT/ybAiyR2gbfPO3bwIoo+qH/Kwmt8BZnMWE
h7Ey3S9K9kWcuvX8VgCTbN3tGp9n66mgiaP+ZbgPCHGVrq9iAEiPR0iEak1rYkwM
jwC4vf8OzhEF/NzzBLjmDoIEZsw8mzEV+qPijGwYdYQwrPK3UGzmyMPWQIIwzLE8
OLEsyR0W7U/e0PoTnmoHKS9RDz3GmSeBAbxkBxh1izppuXJfW/2PDHjpYk9/HI9O
EP8iiJS9Hn59bf29GuvyQGdX1Lo6xkCqfGz9OXR7L4ooMiuj0gblEjXMg6EiTETb
B2Ax3CireMnLFTc8zKcnjH+IX8Q4WV8Wol2jqW+rDjLbjMyOP5/m6/f1eQwYvtjp
m49mntk/OF3QjJiG6t5bpw==
`pragma protect end_protected
