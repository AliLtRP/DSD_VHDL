// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
bPgkAxiuKpu4hBe9CkvWAaHAbxoa6vgrRazEz5fzQSJ9z9Bll5dB9jEzMzdr5i8HzUgncA66J32Y
4Tif43eQi0IumFdGc2APsySPWczuYFWyqbxBwVE1U4OsrnyVEJVMYWnprgpZTfjaAmT+sZRQujjV
nG+pafLP8YBIsMUTAGOombW232xXsPr4DFY7ORg332AtfSEWM5Sn0HeoHpHvTbZe4gbKxkaULcyA
axGhUCt68ZzrIO+FwsabRKAVZPxwNBMKR65TRN23onerHZliS0fxockUAH3yzD8rNDGsUOaEsg8v
aZmYts12A9TTyxcwH7yZZsEUOPDLxkWnms/t6w==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
eea13/uT2tnBpZ+OxpFoKpQLg0Z4PPT9T8WADYll6lxwP7m/Ylf+aWmM/hvEgxcUl2FRCzBm5c0y
U6cVyncCWRJsRlGm0+be+8g1xcNTeJ6LxKK8KpZ7xcF5aSJERb/rty1EAaayOvItow0CwakxPVoe
/Rda7QmMfbc1RjD+Se1RzJY8rE3Vb3ac+Mov6kU/f+0f4QuF1UfACyXaVkn2qiHw111bhGuH0jWl
1X4s9pW9juullXy86X3sNZrdox64LHAXgsGl4wZG8PQcKAKq37f9eLR3rRCbfP3HGybG0QlXkDuq
uxzxg8TYjlHvMpCrRm9rz8JIcDz1jvgAZaSLgcLoxlUVRnFLuJ+jgKJr+ZMIg/MdmJ6oBVRtSWSV
5ijad5w+OE6lHB/uuKuIxZDFQ01cERVlHtzxUIdrAWPJOj4eanK49e16HD/dGRRfgXrgzHTF8ix8
+qNCjvJpMxitwKE50bDZpVGmjZ70zmJQlIyUAPIHeYggULKb3/9MceX4eSCQMTC9opbq7z2hRRW6
AoXT3HjRPwL2SYpIYOHGqIPFEXQvZ2EbkWP4azuwIs8r3yRUrR44Y/OMvnR6wygi7BIo6bxQpKlQ
i8IEWvhYknDv+tDVCBA4jCfo2zKf6DnN4JPtsJKW0Qm5VpHzjr9Ng7yMxGqqJ82qAZ4wEC2bMDmm
UKUsw8bbqUWrtpxvJtLAhawLzDXW5znJ1uAbgsaaMPbAEwgZ9RyFCvZMs4m/qIkKBEG+kfBLSYnx
qIgzKw56pFSI6mjjOC8YeUdrq5UWFcrslR7lMlafhqSpyBAKKOW7bUeAsKgWKvHvQY4Z+5ExXs0h
kwImTauWpieRscGFPYzz5BrnC0D/YW4N1VfPmrlxPSMdaH9x+qvN+yUyyW2Mb81+lkF4IBh/YnUT
ma1SsQeDo59KOylTHYWa+Z3EOPSD9y8wJZDYTlXN+0omsHWNGS/dTLiwayiO63Q9ODXdGYYhbBQq
IHI0xYks1P5uGUxOu+sb7lGWtJ0gExpbtb3/RW3p5AizOC9dsRoxeHMj6WB66rcb25zYSjym5tVG
sWg7tKVp5NylDH3ay8neKkRL/He+SmgMQdqlhmuWqdpQ6Mn3ZmJoEUK7v6PhPH4lhTpMgl+bBaOU
oTvzJ+V4+mUlbF3tag3M9nigD9MWJ9rzoT7NYkG9TR9gAriUr0bNX0Iou0mDCa6pgyEVC6AVZikb
ubkiLAvks02Lzx1uIPxcuCSJ2+fLRFOQQHd8O7F6Kkue1NHuyOHOiZ7snL1tlMvmu3O/9rBS6Ng1
+whTXcXCBi1RWG+thlXVWUPCYHdn49f7Zc04Qap6ofLTMwWtbvdAlfbscjB2y/EYX8aI4vTJI43i
x/SX6NEGeUQcxORmqTk5A2CYrTHSCicNtZtHyC3iwYd49J+0Us7Xx8fQF1utq4d9X86aWgru8Wox
425KnOV1UtWEZMC2a8ncdO7foUyALkRuJ48JXCdmiLMPC/uzv+9MX3L5Meu78waZBd+SSSsYqaVR
gP8vsDV0LzyQOGFoyjBvERNadeeXjEnXXGEjY6jNtdp8msPQmRGyaYRVRN7LfPoXamWEOBWO468W
9dI4Ev81Uscu6r9PawYxvVHF0MrsyxkZpy/eVXKZWn7aiHOmdJv6Z2uFScgB3R53jEiMSGyLV4Bp
DNilpHRQsHdEEgRr7Q9WTCXz/sULqXBJMubo08cG4bGeEySyycaoq1qrY3zXtf7YG72+diKoKWU1
ai6MWeBf71dBPvWcZFtGfghZ08f9l84hcCXGOPNbqgQreHasnCC9rM+EgH6XS1LzyGtGZzPM+jls
vrsItUALGypKvpkI8w/53kk3iesoiem0S8mGFBkPYKiMYx2i2w6RuUaRVro4uEDw2ioyKKkaKbG2
5lGNufAshiQOwfja1nl7XU44xrWaFq5fmSd+7kqtrc6mmrSKGV7KGcDT8G2Ln59qs9yHg9b6s8p+
RksPSmgAR5heVSV4cYRQs6x/PswB1gvtJ+ligzy5SzfOVir06sWJESbtTtUbcMfyt8J0gWsBSr7f
RwzuxDkfHdrqWY+/dXOtvfxy3kRnjp/mqmrVHXa/fgb/VX7SHMacvPzKaLNNYetFP2Zve1XbdHeu
jLkeAk8tQm6foLc2BNR4YjJ+BfegYMqMF7ppUmqRQCCNBFJ07cJ1dZpOh/1u8TsSSdAvs5ev12TL
fF2SRC82/uzrJJ/PrcW00ev/JI+UjsZQc9D0XR3OS6DGok5vF2uUnQTuxw/9acEh43HK/JWKKA3L
pYVa0WdZxGHZDaThYYPdtCGcythlpyCKwbi/i+IxbFKb3lu0Tk5H5+sexpeGulhSgJlJCHtN3DCF
/uFvPvp5sCLnln+J8YzvE8xxYyWST8BdaEOv0ETbomCH5Pxe2MQsCW0yrIMCGnNfHdZ79KA7h0Az
7mxEp8CN08q9K/EYryD76kePin9nt9ASMriBRiKWKjO8YVEnma3+5Ya8SWpz+eI6exWhZ49u7mQ2
kIAjq3GonagdLm8sGJ2I9m1mRullL6tCisljcXKklJNXR/Cz2Mjw1F4nIomU2JYMYV/1M2GXyIYU
jmTiIhPLpeeZMBKK6mtVMh3cmLh5iX1wFi5hZpbaIc0BkhuUDJWo3b3H1NLdj8WVnu/YY5YDMNmE
U8uRQZ24UVt+fdciInyldG4ywogu9WbDx6334Shq/0Nv0jIg4/ay8fpoNpFWftYDZpyGZBpqGqWD
b01Emw2ySgVuDOL5wN3lRx2bRMKpn2HXbPL4u3svIA0MUKSNPojI/9bnE57hh/XbrCCdvHjryAdj
rMo1M3+eYId1vmtFex5oVydxDwBu72CNbCstMwounbWQfkntnk9WoeKOZ07jLBfr8ldXl/8LJfDs
rvYdPcTAJkxgpFW5kLhnetYKi9QEVh48K0/NRCWw+JwLRWhr8kVP06lk3bQXWC2QMX/nksZBm9K4
QY4Tai+RHVO/uHwolEOdLFV9v5hdMMYj7RWRyO+BAdlKicCuXtiPWm35npJHAyVRbR8ttcQ8F+zG
sHR8Nfz5ywj4DVfA5EAVkBJWwjEOORK07M+WnViM3htQW80SAQ2MhGMn8bVFMfmrMj0dGDNDF4kc
xRDL1LCsJg+0goXCvsAxUxc6CaBsX8GHaslxE5Z7AKgfxp1o9x+Z44IM6uzV7SNFw6hio2PCxJJf
Sf+jMghvpEM+b1ap1nGBS9pzGM4vxIgShjpXd8kqz/IqNGaelk3TOxKb/6PuuR4ua9Wa1XOL/7P0
S4blzo0mgoVsDPjjvtxeyER/vy94MLrMrH5KC08HSyvEMVG2HYWXVYPXNKCxtsg5Blxxc5CZSg6t
wZVL3f6NLUYc0HlHG1XWDu8+6jczxCot9Xr3Orkwn59nnVFcpvGCtHe6Gb46A8u1SiFCamikoX1N
/yDT5fu2s24+WwB3a796GHB9a2Hgbk3T/qZHJaz58buHulpDGli82F9Ihhb3wKrGhy7s6f6A2CiH
geMRa6Ypc2FpSgZjVZLPuZW1pkIIW2rFkZgCFUHzrdy0W+2PReB4GVix2qnYT3O0GfSaq+yj2mrB
TQmTlYYu4QtLM2ON40AuLcgGv/xQColy1Nd3JhGKtqcgc/e+kN0QpSxleRdaqfePTJp66hfw6reP
H0El4gtcODmL/aDAAd3NJ7xqzXL2V2l0m2/2juTg7PO8Vck3rRx3Fst5F/FCZmnjK8NIzchdAwce
MeKmFsQPwVt2W+eAv/CLgKOQJMChRyYDbOGhDDGGgrWGpSNAyGTtAMnka8WPGxum/FVoIzG0IEsS
5QLgy2tZLZK62HjxLaE3N9TCwCtUsM62JXy75/iP/94GuwRo2En/5PJV0puS1WPfqW+FeiAtGTkU
/mXNmcAvqX3wptuSOnHnD59N3YVyoIKJej6saFKphB6dkbnEZChX8pPda3r9ImsggVuA6q1gJBrs
557aYq+XMmYax4+1Ph6dWiUZ8gmC/F2Zd+PFNsuVMmSasSo1ttIfEwBQOPMfjuyiygjt570zkxmZ
T7i1oktELx5nG14HjpwGIPWFAeMPwfsvW7QXoqSE9KWVjr+zjqHTmKKK081o3wlm0RH5kwkbgj+Q
dU80pXHgiugNZRctvLlJPmKQ5T6AT1MWADtAH5ri359ilFp61UaahBWYfnSkdpQz/bgyK/5xE+iy
rF76szRtUqOWbPalMvKpFViT0c5UU5OrS5XTKDx8m89T2lfFDTx99JUaH2vE7OH54Qf1AuLcT5Lw
IuE4aKpjRnoxQq0IGEWALDJ08fkyeC0G0BJ0UmjeWtIBQwTPfz4/IIh+BGzD3YiCxyuAQ4Y2hmSb
ZAJKk+kA8DjvTRomju5q2xPIHLt28L6/qD/q1kH5Q1FpqBVWdKby73E4QFOKxEZ7ToVh2b5CevyN
ui3RXe5DVGeJ/4bN/J8Ub+541U+r+evTnXlMFh/nXSZXPhmN8WhA0QXYk6i03aN0c4fN+9ybB6Mm
iZTawSo6N/7LnqqBpkiWC90nyKJ8/iCoDLNcSE0Z2K9mI0fOvl9qMOZ9Zvy63rPERyvYmIwEiwi4
IKBG04clpZo5gn3Vplwi5WBqmeZ2A2WKztfoc/uhGA78zcEerQkTRXFRs/BbnD7c1GJ6qdxfKWmc
vKWfdsPWmcF2FDFOVtZf2peUav/1vHUYq6sN02wgAmYIuR7EFM/y3P1T9GGZ2DDcenVfq+3Bh73L
q9thiaWsZyE+HpkMtYJMa907oIaLqb9Z27FQkj4k3nbcp1f5O7q0xDkzCIVnNZe3C63Mf0hbMyoj
Zi9qSQfFOFaGtu3toTs4w84rfhZrpBzCEw1/Y+pI4Ug2Myv46TXXoqlRTi73LKIxjN/IaVyXlE9i
0bSA40zGQhr2yYNOQpzAkXr94WmTDhhFQJgpzjuLcXDOxK24BzjCUb2H3ODJXsTfWeHRKmejjCtg
p+Ntq/JIFkvFH1FfZiEIWSqrHt6/u3oTP+q/c1phHwJsy7MiwUsELCaJVM4sycAdwzWBz22+6DKy
zE/40fwKzSjkIREu7uPYX7oSSoF5X8iJErBayJ5WhPI6DbcZ6FKlHJI/I06Z7rUOZifiHgccywtZ
Ktcjm1xkQ5KWELBd+MDVec/PzjziwoeFo+nXoxc2WYrcHfjgVNvAPfqj/f+CuEAbXlaI8Yq9ygJF
QQIc0dxZ3jtS6XT9b2BvKturEEYcMeNRFZKqzfR05Xkt3YpjXsVewNCYeEM/4qlp6xh+eeJRvl/2
O6a526m7dEAjQ4VCHEvMycJuw4uypuoVGuOcyP/gQ7RJk9pS2/lTwv7eFm6v0Au5nQ14G0DXj3uK
cEHxDZw8qKZHjecI8zORV07uMYPpxL7uz7kuMLOAjsOSg56IOn0Xw3qvrOGrQMW95CbFq/PChy0g
fK1uJEmIiIL/uoqtLNzAF1D93QNBziFmZZGhC8mfrodNW/KX9TLLxJ9g+8qdsLYYoVAuv7HEYwGz
Wd6szTrIhea9VxFbTatFBeGeXOsYTo8zKFm3Uz0J8vckvH8245lVN1nitdNNL6qu7drN4vpjpVtX
+47iIbWVWKf/iaagbBroY+rvawPMYjnQIcmTndkiQ3FVl9KTExlGTKmg3oGSo1yhbdEbI9IXuEZT
OO64k1IeMCjT3fgz98ZGhHNAgFl9AfzUNHzqL6k1e1UQzC234V8O1Ldes0XxE8TCxvIBF+dHropw
/aKIgb8H2nmakDzFNVUIkn8orNJ6UFtI19eZA0k2KZs9zYaNAEtu6cWQSBNJ8Z2bxHdk4bcNCx3c
lN8evJUNV7le9LdwF+BQ+8cSCnF4eVV8dxibe9LGC1S4SZIh6U08Vf6etDf4pPj/hmUR+H8Bi0b6
6DQSAUFzq8xBlvtQD6O5NquXeBp5W8cC32Mj6MPlj97bHU6LppuDps98pe4ui53adicIlef+yz2v
CO9sMmOp4621og3k0Ct0AI0w4jMT8myeP/g3j1vJNehDBJkMM9fPyUEYDbckwBCU4gLB53rpe6wB
CjKPnoKJUZxbA5ayFIxk4WRKEonyWKHqfZ3H8zF0xFPwj/fzG2/6Dz4NCf50HR54hKZh7wscS/u1
lUBrsnVOE+Cto3tQmwjmiyftNPfLuxVwsEEHYE87NcVdGZV01vyKzwMrC8AMirrVXufiIoK2wtKl
Qoa+N+c8+MBafBy5iyDdtOMEQC2ZQyZDhSeBCCDpD0wBapMjVnXoRgidphkDZbYhMYllFTq/kUpf
i8CNN4OakIuSBRPYxFN92WKeOiCrh/91nYKVb3XgQsv/EVROnppeukOJ9TdrXNu9EP1tTvc3djAl
Ot4xa6tl/cWTrSeXgGYJ7IMptNP5RrhJ7/UPyYk9zBxXmd23t0Sih5sEK54Mw2zkxrNtSULPsAsV
e15KsR0Fk9zusY92lZLMl2pZoILmRPkrsv/Vdzafk3n7SUw64do5FKVaT+th1oaHKxuK2kRVjS+v
xhUUX2QFk8TtfoYMMW0ft1yVI66UI5KdrTqIGcFHFg+rDPm5ysVGVUO6W1EurNVMlCVisz7Ptq5S
8nckbu7QzfQqiKMw7l+zKjv76H39Y2I7GKa6K4g018w6HUMXP7hn091eUSfLsEKE9F1PGKkvYipK
ysPBqlk0kcHLbFd9araA4Rv6LOksoTS1I4otgzf7n8ubc/XYhDvw+1Jp1VyhLp5SI3eNx78kB/8m
Fig9H0fGRYUf2NMK5O7DdIGdqLcr4Gi1mccZ8jM2KFeO0ZEfym+74xHvQguy2ZLjzxHBmPo5ba7K
b0iKI0k98SBwzxGETeFzHQ0PdDXLJhyO5Fz4h8WSucOYwZdjE0h75Junr25YNtOgpPfCfZyklQ9y
H74IPFUVzRUIhjfGPis32r1xQiTKxB2pNoG3/XiyLqyWOCFmUXpx1qy1H0spRQXmLYCDWvNK6OPJ
p2n4KNwg/bqb6pib3P7u9wAkxnu56xwy2MBSe6+M3snFCVu7pbAPeVR5fu8kaSN/ZqWojJaIOCHq
+6o3E9qP6/q1udZx92fW5GRjosRAoD2FOwfjyr/85cNa19rCkNz+pxfUBFSvlZ4SxFJGI0n9yniF
12etn0eT2PcZMjNNAGL8oZYlXlkxaLDVUbLz2UY+KozB0jmzggjiOqb9/HmTJLszJfcRPdXSmJdY
yi5NMF8MWP0ET6xzBS6PjbbilZd5XDT4vQdMvg6bpHY82beINRnHG8IRhvtQ3NwIaAGdt08yc9pn
1Sj5h4bHCFuzJQeU4KXc7J6+ALCDkX2Pvslh14XVtOvzPCzVNQs2AsRiwtKV2hDkWWiwFlsABtuQ
REnweEOEFdeO/bXeiY4htgq+Vj7yJcWaPho2I1hz1zVKTtKT4sxPstQ02Q8p3+gNmn5YRl0mnXNG
rIlzNTBR/CYdqWGu4lA8LYBysU/YJ5W1mF5Saal7NOZ+B2DMqlNTQ2tEMZzAfTiGWE/Jg8FHR15c
CtMgSL0++Y21haXoMPHK46LAbctPaAqV/UByqWgx+d55sAv1HgVjjhTUSIh8uTIXehef00qj/S7V
O9nw9z54wfWf3Qh/K91cVl9HYqOXOvmNX/HucWEZ2w4RIWctkbBz1idHQMXF8CuzDJYw0hGag2Ax
D6MA17ebogbZDePmEgkPU0//4TG9XHYho0Mo2CqcwCbFxhxf9GU+mZXi3i3uuYPBuY2N/nj0AtCi
ek3bJjLLqfE/4uGMIep5UG4ymwrkL6KJmJBO+staQKbQV5tA0HmSuFxrtgTOKPdy5VNxUxUMGWop
nhY/Sq7L6b1dz4xPilQRuBmwhyCIy/IoCDVAVk+ERK9ZCi2Cs/15K4w2HjFy6ZyZuPJMQ4EYl8Sc
DtpCOKQXWaxeVOGIIR1eySJcuscfYD1gkGCFkLtisBqc4eaiFddjbJv2l8gcrakYYN2FufamnuYw
Yv9YXMaEsX6L8NQiQ4tmdDl7iiho9YaGHPk0d8EyeRA+hdPb6/LMB5dq2uIHz8QlVtP5MuwYuNCM
6eP9L6nHoG9Z3YZWzTr6yQH844cdANFwu1N4+T/AW+xOdb7nixCtuFz3c/lU8IVtrwGkUsxNLPmj
l/Zr8V9PQVnWYLQKu16fY++7P3b3+E7KsnkTwq8RkSKkqK9Pwshkep2PO+wDcIPNWyxvj9v0H8wT
Ye15YxSIvK3gy/zrJdXzxRFiAXCToMsUmeUN0cWgXBOnbw6njDFDL+w2KsQ52fgueqLTCNK42aiK
VYwQTbRLEyS8YNs6sOPB4vgKe0og69PZCNh1s178PZvyP5Xmzn51LrdLyCnTmoNSx/nB902WjB+P
fdSmN+TS1+I8YT8veCuzMFeIDtPzDyn+Pou9UIJES3gtDiGKWT0TDn3omhTFVTt972odfAKnJhb7
SIAM2DhgQmRqx7L+NLqrd6NpHu18AaGUeEu7cKVaLIZPaT8C+HyiKCo5cjVx7dJ2jAqN1FPGC+3B
rfqsjgk4yOUX8cdYAkB8S7YJhjumo7yu0sZsEf4E4fIv0dBzoVO4RPMt/54i3agybkHZKmRLyD1b
+d9ZjN/EOGHwYBY2jFilN84qhbT+d9hnal+KP0/PF1JcVHI59mOyq//2JM/dUMFl/U+4Sr+VHbmj
j/6gt2TH/XOR3xOW2n+2pQ3TIUnFUiVYmEV4of1PB7vjfxTGhUhlXRlR1LOASkFn+pQNAhqmSHnF
4m2L5IKAk0cQEVMg640XeUS/wGRpz3d/yNpgDJA0vB3KDf1WASLm98zYo4tnG8W3/JF1vcNouMEJ
6Bd1yfAcjDAYrCj5gcbQbwGJTiF+aukXerOFAWRp4yCVm5UpuYMVkoC9JfYClpXP3Wr6TuESNZTV
C809fYFDg2jVFg/Ya8XSIz0l41e5BnbTNKCcPqOCdvMoCtWgh/0aFI2kdwfqdD6uw8SCh07dknMn
G/PzXQkxfb9hvp9/t8wJ+KLfWeJOs/FdTJlFwtcdV7RLGtxvnjIKmCu9MlEZrOJfz48kmhbtCvBr
ItM4yZpkdCLI5k3Hbj7HlZpN1SOCxqKofbt/HK90cq1GJj8OOAexuD3VTI3/sBktFODvgCagaALy
t1S4ruRmZGecGvZB7SEwD/1BmHPznzx5b5mhvoxrkWmJwx8/tO9YEqlJhDntOB+cBVPJqXKdUCWG
6cxwAMaw2i2WqujKrhL+zcfK5m7UwyK7Pvv3iAdVF9nBVH5gRHd6MZa3HJzKAeNV20gCdVBD+RQy
Ie4z6EAlgJAx6dHCz6BwdNkZkdSvW78WyNFVDG8hQH6CXYlqJ1VjF4OsJGXL/BD9gDkHNtHn3NV7
O1/z/0A1WLF5Wswo58hoa/v9OF3IPy8n1zDAgBbbHEIMl24rhdH3aihvCd1SrQjgmOUt/GalS25C
FrdufwRODKDqyTS4sLqwi/bNNr8E1lBRfW6v1nBbBZb+tTpgGrlpIQPDVmIdOQ8mOWGLhrKBBUQa
qQW3sqWdHIdqBgZgPX/Y20IoG/ghQ8ha0zqShe7GBZJ2LMY4AKiX968yhdL0lwjdonyExqz7/otA
reorHu8KfMvqbLSPde8vohTIqjnRIHvIs7wRsm7e4j1oB23qQU/UvgvgFM8GeiDDGIr5pfCXgUHO
CsNJ1o1Mgg1a0dOuZbzhs73cVkeuqiNHryca/PpDeerM+Ez8PCzwLie6uhqtpKvFsyAxdgxb/jzB
Ld2GdH3zBOIk2ojj7T+X4AwJ8jpg0Amq6/Ozo1Unzk1fJE2vYHaf3k5tE5tmNYx4h1J9vwo99+cQ
dSm/UoYbVO7Q99g3s/cuoR8CxL9IUuNx38jn8HnJYCsj68Q4MIGcW7wZTpO3xdXgmXfAtrOe6JsU
yM/A6RAk/R5FWPeHYZAFx81WJY5Tvew+CK0nrTWA4EvKfDOQaJifmzGoj54ikMAsJuu2lo5KPoR6
S1KHUIkREg45LBVwfV89NpDcX/D3Hh99cHCM1zhgr/M93+UEdAfv/0w1yVzJKJ4Fba1TYcUuHXpW
X8kCFv/GjVFg0x2jA94rDkC+6Ar3Rrd3YQQH6mGOy0lIm6SHs4GPIJ7vNc+SPt5yp4qwPReHH+zk
7UCTj/NdZKfTqyX13gHVfXJkMt875lC5guIzSOBAxjQLO76IFf1HSe4LgQxijwxDLI7ZNlaYqFSm
p8b4Gxuy7wdRPJGOwmYVg+v5RkxbhTV4oQeVovP7Pa4MjH9wT7O/G1B0rNCNKqPRD8mZo7+aUx2u
x0gZsu3JJI+6b6nfjM1MJhALtZZ9a5vd2ZbXPQYJf95LNkI80gqABnJPWJWzzUmrHeb2fuOx6jKS
yW9OrASVRTe+PfeI2H9oOJBgrxAtB3BkKKpiVvAlU5mqcc+Fba/rCfEOMrzZhZGYKK36IZIOBCNq
nqQEBG6TwRXjpyVSZ1NVZelCuiSGQAraEzhYp10Lzd3EvR8igaDJT5mV4DBpoFfy+INm0FjmBgXl
8Y2AAU5KNB/vp77skOUiAIaOpXx89mv5xyTyboPxQ+wZY3KdHwBDYGe5STKk3ydqXRdtqd6rklDX
JoEBV5V7D4Ko8oQ5ZD42EjdDGvhSoeB3uJBgBElIkaMya391/eBkODropyodOh6l572UedJnklvp
vtLgRgtq3Uf5XQ7QmvvnH28vpN8kJzN/4r2FO8EheaQVh8ln2/GBY4oYPEp/xoUbdGTeyewd27dz
f4MIvHLI/ViVAozArKRHCLXuWk9G0xrdw4oZDEocu9RQMg+LL9wSOIrvGqS4VGUDr6aW7cmfh2tq
X4lpWKrRKrLe7CZe9dp2NtWr0yqSNgqJ2MGAaedjvW7Zeax6ujYucEau1gl2hSlH8XGy9J5BiRmr
4knd0I1M7IvsrK9JEh6Aw2402aRICMx9yyi5Loot7y5nwTQnzXvTWour+pzYdPOVpd+qrIV8pY7U
JczgKOMGUWt/iBVEtrb2nyBxedQFtHzoRqB7tJVgyjCB+n0ZlAy77fSaOPx84bL9W8ImV+wJ9mgX
DzZ8Wk9GsT10Makezb/j7z8j+kKwJRIbY+ybs1rI435LGsNTbxo5SZjY3vvLv3DROxX08dGPUe8z
AGBVZbFGILEXFfeRS1OXhNv9W8IxORqG5FcacF1K6QO3Ju7yy+0iTrQjw5mMhL3ZgjjQmpgWX2P5
Mna6eNFu6SxLydOtzt5FJGdg6YuTuNBNGzPMKZ5w7Q8ojGQ2n16vQNy6RGhXemaQqn+0kfjElLPN
TN+28JLvSC8aSdl9/7nR+f2qV2TLBHFOom0sYnxoxyc5+exeiVN8YmfOsHZd3AHP8H7iXyXE9BzJ
L0egx1PLFJlKEF1gSbha7tlEgRYf9kGWlO4X/4xlOe9kv6zlnBPOZk1n2Lp+dXOhGF4kOfy7OCXo
55ny+LajKjDv9Ve+4qMU3AwBgUrEFHFwWU96ZtJMZ0XBaaLZxlxUQ2ul5Nq3KObGQUp1MPWvKLa/
WLSRqDonVnFwvWyiWAlmz5M474FjIK4KUvkSSgxaCF+0LWwdVGiGLx0owRXLpNiVL0HWbj6cvKpl
h+OJJBLNvD819U5aAvHIBzjhCtwXThAGDeFGOBqBqUTsXA3chHYT1chOenrZSpId9B+Y6hGA6idO
LdoQ0vP2x6Ff/UPvAr04w+Z1wBVVv0uGAloHMWC22J4SOCytJXpuRqLullNk1nu7iQiwYOci2it0
2HtVPUHz9GtKG/56/y5MgKwYeAyHFlLxaWFbHithXXkW6u2D6JZYCqSJcv1yXeK6mlGobEQgNZ2z
o9c7/TTrC5nRP6jVHJyHnfoveHJNCYEvF9V3rcOcjOykeYSeKf+acoBrTI00xeq95gzaETEqzP82
i3mbp2lyH5KTu/yEkmTRQf76xiVFMKLsvz7hEeH05aYbjNUVvV6ZwGNQwkyZyxQlBbLY7Myz5AHE
O9IMrOhTaz6RO85brvAbF5iU+VHHI63DpRqZdJwoTpSO00MsFSZIarikKxwEoDgDsUEx78Xxfnsd
8dkFe84qMDVaiymkcKEvZDKxHa4Lqzn4FdrprZYEykTI/Oe2hyE4+/R0clLCLVVqJ2739aW9zFxS
LC/FhGN3oLmFmoh9lOmoIzKHKZYAr70g1K1wK0+KgTvf6GRirCPlRVG13dzR/FXfRXY2m83+c6Wg
FmvRCyEI9LKFP1+u3cV6BgdC7jTe1h0AaJg/soHRgHCQATRgwyEdf7bbceOD1Z1d/Runi4MD/aMB
SRXAuYu4neXsHZTkl6E0sPKbgwvpUJ687AnFa9YJuNNivRMmaBb3Yo/gvclAaPBG0aJWMvctp4XP
NjX56kEZR50HmRBSLPF0Gje7f2Eye/zyVAINkuHrIMVT60hSrTFuqx7ibuVsSL5l2wEqcP/3FWWz
9PgVwfxgB38/rKAeYVfY8rvOJ0MpRnOWv8hisar2niPtLSsFVDlEbntrtg8dL1MlyKRJFDR8d6hY
Wnl9ZjTFoqg8tU+QCdeqlqWTRxRDfGe6XIyKFqmkmhbNp8nZbucIY1gYoDQbKexcye17TmWg1fa/
Hf+YxwMIP/p0DdsfW0Gkq9iHO8FznPioBrFQoiTnZsj/Nf1AI3z5yy5zTQIA2e3vFcewmCs3E+Mk
SBfu+Bk/7yYARhs1XLB+BFqItk9hVUmk/iy+whyPjU3vOjjWrDZg+s+7yNzy9uq+b3S2JovgMmZM
2D8noEZA3IBrKYhIeJgZ6NLYIkC9Ay0LY6wBYJtTzMkE5PKLFusEIwIJXb80lOrU2AUsHQeZzEl0
y7e55bRol/j8Y+A+t7txUEGxoPqHMbz1JGVpJ58iZSJPjnaAfuAhyGJZkpwd3QckElCE+gNtwUG2
+EJ5mx3tkWNNFqXCCvxSgmIvoGE07pp5vFxF8jL6qwqzu7VFjyKIygENGj6pQsOQZtiy2FEur2Ex
wnqOmDuvtABcEyg2LOHo2aGP1LTMXgAuSDsjXe4m7tevbmn9wQXmMiO5Q3/oR6ne+opYJeJfEwUs
7i7SkPJRWpsgu+BkcP9P6pIzg6SFkZHS/PqXllfsBMzuVMbBp9cRQ3rm584RorPRSViDVs+CyiGO
DKGgVUeL9tERKX8i5VLoAXZs8fXRA5pzIqWFmY2JUQCFchuXITXy3mjJcsUvMivGORcMuSm1hSr5
zkkjUu36crEE0Bb8NCwFbqqRY5Y8dao4hyrhb4ZdkUKpf+yzvlA4gXY9kX0FvX3mw2F2EUp2KFVt
T6TY0uSMSE6HvHRnYbKYoui6zVuDKthU3LH2nIDSWTQXetAiXDi5ds6IMLjiy7rzZc/DpQPrMVhA
e3Q5eIsCHfoefSVdAlGF3ekwmZuxxo2aN3Rlh9GMMHZXQL2NK+GG98P7q/LXTfMOHb8HqAQ4PYIi
XqJ5Byx3f3Ptf6ylk/sH7kGZqSQZUGOZOHI2Azj9/nhlBWXN98ytyftiuCWyo9AsbLhkE7CdZl6g
TREDl7KFMEOVJ6LoNHFo3IYjvAtBYKoSRvGgnc/OsYKqQ0R7bDF+aIdZJdAAa2WP8EllbSx2wuk/
2twNwmH5aJ7G8MBQ3mz9mbDDbz5lKGAJ8P+b8+T4Kw/GlenKepZeaY7qmw6RsjToh/lqQkJjM8DE
2ek9hlX4Fiurr1+rzVDj6gIlfXAaK1gZDDq9qsB6+HJUKGQw5Maw3jjrKJMvJbsQxyJd1vmvK+PB
w8RwTrlu6qdOlqT6NkKGbzJky4uLT/rqkpaZvKG3wPTk13KGvaHiVF3N6C9YTQAjgjm2Pc8Jmcc0
XogPSpu3H0hBBE0XieKbFLc071q0ygAxi/51GXBRctore/EuC1sFZOezRrVo3cVaA5wuoiNidf4G
GTgglBxCHsT9bC+/dnc873Fo5BHYdBVuiWyzdJRL3d7LqIKZyetBDxawfisZInI4uPSn1MtdTjNq
hcqwa4G1SLhFZxsGRG47x/pOFDkwfYkJvbOjyJwmJFEl1QL1U6VDZSBgl/3gD35Vg748gLpF0QnD
jJevzOvst2k74Q4iWYL8tJQ2qQjAsl0Iz1IHxlP6xTjH/EYV9cATXhojvPgbM9CYj3ioUlDinjXi
m6aYe0VNfNjomRL5b5vZUyiK85lImDVgHlVT4IyXorBzeCIBo0Fczc3/9vXIc++bbPipd1wNtgac
hyUMF7PG0/KgQ8ikovJTeoq2lRiJcEvec+wBXfLBbj2JNv2/GLCnRnsZakFLqi6LbhEgF3DgLxAi
sVPCicVqxUTFYn16bIQFHxB8Oz+3+lEsyAIPe+IhRnIqziHc53OnOBesbCbhXjL2KrqCpWj7iH4N
q/oXqwmme4a8AmDIrb8UbMgNRR3TLGb1C+SqCp9nZycax3/owSbfQkArK9r9y8zRQslyuFf0uLZE
mw4c57vvikgQamAEEVsEKKOap43N3yxTUqbk93JAJW+1PNw9O92LO2lYOZ1CURRsgd1TnTw9egyN
ylYxt34yNbQD/LFFDoSSR/p0mmIKasgr3TeaqCdfiAcV7wdkMNnH5sYxbUkP3LfEiNEg5pNXvyt7
TxY1gUC3F7+XkIWhgkoaBJHXSNHR9wqfXy3WOa6KljGMqa/KkRJl6itFBgPJVMkqOSl3UE/YuIf0
l7+/h/oW1q7hFNqJLcfjBU98zy6rdB3o3jUP0DxahB6/hf0i/QB9BC5dUFx7OSI2+SeAeP7yXnAF
AUfQW+yvgHBpn3tH553x/6URMMERjFcNsYT1uI5T1FmpKrWvhLzjEbQt4GKEcJrOlW2bOaX6ETVQ
SR0SEk+z3bPHCLkYymsaxeuwh43OgC8thkWyC23citi/U9P0Ly4aoXale5IGu+1OJx41bmKB8NU+
JJl5JeDeXjcHqmv27gcRN0Ko68A8iw5fKZA1FJCIW0XD0CV58SGrmB97/rYqs9ZUjIBFTnKCEflJ
XXqN7LmMdlVTiHKvj/WuBr8U5wKAMDeIId9vpdxYtfEi9+pLJqtC2JZENHThkWKu3S2Rn30FPJ9x
Mu5LPga9jO4RJtSvKCCLJznc3w5I9NORyCyrULmIaccNSvbPQkw1hH1G0o4t5thZQQrBXvPeqQ1k
BLY1mzOHdER6UWJ3v6EqT6b1aKsbfXbXTufZh3PdmUt+sO+z837ef1yJOlYbcK/Jtj6Vom/6GUC8
6FzsGKCP01SXy/havk9aGQXqC4588R1KOTs+fMbbHZ1brKyl/Yni6aDOVU4ulCD6xSNuLPyr29Dz
Qjta+0GqjhTCyGPzjz7MMNeOLpNiTIneTdGL/nRgINpzk+eAGcSw5xWebn5aqPOlvsYQSWtw87po
uCZqN/FKGgSaMjUViVDRf7LvSbjxbIik0n2OGC9Mep5Lbs8gd4Wc0Afxr26lsan70nCxL3oO/jW6
W09qDO9Q9YDUUS3Qw9BnTJ9LhJK51wE7yRd/171xrefGoRe0zfPheShClalBcksrHidWc1xQ3ffz
sRbYCpEfMt0CLz9jlgtrS1OwFGA0wyHMXDeaJc00Ch9zt1tviK20pb7Rrdh46vxvOv3AvNwQPowB
uFFPCdLxWReKnq8b+TuD/OXeKoO+p2GzsVibCawgcWfZjGPmuy2snJqz7zMAPirxFSxahQDcjD7B
w1zMvQ95d+/NQfAcFljSsTS47mJ4b3OBUgavAU742lHTsindIyv6wc/O4zPQCawBD7ArwhzBGOrp
GCi41B8QmFt/C1jE3ZFSUn3PnUEHQLiooslNU47Y4Kqe6ItOFfrOYx/2Ock8xNRfa1g6DWkawm8I
g62NGdks/9Y0DGioFs1ICjiUKQy3K82hpuFQVefRR1LYskAcpFDQPv0cO+Bv9UH7BxI9bzq57NIW
RUkh1PKw5CXdMJ/UlAnjpHOOvftbq4RiNpgz94HDEyikKJwos+Dcv/gQHEE1S4/wlTFE//+u3UsL
YAOEsSt2F+A9W5k5+kMvskyYUWviC67hzYZg+aRY8LSc91xsqpJ55Dvo/MlvQaO18nx/n65nSt10
55XjfB9Bvu2Ufg1XPYKfSYpNaAwse+sEKejKcpzcRaBCTkqBK41+nxXPDb5QUUa13KLPZAYQvAJ6
NS9HV6wUJDx0XEypBAJVhcLTs9sGQE+WlNJWWSHHUoqv7p6HHy3wdlbw3iRS3WZvz2wZ6p4LGmWZ
xXyLy2AfDVK/2kOdvB80c10EwapC/SuLCS0QBGAyTd+mzYDxFNY6Szr9DIwjUeMYh8kB4Qk7faZ1
9LxOVRZC9+UvJVUojZLs1+o/TRJwJdRW6QIJyqs11gOiZZZ2iRhF4j9suB6Ku+1KEPlRfgSNDsyD
r+YakvrPFnfOmnbUHFNjPhTjH83NMGSxrszj5Kvuo3GNT78OgbcrzR2KhHAW/Otm0qArh4axdQTC
LCNFHIVUrHFCrEZsLsL4gfxf2K03LGm0RSDcwCnz5jPzy8iQd9GO1MNm8T3KPaGsIvzPn1H3Tip6
dUjJLPKuhghLZq4wMI+7lGLypjE4K8SCk4rydWoS7hvfn0drpnOrCDhANBriqiMxIIWlff1ZR/lX
gMkXn5h9D56gWZB1rOcVEvRvoBVnzqDR2kWDpfNdLg0FRATpg9GoLW0JsW/Vs36uK7PqMaXUfCzj
iv96aYgE+44Z9vS5TjuTbrUzdwIkk4tl8CdGVDzRguuzN8kYxkdHKL49xWkw0DPPzLrYRLVtI5pM
3HG+/J2HjTy3g35Q1Q6DJNlOBPDgSv9jL3QYqpPZEw6Jzp1LZBgiowYjaCkg40BKZFU1h0GEL2vZ
1BGamh/kzgShwRm33ywAa0SxwJzpnAIfbpyUckUeo4PWQad2vlAGhwC9N/sNIIjFhuz2aCjvuiUX
lWHumzdsVMkHnSLGYRX5/H1L/loCGQy0yHRDmn7tNhgysx2laAPzKq65iAOdzM/FMsYGEaHAjB1w
iCaj/I6TdHUYLxx4IbgsCMGnDb3Thpz6lO88XfC3wz2q/GUVGtOOtrO3nCfkHdXyEdozE5nE2oDZ
sc958jZW1Gym+xXSnSFbb8+ww40N1hzvxd1Qzr/0q9wOSAmweY2mU6vhqgWfTWwMturGV24JooTK
OGAW8/+YNs0b3T6vNXUpNRKC1YY1BOJIPCO5/JP3N6bGtIIoR+vqgW6RrSJWobJt7HP86dNGQKje
pqfH1RLy+KreuavSvXFjG8+LbGSxf9u8Qlm+AXvRsnLPfdeGZcqdGw9SOL+ETiAFxG/sf+Gg4/aV
H6Hl+M3HRMRV//FbMvxcA9+6gwv9qiuzTYfZiA2ovTLV+YnBgu1fV08SWdSKnSLTP0WNh0m9AAHe
bUlOf+PdBgzOO0xrQHdhthuFzV92ni3kmg34EZ9D3SCvoZc6uZzi3AC/lU8XbFxRZWNHHw+tPHAE
ptwtX6ihuit0CJqiw9JcsZzrBKZZlFclBRF2ABh651BHszHyAywJ36zJwVg3hVev2fpl1vNwx10o
QdcXvE/PTHvcXlWSIQxR1xu0bZlaxCSDpnpGs7o2LlsQ/c76naGTFOWfApPhOVlKhalNobVGE0QS
18v8fqPIlBrX0oZhV5MAVAXrSd1rKry35ClTNiNOFIpVut9OaPkYyKUq3GhBXtY9D0FNclsnTEkP
4lhSRKRbAXsiOLBZaCseHBgvZOl8NQdI+DnqLk5L0UvMkT8qPJNdNMJO1ENtCBOz8cfcX3/PsEKC
JZtCXR5XhmQ/EZzeaPu3rE39MwLY/qXko+CPQjLDWfDKrXrriGDvhdfA3nPOWO5kX4lU6u0xme9w
ESRlah1eD4hrrFxH4XEbQ9mhMM9873OK02adKEbtp2P4YnS6SHm7kMjemoWGO7qUOsM9/P+97Hdf
NkliNAQgk3aqGEtF+uHbwfJovRfK5pj60tv2cluUQLuJ2j1EXokiQkWtuMf5oQWCMB3XNNNHhwvw
hagSx87QUGydZ7y2MR2jfhPNnx+rKwymefsNaZGCmglfIucRIzP/crU4AvU+Z1q0FMiM9Wkbi/Hh
WxpqV/h8Vf8AyYR+BSKvvd7zO8I27gpOZxLwRMKqgcLUQS1pqGWUrjiy3+Tj8LKdNJ4rfZPQ4IeP
pZojGQXF8eLG9bTDAKSOH8nbdp/2iLBuv1Ve8CcfZuMLwNH49ZR8M66sZoXF7vXE5/bL1z4IS5HV
ZG5u4iECGqj/HAY+WAuZ2lt8p9shUFE/651He2HRUXH+dGATAR3cn1idEdTkxECS+flWsKz36VzL
UK9wbLTSbbMh9tecNZXE+LriK9gN2F7YFEeoMmAJ7Vhl2XC6+mAV5WfJertqlu3fIFha6fzGMGK/
q42APdfpC/BP5x5DT9l/eF0FHqq3tPoQxJ1crrc5ZYn0wwZp7yzDh0DOk9nMutqcA8GyQp5+4TVm
VvJBs/M6ftrGJrCkj5FP3DxcFpsJNr8E41uei+TTfR1RNmikoQG6ukkBcXZG/PCvlEcObhG1xoC3
mWATI4yBd1ypl1wv2xU3XMjEOSojU87XU//F4UmQFNB0vnHucFM9W6dS/FDjKq3yCdz7+LqLQcH6
/QFQST9unliWb0hLHtj0FMk3Wc39stJ85aQxzbnjsh07bCseaoedN8FktkVnke861eF9ocCAlRPh
c73OTe/BmXUiXujJQteFWKGdLmSxWynj89G1DMKgy9LRVcnv45osUvCjZL71F2Mr0Q0PbStS5bcN
L4KMFc1e8y8nuB/F4drAzo+v90YIah/FIPeWXFA8CzhjuTRW4XEYf6vrj+C/h2cS/p4+la0xcPjb
B10wMOsidmvJkDCHzwu2vgvStO2gLM1b8mnfSZWotbtUZbooToRWGzB2mAy0cMhBAGLfdn2Kk+0C
2FEKh/U2p8TIZGnHfLKfOGJSNcktPY5kWCN7HuKRJoj6f3HvsLMrOifRqYvM1NU4ZTDnaKfEc8J+
zJPiReIyK15iJwQgSEUnytIMd2HFYiIg1Gh+kr8V1cKeqbS2nEDVZTnvODKAg/nCyUsbWOfZFCRn
hjQ2c3xlQ41KyTDb3Ep+88w0tOEGiRFR3Z0ACyNQXEQCNH8eJyaHsx7obZ8J87QRgS3j6tC0pjvr
11EsWLCJ6TcMrHPPrnEYVC6wML+1M4y5sgYPkVn9nKPiSR1CoVuIs0XqXss8KBbsv1bQYjUxieHm
g07Dq5cVA2ma37PMrUngiSYzdIYgeJpzDhcotYzypOYfNd9ZRXcPpiGk8M6h54KO7LJxFs3ohEO8
MrVix+16Yr7zvdMP4T5tNidOTh6nkv3pcxibfFqKqJmsL36Ji8+cZa4EFC0dBy0nzwbYeCrnUQsa
IZgBm42Z1le+k0T/6/XOIg8WwklXCPKSxLzpgE+ajaR6tx5MCcPzFlR5ku0a57wYCrKGGfjDQECz
qzQQ94AYgwG0b5MrRFsg/gRzDbmi5eR/IajnhbhNesS6qyMjzgwL2Mt6k91jR//UC/jUF+W6+VfU
6ME06doRHttmcoK5FMp92svAAUogQE9l/KjZQ8iX8q0PwWTn5Dn+DEzy+0pB7cT5lTNcxEqlq4Ju
HbL80R1oZUAtoqjyRa+FxT5VJdIZayhpSdX9EF2RN5BfpajDXDlswwcWNWgQ514P/eEIsNAn4J3j
Eo7JKRTkJcYRlV7IcQL+VFd+L9VoBVlAy5ky/6hTYZW9HTfH7RjDSqEfmgocxnbEm0Rmsn9OS0Ic
YHzhoxt2dwpJR5Bx8XkS9nNV6qVN1kJst3oVC5DA5oZF+4e0qBrkRtyXDm65dcu7ME4W285TmN+H
+TAPl+92Gt/nQcO3QW7rl/nropWR4Tf42G3WNNDCilNR4/mKPzb+YzFGi529MX1DsTssLVVlkBmi
0AQ0wkh9kT4FYtDd00FC2n35YptAA5Xu3BxmFLVO1dW08e8nr9c313iSz27VrnlsSJ2Of/GD+u8g
Q8iZRZg8ShyrkA/eVFo8zukejJZHthJsO3IEi5W2AFmAEwWye4F9BT0bHfvwo4GUXGCD/YHkk9NG
Ehjv3HqjjoQ95UKjS/1iTJA5iGAF5nwyaqkGb6kCvpKpfRiMt/miInDzWOY5ZtTz0QG8Kh5UVMK+
BNA7JroJ1/OSL//AIHCwOcwLAo44d8LBy3hiEvC+JVfin+XDKQqTj/c4oQiHrxsqsl/hECQnMRb0
V4MjVceSI01QuZjmv+CzkFStyuWyBoQRS7Y/9bobdb9wybSkCjqsKkHF30o+b5k4Hb2ovBvDkTlf
/6R0YH3csdem98K6rdjoCPFBB/TKXoiPgmlEvlCRJWaoyfYgGrwnH7N/icNRO0qdJ3lLnavmYt7T
URfBu4GUh/jrmNg/ak1hX0erDthdmE3b5IRhPxR6yzo9MSQKA68+++Em5u7hCi4G0IPlRHCB2SsY
Wr7s2VN80XCpFSttYz93gTnfEE8E3bVi8DAtHIm66zl8JdhDrxiK+/7zawp0gFlm9za3vluxT3Xu
VGvOhTKQSewl+JcyK0cYahXwBaaKEQM4yqZNEzJXNvEzcE+tEA74fb9Ay07v5iyR1ilrhDdP9KTd
I5JGx4r6+bTQQCyUtsJkebO6VbL5hrVzeHMTdjk9qsSYwBGOu59FQesfIA6mN6cQNeuLT+tkUSYE
uZyzvKE1X1akXXsEmmTo3vcD5Mh/byJB39IWAfWl46ec8n+l4+U/KOe5OJ9EVkkiqjZd4LOyybv3
trACSuJJ39XeBUCqlEkJTrEN5TPByMV9LXqxpND/6aApxu8dPBLhuHpo9Xiu6YoM5VHATLTFWWZ4
zEVk1+5yw3Cj8kSUcaoWgXDfpzj252LgWtgAwnmvRZ2SUgXNNn/kAdYPMa/k9XGHuULKLUDiVMAK
3om2VQSbHAf5n5u1fQXljXwBWQ0Y5rFHybMGgD33JtMRzjLQAOCe5D94bwHDf0pA/8Dy4e7Po6Wz
5skJmOzqFnG7UAm6cYAGWqY4DUq7VwE2j+meD/Lomv/sw6erkd/XFRmXMqPUnwIz61GsLLwc67kP
V8xWoIQ+hI3fImvJLHAlVIkV9RR5wPlEeicnTU8QM9dOuYHlMHZSW99H1TxG8wUYtu8QHCvqO90Y
OOSFakCUmv9L5EPnZeuqAuYAxEyTsBBnQgWeHgqM/Y/AC46N4koAnnc35SvM+Ls6l5qgoBkiS53x
pDPo7jy7cahPJ3ifqt9pnfAcJ9b4vrnwBejeuWj2JguzgpH9DgQN8PXdoNHOU2mHlKx2VYLcw3Fw
UomUn5G7frH1PX5y97USAUFcgv+/Q2W5U0X1a9snHxHfPPndYvZ+KPuHHkxr04dNNnDNN3XmTN0B
8TUGARqJzikmSW2f4wVzehAO8IRMT7e1r44FmBTOVMl2+CfOehAjOWP8p3gOYDF77FSKixJlhE0v
IJQ/QtsEgjHgnvYbrYzfUaCQXlsuKeBVv97d1ITPtZ/I8x2xtIO5EzS6I+izoUfD3VDp5rxrt8Bv
WmhRS/MfSlfBCEnfeuvKgBpsh9Wd1sSZQO9pog+7FNI42uSIV91+il+CXfFAS8M+rQGqsi0TEdRk
UcmXeY7Dw30hWseeUUDVSBCuUnUoBWyWVnMe9kg5AxFOygV3LvsHKLWQPjzRbxLrq7SZ6rGBbpUZ
Mf8BHHuwMB20yCknleoP6yMX2UtLDvrd4nJ8y6zDWGXlAEzgKrobRuSbM7SD4mLhy2aRc2UctOZP
VhV5qo6LrY3Kq0PaEDy+PHuSs1Q9nJpQVU4jBp/4TbpKg3uY1t0TDpNkdqoILQEfu5XTFS1EIaG6
6VyYYf8wjTjLSOL/KpcYdDbPBUh8a/wBaj8e5c2SfN1ucVlbnsSc7k56pOcfJlKiFsjyiW+RoQh+
qJTkwD7AGummcx7UQ0plO+R/D0AjUkT/FFdWvJF6nfTOG3n8jUhv7kufl47j8fYKQz8CIOZln5ah
6TMP6BRDOZNZ+5oMc3lnYvKKzc5PxrNezlV9zXs3jIITFP5WI9ZwzQeBeXfLHrOhLLtO2rE6xscD
lMwwM2QRF6lzyNIEQ+zntKiw6aLkP2AklTZndrwqhrodoXRysizvQz/RoZsDAsMst7u92rRmMDq3
66zZHNnZP1zp6E2Aijw4GkUGpJEWmcEtinuuP6Y2OFjDSA9DZX+NqCH+EoLVvu+Xlb3tl5DhztN+
+bbvfHuNDKEHZDlQ1dUH5TDf/GGps1Cvv03SXxrUT8LB/CbTUKYLEJIgPmHtPAkDIw+5AFviRHaE
J/E6uBauKGr7EZ3RNwtybjGywl7T7MZBziDVNDizNm/5xjO56HuP9ut/kx2brP2ynjmclV+hpo7V
CqGBOWsUUfdIjjVXmwUSDLOfb87jdt/93zjx7QR8cQB6wkOAY84z0iYfGznunoebi3B+DTsBMDoi
ylYwj3LcHc1ZvRYEOeqHCpcNgXPfjaxMzyY20C46B8TlWZ14fCEho3+ge/H51LJvQKJgJNFH2Rjb
gtdT6ZHQXFHNQd5NVrzcz06lQ6Qbgb1SOnZEdibV57o1foNzxosJ0h5Mttw8bTligIs976agCiHB
BUQGE1cb3nzWAe6ty9ttizIi0tII09i0HWJVl8XDz7qXK7R0lELL0GGbG8uyHOe5GOUBc57GaDUr
k+sqyQOCjoob+e3zopAKIupujFGodjVExaQlG4clvqhRFQ0GwXH+Lglwo1DrIdZIJ1n3XO3XuskF
nrlm22nzcEeP3n5dS88P9mXgvdAaMg4T+w/8rF9XXXrMH/zsHT5Q7NooWoLIvnvDrjdZdbvOfAJl
qDQROB5cXse+fvC3bLp7NMr4gBjDLMWqa75/HWQ+Gw==
`pragma protect end_protected
