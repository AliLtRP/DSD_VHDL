// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:47 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
tP+x0T/V3OZWH9a0/w6zseCn2PuoXiatQnT5Yp4B4pcvOhG4ENY8Yq4of9Vw2KZP
sgCPVFudnP1gsjONvfYJ2m5gPQ+JZdjLsAU6A7/sVl6Z6PnzNSkbg1HJ/V5ul4tU
I6lbcH9b5z03LhIapNlAodSAJEJcfHRgpmCVnsl1k6U=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 42992)
ryJDLhur+xfL/m5KU1PMA+32GZbqehwSeIirlXbX80EEYRlYXegIbwodHmFRXFq/
suB+NVDNIGBdfTvx0pFp4mwIBf2iev88+pP51+A98lZmlITVKWHC2M9ZVpL8uaD9
abmiNSm2Uu6eTy23regntNqNV35gEIXq+/PLF39/QztCb0OEN6wQ+8Goa0/mesPY
dNCdWujv5q1AVrA1myymENT4Ijk2wqh1ilsWyPnuE1p6aA/2IJfyZko5xsVqDB4C
QUykyRRwm5UqxNvnpJoXT9EEfkYHUTZAksUZcZBxrOLoElWbZ0E2VA2CCr+D0+pM
1H2Sa9W/pFpG5xIN8iKoDKFao7RWe5pEewhJURqnlFoWXZPC755BI/9qQtzDCiFm
v3I4pDoM+FyW6SYhcnTFEJrzAJsbid5mEFpn5hZyf70w0I765EwQfr/BTOlCjcYg
2Tn3Y3Ek1ueNtDPASXNE5xMjuPFqy+Ob1kxj5iB3utti+PmntFii0svQZ12L+kNT
88PGCnOIymguPVaWzqG8ujeQ/h9yS0w+hsDiG2+U5UEPA2LdU1fPrHepZInHj8Iw
UQN4CLUHoO3l5kcGUdbsifDBxZpk4nwyfOSjS0KMMd6oHuTGzKsTafnO7a1Wa5Nl
3nbMMveXvHLtoDDbdwx3qlvvpq48NmM8PbQ8gj/9rmW6keuEiIh8Bie24Xt3IQL3
DQByhk8OOX+HgRUAjSOkWmWms+zW4l6xnvm1hJVwiDYhWy5OE/aZDu/jVYcVTfNA
kbY8LxI6KWcd3z9Yhf12AIyEa7nheiz3FjBMYPEHNUGWpRaTDdtQDxIqiRYtlgdh
vzAg2FEzRCFohmdzniIAfvFDhdu/hLKdG6NqaEDcYnWfAAjskk69KK7Dvlb1FDNk
qJdTzOm9V1af5EJ7ViQiJoWrqGh7TzNXMdBkGhpK28dz9LpMqqysiORVA5rzv3E+
usC9oqy27X1fyvooSAPD4e1NdQgoeEYVXQBXboyK+gzGyC4ilO/lROXWJD8RcewR
6KN+Y0lnB6jMlTeWOOwDLc5O9OjPp3VJ4KINn2RVNNXDnfIlYHUa5ImeC2IF7Uiv
eJ4tSnAfbmAl5I2qgESUcLu/y+S93CKdjqruojsHnXCUNjK/wDEcoqi8MlX/eY7U
OOlJhGN0WmYH7KaxoEI1xNbJCaIPQazzJygopHE5owxlqK2dLKamOyU0Uz0SISsb
9wMh6ZF8a0GRSIWeTELtEbdBZ+I2ZnmHCm6OzlisYJR0K6sA3pgjsQV5mmUk7amA
1aGHPqwR2FFah+7HRfAdDwzv6/MTuvQ9HY2aSYx1lgPEPQ5XamwNCCJZTBgURjVM
4tNjHycnnD9wXopdb4d1sHar+om0GLhwaA5OISRlNx2kEDtdmYkAh6MJlU7KcxrS
LidJ840pKU7vhdhgC11lO9ZRIIa4z7rr2QO93HE4MxR02E7XPhS8qmi17emHbJya
AxWrkIDXmPnlXcNJcg3tR/gowLnHSomhKkG0ymk9D1NBChmIucvC8/4s1ssJ1pzz
AfCycVoLrTaQUGjcD0EvAH41514JwU6zVC6G/VRrrakhfUrDPGZrtSmXl1A85DiD
IYOx9z3+5KI/0E850Ap49kW+BJfABDwu4nT2sAwKM7EPdZp8Q3ZehuoMpDlhyHPF
VvGGDgVmubG5E7IZNZMU5URQUFKMPwVPVJ7bH+NHVqq8wWwE54n4oX0zWK4slEQZ
daH/l4Efd/0ICrkv53Z2YT7wanOJCZiU5Jn2q3vEWNTYBgl+CmNDThQkNFeiZL2m
Eznll9A0m+chAfSHDTP82grRDuxt+Ej9oksznTt2vP9w8F3as3SA357Ma8TB59NZ
f/PNznMKVmenNzAH+df1oY/p2YczmySFAqlojen013UbvUpSa/s+HQ9Y0qEedK3I
XOuppETvXBOJrNniIbBCnfmNl1jHzcNiVXPE8Ttfec/kY5lfKJ3UThlO8o+0FMuD
u1Dob9mFMsYKauhKdcvFW0fLH+zkfvIyZztDtE3Yg1G+wr6lg0RjLJur3lkV0tUt
eSmjk5NNKhx/iozW5cujwLVxk4eHYBW6xZNt9dL6EowBfdz7XxYbeSil7UxFQ3St
XGOaMkYhn/eIvxKvCoHWJ7FSQm6aXi2J0lWkFiE/If6o6FkVWszGm4u2dFM2itn6
hV41ew5CV9bmt0ei6B/1Tk8fGq1wgAhcG6ZC3S4LatUzEcjQruw5kPaeJEl+rauH
vgejZsg55U/ezIMsn4Q6cJvVzMS5gWIj/mRjMNVXIo3DB+0Mj1GRfr8OW4IFzm9C
5jFYr+JXVg5hq8bImFNweRgl4vmQoKsxzyq2G9ALgQBSmUj+8vNC/JY9lALZ/pc8
BPU+gTEzClBR9xrqSCmP8rHG+ieNfyL7qrKyfYXAZhO2rkXUjBvbi0nwJR1sJnfU
nEd0A1JLTUi3+HX6YV+Uj48zI9H0jH2gXcTxwEW11HnGfcePIv3JHZHt0J3424aG
F+aP0phQ0Gp/HK791E2m+mK7DC4kSAgA+0pxP8wxSTA0sFRrmi+w7JuCl8FzZt0Z
J8v1Y5obgG6G0u1z2Mv/BidKyzs1b2KJdlg8ZinA+YS6ynq90hVBUOQDkM502xWp
j+S+vPRs4iA+04tmqNlxC3ueNGKb3eF80jpX3HBZCyq7lK7oubHeMZ7R+9tFbBYh
LNosqIZjSHwcGp9YeJFsaaIw4OvRd8Cq+n0TCkdvDU5SU16uzNU+6Je9YB8vvgTV
HS9eqpqGFa0RYNTDQ+QMjFD3iugwV+AI1IVIeYXsO1VybDMf+Ma/RZ7eMh7g5Qcs
o4pHROtjNKyICFzKNvuOEVZvoL/nODrvt/c8UxJAYUxFjE+Q4G4iz+y+GsLi7v5/
UK1EfKbki7jN8Jg0Z0kKOwU+LYdzX5YKS+2Czl3aEtg1qPTtQJJARjTQJbh2ceZ4
NZIq4O/fxZaTfFNA6ZMxZrFoJo9Td3b5d0t12WJf7ZsLqWrcW7DBFrMXqy1V7+Cv
qumMsdqI9PVXum2AnzQuUJOewIY0Zw2Zlw9MFL843yYTxcuV3JolG0v87vYbjccv
ffAXTPAy7PfgSJBLczmIw7ave/HPOLw4VKTL+wniNFmloRz6rymMoVHhETM250lR
cDwm+FVrxEfAFyEGz7oVv9IEMp+C3E/FmDe2HJ56eeSsNv7NlLe/GHENNngPAoIf
ldOVIyr80eSeu5qxrx628aIvXEg7fI6vibHjJe7B/rcUdMoWXCg2HJQ3UcWor8FX
ybPNu23TipoxOvoWJjE1BzHGr0QBJ2XbgafrqyVUa62qch8XCwzXmlkjQH7gQZeu
9IANIUWVVW782oKl0kqxnRwEaMi4R4M+DCgMUjOG+sCv9d27tAEdkxnXZDVnbAfa
BP7m4PxHDIv575J6iMyR6RXmkV0Lj9vXbcmrCzzvT48VyDd2V1Ckvgmb8xzA0TS+
vQSehcW7KyrNUKzHG2txVdXLm7uKeDJ0aQU2PdyIKmwoqstwpaJmJuI3yDhe4f/h
vYEstqdp3YWFe7SQS0uTz0ckigVRVnZf5dyfrdSZXorANfdAEsnf8mc4naK7/hdc
A8/xsAwTr82xJF31O59Sy8zEmV/p98KYcq2yDG/Uj7lfAS7i6RhyoDtr6xXqwiuT
QeD988hLLlXt92f2f74dRFhcKGNgF1juuDPbhxdw3SqxK4Anu2tcIn2d+MzVYm0r
5+IlEkFUYHR207o67K7DpqeyljohOeGBYwqxPW3dM8g+GYWPESQxhi0gWqDL4lZd
5Hao36qb8SOdMvsU4jJZ6RC48azL68zeAN6hDg5iJ2ARyPa1BMwAJwGbrW0PYtBS
Jg2iyRtw6qHXsyhvcI572D1OL3bd6g19RtiS0qKG4iYYdttW4XLnieKCr570RgB0
+01p7W2NB6P36niONSNar9c1XD8jgMTwjADmkPTyXwUhPQXzICXW9MC9Cka019Bn
amnCagFaZF/Zyk29Q1SrHRQYazxm2+IBd/kRySGiJHFh8jQVc2op1Jh+7/KAKQla
9sRPSDDl3fSXW7+AomfOJ25LGO4aZvWrwoOk/lYhUZ07qqP0/K6bnYyWpkRLZXYF
DNSUIbc+knUayaZlRiiMWGfMnjhenMEGwbD3GpvGz25uXQ15JfeJRdQu15lSYb5O
NuK6yA4otV+0MSg6J/DEkijNXzY4IIjXtGVot9l7ZoNa5Tv+eiZ5CdrpQVstqseh
p5cArz7eiQAXEG8SCLHYOkbrDqglTrf81/CnI6iPZUPEbgAaC8QjfOVCaJOfIa3V
353eCwGUT0EhDUAlPh9dqtUbUrfuvPRJ1hZv614sNx5jLUmoFh5KObMmvYFfDYRv
Hllh/Xx+/qQp1eZ6Ch5kxkfHcWNINZCOaC/UPK1mEBJX02zMdRnT8LOmjTinjj6/
xi4KBsrU5GbohUOAmQ4dzCZ/xRI6ArAkNVLYlVcR5CDl0MjRZmdzyClqvEbKtWci
K13Miy5jfX6yM+GQl7EFtbMqjBViOFbuCEHYsgdzTCM/8IJzg01YgQdM6YwPzMnD
mm8/QMqUmbVMmVHWsSjTjIxrnsPtFzmfYcu54RF4NDPu9Wu38feqdVd23FhT7p4J
if8cN6bPB0YHIZCF3ODGilc7/dnDVsR5Qwt0g4/uuXohXvk8u5GIlFzdIksJDUO9
ypb9mypnH8MgfPm/LWZXf6zbrQNF8pwRNe2/qVB9bTKzUU1wpB24EJ0MuVo2R5OO
q4n6U8YpT1s69j8mGZOqqgGgErpTRO8xl9yp4S6DiMC8AqKeqKC0/5UWFQkgSMpL
ldJRDgj6quyb/x9uCyhn/FkIja0FiShyQYbGOImdyzSfn1TvHutdVOB0wVgnF/fd
KFP5iUZsWEEMFLamCOGf4P3nd5pyphGy0AHFH4YzY0R931K8hCsNSo+amdE8yzNs
RDMxlY48k8bdHSwsSgmdK+oJ8lqEZTG2FrBg/3uNuw0PaOI/zmpXprMFkSN7NKxT
k887L/KYFrHA17YKKIU9PDInr5vy79+It8xXyNmbHi/vMM6kZm2CfOwJXI0wH7dc
RcrMSmKrgeGybwH/RCPTeyr6/LpdWY650eLxxdwQ8WeMg7FhZUZUH4gQ7W4lGWQt
EUMZZe45YJbgH/gTCo1LblIP71WXrICVMqeZGFJCCu3UFj5yU9qwyaYoQgw3Y1Qn
LCO9rwnv8r1IeKm2eG0zPYat7w6jCvoHL7Iaovev6pIIDzkSmqNc6Oin9lJLPW3e
8vUTyFd/6CEH1Sx0zAss5r67gVQC+y2xBfWL8dusBri+hSQ2Ew5Mypf5t6/7c7Ad
TCZPRm6qTkAKyYf3OLvgaxzRyuo4XBJlM3MmRduHyW9R2Z52F4oRQtgG5RaUP/jr
DQqFkfCF1KdnFwv3fASab+z5JcHTdT3YdD+OGNDF0/NAcUF2GRARewJ9udH4KUTh
VAguduzVgE21BkDmE+oS2jrjjQNYQnkJDTYXKyCPz3Xg3YjZRhK6Y1tzN2BTDiVb
6Ra1Mc9qghzDwydbKlnDYAUVrrADhMV+7SWvpdPiI9bbC3AtQpg08nis859c0YLk
tHbNvMF4s6uZtSYx726hUqhWKiYsXquuyvNBFORVJUe5rrrfTfMIhPSlFb4/9Cnr
Vtz8OvBAyuw1qGt53fpk47FdGRVmznK+oLHo1j03V9Nn+vd0GTrWffFIaeBVYz3M
l65La0iqLEGNdxgRw0ZPm6j6y7LxNp5GJn5/RwMoqPGNkHYF0i3Glz5pGem7G5XZ
fZGqi4gw9WZ7sAWNXyTnLO4chnKXqRBQVmL2gPbIYIczgSIw1Ckcs6bU9Tc5PTqx
e2wIf3MoHlVQpuDTupZO8szqAfuA0fwd+njBLwRjBPxjoBK0dR8HJRdklhwg0kw6
WhkS9VEaFpwcTp3Bro9IIFyiLIUoiMQJ/Mb8NI9e/rfWSgrQrwqpcLRc4ASA7Y3j
yWYERpDCmK0GyYhPnBdVkAosZmqBEkRcL+iyUIgMpnAhCAYUS+IVMPFEsCCOjIbJ
sggacydvGph+UK/mGdxxXOrilm5ucBYHrdIhi9mQWrWLQl6+NtampIBlNJtpn9FW
tgVec+/rAUY/x00kcXXh+IpJ+SfO1L5yv7Yl04bGUs/c3EPENG89/0ppJacq/Tsm
a0whMlpLDqS8WFwIy4QYBAfxEUK1D+U8YTBk66S5NPowFpd5KKD32SsrZ877iQ+Y
bXXIuFjftPntvR70eF+KmPDmSZM7RdPvmXyOcDEY2zVup1VnnDCulrpAosUo0rMo
LN1hUiZxCY6/HnpneAH32VB75V95Irag4F8vl9O7fiCid1bpa5LyBygjVlSOfkcC
mOA5ud4W/IbeQOGh0SLif2dCfCrdaV3Of1gxrVigB2JqrTMRSaz7YWwmPa9FidLM
5ORDMs80BB+p0z9FaX3f5jcf+VuaCQ7ty5tfN07qEplB5JBn7EvtRZF5Hebx3iPF
h4BgmXSyk+Fl0E48amqjgVfNJPRhBBZ1w4APwmjpgpP4It0YiM59KO91L7Vzq9+t
PA/PumDNHy6SFLvKNKzB4BTmVscCnXaWK2tthIebfnkkrqupko1eXQQrhqMZurWQ
pitj1RDUQKb8/hbL6AQteIgMocAlCFIv5d2UuyUmwXDIttp60bJn+nnPYgig2zG1
8EbvyP9frMK9BKFR9yACi7Pcc4878sZ91YK2HtPNCo2edRRYB68nRyZsMVelxnLp
Q+6pYg5DtHL69FKakePWFBBL6Eg4RRP0rcRJRwAyWZ67lqVEWN75yjxlGgbmYzj9
wJHLo51EWLazGnZj0OFiPaPemslWTBYuwjIxj2QXJ7BS9QBatF3RbA+/z2/IfkQn
w/BSomdTHS7T30pVAvsbTEbj0D6CapKThDI46RRzT9cIjgZkA20D9+FOvq+jCZRh
mGFZc06CwEO829p0ztQQlW3Eji+WaBeuN2CjrL+G5PgaQjNvlxZobyohGDv/EdI9
ZrnfFE5BXUS5asbUDWo07GS204ZBeIT2yEnLaGwRIr8bDdqHYhLb0WPzIuISk5cp
eGNT35N29NiKDJmI/0o4EuBHQVz+AbExQbXIWOSKYpCgELclvt3hbiM/qKOi8RN8
vVIOap5aVi7klFMjcstLTEhphxqrOw/R+3t8WOFKk/mt4otNo9knituBQ+Dduzyc
Y30aAsu3YXexFlFLX4ANPvXSS/1L/z5ZgNgrJZNQrP5rF+pNzSsZO4sJYRzg9AVb
9AFThUihJMDwCJX0iemOBX5jfip88vSHzURKxgBFTXzlyXwRI5S+5AUx2Fc2utyA
5s+lQIIg7oo7mqRkLoJRJMvgjrCte8R/WriETvflfP14zZsMirors7Ifz+939Tlo
KV5iG59r/8nwN2nYGbeNfpnZkGkpvMTsYujHPWRWUEZsvzhdHQQ5faO+uwMxJjYe
kdmc/pXjRZLbfTO6VxYms8yUdgulLL1W+NaYhL6LSRXRYR3JCajTL42GoRUtSU8z
+ynHXB88ooryO+r9cEsxLNSMJsFJy9SD50Jd3B1YkE4kKsuTYKHVWH8ap63a7d4k
Y/19OVp/pU2uDYozGP9ESnUuNDvPjEyWPzRBy3weasg3oeO0W7ELNgOXyTDkfH7N
YusWe/ANYLiHweb9jOaE+VZciJ/zGr5HjjHwjsNScAP4lCxuGpKEp3SapkP2VUYl
JxtSkvWDrsmY8Ssggsuy5Op1bZWVF8eVaI7ay9DvzqKHtitKdcQVgqLvM3lMDPCe
OnjpFSbtGNrqIqYlJkY+spUtZuemUnLeK5LcJUiTwpOt1l+36nAeAHsdBD7lkAwt
LujA5qfBd3VuJP+j7TApi2hJqcMrPeJQnOLkvR2n3/Vq55fZuSLv/v4yOlsCk6oA
Drkp3yHXhptG0qIqsV61sSSK/6w2vsnW3rw2zviDt3it2z/kFaa95IDCjewzy+aV
upRB9SL+Bp9AgUWjpD/DEr21IuFWLpLvd2xZldSPGnvLQtQhe4izyNl8BBmZhsj4
Z53MYXV5mbeG1PUV74r/B3OJ8KYXGco/Haj/DnaD8gyWnalpMRY/zANKxOTyF0qV
8IJwcZ+N+cpssFFeL+yepL4DoOZRzN3mydxxiMN7ImikG6sZiG2039LhLdiVJwfm
hB8QvkZa2veTiiHvHLUazrqXgMEfa+xw4wZAxxrr4t1PZUi585Al6GHwHz4BN/7U
lqB1o6WpJC1XwGh8Y6luZJW1doQfuXY1KFCwIuddnZCqZJsv5sA+5ITjKIIoO8si
/efUTiNAtlFWCyHg2hFkAwKmp2nSTb6CuNzJPeSvZ0OXazv0bQvEIfb1VoShNk2x
8PfB5Nsm3vKs1E3z3wJmNauE5szQ+5rRftBSgMLGUvGNxrR7rtErunqqxEJaCaIi
ZfuIABzjs85E8ApUgfBIqG+gTcoF0LuwuQBpnhH+NTfYimATe/a7l4crvckgGh6S
sFiwNfaJRfZ2exgctl45T7yP2m/loLMEBsnFSlAMGS0dbmuWSxiRFa4tN4w0a0Ob
DeU/fExFohP/ZOB8tb0C+P5KF4vsoiLEw4UNoKItXWT5flQJujIP02R0hoYq2rfk
0wjXeipJSiyzpplscFiAX7ujXi/deppePd2T6k8JC8CiwjBwF1JiUeLg6HKLiivd
xaOh4t38NQ4ksnG6lXaD5iThSKFm4Ggb8OC8/V+bGDLc11ch/NoeiVAJg4GAiLPz
cs1JqZneRKMvxf+q/nmlAO/TnTqdaedwNr+adwR4JpHjoAw+SItOabavypM3vv5b
ZFY6zvlP5NGJCAXsiX8FQKngoPSgEebvZ2Ia4EdOh0WhDb3SooIhXuxohrfjw07+
XPD8soEfZJ1qKwM+2taIyt8R9jljbRzKVeTiSPRURC1iCk8hvzpJzTmAHY4u8b5v
j3ttYpwl4Mr7Oz8NlSQwv2qnJFhwvZcBBsmRO0aeJLN6izh2s8Pp3G1YWuGzoPD0
2GRoGHljXaXbSIavB7CfXKgnJsxVhs921L2xbZw2IcDtNth4raVFyVkirmbqstJS
p6RO9lDH3Wnv86ybNYg2v48yiwSWUqNd1002iVVQwHEnl7FHrsUZADdaqUO7RFfT
NigWl/PxNzS9B+v4pq3+TzzIRcXdy7yAiiEe3X+SoKFPBBgMrkF+lsXmDd2kqUNa
dXaY1tUIXSGlZA32P+1wz3N11v66Hd+HG97C7z2iZ8eXSrhXLfn0nXnhIZ7MS/16
AKd7TYP9fy4pG1P01yclJ0A5jv1btE8iyB1B2wzJiXiMwtCwGJABJxo7CbW9iX+L
V51HNCJ/w3zVkCwQedp8+ozmWOJgjjWgXp2FaLqnyVeZHvaSg5xXn8wC3+1SOLDD
Dsr5F2UNQACjBMfgIQFsCxTP5bY/oEZp59+B97fCr+9sFnEjegLbCp5EQ3AszZi7
YOmer/kRJzevRdBsOWZwdIjtITfUik9fm6dXEpdPEFZKZfIUl5WC07r1tpm/jkUe
eiqu+hSXh4Fe9Y5vAJfxGPGnw8ENP+v/r32lDE6QnkV7m076sg3Di0hB0Ee06SXw
BZcDoI6R1shfQhYUXy7gSJxsT+vjHCZu0eaXm2RQQMiL9JSFtC6MOaqFrh6xZBny
c4ZteDe8qhGlAHgZanYNvYRdKSMrP/wXk2HHamtQXxOh1CeEEMVCblMzFsWDDtwt
wewMADHBczxAv4lG7Y5/k20OIwjx6LozVUikMnPGXjJ7XO122HYdndjQWUq8b6Du
KHf8mnAaRddhj3kVMH8JTcX4wAFMBzs7usdushiFN8tt+DLSHIX9rijFoOcrllLX
xbpOj5yjnJ0cB1lnTs6/ouV4kvPNBQT5nNPVfjz0FNwVcPEPSktZGg0GSaYDEHQL
qsx98BKRtFJNK8ZH0Q7I9cAMFQuhqlpRUeBOdHPu+/98RVGOuyFnEvn1MmQYkPfj
bCN7HAzGzgCrgaoe4P1qBixKlVfBvD2VkslIxaaajGLw+BmV42dcExyVMnp6UekT
w+WctIndd3dCkPTqoblc34go41Ryr7Pv7NRIuKRrmNYsLzUzH5GGCTnyUWGyDJZO
jpUVAYA7daNrFxz4/J10FVsis1kXCEcXV+9JzRd8TcdIDY8tPaUGKSCOpMKdGG/L
765jyQmXUduQR8mhJ46OVQaJC6JM7Hknx48gBh6BC/fAnjRTDGgLLtS8wzAAE/Tz
tKiaeru5NkHwtw+bo1pjW0EoYexFq0wZzLtsqnC72Ocqaj8cpAarS1IeAh//LufM
M446DgEF3YhRQwaOOMJJyfNMPNwfT//Wv0d/Y2I1axGJI/q3xzwn6Xh0gMrXg7Qb
EnPNsKmb9VRiRyE4EuhMmDmFguyitBHdd/p/jjuvBSefDSWFHlQ0ro/AfJaFNI2y
CbRKNtFhTeGHBTKdCShoQjkRvkE7L+CdfEB2YL7Yta5Cnlj26UDnRs6fjrzTpdd0
yd8LtxzOJQdMByuo0LwtNGFh6gH6Tc1dDwvbPkb7HkD7WzK2PFejuGB3s9L3v69A
U1w82WZcx5LCtJk98QUJ+IrwFllogK8aIufJwI4NWVgcZOHOYpgihMdRcexYqpKa
/zvphNhdz2CZRJwknlvKI96lVkYPsi6AkhUOxy935A/zSqxr/TRas2zZr6KlZsRg
fs03D5KPS7F06SP3MsYgxXMxUUatzJWctNLSWHYohdTShuFbGY/3VgN6y03FG3Ox
uQJ2n23uemBul4rVNWFzpAfh8/RZ251PxrZbBVgAgt1OQtgnfzlwNI6KIQRtiHHH
FUuMfXYrpYz9SJnb3qeC2dVVaCA8HtiqL7KBGbk+l+YvmRj67jEbNajW10snh/mR
/dZ5p6RJTSRcSAh6yuLOl85paTjaBRVg9j2gWyqIJxHo1a/ZWlaw+HMESb3JMR5T
UpsyeMJUkIgSaUn3JrPT7lr/QMYiodKlvFC2bZgMeTKw3V/KXPFsTFFALDwcO8uD
o3mvaXSdlsEfiH1+2a+zWI8qJVeR8/KUkAZfX4vG/3C29Sc5reZvaLSaR7vu4yzP
5z+KgtB2YS4lrihQch1aepMo9gZPurQ+hQO7Hjs6vWf3wC0usKKtGUzdH5Bw5ogY
7V88HQOGY2MdeDY6h5JL0xr68beL4uXK0NU1Ex2oSftpvE6BQA5wK7kmOj1Z32en
g0OdzqPbpSyjHONg5esackseDdUJazqffsjNxKNJjZ/4rnKAuDrJb6iNI08cltWW
aRHlu9P8L6agIT3819klO1AOlzgYkdHe1Qga8chmsLTpsi3HdQFxfV0tQUWFn/FS
5uzXUdhqVrlQODk15aRQU9v8c1fN/ZrazHoUvxgLal7Hpuq4irwaVukV3fGZFNMq
LL/zr2M8D/MLJIE9+AfXk7+zSB/wNQfFKf10B2M3gyjnI2Kx/PyUkQSmdEoD7+Hq
j+MyI5xDUJs0+ITUQMnDgj47saoUDuEW2DL1Ow6wGOF5MAMdyv8OEXkFdc4QLqAa
DCvgUPN4QIzEF2ssm0W/vuyqVzTPLlzRaXv7lQO6j73ONlKgSrtbU4awMMeMTG7e
Q1ncNhfdjhOlmDfZOTJIrtuJQ/mN0GQhhYTrCxdDYPs5BJ7JQAp+UKuNrH4kjz+K
TcJG0ksv/RI0cQIzgDRkGbq/jsdSbgi0SVtFmDhZrGZh98G8Xl2uyD34TfF0TZuk
GyA2rL9pTHtrRsegSSrQ6tfnHkyF6D78PTj4jIb2QudCNfRSZfNa3xMfhpOQsRw3
d+WLOHphg2n3vEVxmKnvTGCoR1JPQoKMU4FSLXZTZS4fIDkCwfoBoCPhH9+N2OyH
BJ+u9dOy7wPX04yRGbKGKjY9NCzdoOtvNiJb0fLiw3nNLGjDrdCPpNZXiQyr12BD
Bu1IBtuRVfQPReGPg7NjDYnVFmH97TAIGbXQW9a3pplP39BYLZE2fLaVmwa5+xJD
OjFa/n9rjtaLa4uLBPYL74fmVcyeeVzxW8CnRc00WF8yAL70KRocBlbMkqwp9bfQ
hjqu+1HO6mnO8TuedzqmrrbIVt1pko8VpdJa81CEg5TPJ8MCrzjoajqA7klDQ4J3
N4UQpR16QO5vcxz2UsrShcii6HiHiXsRuMc/dIpmEyrboKYaCBfH8lpcCVbAFot7
X4SqiABmKqx9iIlAf5lasH+TB5xhviGbZ/C7s+wRHrmUD2ulb1SLvZug0BRQ6S7p
E49Ejh74DuYfqvA4saB60uI9dtzXLlgCSN6gSGiRetp33n58qlgKzQkv0+TAUDd+
cprjOf2evYjOEHHtybjpPVziCQJekRlenHBA1fEp3iG/GSFnxWqXIqv7TLCOQ79k
O2V1sOdoFtI+H5BIaJypO3DUfKjOpsVop4S8LLR4G/xobg2QF80JLgY+W8c6D4ra
HnQqAAabUhXdtfG3Z0ufBSSvQHKYFFtfoPYve+CZExlDOLQayweYNO40xdgK9pL5
rRktvzKp+aWWBR6U0iH3FDwrU34ekNPy+hSbK4aTJDvsreDVxsm9of4oziA0dkH0
oO9FPR6odtQocVwYnmT9RJBprN0vSJHYn49ZWUEwJLBuyRRxy3hu23v7Le9lapz/
vBw0zrhwcSDQf6AsTilmZaFjXI7LuUxx8MQs62tSxQVd0g7NBgeMX4HGbJyHw3+U
cYXps4ap4SgCpCODg5uMIEy0eFiaov8KUI22YXYy+LzYIgrc9ZfDW3jhAKx3yfSv
NWabv7L1ZRz+gvG1/bnSmUhiL0+V3UkRxzKN2AzlfHOD/ejl0FgCUkNFUegil7Az
l2OZ44gMx3hdl7zYUyts8h/jUVmztOhFtZ7box1tvr9HPq2kBCP7rGFl7nByP6qN
5GvgjweDi7yljDkpVEVU/KSSlTfeAa72VMR2wT3qMPHgiewQrye9VXWtAED9H81N
3Qb3uzosME64y0T/7IRcvR7tuqYSdWyWNn4X4W4XbLfgXDKMVzNcdHVqeYfJKIUC
oniwTcaVF8i7Ui/z6ku+r82C3DJDA6SiNa+kcIvSK8Bwz8TP7C2CB0H+Gq+/HN5t
uIElG2fiQpwZwJuUSsc6g1xERQdWzqKOI1f27mArBGEi9t5SrtBVGoOYjpCrvW8n
It05G4uzeJHRu32EWNtvDTrhMiBhPssp5QPsx+0jHAVwUkA5k8Ec3xe+4I7ZHlt0
+FnGg8wJN4WxffE89x9Xg+nGOXsw1NwAMiGmGd57V9Yx8DhOdMyYAZgDNfYwCFI/
HU5xHC0RlkjEkMlRgYirXKLfaSWsd1ErEPXg/W5JiUZOuiVV7vJ85bjbF1VUTy54
yHFQwwRPmX5VmFBPfNMePX5cR92GWkttMfvIzG5ySsSK7VQ0NDwLDssIFCq0A09G
EuWTPEMYaGmRqwAyop1RMdbRR0ObajBRbPFpYQkYlKU+sgfRgFsiwPSri6zE96mr
eaaOuvkFuh7ZuAUsfTTKErm8WNKgOsfGUERwO1ks8fa/lQ+I8XAdSNMZbwFRhPq1
QvQuuvNwg8KzkTb1VbDQ5kAZp1K2l/HsLl6J2JtLtNfoHAH8opLiwWBe+tCxWeaJ
H4uGl8wGR0TdSI/Z8RI+OYXJ95yN0C+FYRSEYdUlsscddMuOP0UXFzM2oH+Kh9np
sWNXvn/6WOQuPMiRk57A4MVYToyxdhC57m+SlFuvT9bWP8aMQTHmAaeCDg/G6dRt
clhLV0yF8gR7AJJIq/M5uw5O24T9YSCgMuobxiK0+r4RRM/DdbHF7AL/Mxfbhdbd
iEougM00xUXoYLKDL5gXmxLYOUCvBz6tFiaLEFk3vWifvN6x0fgxrQIhQt9SfjBf
g0rEzCDZf3qHN7CcIJENsCae2MqSLTHnM2pQGdjAi4rkRAcRk6H108ukgDdl5rOt
IpLYzUlehuy9fsMuliUQ/kPp9htBLOYpvQBD7jakenBkGErsOj3TXG4h3Ww29d+v
Dk3wIG7Q12EYklMgvhrwFGRnFv33Kh+v54Z2kf3qvLJFNqjOJYx+hluIQP77iQkE
IY4tZECZAS6l9ml7dsERvQ5GUgljV9iYUYnb2nNCRPFP5ubV1Sj0mIKbc6IKa0mX
gFZOFQlhZgIH+raFNakKbAXk+XNiIAPo6g+NDJ6bCjLvYr5yuYuzECTK848eOPKm
aqOuMVqFS4VeAQLUZZZrAjRflng3L/6Hn+/Dmp+Z+nmgoJC4Mr79yLVqitBIwit+
J6PLZxxXRMVk1yMjZigFk64XsDHHDVtqwSyybQBrQykaKCdGZIpEP47w5fV8yjoY
iyr8diXd/KWETfFg5zWYv9IVYR5FH3a4Q1nCGKR4Tu0PxEgigURt4x2Wlo0KhjPe
P3QSmHVx5COpqmPJWPIusRZajU9mKYI8JAKcte2E0jIF3Wzu+RrErlPwawAqJtVc
UmV9GmOY+qX7/1aDPyA5TnKf/+sd+5ZHsxPPQLtGXUTasbUcOo3+thW/mQKqngRB
aRU31u7zErOHQEE75LujblGDYZXJAagRxLRQeaYCZXvvaYpRGM4cEr7IBLcgIe1A
xhtE9RV+gxQz9VrgdnrOHV7BpF32YNbtdiAJBL3bEw2fwxT+B++5U08pFh/dMqfr
wbA5q1S3DTmdDuZL+uesE8lql1l2OtDR+2MMXE8QwcomwOH2PbuBGJmvVugjzFtR
QTDb6JQstX1iInPV7hMW02RThg4QAsD8RnJc48OvfK5ifezztUKV+Ooe9kUX4GU1
vYhyVGikmVUAxp0bAFvfb4R9xv6Kx/fpvx8i0SVaXzyH2/LiTrL+WfNuBakM39ua
Z9Hu4stxxY0lg6fm9Q0aqlVpx3fZHfw3xhLaRJ7qn6FJf6vDNMPNszY4eu4rItEv
GWzNtzoMyEnuENYB59gTywolkDxPHoDxBKvGluxVAQDfp9u/3eEYFoNfonol83p5
4YgxqkERI+ThWFzTQ5ieKo4T4fEc4QYF6FmCA58BME8TwKIRA5oDHrYezxhGgN2C
Z036Ns62Krx4mLOSKC69/99SDbKDoGpQOm1SS8ER0IfrXFQ6MyNIVk8BB7uv88Zf
pHDPC/OvIshDvsKw+sv2PJZrIcWKsDG7d1TaC5M70pirCETsNVlZ24i5VpD/pLSo
EVFMF6FU+C8rX6exRNcj4lOzoOYw8pk6XDMOdp8E5h5VfU6QBW2F/ubMApczhQ9n
+9mL34D3u8Mxa52q8RWoUxcBf9zLRIaZ4sxUN15fMO+x+pT9BmEuRxxh7HaUJFAG
LuCFC8QQ8ROQBM2MboYJ0RuDUsse8KevUUMEHxOcoc5yFHefnX3EfVLq27Rd95bd
NWOnRoMFAWTqRKY3Np7MtUzqGxOgJWoqR3dziZ2Y8Dx2PiDBUCcsRQQ0NUgbCA/J
uzJ+FQIoD9JQWuCeFDUZgaR0WwogSxue5hb3mWM8QirdgzGaaXjD62ToJmgSiU+5
p7nbPSdFS7PASWgKNQXOi4q4dtdK3kMQHGK24nR9iX6g/Z+K4qMDQN1+j0uZAjq6
hR8Wm/VRsW+/vUCNXH8LEeepe8ZB/aWybek9+wr8PDCF8GCSMVvZYuxPNtUt+c/8
AWIcjRUca3BU3zKnKI+atnMs8/dqKfW4/jJaYRlW7y5xrtefPvmGBAZCrPeTPF6u
fVPSpfz37iBDMvS+kAwqAF4a6Yp9vwa6XN+BZFbrY/Jv49pc+3jKAUC9zwtG9Ak/
9MgHMkPnkjdgYsrsEXVwp3aKXaaVY3bC4xMgfEPVysykgxA5ET0dJxytCvG3CBL2
wXfXRqIGsdSpWUhYo7AmUeop/vmtV//5Mq+dW534VPQC1QQmOg6ygnQvs5DzMzWP
//dc8wJC1eXWuoiEYVvpqvSQE4h2zOD72sQxYpr5bRPWTJKUPxcOySTZYQ4Gj3/t
6fHMv6yXvCeN6hAPFP5wp3gVeC4vWcf3DRJwvOvdYixdzRjjMKQafmqLU34uWhaV
/gcOL9cxKU7f8GmRdGlXnZQrtStGC0oE6pdCl5bRwWqf7vUBjt+YDwDKHw56pr6Z
N11MtCmxzM238UqLFF4vEK2FG9Wb6xutBB9V74Wg19Y4hMHVRpYSlQXoPsG/oOS3
SthgySmU/J1cWDSltC+1sTuS21tYwoghUQ5JYs1xgQGKja3C1R/C0PBMcCIBclB0
2OOhYSpDO/77Q3KrcIw0nwFdczSiJR3rkvKgocRPpohNzd90F195zsIo45ykaQsY
gOg5C8qdwXqNXHm11cF7Qrk0CuA2xPgYMiKpqpGeXeO+zGbQiW4AZ+GY0EH+znj5
RRfjkNLFVBNCpgnSoZdmxWIIcygcI7oJGekj8ccyPMiHUlMkQqohLVgpJuWpzflz
x+QypX0osHyhZqiAy0s5NFReTCT/m2SV65n+6+G8UkSxEY8Sjnn/r4da9DTO7nc6
3yN1mBSQxk6eL0GSrE0ymbaeaYJAZCDM2atrRF9q/7efObBUKakyyb5GQy3F5FdJ
0g9plmEm7g2Kzujw58ijnPmVJ3nuzCMwqpHKITRQ/q1SE9FSb133ZpOOMHrDJo8D
bZHQrJUZ/EjKL6HwZguq1JnZlU+v1WWM5X18D8i2H27KMrXbKAWDlIM78mBKxN4x
elc1PacyQcKkoq2zWb4+NYAzQJj4AOVpaZYPMkIUNkK6W4Ft2EyIX17/oTQ4G2GI
UAGovuvnBmVn5wdX2PsQn4EY39KC40cjGw6AkLlMJVz9SlO8Y98PFZoIKcHh3TCp
3FQCAHKZdT7v7eOFV9K6BvztvgwMPl8fmdMOecYmIrkAFkRKjqJhWQQG+9jPrN15
BOxCYbxwwCMCGsQVk6v6MhSYKg9qQa0zdeJXiSPXue7J7BXBrjQ1JijH5efII0v3
2tDxgL3/iT2Oad+MDdD9TGFpLQCYC4NE5Ht4m5LTsKZ0ZqwSok2n+3vpgvi6MswQ
SEwPd61csAkyGk9yLDmf3c819vM275pGIy0AqZRyHbxaBOdLtaOzaI+kjx5I9REd
CGVaW4qFIlrhgh9XHtXUzpi2z6qgljtyKzgT87Krigrmux2/W3F6VAxAcREVl1xN
kZAAapiROCYcZfCjw7TFriCaUF6QkfLGYi1h4i31wK4JnYGDg7tqfOk+5twX3QiZ
XcqZh6NYCJh4ul+FNO0QKf+E6qsP+0A7fVKBxfIs3/d16HhDy/TJEHSnmuDutIeh
ZbWf0oPpjEB0YmaM7R+VGW5IC4/jDZ+3t0t/FYUBF2wn/cBoH3bUz7ZfvApycCux
CvlZhSYrli76oL7/ur/6D5q/i++D1jHdw3l7gmju/4H4XnEPz8kHvOwpbAVMgsUu
HUeulZy8/EEaxBX6bYTfx9ARj2oU5OXtdqrsMm5Se3+slvakgi3cfQhW2+hn6SnY
TWr/u4fBkwBoidf0LE4j9bN2EsibopbbXFpawAkX41w+XjrZZkMyvscCwHJkjLvr
K2QN1rAyTHDB4ARPeM7L1oIsK7Br7JlT17eUArlPu4kXKwFCrVmiJ+/AOHVTnVwO
Qdx3nlQcnuUP8e/dWNysubXrDMqzYZCDoC1sHpjHIzNhbdXjeKHg3w8n2wnfz9Ak
URYphHDR5OpIZLzZEw/HdA3zjV1ppY2koYN3dE+PSaY+xs63dV/EOPBROpAqqb4h
V8odBsCyklsN6nqy4t0U4ZcimOt5aRJqhl/Dvq6k1OI2XAInFaCEVn+FVG7DsHw1
7H8O9+lIlJI1icEAPI6uHfqWemrGZgnWuyBxl+OqT39i/RpDIOTb862ASHdzAtMC
UqljdbeILcw/h58v41LGU6zcicoDcXr96YvCuZXgnMIrZ+KtncnloBeDRTjX0UbT
UEUKmQgpjr63USxuFVRb16x75Su5pJnf6Sqxad9cXW+b0+AQmTP2AvVYSp/uURj1
mMY86BaIcbzH3wmJ3nUMJ4IiaNEed4UtoKuLHD231A0wynQByqqEg2oxK7OWkJ1i
BXAYAqqB9TILLq35OUHt/nmKlQwpO1osOFC3qmMoKjYXWiUFfglEMbKTjptn1HLL
SGHU7xCSlBRMgs1nUcu49xI7SrVvmo0vz5QhUifBnlV+tfvQfN0p548xlB1VhGpt
pSJ/19ATacBGH1yFRlRnuodEjcFwi0jFH7wEq6cS0vQ+vSKXkyNA2RDV75MLLXvJ
t0dPQoJkk0nAEL5mk7lc8ZdVBtAeyINerAeMPBxsfCAuSD0XIasmW3EjSHtFWzPg
32Jy2sk5mxz70uwARocnVOfSJjymPCQnHdOzig+yGsjPpHhxZzR02mjzZhablNeg
qTyXUjn1RXME7aYpDOg2JnXOrqO4lOWCVsBJmUYtR53Qr8x+YtNLJWE5RNN2mbqY
9/cf0LTiauLIMKy+NDuzaUqVbzNxyrSrnFHX27U6gePROYHFojoMzfwHXDbKHY0J
PTN+tF9qhSGG0qvbI6E0TMfetLBTbQaWOci1sOr1877JB+I6zJJSSE9cQ1Yz1u7O
l4C61wOcgfYcwYQmsNxeSGr44TXQA1m8wQ/742zkGCvsnQ3RKo51Mwq32cyluDXl
llEnz6HRccX1mK4Hh7WxftA7yJhoezJaqZ0DtlGix+3YIBHAlOgj+NQf2l8otPGS
o0UgEEYo8g/aYKvZpEPPqFyhZjVpQ04u76/tFsiJRwYyA34GTeP5L396oGLkmt7F
/3HARW6eCnvCeiYxNV1Jl+cnHG3Om6iaQMtgKRzhwvsM7Q2+cm4DDUbh3ysGZDyU
yt/+cVUEAu8OpRbJs+aAxA4wp1kuh2o8SdPF2zktusrLclj7caZmPtqlenY2/O1B
/qPMjlAFaftK1v1aF3ZAyHXJheG1/p68Wkc53t37VeGdWLx0PovDGTWRVg6EsQoy
Z5hYLCy/wr+W0SxkPGFc40DIKFHtDme4gnTNtxyUInw7CGNOGa9svJE1KCljHuf5
X30lnE8SmsAy07GbqQIWUKc1fKrvApgus1gVLIIQ2r8xCPEmbKC9ltZx0EaAccl2
X5ooc3NUK0o75nsa2bFvjapFIrFGp+JsAPreTZ+xw7/QaveTR7GE0Gz5S3tD13sn
xbvGPALN0D+lAfoD5PFFhCjiFCYjTrPqBUu+mvEGbk//et6p4Z+sQi6LU+lkCNBW
lrrp8c6Oz8/hj1K3yLKCWgDl0EwmwgolfHvLcOyXnsEPeiwrjXiSi7oyoHkM1FCJ
s/RS9/csZXgEiRt/0pLoZPN7FqB+5eSguc60hG5QGPR3Ts14FsuI6tJKGGcmkFYx
DzOiYvlSPrdtL3pWfa6y22TZf3JLRAWkP9EEi3QxUKxvdN9crj4p3dtOJdwwB+Y/
ErIKWZAtPxNI6XyL1WqAj8yeUttD9vjjcQUwd1j2uH4s1fbWowqQf16OoEy9WWNM
2FB6baOx/HgI8YjHDasNozOdgW39VsfJLlHIeQT1coYX1IMdvHST+7wEez+fHtJh
mmJmkE8AQqLFt8gGCZij5t3taj6MRvrXZT35yasz8Tbvih32ExxHemJkbqB2sVjb
MrZTX94b3BOl2PrdBBZFafg7tW0ua/4sWfyd87/DRxDc6CSlR2gxjKZKahckX5l3
k0Jc0M0xizxmdKuCNsYBCtLapD6VF8A3jxzXyyZumqhG7Z3MTvuC7L8CDaGdWFNY
JdUXpBd0uqZdJN0vc1+S3cGIQh5GIwhKtb84ERH5OP9GxvhstzPzodhdm8GFR4pc
28xu66ocdv87mkL0/iymBzBYJct8yMPuqXFtRJjcOOVHB1wSM6XMnfCvXTXyi9Ea
1C/Iti3KxP9amJGWY7+zzK2+45EEwTtJFKZI7//WpU7FWZWH6Ywhgu2lKZniIGqm
EUpPz2/xm1NLt0bTxslK1Hl93OaRtKbk6UrTD/HROzbvQhoiNeivZqvs38qQWQ5Z
GNXE6Qw7W9/pYNJgPB6fYBdGED3jMnKn/Zgov0OpltohlYnm9PZGs3IBVOprXSbQ
0pC2dc8q7ehE83gYzbCqEsjIJ+P+QV/GpP57Rw9tH6vfp8tw2QkGc9A6Nk0CE2GX
hwGTdvH0C+mn2WkSXq7R2LvRcLFTeVLUvlXfS/9TjZG91dUp/Fxtmx99sdTo0W25
D6aCuSENeGLoPaG6WJ9nnwpB/0S1cn4NV8oT5fa1oV6srZQJT4JO53gWbMBuVGaw
3o63odM6yZzv/bP01v10ZarRQCHPbVSc6Wp3ZTYYJrAZz/dVEgNOJdvWsHuOMzqn
fHUL8br8sJVtpF09tyasIcnhfblNloWBFlCT9ge0JEfr1vFLZvL5cERF16L0Q4/x
fm1jLpiPk1YmlD4HsEz52Dk1M8C1j9fT+yiOGbcelQM29ylG549IdRcIUTxFLesa
gxDb2nRDu4kGpoedzEPXpgNKddT/g5q42EfYMUjZqf5kt2qkXQlFDQTnfmLWCyWA
/aQdHonUngw2PNbyzc0gqgucMlZ1ciBQieHwSKCuld/zM7dAQ3V99KiIAuHevwmf
VNTkywSLpniZ+OfipC+lmmlS2KEgKWR3w2mA74GpsZ1qRwEKErUw7dQDIzNWIqVZ
1t3NNyjhCt5PrWb5FwWrzeEv1nLBfPPgLtq2FGluU6otdBardDBpqRrc9Kd+ADUN
hCQhk7bZU5LtmC0bfL786tynNQDaQ4j/Xi9bsqnuS6X2mwzw5lxG8xEfiqF4w5Jq
7TF0LbCCbaUxCoOlV8FkzZoBpOliehOGjHMfqLhTX/BaqkeF4q3FMEysp6jrUu2Q
LrkN6PgZPV7UDEn4xQoa44H1ygzxk8oBGEHlydpgL4xOxQxzjZedtA/CDdLo0F71
+lP2PahzuecRLHEFNFBqgHznZUqNbwtDbGUIR2OPq/JVSZLVo8PC3rDzDDuCJwq5
Xsb/nUQA4mScHG2Q6FEIUHT/NAwPfunXMmokm4USw7EC1t/uPm7f3plxtlvDB5jZ
FAbgCs9JXUtgSQLenbT0G9tCXzAOJPhElF9ZD1F3aExJn0YyXdUKOJKzF/PPuSrp
AX/Uyicm6py3zZyoM2ReRwRYHn/2k+of1ff457K7jIfsJopC1CCK4jFMQ/ClmZO4
Am7hJAtfTChGnGiJkSPLhHkjsMtV/jcQx+R7rAML0hBV94adcEN8KVy2bSZTo9b8
xIXXvCa1dzoYkSSgRdHcMoTCpCL/3si1KwCVnGefGNTPlKUr7h0lrELC4oCiY7Qe
+lNjCAeSa6wmszBqyyF+j+TsOYyG/glqMQ2EqWMepXojPQifeakgAQeJ1cFZhxPW
rfj+K9g8pcblwhXdANDogKOT1kNRBZOLZIcOoK7JN9CZCb5ZGPQGR0PRw9BACAfy
LIM/hWTUUjVzAYP00CzdriiPR8rrpDFWqNXXsUOtiWMKlIoJQwxuHW7u9Ia9WD8H
hRScRDd27O+DogmJJ2zu0feRLxXFizysDPHVStEr2EnltZQQnyi4vWaA3xn/E4KH
1zJawJABmTO6UkSywb1mKHiQDi9iymJ8CyOrHKqdwzJVPIYwEnnRuAHJcNHWCbR6
gxCRofZ/Zl5ySgNzxLpAO57eJcBQEZgf0pY85PIjM+3eYu/DXSJYydi9hKeR2Y6V
CxU6P7BcEQzqy2Rmmtrdlo3Yst9o0OZO+s60aQ8dl4EVg7MMUqBjGlaP4EIdpnRE
5VKMgZqkUZb+KYp4cMfbhYcwAuoKWp0ZUy/WgtY0q9VTUF2bp0h/v/LNTpDjueOi
q9o25mQm0nQcA5fgCZzufGDfyFBPabZ2PMDKQsjpfEmqvo7sSX4Y1effiTVLtMSe
uFhHBlNQiuA7a1CtpDSahrstpSzRuCgOSkQwYRfrcIxx4CuMdPlH1sr6Wq9qoeSG
VGLQxtq0ObV9GIBmNC2rF4Umo3Gau4adVeSz6Qu4oUCmrul28Q0pmC+ZAu0d7aAH
B5Ch0TQIl3qIQV0JBH7ya5dngx7zDtNzLUjHbS+cliuMQO1R+JBpVEsGbA02jXAd
0egmW8pUW0zGukkBhkvhyBfnMby22ulhOnSdEs5XKmaNjHubNifFg2zRCS4m7F48
RQWaTr62tCtYtB89YnhckyS+KEafhN5/iYUFfkHl4q5PmzlkEJP/HntsqIzuBf4n
57frxiPTGeU3lWxSL4GQTMhOasJB8jhMhYCqLhGRhTncAaGJ4pAQce4qpsO/8eiV
xVN/hkKtenvK06OMVpncnegKszvCaC5lR7s7DAFxRGV9iY6RaiBJvMvoePbQFRGe
ImuB6NBUBnW3WE7KLp1EgtGQnwVbaIYSgMSnOhwfdMAEjCe5mYEvnlZvM6fsW+nT
0zCOC3qW8908md5zvAh8BpwDQxv630SQJARM5jCReKDiXR1UfbASOpzD7aZ7R2Gs
lCjccloYsWuEn4J8g//EEj+95QZ4mjH+et8cy3SBK1hlrJBLmaHiExZW2qmdddkG
ZhmdWbtJK8dAj5yxpayaTgSMGZAHaJ1GdaGFhlLcQYzVpulQj6mnD/cscBPVzJ5A
FM9RQFReyo8PKKSfxNpBov4zqtRSoNaSr+xT4hbcjeI48PQZOAwqKv2wSKt5ALkm
cHcuJJluNTUcArTsTD3YvcQtcE2CYyYalz1uOVKrN6afYG6Gt8viqexzjxJFJefs
rxBFtcNLiROqAgEKsuMG33xFnNpIsbhFP4ZF4lBisIFNQe6criOvy1VpEPFLeoO9
E+1GIw3cYeYfzA7d+bxAO9eWSZyw7VZ8cOgoksxDzX+pwAh3NIS5XDp/jl3JLK3K
kiHFr/r7e7rzfXOrhe+hClb16zwqiqiD5KYD4b5mqdcrsuy1qGSe9hr+9fKgvf2Y
ZGZjpfpOCkQaIdunI8Fl8T7yQsaFIv065TbNVYnXpk8RMT98GuGCxyucXc5540sF
ZKZ57d+kJwbTGRa8i/z3QeXYTgL9//9bcEw9I9kQ6jLX9cp0R+geBLOt4RNhWasF
/8QpLuSKeiJHMWPltFZdbRo5Aiw9vpUKfQeb3DDz786AzEkWyx5M2aJZiUzkAmJA
c17Ffdwl56br9JN9oXm3FgQA7SLu0oQWtUP8HjVxDCvSaiRF15pZYxJojaiiS/Df
MMexDHS5AduMSBimz5LnsMbaL/GEv9j+TkfVYwJzhJoOiNLeiknWfVIKodv9rv4o
zed/CAGlp6bIUoib1YnuuopeWwpkS/pI9wCYfzIt/zL4z9VpjBzZkfTmbejucigO
8Tk3NTcrkZKh2n9zbuO3r9vp+7dZIrUEpe7XFqsuAdEsgn9S3aEhVCMMpFcxP1L0
DRwJiZtPBJGCxhec+54zvB7kvkqs4y8UdDcFuUgIvAIrjEjGUCQIZfaA0hSUet2a
p9MBWwIGx8IkthvsnWJ4Klnh6ixg8i8T/AJ+sqq4afhOrUDgEoNg7T+SspWNQBmr
GaO92OscZLStHBRoOk8SyR9/g1x8R4z4X3dUFlml9R2YGf61wn5X+umI8e6wZaPo
kKLuiB/sJquYvREW3lfnCsRfN9D3q90ymrP/TcAfS2pvywWclE+yuYH0wc741vMT
y9OxulplNr0X8BP3qolXsqmvrRYcolDOtbCLvUuR50lkNCWpBFSaciCK+sHpiD9c
hRrjYaTPxC3zFkD6W/g9CYPsf6YTXW1ClMpjU3pLPT42ZKA2NIEyqu1pAdADcd1f
3FBtY8wnwO0jBdHB8Uk7mZzxjLttls7oN+4iKWxPc/CtjXNIEnBzrlLWSC54t12w
4K3Jj7AekENpXSdPCKK9C6mBZq+1rSoRJcUk4KN+E5ktoTYAwbRaZG/J2CQO+cNu
EQeg3jOqGBbXAsOCq1VIXAim2SNjr1ApLMK04O8I9alf5ZUZl0ENrqpVvoT1H2by
6DaYeQ8cB4PVkwOADPa9Fah3z5KzGhfqAET8McYv9Vfmlzd0au3JKJEyo32Fu5+a
43+hWPcAtjh09Ajy7ZCeBMwqu07t9C9PT22b3H2cbaHAsDCorzCpBPZK2NTTHYO0
9+HQvDVnuUPGiDnMZYnUUOb8fBuHq5fEvRMVjVLr87nX23pHB5/ZY5jRcc23tOJr
jwSqOU6v4Znl0+YOnbYpqPnvOq0XnW54Lhb7YegPRn/tkhEFBYaCVC3PVI830ERd
icoPTQk/Rwr4asiFGMQyr7xvTqRxDJUHB09Cqi9k6EGBccj8ZSmp250aJ364L68A
G1Zkf3OD1dOzqzA+0vVYuCqOhezbEKCt0RldA1TOhMnHpa/rr1AqkNMnZSq3htvd
ofPK2NZ4e8v+ZeRUr0E73L931pVsTl71Y4oxB3dkBLei1dkfLAQCEsDUvZSwWF5C
E05bgt+CBqh6zxU9sHnDu6sN3qCHI6WgNwPxny0WPEnWq2WDC5LP4NkeCLUxE/xP
Zbb5INPgsO0NmzF3iOXOuI1CkUlxHB2B30ROqZngW+MkqLP4C8lgOqBjfKYmTh9z
ee5vKW0kfADOGADc3V/6O48M7L8/aDgxEgvY8vwJ9Bf1fjPbc1yyhOMvNYeFx3Ez
S7imWx12Riy9nSFvVhsHXFSkkIQQY4Y7m5rpcemA391S7tAX+JYdLAmt2k4n1zPH
5uv9Qw/jjhW4oC9Daz7IYxLlx447gKSeqWdmtrE+Fzi/teRk7TC8DV0RfoVKlz1Z
MP41+NNdRfc2D/6+g4dFs86ac3c1lgIzn8bnnoQme5w2k44nY2TaXUivi9isHerv
DL8oJjk5PmlWJN5u0NINHCBxySXYkciz3I6e5za15UUHcdxHTpgu5qGNfbpE3fqV
ykji7ZyrEVRC9PtX1fmxO8fiimgof2xT7IloNsj/IVUNNoFaLcGGAlhy/Oz0shJP
3a9ZulTj0v9/tRebI+GVpzLPatI02NBn5/tVl4nkuFsSng2IGThw0ujkQW9NhPlH
L0ObAKDKj4IaudfxIQv6wDXERadAcrn755ksM36WGaLiQZ/1Zx4zDL1Ae/ussBdB
dzJYh2nYxXaQ16NxRoipVoKkbBds5T0DxuosGlphvK2zRS++bpn9jR3ZBtT0qYbP
i0pJQjcs2DznnxZOha45Y6ZUdDHj2OmfCzxvZ2S4YJIM29kU9iIwDP7Ca3/wt7je
AhYXUCk/ks8AA33R9ZyrAnl4HEeUHdf0PS2U1ZFggWKxhNk1eT7Y4jUS2Fw3QGTu
QQqu1sJknEx9lFBlYnF9WHpl6ESjpIUKU5/A1j49Gwwzt2AsqTWT1Hqrk+KITKxJ
6sU9khnJ8En3rGu/34jwdFKyYgaIqfyICxl383OsiUWzvSpUAeQMETJJvmcFdLRf
pfR4L864gFDMpNnn6IAW8ylCovHeQRnlxdOk25iSTqoURsrPSgB4zewPofcaq5C2
i026hxwgd9IgAFlJ5x2ld0FZ/j+GBhV/HvI8y3yuEONhcl368oha51+UaogXuwzV
b7Mo6+MlEpu/j9aQ+lHhyZqb/uTGV5LgMwZT7A70A1hBFjbvyAXwQcBlpVxCpZ47
e9sSgyh18844jBR0I/aTlJJCG39jQBpM9gBEfm6jxmBVG7NQYUvD135uZSpQGvud
CTGBre8SKNGpVrjkzdKrFZ3gwcBNWbx2VD9j3wjIZQZmfG7tz2f9BUq27OA04cRY
0TtPp4L84FzDQi1aC2A1v9ej0AiDNlgZZbDvw10Y04YafgxWLfcHP7eA1DPW3IVV
0v1/1QX3IVE8qf6aUJgd1LQ3BA6XN5WHpEr6z0euMNKX1TYaYxkLk1sZjwAi1y8K
4QU8eHOTmZdzJ9jpi0u4ckDZ0RddYkYHzwpJoy215CXXP2CqhSq1ffic8GpbxlXb
759bHaKXGDpwywHQFHjWxlIltmuLVdbGNItQBrX7N4gcXmO3z11X9irAvAUBXPO+
E+n6edlh4FFdC9grW3JgBv1F7OvYcrlb+gvyq6cDkLJ1ITSeIoQCG6KwoXrDSN+Y
Pww4h4nYmdMXOpAi4ar/R51441r9zVGjQDyB3eenbuVx1XEilIfXlUFM7+x1ZXYz
PSGlTaFdydqL7KcWjR2+xneysFAUoJ4pvNI8gauc+nQ+GxkPUFsohnewUOq9AN0a
eEzbciIDrMnyhG2J7A+Q1wRLA9Ljwcw7lMtAyaaZW7ZT+N9gCDAE9BdvkRwew5B2
urqOh0tLUh+4/HlYWLfA22NWkbSQRFW2ilRdVxrnDor/jaaHIHdFS6U9GgxYf7Ie
KAZMqVX2HZT7QfW8jmQCyw4h+mywZQk5evMVO4wEJ8aXmJKPfWRop1xNNtXtUoY2
3wE5t2trrcCVXe4GAsTj4S8wg74XnCAXUGfL2fzKfDPQ1ARoenI5o9Or1uDFPZGS
0JuB4V3jdfXTV8BK+0mcRnj+Pyik9kKYzlvJKGk6lAVR3e0EdbxLXWUUhDYBz6qy
HWej0B7dJH4ODEer9PCrhqNA0ySv6xH6TkTS3DUPKSDc4SyhJU+k0G7iMlpt7A+7
qBTiFfzR+4Byt6f12Z3QNiS/kpt3NbUpJs7DfP0c0u/QdzYV8ftgqkvG6RSe049m
UEBGgrr2Epd1G+IQlJvNL1FeLKPsPHrT5upNz7YjsXws7KYojo2JcATloVwQvVjr
hSNKa/UMnAQgWTIllrlmAQJ50NEHggFrPPqa8iF6TkX6vL3q4BVR+zmsp2Q1X3pM
ezdpj25XZ+zxrIGcpkyNDSliahLRcozv+CtZ0wP9LzachcZwVAuBiSKpAyjUF+jK
2F/0Ds6DpNs9ooY0U4MYFCsklzlQ6gvFklCOHPIz0ZB/bVQ8Uv5qg7M8ydzx5Qb5
nefZI+GuUvHdiiP8pdo66wbb5nP0qXgHx+XU2N1Ywx3NBYB5ebR+VrVIpjVX43PC
ocR8WEAm2YYbyWzuzq0shXI7hgI0ABRnPapj9iXHLSY07QWqBsNB4mI3Z/WzQ/lQ
IwMRPhmDyFNeqdo4Qw/6hdTXZyyd4ZGoEGtMnRjp91+6wwNgLtmCx5DGkSGlMGr+
61zK0I4MCc20fkSwzCQMv9kdi0I9obH3E0GITMBvJs8J1UCoIyNGSrt2rgGOqfCN
NS6IPV4HVUuDf/LXG2bLYh0sfD7qrpdeYh0TRcXitnSjuYAOSlYVuSdaCj+VOiAT
wketo2oO4Cvf38mKf83dSHOlU//oe9izmCkR516fe+IbzBxCUxclqKx4PIbQ18DC
wf2J+s5iAvOmMbb7+yB4nk9Jb5bIqeJLoT5PvajdvT8JoSAv+yymWEiLZXVy6hHY
PRbuQFfqMsHSfNacNm6P6NSZKRsM6NqMWyVh6Ejmkz0sQtI/PXTUs/gSjwiCXEqZ
uBrENKooTSXEM1gIR8vxvtRAuZPlcrA3LI5O2S27AWK5b/Pb6HmtxWuGrxHmI54t
1fuajhKWa18FGQHtOGVEY+Tu3NVg3ciNOjBhqH2+FB7fV6sLEPGfZFOyLYnCVgnX
fOlAkRNIsBggrVhVGOKTU7Xm3DsOvEazFNTfErIxl8Q3DYEfb5ngM1WnGeEjtx4t
EJ+8fFFU+ddpwM5pdUfaiukQI8ESex46zNLp9J5mlY45Kr5aZ/GaAqT1d07EAycs
CKtJc1pfx0t87EuopI3qgqvQddhHQ7q8WLtbGdA6cSBJkxqmr3wcIhAZu41BYboC
tWq2HMOSK/0xs1p23bpZJjbFACv7QhWsYOPcBgWm83B28q3z0iiJm1Ay42o4lYSo
a6dc6N5w8l0/DYdz7YIQls/K2859v/4mMDIfFlMcIOebDViSacvJK3c8/P3ttE4M
ULDbmx6mDUV8H1JtmTTIl9jUZdO4fr92PbQmAv/W21KFwwIA4/PEP5pNR4YqlGNW
01WERnahqIH/mC/FRa3ipaTrp+j8KJvpB8btpHXTi/klx5WjLjFce7gph80Flg1R
2WySFDCG65lmT5qg6/uM1PsigdopOg3M/Iq/Lspc5XItN8qwow4NMZFfLC02iRdX
YfK7DqrqKw2W8Tj40HNCqmjsB/N84ObvJDp6OSFFFlqjSC2eAwH3McApFrd0UEBE
GcE8gAFmHsczRCzMyLn+fLX4zr/yLUIveQQlrQfDkoy7cEMDlPglaiY0ARQ2If/z
DEeDWK0VrC+aP5Y6jPo20x/NJEBRpwhu1p2ULCqRmZ7kGMk3hlwqdd5/NDXZjxuZ
MoDoh3x1sGRcneVQB1HIt+ujYygOxBSaGrrq2MdpsiPDQxycbQPKpwW5KBLdS4Rq
6suSDLSn2pXYyh59z73k6lvnmEP9YjFmai7CU8B3DBqVzUP+wtbFC1jp9BFgiw6Q
tbsQaup9AZUHzgmVuT6Ri9Sw9DUgepHUZuwTlU9Gm+ZwsGbGdts09t+BX3DcRkBw
FlcU4W5qDtd1iKdPDmPSyxrLs3XAK6zBHPVmll4q+fA+Jd02b/EwWfF0OrcmS7Vk
ZgequuKmfzAiK0HgALPF5bXqO0jUavKhO5cQvvOwEOdPWr9nNl7c25RsPFg5tNTE
yXEUgM8GJoEsuOngTCcwU7jGBFkL2Y5MPV/PWGd/n5EztX2/QHW17ZzUqlmagduo
lk8lXKn40d+OXZr0p9Mwgc1VIywagdwuoIh1xcFk4xH+5zG8qL1TT+JqF7wav3W6
Lhz+0YV5UumJISUg0uuE+iLg16JD9N3NPqILmxL+zv6CQxrsv/rFilOIsKjtqVhc
7WTYW2u7uM1O37IirOKSLLcfXfDhFxeXBxnGSu2o/oRQQBN64tqcbCxTVmEcCm4s
k8Fkqu1OCFgbCzcLR5fen6yIv+aZm7noEpdzutXqT+Yba3Z+6dWqVTMoqM6ZnaJs
taSKmmQiL/9r3yu2X1eWkFxONEM3736KwqYvKPjb4hUiOanakbEO6pllsYzAvlK+
IAX05m36vvsbVq7CeZ38R+0MenGzXTHswsrw0TXClqHJY6YeNqkHxDIGeZ+DlcNS
VD8U5NlUmv+PqSi8MRTo0tTqKo6RTD93nlraXumQ+GDh3YSzfgHg6fHwguWV5F9R
SEb4SaF8JBgVcm6T1/8R1p4GTiN7ZDltHMf20F8eZwoTPz77aUWnQr/LY+EE7/p4
KDMP2WPTVihce0hGLB2AogF59/W/2wBQ+Wjng2t901IavXTkN6I2NEmk5d2U48Ga
3KR6fQmnN1+PIknbeqtMZ0pCnYsxyhfXaYIqx29ZEqtUfjQ3smO1eQc1VrZWY/rp
oSvggjSX47H23ckKeYjqbKQs+vn6AEU/SSDCCwNztgfvImetoLo1tgOKSfOPI49c
jPgjQjq1m3Xohxn34mI4kBJ/hbNB0YdWZeHcFrnt9Y+vWxWWD4jnEDfAxIbhPhFj
neHTLIIadLzn6dUAVbaJnLwwPr/ZRFeXXKeusfCW8WLxKC7D1IBKj4UdqC1t8+it
4uCFSHZ/QRwBuVM6Rc8B24r/wfb5UCjGgAuN7O7XPQpDG0hZbN53uwK4yhyHlc0u
g0HAwZKeQKuHA6O4oMeEeONv2mkU71GjurGmGQkqLnFhSs3WPKmqkFEmkSD2rd63
/b8NOnPBZlzedxAcjykpgZLPNIzh1rTAAWHsCC4RwkzOo/heYqwr/P28CRvzPl1B
VBWz222JN0ITO3TvCOt4sLTxMXtRArW7smpUwSGU2vE0emySN/XhYn8M/6xzVady
ruwN+gZAvZiywLzq8Pc8P2H68/A8fehnNtvFf9Jfh5J3hJe9VUHOG/gNdci5N7dS
y2Vl+QWpvVKvQ43s6N9sz0nRCVSbS/R/oVeawQz0Ipj5rl3iG8IUY1g/R2BNbVCL
3gDRoozmmwic0cwSskVdsf2gU4uEzrtY1TaXQjvmFYZRAn4zwByY7eXmVRdU+WRP
kBBSCemiOPYXTf4tEoiSM8gmtzepGN68ts+uiUI+DSiYu8vf929x/ADPBKgBuJ0N
AVz+cIZ0eTTR0d2N+63mkeQjKcu3xql4wUudXct+5I2nfu4i1U5lJmmGX+Nr87Sl
r4BIp7P1ZqjBamKbtoIcWRBhbGUHhrMqFsfbn4dYnX/9V8BV6eDPsJMjDWUFZ1Sc
cM9+iEyslEvCAuYC0LUTDA2TB7G91O/gB2TcUkkKep2fPKGHXCneVG52Y46PF///
/45v/fAlVCeKBM0WJiH1L3kwWF7VGC4L9s72nTNr+M1voyTYe0VdcVuqbNNcIvGu
w27X1AHOgYc+95knZ0o10AHeM1INTo3itX1QshM0KD3lVWSM2SbxElXQiy4xloIx
uBEsz6KMD4by9QHJLsmS2agWMvJyewzOPBUx2oZAWHdx9og3xHcgchvRnBMaspNd
Al+iUobFCcEkrx/I39kg/XdmQSYrBAoNWJWd78CWa9FQZtNjmhnCV5PLSt60T/E2
y/0fjYeRhp3vSQIQRnYzmAcJEwy3/Bw3boLcOkwfdKktJKxhmWFA465DMGSzp+5q
Nhnrnb+jzGBq1uB9ZlhP4KyhewamsAq2W4XziIxDJSsrRJ5GEVuc42I22d7240b+
2ZaIRMhNPHlMJuZe8oVeMmhIRgI96nZwaiwXmK+mFoxUDB99gxpy/4tVI3ZWnTF6
ny3XyBX9ItrArYj48nrNEy1vC46BvUvHeUelTrLm0u8LrN9BXRMHsaMQWrozl4pc
/AitBF2FcPNrqYXVjidFDbCrvilV+MLMMPGG052fps0XqAAV1MLkSWBpPrLOADhX
/YnKQm6GgalXkt3LFuHTgqA66NHoTtuDBpWCXBXn2a7+WYN0cXhFiuvEuEVP3I17
b1WvzjX8gFxqg8kMpBg0fDVg8FB5yVfOt2Gvs4MZDCUDkBSaMNWXsuCaCOHvI6cg
VRWBQyL3FrCn3zbUHjQ86JzRsZCCQ1CmwKm0bwV9VFmowlyQptLGkCP/pgtfd60S
+yFX7rzsg3WGuWehAGNlmt/TBYv0aXC2plmtnNaDDyyIl7iFpRT3XoJXJ1RK8JUp
eR+7N4lYSpaM771puWSgKA3pHTLACtjLneYSWhv4ERUnJsfQGnkEFmSeTxnomFtz
2ifX46uYgepTkBc3DEQvqh5YwPaBE5zfNFn5sDywEWV+mSu/9MT2KX+dkkDk1WA8
cJncdkO8ErLu5xz9QVAfxYArcuPgTZ+80YyV4fO6kbW3aRfW1hsZQ1qyXfzNMcuH
BHc346Sq3C+XjAkYMKwoazG4jDxhvC58VyFWGHNQyVzHxmoPgdNUpdx+07PSNLru
uelRFMCxLsObSWd/uLLarpFoiGpeT8hwhCbWkWECYTJ3XnHExCNNq+UmU/DVvvUI
D5bFwx6nz0c54m0D3/K+suzIX/w+iVsNV0xKxbPeaLuHjCRYlmHyxeyrNYMRw6KC
mM8TBhLhNL7Ri1dPugsi4ulBG3xMm/1akaMtnYaryeI6lh0e/McFRFOSz2IumBYP
859l8aWFjOHqcPSXu1X61fNlKFyrMVl6tY9EssWlzQQyum7TAfTsfA6LnPF9uR/8
jTGzNifF+YqLZ4lexo/y36qjNGQ0YSkSP8H2benDU87fNOTyZ1cEyyIgGf7hUqxq
PhxeaSIdVg8x8EOcx9AQ6whSFDP7Mb4PNXm2a5kystDfeA2KxRSX+F55Lt/aUIsg
Uw6uzbKlfzLoORJVKcS1feTkNFZdUU0pdPnBwEZVkkuHH+Y8qXRQo958GQqd9rAh
eR3RAbCS60zHzekM2cocwNTpYcFuAJASKsdQgU+41XU01uJxcufdLbSddWgO599X
pFBFi56A1H81OijpzoUk3JF4Cid6w01yz3V+EhB2SlnXfTnVk+3RJkQPoEUcCLWT
3H4R2tCZnOwuCswIx4PsfNnsPRHGHlPNkrzGFUnuJ/qUBC5M5GMWhmG3xSUpU3wB
t2tDZPKJtiUpVuQ2sLHuMe8Ugu/E+bHzhI23RjgR0fSCASoNYQuX6yG8VSUabxQy
AyxaYSxqxxKJlGvHJUd5e1TqkdAonTIFV60a6kB7bpjGouKwwRZ1HQRnoUKVqGMs
6zAQD4p2psWRKxD95j8hvxMFvqAPRL6SbVzCDQD9RnFLPjtzGR7B98en82QVLRk8
w6gDHsMk58wkmaB0cRZKmTIcfKYz5o+orzf5qCJaUEsAlyJsucSNheDly+FpKtFo
0JVKfS4TkZya4UNpvAJmT48/gKrys0Fm4xQuBulLHbBcvpT77hj+W7Q2NUQBQzkx
JVavtKxVDm/p6zf+A7qBtM4qsAbsO+Ou5B3qy071uLCkkwZE/OXIuXsXDGKdPhBs
q0hLxMquOeWGPz7R6S8yhDpuLCcEVfmlakW/4pJGKdkhwXhcNDZ/l5RHmnOMGpVm
969bFDJCgGw9z0YJuoOH3e3trDDVn039PjKST41TkkmZMpVtivWVaGtIg+F5irgL
uVkgt0vc7bhWi/7vC478QiWAZchNzm+0/EKpdrZnTBDpqemnA4gx3Lpsq3EhCTQF
jFMn6EkaNyvKA3jqc6ej+VfS5DeFZicYiPQOedcrV2PbLYoRB1OpJIWUydQtoO4f
Oz531sd8ylb6bqfW/HG6maFSCFjLYDOxMU8ctw3Za96CX2+3UejB6DJlsHjof9m3
I6n/A32C49Uoi2GxsbMzG136z9QW1ohu1i0x5NS6GRkFuWERFGs1sOTKeXKf5W+J
Km9d07c78OjC51/40SPpgzQJDfLmDm/O8lye/tYcQVzovnrSuKDpQSkcJPHpFLmn
qaYqh4IAS3YEHOnLtviIRGMNmmKlmk/GQhnToei2Zr0EcmkcCUXypGWkZcA36/ab
ZAkMPC43SqYgQmYrb5Kug7cn8kPMJRbJ6SBIqgp9oRUAh/+1ojqGb1LCNTgfShc9
Xs6Cr0Rk4c685Tj8T78DIY+auxhG5CRx9dB359+z2lS98jueprhwBTdZCbS1L22C
F04nI8SaVB13v+fwvocuErLEKatONoIz4vfFQR2EGmbbLpozSFOS62YUDr5ecoaO
ZAeCD9qNiBGOYSyeE00AIEuqCAA3fv7C+4aWoyCSqL572nbLXSI8CN7dslbw+Vzk
VJeD8Gx3uEBHeoH1ICc5T+AoiHhqDP9F//VNRIptG3OGJenpD2Aa6+hxgJpeO+q3
iRIZ7zkYirEvAMSwFAUHxEo6IqYM0v1G8cMchIumFmA1WMocJ/hltw7/HjWbp3Nl
GlOnpMQ3d4CHmpWMcgDo4K/kxSuOjG+mE1t4XunOsekaA9V3IZZUeY4ILxD9EReo
U5rxdXCE3qpKyQMKjEIzUpwDuPCjOVymSnGyXtxh4KDeFTWycTCqN1XJQ0w5ps7g
YUNo6IIYI5a1BfafrHbB/m2j3Yg4RGvTcEXRoRkyZaxGobVUMt3dqFvrWMkxJWu7
7jDhwq5rQuG354upZSrmMddv8hJEoAlu4QsNJrE+oYbSUAZj4CJEHRNQ7FigUIoQ
sd015cJZ8oOrSevvVPDdQnso3iqXYn5j74UfmIGhUsJFKPEFEijnF5jUzYufjNEj
vcef9OviuCo3iqC65a9qMlX8MAAmx1rFa3kM63VEgfrhyiYQNcdvW4Aqg3xDMcpK
JfVDsjt80PwrWBiUa7x84zusJBF4RXcUcShijz4VwVEF2zLDKt5d06ACoRUDbT3i
m3BWJLeAexQsm1T5dxxkgK5ai9THTp09jz9FZ7AKFHV8iSCUuHMe8TFG+I14IwnU
Oz08uYI3Grm3FdH2ObP1lqCCHixp2hgsXujSY8SCqNfyr7WHmM7ZE6MtU35JUeV4
ya/RW4j1IZfjbT6FR46St5+VfoC6yNzipPvA+rVnNo895VsKY21p7ztvUXhmk8kW
m9gli7SLj3mLD9duNY8uaWF0WcaDbDNTER59auS3/1zRYQEN6cyhkim8Uq46O/gK
KZ5D+8R9N6HhnO3y5GpoBjA8WfdG2hBJAdgbqOqMKKDYbBXBKBRRnoA7vx++xW2R
4bp0h6/rMZMGPeUmi/sIgt/EoobGt6x94vfAegFhnRqu7n1fHtnGjGHzfSKnSMp2
wMI8ABo7KsR677N6sabBoQULefyFw38u5G40Tk8dIgBgsWQGGGxHAx4szeTWKVjH
0mBsfV+fD+xtwrDYPjA3tLViEUei/W6Hwil8X96XDMWImVJErs7IOh1Pu4Q18jBv
Md8kJslg32SkClJB9dwfCfCIofw4I9VafmvOwTXZHFe9n/LRu1ikPi2yxAQNq239
YC6ozR8tmrmfMuERASX3aTirHuer/Bv+kbPR4bLv6NWZtk6YfJE2KUgb3BnwQfBx
QXy1UiBP0bkMufgG44rigBMAN5ugiGN5wdcYV9p00wAV1IZbCBDEj1CsRs1I5IJ8
C8YXz/TUM5KctN2cBLIHkpxsjeKpnEgZp82rAaCZnuxY/arF/QU8tIBibNGpjUwa
29+t1RjnkC8JJGV3vEZDW0mBymLwWpUalpBN3Zk1+JPfxHhzoiYKnkurfqwf8eZs
Q6ITJLRrh1LUruWra4chcC140SosOq9mIXeX+4pziBd3LrqjamaKUdHmtmoX6fn9
Ipv0yNt5uJTicTAzxmr+1xWLOdg5mFW/yBc+dS4PDhxcY86au8RclobW5cEfld9X
QYOca4DGF4UIm9bFKyzg5kal51gWM+nBSa0WqJZMg7ceIe3vt+FRmvkkb23V/Mht
qtzFQmhaYG3rZqpIzwcE580NTSxDAYpD8l6gmQtaaFEUnszx7rmeQz1dNExK+qmj
FKZ7iU9wd+VuGC1f63iuL30UBfbUnHMTBB52COgIPns6OzcNjcJawnhbjdNDkWts
wzl0on81ct6bJ85adwkIPCftomZldfXztQS2FAE4JwoEuBCw0uKHV+cK7L+n/QXE
Kslcb/eZYLvMmAUlzAzJt7hEyg9EHnEYkxV/m3k+fYKZLwgGeFtO4uacifvCdH0k
Ql3iYpj3ONSjDbKiaQ18c21oA7NkeyZeXnTB5zvj4JQ7hY/xAI5qmYlYaHWAocen
QMk3tAZmUy5f9xYHzqn0HW6LI9ZB0ts8d3aM5HmYVEjHu9t7JkwkjoJi+g/+9XTz
KMPzrXHaTeWSKok2F86Ni4yiroqYPOiet69Yd8EsQPFTqHBv9bkTcTy1pxQuhe4Z
aNx3n2n4B9nX35oVYxwHqc6ALMx+2laUBb2+0p7IIMCqah/2rmmbEcnxxss5paZi
pfi7I1kNI9zidYgfb4U122VirboUNdE3MENYTbPfvDPQ0QRgrCugev6NULruUVUo
oJlzmt6rVIvWj17RCI5CcPztoPaKbX4cnUUJY4O7/NdfuDtNOpjYwlZ7kcdvnvbV
Kr13KmaPouvZ8WSDVmeqSRgqgDDWQuZnp/t1u0TfztNGpUbGfJ6ZwYh50s+qpEMB
OScHoK8Wiar9+bVx7XaZ2sGN+1/tjeiJoQdX9OO2o6XcPFaFcBEdPalJfipvAw4Q
Gs6t12bb2ZqndqcvW3DTq4kZiYtot8++Iem6IW3kpteBj/gUjEwUu4v4gE6OdB/L
6XRiE7CpGnf8llkGi6RZquYhVZvXNe33Ep/+b/1o8rvIuD53yCk9GvUbp9SjU8Q7
g1WutpV0UuuPTmEJlTIYHMxUiJaqlBImO9fDErEpiYlVavQcPXx+85G5tsUFhpvl
hp8M1BSy0DO7nRzoNyLUT/g5ZPa5TTY2OggTUFndnI03AgEtWS5MMqVcREuLL2UZ
UvaC8coiWPhj5ERQ5WM0EVah0KKkovl6UdhVmojsaFxx5KdtQUsCfruCoDFyb9Y8
0QNBkPumebralAD+zNDI5i+In0g0O1O5wUBMN+IZcxm1H7PK6q8zew4Sqej6aK0J
HAz/4nXaYfeWDdPXBZJc9kvrR7omi5CSkUqLC+GJGYV2+FWLuzHCU7IYjLq1ISus
9HdDM69+ucQIerpoC6zQSjb9neT7JuZf5Cib5rZ5WPnsbDIC0032j5gcfQw0+mSk
klRVF/EQ4BEVnGpI5l2Uw61C/YQ6knh1XZztISax7mExjpHbdoWt746dyC1a4Nlt
oWNpWdI/Fkr/4Srz5hqqHtDa7EvsTK5El/GnBBZbYJYm46I2GDQHynp/0T/folRr
mXt05XbwEn52hVRzln2oMjTt7l7jwKypZAvMwDRAGcK38Dj/OyjZcZXB6SkkQ23U
lw3b20ng42G5xvoBiNY6N6Xo8IXdU7x7OmOpz0J5T7EFNcoMiayj329rrXhkAhBX
81QPcBwAASSbv7CZ4Rk2qdIW0JP7zrk77CgYh4ALVnAfarM9kKkbDjWhKzCruDeN
lK68d/3SceprV1zm1Vxn/RMGNeVBdobpQDDnQhexutfNvHFMSmhDVL4J1IYuXD/k
VzErdwtC4f8puBMgEqDwG3DjKsOAmD43QhhbSe17nxwmLzWC+Kl5wYqdzKNMNtzQ
AEnJz/ennrx/xLqAVGJ9aQwRCBmouPAoNRlF4AVeqVjMxHsx30pAdwG+wDlGrStF
dzUYmfG6AS1vJ8FuMtOp6/Kcl5Bknt0DKoVkzLDOgXY7d+6l2bxUYm2SHPOO4V7+
jFCzV/XGBYU98lLUE/LcRSdsEA6TKILcOk+NTm86OCWVKVPj0fEF0nmdXloSe7Wt
kYFvK4z4cOveTJ+YiwRhesnsRnFQr/8tyMeultTDk7XiO7ZyXPe2qurKauLTgC/f
HGt5NVDcclNlQC3TwNeZ4Vh0d0+09yJYRs/9eDaR0UxoMLLpVYX695dYkSmrOjWx
2rUZ1jZ/3mJhBayxmbp5J3VYDF5E2zip6taned1HPX0z3lX03PkZ+VcIJ/o1iSbe
t5reG3+hAJQ6jWOF9z/vtHIJBXKjabxVdWN9Got2Siqc0ou16S87tMR9oAUp4zia
uwyA1ufVYYl9HGPM6EbQdPoBeH5tYzQRjn+WsDh+V7CnyUHRpXaBZpiL+LpvUy14
SS1fICmAQI7GQBBcnXI5qbjR5BrRuzbkJm1wgK+EzACgGLDRedUBXtZBuJtaxLLm
3F/hxxqMntJVl+K2phDmBcChiwQGXWesWaJmdfAiAlExXheMRg+WTjLRW6mZUeZe
fPkfIrhRkktVY/s4I1lLp2jQcHC9zyb7QYYCv3ZeeJAYWtkjNMQo2rZCWCgRhTQp
wETYMo4y3FEm0/WpuGuqnlrx611rCIupxIiZnqoztsBPyov17uhWN6ePMcYOwop6
ZoxvrzvEv6EUfFOE0RUYg0u0XrfYc8FAePH8IwbJiWqSuSQnZcu9qChMWZ8Mmtz5
GhwHq5cw+iZ4LYMrINC+qT/nvqX443l8pspEz74qBao/1DMny8CjNvNb4sOeAT2a
GHrVR9KrKooGy5ra2JsulYreVF07HSfh51ou3hXrOoVFuOZteLsWrwZA4HffLWbN
KO8fH9ATz4AznZz5yBuwywD3bSFd9kg+P5L4Ft8DNkVUqVQK0R9/T2c++7R5L0DW
XoEdfzE/MzQEJl8HAZD7d3BJsN3bMbcKzEXARna46nJez1DggkaApvAPjfbkMhAS
eKtdd8OhXBRyi4WVzbesUvHTB6AOOjc/c7GbDNKV5xrSn25HyV1bLycXeEjmku2O
KdFdClNbRhdXfW3A8pEd8H5ZrgGagTZaamUUaAST7ChB/prGAiOaKLnbrRef0na4
bqL3bOnKsbVWDOynO/4H+CYHB2c7LB0/tpJoX2aWF+tOofDflmOnzrESE0BgThA3
sfJ329/SHFJ6llBz5xci49IGtT2jtktOg4gU9vL/1yT0DF0Au1hrKMxC/4om82IE
eoJXZIp+ocykJ9GiEhLSZqs2jOADM9BXHL00V3xfs2SiSs+dVs2cM1dm0fRanfH4
EL0F4bh0TIEvfrt36XyFz+GP4qhVrerT2hhKLoFTdeXpJOluOtBOrcxx0+nkJ0gb
LGc+42jUeZQ3nkSHzdZ3/VidUNC4GIJnj32M7QodStVKEIPbhZGVaK7NerNuAct1
oICzpf/41nMKjx64fgAkt7qZ6OyyyOqO/eMlh9wZu2bOYJL3tfse0LuVcBRo1EvS
j2U+wKXhzT0ntmh+CIOsVCMoQTC9+gHxHmxAmFpKxvchcXz59/vOnjC0irzRkZAp
S/fySXT+3t2sTOXWhvseKJEv0QSDqTUXlUvbPaM0Bqhw7C3SYwiMOoh7txQ2Zj7p
Wg+jhZPAq58tAcIG0zVz2/UlN0wIrSftypjs+SEifli4E6ptTLcHi+6NEJYC1Ycx
ldf5FC/Em/ltMohwg3ZnG+avamPVw6uwdziN5zGnl7PCWnvhY3bP4TPB+IZUdXxU
OcEKmKgmDpQ0nzhaphJnE6fE641KLci7ONOPqDzg0nkpK515Tnankr3kOyNkgsDY
EvsDZ870nww7aWd6pi9AcYqn1Djx+GhVVJguMee0OHRHRdprK6HSVUcuMaRnCmYz
oX97P/j/4wXuxRf7oZ4ZZ4TdAWeqESVyfRo9u075muPrAuxwjPsgVXe7586D32/Z
TgadowctSt7/VvCjHDyx1Fj105ICx/tNCD34NbxwXtwQuf0P4MZpJ9TlzhM5cHqD
8EaCTqpYaGEu54tyljbBM4ceRmdjSdNiI5v3O9a3V1LEtRwySH7Nk3rvzmARDlmW
J3XEyZMw/81IuFRQZjyvXpxnM6/dsEdYpxgOKPhn89wBCgtCzonY6ThIjKN4+Y+O
Krqg6/eqbauFi/G0icUO/WGj4Z7IJT4dIZRpVTl7CQ5TDFElyNvARB/4CWUBf4LD
+kvGxfrcbmwlu5BJ+7G1IianxVVQhgq8Q7t+MgZXI2TtydGR/hV/ZAisXBX4mRrf
II+TiClmiU5ragWelTzwjvZHyrd5XAPFoTj/BghnfURsEQnGtI6hzhD+yHJm6/Ow
dE2ADM4bY25/NVlNPyFv+TIYWmDflQpBx+ncJZUrzsFyfGgLG16YuwVKmhGqTutt
WjrMAU9JihvJS91mYdavsxnPYhma7xnrISd9j5MmBMHW3+Eu7FrRvfOwIj61bNKr
ffJrVC8xMTUG8QHSuXP+RxjVvMYR/lHtY85nfg6vox51cfXdK/gb2vL4/kqAQi3z
CLDi2kaRx5sOd6hviIqaiykdgc4HVCqMDgAKABFwdNQwZNWEhASf7dygW7ASk4FK
5PS0SUHRIh+LG//qm/vkPlpH/sRWWqUNH0mOdLbkN+fokIwd+XBT8VM2HpProHhH
h+wL4JnRBLxVvCCpmTk1EauRg9faB9rImVX62lGLuITLwo31x8wutOYYjS+xDMHB
XjGdxXKIQMnmSrosk5983Y/cSthayybDkdGAlwys03W4F8OZ8rc8hkFH7HqFMAZ6
vmYBq0oiElLqnvjozoubNRzwaXSdl2efwfuHIk794/rmT4gMBY3OAuItgFUvTiSi
W0K+fu/92eUDd/zFfZhZLLCtMp+oX7Gsdkp9uqE186k+z5bb3LirOYVCk+/LPp/1
YpyQvgPIIu1XtABJSAjlEkZRhNejH+ackhczuYNnvI3Vg8Y1OGxmF80QCSefBuFS
/Vm/aLOH1K4N1cMccrkeLYGgap1nULePesKQnqK61xkYnAP5oEztHNjX+mqZKRtc
chl3Kyu6mKuSh8gROQZTkLEUdWZU9uxFi67bJ/GJSSAwWZ/jD8/OWUs4NpXFq1Sz
6QDGc8YEzO8OMKZ2A4BomE5BnIao695Rz7Gl6P/1IgGuMgP2gjb1xktGfoqn9QBy
MpQEur5U1Ttxs+8oKlEarmKSVES/5rn0GCchzjIbzKv6IOPy1bW5ZWnysUsyVQnL
n3c6XLVsbYdFZiFxSd7uREKrNePNRjnaQDQIjBwGT5X1sksMrVQHbB86HmGx28kE
OiMhoTHuNCkbxqiZYfW62ShcaH94gvygjNO4dxMFyDRdvkT0jFyp7XcIjQcSIbNW
aeUZ0Ea8zlPYHj/shaipz5eyYO7cQHm3Wz6qAucl1fDXrVhx+9Rt2lUwOD1g7U6u
TwRcXAo49f7pDkSxmMKc8xaiDa+Opszsex/ldKDWoy3O6qL72aOFS7uiBGIoks2U
+/PE6dy2E9Lb0RwIJj5vv6m8DXjPB0WiYKioCZbzL7ILbg6S7BUtnJbIYiMdPF/p
ILpXmoao7+EbV7HsWwrBIEhw+OYdIs3mVYlTEb9gTyTRUP5UJZJ7tUUERw8RP0G/
bUFJcTTm4C+BePF6aNFZQl9etoKcqVSALshIN/M5xR56Cd2iDqyLuUfCXyGbIbEE
qcWZq6SSzDI+hdppkJX7DyE0PNiH8x7ASCNSWmoXGSI3PVHRM/VFPUVgyAjB1Lr6
SwMhgyHTuEjCIpK1hKluCuIwTiUCt1claz4LbSgxYZK4YdLvUQsweu2xrw8Itm5L
nlfykwnqJqyiZpYVoKPFTPNqOump8P7KbX+9gHDhrkGhyHg6Z1VF+ZhjYKIBL/FF
PFNUNH8UGgbz/UUK84eQNiKX2TU9H77YODFv4CMYBZd2F1+lyAF3RsRl58NZLyP5
qzWN6n3pMq8ek02t1fqm0FPe3YPZYGgcEdU/AHeuI1gx1jFaUSCY9qpupruBI33V
5INgptSxeQz0F0lD2a+hztP8Y6r3F0NzzZ5/r/WjgCvJKvASd66W1AFfT+V1tPod
bixf9rgF+9S8jmcORCjthN+31XVOXKwtPtLTVpFusFIJ80jey7RQHaQ76i7qi/01
jS86366NjhZvNcl5F5jKozBxPPmjaSs06uqqLVxenocLlV56ij3zpH/HMj5kDTxJ
x4Yt8yEML8tsAqVHT7Y8UYX6dCUSwAqkcDARO96rgHu6buZnz4wUepNaiYNFOiua
LWhzDKb+Rmcd9+Cag4QScN1Teunj6ZM2MB1ine9YfczCh/6kRoqYtd5/Kj9EtD8v
Wd+iVQfew5v60IY2CofL9O2zC79tlUem1G6L2rJvveE3S6xjy8mA00MSkrm2o9CW
ZrVKHECZyHKL2OTvJC6eEp3HVfz/1N56j5BIY03yX9nh46b5TyKDQSXOqCxKBFgf
zVtWfY2DlVN72Wald+4rqXQ98ZjMbteG5gz4eqE1XM7Q75pikCVxk/DyA4vx5NmQ
qRSDr0oe2Xl690S/b4F6QuA1iru8oG9bLZNO7ByV7DbL+TSUDAJcaYXio77bsyry
oo7h6mqLmZAgaf+aY6q1K/K+qhh6Bj6MB+rktiT4OBaEziANdHXHKFRfEg1AWmyf
13HbzVuzF+M8/iPuGZthP5485/x+qUOhKVtcxOrYPj9C5XpftuG1S2tt1fFXV9Te
obR3Wbev0UKDoNgy21+eBkOTLonmC+EZ01F6vsliapjWnoBeVE9MlX0bxI+zDqpG
nxSFLPTm3s6WiTWXSgcWZeMR76YZre0XBbnIZi2MMWN5rvyxzGXW6NdwSW/wHnHw
zhhPhiRRCiElOVYWOIipbmfzZ+qG+67V0+kwdBwDPAYM8f79oNPFeSn69b6bE6PX
kQ7rWVzHsE7TT6N8IKC4wFzzcbkmTDhNWrQoS62bLhDZiAQ7e55nGNG5Q5CowfJW
b/S+J49t0gPkJpLT8tC3bSF7L6lPwI89yw5qqhmwTqkvX2WnsavJ+BI/PK4UC5ci
6gTH7eMMzgTAcuQE8bquS60DDxRRx68AuhJNKwSQVXCFjedAqhWQv6b+jsU250rS
2dzRBtzE/3xrYV4bmGasmrX96VyFv0iWbj3GuUfZ6VrdFbFBeBHI7j3O73979P/a
ypklXApyJPxGYyTbwEt8VxRzbbLb6tnzFPdkxxyv0dVMu4h9IOPaxqW3n9922cNL
BuFJaGgcJi8sJEADFcCxuaY0T0CSp2CK2ehhI+kJbLSxs6pCy3oSTGfyaK+4otXD
gfUkR4CygO4R0yKE6F6D8yICIWtXecpiyFaCB36/km3pTOGYDDgtJWn6XxJ0Mb+G
y98AE3TfioXgYTWPe3/outy8AgYbVR0KA9l9JIc7V/FaLXO9W9XP+lvdXdsPEQl9
9cDp2oFclaZhslJVW3hJ5arw3ESP/d9KuXphRd5gQABP3+M626F+Z7HZmie1Js8y
/rqeUQ6WpMqWz75VYOtE/gNlcW6rhyG88E9Ns478URd6ysDkSsAz6OpfEn2KiYgb
4FWemhQZrWKQRne2mbrHJx6ZvZk5dlEw71qqa6x7a3Oi1nUwMThfwGfD9yqqf4RB
eLckDFibKNqCWnjq8TNtjYziHcNxgeJh9ta1D4LGxb8gM8/obpzcO2RF0KwP93qy
Bpc9hgbWp8L+i6tZGoxwlREmpR/AnFpLE09NjJ1ZpvZWOXi/GKLQLF2N7mzzh0lz
F2skD7jfr9zcYVHZkf3dueukUwgREJV7RBcoYTjtzlEGFYVcptraNPIbYSt5gjZK
ukKUPeYZg07fWiLMbZerjQqwhHWtne9qb0VM1SNzkB5WvT9JuMXxT739NQvB783P
Ucb7mnW/OC9/2j9f1CxfPtOYHQZb9vk90UeWLi3nTp7QIbJ1jogVwp0S0vuMk24l
Cauej5322ZOQzjNzMSTANau8pdgsePdIWJmpp8tdanqcflYqTHR7IhNpRwql05oA
N4QIsKDUB7gNwBp4o7NtZwmNrJsnRCpZbZSef0k3cMybzY6fiKGD10M5IwoirQ+t
uXUaqFDl9040OifGs/VOvzFs9nilK5PmS3GJTl/epdKK1viCbuRfhHmGtd2cihfD
BiUMLi0AX+nQocmua4iZ0VocgK3XEa4JMdXTatVbvFbRcJ3UCBwW3BG80RXtLL+I
CqaZFnEdq0T5xFWrCmbwfGDeq9RhPMF6CJPPuvrv3Y+3YvW45Ono3T8ox5S7HSgy
TltU6wv7ErO73SSVGGmmUNLgVrs1WZOO48zGS7120bNeVYDYNVPFewoyflK+cMaE
vI+z0xscVFTRy0OdOl98CMwwvvQjoLPINk3AgtrKTPgMXSHOq1YcQ8xJcHrl3QBZ
3BKU/CUdWy39f9134/BxzdpMgtwLmRA5er1aET9/arL+bWzoMuOef61ySC95L8ID
SbJxu/zsi0Bcw85W9fJeHfspBnFEhuyAfiU/J51fPAxZJ79EVbG2YKa/HVxPMjTn
4ikBjbkhvqlGkJPtn2Aa3RNDSLjZhUEu0eSoNrdVZq87gdsD1KuVYLWlnWk7koBx
QqiNpe6U/qyknGys8IQTAuEoQXyr+1fIDi5rbe34d82/h8E+6yvcKoLPqc6e6K68
wxWR/v62Nf5EWg6hk0F88eltEb/I7ik1hOwS+qxgH7KEDNgRqcpBM9wy2N/qm2aY
iEg3Vrk8q5g6ztnjC/v1XhQZy1ZOsQiC+aQb0jS1/0RD918iqWyyw4oehXp1+3uC
Rs0ZpAYBAK1qcjvf1o15yg3akDzCWtE1QTR8q0Tyt6iQAEgspvGOOj72UZW0WMC/
XvGIP+qmhmhFB8Xh5ww0W6jXWCPunJdI0WerhnJ7jdNFwUst8rThRuA2bq/jMJXF
NTvbrZLcIPtH2P9xRknDtPA7rxwCJpfYwnLa1Ux9WhFLGJuzD5R+tlVJNM7ONhIp
SFcmdrJYF4IeXO8bu/1R0Rwux9QuxWF57OpvuVykHsFSsHGsFoUWqGxNmgs+RYAc
0NeGT2CuUYoqovyMG/sU0vtoiKj0V3zUo59V1C9HbsDmQRAZIqTCCYAr/M1pgkFg
X6p4ZkKN10OC9P5Fy+nofwkP8GWHhTcnRXeNhO6u3N2QkYQp3k3WWLpHk60yfr2T
9RfQfciYDB7ULHW4H0e/2X2XrrdJrygG/+7JolSHAYe6ApEJrQZKd/6BxG/GO9ZT
K+qasgBW2ngA7hXMaaXfQSc+kb/vpwMD24cjJ/ErhjbIunRC5M5voQLnWlbS06FV
le0VWG24GO00lpvbOJgOA1+uDPifDsWo3f3giJExvQ8VnY3iGG2cji5p7YV9pFSY
RU41j2nkzd4K96UOAsTXftrwmUKpVe6hY8a+v2rhRcfZBjKrYa1K8ai7RV4FHyHe
eq5Xiq87nYW1YFvEYjS0K8UZfgGrxJlX8jT1U8nmI6ZeEkG9RTTkjYbGiXoUNNWw
vr7TDJ4qsIiPKM17rI1veVFIaaMPlFV9LqRx7eGUmQSWNjUBKVzlq3F9TmYYiZkN
w4utHDGTTGi18wcoSUjJke6nGF4YlCVhRwFw40cj5+hnVRlCEc89eJqkrFeb9Je6
JKd7pyrpYaFxiwajnmAlUsLtqktQadGKbYROANiPRkZlti4EMKjUjYJwwgrm2mop
c6JTXzQD7Zd9fwro1B6udH3WdfQoHQkH3/jDq9KrulxeGKHpX/LG9wwtbFPaqN3s
QsuzNI3WeavRK9qJv/x9XQk57HqkdLg1pKdc6AfIoaDcOgGexfQV1z6EUmsk9wkt
4UwDqIH6h3gayP1uvpuHCihaqdYV7PLnJ4kxB9+n1AEXqZB7tLEJZHrVUQMcFABY
IPsfYti8ewP7ESPB3nD0KmROHzybN9hjf938bV3xjsGkmemhhKNIy6RrFAOLqpIY
IeIOY/iaGWOBWy2eHW7JkY7wiv97s9SrWzI3S/CsSHa2XajuYW9vJfUjXWC5nIFf
RGWD/GRPrmCQRVyxEkGQB+kCRiHGyHmo1fS4D5VD2WeWBblfduyjsp4P2ncBv09X
lB5qwsxke0SV6us3VaOrzwuyCPFttGYrcDPJxmXQ1vh+bsJ3YhCGar1lWEO6fgWz
4taiUSugMNDifR919CJ7uw3qrVicOgQGSfhAbsi68IPWAgwjYy//9NbsX538RpH1
RbR+SWueylcxD1REKPXDd6G/dDQ5PkIN/IP1yigRqn6Z9DRld5r9AMjzbqtf4ouj
Y0rSexenqpkoRkJ2XC7cvWVYL1/NdxJRX2rM/tRY+86jcd2hLOpdb4j6cyWi5Efx
8jqltpR9T8RpB7DxEYO7kAqqdJoWVMpME21AX2YM4xBn5O6+2zTKE2GARXrjzD6l
t6YTZBPhbcm3fm2pHR+7/0a/I6dwB7S80ZPGAD5a6bA5nbdWxOQrgjqZ+D/LGYd4
x5YvT5+9gJbjpECs8nUZx+4lGemj8/8SqVCClu6+XvfT5SlBvRFfymurbSUdxf4s
ykaZy3D+T3i9bOiARiEPyrHNv5ElmGRT8CfDRcfEQaYyVsWU6F7qnuk+ZWf3JDYj
aX9YFSXTyPftg42lK/KYWpqAl/az4gB68R73N1SkHLvg+HOh//4XkgMljZiFn4gS
MwugzdsxM3PTNM5IQgkDO4UiMnzlSXn63y4cAKduCQfHDM/Dem2Eey4MT2S6L3vm
i59XinrtRWV/ry5kNfHoYZBtLIjS61RsQYt4PO6mkYAdRmWB1iqBuw//oBfsXrEC
p7Phs68cck2oyJuzVXeb1SmgTYV4jYnN/vt54w2jRAlzxn4BuMGmHBQhZeZrMlej
r0jV4p2C+95ozU5XZ+sbB7GhGkEtf4saMUbgqYwHVpnBlkKn0jSWrCpfFKjNx0jB
dDt/nCVeDZ1PhYgrL+0oGvmk/BTZP3TWyh29B5shSpnU5I7+kACr3PXs6UtTjhfd
hqnUiA5SgEDgZMEvr0qXDpjVuuim3OEKab+xoqCAJ9fxb8QAUkGXKX++Y564vbbq
f/nd9FnPiCXwrSVztM0Qn9l3tMjnjuoWHGq//URvaQyr1osMEMpw55yD9LOX1zhm
OIFJfoKyRey4HaHNnsCGZr5r8tAnVk43Cxy7FeeCy9eFvTuRsAAjMbTYl38fiE97
BEVPffHMcdsMfDhH9nm3J0VMXZQAVpo2vUFozuo7+/xwSpoxctlTqnIAl8ASZVFs
rtw5FOFYwFaQdWOq7Th0W9zQxYA7TWkfl/SbitUIFcRROfvOOin5PFGcZTVlhZkE
xCFZL1ekkQ2DcHZAcaySHt+QydxyEsHZ8cX/dZ0kpS0pKJtcWuNadmG66PqLd/LQ
Me8eDNuE3eTZNh5D2TtTvW9KGxNfc/DUs1Xc6UjWRnYOwJXqY2Yg4k9JxAgJtWyT
zjc7zK7sOlmGsLAa8P/rOaIS0Hh0rW/pJcoDUN4qHUcd/2b1fbYWpUeTvMP1uDfe
n0HaLNKtg9jViBcdflrm0kCedAr2nQ5jAqDvBQ3dddsyxsdV6/fxEoLVrURGmf8d
V+3LbDhsdi+IEdBs7DqYVz6kdzHDamITJYQuNa+VHDNns3O0j6/PJy1AIC/c7y41
5xbMPSfzGvnBb6JrsyAuQ3bpBtWmyWJx9w7vJ1ub8EQU7EPn7bzeV+bALQBVrU5t
BQvU6dJAH51blnjccVVxZCVFRoMiRzqn3aZ2AQGPxO9q8zG81hz9bVGU5Jvap0rc
Eb+LkQ9F6iD16Y8VWRP/pvxb3wc8HPikTulKQ2mdU5J+rwqPXQ1yx1pTFy54Z6Ov
L692vZh0yF9F76K0Ba6uKk8KpRGYIypYo8H8oYESi6cBfV4N8le9IfaPRBI06Ewc
ZoOgpzMMVVM+WxVg29y2WjsADYT8++S61zCmMKS1blJlzG87Sk4uoRnQQjMnucaX
vMYQWBSWC4mnX21q8ooRu3O9es319OxRGqQTCOOiEAfLgpYyXr47LI3dVbDOsbKy
Bu4z1QiOEaS0hrNJgY5NtnodJzKqEeFDQua3u0O+H5dH/wYVWx2tqViKCLH4WpWL
f4pN88JmjXVkb8foJDEJHMFOWLVbl8vL4q4GAOM9Y0/dPLfFKh7hBBHf3IG7pXiW
8BvidN9pXR3g0zwkhJ5VxLFSgxDinZS+OyVZgV+y8g602dJliNOjz1KXnWJoctWx
AermTnDn7EL4UJ1WCf/lLrrRG53VVhHwF0AVLpaltah0l5Ivy071ZIX1VQUJEiPo
PIcrVwKAmC6rWXNKcrhErIQcyo4ITdLXfPD7uXgJqJ1TWultDIP3hzjTM+f6TnaQ
yaQ7V31n6/Duj6MNmOb/D1bFofjIxGrYeHP2WHpIpYhmpDkpuKTrhzHjkoz5XIyk
Y5Rl2NWDo9WyNmNfYcPQFtZWwFQS5vgfo0PgGzD4KmBSzkSu+Ls2j423qLbI1PS7
GPx9haSrS7z5gLKbrxoA418ctMCWcARM4pUjJpOpEqQjC0pc3N3a2pw72c4cORLS
N68n4AiO81BjgcWRb1XKo7MKGszltSzj2AqCwhe1KEGHeL0W2q3J4BYgt7kJakWo
eNikgdtNMzbhD0iyuGKRNGjosqm7IGe++5TZRFd1+QPoPqulAhJmt0TSJV0LJQMP
cdWwB8lLpJjoS8pyauyOpRL0AKVg7ghz2ZWtGbBv3MO8xxpOjMsU7eGsrOHx9RQC
yGwVjT5AZwqQyliUT9wamN3WfFwfTqSfil5fsA4HmdtIc+Cc7w3rp47hQcl8JTXe
wHUx8NCQ/1vds3B6lzEi0yev08Xk02dAzGN+Dg8UnaWMq2sQ+Ns2uNEWAD898GRL
y3np+LAQrSMUMKFpJ23+ZOa+4uVLe5vhF8om9YKYYRVQiW0K6t/kjj1j4GK/zp+/
ykmjjpCrRCFQOCTGVin/VQHViBM8ABt3KngzvU8WvVWiJ37r6FocRuU3ZSEKgaKS
hNhyZeruuzSwOgGJaElD6GWJHI1klSn/YFtmSxAMk2iFGFMclL76YXxIr5zLBcNK
ZLpP8D6mx/Ed32N6YMb7I/SzSSi8lpUL+WPBYwp5yqiT1tj0cYY3jXCeYmCysrV6
mjbhNPIuaoYTnpcmJiGt4iTsu/DKGn3PZaKgCsRI0HwS1H1ynkpFzjR14wm5IbHS
1Q13xqWq9AH74UGLjwe2rgdxO3fwRrKzOCiJTFv76DUJeD8HjAWiXVm3lpcEOZnI
HbU6tNgfoUAqgqOWfUIbMXlAewPdyqHqJnS/xXRGOTLUH4/1NRHdv6NihHToSO8Z
JRR7uOI+G+uHxzPzpijNrqYtOZQaIm2Ipwm4SBLAsXZUGF3TscufhywSc53LqmKC
mYhet6N6LtjjGqKXKTQjpa/7ooKIcBLC/URcI2MweZDc5G2PvXWO+Ky9ghLjn0Br
jZiva0My7aige8Qnk1HaNKSbiCJmDUKLcT3cMXYYX0EHawVLTFHylzQ9fmRCQ8Et
ONPiFUZc0o7ITSiQhq8eoYV7WaZdEa8vzArIZ66MNN5O/Tq9WOwHzfx7WY6sbo4/
DcQpunx5OBDwm03lNPXepSSr1H3EQ6JtCqjkIDrPEYsq4MzsLOqupQ06JeY/6ynl
dhNyZFa5AEvITKwOUQrUoDlrIC3ekGcpW8Xt1i6OJtSwP7bT9DLzi1qlQkxgaPox
rHC24j9LjSw/v+3CpplpxSAB4t08IhyP/qEMPlPoIpRLbsEZLH16h/nefPk1L6Cu
WdnUGnOESaaw/pURIvI2N9UjcsQ09I3j3nIZndJZb0OVegDBYC565hx73xDivJG3
Q4lS1sKXJ0E23ZfBQUd1oZ2bl/aYaZOwhNRnWcfAeEs9YE22eQ4kDnKSN3f4Nhmq
32MoiuURJ37EIy3agA01JJ86upgNeyLC8vPluMTcskg7sRaMv3LnwmV/z+BYEysp
0ruZhoYftBOlAh+t+AZAecr/A4SEdbX/0d+MpP2YbB4Kt7+ni4zRSiNagPlm5vQJ
sMz1JSp+NjqLuDelkkrBWcqMr6zp4f4QBhubquiJ3ZnAdtqICT8KZW9hzxPNvWJJ
ko/WJnVHTzczUtDMaE0uR+vpznMgAttL8oOYdMMN0OqlWNnCSCgjwJfJgmbY5Lcx
IGEp6mizCUube/H9KKy0OVH170NoeUgQxICdiwoANPAgNyawhkLYy24oM/qgIhtv
eigduaynmdew7a7vqi8kaQx8pU7Zzw3I0J3jAEBAAO9qKdVWcpBGned+8HHws/FN
dpadcbV/4O6T1+E64fjeWD/NvpWXZOm9545e5eSuBYcmEyFZuRHltbh10dNAn8No
MfDq/OrTCfXKKck0P/16G+y//PXFow1V/sEr4PrMP7ZFwUXGj/RL5DtFIVI8F8Wu
boJv5GftMLLofh2KicDR0w6+NODMKbsBkzFiCB8kMfCAaCoSOXBnDi5Nhv6R0Waa
KlyIt9W2Ar7PZShCiUfQgimp+gbd68eGLM5KXqTx8vxby+7xPnTC25yOFBOrv9J3
ZPf2egmcggTDpkG+pOhWma183UuMzp2qzJ1Nnh3IGCHgUWkdfDDkrhvnDKxquLSb
T8oCiwYaGChhS//hjGaoTLZvRLEAq3Dr9QxH7sNsa8E1D9kazgWEZXNwSJMvELxD
IKKByEZUFhwtMKuTnIOwTv4kCP8iCX1h7+kNLtWRSeNXr2rYdsBvMCQczSQa+yBz
14+3P4sX4a9vnO9WynuRlSMHY0nn8/3Lij2xAd/VgE2vCeN1oaI1fAQxcKsiummw
HmGotGlEekleh3KhQl5RBwkqmcVWUWEtYIAmS+cnIKoclzP0EWFIm5ljbaZASw7v
lzRplTLzMuAl9KvzAOLfSpHH70oL4jXq38hOuImVNNniadrzdQc7Uq9dckIrmjoT
UVCn2XUUCm+38Viw4hNsRIlJsXRWyfoLo30hsz5Mb0dEmiQOKAS5MeEmbNBkfPus
GCpDyWSnSzLiNeaX6lk+tDKkmUGGPVoQD/fl2LFnNtR5SfVuMy57ZQXRFevCndya
Ypfg1zmDos5coK1stkc7qNtsnSwyRUojOlM9VIf1ssrYecWkfCFwGngHhJmpja2c
UQ9BW/7h9d75yhQgtqmYd45NJ2GJy40a8nGSX6osdbJK/LzPQcs9D1kfZrh8+l8z
6fYUV/ci0VodRi37d0KRlaEzduKegPLk/Cdgmb1tVEsbxYfrVU0nrc+CqOpWN6kV
VIDcnL7u51mi60kVf5uKxLgV10VMAdZxH4OYWYJr16IO3ToSA8/6h+7EfGqsr+qa
ncufmwesBYUZINIlisZDeH1JvFU7gOBPJMSFpMY4HsIq5sDBAE1Eaa3jp+G5WnRS
6gF/+T7NfsCEKxH3MqHq3HKkknzLa3+M1oogEiqLKnzJz+Z3WegxyT6KjAh5+2hR
Gr0n5w1Y5UMX68MoTXk3piA8ZZSWPK0e/9oB3L9wXQP8ZAoq41ldgVyec16OsRSw
7TaeM3dZrO5eXcmIX4RcKu5uX4E2eWGkoNi/mDmM0R76MflRaPWml7ln95JSCX8P
KvQGGPT7MA0+kVnDohk1myKoQ5/LOdsMM1EZ75aA3k6Au9LaXntcoDzM7HOpES3b
Anvry8DI1Q9bMO8twcDEf9Y3B8kD03Gl9+gU2q4kJYfW0y8Z3cR98KOM9nIZ344S
XiC2oPnLzMgZoIYxGCaFqnGvKuUSuEzw/JKdLqFEZzYqSYQ9iRYXRTW7t2MwDsQx
LJuhAewuV7gd97wj6y5QXAexw43JScEKEcCWwh8i3DnwyB5OWB1eblyp5GwR6Vb5
2ja5/VeElCOoFsVMerbfoLQvvqAqpLJJIayZbQ/6S/xxxMXaMBHXg90qiPxw3NVc
1KIbMRepu6262+b8uQmw3KftZG4Q0sWOOS6y4QU5REP/Uw9HW+nNAYMVPUCSW+b9
Xz3L9nzvDcDI6PMQJJp2StHzszNlBxxToWivnEx/j1vVUKSsyx8QAA+MV+6w4Z2/
UZ0hFTeKI8bc3XPOA6posLzBg0+xJv11E93CESiv5zm0wNPDliY2OCBnARA97jlE
yJwX73HSpink5d0txE1R0wq9XaLpkVJ6g2aq1TTdZ+wPRjeBxEbdkwBssuvzSQop
CmWBpWwth+SDVUyXNB15Uxpz2ytpeiFxLZP1Kv0ledlSC6yrOce8ThSyihYikx0S
q6N0wH9k7U/XEfUwaViqsmhgoPwc9Zs/BnwJocqW+JINMyreDOBJx5kbDpFHXSmY
7nBNVHY/1UWHd2oQ7yHz7/WvgVdx1QFq6HN1FSIDkizQfJ8hLlU92HWoVb5ExaXV
U7eZMpT02MAosFa7GGS6KWgK5NgAUmMu91kQ6k1Ep1++WzM/gTSPoxqMS4skIcSi
guOtbR06LQ/eSplyJtZh2aTrW+BuCgUxkcCGM8puGnjEl5bysvHQ0fK6s1KOBY7s
ELWzFAFhsB4Qsy5/i+5rrtDvZsl00Wlp6as2y/Lt9kuErNVkZqBWgI6QcnLxXdRe
wpBKLZQ4rP5zeq7TUYAZ0nI77AU4ryqaOCjVwjmSF4LDX9z66Va0iB/T1zUwXDum
Dplgj9+qe84iQwVIsmGQ60RAwqjcMnkbGfBGR7LaGwxNJcdg9K7GnNVfhbJko0U/
NWK4WWIF5TP7Q786TTs8oM22O2iTsE9rLl3zLNxrO6tl5hHNe2zwvDnVE9zPTkiQ
lMnR28CArrWmVYsOSW68pP8nyi7/Gt3siANMfqx/VcpMJtBOg5duDcTOURQMgZpv
9yPt2OpeGvIYI/7g/XGdklSewi0H0amY+IE+UyXOTC2tBNcUFqZi1rss5y4PX3SE
16P6+jVKYJXfMu5nRYbtw8dWkK7V56coxqTa9RoGLDQ0R+i8OtZYUrqaGMunT1pK
3ny0+805x4w3K0XJMBxNvMs2ARkaGjrb3z35D6I02CglmkGwD7PAlmIK9GcJzeby
ye25edxetczsIuZuKCPA13DTpBDSiD3Cy2abenBLtvJh/QHyabWhxjwrtcNSqQ/o
4i7Sn2B1HlqlOcfpk8SfHZ+SBsZlhC2BMNI/a0tYCp945nfqjO4Xv0tIRw82lP+n
njs37vLtiAzP1u5Mo6cQzGvKHADxDWtaXo5iUok9GTT/WLqPHkSfGxLrBB9FXZms
0hycfHb219BsEQCV8eaX+1oOkNQRKntVKXNUkfx2CaeeVn8BTp5i88mNLQ7g5jQ2
/b40tZWUfvldzRe9I/kk/Re+gCq/KyXmiey5hRj3qy5YiIPWWCVW0YT2j/IlK546
hVo6MnuZdVYbKeTj3DrijAs+IiUrWiDp8x2ydfFi7rHTG1Ryy4xCg2xeqmQG1zmc
czNpsk6KrEKTA0DSP9WHIW6zd/5rN2JC0t750GYi0WI/EBmj/cDGOxUUlfRRHv96
WDDglJD4m65lcj7B9KPIYFjj5k6chPTPOJll3qaI6lXVsxokREY3IClfkcsMft7C
ZDEDhgp713A6zvCcq8WYTMLIGwwuS8wgHFwIrl0xgAMKjXH7tvBgd0RTQXv1QxSp
Rnpd3Al+7uSEW36e8N01TvHXIRwPegNgC6oUYLH4VZ4/15UFKh/L5fa3G5clod1J
PjXPbI3czQ3mgDsdjpFAMrgnWNHenbidMa2Y9AzIPIxNzOCJb0WuoAe0Sm05gtLd
bocgGxDwvhTh8uZRaSuFDHH+4k8tGdlUboE4enM5JpVhFPqbkKedmfHi4AcYIVaL
AvQpct760hdWf5bYBof5auB5rmDrVirXxeYyynPHddgfjc63+XVeadCy9nQWMBaF
ViugQFhYbtLvdHB6AAcgxkWn9GEooJCyL+EN7UJngnwkWvdNU+foqkoYRkpYnI8u
yIgqHWzbwWfWkHvubT98mzJgElg23SMBqRVQMm1YV74zrV9CBLdMf84pMr8UvzQc
0Dp4am+Z5QJjlL6lZhXf7QR/36SRJmn2TNBIwl1bdnzNMlgxL2obQdoS3A3hBxYi
OapiAudT9dFJz1uEgwG2HBIZviSyej5C2MtBq6m/GIg4euXp4Cq3bQlK1wYZ902X
eBXNwNcv4cc7qf2hRGpgsBFjmTHQsUCYxSh00UsYtFwA/Nu+S5useUB7VKVSwZg0
ZUh9nmYMnbthUQQawL0hwPZRLplvQjNnmEf1rnHd+W03ZWqG7V0ztQDXW49My89D
TFvUJFeKa5KQiGVf1NZwGtFi20Y7iIcmFR0x0zcYv+wm+PDxVmMW/sYJaZDh1YV8
znjxp8XeqNJWzn9qNqcKTGRTHf38Eu9bQqkjxdpPgW5mQgZz/tjxQn/rHEY+iIxe
QQHyV9lwDW3HMoYpPVjPnSH/i2QnR2OLmobOV0I2JaeRjr2dMVNpzEJqDwh9iT/N
7eZuGpeu3LdSaFcV81IvjMfMdxcNjbsOi7qqJMJAI/C18HnEJFRo6SsH8yeWKdfU
JCOD/jzGqEqjhEFA+ejy4EHKolmyys8+3meQDs2SXuUTizH2UId1OhGwY+TLsrHs
SlpWNcq3sy1YSKnhR2MG6u7/6RcEnbEv8p3moL+dENygTajXTXg7j2awf0LKJeG1
W1FsRyScTNAr2dUDmOWpke1nYeBhGhh442oza/Lnq86m3222CRZPExxEo/PpY50b
xwbKiRLDV1lMSaZDrgqk4PitQ/rOXpBDvGNZATzgf3s5TQ07XfPtjv5wVMuEWaWX
PaRV57LsCvCoMpRO9MGaxZJSbuHmu//b5dx9iMHXNUfWSEl3uMsQ9ym4YkLvKuXl
PunUPRwOXQgwtpNJU3tcrbmRf6kQAHniIL2MUMWbekSzZncQ7i0+Ltmff57WWnGB
kgtB9e2JZBzKn+ieUmAXKup+TbE2oZmszkfxk4qlPRLxRc7qvb9wBfEnwv9FFMb2
59FcirGQSZPF+ErTwAvLqG+vzYckOK4KuVw8hLjgzMz3NV4FheGIg/vwFno+HBrE
3SPoJ6ROtzzrJwkwUQ+NsSQ1c/i+aPor1x/L/RtzTtf7N9KdNRTDJJya1d1AFJkg
c2EkVez8/z/fSPiXKEo3w9nr6VPpkOZH8kvubIrE30mWu2+UWRrr3oIvVTJhsEXV
RFj+CDwYloJ/zRE6D6JTa6vBiNl1W9p8cO0dkY00+/1ntEhWtb6pPo33lCh6SXl4
v1b953wvSZ1CMJfdPNzqFIft3covdXzwWxQo6qPMaLWPvmdeBJXe4cTSbJwzzsHs
iYZ9PqamrrGWbl04nR4Nwz065X54Y3KGJbhh2QwcCfa01ZkapNtKoijVqJNpqxLY
A3RQN723kogdZSzjC3kQM+XsxN6jTHjPeh7Z8sMAPMziwMoqgfghXUINTKaaF54M
1PUWO1KzwHFGrPUP7KpDpgbrl9Wbj1yDrEvJWRdZzK6CUMEYtNR49c0ZhzTpjT1B
pHccLpCp2oAkfN6ETz/frbPoN66hNGLKCC2lxchnqZsqwYxO5+kJayi/FuR/cdyF
InY+fDPslXfthpkJEsbRfMxKnexhiWwDSrC+AX2b4d+tE4UmZZKHdfVwhCfmmUyO
JuG+5g5xGwZnvVge54AfzK4P/U9K/NRaIhNVSVrcYXoxTGpKirOrq7jjYHt/EKPP
Is6XbKCNljgvOV7IH7XAwODqZLAk20H6GGUeDvzIM6lhWGAbwiPTf0qtENXtKORb
bEH/CErBptvyV27e64SyTFACVQLcMVNo4IP0qpYzaHMjKrKKDRw8odyKhhZMOQL2
OdvVqKi3GdRW/sWSRhEDvgYicI1Vla/wIoA0mJR95VlmiCQz7TQR6QFNcpARUWju
vWLMI7rOptM3jrRG2ddloH3dfAaalsBHa0JXcef8WC9XYvy2pRhVj728JX4vyoES
CeM5bj0OvPwTVcxFHTOSK5S8A23xS/bwD0kLfgxUWi021eLYGvU3aLk0ZXEN5VCt
xw25+pOUQL2XGCxqGqSlpHVHkY1sAdVakhDQdcPBmP6v6O4o1nyjD1iSOFiFVisd
X2dZhKWGES31hRPEtLbrNFIreVdec8r8/Xkbo+j15R/2SeAigGBd8Tt6JWDEiP2V
CVZz4MBQWavo6xTcYcKY+UOrJOejhe/FvcODqGOB9u1OeULM+kVmKCbxohF+56IL
ZD47sFzaCKRvjH7X1yAv010WZbnTewvk/nj67QdpABF/t4yTMpUfZz4q4He4SI0h
ZrQqdR1phxzAwWhw6F3wCOYJdZTGG2adeRg6jBMWyvb52ofqv5QILuXovkgclS0N
F98qokOqc3xyhFr5uSrHZ39RP7zpFWIRMgO4w3fF4awT966GDHkIdoWNWpsUrbnD
1fo7cBS4jVlNOElK3vnFBBrkXadBBS3tuAmkiwcqibwj4DKN4obYrSpNIVUPnnpR
OWMZtTivGqgA17ic2eBdWZ9aOi+TBwD8GNgX7d03OPWIIb64OjR6f9nH+XHRrEKv
qMo18G/zaHcDeb53eSFxbMMjFko5MjQ8Qfi22aYrrfeIfXuNelNAtr6/m/bk4E+E
l3Kn/3D05NxOMMMq/RI6kZ2wbKXkLwE224AQxoboXEW+bZ+JMX6kIMkexOJO6zmA
jeP6aV9bR89j+5cvdz3Mkx3Tq/cWG51w7hxcRjMRrEBSq3AS8fTjyt/+QU/ME1jA
Dnwm3zgzX07RMIFkldSJ58qzBbMhkG9GQM9BIp9ZEDTzIoGDmhxxIhwRwP99BWhX
OTI/OnaWtPMVZqSgJ2hVEFV9A5tcz+P/2ua2msQxMswA3ZE+JoOZBYE1MWy9THYo
rt5536YwJfHg/sI9abEaJMgtRCZyibjgNk23JbiLSZfi/xdy/ipIcoyoUntCIMvr
2vmQgvNonmGLDEYmvcN3Z8ktNqm038BIhogjrVmQRgp5wGR/zOy+K/iXJtfSDJ6z
hpVDCShXarON4qqKE7fg4H6xRSEEkbURnYYb3wCNQxy7lHUJ+gGQ3o7Oo78vRKPR
Wh/czdLkj3u7IgDsQlysxkZ+YMbub2bgRaFepVkEOxQZmFVSUklnZ4yzJs5rPJ6Z
9e/4IUQHkptD6E7lvYl2ZkD2M4BhxP9b+TUH+PJgn0DgksbKM/wye4LCAfORH1Fl
AWuoKv1uQhcBVJNfbq5nksq7U7jUKyTI02YtOuD4uJH4teJWrpNxbrZkbLYHRqTT
moaze2qb+6+Y7DsS+wPp1XqAgKSc9gRLacsAxehWKDem9XMPtKpKUZRZ3gMVU6dD
7r1UdmLoGkYR7PINxD3K5soDPyOn7yeHUn+i5HTkdfVlF9IZ6VkVGs514Lmw6YzB
15+RQ2U5kl0GMR6Zjy0zwudnT8Dal5r2LP2Lr1V6AalbpLUleXtopkzjov1MUc8P
eduFNipol5eVqvr/dGxjSv5fl1j6pJEa/D+msN6PqjmXsshEnTkbJK5QFoX/Ay2j
fyNywazBlPHMU4Ym8P4d+QPrUBIcRJ2kHsCklpj9muQ9GDskHIewBG+YqnX+MkFS
vw1rDF4qI0LTFv+Svxck/3FzDvH/e8VY7RkirIisAg/5rKd5/LrpExHx4GvBqDWh
yGtMTiDXdDNa5fIxaRKoUp0TgnatQDRnCn8ncqWmcCq6FCb3HUTnGaxkJxKybsVL
3nAfHN6GZJ3F0QLULkuBH2p9kFZma7HxI+dBR20Q8JsoEl+hjFewN2bUVyo4RBWi
Ze7aqjcPxjJeozRRfczG8Q+8fNFmq8EZV1COIw57VaU58ifolf+8bOJDoySlGOAY
ZUM7aBiKr8PPg/kmcTRBlLJw7Q93HlfB9l47H2OWG+npz6JHRbGVoIJkhWuLfZG1
hOOSmTOJDKC7wHp83NW1uWCLy/qm3wxKSMLkgTKQE6EHrskwRQLBgcvUMXJoI6Hq
vwtn/rqnMuFw535DV+Iw4qhtuXsZ6fOvkbZe3wSzCpb8ZsbIqVUtBKBzp01AIDay
pIy9AbTTIeWGhoPgCTbqWP4Svhpdv/VB/8cpy4lSQ0s+sRKYuipRbUOnuCLx0cUA
l34JpIUgeTFTsU1X75AKZFI1X8gI5G6BQcRj+foT1AX92hcLp88jU2xEuScE1BIJ
qQ8q5KmVPo09pPWkwHtRpL2/J1nbBKgwhLaGYpRdtpNWvjUnPs7GAZw3GuaAZ3sU
gQtb1bRb8XUPiv3oUHxHwrAlUXYOzidCyBkxR63DiZFMBPb7jlyWlH2lO3QlOJJU
y3auevL2xD7B13bJkGt8/HnhzOWGIZiQ8dccckMzlhsJpIFLMlQlmk1EQTNdwuaS
jZI+A7Oiukabaz/lZgj80Zlg4k4MVjMtSvBqSBALxo+ys1TxQKufj8H8WuAgadSZ
0eUb3exfBWYOd6vHAT5hRhpJ1H4EX+HMKqcv1+aEe0o0eU0CCa2X0dWGoqvrmDKM
GWRlSDyWmb7omTlcnl0ud3++nEu1TAJYtw/7vtd1wmypp6VHh3TNqHfjBlN3XNX5
Oz0kxxDPO3aevSomG4QCJaDJ6WSozUbprW+8WMM+yMHs/xSaptw/I/q83Rtl/1t5
WGOT+bqtH9KgJNq+QMIRg11aVMdq2MdMeEI9iUzvCaXOVcG1eKdJgjQDw24cl9Wa
vvAs7gAo/Mtru9kNNJ3E3Et/sZVbPAeNoT0eQMigIDHeSTxKGAIckGIIA7SweXBl
MvP4DKVrv1phBBLDT5fQDzGJNz0eRqahgq4DsgMI6QBA6FVIYoZZcq0CxAmYZqtb
WISeFeuY6nhozQOTQTDeYgTS+SveEnB9p6CHNkUSDjo0cSbREGxtaxKN+uUeMQY4
7KvdOQMVb8MuvuFvjj9uKKfRHpOUnhJwUZcwPleW17IgKasWRbGOf4r4VQ0smUAp
qmNq8WbifoHZmOgcPTy7vEhjygKPckHUKX9mtfZm55fCerZ6ONe87w6Htq1RqssO
CvmyPPDYcLLIY7TU8ZRUqaKed1UZ92HRzGyCuLIJl84UeMv0d7ZVrvJVZpFqHMix
Lf1V+yerLZt6PmArEWV50z6oBH4f9tps9PoUxd8MGhqMfveWrUMj7u39E8wSulQ3
vQf+M4Z+X/ZTeCiLznj4dd6oLWngHggIW8QcBd5auBLz5789PFna4ZeBHTK10ilz
1WVi8/puf1IjHRPoQ1pzNvSjDi3GqnMm3aW+PhtANJ9ubY7iGqLvaFkyulq3NaDw
C9xbk9+GHJuAwmBQl8zgKhi3/d+YZdfV+GZN1L0sLeMLVVV48lpbhhVIner8aR66
EKutsijBymfSG9/AN2d/YLafrrthECskHZimNTEPoFDdWaTkIj/feonsjL5yBOr8
rJ5YAXbZni5ttcR4BUCqcn7mAJXNoAjwSLtzh+YI5zQ=
`pragma protect end_protected
