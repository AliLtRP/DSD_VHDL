// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:17 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
UBkU34LHjIeUX2/AtnKSZcBzfklC+ltBd1T8t7/wTxh9Et6f1ayQ+FOGGvSpSJW1
AtXlIIhhRqj3tIgGEanaXIT4vq+82cWNU/SThhBce0V7OkfOiB7tfb8z74yJiUVN
5pLQxRJ0rJbAc7DzUbB63H7iqtSPkSVGL3ATmXnU6rk=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 30208)
aVe6PltRA31d2qE8+MmsfEls4AsaxondFkaJByLFfpIo7pqRViHu2MOhX8X54YJh
7tbI+0OBZN/+oVXKer5WTKScgRQ1mi3CFjktJe8ICvn+BrWq6WOiI6VVDp2f+qVS
GdiYqUIO1IppREs2t7pyXecrdWEXg+ENa6uJrMPVHF/2/70zFf6dFs5YNeXSbPVj
JqQJ4U/wAgVb1QdTwSQj7fmgaxFQQCQp0DmB+UOQJoouK9KiX4int69XF6grVUoO
cdLbgSlJKJhQrXnKEzpAYgfzhTAJEXJWLEWYkR54oOh1oeUEiQM9CcieiuX4XUcN
SdwNeRu7zUCEvK3mJvfgO9XJ98FKJHM3n9awQwFryQ8S22Nt2umggtBvJZ+9wqrP
3NQ1H9nta0ZLIlvTFgGSeSLs6hDvaW96cnYLkDJha9xe7gFyw7CyzkT1QyPFD4WK
0n5Iri60caaZFms+yeCOA49rMDvyZA8CE1HGG88jcPImBFxJGUXYTxFMauaZ9b0M
3iBoRKMSHZViFd92jc2kMUX4UJrHLUHidIgwJp3gtVHGbkG37+SunWV5f528aANz
pJNLrLpNjzhcy38rlbll/OK8zhllcmNmVa/ZBVcQQpa3ojMMv13snTiHjEWxW0IW
RMedtxnKWUGzNfcxdPOZ6jlsSy/SdygdlK3rDkhrNJPQykX+iexJ+POne5zp/dNo
+XMt4RFf36Pd1SC0NJ2rAMcr8UNGe9G2hu3BZGKWXU7bQxFhpvlUuSX0JsWRcOt7
ukSIy4L2aiWQBkiqGTVwJ88oTfm9FXWKD9zYYrP1jJQ+0pw5/85mLKVuAdMlLWbN
0uUmjCrZfXQaNpjjT3r4jzBilBC0Zidnff/vTsOFfZzKKndVcZXFJVVfG5lPzIiE
1KcF8nSOtzlMs8hJocF9OwABbkNw/3VyvyHKbpRQ8PfGbf1A4JR1Z9Pk0RoYypPy
075NLV2LDVDEHa3ZlRjuRAm95mPhLv6T3mo4ctFUAMs8AalARvo+mALoueNfT4ZZ
iIGiJQlX6eN8pWMQeXNdlRaQWyd6OkfiDMQGmu1Ai7qXL8JjejG97N2n7Yk6qrAU
GLWter2wlB3BFtByTaoAezqwdeIzuIbXpH25ZSydE+p5GyqxRyEt+cK3GOMXkyBd
nhFhPiQ1LwtDXxBk5V5leZqFIldmXF+zc1Zulozy//beoE929h8jJdiHl64xKTkM
ZQjKCLS145YqGvT/FeSPfJTVrQ8Fieseab25pWo4D1GfREjeYFXS8SpeWIUa09Mm
hLB9MxP0qV+eUmb+BXeQTmiSuHSvlyruMb3LpELKzKRRZ+taklATBk6Qf5/T327J
eUQe6qHUe+veb2YNsDZclC7LOihew1f4AjwlwccZYWMjx2WubLA1wy4kuGOPmGgN
kV4SfdKFsHiAYI0RHs8M5FqN2BiXK8fLsZgY2bKnH6HRHCT7JMuVFEfq+KTlfhIG
cF/w99gAy/X6SZS5fPxhGsAaEEBl5LR82F4IKbxIbvKZB0wjyGBY3eXRjYX2ZZPT
WU43cS7+MDpzx/BiTClkXFomu1EaFUOJE/CLyE0DZPXLneXI8JdfDUIA+vc/VVLA
R4j91j7o+PHqwgbOuQOcDeMmZir5o4EmWhj7rmuGBO4JX45wXzGGHDEgcJK/pCx+
00756WIhoeSUttbJ9qUpfRmAicFa4vnkbPu4lvwkh1yVZNUx7DxHOJHHzcpTeDXs
iOD48sWHuhBvVklcwTSS6JgfQM8wiEBN55/UlGf0TJnIiET/cd6+BWdWSY0uoTk9
Dju1Dn1i6mQC5wH0p7+Jf4TfnA2r4ohFsN9myVX5G1/+VPNacZojTM66vcu5r5Ua
Hr/srEgKJc/kv/nQ99/CwLLZ23DOcvCcyUE/Z30UjNhePIFQVLewiLTaw3Dvwugk
tfhE9S2VFsFRAuNCo28d3FFzqyIe2j6nY3sIt3taBev51n7hJZqm3Y/pEykNDOaR
EQK3Hjet14+dAAZUmA6YByMicMu9eDp6sQFk1mHH4WCx0s4WA1Acu+fMG4U9DMZ4
EhOFAPtkknwfCdDVFpZVaNnjCgm/YZvUNVrXEWg38V3qjPRKqVffQsicuVfT4/eS
h1OmaWfCWlt6wGrBUf9OL5vz265aCmD/omDjhV+qM+GYQAggv4ONsvjYNZM66Wjj
RawTNXuF6nCOTdmqFKVDP/nAjY/RbTfnE4EI/L4/CQYHxgKd4wiMKeGI9YxG2khV
rekBMLcPuQsAWW5QpquFHLKI0pThlDSQC5WgfXksFaPv5ES3hVdwF1Seh9l6bfG/
TH2tR3c8WS87RIpAp5dDBybRNU6Rb31A4pnYjLHH5srlBgBMLp8a9/0bKUi2OvMo
P0LScYwZ+DmF/NjieY2N96bN5ePpCRI/oxVHGSIJof+0M1j9im5gvTImKs8eIB+T
XQUcs6C0W8RC2TR2SbvP7IvfSZeA6ro69Y+LfbeOCgkwLqGgtWfmNRPObp9ov73v
ltLQc3jhi88U46rH2eP8addlWN6XiiZ+E9MoORXGz/qSeQ7EEtWy4rgfk71bAk+z
MqmD1Gdex9e2Gi/a2Tzbui/Fyjul99zjykuhtIwKAFkodXR5hKIk3xJtPX2Y+4Wl
QC7EMvQMlHP0o0CODBilZLBDol8YC1nh5AsGU6DmLG6LZaRjjHagxgha5r7kAkvt
5lZi0nFJBiTFI3GTvoDlT/cZ2A1vQQRIN0qDO5lgxop5Mz8wOcIpWCW8ZFJFzenM
MAiC3ZCNgVJBaZ16COYE7YNb7o7JUZo23lGvQsMkyDgO4A0PC4fJ59N+79r/vV1Z
1Xg7/ftuXW4RkhLYfoJSaAnX42DM5V/yaGnR6cUQnlt1fHdAiTEHZMVc1zivgtgZ
anBeOCNxD1WM1Eadvqz92voYrQ/+zaLcW1cJELB5uQUZW0iA0bIot/13qRvo2hAu
ra2DwEBrIdomkVE9vQqYc+nw41WLxVwbJ2a+FIu52xzIW4MwrL4CvJL2PeEFOhHW
5ZdNzJdae5hSK6rb8EOgpxOVbaXzEHUoCsKSiEo7GNDQnUDGKd1o1sWjBtOIQns4
23X8OtjDebYgA7h6WmKB9IO9pm4Yb6NZMYLjojLNZmlCvMSUhOrRmLXUUgS1gXP2
cY5WaEadw+Z2tdrrVc6ucr/hiPJ8NvSTyG/Ij4J108suPJJ5pgq/dmPeIDL3Sxi5
zuNbB58+5uVIkErDHhyhRbNEW3DIyJXpll+qo8RO5vzN9a/Lld5J7a6tnxfz+cmM
XIkVQQ4Yytp41dU30RKNUQ0RZaJhhW/qqlLzpYe68i40nga52h1UxoP1himErFxF
3xKL6PDdtNT2XkSdt1EusKL2hOC1fQkQAwV5yL2bpTc4zma1PhguSa1X/i4jdvc4
TwwgYnnKnu/xNYaNEvFSxR3yexqqeviELKLSezuZors9S3kUPL8jY860S/BBLTh7
QTkL+rwktGpGpOJswv8KqL+1x0orKg7bQlv3TORypFmF8EUyO5Qd33ewYItWWSFd
kB55+JGAFpxkiyhR3hkGTMd1iYlGoCmItPI3710qkrt3+6SLKhmLG1ZItM+1G/5N
icDtQfr1TuleWxoZ12K0WHBWd5Rstwkf1QGR5AOO4oyqEbjLmDJ+Kzg77auIviGo
Ewu+ftxiu8S7IUoch4fOCOU0RtAib9s61dyUrZLZWTwAjUZ4U3KF3zJZfd6v2aoZ
us+sovw+BJwhn882HGl2rYs0V7UJ2xfMtcZx+U+2v92rpwZZy7jGhSp+gNSFmv2K
MYfpR7rG8hXFWGnbog1DV4GA73wxZ5eYH0dWDYk5/xdTK2M2j0y8dnDVebGMe5N1
Jk0zUXQRvlyi6UpyMHC43OnSn1JyIxPvsVnZPij1uja8CQQptJspb8T8tNdHmgWz
dr9ISdPZuPkzT+XGOJ7b+0lNFVevK1E0vOfdOVsXYwxdNKgPABdfP2Nse5jOn3lg
cbcBY/YHc5vInoPphfXfwrOnjR8Wu1zNcSPFOGB89zqeRufEYkbafYFqRXkVd4uY
HRxLwwVbPNOPjoSOrEcAJLOWr6+ptuqfN1/k27MneBV9Ene/5O6ztIxRxtLHvDr8
+HifauilByHOeD0hePC8aZ9dUnRLYZ/hCOzjAt10ij/bo65ELYy56HEerl42PnjJ
pPMH3W4QHjpbIQzO/LIuUgWzm/z6x0t232WM4vCZMUI/ckXPHmkvhFG/4UW7uH6t
vBaZH2sbyd3DyfGM1xA9rRzKss+TMGtVPiZs8icizvpywQHkhf9VZ+b8tjbw1dIK
gNfmfu+Ovgj8xyNlr68Fsc8skWzfbmcHsPUwJbQptvw/3jz0bSVCOTUzDBPFn43K
qGfJ8ZKbh2S0TwWmsz98YozKPYkzaFEz53hsTXrO4rMSfIUrSMYQHLoq8C6gagzT
W6eOWsq9xhMjAHsGbvIJG15iQMdDyyxDrdMNNk4GffmCLXmGandd2OX5Wzhd3jvw
rqpXfoyKfA7V88oA0E3Tw+hMo3czLX3IN4i3ARjvd7FmagG040XUaEzhk9jtat+e
J2BRLqOjOimjOYGT0J9A7itjKapUlIZCweM55RhcH20J0ZXN35Z8KCVTypuAaYRj
Jfp2Ti6OoafEXGbtZLPxuLbi7e/93UkP91ygWggiAVjIQIZPst36/VtAbn/CLRsm
IeCMUdDALV3q/dkqAguBe5TCEaHkaX1qviQUAwVntTybxGLLYUqUfnfyYEMkAlCz
V2W+5YUEalGf9paDzbjgXT+3xqaU7e0YgUr02czkKX6rn00w6i5vKqZyN9soS3TC
3lqB/BnYOFQX+Wc4g3CAtxG4xDFOBT0RlgeZqFgplkAZTXWAEZ2qALFpgC1D9+tQ
jIHyWBABUGxt201ptom/FEJ2bX8VD2p7bXwAPxv2Y6EOplB3Mx+14IalZPqou/Ri
n/e+jKAFx4ITAcgf6IF8m8B+mi5fXNHImigY9YWk77LpJ05N3xqOHKjUmhKpH72t
tMBHOw+FCR8odTNDmjTFzfUG1w2CajPZN6nMMz1YmKgyiB9t6ktNAmYC/iO+sO4u
FY5KtZqX2fur5/V3jsx8JOJtCrSicsZPHxpf7oWOVauniXF/7j/qRbIOaqULROL7
6jyblvnVNZ5ceLtNIc4kaaBqp6FA1bQ9tYA0I17nbPyeHozcHQ/JRmdD0tt1o55Z
hiXVZwNPelmDWexC3gqYtMxH2YTIK1YkOo4Vx7DIP0ajrydeEwiQvZUjikdoT6aN
kwVdvlFsV+UKEAgnxrlqYkNRwvG8YI4oyJa2656JqjHkDNKmpDOQLkyOxzHVrRLm
AuqNtJh5ElT/DhEXdlswdcTb7ebU2PhFx0IpWGKdyE7J3lpAnEbVdLWIc9sihBij
BW5eeivqSTz6dYumZGugL5XpCj1itH+Tc4FKui+FXLvmz07TY3hhGAfq0wDm6uID
kBWevoz7opss7qpsf7oqfZvmWLORGxqHuvJGJLJ8bn1pP7ogiSAFka5PxvjSjwk8
9/6NILr+EhSqhI6ZS0l/anBii7GgK3kOdZ5eaf43riFXBucz/tilvhum/2l+roX1
7JCinqaT6CI6fuZ18fRjNIUbPeFqIrXn52YjPWQQXTPto5YPTeVycIQ+W95/l+6D
/EMsNmt1nsclUMSp3ljD5sqkhgdaL3GrikVVGYURVRZbO3W8ZplFFZ1gpjnjmX/c
Yfpt+8CQj95uAekYP2P99LuLmLewMqWFgxdzH46iFfpXHW2nEJ+CXFQoDN8dRpyX
9wSPSuogNjsWr0JwsPIJQDQnBx5IXJxDr5fi5ybndsowxARlXtYuWMbG8yFrwK1A
TiMmf400p4LMXsQLOBsnJms7XQNZ7kSyX5AZeu9VCMCIVrYBNktfCWDiecog/jnr
90x5EHVQf6LJCNThzp3DsX/fvu5WPtZrBYzWmp7rqRrGe2pG1B5eM1RVs5MRsNgW
uA2fPw17lNXiXKzw4Hlyp5k0JSkKUPxgX6z5hqt+swvbEkfSuoGnIiv8FSSgjt5B
xohGZcrhvIq0Ub9P+WD+qjwn4UKESwIzwFCkiE73Sgyw10rwzWAPVbptybQ5qPV5
kDH1ECBkhNSLPtpM44/sg67GW37Kmxb66YlV+/wxsmhzMYbV0eQyvgOSpeKyaFxm
nbBd7oOYmiCfh62UO9KxNgDyZheb3FE3T19VaUiIq8b6bsQ2fj8XBM11OF93nlZh
KZnQayRcw+NPnUTSgbisV5npty5KWlanPKvwXKJQmXdOkT35NNWZEA0/YjKd1v99
lU4K6y1goJNEsU5vMFD4NO6kd9T9bhcGCSbJipPMX8l2gRbTqOJHZv2/Dpioklhw
D+TUZ3c58ll36FPdG6wnuEfb5nUUIxgFW65dLS/yN5xHTNnEbEhQOLB8Sqrb9niB
irVci8jW+y6o2ohqn3ZWvG4QPMtYPoeDXWPrrFsyVHf/tpVk7cARwTYCLC5aMMky
Dk3+gdGGliYIqWELi1+4jYEcJFjuBeadYhVoTtyeVQNasewFtqEDb6m86eMkHepB
jpbF5ncVkGISMWGpbzLSN3Wb2xuu0qEyql1cRCee9g0xjeZNdWTYiZ6aO87zIp2K
Zc1esJ8j7xz1Tpno1od7hB0pH8Ytt50ZxU9b8WeEYow9n+qUnTVIWObu0zofIpTv
LYvUXuc/hjj8m71KmHXFsN+kmN8yysKCluL86FwcOqhPOLxTPxwxtW2hMi1E2ZK0
94RWu7hFREx1TsbmU+OEp7k7NJAFBZi2J4AxFi5JGuOZ4EJtD94WZQV0BvrEFiSl
rlR1dv22YM+5GxDphJ1VYNAJs2AY55zn/YAJhIr1W3+kGJl5m/pL92stv5N9iPxV
wlaQey95v0NSDariZBKzDym88RinsHjrQW/RZa826uKCGzWvU60y83E8GkaUg/XR
8febuBM85Mbr/IkNe2gzSz8SQzGrGcILdthJrKiFaEi6PuLZFb+rR8tRyXLzgANI
MXaHpeUrVG/ZhoJTmhTh3/mOm5hlGkS8H+B5w+2DfuCw3xWDXrSnG2O97t+pxx8a
BYoG/Ms5+A0PQA7tWWoiAWEvRVj1QVf9OEe2SPlGE+AqTrCA1Gajw91EYVLvnTJg
IzLpSDXepKzV/GgbHce3OtSa66AyRAI6iruEWBYlVKcbiDfVYhbTNp1pcUYjBgcH
ctLoO5+/ZqB67ptmYIqhfV8bAyfzYLF6HEgkiiN8KyKGINBOxSK8IdszrmyHfXHP
SyGucGQB1czX6A+mqlC7dIeRSeAa6B88S/iB48iD6uLIdw8IgVCEj0gb1s+dtxR7
vje+oQvCCmMjq2EeHFSKAHPwrRsBmsFqxQcP3h0hieiQrEPJo3TgYvY6mhpuYSPp
FxF8yLNsSbLgW1H0jXnjuU+dMoIMSFVKRTcc9QVUPajjcf1n6M4IawjHpX8pizDG
FobZi6Bvhpi9doSI/D7JexoUh2NIPGiUXFwsAojXuAJxxhAb0WqEOpW8jqmAJXIy
co0vaxqN6xWZsTwMqb14icsB1xw3ivwSVc542FDpQJ0Qzq7UrRoFc7eabDqZVMCs
qVPNADc/YfejWNbqng5HZelSm6ImduBtnfRhtF0yw2D9jQgAElvi/Z3RvsSGZSI2
FEH6DBZlnbcrWMqDWVrX1F+6d2mYf3VMFV5/57ucZ8ngYC6DlhT54l99hq/HNLs3
pBeNE4k+ASA6jnD/ctY0pI4xuIgVbn0OXavUWVSb63SxkHcymPH3eCYDmElzdMFS
UFNvaUcpGRsPDfPqMDiAb00GkjhsMAVFcJ7ZG7sE1+nTBKqJ51it0NwTp93vUsuE
UWt3HYqMttx3/soSro4Pmpg+yqOPQ3YY4fKvx0syxIxzSSxrgEIL2ErZkz+psAVH
WQFfPoitsNqbeF2IGSFVuyBielOHiHPvs8EXz/PKNIds//dndUSCjJ8t8YkLVir3
ySgFCaLS76niY8hrK9tltwEiSUegITHhQxpTtxXT/B3v3NBy5gNU5VTyMkAzKXhj
WmhJaBJVBtGDPSrWQvOIXxHMxatrWaMUkCkXWi45UdnM1a81jFXJdOcs+CmeKCxF
mY4P4VE4oqaWCoOZrpUhFaPffHKqXs/UrSD6U0dnXUabeSWe2OulMGWk+AG3o2C6
pwiuopMY9VCeVz4eyRGA6Ybt2PCktB2pSKDkkcC4nQzvPhLNaT314UR1m1gNcLmA
C72ogsEglDLrYPtLAyA30kI6aAn/KHbrDL/py+bKyAdjwJy2v5MvxWA21FpbAkec
kyHvcUCI4yo2e+bU3CBw+EGe2MwPXKTQrqQthB69DUVa0XQX3Ak4wJKLxNJzPCAg
HxY2O1UtczURaERzw7SdIeaB8eWuuwdjs9Rjrwq9iUL9tLAk3G496lnhYfNQhDMf
Gsn8WvaHPJPvemnRa1Hm65esDjbTuAT+o4iKIkf5Z6WwNWKmp70H3bv2qWCGcSbX
kbX2/EDmj5uQyKtD0yiPnZXP2NZL7s1KhHGplAdhaGCUgK3VOC8MwkXRXpS2McYA
D5nOUA5UH73ruKQtR4cfRUDfpPiTgSFEUXaEbUmBfJUM2RArZYLUn3L957284pYt
TKf0YdoEdtWA12V4AvhCiLfFbic03tJB70lzD1mOPlYR1DPxedJJw9j31cPrDB/+
hhE/5WPhi+25d85A34ICcDr3Ft520ThWBGM+4BJd80oiTW07RAlII4jPjRiDzfj6
yKyRmhpfnFE14U1aoL12xoVeSTn7lkzJn6pCZi3TQHSwUl/wZmyDhNBSdSurVOCT
LUBmuGvA58RPfslCZxyFJzje+ln2cSjGRffNOHlbYMmKUIMmlfEjDrfsPvmpBbZM
cpyrCTq6mL5YeVGWdbHbqDlXIWkcm45346jkRikgFSDXl+iTNbdThHI81yp0zy9v
iI6Vvw59xXkhlXcOvpkeKwElD/3RBKNaoIPB1geRgSdlPS0v5GZiHbDgGXFp2cPr
ukwa0qqGU1AeJtyJHWPeYnlQGGqPB1HY7G5PrCYkrr/L2YyNaU+pPulccsPl6SD2
/R1N9LnH8GuNUDQfd1EPwdU7HBldr+0D1O89MU7qMWGis/NWN3vaEKZm3ZSMU77X
K4QazTL4Opex938edUuIhLaRWpPNnDCFIwGUE5S6vxfWckXgo8nOKjpgcxSXfBOR
cah+vzbHxTJ8P11HAD0S1K/d/jOCCQLeOl3rud9LA9cpE08jIn45e5Z0voaLRIfU
XTTUB+IGDUyqiWR3EmQewrk8iKVqpup8gGZknA71STOTupRVBXceUI18pUsA+MCY
27wibh7ZWiK7me+Co87ooi/eZX6oKCiIRYWfIQuAp5kR2JJIzMIPdeYHxvxZK27k
9GEE5CFZ0M/ng7RsPYX4QEEa10Nv7xxXO+AOBgCDbq0VjQW/RkLXmD02hFQkhXbf
jwoGHQra7v9keo3p6UzxJmCYy7W4lpmL7FK/+Br5GOdQ7J8lD3kFpH8JvPvo8v3S
EbFrexTmo12lnlH/iuLlwdTqPwFIK+eSGc5RQiBd/q/yZCItD6NmPsM0fQ69g8av
o5bp9qSvkhRNfEW6R+kFh9iYT8i05xpnUvC0ifn1HHOdmynbMCSYqX3/EsbHL2Wq
HYXn/2ZZkPJBKBys6AQu8mIwtNwAw6MHtKcuF9yfNHzKlt8C5G2wq6RJMR5pbD/j
dNPqh4hOTXgzzeIbz5YPIIGDCoWtyv9r1l2D4S6mdTiD/KEr3urXVuP7Rlax4lhC
7wCXfOxDduvmOluQzZ6seHHpQYyjNix6C/9z9XEBrnFn57Pz+8UQWH5BaJS7JUTw
6rcengB4VnQCzhbO/F16/SpUtvUuGDVD5eksiKz/MGQfTx16pwIO6tGLSwvNPGvj
Lf1fuqaZkNAwjWPB0sTFR3pY/AaBKTqjKcqRtq/RrBJgB8eDeRSkvvbRx6Zj/MMQ
j7CqPQdN4+trKBcy4PHycGgsrV6uLjuoIEhjaZhakWp/lhezM9OuaHHt2KXy+VYi
I5aN9epe0f8X7JzQSwS0bXksrpvEOm3gLAGBS3AYB9qGZAO4hYN0UF+sryoMrw58
8NTykbubrEw10DFjY3Hp1UmU9Mp3Dhs+GN6xQZil985DboEXGKa5W37pULhGlu1m
As1GgfwsCxENwD3yCq6sL2QX7pSx+kvkSLIyCpt9tLB+zsYMzRleHJ5L01gFmc/z
uDqtQng1jbApWAT8JcGcVKaTKBhKoaijVn4vGDb5laAvQJ2f6l4Tm9Ws2izGsqCS
EE2UL/aWKRfSXP2PPY6jS64MRBP4AQaVyrVOvs64p+UOm1s+dd1fQQzSuF4S+DvR
YDvZE1S1H8MUFenoI7TbGTckAR7gQOIJAFe/2PDMt3nYj8xmsERw91LrQdE9gRXZ
0vVUo1w9CFSktEI7AsIua/fjqayGoN/nNGCHxuT8uj9mYiL0zq3O4Rumx+FMqG3p
U3M30xsH2/9Nu3qoJDbmjkEXRObZQ6tIcP7BRfYdToHK3ddqfv5Aot33SbJBxas0
5pwUeac1hDkzfqf0+Bvxq248qfUumn1KFP61jAm1ajcnLH8vlKv6yws+MI8CbBt8
JVqliqrst4n2CXpinkBImEM3EfhLrAWj32OO5XtFCsKvq1tQCKusO7nzGl5hLViR
QVUqGBvA6NBB1GcN6lNjFgB9NedN5jtdhnA+/Oc+1nbjQVc1fFkKzXCSQp8x1lRu
jyf69PXQvisYPM359UuR9e62mvZABIjsLmCYZml1f51RjnnoPmHHsSUy/Efx3ndR
QfUVW6I/2pzQNOXlx1JviWpM+9obDQ3vGvJS0mSZJzM5JNnEX5Bbq7wlsWsCVumQ
DFKnxv9YQDfBCLbkgIB0AIWFRA8CSgRkj8SEnXGbbw1QwlzzwaEtmMeSWT+Ul24b
0+X7l6nLgQha7IN8GrN4LVPRBMpMzqjgywzlYmVdinD0vjZhek9R90VgV6xwgde3
AybIxS285MhAiP0Z/GZIgJ9AJxbNkrpKoadTzt3ee7hreRR4e141Dll/CmqQ9b+P
utDo2Mrt/4yYNQA9eLRCfSl1MuyOq3M7pxTZeIVwCuQXXjyF2OQVqsnxQjT1TYZi
DXp5FJkEkDQkr4vYUBcMpfoIwU/huME4MV/QiDH1azh1NhqiCyahOs5GSA/GDbH+
Kq2SoAcLgQGkSmPzU+EC/JztUloyu7uNiOQ+mzTz3tNa7zrjgmv/ZChXV0vI0bQe
fnlzkkSKu238UDHPumygsbNKmN3KuzoFAqziak1UnGV17ohZIwMn1fPum0/vkcKg
FrLp9Wz1PQNt9P7G1J3z2lntp/znZxbAD74MELsHK7pgpzn0F0fgT7pgHinZynFa
BiBkG0RMHGzb4IrkhDZSsAIl6hTSc75MwD3UoKP2wiSUDoQIWMoDN8+E83awojYE
B5q0WGq01LK9IzfvrD9bfKwrKbq+gr4DFYzCvhAibgrtrV/n3NUbk0Ul8DbrjpKy
eszEsqrZeApGyLgVrxtbuVICJSSYyeqGDtBBnocXvC3Z0FYXM++ZbQYzwehuywy6
GBK/gOZGx+9bZg61Q8ijdXG2WEsfjYZnx8q2ZFvKts7uTSuLyolPKNyNFZTc/sji
Vu1KDW4gIFtnPmCGvS+12CKSClUhyDtCh+NW54hJiQAQEUFtZXVSz1YJqCQNkyI1
rLHBmXSoNXZL8Lnj3c6AGZWT2BxuAO8kZXaOfdaKmdo275VkILH8hUc4DCAw4Q9d
p+gTFpRaN60lJeTXef/vqlCdsT2JdVOj5j9UKvlKEA/ER18tdmr3wSAATB8nVMSL
luiEtAk/5XQRndiJ6ias1yoUqokdEB63lAkz7HRlKHb3tGqjMk0QddugxAVwiRBe
/e8X1rzrku8Cdy0yMo+zMLw6oIK+/Mw/e6N720jEZ78qVwTrrOe5/BE1Krs6px7t
SkbmImz+i/7C9AdSeb1TbOU5LgVorSaNMdApQZatxgEpYIOeUjLuU48jYc9g4g+U
PUZjDI8WzlJL4/41S5ln2UzHrt53ei/rTjGc/RpX0H8MBi5PjDtt6b03v5ZMKUnu
TV1AdpHk5ntzP6iiMfaxLwnCt5ZC7QNd/rA5+5htxpxChTFSRZEvLfbU/bo850dM
X8lErNP2Rm8H2Q+q/ga5SUjF5ynYpKRp7YZSephiLQPkdOBla+Zjsrw5Ir5+BVEG
96mEeUAkJURG9P+OH0h+ylrxbI0qT/DvLXvqAsv7KKA/9EEptZVm9EiYzFhZ9wUt
V7xVGs/79X/GHT4e/9boJeNWaHBXRU+rzRjdDxd4re6qN+Qu7eoRL3J68ycCmAnN
Rcs5ZODF/UhFQcONEYxqKAoAe83WjrgrQxDr+gC3EqCaHVgEZLUB+imjvXX5Z+B0
bN79qwGn/QETJpJ90clrVXnHoG19/t9MnfX1oVo+SCrmKlZOwEndINFxOzn3xJDQ
d6EJukqEHvxP5jRWJYT41+ppZ4Zeb3SoqeYjT1pyZvlPcY8vFbPrRpyU4tpxLbhN
IE6hQrn8dV1f3AZeR2j56Q1KphiAe7J4jZcEjjoNzt4DNSbc2ywdhFAk5u+fSVcw
/OWsA5TztnqPDppwwACuVn/T4CfweM/B1bUHk1Z2r5VtylOJVb5wEzjkL445oVtP
f98dyXese67nSKb173wX+jqKoUiBpxWNtNaFHR25HBZmxaE5Tc3zcxCrLNxbVAsd
lr9Epm4hfdyoV32fDfo9M5grNDp5CQITlGKi7tLdzEaDuiSSZ0lgKMZ+lghTsqa6
H1qUHnWkOa6mA6M/GMk3pLdlmbt6JMFMevOX65kXPWXS3bsW031B5tMyGXyfv46J
SdpmhFkG9sb16nJZcRQtTVNbTDJ5SMjjzmaO343Mw1nYflUR/xPCbGmKdsEhjrr0
wQDoKRFmQI/zF3mmenVlIYWK5oUg9KTLUfB1Zidhv8YTdG3SabSx2FAG0/CpaYWs
o1B4AebNCkeGBMjgqg6hq1Znh/zdPQKwa4yX7rq9Ctbrc0JWPlCBihjRKKWHMABr
fztHKoAhcDhkjvy8CSn4mOl6o4VOwFySLhwD21ISFIrgKxbzTkQH6DEOYYecr+FA
Y+UFyXImvg3wNrjLQ9LgqTnl2wWv6xRNo3lO9yhaakjxBsrFewg4N2Se3pXIo3DH
IQkQjFVeqIGYOB0iXK2EUXlBZaYrj+nMi6Of0mp2RLl5wDHEYvpD6ii2oPjEIvJ1
fhe1AkXe5Dk8YOMlb7xRSxMXentYEgq7+/TTBTDB/l+KlyLwph3pdK+cqhjQqq5N
rIyI1O10aPN33mUsQ25neQC/oxvIoc5B8D8pOdVVgk7jCu27lExma1Kt62+yW3Ba
EvotEXaETEZHuanFa5AJO/D2g9YM595zZAyT9VRj+jDhFcvtwor5tFKSTEXU0szS
13bx9ILOK1HGoJV+Hiz+aj49oPhbem6KZkg8/uBmoM9kdmD1awH7YwXNU2LjXKzW
DeOo978fp8R8yd5Da76LtVFq6Q6xUZSrzcmKWz0ZGO3sevcC69UKhg9Q7Ny6DmaS
jg34UMk25VKzfa00/VGaef2fuKKzcw3zLGjRNMmPDs1kJgJNIqxEA9Np158ziZ4o
+nAc9fjKTlYiaEoY6ucpv6aiIG38YVvBRkFa4bNOVxhl6UF0kFoKxhF/HZMlCfYZ
p6ioxM4O17om01bhQcHmXH8dhuclEaz9jWnegwmHcDVPQuGOCA1Z+cAIK1DpBm1V
eJ36z5KjzHWAY+gclLclX8FuijrH+q2aGWglUXqqGMA3w8v/a/HzhEMcCCV64FMq
4yMY6tsZhwukHsGkYc/IPbdRNnSfcKD/I8Fd/GDrxpPHsZYz+/lerP9JrfuJTZuz
lANMxeRJV6k/4FtVwawXiLmAihCYp5quKaW1t9fkYI9ODXzovK3c6YWa0J+ZVjpS
L7ujuBjo7ybJAv5kMLneXeyKeeDgrjo0sDHoenR9a8AR1Qlr64zBAiYEAocQAvd5
VFbBDuAzgkLRjOc4kQAJQv43sGTaqnqohw0HqWnDJcEuqLoz6qAFu/iTjSJy9x8g
6oHex7Fkj3rdbW+4YUovw67CQtm8cB/y/mrzk6GoQ4T4knGdCzTYHSKPA5k1v1mE
cFswFlvRK6ClCbDpdIdF1XCSk7eOZP+6oTJs2622VYFDLORHKXRJNAkk0cHt03S0
avgcW5D4iUaViWUem6eEV6AHhnny50Q41Mzh5iVQlZ2SLG3ED29r5Txjyd01o2X2
fYrW6knF5WdqvN/AObfvO7c7S5NDCLIe4h9Y5GyF2xGB+FDTj+ZGguQzgWw4ecD6
uosdUKezHzzOQC+IBkL7yYWQgV+uDJKqTYBzkyK0nYiBSKb8+KeyS74fBhdWkOpa
TITWQ+74o74mYTPdhvR8r4M70Q0OtF6shOYp0FkPWqzOsZE5Yd3/lttQRp9gzOFP
rqg+jm4YO7ZoWe9e0WG5Jdbq2k9Kwa71Ha1UI6go3Xmpmf/Let7EEJV5uxELJPAp
wpLKkPXFmv4PnBPQxZe9pPydKiPSRVO0p40uYvTuTdUklVEYoF7e2PPPFoIPRY6v
+JH+hMft1ceCzEqAxZrN4q+YUnSnoUnyAjl4cpmovUyBw/wTKhQc4aLsyNccBrGv
80bhaWPfdGfCqNXc1C+GWlfyXZg5B2B8388d4jXeD54JYAl1B5a5QluVKHCRUhjb
f5OM/qvEVrZ+xr4ugF2xwIxdaNiOoFI4/w+p+ETXHoyzDrM8d1R5ssgHbko6tviM
IyHLVnlBLeS4oORFLXT8Q3wqjuh8DHJpXGE9XjPX5sEnqY2x6rxfd8vhljvQHYQ0
DlKYS89sfRZGVnIpbV3B9h3dhDEb+PstdCNVXclumZa2elZD4Ld02ATBJZFPpoSb
x2g0TacswAtMQ6L+mA8xbU8pyxF54fRyB7oYM9xzc6cYMmd9yw9zDLb5qV6TCJI/
aVSbhUKyBiHRg/lAlHqi5ZgfickwE+TR7njaQ6sI7OyYEl9NOxTjcQITQ9Wzellk
tnO0C8Xl9I2n24uGxcTINRA6+QYvBwlOI9M46BbD0EoGy0Ub426UFf63w4d6pHwc
eIplDykibhAX+LsoIn1nm6ktVyVAkwpr9SUUqo2Lk/qnbghJp8VmxNL15sB/PnnL
vvp/ejSqNTwNXV/MJqmsk6dku5TuZySdYd1Ytw3thEV6irlDVC4MkVk5ZyiWcV8l
HvHY23ZFF0W0wwxuDJuiaEY9qDVBVO4Eoy+UGkf3FTStGloRK8q4hCd59OS8ssXT
Jr2YsmnQofqQJ5sgtMh5zkSy1QAVdW2N5ZBtgyzT9eaIuvT0tUoU09kRDPJ32mCF
+gvVLaFsyS1lMyKlt6b8wu3UiKMuxGC4buPmKSBQoW8+lZiovKKW5bmycCD9XguL
TBkeKVIgPUYpkyM57vNISpCYfhMs8jspAjwKoro9eb0Kv6CHBzhSGLquYzUdbcfK
/+FFZIXL7V7X/uUE3l3a4J1SkakLfxALC8hnDKr/bNc54oBouJXm0tytqBpz3xWX
O9TlcvIOByl2uxiLm3Zarw7uAFX22LTh0qZS8vl6ZxbNS4uhDZKM6szpvc4V550G
Ajv/sJN+A7LmnVrnD7gWDfJscxLQfdvrrZLK6m8JQ+EP+iD/I9CCpKtEaLBjARFT
fidHuSQ3czCClrW8hNXahyo/HfJOZExCsZbFmhea3jnV3CbRiqxngL+ZIz4F+ow4
mmnaxSyDi2HzY9PH46hPSmPy7Dru1q1sCcXPbV2a7nivhbb1gueKsnHROLS1BL31
dQbXbD3l5jXm5zx44ktXG38I9Hk/EbCtblhfxwg5KemQoCkI1rAvTbzaIm5eatC6
rP1EsF0XyBxMzMBDy8EbsbP2Mgh94gHLABfkWO2V8o4KWrrCZ/bVG8ubiQaRzY9G
6eh5/dpzarbvnUfRFtDQ5sKCmxRue0wT4U257JMgU9o8JoUfeJYWSa7ygeqt1b3E
yqlkh0J04eifK4nWHeQSHLW792S2Xr5mwqmJNE4w7tz8mJfaE4nOZXGdSt3y9OTj
T7KDiTodbXWAkyNH95yzL97jsZAXj0c1HIZCtmDXQKD/MRwI9m6VmTRM7MvjhvSQ
cURUVZRhZ+7YNmNrFJhT/aDh4dSGGfa9HZDexbGmCuZv2Tal2VUP2Hn/FJj8N7rR
PrmjfsNCE/L0xWjF/dB1KnZCETa7RXzrd1WSeg0Z7Dfkd7p+qCQDlwWXsu7EvJ9v
vRv/72UO0VHFlMRgHQGDeNnPqKxU624tz9KEXBZKOWBN8mvKKKLYkiZNU8/6VvhP
YL5z7YYS8SjnRt0LdGwKSTuDrg+lA+kwSbqwN9/ksi7nQSODabnsKYkvnlAFr8DC
IhJGgcK71V4mY8tKwyeOntRQjAkqaB3BsdVErI96YFiZ1zTNeXSFe3dOwY4LtDxR
LV68ciJ0fhgfRbS6erwf8UsyFFDds/lC15llAbdLbkAwZBDSji06C6H3mmincpez
j6ttQtrdfNAypPZc4EMc9e6X+cImKwD1BTOX1IWcsUergDu3mJOOrTc1VHRWteOz
LERrlt4bmqQs1g8Qt7ctPmP7Ak71QLsPlrBxxIcy2olYQtq4BbK7DFL86ocgGE8c
QR7Mmsc0HnqXRFJBq1gzgEQ53j1vkvgvEKx2AwyMiu5qhDaqJit9/A9DH5jUsKxV
IwxV6BVIxM0NUYNeGTuAf5+2jHQWj+rQou+UrGsxpfiHfBMUjHoJObr/R+Rp3Kfm
NVHGBbO/t/9vNJt2Q2rpaz0fCofBLK3II/h6Inft/DRNvXUBh4c+OPl1JbqAlJbx
ag9FNc8clzXYIWG3vKVuSfOq7U5FCFu3I1QbWZ9QDwvQ62VAdnZl3qizZ6SZMptY
LlN/57nGgXF2/8m1pre0BxLatD9EGe1aaxwzTURzdb8cE7pTnzE9mqI8xuxLQhDN
v0/TExMXQCglA65p1o71hNlRoi473u4dx3KFxQqIaHTnoWvnOz4h6/5w+ViSbVWF
bC9tRW0ogYeMQsnc5D9IhiWUGsKvGRdfkxYx3mfZSogNjPj0IDaSaR6dcEn+ZGpm
ItTT7AzKxSrX0/oS6sRdemijmMtp1OHmFyAPNBZp6beSCY0f6pmBGSeXLHN+zGxs
3vqHZLc/k3yS5TrBJqT6Eo18g11ALqnI8fiaj0KAjhy8gfPLzbIVVNOMDM/2eaE3
ECUxgvJweXfwLnPBve94EzOconjhMUPvkWDceQKslAFQLVG4U3ZH44JqbiGHRkg5
DDqs8vntYnJmAwZBrbbElXDZiabKCI6Wvj0jUUZUAaP7EY8mYFpINkZd23v9y4D4
nwsOZx8SH5ulc8NEftcdcxqkZT3EnudKebukO2qLy6rlKgb+kFey/9Z8TG5OG254
TdSpyEbs3P5AI58XHb92Dq6ghG4FDtkCjvTfcsy/smmXY3yeoR3rpgesci055Dg9
Jdsvu9IHchceSAivcc9XH6AbHjHQPaUF0wIv5JA3OiPxJ+kGZUa8svjpFmGZHbfv
ZTBJQBHB6iVk8C3A4KiIfdaQDF/yAkv2QO9CrX9XeO2rriyov0LtosCUm0uY9/TL
hsHzrG6g3KEvaZuISdkGCdajZa3jCAfRMO82u+9ZlS4bTMrD6by3k9uBtCpR7nnB
8EO6HBpMQXqeFoBoaKoG1T7tlKhdTBAvxpPus1CPLZ55JERMJoZ3woSA2LSPxTV1
TsTIL5+Ls641wqdi8S3WYZPkgmMX1yQRAoem6uwpTtphC2cqPaudYPd51OOxaC6P
mM0hLc2pHBtaMbLItJlJjI9yeq9/oCnbesyAqNf0X3dMynyzty6JGA6nqvJbslp8
aS5O1M5aWIC51R61oT5kgWJLAC2BmCaT2jBYkZ8+4mrq3vE/7ZIy/Pxk56R5vRU6
/wpQ5zaWje9XJ40Ig0wR476YXrFAfBrLLXlGit3K3CbgPwMARJFlrwR8XINtVZzN
XhhAyGxOBzvynDmg4hLONQi/uRQRXlFbOiIqEkVRxKete1RUcxcKoh1vZ8hsnsqY
Xz22XLSuLPjPZIaAAZruMMHkqGpgDf8h63mPfWU/bF5bfSQ2CZ711kJxXY+YBdKY
+sqZ4ABD8EQWZJnBBx/iHaQbQFG88dmrNR6azK+tqM8X5LKTTewZm5mHus8/U8Qy
cOp11B3fcwx5h5SeoiKXggHl0Ihe7gErayNR/Ql11qQaYMFtZyvA7nhD4Goo6IdF
TDp9mHXySHwmG6XtRzQmcNwbB1ltdBV6I5Box77TsD1A+FYI6LIRcylv1L8scAT7
9/eWBG/tgBJdvM6NjRI10fh+EtCDRjzTo6dV4Y38FTS9DEPkYYAx1XrqeEdnnwLU
4Nl7t2I11ypivtv+di8Dc4fEh6MeiHSZ0fjh+4+DW2iYypMZNpW5BpOvotVoWgx0
mx0Wcid3q0d9ulvIwVx9lXlaBOa0gJUU1jm2AysXRpWhdx6l92DhMAwrLsVtn0MJ
09Oz0rLJ0H4puwgCUdlhLtc+ElZ6gI2hHTS+4Me5fomiUAI+ZCCekAYVVMLRv1qq
ykqS9dc43c2kawxyCj24laFKIcvVMxAyczfYw1gN7Tj3gz9ulWBubx5iDGNOFstq
+wjKfZ2lebMIilM+eBBIcVm3bvnXJH85yHJSOtj+nx5X7wRsbbY+uSq3xFxNzENG
QMVWAH8ggfctEsZOG1OcUtLhby61HhRkDRuRbHHRlJSG9LpARN0agMaZOgWB3i/P
ifit1clTKtDfe3wAWVBaqNP8vBuQqNsq8PxJTN0S+IsLLwXfNkxMtZjgTvqbQk+f
oKXGhWcQ7d9InvWpSWhEjQJwws2dN7ks1+8F0SCXmqsiV3ggTInChb4CY15AUzGi
S01sbZRuVSdzWIv2BsivDNPnxkJ906JOt/rbD+7cEVuSV/lyyVqWQcTprL95BLTd
1JJL9QHRCQpIxRGyeh7z0ZCoy1ECKQg/Wygi0/vm4ewV1kUdTvRdAWrWy/qpqyks
6M9FoIx/oco4qANZi0QyLLGrtN38kIwYzfgUaMuWCAkr9HyEya7U2apH3yQXDTY9
2knZZS5emnuShG3HUwoaiSGlu1RzIj2fdKS4zNEbiLv77O77YHcQpH8yJ1T2pbuQ
Yf5zYGl7aZjcFGQrYnPXHAswuBJuIgnha+t0d8CEdlJyLyOG3eOLVv3p+jW476yY
/RgfWtpyraq/4clobJHnA7jEoeYKmwtToSmNIRXGHRn6dsswReDg4kNNy9n4XKwL
JQe7AqAInHovI2YAQDM2gaL6SNY+BoUkRpNWHqC9caIRZ2rnlf/hzPZwtJUTDnl/
U8GFPIeJSEwBbRJWe6ZD+fT6GVbpu4q9rBbA3SaYn9+vtAcLAq4Q9/uOMtlS93gH
wkh+PWZn2N6cMXdmrvlvy9BHT1wHR5ZIU4+uzQq5uhe+L0liK6lb8FeAazI4pfJ5
+g6Wa0b8lPQpNkeYdmEGx1zySyRY3gpzzJzICBUdcAfp5igm78xASIIOfuTxg4Ob
x53iJPNGQnN9hFgYUCUprNJuEP/D3qELDFyABYmY5cHBbyXCaq7dZAH4DCfTnqAd
OdKq0k7jOikB6YEelxJZ20FtufDjcwQUzKWFbg9b2NktoPl6xnZEQep4dNgrCVyC
JHqbwPpd9Aqjg0hyybME7ZPIhDKOHtzdZfVgAZ/uBzJmzS63Dzw3B0jmGzQ8DWJI
6uGeCztIetB3XgL5ii9tb1E71kOb6TIVTfBy5YvBV8wTjymZNOvpXghfkad3QR73
+wmdo4qmCpVXNey6RhJeo594tflV3tEJEBykP7Cda6XF2rQ0WJ+iUcQ24mA2ImLW
czdyVfJYof6TH74s+oMahF1TrDpLBUz5xtWI0oPsFFurYrQc4LEel58CPSjiSagl
vCZgQZZIHygOeGrEkWm5dKs62kqTU+j9osEMG69xC/CiYJrrqwg4p7HJo659Fvp0
RDFa1O/Zmn3uyRryvkgW7dRdfWdBxh9Q2hJ3Kbbb06ztqLfEFSh3NLhPLUVE8pUf
BDiyNNImn9QCIMXov/V+6tmoxSKnjKvWCiHBzT6fPpgdk0J1J8lh9JYFwJPRhosT
4Zf/JGO10HqXCtRB1oh5iH6axfi0zY/qWisUT4JUQjk3fKwXPWfDmIl9FXaiyenk
06oU/lxi7cAAwSH9h+SaqB2ww6s+qvFBnljwf3/9/Z4e3BffiBFJoBSkqAGGdneW
2A6kjEBLjWZ5o5ViDsRKBKIcHnk6zkXp73F93qtpwUZkQGP8TGnjnyb7zLpKC+vY
DXfmyFnMVYRdkZTZh3FjcjhfNjLCqbylV8YzW7NgNJEmcw1aK9Rq0Nu+SOuEG/q7
daKZG0w180fg64kz1j3ZtrGAcVDjB3M54gI1nxs8Mvoy9QluU99g/H+WsfdOBvsV
XBnj32hWFKmtW7515Ld/MQQ1defXD3zknmVORGMS2vfxfW4cNfJaJjejHFjmo8h8
QBn6CPhoJtmoqtq88BGg9DpgEDME1fEQPGiTYMEsHeEOuqVX/+ow6QiG86BNDmGD
TIvo8/2aduMZLOMqWB3jBXw29p0phImuLlj+1V3TI9AbvmrQ/fi3VdPii21mxz2k
Ozpm0369VJf+x1SmSRggYREijxAfIDB6Bah4GS34ewoHi+NCtdGS0nQEfC9u+IaF
7RteNopL1C3duE0M9HA7fK3jMMZhVUJ0QbLkM7LBnYkiZXkCCitoQ8Rk8bktHC8a
mzbgUV6JH4ztwFL5PuOgIC9vTUd+9wXM/LMsMGaFwVwzV2rZXdKlLBM0NoproIPu
4k/d0OoXz1wkuRnqx/rp23quicapDQ7zrq1JjtE6n9t+79sCnmWGCxiT2+VmDMY8
VVhs/S/VYWtTVWVlo0BoQxiC4epBrOmD294epYeArJoGTlz0cfLcOnAyz+U5xt6I
bsYd2rqzaI/2gQoW11TQMBn5vo+ifSahvf+Yzvuk7UCfZQDzBkOI1br7kD/ScpXw
CEJiYETEGtRFyLmLC3Yp4zy1rCFktoQNR/2OU0U66bamrC9UsjU0R8UzHmWHCe5i
kfph8VTDtub+SMBSVb8IBr13fgZ+lV16OcB04RMt6vtRoimDUUzWpWPRjfq1yJmS
9WZmr7dwtjjkYzfYRaBp7H1ao1xwEOMmBJHdN120PFvCtJsSzMMaYQqX6NN9XcXl
16AQbHMFskbfwd7osGsBWuJiuRKqOLbWLj1OxFiP1xyBPgNxHakwk9gBObFcsOQT
yIt2KXIsVhprbPhNrwWve0FLvPXTkXCTYh5K9ogxhiY6/7mlCEO5vlQf1wtgJrgX
B4u2GyZani5DrhVa7b2aBlVZQB4wNq8IewqyotleSiYpIZrxnOyHKc2TsFP/ZhVJ
iEzAc8g79prZMRTHDRMzbUDlgp8Y/hfbYWg5GuctuplBhB/nwYCYRyMkLNxPSym2
ivB3boHwVk7l5kXCSWSm+BbYDq7yrkkmiNAD8EicY/bbS1RETNh805xxVeFKtJ4b
l/HSLieUXFMuud4m6DuuK8DkKRdLA8S3b2n8eD4FGEw8JHM2rGIptexWHpy7WBtp
/yecfLe66h+AWNWk0D8AZFzjqZbqwg2eOblgHMzWwJiUKZ+n3etivnHhHCQocGBX
69ssjmgq1vscVcwQhReeEfxhhlnZaD9Rqishy4RTeZQZtqzdWieZI0vkm54iiMRs
Qj+aJhJoFJz8jwS/ythDJaKRH9WXHgdOwxL1vJ4p5CjIUylMrbDMs2wsyiCmYNw4
wbPDcqaXfEXTc2Aqx8fkzRF5qOlzFmcgQHUytbKBXvRWlhhgkNRJkUf1w32J0x3f
oWaxUeG3a4z2LQm5U7E2oz3d2ufY6Mz182O59sRMBCSSnXJdtgBf8jJJ18zX4Nmk
T9iLjSOwz730QYj6n4NPys6qANmcampF5s3Q/8b4ypentB+TKnmoillwENhAaXyB
VUqVm8OKuoRPW6RLYxWI07jWaYZw6w7wFUxeN8N8jT1BG8GNdWKHgD6/tc+qk8aT
xqAuIxBBozBkHsxPkhFqVHmHFL7gv0eDBYzPVwjqSYkYjzbGu7OPATps6UiG9D22
FlJyrK9TDfry5eh2r65ySDdXX8rfUZEQf+vO7b9h+nsQYgSq5I5j56M5yxmrVVhX
gCNKimG3/bbgKJBM0uQ0OUdYKRBrtfSmur9w4JoAX+Kb1I0lSZrOm6Q9Zok1Lzqu
/Uq7AQzecrLHYSspAcnVi/bQ5Wa4mjnsISWGkjFkdboS6VAGhEHRbIqoSI7B35so
2Ioa7GdK/fjdXaeGTz0wKc6+7TFadU+9QhsLdhKBzyJaf6uPqPVlL/73lGaKQ0kk
7axzCYpNR7Z/Mj71HT9Zns9BQuHhsSIZCQ1LPZ+jBjUQYPxF3VOKKMWG+L0TM6yF
fyYLrYHO3s/RACdWdwV4vPdnn+AmQwSfaZ2Si0xtjEL7H+6/dR9ja2L4J5B2kCZS
p8vgjypYaRy59zeizjbDrLpoh8Xk18GzTIVsNEiNGHyCgC5jg6k5dTa+mHZReENC
30xZcadnhPAfV7NBT4NSP2DQRwbuL6s845+ZeXL6sg1NyegGUAdGLpuG+zQXBSd9
xciP8VrcCfXVfBnu82GTTbyz78q+pnSth14MwMK6ASwP3d5Tk7yTBHPsuOqQJLj4
0NYhlI//2uRc38I3+G3dUfRpzNUx+YJbRLDRzBjSVOrGYCgH/c6yyU36WVlumf2H
khfotNjKEAFFUbcDnZIVzjM9BCAJ+zLpK2tyvCD44KR2VSFbVRoXCktJb/XEFt5L
5oRhe/AO9KcSGM1fGZQqmeqPBJ9z0rBk6uDsj6wJChelxDUzV+/Dl7gPM5VFHs+h
FMHA1s6Wczghy8KDkJxFR+Rtg6zukP8dWkvioYIYxAAprhARdSlpdUJ0Fst4o5jr
/+FETl6UzR0325C6WIpQ4WtRrj1N6NSywVsGfZU8sMk0SVFozaweOrls8u1l01F/
gXIvJNBL9xlC/ReVPOqQOgOl5WcrxYD7JMcZnfjYWlgI2Rr7s3l9iKXgzpnDxTun
MfVt/aCq6Ef8sOTnAzuPSMs6Kq0WotucxwbvcLL70a/JjILzRpH8HVT4gXjk5lzV
j/sXqVdjM97ZLKZrLdArt83D/9DsYDNGwPP+dgLoEZ9cxK3hvI8NDFQeIJ6z6L4L
7UWceIKNA7PR4tQLjqoU4QOB28gN04B3EWZB79K3eUsCgkNYFpw9r5LWlsYYUrye
9fK3w06AgXpdZdSWHM+YmCKCrHpySWviGzWXjV9D+oToRADGYY9VyA4/0N/p9dLs
DHGFeFa8Oa6bxuaRo/RsuyJw1nwm8bMA2X5Wfw3OJ3rLEQM85S8yJBD8V2TwUv4F
3rps1ebdm7M532n0klwv+3RKYNrZ9yjhNmMlWcvzuwG/2az+MdW85gjnnHJMgZgh
MEePVTgca941ria/BKevXz8EU6MW+U64whe1Yw3wp5UH0T6Kr3q5KEPhhyxiJMRg
bdm0Hi1ATXb+gBtQdNyIQPEIT2oPDXg/I+K9A7Xx+r+sM52AScFxB5YYNcEyNxpD
K5LkRviG2UsEI2pzLhsBWOZje+NCO2R/9zn3QX2bUAqoY2myc2rLO9rpaAJQFeDW
2e+ytf1Q5cJKF0PA94hehRcV4EDNr60qiLyVr+upovi8L4f4aapIey8ObvCVwj62
DPBSDSRm3+3mqAJ792R7MvO5ejaT1A0/9z12b3jAeKjnYsZedjuRYAK5UPHa7tMs
Bs1z7JfSSKaOlna9JT7Ijj2VcVDqXCQ8030fkmqxtB6D/wkkQV1FXlvo5QiwD51r
KA0ouJCwyE+x95IPDpNn3TaR9Ateje5gIMHY3cwDR/SH9oS0GcauswlQPqcNIXhm
jRI3IjV4kiqppZtwsZ5B7j3mHq7Pgo88vMpMQY5QIO6dGJwsZWAQF8/73P2bK+ei
6CZKAWIyAJODVk4Z6OI5DEQao8y+3gStbb1v30sqkm3WOpy9G8aq8PjDyTJiKqHV
Us5Z6qLkdKQT7nABwMKx81zl1ARdSU/YR0Mhg47LtEjAPdCz/IF4MDiwS+wvM4d5
sHWtLZVfRdLJSm+aXoFdCZEyWs9dDnaaPZesYjDDq3tcxq+GDwcNjrA5SWj9FeAq
gJgSKXm6nwWvS5hVqlpdRmFfxErnJRaet5hrt2D27WnnPMs4tH2KerVF/Yg8i2Mn
cQPV3A1fE3sOokBjKSk5rTZBhq+2m6G18kClCtgCn4WJpzOEsWNDW4sC+FTX8Kat
cf4dLfngs2Kpsq0FM+SFXKfoTUbXPYoUCttxJqtPmMZ0H9kQoiCHGEIp16o6ewgV
4GGR9eH/0cGu1+pSvfIAWgUp8x72NvOJI9xHSVOdNFeJ842xaqTZnQRMo9u3TFMs
yf3AfD6l7rBRDOVAo3VJheyg9/F+RDT2u1re/DBZdHgtv/QGwrPdZpUlHL/wQWxu
iXjYWriuXvB83eYKTkeztIFfbbcQOoYIUUMIm5eYWjdmfSMHP7YZbgumqYX2Ct3B
Ya9RnEEqcsSlHVx3Ly2NAi9v7xEdrd/m4BF0mz3/zemlwOzCZ5LxckC7KmsXA93J
M28yn/bb3b/ienbDCcpkoDbn0UAdljRWauVYcRabW6VzFFozRYCNSmZYioYRECqi
g6F2a5Tjbt2Uz/aJkk2jQAj3kzcSEsPkhZ5DoaYbtewEF+VMQo/NOTwU+D7tJqsH
2CNM4LuYbfNY0Smd1NLLTWX/L5UMJGEGxIbmzYVd6E88Zhn+5K4NbaNcObc47mZj
EZhpUDvMqoxw/Sw5W2fKWYvk18A0FcFhC8YpBdMsoERURD+yWO3eZtO5Zi2dR0+O
32Rqv4cFHIMFZ7nG2+3eH7lRO8u6GGFuha/3kvm2RSkFGsfI6cjEN9W66Xk00N17
g7P2FC2xHmtr32YtJ+M41bVD3TgWcvJzllhz3PEq93Z1I3PMCCsW0/oz2Q8/uA75
yXjoKDm1VdcUQJl/FxdJ7jnKorXirxE58KMd79iDjKFQcYQfvrmIo2kcWp8zCT8x
43Cn5H2t6FcJ86UOyesgJIyMZS5dHe12DyMGv1ZPvlLFEqkFCyouYINx22i4oNZ/
4zM5UAkT7txA94qVpgTaJBqMLkoFWZxjXQg2daKJZdXvI8DCTP6iE+VBKpk86qP+
Cwz7l65KfiRSFq/WgCPBPNUxv6OX010BtoT8DMYTGnGqCab09ojWJ1sFUJJsyV5v
cTktJkmHFTfXJFUNu5R+d8NPV40FncrNm9i81geSbt+6VOg7gUUnR2wdurVqQAm6
cLd29EvoBWllKcTh7hl9xoqIciZTCddRbyy7BTI/mFHmzIE26ktiVSBzkfDgPITS
LcGWmDWCEywt5seigowxunWiCUF7BroQjwPtbVEVh8qvZeALahXcJV4sqW6WuNp2
gF5E4t23HzQ46478qwPx/4hnGWemakpZM2W3OBJsQdH/vrq3TqXMFbuSyX9Ojwfa
Jm9EwvUvXN4+fwExXIvnC9Z+LVBD+kFqsNrgguDkVWMRnE8YMRWIvcwVBUiGi4Ao
fr5trnRzOYhFWEZ9YV/iqjm2t5YffqDWcP6sgxyuutYIRW22CB6qAI1l+p/hDmqg
Lu5NC4mnncXwLBAVzX7fxbos2HCmKvtATNdKk5joZMXhmFul5bbYM3RWHbTIXHts
UUUF5G7pZsV4tBxoHGR8cH9tkcMB+kKQJq6v0ndebVuaej80Qs1dydEm23bTf04C
+eidYmCS0qYhXpW4Yl62ghfL89PpglM5udrVJeHLu8Xz19vyrWV/H/kTSYz+d8gT
veMLQVlL4fTp889a6a04g7KfFpFCtLBfLoZDLMavT/DfetAOw4/Rgux9s7lIdSPt
yvP0hT/XAd0LkCFKdwCJi+R+AKLGA9jJQu8GZz7uDBye5Bm8rXFzZ8RJLtLoSdeU
xSYM2lwzyiAVlseKaLKWfUx9oKUWj9uRvvW06OLAvoLEOMBQdSOEoYOW3loGoK8p
SbBGT98sw6idLQanrz7fQ4A50u7oKVOoiZlaHpBpYqxFU7AC6gP1tIUUMrSRs5EE
WWw0rYmfEy8aiGQCbiYYWFiX4eqP+aWUaSlpCHJMI4qwnuf7CkaANXX6w7bd1lxT
Lgp8obStGymgkKfR6W59PnB0kCaDJy17mrsVhM/NwAe43bKyzQOT6b4Bml6RcTo7
f9thnJKZdoE3hlGsuxxCRfTQ4lpeMcHIIfRthtUK2yuuDPZjm/+yzzPK6NUBJWvL
bLbAR2vdjGQCJ+IjXEHsgiq3+lRAE8a+X+Lj34m4sFs55c/Yg6wdmd34GzCxEVag
9abB4RbWLK9h6HpNn+clucZM3k+EF/SBuQLh8I/RZkBUVgXlvGmTgvy3XXxubTPE
TdYare2R677ihhQET0uYDS7RrCQVtigRXCHr182xpZ4CVcaI/de7GWhDOfLr8tD2
wfbfj5+DUHE7rOhpJ33pB58MH81MsxYc/7wrQvHNgxG/skjEGq91l1CILSo9IvI8
/asuFrwtrVjK81Dn/VQ9L+J+rzNMwnv6hUaUpDV2XgURo9MRqCTGvtv9BnUmn+5e
REceix4/0M9BnYgZOgBTtIopNBpcYDXX1B9L6VRcYARIPoCnSSWERp4DytBYm7T7
XCKyiVp5Eh5bOLvC01VgrZdKFnIWUwi19cbojE0uiiJmjt0H61RE6pThLRo6Z/4K
DzCrzPPpm7MaQyCcsm/MbbnFBFa1Kvu8Fdr8sp8JUxxnTBPOsqug5ZAZYQzhkMpV
X9GJz3gVk7Ox4IWFCF+NwXmxofZ7RMToFDUbBb4paNxtkjEynmGGA6S3ScCdc5sr
xfOoNruPYQcanM+vAYIGIgCXmNhf2vqw578azHuwLb9gkAMCt+Opd+Z7bRf/nALL
T0XMFh4bHe5e+txBG+IJCVTl2+afMIWo5U09mCFAwIKSJLBScnHjzaUlpPGt1fVn
rLZ2usRNRF6aaj4ULlqBapMi+qsUeLdeWsOvMGImlD9tpy2+BcGl3HQAXjr/Bs/c
Jvz8SScKc3PhQ6o4iAjXasxh9ImDPm6Y4DuumsYNsxHWXwM6GaPDcNOALKUXj5Sd
Q0xw08B6XMohnc00ERuNKZCQx/KHm0hdPZ3gwtoLyt8zrlCruYw9SGxdEIrZsM5A
daOwuwT2l+nyzHsYjS/g2ST/DScln5h9oQV1A8z6ZVhLehGdm6Vav0gyNZRwuFCZ
UNkZJhkVPBEjsyVnjWhGzpjriJE5vRMZSpKbRjtGkTjDAWHbazjrzdkDVvYLvX8V
eS48IaKepz9hi8xPsoRV0yykZuCR0MMxOIqsLP8CGH4tEF87ZhNvxxKzythBp5xw
gcMu92Pl+NI7XtP5LDt6maRUcLRfEDCGwtU7ERT3WJh2p2YKfhzIMShxIzeQXegY
a2cGFA5VKmV0zDU5wj9Xj9IMLCyFJhbFWSS+zhPCppAdF19O+fjak+AQ2phaTZkb
u2g913EagRt1cp8x0FDU51jJtU6asb6xK9MzmswlQDxSydgQT865D55inmplQ6Ta
sYqFGe9ZtLX5BYyUBneTnPLMTQz3ucUB/ZaGxPHvkhf1U/2GwGhNpAe27KLUr+q0
+83QlkrugTMkt3Fi7Er7ul02SooTu00aKXeYGHYp1yHWXGGlmb3p1Mf56owNfGem
AWLvmYejzMx3mFqN6iNecUL7CHWbCcRfF5raXV9byQLHOeO8Zw0D1A1VcQPVWrQz
I8pSZqLLgi9vzlv6FA9Yyy0mAxgWWtPtBSrXD+Ftx5KtxG6kqNdO25FaCR2w8/qN
MMK/uImdmGPDXP0X1UBTk0LmDgsXlktZsra11dKHvCCftyZtKv/0TjWIwktZoHon
t0IYTPxoNUGctUeTlVaPgt25QbT8Y1IHgH7TSMz9Uawbuykpy6jUiSCp4JyQuMYa
8hfnpE8B0qF2fFltxSVDHBAQ1z9JKRElhlT8Akhuljj6cDvj9x6/e71+5bSO3hW1
UiHGHPdaDaeOSkuBZTi6IN7kJU7QHKuz/8ZTGNSEP2/LeyntM8WEOC6GqPuId/HQ
GLuEl2WoMALQk79MNoD8TWOcSu2EFmomtgs5FfuOD1+Fomz6J1pcQh6QKgoAT1VE
+Nz9ZDlbiwRHnKtkIDh0s+WSHoFBb5384PdTDqxcF4wkMWmEEsFe+UALb5ILSnDR
fKNnAfOr9ijcT0jgHFwrRRNrHc7OTS+McbgYGEkObGKB6GcLR8rRGpk4bvA4Lwik
/vcf2KoNcekhJEYFvJGiDDNC9fANmtmSkWEsmTHQXIjSbBg89nsUNcfTrSORouix
V4uIPR5fPNg0Dzo5dtFs8ze1/7POiH+yE6MYVDD8m+3FvlNcxJdVub0ZRh1ZXpOS
RTccSG+x1yJnhrQHkkeKVD8OVEKddFnJLcmuiUZlmAZSColBLQjulNbCshF+Bskz
SdymsuK2FuDeEsawL6zxxo9LUmsk/ImN2WphFyrwuouEb0po+6GiMQ0FotSq2OJc
7ExBvUd++RAva3p/kI39rRjx1h7ht8jgulUxTav7NEU/iI/v0DD0UQ5Kp80DzVl4
VA/eFIG9KuZDkXXHaAXmMzaL9c/91Q/G4gUM/WxHWsGzvlCoYYU0+j57a6qtxxZ5
9jaa1P7AKI+rugpQ4lQnHZs4JR5a/rl4FYzWKXQdPYctM1Lb1XhofBhXNZ8s1OGM
mssChBoLxSXzEJJupVweItfiLPmLdOcCemeJLxN8IZ5dCxAjh4xcwfpUP79Ig60Y
+wBjLu4937cx8vBeIHmpZDT78Ng8VO0pNF6KzpKfzJfF4PEtYZxtATJt2MH+TcAt
AStcs19Onu119vBtkne+qDky8twyQEYrymcfRc2uaMYbIqdv4hQsUvNG+gtQlX1X
WlG4rv1qRLi68lmHlWOoLTEouduntjRlBISmAMD4R3YFhfSDgEibKoZGPUoNMuV5
+FsP/IDKl6v5GpZhncIeKY9I1OdiurZk7Yp1hEC1a44N7VHjRlnl2HNOgShrQiYj
Mg3zk7nLa8CS6bLuem1aU2ggyT0V3X5aowr3EE3hwcU4tY1mvisp8/bvj/NO/v/g
cyUAMgiB4oxZWxU2kYM7j07R8/Clc1nDGfzNVXi+AeCWb8NQ91C9UEaIxNawAo2b
CtOt6oDC6bVyQLgpo03zkSwK9F8r0z+kP4QOqFFlaauz5xENyMLr7duuPVL6YHaj
dDcTTl+3E1IffMymyADXsRI9Rv3Zv9CzwaeoUeYgItKQ50wk9Qx7f0lmJ7AHDT/R
kd97bLbdzqO3Qe616Tj5z2ZpKplt7NHOUaEWBHff8TA1rHGKsejkvheb6JbCcSoH
XNwDCAnB9h4IiMTCkwwC9IzvBHKmxBf8PCPI7AohyrqaZiajOy1kpp5CxepnD/aC
DQvBERMq9BDUk3SRJcxh3Zbm7FieNxepGDYRcTmk04mfdSNGGsCyG8kzdiHBl9mU
enDWo56Aw+d3jo3nxqRZsHp/eb73upgiViKWlqhVMpX/jXQC18st/R8Ro6rFDS8P
rC887cQpmLmbK1F4y7p9Uh9Whr02fOYgGYFu10fgkH+NxZ/BA88etUn1MjW2v+dl
FTLq7tgqpYiNgEurcnV5438ggWo9Ur/bCFUHYI444ie7sYeOr4oEsDmDarfwvGzL
fwTGur7/Bf3Ra4s1dM6/B8disv/ZR8/0mjQQOtfVSFyRVYGLrFpML+0qjvkr26lo
FpEgAhSyU9UqgHIyZ9Qsx30HLoVrakIm3YL3DwPLEkxsWBE+tpVvvlKfOV4NaBYw
7WjjBTCNCj26OhC4lEfs5GcGhXnNUCtWZBz+YoI+7evGr1/gZs+WN65JtyJJOzbs
nrL5N1XfvlPnONNEt3ionN6IzTrpGXtBPKhjr027r6Bs/ddJRzYsAkNgpckdgJtn
MsF6nKHvDZ7GHOAztjivCnKYVT24YR06h5wGQ0LICEcDtEMsrG10VWB7tSdr2jJC
ZOBcpOdJ/KjePndXuRweIEwZ8YJK6ZrNqQJveQccROKypOtnFXHqh6C9JwzDgGqY
BNBfbDcQKdAi8c+rYni3cbTzMGFmSzJJQAZXvirwZwYvN0CHMBydoJobcUnS02Oe
NN4KlJFizYB4iEnmKSinZLR7Ve2lVVGPAIrO3vUXepFoAi7r+ZiFeH5Tean2Q0iF
ozsbKpCvvjuivnvJealfUw5+UQ+f5aF/rKPDbealAaQCCQPcB5P3Ziyfw4lGO9+J
a/kMPdZwepOpTfty45l47QRludRNAotynSouoRMWvAZmAgpeCzStRlhNtt2pg4Jr
gnxrbEtmwcTIKKwjqUo13p050tpKWcF2FUBa/g7G3w99CFTKrpfrRVGjVpU5jqup
6i72OiveUst8phAY2kOTJq2/SYrqwGh3vFS3Lhts/RNHyekRRXriUxpukHzxlYo5
RoUfMLSFspwuiEjuSM60si/DVrgAD5tZjryjfWD+A4rDnHJw1NOiW3GFLxMMl9hn
fLDSX6cYCl2IFrTan1XmWieLm9yA/yNIgBDqAU2ums5PGmZ8qv2Xkpm2LoMM0Nw4
BKpJsNoYFy32j+trfmUDSSC7tbUT0mDfRYCRVjlZOURlALsrx0JczuD119GteaH4
rYG7IKBOpOXC3x2r1MonYEskS5J0qMrqSBjBMYyN4HfgUnNRpdprUsi4QGCKiX9f
uAMZHoNr9mhCGZKAgsLbqoHBPMtiFvLgC742whOiNKSKrwOYPQDsuA8iNoqwXjxI
MwMS51ltXTNeZv+nlAGRaK75cWnOyFzHqGYmF1OHTY8xot19bybouXvTXcCqKZ4n
6SaZr8vXS+fHLHryQtCQMYJONq1PuIrk+U8J5CvzSWGvbrLWzB9G7KfZGGm7MFAF
ZH8UL50XPgLDzaz56YS3lRKsswb7vjjviM9oa6yYz65zjAV4yg91Y3Dehm8wyb82
mfILYjQq4G8S41qJP1ci/bZ7tr59abR8QpMTggsbO+7Yzj72LGn+2tnK3Pe1i5xH
m8wKZwpTKBER+hWFt4bFt/D4b29DKll809EvswkZlb6g9EnhCJRv1qofTxq9D38B
9vRPIy23+mw87ftiPXS+rSaqwhrriqbXcltp5g7sSjij3kiEYKYKfZLief8hqrUG
N5vO6UG8EzWE15PPNBStvHWqihmzZWHb8x8XYWH+N4yZEgbZhsOrxcJtqCm8pcZX
6feYqHeTBED3vE6ffDA0CU3vzji3EtPZCKIv1HBRhJYLmUXNDO1i8tDWqGo+oqXv
ty4Xppf4rpIsH8SoK6PGyislQOYqCjFeUmdsG26eR8lY6Syy/PFwA5gZVeYLuMnX
/qnpjcmp57cEzf9IyINAMxbdUvUr0SjlpYxpNbZRUC/ms4KaItz2p0R6tgd+wWP6
g/sA0qEw8AZGTMUHJdFI8ji3TaK+IrawePUwjW3KigQk/RqvGLtUvgAjn+g4tYFz
qI+bcbYPouGVaHPxaYcS5t9M7jN5NUQ7HsXPeSvB1APBTEfx0m346gVp2mKolt5z
MGS82zgmcWh8tSqo9zfEqvVOEaowu9OEDtaZLKCBAdT1W21wPfaAMWhiawjW7tZ7
XzBYbayM8OnWM4uZXpUhdfUPQ119nkLfEAnRoP98duRggHfwLEmwgJAf5N6KIYPw
YFz4brJYyi5UCGstsD9Yceh96x50qC63NAoHTRwCZn0zy7xSajxYpUeZZZp/Y65Q
/Gweijfbht4rQAmGDNQUVn8kf3T8PPG3SvxtqXk8h8/pfpweHgOO/pCtDWKQf5QE
dI936tESXgJH1qRVjIjzh9QDxdgWvPlBLYOX2qQWn7AxiKs6Kd8TjBsVZOgQC/9+
EOSbMp27AZZ6HDcNw0hksUYlCjpq6xWfVljQI7G7HALJukygDxMTAC4BDMEO/Hey
lqJ2hoJBN+oCrKgdCiuSzWDhebYzBX2vlc5I+L3U6K0DE7yzh4tFrNEKHUfzNsCC
zz76k2K5uyhnTiulV0KukQvIjVw+k7qZmet812gFVAbaMd9kjVSE4FA74Oh5vfl5
KFlyEUY2ZhN8sWOHIpFIVtlZ0grrJWcP/m7X6kSJMnb5efupDINYGb7mLsw2OJw8
TBGVVGAf+QYl4qJAnjOdJntJIRL195qAfI89Bj/OoxsdseWVrY59/OPp5mYXy4sk
f0rnp8WbUnhgkEe68ctwdonJ3DCDwOnrGaJS5wR8dEuIOMvWpQHGabXJmFkSty35
X23vYBtsXWtzr7QFBkpEmBR157TrRGmNJ5zP8XiZfEWvTvdJpow/kM6fKOWSNDRR
hPtWVNEun8ja9tRQrOH2W1bc/LZd5pcP19N+MiPDzAclRW2lpt5CKWHjRgI92oDJ
QNYKm8azGqqvEWXoN77tcMMbguzOlMUdjvnm1cyBcqB8LwE8cvg1S33yCq5pae1S
4INSeD9G8lKAmnlvREY5plRW51d7Bf9/ZveAiktHfBbQ3Dho1TKkFsl2UBlJkDww
P9XoSxII88Y57Dwbyc85b+Be/ke2x5sTDny1N1K9JzNL+qu31ewOJ/GIDg5nE2ox
AwmQywufddEtIul+O+BMPo/G/yfUe6OXumOblh0iHvpMRt5YPLeA5Vqfo2P9n2AZ
k9r2CvOzVRA6zdRsdkzaInQcQp+ob+WP8ocpggogalJuJ4L0Q4H9/iaEDYU0UDlZ
vv+647vufVbe1l3GhyUVJ/3YCu/X+8oN3mhM66jVjIF8aEPHD+7uMbMumWOoyB8T
nGpL0Z0v2dml4ZcvLsqy0i7lUWzlwQ2t0KcKLI93Cg67yatZ9D4Q9L/CqL7ns5Td
BWVpsMHlzTLPrG/hpDBeNL+Flltde1e93hqQyhvRLN6NS+VYQG/nB4SaU9rvI8S1
PHSu4khRyCu9SwhMM2MflP96gbmHqi5vmJMGz39b12l/enbPIBwPxUqbSYyjhfZK
sZD7DWwZlPL+61AIIKXV/gczN1doml8luLynNxd/exRFJN63tWlu3M/sptRchoyX
fC9xU3ITUi5+F/qAx8zXMhjv6dWQI9m+6Gt9T3J/+JtQG6qHseqZTjzWlNXSLSPi
R+cO2nt4fTPzGWazJuyiBQolHvhMoINCke7ouRyWwejafa7xlZKbB6sEn8FHezW1
cukeFNfyq97iX4fWypupM5JNNbQmaOAPJMi9iJQCmQMgJjBwkpevz/tQJ2n4YnVc
AU5walZtWJUTz6ZU455BsTweQF3WJviks5+Wp8ofbrWHdAjyN19LQPCHkca0gM9k
jOq6tdBAKLz+NDzrcsarAY1n3J8CmW5T6TFC72Oig0bdRuTlIkfvJvEcu3YiO2Bs
PXmFpMDI3pNWm1/iE5SVkePdI7O0RwQBMlHMFuHUgNif+7lVXrsE4ZBnIgE/+/y5
imvZPV83dlzJuWlMnqkKqcdYc/KShS8e1ZccmfSzXProeJCJbfNrpxfV8+h5KXbY
1qqSXUvINYGyjeZ42CpSpjgMdh9MAkZ/blKqrSz2knbQ2vvRW2N6QSc265VLm8tx
B0GYrog+oe8Rvf8TiRE2njuINTESxy8vRYGm2OoiRborMeVrt7mN7uhDWSxNzIAz
FIIIWsObZIUCUPFzgsrcwCrQSH+5i1Z0/gFWX6Qrc5dQVrvyPcOzJA71/UyBRHIq
/tD0UgO+VPu0Q1TFFJDWs08jGdyNrX+Ar9j1iUT2kXrSD0cyT64PUPKbMMscohlA
4n20Elr21CLRD5LTXnGiF+rBpomc1i6RbvIZpH95VoSul9Amk3xP0kuvYk7Uk/lr
GmmSKrc8WAwCbExpsTHFofT+LUuX6j0kWOWcM2lTFwTZ+uaJaNukuR1kEG38g7jk
rNXfyKpsA+h4npBJUV61RSNWwWl9JYtBjcAJg1PT7ClA27zYqKuJQe999sphKNpG
6eLxub34Otsok1immUH16uHLJIGmnoI8WSjSAs2vkWNqoYxF9KS52zXYbQQ1yYSF
zw885J8mbtzRT4eqYQKS4LPc/7bl25xt+1hx6MqZQvao4LmjMshvCm8fz5CTJjhq
u2Cec6QQYMKxmpsW9YKyrQXsd5YmAGzJxAgoxp+1R78xrxCKwOU3qOhMisheHyY6
0aFrggPwDMM/sWhgKt37IlUwdsv/YjTTEmjS79B2Uc/0tVQiLCnnPes9u9o2RZk6
X8GfkswPHuY4WjTv4Uliz9/c/dDcxUeP6QDptrvUzKPElzwpDzSXQIzmvEJsEjYp
Yt8btqrVpohIa+b6lN9LzWTXCNXRXLzTBai3ahN++H+w4l8mXtwIx9/cer81m+Tk
fNXFoW59Rb9cZKl7Rfm1cSLWh1QUlYndf4K9XbsmUNukRqYdpW1zjKNkGvIGhgFa
+aClWYbJHIUScqmIhgM8xBSHKbKaGkJwWwUK2v1z1wQa88PWsoboqM/puk6wRmub
8Dv8Zf3q/vjHFF4MJkOdGGdys+4Ap+QzFbcc7ESwOH6qPUOrgKeNIXMmkwd9CsFz
xV+1OLyQXclq4XhO+7sESD3B1t4ZRrXTWDRpd2gTGJ+j2LbHqNTerGL9Ryb2TkKZ
bKHZX4IGfbsm08sw1nJjXlfZBbtZBN+yf0+AGYWokA0Ancfj3AgeInwsZk1ueaV9
PlYrtfTCLP9emBAKN2cvBOqEvsuvkM0O6XDCKkejUVc3zotz7HoMskWSSwGtDlM3
Kn1n6PQ4ZMiV56uxchLhtlPTWNRHC3AI7rHiztn1WlKBOJ7PWH2kpsPffR3sx6g+
BnihcKgKqgvTscHAjS7JgVOQZm1xNfD2GyeXqeM/bHkqYngjLLZVclhayHFUHsce
3frXF/uvXku45zBX2DXQYy2w0t6ujQZ/86cyV2TFfvb5PhEVagG+0rE48hicMq2s
TyiVyrPJhJbNcsq8ZPtuU/y+GHTsEiE8Kun4OYtXzggQ7Al5jLFIfmHPEyGijzbK
RWTNiiGPaP+m0o9ny6C1llU9tkLFnk/B8YLDLNjxWX1SXeNDNhxdI6xlAD0/N9IZ
xEEeYwqu36lNlElBYpuYrYmjUyebCvA8D7ZoaRow6O1xl11a4o6Yzl7yZg319SGb
0pNoANTty5gwASGETvLAx9kqi1qxExODXheYccydFk47AHXyv6bEa0pkwBJWneD5
qEMl6ewUPUVG7jVThkEMsaMXnFyetM5nJ3C2o1pltIESe3rLgQEBAfEtOWjzc4wH
0BXjC02gXoC0M9U2IhK6a02JutVPsUBQ88OAKqL0+cufBEt0cXsAaUsYIMlHmLfD
N+nltr74hCAoktZAfv058bnACQWbprZHC9Qe4y2/nKmTESpWaOj4S7WNs33qaJdy
Lx6nRsut2hoMqHeQoCvMoOJFXAUxHjKFpWTiVNqIfVnXVEoy34daGWgG1Q893DB+
oCo5GPJP6KVA5yKejnuIsHNMscbTloCpeUxDgrGj8kjWrdQ69xNPNZqOOdjg5/qv
sYCg2lpWygJhRLsOl4+hgllgEchAWe0z1G0L2y0h6byyCp6xwrUITSK1/LCZkGdJ
dDiJ5vlKJMX8/OGBp6DcMzqsjN6K33hln7EJ8f5lFkXw8PR5y/CJ8lj1UU73n8Cd
aeMfXJuYz2IDxZB+v37wajbwnD8LA8V8Uf5P/CDahiZpYMqtw1En4tiNGlcmv+lg
QKxrT4/75jDPkxCeyEyT2NlUDoGzklm0QoVLwgOhxgd2J3Vw6i0waWIU1T544DUl
uYO85ZLzZPcQ+ozO6JlowU1bYY1/YDOd+Pr5ZgqY6h/FO+qQi0uODHBJb2PKPOg4
tS/KMrIPE/es0h0yMgyicVUtOLYueez7BP+azboQq4C9Y4jHiI6fKkqpRmvhdaqu
YOsjTdrfsqdZ2pbypE9C+QimF095JgDYI6QP6CepZsRofwby9iEOW+8PpxFp+uVq
1g0bDteBdS4YW4Kn73fad3wZw4o3HXV6LuJ1BQIrMgUOZLJUJfiCUkAH9WGriHvJ
CPd3uZUr/yeUixyh5hLp+E3DTt2j7b+OF+Ya667FzqUOzROHCKmgoMyJ52xBMkwO
p2LcNKUJ+bnWX0A23UWB7yNlVwvMlXCAyRf75f37kkRlhSPzwrAat6EuNcz59v8p
MIss6oWFzD4OM5mhij+xENCp5vc25yKjZVhjfrVnJ5MoMwii64yYmnag7pHvEpK0
cL1vwXvrtzQtTnnGEW5nzGCdpOpvnZV0RHMKeaIBHW2Rj74O413UWHBB5JKfdgho
1WrIa0blPmsob6NQ1Jj/RodgpaMO3EIEWuyt2RA6QJ7QpNCS/Qg3rxaAkaTQ3ywh
95D+uKILAx1RhOLzbmDD0RPR9CXJq2FbvSVYxCbIEm5e0RuRHI7HxPjK5WwrqXgg
O3oggKlbd+JoSBxe8IaNZzlrUU2FFnHA0h8gqBU0dfHxKvgVmmwTp2G2jq5USMY4
WNTkOJxev4qek8DmCFQEzozdWagwBASWRDL3nNwdJCXwnmo9EvfJpuZZXykIj2vq
S0K0hpjX7WOjdFiwMi6vGOrwi4wIKc4XydUkpWlnp/hjoz9oBYHKYFSeCOmhYGVT
gbN+8cD6uWTiyRV5Lfn9Af9X/EXzGXyUnrP/BFKnDjo5/jCCLRFgNbFpeKbHAWit
m9OWZtD50JcUvpzao8D5ox746SnnGi2t3MxTQ7en2aWTZTkzkvPyC7s+JSkASzHH
jJRn6JLJcDpzRL3CK5rgNkATYb+NbX6eDW+KJ4kSzl5Tjhu/Eon/4Vw1HyVv1onz
6E/GaWMZkH4Yb7tzwuYII5szwrfGlr3R3/HhMl8sEpCme1DPsgAk1JCbY4/kIeJx
7ar12oVh76YAQlgpMK6yJzbEMqOPhnYunC7tkwDJ7o/WYMpfmoIK1vrQOPLrACMZ
9AvS1LEK90sWp2Ty25SoTyCvwoyG+CAfz+4OPmFoRDMgwK+saI/Qx6ZzqzpPdYsm
C2pO/5ZsXP6K8wJzOYe9R+m9kayGQDgiGVldIkTXUZ+IhUE0u0Q7TnVbHhak9UW7
9AHJycYcTNDzkPkjmMR5CQou04pfe4RoRQ52fPM4cmPS6CXGYhc/jzk90fyVTgWw
ZmLUMDYc1XdiEEU8cISz1XyLIB4zeRoMNwvHWTHk+SQ6UwRRydCumCVvnRaThlfN
9/mRaGVuGvL+3+FOIh/5yrytD7Kn0IjR5IyYctYBpFInCF0N0EWy3cZmPbY9grO+
yNoGTQIe1gIZ0jgNQqPaWibeQVLyp38a+csyOuvgIXFtjh3PJN+bKWP7aqrO4Aob
UCScbnOQCjkFm8bJCQ2PjVxwhl80SrkDdC+9E4mu1agzlAYlMoPnlbAeev58xxPr
t5XhfReK2DajKkJsgvWiDbkuVgCzyalD0ZB/PefVvXqK5KFoC+El2hR2nIyImq+E
qsGHd5FLqzt6vSjaD3kDX/h2XhTfLq0pENeTW/Uwvwto1xSCPZfp10c8uysI9KeB
OsIYUFchWtL/SUt+vO6G41pS1o/V/QLWuOohoHJg+crGi/AUOTPknszYppAi+GPZ
FYDUTCW1WR/Vic0wsuuce1DEZXHPX3hSGtm/r6/Rtp+NcEulBvj3YJip+bSrBNRf
TUFp2BDsZML72oP816m9h/3AeTX/MydsDNoUWjS9688+37M2hKa2Rq5+PW5y3jI3
7Xf4dVPMHOTr9SqZTHL8lMuqQqpegM2eUafgHz2zIvebXjEV29mPtIJWYEPr761z
+DKEExDhiOP2LlBxoWU8sE0ROBFLmV0yFyNbS0lmqvXYmLa6j6/FVaJtR2WNn/ba
8LsOgLnxEHiZ2hKLF/dvp/rf2em8s09JTF1Um1w4xKk3iATGkJVsd4hQw9xCf+Vx
P4QWK5CvSfS5SnY0k2zKYuCFfH4T/a6OecxldKKMGMbuiY7YHE0p9buOyW84ICeI
DNfYVsKC1pRPCrb6XJST5WSdYZimVRgen2ONlOXT0iH0L5ZtMeDSqkYW9JzEftUn
p6UB0fg6Ye28bMiab3RiFSpdeKBQausYQAwxVcrXgZzCqf4ZMJmYeTOpfs3pfQSd
wBif2FLbshVM9S+yV27JIvUdufcHj9lkuTH4MHfamNeOR0WIJqMolqhJoP87ezCb
sAVrJQc2IxIqJmT0lpKPg9tl3uqZ34V/JzX4UWI6XyFV+215z/i0t5g4G0XKgY/3
/2PGm43m+8W5tJ14IEvuxnnUjgJsHwXSiijxAYnAsE9dbcPSaQdDt7gQ+pNwmMwz
cT2XMGwEaS8xHJ9cGPwxouSL7vqNIf79qAt2NiUEkF+eTaYLfUjkNOrEHc9Or/V1
ozNYwG1fgGF4nLBIvlUht4UewOiti0WlxYgHxRgbb1JlwYdc/OXPHGUGNZLfJWwB
Hxlw/ng8M+JBF1EyEWAA+M6WZuauJLHqSpkoznRV9mF4rMRFnswSKjDnARrS6cZk
BAuUXlVKEc1otY2UffFhXOYTjZjVEOq6X07SaqwTFmV2+ZUVofJX8LI+VJC1ttaJ
FUlpttd2V5gDsZBpjMhmzn1t1FXk7n4JovJIo2A2RBVpOQmCEf3YkXT9T0sZRMBY
74KVvKRyK/EaPo0Xeb8+gSJ0yiXmPKSHnJe8ZS0d7T3uMrT7nIRytqxFvjVMY4FD
+4iOnao3KLHjOVPdjiFjG+eSu+TJVu1sT+iIiZivZcptzBc5ByH8+ME/Ide79Z/w
LWmsDagLCm96UBonoOf/nlMRlUO0eZFpLbKXJ54Utl1jQLPSo97q/yRtn2i52JhV
nzk8+cO3PjVqpTiWfcrhVi/3Is2QBIq/kyZjY9r0eUKtnL0SPcSHzRTPTVtA62L9
ZdBPHghSrMYheWPRbLtjTG1wGNAfw823odF5Tp2LqVJJlQqaE6nBmzAoKn+m/jiB
a34YLYvrgGwiGZJnoF91wiBFbQSvXevuua8Y1Yq4NAPFVuU+NcKHv0cRo+yLByCl
2iA7uI2W1CWlF6X7N4Y/PKQ3JdcQJcYZ7oJKlFbxGS1oVOX/ATfbOMyM4Oq71vwP
dwscVFPkSwx4kc6tV9lYZdDCTVHcoFWopn44oUnfiWG7roxq7RzKhRCiRShlaxU4
GXkZr7lOJnIOERxBQLAhaymT5oDls5jCxO2lLMaN6B8kt267pYKgULL2eIBP5zkJ
LbpiKd73vdWeR6dBRKf6DdxSxg4uS0Sq6gmEcxHbfpCSHnt+Hg5Yg+G4GA6/zbA3
QpBz2cFzA664kvalaLr3k0x74kTKahnC+NusKOMB4FUoZSzwdPt5YuEvMPQZmG0D
3EmU0epOieTdcHRL6xE56Z0Xgrflyw2OiMWsdW+hmgXVQdRdLK12emANImpp1E6R
Dz+NN9ueMJW11HDZmEb+nAYzGhEwopgj/gRZgQmQhvwvCyLiI3HHv6P1m3N8hNEr
6UsFhQfvvOa3hY88X9/dVnCfSr6TA5pQ691aXdrzYxTlvV1OZxHj8L27ddsYo4oi
pMuh7B9FFxbO/lK7k0MqjZFhDGu/InMglV8xhH9TDie/6rCSlx16vOt+Ctck3eEZ
9+Fgg7vHot2nS4qXGKFMDEEg4rjrHt2mKDVY3QsgE5md8EDW1u93fZb6jksjbSoW
yTnVK1Lytlyuk1GJ3afBdK8PtAuYklLuk/cD5w09NW0JoTEXzAVDY9mNxKqZQkUA
8irJEex6IP7qstf+2v64dExEr4AVRtasLKadpCvLgiqczd2aDoHrYERDQsfvPn+m
sH065VWzqraRmQ9GEIU+PI3YbnNpi7ThBcpSQvA5dki/RZVM/kuo4n98Igr1ej+e
1Bj7Q2YhIvDbAP6ZHQZbgDJ4JznQYlb+8lQzpfQWEgFZobUbXa7EFVohZfgPthFL
SstiK0x8Kfq+vZ/BcZUPUsWm7pDg7lUYWgGhH4y3nK9YqnxnyJU5NQg07n/E3afM
jiIderq9W6A2v3ranMRbTEnuPppQvnKsX3hpjqoGDEiEIozggrtI846YfNs9xQ4y
ghqo3ah0CvAM3XGXXYyAonijYKS1+Uy27oPASZJC2s3j57HEqeELJ7SLu2RVKpCC
6uGjkOb1IwX+Ob2FTjKehgiv7VG7b8u0nlzNy4HpPu2lTcqZyKKyu28viZxzHAqY
Cx2odj5tmb/O+9gtGAwV0Gx1TGEnBHY3ibvza+8Yu/pILuNjS8sqneFplNaJqyxA
/Xu6JglXKmpmdkx5tUWgWFImIdE7JmTHl91r0FxLM62DhEro6S2EFecKMflcGNKH
47zkqugkiIAf3NN6cgBh/UR2gCAgHdyLQo/Mlf2H1XiVsNcF1563ZXNuoV4MgKpe
GXe+eAdBg9zXGRLSCLWTdB6Z7iZWQF2R1oLAz3z2SUt6owDtHils8Mz8dV9/GaiN
Rco0G61nX/h0sjKtyl1uO0UON7Z2o5ypgsY6p8jLuwJUaznTfcJBBnMd1ehVCNPP
RucDmsXoOGrGHHfvDtaW0g==
`pragma protect end_protected
