// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:37:13 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
J9XpgEMXBalILTf+aryQYgboqQcXAMcJxKH8+TgBiKzAZqiE7Z9+NMLnuY3T0Neu
MbCsj9eE4FPwtsDHLKPLgKL/88KtCblEkBcqvl2mugP4PvncuXzSFsc3SzH+rM5t
TUTBPn9P1jXo+sO9ZSzhA+4cvnZSgF+rzEKji91AUC4=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 3424)
2GWgDm2yCO8ackzDNzzuiO8NPh8TSiRdg/Zh/OYHCmIsrsUhDcZFIMQY1wiERCQF
AQ0/cCdjMe+IaTbu2+yAnuIOS0Q43KqM9StC1axnJAzbneWuUKdye3ul8MrT9qt+
mOpJktc/0L5AE9d7thIyBKh3OHmrwWMXNYzmjJRGzvOH/PHaJdy1g6nU2DnfABVr
GS/3sG+1cZRatCk2HP0i7Gl1HtHF0Gugp+v+jxv8wMExFSyukXCMm3RCop0zhaZU
XKeSmcSLJcbhAHCKNBVSdUwLXe9Vm6/vo38s/D1sk3ms7g5tVvGC3W16mYZ0Dbj5
hndDU+k0iXpDXv1sYGkC0iXhpU/BALAaYdkrU/tCkl4hd5AUQ+OXtk7VCuA22y2d
OYF+9or4Bxi1klxTK7KLLEKZTg3rW081RH/gy50d31Z0qS2+jrPWcUxQVWOrVaRx
76VS3le2otIDbNJxmkZQkhPdldWvd3CPVqNp2LD/Dn2LaLDdSJ6Q/zjcvFiSNJjc
qh6kOVFbaxWi7uzisEz84FPabaQut0tjJxX87EPw6Hk0CZ6F+8NzYtTecBFso+MJ
wq6NIwnzzd/VOKcAsCkfE0KdVWQ+CiiOUQ1Wec4u2HB30rf7P+tdFcA6Swhr64dv
DJYhfX0rQZoW8fuM1yNzeUFupip9+CtA3mrxCqMxQmII29q4xawcnAXbCD2D1AQV
qlSgt1uNS1lTytSZkRrDeib8115n58ooIqU7F+j6ax3CU8OhjB56bzuqMc6ukjGp
uEwEIGeswIiLXiM64Ohm0BKEU5CS6OEuB+IkSnwdWwvqXVFq8bIVqM3092gdQRfn
PGL/KaiKfDksd0PwyDD151UpbSNWXIsmIS4b/dZj/da/c/wQs8+fO5ijWe6QtdcH
vbRYS19hTkCGvY379GyGI1L0cBlH8MeSQkZthgVcnFWboaNjRGkaeOvG14KgOlI9
ovVERnqp0F9cs/Y0Rial1RUWqSjbCIAb7lHi48+w8m1V0WkwgFKmPD0xJkhTIkVR
uBiX4ErwQhbUIFk7JWScVidjtZErCVYdULNRWDt/PA9MltzGRO7o8iuBCTNEi9Na
kfOkBJVp+kitzJKcfuxmTGQ+kT8LFCvK0cGr7L4SRWCXk+wdNPBKMqw6NApx2BWG
0W1AtAYq4dF0iKzxwwevTAttj3XmNh+jN6pDlZkfmN9sGdj/6M+38poNYDmZv0kk
+EepscOvPCpZeZLV8OArz1TFjNKXDv/xI5bwqDGgg43e7yRdRctyiCqvmP2HKTku
gYUdFavksXeEufmu6Fc4Op9FXjvOZ9VzOmK/HNkvLCbnnxALrQcIQ68Aoeg+22EJ
8NmmbNjMlNweqxyrUJWMAApIT/9Pn0bnAZX0dvRcFrpC7rpRvs7+XWsJkMyDAC43
P+Rc8YJprp5thkKpib1UpJWbqmWp4MFgf2YJqqcPCEcwphYeruJAi7+K/7NqoKDp
lzT/MSnSB3R7pLQvNhgJJ6ioRH4kevUpCnhs35GAiXeNoN0L8X/Viu5nDfy4DHg6
jjHuyaL8O50LsJ3jVKY7vBQ44HZhMYcGTnVv1An1qzaRvrb/53tELqfJZUmFtE7V
kUh9cI/xf3KtajgXuuX6Am3U558V1TDOXfjRW43X94vB7Jw5+esw0pzOHuCVtTFT
sYvVl/m4xASOKK8Ab5/N2nZErv9EEB49EBOyn6lyNpU+zVT+xLmhxv50iAMUjq9t
MTzhpGr5pQhSPC9uo4iMnzIIgguiL+pilnxFzc6NAjmNcPNcugL6vQgK/X7V2+l5
MLoF0nFMoinCIEZw+gw2cuzcXh0IW3qLXYZA+c1n0t0XkHTvOYXRISeSPIb6rmp5
IOnUpoVWmHpVkaevJEdnCsD8yofEzh1CHiBXFL9WjyvNC3Bpj+hWfyQtIYPlJ2M+
pxXWXf88ARMb98zD3o6ls7BJSSnrWW0tqeBgyCjrJuX1wYwB/IcjxcllaXrTvI/J
axfRCHIoDkaJk57gumEspbZSR8U9Ia07UWm6ihMRQc62/Tnl8i/OuQJ99U5PX7bE
PY4x+wh1OpvxIiQmJTyFQAK2aT0f+W/n+9UoTnK0OtogVbdDaO7AnBT+TveROgnL
F9DSKuQ5yU6Tgb3BDNGO2TL/X16r3ZkLW0Qaoe8STQq6qYOuZWsCA/TehsBxCcKP
Vsg6wWQQN3/ggL0sw3ygqOeTkktVMbXKZaj5u6ny5xEgNfEO+qUdrAdR0foZkyoC
4382YS1PKv8f795TvsR5JscFYVSOfbSchPAwbRJxtv+fsnIIWuhMsys5A7/KAV8b
aRPWZ80u04vK/KQPxauhPBBTxQNNaXHP1BOmUYHIXFppiyb/WUHOXJuEtQ3ZeRpk
QvV/rOGNliT4iiNKCea8zLyhdQHIoLt2iGbmHlu2SFY9I5EROTI9IZ2gSGeWy2UU
PW4vISqKVmZay/Iutw4psvbtqHTCGIih6q6zbdcigU82qC6yaTnC+bnCwEfyKbxv
4ogkTIoXT012pCnhJ8vuulUenHzgI7sjccFHKGnp9d4wNm9W0xys/8pIL2SH1Uuq
kbr6TPsU610ImL20gRx5F/7rmcg06hUbP+pUan29oY8X/Qfq2Ci47PkSsEDVApGs
FvZxWgjVAHa5Z91FEOb17qBrY9KSaEETFCluK3zWl/0vCRp3bkKvQz8xG6xDmcrU
mrqWSzVg5h7C/Ayn9kwr7czCrPhKOhydxv0XtKgAZo7IDMnQlIOAZA82AlEmSYyn
9ni6GbIP/9mKbTvTsL8m/VHnrvSRS7DraTZnB21OJ0H1h8A5q5fPc56cNQjtVL1J
qjGqBiNYasl7R0XUf9wdbNdZ3PVEXAA4ukaYWBnf2xjtZt4o3Xo92CiwPwtdAmjY
xwW0T/TLWboDUZ/y6yrzo5SRW+Jvu6W+lDolf4IfOCRUQkRNoGKv4NJfZWcO7Pc8
R7qRD/Y1k2qzTz/6SsIZj52hc40pCvhbzAinBG80WrEiF/oaMfiRwBLQqzWcWHwf
CuWbb7sx2tq5SkEcMa4ZNJTUzE4aOYSwZRuG3cvlh5mqB2FD896+faVd9QdWfLXE
AAT7+UpKCWdR6/Y/xNn8MKmguzf3MowaF0k6ZDZyN3B0D/tjQSfolTwmwT8qkzUu
AOz31KW7hDYd2WiWVlecWZiNHSGnM09TdYkt2kdmhxdDrLl5g7OymrSQ9iUri+/K
8w951b2R2bSFwugo1SkXYCvsYUVEzpQSTWWoaaNJ2UHMDv3CeqhbLSKYxCOpJlEF
cowpw9r0dR0ORUop0+PDwmPvDLqtusQVPEEM/3ArqfZNPSOgxnI9rOjeOBb/sXYM
lGsC7VXNRiic3oIzYdwQX4L3kS0sSRa26rALEeCaqnlkyY5f1J3wM7jWSJo0c1p2
/5rcmwFNBof63ikWz+j4w/o1sIcBvP6NM4q4DhXitvgT76HJAXQDlq+xObwv6ILl
P7Ww/T4Bsfe3ABfXUvQ9lIwn36htJ0Zz/Kb4tC2bD3nsro/uhEVnf8wqVsZWH2Hn
O5XBv0zNCwFkyY5GOCINWU2m0l7wgHJEQGejE4upFqef4khV+M1tPvVVE2dXSMyG
K9QthpkArs7i0x2vXluXzT594A8deJaGmPV62hEuMw1HnCwbwhnhF2EaCqgmQzEm
JXg6UNOy42E9ldHCDg8gvWee5EG/lPt/OVv6ipkQSxQPXl6I65mw4nQ4Nf19L3sa
lduvgxy8B2vOvNXM0I5Q7VMwS3MfghEv3Pe4PtxhKPqk9Pos+p98Wj5AL5tFKJ3I
PSvPVSUTxjCJz8CRc43Wc0EQMsrkWrs8UiTtzcUWJ6LHz7ae6JHKLwKtXlx4TZcS
Qqbnn31kEWwzo+UYHfTgRz0PZ/Hf6oEWO/9ED4Rgug+JOakQN/soItrSUp4pr9Ny
WEhlxIIkV/ExQQBBhnt5OGeq4Lb/ChJmer9aq7WRhpJj7gKe0qYoyGWTfaWH/L7/
1xjnqmw6fzI5E7GnZI/OVm1iA4OtmsagK+hwaZddjVgcjUtZnunoiduk+gutsai5
OE1JtBDH1alNYFv8Bt8h2N0WdNIWY/VhcIFLgxmoPGAFI8Efv9jFUpxTvb4PQ0fD
Fbd/CVbRfr3CqNYTMr23T6hdsSyzR/RKB2+YLbKdCth8NBGZRlrV6vW8j+ip2fpl
XvRoa1KicllJHaKqszn5c+bhqjNwadlui9DFefvcesadzVx8dKusJbZwoR/oRZVl
pb90LqG1eiRdOQ0JCaSpXzNlPg3KvHWAwzieeByUz3QJYGn4B7RuEevRAIKhS9sL
8t0MdQOeKGkSEZ8QcmXev8WzmwQsLU6sJ+wcl3pghhuAp4f0F2e/IaSGLpeqGsaN
bu+0LJi0OnZ1dspw7VYI/OZg0bMj5uTJAg+jAvIj9/v2CSbtAFYlGE5QhgSUOfQu
4RE5U0vQ0dwcnUXpbBqV30Br7DwfBRASA47k9RrewiscMVBUE7cNLWC3pXbhsZBQ
oOtHoINrTDH0TcIxgCI25q4nzl2kdzFTBKGqVezRWN/TmEohtLyPVLu65ySa6pwf
3BqLHK+5f0BEdGJt22ffdw==
`pragma protect end_protected
