// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:37:05 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
YH2IGo0qv//gczPTbyVpOCTyl6hgvCnBxknkPFOen9cf86/eCpqia5yDIIJEE1Hc
pWB8iHr/a9aLOJNh+409yvKJiuCSRlYFlR7+zhaVXmB46t38p499yvJS+s5FhEfb
bbXpK26wS9nsqfVCKaFWWVgVgDX8yt8sk7z7Kg/JjeQ=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 25696)
cZtcibZ6QBsuaRNj/Md/Bj/M95sADUMC6m+prRk8Cy7u3jSBZHDVJcK6TpTsy2qZ
6+YpK7gn52V7ghnfqGKw+kGxJAogsAZd35i0CBf46aOhhFCQWprwTY6tHFl46RSo
uGk4N9yavqorQFlTaYQzqBrnPyX+JAlnN49S7EzktpwJ58e/gYcUj+nCbed36nWK
+oaEUSv1Ib9fhMHi9jOTOv33T9ZRpRF6f0fC9kbTvBNpZDxcUNFVwJgGOESbXM1r
OIsMfu26QGbJZZDEUx+a2DrEAqoNWlrHyWvLZHWRdmgtilGUvAB8AS4/SoY7uILI
OEnFEAxGAjFmny31erB4NZVhCtvwOBbU0Y8c8VqSsQ2CVO59ez72TRNf5wufVI67
G0L21Hy9yTEQYx46N3yBXXndK9nWXrWax07svuck3D/ggPcSE/QVO4Fcm+1zgnVH
wU6miZ92cDhVZhGe2vitAHYX5ax92o8zix5sFBPvQdKv4xfp+YCvrPW/Jq/hlD0k
h1NkNEG120Kb1FUvYURK4D2zEi4/CLav+B4jPPMxoowtm/S9fNeuRj+luRAFtLzW
IIRbPx+DqO1bRA/ws7bThzqyCYbFgLye/QCo4ZNILZmA/tK14cVboxPKHdUppXc+
bden//rlXQ8QGLLwdyonfkHNpL1WsP5oJK/y+mX3N3s2KTyPNgpamw/zxzywJvTo
uGJqp2OtukqU8OP+uWqsOjCo5FPSukqBQxrabtLyBb3RNDiUCwee29nRWezvJ3//
GsJDj1LI2jjsWmRltpum+fGu5Z48qlNKNWv/KLqIaA8B3a2+4SA/+BaM19vrkmSs
4d8fnM00fW8SEmn3oQrQq5w8IWy153g757WMJYvFnynJRe7VHuP/EhnP49d2D+Pc
Y5lrGXhF8Wv3SgD+PDVKEMSfqFQfYgl+oWZO6TDBO9LP3koTIeoIwfNf4hdCzw2A
ATHnMjxFXIB9atf0nx/lTupc2FM1cNiFXRiqTdaQ07iueh9BjJGtmfvpv9d/skyu
KEQWfrAlD3Q8kWft4vVyqkqsb6wLF0B72kIgke/r4aD3UyzbZE921bKxeum7qX5S
CUpK2866RQ1+wm8EZu7ij0qd9TOvlPqx4DkzgLGrIa3rCHuhaDQ0G6kM1I62uwK0
Z0EyIuIdgqvbwCwDaVtPMCigIzNGmDGQDkFoHC/EGGIvANalIwGjpshiOKozJnAo
1zivJIHg2/NYSuoU9H4bAvCdQop5OGCF/eSTGRfwjK8cC3R9Pz4oj8rL7c3IX0li
hS6G6AmuRMz1Nd5BuGNOW/qRtlIrAbf+DFsPmJDp3bHWZgdc8yUeQoYgkRCkHjz/
Vu+URUeXZIk1cFzzTI/T/eObttiHcAIyCP5W0ugMeUl8qVf/eoK/cqNGqRjQoSh9
zkXaDACBbDfRzqQ9IjoxQiJW5eSHDXCQlgDCMVyRdNFvtzc8vvKtFgx67c3vTUkb
gNpmov2m0cKC6bGrd2Y6jaSbNSv0T4jEU7lquUU5YIH7jqYiHw2ITzZNNZYOeqLH
sryw4zs4nAeS7Jmot89R+7Funs48pRrD1YXzaaq9w5OKnvcbdzw/LqcWdfKJv4uR
YkaKTx6vQGYOF+klWJgOgT/PKDM+ev1zdBdUjNx7gTiKQu2eVKpdD3gD3BVPnK7x
8g9cxhNYjwrAKQKgjArUo6vYK83/qJ/21pBhrQSskd5bJ681O6MY3KO++4HYKKCh
B+g1Hmm54yho1qR9sys3BoP+omiInzvdyu8POFHkK03zOlKaqZQBX2a5KMFsBA8G
XMUfeQPs1HwumJxdO9fwpM73pZGTtmnF7k04OO6R7dPGIC+TtNsmWrFRzPmIM7PF
Zn9WxVB5LI59gh40FLyK/To385FGa+SJZjelORGcssbi5tBv3Q5KhQxOrbXV+54M
CptTMRVdyk1tzUSDcR+E4opRQFKpbd9R4jU95EjHtHUJklca8HYeILEMJWvmqUdJ
YtGI2yex2YNO0PVYF/hP+FHEoOfEo1WCrjMoAo8LK4cg3CT9tlMbq5GI2gl53rLO
ruJycN1zaxfR1byAxbYTMyqckJgtP6yox2OArF+bcD7mkob/qbXWFxNuOxNzoPb5
IZ+rwS2E+dR2dMtGhrvNTOOqvPrsS7/lkdm+M+Kpz0LKdG8aSn0oVd17Kov/Xi1d
5jElao0t9SYojkisnK+XafHYPPNhcS10YEOPJ/43OXzQ1UcJf8cu5VNM/3Us1rqR
igeeIF4yFG06DchYbG4Hv5IwifGfaDYhXAXvdAF+V+YCn/+CV7m/XxrwZ1oJUn4i
b6RbYxz1bwNGesOz5kb3eCmKey6gLsck1CbmXEQnDMU869opWTaD5OBtzDl5ZGhS
DXWWKqt0L4SrV0WLdBMskZ8fOj+E39Qe7yCQzWAJ+uI6V2GTHTnzsIHux/a1yeny
PExiFAB3D8rskAxEN2rzdvH1NVOu2r8dFF10G3uCu15SZIoM9Ofl8/86AnoX9y//
9upK1mH1l28jO0A3MvX5hpKibFxqq4RTAFPAhlN5lyvqpCscGXuVrtKVXcU9qp/D
6uAdkEeO+idMjW59EJmHeG0kLRyWiJir+Z/ZuWXkxneaoIfZmeEzY+vd7wrZSTYA
whlg1uU/HqmVyRHoSRUzYext0b8Rh8Hc2hSiuAQXjqRmCysKh3hVjfgDlBA/+dqh
bf6aM0zE6C4yRL3WO64DMyXxMvu4VwqMAGpzuh0uUD30oypgGS5Z3sVZTDYKXHEF
Zz5yotu+Z9tBzwscMA4ffybiIccBfCM8iUOUODDhXyw0skFRArTvlksIKQatHRYs
cPYWugh28dJCjxM9YHmmI5HBDSAjMdmUBnRU4UqNsXwyTT0wvhPy7m7ZqhQOlTj1
QqJCfqesBFyHLA/YocI6MqikcP4uMwT9F2rOvdw+kSNwpyxJPZesfRnxVBDDlxHE
idMA24zpr1ka16HjFrM9O5Xq1ZFviuJwo4/3sFQfi+3KaY0zmuqzBYpLn+N7Hcy5
QJoOMuPPdFJElL+zj6T7ud2iMlIH/N6gVHiwNL2TZ97aa4n4hTnxpkzmSHncVL1m
kIePmx8eJKBBWfFQvOMosDhJ6N1mrd6F7FxG03E0pyFw+v5zt+1iJBL0XQphWuKR
LqU9g53LRET6Klh8Sk01jQRSnXXphobb6PNYSPaAISqVLgY66y0TX5Niyq9wuTOm
IXqQskb/8H2FxBXDZ06G7LyGB/UnCxLWARhlzGFJ3oEc3o0W1IwMKXEeAHh6vXZW
Y1OcnQSK+ESHvZ3v0e0MYwbgL5hpr9aWwlLLAz5WnAdXvdmJ653XibX4dMsL/6b0
6chvxeKwhw+MRgembZQXPWdhiMQDnrhHecZBOvecM2Jy3WSZePuLR/nJ0LJtVgAN
p19tB7aSeqkn6QUd8VjpgqewIwliZ5gqOTx31xjX3AkO3nwmkBMyw/UOJwmyEyh+
QLLjyOViFbRdhq9q9RsCMrYC6NvDoUPfy1xtMGi3RND9IeoyvW6iDIYm/cHAR38f
fqdGNIhCpm3MKpAVw6q7TY9lug0obF3gnfg8z7J33xPnuQ6EuX/8SpU3o/NJjTrK
PHCIkdiOIduzs9VtKgKNEpPgG4Lotmq3hpUWmRocXNvJplLVgwuKNI6yrLKs+RC+
zuKLYgFyhY+0bKuuj73GinXltPljP4OHRH8ecJ8htWTNM6VMpI2HbPswVhHTPOsR
rc1bvihg34n4vNjQ8YNUDmOkTyb5DxUQkZ4u/dCR58ihMmgdkyOojC9lsQLL/f/Z
T7JdnmOUe57cx9POkeNXWHa0LqR42oKFv/v4J5HMAi64Do+ozaz5p2xAnTRWZLzp
4ifAa5aBQkyO1TYqH5hfOPh2LkDNtB9tLMqJ+inuPsnxiobeihu8x3B8rsESLQNn
xadbtYn3Q6H54y+efrjjCKnW9Muy4jOVO0NUknRtUNBbtuanv2mXa7vrAS7Zqe6/
aAjQoc35a8Uw8vI2nY67Jx+wzfkua7v6+Bit1PNH3n03sTzIszWKjSghlSSHcxnC
3ZNVa0OoXFs2ikjMLCrS7O3TwmEcn5TMj3UZBPBmf0tr9WXa04+imAwb4DHX9kjj
ZbEaFelBy+4DuOmVRvqZ96uYZjlKRVytyyumTw3IAureys3ohMOklkLnxpxU7uSI
RU6cnaEKrkOiXUUgq0y1HmX3Em6mIYoA5ITKGAVCQGcIv8SAW591b1Z+TtsgrhnI
khvjXYK45BJmG85DfpJmgTm7/OVylFqlqHQlcRDscc3ZOk3MjF55Hch8Cz9qZKNl
hR+Z2OZRHTcDtPuK+iYTQqOYUiiPnBJjYWXx65D1vF53zOkRykHXSbDtEt/sNmhQ
XK7M3RuKVP6K1T6SJNLzB7pXEHyHMbT0FGPQiSgfjw2KEDspUMIpwZ9ZmNbm9Sc+
OduRESZPny13jRIEXneV0ffwoGAvD+WPEBHl5c5TJpJl2YTqEZmwfuPBV9tmWhJ8
EpN9K6BZNYAODTJkbMiRErF1Bjey6Rpyr33hPFOATp+37qdWJXys4QkEhXYYjS32
HUH+9gAnGvpaEqZcr4QUjSAiurEUqZVgJA6z3f9joDD7SGoZoAd6nHgf5R8EgQg2
SbHXp29zQW2yj/y6JtXfG2g7KzcfyUpFPyMlRE9+EKTP8HgRjRfo1EYdd1Ioapjd
U5cKfPcIuH13Zf2ojX+sK1sZCf8leSfWy+ogjIyLfKmdhIdAA1UKaAbURTc3/9tB
V500M5V7xZUm/+EqZ1VriAEDl3KR6TcNrtVlgyspAPY7DKtOoG8WW5g2GZkwRyfM
gIResrrxixnEKGxFvmIMea38netQbyQ6lrWfCK1hqPe30DnaufXMzRFzOUUd4RAQ
kDARcTioamWINaKvsACwZgjIdUZ/UYezTkk1PRT8DfvEbFF8Z956rqeAX6wFomde
2oCByb6FX1aTv+497aX7mbSWh0TENyPlCNMk1zA04DU2ERwXPKmKdUXCe9dkXZl0
f4JM72CnmLek1lU/I4pqGlX01IfbbvsV61MIkZgrGm3a9Zr1KUzoHOWy6F+FJN9J
rdjfkik8erKT+QJdYK+v5s/ACwOFoLVzVUI9D6VslF8nv7zBzSrx/+HulzD2iU5S
JCP9K37Lnpe3MnW4NyNnmKNpljznR8ZZc+YFeJaSG8ZuH6r5frLUfErtRLesAlbc
7i3BYn6nAYTKWr5wCmsJi69ZRg5sP0ovio/6m913QwAC6J8uvsKXnYLG2zG3k7y5
EY3+1kInLDzszUYqg7R56XAwVCgaCCxRYegttr9pLRowNUZmDmur5qtnlW4LCsQE
4OSEiHZDpr+PQXZYWCDFPFY9ppGUVu776nDWBHASq/iSNZTK//nRLjDwc7nxG+v+
R34Mu3v9BCMmqtSXWQx/0eluxfyXBq/G1Tqc9rs7UaJybu6U8IMWDgt8nEw7jtDI
sPgARkeAUembCLHDMLjcTqbdIsXQa4GLnR9LZsTMb3MBxVF3kWYAPsYp2CRJ7YRg
2EgymDSAtsfndJ8LvLQnD4itcSQtp89mwEnva+WhIptUt78/jyR41Xl1XKVCm2/g
rrXElAumHNblWjdCzoflLrulcSweiou95JIZ12hIqIvlGI/7M3+7nFKrZRHqKR33
3AbgQ59wrAL8RuH0B+lOzfKAXAXOFqO4bdsY73mf6VIhyo9z3gyRdPCx+MWw6AeM
lHH0iirCgPsKpRCkpxVMEMekFqhfse4D8EarL9bT25/91sgcSqj/ju5Jr5sX6IpY
Pseq2ThyTWskjExZbPuhZBSBpa24GeycH3CXiM3/5UU4nln8Y5yWjsXyH04E06iS
CjK8YnLgxq0Kz4cZy+RriaPOMylz8W7Tix0zkt9kr+gUYOFGaL4P5D+B5RDWqNfh
dzZuhpsoR5g6+vJfkIj5CYJuo68VCHG2NCKoBFGCwjkkKT81wCgc9h/xpW/2AvV1
mm8ISES6ZcvN9jzqCRoCYIuZkPTosE6FQcdto/6l7jT3PEVVG2vN4WM5stYyu3p1
fDWxtk+th4CpOU8cOK2teRji9OuEYkEfwVqoH1GDegJ7LE9wb0TaPOpUrLDRCrgn
h3qQNiS7OT+EwYICJbe0tCFITm5TBpf+ZtgxWKl1AQMfA+Ic1nETYJZ803B9LEX/
oqvY/4wk0M+yQeT/o4op8G74zLYGXrHA0XE1LhiDC2Abz6TSmpTeSfAZU5En4Tq6
0TFNp4yVN7ZBLCBI4F6+1eRd4Kv9ci/cYLnUvifuv7jkogmzzTFOLgNERXz8FjoV
tlc1pTReRsipVIHQbv22OUVAD8WgFgI46tmhYAc6djCkoOL6OOLI/72CN/zbep06
DAQDRVxnz87dxH4LI+DUC87f1sCY8oA29ukfNSGRXAxLFqO2gFaWHpaogphTTyq1
agUQBZZKk3j76fcj88fDANHf06wg5H4ZgyCXLNYTkcBcm1//VQCnZaWOJuyWHs7b
pBblLRmiyKZVy35tDJdG4WcwQQbZkULMHv5akX1UPf4iqL/w8X6aSClQ0BAlmi0k
+7/ZIkXDT4iFwWsdPiFKGcVr89vttFNFPaT5+kzoQLNS8PCI8Y7reerYlt8pEaqB
aM/TRAjZSUG00MkiI0I7ZOzsDbqkHYJgYMYPwd/F1XXofBQMwJsNP2lwtnkpy0qn
mUNAzwOzI6C3MuTq57WX3/adVGvrqvtxPKRWdFbHks8VQscFQtxu2q6StEsbY/xU
mnqu0U3XY6gjgs45224twNDdYB9UNpNqJLmCuWHGAbCkg70Xt8jVKcAKGUOzZp8x
hc0ah9WqQfxZODnpm/7uaq45nTq/ljxo9XwpV7BGWebf7N2PqQaaDirTPH0Te7vJ
YXeOgxbhMeLyM0nZHjRiCdaNLkCK6GneTICE3G49W698gghSB6sHK+Hklz4jN1wB
Ngt7ubHc3FoD4Ni+clhhQmXtibOrip9EQ9yCtDim1vljF7+18ye7OaBi6d05BTp6
uBaFwXxfsOGUrmE2PTzOEI0VfindaJwMrAWho6kuMER5O0FlJYF+nH6lEmB+PwSk
4UXyKFT6e6G7Nv23dXxqczqJ7AaMit1IWMT8yelHweM+47tXy6Om2WbwcRFinKIN
5v2/QXSViUFmTYoQ8kkREqZsFErUFaezHWIRpvwpbwiyhq3HMAgv8l3xnhg/B5XY
3HYL/142xcv/IzfAXYoVmUEH8lfFTwnCA3I3lHaEZBbVj2tZsA0BVAyWwY1RLLqz
yS9Z1brobzgYFGL1p6gpzFnDtGEk9g2NuKuAP1H3ZNQu3Zu8voBew8kZaimd7y5e
df5eWsZG/DhfIjV+wlHHY0T4hMHNsiAnkdXJ53XSmB9ehDzLbjjGLES7Pr2FJltd
3RIUi743Om68cOKAIHyUnK1aCpE8QpgqOkoTqypPfxrqwE6X1NyWTlfNAZ5oFi9h
e/VfExKTU71czXsHFnJ/9T89tXzmZ0tMhmY73H+pd3LXbcQflu6H6dHPFqnEttEu
pJYIE7vlcnuwxz427XQtjZr9VUsy2RUtiprtftYtxvnyOpZ91kW4642BDPIYY8K7
a+Dql7k37SzyzrqTHWk9wOMl+hxjvC1g0ty6juM3WsURksbgkfbma+S1eYGSfb+G
Y5seZhtqsbrKgFrWVu21mPPjksp6weDQP5haa4uGhIyj2Dfpe+rxSgyD7zBuPi/N
6ax2rn3gedVjEUGfkVbq0WpqvYARIugVhHt6HJWCJnevmZCGl1cnjb9b0mhFkn5u
LcJZprB4+7QoBvA8ARN65ooHSyQJM8EoDPLYjAJPPDUQUIt7ouhOk90ncdHFH7bn
xpv+ZqjThKm3/CAM1h8nbPD8qJ6R1FKZPVx2RUR8Sr/80M29wedLSo5Fjy2TUq1g
sYQxc8zEK2b5k4C8nZ7lcjhOF5abbYExyYOC0ifQJNi7EZOc7NR2pzhubQ7WFuua
7hilr3dCtUaZieAGsUWUDSaaaYKok+MF7NoMwu9khwjPQ9xVbX6/zOiax4JkMnSs
jNXLJY4BWFUVbk8b5ZLAfvogoT73K2sGYLM9yhrnOFE4ZknAPhqCmSIr/CRn4Ukd
FeLI1WS5dYrg0S7d2HxzCMkEZlEnw9AIjnit5J8dG4poiBhbmXrVZFxQ59OlOi2F
2DTtSICStqkQvqWLXG9hszTFe0J6vcmwt72G5VzCBFxbqqnZ0P6rh2BSdzrHuhtl
vTG9Ysm4UxQPSy11Ir6u78+b/ajK0kuubUQA98Bd69OLArly/SA6pT7Wjg2Ly0Hl
XUA1cOwLcLb8VexWUCnx9Zt1sqkxdCZZ8NVukwK+p1+othfx96spwUs8yl5+SlVs
VWv5pQ65QcLY/AX3KENj+Z2Ufdg/ZfNJG+pflaYS3IVzVQiyMIhGTvPiJf5JP8E6
ioZ0J57UTyfrrpFrVecEaIn/tn9m1V3srpmIXSAPAMEQggYk3XOwtZDaUwwr234O
L2o3K7SpTOFYeBBbakfjlBvt0nX8yx/nvYfJzzXHiOSQfynRKM71dI57FUADzfxx
2ycfeIvo2BWsjLAwiGzlQ2R9O/Oso6sUQso5MVFIwQ8jJokK4BgfYo6ycL4Q2U9R
Mm+pZMMDEIejiHcO0pt3Ktbw+3blnWtZnwH3yLEnu2+vpLT6SS3gEIP7XPsHcQkW
oyset2b88dRHQ7Dt+mP1nQ00BGgrD2KujPMRRk2Qmo1OQWtSUoU8KaHO3g1uoFU+
79/DLbL7KKwdRdl86FBZBrUV2PKf2aPf72vKvNPcQXFx4w/6+A5SwhjxnxrvjeGa
yGAVg/nn4j8kMAR9aJWGFturJr1VEK556xyksLt/wZa8jTJBf4bTmm4ZcghPyTnz
vm7X6N4/EbJOrvLRtLnM0VEiAfuv6S2HDFcXUgpbGWKlkZT6/fgxc8TzsNIVkOuA
CuQ5IO6Xb5zrcYeXfOWmKLbpRg1rbwOQWqiAguydkm0cKTApRUkpvlByLVivJMLq
LuImkzErxuMAht8x0sv+b6H/l3qEmtEDn/VutskgGsMi0I1+zUHqGbbwRplMA7YC
cQq+fCMopGPxJq6OMWN2qCAhVoU9vo4JEkPgT8Wpo+pPa+LA4PFPnreWhykrgVOt
BtWWEkuog0Buvcqp6UA+tQNpbHJMrm0DdZEspM6A9wvIv8DQnIZc6JLdfdZrAHpl
v5pdq4bCFmJ7YZpVFBu1hkiDF62FxR8J/IXP3gGsSo/PsjoYHzk4HhxDfbb6nTTD
KvSNq1J1tv/96yuPsGHpSyg2J3oPh0i8huiuAwqOkpqlHkCBDJEhrK1H4cbs6NIR
vea9HzBVZCYlynGvNfd9R8KsjdcArbD8L7bcxPJMnYz8uRy5x4CydES0y4pIAzi5
iW1bg13KJklt9zAxfrcNpH+f6TrZSLtAWrsKTHlfjZFnQByrqZXFjJ4qI2rz1bx3
9wAfokFTe5mRgKsyimqUjCK0iKkeqCcmEocLXSxGXh/o6MlixqY4Em6VRBRlP++L
dAFjYsbx6agAI4ALRYLHOrnh4VQPFdxZ4xoLhr664ln3tiKLHILBTl1ylGWYTczd
G1hiaWUYXws/3JyXikpNAn6XGCcfEe5wQO+tGe6yt9ojLNcAeTG3769+KBe52UEo
BKuzwrKlQvFDtsTb/ks1LZeic11FAhJs2cZDxLVzt8TZts60yMTaB7TrfX7u3j/t
OIHPhmwxx+o1VDopuNKnxzoaNN4hisieDPVeh8NA7+s91ECoRdUCUXn1S4bCUWVP
BUJCWIqNcOQ0APAKYVW2z7Uu2PSYzkWH19iGdt+VU7WCymvwUBNJdvgALAi16v11
8zataoaZZ1//e68kGRvEzrAed4W4lTiEYIy8dNBzmlkKSqiADrcR2TnDGPbw9Nuk
qkz+8ACvTmOuV/Ta+P3WR32GuLmYIzk8kjlRBo1UazHyJRWC09kPfPHU6kanV5c+
YR4Cy/kNNZJ5Y8eMUZX5xrgxgcxw91IgyofahXmLBFNP5ZkAnHaVn/+Adf7mFTrg
yPq3vjvqoC3Hz4eAwGnoiuFRHVgjJJf4XzPITeH5IPwHL+MFv9r225kW0zONFqVZ
47N/L7pw4N1uLbVxD8I4RHAIcmznzv1iziT4hA57BBRn6LfbHCRAJlJGY7pPQVkI
CNw0R2ViY+MeGkW/kWDCOHfFhB2NGgvzMo5b6cdRj8PoOnZ+3q6Dmh6KgSiIOaJV
whw6DagFgfG1it1E1tqIgSTL/p4e0b/RQD6k4mFgG6hZgkkWvJS6PvbimZtQSPwS
9vnfXFCHolvGLubGHB3wZnTI/CaKKnxva9pqqGnp8RRCe3RK5hGqSlA+VgNG0aM9
aEyqg20MI4NxQ+vxY6pHQWI4Bb/yHv4SpP+t5Vwu+jIsEWVVocnpK44kVjLFvvHu
SVNQ/lyPV8xWVkxkvRvi4Wn7PxcHsuhWbwvog66yGC45Dl7AAvvtTLElB4l7WxGK
1ZB1guTLoeYX3ej4FGTmbj70oyFUljgO8mSMfgt2SzWYT2UsYKm1iBo7VSqW88a8
nzsj8eStte5sPz8nz4ZwQcC0v3QRvGqou5g7JRsrFrQ+9IrK176NEXMO0BdFpUeT
QeshNAxiBrRBlv6AidSoP3F7x/WHQ4hbQ++A86AvvgufRX2OLf7Nw6BOdQXpTqrY
3vqxeBhOqaF8sofsv+jp3P9yw/b5LnWT4pmI+DAKNvbMZ7sxaopkWRxd2almW0Lc
olG72nCVrk7LIIjcuURcgNxsXQfescTt7Wvb4wUAV5xI7khdrweKffEh/YuSrVqD
NrtDmgZQRfBfvtqPil2Rng1zukS590EfacEjdLt6RZHG9M7zM/o9QCTKM+Dvg92s
DhnuZ07he8fTKK95vn1UAGxRvgNz2A5ww8oi6JNPv78rnovU6SVRhU78n/b2h9L3
ar80Dz+SJ8hwVSORi+ElZSgsLN+B5u/WNrJ5s6unHRJTW5C7K8/n00dNw2hfBXSJ
3V48c1rCXBzjlsNvJDgXqFmrqKxJVlWEQSvRvndVSYwGXsmmNpSDkKSuOEQLFIQE
Ffc3fn1XBQ0VIYnstlucmWONqZ2PfZeVbRcyq8k3Dm9IQ09qliLW2pxtUQMDksMn
3f9ryYoeJmcnBxtgOh9tTNknqwAx9doeh/tuD+Xo71PMc+qRx7CNMGpt1wLjRURX
Nx7xhY9r0RBmJ32VXYQHGsbrhHtGZMAx3evrI8gIiRc2reN6vudNeU738NfdwwLs
RtDs2k+39dOtgTGU+2CCxqIpLoNfHJWDmseEnLAgT+ljusGYK+BekQD/geKD2cxS
rgwpP6zwlDbh4/1YUiuFEHuJQ4A9A70YoGCEd442+jSsT3gmKwLEsnH9/vHFJr3a
3ffTLrHkRWiGAGRrAmRbs3cKVt3SExroW0vsN86kvLslaNhIN0RHWohleMlPYO6S
lgqnIJS3uBVuW9nHLccIfuWm9zTHzWKrYo8Pa8us+aNM5K9M2W0TywdvVMEBuBhT
M2lNf1YChWCyV1RHiYkATfVcu2/6iyAmTWYgu3sKUSOzvVmK5szc9i99T6qopXjM
0CxPnKexAWRTD4qAUB5G1jiPvlLUJwVrNro4GMVluxjRbQWy/uBFM4+gHillTqy6
yunpjAHQU4l0LsX/ek0iH9nJ4gRhHbPqpxEXsdqHNVn3F4pm6luPK0rMzcaMdZMP
mcoN6G4uZdVQasj3KbzOSN9kwKKaGoD1xYwbsqTiU2IKoURu+PnhOE68t0qvXz4c
7FUNPkXlqVwtm6HftWTRlxKojhKaUcGJ4Ar+BD7ElgesT7QEmMK5UppWmUUyQf/G
6ueJrsHbamPuheYCAq01xrFRVGsMMaogV1aZRekwWCVWM2YCUQiBX8bbQHO1aQJW
QtXPCmrL8O2LhvacDyR7S9cOSPJyVLZ6cBm8co7ji1B7CdkpYeXBYPvW+GLWId95
9a+O/h/qQgjW6Bs1WmDJJazP5F9dYrO208IcjgaBiMljzuhj/3VsKBgUtb2wUu4t
l/GO9yHX4A3F16J22WwSnctQsimpmWYnA/fSIg4+UViofkkSOMaHpzGBOFnwfLXt
3CK9+/2cywmboL68D2PTUnjaV54pZWcgxoPow9fpIEZsTjTQ4aq8Vz4LgpajUsCv
etT716VbpEQ+V6dqEOuHRCYp4fKE7IDRQf/5JFCnZVxldFNpdFf5HprUZHpKFS0/
xOd2FmWPb9WKtCL3SubTfn1ucIVZN+pbx2OFbW6K26k4e5gY1Zd4aglOxaKrMPfB
9EMfRIAjrZNmCOyIWBtMWA62TMK75u+xcLeNd5BRkTzMJtIWCHQB12YvXuCHNw7v
fp/3SXu6e+cwqq1zkdCmQTuSBdjoGsBMpTGE8ZvI3dvqfLdlElgCFn5l1gxFcbmA
lm6cxQgWeCXnce/E8poyaJMa/dcFkJVoc/FmBkyyvNk3FnwXFeyXds9DugZxdePv
Ok1fT5d3X4d0A6aoPBYHJm8aOn3R6FhVXV8e636lJmWujKHMtY/kyvc5A1DltVA3
HKlQZNr2nyg1J0IOHwcOaZnBFEzpw/EpKhCtP31UJw2+h3t4v/vAh2W8/b/6dJun
hAGzSiWaji+yqT/KFAadh81IpXcr5bXmFfwq0v8Iv90lnxApr/mrZLFcEpbxC99a
2S8MUcRUk2VSAQPbQVcGQ4LWUPrtskc8DfH4gO/COzehV9cssaAryha8rhPRu1pk
DjBprAzagufArnrTVpTII+680clAKpyQHLTeQ/kjpo5bspkgc6CxHTdaA6O+Z67F
i8rlO4n4hQb5yKyRg2LSZ6OIHCCwfv6f5+3o/qdCdOzcahVBEjPMh0bqGeCYpZqC
h4zw44B90g+eXKlL45TqhP408yzXXqLGynlwU7NdgARAsxvv88JtOQO16l1ew8AD
8AAfSyDf3u08NX8VPLRLBI144XzAoSGCoAxaguLvDjnWcpWR1k0QmQ8uyazxth8d
PQfD3iixiR8hTRkxbVxVoIbLHtZCA4MPcbSII+aK9nbP6dHcaucgWOxnGzKOJITE
IPwId9Wg2IcEJusmfbTTVnmLRyun6dS39VF1LI1Zci6iyA3GTjeWWZ9Ky7/Oyi2h
hcBw42AKoY1R7SQXt35v40k33xvB2oD+32ryzgJSZt6RWg61KNWljFAEP2cooyBb
B3TIN6l8SBsNbxYnfPMv0qCpeLp350291aWDI8HJZh85BPPMYbCbDDoSHzfm2UMM
x7F9wHbmCvQhFYvulbmIglwxQVPqqWQxr3VL4ftM9oacFoPUWaZpuUfaeXNbmvfH
xZzz0nBJ4yvTgpupmKB/UJCMx0NbE4dmbvgd4eu6U8UroSjoImLo4ZIor9lKcM8l
KgTmszSbZRiSFZvtZZcNdvQYZ1G+Q+PnQsyWS8ZKq2llo0OobahRoO8K84fGAoUL
58pxfvTrV70mJILrkoGHuAoniD1DLFAmog00cE2u9Zo544DQ3+rYja5WOEUzpAtC
s3yWGgsnp2n/HoKhnOGQMuU3NqrOZ23l7Ic3uLn07HdynSDqRd/zpQrwu5iiat+6
D6FCAlIr3kTxXXqGykkWrhDprYOQtICyNcyyDm1rYj+jXzgqTn/JJjqD4qwcBAMJ
g2qnVDK2R0++vK6W6i5v1/WaQyHLqad9K+XGZtI23GGtQ4KVO0r0MrK8AMS0wf0F
4RvsU5YO8Hpl5uXh/e4Y+/EdD2eu7HXe63vP/jgGB2d2CK15W05/0I3CkzvwK1tD
0sIQRNbj4I/RE7HN5EXWL8gmFg76QF0MVaLkRPz7csBX0dlrA6BswfFUjPXOhLLg
1YJ9EwEtY7D6tF7StJNUHZdLLA1x91/Y/l1seA1ko3xWxTyifVpYp67O59yt1CHd
1HVLwNjeQCA+EyjDrqqxk6SLnB0GJePPHGMXEIDJgjV/WXO3o5ZLs2pGS3NqR4++
cXoiwHP5SxXM0ZfbEaORzmxvjq4UsTBl83qn5ypzhPBnZ6OggHe/yWpyneRhjvQW
aW3ZiuME/cr6V4zKKIemMPDGRSV/dVYH8SZ29CbzzU6G0mv6iRyqEh7L51A4ItBp
dBIi4VoWeTgZuDl5rJAxr2uxXwT7ma7qyddNKtfLAntpQfdaI4E1LzGcDrGu9c5Q
8HioIH/hZeqImNTdoK6mNnp1ueLtnBZwcX3I/qNOOpAE2VeybW2AQTX+U9cz5bLC
4fRPx2v3sFPB7/gJ1Us57T6S145q3BIAxIGLmL6KpiQesyb9iD/hMMS3pOJpEJb/
Hz/xwu/R4jXDq4wVvZywcutDskkLjefnUEOt1KhZ7ccQ7LDwDtuF03saISLdMveQ
arOGQspSm190p6jw2yvdVmqSFMmQOnajGRnIgOs5Ula5RNHpeghzp4Ueg5wtda8S
kd/uGGRpzrg/3OLQaddmZdD1pvN8IKcWCMz9VoLSPfQ0zbl9XZJSfQXHLYkYmrgu
2YMrzseUmnHXNimWvonEeZbkrQYGUPuyy0mpaAZLsvpl3UGvrklergUajmwDE7pa
A6NVw78/R+7VjZcnsexLhBU1gFxsW2OGfiCCRvob+fHugyOjMeelQYWTZ9/fcPQz
H0Bydivg/AICgrRSZJMQ60f7sntq2TpXuFJ0eWjQvWIs6qwGMCc+m5g+zso+3c/S
XUxVQIDnrKl2MZecWoEfk2F519FHy2wNJ7CwN0N3ksVX0U8JqRBdWS+nM3zAEGJ6
Pjkug0ODQX12EcTc6+0Mc4TBwJ8f6lOMODDqHjqrA4QBJGJZOylFv3SQrSDLqeAn
N+H+fDr6em29Kx9ZMer4PJIlpYQtZqtz3EXkNJZiWyagsfMWoMZTN02uc/DgZt5i
FfSAUrFtKahycYSE+DGNWhTYhY0SXT2pNsbOymwlqRWtYBT6/zGFp4eklmRxrnlV
ZdAr3dXQwmuvVBUA7hj5Q5W9tLmCgzWpzq86QKjN3HBH7JhKObnjkqJsvEuO5RIV
E+fTmsGLwNs1L/0v2IuBqKpGTPRLz0Y5/y/trXxAdBJfDV9wrYYooUesXf0IKGRV
epLFDVEDcEow0LFfpM5njzm55auVgvFpCyzFpwGUMY5epwpyO3aYkQV652XeLXyg
qNj8s8iB7rqUNMshM7fcLWk8N7rVAajPX5YTYzW8M7P4VdTseOMcKeTjYckf4UYS
5IZ442yKy6S4/esCnG0DY0snbK6Uhh09kpmof8/1FW5OvH2AB9J++vRIwJJiFuMV
EHdWVRBRe38nUPoAK8B54hq5k4Q9v6CeN/pB3BrxeVS2ExGqtxh5Dd7t68CFIOAY
6+XMRv0G2FkO/854FWKwfwZ/rT/WJJuN8bOvFV0yYPOoB03SMe6JCKdTesibuJ4I
7FGN4LRh2yzdt4tdhjtQWpTy3mjxlo5gsg6Zvn5sbg4Dc2m5rgCFsRNF1s1wIQqS
AywihuaKL40Qc/uIO1OU5b0xoomi3Xq/JElwL+s5d0kVu/QdAuR06u7yPHM3IPjX
yfvi/aNWlF5yDQCfeJhNvOsM6PfKM6kzC0HUq0BkSJA8CazdJ7Grme7e3pqKNklS
cVsej+FoxqXpF9fTWzrfmWdEDfnkqdrW1Mk8D8ElRLH0TEf8fw0bFm1UYXpMwH8n
B5TfHRcmsYNFjZay6afe2Q0Qk3Mqpngsf9nR6hcNErwc4S7aERS5R/eLTpj46rD/
ooeR3shuQJGIG/egB3yykHZFQzlfBU/3tK5dyI/XWwW4hJbXE/iH3kLh42DdJWES
4/stLISkmBrTwOZmon5aKKsA2OiMDF82BSitubghzQnSycf53PNBR24Rp013BfaU
VXW43U86ioTVvqJD6nNyw/E15iS16XysoHe6IM2ZO6vFBanHeLBzQV3LZMlDcQcL
12W07SyH1YJ57vpkKAzuE6BWg9Cy35pSEgq3rl3qDsortDjMg/9ipeiLxfYK5R0I
uCVdouME0M9BqSfsjg6EGlhF7cE3Z2KuglhdinGjNWpGxkCTuK0nMXPP77jIiuDw
L2yD0xji4RONh1AdfNEWhjt51vAuPs7YquS87sCLDiuVHaaRIxHt7P9P636YjQNO
joA6gGHSE+QgJtfMSDnRAFBDVGEd/ri54pwbo0avpx5ItPQd/yo2OggYg1gVNV+T
X0G4cepoTSdvh0MY4SqQd1rUal4wR+CtjeOgi83cI51ouO/D2TpAdxv1/TqCix5J
lWsdO2o/X02FlI1+FA1xVbPyakLTDSspnPSBrMnggcFw+zqQgTLatlDff6+Drrxh
fuflX6QFYk/DgUDWuebIf6OBJWrbioNZIQNNXW0Jk3uQMPP5XRAzeeCqfogC8f9/
/xbTfG/VvAR0G07shOBRHM3qcm6QYe5BlC86EgBY5iLYylbCk4oQHX4tLEtvNWWC
/ppSTHW11DbAWDbSfW8RqzG1gZvri2oQY0KEwC5xfFpCyu7hMLLNujZwT81Pw7ty
kCCdHqL+u2MSjE1DyicmCUpIVydZkU16QaohD7XbqlWlnq4sqSdtTJ6jG7OoPhv8
cz2zIastYtygUDYK6Ga0f2ImP+RUCGcVNpu/nVehnSFnilqEneq1pvyqZVQ04p3R
EaAc5g3KeJQZG+a61dAwVZZLLHWhDcoNNaPRpK03jnBV09thRK0dJVWPychfU+qs
orlY2f9qfqSFH0puQc9M8CuPRWnCPjQ3Hszwt35a881x9jX2gl5QfDaCkYCppGTI
Rb2ez3pOAUSfBRj/MiSAe3XSI1rp7CD2XyLcSXZFMckk2IJGfYiEWHqtdqYXPfd0
Ky3NzxO0fu8lWw8Jnh+fxQysnfMnYj/g9OigUJWEw9J02jSPMYMAlnnArtTqYPgA
pQ5Sj6blf3UbZFyZbEr4dpQboUWp2J/mX3GA91XhAHi5dB9TWaj5zSwosxgy1vLt
1DO8dJzgPZoScWO2AgLa3MDtehQi7DRYiausdXXRpiFPt9sPx3Bp6hgsxiedmD6B
E1GbZ0w4WSt3tr9ApVBoh8uZMfrtbAvb1XNtSdCWqUsmaVvnZD6Aio26HlWXxVQ1
4zehBFjSWpc6NMwUUYFI7PlCZ9eLTTzFUQNFFKSABLys79VRbcIIY2eJzvEc2jI3
JOFFN1ro1avZ2g3KTooI5O76XEE8F74JwnOtDb/Zyq/jB30UbyYPkUzyULxqjQ+1
kTSHPd+AUJa0UImaQOF7MHVZkVHq/SK/aOWfTa9C1DJ560HVli5fV5zTHn5FurSg
D6UID/xe1Dw9tI/S17uE/ec30+bXdqgbN9gcH4sh037G2qLa1X98jvQvb/zOC6oG
JLcuPZ/CB23DNoVhE7f2CHH1w83KsjxvUgQyWYb6ARt6sJ3huy4s9vY1q+JJJKax
AJfL+vfTEQhoy4i3gQ1nDfZujU9XzyW01MTKDAtiuiW1PXgzdh9mRS88AIZR2dLl
IHvdeE6UJdSceIKPaQlHYDuz8q15PBJmaffO2NJkNhxO+bSgEDGC9DKOLjb4PoMf
3jmx8xPJOlu0tIeKPoRjkCh0rrjbiJNnzdjK/V5Crn5RQ9ySIeQVD80hj1BShHPp
DomGC6+siroo97mi12U2mkvWPOueisq4ZctcyUWzfilXO3dCwxWa/eYYW6F50wKW
hO4MQob1Bp1iLu+aeE7SOFwxVukJfh6scrMBwb08ONmBbgx9ZjIHrGnV8iFTKL6B
ULEqudf6EmtBOCS5amnB9URTOpGjLheWo/JoN0AVVM/nrviU4psdDvgWqleIAXiW
vbZoLf91dl+vkYtB9kgcBIqH+foKZyPzyr/pnlhmLu7mxRuHqKOVFY++MpIHwIMP
RCJzhlT9g9SIJ3ZFhHnu+X5j3a/iyQTVIOLSBkEdc6pIaNaVBx+mXn6QBau/SR9F
QL1UO86JJZ8J4nPV7zJr6lBgOCKh5cLxFECSWpyQdv0EBxMOjcU/DUi+WGNoZcXY
sqQ0DoyinUIuxTX8RflppIYrN+Zzmb8E9dmuKLdy+aN71Tboe2hWGfNy7PsJ9MHn
ym8pJq6mR569/75RgoI4oI6rgvCgYawIf0M4s26vHiliDvVJI+0N+spTBx7g5nqF
K5Qam7vB+peTUoq4zN0WOWxoyMZzgRpd+8CkDO11/VFjMqCm2NI3j6PUiDbDZThr
ogzqTWxlp/2KBhfHp8oMEHkCP59wKno2RnBpNLCJHV4t0x6lp1Jue6XAOJy/PTDk
kCASVV4RqQXjgQl8xH8+3ExOr+CFQGHLrkeNWBYgzM2udvf1C8UpT0ErWaOTz+l0
GwVaLRZHKjIYyOXMlixdt8lqC2JS2GS0nBb24SMW321nD/cGWBAS05STxpThmp9a
DM5GjK40msbcTlTaes44MsowVrvHqoOg4T0425qP9TdBtgdRCW/CftFqlUuQt+sq
L+gDvoeNbVX6eJId4kSyPqKi+7Pi0hO2xFJKvoKDn2kxSmQFrQMP8XY9TBRUDOMk
w2Sxu7f06iIvIg0SR1+LpXPrKBB7ty+Ht4nUAjwt0QTslYbhroAKCXkkJ3ZFP604
osE9lx0zdat5ymBssdT2/i435ExyIN0oRxi/trCRlLxgSSJfPKrLejiAQUQZN3dD
55oTz8bweRQpaxCr5CcE5fdHDLHA+1DUEwW0q3yfPgA7OAntSIYTpG12Au635rrv
R6UvamlFvKYkez7VOjE4t89pksd+ym5p0ekiwfdS3+0hR+yObJ78zYiVutT9+Mu1
BSTWdEgehd6d6JK70YEPUfPbQeDC836cZVUjmH+jq+2dKluL7Oujwo9L7JeSBdPg
z/6SvyQWMMwlBB4/gwtMog6GlpbqvIf9NXf1udP3eKRKmLdBJeQ6WZJ3bvw/aRsn
2p+yE+/R5fpvUKY8u/9smm07Q5MaibYYAuviL+KN6uup2j0BdONSYJlSlPwwxB49
XGgwIf2ZoBD0Lg8hxOLV/eDvYL7HZ5Ai0keE9aaVf8S4uipiispHZMpsY0szk5VO
CYqe5JTvMU3XqlH2FHaIfHzU+xkpb7zGqViMFbQlCiZUizEukRQx43neiJvbpVlo
GSkwk71P+NIo4UQ38btw/fkVqzi9SsfhneJUfCFE8p0/gg5mjhAX9fU15Rm5/o0W
Rk2es9enq13xLorBncPcjMH9fAFXm59Sp9cQTILo/2lWtGtA/atv1nlL/otXjUW0
bp6FyfVxP27vooABddvdvGiyp4vT6pXy+ZjP9QQj1zeiV4dtSsQx9B041XJOfWE9
CcokE0VZDYXnk1OfjttmCh6SA3SbcstOwgzg/HerQIqB1BbmSMLouDGY/XY5ZBU1
vOPLf1H28xNDO0MalouyeMl695iP6zpZITc42wcdOB7gE+xKyj9xL5Q2VVdkvkZO
ojLs3NIjQdKQ6sPE7eJFFmXteiIh0QICj9x6qGjIHksf1r3A7sKP9m4yyXq9UKHM
7scG7DZgFezWl2iBp5Ol/k6o+Fc8XdSfaGwR+I8KEo8QxIE0yO0S5/rIcnbOXnq3
HMyir/7GQ0HLkEAuBAeVA2J9h+0y81pg26y2Jh3MOItyCszYoAe7VDe20MSUSN1z
Aq+zTKCgIWwgQRytZk5kB+l8d9ljWL00Ytp9gQjRToAV7w61DS7/pnll4B5Zi1zu
POWJ7atAPuMHPhvBWSuczMjqfDIFtcO86IP493leEnW8geEWL988bUKVV+L5oegx
3ncSUklUzsMWzFIxcMCtZ4ClBu7sbxATAH79o7geDBbmyv6nDjRfy0gIoj8Tpf3e
dKt3EpJYAHTLk1ayk/ZvfjV+o7pk1AoLzv+EpjLnJt8n1wuDrVm4S3O8rJVGhPss
+iaA2aEL39FNT+bHKSwTj/8PGSp8Lgkc47p0GJug2UOhD/XV/LPG17hCjJ6IXnWm
m+EjpU+FdJ8n0cAhuKhLNB8Lc4Bgd4N9JongONBijlU8hQB0lWFNk+q/cfI+xyRA
peT1wM/QaoVuOAnus++v9iNi5h8yiMxCjpDLadxm5zcznYF2S6QG+q8nkKxc1DHI
aLbbyybJobId+OmNZT0BTNKxZLaIRD1hr26xgsivnMuIJHju8H48fizh5YhD6rEN
1vlFJRqwS03PE5NimOPKq6TT9/5W+nB81DFLO9pyQG7b1DlsuHXlm/9k3cj0SMgS
Pn2LDG868pRf2qTONo6OfSDYz/SNCRiyCxGvIPvEhDbJgDBgA1gMw8r1b0EgUrD3
e6YUvoCOdjK/pvrd1Z8emh2PZm4n3/SwQAQBXWsukLUJ4dNGmkiDZ+8VNSHRYX1n
wwOm/Bhbzzl29mpQ1/yb/ss3XP+s401Ixseb67IiDaaNDqHMc5HIwiSaf1ah7oaa
np7T3qC6mt8sqF9yEiNP+zDF03OcohNEKYHjzyGwWqb/6xzN9qGVDDARb/olHKsw
Ty21jlWzg09Rjf2104yAAuPblVdiOBPs8wS0O7seGXSwJ9x6hfCLkPtI2cOxgCM7
hQVVDC6j8d80Rfjd2cMj15HOt6sGN3i/7HD7uIyftAZq3AJxBVVu2xvwOoU3TLgs
rCZCQmpH1AzKny2iPE6mFMWW4ZM4SNDNy7TSFbUnh6yAfIBvgkom3X0yadRa4arq
S7eLOtmoNI1zlxEg9fM1dbJmLRtARoxHXXKxCa6ZXQXZB//SCZwn6/mVkKTR1Wx/
ekMbi1mEC7sZBpO0sTB9+4bVvDo9izYs+vw6ExP5BfiiIps+xfDatcpoTp8wX9i2
kYMkUj7KIZrwjE/0kut3dR2ueqd0HCcaOy0Bc4uJkU/NOakBG29U34cVgS4bP3Zb
qiJrviKj+RRxH4tWkoXxfBIEJ9xDE4SGjLb9Dewqe1mKHA5spspaImZD6vNNIXAv
cGP0B3YjVvaw4NFXiTvq0TK9yRCWUChvfUT3iMlzquGj4DAs1z7xoJtENir1sbnA
r84XuZjxdgo2JcsIXPEmlptQ0Alq8UtDkfbGfIHFfd9w5qj3mZci6khUr71DO3F5
I7YidDGt5f0b4KzrKEY7FOOXBx6CuAWeBTudZJvLF3q3aN3T25Qez1/L9Ia9StXl
SWH4qDhsqv7sztt6l31717PMgXu429GpwBbx/YjgRCoD519uJv14yqyWZyrw459u
VkdoIN9a5sluitfIplCJN/Bz5pLdrNI0DNZRi7g/MPUEkwlLutcWKEIIBEep4Gz7
lZs1HzUp6mimrfeB8d1N++6SyVq3jf1NmDo1+QghEPz66Ddr8GTD17cQN/iChIyI
mADgSp/xi1moIr7ZxCh2kLdxnXEtCC6Di8mzn5SfwrV64/ASzxeYRMK04RhUn/jO
wJkoh1qgJ0ILY5BQT5VjO1UwFu75V6CnL+BL0lTWFgFZPNlLUdb8Qm3T+eIRN/h5
Ub344bzaL24bzxKU3GkkJW39/qe9BWoM2xnhpgk1fTjjGpZz2Tz5pB/GDdLB6z0N
4RuidQtFM0CxIju5MFN/vBNyq16DkO7p2Yi78rOJ+OccMk/0gN4do0OvXpnC/4Cj
66p4wS2WM3jti9/jpuMNsAZB/AUc/mvS6qPJmHdIWE/JflQcZFe7aj2zHqTV0ucS
v8BenCQ5ILhM+6aR9HBHtEdO0iReF4/Nvhl17huLzqGnNDkHDtgyogythbcvzlLB
ea2ZllmBTgRdW2X52X05l2eJyuF2D3SkqtOvjty0MsyaVY9TdIsIkbl/4vVoWqLN
WoF1DwUPve143n5K+m+o5xrPv9vz46qyy5OwYUEdcUCXqB0ra5yL+Xhat1aYZfG7
hMU0XXtyPzV7x5j4Z7RFh35RtGDbuf9QLY21LixcympMBthW54BKaCgBYtwv9PgL
38VvU+RymFR/A3lB66WXhlzODgXQKKDtyKFNJzixPVkOoEWAuVI8R6vfxcaj8jG5
kkUu17GJ7yEO6GyDd3G5TNE4CGp+jJaf0PbXmiZ7w8qOV3N5Vbq5ftlRppidQxFr
EfSC4itIjJb56tglfx/IwqP0QwhO0wdxLjTCpgl/BuDeyHqd7xFoUzF8AjPHeYp3
vlyrGD3UJKEdzaHYrqMjEmp8obZsvPNl8iAnVI4LV9vSI8GwgjNwohlCOTu00+z6
gU6sYIfu8RA7ZeaXJNNRx+WSq+iv7s01PuJ7nY+GPxTwa2fBeChwWYzMu5PF8QzU
/bVsuzqavhlhky8SJHGwu+u5g1q8Wa+fmZmkyeXVC2v4XKxa3OYb2qDfhJIINxTh
KVx3hlZQVIQ0hDzA6a4tAwSZ6GvynlF4mRcANHr+XQCIg2QAElkMirwro4KSEpAR
z7b6dO8IxXJPFsr5d02FdJDGM+vrPLAwbVdIUugJ0htKSXOSpjq5JzKvIk37y3Th
xTT4rtV37wPX28S6vpSE6TM2tREQu6Lsd2qyciuRfedj53zGRCEwKjnfabVAAf4Y
sYlwSGuhxRwKBkbH6GTo3f3BPth5Dzi04ChkFZmjluKFAc7HrRDwCA+MNcWNVyXq
PXd0SF53oaQIdT5XIqHAtNRpbhl5+ng1rRwYBHvxWX8YEIGWbjgmaSIicHrpUOuT
mO3ArRoKGWgE1FI4wlVvfvm5Ncz6ZQoyqRVV2YxKzWjugh/j0Tsw1hZ8cJ8hPjlI
H7fiA4exqW4e5lus/ilTdBibr3hbK5TNH2afIXuXUXaBg7eJZIGhQQt+QJz6motO
UwqxaDsWI2Bzm/RyXEExSw5hV8vqyFF2wxl6hIqTJSqvfH+4WvWgbMp+1PHj6pyf
S+dtpoE2/Nlk839Vt4+UDKgXFc4ry6nVecVoRkPu4AfTzSkSG7q0UQaOdEKXJWmA
EEl/feLp7TZabDcKH46KbkhR9OaBdttRJm9BU/4LX1XbpSnHi6qOMli9kJ7YXR56
PbvV/q+bsGUVQ0G1H+hnvb4rfHA/bxneGQG8cL7qA4oQoWly1p+XI46oBPPI47IM
E82FjCmgDB5XLIk6tRVJ3psiVC2aoiHs7wDFzjfScO/RYDWnnzoX/Hgtu68iLpyS
7gYoQVsCeMikZkuWiteEO5s2jzB05Sd24QHMRxeGG8rAvZKWairyM8TSJRNlniJy
vgS91LN5A9N31a7NQ5by2ydEC98nMUNwD7CKWyU74CSovuxw41aBzmoAfzp71XYF
0evLYBm0RRaSUVJOJxuM3IBTBFQvoGjoeyzX7t5W/DNZGvh23DxJM0wftzBnQyRX
8CdOkT4I+G4F1bEcY1lkSWgt0ctNOMORxZ/s7XiSgmCrF1SoX3O0QLG1l980UIYs
8Jp5Ty4I+Tjb8QNbDoDxIqmS779/OOMwgD+qMnd7HQhFdKXaQy8LBY6jWy8+OYtA
OQttwqb/yyvu/ed/htPUrGipTDMPwGRqRaF3RehQhdPh0x8re9XR5Xx+xFuCHccv
SmOeblAWRDxbXcXHAqDLDak8vQ8LvGKZhETKsQ89Tgs8DyNqCpLstZxS3Ia8n0HP
2Q8M0n89/Je6KCpQouCszYlOdUwqxTWA7NDNrwpXb6aOGIfd1K0QD3ugu2SJYDHT
NxyfLCSJpn7+zIpNsSWaYsKRepLxPCNFkik2spgG59gXjMQD7M3ClJBcnJhIxI1p
W3sypO1XdJQXw5Ep76V9TrZN7ktkHJD6u7zc4YyuffcZly0/W7obCv5ulvFZ3rDb
uQumMcGvtsjdnlaFzCSeJ1grhBETpjojaZ8ig9rpLgT/bindqCPon6IfppOIQUsf
kMg4CPsz4kcbsFJMFLYZRX8gtM/+FS8roSxbxtB3ZTSl2ZFFzqEfzNfe5Hk1hLnH
AlcR23o7zW7Pv7N+Hwd35xCKCpKoMj8cbf/kEqIW547tIRr4Qk6fiGL+gepEZhpj
9YInJVaWLkNTow+SDvjGqm6dYpWUMC7ySO2mpntTtI67ySJJ7SXtDF2r4oGm0Xm+
qvZkQIRxvw6oC9GB5uaMq4Oz96unxRk1kcGbOS0W6HJS1ZkwA5NpPH4I7xWuJzgY
Zn4A+J9awc9buwh55osOZFoeE6Uo/tWeXeII13pbKo9kgDSJGurFVGUpmY4rD8Cd
IaJh5FW/KnJ9j9ULCm+CmNhibE0FRXNPiPyqe1E7nX/fc93vBViB51MVTPOJK3qn
OL9tZffB1hyUnpvb4+gIJ+gnSQc80grD6CE60A5mRdeMcYSvDO6QF758PKMiUG15
DEDqNL8QNFkLfJmxosgHMtRQ+/XSOZA95OnZeDHkPxgQdkxEUWlC+Edi4tLu34TQ
JwH6YG6Qa+BUXDD6WKLjs1AG3zs3zblLvLv97wN4943Z7odDOGPjz8nXyrrlzx+I
H7sMf0xhATtBAbOR2Hr/e4qNQDRsg574motJ8QwzU6mCLnDopf6rmnqguL9JR4sh
OA2WzyneRd/pxiqogXWKWLmRLU+xGYPFWiutOU6Uj+UvbOaeDHGhJw2ix9mR1bOV
rB/7p3V/nuO0AYHnBg2dZ4oT29TajDS/cfUMF5TB2rRbEySYIkV6NBoqEUmQyBUs
mQMy3KtoKQNfZYv6CCOuSbJ0GrrGPNTPAtM1Wub4c5NMGuVJ6di3/IKMY+B/a1mv
g/9sjo1/ga6W2Z1D7jDYhvHCbyGAq1jjyE8gSApDjPoec7kncCVtPVCngMijG6xC
ey4VYy80d2xLc2RfbDrhJWQ9I3Ws5bClEuBT30foxhxCutX+feyUCmuNvfpyrZQP
e6n5KZmngwlItGKmKHR4gZvrluD5nAQAbwcad6xE0dK49sx/RwthlB4UQZsdawf1
GpiGSFyMCPg7eFz76edLjN2qFhVZhzx/qtdgZBLjvu0VGCfo0pus4HN6JRp7TpRf
E9FPVwfp+k1/UmKP+ZCYCnPsFhcysZvwqrQU342ni58k494aUgkw85mTgnKng2pr
ONb3Lz8y094JHUDRD9YFC5sxFIxH3KoQ6jk1GkIgQDXjHdd57h2TpuzRp+5r0hZU
lBZeyt2QdgqOj9H6OJra2U/n4E44oN6cijWP/3bapK8bi+BHsC59t5wX92GuQ7Ou
pdvprDC59Wu42PF6m2AEAx0DNdOkhufAD5eWnVDZEkEC8D9vh3BEPD1aJwMWDt5T
NLLeMc00BGWpu7UswEdBwv5i39HYh+ledd9qd+19PLCjZ0ehLVSS7OWd4/xyglkL
MqBdzyJZOL8PYJCRU8+oRbipnptJAwaqoOHhP3A06P8mqmqmyp92d8x70d5ycANK
79rxXUCGse6qNe/YHcwDDSxZv5iTNszz/4gWts/pU5OeX1aaTmseCqZVaVnC2SHQ
oDgVCi7rsm769hYBglLR25fNvw6mfjnoIftZ+sFax7TtUf8LsjaQd2/aGBGGeUS3
S5707UCEfczFrGgA15I/w6/DVjPB1cbknk/nqR/o9bcNm9RWelc4wfagt4mi5pXu
EUx1lcFV6sS5PKFVuWgOVLjEX3wD9jhLJHlN3j76bvB84T1yPvLZyX/WqQAYT0EJ
G22VfKUV9GLfFxBpv9O8JiYpHcBV/BYbU9I1wrdelw5qgH8v2S2nkw5mjiat5ya5
ronotvLOS0kajJPERGUca3e6bm9ZFH4iT6YnXM5hERTP3e5RHMN+y2GKjEcE6/+U
WYeNuFZJixl7GVK31oi1PqqKrUWPOjO3HjfeFPGkUZimzppdrazIGjh5JjGc/qyT
2bs8f3du4WmP+2Baaj1PE7KRTq2Wg1zJ7niNfo1WoIS+KyiwDLuQoa+waZ1DlaKk
8ElhzR0TtO0S/K+V30D+9Shm35n46bQkjHiDHIcDNqQtuDDxak3TYWLyrH1v0VPx
1bffl+vAdhbsPcV2Dv0UMdtZXkft3ZJgixScBpPJuQ4xiBUoZpW4KkMObf3+C+du
mg305f8KzjXNeOf02CmUlvP+y4I2aqhYuyV/abhRkX9Mhs+/IR+nakTNDNLiyIVN
CAowijYRFFciGqzL+bheIDcROKQJUyrNTC2DRFJqiJoyrL1qn2j/7BmXalZuralj
vVUmJPX/ZHMIjnwtNbteFpfPtHqioF1LKHDBNrstqc4tNP5V524RJcPj4YPTlGky
tdY57MFDGy4++WtPhXey8M6sEId7JIkH2GPVrmRmYdXJSBVjwjUD9BmlCpkPH1po
b01+PdLipE/P59+E8NVvqG3Ri0jWktOjY4vIxgNqjpdkke2ktorn8MhsIL9iPIF4
1r3TRpZqhykA68rGniIIYt5aL+GRY/1XlWSbwhrrvX+pFm/FqCHQEfdGFW5DLzsx
iaSu/3719/41dmCJY6Sd/CcOpRcl9iy7nz7SH//xuMUa/rZhiZUrtuWaX2mF2dgd
Uqm9IANLhHDOeeuXJkEY/0e90yhxBFXWTsDBwjvcoufoTkvcvIzDBR+eGYB/nPQe
zoOWlgYfTJeeAYh/IZugIW1UutLNR60m7yAjaGouVTNK6iThamRVdIp/U4D2CHih
FiYOmjzYa03b6lwSzDgBzofqP5DtWx7ASkGp7dd25NIpj7bTNvXnFA9csQPyNFQM
OTX30iDPgmFerXPey/WmKEuuakEBcJAqC2ZnGmnLj2KhC08QNIXondXvZ/sFeDw8
Px1LjhNqfbVpBXNMLal7Jd75D+fIfKlod8s87hETQWyVlBFmIx1/nQJ4uz1OdYI2
2uX46hoj7zJvHuHWpxi/BzrSf+hwiPeCE76lh93stOHPJIxnXSHEMmpf4cVzN6I/
yywTCFD9tpmnPbYOANbCGltlS/MsEt2aDX1CSwQJR33aJxArIUnfy6uQuTHiCGnD
2Z3Te9Tho3d0UETvahmXdJdsyJU8Ask8GtIYrx11CoigiDLFzYBar8jDA4r7evkq
TfNHMjhfGfaoaKkU96b37B9dcFKUhAktzbzxTLY5UMhQVQ2Zs4mMU8oSoxorD9bb
l84EYSILAq6o1MoaKsOGX9QeEdifuhyAYAfhwjy6fgrDmze5OFybL0wa661tOrjD
rv1CK7jGrLjNuoF3Oohyv8Slq4NsY/wjKjO7ZedQeS07iFtRlno1EddB5vJGU0hl
czM1LcfMP1FaL1gf/Jc4je9FjY8HDjhe0uBp5y4s9HlKgCBNRrOkmYgI/FVhZqLA
MojOL53g8gGO8Q4g2j0VbATk37TloAvM+LiVMwPjgZmKZVakvPMQ4a5UtnwYrM+C
YOfDreKKvPuQXjXCsxBfXWlqkzDYtVUHVd7PKvmYp28nnovDgq2eVCOA6StmJQKI
zDy98ZtYA/2CfHlHnngWxVFwGgGXy1AM7bS9CaAcf6qzpEPjkmtDkhM/e4kk2DJN
M/nGZxaTQDPBsaW8NcvJVkDQmvrvrghrlTN2/dTTdM5jq6vdyXUK8RBr7eb5qUeF
7tsePd8B/8fCEO8MMhI2YTloHSjPPCoap4VswLQTniXMAWLtuSRTtP45ZyruuGKO
McGmKZsvogyskNZ/zEU+HQQ3r7LgWUkD8lE2gxL7cuGWdccb5Giz3cH4pqzSQy3M
NUlLXEqvIEYcXgUwjLtqskFrO9+Xg/CObyCTNaFMT0zJPALC4wpEFZ4wS4n0Lstb
+9mdER2XsD9V+QXcdqkBUWouuZFufBHIohObNgBFV68p1MlzbSKOTUj/3Uz28tEw
0QwMXu78PoK3068v/T3SFAx8AYwwaMeeRsknkqHlUImxBpJAMWqQI4vmt1NNjgO/
dP7z7l2VKnyfPvTUISRT9+vKWPa3bMwiluzzNkwPVD1HhrsD8otK699Zs/xGSeav
9K4ADPFFMx702g75ip8HftO4/WvXD8Lrjg4PIa7EUvjcnqh7ZSgM8ZmHBgvyy6Mw
Pjc5umNDaXAjXeAfxA3sWJOVGSxmDbtxNsBZAvX5TU+Lx9vcsaIMAG+4wyNLM3Sj
rit4SEUUN7ZubF4r9synhwgxAcnT00v7rhpF4uLE6GGhOlcADOO/bZu43IYgi1hZ
0oZ12xMKULGlRZs8LHeJQL/7dsks2Iovz+UrUU4/JNY1fzeMFQoDFVdg2vyxRUHx
Q1KirZGZyNt5o0zyNTf4XoI9P0ya+MAKCVBjCZaPWz6rrslYKuW1Nnqkgi/arDgg
XBgD96zOf/2UeEopAOTbQCUmLO6fwisxlpFwbvgH5XGChJoioW9VqLP+8dRAFNG1
xyax9HrmgSk1vTUevCwwuopueqMiMSEbxtEhNMh+Clp4eAbv4uVsalw1HONAPaVF
7ydb4hWeEJF+FUW8I/HIldZme+PFtdWMH+oOf5a+xf9sNYYRrIijR/Za37uXFkQV
LgnB8mnx/UlosVjUqNV8XEncgkCxhUUzOF9xQg4mYM/KpAFhoQj60qRfJEFMt6RM
SvtZVweGDtWdUHBTs3ywauA9qsHqQZ5cKbBfVwm/vdKu9tlxOLWUUxRJOfyYQMub
bTFjbc3xCbF5Rhjew0CkarH60AzQOqk1UacXXirQGwhKl++Knqp6qE5NZLdcK8HX
/ymAtTiS9PKKDt4vytQZg/+ENGwelc6sn/FHJE5fFuSL8tux6Ow2OPAX77nRaEUK
1p8lA9J+whxA1qMHP5kS7D1cdNk5cYeXk6ncms/vOhgs68kGAfwxrbwUH/kUvhrX
OQ1AXChbslMNHbtZiePG6ZdEX2vteAI0Q4ZG/786qas9nvNUEwglCORzixMHUxE8
Uhi4ljnvE0qSh8pTN19LZRvpjXrm6ph6WKH6mF9cpv7UdhF6I/XTkx2fKJInFmKE
0qcuDpEOTinF5qq5jXffpwRIMLD6brMnsoZ6rpl1r3rh2Ypj7Vf3vgVc9yw2y5Ff
r9HqYLGy648uZ2F+GnLux9Ehb5/Ctybh+Ab3RsyfyTcBRpmV9t7fzHd3/PukLash
1nd2foyMzsbOe0r/l3KEwhbcMf+yZeJs6/f6A2FX2p+3KOgqmFefpAZP1PXqiKSW
+dz9ppj833t6I0NHycuOHX7dRdWdlRoQu427dYrOy/7QQPuu2uLKcmrDDBwTRicg
fVrflCB6OGhaV9ntzMDdmyo6KvCWJYcrtDMrIS2183I6QRXXME9AssrMtc0kdNeT
UPHSPPmANdabRm6ziFCiu6oUKrraWzPml8MlQWd5giwQKOqrUvXpiuHjEV5Njc7O
TElVnU5f63gO7tKPxbrWlZSHjG/UKcI3wY32b8k+UtrON2hpL2rrGh8cAcFYQG2F
2TYecde9gw9Xf3/hUj1v8tw3d0U62xOICbdEC1FpNl6Mr3HTu5zA6/ZgGuvrwbSL
Ze2V48aMrXgCcDBOhzybq0574q/7QbZjalyR7aUUlAi/XfeHBgAFIzzv3/G5sXks
3Abhjo+wLmErbFPT3ccsQ1374J8/y9mNj78cszmipp5W4A6O5J7DyxW9cGuwB8Go
8PWakjm1TQnjtFDsp181MoB0bhAxnf8d68kundD4EF1ifP9y4Q+mzVLxDkObtuU4
5Il219tTFTglBS4waDdEo00f+/p/bzzakDY7Ma3NhhxcPd6hpmLOLrf5++MJlDvJ
1Hy94FucSAu7HirVICmzOZdWEbeIuZJEUB49JqbUeuFAaxfX9VOk6XECv28iwzUb
ym0i0UhJX6ZoI/fYQffXPWjDMcwpwfik1rOHDvsz7rq4Trs7ID6MDqJT8Sjd789H
/GsXVnqsMV3+ziQmZ7RbrKQqMkhxla3OhTQipnY36PVLH6/eCr5jWlGFxXbkx6xP
/t+IVlLTG3keGNc5Zlr1D50pBgUiWFxeDEmm5O6aYW0x+BbusyJH8EELbP7B9LEA
LuMOwKgjV0Vafm/V8MHe+cLpkKbz/wnQkMgISMa7+f2zUcYZcqEJAYMTUXcU/mLa
osQ8jnDupnRG5r5uiExB8DgvwlnI7JKsQ1VZzf/Yupko85YDvTR/bBHHVvXtdOar
Yarii9yepFtDwrOWQM/HAuxP+HgKMqXwdbOpOpN1EDtOmLhfx25vkrk3dmXMiFFA
emqmg8cpOjY4O+IxmYWJ1mcX+NlGC2Mnsd48Geue5VFa+qUI/PrTzB8ZJCB5X9et
1c58UlkbNAtCPV72PQVVdWG7sL5GBzl8lD5uEalc7nlDGKFvWl8Wd3YgwokF1RSj
/dAqPZRlBKFClQ7OxgM29VCfU5khkYbnB/ldqGa7RcvuMZlVwVRqeRvpGxnBFKxG
IcGyzEJR3zlELk+Kty90bSY35i37+X0OOOp6TPqdcMYalYWeKybvHdFPn+up7CrY
Ci3wdXTSfychdzS6mfgjgfUWGkCmgIJxxXMPF6LyskR7oF/vbuqcObfEgRFKdyEY
nnzGPS0y4LbFkTjZ31E+qhbrUN5Q53JTqZvVcgJeIh0WxR3WBtYszV6hcKb3aDSh
q8LhrymnueOf+/Qmi/1E4DUeNIQGk/uDlBwZdFqOAwiy7zflSJHoEqDnRBgmvOoX
AjvLAQvzGmzVneQGlHO7CD3xeGJM1Bc21qdW+eRaO91q8zuc66gW04ECh45w3nkt
aewJqMJNKFLIrh5aKxm8fhvgExwh0kAQmC7gyAJsMVv5ZMxakfS/5lBq0EsSzkhS
CnjjpYlIioqEEyWg/f/LLmPdswWLfYJgS+e5NLRxoyAJjvftyuFTnKLa/bIgNeER
A9WUpWKcNRxaHWXSyn1UWvbmWQR1nWzQ+g8Rfbgk9ZleqVTROUAYmMfC72dUZqea
Q6QBXI0kWS7JCzQjFhgD1nNh4K8x8QJFrqxcC42qN5CkYXyEa2Tr/1DYEzbUBm6q
EbpRiOya52fThGdqwiFcGDw7Hca9Eyg/+xOQWE+58BRwDUBJvBqC6APWawmuVrfL
e2VExuoPIli4HmHEoYi08KwIRBw43wre/G8+xWxhXJv5EKwaDhqCjpPae95+l6QF
+XKtncnnb9quKW2w7L4mBMqwlgeWAUoVs+wJA+Qg5/DSDv0RdKJddZmyfrXB5Ku7
sgayUd4Le5BG6UQxviwW1IE2fketcWSdilB/l8qDw0WKahpfo0nmkMZDMQ43z7ex
v25Zq2J5wExa+XrKQP4s9U1Tpp/ZkFMuO9JA9xOAiadSvW4rfV72hRBHABsolFhB
72UTipw5zg0JKjIFc27WbkAeABphjWHyHLxDnSOtHcs9PFyaFef9RFoOBuaN/f4f
xQw2Jvnf7hwqravSLWvgSAbRNlWsqcpk+NrjwoHuPCckLt9viYZHzyBiv9shm+LD
1D0e/5QiKkrmlRlHevFBzi2QJXwJgLyNJVBlZPDXSRP3Eo58F32Leh9JhrTPEY3Y
sc1b2P8tfNE2MG5cmn3s2/FOmAYypYtg/aPKnbMNeBBWQ95y9xo4fuqoDfqeXY2W
JZhk6ROB7qGLmJ7HFx7Exbin5RF0U/sqdbesK64IQe5lLPW9fazfxw1FuQijp46K
nvPcpYfX0oBpe7pg1xz82UDvns3fYBMcXJh7bbMT1rDIkSrYUVxvGmzhL98gnSgF
LCCjM+yPPXUmVgvzYEkOZ0XxYf8GgFRASb1p2ChwQ3kKpdBDk+9bUDldZUFZxN8t
wEbgtja4MWa5wmqcfDpVvhF+v6T0aGOfRB2Jj8aIkoX2SY5sHH1MnUQOdS3vJLWU
s/60apBlVcRTyqewd5K+l1D2zTDyYp48mK79u9FrKmcD1uo1DDq3WxmdWa/+P281
eQWkVlN9bNo8asUZp33TgCsNoUmlKeTkEvYD9G/2K5ySPYl0OcCfN97ZN/9uQ09q
GVvAC2egQVZbrJJsF0QORb245n5AtVJBZDjIEhxtaW0lFofVL5cxP5gu3mIiL3uL
/LXCHGGDo6nLZI3H/Zyj9ri0HY0or1XrPwSTbnCdZc+MICS7lYl87gl8xu2Erz8B
XKXYrdLenGb/RguCFTvnXY5QHp8DC4q1VsXSroEo3imGGyqpI6UIvjfuLdznjJUx
0SxjFq8GKmoqHvP1+NVV6r/dQYXINN1zh/wlclZd4tdBzIWRIX4gIsLlX2SWJxUi
RK1YR7Ajyzd0rFbLZ0zAgRUUGUh+UfDXz63DSdHctgFnE9nwHL8lq14C9BED0Rdd
32q+ZA9AUULXP7V9Xtxuh+iyhG/B8p7zpzSqxcEUFdz6/QgRWO9tVtcPepm85FwB
CTHkN+h3d0N7xe3gQI7dut0lBbnwkyQPjKvAuDB1By4VWmfyVnzPWOj3PKthpgS8
n3qpHMYr+o/vqPPEEwBoJV/Hq1hDkexSnWi/BYlpwdjEWqQJdkunEH8ESLA0C+1P
o5blfTKJytdYSMXnJIWyFecdPRla9RdSC6k3UNk5fp+A/VBp9YJZpjjAflAOKDH3
2zvncM4NZvZ4G6KRiUjBcje2smZZVKrQYJ7e9T+dEa5qZuvmMUWwwfPSNoXJ77sQ
Mss3duIVlK8Y7GgLSFwDL8dTR/gfXBa1N6MdXX2JXPeMdLgTXpxExjz4xcj4rJ25
2TPiQOz1DlY1iaHZFQmCllvN1mXiEVo/oxWcRl06YPyaS9157CHivtewzSmwnNMY
YmCv4U04pyqKR+y3Vl1YzKtqrFFQ/r4jyTE+tx9MZ7WfQpdnSGoXYLub2yToRk1m
s9eYfZ9M/EoXX/IHoQHB932WIt96VX3x2/BakQzT8IVZJd1oHSoiQMy340ToU431
aeB35/LB7sPQwtYHNyVDnwqam92YW1ljcVzK+GufwxyJdUFPEzjQuu/TYThdZgWW
CLHi4MpRYL+lAEehdTxZuxBUzm/PYv96R508BBRYcbtkUOH3KJZPHBAEQjOrE034
+OgGBvFhFZQcW/0aZ5BE1ol4ofcmQCDwEF2JlLLej19Porw76/5crMzLImoLpDOk
N27vCzcTXCB/araIAYxIMS2kj5zR0MdkDlwTI2yPRHFdWYDuU6Unr587ih3tIuwp
UDj1daqGzri9Dkwh05k+9DWMOSKk24SQgzmVNQuOfoSKQElsYzAYKNboaO7cswv9
IHJ1zRKIvOaEiKfqRx4Yxwc1NrwBpGET4RX4tab2wKkyMUApT26H/yIXrjRG12GK
Hdu7DM3o2roSv15kRX8V9/lfXMkazqJluhXS38mwhdIue88LZggWO7phnEPPPFdm
VEWDYNkyqXLQyJ19cVddE0Q11Z94IkRzNx3RD3LuszIJCKJGF7Jx72Nt33TgVq5S
nla95G/wowMIBFp4OBb1bbpYyTDtmn1eLg/BJu0N4T9KZuLbe3N4B8cEQ+iz+qcw
nqw+gWc/jFv2aI6twJ70CPmOnYveIy/pZHZx4X7w9s0c1R4fiB9vkaAs65qXRmVs
YuBcXiYJ+vovH57jKEJ9Wq1E9owhGWEeN5h7VOeUGR2CqI9AkmPoa3B8pWToAaLC
wNy4WQ/8uLJ50bZVZT0Wqh/lxKhofWsfGO6af1x1VWLzi2GQ9jCpZO2ZLFYOkrqF
fTbvnqFRPiY8LR0zjn/YBZOVn+jd8yRkSnWpn/64i+xsLqIwMB6m5yBDWmkQ3I0u
FSGbe795WrOy1MkSEaoKcZ70jjc7D6nm1+988Yk+lpGRIxgYfWFrrTK0RVEWhwPy
Gp8JV4g9WsyZ9tKYQHlMZEkIbrg8YnIjeJRleh0517ya5rWYpxuqgSgj6285oVgP
UyH41NRyANrCtxbpX/AWPUZuI22sqW+DuUP03XlD+CRPQEDyYJlaoeHJi/bP4qIB
7yj3amTl1Q+xkQA9uWNhHu0FqVl9RCr/cMgQ7ynSKC2H+tpvfbzPGVbwzMGh0QKp
llO5Rr/IPVjYwsn7qO8K+vycJF3lCjNOXFV+61rT8jKZU6KrBxmQMF5PuCQeW7xH
4Gv0ZIKti9Pw5gU1EKIoqq7enmYI4XSs3cqTPznFcHVv4MGlaUakYgQTXoMTGhHd
nAbCNjT5X5fVzgAKDJDDpUhrK9GgYjcq/gCunAv9SJgGV+UWBgn/u2wHmvfcODNN
y28pSK8sejUBNpB91HQwq8SMR/LYLohPMR+JwUr6fYut3D2t0tv81BqaId2HBgUp
l38or8k1XznttaOda6r3R27VlFkFNtmRVSPvnCLtlGP0z2grZY8yrDp5efEytWyM
wy70dCLbTwzA/OAY6GwuvpAq+XW4mE8XafOmsRYVgNcHDTTM7iXtpaWPYVIRY2AZ
R6BLRaLlL631TgfBBASQhNOOYjWfiNvaJX7R7qaOjWxvd6DD+t3k7xPW3xR4ezFF
v6Iqqp+GeyD88RK1Og9tYOm6nkkW0ymuGhhxi5iKH8pQbhHVXXHNipfDAE7yBFTD
wEOVa/iUXLjJaWWtyEI8Q+N4q21fAdj+TULmtsxgq39Oi3DBhJNbr4oNa6cfyRlA
9MJn1djLnTUX+zFwMQWjzx8AXzJ0h30FT0zc3ZlSXBGD9/+xJrVS65OMtUhMnHAi
jfvFLmcxThS7NZE8lGrRnZmYk+zjgNgLNnUoi7+riAYyFJmnVWrqecAvPp9asLr/
UqtcEsZr9qIz6Lmf5s1VRvxe/OfnwV3X716jAuR7qwsFWPCMwQHZtnIXCovDwKc0
+IMOgllY2KaS7RH0zW1oa/V7PjIzw0bNMihkXE4qVnr7yX33F5AjUbDawndtqoJf
6K4+TLADBGBfhbHSgyJPFg==
`pragma protect end_protected
