// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
IHCfckRpuSASfwkGc3XhMlSbYZN3jD0aaFdxN4k1XW5s4IAmO/qV/0zkipIskr+1j95PYMs9Ze95
CgNQ+pOam3kCBfeJ3Jz8inEIjzj/cWhQcOXZcQj7BE1TPIqqe0x6vX8BM0Y6HtSoJKaoY+yuyYJw
OfyNf4cp5CTURBF0eNWTE3yzymz3DUNEivTuW8CRDwba2Nftk7hDLqWa3uDrwUsBcGx+Y0Ii1aDW
eSkiOih7CP+XlRR6uHugoYhKjPzwTDws+DYbN48eFl6ocJRz3QB31byxPRL9EoCBRkuxQ3qBXrhq
9xaWacmEo6JMKTp1tZxNAilJej0aiDwaWSM0Hw==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
2NWejfLMyTzURXImEZZEIx50iImZsjRWzdVB1C75zRLE5W1ScSVeQ/bjRX5k1Rb3C6r4dKwq6swB
Ah+aErey6e8jOFo16Fjp2BtzfEVJ2TSMHtDnAcopIecJPF3YhC6FnOnL2aW8063CK4olEXR7rTB6
B2jxs1IV5L3zyzJJ26wr/Qw3y2mkwec2R6b+5NenROteG9DyIs1bGM0zmR3DvPYAo0+vexRRF510
HSj8xCg3Mu+hR2Wz4Q5phJzP2kCYN88/oA3wv0CflkczkkS0K2UQfhOvFiWRrpiGWzspBp4fhVln
pvsxodYWVIgA/4Q0phqkD3VNYG9rUcdHUEhyyu2CHIJPEzzHhYGtu+oQGkY4IJ3I1aj3FFoZuEJQ
pXA2ESQQBWhpod8OEcL9+zGL4m+3owR3HUXB1NzEsYySypm/ADP7ZRW7EIVdwTrlXUB2ASgwVV09
/rcH9mxJ1giTe9ovPb8dRctGSf3m4iqRNVylZSy/A0HErafTwhXQ4bfh99lCF0z7yC9VCC5TXRyF
Q8DTjCx2UzXxdLumEgpGkUgdvR+sDM0KlswP0RyXtVTKvqI3PFG6gF9ACiSV0aIjVQHkphnPg9om
hCFlppJw/e46KPKDD0XF/DvmthL/T5ydPmDw51SWgqTlYNP7tluBfVa+/4kR+FVc9RC9roffQbY5
VdUkWaRH/JXcuHDHSTKevoqHG3lR/QJ0DwcdpsNB09KG/ZfEdxT+MHPE5TcPP10TSBto20O8WnAN
rM0k4B1ECgQCB1KmkRzZTOjQ0dyG1jk43jR1MrcUgimx2UxwU4u2j5Tl4Tzw+LuCVkaXnr1sGoZ5
/xycb7A7UpOIhyQQODYgd+uuWs04ymz07x4xDkgof1JsX4jMF0dIbccZsMl+qjWH8uIUqqQqULe+
WowmwLufEv1Prx4kiYh+szwGZG4IYkMYEHWHP2Rkx3CdDjLoq3SQ71xOHpRgrh8YD9InsU81gMTg
m/BvvovRNqnPEy3PCgYBsntwlunXtZff1t8kwT5qioghNTk42RcCUyqk81Nn1g1qvOMSdYTJVXq7
E3/rehFpLRHp0Xht2u+p7rKHMJaPTgiQl9qgWqBVL1h8wq4aWktmZpf7QYX6slldKSltWTECu6Zb
poD1OpoSiYjq3VWIKO33hQ80YH4sltobWi+nag15qntkZ8hDWkMr0JNKMECYIjDs9T0DvT3UwlG8
Bj0jeSirKV1aaCHPo2isOczMwvW3eYdP3pXcpCbR/Y73NjnP5OeVfoTJyt6W/R7E9Jqu4y24U7Ha
xvAft59mcdnewEqfz4rf+4B4NBJHQdnwuvmbRM7JqpfHR0/xYXUO9FXIOCHmLqWZcFPfSZfQcj+w
aqkQhmWstkRRJ5be7JVjJ5qZ9pkthmeUpdLNu1XZrTZfFCb63gsYIm9QK6xbZosbYp7x+vqHx9mX
PwJRvSo+Y6SmuTo5+lMMzbSb2RUWBvu86OORLMVYUm0DNDF78MrmDk3m5KVTZ15iy1omDxmQ3hyt
wO1OirbcPJR2PtOCe9tfPRU1ep6XgtN0Z7P8xbVpfLG30dD2u4aezGjV2ZgkVUbLxHWtZm53u+fI
FSSwSuiN9JIZNpp7Gl3Q5aEzfcjn6qRIAVSOBfKaH/njDYIB0In6kR41GXmtXzSj4nn6v0KRB4Ve
ue77qIH2R3XztMj5F0lrfvh9EhlixBCVGL6yJTaP9oiWQYTrnMlB1LSLpo46SfXbjEkfBsv+oRhV
BnnTXORJc8P6qYl9XUzTo4+B4Az+YG4UjIIIiBUdU0KUsw+H64lGiVssMSqpp+nyefi70J4uAsfl
haf54WFXsNDzF7phIzywh/RxFxhyp2rBF9BT/WTWUvIb65+wZRxwIONZ+akwA7K435r4ht8JI6VM
JKkmZKRPDY5aUXE0Y9tklkHRGZMFml9HHvNVouLXDNALqtPaWd72wqsrI2rwKt6UmAf6KMUQwm0s
MAPPs6YpK3ushN95Kq/83sOGS5dEs1NckbGTWR9fHKTO0M2GM1TIOKfvKL5DWBQSufaVAxBcVXrN
j2t73ygM8N8raR9rMurRgZ0Yd1PvJ1BiFZyOKbKOyVnO3beZKZXIkQr2ikl86pAaA4+JlGs8sUlQ
t6Ad+pJTSIZXDLxiD9yIJqjAUtBjQBWQn7i0Xp3Veuf8AU84HiuKBIYjds8C2ybIyVhAp9thmTJD
cBhGBxdGvkx2lvIyrWSFV2jEZj/dI0pVnpae6F0jx7WqJ6rNw+P9/QW2mpQ0cXkmzc2eh/d3iNFV
t65MefNugtoiMkHR/S0kqacKLBHzFjalpUA9qc1byJUcgBYXIUJso9Y4DHmtnLDb9LoeuKY2ksxT
8l7nX92FiQFruqbMsV6/hnNRX0DP/tQxq/k+12WaCqqzcXaGYVrNh5haxlgsf8auxLbpx+vM57+8
2X8AlIzx29fjQ6W+6Jq1oLXBdnhvC38S5OvM9zo+i+hEymHrDXC1kTYo4u0SKCz9k10Gp3omW/wp
6hJZhE7VgxecVMnltyuUWNWO9/4nut25gsGoAPh8TA1bf2nSvG9CJLKMXXb6XnAaPHCLFGZmBAkG
+m1aAO2KkHijhVJJKwH/+UYuplGyDWJUvWe2+A23Vgwa2mD5/4rYE3LZxno/JJ4dxNdSc6UsreVF
wftt6qy2XDyXML4c4KmGPzXu8WNm93YEfGJSggPs4fVc5hKfQZejDv2Xzi/GK56Hr2IZWSTVAeH2
8oeynbZua29dWyk0HB8ynJtwwwcHrM8F/m//ZJBBQA6/I2y98SMMUgDd+SBz4GKdCpXpGETYPTXK
HfT65PLBc8orzCQJNzCkSMa80bUPzNSxbqbiWwHDGv35fqBLc438Z/jr9qmcKTutIwi+m2Atoov1
5nLJk5b7Kc5+EyTEE6OsQDYMKXmDNxW7ANLGFaanZ76t0Pkdd+K63oN7/6QmUErKxqtZlvei8SyX
bYQuGXOtwfVSJKaVV7NoF8U78v8gym9phfAMEqNgDUSNnaW3uhOnexr2DrML3g3cqKtPlfRvgD/f
qx6vzfMoYG4PPy6JQCgFuW2jG0nlYoml75UOYN13kX0dFQyaw46I8h27IX+q9JHwXn8NVo6qIW6r
7gzFE3pzpTi7nSQpYGrA8LudhryYfbn/oGmjmpgcQyi0LRWZL9H9jTS1BiOD3p+mK30GBCGCnC/D
hhaOJGQdDqj4sNRvKHe6QSZb8LhRP6+TpTpHcAzyLA3DcAIW2M2GuhSqLPM6mmOto5R77XyKPCbn
MifbJWwdcbB18FDipHEaJk6OLuqqkaCBm4uBSsm5GkdrlMsibIdzyFiQW/HTW79dV40NKnp+G0z6
mehqkiGRywauoWeoEAuflK9+T5x8BVjgadIZhbxCiErcVHbTGj8SRWOYQz8xduUb6kCGqPbdM/Qn
PKn31N/9fuMucSnmJ40eD2Pj4/V0A4GudiB69i3IMVqLKQ226MaVSGDzlW0aezEVjaXzRhx4t1S6
fC21V5UCfbejaeNeI6swS5zkBT/6DPCPGsTkSfIVL9+pt+HOxJBowP8t9QI6n5cRub03D5AHot20
r7bQlLkkwcttoi9qLJ6zXwz1D5A0QhfXrYqqPd8vG0pwZSk8/1/MD6zynVgkgi6EbJETP7NNA3Ca
BUgn64MKlSBQ+QXmp34DmVD9m6k/7tNct+99cOJ/a/iXfq1PxrX3apcdu2b28335WWS8yOFL5PKg
NB82/k9WyCuiBUT4J3GqMhSf1th/u2ByA4sYILnGnvIWPB51+VEpVuKwd0dRIOeMKQ6r6ZKbpA8U
o8D7uPm62c+s9rOUP1AVNHfi6/XGLRTsT2vKg4cg0Z6BSKaBmlLBebys8dnGt8LheaZZXW+WjiUj
AZOJARt6Kpt8e+zBYbsU5kHoERDUGBZU6yCQ/SUCeMtbJ/rPnPUQJPz30Xjvn/Fc5E9U6ff6hhEF
JpvvP9aDZmeDx1ixa1fAv32849/qnc9eG8Su6XfAy3tKZKF1H0pIgPrX3+p63reIh5MubcqN2zJ8
VT/lkdJk+fxKjy3RmonXsHX47iD9YaU/yrV3NnB2LSDtwf/mSijr99hRHsg57IPx2xfVxxl3Ward
iQiGEB2/CQt9UqixtuYRun9SyDCJK5Zg0z0mZ5+d1DRiRnhlZrXk3tN+DzUzcZaq9/iBzk8f7Y0K
Qm89P1sfCm8ihy7Wop8pUxNY7/9+VYXkRaaHsY4yJQNLZhbIiyYch1/8FXNnH+xWkvyDXcy/Lux+
gysvXYMwMkNzJYaHs0hnFsoqLBJB7wXTgaj8WgzE79dfjRNCXkrKK+88ggIo6tSUG3myIDoIZ5II
eKLO911vP6AxlHOh9TG+F9GB31Jo3ZcKaspk+wrP44L6A/SjjRYu8BlLnEkBuG4eekq8dYjHWLfD
ufYXeN1W3fL3mh7o2HLKHAmNZcQ/DLlWmzOQGJljRZFpkZybIbAKvhwSj98t5LnH43TvWTOx9aYM
DiDMmNy1938p7ZE28Ld9NuZM9oMJpKuFy3lZiyFVg8AVTHhaQ5lklSdMC2UwCTRpV29Gng8XIpUa
j0N4BLt76jgLckC70rakJrg3RzcI7e3ZS9jfywOTPC0EDTgR4weXHrjrbv9OKgf+narEw+qQLV7b
Ow4D2DIR/qS2g6wajmORyuWgB23gEtum+d8e/P8LvcAJwMpoVst+U9SFBS0TUEBntnJb9edGAoOy
sbWHcT26hgqA2AfKLZh8zIx5EC7EJ2XtRQN2CcX/Ddwu66hVWdCg3n3wGSqGHVSyZLIHdNwl5/79
WcT0kLjXXuLV9SyaqMpAKNjQIUUM96So8zTPsCCloSdhv2ADMe79RyBCcHhX71whz0AOBwznnQHU
GvUtxMwe/R4fKPdgBAzfHQK0R9jvA8Zj+dmLAKI2uI8k+gF1x3TvVsEIWC1SJ0KkE8FLMqRT1quI
RcYl1sHcRhQBmQFgK9PqHZYzAJvEsnhGwDkBI2BD5lgvoi1exsR7OW3/JibD1pYidbutWTirhKSt
OFo4Vuo+HGh+xU0jEe4R+LWUNmXuHp5Pcir57tLSgkjqHAjZveai3SPbZ1wl0IYJKLjhXCeHuVz8
6rTGZyYnxnOqA5OlvmN1e5tj5eob6YdzMQyPRiU4JFFKp/Uq0TdMScuGFvMFnOZl/WhD7QgDxNn7
ndwIs44qj4Q8I5W5QTzcQkaEHmKgiyHd7A4K+rtkFqDaFTQAy0J/6jS1r9hdacqMH+MD66J6CKp/
/OcE8FOCVX2+5t8xY3yB949Ul08QyjnKMf/E7/0QQe8LgXlAFphUH0/eOwCTpszzH1tG5Mb/WCvn
eLR1p/FF3ytQlpTYiTx9Qw/ZqGpc4dU/g45eVpVkbVDbCj9aeDNb51M9shyGstVWS3so7LhNHlGu
4zVO5y9Az0Pr0g3h9mIop8tNfObTrdek0wfoaEkhQ7GnMzvSLnmoneTQzZ3PriDldJn1E5Oa5Bii
WhcLoKMHPN9uiC1/IGbaLH1QB5cs4e7yY5CRWKK2EWzQf62GgPpA/0+9W1Ve0t9q6GT8EuOKgeNW
Jy7nfUR9D+GKH4oHlJcG3AHYO8vPz5vATTdgmBVLqmZj1bumRVH5c4dv62sS6Tx719xTVqcE5LXj
HsSYE8zGvKmAa8hCAtOzPpulW8jGLKBn6OlmYi/rp63CDMgHRFm5lJmMpO5kD6Earf+seuVUN6rs
xHRwv78Ncd+/XnkU8fVW+gtq85oKCrMubQlcUlR93906dZzrSTDwCvhizjwZ1Kx4VAv7LzwM2my2
hdSHbTrb+/GPF0rYzgNRdQmzJokIs2EsW2XxHYjeMwhqkXsEK9vs6rkbdH6uJqU9mbmcqe/+h0qC
tHey6NiSPMIzOLg/yqgpoFOGjnfKFuIPJbMOElrBwCI99rCqwXP0iJvKQyWueeMgK8v5pcREJt4E
yhnsBNhllIclxHsrnus8czStucPftJ6N5paJG439hI/NiRpYguwkkpPoCDxYSm68+qXGxcDHOHwa
huwPxLl83zBkW3f5ezz1Lb0JMa064cHegCAFMeUGgWtBIxnFPDw+LV8wuNCdPHpb7l3+Rmh/h1H1
KxQgHf1PI5R1jKZejlpOe1BwAh48/UTBEspROaJc6BLqf9g/C9DgWuvFf6eNPFZbVTAvEUKJhlCt
DeM0oZSLJiiaAzo4/BXW+U0tUh+O6ciV5PI2dJsSw5KiWeyZMEr1CF1IiLdLGXQUiGm0AVaQoa0C
7+z+xS5xukaIWl88Vf8s/3kGjZS8Femzc7ZH4jEIc3Kr4QrfXXmej9Ru+u1Uag2EXeO+1uBTP2em
sG81YgwNcFymiCFroZgm0cz2me0KSXc9sZ1hBWCaE4pQH2z6tpIURaqHD0xUfmfMAmFnbfY/H9Md
A5Ce1qXUAhstLEzZuwCRCGaBGUXTDJUVLqLTLa30GLdFB9KTTz0NJEy09Y510lq9jKtJrsHrSiMG
OxXKlWRj8yZXBLCFq2XVaSv3q6VMdQwlA4Rre7t++CQzpZJMm3KGySpi60KeIbv0PwwX/9i2mgWK
6OCr+y3TVtcLvChwMf2pRIyQCGIQnycTm6fdLLa4WT3WpEa7Zh/tjPVSdG8tV9d5RhxEdVLKY51L
BV36dxSWQ/p8J0deori6EaqUIHH/8iua9u/HpYNeX+Hc4KOuGYxBLjnrAOoI1Uhc/ISljAikUQAi
tVWX1e9o3pcsJ3tjNny/EC3/uM9Ohn9m/xWyhkqNMNzG/Suf+JTOK2rnpxrG5jI6nXme002QKuT4
Yrlqs2Jqr3MBAv1p+K3rh7y9BaCzmtllJh9PolAIRaHFL8GXp8/gJ6/YYv0168LoCJ3SSLdfyvpw
XjztDDQ+lyq6jRFvcq8av1iQal50Ei6cek8X8KK6Q9sEXDteQ06F+rpGObqgH0bLwf4dNvTy7P5p
P2kxgXvA4m2Xa5gXDh+0S0aql/U37Av0UopDKCB61islJUpuvwlw6MVuKvB4oouTRndIB/DqeQgV
nl7QCr21Xm6M35q05zTlsChSOhYAlZLCW+oa7UYmFtq4rAayvRc3Mm28So7EW4XdavBU/CAG0XRL
AaYHe2nYK9Iy7u4r0JWFK520w+hb+ktuOfXAdyBm59AE4m1sh8FHiYpENn1SDcaZ7FBPQHQYH2m8
TcmMdkgywJpINXQ/9Sb4JUfug+w0ZXZHf2Stpcpjy0iO/X8/1XotKN4UvDMuYPR8kQmw8uyrpnoU
2YfHQVVhGhrKIiErWL4LOsm3/TFJy8vBmz+yx/8yJAVbErT2uSra2z3VPYIAwtX7QEWEYB0BGIin
HKVfGpCp7BL7eLixPGF7naED9HMWrbX3FxmtCqSRz+p0IaUek95T1QmkJ4hfB4Z19Ze+8wsqs6c5
iOb4l/rPnhVl2c6gL7aJwGHnUvmtx/jRofwXLAzQjSRoQJ2grxnc6bdfx7HWZdRu7ft3MJDwr5Ds
wVTDOCUpRCNwn7IXJ1Y29NiTS2wBuF62MoHXt6C+Hll+hY0Ce6kSrlsoHEZT8FHMLYrjAE8X4jfW
Tu1aVFejqTALcda89hG9Jf9KkLEVugS3UmVeGJGwKN41fLR+hSIc1tRwOKk3RbhVRCK/uTM2VuTi
AvxZyWINSjZqYRvGyfwuVkxF5tUnW1+8e3G4MlluFYhBMoX02kUASLMr0eg/mxSGZ+CI1PWiw/gI
/L8qEzYDOBwbJ5AhPhLuHJUuKDmaBV0X2q8+GreVJ9qjbWezH5LUtGlY8FZt3ERQVrpvhgR4i6b3
KkifXhiGpUDVsVtKiY+4p1QTpnE5NnLbr5Kkzej5wu9oarUdqti/eMZpRoRxRjQqRv2N/sWXyn8C
uMUDedIuD63cHCIfmxuSpQn4dy6itjx0s3FZRKdw93eqtdHIo/um0DriSXR0OZjMsDJ4/vaF0xuZ
hDIbSfMBrQ4YnfuR/9ofQlHEB8X4HpN53rGMGT59h2i1SG7VFokreuOI6OWOAzdY+Olgn64Odc4y
OM7lEjGL4iKdHoS/2cGV0Wr8WBgk9wRiyqZh4J2boPRNJ72GiZ6BxGz3SqwcWBATApz+qiSi0rP6
IlimvtQVWJTNNU5X95HKA371a9bBXV/Rvrz3RPctKL0DsTUxD0totHKw5QyYVmpB6zd2NpTFBUDu
88ZKbcBnOj0lj2W7ceIwu5q1DQNPbM9IyEOU5Oxviec5N8Sat4UisbVlpjSRMzrDo/P2QXcdlsZh
tz20l8mp/hEQ7dBYYKWho0C6MzcRVl/OpPyU0N8gPCjyRzQ1DD1E6wE83ZXw+7L9uM9OQ+92nRGe
gX8iANSITr7acM83ZjfxtSjCNF/439CnxjoEPFytLeey1BHNYiL2IqFCzvYpeWRsZda+oOhSKySi
nGh1qd4jTBq/iTgNo+R5LVqJc9JljA0pL0vjJ8vgSf7puldwgGBCJI79xPBK0gcJ3nJOR/3OPZ7d
a7nafPnVjzrQXHeAveJi2Vu+y+2do2s6mRhTePr/3qUQqi8qSKy/TQPStWWw5R4F2dRnkYNSmwdx
F+rMRQO90DhXw31CTHsdvRBixjBlhnFZlQFBbvYdZN5ucpf5u3g+WpEEZASN/RM0ZcpLzfY1IAJR
zpC9r1UgtSjisHTF5T7KirnD05LR28UedhLj4DqBbFhjDOyWaZvMQ7icDldqAN8Z+As0Qib+JhLg
mAp5BIfMHoX90scqyaLb+K3J5vWhJ//e/pKzNfWdHxssjNbtRU1w3jLz2KkXkoJX49yeZw303TyW
sgg8lwdI0BAycAYwmJAl8aZCQ42+2ogByUpk489OUqMRrCmxkqLd9umTbwqWsDL1VlntCFNO4eYP
of38nGMkMrEDclUtq/wCIuy4ozHGLMqiYWHF/K6JQduX186r+9KkDdPa71C1PlHkBG2Vq1Soe2Uo
YRCfG8c/WTwLL/n5gNlhDFHbVyPEiKWQxmRE59Yy+wivzHvyWTHK5E3JHApnTVISleE0rWMnv08p
2gurCAmZfILI4xj0AURzOo/TCEdG2Hw/B4AkzpQ433qPc3uXyHJ0QHqNSAe+IyW2bCNZXx+ip4CB
m4YbI2yMGevd82kvcVHSXo29ksFfauVYktZ/lQA+mfzvWvXisrtOdGiWKmRtiW9+sRUW8V+vmvFH
vbv7EYovD7igMT4Th/pRRkDubPlkuQoVdSkeljkf7J9ygsbToCtrORMIhENsQY5zOihIs7vUhH5v
stBlO0fMb9UbZ2mJVgdQ8MGmxurLbo5aUAHSeic9jpP7ngyfLgQjaVGEt7ylZxyn2diJfUex6N70
UjbcUKv+xh15JdPau/nbJSUR4fDc3RcMV4i2ecWRteg/qQq4/qepgzuv7eNrOurf4n9uku15romC
q+cPwP2PiNMgAZUT5NOTphZNwDGkch9ed6a7b8LVlf59BH0L480Co3LYwh1fkWRWSoPzyIdTpHVz
QJgh53THkgIyTMNy9GfCiknUyxzP5WgkPCI+LU9yHa48mPx9JpdcThF/zqvDFaJ1PQ5tQ+yYl2lS
YleFEZT+EYeAfqkFddDJIAUgiXa9E6DV7AZtqGbbgM5q+9DZ1Szk2HDdgs+3pJPKXU1Jqcjcs6Q5
OEAyljs29/4PkFOOG7dpXYuLcALFuw6sGKwTlq3sI9aIE8K3UT1h1uxL7anRChXZlFLUAay+I6hc
Vr5h8It19n5qDNMgdiZtcIX/VsH2sP+6T5Tl5RFuS+0ZnGxdmrmVC+zTYQuHCUSivIPgxF1UU5ws
ZNLZ7CQ1aYFa6aV2fzuHEbtatTZjHH64bUwZo346UaOr/aGR9DUGsAJKDz5cwkjf4nDHrf9sRMIJ
zV3axogq3pNmyNqfv6gdfG2TecZqOPEfyPPPDfGnTskSre9uZCFKo7zw58oQz2bkCCEpka7OaBvP
QVoL8jVvImZbcla3/KNEIQB1n3xQwNaI52pXy0WLZs/e5dsEAV7d23pzkxNUEhiChihifaC6prso
3E5Z12h806eSdtTqGSyQqfcdMlvf0vA7Nx0DfGecFNoTNVY0CfTpGX2feWmsCsm805eWejGrodjD
S+SIFQAMuoj6hwN/9S5MLKkKOyL5nZNlZB1dQaXraN4AzCH27xDY4o6b2WKSRTw3jpoTHSO/wxu/
LB1xJZJ9LQR1cWok5x/C3yMTh3ZmXFJcxAmd9JF+iWrTZ8QfgBYFx2yPt+baaLpGzX30zKpvLq4d
CnFiE5mauskwSyVpvpw4f8hwGkjvPKsmkPasI6vrhxaDX2vlfVWXxHrG9OFZQR+RqoKlG5zuY8B1
58XFnjf2N1pmy9oCSpgB+fR4osBhnMuHHnB3OudKl2RPgIT3haC8Xzey6miYqszQ2Eo9pXU+J2+G
SxlJVVAldH2Yk7+gGv2IT+4GF4umav3onyfkjr01S1AXWltdTSX/xybPL/P+hndXbNVmZj93ZlvB
d9P/0DqGmKhuQbCZ4jPae++BJtPCkQFq5QB5gbMUvlqwqjR/GamjtIigTvyuoviOmz/3Rge+68/h
XGVHLp4o0lzgsdBtJEARSvKvskCvNaoKiCgVQZPBIZIQhE6xlUFBxHPEU5pI5JukY1IBSuyiIiaa
Tb9kygwAjiekfzfUgY+VEQoQnqcyWpScpyY9QQH7DLc/Dt7aLt/bAHvOcagBnjyHdApu20BhbDVX
HXTu5OmswGH6zK+OO0RCpizFDhz1lXwjDUh1dPgegcUFiL7I1lqWaTGAD499JQ9PAM+scGk3+1x3
hJSFX9BoBVECg18qgJM1G6rOo0ljGLN8HhHDKtV3W2CuoV8iUmICkfMy9K2yGqOvKkLfsj0Ewf5s
84zv0eu1Z8NvmSZJJlTewIkQQ7rDDUpZP/m0NMLgfTwdOReJkIDEWx9c61fQC72RQQc0dH6ghFtq
YarE+GXMycVIIxldqO2jscAHh/V5v5vY+3IOmvnOIPz1L06t7nE22yYJkNW3bgcELPmjuMLAoBXy
neRrTesovsQ2tlOZLkZgaY7E1yFolPKtpmbG1XiNbDQpvJ9TVAg/dmT/dR61HJWdJpOhKjFjVCBH
sjeGec70PhGbUTFGMjQXdka1mYYIPMg5TTEu2uPND1/N6RDDelWC8vqNIdTQ0ZXgJo14YJgYb4vZ
jam/qr64XGJrvLBQ2+RceAnFqzOCU3is1Ur9IbcYotSGgebHIsHi4HOJcOGHx9ODsRv+p6Hvl0HB
SLgwuH/MWsNcq8HF+fy5Yiaw1jOwvDHL+jmLJtuXFTcdJTPvq5zLXxPPDeZJaD6RkAV6/HC68HrC
KiQSoWu17IcS2Ke3TcRgczBHRCgd2TKWRK8s9vVNbRziuR+vQz9+EvB/1QOsmI5CVfVWw+Qfjd/d
iwJ02AWHwtyQtAyJH2n+3hS5tdoYJh2tFHHZi7FfQ3tSkAfUJuaNLtMVLGpNpMs4Vbi5UxCEeiZH
QrPkGc/GImprEpju/8i7NEb0/cghCb1MwXcrzhjZ9tCer9qGcoA+z0N4JQ5Bt//kIURoIxxPGCiy
/0MC4XUt/LObZulW1r5hXS2JnGeNZ311+qGlFvTRdljunLkml8Ax+Utrh1Q4BHXHkQ0c4Th44wll
4/nd7lU/xAVEcYlQRYL61Scbhpd8MgUCep3f8KP/3PnxI6tP2pzHMKJ18u5uE3QuNCI/x3FhJfMs
/3QbPukl99enOyRPhtOo01Io5Fwjap05ZlM4GegTg+9vJMRK91rqTNzJvClslCYVtxVg0HKXiwlJ
3T3exus8Tf0/94f0q7V8UIzfOQBwo0TonHMkRlZ4XP8JQkqfD9Qfact+Q9+uU0TDgy0fhj2bh9Ap
8Y9DeLGml03grG+5lwehOSwuFYjYgXZpUhl0dEflBjG4G+shHQwXHu/E5sxy+FFkWlVcm9icQXbQ
3l/xBm1XrJdXJJRPN/d2JPh5Gw+P63ANSyV2oCSQZ7zSqIJlUIiTQ6e/x3hi31jHmul+dsYqyMo2
/E5yPl9HV791btzFp2yV9rRO44vuxvFrUMfDR91o3k9y48ew/x9dPpAkxUIQROh8A5eqZ1glZQlL
agOIUy6TYUs6REzHptViSjkIKTsTiCyJtEVaGr4Uqsxk5Gfsi3jdZzNhpdRoUgyyQc03XYvyXeuE
vq++4VEo2jBjB2Wfa3eShiXRqZPmowH/KcYs279WQXN9fAdaKz6PLx1ruq6RGEWqyLailAF2oHIo
TEHn8zltEioX1C6xhilyUfOakqEkQr4mp2hsENeM6FFI8oKShoqmqndOyz38j00jn3tDx8/i+W5G
C7tJIkgHUiQ1nI7I5YJ0lFojnrBYeVGLs9+6nV2Et5gg/nN/dus7CavILI8Y81LhiNMpkf8MiXzc
f5/aqHQqqkXh2ouRTRNx5oKRd1DUWbksyL1HOpdKN7YV/uf0ztDG133JJRGx8JKiJ8NaDMVpswik
KHd8QoFIq2Trhs/Px1PJenp+d1ie2pN+cXkLsy3wyYt7+jkIiW+LW+mogkK8ZLIj64tMbJ1lvfYa
q8LWhvx8MuzlYGO2JJ9Di81K1UFXDPUI62SknnUDCWPrmO+/KlRHVIBqM0x7dE1Do6H8dnniOQ25
E7qwRhu2jWZVF3Es8xc2CKNsYpiycsdnV7SKQHa7v8D2Zp40sn62ShTctfkzfY19gxMXI0LHdsyM
0rqsbg0hbNEAKo86TUl6ogjPm3uPAzWF97AMMITTG32WfJqcF1X3ldOaa6H/gbQ6XU1p3b7FWKly
3NKXbGRD/OWcKce8wAVJzetB4Zj/3PU7zxdVrpoMfE5FOWKLkaftiMRHfnLS+YcT7JY1fNO9bMMa
fqsmRvxCBak205Gd8Z9CS7bf3uKgvdpyJxY1CwMN2qowm0yWgTEo+ERljREIaVRL1betgGKmPu9H
2JbxDeEGb+mPnD643udzC9r/TCjAbLaKjEcJ2hNxUMuUzZ9A4EcMY4IcohPQIvgN/h7CUtUMKlzx
eKaigUgmXsKkCzzCA4Y2MhmSMsIPv3xKrcOVvWeUS4cEEagrTz0nG69KI4MLG9adou08eKDoBvbO
F6ougJjnLvL0SsfsbYVY2jfpEMH/CLfOs0S/1exKnXgWUC6W7YFenPBgDIcsLBDOvPIdbPZOZD0I
vXKHlk2vTylv4U3RAml15TkOjpxm26BG2xTKRpUIjv/WMDjB7VLK9viBHNyzEnLRqRJmSKppPw7L
Pb+Hov+VG+b+gVWvIjpu/n8Jq2/uXpQow3CMYm4pQwH+EUWTLDh6dkQGZhAQz/pcONDfx875Q8Wu
YA41f3Uu7Fx43aZ7qnZSfTx/5YoCUIOo973jZ/zciaSbJMH031YXrFhTADytjOK2K9iLu6Vzudj4
xAIj5X+RhVkBn1DDdPpvZAEQOa7+t1lMwJImn96KPgQsj8ZrSjTIjzrNZ4QQg6cEueL2UiEDFZgR
bY0BmM1onj63tF4jiQqZoibZMCRVPs66AFcBgD9F5Q5mWEpFo6sVWi1GX9gwDiB3nfLJ6jh+4SAz
hJmfWjInn45LR474ys9ivzM+A0folzus6jviGNWFnX2mn7mPdf8Zd+bgrUVgQAjitC7SE3Mf2D8s
nXd2GcYB6tiE1UJyx5KhhJh8S/bRx/s9nUnGKh3aXb0gKpVBXnt4rV/twuz6RBMtX7aNmAi1N2Ai
ntDE1ivV9GoBvqwzKXKeB65MGvYs7tQqJDH0dD+ZlD04oxYlN33AmZuQCdjVsD38rhqe6w28lZxo
sFg9wQCq5B+UWzEqwMLw6y9AG+XZz/RDQfY30L3IET3NR4hLUp7+6DuZOyl1rDcuveF5TyT3QwtK
vfv8+3UveW+YB03NdCWk1H37dO9zJhvfLpHUMeH0ExAVr2qfLchLgsgmmMQ6dmbSRMCEE0aLg4ai
BhfPGM+zWdmd990o5beN68uzTMhhT1gJTLupk2PztxeiidJVxU63CtE4Tksv0C+KADPJDIg3jFvT
FVFqhfflXtWqMEk1dmHhL4WVW4qmTE7u0lpOIVbq8mdAyJlFtfDPXaeDAjyHLHbQTcivJoyk3AQv
bueidk63//twra6h9FA0/xK2WNMdlVp4o1vZ8vQ1hP7Nj2cy9g4r4bidOIXuGABpISPO3mHG4bkK
HVE2TXhPx6HyM/vXtb1hZZXy461eTOCXQuvom7Rwx3LZIL1ledr4kwDPSne0xU0+jnRMB5w7QyDH
Y6aiWAuHwZn2ozpW4aV7tyIOoSBzkMCZgphXaWlEMP0mDxB69um4wWE+X/fNH15Q71A4LMJbJKlC
bWA7wLFOpka3bwHiJuLz+t8pRx75n1ZMK/QgeSSobik0NUBI/Ye+BtuagQPeEZ21DnBW5rdw0nYG
weO5XbSsKceGg/259vQWsTn3WoVsYoDD657SI3Vh9h8otBIw+GE9lc9E3mhQS04BsW1GZCZAyefe
N/4qQLEKjiVAfCZG0bE/aejrXEtODQDXDLNRKsExogQc+kinbS3pbfbC95CQsfNNdfxg6ozkGz8Z
EMyJLjgE3BmYKPGiHuN2Mboqq3NUYDZv27kxdh0srXE0G2Bdib+iEueTIFmDLWWZzJKQatyMWbkA
ZEIkvHCVg2tqACcUs0pEdkdY7JEhf8XttTKNi7uu5BBGw6SQ8Lqr8CnVGw86mdJrZn5vrB8m09mK
BNxJJKoWnmq5uVCM5Qp7j54vTFo5en3xF92vxi1PENSgbWwcD6OtA5jpjcg/ZvjW4bnEWeUlpcDX
/RXOBcGpyoVHjtZNDnb2NfLSdg6K0wwhSMtUdsEmoAQg0YCwjQmpRoKOo0UrMn8nj4hauKWmHBmS
dSfAXgWuB2XKT3JkuDc872fbgIjDqfStzGIyCMvV4Ex90FQ/k0NL2SpnEsvcbB/SZmrVRgcJDOvD
4J2SGmuT8Z6MA3SczxLgs6aw+6PmPOEpWv5AGV1x9qY7Bpq+ZHSJBTsxlx0TvXaBW1uydFnBf+hw
8RgNTEXsxvll7kAoSXkYhyXVIWmhb/d+B9Oo14RfM3Z+Eb0Z7qYKy3NXOsASkrDxyPbIW0gcmjyI
sxL/MRe4WpbfV6mzz7wRZ+nL7EP/4/1yVebtdUztoLsnERgvsvfRcGYnSd7WnXPTpggjuviTHQsO
JaJ/exapzs5nNG9UFQH9bZG8BNqa2svHHNWy3TR7Lb1+M+8Tfj90aKQd9BQasXUFPgPdkhgKlCDc
rUJOI8mLMNue2upXNvakUp6LSnyauAxJ8ruD/thaQ8JGWGeS/+cLQwT42nxmZ4AuEc1090OnCRQt
Mhp0zplR0ZXIO/YtJZhPfO6YHiQ6J6joEveOUChGqOw0SBwTwhWoQ/ScPJzzWQDVMoVLjPufRzHc
fDn41AmTcs6t9IX3gm6/8IW3SAK+sbiiEIYDzSIWqDP1vAEy4YIsJsq1Q/KAxSXz3/CicnAjk4kz
A5TzmBE7YpcV7V/6PdjmWqmZ8t7agMl/XiI7ZnMbekGWeqV1lXVcEb1MDXKBTXF6lE5bwtGEjAam
Z6R+q9pYMhoRBcBl/HNFwJPGjRkN8wYIfmkD3yR+0XmWI9doJIbmYx0HW2uq6ceOmO1ULUShExTk
C5pgdyy1GOAhl/siNYySIjSYfkbkpnJEir8jldwgCDrhSYOBinKkK08RcrqDWE+uR9T4xY6ipoPY
eUea8PyRldQgQTg9/hBPSSyUGiXWf+/pE/vrQqt4HSw81XRy2Qei8Ffw55UUflatDueT0yJPxEPO
jpJ2Yh4GTv2s6PU7bS4gnoXjl5ZAHCsSdkDbeZQdEDgbBJ6kmkYtKnM8w7j5USzEMmrbahXvjank
1KbMJpnIEakMY6p6XUwThUlNIrQFwOYaQh1Q53XujU2o1ScvJWSSerC8zcybYpmIzifyK3roxvz2
h1DxL+Tg/t7b4VX8Lb1hyRe9CUEMtBiqK6In4ZhWrHQHfqEdq2YOjCSV1w5K8L27Dh1v6MCVimg8
iPgHqBPWBlm31goMdB2CMCIZ8oNXchGfz6sEeFE1rJ1JbgXcSSIwYz4j8K6jqJgFxkP3pLUrULvA
9KniwUlrzYjKB8VO+dpugJL9CdTSh53DtiOEz1CEO5B3mdvxmh+yZ5ScNT/f7p6MDihB4blXt+xF
jreMbAtZ6Dg6HNnMBNOoFW+1MksYu4yb+l7/QiSxTCAGsS5I+PFzCUAFtoCYjVN6snH6iWpmiCmz
DRQRMlNzOJQDddFlSDdG/afA9rpJd2keCgq+kCRJ4lTzQBOj6qHRfps+RXoCGWD6J6J+8V6OTWV4
ZJdrg1k9pnViITSo/iptl4odsGrGzM+a/cIQYBDdcRELMcEdMA7l4O+eZpFQ/DHvJbqU8Nz//x4e
RcsKgNki0UPMNhzf33ZGrOZ/3CV11EiHYXcoXtlOp92WTvhQcvy7ke57D0JqaZPnG258811hqCld
DvA6VcmJ86+oGQpuH4lMhTPtkROmWL3ixQNnJ1MELxIB+E5BvbQf5N7jwGpL230ifxcSzu+6VZ5U
3Y0Qqv2xGQ5kQ1/x26MlPbzzJbzCwXM612N9bPI33afYaSYcbjDIFB2STbkNp3YA5BZ1HIhFS7GU
m8qaektVhC5yIdctFGGgewrabuCdjIcZo9UV/MEdHU7qSs2Y9EU93S0W5kav+6fyk3LdVedNmCAa
pCbm6UVey7yqJgmD0AKUE6Nhl5QQ526lKrkA82STawMf7ZU2KL7i8rkTy3XmBZOT2AkxGsS+06fm
jt600iQM0Hbq2mKKA2jEeFhMPTyrjQJHSNoUcZNtFa3h6WUtCQSPRmBxil6ydmr1o9BKmkwEMlCi
FWhXR0IeCvhE7PUtDsGMN/XD3U31QdX9gGuEcvPMPP50Ca0ueZzYhDJLXR/3OwS/wHg2Jm5OgM0X
NapYzyz+E+wdaOvp4DG0A7re2EqygUZwa/IN9DZzDgDdpnG6+JQ8zrg6c/swmdCRNHBNXr1L/fOi
aAApGH3lGf8ZmWa0dGwk7aVqNvG1JgYkbdXerENcuUnGH6wbmvOzkN0cVMUYnXD5SdSaeVKMdOSw
+/P57trEbjDGQD0E95EnjtoaFnk2DoZgloZez636yCc0wg18znms+dftnLNXKZ4KWOXRlCd/gZx0
lgnqcIiGhzJ4jOe1NOtpewynzaJqQCpz1VCmuxGZ/gUQmQ25LeQOVWhbVeERAmpYmqpdd2i5p2TG
oGoMi59OKBLlRrSBaiAnsa3gIHBcUOt+YcCnq9F3WPKdaPUSfnwlkAOjZ3v24Tj5LGRNT23+jXZF
Mr8XuwQO93IPlGF/nVr9Hgr4o8dUvdCRqdEsdzqn631V4/n1zw7G49c7qbxz4XrBxDs0ynZ9SmG3
pEmNsqTZ19BD8yrmTiwwc7y9pEgOxlsCfhXrJUA/KilIFYlF+n21dpWubEXy1Zr/qu9fY+4G/eVX
Q6Ucm5bqnWeItQE7VzwzcMX0Ds8StbiPtH5H2WlpvnXB43ew88g0OXAUWAqZKA17VqukSq9+6Qdj
tRDfw6UfBVt5ITF+a4M84cBimj/amPPsLO2tP+B6Qd16F3eLnJG92EWagCAsWC1w0qGQ+/rn4gMg
t8+h69drrZM+e06mHRiawiAlrUUyBF0/5ekfVVws24XqjGc+rTQDXhLlSEJg7dO1jwdBNm/5z6b6
T80zKpXE9OXGR3qNVYr09svRtcjVB+6gGJBSC6w8alKrM9+JDiLCNf8DMhNpn/dCi7Z4gYgW4xbc
seJDoj3A93N4rYSibTZVeb/f44T26rTV6k5WXOxlVFF+NysyXHMtZmkN5J4akmEdZUevTQBUFMcC
4/iX1+fEidyNRloQ5MfKi4QvcmxO6/bMzMu8QVl2Eq3MPR3yr70bm22e8lue6nh1mSALz4MYVwci
T4geJRsLDBlz0D7EG+6nCF8Mw+tXGkAtWCWJN0SIgDgLxFAeqOSvfcdlEU7OaiT9QlbRHaT/ZVx9
cW4yyJs+AKlnOF9VGM/QNedXHz0ZpdpT+pJESCdOMvE/eDOhdUJRwc+7aY/o9TWuqwSRMlpyp9Jq
yGmEiFGJs3Y9A/A5n+QKUXVgnuZ4y+Leq+yUwswIrZ1VFDLR6x6RMyQRGj+dtw0S/nfRSqavEBO4
agabcn5SNb6c55h7cORy8hjGIPQ8FprE+hWW7nmGPOEPBz3ju/jc8PheM9D5jD6njexvVDHeFOx/
eLUmXlf6a1coq1JOsl32Ll1Jg45WerrcoJucAe0phmulTdO6o93zsFPxOOOK9+RHv61RfvJBFK6P
JDN7/98MJdXOq717eJOvFovk9IV4HzkLky9poUaB8ivF9UEEdUkOw0XteeTmT1hOp/aBBL2ONUut
hcPBeMePHzA8O+efuiG9mj4MuYrUT8SvjRuw1JUE0G0VGYe/umXknNEEjidw2Nyf0e/S5IEwV6rS
oUm+Q3UJunV0mbaOQeMXAJVkH720tgk2uy72uhBDk3gd9XaNara3TswyY/U4kTzMijHCKOl+Hn5V
KcJuJa+NLVzXOstMpzlcjBsemY2pGapN8Vi/UD2JqPXF/5nbM4s4Nu/6LgDTzPgJwmfdY/Qu0jiF
kmJBAVx9tERobY1fY+ZIcb98eirAI0mONDbqydX3/xgfWgHmcm93roQ+M0O/UWCzuqUEHlocyEOA
+p+ZNkVFyS+URvRtxXbpPuDJ2DAbb7y07m5PIE+BRZOqFhPeQzhSNuEOQUaeVC6zaXXbpXq9Rq5o
IRbzCfaewHz0WntslK23U4spX5YfANWNg04ltLR/qg7wLeyIpPsJM9l3xOgH2PtmfBVrTUF+5boX
egRvyAS28HqM/LENSTJc2EKjHKYP0GIPdD1RyH5Jk70ed5X/hXzgdHBNcQNuLvXJN4oq5cGSDZNa
9WFgt8eccLT5XgHXerasij6Dv/sNFHUaVgbuLXBaS5bhNHqfrmQxzwYulE0wVG199gTonT6JO6TO
CJ7dT6RV0+xoRhWsTKjhpRn+L1Z6D0GCCWNvnF8veR/n6Zy0zeUw1sLvfr9ZVZOAoilXexNvLn+c
4fIQOTposjK9BkCXsLcNYppC0F7aEMTEarZE0O5O+sJMd9M67YOiAZfGGXkWRLP+vr2vbqkRp8uW
9PLqo1+LbVsRsEOOBwkiRAZmLNvyU6coEcD0anSDVbXTpSCiJAfzS2s0cT8MRAPOPBraL+fLRJh5
FOikplffbJaaKRkYQjaVYFIYQfkOqd2VUaGtfGlfHA5QdXHZ2nIB2RMvrtURpzBhJbbKnKJxJHja
SkRPc11UJAdr61dgfF7A0Vr+nmL8OieSTSKvb/i/a5yOn/4CVmUFoisBm6pelGOKDP3NcwA7+Ezg
XoobBA6e7ErIIIQRxgIFPYkDgHLMkbDF4cvRJEB7ii4zqhV51/+fRiPoEuxlDzlgqTtCKc1f/4nM
y/jvJdiDV2L6oar3BLRNuN+ZQXdp1lEJEA97nV1Hx84er2sVlAQuR8chmZafgRNs2hbvOzGGdAXH
qnHWQwJjuqgDoczVxW98Shzt1B/cM5CkSRjWoFO6qWUgMbY38cebLunmqwMxQda3Li3mrqz/AP7j
3Z2uk/tLsVakWiPOqkrm883NBPkMA6CyislShluyRC2GJX/l3qN/qtE1zN4eu7eGuGe1tOa13Gjw
wuwf6fbVVYccNTD+QhhW8QE4pjj3yEjZj/aDqHCaZN4atYvvWhXG3hkk+qTfiuUux7slspLbDASS
JmmF+of8UVzIikIe0gUbZDunZqgIuqh4DKdYPYn1NiKPEX/UbwyEsoK7WzaxeZD9Qu1AL50u2HLV
efJQmgnjngfA9ERGra7Wx3e7fCZOxDK7iZ4asUT9/Q2vkqmcxqvog76yVy8iEWXrHCgIvjPTX2wo
uVYKL5L19xFxGiesE4rysWhuhZ4sfGrFJkRRCYOGAdBF098bZtLQ/gSU9wA49NaMNVqhFHU0Kl9Z
yGFGIRD9EwHtcrNRzZjez7lUcc3oWcvGfR/qLdQ2UwI2FZ1guhM3Za0DHk+ZcKdlckIYnZlRortC
dAV53KFU3fubKeLM8xeP4Y+g9eZLb2TQEUEYvbif/QVr9DZVcJOBg9BgnfbU9MXzPSZsFgR4K8WT
XfZ1S1hp8GkOXd2Xp4QSfml5w71KLqWSvSnUJhxwnwTN7aXGLVXYo+oX4wlo6FHivAmTqBa1Vwx6
qtRmUo9k1cRuziIhDsVqtUaxRT+1eryVnFsuwPFPL/0VZckHdCDw5TqkJLZtftiUCcQHCIZALvVy
CBatPNEbx4mzQmqvEyyup/chVSrFgedutmvExyI0ADCzvOJRMTwN+SQzGSEW6HecOtcushLCHaPY
5xQKq3qZFMdQd0TmGdiO153OyQnsdMCvUV8VXCIh48yGQ4EAngzGd7bGIcEOejsMEiEU9p/m3yL3
mbfgluuRzscttinv0EJsGLhzbJOmM/LXWnfqfr0OWVeqxtwQFNrDYaCmI0n70jfT2B92J+zZasNg
0iPuDv1aVzgHh34dXtBV8+SfjVsWFPmDUjDb3E2IFfIwlhoXqlQnZEnVNhIadaWXx/wF6dFJzY08
lJtjDzWFjce2u17biU47KhHYOMfpHAG/R3e4Gzk4zp4Ot3uWnF94UPtSctSdee9vD7V4NR0I9IvV
Wmhwp6dCBHL2GorGaztJE/eP16lfluFVoyoNBPrADoX9zfpqVVaIjA7K/PO4z6Ciz6iAocXErPka
B4zj9gtHwKIW3NmFOCdmnUzirvWM9NJgCCXNz+LEETbABDJ7j8xZG9scQo2btDTw4iCKDJdtU46q
TgGTOd09RlkZbyIfZfCgZAsuiKRSb4dZtruDIIWGhsydfmLdbBZQkuSVOhwIPiSNM1MZ22Sb3679
cP0/TXn+2iiLYdsQr1TSY98CdJyBcWfuFwcJJwrgChsvu04EptyE1TWcbtvtdaeNM4jiqsd2wJBp
XCxac6jtKSASsg24mEg6us1fB0csD/KaAv94uLrPD4fciltlJEcrWVWi4PrOxQ/mV5oYi5/ZfFhn
y+80wxolZ/KGX1GtAPzGmuKGfUIC4e0dFqIpvDk817k1vkCbvM4wWqxBsIHwlAeIXF6W8CO86/CL
cEWHfi6VkW48y9a6cnsJ/6FsS4y/jLcU2hAoqsx6r0gbjnlzHqRbbUzGpddnn+Golw7tyPe1Ns5y
eK76RdST3oTXNxNE44iD/EguQ3NY+I6m2Gj4xf54DpGqvFsJZX1OqnQSFr3FD1h9WBpLVQBpWZc9
IWG2ruRk430STFEOGM0XLmyNmw7swep71P7ACxnCRusCvUoBkAuRfxrGTnITyOdUAUQRRNAawdYc
sYxIvXSbd1r6RZb0xUYLmjDoVR+udk+eH1ijOiYCGsUSRjzY0xrACYq6Lc9eC6gyKWHtgmdVk48f
Ytdu4ecfilErAyMAJO1Soq+HxibN5W9K+WIlrfVgsesqndl25mTgaIXl71JIwCKp1swt6c+SpGLQ
sXUcZexMoySljUhaO9o8HuN0qPP0XEaoKJv+wunY/hqXKazUq2W0uYNuSb4dELTiwpbzKCanaszo
28Lc7zyESXMRtEg8KBkrKiXXtdfbdKliSrvW+uxnc9A8pU80h2vZObNNVDXGJz8qi3unqvoHLVP2
tUk7VcIYXeigooqF4kHy9a8ntcObkvTMTTXO/2RADBjgbopeIYjBH42u/yMBOJJcRTz0cXsLI2Wu
ssDKrmEPINgW4B3a6y2ZMJlWXBno2ILrJSAwAwyM1zOp+7zPi4fhjwRUd5oWs2TzW4gsstqWHmEo
Bo6H8mqGk+HdeFQtEp/eCLlJwHwJkIu7jmxK+tvMi3F0P8LEmx4VDoVR24OxyF2fCFBrZn6LR4Jl
azSJRGalTgKErIaR+sRQQMf/d08QNCwH7voUXKWAvbyUZ5nGh5XzYTHt0z2y0kbz6C0dV5tWD9GR
rGACCEaHwWOzk5vgESGpaGUCV960zWpIGLdk+QR62c+BSJn+s4OmaUqxWY9oFq4MuDIUWnVi71jd
Nw0gLMVXifvK8UcZ45gHBxSl+GpspITuw4qCEDRrHsR9YvG5BNlIHvDyDD35iH1czLxIUNo0X9YB
qxqOWq1oQtWhK8pIRyT3wM0iZ2R4vO0xOXugSaB6LYDE0Q3COs2KiDq7pr4voowGqQfApnHk3KvI
ApTw0+9xknNSYAJ1i/sP0T2lA6C1um+oVgEiyXfCPj2KsesKskJRVOlvzVs69/zo3RjJW5BgQCxO
W4EI7Krmq0AmXbj57nzhZj4n9en6/JCuAYZJL+t8yqkEvnhNMBcgAkG+mI1Sd1SQl6POs57e1FRI
FqOEdVWE9nviAIsqxTZjswuhhjWkwcPIDAlUBKBYwCLHc4CjYFKFSYr9qjTiQHB3YPxCHJKtd2uG
Y4MOT+ialGxbObJsi8DEvYWZ1mCWBwhW3WMfLLmMB/UbvgbCwE7+LrQsi9fbC61D1KkTlnGhGxEF
H6Hqk3PsgnWMn/co2UL73ZQj5phSUp5rOcVGE4fED5pIhic9RDQJD6sszaOokezcu09+FgQ0HfKz
4jY2FU32Y/1B22aBlC2tFXlka5Is4WPlJyGlCIauQxePvaMTqAL45T7WXZcyoKM2Su185sGKhB4V
AGb3cL2QI6mt9IEvyCqdyqoDq4aZrYX3nDJgHxczZUokvo76G5M7oG1BMoxeYl5IXLvgQuBr8uke
vsHihkDwqMfzasvgm1VDdYZfhNQTHAWUhbfr5lROKdMPIoIKg8OlRv5Q1UicR5avenjOmKclgWV/
V2aCXePowYUCYA8kLvWgeltjvfqq1ymVWLh/A6sSux1mWPp/tt7f4QhYKujpE3ybJK7670+mw6DI
8El64VJqpD2N7Zd7B59N4EHAp7ErC5NKo4XQVlBXzsk9J2YrCyxER7c7MAF6WShmX6Bj6usrXUn4
EQZfuH2bGDa97fPmJrv9/ce5Br/CgNFA19fO1eoLn/zmTMTwkbBjWaZ0UxhwZbiCX36yPYnj5BGX
iS984miwDTN/xSes6gIrfD/SNTaLEMACakQ6NnlulsqeIFz3Mdd4o8yLoVUEGwEG+M3rYxY8ciBe
z3brMiJvZF65TqIGRE2aBifGU5HrrsHTi0rj7mEgPPWg6ZL7CNhwdwhziCph9bUgH07w7566N8G8
oOtsQ74Unwl8wLtO/i6HOQ4iZWQV3nFmvaLzqONPkQCSk7Ysu8HsqonIOj8ARpaTXNM80tCMMLhv
bbsKmAlmz+BtkyDmOJ1zK/DN09Jl1j5B1VRWSc5tpOA6fzME7LCun/TXf+LBYaOyTDe6nFhCg5n9
49WvYdkJJ1bAzH/Tuf4AwMQobKBrcCoJf20+P3HPKTMN92ICN2Y2AwCb5LwuZDNlQvpiWkjlE/Ez
rsKIAmXvGKdZOYQo5uwjHCVjulTGp28q8gsF4fKn8JECuqLVGYEj6QPdQVv5mdTkQUgfPirABK00
CZKo2VFlKhXv11jzN67Qv/lGPzxTo8WeoO0p22tvwjvUF9ecMP+Ggd9AhQRQNCpgX2WowPn1DczM
FvQcWswdyfnFh4YVnkY4P6INoam38nbrivjv5z6EisUOP8aH58sidDNR4lK+REN5KHiQRkDnsfkN
KqvHHw45P7uFDcX2A+EKxF8BPrDJP3uyTBe3xBlOaTzDhcAp4BClwuC15WDWz3mktTdA+09QlkTx
K8MfrWPef0//RVLT8B3oBU+FIxJkJHy4vA5YiIiFRqTYoghOqT4UFqkojzWttydgeD3X9Z7Xehp5
HXG8UqUfr6Z9MEl35aAhMf8nM9j/EJNIw4DgciMkqX6Z9mpYfCN3cMIEl2+3mZf2rn81sa+G6hZk
b/C0v7mahOM6jLBiohp8i/nqxsmFi1EbaMACg2Db5kNepLQtCNHxSEnfq14FXQBUifjZxf+BqIHt
X1oCfCHwL7wtS8D8swwhCWXqTLoiKsRHdljbdwrrXrT5daBDkY1d7DqlbzX3x6D+Wx0NtRjaRCdA
sVVDCj6JHdTwmzXcfaw5xySmFpQyxyEePQMzYH+LiDEu7Lb/wo6ff+BwZBK6nbdQOCltzzeiH/ut
FKWwlAXPNyRfNHtLj6ldsc2JRdPA0+pr3Y2taA1OWEdD8VhptzJ7ANq4ubNCLkMShlmyGgFxHXa4
TP5YMuv0K73fNAqwT4/tM7A5R9jCPBULTb6/zN35L9+qr1jgGed+b+PXF85jNNJWMK8o5eyVHEMu
Y1EQYSqJ6YUlslPZfSgcprd2sXswNxlGNZRwxw2qxqbm5wzXl3HeFogpgfUADlxX6p4mrwiAB/1l
2vSYLenI29chpHGPj7KnwLvVghIPN/9zPHGHXY7r717GX0YFHW0Unqd/PsHxLNNvvCWrP7a9vtb6
o9vyDGm1OlxxemySiwZHfdQh/lMEFk054qRaqniNjHHdIwVSbaIVOicE2l54+k/xhC7l9C1WX7jM
xmPobzaxRZjI5dIuFraO8qW/iXdVgtTbGtjHvilj4dnmjbmLSJnixZB6jefFGLp6voguKHFCcbA3
7LiUc7MjWa3OvwNlUfo4r/RBir6nNjJh5xhXN3AK6dAnD9f+TWuK1BLe+4ROTsKOiP0KRaqBfyhz
+BZciu/JWZo9qc0AtYMo2EH4MQGhcmlzGkwgDmZxytfX8++ETa1qObMCoH5gy3+n9OSY7XqgYJ2M
rPE/X457SWR7ZIGp4ZSGRx5RLjfNlkMVEDOSro3aoMx4wy7fz7ACS6B+rweHNQTqQnkzM0Tto2mF
3wp+EVH2uX9YUjsmiJNFSyWFsajv42xWnn+X7+jix5IDVRuT5exXEJgMvwpyyxVO/IPxIHpoqhWf
k0YSlNtGmM5N9/f3ezDmZroEVCVoqQYvV3tU8lQODIdqE/FJm+4Vg4k/f58yi0U/hDf1DUHe9zE2
3LQJ7Th7nBzG7Q14zZcFHpwdx0u0d0hBiFj94VVylQKku2jusi4j19brhjFdK6+CseJzIBQRH0/H
j1mXvcESiE1DJwwIWPdQoLr1ZW8E2lMub49rZwHHYXfwooqovGTQgbNQ5YcTOwGXKTOY09S52U5K
jlCYxhtLQ49oChz7Y9vVlHrf/o+yB9anv18OOXrM376LXc7hhhsZqwP90XSsvFdW9OiQmDU8TCVx
RWZSpvBbeKMA/KoM0ozR2oJmry4gIL7YNzUtU8AzkzkJam9EN147T8bo0p65FXD1zGHBRL2ikhcm
jtU28IUom/641PW1JKu2L8S+RrX4pYJ41sBBtb08oOEpSLOYu9Sh3L3mILobadSx7de+Ahufnpk7
LHOg+e0aaA1bKBbI6tWHskhs+UwZyPR7eaxIfJF8xz7bDcHLsqjp8QTy8BAi6ZPbOhR+7OFFdyeX
KUvT/sptlxEDQQEYGlMtbQU+9g2vqpuoJlk+yudpFqQyUqagixIVtyZI57Vp4/+2D4frmMzzcSAk
HXiR/ERYzxyWZCUNahTDAo2cHs+E0HPzo4fg47pv37GNgdMWt2iVY+tFezKnWijx97xuKVg+8z7L
VCQ57Z2cgoRDY9B/gLx5yD7IduKeaRSEn6XeN9jy4HHb1Nf195F1yO4jFkzrtMb1czmXA4FMBKJu
JVHpUSgLsnxmPWsI7vzFFaZexuxkHTAcGCkEU8z/w7QAjJnAFhof7/afjhZBMHee1sNgezKbzwqp
H6iF/cBo/bDXEg68xK0cMkD2zo4ogSH2MoDbaCITLkxmpS4lnU9AytfRS5lnWQwDu+ZYQ4tJaIEr
LIuvln3P6ma7sXcc3egv+OLlPfJov9OKmvfqv8nufGdvBn/ChklKKHBeY++KsaPBQ5QylP/nILuK
UitZpQYBv77aDYlBz3WdQRh78ZcD+mc2wbOp5Ce3BWfxDtJOzl5hmbCkALy5OcoQM+iCP1YQyNaR
oJeizDC+FExlCp0UZPjvqmVKNFXP4auCEXqXkEfWU0Xr+ZVNrLk9m2LDvBeRQAb7KwCC2dRynpS5
tesF/Zu0OMO44qP7lPQlJPa691UyLs4l2MfvJq9kw19FwtA9ryIpkf0TmlM9phJxEpONVyHoSWlk
Yl1s91fhLRLF1A835ugrn51AynidozWnJt7Wz3ZXjKSn81FFmTucM2fzz0RQm7vIgrTeTwIRzoUt
yQgfKZ64tfmYEzY+7VewyoZ2ecY+vkuQPfRm9/vCeLDZKmRvmDgYYOToHSJAv0Ntwts4Stl1DFvQ
DxyajdcE551LhuP4JFPzf9ozTjxlSACDQVv6nTV6hIsEj3f6WIAvRzL5FgTYRbNQeijPc5GTqYSk
kTqrhwgPq5YcrWbxfsxzJocHJnWaJ5Frljlef8CNDlRWVkyk6Lo6QZ4Udin1voi8TuCtk7qkv0gP
TjlZ+FHwz8AhkvZRanNVojsBUJxFoKWQOI/mvbUU0x6+mq2t1eEdslqqE9gh4/TpTp44Zn+ik8Hy
f1c3T4EQW4XQ6BMsq0EHkje3Xs69PoKva7dSPiFQuTgGCW4JAeXe3YkvUn4YjvQD9l1cGbLIe54O
4JTIg0/cn2FB5R0eSDTq9ELxJAgq6miRN56kCmxGathXyB2VE2kpvmKiNRuLd18scWvO/2vqe0sO
77unFIwirjKgkqqx/D0My0ZPIaH8eUwWLHSXjT20RahFy7v8PljezRV/lr8LMGH/Ro15AQaab675
VTu9Ifwjg6U2WQyMSoqNKSDv6UXdB/DYsqfPh32eYbHXferk6V1d0bpRzwsB1UDyVhik3pIlCjpB
UkShcqp4rx4jSsp3Hlo0IWwl+hF9VfAhpEXV38yG0igFt7DENyLR+ARBnb36gqcHNNCrs5vDdaYP
Lqk4by5PH0y6KK7ZijGcxxvO80IOsSCXVoIi35Sejq6KYMb2AvXsCPPHr4v3AYVcZVfYr0PzFKMp
T0dH9wymJW4brXNN4eyixQgcd8u18+Tg5Ce/10V5mpsM7FIdrRupb/YjkfPCB8AKd4FLTM71+sUE
SKwGyIJS8hQeddwoZEBRJCdGT9a73OmPmWAsBmcE2OHoJfJO20sNWv2ULJ6Sp93NniLSuDZ0Xocg
m8r3pRjAxm6HYzk5RekGpfWAIZh8aIxuBVFgHALAmZDbaifKSyb5u5HSOtkwft1ns7O1Z+WL9ttO
7H/dvvmLI9Bwqp40E1bPRa5+NOPIWmuVdffa9/JUP27oW34EXfawB1S/K4GgYA/eie9kmQvvyvEy
qiAD1LgKx6PACPLWrK73X9MfiaHaKwEi4EnBBxn4ABRNBR0a2mAi/EE4X0She/uC5Mdr9RlyFNXG
X4lA7HhJlUT9YgJqkGg1beMRQtqYE2ek4edMDGYLTupVntu4enWlS9K8HdI8crm0X8iR0G7UbdGM
Z9DyL8MYrWW8StbcKtYn/1leb2Kdv/Zr4/O3tYbkCj0/mjsohkWvHXDEePgKLZ8bVTjKmZHTCttm
Es9LV60WXoZPQTBSyUr5/ct2U/0zyRq7un1VHWsY3frOB8YNhSNNMbQiYAr5QIPn6lpCZK1mvCN8
gnNrYiLYzFXxuCnC19KU5U161IU4p52PZwcfVdQy7EIDnHVAaOgK8pNI3ESgJO8jYzFTeh2lKuxI
jRSc7p7rI3UBDkbh/o8M5DNre4mwQUzFPHlZfbfKGnIULjJYEjNMo9IkUrNUxL/F+B/HSfzFRrOq
/wyr4bYxjWRNtHt6V73+F6yMtBJHkuXFon9BBT8wxei+ynz2KCytEj8M/M54KgCH2ejvW+Q9fDpF
RA/31g1u0k9WZd6mQkyRhTIWJ010u0iQng2i05O9WEYBmDkHmn0TeHTD30DhOZ24nYIiT26ns0UU
XZpysMLlK285IhUTM0OrPrFvtFvWNgMlLEcdq/oiOOCQdsvpe/cF7vCmORgntdFYYw2dcJ1a/+p8
hsFZzaKbuTJsK87TWji1ZCE9akVznMan2Um1x3K/5hbfSru9T4NnBK0nEyFVkWylkl7mTr5TYWur
Lf+4V19GFWNPXjZoOLwG05K1DDP0lfhX8eHj8E0ITorlt59+xbTj1X16BfmfNG4XpT9K8V9uPTUL
9ZyKd84X5YupGyQHudJy1telgkAE1kn3QOdwAZLMlJiuBHUZBUILTv0uIpROuh6FhKtywm4tRgp7
Dkoji6cIhMGZ2KLXj2XeycV8yxsm8pzcMNjXbtXNV0TBI77vwIrSMh6o1fyWa8i4Wk6577UDn64x
cxgUN3LzX7rkhXcnUv7EkEPx3yHfDMko1NmCV0i5ly2ExHOfjCAL8KqVLNkLFFYK4Tgg1LVHQ067
3dCDvLxOlrqKDkNpEBXAh2iaeZYZtGgC72qliUkzas08mq9qzmVr1qhVYA0XOjFv2Gpk4l+j/Njd
yL7v7vXu/Scyf+M6I00vdeUFeKOd3j1kRS9AEPRo3Cs/11uxvLq6F8vHdqecVCAuFWx5gYKS4yUX
4JC0ViZk87IlMMoyO+1JK4u8O2+s8zaZEvLKzpAijkQS4tyD9SWn546FmbLtik2sO7Ndwl9mP+z1
Np/BGPvzc4tIaGV9Z8I0yWyBLAO5XSdErJfPIKL/RZ0iKtl2H9LJ6yUTC+N+Ui3AqJMYWqqM1bAy
ACpymaezWxAkyv7nJrazKbCkGKWh5UNiakS5aFfbizzK/YCApfTldoEKNZdqS3z1YGkslMvAFI8T
xjJNmrG8QzwOTAMZNCKoUOyEDZN3urHE6zuMifG7vZuJtoHFopjGAmlN4pJj9R1IgoyqQ4fFKMcJ
sh0eOwk5ayxaOSB/7CEbP1YdSa8HyLabUtXPfSDQhs7UHH6pb2RyH3uHLWJGspqL/+utn+FL6FMB
ZwSnXtRlM98sxdoPeqpPoKKVfUy2IrQFWoEIcooKuihF8VceKPgoP2mkiO3rmOzSbolI6rVURZ+q
tHSzB76GW+1K9AHlpD1ojnXi3nyqIqB5VsqLTY2HgWd4ADFK21UPLYpv7PsTUo5uONfhtgYfyywb
6Hv2c4+ldLK0tu9SO5oRpn4zpzjFyJVUwXppmmdCFEoLHOqiEqT6zfxgHEJbhAjn+x4VM+kO6LUs
tZb+QcrWGruHYdXEEzhWamxxc9YPIGW0QB0eE1Sz9Eomrg18u789CbAWk4Yq79DNpVMkzA==
`pragma protect end_protected
