// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:31:36 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
YXPSjvblpJJmr1iSiQXCSN11jHo051RM6YBcoc0A5VWl5eGtJXzj1IWY6z/Ih663
d7fmBrncX/wTTKGQV9vi7vZ2+JxpZI4X8u1/LbtLoeYkmbf6uWg/PlEPwdHNku++
G4zYyPOqJvL99LG2hOcrFUwCI9tRUK47ZOnQxqrRGh4=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 9808)
wnpfYJLj3r+qpJQytfMMQM46STQMmMuTDjv5d8httaV6t9u+dvMEWT8tuXdmQM/A
LhPy3ydzdnTP3tW883VKnlCUFQGGfO3cdL4FccSn59e8Y4eS0DtU5vA2HNnCPQI/
+nmq6R+u16Lyi+HhUpaNV9wHVyKiRyQoSPRESjjqe+cXEsnzDrpk+VHtdJShWE/J
p13SS4lNDPRhhcor9gmKfJa5loiTGTzlDjB2k39B7TgFQiGFXGoymOuomWL2QZc9
+GRYBSflbFxacTQmq6onOdEcRlgiZTUOg2GRWamfjoaZ1EIJz2lGpZTUfkNooYSh
29cvy69DRc7GooY/f2MrTiJberCvWc5ZLbnN2jB86LwVDi99yKdos8J7cWv4vYIS
eKMbH58/Xl8E8gsuj4rZjhTYuW1REByVYZPj8KLshly6QrxjtzwLCiEWQw+4itlm
NJU5OuKdbd2offx5WRCB7H0O661b7gXsVGtLuWifrwNSOjR3i818g5W/5nEUdbrh
mBFXyzPKw/SlmRHMPGCyBKRysecNiZTanIwTcUR8YpWt8uS6qtRo0N+JA8h4BcgU
HBApz1MNWluC89Y8KzyWI4WNoKtvoKxg5lG9TccUoL/6q/cAz1Edrh+Tta+Fd6gb
vQZYK8zyoE7M0fhavwD9kOM+TRnl0+AdGf6CmMgL2jmo3S7elgVBGblkK/68VNW/
BeQe3cqminuAQiv2GBseI+ramR2/YcTEgeYCzNOQuSPC3lxjnZuAYedK3Nt2i30v
R/Rio/eZhw4A+FFAF4u0+uwJyIypN5CnzC6Kh4PeQjhA3/1flaZYsF7C29bKOklD
KDYl09Lhb5jZ91ObQnUjapamVbBn3ZEGrbxQGv9nMZe2Yz1Ve/gdWEArP6sO7wdT
pXwl1dJdkJzyGmxuWmgxpqiUgmdrd6YponOpvRb4UVw/Ujd+jR6+NS3nBkGzX4Kk
g2rvzmFentFd9XBtPuj4s/NL7pKTdMC6VkaVA6m3g4adB7Cdrc12H3ng2MMAp3wu
0Lvp7Zk8I7yoBXAXTxB60O76W4xwAnkEDmSnJq+ulgwGRBGzG1MGfHNXoB/i8TmR
DXFdCUTa6CY3w8l38KqRlTPleCa4AgLhZ1lPBUjX5TW3Y4dHJm+B6xNjK9QS2+Q6
/Yo/9STZehN4h7b7xR4KNPapirsfiyEn6Y3prDHOqMtlxpBc1iUZGMnED1Ijp4tt
gxVvYzAyiRljUAvCow4I3lrVNTmRMGegZUYTgHM8PLDirf2b72LQaUkSICyx95ac
ueEwtsffTaQJE1mXFVr36SGYpe4opKgTTDYZMIvwTYEKk84ehZSu5qftb9cyUibU
RN94xnynuHEdiCCTPv7Y0dZ3B2+EKKpHqoKkCFIRLZlOe0D/Z1/FtkAf3uT1J8OI
D+8ybUqXayl7LqG0V163Plbl6sq6acMAylzpJ+7JZHtMsVjuA9tb0wiZaSN/TGpy
GVYDhJWx/l25/CBrDHEdkBcmM9R34kjDlo/6CF5SFuVV67CtjarcmTJ5IpTnPrYf
JZO2A2sVQzRlByF4c12Funjbxn74GcIm2sn0al9gQMAwdeGwNXWNd3vuYg3+s1eQ
Bsg2vYp5o2gtb4NMOCpmLenkDBASW2KsJykvz3Y4vayyJOnzIPLSWeqwrKIopK/I
MjFOjrxknwt13hZ8h9CGWdTHMmJtBl4Rrkd8WLCZ6kqQcGsH9grtm70W1fAX8TEW
CV3XaySNo2OfYAQIds11lXg2xMASnQWdl+N9gKZZH/MhL9wBZMfHlPgNlI83ppAQ
uk3Fhb7IX/cz/UC1xj/q2ha4ldVT6RNAm8N9j5d1RdjOszos62clvPquUxpKVn5R
3dp2GWAmSFmFhuqiV4KIRb6uyfYmLCA8PpppxSs9o7unsD8BSPtWxTba+boS3wsS
Mmad5tALVktItIUhVqW9XO1mo45e0mfOtlgRAehPnIbzDUMiuVurXccCoHywKTFs
J6kj3yZHm2+3ydMrDqDp15NRSpGd8cKcso/KoZ3Ea9lSq3yWscNrIwuxvbLmUIsD
EA//iptK4F1f/9j62BTuOu3QfcnuX4Yr/zmPSP3cnMJd80vihIOfGmQ0piKYsT3O
Ppza61HXWUUD9KsnmXWJhgYdUx1YSF76kk7x2U2iKoXzisgSQuUxdpLSE3trtdTJ
E5K+LH5xouzDMdlZ/sT4YSAIJARgq7f1QNjnQ0vP44vLxSN4aq4c4yk029uGZOI3
tn0cgUwYduJKQRd7DYRYBjsJI4X00hL9wI4qTXAKQLTRefxDxwhsTwpptyw5mEPU
feQiO1aYqK9H4OrtEzeV6uH6sOdsmxP9nJ21ft26nlsFlD08zPQfwm9m7C+1lYIA
JqXJ1h54KB9EL9gWqGUNDBojNcGAvmMun9xcMr7Sll65WPvwKKIj5IN9DFeHYv4V
+LvszCnLLDpyXVfEHNloDOBx21X6t6HcDhXk6OHBHmnwiuCPaNpSGpHb/zLKB7hK
5S7q/VpGGxIPodFGIXUbKnrINv/g4H30iEYq6tw/TQJ16vjFEnsd1KIaF2Pi6KY4
H+0AwIT6bEJCFozBNkkc3hcdMZMl3kDJMKkdx1JGoPHLdnNqOCY16VC5XElV3qQ5
Zxlt4aE3gHV/TQzIgMuiAwK0Z+9L0CctdMy9DL1XH3rMokBNHXEAfVkikP1TtD3C
GDKiHeMdSfxFlwcMZb6hSTQ6hWUbilgfrShK30W2Kd2vFNu5x1CFWT2JIscFLjZU
s13Pb3dU7OMfCjD6sbIBIjJoazqgugfGyBk8EJfejCfWSb4OIaPqgZDZ4d+mX53L
JMZsLn8jMrIL4kE8baDufiM4PWax0g4K0CGbv2+3qFavNC+5oD6YLHrJmX57fTd0
vi7mNOAEwph1WWEz40D93mn5dUi9mGOY/M/vn1A4vkmXv2w8rUj5EWW2bpQeWuyA
ckSLq7G11oRny6QTcneGvKnX2vZyhhJ0vawk/NEfwPZ9ZyshwB+orwJa762uWzQ2
eNipYOCztSdbuzxoZSar7PjAgE+yXEBCw/I6N15jG9GfjZ36aRCB3POfe2VRgMI1
ClFuhTIZwaLS/FOlzTTgc2R1LyaQrLGYIM/p6mKw1S0kyXATxbXal9yQQJvmm6HN
ijZ7MvQKITMZ++NrEmg6t9H8amzUylNGjRS7or1GRAuK630VrvV+6OTfUE6lzqJz
BDHrITRgKnT+eJfHlobI9AKraGRYLQPL+eFa0kLzPpUz1JfBQ2O7/67YeZxHcadh
f2rcmjEF42lvZmscu5fV2TM6jheoIuHsGzu1UmngWsop6GDKcw4tlx0TU9hJxYfx
fIl4U7q1VXJqLEzCrKScwqWPTxvIig1CXMFb9yvMdKgu6WaWQEnOjzOmPc1h2RpJ
ZspwfjKk/Lv3Q40xVBB3G1Q6CXMnKIaMoIG0UHAV2ut0bVN7xnpcc8gxNUUqVPrN
nKX7cGNkGVGoOGrNROxGu2sjyJcSf3+pshUA1tOmcmDtPaoI8MV25/yECQJjqvzU
6e5QVHmUkjhQ3acvk25dxjZ4NoJqst4EBIoNtWqS0iBjSECy2cTPAcDVUeAYQgHR
lxZcgz+Knjn7Xsa/vLy4VPA8+af3V6GiR9qnEWOpCl63Fuw/NcB1YCHI5Nn92nH2
LVSwWc5GIBqsnB2vyBVU1+jZXVgIiYvw9aWKlxsrqvsnie1HI6o8XQKFaOScB1tZ
k5aNLzfrkhQXxs0H+wtQQN9+e3yz+ymaSYzfx+ReMxLpgFj5PlWqc4TYHLqOcIB4
Aw6EIX9JPfAudDuc0yqcigx8GX0oLQkyI31Ty8Fi1Q+6uFG3fJaoxGTfqaF1Ujta
OnI2ydYPuDYbpX9hU52mpr0MOw4qHrq0TNfY1KYO+O/qjT/Y/kXcZvGzJaOa/OBQ
3iKGf8QmFKR2lJtfnL/DzX+1+i0QUygCZBzO1Ta0DekAa2OlAmgfE9psS9b9+zt6
lJqSoFjth+gKl1wHRvrYcmc01z27G9OmwfZk88eE/kerv4PkIE9uUUqG8wTx/deQ
FVbrzHGIj4tEaijAbmpUFOYpPuUoEvZ4jukaBNS1bzWoGko3DtGy+VU6mby4ibNe
GJ8ggWMoK5eIJ05zLcV9uJj2wMzTdKopWB3/AS7eqggYaVfG/jOxYCnM7XD/Ep5B
oSytJ24ccamecojv8+hczAdbYeG+fQ/qLlddU50HIn4nmk52oxeNE9ewIbln0AXO
41/G3dDsAeTt9vXroO3H2w5BimUrsQo/XxyQmYfXBASRmRmm5K5lJgxVDp/vTilO
zSDmlo5z+tvTWveOTX0h8/zPdUjqlQInCWxYnwqiZSaZJIzCNtznB6GugFsWz4NE
GBMPrPZdk5jF17KtAkVKXnj0IWuq3AME+B+gNvqZ0ggbfam6R7ah7BvZ7xlurnry
2Q0i1YJEfq6W0nmnZkZKlGj0ZTA/K5SCaajAPwpk/+AD0lbNwVcFspCJLPTW4BZf
mA+IoLatItDAx3jPaXb+KDgleviMEVFwTpPMSaJ1J4l03WpxfksZ4dXrxT7ClWo6
1Y+eLdkcmynw08ot9rgMZTx5SNdBKS08i8dDLqatPIxYsKGZaC2FqlH9WBJKlhrq
a8T6dFG888RNaa0Zefsk7Xihr0l/SJ/ApBgpo6WU87fKSQeFhkceqLVZmd4uSxWr
v9x9p8By8PN/EoLeLYwp85/MFXodcxdttyssBGBf42Ryhyc4hALXACF6MC1SP8UC
19B2BsDn4bosAbSU3NT2eGsaBE8RLoLYAIXwOaG8EhvcBBjz8pV4jfu4/XnUmiKX
axTfU4HArGqXzhiEGySG/yYe0lI6evl0ZkvzSZOCKrTnptV0gFJQLOHpIixbnbpJ
bWNzIgzF+p77NYstibNrHA7ZZ+MTDjSCbt//YAOyuXDxxqXxKt03B1gNUIhzisk+
czmfmActDis9s5MpDjASBzA+sfMdHp4I3RTNk96txmpYkvJx139bpZ5b7/iD7U4m
BvUVnoGomvbyTUedyK4b4uOpzZuJZazwJhUppXZSJibCQH3aa+mCmLnLfQjMhwSY
DFgX40IAKseiEzxmZ+obslCWjXY8bOENBBC+P5U9VLh0cPqygLiS+CXPa6g1Qe7/
uSLoUbdrYACbqZDiGreT7wqRs2YXWvkaV175ZLsrDLASuCL54Yj3JAf7BUE5OS5q
pBgiBX2i4Bf1QGj+oGC1Xit6/7NGwe0UvIp5TpObLUMs+K4K70RUsc43G6VwgI83
B2UBBkER+KMrKIKVVRp3lLqsORFWnxy2s6pcIwodIlscHbuZkkrZpo7PeVPCLedM
FvC6IPD4CXqF52LFYeydK6xHKZxBmyVEoAixsln/S8ZsWZk4qvO/WPo7c+MOM/TL
oPU136g9HlMaTKArnii92sVnAqeVBBK39gamTNjXSXrrpJLzv24AIp1XAGiJumvf
jO1PKkiudxlluDPj68SFTCr0RfPZ1edEJg1i0EAqfKJjvD5mj8zpARnrCwuBLdrp
fprCO2H1BM/FtLIGPpYQH1nnUkSCWfxpBC+ppPYIb+HMlPshfKp5zd6HFQtTeaDf
qH9BZ/FsAbZSNgrjFNS8KIsak/3vBWSbmVDO/jb/juyOqwN3rKf4viOX514NMGuM
bckT96KqVPJuISnDIik1LnS4K5IfAhilTq0HRx0frtawaURQ3mrPRElGcEzsbXmt
dwJ51NTG9JtgRLRyDZ7GJa2SOpvrO4Do66ZZXtCRtEgrUU18D/80kdQHODGr7N8F
N/siIUe2mJONfzoUwdMQPQ0geP5f10zQ8Q7T+ynDlpsJcSd5fvn/DXRdyMAWWZED
WTE+k4VF9vmZI/wOkTATOKXdyYtFbpOnS+aHCzoxbI8hjTrHcYPBEi3purfLvZBq
hYzXtyBZvzvRyYVupm4I/fwf6v7opgYWFR/8t19djVz5F/mc2LmzxAXlQz72qh3I
IQhnU+CdXUNpWQKHvoSGtTqtDGUFgwvCKP09Re7jjdduUsZyPIPzWpJ38V3gPZ7B
sqReOi8H0/BHA/++gRarYqYKpM5WIIzgSi8GrCLxwK9HYBaiQJX8ofwMwgBxQXKQ
nOrfk6zKgtFs+P7xlrfokSyGxg2QzEEjq69PjQs7FcRjasLWRRfF+zKo5SQw+zMt
zlp6X7k4/usM5lzTGFSLkDZzqudcM51bnA/gS/9N/z/H8EVAlBYZB83ERNRbDpZ0
wL+DyA68SKP3DyMxu0Hwgg1Ozk/8YJuPaG4ApIvzWcZiqRg/1M3bvDP0ofbqqL5S
RbH1CUZR2Qfj6j7oet8sSxhNtoSCF7PO40zBUgKqO0cDRLVQ4bqYd9cH6reIH7gR
4l3p4NbI+KH3gRlL7LoKgEImx53oK1xcp3c7fGZGGgZDAVNhJKPK3IMlny61UPb9
EaaT0DN+893CQNBoOowOYrPyr/DecoB6/p5rCDc2MzAIi/McfiEaNegJSN+kEL1/
0WBLB6dB67yGmvje+5YzcOMBcoQXyGiLBjOGEk80NonrnpTSVcleL/4tKTOM/op7
Fh0DXz7iH4p73noIPhbC6mebNK9pQhEOpjFXvUS8RG9Kaay5fHcdzDGVjiYBaEre
j51KF8QKlkHBXrswWnKIrsqvSEmmlr19Fi2R2mlwD7fW6maPCaYHW6RJmKOqqMhc
OG2HVaxefjLYXU4w5ADakIQKQ+fVo40Cn8Ysq+e/1NeLsPWuAjjIIGbdrjmECj0n
NbNXZV59dyXjNbnjD2dayyUGa/EHMZBTrdiTj5oKbQgLqc8fWtmkhfhcOUgRkWMV
CYfG8zO9tWptmeQH+JzRJj3UJKJkeszuyjuMufeZHx+ATYpHMNGj6vkW+SiDymfo
RhZ4cL5r0pw2MaHBYPwGGfqWrst/PRug+sdIgOJoY47l7YMy2gK8Wzg6YmBJGW6U
fO+567kZj9pfQaiRucZ0RI3q29ogtfaAE/40NmwhCXVFpKNsXMEQuoPoK7Mg94LG
v7RA5dm4BQaKtVFEiKVOYxOFY9FRg+NQBoe6burXeNgnW+fJ+GgA6wehpgL63KwT
5QdiakS2Vv2GsDT58jrb7k/5UF4gkMzXyYo6jNn3zzQ+jaMhrdcqf8eBBGqRypr3
4rn7fuEjXYwz9HrhS0zp5stOR9lwt6DLR5FSfXAnodHO9gtX+z4kaTLXE94yHTdt
MsVCgtb+okR2raAP0bjtpEw7SGa4c8Yi9cD7e9fPkXGyHrJd4vVEhD490hsC/6xu
paz8AOtOOIV30Ewv8c36HsnoVf0X3CmDkrGdATv8QcVlgga7q0vVZGSuV4eM4B+r
Msmi2JNQHT8rLxcElRM03L71/fceldvJN5CwuV0pZue9YlnPt4knTOlU9hFzHPqc
00uNRa47F9xkbEJNJQQb5IqHk8PvAJM3CapSiSJK9ng/cZbpappNjheaANrzOw+d
8K+CPmTypzdudcTcwso2lMLMg+xWa+BPDVz9Q/CfdLe9r85WArXbhKRYZkOv8k0k
rcvzzMdzEF3+08ng+nsxG/XKWRQIUW/rqlUX8ZsJ1/dim8YKLkOhDY0nHgiKfLn6
9g+tyq1HqnM3Dhh/iZ7GgM4T2pk7js6e6F3RXPbLiYqR5fKmBf0kiiLYWL6gTqYN
csyaq2XmayHGiXW1N8Eof0CcMZdm3Hrm66TJNC8rjIDnMZHk2crlUKBG2z/kmhNw
2UG1eKYuqozFto8ehZeS6yEGa2Ins6YioI4HZdrGT2RRTXy5XCrhgAMvwRv6ptkw
RvSaBleXJsev99gxvSaiT8Yg/y6Em6Y8HLU5G1IdDdo391mbztoYPpNWf72mG5y4
X0xYWcAGLjE3zdXOjLBf7uwapdK924E1II07+LhWwDz55RN4QpYEtooCTzw4c6dJ
avsM6Dg6IjfdBaypUR0cviHGniUENWVSGgpdmsU1uaN7ZJ5L4Py5Ro3qlVe0v2xf
XBROgv7/+tjNTeEc82gmDNNRMWtjkab5qIpozsOf8lyQCLvJwGlvOe1K33GzhEoU
jM+R0qq7fknLkrtI10HlrIrb5C7uBfixkiBqpIzimTybHYgOvYbdprlllKpgLvTL
d9kjmzP6S4ikLIU7N4k/SwcgmOsR8MerU1rxYS4obassZWjYRc/9+Qenmx5zF8+1
Qb5lER8o33FcHw/mnzyEHaf2OjD1nxbwC0urZ5ptacJnPx6v8pjc3LOOqlngaCRH
Myk4bBxzZkWAKPg+6f11HTu2FNBtcoY7XB/5tVWBTLdm3sX7wFzKEpZzw6eq+mSs
6W+Afd/wo+LhBKwKtB4FimwHpuuhWj746jqVI8AEnw7neOwvHZMniQHnAYBju7Bf
BUHD3OTe0k6/v+jxmZVe4vPtwIcC/gB0do6llp4ZXxMOrwGZdvdV9i2BY+czrXsk
E/5TToIG3cId1v32epausg3jeiTqyaCfOuWH9jH9CVx88Nai6Q9Pe1DJj/TcblJl
iHylrunT8cfdMmaZJa0K+idD6dvF+NXGtN6yNdCJI/QrSt5mgldokct6e+onzFip
gOGdSpuYCe7bfS+EbbkMvyD8MRjGhjDVWFxQO/SHNwGoLJVp2fAKBzLu/tKglIJG
LkWWERYFSbpQoszSZKMUIEGOYanEgGiF8LBfs7CHkDPpkW8zM6njqVvhhdoMS57k
xCC8L+9Mw7PGYlF5essluN5y5HbkjvlDOmb8nUHyX3N/nCXk2eg9Et/aRXyhrWPf
hSGtAWD4361dMk68+jW3PVUc2FICHaYcGcC7Jr+uKfflboqWQZQvDULLAvVFkOw7
MiKrMAGJi6iFl/EHHrnJcf+mpRnQcFD321SPKlRcEJWxaLaTRXrWvxcFToWfvxEO
w4eqr7ygJ+WFxr0qKbWfrhmOvHJ0drDTMe/kCCUTX64IgWinFAAI9yRzYXc02P+l
NPHqosc5SzS4SVZwbnsib+/dmi+T/L2EL4zaS0AlVHs63+ooNAgPNiIhhTz0WnYD
uzd7yEhDmMKU9e0vjuOsleMGRXv1Ftp7ata9Bf/vDh55EHImnuOrXhADJDKKVeQ2
ziLtDHfVMmpojGlW5UM5X5sZ/JfcULr1IUs90UlewkIETLe8UyDxTcPYXVmEygzd
7IMKOIybDqPvvXz0yy4odwxdzm9XIQfBccKnDkjOwL28U5b/sMX/aNRf8bqG3U6I
7JovdtFdhAOoLPEh+vOeGoKRgHfHaI7p6ZaZAfn53wxq3VF2qgEZ4qpWXLr5DYeG
mXJv1aAr0kyCSv6QREyAI4gVovDf4iRqGMDbPPdPqVFM7yLfYFl8fo6SQkolGfOS
ZMqM2rjtC86RDzag/HpvQCAZpl5VLzJZWWWRDxqN1bxjamyJYVIVupoMHkkJz8j2
XI0x7MiVdIQh79NC9FTSPG7JHQDRnU0yru5XuSPsjTlj8EPeiFDkl61yh9TEYVgy
8gi3Vg+nDKBnTLjn4FnPJ+YpvYKwF74j3TsdDcTKI2nbK3CoV/mcB27buVfr2faD
2L1Mx9mbqB8zANUc+y+rcxMbaoOhVi2nU/K7EI2b42OKs0cjqb6Dcj0nol7oe/8V
RYI2pqMK5LYSbmAAOk4WUbiFuyyroQUvPfqj7MaJTTYme+LIOS9gW3PKoqxEEQrU
A95T2zBipKbRByxgw7jan3rY7bSoP9cpW2wrr+734uGyEb1nnlK5DcS0Uji9dr6z
LKirJ4g401k+6D1RqnlftrT6mIqFWhtaNJQu3IH5q9BVwCY6vGlbGHvJ5z8BX8Ag
rWzDoFljnAhT4QWfmR7rZczmvuPeG2DIEn77oPUmXHAwXK00jZdDMB9aJagQJI8z
vbc1VV1wm1UpZXIeijfAsnQ6ePqPU+B5c8bWm80jOSRVmhE25K735jDAfzIkssJJ
biqn2z81nSbCw92LrC5LmMuugN8cJXtMlQ0vHOTQHmExQfNyP/sa281pzTmuFzq/
RQ+AiRkWXP/OD+ev2/wPqzDQZP6w+xMUIjqmgX8Xv1iafl2we9Huc0Pz1QYxVNY9
Mtz0vOGDoE6prpZJDyNr7TwEl3fWCI6i4yoKLmhdVQNcE4KRp7G4db/NmjwCcfSN
9oGjsbmPXD1u0irufcQ+0ImR3sGPSD2NXs1RgEE3x+735TDcoPS0ftAl/6Mihpwj
kJ3CSfTCYZ0HxII3f15FYYK4ooBCwuCv4UJa/SVEUqipugdFFNdk0tA6hZac0rla
GkQnGtDUqyAdKKY+EFkYas+Lpfkoflv0aXk/CGJYH9WvCYEtZwBf5nMq+LgRaYJ/
w3OMEA0EZ+GrNxTFoIkTUJ62mQcsuYk3UkUOV9+7A/T+4gW87EZTfFBcAyZlGPIX
/lSnEqgTThOygV+x3GpmG5dgLrvOy7S58cVpDhU2nN6fDt0loZYgRw7PqDheLKpM
5NPIcqUU+4+qF3YTlTDeGR/VkndGK9dQbMlvxITw3m4GBfE8M/odxjcUm+I5wNY/
Ckc0XQ8XKkwiw+sqJeOxgje8mGbmIDtNbqctYZzPcccrVAq9yywwHRcjfZoJnBtV
60Q2Xzanb8oXF2Pd4Pjikg6VCsDS7RxDEwbkhYFZYsbcVMnuUjX60HHFZMzTXPx1
jOQbewMpgKIDHDWYmZVs1K1ta7Ixwmi3nsZY51AHi13vCL1Xsii2+9/jt5sYNfvQ
ggxDgOdqD2d26z5wCoRcZE5lqfLr1LezVv6GRfYK+mS82KBrUJAonXbHM/WkYrU0
OBlWjDYQXhHIBneMpcbD6PInVY0b5mlBdcs7SjFs+gkUDjHSud3iZ4tNBI5xg4C0
bvvo1xBHouSRNr+zcDMdSUGsQ9FLcXOE1f5EqG4cDMmOAvcXX5MN/JOaY3RWXgvi
1eUtR32awhdlunK2qoBNGMsWdsYkcKrOGnhRq/CS32BrdO8vACmE1jhiVQz4SOph
P31WD/HhKmwERJPMXpk1j8wgt/WKC6Mp79/ETg5rgV063z9fFyuuwANz6pRU0pOd
vYtvw4UxTrkCI219GkWibQUKynXF5Lczp2LDdm6/8G7cYnNC4F21r6s8ioj1oncW
vuI0YFepHdFZsTmvHYrPNYigqkG3nY19ABd9FTgt42XkJ/LcWonlhuwDU3VgKJPb
KyzQDNvU2UJNj63eXMMO/iqHBakWI4Pd9YExib+YznWFbopBQOiYbiM3Mj9zI9w0
WPGZnkOw8ALkyYpTpaqDH3Rt/0rPvtusmW8uV3lIYk33R3ANSlX4jURMqgh8CFsH
PzhC6fLAW3YzRVN53d9ina3XslWM5iZ8Ts84r6HMmwxCPDvydFaQWtq8yDLUxoZa
K3oE4wlwAYw2KBDnp6p0KVu4DWvTltviGf7JqICwHxYZlYMPVyeERf26ncF1p7I/
wo0tW3p83w1xG2LS2L4v5mXOxyXfRNPkEFQLhxobYCsopnk1ifrtrJ/m2XzKKUZt
tESim1mXlmWPuvp94eMi2EpOVhH4tKH1hYMTnZsg+LqTw2BSezLYbEh/5reCEuoh
WCrgltdDgLiOyQtLq3WfU5dezIacA+7R197BsmJRmByTn9lLRXGhbVNExUrBLrh3
MwPxVIynyZY7eaTRc2L0cyzAadcr2MNCkuwSm4Q2e9rz4Z0T8PfQyIPTtkt09K7q
NUgnqFPTD7IoT9xh3O+Oh+Me4xsjw5eGzG34uQKomnXpV9RyT+flKBFOdIKIYPqk
+tULC+BDxWbqCVoKdpwgxE7WPn13idO51jEhl+2aNLTUsFFGgeXOuSsLpWsm7hiS
zU+Mcuc7rweC4cf4YADrt8fYlP7qHfeJ2pqOhgGehf1of4mxvE5RTEG62fRZZ5k4
IlCIvuV1bM5ZqCHd/PzEijtV+qzLiJQ59/bhWU80SC1o4JEk7Vhw7I+OPM8mn71w
t5MBfSBYwttE2ge618riuPF0yzHYAoikO9L2eHRGx5Og5EsfTarHdcppa4WqPIaf
bFevvGRoaJKhQa0KRfZ5Y99oFfb4HZRi/GEboVva5ZUucAMviL83vXIDiskvIOE8
kU93s75WlydBkjnUeyu8sIJEd2xXH8pv7i9wybcv3mC7RpOnJdHk8XYCLkND91v/
wOaxPKN9jDZyFao1qoihjCxokOA6rOEWAzebNtZrKPTVVZzly/LnSKi0bqhmf1HA
vJZYcX/sRwhYA0559HjiyvDjDOOVEdc5FUX68CYdVR5N7/XUoPdTUSeMSuDy4tjq
N58At0RAtHIe7MviyEvF177lOKIS/ufrp2wCKkrW0w24L/I0Ehj49EHHMdVHgGZB
fUnvDdo1+U97uNfYwOuoIYKQW5QUbdmPB6oMLGUbl02bHqAZPmGxLZnc4KhzxFdL
+GI7fPNlSx7lqjmrnGNPAMu4vkv6KwNqOek7hzV5EWEtjxU4HSE2spuFbPCcs00I
+/DjtDxC7RtE1S8U0A3i1UAzH53AodwGiU6HqdT4F8e/wbJQBPhqAOYPFmovy4fc
BtjvwBkDJsPgCXcle9/6a4shypOqD10/I4b+5BahS9maGbY3W13p0WaTAIC+bsu4
mb2lamLUOiuMBEcWBLTIoJ/5jEkhfDKG0WJ21xrFlQG5X4KIRgbkSFbbs3Hh8KT8
FE/OXEdqJ+xFxioY9kyb9bjGWrzJ3Ok4/lFdTtv4HJ41LjO6+1dWhKEy+hkcuYJr
26dVbC3bDUg9gNgd+UmMFXkSKltT/SsNdCXpj/C0ap+M3Rh9E2IRRoU57mcIM7D2
wef3IhgUJ4QGS2GmE7Zff8j4Od6YtrR+yUV3fGBUfm5HiWOzAHkteGaH8PsfoABy
Fkr0aT/rhUb4MXQCEyxN3FWgCkNlv/cWfbgWT7Oy4lbtxoHal7E+vBkhJIg17fpi
kXbblLjZhUevj3lmRnkStSfrlqjdFhBdTp3u8ZZ5HNECrSks5i9AThaEIvh9rmlc
y8wvmRQjgApyGN6bkSp+xgJo7GwU0wCfPH2aYdEPjXetkRyLcNsyRh7rgtRsPPk7
o04PG5/kjSNkzxwZSje3184rJMb2Z5WJa7deXIRvGIyjbNBvXiTyPFSam5yeMg1H
PtPmmtYB5IYq1iFayUkPF09UpGP+539YdkSH7/su4uWDRsKzVYiWD1jHuP618aum
YbzJ91D5QQppm/UZQrtfAA==
`pragma protect end_protected
