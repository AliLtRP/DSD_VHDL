// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:40 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
SzwvluYPOSuNPg8cqn4ViPH7fAwKXz9rMDaJjjMf84cqYpiZNnCWn/ykfkcQZR0j
dInsDw93yjprQ1rXW/wrKD2DvaHBXzTDkFhDzYIkRHh3kR4kAYeAZuMk7P2zu5zi
Kw6ZhJY4xy9c1ZrT2yCNdsAm2K228HrDKJgp4477mwc=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 14560)
VRdLzzDW7bfVcQANVSaGDtkOq3vLY1uBt+57kympaBojMqrZeMlJCsnyYNKjLpHf
0HaxW6arR9ORHJLqnn/XhWBwuCkY/k1alv01i1P6upVb7WhWZrUUCphuje6Vay8A
ucdHrdqlCkmYYEDtdvL/l6/d12J8X73vyzCpMkl/t5KGmxGFONPSV3GX2Uzd5jFm
ObwOHn1rj9joxxmxrjOnkR9yqkLCyMaigTp3f0NKVS7saku533WEVaCZegk+voWa
NJcl8LB1s0SjrYC+xUMnTR/z6g2abK7KZgJxjzuWGIMGQ17OgAv8j3oaGmFACXhA
f9so4HDRaeHkS3wrb0iVp08+ytk4j997lb0mfk4sjeswQ8qayvwxrbmogDgZ8jkC
LHOaI76Kit0dS2tOVhf1ysJoVKcR3qiGflFNcfxz1wT1pbOHwtMRXwVptjlGNesF
PYtsVj+NkM/RdeeZJmMAeguj/PpS6L0HbDQHk+eHoscHL2ERfqy7a/cK53gK4ujc
a6iwDz2ePjoGk8SUB/HR+NEhgLm8dBZBkcp2MuRSDZJzro+U3sLHWIrRR6KE9u4C
77yOxifLQi0ZeETb8kGScXR91PnUM/LsWUgx/sm3HddLmKeSPnA0o8Jt4Ul0Dngr
dA6i+HC3q9NM6TnXQ8Gww8AWXUmaDwcq3CBN6w091s422SX9e/no3U/AQ/GWr4wX
9Zoh6GHYOqJSJbkxlxQFGBnksTA+zXPSiObuuhMfjulJF2e20pJ7FX41p/xcT/Gf
cPo+ZGrtwY41bow+CIVlnc5FZ2aLo+3aJft8PBNKuObfQyUzyzb64C6FRjHfKilX
ztwQ+8m9sIAZtbjcZdmOdetVhjvatNMZA2w2BC+M/noyeamnjI2ugHlchBzsUGe8
JDQs9IbRmuLblnIexCL3trJIAGjPcQC6OFOfwIGSd2ujpK/CVPHNujK2sAF412H+
ceVtfUANVnp1CeL4zLuIVeeMdapu6K3WLHZmuUtomVyjVE8bmtHwSN69n41BlfD5
iOfBLPElIZ6Op3eXMGdsNlrznBiLFEJ50eY8JtWTFIgv3G5EZ6PNDsnYtDT1kexG
f+L+9IZsQDLKzwbjRfqi1poWDJoCVxslUCjiuV3BN652rW0Z2IPt+S9/Ojjmxosm
2UKyu4sHSHxgcnIsrlL5gX2hq8xKQavZETujHNmlmway/OBCdcrOSTtm7glRIa3m
Hj3feGkSEXXvkl97uJ78t7P3vc2b88obNpSQmUOQXNO663rJx7R5ZFhn85yohH3a
zGbxLidtGcqOBsGn6NTTjyydmoNH3m2HsNvkj6wHLjfIhx6XR3w4nJq4mNsyFwIm
oSIRiRwo30025rH912QwlLaJvQ0UfKWKuv9vMuH2i00r2zyhJhZULe1sv2cHV1Yu
z5cubI5WygACLdPeKs/473x2Jgvk5qMFMS5kT1r1Aruye6Qhcsj1GtilIiu8Vvdy
U3Rc7lZQLUtQ6b2O+69GyUrQXcovGurWX4BaXxsGKsYmXMxElfwMrQdirfvphbQ9
VJ4968O6tSeOyRDycXFratv37KBZ3pIzqsCCAr6jWGvRu/BgNLoxzZnohovn5Jp1
mzAfvr+k78zozgrQvmc3pNM4XCfkK2PKjIb4D8TfvYK9UF7FwG+AoZ7fBhk4oB2K
9Bl6vP/S5EdfQ3hkkqYPgTdatkroUjNMTS6MtsSJUXM8My8tvaU8cMUeM+Bn2ObI
aEZ9VHhj58xxhsvlOjiaMV71Ks1eLFPdCl1f4rsfgZW2lkGSu0mQlGoaELZuhZS+
QH/rJlG+glcvRS/l2T0r6RbmRb9mZhtL0iov7dvCkNOoK5Q6NcTJ09ynGHQoc2/w
Uu2hbcPlK0qn4x9qP6vB59A9lZlcizXy7MzULyZpe6Aa7aHxIuJu0KXGyW2IzZMh
GhXvd3fb2ACBSe/PY+SztWd1RyF4ZhqeQj5xeIzYziMJI3PeigczqkYopOhuIVDo
3Dad+iNBTp3RbcFZI8HcWQYfjSGaLou/occNVtKd+IxyNWc1s22ic+Zp89N+FDOD
eoMITCQEQy0mhKYAByRXga3q85eCg4meY2RtkOowpBdrXKwxrKcyR2cWREk6+I1g
G/5/YdCAJSTMxn2ygkCk6ZufITfW4F39EABVQ/lbz7yd+jSn4PJy3SnPnBBS9Td5
PVbIczdemX3glNLT/Njl1gq0WwIYhvcJLW7pcKUpg8wHcr+N4InUIEMYKW2Tku05
d+WkupSTZxVHKrhykQCrIzfYRHK9GeEGtwHyxZN08NhqsaeZhTV1fRqXRV0EgpOX
AX5vGU2AISxFSiYq1U0OXmV2TxHA70JS1xUbY0mz8D1Bh4Oi5/zdzLSIzMvz5vhh
+fBT4+kngJsxDlvV6/PM7zXrXOpw885oWOqgiDkcx/un0ZpUg7rar90OpGG7P1K2
jt1tzkf2AINNkLo7dIydub4ju1mJBX8GmKJucCrTYKqKkfNmVUwGIHFt9PX83DXo
l/Zmw9gP0jTcFgeuqsQm6nT/4mWhaKZhnEqs1lNrFl+3bMggMaFGMTfe5g/oWlyE
HNR0Qwx/V8gi6svam0BwjroUehKyBipI0yBYjDeFlfnkAYaOFiVzgb/uViZcJh+h
5OhiUtoLck0g6PySt4+4w4wZqcezu6xDwvTnfdtfGRkhrJbYr1xManN50gtQGF+M
57MrRL1UQtW96Pttppp1G0ZihoM9951TI7Q0Vhzsfm7Usa8xB0L/KdVQ27KIXzQz
j89QEQjRVUbKahAEgCkBFrMhlxwRVJBSguHH1QuS7AWqDVV9uL1oyh/L2KyCzoFH
nseKR9OM0eV+0GlGZ23GYM3FF4e3bgMgmaJ/rCIVNO9Zv6ua/esO9ChH9CPi5lD9
cUITPnLy0FW6CR0iT7LAFRnnUq8gjbH/380ylPSwsp+6QCUt9+vFD+SmJifzWkKJ
fVQb5bOKTkCX2VNTfrjnwJpoCYhllH0g0ldm4I1BQxNY2un07U695rzvWkjJqg2W
EhYy3oYWdcPr9ppb75wfM9FlA3fQhTzZpsjIbrNWqnZEkAu/+JyJiWEavy9BCDdM
UBGGbU3Vm5o5mjfFBu9z3t0b59De5PGob4vrgSgF68lirxvJ/2KZMKAId1o0olaT
IXBhjTJNuaeJmzvP9l7QvX2tY1NEC1TgnL1H7BxswIfVqsZ1tHZaldx9JXnO5VK2
pTwpFVKHawi6ODZh8YC5KSJjiFX1KBXENsXAtMCu92IGYc9vYlEWtOWgAV2kTmFs
i8tiKpvPO1p5NCZibhM+riNoycybjcrrzIFhGEqWZyXFyLV+LRM5vq2QW7StPO4Q
SJeUxTIoysxAsx/byIICRFsyhiKKWwW/Wj/2xd84si2oGpw/SceEQl2EuGwxAAxJ
nRZ5fNTjWp9i2UrFYMUHDOYl/qGJPgdphPMEk4UzRxIH2x1VPH0WVo/x27b39x7c
/0IYpSKadMdMfwGQi3/D2KmhL5wxVLJb47JMlsDKLhzZE0LayQHbioaz1S94/PGD
ZCU8Pc/xmk7KUAUPF4sTx0gPGhRrn0rX0sGtkm3zJzaC2UlhiwD3h3/M/CS5o5no
XpzudctV1qucxTY0vJ4k7ZyXFU65iOF0+j0LNXavlKz8erLSbnlqBRXTraUq9LZO
5J5CuhAGDw7NKtja7OdIInVrLdI0kWg85XMyikUtLL3fk0Sei7RSkbRoTVt/FoAp
fP39dHVIoDgE2TWZxwHZHi2PeouSMmBeFgg5z4qjCBG86tpa42mwhqjoW4+ZiTo6
cIDWn6npf3McZpNXml4orpokiVKAynWA8CdUrzzdJ96I9cK88fav1dOW6O3f/5V4
mMUF03waTSRKq4057Z770bC70EcWZhddWei50JiaW+mRSZJxluX7SGZE5Fdqp+61
7xFWa0H3OQqLJ2PPGF5kXoei/0vQwP/rZjsLWzhFcfyNU/16E9zT4ZD8YMA3R9AO
U/g5+tqB+jEYx6NUjEcbckKXfKBAkeHT0KuOg8dIi4xq6OVqG8xRTH5hBoaZCab5
1xlVkt9YGz0uhzMGB/hHVsAtVv24EG3zZbtBelJ7uBmbK1wyM95RdSdwKBnxKJa8
9dc/Nm8FH9xIlORUwS2N5fLfbYIePkZxDUw/fAl3Wg9TglRmNfF0SZkBFioeOCfK
0JtSNzakuJpLDh7w59mLWIchHDmJ3a8lkTUB5R0KPMsHhrMAbOCzbGYTC0op7IO+
VFdJRsk5PJJu1p/spuY7Y9lKIClL8qfPd/aQ3ja32xNKC5GqR69iMSyPFubeheEy
5AYEhD35wvS4FYxKnb+F+4JjMzziK+Oxx3nETYti4YtHpJsBEcNL5DqT5OSPJTjK
snfmOQwH8FE9QrZkaVfR+iK57CvYsbSZgqYuaT3RLDeAVHB1H9ejjoyb+kMzCa1S
X3sEUmTEWPLwmHDC61IVBxY9FKU7iDi/yyQvwO7d4xIAFc9HYSuR2a2Klbrb5o5J
arXUSL5DAtv/Ap+ncXzMBktgmwmANmuMPel428YgQkQatZ8YGMp+viq3eQfdxa/v
KRJuySAx10eml8U52ylzPUZ/X6R/gb3HVJugU8MiQzmX4qabixgpuQwgrLkR1Co/
QTn3oTVp+NujNHqIYU72gW2qFiMhfDTAF/eWGeLbyxx3MF1hOuu+fw3DmQBbC92U
2mvnpo7pnRb65nXmAv71Z/lXKVv7KFVJQxGfXKdnPmn0ZSL7s+zLbJsAc1K66488
p9CotaUoyF4VCk6BcwAf+IxFXnQR27KUZuF/JbRc6kQW+M5+WExB8h7YDONrepIG
hPz9QI/HzkMNbzwMjm5B+vZ/iMgB96+f87+YidsAqkvFmng4UZh/ddItJRm9z1I6
YujAP4QCuGSE6mkX31Q1+k/1FX+y2E20cm9kUnLK74oYv/VKmbcYutRR5cyIYXaI
ATFAHd6DkJQrtFwlyBHmFBt0A23XW+TFZMH+xUpV8SBTqtz8WLmyRfLGtWR8Tl+i
EcOTsSXvJ/RBZZktXb4ysE7CNuskf6bqXPZLNoZXp1IjKKDWYCgLGPjchF7QXSwF
FXRqBBXnTUViMkt42Rvwv5eOh0DuTa+LU8S9451dvHf3sg2ixZa0QTyhJw61RHuS
V7FrEdvoRSgXfv/7KFjfrsfi/8ffBd1Rdu3idwCBy+u8cMXkTzh9qHbITSWepe01
Xn8jftE2C936u1ZXmzexPc5qWAJOY2ld8fL6ie6s6XvQaqDGdAJmyAKS7PSK1yLs
xXW1TpZOgnQo5neiQd+dPFeYZrt74pezj8y7NzN9p1FbdxrE0UDmbF7IJZCCfawh
6N5yH+CZNZ7dbd2MuMIp1DZT+wuMbfOVbgVrPrWkfRggj4twkd4pzbhTeAtCLI9m
wmxsoXDhIYSOstgcf3RXqjwQ08ukqYzt0EsqA51hoG2YZWr5wpaaKOIKPgBtum1i
WOli/u2WSfldwoMm2xdJSrLr/1sUwzQaP76PEUyFceQmrUzWZbbpdUJtRri4i04g
I5B+4DRUdeWltMb/Fb5u+OgbnF+63VVp8jmYhzmr55Bjy9fnjOiknGfanwnePyP3
ojVrIyhayaYpAkHKGw59txDGAQQ0AXV3dfB7sQ4HzGqhSQyUBVEKyXEPW50JJrt1
EZ6PWaAzz1rH6i3f7qEDBH5zTBWJioCYZPyQ8OJk/myHLm5S0CkOfecrbOg8ubV7
nLJFshnFwQJx3cT0be9bAImZblPpKsOuHB1w1/n1FqwW8c9YaTq2akot9sgCmDes
gn5QOqR/BSZLJ7Gjf8u5wagz2GWX8G/wMlSTY8zMenX9ZZPoKowaHVLcpFeehmk7
HFnbOVmBD+ewEs/VwGfMhHHROXLc0pdtnN8kKEN090kO2rZ5AI5kG1szALwZtGDw
CtVUEN5rBAqXOTUFtonoOppQTc86ftu8kqgDC5Wq+d1UcM0pU7T9ghxOjTjbTnIM
QoxePVYveyXudSb2NTRO/dL+PP9L5LLALg2WYKbpO61ac0czSyiRTUTF9EkS3Vch
tKbwSkWzlIHaQwXYuh/76sdAehvYkZj7Un5XEinVqS/7iH0YDlOp1kChH5qJMTsu
aJwMdtz8yqiUaRSbwJQLgSsz6Eqotj+I+WhQ6LVDog9eqjim6/69rKjXaY4yd2Fx
Dh6Kxcxmm/hSJSWuPfcK6TQ8g6jvX556Hgq1ZWmxvuvMXpaa66P1Hp90ji3s2cBo
QIp0M110RYdY7/Ic68YFUS6ztpGwyM/UJYyZj32OIQIzFb8i6jXxhivRI6Y1SL73
w/t/JCCK1wHqWQ44s/N0536Bkn1qXHjqzMMQYqbsbGy4sEcLQ5MnZgXZTSY/1k8K
u3o5VuC6Vfd8wTMhvegDYq5VHCTyXIhjU/AQEEm7vaMo463h+0WPyxaY5eLpW0Uy
Fd6i1ouVCu89eSPzexf1RIjI93w3A/XVQ8Eil3vipnPhlYUrwR7DJwBKiiUi13Ff
BuDkwEHqCftEzcfTinTccqoCA43T3UMDGlokoQueHXYUaOJSXJ4dV2M4ANDBdFSU
uhwWCtHabktWubjinIQLs6ca4KJObXqLM3pcetTCWWkbcrbM+iSwKDE5q+ylNcmR
1Jt0sn9ScFlYcR65EgR2TbFW92AiP8fioaYwwqB3xGGL88Yh9vdYVZ2k86bygZuU
vfy7ADLmvgMFQTeu58iD0afwWCAXMtXDya+8bjLPVG0PKiCygabhRDzDhyYbC+dF
jK19IRKXsOKx+5iLGoULe6RpSeLIrJqKyAOz2NA1uDp3amVPULMDFmSR+ZZtr0dn
gdBKc1TAq6rDi/886nd2L3nsdHTh7tYGNmh9RdH+ME5jatdjFS1MbHukt7R23NBI
YQt/o98AF14bbetRgwLPWdvOf/gSPNgoTGt5TnFtTSjvcuQ+XllwUnf3hdRmqMOh
10La1g1s1E9QIb/p87ecf+L3aup2VFGBkbMPdJ9q73tDfqVuzRn7N86CRMWTGUB1
Ph1HdTpImp6y9Es5gYlXLqz8DDhaViVqItJVvp5t+xaiebmdw0xhRxggsU5Jy/1m
O7JN1K0xfgp2mB+LfWOtnm0o9sj2mxkii3Liv3OZwBvTMzb7mJnRa5Iog/wI0Tzp
9/I/lFiB0naZPgsVuTg4o1oKPPBVP1efbkuG7U9mOAHbKGFSLo0+FGuBdcl1zH7D
fDET6yGywsGQ8QimxVmpQ1LvzwGYXaD3VjLmoChiGFd/w5Cn2ywN0GSA4W0wd9Lx
6UjCGq5KcoPEXlavfh5Jjj5qm1SzqcTQ9083zUsC0AlzQnRn2CW/J15IC0mhO9uL
HErzDKLoxasRnqk4eTHxFn3GiLjiEC+JtrUVdJSElfXGSnLUfIrRWykniS2F2Xk4
Bq6IsF9LizAcidg3c0noFtMJIMecEiu8fKp/v+e4ZOQN/OAL1F/923bxbLG1C7lK
q6so5GyyBTN2ox9W+y25YH0EzZtS1oKHEtOf0iYLI7Tn3WkV0HBR6BRiXVWsRJ9n
AbyYogGe+I7IV5qzTnrqrvedI4ulqV3IFBUItndV2HOyrr9uNW/p0cY5o37Vfele
ocCYuKe1dR20HvoN3XY6erhkujhpr216XeMg2YmWKNlPaGqb74bPpSnwp7Qeb0V2
/pSrbEfsOh8eka8Z42a0Iq7GssHHtkFcr2GhjFq5QFNRQx9N224HFqWVvg+sJ816
1OrWWdifDrYqsBiHx3Wx3cK9CV1dJpwlssM6ZvycR7WQg64gjdGEeqAprkHPMdtW
stB09QxPh+R1EnNV8dyBYsOgXJw3gupVEwypbmHhV3ulqajPDqg2WuHozj0fRJ8U
htjORRotBe8J/twLCGE/2PuGdV7Ehr8cO6b9dbHr2vIOpZAY3eKtZvTNYCqCgsrf
kMtCGEozVn6Gv2QjmSWCZtsNWl9XnvVyx54tBqOcuVX9pWeAP/a8CBYLwzKvGwbB
M/JKfRFSaSG5l3u4QpLg2qBaVvuu/cLpUewpdmJt+Vco4HtKRKztMr4mKHcbS3sH
Pc/tNx2T2f6OqjIcQFKzx4o2zmzo4py5KgL9Uxct/FzDPl0Wk3axJwv23ELIIptS
Fc2g6Hm7oyOAPpOcOKNcQWZ2MFBwLMZVdyZXpmF4FvW6IzhgL/MiRvxkdhKtVYnn
MZRU/ewIgw7lEdBZbmX1KbsLHpnaQwNFm3qJnkjPGUOr1/g/yJBnIumOWwDJWvWW
6zoH4VjAT8ZF5F6P4w+tPMthmJxs7L/87qn0BQEMf09NiZcL+4A1JKOMSuGpCGwg
VrzcO26WfvFcA3QUB1Ryexp6x2mkNkv0eIpT3g7I7YcrYopuurH6vYcMVdQznq/A
tl9Uw9rklE2zLHPh0rzcodZexsRODOzF94GTHdDJbcNZgyQlgIIqRKJ6f4gaxqfK
EWRsbe22MYacgbCJxgArABaHGQ0vYQXBIfUYqfxrloDTNJjvGCs5qEzkROecwtBN
FioOSYZ2cl5M7VPyonqwPcMgPOXk/O7PnXEAJ+t8JWDiPm1pckZuj/Yao4zKCfua
ilZYKgDrAQQq1NZqIqACh3yQX2fGqWCA8ppg1ywGgMsIZd9UmTB5smlHFnQ7gcg8
5n39TgBJDUrpR00QuUHSDoGc6JGWq7pTPR3Z3yUkxMQ87tZgFln4MYC/5ZWJCFcW
J9ISPxiED7EuZCZ6V+YshY2oIlCW2W0Nu294/Z5hhPyzbqDG1u/GozaTxN2vzBJl
UeKrRaEiozbDnDrAIuVPJBU/EJAbbJt0YCQxPETTk6Lsw4dCtWk+qM+EtbhaI521
87yG+p3c9+1AS28aljwjC2b1JOfUdEYohyykrA3j1qbx9vWUsVRgd/iWRcQDQc0Z
LTcXgR7ak6vs+0zpghfERiKw4WGiElJk2cIKCjpG/vVdsEnh5mA0lBGZtoqPQpK7
i7ZHAhVQHDtNBwibJTkXg+N87gdxyPjVrmwk7L0MDddBPaSUJ+nctyYsw9Puhqjx
t4HxOX0e83qOAl7z9HX6B3o8l1teLwW5BYZ7BaHEFAGCFpOD1/jNaLHotGX9bIKA
gRwwyQobaojmyR4aAw/sGZzwOQFIOmpwcInXub6RLxYYTcwyhGk8fiYsOIAMq2YO
jOYh4YjqZ4FPoBlrjPMIrITqEuZ/2yuKe1g3VtwDBHW3u2Dgm8XfimocLkZa4Q1A
/8ti+MEiNoIciDpjtiPEIHZzHiiL4Mwp0RMWcI5IDzn3qQL9H22G5auNxNUVXtLs
g6NkOKkqJi4PT9Uw+1/BqUZY02hvAaZu9PqmVJ44hHK6SHhdohil2PF6HR15PcqI
RJXhfNCSketZPBfX1dWwdyUiWvcCWZHNZrEz2efjm1kb/PHzW5wZSHeVuRzW2AMA
eLq41OKEcBg0BgmWw6pth9bpqfT/golmhTP9807qDrfepCJTlyg++QiLPjeKVeIm
t6mA1Zf9LseZHvc4aJMJeaXEbj08GBy5hF2RVaB3YH07Zio3JignJK0xo3SaUrmW
rC9TxZFetYEBMjfCY5ua7qqYdrPKGLyCAbeFaaJdYz1FYwIpXDUUPN0sDpPNoXnz
fd8VdoznxkjRegU4udBFOJVab2+kjr253mf7gDGJtdOjuKNm1c80oWh1+u79mdiJ
zOpECSFOIj9thD4kzAk/DVwWAv0pweXABWOLh6STRn9gWCyv12X5go8nGuelZViu
RFpvjpMi4zxAmmF/XA+FbKQ8YVq4OO94qc3yHIHFK8fYk2ODXkHS6bcCIZniGr19
JUt/1WiY8nU4fmO4Uhxz6nYm88DW+iMPz9oXnDadjCRJmbgEKARYbWcuzZCz/Qf4
BTGVuJn/6SWQdpdR4ObycUrXwU9dOIqJxeItbMrx/DchoXi3FI0j8FdE++W+bK/m
3CtZGkVvEGdtirWo0QRh52jWxwoYr0Coyd38QGmHeyAzrkStZ5bqhm39WvbQNGW+
JdAbeeGa59dItbo40ceaCGZu1TYHTVSYiFDM1lAZDkoW+jA3Y21P5W11ZdgUrnOo
PLvztjLkxYOedUlcZBWLpVyZpu6m6hD8zNGJJCTNH7xdFJgLcrYugnsa9BiZ5jcv
7Ujg/P85uXO3O3BmgTRN8MLBPgVHBbXKofDrOIOzFlr94IxqRJ4pgCXEsL3UGogk
Zrk+XqRrBw3Z0ZOtPMbwjQ2ZotJEHo/Hxw8Y1zmCa2Z2/K5IFehr7WlmJZuOV9pW
ZzTZ+42olb1O0ysLhKIxArtHm8INQnkB50OaG4lXN5McmTtX/PPMEzwbQ//vsikp
JURKzjrL4hHwA7RDDFXlVbA8n8cPcWd0gulHfMeg3R3k+N4T7ZsqBPV3S13E43Xt
+Y+4szHQQn07tqxRRA6NcL48GvgzgAe0ZXaM3twM7qa0veWHIUTadX5G2FKrS52Q
X72dl+yvvt4TsfnSvMQedyAel9zlMrEuRnfxKm26FMoqXMD7pxStPtcRvFZCNd9l
NWGtO1vvxVV1NjK5UOiO7NXtGXxutw731pTCMFfAA2O72UEdCce02WUKlWmkFcDi
3ADCl+8gW6siBUf6T0zP+KyZq1ICRFTS7utvjqU9lj+kTwIDpPEbXR0e5n+DLUZ4
Kole3DVTGyP/uwVD0SCN5oGwWt534WZczVOmZMmSfM7Z0HaKPi/w0NLla6h7Xlyw
AcTKXtq2ahyEAqmAKcbRL6Zjmsbfj7lHct/ptAXmom98vnUqvQe3Dt7WWdRDS+nz
/9ehnHR7PS6NXIx3okdUIdZXYN1bLCYgF0SD5SNumS4ZwESM5Nd3doQuc5BT7fBe
aS7FK7JD4Nc39y0BtiM+kGhbt3caMMrgn9WyLdahQ2LE0+j+/dUdMFpTU6YHsLop
u4FhiIdpQNniC3Kf8lGqK8TEedoOvCvt+cyuDN43yO2FhV+BhlNAQx8I4hjOAkb8
lzWgtUCFKahNFfIfaLA8iiqugVp8ivTPPDez6zobUzVN4NnAuf5VVBMCudsmq531
BOMXy1DioQGkRhXdacUk0zxOA8PvPWFgSHoy9ECwvu9vdMw8VDEiZAgYqds1pUCf
xuoeCaA3npsaEMhPhqxyM/T+Ip0cVAn+822T/KNMFQgOtDvNc6YyfvEqa62IceAd
FUZL2xTBWWW3YAJjwRcfblC5l+PrLvB6BQIh9Tc7vSPEunOyQltcscPudfyq1va6
KUfioy1tC5v9F12DOX5NUE1KyPN/QuaNbBajzG2SCH992cdz1HyjK9Zi8tlmXfIu
DhL2K3vkREv71p62ErViVB3z5lHpUwPTT7K/r6gUWCC390/iPbha11VnmeyfzUh/
ehQ1Pql4eGke2hoQ/HYMa5rkwGIoRDacs5Nkhkb8H/G3W4bIq7kDstD0U3nIhnyU
Ip94ocHUEOnCMBJqXGAPwEZWZt6l+SDV/JzGRV2YM2BvzgKuViR0BNOYPfCMjN32
W0jpiNlgow64SxRwpbAsks4eYcUNJ/rtfDPJJ9JB8mZiaURCXNEwt+UYTS2EuVkB
PGfnMMvs5xW4sTUbi4zkCcsr8nF4qoRvx4VgIenhVRTjbxNVaEHNsoJMEEuThc4c
It2wGF6ZUsUrhIRCyjpSY2UoriWcHREeCtiu4+l4MbaWTYe9/5GlF6zDo24oSUPa
hDa9kzmfRTY281tXcxJtK/Jd93q1TIMhYQ7BcCYHg1ZWwr00LSvMFUJtOW73tdU2
9fYZtJMhD7DlfhxQXJsYXU5zG7Y/5NZeBB9xHf45UY6/Bp8/j883yGRYlvn/b1az
v65BRQocSUCSfOXitXByYoIH/Ze6x/6+wTUEXQucMbv6LhNG0npsF0oxJqzrHVtN
AZUFEn9MTYB5fACgiZp9vceEe3SzcneCciTTQ/hO96fK1R9xL0qOl+Dahu1lSHBp
0/TO8UHKD1kc9zWAqacsLw8hgb73ICakvJTS7ZQ/tY5fWgbT+iPQrlM104GT1WuS
KYh2DBzc9tAF8OFxXemCkh4o0ujaA1Rssi5qoq9B16lIWh1X5ZJncb5UcXWDTaqW
/oOOiAu1UNRFsQWmm2Z/pb7WXY5cB9Ll9nEHRsgO8LyJssSgW6QOKxoXXfOaRSsd
6U4u3lVSu/tZXDCvPNOVwLGGfbLFYlgWzrvqeAs4ieDzjb6driVb2/iPrf0pcL80
WMwBypmVkScraYl7ult/ZwvTVGFqWII/fxk7Bt2xwy18eeYTsnzsrVsIEQFK8qDx
L9eeQo54BV9+u1n2Vl0VL6eEHnCZFIZ/kDYeObaFitUrgxByiuHSkrnZ+ZP2rk15
quvgys63oK43eIH9UzZzbSpVwNiNC3e1PgMJBjNXUykvWQdD6aKVWMeAB3Ziq2ze
ETN8QYNyJedEby7OowjlW02YeDiZPiqOrZwo9TNTgQ9L7URXuhbAI0CTl17DGaP9
L3rp07J9IKcyELj4n9vkkNRAcESXZ9UbqHoyh06+D2sdNRL11nL7A/CVyJbyzmU1
rCWtxWt64cRF0AViDMBe+THh7as5GiEtDZipW4Gy7TlrLPsSYZlGt+b0rox7Xg2m
6TgtFhmpLli+vwKyGHtJvxlnvFYIpXEZBIfvJdgQwTvqPBztOpiBOgblTaW+/PyR
QgXPp4FdTxZ8i/AiEdZrO/xkV+gUPuifV/eL+yGDfy5euUHPyMEXO0tE1uyy1FPn
HPYNAhGsmU8sJyQuGGBF4Uht6trk1bwFoBO8qRHBkKurh8rDwMPpbemjcR36iLKm
nfCx7vvdsXBsEgU4Fs7kTdY/dC25S5KRJQn39kNFHfqBqeYfPupRUxVArp272uZb
USEoNCo+5OuHLXeQsunlVtTB+qd+1BUD08FIDmA1xciNBXcD6dN8PiEmqT+MePhL
c20C71xygmQPJWtOIEmEsKoP/o7JJeqqKsX9t855Xk/oB8gOvqfI/SBov2KqyU8l
nOU8nmnbD5UikAVPOl66xjyOQUy+wbcL4Pa8tIV/203+oM0t5u9edz+7TcOlsQID
JV74SsXgTEY/Io8BKA5aJqhOygor2adhjjMK9xVb350fA9e/XY75F0d5mwU8szIP
2hxi/fUCFsfkHcWiBN9rEgOtP1WpvJh4Jyo64zcVqJX25t3IInWSqLkkZy3g8a1X
vSvSJr7KfbpYlM4lXZ+Un/zSuOEzn+QnR5AzLY7VxvNMtOCgpDNIF8S65WfKtiga
TkG2lqV+D60AJyDeg1z1VyMFKwj4TY19ge3bvbh1CBPZ+/4dmntQa6O7Zb4shjpK
nA4ENj3uHiC+GqUui1oDJn5wMEVhbawAfJHfolT04vytEPOxqD5ct1idPEtbwpvz
JFfRgkt770ZmxKmVx/emKwo5NtDuDQUilhbwFsTCA1SJ0nqvLSGZzJri440/fJbE
7047Z0WL6EuKLsnJFnv07cwgkCet9SrHBQeUL8SaWyszkkmwmOaoEiZq5K6gl9Yc
YNF5aJDvIToBBC2rHx2m4kyym4NODkxq4p5ROkOhX/VX7jBvgSjMSIEns+XnV+Oo
TEKdh5On4+LuS29ymulW/zff2judI46brfcE+GpVvX5Oms81YZ1xvnDgOrroSqO4
po/sd9M8acxGxGX7SPN/bGY3Uv7WysDc0RNKUnlAkwXDMFIEmsLeDZWFMoDgTyi/
/Wh4F2AxRdudaPUOEY32WRRbbgP6SSZONf5wGZ5nFaA5nfvozbZil1ZE9z12Ab8T
Gbrlr/e6dYOVmE+SbujM+KEjIdos36LEZi4pGCdePcHmqCzYQoBY09Y6ibhuBtBu
ufZI7UH4F3o5w0L49SfebqJQedzjpJhSR8eoxXPHb98PuHnxqNVRCbnqEaMj158X
/tuSPOEtaxA1tJtrSZwh9BE3G2+yex8TpHy4KRdlTstmy3p+tmABzUSbyhQ9Mmw5
SsX5JNXm1sybqytsOdSFNjuEiFtiwbWFSonOknXTfjvZfpCAU45V0HJW46/T0eB+
qggiriecxO4LxqEiYO0rJLwQWgzlPWPH9L73A2Uc1EB7DvMo/cWfijkiPntEx25j
pvS9rqdW3aqp+qjLcujVb+gOEedKcQhoFsC0+L69qlkNCrK2Q3CDMPiDMWdMHtXP
2/9V41Ltwram4KNAUTl5yi7McBmfHTcqvlo25xidI084PsrH+qVwJNNo4MnzHaQH
RNQEQ/zbEtjjxB3LGEOtD74EfZ1fW64WTi22qAcrulHLKhwPGMJ/C6cdvE73sHBO
EnmCADIzkSiXVZSa2tNiXDy+f0s5Yzzv18YFCTBGDlPfKFiaiEyWsh/Ly3/fH4zN
6C1/nvFdOsOsZXPU8Bt0+rE7JzKz60/Z3AQpy4LKDEFehRNGmoq5pRRTan9QmshZ
m2soTwa5i+yYB9UWkvV82t/PO6b+hjr64KIFefeqvhOC9zdOBoCA4ZOVHVIXIekX
moD2nd65Br87nRIbVj2GxblPpO8A6ErCP4EGIOpuo7s3TkvoCHzuVlqL+r0PLrI6
b1zYUjY5OIEMHRTRwZOVAx5jxMqpoVGF/d6NIMQ5zsQ2wtnWhZryUjtap4QCi+iV
gjraSaabuaJOfpxbpdzdWDTxseqPRCAIexACrwCX6mPZ8fhtnye5fzEa+f6IKq5Z
BmqDXeYqT+IVkM4eeJIiB3YMik+GJ/9XGKzesYHb2ZZEdoRTxWT+HH0+tSyTUrAE
2r92AM5S7OwU4N6AXFjXvaSCQ1qaqUopmhroXpI9H0UfmMQxlipzz0HkRG7+l/j/
Iv1LIeT25VRvpGVVxTdAf/AhFcCkTKwSk2u9BW8Se1viuYY6QNoORQgkAaCJ2H1n
2Yb7lyEDN9TVbXJM/D8aYnRoJeqplbDl6AgEVTvPQQNx1lBNlgH9enT1OSdQAPNl
YTXeQeWSw9enaduQ35w2zshaJglzfA2QLc/WhtXSfa/H3uMJz7i9qbttb7MzDajp
uOQSqxQL+5kxc7J0rA+dypJbZmUOSSQNuVhoChpZmNI9dWt1jphpmfkaibF9+xcB
82+bLVT5N8j7g+v4rirslt289b/1cHI+pGjcHx4zmOQp3VVOTCdxFwtAzu4orN7N
JoLHRzO0pxinszSbldhomcQAeFrrc2umOlRkPmegznO1JCYBHLGtBIEdm1m4vWm3
HSvfRk1VwKQdhKbxxx69amTdXx8ii6tKVTr6RwKJ4Du/OD2u7KlOfZD/a3tHLvM1
iPlQcxjjJqSMYC8cF8y9GQIWGcxwsihX13rpwmSjaEduyDAGOohnenzOfiMmtjLG
OlSx+kx+/LYWiB2OUwnxJn6nkIzSwlvqUe1PqegjJ9/ctTIDFGnVWkx/veT93Xu6
KvYzWzkpmH/+B97wIblGqD1lSYWj1DpiTEI2FTBYUaWWSgcC+ZcM+gg84XIjJ01Y
z2gRoz2nKfOUIEOlbY8F9df9cVTJCoeSH19j6eBU4H8s5EtDrGmPpAJkBykBnM/X
Exm4PDObL0wYPnrzcWuBVMJ6o/gcA2pQB/HYBIUMQxm026VvDr7brP5zi0xriWzv
3WWTC7gjB4hWp0PMzNl1J84+/4MUfioZAaOFnvmlVrPW4dqBtbOyM6lGNaQ9V2Dl
4yZDiJcA5H/1A8eT2+Ierpg4LfrGXAIZ0yNyFQWZr/n3yaz7JAFz77wlTbQtu6bq
505g+/6jcRkPJHt7w/yUJqKAGRB6idnnTG4S7CHMPjCGKRBq0VJimI37QlVaagD0
+dTlWodWnJ6/9d8GUvXpN3rwQ58FOOd8IjnCeXTAOPxJpan9zOhNNOpzSiGidq1o
4OKPtAchb56X7kVCf/B4qMLnmtFtp5p+NYGaC+CcLJcZ4/BH40SzGT3rP4ejlbXT
tc1PNBgXJGPtFKhQh6zXaAHyW+c5RPGbyZrMi+2A/QnEOEsdG5L+31rPG8gr/ZQm
h/4S0ygIRA1bY27qWqbOl9fmiPme5stb/XJpnEhnloIthGKKdZsM7RSUnwVXAvyh
JGKlrzTbGx4mNrJ7p8TqBPRBFEcVYK9HtQF2n4OlgZqxGdyT4izryHjuyybG3MZk
jLh5quH0EF30f/rl5q7HZVZhLdBfX/JiVpCpMChDTRk5ZPf1Ua1Zy8FmHFa3C1vY
Gd9NLxh6NkBI9SsvNYm0HEAeppWvarjaGD7KBXCuashv9mlXXRoJv8OtSjG7ai7I
Wgw7KOl2bmSLOHIVsdlb44Psgrt16j3R7NaeKF15ETbQA+uzqpOs+QA9JpKKnG/1
unVpVZtSAUMLgmJ8s4f8HORFcFkdNa3ReTMdfYtILRfp4gXIF7emjzzX1Y2J+FeR
qOHYQH2UnTMa65xeYSMHPL+bgAL3w7ddXi7JnPfwpwtd9opW0NY/FcQEsJmtb9Qk
n0rvmB9tkOrptGzBwnNih2o4FnaD+9VHPRKI3PE3VKRW4jhvhU+rRc8j4Dty21on
G8XGjM8r/q0Kb/EYuDHhZc0VjeiBSP5wJYC+NKwGK+8GWPPg48c+nRP59Cb36L+U
LPTixD+D20IrmxMLog/OQWA2zqBH4QF+5FMwn7eTrjfURvO2VUiFKvI9pBvly/iU
N9FNtVAzNAzRzE2Qy/NpgQQXZMQyghK6mOIy5GiG3ukT/geLpBK20OPzT3lHWg/i
nYT+bluIT8ASDotLpK1ySIEgLPEKVH5t6OyBmWxCuCg57xkVAR1aqscfE8Qr34u9
4waNW5J05h8epjw/7Mb0Cm6kWKv+NDwrSVF0XGKhnglaidHX14hZ9wIRc1jHEKu0
PgEv4XQmjYMfTqBOzq5pCTiYEuJ0KjmGxwPw1Zrmh474wEq4EGgS7aKPU6HiQPHX
FNIrd1CrPg6icBOPL1X+5t7HLwy9Np8B1sfv0QbvTz4wrzZN4HIOjbPrxe629E3O
uWl1EOab5LjjWH7SG7wNgfOBY2DBHhIPwxKj6pgwDrlTNU6KsFEfpcW86d+UYJu9
7nt0GehE3meaUaV/9EUf888EwzYdcMn7KUmCnTpA/l4O9P5cGhJaBuP19tU8pEF2
zt5aKSwdmL0U0r6hQimo8ezjfnnFC+eA2rfXDaDS4jyZRuG29bqEL6BXKJebd4g1
ThSrXIpxYd8U/6syxoS+TgZCkTDDl4Fp36NZuTHyOy3iIciH/hTg4xu0rP5KjfO+
edvbRSRYJxFkys53IfMCH++SHCFSnhUVXEisxPI8PhEVfhcBjLM30sAQLLbRgZ5I
KtxzDseEM+1oix8STQ5IRix/AwAflASrOL9gZBK09wlNDKV/2Rksqys2xKI9KR6H
8nIkkJuRmJxuQtVNwdD0GTMx5byeIIIqRlIl1Ga5glgD/R0PVi7WZMURSrkY1z4P
8VCRBDe6JbdW1eLt+ZsXUbckHQjV4A6NUuoX3dcXYk8ILSwCH4pd2feXpofnJSkl
zvxgFUipCWvqLU3FQAENoeOpMvJ07+22d7Kb6gAijGJeUgU6l+0e6LAlkmxiFXFk
lY3B1RF3nsM2OQ8SA5fsjxDaxiNmp3+Len2KbGX2uhoWf8YnZAbeOf1IKRot/kt7
6vooTkamowPbfqIn0i4g1gUQXice7fvYKYc6LlygDKlRC8Hkbz7ZTkE8X1iRTXlR
GbSaPhGCioEPu8YWfB9nZi258PG4/agHxCqoIJvXsCe0KIMpJwkQi2cjCDT55sbx
wWXaZ25/uEvADiHaUuyt2Ch/FgndRfrLZRBKmTSVk9FQG9LLjAJvoJ8qUNkEZeEG
UExyuadGJPiSZC755Uw2gc7JPxP0SvhVG0K9ZbpkAqGq1w3yON4HBMS+l2qIi1aS
BLlOFGzfM1ZmsTZ24Bc21a86FlWFvXQO34UU7oP17l3oeTrJqt6Nen9YqvP/ov3z
Q2AKVWEz6t+Uw6q7S6kWnOOLWLhwgKCLKwuaN4cBD+b8ia6Tl7e4WBcP0ytz5rXv
v0IfyjqKxzQdPdXBELZBPeReL5uI0A6C26D/NcQK9EZCBHF7zkSII8z9Oz5aqO02
fT0aAvUZipyfO0NoKox+3Wgz9u1a7rEAKYiuNoZjB6tyURXyGkbDCkECdHJWqFO2
xJY0P/SG+W5sPJHiL1KrWFGoYuZVAbUi1ngNfCTtJ0blyYxSbmtbS4B4Rsag5uHw
EtGMKPlCDXSP9/c2UUpj/4EY9/M4ZeKYqOW5AvAelsKZfCTbY8/0FemgMkG6GJ2F
kaLYErUgC/uj+ikfPjLmE1FFeES4uBhgaKDdZwti6ugWDFJxhbdbx3CizJKfyyPG
sbbaFo5fS8C4Dt+86w7AiY1AEPTHdPxtsIR7y1RuQm2pYm9ZT4gFTcl0JJ83mRCg
NBhCKWI+HFxzFNFiDTOBd8G41bXkSLZgWofCLfzdEndNLzQwp/+cQSV3ibxmdcFj
RySE4i9P/fQ3uWpA9D+Q6clGpN6fbHZUehv/mchaeXp/oeBlL4ORphMrH8Ys9ITo
qa0xdnIuEyM+WKwwIZsy5s45AbDpQoB/xXgRirkpphwJ4/FasfsVlEHl7M0ONUji
HJcilNhJK2sF8u1sj7CxBqzaje/59TYZbpxyHRe4Q3nVT9XqUlVUEu40h5y85W2S
BRIuIQcz4AupZZMX6Zn94uwFvbdYWWtdIQVBzLhFmr9bXWBAT4YcavfdVAXL4vaY
aMmhlNWazNWAFSNDGsSVBzf+bw3xjNT4S59k7W8s49/LWTC+AeGnzHdlEsEEC7a2
EHurPLxPEQQ27YZEpUsKrzqK5ip+Hgs6CaKOdkgaVLbX/jlx+fKXEMqM7wJMDvzA
WewHfgD/ziauc6NUr5QEw5QbdLpLpThGoUgoqG/d/nGEGq3+VMqgtVsARaJfjAAL
2RSRaNQjaQsGLOphRRV7tHTYhWtzltjkdJSSb7qPHSo/lRCq64uhXHK3fhvMDf9K
P+Sd6ZiJU5EluSOA1U6Kw/pzXqjBBmsX+6scUrR6A+voIYfWbjsVY7sQ/9+WAwp5
bi/kWnqhADDweOUjRhtGVIu5gMMdXlsXBXz4QRaVIE5urzUAqgqSMl2MbcZYRtKV
CGqawMpZAtA+3zPcLVs1tGba5kjoXGUOUmL5NimfSXbDFJY7V4mKELvb72Jc9iuD
969mNYlh+7C2j+kS2i6DneEPHKccyNlaFCZNEtvu3w8fC59O9zOD590G/ik123As
1X5tj8fKt8G7aQxFy8Wsvzblg2qi31C/c439hOj2MUlf0jul+eVceHoDDGZMqups
nKGzOJ61s7Csg3yuWbTHU72omhiRWSAENMc22qNzgGgNt4V9LQGPw7GHbNJS1KMh
/Ots2Y3tZQCprsRLEtCRJVJpdElYGJE4FsiN2wMkFovwCSGWhTbPhm7g0a/eXGPH
h0WuoO7qzn7OemrC7SKOVjpHLAArSxu39lBsAhCGO+aaD8lixO/TAIgsUg1913AY
Hy479AVUkbaiBnTFYsDS8comW/eyptIXjy9TjtMwqmvQHDJNmqTosqtL+8HT2BVJ
t/cugHZlBoKOhUKoqvOZWQq3pmID35Wj9+nID9jut6T+DXcR2//vTSwQNOz3/S7S
U0LH4StwbeynZC34ujZtUA==
`pragma protect end_protected
