// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:29 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
L84AYoqNB/inpz4fbnHTvmZvh5x7fNd2/RCDHRTFrcC1yAg9XcugHEmDIphX1U1y
/rPW3XRG2Z6tBkzmP+bAvULmjauCnIEFCnKIV/G+UmuYKDIjxSArL4WVYxeu8lb1
Wnf1ylwpR6nF3ehPT4YRZsd25FngEI5rTiyLFY80ojY=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5696)
jW4zHOe8SAUGwuE0FKjR6KBDDx/wuZi8LpbyqehNXb/E+FYOvaNLiTtzyI2o7rLp
isIu5+r2Ynp7XC0Iy89TY9CAjhmjcCIZZFkSbj2lf1+QKE+4IxhB+1A1uYeXctw+
sDvIfKsQ01HGUli7fYzeo7RTQHA9XCVdk67SEqtPBPRC/mvLJn/vQNuTXYY+E/BL
+6asR12yOZ/LL2BKSxudIj1bb/wovIKU6miJ2DnKQP0rlRKAq1Y2ZUVdnb4V2GIT
Egy1yNZcwpLCe9VHhz7MKvbPzJbfkhuziA/TCi/CsKwGx9hVdzX6NDioLLq5OH5O
SGu3PHSAofMKySLAcqJHDIWrOUXkOKYL59IywvLUUMs4bYTEIrkb+S/9e3MI6ufe
T5esZwumAHH0UrGdh5JlOSLTs1Mbs70roG8Sa6rIwDEESyRSH84KCdBFF5q2hyno
jX+VNphnqZMP1PVwSEAUVXMG2TQwUPbHkU33wLiWtmn6VTa9yb8Fxj4tCtQ4JHgc
04zVb0r5GLqqJ+0PF0uhuyQSll2XhWQmPQSF87QuZJZ0nOQ8xSFiupz2aikx7tl3
02XupLGLGXKhkKhDEx8jRtyLbCeCQ3yCX5/Lz4FmQgi4XAvjPWozUzeS1gXMJ7EZ
Todgp07+odRp2v672HVKDOo7GfNukRQhZTK2J8oj8TT3hCcXKM+X1Ry5pX9Yikr3
o4QcH7Z+OPDshSGxhSIaURymcuZFClERVJDXxN6SRwpbPumQNAZsFY6Cs/IREcyb
z+QZQ0vAlM/vSKgkVMM3ETlTizrKJclrzGS8TK0KYIjZoUKcRRkAY6BMNdug58mr
DuLDCYyxMGcrcgF9WorcnGQMMWEPwLIgxW85lNl2yBRNWOAXtKubnNKoTmC2NjCv
Am80jcHN+b8M87G9D+PLR5LPmmG09fGhc2VCRINrlbXvJKAi6F3k8nT+5InaeiTT
nGa1IToYDaWMgYTapow8SfR3g2+dgQ/xIuIUa+Wo9yQ1KHb4TgI6iannVTtegLzU
hGHBzKS3yKJROX6l8qMydCY5sdgghgh48PTtLpZ/K6QjdqPrcuGjnwiJ8+W1ytQw
/YiNl1Ng8lysJslC06azTaCP0EDJgeV0UNLqGj2DQ8kyxgcBdgXiZ3uwD+ppT5Et
WfYKpOzX1FW9cIx616q7RNeZFHdsCoRgucrkGiSqpbYfewxE6yTdxxy+Hq0q4Pca
P2uisBP9auOaHfop+hpZDw1mlrPc15y1KM8ybjL54bpA+3b3Gia5zqD8VQiWc4iF
VGpKvH5aNgZADY4G9caEL35nLZ9+SsYk1iYDgu6XpnoACT7iu/Y3zRPoplYuctUi
JATbX2fkENEev9PRIuYFNK+qHY0Ja4kqpY9oXF0HZdnBeSkyxDLTtitkR5WTdgOf
rMj1UsgQdXBgYZt2DjbEoYv4D56AQfPfnlTHkwFWPjhOyBy+6MuYkLZvMEuL7nNk
z517PMqPiZs/xECS8nMal5JP4bInR1osj8sYO3MHT/nSOKRgGy/VEdpmqDzKn7pS
AOptPThaXxcHfmrvjc2AIg+oGrPeHV4n4oza/SFr1FCBWEK/8zHGUT51RjMEwipL
2HNXVDO3d2iNf8kpHQ4LyYNc7oNgig0EZK4DltSYoSRpng6ibcJ1SIBTGGogvci0
1/yGKDWWKgcCzJh/1YsOCcMQc+d6i5BdNoh8YOMWAwzz9UAh4tAHgKMZ2LVJ/Jyb
gMi2wNmwJbf1wJD5po4qkgRu9C6kxDE00Gh4afVzZhcxTKBqPd7i1TpPVfRShNDQ
cHpbiYHz+dcYk65UYxQ3sc33dIk+r9Zd3dEvlE/dVwX+zUmr1FeGW/R/nWClz6up
iFQMmBlGBZTb458rI9vtl3gkF7iSNeqHsyCQXuNDDw7gQDuCf637kO3ttUriPgnd
MXr5Df1tHs+IR+3oRxgUjGRTcdaHHU/MlPbR5zmBf3Pbmg1t7sEjkA4yvE0vEgNw
rma2q0iO5OmbOyHG3nP/ws4i/a39V55+dIOCj6VrdOkRzy60R95/0SgqeD71YNgY
uaTUydMYHoViwb5Zvf/FepT7vC9R/eJDffxTEus/PVeQgXZKwmf+l/+vC7yNBRV0
DqPhlFCxvpytPi5kKA3lkOB6A2SUjE/aR1rV6ED0sUEBVr+5LMOeeVAoIugQsRsq
tUxtFjEWXYzlqT/SrIv15oosa/ICoZFx7IsGblZdIXlkAdoLLjNKKw8r5DDHCz0N
zCHTZVlRxHZjaF7JpKC+YgbJMzugqdb+ZF3nwSPyOz2d6tjXHnvXFN+36P5Vpwr3
Q48Q9TRQKDPvsrSmaQ8vt45qkTZAkJYiVe6aVfi26vv4pqxVgZdKyXQX4fC0oZj5
LhgAdJaNBnrvWnic/hEIRVwDDRKeAU1lgS8Pb72apBvBgbtqAY5P9ZBMrdvDG866
ZSU0ENo3tybApQuDWNh1iktQju1ELoPkiuY9ho2Z9KVdLltENw+/FGCjlhHFEUNi
NtH0h8gyKfNniNXtB3cYbdAiG8T0q7bqRIzoOaSyDLrToSs0Gq0SAijvTu9RpPVO
Xe0g/i0oOAUKTt482BeBXcHyRHZ69AjNJlkxxmUCMgo9QGTvjakNPxitIf9eK4WE
EwuMS+QxIFWpSJgDQg2TBEQmKMrxKya1lUAT5OBOkY1m31NOUjzKkHS0Mw8329EU
pgSOC56kmGYKg73hYRTcdMuCxdOXPMB/Ka4QtpecZOL9tO1HUTsMCBeZIixnXPMi
hfC2daYTHpdRG98/A+fz8GlXeraeeGmUREwUCSpxXVMt2bYKmgj3cvW8JYBddLFw
4tB0Uo/flJ89mfT9oYUuBcuSlBwl1JNE29SEIgslxYSKbDDd5MRovBn49sA/AEur
z0parL8BcNJyggg3/qx4EXYUqQRb1hqQ5EyxbER1WXUUQXv5DecYk2K2bWWtrvaf
vMacbn0GUahUtfV1hqzdjjRfNiXdtxmg3NWZEdc7fs+FQeg7HxYzfgkt7XfJj6Gn
UsCjbEe7rYttFk5lPZQsCdIdT9LkXk9hrAgWNFmZQ2MaZxJfclFMFA8NAxZvqLWO
cRep0DKgmCEIrTlDti5O9Gsk6mhzV0elo1cH2jcjlnxqAmLMtEfCo/YRsOOItotO
lpvOTsMEXhY+57nm6M0luKz8n2Ondga4/gp9eNTebw/d/iHamwPonBf1UwxlYO9P
uAm9dBJ27c9MidduZTAcCcJhmh++jQoCcDdX8QZO8Q5HLLQ+kSB1opSZHEhwo5uS
z7FaTRjYltHjaOMaueQXpwr7PUJo1qtaPgBjhejuFvUujm+sfK5JxyeFA6uB1U5D
VJ1q5ooI41D7ib63R2ot/AgO5+UeVP2uEG7Jhz8RQfj+VgkWBDS+X/FGzra33A+Y
Okfz8CWxH0+xUJ0XE8lFfiyd3o6RVMKol9hdRiUZx7FATcq2Q6uFgPH6vQTKqoiv
e34LzczdIOgYUPOLPDCbpru1B07Uyk8onKNQsGqLwaPsOD3R2tYPe32a/KchlGQf
Xjvb2EUHNzaS6vceGwh0ZiPZgjtLSRveboGLRvIT7LerhTzzdNqkU5EwmRtp5XOv
UUQM0B4QBT9kQ54aJl4O8z7/sMsl8Ja/vdABwMx2zHEs81JbKzKazj9jgzSSvNqy
IE8fAQ09rVvEEA0rF1Vpsi1NeNAE2ps+bwJT4PYU25+1cRXSNGWpKVTagHm6hqtg
E6QmHKg4GD8xypwQJjpdzEGSBGhjG88070tyGZvGNTNmDbhskAtxOlmG2mWeD0rw
JrrvYBsNP5eTvYczmO4N4hD2u/k+r7Hc+PLG96fzKd+E++e0cp8QsO1QZLcvPP3a
DaTrh8abD+6NyTo5GDQmpJaqlFBghzbWvUaVbQpGjXirON5BxFYFPCXaBwdQ7d28
AzgQgFF34Fi/2Ak1gv2Rg0M/n24Yfygx6VkrPtdHOj5JrjFeN+QgSqiEdOhzSEkl
iekY1KpIrGX8ym6sm8lriOKE4RzfzWyYsuXn0TIG1qw2M9+CQQ+MKXCcWTUmT/Y2
ZX8xXoHsuY2gIy3dHHfYxlha26aiRbgZZouT15KLdLNbrA1L2F6Pis/yHl+IJU8N
5SE7mJidjIswLffXyJXZe28tm/Z5ODw60b3h+4FgIAYj7Dmcax3XnYWUL3wvZlf6
ReGiRbgRqB49r95RmUxzeetjaYxb2EPY/73YMUY6ovdplVA58P6dF4UoXEdXUQhV
gnvw4deTHK0fw07S+JI8HQLy8vCH05Upz5G4vsj+weZsCmsivw12elhcPSGIqaEd
/ODZRKHOvZcg4WZf8pPJkssVmht7FrnQG1dKEioui7s1eJL7bRBEkCWW/lgicHbc
X07oxsgiS2ZDThuZBUX8UcF4JbEuthh4g75nlHtTo+RhUtX7Cr9S3MOiCyDmhLDL
U8nhQ9xjSp8DZAwmzYW524or0NvICiZEK37d3WVj9x/kXYGh579/OJAk1rgzWqIy
cfbKI0z6TTFBnKvOM6PJfw3bRdteJO0TJsXvaekmIjDKyxUFIvu+ymm5oy+zuLzR
xcah7Yb7Y0MNpUhCbHFcu5rw+K6Kji8Dw1tp8nF8Q+RxAU6EU+/tIbI7/uPP0fBs
srk8fa5jsaPJnuuJUZ26GK0FyhffHYQV1LZMgcQcSC3ljLTkeC8VdUPSrcwYAkCE
EiAzNgfev84yhUCWcLVzwep7JnlDnH09LiMlbtWu6CG3TqQJ0e2XfGfg4tTOXMr/
2gZaR2h21CTal0vw4v+LHiRGh0e+OrWl3ilAYvxX9nc+PNGRAiRDicO5jtLLUkT/
ygnCKOx7vR1KFd92pGLdT51gAiDWufCqWM5cFKeKu83KepFPWMJhpzQZAxdvsVPI
aR0JTiA9+SofwMYMzbrFmMCrJ71InQ3oQXVbfLMPNJpBoeJ83qLsrSNXX3FO7Slf
dU2UAYWFspuOVnbXbH1ujY5uYLNzLnvKY7PbdjsgdqlFeKB5DsGPVCVXbt2JGKD1
HqpAG2xqlFyGU9M8qsIDwH1Eu9xReUftVUT8aWtZjXRJWfBEWxwtNF/8A5HXzq/E
jTrO19qc6txN9P2TLRvaZEvHvcny93soZ+jTgwyl0wGrqA8AG6Py4679gru33HX2
TClGI97NC55YhVp6BAeJKShCgNbnTLUAl373ixaTpy1eAo3+NeenrYtjsM1hnWLL
zOCrG0oEM7VdOP8CTXQ+M9EvzoPNFQVGEQAjG7vQxLJnPdx/ajxQ+8PDOG5X1Jap
GjvfulipSGqYmH3drv+jdOu6TeMQeL442dCi42jnxrYsnNTvdwE1WZfYgGTlf1wg
vtYFd8SjwVzRBJeE64RAYj9YV1i0qRgWwDjG8eLaTfB/1+RrspdGtx0yCAaH9QL/
uBuTGDaMR1dq/Udm3UF3fSii3vsP0Nv2q5NJxWShgpbnPCAuMCTO1NcaAsGmRjOx
r54P67V6zyvAQ8QoeOUlI7g4pGLYVms6t9XwDM6n5108cnNPrtqHNuYNF8A5qvsH
j2sdIDnbR6hIg5eDkalnHU/G8RcTGa3LnsISXxu+NfuDLhw2eSM8UZPz09yq/Zgb
0LcD7vMn5KLbBxA8RyDEERo9xNceMK/+rdrJeFsygT+2WFEWXK7fLSW51UzNluhr
KsRdoqK3+5LEuTF6kclrW+jai9dEWL2Tx1cmNdRlqW7K2ojwAw+S+2Qs2wKjwP20
Xd4dhUj6hfXaQC2tmrbXkYt0BhAXebfq6h5vXcmwkDZugZPj+7vjWL4VhDjoeWHi
zSwJd4V67xNAbBVMVlvRhxrFCDZ+ZfH4773vyTVs1cGWPgPGt6wKHjH1ahYNttJ/
eEG/5A2rjqp+LsBfe6pg2uePuon6xEoyNAUnGRBYhfecxazywzrxmdU1F1VsmLoR
G23O+ej7F1w4A5/oLALBaWFRZVFehqypfQRVNcrE7b8GGvxhVAjIcwtz7TnmCj5i
tOQsy5+rKnaE+cFus1DfUmCOG49p0xd3w+8upLc6GIBzIWjHaX2+75Tak8xECNIz
mxF+KXEa5xElMoZX4jvXC5t6Fe20nerrY4itP2nZT7E9p1Q3Y6mPjvg1RfSd6h+1
eJjyav54IVf2nr5Gn0kooeCWznZvYIYheCoE2cEYRigizvGljPdxBWhJq7+GAAS/
77lDD5RVvKAZLS6NZB3eL0ukucXbSx3hN6D+3wLZKvCaCaDYvd8i/1ikrJSy7UC7
v8aYOlOD4Gytf/Zw6VQM3smJbYg9/p/Ez45ayuCEVWzboaYWvrXrkVcOqHFZPA5k
DlBDAW3cwQw0f1/v6SlaWAXaBgVEFnz2NXJ1oGDIFKYYE+fELdPeWwj2PKKbI7T3
/9b7RxSS/pDMSyLVD6QVhrfMcxsiDVa/igVTvqA9KCbqFzh6TQmazg6Xr0lC+xBb
jC6AwWak1ljy9vIDpLaQxBZb7cPHSltwvNO7HwgctFw0cGRMiAdPCLjTuQrTyda/
cH0m/9P1pZ8xdrVhtW8GfzaNBMsVmzI38Y4hZH6FPoGXQHYnghg56s3jTdWxDmnM
83MLAvgYdr/4OUlbNepvJ7Vin+3igCvZ6YyA6euitnDl08SaYgiTMZtUrCqzGnpW
lfRQDJo68NxUysihG+pED/8I9Dl9UJC3bBiliCYdXXxNoLIA51hvtEgKvg2MWPV/
Igos4Wb/vM0aVsIRnS1VGUxTO0FWdGKHfbiQBBLcux8slrSGmRo91b/h1NAmJfsE
l0Zg5e1BMSaaZ+DdQbsJUf2hXzn82wLR24kgYAiCZ+FS11+uDryDzW+6UBNHNYVP
irhiU+hhO2TqrXeTRnFmhptnsGHnEey3fAuH2AjhFUzZDx526efRZxuJb1LzGP2n
W78ONV5E7YCczKTc+VbMTJzcPTXmbos/P6N2rW1b1+1LrFN//6gKdMpxFFE10OCV
kKdwtc6bfDJplVMn2aJrN8yM2BygU1pGzGc22XdFlm9TUNW3czHFqlEjaasu17CF
pcEOzsLbTjYyfTGuEUSZa4d36EeQTap+X35yDwUct/I/uQftqShAuKmnET4C0hn7
+r0Mw/f9j06S7S7Zp2T3u2n8++m/q6jVB0lLWMDaZoywE9adUDhsTNRUbCHkvVIh
AAKs6lbWdJGFDlmG5AkuuBSxX/t4dVFvjUoPvHwLOqVMrxt5G4g693ObovUpCtiN
73DV5pze00MY/IjbP3TSjhLY+eeBsLTUtoV9JqVvIiPJvoXyg9lWj83v89ZBG398
4JtislrxuX+M5jSkydiYImo09UrWyohQYwdtiKtO0xLyvcdEYH1n7ipTHxctyAEu
8l0N3rv0j2OHqy3fiX5uuEINGH14l3QgydKv865RLDjSUVV3rs+jcvHImzkVTZAg
2jVjIFnbyB8I+7+qW37cKsb4cEF0HloaCKkowJ990gqza9YQWXYi9s1G4zRbH6AY
Bhholr+rvNrkAV5HdLgkkVeexfCUfBg15IHQr8Etuog+LSjjFKBPh4w0ptKib+B0
L+/0A29gAF8WqNWK1cOlBUYutO2t+GLCw/wWhsRexideSvpdH8EUlDpajuRy3ohq
lVNj+96dJ6Ljv3/FcOlPe1BfvIQpFUaCEKNTulSSMzY=
`pragma protect end_protected
