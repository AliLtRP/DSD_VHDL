// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:26 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
U90J9cgala0yhYVnSR6+1d+xOZ4umod/FAiXbaHGzNuSeO/iWQWC+MVvbH/dbRMu
DOtFsLUaCC2BSn0vBZSQ8vozjFU3hR+FLenD0+c0eVTSCckErMcrth8C3yc4jNzg
oGSZzGnAa6YmqTKMUl2p01TMAIIHyJ/p8cE5LKv8mTs=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 8448)
ulFiB96XruhHI2HYHm7YJUrtii5AYDEgz5JXbE76B2u328Zl6NCmjyd9tUV5Vxxf
jOQ+fLuUoXEohC+WCfIlynKE/kCy5dHYG36b0UOkMXmFZeACgtxCs9Ez02nudL3W
qYetlEVA2IkXuE29KA26yCzcYh8y1wcgp/L3Zvo1Uhq24q61IvKKzwvxy6j/nqjB
p/LMpXVsfZnIxkq8U5472lO/Pma7GiEHgTC/JdDqomoue5Lnfx7hYBgXdLlhu0Db
JNt0BbKuIpIlYXQVujoa+fseQtztSJWEQ5hF3CBbj78UgffTQpFR+t9Fg/yqcRUG
fkjPoGp5N41OqNDk4SwFz4ER9LT5e1CFtGSgg5oTSD1AsVsPj9N1+nD+feTqnF6l
ENXk+arQ6OV9pKc/RY+pgQeJ5ccSrYEjXsWdYt9CzHhQM2L96vkhXj2tPRz8enSH
i/qqNUq9QY+n5ZKT6RNjg03rZr1fUIK5RahAbgQ1C5O5Ib7HKAAW3XsNdO8fOWVY
H/Kd6NhANtnj/nhkS9wPhWleFB62QzjX/njXg/95EoErHAlDZdjmphgNT3LwnXJ6
bXGyJlnTHjFD5KULKxpZRt0GDIOnjiNb6qERs/15nfJPp8yPfUkwlb6SZMWoUJZh
fNuIFIg+sl/yBSyvb9GHl6p8vfXU6vBd9YklOHwPp3Dc6P9HRyclPgEEPAwpbCDZ
p7IU6qQ5FkZoo5bej9lg3WRvjuUFa261yfMQ1bZk5990GmVkF9b95qF6Al7V0W7+
fa8ORtDlWNANfj42QCwcAoBT/Vf9W9Nuzl48cukp1q2VkfZVViZVwywm5JqBTclZ
jLf8SGgIXarVHKwd2i6z0KoqowlZArcbHP/anPyA+S93xoTTsXGVoTSvlkt+lK+m
ebZKwyXtZjG33AlMMFIoqWg2+oNeBFfQxm7RGraV+0V1qPAOjdqyqYHTuwt8LzTm
Fz/V9h/MVDHAj71miY9W5lZYb2ucuIXNZGL1Kjf1tVT6iCocS8lQ6GydiDQT3YHD
TGq47INwBNpXqlzilHCvaCR37yk4TB6GG2g4zUsFEnbd7OxhCM32NjW3n/Kc6+Ng
gmo3zcO4iJqSh/iS2r64C9fJcilhAQzJuvvBG3G7lWmXLygmHac4jxYUH6AO5/em
HnDu3dESvfYzZG2vjvsgGomkDNn2X8CqRYpiPGh9JJXrvMwAvvf5Ig/u5W83j0xH
vpiCRPS4ShjuqaancRb0K74hE5jPm0iEHH7DzrP6tE5OGaIIXK98MJv9jdtDVKTb
LRV1V+wGJs1wm1qfmny+EBeKEaLIzxo89fprk+IiMt+mGqcM6ZRRoxtefGBE4hRx
UDAXZXregr5+y4XVcntLL+S6n24PV6gfqisMj5jSJJliz0Sf17pb7Ac6axBM2i61
A6edWmZStayhYOv1D8/f2SVdC8o8+jz3WvAGQIZeorNfKEC1ltNtrKCZDNbp46BK
8I8nXiYan9U7YblsSBCJShUQckbLhGYvrB1bZJ0QeDmWcVXsPrJe3n5A3rWtlacy
plVtuL85k8hp3+xc5MiDrcgsjkxZV97yurLs3QJnNEaQjbtNdBSSvd+p13Qc8ZV/
jqE1FBKVse3tXrpb6XW9CDhSJQcVfczD3W+vr3vM4yAG1KVrd8JEHSJflE/BHqn2
ndr0O9rbRbEkNxRotDcz8RL5PttgQIem6afBVxOhrBrf+td3xOFNPb9fBVTDKNAE
U28ne8bByPrdyGUOGK8liaeckPrJMsJw73p7bYpPZlnLG2CMAZqiIVGL4rvKXAf5
xKn/DDmqZZmSIM/HHMNSys+elz2yQ0yzPb8o1vi+s59oIgz/KhOGNcmEgO3eSew0
TTEPDhq0+SjsHdzynyHSPQts9oC8dnlqizlbAlbHEj7P1iUyJzdEYLOS+3X8GqoC
KZb2rCKvaJxKNQmjPmlvh9WPQyj4voWfzjzboY7iETtCNqAcrObqnLccWpyNsnEu
MdAxphhoYLUyfz18LL6uZsgIuAwJ/B66/OiiFDBXSyLYV9DhSoYvJNAOgIBUi1eF
cT1JR7GpFe3MCH+cIKhmVAaJw88LuAwV1zMq5hSEho8J+tzAwuHShb6gWdBWxOMa
4Kl8mOdI2IzYRNVd+TmpFofZLa4cfwN42v6oxUoBTcHNTPdYEpt5+pr9WK4PsGPy
VyIWg3oDc5T+1Lp9Ka65rNOyUbtJlLeLuVq39yHmn4FdcmcIimsphgbhvJDSAOPZ
V3MRwxzpxIxN79DOPpSBcIxwgOSBAQPXep3S6nNjcb+Uqi1cnTnIw7tuN8pJO+WF
S8j7NahuRXeq7FHCANGhck18sx2sr1pcqIZblNpi7ajc3vDV+ylkHI1xNLCLb0QQ
c7FL9Uvxtbpptysipc5wxNELW03X62KNCX4941ExJHzAX4UQMlRYOmukcHBbXCGP
xuM2xnzGN6XRfYjIhMiTjaBmeCUBB7arDDlRSOkmbFNSjTqbT++UhJTJhR+KoSW+
U5rXwJgAczFr2pQpc2ITzzSKRHXeZrqygoQjk9GrVJqrEy6+PTquLTZLeUIrSTd2
g/90qDuUEajiXQe+d7iqJQbKfCChVO0bbSNtPjqdu2xAbmjY6VRh2XtFdV/HeoEw
E4eeuoJlIPA9TTsOBwj1aif2cy3jY0NRy1FjBhRCPY+Mahgtk6qI4hRgWspbwrUx
7HpTDaQcVjLpGNOoochcl0QKBqHFOY7YOaSuA0WzZtESq4W/RDGdd9oHcwxCOVB8
4bTcMrzsKbCoZqPsSt5+t72uCSsYiT9JsP4elMXpbHIMUeYq4HrquORXjMaaSe0h
VvYbGn43Hxo69pi1NJ4NeuNFvSXnTsFSnrelI0xCFff/AYl8t9QItGmsUmRQYwp+
OQRdP26+qUBefcwBOur/msYITmZXrRWbsUPqk3xZR6FTOg+UJ8QcZVVLPM6lvM5/
EyicgZ5RS3uX8ekWAh2Jz/+pPolzIWXDwCMfT3zcDGbripTA/x+4yOkKsya9j8QG
j/880qUc9sIONrE0JA9QxUT3Tx3GJkNQw4ldQF7OuF7EWErN6Lyfs7ObzoEN3XsT
UBbf32w6uwptux7ZEEcjQRn26btKP0+4XPYFXPPhZ5/ZtFPkFagP7cjVRCsj7LT7
PBAB7r8fYeSl3VI3SGflI7rCflZ+22lpIkmo4zhJMHXXtaS7kb5nLL6UWRB5q56k
sMk+miWYV8j967+ABquSNxjxJz/P7W5PemZrQcnQ6iUC2pJ+f5nw9/+8uWlscfFK
lBLbhVOGejboVcdTI2gbgUybvW2DDZ/4tr5gVZOZb0ExzeX3wJOJZyqi/+ySgXen
Z89m+SkQcQ+pD7mCMltBmi+HwlVTjUDQ8+SUpbUcy7dXtra3uiyAe5QFeBhalmMD
kuVO47oGZqGE7QD7JnuTnlH0p84CLImsgeF+EB3zI8wqdErP5riPi+v1xJCwmyU8
LM7FJrQJo4QzXsFvtFWb3kcxoLg77Z2n3ZQY/KvRQ/ZprfM4OTV38+y3qtD4fviG
p8RWRTQQ/5Q9/ETO6pb9HzSxOxvUz5yNeQ7SxUQE9s3bdORgDWIpyUMgJlh7fxEX
Ntwfm/op6kgLcsIrqSGyEZtIf/zbhrqd1r9ORKrkU6yEojyb1GnRZWyYP6palQRK
wzNoKlY5n4pCChAsfC9qeyWiP9s23Y3qsKD7lavKEwYdj2T/A7pGztd4g8oOeMwA
5c3wy15s+KRbDw0pznJ6iHm1d74wGZodAGR97rdpHHjL86L6pu/f8n3iIuzC1zoV
7+CDQl9ZKF24FD+oazflp/az9Cus1pIA0sojIQkVKvvfiJUV7hgLd1YwPmUJNiRB
5V+bS2e1Tk1QAZd0nTwF5fp5AUyAYapnHjDLIdbcoHvbi3qGb5cq8Kutp562G9fS
gUD1TGBMiiWsBfRGrHgna8yQJ0/PMiIOA2OgOP/mMsoynE9RXlwTKqJq7mDTPgj6
/IunRxfh9bGfjCaVH7smKxjpdwVWTx18jlWnhTO08T1f5fGduUdAbuQjrglaML0q
BQRy3jKzRE+yiLta14HBaAFNEXz9NbHLEdFYHgGytaO0sstkB9mHOPH/S2Hx0fCV
6FFlpjlxvJb6ZvBpbBJn5QDzfqLYz4LXc70w0rtBoGxaaxI6RDrgjjS1tj82C/Z+
j8HL56X5ryL3QHfzbSzX4VPhTVRRSHwWHaJMPAgN97rJqO2UggecTUxJRR7Iyl2c
o/s22aLA2OpsVzxst4bDM0EsbZwYLDJJT6DL6coQkDTH3ETHkdUoxVoPlVw/Dc9l
jw9ghPtNkyHCOV7A7Rw9pNBh1WsV/m8Vj1SK60aitong+8aq0PBhUS5UT2TDAgpu
OsHnvbC20Z8f41WOygEktCUBXUa5gs1KboUc9j0ImAUUnLmK9ka/n7ON1LUTPsyg
hDXxUXNFxBBP4i1hSoWlWvcX097YVa6EZ6w3gSY5K6Fvwn2HtPoz36y0YqdegjQ8
2TBfmj5i6TP60edUUBbQmtc0cydPk0k5Yb/rNh5tzCWeuUH+83BbxMLBcip5y9Kw
RIpJ1hNSwTnTwYkASB9Z/K2r/IQ9VUPLmlWadpbXutU2FQEI4Wn5C4llzZVOA20Q
DWJadyILtf+S2MyWPNYxXZfZk5ZM+VsO8wZ7yHGx//u4cLb1bOLZGlz1Fnm+BJmj
GuV3AV8VanUW9ZKbQa7mM3TiLWX9sAUW8DyhBxIlfohaEc6F1g1GUPa2Cczbk2/u
iJbgColAMS0IPkLlegLnYk6d7iHjTh6GgOqFJ3186pD0AcHUza5CRBatA38et1uT
qoYmOPDHbqC8KMu+kHLmHOnbzNZrHBCfHFaOALX7Vl05RcEMTK2u0IMQoqTpP5K0
Lu2UAY6gQ4guRCInvpGZl01oGrBbn9yBX0aRUB7Xn/e1CN5s0s4sLHQB9mcVE5v4
5GQtlPaOymUkQafYitcY1Px3PhWAZLaGqsibgsYjNRGuvVs6W3571oesdEFBaqpu
Z4GDRmoKMrihL6jHsQXKiWgVhS+I3CMD1GVgJUBoCu0ywKVcYK6VgsRc2TQAPcTl
Qf3jcBeFQZXtgAMxJ8gi2I0QqHt6u7/wlEkI6OYmxj6qA/0WHJGHoZ+8sxmwFFKv
gUBQQbPs9EnVTSy5f9MGdFlGNrX3Zq1i6ytSIHpaM25GicoOIjcJHNRfqA6/dhvD
OjDfJD2H1n8YnAfh4jDLeTrsluwzwQRjA0eC/mNw7lgW0QKoGvViyl6RyyWojD6L
TvywfvuXqAuer/3I6ms8/abdT3XdDbXvxFNWyAlhjSsvwASFQbXyMitWXftAW9hs
To84ZdXXyw234qP80SuPtIrri//fMwxgzE77uyLUEGJ0Uz4IurHqz7BAa31SjStt
fvCg2LBZVrEOaxCSHxDsVmEgSpymflOTuegBoli+5d8FSZU2zzx8jGmThEUiRib3
O5PCfd3FAzWFahn9WXCKQ119XCE7cIQr99ug7P7DKVQYKZF8of9EC3nmhA/ob4j6
SEqRluG0q5FthiIHjTx7ludDjxj4wVLSGlN5EjNqbDJRHbbJ9K7WlproLYE/0MfE
o0XLi6lQhIN3OyHcUo8l47CDswKhrfeUPPutOMVBeJHqI+/Ec0qwStGxQVuvLmiu
0jqfMxWxvVn66SzqGOzRfUyvBAcV5HaVo4cbmzxdHFwBl2X/X1ndB+Tm/x9kAHH4
FjrQr/DLDOjP6NHBqFeMiyA+mWTAu2FJf3K7GRgUhlRlz7FTHXUnlrE1+WYqEBpH
Xu+ioY7jjtLB5nW3h3TFqCBCyWE63zf8EfQMGBsIVlPgVlOLhaHnEnwOwAIX9uFJ
ya58azl1If5KsdBThDcLRPrWdxTpAFP4M+v+5zkxKMKMQBrqm+Qi6m9AQUOO0SJy
3ilitYp68G0q+J/vYw3KiXiX/u8QRf/F6WOXnB0TtHY8qKJgxqsAr6ZaoWsZJ9U4
wwjfcCJSyWlK+Z4PzZLxdBrXNVtf8r+SuApKSpmcj5J/26Y1DZpNcJB0NbedHr8g
XtQYQEK8+RvlWECaU8oB0CJGdVBBQBuc6JATdU8Ack8cDPL6IKlE5fToS/qlMAT4
T9O2pHsEif6Y9/xG8oKI+YMwm3DiVKHZVTf0qckRCsDTBPFSmogJa5x99PGRlTmZ
aGYNWzgi5S5EQhC0g+PaPux2kvo8SwLoHUNr0u9/1TE3WuOaj8li+NmturgAqSYq
BuUZ3WA+pyZ8FxLBHUG68vgdswdqB6ajNC5oWFZ0847IftQf7f+CwEcJh6liGoVc
wJSKCsjZ9LIJ5y242irUZ8DsHzS4wdftziPdJmOm+cv1CJLPgv9dz7K5nHuSdoba
MwLAtJhvwASNZ9uIL5aYyQrBfK8kR7rJaThE1OQ7HGQLTwogR4MaYHas3LHR5ieL
X6huaUQQdrvhqaTBveLzEwx312sIQPcybWF9gnPSKj8XC7a+PxDS6+TSWJfgAtwi
JEOHQGL1Zzppb8dwRA70467KHa1wVDa1FfMolGloI8Q8CflbpueuelOVyt0LP55g
PmAm4VolOovXctIXWRjn0t8cFb2X4/Es0udp+jktNMGG2DqIuW+ZfLrJicCkeaZ+
5aMgZi379CbxRWABYscALSc62HqD6onnvDkFAOl6aBk2l/WMuieTWMX4jHX8nsnS
z6uGy3nYDM6nYKSPyUL4HuP1KGeyJQVAf0mUdjtmxIa6cCtv/iVdEAc64S5TsoPv
+46NHPVV/mQ02WPX5F7itRWn0Hu2XCUEnC+JZLgxsFBpmqZO7DhKVZjraVvWWKEr
ycRcOfCYCEMHppLZ+rOWDhypwHQ+6nFVlRg9jFzWiK4bJn/NPcn8q2P0QiYXQmtJ
BoUBmQbO2mc2LdpcxyjIVyZ5txnIZzU+QKf9ELnA9X/Va/bFARp8bVH7Kw2UQoK6
IEUpM95B9dDjZToyR67RFb2K33fN/FOO32yxdQ1JekIfl7LS1yUf+eLawASkEqAd
YfPTBA0MY3hgmtllLdg5UQ2lE1jHmRfPW+0sV/U82tvwSUjMaOgMFQWTzoJyT62v
CFH9Nfc1M9H2q5KT8wxvKvyv9Mtti25+t54VuDq7wmBoTeIMeP1WMBhgWRUloiIX
izhjKV5oNPJuMKGvvGJo+Bs+F6Gl5BN4Ei/xXxSdB2YXIuwJNnI0Yd5MQcHKy4te
MWQUczDgatoIbBgOPyATfkUdvZR1nKCzgXZzuwgUTXy+UJPm8j/OUSjxR4/ff7jL
Opfid5xRbJnz7sTGbLm1LPaCunSHLJVUH/pcuxc9REKke42FoD9caU6FV1XmGOdn
Yr5T6oYEXSX9zjZpak0YzfAz0i0GJIEmLEyHlzbFko/+WK1lUGLfNoTS7l+lw6QO
ov20+c++9SzIZ1DIjQt1ut1na2+WzYV+UBWI2+dF1M4CjMiE+4KKvXS9UhmJpk9e
iLa+ug5OButIIHqVCsJqMkX3jti6NwbkWyqKQGpn/9cgev2Gn5i7OSCXUyO8wtpQ
CA0P/xgmx5T3iD990NmLMs0uurmeMI8RZZY0vtlpQnP0ABqDYs9/fctuttn/7NAJ
eQ9mvlIiSi0wAL+7dCJGrm19SAxCretswHmA+27K1IWuCfA6tJEsqci8/cx0fXtT
v0ja0DOvez85JrN99GJJCUv8eoazPLfYCeTn763vRtD7WRQKLg8gkzfYEvb6TMxX
fjfC9ripM+lQi2USbAWoAffh5E3E0SzwIKAnp/QeRc3UD7TX+6YHTZ06BhFB71Ba
KUN3W33NkQtKucB8yFMEMLcJwBPyQKTsva6L4+f7sUFJmThif6utnpnXBAGZ8Uao
cpdXFFTeBBkRDiD3J4ElbdrDk1UFNSBBzothriTpqhp9Jp0gzHcHyEPWaU4Yl42q
Djqx0INDtFpY74Plbe6SsqZY1KP8FV7k7LHkbQMpPixQ6KOvGh7g6Pt6mSem/5Kp
KYSUVIYSu8t5bhmUHmwPnUdcK8QmgYZg4zD92l3zkM7AcScOxZQUFoaL0hjzDfOp
RbtdE5GNZ+ZG6HWj+L1OFltvO/xFtHI8/IpTE7lGNStgcgU2lFH1YlbLFNRO9+Tt
R8TKwlATXCSnA3xcxD7k7cNQbwmbSLjaUWLVsDqa1fvyFg++a2fAZCCQWb43dV3i
GmZw6htlQi3qxWsJmFjfldXWvZu1VO4xt1F99hkBXhbBujq1bPyoo3FtCgPTkxNk
s4OMkWAG2xEeQIb1XqZkis6IAtvBxdAwinCaizWZsSySL8tKv2/IBm6QvT/nRkrR
ug64DNXthBMiPmx8MPv6WZrQFU+mPhXiQG1O24+vojdPK3Puo2PoCr+Mj0OyHBmy
x3/QWuKlg8Ra82g7vsAuo1gCCxpO783VCGj7zOW9hcf2rE2rl9Em+Pa1nwczYyBe
v6iXzvnk++6MA+9qQk+nxp/3XGxsfDy+32xM+uvrSc57qqQJIK1hX9He2orV8xts
lMmbE7qQX4yoE0f1NAi61d/cE6pJkmHYCZBw8eHrWe1043J+0uQvzHhA4wAmpCT6
UCBLdQ+GM+vQ/qf75adAE6bjlp6jeFeSpzGIHX7RNY74vASQnm5NA4yKtbwbTFcZ
8ZyAbrafnEU1tTq8Yg9vsrSSnIPvQ0QTI0zX8jb5ZVgeidb6XDJfiylrkdNfYqUI
IPobW/N0h0wtF9kdfPlNalfMc7Z0SPTsIFIjwyt8U1a6+WhtEnjc64tAmqqlXxAa
AMU+6UdpIAAzbxDSX1bOnpGom6uJwbzGsjgosXov/DNPVDFzffG92t23I4esp/nH
M5yAwpuHxoBvhtv4cCxLfPJyM815m7HqbDwa9Lq8b916xZMb/0JrobBxw/CYmRlh
+7gIjku6ZgsgGH4LWp+C4UOvz04Br9ULsJWpK83cFIRjc9TEV425K2bZjn6kr6Pg
9zQg0GChKyPh5ztGwbucnVu/Hd+p+ThCZ/1TTJxS/4P+tHGXM7ypGk2vJaELtjp0
HpeJ6SOcWZwIQMFUH1lXKYiqSneB8tP7q74muXtmobb0PJsKwjlRakzbPC3cuVFE
BdjVCDnbCbu2I6Jwpb6rEEQae5zzUbRnQdSegFAbtFjmPGYNUGNrjAE7emrlfNTQ
cQ/DFOR35mGNSbFLRKL/3f8VmWiEzS2cMTqxJkAIoCqYNa2yg5TgbC1J3AZT4SIt
OakS/8qlN7uOZsuSMhTIiipn0nnhDVUTTnUxCxN7H0wQZn1lQyW2KTSAzUC5gXnu
lRJZt7qXCp4ynksOGoviorjONXK91ZB6Zr068z6dfRIIbarcB4+nzf4oHFJLbDSC
COBm6PalGS18OEFUTqV3yxN09ZD2AXCbfuBiLJKr37ZXmjI2LBIzDpkhwDFmaN3p
GG4wgyXFpfSvNzJljJZA200hbuFywv3VSVrE2u6QvmiOTYSuxZIAj0ONnnRziUTI
kIz12uw10l0EEd4GF/X/wDyIeDS8w76DK9JMSXbjSP2e9srUaY5KfzX5sMQUb+au
NePoc//J5fgOtyauu4jifEiAblCooIikY5iZ3UDI2hbVTkGylt8DmH2Qf4aA+GER
R0RoHUPvbBC65mibwsT+vvtQpFAK2jpVrqcBUZa6sdNJTg7kRMMT0GV37NqJHhIc
x2X3qnLKBA56T3tJbIXq5cYVb2m+7BJ2c576j3tkvVsTln26FXN2jYfV5fLTei8g
V1vso3nZx6al8k27bpak0BidthOX9i8zF0C8Wg9PTbJF3IfTsxKK08Mz9IjJ3kZO
sXAyZak7J1XGIcwEV49/wKSjCYkr+q1Uf3RyxEM3tX6SOH7PWuzrKE73EcDGLhN/
nuJsIwdQAvZHCNyNbtUkVpR2tFFe+KkPE5ulNdjZI6Urdz21pBED/aA3D7jkTIXC
JFcvMBwh1NPBf4OIo574MLpkMwNMwv4oQtRXhaiwi9+wRCM/gKxcsPtDgGgYRUlP
1XQLCm9wwiAuFOfvCvl5HbY2pAL5V6E6p1aLqIrnjZ0WRYbCap03zL3wimxIjLak
jXDTzMSkst6Y/aiwpL5BSoM4P4Bdv53jAt1zbZ6GyQJdzEBztJG02pQ1ZwR86b4T
+Ju94MmWjHlxUXE1EbXz9OxLqGpFF4Ir4ShCX98VzCGlENt60lf41tpITIPe0zaF
u8IRNRtIl3JlAnCwsjrflBpP8vSR6gHxtAKOiOPvJdS0Doeg/kioyZivLGhgAqws
LV6wNuf9WNRuATbMxkVT9vhXJu0OF69PsS36eye2yvWSiMosmUXJjTIWqWrFq5lt
EJpWgk1DZewHnOLI8VnW45RVY7OCgTkhDGwb4QGCFsSgetTfV54hfG/6t8OCdwci
3xMh3o1q+a3H+lTfoR2rdmoaJcSM8S8sP5F8CvLJmy6aDi8M8KlsqZMevMmeua0Y
105AQWHVlvuc8qlbTSDl9TSRlu9LCF6nQuacUMiAcEOrZAEhO5hMvO1IfLVeF26e
0pLe2sTYB71QeFN7YvmhSdYcKvR0gtVynIbaL8N5SyYlu9gmdRZ5dITMZfdGSnSt
67brS3dwc3UrfNW/q1e6zjTbGs60RKhqODHiYcxk13V9+t/K1bwT3p/2oxxie3pb
p/GPYAT0FOPgsmxAUQL5TLvuc1APjMe7IEEPD8+GVfUNEqBAcJ/xm/IOReGXV3dD
Om8PT9rH1vb5ENMefAvIr/Ur5jr0tW716RURf8UlKrMgs5dTODhOsEF6nQpDJ7y1
qSWd+fs/2rDiAdmthx4vVgnATSh15YA3WTHhzphQAmYqC/GRE0Uh4oPa9jpymf0a
NV879pUFQGpqQW9tJCDnzG0mO/T3hFS3Ufc9OAfF8bkD9GYDDDqmD60lUdvNSS10
zhxMyr1jx+9AggN/kQQe7XRn4Xr14WgYVwcHAsHrYi4iavyVUD/5K2iNnDMhUxVz
IC/DUEv5hb2F7Bvbkx26UR0PA9LPTIFbsQBFKmrZ/0F4fjfnpXtJPyjSoRze8LoY
GgglTGxrkL/in+hceYaqXtxt+prI9SvUk2pn0Fdg5H53Yni9H/zvGG55z1RA53S3
zDFnGphPDmba1hsot4qEFcqhOSgkv1q6Pkk4tLwH2UwH31Ah0yqCDEpSH46FBFvz
gW6X7+rDN7BvanH0BUYXmwL0uEgV6OEGfEUrA1WqWRDT0g0mPQn3omzV3FwGpkVL
qs5BeFyLP8dH4RhNY3FEy0L2CK/WnbuKa8jzCOPO5xEvzGtd9dMJy8F0hs902D3r
Wcezj1uGANT0ERxDuQ+JUKbvF+vK7BG9gfxaDvrn09IQiQzdnAJv8VoxR3ffWWKS
`pragma protect end_protected
