// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:21 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
PKPT0GY+4fitIQ1cN5YwX9DtBg7VepSSgOgnpnw3GEbhpZUE8pxkI2aIN4w0I/vg
1QWRCg2lOVJJHMIvwRzPpk7fUoKz/0+NmHqAB79HrjOMeJ13nXC6DI6Lzf3XGLge
++SfxHRxeQGF6m7lpEmzLkVL7MtNUM0hr1Wk9j5BI+M=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 40624)
UjUAYcPoWBdX22gIS1ZcxkqqB5iAegqnZSqBwsl99TItCao2KbzZGTepQPw+Xj9q
Kuim5yK0ZaN3aoeyRc1r+E68BcGc1dfUrCgWcZvyih4xEob4J35jcEqRYZSsMb36
Ix10dIM1GSg8CCQK02hlXGZiV+7JsC5flIG6Kjd3wFjcAwgv1MYvUFzmtZLBtGQw
UeijDA3ihkBB93JlU8VK85MIBwjisQ2Yk3BEKGJHag4EmPXsxFwou2QkOGmMX2iK
D6biMCHqZQ5MW9CE2SjfJUAfhfgvqDdyvvNu75VvV4/DDBj7edWKqenvlyXDW+dA
BAg/tI65LQMEWcE7g57hn3SnllHfHC01wQD5s0z21p1vM4fucXzTgFzRCXMdh6nL
G7Cp+GQXcQW3J5IjMCLev7mM+TuZsoHwEpf/LQaCtH86D7eUToHFcAMNAL6Fx2HK
56IpANuj2JLUl8aJNd2VlFlK/sqc1pL4kl2MVbTZqxvQ4ZsjgFuK8Hl1My/VZ+ch
Y3Grg5Rr5aWCRpO/EBJSN7v50i4AwBHZBbG2CVIvktK/csvwZ6qE9HPKaoMMkBBg
PVjPhKOdg4TvthVSkUNOQZ025AgBOYGqM46xsY4TjHG45jo5YcOEhng4qUqN6t4S
o59TGrjuix2yhxHgGGJVtBCuug5jXFKvkhmQ+9ST/03Vu4DQewC2DO6OAfSSoLlR
Z/UbISzMKfUjGQlMcwye7cO0e22JyrSaYj0r0u5F3dxPGNEntydpCSTLQvfONaIE
SCsLMbzVCP5cGI7ZbTNyv6pNHOJAHO2/ZCAkRNeu6H+Rpg6jsYKr0c0KaFqWMzeW
p4UbdLpoarmcbmI+0hE7CCAOzk7msvGMZaXEP14+Oh2hIipnBNx8iX8P75zXgkZp
HkaaYPpf213vQk95gezts924ahjS3W6cNxOV5SEpKdHiqy2QM7QsdwiXF+5OXnEk
YdX7fFG1zu+MfjvWYmcv1WSLDAAVuSIarmhYN+cd/myNMu9lvMYBLrQwzjC+hkh7
b68gOgRi28s+pBJiF2WqK+kRUY/LwOnGjf6tfMva0KVEs6B35E8LXciwhm5jJZxv
X20gd3+uGJpBU0YZKLDheAcbd5MdlhF4CjGlXCM6CJTLXQn79lwVIeWem3GZxNe+
5JVViCt9J0ZrJyLxpgkisUhDtOyvPMAMWYVkxbPKA3Ti0rvoCk8afGFahvC+59wR
RRyfoRZQxWmUw9i1EZvYkNu9NfcdE87njMzcFBI/gW5IviDKyi8daPzggjo6OSVZ
JGXMW3hwvFZaxkyIl0DD4ycVrNCbGtgAVsO1R/WkQ2QN1/26quT00lDEtiXHF35k
mFUQtUdFbWWCDVMSfhPADUevh5fzvkPrDd5uX0JGRUCfrgkVLTNOhsIBj14dMTIe
b1Vxo241enklDcdmN/xzVQtbxnLPykw4GwnwGaH9QSdg9W4zedekXxoQ+ls4/v5R
MVrzWqagXCpMTc5VBYz5CeK9iQJ1U+at7G3rm0RtxqwhrFmd+Ou9EJ5bsztqqxmR
YwqxodwnS/sN6B9Yg58PWemBFtfqKGYVaKSIEB9PnGqd/Ir59F1+4bGNSFGjgbA9
uqdiLW0TPQP3ROvo4XdhorQ8ageB3jjHG32uJApq6IOAVYu4BFniHqfFBjLRLDTi
SsFx1YIiU3NMjKjJszKVK4tsfoXx5qmU4zrxREjDLsXncQno+lJUHdKYp69B5QVZ
O0AZ3u1O2wl0SWTpomigfcXhq9HMkBmPhXBXppFQJ3OTipNSwlYoQcV1L+P1wN8Q
sh5AoLFhPrIrbC203f0364e/0tjdDBRq6BOr3XvrSJwKBibJyYsozo1RyW1nbd4h
zvqvl2CUezHh1oIUWv6m2VdjayzSHM5+cMyJHjz3uiM61ex0vDx8IhVYzdYxFkkf
2Kp8HvzJd9vj74RVp+t02sZhXWT94gMm0j5A7B9rcw43JX6PrWrfO2uydW5MPXaV
AedeyDbGNN3jGBR7+YFXLC5GsC611D2W8T/UmHe69BTBWtWaqNmf0vR8TTz5tH52
7Txzql/wtIeoAzX0TDl0O6jsC3Y2dhLW7YqrRU4MqjO9BsWcHxNigWunwHt9Yj2n
lYbonrOlLV3+dPG/ygYmjAZBonv6b8u0mOcoo0G5Cg9pzl80gBeNUL0uTBZ276Vn
CsNdaQVTMgbwVp1XNy4izZVjKt3GhiZ8Ugc4PTpmFtkxm15yArkxgnwf2ShZOvgu
5+u2Yy2KzNPGHlsepdUDhS4As2+QRgjAG6y7UHVhrY2bvxLiIw03RI2A941snaeA
z66WGLvtYq7z7Fcbba86yc4Q6B0U6tkDixfrC9D3f9oYbyheUl1cyzjQype70NvR
bV2Hu4gBGTnJc4W+hTgmkrJoV0MPcjzIa3EdWkYRerZI8CCu8t29gWqvqun7fkX9
BJZ4rIyZghkUeHoWeL5cK/r4kxM7KYW2C36olPbMNBAAUbpP+CGUwRpW7fJgsctZ
8h1UjYIyhIjyMXmCZk40vKlpOXkHstzquTlCtcxEzR5mfgmLPUUVB08ej+tRRBM2
pJN5krhlfiw2RygDE3klEjj42A8c0rU+wY+IT1RIe9zNajQ3LalILoMbfuAoG1P2
5y2Lun7j4tc9esttWb0vEMamzT12W7ueuJw2QURaIRIVigZbM7qGSRYi6Rdqx8yq
5QSMLAV6q+1kCz2WGyRL4jkX/rYM0k4nf0O1BEQMdflKMr7CHEpZ9ujOWhJWX60T
8uf1glErRwHgqd7w2ZL4PIy7bEGb1nb4x1Dt/g5Y02nrZufc8nTqgnEv9QhMkOE3
zF3zbIIqTHsP4gLhT5x/BWRkxClUREda8ViZO9sjaMWgEHJA8kq+EHd8TDVZzDRt
oZ86PQunquhCuawdrH/fEw7QS1KriHZZHUGTyi73EuImFtqdVfDR5XxQ33YThdXF
JisET8whB/iPweeR4PwVqgXXqHOYzEk7NHmHd4D40KzQRRcu8lsUykVT+c3kwv6f
Y39cngZVEPHj++XYkj+IpNvT6dQSA6qXc1LTPsSswnPHyMfV+WnDxQUqaiv0ylYX
jr8AICSzekPPcj612vK1Ot1aPc8K37vXynkKOxb9Jyj1/aGi3C8S/tCKSlFs6+eo
OwciHUOMgf3g/mVjFyFTPBnv1hZQ77sUnN1uySBJnydtQn3BJVJw8AkxNqqmNv5x
n2WEqGAaQMu7bUDhUOtxak2k3A5G+knVLxGmvpk0RZw23cdFcptlzM7ND1gvfu1S
A7bJpcWgzMy5WgEhiGKd7oUaJpJWqFBJJ+CNHL5NCypvl9GQO6SM5lYgHABsxyGw
flxKY8igYKZEyEymwiyFHMQHyoQs65COxsn9svhjgLHprYU2P3gQrMue6dxO5a0K
wHYhaw0ZUC+C3yh3XO6HRRbWWM5QXeovCvEcJw6crXEysn8vKRHUNaGYlXhQDLxp
Qs8wvYtawAZbO7CHGGYhWJd5C0C/BZEper+vd05DWGmyGhsaezq4VgvlwEz5Ekhh
g8HyUWTSRO5wC0rI1xK6iCNQ1HHhO2t64VlwETYPQ0IzlqvPDEyH/vkfXVDeXGJ6
KkusEukg725V11YixTo4NlHAd2VcpgPHsdLW5HCpyzf7J+UuTGA0tNnWHYUwrXp2
vpGtV3XhHl7fkGJGsckfyYBvT7W/bi48cohOwBwJy0AW4N86Q9bSzahovAi170nl
zL+tWDGkQAcRvTWEsyLQDWqd0vwwLFsu8dZPFT8iniKp8xlqrVSoZ0JOUBT7p2eA
9Cy6GvbIR+GRMAWuaypsZiGspeFBKMslaDAFlOu+AH8N5XRueNQmBrJNJxsxFya4
p3WKjwOs1TF/DLLZicXePNq+7sQvstNUiU7Qau6fnFnyPyAKwahHg9cr/B+5Vw10
lDPwJn19fTEA4ChtKqmtyPuDMv84PywKxz7tD2FERWpEYCsJuGzwF5flAgkEd+ZL
wj1ReagzdHjs2tmi09zY7fN5WQYjZNmjlE8vwb+AVoalgVV71/RBxu7a2yUVvX9P
YbOpC03CgUvYwVm9F9oVVEfAjr4yjMDB4s6xvTaehQkq7cpaoda2luWUG4uZXGnb
kFj8lVoSE0wQqOUnMKDMTrDnf83pf7sNNHqJGn0ZZ1KRBtec9DmCOziLjb0WShW8
8/jHdwUyFktomSVmIPpQ8eeALb28kdPk1ds0SbRDHJr2UmgGKQ9kQQMBUgVMsNpp
08+oUttz2tXS2MCoyG4K57uz15TFoz+W0UI2CbQZYWh8y7NuxXC5DOkTc//0KHsw
NEXGqXoHg/BUqvvfuYSZM+EaHOhACECqzjwPY8jD6X+KG/assJIuGf5ZwNLg4KOO
3UgsSixuFowLg8O+QLNfZ+P/FdhLIa61OsrJMHbIe3XN5iRBXkqEtTqzO9f9XDik
5yDymH9rp6sBkp91Ztayg/ddL6bEd5pyoo5tNlB9aveec1ti3fGyXR7bDu/HCW3T
Y0jOZmKAxnaoh52BVmpvA5hJ6blZWj5oDCLlcvqjoxw8txov01Ota+UQrujc0mzU
cTC92luV+CEauRu9bfotEzLnN26ce45IHPm+ePZX71CaElUZUEuVi2ToKJo0447G
8JsdPJdEAxx0/X3mA0isqqioqAiAU5+oDEEm6l7kdRWpQkC7LUUem/fRrD1zAbJU
lUBlUctPRz5sj4et/94+pGDKEh3m4m40ZSgWCL6nq8+KrOIijxy00B0abZcYFWmD
d3exktkqwurElNoKe50C1+HU7hwGcNo7gNb5P3OpMzZbCbTQhDB7p3ZD82mi3LUG
DXeYWlpgVeONXGwqAecGaqIHR5PSOTLbtU02eZBR6obiSSUzVVM+vQBX1c/hZuIM
uES8ab8VJmCXvQ0l29CFZLysv6sVnvfgAlb0LEnGXUeLDZXFHSF5f+iYTKHUTk93
IZ7Kte2zU7C6kgaXD6ZmqzqFVOZ8MI8afvlSCkWko3rrN2ziwxuci0sofPoEuf3Z
TVrzdOJv+bv3TiNyfAShriCp81+UTx6nPHdpL1i1ZupTMYGmyZcOaqY5k+0Iijys
/EV/3Wxeqi3A/g/zS2EQp326ahmPVw4587YSKXbViYyMn8c4wwsJjC8Knivh5T56
GaYm88rExYux8rWvmPvFqXChLuTcMkSwGrqelg4FPpj71LIlGjxYHwwokLHCGncy
YiEYNM+wNCe3LaxwV64cvDGqbnDeBGKiyNj1mPNN7W1YCf5VbA41o0/44Q5MtkRs
mV8SBb46l27PZKu/aQ2VJHPJ4WWT8FpeXwSKRLD2CU/84vBmJLvSm3toweQVAfGR
p0LWRAKvhpX267oGxHCMhCS2dGa8Ts8/zRYZiTZMciHbnZqd0hpeeYvm+xxfpBuy
Dbt+CIRfnNYLLmqFadiROVjbhohqnuK9sPraHFpFyEaSnxE7tpBOCHuMw/rqLIXN
J59rqyjwQW/7rKCTYLmdp9Tm6cgkYIda6sx9yDF6WhBu1V3iTkEclZ2lj1fmjKqw
qvahW8EBHlUwSAScdxmskY6XFe8bHGybIgypFAaNWOPSsURE4G998er/bgqOYxdR
/Dv92HqS5NQ2RpzkQBzE5WvUO8Ejjs+GQUK954tiod937XKlg+md6QmlcLSvGRxI
y5a9G07tkxqzaJSTJJ+u80qXQvawj3fba9XTsslIIG88lDGSXt9xXu9+xZHrPRG6
27Zkfian0eMowqDs5Qcloo8UKIy0tFFH4CoGFukbeyq5Vif5odBZiE43qWICqq0c
3zcDLwrnTK/D3meMlc88N+gxt+G4PrzVs9el00s7qpkUyPaj3Jkqkkdbs/WcCHBV
RqGNSHjaN7HLLKm5sM5FECWkJVLE0IrQmp3zpy0ZbHWK/voRZZFv8q55NeuS8B5d
aKJubtsram4X1ZPA5dCohHQpQ8si0xqJe3ApS1jv6mS5J/YzOTdy1oTcexAX3HXN
r7vsYiY8e0yRN1swuNJ/kfNJgd39m2APDinxX4oLu56nL3pZbVNfDpUUdJ3kY9pK
65gyFpj63y6+Nrqhuv9JbX2JCauco5LtTSzFSrVI5+A6VgIyVFoBOsDyCcttEX1v
+4+QZl24zg/FS2YLTF6sDBvm57cJE5PF64I9loMJQL1hziuM3YNuYwfWAOu0mboI
m7ayd05n2cucJpQY1rNb7w0oe0KEhOGY9u5wn5gGPfQrJAbknamxiE+dqxs/pg+J
i9WG+oKD9AkHCKy73Sylou4uh0gjr4VM41SzT8oNvznakfWXmIo04fYlwtUrHu5c
yR9p0ZSW/WXGyx7DVGRW6gwufO558Rq22/B92csMC3mgNUQfWG6Q5VWZP2RGEOXs
/mQaFKthqfkTlO6X6Gv3Tlle61Wwdlo0sQnGGKwUv34W9f/dRvTRXPk3YKvdJJZp
/AaQXm3d1NdLRG+bqn7Pots43DcxcKvRpR0jR4lZZ9X1mLDZRmq9a+uzCwaNwgFh
+fFwIhNEw4rUrLGFwyVTxbmry6QVQ4YC0rNiUZyo+gceJLFAQCMejGdpnN9kfMBC
Q0Gcf1LdbCpfXqeV+XUN3zs5dSACsyNw3no9Q8nATr+irQBUKX3YtF53DG4YCuhl
Cx0Vt547v8739yyuFyBSYrm8AtotsL3AD3c2UHHZWno4ncQOCLbTjbc1hTw0EZIZ
yhmps8F5pifxSSS6gB+sqJ31PW9mLe+R8ynFyk86YsjYvtfCTX3W+AQB3PgtShXT
MiP9HCC24IbC2Bz+wcMdBCzpIgLHSrKTBEG/9ovg558ZaexUfB8GqJYuxMg88h6n
Xk7dZKcQP1539BIANCCAoimnbLtS1QpIKatLWSrH9dmZeyu5oN20t2IsWZAzyrT7
o+3n5eQ3PIOJY7iT8e4uM0TTHLOeNVq9NoCd2mQ/GCc21zxeZrrGlV6KH6ZRe6O4
JO2pPiCtoCnPzNG4k81tS7tdtT2HjG+C6IPdwLoBUL3ExikdofsAyA01rwrAsP8g
Bz09k2sDnxccc7TeMSCCBBpk41Yr2/1FidU/U4K5Wpvdlt/59ksilVg/IyGyKRfm
leEIpSJ4I8HGFj82kgzdJPN4MkkIXXbEgaXNpzfOTXwnx1ZBPVeQxpBOlo/HYea0
rJmGPN6n6oGK5grzbvoOfLISLqCZ44D/P8ZzqCDlrrKs0FoRe0EkuP9X6ZBwaqf8
nVhtgYT135g9zYto+YrJ+p3IKGeRuRKrvRymFqr6E8CrW1qQr5SZfGHRsUpP462F
/6hMITfCkJfYx+/cjAMgVa1q3Y7SSJi0vZC5pe7NgFrJmX+b5/n0+pOEf3HSxPYC
JoNUOxMxKBAUz1CbqB5pS3dSONdsxt1XnoPB0BOADIiBiCtJefZQzkpO7Gwqxj2c
u4x+9fioN085JHjuNPhLVtQrNKBX1eCprGEB0yshOv7yagU0zG2zcfsf2VR+ELJ/
vkHvwvZ7mv2nv27/zU6mjO28zZjjaUJFULkyUOjWcpH173bWXkyG9A9bqRJigb7p
uFOK1+ocp3ptxgCMlTyiQwqw/5lImyd/hYLhakwCxb5dzmxjmQCfLwix0x04u2M+
+NI3mu7R2/lJGPB5WQ8NVWAOAxECzkCVXYP260oY/Sxucx9eW4dJvwgnO5ycGhCN
JQ/hRpDi2EaHoEBeJ/K7zpPkdc5Bhu6OINXvBBUW2Z3AYEqX/dnPoxomjb4z6tLD
t7YxeSvMc0wtMAVS75qvreDcqZs1mTMF6OschBcBSG98AcmnHdHS5oHmbpvEyXFR
wHB4mhh/KY3VwzB3ZQ60UnIVMMj12zIzrEOlxtjmw7PIMzC8jAC3butzSmUw8yst
8hzO3Nd3tN8ePoYUK4UKnsnmSye5ndPue87IS8Ky9hj2VFF+vrRRSwxkFWukW7ci
9r6sG8PvGsBaMjGReMYD0UCvJ1jMylOVoknFSMyYpPgeayCj49zWgmrQXgKnBodU
QmmWTnSPYLuezfIL7tfkb705XYlRq0SPK+pBZAdw6BZ0tPGvJTjeB2ac5rK+i03/
mG7hEeA63nfJZopBRvKeLTIFWse8kGR/MG87qGHAzvRJe/m9f10u3aRLA41d/aod
xz/n74d2kp610h37kxaXOhEJ11rS3L0jrvpA3/+wQaGhTZ+yf8fh1tTJBRpHhTlT
s3zcSQOoj16x4B4BqMLO95G63vjDfmonOWeWvJ5bEDIp6mdV299//ZTz0uPp/vjl
PuQ/4nK1IOnC5PEFArz6qGcYfZCC8u6kaexPx67q+yiQd5mgXTGx4vfbRtuUq1qo
L7qkjIJKAP9rINX4HODAti0xnlxWqoU4ugMX+Cepyt7bQj53WwjZiELxDpNApEwt
oOrgIH9LFm6xJwnExw//3TNEx5bHq840lCknoqFXn1eZshOJMTMtd+sXHXFeH65q
BQ+NQkOtxgdp4shlryy232kF4VA9Xu1IPqtLrTfbJHg8dGJLunxSmNeZWtZ3aT6F
3DrleEEYADmYBGEQvN7RVM/ZEi32I0THFNB4HMe38ZF1a2ho+I4Z9Iwulmh0ZDR4
TsUp/aNa4zbyw7znlRoh4Tjog6Sayo5VCj2rUNBgQK3VPhdr7rLVQjsccLaDjhs0
+ME3ISn9i1BPNWmn1m0XpbzQJTpiTSRiQqzbSXQ7elGpUgPct1Y/gIMVJVVCd90A
w3Obm9c6kqEUB7EXZiHU5tSq1xp+GCcYZnpkeMJzTan4qJpOWLmtf0FZCELK000L
/Eck0i/X2pzuvmo/v5nXILKmpocWmaGitV8zZZoV+gR7fQ59ldAATFE6nQr1teHS
EvFNx3AHiHZd1ArESEqOS5VvLVA+z8Kor5dio57ScZ41V6OVFgk/P9qnRfCyJGWX
6HxXFAUbwhlr2HLLIR1X81lhfJ5XjEzj3pLU0lRUond06W613CthiSsORzjTL8tD
HIw5cW1LDHmw5UC8ryByIzmQBXIZ/qMiJ1+RWiiScd4wabkTHyKLRBusWxUG0RG2
KGLXisqw09HPWDB2xm4w/jQPN9rSbhvv4DTKimawCsSjAviO+DSqcnHaXseL5Cu6
COzLDMTLs5wxjUQ84GT42UOTDfLov60NrBN7e1UvjeNKJtzCAlTl/sstq8Vo0YUZ
LmZnY9Mapfq3SwTNrheAuOeRVP6WCLX9Ib3TH6zHNQawdM2mFgnt1riPWMMMy9OF
m+d5iFEDFu96YVNKU897PnZZgoR3CnztG+CeJW46VzP4iQQt8a8QY+hcfA65XZtb
Re69MvjP4808oW/Ig0lXPjvhf4ixxa8NWPiY2ZSNrBUwNoo/7sOdaqP5keppAAtk
AxNLR+gjXM3kPmSWz+NkLJND8SLzc+eeAkZoWRcaqagybbt+Qacu+OHXgoEtUCOj
4eMLBBGUwMs2EmjQMYG6AEwDOvJvFZyY+h8QSiAUFAJ8A/gRfNuUvtWP7JPpS4on
kOcOLlO3jRDj0gAz1APeX/MrDfgk9IDUKBUmkLtajA4z2dVnFoxPm5Na6TI78xWl
AEoBCCrpOo0Chii9iijVJrctNKUpTaLC2hvfeelYR5IpsXp9oErsbOHTCAgWJxoL
lbncJSD00lIQknxnmSa+lK58U4tcD4KDQcrgRw9FjGy5mcKT02S6owUTp3Qby173
pv7ozsc7XVSBJA7DdiELCXrpMO4KTNf5dUn9Z11DYP60CwaGRy49tpkQUw0EuK4o
LpkD6fN1qVtHzFHlkxco7gWC9aFXvJfGfilVMB3lRNgA1FT7UmGI5c0rppV37Zvj
ULfl1SQCwrVJeumVbtizgTEdzP3tDOajtpaxDex7iQyiUHsrbucp/saR4QsQeRc+
nE5BB55KI/4SQ+3bZURzFYU6Ptm6O5DuNIZJbl1ePddoRL4R2IARosptN8NCJlB3
HlRLBhqqjdWrYNzPY77446Xh2N+L/sy+FlExpqud6NtkfmyQjvVF8KTT1LeP4vIt
kKT2S5Cu2eMX+dTbifBoa1hyvTq2k/+Dm3DiU2oLiSSW8oPgtBPB9++2Vf4T2J/C
YcVPF9w8RRTYzo7q7QetnRJMlotT6NHH3ta/8oGEoXOJhIoAJzaGkg5PYSCYV+9v
mORpBfQPzOeGxwiKQBW63iocawyRSY0RGQH2YT1APIaeGG6a+n+TYfHL62Naa6an
3V5WwAPfuM72xQ2GJOxgw59/yi2LT2SDk7Ie4OS+e4useVHjYbbvDmoKCVXoW7fn
CVOBxtLAu6aHSryEH3LjO/QIWmW3gERCXQiEcDVck5HSyFC/HfbxLUqDrSX/zyw2
sBz+ODpQfaTa66PnGUkW631FwtqZ8yC79FogWZyr7uz69iGU+cAAnPys535pTuov
PFH6SXoDOUkq5vYcT52TEQvtAcb1L3zspVMyybKNuTgh746EZaKNgUskz93yz/3o
bU7AGd4obEJzJ+YHa6VCvlqG70ushVFMj/Fx9QbG3vXuB2rUvrxeQrBj8BxoIHKf
DZ4usYgrK3kIZLvgOMt/a91yMp/XA6oAz2vYIntzZ+6SUTaeKbCiAVKc55vVGgwr
JMF4Wi/u1CPWHGy+2ed0W8iKb4X3LWPXriRorOm71KnC9+X4MzbYHZ4FFp8MSeGp
jzU5qHyYsTbfVhNpQFSaKE6kB2GhDNA6Uy6wl2YS5XiqHM1fONDMGWcOQ5VsxOzi
MwILc+3ITpB3cCW6qLDqKKaDQHO1lGCFZruqxBunrVQrlpiZryW/SaDD+bnN8RZJ
PNCwGNg7qeXjO7RUOrcm3VcePll4/hadc6vU8cOitHu04zmz3WTpQNnQCRRj775a
0CMDQ0QMW5c33HZOCnmjZNP39Jq9WkwwPzTYyacJ68uzp+ovEqY7XBYrIO5SbNzy
eN/19nGorSAcsznFysjh49srfShQSs5y3VV8OTNXxjwotObKrXQVi1kK3lh9m0X1
PxReF6u6PGooBc6r9PgiCckCBKpA9Fjw5S8qPdbdjAfwFcw9/ikr0eccsfFYxE6h
19WxBHZW5+qQT3W8cpYwDA77u06xAeSN7Y62KXASfxPoOnOol11UJ5q0LDfIp6ht
AZEAxFpxnHSqsIaC0+CXXzcuFZPJKqpB3vbbtXmFl+XV7olBUZjkPd/K9y8ANANb
LWVweweTXPzNEP4inZ6SLq7gF0G1xZoCdG3xSbrNC19jp5NEsrqFRs9p6shPpTwN
2kyGx4uZ8lkzk2NY01ykpEFx0vC9GZ5cxaFHCrdBDD79fiyfvyC8Iilm836ZtG/3
NeEapX9F9WMKrhIPe8dwtgCrFBFh2ftrH2TcQXvwgnJrb7cVrRk91dwC1ZpQgV6A
LGnYrXOqG/TSTNHzT98g79VxXE6ozCWzrAGx2yDkDLrJJqn8FGBy+u5tmM4mnMgu
/gcc1F5TTaqpWffofHT3+lKb0Un3JHHbf6HS+zDzXg6bBdsDONFv7ErkqmY5ziWg
66q/WU+F0oscKXxQNANzycGkiRR1WMUy7FTARWNii3eWRCMJmTYPLNIGXvJP0q0s
O15M65vmq7oQC85yv3PCI4ZKrvU33xsgUdPGxhavCNB9VNlt1Uk1ZOc8SmuEdq5u
aFeDvCThvRGZnEzD9H2Av39kB9PD+eeG8r2hd5CWYw+ajGWWRC7engxWfwUEzpT8
CdrNICYrIAJ/+AH2VRcIdvzk+2XQhKgbw1F+FYlXBAXgbO4udLkZiXc2Ev1YjOBR
eNsnMvaszRVmLEDHwB1EDcY+nj0245EpVr7EcoYrLhJ3dWQiCIAD2ozSZ9eTsiqS
bgKhyynvw+9IdeqO3bYyioS54gkE9dGuhA1PvyheWScLPNRyneFMHXgyCFMDT+vQ
ixWJX6JV+hRWTNBMAJsVOmEBW8eRQfm8B/Cb6mSK/yByAykx1BHEikbbeW6mGiVs
MxrNM1zZ6xC02fk4ABLSPI+num/+zQKDeb5iSuv/M5olMRoy79LS5rnSrfJuoizH
iT6iL9ORUia9VW4ewoefQv15KAxvb05c7CwcLeynUnYRwAdsoxD4RZHJF3rK514F
JdnqXzgjjXt/hklVJqX/pbQWrLK/5/Pa0Jfw3yjVNjv6zNOdW51AVwR+gv+4rr0k
uqVpKGBIJ3Oo5IX6JhX2sHxJQfHz36wpWyp41mZSegBkW9PkZw2ZfA1uvzgUlIm8
+Drs1k9IT1KUqTM3NXfOkI4Wmt9dV53OOLxY2JDlUig0LhMNDcntyC14FqGlspwp
EWfMzSz1nOiTvsTOauJp4WpDLXSSk1ixmUs7zYOTjda3bCSP2THk/HdFtG4cjQX8
5v1qkM95FWCQsC3ZFZxOjYgUVclKYdO2MSvFbWEr6jE/06O4ThJ3mZKLsbnHnHKQ
cIeWfurVnriFDEoK+5TphJn57Gs3C9xJ/W8hkESEfPxMi4nYMKqSMJtC9kgLUF6A
WGXVsIEQNP0CXDpyi52yO0hYmXW/iqUlvfGK1Hk05lsCbI0GeEDsm+QKqghnJt04
LhpSlcuynXi93aKGLIXoGeiS5X/AMMxmVQdC+8ZlaU9JVAoqQALdKMYs3AjELiA5
urt0TybEaj/h5Kum18ggSQhMnyVSgXHiwyZiXyZB6setdrjB6+FHcrETAMn9P1sL
Xb/VJWgHmV/ISqo1Ar0ctvgCRjP9rKWlRtT+x2PKRysvWXlgQ73YMhsrkVByqIs9
u9gR/uKaTVmSo0r0b6zXWLbIAEawJ/H47DzHpE7EvciYRvXePYq0TkQ4QedMP77Z
Pt2V4GuVrJPKtUcXFzjmuNGXu3rgEWnf5jimHDNMOSUEItkVmdTLEQYQM2SBTMQZ
jL/rPNguX9Yz0IcRpr2in3NdP4MI76yfdE9GTPm6N6ka/NtiifjWGFQXNp09vxkS
CKXncEQErh/rdYGsXKs1x5W98z+aLu2xROv7cXU9mLRXl3G0qqkyRJMFG2w8L4He
2u7zDmJHFyz/ziaCHraSNFh3WNu63PRG1/whPzZ5PNLrzUU1lQ58FVGe7unKdrd7
cosGNBrm2zaOUPEUIBAn0FVtXWi9Mhm0JWu60kiCW1DZ0VjKAljRcLQKsZ3FiXAx
K8hfFF9x00TgFJZY4IW8jfgqa/q457gFf/+D4eQ5Cxs7ps70+lvLNpTyqwMzQtG3
lOJxIl3HfArt0Y+3b2SrcSZt5j9Z/CkqYGkJinz1pdWWI9blmuzeOxAUHh+z04Dn
B3SXzevA2euvaiUIWQnzq+EciUbnz454fVykoWtun/RqL7TnGWO6B6hR5zMs2ZyX
2T903j/0Pjjx+XTKLt90QjB7xDUPqy89LSXGxCCPjbHUr+A25H6aEbWq1Mci3MM5
54ofzk5V28ZLR6xI1bJtevL8Sd+f9mabTCTBL1xarhCeU8pZEYMrYQLhAb6nOj5J
4OD1N8p8g2qHFO+gs97fDVpyaumg0viuKoj/A4UzcmExnK46wwUGMXD+tUCn9VZC
xM/3NvygHrSEkepknN2VjpW98lUG1uRivVPSkM4Eemldx3ZiS6jggpsPoKVv6kGa
OJnhmD3fwJtzifFSJR16TFH308DCaq9tSvPdr9EX48mMq/kdYglMYY1TuUzMRTkJ
Hy7vULtLQWSav9QMKYHT+RxvVWfUopdviUHqGANnAUIZ7VhBH7qNQtDt4aEGpAJM
uQXMTLBo9jj2JePfVdujpCZZuHj4fLQBgDj9nPgt01BgY47FMkZWI9QpER+0B3MN
CtnJTLHUv2AzfaUOwyj7PRk7lkIXT8yX3Gxs7SThvJrOC4QVsEhjb5Jz671Lz8X3
Kf0N7z2jVgI6RnQ2ONtzlaIT7M4OjhTBxaCVKPzMCTGe3iTKlqWuce/Ydy2bmfHf
SjegY4eFBJ+807a7J39KJXwNELJsiI9bL4997rIp3tiyEUQtUboBxlDnrMeDs+Ur
UvmcK76jWOmNVqJgCDYawSsL3oc3w5CooohlLmTc86FsR8wWX7TGgvoNivWGv+A0
t/oRdZj3z+0+Odb+VpJkxkBe4qnRLqJe54VB+zHLsKbrxZDfnWWb2HIp4j6E73vD
CTrz2RwpuwabXJCRcj/GX/TK9jrXF3f7uM6ITK8EYTlS0F5VUff01ciRyXfiRacJ
U8GeX9yGtsEPulYXdYRxG71lD7thiZcf6zQy45s5U+NZGNwvvP/c4hAF5V20gxIB
isvtV6x5eoB2bBSrihWOsqBuDKxiDCZZHMwipbO8p63sZCQYxIX0bgmxBuByDjtG
u7mX09lrAQLTGmO8QLaF0xCfT1tbgIvobzuh+ucweN15o+qbYAXSlT2ABhR9/lD5
VTFpk5EH1Bv0BFDhqvDldougnV5KkgACD7HUwtSU2LP3tU7m0eZNHK2LouQRmey9
fC9Wqas/3vqmOfmwR/ofQcg9xTgU5gdq0X8F9CNU0t7ZCSK8KwxLJg/Ysg40xYi9
s0D7MHTnlisrvGfqkoVav6P1/vCAVbYYhLLvLBxV93HOgb5jXirqIti/IE8+wh2f
NomeyhZcujLjynWobC2PAoiOHJEDwicbT+FPaao5kXDglCsbM4Aq9n0A2vKto2la
9/b9F4FnzlTEryq99Yo48U4jgR3TG6fxw8CT4mmGNOp262YRVZn3q6fVGWhoJFgH
XkOPIOtUECGAhm/vFpqgfZsX2AxElKNEbNesypvhcIsdCot7JzKRaUBsnM2w6m1x
+Ken434FpbX6BIt9Va1p89OXP8jaODpBhUA8beXFUidgQfxihYc04x/B31aUuDqt
77Zio53yt4r5aTu00vJNQrNTTv3LKHRsXa9/zOY67lND7NoPrOwnSOEtls7kshBA
RsFMWE+9NFjSFF0jX31J2Lb0YeVNSVvqRzPrAQirD0zR0fOYNuogHe+skALtD/ei
zW1X6sr+vlcDWCVn0utom3YvoIjKoZwHhwlXBsD4TqzGmDa6MGVr2ANy3I1c+NWl
CqVckfeWSnspv6TTe3kR3UNffVO3aiT/NrawqTqz3zB0/nk3F2UpQLrFm56/bdUR
JKBG+onVBEqLZL9Uu5EyAMtANPw0rYyc630Nr6RPgzp9enFD2CyjnnypkRHeQcKT
gGr6l6b2LrnLNbrEruot4nyMudX2Id7VOfVWalxA1mvAaVCL4BwC3ugxiHJcczYQ
Io+9iXMKN/uYezz+lmQ8NTkmM9uxJ2PV98MjpGAYQ/EeBvlgxndAhyaDkaDaHNHA
oiGG0eI4TzHTfOzTOn1Y+hJquioIScpdPRxidG6RpuAOUuUUI6hOsJOQjE7eon8h
qTxiW9bCiBHl4tu/NFYIyKI/oa9ta+caZCjpLG0IAxI+qSRZn3xdnoapBB3AjyzJ
bqvTb9OQ4dsD2rmuYpDSL3NutuPckeEDp4xxyVe/T9o2x3nQAGCxU+9OLgVE2RYy
9q+u5W0PIy8iBCQPdMrwFh1ccDHSebgEj+afElXYBo4Dy10dGxY4mocRCbfCI6gv
JxAiMM5lCmSapICJPgl6u/I6mamolvpjSgoO2GNURx3SCaUkMQG4/+VA+HxHlAT5
dR33Rk+QypyMayoGqAvO5/hC3VKNEZxvyxR0KnIIGqcnvPg56Ao3E7Nz/at17EGB
zCRCz3CLzxkdIOodWRlZYdzHKg9uQcYDM+uTPYU7j+M5Ih6T7DOYqdnpYf+ZvnYJ
AQL0Uj72ocpDFnmhaRHlK/2WHB2dYZwiV8q9Cu/A8EJtxHsMaWxxxSQ6fE7JM1iB
kgxn6FyPlM6KaSlml+n0NP9lOJiQxOjj2nBjty5/yPzQDUV6l8JvHL6kj+K5tYUw
t65PzKLFa8b2unmfXiOG+rX7YhrryW3l0tXw677d7w3p6OqJ0S8RRulaZw7Dc7rE
2VD5QO0aSW3xMmsEV9z2gMQ8U9+3zdhdh9/seGMrqAGuqfdFziBx09amaN4jCDCR
ImvOBG8ZjuKAIavjNM1ckonUBSwD9AMKW10psspvTqMdVi/eSrhuVNEqu789rmDq
nN/qyCHICtDBCdKzSHphxHiL7hq4jI0qxGX7zqdSC/dfz/H5w5tBV7ahVjz/BA6V
7YKp3DM3TndDea78W+G4lXUgRX6cYpyIqrat4HovRxnqil36FFdsdb6T3GlYjDUg
FyjdxZuFY76utIAuN/ugDIv75LIqmUm4ZNjvKl3uHE0HTgI2EdQ/JfkeahASS1nj
WlzB8MB1vv49+OxUWV/sg9IJ+EtCvldtk2qbL8OQ1anVvmeaTlRgb1qzmOztIF7a
TJoocxc6RKWX9hZaUXbvbGKOMMDnu/6MKoopc3T1QcnVSORTrQBG6Evi0w4WkjLB
Ce7hzx+TNuVan5976tTZKuZczDLHzKaOgJzeOT6iyyHiG0d9NGsA48JeMIYpch1T
FVilKmgbZQGz1Q2iOYukCk4uHof61TDzoNe0yqRldwHqN4Lzl2/J0RQQkMgbkIz2
tO48vGqlpREbum4j3fXHVQaz8zbX07mD50r5HmhlIs366d76cpWfWaurz0iEPGDN
lkkVqHWIJhCBMmTjen5zanEHd28RGhj1e90tyKsSLm+DqYngY3lzqeqIekMCoSXu
EOGwHLEPyd/37OVTJk5yVHZ7DsyKX2ZpIpdJGqsWfSUPcl1xQZYiiYbTzO+4Ho8F
n1T/Cx+628NdVW60Yi4VEyI6dTotzUXJ++Hv/Z3SOKJqlnb+DPRa66OCj8SdK1xj
FCZYp3ufT5w/Mlw/7Ou8cWriqKfcM7Vmz2RpjqqSLGXMhbgaMna5NXx0RVKO8Vzr
hKWbPN0Nb43tLgCiTxCeU03kFsD52A6vYpQf+UbF5Si8RX5XPUcxLo3e4IjoT6sX
0dEwt+C+7M11heCoplK4H7SRxwW4hstd8dS/6ETu1BgrbDBRs1TrM8kvaU9Su++s
nSCAqLsOF3hITL29O2Rjq2TVNpyjv2RN/Zx8NvNZnBHiMt0WC4+MeFf/b3CSBTTy
6zBsJ8+DVrpv01DSRvxQUDgQarCPH4T/Mej+ZMO5VIyJtDue6E8UKz8g1q0GBtJe
0wEZof2hlriuMOAF1KilyU9Q7RNlPK1ooTeZRu2vgU66hFN2TAqxhw5EbC+s8bsB
+cg+gMb6B6d3CTNP304JMIQNw53r3JodjWCCSLIMNlwwvJVjcIvg4wKYy/hvimjs
MXJEtW8bGUG5S/3Lueo/nMkceRPds4aTsHXoeDdIMnmNLbs3igr+V+8U6fo/SNTQ
a5QomV+pd8R3Bwe4NnaCqKVa+l/0daM1TQaCuUllmlLhxL2qwfUyMQN9W8x2fdMA
3yAyi+lxXqlgQ91qngiQy7x+v+yLP7WDatQYmuwI5FscamZZpG+QH9iWJBFUaMVc
HJJ1LFe8Hg2aI+o5wzwBPoqso2tpJT+FUYxqUDXfrPaZO/ft4IQbjgwi2BUSxx1s
m5WQSC8Py/JvLHzBMVwIRbOUeqn9d1iz52P8NWks+bsB58Kr2YcQJSk1fQ033XfM
k+49QFn+l8UqRIQ8BtCtrku/yWasDZPWpsTIZJyCi1Ymn3V4rJ9P5n/9tayK5mmt
Eh8H9bdgBWlul7wnmaoSSMr/+liESPpCQH0dAwfJVFVaCnaKiTiKh/HAFRLqJRx9
HAWxCxbzNRf3AMpHSH+o/hrnndZ38IJf5yBbd1WfE9MONC6FAqUA6il31UUakc5l
ELfrd47wLtDpkmmRAdsOnOHdJsij48SR47938mWX8O7ithVi9LYFKGJ6yiPcN6Xp
Dzl8U1kKGuk53tbxilgoPeepYoWS7x/+aDGKg4UURfHCAK2rq4AgsBlRqxalFGEy
Tn2n0G9dBPVH1wkTG3Aa+v5/SxV6OQkddiltMVYyeZrmTO3rZ+BVXZ2BFlF5IY8Z
Wb1DDR5rv9uZgUXUj3dpIDMCC5eP+cV8IlMBXkX1uOrEY25M2Otsod5xXpo6ixmS
lcWk9AQdTvcyTOdgAiUmmL+J9622nxQbKnKQbXc339LsflgGOc5MnNQ8rnInXB69
HMKzgJtjwo4CVJAl0wwggpARQbQOpUSi1SG6YQDzYH4IbwgPWq/q/at3wAr6rN+B
ZH9jc6DLYYRb5xho/o8hh2VBAMGRypBpUaqYUreuT9vJQXm2Ut8YYH0LYvD890Pt
XtJPUNSRMS38Zwwe72Bmh7Ye4kxoEBDWg2Zb660f1A15dfhbU5CKEWVHzWvewqOk
6i3Qe+4hdYlDdhKYo+RHC7XBoHyvO7tY4O19yhLACUexmb7/8Tc5uEKMWagDWtcb
jJKQcubeHfukbSYgNBHBv8acDxwR3nZpVneoIWNtPVHStrOA1oQuXq8JctxjjClf
B/TRuMOUOCRQFtuJK6invDLOFl3T/esP1I4d6BS1VSpmq5rmdBL5wOS027bfSr3+
YKT0TzL/BxOrwS60py/UekbFPdypbYZgDAuHxgea8zXGCnMRf1YIpgEGPVYvqrrB
CV8bPCJvR7465qhgLaULjOCuN1yc0wijaXFjhG6wQUjM9Df5Myf2T76QyE+Tn38b
Oa1sABpT2lAJ84vj1WzoGsyvf02hQ4halVCCrPMJyYwqbF60Yr3e3cQYnazfkx1m
JEHrLXQmUoyvr2kIWpZaoaCArUwgSsVo4yJDYKW/36VZYL59b7YLOAE8PZAlVEHe
rs+MQzZ/94YGJUsAZwIHvw1MBtnI3K0LkWVy+KeNJZ0d61C6ttHcsYgXwVSA0HJq
ufPELJhTGXKFK2a/Hgstu2fhbp94fH1zFGUqfUE+SAEdzd/DznKG+3KRWMR9vpXH
uadq5MzOzqVg4GVn5EzSU+yTGUnVIOAx2u3YHQa2J83Pb6nAFq6aQofCj4yJBHfW
q8lZ9JGhoiGmk+qzwBcj/0+H1d49Mvv8TX/pbvC2dw/809Y4IZUGqa8FyeWjs09z
zxAOuRSThRkoJ6fnXLB3DT9b3Pa+b2iK48srL2SF0nF13LH6RemZU4kCyaYosy6d
tv41zG2I4Z8oks7++hk31v0c3N9hXnR2Nd+eMyIcTF2OCgcPwgO3Gp84MKg58ge5
mGy6RUd3XsniJrwGXu9efqvYzgHAjiXa3+xd4IzQyASY6Wz9sYtpLkYreyxnc81/
/ZQmdPJ9b+35qFRcCmvp+3HyswygdJIiaHYaGmPPTGY8sZuGDYCMSLhlWvPjJeGI
9QFMUo1KsSptPEODtVa6LoavH2WJKgkpTcSw/pIOS+1VB19h94HxZR+0XHjndKY0
Q4vHoH3c/h5mPSTbONg52RNe0aUAOEyYNp5X201xuu7C/ALu2TspsTbIYtetFiIN
SWPfd0mejuNB+ZKjIktp8RgASolUx/j96ZupNwcHJUAg861DDR16ppegihX13goz
+N5SgnBZ18eXUUuV2983pwyXdrTSLiJNPT3ARSU+AbBNe6ymLfKsw14BK7xyDJif
0u8Rt+Jp2oXtqAj0wf5xyyU+JOG+WAG8qN2eBPBFjVYjLUsH28S41g2jWm849sYu
kL5dQvCZlsPZf75+TucUPadibfixKATLd40LqRL5kmBthV9DIgGmvT6OTFORU1oV
uSn0TTSQ9tF+N1WtEpKfqR8Nk2PiPdAncVn+czLrEdW8JctPMvyHFYu0QJRBloW2
Zz6zqzElUwFfiHxnfRKM45cQh5sTIpPg8afJrDMKAvTquBpmShXLHSqkJ0A+AeqM
ZFfFcSsaS3kEUgYsohfc8W75Q0wDIAaO/mPGsKZQBE1dijcGNUbDwPrV7syRLcMH
CmL0qTTzuiOecRqeC3wfhrYUgsH670AnQKjwqZbxt3f9D5/r1h8A9gCWRzEuR84g
d5Pu81AVkvDlLH6Ku1i8WVTX2qocukUs34n2iMIvkIiIIJrCo8Nfe71GWXPnjJsk
io6JJX8EUVe4rkywgFleF6xXiN8Uz4zH3WVJbyO8cVZrJWWGhzz+mwy0PADlA+cJ
Sy6AfyUCUNGlaVTzrgZ5qtQ3IBowQMWMibtGomZgAVzTa//WpM2izpdEki135shv
dBGjIxdOfz2fRfVXcKjLLjvwpnjSNIzFXnNuMtlSY+ZSkzLoM/GmkMEa4+sFeex4
4/3h8cwExMJIWVGPeKCzdZud3PLzQh4lQiRhxIuEfA+cIexauKxgShIb/cLudtI2
Vh1RPEJDt/oTe2yM+Vuu1q4vITpaxABZ+bL5K66f7SZyuIzpSfuhLzkP2faXcarK
36QsoHbvdVZA6xxJJ13C4w2GvDWxHlbl0wBNouXzyDIQez6s39sP6S1mkW9D56Sc
Irj6rU5huhaaIUwyCbM+b8V8wXeIIZdxENjATDytAGrJ2y8xZTFtw6CAjNrvgOSu
dZvfufZ7PajPRKnyMh52hefmc+XcyeqhJ4qPcE+0+gvr5nfuwrADOKfLm9saLKt+
uyjNQOz3wR3md+FgL+0xNiF3M6LOyoSUAh8DMLsvZsg9d7Dk+aj5B+FrUS46FsHh
TAqW9KdXR/KmUAiXlXXdF4naQ7eg3l5phAL3mlXhQSGZyY8wRDSNgtjfOwoQ0xQo
6d+sNXCyRIQhMl43Bd6tvndP8oNmtRBi46LBGUJ3qml8I9dS/sMWsW+68Zojxj2r
c65kkaf5jglU3pXvYOURSR/FbWw3HeWmE8p4Axd4Mu0DrH7XysjEDNucNPvk5sbx
QIfz4UO8CrBTmcyowjyYpJZqwMaMW/FoiUtzTkt/MXU4D0rZ/BZ+DtLkqH7gb4po
ichb8Oj3IoPiIl+Au6p1IJBo9iQ8+9aS207ImhbZ+rDmq0Ma+tgDourBx0kBglQK
bhGiqIfdOsI1BOdYkdSMk9B7xPdKr5ZnFx2VDpubRc8NaCI4KMNQu7h9i73V07cy
QoxhygvqCA+7l9Kp1NWM18Z+uGe1Vw3F2Y8OrdZ9Bpaj4IN2jRKu6D5av+JGCF7v
K1F7UnumNA+uf6WkaAhiRQIgansRcHzWw/Qsv+nuW+LI8xe5n8auD/nXJh7SR7RV
gUNspSpKVz2fEXFpIr2igV4avfiR+4iS6wWAAjWX43CNkYhXTooZewKnOkdGJBAT
+YEea4oEFRvRTAgJKHmoDB11KMzMsMnzhE0on7QL+3T0w1eSUzSDS7zueYE6Q2S3
HPsA1GGFSqeC0jL0BuVmdyoaAu4XIJqzri69C5RpQ4K52BP+CUSYUZl3TqPDUV4G
uv7l6s8KlhItZciohV2jyaFsGjBR1Kl8t5DbM9b5lkkxBOUGsqqx+KBtqz0kXUqh
hgtCbgObtS5shRrRTPoyi3yqMzLROE2HGM3kjZT8CVavJvjrCR8OkCML8dlJBEi9
Llz4cfFLY1saf/nbuHzNKg0XNdF3jbtn9eKLI8sdpU1BFDHY2x3q8t1OsRWlcRuJ
xxwh39y/eD6JxqljDEz5c3f+iqSqQc6kEC+6+wXcSXLyCFU0CAIFGUVtULLGCuac
RWZdr3t1/imShWLL7mSrCbGQHg411upXQG33mvUaaEmx+hA7B/0AjAB77wg0tCng
c/4K7VLCps+xDpi8gq1rhfE1yyTJaGZ8G22sBxWz5V8ef8f1+DVH1ojJiIx8KBof
wMUxjV7DYss6aNart9jIzIG2aShQAOXrT0yvXv/mQKLJEcJqfc2of56MYbKD+v37
TXL0dg85iv92+/WcXX1NiwQj9mEN6V9FLmvktbo2i7WrrttzfYgR6qQMfs+peLV/
pYKyGjkIv6PjmZf0Q54hjfVsF+FXUoe9ouXwiY5oAqNNKuf6F4lEgAsmL3X4bB9s
t0xjpuL3vYPANfF8RODOC1KH5CoK539riHcJ8EN/VxxduI2fO5oT+1yYkeA6it8l
bcbHw3xWUK0c7v1F7fk4+WqGBltRZrdarhX4kniIYy5UGbc2vmnCOniX1KaVd8P3
WAx79qnzkroluNYbxeeOhF80Yl9Mjx+ofJoGlXCBcgruJ/XxIB5kMw/5HoXxyhIw
TeIk/MRt5T67xKntehcl/iOoDdfbzpNndMUz6z+YfL4ckw/vuq97C760ivBn90UI
uyNPavSpElM2NUb0sEcwsTYH/ie9b5aVtuIBS1cmx9jB0lC4k9e6syfB1z4MlB7m
zEokVMhin/bqHXrYaXt13htTmMN6gj2NCT3u0zh/WRan7fvLyKWrVhLfLMoFWqsm
AMGQoZcL426j9/6RIFM+xqpftRBG9z6Qwm+T/5yiuItoocInqag8I24pY0B5k+rv
9IiwKfvtWZ2RJIh/TawkJ//bJmZC/AG9pUlpzkV95HhcFNOG4pMNAsjQv4hsd6Mj
kVfmwPQlX1vkkJtz0vnczvm/Eb1e3NIw6EEleT8neY77dTdOK4nFV7ckaJVxMwaP
ECzMycMAB9V3AbzjeeDf+bi0B8shm1UqHYMOfCzSDelD1nxl+bjfZmJj654Ihl20
ncEd8FKgZa/uXBRRck/RvWx9gUpNCiOWMU/EHxFqLk3pn1mJnWY+zLYIYuJutdYk
Ev9G+2INMXCxMiqqq5jp/DzxW4a9Vqz+qjd7jNDct5+eMuseHr86OUAR50DaxoOU
2SC/l+LpRfzQY4l+jZa8PNWYi80VSIKZz3USeEcQSq8OARzhUqC4KlmwtuHkOv92
HD9N6GpMp1zt+qTnjx/Y+guPC/B1sFvmDk1l7h9+2xDNqE/nHqrynRVUdbvg34aZ
7S5XmezEw6DQvu2f+GUEVdvGFDg8toXGExT+dUCad97f3YTewX+fxbAPeVywDYEs
GNUW5a5wZOeWxAppldlYQN7KaQSZiAtxs7MijDd+dZaetBETO0HEKE8YRW2Q1PFh
yykZb9ZNzWMdLQTLKPTRG0XRf6g/mcocOeQbCyeih58Fu9MB2Wm8+2RzC7gzmseh
vkIL/v5kYFjSyVThlAu7Qxs8pQUhw65wnAKssPjxrUMrm0VfdvYXpRYpgu9ReZgQ
T3O6PDlYfWFnaztG/aGhhcuU+js66znY4t1x6ByitX9ncmpmVUvHVTf9zXJ4oSbT
XdoCRaPS0OqVMW9Aux0jIVgOsFc53y5cN+iKKAPjM9jAKCvv3FZgNvBg8hy8ba9x
VpRAAD4C1cEww80XuPOgNhUz8q9piEgi/zCaWE62rWVPkIoA0cYpibXbgnFqoSmY
YvEvc3B/Uz/8ULiCZZAG0ffPQWQzX/JE6WYnEaf9G6hLDotjBCkLNgYV/Zbq9kfh
VsOvoqtEmO9wWs57AaAmR/NphK+azPRxsY/pohYTL4uaiOseKAnrOCPRUEuc4h4U
04eXprSjXYalpIYA8YoMzQpFjHosN6uvsn+CQhFMBVZ4va//qYGiLoNl4wSPYZLs
JKFJH+fS04pAXZtbjxNMMvjK5a3ZUkta9YAmlkt/2GHVY53IBZ11H1x71BGtp63g
gU+TY+nXKWPH6+fKoBLtNVYWxEb9jP71/3dH3g1vl0K7BM76IuoOrFQkzGxDe3Ww
8Yeye5Ys1iS2zi6/0BxREBW0pIFyNuKwDo4XahyJH0cvr8VH5Gu0qn0u5EDcFyY+
oFpfoA1hLYTP2EQHlggswmoOPWMCdifv9/4GQvembxUUhjRtAMmdeCXeoikMi/x3
K9WkwCcjaModlgq6/HrtlE05TE1ZR5idp23/cfH4T+jj0DcLoCGmUKx/NfOLEpEl
W/Ex10yULegoMAZabA7xnMEhyBd2Ydv3g6Uq5paItBK63OpXJAWmPs375/b81uj4
JnAOXQnIqVLK887jUFudr5VJD0TB1ICDT4nT43LpEX1PMt2XTr6LecFGeTBw764L
owJzOTBQPVm99/8Gq+53vZsXQY2Uaz/2m87/TxMEzt2UBmmLL48gGHtr+P6l2qHa
1OaNtXjpWkZoo5sBI3lKkm0WTv9t+Pwiiu64WCrylNB9CTNHOF+v5XQtZj2gjv19
fAg20JasGMGAdxfkTl6vdRhk8xFYkHSIpcOMGNtc9AR1wnBqJR1e+lbAW6apoyl2
FqvZ5v83RASzxEWlg5PA40NFppVgCEVXy3GT9aJTRhMF0PBupySJX/NHpxkM4ZeF
1uR7RY6Lu/ex5XDgGodeHipCNjDURqhxrO6uKzqGn/oWGEdzVSguv4+4Zh75jidB
2EQPOFGz16zRn9w7qUuYgldjYrvT/bCPdJ5hmlwzYNlgwxDBcZwvyHuq5EvOWKm0
leKtfIue0BzSs62vfCm3LxtRodfrskzIzANM/Ek7kKtxhLATDN4A4SF4KR1sWK8O
KZKrdR4Vpj3Y/ER4xorol+jdtZQZom/cOLx3uMvOi5agasXqACE7KJf52NbUoMdo
jSJBcMBbeeajlI/XRRxP12zEKJ0FHIsJZf9CNmwAtDf4/EZzGrvVDqn9zK9oh+U8
ULJe6otP1bLH1r9acKmuUhLycpdO4t09z38pf9Kfh259iS4DR9HDBDEpz/i3tPVx
iqOL/gifJ2LlH3qFCnPQsFTrBxpUHIhgLftNJlVzA8dowG9HUVzfzDBKwPO2tCWQ
HPBBiJ+3ZQvQ8Q/VG9xMoXN6y/kLnJ0/9+ALdBg4Kw8jd0f6pnN1C0F5pi0c4NKk
o0mS4P86QYjMk2SY47dhaRkq1QZG3Ji5cDYxLBtUUfcj9IQOdtfgorYEsers9auF
an/0l/sZdKBmbv+0UaJSRZ2KMkkbowzYwwB9vXTu+3sV9m/3KnThyOvy4OPrutwJ
yTx/Oy8rIgZrY7qQWQ14sFpJdRrBtP8ri4WaqIDIaBb4ryJauaNGH0BXIxe78Poj
bbZZA53LAq3q6vgbyB9UcLDkqv89iGmjlvtOwrbkETXeeAnOJVxBIv2wVRbBr6um
Em2oYA32lrG8qdEn9iKZiIh1ID4CXEJdw1lB9g0eoSakNwzZ0F+hTyP1rOvXQLPv
RdjVqv2fThKa8MJgUnlejNcRNMVG9DewC9pJ3UgCmU3h0coVAt7HJ6JuQ6cc0UXA
SmMPgEtS97vRjKPYK6f0Pmk8b0ugvBxtItpPJ2yqXAMgOOErFDqO7y/z+Wa4SLO+
Aj2AGqbV4R8/Ye4sYzlXPUsNZEivItmo0ppY6ZcnI5f5EgO5QRZDBpsfkdn+rs1U
8RsnZdCnM3Y67BAdTZfzsa46YZDKiWay1IpYyojfnk1shAXm76DsQ3vQG5RMSwuk
gkCFdAnURtwAVkgm6ogo1cQrW5E4DqrYdTJyi1e86v14yva0LWQRN8jZ4LlCv3kz
lTSnbE9T8346Kj6W3gesU24qpFT/o6ry7PeYwCn/17p0Ej0ihaf9mWB3oFQoa+RA
29TQBQQ9cCbne/oEg85XX0Xx1lFouIde4+4zYktejC12Kg2EkiVtgazpAcByV9XU
TYUh6YF1a4LryJyjs7nQMowL+npGOQkHvb62+pL0vvZaIPdavl0/nOagSvvFL5Xo
Jka3QiPRzRskHLjfbRWO4nNFQfInN+81zkcUALgb8Ii7T5WT0TwBnMKLGYah0W0L
zRtZFw1zftleQAQrOSnBqEcC90zKsb3d9/PrJOvmxG6UoZBZP4JU91RLUgTrBe1w
0e3X5mRWsF9e1gKJt7biMEJCEGG390zuoqBkIad6IRfMq5QTFVbv+FgeN6D8ODan
EK5Pi+E4VgU1maf0i69wTtFMNsKzdXq5oVmpLf3TL6dnBEN5YdmdVLN5lastulls
/euAk7Waxx9wvJj7MgOIrddrniiw+nNNxvQ/inENujkd203dQ3PTu4PIppaXgrrQ
KxH4w2HF35Za/36QKDx1b+J0IyCyt32X6wcH2+qOY/YJFc8OgQSr2MOuW10FjKBE
JRSpQxhCvywlDlBzaC7gRAzTXZyk2BBKtlCutaU6fE1HfdY2Y+RahYellMjq8o4Q
8ymMjSWXuF6LZaaPQv6UELkaHSyl0xwK1IcpLMLVg0XwVRP4nyrW4vmG18TbvhpM
UaQxlb1MCBdf/LmkEK1T7+gf5ZAkorTY/aMHAa6j/9TWmOrHvOUJvTX5rt7ghmWz
m+yFVc/V46CSi961ubAVcD6oq6oV0ebhKin5ivQR+skbhWNUxSCyjBNSkhFT7IgE
BbJNhwdCmPItqXUGTVhfZL7Ssrt802OwBr+4PJATZRAgsOim83dxDVFzGFyhXDbm
IJ7inX/PGUZcWx8ne4Veiho3JE4VrxkG6MIi9Xmd8ZmbKfX3haMVXQMAk8YBfIqf
4q5U4q9sWMsoNE5CPFJK14DTIQwDxwcWMZc2QXDJ+c/EWb8Nvwv5PdH+BBGdRI6q
4wapR75GIMlGy6h90/1kSeafUr2F/p+zmokQjwANshPms2yzjdwORtnZaApyETc9
yCGl6BDZ5bhsi3XbVNPPNoaCNrQx+aNd7cZNsD6nM7bIgpwSxXy9VkiR/wSinF2l
vEUvcVxOxi9nj4t3EksGwpYLulEhkKt6Y4sQ8FzvAX+FFZnAsQXltd2TMt8Z5fF5
HYfUmImNthVsqBihQ8VHeEib9mH+ecaqlh8ASEq4+YFF5oLQHs7m802ZT5xrNXuT
attGgO1i5yEi1qShczd83O/PMBXWEDpU2Tg4/IMBWmhXtEkH76pdHMWfKedzmgOw
UvmDLyZKgXfk9R99YOc7Kvlo8B6KYbMNIELQDT7sqCJIe0w/DlpqsCAYb1wt1v2W
pZ90P53qV7bWYXoTppfzoRoy0NvfgIam6LNROrGQc/qcnFJr5sUYt+cFGURsqYzn
e6zLh+Mmbbr5cg28aS/nf3R2M0p5PjtycnvScU/O520qFK1EU9CK4r4oh9qYcdvo
M7prIf0RX1GXnBhJyWLW4PXsPBRX00pjxT6lR/h7wYfnd7sOez0+h6WURLMtpYTr
FaWWlaXesgrWPUY2FxdYK4+YWUqEWuHKbvIEdkSHyuXMy/2eKRDmLXajn5UH6EYB
1bj4FdfVQq2agh6h6BjRuUtnyS7I/x35ew7ym/MyGqUmoTAG1dvWPRmq0YbsR5km
szeAuQbE2X5XNJNSp9aSSV/0wFqXuVdqDri7beJ476nz0H6UyTeNea9c4aqWyePK
V5xrWXjbtoZhM+eyuvk70LO2dXeTAbt+KM9Ma1NBeKVK9DgSQvBomCoGDtUPKKIA
5sjPxj1sh/n+GOu5vH9dMjuLDLCNt0mXutZs8HwXjZBc9ysCSvaw4gWvMGv1Jpn+
nhhOr9QQYdXJ44By+fvgPwhodWsQImDQCLhRTORr45zCDTmfEGxHXpcVOa+C+q4R
6BluOyXnB5+Bo2LKCxZqxwjcbSMvvBVMdFFmH2fepToX37DaWSsZRrbUO4poAwVg
D9jQSwpkOqigu/Iv3tM71WBJO3yBys4EVyBg/JGuSk8Tew0xg8FKF5Ki94WXJ5Vo
tp+hz+EhCvIR6B0ltQW0CcV2NP77wXIfTCaXkNk1L0TU5bcAQBgZbv4dVpMsKSUz
kSYU6wvH97+fTLhvu3C7LU/XcjUynXPJQwqD6KO/rxkP/udoHrzmRW8VA/3lVnen
v51s2q3HdmP0vHOfu8wjN+1ujBCAD0fXgFCCMVmcLZME+qm6MqT06cIOncPXCmps
p0saRhAT0atn7cIeHJ3h3DniKda5IZDd2KewGVQfETjL1d7tgCTHYFY3NiycggeE
vOKKBq3cYci0d9v6bn9eXbIpOR43cgGx/IFhyvLwFhQNlK9N4pdKSytYYzIt30N6
x5HxyM0T7tHV2jQ0M5FUQVB/XNwyJnznh7SLzyE1lmdEW94QNWNpZ1jj5tjzX/ES
hKvEaeKX/EOJVwPHngznw3ZHcMOLPi/nkYhGOz3gOhI6r9V75imjqNsmagK7J3zF
InrELa8u3L1P2DFrLL7i+65gTP52N1kNIIVU9ROaqRVzVzEO/FRK4YTNUYHKJzgY
tqnglmVOfrUrCwQqJyJ9jGbQeeBCq84robLdQeKVY2/xDODtDly7QzuP//51rDhm
5hugRmH+57K8GXYi7maYBNOp3lY+pBvk3cOkaWqQRiImAQnJQtp9Y8UqfDXC/rBK
Lqna2z9Pi76+H7rC6UW+KR6doNTDRcDYD3HSU223VKQZRIoc5j5Eq+uaEoA16M/Y
52F5FgbmqPE/gDI2SqtHvFD3k1jEC7myGwSra3ft9//0jSjJuBtIgBUrsPo0/9bl
U6E1sSaeayj2eHvVPtPS9ADmZKHf18aQzlEgHSFVqYbllusxWZ+5KTeBkQ/T2trm
RfeR+l5tWP1+Gmb6P+A7cDsF958lctJGZntcmmkKTzci00pYK7abnEYF/ELa3q/c
DgZcB74vd8tJxRWwUsyIRGvBO4csWkQ9egamS/W5hFEdrbMVsuMaGC+1+IybrTvQ
4Vg1gqUYy5pMAAYLaLMNJNi9BE+Sp3KTisvNHscqqrrbzMXNuTiQEnoUPLgwT83H
sRE7Pljo2kXizldyGFA1wC6fw/GxpeCHOp/Le1cDfehqfg/bsoIGjLmuA91Ij6be
oMG+o4hPcqo+wzzOmQ39lFqL0J4PWvTbLOO5ancX+a8EvNuKhLV2bfTzYw60DRrd
CgbOROf2XHENYxKqrH5svGlysS8ROAPMEOQAl6m9Xo82x7T/N1Wum+xbEM7YgDHK
p4q94Sx9SJBIM1UpVdVQ+hCJIJijKo/MeGub3KgYLSJAhmuwgCNBBqGMl0Nh6lV3
y6rZaRWmGZwJAQRE7X5dr/zyipEs3YJfKPLFz9naPJBAbzzQvcKOiT+ntKtwPiS1
NBW80FAOeQMafqt3RMI8Moid6/S9cb2yfreG7/ijL+D1bwq47k9whoI7RegbWfPE
3mJY/TB5+hmuzI1dPZ1FrHoZ5uPp0TRDVznieDkXM5g7GW3zb52CAwqmGuDyBknb
exB762ahlFjX2R+ReEu0dFrOQAl8pj3PSfd3vKhBkS+SUvxccNQsgljNAy/rbFdu
IC+pD8yEJSr1M98ceasXLNv6szFszuT8eZcsbTLXVXVt+8kREXKDP2Zp8Na6ibXn
mxb8JUX50VlqEIxszZCpYtmTvfmaHZHo08PJZnDJx3a6LLRz23l44oqD6gY/M+7g
30yYax4KjqPcIKA+ldbGi0eUKrlYPUpaWS8zWx0R3o30RYB6PE76yJ9Nl16NFI+x
bFTLCRKxJc7zaICrZwK/tqjs3r8J1yA2xSB/e2Tqwnei51P8o+8QsTHnD68zjhW7
eYx3bqjJeoK+pLdcY+zi4ra3DPZixKrLcMc7UhKqXbQPRxexPci/LKmN1J6HLk8q
j+XibOLrOU7iYODtMHg52xrZr7F46SdyEy0pEPj8OYKGOINDA1Mtat8QYLo/krwc
UVn1XwKFf0kFdlIeFVxf9gvyhAcICvzmFDL2YMNDFCygChjG5+WBxqEOR6wZ4EBn
AYbTXDHG90YBtEys37TaEZ8FZeyLnUtmFhd2gmjGOQOq/HRshzsD8XlimRXutJLd
uJ6AzxHSPEjAKebs0i50MsIhKi3bICc6KThs8dHM5Kl5TqTnt+p27++qLDK915+c
q/OF33J7oDoYflOLmCgTbp2bfPTa3XNgApXr9Yt1Dw4NDPhcUW3fYRwZ728UZkHs
A3/GYMbHDccbnPdDJXw4R6mldDMRltKNkHZtekJfD9smH4zU57WhC0v/AVAGBYWb
aY+Jm2kBwBOUnnMlbXIramoxxwSMJ8iKbbB9darFPjFn6D8wClxGHHtvFqej6AIx
5M3eSlAvS5YVpU4nznZxPi7KmvpUNcloABpchT8NWDpDtXBgUOkvFWDdCzJXv+UI
vgGRaU67fY5JeI/45QSDP2JGbIETeRarYYC3jmAXAwkA9pXKr//+sFrc2GCyJ2y/
w55UKiJyOY3vx4EGvkWqKiugA2oyyn1lIrvFQd+buNt2YFPlHJJGav9WHGo/Zm10
gmGbNtX8wYi5iinbQbFBslzsuGLO8VFSM9Pm8sVZxS8NIlOpsUKeh8ijD2QitH/c
6+BanFql3TyKCMAjgV/aXEufgcM1apSa7+mO+cQkKWGXsXVjXcSsuMMH9VgPFB9L
t3/YFL7OFO2qHyNYW1ccT3VA47/HIrGnFsfHHj/377KRFnNKUHtcrhlCIBYqV3xG
LDigMpyIF12DT2GvGn7ri8b+WOSheqo8b7+KFYhI771VWAL3q7ue4FN8Kn3vjMPY
HTFl2qpj0Bb26aOXRmhumbT6VyeEWAzLypA1ivDNaGYP/v86/r+U0BmwZhiMDE0Q
a0GRuqSe+McekduERRia9FySWpEmgvw8+It28yuYfDeP9lwgym07QuDaKOOJc9WJ
bN5Zb1AVbjAbk0FOac7oMUggBqGQKGjQYR+m7Qoos33SJdCCqa/yfd2FLkkkt1lK
OO5sCJcmIAhdO36vv1DnQ3D3WrFbBYTR91I9N2LSMEr44dThl0MVFu+8uskDSiVP
Szkdv5DBgR7ZyAsYm7glFjvzQdmcI9c3gxdMbN0hlQkR4jV3KRCFzgtxx/lSpJaK
+y3rm8/hSuakL91IxuRi2zrealyatjf4LwbAEABfvyRL/JFtV6J7nJayKZieSKYU
7W90LSw5dQBeMwjZlTuEEo9TAs9vWj/TfxXJO9Gv6J/UiNiegkH7r1Vf0UvsgRVX
D8CFj+rDg+TH8nt5erWboHMBixKP2DXvr3EIyK7Vp7IJqjpUgFMMsxrUOAhb1hpT
OHH5MJhIrEN1sltx9Mj27jcySohOWUIppZ7w70RBgWWe4hFOt5vLtFiwaN+N3Gd2
4fXADeNDngIcLT8gYLFlZ7cSEJZLoWTmw4Y0xxNZLnf0cpxACWb7Gwd/pZDk50Ss
oc11WNS4cJqjN+tzRHwm/St+pC7VcmSBtcwJELl+p7PpVHLAFsYF1fyyZxlLuP1Q
ijJOr/XYazqzA978BYQvEOw1xvngqhParSxtV47YQ6serU6DO1hnvRelO/Crt6pm
m69wXNiKTlLVoDNNHpUoSTOhne3sVzGA3TiazZzxe1D4q/lLwmMh0bTy+QCDk8KN
nJ8gLbGajYfEJDdganIHFXxgGv7ecpIf9wnH4rUEi8Dm2aZf66bwUtddzN4KzJNw
ZWOKG6hm2gYVsoaOIF7WsbK9FuhyxymkEUt1KAzsUs/y7YD25uWZ3v/j93gHW+CF
9ebvRH+SWFrEhmY6HOzFFwqzu/zDPgFfj8kevBqNSVwh+4vdUg7SW9qbnW2DKfPI
OJ4poW9jTVvrB3EP64IlAiLilNDFHkWsk568o5DDQJPWtufjTTrc3lCVDKZPdUnp
arYV6UlD3aGj6M8hgHqkrH3ZpqTE5ag5H/15v3x2lt2IqfN0jqbtjVVzefUxEYJD
n4sXNXM4DKI3M0xsK/WSvq5tSWy0L36Uhtn4nkIXyftqFgEgKb3GSwd3L1tm3TXB
KzUVFdGDg+yraoZdPJwX0g8+ejby0dXYNYn43rbU/A0rYx3wwAovLD8DxqjgZvlK
wqgGfPu4qAAQcBy7S1NjxJd9phcC/mMo0LvXZZHYB4GfKcaeMHcrXTgudzXhVDJL
WE3kGCH0Kq/5K2rE9ff7WsLNx+YHNG29Fp7SdqiIyXEHC9ezsBGldnTsupGdYvRP
AWyr1l6SRPYI71oEGyHppWarajZtL+0zzMl5IAS9l3co1A/FbZ1Em7GNrCW0umAW
S5cSKWhTsAySiZOaJmqzK7MANa0Qka81prD6uTiiHvTie2vh8IcSZZ+qnWw7WuYt
lFioreJ8GyflI3xezG9DQbb6EwV2xzgHm8ylHBFIaWJWciidfzt8JMQrxqCQj15V
7kCZ+gY+zJ62o2bsnPY6iSVSlVQQyxZoajP8SR9r1eO1HptNIEEPtACZk6L3RYP1
3YQ2x1T045cDo10RcGQRrk6O8+jWI1ug0Q5VwzwCOS4MYLxY2+5QdA6qG1CFtX4z
sInPDePVMIoLIgd/PO9HPvtRb3QG7uItdMJRBnidWUT5carcuTlF3h88MM4EsOV7
NwcA4m/iwt9uR6SwXAdRE9MqnyKpHMnXQ3Ut3L5MKhWImQ4jR+yiVQ10acCd6R0C
WbYtnH86ArLEECnX5iiIkeFW2Ejkc6PAcEV3FtH4N8KC0fm/UxKHLcsTrg98hM+A
7pqcwl/5XCl4p5059qIljsfqyL6Fc6omsUKHAkJkmnKTXP0RhzlADwnE8MF5PYTQ
0olsHkDRNuCX3N87HfP8GWFCYTjPSMwsFQgcRr7diCcSB2bwjOXpxdgpctO8gJ6D
PiCk/OihijaFAhen0dRLQCr+msNlW+9RLuT2S+cQCOLMoBKtFgphQixbi6/TJRUL
uTjzQciHbV7joVwsJ1yDzByNP8Z5E5WXF5J1T2vRHdkmP7Jds4BoqQHvC88zP5r3
VlXzEftxkKD57mgN5yW7swDZuaTQCU3HPVzOkEUIZqI2JKd6LeWk9Q8Rvyc0bgX1
2zJDIN2y6vEvEuqESTpc6qh/4q6VcrtkpDkCsnDt6w/vPlGP4ej3sZoD0OPYZtAp
j7O0ySaKvBMn2Uk5fH7S4AxrO89TelzEx2lr4foR6cvB0rcf/sm7r9qMvDeSFgXP
vTxdac/Nm08G87D0AvPSnLcF7oNvC/9WGlf88WdLF8t/MVYbOn0o/Kmanm77LB6D
NfQ8KAQJbfFTcDO7h4yRMtIPLCKoaoPoOH89Reu6x2gDtgyLgAo2lShkSaK6mTpa
hgaVjN1jAatu+/64nvFCLQQ97McmYcDWxrOKZwFoOo2mefRdS5xxw0jXarMy6Uug
6livEz7szOhx+vz8tTsJOgw9hzcQXmhI0IhyEceypPJMGXTOB+TH5lzcqcuq7qE2
j+sz9+rV3pwsfbSRJGgIc14EiTl2A12hne3YSwBwuaBrZmvEzcF5rSahYd5gc4ga
F38xkLDp2tHGJwybOMYG70zwB5k1/5VS+LBI0U6CCifMvXYiU27DUnwkzRsbX5EH
5gDQ2IhCZskpcrAz2f2JhBwyHCfWbSKJCBRrZfFkWVUNalH4dToW7aCO34VDFM/q
cSRf62BRVRcqHwgpS4uSp2wqn17pohMcJ2pMiS4yWCBKMjWh3Z3JrTtNUBDy7xLG
UQe37rf3wuuf41OaLNtekV38l8iYh+2ziWcoAA1ilCsGTWqrr0LMO9Lo4UMwltIR
mmAvMNfCb03dsuWzmIQUbWnI9ccE8rS1LQTc/xvYg3ZDNXQGRHr83jNbKxI1c2Kv
cJ1AfeUBc2wk/p97fSqepYzeT9l5MgaHr19pVF01QKdy2xpT8M3/T/VHN54Tp3kI
ZBnFwwmGZRSoN8TZL2uyjq2yn1zPZUvLBEwONjJWu9CI3rEwF7xP9lvPnrjvZYqc
1rKRNwyqdIAzlm26okQizVJP6up4FQmLcqjwAYhjDQnApiTCTADVgcrPVSJGwh7M
SjLfJdkHdGnvT+uAW2mE24bEmJ7zFTgyau1jBK+4UoylD2TjIx9HhW1TyfbXwKbn
XmY2CFwsYNEVLGPuQczPX6fSkjARMqzvCFzjXZU/X0DfAjl6F5kgfXzwLs8AO+bG
H2gLZ5G4c0vG67sxqexaX+GGhSndPSYuOKCRt2mbdm3+dWtxSkI5o5hsGJXtwvTm
ZfSKBvZiMdQnPS53O9C2N1qvlz21nTAQ3Blo18mz7wMMjjnJaJHkz/iZ7yrMB6yL
jH6STzwHt/W5ZqAtVaWdlZOZ2l8MUih8k2YJQR8Lya+msbO9RO/X2vZF3yTU+TQy
LN0F+u3TBuLlz3p2eYxw+KxL+Vug5asxYhFMhyuQVAY7YhCrtcha53iiczfKhaS7
t0QGpy7m645W5r2R+fA9PLgZ6/auu7mY7wa5e8d78lpuoP+vkd5ln7YDnql+/L53
ixCUiN9TTKhVqLLfNPUvkZSB2SNYG5Uv7Uqo1a3Ono4fh2TDGMfrUt/2vc57EMSB
HzuFAHloo1JHLha4IbyMx/G7q2DYqn8w3oGC/1pvajhlbcj8XywkK3QiILRaVctF
3XyXV1xYICMLRlbDqN3iMJZPP+nAqaKda8kwmnSOKANpv+494iINkcULt4SoAh1X
TKKa8BbsyiGfAwiXzWrvDdOSGpWUTeoHsuLMyZ1BkIFyEHF5cSxfKb5IAbOIP5Hs
qZt8dPEwGMJ8ncP0SJtMVoBN0KmmUMUhwgaFghOocazTTJqNZTjtp50nzQF7r8TB
YFJtHgjvBSP+mx85LZwSjS7Ehxt7MRlGZxgftAmoYoYyBO/UVTnmC/dDj4lKw36T
Fttt3ypxNIOxMrS9xl4L3lQHK16Q//zVfnLtUSb4NQTJpLwWBmEo4SwArEWXryUG
t3kPGFrjMwMhvwZP9Q2CZJAfPxlJqyHHudLTr7NWZmZeHUAkA/PgaxDTWWDRquZz
HWSVGXlzKnrTZesjcqUh5hUO1xiiyG9IU8GtFNR3GzJ/EUQ/X/rq9apocm/A+hBT
Yd2KcjsGFiTkMjj+yapvuYEdBU34Z8iyXRMVUT7xrQtJRnwSZL2oivSPowaUS/nS
8YW+O454toM/sZxwjqDHgevQosOymFydrJt3BuccuX4JF7b2TfvYHEnIdhsm4iiY
ofm4dCL8M2qO0D6B5sdMu5tcjJGwYsgvR0s5CB/ML2wyXw8jHUKCect/yUgnl42C
KyCquplWCcO001roip9NKZXAX0bIAQXsbXXl6oF0nGHCS9JJzWb73K17d6HZy/2A
gvyA//8O/M7GVQpwV25HUdhDGvZHOIj/Izlluf5krXCq3i+oTgq+0OrBM8mVBFyj
wZj83VtMICGWf7TMFIMKbFFOx+pdTN9zBA4V7tdD4yedRQIG0ALtru43LOxDYXk2
VwJovKhsPLVZ5Q9APENXzOJ1nbzYTYg/3j1+jVgFRgNbnVf/R0TxMZ17Eeb67vKh
xJDzBYPCX6GPtSl7ea/vaBWDAUj+n2QAnN6twi5pdi8UhZOs6cwqWCI7BNnwTSRQ
4p79jUYDeYimGTZe+XPM+eI9P6zHURaDiOktKv2IfRdCqoDttSshzoBKTHnUd3CA
b8GH/YbCpTJ1Xe5/V5bSCXhDoDfSGQdAMaSkfNwohhNx3nFaOl2OnfXErtkD4KWj
u6H7pWP68vK2EvIQWwvRstY2cV/inslO1xWPZ2AiubBo7aHWtxqBTaA3qxKcbSjA
a250y32l3akFs+dsAnpuqDwsRxp6tQgHPGOdcpEwrmarDHGHMwkF2rBcg50aa6Sj
XTs0ZD04ggwzg79G3lC0Qkb9o4s3ZWz//FR2tYUFILmXP7P+UwTaZSxi0Oh6J7bW
2xoQECJaCkx9BIhIsE0jKPhmoi0WgDlbaBFR8Q6kx+KLcgE8VEqQhRE87YLcqYHg
f5wjmZ9V50Mdnvqjj6/HlRGCwT1gMlVJVOIuhj/FS7j++Wk4+lEsY8fgtvWmlzje
rNczjYiQ8XWQGYuTiPHT4RQsQFkFfLd3I1j6VVD5r5r4Mea4j+H7i92jZuidcSDL
xYOLKgszLoCLvdh3a4tBCEbCYYKWiPIEn3qjzjB7g5mnJWWqyNM+IGgsuYi0vvrG
mQHXywjazboorXnHPXkgkZpelGDafbx15iD/vJF0VrUIsLJ0MqglUROPjCjXJepc
ffshxf+yBg1/9gUzB0p6uC63AQNMjHRpY8VgfgGaGQy9JqdiGdNnti8SpbEe9DBw
Gre4ZznGhY90pufRQ7TuZcQCqyERESFaSl3ZzqUfdBtf9YddIheWNp1TwFxY4V6T
SwQJLGPqzcjpznpzIDUuyniI6nj6SNUhHVHhYaviZhxWIDIXmpOlCySWOF+osZqr
ROaXaLeFM+qUhb1lDg1osytEquod0jBR6k0grgWc6WESLX1JXFGNCmwigircPqnJ
7gVxWlYiTkZKoyiIx/MBECRCx4PAUAxYcsVTgR3AhJMt/eJgPO0rJZRaPeWWyDJ8
xRErqLs1YbFPA1iyOpwlAT8RQeaohoCFzVF1K66YtUgUxZgxtDZufTuqZQia0tpQ
FbHGPu3sWldI8k442W7ulqBKvr/xMKeCnh2aIXS4DM/lGytfr/omOFsK3+if1Uqx
bsfRPwUVfuhSt3C0fzduDqwJM2mnWoHZiOsiISGle1eKWj5q/Edy6xmjR50ze0PX
RLqeGwoDabibH28hbTb2HncgJPytZINRV37wz8xn+fbbvNv6/6kCiwWmaOIX9Kib
LN0HiktrrfejiICC112x1wrVLDP1fmKp4o/0dFTZR70fSpfNyhRAaiiIVtri1iXo
j5QEyB+cl0gc4pR257KHmuA6zhrzL459VzBkYO/z2UfuJTBb4/qQ2uSgyMjB2LoE
s91f6FuvZ3Y7rx12/wgnpm44vtldaBRQzUF4B6nvDVJrxMlj17uNK/0aMLumuWAM
nJi1RLYUwVJl1BtN+rPRYEHKsMb3amZzs/VLaz+zlcYKyA1p4bFt9q7sQ3x3FQgp
Rp1KPihTJjWKQGOdGFoqGpOVreXQhrzZLh8b/UeKfO4r44CnuT4zz9dwoZIPUM1c
tz6G1tCgihzAYpHxormQVK0wESrwRjPMw2+Wpmsbjre6sqU4erfDNBorGEwxwods
/Dnbj6mfrMuiCe53Up9TaMWd4kAZ/T0u92tyLqsuMFAq3+B3U/luCXnRSSIWbKYc
ftfMmkKOvMDPtMwZQ8Hh8q3Tg0o6GdUk4LNDrkdVuyrmI1xRmHrZnFF3zm+TDZ9f
CyiEHjh/30krMd8hl6tDR7EiecE0bRVt5DJ0Jh85QlBMzMRnYQbSpMaELonfTF3y
eGJYcK0WJL8GjIjKU8r1oAnpv9l7p3yov2bXg9y9CATmzf74TwxjHZT20o6Z1zA9
d3ogNBh/J0rjg1RiNipXs2VDyH5nri1ydX4nY46hiBXe2KE+CHiaE8vmV/CJL1yE
fhCRn9I+QhgjIE6lA46ALVQGKisKGfXq/OxLRDeYmZ0TMQ0GJpthhxHh5HVFLWAt
nEvZS4OmJwn999+p/IkA2iy0+i0M0Oz0dRJyoAnQygghCQgj7Wm1aKXtlcv8edfa
ld0AYZuA4mzRWt+7rixJ8GR118J/ToJoiSYxzzbF4BPPBWpXhDjfhXapPua2XO4h
WYBXcmY6gqEVN9w5EjTnt5m+zhirpgQg8DMET9fDxmidu5NDqGcTgcaIZhOdzx0p
eRnJ5GY/sSARakOZcmRLOi/IzZ3P61G1ybb9jvp+RtN92z39bHMGq4Cx7ybmDs2Y
zPfrkL9t0zgldmihZaPAHVNNCTi5ZJifmt8X9CMtqm5YjXYd8M/oX5EBTmwl7qsT
HSi+rtTBkAzLCtNT1gHM/deHWEqEAWnGR6AGnIuc4MTCq2EmK14LMody6p6oEzKq
T07OXujgBR/TPrq1ptgVdbKZaaxVSkvRKN6jvLut8iMFX77nYullelyfKiHUpOyt
Z+R2jV3PnTnxds9HWnDPsKBLEpuz/PwaUv3H+T+WYVcCPQtyemxXYWs+IXr+Pxaj
VgYtOcwHzONZHaNVBXHiywnGJ2GSYRSeOHuKVbYnBNJ+760eIXpzkOK8g8wFREbv
KR5B+Hb5I17MqNu7p1dYkLx+D800Wtpql6ErJ4I1fKBURwv2OnCyL7uLbdIbIsb6
RC5kO4xg2UujvIzbN36dFu6igCCjojsEuXnnMHu1+uTyaCf4tgQHsmVsbCpl7UCq
eQrxFSbSQTM1yl+SHO/FktpU0W7rDl2tMvi/mSxL/TuSVEbQxAhI5a4PMvus1WVG
i4AQn0htnqsDCfegJvUemP2zMDABVHNboDRx0j1j05Fp4/u0/OJihLZi1nrKwE5c
m+Fg9Kk1Mo/Z70ocDzW+E+vHx4YjEup5AmctWl+/6s7Ucnyj3N3Le/rWyaGqzJ46
8mNoa2oSQsdaSnY67+22IFOELxNe0qor6pavLSZSuAtRa29bJ5F+noypBdcgVhrJ
nypaPoYmnyOa8d0nAxeIyVmYAWMbtO2ocebbfNbZCvFfhLwVX/OU838lNvTMyq1f
ptUrgQ9SWHeXFYzVIPFbP/Uufp49Ggl/HSF7647OirwSbQ8DlcVn2XaH7Mr3mKrI
GFMYWBpO2AXE4Yar4/HRXrxtC+zglnJeVQ5uMFPPmRLR9Szy0apDpiTdGmUF0nf5
qQDZB23Ujgnn4encdW2lR8cIaRntf1Zn2jKRX6pMruujcBupXVsmSqarXgDlQr2m
uo/pReTDZj/72htvYD0spGEXgilnDryMgZus3TEnX58Gbt7yZEWmV4/1YFs54c55
knMtk5MAkb+JOsiR6E15aQCgFWERe0rvofnkq76NB/P2bo/qrpzfncT1lY4tMzJa
ti95LVWeenvYKqq/37iDq+AfIY9z78de3JMSRb/3ZsAqHx7kDa+pEkUGLJEsQsb4
9fkKGv9xZvVk8xpvvuT0SENCiEgLSq/kzCQWZJvvVDF40uDBf8T+DSONZhiHxky8
0S2JXK839wNM99OPShjJVprQAXv1ZpGJ1w5ohdnKeB6BqUjFumajMZnNWRyRn5kQ
hLPqRF1mN6nduvMekJmoP3OrQOL/Kq8BY4WpFT0hnlz0clkORFHVPppk38u39xMd
N3qEzBJP8t4ZOX84wObdZqZGdPZXkWbRO8/q/g7uxQ5/o0FHEh1+39HP9Mk8LIz8
q1/Z5cSUTCluiW5wJQBqKpJKvgjTuEJfGPcgjzH/WTbKSvF1NjnpqaS4JC9Ozu1e
850J3l47P6Eog+j2+9Hg8LXEndbRzjIeQKEjh3OhMqXcv6qTl1KEXKbVuPKJbMW2
BjuzlOQTWHwFRJ8iPbU0T7MQSH80Ktb7S0q2PAIQol1mNoB94LL61wgIxKVbPEFi
ckdgl7X7nmnOKkzNugFFnq967V8iOcXnJqQYfvt6zqQMF4GlahLqqrYRCAk0um/C
rlAE6c5XlO5Zf9ZEsemnVrMdTQb/ADiYRhHbpl0zvKXcv2IpcItLhxtzWS1cXzs+
LP2hGvKoSBbLIwLAXx6VzLIM2Fi3PQrDxz9UBjbq9j9CvRKoKnuEh6VIdN6my4ff
H/0tJBtPgIephooA7d2Y7ZAdFoDAEBsq40RF+M0YGpL4pYEz0cZoMyULzcVDzll/
f5U9FnZOwGS7NnV1ULqJvBQVh8v4r2ImcHfWdbcBDtMyQ1KEKmWZNKX0+MyrOE/t
C1fAt+iLc5GZIaOY0D1CI7v4Sg0wxurxlkYUpAnujYSj9v7YcamJ8CQCivXqKyve
IGiu4n1qptMC/DWrlfzuPCLJ9f2k+9z4AUqkiCYzB53Xo340W942FGV1ga6Iy9b2
EE6ipw/qc5Lq/povH7v3cB+6yrvH+eVs5m4uZMmCqX01BphUjWz5XNUU9SLwlDvP
fjZDcZhqmqyL8uZitw00CcDI2LoVAD3XAVZxXq27LzWTxc5hLgMVcRNIOuKW++dQ
2b9ptUCvrKCr+QwyHooa+nfNu+KfRda9xPGLvXlz2tC3EikXR7/2sqblLyF2c/Je
DZc3sR0DJcA3Y5Cs8zyVCswTmZBn/mH3apFb0ZJu2xp4XX9FGX/rKlUMmy5dxf4i
jkQ3EYE0cBaL8bU9vN9vt9VJhkqZTli3veP8oliwjS0mY1VMYLu6wbyfnN6rQdE+
KLeHSBGHd22H4S6eUOykVVhOQNbM/lkABfEV5RTBLAvc20HosG8GEtQwDTfY2tIN
fywZIG4dK5jVpvJXw5SFL2sGBMwbVm+Nj+y24s92zSfZ1t1iW1Ftcbkyj/v/HDJM
UIDbGDjtkISA9aEP4Gno7ppQ6M+7qk1vf0baZmXK5bNXIMYmVX/OxaaYxqGjQYWs
EV6RtQlUDEaXQEuWguag8ATXL6fgDYlzz68lT2G38H0nWk0fbNPsreZgqGZIRpxU
PasFUMYqViM088WRWWKSzpzOK9vCJcNsxNf5TZiJ9OJNv6DyonMIF5tithDTaH+l
/bUhNWsffQLd/U/ykXE96NL9B+Ynco9BOiA2WnJY4VvD2kA+JZA4A83Br7FGBnkx
ZIgpfMlREzlydF9/L9tzb4ydPlUtC9O/ZMj2sLK0+DLGYQQZGvhCAbH1lcxqfT0y
+WkJugbNk+DxrFu9yHPoGc649GOqyumW0TyZqx2JWpXExYjwE2EqXcZvhTh3Z+fW
3zzfRB8KUXabC7Q8ty3OPGJb6DSYZsyTSWSFGvBfNqEUrX8YP1435BpE5BAMGulx
HL7qkVmLYbvi91ATLkBnYNREhJzBIZRoz5sUr+NnEi0PjbEZebm+a/vP+HiJ9PZt
cw93se+hTR95X/5jSYSi+oSPrIjeRBly5LDgyZ0Nj3v692fmG6bq+6CWlsEYbL1p
x6BKbi9cTGJ8npPLEKcaQ2ohRheZ41YFc7cS9CNjNnMtcFK2s/T3ntduNoBcnc+l
LpD1KvhR/ySkymsyjen5EvEO02U9MR2SiA0bf5EN2lembdfAR5a5Lyu9wPy5aOcL
Z2Dw6KWcUgaRg8fvNlLxH6bRiDggjQJQMFsGKSa+ng1l/mCSIvt5xQUE56zpxCN/
DAMZNobJC+s7WBV7MZlzBINtKwb2gzgqRyv3MtVmqbd5G8Di06hdGX/vn7Zq9jJP
WX6z6jV3WlzDppUHO6BDoVe0gFWwrzvL6R4PUDNpEOw/k4LjtXJoLQMVy7sdKBmw
ypetwaCmcldkpOpQtAqtV7mH2OWA1DVFiXeIExwHWp7cwPdlxw8Z8huaAyH9KiiK
tBl0INJifgbAWTl20aBzJdlh57VbrULZGuZIVplvmruK0Fv5Sa4J6fopUrey5ANA
E22Rt7K49TLDHLr3EVN1pp3m1NioO+SHS2TDh0MVTm+CBr/NeRGqnEs9g4hM12t1
0xdhd/3P3OxyjZHfb3DnItgDiq/+dim3VN2LaxBW6OugmrBgWe5oB9vGDUn01t1T
SSzdpoXEx4aRuxcHYScFZhV66qMcbljQQmw2VzURnNqgEqFIc3sM65EdMKq1TP5A
/Rr5+hTpBxDo4XeMHxgj/LisWSIwMnAb2AEM2+3Odi7GKjIxSIN4v+IwCF/1nIDx
CCKsUBOXIaV0DhW+C1hgd/wB5Z17MAgkFO/VtntpyKFQHt3KVcXqu8GHBLQ5EotW
srvabC/VGltOlouS6ij+W+X/CyCRgU71MjIW0qdkgZ/irGpZVZBf+G+pk83d605v
8gHjrk4RWB4ig9N4ttk4JG5WGL2lEr3k49aRFs0/eVvFlufBYZjifwhMUd/eIZ/D
wkNALvxtR0TsD/j1LIZXaXuStWHNqDZ4Nx+gk9J8gumHJq4Gy2TOPQiaGdYQFB02
2dS61Aa0Lx7lwugqIrmVmoT9DPjlxlvwlvEN479HiIDFL8NyswOBFBICftDwQkqt
rkvBi1mgrnCNu9Llr+y4MxN61iKFJmBj68uG2kw86yrmdNL2uFMbln/Mf5Ov+WG5
JGo4GRuzfBukIPPdkLaMPpFEVeLoIPYUanSLUpBFzOlujAp7jDLfd/fYdutR5wbK
jCxoS72jPoFXB6PwkHkCYhOvY6bvekKZaCD9RVanvjiE1Wkskw/V5IlOYCLdU8VF
4kqwW020HrTqkvJGC/JLV2D3cbhkRnJwYMGUX7+13uJ4xPrfPcJE5+xUUbBkVRzX
O42QcQS/ZiCibFYs6ytcwwrTBJUf1WcIyhek52FN9mJMPsZQLfB6nyXhny8C4Qor
luwkWKeQx/a3P7j3YNP6nazPJkLErVSMocyqYw7qJTbowwT6BOtBsZNgRwCxqo4C
D2fJgyX3RHIuH3/8Fqs/ijlSsZMa7+vUAYWmyTqH3lMEylWI3D2iiXSCq8nQJYHP
O8aScSnSK1PRewkvkDdEK6mHiHQlpNL2kPb+vWVhFowvknFj0qVsq9D+tXrWZq/j
jD0GQlVayUe2SHrrBad8e3JZ8YLJeUPJQpK26Ap4WLWE4J3Oo+r+L18RSO8bY3lM
943ZWI4tgxU+KEFDaNN6nlrb6Ij8wWpaNcDCwC6EWC5CDykVFJYX+HJXhryfaNO6
gSO4WiMHTnXb22n9POkm5osKmKnmkyHrMykiQXV8F7HtfyDOMKZYkZNn13WfcFzF
OQdO0r0wvaAk4T1VfrKWKVlTLVgXo9C27aj2ru7TmUK94pOBOevxDBvBX5XPkXLh
+dY4l0qbCW6R7P7S36pZCn9uFMFynI2vuInKxuf9mf5AvSAVn92sDlf9p9Bo9pKC
5F1la8SUVlpXl4hYtNmUoGkZyZOt30NX63TogdqTKmI+nCsN3LnziDUbRUty9DQ3
heLjqFdgTVHeSsiWzxNRgonnMvsq/yvVhikjz+j9lxgu1SGJ+bs4Mz3b8c71c4Qj
mnJJnxYvSkAC56zJzJBHiFHKPKvwaZ3kOaO3GKeOQE7O1dXFAKITpUhOfY+ufcYt
0h3w2xs+yPuH5pjYr/A8JTF1r6TyZC71xzXtIAMNNC+lKW7ujEsShEL/JxjSBLmc
RbdnefaEIm80e44bJkh0KnxOdNrIJm1ja61VRML+XzfWvdXFiWbhudsfArb4X4oL
l57ZqX4W/95GvriPW9uGCYhsgA/REKj1Tk3b2zRSR9ZpSbtdMsOxpvXA6Vxvf/Qh
jn/zcpi0VMaVZJl+C42MJHaROSXx0vN8jPzxhIXyH7CFkTvSpja7Q3y66O7E7Qhv
S8ruv4hDyeK0Q8Z4oG/M3/j//bSe+mJKm+LlOrSqqeqaCcRSTahKk4tI3pjKQMp9
ZHz/mwBdRKUEAd39tWkwUfAKYRvsSAQzOE6NedP7EAPb2DeWuIyCH8bAH3Pgjc6f
tNXLMuad8Cxzh9+9YpKA1bhcD4QpyIVEYvKVZBiIpPJouWXGf2nifexi3/tk+yuZ
zQ8YL/3++TdLLhvWyyUc+me7asRxXRucHxZphzOH1HQosMeQxBnZCiZm9qYjUecw
ASJWjqUzTSDgV3lzmL/5T7wCY1xRBgqaktt4OBsI++6vDn9+fXYoKGIvBvKZmULX
7YhLnbvwalERj9Ad3WkCAEX6kLKJYju1SR6C7jjvUN8tEYFVnAdUHbKuh9ChVVGL
tivcxAAW+he5iiphseA6T5+2QPVEWJtXI6xFEgR6KIR7MrS8SXprE0SK1QzKHD9H
N2cQHPXopsR6VFEtmq3aZbLXcG010E5shU6s1CWpICLqhf/YlTFPxpTkg1p62OzK
0awi5QuMlEfK3I16iX2DrEEVDUPO3R7dys3aZfkJwL9UJt67jW2/Tr8Nx+S77ib7
gC0YjS729ch40/B3KGvjc9aaV9Osw2VqZNxzVa9+o8ji3RuJW1pyOv3d2GkkhIPP
uT0YqqS0DYmJlF8ZOXZeE2Vx2GysUCZWaUcFlYyA7ygRwYSOl6n7z/XyPHE5A7kv
eXpW/PbFwwwFxcY6PSXwghROd5vqmJQtnhEbcuxeEgMyYdP61GyaBlB/TxeraYEI
L69jlWW/x7mbjYYt23OeU6uOi3+5JiqMWRr62eRc76flzOMYKPgX9G1M10vx3gHu
xUqlvxnawEaoFOQxncwn8U3rxCjMju7sCYv4N0NTAolznQCDJ93ES9wfFZ4PFzxF
lXCMCJ+USvmeLR77q9PkIytzxII+lwHHnEhCyxsUmpgHufhtgVXttXBzVAa9eLMp
D/2hdP9s4G5JDi5NimO+VM5lz3kHlRelwGDn4WT4FB67MedwpsyyBshvCLturdbO
jZEencvQf716l3Dk+28QLq8N8Q71lKJx1uhlxhuhl4VGBaVl0Z1u3JnJaZiC3Kzn
e7JdnvXf2SmPvUrLzH6sTMhYvUg+BELeLZHKq3IaSqFBlq1T8TD0+hrw7FIqZDTQ
FpOpZD1k//7urV8GtBsykbrrE6fXWOgOGNRIFhKf5+PJti46acFs7yAKlIniZpZF
9HxT2pP8lq/JOKfyeBFeVShBwL8RNFXXM71VlTWy2KCh1lkLfw6B5Cgi6vBY6PwG
grH+VSScXLmvBT0l/AuJbudukxb7b0L4Yx4ZxeiUX+/APMc3E7RNmLPZWNb2gFHJ
F95hfmH2cvIKWZSmaPZWWYMH46bUZC4OKRgq2Wj7+zBRLQLPmtkzmJKsyCr+Bzh0
5ZUOpDVQJe04HN6+n+LaWN8vzIHlbC6tNkbMDMq1D4/+/ykhkmCrwbxytwtM5/Ry
0uKNt60DgiF/4koMAxHH1hQdyswRigYxGsjPHvG/62lKnkVJkoYck2y6CNIf+RSm
Fazl6HYGs+K97c4GaMHPUDxSGTiAJ2KUQ4BoE0nqyE7xvo3jEIyDeJ1cwNjtTDwB
2oX2+DO5kLTn/Yev5xDGaJboV9LY1CQApynYEE5ZMq1InOt5bZ1KZKfNji9TMC6p
l2wX0J4HJmyi53osSwS9ZHtSwBXoMprOl6aUud8xVMteywFzKAq+2TTnWCcqMrdg
dAKDm8MveQglYyvS8jj7x1mfdBlGF1KLmUDyhWWSnwzXaB/QMLWNmKVsmsqNhrJz
fXUJyijkp/ujla3GKvb0iycy2BYbwmgyV9ohd9A/5za4Z857495BdiOEZ2aiV/q5
cVM+sqcf8WRrrwodF9iV0QU7PVkuZBKhn+XNZuluhK0eaJCO1hlXPht3+CL3t2tN
pd//QOi8IqJoOBFwwP551k7qIGhgRdiZsHfhQBMvmHAX/7tX/v5DRyO/HXmS6E8U
U0N51caf3pGjRA7P4rIUwH7ukuQjzIUHaFc1H3R7h9jjFEt5t3k066Eecy5eK65f
vR+D88rmUDHXvl76Lk26Ip7usFVXpsONBzgHFm20oKYDczo8gSdazDuqE7oXDU4P
VIhCxuHm2jDxE7H9cJzfezZPYsnPRBGO529zQi5FpAehm+upp0eLGcqJz6IlPyTA
a2SWnNNfX79AsGzCfvr54SYxE9q7jYBcQzI/kQtLXB9EZv+aCEpatlV8dO6kag3T
Kci70+UwMxT4v67fmY/+PRBnZkBCm55WZUBsJfjYjKqNs1jWLmq1FhbM2pNFdpt/
tOioVE0p10YJ8PTAdXRSPe0CQ3gs25/EAxnnxhb/jfDYabLSoNO5Aqh+4OfAZ45e
HIg4D06P+47GjI5WbkVqgN7ck7fKUlV9hHYI3U6m2jkUTGcmzmZ3nBYQx0Y/dCTH
cpLbWeJ61ZGwEETRBzfNPHeILvIZ4/h4vDoYemT89qFYn+awiuWJP/fOYKv3fU/2
ZR+kahu/ogrNnsy2kGAwkZqb8pLqli63xPkml0gvFNDjCDmf+pos6QZFxYSK+HXO
DULqGIOKu+88r9aa3FYofPgPPqgc6Ma6aLSVw+AXML168aLrJX83iRX//+TH42rH
opRDzH9WUymdUy/Yyh2bQth0c3/EXV5kdUrRi2BPhibgnaZP22HaztdrZXWG1Jcx
M8YMfO8Y2KOJcUGHIo7rydL2kbZIbNGndMtDRHBRc+SzWGlvQP8QXguuYgcB7QXC
/+GbmTMOTU3k6Dqay46k2otijmc0UUqqhae0f5EU8qhdq422cT4lbqMDN2j8SW76
DZMoF0rEiKMxJUOqvMhjVpmcdFKdj5RBkem/7wtnYkGYzeG9HtWZUVJ7KuUAULyp
cUzzEqV2XBqXH5k+vyjX0NV3qXN4q30DCbmqOCzWSDavZWx9sP9RyCpEWtXNDjop
sfYvymO49O+OeC4Q127gV3TJ/OEccmdvVh6uBYwnLlfnoSlRVxRP3iMEkwZlrhkn
0gHwP238sVSig7S0x1FzjG4Rw+e3OM74duJnBGfWO5KejqeHzttGuSfUW/waP3G2
XA8Z2b9Y3Bg/57P6g7pP8q+XEcm96O2DJU5avNqRoGtXlXF0e1o8Cun9GTNSuzAO
a7ej1u+g8KdHyNPT1wpAHVBe9uogcf6xzjgUe1SSiDClGYREnT2HreUVuGaUlEOh
fyDvuggkGC867zhwSQOdyNEz3utn5wjt+O5B+yu4RloNN/xo1ljAqe3USkGljTmS
VtN85yG20M2D1b7BN52q9saZL8C1Vi0oPt3pfemQ/emUEKkxHwx60AeSv56wAts9
jjOaVEVhKoAv2WKnZZgvumUCDcnnqhz3WTbZG5SrVY2S11nROR2yRhyJEl3d4B/6
bvXKo+kq9XBSUJ4NYXYEgQVALSsvfl276n8GJNVKTQ+paZWmHZqNxXYSY8JOXdwq
MUN7iVubJ+7+eaXtg7RD2QAgOiFz7rCioXjIXhdh2hdlXZ8Xray82V8cuy+/eqHp
QWcN+CK8NbDLTOnDDNxchTkLgcPOgVqfIkRtsfcG7vHTLeDklSnl20JibAcUr51y
/5ygL7M2lByAq5XaUZn2yRNAExrO85S8/7+cHpqliDZP6Z2Bxs2ABRZif4oK/JB1
u7mrfQV3UtHv8DJ2FsMyK0tEwyzrTulJLW2oGhyTGwCE7V1stcekily5HKk7Scp7
0kf9LGnUnuORiF6Axm+EbOIQYkZz5FWzpVxJUVrKL3GCo9cBvMJcN3nICh0Dunwt
uJ7vo+l0KZEqHtc1c3u6vTjYbae+Ftg5pKwhOueqAlKdgkbdPBy73Ly6fhDxCZc+
LeCxQHV/JwTeHvntHULM4R/1m2CaEPB/phYyLNdaGPuUMeuI9N55+R+9kKO+CTYy
0px0/gcj0I3Xf+stLe0GoZ555a2hUlGvTO5eivnH+sWLD8RE39BLJzfOjCf/ZxY3
Z2o9QulaPgByMbQkGBE14F5996Ci5nxtEWteY50zy/obP0Ceo1B7LpVFHqwy6zb9
R+qV9T8t1MTnd1Xpq6iO0B2TERtjCB4AwQqsv0rPt2TfpSznyhv/5dUGupMzjq2w
PJhFDXgPP2gnUCOQpnzkWKf2WILAn6ieaERtwexpJe8CeX+1h36TlnzA5z016nvf
FTSGpm8jNtySzpyBJAEhBmNUT/mhv+yEdu0if1tsKSdQ8AuvIhZoAeVS63srfBeB
qIg0wCJASw2GWISrtIkI7RgYBBb3zYVGmsXC3aI9Qsv3QO++sN3NWPAJfM/QCrSn
7yrevN1/DhGe66DS7UN/1hmmjkMcC58ETC8R8vStdV+lHPDVwrqizJPdQGXdwH1B
2c58wx1sZ87F7nKaR8GnDURb0/RZvKZnXZA/yAXKX6SPLqO9G3befzVcu5GZbGCT
XDIf0d1ScZ3ihy2FeuwvSbrIFI8mkJjU7zclHB3bV8nenBBU9UajL0kAEsLiBiDM
liiauDZvZNJuGjb/MBSL3icYp+1dHXJG2pDKmgpkx1aI6vg2qrQqMEUMsfrvSDQs
H80fiFHcGZIn3e8BK3ARSaAoNTrjdOZU+JUhBbIshy/waIUo9zEwl9p42SnaTrxB
dwzy0MaawfK5igRdWXPrsEsBoQv7BFbPiWcvWIVZ0i8lXJcLnUvajKAb/VW2dKh5
A08kaSedO5pX6l7U6xjHZto8zAmCCNeLfd5sMb4sJrXVf0K3rG4BWw1zJTcKYiOp
vDf8sJkDab3za5AFBg8P7yfjcUpP5hG8o6FmfX950zFr9HUgKoaxKw+6lHx1DtBn
5zHN4DOdk8LdWl0oFhT2byd4Ju0LYsXdqIkCj9qikFWx1MRLwLmcSQKjDxrcOPUc
bQ5mWciydU1869qy9lSdWw0VDYix/QIa63kVqECjPkToi5akf1bqwLg7ND+tMYGt
oq1gVj4SoqeEPWxlOAZImajEd1h1xZabZfKB4l1WsOnMkQcZVLzfEVNxcLlNlrPI
gg/HTTCPoI7dSBjxVf0tIwRVoVZ4og7UTzep2y/iCZHZgHqUS32LTtNvnM7JWtMQ
Ie2aC2g/APpGXDNOXGVvZGSKqB9yMR6qT5dHSAy4+Bye+rxaVQoBWGDlIDd60hXD
/BGbrfCvLdaO3sDWB6kbMwq0BaY/WDFpka/VG6ZFPmiYK82Ab8qnEH4qirbuz8Pw
4UUg7FEddFjQQ/M+yvcdYbkpkofHshmTBD5/oQVGe6Kwe52npJ+4NTUFcYFlD/WF
vv6kMWFTOw64n/vcCiKZ1FpZjphrxbsMHC3DZPh4EdhSVWoGS837xXh45clq0J84
D2yKsPdwiz5o8D5QlW4mewaR7f5W9FqGn0szW8Gv7zriCDa1P2OaHkD/SdUhU3Ic
SGWrwvWK+/KKLQa/4LYFthQ4X+pyxjA3VWVUC6izoIAY/fNeMuLpxwavEJjtBWkX
DeF57Y168g/Yjj6+Kx0rJEWfFx92nu+ep3gLqdsy7NEh3RsyFXIKKhCcg02UkX6s
R313CGwIlqBlEnzUhCoiqFlqAJuvuiW3RokB+5wdI/MgQmdw3XEZ+xKbf8XU+NW1
JPtZGqy9YZnzfJr594U3opJ8q33L4q4Xhu7UbIVg5R9t2oQWuWPejYxbP4/RQwD6
7EZxaGiThyLgByWDoFPq+71iYLHjGCzOlQVdo5hayBwCOV0v001lEV5o7d2CPCxo
xIU+F0vfqVk3JWoHnZHpZNeQlDH4C3SOVqQZjfSvjXmo7OPbo8zVWxwZUNN0o7lz
g7YCi3LK35dW4QlefBrDelp9TyzB5BLuZXJsvqfaThv4v0+1cLGwVSv03bcShf+c
h2G/wLOqhDpnqwjdslzCBaNmw38APtIki2ZVCfmMc6jCmFFhQASTzaCtwvBn7KNJ
U9j479SoIFx7YqqdiKeGK/5CbYNjlDSMr3wNahLNVapjVi94gxJlyUGzw7TgA44G
YdUEJ8Rq2r969IFECREUqAxKlEOW97dXLTEI2siwvmuB4pKZkbXvfrG2YBrWli/9
mwz8T0G+bnPZz+vQ4aK6Jqu7t0H8mO2pP8JWEClK7HGYVHibQzHKaeLXgz/pBYo8
+IOhXzDQ/jsFVm8g1RFxNjC3k0GscOTbuZztW/JKI1TCCSWWrFpJvLLYqblHrD+M
vZwSpmKAoAFuq01BKIl5Gdb+QjawKaKkAJZdcSy1MHGxwE2jf0xDH9Ld2G3igpxp
69ttjjc7qJGxHnBBUpJ9He7LCn9i1X79LS1qvTxI/40lX8CZ+HcdKY+dfpyCsmo2
iDPBoTZQ4Y3PsYRiH0qjAd4v9sP4oZAUYwcxWEYHNCCWmC0+Gnsy6ODd/aOlnjkL
CrTSuvwfo2/9WQs8mPEVjlIEm1Lizwap5Z9SwMTXSlERRXT/nTkCUXLRBfJJyA7E
W07srr3kcVOjVmv2rvIZsre7Ef+EtyL1vcQjLxhMvfHLXiOQPHDqM3dilg5GW/fW
Ox7pmskZ7lCbyAz7PAa7Q7iBJ35792F2JlesaUiwmdvjMUtPA7A3Opye+HKWwhcj
YmOrsNyMtACj7ZpkW/W6yVCMZg8oHe2r512fWRY2dISJJ5YPJphfRXbb+Oix/6WH
lBtQ/hHgdqqHQslO0i7T/M6spOX9e3CA3yaD/xr5GvrQD9Br2ZRkUZa7TQC5JsBU
ffNW57cTsi1CWV/fY3X/TUHN7tirkBR9EP3dzPFOAiDIrlMFEhx7Ym6PcpvXJ0OZ
zWmetBFY0xW3gdV/iy3r6F9b8ijN40wqfBwJqs0AQlOp9WfWnXQ0759HaqKC6wNV
iyWQeSg7XJszepuByN5UhD3vY7w0LuRm/CA8556UscWkO49vBb1Q3ahlV7p/yH3x
aLaq73V6ep+cIj6UxEt5pCyLZCyCqbRkdn1boh9SeuAOsvKXpgQT2RvoMI9JnqsF
wOnz5xAEeUn34u+TQB2yMeOeNfig0cbH1SOE7dAi7+TXbnPI1cAdojCkq/oEiUy4
ILu2p+IPxEz7bZ8SSgS1igM4pd8yzcTkZyuGJZQ5Alq/djIdyqWtYS5KIH8mkd21
cgm0vwO1oUBk8wKEMVm0mNiR518RdXeFsbLHXrAIyR/vv307LR/sCW6emOHSlbm0
/XHSpGeWcKtgDpKmUOW2df+W3aOljVI53eTvt6yz97DIv3xJLjbTe0icBDkvqps0
8PPbAep/He9dJU9NdgeutF/uUSSZjbqX++aOwpc3Gj0Tut/RDySVIeZnO1cdpEYF
cUteih3AAHMdPrJ0sKm+objiJjIvgUmMD1D5FEJBM45EpcYLUFNudGTic2U4lg/4
5sWYoKo8Dbsi348RhH7CazGNFZ4L6x6wqi4xYYVLg1pR7uJ7+R+tvTxim/TJkbJP
81M5AQwQ1UZF0js2lA68mjQiJoeBI468ZEUxoTjZYhTAanRLKXWah3TwRAa5hDmo
mWr9W7bEgkxPG3WdVLJoSsesom3yj5ATYfKc+yHGwZlDHtyftzF0B66hRRbtebwV
2OnLZibnFLJ/fw5ZIgC3c+2U//PQI+9WFGE11U8tB/UcYQqHcTwNSXs3ZnhKVhdP
rcZyOy2SfwbL4UjBTZkI+WTx499XqEAn48bD+tbizQY/ATSI6pkgifEW9GaN6Mya
mekSl6f+s/Z5Yd7sAjWmvyiE+27uWXyb9bJ0WYhAWL9MRqCZY6Sy6H+bz1mY49wG
3XKVstIZMar/zlRc+em7h+ZuLtM1Ry1zFemVvXSECnTSGuc2Z+6tK6dUeLl2I05+
NK9U5BPaRVTY/IRXpKRu+ZifrOzoELKi6Nl8q4z6jSKw9nkPG0rQirh5nsEL4qs/
LlMwyTrNXJl29y0nSCYWPqh7O4VCS4kI4UbHlJrV1qRWq8wsMT/GYBqW7HAzkxpD
f7/wSDRYJiUpsDeugELZQoXatPSDyPcULlt3tgYct7/+IgkFPL3GXqft3dHO5fwu
wsG9YLOCjtIWdERsqE2GcMGS7BTT87rVPPTuiX7KNewwGBoVAUO0KPYnyzqR2z0/
ki0qmvxQTXqX22XCP8h+5jxwRYPYQps5EW4dQIItLWYqqeh5S1E40g2bH9zIlDQt
rx7ky5bbHxqVZbFBnCko4Jg52criob/w/UodeKf39wDSyMpyo7fjUU3/Lckk881j
AE+y1ztvLNrKNqwoLz4L/TI3hkrIlpN4K65zMfz2EscmKhbVY5hB3sZs9IawPYeC
g6I7r7rmlXJtCLww7Id2mK5vNDPd+4/3t6WZjf0ryDwhT7Kekhx1lxSrIhidwFXi
1Q//xGHebMFKtG76ErTodJUcqU/C58u3WALx2hqR1Lu7J1uq/2KndvKCKJTxbflg
Dro4AhbnL4XgLKSHZA0S1Yxs3qEQSKu+u09ZhOgGEG4qLZBnB1P5iR5YqDPgKGdC
dMHsNBATOsThyNlquObnOKB7iZuf8fephMiZ0+IT0rSDCigMIkEObeyVGNN2HWY0
jRP77XMaTTzzmAi/rafOiJTQIXG72+Dc074DkuAjgM07IUin6QcIT/wdzT8eyATT
/Fpwk/cj7UHMJ3jdONvRt2yV2gV3ofUe0wWXUSUHQW/ziyEvZUNnFhZuuTsMBafd
QT7RypeepbQ2e+EVIluEcQTOXXTlVfYBaAmJUdgAolkOD5Hx4Y+16hp5su5yCgpq
E5PGAvmfnmaSBHxGhWbkHPODyKEPfzTOhSaC/GV+jY9XAl93/XxJYdisaPMv4PpJ
u3+VUEYvhs1tWgXlfzNOJUqd5tBCqFqSxV0bviURfEXifYJgU8R3ivUS/bWMdFDr
6vUXwEy7Fig7zU9U8jhAR7Knz+TuMm1EgNjX3t6bQgiqij9g55KCaJoBLn3NzQBw
W48vUDyBZw0DJk3vassjIgSRSVdZBd8CfHKvo9aA9Akr/lN6vYJhb/RqRGxNSKEZ
JCIuywAiSWhF8o2sbzFRHvScJa+0othknmxW2N9UVxsZwHhvbWORBGzwmkUlAn8Z
AlMDvMrKqzoB5WEkcshJqNNPEnQxnGnlK01DG5HAvzPpX3oX1nL7M2q41lSieL5G
SaroGovX/IQQXin+HRqSbknBn1DBij3cBP3PsnLbdmh5vD6WUyoVEyNzKbQLUQI5
3xSxttWj5/wAlQ+bKGL1MQvqapUSxxoEvqOGusPaZuVcxM64oO00CjCRvIJgDn+e
r/+aox3lRbb0zC0X44NUh5VukyMMIEpkFlGNjU5xNYMS81IpQ9RAPShtfmh9b2fd
OoIpDNYCh97v47WjCCZZLtlMhYeySK9SezhgMvJkAZfu1l0oXDNveBW0jPQdk5jb
xPTa2pJdqA3aZ0LsKFJrJS/Wi/jwk69hilej0dbKRjvOf6a7NiVIvpSOffgfBKRW
qDTcEFDM3tT0tordNKl6lZnkK4arqNTJC4L7EQ2SwRzT33hdWnhz7VrhxLFNl7cH
GeYAlTzzYrYBGY1tLM7/q+R033aZm/gjD6PKS+BEvQR1baEZpPK3Z3uM5qnfy7rw
MVMRlHdZuyxEps1jQLyV6gzxJ1sqMTf+ahlC+Oyth5hn6s3XobaB3exbG4f+VicL
363kHp02DjXxAxzeDH+LcZvizI0TNg7ncdotkXsftH9B7pLOYxXczMtb4BZRAJCb
67q/jWg13OgcRNBDlKAXaqKOvWdM1hxOeDFmodeXLbnu4Bc2Hl+KiEF9eImBI81I
IeXSqLgI9d3VPGBDs4zO3qmhd7oO4JxzQ6yA8+TI0jOvt3fL2ch/YLZW+ON4unjO
XmOP/Z5hv22a153v0JWZD1hISdf6dO0QrOpwA2Ti3gZuAaEch9hVb2ISSct17FOt
5uHGw8hbPqCVvMGxJsq8ZGjKUSpOaDnf0MRDZZt3V3YG/CgJ05fLUQu2BAp8ECSH
LirvEJkHwtMdo5yUteSDqnGNzchxssYhpqlGYskgAAf2aQfhlb+PQLVYTs5M5CzR
Il58cbjI0vERA95JvwnfQv3be/rUhGAE0lM68SXIqkiS9wj1IQME/lCeVsM4n0Bc
mYMfABgGPdZWjo2qDs2eYWK/o+Iyhit/pfNJAnT6Q7xHRYIwk35ZSWY76frnrV+w
HPmLEmNP93UuDCMHUOcAdeMecqu5ZbLIezvj7HI0cMHlOFxaD1vB/pARjb376sEZ
37/cfwe0/KSllbfJ7iQstS43pQldMQgoZejzW4Ag347A7V4zcCGyMWdzFC1smwav
6Ah/lzo+W6sKs+XUbNvocLqkKwTdNs03ovu+5adHp0VJy2vnhH94NdYXswOq7dXB
nk6fqtsjsQcTcTjbtKvslzIal7tSRRmZ+hvTLtt6Nv8DfJ7M2PBINsaB+68B8F4s
FUdbVXIwBuce13LAe/75ULqQX+35j5yGIu3T1ZSNqD0Md3BjkVAP/sjKtbzgB2r7
ZMI5X9uhg6naovrdc/mxHhBjw3T4mtDyhrQkBu+AXNmqPiq4LzYFV2PWYcvewH2/
4YnFjKz36bzlNssAID2dLDMh+hlpTrXitdHOqdHWQB52GySkv4pY3rSzpN9eg0zb
k5Zr4Vf2ALb9h9AyK6uRW0REKzvUJQzZwdaIdoOL+72QznmZYSiUPSXZNQfmPYbt
qRIwUkVW1lVHp2RzXBksYImXtm/QiPYLePZwWkiEAYRZDoRJFkqe0Whnz0uiRyIy
M5kosLAd21EedPKaLa7HVuAwG+Rih3Re/s+y/+EFF/D22lspChIc/Q6qUp3iK3ki
LAUxvO8ANcLIEdbbIM+0X631+VGZP/uLFLcPb8Tu7nSKYMQIVM9NNUUZjWkCr+FL
ey+nNUzuZS6tAFJGWEeSaVZOu6YB+RNMqyRPDxW3fdjvna6Wf5qD/L0nAmjw7J3y
bu1jLmANv9C+Km8mEbiqrlQimkYEqHU54kcOhx057Jx36k8qXvr9JFoX7pXmCq2R
OJqyZ273Qkx0S1wSmyM9UaPAPRdeGCFL5oFzzcbsqqpvhjv9Q6q7SqegqGuuVBGr
FU/ohvhe9adhvhr2mYHl4nLyLSESxsBtoepadJPA2fmy22n4epo+3ijdXExA2WV4
+21gC7s4Kwn8WAce4t7CXBBd3o0NGWuMJO7t3gFNlVcwZWyWSbKX+jLlnsh4QAMR
DUZ8LGzgdwXOwjLYWfoLD2cexrHvMqDyqp1EwsSHxldIFTY3JNqB2Ok3lN3JJhcc
bc2sb+JmVW+pPGLVPSL2qLik/dapQIcDzdoKcth6VqXiAAxsffeIiXeXslATB4dD
DRWeY0HKk7A/wXzQ3lAKV3daH3OMlNg38invpJkZnVkywK+BPCoaCIkKw2dLv9AG
54fGbqlalJhS4E4YgNx/UE3HW8d/Y539z/lh9p5WhTGdmb/In2IAkiXXw4o/0s6Q
vE67QOBFx8iaumRAbtmC9fsERtr1eNDAaBND0l4TwP3ZOuSIXng+3I9W58jOgTib
sXrH7NjbrbLc/PvBWYxZL9u4yFZ+ec5ZAheVS2u71/9N+MyJ4uBPIA8NIQF2Be6Y
PIkylVT10lJW9XYffy4CKkhvpalYEGI7RYXfEQHmtS6egs8KJY0KwzdpWe5VpkPq
2V+Mc0k7uT3uPDdXzdTnBWOYmzukHeJREgbOylfzo9x3aO8fEA8VITXY34B/CjSL
sZnu08HEqjGhfRPYDrevDlVv/QG5+7GoSNuvPG1+oIxU4sKc3rBWGFlY+e7rHbAc
cpUg4uZE9fMPAOKNGrXCNGsw+UDqvjclmPeo53C/8HMSusSkedSbUxUuVgM7p0SY
lTDyKeRrrzWSYf10uaGcpEUlu8BpAx93UD4npO46cFIIgs0TmtC3HrrSkn1FqWIz
K/oaz2O1rAIweBwlycgMrZAe0t1J1C45V1OQKaI+pemdc1xJqACysqYiXBVGj2lL
L7rElQm4k96L6nS1jSd0ZgxJ0X3wq0JeBqxy3maxrJBTyHOA58guOZC/ZBnia9dd
86QQZjIEw9/weCK2dMrxtD3XMQWEtvhJKs9nmwG86woaV0KkK/aYuGDIZk2nNK4Q
PTa5JPpVMmIynCb+P2UQdw==
`pragma protect end_protected
